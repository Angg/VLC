

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
aEqvcre4Lyvq+Tt5PXDTwx71ktTXYMy4x/0E4dKe9BgxVOReq4m528LoaLIP6GW+fVGwy018LBOH
jm1+bivxEA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
QYrPCp2aMIlbBfuPNfY2dUNw4w+QKreq1bwTmXohDVK/xUEdLBItloqXSCGC7+jUg/Qb5I85f/Ah
KtJEJyCziwj6IUpMayW9odpLYrmaGSusKTx06OZfHHMO82exXNzudcAn72ELL03w+v3J7Rw16Yaz
qLJy0R/MjFA4OGOwuMs=


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
WY4Zr5cvsgwcIO/1W7ZGRcuOPxuu6EPbRD5e9/HsVO16X368aWkQR33DvIRaKE6mu6z2j0ahwjZs
reKraTCWpXPIX3kHEOQ4G+U8/pfBNAeLu+gHRaqilAs+vw9yv9whz81+ixVCKNNcRWQOTvo30pDu
skLTcm2m/QQjNLEpHtQ=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
m6613vAd4+Ikpmzvgk61cQ3LztOi3BEUS+a/u62stTAr62ac1zeSm3L/nrHzan4UzFg0iiv0fkQI
HlLvWFQnraEvQEyI3HNvXjW3i1zg2bQV+yu1q5XCIXhmGlzOkz2w70qM5ze4T5v98BsjMp4dYmMx
A5f4dpYgpZiFnTGLeMS7ck0fB2IZjiquePTdi7jgm/IG+qLBUBUT8dNiDp8GCdQcgG4HweV/m/jI
vG3z9EfAXam/6EPH8epbQzdWAIlMPFNElVQWIXYwEK7n7IkwPHcKKy8h8TIQQBgfI3+K1o6wVERE
QWtvGEQ9KskjsTu85uDfcWnHbHjSbT9CjOWhQQ==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
akC0NqgvB/U73AVdpjoyhrtNQqSO1F1f7/iM28U3ok7yrD2+mcT2y/A9xisbQ06qgSdVkeeZQ/fM
UEmZFdpeZP65dH8ladxkyOXEBZxMn5HBR6Cc/cxzHpMOCwyqreDrscOV//dRgt/fMDUdAzVx9xAF
S3wPRW/FXBzvZQSBlmnr30bFT/LL4Cj8vJGIP0+tX4O1SFvZ4wHGKlU5KqTKs8dVxLyBzSJGBQVb
pymfPPn1F6nJ0s221XFfFykuFYfHfCrSyu+wvMs87eFK5xuSJUkyXUmL+AeodntlACtqvxNeG53J
I6QuD4FQzVWl4npAqVztFXpihv43QWWvfcc+3g==


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
SbRxC27qGffCE5dqvP2lAKXlQLXs2E8yapa9AwWyA+r636Hw6fp2hwwnmJLYUQJzK+qMT7z/eV8Y
OxzIIxbpnjsdHYaEBRYqwROlVe6YwnZ7L6xK5KKxX53MhhFuBHhAxWp9i8Abwj6PqlCffSngelnZ
dnsX8SbNI4PN4MqYSBwgphTtKUTWu1vfLq7rTdNhmsL/7y528gK8mIQQ5SkILrzE8DHO+vA0WuoB
gDK05L8J22kNnh053JxW/y8ZxHFerifahlKocYNdeEgc4mj1EWLlwOKC3M4lBgZJ7fZnJl1veWSN
xU8ddBWIU09TNJJQCC3Tzn/0bh/v6jX6rkbLQw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1022992)
`protect data_block
A3Ou3c6bvypPqmHH+ijeb1RQBuGsBqS9fNKJna5DJ1rK8wKYUlaVV1rtKMcBtetFRX0nAVg6Z6Ko
YnqIgLFewmGozSrX3LP1NwgxF8xVyEvut3701tasjIFJbgJ+3jkI7M4VcHi0vocS2LvT1VlraAvt
ZTnXHcWrv7GhP7N4F0KHa5yshxL82w5nr4YmEl9vcEn0ulKY+2ZfGTkdD/caM7W7SVvFyqGUJp65
rNPI/YFuLDb5YJUOrLGqkKM9Z4W9kojJqH7WS0Sw0OhSqmEpuyHC2XE+ywdM+lwCVXdlSezibFXK
qHr1myTNnAI/L1+HsLuKnQpsMmuuvlws+IvVK3UlLryL+uljmqo+aiT1SnSAZctWz4sxZDDPs44Q
dFuu/acsMMTUIRCLzbq4n+t0Pbeel3bjjDmuJ9COMEJeGemB3bvs134ic6Rd1MjAq5SBWFiPqxVX
wsqYi6r1BliHgF1DJu6Nvb9ArTAMKehOOEOO7mU6HCGr7nEe9DHGQiwVhFuLwKRr/4bePEIDhbrs
0k/MCUWp7C6ZTLWtGBVIxvaryUGLMFnPK3QU/eiOMRIRQyoqhYKvK+lb628jwmJXeTH/wPq4+UBS
cW/h6Oas65932tq3syZT0Nd8AYPUF2BBDhtA7UuJuGMDY2NUrll/UynjR53pG65DBhjJqPM3kq1O
DqEzm0z6tK3bvUgkShe88cFcV7/gEn29+hIiky0givS/M50D6vFijAmj7+cO4nkLEgyl+EVGcfKK
OF0fAHzTTZV5lpsoHUo6R7uDKKLtSGXP6lEkorJvgB65UiXhy+Jo6nUeemzMbQ9fzMi2w1w3UYUz
Jo77SFg1a8e8XNxQkzO7nWWHRoNpZh7ibNHDeFyRQRnCt2rhnKzQKcVlPUt9lEQV4eOqc352u05z
JYu/iBjII+7TXjzjt7P0vXmZRb9Evm3yfLTwJwiZEFWpt5WNVhAVwC6Q/vfrWPJ9/Cpc24O7zalO
JPmayX+RASUv8Ct89KmjlcimyCDfBfFffFIj2yyikBAlujKs6MpyUEIaw1GCOMWWBjuh9E3kR/cV
LFLdtrHRQJty5enLi2Y6gjI0KfCoHJNXQsQCZiImbNHcuXZJVz7v1f6S76HNfmkIeJuHTC8NDj2t
QA2CzqBZyXkNuSZxFB9wS/l3JEpdYa4I0pzP7QladoSGdGcZvh+U7OzWMhzleFsnTqc/NkM4DePp
+cfltKbVvCpS0IdunoKQ0Tv5oBY3bGyyBTtfLQr97T5GwhwdVVrVf2m294gZTNHfGpyMrZOvxaQh
YFyQZ/v3is7TDLH7aFIMkZnyoN0F7CSA6XNaXn4cSZax5VUKaasMTo7Ix1oI8orxk2Kox/dlrFmS
hyftzOABEpnXJIdQwAvIy3ZUDyZW9M5nv00J5QxX1Kk+bpqoXXS9cESc0B3DenjpEoQlEPmrpMpt
II+d71FbUyKgKHVJxqj63wH7WlptYykLs4AwITPyLzUInkTVdl/qVQDtzmfWiERsreq75Y2SYvDk
f8ExEnpfs4OyuLUQGJNb3Q8m76wZCnlw1HJnY5f6132G6YBXrBdMR7FSlFQ5kDgKHm2C/l1luamd
xdtf4ev1seyWIzX82YmINNZCxNfkc0RODgYoZbielD1xfV+AA9u1jpRlp8m2StbaF7czY5Fn67me
ZGWCSoCqCEawYx2igFhELPmfnjhUy9z1T9tAmSHHJRWugAAUEHI3EK3iETrXAHWJPlZT3kp3jScj
wiFWrv+1jr2m2wSEEDU0e/WQbwTm3vcjnUJq2/zovJQY6IZyZOn1IHiV46w7hHpG4LARhblzvXLg
jtEX4A16VoGH8oALXvT9OfZjt6xgPNMLfuX6FedpWMSu/tzXHV4D9LoiT29+QjG98+v3xUfvwGFT
RHQtvcNhl43zU9TeIm2UWQDuFKvdlKfPY4NyhJrM21j0YLlIwsGslbxnlyCH92yVh8jearANk/LK
kPt9mnna77kBcpscqJ7qQQe/ngRGqh8TP6vHDCe44ZLgdGTsopYp0wqSbFjRspm0CuMk6D1Jv1aX
TfjSKaDYp0EMnfNxK+y3C8RXmY4dCU4AaAjwjxe73kD4cdmU7gTsq0XCtSmgnPVFnzojkRl0v1IZ
j7fn1eZ9iFtIUIEpJH2BrOToJvfo5lf7PZseIyQAYm/RnuKLAaSqs4vErvvG4GtfEhlrMeTWVwGM
beM2RRxQ7cgkvvgVASEQg28F5e7E5Od75pPAz/FdRlc9XwZboQfYaCx1Aih/auWIQ1qMFVu40exR
CupU89Zo6eGBSVpvMYFQGEbSN558KEnRzBFF2b6iT42wmyNXB52+8rMeutFLPnAxZ6bFR0q8BywG
ejMCB3z4/IyRs7GhYqck4LI+pA4q0TTpD//U1rJRXkdCzCMkxPOVbNLQPP5qnwWf9SICsWMGSJYa
n19ISBMy/hgkU/32Yrwzp9ixj6wyav3ulvBBYPT9qJ5wE5adOU3PejyZ1i9v7u7yiJ9lHlPhS8Mx
3AnuVZfN7B75/tr68KzRzgqgRT+RkMx8MDy/uyyUM4/0fYKitZDtxJ7gyXokmRZ99mK4rrwpWMom
yf3pqlE+CUB3jqvLTKbOTGulIqDJ+4MAaTWSV9CcdOymw2Nl3Vljl56OyqlSfUAkhnTbvtf/Rdbl
W2EtSFADKi+T4UXKD3F6TGMJG8ns+l/jzJyyFFgiTUqbT8x8wxc+vpsdR+YP2wdbCazwxS+PWCRY
YwyWksY11h4Q7HRzp21x88l1dQ5/Mif7kMvF4L2Ijb0EN42m9WfcdEnE6E/yhw6YByXoCM9AURtW
dwuPpBwwpVioETkM+4TJucLS67aRNSLFZzYjis1BCBGJ1ZDNbd670rvmhbAbCnbb/DFTIhvwaMZW
GdanNUJgtIYg8zqKaeiZsLd1fQAY5rWnNaOHEtoUpHCA2mZAhVYIgL/A2mQ9pfo1/p2UQhopwva7
Y6zhaHdH826tkYPigpMkPudpNsP/jjG6elDu83d3PPHwf64hzEj+NwOlNfQzMGg0CjUqIwens/S7
79kmzCf8urrzptP+znLrqB4WMlJWP4cTLjp76V7MxQrucEEGUn02EIRgpuGwxd1YlvLRfRgHVU2I
hYxWX2IQfMpZs9eiTA6mehKw6FBqYFzxWv6KBQEY46sAXSh7uJMEWQQKRqAWhmgzyjmjKuMRAwQU
INeul+tV62vhmQDcxnTgT8oGYrIxH5l8nmfjEXeTUTGYKdc/Ll2ifAdOx3nBNYrVQK/ZqsHrV4of
GQ0jpMHu7z+lH+6EqwRKHhGVUMuaOBpDShBjce3lmtncElXlWV7BqLWfwABNKFApCiI7irQCZT//
gUTtRSO5t7XknTTVgFZ8S6aO6mU/OXwhtjRB4n2c5fMzQhR/pGaoq3avsL96IG3ImcWtJmZblm+V
6vFuU+MIrN7uH7RUcOztLbhsS58koJb5mKb94Q2bcmhi5TOLaUzPvy0Ntfzz7TaDU9fVnqZtB7kQ
29ZIh7n6Vig6TF4LGUHLYbZNztbvte4qThqw956eeQoyKMF54A4QgmuLR8+s7i4NZjJ/oeFksbUn
pOdPSUK13cIRs8ia87Ed1gengX6cLunLqnAh6KvCnv9tKrnhsI5J8p/ievHrgZcvQiVT0pxX27mV
spZa2xT+RElIByGoBSOq/2qVYhjJ3Lim1Z0VvVuA0sEuAi23nDulSvtgacexV7T+H59VHEAgbLON
1ghpB+eMnCAJ9fJapjbAI1ULeTLC4t6yEFZgXVcZM1T1Q7DrojDSCk+80xbQ5GnMesMzgEo72ztA
OnL7SSBd9DmTxLtGMxaTgnXnDdqSuNIpDn6Ql+4whZ6j/kQC2OwKlWyXg4Ao9dW2m1uGj0OzUK8L
fAN4BOyVBCqbIa7jjWdei23MdDgPuGC0zag4axNiOuWvQ1ngtPwWv/Whc6xS//B8avfl7N9isTKI
+DcQ3/CectUbhmFcZNQDkJy7VLakZDBIx0kg2VF9e8/3yrkaXe6k1GP8MJhmLY5nVooeQQ+IZzj/
hdZoVtYgvim0pnegrxu9oVk/3SCpIx/qXpiTOfJcngio8AauEARk0GcUGjT6oDgzqSahQBrBtE29
yhwDNjxhJ6ap2gc3GTGkj/hUEsPdikylQKrAQJ8wh66fIiWFKsMqqxYUrGgHiQVHFhybKOpznk74
0NfAnsAtg+vmJJjytPB91d266YY22GEnuzAxVjtV2/CYxIyRrR7cZQ4cziBx6hiuJAOoXuuFxZm+
Oyycj2x09/1uDVsBn5Hn2Vixdi73AvX/e98C1fydRvL3DWU7gfyV3Gqsfykkrh1j6afok6GQ63kH
Rt50dvY5EYx34ofwOF6nvJZg9lWrHpBg8PB3bk+oLSsxpWlSRoddsSXvNfCGll8HPUr1OR/V0qK2
I1gyE3JmH8Cul6advpgCj1wJDAZjBF/6lwTwJaNXF87/bFJno0EZurDI9O2UsZMmloam5FIKqY3l
kkCOpKFqX7TmlgzdS7AEg0ce1OayiPAG6GtMnI+kvZUcys8FJutlvLQA80bLIhQ+r7f6H37nZo9r
f3UANFXwFQRRcpFYwH876N9dpNWZp+7iGrh4roC3R0PrSztmVAiz5rCEC4JD8Ziv7dAaHgsSm0JG
hMsSv771LnALrwmLLwLojl7yeNuS6K5E+NCRVMhgj5kKMALx1/DMsyv5Q4nJKNKtW0Arvpahd1eB
iAkhUBUoGIee+mEoRgugK7uvtQ4vJnyxRb+aZWBWjlrNLEVN4O9RVJX3lSjtQ5Voojc2x3n5/aLn
wh/pZA6yEt1St+Cioc5Epx8OceXTSKM+g0nV+CyLeTKDAbjOkcG415GOvX8v/fM8lTTgxkAxpPvY
qwSL5yBq0gH74Ck3EPhFfuOwSC9+RpcEeXAMcNvkbOVltFfQFN57HI0A+ps0kSMpGC8tlyJqOnze
OuajQQS3/uzkUCuqVX1ajZDWLVmmyvy4MbT53IW74vtzPGiw0P5JrCHr0T2Ffs6QolwnIFBYeNdL
RkgljHHl3+u3wu/QOGpxfw755BrezF3yUlKX4bXWwNyEGnqCutM+0j2rdwnrKOXY2JirXJY2fVP9
yWptvakSOE7cnLu/ubbPgvEZCrHk4X8T2wahhRVPjmIdfWEUIyNnLUAjjmTdPpHmfkKdm0t038Zc
51XTH43Bv5sUl5ur8WIJ/NHzT70xh/3dafoi0H3rNe0+w143uh24m6VKWJXpRL0KknZ8H1FmMpPD
UWStyM1TBeTYyCAjJq7OEpIZ73cO/FLyfI+7nOWQta24mFk0eTtg+q9k1WajCCMpPtFtZig3s/gt
XmR5nlPZze5NP4f04wQ5nIV27dj/dm5jTZXU8pk1gz/Pn4U0FqDnB3mYK/R7LkS8nkqTOAZsdt4j
F5w5uSu1Fn9c5YTVwGuriP9DDib3iNPEAg+JVLftYN3FiazqJraBPYV0S4SlQbxxfNt29u3nCj1g
GfYbc7uKHbR4erUQC5RFlzTk9fG5nfAqZ6vAknDuYQ6RtL9ZSNQ2vOoM/gofWWe9F6baTQChhLUi
MgT0oBf/Zvu8RbvPGR783mBgiMcQOzr8A1DQoFjDpJyd/AwWttYyoBrCKng5c3+CQ7daqVrgjDw5
gSTusLCQdZdICY9QmmUnqZ2wEnyqHur0C8Pwag+MMbMX4wzhUFyldWvmxYlGG9KIetMYn/pWyikh
pr3Jm4EYs+6JOTuFvSwKR2mbPiiZ4pBZOaD+YSY8eq/B8Usv6ZDEGFtHfTxhV5JlAgWDuZiP+sp/
Dcx3K4VoZNQVmzFS7t3DZJRLYUBFMh0TheDe4UXKSd+bYa/GHQnF7HoRjMQejQ45mBBu7XhjOVGQ
k8MX+SYLjPz22o85nZJIhedi4YAgxoL/FSeptuXDG4ZiFMOe7qVRvty+jP03RpjwLQiKbjkKqee9
sUhSWZAAwqCrP/30NTEx7h71byhg+akH8xXwvLIHiDHXWc/pJjCVh3cScEaMUtZYyEVDkscPr7w1
u57yDAeIzCNfLrl3z0Bg3ysTGTBO4bAyWR4oCaWRD2ga2NP4swwQRpJ4912gcY5JDRW7cGGuH5XM
2rQnva4gNpZ45Ep8sVJFBfzuvdtmyNHHI0TdcVZnr4Exyzr3ElHqJBG52g9hSWaAVoW0eNa7cYzM
xi01mMch5XPN8Aim7n0+6BT8YqEob8J5r5CRlZey7U5VfgXktg9NFHRE12VaXGqgoHtsl+HjPk+e
+VQFuorQY8FV9P3KMvM4O+/3rGA0DCPTN348hoc07j51izN+HDKYMXO8Jq2rZLG4AljIV8CzgomP
7BdR2S7IMS4vrDS62tWO6qPyfKAqjnJ8JPb0jjMCwdHCjBAvVMoPml4utD+xFg6heZojlqGOERZP
wdvNLe4FtUxpZ3xII5V8WbQdnc06T2Rcaa1BJRoamOtX1pICydAFsBbnNToM18q3oWO7G4qnM7+3
5UMKT5TbtBrMX1H0yAJ4TkwjJtd2e8BHvUoYirMO+Zh++3pRgvUvU9/IbmruLQFzd/14ytun6Szv
wFpHeuIvFfH6qtYVDlgW85PCgmIK8TBg3sqLder9mIWNTOD9vSMd5Myw8xD+HosS+yJKjjDsmm7n
FqCDIFyTI4UKHWR/r6pK6KQ2pZ58zb+mCET/EDmt3PTcfTAdbx/TYI9D/g3WsuT6VJh7BBsgXegu
A3sCNiK3Df7QLVcTUuwVZOGbXT4xuifQZL7ApOn7+OSzNUqyl0tBo8vL3UlyvbqknUPCvJAdC2ib
fWR19arHkt8kb40t7fwO25t4cgFyWopsHiUlxjI1TDBFr7yTd6pao6y4HNnzbfqbcveKYX0ROVlh
rGyXjwSmA0JYB9VZd55NcKjiB3YIA4Wd8es3pG0fOmj4D+p9mFZ3qrXxqQ94Fb8o9i6/py52d5qh
QWsoIEKA6MfRj++Uy91hkX12Tm9T9BWzyo7u4n+wT3Mn+9J/FDoWurk79kkwch41CNlnEthjMGwM
W6ass1UTasFnpUHTeALYO1KnSc9qTMgIViU7fJ5DJT5mLzNiIkU50D7ecFn6A2VMZe7JTY/D/OcF
pMsNMZO0MuIIuVrx2GMf79U7hNp3/aaGzUfJzMrLz+2wEHfi9OtnZ8L6YeFab7Io2B0DPYNEZO6F
m5OJX+vxsd+nLhwCb2lFjYBbuw21kWE1ePAAr0yR8N1AdsHIFnQqU7hmeONjf1+wJwbQcaVsGcSl
6dmK64et1zaIBlA/R97nlCiOpOkY4A19zo5RBu0yASIJkc704Js/RVVeB32q00O9jz3cSQD9wvlr
h/UPjlnFsGgjf/nysGpjqp4D31CrqyrrcRs1My4Lghb8BszziWpI5mkiNh6j5ogna4PCHTyoC8Gt
8qWos0esBg/whyjQ2074Wpj+niXqhxg3jdkmH8Wl96x7K64W1ls1TTBSATF5Sz3Rrv4rSCF3uvCX
O7Je+lAFbmhE7L+Kh3zTvY9rMwurS4ZSfVIrwbb/xoJAd5RmyoOpUD3dHxoWQjtvGiFUE6xzkH0w
8jexXWKhrddPJa2g4H/WWyRsgSLw8czR/KImfmxzjWOVKjg9gEJGMlR7uAYIcTsyJBnk0/Td0FJn
hGTXcblvPTnD3+Xl3XENJs1tSRHy6eq+Wc6HnLmZMZ2/c+Wp6nhjnFdxeAKBN1NpBMjtXLs29T7W
iEfGRn/GnFgBUp/2BvDUZuON8l87azNnUf1DlC5l3AVQPOS51rW3xT0ecF4wRRTA4tlHeepf89Bi
AiaPA2OvxNiOOrYscvusmjJGXPezQlbIEbcyvvlYCPDvTw+SH08zlrvQ4unE4WLrX0gP/ETi2r+2
ZfPMXFSxijzVw6aI9uM0fU6RFK+CP5gdfr4gnWWVUKWsyPipi9B9gmvbfrmivaCItjP4xT8h5fxv
8U2cpiz2LvIcUnlRwRpWG8B9+8SXQ8ENe05G+IgOGPbTZ0cTOzcPWOXwyqrmW5vfihsKdAxmi2Sd
kF/HzDxjkI/ZAHByHEaAX2LhuaFxEFT4QhOZ57o/J6PXL9+LavmYlpHL40S/VReskus4Hej/IcJd
JM0ZT/zFsoxO9ZknyMslNLpEkoMXa29DVlJIIf0ZlDHYR4vYQDt8mKWSTjf/HWzNCh9FgUZHKgJ0
o1ErgaPSw4arREGAfP5jfgys9VOZHmD8lJ6P9Ho9OX2XSF7d12P0q5QR6WyHXPgG7TwLaoEhQV6t
zxeGd8j6YhU1702bFDLgQiXQ+UKVmiVsR5Mjz9v2oyHl6OR9hJ2PTW1JLqTvgz9f8TPr6Ys5uDkk
N3u6avS94fuOwAqZ+sxBQYM5Tp+NIqEU+SDwRj24SiaVNoQjC4vsmJ1ODtBw2DkobzWjGQTGfux4
weIox0+X0ohmMseMFIX6BOVHj/G1+00IgN+0F7JdI7e8ZZT6SlBinooYpbouregjW3BUCD7Eo8Me
57k3t8aw57GNL/nzcz0rKk044ioIWKP1Z4J1mh0AdPlCtHV0g0xBq1iBfCwoXFTA0I6HJUOYcx+M
QLO/hJu/YyyeSWts2n9RYDcf0xPE0/z0e3Um6s/PuE2Vi4JbmpXMoPdDQMJKrjQcvgHy10M7cuCv
Av6JcmpMAHDMXXQaei1RU44ik1AIMCpCjME9KsqrnApHfJL2t2c5HSlwUD0MK7bm+/Vc8NXbJLKN
DG2lyfSoC+pgy9JFR1Vu9UKXCkfuQrDrKFKvD8VlCwvYcleKL7AKbkZn4B9+FbjXpz/dDVbkCTFK
nVusaInX6XUYfoQvrL3swDQzPWy59fF5MTUM2DlMPuOUU0F2eKFWYNeZtC+hssr9MdK8QJrhPhj4
ynbBU/5BV+NPNCrsquMJ+7GE7H95u5Y9trgFDRAWo/Q3wwr9zb0pcu1MbSCsc3v/uwZ9SnYx2lvy
Oo5KZJ/xctA27HY90G6rsG4PnzsINs1VGqtYURqgjVlTJSksV1vib1sUnlnFESyxumFU+6EujLV1
Wf7vyUB1zbKOXwQDm3M7ZpOPFcjG2M2IViwiRI/0mAUAMGTZz5d+/pooD/cxOHgOWsZc6cuBaH1e
YE7S3FJV5r11Ybxw6XWxWCbT1AYRty8JUp3E2JKVjP8kKw/4ltngp+2GAKzpzNHiwg8y/rtTgMZo
W4Uw/5LfuhBh3dT/7JmTjdVcGCQ+Ibez3OXcKH13ju+uqjbAVt7lZLm3UD93+OXTND+X6bOrZI5c
F/nPUHVNIG4i3fmsOCcuWHbAg2MJqQ9THvqW42M6eRLYkFgmpNRWaht5glc1nMiqHB058Au0vFRT
jpXehJVyAGqkcAxoQx1MF1wJEq3bcEs+2F9TG2mJcSMjKEUZGn1dm4Ry32smFBkqmuzCZUYyDlHQ
BZMZyNJycEaEEaP2HCXar1FaC1RsSS9mC6rs+Z6FOqDq+c0BdLNUI0BvpmINq0OBOhGgQSZTzLe2
/HKDf/gyRsimT4xV4mP6Tn4BJuDqqbvjNVofo4cZGpHhIyX2AJnrh2sT5O0ReP4SmPKwrk5ph8oO
Vqh5Rn0duL6GxpXZkKI0X/bvlMShHvvcwfxnWtu5N66+2P4sSpQZRNMZeGM50DJ6Eh+wJkSiH0bZ
wyGmqhjws+yMZekPE8eBWaLF6u7sFG7rRWQLC2yT4fPmPDLZ3IYd6fH39SuGOkVT+9HuLx/goktv
mJ/Y18Fu2TqDlIZRL1T21fI7+sUkih3LNaf99CvcKjZB1n8md3BjWTUPebcVPvJy+CSiyRe/BCfl
gtJ2G6PT7h4ogWwKlzcGwQw8uP+wAIH3MPav8VtYQOrOA19fOuGHezvpG3u1wXqo2VxRpdTMworR
7mZ0J5k1iixFNwpVzu0K7Tg0YvAhHFjwP7j1BeTB6KtBOIAVUl9o3x+aTLzoxfh7VFlWtUcFV9TC
xE/8XDd3jogls7iiAhDEzG/SYKPxnvW7RTK2FYpTZXhR34WgvGleda4dwFdbE0E/tSbWyN7GQFBZ
ReTzcRa9Ity7gspkOpIviXGf/ycySZ/c3neQGyvkZ+x0Txkk5T/4o3RgxWdu/BK7sPFtmAkvOtMS
v2B485a0YBKxaWUWDozk3GLwj/H5svp46d06NKWgGmUIK5f7xIIebUO67YHWUtXBrGFrRswiASP+
t0BlXLrFA7mMTIA+okyRS5NUamwUzeZnyzQ9Zul31fA1mjOnLG+55a5lWZYKflEpvMCykrtaczQT
sJ1NMKwY2CdU2ePq9GxBAVJq1uhMoZPZSyQRduItDwKNDR09BodrJw8IqjJxw+/okcl4oimJX+v3
DsRJa4DDjtGjNbaC127+oD3UMvlZt3oOF6xp5i6XjIuDBDa/SbxXGEuvqtDGNx+QuBSpR+V3Qcn9
oabftyxMKuFMNtoBMbb/C7d47DUOi4cRcP+qOW1XqZiTRMmi4/MDjoA4aOV8VpnLxdEHcC2Spg4T
i3274q72ragZgUZ9wO8/3mBeoJ4eF9Yo27KNxIN1rlb8zQU5Y0IqnES5kX+oVWDM7591IGY/q/LF
Eweh6zophywWYS+1vewNPn7ljJ0oOKRFb+qOV5Ox4Qd9SPcEzPOfAfPRWD4xfYQq2ddC2lxfQQrB
BTRo7lYMnUI/X0vbDC5HRy3m/otQzRR14Xw4t1FQp+b2sgsvoHQtLpu5GCgKHVgikfBjfNt7gYhg
z3rhuKF0bJK3X92lVKwr5pAQllr/PxXNOQcX+SEahz2ckYeIOPFBJdMAJIaMDuT2ELeMrt085Obf
1TTgwYV1w9e2zmARsfhCcCDNI3L7GcrrvtfYRpJcZiO+CE0NFrwZt0mFPrasudV7jPj7R6W5Vdcg
+ZPWFhpJKpKO/neI5UoW4KOBt7qJjaKGTQUrCLYqwyjvrXUgYNQPgtip3c8tH84d1bD0E2fyk90j
YknDhzULuW6SmMkszDtPUNUkcwsGwTIOD9BMh1ylLd1Ng0ulUep9vbLymF1Z9BEMflJsAoXiQNd0
fOeFsoz+IfuVxnifpuAKB/6y8fUwHwg9tkPiw9T8GHFjke2yM4MXE0/ZwK8ENL8+aEJEC+79iQyY
LFLu5CxFriw8Z57TZ6+NvNpSDpZ6yi93oca9CbreuAb6lDnm5gMVXKu367OdXBEcaBXkoJNs/L3t
52NEpiT5TS4gDsZplbcVyMWA36juAV0FNld+s0rsDA4uq7EM1+ikasKSAsaPqR40JrC8pdONBzhd
38WwGDCzIx+vVrIZPPNP4FR4C7yFLXnxHoNOZQsEOyj2hDnnJMXMe25VZDH642k7qVvHGvhJob5z
ZrCyaJikz6+oiIKrsIDa+EsRn3pz1Ulr+X0YT1hxgcmbfHY1RN/eP0Cuwjuxgg1xSKH9D/XeMLDS
ZzuTlSUao2KBnKpxWsZXQ2wsdFg1SHIfwqUON1JTvg/ROS4kAyL6AOJQH4qR65shbyvT9mDGagXE
d8B6wMOA5xbtEePoCDqzfy11M1J57hOqmL6mq9MNvcsddTp8qKK2GWdP1e/4itqEwb7by2k3cM2E
9W6jkDU9hl7G4WUdeg0WYOechGZP9vzFB9ghPnrdIpKw0UfKZmCa0YVXUEIcXSJ+QO2C35V+a53/
+LDejbrdqSHuHFTvZEux4K4VWaCIZThwM3swpcP2fkZ9/7vqpBFTdJ5LUnY6Yle4shEyRIDLOcd1
AS6ZNhf49c+yP7sG7foSqpJgITyTEw7auMZ8FrBdehPU260pWMF+GsTQecStnLwW9dWi1Awr6fEe
xKEG1pkvIM3DgQB1IMxRQ3Ifg5LTw2lu+gVRyFjAvZ17YTmWbx4nLbxUEUFDjVhQ+qcAfnxMcknu
VI9ti0nTBd76x9FsaFrWbp4ByYQEZwnFzylfp6O5lM4Qxvb1fcPhpA+anCH74/Zm+NhooX0VdU95
NRIeUimEokGwNTfjcHDwCQkSW8Yj2bUrgw4SJE88MYYJtc532q9z0bXHlT9/3DBlBEm51bj/gtUX
0eQ4wMYFjMCsBvnNu8xylxCjnjnfaA7hvcrpof4VoQqa/Gi2t3dKmgVq6tbChi6BcELtX8rGDVUA
NpI1xkBuX1P7tQOJKLuGX9nQREmeo6CbCrGVKo724jzj1bvXq5SKXumxeyA4lJtnXsArfwbJAJPN
3QXITMaunxYLvbkCIEFqsk8vnyKfSkoOePhMXmJrDuIeNuhGB1yzEWMx1JGAcWZIOxBS9rDyd5pf
dPI6tkX4OM9BM2MdYYWSwmNjB7YQItA4/OWSQAyGXzYXLJUqE2sz0oKLYglM2P3PrCO1oXshQjtp
CLceGAWnUgZCIs7/Hf7Txw/S4M8ghkkwgCLXWJdPVeleTx1A65V0vvjxf8PegNd4mVLl1FRz6JKR
HWNMyGkvQ/nC5VhzTBj30bR11QOl+phSUbD1yPPQviW5qYsm5FwYwaoQmrGL4AZfiVjJE6+IF21G
aukWZEByTcq84KIUFL4khuF0N2ar6ayCUzSilr/8ySW0EMgEujUxszpe3eUouXvi6216bgHCBucO
TEP5+ebHZh8R005DmDfz77FX0EAyd212Cd3A9JU+u4PJfmmVGutcfTbeXjLyARkE3SwajHTdEPbd
BZrbLr/QRS/5xOn/hcgNvbvcW+0jhIq7hfxsSA+/Ig9bZud4WIzKHCOLB+XVjuIg34PzXYk2csnC
fcqqHNYd9Xikj68nNBQ+mlcEfVsYLsc6v50T2c76kMr7IlhFiqhEjiYe5o6X5fali9MXFz52EKhR
BVXUK0krNl3KKiTO5kotT6VU8nUVQ1SxB7F3g4t52adM8m1U0GbLPJAYwWLOkKHjmzVdc+2VB0QI
msPaghzx5vEKua2D3Hh2qA7Bh9SstowqdhttVHhl7/UiVByVh6OwZ3YmsNvNIDOmQSHMyOs6Lz/p
KEo7zwIWRJLHY5e28o8BFIvrYK8kZhh9C2xNkjEZQHMHhXC6Gg0lo0dBwSEePt7Ii7gx4632qPhd
+M9LJ+Q6ijhxCHcxIIYeAb/yFojB6vlzYuiURmhDx17SSiRdz3jPbH1tMEgZIkDiv1U2gbReCDba
Botm3D6rXg3hNKax89Lc3LPNWMyRWYphpHYKdC1sxmaztB411wh7m2/0dNVhW8oYb4DOU7fOmixY
YH1efF3960p8u06cqtTTKDOQJRAk2gxynOuqaX22Dv2zzztEKN84n6ouE0nqxnkvgh7hmAe3Ym5q
QTYBLBk/FaKHvKaRDyFoIGU4ixv/IXPCbq90RdVfuwzdbH+mJQJl5nqn4dX5PhXTYLfBJW5Oiqc2
Bb0LWbXTpjiREkJsZP/plKMhoDlAuzgtINCKMr3w4Og6GF2H6AmCgZjRBfgFsScSue6GFSH370KE
o7ndcfp7oNnfqnK4Nj40O1CEHjgz9QL8J+UP0c85LJ+0oNjS030aWk2M5+i19idrzCaNOHU6mRMj
fuiyTs1JHw/okgqwnB4R2ymfwQlI1tmZNKWQ/VdQ35L03qkcI55hAuVN0O46xbNs2/q3L9GR3o6y
/DmVYZgeuwIQ6Dp6CAlyLiKWVhRIIHJG01QhMcuXIb8EIWyzGR1ioKGu1vyFIXE/+ltbuyG4ttrR
jbryBcRiMc/xD7jcCo57hs4UsI0bBwkB/7FgvuTan9rLfN6tDbCu0hqEezBohR7zEXD/z49pzquM
SkMuiqYWJ+LTpfW8oEoJSQCTHRwRjnZfKgfgsEEf7myUWVgXV2fG4ZjrKLmCaMwdydAlkxcWlS1v
dkU2fVPUmqQ/uAyzrJN5jbIM9p3YhWJ8SHr0N0KcPRoxEqwtKKpnsbpkYzizqVpJKcdP/qC6ygqC
jl/4AHNp9wYd+KGbYqJ0TLYXx1cbf2xJoOVivvr1nYWKYE2Y1zvtCI8vZ3UgYSKsRouBG+0lPq5C
2CaikmHdja0N3Pgk3W5QJEXj5OIS2vIpH7+fmC9tUjY/13qatQTFiU5jJ/XAipH+ptFrgQZuucqs
pN7ro+S6Xx5gMK2scmjCWndpo4ntmOXRGg0B064JhhGT9kwAyy4OoV2fwhOaZAAa3qBk/yoCr/br
zdzjzlq/jSG2lZGDMBSqlZ7TBWbGBl3C3UqcntLSjoh7XwnlSw02eJJxJHqC3kwaeqBsG6i7CKzg
Vm871DA9A2Q0EryJZJw93nN1MXDijpxUmD/V2JXQqMUf1BpQHNtmIKTlvA/JPekMxgADighwPRv+
dGbrWwdkHk/E870qQgGmcYn8STbotESTR4szTI5vHdY4uMnbiBxBCpkKzKHwT0+K4F4yoKONOjzg
G65dViU6R2DYp5vtmHtl/KgNQzHu1VKGu5UmpI4iry/JIp69+vLmvHpkqs9vpxkCzF5Nxh/c8A/R
/tyAhLPENRiFYMPalA/s56UchiuWLu/oPrDpzC+yAjFRUk/VbZyhtX2mJUb8zoydIUadBN7AYxI3
89+8NlPrd8kcPow5FOWFWiq27kjKYZpSfMIYmW5yB51con9DnAbphCCl2Hg+iLgS2qakxlQAmfrb
e6BaNN2xQ0MXrzMqfEAGdAi714YVypbDl7tFrZ9HNBpUTrTfidOcN/kmXcRCO6103+wxMpQs9RWO
BLoifr7ci6jdz4hchp5sLk9wknXsAA6YbzsXGP6qyvdlvgprxchvILByblF9nvSaSrxN1IlCnX/l
xye5sQ4FyvsWceWm6Qb2dBs3ajiXmOqaEWvbSTYy8yCUPNZjPOYazqiGdcDKS/yI1t09ewktUyFA
CfYLhInlVNnpcbPxq19Ch1zUWKRHXzKWrmDLwHolbQm2+1a5i0wZizKZA++v7UAkbkZjFp+lmog6
jy+/EI32Df3lTEajGCNSciPOMSkvZWlRBtRETm7v96s6D6HWluiPXJQtY0vOjPf9uJ/zpYnd5LEc
/m46oTNVlxOp3CTSQWG4b2a6HpPiuE7qNeTYnOpS2/CdIzx6uFriaIK/zIXqmZkdIp/lttw4d9oU
7AU3fYKrxFPzK/z0dLMKgI23rVe8KPDfPox5u6r4Z5Irq6p2I1MNb0zhPZCEYOi9luBbACYfFPmn
lEh4lOLdn69gticEa9QqBOcqITk+cp7AwH91r+ecvVqHESQHNICT3f0JhABcSo/2fl3TStSTW5hv
5GDWYtbgo1lgVP8XDrmupwwiaZpbeU5TW3PmVnDEVMBS6sVmFgUNYzsV1LRUXevFFrybGY94tDmz
bSvx8PR+nd6PVekiSAwXdmMpK4qdnub2Q2Uuf9GU44P9zJCyzolY7kY8sFVHEPoXFGl4KxuPQ6GW
rbxCm8m89f3bU2tTRLnZmtIy9ZHlH7AfSGSWfqXH6cRRpIdDZVeCcQSXyXqu/MyNniaA4ZBbPsL2
Q5LNqahp+3o+/CecnthXtEmiKZFwHL5mrQQI9c8+yiQHBpwPr56JkrvJJ7b0jD36sRKj/LMNDG1k
umf6s70nBTPDlyHHa6F/enZt2jiR3EQ6J7bERlGtjILjNs+OKa0oaXPEXnhiZbwPef4nyZhWXpMj
+FxDicd1Ww3l7HXW00jbT3L2Rt9q9LE3GrMkA0PBPwed28fZnmuIRHG+Rxx5PdZ4BtOppkp5jQNe
cvbot9fJ+mUqTfWSrYIKGG7C45hdmiI3dVDm91kd0O3DjbCSd8Katiljeed2cEMT/gQxF2NwYBN3
PLn8nKx9r2BlM6rdNF1OljHm/flcGIOhZEbTmvIfejhL0SYrmy3BhEH9J5IIgoMRFyllOfmnnFFL
5D8vC2KE6dTDIubojkzTh9p1jQgZhB+JZw3E2nJV01bDNOqCAUqcEtPWhW7GoFMZotXnfXnRIys2
vD2wYvYZ9HeylACT2VZnKovm3gb5rCTg3uICZnXcLuw+YPOEYSdAFRboPJ2lixoTS4yowsJLgYMh
xz8XQvwYoHxmsxLe0UJj5U7kyGEqmpyNkhP/Na35EJBvDIzz6H0zEyfGB4P9czYbCzj1cmN8vQ8x
iyapiqFZdus37+qRFRIogvIKLS/0mJ9HSmGgqUQbRkGcToxvJixY+j6SjiVl4ryYKiLhpZKuE/yp
aHv1ajWht3YcQt15tK8GIVecnVB66uflctJs5ffTPkcJTA9H5wOEIsTxEr7G55/PomxUeG+Y104u
z6cuatuu+dKIbRYXgGnlKNS1jZMrRonBonb9cREEPwovXXSAUcWvHbF7fnDom7YqmIlcixpa/15H
9dW2RZcf9fUQOCPaJHog9DTplpWC4icXleUdiIZ5MBv0VGDePnfN2V343ziqC1/Jn1KhrWnaJ503
b+xqD3A31B1CnIXgxtHpEono6imf9FIGnjCD+cIu8OQ4XZ3yunbRQJHqUrHOLcvZlppZ5lFvJKxn
LhVLMP+JvnNxc5cE2OJ5EGEiHgSMMZuvEChs1w+rhzJsEIOmNtUMLB9JbhVxd6KtQ67LYh9ZgpUf
al64Feg+iZZZ/Zj7AwX9rACGU+xqLBvY+BsqGiMGJK7fOmjw6uAtY8yFhUk+YZ7G0K7QX5IPblop
iuj6D5TlN0EJp8G+1uTS+0waGPbsDTag5bZU7jJ/SNrY94Ov8SZlwRIWtbnQzY2d1+t6XKUxZsnr
nyNUxepc8Edrupz2mRatZ9nZjpx3uG4ppV2bSjpaBeCKTEPd/c3IZXwxc+dMAzbuuDdjNJtuSTEe
zvkMWEBwLNwx06ZnXvSfgFThofytOnE3owlCP44AzGAPq/v9ny05JwKrI8wx5Yj/5fzybXLHIoAI
xU+EtRSP1Lt6RXH+hrm1faQtDoK1drfn36luwtRj2lQH8ShzoKtLJ9Xnfu0jppzIQ6aH5K0q57hb
CPDPaqAbK7iswxrbuFO30s0H0MZNvc5LXvxxnvh5lH8Kc/AktM1HHYuWQ45RsF9kl5R0H/T/ddg8
3Wa2YzYa/izbSKlZGmdiZCy/AywSRFPoUbr6EQhaMIhWuRKPvxBv5flAqqHrqln0pzs5oBZOu2Dh
H9CNE1d1sacUrbCPTBY1+HeH6Alrr8TWqu+TVyFo3Y6V6IYFJV3k7It0tmBcy3pUJ4GWzZeziH20
J3lM6CFl3utSUF3pba4P+SESGYkzjN8KzV8z/Ww1nN2cNhlw8DvGbS+2W4LFZXvOQHsVKOExZx3c
Ks4cjhQe0OljKRjFINmGLAF/hAYChqSCZTHsxIraABhxwjxo1BecdCJ0xw6gKPLmsyM+rKIuH7XX
GeF/pJ0y+TY/yqye8WexEpZyzrSLLNVa2ddgvIKgYdymlzgdTC/lb3J1Obke92voE7DI1MNmRizh
Q1L1Y91EkuvS1qNVcwQ1lHVSgcZAvFUUzZ3LKHgXpmv6IPmp4jiacIfzA2fiFjaAuLzfoK+BR811
7A3wrdERZxDY0AjOUbMuLSPxWdzP8Zz6G5CTZpEgkLyFcPtjRMnxxramvfg6iOluaVYIKeqbZepW
Z5cfV+xbdozr1VBHrGilYPsogXEShFC1NeCqkTlH0OK+BxocAdxCccVMjeLxUX26KmVAwCboEtaC
vXBLc30JTdV5CoJ/vNHwSFT8UUSqEF/29k9qdtMjCmKFDXbK90xazYOSHY04DxqSqhtp7gnlInCC
iL6CWTkKZZXu+KRb/SEL8sCFn7q00dW2fKM5dz7QFSk1Hl6wMp9oG/gWFtvwoPo8GEGrH23qZvPl
E2vdouF/RIcwUoYr/2ie+9TQvMo0OEErdCUie9gzbHLpYF72c/g6eENOVL0sz/bf4r8jHxT8bYE7
fUi07F3NunaNlSk5whK4/fWJgSCiEXd10N6fCCKBXmoTJrZ+G4/aoSQDeqME/iFjQ3c3PXnYatnH
pVdln9+kgLxBnqwzbW+qllFAWZu5PiISzC88odLU5MLPVH25Xjw5noXYDhA2FcCtVt6Ap1BUqNVE
/esgpOcbXYKAR8Y0RtM3d7z+WXJOTZgY/t1yOi+S+tqjdpSCy4xfxrJr4WP9vhBeyoplXHo3/8VK
csaEDWWXIPsVvV91s19k2W/X330bVpJCfwpZZsQkQrFs4m/urU1c79k+B2yN4LZ4j8B+yfTndhcC
EEx3leXh/VTgofDs+PViqWXC02KEGPpKL8HKXRoJYsTon9LNez78kUDFyfIn0OflmqJSbywo1hOb
TfCADygl5B8zWU7wXE67lUuelZZoiPUf2T1iQvAa85u8RQvRcNcyhYUHsYNIV6gwKg2pXpqYQO/A
jP4bKXMCmzzMAJ+mB/FN/U9ulhZOXDhRvuu9OhAFvxS3ZdjVklPJqyLlv436dSL7AA6JShPFrVpv
YmKOKtdZrgB4LXjwoqoaa+gmSdBu/ktqdHP3YUL+/6pY7+hcP9JBzAN3hTZMUnAQUQCG58jRjreY
HAwBli+rnwklNicp7GIGz95JF4rJ73duxF6DZxaJutUcdDoVE8Q2I1G7L4tWhZb1q6LxApEnx4N6
DJv1t+rYeRTV45bzgOJzCAREq6daP97p/feJy89cGKZ1TFny64bG5o90P9pWxtdGbw/iWIRWySJK
RopS8Xrz8Y8d9slV2YhTkiyafhlo/wDqHz4rloNQZFGfj55vp4Nfi3eyPO+gMqPN0yLvEFniurCt
lQtRgZalr2l4X++RUBrU+7AelnJrHjbaFjJ13n55y4QjNk8WoNL/GwoofyoqR6gEAHUmKaaYbWS/
enwVwcIrrJKlvZNNfTr2agSLdOdAOUS8XPoPE5vcef9SNX3TzkOtK7ialq5VE/Qc0Rd8qT2Qz+Cp
fQ1Pq9y1nrd4bClDjxiXMUyiXMRs1Wv3bc7RivjmVavqJgOJer8Hh94TaTLtF3zhRgFWo5FgO7Fa
tpbIgWk4Eee1Nc7zxJs07+5H8CKOYTD1Gae8dqsMa9E6ICR33Fa293+QiBPK1lMarFmKu2tdakIz
S4ZvNyImIjamHrrKf2UimwwuMvGXaKhLSJPJvCvVRYlJUsFGcUapggefckeoiCdB+GwPnRkm9jk8
f/bR5lGud9we6HU+tUwUeORxcH7X05wI4Wt+LC3G7z43awZT87zkV3bHijJotfZsmXWxWqsfv3t8
xwXY9Y71S1icyUsoor8UUQEPvYgGpMN1HruBOQv5fUG7vtCrhdrbjxHwMy80Z7CIqKXV+DQFCIxT
k7MLWpDbm2TowpuQFQSChhfXPrZ6cho4jJxRnhXQBB6FQTx85GgJO146OlVCHm7dU9mTBkLWqAiD
VP+Zfge+fHrS4tsJdXUi9ebiGHAjxt6UCIdez4yk7O7bUSjP2Zhy3q5pcAEtbtUbBT+sI8pYEWHB
2tkvyCKq++JU0WUtXsTe4oQ9Ubc9+kPXatfazJIg7TI8kjPYix+mY0AS7NJEQd5Qzi++JsHAZCBo
//PsGemMTO+D97acrl+IxODYRdi9ZPPXWaUidpJcyEUjbXvdoTUXpk1GLJh4xQppCQN3ayzdgKzy
IqfyJVnKkzBtwLGknmypVC3vHgRkDKdpsYqq5C/ViTU/xdWFUCvBiOHZexdIp1i/QMT8CF7xyTjQ
h03pneCd3rZEvrdzd5caWiR0S5oY53IVjH3ersgQtsdvev9VHnHSQWIon5oh32QKIGYKqAjvSGuh
98PYSF0FVlrKvY0B6F00UssJncBoVHGfkoNvzw3usS9CnP0P2YVw5iMQuLZE70PcimHlNQJhoAhO
+yQdD8zikB9XFRcm1wTiuCdcVbCCEnItkBlkMleT8wR+Q0pBCfMqw0RhDrMs35TGXl46bGFwWc48
5J/W7xhaPwIyqz+rZdBiIx6OT+duYiDKQMhrvWuQRnJvRZY9lxs86U29YIfxxOgQ1RCVcNilTXoC
3I6agabH9iBktYXeTJ0q/X2GdH0J2ss+WnXBQG2WK72R4HjzofGy61IEPBSEm2Q98YUBntGZorpp
ywF4OPPKaHdcwR5VcLyvWSxL1sJsT7wSGiKZZygebkZt5nnWgD4udr6wlcGTT5PKDLXL7JdsA/xW
7XXkdMwaqVxjXnwp63fbJ2wFPfUOjUlseOFZCtQ1O2UtrEVhq47wVmzAYQRAU4+46aZFSS0m9PJE
1v8RzbFsFrWlwFLYurG5Fnr3G9MDZP01kWykg/Ky0H46Zp0P8GCtOKL0c7B9ejNtve3ubzE2Mj90
9Y049JAITDliCAVrrZncL2sRqpcER6mQMdY9n0Hi128rISraFwsQbqDNWg8ZlD+nGPf9tTjLBnM0
jeA/G6CM5OoMWrQFrP6CeyFYFT2xmipz1R1ymIU8EL5rwTd4w72qfa/qfWmnV9Be+forLflBxcKZ
ORytGpnoEUQqCn+35B3oK/eq599na37ri/JQaXTr2M+27K6nqFpON1R/h4uZ55j6Qf2OVRkE9EIQ
3hKrJPvjMzkoOWb0dx6la7RsJ5PNPR2ivd2R3CVKBZ0Tt+AeGf5O8d5LfQR0fTCDpCF+szTm0hmG
wPqcJk11p0KQkeyH8p0muk8xJ4VVp69miY4jQLH7adldUGCB9iK0FkWNqU5EqESPd/knpiBwTP6X
jCF8y5xpRVaKwTKZobybHvIZ6RUvYfU6dqEKi2r4DcsGIY5yCHX12VbP456cNCe7RWzjkJcZI78v
8VrF/QMv2D09XtTjDObnXZy2iyfbxeVwVJfJgChZg5UhJROPaHoRQvezjF+kVJd7m2WTSWWhYirb
H2eUUMLvSz13xjC2q6rMCKzpBUPXAoPuvwWrPtk2fp26KYSKq2yCM9UFCDXtdw9twKQ55h7jaMgV
0n0XTAgqEutq362ahVVjkl92OSzetCTjpC+W7PW6hiKHCW6Q2/TtoYhERcPNJsxvZ7TSViK/At/B
EBWyyOgHdnwvkW7ynzSo9RhNQQpZi8j1qzWg4G8JUojgRj/kxvFO700IlqWFwC9/XRuXr8UkTv1q
qy5uarnWTyh8cgcy7QEe1S0xg1O/EYZXSBg2N6dYx2gzDUPKj4fUUC2UML0jI8YOxovdDt6osxnY
3bY4Cr454GdIdCYtAvyQxJtKonUeZm0T6rngdXQg6K0RRZEdNqB4To+86YEMYW3VDGWO2pmXO3ZE
DsK2fhEeWcbSD9+zCsYwoKf3JdoppoFXNATsFGwPGMMHQw4dzXzM416vkpTRWMicgk7QjZXAejWs
sCKwhp+z7G1SgcU2MK/rzmspw3XmMQuQERrNRaspoOYwMnC7UvOsU9EIv6i8U/pu4h72wxJZLudK
0tetgyW9tE1dPon+K98oXt58ZWr4JMoIXwzXsuPqwW/hiAP9V5kj0j7T9APBrwC3z9AqkUobG6sN
pT//w3iVe0/k6xaYqrFvj3Uq2AQvY31eF41dJFwgwSKGAILhUmluVqiOUlhFuxQriJcxuwNJNWZS
BSBD94mCyQwfdg/RDT2tzQnLJBT44Hhmyp0pma7GuMjpKZfnS4s2jB94uLgkmrgnvMZEoCE1TFca
cdxu3Cgg3DuHKlGhSc9tRps6E0IJqLmJ1nqHiDy4zJ1aB2vdUKu/6rVZ2+sxTmqVr6QGZjtrtM7d
Ht+jqZWs5L+rrfjnWgEaTpxQFB889qsyP16Y9rkSRIctwMr+iuGzcFoqjg3bvCoqXc6Dz+Sq0rgu
uDdPtYVBb90MTzAA5stQW5wW4up6KLgx7B6u3EAA/6SEmxwACrJCT2neoGrNNR1hB6b09MgoBd//
8uao02wq/UvkOTpdWKllvmgfDMJPZqdP6ceyGvKqDV4PGP/u2DbtW6tTayp4kqgK/fVq2QV2FOVN
flDmUApxw62ymLLb9ckMPXccSyAouxD7b9ZeocmPFcDR955IN/lhup3WMIX7ZcUXb/EXzJdqFMer
4dMXoZVUk5gBxhPEUbDke8EJ0hMcx1rz2UdtvlbFCeXFYXPMirzg4uB9CscF2CHsoE55WS1V2ZwB
uPf+iNjjgkI7le5W/toSVtPcd39eTrOJHsAlWDcBy8hwIvU9haXq4CH3D4QmFrOQkxZ0BF/A/T+O
fCvr573N8ePfZYrCsJrTI4Cg8QyW8fpq235zVuKH9EQvS1uZ1gzkbPqLI/WZSL0kJWSHCM56f9c6
hB+e8rXRKoX72klF9VftfHw9pXGlWb64Gv/x+seAxkC/ycFGztyDZMA92W3RN9UyrCKDbj6djDIY
Kfh06HkncJDbzcoH2RHBjX49e6uYqc1PU91Prvybn5PKj64H+CeR9o//BzTjFBYPekHI9xgMxSNq
o6qlZusxITINWshT3FBE828A7aMzjEAwZA2mIPlQmzPhzSb4/Ekj6z7y8YQC1OEVXG+U3MpXKJ+R
uhj90t3oBIAbW0Squz/3lgrqfmQVSCCVJuIwmSVMg6cpj/8Vqh17pNJ1hUwqYtI7RAgWfau+q894
W86prmnpDj7o7eZWeQAOuVmrqf2QBikYfyV/V8B+o5VYUbrjj3zme78i9m6jXa+hMkDqetkqhRA3
+5bEL42cSZ+lFiYT4AqWCJqEKIhoNtYBVDvfGNWN+RaszON3/u7Ps33SREmE3of+uqSZbM1oxMMa
wY2au5WPnOx/PbGFHDbI2f0Boa683y0+C/33Uz6aOmgxbWGA/J+SprU1gewfi2n2qPyamCSukp+K
y16V+aPx+wtl9AKSbsJRBN7Q3auUF5TDqctEuKf8yxMeRQ+2PpbQFZDzNJNf6efb5a2q3jus+h9q
ljlDeGPyhtGQSYztURWFQU8A/fBeMDZ3y7FVmhJYc20/qGgywJcFrkNWGTXGUpic3aFy6+JFXtTh
MYsuBqeZ2FUqKV+4tPSutogGzHiMWZVDLb5L+lWmoOO9e24BBEx4gh3SGKYrZF6+715sqAykJSjb
EpC3Vf7ZPF7a97FvVBBgwItQDZBqxtEMTKTpi1+akTkji9YPcoNLPPq6rxwhvZBZZ2DIgO7V/lbN
KRFTp92EapAHeUaRl/5UoPzJY/aZF4Oc3pWltEZeUMM/VMAQG/0o0DH6STEYmxasi3WJ+HTM1cpK
269yHAbrqHUXzVci0OCkmHEabpB+VTD9I9vkiVZBtPqqvZDeTVJFvZiWBhKhOUXfx4pWLyuO0X0k
hxVwowbbntFCV0NIHkIfRw4JP3knEdlZc/Clfc1KlAmIVD+Dz0JtrUqOZmx+tmoKFabjRtgmro6i
jrbWuW9v6xwNIbs5BjIq2GdU3KvxDWY7XTJqczKCLGse2qRWC6y4CSnybh/8I9NWv008RNkC3YmH
x9aMJgNMLDiQCB3pzpgqxlZODE6Myj6frhHuKsRhikxh8KvHfEHrrM9t49+dGld9gtbjQRWYwyCZ
0Y5ZT5kpw/6Pnsd5pJnDiopPcRyL0ErXkiNOYU2cKCPsvyXl2K4esbsWJDjM+hylgFI+4CTePEAb
u6pTcxbO2aJb1CPju7pm/RuOR+xOSiQ3gOnBXno1jM1OPabGurun+MBk2RZf0f0BKdOMvia/ZcVK
RZw4LAdn89o+YoUs7grB3hc27/wM+N+LPWUqlfo9UxV2IXMjMd9ZvE0kOBkR2E5IxHrHLtvfNxiJ
bsrdJRLg2TTBTqX4HQCpHfiAzx4JO+02B4wM2u9kIy1pYTlSjP+3PfkIOQQOtRoxDV4S6WphwAed
pN799VYJxv8ZpyLXQW3lBUcC3Tv38xA0tpO+BCtzcWb1rQG+MI1JD0nq3hB4e0TFKqvmrw1yo9Ao
t885C0TR6ht2R10KMjTaErQg1wKqcazIc8/rsgKr7ygJN3LRWuiSeOJQH/v2aeDZ2DFMQ07o1fJw
0u/nLR+uvWuqpgiIddwhH6R6tx4usLzkanxjFrYMRNKSZFlx9pgY4uctGPQ8CFjH0IizbZb81KYN
2oDjCm3EJ8oYVVYpv2A+Nvc43dmBhnfhSoNzS+xGLHFTHVQZ6+VUq2n8nDIT9JwqXPZpDpcd55qb
0+ngipqehsALngGO/XtaBVx3RPlPnJeV9+6b3xQk8GrZbUSeSFokV0mUng4dwyjXmIfXxLNOzbdc
GGuEfroDBOUSAcSJ3RQg4rky1XK+KZQ5qSwLRmOPgK49EwmGEA+mpHoRS4a/3lI00bQmmkvHYarL
f4bh9kbD2hTrpbfo62WcZe0G4Pa3unPHH7SWP284x91+xvUPO1keZ0o21RfDpGg6JxT6Rw6U3vo0
VDMsyjEciHBDeBtxaRaJ2/hrJa5wNdihKBbv7vLFVltYqMsp9+ANXXTNmpKYRIFz7XuI8546NFpo
yhovStpeXosbfnk8nTMe6nwGL+DWMXBL96drE6Wm1OonmzWbjD0YCyLUz9QOJciFTwbGG6kqLPrj
fd5kOkIEGQPzlbW9U97tNjp5PXvnbpRkIt9gNolBUvDYK/ZcdfwQ7YFac9ELxPcMg3WkFaA0KerX
b54MaTVKu70aVI1XC4S/Q8a11Be0Eu/PMWIU3Fa65UHt6qIDr1fwpHuKUoEy9LkncQjmVlZU/8/L
V6J8WGcjd+mjHdIZEHZxhPn/lUfVYjJv9OiJAt+wL0aN8DGQ5y4fpkve9hmH0Qq/Mv9SdYI0o26V
th57ZjEL2CwYaxsxhCk8jLMWyPi4NazPBVhm1I0Hz5HD5dkbpeIZbg/sloURN0koZC7gbX5N+ZQK
oU/pqnwV9OBQ5qBWFVm1zyTIIqj2INaoQ/uSahRgrJndv/R1n7p55CMEFXozSrnPLP7ej808tMo1
YHZWbvzVjsdNSE9G7Xp8juCtsdjTx/Y5C3ag79xR30VuKnPIX1wGlPo5gNHSxkOSLMPFN7TBCdHp
c3lvdgepu4AkE4OQv7ZnHZF5O4hZVHcFdyPtAofziez+t/Q5YfWSeBk3vm1gM9Mwkh8hUvvOSp47
+toXU9be0HzWRPWOFjoaG9/MWFTSl1AWQkt2ukw03Adlapy/IRo4v9Oz4xsp7ozIP9cIyt/M9ZGM
Cx5tajS24aanHQ3ZAvKeJOXwH9E/59l/5aipqxxKYXyzxd0CuQQLsXWozlDcLFhbMCsGelh6nzK/
Ws4GfWpznoBBlKjdGUE9wuD7SNHoD7vfSrJ4UH5GpjYseJ+matTHAEJKWXeDukKnynMEVC4VlFus
FXDqPIvrzDlJHsmONnutaDhU8/Kj9++wHY789v7AfcvUyUFyR3Xg1IZksJYJEBtnDlkYtuqHn8hq
FmfjeAepQUHtdf98S+KRp6+naUscherdYgotVGwbpm3lZowIycWin8jaVu8UuQFF8Bb4w7AZKUW8
MgSsG4wf+eY7Gs0mMLz63ARe6RUIS54Jp2Ul9o7R5MiKN2CT2HxaaHOzmBLLpHaFwADUTDoLxMRN
9pNe7pE4kLE3BuakQJK6mzRg7JAGN34YZqak0DMPSgd4hSUT53nZ181M25zt5CC3HTPXuXVEoZLa
91SOyJ09oKHoy0EIlfs+Q5GLmQrpe2INV0Dw0fmQWpRqS2P2Nftc6wjLBH7YWIcQJzy2StmFQvTf
i9e8IIdufEJtV7PCckko7V7Gx7mFihq0AA9lrQEybe+UjVU5K+x29wHRct4kjt2WA04cpxvy2q2T
mq3kwT8aFift4eTQx6BiQtccznZjxomAjXI9Kq6H6oCFMR/4DnH34SadqDvmMasceC8sq9FhKF88
0EpthPWi/569AvtFohdDgRP93KVZP0HlrtVMLzrGN1XJN4mrrlcq5G+ylU2WaUaGhCimG1OLM1Se
EcsyO6F6O3NyRfukwJat0KmetpV3TjxgxyRtln4ijCQpKB2Xou10Lpzuaa1fBjG6pJc9gnUpt6kf
IqzLhwjshngYiCo6Hlg1Tn8hn830H6ef/WEi1Kb0o7UiBscj8iA7+/euLXsusG6spbARNhR+5env
2bZmbtaNNfhuVGBdRwjxdUZ4+zEO5dtWZYIvgOTzWktD1sv+R7Erj/s83zaAq9rQ22feKQ4/CJFN
h6JPSWaajCQ4QqBau1Bqftpqrc/tCBl+UG6g1r8g9tO8YqJ2K8BBGb7xx3VK6q+VAg7Vsl2/EJ8G
5/CDQRatB6AhbmpShMoUlmpYz8A847HXxK89hJpk+xlWcKmeiz1Q84NiGW8bILWzGWMk9b0ncKEu
LsyP9lu2P8sNgHptd4X3RtiemhOKTeLxhh6xoVPZRdqcd16JrGu8NSVE50X5yb8yCRyRD+84O+97
CXuviiXG9BebFrD0Hff746ttBNXaBaqftVF3e7fga5m8YpXzSDZ2jcemNFjsmydPBEA2X1Ag+GF4
S0Upt3EvSd88AARzzyFtqL6pRURHBlVkixRtTvyzS5/D+i8VqD1fTb6bTkSIkWMw90lFJ9kGf7i0
kLEvzRnUyYwqH/jf4UpzwUe1KG/nmBBsM+pR68NIn9Mcyx2eI5nGfPGBUzovewQBvOq3NoaDmcVx
/FQ/248S4jutwcLeUdvUw19zvypnvNC8tjzxVde370n6SprYhsLgOU0GloYn4yKMHb/I3JX2aDHQ
Sv0w3WzDER+wt2QFS80Hdtql+5sbIo4SWbnRyPIsGT1d1+MigTJ7Atl0yIefBzzinG1KD9UhUnnv
U1ARamjfXY/kCzitM0lYPkUOO3IWfVClqgC3IBB+ZjAZxfMkPS1+IpvDBzSKocj/B8dYjDAFKDF1
Oge9aaFA/K5NhA4zUJtMYgAsbUz2LD1h1S8DAo15Skj65ughGXvn7Blf2FXd+1slc+YcbWUpZVi1
cSQOA06xlRTiAYTchd795w8FGD6Z+JylKL9+EwCYxQMiKHPTeVRgwVQzJB6e6ie6ObB/5MKY8+I3
DcyK1rk/cG4Nidk85mXIQeG5Gvv25/o6Io8h2KHsfKxtrS1zG4dFJokoU74TUC1xSpDk9SYfi8/u
IfwrBxfIbVB8pO+AjZCICguj1LtU92njPmgvNQZE6VIVEsEBQ0/sDpn3GF8ZriUUquUSiqPp7VR3
sfHVkLQZlQW4mB5XiqdtEQazSTxjdhQAjOLAqXGN+qlAg5DmBYCgFz/+GfG5IUDEVjB2+p5l57vl
Z2nNfIrz7RPsNBcXDIOID6FttVSPNqdnwZh5LjV65SWTOIB8pGLpVBsOpIcuD5WIk6PcFzmjttJY
WUtD4J++K1pl03H6aK3Tdpgo3sWFqow3/NTglFLKwGFAzQxkWPO+3wc2avwWEWJ+BZ+79JLOjgTG
ySRUv6oY8WsHJyLyxTJiSD3Kp1Yd2EWgrDLtsftqjKnTD6P/VfxQvqL8cClp0KZVOUGVRqlnqGAM
edfuZ30f08HiYNTQCsMGBJ/MmLXkpQwnUs93iuI5abmU3MRMSmSu+Dwi7e3P3Ln59MbHb9mRA9c4
yWGmoX1D7j5FPx1mQXj6tu41cKauUAHJT7cXqby7TDsBQPzQLCQzw0sE4hDQ63S+LywBx4aO0cuL
tqKjTL4kL+nkmL55v2KNsy2j9ve609ep//8djp/4e/HGhy/6ODHxpBCx5+UTsFd3EbdI67rJp5qy
q/0nqFjoTB8G+7YnTBOA9spnMPyP8T8i2egO/HQUHJd34hO4cW44TFWwKgWmtJoWEnR7Rt0nDHxu
6D0J0rMx56TkWQyMxaTmpbVoJ49KAWoUQB+QIHFwYHLvD8Y1Lw2PQ/T+RcbQjKRvxb7J/0STAfz7
iJJvp3KfCu1SrOGpSNi4Mx4ggJ6Ug7YDqjAFO7SLwZYCRK7jSBaYg+fO8y2sGpDzSVUHgz13mgQh
/TSJb4CnTlICcsmY6aVba50pO2Xj70JyDbYU++yMsLlyl9GrwE/kuCyoY0QXd9t1+eP2/TmxNweF
NCZ3QvbJnpi7MkTJb3mscOR+mkSUvi+zfPKrKeaMepsrhu1tBDlO4U1rXf9d5jxBnDyvaxNQzzTo
9zzPdFXnS1d0Lrl+pFZc6WFqI8n1ITb+UOq5ij1s3a3UR5OgJJ++daWdOxRz1ZyvKlKSq6wNu1rO
Dc5WKiajqLP5nW7R3VpS5MIIpjy27UgOYLLm7IAlPmA6L4D/9fHYJvxERrCnsiZBPkTx8m+TXEhq
qxIwTbQSLb+kHD+Luo1io4iyB7FUrAKIW1wExlyIO3MdSPYyIGh9iEzpK+zSe9Q5Fvw8znSZJ8tL
uyqLrJA4PTnXd9ChAgzX40uaGQnUCNaDbWiiq4Oa5Dtbr4EhOtsKS3knqYQM99WF6K8LxaX7K1wq
M5NIvDlaaL84DqNJGsDmZsziKM490paRRCYwSMFnnavAHS63mcjTuk3t8VX/xWi3HqcnO4dlpF18
juAm1tc2ymMdPcwADO1aEDUfZrKN4AT4ZhZCrPehR+euryFOJn+mGZDpQnqjlC8QSIZhx5bSw3gV
yyc6fwYDJ2uJaEY0EruZkkQL6gAoX0ITEW3TPLvVAl3t58pKUEu8UxuiyE2j10GBj8+8bKsKI5jJ
OK/8z8AgbCuE+Y1U3f/UJAD3d9iQDEFRuFJqUCu+B9d0RmXhup3sZdqlGExzo4ERP5G7YQFfro64
yX0EPS0k5su3ZqzTvGoRW1akmxO0hdV/f9XBuX9cN/dvVEMb/irlpG38W4B1r5cQ73iDNOdvrhnp
HnL69OnP108AUqgjwwuB47SgwuvO+9j9r7NVyJan/mgSHnd2eMqmcFGJzmK97ntsGpkp5G96hJWu
WjV5vg9f9CeudHIR0RJalc0eYbeuZREYissCbBsllTAOJxqbYy+qCBakeapHaqQl4p3VtwYTk2m5
QQ6Y4WPfHy5gnZh89FCfLEyfp0W9K91LsHwF/YK/W5udx+t1L+nzx5il0D1u+A+kSgDPxS9DoUzq
ehbse+3l1rMLLSlUjfPi8JqXDjibCnYxQSkSqVODDXO10qvz0I8HFo2HnXp97k0msh1qOpxQrQEx
bfaCI+vC2jfG96GfQ4spPeBAoILV1YMTEcJvti29u6lYIFU6MgBkHyzcgsFMI1lPkzvVVSewRljR
69d94+WWBPT8AE5kxX4HI8ELxa6bO7WVeC/zHv7qU39ubRyFQMS3UphmlXsEv8zbQLXibBJg+m3j
NulP8vpWEQcxyZy7kNl+R3eybtpI9WIkOKs4AWNt09CcB4cDIcK/jIrP/egRQSwabZPqgKEt/7H+
2Axu+8IIv9hLUS1NyFA34gA0nD95iVNN9IAe/M2Uvph8HhEYbk4w5ozkz8Qar0Apen/in+MfgRW9
NuxzR0RvNeWVfpQ7jSN4Ono18Id2QZaAOP3ry7LdIzu6WZNOVw4l2KqgCFtCaLcHadQmYPD2oPD0
mtvIZh1eOOTLbdvzQbfLUNhM7DVztSSEkZRlqQDRDfhWc6y8IOtrzuI0vY//nWTFGP1w35BsPtGi
Mj8CWGYSgbMXhqYlD+YcPZgbb/BLUhZhCmti4LOgc9XI9LG+x38CSrV/u3UfB+6ukOIX3aEgYNpB
BkZSsVeyfUuMGcO6kgaAPRWddNv2cUhx4wfHm0dMsPyiOD9m2FSgxzHeOM1bejSbtVdHgHxzxfrW
j3aDYLxxNaDCTg7Nj56BcruPKdyfUKUIalMHieVOx3KN/C3iuQxBQgmqFLswOBQ3HALrQb4tH0tf
W5/iI6yj/NuqyKv23Ed//V5cxFMGuRJonkd4m8qXTmuvJmvv7fvOgy8ZVZvlAfQeoHisaWjjsSnh
OH8LaL2OZtG4QVL2y5ypaadiWaFBwWHE3d9otvk7R9+6cW3PFy0q4mZh4whkDnzhOaY75fI1Mi1z
lvLC7JD4SKBkSjEZrQqt6qzi/JrZNAMbT/GAUzT6r6ZnJLjbFhgth1tpGzewYmZ2A/03+BiUaVAA
IsiIA7O32feF88GhOeGXMomPDFh9K5IDfT9Fvk5SSvUvXkvTmwpnqCI19tsim03iPQBEdRrb5r7D
M5B8Q2SIC+oWBHOqBybVXNXae0YWj1C+Xg+aii8n/2EN/OSimRai91XU6skfCov+bMQDAZePJcLL
FlfBfUO76Jnvq2l3UCQNrNbKUb/kWAZaRGavF7f7ilHdi00TmEaj6c+u107KceyHUHQhsyJG5/Dx
Cjkv6rC6itzW8xAY+VtLCkqipb0z7d4H4Yhi5NA7CW37fk7sWJP+mvl/hxUg57DVSv8reo9Jf09v
v7b/n+UuF+Fuu143jVVsNeQzdgXS8TalW9E1dSPO4h1m+X2PZscxmGYo3jjlXSGcnOMqsvTYrgV9
YTR/gE8DdhkK374QZBzKF9jM64tZiUA9x3JtbGHgvbDhSyikEBhCNqgZttUBbNWM9mNyNz/Uy6+M
mGGBoBvAXYSiHfsFopDsj341sPFhA08dBA62L2xzrOR3BZMm2978qd5dYj4YONp/d6KOYqYgIm43
M27z592Jc2/YJEkm3WJaGu5EorbOZdPcZPJ7o7HMo1BEjGQ3DdtEaIXcRj19n/GikRAcrZHOugNF
DHOOj9AnJ8Sr4M0I3Lxo7kCvgfCuvOUCFs/ul5q6uapXZZIo4MrVMxpJwtKBC6gS7EcLT1gMjxqe
elqXSfEX1eZflgqFpdQztqTVrZ2at4RSnadtzGpC1C8c8zWWvGohZYcaSw+ITm/zdgbU3eGzrRQa
A1qgzEfs+gV2EFE2Z98cyI/NwUM0KWDQZOkr0WxG2MEzlfZorVVjgfOTy1JsPlsmKBjwel7JI4fL
6moWBPYVnwrGYVAxQrM8fvUjAUnL+T8GLcFmGppRgx0svDg7XxCiO7o6FYI+qAUV4uM6c7x+bUsW
FyrfLYPRhduQvBQVzCL8VKbS5t9PpU3xjDl4rF3MRO2T+Aw1pLMZLHFQmUSF/o0LzVgocEchwqcC
A0A/c8hAXJMO+RqajCO7Wl8khRkZmoDBowJFgkQBh13rVPWr1KDpaeidbQjqZ8dvcQ4D00vcr5sP
jdM0B39kbRUAuG+R4UM2i0jeJasHRZ2Qx5XK5wbejoFlq3x4hf4pVcFHpzVgooz8kIUjmKVeNIVi
GnpyKIVcsXrqlgJnD10DpdKF3fFyk6bgFDUn761ZE9cirBFUw5Hk25ydyxKY+CtB8HmIa9jzVUwY
JXR0/JvJ5SLHPQ63Yx6VXd9PcXG9zSD5s7QBKVy6El1bf72TR5/e6Y/NHvkwsctKY/xAGM5cM6os
72AnzGb24KYvu4teFJ7CoVAXN9nOIYw2ufWjI7DL983LwFp1tYJByySIEygievQFczDdrgv3XmhK
vvh3838KeLqPFuZ7mE3oi17wqZ+5S1pFZBG5iIJ9MSpqW42eTZLFgJFowpknppEFewVvgdE/KFJm
QYiLne40CwHvBCk826vb31o1Y4H8YI+9qCdvHTN/B4eUN6/c7QTXbW5ZDTKNSQs5161FtFDJ5n6M
poRres+JIlPA081s0sklNYhiwRKzXwpEwwBAzW/U38t8OE3ZDl15wJ2wu3WdCEjrU4tHSwwUr62m
GKEpzZh8ALpoQxL+EFlACndNT11l+au1a7u9bvkg9MDkFFe0FRdBOnGaWDdC/f4GtSxn0bMU4lQW
6ksGQocFslJDhw2VFm/WgqLqOv6dnFg5+7AJXaNwrfPexW8S7q13Bmysvs8c+ZGhzIlvNSc/q+lF
/Ok7pmPgtDE7I3RsMqSYPD94gb03XIiHz9er3duSCH5+JaVGiwnM044vMie4221qVKNfQLE+1uc9
i0WCTZjkmZ1m7EUoHs+P5PuixOLxO607Pikd6DnvywQ5TpkB1c9jnkSBu2jxpn0f8yigMAP2wxp4
UDQ3C0Spc+MbzB3XP4DpOiJCso11DaV7npIYYiqq37Uqa+Y/kq/wcC7Lrrw0IjxUZCnz52H6hhb5
t9qPDCab75GXBUHZuG4sKYZkyZWTFVSyfPesrQRlN0/C950clJO3OiENoFDgVfiT5a4T8F6WiSlq
CXRwYo8m7FUp8VutJEnAnGRtO/4XLQ4KY5ez46MSE3tRUfnju56aHhqThENzyYJ8sEr/GOMANDTb
IcEPIqmzZ0YhTSWf/09UtaumHXHKmWaVgCI8WgO7glxSoRZ7VUJvsnnvT/tKV9cHNoqZUX7NfFf/
ZeVUZmzgsFV2jush2pUfja7vF39n+IhpBEYkVpou99b7DdyyRM3HM6i7NK3mqO+AIFIvi67RJimT
XARpzNLneo+ozGRIdDiisxr5l5WB2lWl9fG9/bhtmbSVYSjof+icK54trSEgGFG4gB6wwdCHQXXI
cNk+5VYlNDqWqmp6qA3EUkvz/sE85ArUNGx7UVSF55hwOtNdk0zki5AEt7plhQ4JEtU/oZvcSwBM
/6sG8tzk3eVT6mdg56s1pZmZ7sswbRsUdw9uDtQ4M0lJrFmXQNY1lEljDqOnLREk6+4P0ciZKDuS
/VeTU9ODKZWrW3WwLKhj0zXkauuBQ3q7GQ+QOB9S930FtmJuGRcJKo+sb/OGmbelQQ79S9aBKGTU
pAD31SaPXq4Q3slkcM0OpJeY/5fVVKCN3sEPfPuunXNnmReqmhfnNz4+QhUdcI8fMfrznLoypUJN
RhvxSGADYYO+E8RF3pX3rx9+e7A4DGK6DWUG6qSqeqc7HmvWPKArail9iMyaYIiFe+xO+DWjVQoF
EYKKbxojYMwwUfFY8M+BpUuJy+u7jmTMV7t+8+41jkOq/BPubeZLddAZJRM7/Aul/0n22W49OQRf
3jeHI/Jmksf5nu4JsIF3C8a1mI8b8BcFjnVcpFdNrYrOVZhFr9dbLkxObAaSHwSNjNlj+H9uxdFP
5rAuv+HdA3iK8xcPvG2J5M+236KHhXWGAPDRp0yCcDys2Hepk79HqGKFR9eIzrhGQuIH3xq9towT
ZeNndXgO0qADrP7l9c7pLS/oC5zjjos5D4jCQgfNu4RZmd5V18OZM0+MZQNg2NZXI9htTJEEM/pd
sXG0COsOt5v/TLIQ424d59g4UQHgjY74roX1uffBnakr2mBogMc7SqdOhqxr9qlIvr1u0rg9Zbje
+ePneiUPOxjmSFDtMLvLiMZmLxfNUVFQ839JGR9NK+EKVThkNCB9lXrsc5svBqcriCFk6ObWOdHi
4TBWVvBYI3CeWBhFqtWsgegJYA09HN8R6jRFrM4cssQ/SZCTYUMO8s/iZQjFhsEAKtEilAY5rswW
BDcLpf4W8kokvtMC4+6Cqb87Pyv8ZoI0m9Yx4cP7XOrdiYSRSQQem7xyDd6LzD5kp0H+gsBMXICP
MUm2cvSWgoRiewM8TpiBtOCwiPHveQczv8dKKepVtoDr/ZZm6aDt5WzzE9pLbeneX+SI5nxOgehz
SDJtqclVce/LXlBt3crUV+AwMRXkyD3mvio8Oopp+wtGq3HEcLfzxIMiVN5F6a9fCFEWQFBWHDg9
Gy6Fa4uVs293DVRHzue3xfvrLHecpStz5rpC61u9NmvQpRwVV3iTXWELliNn/S19FUv1AbBCNfXA
Yah+LZZxo7uVnSTeADqrFQKu+MrHwFN+tJ4HfdG1KwrNZQ6A5MYg4ruaEQ83l7MhAeQjMUpnddlw
yJTszO/CM5GFuLTS7NGe+uGYh3bKNFwWVZ26GZiUxM7SjMwp3PlgKr181DmaT67h6ECdWVx2/Tkk
IExCAbpe6Yq19Go01QTAxms6kGNlqx86n32NyihZoBQh5oHIFrD3uSeETZ4m5K6O0h2vzLw3/DHP
CRl4ElQG4le+fYj0B9gLQ3jA8/clSGNC+//DTdNt4a2r8HO4bEUgr8cFRLmcg2uLQY4/+IA3DKni
A+7nONQXjSG6866XIJLQ9So+anWywgEZgRkDUIpR8gTiDtgr71+ym7TIAagzt576dGryWHFoe/s2
bni91ubks7lsicsvjRf654wUgwf7Z6zgbpIixUsUQfGBCtF+91D97Ok6JMf9nNTEcQ2J7BYYiZ1J
iz5k+dS1O+Ve6x/AsF/9kHMSLoXHKWaaTQYI/uEoxWtcTNdxaMZDhR/5I9k/R3Qr6F8RRwgGOMmf
plw4jO1O7Z+8cyKvtkOK7RgZfyBErv9pCF5LFnduQOvIb/Zxd8OuTxgCsVFQKsUdLYCgpbKLsd0c
oq+t7fpiKV6q72sdQk/YVR2C7sGvxEPOgIMkoOn076egbHuY2mgUuPxtH2uzkWaMLmSkrgB/74Y8
To6hvTbF8fAmUeK0poypD9OfFD/GoAU337bLBJY7SqxTNJrVjP+9SDkYEsU3go7cpNCE7nwxg42k
y8KOnZFzsnvYM4mRKj835QaPU2JJ6v5ibZxiZMqpOX9ho/UY0jo6cDbrc/APozuK5pjAW2G/+CPV
YUA/RcmEOtyxZesaOGlJO97zjllBOPuJxNCXlIwtaeHkgeV+4McfejmVh3JoJgjI9jkF1i/pb9jw
XigAQkeCA+iQnj45HOQxINwbrZa6FaSA1Db3eaxdnhfTrQOjo+TgWBCnjrZ4xbCM2KvDs7PTNrf5
MsCdOow15c7u36JGls6iMHxbk8JgYoxKyJMPBcJiYME1+w5hOsbup8Qi3lswzdafbiRezxIBJJKD
jcZ4+zM1ArunjQGNla6GWuBl2KxyZqCGnVyO+Dk0yo4VGmdvOcd6Q1I1RGVzbnKoCx+J/4EbPyBg
KdEGg3b/0upx+A54QD4RRdkMpqXrO+ivONR5L7J4ARk8kvs8w2NScBuF/UG2778HTCOpYWC4PSlo
n2AWklEsQNwj/olfecx22UnLsdtJ93F46Eq6MlMniP7UnOounvJt8/ftopst8u1VjzjjYDxk0KHQ
ZQBVCSwMPgV9/AKVUY3riVtPguwcDsR2Qog/Ik3o6hIPUVw04hp+nyxuL5bLZl+BpuAI7wV+UjN7
x5LMl+iI3JQlfYR14EW6UsZ1jk6eO2u7KaDIWyBI/NhBljFsYPrOkivnB/ZI2IZxpn07+5mVLSPW
RmhKMZMm3dxR6zjd/h4pPktQClLiNEQqt4OAR9UeyfHrLeDze4KcqmdcqsyO1FKSlPKHwf0EbKJO
IeNPjh08VV94OdTck/fS7AdM/5OSIfyWdsSytWWw055O52gj7xulM6NPhn8PR4NjnAcWWBDzRaWM
yGWdqdQiqyq9xL+9Lh7o6jLZFoLkgBYuzb+Bj1pAc2ou+JPc7aKKPvRsFl0yrC18khtuaxt2izLw
q4ScxAsmigR3GJezkzurLwpkMkJwMOa6fc7H0I4KYR6igra3J7P1ErA4GkgFT77H84leoOS7KqzH
CmWk+h1ba/JcwDjwxuRKGnu8v66sPP5VjBkH4JM0SWX81b2fxvS0SWzKzNOhLjMq0yCSNVeOO/4D
KJ9QuO4t4RR2sO4/tZfogi9RI1AcRP/GX6mBYPiYTtxneHJq+52CvBL4pdtm6Fthx61d6G/9BhnO
HMEOVkSLOZokpWn5qRTz9p8oM9fa6kPjM5nXhOcHEQSmlZ4/+K9Ug57wLPsrTeIWbW02sL70L/hZ
mDG308T+OJlT/dCN78kG57W3R8kZ/9UJOgy/7mtlhMUskgf0xt3KYxUFH4uBHkzs5Ce9WaLZc4k1
bt99B7vFhMoD1ENciU2zVYkKM6f4LE1kMCJJxf352bykKjCKXmN5Mu+PcCJ1D5cB16muJ3ekbJq4
9bFp6LklZW5QzYN1A3mtSR/GPMlg+G4vK4OnSlgCgMqC6Xbp6eJV0StcnKai+Zzkfy7RyHtX9Vc7
TJVtgeZVSyiycsDcFU3kDTOe+oTJ4wFg7KHztgtw748v5UUHylew2866lHLW1cGH15lmwFJlVQTC
a27ue6eI2FMl/0scyJVSvPRcIBUzKLKNu1l+2J7703oGOy4ZQ8Fwdp3x/NrpdRzHtcsJDnVWXVLH
ZegRuaQkUe4NFNZGT6SKv3KT9DggducPR4440PU2wQvvcZJzkVGBn23Nvzix8uxnpZkVtvAajAGO
vxVJCa3CMm/1EgWRbC8NKl7SluBMmv2Jh3xRV0XVxFL31jFzmjhxufmRW6sjs7riB+1i7VevAaz+
huoUtO30vCk68aBo31UfsAdXGhU1rtPUsO7DIJQd0CHk9EwV/eNfdV7qVz3a7OiFKXXPfIGm418W
E+kOMF15UPnhgJNi/Ha18ko3P/iv50wosWSJoszVs01yL7Ywdb8d1P/PmmLS6RqHWsh7JN+rvwTT
b4f/wHEz/Z0wSSQPT9Bk9sZyHijuvnQnrsP/6LGTRY0LtrciNI4Nl8lOmJSLDBNwQBIn9X7WkajU
zBCkzw+j7nFihg6c0QLqvcA6sh2m7oWcFReFKRMzdHfbc0T4VK++T3qYUGWuU87JKaDDKCAf3pNt
laZOvUDBJYoX0T2DSIeT7tC8jGjB03pZpqpO4xhkeu2Nf6q9a0mCfDR85QFqi9tM9tYzMz6G2JEx
f5eBGp+3Agid5gKj58n5g9JznORI/zhQZ+j8rHgD5/Gvo4Y+++Dzw5Do3QC6wFrql2Xc+kCz1HQ/
PD0cKxG+b75L9vbrVfEVtW7YKjj6DpBZBEw5Rux1cVyQk2YvW6HOe8FI+VBinAXqcIEk1OoefSEY
xHIaq/MTZdj5ZYS4WzhbgyaTsmcxqud3o9LgFRtBb+fZ4cm9X3q0CsrhVZMW36VPO8ifw2G3PWcy
bWoSS4EiXJqrAwrBzpDKTc8/K2I1BFf2unQWRcuGqoEm4TbDzVMkt+z5oEuFHm8NkX+r7wKSRwhL
PYZv0Y2l/tePHY2nrb5pRCr08dgXiGKub6TWlkJeNlRVNY45zVh1uEgT4hO3pSCAhqEttTOFkpVb
fBPai8Hgxl+VYuYCZaRUcDAej3BFix4DLJfj22kyhsbFwZlBaAcS3M52nbqEbUqsidN+kH5xuZki
SC6hQmNyT9kf8W/OlZDhpmBX54omHKX4O3ks0IE6NzPTuq8qta5VmX3ipn7VUwGsh+KUx+BMt9Rl
qsC4ys+LcOhmi1eEWq6QO5vm29NibAvI1cDikSRAvEJh6L21iDf3Hx5HvFWiU7+lmF3Xs24rZv/Y
yG9xHrFjLQ7POeOQ5E4vYOXUDtx9jDDPLRLx5g61huCDfkKMRiuEfTDLmfmZOwBcePBHWZPX33WL
tOdNe7SzBjEiOlWJzNfqPD9fWVxUiaQcYUVD2Hh7cJnmIDlTnLobaEwH1UvoFNzi2nOenA1Iivmr
ZPRdSL911gHedMZeUjRaoTvTfc4XgRHiC2uIEIYVfIA+Llw9FuRZvbB38bBePLeiqmy7lLSX7w8V
LYg1xBiVtK1uzgid93GjzUicZ0/EUJ80IcrDo4A/ARCtusJ73bAT5sSmGj2ZF/B/qavS2BKJVT7W
rheLcXL8wCIYyrTylHj0vHV0MSSU7Tdt//n9bTEb5z3KRIbyBOiOrALv1/Z3kqcIEj6XXcbOOZW1
GZHHBC3IFsDs2pvk2tdU7Mr7/brv1upOySMj0NnC0i7+UG2KdnGyMp6DLl2pR2L/BHbLN+9IGV/Q
emF2PnJ/UHYyXlFd4uAAcA5BdaBDfKSTTrVy8R8jVTN8X/RzMewT53Qwpm8MaO+uvJvD/7lKz63t
hGMc6Eid8CxdOLMS0U3JA0RqoiQNTTTjk2J7+Zo4V7SMY6zxsRxNpf4Dct91I96AyPZ05CPW1AbH
QmF6eR2u/oSBJCWDoehpTQMUeuuLa5HVBN20TCn8PaMjadTkLlAy0ukLBOYunelvKnf9LFKbi1o7
pu/7Bx06fb+6dh5i6RExnzS/rAolLG/7alO9BQ2O8vWLoHyH2RWe0v0f32yTwDDYsexSkpsuxzjH
oJIWU+wkP2AkGuIup2h0YzCWKCgAc4SRkernCUt5kQReXVFRhAPIhrAqntELmrcxoCj64S1n2ynC
YMFsA/ZlXdGEnDfopfxYs3+HlZaGvwjBLelaw6tphwVM/uZR+NmJDLEmMSVvMW+lrouOhEFm7wwi
udCkUmgfpglmJRMLvo0Sla/eqsyCfuIDOV22OVvKoypRbRmxTa/gNM6ipMhvkH9kWdls4v0ifw2N
dFIv2rOcgz57/KIybIxDhRwDI4IoimL3UvldHJX3nUu78JvYF78mEWdoj5/1eLkJhrKluqei74Gf
3n+BVZa5fr5WuqwSI/kDX3xH9OEmO/JLFDpBm75/h4JyZoWgfXTOJkc7PfM5OrTbk2bgRoAaH6VZ
Zf5OfrSMDJIY117C6VMgbMIIwvgfbr9kdqSp+kdAEzGDrK2eJlFtB5UwJPq2vHhofMaLBhh0Y5j4
IcfoJjAXu1zYMx0UaTVB5at4zKWBMdwsynxRMJsNji14UdygIqcOi/bxxo8RXjq35estmh1ZTlB5
EVGdyU5IUzApw2558T64emgdJejWQFD6kxCFAw19oyShQKp+c9hl9Wx9juvEP2KTAO5ChM2YEFR5
lRPO+/qOTF+IejcAmdYoy877I1UYfEfGBtIGvMzLNSRxOBApvvGYyCeqmG+BQ+qaODzAWbYjkDHK
zSUZHRpn5gKhVxxGGr+VVs2zV41x5LcPMZhPHrYriD2F6cPgKIPyAJ/vIY2jeTd3xAJnNRa1S9j1
5a+3j51TZJUzwX70tVRRNsw1DxbKrKsgtMRkjhLQ5o1aAnZpR7ldNFq0LhXpefrUkU8HCAarTpnq
z3AZVAK8UwR+atP+GqZztRdUaL6k2pq7IlwUk64TVadPsfkHAzHjPn/4ZvYbcCCGS/1MIbj9HYpN
twgtDU0ItpCtcldqZf4qfgjSeEXV9+0Bg5IB5DePSDFO7f4RwBhKiR3coDFby9UqyefXOoVqPK9d
KaXTH05JojxHHT7R0s9HgcVniexXBtQbNmjiSYa+nzOC4kwllJNedfGjN/adizlODr8kD/hpYqbY
R7Sf5Ac89bF4xl7R0xE7HUgXijF2Xl1srKk2ukNYuPgayaMddNdlr909NTpFwb4Vo0hOXU2kIyGr
gdJVYrLcXMIg1ZR+bbQK89hxtKQx8a75n4sNktEX7f/S6JCSWwEZnfr6VliM5XZ/LKhcuLiGmXZV
0HNvN2ggzYd+JxGnHJNBCA55mqHeKQXQ/bDuG3sNVetMuk3LxGy3FZg8nWvcZCWXb41Ez9oPdHTz
UlZFNXV3UOEdm/im/NR7DbjIJJtv53JWNqMEmSZwJZXerNs4Lnny6JtB74EW2dfGcSOSN4Q5tK9T
y81dFDrJlG8ls1YFNlUSlSlxFhDtTn7fcw0oSuRVUnJgoRKSb16qo+tg1E3MWpyz778iTgzBbdlh
PYmxaDqTtdxNAsJ+MsH8jlkwM3+bsfCfLPr8bJNBF8GfbU6JOioT26sud47S9ExoUqRhm8AUX3Qu
PuEidsbpmEk5BEsCmm4facxddHGnFHmmOy9xX3bB5IWuFN6+WkyQRWY8HNdf3Hx5KzX69xVt3u6G
9oG5u/xMqGDNvZMz4WrkdT5+N+D60NJYzWsiDPK4XIGpq7TFlaO7VknDqu+jy3u/I4XsG75AmmhU
sRjhwAcrvTLY7/r+1wpv1Jr5Zs6LpK5WXiovr7z6vMJhQVq/MrBWppDQc6a7h+EHxo4ABYLu6YJ8
/qwp7Hvv4Mlm0WfRHQ49wAmXH0htNL6DuPvKv7fUXc2sajt8x8soKaU4Bi3dYwHmob9Lc7iFhtTO
sVwVHoQKRSKrbkEqPmQZikEt7sPNXzmIG0kqhdNiRhQ4OLrY9PL/oHEVLI8TJKFdIOLWvoIoQEoG
0hnA6nrB4SPP4x0rJ9oDzA6s1p1mUbaec4P9RDeSILU1bvDysN7/FyuOqf9Tb1/8/hNca8BaAw6g
Mqr45K1xjfFeq675O+uooK2wzcq/ML3SQsaBuGyF189/OioIhz7eM4wI+tyXSgJchLTox1YJtJZ1
GVPBxI8E1ZbvBX4Ue4an6DxyacS15hbx86BWMgGNn5xtouA6Qp6digJv2F3wA5A3KrMCol9wrYwf
cbWPo5PUX1Hq9+0qBzwPeFQ2wT1029OQPScrEu9TWVyp9Iz53GxrBtU1ITmmPwJRRt4l2LyQyayJ
BJvv514VQzlm/ff3UM5OnhOGRXpAOXWWjOpJDdgR16uD137gFH5Hu5KHVymQI902qojf9NJ/yP/6
l1Gn4Ypp/xan3PhjBrP565vWTK2RCFJ/cnDdpqG5Kd5ZygNTsCOKApXa51iHonq7g+C+PIppeaIa
cn6+rY5jc+hfinulRliUqxtTloP6VnwYdJuVhX1/FLLZsn90P2uuS1brtB0flvFhRp9j8IB33LBu
APFQM14en0Nc7sPcOoGaxmap8Pu55Eyk8Ocdru54PS8Yer/k0dTxEy784XsNEal6KkfrjtFh6QbV
nS3xudQVvBrLX47ZvC0e9NljSZc/SpsWX+eU3WdECiR6LVJa+3iYnkQgWmleO0cMmNp/6ym5TVrZ
FH0PvmvH0opGKy7Rk7fhcvL4I0SV4p+ZSSBZkhDGbvxDXQ44eUvbDJj6reKQhWhiPEhcBbQRvUIm
aWp6l+QgulE8a7QNfX7208WTE7Zrqyk7B/dqLF1ml888QjTOFPj1o1Uy2EYw3PjMt5OAYE887D3u
FuKk9Pq6mu5ZAb9IP3vygOWM7s3dh4MwnDa0o4zLHjEAeuJPqqLz4okE5KefACsoa1QGemW0PB/A
zid11LiMg9EFx04i752i9nn4o9e4epgBKJMqmq1LzH6RNGEtcQAdfa2lcxWVvmJVSz4zu+APj3F4
XedxVLmM01q6MTQghg4/ZM65ZA68fZgxHgNkO2xbPkoOZbLqC+PcdS6ZBIKs/Zj3wZyKu/zgD40Y
AG6SX8fkcOidCh87T0iMp4mraCBy/34Us0CwGlcz1ISlHApwzgFtV2LGL8koyQ2j0Deovd+dtHEz
Gp4M2swlEk6KO3uA6cL2+Q6pEkchzbG4AzmyWfgAz7hCEh27jtT/Ih8Nrx4DDbYKCA8JWMUFkJ+R
Fq/yHqz8/rHxENYIgyFLIG+UURIQNh6BhkEV1HOqJ6oxIx8DPlqBQBjFPGDoCtkK07TguIx3yeNF
0PpYtRzG0362llHrqyThZdCsORrx5ultH6NK4cZs4YguJ25IkfFifxevGBdRm02M0shShHn3xBXO
t/1Mq66n8bSkkWuDKDmKMb7z4nHMSiBU2RSHgchOBj9BSP7BjSPOi7W5Tf+ooxAN23ryiSfCl9a1
9x08YCwmkZgd91TZiI7eBxbgghhzpf2QEWyLXheTP3yKWA3h+vzsyWK8z8oKqUh2bwW3ZLPYEHdW
vs8KlqLUoet2bTiMaD+/uxBpqH8+Pvy98ojRR/UNoAI2YuMgRnWtVAPm+EDj4aCjEoeedrgMOZCe
87Wyt1+qkfd14ocCiOhsdw/0zGl1/OeEZGxLS7vjR3EyVLKUr4NlXno8DGEm+2ogpnsUFDEu2Hqt
DbUIP+GG26j47TaZ8xtneaVPDulMClP2k7rZyigu7Kv3UYtShK32v/y1LV1WNPf2G3HzWZH2PilC
Fy+dym8jQsO74FpPe6jwqsLkfXgUgZiFwzknx8yMGjiG0lmL/ObZSNQ5vvfNryIuzN3O6AB7k/2L
qWa8tsrPOVB6gaPwf8Xfengok/sBawu2PaRPefR1/WwLNGeHAX2BWprg8h0GvBavqSet5nnAOv+0
UZgiBUpH2xzxqaN+mGLooYZOIoaF3q8eFMl9Hdo+58Ozn9rYGRMoi5AB/pXguL/pFZ+qv1axt0EF
CMJ2zlijkobMZnq7oSHGU23RANHCNN8maUKvpAbbqXmJtZRKdRTz940zYN/26l2xPBqamxBWprEw
DdTi3CE7pT7r8NfpL0XK0X6+CZkRn5LTm5um0a4POOyadVtoq08tc9Py3PnroSOUAeehDXua373T
SdJFDg0GElPYzYKyro+wU4RiiMUndiX3+9c4u7aeDgXP4sqwSGpTLbg1uygd4VwW8IBEq1JPk+Wi
esufs81MMukNYyne0XfevtJgt46f5nIAZppax3wCYt0nqPzJPeTjaCmOWDy18Kreo3trSKi42Bxe
6hT8wjm4TTmHyx3AbnCpN5yyD5O4gFh0vqO7QXOUa+Vyqa/WOoY+XdgLillPenZRYD/XK1mfpCN3
O0h4KbNNRm6uUjiOGu7O0af9Fcz9ROccJ2T3JzJZa6u8kOlQDiryZlf0GZzIdjLlODqTTAKGi1Q4
90se2FPVa95Ph44TCwfwUINma9v8BQSiqjVzAxRu90+W6CLk51ADmha6olMbgzwYK2WjaL9x4LF/
LiZj4xDFW6+DGQpOe6ZRVCh0CeDpgmS8BUDoOn53pVtB3ffY4pkfZNDgncGBgcavMFdspajk7z2s
QWqxdlM7wUI/XiL5hx5oJyIj3eI7Ns4Mt4XFUBGwIFrb3iJqh42V4NRJqmkARq5idea8d0CYxdNr
P7bRPwIf+rZcQTa64tbWwOeRWc/b0IAkSfUuMh3aoR6FwNR/roli8Gv3YMefborY8+F2afdRk+NP
VnNkBRrLUQj/v7AI0vKlCwbTdwD+iMxdV1e2E2K5ANDBm/BWqN6y7aPNSdxmJSKcu/T9QOIbYHEa
/LTPHVO4992WojQBMgNju2nirU0PhEsEzGz5ZMvHNbxD39+BzxgxzZ1lz9wjjVtFE5K/cKquNR11
5ut1WdKZz0W+ulieMwFLMgoAIphL2o3We9sg6ifCSN36XBKWQYghsqih0flUDObweOw0CK8HrGGn
2uCibAO90yWzB7UE4GHgo6hgjUaPhVhUdTwKuuHW7IYrXa4mxVfPGVkbklIX1/uLysQ0lJ6jt7by
0ckA7Cq5+dWvMvpqYcSKIUnEJ45ABRhap5QLRPSOmwqFRaOXi4utp8PORAEDhPybCORAFNl/8E7l
/fGv/m5UHp04X2GVylJp4C3XRhvZjkQnlybABRU5jjV6B/L//T3CDSgXtSMyovzDVIB3h0yZyytT
ZxxniqjdVco8LXDs9j9qmw00+p6V0skYTQWtEx/aRcRYNyCLcln+3Lq/yy3q4h6kURrYdfiwp1qo
RDSm7PZpf5/dfo6JFauAvZ/hLiAFqFDkDpd8rjHg7mrBlmuOiZxg9OUmCt9H8DolLUTbFHiknAfA
dCVT3XJWur07F78j/VoXjfLa8yTuDN4TraYjBJc9V0HU2aYb7rro1GlbqsIggFCAHTxTVhNNlTyf
O2hrJLGLFQ581i3qg7nOjPcNE4Y+LP1/uRdCmDSPPDX1K0gAm+7rMaN449G9fMZITnS/wqjBB43p
ZPIODoqXTzxXZyaz4AJAc/rRH5zwlzMtFrkuYBVq1/UII9cKTa7+IYQDgaNwRDgF61zVHnnnnHhT
/NxkoLFr5stU+7ZFkTecXMi0YtLwIWOZLr72MTjFWsUwKjq/YsTJMuMQ7y4dOWFN0r7GNas3y+kr
PH3lelrD97PcJjjorW1Iuj7lgSxbQWryUgiwKvo9wwjvlxcJTuw6gk3+pfBDdRLWaf/wiO30s3Ov
1FGcM0l6ZIzMdN+wpvM8czD/TqxWTSo/0L5GSHc7EWHh70GlIEtaSN4SlM/zQ7kkMYql9zuj60/7
PhesrwI617qfpg0kOJ3nG8uBzxfgjYxWyEN2z7ViP+vjUT7lgWnYT9nkPXbcwRwU99wTjP/NqIdL
ngXA1SYN25ZA6V6C+F2CSRsvEc9cTJKdQu9eTz/WUoop79HM9+P4aBjtAciZujmIFBWeqn2LQ6rn
eaXVHAiOYWYJQuwDzec5+PGnfFbQ3kvLv1tIvzzcag5qWYwE64pLKmr4uEyscQywM9NoqbvRxI2Q
tuaGpulJojq9JrxODGqUSKt0vWAUyK074zwYMBNEC7W7kZ6oma6EUss/XGleJUE0lJhlcxQ+Fc+A
TdvDjkGPwxD2dArIiCKO6e0iItpa6RdkOHV1SU3ChSfgZ2LQ4rq+7S+4Q0jZbBh8/A/26LU7f3kp
xja/ZiurGoqfG09tnqh5sAZ7+/h6s/rQ1ro9R6LBI4FnBGVC7hmrD9nVjy9KXQeysN2EZIPkJG5K
N45Libfu+q3titZSrmpYpNx649Wfx/nn5GP/Phpswx49EAzEpl+mTZH7H0zTYEaUvz42uIyndkIb
PsS3dOFAqK2nVl4aIAyGoNk/lvGADMd/iiE3O0idhMz10aV4pXEEvyR8Fzc17z8Rs/TXnwFx3bbK
Klnn6RVAVBfPHcGcEehgYzDCe27y4oq60PrwcKWPrTnwzj+RgOd/hX45EXJON2TDoU0vZ0iATTka
r9eBCop8ygj2leLWDHXqiL9vLsC6VYm9Ism2iHE2rILkUQZLIV3ppx/3TiBMyVVau3lsgUuPlDW7
cAQZc9sTcBvrzEu+0LUzAak2uakAn6DSw27qCbgrcdvNknVEA8WEpNF98+G794TbzVy11Eu/1mnB
+fKRgAnhAmHxN+6hawSR2ix4GnVIpsxuy3LquBEvv4Y0EfviGV0rtB42s5MjmtdmUH68POSWIxam
pXl6ivxn0CVCYjsWGzh9UBxmA/Bd1AU/qQDhe5tG4p1SaVCbfOYNnUbs8hK8Jv1ald18e5bnySLd
zGscqdDpZhAWXeQrrBMa45LTz7vKyjMxqEM+ebz7klB0rQvSfctXN2osG7dT3GK7FkjCR1SsdwPU
AsEqw4cemcsUsZTY9t41F5Yhm0zECk+Ob2leUi3joUj7EhwztrEnJ0s0wMbV7LXYyHLJ2X4ywftL
13YOWkDr7qcDFV8ZUnM+1iNHCpHR+3/czZKVJvpx2IhiVopaaz0yUQwjJ2lTcm+N0IVDzQCdjHE9
trQTBPmA31VOFzwfovrs7wHVyke4omsiveXCmH90Uyeb83dE6jMsPQRMrnEsk2XGefz+gI2Szv5D
A/3Gyx5ZbBN0pAmL7fY1VPdWHExOUTa/fpGMfNqV1Pa6uL8mUe9lQIOKJCV+QOBg4cDdqUxs7mLo
C8r2IdB7OkuDN6cJGluPP1ugdEDXihMDSsC6ODhkL4/M+TNRS+nPbR5/5T3mxsPZ1tbZJZyjnLb+
DuKZM24IEhPWpaXQ4CVDBx+xkIX9YCtt0wyHvobCt1FSg3Y2WwDitM4PrpUkpqQR7i0CjT1tLCbj
IFh/miQ7Bqwx8xYTp9dBoINPN1Ka2zZOivLPlqpWqT964xasXqhvWNOFRr6op/oeR82xcYIDotyK
xumAfPsey7+Y+0xcCeKUJ2DEY/InoNVu1omV0PDa2cUSHxDCF7ao7P46Nga3aQithYa75rRy1qpV
FM07miU1nkUEfeplWEgODV8mCCPRm76tKb0S2sjXeMzSUltUefycbCvGL+V6oosLGIlh2uZHcyoJ
0JQKNRAgay0/3CyhH7qFwTIGMKNhuAZb25wp0NMW8GgvmC3AurYgFvl7aAhPxH/rO2S36EK2Pa/P
njdCFfXPyui9G6W2fHevFBBpYRxwBuZZcYfjPCfCo39X2qpr6hrld2wyFTa8o2EKEAuULYtUMMfu
dMWW82IYGk24CDfLUKr59BV9E5UhJqT8Eax9O6GGQKBzpV7RtOZZb7eppGEk/9q0MBHyougqwQeS
/ErD/FHlbjsm8piIFVEUD22Ypd4vQRxjuoVcgHMYG5WO4FpM6Wm1A3vFd1bplHXpiCALvOn+3sXa
FYvu8ts2eyPVA0zrgV0lKIhmtHNwIQ1ZSf82U2Eq75Mee/N1BmSb/igP4gYX1OSaX1yW4jp35PVq
NI3G6VtPe0v6g62A+0rq5TO6qXVENUVfX/npkKRCiR6RXrEDFZNA1CoV8u6OAK7DnG8wIYVv1XL/
MONQCy+5/RGUrokLNZJH6KxDwv2qroTD7Ckc9qCOf8lW2MBVWfds+WkwVS3Hh/VGUviwbNEtbZG9
xhSSQ7acAoJa4CFxL5/yYQCv/jdHSttBXRfblEhKp+c2JoTsTtIngoL3wCvyitldyenFCKGZ9w7D
rRMESWYRGa+GAXpa7Fr4/XhjCCyINABDYfeqidKzlQtwmX0OBHZz4UIhShQNEMiahewMrrhVgEgC
bwNuEwQSnxFvuGdxSrfBXtBgAWX/7HJFwQPjIxujp9aCqH+RjdQfU8a/+qAUF/Z9CSx+KqTWMlwv
1ge01o6btgsEMwVneGfGcyE9bkKRj7YGKcxF+va+v6oakzGDOVKEuLJdt6XRQl8SrNk6uBlWA6cP
GiRbJXCndXS0dGWHR3W39dCuBS/Jnr1dtrCe7px1A7FU8Y4ivite52cMCUtqhk81pfqsYe+FpeAT
FDy0WBm148Vkk99sRfXOpmv/ggm84YHH4Wy+yzH0rzPhuVQSVkBo8/lO0dijJuZxcDXsbs+Vd49V
lGLhGZNpyIEXB9ahjnos0MRbidHmuHNNDijxAkfcH80eAA/2iRPy7tiIk3nwpSyKwpwkoWBgwho5
ypeT83wIe+KOaYBV3ENLfhnAOiCaJwnEFQRMttNNMh7Dl7WmLeJf5LKg2uH3oyE2B8LR6cAiKYGg
kCQzy9S3EouHlac3/S3DNpDRetcygbKjEZxqCR1EN/Rgd4A9+vs1Ac6L0S0xHrH2WvwH6mbxrI9n
T4+DpedJlwscH6BpHA7n4Mh2w63grd4S8LO1RsxWgtLjaap1fVsZrVScInlnC15+Mjvwikii/YUU
ksnz/cVKzxnAsqrTWOZQ9TrdyXdYg4z/kCxsBsrWEA04Fsw7VwBgovdc1rk04ZJ7Y934DdgO/vwf
E0EhPqrNzmt8TBCmZD83K30lMagHeulx12S7Yut51KnnqqyGOFuNMUsTLvabykxgODK/OfAem+OR
/H4Qp9OCnl0dk7gzilmrqh/8MWrXqVMTvs/wInfUaq47lXBD6Jojf0A9FTIOiV+6P7QSCudMXzYU
GWolBfkc7mSr5+UyBNuzKzpSA1FUSg/4AbqdY5IPtlyPU1QPW2T+mKkj4oTEuniZtKN2oUDwbp2z
hxFNa5ejWb8X+A5GTz8WSIr8+YFYDjSf/LWJCkjybOCuglkxkoc8gwVTN5j4JmI7Ueh8ZlLWOqNb
8sX4AS/FeEElH/GHvAt5Lq2xIwhFfHCINrxEJ2n8ppXAQF7vzMyioRmrfu9fdugiWZpfqiWP8dXE
RPSiEiOD0pnF+nqXph7umBzsjTZ37T/9TuwLhkoH2aS+Z9/0W6G/dqjRpGciHzH4xuT4mLYJH/Cp
ryyJ6sgLBwUj7/QJmmTf7RUvZkpSEVGNARCjvozoe9UrE9lVs2eiERQLt/3apu51clZqw3IcTTPd
5zA+ku2VaFSZbmjFlT+RzSaUg8tZ43qZpaRIwaWBpYJ8lYUcvd5s1G/iw2Pw6TJvpnIRybKgrDYq
297AvU0OskYUIU6Ce45A/53jhaVsWlBgPBYm/vJ1ruZE1EWIRh7yQclloevK6pmPSfLtDmaJBBc7
KWfjy3BWSMoMBfQ84vOLiX4mU54ORsjrRtaZAhqzugL7ePJZc8JW4N+9TSmYiFmNFQz2yQI25pNt
5ko5o2sdGeItr1F9b9ee6qUPWI3nD1vdVegqPpkc9g+oqS3BbC4Tx6z4/N9WnMpqdmTc8L+9w+AR
55CI1pw2ugVCuuL8Mwk8GFjfdRa+2aA3YtRhEk4iKseVsu93oSNdeU8aSxWE7u44GNkV8OWI/hfl
kShyYCezh92q2K7SL31FwBbvahc0ECiTsOecWUidC436wPABxVOdf1pT0An/HuDGLl+8obs45afF
7K0xYl37+ox+2xSOEnq3nEcBh8DZ+vnTuxGza8KDc2HgC3MciDhJ8EfBPyNa1r8Zlqr7TZ05Bhi5
AeQeuNtHvB9JSc3aw1oFwHkFN4u+jckktSyPtFaKo3ItYZ6PzU5886/VZGif6esnWhrGckSoeyhB
0kXRBUV/p94+nJle4d/h8rE91q3DwSOwBmGYddJtL2RppQJW/qbHVriwExvPkAPdwvIaqVfbn5Kz
DaocEaId2b+1Aoa0Tfxl5gDliPPLk186a318vap6OBk3IuRe9WhuHoJxELQPWwoKMkbwV8+TGK82
8GQTC8ejkZGI6VazKWvwJ32cqsf5a615GmrVph7HxGie6MBJA8LTBMmUYlYW6/Chx2Xpghgb0czk
Q7rkxjNlJTNKGpG98V/j4A5u2TNXgbEIkE5mtMOZlZgnQfRhvakCmOM9HyB/w+MFrFtVMbRK7lC4
AfPqwnT1v0E7fRdh00wU7PS5UjtmONoI7wLm6WFl8W0Wpxcl7e3Nd9zEIV3dj079caXjxc6O47yt
V3ClEyPEoBwGuWLI9AmDeVWF+1zGNnQqvcLaTgyUSKRYMF9fKfZSvwp/ZTDM/iBWDIa+8kbrNtt+
22ni0hjbU+dVVeh9PIQdU0TSxTmODPMLPjkdJ8bRaEfj74wLOhr4meijjpcboNe31C+chImkZ5m2
8QZuH4g0pRbZ/Qv6Sp0ncd/0VF0tYQkmZnu2sZ3oHkpnS1hL224gK7iNJDW/uY1NmN2ZXqNfalRl
X+cV+4TOG+MmVfJDge+Ki7J1Jq/ssLRNzefIXFyMKXJqs9aqWB+sV86Iv6QbB8bJLzSAu5TOaxPG
uUPg9Br385ifo68dIEdWfG8xY8m4iwD3AfOY+a06xMAgEfbhJNdftXvRykL2gLgL0LJ/WtjxyVJk
j/n8NV3dFj4S3yEIzuEJyL5PU5yIPctQGGPMjgn/tNc6njp6dmdRxNtXO+qIJ2lvuXBq4ENKvrgm
kR4qLjJGq7Vd+Vlt5e8Jc1J0Q0nI+WO0UEnl0/wds1q8rMDME3RUfu2vUtRG5GLWvG13U56Xi0Fx
l5P4LMW3umjVBOfBFNM5lP5ILyhEOwR7hH3EBhd5m5jHW7eng62qghyufwITJ4Q9hME7D2MGmPhW
6qYMgu/JUx/QoTyCPAYeo01GJhcMGq6cBUAdUF1/PwKSXRKJjDb/CG5dm2JtdySTE7EvPYOCUH0/
4FPkBUn9RwKfHPoRmvxgEYLoQY2z46owRuvLZxyHJkrj28u5fDz+S8lP0WTzBxJzeHNoXsmmzZXC
0PfNiabha9MrhDafjLpdTb2An7Hpi3LD1+8jVdgHj9xxrz33hgF5UeSPYwkO3qWXqfyc+sGVEGTq
hXb4k1iRmcb7TO3390WP4XFkzcB0vsTUeLg3WYyoM+QspxX1gKNfvGuBL954A+7vWcQgeG1V8EJv
my1wnLAG1iKkuFsjJXVgzr7ltjAMf13qT1kWe+R+32l0NP9RzKWcPJ4SLXtIFDFHmk9jx5yi0l0T
0V7KuF7A4TeGrOIPRQo5a5OYZDH2OJKFuwgIBW8kUpanXZjJgkn/zmZOwTdObrUX/xB4r49ynlW1
f6iahv3BwCWKRguqHL9DyRYJhx4C7n5UVJR1REIkEpxd7/Mrtg2EqgnkThhWi8NrDFaFVr+I97XF
P+GuP8Ep20Ycycbk6frhVX1OM065VbVeOs8NNbWtsuHbVwxD8EpYvuzZIai/qO+nPj6zmKgr5Y4H
XaEH6thfoOz5CJzV0ZSAd1o5wAvDAt1cSK8IFP/Y4vDBtnzpy6apwsi6TSEe9GS11ZtSPbm60hX/
JWn1/LBIV+3/D/7+oNcOiL3Mq20/ZYb6AQKPwZolzxHcPJlTHlEjy9Hdq6UjD0o/Du+Tlau+6AfR
N0kKr845GbXJ4foMSThhNf0e8iRP84Rr3FD7y8kdeBH2vWgvbvX2DywADJI4SegNZ9+JpNitcjYM
/+EELbOgFrxayJ5y93fiacWfsZOJKKNIYtZX0nmIz2QhAlj7X1xe2xbDg7JrjaXIAaubzrOXTXJi
Dxh/n6A15GuQF0ChQjh+k0zo4/3w3CrF9PKVnLvwcX0CEvR6/H4e+5EJl91UwLDC0kHCf00KWBEs
4NEdPjSeYYwBtQ/YdNr+7I1x4NmqCWaIbOa4d+bWrNn6tIULXM93I1LzP3TWcLjCHsHQl6EbaDaL
mRV72Uy4T/kGMpsk932te6HR/RvQnIgn9NEbfJxcGeYRVQP6bzG7q3YlaliGp2AjniGPRlzICOip
0/KahZwSD1t879i2Ez7jp4yJSclM5SSNRRaI19MJqPqh0mQkvapIu/zurrp37FKtcw75FnSYSEsw
CHkSMaFLw1K4XrLQB/skbYsKwBy8xGHjpHAyVi5afWqLKZRHM58Fjhgt7iNWUOGpERdeGD2AQyZM
CxFYWUI7WJVItrBr/NVJARnNxSgsmI1Nv7zx4C9N+yUYIBPdE9FkfuI4ZOaGi2l9PL5UAU2ioGoA
3SLyoG6msgvscXV2BuJEJyqWpfIQnGVN1R8fC1YeF4kuBrLk7vX9At/UjMDVfdaRpFl7o5B45am8
iavE7qiRK+LAmuOusa9DfCCAYbtrRa00Eg6cIBw+qsSh7XtaU2qLlwNVhunbPDQuYPHEqnOrUdp5
PKyeEAksPTwPRMrpi0wz51unieXCufg9XFzewRp9IpT8JPxVbU4G8bvCYYxSUCdVsyFIXchzS6uV
vW/qCXKvnMDLj3nMeCB/bJu8PAxAIReziCj6W/mTmuSfBF+t/iv77Wa1myBBVMeb6bmdtNemX+mR
zKLeEiba3Dm91fxazVcZL/vgAbDNpjs5WRuiYWMfqMd29eKONMVMVww8CWIjkb6wD68GteYJrpcw
viO57heYjapaYqRyP9A39d4xHF9jvee/pcHU+G+z8WU3krPJUkxbYCsMTTnoX5yMFnUH0pP294T7
08kB0CatpbCqPv3NC2cNijjymyNPpsdVddzYw6pRIvulRU5aDrlT52xKOQIasTy9SkG9KI/gqcLg
rdWUxpF3gtKKVw9gbNbimT3JnVFZldsLk9MQu3o7H08+AMzkbGdsULrjkisuQVq86TJaGilgBrdO
6PAEyINuDamO0u26lPJaW+NOMoSGIZQJjyzL7s9s6he6IAim4mR5/Hm2IaldMogOeewkAgdMGPmj
lRYXdhV7Mx6YT7FuMGtTOHadOj4c+8ulObSdPhIUwNMZDk3blOQ0UQJbQYdfAm0yC70zkAwmQ7Y5
bVyi9x16G76qdQVlkFBpu0Ye5RV/R4Ec2vGotLDtWPLh2J0sADwDUhE3uNlTdpGx3xl8lP5hwtwY
H9LW1nTCZdBCxF8nQmXPUCIiiTcKWBtxEWMS0H6fgF2YzLQkjD+i+I8nd5+7fCfrVTbfvGVKpu3M
/w03DxCYVVOiqHCmL6lRl2dmAxbfZGPrYvfwo99c9oqvbDvVgrSHjHmLbkOVDdbbt/LTUA5CbQkq
9YH3TqbV3hSjxqLp5VsFCkV6YI4y20yZSHVUgUis62vWmYUvA6NhqFeLnPpVvdtQCX8O3WSFBodQ
8Ox3i0XiB3Fuuy8quZ1H2lRHBbze9i7E3a7vSEWPs0xoAiNSbKs8ow4bztfeSKtCOX5+oCUVYF3s
0QROd2cBgD1vsp9afjv/l9T6R4aAV2rt11gDsmlOqlKxSoSaU0wWE7arWjWARNkkGk49xhfKdXcS
2QO0BZwNKfZWkI5zJ5Ch8mHp0Sm3UiL/nZqp7DWvnGxx9U7PITbBJRfCahbqVYmwGdh7LRkuCaLg
/LupS7jvnlLZzqGOZsqwA58VvZVjfzII9oGP2mGrFWU0wwrgwNytBRBHnr3cNvnY8mPcGcoyWEiv
S38XWmF5FtCK5bnsBS9FsLdjUkoNRinRgVmwrfPo8g0C5xmP94HIPm4JDDnSB4GbSaTaEarsNy7/
oTxYW9eOcMWrtclXRvrTp+4acXjmyLg7wTO3XJjQV2cveaE6aFAFbcK/1yu2C0e431WcJksiIvf2
7LfKzqyJagj3fpJrxihjcrR+hhmTm/TPz7ibJ16VEpEN7Alf657qk3h8hYIYIdbc87rWyOuM7ySB
wSwTEW9kfUDU5GwAz2J0tZgbYd+146FP//VHlbDBrlpxQat94yZzAtRg5CgqxtEH05svk9iFoMas
S2PRTD/VyRTR4rd8Mj5B0o3TcAUPephailrzgJweKA5AN7uQV4Ebw63AZmA9v6QDXbjRuzDoi+wF
u0V8rCrFg9sukEzHhZpqmq48yHYmAbydKdo1ZUgNsPWk98/9/4BsBwtiSa335B6N5W9WPtSFIbAg
ueGzCIKYRZy5tjHZHWptm4Et6kgbDTQyFcBg32u/dAz+oxMMaNtyAZVvW3b5tRc8iJ93Fb5o49or
JCD6gfPsUFMpc2GeGiWk6Tay8ajLNp16YLzboY2Ck2JajQ5U0/Rb14ZIrLf7tttzffgGe7i/jsku
RCa9NoZirXCsuZBC0rqBDA6PRBnPG9IpyapcORoLg7Kit0bDqNMv/aZtO5s05WL1ywsqr08R+sid
/7466CUDmgFblLEbx7H2lTWllmrw4Gh+GMcNczVQ7Sg8eSZCT9zkiRcaQ0RdJd46MigCiIp+eL6h
WIapx451U1/WPpT3zGXCTe91Nf/iiDDBSr8v7FN0lBv06ujv9+ZC0JBablzeBsa++FWgo2ftZ5mR
PbJnkE3tSVOt84wc6g9qdb35puZ4O6i+1HFYnjBC+B0uQHzVfCeseg3c9rKUSLgxnSp6ny5dWcDL
lh1xsyO97r7NG9OwG9IK9FQdL7tooM4oGEaBcO1iR51ny/rOPI/wVVxug0fx9G3pV4zJIf5XoPOQ
yM+EBmJSwUdhL1cYnnF7SSeQCSYUTLUyvbNUkdiuzYpfbFFtbEtPXAWS2UPhj3sRySrbKyWJIlzd
kpa0bHnmhYHtBXS6EmulQkMKrfg9Biw0tWnLTotk1QZmajiO+Fg7sIHcMH8wA7U3gejmgHAqo2eC
Kt7ubAzzD8bapeUR9rhCjrXkH+piZvOwBYhPqnK8IHRxLkj+pg/g+/lkiiSo6+LV08onnrZM+DMS
AM2el7YbcX8e2xNgBeIOTafq/lzH3Vd/g3pxWIveqmXJBFgHNanHCY4lX2gHjdzNmaaVyzMsO+7u
mlYm7OpPI3duBMlJIxHCKM5PNQGM1MviFU4b7t6FwNM/SB9sHmi65ySQtXm921CzWmpU5f8dyEu5
qQOvmzVANdHcUwTn6ui++rurszhemS1m/FcoauYQfCab9KOqyZ9HIxXSF0m5vMqnWipJwFlaEVj1
M3+XgbOi5sYqLDg3yuX73PtjGI89qSN4aaQxxjxDdE2S6OTAGKDeBotK6UhS6NIvMiRFTgw9QdfQ
2kVrUh0lphzQOtVfrujcHBynaeOrkihRuejgDiLpfN+DiUZZ0PAWPmXQg38x2nBGqqnF7h2mkK9B
DcJK6wFqX6FS/zW7IKWArnq0J/OhhUmwbPSwILzGhqSSYorx+3CjGH5mvYY8gw1+JavdDBKjRSlx
2f26wrmXWENro1awIrGzWw+pccz/ihem/X1W4ManSpNJHdsT1R7yEV98wWkIjFJtpFjixL+xPy2h
IyBNH6ctRba3nXQXepQvOj9rm2ZNGWmuCS9bspGQ8AswUus5jOBF46eSLJxtXpL1FWzTHhLrt7AJ
0uQmK2nAzaI6+84jqVTdj8+KWJO9EmXDXA07Yga711wWBrrsG9tzJ0Y019nC36icteum7CU0qSDx
giN2ISOC2Dk3VIL6pZUha7SJUwHI5+LVx/K4KN58s4JUhkj3M1IJ3/87itov2XkaKVg8ASeYUTSw
JYL4QhZiak0yzKx1ZpF3VndfPR49s/0pArqC3LuR1kP8hOOLAsA8KxqivGli1qFw/d9K5cLdXGhM
dM77GI+R/FiJjHQ2euwdJgjA2XYEcpiSTGH9+bO09X1w62L7lEiSSVcSoc633RCEHj/FvOVNHB/4
GfW0FEDH09GUOFlVrQkgSJ26+OnxmNKjFvTxvNtqPNBGwgzlVBLCvt+OaE2wdNqNQtgjxw6L651E
6QvvPbONvS7iCdcEAEo4bgEDDjRxGQW4NGZXNtnKm+RpXhEaqaZMyPyV3oKXu6u83P/1EMcVe/Kg
zBOUUAH+x6u+CWV5eNMc3cxty5td2ViqAxWNgHyRRK4CPkxTFNtvCOBF1arOXPI5tFdSoyjpzY5Z
QatKadv0htgm1XIXUxv6hSKdbSYn8VKlkB4nvLdIn4/yLK3ImHweTTfg01TGsoAX+ztqR0V+nQv5
lxjpunIC5hN28im7Fm7i+uP4+I1rfpYYC0xVbrMHpb62/nkHMDxS2w58WvS61Y43+ujlezyo67bH
p9Ib1C0udsgjW9PDTTkYHlHwr/lTGNvM0oGISTXNWk3wJl/4UbA24qyj9Q5ouf//zckOLdGDr2Mq
k+sBx56wUhOpClwKQ7OHfTnIq4rD2Mnbtquvtjkr4e56TyGazcLIw/Sf7kb57NU0sewBX4JUsNVf
ATH3IsXg/7yJlKb++bbNvf+bP6y1f9XPiCGkM0E1RnqVdYgj9HhYEgj2HxQdPVl2eYFPUTfeIaJ4
tzEnDZB517/n/g5pWStBX81oigcFPNqkEOMnBrnCnf+MJfhXvBVUdWY3jLX0amCyvWvLUpOD+KPK
T/6GlYc5XxoF5f4ItPjy4CDFAMytjtjUiSffcEpTwARqJfHMpZK9OiU6L2eujbZFgfldmHY4QYuj
Um0XQaQxf0qD1lQaMQwSbmrvtW/G6DdASe5ftwoiFkD284iLhg49fB5AJJsFnSPmCv7Wf6oIhVcv
U5n8jpVsMBPwor01mBVW9ML7iBVUc2t4BpVGlKcPUQBhLpIjzAIn2vwMcMNeSskQNh/0MqIgcADq
zgx97qmcuJqY++yCUQbxyG5q2dJELyypzaqWkoNBI+6tbg5whg23mzpqjaLU404zgG38Tb/hCewY
j5Sn75gGD5SJzamHJEP7bRYBC91A/JfUhhWN0P2h1Be1BBkJf2gENnZDPJQ2P1hGQkBdWFW7/sH5
k1jhzEj1ov8DeA7l3JZonctuw/9DSpjOuIh9+L6E2oNGYq2iyylSViocqoyKiLZN6EDmgUOtZtKZ
0oSioQOdffmrxzN6wQvo3B3BCuVaokNLuSF9F9odG07d73mZnGxDo0W7lrBvXGiIgbWZ3A5ldpXQ
iacO23ehGvQxVZrYlrNo0kskvYJ7mPlzzQOjLfiJwEOmHvz6lF4v+2S++dJ5BHwTCW/csOhJA/Yl
2sikdxVXvSXo0jkUXwDrPXX0J6OlTubidZvr0yCGJ1E4y4Urdys/7pekZyaT0ptoCxqWl0gFl8w5
Uyjnmp/hcV2P8GyBrK9cWUV5LGGJJWwVO59kBby7CoMGvjLrP2vWiztkK7FML2tWZWWU5sduCRlL
vBXoPvfdgge2rZcsRih97GQLLt8WdLm2m6NhYs1M1rYL/Cz+bKr/5j25lvUQAzoNDwb6TFylcJOa
nYbwbrqjAPWU8nJxeWT1S6anYWoULDZ6J8vQ5cWAHisPKFZfA0jyLSRFMBUVEs6P3OrEbAlOBEd6
znO36n3VcOSH3XFeb34NcXiXRWm3CgHoEp2OC/R06bJRK1b3+l/EG74yiyKIfg9KzAI6J82CSZ7t
QUTp8C+fMsDdDBR4XWrpzlWMDSJICujQlZ0cGqaj+RfwugtDy9TsT7/QWvg4GNTZdvDjk31ykusO
lfYrg+ytt0Yy2pw0V2bMiHkRGAOlcXkcYX6tqQ6d7fs2BeGTARBjFJ+s+4nc+X6XWYkWxHaR7uhL
DhZ8cH1CemuTHQeSGDTv/l9AOsjZGIislu2dZLMEFBVI5lTHGYgPJsPqZnEr0re2CAdn6aR/STPl
1QP/9823grBNLaBhBDE0owB+aNaDnKjBSnkk2CrErgYoR3lsqzbMlLRQLdE/gD/6JNmVqCN6cuvG
0JTNPuAvMVlTxdJpd4ZUcJtX+nVknpZdn/qoxe2qbgqS1HZEkBLPPkYQF/EbCxhVBK8HRUV1Lss4
DRkv2wvJ/iEUjCRAJ0vyCXmZVibZiGFpLpfqT+bKOmK8Jl5PW7tVWoBYpopTsi1RJBZ3s+Dh2/Ql
eTXoD3kvzsIWSofaQDXJx7rBqJieH7iabEDqQqv50ai0twMFCoJDaD5clwQhC2S6w5stQc+Nm/ur
lt8XxhsO6fQEJ49pWSnEnl/uoerrtfeYabOkhfBrLFip9rzfVS9adjckChU2nlBfXoC1xQXPSH/O
a955Sw03O4D4WY7XLcQmFbDoQ5ZGfmEcDbw4uWgVA/QwUt75Iwp4FiOs/sC4lfmXXHyfEMAI9h8N
4hFsJ/mBw29WX9zhC2soFSMv0LKia8RagTYXY1PX5HTt8ogRuB6brwNUYirpyF9pH8SHwr1bvh3t
AGEoCQoFN8qWPozVYzgzp6ai+h2tJVHfWyRRwUiBc77TlkkM1ira57f5OKl4WS6Vyub4K8Dq7MvJ
cfb0xAAGSIT0J+qCOs9Bh/ER3rRZj7akreiArGoBi8K82JhkKyGPDp6VFBMQsQ7N/MVEE6h1GXmI
WQA1ktaDAzax/xDmW8HDTrdE7wPL35zNJSpi//ymiqN2QqEF9qbt4wrxel2WDMqznMoyrVWIUMxj
NYfs4SdT1dC7cv6FgAz7TF4++oQn+WeKpuUR+ZeLo5AwrcnbxHG98eEs+tVQADroOkN+YbrT78do
08bZQ/GuU3nGqmhFwhMWRQFuLgucFdcvfxuejiXmKWZnjV2ulbf43YMLkdYAQudTvqqaALcXEg8R
r23tmcQF2Ujd2Anwy8wm15QYMK3lq6EX6FWt0LshcOCuTTlNj3y4uct5AgRVzIjOP8U0fQDoilhT
qHz0SI/Kgw4VyheIYXRjuhhC8Tx1zp+2OxVvzIL7lAXs5XTpNMUKNDWGGccBKUCqkx+/3nhr+glg
7i1WdhrVy1zjY9JYbOMUGEsCszYO/g6Afth2aqqODn0st6i0xe/xjoH9Q2SvNYLde3NrwLmH3yKc
pdXxUY8k+xgR7dAIGMUA/RshBj38dHtLvwTj9+wiOThs9Rg2DhN3zu+VkkwRThaqkUWiJ5rYTa4d
tJEaY7HNUYVzhAQ0bBMFNnRf4uqMqQoUC/8RQuF2uKTYvnqMPM2Lg83c4Edw7NnRMjVQWxceDIlx
nhSqwFcR/a+k1CNBYvUbTJ2KFzuBeIflP8anDOjYo73fejR+H4+jcEZiTsJxOurfr3mL65Usr5Le
INx3jK6FqOWbdfAIBHRU/mHji2vncC3gbLDox03BhJjFuuNT1Ha259OmupQF1SXO9J0tn+Nxo8RK
tcOfxwC3QJcNSdnOLQTMSg2R03OxfQmsYecbk7zUQbruOFFris4rdgZGQh8CB1mWhXZKQ/Ioh9Ze
Wc5GUi9b3COXF/Ubj4XQvo04y0bg1zM75jsjXY2E+/NiET+l6gMgIQKco1BBgB1qhnv5ECRVkQBL
ho6Itb2MNNMjfLKoFQotMpGi2E5Rw1gyjSgjEIKLLhBQemkBQ/NCbHejLKEHn66EhAArwyuoAFpL
OJbi0dMB3iDocLCnPMcjI9ku1NbgBtPQf/CusIPMkWCVVIwYtCuMy3PIz5+8a9AaWcIXYrbWsR6T
ZYzAIU9AVkbl6O+mGc8kNZgGjr48I8AovCVi0JSnluGGUG11oKybg1sCxC6F+5KNiTn/gjbhPJMZ
UAXl4eS1eXMg6UWZxHN2+ebsVuZ+CxIud7C7XzWwb5WNChbvYoXCJjBPi2Ur23ZRRzrnWNPX2Q7m
5RV/VteUrdphsv5NXmhXm866vozToYHvNQyqhKYxioLRCagy9LSiFNM7UrnYjEnkiM28n21NjXKu
xc9WTvFzue0xBW9Zyu+VjHHRSrXmRid4cIilWDnPxmCgTuyQ78rrZh41Z2v5dQytzntuBOBt52DO
d/waNnb006Bx2l1/jU2J/eL0hPwBigwnBN0gUmc157Muc8vVO/nPvyACIA9siIInu497N/PnOXXI
/tUWIMtgDRqPo1GAB4lS2hmhVmIkLug2zv/n2NMvvHvy71/ttpqYufEFolMGqnO3enVp5Knw9LCi
tEOuDzwuCSgrZLVm7uq1vl7TVCmFy2ujRzI0iSOaOp1bGQx9EM3AcVAcIAFyevfvbOY6avG6SV1S
fF+es9vv7v4EmgWyzVrWmuLwO5OddxVjsqgHkD17jYwwhlLfkaaGNyX8Rov6FuM6dgrT+YTepBTT
E7AuqqDvb2ylhGDSFHRElVmp5DLmjrtK1Jv78o6kRarxzFyCr3PrO3IFuvTbX9WGBQ5borLXj3qu
clVPswtuzditWVuaT0+s1jQWuAT7siJEF+5VJ9d/Zh8bxtbOzBS354H9+oTlaQkBn2OGZLkDcZtQ
ExVRqVFzMyfICzoXx1KbTZ4PXcLJHfz/Imr0rGEKpAzi1yq8BMwqwIUQ3jEnK8BucZjh/UBUBWvQ
qjZkRVgvVuUdG9Gcq31clri3sGRK2D3HPvOpeXHdxnpP5jYD8x9+IKLIUjrnSCBVMDsV34Va+4Yl
t2y7zOxw/GkUC1G6+K/5roVXrjZmFfXG6EnsHDvp87G/IsPtyVj28XC7iDQzgN8rwpzBsEtvlrsd
c2fmP3ZtFnUep67yvhHTzsYwxYKy9kPlZEd0tDvHyVVZvwWZ2KLBgtBKtN0GphGTI74mEKTZfKTN
mP/gsiP6WYrenWQ/iE/bQIN8xTVOGlUzPAfZ9qwMlvabVwXipWwYoZsvQ7wvg6oupMZMCZS7CCh4
CD6S7gNngdU7XUgpCEvbQaM9gO1KnUIcv9SpJaR69lavXs3dYIhogHB+K2LBwAA/Mb7orh72SAlx
1MEhuIeBzmbVvuwDFTuEGeREw9NewA4kSZqI7k36ghn6piSD5lXd8fTp+AXmDJXTvPTAbhSiN644
yGcKlxsH3sA4N6Os1SGoBMEZ138zIlwjp1MBaoBQ2ZLXjilOvmBD8v177iLiqz0H0lsgqZiW4MsE
0sxE++0KbriIUtPX3ayujpAM+vBpWVngZ6iBAD7DiP+rpmz2+9pIaybDIcUuQUmiWLW71qatR/+6
3k3yrW/UZfohYaVRFDjISf3ealaCZeSBymaELgc4yvuSgw2dwLQvnAIpoic7ZoBv+X7D9CkUwjhP
7KrYhbQg9e7qUOD9g8PIPOzyQUptSCzecEYneB7dU0bZFSl9c4NztcQ1hF2HoebruLh1TkEHhIUI
c/z7UgzwemxRGvyC7RV0oDd22pfNsN9VBoicPhaRzLtv3e/SyFRrOqY7m0iu3jWV6hk1esAmWlRE
Q1omcfowXjlKDLeEozIJL1mGJAFiz8757xUc2fJC7HXrhbW9WROQ4Ug0Khh8e5j4wH7smpdxYr0c
eeU0BfKIIWL8Y1dQLcAAUIz1yhiEM0C0Eb692l8488bH44zkEY9XmI0Z/JX8v0IGf4T4zDjCZIpw
H4VSFVhHYpqAGX79AI0K/fc0x+ogSj5iXlFnYzZWqJ6/mhinjybf8C5z8Z0MMpUNw90K91B0uXT9
5gbToqomWtVAm9NGXtSfYSSmRt/tYl5cZTBFPjJVJ1415AdJ9iXAGuy1WzG+77k3WZyuiDr+YsqF
i+KJ4iL5J+4UQLVO3zNH9/2LjtKxxMAx7MftK9OFhGKTbN9vHXwKkNd/LSRTZkyhry0XNlBRz5Kj
gMziuA6p4QonVSym+e8b9COcKtXgtvfUAg8SFkF/ey916xOCWkpCXbr/fT27UtQpg8hYNttA27Sd
1NcdzxwXNvaXDvRCHdgYuZrQa30nVz0iVEAqI4kk9DaAVH3IvlXHsgwKrpajuRh2LhWQs4deyzs2
5p+ViGiq+ALtqR7AQEryXTZiSvxrnwQ3mcO2jmeGVouT6JUco3ijRxBwQntG7LVNdftkxnnHgYP6
9212bqfC5F+2X611jhzHDKLq5ZU3tPAgr9/qGM3I5QuycDlezOvyop/M5osnO23s8ki1vDGZnlAf
OnXuwVoC6Rkx8v9E5FDwWftvbOCbfVYizjua5doYdMGJfLMnrveJR0f6xpUcxI7j0K/bCVWvSf9T
OXlkaZDfmsnLgPxCiWr5UqB1QvLOyd/U5dhusVxRIcRRipVTxza7vJv4UQYoUiICTERrecfws/WZ
2+k+tzjiXKpatxZRWIup76e+pCMGj6fUAcBDJx4klRDuo5nfOvwv1xfJKJP9mqPLwPgKLDVrhWZn
NnS5ciT27lmudf3aDfuLvMXE4RM7ICHcr4K9ElwLB8TKJeRyvhPrN7TG6/swUuTUoMzyE3Hr8QmY
GpwT3iWGLZGPtBvbEm5lOenWiwxmr+j0nragFJSJqXfrFW2FHsavDTzvTbjTczwHcjQbmmFTt9WA
fcma1Gpcqoo2JKBffMJrg0WazfFcG6ABlGANjJxSIyiqHpGK7cn25uP4X437fAm5vwkQWizBjaux
A23cYLWVwlgIqd9/0tCx0GnHQ+Nn0rQeQDlwbGGI6k0orEoViLiCEodrdxSKjCANCosGuG+M4WH5
Xne4PtFL9FKp71PDdLe6T8LVI36wv2nashJIwtdA4RbYOWhcG8cuESAKu+mt73L5wXcLaEEIbLNm
b3IsquD9wyrlAOcpRc/5IakN8lEmtALiFsuTcDuP3vqXwRU+XB6EfOXu4J5Z0kw9mzp3Yn5IyICZ
Ebv4rfcQlapqBEgK4IExoBJIuQ29gT6U1jkVnVdqqvYD+iL2ODdUjVyZDgSV4+ihNL4P3xDVeD69
oag1UAVkl481zg+wyaqtqPhZ2RL2/S8YumWe0lDcVW3ExGQDA0mIh0SMQ95yk5ahXmqo/K90TgqO
p5woGejOA2zkx04rhu836wlQvRdpYOG6Jvt7pviHvnl/8rSyW0TsFHCxq6tQqNzcvLmC9O5dd7SZ
RjFz4gfNJykM+r88wuf3TNxejVAfdCywNvDElmgfpWxFRcg1cALpT7kC0N01vvdmT35II7zp2sYC
yalCYvcKyQ6pvtpP3HVE/MyXN7TgPvIMYHp6ZcMHpuaoUtF4lQC8MZc5Dbh7eFt7dQGs+h7GdRxR
FhLQ3jZaXfHpEEObZr2S1L3xUgoZ0Np/FgKRgdcjtb+KKRALIVmMetQ75yx7AV1njkrdpkB3pcKf
nl0cTANlLdhVExe4NOIEOIpNUBLOt2kalBDNk9NrI22N9Iqr7RXqf52Bk3rnsg94fMR+l+jnfHi3
WwhdZe8kmaw2bw+Gjj/ph/5HtGhCkY3ry/Dk3eyi962EMl6uISFIMcvwjikrpb6BExjH2I7J9+BU
fBYfWV4e8Mq7cPfelePIWpv0xrIJ1nJPb9N1a32mC5pHbvaxAtje56nnScDKDVUwT5BGM/TwkGBZ
cd65ga7kCPm/JCi0IQvKwu/iDpfsvbnTuOiC6gTTQ11MFtJKYVucycbLumfL+bAii7Z2vx6zOP4K
vAjmzY+hmnB0fIUNWURS6zT194O+zg0Wfor7GMKyuF7sU619yhIBJ5NAudtkDxEt3VqeF1j1x6Xj
lzVZNJPTvBb4ICuCdGPgqhWrVf7d/k01C2BWUIY/mqEL/K7CBIkX18o3YNmDzMj97A3C3YWpbOam
3ESM5TM8Ih8GeZAWg6wqheCvGAiCWAJP9+z5ENRF7JDPnnsex0fShZg+qRm11jdrQVg0jchmcZln
sP6OhrlPHSw5mMqosnF4T+nLNBnARpN9l7hcJDk0M9Y64dSwLAMNU8mfqdg19Frjc6nqCIBAb2KL
P8d1QyQymLW/MoChsE4YsQTNMVo31C3K8Tq/xEFO8QNzrAjJuP7XLTTIYw7TihK1bxKac+kHyyPp
1I6AhTWul+jg3nfCBiLpy8XfezOvYE0YdUpvaXU3ddSGU8fXwpakZdxh5dKkJ7K8FWQ6qR7gsw95
TGrUqEk0xVT6ryBbjTDo8J70L8Ot862s3JDmX4fCkRPimNA+IP81m24c/oik/hqmWCwgOUoOcdsQ
Z5k+t1LK8PzlvQtX6MPPTAzONZcrueHYoBaCz1tybIdlSUef6nmsDuseVvs5EQAtgkxsc1VITnhM
0RgPt74FGHyacUT+dKnQP/m0S6YvFZpoNSF9sMVJ1PBdj50DaOPSxneH5vV9rdvjD1JDtvTfXoUq
RUE6+ZV1ZI3dSQrCG3MnujBfQ3aY528RLBp+libNCsWcDRB/VtT18tVfOst050V/o59Irn7LvhTr
/6HKpYptpPhJ4Gazp8uuYVKKrc/FRgwQ91NN6TSj9FNUxFcHTOBLbIsKBBiM2A0xFLSdGTDPn/ko
VpzG6QhLOAxQUK3qXtJHLqnXIuZaw/kLsY5ujojhUMrOnrznT+kd0OZ85seXutM7YfBs3/IwL4IE
VLOMlO7IiqZf+bW1eNq6oOTlYps1jaAbgwjbkfs+UpR/o0+LFsZLvMb0+1vF/esk8SUrkzqhtXrn
gYqPg5LthQElcDAwv0Oq/zdWcXgp0SoY1uZpDhc5b9fX4CB09Z0IY6GI7fB8IxkSfvP62HFk8hBG
q/UoEDb6mhX5YHfeOBW9WOjU4dIBjtMUfiZkLaMUk6EnAgooHAKYPn4t3NSQ0BwtNZb+bmyFI2PZ
sBbu27qOrMXVtczxqUIVrSI0D6yGSfA4hP001cXGt91uVZJBacc7fxzmX6A9fZZaW+tO4mTLl8oC
8+r6YNo7+lvuogMK/iutViXf3FDYMJnyisWL5ac0ObhskMG7pP1ooD/Pgsc6LX3dCHnCG7nwLg+L
irgj809JGA0a9CcQOqkxyVtD4kTVqq6MeRz/wqMRRSW8PqsNe3wMV7Dos5M8sbVKTaRwhXgAvJo6
TSNolEmWhgOZkcaIyFnCkvYyVT15aGWaCrUjt21zm97jTzX1IaEv8WBNXvpbToUVuyCCgNxS8Jtm
DcocULbJdrz/vYn1abumCAMqQorgwi86AoJEFSXocP6f9fWNnzQMCPNIPD5AOMTwTdOb0ik895gQ
+1jX+vrSOnBpA8C7LaDCt9vZN0vcRvDBx4Kg7VBGuUcHbpyYdI/8hN11kntGejvL4/AFEzycDPSz
I1AkjAM7mCc9BU1uQCxcqqfm6+2jDml33zQShc5ATpVRVPHqC6j6b6QWS33edF9JT2yFUBMaYLQS
N76+1cpKH9r7+kTkynkE6bd4xgfYxgyNsZ8ArFYlXzJrUOZnQFFXkBgaCCa0Gtn6i/8nu8prINnq
SJutSkqIvWS9xjnhYSoF9m4zQJRmXlPFj1IJ8ztJey1uKrfOnXm2NVMLJZffEp3NAyZVYgRLIgNd
kZFGgjuyhdFXiy4cBVW6/IPHaGn4nIbJ1dbVJHK7runDZVXXWGbhV3hi3aWb7wVNGn3hfv1jRKiT
We2gkwX6cN0qKyLDrOUd51LNtCJAnz1i8ayNrLzQ10rHf3TXbWCI6w6NgH7Io6xi5X1reesQrWhW
MmA03Ryp1F7uh8ENvPk5qoBmOxhnLLTU1NBPYU50kECH1vRcJHllfXsXrThafcHojT1S+GJCkBSh
9XprSnBUCwb3pvclwcRdGHpyDk01h33Vofw1uBtmH+t+oD0bIRu0952PxQ93QD/87S0tEIb/8uIe
A3u7SMM/VyMoObDACsNB2GlagnxY+QmQUfX/L8kjMv4pPTGvqbSkAzzKgU7yFpk29XpHbLIoDW+B
m0Rfe4FML/PvnxVM0oZvg/p1GIXWXbWj3TtLX904reuB43cQNeRp1NC2+f59aTxBCIn+1UsvMmNW
3NUp/qfV8f+nvTTGngXOKi/iQcBunt6ij7Rb11KffGW/E4fFF0k0gwHUZRW9biKPzo6iQBVGa3H4
P81+ma2qawNto45KuOdLlC1LAHFN7Gc+k7fMpa9ObGOuli3Ut4f4lLOuBk832NQ5HMMtRIqpFGrT
zjBbPROS478DgfGftT1dTLSVCGPkQ3Zir993Ly0LW53KbA7SdWG1Xs50xFIBEzWdPZT08gHFiO6Z
7UOiM0rI5qhYhJUcIvKXqUBsXv8hXweuYzXXA2FkPi1lRYpvSdT/4zxmhkB6JEIkip3YW3keuM0L
WKdEBUog4bAg05OTDY9EjpJid+UtioUJKuxz8fVqAZHCr3QUGbVZXCCNJgA5VaSq699PDuce83wH
uxLgCh/0pTgaQXMGojIFo95UcRM4BdahP+ePSQA6aL6kWD6n0HUNPY5QWUniMAx6DUAvHT2N27CX
EbCPcPbJWB1VnOIqvuogGo1X6V8Sdjhk7Ix8HBk0IdlevjK+o61ZHiQH1p0bn9N0+pSJGlNBDJcL
xXnj73GOpzdHK4SfKj3MWpgKm+YzFB2oBh+zWuc+eefqxPKxtN2cQCnIim/lGgpfisF1bnJHc9S2
Gggde6+uhRfuyn9W0o8vVFPI2NAH2rpubhv96bWHZgT8hNeAMm/nzqVVIoKgNgzjWOhx0cuAZ04f
zZblkMHkkULHWTTCQ12SGkoIq/auY9nhEgvZiClGoNvmUvLSbtru3R9c0FTigYYm3RNwHXFOZBeF
l9w3Aj2DBoznT/28hXhm2FuSBb/Upze6aDn9JrDrFNUNGChMe07csPIsarT8xK83mdeGYb/1cB4P
qsCcOCqrZmjm7P6ELzGD3xzApioSq45/ViI5wrX8kEdQ8PatYgKWIDKt9kZCVAYC+vV2urfRHyym
j4kbhVeVY+xVRTYmLaIuQaPvxoIXzdRg+nG6qfnFxJg1nJO3dNKBvcTFQH/cqyNdtvR+Za/rGGpE
vRx5F5cDUupJaseZr5m+vBagVZcQ4pjUajN6xFu1aeuZ9ZztxZlNjLt2AYs4zxK7YVh+A4mkHjH2
21c+c3w48EbdHi98ChjsxF3/3o921rbb6hjK1S3XbXYUmQX3ssmGhKJB1m7nk52ilw/loQbg+yCR
DGBYE9dh+c/+v8LTMMXS0ozd+FCIheWzFzUj25/4zqBCDzmZn9nMger1UDugyHExCJ4zgg8Hd3sa
Khar7+X2b3ncBiCZcjwJB20ZxkRP63MbxJYABHLVt2GXra0nszy3+zryCaWr4mDH4jaM3zkhvw6f
edqNxY3CExc77TkpbX8EEK2U5vqP6CC31OhyaC9gAI2w3V7IHGHJdhlShUaiLoeqIAFEAgP33YPk
DCyqWUQKVxUq9T+CWTxtXc0V76a3qGLTp2A9TfLYi7UnkW67Ba7JGcrBONWgNljQ0DTKqOjpaCsa
p3+N+WYiZtNvccF5FlMoMdBnBMvFraVwVN+FsdQftUr5G1eb1Q5cQaAZCPHv21yCRaVN+CixeNA/
7oPjG46x5Kv2HJ39Kk+K6oU0aet0gPbx3ESteAvkXzfoBF3Z11THN9dy0eZZAxAVmCxVABpH+THw
VjMGu/QvZHa8Y4JJzyX3YK2zSt9v6G3zRl/H5xDnF5GxjHOyio/+7oVmRyTeJMe1OEw+oYO9d79v
8H60MT4kgujbystz1Q7ghqnPjR8HXI6LpRgey5q0BJK3gJPTNUGCGJWFedlQZVs++GfsnuFzk7LY
OngQNAfDE17S8j7Bpkd6D14V54OhdkLtS0FB5XFzTQ2NC6hs5yN0Guwnb2fOohEvHRIIp2KwLOPX
eIxOJstWDMNEHglxeh08w5eUQjiD6LqaPL4SCexX8GgR5caj9J95QQ8a5814NjxmVpN37xZpbYv9
n7JM2v4qTzKWw8dXrjH3yxbFPtrd1f5PhQPKklJbnsZjYR7nphzuoFhvzT7LOcJpiKzei5uHVRKE
ym7jCb4JuKkV9IjE1eEGD2aPmv5tdp3jxiJhINF+BSu5X26TPLFBoAGr1tj55es6rqylaiAqsQmo
xxRS3q4gVU9M63WxYgVCA1/C3U5ye9W5/Ur8HLW9wxA7OjxNe5ixitMSgNV0+JOG3a+emqigtzDq
tkhT1KRyWsKpt3TlIzdeuzSljnpQ91EfAxzDNWXdDHRDiT0XTtkW6QYykx6Z7NEzNy8yZW7EzEVn
+4DTFgImayV6QUAn0cwaartZcyx2xLYBfiQ54snS7AiWX0weN64uXAvUQfSbRb+mZaxUm4oV7TO8
hFMGG1bq//Xt52qZrSN16cC3FPoT+q1bUSZo8NSeP+r5CCqo5ss6FQoTcU8BJhiENV97aIG2WPlk
vTRmrUroQz1ez0TNyNN+S1YnNLYsCn+hoRov8kRhZ2qriHkhp57p2BCMlzbsWcdmPB3TXN8cI/q8
irXCLVoOwmYUVc1JIJYlKDtReRYltS1Tg/W0DxSYJ+k9p09++vmfVAaFWned+5Y3nVCtSDbRgZo8
a8FhFp6mbBII29dWX539viPSHhIBCBh1ZFGe4G0d6JJm8SB+TszUxdFDJqX7OTPz6cPz5r0ECxqO
rNnAL4NFp6eP2Q9vZuUSXOnEDcAWJJalFbV1BE6MfS95qvuDr5Wq31xisf4ELDY3aLb4W2LeFSwS
+uXk5mBPtTYfFXLXvVMd1KYxEyAi9baU2VDeQWzH633eL5P3ZvsIYNLsNbmQrPPby13IuvlcmEXv
Jcw53nh135yBTJgiWYeNu43oRbPDAGIPPfImqSu6bBjApsA+2y2BamREwv3I563oKHFhwIDBcJTD
C/u1JQYXcjdc8ksHfuvxgdgV/dYQH+7aRkx90gCbYsgccQeSAVBQe/89H63rCwddyfTqLVegPaLs
+8P+wSokAhRH3XCbJaR6SOVz7N0dKLd83NprJkAybmwounbgWJgWUfY5fEahtE2jciUmINGcsuR/
afiLobd6gkNT/ePICSHQiuu4nlna5Nhjjs4bUxMc5ACRoZN808zk2e7RETc4mQ37zIZmgvgVhq4q
OvEMk7d2x8U2zRvjb68mJy3qIUK34r2CbfWEvMAF7Itz3TVaHyK6XpWCSBlj3jmhUxXI1YobF48W
rdJ0jjnvmUaDQk0MP5uzfvCvurBjkx4MeId874U+xR+jEGrNxZl/QS9Yo8NZ8KoUrOuU4fXRQ0Mb
XcLJQkM8Fe2jJB6BqAM9ZT7o3JT85c+OYP2KT364Nj6AVMHmm19mlfF4ZbgvcXh/KzWAdRgwPxRK
nCxspMoxPyLAihbFDJsknUwS5keAyb5a0pZPlv3fS6LGx/sWlseSVY++0kF7kLU9EOGjuaCFkEOn
a+qhLJuZVVjdDBeYOxVpHE+K0ojyjEYtPg5fYJwUNWicf0GgfroYCB5bPZLIEaTR9cLSEqAi47u7
MfXljZzTIONwmg27N/jrzk2IP88y+8/7G5DJ2TGXsoBLniu+j0kgapL758BpTI+8GHFcOP3k+3T1
27IPIYqvmK2+o5NDgCSK5RJeilSfTcrUfv1rQV3sRiiMyRFi3M6gpbE/feV/S6mlhGa4w500Gn/Q
5iSiiNCr9RGP6RQjq1dZqWZLYh5er4N2KeU0IxFKa81QNGfWbqYIEPMmDVNdgIY26Ee3jjKBGfpS
3j+DdYM+oeM/iXQvYjD4MxuiG4UBboeFKTzg0Vd4vQ4+MA8TvhC40MUPjRnW4xpD9PRS4tjYlP2y
R1YZ1KjCbXAzrGfHvmlfRljKdGpSiFUc61JzSXRxTDhzcOxe+xPyDicEYEnw0tJ3JYL3ixrkFJ8/
yrv+Pfm5JuYqgecKV9isQ4Nq6Hk866bfUH7pWkhQhzuobnNfn+wtQlTzRaymJXiEMkuPXiL6P587
WznTMbWnC7qyntgOwBDwRez+nPtALUnPEJhU4hZhvoKmUgLmJOPZeKKNRxRVlhygjq7tB3fOfV04
WMB2H7yW8b7ARBh2FzV5M5hY4HK7Sfh3gi6xIX36AjeZPkpq9L7BmJOEFcFB42TjgMvBe9sAg9J3
iYkjtRJJvqkRai5ThYMRzJOJ7ruMW0CInvRJoKugOkCHln9e9fCbnosHTD37GgYgTzBwRTuLMEu6
Y1TmVnaQ2pflgfnsO60Ha03BLmErI2ufY76BMQl6GzzVU7UMpQSNtmbf3Ph0ISckZrsn0NMmQXAP
IT8pIVIs/6klDagwMMkjno7/RcPwEpVEzAOKSaSR4gaCTkCWG0VR+hTQrGxd07agQTTDDI9jXU0o
HRls/ai3BB4obOubSF7X9jzv0/D/RVclF8YPakde2Jxa8J55mmHZUdGJQ0zQlGOZhxOse8J6dSTr
dBNEgLdZODBPfx3rn8+UWIdZWg3oBdFqYRA5a+xXfVinYK7ZK0uzJZrqM0LA45LtSxVDxDeKgvKj
QVdzOnEfc5/DuTYi+6kLH8omVUyvc/BuWPoVQH6eX2BEub6xYQ90s9xNAcry3WdBRrkyL0Qee1Q8
OecGwT/T4KyIvGYz3vT0sNgc45BQdFsWuh1tw7VKaU2BP7xGnR15JTkDxeKKhHHK9fKW3JwnwDfe
WthsRdVP267end4Y7x7vSqt8f3yNJbtAhj50QUpJl4NcgrK3zygr0U8F7O0i+/SHMW31Fz20pJkI
Wd6GYAQNOP5UUk7cI/NAZceN+kgy0BGIHDdiCM5KPNh2o845lV5zWMPKSh2jeb05EIwUqZOTZlTA
gqJCu/jqLI5vUW5DbFBt+G+hzvd59CPMwHoKw++vgp6DkWMssMkCbqBGTuW5HcR4JPphjPyj9lQL
g3qz8Ai2WLNeeIJ6B93MUMFcEtKeIGvPw/mu//c2GLS8IBBPOGKMpl4PRhq0g6zPLylTzRKNol+l
RJm9HESX4xnAc+K7/u/Ytwfz+YwcCnrs0hYuP+zd0/bTttpwIBSK/Y6Z8BoIl7xIbWMKqD8MvS3S
BxvI3zv9yh2aFzRKwh4vr1HduzXd8cSo8j5bPaGyS0zXsjDct4NzcH0UKGnw8NiXEDaR699BZ8q+
7pl6QDqS3zyVn4qSCfvsggn7BIy+EQvdQYmioRJHAhaUqR5b08/fU6CogWVhEmjC2PbmfAPsPcI3
M/HYLmF5Kgj87CpgWRguiH4Rj0gTKOHI5AAfNDOXKb71NaX+NjbT8yaH9/nNmrTExCXi8Nxg8Osm
0GUWM+hAPpXJzpaDTqu6naJI8iwcEOamA73raoigwPk5m0vqBcwkpn3aTDtRJzZTdoCKwcmp7wpK
/5SkjBlUQliNoVO2F5aOG6GDUcbyg/rSnfSZYeMt+iVIyZBZ5dnvzq4RRiDKvA0MiDTujAiigMt4
ym5jxWtEjP15iP9q0szx5jE1tX3PRCOAfscN4SGr4Fw8KHsCC014lsfNt0QUiQKwcSiwQKmI1FOl
yQb0u/P4s7PBTw5xdqp2urCOLDiOw2a6WhhJ8b4tzD9JK5TFb0W16n70hYe5wJEsZwQJR0KU5AXR
XbFcQqUPJXUuQHFZH5ZVYJ2DuNkbXUSXZSKKBmXjDVbLMEKzwG9PZwRgdjlMVAk3Umop1kNgF2Wc
nlChFTHpBBrMJPRW398NTTPZTt52zNCU5dqFU6FiCdxssQoSIjycH+GiNZgLqUAQ8gwkE3L+lQDk
ZP/SkSByu1t8sIY6WpYYB4qzV3KnbZFOu0+OBaoQ8OfEP3I2CNAURWaUUu/zDK/N0nyAvVve9FjG
FyAC1hzFI8ScgyFsSmciIARITYOhOtBwSSkeRALp6FcecO0eTqrHhMCpbUjcUaSoEPUdYPjPt7Oq
xn4a+H/A30/CfUK8iPUyHpvZeFaZOqNAg54oBCUqnjK3d9kV0Q6vwO5mHrVwDbWY6IsZWSul7JY9
hk3C52wUSknR83l9fgfI5STRJgndrwLVxRyylWZUL2nsIgF60bicUkARBkjxRzwQWHD5eDWEoiDM
a4t8PEsJ4G7bYl8vmDWtu1PxiLsNqGXGPp1tHbqu1Y62bCveQ/J/sBFD5zspKLCP23o9NgZtzkHT
AxaA4ZZbkeWXVfe8YVYk7qr2no+Wzc7M2HXrE+VpBVFhUv0lmjTAGUrqUgQqhRjlZyDiaUqmpgkp
wbhYNjlh05jzOXbpk33FVwu3lzstpXPUzGYNZCKRA922ygg96C44lw19F8uR0MJNa9/aIURV/rE8
L6hj20MFxa3PYjLl26IHrFInZHrIxFyHiET3K9q2PpZSk+1IrPn296LMtU3PKfwNkulh08V7tmMU
Niudz7SX4rd9tZcF+uWy5xoU2Ui7mWOyu7P3aK2qRP06ywcZzIqnTTBvVutIUiwFSWWGIhB1ikcF
blzR6/KIMwvF9VtiiYFPpmgStTC7Ihe0mwOjZR6t4yLFQrPe05yDOhE4gCO6hEj7aOXI7IeHiT3T
SOmEAI/oqyWF0BOjX6K/mkQERtbNIPNBtk4PXP3/g/vxZUgkEw7EuoKxiBdLy4DrlxkdKlxdi1/u
z3LE5BCmZdERvA4itOV1Jw+nc0rOoSjaG4GPGuPhcFG/716SdXVV2JhaF2EmylZgk/et6qc99sCf
t5ahyxk8SWlgZE2vOpBtOfDDeN6Xl+qA+QoEyZPfN0XHQQEghaGjar03rlb42sxGVm3t2sh6OdFW
j3Gm6PGbTd5q155CfyxltCo829mkfOuXu5RYeVk4UwWR6MgtSjZOzJp3gRWINR7ztMbW7JSNoXvs
0yFY0X5yLIGJvm0k1fP34jgUEOk7KIPQwc+pGC+zVS5jL3PUieQHa0W0wbDp42okHcUE7qPEYSbO
m3+XjXhirMLSpJcTCGvRnfSV4Lo4znyuNI+7eZ5ggay/kx9irrTIFqhE2ZNjR3WtJ1Ltpjol29VJ
xpHvomOumvcglipdGoaszYMSRlZNnCH918dsVmV9bO8d24bd4OfZ8+YS4Ggctk8fGNjE9PCEDUmp
6jgpHJAhJqywbYVeCH2lqA20oZgXsK+qbwjQw3sSEcwmzRBbYqmWbQyTdwLnQfrw5d8XeiBibebN
4+GMIwfvmjVMBlCUOgl7CpSbxSB61UHtiky+cZO2qyCE5HsHSca7GLzlNkPJQt8byi/GIakueYkd
bibB6nctJ/wk0bSzqvuz3tlewjkH0HTrC6mQwTiF3tiADswKwqsuvP6DU/3bZVqEN0sAPeQU4Y7/
weGDMnsQ+48L2c+pumw4k+Ux22fQQQnihEqfovmvLxWBByu4SAmJptMWDYgYcnx7+Gj73YprK+f4
MVj8zzbTzV+NCxr/L2wAb6nm3gy0SEepHuSUZn8DiV017ojK6tPw9hWsDUSq/d6MMaXEfd3A6knR
DBrFI+X7YVEPDj+3g3a1vF1hv1eSKl5CEZALbWpNF5o7QHuSm5MS7A0DfllkTyIfdOLQOtYwBqgh
j+Kli5plPp6GxPoxWF7eVVIMcqGpfIODlfKp72kBK4LszCVj5a4JMQFAha5A3SjqMNYDw4CeCvG1
OOy8Aunw/GDCH1pnUkj93qO2IFMl2WVJK1As48tsTTu6nZdAf2ZntJEMIFqEyCz81U+glAi1CblF
sLEltourObkCDl4G6Npsh025yetO09uESt+ldIXp60+8UNYQT4Tn3M2VAx+DEdfL0jCozkydatmh
l5aEZE1EbHn70lwkI+P1hTo/92rN9g+iwQdXuUtVbgEaL2EpEAGLhquX0NUfLV33G5w9wgDtPbT3
GI/DpEezG45WAwCD01jQFzkTVx7PxID38tMmme6OZ38sGsDuDTxjgVYRE6W89a7gU+vBEe/vYweF
6ErnPNRLcStLQOC04Dvv8XkqEdmm2zLxSM49l3C+Jp2o49HGx9Ci0ZFB61rxXFqkX2BJaB6sWGYt
JKzkrK2otovI+n6kjDc7A65Fu7lnNxbZ8y578Wio7hRYMZ0Y5Uhu9IeV6c9uXu70uFxADihvkweg
SRHlYr0IRy8GTLtn55D1tZRy9jkKHOYM6DqU8m631uPmigASEuImFXt6nP4+f9NViYosaonDLaif
u2ehqsH2TvgEXSjt2bUG6HyPtXRGWkMy0Kc67bxqnQaTd4mYDbTNX5oHv3n6P4xXtC5AOzi4gxxh
9Vu22mEKU3oCiP3EehiZPeJ3NQwehEcZNYfF/rUcQ7+1barckIFNemTxYuZww9cVX9XYtP/WDipi
e6K2J09HYJG3Locr1sKpEpnrXMNZDjK/sZE8kOPKleyShWSNjTa4TjgzJZONZqvt8F0+d4A8tKof
WLjsi8IV/wpNo4gT9ag7eLKyt/ekhszFt1dst8vawCggs34c5iNRYIiTKaEv+83M8Uasi/1KZxb0
eXPrGSKVn4+T5DgG9WaeVldctViZ+lG+yM468fsmvI69NARcY8WeEKY5YWoJZe9c4vutE2/3MFOB
RHAU9XFZ4h96E2eG9d2rBRwTJz6V++LecK1XIpDwcUHXNW6TMjHMR1EA3BbHF21vjFq6yd4Mba8D
xqn4Bv2Q0DuocnSW91v/xlrUq2m48hUw/BM7oPYzlL2ipz22rmHON5oQWBugmix+0+PuOiNoXM4t
12s8UNCOjpbzRu2VuMP4nOCI4DqIz/e/n86hglcn80qeuVEIpz6DvWLxRxM6lMz/lkONycGb5Pt3
ZE6thVFGrd091jmcZE0ys3J97VXh3Y7933MysXC0t9h62Spro5ZZ6YCNo7EUcsCJCs0Te4V47xfG
Pi/NHQYd5KVYHJDxb6vHxux2dzs4vup0BOO63cVRtYEU1rtfb1skMMorXCpcaJuZ0pykzVamw5bV
L1WECkmZ1kwNKJBQXCsFRS9ZgELfxhppGG4KRlKV9H3+Qi5q/kvY8H9s1RocrZBW3yxcpLM7g0bx
U40PgHc5/Jl5lDT1ubtPGjVirD6WVCrMDRKRqH0N/7ev1JjFR5uZFtxJavL6Q/j5PhP28V+QraqL
3+u+QVdpy9/A6sSnZEs0ucL06WDjM1sJPBXLM2fWnwF136y6nJcJB44JFSWLhKtvanTDoTLTuczF
gWF7tBgf9Q8/Fym75mFP+kBsj3bbQ1HHMpYqgUbejZK25htNo6ibRF/yLmJyXTXK0VTsIOPh+0Xb
50M7RP0RsMFTxJpKKZcgIsmi65H1I1VM0HLJaMvnUPmaR8Sm1RKHjMBqyeY8+z1omIfnuNQKVHc+
QXITKtBJLJoAmYhlepli7GnSoqi2UhN753+uRHud/1zl3j/wi/A7bCtgBaC3e/cz5eavuZ7vHerp
z57BQ6ywwC4O90EBLLOkFyOfMhlo9sMKN1/dnM8JDIu+Ufs3aUCgjmOM2cjhPG/e2S6EVzh1gezO
w2cobN+VyNr2JWSao9ZS8WP+XzdvBvclsRWfjJMf59SZMwuWle26X4rUEfAOaRWuNHkUbD/PyTrd
fZGzK4F/dGbt2hKSxpYnU5R5cChZIQ0zG7vUxikYM0/5ZlRUW/hi7eA2zGQ50XLW+c+ZvCLu9hI0
iWSrOIOFNlwbARPtGM2daYTWq7hAj32VowOwOj+DTemZnjkArVFc4kp8NwKB63tpJEI3zA8wCVmR
1+VwY2pLNbhySXCXeW8N0Ie/mbNWowETSNOGebCDRZ96YFaKDXXSYaX/7wQ0CRVFlv1RBEdXzVkt
gcGw6xkCXJaO5LdKl6TLw2dnA1LWuvMPRzWJ/kQTLTGT/MN0rOUO4JBAzXDFYVzGC3daW2vr/gcr
lg9PuYFxX8zWBo19Mw/7ZmXAT4mdzJdmRBENRMOlNSqo4oRdcgbd0hrSMztNGC7bMc7I/mXICPW2
2ycuZbK3Tz7VTvAXzmrvdiKc+K2iDo770oVYPbClQkqZImD98xsw7UjXWmPAYshfxnw2o6bmNlEr
zBMD2EHymZRvxJ/9hsDtugsLvnY3LGl+3qd1paOAfkjngjWauOiFAgLL01m5s2kVl77ufulv0zsQ
Av/X73S6iCpa96KjkyyRIuQ5TszJtkawK3WuWVllXrr0SoUAw3JGnnj5i9dy/DOGpNQaJXXb/v4C
cuCww7mEvO+IUxijGKqQGaEUwvKmNQ9As9tvt4KLGEr7KCwRqqfU5hr2mHQFKPbuQZvT127d+WHr
uH4uEFVUNpe9jxwNiH5/4gRZI6WBQdSuCsRLEzorSaIQdCjtRTAaUrOEueKnlhNq0YJJTzXoleWd
s8x84Uel7vdjklWQCNTiWcFsU1FHs3dFWcDNkU0H17u6vojmwBHRcpS/QSnwa60l38Qa/Yjlc8qu
oJJst6OqxFSF2cqrQ6GU3BvChKsdiq5/SpZ+c0rNr8el2pbKPJuNf1HmCXsq5raAFzKvol7wzUb+
F8VLwGV9kw1Nv8ouibE4ZIlSCcpu/hCjCAwO3H+c675xXsXnGta1cBdXOkLuSDJnvYEountvgqU5
kWA20POvACbpFueLKj3lb2pKS8HtTsApY9Rr0fGjDphw0oNhE7sr9PycX4Yp4LhWDA7xw8kggU9A
4N6kCU2QudLKjSyku4CGpYQ6NCRcuVWfrJOjmeBkOAvxFQg/mLQuLqlcJRDmYZLLJ6umV+DA1zzn
mh/f3Z0Id1m+AKaTwHPwIUryG+QhA42Lh6mHzQfsZe/oj2GvTILRHEjQR6w37XqFQq8liOa99doO
VJgqOh4TJpzp22GQL2kyfF6vqqScMytsIF17T+/aHFtXdwNF4GsUi7+X/H7NTht6GOf8WYyAf3G8
JwzlFr9WuckCCJuOLZNVBzhD5cYBIVASi0kp7B/hedKr3EqnYLYGcteCO+n/AnVzVpRxd86aAiJn
GL4amNceZT3ulg8x+HQt73tGbQ3aYPe5w1wY5LrMAuWHdK9ybN04HlOEagLGrWqNpJwD2h06hZPq
T/vmq+3Hu/935AfKxOOQvhKgKwttH0OwnzC8nseGgom3tvIoIA5g1/TEthHeIB4tAx98bGbfEfpX
DftqFinwE8iW/mTxH9r0/SoPy2OPrLkxCT4E21OcbFJhFadeDWdU5eGydjQrbzweJmPTggtR5ank
La3NP+QbVQsOAidieii6W2+2inM7rdCrkZd9mfRDExfoqv0JcKwKRz3WTR9Q8usgvulVZ5RxeALJ
N02oSL2djoycqnrhO2T5yqM3/PlN9EVzbTgDMAYXlcgqZBrOOcUenWyB4eKzos6+IxYqRjWlUz2b
aHB0D8D9NglBg44qeqnl5iWFeXD2vya0JloBxoUMSjoxQG1Q/fzjliOwhSyrp1ueUV8xOh7ksReo
shUBN+dPSiuqbv/L0Mxdmnn1JDypfdNlUOc/6WTV4gYVoVW9aoRY0waEQaxlPUbYRpco7Hf17DUU
yHgncNriY6bHO/gL52x0+3l7DMw5oqSGivrwlx81KqYW+3kwDZGKJdsbiu9Ufgtj+G8BNXX8FZwl
v6Rvu38g+KrxpcC48WUtHnq8ETpNBW+sttVpUWTVlA3RupnsPxuNCSG4AJxdoyzN2zMhcqrGhQoW
WyVIwwCmayqfHnA6NoS4Z4lGjmOxFyMcZ9SovH66qAjM21MGfHFhzFBinX4U89JSbNyNor2u/HJl
GDMizoMt2DXrtc/6WOOeHyBHvk65XJY+4DPqCc/oJbd3k4unM8RRpqPnTobeHTx05vFXKZYbYHEw
SfqCcW4E3UbL/PPqmw4siksF6FSBlmc+I0RTFMAcrOmJ08TSvmVpUJ3i1I/Ic/i2/f9XTah6/lAD
mTeulFzPxWg33Y4Cj0j8OgbDGCsrbjA9qs3UJNblUfxHJWOaN9uaSShxxvnoFmpEVFR3cc3l1Snm
GoYqcVGDUQSrCB/EZ4BkjUjs21onPDXg1bKllpak/ACpHRmQNQOgZcATRIaQWljeJfTU7lmh/ai2
92PYqZXXklvE0PPzaJ6HTbjmRf1cpcPYb1sd54ilk+DMnXsq9h8iVQylxqxhVazVB6uzDIpaic9D
jxmT3DldSB/XZwoLDfXoyQv/rtoNntw1LlcKU7aQljNFJqfJENyW45vVFipPgXq1k4iNXwuhLYY8
/1VfHljk8fxB5VRUuqTN4pUlvS8jYg+X9o7OdngdLgZU038J/0288M3bDFlUuWCs1sqMIg83NY7g
YhfzXcIDGhyBYmbH34fMxFhmkqPC73hnvRLj2LPMCCkRvdLzkNPWExnMx7u2uAXb/lpGZq5RO6qj
hkN7IQkxCugFbObY9kOZt91bKiReCBWBpk2JSvDscM3IUrcMcCb2JFo1XSpSJlBrwgE0GwaAn1Bi
D1O33yhgBEoC92EDlPYALi3lEDN6jOtJhAPqj/A2nsivZQEzi/6zajBduI0D7bej2IcI7Bm2diBh
brWcJNjUCtZu4ksRiG7phyhvhXh81hS6W9xqsOjkXai9flNMHEZgXiDtv28Tn7KWXnYFxurH/Rlj
Uu9ybf8SHgoA743hq6cu1sJ+TDAI4WabyFNDbgOP04Mj7FqVjMmaK9WrwMvXludY4CiaJsoPmtW+
hm6tabs0/8txPZI3jVfNMX7gJ04yowqywBNDfYu31EyyYY6AcTc6rALLowP8hHiZd9Q3AKmOKSPD
fyXDrQvvB34KxMvgG9+X/ZZOR+67p/HrecUaufKO3bTbpa+kH7Q9zE0QjyOpGkbeaJgSPOGQ1A0H
eB5uTb4qZm59dts5SiT+cOYKcJFf2fScLiMWKzvCnlYuvUVf/steEeK0bHm4eT5ubuJjnX64eUWh
r8MQGOijj2Kz+yXnzPOsPEmCueM6ozAntM0b4v5U/pZQj5Jz0Y86kqH+j1pD6TBX6mbOtDVAgGdw
DdhkzZ9APXJ56ej91NyELXVaHiITi0dKvL1iKBCa4CsH7J6AWfaW47X+v42kKKvazQ1Hw8xo49H4
6Bdq/i/9mkLUCl0ZCfqx8Ii0FHTmL0BvDUUreG5DvPqkD5z5nsB0H/eKHIaI9XT/amPZUZ30+u+x
1fg8nNeI5GKYlDmOr/NNu8vUyJAGCEkGYI0cBK+UOGWA16o4g9k6Ue3T4ghpLYclPtnHBMo3s2eP
yVAzaI6CxP19X3nRINP1hrT5KBv4Wd7Q4Z/ZhDtIzGdA+RXst+G6MV6C/YhSc2J9LpgBOPGnCy5B
jSnaiQzv8wRpr7MMTdRgPUnLTkAeSBHKoYGMXWC3f6IwpojSGDqFp8tMSv/WMysj7NqCiVYXFRLB
91i6uBHsxy2pbanWmN4I9pTQRHLQ2ERqqGorHcSy9+NfLbOUz/fpxQMs4f5K4wX6j3kAY2pxttOM
IeYV/pm8t52YK0I6a4d7lgC8t4yxvwNGqF400JH0ebXgi3ir3wNhKyxaUPluhnILQK7JTTDmlrYi
vS8XjjJsQl/8zVeJdvUfdAB/O1D43Uld4Z6HbppYpddOaEBgrELKtVLf5VoSLY9Qtrr9uC5y6WH3
ZY5Lh0vxRXYIWipDYKC/WS9B8Ew942gTSMRtCP3LMJ7p50n1DGuR2f8wi0N7cbhIdpDHfneLseG/
FiT1aG5fOBB9msBIIL6bCxpqRpYaInSFJwKV0JBlCgdwKWoz3hHcuzzyMDU536kzQ4Odiqv2OibR
gPBFAIvWy+pctuIK9KUxaiAnY681maiHbaNpw0ZNySMig7OrvVqdMLQ2olTQAYHCITAf8twzppZM
ni/FpCAMdzFtmqGNfpHaLewrr9RuzAhQA1uchm6epsnKlcTWYPxVLYd6qdYYrFBIzI3hI67mAgtj
jfU4vDWmcyEltqYDIL6t0W5iRvQqzP/pLt8bu2DbTKI0ZbpbYDqGewn7S22+Fhtt/5TCTCe/pNmV
D2Eoo3A9rk59eL3biH9956EOJsa8VLddqjjOpXJnCXi/246WbDzpHdCFDgpDiu0tYEaA3jRWNFV/
xR2X12jusz6FZt27mbnpUh0DMaiCe4RHVs+PO1qZosrm/0PeRUHSnBZtrccXAU0/94vuqLKZVeb6
ERoF6zg51a4Ox9CnYCxmq4p+TA1warv3P222EpD32S8z9WWX45HnI/blxDDG+kAvlliT7SuWtYt3
y73LlE2jxrl6mzHx2mr6GmNoDnunl9d0iWqxyIPZ/oRc2fa4nJy7/4tEPFFWj3GhmGODcFkflIxG
+aOx3rt+rvdlzEQ00JrjOvg7sf75WWTfCKTKURZrb9Nf4mj9SvMmsqozML8AhLGscPnzaWajjCB3
W1PhgoQSHhYC/sCd0txRQoJZoBUSjOdhEQVWBxGowEjEeNyS4Vq2MoL3M6J6JKfVPqUnYOwsijUN
LOdIfUx+kkjG9tJ3uNzoBUOeM/0Kasf/54r1/mptrDWq9p3pJhk5Tk3PwyFMOPuiF1XG+Jqa3kkM
PeSZXv1x5DfsUir6jXOFFlIxt5tdnrxosyecdFpWTgGoFZDepn6IKjJmheO54Fdq4BVhrptOZ8LR
a/5xnKVJpfHVWDFQLeD8TueI9yl2xah7fD0or9zDnGe91nvITjU/tiJwvJi1iC4WrXltDxzjBIqd
ACunpa7Vpr2aAw/tnL2Hfx9tYM3PM6HvWmt8rTbwf/icXeJ01iGxacefYdZRddDtXUD6+Z4zWZFV
t4Sc6p2Hf60I7fo50MT3xzF395fqMRGkGnHGMZMr4PAWycEul+iasoycketCMa6m00ezfmTTDRyg
ug5/G3e+v6QFvvtcwY7f47DYc2sqiZqHAMZpDKmtw4Ok4HqZzXWme9TQpwHKpHnJx/FtBak0+lJy
qATST4dZ7inJ80DmYyJP8UwC112QByAHlK80UITmPMUAeIv0oTxl4NE/t5WuXXhZtsJB2AmMBZho
Ss9aEb/CN2j/rdXorWCz+smm7Sn7EHZ6L5XMP/gcJK4JYyXufMxo+59KUJQnrs2GzWgeetN42s3D
2Vgg/tQVZR2qEj0bTLO4MlnGur873Le1LEHCB6s2gqkPQ4uSP3JYLALKexHFvJt/5JKfpNhs/noH
ouP+xgRJJ2NM37zD6+1aR/WpRMlewV01fnns4pTDLHDI6tUpwRumwsLPSx7lzJp7Pg0j6WKuqLgA
tROHd5V5pzT6rPdcc3NIdpXVRK6P/1FKPmubUZHxHuacK+FXm5Eb/hXdaZO/eO41c2E3/hPpEkcE
eT5NWm6ycfbC6dXXWAtYOB/CWxrwn9mZ9+PETlOqqQ6HMV4Oqvmj1ScrYtArLH27fG9CSWxHsunL
cRxCud1xFGd1PKaCoIcdE5qa2JlSki5OBBHv1GyFNeHvJIGoJ1jiwDipFQ2DZvBDRK49lPeVNAHe
148PCautMVQRJkQgbcxz+jbv8LfacMs04PpNWOO38oywutFnQrdeaSPhNE7Chyv4K8QXHNwiWp7Y
6dNB0wAJTyjTPnmmxZN1Wztd2iy3i9I4rFw7AFaTK0SdmUgIRDMnnG5XgyYHrujhxmR6we4IKn6J
xnBm1k/RKU+UiX9Mp1eRFoYKo1Y8Sa92qCDjmvAy5QJdwgo7+/rNTiGMBGIvHMuGcYKBNC4pLo+6
FI6KRZUH6BVPYH/eVW1S1VoSNpilo+F+p3aeEJFhwOCnceGvuxVRKAHDEswcL0sfYi0Oo/+Vo/d2
SpGx8XJLQa3xm93nQgfuBZu6WpfpDFeZFJ2IohIsEHaTXUTSyzX7yCyNV3jOBIopQdGaCZLILXSj
gyH8X4JcZ8T5D8pH9c8fgCPpMYMWzb9ctDFdVVCmTXZ/QsjwOJ/Hw1DQCT0McidAvuUt2SKunDmm
r2ZluSLNLCi8Gti+Tq0Sx4zicnPNkUrlcsvPGBJO33xuRuGju7RJcoiDhr7uyV6zqYgez4BFNnJC
xj/zunMLg9j92M3Tsq6q7XtvNNIR9B2mt3tuauLy/AIVpvB1mKaYDEbkzNVSbPJQWIKKeUV8TX5e
jfgRQyMLUsDJEQshWZI0e21uDr4WOv7AnzletF4olSE+FvzOTUTG6NP8Osy5d8mgJJvFrWga9eQz
6TNaEDwC/Vxt1e0k4ZK5zH1mjqVo/I5kccsUIjRkkojfhB1SkAyoC6+DD9aGMykKR53Sxh/4UT8X
bAKWNCT6SezFiPxeeyref5G8VOt6cvrCnE5jGGjyW/HuWT4CESNxrxMBd/rvsnjqectIjpPA8r04
A7LuZGr/i87jQMkN4xrkdpnFKw7jl7LAWpF+9eh6sfyYRpMWEcrb/+S+yTSMQmOtEQqDl66skIle
pgjTpb+Ks1sjEpYgcGEY1RdejUzWyRq4PM8Yesmp4DaWKdz4KTT7059qti89nhC+To4czHRGP/Xg
5judkn5yD4nj0bd0j4hN8KRJXGxqFyenbHdiurEtbnvs0oUmcYTAI0fanPwzZLGLyEQsIDtsI5FN
M6phR/r+XolYYSGXUUTTHnbc/Uq16qkiAiErh399moo3k28rg4WTXv4zUjdqrM8TiSOoHFcMWCfY
MJof3h5ZlhDiabi6UA6sW6fZJOMeAUzJUVKbDIW+ZPTD8Ya/jHtNaPOuDYlNQRsLWmunj5f/mzhY
eGe1Xwhtkuu9ID3YDQvXKB3qPw8U5YOO3vfmYmLvPGYMOL2x3oJ9/U7Cg8pmb6OXA1T/C5Hgyyfo
E4P11NA/VT7BxNxR7lBbeYgAByighQ/r4t0BsAST8dIrdGvuXR8IjCw97ysQ4J7QJPkzGeFwFxVp
8VIE1HZ8j5DM7/5mI+hRGIQ741hO+yxnCswsk0cNnt0VSsNq4mjv2ArreNaL0HoHjKLV1Bs4+Z8T
Oz6a3BmJgiEUR4jMZhwP82l26Q6+fK09O/1YiCSTCamVMjTXjBox97F6s9l3XI69nGpQzTuvRRSe
zVKklBIKDouByeZWCvf8FoyAT7HAaBDTLTOZgSo/Wzuko/aYEcoqd65jxIo5hf5+Gq/8qm5cI39i
RwB2Rh7w5uqD0/wlhSNZorDw60XsmSP17PkPljh1c248dTNlUPEZYMTxK5EpuJC+iyPR9/vlab7K
S4mr4fOfjQRSy0fUJw8MwaswQl8tcJbYnUBJEH6u+Mph6nvCg2kmFjz1HAOm+sallxSu/xrwIkOv
Keqx6hrmY1kl00mlnsnu+65FTJ8MU6P0U/eWuhlK7bfNMp72ZFvBorcTKXfKT9UsTIIPbRizE3As
OsrvHn/GGTXQsg0k9pMVbnNmQcPgnvmGYOqbTIF1+1YgB7BPechjVU2gegPnbKiQ6/uOwwCsBE80
XCn05Hxp2SjwhvGv2H03qgS/C3WIoJEJbZ5MBvSmYCEPRgYH8Ep9hIZC94xcO7Z5O/TMA/HYbrVm
4XzQA+lW1xkNoMMUTENUxkhPkzdLwI1Afy0d+pSrPTZNNm3ldbqYURR20krbPKmD9mR7wPqmu5KU
g/5nqTMhukF+mAUQa5u2zDKxnLYXKy1rMLbUjJ3XHalNjP7AE623VKQFeYv2OIi+KCwmlnI61zoq
MilivFxeZ0sqqRMlYw91rGoq2TfqrQaZCcj2hhDcvVnwS4TCBr1Vh+abPRBhjEDdQVd2gloBOiPG
tC43Gkn4WvRoYYJvEghntuPPM3/V5NAEknxTcJZPnUusEvwsXHX3v/hlR2lhwguNBRbDEHyxMMLY
XGw7qfHYuu6vonm+mazWf0YsqNgqZxgOq09hCXeNKcGeRyn5QSRw04n4giFwVSRt51jtgOoiDFDD
cn7aN0PzHqqoyaROKHCM93GAW1Mmo4lYsljK+lPX98EZsre3mvhYs/GF67l8JrKp50JzAhyhchul
e0WcnE6Z074WmdfjLwx4vNmYpihKWPr5aXS48x2bK3bozwyx8BfyFs9VjQ6RXbUyeChZFPC7tU7f
0drtUvZpJEoP0YNv4INMzabu50cflEy23c3S0qeEK8+PI9bSdNxB+yFVDAOZFJT0bkyhmcHIHkfH
tvGmLh3L5fSFCKXeh429xsP0VN4/j1uetVjDLNXLkLNjvhgmjvaDnx1J5t4iLsv9J8hDbxOz41+i
PrKVcFCDpjepnEng3fzBBCGPe5gw4/a8fVdR7myrJKg5mP85plp1i0VsH/5EzapWmHZ4LB8hKYbP
YFYs7oweBx8ol85a1dxEzWx1aulS83BIGFdDpruFoXEmV0YvndNlY2tHkb2RgdTjyySx/ckCRLhC
QrL8fevxlTkgG648ifxVAcNVWdKWek3jHFEIEVy/kPHJfGU956LMrXgWNVUuyla6EPGvnCiw0oil
BsmONykmWRBAoqUPonDBQm0VtRNe2mqOFXlUZA4c2szUoqJGYJFaNGSPIqRNHXq2s6/0YkREun4u
Dqct2+y7Ri0yjiZQID5AKcQ+C6WW+wI0g903q71/zNKpVi6miQMzjp9OF4iFdcol0gGlV/xIc3RH
RmhOmyxgZ//vog3sewY34HBku4SUjNK4XQyRrCXA5NE73QY4f3Qa5Bh7LGboaqq18XYQTWO/QgzU
RZRgaeUFWGjzrRiGvKFNYTyekWtcM0zP6+g+qCvUIDPEzP/w+phm4dSi7tbbdfDRNoQ385kcpPCu
M6eVUlK0Bw8RJCK+vMK/qSOra/Lh5iTEXmG+ZYMuxLNQmzHcUlDMzCqWCLZJNdiBjaTZw/0P348R
KGS3oedVFs6PHD8j8xpherUK/YblFyw9VaubqepfKpLMhVI/bRJkqmiwVegYqBwjq1oM2wMy0l2g
r5wjTVwSnAnAeZXLzljkewVINF39gRx9Ye9Y37Rl1rRc92kYbWXvdA1eXhPaiuGPSr6IJzY5rzhE
VU49TzVU/ncVKLI/hngaeJfUIbJ5lOeoa2muX6+uYyDyNLiL8kmjCFXUHivOrB8hkSH7Ic9s0G5N
WWDeooQJ0ni3xGHFupjLbob2cH5qiRSCKCY8WBKTIBst2Aa4mVvSTQu67Z2rB+feSi+tPZQ0q4y+
lSlLJoa0y15RyG4I/UxswyOwr38yOJYSPCpigL8QWp6qhomh9fb1XlN0p4NsUSx2Hidl0ij+YNFM
hit8KiTXchilGNdxARXTOGemGBlm0e9uwicpnL0SYhFHGGu18dOAkHQhkWeAT7ltizZvmvO7cGm+
egc/KaAYPFYFKq1cQTUu2IYmsbUQTJMf/IYYWwpdDxpB45Gg2B/Uvsgoz0ylWJ0DpDecSbb+i6cU
oZFvtkR4AjNZSO3tGXdm62KZyWF3/d0OIwOkm9UEEknCA+izmbWhJqD4/hl0oZPGg3KIzRyvQH7Q
lhgZccHGv3n4+ZJbhmlcYKnrZDiXoUYIL4fph989TnV2gG2zqQcrCJMdNK3BHM7w5rdhe5TXrK/o
PcBuSPUkloHDU9YQ2DAuVLGGYW0XlrooidNcQglKNKBqGO3caaZM5OLt/KpMYZEgA5L74BNG5cSt
CEoItslK8chLNfdJ1OeYvcYuvISK4kBw2zB15sVIbaHNOl1GwhZoskT6t7ePjdiXECwa/fNPQwJK
Jyii1QEj+zQ42rrZhly6kL/HowO4OHZjX+wQDRslocsx+RkUfDLZ0ViDxAVonVj9NTOXiKHDseUh
hUpq22yPFEDWnOLIO6/VqKrmoP4QVjjXiz+7/Ipf5BINlh4xh8Df6Tg0vj0JEt3jNcNyTIIApL4Y
aR2qIIR2f8WeRf4+UUDscn4NbBapIfj7Ln/Peyc3oSDGf6z7xfsWI0V8SWohFdV8CTKG0ZWf05zB
f5LqVxJqASxVcMQeRMR7ZYXatbvg678AH8gaXfgOV58TrO9yGD0c9NR9trPm1e8onUmON0xnOn6B
TqrCiAEnT8qt2XUMbz7XnXoo4m83V09zvOac7CnoORUcyLg81qEh6BrqEo7FmOmeIUDSs122jEtj
ualvCf4tZO/ENKhmfwwxppOVCx8ZFAZaBLRe3K26mPw2DOBbQ4faoT11Ydw7lCdFD0lQ/QHzJdSz
GJqATIwdBpv+cvkVYJmid108BkUtoOJATugFVMfigbByF7MWu3sMobn9W4lDMfGY7SWDtPynXib7
DbZqEm9yzEAZ+RtW/vikpPvM8URjfxW7et4sBJwZk90ihZiNekrtdsQYfcKzDRgRSmABvecRmrEB
pOf9sOR3CR7cCPS12vXSZ9NlpTA33fzdtp25NRwkoDiOBR8R0XK0qnFZec7Jjo8GtN7x1yfcKOCJ
kf3cMj5Zhub3x9z6o/+lLI6vEImpbZR7cpN+AqRNYLZycZcLcYwuiWRm9zkRyA+5mEiyQVd8pYJt
Qyf9i5f05n18uMqd0aokSv/fJM+7M4/4fv01A2kNpGX3/PlpgkdXqrn1traApXE69/ZaeBN/jbYY
jfYGfGgiCfH02eWwmBuWX3VKvXO9EXStLK5S43mMItwG9RfilrOEJ1yzQwe/YsS5LyieMnhZvj3v
tT1NU/rN07VHqJdGAfsZzyotVF2ma6YVJtpQQ2q/ATlxfzYIV+LvS0Ka/P8zGjLuJe//EedgGZbC
h5bu4tvwMrMHmBFW33AzMk5oWF8lHGXF1pumqtXfh5NY3eHIbxofXB3YkCYFeWtUB/j5ZkOhMk4v
G1wmujdfatCR0Zk5/puVS/iGjLvh6eqSirvwVEWLV0V/kiGUM1JAwrCxWhyclEBvGM02OQ472Pn7
YvlWnnNjXFoaF9WJlLKnekVxIvXXm0QqOVlj2FUvj35512kQTUUmPaTOLsWjx5hPY7f+WZASTs23
8vR4EJ7vCXrv+jQ8xb/Y64ldKKE8rItNhNZFtBVmPn8nRR8t4K9fLEPuvDqwLMLkmA3tDiIY7VhL
ZIj2pNfWp10kDyU7jh/yaJkn7MzjfPFFb/UHjns4eozeyuELDOwGi8gYYJooVzW6KWbR2VmMwMyz
H1oAYdmltkL5vOTLKASYZsac08dpXi/MYO7fnzNQPl7nZNdjowh1wBN4XGtm52d4nRiRqyKuSWO9
GYu0ViZnaEZg8KmkoHv1k0pIPVYbuLiip5VrwPd+Uiv2L1nK7lwn29K7ISF4tCrve5d2xNsxl3c+
6SU067obgK9KKKIiuWQhp7bcSGYABfE0F/kxcePpI4qLIgeTTVr7Am75TuGVMs6XNptgSt5s4m3v
Ijwa4KylaM1G93K2WWoj2vWEwtQXS+0mIwFYeKq9DpCLFPofxs+xaiAreLx3wnzSlhn6Z3WIaHew
sWGWTCYfoxyC0brOUb+yO/ILqr2UxgH4Qmd0TldJWAWxZ1JdEF3E0acgR1i3VLleFY+hCxwPdy8b
g68tPCiTs0Gm7Bhhk22vaDRnLXEM1RQX5RBiKT7sGTNxQbCZFi0Gl7DmFcK4vMdl86k0+h6Qnp15
ZbWF5L0IxUqkalLREpq6QB7sbxhUsYlih3xGFkiHWNLkHDC2A3kHcJnbXxgNwS53a/G2ktjSKOdm
g1oyBvUgMn1DMXe2wVkCkYkMYDthWBOXa8+ZJJ1zYvCS83+puzA+z8n1ipEth+BbpmKNRI/lh8/N
R3tazFX/hLLycBdm4S7oQ3dl/F3f3yZFGTKzLMhjMtW1xLTCDw6oHObCXV0YjxyXtwJdDmmh98Ws
un4O5K2Hlnr3JVzRDnFoB9PIOrCgNeGxvJUwnAY0Yc7YXa6CQHE7L2E0h4Skrtl6LR0dYBeCVGg+
rNHAweH9+8D1xZRWQthkfQ27BibCng3v83Q4LnS5pPl6LdPpHhZPDXwYfkkEthDo0KHVOuSU+ZKl
r7ry6yUkxW+EeHbxWgC+/OF5Cg8ICRP9HWzbpjsvCa+QUcfiop9jIHKpTaJhTJXVBpmNuHWQPiTc
0sRdHl1gsqa4TGFhCg07POQCSlwGEcQtHZV527CJrxoubna8eeD2zqAPWNZAm3RBz+xPD7WuGsu2
QOMzKkPr4MVG6Y04ozcfislLRVlIzER/vn3yoftmu66tsoHf2dRVTQ5csYiv3psGt9TV9II+ZKQp
C4gi/DbWa2TEvajhVD3Z6D51fSCch5HEb0ucOJFXp3f3KVSJIC82BRx8GPa8F2GpByikLSe4sD1K
ZBt4EGygqZ5/uof2B6R+Clttljmty07R8he9n1fJVk67Oe7o9EPLSxuHih12Pu3aXWLPsy4i6T2a
+aDNI9SqQMGY50/Pifaf1Gw8mVHr/Ry+YNYlCUCFbOqtrJwK64QFRcu3XH7Tx8iHOApCEeTOPfQk
pILQWXmJmbWZWiwqNe0Dw7tbO4MFetJls6WEGhBOITOrd57FMighSu1E4NAa0cHeIIlOI0V+pGE9
nYVFD4MzAw0g5zt/v4z7eQxF3mi5JRiuBcIgVbO3H996zvIT5oh5NsxcugvFXSwOwj/G4LKqSUGp
fzh+vhX45sSLsYw1Nf+epoK0pvlqAaaQCPapwT8DsS4rSA/0A8lV9s13Sm3rMPRs7BYTR/xHDsdO
WnIsSVnJo/euhGG9FsNO/hQhcrsl+mtDFNDmuZC1nRdEBjVVa9jp0Hgg31cwtHh7UDmBLaQXflrM
KteUDbUDcxzgmbcPis5u3KyC7fUGz8lUIdGN/sSbOXf+H6768YdKgQ0taPaiibELmZXtCKNg/Dsd
wqJrdYQFpWs1qaFURC+s1lFYdDcO5iCPxbnRLNV9fakW5OHUMgiQ2o4WBKx1cBlGDCWZyfizqAau
uD9Kap0BquoSCr1x/r8A8wQMRl9pk/Iw0GpRgVTSmboto/E7Suycg/i+bl2MnBanNE7vDIzAIgbp
v3hXIuChgdqaeuW9qCKo9qP6uqB1gXTGZTJVBk1NFhDZubUPuggUGcR1bJk0VktjPc8hPw/5HfNz
9JwaJ8AD9NTv35QVYyLmYyZqOMiWEfA3IajPFiK5zVHKdsI/3iPH3NLafbtRRpxHkTNCwtBH3d0Z
vbGXGO5Y1t1abTPRDl97ryWVsuMKT8NaPZQxyo4T1jBJP/lNpdODO0vQ0VcObQJkyhXvxQ/AYdv4
0CbvzTDyajoHjT+yyasVndI7JF2lFSnNszhzOLA8vVf6jFMbFKp2ymTe2QkLUaNXZOMd95jzvD30
Ni3p3FQQkKN6eLRehdQw2XV0BAbcHjoe0lSAvGXayxmrL7yKtcqtJo3weUYuVjZNbmw8ZjlgDHma
wHOS38Tb3L07bQLTh0eIg2gF99YbABDTLBdSb2BTKecxaYss+38BBRFTq0s+5OAZJDJyLEuqW02G
eP8P/sP/Yp+F3Mhl++DHZnjYL4jJfsQjtftgbt3s3VjbKOtlx4qA8gFWtBAmcckH7sR8uvMa/Nto
YexdVzeT+oANw1Hxi8zKAYHsZ15py4x4ypjfHsf7uwwPvPYOeJDkAHHUL1gY7WiBPjkToCz3djSv
yyUba7LZx51rQPksaHGyD6yZrqPAatWEpw+D9wLIijWfABidrgr05WgnmS9ulOtL5SVZ6z1173wr
uscWeAryA7TerZ+GqXRLhJU7pLo1mufNfGsouoJ+8SFzHmcFn508CTfgHxtBADaFO+ubd6wIvLPF
jUgO5JnQi/48ykr+4uGbhszC0et3pl4ZsSX9uG80FBM5LUkewi2JscuzgYCVYLRIICZ0I9k5nN86
AT957B4Ug0erw7qvVlmmi3xZepfN/nlACu/KfU8p7ZjyBSG4iKcHozUUKncpL437/isDiP8sbLgh
cAYrL+/UW0DUiM8ad3mtruIONMABOJ3nEZazcaTVnoHNxMkxOhiXJ/JEfsnBsSCt3sRtXTi1KOiM
FAvp3zdezMMaW9CRq1Qf99OceB40Fru2cQcW70kCd/vZlx55S66yIVcEusy79oujcOw3p5uWuGhh
C7NKwQNyYbGmMd5KS9LrlPWboygXdhYJO86un1QOHWILeH6q+sMRDoE/+IVndlgV6NvlAiG1dIa+
J4z/e7rFC0TcUKkEXkdpdW5D0DNGLx0LchoU4P/Pi8QDk6ruw4G4t+nUxVOaW0ULgcRTcYdPcBEC
bZZYO3PnbbN+1V9+etvAgAV1+3k5HC3l6D8zOsbkifjd8fpPO5aVjjyoiUtjRHJpb9KLTuSjlAtf
e2xVfVg4ZeCGqWbgKdXTVVAwzXLSuTBBIkzu0dsAH2ckLF0w29fSbZTQSqsPH/OvyiBM1od4MyrC
BeMAZ6R6eGukEDh98epoHmTt7rOhKHYopB4WnDHthJW628ETpC/d24i936+T0FdoVkvIJNKdnt2d
CJX0OdvGYs7bXHSGDNfdSWy3qYtRP2hezabXUoGQExo74+HLtW3Ep02JtsYsi1Oo1mXpX5HelpOv
dTEe56tGa4bnuTaIglD7+VsxGOP9GAN3sxcdSosg/Web7/XwcroSTww2emCjKRa0MFIuYvCo7vmj
K21oEfIY+SfrWi6EgKJkJJnEr8OKzYFwe4H657tRgR2ow9OtcRpudFOJzSZ+bASz3hOhsUBcHM1g
kPMm/BhluL8WAWN0zGyqaDHDO/G12eJuQB8bqLFGN+jXJMuWzL0NI82hTSv7AlTRI5bt/Drn0gXA
hlqF/SUHHl2JrcxhWZI+13P3F/WLN6+LCHHtxBUXnk/Ghk6liSakrIioT+8OVdFdm2bWVhXFIuYW
IonY1CDlNm7aENSzu0QlyNgFUUF5hMtNcMKH3yNIgfKDxWuPAeJdOp7z5z+mhsRJFbrkoISOuZGG
jJFK472ysm4G+E5TYKiFQm8HpWj1I7QMct6NDDLe8hWnGCzrGDK9p32J7YCnyJoi7S+RXwHJeNKO
mroi9QxOisaZ8jwPr0ftsCGpGzwsaEzeJ3xctq5roNFK3ZtnMa5tAWFtZNaGjArzxdrewvaMgfJ1
sl6i2Kvpu6klFob70CDa9Q8zW9GX5HHx5XQT1VGo+hvhT03Bw0Ht859xt/XfGXeoLs4wVQoGbTH9
U3veEq5tAL5nDSYn0StesZrUoMvihOHTuvCLFjmf1D7J4G83aQLDdgKdS1+dxP+ZVLDjwMt4zu3w
fTQ7pB6a+hvt3Nd7fW+3rRD03PF4jCn1l0pdBZNjHXgEPIyLDjryuBAD3zfeW0utGaWd7DQ8duuw
ln+0/Q/awv4/+I3IPqibbzaaRUU6mQ/zroP37qA2uVsb8Fof3h5FK1dM7POKSUdL0/3jOYHqLaZx
v7tvGYZBsGuXxROlKxGVqAqd4dYuGs+Nx7PP8SniUyDFvYL0YJt+1yRYgxNxvTt1wq+704krac6A
fsv/TITkxnbN/VFUp4mlLQc3Tmkn6EUCp1SGguHDvxlp23U8e3GsB3BdT818B74mL9efNA4R4o6K
RKxV0cOh2tnx9vfSN4hGwt1pLSWrx96nBbYHxu08UfQhhvKjqcSj2tbWZKalOXrmEWNfSrzKvb0s
QfvYE1Zhk1qzcnUbngjd+/0RHrSxMdrQiSgmbzJKSuvKzp7x3ALYaDXK176XqumhGnM55ERdsbEM
89CCKx7fb/2FA5/S34WmyMhTQfln4CN/+3T/zHMTUmbCOqp1GniYn6LjnRC+ass4Dyb7ztUPhXNn
gTY98G83dsWD1HzTNWl2RTgbv5IoTFh3qKdfeufJUuaz9j23+ISWE7WqJZBus7h+auRP7LOw8JeT
MZHpYJOfneiQa5Ss+QVaKmulG+02CsyBexKsaKEByGiz6sy8giQITOg6jZldU5dhdaK9ciBYneBQ
5SH7uC2DAOt/ufBDqe0KKxb30E8yvSEQgKoAWnxB1EWlzaLD4vQXq3e9WbtuQhMah90IT4Nb1mJx
V2gRUFunbW5q9CCqUHmS7oYuJMpTjbht6fscea8oRI1pe5HZkj8ye315dJi9qTdti37iZVYq/WWr
ijsoHjIRzqAIxZcrJqc1Ezd1e25z3PzsBsTO/kJVKUbgKO3ps4W/SU3Bz0lfVXl7zt+TaEBojSgE
o2dm/YOKf9I18uZ0t694oZp8aZSrbVNcos6sg3jjd6qFrFaMZb1X0ABy7fHn3ghW/3mwqO0qI04M
MFJoCDHG50qp73XeBMv9jXYUMpY8/LOajn08DxSsjrQ3Wu4xnjF7MLrCYS+bZdTI8uUZVr6zdoEX
UKD4cJCGKbe8wjv0g4dGCUy8KLtK/20z7P+sgLUf/iR97gFCz1YOK3jUKMwvA7SEsmklZ0ckwJ6J
Y1bCoBKQ36tKfBfLsQejxrtoeivI5a5BMbOeIAnBq3aooUDo4mei2ctE+DAv3kbJ+PMZsR2DMzlU
1jqDX+LhmjK3Cc2DLRq90xUzVg0fC+mdDW4o7mQiPXMP2Ub4qEDA20McOUK4SM6jGLf0IQEjtf79
BTVD+JC0X+Hv8gMvCUqPZok2x4FBrz8VzuUrKvR/KuNtfyzPCHqajUQiYuuOiSLCvSgVnov4GFuT
OeGupGOeFmwZznsp70/5Gk3zaOh2QAtZ9rk5ZfcfX8UVmEavfSOXoMoxXjY+V70pUl5RdqxCuxYU
7Y3o6VmMxqIoz0nMQKRbTcKTMstfBgsZDveWqhRmGdCEiD50X1p6czHzV17TYu0+seaJX7wSiSY3
gwECwFaIb4buEU8HYsur6sRoJZnzvZcAwaFo8m4nWO2tZzzEy7mPqnN9dAYCPaTqTENGi1o/zeSq
dEbVVS5TvGVspztfNY5baZ2NJeeztC+xVZqWHTxM4l28bNnICzFVmMPgorbsE8Tm52k3wGzo7SqT
DNwlFNqmemFi7RbYhqW7+PjOvQRZCFvKuyoEyQjJwzkTVsgxRXE3VEAEPV8tPpFe9joPHaxmo6df
QwEhV3rgLxwWv754L+dg83KtnNphO8SNsHF97u+xTacPJU4fnu2EKIXqP+afrvqfQ649lmaQ0voo
o7+0lufAiibOAYSVUbarhWuClHaCmystpOtcky6uLdrMpTZejIcskSyU7iadkzFRM2ezYH0cjOhc
ziWyr79qegTz1GQz/wkH6/s5apjibySUmB5G16do+GNVv+vYFVOLGBvwvXkxD1vS02vVk53Kgx3U
KqOOKqPdPsUP+qFz2Uhz7AB06ui9LPudkvpn77zeZIDD9aAe/Z0ubMX03KdjTi5sxDKb+qyX+JgL
sjKTRp26iz6HeKC5aKzez2vGcUry3/jYaEBcz//UBHm89XfB7FCbKGeYCtf8tiDVOHP01Ti5r726
39ijlTvCIpoiqizFCsdA1Zr023cmlDj4DrjTcfebiFpt9qHCw4FWYy+sk1tMhc87JO1wh+Nue++U
q8RVBhJnEvHBsYn/hOv6lFdACNvfyFPQCDP1PNwFL6E7OM7uWfNZ1XbOPUFA6f/LXuOM2J/pofb2
VNtNsFz/asj/v93mhTaxjxRpLQvlvbiWx8QQMhImG/3tDUjc6MaR34vVdWZjOTMr629vvf/UY7QM
kopVP1mzzQ8ZNrIQlaNs7WimUIotI6xj4+yLGMUsAb7M4toNyvJFxTB68x5Ws4MdcCfBjJ4oE5ji
M4bi3/FjDJBHSfLnUDvaHaAyCL9ewuC/yDrLy4SOUM9YhSfHfI8ScXlPxmBKEDqLE/jkOuhPQiPt
tOdjHhW0xe2OYxv2osHJfd3cuzj+xhYLefM1CDfRdUvjoVhBfiLU/hKzb1Y4ieZiMQuAJG2xbE6T
tlXSDpqKgxNB6aPprl/5mC4t+nRPYv3JacxOnSGnT282fq0fYPfNg2FckJLZOIq1uVumLJaPW+uq
PBm9vH5yxQ3Pa1Q304C+0qqlsxcm7hubGWbEvAaK+Gr0iocdEw94pynC9lVFhhR2U557WdtMqAED
vIzdQmHddaeyWVnJq17B7oxtaFUeC37BMem1SLsH0MK71l9tFc9BQt20VEan6a3sKVRL5edRGhTT
pTU+CyIoyoj8vXzD15Y0UtG83jNuj98UNPxlihJigRd1hW3TGQZIwU20y+CDRfqCL4GB0UBzNV5r
BnVlNZAttBjkZEU46WIvcCD9cbuF7MOtIL3qhU1vkCe6KbY1kizGX7OGAGojPL0WODWSjJMY+OjH
+xBsDgZ2h9Vi+nisZ08rsbPOr2PD2vG08sQ7S3umfJLeKV4KpfYo+q1mOpRNseOiXKr0CZR/ZclE
z2ffoIV0znaoLI4wY4ft5bbo8YO8RT3XpLB8MERBEZOVuRqB5FmeA5Ovz81+hSS+8Wu2lRtnPzHD
zusQD8dzi5TLjOGAysnc6fDcCsN2k1qnxdlcYoE5wFTck/lCoWe2ATzwxoDPZxsGYqd3L3QXrJGz
NUchEP9mtgRxaSR42J0GUfVD5UwB9nL9r9/jMoalPadFgChKVNT+il4Wpi4KvVYxcEuppWaBFFis
g6Z75VdoCgblKOta11yRoW0idATKgyVhPXpOItPqp1iO+E1UDQ7kgmu7iyY7Ve2U6Eu67W6RULrv
aTtWzRFDH8IU8rRdTzgT7OMPnW6mxIvArckZ5mSmoc99Yjf2ic0mNKW0bGga1RkQysoWHU1VuOjI
lEqAQ0XrGDeuAKvtAi8fWrzuTd8NWPnR07Ku3WaAf0wDfa6LrRlDMFHIvVvSCCVr7xixvcN4ofyH
wR/dH9AubFD0YNDU+LhKVMwXXO9zVlTBVamTJ7aOXk41P1duw/b3/yXISlq6qW2ZE7P8amKbQJrp
r3Xz3fi6zQ8eSkXdCX6+KAcTpv74VgDHtMhM4qHw5Ws+R4SwRCVOtBHdbMg7vb8gNG3rDaP8mpXP
Hh3zmUGY/Of40mhqRux6N4FQLTHgGSiSdns00PogDclE4Yyz9TljH/NeeF2zzeXnbwpMwrlJCxei
aFYeJzlcKAnyzSikA6rXGfeTSiQLZaUI3M6M0AE7wJGeh+cHTAPUaLLA6f72JRO7QoxZXqBKy/15
PqaRvKOUwkD7AkuO7IhhD3oYI6J1kHyjISvK78l6IbzVRBHBx9UH2UmGHRQbMVamvaBpPqtOeT0M
HoqB3o+4c3ZngM7SVENX7duIX0Gozt7IQL01tCk+abJIWiAIx0LEbmjaYBkc6F2RTtDcJg1SEsxf
UbUujMTAF2/cpSxmVPuXAShasUbnM/zNmf3k5rcbqJjGdysOWq5hm/1dFy0k/OpdtkKyaLVNLeXj
Wb826ydq+XVXfSItiAd2ANuX+WRGAb9E1Vg9ofpVf1/rMhdsPcqH3lBvR0s7XfvsaU8aDnnrWi/k
Bu0pwl/+mUTyxhFhmRQz+IHhDcIXAY/gTnWgwxasPxT/EepdkV9ducEDH19r7NpEABg1bjG7IOHY
q305csVahnDN8KTjF2/jIzfJaMyaw6X1iww1GQujik9Djq3VYwiqrESsQU6PxInX3nLxScRgvHAv
AmNOV6RMO2pn5NYfj1FMuofTf0/AKlpY4tmLEhY3dGdpWy9/H2O5nZnsi+cWXvFX9Mv+Kij9KfaT
+pEzQPf/Rt13CJ/pBGpeHjvddTVnqN+b49cZOooUIUuhRIWf9wZj+TbkCYW7+zukVHWc5zWOVPnJ
TS5fXb0tAg/4cv5d9cD7YKeP9CZCa7JA8yE/5PG6f5HRAZV12cpsgbkVZt42dKwYG+zSCqGNBy6g
JLJXwDxFvyFd+Jj0Fy1Gv0jQsCh2aUK2LmAPx7ZcS+FbHkdV+baRdt2L+6aAzFJ5TPwPKGkhLb3o
EJgTnRxxSB+psBVF42k3A3GYlExDkroZLiXmo1XcxTYBHbiRb64HWRseGUELPwRr1nlNe04ozIiX
uwj+quj3Ig1QscG7MOBeMJ0iiGeFHvsamleQFnIe7lXs6yDr66MEoZrN1UwU7Qtkm0P6X9J5Uan2
F14OA+7lN/yuTQTtoh9lmBG383Mpt0wQnDj0qmpAw5DD0UNza4b/R6M1+Lw+LwhV3m5pSZAGH9HQ
3JkxqyFNB5pf5+jwQ1jwnj2XZB6a710J/f9o9O/2rr1UpT+KHPrRfhrT4H9j52EMra6hnfrFYmBS
yRPgFuO6PAEt55Bc7h0mrNLodqN44XVV8KdL7e3pg5IHncTC9IJxlHb89A78xIAVa8SGCN4TGGtZ
lrnLZFIp9J+BtIZRnirnePgfDBJsK/akp9Y1CkWhHJVs1HMRq44DZ84SPG7mBzB0Sh86Jlvt7tXe
u6rWNxi54R31w7Hp5Tz/Vh3q5G52iOmtBuAhFT25bH3+OgDRWrb41FnL/HWtzbeHlsN+bkNbtRg+
8nE4r7BZ/AKhzbMVAOC+LJAubze4aBW6zUHXU9uY6Vur/N9RlCB36BdAESRJcPKPLVVMHiB1H4U2
CZmYSuopfKuOw8Ba6PnspbIivn2Ja9BG806o7nIkSpo4BBnP04FVrf3wTS17x3TQmi/jq05t0crQ
ykXaEsxM8dE85KgggGqTpBqDh28OpBpwFTJgEtWn1nKbL4G13zIjUy2SUwucaH9ywhJ6oJQ4tMxd
URbW9Aclp37euZdzKzZCs0Y1xpp6b9jPJo+B2NYx1nIofB4+2pSGPRgjpthURUoYHCsgd6L+Fb5J
nO1JxTZ3+UELzW/KEl3HJnE1IRLkQE9uLEdnGkjl57dhG+cga9xyVnwX11mUZOAAQu1pDKSNq9W9
SEvuGRnJ2CuFinmUDyMgoo2hXhqARnYTO33faL0/Zdbu/nBrC0sLJaUqjuERKvN6X19aSvONI1X4
JZ16zCmJohA6QL9PDko3KM+l3V48wgoeZSXiM+uwANQi/U7bLuHdn7z7hN6GM03JcgkptzCG85Dp
/7y8w8GX/STbXZ+ZDTxwcNYdf3T7giPmehyTAx7wx5SKan2o8m4YktaumbbZi83DOXnXOICzQS1p
5xN8InFK56TpLchMGNzUapZ42/lmbgKFKiitkQ6NNeHzI1sJj3Sw92iVzWD7Ahsnue5EVrey/LxE
Ws91RXvteZBo5imcCgZKYC9Zl8lRXezeQfmaWHB3Y48EpwltNi8srvxiQY2/Gc5rmrDAkRekuXFJ
U7bPxuUHwA0U2e/nt7MND8slT8wGtinBrZ2fn+nPBE5MbtdZZdQcssT8DdPA//kdvRC6Upn6VF/u
7PmmfE1OYuHeEM0BEdQU4Ed8fiJFvczURgX/omrbQK62ySK9+AGQU5UCFZB4JWS7mH6LzeGWDJRr
+rO6TFlnNFj/WL5dhaNdwNRNqLIeBW3o7RpR9JrMGlvco6fZBXKLhPSssa6DhO89dtE9mkIfrD5k
uJUvtlhBtalkyUq8G25HWllDBDUz7ZujbC/XPAF9LJAE83TgiZJpK12pS6LOVyF8Q6mJwWkq10lx
KqTbB5NCGMcrJr7Tehr581PWlFLchg67Jc0ghcTZ3jCP1XlUH1JH421c79/7IRt7sticlwOZlt/e
dGtUJkXj9wW735AAZs8dW4YoTB7Cv1VNH/v9VswojHkqsiYn+Qb4FJ6g0CYq7b9wdV6vFoONUvrV
1JZMN0CJfydblrDSBNBn8x6W9iHk+u0YrWWnDtuWe2BodRLvVKYEDVoZUdHfMazaZy6DlDuHY/Fp
qslyQaQwV2TSa62kUchDo8/3YZ0jeCoeQwUuSH+l0eRc43dmJOOu3x9n4+X7S21TPzWK7NboJVwz
A4qhrt3js5xNRVO0faeiUmc8kKTghyA78RE+IGe51yvTs4Q6uvERaahGEHlOtwEgx0HAmTUYuqiN
08lYehWiekpkhew/anGoYWPN7FO2hI/7ciBUWwTZE5v6FHtK2sQxWqYdIIA6jAmnA6j5gynxP2ka
XUV0FMnsv6a+Bs6Cm8eQDHkxATs50ePOtTgk0O9FEn9/2jrwsAKzPazbLvSM/oN36nbFd7+eQnOe
xPcQCN0PfN6SmtOhQtiNDpCta5/VZBOJguKEpzUSCEyLoeods9UvHO7NCFW2iw3mZPwgEyR6oC34
iztL/5yMVYgdfCiyCtY7kMO8AKuAwUQb2+KvsGR3N3TisEo6B+GSWq9na5kRn+RhmDL7i9298Sg8
blxY6uqH5casv2C5gZUVRW/mXNUtpZwtJZ5IUXoUBwsTBdF/YiXXMc4Ji+r6SEz4I/sLxTvwd38y
rTeA28kcmZi0spBsnema3vvxFcu49oecTw5GzirQCI2sn3T3pVnNSe5o8JPpNBDTrN0lWq09ZDRk
SnD0qfU1ISLINNNBSvolGPnwcVZh8Clbj7v0qhgus7zkwrc7IC2UaWb+vcsQz3WVfUcOAMDki8rY
2TwCiJz4SOYTpTkRXCtjxg0D+07MSYMGmJ4Eik0tq9HflODBL2aP9OwacA4tIVZVTu9rZyGf6K8A
Q5/oJmEiz8AphlA+a4ZrePazAEAB2i9lpaFxJwvrjBn8FbPacS26VtXENsp3xrXzdbqEPXJAbdvg
bPCPavJJlrq1iDrBMvQ3NsuhAunyyejJ6u7PufKSwsur2ug72jDuXf9D1TqGvcJOcwPxDfO05UYc
BMzOg3kl7iBywmSHkgGCBXuauTCOecNT73OxCFA+CUW8AWh3FrKF36+nUBgIvvWJsFthXWevdhjD
x1g552pz9wSNyt26o0jXxTmUv1tsgFq+3vED06ekkZMHFxPHWpKJbYHnMbA+aFNjQ3phy8SIw/3s
9nFpSIbyp10R6yMGz9hpzarqdUN0hnROdbYvooEAhruErN9EeSXr02CFd9I/gG5BVRcRzavE6DIb
Cy4UcOFRo9mvlhYvtNmATvzoyEiTu+8m+pKPn/YocVXaUFeHm1UWkhBtk06Dc+MdEUKKUo/cKQSy
3S8jHskxt6RrYbYmy9RIHoyNF7cNn1ETUCdpsB8UXVX3m5FcBwuURaqcD0jMf0oDZCPdR93xmzIG
nHTl3QpBZUmzW3Qcrh2NG/K+qvCaLtIRngsfLQHSjrqQDgMgRfh9r4cZS0eFSB0mcUg99Yq9wXcD
elASLpaLmxmUwLQUCbySvy6JRWeaBE0pzgqVsHnZ4EQIl20W8kN/x/Ssqf05rgAk4PiVZZ1ImJDk
OFCdKmcF35JtLijCcYDp26gteIjJEMhSV0GH9L3dNj+7ZDenBB4+JHnNamg/Dvgj2JzA1TDS9esh
4kxckGUVi2LoEOBwwHx2Wc6e98h9huDaKmJ5GpCl5KWRM6KF4NaZeUZ+fZ/kOmau8fuv57/uRXUO
Aixx3WLpmmT56DK2XCB0fXj1Zp61TMNGMdgzlmHFbC7XDa4RZ1HRPiHvdCpPbT9wEMpiv+vLGoDt
a1IJpKfp9p1pPXYpGE/jWUU7r7Ej2KtC1nHQjxOT1KKb2A4kT19cQpBrA5Wdb1hSgkxlgVAiXZAO
x+lsvQAMSDozISOWyWkvI8KbfUt8u1sdZotajiAE9qPbwoOaXI9brr7sNnxSKvVbg5IfC1o05rA4
46BUp4lUFe2PtmlZ2aQesqQ9UpALKqoASvR5ZHLsL2H8bxifMBUiwhG0xEG/b+KALebb6vI9sW8m
5xb4rJ9DqTIcCGxuXYhzEuBW37YExoD+FDgmE/kwKDgBoRfhU7Emhzb7rDGV/UrLdqN6V2zAKz/j
ZF2fVmxwvuB1gwpNKzQShgZZH+iI4NvnLcgriEuRXfAvmE0C/+t76nGUGM/tbCvN4FqHfW8ABrVD
6+3w4IUbyFDbDWukaQRskOBJi+JjtvPVZLXPEh8vRh3vL8yusTI+yMYAdmsWnUpaHCQGX1QQFI9w
StkxTKX3/BohsDrc6ci5SBMcZTkd4WLW02tOkjeV5YtfDLuhZm5WWP5P4GfFyejkYzu1LrBllyTR
CbeK8H+MM+BBMbPaFPDzo0DLW27A6ha9JyAztQkDfbfbAARCIrYpluCLdL8DuImUm/ajFhMdaJfI
QOqtTnH877KMfOFPuJ2nyhmeHRgC63613HvUQj4TiK0+eXgXjpdbNcakzN/jMa4AWM5flhqjg/kK
sKh82JSwsbe2V0r3QKa3d9178n5UZdcyMo/6e7YqQ/ZCeQiJiZaqdhNC3shJf6Ts7LsN2RAzBePx
iDd1s2f/ODoBmBGcoXBN+e1bYdZ+MEyX65vvoJINj9p3/bP0HwtZoOZwUrtz7Sod5h1G5RZJHz6V
hz5LJ79Et71Pr76LvKPaVwfmy38hhV+UPJltUiiF81u6TdF7EDmO8Pyyqrwlqd3YHe163O1PPr9i
ju+oxWVH8wFgaWtWx8qZs6yhhK4VeiVS8yBgNNYHF98t8VnuBKc1btsB+u4dRUQ4YC4mxr60bfSl
0dnklOx9hcvdoPjAJxH+53zA2aVmxvOEGMWu0Jv3Clx6YyYSE5dOThl5mrcQWpgkvK2vs+8kzVKN
CzN9k5a9TTs1lukCE5GMZsikQEFtUL45aqXH2XBYessq82w+iVG5yZlw8iZ3K9BMj8KaCKjqvjrv
4c3Q/YKooqqDuwhJM2UgRQXC+Bd1+NE0pdGPtSytdUwt8VVR1dGClRIh3JlQnDuhVDHDjfmFVOAN
pgP+80EjLgt3I64Ibhu79IaXe83A2r0Z1kR+q0W6Eodj6RZIXgkitecf5wrgLqL4NOoRgqDePoRw
8/VEFVNSdg7Isju+0oZis8zzbZH2bc/crRr6IVLXjJNgj9c3Fl7cI+FvJh0Nn3SCy8ifqn4u4eSa
azsVygOJKtEicg5IEM+J9lN2xDbtijsyVioVu4Y5BSvKkPwA2WNzteZF/k+21LzFOmxiWNzLwUVb
/ZP/hTGfuMzqIuZTuGivajJ18cTIISqiweLpO6U34a2mxAwkTMSf65+AS9tvxxyKrqRFtXhGxSxO
2hGH8XQ9yZQHqSny6/3vtCceJitonPjAXtej6vsEWHcAykZu0eEUBceOKGNQOuXCGaDr81fGNhUJ
bOTOej7bTGF5mIf2v+3nx2qH7eWLsK9xr49tR1KPTbZ2feUBoYRv/UtT9uiZjDSoIP6GcjKofKES
hoSukMseNTei5+QVRl4RMjWPFfM5mLuVkSYQ+p2fF2wyRzdSAPhwRTtPCGVj+ToGSC7SBwhSLnfi
2lWQWIPQ7usELEizNH1+fTv1DL9bScvoMHLmBWDtgGnXvelkrE5vm/KYp+aJq3OyIFsaf5xXWgqn
8vGutIsbAeLz214fNeHjAZsvJPQRtWZEMYIelsbV4VxD7gv0fvzmOw52TVvRnOm/PKFIRan00pUz
Fl5+JC8m8cpKZI5LvK3oUwd9HbptEKwvvjoFc6Va8tSuinU0xtI8Z/2GQ/EyNgatevjsbzbmjDqi
9lEGHJPsnHq9kbR8GamC8QEzOmQXpySz97HXPw0Xvuq5MuEw9CSoLq7y/VAQhNCwe60by8l5VBSw
iRokCHokTRYVVdSlkw9a1TsQld237hOaRSrzxjEJJEI1ihCLbT94+xcFiSzF5LliDlwNBWpFv7O1
VYCuMl7eHDDQCBFc2F+k7NEkU2Y9Hdb3B3Jn6J/ctT5ckiDsXDtMjkh052K+IcOJGepaw21SnY5U
lBN/LdUI80KqZs5Qk5fc36/4MKpTJ8s0EVzwW6Fu4VI/EhJPxEVbr3f9g/8XYgkTBaorZ0apkFVO
GR5zPt6kHJY61XKDVsv/l3cTVB68uIkHg52AsdOkQ+cAZBezVzsif9lZFMdftsxe7lBNQN7yM5vx
VK8ExshwuEcD3X9cxSHzCfVm4ct3hPYNMXC0YRzAy2NPNHLxeWMhVlb3jjLP1G43ca2n4/mqPXiV
VRxBFojBtdODRiJYK+aY84KRZUUBS00bsg+PyLD3I9X5wNlPmVStDpC5TXFEFl5MJG/0NgD1H3j1
Z/99T6v+gqmqUVN1wexI2Qk0Uw6cykXcL5yN6dlD7ahXk2FywYAkjTmUZhJsWBztPG4CpPKTiEN8
EeIwJOIe/sm8IWKYljjfjhRQ6DjWxBODY5ol9tlq3OMNZn4DUycOyHMlclXCITWWNxUWAKh1n8Bb
ATCZWsUi6uVrbnZbz5pYeGdX7nUmDmo9CYWSCB5T1sUiKPexI6MqtBhkYWuRjVjWTLJKHy+w5H48
5NX9hergZaiyBFwgJAE3aR1CX807XMQbatnpkUVf7AlUN4nN/iWu9Dn+q7Po9PsqJD5fVrj+i2Ok
I0ErEPIH2A+fafRsukgFuU0Qy9YRhqVAdhAZHuEQ9FFjARNBUYNChaqV3JuLlOTtnHiFVaMW3afu
MPYTZf4Rq5kGpUHK2EFima7pqwP7uxQzG30Du9Y3zLBEEW+n7vBvJ+CLRQxk6+cSzkaHvVUEy4P5
BnRiY9vd06gJ21LEw9dskNkTtWgMXtLZzy9zLp54cQH4d2jBmI6VQXvsPxmeVYtuyifuc0qRJefH
ccxRmew+IwasQAiMXK/D111fC68FQDvTUe8txmENsXXu11bD0UEMpEygIq8sNxtC24vK/r/EfBNc
yF9tPr/PVUeF/pSgx+b83eChOcDMNVyHRzKqnWjsZwuV2h0gs922KGLQIKmwwyOYIyhofnd9vfVg
/n14KoEmmP4Q+ty7KkZWWWtWtN78kqsb0PrG6y5g8ckKP0LiVP1ezdTnSpYeyEmzmY5E7NvucEeJ
Pbw8/WWtSLQgxGJH3WQ8EP4FI3y5Rnfy6/gXecx7EIsfDWlSBRGWom2vrl8cpbPj3bwicGWd6nH7
2A93L8ej0mhIX6CdxgDHa6I5hb0lPGDCuGT8kCdMnaClizqkWKaALT7Ew1fG2FVnePbqrBnTEcrL
R4cbTlEjfuIa1nTHMY9u8x8ObACBrBwsko5WG2O2F6zQDjFYLPHAKw/nrBSn4Ab1WmQQHyyjbw8/
a3KDHUrZ9RhOC5abWST8UJf+tNyC5WrqfEkAbhwI6l81By39+rd9S8AvBAmey2tOCFx5EiTAyr0e
osR3GccbmCdljbCIRAVeFtWkkKG1fmByprjiD7UA4rDZoMPog61uqqu4HpPSitwOOQt5TmpCFUjJ
D8emcwtRMacMgz7sUIehkrhrRKPlEyK4MZhmqV9GtpFyUa8dFpftZ+nUWnqdCpOBoY3x3c90dCqE
1gV30fIYMOJud/o74unAkqSNM8VY24zQ4pirg4eYsw8Tk1LzVyWZDTDhDte4+arua0Xn4589bLT/
LzBVKFAH9JwKdNyfpWFa3E6TPNrzQzp9HllfVZONIP6ID28xroDxbCUVaARiBbTfBL0j0P7JsZ5d
1pBXxY1J3q0oN/ewhCeS7ZpC/CKc3HCcXQz9ekbedt+rxX3WQOBNZKHmQhm4YtDXjWxX8/KBrJE7
aX5HZM0Q03eOdvOFu2E2uDq4/XoeEDIGlvGomU64nLVOWM1rg5Mihv7EK8USANsAyo7xUA34iMzi
Bk+QheENmAq3RdtWxGf5GjXdDhWihs6A/4h4wkw1Zm550+QY+/yhRayF0E1cDbLwyTKhJCAhdOBS
s6/G7jbHbazFHAyYe/MKOJgeSrlmc0pIxABufyocEN9dZAgl7FQ4351ZFQAFLggqHQ+BcLws9gc9
njSs74O63KqMbHwBV9sVVR1Ak7KwLKQsxeAzvrxtv91vry1xnL2PDCScNcthah413vV43xcZzRbS
8FSbsFdPcAGzmctq8VeDmAe1J+Ej8AIfCsRAoidIvVIEQ29J5rR4Fbzf3Di+G+/aCnEk6HIdHeNt
X/+pyCJWAqOlAa0WbHrwF6iiR+rTfV7B7Cx1YbdHKLUxlXimVqVgUVEJlCAE5C4Rfny2GYzKJQdN
7JbyS1CpiAtr38jlZ5ItwRPkt7Rgai5yd1Ay/oNDG64Mqt/bgoxZL9SwAhPx9aw+YAVA4Qx/xKvh
tMkdzqEYyt/oOaXDvvc3FSMvIfu5pXvTGpfhuqQER+3WPmIMKAxL8Kjzr3QuKlvXJZNOkxNQDBU+
a0+t8hGp42KkxyvxIDkTeGWw8KcMoCSU05WKEXrw1KHSgA+fDIASAl35cBAGd6Jou1A0IdWdzKGG
1Y9NhWA1Y/36NI9/Sdx+UwySnZr4lh7eqxGmH0Fq897vgwkyGXED1KtDuQ3OvLUTi+j5/83Tcyjk
J93l3hbtiYvv2HMJpI1lC9PSVqqvJBonsSM7DvKNroPs19zxoX1qO+6suZ0V7QC3csYzuU7Tp7zC
5lSJ+Zbd4vQKZLgzsds7gKryx1AoD/9VY1y85AroyzhifxHIwexS9nHXSTPPAnpH8gE3z8BddG8q
0aVz2TocMU7+ptrl5S7d5Ds86CG/2MG5lxhSt1hdcDPto1B4e9Z9AiT6vsbrC61BnZ0255v+HAkL
LXuF4i0/NTgjdwrHQ0ouWm/UA+xSgc642MVzhg+ZQ5SVT60YFVg5EjOYXTltP2nHZNYNezmkvODF
okAv12C86i+JxO7gWTJzVsVjfUv/a48GqWAGPhv4mm3S4+9wbYsDnXccAOh1BDKOzNr/9orIfbLe
hUUMUJzAZERzzThLe7mucuQuMnHWoIs7nJsevvIuVC+Y5AnJq16fHjkkVOcmHGI6rC1/t4PonxhF
lEAiL8jfAMO89xbKLZ3o62H0FgLnOZCAvYB7o6yJuq2qI9wPpel9Kp/t+cg32VWgBbr23AQ259W4
nJgg+0Aa5GnxqO2JBF3HYWuT9LDItqwC71nEtX3DjNCRsClfsjC1Ypf1L87PG/Dp9xhC+KKlOydx
p3VtTTIJz01jG6Io6WPamJoP3H4y7f40iVzUzuw9nK8XwnAR3QtJJKqDxgFennx17nHWaToGTrTk
d3MGdtUrvnJePHyCgBe9odJIR0/2RRP1l1M62slv5ReSa9sWR4cf6HamfPWfq6BWKG3/7mrAyf1S
T7vVoAuoN8Miacb2rkdTeXl0zSYYIKhtDohRjtiqPFuxeP0eQhIogsI0DCIaF8QLSmWwn6a6HB5S
hNb98jjlK795o1tCW3k2NYuuNZBkWj/ijEXPjQZiBjHTuk/SQ17nZ0yDm5kpQit+8khRTd5I4iEV
rieqmM1P/GJRgy1N+qi5S79lsMhsFL2kvaTLU+gDzA431L8nTIzETE5dsjATtR9uTbvUZNAYjZyK
18dc89Rznq52+Q9ZvzW+M0tZnHZegiCyBkUBWVQd3VwfUZyB0j0A5aVkpWqFe8HFri10LQHW4MCK
tsTwkGKZ0YfCQ4dJMhXnf/jiDrcjXWt3On35rDxGJGAPcYgjjFlkmGDI2VctlKFrPw5KkhbgWGj/
FcSHU/g8yhR54mu7MR1HvQJWYCFg5mFmXr86bkDlx8BzFt67J7+GtZA0kdUXqRyB6b1OPVHkaJ3u
nAgr3oWqPS4+z6Ds95pWc5B0Q9bu6GJChhAYEaHuiWXtgRKYLJGahfzvqZUg25TIgTA8K59Yqef+
LSNrwcYWjwOciPwgwK30pGUBeqzz1jK4/pAv3Hi2dethG3PGWDbMUXP3gJL9godSlIpGpUw9NIXM
P2QURKS5R6/c6PcnN84sOjmx5aee/RUC/eAXoTF/UhekKayDraZA+fVRoWQfWAxjh4FIjXnq2l2F
4HrRq6TZ7gUDF0r6Wn2pm57kuO3g12rZ2+5zG5Hb3xYF8VZKwgr/Fk/9JjVYsP7xn4uSLNkSdT3E
sclwhDdxgodKc7gVQC32nUQjnGXy/D93H8nDZXVEnjQEWtJ79F1QIe7i/0AgcLgU8ElKfYBenIyr
xawnLCRr01fC6mo/MPzZ6y5ODiP04Ow9gfu0WPbAhgBHSQgiwu/x8/5k2K3oIhCjecEl/NvVVZKe
EUZ9ZMyzjVPpK+jOCBSxJxNfSRuWV+tMKXJ2GCTxgt1+0QjP7HIRjnOqwoFk1jh+6SU4/9LFkEb/
ylsi8GzgslWTq6TIrFDieNtQyYI+fMT2a0d+AftBguzApuqGfm9nY+LN60cnd85QDdschInj1dy/
AxtNopAbuXQ92qKINDOK0aMyRufyfM0Br9Mfql2uP1L/pbdk/p6Qdi/fXqQ7L2a35mCLIrRSKAqu
hfnsQO93tMVU5rJFc6xrE9maufz2bGRQzW7nt9oJpbCfocpSju9M+Cvn/Tvz9p8feVuli2Hqe7rk
U6rE4sYRRwiNaMXBFqqaBKusx7Ylvxv8b8mz/7hvL1LY4EfrosAWmZsBGv39OnwsE+eHnaYELMxh
CsgRCJ2HUj3YPtGDR0/lndtZBUsRGoFGu9ge5IFNHRh4hZmyKqzTAbrK1KY42P3wiOAUD+Lic9W6
vttp0EWcf1zeMhoFL8JSbI0vBLMxiPKTxtleQAjXW5PqeAc7JSmM4fcZVfwkeWBQHUCrhMC9g4JU
QpZ+7Vn28VeML/XMl1Q+9ooQqIjrCB6KaKhh5MN4rOOhYQc20Oo55RaSnZtPaajqZXStladcRtyA
LWEECkNSxbcxn3yJOtVO2Rd7H3HcvoAS0EDhb3idiHYohOvfopsQafyHJLHuc5+cmIw0hW9/zF1h
hsz3JuE1DJf1DL/YQB6V7DuvnT0UESly6ZxwRwatm492ShEAwCkcs4yYeUQ5oLXjao/obMubxnO2
48vLtHTDnES4OIhSxPYStdtdsc64RtdQgZNoqkTtP6jyQkddvWchOgEiQQeM2RWYJDu4/KvY6Kev
tMM1bTfS35YXhxbNVS8XaPVHQ+AQ8Kk6clVKT/nnAE8TkqXbOTpVgSAAhfyGUhXvqQvNiPr5kKmy
mBpSokji3syKiksVVFYBf5MwV+AYZolqNbUn8Wru2HbzcjEseUx/aKBvtBboWo2qOz3EV9vpZi32
lFqgdEekXop8hROyd702DbfYpOPrZ5hHsFvo3C+dh6lYfAujri9zsye3GzkwxcocGURx4xi3r+Gj
aAEz5Uo9SH/CNv70jKT162TcFsUiwiyatZsKA9pwI45uOHsbNo9FKDA2J6DYNzHWJoW/2uAxGf1s
L82pG3FnHhui11GflIzovzz2WiGL7ku6Gd1zv6XhKfiv95ceOnApq+qwYKBoNk8wrqVcgbMI3dT8
54OzODZZhH0Uc6hn115QJDvQWsvGTW0jf1wzojA4kHzReHUFVLJSestdXsdQ5upUDZj3Zy299e1S
zDPtCh/qpsq1txwPnfyG/PcEIqYeaCtjXZm3a4VadN9cvupPi8amORL57C8T1fc0V8Pzz85bL+3t
uylf7jQDHfG7RFWeZYa0vPWAUU/xPRYZbhZtwAj17PrpicMjVDcScF5GELAaYMrnzbAqZt3nRu0k
2cadoIydzBtC09L39MMMdUmkmLVM+4qTGCPC8KjTbFeFKrwxCDvrKSzat7Hg62pRs7bKvMR4Nfv5
H853Umm0v1fcLSunS66abXpkjhnQbKmAJ9xLvKBzqOJ+2YNMdRaEyuzTczA9Tr67B9dPkrkniYh7
QjDi4r0dOaAINU8Ruzt1nq4hY3+/m/LxyXCwxp7U3JnbbzifdbVugPQs+uw6QsZOf4YoAzhtEfZg
DiprddTerrDSPKAbvpe5V0eizZXuugQSflRHbqo/Ds2P1QppH13XjxWbSo2BRDO/i8jphwMZeMXO
gFKt8laEg+vy4ublWFkkzN+secEYXHiQl9uNL88GkUNpFqBUPZJ8T63DvfFwlaBfZHR6SdUr/BAl
W7INJd+ETYHThJuSc+QVEwPTZD57lfQfHfuw9grTk4asgl8fH/6KG6+Gum4LKaF2XOLLZRwSrA9U
T+rZ9yH5Ng6uWhubZ6RtII+gWsVOrSRBrBE5BYEvPQ/qqvhx9MkS8zhoDvseOzjRlNNIU47WHPSP
zUAhMytF5MlK/Tz2x50HhybawR3X3IieD0SmnLTsyFTl2Wzz/OvYaJPDZbx3pZ8IUll9RahRcize
m+ln9UPM+XggqTqtj0nERyWE5eCmR+LaDJuy3jiEqzD+x9JLh7BWwvJosVM2tosKO+XqB1Pe//Cl
/ysUBxHckM68QIE4LIgtpSfehCF3TbrsDZ2RDVKGkycB+jzBToYVefRbO4ZuaLCKggrGlpBIHGkX
foYwzFoaa6wy79V/O4xUwXNUfD4lQ5j3ySVVwmkdvtcMLBlAgToyuOQKHwZqN08Sw3wRw0FTZsY5
q2zsEeapMdBglMKyrMUNh1gT97aFYhhPMUAbCqDAN4UA6naz4ZhRuWHP0wdKlThV9oFqF9Rt3siN
RTVakroomlIDH22cnFG2/oKaXVfB8OYMUUy2TdqarrAdSE/mbOusAwmkosdBzfbYxNfItpyCTrw4
7yNP4iBhH5EdCXNDwfPDJQp9qdUCD6lzTVn9zNMxPjLiVVbPwNaOqGjxF6ajJ5NBXUZNIUN4yhLv
11UkixSzTEaF+jVL0VzPNf1fWeI+ezKb6I4semh6IE6VV/fFD/4jGT1rjPyowZyxvuqmRV7wA9Uq
OgSFfSZjDbXz8gFz3VTLvGETTq4K8m31hbmLSZPexLcO4FKiur4DLAsssiYL5L/OwKNoQ7/NqaHZ
3LTAyMePebq79+t7rVTeAci5SzzhycPKq2l5eEgskg+43NfTPKf+KigmBuAfDr5rL+gZ672wz1yH
C23DDE8s7PI8Ev3Gvw9o2pr7nY5DEAdrfAiyODAffqgIA5r4lt0XklWenPphQ1k204LXJsa7/YVl
MBnNc2PyfTLjssuo1S9I2q5UMWgxblqumH7f4vc0Gyak1fTgrSWON/ZWATZPVciEqewe+tvN/Ckp
59Cbohf5JbKnHVA4c83i7QNA3CDWjKHCZrsmCWEbVBl0FH+Sf/VNqI6qUndyZBySezs3EioOrR0x
1/7fA0JSd3dilj8tILnpP0NW/kSAsMBC/Lb8lorn/51ruqrPYV8VR7rsJIdpEetHMxDoPMikD9N4
gW9aBWmojNZwM3QwHvIybOjL6rNq5Oj7jKEcPeglsFI6Gc2UBPaHesr3jX4YYOt/Y79QtjUC5Sj6
a+m76ivyGIXEeYfCEA+2BRUP1RCA4P95szvXzfDh7+TXI1/f1PBBggCd1f+7t1QdYFe8JfMUEL9Q
6ya8qXOtTNTftujRp44XdMZjrskJrd8N4Vt17UYN3VOndDRWW8NLOBzsrgbfvl1PTLHHzwBFgbQI
KnM/Z0REA2T6Grp75NLkCdDAzYJAD1piPLzru2S27k1xQIQHRQwJCi8RkcqbtGQ6IkhM5rraetK0
GV9rWo+4vpDvq194zPUy7K66/QRM0K2gy4ZdW2EkMq2Q8rfeWxllbU0fou6QP4O6xKhzDCjmhY3h
/eLmvp5RDNLGjVgZgW5vPlVwbaV7HxvxLebUxai43LmtiMbA5I45p7mNTsJD/TZorxEyTHNmaKd/
WFisrOhSX3OPTgBUnJwSUu2kySoZmRgd385xD0RmyC+7V05sai5DrCwlozi4xptRCrN8UqDF3IPd
oFA1TAZOgpNIZ/uRycEAqznu8vCuXN6LWWmj1+OqHZkaOfpu8NV2W/4jZMTOFDvl4C2YLzCaxCb2
1zA3qLUDwAiWxZfb4bpZNij6p6rLQX16lS0z0QdjqW6ajMzFATKSFpyfgAz4PVQU6Q2l9EgYnOm7
/5Zuf+IRR8l21mEbDPKGBhzIYSL4Q1nNG8WyXj/F/FZOeAM3OpClSGTJB0gbNk0Wz09qYCoKj0hL
FwDPI96LZZ17Q6uJmlzzIEOcUfW1eikbs7niGoLUuZTeHlM5TromqQn2KCMQZZ91HLH4sVVnfA6F
GcLITYOZtQElu4wrdHaXxgwMaZYe5yi0d9TKzcmEzxVH2D5kAfVJhO38AxXfx2p1UENTOikRPhuq
Ubn9QUXYpZ0T7HxuEXdHqELqlTaNNJR9ffKZ+xlAJh4JugqHQFBsobt/ceuXlrvfk3xjeOSodNiD
R8oTUCa+L60uySiiQEy4NINxRZHcighBv4Hg6IlBkoMgbNmrxF8B5G/1G+RbmkocL2ppvUBUu/o7
qfhLNGjnd2EojdqjqGyyZCZwZPsiDynX80q6PE+Gy1prhYRSjOwDEgTGL+8DC8WyuMMJDhhEIcnw
IiwUGbag42IETj4wfVs+MutXph9uJrSM55rtA9tjn9iuC94zaaZ1VesDrYaoecjl3Rm1BTDlXe06
6UKw9QZuTGFkumr1kp8swx5gv+2AiLtnbWvlD9myQM5MgUWuuiScubIS957DeFmu5dljhqgOkA2h
VWJtLN2WU3f8ZoTSPQKRGaTgGW3e8sVH8gAl0kVsRSnb3vIUm9ASQFX4r+WRvKaJvZ1xbtBYva2d
NbWQU5f6an2K3ASedB3MdnudGoGbB2SB8tNrlZblnccP/fbtmgxUZEsM4PNBFRq5f/GnqEyhnWhn
0U0Kuj6h8ZVc+U+H3PBsT5ydtfFdBV3vsSD0fyxhJ1JnumfW6+/S9pwQ24QogFuJuhmytXcAUm0z
KlbzWHaRa8Ii1tMKnNgwv/XpjuFzC8yL+DaXYGvj/fA9kFaSJcVNO6ZCtDPXNnXLJYKQiIl1Ne+K
8ITkd5YSeQZ9ZFYspSxZAuK8JY9RAtWke3DJL79yu2Q0HIhma6SxQbjXxLXvK0zz1GVKX1QnUNcM
sjb/I3OHc1DTn+ohOldGS9ewEdtYeUA+DyyvlPWDioqqqDI/hSk+CX5doti/szPE/G1CANknQ+1L
9v6TWnMpzf3GLRcNMxbrXHSH6GRtnwrbdkXydZV5ZdP3fcYK04c0NXQZHYn0Gf+cUMYV8yXob6yr
29q/PJRs+6fe0AtA8TvpzdNTbTukoRn8n4atuA1b8nM9kfvYAhccX3t7ujfjO7Bf6UwmNjDE0h5k
rHpe/JcNqzfdZBkPJb6slAHCUW2FnigDFrBir3tU2xeVx7lRb+qFCIzESREfGITDZ9a/kEnHGPFY
uSfVTApJR1gON3/Wv9ywvSv+lH4JYwpvmSUalgSMmJV1Go0i1+NnmEBqpekjD/cxq6ra8e9kgRoS
fZpsXq70HMlZ2pS7nSSG2WJR8ujsunOToL4fnjUuZxbV7az2uW3Qfe9bVowY/I3kSFxbjgcnV+NS
/fUsw52LVNmbrDngl4W6jUbuNzOxltfsxLf9nbuD9xEAqqiRL4Z8TRIqWttGnkkzDCa592LSufnL
zCMUO0MbQKE0huK4JUveN3QTnnk6qlOM3X5kh37mT20oEeOMW7jb7RnMT63TeA5aLSrD3s4AlF5F
v9xFgwCk7E5q8H8rHwDR3S+2SEWIc/AUqiD2nWmAZ/NMOdqMvqlsMGs9XF5oUnpKhDvI85uX4tK3
yvwLQOZ41g7FkPWqKDFlsDs8/ZFRfMDx+rL0knjw+TRbulnAMMqByUz02XZSDRMRS559sYFH8md/
bPAytHm9fPiPZOjT1I0itlAwdKRX8l60lHY/jiRkOwbCjMJMB9xHX/da+F2lfQ+/lCggVHXIl5Bj
m1PEkXJ+ClKBTKOKrj6HraFF0//KKgrfIHVF784JC5ofEqMjKeXSHOIspULovLngS7q0fyWf+xIG
V6UPBxFI0k2mlUdE+0Pz1J4A4VO1GR61RZwja3IjxGeTabPD75tvETR62r9m9VfWw7wrL10tpA6s
AUSHifhI6PTemjlYiOXnwiW5DoC79UJU+y7xDPsvcGTALuYzIC7RPEzTfg1nZEyBkgy9E+LpRwXS
KjkGcZ9Gu7FFYBgICqq+0wELywSzEZhOPLdsXph3qdEN1JlPvi17yaEC0VukNvPxL/YjeRDHdKTr
WK0ymgbzmdY0B2BUdfIjChkOiGZRPCQ5T4mq5p2BdrEUmSsf5RQmmeh6b5jZCkcYpBfs12mVmZ5g
WWF9W18r4L3H9BkKnwbocacNvzm1AVRnyy3OIz5UnyKCr4T2cBrzvDqxdexjH7zSAm2SgCjKRpbl
iqpcdwGbuACX3Ns7j1lQ04GWj/GnGVXaGZdubqT/hZudBaf1OrsAf85NWvQ2AbTQMhDw159+Om/3
D9tWe5J80P6210VTcRCXUOs7iDjuHOHgu7Ng2HOjge8sMjJ18X/XZvuy0UiUVTIGLldAOdGKy3jP
wro2IrZqRObm1qBhX1lUYgqY31l40byeSiXF8nMob399UCsVQgRgOToj6PVxynqfI0uTyRHVIp2v
gAfgdKhfbPREa5EuZ8tKjH8DP6CXCJsMwQ4zJuZuPzsTxU/yNwyiQJ1BGNsFLLM3dU8oZ9ZdoJgi
xr2zHJ0P/Heitvi4sMQGXutQfYxSBqpf+qNCT4smo/YDZZPgpiBPB0Yhx9zv29E0508nLt0OYCrt
eb4duvnRbQgPeIytvl/OFRGiL0m3D/BIXu1sM/dcXSkGmwHFSrM+ea4ZvW9TnMuDDjuVMQyxuWnW
1fYqVAHNsCTdVXGfXf1ndXAOB0BdMcHvx1PWl4I5gwAs0qwfvlFKnSseYRsF07AzO1E6a7HoF/dR
pGf75pPK4iVCdH4kwKhLKCfGm7JgUazanyVZyt0P040o//SPhhCBcsTbyFwZz2YZr6xpE4x+IJBu
G3AesnMNKEssuyS8tikDNoK9yBJcIaMgeqyAaqMFk6VpKX9NVVP31zIy4fuyskNfMAl1rS46LxQG
eQLnJndxFdsVXJi+Nr+EhOTzRpNIlKplnz5HueXvs4+XWYmYsSRgIuYqJP+1QftDT9Ed8s4FB13I
h396hBUPua3HsVv8x21mU2OxWHO3wGijkFe03g+BcFZzwW3rPeA8kR4OAYriPVhJh/eWRgJIeUE2
OvqIjHZQPmlSxTMof+Gdpo6yU5mxBVkp28qhvXFq171FTX1jKm7TQXEXuO5ndbZKkhf4qMkdSEnz
LYAwasw5VcGb8MFp91GHS0Hy2lQMrNG/LHDMsrfc2qTUMunJU7qF1cMrjqKckh0sJ2eNhLZRHsP6
GNGdm98YRJjL1ZwFMU5Dr0EjQbHkFAe0XFbttF1P3+C+WtDGq+QNV30HGzwR3ymUqJIxv1zJn6Jq
QwkuolBZK1fkltPz8hP5m+fVsIimgobj4+/4rbH584YJKmYm594DO3Qs51zsnijfNc9iKG8b23qB
xqQdTkHLjKtySS1Zk5SqVQQ1lLCx/BWus+efT/ubmhL3T3SdFrabFHjFqGlhkoPab38E8MWCuAVt
kjkzqgzuk4cBKpg8Rb1LyWTdDS5+6BYt5dQRJsDHteHDhqlRFVy57niG/nJel17waRAnVZQRfjJ/
/e4+d0LQx6ZDcnA1UxzfFoKID2GiR5iRqPBupwxCmj51P4cvLUkteFXSiyDnoV5tijNj//WLvrDD
N11NPghyj/fatmpHUIdys/mkZj3+cz7wc1FHa8QtPMssPGRbgoHS5tgn1u9iVON1WIubC5hIDMoB
1r8E0JRHyf4BIU0JXziZui0NkATYpAbH2vJn1P3BJOp6LRNhFsmOg2qzrX1IjTvn3v7wgdTIHqZo
CRTAr2ooXYYaUqO9r3vArjSMUcyQTJTUFGUzFXot0WH6la9GIEUG5tlEhwFtHCot2CVGdJbIpJhU
CFal5M2MQ5ILbGu/rw7mGxYGix4CZRhrmh5ME1s1uRJ+2+ukZDRIJIiGopU9I5KJj4BMVZHVxUkw
n3EnGTDMfgukAsG96aAJod8Tm0+9DCIOCoD7WjbEb8m9wIuKLqmeSE71V/cAu81YAkLemdRTpu+N
/EvQuH6cBMsiGWQE1ihtcz+5d6cXPuVM3BYFGRiK01dWmyRKKW72Oft0a9cP/3u9gU/wY6JQZtqd
gOdEIBZ2XcnQJhvTbURR7dmFwvcQ/35T0dXfcsclIcg/KBqBSpUFdqbZxnejkiasLakiNS/eVN3O
FXZ9hn1dsi3QB24TXzoRm2j9OElu3qrOnIUthA1IOdiE+Uv2GF+XBDcwZfB7dh6j6HPWRcbTzKP1
Qe+60EW3vzWaf2jWn5XdKjpX70+CHWDtVO4ElEpVvsJEk9yKkJKA46HruHs7UpOezIYr7XJfdnTv
t9I8z8JZF4FKbe20tEq/7HXHJw+qfHD+R7mrbgbVKemAW0obRwMWmD+dwR9G4gXQBfgSQpE+/euA
Yr8d1r0WN9i+QRL7xEW1ediyB+7Ujz/DIlp8QhQRFTdji38jppccQNSAKbfnALCvS0W1eP56a46F
M0XuiVUH6Ux+qaB7GA6wSaQt8uUgypLmfRtBaOcKl/BZDZuQgC+FZ3yJsnXVncsnwUgHA/j20piI
/wcUtGGhgHE8DRFDTzvEiVw/UEVNVPiqgvFXZA2KPpzbfjaeAZeLZO/GusP/cCr4Tf7cjZwXy/S+
BKIq4+JAtKscNEZqgQBm+IYITjXHC7SfSDy/UhzxQoFgcOQlJ6kHxX4sAEs6qBAVsU6Y540Lqvu3
GTx4wC5A/ns3hd/IV1LDoA3cU0HPPlWHLEb6VNBDZEyVDUAq70wzs3rEjWOxoKHZN1rvRXGLhnGt
QC11AssSXh6d438NqYJWvMA4tERRA0RpyvbA8zzRL+miptdcnf2SGQAuY+SIiGzBAtv0YDjAFTQ7
arZSmbUrNZeFVPWrn/9ChiW3tSHg9e9syWUIEpucnCdaXdF/T/vQS1xQSzL3ZeT8o6AYxxBn0NEB
yPP2k3OEIdHeNtqLQaBOn5k59ZMriiQQlqljuoVINN0gaL3WXiRA9bi888Gtn1MAO+rJ78Cuz1WV
PmRVCvYpfAOeszh5fPnld2E8ETqSAkgbrd6jmptznhrzjopooKhihYBoekjvX5AulvuwmhQra2n1
EIHdYa8Xl4WlFlHjTh/rAhb43TWPjHWi9AXis/CDFJyVX3umY/QRWVEs4V+TJvu23L+f9Ogxv17r
HbBnb1tpKziXB0xjaWSXn8RqHXgs0aBFZVIlZyhxpkTi/ReAYPPje1Np/OizO/P6PAF/Ok6xjhAq
2QITSzGGk5FEHNWR3dSYuubX06ib4zafPQhb+glah1+gRAnwpXrMrItNNlNlC3MVzh60BfOftD39
7Cey/ZJkOvxEeo4HSVA65aKHXy1NjaXSewui9Rdug0s9NzCD+6KKMMgN/VP1Ev4cHhuny8scbXhp
hws8A65VwHzDF/siy2HOId2vI0WUGsFxEmxWgPoElNeKpCnZVKjjBPGKTlkjRuJ3ZOj7FBwrHI8a
PKuue2uSdQZzHb4Wz1WKAeE4BOLTQxDELOKzjxwn76KuMUvatPHKg64kxn26QK9/o0SrWUguiCpd
GuQPkP24GT1UiIviL0bfkzk0j+0wFvtlSQeWUrLeNjlVrxJzM2YmdUTSHh/nF1NXKZl9rTTcBYd7
cDEAvRSdC8X05bMpdEQgFC3Jh37Ii0xobFleLKebOTSsFw/5J5zH2SVQdiYhjTm5ruKQQwwXUcWC
0ckc03IoVCEI/xAhFrSl6Aip9fANb5wvjalJUjhRbspZyz46I3HeMrL0G5g+OZHhCqAT+dhvTKPO
rDSG92ZZiAdyQR3PYi3Tlvz0tpnl0rHNovu/8ag64RXU7vGgbtVUtXNYh2+GMHoehoZs3YhFk9Zf
KboRBpf/ex3/g4RHV28YALdaZGGxxaLgfW6Mv1MrYhw0mW3gaaHzf12AW2RqXq3c2V5NHjrqy7kn
HAJN+59+V3DwrBFwKqLMcxPXyFb8kDEH+Oq8hw14vfmD1yStdRP/Tm6RmfS9tQTIkC1kZ8Cn7/g+
yTypzg80JG2bickT/gT5d4/aVSeUCnrzTzkwkwsrFQmZ9e9Ip4M2BtY2tOMT+3tXtUbs7JrQta1j
sFrKz5fuJnI9ifjwzIox7AlAChLdNMUjNpWkhgKIAAc9reOj5hyFO/fX+ZIa99Me5KPU/CYc5GB0
9pl0g6YqKlL11W/YVteEs+k1KMajKq+B0HflD+FEjyGeeYPYt8DMGn04xdeEyEoZMo1OpVwCvwsB
WQviEo9y1q5LYjkwWLylO78nFPbo10Q35ukjALcsNTD+FqcyxnrrXMulMFud+X0ncZQSA+dvrrJH
FSCRfCLIym6bicYcjlLYjn6/IJApW35r7AqiwRNL9BvYIDHEFtT1bCtx2nxQ5KsDGK1xGzYQLRpV
O7P2e67w4YCurVAfy74CY/10YL4IDTBaMZVfJtts91eJoRzafrXfvY0T/Eeuan9DPImL1dclVRtJ
qL2GIbbreG8OU/SU/66WzB/Z7YQFqIPcV2sYk9ycCsiMdRyLONYk4xRABOL4gSjGzpwmgJmhSWIP
uDppjSk1QioIHaZlnzQOfnSDOau55bkNRaIFtW4qmNHlI4yV23TTqmy43D8UNIoNTI0XuKLW0TJw
gwhE3oB6lGBUtfC5t5qLv63zGGgMiym0lTsXIMzaQXRurfrdoqUYAlgGpLofB2rsETUXcGP9pOYk
KPVTmOMTUlDBKdsAGTwkScRsHQojVUFfXb5e57X469fLO0SpsXp0Z15WLKXwDUiilqOQjpClakHJ
7abJh6QIW7pe9mxRSqljInOcHwrhWGHeVNbvV4YlkKtmuqFdN/tvYsxQadjdXxFQttGJycGN2Crv
o2khV/YXqiHhkMk3u0hCIaKAdDUax6BN+MIzmcO8nLSk5u8VvAnj2IJWCCTaGtIcQE61xPXeeE2O
VgU5Yq+FBY7H5bh1J2cDmHmYp7Lfh18otE5D+HCwQxnTe5/wUf8NcP9yBhgpNEJF5FNOsWRwfBV5
2qAFa3o4kR0c86f4nv1t6LmJBnyeP6tU3Wj6m2Yq9wBOyzpmQ3t4h+LciQJU0Jr1CaBh8IhbjnYB
7jLvSx6PmUMzFdCXbRAKNcmciza3lwiA+o+V8oM8WO4DNyPdCqi493qTLCQi5Y7MbK8zvu3nhukx
UIUGw2KGim6308mi+q05bDL+9DZEUIVv9pAXWG7AS9JIq0FwBuPgjXv889lbAuNsmHjoPs3cVbbK
Jk1wMX3+5F7iK2Pad6FjZAMFuCsKq/k7qZGNpBekivKz4iP0B6ENoLOltOJeDOqAJMRYZaWkxa09
EM9Hgxh8MrMSq4KVUC9aCHamTKWYxmkxGfOHhejAOiccDC2tAYi3+gQllB9TmiTCinBVp78B2MRm
Rm6l+sSeZKZ6nkoWHukDSkGum+pIkCdXiwIyWcw5CNEkLON5+rIxAfOLX9wG1zakJ4rd1A3wofaM
4ZVq24YUn930pP4lxIiI1ZZ+f9tKabBmAZbCHkg2ehklln/tgYYZ+d+S2ajfR+m/w/n6dYHeH2+O
+hqZkMMQf0PwKfgA8Wl46R6uuyGb/fZCuOGUJ5/9e30+Z9Eh1l0AaQIuKhVSF6ZbK8ttJKOd40qz
GaVXx07/OQeanbCbQzizWYgH+h9zxnxDbO5s82mjbHuilC7yS7y5faPYoA32rC1EclSlnc3ebKlN
boezT+gXtIuB9B15nq8iNGWaZYvn7pcW29SYy1aLBLQ+tjHylCqcE7c+GaZHW44CqFtdp9qhJBOk
6jYzE8Gy36VUMejnzSJ1cIZTNwfLHcSch9QKBElLGS7XwUp3ddUEdnEABnBqq8wyITS+KdbXo8iS
m1C6vsIEjSYqFqNm/qfm0ALBWiei8s5D2iiQHoIVZlfkSCVREiH9w3waeR0/NDVoPYSgltDW7ZXa
g0SlX2Li2QrR6p+OjZYzo6f/F+zbD6kAM8s1VpWQlh5PgTwe8RgdBAdKogoL/XOkY+mpvT/ALkV4
X81sJ3FBwxANey9osN6o75LWPKwV1v1KtpQZVmi4yZO8HWilKWDyGNdrDKhobbcjfxeDXpwDafzv
xa4hsqFm9lv5LXyyXTS9c/OdIWue9Rux4zOIEtp1ffqsupH8ixAnqoMxx7ysOOSzq3XkkQxDaahQ
duCuHi9JDxddS7nn9Q2RoxZFdmRdxJugfWB58qZSgMEELgLkCkdIw53/FRCI03z9BGgoDc8yphaT
IJ/z/uiswQdV53j/j0Wwnj31cSLEJggKNcuPug/i7k7NCEoXQhcEGHGvzjYr3i4dPYVVnaMW79Ac
b0FH7Gtd8uYvzs7rBs6kW62fD7fZ8HVLBL29FiQG1m7whnJqkTomH2GppPb3VrY9ycM0gsHyZ6K1
oy+Vi8ig0nVAYwMCJIBWnDC2zpr/hmL60hFnkw/7slPVXsSPy1NfrxbrDa2n2z0rWCDxeqWsUWpW
RxUad+ouwLJTtfKZ25iu9Yw6x3HAJ9GK/+QEbzmSo5JViDieAwHQt1WffgCc3AQbICcYocb4fQQI
cmcdFUxj1139vgyD0IZvT9KZsP3j8UuU/WsSbH91NlKhJmCMEyoB/5PbHjd3WIM9qmoh39yjrCop
5mPrS+WXKGqtvxnF4mZ0YscXPnKimJ8PBUmpmnA3xcbSaeVSs0/DToJNU0PViPGTNd8FXyjnXmgl
9EC2kk+5ZgMSVqiIIWyz4J+zZhSosJ5oFSe2W3mbmZemecoi3TPo+rrjj1XbPpVTaaFBQPWHYv45
vT7EvFyCYdY47r/uiYQOogyBtA7h73cpNQ7Xvu1terBVdWarXJ30C6/nqVZbK5ZRO+io6LuuwrhI
lCHNlNYJFJuSNYEISIBpCqWjTd/5p4VOBq4/WRAKtdr1fwFcWHIvxpRm1JUBzrxMoIDEeS/W47KI
58/cHUThxJxII3sA5/JYC8iz5WX8EuHl1YWuqjufVPpghctjqOx0+jH4k4XI/Ejzb20mk2EaAfBS
CuTUDvyznGRPxGn+y1+hxq+TPdzu8bC/XvNKtZufPuQPNaiGHycSSg+/QxKczw09Fvt2Vndtnhbo
p8kUXeLe+3Gj2lN1kBfIde2/78OQsLVX60LJzZ26fD3GddmWd753Kym7Q+ElX5IzTfRV5bMi+ikV
vRjXIBZJ+fcEvjj/5O8nu/q15nYAtzf93M+9hLphEg6gFjmLcpBWJltDJxYscAjBysQeMIJnKw6z
yoV6spEnoUKsesbpCerGJinZUDcs8ZK1UApQVh4dKv/MOte+BWGzHPsQj6tN7AcO9wPJen2Pns2w
wjPk6Oo5zR6/g23KqGl+Ku74O+fsjaGXnaaIboSGrKc7fq/KAboh6dIVqqT1rUUPMcybzjPWSW19
yDN+gWVO33PrLkuEKkpNW5VJDtW59V69pHL7YDZAc0sHuJCXkos1iCz6iVJh2oG/aciuiaS5qSmI
/dTgX6NYesa5eejo+Z6AMQOfI22ccz1iy1ibNsIYg94gd9ZP9AADFLDCwNpVl2PvZDeiR3Xa5w9d
avOK5UQ3mP1DiMv15iERytl5PqztaeU4nKAlmHEXTrvRr1dT8HtuIneNEmh3ZE+gfWiNSr77BuxM
YlNo6mn2PvVj9Bs56ohO2eE4YFnFKJPLyw65k84qD4P491ia2QIbwWgK9qP7DLSQoSsUZnN79fRk
rQp2KKMlnwIhZxtCu0zAthVGUwbB7DmwpZ758oPEc8T4TJH4dhrqGRATM+ATV1IIvYGMn51dMFOT
BjSRibQittG6Wsam9da92eCHorTQ63x2GlzAsxpkyBg2BM06XDKrXctn2YlWKlkNBCgYat7fE+qv
vy8WPXv/R0vpvrfhwD7sdiUVeNO1Kq9o8fz8yFZsVUR3YokVaVSE8YeIlc+yZmSeCCoRmsg+mEQh
1km/IP7mZju5+m0Dd4GjySFs2b5thXvgr9O8epXMkVm9nr20l7F8b/ywof0d2Bc2VGiIQM+D8LOV
XWKtHBobyM8vvB9Zi9ufkqin8ZidtvM5b3Hl6GHhXGC+gsSuPUdqvbZ4h9BL+DeVY+9qKCAd8D4b
m8+0brJKK1b5OjQwx/scOMs7Z8gr9Qav7iI/ZaU+FyqkaLfBqU4h4n79L0gBW1GiUsW9D7FNPerT
NyJZurz21lO4rwFGqSNbzYiOCBloo6cZNtUjLL6CGssvqnjikBsu/ZyOIXPINkzpD5CGhTl/5av/
T6Nz0N0+6LQ6i0MzdQdD7EZaTGKr2JBDx6dbl95xiq2aA72yw6g5SMgU8NFGgfQgqETCfv+iBSa7
ExtBZrz5WP2sdmFgPC20tDhb8MBqTL0FBMLMqPGpNwCG/VvaqqTj/SmcJGptgPMlFN+/d2lnFgmC
kfK+6Pyaof06QbtP8RaJglXQFta45o80/Bv9bINpO+ttvvz/ZeKLHH3SBj71qPDsdPUKmr37+t54
jSpq0MpxOBEtIMZRui/kwVq/4JFlpPPHV8oVLTwmPwV/KcraQGpcs6C4RM+Im0eCz+9WQzhJaKtL
NnTsG/SLTWT2qfdid94e5et4QMQOeWX65jnajRv23ug5aP/D9ItUVDbM1TPyKKp51fDLWywtJ+fx
8abSThYi2QOuv0MkK6WQedqLPqZhPH0HjhiOUkQVz+KuVQsFuV6Iqf68RyDDgOQ82KBtQ4n0Y4oE
l/W/RMM7lz1YlLBkmlzZFwgPg1EAKyPhYfVTVVBINJjY7FZ9A6ikOWLCCSZB6DosFYElWn46XWT7
QSgoYafMpgBrmZcyZ06GI3BAzqk1szyxNK2iAVPalV60kvW56R22pxd9nnun4nJf1QkxVHESupMt
erHIPxHjy37eULsUd4Wd4OtNoVpSOELm2N4RmL93mKfH9HFntKfPG9bRzvP88i9xmWZr94YCvmIQ
5QZGQhtubWwGYRPwvArGR/kilXGsdrlvOSZlfPcSYArzm3VnUqzvtwJFVDJgYBJJFKwI7M+ktMKK
O3JCnlkpPtu7og+c+XHOF2ENEQ9/o7lEKeSBqK5FHcSgJ/JMFPPClXl5b+Rm+AyFfdzLQhVCwpNp
YV8lVGR2cAZXg2qTIuvs/FeCayydjuv9Vs5kFSPL727fLlqvB8aVF2ktylxWZoUTMdB+LUcaR8fC
Y++RlXs4Rs17xO9Ia0X2dcDWB9lQIMdeYXSM8oQx0lGJ4sTYLGGyv7uMNCrBGw7TG7DyhnJpNEce
tl7GDxTK+1O5ito/yKQqz1QK9V6tVRL2GrfgX25s5H1N4z39yW2cE6wY3wLzVLwSB9O7XiWhaD29
phHci1ZKY5vw0fI93V918Ctqu7VlllvY7A2WlMq1NI5lnzw/K2WE5OCqpkgBmtSoAlvW0Bbj+i0q
p2Qj9F0MJROEHtcxW4aTCDgYM7iEdyE5+wZugRYGnBx2ldG7ALNpsLzSkOus3qdkm6y4O59Aw8F3
9IgMti08Nt6+IZXbxqPItWHk/Fvgo5B7fWFNNVR59Lg6HB/UigWGnDkwIGOrEMIm3iTvvODYimWV
utAIEjH56tQuHhR0xnOnj+99mbpIMqY48kXL/z+/LSY4JdhU04FEwJKp6q2yWlp5EBrNrVSWAMbQ
EUhQlplZNQotKDIV/XzTVwdDB/zZaMAMVl1vCYFU7/LmPNgn18y+aYjPeFtYHhZbeZ1oLYMQNvtn
YY1el8y/hoghvh7TS5W+bQ90Q6dql7euQ7q4FK8NWAA1VA0SxuYrypo+Fs5NH39+BBxf0Qvp41Eq
R93nuYAiBz3rAjEAMM3iZ8QVQpuSx63C2fO8a3EZYtWyedrEj1sABTrHtDNtEkY2J+1haA4GOxws
TRYXj2HudaNq8EpWm0Hh59I+SdhXkUQzejeDrge5y8Aoi3/1tjf8BtAA8m+B8sO9hGPszFr1mKAs
r9xGg/asH/ezbDHOeNdEfqG8USLwUQ1hVrWAxlPtJt4E++7wTTFTzL6m4eQdQKXdmlILRZHXfrHz
0c7sGunNDHoauNXGgcoW8IeaQuOwtfVaGBFtNMvlflpY9FwntraWwO4ngFYGUj56AIt+WSG6BOXZ
pMc56GTeqXjKiDM27aClWAXT3/CenZF33qtck4bNkVLiLJuPnZf6W4m5DkMmlhS0/TZTzMto+ZH9
7AJO6Fp4kqdkjg+oH7vXcPE58LRir2jaQtKnmHbe5VqBJ3exYOWLjp4mQahel3fvFEoFIIVNV+Uj
DSmf0/31cgCat9Iz9BqvgZx9xB0LNXp+TGmMvvZh8fx626xe+BF6oM19CX6ckx+vFDo3WFxsnNhV
iK29KTtguAXxOsDqmr8tqAaXzMYN10k2QWR62+JDmtIfAZAI+vtPjToFLOBFiDUyO30zESz4Rt3l
GJFic1xvOgodgXBYNfKShIDxP8zNLF7ViHUHaDmPLx58kZhJ+o/aPE/FRjyAqn7+rIYmQOQuJM5S
9ioiA9Pk/l68ZedHE0zN6aVbYXJzGjCSd3Vux/OwxgcwEfnjnxmgQFe5L3YUFfwoS9CRSsasK8OW
0U1ymHMwkGcaOSf6bdAcZvbd3n0o/kWdpU4ot/C2uM4aZ1MniVD3+yjc820lXfZ5Ubd0CfRvN+Qz
pBdovVqybEdmE45oMhiiL9Oaww4VB+B9uTYfQV/LG9d3zdU3oNdZH7EuMJa0dYYP7tNna2h2E7mi
W69DOoabOqBPwiAPmLTRCRuBra5AJxLb6p3s/3qyJe5izFV1KnirCsiRIihPlfctwEXfXyIzmn80
UfaeJXvGxwLJYr0iIsdAuagjQUPj7Yqqgvx0qLO67VokT8rQyWcXpG/1WXdhmDNe7N/rELcjCi08
mYLVybh100WkzKEcnDLhFons4ilexNCMvq/LaWy2E88ZuwlSXlnRek81bS2ffvNCYrnATdty3z3t
kieaY20B+2rVPsFbHRZ9nYj4C7e4LXU9E/0SJrS72mQBX3wQceuI/LhbefSeXT4KEyakHbkWX59r
rIcKF5Wlk9a+HoDx9drcDLFiX4UhU4eRnEXjI8mAs2sEmCY26McGvv+7kdOdc6fOMIDHfdK2QPBl
leX42NSzoLL4QnBt/WWCE3+7m2PqVrUN6ObxMNCkEpFR4HNAVIvzQQrXQgOxR2JntWC2pKyVYCfz
FffEale29bTmvYaQbhUYhqiWgnieiXJOHEGaEPgnOr9155/fDABamU+710XGPrKn9+sYT9oLC8Sx
j76+sRsZ4C/ad5+rALGVlC1sN/u4FK0AI/4K1vLoUmYSkkXfx8H36KwaBYLQUJAFJO5qqoEJfqvm
RSVrZcRduhWoWFGgmqd00sizaBTlThA7elOahEKgRHKFGSMtP530g80GcUdpj3jx62lCSv1m6T86
v+eRw/SiHK3bQ9Y2fXiFDO24MDL2RCqYlIzdjw7mpydbneefllYEOOad40C031duJ8/VZWz5mObv
wQL6eKC2u/unmAce7G1bY+v+HcMzM6CaX3CuWITKOSy2lDnLeYuq6Z/MzD5Nf8J6+Fr2HkOhfIJX
PnGHmFgUyhLu1TqSKnGLXu4RcDXWYMo2MC5aL+QGFy4XlaA2xbJGWhCJL2g1uttlsvDxNaPf6Y5x
pKBVt6jEEjCuvw0pVXVtbWL5PH8UT5ZUv4x3XA2hbfxmMb/uErxZIhrSJYP1VA/fuVeQw3Ch8Wui
GdJ9B0cIt3niEUhVRUygODDlSt8nxH0+2rqNQ1SA5KtMmEMD3J9olUIjFW5kwqI0GJFt+eveXfuj
m7Qm/Xs1AWUhpL+RrFfNUlXMZoBiUROt0McLcO0Cv+aof7ww+9C1VmW+jWulqmsfls0nwGGpk7fB
TaNOas+EJFRdy8ULQiKXYAunCK4KK4cZYuSFmbwDp2V0MCOIIdxYz5VWgd7aVOTy+z4HWQgX7Hb1
N3ZEpnEe8jhFIRLzMPQzPcWN36n5SMkhGAnr80nsKYvp3SHYfHg6hLZe29URL5X7wY6FaX3rdx0k
A3Z3t8op8l3LFdEJH9xN49qnUIImHuEPGfdsmCMxkknV0csL3tKXGNXFbhwRc0tT8aalOWi2H2G3
UMzyX9lD1KVpH1X2wvZQ0RsIyLPrUYfjzXYPFj9w+2R/W/DHXS8rVl4Hz31zYLylr4Yym9Fyh6m/
SFA1jGqmOoMZgdR4U6WoaJKhd3lBF0HgtcJLtCTdK9RDLbOsG5yfos8qqVxapxQmyeBpjJaVKhNV
dqyTaf3Qb5wDfCJlsgWTVG4ZjPGzcb5pOWyn3B07NJQxukiYtx9t6vqXYqvoH7TP0jATSmuM91iI
RxmYUsgNQL21sKabfbdwkoZ93j11sStqLbx96SJYfbipAXBY0sFYblgniscbqbWPc6HLEsYWUUzV
Of+hFISenmKVr1M9xTKAGn9xYCZn1vf33Ry44UHrEBLmPUlfvY5zf47kttgKltVm1i5e89mEIFnJ
D4GsQt2lOf+9PA4vIINhDpnSrc6PEXmIXUl52He68dyvKsqo1n6tukFiMIXawXWYPc5Ib437eE1p
7qaekia2EERVsSfWsrslchC3emlstJkR6NrJDejK/nVZx21IIlCe8gLwF1Z0L8JF0hvzPFDFc0ZK
jCmBJOr0KKE7AcHcigoNBUUWkWbgbHTt3gGfpoUALlR/tQrmRkfR46GtlKelPgex+lV2FnipXPtM
k0Qp4Vm3Wdbej72V1ZpIvKmvbr/hrX3OrYVsOOrGDuj4xzULqWX9kg88cjXTGHn0iLkJ5jEKLMWQ
UhDVDq8ni91q2Fzq6mO562NIViAW3cw/c0WIHV0L8GOdVDbCQ1SkwvFhRWOsUVacqkaUqHfo0177
I5H/M75/NIPVnWqHSl7htlPSMldqOfyRlY35DLhOMi1MyJhrMSSvjtf3XarkyqFZau+mgA0XPZXy
CcWw30W30i33OMNx0YMsVRQYv7f8wIm4b8QUwLiS6PmjAqUkRtBN79QEZUu5ikKzwC8kSWDnzi2J
rLjasKm01GpJPQW2ZD67Py7YMmI6xP4h7PDLGC+lOLSKzHtExl4VukEV/bpiva4TnlOhMvdkFYTE
s7taB4JMo2q+Mt/6v/IIYO7AY9it5sW5qajORn1hcJjFn/m/SJ44edXQkM/0gkGvNE6c3J9+sLH5
QP/yBnTaorkFe9i70DSjfVcfTTz3G7T9bFlonN6gXCWgVQCYfpuNGtQpATu903ZAh8uD71y5xcaO
mN7+7CgDSSAWjhvkZwAWr3dsLIMAcuXCSVUmNzo5ZdiLvtgobcXKXth+jmCkITUIEZdoTslBqOH+
9ZAwUR4E3nwGjwkaUR6HkfBLLaBcvLh1q+EivSMF7BWf2BtS/i60pQ/Li8lARdvqaNyPY60/Jopv
XYfOMGXxShtJs68t2JgnvGmlPdCU5vDQGIF75tibtf21MK2CxIEBVG/DKsmt0QzLv5dJ2tUTpPKV
+/pDgWLgdanZ0hw7nYZRyYhfmHeI16yTpzb2Dn1d8Yoc310RlA6bhlje4e0zE9H/oI3CGpnetFkR
elt8PphsvO/pX7odQxNPhUG2Uo76HEtqJkBg3+2GX3mT2xSNKKFmU5Twmi5Teb7b+4K2NRmZCL+j
PGcJCLOy3g/555SJf4g8rmD281N+jZcakP6pqNQBqguorQOF82EiPJla639u3t9FrGTZ9bp+GFaO
Tdk2EK4+nVcOwkEjfcnCbgHv+KoRgxUzksDoyUn7wfGm2s5WMGBBXIr8CHJ/2kZ0DSG7s1cf8E8V
Xxf4W+JteATcaSSVt8iWjIVD3L3CtUSha9UwHTtQEpkhixEz4ktg0pZb/JjdtwwpVhVUokq1JlZn
3nDj3CT7yyYrbTmseiXw2RolioU5BR83/gJVFzkwMKZb2Om+RPYV2gckC8dAvchagZgsKvNvaEV1
ITMzO9e410F48Sq6GpOyG8O4w5olJ+jg3PYEqDgHJaQFZX8h8LtpN9oR1fgu68bDXYgoR5e8nOTE
uKKK782ascQudf7Ur1zLTigzgUWxxjs7RSyYJDLDrMSyW7KwMYsHoIOmtcNAfF3YSMfNgweqeyKD
x/fDgU3S92pLq0/HV/mnqmjtPlR+0OshebQtZ6VrxYYKNGZ/A7WrfP0r7kwAV9i2wmO5nXkqN396
5Z/u/aGMdrDYj6LiluWHTmQQy2xk5AQb1+5Can8bZlHP+JEFEeY9po/jTLy7MJKDTtIw9RXAaZC6
Yied5f3nkO5WgMh00/8r40+3cB0fkSzZmFU34zoBj93aXppd4F53jFNJAFyfXSsZVC6no3lSqkFy
d7Vv+++vhbpHrf/Df3rUr8fDHecAgwL+6LKPL5sI02iDolfCHl/zmmuzpyIGuJ69hNERN0IXGcZY
oH6VyOHhUCni5e3vvP37o7iunajpEVgMu80jd/oVlKeDknrI8B5/03EZW7msY6RWQYL4Id3UUi7L
l/eCGWDQry+jqSMXVq6Pm1eQo/HEWQVeft+Q7XKFeOV6EA557JD/CLnwV37vtbmDQasUCzMaXsCP
mXxvpL9LqQO+56s/cPDCTLaAMFwOmMzCfGm4BcFOKbpFZPzSSF3JEzX1SWE7X727lOA/TaZizmhl
hqbzujZpOYHVONOcC73Djh9BxSYj0ynELCxNCHZJa17VB0gtgoZlHmffl8PI2pSIzswtHPVIWOEp
m9kmh/+5C0Le9bTgXI3rJw4/I5MgLvgyjGcbn6GhaPJK86zjBHHB0OFklcXIQH29B18qxUb2HcGM
55G9HtFJFpzm0+9aGS7OiYyVpFkBytAD2zKHPrc1tgOteNaAMbEX3AU00b2p6yyQT2qM8jXinDvR
MKsZIycNrb7gu91A1y2ZGRP2BYfnYZUqJCqAMcmCNyGpC7dF2v5ODLzjO+vDSkjsVsqpjejCAKUy
LTpADsHncCoxnKxdW0lz6KuyOOSdl+cnd8VYZ/WDuPHIB5mUFf3Q2421jEnPpHxdpntjtE401k9A
C6l9gH+RUmlsym5AmfaZDYsCLsdYw1fGceLomz+j4GzcwXNhP1V8p7CReQKruDayB4OpoUjpneyo
OlldOCBwQfsg53egswDusTeCshY8+rt1qU2DCjrMW5PK7IF8xw4ifDnFglVyEk2jlPy/t4cQTPRv
wiPYc89eSGcxqpwtW+f7fPu1Em2K7dhnX+ZI0XuXUaDHa6Dw+LFHb16H9rWjOJPgFWDdJDUFVes6
vQhYzc0XTeuJ9B0UqdokHg7pulxoqoWgc98hKSbPvSWTUCrpnpNFK8uBMu4LHfjI8hJ0PKw4zqAK
7CQ5zhf94hGNC/3mbuKtmmoc7z/R8SNdICbIO/zjip9rHrFPw+/o+HNZmZ159sw8IzJOJ4+oCOzh
A7c5s8ZNLUh5NJI7So1R6gSUyYTtGVXD0CZsfZ0gW8mYSv9qZw7wGpXoRNLmg5bYauAfRUhUa0tR
xviCwSmWGgmLLmdPMTz7QtjnJOcdZ4kh38rvX6K3SahXs22H187blM8V3tcfu9KScDR1siJs252B
aCRkg0+Ch2RCrw1BY2Cx8Hl0EDjrsHtfn0Tu5ixWkL85uuQpOkb9Qzr9oGr/DgvsfppQB0ShRm+D
w5VdT9rtBcnO3c+SHLDM4EVUliw/YtrYtQ1X5TqX1wupWF6PoBhz5y99ECcJPXMAJFAq2dUwbO+E
kerkCrA5PY5D0hLB4Qh6wJ/o1lU03xB7ZKHNDI4YFCJV9yi80GoEAk4SJ2pxd4Xmkp+M17F5LJ+T
uqqFJUMkc8pxMjFY83P09h3A7dovunW1NzIl5fxPyyPcVYD8Y9qKbv6T2gp2CuKwx3o2s1doP+ut
AJ9MBs0qh+TUnf+W+ya/LhHU1LUfihaQSM5Sj1VdQCZQGsrtEVdq2mVyCuk8//fSXAtBahyqmkub
MpktRxq4oHvW/TCfWPaJ5KIHz8cQ71VLow6Dq+kPAp+XvY8L+DeW0D25mX8G0glMqSGYoCh5yP0b
Ng+jxlAfAzefAPzn+2CAV2CIoSw0Nycm0ufQ7WHD0kADKmMOnRpp4AkuYj0sMjShyEIjr8zw1XlA
+mCYUcpIQEMafN11efLinCpUcdb+/PyiupMPQ9OQf537hjYui+65R+juPL5yxSUvEdfIXNeIy8/z
6QlMZN2rYRQguJFTk02Xyz31PifpWXChR54c3rcYxbUbdC6N8hxEJQtKgeEBGHUH1ftS4+KOZdTr
3BK7wqz/OH28ZYQwqdudb8dBhW1bcvfBuYWFSKs3j2/WACRT7CuVgZS6qwcUcqbX42JhKcCWCV6V
esYPXhiAOwm7rDv/WgJyMARZjGMefujY8c1FU/DOOVbHrJKNDc5lQTm9k5yPjHzYdPl0pr3yHK3k
R9mt6e/4xe1p27RORKRDqU4S1Zgrazew8PBmQz1pLuLFdxwA9tkdT00VxjGfQrxJyr044UZlDiUO
+imXPCWzTSGjl7qM/NxWa/oOUm7D8EoL72odTE6PuTNcRofO3QvT1yZL4eWFiMNeavDv2zEWNjVb
Dov+I4/n1V1RHOINV2wcHObj0O5AWcwrDUcrkOpT2V6zVlsVFxSpT5i5NBT/nYQLAK9JERYKqT9A
oL7uU8/WQvpH+BuIUWKEaHDsP+qNj7DAMgAoN8DZZYl9hHZbXlx+pqwrixTw8SO29ssjawtboquM
ykQlgofZ0AjbW74LUGznqHhIzRYj3bNBJH65DMMWsOw/0D/Hoi3b9jJuKPgWQKy5pB4A/yJTgNSh
JpPVe+Oy1YRxyxPf5RME/PQ6etVwYRb9xjqoEBFCiFOzcgBczM0Ww7fnNTuQmW1+v8aqYkJoGTxD
iWIRShfgiCARbKPmWg8PXQ3hjrFdjB/jCYO886Vfo8/qRWW9ARP8rentE+nrg+DV99Dp+JbVu6De
2WvOBm93H8FI+QCpdxCArnaZGGutsPzwLSgOgQxRe2XNz7ouS9FLvU2iliSluQccfRPrW4UxxW9n
5/oPAWSZWqXE9p7iBEx+DM0AVbearCivDa8TeBoNUztiMCu2YKYNY1c+TdKIXWviyOzp+SaL0X1g
2pgWK6pUVm3iSDVUvolDleg6m/ZNJotyh7bn9gCxjVrQqQyiQfxaSq2MQrXtEQ1PMczt/G5YbH2G
vSn9Jpao29NBLqkfNQ+D9ULU1Lfn1TrlqWHKemXa3JxOu8NSlS1VMoEupvyc9yMzUxT7yfYPnOA+
O8l7K0tSgjcjJneSgPlzSjMr7DlErwQgksHbo9WVOf8z0Z+f2/dY/w4KxNHifSnjFkzslbbhHwiL
NkCCqRwNjdeZwuiylJAbnwmIcOcQiSydyAHXxzG8L7gE/dyzCbDG0X5OhERurOBG5SjkcaK4hWX0
QRBDIPzB8sPMI9m5tJ95Y1p/yp4/WKPymzZopoBCK4oQ6LAdyR9vKh+92wO77TGA6T/ZfDK5V7Vr
tlkkVRKcvmJF3YkGSmv7PLajMIQ8cuHBjZQlom3rMcGhK7SkC100EsHqNwRysedw50YVwkTw2uHB
ZjTSZLgy2Byspk1xHJ45nkeGkL2DfG6p2gZPkOutGeaFZbybisJB79R/sYDa/aSGNOGYdXLuXTJI
poDK45zVZ2IYSBbjwflBfVNkMPAt7bkr5nK5BkkkcXffMZTulh2JWct0i8/8Ci3E7aAv9zJrtRCC
A9GbBzmpSS5Ly+CVdZSaaMwpncGGCHXBYDU8AWCm2G95Ypyio+vruNatBcGMXQ+H1eSZCCE1Aa7z
05pwkP39OsyYUBxrl7OWEMREM0OGUlN8idILRQ8np37voATEokpgn20tScKFkcrCpT2vHsVoVuYb
GiLiRNiKbceV0sAx5DIIJgfapBxnypjBeqi90qXm/Hdh0HMzHbiA2dOYWeB7eVqquS9MyjUby9b/
XINzAXBnYhzYx6x4Up2kI6GDGwqmxxHfKQAPKHeUyeSj+UgQ1C+4glA9yqyu8kSLB99AZHyMLj+4
CtlQ5DyIAYmOaiF/153svrUxgEtSaSAqAr/SCH4eV1Vpdu/YPnfVgjk2E29j3jYZe4iSE3ZcCb+i
AhhBCNTtKnz8y5XyxmRduDEOs45eTv9EEte1uRT+JZo4OyQ70J6M3Fu/b2ykm9nOMITQttF4ekbg
8ZCk2fyaOO5JUWH78RPZm4gpMjFTXTTl/HS1EXkm51uDRUVW8KAAqyvG+01F2RsdDWEjfmX37zYZ
99Nkkm0/vv/20dIrQmKtzJlUP/sNkL3FN9eRlcutvsUJfJIFHqPS8TIZiEgCZoXhgRi2CvCBv1xV
OYVKbKf3yVHl4emk1GJEjaofrkzDcuoVjYY/8k5jhh2+DgA+HOsahCeFYuBspOmG8x32g2kK6//R
JiUUqOQQedQpjxCvLAJZ2Ghf3zac5wf04+QI5XuykNlA6yVXN5jM3QmMsD3ts0ymLSlJeu5Jnv//
13D2+XwO5n0DmuJVIMaOWNJ3MySvlpQoGN+jYgknURpe6WcjhzfYvP/JEOzlfg5071WnJf2ZJm8y
RG8I30s+ZUw8VYkATjBk3PWcug1zzUTgvc/hC5hrT/HyR1SDv4voJiFdt1QSK0lId36Jc4xbwbee
6i9K48l/h5WLgPlwpKMMfWbLDWPJwDRl/UnUbDvbUXeQz7FspsgKoEim5HPKtCrYW5hPSF41MTHU
F0hL41vKM0TLEk0oEdymwGHluSrjG2o4tRolcpxobjH5rwaaaLhg4TduVxKLd41Dubikl5btU8bd
GKixlsC7oxazWhJvLbcgR/11J/G2vBE0i57EvFy0jp7GDnuZnkLOrd4tpJmMKNtfQrzQ6pZgSVMR
jgLOdezXVabsfUn2I53Yhg8idh8kdE/9f99v9OecVztuHLuwjG46Z+W7WbIHGDy2qmst9ndtP92t
Ay+1FTvcWB0Cai4ZFi9ARbwq8PsYrf1Xu1P67JqsXcNa+/tB62ookHFPx6kR7wACuW9+IPRQ69V+
Dl7uvNEAcg5yuwTwhXl/irPNxrHhENm9ZQoFueIY47Hb4z11RYZmRWly1E79FeYqm3MgTzEV6C1k
z2Or3mLntvZ5o29D3q7WCEMz49FRg9h0NtXA9BiACFYwVSTeijRXDDo5P71vWJKrBSeqiSqxGZsT
oePFl32E0bUptn08M/6YLXd+TnxmBHHqwisBLrUSqoDe9yyvfRRg9ir3bR1j7Ds/ZhsBnx7MNGyh
908r3YE1C4nx/J248uyIBHYqgxZWEo3bxixdVuz7B5VndtTg+Z4akRgIbvNyL4w/Tkv6BJDmQKIh
drOKNw4gfMpb6cQkkmn1CDxFSmjwm02U9gQ3BDxwEYzNjbtYWwoEtEbt7K9r3/40CgQG+xzPMUoj
HJqC5321nbNBg2mIZVZ616DuqRe+mamWDNkufQZ01AGL6p7/wFX/BvRMC+OgkV7gAV/7RKa41eKh
NAeLGoqkMqmRc3tw44jHJJUXyRiswNO3JcXpvjgKd+nnTO/e0nDEFj/XpPtfiAPf0F0PY12qI0il
/L3Cdbr8+Nx5O+Wh9EcUFvSu9FvoBrxtlso1QWBgbBhBMSYKWSR+GlE3VXs06Lx3yjcRpPtWhIt1
47U5Ztl2oEJvXB83q/JibZ0+Lo5OP7ro6Hl5m4p7RWP5A3rsXAkSZMudakjibOt1bb9lVlhMkKA3
064GoSQOmmeySsNSspao/xQ7UBek435ojh9inetRbjxtF2B7icTyLWOs4dG6aozYOgrcOe2J/9RI
cp57PZlX3wQu+OCuTrCVXGmwNuAcsrAUgPU5r1az9bK4B5vEJpD3w+DXLbyZSSYyEvvm3F9FXr/c
c+mlSB4D+h4ktsrzKshqOa395BPbqUnEGcQPXq7EMnkiLms9VFsnVYjNNs/si/E0MdJP0VsWhdcg
2UiK9CLlq9NQ9pfm87MZHDgukdSRif7T1jilQMcBTDWbcs4KcDNYr6KdmAu17vTUYaZF+PUoJ5j3
ZQjpVjnVDfM4Jw1lX3Mm1BiTDtAgZ3ehR9fTicrAea49eEImT9UdwG0TggGsK4Xlg8+sSODwrvZ2
UJcTCZLR//nmpEj6wbrnCpaRYlM2X6HABLk8o1SMxXEuyd/IP3cjWMo14nLB4mxH9YNmJOSoRI0Y
qqznK8r3ipVI6P+plksaU8ysg/MgFacx2E5r/nkzW5q58XczThlB+kTTFXisdbRt5OAcYstzOiEv
uUE7nlC1AR0QnOWw2KCY+zzTcduBfdxJJ3hUjES3nSTzf5Iz6zPRqZJSsA0Ul47tjpqlWWhyp0qf
gtmHR28RuQJu1DFwSUuBvh7DKm1wUHRbkNbY9fpfl8YReaXrGOd5xExQ628/tZHZJhmBmJRmAzHG
jBs2CbzjSlqwX+iWLN337pxjTGb7JMRBxFjvsoRB5i9fRp6ikNjA7dem6mN65K8IHrQ1g6D4GMc0
0ZCt8PIJLaoNSNjn0Fa1hZsojodY2GxSi8Qf6tMqdSgJKpeW5rDWIfBU9JZLsMGS093A+W3qbRBt
pm1T08x3OI2BnyJ2m8i9tQNWiCdVXP455yusgXaf//pMrvBSMRQkPPkDKu2sSZF85Yy138DQvimR
d+dMSCLKbytdHlNeiXE6GyKEgepYxsq+MNVToz57aRBOwlA/X07Rr/5AcwzOKVowsnKF3qEaLd+0
cHSek4sNUdE9SCOH7h98vvCmuGwcdNyHU+6/sWThPd4fyGJ/8MMfAzJjNfTSJcYapxRf2m2AbFOy
GQoYH0Fm7XN0rbCRcJdMRNqYhM/KKvGyuzQdNbmGGTyF+MTwhH/qX+sE2rAg66K+F8GHbkZsIKSZ
Jwr8UWDT9wvemGZMFJWm6VVYWkpk3/9xufuYV5LsLGZFpF5GU3K4dnRRYfi1/sWg/AD7zUlqfcPJ
4zOJhVhBIlHRZi6K1SulFHd0dsg0eZFi9ILYmyzjcUKcGo3pyc0E3bFgEvksH4R8rkzb7J+CwZgX
J0zDuNr0mqfCBhaARMBfUU5xQQCv2s+fvf4JzXcTH8fBH3SQh2HlomkjYZy3CytDToXN1Ube5LAw
TN5VHiAbrMilbh2GIeFIcRtLfaurivdf670DwDDJvpeYDSfO7hh6fpBHhAVBBeJO4stPRJNhlYDr
T4uSUQs5gizri4oUhPYXqkbRNfOqsD3KPhRsX/i1XWAEsXW7FFZ2TQbNSTKxPtxC0BQvrjR6Wqth
IqtY/UB48MlGnBXf/GqsNL8TJs39hboX34OTeQmHu6ywacagvP/d47C7iPI3RRD4tmgKHvYxNRRI
hUzxpTlTkCVwxvFqX83rGiJAa+HKKnGKk7DAK8FOgHtxm17p9xgTnaIRsWiRhuRLr6Q+KiKxULj9
EJ3HwOFdASuNXFjOX15XeHBKGFHFtPKixsViA61n41rysMSYE65lICcpiiP0qcyxhM9nnGS1ZozL
8hS7Ta5+e7YCE+G9bZFlZGmEVq6W9W8bbkTPlMdVO15HA9NDYOORTuoX8AYGrTi8x86f0srjlrtp
vn10f+bHens5yLjhPua2ybSr5y3KKzmvxmjBUZHUadDb8H90gIQXp19/LhMfseJ46CeMH8AvBzun
BOQlalAHuTxlW2M6xKpV1Ss08OORfavIxJsXB/K32SlN/xTRWXlWCHU+tT/t5/3QDZLbsC/8LVTf
+HMQTkONeN+laICrbVWfBGRzQanFsuuYwmHe2N3Il8W7pO0LaqcCi8KsDkQheqNxZfpKK6vAQ2Hr
brlHEuQMWLwxsf3XSTvqM/5t7/bmL6NN2xEhfTGPg1INIcyEn6jGyUiqm09LrPSkQxgeDCY0G1mQ
DkU3qzBlUAiZKx0mU20QLiTIVs0LrKMxx800EfB8C6gIRsTqmbXm+zu+eA+4TYg/NjXKYmXtykL3
K7WF0LP91ICfU7oDs1yhg/FhNXMCjJkzlDzxHvqkQSUOl+welu8XdvXqza2Bsem/mpvOBBUD3zlr
cfAJRH5un75Ah/m1n7Okaz9x14kjV6zdq2pGQwTGcFYYjom/tvmnPIYbNMuuHxMD/9ho0e/y+ihX
cbZMDN6eaDoM1+aaYtFWR5WITakRPvVVrdKmTyVITbZU44tM/2T7MBIIKSqNI+gQnlOxZLA7GJ14
WEFx9kRmkuPMfHbdqcnhyll09RpddlR23e0GcNtmzLb7WXxFCkwdjRuhjKOmqlArhE48b9WswSqc
gf+yzw7wzQjsZkFBh+cYvLHNgQvcxq7es5MuFleVR/6eVbEsnJXkcwPIFp5SrWN5HjPeWVG4ppO1
EsdELpfKIj9owURVWlxntYVGhAV6P74Nc7Xd0WafzwggwlSQh58kSMSU7zCakcea+cdQQrOl0SGM
hKJQuSs84bY0Rh0kHRLVu4Yjg+JvC1Uf2BpQ6Ozfe7nTCGThtFNgT3sX+Bn7av2CvjuPUHySotp0
VbXqYT6xkm/Igf9mXAVL+bdhWhc0Rz5DcmDqQ7wyZODkrSYaS8fmjMHdAZdaOpfDm6VxJaFd58AA
sbPI1vZQsQbANMSozZ3+06v7VUUl9iAJnCrwydMTqbmt9vEzH3+VgrNa3S1DREyqr1pJIO36zFm1
OqfO7uOZogrb/Xa452w5I6j0kGP9awglTd9B5+BOKhofNCRsJWpsX3onhRrm7guTHdx8E8XNY25j
l/13eWYyuKxqaLJgouxlJK92J/gRnZlwib3irHSx4YmuJ8qf03bQbgVVxxTTj/Kc2rB4/2EHTYv0
rwNaY1P2mkKIsWQLmsBAzhCNiu6gFhgzEYxyabs0fWb4OgRah4LYFEl78ILptohQ+Iep2WwxZ9TJ
77KjK8ddrbgGE8pP7xytdzrgxivS76QccgvxnDlUlG8Hwlx7HXQI0wcokpXCcsYA+k8C3JA9VkZV
7T+8laDPk0dbXnuDfU/QLHrrwP3rBScJvA1+7IbplNi/VQjJhs4kf/ERA3Uz6bLeUl50SniT8+Pc
TqYFvf1zbOcMamGxUQvvhK+kIcWFpdjSrWHG0P4Xpzhm2pmVyphjKtZ4cjUaXQFKlVJARbQ8TqJr
80lIdkgelijQtsAMKejBS0NhPrr1jPmgczAtrP0Wckq6UbgSVjiCjx7sVH6Ix4ZKHpcvIdU0Hvn5
GgSh0ginlvQbr3kilPxeLntJw5yjnDeKqF2YK+bCEzGs38qsSvY+wl60oN4dbP+Jwpkf8NgWX+4Y
jeVtGPEEbsGAKaekHIlkXm8oJqdvR9PoFr1uibdqHKNIv5lcJYtuH9kmnlJJUlq11mDFL20ywvx5
SFC7izC+7noGGn4cZ8b+y8bjhQ8VT10cHJ4NgGFKJ1piAZ+Hp1KdLR0RczZZ3VE1Ct9AMmxhIQkf
9HfhURxG+5DePWcV5V4Kc/6CecTymBs9cH1gZKrFCeUgQ6WsPkY8VgtI1MGs5apcmuGf3vdFeHY3
gemb3nD+CO3wfaZ9CYfS7pEk4zcGPhPVJDWDNP1P6Gw3r+n+yOdzfA5YADPh50DJuEBCPBx6oIme
oL7A9FUDFQLGAp7LeITGdqEC3VqIw2pcX85x5cqLBT51R5DyLhgGUqQ0sjj2oUXFXEj0phassHtF
X0CtvWBpGYVnAezIpbwnqIpDoTZ2hE9VtnL0mEjZnukzf3V2DzB9tNGGdZtJIKjrhHaRv4fuuk8n
tBU+RX8hzJRpzZsXigzQRLGkCsLH7nQ+TKDyGjf93XtJzklRSWCNHgiQlbIG+feEcYXfaH7Pdkdh
6UPFQxagYo0yuidgodUWUpBxHftglexgrApjb64bgdtfIrHWPTfsmJ2nSt5lEKAvxrhqlmO9s74z
D0TJvHTb0VMI1hP2wHdxpGUbPXYAntGMc4l/qP8yY0h4tTJGy87fR4WvJHyqD9CTmH2njgggh/Ru
q3vTjCLFmxxRYg844jcynZ1sdGAaotaz4loajqBjjiACcQE+3l7kbNLj5zVlJibX2qiKSgUEKnp+
8xbOmOlUcUFc2Gxo+lKEOWwl+6fxAa6IE0EhPSN94iGXoFZGD0iRPvkq6CAPKNTmreUNoBil7YGm
kXcV3kiufQkPmjvqaQUzP0DR2+ENzZxsdHJZ0+ZjG7MIi3MJ4qalgllCi6TQ9mc6J6GIKhM3I7tw
J3gTfO2Sbrnklzk+XEHwJaN6UQf6o+j98Q0q0dv9N3arNy5DIO1ypcjYEwYRZveKd3EnFQyA+ynN
AC7z/NV22wtqW+wJF10AoV4xU9ClEBAQLKp5GZ7t/wHg/prOh24IiWpwWdtTqg5/nU5yjWrF33X3
HV6AphBTBbq/Xgcyqm4dcQcTbBkJL758K+mhv3yPQNpLw1nAbRG5SYTcrvpI5nGoABKZxQJDqj54
OobnwQYX2jgM/4CGn2NSD9jsWteMBw9Bs9bd/Mutv46GRKsC8OdYas1NLWbyu7lVvCpOmbpd9YQv
5eCwKFoCJO/TyOcRkLF/LmiSKgGdBVwNwXaZjKIH3IUkaKypfvw4k1kq1dDcWIBn2x/rL+PSezCy
MYbB8YU1vYI8bxD2y9cpRTFqF2yoYoU2VYT1vCnICuON8FqUgyJsuwjpnZUpC1YHZHi1o2TVTGPc
SiMsdgquTo6LPreHWMLXPTd8OvpSvzcX00tVVUShurjzrtvDxZzrCXxDWhwXAY2c6iOcQNb4F25m
qbQ3fW9B8exB2OhYKIEI3DlnQZRBTLPRjICgejIsvYaUS+Am30X1hzSp3HFMEtRO2AN4XEj312t/
a14vX0yC0a1ATSl3xYZMWg4joDYgJctJI9RnQWOmaSTb0SHlevIYS8i1KIp4IHVHjEP5aZuB8iLh
NP+sy3z7ymGQSQwLmmLZFrU3RhKpsCFVN57/PijCOxioVUvLT/C8sWxczAYi+OynqrUiN1/55kX/
yeWw7ooibigo7rtUbbMEXXbkROTvhfPK+PiKqpk6h1oemTB/gncQR+X2vJdva+5GuzzE5l5uk7AK
+2BVIOxOvpNjp9aq2uQiS9xnQlMGGgDJH6k5NadN1WB6BE/SEF4+BPVjPDZv7Z8s44Qhd2uqVreP
onDJcnNVHFKbLeTf9qQHOjGb8fLeFIDIKAtwTDkmsvahRvpVIbV2bNyyZQDaCepBgx6ExLVy8M0K
gBbRu7sIYrNnWUHiRElXtnq6U8y386ZfDU/Y+Y4MwbNfPKFcuLSTvvZjK9pMIoAp4kZLthta3nne
oX7tnK29I4vubH35UZOxggGz9wu6T/r/v/Zooa7deH0Hn8YDXLVWUKUo7APMb4bKKVb0LMswBvVX
LX4qpAhdVMFqDjgD/yxa6RkRs2opFAoxhsIx8xOkWjdYCMH88B1qmyUeIwc6T/SI7/EJ5NZjNmlI
IGroiIIwk8mmSpzUiWz0WKH/zsFShWDQzfsNZDvGbBeAIXRBee8hQW1f0AsPBwleVKDTtvvzTRdJ
N2pf5Qe0KCbUjR55c2PQqlxUaWPQtuXrSQhxXQjz0N8bw592k6RJnhkAlgIbxLkppaE19Ewf2wK7
8apfIlaz7mOrhpbHU5t1PbYcYmzL58DNqMOCMDPnxESx+XcDd/h7mqdRePUfte0M+qIlFDil+l2L
VWSlFDEsZvwkAXbSVdS49suWpJ9Ade/fdSgrL01vxKsuK5iIg+MnN94UYOCMQyC5smc3/WyD1OiU
M7f33lmPG8EsbCtxfGkYMIhynikQyU3+F0+BiECCqPmAREHM4LwUzuC+HQQoEMUMQ352pvkXpPW6
HnQ4qGCPCL4XPsjw2LltJRrKVNRih8piN5SMREfxp4EsvIyx7P5tYTaLu18ZTcS5t8wyq7JdZ4lM
WsZxton6YNhsGCxlfTjh83KSSa/gGdwIcyIol6MODnzYm9Xjl39EHKQze9OE9W6DMnaziQlqjLfR
VWvkL9robzT20TTwhcsrpptOrUogyWexBB+BGl+w2r4WvSW2s6eF3cX9/unbWTJbbcAtlT2dB2JX
aTyoxo7b8D2tdsg+23QVpEUgPzt9tmkjqWP19UE7DyJeZhjnkgCrbuWX7lcPu62Jst6SRvqvpv2k
QSNsn7dL/UHYwJZl81N7fjtmKdeqSKfE/fLveMiKCQOcKwh+3z6mMSQ57R0GHS2XI6yM3Ay1IP7E
0NzJNv/38nc7h/W0AwIu/YwAmt8zgdA6uB53K55JhYXjFzhqXRkU4LkoalfpjQO5N4Wo/Bl37DeN
Ho9X9rPsDsvriKXA3qM7uxXLSqJgwKKQ7FkOiRl4nNlYTfAQfyZXtGmsRWhIvMYwcg0+ATvVeU7y
KN29nnhnhn7E0jfR/K6dlu7+H9tU/nc3h0PuBqorZ51YiTlpYYT0CIhMCIighC6zBmxBaCCY+UL3
/qhvA7dBlAW/aoYRN/AfzlIZlN/rvEYWAiXsXfZUvdfpllHNPQLBWuiVgeCO4lMUa7aS2I9H2gPs
XkVSqH121iC8OHfCJmDvVq5DcuWsQI2WuDBuBXzXElsTHphPOQUahh+gIaAvPUkAQcFzqip40CzF
Yd+Ykx0IFpDZw2qajjX/UIwVSMjR7PnL27EZacKaU4+iVsT/cBsBKwx3NB+ieRepRfP9U0RrqUyR
IO7twQ9WOqwuSjvm3AyiI+tYdebQshk1CZBdq2us8dcm5f+usmA+VCEFJidBLbOrPorPNXzyrATT
MjINhFA4L8dT+UHsf1AYBzUWndiiu2NiKk8Bz/LEQdQCrdq0NM1u/NF6EbOocU+S50CI90dFsx8g
g3IxxccHEmL+rf81H8LUOI6uelQjslZJcMnhi/ww5RlfzNoIRuLJnPHwKm2KpiPL9ZY/W3niA2xK
x9YDByanzv2OxgYDFHfqVP5fHBXzpil9SPqDNGhOD3vIuVP5Q4yQGkfa1iaPKzzivZoqY3y5md6c
0tgCJKmT+lB64NIu8cZgMTQIT3KzhcTfoRjTFGIKXYha35bcHffCFyneheN/UPvJht+FzwRHwKSt
UhEpPr2rhrFjB5H8ki5+9MOaM9W43YGne8nD7Nv84t8qhsqMe3tRjBD3lLW808WmUyLOsyePoNSB
x8Q/AJsoz7OjFFxOkuUJf9gS4qCDPFJR9+Ds8SUj8bQzZH+90Fs3DTqZbZQ80Yt+HeVUjD2ES7E3
h+a7x9guh7fK4SIS89e9Pgi/NliqD/nDu0BllOA9GJf1AlmKhxjuXhH7OI24OXk/xbTs5iWeLtQq
J9vvOQy/guLkeN38fYad+T1UzdClvJtQPG3UFwmT/AH5XpXGZNhB1ehJ8NpK5QTtDc376vRTxig5
WBaC2U0n56iUUxD7w8JfA54u5IxjgHllYUeA2HK4Rv50NQcz3x99uhcwb1jNO8oNgO8bSDo3CbgL
sr/2/+xp5uSdbZDL/E4jLGM5qnaEkyTdjWJy8v6TpKvqW1SCJ6EzE5Ricmh8DgSQXXjJju0gyY/5
2LsC2ywCM6sS0inEaNKu9UGTM/DF+pKZlHDGrkQOWNqj7liP7jjFcotSiLYIxYmfFAgSf+z3/6s/
PzzwMi3EGHacUUM2gaen22OiExx8+dCWRXULe+8NfDB9UfbONXGq7vjIl/cqjOl3Pkj4bxEaBZUR
ZXddVmCBb6EglZgncsRoqnZhH2lg/S8ws9NgTociakImRMyd/HRjBNbMxmjtTcEVJcMYuUhmz6Me
7UlQgLaR5Qy/lsDfE6bvJqOjRYZhvdTTslXIDXNSKaN3AnRS6+bgnBXmd+LXWZ/IYwlmgC7l2qjp
MB9om9LHwHzL++N0Azk2rbsU927Ss/RRnb3Gw7n+GSZ+M2pKhofjvtQVuGqfXHugct/kXo+91vBf
G4/AJGsHx4+J8z1KCTVJskJfqw1UDLSBQyZglN4DnsvBLEv7v+2rXC3grls49WvAxf5nJDbmqQ9p
5+hcFY56ygYBNVkxJfXtNjzmUCcVWry9y8/Crc3Fx7JW7LTRcII6iwT3PctugSM+Aew7g0y7oxIK
N+J+8AEqwHqMyakHh4oHNp/4LWQdDnCGKYhZBuNTMXTu5Yxvsf3Ts1LC8MORdVKFcLDLzvzksqMs
206IZ366IFXoNV8gPujA6A6jy8eqSOYc4cPpRl/0IV0vEJR6cBIY8rYx7RLru6yv0vf7TCt1ZJKT
oihBT3MUhb3+h+k/Mcyfzh0EY7C66klP1vI26w6hE3h0ZO6NVIZYzALRyaKH24j24jkbOgVaEDzE
pEU7rxytVc6O4B24L3G+7MxPyusMSm2FqJkkTXtQeOuiX1D9AKIsRooySx03d0cm/2kb7/sD39yU
GWVm6O3rvUfdEliCAvYGwNHPtZi92NlfMy6OFx315IPATdX9PV4AezDatUBjFyZMz1mSja/CYeP5
G+cXoh4gwSX7Z5hzGs9x5GXg85aI7UCTFL+yNsp6s2RhF83tIG7Iw6FU0T75ZY+GaSl8DZy6qa1t
xT7QZ7SmnKI/o23PaJhCiUTgr8rBMjS1ANP2zIqGEGG8Buzl4wGI7BWvXcc1V4gydM631cWWEebx
IVVag0bUNRZi+4cNKghfJNIwLd4eoPcq4DRtBfGjSdCRt/VDDRsrxUWJWBaiRTQZ6JE9pFtpshoA
XsSyjrfc66QiRoc79l7R1nGG43R6c2266Ei6BjJMCczpOJHUgPmw1xADcbqZQl1x2mIQZaG5JKbL
sEFdah1OmWtAP5S0B7EI4gsoy7osuq4dbBJ6VcS8TI3xiwRyrZErQYyCKj77LfHUibv893UkSsDk
MMPxPkLwuoY/64jNk+ksbhiz1lL9J9QiN3nkvne95O9tPpa23kt+OqhGt/6zqLJTJ7ynD7UEqx3L
aWXnMxEhfm8D284Y9qYVpUvsbvLBWvtstvXmXQoj/DzeSJfG2oFqZZL68gIHVbBxDXonyojQSQtU
BzTKttvqpZOG4B83tUSPGWjC5p7UMa8QZ9AccOIw5vrxxoKFh/Po5kwBQR4MTBqG/jtICQurtDuX
aKZTY7pY1S/8tryxosYjt6bk3k1cyZMz+5F61wG4WG4k9FZTaMu5LqY+7c6h1wuiVCjoC6x500Jq
qOZ2nb2cLn+GylTZ0kCcIF7RLhCreD5iOBp2EIA5DsNekvT0YLptFk/YrELaXfoCqzbOfJ7oHidP
JwvKIDRBhpGhkOsvO7imyOI994rc1QALi/7xh/uj9w4lJZI1Usxf6sIYGYIv/LooHWySNQLbvYrE
wU3UCfRpg3j6gf4dbd9kIJyCIALR69XjjaKhLwJyD+xk5h9RZH4Mz1x8mN5fN6WEfrWQNuR8lnr9
h4RVmMbGCUO2aNThA/1jvcNe5BOqIJ0BX0gSdIbdmdHx4qxTa/jkr659JvrGA9sffNP4s5oURHut
Zr2cw1KkOE0Gwu3Xv6T7bmhLSKPKht5HGJZENwS9CxUJTqi7TzwyIEOcKhL/qKjS3+r7Ps6vQssh
w6MFIHTD/vAhjRT5VtCLPLRdadZuJOT4KAaIcLj9Ky0vg+EJQVFDgv6XHopHX/0znwjg72QxYs5Z
zgZP5BtznxyZ3wumPunjEUmiJQyprxAnL1fLDBiFwGgzFDMlst272A4wK7tmTSbpJao49Vp9T5GX
S1WNf8HBCRpqdG/KDW19+Z4oLPFyadxtzRzd54NQN9clYCE0bWHoKik/eR3B2BqacI3B39j9A3RC
MmbxjlKrF7LZI8/XWwAAz2R9imf3ujPYrzQDUIAGH0tJ8JIvXZavoYOyn1ooQcPx0rRcwpPpK3HJ
BO3Z6Bo9mt5pFOmUWaXRiaIWfBl0ELCP8pFfiNYgWaMH6r0QAmQpFHq3q1072oXtGHPKdIoE8VRc
dUiKKRikPPSdKXm3KUnVuqkiQsGcgK9ac1K+8G8lAzQdkHhVf5/dEmDNuSG2EnzScGZ4D4NVsGuS
yd/3KEWma+1zrNc+ZQgDo4M92msKfaKewEsCC8sWl5BR+xvv6/G8JylTWk6cwhXCqezEHZ3Bjjsq
viVVZ0H7tXVp98myUlk2MD+GU15/v3ORapTekDdy74sB8cMYG+nWS13V2eNhyGDAiGr2PirsvD0Z
QYOQp6CuL8RAZZOwSbZ26duXAVk2f+7K0pyaeBBX01fSgvlnfoIgB2JnUodbdTasx78kcGiNeMtu
ajKex6Lrxmu5EOVi/Se4z2LGcQ2jxJu27KpzINq1l71YugJC/hQHjG7J9APsXXnhlzMYFeLBT5Yk
xtW4VcB3VvIZF/UTEUGcb70mKxBlJIFfp4a7ZPV06FVzjQET/FtfTjCiK4bYdkWo66r6In0PyHr5
ruBzIBVHqxurM7GVFEB/YBYu4TleOELBKl4F/5Df3ge9x/YFWI0PXhKgE8SChJLGn600ZLJqhQrH
35kBboTjLdzIsCSLMrXlQyuQDOxYnMf57snwbbyM5kOH/rqLhWuSDUvlmNwI0om7RwHq/p5jKpgW
JGySxdAUa9hYNZ/I8IY/wSrIt+VDyL6J5HI0AAHNysNYQQvMjrmZ4CeVwZVqm9eKaFJ+GzWvXn22
43KizbgO+8+zh0KcPwY7lcFdJJL8TiOfcY+vMB4voiyu6Xvijs6zhPLJtSlWidjaO14hZaOGCmDo
5mE4EikkqIlI+/uh4axD6d5KBEjJLjkfCk1jwTvAVCIujbsVuxvtba6qfSSOSBYLPgruI2hYWqGl
Czv2lcaNcMFPLqWupQPuWunynQS8lrDgOn2c+hx76ebTiDzp6SWwpT/waIywIaRH9HLQUgYIfTDz
m9x6yyOhNH2/GQIsfRXK2nZ0mhw1ddqpfMoVGAToz+AIjw1Y03qAgNKKNK8eJchrAUT3dck/Lbg0
YMjfZDc/9gQbudrnSP6TgUdrizwhC7wtzLzH/Mf9zJSsC9eDbM3nknUGzks/YGxZPaVdHAh0UYUF
AnHLHdUK+XvidICe/8HRnkychC+ZOiuNJNWT1PqVrxZqqivXlTC6pTUI6cIR3G1Rqjp7dbLqQ+nO
hnAwJ3p+3ARd+LNFqyC/yWPyCoasAb6hgh+QeP7MBV3A5FD5gY2xT36butKBGVjScSnQQXs0tO6R
NeB3QyF7NBpM10XpQOUmNwVDWw6tQO6vdvW6kVDTslV2q4tKnitCn/OkZL8tQgTY8LgnxbdZ2UzD
XoVy+Q1aCqJ5FhrZvoLaY8UD0r6kzkgpAqyPhcbgLrHa/fkX0CkIfrvqHfefVBkn6r+5k0Ht/gyf
i2Ep7N8VbcytzNGKniO2fomb8woI0KKbYlPvaHvL4eZpWfC0ILbDOSCEB4G6yoOIKXAvdzvjLBjC
CrHJ8IFwor9KNeLI/MF0/JoZs1UHHaB2oEA4AhHRvSQ/sz9TgSePU6h6Qx9pZZnz4Z13E1jFgReE
x5n2TuDy2qfr5PST6iOioRfN4qfnHtTulg/jglBPhI2GuqFMjLdScxAjk4LiJBpfXE8ANIb4zVZE
DX7ce3Uqxp+fjR0KZd83mkHqdjkyX6VQ9YgyWKcQMA2UEm3MIsvLUw9K0c5/cpbGIcdsRfXNRZzM
1DsIKyNXn+WHliIf6l/T5lj/3hGMXIMnAxQ5e5QxNidV1vvwtYoOADWKIPcoECu5mvf2Z7nvOs5V
4MCprG6W9JnDIcTyqd1SsVsmAo4BA5StTpaK6yK5a0rzz24kN5oWxTe+mDonBSGXAHGBSq8Ugo5e
NPbK+yjjiuykwpkS6cifGJcT9YWRUd98jvb3jQFOsY6pAwfNU5BFfc5hJsqxa7YN+CdxOPZ9viOe
iMnDyBOCdToRMqYRn0CfJ4G0KguMZPvYVBRAdivgK5lKuwKhQezcj0ZiLT5EW8CyjKU140V7ddfM
zKkxy7wPgKl/B0WWW3bHXgsgSAw1rkWtrXikbxhX94kfFaaZdQomL5fb3JzX1yGWB/zLbzNiak6D
bjsgzBzG/TUs5QNQ8wEJYkU2uEEqrXQYKX7D8wRyArIyflsJNdSVnMclv1BJQ+QH7lTLiSc8kWj0
xQfE0y4tiawSGNNnJxjcYJ7l/YUwy20ybcriZJrLDvtXCTDbdeSqJMBz/G3lWviWrqnQCH5XYQCF
t+HjC9NGHkzpff9J2a+hrwJF1m0DM3BrOWrCc7JWRilT515v9SfCTS60h+fkW5KtH5K++4KehBXK
IKb2DIlu6bTc2LgUIiYx/YJ34xRcGTnt/IgMM/v1rmjlN2eonG+eqxc3vFfIBehzsP9bSSwaLCRN
yE14asNm1mTJbs3FT8QIfOnaufNA9gA0WwmZWuneQwHtV2KJBa5pnQMWNeRvgNJpVVf3NZyeODTS
x5Z/A/IVZmJ6MIA3GZ57NB0e1dTVv4xvRylcUE19ikNPmKUUyTUoP88/zEU8HFrL3KJazC5pppP4
SL6cKER5WXhNYMPFw+GtMaOtTLmhoZQ+SwbYctwINWHWZ8B6gl5Os5ENejnRDkcdlxfD90N8PbvK
35UIb8EjBSvpRAm7V+76mo0SM+b3To6Uk/8X/BjNOTRNVHlcOe829jz8uhNBnxi+dcQcGHm8vlY/
QRAIZsazimXp36cgzFKNAE4YR5h+k7jH8NPrqG43JpFlxGBGSHduCjJ3LLqI0FgKTvFnxcQQPO3T
+PS9Heh8bzG05zCk3WqYtzYw4xSlZ164kM7zISU1ucDnuScumwMZcL8oDNstezTjZmht7hb11ME7
9HEOT9cfHTNe80nPRyuRL8khQ4FNTO3Zd3V9BDUeN8nrAV8CuhaxOViheRxTxGN3UtAVkJzKuNnP
wmhZX2q3WZ7c7Elg/SETnEmmKoygM+nii7HZLXjP8uDWGFqG56BRS/SNgRjom+k8nua2CljSI3J+
UmahzPqkhysqhWTXvi0NS0AbZks7CXlW2s7SkgnpMAjD9dXraswlWiMiREIMeO/gPyve9DppmCia
1reTgTXg0BBbmRcibg7sfLp0FeBccSlEpXffjbILF4dtqn6Z01uY+ZCZAxjMpcR+7bckNjeWN2Ec
wsm59B3fj/+VZyngfo/eLjKx2C9sbFtFpOKuYj2zTnX8UnlrujN+kwSUa85C/p31mSE89GXt8V8c
VTWJMiExX2/ygLCqFbAyedVdO9A5M0ee+hUq5SrEKOaTSCdA2WINRvnFPXLnzGkhUQtfQwar4Pf+
QZn5snrJYGRmr3bfcdP57mNitRQnxasm7NvE08EPhlNNBPwXvd6ou9vERgS/YPsisWne+Bv4+e0A
obeQl2iNdPJW554V4OKB0BLFua70bJnDFOZcn5mvw8G8GSmBZK0rtSPHl29ku+vaU7CYkvJB4Hid
tJni8kbSj1JvqRH9TmrsiQHHcyTPcVRKHF2xBpPWseberAWrsQ1Y5EH+YCqesUQ+pjD7ID/VHzUt
ajuJH1oiy7gB1lZqEoKi0DyAs45nFN+B1DHQ39bh4zymatmHky2GuJFq9vmpDi2Ga8J5tY4tpiN+
x2GN8MblVoa6N/YeXWSqihrDLuxKT+1XtLXzCNmT6656XWvvcs9X29Cjn36SXHbL5KbfkY8RvOZw
YCotD8SBSO/KbfYLg90CYVSU8AVkfVwgBJjHeICLADTwlNFHWNBcuRuz3Ri5H/RAk+5z3tsCw8uI
zC2qP6Cg7l2chIZH8rpWGc5tilbhJ1UVTzQDVjVClSItYzrLCxamhnhx0yAUO7wE68Z/7InCBB2e
EKKc9F9g7wF31RajQeQ0tSEexgeP7ZMpCxHg40uzePZOO4D+O4qU0hAsQzZE/mcc3v4/uPGg5h8l
E2tPYLxYLvzWEsEimu51RVDFyxkd+qFd54F3fNbg3wFvkBvPm8He5umVzOgMYCNIDRqpuYdEI3I7
SiFH6UUVuRt8V7CYDIwi6XnXaFDtVIe64iwQQgCdFnSfwXPYJoEAIXDVVEFSg5Qe+qYOirXTrfYP
ZfXyxhKqilTnqCMvoiuZ5kgViedvvT3zZEL18uIars7aHVQwXpw82kY6SVXyER2KazdD9qXdL9nb
OYc4ngRJhw9olbrRh/nK5RZd3Nb9MccGAGMgjBRmBZ7ynZxC/LEQ5NhkxWe1l5glDexPMN3aJ7Sb
uDY1YvJuuKZodS+IKOiuHYr6ft6/Ju0mpnHVgDgUcUJWaxEamAQOX/06y8o4/EvB7VzLTLv5WVM7
n8fB5LVFbBh6UPO5onQs59o/XuhooFTVRII6tXPnOtjmatJsForBYZ5i4WDokGAE7p+OyekzdYTy
wy0zlW1U9uHhF1c1jxrPcdSFcgWwVYHQys7X1CTDtvDnSfaQ9z9ehmBIppYlGel236+waljooJ4i
C/hIVOxotJtnekehDkL+8WvHaHwo/gY947VvxthuwSkHdgCMB2XtBrq4IcRLWYdhbny/+WRRf0SU
w0GceZq14V12L0Ylv4HtvYMD+3O6n1A6ZjAdlz+DfzGG5ao/dghA5mfCz6I/ZeUIJ4d5WjHzdal1
k8kiXhCu5Jke2xzDqGKDTmqbk+jEt2N2LDVpaXNR8+WoFmQtT3G8gXeqbNOQrEPez2VgX4C4fNrE
BZ/iAm2FiTxLAxYAEmv8M9XUID4zaetaS6DVu/p+emBZkTKjiASB6M6UYMDZxVKtRsjgTD9Iuwp1
Mp6lftgqMfq7ZWcreJkIJb0nwBR2LfU6cvIPSbagqAwkIlXUkYE7a0Qxp9NNMJnLzAWcUkxyOOzD
Rbt+mURv0iBfoDZ0svIw234Xl+lHdJLoxfbuqVpEsTPLhDFzzkctPlS6Cp5rOgjLBqlEGoFJ80GH
1GR5pwoxQbozUNdypt7MSyMwuiL4yMbe000GIehLKAGmPTDkwVdNMVnv3RpzlQFsEtb5VywbpKFe
N+jEf5EEvDV5wMZOyVlP0mRlsYlUtDUpxauv8evvhKbPF99zFC30N1H+PtIBbYBWd5dW6IzSGzYd
6z5dHctX5yFFzoZ8W6soSysDaCDbMio9/5lYqgVyTsZlYNjaeFdX7Pt4pL70/XPgvGwlNCWLoC9Z
o99HKYnGrUw8dcX3mHsxYJGG6NYDEmj7dutb4ISJ5OqLlxcLgpEmtq0t2GurPtx+Y8qZesZhJDm+
L0pbvkzzde4WAQ5H/iNlhbqG8o8/IFLuN1w3pnxzmM6ZN/AHoah4zWRz2XmWbMR5583KVMyToWJi
XKBK6rOCnT9JD1PZxxdf+bqlB/GiuyPeeFyQgsrknN5jcs93zY4T/ReMPBdd5o8B76Q/E993iivS
pxNejyY3FZ8eh1ILuSM7I63FE2gmvEzwEZdQmzIArvx9+4ODRzJDAzgV3tIT89iSEpir89fq6WMF
VOxJb1IDgQaA6pjtAZUJ3j5g6p+dlWbf004ErTs7wAhhi0/QF3x1h4vphLcpqhgXw3HauWsv8Q1r
SSO2gJNwTngyuzGRXGe/HYcvZVsgQiEMLh8Y08UoYVgcEltvLfDd+e2nXXgowOp3aeJoMZ9PFfo0
wfOy5rI8HSxXrqWQQ4jGn3QO5X1ttvrXevK4sXMEUGaNIxpKPEw2eVDrd1M/EJq+FncnIW7OEX/9
N2ja7F3A6hHSD4LyjW7AC6Qv7Ie2XJVqTNEJEVV9DjvR57G9sD0m/vweWvtBYjOyBSCamyfeOhI3
YlzFFd9sFZ+tmfJHzxGJ3mJzL6e9UpxoPO8lfea3RNMVrgf0BySu54eAgR2JYRCvswB9Focv+dD8
okQkB6JfdpQA/Uayrzl8QBaAmBn7Rzp8dX5gPoRugqQ4NE16dL2qwjXgVNM7tv/7dKD/rTVawWSA
0539HGNpi50Ir7iAcXSjSPbrAYaYriHzVxbMWAwdRtkOTQwZ3JqFipRLCZUEBa6SoJJl/crMparP
9LEMVEDL53sgQWmtmj4bvi+cbqJjTnKVId7w6h6CdBRXwsU3gvoFLiw/YvL1E2oufj1s3/MeD0vX
9dI6ympGI+3eftPg09ijsRg/elnbw/FDX9UPRN28APMKs15M9pVizjPMjvduEah7z6skeuq+i3KV
W1hGA+X8jCnBmCJ24iguZjwhSZQJbD+4rh2TAnXmg2H6aZ4Kgop0/fyGIysoEm/a3vEUX/44EwZ0
dMteW/XMiCM9GAMlgNim7ed9DgVyYsGEWtl8ESKyxwV57bKK1u99SShLkFvjhmQo547aKSaOeUP9
2o4xtVAZKVQMvEs4dDw4lzVl+JfjxmCia7LJKZorTOixEcsaRjeUFmK6u6Cg4KUa+LUhtbwgAt8m
HUeXFvN4f7YxaXDa8tvvEYG2J8y/WK64HQBA/cIa0yKci5oZde9M3FKbDG1ShGeUBosMF67zdT+n
nDIzxa9peVKUw+AbPGwtxlokMlIV33QdavO5M/2pqpB8WF5eoiTMPHjsF9/r5R84V9Qk8T3PXRwi
2UQ11h3LoK/dcc5eDbsplusMrgSMfkw5CPlXRp9elHouwj/wuHxsNnafK8vDlOkybG1EYLOlHsGB
VZP81q72T7fZCSPUlWMpJpohM6IJxVp/ertH3XD2fc56RRnOJz/JhrUOJ085TzfjfvAYYfUqhIx+
v3kuRPgNw1fuDy0y+qxKJ60tKIdTDjAUejBQ5MfE0300bipDOH9w000VQNFmSIhA2xe1MMiB3OTm
3U4c7zKT+u40X4DY2vYntJ4Jx5M89u088KFMPCu92/OjJhmbzfVc9Ckbl/+PAzkQTzogjNugdFSL
VQ/D6llNnr76gZDggfagaP1QmZsv+y7B9IkUL+9v7IPQ4WgDzu7ZkMaNTT63ywbuESdY9y5SpUW/
Y5jNBltapZEcn8tuo/hVy/xzJhLfGA1S3t0NgpGbaO7IWhUQbMfsBC2rAx1RtG0+aBSENP2yxodj
f0rmQcnMSqE02ccqxxzhUjpeUOogTanA+HNvUBhLd3+oEmgG2yV3XnUycxj1q8bpcU2qZhUjnhQM
IK0OM5CrGRso5j9Sgsvy3mnunx0epN6rfUE3HRlPjAsgQFZGbMN+2FcyRFHz1cwKZfe80omhSitg
W5/4TlJOu66mqP8vALeCSgFDbOYNV9cXg03AM+UrlflrIMQLfPRpxk3BTku/TpgRvC+9J76PDDTI
KRaaujJ/YamV5+9wVKONQI7j7LMCjrKDWVAHcZTD/hPKWzmhJEkuyusY1M81CEJPiX/O+odJmNTK
CtyPa8U0Ipm3xEIHoHbYYmqT8dS0PPWCizxby8AluWgF3NJSE9X9ezxi0iCQ/xtir8TI7IlQacTk
V2bjTDoxCmHHfkiJL6sQHXLrEvvb0oBZD4vyFR66lCfsKqiCWg0+5xHFV3VhSas7V7BDBdfK9BXk
7Zf3CBI5m1uDL9BNSFhtHIJnZUnyzU/UwpCbfBA2/07/dpfJKweeB3IGQGgBZfUzfBQIJ9qL2Kou
Rc4kS+jVqoDKv0xe7J0k4pEgbsg3bPF9PV0CpzdBfF9ObZ3hfrQ+xYx4Md4AK/K9xomNQ7IbCJzM
JTU9xPAmW+N4NBmZnQnJlk0vBw7pFZ34o/ZH7O6pqgFpS6F/OPVIvG51t7W4RhSkCbkIXw+t6Lin
F1xgQsnoGWP8qXWtBqJHZdEUhNNyC04eCS1dKmCWI8biiT78AD3gedx4nfypQWSVZ9WvP8H9J6ed
xPsZ2S2fOCLi2czuE2KCmVqC1BM+laW/9VgaRH5yjwHCuNxlhWAqMPMToFPqhxKwWsdpnIGcgoVs
WBFTRVpQdkEkPWgVS3Qq4RHOelbfevvw2a+y1yD7zf0HgxVJGP3WpTo7LEtMO9eMHoCW1YeyhINp
PTxcGkun3Bplhk60PP4yMDjsCfxH8szVxdToN1BNI17RlpD41XH9/xPlRwADofHZ/D77wxRN9sIV
Or/xgsCCedx6Eqf73KM41HkgHMyqbfs/mR1yzGi2i1g0mO3jq2PSXJg03B1KGHwckZCVfmwJMKRT
1qUOyFWVXAbPExy10x0WEcEiVvN2xmzY39Xbx1pvcpvgLDZjwwRxHAmvsRcLxIeoE2QrTJK21uhq
5offUXy3K48xIqmhfpyN5VbHUFVxISvN4oxWIGl9ITjm3NJscvMG2NebYvTZdVfDt6/Brdot6ug/
FMzEjPqngOZ/Q3r0IwmMWVxP58SOeWES2EigPqNDjuRgK2vg2KGW3qIFIul5XlY5/EiVerj95Jd3
SGMeoF8AY0UbIw7ZpM06SAlajcDJEjw7gzYfLnkKr89lOvYw8lSTpEmfzhiGQueRpCuaMNep5KEf
F3+WMWjvxalAIomLCDjk8ETIv5/h12bIaz0+1hv3Kqgyahv3rxA8yuImjQ2+MZnObcLig2Im1LGd
vKqNDdgqS01xeMJUitO6VKLkBuXlC3b6KqiPIUoxT8J+aFTS3ffkTTMmYG60A/C1IA/o/P9ltwqI
2NxZGf98gCYItwaKKNxhJUhTfBAVeVRttAObAnFY2ddf7AUTtO2TXR+BsUXgDDHwHO1rCc5hYPKY
SF3tA2o1msJxzbGseLk4vhwffCrjQMQu0lcbT1rzRniGlKzpskHaY2GHYOKSx1Y9H4ZZc53JExkl
ZxM3pWBxmQuTkVrShOnU//ZrLg7wKD8bwfhDf5dW8w70I3+Q5rJpMlDxtViP4jQslqF9+ELyKbDp
1ScN77eIjT8804Qceq60bcsp5qPxBGl+0Rala7oRinT1Vivkt/qMEGPRm6sHzm6f6+yIxLrw3jTB
f+umhPTy5YQls+6RX6ZAgNOBQ7pp+RtqZugxBtMEKXPhZ2RbwJLqLGQ1jdKmHFLKwNw6IOuOkA7W
Bj8Hmk2O3pcaf+5qLG07rTofRrPowBWK2pdOB9F34W4WVIcA69y7+uZfELYgz7H6M0MfwjoxBs2q
ctbf+U10b7HSXVFF5oPL0xiiXBDx7jBkt2pjqiG2qRBiZU/d9FCMYsFczwf1ksdnha5C+vDog3rK
BdVF/9dDz1Qd447ZAtpP0gcs5qiQTwIcw22HUvvLvJr85IRIf93j4ZQE+X6DlFOmiQea7sj+4RZU
2hL4psf27KKW/2JeQy5iYtr3GUAWHZPDI5T/Zi0Tjr+2W5TNqCwatQhVlswtwu9X7tdgezJmy0cS
8njhvr52n8NeruJOIjFas6CU1V32fiUWngMHeLd6FjJfj2aSlr9vzlws6Q73ZNgmrb4bThy7o9Yz
aqVr7ixyVPHqsmUOQDarr7GxPIBm1xDWWV5DB2uO+AsXamDMHLgm0GQCAatBTU8YgVP06doFp7Ax
CrzMIQJBQtEEojILtDxXmuNCxWvkk4iPHP50Fqx1dSZV9ZFAAiUNY9L7y6bSBy3lapGryqBD6/Bl
K9ZDcb6n/qhuMBdRb7is4prpbAqnUFbf6Q7DC5mUqJIEgAkY8FcF7APxcHt0FW1JNOlPo6CsxT8h
vW16oA3nPhJY6FiMXezjr/TjrZWM/wZws3jGJ3krByVCwfPuX1E7YJesaTagtiKbrMZMhM4rspvT
64FeJCFfj9HnSNbQ+AJCgxlWvYLy9nHvNiOeJpRGga/T+BmPnln7XY0m6svhWd6R8YbRSQ2b4dum
hKgBXrjWdZbyS0oKI8jRDRvvPa6Mh5V4RRI6o2pVXp+UlJVlCPDfXvLOk55HbBVI6nTNc3RkLKMY
Zsp2lN3nyj29YgzBH47brgdpg7P0I+l1Q02sU8wYLAswcXnp8DtJaeAvjpPMZha3+ppFEAOreDpa
yTFiV46hmSAufpU/xOoS61Xnm/oDAuOLa+x+05Ym1brJUJYlp5pDiLwg7uUnVCEMkDVpAl3el6DY
G0OS7Jrin9RGopQsQYmbW9hX4imq0Rw9ThcSrdfabWmCWuvwQ4zrhL45a0oMEYBd5ws4ca9Aq9xa
vajUGmBZDdl1WcAlrgmYWWtJj8kh1Ke798ALkysVWdvfT6pcdCR50KSjFac5r6IWv+VtOTQg4Akn
ASCVJy+6KhS61JbxKQ1vZh66IpUQ9kF3tlIWL+N0IrokJaQ2cDtnFM6GczX+sBHduMDatr9h2l71
7px4GLra89wW1mOfBxj+Ttrr28Tebs2ayvjwPXmXTcms3iZlNRf1dIBuseZfjjJYOhEj116y8sJh
b9hdb6OOf6mlr1KlWnZI1l0FpQJBsElAAcQ4emQ6xFqTPAkqJ+4fmdz/0/73daYQogClbxKrwt+6
MqXPOlnW14evPJUX7Ywk0fP+H6aa8r9jTHwJlf1Y5WttbBr3Cuyu3yD7gheyK8I0iAvPcCsOP+8k
TKoPxn5f64umtOC8umQ47Rn60UsULvbvdGKg0Wp5pJiX4YeA5oNzUK1IanMY8e5p5rj8ZpVjCsSk
ehlDnmfQ8jyaL+AjaWqdK1wjp/MWhjuttRb3crsrtO1l7i4IIuiATO9q8SJIJEog9fMrzD5w0OJM
SoJwGlmvSDZKrdUCOOFCNVtp+PMmM5QtTB2e/buihHkcrulv+GiAG79/Tfl33Z33wG8f3sUA50rc
CRmUu2jYAZ+mGynA/9suC3aunqvLNA4iq4Oy3GgDhGWAObp96IMyJP3NMVhTook71MdufLUnL5WM
cspWvgdLCsn4AX5RAslNbWQTHln9eZVgBFC05CT8oNz0MAC3nr7YXvxJyWy2Xyres4wnQ5zki9AH
ivGqtLXbg2DBGR5pZkPmhu40CSwrrfsU7mDOoHVOeJb6+6kQIwcOIqAeBqhw2I7KYtFd7+UsPRuS
QcgUPv+VRvwIj+zcOLQ+quIIxKlushlXOio1R0x9ZdNECxU7BsNT6cogKq4mEb6FeidzlnerPag8
a44mUYiIGQUrInMsWbF3hwMfJSOwYqyZ6Yl51vrOebPsq5Xqnxfp0PtswKz1sVoA1TzcegRnRpCW
WXUD2K/57AJD4wPX24IYeN276e/K/hd5l1l7Px9MAuTkTzKSHLpJ2Avj2ALby54nqSsZStITVcNG
pt5Avqli24qiWXgJ6kZTK3XFreelTfRYZQN2GX6+6Hr9OTVmmmCOY5Wm2jV8AK9lWkhyL8obBzoo
jyBcHA9uU9cXleL2hGg1SLEUMkJ3O18DrM0w01BrIN+uCfMV4zZHCao1OKy6Ms2tu/x6fkl30Wfi
OlZo3nxmnDvuro77In1I2L+KrgaABkThI1Mt/Kd1D5/XxMMPwGkVY870ts8dmKA+DaMUb9W6Ocgk
1MLEXO/Y/hZfqlUKQQseb1NMjNPQIQQmmWC5VwfDdLu31bSdvxM0VdY1AefbRrPSqYLt7Rmop7NR
1F7+BHt5hny6N9wXz+4uogCqH3wdvjBnpzu9CLVIgWAdn95erxH67tHHIQrxyp2laEmLrWtOlkQZ
RsYzDH7cYgJxutdHnhjlcLtsC7jFGK+NGV1YrL8Z4Eo/MdsRNITkbVobq1MVsB3dbjmRyY8wZgxa
Gsv+wmCcfK0RZ+6VLiw3nQ/uc8HvQTtryVaXqTRuvboWEkOyQATMYSOMjTJXq/fYbBHM+6V4VMmt
eSyo6n53V40+KzWu4n/hx9KDUwadbtGkH8albS5uiruzT39mw2VabvJmRRD7q2nidY7eQzqcWjbD
DYI7WwConqGm7KhLgVNMJG19EObs/NMJypnnDmI4vvpCxTpQmHfoJOXjWlN19PSssf5X5M9LJsGh
6G+AaNZWrv/U+29a7TT7FnIGjUxsGo9ha4Rr+8V62kQAq2TRIVPSOejjJkzjrSJUHt3L+d+yY+41
xSjFg4eXnSTz5AbBpmT9TYfq6jl3C6RG6pl8c6wvuRoIBadsA4Y7ntdWb1tIIK39H4bw0B8acof/
WSoMx/RGpzAcaBhnq4me9y9JjFB47+ZaUFUp3uIziwg7q/LVfnp/h0E/BGKDBm+mZ1YQlMSrsS+j
tvG2u/SfioBBplHGVXbzkQCNK6B9Zrbz63TNs1zEoy5JiF3bHCnQ+XydSp77T5VdbfmqRYJauuNq
pkf2Ip7rwjsVf5eD45qSilMwioMAM96PGZaxhifyfHgLuJn0+wfLI3AjEIAVqcUHypscyHfRTGwl
mw+H54Oahgef7QmiOr6TbiPflcr9P0FiSjzBgM8q3tP6rah9nv1z9ldk1qJR9y0A6SsaeM9J5rD8
rNyyfqV0ur66JPOSBa01ZXMxOI7itAWhnLmzk4iADR0KGcNSGDJDmQeNZo8GG0LIYm7m18jrI3NZ
0cKSAZbIhu/009jGcxkTbObU5TinHEnh+44+WizqiajsecjJvyn9zBjt9ABTSDgsjVPwOIFpuO8d
oBa4+Gw/Uwy3mcTmqUPSxjTEWJ2MVYsjEws5iQt8Lk6TcmnktfkSJkVVcGvGn3fmYaHUbICm0T/I
SXD6a1B+6q5txdIEhbNwhJvU+1ywFOMkrzPl98wzIr6AMtNK7Ki8tgVQFfRz3YS91qOQ06yNP7+y
CCU86uZmkGw1zruCwFZp+Do4+m1iGpItvo0iX+KAnXoBcavW9ndFcUDS/dWFI8Plc6ZV8qEm1PBY
CMUodnA2TqeuxH/l+dDcc/7wuD29Q8g34VHxzR0DOeqIJP/BLs1yTW8N7mchqOO6uJyRZXnICrg4
OHQlpp3OlgZoEh8umoc1xnmc6k/kQ0jELL1ek4SptHD+lWkj2jk2OUzuEbARfwXhtYqVY7+uWMVC
FJR1rN+QKyjBEU9h+hLI3T7llWG2KZsJY1q2PVW62MMIYcEYWVjDTjMxpjmunTGaBRdyxTFtIpm+
JUoQN0IBbzNQdZI4Kwd+rr7Seu56lG8HBf1idEUN5fV4xps3DtATfLciARI025xkxCYHylTiThFz
sK/oG/gvkbkACUFdrcWkUcgaibi0yjM2JCa7oeBiMILdOyRxoGgmXvkgpAUc+Zd2F2FwBwfF0JcM
m/HPEzSRrMcppb6L4WfigNglvcNyqqtaZQQvPGKU9hydf9ksaJ+WdGnefqSJA5ZlELqPO++mzZPZ
TkmuaHkiQ5UvuNv0h/eTddHKxW1xCElOCc0R7upMQLPkVq/VAthrOLoHMyOnJI6fQxX4APaef2Qt
5yle2MZv9KZhPZ2ssuwkxbv0Dzckd2wtuK8aZH19MWPh57bxJRVy9n7xD09Li0I7p5wbSwSVYl8o
WYkiI59NyJY4rlMAevB3JKFq7X3znFpZABvKEOnb9Jy2Ah3LGTKeDkRErCV1cGXxt3muGFVC/x08
Wm9Y2ZlCYHg8kuDzqWSbIbCHkC/A+fGbiLAdpntxKURF4NC8qD21kWrROtYX9NW6cvw7I3lV2RRD
0CgBFV4YbUWM/pf6REizHYYcik+jDma4YXw7Jp/yGdmPn1hoNMUOtATbojww/nINHRkFeRhUamJW
atSyPOV2MIeYDW6IQVoDi9k1Y7+BlppuaIfjtulz29B77h3BL2dyGiZ4SdowzBDGZKTGJk2hZyla
aLpbNFBbHWDMuAfn8qAaZz37q8kKErmV9OxQiG8d5ukHJGVcPbt9jNs+SGImWtdg6Sc4Gth7hc0j
KLSUwK7cp6Ty6GwELScsTO89YYWLGoA+SBam9PdPvVvAyedUThN8J6crEQlVlbk6ErzCpemAmrz3
zyxF/s+BjO+SJo31bPKmSi7hjY3LEjPXSEXIHBL5iqq7Za6dQRRSiiL5BBhYlGhAOeMMNwo7jbgn
3BCLJaME4d+gK9uiNGVSWPfQHvuT83u/qdF8ZmlPXTql5AeN/RAG/Hi+S6eWXn6ESKydV1vs6t7S
cnpc3yNToyhxbZ6Dd+lkBJIM0qdngDXB0dnoLMGwTOfZnwiIrybDvpxn1p0WBnCPFVpV11qwzwZl
4EsRXjMtM4b76YEIg08mbzqSs5GNu82SjxeZZ2DmT/G/tRH9OQzrhYH5/Nl5NZUMZTqy93o0jWC+
njsk6TuPI1Qlb1kFi09JyHMzG9W/vf3JhLmDGwKFneBh3aDwBQFSOlCh6J87x/VgTZs2vsBZjuTb
t54oR7aQHk6ZA4V2cJNCvrYrtLj8HLkDF36YfdxmHjOZxx5q5gqXHUIrkGqxaQBfC5D8sXuP6NwU
wbTBfer4hRfeS/szDNTS0ASuS2vo66TWp5vF3aZwQuB7Whqn5QQVbd0mgvG5Jr2/GgqX4n6qC6vX
8Vd+wCQ5Bf8e9maDO/flKfAGRZDWBrJTpE4CnD2ckZO0drNLOfZTovDRJApKg/2fan16Nxu8uCR4
TEqgBpb36a2o0P51119aRCi/7NShco2sbWMupdzcJjAozQ2P8XhZzpRlG143xbvtbPwiLWRGyKuL
sgWrEiVqz+4Lbwj5pQx8I32qoh2docYwd/XTRWu74cToCQAYSI7BM3KttwoLcDv50TMUEpHNpbT6
U4fxNX5LnvFI/Q+aPv/RcO9Sx6HBxuLEUbyQb5En5yzDLz6Yq9t5Q7X2hxHI+1oUuNlhlz1RgFxk
r7ErTyMLBMXfHfQreTUUpOM6aJ1smqpZ6Fp9LZ5/b5YW1FCYKdrCylMjoVo9rvg1yLyOsL8jMeoc
8PR69QPZvH6WAYbBTb4gFOu7K6J2uP/8ryhxVThYMRDFKZ3OqQ+lERldm/KXXRjiYQzkanYvUr6o
diDa0BGrYFUpxrVWNerDqkQcruZBPZ/9cqTiLAdHZIBzhWrEb58WgOHJmahSDwlYOuSQhwIUNVes
bPVsPMw9bqCbgS4QSJ43qi3M1Cu/SeP8inGjzgW9cJBgpWfJJy/K0wGnE8THRV8TR4uTqwvWqKq1
TygMQvkFObqSWT6/o6NgukxUhLLAaTjGKMEWwtVIGvzmPMHy8+KELcwpU+vQxUwbsKyEANVB0x7o
XN9qcg8SFdPO1Nv5LHcs+GljvstIhUNOc4bSViOCVsRAWoEptiZSxJgbkf7JjuWz5OicgF1sQAau
sEql581jhqdZPGl1JE0LRPiMGp8jdNMM1uYumQLdcLjD7I0GY8tUlyEsEprx2FSk++zaW9X9jU9J
XiU4lBQMwnD29iZcdJUKtoJCikScQaPRopJ1gjLLbQh/NV+qQb7vZICiczTU7S9YhLojrs7fgUQE
jWjpcCEVUwWTBzEO/28L85Cpb7D3IMIZ6BlEgYRsfw6JJh7w+0ddvJzgLSDWXMv7ETjuQw+3Rl6j
uDvcDX/g/Soue6mTWiTXBLJSnrCTlZoVNxV77VSOs3cnfXAvl0sj38wg5Xz/NTO5WdcX80+TjK0i
XfAdSoUn8QqtHqgExnoxQQ/MVduhtQLPmA/Qp6eOylekkJTnq3EFH4ozVPR0umiqigSM2F+dBtQm
fWIpQhXGXhvOLclBmbRKL9WYM7sfw1OE8ItXZiLCstK3gy7frCnBpAfGmaRNR44VGDmZb8Jf1F6S
TV4GNG8w5CL32Uj36A3UafJTioKywCGgHZNYCDTzXw6YhPMw6JuTJ2Wz+jPYnaOSTyriW7og6SlF
uu3kWx6m7rZX/BhJEBCP3h004GuSrTxJ0QlRimrlCoNAllEeKS4z0+pmSTOhYg7GWn2z67Oh7yBl
m0MXatQuQkXGmrQzob7TWILndpSc+X/gI4JJB1SJLPICMP1dMclZsGxRD3aK21bc0UAvyX9hlo3F
g9/oNWZ46gxF7yhTSoPulrnHLYnqQRb2vxBJZFeJ7Jv9baWslJ6uJlgM5H+qoaV0yNA/8awreP6i
7K2/WcXc0N26FJIiY91la2TFxzds5WYcY7tlSYqH3lKWxewd7kPrFIddyO7D0R2aGlAPz+IHrDLD
8rVLmyrWwOtVyvI7XCdQ7QnmKPJwVT94gos6CpHQ2U/yKJdR3IQNnRXVwMWgZ3CoUJI+j51DUi5i
uBT/05VdxZSQx+Glkf5PqOSF7AfUMvEfowJMw/4DrrBX4wt9Rw5LOkK2KeUUNSJU7CrAaWsDCvRt
ihXyAApdOCyXaUHJe+LyQgtmBuTt4wGuS2xCJl9fNjq5NjgB8pkvwJrgpzYbR/9MPwYHzHjJyyyF
JhfjXtnF0q76B6hxdFkz9G7VtuXQsUJJbg12QkG81hD74aKCb54QwJVYbV1T93Qd62QK9XyoNtZu
UFcPMoJ8lMdgPAmYcbW3h2oNjdD1zOeMrvU6+H2YP7ZT88X804uE7Z2MBcXIDRgTcjfQF8qEfu7p
vO5h/3byiWscu8bMb3SDviSCij7EbQDRg0NhIzQY8TnPPNU0AN13KoWQ8D2+8y7X14O/Ai7hJMFA
XAIUCSJFLqzshoYwthFGo43EsMirSwBst40M5f3XSNu7VJF9WYqE1i9LhrG0WtH0BxjO2p3Qt7UO
8pjm09Cdo1eDzhvmzmHcTg1mhTBDqo9KmEbWxopRVnrKwYjGCgUBXBPYXifICxWJz5xaa8h8Ds++
JISXjcmEhce4qHvFik2L+32/W1vHZOzTZR9lSBHUztKZqwL4+7B9rYXC4mD81gbMvGMFFNYncC2T
xcuy7NcbROZxfaFAidN/I/bWuZLkjCmA1X153/K/iDk4MWA3eUM3UFm4qViLGwOIW1axaXpjJQo2
WP/DrmqCNe6TtQRJ9aS4wm+DwNnPB68C6399/nUQKa0t2G2D6mzcfG5E7NMEvw7XQ6mkJlsxIz2H
kwdzKKXFnIVgqLWc/mpdzGWkOOfeupuGSGT1r2GNmXsF//XMZ5zW/QN9oazTzNr2QIRnQt3J3gRf
Ciy0beaYKx2+94AM4iJZYoT2LE8LBOk/sHRd57Y1Ie2B/sDKpM34/M1gANgjM8RABY2YPhaJJIUu
U1eg9aM4BJA4gQgaM6jB3U7X15W6dcPQKibcitGQxQyifztEF5b6Id4qd0Zkz8N4c04X1oBsPl9b
IjfjJ2mk+aVcvnm0AYj0mM1YRZFJqSMM94vcgYONyKtjkqBPijYBy/1d2AGR5RbSJHNoiyVWg7de
ZnTZEarLce0Ev3iUF3cEiQdvE5RnS0uh9wB6/tpfx+3LgaRIZ/1nAnUsX9qWnZC6jt8O+VNOoYx7
PMcyiKhlPdn8fWrH6w3xN1L1SZpWxWDBA2fy0DPUnskPqg3yvaK3cd9aqFhN4idk+bBFCyL0pxGU
h0upmfGa9U9qNJNj+Nf6NUqVLkjuNNv/9w2XIleodlUHTGHCaDDxZQHDZwglaKeMdWEpiMtdZveY
a2+cTsofSnw+mfyhL+i3c8/YdGiD82WbOTi81hDFnFWJIWp4iRMzcqw3yVoWU8rROY8HUuqJnTgD
zFqSCyAWFZNSDrkNUiHN7QdDCxr7E2myI12nkpxu2PhNEmzgGipvMYi/v1mE5+P3aUz7sj2z62qw
kK3MTCPfKpD7kyc43Ki/AcIteKyUJRy24hACPjWrJF5OJA4LcJYvXTC7LDosnhMcqmA0alRtuDDg
U6vEOK4TBBGeWpYjvRhT991LAZlH9vH8MddblC0RReIrxRIyEecNos5lU76TjHh1w3CpMeioM3QI
VzTulcae6LYRzs2tPkMo1ltu6laleNFt173RieDYbKpnn/mu25I2B6VZ9Kf2IbITQkR5JfeivkDq
QxiYQsTLHQ+blkfnETzfCGxcuraVqak49FKT/QdnbPZEHyTIrmtpn+6ugUVexf+4FhZQvMCmorLS
OsdUovdIV/RsqDgOW5oKs3ALufd60Cg6CMSEbzN1W96cw9fHFNpxwKkxTdbt8bjJ2OR15SrqedV6
2U6ywBQLBmCbQ4+3q4oe8RXPhopM1G/Gt8U+l1j69ME6bKiBew1at0UwXM+yKHfu/CanCMK4p/p/
iSgCFSUmhOcCAoMxjYn45B5Q8QfDapTl4VkSJ2tIlQZTYolMDyxQYEVejK3ZV/pUVGGzJWRI/yf+
bcYcOCkVeQxH4s2DAVV/5MsVN0xLBCTEiu8Qf8ympAu6EUkYndsCxmRIdu3S/w1AZz8mLEyhg6hT
ftcHyjgKLJFYD0rwBt2jiOGTbxGff9eCpXa/nBo408IApyTlEHMHk5BWTa4ccx9X/sNgfh+ZTtRR
kqdt7XZz9baxtKG+dFAN4X6LVNZY53P3LYNSk3TkrreLt9rSKeRC+W9cb7vTbalXzHTcG/hdB508
shxBVsLrb4tPJ9JYEJAySW/iZIEPfQxJ3n6+qWecegR4R3o/7ypTo57fsixuJU5z1tKit2ApDKus
2wODx7gxqWohHqAbOxwgzIQ0+CMDeHYIdIjn1xraNBaX4jseDfOxqWN1/Kz6C1+yFnDBfoA77bDj
BclkhGuuwnOGQblpKqi1MjPgShX+KmipMta682UFFJeI/+I2iZFVXr2y0nZZpWGtKn+VcAc1ImMp
Kt6RE3N0IBwGAxrVJ5BeyifW2NZyiuPigruCkYcUuMf0s2NLFReGaBDZiWv61P40GlDD8eQKx+cd
tX03En7hyN3ra4R8+s/ZFK3eQcUJezJuF7j4UiG8FiQNt+AkLzfBIL44g8IhPHEd3mlJSyIY9ad6
gMOpavFgG3hZrG8BgL7Wik5JrOldig32R2WGfN0YqeUDM4Tq/YaavjYpneWplf8KnrAmRT0YD94u
x3atmiLKdMNu3vG4L//5eap9UBv3pC9DuY9sDlafoAOF0DCrh34CJdqcd8XEcysp/vm/7VdxbGUQ
00DD5qxApHo98bP+jhEVHDbXf92Y6jE6YXlsvBq0swyzFuvwkWu2E0PfSQae3OJAz1cwQaLpVs05
63cmN+QY2tL9S087tzQQB3oJ6NEbRFZJvpRkMYJ3Shtjy3akNAcYomIVetaXUQum2M0a+9QwacIG
JVAh5ZZMQaIyWWWFJi4Jopgsojd0eGldOLrxEeI3knhtK/XSXFKaZkgRzXyk6MOcMhoqGftMV7dH
fcDZ534mCN6ws6vPwp12mh8PxsRH7dFd8wTQxhrdy+/K/A46chsCs9HCSfjD+0xA7zK57tphfBer
qPbOPWusbgtiYBnh37Wnqojf0W9VIcd0De9u58nk02v7z2RfRXN7CHMZg363nTJyzKCVQWyr/o6r
LpKKOnCMAP6HsKhFmSRQ1imQmNMm2ldKpaosv6K8n/m9uNb8noSS7nMUhPir9IOJvvG76IHQ4N7n
Q5bjQgqzzuhw0ZdpOCdL2KDLgI3WyhuadbkU2EJV9bzcLSVdSMqV+4IHesViKQrZelDTuiuY911G
vHgHYql//KD9lK280xrRyO8OCWNHJB2yvPK6WsK729C4ZTXXtwHWxRcUTuABLB76LoWAibuvBe85
Y19wuggipsvkX4nhq7QOMPv0GLoareHRQ0mF6m3RW56eJYBzgoVN7qvnslCVGCaOzsgS4UjszxeZ
zpOesXRED53qe8L6ClOXQxf9emvbez1u589QHGoxUfa85mqhmpnNHGAFg0l8ceJRqoxoKfob/t6e
Gnxbkv7q/jRSudOGgU7kEQkcqsXBLD7U8tXcTDTjNnaAsnMiUoGJhKxggX3C7Q67u+X5sF5vfAy8
g760jsq1ySJlQcfoOwZAplvcn7PK/gTsRiMfD9dzOK7vw2CXTnXZh0s5g4oiRiKS/+gfL0+U9wio
loQyhMipGfE0SUkG0ZuzN0ynAssiLvqUBL7zY161iV1mjEaLpedCGjRMJ5xCLLT920SxGB5BDv7D
lm2WGpjylQ9P/IXX8ZOCLupCUpa0V0FjIFc5E6u67Hp4VtD6KhCbomXSq2tp3rewgQjCVWh/SXVm
+LykvKMPwM/dRyZjE5xFBzGe7lIxfELFn85NPDMBkjZwwrFb3V7BDjrzd2sznQWrACrSAkqJnM1X
fHM4VFKehXJgJBBSo/8ziTq+67ZaZka1uvxx/bOpIR/oMriorn/a5O0SFLsOEWRcJAoL3op/lnim
1o2meHslixb3bXh9EH/dJDiqY3jpao1KEaAjtfjxHU228fsdUIBw6uhRtfUYuLYoismg+ZHPcCuT
0eHNC2g0TUi2vq1tj11OAFa8CgzHceUGPpcmzB5ed09tHYIYD+H4ABkFlj/nft9dbqiziY7NasKJ
cFPItapTnwRpCCwo4rDA9YoVc76P0231OfnRkOJWYXn1npVKp0b2PnudZKldMhHUzEtMzFnQwDyD
/PJhWCGY/EAb4OhANcDsCIFOuuvWoGMajle+blmAIRB2AdT82jjMovrg0yMZCs0jjXsUZ87JKFXH
ShfsK9xjoW2hgS/gP7/bbecy6UzCutpbFT2MLXieQ7tmZqUFUnXWi0WSFSd1xqtLg1Y4PL4Apptm
ZM4GlYMPEvKJofXLClrG1LmqiYRih01JYokidCq0X2Rf+MSZkspYB2i//SPKa8qfmzq8gQFMi5fI
CUbazYClVlkGROEi7LFTr3fB+GphVUX5AerpT3RydkLD02jRaU0xOJ86nvj2O1oxzYWSmAQr0Dap
VkBS0i1jcYgFbpP8iDyeyF8LTTy+Ag65IyNMuVWC6ZLjM0ssx8wudZUTr9ULzctke7teXKqpfW0W
D7ZOTJhedcpChPGBXDsnQFAi2//GNbkV26rNf7/Kj08SkCiGzNiXsydd9BdvfGX1i8y31lSNt378
+TEtPOwxtQwQbcyMmi+O/mz0VrwdVakrW29euhfbHlorOH2PLmv9tU040hxl8m98BtamcvKInPY2
1E4g/hZF1Kf5zvPYH8PPb6ZRAYBM+Y2heWUjsKVgzqWIWvvunivP+X/wd59nrxAKqBtiqPxwZATu
w/UoXkksAfV7c3XPi7pYsIYWywKasNQ1MxBLm5Ib0i0xQiWDxRg3UK39xZRCRfYjK62gKvims3b/
sc+nxVcdt2ippGZAggoD/zftRb869+GuqbMSsEwEb8cLbU0y6dgMtNxdzql/hotaP4myZa6DcUr1
Z7FTC/e1zVUx+huPRRNHlBhsZ/NVi3iUOb8IjD6S250UeDj87B9rqMDR6KBxfC/DGhdCavH6QNx6
lzA2ZPBlXlt0WLD40BqejwUm8k/SPVCIK4HJAITbAVABGvQ5H2OlZU+h24k3fI8A5NXOa16jGhR6
tsVzi9ZKkBJHbgUu9OgSOoVliGWeQYsb9In7RwhvbGPSYQhFT+17vglpFLKMAY+VFl8GdWxWPSCt
zDqXbCmAJfsom9qaFFoS3UPdbbI2tZDDHvYiD+2tCINuw0U0C9bdGM/DSVof+OqINl70/Enu7zYk
mvN3GxumwfyEnQRo/bZnJWCxBo5OPN7LXpiCImnGJWdi0HLRA6Oe8663K5JriR61YBvI6rdPk04r
zBlH04Uu9k42y7xtMMbXngTvdmai1lBoZ6kwO+fwMLTHV8grNm7gPpbZ5/fmlkKyxHqQogO9aioy
Orme5u+AVzMvkWd3dEDgnfmuobwYQm7nX+NYLPkPdZpOdWdQPwkW16BFV31w3Ridsefq2pZW8jp9
2zb9IxnPTDDeocM2ZApzqCpRkophJIsaqIuhZ6J0i5AMZihJD+RlG+C918yiPLw7UHKKWJEdskdO
Z04/MnXRnK7qPKrmfkPkKIdwHnNXXFe57zcCEbWQBetFAqfnEecQvW+Ixina/wsE+8K+L18gQcrG
lBKzCL1Okouv+7BmGYuM5qugXMKgx1XMr5Qb7U0saKMd3oblaEKbHI5ovFhhoDZwwMnEYMypdUdn
FHJZil09f5jZWvv6Za3j5dkh1BK7dzq2Dr65AecO0SVAgO77Bg13D7TkM2NVZNGJ12Pn9tWu20gP
UngGlo5kPYcJhTSRRBzEi+OnknGsxG5Yv/Y0H/7rWcjVjOfVo5iXc0R5Vc2FWajAF7bG740Ld52M
aZN0BUSLYkxMIu97Kw5OxIGFCwiC1sgs4+O54np2r8TM/rIxm73AxolTXy86LevMI1Haci0SPrYM
Hv2ydW80oJ3T/yvdy6UpiGhlIqu2SufQj1jLhsmgV4s7huWxh/0RFhDRStx50EovlqH/Tow+ZPVC
SXchgM9O4x4KH1ksN26YGvdoldGzBB9B2JSSZwVAMVJvEK0rDIJGZiKiuPdX7YeXuvzmkqQprB+h
hEZBc1dSOOJiulCpiJZt1eH0pvfpKIIca2S0/zMT060CItPn2jGhiOI8GwBiEBnOnqojag7ISl8J
TI2jRFLB6UFDztWW+v3cNbhs6LVafAn2WjBFZG5RmAa8HYRGHAUaZD0N9vPzDKA0v2EPIbABoq5h
lh27m/v/Poi5kiV+FD1RJmzxUXl5uPq+C4ZujQxeCDM+6nNJYLfsWZYQmtzuMzwRV6EtDxrQOKz9
BiNP8c4fb+nt1snwhXHLyr5H9MZH6vCrbq5WdouWPWb1jZlacO5qfDGgeLo3WP9wYzJ4o8e91yED
qK3ulLVWOlUYhpV24jPnfOcFk+CEn0yPxofhTkkZOXnSBO9yEWsNhZX16Nfc3Q/Cu2tGL514rwaU
HzRVPAtujPYQxEd9h86d80Pwt5NSK97aBprb5IW1oi3nhQIxkEL0i62jxS73/1Dyy1fyAQt16mt0
wGP73+XpBDvgTU49vz9vgyZ0iETvEITYWzDGpHX5+E5RaholTAD+LqOcll8j5E6QkiGIHwX+Ik4S
Mwgt9AYIfNQgopGyde3bTqv1NTUtCXjKKgSdW0T58r4eKYOPVptqJHzuX+3XUMwysaHVwENlAZzk
UJq2BQs5N5gtHQonI6GKAxBgneRPI5YqsTv5clygRIQPrgbC6UkJjvNFGrpACFvmQmDIWtuiELep
PLrvJbjI8Dy4ceOCvxLWYw2ZQcuh9e5mtr4ahLD+Ern+3oO4HJInfbVgFrGh1GFyxkItf8rr4FLU
TUOVG8+gIhcEZVCqhn57QUDEhxUICEPrDwyZhPeOFevYpklAapb5ayVknNSsRUwu+nky9qePfi2x
6Yc4MNfZWmHmEJG7YL3mVi5Kg98fwftFJr2W7pJaCXy/TU6fwbofrhSyKKarj2PcWNu0S8wbO3Fa
kjrcDx4eHkQkHmrTzgBpZr6riRMlUQdHg580QIaanlLzAkpjiZBZroSaChSx9c+3VgSu4lYeX/qm
Nrpfyn4I77x8RpdhkTRmfB+rbCkOcgMeCTRrb6bKaEfest6zfOi6RoQNqd03ewzV1nhEVg+7ulMT
03pV2yuApZAAwXh8rBI5bQpr26Nipp0fIfeXXdv2wwaT7m44+1q++rpKKwUD2z3u3+uU6qwQgSOe
malwZXWQ61wNjUE+FXsu18/rQJAxDLl/ZhFvP5vZSHH5mBM5icObqowI5diQeIx0gNpHHd4GZYNY
/ga2MEt/miO9w4uUnE/LU9vU9N5NLF3bhh8IUYU0jwsA99lZQ038OriosArGRv7vOLZhZBYpZa5z
QyX5VN3S0g+sbfmiwaUnxn+ClC9l2qoFjgWbgSDmmJzZcqd9KnOOG9EodJkK5OKzw69IXQaR0PbC
g9R5fJ78Yk/ijTz0YtktJ5s3Pt9mTYlYG7YCdMXGHrX/nmX/lETejU3lW3dpQADi5EZp4pTFQyvC
v27NcQIsBaFeX17VXx5zGzDxwgOSxFiKOqH2zEgC8ka2SIIkEY1c2t/MpP9yprt/GklCIQZG8m/h
gsP5aI/x2CSd+HEZp6BoHylmxkFA4D9/DrXLDoUOreyHKh/cPrKRIh5e3sy4plbp/Bz1ZLgbfkju
bDkdqaGLkRPNzqXgO8UtjL/f678WGoxOEX4IyhxXDvqFXUROZT85XuqYY1wtMJSiJrtF9usOH8Ms
il2kg5REI2PC4Ix0MF5LUBpXvnCok0ma06vvTEG7do0xE/Eh0cpG1E3J0qPUYVPRxl1hcKLtfrA9
z6GD1dVmMbkciyugDIYkMml8E9MiuKepLHgQPAQ/Ghilal7qaiwjICE+NL3j6Vveerb+Ah1L50Zv
aY9To6bPYyltUV8/1LEsW2taMPwjxSJp0JradEXWgLhOyTiDY9pVNtOBXtevhAzfWMs3wTVgnDjR
mDdZUl8iPyqyS1CQtk1PHDEdnXVJOUJD1VKeo1i7YLBBdIg22xiJD9jyA+F9fR/bJFw/NruUEAbG
x+Q37j2kNB/EYxtRJJOxcAD0AGWVFldmMgNIoBcT/s62dp03sdFM755E9XGFIauT9ctv5Hx0RxIt
5oV/kYRSk3deBSRYD+WptCPV34YyAELhE79C0RKjir66mjiguWCPQoJEHR6i/I8ZBYtROdhM0KHH
/jqlq/bhl3KKqqOxxDq1QFKRg2i/dAU8HvZtvwpZjCCckVcSHkGIvDoFt8wTSf751Tk9lGDHfHo/
VEZYHLP/zW5ISoF0/mordJNIoTNYkUetViyZ2Z6KAPFiiVx0FphzLRjWZ7b2xuXPnLsgTeI5ZuxR
r4oys/9DmbjdZNL31S9OjmaoO45MuqDSvp5H+PUuHebAWvdqY41VtVua8hD0w9/VA6sB0RPX8X28
TrH3JSIdsF683Hagrx3AY0h/BEWfF2r/4Ms7m5Xp8ILtMfENODChePW1S5RMLlLn8d310Bk0kl1e
JR2Hbe9xfZqp4JiES8KCC7BHbyrKtQPnndV2DRTprQ2I2TuLDCnBVMFE31KenpHJih0gMfvOxQQ1
mzaR5XnP3mTMjop1aP7uk13jk1f9l+3uSt61ca6feYLZcPumya/svALn+4A7Zy44W6JyLaBQv5pj
tsFPAR6Wrj/nCfIo6OdXvddZk4olpPKqgb9hM6Q8hcVdP7ufaITFAsBEIqa0rU3PoT5DcXZptBvB
jBGAQiuBcXUW10AeZf8Fb9sIWxureRsBDm9C0PeNC8wNlXWMw4blZMW/bfQB/FV66ugX9nQokdec
SxuUGGOW0riqRRs62UnKa4DXbYfL8Utx6470+/u6vgAAUy/ULP9iQBjaKWamYrbFw0cqeshCyEoy
pSZE9Cx1XL3THyCPZzJMTERTcNJMCIeyB734NmegA7PiCe3FveYMPhSa/hXZzk6voukvW1c+mvqu
5WBu3dqvsOebKG8XVXUZkCuPIArxvS3Ejve2Lw7lzJgRAxsZP6f7kuDvREu9iI89LMImzq6IbpQb
eUUWM+qbiCcIpP0pgGK7+fYMH2TExSGlbEtef1IFEKYvNyY3ZX9FKIxKeoDpnJGZ4V8k1n9eJLy6
7HN0t837VGO5OMGP4iNJsj3kw9YnO5kHmOAWLaam4s+bI30dRY5tz9pp6tfAlVqlEo+7r4AMEW+/
+UbkA1Ev1vfH9Ev2rUM427UuIALrGrvcNIiQeji83BT7T2XubvX9A9DFsD7zudOdURmY0s+LSZ7B
co36Y5rpu7MompCMM/G+Cvxrh2gsZ+kW+u7WIjC4iZLogTF2n2YFytM8P1+LE8dFTZsTD4Dl2WEH
ryD3SFEACOMwI+gnZ8ja0Fks4VcKIzyAU1W+WmU/RV2cp4yq9VtSqSKMSDSsMI5P0KXCTBLP4okJ
r+Tp/bOPiFstpfSK7g9NYCfRB09jTMAXhOcm2ew1RDXGnzWBaqK3/xalpUmbKqKpCfeQIWbLHzrj
uxGhT60UhbisVn5tb/n6RDc6ddSFR4mYYTfy7aulcB4/9mXcKRlzCu/XoKynKp4BS4ssEp/hUnCe
wSFVYtR5TKZb9nHLEq83+VB4SXNIsgHUEvKwNrb2p0KqQCskIYXfcn9XCtiUN0HLJllhjduIgAGG
nz2CiygziPNLZP7UgB29R5f+nMDA/8yHdREXlC3tJbM+kK8aNXwETjFqdtrHXLsw53noNn7OlIat
xWwc8iz5aQbJkGVIsozbtXWKV752VbticwHw2YQXb8k8wsjASgQuNVnCLus6fXhoIEH+JMo71XAW
xW8CbQ1/NBQJMj3RrDeJNr+OwvvNseyygiWXufdrthkxLunTckbMKKb0qG0eeSVBnQE9NkLTqhZE
HDmtfYNfAxEwePYI/0TlGnxbAQIy9MqeGaRiLZze2lCrCcnvv6/KjOS/9qCrvtxQdloKkBE9zu8Z
Bze/YruHUU4iCjc46B8biWSQLEMKKyk+4TPPZt1O5sZtv9NgZr5hIwxflyFd+MVsUkRFa/QZbxCA
MwhuczaWIDio46YbbZeCJcjlZKICCf2bpVNxWwsPBIF3KNH8IHPVoIfmdOt43TJM3eauuKOwRePg
+1I8KJBZrycNPoEfUOsIL0XYxX4qMJvDRpGszrUBXhtf+d1ICGK+6qKJDD8Hz7PxJntQvZXj4v91
IxHsNhoa91RT2oqXt/MWv5Kdt7O/hGViKVhWa0IZY0ehL7RYDUAk6ZTRwfKY/GQGTmG7fqFuNHP3
4FjNnwir05mIOcL76HAx0Hmum/mVaIkNg3jsVAfw8KhPeh+hw6IzMfwH49kCtGZw7Aa97ITunAXp
CwZpZb9qGuoxt7hQaSxp+yqACy+8IZ8fwnOraoQZj2NJRsgpqMPiozG+KGKFwui7FXAiPUwJyKOW
M7m4UXd6K2NLNUpB+cqBbpvz+q26WEgzEaedwuAE8fqU7uJgvdGXItDJ/tqnEej/SQuMGzoCoBGT
3c+7qexDJIbWZXqEX2TUtzfCHmxXpzvUjigTIbpcwq5i8lu/i1K7Nhpmq5Ch1c5s3gEqZLsrFWfm
byCwy8AzVFpdGDtoP0JbfRzW6Jr7u4v31/spGrpZPA+r1fiMy4gmNjbPWza3mYhtOpTQvmgk67rv
cmzqtfCS6gw+A2ZsYTuenvct0D0Yvzvk2KXq3pdXqC62RY9vg5CohntaWcNERudCsoEAejDUJAqW
y2XNcG6f+IhcVQFjWjsbyud7qFIISDeCNMm74nOchCHXy3CPaLn99+xIJ6V+tmPBRv+04I1mXDmq
Z0RevN6KZxMA93jUuWkvMYmpE7D7jdocE0dopz/9kY7X3ZNEob9ng5vvEGay1Qa5vqJKd68TF7sU
nQuLDM0O+TQyPUl6PXA/UtopeBIKtq42Jj2ulb9viZvPYJ3QyIgN2YtBr6liiwmW+bXsNNhp7mz8
b8RF9KKHsBNkSTgh6feZ79oM9fOCSa9uN3NGifZXem0EegzyhjMTV3hKq1pvpiKN8aSENaQDAIQo
0SRQOzil/SVDRtSn2ox9eb32u5ZF9vtxvKbEauCCwpQTPEiDnm2dymvbMWobcoaphtfmWehSz5wF
XnN/kSKbraL6zTr83YnqM/jhUpqX79Lic3uNfII6+noaS2vBwnXRolic/6PNlEMNmKOTcD+p+15Y
3aManLteJsBsifvVKjjw5x41kOakOUPGxptlRq23v4lSjiS06CZSeOcX/vz+X0tjuydgnic8eBO1
HYOURkkVULuPCO+I+Ve8NcHu0zMEY87yy5echnNsXmV2kTmQZS7FE3RRdHMwLEwco4+RFO6Xwe1B
3pqBOBeRIx2AQfouwsPMcr/qgGjpD671Z28F3kz96ADFkpLGZnb8ce2KOdIry4nAMaX7Gn1JetyG
Xmc9JFZtZDgjS4jDRRE9hVDnfBZRBm0TSaFYhXaktEXOBEeKYBDuDYf6yd2ktTUOBKeEokmPPUzn
wiRTWLe/q3pRgXgMiftLBOPs3p2uX0cmzlEebCu7tT1RmyWbEy+NzbhLYwvFKJQC+mTB4p/X5Imf
4cbJ+oISawHNdbYyPyfUJwECcnxKKf9rhmdf++OVFA6K5+QY08F4SbYHFPh+ng/2cJLbfARgpsLF
hOuBnNOg7Jcbx/Qaluje73ZNHlOIxD/Vqv/MkIpyXyWuBkPIAaiS3RAVIcm5ecFOw/XuBq6zUyFu
oj4qujUwz2O7yjv5FAPoO6EcUyiZxVFDe+j+6jOqpYkN37odCNrWdZO0aI+PbK9cmXmtQfL1SsaV
Q4/p+QcJ7d7m6pRvvSxaElsGgGC39AJQCvSF0CvMmy5Ux5oOycZ0e77CUW025mlUC0uvh7gx2k+G
gK0QJgYyhldpuqTiXvuph67h0wBuJxvkLO5WEExLIOEcex3FCMlX/OYG/bEmg/pGxBv3H7ldUxwM
q38fg+ZKPXmz/XDGrOitunMPVHRMi1kecxFSNyzLBR1hfVDQ2gLtEGEvhM04do555n82LZHLIyqQ
dcdTpIli3NJ4bvJDkYbRP1de7dGUH/CLYZbZJ/sxH/if70GeSnnfziDk5AJY/3VaKHPHkgljBIu+
GQjprGXex0Un0TJ5hHUJIryGfctSKOJbVPM2O+0g51yNCHkOzR8iXbnxS328mrvJX2E4l9JwGR5+
epVsodVmUHAzG4stMTjV+nZeDa93yRZRezMFG9rZXf7+kzVH39W2wM05K+4swUWitYBHFELmY+Yo
f6rYf6ub8ceJRqo4kQdEBGHhfu4lmM/igiX6WswJYZsf1hutyh0XF9Rdzz2QDXV5yMj6CqzU7MCQ
BzYq4zgFUUdg7vVVDwO6SYiLnWpqEAf7J5zz6NOw+ODdd9dKrQMZf2Z5DQ1zUQFp0zug6hDExLfL
SXF7V8yh+JFJiypaDM1sUlBPrML5/W4jj7ANu7gRv7Ejy7uuf+SWvPsYKHxD6H3aR8rCvNpJEwS6
RLEJChxgUP5hIR0uYYE9bwBFSrxiTMxRxtM/u95f6/Sw9S67b64Vja+w0CTFVRiY2GJlTA487cux
KkOIg7VC/cKpTpgWqYkwd7lOMd8xDcdI14cBryWT2M6qnouyeuQIh/nRM243MBRK9kHTL347G9Wb
D20u3VtsqmpHPKi5VUw+imqlFQ9dBGl7VdcYsusRY8GPdSc6yeige5n41TfQrMes6cFTRDZ96h4u
c9Gzz42/cr96d33oa8+oR2BUROiCUsVKJ8BHv54b0g7Z1Uok/OVuoIJ6W0E5dWngA/RCCQoF6ac+
hRT6+eKIA2l7Tvi8Z/rfUfPzvJAl7ral+ckOFJc/myCDlbN77wL+UfN/YrV6cd86DYwUORb8cp+u
quqZLFKujh2wFmu/uD+2JaQc27DlyTPnh3oUccwUsTVNG0oCVopIgTzGEHqmYoA5NlFr9p3cfsWe
ftHhwlVOJ7E2BIA6qorWPSp+W1q3zOpYNlTCdl1g6poqCam630WhxeHeM9SCxFRZ/KbfDbevDLux
BZoY5SBCGwpbD80lxfh1O/fzdDnCyY2/UClzlVZHvm+S8GnpWVVCTtZR4u3iFUVh56hHq9OEUPCq
3YdjnxC7OBkfr9bKLXiPxDwNE68hrrtUR2ZJJFQnU1otqHFZ5cf5yoT7Wdpxlj8cHBoohncFyWde
Rc0NeuAYmBof667wP1092BXIn5njC4YRMYdJN1ffvp1pj6+0wEqtuFIl799EMYuvzYfOHFiqKDhd
CDPvLblO/eJCzk+nKO9vOEHLGagaxNNLIekbkyVPJoqiXddiDKNsY0/Wp9i0OS89cMc8RRntv3TD
x0hRJvisPzSTvQZipN3S4x+AXCGGsfPG5XxqajbF3HSklg2QWim6IXMEEzGJjOZISP4Ya3Jvw0Hn
/pO8r7gw2hO6ialj3npL0taMN87AQ6sMPDdErEGI9Mq5MOIMfPCafDr5pv0KBUPuSPV44tRloyHh
y15gk5eoWgOwr4LuW6huHbQxJEoHqBfKRfjmdDJlg6TWEnX5KX51+6mhWHdtSpiojmL66YNYpV2E
QfrXTT1+m1MWGd4VvTvp1C76He7qhS/fuL0xJjXzyFqddVgv1Y6cbVQU4rwTdisptnbf8xO3lZh3
yKo4XFVRuw8KtegxIgo5W6UCOfanN9teTjpZ72IYbXzjPs4Ncgvt3q+ugCWPD5HqDt3DFWZvop65
smt6FnqaSdY8A2UO5NSVc8aCxER9g8Ug2/wRvMH2/h50lnSHDHi9MGrLLNW0QgMGpOqy1X4NBZ7V
GX5irjHVWiRTkvJ5uO4o9iVU6NKNbfH8EzDX29xppP7v4FHGuNUT/D9KcFwG0D6LDrAeLkz0BqgJ
qrzf1mSsP6hn/98wo0VFQOVzJh1mPbZIjXH/Cz73ffo8N9HSuS2zn/kAprjFgZJ4DOb8Lzw9IwFm
y56ADPg5HXiZOY2b8po4WJC2bmmJc/EhMA/Yzl0VxKABRicuc3fw5RMfFx6lYw1Wgdy/WxSHMo4I
da2T1uKgT+ACQTn2mxt9ad1Rw+rz2/jAEbt4tqNnVvsIDmPbmSrYrDu74beVlR6vPvc5ukWPKNTm
1uWjYHxR6Z9kLVMeYuDjT4y75+N3S4JRgMk9mOXgYAUeTN5frAtFQlAyKgJJ4vy/D1DM8a+ioORA
9QFhkiemPaGHu2l6NGkNZFTGGpwlv2s9nDyLdauZxBA5ry6D99GCCz3xtsdqXrrJkwUXbJgGKzzA
qwN1vkyU1WBh3fJH7rJJVRDmvqp15BQh4vnheXImmEc8GuVBDKz/gabLaiG886lXRAQnlWdPxTK0
KJpDVta7aD8V+LYHuYvyAvLooGbBKctE0KP9IXP7j6GFsl+g3I04MR7DcTiP2TIVoZPIbzMf+xp/
TkFLwcQ0acm2BuewG1CHV8+uYKpjZtjCBvXc4N4NPY3lI7uCnGqqme3Sd7YLtCy39f+BgK5D9N2P
qdhQfAxIjGp0kdmpJ62CDc5eyoJrxLv0LjhWCl2Fsp2iJeIsKFGl54+mmELtSsnKfuCMzit5rJ2j
maxtdZex6namt73AROxXESFaKTSqmQJyIWP1EL3HjFMyhroL53MxwZ7tuEaLLpGBsfq634WkTtky
LpiJ61iQ6Qbrfd38UnibcCEUxdCZP/X9153qcfJeY43zMwaBXid8iVtX4jWB7W1TaMgTndN00c/x
bZOHU0MOwe4JtHDHT5IPgfJqpImhHcTioioOlixWxESomrT5965LlvbHShqH1djAUqv1pFaRkJ8n
wtaFydXO1KYj46KKbW8wptJPf4rY8ZmDe4hc2uF7pxhnplOcd+jsCPcrfblt/6jhSfMR5ZLiDaPY
7UagTmF6iMrKfRpLxxKH7Z+y1pa6DGGzofTHZFo1iHapKJ9IulHlKWmH/H8160iiuaKBFZABgXfK
P6u+3+jYeot3azyIiywDd2U1XVSpHllVLA/Fqo9KTrv0VCy37dh//nYfptJ9+V1121hbFLL8uvAa
PL2kX/Mup6a7M9UlX4tK40RWbHzgBclEK1SqbuEpdQtkxm4Nb+cFWAnadmmPDfGXjVQ6HyG9vuUr
ndDM1W1MiQ3ZU+BKjFsZVVluBclbOJhDMPnivJG2NJ+5BLQLrTsdiV4FChYA/39ohIBH3BQhl5Dp
fbCFr5AZUjZseIzOLjcGdU1o5zjxZ1s5OyVVuXmHBY5CY5Dd3pxyAz26QkoZAfktD6R/Ko+Malvk
DIEx959o/JbTRPmSkK1wREirebFFJ1QTipIwHGjvTztj3Hd28SF6aQjE8QFoUM2r0TRRnx8mrXZy
um+4bK/jpcTLO465IWvM2mrGzUHVQqsImw0ocF4W81UlK48XF4Xrs6SeJsPAz+EKU9+rFr7O5GMA
uWaSg5NACxPSRq3YBu+kcp6kAV5E2ft/d7SYj641xLVOQIgo61vLZXlReDrGagfF36+8Y3Nu7Ukm
A6/U88pXFzASQYMgLSni16jbi0UMuGpwF1d7Dlm05NCzvAhdspoIbFN9yO88nqJfI4Jfr3cpG95M
1c2bWkeMX5l0XbphluOQSdDfp4O1CETD4AG+KhDHiW3HKNHtExlxLM7bPt4jQcWMMdvDttpHlBf1
VRYvUppB0FNeUiRE42nen/R/YxD5Nb3qqVA5KbGXFf86xn9wXyQ072z8XEXQ35Sm8rrp+as25s6q
Qpu2GXvkTG0fT2iqsM6PW0nogMQSrXpQ5HyVHEDMffuqETJ2uUotx4RW925x2r4MYOcV734dwVgq
SCref+6dGMXEarqviR9Uk8Xi/DnerprXKtnour8lEHOPSCegBfcvjCMF5d5wfSkeXuhkuJpf68Gn
aeXYRBTdqHiAgfltoMYjcoRh3As2ip2wklT6qrHq4PdO7+c3jA9T1XR28db+FG8q/9fx/PMcnBIF
rwkm9jV6oOyyEP9ulMef4nHpWEJtsFKoAw3FKSSIcD248mtj5zGSZ2t6R7LD6JTK3WpLK7OnR4/4
/0Tmys6SkYhnTzBhGONLnZpqhN3Y26LrtcPvpA4l6nLtLU15KbX5jAmyslymvxfXYHWZJEG6LiCs
F2e/zCFHgUYNYLKWcaj1DGy5sQZ9zKBHH1dl90mHvnAaD7BIbqrHlEXewu0m+xBKaPi+oqz8tWyE
tQxMDmAaFBbsi9d90u2rrx1ecUje4z1ptJO3s5UorF8T/CwNLuA+EmQKctlVK6dsiQ+hqN7lz47E
ATh/8hQ5f/sTwpmY31j9pVPPzM0lTTWiZZJkeXhChYFn9G9nU3D1l0vdOhjhryZgDat5fvZALWQH
dLuUopHPYhuouP5SWqOmps5WTGYI0pfLEx5sKxzlzEiego042M8Vbmr9xrB37PJ2OJZ1aMNfbbjt
yDlf8k2iiZKVgU0yNV5rnTSrQc6XGPQK2G20HZwnRBdA1dg1zqPnVuLHI6neuUD/NiUvsYKRhada
xb9WbDIOUvDHr0IPsKDqBcYDdaAWa4VQS8YebIn9mHivlCM+DfC5bNfAnn/ar3BbxGKbw1v/qv/r
HeaawOjfDW8BlZZYzhkwlUn6WiMJRh/o741C726aOXnv/RBCMIKWZukqiGfcMOTx1KASk6uZLDm5
/5tBUg7RjxYP16RD27NALVT21fal/P/ZfMcNYWwF0HKc6qyvyvclzYRbY3oagAYVx4Hl1SV9LiCX
xz0Kbbsi5JlE3JCLys2dzvSQYAvM8fE/c5XvB0JvGMSvmJbWmUzVlVgxW2iobfg8td/fkWx4EnyK
+AHnLBt7Ot2s4DxVc8YdFtrHyveghb70dsavJo2pA2vDTrlhnuXrmXnsk9WY5HjOoyF0NFRP0mGs
fLXjC3bzf2ObV+sKKnuzcxJx+y3XBQGvQ2zFrNp0cCbfWRmKtfgXpHdR0RqN05eeL1G3k2JsJ5TE
Qmfiy0p7NVjYf39nxr1GD/IwQ67hHhhfx8tHO7YMJvqjgd886u8Ci5ylOOnAT3GgSHSIT6bQYGSm
T/oTcfJYB3U0GJ6gmWsTfgpgBAyhpB988hRmo3M3fpd/YYLbKnSngkKc32Uvd7LEh9YS8y5gRjxX
qVN7ag9BKeErwQYxBmcHzvpyp7/DG+p3/oJ6OZlCfCU7hCPSdRpH3Yu/w3fMl8lekJ8/vIEb7S4p
GC08EfU2SC/RvN53kPs9E0CwuCMMkQsk8Q5RXbSeahr+fZw3NkLE6u+FC9mPDnPnoVC4VxqDThTG
3MJdMv8JH+4qnIeHYGFlykC5giqFZzZs9WU53UMEQ3TDEabOoZaUa9XjJ2x3FyD0mP+8GhdobF62
vTAKnMQGN7pHMuFTx7ciCb1/VCZCNdaHeFNV/Jf6yYM6Y5scfivlmXfk36e0lp0/2AcFsblj53B4
8YEZjweqaLe/tbIVS4STMjE+n11pXBHepNT6LuppNpw4Z36jeCLrGOgGFP9PbCB0Bwh6kTrjMHQ4
5pgJ8WK641ysKA8k0rXyJCv3NGJH4zXTEIBSIhVyW0cFfJWnPHk9CbY1j+j3pNq2ZdDSq3tcgZpS
kdifkHEv2vqgT/wQxwhTKCvlj2wCFg7Y8pLLHkE5c7EUq6k/JItpBgttE8002RbmIo+oPe5mVyfV
qwRvNSEmPL+7RO6NKdoKLc63pppvv2Sin/nj+zM1s9gIUtRR/GiykDI6UC8jSOfm5YPF5V/635WU
ybQoIVYQ1eOxRyDjhY++5lZYXfrexqiVSAvkQe0v/854Xt1ZY3IMiRvt25hGBKRTteEgclV31rT3
vQH1nKwFt4WceC5ovB6HCGQx8jsqrimmqzSelCAiNtGTZ8IQ4NWRnPfGLv+JK/TxuRRj8Vlew9CP
tsyswx19wiScld6Moqt+rzhhqxlDxL0RE2/SQxtSbe+hGa+pAiX2puaklQ9UMYyTpEuQe8QzbILG
UqoxJvclqVGjyCeKrp5K3ex1pIN/6QvIsn5X+tQ3qszT/LJpNL+bYP14zSsCeug3jms8r325l8Nt
5DtZGhCw8j4Q3SVz65GZQlBPq/vHR1kNKZcCXxmqTcHJJC0vGdrF9onovGTNL/X7fT9zERNOrl7U
mytCv0b4egjMcbAeCSVJGpqbj0JdP4rzXO3Q5rPQue1jL+4ls7IIrWdkMM6Tsmk0wvhcvuQsZzXE
h1dAiI63AkcppKjerO5VtqHRTO+QxhNULwrn3WxJCewJK3Ok8n9lXxqIaGKx43Yiq6Zcrjx4udGM
CSHT5KUTSlnIwwOTBXcW6O9XZyjtMUn27yhRygTfQ/uHCk00gtYdAF9NuhbGnIkNsntK2D7vTdLZ
GNw6/pM4PXnnZl/uU50hf7SMaAkAq5Izrdd8wsb9AUAV/ntogufVg2fCQrFscxrLkNzgflqlDtYh
g+j01pxVetmjnli8VWAb5GsCigdc0JXs+Z8KKDj4/QXUakXNmCmzbEO0gkf1a31PaSqIlL8O4WUf
fKT2awgnifgcBhHAtIX6azk7XKJ1SxgHa9Hb6DYqYoB9LF6i2bIqQUkV5C5cL4uOJhnrzUB5xkBc
JKELCbrOBCO3kzq7aK/DC16tJUGUdf5ta+H2Rh9xHZWYVk9tZgeKuqqmdIXFSHgNvTGnTxagFM/c
qUwucK52pQVEdG76a4Nc8CT9UgPbFGVAMrj0ADEdtQFm/SHw+Ow1oF5EdCWdJGtyHI5+enBJIckg
JntWFxswuGZkJwG/gYWpjXmeLA1Xw8KHzNhF4Y+9xn++DjXBfizbJPrOleWx2eJQu7/6sKomeoUO
cxbtEXx3i9gZ6/jQGOEKE8ABIM9rSqE7K5Xg+s563wcawLkugFruSauOy8CLWxczF3RDo6WOekes
fYKW8AvEasmXIUyue0kESLPhn5sG/2KXKOI0G1wI5ySNrET/OKDiyFBtR1mzfIQMsx//zW5z0xPc
kpoAIjfiTWi9KcpZhtnPwPlmxeHxshHQt7oDC/7YOwbc7cAgb1IkUTc3hmsrTYz1pymwfv4rVPk5
yssFBdfQ4jUPn+Vwm8m4zn2a+0ejz+rJaubgO8YX/kUlZogUXNl7HwHXEBeHNJjJ9x2r3swRrROS
zDc5s+YyABjhdxvg1K84qZSL0Nj6u1cArastKM3IeH8FKfokQYXNmvB5tev1/TpFMpkpwN1ENjN8
O5NTfA4y5AOjDSmHrKfbefBVMw24MN2c6Gim4zyXB7mNsnHqh+ekN59xt1pPMjVERdGGTL/XZ+5V
KUactRozVZmSdH9Lm2QNLmQ9x8iKiO6wZjGzoOtZMB/eKiAKhYeWTDV1/BRCy1h/py4logjn642S
swGorL5ifjDrLAvohCzISEi5zIppv+dWqkz0SWJ8FBj63MFBo+Ehs4ctd+FwGkz0HeL9OIKH4PkZ
mr/GMx6fPaVC1smx7ArSNZwIxIdcRGwmxgjGkLDV1IOuf/2gtII0/KSh853nfg5b0yGKSmOZo/Lz
Oz/dIXT18z+i/riGESukkjgZWpLgufIjv9QSCNjJOgY1y0MYfpCusTffauBlf3g89QzQXEXuFDMl
hXjVPj0/ukLUFBoc+dVAncSOb0wkMel1w6mxx0M14rzFdEALeCFojYOmRMIOBzeOYBsx9J8iNX9q
lPSkbeoWVxE0BWgeBYdpFh5wkotfeL6EY0XQWyYG5RwLm55yOK4SFK2xaF4d7D0W27fIzrV3xZaH
g5suoos8bIQfxlvwAM/WZPsSPLE9uQ8WrjoI4IKJzfSMrQ8Ft4eu39i/56hE7cHprN0kwuoalxZc
xIM5I5vC7SQRR9D6wGEqZAkgxiclnKiZm/x2Pimvgr3bZctgfLtZEUeqNGHeT8YcbwzOkQIupDof
qAK0PiWVUy93WRs6KL2Q6C2jceGrlBVUC33Tf/LG9xkOOmZpBO1+Z+tNWMu/zluqwHpblqUXn51m
LfyfdYI3HlF2d9uIJVK0MI0VVq6jnonTxD6pynDZ3Pdpz/cBoNVGAGga96nIQS0H5BltTCN/VZ4+
DKadctqeBp4s07/3mf+Co9+/lScRJZYCZ7ftWKB+z/rLeGP+0SBWMAWY5CHaRYD+dSTM6dsZwXWI
2G3OyN7lkPw4nTnD089K7AqHjEGwxCJYjcKgMz7npkFH1VXowg6LSbVyvM3LFKjIxoI4Fzve7mUb
It1q5ZEjS39kJF0VfUcX3kKVjfxR7EyHi9hu0yhitAmUrcfmqeFZ3bjIl4s27jkUyvzcNapeR1e4
CMvcT7bH2ueEw+mq5PrWy8fsbKNGq1IFIrb046pCZDPJcXj2gOzvUP3zi2Bs/w4OvkxrpBvmfqZj
e+lY5cv6om17xbrOt2NbdIwIr3vP7ZpgiW4Qbz+r35YiyeMIUe1sSEXkXxvmpH0H8TfEMZ/pNE+V
Nt+SLO62vli2F/7R5EUB1SznOig0Hd+TYdH4N+bh9guYng6hMBp6MGE/dzQvGY5gJdDV3YDf8+8y
qnVGJfwWqV2VC+FKU3bRE7C74pAV18abc+x2CJMsnuF2vOXqM8w+gJlChCRMASWzW0kA2JUA8fKQ
IxgJ7yWJy5cifeXh/ToBtzF/GDDFKMCUGHKlyPD8aIUn7jah8hZOOzOSH3EyVeYvkEqLX5LQO+Bj
1mCjKz2TtAYZ9IDXtzYMtfdo8nX5iEW8HVpcMbLyBvBZdcLGRo9/oG5oDH2UmhTanu1pW3Pm0BxS
VE/HcTQV5SJGvGpI1XdkH68TtDl4Ysh6j29Y+nBOVUcxpz7Td3MFP/wGqUwaPfuOt9DfgCWyCAqG
pmGSVd3BPLMwSjtXDrUPge2fBGc0QqvlFIQ2LZT+pu+NqXExSuMR3Z7+blv4SkjTLdk5lKeJi9yD
39jNQQ2NaNpxHUkmF2ko7bokUGj8/tCuOcgpA2gBwc7q0VC6hU8zZuvDn3Z4K7PG25BQJhOboW0N
ekgkGWtT/eb0LNseagH9ggWUEzUe2rWw9BqxwRENZc9dM7H4hxZab6ct+DmImYvDOq+XCsW2mC2j
h9htiGSLvMWZHpwQOgnK+B3jYK3ezhB6vvfW6N7OuKcL+nUY4cACgXUKNPZak8D16MjlS6FVni9l
s9ncla0m+qgvrt1X4FTLvX6OI1yEQZGKdFiPkk4oEEIdsiB6psn70SiksK+Iqg7ofV32UEEpYlTt
qjKNRcEeh1azKWohzuQub5WW8Cyk1abse9VtnesfF2tenjZB762yvDVHmxacr5pr7DINgV0R8fpM
rXsgSD+KkUmKEo2XcOv4ZRBARA/C7gsf1lUUTNLxTyHcAMxdecvqcZtKUKQe8Q90gy0DWIo+G8GL
WmCfsrMbbaeSSfwOmM6zA4DmerWpUPMtpNHVhgRhhcQEYTyi7Ueq3UOcQsSq7A4MEp6RNanGqdpW
HLp8ThJuALiXVy7KKx5Gx2blVX1EdQ119b189OvaInMmVE+xI1x1eq8EOjQKLk2NrHTapXoz+zg9
9tdHjJNA29c6xPolHaZEx1hiMm+VGSOFt4N7LdNhda2nUyj6kST79TRmbvN0/8PhC7HRZQ8ZLzjd
BQp5nXVJG7uMNeYtNvSRJgdFdlAoCIG4CmmmwPsKSsVIyMRF3J7iwHjxcHClHa5plibXjBuE1rep
9oFgNmTwXN0jhxmBhUF9zCgOOO2l6NCJvi68scevB119nM49pdzSKVulH0NeqsB8kLmHCA/fAWKg
EeAAkarHZbOnmqMbElD1f721JZYrZE/Mgo21WJn4qj7QJSG8DwnNzJ2u+gDA8HTou63BdjmR871R
sy5sWQP8k6r/PmnblhRnrlpaPJ8z8W1+XLVc399KToAI2vu3QOLMFGaiKmgzwdnKFX0QGgUzj15m
S0ig2tnoo2NjL3flSjmDC6zsVcA2KObyUxDGFWXF/4M5MlsSSq95tc7d+fNXsR3kJ9AOqXd+g5/k
s1FntzbGCufx4O++rGaxRrSJQqxTui7aP96tnPnigjy0c77UnCMDYDsl011UZbWYrv7GsV9LbkOh
CH/grID9bZy+M3a4cO8pQgI+jNY33WGBY7x5cLVMYFlLiOLigS47oN3HA8uSE5LWzpAJLG9hDq6L
aJTDMNDuOc4tXzybCSxfzlrrk01AdUqeSDief1/65b6hF6BrsrFhpwY4wUue6f9Gw5xZbnqsCBRf
0PRGm0GLIqjB+zRo3vWut8oGXFISdhs7Qx8c4jIUkzZosbM8cdlOVDXbDofbghPLOo/C+F2I+Own
LqBF3mJwREn43wZMkoMIRM8HrfwAvnNievfcn6pKhkjkljXFmgAmv5UubhZD6t72wfxhyGxQPGm+
uWLnkEKtj2DuTVVqdLTvKAVbcJoI7OdT4m/JzzfccrwmrVJH08Y/snMmZn2i5+ngzI5+zOTcEJln
S+T/lCAI6BeQBD3NTv/AypYstvSjwEsMxuPG7pibfYTq93TbSrvEs8VjTdE4SkufiGCkEAFhz4Hg
fi5mph4c8XA6d9KE2fffBCYFgv3eTXATEcbE7kUukw8xwC1S8ijEL/Dos5vwj/56+gIHEbhwDW+V
3EnIC3sSekh6jumiH7gd7yS0GUCa+vvCN6ZrtmeesuAFoVEGwZ2VJECoNLkXUCKXfTzvIG21pRse
jby61F2MSIz9Hq4eyV8/TtSeVbcIjpjL5q+N25SOlqOTrx4DnMdbthn0Gvu3K3tdluz5XV5QIhl4
DCsG3fSi9gqzULjdm6uw+KjHoN+irTAO9+KWnNmpeK61BJmcBKYCyY9w9ceN6F3vPogHHus/P+u/
nTQ0nmRB8rX7Jbcva7DE7xw1rR1w8C1bfRCJoKao/SsB++jRDB6Uz1BwHA0ASJ/WrJj+57Siyend
3SoTq3dKamPE3WyG1yPFeRhJuA5Epd0KsSg+z7qekPEklGWUd/inMer9B1zOKt4nDUhYdHKzpxYL
/H8zLH8YDUxAdRgQd9UH6bTtW38jjxDAg55Z57yJ2Xne8c6ziWEL58Z7zMOdEAWbKG4hAEMWlhrC
sRgX6lE68GaLPZ2ZpXMmqxeYF3/RzKJD/MpwCVG4KV+gfqknUYBoN4ZFRFxHNziQZWLCB9d03FXs
n/hdDuT6iGEbyBHENR5MPKdkLgip9piijyOne1yhbffWVh/CIStVOa9kXWQJ/BKFC3Y+EL2C/c0b
P9tw9x4q3to1lYLIApULZvPOiozsrLQtnOzOQix1MIceAsjQ5K1CHQqY+UYvWAU82IhDfLxTWSPt
kH3MHertvDeO/R+MiqDYlXqz/JrrPpEYcfHVzc02UtmRTArqxzD1q73n9/+o1bfGUVLzyt6MjskI
GyULsDEc6/NFItTkeVqG+xom9l1IL/1n2WZr5/BHyfI/uFW2gxaiLZArhbeMY1455gWRizFele0i
YXBqR2D/kYy0sAWEUdbFQhOvEcB8Z79tr5AKFAknr+NexUt/PnwIYopUPRcIz8MlQwVmyo+ZXCnF
yWfjBpJhvv3kdA2q9tin12vMp3/bQjKxaczH9287pP2RXKNqSVGtS6jk+MdsLbpZFOvBp6ZU7HRn
aN6QXCrnjQ4/ZTYgwX8yMUNovr3sSl+PNk682jA+wdRrMNqL8rt7YzRiQ3F50ANLUkcGKKjiaQQc
Cm1kx8nSI8NMxRn/ClAHgrS2W3zQP88Uluz7eF8ezzUvRvF5araBd1ICtv1mV48FdvVOsW7nf+QN
VwOicno7P+oS9QYsA84gMN2I6dMLXsegZjfF/mxFMhaU5+K+F4Un8kgvubpBpbg97odN/PAk12l+
FMHgmJkbEOP6ZS3AdQfsUZh3zx5hmqMkYWZhym2o2mtUizl6sAY7MBGCQspuBgBunD0qSEc5GwT8
oeZmlmjwvpymb16z/0+wfnuNiCDKXPIrUwCXcc8TiLD1pmN+YMWGKlddHYz+f8h4Dci2c2/HhTdk
kM1lLWEaJMpjVeRFL5VJsBrZvsoUYuos8U+TLlUQ/SAXW7t9MtTpFMljxH7Lg11g2lyB2cWtv3dX
UBeNMc6f6LGBr4wh4EheB1mo9uCcpqaimg8W2f+4FyJjaR/BlgU794gs9vwwDT1vXKvqCKuQO9Kh
q4WXzRESvQRYSBdPl4Uk9ZUXyAilD0z6Ve8JoKN5o2nZmYJvMPq8ZBjL77jHA0k+46n7GzOEwIuS
qxN8CkJiJI6jONHNj5oSty6lmQC64hkEGV85ZTeMS1JHY4UWxqERpQRshHU7gBfuFDQUtz7Qmsxl
KNdv8GKL9XfWU6bvE3YIpqHSw/XkCNk0lbAivnKj5hXwBNsqRAOUuNFdPw83XhCxDiCb1yoTrHPF
9cDbNv7D2SJ6wBWpbzVZZkW17VT34S020fLUJm4Nz3tC8sX/MEVJqODLa9p1TSXCD3TqxOwdaSC4
wHso1aBU6bakuzym3LFkUrVNEdrJEgu9yCxkFFOsQOE1MV/LEQDU3TmzLE1qleAJyQ/7ZavWrG37
2sd/Y9iIHv2dRlzx+TJR47qBYeAXQXxB2NPWWMo3BXk4Tl1TtEMFOLdykj1mZbs7yZx5qYT0YMyg
QdYxGHlTrMQmMaYuYdJtLdpnhptSjY++z3hKEmqZURSpJkL0erWxeGEuHGbVIDWIM79aVleUIYNI
Eb5d08mX1T4jFMEc9/Fzk2HCdHjO3PkIu6FFRiDOLSppkjPdinUk6v7rDgKQiYDiR/Pw4/m+8rXI
zlj4J/TpiinbtPMmmnwSF7H/1T6E0oTDicjLmlGGad3QZkpF+pdbYLk6p9W/38Kr2hmt/INpIPG7
wqXScHHpWIryME/YJfB80P46d+O1DkY5KIMyZZWUQPEu+tA4AjhNOylNjR+fLTTts0gpmfLcpwZL
+LbOTMCTxpq6A5Wao7DAbgFGH2AZtU+dSy5hU9mNv/dFKQ0PvNHjgNDz8tQIfS/B3b40acOGMgHd
8DHpWIqHjwhDzTN3IYkOu8bl7ZxOzFNYqV7axMi8WtfpuZ2O8yHzGVW06G50FseGpOjFHNnHyUfc
6Is0Y4/jzFE961CO9RWWdsf/SL86tgFDooCSjicXqFJyZSu1lf9L6A50iFJRP9ogo67LkUSV6+qy
G/jO32pJ3o+BJ9bEQjHHjubK0hFUYhrF8qrv6lzF/s6p4mhw6OLJcFsU3hkgdRV3B6/TBhmdBfWY
V1XGV5621Zq0ZAtY/ts2K6yZea9E69/rc4n9gUjlXhb+01XU43I8fETscQvgS+jP5c8OeGYgPCPp
b0gwyaT8SJR84HQ3oq4PRYiKtNO4nfjw3+aLftXHLZ0I/Iz3SpwuTCjUEn/HplkF5dKwVKbvdkTa
H8oasDnIuhyPZ9MT5YGzPl7lJ2YJlbVqrJPWBvqYiDhaiZe4xLvd2sAAD+5KUShALteI9iGpGXkY
gQf1M0ILjY5tBNO2UgGTEv5zCkzB1h09e1OFu5NW9137KXaOARQxz52t4jitFGP0U9ULGeTemle1
trtAyBXk0MtVc9NGpamdNmkv+JK/Z6sw9o+4u5lvGk1ifcKWr6tK4wJcBeMsWLCartZeNpMCUBvH
6He0Jjhm9jB7tFsC3EnEOjeQn4jhZGPOOX12vIOG+LE1YV/XxspRwYIYnF8WG8NO+YlxgJXPjY8R
uwMZ0f2/7N1DywKmFCXm3HVEbe1nNoJDEnfksMZ9n2RJj4StxplLot1J4EoFd7Ru4Macw6OLMVfm
R5vh8Y4uLci3C60L6EyksqYeh0urxJ99qTee1I2v7H0LAgcAZ6aLEM9gmGECVvbKoYJAEaV0LyCb
edBq8IM7EL1z7biZuBw+fUEfYOChSsx4XCMGy76VfWL6eoH7zv+RcY73DO8W56tWZ2z3i6gFOcqX
hEQVf69ZhYbLR+lHOjozDALRicnOXQx2Lqup0AIardA5LvWv+ZOEFKurV2cndcMCYzlGiBO7xKvi
enqKsuAQuIH+PIW94CgxJaysz9nrZmwTEi3pvkjESmeMtRnrw14JFm2nFH37SVpCmDdOyn/emWFH
M+3gVOKYI851MOwoiVj+YZu2J+EhjlMhX7l2RBW88Hw+WXW6bFGRDQWo1j4qzZfBIVqDcT+M84mY
t1yZrfKu1g5N1r0fx4FTuY7ZXUcf9Q38Fh15IeAKPj9xvB/2PwQ1aY1Nx2WW/8JW+I0WgsvLN3Zm
CK2/bOb6W3Zte2NwrST95xHESs3mL5yiNymHnBdQRWkCnZvsOsh9Q6Pych41us/4x30Q6CQQ6JG1
JQbtoDFo7yG0KAsaf8Ztic+tJ8XHrFa+VaUZFHXofGcOsWBUcq/X3lDaD2AjF4JXWd/p6XbS4q04
LVAJ+8B8kt7CZ4arzyyNGihC32cFqzLCL3WIzqxVkLwL1XdFp/zu6dCdNqrI+N7+2zdB7NYh9j23
zNTXOrgN6KThfA6dcuuOgraZSphpM22g4RzL3MqNnOrc85EkEoJQhDjguotCosvMMKgiy/FkvqME
2eclIkoN3mi23uD7apIfbqmeE++qNHQ7CsDQXWDcG9cUb/H5hR6v0RIqOZ6gb0WBzfQRrM928CJ6
+QaNLEgZJ0qjb1i41LKnt2IjtFnAFoR2pmd0ULHXaxvYv4f6mRjLqIanngkNHmKTifendvI4AP/8
TZSwjlU9KNtLmW9jZPUa7xjHamivEc+BZgM+enOExpoBh9g8A+SDifvLSB2VgRRBYFT+epCPiqgN
8ZrpF2nEze/5iegO3Qif7qjBD0FuUbJhCKS0HSZkc4+uDLdZUbSuhbXPL7yQfHmpACMeP9zvIdzW
Zm5gGL/w5DnBLrL3jjlgkA570cIpADOOBg9YkDDo6dueGJqXJZWDDtPVYH93K8BOpwOhtM2wGkq5
JidhqPxl65Ebnalr/a/Jb2t3KDexxJre2IbzHMImOuGMyZTl2kKvsEWy/FwpdCL9sj2q9/p2qO48
3DAuSoqnijvzLDXci257sYClVgwJK6k1PpGrZiHz2mcy3eLEhZtrbABOa34ceEy+i/mM6f42EE+Z
95+hXcRNUAfG4SewoUEJan6Go1GqFqIJh7/rqGDvPauOX3EPSQc8VAtd0xKQql3lOfne79PEpDXY
EWX9ixXqTiIIBcfXQD11HOZhXdC1LqQvigBtFpuADAwtQRA6m6aTOEnAOUjp15tuABCRTJM3W6nd
Y2nI0jFmgurFmf2mSzycp8DnHFAC9imqXvia3ij5ZBXQv6z2yupHfiflGhaQlxHHHe4+cIkvm5tc
nb+Gtmj33PuXAL1OwgBLbI0C33jtS8/Sr3akjc/3zKZqOoKDP+k551q5O9jN0Vxqwlb6s+oRVEXv
dCuq2LYZfnnIuxfsYUaCB9JepkgGtL38TH8pC84DvpjRjc0FLC4CDyO0pWTwQGLNFjhaeyOHkRaP
XzN+UkP8cAZS19/bTxudWcYpdaA47fPsBe9/q+x/djToh0nWndpwwtxOE++GbKOp8vwU26L3oNU5
75z4SCevtzsAK74ctb2SzC0egkfr+SG9CgH/zQR+SU8Xbl5+UiF6IBhP1WDi3fanF3+Iqly4nBOQ
SkRaWOtnVh7lyZMp9ZURJ1q6DhZeaU5/U+uboc3bvvEm1m6NByh7uZYMx38fhmft6y6YefUCN7lx
Qfd+zCLUssXTcikMk5oWydSPZaO1SfzZBiN9dPh41Efj5BwG/GadpGUhrjPJ0GQjOwGwc8GpEYdZ
JliglGXozEkzu7SCw6EQUby/H4znky5fD9sERLdX7ey4Fi3Fo463WFzVZ6TJmhs7VrpU26w/Aly/
ytFl6TZf9pFMJ0TqNCDMysKcztopNlA1LM6lEITkuPrrbg0x7kikQRCe58q5Bc1jZs7lqSpordCY
18xovvJ10hO0I1YGNjI1sa65Law+XIxEA8H1N3oW40ZKpdg9DUkJsRtoEWmM1NjtcVmvNg6SW1la
v/4ISPKqINgQgFi7hi2a3hNtfcVeEa5fJD3vgJI7U6UL04kTb8gtF6t1i1wjiuRAQf6v8i16AiLS
yRGS9In5GpPF8UQMJodrVtiW+7xRGINiTK7blHimbnVHJZZ8s+H2Q1nQ2rY51Pq+hvZpHn4S4hNH
zEHR5UkyJuieKhGotLbGQ9rO63BuivObS7hrFEYRYJ4ZjbKqlOsu/AFcaA+zZMyUwPMDv2jG1GaT
6ze1LA72bNweYrBhXNd8HGTnJJkzkYORp5jtgvQFoj4/2EkKE5EfXEFtfE5UAX7mUPhoOqQCAM0r
rmJtMyomLwdp4r0fSDaiHVx9OcukQmIEEm9CD216mgcRJi8dG07V3Q0sP7eUDfzhIr5MnvEMmnx3
ZBEuAeB4XWcZ4f+uaynPi0K4j0YjT7ZfJuYnDFgCX7VCPy7P4zvrpwzHZN0fxag9+OfKmN24VAHq
jThj5J9NAkFGbOeeaMvxptAV4tW4AmwubnRra+jagJem6d6YG47RYU2DV1a7JlaGIjvWMI/T4erP
E6fYA3E4wGPlHUhUCvXiojDrtaytdiaBLER87sdTAZaqG6vNJdlpKfPwpiV4nkTpjXJHnNtFCHnc
0G0RtyhLT3BY7olnozt6g8fZ7G7XBKAhf2rZkOKCoTi3SptVgbfGeD+ltcl7/VmFMDM6I98iZdZ9
DZ48zB8z4QQborRfV4myjbICffXfOWzeUOWL9VMUyjcnNtEMtHJGlTuxA9oJ2v6NikpQ4RrU6MuT
06PQ/BxGkhYHAfY41lTFF6M6UJ2H3vRleRhZMGPL4jiOuhei819oDN21j5xLZlQdjLPx6YljevNF
xSJMA4fLk4lQMBk4MCwuTng+2lRoIcFV6neZhsf+HWDNmzzUqiNOfM8Oc4DZvNh3IPypyDqi5jeN
llyr92xJamteJn4O1DVYjKLxAiBSHlG2nJv2xTW+b3Zd+iCMIMmzIO+a44+t3ZiNlFu6UtB9jooC
Ehibxj2NYMgOatWm9b2Jw/TcUpK1j/Y9de00CEVHGN16dpMuyGSLH189s7kpBSTGdPIplrMnVGvR
RFRYvl6BiqQKXpaiiAEUOI0N/+RgCJ45i9ljKBahQe20J80AFn/SngAga8Fy/44Nmb/izhjKnPI9
HP3YfhnTKdyOEfyl9HCZy2iOm7onNr9cn9G5LDWAmOsOeoVU3sYSZONz8GchuchOJ8wndUF1b26y
sMoKut6s9+Kjz7Ma9CpV6KVDw2Yp0EHt9LLLpRwG5kdorkL7Kl3Hy8lcBOsN1ct6CD2W4ucTIvW/
c0KXJ9kaz24y/2OQ/aMZx3/ToJvyeGwwZh/3fyS+lwpr+KBIIz8pxmmwg4Oxhgp3ypCXrtXzmT34
RR6ZqdupK57PlQ8M1c6cQ3BHLWWu59zwGW3C+11J4yX7yRyNQWdYw4ZI/xpqhGQjMT4pN8Ct4SxM
7YT9rIiMC3U+Ki1w4I+exRADpe/9X5nAHoJU53+anr7UZFWfjNk/w2tSn64Vl399pRjxhswV9akD
0+QVg7K7qxzhCgtC7ZnOLLWgVhG4fs263IEbPj3AIRq9/pFmJo9vIGpvahK9B1O0McxYMuBU4UEF
QAb9vbDzT7X0wJXsXbvN1JBHF6ojOfotOBNvVEqOmSLPMV3keaLllf3Igleg3bQ8ZMN4XrBAhxPI
CgQKw1FLNeufR0FaNLWqwmdQWQB6aaPTPM0qVzLO7m0uTbO2DO9uFro6gfWOj4u1SXeEdqn7/lub
yqBw/xE3nUgBt/U+rnLLngbD7ri2yabPKZvynkPEPBTzEtc2Sz+ngtBSZqxMuhl4P4vzR3QqtMYG
vmNhKUfKxhyTZeRswzMVmBWHcJqSZufCZWj7/jbr/i8TnR1Wq5rXlz1GhI4UL7ej82sWt/OaFvJk
p7+kEBXrZZdE0aqEqtpvzMfm5Z/8IL413uwsJGLuxeDkmjw7y4xe5nZj3BEWNp6cbhfBufRtiTlX
JYs8VGOptvT8Lw2mJQzWGsekFNM5DpvegTCBlvOVMPO5PyKdt5uoUWT8VbNCcUWo0zTAckW18Q3k
/LB61lrK/cdL3IxnDO/jkCeTs54ZUzzQ/qxjpau5a7J23WOX8UXEam01yHUtpweGuK/43kZ7tqiM
eu7AcS9e/gm08KQm5uNIFt4UkCkR9Wgtntke+pFBhYdQDa0o97VvLLX0TvdxbVLBo/1fjfgrNjUE
X/yttn1Meji+WS3Bs09uSL8mB8ldCVd2wZcN7p52RMBWx4td+463uJzEGjKPmKcLjnfChIDq+74v
24djeueCggrq/u3zHPltYRk8QkZUC7RpRiKhvAIO8fujQ8LxdzKNPk02T9vYA6R4ZeXJo4Ht1sQw
YYCzm0X8r6gehmJJfdK0DG1bpMBn9i5nnc7MTLoS/ucJAv/fKHxmxKXEGO8kec79PWTPksizq1hb
D82ndXyv3inDHYJp5TFWypCqmv+MyBku03vtkzvj/SMvJrxDA9B1sAc+QgUxnFI+RjM2GdC19nWc
pT+2B7jvRCxyUDN3jrNYWZN0S5E5QAInMaJIUQEXvBtn6peTkG8U2JVhbToQUOGyajRE3kk8BxHh
ru/T8FXzttNhoBFvSehVPKZg8bsgDEsTtVP+041Lt38VE6SDvYMdMyAKb7TvXUX1533luKLRhqlO
fsQofNxvDx8z+2ekmwLZXvYyglWYGlBzueGShXDWS5GdWksfzo8LMlr9MX1Fb8vvyja8gv7gQsQe
4mI/2TUROmp8UkdNK7eazgxLv0iDf6VrWwY0kFaKafKgNUDDG5xlog7WSih9K/nxTWMqNCvlao9U
dbXIPlNiUrHdxH4jxPxKYPcMHwTXOEQjRgowDFQVDInLWnfiXddh5qymrJ7y4pGFGGyCufzp7ltB
SQ/Kp/FY9USXAATwfCkCj3BdLsk3rt/Iaem137Jk0fwfL0tikVPWmipgaXjo0Grro0/4xZ/0JMVn
jVZOADk/06DAry4eXeWeebpcSF3trTwdOHIuJwM4FtgTU7hdsBGnK4dnNm0qLwFTMNGEq9Yk30UT
u+o0ytk8alhlX+8oYY+A68Qc2/P8i+ph83F56SpRqcPB4H2UrhyR5xc3oztVKa+1TvL/Gl3SGzzH
XAHqI2SKjTEGajFU5pPsBA1UuTIacx1S0ZUN6Y8XFNr7MmBXm0CuHBCaSnUgyxVptg+I3JzUnafu
tq/CGogbNIKZ/LbPZn6OGymt/nJeSDHxHXWZ40u3c89x3s09w1EaDPPfq44Vuxb2sMnNBBJV0y0Z
0ZODnVVSRA5Jle9+TiUnY8dV2YthRR9Hq0rCtWEQLbDiObE80hOVcWxX9P8+vq1DkUfR1yWlJYBT
Ew4DJxGdWfZhxLAmhFYumoTjqR7HuaG2Hq0eNx4drEFIinTWbfVrK3tRwIUQEORcKoVXFcR2fFlO
yr8x4hEAfbhUz25YptCFOvXu7AM7hc9o+zmcl6Ir+GbGCNXKrFYELnv+N6dgraupNi/9jwONGgO8
hQPaEGddcWBSwvFzXYuW7Si650cXCQ+L/4ABKFzF3UTsQzcIhjKun4x++IM7ywlzX48y6kPp2sdq
+XfsDOrm+Z2fsSNehalepdKGHasq55rZnL0TJBHQh2dfzYc0W6js8/m7QAiTTm5UW/3HtVun7+Gk
wf8/6uM653i710PqbpP9voe+GATi77ztKRMYzKi03adrMkiReL5TRy2Fn6OKjFUtzAWfkNJyYiWS
Da4q/XAXhDgtxQVeaen+upZTgpfKCDoJSW3cD6kh5nB+C0cfxEbb6sL8jdfvekjnEj9btrP1Ia9Z
LOHFRGJJzoOj0ru6MQDgSPNh6s135kjyzp/r1ovQ0hL+NXH5pwRCdtlJjiQltdoJTSbh6bFXOLTH
Uj492KZbYKg5qWSaclzHlS8uVF6RG5lJqddG/jZ4eJGuYElg+qRxXwLpB1/zzv2cPAdiq3O19LZS
l209Nak/lOQsm7OyZiVUEBrFEItPhm2AC5HDRaZZ8dGNdWvtvMEkCiexWc63KBkH7hiONMrOnRmV
7b1j5myh9YWUmnsAxWOvb2osKSuZiUG8ILH6KJePW34PXLb5duLfAbuEtWPjOuYcMs6RNVYiarpn
tCv6igUE/9O5dlAx4/Ud/RRLeXyyoT5DbUYEvLP7AHz2Lmh7A0JvsKeo7h4XCTFUtW2bQ7kKPlz8
x9ts8i7s2YTS2qqRHKWh0dMf6IqN7gW2S8V2pAooIixwnKLw+wxqtaZnGxMOHFqenkoemznLTfsv
qCncjZFsBv3j63Msdn3oP84sgP/4TPt8xK7f+9VeM/ZzlUjlQDlNY12WvqJuXNURZ6MTJmyUvw7G
6AoLo2l4+IqW/95PnUszwX9LYWKoxFcdbtEpGQi5P54i5IClGHwQQ2WDCskUUGzeoNr4uvobnlow
VUrwdHvAbTDc4MfqDBUiyo29sPtJDcbQSyPAX/K61mMcT3x8zfDtyMjv1GqtOOUHS/46ed0BSLOw
0FaywMfEenrlKvQq5v0DIuzvuxoURl+MwK5RL1+Jg/Q+DLPgYm/inYiWMWTfk2cXkeUfGCfgh2y6
RQ8/fiyBXchnoNVqoh9ZgHtywI4qih7l7iZzy4Jod3l4nlYhx5z9YMaEuz4tZRYcGM3h/5J5Otg1
RGKsksWmIE+0PKamf7kquRG8PU5oFTDJJEJFwpKu0qLAPpVULZYgGYFK+0LePwyOo8t/oOBkvAJx
DNAHSeKfIwHwASl0CAqinHHUqHX1TU+XtFM8E8czDAU+Sdm+w6fzXHCmJyjxR1ItaNk+QLL5PdTq
WRukcK9HYj7L1ZTKvLAtl52ojYhGIzE7UYhnmm7VWvE33FM4LtwqyXtsYp79GYf7w26jV2BKpvLo
BNkVGJHkcnmgHxsu86n9hYSPvf20fmMxMW0YmnYiRFQDIpvUKQWPff92PrrSzGtV10soHxiFuuJy
RIGjxbox+o63HNBhTCKjiu7MZEJWP5RLNoApCAn4esN5wAwplOt8/o+OoU51Ic6MLMz8zlF3bBO2
jS0Z+Z+H2Dx0QQ3CUjg6/HOzFbOsRnvWHVgJYfyBqgixpCHGSCsnjO46t+Lf+Js0nFHnP9Q1HNkw
xPxPo0F7GF5zhZ+J/FrMOGXcTnhbWTZnOplL1KImQBlndTJLO9g93YJqMfRVckSj2gWKd4sHCmwr
KLyFJKJJ5Phhvb9r8BWTEg1vxnzPQbfmBSHsEyXI7rmFgRNQScsrunj+sYRT2shfgg95jqKyQ8GG
H2VdX1PyYQnDFq+1uXxLNdX17u13YONErIcP1RP2SP6LVEhCEXEYPrXYLguc+4rF/TnmFVr5RO8j
moNQYSmcI/jve4oQko7EWiIpapinVr/IV2oPVa1fH2QjDDxHwFJCJD5jEsV7OfAK3NufycLE8Mcm
rvL1PMCuMGvid11s2mRbarPDTjeHsw9ubc3dPhQV7HjH8CKo6EmpMYt007Q1DentIgeTSHD4olmA
9eABGN558SAm4FsUQD+LfbFlNM+3BUxHwQRXmcvNipoprieDMYXB70W6ddDE16IKsKkPNDl6HwNd
KuA2fIqkmt2hmmbnj5HtajXQfRR2biNgD85oKEhXqIgX7i4Xwk1LWQ5PBA/LZpnt26RtLkziVO/W
CQ4iDPgdCZOHJ7N1Z839vmCBnXOQFsnxy9uTtszoGX7hgsrg2v/R08GOapmvha+Z3CBdkpvmt3Ht
t3ypRaQznn+ZHoUlvcxEkyBIklfSpE/g6M1SkRRWXhrUQxNTazQJYqR1GjKlKQDVwuP3UnzXVRmf
A8RAEQ9VSaBh43VuraT1zpJ6TlRCiI/Rqm+nRzu29mdmGUYQeplLrkhdpbzg4zjEhYmnJgNsOhG+
6rREgzuZNQ/ZuzSyEF7tt1BzL9WCM9j+y1euiamNj+PxPervRdFKtBmiLuN0/ZXtNAWyR/EdN34X
fpRF5+sTArz+VsB/7XkHdMNzRVaDf4E5ChEdDfb6UaBcNy1dOvwBpxWxWvNn2uit2Wuf0UUcLar7
+51HGGFJkNVnhn5lyLFr0JbfMIrekVn62JVFDbH+Ht5ByKLVB2vuYmpH4DbG7s0X8HWrk+3e4V+p
XtfyBc+TjV7dxLMJ47bnvgXNywtz+BuKgc7bVfoEdJ1CDMX714kSETAM+zzG280AIxLeZ7Ehv7Xz
qkF72+cPXAn4TB6AM39W9Fj/+fJC5+maprWjcd7z1I4w1FcykoMVEzIF9w4a4iZHrBiZYlRDolvz
cmW8ijsgCeiZ0F42OCiSMJmhVhF9WggsXmZzoSreTroGuft/9B1sCGHchxtuq0UCAaZBOJctPiky
k/HGGKRTOosAa8s7BmyJZW1pLq/qYuNO1oZq4lu57wJgwowtpkAYbdIn/PyLKnJUFSOMqUtfkQP0
/Dw3Zq7Ht5rZckU1WXBt3vrcFH94zNYay/kKbKXXX3jPFJGfRSPsC0roBY7GVmC0/0QhhJC6DJ5j
vqKq9A+qek/A5S+X5Z6IN0BtysjlqnwFcRCKF/6boNRA3g04Dc3G+avu5+USwBJTO6Ml2mQvxZ/5
fKrYeq12ikqC/hBmtI16NZ2R94w/P8WcQTPiu7Jo6dSTYYWxUl63XdX06hy9xn7RnQ51NjhBOZd+
t/kO7EsBF+kLrcis2zqT+2crFEdm2SgdhiUsOMVGPXeYrR4/a2h8xbd9TTeiMETp4XtJesR2WzOI
QIOtoFDjKlZMmzMGwjxm+4vG+Xu8QLcCA8VPkDBe/XxKPl+kJUGOKZhGuzYYHGW02bFz2SB7zfQU
1o4WTTp5e8MnyJoTFY/jeL0n3sJUqmofxuGQr0bV66B7jpc4X3/o8By7DQ9pXXjS2Yn27o5YuQeb
CjC+ajHhy9Nf1ei0oAsLQsaWWLmBqrO6PCkqbpp/tYA2H5BMyX8+z3l0wlFqWyqWdIvSiNYJUcGs
XWQqT4CWS2A7SKEY4BBlbjmZmburQixc5J9u7OLrfqdQWNQ7UnZQOs+RMuphvHhP4VzoqZZLU7U6
jBr1bldivYJegGcq3TN1usKMRDM6PX6G3g2NxOdmLmY8PuZ6+qDLTlHBSevRnJmbzkfhTJer0zOU
ywySBWP7jB+ow10eTNA78wH31VvN8KZkl43Fl6aLO6rkzsEDjxbP3RwOWKKpcIi6YWl4/PB4bnPQ
WDwIEZ87/UEMB6Px48zombF+vaDjCQ/16B3GBN3DRyapO7s10VcNUGf5z5ytVRNihllWhctOTUun
Jx0ZrGVmHBgcpob51v1rrEy/JmHCQSuyScZc8x2bGfugVp5Sxb/iLOWOZRPQFOvAbbkbXIy3/lpN
t+ZpzDI6ece8dMsrCdv0J1Qb8x+d3KsTA+g9L6Dh9mWFSixOcORCvuMB2oRvHbFIHsjubKoHNNjc
o96LF6m1rGKqh/UGB3Cxnido/GFx+oF1yIpDcJPHRCIpwHiUjDIFfV29rw3tEGDwkGeAPMpAH/Q1
D4Fe59MLowrE6lxr9cirW/ly5oEHKfZaLEEHZ5Y5iG5opBjbE8ayZQE+IONP4hRY5YVnQewpRBJ8
7whABQu5qe88Z8tVW1P73O4Q+op8ObFmcjEbRTfI/qnVAotGuKUpYpWFLOk5GCdkXKcOi3k21hyg
XQYJScR/kpmso236X8Q3DEmifgtDUPQdgExZh1pAqkw4C6qIgsJ4RMHdMW70UURqeHiS77T93eWU
YSRZwfggeU+pDECO7a3XxGm4GxWCqzmcvTUxTzh6Q6XmU/uSNMUon1Jglexdcm9d84QXztsLYGEY
826keJ5rVmULPBSqoD18F4nMMqQEO58fipX/rcIWmKNoTOo4QFmti8vXD46JKZmaB/A2ObYVluU/
0EMYDVxpri8dLvQ83P8Gv6+5s8uKchImXmqbxEtOghNv/zZHP5PRr/46Eu3YedZottS4HhkYo3li
TG6FjsxUKWZQF1WCEJiMdrVwDkl3UEAU1nYBulrpswWZPqx3neKoAo4Tdvz4XMiBtIso3DvxfKhq
IqDEzxo46/Wt8vm7HAEfU9D+GzufPm1FmciRDPkTG10GU5Msr3gDfcH5vxWdc2Yo8iFS+b8vu46N
Y9H3mbJJZ6XUQVYhW66wZtIyx7/3cRtfR4k+BljpCQ/4BvSVvaRyV30ph+2HExgIMdBINgW/o9B7
7WkhMQkv3QVqx/cCIv4J1QOxSjFWBgNI3WZpPDDbfKibug4TdchTOCSCQOD5KajZg1qQdSUncUMC
WWs3TlZPyw66L62nIawnEJDUNNjrtHIn/WIj9+s6sDUoiczCtBcVL6CKWuvSNTIrQsbhcaZvejm5
OOH9GzyI3Ob05tH7AEc+bvatyducSJiH5i410pyLnGsmsiXSdg1fpwVdvS8OGbCv7dEnjF9MCr1u
sXGPkuCQV26lWV3CD/ETscfm7SzBKzkrH1fyRZTMOqUAxp08NrpxyFvMdpxfXYCxJZCaMJzWK8ph
h5F9/7AyikFZNT+dRuDCQ76ggjZS9DoIM7wnvAC1nvMsVl15y2MiHyo2jUUZoCZ5M511aZFjePhZ
VO+HkZ5K32Vog/78xEgbu3WyQysI7gIAKol1pQPcto+IMIlV1rPga9QVnahiOHcQYJkJhJA6zEj5
RZECMx2W73+Ems9EjLqEhwELeQTSookdcMOD++tVal5HW/qIL/luf+DqLViDvvS1fvZErjM1dfoT
h0WqJm1xkS/KtKg2V2rTDe8zI0ayAaAfz6ih6A81/swzRR/n4aFLdvWPrLXLtMstTggUrThoW1Tb
vHBHWqqMsKQiYT+XAYQzn8RCtFGrNI4YsnNdkxO7MiM7aMsYbHesy5lvuGJFXb/iDq9znf1cFhZ1
N/gur8yX3AO2bVixz84A0WBs/xBtzK7N8OoCiBXi+TRPsMO806FYwHX9t1Z+LQP21hrzVPD0Tuik
Y+7ggLpU8TB/O9d+QDkYxOyTtTcmo8JWDcGCejAfv7DN1Ft15qywcDDSmJlSz0qlAlH19VO3pkRU
60apr5eR2U2tDnk6z/SOgQwbrrj5eb/ttP8LjgfLIqkDpUpukwq1pwMU2Q7CxY7Y+mSIcBtz0EA3
qzNAoK70/w92/p+pQRCFGwa++eRGOgkFouq7XEwsF3dg3NViG+8l3PQ22LyZsY2ejUOY+eUZZEcV
/mvRXuY4NkgFN06hJRU88lOd7u+YBIqcAMXrZ6YalpVtRGpTVA+hH83NkjBA+KdHmxUzJjGHkk/C
NpXTyWXvO39AWa8bUz1NwMD2O3JmxPsGUSFEJqJnU3YfwwQeZgeYZhfPgproESfbVC8kMADTfw/N
3afARpnRQgcNaG7YLcl+N1Zkc2dTkKbzy11D0biH+GbkS4uZenDNA1HQwQXyVmokm51YQOurB3g4
ae9bGp7fhW/884XkEMPGlPs+0kN/RlJCr1UTOYlN/FOb/9viA52teE1Bl15SG5a/4/3GjZ0F3u4T
Adax6cfRbup4kdLFdQXCqXmaSVrmg33jxGHkJmQnH7fm40dSOFGkMAlwoqR5lNqKUNh0HC3Kaml5
ghwaVQRbniyuTm1BiQCaUodnvhq3szkcMkcjaR+/bNBv2lZJ+b+scrRKHKPCzKrLJqRUmVBjp0Ww
Xr6axcu1jTiEUThDF0omiOmvci1XkCc2AfVPUWAcE5pQ68ikDKVtsEqd0TyBCYyw/YykA0FNjEZO
aBBritpy2AObMxG4em3c0JhecrUvzi/53N3ilfCx7Y36gEor8zdNIoX3891YlvSFfaSX7BsYMlG+
PY6HtT8LQcPk4Wn5U0FhlBcyvKVvwIOnL+WSRk7rqtPuzKmTVK2E5e1mlfd+XqiGiXiT3yV8KmG+
PstGjzMxsJn7FpwBb9JjgKGZnDObx22NKecuHbmw2uvWEMpUpLFPX0r3OY9Tw7Eqdy62hUwqbCGx
tizdH8vMplCDp79Ox2mR2TPmH2mWOpAR3gEsWZg63ZzQGGCdJGS5xyL3cgBQ2rbqezkp8Pead8EZ
cWVMQDg5REuncJCIN8hlRu8rT30eMVA9Th1PRNotcXyLHjE0AgvzwtOOFJwqQ6JgWyEJ/g3boTk9
5CfzAom85f6kTvYbqPFGrwHBT+afNc+BVAa0tGYkGd8SVGHPAiQ8SB6qgISxKJurtX1qdUPzPoTo
CR3oZRPN//ukwOHNIVu9Q1CztKxnkEiHkxIWqcD3s702BmC0i3nLdKHRYyuxLuncGtUxFmwxePa7
ng+RxrAMVBCqor8NPlCKoRl7oz0J06Q+iYM1PTwskaABFhQw6+3iHnU+HDl3eEhuyMbdn7+bjU/d
tROD2KRqGdvGwrnkCuSQxjMDhXcSQXzdpfD5+s9Ks3wZKHlxNcyAvS5CSxUXjjG9seaHnKYyhYZY
VT2RLSnWd64UHBaZGa3wVeyrinM5u6ixT/W7qcxLBIUXHW2FaUjMiTb5f7CMPS2FzParJnNJhcv9
ayghBYl+6PG/sjfc3Va4XvV+L6NMsJU+03dfVJVmdrOMp963PeHPXB8X48WrUystqUjw6oD8ehzA
KNcWe64vpetayeYrDyc7UmCJYIqbg9TIgKoXUp+au0Hpb0kwbRLwW77+TxmfoGj+SIgsEM6KPv9B
IJWb+/JF/z43nFYX9wOoQEeoYvO21hbX0cA/zR8HCnMWJR3W/mPLD4EybOk/bTqiWybeK69hueeG
evgSbvvKMycruvx20IxCdeweTlHTyyQGkeg8O/8z/FkVUOgNI3hpBjxuCPSlVbE+bbbKQb7mqGFo
+bU4n8lEI67FeueHi5M6VjV7C+7Y2IyCkn47f7kmLVFBK3W9T4umPJF9W4FOUiCb/M9yyIhLgzQG
W2fZk4QoBk5bS+pzqEFNZ1+lnzHzKUJawmbw6g0D2SFm0SkvN5LJBenasKYgLz/aTbZRokFoRz0N
MWqiueAn/jybsD9i5rv5+9Da3FHebsdpXWGM1oNDfQ/1bWujHsKfjhKkQ9JwOqQko2eeU81h96VV
2PL8F9MJ+2dftV3fqchXCSmr/J2rWNm7dgOFth5ldmKH6qxFG+4rZ3GlgPzIAcA/4KBls3M2MaDU
6g/258fyfC1m/VZHy5QGVlrS7ZEqxTarnSHp2NPaq1mMvr/SJoCk1Tmgoabh3P2qIVGLdFkSfTPe
7Rg4hoNwFHwuQP1uvNTxTlk7vhHnX1FisQepLo+XS4ewaCWoLhLfBQpdbqLBjgP+G2WOM12Z/rjJ
lQ3NJW0fxFcXqNEuEl/5IOcTiRNGbrbily0iSiBw9q8aTdRIv51fhD3zZ3k1WZWO11Eqt4GjTR4t
wuVPUgA0nfWqgLvXW0Yy927SHfpnSJILZW6My38rCajLw3HzHTGWNBdq3pLnZUIbWVQLPAOsBXaR
Tx5OE6KdUvEMtVEo1wXpMFt6h70QAJZaPpfULuzSXR3Fr/ORjkOH0aUdhqT405IwlLnALidWcvCL
CjDDv/TOB93xAPZ6/wjeWsFLcpnXFDTsRXKHZoTaNeoluu8N9H5/tsZXo0fnV7yabGL9HhhSMgkT
CfamZM065aHqdMKaJ1oZqLc1rQw6/D7UgDe8RIkTnFhqZPKalR2WC7hJOo8md2Gm9d9eJAzwaorV
/nW28P4Kzu3mk0kGVburKfzT3/AawQNpoCXTqg1XmaUmDX9vQf/IR/ttNWrahNAGZEr9hY0aSd50
CxtroInVizDH0OdVHaH2xRXGZeFd15yai3UY+NLKfFmTh77SoQ9iN/lyTJ566VIR+GMhgMVY25l+
LyZDCPl6ouZAHnMRHmlDSjniXTQ6W4N+l5rDA3tJ8/bwcFqKM95Oybo0XSF4L9qtY8YkFzEtiIy5
xTCooYoJayNHHRi4qD0t0SIImBzV25erzeyXuJUPxkF+/QNm5NxH2Jst57z6bL6KypdhHVOcAsMC
cKdj0l3TUfOlTwclH0iW80ont7OYcHL8M2fCOsylFimeYX+SNXZMqYeSWXBrQ4ZAzR5n/rgsgs6U
cvOtA/37GLw8xl8Z0ggd91B/Of3l08v1szfN/N563LpeUqEYfFz1Qu1T2ekRdMHEjfO78ksUrkwa
78BGovl/gc9anYEwh4pYeIs6OKY14QxquzAHdIonfhfB2OpRiGIYn60Nz/8qqeFYsC/OFEwJb5bO
iG894fWzmvlDowtPwWxHkwtLYX/IcRBdowKkjgWGuyxB8SoxTAg5YYgnkUclI+WY+HCJLEwCNCi3
5UPJr9y4UZ5vtviRafE+CqXAiAbDR2dg63OYCwUfMg5DOwfFLOZq4o41ZGCmLQ9SL7Dfwjig+VGc
Cx7f4Vvvto66DuPZtdB4HpC1dJSC64oZ8lHB4/9ZFBVNKjEh3Caabw7mXRF1e2a9goZxEfGG768p
vY7UeEXmXp50Y27YANJ2X8EUJ//6AyybGJRmX3Fg6WbAXhzXn7+Y+FmI5z5xKKko1tR1P1Befepf
dIUwZYT+IF2jjB14yZssd6qTDDRQ5uptAZ39dPXqYuUTE1SBsBvYSwAaZsd+MFr6BRp6RklGsXEJ
Pl64KooRHMJ7/OpzkPfyLgLfGaLoH/sB/mWfCXIBdWYiEywfieaPz/ppwOt5pFZGNIqmO4qnc9Aj
e4vRQVIVBXuo6Tl+J3nLJjmimqbsOBMPp94qZqElMju33Bufw55rVuYxjbpXFhpXAlu04tbGfOWa
MDPS1bBM6vpQDKzUtw+ppst0ZlaohJS5MOhx931rXAFkYsvqnSf8jgyDta8zOqL9ug+3IC5CxeH4
2wHTNiSscEALZ6JPW8AbnNvxJW8HtmtKgPvvLg7AjBtYLr9tMfVr3Ne4ZDXBzIv2X8ScoaFcjTGR
jHgigoBu6GUYpVZCWRCnreKq78gKm1zQ705Guvm6dAJhZn1uvPo4ctQo633+fGizhHbRJLvqdTH/
wOCXy1+5qS7d6ahGLfNPGybbhKe11edsWSlvbpbc0XvQ+VGNmMkA9UMXJzgkJHEdxdhhphlP1ikE
8xK9kuzorWsEyBiCEFQ3vFRIKGt/Mb0ZrpraSd0fomYTCWpFu+fBzr/sdZMhbiJjhPt6B45vPWH8
sQJeez+X6N800XArGOmFjopHFnbS78C29aRmLeC0bfDESbQ5MxNUggsoynkRoemaYQKCoO8AcrHD
0O38qLfE/wS/StnEC2vPH10ciYUz0eKsWwZsL6ByFsYuqKCHN2Z9EpXcSx9aFk+TOcqivvU6+5mJ
gvpYp/5e4r7mn818hiFrlu4f3UDfho5SRnjz51l2ywM3lWmABX5qPRfMgW0qOHXystd2AuPYcObb
0HO6koqyOlYGet+MO4N0oss0xXUFviDQbhlSNuaYsbl+4fr/QLvpVAIYa5UttrPHh/hLJujFpe4d
hhA/71o69xyfI8hTBGfOCHKOZMyTvqjCRN3IvMqrRNT3t5Tgd++rkR94gZWvUH+t0CWKWJGuacNi
/MN9qEUENMDDF413jPjnf4fM02zcxZ4xdKQo+fO+cI1FVrY/vhTcmBIlOCpf/iDa8ZONJyzQTdbJ
m3hQDwgADxBnvbbbpUngfIzvz9SVY6F6dkBEkL1uDGAAR4ZfrW2hoS1t3/rgmIZsz1Towlncn6TQ
hxRkOE3SFcW/doOmTcF+ToKBrUnSe9DQigJWAfGlA3FM76sgFdMf/NShOErPvv5+EnRV2/FnayNy
sBHH+KxiBTAu/M9kR3aO8ELGcG31Jmty+P/3l3JP++njL3VOaTBTAYU8hlliMDq4X+6ue8ASlby+
WEMcAbqtz49WS/GcbgrJtzumGDaChiBYm2aMiWAmH7bSdPO8Od1OiFYUXGm//xYFZ1x31JWMi1d2
a9KKP6DwzncXnaSxA8EHRR2bbHsuyTKJiuqoIRTyFG1GEJTBUaITre1jboDH5exHPCNn7q2T35Qd
MSuS3eWeWERI7zt7wl61gPM5XXFaqaNdWDifyZ8k8AUcN/INgcLrPkanHW2wPDUw4uPVwoIWhQV6
+AGPHUSM4Rw/tA+rRBgK606FfGvgzkySXAIiTP39UCZLNZk1I67mTVWS92q349kAQGIIzWSy8xej
D4/xV+tdbvP5rOQVzRDbX3DPc+5sRBRk3Yg4B8u8SDlQDqxpusiedqQoBb4lx62EtvxibfVK2jlp
iEP//TFWNX9scw4Sp7nrcQb1zI31TANrq/GIW1LGEOWkFvSsKD8C0Q98IO5l1ifYj0FGLugMztqU
6XpYvK+SSsb3AtrPvOIe0bCp/5LZmS3QRg645kNjjCAVDC/MPhxPV7ClTfY0kSfvGD9Y2pFosVHZ
xHxoK2df7UanCbna0F9UCsLaeIF6R+GRGWD8lG0qopsXGZitkyHbeiHWtEch0rm2zaaT3oNk/Z2S
YuopmBM+2NuwHzPzIwjfuOD4qwtPW2ZFQnkRNSiV7IUkyPkRH9DsgDDQCsnTJS+mqwsWwnhqjcSw
O/s6tJcpt3OB4vBm/QXXz6TlcGagICmIB3wTmsKh24SSx8bX/7mpcLUBLo9DX6yp0nR4v/0kjJSH
meydwLEb1WR6zykR8BjIfXGw79eecC1im2uSrWy45soE5ouxNOz1wlnoPsu/YHrS9fENvj+vWEGC
j2Kkl9lsYTw+ZL3UWnjU4vaJM0zCiGiCLNUK+H3yy4dwS1bnFuTGIj68iR9+nNjFeFuLOSo5c02w
pxPOYV6921lVkusS61Jn7q5vQ/N9gD8I3+EO3DRzW4dAt8pPdgFUy62ySnFk8fbdx3cP2SIikPHN
IsbJALEbOLQ1u7iFCOsJTV5Bg8RpjhfOdgxuKrTBJIDnmM6ORhvOqcwoLnXxW1fDaqCwMb4SUL97
8lkvCgFypjHSw5bzfc5qE4QQ30OEmqRv0UnAtF37GX5Pg0jCv7CN4Di5ACIVh7RwItemR2wFFK+i
lo2bpsMh89Y/up/LUPKHKAlxuYz94msNP5Wk+sACu9SO82iJdqAyJ21PvTBChinUhkgMY/QLmiOF
Slub9t5KKWs/012Ut9enFN/f1+mXqDUhBP79Syu3xxPSpRgw71qBOBvOXmAqysVd3L9QzRKMW0RH
5o5q8C0CV66M6S3AB8hKm/OLL96caMhoLZDqV6fRaBN5bmSoegaA1wUUIb4FPGYzN/TQ5oImyE8p
cs76S+nUkkvizq/snsoqAnib0YNSmYCqZYCmB3vDr8v3nai6ZE/3FZua6RFULNgpobCwC+59CFc4
xOdmNpW3a/zgTuAhCYwXMJPm7+Ar3Ue4I31KqUJVjsLHzBcZCI/JbDoWkHMMdUhDjn+iWnzVyEaG
zaoeATY3hDj5WVTUPjK51AcSjVm0dXg/rG2qNGWWdKAybR+pIy5dy7NHp1oYkxDan60JSCgeCLM1
aiELAuZP/P/tyV7i4G7lHx9SnHmVoRlv/+tXlGMMzaKPWK5EO9EuHd2gAFMhWgwSupFYe7dM8npQ
J2Q1h348rTcpK1JM4j8von3kGZTGEle8pYC4O9PlABR+pEsRe4EoR79yHNc5q37Q9/GgO7RBhHTI
nN3S980n2lWxPP2gNZjqhPT5tvKmQAi++jbFuOAbhtBvHHE+mq9E2/4/4jpiup2/yaOPLvL9kEpw
sGHtjAcohjBu6xeFA9kgNCd4m1IuLz7SUYMyU8KFv4+sVHxMuF6njWcOCvZSfN9PYWQl5QlVyWTR
hmLzVj+ve0MpHHR4sbC+C6JfDhIBRC+GTPu3qgW2izcSE4SdvwngL+3E1x6aepP/C//MESgA+tgP
IlaLiB0eTkvL7buxXSlGLjggewuDcA9IHHJfwMQZ6iHEA2z71Ma1EGKLXAgsumaJvhbAKPAfsjXn
DtfcJPzaV0ciN9vBau+v0z0+aMl1zdXBO9yTSIFkA6KusMufpVv+Q6y+sW37L81bfSlv/Bllibk6
8l/PvfANKods6vfmPvw50u0HmYWnmsXVBZGxAgrAlDdFfdOce0OhFRsZ8HUEqmNmyiGMlC0Py4iU
rCqLHNH2y/Fv5pwaWMd4SgSWvC2DJQ/5krXNv/6sZy2zwQNtsWiPw49RnV1Q/pGNajn/Da2AncRQ
WCFPQ7tEkV5tmX9vW8vymM6xUSmagoeRVFWS5wTtiXcXQ3Uoz7NquJyhLVPx9vH41bXXZVakIrRp
VD5lB1HQyqlVVM4P55kNlvpl0wH3Zz/q1q3UB+p3Iu0GXt/zvhBkqukslUs+5C7fjgcdeNVWYPQd
euJNcaP2B5tbDaQhg84YfRReLANaQI1umpgGM5yw9vc57iY8dBfD0bT6qbfJYja6hIjzYxBdCe4W
5kA2ieNJ0E47cUFcKCgyl++FjGWtwqMRlh5yswwOaEdYHUufm9c7Emdz1RJr1v+MtCnZ4GsSUbaP
A7SoIByFMe+vUef49GlOCAXgXhbKofGOZCmbmZSDAScYBJqvLn22LtDNOMsXgzwuI1v222OMZt6/
1WOEckaXWPrCwSJfGJC0n1SAXGxzFTyel7j08/39aj9N3L0niyOwu3Nq6MMZYipQ5hZs12mMfVzX
0Kr6jdWZjc41XpQTJZXYZN0+FrGQw/r0BRTAKEJhu2ZOf8/vC535yOyBBwDgZf1DTMV3bbcGTjei
pyA+iiibcMxXC0mPOCZ8Azrre3mPxbjsHWQo8HKQFJ28p0X0oGurdLy+01muz+KhuVzWuHd2z3Y5
ZV8mSXhXHB5p0zkKZD6YgdKHFednFiedWrKATnQMLYbGu6kTS7FTDvTaCodbcT9EkbG4+kGRhc1C
BVwX1CN++ONATFZ7D52S6VRgtvKFOC7JcOavfAR4rvO0RU5Qde5Hw/8Xa/88wABCVxu8Dk8EoF0c
9jfShaxxvrF5vYvgLgAMH96tWpq8IEabGkpFUQaj7bUCY4H8zcSMwoCRZ0fQE5Oj7+ojxoIulAhE
KFiPTFGgDtpjr7jFQNZdZLh/l+Glf6JE79LZgzIzlwJYZ33fhYgyBZ2YRQ0DSjQ3aJTHfPnE/4Rk
rj882/7Dp105Ziw936WnrziXhtNqQ20b03LHsEYsgeI8VJFpzSjISrfslJYNg6wQH/tpYcAPchVx
R4jCP7xlr/bxxUnrtdToTYpbROxoR6QZkZoMDLkcyToFUAZPXZiAz2ats5v3xu+Lu0VvoU6u7SS+
a6gkrEw65hk7GfW0qmT1yR75U2Jtfx0vCAnB74ilCACHMoV1Du9vnJ0tjKqAhlGzkdlqZhe8ao4h
EF2LN4tq2lLMFRRpZ34eGDEK+MyB01bNC21WTI2ruNf+a+K0Q/gx7tjXhu5u1Mlr1f8ALKKvkQRv
EJjvcUHfnO3ZoQtBclniIb+XSEVhglU2ekeNYmSHcftGLCMMvTYHyjQPRx6fJ32buK9gcWNXnBWF
2iWR8wtw3X0qPj0U+nwZal55ZhdBwHfIqVP8jq8+8w7rV5swU+mJ8ASwIU87LrIPSuXSA2Id4W57
OfTxzebfsUP+xtw9JSX6GmGeO6PLiJ8MGY4Ed1nga418XkSH9sUHY1rX0uWIdsn5I5hFqGvMf0lz
TVYAIGim2MJgrUmlQMw7nsBCMwy9xsG+s9w3pYwhes/JvbYBk3BUaU+W+joXdTuesiLma3Nr30fm
VzRPF43S/sqJeMGMaqffHz4R1l7VN2EqSnnjgNw+v97b/5MBYQKc1YfOxJWXrLbsvxhoo+SNPJVz
pL7FUJKQT0kleVSJZgD4nYSnxKGXU0Ep4RCAFxFaPaD1H/478AvvipRmLHjYgs68RaYUAbrUmxza
vTEAuU/ciSoodkKubhn0dGU8gNtMJQrXi9jCVYW+FLabNr0gbUFG8pBwNMOrw/SaVnLGlCM7Zr9V
Xmqoj9Y7PztCc+x9+YFLREqKVCoTk6pApeAUl+nUpIwsedA5/8091jz7AC/sBrjjGAanVvunhb2b
kHSvEE6vdgJRSeGbTI3aBMdqQrEHI+r1YdYM756dypkXEsfmg+3yn5rp8MGdTgbtKLxU7RC5dQmY
5R/XVK1enChHwV/Om4LN8eKNiy1lm4ZTWIjyoNlAKLPMbLaV//i8/BrlxYJIQRRy2yZi1/8Qt38b
tp9y7li1J0P1+Nz2CknGQPcCo+xYxKT6NWv6fHDVA6kWCSDyoUtg5Kd2xDDP7r4RXUBW+CmCVhIA
E1J1BS6YHcSZkNArHMdvSfDj/jf/jbzWM1/8y4gM8eCHYQrmuZqOk5wDlmhu3fA9v6LzuDzLBOyz
QdVV0RBq1Mk0mzVybSm6NDrxuKIiEnpfiXvTgbXFV3aaDh3GWTKUcViTFen4c9q8gDpbkCaTTYL8
Cxd3rXkNzBLe6s7jM9CNfWN/qg7Vlo/lTD0+cFJDTJTrFd5e//yEcnfVWH7s5V0UI7/15k9IgvWw
/nQghKI0qjXMyFpl2k+fhrOxpbkNU7myoJHhax9Jw6O5SnZPqsvePOWO0p64t3dKdBzopHuQzS5f
UaJ5nQ0wYN+MR+yaivgZ7yPRCg9MB6oHOlP9nNxUqZKm19ldZnZYnL5l8nT8mNmdAd0YRbo82Jw2
BZfDQtfHp32N3N2zblyFAlD5DATYR3uFdgftHDi9dtHc/AOT2+c9U8g1TbwBdoDKtq+njFAPvevf
rGoRIMPj9xIkEOQ4VrB3i9B7r6qY3DD7xZj8bZ0rgtAO8UX2Vv9NjqLmbPz2srwI/prZP8M/A036
esG29QhcIWpeffd3bosEGG2S03ZrSvAagkg++WTbEoDiuBtjoAbYf4X3mJrSk7BLoSX/zUcoIbNZ
iCxx3aW1K0zp2QaflAB8xlXgT0GLQFW+aSP6b+gZId4KPeNxXDgKV/gzeVkVQziJXaefWzFtwpfO
iRTiwzJs83sWdKxoS4anXtuixDq3ilcyotlBmYEQnuz2mZSMLT2+AO9mjVRuJc6krjmLsE3dS8Jo
HP2lfra3lfrAaL/4Ysj+aUm9hNbcL6dqkzZfMtv1Jkjkx4d2HoR6VHRg+W6///wznpShn3/oWoYU
JDIO6GnKsuv39G0+N2/YDEUnqHK83vnPqx7B4zgk5rBo0SWiOVgTHg620XiBCwYrdhzQxSNduCZL
AHbjHTOZfDiYdnNiQ9z+vhkRUiZt53zLXNSMW4lDUsUZN7gM+wdoMq9LJAdtYdaSVEoMLc2LjEjh
9ylfYcYIdGmVccn1BPSCX6heM4hW0rOsEaXllwcrfZqfQhzAi8cR4OLC/hv4TMltLePzplWBzCVe
KRLP5puV8ca3hcM4cj84HohE47ulRS/MK+mkToQiKNQTzgvpsZUMgHEaNidDHyD6Y3nyaShc5n+B
sLHwtqbWu0oR6QSFGAyCPa7fBJngVcEgC8aSypXnoQnIvYTLbfKXh6FnPLlvyBtG7UF5j+IzM7ml
qAnownEqulvRgn4IFgvVSd561AjTiL+RH1j6UlwonioYHR9B9FkT1ERa5pX6M+ZOxgzl2f1aiCIJ
U3PGtxtZKyFAQisMOD+DW4UfklIrxuq3jrduVbsSLLNwIh/HHUqQEJtBtlE3QN8t78dfq2VCVxhI
xjqiVpx2Kaw2dwg2FsRVF2f1SxvvsWP5WYj6qAqicjT2/wrh9OcvZEMSnSkBBkpp5/dG6CWlI9MJ
JslcDNBJmGC3GHQZFc15gKhCvdC9jxvD/o42ylRLLREvxKn9JR+VPreBHbUJ1hWxPjEnglPOFTL0
0PwyDIVl3rY55HkTDuMDVsX5az5ZbFUXN7oE23FT7HWdqQCBkdYDkqya0Eu2sbw1nO41nwTy5Gse
9oxrdoXikjHudCtaYkwig53T9XwGbFSDhirJZ1TozTkRf2Nq1jnLDH3JljADNYA6/oA28af5IawO
Bj25LVM6zgU1Re9Tgo0ZO+16XEM0Ls8lTarUg6bRIsyh8ssDONB6ZsGEyELlRo5zaMWxDT4ajLca
HNzkX1WfJDZseW6gFU3w6wFu/jHESHlgH0cDUFSYhv3/rJyROYJfRfoe6YNp9NjTFaknGuKqFBki
tItUA3lPC8FVT5gghURinmzaAupkSxRR/zxiD94dCkohbfO5xybHqJjdhvxT2MeHJrmuvSIxytDf
b5r3d0pJ+/ZzUtc14D+C6whN3/4HZzHYWgN5AUjFFa2jR3VY10Gn423fEp3RtLaHx8gPTTjW+r37
64k6+AJDF8TDsdTRvSqlTZia3viiqR4YBjY4HqgbBBTD+gVU/5BziXscnCOL9PvEVRPOB58Ai/ss
+UYgNuhFrS4AIZQ0XEJ5FpkP8jPqaSUCwHzIdBg5GsloZweecUGoYlNOiL28yxJZLWAOVW+XyMya
FBXSc1CdseznS8dmfKPJ5jot0JiChdEOqpN3w/HPwkQLikG5CCKDFhnR+JSraOg3g+z9tstOIFC4
niiyYh+iLx/IEItWbTcE1e6ygw7C9SUNa1l7BkDn76Q0/M+hwfa8WUkUlUj1uhNPE+I48alEHLA2
OO1T6fyzxuBALjgbPBRS43Qz/tqI+ohGrZl90rdATy8L2JMdlUPd79NCvJ0+bjqTwaCtSP727hKi
/7Mv4JLYTZLKZME0h1K2uyKu/TeS8jBOvKjQqSQ5dUsfADtjgblMXzqWb+JHy0WLSYydv/XANk1U
KPNl7skjvDH6UrXDVx9eYsCU/0JZ2dIiyNiQzuh6D4Ih0vx4v4wJtfNLU2XCOnO5YU+5IrjQ40KE
nfvzj4clZBz69u79H0hWOYDPOyF/CLsi8lKryCyDI8vmD7crffQZpHvB9qA5FnkrJtbzutm9uqbn
B/2rrpmEZ+1DZcOsI3D7K249LRqXCZ5nHg8MRFdP85OzhUIJVYnUN8JXQ+ptxZV3AZjx7xMElDxR
ttGhIwnWiXXExTk8a9Z+9E8mpUDIA47fxrhBcMKsZamvmwQ4zs8ZtXYMTO8XYeTF3HvaDFnuThk4
JGcJA/K/cx3GW8BnBl0NmsAFxW7W0xHE1a9Rye56yvQlnyg19Poh7tYtvI9rDofR9YlayXd9/98W
v/97K8ALygyau9+BUMiK9lAdsWhsdQUOcX07n+OKMEW5YRdH08Cw7zAea44RpPbLMk6quJh4083r
rtsZ5koMv/1lfOp4x7y5ci1/WYvS3qgRmTeDftHptJmVT86ebEqFXsWrMz1FtouPZVUzw9QTILdr
xJ+HD1/+qs096jKtVpwP+gPgv89MonVlJALan85R6vRIGuKMBzcWdMe6vbcwtAoLVZCH+lpsW5Mb
N5r93Wmz8LnUZxbJjZvbtJH1LfMLVOUw8xFUqOeEUDDG9k771I9GT43rDI45DlSwuBSgThka4NGv
dAkLx0xV68QupJ2MqVY7I6OljoFqr511+tVb6mBGilbV4tNy9aOLZWP2q4Ooa4/QhjtPHUc/p4IS
soChSeYhXA1oVn7rTwooJkI4lSD3RmvtQlR7xoVBWBghxscDhkTfBNpUp4+GZYkXYEuzr3fDLWPW
4i9ZR+Yvnd3VUx08UxV0zXvRIXguFw6xm3mdTGjsfBPVRcoJnQHocrEkR3VIjritzVudEysGWVGj
HZEFlTDhK0vdUdwbH2LJeyhOPwtVDHs/gDEZAyLi5QOMO8QXpT2La7P+La3Op1v1uQvszqLl6QM7
lttzaw39mXBUPVuUqFPn38VBjogUAQXHk99vdBuKTJTm3OlnqXXj//MxdahT8MYSX/inAx9cd6PN
P4skwcu1kxO9vt1FyIR8Ruy0SdLOm4Y8kAMaC3R31qwLCQH8+CIVdm6q08UAZ1JVccNKSVkAr8Df
Nols2oCCKwlx6X5lfq4uHPzqzuRyz0o6l20DNGRlMUrmKbMoYdYka7G4fD4W1Mz0LvvoxolBbrNP
iSeoBg6UHqKOI2yNxQIgwLBFyIjc4Xj0hLi+tImiWB9u5NPWk9IB7tH7d48hGeS9AeNy6yzXA8kd
D7wG/Kt2lgZXv5H86dfeTIM47rJMtPHda7MF+sxVOg4es8WDUC9pB5BU4ASHAoLtlMOvdlNt4qds
lP/VnvLnDjIAbpSNRwN7sYy99DFAZme/M9rkEUTLzDsOb6L0sKR9X5p1xWwwJC0HeD+Zzxt76rPy
SSK3hKwm0at2FU8Mh1RLu1hXANjN3vEcimVerGHlrGwLEIU1tVYRPjzoyvfF3N5qoeuUnWfv3Wg+
YMiXWOswzDgZJATLI5+fB/j2fMUis/FxuGDsTkQmETUp8v3szPxQM6b5ClppNxAq544f9mxZ28ZP
viXw4/0alXv2qkEmP0AgQQyw08903Qmo5wYPj5qlEw9Zly3a7DcOLy4lL0wDJ8IF/+2bWUthjsMU
g1RNQBIhe/hWfQXbTp5DYDHwjj7CBx2DPIg1aDnISsMjaxK7d5FLL5ATUy1nqAHkEGj1urQnfksC
X4mswJFNC4i2ij91gUPKFEdTCSptTAhIYBp++/SXhvO0SVcFpb/hxk79DKr1yUI4J1Y3jeha1DUp
FaPkbO1i9CO3GKcWohKt8EJ5Et0IVaOaBg1PHY/mUAlFH6rTUWURX2kEE/PAaxFyVk57pKc/pcsY
uhj3GTYw90ODlHrlEeRgQWiW6G75zlsniBtLgrurCYlwvWNK8xFZnzziYrtbI+1z8HYCH4b3Q+ew
9w9IT75MNbf5Bfq2YvCFV36NREs/MOC50lf6nCXa6LZTdisXs2wKuleU2PRywhoMr6rYF0NLaqhO
y3sG9N07VMBs8CLErQIVmAqvPmwNBFsoYa6sSMbPVnkDufx/NdO1pJpYzyvwToTeW1kF0cNrSDyX
cWZcrapXnK3IAJSi5E1oKqqVfxb0NEWh8g7utkMlINcNzEeUC5qTjkCK5QaGqVslSDFYd0Qz+35f
uSDFVInrRUSgiGO93rrZWxtDwMLG6QkYgHLjMALa7AgoZ5eRaXEvI7OYExeMDPL6fa3MH9uf0lwe
8C6i6x2u7BPEkX/UGcWZumylXDsgI0aipVPYJlMg9OsEGggiDdj2GSO0QijzLABhfeXoQd4vXoD3
NYviNO9e5+WyGr0REcafjQQiYdMqpk1ckbc6llpjk26XkqNHkWRi2V48bSZ8osOGgCKxNattjBRQ
KKNJ8j5707wE8+UCcq+ClI2/M0L+oP68XwverLCrAcE/infpKc+rNbu2WJX8gt+pcVy3k8KKto/Y
MpQKK1HIQ0imUdt0dM6OBCYL6kTmknVNjlKAlBcMK3DRBH4crVBrs54w4MyGLbR5fgq63IrKO7gN
Y2zloSDAzdUz7yEZXUDmrQeBdN3DZ8VPdrVJUkI7kgkr9DlhAFGWmjU/+IMo/PiX20mPmJqZeKoh
RMa1fM9uqWsH2McOHH753e9d/kMbsuqXoDfHWCSTXsnffNhu8SFyAU8udOazlxBBwP20lnT61sLc
ZYSmhUlQ09BJbv6h7zvj3ap8LiBsE2feOm1bJsH83ip9Qxnmavhq9Ar/UaQRd+41Q0ydO2KAnCeN
whjnn8TAGm/k0X7R1FTKp0PTViwdwWrvqttTGw08DyQnGDnEWSLkT6N0joIt8yr1gY8uysgzVOw7
ig9bOkQyZ0VucYJ64hh6EKMLY/lg0OQOiP06eW9dSH7NHNWNW0ORpYjdiiBrzWJ6DWeCiIgvF+dQ
WobMXqy20X+NRU1/J9Pq60XbK08jwHvk0+V0ef+QoDBlE4+Ub9UXHENOLnYZ4ysyzIzrjlKf3aS/
7vduAq1bbDnH8Ro3YhqpfjZR9dfpbpWGGBhOp+u5goOaG/7LVRXDfFzzNZK2Z5O/Til/leflFg4+
tUrjpXj1M+LmwPQKfsDNsjycrGZsCDmKuPVsDmyYbghbzloeJsgpoNVQbAUnbVKP1ukGw9F6kJHp
+9J8+0LkjQ1Yni0/IZMU4WaS3zGgbhbvthk9Kod7nXK0YCCywV7oEEt/tEsuDRj8fpkgUsMeW40H
a1pNIxbwSiXGatGrDmvcIK87eaoZFRWDgZ9Kl3NpoHfaixMKFqCVVQghg+50VqceSPhcxKozLKz8
2yvxnYYiXMy2RzjJr2hptBXZSKBDae4DwlrNVe3zzBgHNALxvWhZ1EBp6jY/KR+UUVBkRR21tqfp
vYrEJ1mhD2KdlxvaRlpFwWuk6+RF0c1lNoB61Zom4tUBv2xzMt8SECeoFMYaayqHtcnw0ZixzrWT
uCh+tyuN2c/hWyKDatfuhHWAEyEP4Xjq/i3sjI9yHkyJAteDHZQ/PTU6YIWq526kuCMM/p2s9nPs
NlM3YPC/0Uyj1vKWgVv26D12hHcUaFvXdbk3AzzsNS5+ZlPWEpdmWhi5sI7I9m/VG2g1bx9eRTDB
GZCwDgx+wrDsIR5EpEqu1sWa/KX3zqaGFUnG4eAjCOnmG4nnwJFMpWXxS0H+ZaRglWR6DGa89zHw
xFoIvNw2zBj9xIac3WSW80vuakOuZK4Vvdg7AJraTwPG4cjJga13Igos4yCBAKQgeBk13eF1rwu8
EUpjuG7IKCstX4Up+tHIQAgG+ZEXtO91uERdSHPxK6oW3NaG1qgBkF/TnfMWN4FQDDXBGqKeGsDe
nXXbob5P0s+wNy3vuXTsJQZuV6VGBVKGFqk+3KLi5MAGo+kIK7aZWe0yIQVXFJxuhaYbEdPr8NaO
U+GQlNVIYX4iySLL0ParGwd9kzfHZI4+ETFLmZzs6FPi16lrDOtlhoOtsanuxzdEyq+q7Nc4i/5K
h48cqudIc+kM96NV++W7DlMm78UzOGEfHPioH/oMaMCK0ofUIpzctNiQ78FWFramB8sJ+TKTczV3
Nvq3qG6ezeq81JAEwrY2rJmt6UGMPUKau8FtrqsFtljJISmrBAAFk5GafrDmlO2tmx+39kHYY2Ur
HCp0Q7u7tvOjyP/jsZZBG4nPRrWTlOq7Smb11g7kgKpGh7lrNsQ5tGOeaXME+qY+zShILsCeKB0v
lE4nB2I4E0l09EcJVMrUp7z49E8LhjDwXPt5AHO9FEn4rPX1aajJzLmEu+o/qOL4aarDuiHifkUu
3rwIrEHyKth1gr5l3EVjmCKIpLBA3jRCF6zNxNUPNteaR01Dqwthr9If/uBAk358b424wsXdMsOv
czDsgyyQlNLLsEJB7L8HMcTJEbE6FmsxOHlzYwVQsNhF3Cyc2/OHwOPWO29li60xHdg7I1wVpYG7
tL5N0Rez2HcVpDiLmiexuRgv0bdOTEfpr+FVpPYXHYUyi+xl2HhuV0nj0NsX6/XoS/w17+8nT39P
KpOEikYqQzUpmZuRvcOx+rK12QV2p5BEsl6ejwEFuVQZMx+YN2rp7iv1gFPX/UshWO9g4nXeRGIY
9qDHaaJ8otqUZg3J0bVtATt9TtkNJtryBY+QFN7Cl3vOq38AtHdMhLMDABHfOBS8Ut1S87oX+/RW
O7em4OA6ue6kdIEtg859Gj5FCytjTAlCwIWSXfNTdaNkRo9QwOoiUZN1TFHdNCKgeb87jsJ3/7lp
jf0wSl/ZmuSNrv5Zwptc8gOlE6/UM2JMzDVjt06bsbV+mm1hhQ3wnkrMF70Ol/uexOaKdxGZcRJH
j19U4q8rlT7i+aB43VA6TR8ltLowfyV4LQaiFr4t8KRT4WY7dIui6GlrbLhEMLRPt2Vc8nR6AP8D
yX7bCvOlCr15hu/kh+yBAmR1max2dzA88D22SQMTnXOYJR2xYsOOsL6cRn0IEeh2/BNyqxBnOKfz
XRFGjoAiqfiqNroIhoT5xRYPyCipuJLgjAf4CSIeaDETlRpnSEL6gle36PS+wHGjJqVAjXA4E1QZ
w3+GyRymkHTCJSFTw4bbPwISuKbpWYL2Qmo22qxnmFYxnsxmCePozC4BZF584v+3EsX14MHY0/EA
MHEdYlJREhIb/6F17drXyeG8fjvPxqRVMsLo9l8tR6Ib2ijbSsj1dZO5kMopkC1bItMkm+OSeaKO
WvuDP2Pa5GYrOGDdSfDt6TDhCLwYwvurBQQMutc2co6h2rYLNlIdKnZLU2vUjot4Ap7AQAWX4qV6
LF1bUrhJn2QiXVFLQ0oje4LKXJp9h1jj8uEpOUiyWgggvQssPzJZioPsV5Obo4DwuvAEdIie2zqt
i7nq0433/h18UxuwU/4Ba8jRYRQWJLyMy9Kri3af7C3Vaq20zvGZ7k+6kqa0zgJzclDTIsMbMck+
o56U2nLJ6QRN61XS2Etiy9z1eQBEGggeky17N7bUbCV6I1y14+vQ08EaCTSYxxS3KEu/dsnwr76g
aImD9uWUey0Fy0oHx9pSHL/bJk3K0BXy80nla0k/ncQCfxClhyiJ/tzYekD34KVmeHcpiAYyQ2HL
aoQEMQF83N+W/Ul5Wi5FPLVqL+IzzlT84e+2FzDhgI/RYXyzZiiDyonAO8T67KfEIxjuCp8045kv
yof/kCCetVG6px9c2+acONK1V4hWfS++n+Kkq0zq9UcQ4MTzQHuA/wUjt/hP4PgAH/z81i7odm4X
YMRxHDyVYu+Txdz1Wb1o5QYFeSwv4zpHhDJA4ZuVSUCtgRkyyGi+KPTf3REJIk4tUluYhRELUuI0
/8FYk0OZx7UT0Znky6jemMiFsNyxqsCkMWryLruYS/9zSSRHoLZ42FEt3yF+7eUrV6Rxg9PaaH78
hg4ZeGhfjxX+BGgc+hMPXC3tvqb1ms1Yro1TYUaO3RhkkQ01HHXycxuTy6dH7bmGGCvBxglDGkB8
FnilQH1zAiXgpSl1S4XqMXdrmGLLbtyE7m2iyzPYT+Je9/AXq0fISleCGGqJQpXdY8oEglZa+sXm
8W0Pl/VggDZoN/RkaAUERfTKLnNP1kOHrBcLxp3igWYGRALx6TDropzpykA7Xqz7bXmAyuohmKln
UQfnmNRXnwWnx2ck6qE2wXByMnsAS2ObU3+SM7rGLlb0hXAYuw74a9WBV+aiLjfCG9SfEO+Uo/j3
Cr38O55+hwqpM38d+H6kAYWSP6NU41NC55Z6DgJjpgK2j8B0OMP7RyHJAS5UTHw6DYGM59qEe0vT
mqVAWih3cBWXLp97rKQ/XRBgx+zVw2ZQ0d3MvvnjbtYXTqCfchkp5BrvK4qAXP84bchkezWkm7RH
Pi7WKIesKxllAwyMkycUzh86KtGYT8mjveSQXmpJtDoO4I2zvj6NStu75tmx/m4RVXjirGor66+8
4KuyBeYXsTsU35Fe6arxVj+tTMXGxopdihbCq1qUIZdZRqCdZ8dcfunDRMRtXsBA3n2FR6xR/rvA
+0OiYnSzt8ZQmuLjBmS/O8+gnIJg8yFya8ORYYc9hR4Jp8Ggo+VMWObJoY7J4EOjnyIPYDZTR/Cl
iJ3voMikHNqkEV8U7TiCUrk0wOzdCW8gvT163uX8ELMtmnBCU9mSu/Ye7H17wmt+kzfE3cRgDtes
JXwAQDQRt6g+hbBdOzza2pouU8mTYoKkUGWiLpoc7eGvDOdG4PKmYMkzVdXOs1FsMU8pxk85st9q
jlV1o03UUWGs860Io5fvVb8xZR2ee0Q2tHKtQHMvfjrpeh6sRWDjukFC5F25XZCTttrqJAHJMpuA
96jFpff2Zi0el3IP/2Xk1aC/gzst9KFhNNPpA24JxotEygDbGb0zd5uuzjIDFElCSKV7DGq1K0cE
5K6tD+GBWeAm8TgTQ1LpyEHQz1V+H/Pnr4W8+8Iv2oGCFjY/qMfd29p2HqL59QTDUhdESKGzedUH
HCS4G5cSYG4Z0HKuy8A9V5X4086YEWftovw7l0cg3Uf6n8kalXHC/mIW02qFapQFZufas3t7vRW2
UZROiuMSmeYrOG3lTZVE4jkuOHLwdFtqCbtojzcU4BynJbg+XkAW6dqI+0hJWm97j71ALphIvrsj
snGHeUOL75enS3Drqb9YkItcWnhwzGeNJcMvz38OVjmw5+3Vk7D1Y+QY09C6zbUv8wNM//OUckGG
PkPKayX8psfnTPCPzR80Qu7sWepATmKtOEyZpCsvV//+MYwVK/VT9zTQMHrulDUTtIi3BWa+Zlu7
/aN5H7dZO+5uIZV5+0ziabTFmwO1c93SRdPjTqClzpng4ID8UYo45JnmYvvyV8d90cPmFGL+riE6
1XBhvktODplMjCB/+YjygwHCfj2uSi+ibB6hLxhbBOPdCJopsv4SjoAE0BXdLSFYZI1w/ZazLgzR
HlA1ChrktNlEfl+fa7N6YdwKVWWP0+bqry8xqNXTjYHznjN41mlxk2gk/qSUXfH+sEywC6BpvOb8
hgYkchhhzcvGY1Zgch+OyJ8TbfWnKSPCvSPhOMk9Mkk/I0ACGIwVeZlfvEX0FN/23VQOsZMvTj2q
UR7gqKu8D+mFZo9FJKANDEPrNsZRNdRcggyUCVs+0BoP41BSSbNNXk6KktL3dekGyuvoT+xhpPa6
xqUV3P/OJjwSsfCZOY1l6/4xHdgc5V4le8QwdDuxWJePEUvNz8NJV1235zvhQZqOrNbXlegGJcwY
/SX+aFP6hHK39/rQnVT9eAWSsweWw0Nv7I9TcAAdBBWdh4wVibHUJcJOL7UqpSXzkPKkt0raEdGm
FM6P9qqF6JWZ3vBOQ+xaUFyQFQIaiuziz9ASBN0Xhtwc0j6s5gvlLD7LmM6JgCPLW54JLVL/N7uR
N6t4iawhE8/QMqYdTfKNdm+ctWNKuyUNq5n50cq4qcAauPppVDcpzm5uLqMKhg6YQDKOQGBIQdxc
DgzqaZiU1sB9LRYrDe82qgCd75ITxdIGulfl8A2lb+d3mN2AAg3BlgxsudsfGUO4j/G0Prs4ZSzX
r3W7hcOz7WBeXLKQ7OLMwnpWF6Tm/By4gD/+PeCMLMorxWgbhP26y/UEFejYrS6eb9Ns9bxxP9Rw
Q151WyumfPNcWd+dTOplRFiURC8bxUNGMojz7Ma53clAkp3NGQEqPOgFVy6bm1ix8VB42239Pk42
HBuI13+CuLyJC9t2bX3/gqPyP6lM9iOVindGVhuP4N0aPxKJGWMH0BRXGe+WGNE0jqvhtV0I3IEG
3gTvMLyWbr+NR3QG+HlzZ4xkOtLlAZLQYECWeoizvFeP7ZshyPr7CpY5QBgsGdSErMFTLdWcXPqg
6JZBDqF5uIc3HdF06x3fejJnzegnUyCEfIsNCuxUa3qwdWnmbb9XmKxIdhtqVR5y7QlbCOqLjnwn
HIMPTQ1p2MkJ3vTeUDH61T2iZk8z7OeP4tPKwcqdchikaTkSmiEpdLI18JSrKFraBNoj55pZX9d2
9PyUA87MILP5AJlEV4yeVruihWzDepXjI9wepftTdW9vfqMxqSAsU3VSUwXTUR8Ae8OTqpN8E+Ns
wwO7poJAuD3a+myCS6Mww2oX18fZ8LCtFgERGtrdpuVnTEn3Vp2KQOvRVPSMvIsJ4eZBUP6xgPDH
AihKzSL5wADmr9t02og9gbOP1wDgd1dVZ5+i/AyE1HgmlMtiBnr0cZUgcLnqTcqxv0mbk3XKa+1o
C0dgTWVEbFO/ZbxmJNadsXx7jH9xcs8P44wg+I5ST77V5uUvTvvmTicqgZ4hj12ySNIYdTdsj2+9
obJuW3eY6nVIHdkQDdbtxoEVv7Jli2og7/FC07QslnH6eH4Zy6jJCA3wy+OVVsGXSFX6XFrrDnkC
WojLXY8gxdyfweRIedeAtV+hrX8uIbQG/hFR1G5fjI5i4t6ndMkCrXog0dkHPvGCQ2vQ8ZwWgrJ1
KABxXCuUpkOdRWbK5T2ffQQV5KJVkvRoizsWM5OIBPd60nEAeBCLXs1yawntM1xSLv08n0A1fXEk
4AMejJwgu+55dOQjP61bCBOnvTrNXwxNWucBYS9sq3IYuzyxH6vRRstCxTOfWpn7pMkr3v9r/hFl
sMfkACZCpcrn4Lrk91E1jtFSJwe5OhL6ShKHmDexTALzkIrZAXFNxQOWg+/jLjZKBwxAjnAXuIOU
etygYCcWL+wK5CzW/uH7kYXVuPNaVW10tnVg2oAIn0lHTXVaVWUUjQTlAicZEC6PJR9mu2+ca1A7
fsHJBFZO44yS5eJ0w8Ya/Js2l6mVXfpWNEDCGWZNwyKSWZ8b1DXj4iFB3d8bbZQ5RBh7lXcSOxvP
J7I31lVAUVMwVmsgy2k/uzsVOsyhbACkqDl3Yy1X2laAnZfJQ+eXdEmNFLc05egq2cIPx6jdGcJw
rLIyJBFx8lBWjuIdq+YBozzUBLC9Njatow0noHQ/SLYW8oIrmr7cEbhpn0u8jm4qTVSzLUEzdhu3
1CcnWls7ZQRqsIB7e0PRIQEzwl8XVL6C7FTCQa8+Kal6JL9BEeTcxaAZmRwLwULbvyysgKOyL4+n
JhRv5mxpY4vBIEwjUg+2Z/sjrm2aCHU/vFfNZjhthqgCp2/lN/BgLVD+3g58MWz9RcPrGQnH26oB
c9Y1PWV4QQBCVVBHYKiTajxEGZro4deNZHqD6t4rj4uCVDpiRUaEqIOuPjjglhxoXPF3vm5MKitf
lhDuVi1/wwnY0gLe4qiNHFT3JzEaSpDfFB6wJ+8Iil/p8ss+i/O20tOR3QAO0dq2xsMhm/xRY+5R
NKwC9zpERxvBkEoJ8JNXxAd+xUW6l300CGdvcBsWflxeDVbMhKcR0ACOVN6K8jqdFcxgPmY6uAVH
NeLlTQ7R/oHHG+6f0h1mEfVJuSZ1ywET2VpVvZ2aAm/Un7dUI2deI7wRMmu6/O/b8Sc1fpscsnMq
5SKscX750y+LahYE3AAFctkY8Ez+DHkv4Ou4X9KdWI7frQwQkwhh5OSvV/GlPg8XJp+ePy+rVP6N
yxb4xk2/oA7D2bd6FBJvtwaYGvE0eBROYSDecoIzZYV5u8L9+ktkRCO5DuAlelCN4WM8z1C7ka7p
TH04sBx/v2IzVOx0dEF743Jou6xZw0MW7B5zjytU5PT3yz3CwTb+HtSNkVVRszQGncl1xgXfOlgG
TVr4NAKtUWIDikCHGRcQuFUIs9ZkJpsWyVdlBz/y6d5c08C6ZSeAViJ37JGjYtFQ6YJC4dygh5xh
C5X4mPICgAtIsAJQAzpWyYT9XxrRZjJ8Ndkbj5OhCuHLCyOvDTkLx4AGCrGrFTwffJ/p7y1nZr+L
LpkXR9vdQlKPzCwoJOCbUa+jWN5t1jv7+wkKyVHV+qW1YKKXQEnupvSzI7Ft1XKHoYXTyxaVmgn4
GKyP4nC8Lqo7wYWURuY/obaWe7xZQvLIKBrGH69cyCjM2QwEiCIJ/mjkQzQyYqEQeFBv7l0wHKSr
hzaj+SKa6jL/jdJKTypVszbeaenp3HwPpANBMjRKmW2YZhFodGAqgVshue+9/kEWuzFBVh1jzMpe
OQq2s5/9KgbXAo1TMBCsHjUGAbqO7mZoh50Gv8bqLxD8uU54PiThGM7+b11Il2e2ruv8o5TYH/iA
PsjnL73uKTbHxkUO3CnwngYJPa/4Abgn9x25kW11Dwp6p+oDgRkeQeO6gypG0hkndycDhfzJ3+MQ
EiUoqwSj/jz27YyZHZvtTZRP8vUDtxzbwnKD7Pgze+W7rDic6/jYaJgavf+FxQigUtAuVVEO/AIm
090py6fBLSv2a0D/BGHdwuqw4l5x1Q27wMWZ8K1tLAO6Lfg2AojXBHzXhHSVbIPww1uXsLJIgizY
2JwWGasmbxrBKbEQS+zMBAfqCJCnwUTjGGqduap1Ql+RKFrEZABh8KdCJXghZowBegqoW8hjUmBN
jQUoCaTdng3DhF24Wggv90e343HFfDXn3zWNbQr+CFots+mm8TRcs+cSUNaA47g/+J7TUidwiZLf
drblYmYmcS81UnC5R9GP008DPJn7nq6nqHVNoAqhEaQflWWAuE9lY03dOjgSFDuQd22zO0n6A1pd
QLTZVC9C0hAHiNyO6Tei6x0liIWwCxEv2MNQkSxPP45fk7eQNSQyNVbVqpBPFn1eA+7i0NdkoeeZ
BsPRRd3+0T/DygfLpAdSVSLthn7vfUl7dLK6OYZ311D/Kn1e2bPC6DQbvQ80BLxQQlkCySzNXfV3
Y0MRqfd3EgA2GterwxNbbtiIH2RUVUBqy6Tkxr+xpVImWAwFUke1H9eEUeZdCwZrr9GTicQmRU1b
0xq3Z0vynbvwHk6bDnuu4iD6yvW8lWJfOlNTnH6s/MwFt8yIoGNQiZ8nrWWJmeXmtzo0ftPhVJPM
dwFQKETL7Zf4LKCTKigC4KucFsCiBvDvXKl5l+QqIh42Dlfm0CF2dn1ppoDmVsuIAStMD71mYc0O
oXrZU/1S37FtTppJXJhxorOCNdRhuPwBAG3byhCZIX4K5iZqsWIahk/kIR5o3/gBIYEHofWxo+03
lYLtWpljvDLqy+4GLMjq0GO6MRFesx5uqlAkYRylhimFTQwJhI8dn78EO3r4hZSh2y+UzU3AiNuf
Ly7qDvz1q98cTFG7jx0NEozHhCOVauFLE60OpOx/kUOsBc7ErC1J0P1BZrLn+Un18o6Ma69VeG9D
+zVaqtUmQI4LwfgbHVWVJjW6+XTzlghaG+j/UxDfkGKK3HHns+bsSISOKwemuzM1hj5F15+X+MDY
zisSEsV9CRrsZ1WhqcyIRKEGl+FGf1TWVOzru3bBNiWC9l4WuoVb2oTDda3FtWx7oo5jU4HYH+jv
F7BSqhLR/CBCDU1c7m2rq5SD6fJKIMIT/og4hMpOoU9C/AO2rqfJ06kFMv0dzuxqTu0dAqCwvN4k
P6SamCBSD8ctUXROGoUAete7dGNOnTY6VBOJoyUabxxOadelyRzF6LKBENCSD6HAGS/HLzZXs5Lo
WErP0Fr4iqhMo59SETPPH+lWG/iBalFDKhmATUmM2ZGz5A3jzBNawM6hZXKO9W7YXSoI522iKQZd
Y6BACbaAFdlp7QmvVM71PKf5NsmHM4DieQYD7/a15LryjHbKtSKguvrojXJuS9IpD+kduciiIH5M
eqsex5jt/k6C0uRVEPXMLrTBTOD7jeSOU0ReCA1qTjaRMZJCn/Qo3QodKG6uaGqDJa+aWP8cGzVs
RzbTR6XZ8rnuG0Wg1cV9bODekz6yWD3zFxsAvg0cKvtOCk4cEJ0+LXj5Obad+0dTPuyf0tTZKXuD
KjRxIL+8gPgMg8Tllz2txBUs2hFL4wgqhDvNrFVrWj7bkt0peTKNUmpEOf+2fwiNgros2isdCeYm
PevnfgIDWq4hKjd+icjlhKnva0S8mTBF3iiPIjeW+/5KmHGkRahwACT82WyYfRq1K9unDXKx0Ts8
4aMENVF9wyUjH/W2liOklzg5HCgWxaCu7gH4fk+7e7gJwdhCY70GbxbXrB4Bfu0P3TGwjxzvSXwj
/G/mewojRVPc89OESs7vsSoSxSTSZZHZiRwzWYy59ZUodFTCYlI89jOyGbSQHwNMTgZHtT5VxnDg
GX1smNfgqwiUHd3lCYtubJA4ks5DPTEnnvvpH5pc4cLJtxJ+mP9sIo8e98KLkXoosmqmqhsL8EY/
0W2pbXlpJOcXKZHq2Q8tdg0Yin+Qbdd2h5zBgPudU2Omevugp+LbVw1OtsG3Z3A03KXMop+PJ3kl
iR9UeYAyvnj0s3iS9D/rCNbtrb9Qb2+YJEh0vZpKnz+eOhWqbPPRproGvFdtkM2ldZMOm3T/s0d1
M3cMGs37Q56sCEqMVW9/sZjnrwiawXnK8pyZLtQ87Gbd1q0cRyuQceepuYcAGsowU8tGTWLeL7x6
t9DD3R3xMzKppMx4nWtOM3ts9ppqgd1UVTPLVIOlHyOR4NUxqXbhcAH7i2tvYs++yYo2V9Pc4+3t
JGtnVdQHuc/IllK/Zf+nlTkBOi1dsh8CVewwT1etgRdRtvTILTiE8ZW1mhjQO9mHa1S95rbTakTd
kNNmnoQFsE+PdAri6YU0aWCy6A+7hy1k/gw0IkPfDM3kDzQp7PQDsWXS7VghPSD8NwiSTH93bIFh
KTcC2a2Qmh0sos9Pa/6V8UTsSniNTOvmIlWSNxA3XCgShqkkJy+pKRSXCIbUwarsSPM+7dX6c2As
QHoSjWCDJno9ADgbyawfJRQ7wTduIAhhU1cn1+EKWORMG6kWJewIScLFI0lrsVbtRJNXNfrh0+Fg
xmWR+m3WxRJKiWlAiDbLHKKzisfUcDR855tgxfErYR5dmEK6AYUmIi3qBupw998jFxnC+ua6aXKV
AM8Jf9irZ9mdFCkviuYWwSS3dfF5erdwBUttvhfmlpnEdrjDldhcvy5EeutjFmXXx0VGBBRJe7Gy
+nuNLkMV3z9YH4pX3y1hDMdt4k1pAPu+rKnC5a40+9HHtNq4xXptfuZlLqIy+IjS0ZmAvjzquM2Y
cklBJ9E8l0EvEt5iipRr6wvG1Hw/HhOlqG9umNqTdY0TEAKQH+pnfgOtEQTQTrEW2yOQ07n10U6C
kP6FUhsI05FjNjO6uPXj5YwG2ONy1TynrbPpBKlFbg/Ra+DWerAVcdWFt/eWF81j4+bh6kVDTJ0f
i5jASMEywG38z2IjbHegg3l+atuJ8+AzAhEe9ygj3Dw+sGdJ5WIWb9udXFkSJ6DvHAS2eDhRv6/b
eeK6tsq9B3E/H5/EWbgojQ1cxEyVTHyBNeah+YsfWyN1+vQjX+E/GdqK5FVzsDR9xL+YbqAO+rhi
eDiT17JOmvRp4Q08vr1v+Mp0PnfI5deFhtghIF6c7BPDWPGN2rctq26scpWBZ5uU+6pnckBpg+NV
pEb+gXhuE/By4CyB/va+N/7IHhjIfuO9UyGTjuEPzkbcIRjot7JZ8Fd2t0jpBqKBlXVCvUWKlT5C
pWyRIGUTK29ytUccqdSfExQ1VxtapBZAeTVmeX5U4jSgbgbjvlr9gWp1+TXHf/dEIYKeUgV8d3aQ
ZcpdDOPgM+SpdreILl2CruMBw7NdkM3n5E5SA04YcwiRN08tMhV4fXCitTbGa+nxIUPn1Ef27tkt
jWM2U3vlClFm8R7cuD5NM/PhaIAjk15cE5eRBA46hav0zO3SDrF+7lVFqD8MXT+36WV9X7z3rpgJ
JhxUN+HjGvvYOx0E5bmZqc4OWu5jPkjUShAhj4uLMWtPZZD1Za8NCP5m7dYpOC8Q6fPxBVU9zo57
x1amRRT0mEUPO/Tle8UX+P8JkyNvV07ysApiV3s61qNGVU/BM3Oq69sMWqqDOC7Ku0pGaOFrxrDX
cLTV18D7US6SYujY8IwTMX9nVxTsgS2mb9u0jHxN9lqSnS62mjNVGtA1PqMQx9pG5wfwxU8UTSjb
BdTHz2dqz7+jl3f565hRvyGgE/ijpkZkqF30hLshJ3e64g5gwobTAykxgMhfpnJQCMG4rq3BYM6k
jiF0YAyIKpgCnHa9vXhoUCrx0RrKknNqBz8Q6W85j71nhojt2RYOMbGjQnDqbsIT91mDTBv1rj+9
ePl2fo3mbTcePqQ8Z8u+qfWZV8xlS/KnOW8NA4LhTPm2fIHzr63MXrGkcfWgmp067j4f6hZZoaRP
lnT7U+EVs3NlM2lJfHMzPYR0JKXnN1ilbTHbw6yFsclTEgDaxmt6YJtIXNxRuvrm8Rx95kGjAXyg
WnV5aksmcMdhXKyESZMwp+XVPKKlcSu6gdhdMDYX+Q61cxsQbdzBfhpzVxFLqFly4jIpXnkT0NMa
s79JYOqXaCyUZwgFuAlyiyHN9Lt7cLrQfhLs+pwo4IqHsnpVvfXv9W6drPgZF2MDWm7ofQ4Be/Ta
0eUnJ1EOHqq/1OW6jdR7s5aW1GgQRQJ8rsCMf3pwx1pnF7kNsM5lp4qzCNTNWc0wotGQNN2ymfZC
0W27WEzxaKRHX7tPmAUG5CkboZbR99mLeUdstkkD5Oy1r0+PuatJhBW5Gwg9A4DO+rjtc0p5VxOT
EF6rH3szb6FFewqeZIZImwxkPuKIwDbpESqRilQH47Oh2yiHX1jJWBIfeOqB2CCZEdS9jQQ76d+D
rK+wm3OYAQjbSPA+gUoiMay+1W1EXHw/4zS+H3IuGHb7mJx/5DftHrkDhr8I8PD/V5AhkoGeMuu1
c8mLJwQPWzkH7z1gvSdxFOy1e5CAqhQNfsvcgm7TKQguJ8X3SwRIn3SRCBOD6dBQkRRJ3B2XFMNE
ZexKRHiJwfur9o6tnvLhxGNiiXYhdxvNj9IqQWD/z4R101G0nUgosM5DZDK/rqu3xVOjvsWoqviE
s6kL/uIDIM5bmYkdbYINqjPRWTOKLCSoM7huHrBeQ0AJHMLmkzWxlXgRv28x6KR5Bc7J44UES05w
kcswiD5O54lK5DVrbcLsgRnKxTFgqafYPXYlOlAJ7osUaGW3e56Y/eajKPb+AUYAPRfwa2wjj9X9
7b9ArSAq/HAodFKyrB/kTdlC/UIvSKLQ8qz5IlAX87JP++DthkwTeN3Iv8pMc+Bfex/4iK+Ca75N
Z/IQszL9b9W/YdSgZwsLpWO9sSL5qg5Nq5DPpl0oVq4RP2IgWoaWCrYWsMkEZqwtYTKfYGjsklDQ
g0di0Q6o+IE2h1OfRnSuocNq+GSvxJpTGIo7b+9IdPMkgBSKCmGFY+3n3DaHhx1agRfPQEXKwiLj
1dVckWX9mAb1l9eO5NDc8tJ905QyF/qdV0326Npg9xjyKY3p/vtqvdC8Ks22dGLywHnWj7O649CP
sIyvDOwAygpST/Te0pUQ/SKtRh+bDg6TODUf/vJ+3wO0YRmKIkzf5XFQGCQOSgGVcKETJh7zxoOf
8XDhXLcdEiJo7PW8Ij2CvaMVCS8SI9tgSRRbFn/t6wBBAEHoRzum2UlqeT7N/scXx6ogg8T47Ula
W8/LEnkEWSnNT8+Q9Pzm+0WcJ6M5LmxEy+zQu6orvQDnL+p/f6IPXJokck3EOevBwfznu72zdYFH
LGOX0pldfsNT92uvtI8g0vOc1rxO4gvVNbAZS4xy952tQYZ83kIXVMvHU19bqocF3bjf2ux6A13J
M0KgRitsPxwBs9x6KGS+XNlRu5IomKp8EIlZ2AM5X/b9oFf7Dkg7cIxOvRcUazCkTSjlxrmj1hh2
pBOT571yZ9rCO+LF7HpgbADfseq7mvyRXQGcX9vt+UJD0SggAaRrMH1E2yI3jJtV+iCh+9hXdXyT
KkFf600jz8ijhzHm+AJz5vaa89lbgQxp1r3NfTuGBjGVLZQpSdl3XvgTO+0z0GM54IjqU5Imdlnb
Z8EfNkkWvIHhWjRWfh8Sm8Lt3FHA1gZUaMMFHaYzzfEVzjFOnz5eNUvXZnT0SGppOc1yAEljkhDX
MR+lQww5jjI+3HOTIds7UqRM0vvfOxpJHzSM1gTF37UghE4QeRg3hzFRHfoqtE5LxFqWjKOhe1fo
b4PFfidN7MHy/H742SLxjrshlENZ0QwGaMkJn5gZVko7oLrDgPhQUwRWJZeL3wnpmem2cOwq013H
vcZJOEfhtDA5bKmUWjOdNc1kqFKablYlYPqKlztU7Ck6hA2AgCJz2pyVHuzHzRvUy0Y9L0K90FX0
uvjQh9dEcPTycyhEOIZHuv2TRQVAk3HomdaP2Z5eCbAAMouPreQaIwBPDczBYKShSy+o3YcK+4+n
3uz1uC8Qkm7sa2ZqB/xJL7KKSshIG2AGEh/lYK+Jk4/Lek+FCp+lsVhvJU/1YBSVWxHEJNgypIaU
01DclZGZ7AaBlE/NiBoFAznZcHp9Qns8kk9GK84PYnLjKmAclBsCNhGUe3E3RGXSpzydr59mqAZq
AGCCqRU58hBOjWtFeYNk6GYgyyExudPScMcZL6rohfjzQxwqWGTWLQe7hurouqzP2gfp6xnT9ImL
ZnTmAUXoVfIi0Qh9eKyeKPqYy8bzy585DMfKEW7QJoWjyQclPX+6pZakvUJt9TP0SH5Jhd+PTw4D
JAHRb3LkC5RQouNSrbYOOsB1GDBBY6GS6wl6CILbd0+BvXLzS7HuvoIftIR59EpgE7PEK/EBkgj9
uDUqwqAXisF8L+/pCNPTk7/8mm1rXjowRVOJxa9T46qPrvCOfYzBEkBkSOGneXzh45oBwPY2x4Pv
JspYtWvUK0z37V0UAUfCElDeWsixRgWdQUg+BbgPrkuFwcDK9AyWYlf2e0nnEiSUAfbFCYK4hxSY
TS00eqjgrAlLLZNGWbgt9FoVLTP/3dXN7I2tCZKldgwh6f3GLoDyLs7+lQpGXlErwBb87PFHGT1D
krkPUpEogakI4Lry909+7in6UurL5yhxfLa77P8pw0qwqqyF6Hb1/IX6x+TMtTqUhIbdCQQOmPO0
TcLc/vZUHSclbvgXVuonUSZFUu3VcCFzqK6If3zi8TSzmNZyoQnGxkqmXpkTYtBqmfHhcEc8amio
VZGMQZeMq6dW7D+4bHmOStfITcLk23AflZw5sbVCWj2ww9Ac7Pxk+vGXmaWgaPR3XYDMOQ0p4VWS
oEAGAfk10aClWu5J1GOSHjyai9xhGz1AcevwjpVoemOE97jLXu//Wh/WNrOrnpSx/JplXsZROACF
doN31nScQNcqWVOcY+R+aR9g3nr2RUXXTRdq3axqscLw/r06rRm2o53fGkaOwm1r1Ll6NoIjVlTd
KrT/SpHDZNSWzKI8YYgPFMRZKFIOSpcpLn9GZUdGdW8FA/gGMQZ9HLnxl2o9Kz8DLRCojej4LyxB
tWrr29KkhCUZpsg/BiNZbOCQlilFvFWVZSPxllwsuJITuh6x4XRsXo2ysT6kpqqBEO/uejdY+0Xm
Q1lFDSoOOI32fEg1sufndDRMg8BC0QjIgaW9REu9H7POcVO5OXCMIKmppy9Yj8oyIPfVAWqr2kWS
BECWv0hjx093PsIcIBKSxJSvlhlCHPzlRopndff6higf3UtiibBQKzsVW1vg7k4ZUJez1KFRl2Gn
a88n7nOU13w5j65tvQ9gbqaleK5+1jJ83r2XOV420AXwBWcKyQXonW+D2a3FpLO5brBgVpBaQhv0
sFI5HHf/phMWZbTb7XRcpDPtxB1LXJcb5XD9MgojIIo/5oLSOvwQ/K8KHzXYYWa5f1met2Xx85sb
XCEvldHvbl6k6+5MwCMDlENwi18I43edqoIox7DGMrTSuxqt5rsq50pDTuywbX00Pyn53PUvV43o
LXyaI+/XhMktyCkf8EHK+nAgbXx+ztefLmrzE1eGoDydSsqKraKwg39XNP/MfoXkE9NAijFb9hu1
vj7yKjyukKA310Zo12StVihBven1TmQ6CNRavwaKhumEzyhVhLY7Ho+szsHoq3Ou9mI0cPf6qyV/
j+csyeY/JsPekWolWPV1eIPgB+dTr62cNuSTiZx4IQzYgIArmv53bB/xVdtbVKHpMCO4/b8Pmp19
8YmX+CWUFg14p5krpLjQApTTDY7rjPJg0vhcZR9Yogk53Mi2YxDIc6imwhkefttGBOcu1kbJE56D
MDY8Vs5fgIaeE6DJBH33zF0wTyI79f1YYlWnVnJKY5hImYYao1nKkoHBY6qxYa1fGCLs4DJSMiVT
Ilh9OZNT7QUen3c6dLVfE7RHAp5wKau10vXSUU7HeAb0PRYHCRV1fvVuGdvk1s+hBbsX9/ZD5LUH
Wb6z01sOAH9lTskAbcbuosyYhElq/eF1TRLN2kf8VoMFvkTcb1wE+32hH1cEDIV1/i6kX6GOYFIB
4kChpqOdU7AybeFnrbFGKEykZbk4PPegRUN9vdTFgovm8qIMwAXM6nEIJNBNC9t/r+MDfTwDMpS6
mOc5vXzVwLC8nDuajo9XISasaLvIPn0rIDrIsblRLw9gjmZ4tu+/qMCo3VwAOXBVx/Dsr0skq1+T
YGCtCE17BArvF2jd382PTPNFjqDmXG95kYTsdio1IRpmSQQUZ/HFS+qQUYTNha9z2y6Or4RMHjv8
S9uxOScOhTgaW+hn07NX8Mrgs8O5AJCLiQZrvofyNZCQrqEbILv/Ej1/iTjqYq160sfggiB8roEA
6UpGsvW/yHtH9JQ8iE1Lei9pc7oo5e1x66k7Zv4SEYkcI3jcf9FFIM/MgFHilKk6HLfihNtMu6OX
2UcrFE80C100GJF07zx9zXlrJa9i6lf6+5PbBDr6GxPpRf634gfcfd1KQWgadYtO04SsomAbAUhq
vy8fkMjpgFuGX7hK0M26wDicDCtNfUafErHsIXpnqaSPWtkNVvnrVkMFPhyABjk9EPD13/ClEpDj
sXZp/c+IRCjI6ypMUhgU+jyX6cyqcCesyswTdutQXHwcplpK9XqWaWwzkhD4tweYlUMJwe6qtTns
I/Lp1lwRDTRSG9QafIDoxQak/I8RwdISFTIjcnr5VqiQ0b7243VhuD1Y5QST31W6RmoSjg1sR6II
cabrEphkFctm0kw5ADwp7aQB1FYh19TBmB9p1EbvpSRBJvHG3oWDY/4mEmUTvmsVPCypY3q/tRRS
BXdtU2bDSFu09P1RhlTa2eW4qIqJu8zOfgKZu9+Se7HET6BHU4p4USZi6lAUAmqj4KKcR6gOgp2p
lP9oTcH4qhL3wWH6lQPUa1UGv0nKM8rZ/uCo7zzLxHLdxYIjTaENit9kTmggvJRG78h5aEqv8qdc
SiWm1D/eSYmY4WrTguzyxtj6Figah8utHTIjeCXOwn1GOqVfxKbrq8PCHSfxAQpw+1EFjxw7fLKM
iq6alqQ8UtGwrCRh4Fo0Yu3GfAKMzpgPfZDDUhLZXSmnnJhRuGP+RgAdbJBVYX8YiTRydb42z+YU
dokbMrh0WA0P0sghSplSFKTVYYNiGxvbvuzV6GnoXzOpVW3KYzkK9CDemt3retKS1sNQ6FuTfxy8
mGMFqLttEBaXu2vhewos8rm0WH2ZWDcK7Nn0WmdWayvcr47kZaUlR8UmrUzOdMuDl/ymXpt0BbE4
/gUMXraIfxixLWzciK9v8NoS716cCaHaY34JdJVHl/EsdmaUDSpRBr6HW46eNYfWRo7VGOhbwzPP
SFXHfbGsy+eLIN0d5e2trBBd/ZnJZ/ttkEzoa9tUBLLQ4jDMAzE++ljFBjBEjMXl03jm/9VdfFm0
t3GkR6g3dN3Ci0z7sByDFT4QWqjW6Q+KQXEkVTecYOmE32GDxCWCzoDFcPq/oAeC0FF6b0iNcZsa
8E7ZZZUHWi5IajJ+s0Ztd7w5z2nzSxi9GHoLqH8RMJlw0D9HalEIJ7FSpawxNHmr0uhJ9eUTKJas
jD2/KOYtLyzsQElbWF8danBfWzT06rWy3ywWK8i6mxOcdwFCsTkpyO0hRvyKiKVR/t8SDPabJeWy
2TpC+5cYatiIhUCuUS8JT+Ct9yopqWC3ZDR5F2VIjMkZWDRq9wg8Ig1ErjyuWgTl2l1C7O86qxE9
lbDG1qvB/1/FoFk8xkvCjvz3FGp0h77CbzQAhzIB/BYPJ04dSflusQXEUPSOF/rsDDYVNoz6qTPP
ZuBlrtxPwzFTKWnHnAU1NDcqfo6+8VrvWAwAHEVO5OUkgYagfbSgQhuw0s0Ue3RkweQsHqzMEiGD
EMqSHukQ4rGMqvBD9SPlWfDIb2Xb/3qajoXL8vKnu6zTTtu9H8bj4E3P+NKXKpvN8OekENaIm+4F
h/tFpNQ6iKCy9kva12H4y0vS12Mu81ZkUMm6chRcItkmpIpTzlz44YSuH4qdG7xbr0fhX99n9Z/s
mVp1VNVaHGzEDH13mfwi+Wz6sMUnQYHpdUqA2XEpNF2OS26s+y6p1US8tx7nST99aOH0zb3GUYEw
3W1oq4ekWChs4nRtDzdMlp5e6Lj5cEzvX3CsC24kmBV4LRY8NSW6lIN4YSsXycYnMskCfuGIf7+s
UOt4PqCgrSXEdC4KTmtsYYXCPwOJxBedO2D+uf2D5LXvzwD2Wk7DfnuzoMJZXGHLA6x23S5jMoGm
E+4xjw8FEZ5EjgdfsvPcWYdBRejOru0dKb+ODtpRP49NvqoH5UC+QVnc5Yicceu8EiEXthBh/eP/
AuBCsnja50WW7TJskLYIZkP4ULNCQD2jzE4hoAABsCPsemGAmgqNgr/Np172iH53PnPc1MhZmezb
xV2tq34hDa+9tH4vmLW1MWD8IDAJGk3sAC3gJ7mYJvhNtQAPLoOM6+kRjIzEC+WHA2WK56IRe3qO
aP4OE84NetdJIuHJzG369EEOCI+r74S7HH15cG1bdtJtCnet0OWkctPwF8U/LHUVhAY59x7a35KE
HsJmpk51IDR3G9fG2UqLKyE/ac63cVYBi+34Yf0zYm1/rBPu8RJm1XMuF7MuVRDqNhTK2xt/n065
gfq75Lc7tbo571kYxTGiOee+FKmntMK5caT+kLagPwzeAAWJlDYyyIU70RruIyppFzNB2CKa0owX
jc7evVrxcDIy1f1lalE1RDTGe+VfpaueylRT/kO5Kgh3CLd51x1VyUJ56/NIoACgGulAriMwh5G5
r/mrDNm7WQ0d6liVZnZqQhIazRHbLGGb7B55V4LKQ8S9RZabfN/z4AVqZJMO8Jg3GXDeGIGkEdNi
r4b6U6OSaVvc6+EV4wYukjUIClhLF9+7Cm7WsZO5Q1gvpl217rb1bTOjenc2anEvIW4aeb5WBEXG
izdhWne5lG90nMNFXbXZCIVjfAhVjXMl5PKVlL411/K4fa0sj2MvE1z35x+tqs6P1oH4f7b169m5
7BIYNZvEUgrRGCASRJUllT0CTlZwKQcPcSAxn+I1/59LIGgLRbo3YlAkl9O3HzTed+Z6aGM7bNll
dRevbIf9FSJMHwJRCrmbB3KkpAodFJrB5Tk1MvFht2QyTNnZIKDN2NXTMIrTFCpFbpQHQHXYiiBR
QEu6wXZ9R2r5kc8iRlIxKxcGfUo3zDct1QKigChk+xViHKPyeDTIUZGw8XVxTEU+6MJ/BUQlpuNW
G57tgZchgQ5g3TwkbwUGhZ0tAJVHw0F7Bhb2oa3qEhzphSpPlPGlgW2bUqWzYrnNPIMsFSsWepsT
Tr8zLaqfQ0inNe8b3Z0wQh7I3Osis0GNNxQ3G5+fcjFgLaUlnMbzvZpnXqPJHwnAi5GA/NuPpDrE
JO92vhjAkIw8y3i9stpluAxCKDDjtpK1SUZ0DogrE7SQIuSZU2sL7UmWtw6D5B7DQRKzO4tLfC8l
TaK7YnN8Quh4DM24SpNzjGrlNwwl0cEv6JVAshRE1lNX0ZTJzDDRmkiGuYRytd49xJbDk+kJ/kpf
yFv58g8yxBC1nXWn78bWM6NWPeg4/J2eUAzEy1SVBqB3Nj57HvCzyvjgSLLh81/RmT+VjHrtorTc
aNhDLZCBvYM7Z7jzbWUwdni21QhgPXEa9EYMc09zVrSRyLsnZYlh/ozPdr6AObcubdtCsZ/xgSUx
6gLA1MF74tBfgugnY9pNjQse8jZaMl46Oplzvsktj2RlnU/5msokTmzcdUe+7hU7udR/2uU+5i4B
NeFFzaGATOc1Nc4LQw75qlLqLAWTVmcb/SIKo8VjdmK6Ld9QcKFuwP9h4+Z2nkyeKh2ptDjKXtSd
ewcPglSEJBOQkAsW4EPrN+xqV691DAhcJrv530qyxcK3VimcVdSvmIGnMMdSwuVzC9pGCEiyMgfY
6+LLOxmIx0n3ICwfzePWRmkDnZp2Y2uBxjERYQc5xQsfHOby/M3jxZKJU8T+L6qRsSIHj9fwl0xr
58y7Xby9v+o+yavrcDzNxFizCTafqvsdQ4GEgiEznnOL1aI5YUG9LWZrOjq2EZNGpVv5hnKahaTi
blYtqM5crGq8H+0/Pb9q7B0HlOLb8MPwsR1FoinMWY5wrQ88WpX17nItn7X4XaGMfAdnw95ejVoC
1ojuXMlYmxz1p5uvwFCMa13cui4IRilcqgPQjsi9/tppBIhbIg1cbJZrKApQtILMd9UxhdTDtrTJ
chbXT4sBQ6nqXCeaQlUbLh+HUoEjaJvinc12J9SQsh+v0kTsK54ZChE41O+bpTEDQK16MvQG6tH+
ooqjN4gbsNGmBNQU7uG4PJqgHcd7dmXAZTKWxvo2Z76kLTeHQtnwwdPRpkdllO8Nten2xqf+f50g
OpQh/kpK9Axsc3ETOeFt47QeF2sq5UsOp2ocvcLHFQ0PK+CDs7RSg7n2KtGHe8nm+N/DoCTsYvJi
xlfV1Hf9Z6yFaW+3gn5AY+nnLYGKYZ7uZjAG8U3EdQ8ESTTYEkoezJmx/piW0sqBs9RU4PJ/jJLT
k7nZvN7b6bJF83afxp+T5GNUuwav+fSXG5Bp5/YJz4u3fCiPCDxaFw8K3ln74utsJfPhmmAxuGFE
ApwazpyTJVSOgHmhcILvht9IZL4ZjwmOo9G/eW0BDpb1ZBHavoUbWLeBi1ht1vPkS9xkV/S8gA8c
oD460I9MnVD9rdIdUfhMON14vthBdQu2ZVJIaPf6BXqZqs3Bl33HR046w6ir/E8hkAdgtjf6X8UZ
lGUK+VVqVs/oGIzVCXNlPRPt5Q//y/IQEYRLkpgToUdE4Vtc2TXJboj9tOtstZdWzJT5SON6qIqv
gF/cp/pYLqXC12M4UtEWMpgQE5rcVkiIwEe4t8Bj9t6DQ10ZAamk8mAFbryYAQ7d35RDq30EYTEM
vGX/SsQ7waIOSKPSzdVYQw8oEwTBRDNR5b97j7a8V+cj2OPDdbIHYefAwLYzakjrRKoB0Srm7TD+
6P8I+YxIt1EQvpneq6AtlIkTOpuAzndJap4RI4iyYaQcpH+PHntb36AxtXLiwWabUXg/nuVU6jpf
o2MO+JpgFpsB+326SR6TfVnzELXPGzSu+D3yottRLi6Wu6jnQXrC0noEh71D4lO6vBS5cX4P5pOg
eh5Qs7x4VuPk5Invixm8N+1WF3TrNkZYa1K3QJ7VlIxNHuKn794hJmrgaRCINf7O+DCMlpX/eMlh
8Lcs6RbKsYo2ayCb4tWGcFjD/z2CrWgXnsJatiB/YCoUrtVymPZs3qVr7bwoutJ+aHyJZh2OFtbc
wub8cQyGkrfbZFBZ8v2+x2WNWg6a3dEyoQPP/rZZhbSgtHlGkLeA1RxBn3dxEkvqH4mblKoNiPU0
CnzVwJbgDDAqe6q4HNooV3RzmobJJ32JVrpeqTg5Ct12llXFYkKuBNQEWhP7Tsy/jtLKkJCXjhax
klRK7C9bOiGvk9h3AiTd+CzFQHiA6DSCtzZtyDhXAmYqoOsTHw9MzAWTSVCj5k8OnHEgi1UpKsfD
v/Z9sYLXdADwakfmTEyU+HV2KZ4tR1QUzIoooNjYk5IpPB/Qwocxj4+ne0DfXkakbjtC8sG8f5ly
/crp0lvl+TuXm6IhNupSPPlRNB50rbAUjOPEG+XaD1Af2tJuz7Nzvu+tmFSr3os9u90oVsOOUdDv
kU+nDcIE07UbO8ii4Zl1lReYPQVUsCMeezvDZQv5tXsH+QuTxqt9skKH16GH9qmtk7QeK7GvQ5mA
siiX9SOAhJRyTsTplqWmQnT6bgDBManEtLUN3k4uFwfJb6JF1aHP2K35R+agMiA9na2KLx1ZkMBr
PJ/tasSkR7FrRfOa9xdfKnmEIvlzNPZwKykFa+OBKM+Gv3NTXM9FdOIFW4hfQQfljmuErcMi301H
lkZiJU+higsJVfjJHmpS19hCsaoR6n7PtasCL/ioj/sGyUiZ5Y0MmyxTT8Emu1QfDuMAH2g/xWIf
qNg7TdQqPIRAgivsCv58taO1qR+xsRBgpOTYa4nAUAgpWmNCYJy3lXpttt3SapaxBJDaHiBcZ6vr
eKOj9sYB9ogVSuT65gnhbHEUQCW2a9NiGOXffD0EXmG7N0QkB7vgvIp/i36R82YwD8eS66YHUUOj
YiLZP5HzT2VDMJKG8dUsTrkjrIKjxiqI5XMoG/8QDBsWTTJut93jw+tzUbs7pRoJFRD5yGgLYq3b
OZFzLod0b6Cy1akDy3vKTADX1bqVESdM3PMZ0o614KJBrGiDLDVDn4fjPt2fsvvRBcAthl4n8Cue
7vDqk5M3H/DQKzJB+EdZUbUn2BPdsOOCgy65CQIXsC4uzH+LRuX+pft73rOM7tq6PlMYKM8p7qG6
sQuipPZkmEvZaqJFInbPDUF4KIWiE2uiTbpFGAAYAtW3kv44MqM7a639BJXkOW/T+ZplhBmqZQqH
MYCLEHzgkenKzVW10gEcG0B5e62XxhSn87meEZJBzEwSNTRBjcDrLSQrA+bFzRdRH9yzGdXpbAJp
UpE30+kqhAlHAVgg2u+eKCtwFE5Hx1JEoJRcSHonwSrbz6TfYgxrR2AetzCivsyf922wGqwuZDN9
RfsLjhQir7z/ETZdg+/zdzI4MQSHcYOqftrZNBp2sfwqloxErH0Pv5R/ARbCoYWzQrSZZXUYKDO1
D/Fqwbq7MrymdBqccsmZN6yGcOa9RGVQun03ThneA2201Lp4OEDlXbm7uHOvkUWYYAIOUP+y+X20
NAt43jE2GsRGvlE5hDwkq3pijA3DPPndU+EuUSgPmFTbRrlIUnq5cDGmIMLI4oZDdehzVbnjNmhS
rb1hKYfJg5vWJwSwgPx01evaxU7xRknCj5mtaqaKCgMoXpoNLQ3j7TY+AAYcJJe2FEa61qEPW27t
R5VOaFgkLFppYh2PlUJJfOU+GddBxv0KIVPpCVo5Up8ecpdX2mG3ZomDitv912e30NaDE94xT2Ig
5DzVMT7i398kb1Cn7VHUaixEGWSLpIPEvGVVukligUaSGx08P/zyU8gX9XwiJ55Yhh8wxD3KoXOe
Sr6Bz1G3+FAzrUcIcina4BbrDpPAJC+QvdGVZPelleG68XGCNLsRi/ivBioUfpkmIem4bgQq31ST
WLiQw8ck6me/b5RHEmIihBEGQPANIGYc7d9J0tVPk7jyhje73prEbA1yhEWga5f7YMy9VUaBmLrx
NKfJfi6BRx0ffz7d7KXuOoKDeQNn1Z3giS90hKvvJ0gToCTDTXJ+FSq685WPFrmhBQ+475IdfbyE
gaWQLNJKwdmvrNP1ILSP2qKxFxCTMOM+ot8txU3/S2ozOs9kzQ+tWq+nzyf1DLuJm4XNq8dFsu8c
paaVK+NMisZo8MpO+F5p42PpCwi4FkeKQTEoNJ8e+ip5FnjcvFn37bMeP0MGU1sC8H7wQY3BLpHx
yCpm7tQ2Zk8Ji1It1qGKnZ0fx8AN1O5T8f+nMof3R9mTVPBxZkmhpQLPUNQIEy9zAeUPqnxerORf
JvfEVlDDI2GisBRN8FqixB0XBIaNkTKDSPAUpxx4NuAHDdPR/q/bZYRFBAC/wUCkPQtSeOc9ZyHz
W4koY6kMCcYs5hvK5QBeuLQEY/KSgzMgFPbrZAoloSawKMaayZ+e2Jv6gOcqWqSAkWQnsPLpq5FI
DG3235YB1OoRP5quLfSOG3yIDGx27hSne9R/4gfuH9a1nhfR4W+8FutguNccchMIvVHuAzy6N0P1
TVOyPGTfeZg8n6Dq8FpbTh5DZ5N8ynB8U/vS9zWTGm/JfxTQlNmW89umxM2k3GvpJSrgSyuVobtt
xi4ofZDt0H1H5AlXLi9HnI2DC/gup7NXEXlMpKimyxYlNQGacfa1/jjnDyOFmValbwUtinJnBIby
D5DtTPl/0feFcNxM0lzVH9it5k1ytse7uTW/l+QnjNz5OLwGN1toDnTQric19Q9CbvXOv1MT/F9w
I5Hq8VZdnDsSCuKhTy0s9Tc5BjJiTPPWCfZtgNFFWaDYvekHCIse5OZAe0rGUaHk7MG6E9Q8qfFB
S2vbqoAl/+47jUR3a1RudQBgkNs5IEi4nKtcyXvAQ/peoR5FwAagTElGxbrb1H8bV6k+HxxAUGEM
auDxGygR/r5W3ckUBzJjy8UMkBQo8XhhTyGEQ/sMU2T+uyQYBN3HNETbUKfMC2ydgqu+1o1AG4jF
n6dCq2FwVZvu3dFm3+fPylRiY/WQZFiAspnOk0ujbIlq7JLkZOGtNnjl1HpuXzeG10AilKmKzC8/
+UYLSnhdlBhiIXDeev7ESqaE58kFJCO6ePtB4uIuQavOwOFbem3LtH52p0fueEFonetxJrDQGIM6
KrLPH2akP1jQbqqfI1WXauhhsvgRuh6IdjLzQO640K+Y3KMbHucm424knE55AI4hCozpHDA2iBOX
hWTWZ+L+UHJjGxJHqqbS14XBBy5GYmY8Lwesl9RQKNejaLt0TyMTcNptqNuBUyiYJpM1pkJnJL2q
ZzYKBjngdoKP6y2mf1KKn/xz4lv/79dOU+m5hJASZR/mTjC2qvTKaiI9lmNTkPPe6kKZIDv0yVyL
RuMLEIfOe5vwXItV8xVm1Ocsk1iO9tiJ2zftLGErW+fzyEdxdJzpTBKFogKjtPECprbtucUE68Lr
AYEY3NxEtOPdwcI5w56rgLUVhjZlwmVMh0nSnleOkIFCCc1iWSuHwWKtACivOyUhgppz1e3cwWDx
1z6VQcABV+pCOEOF9M/Hdrh8a12IoZGqeCqb07laFFEuka72yWvGwEGq2AHf/hdiZrpg5rtDpilH
2yT1JlzT3ExmN0RGn8piGa/IwsE7K9/LEBMSYTDIQsc5elBIVmWMta+2cqY3QBRmQ4axDyDoJtK7
/hMSqrMrgF6QsVYBPoG4be7iI0q5q3vikgxordFMG8Qw5Sa8Ruc+BTXbTY/hSj52/QmxPo6NsXo4
ZMEid/OPaRgUJpdI6KBvb0yvBHLlLqOaXU4yxaQ+1YnU9nEI/C9MI3OInX5/d8T/hPuwfOl4NegD
zdLdLoDJZyR+5OPMkrIU/kTU5xQDw0QLoH5EkwMqSZguvhFkDkCbmBpafQOXEoHl6T9YvtwQjXEw
PqCvq3CPgkoFiiUTlkAp7rjdZFSRFYep8n0XDUnWz2AmurooRdejIG+8cdgkPd9cWz7k1BJRtvid
9fJ2BcICwf3iQADQ4AqfEgg3srNdCbIesN5ZfOAoiU08aNFDRaGVSelfysScNwy7Q9hNywFKSAWU
hkw/opUIhBOFyvmMNWVJ0a4TI4WrPMmd3JOt0ZKO38M4AH88ua7kSYXrIOHMA9mCD7c9CEPGzXwD
BQbRb0TwlryLNFZ3AMPfk8hU9X/ctkbhWcuxikCefbqFC6+A40NFDXVeP9Lul0/b7T8qtD6am8rA
iSD5d+rggbXQJyc6OW4dK/ByaYXbuYQDETzOp0UXLwILnOTNvYdjzMrclWkBGitjrWWhjC+lA7v8
UcoThiyjw7eGA3YR7A/1Q1rPd26ZfiDmPvCUqnarw53a+McPqm0cj8r/5QFBrNceqoUkrTI3wxaa
2P5L3v2eoDcKcGC9iTqU9ESWSJzVlZOqAy7J3ZXW9Qk0LqB2N5wI/BfQw4D0TlRn5Rba0Jzg9S+M
O/Uax/utEdkVj1Mep2gCgTqWtWzK+GPcIFdPIL6080BgZUlirzZRlW8WCpduXjRoFvB/wxOM9i/c
i2RFOUXXmb+80qBysTGCPzqgxtSKZuhx070zBeAlJO15QEyDRzijqnY3/jBoDJfPE0xB0am1KfDX
gl2RpiWE43qrZeGgP3osZFj6er6zTkzzwH+GAaFKvL1Su5OUkpjcmcIu2Axlm1odXSdZJPyxg1IY
RYXKk8Zh9s2DxToH7XEzHF0p5lMktwv0DyHorQ+5I0jHh8lEGHP1EOof7ip1ZR7EwZyNQYpsErsh
Xbb/oqzDLyVrgpZ15cGBwuxEMaezVr/MX3EpfW8OdrYhUaowzbU3Nl0e0Z95Bgt04A5JB1oPzFYk
c5psdcJaMRIqIv0K/UD2E69EeMP7/ErOOAUH7ihehvIyM+RKi8hceDJJE2EM/eY7+bL+j0YYdOnj
IoAOsP9NNc3uRZFkcgrsnEvRs05kD5Cxqny63ID8n2chvDiMoR/h/AP7Y6x60qqAs4FTk6NWOmjj
GTikbG3O8EX4wr9bNSDkjKx1Aji+2M9h2ulrdgba8L07TalB1pXo/oRIi6YUIOQVKTvfW4yHF4K+
0ygOHEBv3t546WS0/5f727K64kQcKpllaodN4bUMMzMfQT+hWN2+bwsdWbLTpjsm3wjxpUJqC0YY
W/vg3ErWPJsqqnUrhp2orwYPqI1iH2cLGdNtiAenTTqNYj8LOMf8QqdHRPjUeNnAR9ojnUTgi4Zt
sXzbn5O9StRxiO5P+2p5geB8S3WxtfbExhu83MY8+0AMqaDk8xVyWwhRJ12UGQ6D1ACsjokiNFvs
8q2E4k9PFG9+Lv/45c478XkdDyoMKtJ4gebq/4+X56M9kmDwU3NkhDDnSvq/MhkaE/DfZlUgonVc
kSJl++B7GwymgbkYMvRMgcVI7vupBo2XeE0jG3Wbs29FUhUbHoYPt6D8LPIXrPTbd4jPi95yZUpT
39d4cRrGPPbfvOTG7YlhWEmmZY4TJ6FNEhXIndyVrrgRtIoOyPy5Eu5tRDoS3AN4xTqTmGJNgf8q
NLHQ2YXOwEqI2C372ocfGNBIeUwjx8sO6V0Vs1byBTnimAGtHfHwqzOBij3SSGV0HRBfe5WAse8+
gH+nFn9NlXmtCMX+z5NMLB1SQMev4RtLnetZLlthTBEYXgCKSjLwFXTaznzmbObnmvpvVpscOsHQ
NYcen1QFWXrUE46VP9hCyTL5+Jizkg7F8Xr8E0aeGdv0JGnMcS/S3iW0k0FyKI5ZLKJ6LipY9O1u
/wPwRjVyjDUSsjBbW5dFXBmbtddSsqyyFmOSOM2hMs4XpYumIfAp0ozoqz14pdCFIWYlMdWc/MuQ
proqnrx0lkUkRjWtFrJ7q28+KYkiBM/gYDU8YxfWDAoK0y6bFZcNN0qxmzBnN8bL5AtgNqY2RoBf
wtnoslbrpnl2tUxpQmCyHpE+GLgc9dZ6FaAbrbVYgMXkEfPfOn3AyKBu2ga3bnPfylHOCZSBcLHJ
nrb+Njv7DOFhZspkDWzgGyuUrSII5PSnjgXBT6K9NlMKr4c1Mgg0MWUgAFKdN9H5+OXCg7tZFyUb
O9H2q/ax+zxzRP0nx6FTIInT9PTNk/pce9i71jSmrGvqOOQwTmTB1r+P9w85Dopn5xskXi5RQDJz
XlZ4MtSWCeu+aEFDn7GyQIU30L0WyCqn5p1T/hHluykQW4nVkWv+fcmNmzthoJDmhDdjvjI+JQQZ
Rq3g+bvuRriEMwyyovxDtO9FTlqQdBXj0SZiKUqoD9UtYH9fkkfGoxJJG4pv8hxvC03a6F2sORrq
ADvDhaChFEoRl2Kxd0+Tsfp5uhIxQsXAsKg9zOdhasDygoTp7WPWJLmnZkQjoAeHvN2bIy5R5oKG
dKnudtf/IXLAWIFM0AcR7ptw1CNPEQDxpFUtzCuptUe0wpqo352BRyw0NM6EqNAjxBaFHO9sFDOZ
pqP+vNbBhouVn8VdgeMoNNoj5fufSAMjMsbs+npFHnzuzs3juXEfPkCiUrn32PPsUFFjWVJKaXI2
JC6RRx4WY42CJMN/BqEOdzpUMvLOERmXtkD2pX0ICF3TDs1i0NhZw1hEJ3dKL610cR3AzObbixeh
Lmqzmw5IdBZIh4jlYcHxdLrwY55qHv3qqjqlthrbwBB9HpNZV0mYMzy6dhzeRaMxq8Tje9VVuzBS
2jAofQqkGsaac7+qjm2E6WGeSEvPNSH9/iZCoMOD3+cndn8fARPHOYZhWWiw/fvi2zyRxkM7jZbi
oM14walHmuIcdjQk3qgEABnvXwCUqkmpDw8uykdwvpOeH3jOkjrP9HmX8EoPWC0atdd670XgxvEL
l9x2tVyvynjNqcVqzLC2lwh54/i/Z8nLNrEjMhRixnIDhkrP08r0h5s9I2s05HZti6h0zIfUIK7W
DYW/IU0l2VNNVTkA97RZpGT8l7du9WejPmQlAVP7KrT/CNpXd0STGNqLRW5pABakxSEZsveQGd6K
nknHIoeCQJZgL7gYed47MnlZrfbtXrRQ8O1kR57rtaVQFpJxew4gRzLsFo76oo+xBQRG/9ZuKwfn
ezCSoDqcaBYwtx7oen8BQE9BQwPT1k/CZRg6HfMWlAjnwl08adagDZQFGc8CCzMO1tFznNow4++R
mBbPjrYZeaCcdxI+qK4FINNB3RIX5fWHgyQUq6PAp+BQBGBEwU83atDEXlPTIQc0iEJU6beFdzPB
2o4s2twMIsjkDqnKic/zRhFLBERY5s1j156378DKDqaHcrsAn3KaqhSh7Z7i5OuazxzfQWSw5p/5
Gfr6XvVhGmS6TWdWw5kTlB3pXUnVPZUxTF/QsGUY9ANRSKN+NWG/0Qp4GOf1cd28o+KTKKmIZHOe
AzNBBYok8wy02MbhNUVTvNVbmfAqiAH2jSnTtugU8n3APrJ1FQLzIFHaUPcKA84m5yZz0A+FIJB4
Hxfia7zV6oNlIFrp4X/F3pvDzxfMOtpnaeWJkUWF3fNkuNTKxtCPXEEAHRd2e5MPaMBfisVSoiPR
ov11Y3MRSgkIFE6Lax0b2Bx4IhbRkJeH/ZN9Ww12pgFzoLMtFfLWzOsR+sqalusdj3z857l8ngOt
loO53skM1bd0seqvAjCD6oQckLgSUrJp85bSl5xWvLjqHS/sxSKvcCyzKoCUGhSPjKsX/1HiG7Lf
CIK0BqQaxkwfeIxVtilFenD1IaBohIqHhP8xJdyg4FzfV0yn9Atjs1qU4sCE4SCl0JBknroievEY
ejjG8Tjd5vM8a4u/3EhL+DOR/YUNixoC+dvh/7gvSyAZe4sVpb/ZgOKrvJvBHyx4fG+43zSNS3op
fKxM/yh4deIqysO7OQYSfkmOyPfbhGdq89BmIBlAy2QS61o7jyIrvOm1Rc3Vey9c7NCoCXE6tfIk
cD5Uda4sDlxo6KVuf3vTA3po+HKujLC4sJrSEseyz7By+9YG1zMqqVwHeuw0sqE9s5mv8ShsGjYM
QWbU2cBkhFwBVI2UZu+GVPfrJDHyoohVsRqNXeJ3Xo9Ofvm9OHwaFGxeimv1XuFQoygLiOp1FB6Q
DXzA+Y8FyO2el0ErsUmVOHpaeeFxJs3D+aVLmIS6l1mLLz67oa2FZ5FQIZ7zLfQFtt0mOZPpg371
xHbcfcskouH/fr17koQ06PMSc0Tgc9RiHidfQdgQ6fCVj0h6HWOGDeJsZLbzQO5eEVjpzThZShD7
ULCmL+H8Anm50/4TsUWL4Ek/Co8ZJlbfgdEm2PIgPQZJnbUoYYk+kAg7fKJ/1N/Clipr2apuiCHj
dH3GiRbVfnqjGZ6hA3fjHbiPKSNocB98eFyf+swrGV4jqYnDD1JcMst0LiqIG+wGiBNl6U7kA75h
EjignLLXUTH/w0nbsUlgHf8DdWEvJBcnfWd1HT8jG9KQuCNfdFDqoatHywh8Ipu0qPY4DtJfwzxG
IlcMc5WFodW69R56YN+HRcJ+G0BgbjFXLFvN97KlpXKD0lK3KQLhY/RTOD0a6kVVwam5NoUFY76v
E9D32YA0jwA0L1Tke5pTwDkt6RbkD1O/trtPwla739/tXhnkGwBszojnkKEJ3yyWK6PCuCt6hVu7
gp3zp4mkyvyTtycvjnjglXrgWxuQJe15/VbY7oYuitPwt3Npo2C3i9AT90DcMGJnyBbAP8anHjzv
Dot94zosQ+3jak+OTzH/p2ptzrOLfKEOIo8MEwPVMaUVx7umIKRsXHRb0YADFT/u88dIGoaGJAoe
b/RM0AJdsGNS0JeSdNB+ZJv5pJNBeCyUcsHBJUHy4+/p5sghCzBk68ySCT60RDXjDepTOOtBkMHA
EGavnbyfYqkRvswmJevRL/5CzO8j5hdksBTdirGlVNEPkBWe3GHsLCkSVIzFdcxCaY0yL9RfkGzj
pIJbkV/03I0Aw3NWY364qDwkbqBtEx1AKOl8YG3IhRFGjFlucmpS2sApMziw4Vpa0a5N4mdvEtWP
SRabQN1XUfCgyvsbWREAwIl2OPKyrpJQOWEnpyPhw4tLokBwDFDFEYWPVrfE1b2G1NikRkA35ufa
jeWMdFRv98ZEITzIwt87zf9WScROI+x40Y+odbL53kiAH+9LFm1dXClZaZT7T5KY7kNNJHDbZTgU
CtuO2rB6M4OnZCYXDhXoPfu8hdM4zBBdV9cCqbEdShCo4N5rMaVj4z4ck2aO37QABnXdgwicCiql
2fZRwTQzESLwzC4r6xpL9vM+9qRedFBDkB5PzJKBaEPPP+ZxGfUaZmBSRzggknk4bcwe/A/eLeab
A1liTmVr3eXGROCj7LhYeuXPdste/OQbonDxBxVSkSarSWhV/ln9fuTRLvVCdr/flinP8O5smFO3
EYVBBAw9lklooNxxXBsylzb0lM9KGJKrYdk6nOkPKG46m+YK2Ae1Are4lOOm/wftfZs++RXsFmEz
qoB+kfDhb0NgGo0uWNfymg2RlwyOoHp3pz8ie93BZkFvOWlb5s3yAO9j3m2jGek2ou8tvWGSiW0Z
+dl9EUW2ZwzQU2y95PMrkBOHAsuqNTocSuwB12w568wI3TZs/UxYD/0Br7wy46x1+yUhwqoW+fLS
C4vQKSwEOJ42eFONApGGf2o+sPKWPNwpQIa0QTgBfVfAvtT4hFHdBVdFvW2KXoa88EwQ0ERKSNjw
VpfU27OERudD1iPUKdoNzEHrRCJ4ZIcsK6DEzFBdjYATBQwkLB0otUBbM23nxLys4pCa1Q1vQ0mw
DOS5IO2raIpfffgvQw/PQnLOKVtGa4ToGKwfcua2r7RzXqsAntJTU+CQ4mfRzW8fbwOxtEdH9MxM
GsGxaPS0UN5lF6m0Ncxy4P6I+k53imKe42TbFSm9ncFqE//hNH6xqDZcjI4S5RO4plAk0tG9MLv4
jJZeQFP1DbkrsHn/F09ZB8vsVSOVA8ky/X/jkQlvmW+w1MHMlQUCTwB/c7i5aH3MNp1Gj3L0wl5a
anZ9sILtUxh3J+2d3ofdYPdSjsRN4NXKTqXgv5YmE9oz7v17H9tAFz71Xy6IPwTResB1LxeFRYI+
tXj3wF+21lJAdMFmvqjTC8ezB97JfxF31yyWAKcV1mVDycKTWjeckOzVVvXs2bTVwGUXakO8ieP2
SsTdUSLa53/ywv7YuHL5Nf68/yYLyHihTpLnkXpX90komO0XWulxBg62aO9FyaogE6xFT91Abm/h
Td3NsLAQLj/d2mLYqj0kP5l2Hau9gWEnjM2OKdqULk9vZGbOci4bFw3ZX620J2MMQcm3M+4gQEC7
Sz1G3nGlkJIBYJQO7im0W8zv6+T4Jvc+qobF/k8zJ5c79QEJuk2tPSDXUcSR4vLOZgnLDX51DsNk
DMvm6MIRetExhtSZOR1cZHnIrGqZjQCXZjngR5SVhxHdvRd8g6fVaxGf5YeiTy4W4lRLK6cI3ts5
dbwbh6W31jmNL+9s4Yx929UJ5R0IautspiB8mKbx+3YL6X/3vLz3vdTaMpJPYoLPGsr8gqm50spK
LB2CJF3BaJgQDFv/2HgCxmpekEjRhQy7BiBmnYjvv+CHHT7YaD0JJYuDYsrHfeB7u4hFeKDZ+A2+
bG9yhijDlcM3rp1ipnYA22t5sTOtix9ZCaIDN8BfGtuoDBvRBjDH/LX7fPtC8seEG87hMPLufYvz
AId1mrYbBtVsyVovhF3K5PLWkj3O0SMxV+qa+7dAL5pvaeH+wf45cQlmnI7AQyMo8zvTDOfgVQn2
9x8WYtiho6IJ5R5ZPrd7He2ZD3s8wacuwaHTu4Pe9D2agi6M88Uat9jR9y+qKyx65O8IbRtslSIz
PsLOJsxl26F5eKL1f1NtbjAGLCEpPphZyNTkaPYNBrfm4KC6/t9699VUv8NeI6w4kcyYMnFOvNI4
tgioXp587ECHpZl3Id2YV96/hMhbfceEEyCQ0BBf1/x8APSplLl722QL7/hnqoRC3QHnjsSDhf6N
nXDLjQaESJ2aewASNiAG/YTIumjvwa/78ibIpedHBlgsUsGBInrskBu1cm85P6kUuYYSjQsflC5V
NQx9EUx23UjJBUTF0YR/siWMVZ0CxUIVQqfr9HFe9eojjCpEeinFLFo6ncAxsShUh5hBG95gXjpv
6MTd7pB81DuycAJUkh5L/QKpR5wSj0Fx8vdASomatDUlEGgsC/4wlOvkdODp0RPUvi4cHl2cBxCt
gQ3sVXWF5RCUhJMmk7pdh4wQamSivyLrfSzc+Zg/f7QHA+GN9XzqEcgfqKhxXZ/9l2kubfQnCddu
VCGpi/w4PQyJTo/apQUvElkHgV1DKkz1y/er+ITlwshJleBq2FuyMRD2zMO9I9ci+aajEnlK2cMn
68dmAanV5giLHiZ5PnkcSd7IehYGm1cQ2ZbrNK2v6lQZdsyq9jy3nBFuUBH/cGjKXmHVw/J7XxaQ
8aT2w0fI6yP/2ALJTGDdO7TEeJv5TAnIZQdAXaxHhEMpxIoDDgqv/gOXGv1C+juSsnzU2UxNG7SG
fcYpzKbEjV0B1+tEVtdgetx8MyVYzbPDSvfQbsg5slqDGFdzZhqUEUxlceudPUlJfAb7G4HMroc0
3jKI922LA2tWYOHvQDq5Lk+XmBoC+l8B+Ylo+j5jM7D7nT9ymqRwSDIEjt0vsbXvQY0Yao5HLzpt
8UP8nIrbKFt/bMyunzkXFJD+Y7Qvz/tOd6CUZyU/EozV0EPwhQaRq/ee0rpsrhDpefo5NnK9t91x
TEB1IoBCYRIt1uMYt0uQ7JFXnwYEuKMUVZ+tf+drn56ZUfdde7PXxhGzM7ATODyaqENZeZmOj/FQ
fBbo4ZpJuaOkjlPSzeyJGkwajQjjDuEKqNF62SvJTDq5u6HxhI5/GxRR+opu8ENngH51ZgIv06rO
AQAOZ3UDkrMO1U8ZcPyc/nWSQPeCkJbJSMf3ohtJhl48dQq7TFtNKwka564IEwxP5aPHliABkTRQ
3aclSpx2wdC9L1NuMJgmIDuDZhah67GOoAPZl3VaRPuB6pDJSykl+As/cmG6Vgymy4cn1Wuf4s6Y
Vt3ErfisN0mAe1yRmujGLOir0d2OYZt6J/7YuC8kwzKb0mPdylqqXMe6DJQugLhxFWt0j9M2JrTp
64+QsV4ANln+8TkDJOXF4ucNEW4+xCaO7HbxWecPuahAlZ0fhkvzX+N1FiHdc48shLklTCS4zKze
mZrVfmGk6IjViA2HI6UJe6agrih/k41CcQILBqjh+GEjSQLTpnDeXDYho41b0VY/B2coNgATg1lK
mTxGkJi0y6DZRBfkCpfXLzwwGEp2K+FnOT2KycnrvHSn9bP95Zt6ztxy+qElk6oxOw4SGIpIkwUV
5ZIGum1WnJlFWJcVlGodk4wIck+d9bRpxVqgiEGeNjck3LQGRucjmseEHI2r/LuysTht6hYC9st7
KK5pD9nrsZvO8g/QcfPVnEZFe6hT1iphP8tM3yJgK+oxlh1gkCkTqxfKs1RfzImTPHlfs1BIi4TI
2DYwjsp31EmCmGQa3bb9t0xAGxZQQiQJg7Q9TBKt9UyXsOS+/hMcxH/sx/oN09cyyUgSEpgdR79L
h96koOfdNCwhjVHpgHNmqBQIlJKBXEW/6RlCMLopu7WExZ9Sk1qE7dud2nWozrj8adkU35ZlePlj
8dstdVBmtO4vebrrM4IkTJkw+G7RWflqgvBItuqpdPG34jtcBm3WKtkZqT3zGpmagiUPjyalEI3U
fkv3uqSvQVETtw2h2KEYva7rwjFQEuwUG05uaTuaU6tMLtAFKGKkg4PiuuW9n1Pn7iYfRQ+KGeTI
nSMY63Ycv8TR3RrnkoDXyFz9XKAm/PPyMyFj9x27kQZBSETs3qclJCvtTgF0MFodZ1KxjG/MZBCH
AdoxCf9UOMigKxW1+DQxX9mRyhh4IczR9ALbjRZAq3oT2BFfvckyg7QLW2CZ8jUVFShkREd194Og
L02N7wQVE3wD6UFZ1KS7nto8e4HaXMlazNUvnclVvgoYmpEJdG5mydr0ViM0wxlQ1IT7b8em68OS
vxtwxF8tuq9d2uUES6E2ontHwkioC+G2VKKe73+emMK2tH99jYV2YBdpxScXrXytivtMiYzkKZAI
iYNpiVVpvrSvGhghPLYj+OxhM3Tn89+drc+luRF3FZZTac5e8k8dDAQ7B/CrOWttws729adcBb0R
hE/Z6s063WXVVssP4JtF8ewne3L4RfGsWitlIegvtG+/BX7zhOWJksZGLbHKcYSvHqq67Y/gRGUB
RjDENrk4Xc6PE0nsdepLMtt1WQ5ctMRFLWEfsf0FzXxTLJuKqRouJu5BuraKmOdsRD8IM5QswZ6D
jvDSbsqY8T8r0uUmUu2Joum1kPIFybPpsnURp2fCSMX9Q99vTTu9jxKc3+kQB6b2b/XlwPXa8iIx
FOAxf5G4ln5FAZISrzgAWG+pKO4feWx+qDFpyVvROImZVqxNRJqL076SfZphe7BjK/nUOwciWSqH
KJdxttUJIi2X0b8zLmff1E64IrkxrCBLBj4FTssSLRLiJCsd0Dz6/PFo61jaw/NFjqHsHaAMgcuE
gkbfvaPfZDvzqLjfzHBNsF22szLSRfcC8Faj+g986J575SIr4l0gh0WyBwxd7z6wiF5A005vUvcK
jHzHGKuTtedOYpMPAg62enGMAIj5f4VMthGoT9CtSukTflVLLUGovCNWjUrOORkrckx2Wvjaatp1
cskg8Q1Y5E/Unv6ttsJ3esMZILIBjWmZiiy0qVUddu1IrkDs79YSzR++zcfmp4RJ4IhFPeQuM/rC
0/f788+e6SkxGiM1J3P0IKyW6uHhzyXZ1RQeAWUVzUMaBQ/B6KL+0UvLasR86dWb/NqAVZoKrw8R
oMEKQYvmHRd+lKvDgrVwa8XdyHrh/QCdVq538ZKDlZhodYwbmFNgO1TZnwtxoXzZ8diQ9FlGoV60
yKMWBksjFMX/6zMIosrewwYY1WpmLquAnmYnm+9qstvt3mJ1L9a6uxbCHMF5zZ+8UNodIpeMew7g
YwsmL8DXetx2Pttt1z9jsFB7fX/IPka4g5D8aXOrFOtJSoHe7Oabue/3+JxjuQ2c69HjmLb47OrR
Ub2jurJkgowj/ZcxiQxe89awTYW0sxGqkNZuxrrIqZZFw83u7MgNOvGC+2UrRTQV3nHONc4BYSBS
HpwGcFjdWALqXWqy+h4gc1/zl9ZZRzyVJ9Ku3qSONVr3IUfkGkwy8ptz7nRzPRlA9wcXdD+cBc9t
zqOFwj+1aoSiRpN8ONPt6pHu4R69pdhFE7ip3upmy04YPrnQeokkDbUpwDKL1T/XV4GDZgCRHGq5
jiiFWWgLLg1R8gNEjkkbSpiUuOOh1dVpGSOOG3q1MrQ0Ss5KCQ5FktHvPksq19Xxga/LuKiyditK
1eIuQFbz8aKZn6l5Fkf3/bvBcAWFDw40A7mK837T9S5J5ugouUiCuQJs5k0PC97p4Oh+3DkpGqRt
lzUuMvLcq151OdNDGsgZTCy8GeVv578xLn3U8Z9p93K4KHRF3/A/yl6OeAOps4bYR0iCEXdMpA+d
Szby97BcJs4f+Ud1ShjjUzBop9rwun2MuP4pG5qZvCVvaPw2YLFM69hMT8XEOjVAeVJ1NTD77+dX
f86ABTp5RTW8nlS80khKCLeZ9zOVc4CcKgFRxj6XdbfZMbzOzmXy3sawxDXluAyWNRLr2LrQP9WZ
MrClKyB47ZDSlJmNnFTB2Qb494nOJPOVf00PIBKZubSoPsA8JDM96ICnw0SGG41XPGoXKCSOFAao
dkQsLeIog7ngM8eIWJsBkz6GIqnZB8KfycAk0473hlWFNepC1j0VsBNToGAYzp2nVMaMc4+JLQe3
pBuc6+aZjwiZnCY42DvuUQ5atzPoeCK6JWl8sSI4l2km4lHGACNyu5nwAnvQUXadThUgw/C4D68A
Dx1jIdNBx/vNpFlr5xeRoDXufIkeLeWgWdKpSy4zqyY28SPPQrvN/hG2Y6+BZetQgk6ugY9t5uYI
YAYFIAuATFIaj1vZedfHPWZ6xrQbl1qhnaFRpyHGj/0vFT78mYJjvP9RjMREVkbkyQaVcxxJYpAJ
DUAN90UPYNM++aNUmINcZMe31XPIBHgphTCK1bcT0Dc0VkSW+LX0EOieZaEfapTE0uMJSKC+3HGn
zzeJy2qxny5vtUpAnPTCSZSKulvtAW7eDt6ZjeLViqZve8O3j6GPw3l78hz5BywfsB6eIp5vXBMo
giF6KUh7tqXEF8uza1zlJ88GjYnlWuioJPKeuNHuDnG0s2IQvReq8UajX4gGTLbpV0qVbt5Iw3D5
auljwOtJJeVmGZ5pzGvGEqjdwCV+Dj7S9orLOXK9P8h6DtrOCMO92jNGNXDY+c9U1RFii7vM37lC
wIQT7Hf89ypcxiOMqTztlXA5IvI2eCVnGEQxRjynxl1lfgOqR5bZoxLtSMo0lZjLK33jSFQbP2R9
eXU3gWqadMyFNnOo9R/OroujxVlHdhuIPncLcpe8GxhnulhOnQSvHsdq5nF7jQ19m2OV3r4p6Ysw
zXl7dv6SyMy0AyOvaRPv4cxBKltxK5flnwqvoSVfo9B67eIiAlCJrdlM6Wcop0vbt/fG0h6d2cg/
gwyVW7QujA/6f8tlbgVqZ2HrPSDul7B8ZmCQCjYQyxNprwHTL/wFOExE2IkYNdrhM9ttj4XwAmS8
FJoCwsuyke2aIMPFPc6/CE24I9zm6rOR1e6M7ioPRTVuRZJiNKlAGhA5aK7SD6D7cc8Du5xt/8t4
AA8uT1lfNGpXccCpV7MYdb55xvmzjNDeGGjo6MgUZ8XM7v6fS/pnN2kPvMTuFrulReWzxdoII7ba
8XtqTlZI3LqcByBzv7S23Z7KtrGiy7KAXSZhJnpgJiAd4ELu7IGmbx/R0gvRBtjxzvyD5taEp3Ac
6Ih10oy89Fb4KvnMWMXyf1CC36/a/+WccWdZDgvFlnbL2ptpCZfUga5TRs4GNUtuQiDiFHFWVr3t
jjDkHzYtLXtg20spDkvuhu2MiPNagnLkxo3UUBTE4M54peDl1JyV3Iv+LePx8Ok+m/vbQLVauG8E
6KT2D9uNOB4g3brf2HNg8Gl1hjx195Xp11L8U+tUeeo0CM05UeHcI0+Xbqvto2d7ZPWFG7UZfcG2
eyh3xyhzY1WgCpGgoWXLhOET1JPaiiYcQ1cB9Hx1w4ujUF4nm7TV0/OqQOIxodFD8nTxU7Z6JJBk
BJlOpDg9ppnjQ0HGGGmTI+Yko46LYwLdmA0wrwtJwxbpkX8zuW9umfWz+sXypgjggbA+jVUh4u7d
B1hH0qrTkdFvrC/er5N1dw2Ph58gkGYQAytRml3nZgpRG8/G0oN4R+Om0vrAa2g0hd6km3HeDKQJ
5kHnS1Yy5rZBBVcwhkNmyINhKF3H/6JxRvgSKrUnlN+35Gx3U4Pkq7Gpg8k1XdtT7dKKJPvLaSiN
Vsy99btRnvJ6SZ1rLKYL6ng2RjrvX4KMRldZI0CwHD3Uy9Vf899/RvZMUQpQAC8xbttCJD7ilEAv
AganWy7ZmOTOiiAmthbY2LAEM0h+LX4I3/YFal26RLvuXyA9QflQF1anx4phW9OWNP6edzcGd6j6
w7OwsxRSzsdK3k3ledsUs5pkMIlp+5lbOJjX09YwVathvACbI9ZFpt0atmkBffzR5xO1xXQHmxyD
Tr+Um0CyttliD2SpxFFxuQDHDbW0v6ugkGFuemjQQu3b3q6pRXMYIllogsLA9xLoc08/88i2cKBA
jioU76PEQqyLhQWV351G5CELQ/JAxwwB0IX+mRnK//LEWiGEN4k9YTtj61qNypG8SFVWhZHectoi
pJbqrT9YOgMYA7b4CnyZ4k7BXqkqq8Cks1hH8q7KWWZdjkiD9n/D+YR4Rxj6G6sdKV36EZyJNLaS
yeTSZ0N+nYvAGQvSHe45zdl7iLuKAJb7hVKaE4mp9lv6wNWL2fV8Lf6Eak8HyrtYxn+Ns/ix6pDa
1c8fkGl+pEMbMYbX+FZ0Vx9QVMEwlcFXVDt3fWY5Fh7+ChqhZXY/LgTFePux21gzc/z9wkFQ0RpY
GACSz0MpSLoknKku6gtDJy0BJ17zJelBTgqCeWWyv1F1INCvCw8rZ1Vfeq+Kl/Tl80ZTwR6ABJnQ
Na7xU4ngKqlxsGZM95Fg7d7O+AQBOii/47NGGPIett0R2VVoNzVoj1mUZYTrbmYLzcWaShH78nhR
XljjcpW1OMnC+xV+2DMLzDaOvDI9zUu4fP+OAsOy5LnAVkZH0LOJWyBG3O5T6fyrwoP6YU8dlU2H
bo6MeGXr2HQGhQ0i65P5OnLqTF9lm+Nk/j7nIXrPjAJgybpoCpvIch5ls3i5QcoTgklXkkFmp4vc
MDy6xQxy2UayEJYPEDpxj31maOYTPd4wY/U9qhcZqd9/vEeaEw9V6lsvcevLAc5iwl/bmntDYZT4
pr36Ueu8I9RTL8bdkXcdmdjHsSH6DB2sdM8D/TE454v5cMEQCdMmuqLaSqTpkMWeshxjzhWIHA2o
fC6QgPn4HtvtRLYTkMCB1zqN0blpNLhFshFRcFzmLhv5llW5r8DkXMDGWcUPxnwSYtByDIn25Ids
qRpy2MztDuJWxSExoNvMU1l6SlEyDIcXOz4rl7cmAZcdIxSc2Gg2VO2OqQ/zxNl8Mr9sbJTSan6E
t4aX4I7Nrb8KO1wXrGIS4acaHLa0JmuEGOthznKs7jnwZpj2w60heLmYk7zmayDOMOOvW6wEDQwx
DuNMqDyPu5nTGXN6SmJDhifsQjgvANC/r1Klo0aRlTZMwJhAH+9CY9Zr+Z4TivxDQkbj3l6VKDf6
4Tz2H/B+Q0hrRGqgm6TowgJNexUyoWGLEOeGaQFEjU/ZbJsG6P3DBX4jMqHehg1fUsqGi4Dygu7S
NsuM4KXY2UOALiDM5VwpIirQeqlQvpkxMCcCps6R2IeCAFn8Yc6nxWUG/W8FlnZcHL1nGWHxeqw3
NUCd1PSsRAx4wyjDEVYgzkKNiZKme6GC7AfcApAZcMaXxtdVpGUKa7mGBUJTcSL78wYyJBGu7weR
M42NNY3Ck8Vej0GvIVISzAwiOMHxKMk/wKUCOyWNxVSq+pq9AkRvtkMOkIR7L1wai9cN0L5iJ1hC
L1zzHbUXw3phbi5QopiEJ3PwHXhp9OnF9EjtBr5a3Lu1ZOBUFXfvdEyF7VBtsHLYEyvsYa8IjiW7
Qoa4byZEB2Wl0Af9zGDOLQebqBNt1F+irzJuowrk+KeuKtSWKdvEE/Y62A5W2xslDzL6K7wKfnK0
MNG0a55wBqhp4Dz/AXcsIqz50rDAy1QYxhZeMjEnvvIOJTMJ0sJH/4lqYtjNX13XS77Wbgj1Au+6
Rzh6fQeRtV/lpeM4+ycVAf3e9Lq5a0WS/dVxPH7n0hhBgZBI1I6745Eytud8j4MZZhZvYdo9b+uN
qVEz0CIjdkhidjOv+BWuROkHeiKXaCM9JWjHoIAg8j8S/WiafLF2q/AtdHsqKzWDusJaB9Opy3ss
BoJtcHLEULMLEiFO+rALnXvYMti1POcwo3MpOVd78047ZQl7UDkGydfkjMCTKNLYZwqkwgy1E/tE
CuVd6vsCQ6tYzvN31+bn/9HDFzfYULUeQHOGC0S3pSIJaGMTysN3ayvcuzC7tn5Pr3KEVBrfsOtk
y/pLsbtxeESX6Qw9kOt/UvzxV9AeYIHz/Gmbr6Qkmbe6SVRyXQm/zxArj1+I8NjWJ50lLZ16xpre
a6/vss0wZHgTx5KNvPiSlh9Gzz/POeCdH88KveC/ymVP80ckgOWf1sjrfiFtPjlGRMQcLhNDqSvC
cOloWRQywyXRJhgXF9O1FyCCY2XLSB0xy7ymaKAVrlMbiZWOYMAQmX7ChkxO7rHerxBVf7hNCd3R
U3NwoFqs6HaIuyugHF+WQJtyEJsFx3oeXAfecs128c4bKxvC6ZlWABLx4aCQ2aujH7c4DKa4d4/R
AGhGTZPuQzww0DzYeWby4cFI13oNDvk8cMaTc8N2NhFJrEOiFjp8ewVhuns0eJrjiBUaw1TpRgJc
WK4WuZDgxY76udCS9QFg/HovQEjBiWruiZHhdaENsaSHnLrv+0quc1TDBjH1A3v5k8+Za/6DbljW
nFJhx8U4tkdjzSr8wwUHzlFeWzw5TprRUcg6BHIrOLfGYY2MU4LrtRvc04HjYAiS4lWyXLfsLVvc
YFFvYA8x9Ofm9ndKrMZgETzA89aShjOY+AdQCmmmkEqJgwrtoZdUer+CRdz8xbhbP1LdKHDw1vIE
ZTBopTNNOvCNtVFaIF8Ab1sVgNQ3C15sgaq4IoAF/YveM/93KeLphbz4w6DbwAwlHGUYYT1QVLlP
yI2aREMMHmVLuOfupwCMOQhIddU8n3S5QZYD49/Yl0EPjlA62o/i6NAeMchpJCel/dPCKBL9QrD1
o5WN+u7SDBvW2wY5Vx4tGon6OCuYTWx4wmAe384/67UQnYfr1Tjz3HVAGMJUU30FmGGO7FowZ736
t0/JlCtsyNeCK+RD8Tmo576z1zJfyet8Y+EEXNKnrUr8xPQNv854xQWfePEn2ILKz13ThNmmkfIa
IJOvYHomsIY8ePT/KalDIGTnmXEz0il4TjiRPjq+mIiTOHFthY/JCJtFNWbLzTYRUsauzCdX3iNo
9VP4+LF29rjbpmiCHuFj+DWSictysMXnqOYxHwFa90HISCYab4lKeCnllL54PNryfIT0E1HOZF38
/lOQ1KU11kXMXoh0A4ivDiL4VWzoAYwO2ic5xTWM6d0qhzrsXV02Z3/kBNEaQ/KxHyrttonPR+L4
/mxVGGc7AYA11KvgHutMqWF/S9UmPpB3V9LOX9Ihg/NHjmYHHYNIw/rFwySfFU+Nd+UDkmdll7Kp
NxkeNLMAo8X40sGdG/iC+9I6xoTdu8N02UF4REtmK/ndE08vwswh9gkxtrjLeQRQqoXPAoA/gz2F
bB3r6qk0VXCVjzBAXcAMy+iycmYqRwipxG3EJ+33PY3Zkr8qjfZulVLcdYS1llmExkvhS0dBRi8f
T0SgG3XgtBGXdL/ukuDcK2uSHLyZDdi7nhTcE7E+yWAeL/4knEqio7RHV2L1pD0IfbVRdlQVQfLN
/OTVgX/SKjOn2MIHPOv2Djw6zeXIvGi06LlnO+8zJOWEJU4Gd7Bfao3JrYqSye1hKNAbw2Y11FBZ
/GjLVpsSgUssgyRegJuh9OWrReMJhnp4lWKmCPWDeMEuKUhcfaEsE5oGgRIrWExoPlTK/8MQ3GVu
/WL6VdcFDjvNx2zQUp788cRHEZ4kj/wRk5QaVWSgWSvBSBmLBhhwFf/1pISInNgepgD9L/r/R5Tc
z7wR24BcQBBSp4uhou19wS39m+TcYY+io+M3ZM5zQq0xc7OdSmsagH5EhP5UVQ3Yk7D+AIXwUYa3
3GpTke+ZMfPdKyA7rs5BNzbuWDZlU5/V4VOzR9UJ1dGtpmwOYe5Vqe5Ztvu6cQXqM8LFOKPnoLnW
/jWKWXNv5aEEPa9Mre6f04IJNM5V+4MbJRdSutY9wl0rHzD49AWEhW9B7fAhfCx41C6X6Mau/t5T
eq3fWmIdiPJeU1fAdk5Np8xDHLBjJDbZ1b1Dr3N1uHhYhcEmd0XNCSJP5PCkMKf+u8md52O2r5hk
wagBmTH//orzEjVe+wgDMXsiR7EfvTQFkCGlkHD2wz6N98SPwLBFBAWn7E5HMGAlmvs0UsQRD8AM
O4GX/EZVILpQxMtYzjR5AbfXxCI42KUM8B+GxiJkD0KlYFwXnGe0+Oo+/ZB5nTIOnhq8Qg1pIio9
LxyS1e8qf6coNQOENueo5b6wUsp0fzAm12VHuqVp6VihPiQglqfPzPfY21SrEicdjwB7x6diKdFo
aZRnRFirVmcRtYE3oqAujoC2Pvt07+M+P/1Gl+taDuqiYlHsukQrvMVTQ8ypL/cx0h52Rfaz2r//
bPvNBnM12Pm9UVe/36KXH4lcS9dX0UWWJ6x9iD2lvYStROVy5PNCgfZAi2LE69Oofyt99GbE3cGl
IBiRHOqYxFWi/Nxc5/Yei2xRQdpF/yHFKDj5IDUiFRXm4vGeCAkv69uNq5PV5nrQ1At0WV3gJl/0
zEF5JtBfVYkIS7LXcp+2dFs9gzZU5fvGAWINNfvJUtlIkQyFfwkDlnmvNpMMHqeboxY0GlpZVoXm
8hmvsaY7KCteDpDPQXYuNa4UfEPsLyUtYogpoINaBHI7NLKkunIpDUEKN1reeJeUSqe3qccENAMx
VzE0UzwVCMky74x8v8Zt1M5jlgtrMGlXAzCNzAdrgLO6MU3/1GHHfBs4XCBOZVkL5pn9D1CFhYFg
TDKeOLkmCKq3VJeG00cjhuxAPn0Wk0At335P6wQjKU3BgA5C8Blae79ile9G5VyyjntrJMd+3vjd
QC1pVp8/nnPBWMkybfiIyR9s+yI2S2qKorSzn/TRDWB9/n6vutAZ97ayTONV6nI4KMNPaY2t9OB+
gLHNUuqmBvc0ESY9I1oBO8658OohcRS0b0ndrLPg3I7NGhqw9QS4R4fclM+BfwFbGqz7Cy8MCvza
SphURlvNfXYZaznzVPkJq/A5KKVJbOLpO6OkmCyHoXesKWxUooASYtvEEHMJMwNydkOrls/PGltP
0Widy9VU88AkjFJ6QPqlhNmjMEUSDz22tAJCeBnX0f+xSV0SgUYxZAqzAeTBzXWC57StF1MmlJ7O
ZQZ+XePetuFF5cBHVxurxIlO6vBOUw5sy+H1fajgivolxm1/thvwO+cCgssI82SVbgu3yulkWDxX
CzMeE+HpRL4D5KSZwjY81ao0JLrrjm5PRMw/nwLgdinWz6+cJBJqzFVSl95d8pmytRlBMc7xUPQ3
dfqZLunDPZcCu6B4yJHG16x0spMPoZXto42KeCLou3u+cvqn//QQCHKFBkeJsRcPSyfEBhXFJD9G
/Zhl+D+dFLldOFAnYsyUxE+yJi0Nb7fJ42EWDQ3y83oYbc2PjlhoUbMhy+7LD6NwOtnnBHIG/ZJj
uyyZUU0OPFkqH4EOwGYQ5iBvZuFJHyagzBKe9n+scuTobZcwsXriLBT65MPHzGTibMsV6feJOk5q
gtfWWljmT9jczJawmiJPIqafH6fWZ5eNq9r2rrsJf1rSwZE+Hvc1yC5EdEvtFuPjD+Zv1KoqxE93
WhSRu2fGtDXiGgFl5xxx+xfWVOQlJJEw4/HBrLRBq3cVDP7pQACfv3/pARNX4WQp7hYE148mRkF8
K3vizLua6bE9J6QTrDqLF9llNeGhUXbrdaChv5lHwdon8f/as9EcTXB8yoBc1BnhPVBDWlpmAZe7
N0s4hH5jc6/aJInRmTCwdhJXkWZooz79PiF5ryYLW5hcYl7BzJEXcHg2nnGMcpsyon4F/3zqxWpL
0de4gUWqIFOdv+jvq4flxr8AYoOoAz5zj1C3rBavHntlKk8Is1Zk/dzOk1h3BiDLiQGkQCyRhF6B
dUfJlACdjACaUIYtQt+aXe9ukwk1XvDzLogiwbXqCfgg2ffK2+VsSqf2gLwc30gmabzWRX7OO0dn
Bnjp44hafmz8R1gBUjsO5Um2C38gy9jdphcqQDh7pzWseH+HrOXymxR0Euz/TUmCBUd8cDfVgYik
WJ7/cltVzQOZgTtBmOn2tgtg8xoSGc3TNYqNKK3bWpKwqT3P8Q7hJkhCWtwIX4rT4B9CP0FkOUeT
ajZLAzA0C4p6xTA12VBgk7UxKdszO7FF6dK/fXvqhw5kQbtcCx7m+0LgHfnj/DWYE5XdmKbsdsWd
KEp1Lzr15kLPmnmeDCa9CVjajcAUZtuxtJCwpyHrvo1h7t/Rc9/qpFCDzP8YhVc0SCzYpGOyFqGO
3JUbp/2iM8hsQRuHxvIhe0cK84mFkipgLj8sJdBUwf60p7xQus4pbVlrzP6VHOOZDM6UICxvgflt
fdCdQ5Oh12JEXiJ6jnMASzhJ9rnRKlgAGXQKxJWs4gDfdJOJP2CReImx8ynEmy1r7oqEY6PQ4Hq7
AWzkDpRgBWAXrJxukHlQB++eIkm6riyfqS7IPZ7XLfq4f0rpGLaWgaSi5onU+fbMROYe4vDGom49
kmB9sTqGbeRhYIZmWSmZflxC2m5dcxA4EfbN+ECbO/PB/YpcoF5ilbtvisu2sKW5DbP2S8yNFnBJ
jnbMfe6IAJwn2ICGNiNsJ76VkIELRqSwKGDQJNEl+xdjaJfvLFIeN7QtX6WJ4ShSoXKuqxT647vZ
P8pMB/wRonj1GAZ2Gh1FkH+L8qGG4uDVcfY0u/OP+eROvaM+Gc1mZTxrPCZQkmZPhw+hoFeBeK0W
cdIx/otMPS2flSVMApJ1V0sNgV+WjXCzvPiaDfhYJHcj7ZF9v2teXwNMVvzQAnlXPe4ajDP/LqeE
2m/QK7EUwHf3E4pqooPxX9wiVOUH+haQdReANxaeTxL4b9FpMl/IqGd4a0ubc1wjq0KJLw9MPn7R
QJP0M4hqx6AwCCdpjLwPvQ5aSeMY+4jiq6JNiZLIZrVmqTjDYvK10KLTLzNOHQ2Y0jPmBSfDkdH5
eassyIH+JOveyXy9L6zRxSQ96LkWEuPyIhyAjLqfrWZwS4prihQ56FGZpIOSEPkUQ1SJZRWgOQGP
G6xoHV4T6i1zW838k0kwRxhb90YJfsL9LloSM3a+vDITUVHiIl8lOg4S99oc4yxsiCRjMDeA61z9
BlJcCH9nsHmgSdbGrjTboEzbjoa2o+pd7VEpmsnMIrNbZyWXhZifLyPCtQYjOvvaOiI/cxEiYXDS
5UlJxZPhqxBv6a4GNw06tx/RC4RwRH8eyk68qLgNHchAVIOWovQazDXFTeE6PR4Mk9MPSPKsSE34
KoGUhR6xwmJLDnTHrZ4FhRvAlygGUacPeEJCYAmiFtcUx6FaSOb9Uyskn3yzpq8T3zr4EjS2Z2lH
vDzZEcLUfZBcUfXcvhXYHsC0JC2VafWA+B8TKD2mwZZsLVBp/Pwh9dX1QY//ixgGthjA4rbar1Kk
Qwsssi0OnqlKhN84igmo+cMqoqfP6O3gvDTinoOmNyr7WafOapKbs9DcTdZ0IfelMBPx97g/zOgM
INE0Yb+JAQPAaA3X4WWN1i2I0fPSMudhvTUD3aoZE4Q2bnv32PMr/VTUO2HObqVKdWTglJ/ZxDmi
QIutlCzAKJB15JiHUWuOC+9s/wwuXYrrsNoc+EhxKLtXkhyie+vwii8GpQre9p8an2yeXnG6w+MR
qqjLDrEsNHk9/2zS5lqVNyBYqVaSWEuA/K56oqXKWIAj4F3Zeh+JuSB+KTPrLesToEAvChFLsHdU
X0puyWzBf2aVI6J9hszSVQO56ifa6b33bqmvimbiQ3z9qhV/3/PE1xCd6x2KJTEv+/pWjalc6hLJ
v9ZX2Hni6Kbh/P6p3YTGQobv49nmpOZRPxeczavO2RlF4GSY2a/mhFK66FPyAll8NpyI4K2knM0B
CtH4NteDw3UK4DF0x7WLGoyiFr80eRtWMFL2skXqsTSVKkZ0jA1T0XjyMLszJKwR3LyhddvTsCcu
+qa6aZeZSbf1q+1sXajeSUPsen+9FjsN+snMk7QCX11LSi8nD0LfaWsSOGYCde8KKhkmrO01LOSh
1fTg9tNLF2y2v3X+GcH6AvVCX+FXZw9pm8BhLjZVVLLckM30VTtKf9mHyPl7taz8thf0EvhsG/Nz
Z3CuCitM+JsmM0FrxV0BZ12gbux79JMlm7RPv3ugJPS/deO/DliRzYeS0c/jlnv2BmOpNAkdbfXs
tMmRCT1uS8/MrhXEglqu3nvvLt6J7jHX/YBSV2H37/7Tcpwf1CVw+Qu/1zhqoAwDC39rLevNm7Pu
1A0QTWR5co68nsqZDoKWGe39ttBPIX+kmF0ZqRpOqSor5kSZDzObqAC9QGPDC9NWvNfQKsUT+yxI
p34m3KTvOUsxBSWHBZZzgY5kmj/shcsuOlSM24B28Hq+fqbGiujj9a3w9xcp26D3Jp5GSQnm6Tzu
GXJxUbOaBpz4OoOkRqKaHkzBsOfr5/uVuhYDgrygvqDbqL2G4+SKx1IG+bPAyo9eqFs3D/QLEAU4
FovnSUmm5M01q+exxFD5bOLtLoCELvnIUkwKU506zf7m2Cr6lvi/VfYASYsNK3CXa6rssyv+iKJn
c/crwFN7Cl/U13gvAxEYE8KjbQk+1xtbSha9J426c6MrqaWxnWghZG//Q1VF0UvDJ++Yi7LNmfRm
KXVYvsQ3hCqj9iH/G8f84bF9o2xDZWmLB8r61vm4TJ7/oZRf+UhKBSKYAN+XP7M7qbl2+kxxONut
s2jxNMXiWyCYTadC6xgyictuOMFLGuI7osXmQprSJMYVd5E8b4IyTQhs0Q6ioLQklVDareM9gf7E
tNDPRFoFB0DGrltQwEs0BtgYSvz02AE8Jbf78l334mZFrdDKgRDP4UotbFB4E5/dyzJk2Z0EwQe/
NNqcQgPoX2jU0+nCrP1y2RPpstYLAgtE/AkSAn/YBJNDERSsIod0VptdCEprM1Sz2mzvpLrwfWK0
hLz+dVvvvmPNWCq8LMtQL62n0weWuZc7QUPHx5daaPDjmN3fq/Fo8kdLGRDnzfH+tVdmOr1heVkf
iysRcawGYIr35CLQfmr9gr3TCzmFpi3900Op4jE1XFkCIi6+JEPeyGOol4Vn5aRDifAwKLciJjCj
aVSUSzRjUJFnX6cpNm78ardI8Sr5r0rfGPC4/1HSa83rhZ8Uv081bJ0dyntZzQUm9PxHmdcXxOqJ
3MoD1WywCH0Wp7hs+pgfrUZPjwNXV5cEiGp5Zv80d7N3c7ojOrsrITrFuhti+XWRpTGVq44ucSuF
5CuUyS9QbKku+sQdqUKMVGuL8Y01+NkoPZGeUqcq4BX/tuZ9MeEih4Z9+1J4UPzLNz45yOd8VOJw
zvIW/htYDhWGAufL5p/Ac0MRHxmZjaSVGVcypNva+IwZbm/vUejwQo86UTjxpOzN2JG3LJFkBjtH
lFkE+N8ZtcpQlf8wGYQF6t+UO4PORjeNj62k2uwT40NXUSwfqTb/Wrsvrl6lY9b26ni+WSSdtdKy
8eTBPrVnxlp8fWWRjXHBwPCQI09U8k1/VHuixsqA5osd2FhkKL3bcX63vWBhhNU8NOc+ggqPMFLL
4Y9tzbw5JW2L0N8oBchNy+y0NCigPaBRuaIAOIawYQeFLj/jrJGwyVTHS6Y3aiZpPMMdpofMIHEx
lb7ZMSBJlUhHXmfaF4g/JLfWYDV2ll4mdcnx7UgXcsmd1dQRUTG+tH4omzE42KM9bvHoc5IhemOL
YOwhP3410/gfBCwTdxixOZ4IC5GW3Brs8X0JQop3xCZs2hir0aj5HehUpOZIobqsJdSDvGaeWp2T
T5tIaeh99LYY8PyNo12q3M9iFu9WOF+hEBRPsgthnXPUN6zamVw0V4fvb/eCW861knP9nWaPGy1t
EB7aaBZTV7zzmFYIxo+HK4z9D6nIEGSkdndF+4dhbnxt6ptQFCp62scS0ThcGomoOB6K8Zg54mZz
2VRymgLMLhSvHJHHlM7J00NKjrJ0rmwwFyFoJ9kkQgmkGiJaTL+sExKWMIo1mD6ZVNChDJlWiwYo
lLy3F4srjFoXo+K2vLIvrwdmxFmA3LgT3V3gge2OVAfR5kA7SgPz/LULlxG+mATD8p5DBq9Wfrwa
Dj1+hvwSBvHT7qHf78ixe9Z5dW2M5S04vuQFw1qOMRExQgQ6rR3QeXxpSgomu46DmE+f3F6vg56V
ejGmM1TrtLTi0JtuH2Gd6xHWnZSrtKAHAItSESiERwMcwEEoKUlDTAgi9lgJ9w4gan8NkVTcDyUs
/O2UTxB9L1T2eR3WFBBWMsHQeHkVJN+dyqd67kRHIvlJYN+ELMHbzG+4Ek2CX2nbADi14/pExXzc
CpNtkZ8ccmNGpG4r8LQJTeO6NCthy9jOIuRBbiOl4X434rO02CLxfltsFfYpqUJ8jLwrAIy9fu/U
1xvpt78RZEUJtuDvB9BYoCKAvZazYRpQ60bLIAHLFOeur7WRlHsD2mLcOMVLo02Dsn21P/TQE+Cs
itfph3wS4plbyG7aR6Un9h8cGOxUgTCs9FR7X/7AKzISgpbV2aTFkI08M+yhHyR0sszD1MEDzNS+
0+GYk7McrMrp02t0C0jIjHylrqch56+TTC5jhC1n2LZGtkBL9cpNYDIk0qyNImrokNnS2JLfO+Hx
C3/004mMuw8eFClCmvKEWgx3PdZ0peREGJ/xYkVmH/9rKfSjdtecoTSlnYSWdbKJTpcOleuHLEsb
1FZ6BLRplradz7tHV656AmhcdYpxjlvMfCQHnJVaonJV0UkzudVpii9G/eAxBdYmp8dgxDPaO5i6
A92sp7NKUWsW9+HZYmY3Iq+VswdriXjNMvcjz8ScbBYwrXEQ/JKNmrvFQcliZrEx2f5WxptxLj0g
vyLTIFNgW5xz09MBEfkFyEmJz8yvk+nhjq+Jw0f+mEsZhbpO43TPFKaOI8AFjIHo1R5z4n30abPt
j7R5EsPxG2jAdzSJFEjqA9/fMkU5t46w6o8RQ46AoCLSuDZEMR940m+xV8whG7L+NFeYA7497gap
RjFxw1BqYeWFQaKUw2O4Id/vKHeNlK9oPykMjJ2YdQciKZbes2ESLenAiMs9Ia4we9B1Kg5NTvPz
Her4C3yULDl0FfsWFi7DKCJ5XlAAwvqCCN4gFz8SsGWeVxGStiHnT5bO68fEqXZx9IDyt5jPfSUy
LhoOeHE+zlwGfIDQZBf58mkBOEKDr8KtR7N2Tx/bYUMKdfdisT42tn50lMSACpxeDQJRBWtO0jr6
pKtmMGRNDlX1E3LV1qrJqCfeIBeIe+nNqtI3q6t0CsB/xcGu81ikMY6kZvxFUSC9T8OEMWrcphTC
nx/fyMKFbC4d7nN8wWNt83H6BFGNnz0wkyUvfr23HZJoHaIviaOIpaMjGfXNeeR9zQj6qK6cI7Mc
UcjhDjaOT16DpjZS+THqIjbBrWiZXBE/kaUDz5kicY7pNECsBky9zPDv6KxZnTi/v3HPLya/dxRM
VgUNdj2L0h0/sP/lsNxz3ed3Fjhx9DiGa7Qy/eALFIJysnso4idOCeJ/fZDcbXS5rWGINCnEVYc8
QM0gQJcvlPABSWzN/E7pv5gVEMZwEH4IxxSpGKJGlGVqCtjDyDp+g8VJJnHoG6f295qnBPI5IBSP
wSExzfjh90Aq9JFv6VgUnv16+lkIeZ3X96CPN5I4QWLauRF3UlA4vU7wDpZOLsqDPauGE0QJs6Ao
sxvrIk9JCR4+Q/msTbVLvrGJbfW0x0LqfEbf/Wi7BNMuOlY83VUgYMvPwifn+wuUO2mnrp2I/kEw
gCTRVBSvodVGxHtXJqtaDufhU5och7sFPncloQrFcjHgyxVnHg26+4gL9Uio/bxfKjgWga+ow2Ny
i0gG9kQogfhhA94CrxmBEvQL+bbJrjhCHg77Y69XW7ATS8dKA+8FSbimRXvtFw8JaHoEnN+N5Vud
OkWMQGIBYIY73V/9s+FsR6WhBj2ouWXOdYpth/5ANgkHjtw8SjCSc/IwyFiFYu32UYTegHr+I+EC
G0Bun887BrbEtxSCaIRlfsHFUPYcBYweRDQeaIFlQUiUX+pD19PEa2FV/6rA+GJJ/JHfWF/m7zBI
qAWPhjOoth7m+zdCjYs0LqAN0j4Xp7908SPl59oSMiDIaqINmbW2+hWoHefsoLH6LEsfrzicDZXv
xmZqHGCyYfpbc2dW9et4cK6fEm2uhIUWatXHfHN4k1rx/ZFL2SJOJzG0/vCF0sFsKPpNJkwkgico
naFDGCekmJ0up2e6Fl58Jp7JjKXuf79F6+FNC+wS119pCP5nDYQuFysN2inzQzm+NbhnWw0pLauL
BAFfsCDn2nuDS46NaBNQNvp1d6volEU/SCeMgoDfpDwPynMRpWi06YwDpHna0zhDLtru+1Ej/h67
YsaG7iaebi702m9wsqvimcAytVY4/H4Symj4CaET7NqmzwsukRyu/8Cc6VhOixuN8Tw34Q+eqzB4
30L2K4lPtRRfpoT4O7Vd4hiVRFHqpiIE3iATEqf5b0EEIsZ4svmKN9beDPYWJTFSRGbYy5F7v245
8SI+bCXTMARveMVhAEeV+cmU2xxM/q2lioCl/JS2OmQEwYWWO36n6tfbLLTIpYMJO3hMjUtKtEDj
3PrXGwSECqZ+8fFSK8uhyXKE2a4BaSX2qnd+tFGqWttEjPQnX97C7utE1ChjJojkCEQDc1TjG64T
qQRdwd8ngnRAd1UMsDG20Mb9RaAlU/VWwbBj/SgjEhv4+YAYD64uFlGT1KUIufaltDzdH8JssK/b
fvLmv8EFgeTYAb5hzDKELf5HRi44sND/uMhv4CEEIXMPvGxnJsBSnGf4iGzQj1rEddv7SVqm2eb0
uupLrvDp14O/YOr8v6DVOs703PTKyzDT3JetWAeEDKBFGUOeruXR8WpXWitL+6zSNpNTrq01oglC
d9WOLJKroYNabFJXurM/IucOFCIeoDJOZrUOf1FDQ4/1MZp0MBWyVT6DnezJP3Jsa5RGuOigCcLT
Fcrq0Xz6XkHUDBdTAZKCs3xwrcOldhQjEAe+M3d4i/ZT9TKMbTBH+GFbqE2BleudvszctXLjiCr5
of4nU5Tj/EG1Mmi6x2QTWWiEjNwb9UoNiKnHBa1JJHjZggK6GUv0Ojpn7dq1jHQPItFLm9lJmPW5
ojEhEzL4qFZ8RXIxOembop7cEvKq1ZMTEorKECtjjHzTr2yyOPrO6bCdHHGi1Wa9xiG4ni3v14sg
jPvuNpThje+LmDn3pk/ruRR2xExLV6pNm/mOvsmfI8vSCRhCWjMxqrXj8/hwfJPhmBJ4gLarHV3L
lnXKHQoE41LROKvFEbvZcHgTqfXygqcOoq+5rEcpdmPt1uSHfMDXR+QYkIwG8rgsWmcTQ8O4Bbx2
0m0xOEPKVJi/+7B2Lnrark18j3TgP7V5yjWFmj5TNshcnxnDQU+qY7f7DTONb2jLcyqzyK7Dek3d
TdUzl3VQwPXs1lBM9gWVYL1B7kZhttQG6vvVc29us22JbYgkFGrT/bOsEMNnHA1ZfJkqqWL5cORG
AeOHfg+zJ9AdibVuMcOG1QKlSsG2MviXl1dXkk0AzcOLXaJNiYv3E3xOFhiChwJwNDxZXrMA1MAb
5Ck6KC2hWq5zbd0t3mxQV+c9U3jXbQERPVZP+RPHeQ/RnzL2WNU8mshWLkVUGFBS5/RQ4Yb/g+68
WCb7rcHkHLH3IsxXNCe+R4i+YqHSdg3+Q5i0Rm/arKpmEVv58J/jD7CLXyKNtqvVIoiI+TSy/JLc
uVYO72KLUT+EXk3WWsm4pLiilHFxqDelTgo2JKWNKmUCtEpJpBaW21Asxx+sSgzAITgM9XhstCOu
ngWbASawZbn4j35FCx78Pu2W429ZjLAac0H7aBavD+XoBrCgO2+5gSW9CMoED5/Xz/74vP3dMkvL
0YnwC4E6Nk0Q1kNKukvYzEKSuGoC8PEAJB8oTWBjqXKvwgTsoPlM5zAmMlEhlzhndfpCTVxn7Cud
DMnfQLMnyIZY6WLxhE8RNj7j8gLHOcqXe/vMkSFH+CzaYNYE59uXdZzmHFEuqW7AOgiWSSy/jEhZ
eDnmhTKMSyoftyjDnVnR6YkYMJ1qow1M5G1ASQ/uth+XGKZ4Ict2f66v48a/pydBT5TraoIAZzBK
uB4/lEYk3b9EgLqvTldqR9O6B50R8qeuekArzvkfam+V1XgJvzQyH2QNK+N8vlbgs+QFvt+IR2pY
tC0FCgCUFXZqfYyNwG5E4LIhDK1kx3rM+itqKqzJjL3mLjK3c4jIXmDHTtuva0n9Byyw+IQ/gISc
CnlWl+lRZHEl+3JPDDorEs4H7AHFO7bqPgTAogF3kpZu5cGFcbVeJVYGdXMRftaS+CQxZPisebUR
R6ZyIQjzAPiVgfkF4PR1ziU2ippY8NFMmFZsvx+Ym7DG4gGXdOfVFeszDqXMcBx8l6yS2sN4vesh
qsNwHbT86hgO4Gf4MJgAQwaZHTp4ahdbmDZ4jW8mcSgXML0chjsmBCNqBArjMwmnt9Xn1047/ofH
donRjWoVo2o70W688oVECT7D2QENzryKafJWvf18N6v2oc6+jQN/SFdpQNFt8LwBeBoV470hKBGF
WpCtskey+hxz0KOPti0IFg+uvi6n+S5y0qlh1RkkWsm5OZPZ9bEO/OSZoe+TV4x68xtZWbJjbuI/
b11WrC0MZB0LzgddDjEplAecAKmQ+ixvERQzhLrM1HL8vvszYXBhaQOC0IvIbijf60xhQ4a3Z280
PuCQV35rG/Hv5shbtOpV+7GU4f8+zOtACC5zqtKUh6jdc5UR685Jx+oHArOPZ3Jo4lOof/XCS2lp
1cfqQZh6/lgBMUtezh0o6QkktALesZxaxgVH96aNakWiqLISlxYtMfOWDIjqVYhzLF9U3af1b7Mx
rs68v4qp8LzNH6HlCJSdDdgOskVwFQ+fkPVc5Qf+AOKUtYIXDacqBZbzRCM9/wr+zkh9lWLtnjgD
5yUpkGCRMOoQ63t03+OjtBAUySfo7nd2lukE8bKXHfOM0MHg55Arg8kv2bFoNgcK+UYEssY/800a
wkkIBPMK1ovHJv9eYLY8DD5CxhesyF46GbRKyqAxnXtw4o+U4h+Y3J7Upp6KMDA1Z6J6wFg5h4kc
5i4tbmjdiKdNpnd00HZN3QGE9B5+rg+Xe0/uKyiVtqtNqWlWtFM5h3ncd3ipaa8Xo8GZ9hX9nsQC
cypXf0AS7l+Ygr0UFzGnXStNLCsBaVshcmZ4cqr52TQp2zBla7a+fW3x3ERh1PnX3sm4EHnYJT6N
c0x+PRamSVV4xPPzb2ZWXRIfst5lnMKIV3dK0QNxzq/NZSwVxB3K/Bvp/8cU+LjGCT7NXH9Trqjx
Nh122R0tllECQcjcCfNC1aBhfKAuyGLFmE6dziL4i6y4CM0g+mnSWIMpTeVP7uddsEIuPoSyA7rJ
DYWE8myfPk5X/IPyaAjQFDNCd1/47vR3pLzPo07Swi1EfRKCG9gLQOAe1xt3tdKdspQWJBjdqMQq
cl9oLbIgd9LMkLG0DeE+nmWoMFKg6/nayWfJRiKX5nJ0RxHxMAWqZxgqcXK6AzI3s+Qxi8KiX6SP
NtgwC6KyLPB99uGLMabOyPbx7+tpelquUcXWjcB64GzTqK6cvx/lEp1+mw1OkoWyIAYlGN9aDayI
GNTyGq/jG8GCcoZcYlRZiiqr4LS4FdZmvO9vmyFOIdBsBikU37YWZJfGLcSZeRauhWhOJ16ft+A3
7bcVNDwDGrGgYK0d7YCayQOt1Av8YU/wCBrmnpFfd0UtNW7SFyCY4YJvr6W3d+ENrJoNvgLIXYvK
pPkE1bcd04Wy0KtseD4t9hE6Gq6kCVw2FlavbbDjqy0O2sW0C5LyB/8TnuNlmK+uUYnCkfGBcyX+
zLYDgPM51MeBojbJJt4745qBMc/TLt2j+5S8wWoWKfqDUmDL7fw/ZgBc+aHCa+g4c3DWS/YLidbf
SY4LoOuXQEOzji9ZpqiKjvnDLEZOMRPv21V18Y3zmgtqreOfOiYEbBkbIeBqm/m8TV16Vsv0g8jG
jJqERuEwdPwEanHjDOW+ZauMw6rG8Mu5XQvpwrUo+G8IyU2cWX/PDTprYrnEU9vux3n9jU6mdNCK
dzMCIsLU2ZG3JiI3n8VmpziwF3kDfwAisnNfq4pKY9fVyjhNBy/Ki1cZQybaM2EWCVFRILBUaVy5
EiN6ksFIV3ifnR2MT6CWcI6FB52NseMO7paDf7Gb4ywVl39uXB0C1Q1Dsmv3toyI9wnRFd7eXV2F
b90dTaYpPyNnOyqvG09kkRQ/Fzhx+C5YCud9pjo617TGdkUnV7pArNUUZ2QeZERFIHTBWnd7JUhv
crViwGpFsYWQYQ+ngDnY4aAPHaYN30R0TuMqjetcRMYgCmMW34tIQ/TlEqPtOBIvQwN/Y5gLJ2VV
Rct0DjFoP1TQtjryPUyVKMhR4NsphQO8KMQdPMl6Rp63DBoVerLBMAoiTH1UiV+PBjC2BWuOhSIZ
XTfObJSiZhQHX00tuEBdZ0kBsaCY8f+qSqv6zbBZbuwlB4o5Ot8g3X7cVsxB2l6lkLcFR+ZEccoe
bhdSJFIU5yGsmOpqiRvh0IZXPZ3UZQl1U5qOTDo+f72MqhMAK8MLLWNTandT82se3cIo2iUUx5SM
//7ac+JIx85gY6cm50M1grpTDXuXuGuNw26T+QWoHeVQj7dfiCi6/gYo7uW0JDhZb6t73voLVvmG
JEQppwUy5mA2goTB+NqSWqz7bkTuAM6uGxc8uTitnALnX9uwaK8MZKhHLbhXSQ7UY1AkxvNcKzSB
Xb7J9sQS2nRj7jS6xOu8oGykBW/7Ga3PMxiAQO+uWdfxdBQsNfdEXV6whH51RlekRJ5eClIMbLXP
AA2DyEYdumEoS1goiWIyr6SVZFeXhliQCWLGauRMuYqBOQsNGdKYAqNSuD+7LQ3WphmqTTSTDJQW
gN0WOEYCLITyVl2dhig0m46fzDdOvFd7gMkYbPyuKDFdDeJj8b1uGMl02nY+NchsQO6q1Rsq/zdX
6PiZHkqieRyxkJjvRwda6V4A3rqAdUGCNtI154A8zt+FJlK2zAl8AcxJG1a/f8oUPUgScWFGGbTM
xgNaW+6EHvQ2BJpsO5VwnLFEI8ZjHJm2vG3F0Xov+Ry7UZE9y4K+44JopW1I8at/ZdZsOt5IfdpB
arQj+Cg3IQ9+m1eWwc54HQTKqtQoqR9JxTd4w7jSKuRbmX40JNNaOfAXnLa/uEh3U6XdrjWv7ffy
szr+t6CRmFkla1El0LmMXMwV/uhi044IUpjko/Rs6WG+olPoQ270H1ceML1RA2qFDaaeE7rY08nv
0SeibEZ/GLMQqCwcnoB7tJ01DFISLQmfLqUMlx90ZjKHYo9uJUX7eBV4mL0QqQbnwwGitkFBdcEm
CuWbOroSpAyT+ID2jrPg2Bg0XJnCvejtgjycPzJQTNa7hMIGBq3wYYd7IvNyxImFrF0ew4MPMKC7
TxXZgAFk2Hy5h2MUeNZksomK8Nc8BTZ/g7+qfEpKgFS02HybgiE3Wdj2bOnbhlG22xdVtbyCKcwz
Tr+VF5JVt9R3GzRpr53q4GlyME7YtLtUeA8NpEuM/AMuOrfDsYgLVu34lRfpqxF7V4oV1b2F/9yQ
kSubuhkiFCoJD0uq3wwThNnQzv7cTOFoyNT67Or1ksmTeMfk3UyuGeh3onN1i93q2Z2O9+V3yUl4
RRZCz5LhYVwNfHED0Gbx6p9puxuOmC7ZMvO0xLPWahuVDzP2XbDWHzM/kt9ahTtJp3McAupT2S0I
lzx0PXss6ZPWkn8JIBemvDnNntiYabvm6a95ooZOhbFE2svTIXEHpTt5LtC3qf7rqk5e2WZQxbce
ofCvS10sFZxAOnsvSA0CDQLF4LhySM1H+Ik+V7CU/XD+MkIOhRDCUIaatvzlRuM1VyzNaUbFjU2o
TtJEMIrlVJe3TTxFXF/iVTKAsKxA1I8v2fuowf6Q3NjSnaJ+C6hbsQUXzHYhSUqTqdV9a8wgXDFm
dkBI36n6zjAy0dVA7gFqL/pT6yC+6E5cYX+RXB2XGuzUdozvFVqPc3N0gic5L1sS8VDGHW4NgYrO
WS9QpV+fPhOFRPO2bkb4XjG58UCLQjZyQOwnDJ4CcI27X/SkGPsNiWsvAQfqRllSi2Qa8FA9PEm+
vG0a5kiwqVqQLvPtKcBMv+pAor2Yf+aoYcVVxyzhbhhqlucjg0TDAOYZgOmBwSRD8FihwFqez8T/
SUnMEN7VtjEqqSc6DEwIFGD55WAkfbL0vepVJstZVjG6I8eBM8SnvkGUWbD7avcQagWc+KjxLq3h
G7sM9ZJbmNiDDUkK6Z4KQCH1JLU9LjZixlhTUPg5TnxvZtHWKbkMokBz8hX9WkfjqvdxlWRyURbF
PX16dRYZm9S6W8BrV5I3r+0uv84Vuae+Zd24Tf0FIv04MZobsIAHn2vggiRPrWQhkv61sIFfwxXW
tfOAbngyPb/QgiNjkNaOMZGjc+/ZZMbmbuAkPrlmHr3vF1r3PffdCnXaqmxlWIfIAdAm7FLNtUEa
VnWZ9PdS1iEBkrZfKfN5iH5mi+1mtjAKSYGgvCsUV2iC0W+dCqCpUcLrpMm0vBIsMsV0N6kGZP8Z
XwS9A4XaMJJwVPV9VRAQkK7Zc+kNbGSyqDMPDtGpyvPjBHpkZJ+Y8NhUCJwwCH6fXRNRp3qncAYk
85Y6sfwu6FhXWr1wimb3p4tHOkEJLPWC7uydL+opjr+h3yclbCAeKOxgaUNPqgwTQjNXoI4m6W3l
jQl5uV/SjGDGM288pPSx1mWSwHiuomfFnR3pdXfz+a4Tyv4QnhGelXvwVRehqctLKq13snhiAtC6
sSf+UinuyrwYy2WPuJ5ae6vlT9nIJUPYhZvhMNoIi9uCP2GqkuGy0xDBgHBi1DYgM6e0Ojev3uKE
/Cce8V+VCMrLH0kKYi5bIwH02thclsU0pbsHFeAmT9cwhGnkbzwDU6/YUO/YtP8lqRk9Tk+rzEvb
ZYyrvFnkn+trW3CyX+sqVYwcMoE+k29JJXVG58iso1qloU56J7B486gsLwr2UKyA0uFfXpHFnqNX
hlzitb+xXmci/QPoo2rxY7SUK2vud7gFCqn51UmLCZcOf6UInaGQ0ixcWmzr2Lz8zEkYbLy2cODp
Mwo1uE4u3sQ0hf/WBLFHMeWFZKYcqKw/UStZyu25isTOQiZboC/fH9Tad7Of1Yg7XkkDFBQJXuvT
E4Bbvb/Aj2vS4k1sxIrsvRwgGoBk3HgN18ETfE6jwwIU+vSgL+P9j/1epv1z/YzsQCnceXXni4RV
ePOJUUgMTGVCyYMM7H+QG6C4p2EAATjNE6PMgF4SpgjO7WFGjAweAEif4rOmSVJ3QJc66bTE730y
kLuRGVwsHHXDxXWR3KK5QBUeqSKdnEAS8aZsN2q1OdjBSvCKEF0w7ovWu/U1qymEMQTvHNXaEjMO
P2kxuJU9Zoqpm4F/N4N5U3PAoW5x0cAC+tHxr/eBAhazCDFZpMvJ2AWvof5dHcujtycLJGAjXgqb
RJsJWK8oM5mQ5DH/pMy83ZzOOCBaS/UInTQikhJDRtIM17j/gLeNvcDcUTtBuikWRRTseWVffs5Z
TBGhLzfN84BSZ8BRm3d/uRi5Mzgz8928QRNQvUKx7BaDjPEjwEaGPvmmpdmEu7hU+NtS3+yUnuFP
GToKlETYJ98cyU6wOyRNs4y6oVvMEyq8skDvhYNwDPHyykIzzapaxYBYAJ+bMyoH0F6v2BDmkGly
9I2F6+NoBhi3Zj2Q8fpJZV4FAiFV1fI1XtBvHGMknMR7JvRdbwOMGmQl3IFwf/Nmwo4RuwUY+OSI
YQRV6sNSVNp+XLVXcSR3mfkmRon/m6tO/uhgKYsRcLCyqgcJF2287GTTh4mgFXvesaK6/Y3luNOY
v7nANTLQjbL6+d/d7CQkTT6f3SSIUMqRZyYzH+siR7x5VLgDd7od5uzpnjhoCkgOzaIVjv+57VEe
N4v5Ba5YM6cGwpOIeQeqGuFT1ZgTZLtvDBb3wT89E4FuhWporw6PYWSOS3/7vids1uZIZSV+bng+
cnj5PB2dEnJVzZw0gp63MkajLxHpyorkmg5EyI4L0IYZtbwuaFROO7Ar3PO8uh50i5WLrjyo85Cc
sccPSzAyxM2c8Uu14IFG4dwCqdKN9YVPZpH9RUzD+eOtQOBYImLuuLuMgbupkVlV3By+qJzRFtTV
zdHBGVbs24z3nAsg56SdFystZcvofEar7q0nx2rDt79sdGan/iKUCjWvx3E1jxtwaNSmmDVCDkBI
t2KMNMheIiV0gCfNVmr51rM3qKu4k6L6WMT4aa2MwEsdbI/ZeHuj7tyuboMuPNbf0Fnv/+XTTFRu
7G9hJBLp2QGtVi9V6zib2CHDfXO7dnR2cAUbgCH1e7loPHdxdVzB8Nzms5uBYMVOF/O/5tV04LsW
+/I20Oc2jzJtOhR9Wct0iF9UtkrdK/BQTXh2qnFq1ORSbf/YvOwIQ39Re+3AN8daRUtRMUWfRb5M
/fPwluAYtENtsQn46lajLfPKn8DVzYghxstXC+6b85grCiXxPCLisdaZ6IbkdAcFyql0Ioqow/dC
vIB9laOZ2PIUj7K+g3zzQXftC/tP5nl2PnuM9bGfF91zKC5+z7KuykxgFXPp8CXfHgku7QwE2fhf
HyPHB1p2hN81FStRbPNxVxKUnJ9EOf3Kh2EB1GtTwJCc8Vq7kqUn8vNBsjyMzuV24tXAL0P/kMDx
NJQsJdfn0tiTf5U4UpJmir6iMgMyEuiVoJWAibMwgqz+UvFWSIMAkan+4VBPR4HU3cPxvs17PoYc
+hzOZeJP1zDVKcCgkmD5ihv24KLIeeEhN0Smvgsf10I4slsWG/NGbPVbo/n4DSTBscJj8YQplXMQ
R7QG42j7121C3m5ii8mlVTFQT5796ZeZAVbVG4i9idGg/5TtU/kaNwN6QdtXWDE7cfDKwIEiQaEg
UxF+JUPnkyPjFveuAqUexSSrkpX2Ct4JgDFkwC7HC06zB+wH0Ld+gGNt8hmwCpzYLj88LphzOPg3
Vpn7nh7hXru/7FFzY1kSXtkBKNII6du15P9YuXSa+7pwmMRvWJmR0HV2kEkX+olBqigVkHkYWZFQ
FceP+JhcWXx7EZi68JNpV9cX9PbcsUTsFRVAZeXg3WLCroUGpnRsHKIevPSR/nxXWpYx1U6CTaeO
0adVTD5N+T8NQsqWpnlfkT10WoZjCFsqLvE3/XQCmy2cGeCHwVCHgwp3M2edjFaAhRnrQnhcSC0M
JjpJH29Jp0lQVpw/IZtWMvMVXYezyxORaeqFNOP6rsIuJ4TlkJ+bTZwYeE5o+AU6mTAn0CPUyzVP
4pLWtBTEg7FfkH/V5wlhE0anJSAAaVFEdr0Kjv04Z1+78/TLe192DQv/OgpCTpjhhyi2vp+UjKSb
4Vb/ZIOhQdLHRp8VQ45FVEV2tjTL6z3BZyD5g+irGE4sEnCG5tx/M5AklfE6cwWeSWgFKpjlIx9f
T8SXu40sMYtgKH7ZKloSV7pLbpZxNVPLxw+CjEZmQl+b9JNTvGlIz/0seK7TbhhT0960oyxORIvk
eu+RDpQ7nrfXmEYj24T5BgyYKjlV6fkt1AmdEkFJNkVrFRMku6ubCGNhqpoLbzBsuNLxOiv/xD1/
f3BmRTkik5MMmL2j1hs4F+lCYq1VZZ1YP7e+6j9/48okqRSxIGSiE+ptucTNVirrY/aW9uwiib/+
pVSDMBWEnRk9z/rYgFOzIUImhmBwiY12KKM9sCmhRwPA/eoZALWqbbQK1dTdDntS+14lAubkAy4I
vG7zpDTKgj/y28OV4L0rZu16TK2MMqdVmfSPV9sC7CCurLdL1Lpc2ZYGjSVLOuOrNxyIcM1hMgMv
KUPvdLoBBEuGvkwdY19opTZ3X5hODXCpCPqDvdG/jnZbFiI6bTit2gxFAkHoZd7/Un8p0WhRTUCj
wAeSnfERyo3HlDxrcCTNZH2aA7kGSEzGUazwPPLOJRKmdHYyXG87RHbI1GUY7u7ckX9qGSpHQRsr
GRGPsOHJwvVEpP1h+MdxlG4u6eKBMtRWs5aTkjBpqpCQO9g4EW2Ogy7hY62IPjSLgZFThE+IDj3j
6jTU29cU4u2uMf3OGdR2jhqMM64SNWlRICC/e/JSDMMddPFDuUGCmXq2himej820sbK+2WXCYvqD
PYRAgNL8RDjjwKbKZHVPaKfBIE/X2f8jxxXju21joDX6/VCoU6H2DarrkHd5EAQZwv4HHWWnp4f3
e/tx7y11Fw9fxt7uKZnS8Afw75z6rXbeqPqScPh20folwuwZp/6lD2Hj4Z6QzCsr9uhVF3jlCLGI
mULDte8wJUAQb80J+8CrzR3bTOr4D+zG/obLjtusrN/dzfR4wEKIUqIPptHCZSQTigc/CPYTVUt7
iUDDjMarMtyD/XjKmBlUumRxErId+++mkHsoadhXepNlN33mgxUrPZWiKbDmLrEDqFopOU83X78U
31hjgdVW7guU3c/xDrvGtVpnmOJhFzZ0JsFhkguwQ/JEAT5qO76WBVFdqaP5fWPJ6uhQDT3CeoK/
78fhLXOiZlATMnqoSy2YVKc6IVnT0RrGl78fFVkB5/lQECEwzsCLjkDHiPzr6FBXaQKnkxo+YUPl
1X5iP6jBeF4+/GlITkmb/K4/AYGzce7hggl6uBr1PTIFI9gcPNdiMudn2IigZm+vJjA/aoM9gS5F
uZgFAY1fDsmtp5i/HFvg8BVH0CgCTDEkuJajk07i24mHXgUFToZgz1AOXPIDxZYmErPdLpoc7Ofi
dbMnxQrW4VPsSK+IVzpHv9MJnjUaYJreNRsYCQ+pLcz3MnfP7OvuWY6F3dbGRECjkV8cHFx1CnYq
x6HNEMX2KLpixzxLmrTy0IWGXWZ95FOJLdhB6bSmXvx/i4nrlZq/KJuHcmf5O6JWutSKxn8obe/Z
1Vx6M/woljouO6y61N18ZpOU6QYRIKeJxSHjpYTS3ncuchu1rJ8zhtGbTQgP1MFCGUOrKJiWNakj
riOrTKN2pR2isFyJ9UNqPsxK7T/MZs4TDah9uEPHfO76cf0tctHLfmUhKRuUQmqYkP7tv8/OVEtB
QSDZYaqdAmEXRzkEyhTAFh2e09zm9Y1/UhgonGAWpEbpaNZIBuhBxcFPjEbuZsR6g0UAyb5k9QK2
4xr1m8JwJZ25Hp7UlI7kjw4CDQ4hVfQ8sEt2a8oTLWU0lEmJpeJU+JYFH1e92ew2TPXU4EpeWtIX
SlwVeRo5WgUNKfF9XpSh1vLQyb3+mN0rZDg8GSD+rHiAEI5Nv/rYBISQeKIjaA1RTWPB31J/fnSI
2tyeKRSlqqZn/YCd8RtzRtXwwCNcEA+mnVca1wQecZ2tybHSgdmR29Rnv0CxnlB5ueYmT4+AMwly
TNXa2G0aJ9eQbTtYj5GADyaiil/xRk4bbcca7u3mOa6G8kwrYWdvHgtCFMWWp9s/n6RebwX1F0q0
557RJXREgbUpWjbZpEXiOaU7yVZvRSUhaEWRXMCK7F0h0HCw0X9Iqwc7NMB6obpWjcPuVrezbs7b
JOe2p5tdAdSA2u7yXezQq5W011oZHkXhVDE29nrQ4NyZPF5425W0RY0PzrtwJzzXYQW4s//PmxXc
yHYQe3ItlKh7cDcobcKSFLjDHtiWPhcrvsb6zjdQ3fV/xU26ZIWl6xpjrbbbjigmo9UzfNN4lPYM
EPBt1CTSlBzdgA/edYG5FCL769FJLSYdhyPDuTerjB8IDXnTkQAiebdOx021M3pfo2grajO52HO9
hwkQyo5yZO6t2cHN1imf1ZLR1VIpcM4/ZywJbyjPBGrhoQQYEiPDa8UeLbiXIsL1iqFgXyC2spml
/wrMIooSQEixrqxTmr9HgE3qfysUyVm1ZqtOXwr/1V53N1JXfssniTqSjfltUkIjpkUjyEb6t8Jn
X6kt7ZWS0C2asvpskyYB25g3akMQXKxa2DNMqkM//1NcdyBtPgHAAiei6cJ6Xf0rd5PFzWxP9FdR
BPlno7h03EqKKOHknUEXhTGOdtWmp3ff8IdXyKaUItcYrjnS5e0ZKb2U9h4tg/uOsyYBudwus7b+
cUG2AtDEMh4j+iGNtfQV6bXTqPr7m7pphhYhm+ZIUBNAxfd5FkCOFrJeI0FCj6JUWjTPX8VPVxep
XyF8Ku9aMuIFXYfTcIRYIeVdxeaeEUvJQI9EmPFsEv0XgUDAqTiO7YpvE/xo49eNG6zTuT1TZXQ4
sKDe5wXHIeZRL81LO41I5cx5FGZSefDeNpx1wSgHAKB4RlrEsCbAKOb6fsvi5ytH+VnJy8pa1XLC
XKx7C+9/klMMKgnUJuPinRTsvJb4R3nnqgs5YjCpRYWrRml0T1Ntm38VDaEI4O9rX2omt5VT0Txl
tVOV/yt/4cqZCmP18RjR/OYCY415pap/5un7BX44fLCtNTq1I3Wgzpyp9f22ewAVHTJTWHAW/DfI
ZCa080U1udBmSQKTNNtABDmcZl5e0w2YaKRDDeg/1y5QQUjhidkhJffYlqcPjDC4F3m1PlvkKi79
Nr7xWXB5RPDk0W1LI16/jWMqioQw+gGCtTI4RbG64t9dhss1rsY4cW/6YHArPrPrYSUr9h6T7ajj
OXGlHWTtNoNSClCq45l7cgCWd2hCIoCdinpRUN12Y1HQKq/bh3TzPTQ1311xdGdyyS/rtCSDKzAp
zrsC62SR8SCBfgBFZsigM5vRF2U0Ncr12iUzwgYecz+pVxZhrLNfsrMjwI79bsCaoSb3T0Hliin8
q1hhvZTHsms+2hUyLUJV1BGCrpEQXN9oPIpBj22bvnUcnuBeYU0PLc8998vzjO2NE0zM2GvQhKBb
GsKVAmG0H1ZCnLsVEE22fm1Z7B13f3ALx3ZEidhkewI3NPdSruP7gIKb+rGnzXN6yu82k2/IpgXD
fEJYxPUMZneh156kqkZe0+P6USmh+czmGQRoRc8fxjKr5/OSrURhROnmEBxGWQG0bJ55KrX6hyaa
mLh3upo7wEVI1xgBLJgFShBKbVvisd2addQGwcUoZoyDB4uMtFVRigaDjyrBU+ookvqvF1XUE76g
QJ0MOXRCUVX9ZG9JR989IzH7d/OjA5NedofRfcc1EU18j/JFJ0dv0E6Bis6+b2pr7SqzUDe111Fz
FMqgjpbrpkpknx2wtJcIpzA8+vZpl6Owj9MSHtx0mPF/0TY0o11MFMvuBgsGQdMymBSj/VmNzw0a
iOKFSqi0jN2g/pN1J+MhRqR5TT/HxJ36Z2wIborPRI3+FNTXuEIst9mNXQSoy98bMwUBFdPF48G3
G0cIZvEDob825wBeMoZbtfjVGfRO5Li/BRLlwyXtCorzBTxaEFRM1cg5Lcf4YKPu9DwiwCHN1PzM
bje1fAeOJLUl75OSFG1bk9ygFU5Lkl0DSEZ/t5Kg2Z7Ino6GJLLyqJPpVWhPmaQdgzjWUrKhoEeX
66KgmnXHJpP6idks4k8ltmXQJTMmWW5NorJX8RnB/J+VVnFYW/E2FPZn1T0i2qRTCuxEytcGJ8bQ
7n75QSoGD94HgQfKdxhu8qHZ2sl1mCvB9ihNcnCax3gI2eRBmtxoAjMGCRn8g1d7v+q8ueRjQYXn
yVKZFpq7md52ca6IxOqz+CXTemD1QQGlD0Qz2xkiKjWf3STyJw5ZbvNzG82QObU5V7LoXiMMiAdG
puRkTxUHyLbc937G7HZqvkDc0t4facFe65IlwH8xU0mB+8sOGiuWIN+jxf7PXM9v+y/ZQXESWumG
ku//IzjtS3bOMIdJ43DanxbY7PgPsS4jCz3hk41n/N/89eKW6yifKrJHdr3ED5DZrXqW7s8IvmGy
ycY1pZNmLP2RmbilFZgzUWExTmRIGhNgS4lYdipZ/PQa/RDGCvGS/3xCBWrTlopeGVy2lYDEhsfm
8QhMq8m4jmgjZ/mEUS+1EVny2cFGVIBoWqJ/RMRX/Z0kwI7m3PI9UImkDWqS/V6OPfxC5rP9B2jc
ovU5ZG1ftv1Beaz2IXIuX+RQRvKTeMOBHNRxbjXp7kcpwqrx5tuXVfdwRrQX7CcTtSInpwMtFT1m
/Eeb7A0SUlosGFt7f3ITITvXeX5hpYvgdH44BDtPdiGtsuTTtyNDQ8Ofotqj251XESBhJCXFHGEt
IQOpZ+hyLV42a8+mMD0YCcRkrkom825kAUksqrCadYXjsxaicLE6rrYSkMb+96KUXDiVLwgOqf+a
pVAsvjzI+6g3E8zvWW7O/66LmNIjk5aamdZOaqRHmMJcvtXncuLGH6ynEhYaNez0PZQo9hHRJ4ss
DiWiYUh4oqwGh9Ax4KJgCiQjM7zgbIMts72+aFYgh3dx415IaMcPEuwpEkPimfLPc0cvX8BLoY7J
7ykm7EVotDDmn0aM8L4WKBLSlcBaTClzzZZ2rScISJXM82xncXOe1hoFGcxThmQ9J9PXqI+J8Ur2
oN1M6LP3MIvekq14q4V25NGjAhV5nLBMun2opxaqCJCybuOk5bqG9UIVvsbfDxfp2JCYOQ8lyJ3s
tjmGGsLGBXipP/dg+4ltzUK/4B7NoU24llZzCqAR+oblQiZA8x6KUL1B1wAwI1ig9TxBgVze5RyA
QeDXK0MurkVO8Dw89Xe1eyzj03wyvq0YnxOFloinMNTPMX0UOE1/WhEmuw0GwaDf6VYuZVYlLsH/
k8xNCtK2+oTcdpYARyHpuqXqhB7rkoPZgTz5REG8hh78k3dCy7G0E9hYEbcLjDvOhnWj35TRB6Vs
Jr8XNx6cB2nNEPO0quGxSgLj2GQzSsWciG5XKOSDAalV6/vP+radvW7uQnHxJHJGrQEIw+BTpL8W
ez0BftcCa5IyPo5wmKnGuInoAf1+/vprvNBDY1H3FEemNfhNVvz25JgNpIbsoY7JB2heg30jUd6j
BSJGwf0321WMwbd5cmJMFSx2wPbFnOxVT3N8PDzrUopnHjcQR28EsmgalNxyNTmK0Pybed9vwrSP
xtZLM6+avZ33PQz5+DjXHTuGA/085IkUUKVWUsflDDFlN+CoQ79LTLbA0EnjPymyLibVVgP8uK5j
h3bLfL/tpyrtdE448q8EZkj0esQRa3Ko7jMWdIZcKZlYyhCtNH6T3Hm4rjPrn6V9RW1y/zl+n/d7
PCuF+0SN2+ztlH1CZzsG+1c6/4xeV+P77uQFWKk+DUN5Jxws/AzUIm1AqGnuL/dCK0dIaex8P92p
p/DE2l6YKaT7xZdNbR8syx0Q+Wh19JBTIz8tBG6lpxU4KhT5FsSMvnHZm2pw9MziBCLNBkwQsEp4
/CConuLSzQM+/rT0ejud3eoZEfopVT8GbFJ3t/FPtXFBir06ZBYe/LKD+6DUHJNMx26qL/u/+bp3
ez6Kg83DE2ufZoMI6/bMo0XKgU/QAk6/Fbq2fwX5Wcg9qn5Biy6E8Pz5rwYMPSMOAGGVHy0vEJg+
UduU6MHKt3+Vj5Az4dntaNIURqqutcaROgK3xhthDniS3i5WcnSDfl+rvXurhlHkYo4dkQJKfPgr
z60Wi+vJKha9lYU0AdEwkilX0KFXOHdavubI+tnsvGLZHlvmJ+NkNA/+Qc4T7GIUqCW+tAUXiZAj
K3pL7huMgu8VHmEE9/JTxVq26M9Wmfb8W32rGCiUYboo7P5230QLD9jo+n2BI2/rgqzoChT7LS5N
ImUXfCPcPO0ETCcUBx5XCCIQGZJwDeiADlfd4pPjnTK4SM3DgT8M5JE6/XZMK3/dPfJqg9SU4/bY
75XffiU2xY52fKHjlrkFVU1htosj+X6OHuPDp+NlnIEBWJOA0vDVLGhtwXr8D6GYQCFzBHc3LZuy
KA0k9u51yn/ng9WoFuNBP5W5+vjIZdC/5babXAkZdcqjOYYPXAjDrfMknz2h4zScPziYZKpxqDtU
/WbDuDPyK9JXMcQardHB3lI1JcTT7Pi6DTlXjFHk6bN/apruC3jVbnk66pbhDcEJ4hBPJavR5jG/
wPkfrR273OM/cjoU7+Fi5cSl6p4muWtNPX8PvxPgrx/z1vYwa1Jt4Ci7mkK8ftcKskab+S2fcw1j
PLliYw8qU04M8SMCPfK0x7rpXhU3H1GRfRYtD6qFqt8uAZF0GvNP7aXeLapHGU7Ab6YejY0v6gFs
RhaUkHemG5Qt26aA6bEiSMpE1v/ukskNmh0/fmUguLsuSag5LL5Hzy52YxHIh7Z+9KTAJIaiieLB
Uev2zE8qmBGKlHLZs2QCOBbdsIWdOHlAC2zDdDkYG0oF8WrfCsI+x9+/umGKJTSuspdOqZP5KILN
HpKz3DyO83JyaGe8SiOVMvpILfAT4u4CjPJmcynflLiay5o4IROxO+9wYqKM2ziByt3ko0M7jwMB
urrZfDh59rMWhRD7CrBD2KdnGuPChVfvSdvNhgJuHsUll5VT2/VClUHyvVb7KJS+G3mvzoDnx5lf
n5oiwWdeh+81DeYk5SsDZjAtj5LT53BoRC2/8uLuvw2qNzsX9jioHwXdsxOPpfpHtvObbBxLU7lr
33T6DA01l9U59DbAaaCYGjy4CDHX4DqhoSpz/6MHDo0uT6sdg5rmEniRt0xVsyCjZJ8NFxxOU90u
SPl9Mx0A/VbKUD7xaaUHSleh1EkoYIgcn3mqsmjvAbgBaraX7CbVOJQSXXE0Yej+Vdbx3Dj5ZRWm
J84NUP3yphATtpceFTbNwutBxsq15sBM0PkltMwsZKj+02fbClQH6VrnXqxJrJr98KXLNmxNVupr
SGBBWty+EWkVnzv5VuDRAAV2Uy2n4+lIfBrwD1rsaIyJK4f8y7ryxKJNSRdTttuNlGF+gDgfrG1o
9XZDc5+5a1ch2X2dvmM4sboUuIWsi7jP/UorXhuBJIvlcyUyTA2t3ipOCJUadrVD4BnyTKYJ+8KQ
pb+4Of4Xg2q7vrStsPSRqRPmS6hFNnz9OU1+Bq5KE5xNaCh0jqMiUemRF/tnz8leTuO9zwMcS9O8
Dvf/9VSFm3SrhFynOtZt+vcVPsWgk0mlipkZS593Et5cDwg73+sKD8A8xs2IxHLOEgT7F5B83c/I
fVQu0dyu6+zUA0hFIe0wfrG51oU0PVWkkM+6P6B5dB4dES+OBmQZd6uoCsqO052O5nEuu2S67e1W
aEhwqi/jrQhmxSRG+xcgPPRfzKyiPRyQTbXvxdB0T1/yQ/p7jvSPAP+7hjL0lmj6bMLymqhtvp8I
dcJcno1XTqVFBAS3eZrD/DEPaxD8lsdHOyrvpST2y+CiWxBmqbKjhKR8PWMckCaxJ6WsZG3kXNi+
qWtFi72gpr+VBR3raDfqFJJlLnsr4dURXygOcThN3U2Z9oCLdleAKkHu7mP4lP4q0xi//fKUmVwe
qnqs2knZFASRWjRIAxyEe7RbFHaWoTls4jtn0xaswJ9kfcpBmG5BclII+AzJIh/vcmyoh0D0LY03
IUSJN3fR2GCtRLfOq1ZK8UnshDhxqPE2lsY3yJg1ajK049kxwzr7G38rzQwiXLzeBTO++G/Zpit1
+FLklD7hrcRIuog5IOLDvdQqtroPx/QVl2YFbbT7yo+xITJtu6XxHciSq55Rn8OF66+jvC8kgz+N
YrTXOdRTiVuWWifMMAbPNaFX+cHoaf7KtnQuOPMKpaPlMB7zUCm4qVYpM8fuV53faaeO7zcg1yuS
EPc7EDLOjslNjuUrg5DgSpWFbz+iE3jzQktoBfRq9gyat014PS3IF2PMqC2gZil9pwCg/7wmby4A
LrL9E0xIVzb9C8iO0ibaGWYuMHXKl9vvi+8KZJsplFhYd8Z+UP+4RMF7e/CpXIV4z8sSPUBhqWHO
hrf08tz9zwm6+GFgOjNn4ND5QG9prptCeW0REPVYpnqWBS/2VNDciF/A2OPyWx9a8J8+4Jaw9+8N
4Nf9XlPeZiNmoZMILChUlBTT8BxTowQI2K+wddpScmirCJOgXpLPJmvbX9Ts5vpKmtKbQv0jiEkJ
jzNQFggSHFY1rhYztmD/Z9AHoLxaX82pqD4K2Wx8tn3gLFdCvbxhkUed4w698mbnzz1PopdjK4sd
gnSSadJdh0MvvlPcQKE3kZ3ju/3PM2lYA2yppSJtKx2FUN8eI/cFaI9WU4UD4t1GvGZ+hGhsoy9p
5AGB07UcJQ3iYsy0CmX4cIOPcfWjCPYHzXwY0hnPNR2c1lKRgmf+8b9AuFsDD+2ROdN3J2HJSn56
qgra4pUCqUln9Fyd9CVVdZ3Gcp1+3RPVJCj+I1RWTiB4pe63PKeYGN+cIduEdXtviVaPJCCSNEwJ
rWWFWKDiZQLGjJNXX+AzdBhakbMwqU/vL21JvuoTgDz5Cqu8LmFQDj+Hc7Cgu0+aGMqyYDJ/lmP2
oJpz833lkTDTkmW9f0G3UMnm8rrEzRjFq/17hKe+56k3n1ZvBEBFPYif/LcQgpy4eSC7BimDA7+X
/K3DZLfDL1v1SzJt8k1k1XZE/jFNENoA8GnF3nQ5C7iT9Kcx4Fza1wvSRO3McwmE85FZ8Qi1Juqn
YGutNOU7u1BdKw+zDYVcNaVua1OkR7AQWuETWsMcow+rGOu8oATyWY5arbm6FQyc1WQ2gvgHh0o0
GUWPiRW9nF09lGcXl65JzGst2XAju3IPq8TZDIUEtj86X6HEkKCWt+41j0oSkc/7lzuJNPTH4kk6
x9BQyGnT8xPJkYFeqtsuon3b19NeQRnVSxg0oZ7X2m8Zw4rMa9q6i+REScbuPigPMR3wkVOjRh4V
PsDGzpSoVZFTVDdoZfYhiXH/JK4ftCOT2IEAMP5Lqw3m/RO+OnVPU6JcXYOE0Lh9VxWPHiPZfgha
SmG+1dGfecYO4h8U0KH6gUjLFi62aL6Esw+dv4tIJGKkmuwN/iNKMNM1BcjAs6jnk7G8yZzKOejM
P65Jtq5GIQtE89G69IhiBGT7EyFwMf805kj62O13imlCHBq/q+H2voOyVYU+3Hx0yPh3lEjogTEo
iuFMKvh6Lmfrg5p/TH4f2NXHId4CZccv/ihJq5dBRYanuIJYDnHsMitIz+fI0e9X73UhjnVQZftW
iPEgjHFHYWWFHVbHLlKk0ekOdH9L2FU/jfK0kwZEqpHg0h+1V787G9d7+v9oVQPPDOxxHnxDXTgw
JoWkpWxVjOKVnYc+fe4Y3USZCeM4T33w0ncQQfKymsu44ZUtOHzMdWNmyOzeSDcP41+sSY7YirSE
uikPiwTHNP5l/hLQnopoKXpYYqxljsPSZzcZjva0VQp+gXHpoOPfITtycTHCNgNsnUVzspnb3nWg
emMPOrPpUX032C95yF4unis/ejzYBOQm4X6UpffHSDAzoauAzxTBBgNv9RHHvhVJrkfvcy/vh5ds
WOft5IUsfhFn3Qb6cTcbO/o3reOepz31Vwur6o9KokL9mJLuiTAAvuG2j2J5dFhwMcY70kjP278N
Yb8HCm1UrBGAJXiYT+p7eoeYnl+1ZwDGo7WcVuIlPcFuK1/54TwPlMgnoRcDeqcLu99aDw6pQehk
Gf7MhitRsCuux5pvtDiAvP/pg+12ouUWNXk6nnBRRrkPljO8QHwdsSx0+jLSK2RvdDNV3z5NRsr+
iiqa3cxx3MByY7CoQYG4boxEKQPx1gfc2mwrKMwciwJ9IOOqVjbfRZfq5A6PbM7j5mDXy6Ib3yB5
n8k3xV4a9Hf5xUuhSOfyLmpa+uUQW9umNodAF5U3a4R5VTUfJgJlAcJjS2GRpPlvo6Mk7f2TXfJk
iiH2zBq8L83QQwXonjGUgsZOF9sD8vdQd/czZmqdyJKxImybKN1dqD+FuidfRmPzru62i0D9Lxm4
wAp2cv3rEzKKRJTEnCTlN5L4oaUsuZ/itI+RgBy97P1DtgeEmAdg5SvmRIsQZpVQ2Ok1M/1raKtT
eVBHpAYFGwsaVA9N/yCRiz6MLOFeFTiFcoEdSFFm0piTmtFLZRNiInyApx6/zI9guIhi9MAKQFVC
vv+skWwYthSRnTPoYgyGn+9nLy3cVv13wDPGNPaSsT/ZHEbsd5N49jM5MCJi/0IxyStibAFutJUZ
yNfEhLV1qb58JypGdFY72/QtEfQFzMbPK6J0UcvyNI9fFGSy+UiJZmJsiLL0zIum9MAH4SLATwFF
FyoUaftIwvIpgaUbRQhSNF1n7FSKzL9JaG4MtR8GvmmaPriMyhzLamt/ABgg8PfkALld+VZVQNNw
wauYXS3ta1cCZckt6KxuWBj+pDg7wLubZILyNtffIMxm0FigLOA1BH0IL4d5Z9LxfWSp+wFKDieh
CE1wzFhvWsIWF0bndbOl5z7yGCvF7tdr3ZwkqzPFlYqAlvNuOmUUYQSHj+xYo3TjZE4PUSb4xSTo
/w2hpOFMPhaB90DBoDHokMwOLixngu4veeKm5NJ/W/X3a0f/Dp3G8Tt7Qn1emp1b/Bx1URxCLtDq
69rlQlp1XPeU6ixti8MFgjebNR1ibTHLOlpLchqZH0bFooiPj6WkP3aBsFMAOvSNtyOhm5eqKEhD
KIC76iKAhlLgDgAMQuVmG26YiCKjfoKGWiw97uwJYLMGaHO9xqSW6P4zMycrlIsNJYrv1tu3DY3+
OpaWfA75BSMUuw3LbmmNue1FKBsny/CFO1K+tznBvMrOUuGh/ty/qv7DV4/PZ88WlRITA4JXiihN
7PiFm+KZ4t50lZc6kkDX3FwKthkyT8OBFlgKMB7OSbagTiVhZ7F2CB+Sf4kWiwvsx8/FhgfZxiE2
GiIIB6D8H5C915hTY1JEmtXCznreZMnunRu3R4IALI0K7KfGvNWA//vKdQA/b6IIbKyVZI9LBFCE
HwbrfY4koL44hZtDiIEgwzeh0QlXnwJQMAt1LnSlSrAMrw6rQTwVfxRka2Cz2FzHaI+5TZs9OEu/
iz2makcpQaXxxjKxUd2/EJIVhYtPtBVFAcA5M0BSgMovcm8ow7f2UobpwkuYEBfEZ4k0qBpAhFHg
LgxC6pdE7sTUrdoH6Y06E9cWGU/+a+jc22WP3s/iPDBN0lxCF04uZH4h9qH3m4fJfWbG/japvPjL
TmuTdsLjinVKhRODNfmjtoRMfsgIYHOxaKiX6xSwouVmjQ8ZRmW1Z4FmPBj/BEZ/wBed21hT9Meg
IcT+IOhu9wEH21uKmBGr2nQuVgpDtjWxRpBwJJo0WXJLE5HrBYzzMaqxY6WkAixUSFid4t3BNGW8
RJgUBNnGvkBN4u6HrEpwWGerW5s93eb4Ptsg58kLTqfZcA698Qz7V6llKQrokdAsV6pJ3GXnAQQH
NY6LIh7fkZY8+hcCTcYBhfzbtHkdiqOZGO7xKrr6qMaMGjKTQEURTLseHTGWsRWiGr6460B5z/c2
j9bYMlNlFFYaL4y6RHcClkx+IZlH6IMGsfLsWd7SGYySMHRShEO0RF1cxvv9U+7Jxz97FXhhBAsJ
OQ9Z/OK6DfRIPgEkBpoFsAJGZDiBPSdYEXcbYhUO7rGj6bkP9i2bVeqHlSaovORmEdDnp21pJ0/S
lSm0MDlMZPZv2TDxmX6aU3b7gDw6kHTZRnPiOEpPO1JBo5woB1Gh7M7mbRC5ykM6Qs1Stp+zCgne
6/oNJg+00ZIAlC/X/JgDKap5UKEnIE6fkqH9KIVWRs9d4JKBwxuDousBQ11h/E/RwzkwLzcyo/Gd
Z1xwuMPaqtr5q/oHAngtDdt0WIxwykCtDco1+TigjdKdAuHkWb9BNyXCHY2l8YYzHVPrzyC1CZNr
F/bvtbdZPSIJpuccbFEM34Z9LhFg/lNAiOiVUtO8kmCSui+5PmJF2skJnkJIeEdU9Xk8GmU0r8aU
3V6+NwUfI91uHIxCP69ndAyNO7cbZ8uR6aykQKcnX2eGdlTZd8iB6P5H4tF8BaN9vSJiho+0h/b3
w+c55M26AKmYm02eN8tAqAKXmHhRC76CwJzRrS3AutpI/v8vde3lp0CwIwvzKlr6uA4AkDgk1gGO
29AnJPxZlif+XGPp6gKkFKDeTvEf1zh8k4RtUniRfQp/O9c90Zy4EsSZR68NqAahgydU/6SMvnY3
sLvsPGg+6d+suz6wT7buhGHExM4E1GSusY7h9CBecOtSmnE8cVdwVsepgxFTjaNxJISdxAuQQdRE
du5ytdL0vCZ/e0K2SV/64TiWy0milWw3W4dItJ5BGGKZljlfe5vWPYx7EMlrdlZGyxDA4z8zF2dU
u9cckKAA20Q5bWv0KPuofIcgJUjDCy7Vy4092P6YzOv3Q7tvCCPBXu/TenxjxphtdOF0y1Fodi8S
R/c9qZViKKYE5iKzmfjIWYYu7I7U991WMxyHAdfmAFsLB9KdJcLQwumb4uUFnKwvkUFtm6k9JJuj
JB/EomI0N7Xg7alZdJYl7DgpiDwVQ6h57pnropftfizuf49cu3diY7knRp3y/082qK75MJjavXVi
J4+q6q7QYeMqn1Plm6Qo/uqbgEHiUz/n0WWbtKk2s4nuv53JfZBHjZJahJ4Siqb1NHKRz8XXVApP
KSpzAGPP6781cRJrPj9NByTDPKhm+qNPrJgTq02a+3TQFEhuOhafC0p8ValURUu5MJhcPYZX/JXs
PEoq+zn334U6IUJ4bvyj+fAgNJS7eh3q+b51Pmc9FzYgcC8N8PgRcRvH4ib1KSRdjhQhd8YnoiOa
WSIrkdGRNxmInJxfRFGcvDIP+kyBSsYV99TGx85oPXxvH4PM5XuN6eKKtnM74LxcjP3s8+6ALPRZ
/v86pO2K1T1RSCM50ZVXGz8jaUJ010hRy8aSwKjkWO2hweyOfK6gidWI3NrjRtmHTiOhXDJmyRNJ
YKYFeuuDQMqKeT57E7Qp7FjJ2xmpb8dMpFr95B3WnwyhaJnzT2Pc2fBM0Nu8IO6pxYJfrUgCeZeb
L1/np/3JIau4ZVas3T6TFKyaXVOVe00UwEvK0YeNPOtZTC7Sh1ZiiOrIuY51fs8Brbpslma9yVM8
cOUJtOVhl0cTdcdMNhr2GWERy4bLc7B/7/LqAC0UF800y9tbVfNhrteFkYL4xJ5ufbLgPieYaMAw
DWmF1wX9q4VKkgAfnNDDxbKBdYxlRpD3vm8RPqCuO3+f0AY65QDqfpl/vye2222IUwaFN7T/691g
fz4Y5qcAx4ViX3xHTlzONN/Gk9S68llqb+xyuHLO7oDeHxGZq7jEub2LpztO5o2OgivvOYURAvtb
ADgyWD4BQhZRbho4Zt76FRq9QWmKdHmhexYpGdJSIhRbn2qXmwwvK6c09xIP1XeJZnqfQdPYFNRU
5h60gMdQ0eUj5bGRse3dKQ5DzLMPg5++GXRICLlyFqGb0NlRVEvbAs2HfXy/JDqtlxpxJuEAqV+v
CQVTmLnclBnEAOZjgW29rdqFmZkdx+nBuHuukCrSeTETU/1IvUoochssB3pSJwXX/lF/eAlFAXqi
aLBpTOWQCEVlBb6olht3F2cf0y1W3LESzJxLN+EfySWsHawTvkGYAmUIX5pe/iyCyclcTRepm3qh
Jl4J0tyTlKDsO6XC5bv6Lm3SqmPR7U5qY++dqkOluP6zCjO6VUKMCOc+nxwtvepSmVNQK+yP568K
PEfIMXGMZMyT1/4cLYBFTa9iPoybJLYoN1Oz0q4hTBcsb0y4NIfzu0YlCQJ9cIvkVbW/ldFgfiAI
TCXK0+P7Z2f2cgZlBDI+2nuQJh4B3hlkyxovHlv2Gjw5GCEJ3Wv1Eo1mnBWl5TiVsjHOVfKoF10K
hMAY/CQfET1SZw944PKEchdzdO4Rqf6P3SihGpqKUppXOmIx/rGilp1xImb0zu93gxd7z9FAvbiC
p9/7Wl2dWY2K7COavHvTBkrs3y4fMHWQfIaDG5Q1KelUlm7biUaauvimIAYPgw588nn317pJuYAT
XVpQzvh4Qky/5EObIv0v+UOfkkgp32kgHo1IGNM//8Bv13ofVeVqUwYlVHXjMcvjPf22rLwOvuHX
NESDv+6b/BnBgKyxB7IhdFOvmwXNbBdFK1LWLm8YbJVdEtvvj56QG4rIaLrCF883BvFs8U3BQStc
dAd6C3BVV6t8bFcl3dNjgVTNBXc3SP9ojkfubDcrn6euHVBl7T9nm0CW60eq2RWeq98CQYJaDls3
CYjVPTnkmPYpIezinf49rUfLT0Fb7tpzCPN0OvR8+IJNe6jjbvDOz9KcRvNryQc26CWGF6CXkA1E
QIH6XTcpjOFM30BJuFGe253nfpw2BX12tZJodfrm+89blg42NZDE3kfJfE+0EZJsRFsZ4wGqS9bM
gA1Hob32wLtiyM/5nCOvTMoPIW2KyT9iAU0AVacR+3+NRinKdhUpP5KEFCj9HAKvnAll36Uf/OrO
uN9vfRwMGdzv/j3VRJnSqWDzCM+u+yL096yGVJXBEoaULOwtgwdNkpHAbg5iAF0Eejfkx4qo3Ue8
Kqd2R/hnqDGmJUvkmjPIkACyXXMmX5qVHxKQqXUWzvPB/HIQARa0ZSoc+CpLyrqVZ17orRWv3sS5
apEw3K2dK3mCcbEokhvrnKowSUU9D+ppXrLomu46smDgsV+KfggJt88tyn9/g/IW3Z+licc95BSz
zzV6tARYXBqaowRkCs5Oljgqo/0krzn/YoPRm95dwHPVM5bLOQTP9ApxoImvJd099wy2qtW9B58K
hYw5vLxUUNObGrXZdYCb96bysV6jOirttPrASQjFnoBJOx04QmJRra8J3bIMh2VEd/CZV6EJ1eCm
4zBujFIipDDfEMTZ9JZYl0az+VDywTzFZGvNgmXswzwDOZ/AQYyowbFD0ZthbnBSQ6AxF73m2qfw
ONQ2xMN2RLK0okpvzz0SZLU76udegyx1zvwZ+2pPsIAMaVo48fLlXLw5sv/5Wj215Td1oQSF92ez
F+90h4/Tqj020BFxRZkpNnK623hiJ3Vmjju2mLMhxfK2KR6/jFrJDmYyM/fKeAkY18rY1ksLXqAN
q0bL2lbmOOZj28FycAh5KwK76wnvgCk5IO2nzzUnjXCcHzM4nP8aQbNlcNihN16vCVj5/CS12lq2
7Jfx7m4RLAjdsDCnbEi9hMjcg7Yx+oJQxNV5vUNwh4RrcqnceHr7cXnJ97qyZD1/OjAR5ggz8xIB
xCTAsCsTgnM6mbzw3htBHdK1SCBFZVOBrF1XYvwO764IizP60afiUar2XfortEm9/3mJiE/y/Pp0
Sw52xHbXMrL11odH9iaPCPVFjbiFTZTrtOdto/NQvF2FudZMM6HbB9j9aiANPRS3EV/1PnK/3T9P
cnRl+fayu5QIS66xze6JgmLAZyTXPCW28YRA9Ct2CWPp4RNVs86cbayn0EXabaTOoTFZ0H1IM8ak
Wn3giK3qp9qaeJID5SLgLzuPS1fGTjftyc5NvVqrE6HmGyEuI+WNM/OqKy4B6ZDHsz+TzdURjjYt
C/SO4k6r2buCbWjMXFG5qPnXC7lVxs6+OUCqD5BxV/PBWKPhXAImnZ3M2mIZnBiLQdFwGX8ZcnY9
jI4xdsoqE8dCsLM5xLPkn0hJMjPKqp1NvjAcjQpc37/0qAWfUIgxS9YlVQjIWOMaPfZwqnpP3vkg
btOqmJk/fcobAK72Z7YCPmFCoJqrFERSovZ1sLZkoknLP6ZXfV5mk0fXf8r2q6oIq7/20Hq8rvTb
e0LTLz44g98qDkc7rLdMNCY6dg445NCSwBLdcJs+G6r2SxT/ifF/ahWUUD/qZqRFumqm7uD+Wb/N
AATWlMPAZflCYGx4oYWQ85hTVQ3MM4p5KJ7p/9GUzk0vwU79x0t2TCJhKmXHIWNs8ViWOLPdGO5v
6r2MAOpCH9ZGSXlPYWlCp5kLMnbdGotHd7A44boOZ+QmjDHJIkrBUrtj39rUpCovj8n1m98eDzjl
LyCY5jz6Mx9RyT510hd/l6DxnNuN+lAtMs5v2LvGBUJDbKcSO9QAOzOFe1FmTB42u0n13LOt8EbL
rxChL3R3/5KBe7LcjaMZ3FbRCQvC7pzJCo4uJkQ8SuU/7NCda1TQ2ohez+wxQa/xkZS6JjcQAbIq
R0czGYhKti4aHe+lUkJmmIaPio8V4PRkIvQrFyHDtIBQzv+RZ8NI5I0+9roeq6P3hppMgXQpYDtu
6C0dBdaNUzayArUUJ2vhl0kzp1GcaBdYEnbPT+0fiAh8K+jw56lwc0tG8LxmtWxOzuYbSdDRBV03
1TY57++PPCEbHh/g51d+7AaQrKMl4s65ErlWsWCDTU8KWUbolsA833/yVpABaZwJbeB6H/5Y2Q+E
hO6lKrJEez4/A0tA+j1aEdcSd2RsJfxOkbieuQ0/TsY/mVPXgJ/Tl/OQXoTuQoBBBhBppBBfr3/U
uG2wGX2Pjo+NuVlYlNsOMwXnrmTbZy2wDj1KDU8S/DVw/cIHOODH3Ttsc4j6+vyKV+nZbSOj5Wz9
OUKcrxMWN9Na5MzZWZ4Juj+jmdymOFID33HfJ9sniJ+FcD7AeSo0RVXfqCbE4Pu0AyfJU9UDa6A5
tBCDDKUKvX7ITEJV4T1TU90VoPnBu55JJyCz6Nvgo20S/UdEigmuxpsOjOGrvNB9PkGDEgwrPd8j
fgxEulMaTogXBaACcLh6UUPbrfeiZpp7BVdnKx0wuaheBFzP0IorY6WjG+naUmmdj4EkopnMcLFK
ojqmGeAsjik7tuWpiKYqGqkCAf2zv5RfMmm/HulwFpDpbSseYEw9vNNK+iwzxMCJPC3pW9A8f6Tu
7/zCU03Xq/jvoWxZAD4v88mkqz1jAQAClcXBU6l8mg7x3gq/lwx0S5o0FOeJR6ewoQniIOSODCcA
6CrpxQYi0H+rZHyatM7C2Yx8K7574sKn/MgZfBIhKpTVlfX5iGm4ZceB1cIzV4mLXqqYtPnduxyS
TxYEPTa88AXPCVr2gQPvgAnVTTN/vJuCNm9XrFwRyehdM+dVPQTk+mH69f570AaBgo2rna7PCGay
v2PTS+E/pdgs3bWS0S+aNeEuXjWnCU+bwHqDESm0ZefjuWswXSCeTrAzRWpqa1nMqC2bo8ze107g
yHLs5D3SDxCXAnlircoNdSRpZsgWvhgmS0zbZjjKnZzbeogfYzeitOq/dSCpzJaH+qzU0qtCH+As
t5QugQmrdFJ5fBzP4EO+SMFXYB2OxKW3JwfAlM2rEhS7SrZKGk5tbKZVIbE7KZHZbAyt71feW8um
pqPbtpRPVCxqsOqWL8ZF2CHoLSByu4L9oJHjJR8K9U2vYEgWan1db3PX8n5ZRNBCJ1CQ4S1NwvIc
vhrtQEH8Q6mfM+JrKZSZ9TPZwsCe9I60qQw9L2qBK5Y06rwRV4veBeg4szKC411ZIKWnFXYPYabe
r1jUl0WZGHBrem0hK0+c1u0E2Yv3fs5Z5RQ8CHCVcHd26FURBWgVFB/xFFfhAdEWUrnuOw7VB/7t
6kqEHlLwrswYzCHzbSMPAMhpwdYYf1A/1Qz1P9+uKTEHkJUxT5MPIUFnx4+KAjkLvgS11tSrUAw4
ktiOxuh0uQnGpCJf1S3XNP+1wGPSa5OWejvATmfmmSSsczTYfjXtk4r6gRVIEbb5G1BB52j7Krsa
p+Q+X2eIEwmsl6lJSkw5HkE+cnAkRN7JpOuQJRkvJrsnDMUfIeLb5XYmX6jhCAxoibCjlfEvbUIC
5BmAhPxSp2+k2v4jrHTZDcLOuvLFA8UPjlvV41Yp8xUbOvfgggaeWrrDLwRNOrVTMmMk0umKVLsz
a13mA2RyUGo21PXywJT41E8JEOJqstbuVCIpoD4TpEf/jwUDSXmnK6QoqHGjanGA0nxKB/3uFW1u
7YY1S+Nto62AvUAmlT63f1cZBLThNOe+43wglFzduxRCYSrOajCySO2xt6v7towDAQlVfQKLlK7G
YKwFLoSeVyZSx9nd5KVD9No3H1I11bC/Anb4pgtMhhvQRCfbew9bkYL7f6IYYPTR/l/eENltHvh9
g52HfVba3FBfBxNy1oLUEjf4+l8UYsb9L34T4AwdzDllayKo238D7LUw9/cajgPHLeaaM87PH6dj
2SWTItCNlBPjWNiLlcyaVG/XEBHK0zsI0wRcXF+4AqWT0hMr8u6bi8icZYNZ2lBOrEuXZdh0gtFw
6RXgrJhSvabtwGb5NzxzqMPl0aOv9TmlmzDnjwuxI7MHoRyhYJVDtWgAneG3C8S1N+o7F2Ybr23X
hF6AJovl0Kmq8n9cBI3qknOjAHTtR+rvO+zp6qxUiZ0gTcmvmAlCWQpMyrVA4A0PCnlvYeXiXBxs
bTNg1OwukmFdTZsieC1xP0N0fJs/9Yqrb4jmIE+2tcvNJdu6Wwun4dvZ01CdfIyiwWNb/YdNl7MS
wa+ae9EwqtazxKO0BdxEbtNsACu7Dvad6M9zKxdPQFS9vCN/DLmFqzZpwELC73bhmBLCDtci/mwK
4MBN4U0rTmNaPg9KEh8FAw/BlHAuWdZWiMBTycnoJn5lSmGjTyNxfQ3PStneHu2hqKN3QSzxHsbL
Vqm9R6Xwcoq8BJKYTRI/Phu49sHtk29JI3VzKlw/FlsNd3kIi4zYtiHvNz4KtS/z9a/oReOOUxdW
Sz8mK/YirkSOOCkfEtbWMxaVYoww73d4GyF0cIHNTeYUxV3fBMltwgPDQ+qsR7Hg0hqeQ01x6SwO
70UkkhPdo9I7YjkHbHP1FCwueRbp4FRW19b+NvHyzpbR7l/QgjYSsGJtSzwaGaEVm6C9Ndk7Idr7
yjm1ZqlPEMWeaJLdAag9qSBBq0RaILowbPciHGNaCKXTf1p2LWbuzVR5r3YWgYm0j1yDki85TubY
bCTywrWZCApWEg+zf4fTDuvwph8K1Cv319iJTKODmri5ySDIb9XxHfqrVXN184lEwg5lt3+bxwJ/
wwVg9i74xa3IYxE7H9p8cB+e0d4lB9PmIOYat4kQ26DykQbzeHt0qH9IC+LbHDZu4YOMN5ag2Cs0
FturPpgx7T2bkU3tEYaTIJm1QMsRiTgy0AabzH+TNqL2KlSbM72wbR6wG1MclP3CZlJ5VKWkq2DD
rsUvfsF+THchEsRBEZ73eInvt+BeMJbQsHoX7CGL58y0bpID/3ZbDXfpK8chi/r3MzALdbxEbfk/
a4QLx7lHdwMRJkjTCAjQ9ZByhrFjJxVqvxkBhN3TyJ1IdVngGMdnvvQd3xFA79SYWyCC5fqbc7/f
r5vbCyIBIGOe69H2+QLN5CQVOF9f2a5F4g/eEjy0nGM1sAfe9r/iO7iewr3ugKb4kd6BcKhKq6Hj
QS0axqIFiIMyXCa+KaSZhIHKGMi2T3yz4n4pgHLw8SUKrL7JOBIb+lbASeauueYsk0U3EF4HDqS3
clJOrzMhL0et7h74lAn2IwsWe9JhSa2R3tmebNIqLhZLjr4968/ZY7YFJXoh9Paqa9PUwMi1KaqK
Os7el8TLBS82pH7RagtLvccCY9U+VNUZGpqWlM/TwBAhmouXFg5AU6rDk/AziC/PcbI1MUsYLEth
OeAVCK6p4LTvBA4CPLfuLQpHiQCdqDbpijgUDQfuCmaARcf99TiHHNRXNNmtcvKr8u+G151bGbL1
dUy76ogmDiU8Lg36FWzif4SID7QcZJJJ7iorgnH2G5uE4cau/lmtS5cTkp9+oa9Lk/MlhnWSLDYb
pNKYvqFPuH6QuASrBBF6eIPA0S3ud+vR5t2w7smbsfZiCjsQHX2/AdJeFJhxAQHyE8KCcCW4Pa/C
jhMrGp9SgndYr8rK3/d4jDyScqNxayMRbGFVC9DlyNvXbT8CfM372hF4pMbY01qknkuqgWqEL3w2
dhCrJ9aZ3NQDxyuxIYh3+ts2m7UohTjhbtgc5V47jdkUaeSI2amPGW6pRQPUGF8vAGh6ZICWR9AT
MS+HSO0Bxx1AERq6DVBBJ/aOzCzl41fewTHuzGcLqMoGuAJAA7scB7uk+Pf9AYbNy5DO28DSyPeu
tdcTc9NM/SK5AW2T0C34rGk4OMvhrggXzDQ1dJ+TCf6zkgdiDeMLh/rjOcGqW9Et4ylj36s6X5tu
JXyGAHEDsLRKIBwF4/R28M/IUo3VpgFMgSc7oIULKJ5dBhSgE0FlHaAYNQhashuIdNiZR8s6hMFY
Mcght+rTxLZImf5lTqwK1IGzWZbU31yULrVyFu4r9Dvkp0CvuC9xG8yM/1c6JolbhnmXizO9M0i2
SJBjPIeiBF1uLM9uVpy84IMPSqQYy1MsJfL5MPPc40MpgrjVqgkcl0SP49JcmmfcbyQcmt8OhMXp
eFgTFB+DV5KJkzwINSsmgf8K0BYA9TMJlrLY4LPIIe6mHvI4VsPxrNEraFczVt6mv33vB8pbVoLt
IRNyuQ1fsPOQ+biTAnS50NJvDYgBHc8oj2q/KhP6XiLIAqVqf9wz8C4jT2PHrXuR27H/UQ8+8zuV
by5LGvQcHI1y0jV/NsIwlDkuqZyhVKJC7l3jRBNJTbJKVHMFiaypTLewAEnlnJa0IS0n+fk3Xj8G
F2VERUfZSO9vpNfJI9dVjFdH3vy+mgxyW+RMDEyN819NveJiYx5P4rezBJmWWhJUB+TM4bqbRKz1
KEccqEC9Ka0psReLRo/qYhvD9l4L2iX1DT5ghbY4SGXsMymX8uB2zapYzVLEOstBeySDQJcGdfqC
uBsh0x0WizTqWLZgCf6PmGSLXDN3Cx0taRF3V+vaI2hTU6KQxPbByn1C986udJ588Hjesdwsdt8g
mHJBMjoHAnxcMdaBXxDOUuiLFdlxwiGJMdyqguf30Rpd5UJ5oA1ZfLAf9DWjIERX8MbYGd2LGPwl
EHLr2zUIisi+rAy4qHfWgMs8PzRM3qNcKNtOu1UcQbEv6hojZZ5y2HekVbhEhkEW/Q85+SWNLoB3
oY4AmU5Fo21iiFXMkeyJUyrlLgM/SRc2/h8RD7FyUIOrmB/SPWTm4ZnxNwhDtms07Pvf4xxq6SEn
tfxxHlkHUImJR2Gw6kGUj0dkanelqWjMDgqGx5vDCvG+6iu1gaHJQwr81jggPF8Sz7RjWXeBW0VH
FONX+h93bsrc7SL3fRR+yv74hCvHN3CPEfYWAD6NaJyJBGHKcJAFoo6mSKn//0ClIOqCad6zuf89
W1gHBcvaoegFLk7d9TOZnixK5cCHOEwyrSw0nBCutSjF4KEMEC8HAGwXK8a0Ne1aK818eHwI/+TD
JYV/06QN4fcnFoI7tXhlXaqZwRrJeuIad7sNHvvJrNWfyv79fs3ZfZz0x/uEmId/D/1AMB6JdAXw
3DGLT10ybwjICY9+pYvot5hwH+YsZi49EWXmWNhhuoB/oL1mTPwNyWA0Zm22DfpaLpbl/lppJTfR
glKvHgoDP6sE50km8h/Q3xY/5QRJAJx1PUGqavFG4ccttspL4NDwItd1YtpG2EQSVdFbg2iWKOjK
V5NzYllCJpSWaRVIqBE1PtTCkqRj5C4oeDjUYnaBGo55b7dOELF4bc4NlD5ORMspZhvt+8E/1j80
Diu4S491r5EWBE6BjTLDL2iofHdMETFUNnEtJuYSAi73muPdicxkc7JZfToL6lwpl8oC7EfrmIiH
zDsLseGUAzJNQMPKs5VqoTFvKrGqDptQsq681bnrAzSDuH1p49G4cVheIJZJRytjxLbTlHyaXBJP
pCytqrUVdD/dkHVXkW8NRiJBIBU/TgQ4h2ay7Gi+BvcldBOlZ+CQ+G88FVKlBAG0CXLhVCD2fvrm
0AtSB/3fVzRA181STWFPh+wNmlfVLhf6eDJxcagw2TBig/ixLunoq30JQ75PbIMD/kfqskkSDOoV
SomWC3vdZOsV688Y7wR80a1OhC8mLxHR9KMjrRW8pnDZMxpIeD2LHprlcdYtJT4qwRjq+TZEgJoT
3trNcRRbnwwFS1D8xXEKPRySwaxxWJaXhY02XQdoHy465OxVJcjHeElU/tMJOXCQJuU08t7BDwxU
/1PFSpqiBYpklSTjYItQvCTFeAd6oLcsk9ACdxphbvaSv4l/oVMJiFxc0CY98fdYERK5LsK0UrPO
Z5Zicfs2Zehnqm33kygq0Wn22GfI94bfx3SvgpvQp5VpBBTVkR72bhuVlQACCjqVCNSeO6eTUh5j
ESHwZuEeyPR+WsquORNRnvl3V2WV1OSPEOuhyYhVAn9uT8dYfnqmOLLfCVdSbHgv89cehjJY/3ha
yxyb105j7XO3iVxGCuVy0S1pmTFfn32VolO1KvIZ8lOKAV3d1N5p0Oe2Oty0JqscKNyb+QtINeI2
RY6yxyhKeNB+ukPABuUCqLXSgPrbhjCCuB/GwQpgfYYRqum0/wYZSR1M9RpzPRY7e//eUM727J1k
71y2GJVW/1ePiwc4NlX1KHpEvrQT7cZ9du7eMLS55pDGwq9RrjjZxFN32WAUTCtjL8KRshY3DgJL
ni0S0+MoQbRXhMZpLCg/9xSEceJiT+4mKkrxakecrMjuJhoS6i18LSJuisbFWo4rnrnqXBXb8Ce3
4IFE7fIkxDY2IbdvvuPZLhjgTTF/qTRDiQrJ3kO4e7FzMStRopzfr+DYXI9SoxmcaoZS0whh4u2p
5BTWkYbZBbSsEQCWhrUFhzo1bYslHXNxfAvSbzMxzYnFoiKq/8DKJADVP+Jbd0JRyHBwe1IgN5Az
H8scBbvahtsvah7E/HjIlNqIm7xC65PQOvIWhEy1BVjbe25rTSNbSYhK6UNiPL18Tf1NWD2FyVvF
SfE4OEkyGLCgJHjIAiyIeSjMZ2rARz03l6aB4KvkEvc1MudUQ9eXsNe/7bWrauNeZp2l/9s4niUM
7QHKijrBDKvZnrRMYhxj/gYk0bhnh2rJpZzEG8EUesdpR82MHk7FgdP9yOOUirYGAB02zj4fNdNI
mEhzrwScOwGGppDBYE0Rwctz/VDOOJ5GAxmZdryL2LLou8sJTZOwkz4xlPRDBjl7Y5MIAbcMt/ng
CoEnBLzwTitwVT2xxN5lTUTibrzrtJT5C7nXa/oWiMMP4yYgxqL1SmI/vAR4L4GJd4OvJ4Bwyi8O
0T2+XeyrZjj9pZIgsK4F9R065r4knFYAZJRib5NPnbf2HoWdvjw7t+Xct50IqZ2B6Aa5sm1GX2sq
my0sIprwMdKIYGw3CpPFp8tj+vZFB6Mbs7hYj9aRvdX7QLvClrRPtNDJHlrOPZzUm1vM6oTD3DEg
p2QqRKczNL837I5h/HC90dlFGptgONInLAaknQ0y+DmT3rdiRQj+dhnF94qXIy+TOkO+0pHUHQk7
lKD8/zda1kAYkLumidLS7TtAoFRWMtBFHdxn+bFCTtr7yiOJWT709KSVwwrgh1j6VNESZzMvtliM
jrGOOLa6WiIBu+XKOvNXnlxOC2o5D/rATWKtgKRbSQu4I0Yg2mw4U96ZtEixQw7fVrYGLHieEc6+
tO1qowrrkbhhwXuM4QMOoVgCra58gjj0PdJ5ZA2NeaH8evrgOQI9ZZIgudBCV+8yZz1git8A515Q
HvMaDUkxFA1vilTL0qsGOiv07ZTX0xAxitb9sacsDKAju2OrFbkm61G/9+7SJrDMUv8gjiyyaO+p
fUkufu4paLNn9HcKG2sBCXSlRWXpCRGIfT3lfVp9S0CdkyuKuyEY5HDGutfU97mvCKuoonk54Vn+
+Smol34r8xcUbjut2PoY4di3bWmqAdnhp3W5zvEstm9zve5PpnbdhC2e7BIg1JlH6WU5VrKNtWGS
wquQLLKuXVvXfMfZWgqI+ctAJPrTyQaM2GSxE8ioIsC4PyzUS54Jn+4rsP19MeAsuuP8I/+da0Mk
4WHHJmMJk4ukRmkRLjhLrxawvxlNg+njPGKB/JSEaFxQlnKpKDwmpNjB28BE+TRcs8PXzYPaeuFq
0f1AXc8QJ5Fu+gjaHk9zxSqoSV+HkPNpf0oEWuMPPzq+XoZkTWFNHKIPVCSuBTSxOji1zxAIX/Xp
kXp+i5bAcRLnLj4ewuSRgZOalIyylYRR7biGcjyEsWlHCYl9FCJV32i+VRz88zYCC5km0CBizRKj
O5rICxI116MZnbsN3ZPOlSREOJofPf/+KNx6rA5hh8PmXGsvc7y6ASrcEM80vN4jhrhbgLo0qMjx
WsEQAtny5Gx6vCnd2sgRvh/25c9lgmgka5C6PcPwUIW7kPNogEUulJPb640Wv0uToRZPNMK6oIQU
xMUTXyOMDackpj76q7RbYBcLcGl9wC8xfrFirfohtKXYsP0tICOT/fM2HSC6cGeERDSIn2Uwktxy
x7LP++vvdIsQW+EPP0cPtt01EgODmTQQrkbDjxQeID1+VRF+ccjw77xE61xU+j/j4W6ynTgLSg3q
jU4BcWyy0Nn6xReSyD6AeSngfG13QK+ytaD77tFIB0C9dbf/Vb+hnErSIsKgYHHH9O73fn8Z/ISK
zApqkUDZdm17rkq1Sc7lM2+ZkurB/MTvIvlzO2G4TJRPafy5tt1fGvUy52ZnvQHRAN0XNWDVU7xl
rTKVSFFHdXiVCzsiVHFAA6FwnU+DKu+wQbCsfPtNVhajp6MwTXV3eZ9qYccUvDEh2beePg9NKIgc
BjypJ4++qJ+8OhFyjJWhd+tzHUGqgAswlV4hQiJ8cbzsCIRvViShbeH7+0wfKUwTas1i6+S/uTd7
Z1XeoYJQy8WaO6hgQ3ozczaenyA4DXBll+n1245PfOFMKN7IT2pHbjO/9vBBX6s7UgoHF9RgKiiX
VMWdCgLs5oZtoz+mvY4kutWOWwXY+yRqN8AtQ61Ry3cGW8/WuS+hIpEVP4fBivCRD7DfrXyNm6Rf
SKhSQDdoSAGxSrginIW74urL/TOLksSDlNaxlSD5R9x7zuQO8w5kcO9N+1jQdPKJL4re0s/aQ+FC
AO5qfnZUIrRYW5MWTmrFku9Ucf3cAkg4zINi6DdrIcWNPVGe7l3E7Zlz9bB3aAWLeOhSJaA86AH/
nampz5OSFfEc59nUEu0f0aECz+vVzE2HzW9XEJdxOZRsbVRcREce2NWIU8aHMQmBPJos+2KXXHwv
qRGQm3XPEFAINSmIGP3nwoILsnG8wGknQPLMHkNHVNLXpM0kD9Jl4Z0iy+O+sMxogVcp6qlW04Z+
pFy3pEANSuOW3Ks8xPy4zzc5ai+1L00JT7FS7QpaeMSAKLC7Rxe16CTXjnvb/cT/klcGDbUGuuWJ
V3+Weup3/t0p1Y0tydWRyJgGzIc1vgZHLXtOjADQI3Frz34/7JrEayYdSBqLoRsOabWKNc/GU8QK
xTHCBTKFSdVq27/5hFa4eaCo7dlIzlmjOJ5xPPN16gu2TjpkXyrmzgJsibXEm82uDxr9vRvUJa7i
oS+f2eT3YLAvGFKvu5LwcMh55sGQJpyIfLFbr4vj+nlUVV+7i3nhv81Dnb+Vi6eQVwVf+nBbO7iv
i5ZgfDP3HPjGwTJoYd8dp0RGrCdYDEsKpK0qyNYVk5CoZ25Tdmqm19p6VKqe+9+MSEHPvVcaQcjN
Rf4FT4tr2sViwaTWOQLiC8jWa1i4yuXqXsE64rOcEvtaGe2WRBIHK4hTDoDA29THvs8ji4dMEZm1
ty4ThOrfuQ3e6Eo9LkN+7b06se5qLs6ttzu3EmESWi5a49RpxnIdnF5hQ6hdGvmkLWMsWF3zWfll
5ZpfqsIdKAFpvmCMg09V1etplf4u/q6AMs/UssRyetAVwcOlzkoANGV4lHGFGVFBamZTE4rgSjId
ay/L/uGnVe4a+eRp4vUgh9ffmLuoRblNZ0qtVgjorwZKgLUdEml3uYjobXlooqV1mMu3xhIrp5zz
OyaFj+9LO4cPcm162zx4ckuhYD0f2WQTtXMjKfuNQmQ23tXWh6q1yyQZCV+4zwXCUVT15x6nqyIl
Pvz/XrpNUtZzUUkArdNXFSVxxzG42Zp+cPk5yHBW9Oiw3ZBBeK4pJhlXBS79eOravqyKEdRMwbj8
j6YrpuZ9bDnyc4EB8QVuN1x8UibAsmvAamzk/MrrgpS/qB0Szxq98FdyFr0rm+p4XiCgURMzjDU8
6tEpQNRoKIG62jCu0j2kBmyYuAnBhKwyUVVFqShxq0jDGHoeqKwpmfC49w2KupiZdAGl2Ew0LTBo
b1mQBV66j9tNSWClnnyBJGtVjqNQLAkqLcMNwQl6RMi4IvDPuR3Qqx2ZaIMf/mdG+ur3vfKYzhna
ihGoJ+3FyXt3ODzNx9cRhDJnq3t0NptICwQgpIU09WQIGguwPHI01Ur7UlftO8MkvI+H0Hp9JTgK
kq99l5ZY9/h7devSJ+r6JPLhuTRufzOkslGl6YvquN9WUTISsQLdqACY3HsaMiYahIkNR7ANcg4Y
BtC1IOH3SSAS0zTfam1x3P72kcZb7VF0hpLVwGqZoyhmTrABextAPokC0Z0Ob6UhQEfGtzjyl0ow
TYwcZV/YCTmO29w5DKwzqZzDwxdg+KX2h+0/6Av6Cp5DvfjofBmAYf6hGkj5/c5tDi5pXtFE1WVF
96DR7IACz/1OJPntDLORc8GdC59QZr+mWkUKQVX5IK6ryL+nlavYxKk1Wbo+F3EOW8iA70rWTQNH
0Mzh6FU3bF3FIjFK+JiHSs3HApmSYmPn29gAYy7jPspg1MF0Cfv6KEmlwvhOA9sJQnhJdkvNBBUw
Pv7kS3nT2lvW9JqfMjH9brmW3y4Lc91qs5eYVwJf2h7+3XwqIE53x0zrr/sjkYwyzYU2cWb30k08
fLwNPaEk8ZxYS9nJGujPE0VV7fbEwzbKbxl2YA5LkH0cYIlEn5fCslUmxIChNxclouwKD4CnP3Dy
ERjB0GIEDfpxSGJdGIIBunY9uSX1TysYWzVd7eHqC1NRxuRxOeDMcLn/qfXCVLeeLxf/5mooME8J
C0GgGmJNGr/SdmFjXVgF/IG/NEfZEUqeTNSHI4a9UH/T0rR+WNIoD4VSJtYsBBN3or+0Liys97uU
BxhZmW+01DE8jYLXf1eq/SU32Kq+9metCtbSsBs3mvnecOEKAb5sZ6GAwnIRz3okq2B7ORiwOqs/
OStQwl9xLEb8hxR2Nq/IbfccSB20XR/vBs/X+21tm55GSHoO3hAYrVajwGGdidl+rjmOs5nSRzMr
FO73xpWKRdVqVsznIfqSD2TEKcIKrO1SPq9BT6lZnBavmyTJaUy60flptby0bFAQw6NoOZOIlmoS
l6UWZixZJyi3HX4mgzDzm7gmXq+UvJgzqLvg38eZfehtYwWqcc3nRDKFKrstSGJh4PlA4X3nYnVi
erNtwVeRnNGgvXIe8uNvYA3/DZjo/N39G3O/2CqIYUVcYflgOiJhckGOD+Ze3nMRZYCbWZgYYNfG
vIwtO4qMZr/T3r9VHxepKErXZoLKtaHGYGd4XnhO5eQRK7kNWQC/C8rLBrvexbUa4qFuaRzEgW37
kqlnvJ8yt5zWQNVyo/lpHuiEA9ilFLyqW3fXlwsxMVZu1a48a7PnBQRv5ZKo73oQ2xVf5BstmQKI
DAbimmALJDi/18u+d8kgON4iGz7vq4fXnCE353B9yg2POoQmQFkdTfdMf8K42CVoXEhiVy8H4AmO
x4YOy/nmKTCG+ZRUhR+Mkdc7b+GVtRLBAkWyCRrPMgSf9g1NchnXx4y/iPMn59mHtWceRJMuDx9z
M0CIuhOx5rdMq0Z74mkXqIcKQRuf0EXSkEeCUN1how+bBropz/jUPyjHEusgQZcRXCMgVEYLHQJk
twMkkzacoRHrN5gn1V+evIbpjoFYlHfFPQEGexfBT35XM4Titugpp4j/It3T9JOv31EMsdnWwokQ
+0eDGeiB5ZmZ6A5YyHVj9QeXHG+RdL1+5j82s3+jzunlGMW/cfNerr8UknNS6lSsT/D9g/narUBg
4HRyg4/IoDgCUgOYrheLA9Bp1t1AKrh6JeIyMlQfzL2xmKJv4IgSH/vecWP6J5ZWjSOr44ARRhIW
mANybsH7XmW+y3uCpCvxwcB/4FuqRIFccNY/np/GFFxcW+CBLQjR6tHHKBjQlkYvp6Ev1YU+XBnV
IfVllpqTZmcALBwRGtzE5Zr07qGzu1BBBk1vF5jpAj0oS6BpUT4UT4P6DQsD5fzM/79cPC3BDo1O
QQDT6pyHQx5Su+72MnLta8fdDRsxi+jw70lUXELwX833QyKC7F3sRDxvHoMEr5f4Rn3Y5W/Ynmqq
CgNValUKVK/cSs2+QKL7f9HH1NbsjZoOE7woRC9Bw5o1tNj6QSTx+VsPFLSqgglC90JD6zXJphtx
wx9+OI25fA1mwehMmr4Z9nCSV12dw2u6sfKERAbNOTHTI1RQQXLeeGc/fAbkSwlyjxR67XrLOZ58
0snQoESCi/XXqUas+TOLZHUWaM+koi3f7rRj6CDcIaHApPZvnY0MNNNZ8asbebl649mcl/3BvOWr
3wRAOa1VzTxmLsQcGZpI4yqPi4Z1HTbu6P/slX+Mdu3fug3rvDdKZWpvqqujRr7c6/fmuv3iaMuP
pN6FD9m0owa0brLwJ7lxnLqUy1yLcO9a+Mhk2jhh+yU087z6IuCdeyQQyIiu1zhp3OsfAW3Yi6pq
bcRpEHI+ega8hnxcfK/pe+uBX+WCKmeRkW9Sl+u8xVuhYyeZMe30xUr/8jxrOzd64gQVOAZ1NBlG
dC0ieQyEDBSCwaCnBtzio2bDSDDmIB6PpHHbMM7I+Beq1pXpPZ4KET1CwV8sC9PSnztsmJRDuAKX
3ii/HOLEwHMaIR5gVrrJ0qL6yuy2gQ2efNr8WinbKkJgnKjm1R0EqeCkI4JpMI6b/SEx6dSk1skx
1Ny4BDDBQSX0sfnzpPV3R2f3mh1jppmRXO5eIwM/q2BuracctZThAYYIOWH4PfPTfallwBW5V/Nw
gvOZWyGJLWx6THBsgzPEADfn2543mlx2nHfnIMGQ+mVyv0fVNPihjMnkQ/vt6tpMSRhs3879syWW
9UFCqZ6tp8CpQVYe9MVJKTxVv1v6n8Fgz10peb9icHw06YSWo2uUQxRjASCTaUPQOe5/f0ESpWsl
Qw5Kc2e0yCvYo48cbSvE0jcEWJk3CcmsjNxHeJDwXlDMHRJTcdgV33zo7i/ZeuWHhozmNOqXfIvo
0LeGWhsVpGHAZN55IIWobmqtHRotPzVkstOvzZvEJwOBYbTKRUr35SdGxgnOHT9O0NgOZNcDZx6e
X5bI7tMuXG+khCPkMNEjxnQsPg3UBc5cgmkqXEbRP9Kzd4BiZYiQ3kVmfK7UToPBROi+c4J+WcGr
epJltktWuSrpk9Xz87F/dNaVPG69qq9YkhUSYQjj3h1DVO04y+twWd0L6KUHdHEyKgo0sogiM9Fz
dk+634sIueQsEwk8gXjyXUfqIcircErQFKllzKaFA3jUjixKj71+bK+fhqnhf6ef4A2Pco2cND/w
H8aF5WW66pnCkDe5mFKTfH7f2yGddeRhdzLgzongRi2F9Bi/nAdOfKuT53XCNQEyz1U1JG4Xa2fI
20odgSLvXPKdpXNVF9PkivQJ8v92jjB+cH0UHuziJySsmvNaj9I6DfL5d7Z8JP0STx/PtUr7Iu4j
dulO1pWWnZSLl06NDwOgM8VoSO9x/pGSqah9v7xtqGFoa+qwcGkeJcD6kBqqf/0zQyQ4hMIemi5G
6AKDvHmN+9rKOmu7RinC6yTWL+PPjE6Iaw2bFTAUB58sHNe5V9klNYWb2Sn4qji6JuS7zTOF9Jnz
kiss8Hf5Ax55uzaHoUuN5sPS/mIl26ivG0t22UNWZVXBtP1iEddKkzHB57YKI3QBttfZKFEGl6MB
R3kfabQSaQsvH8FYZZ/DxDQugXpM6T1wsSA/LkQjtIZ4MzgxFu85wF09TckbPk9a+AmAaHA+qafy
dWSwAUVOKs9g1MOiqax3RXRPXiJKOI+PIJYUwAI5zo60WStKDb3ziP4rPZiAsjpyBx20jyBfNwFa
jaLSqb1n8Zc2zDcRSGt8qPq8r3vcCEk+EgiCEvgiuq3Hw2jxCZ/nWlgFH+OviO/YZ0uqIOVU9th9
enXLFvZ/IxhMhssIdy3NH5SQr9yEaJlZMw7qw2clXKh0+lsDLzC5y7T5DZWafjhhRrYmGvatYC5x
QPbsBXW2ff5DmL4IG8q7BlndAAgTcTSaJzW1vf45qPHas2QLoJDXdR18SjtnOWDxWu5AKMcj7NE8
GyzSB30rs/mod8sRNi8WNr0FvIOsstpuAZCc94vUGV6hWgYkaD/N6ZTczkGYKyzQA/5R2BhS2E/z
0CRZxarHhBsn8Zt+8X+aCSlY2UiMBpFPfPAvyAYedmmgkajV2bVDKFl6BIePvdNNx8CpPKDB2RAO
sogCH5gZd2A3NOo4esEWR9DWi9kIOr9ezQJSa1XAwoEjVjqJW01nnFwH0S5hX2oxwkm4y1vZ8Q/J
85A3smCmP9B+/1DtZTElKWfYrf8nHv5fiKDWct532JyFkRPWnUmghYqz7YNK0mLLfuXoNf8OlrsP
JYIPkYuU//OxH1gD5ocyI3U+wim6K6qjei3rzRISELZay6qdgnb0JugxCimUZWitYm05AMNvlUM9
qi1LuETtcaK95GmmwmddDsvhkjL19ctks39c7KOf91P+gm2hZX5yLDGixVzRUb+nmtbp1ie3oCRl
D/oRwSs0E8rpANrbRO/xkEcTTpPosyCVEezvKY/+U1bIrepansiyLcR4IhY0NhQUvhExFxSSXO8+
iViORB8IKJRd6kHPY8yVa12OsRWbK8p+ttIawq8ceO5pP1WsKcOUtDkgmY2TaXLS7CUqwji7jRFS
LjCZAVlqVRF+dTdmRzxT3bxttmN62eePO81j3LPPYIzyqYhdZO6VkeTcEtTZuE9OxrMGoBj2XnYe
wtXKtNAaSnOZT/aI81FQegCKOXGIl7PT4o7MoZD2G/cY7qdmpTngJeVowQmc/Hm85M8J0I+yvpUd
mWa3KDhGlNVLNSC4s4IceffWan0feiMrcZrblasoUEKcRSWuctvQllfbCk/6o4MZjStuIuErRjU6
legrqJr16bGo8oL1vQRDvvIT8/q31KxtjzcvSKv0p74ZX8SBHp6D8qxdpJp73GxgLrCbtmDjAQhv
KfJCHQ1TFEvJWS6fzN8W5Doqvdf0QGdkKnDxqaphcNJeFKNAc146SZvWSxnglb2ww0TAoQsl+Sra
yT8uHoZnzLESKv9Nwc85JC/c73O5OBgGxYj1qcBuaHIZ95Mdr8hcSvR77FksQkthgb2EaoZf2jH8
IPKYdDTpaXmfs2hryRBfd9QsjLPZXNVeyabWNpZx+q9FU59msTjHDHfDL8ad/y1DJITr6Gjr5dEq
1rX+tGq7LapMyLhjxN2K+r7I+3J3mJscy1AG/taG0HmDcVSdYM650HGRDTV2mqfB0+vMlbH5N9K4
78xXgVNyvyIGpKdx41/G0hE6j71S48ZUFs5VFgYRl/2iNQmkWTiehka5f/whGoSnGtWDnfRqLTNx
p1FJF2x+W8Ektff0VHnrLRBd56LZFBVjaLcFEM+kiPNqja6ikSWhHcoCY85i6KTZAPfdr/Kyqa9c
XMi25IM5xvll4CAw6HkCAGQjygAVhklMAcoZONeqInyU18KsUUOOMylXeIlRUmRq4733x04K0rB1
+le3RHajG9DXJATFEPm1AGap+vrf3h9PaEXCtqKd7vjpvt/ngQqfConiD2djb+/sdLKBhC7zVhpL
SOG3n2T4wnxxZsoznKUEyREFzP0HgBzLaPRzjY39SvZF0LFDXK/peiPtJeHhsEF7A0Th5YBZosD9
pufgiIDFsrOrWlOjuzigHb/uPSOfgAGbJe4kk+pZMlJNsi0TLxpBMrjYlIbAWvqgFCFdENfPOjNB
23TPjdJUUp939Y1H0cMRlbcjENWma8ogQnaatJc2aqbrFr+pbz2xhBP1ocg04Llvg1n1C+WhLk9T
xnYql8Z5+GfHNryF/Te2PITOA+uAOfTS8u9iKeYPXJx6UfDb2DlU84MTC1C1MZOGtMmEMGBH8/rI
Hb/AuQQ35uFbxmKegwcjtRwtzg1WAPr4i4AebqeCq0Ta9yCHSD0pvUBlNJjuRxa7+9zoupoG3U0G
fStDvzai66LaM3ziUpuqyZS+n9emW9SIpkDiAOVnyEjP4mgC7vD3t5/2vPs1TuaMBPXbKFgq+FwZ
FMPO9f0odgSG12UM/OoqrsTr41aRliI/GRw1FP0rEzXvrgxUKppt1/2OCOJMJIytU+MCbcG5Ed4N
Rb2/SRR+5Qmym4v5dpvc4E6ns2Mq5S41g8aeM6XHa3qmbxVpe1Zd6DbypDUJQnu+ZmIocg+b/3wa
wINOdkVHCOHbf5grgZO5f5N5EJ5L5Kb9rJhdu9qU/GjTulRMNaZJ3u+q5Kmhuhqt5AQYvGXq64vl
39Pdm+6PumuyWNXyKvlk7ifpjC2RXBtYDn4Uy7WM/cQCLxSKjli/qkMjbGiQtEK/YtCF1+7e3uM3
47fvFvBFDxtED4JFC+i5bra3bf7hX+7l1SwoVspgohoTJZbB55a2b9SMCrKECGmR422UPX3gHI3X
7mQRNGsKHUx4sbuxF3dXrGMed67w0eX+NmLLr/YMbhU1GEFHjOPOKdVmoSk8arXepWq+38c+e/+C
wb412VrMSOk1vT0ddqYaxNQmKhqvx2ciXXus+o4MU4QatyTGaC0pbPIaNL4FlezaS+Tjn4J5qNnA
0Zqq3AnfpkMUWd+qb25VvLQfbOiG1MLbOlH3sTaxhO+av707Rv1aRa/tKKQxhfqhEyp24qmQQlY7
xj/PhnCMLtVTuAa5QJJ1zX+Y79u0IWu+BSyXeJkT8rQifXt9rCsjQnUyW89Y0n9lEdlZfcd9laPi
dlPLg0eNS08SrU5ZINMqWPNTB/myPsYbQuNetKchv7OOa36sqhkuHyP8sTg+GOJa2cmLmGzkB5je
LbosB347sS7/rxk/znZLOoRtiuzHQPTHs+gm/KhG9BvAmL940UioW/IIAPIEcrfkTqD+X85zQiWD
VFUvbdi5/JqzZfOBVr0+ZHkYqoc+SooSigCdGSA/3GFMeouI4uQt3+VIU7ZJz48LauJsQlTMLVjZ
mIyyFRpLGHycBkj/IDxKTVR0G6lJt2lWcufvZhzhmTbg0tCne2mLWlhT16RmWdQNQSphiPDpWM9B
NvdXTdY8rsgDV25//nT94wHbGEyTpJpi84dU7cE0ZrGDpm9s9cXS+W0xwPPVXe0wu91zBfekmzQJ
oFSl0DHOi1mgv5uk/ue7h4bXVonK/Y3FUSE/bZTz5+Kyyl6B/WTcOj5MDBpu7rIj+sA4OhzsdLmG
pXQrmHSaSsWHOjTInGsSXVgYPsYVxZqAKrCWCC6sxlCWHGr6cwqVHK2rvyTRsYJDfkq1k5qDcBP5
9NHr6O7Qsj5zAj+XS05cvOrsvaS5euvuTIej/1Msv8viBxDjduJedLcyAXQqs+0E7ebgx1HTpXdd
u9dfmwWzcjQeV9vxwh8IPFkMujT3E/vQDtTYRcoChjDK4B/MXXcusotNtKYqrNgKPxNhmIQDBa3+
DaQGsEsbHn5332BN0f4l4udJSfrjCixNskACloX7Y0IgELImokaXAkfzxxFKIsMetLYkjACfkfOP
N8xuK2EOj9hckXJDrnJNNB6oESgaNbyrQRu4Y6/hE4LzbKyBttct8Y5ObwBy5p2lpvfoUx6D6Bh2
PqoqaVjyeCd9pCnjNhQHkdo2HiIBryURziAipv0BM3jp20v0tq1l6vl2H0j0Pqf4Eam5px72eohe
M4y8DOPQud7gd+q9AIyHYRySVZdJcvn7wZfLd166hk6abnfbL/y6v43hzusoSjpkEbJjtstB19Qa
Rbgd52nZPfqg+R+2Q7WBblmHOren0ibiH2anHarztYuuEsQN+5K2kDYxqBy6M9JUqPRxyhEwNkhd
zk4UPWY+/ZpyKo8bjN3I5M33W5KxifQjMUlb7SdYBR7LxEboPcFUWI/X0r7yRjSoTmYe9adbFH1A
sG8aVL5IdUCihWNgANpjG9awNPMV8Br8ivgJWwSwIYrmiDV73wjbvDr6d/rMLJzu1Z1ETYhPQUX6
ouuQdKtD5sqIC8LIMWazPPA49HmZS+mWAEtgNEXHQzK5UgrJ6yh2fyILEKOtPJdpF9CjpGxn8zzf
J+wkgst3JE20aZCWOpdN9IZ96caTym8rVMa+m6EU1dmZCJ4VMeCtrItPmvg8larhHWpOIjL75MER
fJkeqkGI1wPm9wVA6bN7TMcHFQbWLUl+MWBC4GCtf4Swgric+9KxCHo/VNZJRAn2b09pqhMo+E3i
nj9T03WIjA7boFpNjm7kbVmv7EJ/6Xdmzb6Hxr5/oLzZr71ccCKDXBhbKlElqhRAePdk9/aiG1Zl
VUvZ2RiWmsvj79sKCO0xH3fBcVlZZNiapKD9WBRhEUZC/pGgzDoj+ZuvVIKySJrgnxaTsW31sVpl
j+U6DU9YkVapAS7w4l6IY+cL71AmVN3HbBZeM7l8VH5f16vPIidtIGQlJVlRVkqfRZv84B2FsWZc
+Nzq8SyWZsi/p3pZncMlBi61amg39RFQIUNZVQSKppEFatuBZ204K1oeMNgwV8G2DltiSMW3o/Jl
w7QfyT18DBydR9LrbzaaQmloFk64yKXkyOVRHQJ9+zA4ud7Dm5HxqYpTjKvZduu0zoG03+pwe9x2
MG4vNVLiWQzo6YETEiDGq+dBnJpnwTfd7kECiCJeApSDstBKTXxzJiCP0C6gm6ckiZQD1kKjg9pQ
ELhdiF+MeqVlS8LJ1/A1zNoBsadOPKrL5CmfASitm/jwstN2u4xsG+mWOvEAFjPNxTWC+EGGYxnq
3wxKBqvf+irQ5TNkiK7PZqaIUQ1dBXyeddPHBs35QBEk0krEK9+3iaf3AM9+YaRySoyaOByk/CkU
ayiU3J0G0lqU+/uEcZGDE2mESYyH8OmwkJl26LjicRU2Jn6ZW/268u0v8kqtP1aggGdNEP5sGOmg
EdWWKufwFEYgPdKAxFOh5ssJyIshQWCV5NJcpaHtIIxYUv0dEVmkjmMslHIESAZlmFZ3levGSOUv
naGNvLmh0Uy9HghLi/O46H8Gv2OJo4JfAbvmx+8s8Ff1bUNPJruTh6e8LzNuttIukwlmZTQaXxH+
O0SSyiNw2NrE5wnNZkyAkEC7ZT2O3prvWlQ8oldoInighCVde3xJQc2360doYTMWDClfbBjMLJDf
RA5t4F2w4FEXnr0LmsFRZewv8CiPO4Vq7QnVkZVTA1izZhugbhcAQ5ezSWVA1f/i4Le1IjdVap5l
4dWih76amAHlKW7O8xRiWNN7HeKKBeFBJ8FSAQHTBCEg2OVUaM8cY7K34+QyWI+p/sao5EH4ZWDB
34lQtnMQ4DPmxuOC+oaZXjLvYxZbJOdQoUE4+eJvPlo+91NaJppL+Aoedree3uHgGmWZVOyZcYX4
h9Xa6Z9ucki4brpVJlpS8ZJ/5uLj8tDA1l4MjlWlA23R2kWWgV4D38gE6A3N8eNtfVZd/9CHeq6+
59gEg1kKzI7qnYs3jZuB5u/A70cuPoaNHP6i4QBqBbxoX9Dpq7lwFVJQNGWZknSi03qJk5SXorLA
y8BZCjcx8SWfRyXxcQ0E5wK1FExZyecKRSkSdyzIbGSiW3kpj4w20T4fBNlRMTB2DLudkxdcIe6+
VuDP5DgnyRNqkxFgWKAEPwQyLUUaHaTkJjdSvTLRwFTNoqHMLIPsE8c0rQnHubrpbUE4jXz4fz2y
j5Jd57Ke3YiDlrx/iJTEY/uwex2sqG/zQRHzS2ATCadL+/hbNC7Tz6Ckhglzyy/7X8GiEIl+FqU4
hsSWLhs0prId+hPSQvoT+idBUwVVwpRn9HXFliWUIM5wXNav5JZfZMeZ7Bk/kiNJbNYrXdFDguz5
R+NRnVA6exxCOv5VUp7QnP4OI+9phcBPZ+ZpoJwjzEgliRBn8dJS3wJRvHl9FDozorHlg1Yv3v67
Qp4H/9Kdch5u90w1DcbxagY+vcw2Ki6yzvt/darEPdgZ1AuXLoU78QdYgr6rrzv1KV85eEhvCLBm
u+ED1MQMP8O7mg5S2Iwp/VLDX+gwu/YeNZahaB0rWA/AT+S2BkcqXIlbtuOk9Qsk/fGG38v4OAHE
qRp8zHWaJ97K4V3huT9gcSvoJHCzEFZ3Bx8jp6uvXtlSBPaGytg3USeYTKPTVZ5bWO4lBlwGOmU6
z1c+LcUj9AT6deoiQdvycmMq0bJH9b817VKO68G3C1B4LqlpCEjpavwKDllattnKqEoxDdU+hXYI
kS4uIs5VDXHd2++W7OvlUEAz6BY9I19yEf3btW0RJd/MM6/g0vvD3C0eC2d2kgzX6K031x/0UaBj
7Duhw63DO6XIl722Sc7nuootob9JQy0rDma6N9vXHxSK9A1H2JBgMIskEJEFaNHZmzje0YiTGgj1
EpsbooLv2sl+h3k/0hqEzeYdiFMdMbeZh//P9Bj7dcOlHfrc/eiTKXebNkOnynyiKOFSSN4Bm8Cc
zP3XI4f9rXrKiO98hD/lI0fJleDTOZi2mT96OplXzTGaFjFEzrQc/itnFtBvSqATdQ0YJZQy0GfR
4BLs5sPwb+JMK2Z+bTZFMhvM4I0utb9004KBCF1h5a9YJ6i8UkyJYa+50vY6BpSGGVifCi3f0mg4
AIr6cUGDegNS2EwHiPyEZr5uu//3DzioY7desHc8RopyFY1IlkNekXV+hH+0ww4PhaYPAKz55rLo
hRBBjKcKG/dwH5Iy1eFU3GnGyLOtLvCUeUtXxjleiofEi23pvLSiJcH+24rjMrx+ozafVV1xl2+C
p/qi06CnMGi5v71pAVv/Fr11SmpoNK8DxezAUNo19tddJch04UAyOXCHNowyZS0nTFtYArp3+f5M
xRkp9nYxv1CesIHXkQwyIecrvH6fREkoO3txn6Fld1NK3UPoK8/bu9QhEJ8a6JLUsnMunrNXm6qz
NFOB+vvZ0P4A0zV4MCjnV8IKAUEfvqZHMFL2q/kzBS8Vy8YDo3HUfx5CZpWXSq5/+duunlvVlZRV
zQOflxvbXkQRWEd2HvODs5UuY8fhJsoWQaO3HNFIZSNp0EjUxXbdbQ9Qsi6cuOK7WVcOv3YNW/bf
sCRo5/l2c+NkvVGylmO9Ivgf9JrdaqQqXauP5EtXZKYuQ2t3Iq4er4X0ayOJyg73Xe5cyIQep3Bo
rRGDMdkJAaulyRt7p2C6XB4PmkaA3fLgDu0U8yoFNLVylTfXWTQzej5qAUursHS+kOnjcGVgRq+0
1KTQbbcx2YrHOtMy/XnvqOr+8+Gxv2o9Y0BQJct9rgRycB0TbGqikR9ukCRfZ0t+PsZAIHrnl1+e
8jKfYCiqFVkOgoQUjy94zIK9DxNy6JrzfaWlsEfV1ZU+mgEklxpT/BVn+y8rNQB+K0GDMtjW7Wy6
P5BPiHlUi3f+fjlXk9U8IDJ9SyARMpkJk6QIR+PuxmrcUSLZu84rdTlZrD0bGD5UOh7R8OvFWpb8
LqMUeHi4nvt7PPI2Og49/jGfgpHEASbKaYlO19lz7GnXOuDVZz1RqDvjhG5AKnyvoTgkOTQAv/Pg
U+vfNlF2ZMohrxZzv3ODUXmY9PNe76P1z/jsLREkAXyEs5ic9SbHhq++DHxClFVWiZv2qIEIh9iZ
pWk9IwD5lBUXWlDGhIzW60wJcPeQdDsAbslEXAcJ69i/N+OnRYzwmf00Cd9jmikkDf+btfQ41huT
22ml3GpOTM4z6vmedbU974wdXBe5RNxBH+iCfhLXKSHXy7Z/vSOHnmkimDpLha2HaqIxgGsgGaJm
MUXvLV8D4MHxIyI4O9KCMfE9Hl2r1tzBJWdXmZk2OAMkP6TbwTeMh5NXP9efVrTZAK3cZJuH1WWR
TbzQ5d/IQaFuqlOtOgc7mSNyNIeXh1Hr/BuHzWRBFfNTwuKN3H4N18rGdMHN3wnOOWJ0MRd4uveM
fNKyRfFMW3XgR/z7eCE071MnNMGvDd4THeSK0mBXLer3pSXzP/8OJEPNXua730v/xQS27eKasyrb
t80G2RSzcrjolC9zvPVF6yUqv9VbMCFOrqeTAUgKNLR5H46FJLEHQh0xeAZM1BD8TlPw93hpZWY6
KjEoDV5LTbJWhl3LdLaqcaItnsLCAEWAyABqpP8wg6lWLUgkZlUJcaOiqCXb0TpzX8QKU7aYlPIR
Q0SJR0NMZCpd5pfS9y+vVmGdAtHCQ4Q/jRxdQC42+mhOO0Dn3KczcsjTjo0qUn0tnnKDnf5Ir+8T
5hqqqsCqftFMIvCHKIyngsBj0IdN2F77NlZ2fVSRSlvnyX0lWjMpRcPsBbn2ptdJ6rH5OeBawBSr
a+v30PzKGSKXMIs5fACCdXfd/enNLq9Ks3EdH8EEIwCwC6GXJnSyimhZt2H8E39GeV3ZBV4I/yQw
XFPVCh7I+9Q+GWs4mI/Mr9w7xMb7wjKPIiHHYOZRWxB29C3vE1ytakvj1IFueXWB1tDcCm5dDzss
qvJJMpB/eVsSzeTunr8xNCTZAs3xEAg0D7TVOd/bXjeIfHXP3yZU40NrKcIno/hxT7G/X+AcPT8H
SSfEQoQim4kD5mIbw6KqGjI5cBHKPaOUsQ85cNVDSzvk6So0elnGNK67e/KYiZBJxV2qZI7Q0QiR
2HbKr8o0NTEyiK1ql79L1LsXY9Q7Y/NggXUOg3fU6v86Gul7upe5xjqkZgF3LXt7AjiTdIMawfc1
lMZM7dznJHze0xe0aY16+mZLfHdneQsak51g5GAqYkAhJoNE0pS/VoctNh8pENEeJZEcTRDZiR7w
bOX8hbNvbs5q+I/PYMJT34C9kweKidCUbZ+dr8p8+Tcpi642m82x9CX4uma/uJIfuolOWSmGBrft
jixiU040KPz2tb5fmB6hcUaZ5PCYs5pqnYK2rvFyLmSMPzcAGlFGUotKL+d6pD2yEZPsGe172KJ0
C7iwi7lmReTRHAUO1vTTyH/fS7HuvgwHV+tUTHi9nlB3a3uPlwUvbcPq4+DsMOeCT/WRCpdOIB1J
SwLDt1kA+09vdp8uM2ohG2E3Y8ao7FKthvVU43VfSCuW4vFhq06kin1Gyz8yzNK7MdsL92aMqsSF
ljZ9V2EVfTyMj9i6bwMHrpTmS86okxKbdqdyAfcELv1d5g24x3DKwSDPCyuzs5h3OdO28bKQN9it
j4RGLRxLU+abepff/JgQNtt4Q1SreCT1e1sCPc2UBhBQGJRj2S1R5h85XCSYpES8i8LANaMT8gcQ
uyZeI7wyuDuP+Dn84+kGVD3kYnCalaCHEkjI92DW9CFK79kxZbOop2Gy3lxutHAmOgTFlJeno3pl
+cCNiTRmm3QLjOv7De+lbZJkuV7wFJ+XmSgPGXOYdocVxxM2oHgzImPQPy/aKGfISsxoohYKqWXQ
PN596cBHDY/S/0m5tqChcyWrrklklOQKdWuDXAAFibUCuB2LgjwVKtBgSHNKczvqDk5QCMbdcV04
ZOH/c+EKjMhP71OAcn1diY67ZhU4myhWEJczfPSCWgJUR/UkZS5xKzzNOpzZp4Gg2jPX0ODEzsyg
0CXfk2SWH8UelhvTGU2l3ofCrR2bfvhxexkHZdqYIKuMm+e4LMTfpFN4nsrO2RZAtSDA3M8DunuJ
JYaG59Hw1XAuwBtYsCe7VZS5yCSNk307btrGxUU1U6/PFoGQRinW/iCgnc5LdEE7Z4ltgHIv9njc
JxbHqspkknlzi8Nnzj6Ms2rmGIcTxjxrbtG5GY1+HME1xyz7OEWkpNBTPuvPVXvJebbboAAYppX1
EYPniv5fSAbZK+bM+XhMb3Dn0t0M3i/GckdRFVOJpGzk7aL2LKo+FV0/SjlkOKptWpFTkWz41jog
pwmWr0YG7nR7gLPfpA5QnBqYryKSYwFntF845zi2d2bMg+X5TqDv5KW8QDnvHEs1TEESRiX3uh/e
l9kIVYh3JyPHu7N2WQunum+pQ2PSFrAz+F8eoe3nVk1mpIEqp6Tk3XeXgIZ+G6hziDVox2DcSsKN
S/r5Kb7lCdLvZqQTsdnGJlF2plQczvo+i5AsxkRxQNSzXp0Gscny7fHejc5jMa69+Smlw70QZQJR
Jrn4Pouih6R8Cr8dRHMLVoJzx5/fxxmJU8ES/Xt5FvfelJ2IMxClTTzCyxqK8eH+Lr7uHScyUtXb
nSslatUZ2zbXxs1oTmu7I62EKNChf/BufFLcSrl2bEuyf4IsUoLRqiPTc6isQJaJySWciy+xsTs2
kAoCNHXvAUX9m0D4ASkUqt5hYSEh5SM6SFLOaRjhJaWxz7ltfSx6RSjfkO9W+WTlurdTklFGzZpC
g/q+wJiTH+rgWRaG7IrKKqNY/aTHmNNOqDfeXqgJBO5XtEqc2VDZPRRsZ35/ipI1lMZcTcbZWpFM
pOadYsigBuoad4SfsTBSAhbbimZGaqJm1cfxjh4Fr8H3uZFA8lvuDoSmSTSbIUE0XRu2v1uQ7MeT
C/cuzQ7YLN/zLvbU43rCvSKmdQ5ER0wCM5ZrkS5WnRIztc5HxATQMFUM9KWETX9QkanYJ2ORcoL4
Uk8HW/ZhMD7Dw4djhZYT+8po4J+jTa+ZRcWN35J4EJh8VJA2EG1GfXMjueRlymtq7dZu3OIrTarl
Yezj4Xo4dTUAuyWKARWwPrK8DPY8wYhyIxWZAJhEr81UYWYUIv7ci6Wy8u4vQlLuOt76XQJ/BmEb
dBRkEi9AfVJTI/e1PIJu8jlnyQ5OkTMGPficriOk/8fNbRYnv23F0+pBrXEZe3SvBqhmHnDaSnZf
CSNVsc/7DJRCH3uBER7HpmEWH84N7/uBL/O88w9Jo6HFC4bjF60sIDkHxpmEvjz+LDi5kSwgBPgJ
64h+avUN7ZCsPEu3M17CiJz9GmUnykEeMSveWkPXLftcpb9ZXKuNrCMQ9JLBb7eWjK2Y06uihPfh
poDPbCEnEk+lWefE4xaOCFY8PlHtc7rF/5oEYKJbyJQ2KTX9rbEplyWTFgwKL/wC107gEqvE3+2s
UTF2Gu6Zi8PWSsKcfOyVEQqTEtnroxx/wCf97NOMR3UOS2CBwjWXbD6B0Wd1G4pVEoRU6fd9lp53
LNs6FZH0k+MFdLtrTk0NArHxB+H8JOqvE9qbMRWXhQDrmBTlH0FcshSfB3tbOyTCGFU/bGZP17jZ
sDjJtONzE7bzAAbCVR1uCWvIyQSwQH/QiAy+pcW289Wm8vpW7OrxtkHUCWPAv5HjSlGomgOOJbaW
jfioJvywgSeqZsohx74zpXftzExK/bPfgx/P+0bZPZefBTqy0LmFeMh3dI60bOkNqPRRPN4rUDmw
oC+rAYLQb+hsEmu6VkTbR5TMIHdn/Ep4YOHkx81Y5C4QFu0w5XCrHEG+MvzmIYSCCmfezqp7+55k
tBWTxuoamOm6zddxbu2K8VNXEg4b+2tn82YZu5wthAs3XR65kJMxXBHn2tuRn6WF7aFfGSB+wQbd
TZJiy50H6C2p+EqWDfeV1FhSvUr3QvZZXMafEjghPcL7wirQQd2DsN+wo9V8hHuzQSoQ2lMvIwlv
5LRyZBGX+CiDiD6HZ8XqjZumKz/MWWTbzM3XyPlq/t24/pseOymoU4WKbViqkoNlu9Ljk+uEfRsl
b0YtLMMC8k3lSuAdTVtlG05d9DDjMO3ZSW2hRIquoYXuHdhKxA3KuE07/UnfjE0gmhgAaGcHtkmK
CvpoptbBhVJ6Qjt8M0I0CcZHRnohw5vbHbX64KvcSnLqVNXVAM4zCO3Z6C2GzXgrEY82AGT17LTI
SgPOACoaEU6Wd45Ny2AG29vWDQynBT4RbE250gZRyhcoS/Lsd8AbyOHly0dmOpjWXCM88CImBPXJ
gbmkVOa3ETepS5X2UJJSGtvyVVYg9YCjTd3XGeoCn/Psxav++RIBBBACwsAiqvRDpZ/ujYye1Oea
37yr9xZjR8YAPfviUkZ344wARFXbghBfVk1WgVvUXkA0iAgcqbsjX3zQIgc4E2mO5iG/kDCjnLiw
Zxfn3Vrvvx/4es510Zp2uZhSOzHcJy1KJPJGTSuD9rEdgE+CWVcBELqDPCIb8J++rhWKY9TZ+3lc
r32YDjrjQ5MtwQk44MGYsUF050pjXzf+FIO/L7UuYjWJ7dbWEg+Ze8l+2zY5WnvWEalLdJ7jE6wg
ZdsepHdBVW8pj1QLU/S6xZlizBeuKK/0CoCpjF+CGP+bV9Myu3OK0xK2DkXt9EUlhzyesyJ/Vg5+
YAB29FYQLyKDGrNJE2h2z12p1WWLRPHewC9VK+Hh3AU1ScpULyTuqBTvJ+MXjSrD3YT17lc6yU71
/FWgnEx0YHipt0D9CzEfCyXoSpscEQjIYk1L0vY6B0NbyX82ScsUIINngPL8qJcUQDkC5j1dXNBm
qa7tir/qqTWYpgEmvpwZ19xOmgQ44wR/smfEdhXhBV32g6g5PVI880S4oS6vRaRVMKAj/ZbuWjNW
DrP0vh+nXCZninkq/gaVqHuq+NbUZZPzya9f0SPuHU0POFwUxstwlU/+vS4bIHXNJ1nWce4DkEJb
QbS1mLjp4VS18z4xW0C2a/DnR7NxuHnRaRF0GS6IJs1PA5wvvaL63qy7njlYfpO3t+n8GuwLj8ph
OO8L7lotCymeZhQX5A5JzmAtJwk6RG22vGvLgkuMWNx2mGTaXJEjvBpBLcKJSvFKxIZXsnl0EDmy
RVLg3GSaNUH3AR7QVElSLUwzWW+Bd4OYDbrhJK5hOqOheu5CxviYRx3fkunwQc3nfnFS7FvDoQxv
EPku1i77Cjwov50ysEXe7sHGo2TLbzQyJPQP+CthxoSuNgXnUbQzzTJxGP1zAaaALc5VLBcAlKEE
VKB0z/LAAU65u9YrHajdbopZzSotH75QMTiSJaKuWIPRKlXOyJ6c3VCUtt5J5Eqb68Zk7T9Mk7d6
ajRMQg1oqs0oLzBwVZQ6ehaabNe6ZcuDFQf653VewChsZ0BA7yyUp2WFabdHHIGiEXySChSFE88g
qtPWw2mPjxgNfies5w3+u5IgxsjjkVJaccWR4SrGZ5jAMACqDUqwmGKrsGJRZQbuJebP/GaWepeh
Gxfr6fXzl9tTPhdePkmdQ6QVDppIstqJX8fMgnALBDiMkuouiXmMkD7fBF11XjPOJc28FU+fq1N1
CdA8k7L5/S8kqmKv9tcNqUHPx5n6QG3siRaT4uL5hWFxf4wEq7rxCpjWNGF9B6BMAvk4Uc8PMJMI
iFtzhtCcdW1ZkbF4gGZOQUEdPMZ2hTpFoy0iIx9GjPp6H2KLJz/IQOs3YUUaugbahRzSl97LQSuU
Y1gMHwQ1gBNNUrNTB3tFdCDNP5xcoSa069tdf99NJRH8mcejy7dzdaeqNdYeqDHxqi5s/8zg2RBH
j57hwdATnvbeK7LXu02HT2jix+hh2KnqJs7XjMwTB/lNpi0rXgbNZi6b+Miwqt6LzLOIkSE+3tZZ
vvHwPcdEind2iKU9r938T2HU0qP0R+lM9pb9EiSg3qXXQuvOtJMRB080LifBd/b8VyPPS02WOjeb
3ucZtcK52PmD+HoPxR0H11i2NMjie4ZIHaHinByPGNCnJls9g1TMACMv4asxD+df25QLfOwlVjpR
wKTHje/d3YPIA4WQ2pzB617A6jQlHoBjAgOG3ApCIrTl23zSEghwGSq9exBoBB5ZB4gUJxD9miXg
vEWGCtaVl5AECHwvBuR+GbVuiVO8pFsjblC4PyV10Nwx5mUSHSaWp5CWDhxvEOX2NfUvX7Ept7Kq
t0+eYCqZRvEoyQoV9n2pj0IxN9mpPMZHXE2CgVIbn/SmeR33S3qts8uIo4T2JzJw6bozvrgZiAZ0
PZLqazeSDwk2dZHXaiDnlzNVeycwZagFb8jGrdrkqnjNBE318v1kJpofOp1t0YjZUjzx7GNGRdI8
/yrbWwkh8shxyXml5Pg4Knpuf33Ft7WK8br2fyHkSsOL08RwloRps2U5rXrFqA4f3bITSFgZKjxg
ymMBJX/g/9anORv09czP/lm1XFaCtUJnXtX9YKd9iEpkwUnsm8s8XNFCfHcn0WS6/HaL7sYqi8DM
pyEwUO+dyxjClq8c95kTOjNNyZpy9sAzD/EEdpDh+W1elU1lGEDlknLQ7FZWmtAYs/KdtuJC3PA9
aWmK4/ja6TZXhdasjqiQDoiOCPSRs4GIgAPPSxSTFaADnyEnF/BDRCWeyAgr2uridXivxZDdmVoc
nLeMqtSs0Ga6NHJWz2asjYRzOOM0uVpZtBbyU4uE2LYLxP4YK203P/PZG6B+3adXDVWusN9qXHvq
d8dFYy4iTe85MByPPViwHgNypsIRgtkVH5IYmQjkruDesPQrrMlSc767+OvNR3KXKh05zn5D7OFN
AkxZznM2oLEfikF9Vs3I54ckpKRts3eucCEsWu0yn9LdTVIkGeYyJH8TbazM0ScoMSgnNSVUuls4
n1lN9fJA522cfuSoHo8ng4lkAa85L/nsU7XV2+1hRmHXWVavEZBWwobrmubikjJ5dDkdQMLoVdXp
vffvU3w3J9VUTgCn8UHy8cWwEuUSz7thNjS14XjY0WZTxqBbyzBaqTiOpWhfnVhfuSBRdoLTRvG+
H2dRHn1w7p5u/tr4D7XYCEIiV4q3DjIFgo7ynTSq2CASGl2Uert+xiO/mWb8oPjox1IuI2/DfWmi
ldPARcdrnus6FE9ooCpp5JCMaISTr2NkM2vVXj5orCa6dj1bzxWyExZtk8VIo8VFGMQd8PxaA/8S
x76hTiqaby3fcujRIUfizc1l+kqbFSvz5ZMjt9ukiDxJmz9+CbHQGKOcexxYItdu5R8dutD0IwpU
8giUYa9YFB54hRvO1rPyzhVkXD9YywdWtirDBpXiAgySAqBb1p9//ZTMAafderQjxGoNwq+uyqYd
wCY26SgbwowrozWaJTqjCCezXmY70dSsLQM+Fa3UQ/yAeYRlBE2iVaR+MVNN0ImnBhH/ZmRdsQzK
nl3+L26g4MNDQglf662mpXRUrcvv1heSRV5+C6L/cuGJ4spdW2rSmzJlhaxIrOKNJ9uSkPGOaTih
HKLY9lv5VY+3sYtAOfMYunIPaNTUI6goBX9aVpD62LCp/k92z127qcA1mE8zzyfs7yu17Q51z2+e
1y0Vwk/9D2HWYvoQtb/USPPLfMWd0QYar4Tu3ydpz1WvE5t1e55JPam0hZIziYOgnHDsCfCn4DZs
2QpF7eH5K5S/IDIKMjhhyYyOgANKdEDSFxzKy0AccjkkHzXDx+Uz21PKIT57DSO+Cn5A+iHoY2Mi
00Nvk2xACcvrbPtuU9S9+nlG+v7RmGXKobmrO0wBFh7flP+uB9tjL8FUDggZFhHdpc3vkW1yiXoc
k8/VE/h0bw0HiJXb+I9gZk1Q3XKbpP/AN8hfPwUYCZXgen7oJbAx0sOuSKNeUhrh28U76+z2zlcs
bDmw/GDQ269lrMLUVDypLNISdGOCS6/CiH8j86DMDK4E6FFk4lbQATOTL6qoTXC8fpwIJNmmer+p
mNVqq0OzK3Nz4ZJtjiz6gh2hOstvO0EeKgAmFe/KIgAKZibU5A26iKmxJVtfq/EBeI5xxRGUJ6Rc
J+T8RlyGx7xesLS7fSmAR5B0ZRYWxNn73V0cRdyeP0igWVIFmxhW8fxBMf8zriDvHrDO5G+nxP10
46Cx2RO3/y6Q0mRkh5Uw8/FS4hvtDd6qHysD6CYa0w4mySTGD3DbKsDJMGVewWqT5WfwrW+DaYAG
rTmDZuR6Uf34SHkd+34zxIMn3Cc7TIuWNoJXX9WyxyceqcSihyOpX0FgGb3Ni7fgy68OaZxSZlOz
73T20RDB7i8zvDYadzPXbI/MxrtqjDhisAXRbp2B87/8LF/b4gXTQMu8Djwis8gVuhuAinmmjnk/
HVLLMkhhfMsWWFkiMJusx4bf0wLuVEFEGfW/4osC5LfFXK+12+11Ia5wNRZCQoMOG/0y7i6yBjlb
k6sLxn755RYfkG+a9s0pZE5NQwvgam3ye0gDRzEJscLasSh8aLz60LpIAxwbrw7ynr+EHnpKQkNT
ctAsS3LZBlUCFpS/0wiU9QoTEPeMa4YvdEW9/f29mQs3T3czLFBwXVju7Bxhv2CciYyj02P5M9C7
T+LM1Yi++P2QVGtpPSbwcb3vcJ1mWYuzXlW8GBEh06xstz9IkVQ7/iZE9lh2AVjfM3jJS6bkZEGc
it9BqHajp6w8LwrQo4Hukf7gFcWctExYHQRVNncjvwqKIJinqvGuLz8Plk8rg0cS81izQkQkGItS
knooMg6LLEyTAsbg/o2uK3tJ0NzhnOymUNkSvV7vTWq9Hsh+ldoHoDvqK+srPEHOgbXhz4lVa8Dc
/viFGD4IVe2eOu33wiTf/ZluCxw/GOafHQobVPcArW8tkwrhlO7jXYcpCGmk4xpaOw7f+4qgBgKZ
HBGsbrR7Bkf0oO1S0rTsQHwL047AoK2X+sPid85PJdjDLoDbbHbV4IhCL4VaJWhDVhGNNCM3fHmB
dkUoWEfuvWkqv688ylueIXEumxny6I9CWp69OwPs6135qZ0lI5NHmFlU/A0BHP92U6AWEsUPkJQE
5EVhgx1EuXGCGxO+ty4ViQlcsGWbU9NhQF2JI4HbRaURzRIhpWNyiRbRrYikgRKnnPB6huj6ZVtk
iHB51csSO6vHqZD6fi1KDApEJRqQUpOn0oX5naw7vSsroQfCVg21VwGqeZ4R+UtVESPGjYV+HaQR
Mre7/tadLxzlZmZYROaYIDs1zP2ksrFwciWhY3XdBkoor4C4oTYjo901RWffwFaJk2AhtfHKqm1I
0n0p9lWV4ZCJ6EzsOq04uhfwXEJwAfTgqjuE3GdRD0B2ph8VyirYY+gXd9j4nXku1757XLom/933
uhrDwKR7OVwgis3DpFMNHMcpysIFD+z7cLy9kZrI45ATV7iIoVmT8VBtEksE0Kc3qLSdFlPyRmQ7
5eDgJo/8WNeVVlFSsH/dGSzFpi2ocNL643WIvNVP6DFZ1W+UZYBIkk6t1VDf0unIkIKHdPc1IXxR
GsOkAHs+yns/6sbyyrAPd3UZPyutL79j7yRbTVDmMfTQ52cCzlBLMdzGJDgi41uEpk7sWjNEYRxY
5tZiGebD+5e9qlKLde7LtoEmSYSZPP881gs7jDEGUfrP02//k7jAcbOwlByurFcX6MgU9eP+z2w/
UNGH2LqLWJnM+yxj86p+Qo+hvEiG2/TK5e3KIa/yX0e+aXda2BqM6Tc4Cki6XBZ8vALYLuP8pzLA
R0krCAv5bcsucfTH8raHCSeOzIi2O9nZkY4sIjCcpP5qoPfM3Blo0DAajVM6Vj3l5jt72GaXobVt
XzuILDvsRNCv4ZcsEX9epoHS73Nh+x7eJX/CJ0LnG5Jg3Vt4fl9HLn2J3mM6rL+2HmvxT2di8k8g
VJMgurGXfhVhZIZBgTaKZCTfDMFHzdmGsHvMEUl3Idd+LQWLNZEs7Zj5sgBMaSADEi8pawT9HUSn
o4hKstZk7GS1eWZ0e7p+FHW+9MD5tN8N5lWBjXd3+ffFq00NU3g6f37N2vlHfo7mcEzus9Yq6Zpm
GovLoIqwnN/SVZmizBHlyc16d7T2Gl/AFXD+xVENlGAe/VkaCAl1TTPva8Ihco4BsrHdET34qUEe
JGKp8VM17sIz3KSDLYedLr4XNfHc3n++vf2BRT1f5y60EXXB4K97/oMJLOcX7F65Gg8awDHALC+m
e/VdrOHgS3orEZGyZEf4mA2uPU4vlnzrTFb9TTvbpMDkeCZ0vfgzTBDrOnbaq5HniV5GOaXQ0DaY
KBSP4PghVdm4Q7wfggOtI3WHtdtMzvR/cFZSeHNC2QGCoxLWabKrqUftdEW87HVAIhqFzspwakjN
IXomURDowhJCmVLpA0JgEIp7EfHYmru/ZaprPuljRaXmQCl8FbiWdAudmS9WjA1+0clekWP4Z4A6
kjbAHN8pFqUkxdKBTk21TKPPTRzE5TZIVObF+U7NY8aKQ+6zcxTH81bpWj5p5xWMDfykto7f6NAt
jxyUXWTewjlyMGaPuPXIDYpLddLG73LTKbfkUoMzUyNzyGs/umsCfiGIR1yj492otumtFarVdSDX
unTJiDWXg7YgBcKsuIXzZEfwin7ofQqx4rzC4avs8C/7AUHZ66pyFcq8mhWlTiMEiaOTfLOAz71L
BilrXrhSrjBT1QPO/2tdQCh99uNbokplzpVm8BejzDrYOnryX2E2kN4B6J5Znb3c0hz+p1/AkUlu
t2Wl4hBNeIQGHS9QPvrjCNEkamyleigbH+ABz6SoOOOPoGqqEO4q+YvX8vto8nRmoEWm5DRzsMem
YOem8wlSiSTyNiYZfQ61SpGO/yhl9m9GEddc+12t9yzVk4s5vr2zjRu0axxDjk73MHewTQVJffKA
js6xMiOLWFLJZu/MWFt/7dHDV8mas2ZctDn9bkbMttCJM42lUqgs27peCOj3ikX/tezrZdG10h6T
Ll1P4ZbfkFfPXDoq5HeNSGQgC7VJ6QG4sn1z8bYHc1Bo0yfwCz76UR4u3f7N8j5PuPjGwHzrWSfH
SVR3lPXrMmBMhjNC2N0+Q9XDIY386WENHOmvoCUeiuBbSAkNqb8b0wrtoFeQ7hsMwjE51UUQj8Wy
fNwMYRjGVBi3Kxm0RuNxmDGWenjEK0p3BT4qrhnQdz63xuMfjlX3P/BNfhZ4Xc94q/7o8ACCMmPb
815XnEf2GBgM3uMJe3AES27QEYwaYAsga93ZKU/kMhv7DFBkZayczjIvVM73LLWFVBkFpsYsqvPr
QSD2xD74/kNlG9IJ+HjYxU4rvqpNah99Y2rSZt3mSwSkech29x8HAMK0OEtsJexAJSq7tSzEoHWk
aH4zFAaEushUeZcIlQo0IHJBv8RumuJNz4waHXRkEeb2hzNGDbtVo2Ff37qVVgFEVclu+jqWisTB
pKsCMlS9SGLUW6UsgQwbtdUQFiW5/B0bosmDme4C+7bY/TcM4hWgb7sJBsT3EXShTili9EZiR/7S
YQHQDATx0jv/OI/VqQHpKtZDjitfkkEqallOJHdB79WnodRDiC5LIrsCXaH0RpKmLs21gYf3D1ox
TWTPR6nvbH6xEwjmz4I+28NxxtOmW/Va621/PP7kKg5e+TlM41N/M/d402j5Frh3EhvL+mB8jnuL
cNEvK0z8051pZ8tNFqB/Mp2zNN4r0CAvEkls/WexWHU7GbT+uIUmUDey2wn7ablKtGGV4uv0RP4j
+/uGEca+OVcjuYjOfpljIs+ujg34GQ2FxZv2Szt/jQgPJsS+RsX19WvkvVzVQmKLQd0EtG1X0U3B
wFxgk3S6A8HFo4fIyMieUgTav4scAj63xMnk6U2qg/ID12pL9IYdZDxD+/jzQNZi2D1juHk6WTNZ
yXD07wEJAjikMCkuliye3aiYEubGaeJtoJAtuIGDsbZmPFn7GFsbsZLDEwHIJ+iUE/zXDFiQdJYl
LtZFTK6btEDenxRmtO349SP67mNEa+wEwVN+f1thJAyTLhUQVwhq2h99q0OsglPcboje6gKRitvx
IeOzDHzWHy3m2frHDD0xeyXWyWBDOfXvA9+pcwDlGc8h08ZRk2Qm3ZaGwf0bn6DPk9INAEyKWeWx
4pgGc1bJc3Cyx1YK1mcgSU2dryvgsZwJdvhagwDilrnvDqPRDM69+v1fSQa2VdsDj1VgEd/d4JmC
MEDU8kIBPm3ZpZ9zerTZthBNaVKAXJvA7rTMlUJ7dRBuFFXL+nkRCr0KgQj9t8BK27s+vMJKOMGd
W0YDswshxFMG69gVEpEN7mlBVtVj/VxpSq7n8uaDOXowb7rwe3luo3okwSgulrlDIkg33NUfyuAG
W/JKup7HR6d/CJGiE+EBRAL3xq5v8O+veV0p6MpCnyIyzDwlP3s5XQ3SYWSlaKzdg4/4KRLks4le
XA3aixSILL/6t+oNYcppi6NMSuHRutiUhFiwWdg3F5yIlmGlcJf5oIyVKow2WFSobiCJlVoZpmn7
gEsfq9x+J2u/XefrRFtsGCG0yTwNhLi+49Q2xKUiFPpS93QDL5sLMRR+5Q5gTROnaQLDFmfbgCUL
QJcKUdq/AH2rHeoz5IEs/41tXperdqVXjqxmOiTJxNT8QG1yl6059g/IZwZWmbTuywO+kE16vU15
Hi+RfoysrZbaVkwdnY9xRFcAzAa1zuPZENC9kF/r/XMvXfOZ7JAOZpQpSxkTCsDtrs8psRDkfsT/
NTOWa4CRRBXykRVJT2Zwev77wxvVudM+zXJgwRynj70Ij5CjyAQ+xtG+6ugnjYycCZFwVYkU5WkH
0RLKlQHzo7PwLhG7y5B+sp15DTkK69qzkoOCZFUDL9NGI4nNczwoZaTMKgA9GGwMiNqxAXdM/dpP
yYUjaHDyvl86YaSBY577GfGnRDbfyxrF/tFyomaKoj06ZyaIUHu7fhyYokcfbAgoBOEzE6i3Gz75
mR4TV7zo6NIDOiuV3vv/c3AKgLv5UKRIWE30+uKrx6GGToyi98OZxgQZFQZ1oY0URmkd48kZ7Rrd
Fp8sF3CsTsiV24RcTFwFo3CGClrzznlE+Q6ZMN1YypkcAhcStCkk0kiVSjcEc4yTwcPqFxaP5ApI
Bvi6/jKYL/UzYPFupJidOUUmJS1Sc+QrZ23skGfPi0AgqeOfy4mcZkBq75hkosAOCRK/HhI2xTmW
DMT7Hl+FctBJ/7hFeqkpjW4w4I/nFDCa/u8PldZiVreOs19ipV19C3pvJAITX/eQNy8r97czYWui
OYEzA1YxFdWyceuK8YP2RYkZEhq2y0fYTkIK1or4NxnUtkjVQJpZiZKgXwFaQVb3DQmJ79n64Ddu
wiaVuVGvN9/E1fb//mXWtBXxuzDppoGqltzR1cQSmiRVshOG3GP2wkbnOAdM9Lu2+BzLogsdUuct
VQ36fe3fZhjNSl52gqbv2f79Ts/Zv75ogDjhurmLvyMWtRIRH+OjYjg8Y4/+7p14ydwYwOMLPfkE
6mJz8JQXxRYXt//8w9bu6cmRsVbYH2cwCoRkLe2yaIY9lcaOj7zA91sYgFsuNuQ9dmHHXRE//3q0
HtxkRGVL3FJHbpmyFUEyLiS6t/fA5rjN3ORbzALqCK9YXzBUw6+IvZ/C4am/HrW0kxrC1Sa3KfXU
dLelaMEXzGi1ip1rXivY+TnFt6Mmf56gUcf23T8ISNsqlafOsEteL8jD5qGF3zHxYg4qgVkWgN6r
JiPElZqV+71/fLronhC3J56w7hnMR5DIUrQX0mtOV4c0eLtPsRnA5GYrHIO09oJn7KlaMhiMBvSw
0vHdReKB3hbljJ17Vm27ruM6h/+LIwb+5puctoVD6MguG4BcMjy/rWZ9GgxvU/cruTtEkqePHiec
7aZTDS73SGPFWIrkiAs1t+E8ssQHde+iFl0mHXq7G5VeMO0zZHm8qUoRjgsNEqu8a3lkS1y+N+WQ
raUawRRyX3Mk0E5eiih+VkCcT7gPIQpuU3ldyK6dwec7zRMGeNGoTz/OmhPGo6Jn4ycMcCDGRN+4
TrM0l13B5TAGCrWJUyo9z9D++ymrGzYYhX3C7eF1z7SP3850Chpkyqzb6/JueILqQ4YohzQq5BzB
rxgK8fyJHQAWekXjcO8L0bL7gkSW7cn5D9U1BYFVxaOX9RN1NMTP/NcmMf2v1vmm1yayUCere0hz
6KUnZaq7TG0X+o4YUtvUHVakY0+lTivI62++g193QAdbKHyJG/nLx8JMCcooMuydql/kCwqESnVE
kcySUvramvHraZs7tYRUESCtkYv82YygrMt1LbYSU+lf18oLz5yBdLXKOk9hVQGK7jQ/HaPgvq1U
25koGh9ABa/wvlVhHbkNn1jFnYFjICVTl6eARQ3Pe3uKcd9kWYiA0FBhzVvmptSvuz5H9DtWSUOa
n1jjIv/DMAUe2Rt7PwJdhrpg1pxk2uBZLE95osHS3G6KB0xv4tWcdKnZiBTTwHBdXtUxVVgawUIR
Gsk2tBPaJJC9i2oDwVjsEGjJiBxofGf/dDVh3Mrm3HrgJp6q/r1T0PkEwXXa3oDeCRl8BBwzbaIU
EOL3J/JT58kZ/9zAyeBJ1w7jwEE0QvQNteESci55/ByEglrv5V3n5bG7YpX3oOqaxZVTQGX0lG4K
H7sRY83x1hqmer1GRSnfUmK2/ioSo8hgp3feM8Kwe8PeMEhmoAkAeRWLz6YzhlmcrY4FN1v4eRMI
xp43JJh4/T+lWdI15J9rR5PF8FMmVNu9XiOSR6NzEcvNInUAViLRIQq+LahEkKfV/i6zrdNQMIaB
rsKqpt+QxwGKGgdDuewadDq46zYAKg5locoG8gMMTfjH+Cw1KpHXT3+NUzcHXgN/5ZQt1MudKvow
JQSw6b+1mpnI0NpRmPmBCmqETvnNUaODiRrD7SiuScy1OzHctbOd1wTB1yOThcDuiHgzXeUu0u1b
a0dnTI1vZpMQrihWmLxei4u4maqMWnX3q6hUWldA5E2EJJ40DvEGeqyd1OrYGyauCyC/bIUFL4rF
YDgBTh59rLhKVGTMXzkcqKPY2pOkg1wnnbqU1sEwp5UGYMW8sk2XVd476G9Za4ZO6lBy/YIHnsOj
erizjn/im1SBYuZSgPu7nKnFOlPO8aTkGSNoXKi09NAumcrYNLdZtoB2KeYb4cqmzJU/cH4fJKOM
ufwWnovJ1VXngAeQAi7Lp8Smo0Z6VItqZFTwsyzhD0pH+wHWyzYYlNYXZqcbD/XtU6UgOQLdbFZp
FLgYLLkbe4B6T/qXya+3MHmMLn9lDnp+sQ+dNp7LE2excZQcXfuVUx8rUN0M1+PNvU8AZMK6xG94
rnyUaOr4qtBuZcDzNCGVOhDxHFVKemPRI0CQnwPUXjVVbP/WT9eJnpB5x3xD199Rs/ZvFyosc0fW
6FjuxLMu1C5ox8o8SbcITAA0YSh23D//5Yiwy0l7Ka3T/qlw3Wc/iWYvkBeJTmpQpz4qagGMzrMv
3+8kRhu1YkzzYEqDV045+oZHjNt72T5MHeUvFS1U4Q2wvhZQSrPmazdYnZp5GiWXW0gOv4+eMCA9
AJMj2P/lNHBVNBW+mUHvRN9ZWdP91WkLOsHC1q3WKfQT8YBSfgLhfsD5FyApPMDfFAzly7zmRFFq
UpnudsNe98N4GBufdtdZOuI6L82zx9wrmmu1tt37Q0Gfbb416rf0DlsMgsuM2oazfM+JcbBC4ULg
KnfZhX4KL7CJyb6aTVzCH8GUaMww5fQiTaoQblYVI8doRVBrqehm53W4YDv4GohXF1kyQiJTe9RQ
kmHXniddKMLbr/CzFWfowoQbpGMG4g5LENC51URhJSMx6hjliTbNqsZeYkEWPVSoKFdaCkN8gDi0
BVMh7W6PWPHAlDeJt9X7hMXmuFuB/sSx58AuFEoRw5nVXzGF4d7YjVa4IftpY6R8WcLPHLQsFjd5
+Gr69tly3grLr+ksBH1vCWUCcJpuh17Ohi41oRlePzHdVELQDtBiSMoYv3+Kj1aqiaoNZmHkHI4+
7ZXcKkesqFQbQrV9kYFiaX9iYUrj8qPCkbhEDOCzcMGvqQgEq2/UTZIU7EEXu/or++abEJF0h+C5
vWkg0qBghijpFoYHmo30TduHCmfnozyyasQVM3tPzR0YfremDneVbeT5q9f0WMlY1QoI8EuHWH6c
HjU4L5ZwUDGG/yeN/iwtM5jlMRLebHFUGtkc9g0877Yv5YmH4/NBXZyNK8dTfIIvxrLty8hFSsFs
uS0YtUyZvSW4M0UE7cDDu3FbFAFSkkxhmyo/IfiditHw8HgBAP65GdgqDCSmFiL4v+lBMj5BgLEs
Upd+twTy8tMgb8lVg+8MhTP/KAfgylj5o8qb3FqECAk9hWO9sdGUFPWE6HZM57pwyr0v2LXOND0B
s+pN/93NIg19CdAQFszuKAB8I8jS2rJEyoIIdKxyN5B+RVEsyvO2l/FycVOe3TEvHOn+dspxK3Jt
1/8zeD0nWUZEA39aIIIceQeJoRcJM1xwy3tZ0yky5HLOkPrMqGpzWdZd07G7jGjzXoJ16ol7TwuW
0vHiLhGslzQOTTYRjWtQOno629jMQxvSoH7DhhsUqNmdDmI6E/ZaEtInTDhFbizmpVGNnC67Qx18
Z/lgCwVeWOVzmTVmD640W/QgC5blA8vvsLIHzDNawgfbl5MG/HX2qrtuxTid2Ua1EL8es+SnzIzc
wIE8NQtK6kahupvAw07uVMJH9d5VWtJtHVPc7l8zYJs6hJ/qoCNRYREQpLuDo5n16pd+tR6dAdFR
ilVijHe3oSqMM4UIZmmrsszGDpvEniHnGyiohhkta0MSVNPCsBTOgqcRJoBDwP8CWVCu7S7UHS0t
eKkBOa2FK4jL8mFobxPWVAg/4d/JRycuASA6eXhH30aaWdWp9a26CWLGuER27GEwcdFF0edAO+A7
dlNAaBzRb0mbld8y2N4pnwQmewtmtYiZzjYlHaYB2M9oNNgakSpa/5hNvv7rf1E/deU3ZNzOkSj3
hTS7vg0ixYI7RHXWAVUpOhd9gYILB11guIjMIv/0VFOL0mxAizV2bOwTuEvhPJ5NZPU/8kQYbwTc
4yEhHPgCE8CVYjbcw6w28Th2VGd8PYN6s2o4MPsd7ezT55q9QhbjSfxPKk+dF4YY+FpJw3yulEId
IqeuPhJyMKrUyO/1lLeCaF4t3qJwkFoeWyggd6n4JwyyA5MbQlpsBG1SFzfuwkIVTutx2nrTJC1p
VXQUxUrWTJRipA2XRB7YybYXJZGeVpN0Ok45MnYC796GSNyxXA60SpMj0ps6V5Gf8di1DbnfAk72
/JvCOhvCtgTq0iTodQ690c+8ZflLLdmAj+3D9X2VTCjqLjIBdAFNuL3XhP/Lg+lDtxP/VK2ZwOic
nQIvCl1VhCXOTHmmBKXFphBq54eT/TQIu6aSvhNFYVzMTWKi1H64yqJ2gmlPYdy6zF5KFRRYUukn
n9WiIxiBMSPCU3OmzLx1kvA0poOLxuVzCwdxwO4RAsIJSDjXf0enfLOh4El5GlzrCiZ+rdDZ+L+K
jYwGrOeocyZI1VRMcsIflhmmtuIz3GK/jHmJxD6BzQe3PwZjzZNnqhk0wU3KCGIdofW9szUTz+WU
WGAEj+PU6KgPYc6FvKmlPg251tzkv6uYeESNnhz/U14B3KCPiEaip+6yuE7BVrh8rmpCGNCYHSqs
/OJaMqThWVYXMEVYVGd7JeafEd10iziUpAX3D2Jt9XCRFjJzEREms/7aW7ne9onydioIxjfxx0CO
5qKaKK3OIMDuZwhhdS86HqVejSuhZxArgZujfq2zKluVVS8D7zSFsqCkhOom29OKaWYNAX6WhHIT
2dw/HKeQYGMX2fgRN7Q9yu50TIfArDgxJa6kw5wDlhmB4oyMLWDvZYBZJAVConoUCQg4JRum3ReU
X/Biq4W/Xh14pTEJ0KYO/yKfyanqe/W4zzaQ7I+9P7fYidjRO+7ED2Xa4S/Hbg9EMTWScBeay8+j
y0dVt4KQYD3qR/wtB+qqc5rdwyDEHwAiD9XNOKHCszB/T9MTBt6ejgPX3/19DMCU3sClcHQrmMYb
VFhFWe76ZC5vlQGLvR/Q6Aq+QgH7Urypb2K98VF7lIzjaxiEjvriQyJnmDtZCEtXeixlWS+NuD2n
YA+nBa/EhwC0zsdNsHO05/gdyUw4r/pykDL+nHuKgneRC7spFXWWI44m0mjylQzfFIm/NHfHAhqr
rQBVbPl1e+q/m6Gg4R8Dn8z4hZu7cgthzDt1m2F6ZfzDOOipxgtwA8c4H1m+re/DDtxGoTSDXtvd
xRHv+UnfP5T+WBQ1JuBjRRj2H2Zrf5rf5mo/AMoXyHtWk6rr3CxAop4wZCvbP3OX5/RGy5AWZ+h6
Z77H2etFMWk0X5GA28Pg569FuG4rYBxixevCqukhiYlCq4iG5YjdxzSEChu9bdXkqgE1PApUfox/
ubBbTdC3fuDzRzWg36KmIWzeLuZYHnjJKDIFRwdEi1kO1+C/rNSSGICdCRy0YYn+D1YAuKdMiEIc
ImhKkZV3LxFuKtzH4eB6zLBGSzGI+suZxGbaEFFq1PRdpGiIETTJ5AC7R3pjdbZvc2Ps/HBt8C4y
qPcnuUlbRg0HO47+bcOzWj/V2WZZZDWL4eWRy7J716Fnb2Utc2iN6kwVHXTdb/y9jiKdX6P3bK77
J+x+war6oQoAZasp9QaNgj7nzKw8gE2GoyH+hTIjdLDqNp/qQ6WS1QgOa5gutA1oh3tYt0zLS3CZ
o5D1DBzYOwwJ8OPa6Krm12XY5BAtmziCYlkPkBjf3LHNxxZIroUQQagHpZ758OR/0pKbolH9sL8f
Kjqe6NIam8R3/h7EooaCsoylSXPIXbIVg8slJ6uqDFApidRmW57xXiWzsNeZ9PlFHmdvG0pgw0PH
WW5ji5Um7Lz0f7BkCxZV8Zd7Fq5x7oZov2AADL9KpuF0u84w9eAmrMC2aD54+l+F+n6toc1wkeH/
7NtlMsb9BlDkFC6scKnAVcO2cbxXh1RCd304chHeRlJuQuglc+VA1XkhgkuYF+NhD+9wCNzMmF6R
rz4ZJyyFQbofciyql6eNwX3RhnijDhntOcn0joiqbB1nZP5yp9CemnPFtF/jpWg31AR1AObqVJgV
ys328tzScTG+hoEXWR2CoVMzMwvOs+SzmhQLFD5dZbWJQkT97mjtQWWiBF88J4uKrxNWVLCQGpes
awA685C0emkjzocKTv/s/Qg7SFYNonU+OESvhPyNn06FyFAjfT6wtNw70bPPO3Ab9w4mfgWWRwTg
RKBQOk6OVhJpK219L30oJALmQTZASeHJxILwgpOGvL/8qELhEizv78hlC7Orn9IZmFUj7Mr/DmCG
J0JNIEJedwwzS3ErFF6ldNlBHUPpCMrCrz1lJiUnw5oGdfirpkvnm2wzgBoGXoLl2xAbisNIln1T
TPUeWdXt6CEavoVb4YTA6bdQRrYdk0U59r9ibVkr9OAMVCq0+e8+79+eAs2oAgESkVsJA6438FVy
a1GUTmoTNLOff5Dw+ZiYnxdknkUAUIF+6Uho3bluNIYm8YYCLzPyegsGyTBhPBZcC7Z0tvesmPx0
ZATwptxvoAoVJLy7WvB6ZbpbP0/QsoadEdkQOExdnMwp8ISYbHFbsQnIwI9Z1FPzj6WE9G9hE3GE
Bh6hi79XIwbYDP3FNZF7DOp26MWN3fx6drJL2s80OLyWbBHw3NV2bjfGDTwhyanrW4+mzOJMyTNa
rkUxWz2hU0gJYkhh5VC8aRtOdEuDFuZO7HupgW2MQpxMeJK+5zVZHuow4iJrgAEYmKUE0BdzDwLX
SBI/8C6nhxF6KD9opsmHAMMDiUhBUQpJQWPcQ4tSoL+Lr17ijOWslQv+Sd2ejGDPnVUCdWJOefZK
JHHdVk+sS2Rqx3XD7wnekOr9vJnIOKrmkVTN4Y64UFN3piGTvXUsYPAUNgYXEBqG3dfu1BgBh/yz
5KbTQttGJFQYkOztzM16icj3TpXij7zXQRy7xS1Gu1Z3K3o3PNemCewg61rVgoCLpDsl6zHmwZef
g9zbel0EJfHCP3yOCnB/G3DL/sbU1BuMe0tPxfc4BdlsHS1ieP2JCeqAJE3tOd6Jy/Ek3VYlX2DR
Ff3lreSZGFrsxuUksU1l66EfCKEhFUHGtyxr5tXmALwhhnHC2AAik3FveJYGQxzJCisYTgvhLszQ
hJR5M7UO67U8tIJ57YEOVbOcC65tiSjXkCt82XcSdC1sXY9Vhz7Nkmj8SOEf2aSI0tTZBnymtPJZ
180IT4h9rPk0hPhoza0FaBB7hjMQCEW9egdC3T9aOW1hujLcJQWxM3Dp7bOKbmqka+rotLWtfbYW
MpKGSdDnyTasxNfM/WwuBooUQY+1MRq3Gz92TYlE+b4eVaXAen+u7uJmbz9ShQMrOpxL8FVM3jHp
rP03v+rAOvb1kNH1hrfBy8RSSWTtosaIoAqwQyxCXzjUzqAyASu5CFhcksAKjblGIobb4lzc1aMs
cbZODTTHroCTf5Tw1e49Qhx4beUn93J3MoMv7Rj0LQm9aFLH0wcSrWwwVaUquUoWJByUQ/ligqIG
PWBll9TZBTYX6O6LlTd7/9pRj3YzYRuCxNP6INzlFiQIQeNNF7Lg6SUiAjAFEtQzk8d0plc5k+U/
qPZ0UkfJUKMESgtTj84VQAxFuLuwXDVhOX5HS1K1OlAbaKKibsGK1K+Zm7TvttQx2gQeuCnj7m93
FYRqonzBojfxLsds4RhdR/575NvE8j34GsQ5KAPXY+CDMm9UfJA1bn+pQsOxO0iRcfLC+f+BzKpR
7fS5p55OXDkgv1Pz6BcO+OkT18Z72bf250wGZ0No+25mAVWvCmEUqShzgZ/wBUbsGDz8DJHrd9w0
2+a45KHQaY1lby0Wr3bwX7TD6+G1vpVYDK7O748dQLmG4Ty4MI129MdBLI3Mv387tx4HDrJrrgT3
yN1Cxo4ziyA7DOADkb51JBVDWA34+Ws02RC4fEEW5jW8jDbwn0tm1TQAjEmSg+Q3Xf8vQlqkNgkM
/6+XELx9MMGdGasK/1ZB7jt10l+kjHIF9tP6u867FqizcjjnQTROQZ2eXdG5hzEqdfcX/IQt3esS
pQ5+hvrfPNCxiYiGhP4mhoGntJ4S1JZclZ9Ek3FYu0j3rGz8EdgIzabjDDxR3zz7hjQAt6Klamfz
IMtWMP4Ix3Y9DGXy9Z1NfZT3nTfVWvBlDIel+gdQtI+dfhhkhMJicRjVEjsPCt/SeFLRoj3Xu+/Q
i3v4Pdb27cExi8ADyvxOBNsjwQ7f0a7r2vW4mYF0tWTo22b0LEvWddWAlcrvR10Ovuhwm6gFRs09
Kw/X74u3dOFSWYeeqmNXnIBv0aUGNrVYoeYcVUXGVt75a08wWeQVxnKfW2wkRSV5SfpFpI1AmnJI
ZkR0lUxTvS5JNVwYeKMLKwIntzTcUVr0iWEyLP3FVGik3n1JkqrSl9fRFdj6hb9cVTsZcfONChMw
SzRDPNhLnxKTxVxTLa/HC2EARqUakyJe3aJbqqiVkE2aNspd2iRQQLzxEDH2NcpcdV8gcQqS/1ox
y4oEF1TNGjknFMr22ZWOyN81oNTxSUdr4viakztwFvGqMMlVImJHjrCuXs0Z20M2HEUv3N0uFFUi
zbw9TkajI3NFw5hJ8F4MyHOqWug7t5Zt1UGAU1uU1k7vXMDZPALZMuis7dUy8VAeuV3n7zlSHG0u
lGEfoDyBtd27ULSAkHsaSY2nulCRpex0O/GaanhWFIhxliZUTWJvJjPDNc8bUyaJK03yrMdnnih+
M2ga4/U5/hiPVlXI27iRpycvX1ZjaGJ+aOahoX3RggDa76/bm/f8u6JB5R8b8mQ+Hw3+BQETibkP
VYCFYRl/jF6KEUkjTnvDiJY54rERS3V+Q+qHb65kOGJGxCuzF5y6lGqx++Wlup0vkEp2jFimQobj
BkFhUhiT6LUv3Vx6NyWISHo+4WtX/Q7ESWK3X4Z/KS5TlZDbks4dK3XgVbRaLKncBBXb8qJ+cKxu
7EVMQkDNFp/UhbID0um9Ca0wJ3NB1VFyKkdiDSm9a26T2/1GPYkUtenYyn4AiXSA9heO8SDfQ0rB
MWcgCJaDpdZJYOt/Ftxh7q8/KSNAPmB8/P7HcvfeslFlXr7baYdLCafVwnpTyX8oVstHwPzRyq+q
Ahp2wleASlBdAO13yE2jM6A2FN6Ku6AeV+PHkXcSH/6SKNcaSXEIPx2Cmk3Vfp9Z8Km9X+phXZjN
8DF7dEuI8eGSJZZLd4MC/FcyysSOXbqcoXLBufg48G0zQroVjlzMoxkYPLaIzKn22aeMYmmUV4yH
9B5Xxs5iq/kOlDkqhLlqKLSA3F/wW36AFzqc+ayleKw48nV5hotx59jRbiY4ZdEEq6H69KVKrlpF
DKOh0tr7IGDCr+n98pj4BjTsZzU3yCwGGTuhELxAiCkNBKXX+FXGIKBrvegg/Dd6x0f3dQt7bJY4
eK4OG8U6lO4+QIFmt7QGqbjAalPALLPfPlj35iD3dfu8h4AC11hpyp7JQMiChTZRFVp9lexx+Iw4
8BVHDoUbO6aOUlb6UbFqz95K0OrKbGgJe6OySDUzPfN+CA0LQyZ2t0IGZZMovrYpk4g6hWNKaJKa
a0g6ncRm2cESwjau54l6lmhFIIYc8sVO1XKiA8ypSoSJRqE73jEw++6jCUZJr5pWcqrZlvNJ2hXM
yRlfV/9ozcbCU39o91x7MYOO+WTT+1YH1/1Ys63ZB7ZIu3dsf2KYoquiwWm+4G8PLjeIBPmYJqdM
TQpEuC27lhXjdVSJNHNBOwTI3cT/7hNN3XxkbJuJeqDNws+eaUqCGyNIAxn48FMft/M5zwTJglsd
H7ffDscPAld5UsJkgk5VOf/W9KrRPeaz1AssDmueMsfD0wLgakKucRUz5NNcvxxWBMZzTjPbTw9g
u6aitWhdvwbVZ8QW2qtxlgG4t5GnHnZaUkbSvbz0plgn/B/ik8+QEmJUbMtb+LB9XxP50zak9TK/
5xBSFWRA2mbAJpw+eKfnG0oCkP3oRMECTcyHx2REHzv6k6OCskppBs12IKFGC0ZiTq881otc7Dzd
a2H1Fc+6C95V9iuHbLMC/mUG5eAPB3U7kFYjxTBogvI8TkH2T5U9Zuv8H5RC6DXz634g3CI0krHk
JT+bygeuYioHYwZkx6rNfB6r/WVVybaGz72QkPzA16lMT/YHdlVnMbVVxkAjRfgR0AHXNGlR+1wT
RRF44wETIxcH8q7jzAmXeTMVhwBZc1JgrSy1lJHR9ryEsCG9Ai/7z2cbrSZ8RerQj+SK/wuwSa5X
XH/v6WceGGek5/J4bCpA4puNLFavNuqimc4EgLXjupIkK5er4+lNXZf020JR7CMS4vnvHfBtw1eL
i7DWSKuXOoBP9dIinrqNU2aI4+1HMBjrKq6TcStiwa7QT/TouTKDXysFgStXO9Bhy/eX6vxiJ8SG
MDFcjAbRQP8TbkhwBoGHJ5RQrmhAcTk0JScCR4eCDgG/2xQIjXTzkFaAw+KtwhY+VYeUO3RNxt+D
0BktcnNby4X4xg7E9yIuHB+JrYkB9ludMP7AAhz4QxMVIvglDnQjxpb8f2+50YUUAN6FZMP8HjCG
gM38EbHeXmFwKTKq/Rpurp2C/J4e+c8MzCko4VRuXFDplTZoRjk24wMYdnYuTACuSXO9llEGomJo
ztL8FwuEVUGIUC+nbDmGkdbVmMbyCgJvDe+qHgj0ujn82dGSIjbyK4moZ5vOGC+WatQau5mbIpF2
6f6CErewdchksA9N1V9ZEueSwEt7kSnt1PNIBloHpOc8rQgCvn3hKyBqV2BF0e6I8hDZPNGFxv9E
R7VXrSM09upA05CGDzf0XbTQQcQEO5TRsqZ044EQQoW5QwKzShS1dfwiMP7Ql5TH+K4ZgtVFMxgY
IK5yIMih7rd7rj1efBl5yfcO3Xo5hoz5FNk4MoN1zgkwFU9wPqbEjCmJRS4E08oDISFdlQqBpPC4
cmp6wgy/HkNrHIvw0ACs1Py00/ykkpW/yhtnzt6MfjYzIFGWznH6cevdXBOi5Pnx8MxxN2AaAWt4
2AmlTu+3269PzlBbedR0UELAgL70PLhE46YtjXttWvBL1McSzIbtCDf5adtjuFEjXY4rWr2J4B2Z
ROm2R1W+uBYP07hIyj3aKp88K/YDnTnjRn7IXnT18ZQkIeJDDZLEfCrVG7RorRBO+ikmzmQLAIkf
G1wWbd2seysRBXqfm6fSAMPPKh8gIJ+t8MFFkNzfXaaL9m0eYSXj21mYpufX9CUPrj2tkpTvPWV9
Er+DZINRjGKRCjHEMGWuyMn2AGnvfaIWok/LBs3RFCYuE9szCP1yjn5YmFV+NqKGs4ao+NmKwcYP
mPsaOudlPIfB6S5rxNWl3zItJLBMV6tDpAZReDGIGb7PSq6AuzPb7YteVHqcaj8ZgKl0dlhslt/N
pXgl4dA3W0hauCvzMx7fqX+DZSzMG39iq4prLURldwm1D91chhcWbPcFWIJwSyL4gYUD/1GH4yG5
0Q+uduC3sgk62icXLxvHDFqILANn4fbWPCY6oawynI2ZY9U2mRxEsad8+YTpek+UiwSkmQ/8ISYv
UNqPsSpjvMEAlifpi+rAHOYdeuNnK6NoMq+uf8t4z0zGdD9PobGL1q4SY8pLg80VanUqwqy7tIxb
ypmD6WBxr044/uTW/eordNhvswExA4egoQr1YdbVuLJr7AP2G4LGbQhdfC1hzWfHvaRDgtn6uClP
hwz79zGK9yGlC3UD2qqCy2kY98JaYK71quzrmCG1lTc3Qby3I9L4EBPraoXBK568PuD+K4Ac+wMf
o1TbvI6hh5r7zzKHuIF8OyyFb1uGgXXBxn1fBmFLBOVy0CA+4awwyVqxocCe31ryEt+HvkbemONq
ssh8C50imZGFYrZ53u3k6lWb+xwK6zlhe1KEP14nVYq/lnlVKitXj7Zb8AwSmIqmSKonf0fzwDSt
iKt3Oep1TJIGz3ZTtN+xPAmkDC49E84MRYTUiDZjpTKU0ggCg88p1bZdcrVBst/AoAqtKrq0VnJX
kPpEQX+Ksal9qFHVgMTjb3Zwe/HRflp217KVX2wWfCUWCMrZ4zrbtFNRqCsiQhB+NDkgRT1FFRSF
rHXbIsOXVHgfW9vX2OxDTEoF1Cu2WTAKCAHoFwILRPWJLXbU9AILPNy3BBbiJRSCMHPwCPr8/Fen
H7Ptuxrb01dkFXMUN+6pn4F0CDmjDpep7vnObq1JkZiVDzA+imo+U2PNJLQrbhZMG1D+NKzYdf71
5uL1F5ltjhIqprkiM/egGlmyX5Z/lh84BjNE8phgjrDZHHB70fqXg40jzN5ZDJpfAFKjlvzkffA3
lUHo4DbYacUIRZ7j3d9IhWQ3BOSlPO3amyeypls2cuDa/q3W4Ve7pr/oE7ZKTIpJyvvA3liOymgr
lAkLeWH2WKH3Wgh1RD5JoW5ZmpziYK432HCTmswp7QSxEmJ7ghvCJ7tHELgvX3hbCMd2NYm6xcbR
qn0WG2ZmJMsfgvRioT7ZTsgLiI+bWXGCgVeaFvYzPewNC+yEDpC1aPzzLeT9jE5RKpIPzc9SkGWf
PnbUNsAn+hwsVRuPAhM2BAB049iVYJZc5z69HIAuz4Sbzvl4hZJHo4NqvMfzxD7jd3ArJZnP/nms
PfQ4Daa4BUPvm7zsXZmcHnfTvLzj7ysocJOu1fPbeZ8xPgOguRDGSRHEcVFwCXmtfdF+m7COszj0
BPdhkNajwfdCsbm8Jch6DBNk1vT7yfKOewRouevuFoxpCAaDYfA83LP4ylR+DRAlFSgJRklfZkpc
4alCpL3By/WtriBk1oO+Q/NCU0+mW2UBuNXRZMkL+28D3SX561GiBr/a94bJgn4B/B/NWmxihMid
QygYu508W/AztnDC1NmNEmI3rMTb3NJB6XjC+8b5fO9OVQXprucssmJCldQLClzRgq2KCkXVdoZL
lMzEKDzzlvgzdYJJe88F6o9LR3morMoBOC1vOgFobrQoSlxjtJLj+laPQr17b7XM5YdxhWhlVsSJ
9axENCpUoOnroAN/GDTKFmfJLivagrdwYtTl3uhgiustdLZGWI3MAO+7uMHnW/0aEoNs6PRbp5BK
mXWJ9WetG/Tq9vdRASfH0qULA/voszXAdhDNsalB0ngZUdd10RGj8Q2ElxBmsKHpSHuvNcLT0RZI
uyOTYFtWPH32hSG7yZE2tXvrjwa38lCvogbzsCN/YPGyldC+wufJ8cZJu86shOl7+KQRAG0thWto
MUGd6CtJ1JFyQBS7IvP1zlhG8PNG0wgn4rWp4bf7X6LM7PQwQUaNUJbFJWwSseKFf2L9ZNdJDjnR
0OXU4cCzcHxFXoevv//Llz1UVkvgNCyQ368W4cNxgGivp416wQ0T8eZ7KRFPzY2PfFkK5SB4h12a
BDRiUuC5l8Z4x6eQMPASBL+NDK2DZjatj9jIEEs5KQljB07Boqj1dy41u6ZD9gu6voaQ0flDpbp6
+8sNtGUbPqWakj80fj35UTJ3KYsqJGsfzNquf109gU41aUdQghsgYZ8O3ih/yTHBrBm2B6/pQlXD
W3+iqPEl4ITGLCwTaW7IdkBuPY0gxxMDe+w7Ic64eZ2is21rtPpg+WSq7rEx+VTtFy8t+w+f12HW
7j4uSoNe6bdoFA6F0zJF2JMIZbCsN/j+D0V1Sw5pw6VZChw3IQBfPY+nepwojIzxsgX8/n4anCqx
FimWd1IThSN/P7Im/IWTN2kg8zdgTYCJznvygSsut9GsmaKa1E8Mru5Jz6d6irtWCOYQKfOHaQoh
VHj7u4wpq24I7iqPJUtzlL8oiSUa4csnUY3qA0XACEvyYXhQdhTtHfrle8x+fvYt3YTZ72hMixZ6
WQ9d8r37fW2Q6XRCpXiRFeDOENWNAfO+JHDk5b6MRsAgGoFSR0pNBMrchOTFUZSjSK/Y+Viv3Tzx
inqrwX1sIjoCShsjHHo5IclvpAjhivwe/6glOj4HBk9yra3ndqztCPhFTBQY+YA1o3aXBvEHcZ6k
qKnzBaxHC3R49tp9rWzBvS70TiHqTt67GRt8FNqOG92I1oYpiFjHItARzM8jdNPnAIAJXUfv1+aC
eWdqnBQxRAtShdrRWm2PKzJDBbfkJnPMoQEaojcDrnWF3kOiJt/fK7/hdObO/poHERAMhbxe62MW
/e3xcN0/rFMomFZbEm95HoF4FZo061jHfbNzMth/eb0RzZsAmU2pvYjN3PDidFexkV+FH4FhIv5D
0lqBgbTz1pZ9A5CQERXTA0y6ZxkBMPJfO3VtfMo7wA1e4R6DD6ZOK44K+/FWa4uxV8qXj5RAmZ9W
legTZcHh7g6N7WnPHthxfzQX8ocY8HAF0O0dZPxBWhIBsxMpAG0dj70Q9/vZMPFRH31J5Q/jkESW
9hgy78fpJJXzXKCZHh4cV2VQPI5WCvNH+F3zlPm7FaYbDa+bD6rplGLXigqUNv58JiHt96jMY9pT
LMJ5ERcb4wZItdfUW1CsPjHkNedQoODY1PBhG4xxCUCwjGD6lOrhtprT/Vyug2VIceGJOqsTke94
FHwNc31c0uhfTElgqyiukdENgzxvrb8Pwp2F+lMvkRbd5rzCFh4PMGkB+vE3QeuR5Xoer0A6qE30
w3Oq3isx6dIGX0VBE46mUi23QN7k3LVqKlZokEYRFM5xLJ5q9UHyELjnj7rP480Tfi1qoQk+LxLa
OxAEAnrSWpJYn8rkJ7eesRdluRMjkyVmdNCFIhhLc8Xximdwt97KuoPdjwlwq6iIr8uWXPsnyvRJ
QlvR2OHVHaHlKfcptpDt3KYkqZFebhOnlkaL6OnTL9jMf+4KfCxc+djcj8DPvF1x5JYmDSlpU5H0
imkfyKww5rDjobiaBrULveqacfocCin7KWhvQP7qwcrxa++4oUKkMglivd8mGda+qSb3y7iQ/Sdm
NDDRooDHrkWde6Leqe+I3L+C9aD4Kvbbq7LJ9zM+oY2jf7IDmuM7I123c+l1cnmFH1ZwFptXbTJH
/pDL7w5p3pwmmmSC/yaNYUguqaSxC6w+HTamLBNJZDRe/YFE79d+VVMu20dDaY6oiIAUCYLzqcnX
hxzPSnIQxN0N5loeTB4ekoZlejsruPlTLgc1y+Zln+EPYOcNSVhOfREHZiDTGS8r7Wcq633qrasI
/1FFFAEWvqZw1RAn7YehBg76SApOSGTk4yqdXURBh88YqNodsptHxj97Jm8Q0MUUcy8k0qWWUO2Z
r8TkiuntQh48rXeCje/Fb0KcZdpO6BGgdqc7DAFnihFnlwf+LmG/p+HJqy1/Qlqf3lZhObAvPIoC
rn9yAkJdoZWHJg3Lcca7bvwk6frqQXuRrqX7Uj7Ps7ZWIKiRpLVQ/OhTLknYcLcerqX5WZ8iGEcf
mORQ6gvmeJ2RsPBV/e63lTjiZ5btH86k8MiUk3MfU82QZ4q8bLMZ2Q7hrnF3C/HqZQ67aM1BePat
GCCSKsunjWAl9UpFuhgpzSWskA+vxweqc8T6FmrNpcYe0W0Fpm2OgzQ44hTdl3mxGQQDaqasXkz8
SfzzSDo+ZOMXPVGfM2WcqLCOnNDu4yPj1+Q6yyeG31YnTmGGigExcZca/9tTgjxN+uXp/ODLz5pL
0Not0wn5Y2l06rUo1k0N2XBgwLcLwrSXXh4Y5A0VEsOu/k8ImV5lQrwCIDEn9t6zgscRtS5TbOVh
LO6F9iCOS2I5kKimjO7ZjINUifta89lCQ4OKTd57adfsSV2g3XNXul3bq60RoW0JMTmH/kmRWeq1
hR10l8dqWy5eC1SS1KY/evow2E4XMRGIZr8fK4HaQWh4lbhmhQoqsR5AF2dCaZOtochqGtjcE+F1
SqTyCk2tAwtLWzYphiUoSyVklNmgtQsU7fjzbrfI1+cWjrXgJvQNIei58qowVeyiNX3fP4jk7h5v
4Kf2DC6vidX8MvUrJStK6Jnl37uklLlrxDzHXdMt24mkyaxclSXNhLnIv5lV9aWf1lrltzpYmGUF
dzS4JHWqC3IrQyiU+Fcn3moC3Gl0Tajb/3embwMykOy/Z88bBqkMfxe3rLqiea1vyft2RyzxDsPz
fQ7+DljEoExzHbqY/5vm5TuJovznM63SL8pjLnCIJnlZb2v5Fiv7YSbW08bpCtYeJgwPiCvO0sBs
uCse0B/uNbjj2MzedYSVYDCSX+Xh85hmdKWZMwfD0sFIBDMd78oYgl+kHC5n7AZ/D4zjtQv2FKsQ
7G5/+1ilyqJZA4hoEzePAn51daCdmuKjVYkH2elMxdu7/JxNPM7R1BXSRs08hGTlBTtkHEW0c+IR
00SLBF8VzZMjD+aXb7cVQyB095Nl1ClAyK3mAosDvrQFeB/zavZ67YrM7Xyw+/HcGzKPMgPSUSNk
9gycLuoPObKw/0JKRRWh/htfi//DIoaR0TLQBFE3+z5CkUgJqmFIbp378P+nPgXXX1n3CZGOkqoW
Cqvk/s1+kwRHo2so0WZ9teL28jC1utw2aCCSHRdUrUku0g9mPCKEBNd8Kglz4XmJW9nuul2Pp5EH
Sis+nNSqnoWjveJALldGy/06J5xWz2N6iRJna6oOmvyErYGIlHVhmLGr0KF9I+7okbUyuri3Xfgb
I2mIvV3OOqWbzmzsi9kd1NeBU4KL1x68TwezXIsYwxN/J8BEzA9lEIw+mDkTTDniJGMVxvnmwTBL
XW1AxAGpHJq6C3FSNIoN9dFYvMItiqyAyb+QeCJ9dYv8B5iTOEiMPB2w8JZULDaxEpGm3FxBjstv
zsGoFlwXyjhOiV5ojnGkTq6Q5mj7bQedM6vsFgugyjlq+EPIyFsLLVBR+nZrsHiw5aZKt/3SpCNh
vpLaus2z1KBOoNI4vffTzXWACoO/qh8MJ9rap2MbytiiwshbjBlLAXzID4r1Q1U+fdsIZlsOIyKn
h/QizDdec7nzeTxBbsUma2bUs9CCBy48uOtf3fqWhS/vVRh+ndH1JXSbKv4ptO0esmdEgvGq8gIZ
PqQst5ed6KLMyr8VNLrjr7ae22BEnHjulg27rZAH9FZNQXIWVeecnmxoXf+QbNMzo2VZY5OTEzkB
X/H/BGyfw4H0blFciZUkPh0D6JPe+S5Cn2XsSezphQd5ZmyN1pMMeIzixI3TnO89fDTJXCRmwGdV
gPa7yymD8omOIwrHPqK/rjzmPGe0iSQUF6aT9Jzwvt8N5dq1MJ4yYuRP2TNaSRUsr5OMTrnyq5D8
qKHg7EudUklwrUAvgqwqMRuyUgrjEjYylFBlWQVJYzbF7Whq0alBDAc8NamDFca99VyObdLjOdS8
bKEvCRSRLPTP9HkYnFa/akiSbudYURFa7Ln/7MY4oK2dvTcuX//IrxOb+dpGt5UCCJJLxpv6ek8K
myy487qZkwdZXxk07UdL0mkt6CibqcTiZkC155DVOG9duQm1xrWRCCY9uE+EbYfOwYtBDTS0CsSP
r+lWGX9fh1zLrEGRnZiq6JDvgqZfac9qoAmMVQdrXKaUDKwMRy9Cduqla2i7gpeRvGbaT138h+bv
1xVQYFDpUf8HH8TtK3FmQFUDamfTkqISf2j7R9+PloX7tgWcVconBkBHqymjt+AB4n+wVYBNVuGV
lOYEsykYGD0Sc9QKYSIRQaSMRYz1bFX5mZXfshvv6ph3LziErPcHMwa+hq50m6yRMlaFYwXosNB1
/73mnjaFka01QOf+yYQb1eBrUUfuty9Ya6rDCZLMUbSoeINziHSHpDqzeoKgLdb5xBjvph7ttMz1
vazll5RjZvQiR+0Md9+K/tz4lx7AiYXNR5cTb+CtkSt3hGu/AqspFx4/ZbeWviGzhGh+FWysI/OA
yT16RE83yXZBxW983i5H++upnPjqWUxaUiXGlckpEOft5LgEMPbDKTKTvfQSSvpLF8n66Y2mWj49
HJrjQplel5J0PHxnK89Cg6AjDClzpm5k8NjdSc//NMmqVObmK5vZ/2yN6nRg9p92W5yf9Q++N6Eo
algAMnTf67cdg4ceIDITeJ+2CK8DxBigViRakoVymYZm4A+9GLMt1vFfyvVTzc9WF+wy1W1TQwRh
RxresqTrfLvFbSsngZwKavm8BhW6NyExc+oP407LCgp9kr4yfAo8/rOoEpqrkvmiJnY6Snp32MuX
GzamadjLp5Mae3iTWLyZC/MO0IDD3CEWxHRs1rqdroK6/SPDTM2vBbmgQB2G3E1YRah5jvaow7me
CCExoD2b0iSlkXMjYAnvm2NLXDYxXkBjfA+E6eDZarB/gNlOI0SWQeWv1bNhv+xgc/2itWhC+ZU8
LjNC2PHk4wmzSwv54GusiX2n9LNRaf1yT5pecPa8OUy0h6qQhC9pGebafRZajNSK/RzyFAvXzamy
LOooDFsV3TMbhG4Ae3yYwQhwKf/rqbdOc/dofzD0yousTsZQq4iH9DgiU9fPTLdSfN4IV6c8zM2a
+EE/LacBh9fRqezV1lRsHOuA5hKhuTvmIR1sH5TUaA1ggtv9/kTGZ3ixjfHLs+/1PgbeMDmNrFGv
ZPNYqS5YFY70wZirkc/A6BJGvVFQQ+G9FlUA94moZnExN87agAbXO9z7WG7I9Ujek1FYyoIVv7z4
l2GinC7xZ17LmWH3G2ProNJVmMPy23SQlpDf3P0GnQ4HVqU5ypIMvlIjPeOtQBd5LPz2Cc+m78Al
Atx1z+cs6X6+/MOa0X8L6B++qyMwb9t3rMXJPsED1srErlZOfmRWPP9IWLHsHwueS1MEH6kw0cg2
WsqFEbWG64Lun4xaQ5eD2q+lQgy3TOS9fd2+PFiLnBluFePGjb9zGmpm02InFaLVRKXqy10qVF6W
7GH0jYLjCy3npSl5leqa1Q0HOaKCnMcfHRSW3i9EuxJOqwqhaxwhUh7QY+//j82H86zsOPD+qh/O
9/l9wOmAjKXK9Ihkvrg1xUTXCHsVn6l4TP7QsL+lQ0cmFepbyJCGzXbrDv7XlnRkMd6oz7B7rZtN
K5OMEmlfwO2NBYMNUcjxyyrI8RNDjh4f7i0tMALYWhdDxLMqn5YGte84ZJCSiTT1YaLO9gs8M/n2
mQVIyGGNeylJVo0627yW3XXc2/B+NnMKuZId7lbYD1hgH3GWrTXALu7ug4HJWDsyHaBjZtcSV3ta
jO1QRnBNxgQfqprM86dDhkyb25TWnZrF6vT8Hb+QjmaBboKaY+S8XyF2xPwJ8VlMh1R+yywcroiD
KaeeoEafyOvGXyUf1MTZwmF3uTHsY6lH5qStAPrWJ6dg3YW+urHja6Rp9mmT8V6Sf5wV4c4um1E8
vuRZzSgywKH4BXDkoEvDiXU7kFNQddEw1X6Hb/x+EL4CRCcpEXEL8uA51VN7/6VNMh9bbytzIRgT
kzEleJUglRnY3TGk6nHB+6VT+BmbHu6AUHhL+QQzAruYjMgT5uMFW5h/fstGq77bWEAkEdPU7gWv
sEl5ris1NWYgsEJD7k01NhUUvJOyqsAxvtVpxpJh/oFYpvUPOv9nwUV0ZVMtEs5pLR94SGTu1isU
4YIkRjw4N2rmz8r1tEdXj/IWEGMg305IaM8/FRTMp5oOLWmk+IHYOJJiuNDUomWCDkLpYg1frUOe
JtgbwBOUapSfwKaGUacx2hxjIZcr9odBs7+Tzpb2epSVHmyzkvYBbk6SYSwmtK1c3xiQ+FCFOkQS
QwvXeRy1hieJ/UHakFrt3iHBRsBapExrUy+sBDpx2mD8uLxKKNuIQVJoc/CREXXqjrbuu/CtXmMP
CNxSKNVQ+SflzDinCHvRzEweklJylJ5GGVdr/J/KFk6v/n+nPsxF3oaUikjKpOVezaSPJxt6B5uT
Fg1LEeBg5O3NW3MAqEEEbb3pi36T6b+1BFU5Hd4bmBdzDbu3cyWZlyUsFB7rPR21U8ijWu0egdei
Jk0Qzc/x9ZwFl2aOY9IHSUAGJZvrOH5eqc/Y5Vg0bIPoqMiF8b+sAbxYz2bOD4MMtwvrttqTJuX5
44tm+rakY7Vk/jJ2gh2GEcPZAxN2DQrsBfLYIeaPiLDr7+AtQ7joICFO4hfxXqiu3eQsMc/UO8ak
MeQwHRc09NUvR2/28mX4X9P4U82OYoTAC7vAsk6wMFs4Ea4hXThsP134K+iNnIqRu8HKqb+R12AU
tCXHjSAFzsAdOvA5OvQ8kIh4WEFxhxgx1xkPH+Q2LvdJHE08ZFoo5UnGCnirmBKIEYCnaahDk5au
Vfkt0vbbrBZGwB0gZ0zhKAKayfu/aBEh+m38FC3N+FHEWjA/PTSB0rYVWOIpdZe4GwRplYZcYWbZ
QLN6XLprWeVGZiMK1I//I9/0wswqCq1fdfDYVD3oP0sRFTVKWeYmgDxOzCzAsl84thhOcSmnXXbS
w7Uj6YRvOEsDIv5bwynuNCZPQLZr5eKna2qsymEZQdJ1yzWGPylZ/38EMCtGQamBPW8K5yQC/y7R
nt43zGRXGcK9VUv/rc3Xddyn1Yn0O2mOi9ktqtCXYbSyfcfNZ5dhM81r/M5/hwNWZkZ0VQISshMU
IiUdtgNH1Q7YuoN+aH191CCFT9A1+h1gZ/9EtO7YBKdO86OA+hWvpEgO9swjiWvY7xjQH66L3DgA
zQaYrXGCw6/63bjGzATS2WnnfQqqFtpZiqMOEqzonwM4HYvJxRG8tqcvk5qJCssqve6zOFuZ5qil
kQsWR9bTU4MmD76FWy/zDFR3Tp6cRSUsJh7Q9HHMQeG+Muqvp8BpfC3/IjGjgzqt5t41UCvjGe7a
TjHorDs8Qsc89ixP4Ym/6HvI2/aI5Riqth4AP8TYQbB+YZFIPjfE7wFAsgLZRuCeqQ9VHhnTQDc8
be1xx1Qn4ASQuN7vC8073Jx7/hEWkiVpFVnJJj92y8JGQVgEPjCxW5Hg2oUnH1EFPqTD1TAPXZc2
FRYXGIErvYJ1fXWtHiNlmXgP6W0XROJT2QD9OEbqogsB4VdZgqecT4Hpx+nydUs5DyYGSNPG+vnV
sSGfnImGOVosAV7GW16pxmsapTeTNUZLeGgfE6YM7GVpmV3knG4uTsBY0d2HFNw/NS3e4ilm+4fQ
w5UN/3u3C5p1qMSau1GcuuIkVptfd/IDO4eS5TGAt4DebX1FqIOCFp/U8uM/pljxvqHlkvLyp6hn
w3q+YszycgwskUupSaZg4461gMtRvQLBdWBtYp4l3VLCSmVSLDepNSNOI/pXx1pPI6wwQgqNZ5Wr
QDNeUwjYVhl41mJzurx8YKDE2RNlVq/WBF5S5Cs1l60UT4ShQGb1timsYTvxOZBZzdougrHRlZwE
rudGg3R/SjW9h/6OMNYF6lbJciMX/Nzu6C6GIJM+j3jQBmPPMG7SHjFeFEtc8n3iTzviHKPX6bjq
r4n5w7npgCg2aJzWsA4LUJtboLT6J5wExX9gKtBSkKhf9LTCygaf0PkucZet4rb3hSotSOuya6Dq
iyMoNwJPr8YoouznMyvlpbxrGH8ePs5opb/d4DYygkcCM2b4HUt2BZR7/a2FE5yPQISvpeixhs2e
bD3N1Q6JE5W9dlAtVKrxJfTyLXlw+cP1IJG8cc1+ELt6B52dqKoC77+kHS3w9w308bxSza5wpZjw
h592xA13U3bv9wOBHMrI7n7N5l1kjSaP1oschyvg3UUtjqT8OQ+YYTSSIjgZe4TCA2Xs0LsgqkyJ
42liNhPVC98U+YNLvLhNt7B9m4ym3Ibeu+EIq4tsaNgRZqRCDujsFBCrFSdWwIa1T+eOmasmJN9N
mMfQLIpYI/QoT09TLVa1dFwKEgIcVq/hmh6symjgHMW4b6ndwVpchklBbJGzS0xB+I2ejqe1XYGR
hXMnBoTatOWw0CEavQsw3KvkBbVAXJ/NgujO/jXKdpkXMytOwqmsKi7NcPci+0nvhz13gvHThhiN
QWK8uB2jNxWCA6Ja4Ps/xnRqeAPMq/LZUhMEHKe8gjZB9+i3oxAm/oaqQgsJkySd1uxhV+nhvp8J
ahymFcPWjJ2Pj5aPbQjqboJME5JgHIDcpj6Vk40f5kb16tfFJzUbU+MsFShV6HuAFGWb1rpLcw5a
hMiN/Au5ZMswLwQeHvWkUzA95EWqtF4Pcfo24rLIZuGWNEUjWzTLItD6q/JhNBdFNQp82GIdiNnR
yLA2L43LojkhZdth4EP6iPqetP65ySB/5d/2K+cj6wKPaeS2KPTcpamwXSyRREvugAF1k0XXCQER
FTT+YZaHJk/2TN/i2d/67K2sVyJUaaaSNFAH8C2WWNEp0lw/G2ujzImG1UPCGEE6wRYvDiY18Ag+
rWS9+kAYVvkS54kjrabf8zyAw7vmU2JQ3XP1g1s4JwkhK6uHLCdvkhUSvvp0pvoFPH8s9Shq+RuH
+G1Rc/H8Cc7Rv/t6u0390ySR42RV6XG+ycy5jjlBxUOUos/OIVQdoQksP6WX8Fzoer6+LxyQO7nU
UHP2ZK5wAsUptI+HRpg3vS4kbaEE8GCyhCv2SyHE8bMc4ZOcwElYVNm8TcqaH81rv3l1Yud2r4tc
EN/Ib1R9Zq+l5I6Ek3+dcaoRYQeR+iCgWTcS8sYz1xR6TCNmvaNwja7DUeAK7FQ145UtS59GLSIs
l07Jl6hczai5Y9jkemFFn7DS67QF02hbtoiXONZO7Ywn/bmUfBo0RnLedne7DLz5/CNBu+/g2Em3
o0SqlAQUNrUJeTbq6VFsvz3uXonRy6Mh8amuWUNCSAFUD/rZsAGwII0+vGzbGGjJ+tQ5ywaChc26
0hKfKLXROS47pZkgux1LGHxxKgXhA7Qw/vBIEgQ+kI634/LSDJHAaRJrjGXUzpZhHFgQjhH/gsST
rtuyeTcIhCLV56F1c5OomIqvTC4xOwCRycLtkosaPA7IdIDTnR6rVNjB0pYl+oLtpXg2+bBF12Bh
6TvM3KwGsZpEfcQjO0sd6R1Qwz2/oVw+dJ8/izxLIyB8mDd2iRRzkoa2MubMgLfY7id7K3pzkdiX
FkFOTZN+u8wVs+pdXLK9kKULgAgQMF2rlFLvvtnmPo6yf/TYjGXjOAX1JbBpoahj6DNqRZXaKAbY
tetxsYjKFGWZiEeIe6sze+cY42JVwbXjVQzi3fINEq/6Edcy5NpE/zH1dxHmFMBarE5EJ4SucfmL
fOs4d+4dJhIWX+Ez/xanwmHyLNs4JB1V0AZnOVq7Zz3w7+KEEYcgtVWdUKVJ2GhY/or6Fmn8VXAP
CUPnGz1ALHrcmiNsDK66XmGnA5CrrgLAK0fAJIMJdXMgD175uq6QeDJNXS9uLgzN2k8O0BgtOB/u
oRrmfHtOzlpMn5GQPjpTrLbHI1/qW0aqz6yK7JT0vfazx2ZHpDYO3yRqou/UQBEGjhIE/4MIb86b
P/OFsu66XNXa97Cvzx98rFCAMMrdsr77+1tPRynixhomouTQm/v4A8xjMbrNScNBpaVrJRCxLgaf
B2DZm/u2XrfEI3rrk9s7Mne310IbaUDtQkvSuH8WwqGVlsOps2uO1WsoiQKJk0ci0p/FGX02E2GZ
5ik3rv9wuEUm0oiswRlDoAv3tWSDoKS28bPlVdpxW8TyYlxGVGzwolER+Fo+XPlI03HnLQBJNKsB
zfkZY4a0TVsSFDnT81WcMECpgbZ4kQEd1FnxJglDVjCSEgGoY/WTq3V5nKJW2k4/ot5SoqbqeVUf
jfgxSWERPEXHn9NGbF7qX3/v8jiLiZdcQfoOKMOnUhJ/mxTIwkBhG6U8OPbgq9M5klw0vVfdcdYi
YHyMfJBvNbvEwpbEMpA5wgwSmv/N/KD4tztJpRbP3qw/JDOcdIxCpESoS51ALshypwOPJ8B7BzJM
/d+kekhTfFCCq8PEmyN4dZRSdWTlUq7ytAHo6+OETwlwb9XqfQ7jkA5Nx3qRR/taqM64iIZhQ3cp
fWBpQ1pTsK1oq7kPfSPBWul9XFctQIIBTBkskcdAItPaLDX4EmYGe7kHMiYc3T6c9ukjCjMxO+3K
73WSoq9YBH9dRPcXz/9nZbljxcfVVZKc9h+y5meodD23k8iqEV+wePPE2zJ3vwEQLlVGtqBvdMDH
pevrRsf40ISkI06/6pUN6kfCZvxmNc/nUPAmKuSuQ8/JSRUrDDd/tmLDWkA6XmnpG53asCwME0R+
f0Rb7nSvsyajDf+TqaA2fdpv+EBpPptnxc5oBzvqskpprVVjgVbpGUGMbSSNyjd1VlIItslaf5B2
F/s+wQcoONmR0w+XYqVjLrg+QJL2w+3J++vTbK+5MNjY7apUkTtCxcX/+V+6ao8oZKQVPMOeRx+h
8AOL1DeRp95VkZFQQAUkj+lLsRPrWml6QS7uGVzDa23WvDoaQLdw/7OR0Cv+hR0uh4lslYGD2tIO
x1D1NGozL4ONa2+o8cVTEI6gODXWf+7wEdShdP9Mx/bSKZHwAW8+rUIjCfbD9tfDyw5k1pYHBRbL
YxMA7FTbXUxvzwnT1TSnr6Sd1pn8VBlK7NnU89Hc7ijvgEcKMAntUp15721jcHmMNNoZCCYBCDYJ
+n26PrThLMWDqOwmb+Uxcsfko5Kr5OKi0nnTJMN4k/qGXX3kjoaDSFoZ/m4gRlVgINkUM2+8roYu
lhViujjYwNsF7L3XBCrGQq7CBOBTO0zubbb6P2Lu7b6kShGnTjMO+FjeVZqZ7FIIZ7/d7v6gEASW
Hc1el638+6BaBb/fuc8YFKPyhwjBdX+d3EidsYi+YoSliCM2OhXZbiIGfrBvyKA9QczDu/i1Jcan
0cg60dvROYWqLTtD32KLh7ZOlIu51t+a1N6Sm5LnPopqZQzCIIHSwBlZbZPvTU8KGipUqoixUn+o
XEcklCIX5k92PKpdvN6x15VUNpxmhDBxactKsXGf9qmKQTeUEX/7TYAnHl2CIeNJs9FMYx2tnYJV
gECzAnYvGhnWnLLFRjO04vQ6x6ndhrpUtZvzJYiwrIIf0MilvgqyxkegJ/Y4vT1UE2gR6C/izGGL
aaLBe9VuVip+sK2jiILj8vESn7bFcSU4EJi4xAvgSryGROVlh8nr00CfJRVUrC2m0WcNxA+D4k99
l7nXuPuvw8ByTeigsYrwkhihljUqV6Yly0Dpn8+TQTBGnuvzRYKucmYA88LRjcQQggB2niBJTaoG
zaWeLxT3uHZlCk2Bjhej4I1a+15QCVU++cTndWlAAWmGeYlf7s8cNGf8aWNReREnF5mhu5qx//0J
Fni07+SMLv53CytzxCEitqRuyBjkvoNvuPD3meYH30fPFhSW9jmtx8SubiSB9cjezDTR1SJcjA83
e3dBT4PXmL5raWH+R7Mdkk3Fkrw23YBgHl9SnhK/K347jzzs4W5VawDGti1c3/8/7StM0rEptyW7
156iPQLh0KgJxvX2GWZrwhhkcsipRbcqmKT+Oy9lwTGrRJ4oM2YWX3DdDP2nbrv20Dz8I4zOtAWx
RHPREPGUBcNj1nfhOvZnVaKCdECVFNjssC6tyq9ZWZjxO3qMOP6WzIQ//Ehxop/FWcKsK8Ad9ex2
EGBskntU4rgAnwx3hJkznIB1BMGsnlyeYqAjIZVdoRvLay8aMcYELhFYlP9WmPFcdMxL+6zqFmGL
yjotjfjIt4z5BG9zp8C6dFddp7+R1gJP0RL9nKk1n2eE8LdXsaSqlRa5BNF7CsgLyYEcn0dhpJ4B
/fsNfsy2kqaW3hd8K7X+FdAQSsopCu8v34SIwMOjO0HC50J/JyFuuvwju6riODHkmRDLa5fLAGwx
L8Ps1O/vp2Q5vaFuB/e3BnxqFw5gQpgXx+awnR5S5ZjZQKyekh2zr0oBcuMElzj2QTzTnQqWBg37
Bgw9t0qO/z80iGZdTuj3UBs357Qe7jO3MNUSK/WuQ11Q+iSe27vNdpMvv8C+Af9rWvLcMA1Hh0Oq
Dr5Wo6J2J93s8W9zBr0SR8BpO42ZmAZcXdKKfIZbLca8rrrDj470yGnony+A/twgy6wjgmJG9Cus
qIzNwxdfb9VBhra/N10Mp05t1AxcjSsGCte2jL/woME1+BeCbsqjE9R08eJCCDiWEXthBf5XpnF9
r2iq3X9nAFdhsg8cYGNEg//VMbW1R+laVNhIvyH8pObv4iZVW1r9bHb9VV7Ug7i9P35dyRtvSYSk
kSnx/NUnCa+1bk038ZvgNzfXO63FYCSkjCL13fYMnASDdasiEJuhRJJskkqGt0OCckKG0aEw9IuU
nCDqXdQeTpZOgLzc2B+WIbKvgWd0pikzLNaA8LSXmeegoGHgJ4ceiBcXFBU+eqMk/DOLpj4G0ggD
LvAYtCr06YiLaNmgbeny8ftBDo5z+nySq5ee8ZOA5kqoMvCBaXdLxRCchIRHLVT9PtH1aIv9cwfF
ZSYy+UqsDs/eZ8JpAZZ4mYw2w7CRUI3kOjp2xmEq3mY0HDdlfSN3rjoQUSDLza4BSHt2gQsWtt3h
fTzY5BYMuugyQpQNWVrHewLBV79xcvWjw+J0x+u7kl4kI00H022JFMjqYt9/lwRE23qpZw4WzMuY
zCCyCxYmbfD2R25ge78551asEv79G/2h7WPPpxFkrmoPBmfZl9IH6efVfUevosbr2GJ9oplT+l4u
kITQhwteJUQdqcer6UH6Ldpg5yAeCkZNcd1tzNwHN18CyMt2Cie3wn06/1HANVTRQP7PFSrbUbDe
v+bFIODoh+zBoSWfIhBfUT5b4WgGwXR6TUmjlDIMYYnEJx3g7ohhDscaZu/JtgTPsxyQlXRjlHrj
LA3cc68U8IQPcTpNsXIt7MnxYkqVjJinMidabYVJ5ci6Q1dtBI9AwWzB0IncZEMrWnapnwdlPY3Q
Mw9C+TMplz8nqPdaNKG1u6aX41vZjLwcMcUe7u9OsNyB1zfmtttSIefACggBGOW9mgJ3zHq5FYCr
5qKlhxgerJGp/4pS+Vnt9h0Jrt+mr0Yyswpqvc/AbcJssWEGiq9PZHgc7C6odwJ87sRLwCcsKfrr
ElRtLpe+CP3LKfpVzkqbSwkyjwSrxLyHMf4/Lmx4aKKbnTAyqf52dg98pN44/ACNUmrawMcvZypc
71zZBy+xil/r22ydiT4n/m7aKuOF0kdrEamHm+l2cuXUsdicq1+pBTUAhb/UeItRgFrIAQI9ZvpI
IOqSzPKyu87ga+Axbz/eSsptMgoyNxCnE52+lFYPgOykH3Vs8aSn/DFKHaaWZILyhdm63SDyRcH/
x7iWCTXb//9I/OPJyfT87V823W5Cdre9mXtYJItRjta9OcwizamtVAL+7gRXiEqfo/YmSLeAdGW9
VNBgYqIm7HIbwSOAjwjH7fSRzys36MD2c/3ma6mbX9P+w35QLPOPpt3qqJ2+W8/ZNQANskWFztOa
9Fb7duxgvbif8pZytkrpkJqUBXRyu1cvF8ms6Pqgarmcsk1vp9Fvqfg9N6bEDeX0kOVF0knVhWot
/x6qTCoX5XAUKjjxAfZkxecrQLF3Ylo9d/DwfMEtUj58sDwDbXUaac2W26EmpUD/B7FcoOuBtKAO
u2G8cH0rr27tM6qgh24zOzUftLWsWHTAtw8ozT2G8z6OW6VlC9GBPCnglz/Q58lKQN9kq6iIsp1h
En0dyd4F/501c/ElXSNX3Bbx/2U7bjO00cAI+2J/9SjukMu5uH7K0ltnSw9AEZhrTN5HjleB0rT+
8BY1PB2ux5T57LGkQ2YjrzdVpYblIsD4ftmkdtja04IBIEtXSEE1pYqPfrlqf6U/We4GF53pAYRw
93JuRCMCcx5B2WOUWBu0Q+M3AFdfi+fePe3ZZuPiMi/boHIh7aqoqFqFwNlJnG9hKSQcEI/AUMHU
aRwSUrAlgYvtPcRQ+NqEUVSLEOohB7DBFZf6Qh6ERBFm6hdQjBLGf3qOXSAq1wcSl6lVYkGMg0I3
T34KjNQE7n8kseqxVaQAO5QNEXTkhgjWjDImQr8hdzcIVLXzuq4nUa8KYc3i2IhHwMHoaQKbN/FG
/PNIjXs5f6PZZtvESGp6DwYR8Hx/IPbwIc02R5lDmOh/KQeH7BA+X8OO4SqaX8GlnyOv8aRE7PfH
XrqC/KwwymPDUNRd0Aa4pNlnz9ckCW6A3S2PppciUInphe+J4MiwYZ5pnttyX2aRdCQg+31eIsPW
PJavvugBCdtOJq198O2GQcGWTNYGE2WgPzjcbzVFd/FIBBwOKOOw/p6lcQik81SEgXkKZ3o3fT+9
I7OlB2dO0CV9oSY3HjGP0R9iu/L9+qWEs55eJLaAvl4zTrghNuzBoHXfJuipDXU6Dqwh9Y/DrOFi
hztWSbpbMpLRNxSwxEB96xgwtaTng1gnU5bWpCiV6QFIyxdplYCyYfdjhNAPISHcvBLTz6hBgEdn
RB+BKzuukr3Iu6mCqj/JkgO4PPW3zP85J5wJCmcjvEGMb7ETlCa1o1vpy28KtUG07zcYXgb8oFbP
0BD598+dYwRZCOzjLxSNX4hC72LX4XKRszmEVZA4ay6zCoFx4y9HXxHgmGuAW+IXxv1dDDeXhIME
28lnKsshAmoo2bvd1lhlue5upq2hpg2i5Yk9A9NZepY7pdIQvI7OxZ+IECrzc7AaUJ16Yb3J78HK
Se3Y03oW9ZJ9uA1vtPX5yv4fLN/XWrx99/LY4tfO11pxTwMCdi9/BtJglX+p2vxs/mMISE++FEGq
83nSXq8qIazXPZ1mgvl1dgysk9WrjmcdkCxuMVp9KkfUodckG+Xnn3MynWu1IAVjY2tuG7F7yhGw
E3p1Ay4f4oAxc5vCFmG9W+pxD9eC8qw7Rd6Zrr7MHHt1HdrpRux4wu7MdMbjXSLzaa54pm+B2lW5
qaWvXILkEbxboJxg68K5wOCwaHU9y0sWa6DFSyqzyJB1C46zylu35dzFddr7wGlIs8cfKXLQdsUX
bRnWMMZAqRB6UGXaXqoTWYti+PR7kx9NvnA5yjPA+ZFyUG1MWplQNTvJzeqLJWV2dADP6rS0+AGr
gVHXl+gbzc8mJV/a9F/BVtZ2SKWhz06dAFoCAr1Vz1Y3RGEHO1M69Fifa+DV5V4LwVVX7lxAJGC6
k4eOuxgr7KTnUFjWPDv+VRGD9Ck6urx07hNJDBG0aco1iP6JVFipmXJ4OxEXit92zDaPcr+VknWP
eISQvuFZE/tzYed8hd2/VM9MNOBBtKrfSaCOOsjtsGEuOIl3YaJvN335X9LXus9cRrWcWUx8hSJz
PTWVdc796LXVDKmB7HjquvrwKtdcG6LFs9vWJJAFFW1Sj6D0/b9w4aEA2HSSUcduasb99jT47FeM
v55NwRotdyKuE5OSTWUFhju/g5zV700m99PZLyrX9OnvWg97khssvocxLlrpD5gQqSW9ngU3qvkM
rixb4GMczDIjBEc/Kv0pvdcwsB4mAgCYxYjZ9i1npdM6CNh/7Y8tD3a2AnMUNdPHkgNL9G8dVnPl
wrm4qOTG4Lc79JUKk70J9dV/uWjeNUyMrGDKrn540bGxKUFKzbxVLnNqndjrQKNNEQzVvqtBmrEk
llrqAMDcYPuf1PsQMWdkGRyhb/WexB//s1T3MYCYh05aZIRsc7QMl7WFH3zNORTCxoxkZQ1eU3uw
ttpq6u3K42G6kgaSaN0aKrJQrT+PQ+ArRLQwpCcRLWBcy9uNOoMJp/vrH275Pg62U+Re/rTQ9ZG/
sLz0TxytaPUu262aBK/BDZccTFgA/8rTylPTb1GIZ71Eif0o0X5hoiHf4nOLCt6D+9hgHBQjnqDr
krAMfiYjwBsn8n40QEOzCXEwJ9VGlshAg04gYEjR4r61g/AIOSb8gu9pPITHsq0O2raqggP9y9DN
e9bc/BQwpBZATnwf34SuXgQioz11eBeAAJAFoTv76ymj9WdFTTv9SDSbROVNztc3Li4C/pUnLH8i
xTZdP5JAF7ww5R4anF940Xv3m7qKTqNtbRSqoOS1DOgbUbVCtKsy2O6hThw490OBi6csjSdaaLa7
q2QL8PuNTrer15h0UbwRxA/Ys351yFVZsE61oJ6EoNfKLx2hmfwIzuZWC6Bw/2On6GNZy3m232Pz
pemtENAN3wZz8oQb2oQcUXs/ejLni7/d8bSMsEHVJyWWEyYNNRhhSR3QkXKC1IuK0WEou9MUooEc
kjEwKWNXzQIzGhtbwlnCBmt1ArxhbgTCpUJne7ln+UxlY66gIusNG/JsjP7I4xHq3rmM63WtyUWd
Z/d+hWTMjEgUn7AjnuOrX/MyL51Q+Dmh7mVRGMeuJ5sHYQ5vEroPpvOAAeZiKycXesimhyRNHSWa
dHUNeiGrNR2Vp54FH2XPMzmfbjDraN1lC/UJ/7vaJ0mamb6+z3dDAkIdKFNKQDV9McpmMZdAHuMH
IGCh+0AUY3Qr0/p/rhRM0JEVSXydZ7rpvHoRZetVDtXmWIEgx0QVdVZrT7WFiXbHvujCYfIcbcZZ
rRlfg92HWSqkS7cShbhcFF8gcNqeVF81O+EVUiUjqvjKmSPw+rogZgDS8IEFqW84K9lN2xGby7X0
GHbahxA3NT5Zvq9HL6VfzFE4TrUVRXi/QXiluavblMFfE5sDWMsrE/djKzfCrvW6g+WSHvdvIaQh
89uDNLlHbJLCK8juNNisrHnbTDze2AdzwTbp2LCSQtnPKtUmVuhX2KfYJVD3wEHI3bJTorKYaItp
cLgBUm3uAs+GjB6fLZW1riN9kaCG33tso+2p9E7JVysOdTPQSaszSct+yNVBZOPsNWrQ8Cmloa0h
9x0Ks7aPKpg7Z+DxLVQJCgqLh0uZGeAI0IUOB67Ja/NJbN2uczZy2WHv1nOrbhlvxDhplrMrtSdf
PaeO68N3ofQeOgDiJjX3KuWwJ4eZRCarKQEcgbSZ5SxAuCye7wMw8n4DX+J1uq39jRanmsqdRnXx
yr82uv9h3gn8gZ9qoZIM6rupxW+x9lgQSzyT6Y3RROVlqdD7MZQxVeGJ0watWPHRHdFDZ9XkVvV4
EsXXpU6inEuhJfVLLu472abg6A63bAAw+S+f29mxglVb6zRrrA/0KF1sPeiXphNiq7rwfPFrpST2
X+8HYXK6oNGWoMi5PUC2IFdnVND/eNoYagB5IujBVVqVltmP+07Yqn37PmyUFaiZJIJMtqyXY5RW
5h9pPJs6qd+l1Kk/nczrG7LLNcLzvuAbX7eFXzbzbGbQDyTZBSqxud/Ci099u17IyxmOaSwc6kof
bw3GqLToBymeRlawMHcANxliKVYNvaKeIiiCkbQ2UQ9sJ/zf/yMmWRwxVWd1tZkwvgtk+2jF+ZtV
F6mqhQjGoRaqrEADPbn/HvAoi7nWUsGqDeUhaWFMNQ7GSlpNB5LDAT+rdHBPdFQi1XImnoQuM2jm
ACcJWq7CsbHlzizc0nEAIdR0woEd5O5AWY3+F44Z1m3y+cA9VSTno/xGlfzZbFpRBd1csHzaI5oE
5tTQbgtSIX3Du9K8BCYcXtUB3nE3psvC2BuuU3277dGshpRzkIbZosRBbP8zXuGNSBX5ONBjO/i/
zp9KPfpHDzWzoHao0O+A3oh5xiMk3sUSjyOUfG05pTPNG1T19mwCGYw1oJ4g4K3D+OTQ94TVALLd
p++L7Idk67Is3vS/6e7AHaDblAddQyoqiOsedglq+F9Ludu0nYAv6EDftrQkFBikY+galiQMDm67
2V+y1C1LGnWvBLim8OSRp0mNSCpHZHcZfMSqp93hNgo/KyTk4lR+LxGVuHsPEqsNQu3m2+AQlVbg
DY2ZQOLNvv25usAyCxZIeOy7W8s+CyrYDnvUDcNm1t05Bx1Ii5GCpny1yYIS+LLYSiH4CPUYB0FH
A6zMKIAKc/hPmhioM5Xy2aQq89YN9CHE1xqp9EyG2DjmfcIShE8fB+7bJLKhpq56bZJij8yJxIHh
6ewRBXXwezuvRZFsIKCrrwSj1ZjKr9d9Wt8WWgd0V+DrDwjlGy7WfuLTfs4G0z0xYN7MqpCpAZFK
xr/P57GtAwVrf6CouikNF4Op6tjr8OZ+mloFA5xH2UGgSX6PeFSSjcYD34PvdV6QAyK4aJgu7og5
46qgNSE4+2xbHPUC4xMaKKmiHg1bU8wNCzHM395wnl9ln/6ttRelVN8g8MnrHbZ9MekbB+qIC7bK
e360sKmKrxQb8WHrcX/xCJUnmBwj6QKBU+rr4Cqfxee/7wDbFTa4R7FyEhkWmBLnq+tkCaAleu5S
ceOcJO4/zLbwlcxrnfiWUrYvMTCvsWyT4YcffHLsJV/c8eLZQ5jXUdXLl0lf3+WiGUYV1blXqzHT
2NIkdGmTUtj/GOVgW/Z6CAfszDN4yuOqJibBJCwz8upWMIGe55WmdaN+8isBJHSUbjr3PRkarYee
wHYZbdj89UVqg/56zp5GIPESg2Ll8QODUIikkY+jcYbU7KBpsyOmoMdFT1LcVFp5gwojXkWHMVfe
v51AFWP+e86N8Rc4lquWF8ZTZkqg44Hv6HlqgVAorbk3zqB7cgsT4PBULj5yMEi25GI+MJj11HjE
XPB9Hcff9D6CsPCNlO38oEYMTceBDjHfeQ7YCqEnTS+/80E2UmFaOqeU0Ezah0KzvRwuAt6aOsbg
9OjK2FxPc65RJYYnMRAAyPFueGjP1uZM3fYquulJ2YrdaBds90z940QYRiqdaKc6As1SArqUtLlP
6TQYNB8FfipnR71UDJS7Uo1qUehhA+GKvgyECAxfWkzjNzy9DeuidMoQrfgt0no5Zv0mrPOR/ojQ
r2g4ReIWj37IQO8+EcezeS+Ak1j2rYVO9ANzI+hC8X6Vk2XmzAwuP0gLqz37kcL9CSrL76ewIG8e
zYb16w2ldQcDbHkU4AKmtNdNXY+77FpNv2TBbPk9B+7uWFNxEW9J5nCKKR6nmmSU1aLMhwmnnSM2
I/iv2J0xM4N4CkyKl/KeTq/Ubji3Za5dwggQ6CF4ncqHTPD+9YFifqRXRSscRufhkUuNuk5X1vl9
PKPVEFl5P278V5YZ0L3LxVopgPcOXxsnhSR7K3TeVtjeCB+xw2f3E+wMCXFWFF+mLoJxI1sulEmc
l3GQzKWbTCyPrkUxu5nusqxEu3ViA4l6pkx5oVCxep8Dfhp1Ri+1FQ9Ehd8cMhcZSXwi6HuoDjAg
W83eKSanwFKMLbN1NRoRcDuJiGnLB62o4oAJ4l84dmUGsHUnhd0F0RgissD2DzeV2msdc5vBEWgm
Fdu+ihBWyDeeAw2ArfKV9uFHwGe6gZZjen+jZqK++awR++uhb45eKd8p6g3ZHUYVpzGQotUJYYCb
cwZhTOyyhZRFum3+htYg4xQDzVWEInJWg7aXy63Mh2V2bQodIeJ8TOBSJBTI5OV+RS8yAzvGDtNJ
4Kg9O/+9EJGgNoMRj1RdYCEc1M//puGKhFtAMi9pgaPUxAASrtWQLD+rwZQ8yHOPdspZcIYJr2F3
65LMTSs7QLv72S8bSfeqg/odFjQTJNQvbG6y3PqP2lCpyujvsjx2vv9Ec8ovGPuEqF1AIni2w1Xh
GJ1eXoXIZNyHShDtof+7paVK8TBcSaEHUObYxflAZwwAheFDCOeEnHu575ROd+vFmps1TP+A+BCG
Cti6XMGLrJyzjy2BauqTcVWL3Ox8PTDzjnZ2vET4F7Mn05HGeLN9H8YfMfz6hNP+QLmum5xtO0my
QrebiRsBpm+uqyh7R6I/XMMG1RhGL+P8zJnjUDDzyJi8imzNVZMQOiWksa1aJm9s5hTeqxN1Fd23
88bql3IYiwnwx6vSYzCZ2VYe+xNyRqk7+abJl9wgx2ceQy2S8Laqndwt5O9Py0wFfc/xhbEPJ6qI
Dv+TcBdIRoJsCY+3xsg2PIyQ99iBqZ8TuWl25erSKhdow+3BLiQR9expD+6TKwrcvnJGjLrPDvI3
/8BU9ggaGH2ocx6pic66YDRU0ctFHJreXBNFO3YOYlDxC8dWAEDzBmyq28vBKiaUTCCY5KF/NI9l
2y5Taqdn2OouO42Pf/XLqpNM2OZT0xN+kD1vmoQo0aNSm8BxmeSR6N5NUe1fUk55sL2zLNvi2hh0
skRmVBs+2zx/32sFvbebjHSKGf2an/0oKOsr0LeB+yJpRsvEYMj19jYcUPUmZg6vyrzsE4NP49QA
w4pclmanqDvqRdd3jJvcUn+1ZIuk9UIcfD2yg5PBVE3pyH8oUGb6/YUjww6SphO96y12uqeHIkVE
5t7lO8XmaYjlWW2DocqMB7JfVKZx2LEwcGxG22vR6usBxMzT0qfvJu8VsSYBOuUJCvvdjoTjixqv
4vUXcSCs+GHclIUtPwRgI9Egkuo/HjJxpInGUb6NXc6pLa0s6qXE0uYF5H9Ywhb6gvUioWFtfJoZ
DWA27tK9sAf0F9smtXdqWceVlh+ckGgaOeAaavyrVnaUXbBgnnOTZxN0YrO7OyzgyjYAEhZLtvhp
261ktslZFHKzUnl/+BWbba2gG20dZRSAN8VzcIIBhIy0IxoEHbFttJbIFSn9vAgdwcLEYn5mjaKT
nnujF/OPsJIe5SSDpBQbaF1bbbcILV/6K3W9qAaT7u7JQAWQE6H9mUouUG1M9ns3T2UK0gellIfJ
o3iBZDbwI9vuTtb8SueWbtS5jGm9h0IZPIRH1a5Ef8y8aBVvOvNBhvhm8wN+B5CmCuK8dVEprtiP
pl+KodLbj247dShMH1GAggMlNr71hC7S78d+vuYP5oKRSDwvC0Er/ik6/mASaB+f9Hs2D8P31/YE
YKtQxdZns+j1dql1SL9M2l4mXn0K+ajL5byqI1J1vBAdBznGhw7v+G5tQC6j6ua8jYmiZIo6kcTZ
P+M/Ia26b8/iLi6/EcS4yjMPW1/h6O6gjV9NjXYLeWkI5ATdN/Llb0bO02MuIaO8ACGw4xGVygXK
rWKLLQfjIKvFYvkbqO304b33hxHoaFmkXcNOXbGBHWyPtL8j7hJHzg3oPMk7aB61mHjj1aYB14me
8mOUGQo6v4KsoNUAZ7jPiqYYLMYHnp9SF1LoBoPJzIvE/strvZ0GSVDv+WYyUqyJAASxqooDAr1o
wwmH6AbbnjeGWH2KkV8S/yTT6tQrflKlAJaMMmJmt7XdCO5U3HQ5DCRGFM4tN+VrRv5IYb7QKAjq
rsrNXP/A0z0irBUYwthxqzDAAVld2iVWO8SJj1n8q5OYotL8nADiWfKOfbTeXfachbyB/UAtESNQ
7vNOIicoMQJZ5cVt0zXnft6Xk24OuEoD/1sIj+ipQDLyYji3DJTPQBuxfIeZhbfkpAZg7eAIwCEe
cKyoOTTkpQF89pse4PpJKWqnmNVRReSa7/V5PlT5o7x6Gm0CC5pZW2ltYdGDnahLBjVdCBa4i90f
/k0losUGhYtziamfHNRIujjmr21lRg/Zb27V/RMbk+5gYyfAuvl/BGAsLAn6WfRViCPvLDRzD1yw
0Q4sMdfHi9z6S6Ka9oZgoxVX0wmZyN1kTYlDuiKkyl5tSpFC5pHa5Z00YExAox5uyL63YpJLlaGF
umvGuQkZ0fBGsrSGT809dEObFpWa4VO0RxhpxAhocwxOnl9c5JeUaIsLVH7TXZkz+e0JXnIMh5nL
Vi2d+Lv+Dqo4Dw/fJbFv8gginTaishhQW5bVP4gWZvo4P70J8gu+6VmD8dpA6pqGsU3TuqjLZ2uP
NM2CMMQXmX8LZmlXbfh+CLFLXbUCft2vDt4JD0ss6xnbluxUxYMz0CKrrGID5qim1BuoBKLKd7UC
DdQlKN38Y0g4yLBotYcTqL8a50dH+vCZ9sXoYuUEx3yovCX368zfDp263ZRn5wjDlsNK3TOjiOCp
qOwXl0rPx5Jb0N7X0GYdDMUlK2mVa0wk6TyshBqj1Fyy/VI6dXsgWrM8wz0XkvYU7yxta/4euiUA
Z3PWTQYjT1q5HFKv6QEh4IRX/tiaTN3+tN3X8AhUO99Jvb8lsjDZxLCvt+eDDp6E1wNUv+F155Hv
ETK2vFAOnZKF5weiN9AKx0hPd3sVL7F1qox0cO1T+2OWz/WCy0myLV56VjnIE/bU51cqv7jkHkef
KsJhKDRTSovteVD3GYwlz1zfNFmbktulrijvs51+lrFy4bRBR9YHeJCeYZc5siGeqY/P7VcxrwS0
wzNiGAL8A1QytYhplwFLucwDKGssLCurmT5WlhcN8FePHIipn8rSjMtSBatqMoY7MsgpTHlD1WuW
LcUZG93F7VmXtcV2bPlfEdCS5ZEj1Biyg2jW3VV2WN8hpq24GCZm2zdPtFktxLPWnwccpkiHzL62
s6bZUWvJ0M0lH++EinbCyEDhK84H0ZI0WEWqjJ5mAYoXWHbVMfbsvryUtuVHzrXMOsyxpB9VPYYa
0mezP0GO98KdCgbFA+ChA3oQ9FQUyoQ4iBei59s/t8Gr0iwf3u58aqvcbcA/ZsFoHC2fpm+ccJKi
glfP364nh2AKZC+uj7Yn3XZYPfdJdKxadzvz1aOcL4mQG+E/eKkaDLxdgBaI2JXuutVF85g8F4+8
gPFbckpqjiJSPB1FiCAETLBr708tC+hUm9eZ2m09XCdwpwb8BGJXuZp+rvYmMjwQfWGi+EONPay/
parwWHZh7DxJsgLkrmwILFPbg4rEeAQoPJOEBRnB49vqsD6yTeXygX5lGwqsOVo0zCdHpY9V99jy
znhUnX4GWhQhFrEb7MjERsrZes9JGZtcw1cYbJLCHp6qoDVHt1BJqlgGtcPvsuOXrF0HPmg+JwFT
7pvLPd2wzdTsgUk+c6HjQSB0XHHTf7hMn7bl94RwnVMCeRocca4FrYfM7EBMzWbmaawtsKqa4bLo
b3epQLYBowN5LgAct2dFMuKb7W2k2jwYkiLNeTyeUbrl85vrOadizLFa3fd9pEcc0/rwNzUUa1N8
lgIeSiU6ygaRpew/SlI3dKUfZ6aOuUAnwzeFQAfTyyPJPiCVWFcxMeFApfzjf/nVzFZqkMX5GbHy
iTnXZYz5gDDtSoHpHL/9F8kgd09qqZzwxZkeVfuZeEWTqsRPeqEKg0RsiZcY0lZsMEPMU3Qwwp8r
OsY0Tddh/mZ72YBjL9UtthQ/TwWwJu4pHxmaV+etKX6tJNfsE0ozedF7yososhjDv1FsZtq9Kwxw
Dm57AnIazu16FQnhJptHF2E9vv3jh66sFbwEZC+iqMZJoYJDJzrHc1ujBdtu7RvhNRHaFPNq3Vgk
pEmpnCIEFEfoAHWyftmCeYbKL3HlgoEa0NL8sS1FKbKK0qY8c4gYGID1xgdlxBjEuPoRZgwKPj09
aqXygMtVNyg6mf78kbxtF0yTiipNLJ/N/2ZETtzilgsoXbmSf2Ocgnu5TBcm8ydHBge76IjtyO/V
TKOELzcrhy+GY8AsaKoXijcnGTpgpICBuJtBqBPdShZ9Nha+BgI8yH3Vuwt/2l4g+egCN5Oqx9X8
S0RXWExZwXmj4KYTT7+vjPIYxoqqHR7YfHlPoxVk/WfDarkn/pEvPpPbUWfbT6SNnZhRNkS3/kxL
eDpnvU33tC/NsM7f3/7hTBqRv5KOS2Dv2dLTg8qpcHNSre2UoEHaUnUnq4ayPc85P32RMuqlsg4S
AwwugneaFQRhQOX1dvEdK+rxkHKvG3hTX2Q/UX4cLC9RgMsgqNT7Tf3m9C/dkcWC9znJGiu1DOSS
zBe6FXg66ve4uwRWzOlIXNbnaXstw5/ynqP4XZENNn9UsQtin//DBQCAenk/8GuuvdwdZdynolXR
0G7fRmGyeGQZ2+s11D5HsBdUthjqnNH8wT6NIjwydTpabr1HbJeJOf8oc1V+Nt31V77iP/Xm6m/5
lRAIgtGUmQdJCdA9GGgJBCX56zg6PVaNnLBUo6yO6gAhXvhGQ/QhpvxdqbGXneoY53O1ijjPtD33
mkryvNnNXGy1JETC9palbU9IsEKkDGg7CYxJgMJORSsmlaplzLa7iWGliJXvWCKME0gpHYphNQsR
omaXESN8uRloy2lYMG+/upe0hNB2Q6UY3fD3ocFqnvrlZYks1b8wvZQYb++LQkbHZU+7rROa/+vg
r57egQnOZfqoxHPOyjdEtyIIbyaXqr7NJb9Xf1kgMYX+oNdHP1Du4D+aXYNOWPwQ6OmFmXUT5AV8
ypZfGLx03mbuMGir2q/iob7lRg/9Qnuw1di33BbT3znwb6zVf+CfZ488J5MwVe5qY2UmUTvaYU6n
PUtKzLnrfng+ZNkaYbQj1I+D1fIMYD20Gt1/q72kW10338Njb3boKOZPYncBm75RGijws8fUHhiA
uRI9wL9ww3eE6OsJbreBfhzZrkFcGpza+boN13E9C3sQWN23z5KxZyzeCBEstsCUy06kg2IvaiXn
2oEjeF9bKFR1tb0gIbmld72ouaOXa/N4ub7n0cyvdojj2l73K8SHOuIaU3pgbkBq8NCfnq/CdCqx
E8gC7ivP1QKmQHgfao+o+XvBqlodM0q428P4TZUgjQ+J2DXCsCFuUnxkj9WBe4hcByt7qDPy67Xo
L7uMgj2YiTM+DmM1uWvKL5PZ3RIhY3IvEc6acy7VxKgrHpqHtE53PtWYlTijcHKzeWbEx8yA+Ntt
MXBa3KYbWjOE25dtesm6L/jBHVlGqHS4WvtV1vSrzS5k9oYLErqYvwr2BBtkmVrYdB0C4wk3yFEP
D26DczdptjSOIr0Ix4MgmYQ3+CjZVKCa/NOrk8qDKYoP5DynWEEkzIeu9rNg5J9TSJxjV7x6Snus
elZHpGNYQsvCMiwwLJelDK3ZgZTHRf07EfNn51kkgCVXfvmUhDgzQmw0WYxpQMOF3seAvnvR3JMX
tJOY6pkOzmtiGY8pmwUoxka4eFbqfPoi7V7fFMvykbAGRpa2DBabIW2XBn0CSDJlT+47RuQqK+f/
k7Zv+H+TJsfTCUMLWi8dP5fDDme9xyViVzWdBroHDuBzgFqolD2b3wl+VqpJ/g+8a+/0pp8fUTg6
HVIjUH44/AlgMjI3w/NxEogIYQ+/HwMclZGC13oKl8dIvuOr9LinO5R2oFRmYv9CfZGl2UylsCjs
Y0xOWMpmEdQY+xTQIykuO8rJPr4hV5iINbMAVQJgv25/aZRUx+krkyFWTYep+We6zm/LBpEKM/o/
2u40vPyF6rJGAgANG8NedJp7PgXHdYBbcG2UekhjMNVlbqSQlvNhbCrgXSXk71QeSsvR4Psh0Cd1
z4fvKJ26Q7iZ4tejkglvhp0pVF2AJ2dy4gWnSN+hEIFa0wEWlahHoG3dfYdzVYoCfVQkZFNrZzvA
vDD+nnNKmTjShHFzlIIH1V8FG8Gt+JIqWfO/bI9EuOgEkMwu+OhZ1H/fUMMlkQlcUvxl/hSchEDP
fCxbYqH7vTgC9/ZDpmUCcTl3kJeOxYqH7sskyLEBwRqAMR+gCS7QIMdlPChVhuvaUZ6JtPDNc3wg
ffNxF15QNb7+mTYuFxjTiAbPdurQVVyYJjXbf2zttu7D9sp/PsOveaCy2O0dr3XhCDNCC6IuTdT+
yhpIBotR6LZrqsnf0RRRzt3mTalKSi5XV/KcCNrutZOvxVj0mNUIh6fIX+181yzBoWvaui434J2z
qi0/dNyIk5dnc8UgxETsJU3BZGMrbWgdYF1C3gBh+t1LVkGSLzkYOEMmZ5efI8RQ+zbku/I5XiUz
KPwX1sE1JrFF5aap3pToPwSCO3byXpR5MqeZ0dMuU9PfD2gwl+9Xa2cgQEHrsmUnJ1fakrBq++uD
lGlb31UUaPKsa7YKzUrS4N/GNLSPZ60rqJDIR0oVFcF7HnszB6rKjvdG92l488tqwNDzUK3pVPBn
k7fLX961JydM1PN4HSV8cUN910qvBcKTtK+Mi+cWy7xHN22g3hhhf7XT6p7Hv672+yp2hQBN/ZNH
fLmIKgLTwDIyaHqf7G7pWzqgFscrfDuik4ixvqXeW/bv8gQcAI23AeOCdThKlYAAHkgojXIUELih
WlIJvlGMWNMU5xkdMIQtS7LsWZQxifPnL1KOa/UFOz0xAOnvWikv/B1O/PJTID6CvqJRn03WD1TK
VAL5Iv2rSv4fVyu/u/KOlPDv6VFlwKOUhy4GQhltcs3UFayk5d9k//LmI09mvOLt8wwXKkjkwE0Q
JxtPRZTTqgBFsu8Yt+Y0LKiM17A7cgcrvXe2shTHveBr2pFIfOzSO5Gg9G6OM0V3V4NBO5rEK8UW
DFwQUYgTi5579rTnRR/JKjEdgWmmEa1kdsPLgXXmL4JwcomWrpJBSRXHcrOlG90R5OvqoaBTfcZi
C/Wa77IkMG3zy4TIz6Gs6vfybMP6ICzmQG+6epDr8xj8SMw0cW5dhA3ztfEb3tlFMm8Jw8oL49HD
0aQ5K6gOq0bNszjdqzY/o8bwMtibij0vDabO8GA4TmQ6SD7VmGAK72/GbT/5g8tgGAFnvKLXdNZ+
Ui3sR06LowR1Gv9gxksY0k+vKq2qSUNBufka7GC6d5kftvtH/rCKTnHO9+K2TiHEqU4JfOdBWljb
aK9BamWdfzHCHhB1KrS4PTzGeTKwnv35dg/oK8nV+ev0cM9yZhrTkmjHSqtmRqg0ZeE55skes0mK
VXi+I8SHAqpGPkTQMV2CvX15nD6VeIvaey6Jm58YgppzrchC5Zs7gNjNPRi2G9Twfge+Jrnv8hHx
HBwbRm9X+WIfhs5ONp5OHcy4oETokX8WLZC5BTKoK2hBjy1nYB9E6UpzH7sVlfsh1oHjvLGXc7bM
HR1KQBUKBtX0++eonIPgDnTXs6YvJB/ZvnvreTSjcNfp+CWJb2kldl0ioSikGJ7Bzjb1YwvjgfvC
9Dp87PAyb7nrt91kAtwe5HlxziI72wkhi2HpYxTu6Cnvaxsx/9H/Y6UYL+TH7L5e1TG768TEF/DX
IsOtEt5BWm+mAP0ueX15iD10H1K2sZonVBzUuJ26anN0tlhd3TJPOyh2Vr8wHLOX5sS8siNMIO9w
Fsamf629QP3aFcPdeLTBlVB0O9lN2HjEVU5bGFR5bkXYKNGAjCbp019gZ/offDrPE9hYZMnFi2HO
nYof1TGW+BC7n50e5VLVnSml8X/CTKGSwYUv3pc2PrkKAO6Iwif5nIbqtjzD5g6yId+OgQxSO9+Z
7s89q93z/ovFxPVs0Vna5mPc3usTE9QzeMjfd+aM8XQlwqZ4nepEV4w4HatZXIMNOZhvQ4tqsDsG
fnvYGstrsnIUjpJMOjP/DSxrw0xpBe+B9mtUhtypl1CM2bt5ZvtL2whUP+LPnufOi/JoNSBU7sQV
th3ESGzriLlM0UVWLFpSRomgVzhnZogNUxcuZHqeTl6ltQ2Pu7xV9k6ZsudzPBzYBaeQ3ZqTvyoW
LLGfD1+vWqqpSgdmCHwPNP5asfgHUahcpK+eEyGFK/6ctSwSXZ+ZtBlSF4U/kO8+kf8YQjTkB5PS
bwnomF4eHZhGKmmTMoXkPkl7R4+ST1LjjehT1idMl0rWOl5nifgsZxyWPAovEjlAN+fRL+7Zboj6
sAiYgVFglRJQ/QE/eegg40RCTq0KCXouT5WtH1P79HIkrV7jvJfJ8dZY2Y+f8lVz3hr4ySU7MKie
i5pOvQaorlRS+BB9vraSQOe+Pp6BganlyXmfePn352idJ9J5JEQUPyoefLJiq4L/OBghFLXVJqDN
VA/6J90iFX4sgT6GPokEnlJqZ5eYZ4eg70SLFhuJoMMEUTRPvUPEfdx25zuKMxKQ4QJfp3vkw6+k
4YHp2pqlnt12yS7Q7Mrfuwp7zhE7VU8RdtxIIqS5NLjaCOjCuS44OJmy5BCqxrIQJnIOvUvI8mHO
cXDnSNqgBPsj6m+f4VW/NjDiClombCSsP5lPV5/EPpw4a+JQlTGs5r4b8BYXHd5n9jpScmTziHEK
EJ9AWIpRI32Sc6GrRe0LNjNa9T+xEvPx4Encf7L4dDJmDgfOz5szm8IMLjAPcpo0Rtgx5Pkjum2M
dx2HA00SajgVZXiGyq7Zkj5/P8mtLToq2oT5TxsQMwrN4oQ5KdPdtuyWULrXiyhMRiBgycvgL48A
Hw7jkWn3fCkBb/8H56AEe9kRXZOhT+Xyx2XjsGv2G03R8OV0kRrVR3nytwksLNE7vMgbhvP20WpD
3SathVK3Faq3Wy5AfcU/RUZGm6mjkiILq/7seXxFFgDvnwbkt8Ww/nzEc/luoVuMRRdUiajQlkp0
81vCosTkSkyBj2dlhl9CucNFsCsnth18jhT2AYDb3464dKyxY9NZXNLKKvEs6WdSUEh391nkaVoy
g8TyL6F6zMK03haMz56q9ytxW7dD50udnMrsjcrrE9ZlQLgUevHwa5O3UDICvbw1niVdJkURuKSY
drgOtq+Ab3vP9sdtghyRSgokG0POhikY1TmRsceiHqOR6Nn1R8F3cpWMnrgB2W14zZUcROyRMlmE
8tIhCzwV1UwBlEFKyTHr2b+UcMDTwE8pT9QEuL7HBSpGNodsA7YuzPcYZw+AnJK5NkK4V/nxYaUH
8mZCZ/DCbmYISRpCcmL11wFcjX7CZ8pqqUhVVS10GDJ/rwNYc5DLNT5zCjBbPY4kKDk/Ldufutis
Nu16vhOTj19gCax+bx33pMQxUdrynnR421rPnpWobG+01X6y81zYATA4YMN4JRuti6rozpjBqgF9
ge/hP8TRR8GUIs1f+Ei3k7yvYP0GVtxARH4zN2/clFCPlIuEiTG0hwqOo+TgEG1y0t7wviySLvD0
Kv2JnCkErUUGPZM4iU0/U3DVGXKXTEFT1pN/Dx5IpmhlYcLbl785JGBvww4Iw3WJIHROnCXTJv0o
vkNZpwfYmG8wFirsZOanZkjijd9hZJZ3q/k1/EzVM18B6QmETAfkTckx0dxPlMrodubsiXCWfy4H
h966zI3KWo67to47TJjeaJ/O5o4TUwgtxUUZpye1zIfJT0J+et9BEz7BALYq+PhI7SjzTx4TUPpc
VsGx8EJQ0usg+FtopAhC3XcJYf57E+EmafXenkXjBcaLPODuKXuOjniqa7OQmRzmmHI6H6k4cFGl
5HxBKsmH0jddw+arFh5C4111EHn2pYIWannjT/ZZJrRvFDFTKTk8LWQl2ltSs6tTRNEbpPpuEVa5
0mhf51niHFtYhmu6J4YIyidgLNQtisNs5iCVn+KsEHZAtoW5c3S+Iq6ZLUfOECZroerofEo7TZFM
O5UxOydKft4g08iNK8W4JH7aaMUBrQwwTWLpocm+I1oGw2Q2qKdRLYYiIG7j9s7+Q01f30ifYWr9
cQdNIFXip96fc+RD8CUe1ZMErpm6fT5moc4uMLsg/IbRLPoZxXz1AoL+1NYv5S3fZiAlLRbFSTUK
Yn+qdIMIXtBp9R/Rn1Vjw71DR5KTvO9qV3Y0dJyUh+w2q68upJXleJwzf0YThaoCTAuk8bdKVw0L
cIby6kmEE86XRscjyPYXxRyGj8/RIv7oTccekDb3/4mJbOP4mNLSRBD95T/8LfDXVors1JAAOvPH
AfCgu0e3cZGXF3jIFre3/C94dSRd2QPaKbiKRFpZsG+iUslUB6ReOlYKA41ynpckWGn6gPnm8ivY
uAeuqUr230GjL/NxajM6nNzSrIQcl+D3grrPmzUNoKzIY6EmrJM93DWNqteiRFu+c7uuvOaRZUNn
G8mh3N1/BdRDc4Ft7wMw+wCK5vS9miE0D3nxVpitYLJUnN+GDZvAgWYO08Xg1xMpkvQVuRWJr6TK
Jp5TMWyzfh28Tdu4egxsg8x3TBYxgUKHShe6zNRAarXATc+CCxxgG40kITQGrkwhsFAu3NOC6snQ
L7rw3QExf3XkiTAjpDEhE3NdZzUNgAuYuYImt+TXrdaIkjWCamJy59+jFUxwkVSLNQEG+OjZ7wVB
OceuC8PBEwu1PpK6gM8HVxhhjgGGnqc2N4MqA0hSotqdXytHovWvIjJ87+RPW1xju2vpv/r01R9D
sjSISzdz6BjYzLGeC+FC8BiCre+Z8yYeKLh4r40s5qlI96bMqfO+HVlZnGw4sLQRTfjrG4UjKXir
bcGkjU5CLlGTWkK505nv4pig79Lumi/H80//Sz07Ms18gxp5FFe7WDc+Rdv/uo2LUGyWei/e5fI0
Ys6SUOMWhmaesx5F6YyE54jISgfZajHCW2OIvBl92Alxeh3B3Gae4zz6nTnSqW8RYSRneq8YjcK2
R/7jCd0FJrb1gp/K2+ucpfNAqvBJg1C+7LcKTEk49qiHiGhQ27eMPW1H1lmOx48YCKCDem8Wdslu
8lFChgUckrI23FSXRidC41nt99Du8I8eZOPD6ydkcax7zIGGd5+5Crf/7tKKGfnUXC91459wF3lf
20PDSRhLSxJ9ai20xZIKirBhVC7ZHVxGNKlBPwK1b6wBjp5FYT3UvBe6pgbzIJn1aXfVCHEGc+5L
+9xym+GSp9jsmiHeMzMRtHv0ujL7mZSFiNnouKax5EZrgIU3CqYnG0sec/9rnImHudnwRHQRWloh
SJWjZ58Ag0qBiDUAHuSKL96eduLyTXiHFnsiAoqLPExm2Bhd7ArFMLE8Fw3tXrMw0ovNtlcwKH55
sgAQ4vMbctN6KW7yWOtnq96g7zQ+Q0hkCo70v1I2Z7wboi/rVY3uPNeqNvwQHcRRlana1fcTUJ2u
KJzBvyKeHObgy2Vaed0eecmTomUfO1T35X6PJa9hR41Ut70l96sBtkeM5pq4dr2Ga/n/azwMCJUw
v7hYc6P0iC3qZv2wL9z5UaIeb2PjvWEwSmWlNleHP0rglYW8iwPae3Hlm5+kJdNW2T2LN8k0KoPK
1NRkJXw/ZTAqACF+hSdakBgW2gSjt3yoihzKvIF3VVXG5/ZIdTYzK3+A7tOB/o7nEQfQ4CHVSNQ7
5Jc9+eed6Ld9OpsfPy9NJGnHzTMAIvlqPLywIqpGQLYMFQP6/OwqPG0bUZZX5zRUAkKKPzR0sKNX
DmuoNksXQAuKVpiNi2/6d/JtCpb5Ki/8aehToS5tpZ4bnlHo1FwtLdMGgXMySnkY+VFhVn9vSDSi
kkj8dKZ1JDSmN57i7P2MN69CsUFEMGh5befCncIVT83dQ+g0ip8lw4qdPSgCUF1X+9qonibSwf7k
yaaDfKiXkAudFerB6UXyS5dBPKjzeuBazYPfBpEz8cBd4HE14DVfrnctIEiPGNosw1NgYMQb4saX
Om9FfZlbHJQkLeBd9fFMGuV5GHg/69zwAY39i3BbY3GvTwiEH36BNDH9rQUv1d8Q6Cgot1EwZxZN
LJjVR4SQbAMssmwEQyQBVRB/SByIV0vB/FyZeBh9Q8kqLwKEdlnijzYO94Al6n3HW2vUyR8QgAn+
PBH3+onwuM19K0ryrQeXsqs1/0sXPT5TKJ/FPt3QMjl9fvHf9gjFe1rdwMr/EZXrnm4twIaRa3Rk
69WU4Fdh8J8sdGuSCmjZQV6BeAsZMUhPrJVicwSnF7gM2+vRUkS3sgIKzeL+53FFe6oEElEqRrGc
Xr4EBkCdF/7qF0YxXXgndUH9sreao+Kab0gCw79FFmwUB9uDmdoBlG3S/4cLzS+08OJclwl6ajjc
/lXX7aocQ1x7i+uj6GRQJAOwC95qz4lr4TlNsdBxbFBuBLl+7OYNrLPLi6wfJBBuvHIcFtxB3Ufz
Fj9Ox4ff89a3K4T31ZbNEwlQr1e0JDR5EsXBXUTxym7Md23iTvhZCIoQaGoOqCLz9jbRjLaD9nG7
LEt6amCMnrSmZS9N52QbPF/rXNAKPDd61RKGSS+ZB+U5/DwU1UrgBRT4vtfs4d9PHX1I0kILzny8
7Rs9fWGzPPs47DDozjSFQsVk6EkIuIkKh+DJyZSOcGalSsPAAcgSDydUmWYXo1L/3ijEzOTFTXjy
hq13jLUZ5u30GuT8U6kAhnu+T6TfUU4sgUJ9zNdEUnvXItxvzLXzyF34H9TTiMUyU1IaFHl6Q+8y
qOtUJ1WEqQHHgBeKFHIeYLeB2A7p4Geza5PRxrRteimFu5VDB4VoWoRtq5KoV9hNsUGq8GcHAma6
xqJ9sdFjeLxNe/brucU81Gm1+1dpDE9nLBdfDcWPBNPteNdDeFX6UDaEO+J9xcH899GN79EB3XhO
8nuIAKhWnVGY4TSDYX9tvPhTiJU+OXUIlpmJgSHYgjV+Cv3dMghbKswHWmcar9iKGOear4dmtCk9
Y/qBGTqlh7Bvoq4VIXrooIRM4/r34vPBt/byUExjH5PyttIyq0hty5a/e7P2XYOzd3nfV8C2Pg/J
9BWd/jcoL7ad7EunS63GZ/+86nKC1+SiHYtvnvxyVmljQpJOm5TGUNkrztmmwxbUBDHKQCdBsYrO
wCXJyLFzyMgnHER0HOuPRejyZ17WbfG0kA2qtir9RWJvWtjtBDMx2Giw12zQcpU1PJY915jqvfSj
5LR/ZjmZqFcW5tMXV8xs6/j/6/FH266Jmi9XzWRCoWjkLqyFvL6TMtuQDCMjb6+9mJyPwUUMDicQ
UuKDSi8+9HKd/U5+YBQTGah9M7gj/795KEwot0hYCK6DYBWSxi9pdICiiPlXkC5jn1BLy1jvPQQu
tvJWJtKalYSa5MsvcDLveF2LDvXe7eFrX7ufwlCQ1EJtjlrMMBIUB8LQ/cIeRqf05GtNfxTwTA2K
7f88LYEq+YcQj9YzkAy+t9/SuDJnetZQ944p1kRbqtdmo4zrXNOYR0F5kMuXNBeC02VKoRRFr6ge
b4HTiU3ODfQ9vZdiPdMWkFlM6ElZA+QgYWdnGWd7MWjOv/C8fjI2s5fULJV9XTGJ8C4IeB1A6L6I
cO8nsGADpHqyQRmuG9nvYoY9Vtl2WGIweNPsSrCO3bqNSspx/BfJCj4Tt1mXTLlb8ezdiRwMb+9S
VxeNuf16QAecUznpW6WgRCoYxzx7xGN1GUI9DTLiLb+b/FQOTg7PvKN/FvODC0W6iMbFV9y6WIvV
oYWbKAzY0PfFKXB7mhs1gmuYxxa5biz04IVjQWRqBgqwBDiEZlh3/MbNp1MOxZ6F1gfBTwy6zxsu
/QARk8FQw8b6oWsPvZ4DEbs1BmRh2AEgpltkDT9RdUjjCYj5SLLjHZD+1kt1LEPR0w9j49XGJAYo
82Y0oVYo+WuXSMrl3M8TuJHBH2sQLY402S660+5BYeHyclREiB/XqozxUvzi/IqsuCCiU3kMMPcO
0F6nqboOQ0Q4KURRoUoizEE3mxNlImve2xVdquO2V8sic2yl/8ANg5AjIq+YBxxIAzAvaCFRxpIT
0eQ09h+2oqKFA3IJ12S/ko2zQbnU43M01QH8qS+ieBtTSwVtajDa6bliBx2dNJ75h7jGEShmBPEN
kgHyvpt4DFKObVIu5G5cMLNuEOa7e2yPruQPeT7PaOsTuT0p3dYdjRooQzaFkwKOFu4m1obX0OJv
3SJXb5GNvkPf9tErXJUUOWS3KIymO7Fnx4oOwu7iCxBX8x3+YQyF5ntLEUEwdOmO0+pDnkQgDBTm
ILHBcereSjRlLGXnu/T3w4fz2ceXUkqffLz5JjMgl3qeuZMlklPBDvIEiMSpq5W3zio8IbesaOwy
gx8EriAJlTimANhRjlPYMzR9rAr4Kx7pdfPXqfZSRz04KbUTmGiyj9qKvFRuEe/NkBQjOx/zvF3c
g2jeq64cllzfgS1VfeZKNPyFZ3yToi40g705qVGZ0sS1vg1+TCQ+CyFFY7zY4j3CEq+tiEHlkC+Y
YN6fNEeh+6offHwnKiyHo4GJr11tN8PqlJoB/tjijmF7JsLvNLu6AmBf4HeWRunRYy33mX+0frGc
NW9IfHhojtCaGVdCqzUw8Ln/jD1XJxrUddCE5Y+VrhLE86U7h1xhZ/1yE3bAKvGWW/Su7FRAo2Z7
cup4ePKelzWerWbxibGBYSEX2S4U3xtLvgoamjswlT0llt6KPdDq22hjXUJwSXKGqYAcsP3Eg2kY
RhN3t5HR8rWj2rLoNZVoHMWx/wx4rtIsKN2IyZ5Iw8kLSLTMoJegmYLC9NQwvMZebW8wwFr8dew/
+D6HlDuyKrK13dWcXbUPGYL+iZsfWR8N+f093GwZJgGyhMfLeKSUmhPr/SmlYJihyFzlCpDtoV+Q
aFoCqUr374XzQ2HC/qH7AXmjj1we3vbJcGOw7ZVHWJqlWRTS/G7wQ+fX1eBIv3id32v8L9la3XMh
oYc9R1tydLTMXpG7KbA6Hn1ypmfy1CMe6OKi+RO0y1/GWVEe4s/5xUzTijMupwZqorlKgzRoPCxE
6xoK1Z1+oNWRrwPazEm94bEk+NdaGcjpL4J5flWPv7p1O1mdSSxpwIbkCYYibg0eys4wgrQ4md1b
8G8ODdPxDFXsIs7bPDj2EQJ7/1mH3rvyKCiHNGyKak/jVYrtEj3TkIKkckfXDfpXw6+AsTcoh9/w
K/RB5JnuQ1cHnEsmPagretoxQ6aU5BisyZK9tcS0CoHHYsBKqC5NM+2LoMXI42sEnvQLfBqvHFcs
vbUDQaIoe7/6O5rBFRs3YGZacwnTohyIoCr9jndrLcRBc/6LMuLevXoW7wsou+fzMBXJlM11LUQE
84UgBRg8K663cAYLFixGGDvv0+mf5AieLXdFML8/p3sfvbp0QFZYSWGa2aCqilOCQLSRPDkb3B6q
/DYQb3+JF3Vn9db5uO1jI6H+2DrfmiG+MbqJVcwWpa2LLgGqJ445rmaF8XtwTjtKspcf0xFunEZH
aMZWAh9f5TzY4UltiDw3uNOFsxLfwYUs4jrkfm6ioWGgAgBVS5C7eVTprtUiHF66gKZP1r3nQbCm
LnyVNgxCx49BVE5QuXip46tHwsXnZj5eKWVYmRr/wLVHky1eYgyUYpSPzZ+Fj4O3ghBpzta3F9bd
2rk9sg41yKX524uD6P/vuoGfD7AU+sruwcr2VaZtQgRq5aafFg4YgMFG8Yae6MW50XtvdYZVZKHk
L+FLBu5FkKbIohZFGWPAJ9m263qCfD5LJijEZxryDV0t+49YKaGsquv3t/9E7dFIes4v9r//QX3e
fGzQ0tpavTEbGTZSuFjh3vEzhT+u0Z77K3ToS2Cc0WgaFtvYZl6CJDW2hnp1LL575xDCgpdgQfSl
YM4aSPHeLOSzAQLplInq7n3kv2MGJz8euAbdL4CZ3k+cufyZtsojhdEbYqbZH0lfoJP53MIaZbqc
4CTOmypF8vr1uZR7AsX9sDxzUobq2JA1CCMFEuBMdZKc4EvX2e3p2vtDvVzNAxd0zPDP4fw50DIf
n9Jfwa/LCzp8lwwHStpnV6rL93+Cf9lZS9nXh9uoQlY45UIGFp7XiGs4vJKff6QZRyieV4D6B533
Te5NyUEY4Py08m/D2/3NRkMfJGKiScpnM6PqPcpQ9WApexkIOCqeaJMHNE5CPTj6U4LXxpvOpl6K
1p3O8YLWCiRnSJpHcgdeBHkSbpcGsdRRVqb7tmy5WX/ff7a69wtQyB/WjAUcg5/+Z4DsY6gwK+KL
HZJXHnlOES9e51YlpT9TQGIx0DgYNwmnU6XJC4vXpdG1H7hAHS/94V8h0TorWH+Gbb+Ywi9buxNL
QdXhgQOIgNQRFos3cAjBlCGdaXJ0Fqgi8Rpll67VxN4FTtl/chtyrXj1i1k2StNPSTjkovxgQsI6
aZVKkOLOUXWYkt4lyJKwys9Cu0ifUr2YA/5ajgbMch1uj0osQcnqjFe7O/ZsKv0eusT7qq8OqFt7
QLMSdtoF/Apc8Ii74UGGUMK94hiSPN5LDYK+2NY4hIgwuky9NgWjQIc0A86boKGSqyB2qUyxEzsR
F/bcLEGWW2QJ2HLl/ln1zD5Q0WcT8M1EvnrtkDbobZO/JfGSFXQVpzVqVJvc/S+P5G906YS3DtOq
/nG+EBJZzSJEzZRdCaef0cNRDyQ1EdpZmtAaAfUqyEg4WDIpPPMJQXyEjC9vfxJZNGqFyW0VTLRH
pXSLs6FrU0Mk9x8zsxrFFJ1HBitLsqp+2FX/WTOh8BjyGXn1uABx7nklIP2aia4q/J8/CNuMMdpM
65fu3c/LXNA2+e0Aw+Kup5avS6Zj9NjWvPA6/34wz4pLlTpluDb7WLEYcv/NJOY/JOYT++1+vA5A
Dh9Vh1OY38UW3lzvxlJemAkYKPo4MUGhEEWFjREwtqRKrBuH3cl3gGokm7JPTUskHs43EqSSHJtE
umo3qioecdj7BCbQpoMQ5ZntabWOSO2dbxUgd92PCmM8l47v1cmUjHkpxNnWgAQKGAtVZiLNr+zl
nRC+vSJRFLYRMHTDOfDH6idJ3nE8SH+QODXgTtUaTtr4PsMRTRDmvXn/hmzKVLnrVUFPiuHj/eb6
Yr5b7JnqVuVZy6RE//Ar8SwL7xDK8FdI5SLCplten6EZShF8tWZLimPEcgLIZXnpizMo4uNe4Ir1
rscm+At2FsayJXF52WWSTa95lcOgzR4gb6N46gRTBIWNU72k2AE+1m0nnl/HyA/qgi2gir/xChWp
2XrHVnhSIiOu8r/iNn/Z/20YlkCewEFZCYHuPxDdyc6+5+KhUBtldSJCcZxvIaruiqQzNichZYkT
yMWVkgcxFstqmmkaP+o4t8GDPDD+EHJ9UsFbhKxT0Fi4Q3ad8iiyV4JdIzbTtDt+OTdaodO4mMJj
7xsZLdanKUlVeNhzmxC4uAKQjK4PypIGiNi4V53pRkOutX6AZNtwLjYmntFia59vDgqdj+kask/j
CWsJLMlGW5mpONoO2PNGHXg8+68e0TetF90eEmu8T3scpwXYqYkD10p1pLhj2bm1NlBMQ5zZsNZ5
/AmEifAyOYXQsYndz2e1i92xet0cPzhzPGJafcNNyLp2e20W//zF2NTXohNKsNK9nqJueOpcRXtt
47VjRC4tq7mlTbwgjQ2sca7oBKe7Inu/R3XSr/5f2Kg7r7DFP1/dKOdO/LjaAQXJiKDM2J8YJcIb
B6eo4/f+ZIK1NzB+7sVlAkDTls53x6UJvzQm2/qYY6Iu5wrYnc1aSVB+4gP/SlEu0sPspq9dEHpa
Cb36KLyj3OmFZiESu65E7QIZOLGZZFBX1NBorTPViRDZ9Oo5GJrg8o1nyZ6vo3NROrOEC8IqK1+7
KlPnO5n9BLgU/WgrvrQF+Ll1UayCoyKs4Ozc8nVq1VX+Hsh6OzqIs9Gg3mwHAf7bheHYkH5EC17g
8i2BCj6C3dSpk1+hApzSrMvJfTi3GFksq//p60B+1a9dEwS2pP3F72TgBP1TP9JXUST4udCIJDOX
IBIQuyQbduJtVj5vPMhKX2QVvZDcOYyZMcQem0IB0ILSOqG4WjX7DqdfPeVI4zah+hV+KTHEDvbV
3G5hUbE05HvxidAEj4Kqzip1MZiKNfWFBTCU6Oc7BXEkRRJQtw90gYIycu43RMPVHMhENhm/xqfG
BSbFdnM/49F+ETMXzJMwHTpzF6oHkhQSUhd6ZdFw7ZebfeLm0Fy8yMkvwd/zR1N3NSVJ7Vth/MiF
6klmdNgv/7tvxbbZI4vO3Uvq333XdP35Za6Vzjr+g/K+7cMQ/eC8+/yzTkQVI6yMygyy3yuz40j9
Q0vnEYhWFL/8kAUfFxz3mtF45X4eC4tJaz721lQ9gsk26297qZmKZt0Mu13EHdmHwU/PQlH/2iLH
NOTcbz4rk6kyEJQqIqSHr28Sl/aNtnuJnKwWOY6TcCk2cIGJvXqpCrtpgmYLDWZrSqN+eTNpGs1S
rXCswAxTeLWDUlmeyyXiJK878vMze/xE/SffsS/F71JUCv5RFjYTWNgLDjEEzJKqBKJNH8OWEXsA
3UcS20RLQEqsBZMC10o9wF48iixvZD5hYtsftTcbKyNXGtJyHBaJY/BtWCT9VXoWilWotjKbkCSn
DCtkDxKELEtkPJ5+Xa1wMUvo6hv7tb8hV5Hpjk0JliZKhsw96Q0YBVqYNQut+KKYq+u65HMdBz1s
LD03fJSupOlY+J4iIFk2YpEQ3//j5aygjqZHfPm83ycAhrYM6zxLMnHvOiUHCM3/Cw4L3y8yxvin
biDOntbmsC/1OGbHen0mWUKKWf4OvYfRtcJpSdr+aTVk9i3w040emWpecx55zcD6EiCMFEFP64L0
TdBPzQHOCU/DN8izfE0XEoG6wr3gBri18WkLE5E50tkaADdKH4PaduuGbRejQP05BHYTdVmRJ2Vd
Uz8V2q+MhPlfmL4kyvqCgl7UH+8eKvS+8HDTqU5un5BVbjo8r+hBRr+kdAD+1fwsE7Kr2VC+8JaK
71cVkJ38TrRWH94upPWspPNY0Y0lBm/yn3a7kSNcUzk5ji4X/fvRTehhFTW1FBaFkjBwIW5nP8fE
aKnUgYTbIJwOtXCc822La6rCbcotjL1CSw+GQuJ036nh5mezW23X/rPYCaG3a6GREqClQzZ+cQlm
qAB2tWop9qGTCSArNeA30iB+Jv7BR7snWMtn52Kz61McQpx+nV0LMLDmHqu9GylN2nfMpULlDyBU
Pgt19Q/KN83AYdEOiptxl4alPsMW4TFDO/+9UzHyR6+8ZbG9WQs6x5AcHDAL+rnduAzu7e0PiLZ9
J/kHXrfFF8qYKCWgTZ28l7gB2WNnllaSogu4OORquOY/bNb+a7lJzSfRnOq57wGI9kvzgClm2beF
cNSqw4neuSKX1yCPVsSWVBvzWhcMuiQd52ULxbt25vtQU4GRlLCiXjZwOJd9I5c+rTIMWkQkQOcB
6RW5g1RkNfjONdcSlwQD5+26BNVx5smWafz1Y51jT8d7bIj/Z+C6uva7b+Lbbc0litwbnom6cNfI
OxSR6STMTykHRXhuVF1y6O5yJvgZ6jEHULL9Qcmu7vdy1ZFnRQE8oR1Dn+m7MJxdJplMYvddtGsG
9xQKbMAFWcZIak6BJnDxVqsVQiYLPk7oLt3ojJZCBUMVvRAFm3xO4AaXRDogbjWN4cYvE+agAybn
yIJdkl4AftSST3USG5NVyXksXq1BW1jmB8ix0uZ3MF3bMwhAZ4xVZ9Cg0lcG+up8gEaqI9sidj7G
kIwpJnRqO4VtcbjAYe5eYCfEdN8nfZVE6O4YF1m6TMXyHrKpqpRqbhHjtPiXHFNrqrVvV2GxmOAw
gkPsF3gU4hVTe9hZPYsa2jNOTZ4/TwPT70qSnLs0l3zFvZ9IxpGHP0lTfZjzfpQCnv981Bn6fPs+
aDPX9eeq0KluOxzn+giTnLGKJvmzYLzcXIIxW7fE3qyInLgt46/Ez9Q6OKRfyCklzkOZLhRX/x70
UcmAc5Rnxrvmv7iUHxH5QoV2rUzxR1via9c74ruwm3RgK8JjdNGkGhnBTN3I4qsBKvGxkobYyHna
idaxVeteJ15V+AmhEobjxleNPOOFRdyub5Xy+1KbzsDVs7hLZ3/f9dkTGBk8Iw0983sWA+ywC7fg
g0u5aK0gAP8XAjnbfguzwIbbKOEQW73/wf4U0xL/3aMlPQ5uUaL+0rNrT5RtustCzLmx8BDgXu7i
dHI+MWSrKbvl3GghgLLe1D80bwILcoNT6zYB9SRK+qBlzM75f++BFn2yxPgjFJJ37uF1pX0AdqBx
w05Xl93cZdxmGJaUvSjWoE2gqm7gmcv2Nr7opzWsEcaQt7No3j7y4SrpiipVzupkwpxkxrU5CaVX
lR2e/MtaEX2dQ4LaJT5a/TLM0uCnAfrDohrJSlLL75nijirHsRz4lOoACHVcVdXqOadtbDByrazC
1qAl3uh1LW5uKapykY9u9ra5FKLrKY7nSJUfFEFnPpP2W0ydoxetT0YElni5F0Ea86eOmmLCAiSL
LENkmTM8KOxgA05H/AVpRu4QXnt9sGkyQv+I/Rz2aV27XDF50ZPKzPM4f8uvamtnfIo52JML6LDQ
Kt+JuPx/J6M2PmE2UuOPILSojXxS8oo1pLfdkizRsb8AIA08O0yB32a7vc5FNAY03P2fY1kYU3hY
3SqWdBs3VJkRKvEpzI9sP+am5vmFp6tOie0ul2jn5sN9btxyLfkLo7YmLzERWHgtA5E6CveCkZsm
L50wi8sjki5jfNIO2KZi0PjZwPSF9w3vGuJ09uyYd/WMG9310dWRhaWKR6HDo3BDniwh/DUL0+C+
2EQFvhJrUoJMewCouum3voZEMoxrzWwwftkyxu5pTV0/QbukCcpN5JyvXCLGzeyf3oQCaKfqg5GS
cnxWckBTXuIJlWmYeXv6hPTnsqTl6TpMgc1SExwO70cZM7z76zUsMBillolNfJWj7ByVJGbn2o7/
tksLwFdTKcpcC5X3m50tSvHJvD0fF5WfwwjEVpISPlxzotCMT/XyCyf+yy8Qt0bBU3fyXsqA2eLt
yOev3IgmiGy539apSAW3tF/PXSvsVM49f9xssTzttv9aF9ycji6wT7LpTWnZEZmk/4iGGzg000+0
bjlIXoSX0oh2GI+fjLdXuntUEtHU7tTVW9aSwkKjoHMLwaUoObDJrXzWSWZhkn1ChCBx1XwWUY7e
wSIuZm/IB5NXBFVRRn9D1578DVDizBcUIPzZCm/gasmsxKw+RkFYvOeVSLDirAY/M5iodcdaPO7H
t4q1c4Qa4Pa5E3bl8JY+xJKN5Zj1P/Xef8A0S5sDaIb6JJasUHwvGii6JPjvTnhYc3fGvezvjJnH
2ukLUepJmJUBE6JJizuc20Rthl9cjB77DtwNbApBO6TlDrUcqtDpzT79cAUE+5UfovwakPj46j3J
RV5kQn6S9fds/FLlbJ/PvsHm5hIfc/9cXybYnu4YqpERneRF16itYIwt+pni4Iavyog7CoSTUGoF
MDEC+N511X0S49WhlIq8lhAYSpPbGIlWt8i8BzwdveEpRti4J9A8OblULLEikwshUE/4GSukaKQU
Hrhmgx0w6Dh9h7tn0/MBKVfDYuwnHHykeT72fHyucMHjrl8tONo3sObt/9hhShnIWGtRNhy1lyWE
aClPdzgNMMPG+vQDn9e1rFewxmD4/6NXxF9IYCoAs29HZ1yuDsxzyEeONwwPKBOLT1ypxlBMSFLN
/laCL56xXE+a5eWVVgvG8iOPBVrKJOKZT8yYGWHJ5c6eovB52Ncj1jxZUe2SirsV9lbYtSEVVXQ0
g/+1i+OsuKOrxWLzJvkuf3kZhJdyLuN8W0K6EEdW8UM2aJrWCSSuBvdYh+YrJBx1PcPbCtFtxxJr
eqkLVhxZgnUfQQ9Qo0KyXMLWlJ8N0dfLsMn63jy2xp7uQPNYTvBj3ToNC3TrlJO3bbgwGNMaffQf
kY0Re6rOE9dkyGf9Vc7LwTxYYsCp5FkjPuFs5aiS9dAybV+WekSVd7Q9IBgBnG8ILMiHymRXskcC
j7sDJwgPfhzTHzNo6/atNVSE8Z9gESMD232WzVzMUDLKaZw+a2tGllmNTTBnLNMF29xiaB2T4bsJ
iKCLH/NFoHkW7HFKcYridz8AyHKx87+tFuXLHHblZ85JAnxOYRgAVy+Zp5mMBn6cDGasGEE7riAD
OnTLv2fDSMXcuL1uvROrOQ+jNmfamPjdCfRtf6ZC3uAtpVNctOfCG+lyReiJ3/e+OVNe8i60fz9G
fOqps1SbhtdtQfL+jbDd8lR6sbjy2dnecI6zeO4vvLQXMuHQkRe/Xi0NMs1ZQJwgIyDMjdd+7zlj
I60m6ReD2qU6/dSYFECb7buGq26ULp1hghgRMP/qOuXVRtrLd1OIZyKM4GamqI4KdBIpJJZHmQHp
8z4xwh9eJzWutM+qlw2w27oljfvrZwz+/wSAhVmQl/Tv35YZqqkIaCgSyt6jSvwNfc/LhUsdLHyf
CjBIkqMiQE3Ff0l/aQuBYIJwpuV4AlgXpxd/5YcHNcxR3nbf1tVdsVPOKDRAQvaZ/PTb/1Qv/zzu
k9XVKsWSgzbfpk6X3pVBl/I7Cx215Xb1qVQFrDmX6lyAbeTRhRaBNstArFw4wftfiZSgNq9EAv+P
5GEyseSUSmvjMLxf1i/hkk8ySAC1nG6+/qBQBLbeTDlm9yAUUJhg/QJloS0JRgU+az14bnOdPCQh
4EL5c7+XPhEaM5jK0sKvbZAzeQYo9LAhAYLqauIOhIZRCiB8LjXeA4rdpSyhVbt8Y6ZHLKJn2ZuL
5hyrFecc5cT5INVWPJsImaptqiz/jxnlmNvoeiPvZdCpfC188VjderpN84mSUB8sFGFwPeTG33Mi
Jiqe40dk1WlSJr9hBdIN9z88N+jfNmWPs94jmE4KkpX3luZefvjJMGFmGnUbabCaXurzYsMIGSzH
1t8vPsYVKidz00H1Wj3bvbLYLMp3cwGbBvqqe2HwCX11eDk8YPR7x6S1zUi8z0sLDcVp9vJ4Dei/
JT6Y/glEVZrQDG10wJ8p+kwGGVE5git46IpVOHskyM3INdkG5EiUGXx9Hv0WaVZrbqBge6n+ZXKE
cnmDqOKJHrB8XysUtKwRgRRTPb8K+tZMGDebMYW1xQ3ChI20P3y/6ltw4aCBCa50oBTLcMLuQcgQ
G098C3odkhCx7zJDlf5ArtdDyOAYvikTPI86rj523fDaLJK8peZXiCsl7eDVAvnQSYrt32PRh08v
3T6ZYevalqvrWhku98aYDLsmCdsJD0gilSkxhB99QkLIycUp4IZVR5SnYICs0g9v9yRbC24d+iIp
lYHiQp4oeBcnKwF9t7sNYUfDXwK+B/MQAK5X8ObMJbKeagl/Mq1p0W3Si3nzwu4U3REiwBCa/ssS
pWjPhbVLCG9YN39ZU2TDLoKuijeoR7vp2JwSRHuPGy+wJFo6CHWc4vmzS0YSz87ziR33wtp4cC5w
rSZvcRcRU5K03B3uqEJgLIddEY1hytBkXB3oPyQh1G0TOhJALoGXVJ55+VXK8TvA56t7uolWW+qI
at9ErEMdeWmFzx4UMLymmCLlXmwWDoRBBZbpHNtP4oa+1+zFotODmFOI9Dy7TdI+t8rAIUT4rWkA
ma8GKRUR2PKYtskLVMgqDWkzywZHz2xqAa4Mlk2Yg2hHHcSEaiNKFNcA/tCQiE8eGvFhzIqb5oTF
BFfpRBuUl2ov8wwkg9QrMJuPdCPupCDwOzHr35Q9w5nYNCngFK07HShtrubp40KLRSMXn3/gIk8F
wkoyVDCcHp3b9+uQQMJnILsuZlnHDAk4K0zNfCH4815R5pYRzHGl/685BnNagLIgyk2seeVeoUix
TIEMJfD1LTwcP1InpsIMIsr3vjCAD2lBC/vRoCuXWDPKO5G93s4pk/ccBlbt33XnP+wjr17lyElR
iaYHILq7JIS3sexQd4V7ippw3xNUEM/yEvxKgbFOytyHtc2KeVqtY/73FDNHI+m4d5EVuHK5cZNM
Z69IF0gFBxmUQPR4o/6JG86RQ+Xwj7GTqt7x9K1UViVemLgjWD8RDXN2s2uxzdCBYHTBci7uC32K
o8f0IvkISthlojw9kCxSIDhuZ9XBX4uh3IcQZtVGTzwdTY6q2rHHtRgp29zLHa1dPsm74QCsGIJd
KbtEqQf/D4CwaBBhtEV/iIvTWMJhFxJf93DgKzc/+TpRd3u13uBjH3xRkU91MBd9MtPEKRAEZEdd
AF+pnTskmG8Wi+EsrmPqqRXXBKKncE1T52V5OQR7DEGOnL431qOexam3Jtkw+K8FWk/9vwAAOxzg
Xt+m8TI4FoaBbpqwiFCEVANZNpvxhEqkwyOYQXX4g6JqR3spm/AWzjXpvMDEYFLla/BNUBu1CDC+
O/qN5OGAYW3zGUEi8/kPu7Z0uVSFsPXqtDxy8zzGX6i944tqZeoVuktvIfzw1HVCDfpuRqHlJize
oVJzGoCSkqwjc8MGCmnfe5Wpcvhbvy17z8LQhk8uF/5rq7Pzd6roVzRo8RYEvdc+OmbgvUc3tjhB
8rV6TYVWmsnxBOThA6ANc0Z1TqzdoV3vuBjhtEw5HFgG/xQnGbg8JLgqJ0SJOiwp+UCN92ecBzj6
1P3IhX7q/gaSt5fR6MiBmoT5QmmsU+5cAbf1S1lGJVcQUEBYGhH99wS4wZPwBg+p4EvmGMKc+o0j
HvKkFX1Ofoeh9EbKkc7Wb+m1UOaye92QATHN1+ZKlk4uSsHjLdfniPwiigT7G71BhFXTXVKqnyFa
5fT9oiiGg+WZfsRgbvqbpOVKaqSJJqZf4ifzj2FKS4e55Ot/NJ2b6DiD8XhkZWpk8r906+ERx23q
b8zlzm/fmsz/3R7vvVovy5rGURiLnyhP1RpcVtT5JqsRvQYTbhf1/kuKq9we2QqQYSWL6dNX9+FS
TLp8NfFC3dgZ01vw874eSe9rzuZ8L/ICSX+pJ63Bz1BVI4AQMDTC+6cHcTWgC6w9ldUhNJ6h6A/J
ST5yxDdfS6fyRWIVBPi8U3CEaHIK03VtitTk6PM9xVFliBX4dz7mD4uMSEBLAk2KGsn5VA2jTcKz
eo1M8+U/xiBA/EyMrbIsNorhh6H4p/JAcaYuTwhP4GOWMEQjpkGC24jKsOJCjkQXGbjVJkJ05SzH
QBjURiFF6CbZF6Yfc0E+937CRo51+ND/GdsHjPOIS/eH68ila/gEZe+d3UG0QRv1nzppBwMNzT4s
XfE/oHiNT8RwrMcxShrEi5aIPi5HaqMP/wjK1XhtMKdTuqbP6p1HTugkZ92c1N28obmHrcHUsOTN
QHgKyLoJbKdKIz6/HnsCSyjRMCN3h5O1DaB2q8Qwm8SKhaa1QXIxrlfZ3cg9WT8dkUS7ySZd8vlw
tqpbub5QIR4f9H/S84XxkCutrNSpdfcu+9p867dDWpfzMD6H67gFEVfts/4CTKA9RC983QFLmkSz
9YcxHYn4GN/j6WpBkUeAop+IYTX1JA9xgiv7rcHLR0fpBiu/d+DyoHH/dLmjWRDx4WWA4W/oN7GR
zQteubf+jyphPmHd1FkEsyyth2UvJz8J3bSRy8YWs6CpVyJyigfCFVXcx7lPA2foRch0kwdvPFYQ
raEF67mInmvAGwhRkg3DUglPxTsQi2bdzV52D6vq7kLVa0X1c3GL5QloDbZR2gGsx9RKaX1BCFJi
L7e4SuqtMCx6wxdM2U3frSTNMGVbfutzl5pfJ3BBbfQUzyISi4uaeoJLuYos6TiETWJg4qOojIlR
mkVLvDivhoRwArnyFcY4tbYj3S9Cu/023gzVMHwVqYNE0Ok6pomWaxuT6BejKR/2duMol/BBe6rw
E568NdbiRdQrlDe/Us6XNMxwOnh+4z2++RaOt+RwrTajWo+Z91N/2ejnMO6Rd08VFGYuJ7+quW5W
8wT8xWzeDTpI9nuMa9DMCqUI4v4A8T0i7PgGcY45dT8aSef0Z8dk0iuieqT5s/6Drp0j0hdoRXci
3Z375mVN3WkKe9qf9O2Iuf+QBZWwPJ/U5azEAoHR+Q6WN5Lrj/XX8Pt9rITT9VOWXkD+Rgs7zHUQ
PC7ATAkuqG11tufXjUNkOj4ySyGCKuSZ3dphQQhDx8IPsudYS3F+0MMzqH7L/Hs1W5ySRQuG5Vo0
Z9w5HNIWzYogCsbNsYqQ3fGGA18AIuCxQMdK8CCSSQAR/KzmOc2M0XwrlKBYqBsKFE8jqwV0frtN
CW5fi6oQO2MCWkkb1v8qiheDMiU3M+SGXWXdYLWIiixpnSC0JjPIGUt/iQrjJXzipTmikj4a0mTK
EvjBB6b+c+2F2iSedFENP7tjO2fuF/SQsUKWWzHPOTECFnHeSjE4HUwTq3jOiFpDLCUJKjHJXu3r
z1Kd806H3UsNFTT1DBy/54Z4oMoJreUygWhSKd7f37F+JJ1j5pnBPEOPQjDdu1fljs2LyW6y9hiS
sRdoFx3uRcX3zQlucIzTcrM5hCVJrhrYCM3aiWpXhMtJbD1L1avQp6kjCrdszoamojJGxohaGHfJ
oiJphx+J2Ad59clVGokbd4TtjUlZmzhkJvgH8vlZVgPSykZFj2Gjl6e01H0DDGoLEYgvTpw5koAq
0Rh0NqHLx/+ON42dQd07k4iPVBrpRTVACdkfkZtKdscYnjqrvhJXr1DV5FlOvd5GB2tyreekMbvG
oh5N2x9qMzHqDl/7Z0gR0kchvpd4SBrkKY4HayoI8WppajduaseqoZSUEvuLMMFCFobH15IsScK+
F9IN7XI+nIGJsN5LdziChPwuY7iH7HeRVkhfcvfl2C+daDPeG7g7jQFkq607qna90LtxFZAv7LT9
1/r69NIZWGrEZxuuy+V4/k47QUPKf7DyT6TNC/5Kk2Mq6gjI46VtylQvMgkM0yJ+i02q7b0vUyik
EvffW4yaJYE2bIbOHLSUslHtYtkipzUt48C3J3pbXyv2xeJhjMbB7uljYkFlCPArMtuPEaJgnCsv
7oVOGeEoRN0ySKG2bMWAIK4hivKq8WnJ6aKxVYjfh/4Cj/+d+nMnWqt0j4WMvLWpdZXF8LABqIYu
NoUpooeZor1Hs/z53kBP9SdcV6my31PdIZfWYe90OfGw6z/sMRR6Uo6Ky3tQeTfoPVBrrJGgr8uZ
99DePcI2HFug5H9bHj34JK+DZGAXf71VRX/tTtANDLk8exgaR54lMFk9S4pUlRSDJ3DoZYQ1dI2g
HHri05eL1brnolaQTqcnF37M9VcQJkIOph8JUnr/7Q/3HWZ+UV5IYdpZRAMeNstuALtUECCUd8D9
wGoKboQ8P1iUmTw7+XRCz28y+qgM83L/6OTIi3xDPwtSyzOF8lhEarE3H+k2Dchy+EFntMnGk2AK
UFFB2dvz/CvR6WqkWXe6DNyeSHYZK0A1wgm12B0NOLcNb23pUH9zpjquapRwAon1SfHx6vM75Iuq
EMZ7vsJVJbFmtnZApjWNC4KDXFOrBjaxR3X5ti9t5ss797IkyxW/dVCX6XkfPnTw+dWUuktO3fg2
asbrI0J5HUI0QahQbajXhpyL2FQUNMvjNJxUIGlEqAQhCQ3lWJzuhbcdlo22X5BByXZ1/L2waprc
/pEacBwMIm30N/YvxdGYxHG0iH4aB3n7BWDj37Tz6MAcP982Rh3WjXLPm5wkVcuanq7S1j7WstDU
pwAQAj969FzuXPh6/EdopTqPi30CaXDEMb7dM5PX/+hah1UmNPaPV2Azy/i+rzCNygfT/IPYfTN0
Y3QH1+JGKlLWGEWbAb3GrHfpjJ3ITu0IKiBGUuEuYLGzwTwPa7YkUXfR4dutZm8DfOdxGTnuP0Dn
QVwUuMqmIsrPT3nREQVEdlxKwvvIgcV6WHa4qGIooQnVZzGVdbx+aOQvwGXLVCqP02MrieymAC51
IDP3mwmLcbsOB6sB7qTJO5CAzbll3PV3v4P9B0EVNilJRnqLy3Rx+Ld2VApH8eVhWzYs0Wb3/BE5
6IXSeALnT8zhRJGbnZykIRO5Dur5pK1D4m6d9DqaP+sXI1jc5S6krMvIBR9qYiJuSUM5kmSIuqm+
Ispyyojjo3E2b0CFZkKG25zLdWdS9xx88R3deTHz5eBGxSNLMOA10Nnbf8AOXHalKD19qUa1COWs
/qki8OpKTPj2RSrSFE7rz40Ufh3APRaxiCAiqM7N0aYyKwABn55EFUkzY/eTRNh2o3thz8YXq9pB
CxYnY/8DEP7CgmRZCzmCylzMd7+pNy2InN2WwoBhjvXAEJIfYbOePMwHzS0HMzkzPdS6jLBNizRp
6G6UNjB9f5nCspg6wyrTzeX2Jue5K0Ai0K4/Z+sTc3Zcx+vAw4TxWNp954A7nrNiQlVmdgiNxVPy
EH1PPfiEICHCMPAnmqJgMOPH/wNwrzQXUlDwMBqEqUs3YFXcEbaUmzIdp3j4RikOdJgIqJKKahW+
rfThCjW8EBxQzAYq6zIgW+3bGtBkk1auvet/0i3Kd4euuVtovaeeecwqjveROoKYt5TmysTocu/s
qe56C6XIJTELgvxVrJKfheNVa3td1oW4CUfp5klREWLlZ02xdQgIEYU27SL24YODEsjrNweoj1SC
ZcLdY4EnnLlvo4iAVHSdE8QXIGRwqaLFcgtRUAEJ1vWCnyOc4nUjBrcu+0Bo9PH1XmxBIVxdu8hZ
oXmrpkay1Fjd2gzDBp3iqhDgkWSF37HzxCucx2G6Pum7v+dvD8s5bFfC2HjyYJsgtU9OrNQWc296
TmG5u0+tJe5ufR5C//h+ZO0VCZqLQDtyaUzn/xxePy4txYy/g4A7TAOeMY3qDntEp/9fEDtmf0Gn
GMY+pz7FheRfrikPMDIiUvIIzW4EbtMEzrbeDkZlcSJ0sUfq6oR7qXFvJE9JMvIyeovJqr1TEqWI
F1Vnvv+wDmp3kuBXVOLcK+gEoMHOfR/tpO0EMulOXQp1tFSyI49hKxppn0jfuUmnSKAv0Qc8wsiS
UR5A0iNH+qCQj/GB0OsJIPzzFTNeAU9dSvttKNa3Qyt+Jg/uw8B1ciYPd82biL9MnXXF4h0Mlhni
bUhrwBa/9oR2Xh1an7VrK7CiZPIXJ6bNYl0q6qG+jXRYfbEE36CVAWSSz3GHzN9xlyH+gxIJt0mU
5PBL/icuYnoh2VwESoZpgECmzziti8Pk9m+Vggli7ip54Tjq+1tU3ocbiFPgKX2odh5S6MJeksa3
SG6uyDWZAVzjdnA2RQJOXPnuMNDYDy7f8iTEE7M2gl2R9yOfmKj/oCu6X+S9Dnk/v/PgDcwc5DgY
6piEYEYLik0P9Erdk1jnuLyooK8N6SaVEbSlG/Cg3T9D7j39JOXIFAW9KROkY5SjvErqzlQPuoO4
Z9rjEehc3D9GLkZOSjb1xtsGJIsO08AMb4mPtnnOd3z6ajnkjGVboqKOGLQh9sZsfiFjJS0qt4jm
DvMd01fZ4hpdC2D8Dibg3k2pOfTReTyVwjN3YQk39GIJL5kfLfnHqxnQjSEUWt+tC3vk1YuXX4PD
g8urQgh8IsTl3AMtXNWqobUmUv/0gUlSe8AyVfjpdl1IGAhYhu8ycJwCdqiVPOA5dw8eUnUsv1jy
HKWC36WqvRxzXBirlqrXK4j3CAXxSjot1lPVYd2oMpXON0WTsi3LgbT7K42nBi2rmns4P67YJciH
N5Vc8h5VEb1CsBsXG/ocrXa6ase2q7HcxviUIIP36/VMipNZDYL0ZmXKcCi0UuiPmeYGqmB5zpK/
BBMSwK3E+IvOohudgGpbtkwmqE16vDwuvOVz1AmPBnps+F+KvfA0X3Zno4beHB+691Gf9rEU3j7x
oMGsY5ClZz/bQYfb5DhK8oog/PlWBo4+mUtvE9mBWXHqur+DcNAAIgTldpypBb+2GYm6vZxOEWhO
qnPZwCzn0m+nkhUWQqp2nQQRd19InCjB3eFoEIvEkrGIr7opyMOSLrM5Mhv3+YF0bs+9f8NBMsSS
8TY+nk7QmggNgcSGs3gGA0ajVawLHVQhw7T82dZYhvh54S/n6CA81KejbsSUZ7smQHGd3SVvU3Oz
6nOLmLaN2HsqAEVkqwLhfBZmXgZur0mfNQ+vNWJkv9hnaBvaO9LWuwoH+pvoBhH+dDEiiA8Mpa0k
IOK9UUVjWJwcubkIwhOzuAXpVDWAaj6GksNek/UyXZfFLMIRN4xVgZdCUvI2h/IVvmAUrhHpPB3v
//oQBkNWIjP0ukLcufLJAAVy15y6rdb3An6ciy3SyMaDRDfGmxIsZiM6Dxuv8paETN3ZF034KuSC
txG1Fqj0Ur1j0kraKDdkVSwHI9l1yWhvU0yMNLJhEsQvzaMF68CsfBxMR9gNx8IhI0r6EoWMWlfa
14k7CY5ohWS5rWoLQnPX79cKp4si2O4Y2KnKWfpI9H0rw9wl2rayUNoLoE+k53id7aYMfVERayxt
wj0qtCWVOds/Ka4AsGIhp8wg+RrxdIWBJ/9QT7JUfid141++nAFZVUTNpN9PQdSQKxbYnDswXXO1
VImVbefQEic8OYNtmrKREyYK6UvHcvel7vCrq0yq0aWUP6ZkfdiSUuK3TmSKcuffOFMhZeQAzug/
iTU68aQZS4pmu0MJ2Rv0ojT1cFUYlzVuHxfCMYaZrwX/bhrcDPMscNPuAn4yPVFfRfjwAgK/ZiC1
EU+7bkSokyn44qGpKhs4pwYXb7eCkzOP/VA+FyEcarCAHrePJqbJpYHO59fYT4w1KJgZNJnJNURd
LpHDfnQbFomjYTsHXfWTtFFr7lE9fPZNA/ue8E3EsRttFDbE3WTr/Pm3VnQiG271ERGy6rIWoPGc
5eOFdVmdqQlhMVPjC12FPrXP3Hr7G3U0+h/9W09Cy/y3YL8nMBzv/F4B90BGZtW6SMOaH3el5wi2
HDxDZS5kmYXae7+U66p6oHGtjeQ6j0I9DU0BuIdePpB63q8FsQbqZPY9zuAwAv2AbnFAb9sR8gDH
rLM0EOigrrl4AoPIBhAO4HjlTrYPTVc+3CXsZnOH9Ujqh9JYexY4I5gDH5/dI+JOWbtiSNGJI4wl
ts4Nnv/8dg2jj4uOe3DwNFFJhE2VYXyN8vmK9o50gMKZGtHNuvztcDeBqtG8gigaQhqWmOf3Q3wu
FJnIdRUbtEKxKiSFg94pqO2HCgwyNgCvLPUoJJYawrP0PwQ7GH7ZREasdwaMJQGaJY/USKdd1IZ6
6qqItP888owR6WAyPHebDSb5vZ070i1R3sTOzvSXTlEeIeNS/hUaIrmqySMTK2I5VxoACg+WJ9zu
E0O+IWx31Pe8Ssbmp5xZPhNS+Xcu6uesGPpcWakNux61SL4hX4+MHVN3aeOkCRd2Qly5mfjbUqqb
wk4/HWyq+3XuMsnACfv6b9tHsmeGy9CWY+hfASTc65zLMMOKSKEN9WfWQ0HN8ikR0XdJMVm5kUtS
UlnqMb08cmvph6M4d9ZHxL6HCAWnpI4g6iOR0rgKzZbpxXohtNDAfmyvEpdswXvYZgJ9J9SfbTgx
S5izMj05fzSgnRo6sddzU5ob/2zfJhj7Hy0OhOr1oexWIeoG6d49l6p6BxFN/TUjXQsVddPDXyEP
RkxJXDyTdYWhy33e9NB9S37TSFT/EPwCJnVFSYsLX3zTpaE8vmaDTpuGT5RcxZwKb9roWF6Y/fer
ZCiEF9TIsInK8b7R8HUbv7PBsOVZQIuR8U5rryy/boP6fLMC4EK0ZkC3ZX68SL1+B/eI3FS4tO0t
SWVWpFHkre5V8XuJ0dGiRJR0uXbmVl1WrXjFo+DleTgFhinLisuQpAjbgqkw97kYJCNk8wQyxcC9
8LAsDEw6zFzCkQshbLBVHqZwUCBw8p03W4TkiuQ50r/KncExbbKTqtQXI/q5LH7OeruF4TpICF+U
4WZFqOBj3b1/8plVNTlRpYWaXDZ3ZWboYF3tM7gIX0l2PsDIgLkHCX1L87ANo9TMPbbz9rGiKgkW
fUq8gsx5GSbRLDjLYN5vapkD2JFxi+Uc44u+IdNNKfXG7F5cb2qIpoBNbJakoM0UXe8ELQxIFQNu
LiBhmSVa68GqpseLkSYM7P8zPs3ngh0J1yFVUv0s4aXtYIKr7J+zNpeodR2d5NsOM9NOOZRAahCT
FvF9UvRir3DYzsyvrjOhZvrypKka+GNq2Q15dMOcrIPULniaq6DWWPSmWt0p/aGc6WTd+v8s10dB
1iyBFo1CDw0fNzmzWoyWc5B1947BzRU3gwAEGnlbZp3R0z8VddRTsARLwQSTEzf5VrIfvfccJ3Qz
Yp1FARtGHdxL1o255mSdK405Q/fb0QdqKNZ7WQMFwGf5avNCMM50c8NDgJozy2/1Npg2UrRsAwJi
MV+Ka06bxZhBN+TmviA+eluB5dQpho8cLh70MVdQYknuI5R1BgEAYrgq8SoeTZ2xpNt1j3Kkecm5
iLsSr1NBjLzpZbDNyi/dxjun+PoGLeP7bLFKgCI6If+2v8gQnD0+qTUgDvE76nsDsSLpCsjkKfh2
7okCUucjFLd1DW1si5NrKDmLUg0Itx+xE99OBl5zRrSRq5FLprvGkFjnrNWjzPj4EEs7lzf5M782
YeQ++8u/arTV4sA1CdeOWhFT2g4aXqN1kGMgxElvbqtLJkatrivvyNNOSnE5g7OBBr5L5bVm87IX
7Gk6MqswU6FhGMmV/AePqlpZlQC/084ntA2AbR9EdVhRoJC0trAdnDJbUW5XV8iln7rtGBLWvhHH
VNfvTNRe+2uHG0CZ9nst+W1dcWFkV6CQzTNguvd3Z6W7sqJg2K/8yqUgxD/8l0wwZeGSZxaf5SgE
44QGWMfEfnXXrcYL/WPOBEQzTFtFU9BUBqu3BwqF9WrLr5TFgeXx0lcoMOL/5hSjWVJ/UH9ExSOq
We56S5UzZjTFewq1vM5npoNeHW7MDK0YLA8pikGNnBkf45SoAs94T8UEzdIoZq/+SxUe25N/zJsO
DvNn67PACGfjv84lVci+VGmLuMJ6I6iUmziSL2E7y/d66DfdNal0spk702GV0v5DI2iQhTly7jga
sEB3fqW6x8t9swSJ7vOhbcV0ZpQs4ka1KD6r38NUJ5Kyx6QMskuiHBKivPnaVSeqX8dAgCgsm/P4
+BqrCxhblonTyjKmblp/WSmJ+G5lx9/Q+DI5RVFMMR6t4Kdye+UIp/TT/vJX0nnya/lGKESPG2DM
lOo4OTaTd4llejJMUAC3Ff0dF5e3hHeVXWqKjBWQIYL+dP4l/MozqvuTBzhuHc+v/NOlv1VxNUgT
yS7btgd8IdQsVMUNIABRtQ4Mwii8bgUEuZRLD9STG66amu83AXl1St2xVr52IcDyOaCx16K4Ili7
UMXUrl9J3dJgtWRZ2BLcWJAUN7TCeuw6JIhXy435GVN6DUrjae26GcI3om7G3R6XdQjj6yucvP1t
lkv1TMxO0WxWC4V9sBX9UMe3SbMbnAYlPSgBMAy/aX0hSLjOjbis6p97JnM01dvhk8l77zl/qpU+
K6PXmfKA/HZmXPxBYlxKxe7HHO0us5wfHf44vSQqpNbMJZ9XHn38EKUBKem0fvw138yvUFHgVWbV
So+7a2n+o3nB6K/TDe9tnYw/CV/fzscxP4VJZSRe5mpP2OzDjPP5XQjmMh0sqGzcg5PeqGMR0ttb
Fj1HzOsL3Ct2WNXy6KUn0LTfHnHymuvvRcLV4UdDd5BlJFYjM7P34KV034Y03l0yYnE+ssRi3Mcs
135FjUoaALJxbY10oiFk/lTch9Q0GNi3bQnVqb5r6h7dHvFcb/CsEuvDMzPStQo8Lxy3SyQFV6MK
cp9u5exrYd5mS20cfklN1LFJK2AMkLLSQOrTwxXdvZRzNOyubg2i8FR11IF4J/Zi5+/FpD3tnIra
aahAgZBq/qsKlTvXREV23+aOyXwa9fsx8yO7jVyzafO1uUPoDW1NZl8i8ltZbOs6Nd8fLbsqp8nJ
mdPoyeW4cl8bOUbS8N26QNKc6OEndLc8OCrv1X69uhVW1WDbND87vu5CIs4mYmx4OFJNN0xOXSaJ
6BGAj5fC0f2swoLhGkg2zbdrXxjjlJtOUbC1EOlVP307Zfqy84o6D8A+Gg6mpBWp1J1zhIqT0oj2
yDBrArG9e/X20H0xja4t/FYcS72lzY7PO30JVhNR4EKX5flsljMkeK0IZt8YEUzkPpHWHZBlA6uR
8Zl1lmn3w2mQ0/IXxoroqA1q1VChUwgAWYUetIjJXvxd+Mxh6Ltm4dcKoiC6pp8KkFlsC+/riRZy
EQA6v6HsQwS1eoP0WX4MBK8KM7wbm5BmVeKCmPGXDZLblAmBBcezTxvo3bt9ILr9uWVuEPiiaDpz
Z+klOPpiSTR2E/UFpfJ2moBKs616txWAsBAv/IfjEZda9LgvWsNvKNAImZ5jGQ7GKSdD+l1kHmao
rzxdhhx9S96z3TAdFGpTDU4WFWslvvoYKZ0oTOgSusemnwHZqKoSDqXhdlkxyZaIQW+3L961BEUw
9OgIZSCiWtlfqOLPU3ZIYENydNNm5u3TwMjsPLuFvOmnu68nH9Si70u3KIuQCHeDTom2GhlGqm9F
atTGthifT3LmHWviWTULMbv+nqkvez+gNWngalneyLTJ/77athBusynwDr+j++8CVIi0GnkWgtl2
P2el+h/QEJq3NZHBmKt7jVWIJsMh+XahQErKK3wK1Mz26ncAY2w5HcDQjVn3P2htA5386HY0jT/D
gsS0qCmpK7R2T88MvgoIRBLnq0f4Mzrt0nq6/1oOi+2o36nZq4lnj+eliAKRd5Xu8henHsJh2Gi9
ccWMv01ipVEWrSEewqTd84j48mQx3k2c02hPsp7L1SvANCv5UW1iW+aDeMNILNb6fwAq78U1yLmg
QdhpKO0x7Yae8gcO6kW0joYAKMBhqcIhd/TdAGMZ+lHM+HqtEUY2VWdvFDuun9mIcOkOGA+JTNCY
pStkVj/R1MLAyWvX5+AsiD4nK5HFuoC4tvo+GWogw0OplJhe8rFfgJv3u8ABtSeQELZmxZIfdvMV
I0n/UXsvGNHTJDv4lya4WAg5d26NEb3aZOJtephhhSXnYUcaHE8i27tD6MQVJQXD1wOqMXhawsor
08wpHZDlDK0HZDqshmoIdSPkWQb2aM0rVhEkesxBiyvpXFewT6ASDPK1ELhgoTRlYeHQqg4eS0NE
6yhA9Bs++6ljuexrezSH8oxJM1Vuo0WTBVY4DDRkjUGtH7tednBMj01deMAdIP3cxQiZCHxtLbZS
aqsm16wFAzcc3nF7AcmLR7laZXHBZbfC+0aTrUe72aZztUWYPKTt3Abw8Snf+4gPfUBpX03I7UNQ
8MTTSZYPfzG8oZcHS06mXGox8h6WfBVxfi/qIO/2BJA6B5u/hvl5LQwVh79GQlJX5QGD3wy5rqMd
05ca7jWVhsM0CVXcTJOlbXecFoqSdBHQD1C0PgNB+MYaec2MJrXi95QMlKcxa0v8I3wJzP1OpxIP
Zi3Av5Sy/GX1epxTzs7RCB6dM1INLIor41ohUsgloAfNg0q0EVofbGMJVr1ezvGsFohdkW3s/onV
jsPLkM0F1tyYterKxb5chvMaAXjSbWXt2N9quOOvE0o2utIuJdGTqnXNo6YB9q+Poyfcny9rhNcP
a19Ruksrk22NmJUy2xBknL1Yo9VpAJgzMq/8jAnF5IKXKfq/1SqlUJZFi72DBU3IenmJFTBzEHSr
+DqDYIJVq8ZE1vtdapNEigvZcFk06yAISHoqijrVa6ui/u+CxG5kouWdJIfnDOfHUowBMKsOwrtz
Q1+8GITOZHdNegUGqQEPoyBTt4i/JnoYHcVzN/+ZpLo6HO9vnk1G6rOVQGGXRQQIz34Jir41r6Lt
Er1/9TxtPLsEa7wDnmQEP+wD5fpK6qNwgXzuGLZN9iDkRGg8wTvyXY9FCx4gB1PJKQPMCBu7/HJe
fe/beRIyOGn1L3ZqxQsO2pYjgRV/OGevjA4LAcPiVbGxlx7OWmZV8eKAPhTN5PaIzFuQMSI4ivlg
mY6IYk3ESdIwtjh8IfgFYYCLg3QrwO34c+eNqgCJrH2zcO/bbid01q1HJIs1Af6icWeWedtqoudo
ebaoHmqSc9R6AptLqXkPNR1clgCYXIk3hYmfBnd6HUiVGO8PZEW1PMekDtyhPQKLGwtPpLnsbcn3
XdT9HS1ACeJc9pQfpR0KdFp1wL8woBPiUy25rei3KpXdDQ3pnKr7ElabalYPqSbXaMySvDyouLg2
Y+qCb84XHeXEfwh94MexAHg1C9ykO4Ua60RaPPNN4h5u3RKUjqlaqw0u3mtzUhbfwoyS3Muu4VXV
AKSEcxiMSNQdX8G9kUGR706h/rliTFR1NqNnKUx91XuzG3fXbulJUkxemuJpA3U8fxdBo1XQJH5K
yl9TLmv0Fqy8I1c1gRp/+B5LCNxFlkKYGenC0fzxlYYHZkKthK8JLosqMgPqSiqkYQHiPbNHHZLV
fEJqJyMuJiJ/ZI87+QGikqNFuNwRR6acwuX3Ly/mkZcrVzXrkNt2qZ0mObADC+dpOUtKknTqz3HS
kZ01Mu3ioLpfRQ16m8qha2Jo+dPIWuWZl2sbGEsPbC1+FC42TdqjLjy65ndiLGi9JxvK9vi8M3qZ
NsUYRe8n0fd3H2+YOJJGB6Zj7ZsWeFRStcMTRdJXCMiLBZj297XEQl2WJN6odo/lq43mpre4/GET
w5tDS+ll3EZa7Zqie911DNeybQQczo7n7GBSMhAUSedNn5rw6SgXO2mZD/w9ZmrRRwCaBNEV/3p1
1tdWLBydMLzZ6HdNC7mmW5LZTfp34rzqnF4VJEuLSJT3pVx0J++Dkkb5GWw1BBaTPDh8XDBr56BO
YSeHjzmn9tR7GQatSljt+bZ22e14j1ImAhTc6awzKNErAfhuKIzIlVsME+QKu4CjMtVN9KHWVWFl
lfS2unzJAfv2N19BwAFBs0PbolzZMlsh4oNvxuncaB6KCcbcvsrxCoy1CnOikT0vfTlfMMaAihLy
I4r9AmGms3qcDJQvHSbqTrlRb5lRy7FCH/bHudmr0hJUI7z4o95fyjdMFNZ5jVr9ymdG8ifLTnp+
IYaxoTXNH9BAhHxcmV7FNXI8QGz25BGIMMoOTWxShji5NvPi33vQLLYc2Ee6LtibzCgcd7UYjCv3
srtXIx9jaO3ANJyIAmbPZ6ryT5/EWTyBDpAGvXIMIhPL1Lc+fB7QAufA4+UATxoD9bGlcoy6FtFO
xXkL/RGssBffUF9uQfTpyqKfT3nl71zWv/hXDZYG49SQ0P3y9boUYwoT+6qWwRCk1t/LkmFFZvmt
jLgvGXJfIzWjO24VtYnGerunlZmB2okku9B+oKYXiYVGFdEIupNMHDAJmLeH63arou7fTC5Cn6iX
BXWrv8D8OXMwY3cSGDoIanUlZGxz5l2MKqdePN8LtDlnGUrSJJn64izxY3LJ5qcQO/8oRiULiykQ
whliF4vRIMvlv2D+P9m1l9CTAFNcwAnGEZlE38h59V6mb+a7Ye4HYVadiFD+5GuHshzcPZgOoKhB
dUjn1PczDA1y3fNC2ziuJHFcschutEXZCA7I2dt94Q+xk0Sj544tbaQPSb5PfCgDAvAS7+HIqEo8
aCCy2LWCggd1YZAOnwJAGBKn0/KmpuBOn2hRzw0Jo6TVpVKkIzTFwlDiW6GsVnDEOCoBc6zFrNQE
r6ltguc+/HRrQ/9+4FRnFa4cdk+ZbdIxx5pdAw+RXR89CNVsV2WdrtI2loMQm/C8mveMuuDGEBjP
JfWh6RRyLH9CUSH13e8jlDzt/38cMVp/TIe0wX94Wxppq1dHQagTjx/hJ6OC6tsvHjpUgvtKzEDO
QIa1wmwmESvX7vmQ4J0h78jLKaaO12y7tk1A9hHmJeuwg+2pEvajj7xp1bcOrbm2ZdhNqKXwwqjY
tCxTp/V2Nrh9dd/kUDC05hsQovRwOI7oyBi6Qa3s9Ay3mDnV9ZgH1sLri1cLjI00QVSUxziHT03e
+xh/8wXUDv7hTd014rkncQlUxaaS/Bp8g6I7DPFlOLeCtnk8iG9a1NSjszw+//hcl+9DnZo6HyMx
qBd8zfe46jaDnCYRdz6bWDT6VhsxZj/cIGiBlrgdaOx01SdCyEcENmYQCs3FlL23zBccc/2+o6AZ
pvTEqwL1peZhNwBYMtnQmu863Om0HrVJbw8iY1vp+GQQ6he6/vLKXQzCb+YsY9I2w0tVHrxfe2Ov
gjbstgm4jlWYOnH7yv2EuYiPs/XES/Zdf+mlOob9zlg5/eWH+mCnQBew3kt+PL5/R7VYAGVD24pO
VnPJ5bCWc+pK6n9TdxpbwT4yqsm5S8Tva72Qc00iHOiPPoYM0ewpmV1VmE7TarYJB8wHYD6l7rds
V4NG/nAf5ZftHw+9vyZudBvF9MjCybxJceLLE1kgxWuOOtYe7HUEa4F4mFQUr4xFhSxZNtiUnGQO
i2zoS2ELEc5bY6pE97qwBTul0Nxgmjt9a4NWKjj/olkwPi+4RfpTe7Tju27EfzjuW5b7Ju2B1k5m
3kuvG1HJUdvwYPhQaxW0wm3HzbnDiUu0JY400T/PEr4Jl+DtYuanYPpdySz8KC7hhPSJqwnJEA27
n3s0FSq2Cy/IQVf7V7H97iMIRMldMeZ55VPc6gSDEmsb5gSuu+eTvCcQIO84dyOEF4LKu9DP/lkC
tA+KFFHd+h/TqTWPoxgJcEfIQW+91KXNDWuk94HgfAAb6w5gO7XPcTIMOfzcJ7dxWUWxOpOHq5QU
Dr1fjr9O86+qYhXty4V+f0fV4QIWse+JMUBjyGocQl81xx9tN84kZrcHv5UB/PzREWZqWGnozB0k
QTc6DncZm3CrIeROtf24+F9IStSRUwo1QqB+FU1vDkm/3LH1UFFCbhgwj45amnH1GGD2+V8cGpnq
5kzJd/nYjwBiZoHRG4GuzROd07Wq0crD+jVNWbNII7Ah0XKaGacbxcy8VYI6gr+emt4JmxnzaFJc
UmZczMx18JKrtDOH8kkpD2zsr/pRBYRFNTjiJ7GWZlLDG4UHBPD0i+yqu7fK6btiTbvVOorcUG/m
e14fSh1UWVT8N9LBgy8Y51eGQLwO+0ukdFgUtxAl5lx/mZOAgK/FGmniRqVz55YrhGexdReSziia
0MMQedAj4rv8r56BcJrcOhRrb5r/rL1XBgn6grSWQXNxOdgsgLBIlqHd5/zBFyC1nlonNdDO4hBE
GqXETyKFQNPcRIJlJumgVNpxbJtOS0RbPVYwS0jjekYMOrxB5xdA3eMfzYqsu/N3oz9dr/ghXc2b
cuBp+4jZteJdFLACDlVIZAzQ34ilt0jsUb+p2LefoQA9V5Ig83R5ATAqa6vg+ccPSxI74M7zogEg
RbuJjxnu1zFy9HXIZ+9HeWvfrbD2RJHTr2gpv2hcTsCyu0g9zUsFlmBmNKNwXr64HEA6gaokLafl
AD/MpeVskiiMX7cyXSWwIqvP1oSaX0JHLpMTt/oMGmjuRQs7waR7/rDR2OsX6pQbaZvOCsLDVxW6
4gkcA4sqInnYSf64ZZQ9DLZ3ooRjj04aswJeWPkur45MWAdCzFlb43aDgHvueJUBOwX1dnaE2HTf
7CAOHb9swtp+1XDyXdAxupzyCZ9rDRsz4hbt5Tv+OMsuCuLNzX8OkO1ySFdct51e1Q/rNMmKjyBo
zduz8k/IrxesX5jBAKfigbJ1427CBhu8bwvx5WxronDH+tcWoMYOvqkA7s7meBg4nwReaQjoP72u
UtU9x4YsybNHxK/00ltnBmTFItenB/o1K2Z1rVJTZDYyVbtk8pihtE+NaoPqHIKGIfFUxiOaZHZb
pggOzVKdLDBbUdzRl7dc8XgDxLVmjmR3rs2/PRMoFvlVq+ux4kxP4s0tW89gxHg9UZKTQkV0fxOE
90wSCGPzNJk7lTHmfLkAdkNj9IwOF23T0jSShbgTfx9szR7SQWyL1dz5m5kCPycFZsY0b+MAt3mT
HF8e6bH3I1fw414YmZwCIizD/d55dV4k5je88se86IhGxPyVjvatPxYFJY9nb7w1+0aWFD1O44Af
fEWa7oV1t5i8M0WNb8pGR62lkr/nrEiO5TRFz5fukoIuAKhzCQPMXHyNxJxNH1o25fIF9CraPcce
4B8IRxnwhcl2ZrXlv7xVdBz5InkSPWehSwLAw1Li82tXF52y9bNWZDvK51IBFPr2Dj1Vcgp0xMp6
tpjlzdNkM4PvGpcgeF483CwcbXpDIV5dFjhfKHYV6JVb/zo+wHUJLoR5+3XvQ4nbkaH+m0ENeHif
I0ndkyXpVWtVS1UBQWTo8hp9al8SElp3bFjxfVGodeU5qm9HsYjzjqNuaiylzM8x/y0TFUkLEkYn
coukKEXlaPyoLWfVib62CLX7t8h0CyL8yg9Jmpao96u7qhpQ5Q1pb5cEbMBQm9GZeCEByl+JZJoT
o3wfV3+1cUyUdyCFUObOBhuvZaLdsYWCUBPFik9CNEYdID8REP5n2HPBIcnt74PTNVA3n6nzIVAm
eFJWaV5cvqg4+TOKObMMWRBBqgu4Cvyuz6ZdZk3r7QptS0C254XEunEMmo3mWtBDs10+lhSJtWay
b07qA4eMwp+r4+P7zC2COw7Qiw9mQDPTxZrJx5DHiwh9W6VSB5sUNF+aGL2Mx7fNalalCCUFBacG
7k2CGaJKNGX78UyVMLBh0IOc+Lo8fKm/fIS1ebqViKXP7+XUIox51V4rKkHq0PamAddaNqFAzopJ
q+vxAq/f7CsNOCyYztW+V7FUOve499foXiEY98Ra+AtGOWygfGyXqKumA0/Qilp2JJLZZ+HYX9p9
+qsykrMebKHmFAxyoB+K+yEQurWFMNZl/CSopjRcN3MYbihqhGRGHmJfzT+izJP8JCf/iEWnzBAf
VtL3mvcgZBy9Zv62//qxVlmGeEwMeh52v+EZQNVmyHON7cePik4CWByXfvxTMGNA92XsBiNzQ+HP
HUu0TOvMISshPb5JoD8lL0AmfMh7nX4DQG9bTgaCMM4o+/8s5JyIJqo/6kWNTZfyaHNxjouek3Vb
WWzOqgTZx4sQyNK1P6ExSjRoloPDRboqscq7yRVgLwZD9lB5nqyJ4tqvp/+uzgoXzL2LAfrlfKQk
C62SqnWXlzJnVaC9yTd9XOdeVwY2j5MZHwgpEVyMTUfDHWs4cJLZESpthSX7TdsWmpIosAu7GtCH
yC1UGqPI65xoOzg8EiOUwcMF81iKZ3y08ATrGus0oKJlgQzmwdbkN/onqf/h9HoGKfCFpRly47Cj
hYLAJAZt/OtHT4F6aQs2ZXxYeFxRkTeQXDmdP0UDNa4KpBlY5cShrYN/DLbPANyWV0aUdxbTODuU
7qFm+d/rmGiIuKRbejR/cFjygOL3NNPCG2WZDyjQgdm4sVXNQ30K4Qd4n4ZiZ4AGHL98/Mmve+uZ
+/D5V4nr1tiRqfDAHO+hbJkHZQUYTnXDBwc426/M3nC5WcSWH96ry241LxMF19ChEf62/B7wGQT8
bvTmc9F/lj/+JfNnWEHmfpyvBuRaEea5BWtvh2ksVT0QZ2cLhVpUEmAqBjnzddRnjCOl1TDBCP2T
oP1XUiw/TSPbHFBbSaAlEH9+zEvC2ejjq/Oourrm7Z395HN2bVcjk5lP7+ul9HG+XvE6PG+vSZvN
b/sicgMtRqh//AU0yuI6Lr7SlQuSHTLilG/XVfkWLq6Dh30MoanJwFtEZyFoXQW/E6xlXkTfZPxG
9CVm0Ej96tsYoD+u0cJH1b7HlgyoCmCyTKtNwkkuwklgtQ9AHQjNrdiJRFwwtWSgSogY481UhBJb
p0kD1N2YFuaPfd6RJmyVm6nRnJVcwkgbQ9UWEQBying2AIg52NsX+IXWb3Xn/1M6VZ11XBBhbr6R
8ijRFXaKKWx+ED304gqV285/zYLzmaeUhHQkPKwqyLLs+JpR/uYK8bEDl3ad1+oLQ3BoKCbYMHVV
VPS3BehkeXlbaxhKAgDorAiVUJapDem0GBr5Oq2GUFyJjfnQI1nFNm3Y9eZeho0mPiQGVX6CIfn+
3tXkk4HSFl12PFI24gZyxPBwuvQq/x3OHpiR+uo0gHtnYqs7MxgLSFpL4EkWbJ3y/9Ms6+b1g/jb
mATmTeVuGwGuVjTUe6O2nkcUUIWXJyTywjc0xMFl2dKUoURELSITY3fEdRBe6T1lXYRK0tkTVAtN
+y4yB+iwugIS8gvrO8xlgMFCrG4JQQkO28RyvzXxAN7Cds3hY3l/rgXlrJ2o9wWqD96ewV556yId
w23LZoWpqEVofi59aUK7nokxO1W13+DZ953+2kAp3l3cslVH5lFntjVQNd24yfumwaEviSNqp4dH
4cyPQUQntO/bBhUJJg8J4Ijcr3RYzg9ZxdnbVX0ypWOeBvIvdLdw6EslYfjW/mnDP3QMly1RZTV9
yLVCxDkfwciJbqxq7RO6tWo9ElfB++zoeJhC7WQ6p+4ltJWw7MytigbfSVHk6ea0ZezXa27KjuE0
uGs6a5myxRLKcANDyW+G3J+UJe+bse1bjhd1sl7WI8HZ0WfnJkuf6GiIyjOqicS+YurXurmmkhsv
wzdD7h3QGCqyPQ1rdX2ciWb2uqOGEqWAT+iBKzBPKHVPrk0phD3N4dO//icKjkenSHEXew5Deu4T
Iu4/Erb0YPdwj5nAJvLZIss69O71PNUxAL1sOGZ/2+w6oSXqjusRDuriKqeUnXHJdUxgb8lyeCvj
EG6zzyADhENJojGe6j6wz7Jpa7XU3QST2obaqD933moHWUi2YDEk0ZOoiyXBucosBT7A7/+gs8JN
7XDkWBMw/HOLv6ZKlidzUX+ML3seEZxEqiRNDFVBSFGtvqdFfqE9m8LCzVLqAZEbDnf1+tbu3f4U
z83wBZX767s0GjEf5BvHLrSYg0gf/lJFoU5DdPVSoOAYgb3/TfujIWOmGQZvRNrwMiVDjQzX4z+D
OZqVu6jSgKEjAap+DXBA61O10k+f7RiXwYfw/1ll8jsZKHr+2T5lMUNMPPSkSq9+wk7t1qxZcIox
bn3nRkvUQpkm2og8hgOQqVV/DPgQOe5CWinxG4IPzigMQpvvHQawmMap7yHR6dIbTKnLDt4pUQYQ
pqMwwyd2RjKkweBZGgK0O/Q8Ie9+PIrxZ/BWUH/XeEE5QEvcZnWdjF1Tsl64XXAt/xRBPpxczebZ
CU8kPatOYIUv1rx7Hh2OUZW4bDujtFau8fLRYHWSjHOkXY2UrBpKR3H+G+za0z8qUTU94PDQ+LJz
CWMNSBgNmganomMQvGhAxrh16M4hgBFNsOyrNM2/dCYAuzaanbEl+dbpTJKmu2hTzTvONqs+Qxaz
uvHcQHqZYw6ae10iGe7u8A9sTxt6qByJ3nT4hQ46bxH0wGWkRQeF73sfdWw0Ljj+9LLMbVTQbMKR
zGXjdmfSrx0mu5khX5oSX+70hkXLFn3JgYZAuVJ5hJ6glAYvdNhFNCzXF4t1VT+BUAFtJ54Ojhtv
QMV3ysWDRzKdEQtIzxUo+vXk/e+RZoL2mG7wFSRMA1JTLqapOqhNKfIjJKm2ViPgkwD3OOvhjCvz
LgWkGNON8u9TtiC00xFT5wfExUNMPcgODEsL6yWv8hqkB/9H5jLFvVudHBJ7wNiiB/MKpb8Z6OzA
G7Fl8GWVw/IwXmRyOw71tQOHfPZ2wJ7AjwJGyn6e077zpxhxA9crfAlcAXZmOCKh9q8QSEqNU25D
HEWksJyo/i28K6EysjWPZt8cMOgOnSOWDRBqEMOhmlvRVX2ljGxMvR/Z3x2C/vtRhDSPSbthVe6B
jgaWJAudDzW6o69V+HEDOjEkEmEYenUvTcFuFU6uqkLhBgBC1uN39y7zZvEZBPEt0VNsV/qgiEGl
kXZeW9n/9MVSoEGeaeg3enWtUlP6xJd4hsY/Y8ZdjIZTyqioaD7+opnV3eG+rORQIu32vXy5QaRa
DN7s0EuI7Lrykc53jZfe3d752DWKIMsdw4AXh7362vk5UBvK8mXSLj5rHRD8GcyDXp6X7XtEeDfb
2zveRD5Ls0N/3aoiQX1BxFf1SDpqRaWNxvIRpxP/Muu0IVYQPnsfDCHViLDK2rXoLEOETluECEZZ
K2v14bspu53xPecjsxTFmBSKF8nM6tCIvklxP12bIvCK92XrYYdseoPC7mwAOzs1jJOLK/lDv2A8
WR3CSBh7iGtYHMZuluWv+lyW8CXUScBHKyrHwJGYgX53JJS4CBPR1PyWBCNQrvglqh36bJHp8dmC
e7JZu3NM5YJPOXb+b5ayIzPTnqEg+0SJWiHSgFeQ6lsZvw+aauVS7fXQPLBbepRzwClUMP8QfIqK
FOWLPOuqFT61tElNM/0t37XcR/cVwxS2Hoc2QcWEAFe3Oe72tpILFA1QC0mgJYXFGO32/j8ZRpll
+Bd8tJAtSMEGIntejTPvjRyHL12Q7fRp4+VL2mtvZS68IQb0jXzppQTpNoeY/V/ALXNEk/5zKKGk
aXOtkANGsYrcp0ycgUzQ//T+bt2rIt/m1vYDTGPdSnKYAzKSGfNp3os3JndrVTJjmMvCSm7V36Gw
Y40s9lJuU/vLfdD9MKg3dAxkvvMlXQEAcVjhGV4LJ+Gub7xMSI+6GeDR0Sa94RyOHiNxsgQ4ZUXs
5N1xi+6OEEoz8iBcpJicSpl5mpKR2b2ocKIu6YuZQ15Hb91TiwsgaTXZ0anj3U7Ve9cBV0oI3Q0Y
h658iq8Xhro4hBYI9Rom9XwVLgPKFr3fxOvYAtRe5OZQzCfCPrqSpIqKC83tl6JszcEy/5ihSLO4
NUSHWBhxX1dWrE48KKM8Yqbdni8/Qw67y/xQjJRntD6D0Sl1Jo9rjN7nvV7/s08/szRa/R1O4iea
Bcvg3Cfq6Iysz/To0XK9zMz0FPcVy/oDLt7ilhJwjiYlrlA7XFzT/FSAQfm3fcOA4Ev9EzXWRZby
bHuHEUMHygIqendo612AbbsSX6khf8dUiFxLjTuTCN34fZGZNbYbCIv/cUg9ZI9Sp895nNP8iZq8
gXq1hqiAnWtf3/NECNiODyPDlX/mTa8H4u1Sw2Dk0bBFetkR0uwRYwy6D24hhTE7jumuLH5PCiCd
KcGO5yDWIps5V7OuEqaWkvJi3Hck2l7dXsvK4KGIZZ8PQaxjepq+5S4vH1OR4aFaGL0ruJNy7Nfy
0YjJPAM425C3bylqSeAS4kJ88QTtwmKty+sjzGR5wtQmZmNhEo4COMseYFOR3Ldtn4snVY6cTpFI
DShMbz/F5icJqVC0m8ltts11FCnpSHX62Q8EQGDeHE/BFcy8SQMIcjhnHg8WxmmiDhTNz4bO9RGT
Kt0apwIQP9E+6c0QQ5tcDg5mYmTG8B/A/swphiZtPEjcLx2jff9zo/SdyjP5fNeTgq8QqpsO5Ob0
28kni98AyZo2PGqCE9kDuWGFmlrWOW0DdG5XMabpeyxZksYVpqgdipbWWDJq2zzSj9w0acysPlKi
2gRm1T/yTzm8VJsguOoLGlsxfieshLFg+lrB6cxfuxAcxmbInZGz0nXU0652HU47chyjXLMS7Qnq
G5A7VKQy1Blwmt7LvPaAjoRzTFS/Wyo3R9UFNxvlWWKAcBQXq2Sai6iBom30sk79BbX8Vy5vTyAb
C/rv1zWRvBBGB5TVBwgh4TuD2arZCI/KcNBYfByE8i9bB3TZGcD9RNMtPPtcLammRh/EGKsbIsSC
dQpJvxe3+l/+JndTa9cbeDaosaBZsfUSHySUxre2gkrA0jTx68gTHUBfIP9XkAmkITcunjFUozfg
y4eBZZKEzO1QBZw5Mq4mJLMx5Mn3y4YCKt85uTfA7a1jRSE5TUEs4ykjZqqd3Jbm2UW5sQo8SeLw
cbU5RwaeQpIJ+7ucByYL8aDELNPzc+XKPaYmmnnb/XJEhApW7rwC077OcGoV5XBhcXzHMmI5Y2/1
u5nAgK4XRtGsFLEZk6J3vtBe1FG0beJWtB0+RYWGlef6iz8GFjafsCBGGio3Z594pOUGR/Wx8HcH
MSKf0OxGXIn1c1HpPheYej4SE5OVdnZS/8IbooB4U42jQM1k5DElhkKWth6b7UwnjLCZPbFZ8Eh3
5Fknhm2ZAjTEozGokXxmEgPO0Bln2yaeJloS54O1QJGQTqFH1KYf08F4mW6CGbdkAlfMjVDpZovV
Y+XWKuTK1pQfrOw/11q6YlUDtVWac0P2Nc8OLlxr8qEBjHxtokFdapY4+AZtiBZnE3dDGbH8wm3V
WTBRPer/9Vo7XQAALhhzexh3ywVYHQmVPw4aGkMBQbkkDYBnZjzGlBX/z51iJ7dTDcgHXxPyuruQ
KUfUwwi/at3Bf8cojsP7pYyfOqMb+MXr1lWQWL7eg68xcvOdqg+63s3HeisQMOLq0Ii73TTHX9oE
/bNKzEQvRotJtAG6m+VMjG+YpUy7a0nlRxpcrq/JQHBXeLoyylnYxtah/tM9f1wRaykVEvGjx5c2
1SRLTosKJtw68vPM1AhFj6eB7wKnkjOT6HyQOuWwGms4P9SuQIzGTtNJm1cdiuDFR2PYuHqDbQBN
5a407inHM2jzaoluVr0vgz6oaaLjbQ1Ja6LbkYZ44mH6tB3SJ4nNt/IfAykCr8c+WxQ+kL727F6x
k0uVyWv/yZmqe1pkIWdIhbGzx13eruZhSvJefYi1ct+Yx0wPY/pJ3qn8r6ETt71J/AzLln5kvgYt
llxrDc9kxzZ1Dsf8Avzi85D6DqZv6m8hzAUxrzOQ/HQ/fttBI3IZh7kCSG26s9ipEF8wz3l/lonb
k+v9U31mn7dw/L7RCChjfDSOVWEkzT9vMSZSrpi2ADx9wrdYSiZMrGmpJYkjzta9m1BKfmKWXneq
Bnq5IwBlS6zkNDZrUo20788Xre4RuTcZ/4AZO81Oc6CRqVb5exoPNetzVwu9UJzQsEJw15BGEXxy
hsIUhI7/u80sH1DB1I3ThcnkdkAfEwywt1UjSvqkwfp9J46BFrk3ayMX75swstKnyGmqfKm59Quh
shZRE4Gj+9+hMeDQZXDUx0qpDF4VW9VgobDQwyel71YP/daAdBCZt9d3PZek7CvTsQ4YpS5qCKlV
WN1EJ7wpU0kCl2/ra8Nj3uqKXKdBwylfVHeXGew6QVdoG0cDByArXD4aU7mHfXv+JH/SOoD5nVB6
QBJto4Zosu6Ogw1k98AlVooXgfvpHD2op+8ads6gkE/3RVjxegeotHCRDHDgrD5PcuW2ZPknuvad
GH5oML9oNhO7GkwWAjRxzDwCVUI1gbclU1xj9Qcbwwb4GKvrGJqJ1VTUCKcUHzLkUQWfSn6ZOVJe
GCWK9XD4DdJvUbo6eXPZl3wGxKED3MwgTZpILLJg15j6FT21x0FrUQWBmh/27tRmEUwc/O1k+Arm
e5wDOkReJbDJx+WFuXtx6RwQeqB0RAejPcpSLi/LFc1uuoxbcFsc+uubxuGEJ8VdxRWeYkaqn7Ws
f4CDs7YWEetJZ+0TcUa7Osn5Zol26PQGmfST4IL3O4woZVJLoRfQGiSSLVibezXRDbEVfmIzi1WD
d+r8zGrYY6ftGSXZMWIkl5/JTI4h0Y70/c7Ly9ru0iaRyx4/XMlRqxa0hEBvCBQQtiqkFbkt1sxG
DNgob01k4K33z+NSOiYB0W7TZMG5++B4MS5VHS5Xcqexy2AfGIbHutPs+wJMDvrJx3WI2IiwqV8o
nAZSTxyYsX3Lt8d3CIwsLdI/jvrmkD2m5Cc6TU5cDAx8OUl/fRFTRDyfi3/rVgipT8NEN61SwTA1
CHmEQHEDUs8WFfgSaj35d/PQHoc6OFDvPjK5nDo4/QBCjGbz8CDiYndETj/poVJWbmUcLVQtmvZK
kDBTIioH6YWRLei5tT+90u4O3EWLctVj5Q1GAMbUuYCjBYvHNg0jdXIo5KZfM0S4pOkCOU6wQHL8
L09dfO3BxQalZ48nlOKn1hNwWhNmkKW35r3ne7lpNHlQyi92J7vMC7iM3YW5rVG8U3Ayr90PDw1R
8b/k16pI5z56of4fYc6SlSWKGliO5oNJ5tQsYTfcjcSDg/RhnmgNfFb/9+5f+7kiuFvJaVb2m8og
crh0V1yAGd4RA5H6s95pkoTa8mS617HnhtUwzLIvFikEaYvDOOH7AhSsGSwdgPAvJDWiVRdtH+QT
aqC94bd41TTPwJx/wLb0DKjksxc7TuNjFPQj7ZNcx7ZCTegJg1Hcy3LCZicUVUVYRubM9KMgZL0l
/fW9qpzMdVzpAkkmBrOMulEEA4PXomirpa0VG5ofL0l8NC/X4SlT8YcmN8stl/ACzn7x82d9VDza
mz7eAtYQ9LOPiXXEQuwyIaRz5dMUq6gIF0l5fmxJ01sj5R4qvokeVnNKxXCH4nSWwfU3Yo+x0IPR
Hd3K2CjdtfL48+CuhyUzWu3vXOiSWWW2otduJlBWs/IqfL+gDwOJ4hwO9QkxVH3avhiNkOzZiPwk
EBVg93XfED86dqH8oZyDvsWMrHeDCEsa3GpURgymAx2EWJkDSXi3jsSLGfN5Ar0UQrps14Lt8wJ5
mOr5ygJ2VcjnPPk/1dX88tV77z+mPcZcRJSRUdfcjWXBYkQsPB3O5rlAy1Vf5eSghayf5pKyDUuR
jaAXFh0cCXDbsBZM1l2w2zATvFkZzcjrRnbVPrXVLYpxo3Efjo2WnAiDoP9zPfL7tuj1hI0sYZLO
TdxJhWxVsYpk/KAnbYzJ6YhP5dyDvs5CpyRUcCxERo+FmlQrkihmLXc/lh7iX8VkkvzpwkfmOFWE
YvyykbWtGgfI7VDiSuaby8x8/oBQonKK4/vgxD8YagyFq7nodDOQ5ejvvXh2kNJos2xFR0/BHdxl
o8uGAvn3kb3xAIY/UHKA18Dqn4qbgBQJMNanxF2dsvy7XEy/htu4Dp3wexFBMqGs40gD4nJIjwIw
R5o43Y3R3Fi4ycmt77Aww3ZdmMNm0f++kY6FfD0YJ/U447RJK6Q+eNa8cYkrH5zMhV1Jp4w0y47V
bd2mAvT4qMKe5EyE2hZ07sd8CAhXvr3EA872zSHlW9fDRNkJrSAaJ+IAYk8Gr7T3afX8WJdYanFE
E4nsQCs/Jn8rwQcW7IzkhvkqCdOF+RPJBLtuYNvR6rayPVE4MFNbaoAEpgQbDYio1SK8o6HoJL4n
UmyDk6HnVIXIj23mV+aiywU6oP+pik31oCrKzswgQ9oZ6ICOgcQFuMjtqGlgZBkdr/UAap+anr1h
x/t6Y7w8JNL6nOKbdOVWDkIAbgP3DrKcC2SXg5rc7MWSvgpjEVLbs57tFFhvK3/XF4t5LAynhBrw
uCIuw5lio/kmwwTdEw4M44hJMuOhMDJCd2oS1DIztvsIGUE+FfPaxTuLZuuzEApLhPY6ozHNcH22
ZLpTrZPcJH3VdA2yDcm8i+7nsWOeVj11oIAU+gIdput3Bx7hmdPDEqRMJiYDCargj36PgWl4nHUN
bJW2VV3OI3fqwKO66Us+zjqNoyYhR+VSB2XZC5/z4kEJFXn3lh4kGbBDEuSvd1b6bCX0dZr2eQex
nTAUPoa+JZugW0yK+Zq0NdKeZ/h0izR+gMDsIkptLzuhfIrZK06y9YqU8ojCxCTjvnfNamR3BWAo
cBs6hgfe697S7Zs/6dcD9m0EDUcgvRKGD4bnF7yQidSnnA+UP4kauCUQm7nbTYR01YXqErTMczPv
1/scfxHGKtURir6KfEIIKx9hTYN03fpwrz3Pb1zqJRICAdv3yqS1+vuOPlujmLf9yCDo8O8hycUv
aE/R3ELTroSUSnJpB77xRMrynkkFO7LdIFTwfQasiQ2inbUE6WIY2zAcsFSiLMTlhdNOmvjDP/1t
EVdbseHH/cLm/A1LZvt8bSCc2jFrBmeNp5B6VM2VVSuCH0+nOfDaNfqJz3rv7FtrhaxTp/RzZQ+k
9uqZkdBnI2vuVbk/XIqVU/XRcTjZNm8+pUfCTBcykxYvn47ewmNVGKfOjyMILwnmjhNfymUFRyPp
RpjXHMnnOAHHz2xm2zL45DQALsuL3K7o1YzPgbxhosd4fJIR7uWgQZtkTNr1A1QQDI5S9DfWkpAL
gsZq+iU5VgypzNPJIdJkKiX2ec066bh0Hl4x5RarDU1aKEcFLziyl7SuZBzz/+wx3z5ijPhFhJ19
AsS5Q3qw/XseoYrhvIsYTcPGXibd/Wj0e/izsVNQtIUmVLDxpSDrWIQkctp1gNenH/enRX+n80Qu
873P7zgdBEax5Qtkg1X9EuUK6w1oKOVC0VqQd6TW+8/OnN4DXOVAywXO/0ZkKP70mQADAKoL0S6f
NM1aQA+0PVRu85J9xetuPHBRR2zGnhlfc8PPDq2ohpb9UIEdfT3W4OKYhBv65H+XAg4vhf0lbob0
pUb4cGjOwxh8U6Tibenfx1o3suLyrVp4Q79lDEMCFCmdokti5xjtyJ+BCoXnGlAObBwIAf1elK6C
An1+8+HztUvWKy4VtCV1rD+7zu7ENc/sA8kzn0EaRNIoW9GbSvlNBYJ7ruHo67y9dVGcFL8dBq4w
HLPukwZ5pStrrVvjUEw9CBWlCZYJW6q8OoJVk9GXLKics3UAvhEX6Nzr84m5a2T6hl+Fsbk4Sa/9
FUwr4GUyOd14X9Pd4YNgQgZ5KW2z2l+Z3xx9CO15TnVW+DeAB1FfX1iXG4Z9EBMQDBYscmLxamC/
1zdwOOefk/v/SYnpfNXqCqRbdSZaowmTFBmMZjG8zAezc4rYsP+/4JuR2o3d5hGqEyokFFZIhPN9
YWSCvmYVWLZoLpbIA6/tHXQFZRTtjOUF1xD5oaQ80wShdj4yFz6fR1Qv2XGsz2p6TSwbh1F/+Mq1
a1xANzuoMth0k0sRHhWRahQl8B8WYIH9emW5EG+SZPLS7ZBCb3WVJzIvbM1Ni+30qbUnbxehAV+o
XGGQQ6Of0V/b62iowsmA3fbhtSphQKPFOakEEv2XXB+65rMFPggCJw7SELwZ2wy8OIGd+IxBYJjb
hJOnX68mn/La8c/CEZAHDYFQs6Xz7SLsF3eZt2SmGYuhQj2pAGLCMqLqqUUtrXgZgUguuDy4fLXG
JyftjegRjsVS+Ki/uHY+S7pKubVc34W26sk0XISugBzAirc+PMnrUdxWE4/fcNrxnyHkEDn8upJM
RSA/N/tL15t8CEhNO0HymLTKHgAfSFUi20pNv/nEx8as3yyUIu3aIiR/CJsTyrt8y7E3Y9UpLTwo
E9m5qmMxloE91VRHTG2xlOP+G437346+qGQo7ZgmA1xYoicPGpJ84C1xDs8JbJGcfB6d+X9GA97Q
Idnph0YgXoVCr60IKwkoa+JmNMp17ES6IbhSwu35ZzWBkDziyfRkfCQzrnxuwSwTEnZp1DDLIFIs
SZ87787lVnnFGYG/JTih5f+zWz8QWpkDEm7YLUb6TbNHDm+jpIe7PdkC5LvatOaTxv7W6HSfJtsH
jSy6odgL9czeyZljyJedjN70SVRYpZbkvYEbfY0dXcL8fsnuXs5YuTJ/DtqT/cdecV2aJHBUjIEi
mUPkKOVLSYm7sUBib/udrMpLorp10ZnXCuvsAwylbhmBf8hcb/It9zw+bfmtVXthTIjVtN8eKC7w
kUNnnqZ+I5iwOJQ4QCbRTHSRkU/JYZlfdjn97qhWYpehNQcRyG9pSwdu9NVulO/MZR1lNdIILa4h
qEDqq26t5+GRmS6ueH5sj2VOSyiQTuReNo/41WT0YKhnRtJp3e6LXubGUadr8mKtMp3hgrhBeu4z
OPUyyClr5j1z+AQmPmSaXfUDQAsKIZL3nH63t01zGVxDeKNuLIxy/1nmSaidow6ib6xmTiIFCAHF
D9u4oGIBnLz27mQ8peZ2fZESUhuEYA86GgCGqXHk8MKoKPdqKJYMDihhpe88HZ7iew4pAurmP7D5
ou1Ji1KCEIKO7moOXkRtncxYxwBKnfpbNm+Sl/Dgu6/ctsrIzom06/3RBoe2rIRMWqI/fN0S5yra
1rSsqXruHHKt6tMtPnibZJLwpm6rITr/2CGHTkEiUKaIYdRpI9FQ9HEdhtwsb4K1ox6SDQaW5et3
DBK9NapJU3M94n13TWHyNtAUGWpUkNzw27+ONj6al5nAQ1L4dnDxVHA1mh1QuMZTSPxGiqBHcYNk
k4nKP6Q6atgHCeuPcAAkwImsXbV9nLldfP+XGdPmWZpEJWUof9wsZRNrnKCoaNBRWIKqdTmx6ACO
m18QCDGF38P8PG3BLltGPoVjk6HgGB+NWy+OV+mi5f7Avixi5AXdCtfqpqVEDXw7nsuXypwwvldH
GWtjiTCxnCVOXvyADxyXVkqMByg08E4GNrkQW4z/JTwxhYnk7bUpeLsX+OuJWYU578L+qonPxG/m
7MJYKv/o4exeiez+vSBzL3NxUG7JcZfYgxixgOjKgp6oJReedDoBo7HgHuFRhT6OSJQvp/87NV30
tUyspmSbG7uZd69y4A/gvh3lL8COfU7mOdWJ0FMdQIAGEC1Jd8Bm0JQBmCdKrA93YWjXBAl5Xhdp
E8WBvNZYVSL8gdEh/4e8q0YLlcECpi/tTXlu36Ar7BlJM8dJKaAKx+8SaRhfj5nvF2L0wnq5rPto
uuFaVHEQofD3Tg9ulyOYd3B9/PSCVxnDq80cxs5T8nT5gYJwsb82wEtGZFMTsvyQFhfBxvcJz1tE
HrJU/4ohvBLYz01JMe7NFsh6yP58ovi15VL96AZ4KXt5MZBnIT25pB774Khd6RMlXJyxqXMeF4sg
NdlmtmWO0/XCyXvZXsK/aeXcdu/g57FeoVk9L/6oRK5MTkq8/qm+sJ/7RjQcurpLWlLWq+c/PyJK
08WWDuanQXrmzUImVdker0i/ghPuMFApC7Hofe7SCVccRBbm6kPldhhUoX8YxY6bEtg+t4A/bsVN
r1nDjlFrUjKKwMCWJjx3Fvw/gtCp37qdomf7poGh2N1hK3HdYIuMtCoCnHy4rYlv54FRoD/+PMm8
brJXIpgYGSAF7ITfEJkzRBupVXxvy7xP/DQXRoXNrvXA7SGqXkTsLsauCRLIf8tsZZhRVNv+uE95
MZcdywtQKQINiL+iNyMQvSh78NYxf1pS0r3Fe7t5iWIKHAwz4zSLBNQ6646dtSZm3got7bcsBSZC
1723rOLJyBHCF3pzieqY1efyWltcFoMxYpVGMNQxmXqIeVAqzWsImso8AN7kPTiuFOHZmoJEY8q9
W4GlZrpRFWaLhntSWajo0TMdnpEdw8w0BoqC34ChNb4TTzA/BVdp4gTM+UEwn5eJ/wTxQGvWoWr0
XCE0EmVDvMOBRusdpDXQLBRo7VWoKW7TJBcq+rr67KEOMCt95xFCijo3XR2ikIVm6Vqsr5yaZ5dM
/4GqpzB29/pLScOndUXmsvZ20UnBcDxrlleWJk5chvnJPlnlF8MHdC6QY6P8fl9b9qM2psGXLy8w
PSiSLeBkBcGGs0SELV26Abrpia2zsG+qcLdRF3V0ny6hAXwRpfGl3ik6WGOm90vaFW644Ul0hKeZ
azapHbmYYABr7Fr6d6m/RdDlfMJsQ1qIHwO3yIE0c7iBZoJ0aNg/7Qs1rGJ1i1ka+nwfsffm9w/7
fjNttFyDNdD6GU5s2wITC5wXOx7q4AVBugfJaibnmb2BhUhRVaOFBa+CbHSpIQ4Cdl6V06hHdlR+
YLhXm4BpyoWVvNEtTphSh9cqkvtzywddg3iJbgXp7T+S5Jw5aSBPRQsgJgNSX+8rS8QNhvGMC1F0
ISxAuxZELByxLVBZncbWEUmIVY9T5JBEfsqBxnG0rktv5wHT/Ac+WCslSdVaZJAQqyRYUdgwDPqo
Gt3OJxwmykBWLQSptd14+66bJfQBxIQ7+hfrNOTD9O5pJr/j2M8ZpEFOcE/rchA8AoOxwLbCvEUR
W/49HJaBQLAoyBcjz20j8DvTnmd+i2bFjgvL6oVFUznD44aJ4dAZqK9lf+EDu1l60DGfDG+NSyxw
6lliZKQwbn1DlbXgXmK2usuzVFdEhSUBwc2b8U6LAdqpmXpCn1iYov3w84iHJFN6AdENIxJMXZDb
wX7mYK0JzRpjTvkwxGT/HhDUgxIMoh/GqVZiCQ9sJjk4XL4j46OQ3JKr6IWVwVwbHk6btbrkZv9N
ckwAQLZdv69/TUF26OHUPwpF2hgRL18ePP/AT+hil3nlwbUbHTqaf4ZEqnCB5hl/xPkzhqFKntYc
ywj39vOA2lXfr83PXPMcDOGCup9Eojp3lhG+Vnk4cMIeWAFBUcuMc8QYHxed0QqjfPeUQveCAR6Z
kNRpFHfroGRIESoPgkx3For2s4Srcv3FM+tz3fUz6a/Or3VTHzZCglJ476wIQ7uhyiHvvNjvlCR8
gPnR+x3Kj3l6BFgpoEA9eqgG2oYoeXmLMp2scVWroSTjWZePwfDLPYyko0MaMHSyXD9hdjFYoBKz
OxezKzA3upwx6we4IfbrC95Si1beB4UF+AeRJv4on5LP0RBTgOkNw+m98kepT7cKtrXdie2Q+h27
Hjnwf2F3QOu/K2706xmiAwgmhPdfTWL6LkOPUgaUNRSNkAdmSeP/cHiwk528VaktKZLvB6Xezgwj
4/cWYSBLDLE5PTuJPQt6FWmSbHJalhdIHgw0gD28aRir7VrG3pTGz34EHsAmM6tUqXcuh+tXGd7O
6Omhefw9Ws6ebhtEaSz94lNxzKLqm2PzsHCRmDMkGWDfFjvewRqCAzTRIIMns0MqQ5PXTVJjq71o
MC/bwpLa3IiTBM4kV++nE7OGQ3dKkUtOwwFWU9FzYvH0MmDvMPc9U+O/YKNxbb/hNrvgNWeW0JxU
x0jIgYt5/o3B2gUUaTx6dgf89pdAQyO3EpRz+YH9woXJzfopvITmKQZuJc/Z4euvXmVxlxwICmzi
XZt/amrre34iY/IaAUgsD5qXFmF2CdiJ+hC97ii7T9auSPpkpO98Bvq8S3dSWFPyJbPpXgzwU5Ux
9IpomQ34YRhhIWHp+UjLINX7evTlyUJUBthhO4Z4sa5Wih9VVd36Urk9BttGPjIT3p9rzY5vV7p9
CBS/RQzAzz4R4xiNjfpKVT6KVnT9p8680oPsDjQcsVmcHk+CnBOqNhMfiw4LppcHrPVQ9Z9OEdTJ
sBZqOrXFajixnJSfiQ16skLlvZx1I74HJpjT49czYNmwwmkRudXaxKYMab6MQEeJVwm9kUGwkuWX
kY6jwaKIP+K7k1Pxj9vL+JOZCKlZZNmTKDnlJuc3h+B70LwOkcTUXBgLZ5ZXYBsbMgta+kVxQdHc
2Vig5l+iPYP6uLp6h/yLoFoFNaBPxSHLazRn0Uj/bA36cifv95RA0DjAxkTy7ClrZw3jKu1TnrLM
MdXx6bk8TNYvgkjFfQ3vYsMLgRTbgQXc3rQprh5RV09r1Rd+K4OOay66LB3yQpJZcwzJemE3aMLS
v3WEjbwlkTcnPCGpd/Wm7p65lrMFMcVfotYNR9765nr62B0EJ/zx54i6H4bnHQWMyolh2nycy1K1
5Kc877E0TLwtEOCsgnKFr1FVYwePD8fPFHnYUq5MU9kGdvAPikOa6z/o8OHnrQ/PxZHcQoGtTt0Q
mBlDdomYz5ex7qv1PK3ctFzsgKpCS13xVRryejSgkkFO2mWXFqrnjVFccAxRP0O+EWvZ0g2LcZdT
F0jlam+p6oZG6XgKFTWyZhDThaZNfyXKiZdevFn+3BO80QzoFqRt9tcJYdY49NDoCP/FxekvIge+
g4YMTkwbxIh9dIlJuq9yEkFVn8jVsm/QU6GmjF+Twmct0mDoR40BEoliKxsn4B4GqtDGRuy0Wxzi
RN6PO3CcQj9UapHUf44Kvy+eTGQQ2ui3NhNSUk030Q161lku4DpYhMISJJymDO+cToo+g0//x1U0
0QQqEF1aKVG205q07gg9c8nU+TPJMFBIkM/G6QPh2Y+TF2AhQRkWy8n40dEWWAdIM8Sm0AimbYOq
DMqKGBW9AQNWz8nZ8tjGJaVbUwStB7rSKHBP9T3MKNe+6G9EE19YKX9m0P8kDlLNl5TNUHxIEoYk
mIBEAJl5lxcN0njzffthBxraN4qDoTFrMKjOosgVW4NZBOofWMSn1kzoa/YnzP/yzWnmG3v2svr3
L63Mt6poahFRVixe30NaWYbOnpTjLRoX+u8U756138+NWBy2C12sgQYqKmAZUTngBLOagGYs0XJb
dqQ7EK9xkSX9KI+cMsO2RmXqOMq0ejEm/wiK7VILKA16AOEbFIco/Xgs2cwxczZ8LvAXSSD3aNZC
vpQAYP+HVFi3JwilRUDDCw6Nl4OWTKFdt6NzWkh9+6SdCS4FfMaoPFpUJmfR+o13lpBMIb7E1h6p
LlvLuEweXHFTVhKC4XdSxJFcND8/0t5quh2PcIpBAxq+q1ve84M1d0rsbXz/D1NGG3fJYZhfnNmQ
cFhjrm+AJnVPC7QAsZU4UyLmiB9vW9lKVirX+F0e3oWmiHUkgXgYZ8imz6rkX+15JN0VLi7NoMcC
OWxwPNMnt+ecsOpvFuG/gc1kacIGZCqQASmhK2x5s3tsT9xtu9CjRZWN8lnupcpGAtjQ10NLCPKc
N76P5whxSVZBxPJlDlq90hTKfNwQhexjcCWN9kbY9TYNe0Nh+ero7DwSU8QKN5iNZu2RFfSFocH0
hsuX6uXUDC+Oav+vqIq3jB4yLzWBQ1gCryFf/Jde3vvjLlnRkGfiiK9d/9waDWNeTpkI2E2KuXU1
mmVWITaWTpjnaC9apbIYTJJ+3KipLY3SorfKgKdiU44Z1qktaxw8sXErZMPspiZ1aU3xLsIsu5c7
FXrss5icMpOTvxd5v6xWSWiIR6fZsEIrc64SYdW4HNgdqvBKbR72DyfFw867NL6fKTUDYF5LqBnL
iI7X8qiN3/qyFcPr1AJk0dXjwafgxzt8mNiLH5n+8iKEgBbmBe4/du/8XJ1p3hqxl1C5do92wAbm
Bp4iRNLgHiTC0L9MysrdoulG6EcT0YZMLYlMRIQ/KtEFPqR+U9lPBbZV3PQQ5tRYAxjQc3jsc71r
0NUDkulRDtlC1GK/F4xSLNG9m5XuxbvZpj8a5f9QreTCmnMM8Jfm0VSZ8T8CjWC9mLP4TeZC/1iO
ZNAtJzIc52Fo7dmtbKAOdDXQ8hnQiVPkaD4RtwEXYv6HUFGRRaWlNiy69bM+AIFzFHz8IZTothtl
NsdgJAqoX4BM9IeLqzfkiVfOkX/g9ExJ28+Up3xw6/GrwheU6Cne58KwmJ31tzui2Ycevdl0a8xc
kG4wUDlVZJaXPrtCP9+V2wuuYX5pqPyFx1zTmrNE97le4b0Ac1I+JZt2TFYqmMJ8dqklRVXl4QSH
aERYBHkW7fbJspIs2FEp3WmTagobErwgqdBUN0hN7jfgtSFCDcjupbkXo5t/9D0bi0+7egExLd4Y
Y7sfIhi+KrgzQXRkPrM5cm2C6t2s23CffnNHeZPrG5c6e4+ngjA+ljuuOPi6E3vjv3orq4NpbONB
SC8la63us81xjU8zw7OzZjW/WUgDpgH6iei4iraRIB6u0SOY2+EnYNa7CE7nP2M2BJqaBROp+Fr7
DiuVDFq3YVW/kaRfaaAh+6J7NVv9HHpAwBuqnMT51cOYMaZOnhTXSftLVkwrWP2QTAA7hoZ9DAh7
0Ki8lLsqg3oavkvPpqT5H/rPe6X5asXzMlJX5pHckLTpJ/xWQWfn5RcnkUBNMacZy3gg7yavLv9y
RaXZmaHUFJN7ZkuQ7cLvYZ3fs5PrbapwxQTqNwkTDVER1mQc8QA4o6GNH/KMjXaz8/JvbMDY/q6h
sq6Rk7m03cuzfGAmdeUMe1sK1GeF+yr5Lo+pAvURv3tSFXeHsdeBVjpQQ8Nwzgd/Vxue8RQEUm+Z
GXTBOhUeQYF3GUWdf6ftqMsSKW31sNSPgNa+PYl7/ndWFFtKNBcIHWJMXj0hHZoG8SO/IcyOrp5l
njg2v4h/u8RYMithQil9FWRkIO0OQ2Gnys7mjnjXuJ7ZamF2hMkD8gt+vnxfcMfL/KkXj3QMc3DP
TYMFHH6TgtBXPHUZJOG8H2UgZrQDrjOokr117RbRnZs/QWNaeEquiwyX7v/ByZZT9CtCBj0UAOKz
Pmm9DvHVNvUMOPbS3Mp1WDjhTUlQVADh8jERKvfBod82sAdCmV2jgF5xJozCf6dDpZEzVhGjmPdu
6aWdTUteYOsBbgJ+DxUgYccYIzLIueJozKMLGIr/uFehgiQUvkvEQA/3NYT7zxx65NCVaMKSYIbK
RrGGJhlMJ9T/1Jq1IJrSsiAKTKsRmMM7qxTc9K46q7kDkzg5lDJK4/d2zYIKir072Ba9exAW659E
zoU3uFZM/EzJLluH7LThG06jCgT9O2BgYsKhfT3dWU5Qjwn/t/VhNxgF9Z6HsEWnHnkAkZI0O+cv
ziIu3IJk3LoAs2x0NZ3iqcV+3fjGGUzvphKE3N6uiOBAs+Y74wBCjJC6/XBS7U17W8zl11jpNOBj
aiuWZ03JPD75EsFM07s5a/PHjgQvZAnah3ICpECYZOOE3mEOSe6n7LCv0PDnFTxFaq+WqfwCjHt2
78AxBk26samObPQj5KM+zXpWp4gg3lfn5BrWPtWguYHRfkvkvBteEWEN4OMy1dYyx/zss2hPCznt
hCaEdhxeXCqwozEGHOf2CPJfWhYUBydb78J+0QHtrfWFkARtQe42NB5ExM63cH4I7HJU9WstfWRF
P2FSFclJGEW0J6NwVjbHNvqRdx7h2CmzkBp2y8DfW+H2V1mgY37VW9FpsjQFSlr7WGkDU9JxK9PJ
wPUNTokZCf4C+piPnGSqq+ntMPDGbs49lII7dOmS1MO/1+JBVECMDTGuknVFyd9JjPV0qbkgKhp3
7KWP8HY5XSI7EiFBWh29pd8WpZwvHTJi4epXCZShjsdzbXVvtZ31Pzm6e3Srsgey3WEebfzgq+Sa
XaceeIR4sDGTYHL13/DSKrS6/U5l7uMW+uK82x5/Cjj14mv41kpAi5Reskq2936juulDEPG7fpM8
Z8VQnHjjfRj3fQrhyGl3vX0+c7TurnMZNkr9Lz6braVb2jo1lPebTsQtdO/Db7IDCUnpbfWDcitT
YyfFIMceClew8ytjE4co5bpRz20mdyBzHv/XbwRUBcdtqdbGDNXEaSKDF6Os+aMddUWhDg40ni+I
cUe0QvCXqhjJoOfu+ZEYTjRKZnVAZ16LCiwRaJCE+a1nFAzaCVo++WTx4YqNVdV7NI4ZchRm6ECb
bT+R9Wdiv2tLxRPhsG374nhaYqkFvR/yM6uObigFFs2vjtYIKxM1HHZqhd1xrsmNItiglMJJUgBH
Jq8R69VSKkP8u6oNKEBxajeWFiSLiIub8sbXdclYbZ8IR2ELpMxmsy1hgEEUsdaFuUUujlGjvesb
Yq7Fa5AZen57lsL3NjnMzk6ThCLbtJbbznFWjwMyuWeP4aI4LKSEIyL7JgmuP3GrZI3OX7X3aCBU
lxXXVJVnDNmodMnfa2BhA/Z4UFb4OyquSA+4XI0MU89fP4W/zZf4p74Y9vL45woHupPcFBCjSQif
RprZ+eMRygRVS/8CaaFrXr+GE94Vi+XbbA/tBPKNq1qjFaRPGMTohqA+f3zKMDCqBFaav358MDA/
VNpEuJFUheJhVSBD10zM4Z/DC4kYLhN6PrudpHkUvr3I6rVYt8q0ED2P5kh4Id1TYEgmCdqzpyhj
wJfNv2zOa7DdZN5m/3SoUhEQt7prHmt5QxcG82ewhyTgUah11k65ppgPfwlgHPuZ5CWtGOB5jAvA
dJzNvfa7ed3vswoa1D/vIxXHJCs43F4al+4W6cW79YSX7SG95p1NrLgBML7sOEOsSUMy7y86P+3+
z/t2TTALhURoEmFp9rvtZDgjuSFVFpmtJWuPQ3GIbHugCMEIp9tyN85q1gUpidfw4NqtIIQgCM7h
br1KeGcAz8lZ4y/jXbcAR11/bbUaAq+I3kSB7AtbOD8DkTEerGr/FO63YjHSC5naUMuNnChkSSyi
F/OF5i562znWaumxLBLObkag9xrLAdDgOt0dBiVxQwL1VRKPrtZwmXCToYF/GB1+x0CngUNFxs+5
1R9BkJKmtQ0XFmtn6ANS+ViuqZcX/7ij2CSz5WoMKKl2tQo2F7vZxXZVmFOO8CI5vSaQ9VHJxdHt
wp5qfnn/uq7FDUU+e0MM2OZP5LaQCicIX5eIoRDhQacEPwjqLrC8I/fq5tYUbL/hNiKSWDXdJPT9
tXF47nWgEhNlAVSeKEMOB3Yt+Gz7MZcPYPCAtHMRlc+fTT8OJOLleeiX1pLeJhXx8CBkZdYcMs+L
UYyHbOnfSxmQuygpZaOuHoEC5QMGkHPB54t9pvdcv5S/gfTemdgKq+PX3CzVvQI+KNmKQRCyyaFb
xdMF2wNSMpO4qZxK1HQtPL53GoDDeEw1klTDfWmDoPOM1E/pfMbbOtp6/PeXiLTfM+OainpP5cKc
U36P9ROyjuhfAZcPLVGlEQB/8l1jI8on3YwwyGDafw1NoZLiAFXVe5V9TFyf01YnbdpA0yEpU7Je
6RNptNC8Rxz94UDj+AHu9Q4+/s6z6JCX6eOh33LAlTh2Y8ll2/szHkWD0089ucQf2kB1awI03QxX
hIZu53anzwcHAnLUywkDcWebR+tU4AypsxAH2J3uAONou2Fs/OHIbIqCV13cURqAiUF+TpsAiPHZ
ojgOIgfPqGsQ533Dh4blvjVYNVTqccApb6Gmhl6mJBkFaT8VneDU4TFW2RkD5qLCodg4X2cnujzg
UPGf65KCJG2pstqMgdNuHGXtsesHeBO6heVxsAO+GPKH7yAfYqBK2JonqwaCxgYLafZiVVe5g/3u
Mjn6lWxFQmMAqCK5MSW3FAks+txmdsggLANlWsM6RbsByYX3TaX06u9MG41dqwQy+4D1y7lnrQbJ
Iqt/kfEcuB5CeHzLFmYCgkmpshQEG45iW66b9PKIqaMwHEJPTir71wvgDaNJ1h4s5Vu6W/lC1UkN
mL7yzSYzsN/B77Oa1QAs8fmojmavTwxXlBZVcoxFp5bzMmWATgYyvH6lrwwqlVHz6XBl1SFwdFAw
eRcFcyxZOWt0nskLzrSDjA41Y2Oes90Nf5Fg6YdlrSt1Gnh6pOiGcR5+0Z96bW6wjG3UcFErwXD4
5qUeVX0dmnoEjbvTd1Q0/A6sZlpH6zr0SesEF0ZStDRzXfdnr+86eDGDgIYlunC7sRlqo1LNme1/
BnlfoYA9EahN43Cf5hL1OI8dHeLgN6vHLydy8gXT4/sMthS/hgpbOyPqdPKq2PYNQ9+FQMzMnjXq
1f4fWTdsTUn1fs2/yzMOjV67xX2gGk6xlwsPuaB5gJz80KMjQd1FxJaWpO9xCLHwrls8csmFOShH
gH6aFuiCW4P1Iy9g4llkezhfsvyp+uCVEYjMAsRbfBhbpUMI+QmMZ+orR+zJBnwCKJ+P/gx9aloc
S6ncoF6GfhkhV3IcCiF6cODqONw8Rh5YyRfNi+bnApWa63fgBECN3DJlrWz7Qr80+Mct9uujquR/
ns7EsLtTWCVA4izz+RB14rCu2kAKgq1mvQO1xUJK0NoMQScV2jK7zzZhjtbSfTecEGWdzNAL7YFz
FGqUf118wRriLJWUxRQIvZyj3xqwQ0o2wXpoDiF6jDNdHuevy9K1UvjAYhVdFoxcUlo2Pp6TLbrm
QAu/KOkgzKEu5gDSPNpwCUqGHPZiLIry7NHS+8Y5ay+scYY+phhqCDxfXb1/b478KaPY7pEG82FH
EmQewmIF6i/elZirvP2+/s8DEx5Jzp6gi1rj2HtgevREhDxp5R082urHqaO4S2mbcj7efjGes44e
WhcpBPPNYzZhawV7R5JbhXvH9IvBut6bK8p8o/3eV/wtGrl2geZVt5m3MGBDSgb0542gWPXN0OP+
Z/v3G6NvFKyqCK9FT3SQ2vwVzCnOS8jM2ZvR62YXFOTLkCtmuI9tGmdZRly837kWC/QJ3+3qm0kN
Lncbi9hMYxJ/vl9Cgz7HTM9crbwXs9IZ+IPa1+sN84MayF/bYL6yWYmaza/SbQrzAm60zmVcyiHh
oncmyM95PQi8JpiPoObQlLym77tHqHInMQLU1+F5U0fYFIXTPwJXPaF6lSIhmNXC/3eES2N+vhYh
ZZ38Mk6FruKD+HLTChmzCrICEK60hSeEZOTlEBcfomFAcZ8pDGsA5P3OeALRdjM3EOulU3XNp+ir
DkYzrN/b7ljwZXZdpq9dioyPpeVC2dWwcPuyamI70E+jGMAOipDdM4FMyTSxRRWSuChT44w1/jvp
CXo9xgSMtwEvoMbPgOHutPFuV7Fo1HAKKCXUAAUnRP5dYylQWxaogjMRZB6KnMGVzGt3Tkilweon
MAQNQUJzJM6MhIL+AJSdfHWU0S7NW9qqkf3AXOC3FWfXxU74kYel/zoPOHfa8RnqXnwQSvwwiGFT
W5QDSSWpSqjldmPAN4jdu+Gt8ZzQNYpJkpExYWAseLV/UQeEifsDR3Qt+STsTDUI1LiaMz9n+bLw
o3PyDhoYoo5eGaEBi+ydT9Ao249cA7fFK3wJfwgaDiJ7C2C3ROb+vhIYgk0w+Kd5GhqYChL1E89j
CQpe2Cv8LSWXXVpvKA1Ymr8Syf4qdWc9oCDSVRlpgurT1n2dwsTX3q/DX/KO8tcLU6PWO2+seDag
PUzDv/gP3YhsQLEV7n0LVM0WjSJzG5MiQ0OdSgir85VstKmecGYrdumG+RhOhNHUxNSm8l8RQOQW
9eiD2AD2k1wwkuxD7lkBWZJ/1eAb3d1+zJ7EIrIgOpBFTwRHyIknt01Ve7FWXrpTPEGoeXUZwXTO
ggOOwmB8o9in6MeNGwu8RqIVJBSBgCY9p3OY2Ki4FLNCT1HAMbFrKCFMFV+pvQgglJLdf8tLQTBd
oSyErCHNAQN6wsj+aD9JGvB+DJCPZJubV+JW98zk1MwlDiCNW5Vuk5k8CuN9P2HlU5A0zvam4+PS
RXIiu+HjcePN4/GZYUSW9MR0XJq5dYMIANbONqHTJyZcwvN+5I0ZCZETELaf9+d8X9o+DTeEOTBy
FC8f6nzUOTYNDlMkfMRPTrEmQJ6eJA/lCFYtQBmTdk8fS1bZ4eZripTCO7gBzXM4pWeCARHAMGFk
Mnc/9wBeEfBb07KkYvaifjR4hsBMWr6bbdJui4R5ySPzD7/W7JlK+0eg0on4EaMnHwtaPZeTSfEb
cgfekXhu236gIcp2UMuTLAutBn612j6eWjwFGj/ZSZnYLTIl4mIn3X2dPy0oxRFpEfzbNeZ1FDlC
XWW+3Y+IAf2hXoyFeamy0+awy66Wf7zxXEkjx0sexf8yogqPvE0Frqp6wG1FYMN00Wqcz71zlPG/
WT/h3xdsuWYt9rXtO5R9LUiVAfMkTjaRUf7vcrCjc7OcRqpQTLPk/FQjec1Es8k7ObnvEHn9wb/5
QLGjGd14zjTjewMnRvg26gBxkTXkD0+ZPLoRChdUuceJMeUlpuuhMdREvXwlmqVHgLyGVO9kI4JD
is5lyPO/qCY8VB/kfj0/yqONKNBD/OJemczqZ3vRICiOgSiEp1NypoIwY1/cJ4cSLaZXjIkcrCAy
SHNTMmeGA6gJbgxaI/Ry6piAbSel4ypD4wxxF1ihEMqf9YJmzKZ6fOcrLNAo4/0hOJ4XGNSYLgNL
TRDiO0WRa7OT4VrFe8WILCwFzyDk3dxoWEFuJpWQFqQ5ynVXxUDG5FOCV1VXYYLJ2+xVXDvUW+qH
BJpR6KYF+y9l0bvJX/8w1rRrJJMppaFqiUV46Z4VOZ80A2y3I7MOeP9fq3YaAovevcbACPdJraNp
yz6tcFdhegr+8L4Wqjwiij7bIq7j6IoebsB2RmyJNWHE9LH0s78JeysJsdrgYdahRx4xT85Vo1rr
Yn867Xf9BOFO+wiW09LHc/hYytataCddDjf4OZJSrToKNf9rnnZr9jB4nhwJF/ImjmwJY4bf9Fvu
K1XOGZT/igiLV1rMD4Qkzvx8az1QFTPcmHWf7RN3dPkaoNH2wPYGf3dxYPqBmC26OXh/ysmkQq+n
W5gWJqUfbfJP/lNZVJdOuK8YwGm4pM/C1UvxB/9SoomXNamu/kPOx0weqrLvOO78alzZn28H3+9v
zFnFKJNg9ZxXyzFFn2/T5IRlDemc1d6WmC0B6co1d3JhNOGP/Eoi7Y40uwk5ZtletLhhWdscoL2z
wEghH2evLqrhkwtEPcpcPD6kKwbQNxgQrakCMUA3gFg/YNlUdfFX2MDQO/aaJofLMvWc9Jz7aQpj
1o7sHjgLLpC92AaW8MrwqFlMUqLchk4Of7y0tA66JbomSjpy6FWuSLEIcrSWYDPC74/Xg1pYpElv
23ZY1nkPZkDR9TJZdJaauoKdko0hTDdDLbFbpoOGs0HkJ6E0k/7pZvah1BrEv4bRZ2Taita4yH3N
kDPRPAIiUcrdEexX+d1vmbJwOndDNlGmavnacU7fFioUw0ONL7SzWT1H44ShNZZbv+S2CVnEPbq5
F41+pB00dDdT2e7ltheJq1FSFjA+0hS6OiXK+4xmWbQXgrzg6qgXdGqMTiYFZXBjvrDT0qM5NdDL
hJ6kSK6oUS+rOg4nn4/1sWzTkXvZzPffxeSF4aF3kbEVqiqh77JkmpbvagH1j0sf9t4WP5GS+7jD
nCl3X+jMsJO2LIlHgnFKD+svSPyPZAmoL5HQSggnfeEq6qrFg/KIsMwvN7+l2qj3vT/3S7Bij+HY
GN2IZR4I9esF1GMNOiX6MMA7JD2/rjjQYz+URXEy4o7Jl6hVKhNE4jG3CCF4JFeCFHN6BWBLEP9N
iLKvo5pj06ytxARIzWHtt4gSgahCnqSufVi7Tbou5IsS/ENeESchVHUTJL2rrI9IUh3+a48Ikm9l
vZtq6krYqSQnyNPNt0FLqobfoZW/25GMaraKVMjSjQcVfAThabfU3N/0taO1EWnGAITbp+1+ZprR
Suofz0t5HUEmwvunRP8ZHoD6907IwAcsEtSUqL/1/cbxLri1Dv63ECc+vaZRgkdIWBQxu4n8f/fa
ryWP3bMXPWW7n89YRoJRYkqG2kMyjZtDllpSli1XJ1jzhWAiNBDjfuNvmvjdgO6w3/xNYgNpS4xh
nX46Oa/8TZrllV6IZwwgO1VdOtxF2K2LGtIBqpR2gqk2nzbkJzpDVU0RLqcA8Yx7tfNH1Clj8bIJ
6A9HVMfx+VIydmnFtdgcJPnPc41pdTE27sR93CD3xyjMmkitZPJKqtG3qJuMlT2cWShd+HRbGta9
e6EFSPldr4lVFsrMoXYowGvqBkz+/c6gVk5yldXYxwXhopySYcoc1sGQ7RgsdTrTXSuhKGg+OKJc
P9G2gdxs7kuCNpyUvguQa+6mVaeET22NoVfeb4GJD8BT1QM63JLIZ16q8pFLWZr0NMRBOuQvAit7
66EknuZZjz/BypcS7GbjVHwBj+D45GVUoEnAdl6dsCo4ql1DE0aQomOwEyHDzVUiWC8bhQ8lhnvF
CgSnAkuYwBrosAndAKLR5A31BdvkUUcqEWIu8ba1vVME3k+ec85CHZyzovexvHNItLhVWUbQ3vFn
gQA2DbmILkGvrQ99IO/4i4FM1sLxQtpg92ga1lSB3n/OnPuGHIEZ8qiJqImZRkElBZv+tbCDITCF
p57pA7P93q1qScdCXnxxFkT11CidI3ePQPyu6TmNIt85UjNyM935E55iTclKbyxr+jMPuKv3211o
c180IjB9Jp3LEmb8+j+xrXVnoiB0uPTqZwxwuT62KDdp++huWNDFzQ5F4W4pMXKYqCbmfzBlZZoV
LOIZhQWArP0iQWEZBm6MGY6JfKbynB2t02nqFROuO93U0UxYwC/yGOWQUDnBd4Ok1qlavpigYaku
X7xI7T5msGyD0BZUPcIyWhgckB+egTdTFWcEEt7J/5AmXL7SI4C0jkcN7HuL/NNkgHQqjMUGqxTK
8v1X8DMV8axDl+iUHkfFcdKumEJXB44H9aLQwU3fBjSHIEez282AKPZVnwlyEyt7t6nrl9iTagEW
vaawKaIWrUeJpzi5rx4t4YyTpjx+pUOl92gxPxxdpznAt84x3pChREvsU7mzWDzX80IdmoNeIEdu
h0mM2cBxG+NeqGL4VgYWUR97I+0NQSuz5z1nTfxQgWcblns3SYWB7UgrQw45+B79IGuJg2JbG9SB
9Y6L1VLE0IJQxE18RPEnpmAOJ9/XYnrQgeV+ldfZvEIyIZCzoxSHucOU5IrL4lB/DmZkkRnfLaCf
SvfZtdluKIbiIRoP0dM/rk59KAuK9fpkGp2gar8miaaQO1bCVo3bvUE1lZcOG5HQKHYw248aYOKR
WOVzW5WaR8jgSRBIeTU+Vp7XCRIEI/0M7RHPS/HP5NG8jW81sjFGJePLU4JqxzJ78PsMlAW5SkkT
l2ssZ0gdakkLZNQa8WTR2sxYEZLgss9qFVmt7gehtj553xBVNBXn91PNnnGKp/XTn99UtqE8RjzG
knz7n7S/XQyxjZjV668Ybc3pxpKf+bCSBVb3k64QtzbFy/I//5EJ6QuS6/4eqA/cDyHAtrpxyvfN
0VXgcP0NADKi77V4Oxnx3N7OcdsJ9KEXQHM3hF79FU+qE9TCDKwXts7Y/smB939OXVO3xwyO0OWE
FrqLYkrqr0E0Z0r5FMIr6f/FTA3Hqtlyy+RJYUDB//eE9candO9we4th26t9Dg58K4pKIuWKNr5V
xxogr8Td62Emaxgz6dNkshusgBNHkDnNG2pdHgRBgk5l373TQQTbXYAPXzGqAJj7EsSBdPbfw8/v
fQzhEOMN1juPhxi5vzxGeHlFbRiM9HP8KkAnqhBBe3q421dVG0xGgsryK8N4Pk8K9dUYzpaYnNr+
wgdJhn0tsW0N4aA3A31hSflR3L0G3NS4hUvNz9pu55lN/pXzHePQVFLQvOwEULwEkA6kvIfhh3RT
4yDhJORoGkW4Mye4Zjp4mv7SfJSnfYhzMLbIllpLx4FEg/beNaivDQqfcKnHTKwPCXWgSU2Php0E
Hm0sWDIEbfEfc00Vh6g9aJA5Yq/aZVdcpfQayY60cDJ+dGhB5BBhNiE8jxb2KG2aNchqqEX+VRdR
Oaaw9p0kBNHquOwhFWuimsArGMx4S/eSH2Tmv6mMBH2f43sPzWbuRimb69s4PABZ3LjyMKJnKdYF
opqXD7/bq7ptRNA7G8XTPmljsLPj0264oVia37xAKEPyHQ4A8xrEz8yA3AG0QVdFRSRN9/NnO3cB
6Ug7DHsjxEJ3f9M+MCS9vgH78nMWN/0wI9QVMwBLv5HH01t2dCxZcq4YUb29mcl+ktdqSW8vpeVG
VjGr4urGJzkmukIJUFMtNfMMkvl49lAMd31qZfA/Mpg1rcXlH30xgyfEn0zDbW8+sROgxJ0QziGT
ygRenYZhcSV1Jczivvwn3WSWZ0hiMC7c6k754wNwDBJvhrh57UpWKIiOPp0BRtAu2+80s+YgLdZb
pHG85LhuWscJwlhPvBvG5YUVB3jTO9YAIRLbviJJyhDI8j+v2U+aMOiF2Q225CN0M6H7XeegXiZG
98Sn4Q/i3Oo9Yj+9Vwl+HglOVv6wPF/HwIWiqybXyZryGhLk2Iau8zrs+qCCKK2OmXH20i1UMApL
aUK1oj9gi0/LSofw/1h+h11uTMPrPS0PhJrTNxVLQSw4yjGVTlUNAB+6y/8Z9As8gUElm0Zb8zdO
SnLRVuCo3gBr6GvoJGe3UQBUUv6MFzcejxZv8rFJvcW/pJ77I3xVDnSuL4yTz5/9wp9hHQv4ZWOm
dffNnQMa9/D/j3GunzHge2/9COBH5gvCDAmpqickHDI+h2kH8dfmU9ECgKlwo8KqvulfZR1N7NVL
Hl/O0+Ko73OeYeK8LudFakDCXVxdEOLiqNC5K+UvfDHKecbS7krE3mBU5MN+kO/YAjiF9Qm2tFAv
AombFJ6N+6mJdaD8G+iqRDvU9AT1ABsYxhcv88wHUbgVd90DGkn9N1e2wLK/3kY4NPc9P8m+d2r/
nmXJA7mPJt3sYUKlDR0lALT4CXck/MPX9qLXFTF2h2QIlsBIko4V8aEfNH8u9dxt+3JUin9+WHxO
oyHRFtvjzUkRcEzTtbcweCa+0vZJ2YjbjkFzFI3QPPeAsPh0LzSuqPh5QtjQ/8W//snprgOaoBmA
P3+SsbjDaRaK6VAvUyZrGiTgzUJfegyefmNzBP2TpA9fI9PWqAlUCQJ+b6qTwKr4O9xjESh6g9G3
Qend1djN3sYQM58JyzWunvZzeHXy4LUZV5QRU963pzHkH6CoYaP6i/fYDSh0ZF+jcF+TB+k8AeRR
3kVSLsL8vhuJOin9DiyMqsCLitV9vwtkuNJr18/epswaBIJvoMpUhVrbKIyhVQDhBjsJopE+EwST
KEZUymZxkc09DgmXd81BQ7Hu5fIjiNRr44AwH6AxJ/hz82SAZQEIvQCvTzMqv1bGSEVK0kdXz8Np
9P1/c4IzCU6Y9Tb4NbreMopnpgbxyrFwVi5xLIqb5J6gvf36VUXu6JbYUa3+hpjyJKZokVbcEqqA
44c1zoJbvUp40fAVaZQQt7E3R92YkyXKnWldLiBYAI9CStmWvhCaVwDgZSTkhre668rYq+6qTWNp
49BCSogKfz6W3SL//fTzNuh8rOfVyI+w6ca7R8aUr59e6FMQRW6v4iuyEELvTJ/N5hLRf5GG17s9
Zu9veAWYtYMIFZxExZt4gb+qEn6Bw8u4W+Ev6KGLoOsMg+7ZJHkWzDiJwN2Om2+J//6uVJ1JnJkQ
1xGy1uVAGGYY3yEMuNy1lpZxtm21xxmIYKueZLesnEN0CTIK2+D0qAWQO5iIq75ree9WYaLgPXXu
oRq+7MWb4yL5Mf4zovjaA5dGq/sYByEeKdhhttqzPA7TNmj3PuXGr3az2zV3NslHX319E85PghQW
H5DQn/32clmfB9CNuMKMX6bfFc17EEfIEQBaAZWiED3d4Sdpb9Ujmfosfh0a5OkvQaskEddpnmDH
yUiR8vylIvDOJBskxwZiNM3BEPo8bacMMAVqL1zRos7RsqFpUyqFfUV2kyZiJGm/HbGmCT49B0iH
OJ2ZnrE44OHuMfpXJm4wkbrBFJwU9/ov2LwW+cPOYXDfn5HGpV46Uf3RUTxd1MZJ1eQPIMjXEO9e
LKUz2oKjEMrXxV7YLT00ZmaXVE++gSpBqKcpH6ARNTKhvYAFXaFhaQhnDyBHDKv5jqq9SdJliZFq
qz6Jprhh1mKDw9Kvj4vEzQFYEfea+eHzGsQWpKYmubhBUrPc1Zbqf64VZ00WuwGczAWTt/EbTaPZ
XAgIJECNdUwicrz2+gjRqUvRZNHZ4hasMNDhOE16A0iMBOeKzyad1UU2hnAoR/NGpTH8o4CMif7A
2lpb5UkQCJzkcSOyUUj7cnwalTabucsRY1IpZ6rLJQUsYwzfxZ359ZzL3vHMKODNo+aIZF+2pMOm
m29Ke2hmxEuB4c5B602XItZ2Mo9b7dTfwmzyHCw8KFXSsFB3OrGZ6st6f60DcP7XEgfJh3TFRN/z
j/HPy+H+pB0+4ptPVW08i+J1tBPFXJW0nL6tfhHcM4GaIZAmb0yOUukUplmpm9DYiVunw3YfKcdV
LWyNJ6S5C4uEsxnGmAKv8aIiAr4rboRAC4C/TFMqGyFv3Q6mf+CwbXOVtiCcW1b8Oq757043usYA
N1Ztjas9SyCip1Hx0ZPK3mCZk572rFc7W2UEArMd1lyvegQtgS9miWlJn6K7u8QRYDlWYyjPQUpn
jV5882OAx/DFooyU6r7Msi56YZ5GQ9djM/NKnnzRDK+kh1hHTH/tQTIAOkUOcSlysUCBIur2lg6g
8RVsE0GL30lWTd1+yOyXkAuyifqaPFxaO+Y4vxFyrapIRHjAqcav2mjVcGZg/b2MKbBjE+Wi9ra9
UX9a3MCjrC9fzFCeOyjuT2osYkxLkBoftqCfXjqYPARwwzv4ZLc3TqDhFiJB7V6dUYz3teed2ErY
STpMzTtQlkpiB0KvS4o3c2nnQgcFirWT2isLG57j58YIGMqvWcuxv2aYM4BILP+iGosSBj6slN0q
20mxkvxt2m4zi+7yFxcU1Q+T1seQLjdXQkPg55ByVEtXRqA11qCiQ2L/r/LfnbzmKoRMJAve2URu
ckoGZQNh4r1Eac0vsuFJtLGMEInuVDaxTsH29MwyAC/Qvfl2dhya3/oviojPhgOIhTydzgckZ5rO
7JV1cD4oPF+gePU/0z9jMWaQTO8WbN5MuleRprVFsAGMcZHxb6tg8ZEBDEtWk9H210f4up7cOmmr
PUgEY1v371pi2/I08y3BV8SpZHZy5Qh5tIWnDGG5sunDW4l0QEdYytWw7g0NR//DHHf5GUov4iJO
tCEdxwHGnxyW+sIht4QQ8SUxp1ELEP6U47sPGH8l+VJv5JrmlKMlN/iqgva934IiB35jf6ZCuLd+
OOVon4eGEJ2PBCcGO7jJrc8Xhsm19kastxOXgJdFYVCxNfaV9ParyfCmeCGMCMRCt9vOcNSXk9Ju
NS35QEdeaUkDyv/arQT2GnpwMkVtzZKk5Y9/9heDJ6lkg2z9zHSGSwG5fi8XFIzG0bEEP58PKgtX
4QtfYcOl8Hei4BKXwgVzkl+xv2FezC0MKzkTRN9VfKGEbFJuWQ5osDl/KbCmP8TDYcLhmOlOEB4q
VpYWO2MndFgnQM6M17nMYZvX8AlmO9XbRzZC7rPVZ91SAuha5d8bzpvNESm/2o5LIiKNZ42u4xSQ
qgQRzSUBDxJ3yXw6zpIU7FZw3wKwnpX+cyrv0PQ13tMTnK6v0KTB/1yG+HVkw/TnzKGH8Ar2dL6c
YRbLBaCcCvia6MSm1UjIuqBuWDu/f7iZWbZtctggvvQ14sOm5VcHGQbUlUat/HIJQSo9A1sIfRwO
2btWXfSayORuZ6XnQBOz1J5tJQ5Si5Lma+mw9qyYQkYzzEUJTFoGcpK50kD4mDwTojDOJ17+9PK8
HO5ueFJObkL6Fg+3HjNoGKY2HEYasTPCbauzPwSeO99PMjeor2Kqy9W365j7y5z2hqdv3RVkRiu5
9Ui0Cs9QNAgpzTANwk4hcWn9mHR3PpXag7qIS3hp9jrHBKUT89cgR0EPMpRmq0ILARH+T+d+t9tS
op7buwkmZ12OIvKqWzgLBMLFchw15X8WkVSTMJOJiL7JOt1COtKzJm/6LufgqNacCoOY8iYMj6+r
mD6lLXXy9IAVAjgYi0l5QXqyhCfTiIbgfCathd6e/VEywizYruUDMnzFznnmHOw5rlMi5QvBN/3T
XrYnblsSsp4SD75HUbn9twRmJFr9eUUDL+NpLJOYyuHvIu9G6DvR4juxKWdcD1T4IZFL6gq2Ul+p
RViXFZ59iYhGTUtVJ8jibJBUAV6KUQib2QUdtpsl70qbcNTSj6zuwjVxwxHM+0jtOhTuUgHcMO6B
Rm2IxL3Gva0PYSPO+QHe/DrJqXRTqb+8xjaF4H46Ow3yVSEocP2jzNLKeRKSOOb7j6/IB85wsMWU
20uDBiykJumGdg2AgFTQbyLVttFr6umV7ubTENl5hyyMDnpiNCBg2JJYuwo1cnvxR8zwybrybgZ7
C4Nginzf2grK4mqXHoxHNToYww76I7sGN01CPYH9M/tHbdSG97UpQpPbc4u3QqDBpBZ8Buy/T6JU
jYoYdkzZCa/epBJdz/aBemEDzxzIm/2qHyOWkj6H9x/Q840yEhivSnbpKZLtTauPi3mRY2j00/8B
bF39mfLdHdscCYzLNfQjNQSvOxIWYfSCg7KZOxhOLuGZndK56a47KDmLwjma5QGoFzPo1DEsvRdM
LE8LNKRGppCIB/FcSy4BcEBTNRHOURhgslH3FjWENWURP8DVAZhQkBYZcQks01lbMaimVFbaLEGC
VPF1x7Ruuogv9xBVPLF4+cjXbZGnv+0v1L2RsAyujaKOKiu3DlWiBhdGoLBWddy24cLY8FiVhoqr
yBIDvZgZl3foau9t/TGR11i+9f6WUIjN5o3RQhsJqk36/2hNISw7rl0B0bUSQ+xuXFhAjBvScXCK
7k6H9bQgQB7zbuPz1P9jFDWEnhLnrGDBNSzuodCSanPkW12647V+9K4XL5AvT21mXNVs5QjOeO/t
RUUohRSdXnsKyF929MG1hB7SQ61cGwVHzLDToXOUdOUgadgdzKkRhXoVexStvVDsYMAknPUvvBFX
TWxG79mPUwQB5dXvnW3ibUrMzz7CqAcA6MW1z4NbAIedvvqlCED0Ehz2mY+09Cz7d3XwtNfqBhCA
LXPjEMZ2ErUxRtwPi1+RMo0ZMVzLDbqQ5uT7R8jrjUyhauSFQpsFFSjXTah9rzijZTCUh3tFtqNn
ZqJ83b32r66XwmvufjHFl7VbYhA9yIib0gyAhtJQa/Xq6QD1xcTbS184SrDzDCReaQ2YrT/SBL8D
matKFBng+sXWKBghbuh+gDT0JPLY7hSDOwCXSYBL4DJriuia33WIz8o6xY6AWHG8hHE4QdDRMJCH
wfrrv9PvqqN4ViInHqAu7asY7ZfrXTx55G6rp9G68K3FU34ObAmHcEw99GiVLf3ZBNQD5gD9EdaQ
UOD3Lc0Tm4bdoqrwXV6EgxqEscLv6TfZdSOKllUi1bmMXToWEPIftDtUkBpZlkyBase8Cds6S8AS
g1iqX/y1Ehrh7AHOsehBRohJqGOiKrvsfXEp0gjTbeASj3ejJdR2QHYCjl2o28GDuIA8HB3T40o9
w1oF6Qp3jP5fASPgykZROVYP0wvtWrg39iOc71LwdM4IMdtsvWY6GX/BRfUe4cOnkJCwbpD4TUdO
WDzvLElJtKWKHSO2itZlo79EBdSitYo39DBLlYrhhArVco4vNssr6s6JK3UEX26XrUFPMGp1NNX6
Pqn8csiFVpqTrAerFYbEFMoJTNeKl2k27veP22rmPWCWlsEqDuu4wP5PwrobYUEWxlz6ceJx2U8q
CjHCmxRsVj9/8QZrHbyVMEsBOqUChsKVeIPpJPB5RrQFQpF4VtM0K/sZA+/vz1mrNzo7PH6264Ew
Z0uO5cQbmTtWIqq657UrVxxhc1Wqyg6HTWdh1cfSFoIZDb+EJ2FzcWiIjRWQCh+TXpyFDZTUEYkC
rTgbw3Dt64O4uhZdaHTOc3cFPGF290w/f9329hoYf+uFgyBgwk5QHJ5U2UW7YJ6T+5q1O3QndcgD
cIU1T+1qSPxDTt7z5nms5akquntQNNHHFzNxChr+wvaIUfxXhinpha7pxQSydx3m3ndLoxldSIHO
SL0r04OxwQqcxB4D15LIZQcc8WNtQHBZkmb7V9d6RKfx43gnhCVjUGniEdTGQf7OlARWhUmOkopV
PKumCGP7fqS+z9Jc2VX0esrjUGJYfvK2unDPbaxQ1pLKmuOt/K/zA1jYutJQwfvdoGcBtKdnb2yI
JNC9w41pvmMB7U/IiSRHRr29rLR4t76/sJDcnu9xrhAUFItuRt8y7dEQY2PQJa5apaFsqQvbhN89
sHd7DvOPA1HeaXr5PWDy42RonZzelwvAYjxaCnZNllNVD/6vGr+9ixJYwiPMjz9EHg14UvJp7ZNI
RJZfm9B1/oIEOPDPDqbERH/sT89XvTYUjdQ4uBEbznt8Ds2QVbfHlKYkweospDVCoB2BB6UEmUJQ
wXJWhMylh7r9tjG16hfRHfW/t3g9q9ma+bpeyivIIxddjqAiFCbPfgkwTjql+IDtBQTpqcrU509R
gHdtsQpwobwX2liwIaPMdJ9lpwoTDjGbwrwl7NnPooFGjqYwTr//cbSMCxJwtZYAmHVZ/gVJPVi3
3MZRtTen4lXbzdjYMq3DJwmfjmsE8zFcDW2zrUhIbZpUqTOVmrorIbtNm+y2BWFyACNKFpya2eZc
PeBH9iLoyARHio+iUnYPNSD8YxoAxGz3o3GMGCfl8g4/YLSnhluQ+OJyyQYpQ3CXvU4b7bV5fLpI
jXXyep8gbSomIvYNKEF789sxw5AZLZycywc7aRR9MCmXIr2U4bN5ecXu0WQt9K1PKG/Q0r31n4SY
cMFe1pL9cXq2snBTlG8vYuIu6P+oXBxJEdPlJzIXEDaqkO+zrODpxEnPDgwlcP2O68kH7wU5arQj
ZB64HPfMG5wW2z1PXjrGlnJEBwhyTk4gc6dzuJo2GYXGsbNZ/NMPDrfnMQNmfmtPVWWrC6UYIrdf
NtcwIOuwvtV8cZpHc4kDjyk8hFqwYbdgqHJxIMyCF0Lf+IbppU+KAd4sn99GzBmRe+UbIaK/bQOR
/cnugUaXJYgChtUOf435rbCo92heF0iRSN5c7Gejd3Y4g8/4O1VRd0ord2g+F7dijdi5XO6X9cde
u6hXbUEF5KtWjJ7Vkrq4wWSYHQJO7Yv3dAyhgVt8/XeAzVuEjdMXXx6kbfKVinGNeclAjfy/l5bZ
10gb/zWk3eJBAJ8SfQKTEDC0UtqYxyO1jvEqrYEjTLQHttj4b4Y7ikr4adVtgUZ/Mtx0xqY5JQZw
CjBmz6APe54AmYOmaC/2ngsYciTz2q+cOPVh6rwoL571SF1eMhglgPrGFZ4o0FjRk1RxE0wUZt1C
4AFk6wARbx3xUaOXYuJ9Spm/AIUjbMD0zGf/W6gz3Un/DdAHBGXdgcy2a+vUTyumKb3UCgiT7OqG
eShwbwqhZjtx3Yxs8fjr2yXWNhP54vKHKmhzdfRFPyoMqQk4YScjQOF779IQPaozGiajJP6MqQDv
38LGMRz/rG32jDwvq96TvD6sj6tbdpm0GrGJ4ctfD1Ud6iRaIV/mOSejbJ10B859Y6XB4veHqCL5
EQ0k2/4hli1x8DFkeLZEZN40pwpRvRWO+VhrzD3GLBpmGmLuk/GP0TRewMvV+fRCiaK9A6werT5N
BhDYrHQuezasGemMwdclJOrrsK2gmbFEPXKgL4+H/gdN5d/vVaJzD3NzO0sAmadaV5kz3PHY/st5
uUFHIL83w3X2oUO9OpdihF0GUN71/qypguBTYKi1exZBP4tcyQW+1dBnakAAkkpi1fsUlxHi/Ubd
pJF8cplLDI9Rn7KeRYHGz1LPVdfrjgN2O1/qRux5z5oMdLABbYawxV6wz72J60x5ezZdBOi/5Bxf
qimZLDTFcDthosPpfy+hmEP4+QpWFQy0DKKgQzJS9FDhh/p/nShbdfqUt3vW8KHwQ8gmo0Ukrj85
KhKZIcBcyIXLGiNHPi9MQOCo0yYreKeARhi/r9hCJLsAXDCdj+9eU0Hvg080XGg4JJkU1JzrBkIG
Jy8mZBTNO65YmAi5EvkX4MW5tq+j2ffWSAwI9rIAEq9qtzsN6FlLnqsGDtN2kIOLa172EkYGL2k7
DENpC/vEyru+DHLWX5z+irzricG/YZHwl2pznrBCJkzIvmL510QDdTcHUfEEiJzbAs+hYJztVGpt
IQdxuAhLmBiZStBaq20+Qsfa1hATWAiVq6y8QWvPiMWCIeaLpNy+TqvpFvVhAfSjJu+buVsB+sbd
v+Tox5SvT9PzTsOkZEFGOATLHRQXjDN+Hi0UMErDvvwzsi9tlchFmIfbcGQkA6JInBkyOZTQWDzQ
nnHUQFumyvNlyWj7qyO7/BX+m3pAd9Vrf/egdf0S9BKcbIdcl+xqtkoFYhojTY08A3zWIUA7FYZ/
u0MgCecmf6Rjtt9g+4T4POE381dVoguU/X6GVBoBDBfG4n8BwLij+dRx5c7/GkTWjfVQ2oYhoVLo
TrR5LNaUWtG+0MH06PcViUxQMYXM1e/+VACcqBO9Tm8S3eYJa1L83QVu12n9aZFl6Z9rTRnZtUa6
Q3XIu5la2jpDwdRWhl9NHAYuBb/mj7sxfN+2n1/XXclmneV5xAWSFplwoxe3/QsWwJXYpYMCmS2N
gF+5VfYEJmjsT9Tk17NRmc8plucOawUSAob+A0DRIK3RuGk6ueBblKUenoHN5vimqV5bxUBuvngA
YiATzosieGgJ028qI5ByRHkFZPS/hqfBtex1mSGesAd6Ug6x49qafBMIwylUmntA3UEB0Kvu2CzT
5WhBDHdefJSRJaeql8hmXl4IFUOnFZiqfJALLdWsYNqutRjWlCYLXv8ocBPuVILLw4RfeVEmxJ5v
BLFKxZCPZlRo1eYo6Q72W4/f90tgzBqSDz34HCIGHhpRuD/jXC7pVXhD71lWBWq4mJ9HHIv+mPC9
BaoD3n7Dr8hUeub11uXz6Wc7L8+2sWK5tsrmDO7A9/XiL1idkBP5oLMJpTPLFfDtATaDiE0L65gJ
cQZH7DRe2MfCd2X6oCp2qo5m2PgeWHoTZfICQQEno2+SEESxCHb4ntXrmjMiIBk+svfDRRk3Ue6a
Kt3ay85fwOxGHfLN7EY4/9r8h2qqV1DUcKt79BwNf9yRh9vMI7jvnsFn5XX9YbHcCts9ItpL4uLk
H3F1tLHHGfnxD7CH0CWUS+d+YgjvlKo2A5YFZ7usRLQzNx5hh4KBIUcGP/OgfRtEtddpCMJl661W
9gS6vX39wuUTndpXEPTrpK5kKxNbJkwlB7XD0YYy05OeWikq285/0sLy7owEpxjFbFjfH/BNRmzb
5RZu7lKN82YpyKHR4mDi2aaALbilFv60xcvx1NedtXzD748iRGCCkTjAYOg3BGbP5e40lfi+tL/K
ycCvgDNWp4Uf6QP5M8VXhA+ymVOtuwolS+3WT6H2MNc2p9UXjvjDCc38v6hcP2us75G+fpBUH4eu
x2he7BNArHkxiAy+CVZMWSHpCMjib7l7TgH4BX+94ko3BqipAXBxH0gLaVrHKhMLTluA4MoVxIZz
T7MBhbIVSw/sPxxUIqfBzCdXqoz0FjDjlVNmp2yp0I1igfN/UNAFqI2KNKvn7RAtXZgl4wXzRzUz
JryE+d57c7o58uy1v8pIrLcT+i9Ps+H+lWlsGLl+7B96Ul1BCLssxJLyycVGZfSbV0uyWN7TEJ5K
IIwf52OXdbEOv4cVHbCnI87NIkm+8JEVIpyrbQryQx+zJbkZkFbyjClFUAC6xtrDPBF0NnpZX1Fz
+/rgT9oT9SDmxkMtOp0pSBYv7Liy6W4GJ/rvBsj2iXRvbpXK+sGKKgMQJBc/xwEkp4TqCMKXltws
L/eB6gHQKTxVXYjYBUmUXQvG+au1+g2Wr8jmpeKPHTfZumZ5pCSv4F8IQd087wMg+MBW4CvpUBG7
JBmJ2KCmuRwFuiTPX62UWQTkkwJ14trNPg/TTzivmbreBzab6QFLzs/i5cIsZ0mQsgXbeCTF1us2
7igiFeeXwqd0DKA3GFtQAgfgUfDeq+f8eyMaYBjVgLNRu0tMG3ZCCzrOEo9ZiWIShjn+nBXNYhui
FGnGIr16+j6Cq63DOGSmRmoNZ41WNuwpow6KXocXH2uMypAqebQjDtTnYvF86JD6ZKQYu2yuXXMY
+IjQ4IDb7SAVoTEakpH1Kuu341aP77vfB6ey5W2MEUdCTb/T8ckU9wvxy6uOVoDsdIKKYAAg3Iol
xCrJ7j3wF/DxtF8a0JHzkzI+wRMPBoCJT3Z88R4W3Z1r8LqZfp/p16pHNGYUEd993e4hBKtNpdjd
1oG0ZusMJnpxCEB8xfdoyfws9nttS9XkIYGERq/CsGkvbjqgxfCIPRNIr0/c27Xd1pf9Tz/rgSKa
7SSvtj5i1pE0nM6K3j1yZfPFeGRsesgC9x25C9xJz+GTIDZGDiknMrGUvg5FSJbYve516T/N3UzG
OsIjEqa8o7mayiZRb/slxaHEzM+ZijWdiUNQoQyp72IEcyOOYftjU6UXWOfeha4yM2ZGNzfr7F5/
jbwZylloR6qmtIhyEOLmYymOGneI8IYC4uGnz1Bk8GmXqO+Rgb4ZlYHzW1jfr4ptbJP3jvBx+Odu
iFebnuSFS3aNvWKph/r8n6b4lsPDPhxw+qfzRrB8wTtQeqkUpNhv92LAPnpsrniGsF+nbUskglJI
AybbtqvqWFMWKv8m1G92zBfpn7Yxk2FgZe+t2Lz1Qcmh6tYF6IfTcKUIuofDohzXiMqCnaFKtXKV
Ln03Ihh9axaoRQGa6z7C76c8GTsYgNvUrJKPyYZ2yP22nDupMEJIfZ+GboKqpsPyiJuq5vMFc189
QyHgWmYP7gI30fGNY6J3ZpLAcvy1M0yCNRFQzmAaNMkFsjlUSMZwaXMRBHIlWVlGT2b3oAhXFSXQ
o4HKX2DQVKZ49xAQtmWCXNuAYw5LZvGdqxaRrvbrfZfrFPHs6SEOYRpTMzglHM/utFekfS7TUSrU
CA3b1A0op1QolN2KYFGrm85rtzQKgtiC8v02wQpgRGTXcY+BAAFJhjguf6fm1mampbmBL/MzbmgQ
9Zb7hbCZ8DuG1AnxALtuiSvxa3uh4JLyoAiGr2gJNP2kRLrhW/uDfpNmpylE6xRmgqt1lVYx4EUP
8xP1Nv/SkWchP22EGHM0nb65BcMnhy9VRbsaLI4cvr2zHnFv4QNPu8oDvw3f7rJW7uHrrQTmzuqV
PX2p42i6wsRnjy5YkNGO/C56886Z3WEWhL8yvUO8HFryRLMb1Zpii+8SsJy5sdPLU7nfxnLl0Lbv
4GxrdaoDvU/IZLZ8SNfcvW67jxTXQ+fjcoGVXk7e14gNpUOsZHB+fkVQHkm6CMSMhic4pLl+gqqs
8ZbnszZDwqVyuR0hPS11exUpL2EnlaTdOqx6Cb51c0YLKpdDioMNzUOjZYuob9vNSPwmWUlA1nJ5
TEVP5KLDm0oryKh6ZgDavLl/avY+yPR4mff46hpPS5+M0l6FI+zCcyamQTKzTh/nbVK1CrNioMg8
T4zZKKGtWRINW8cBPIRvWN1J8PfiXX2uq97lTRd2zu96brBDA0V5ktM786z8rG4mYe73xqxPCWLj
/fIOsghkgo94XIboNpSjR1ZuqjCUcd21d5t1OPLuXPkI+tS6X2rKYB9eVq0RxDoriG8i6acA0qG8
NYTEjybiqcq9uCWr3fyCkBZaBux0A4hGdjdcupE+y17wrvgCk5/nFbc07q9olsBBfIBze4FEUaSN
BEl4uNfWK5eZvWfA8RJHVth9bZX9pIFRR7L1QFrnzAHsTNIG7rUUQJwKjpsAMxczYpCL9YBuxtBi
pkouRh1Yh6+iJ86pq2dS2GE25vSK+UKVr4iOOBNhCUrWk7aOL6Y5BzqnIg5nEfQ8AUtppAm8skUf
IQQxEjm8nr2CUQT8eJMtXCl1gfgdhW76W4CmQ8T8dpJVTj06uvoI1XA07irfv8nAbYxLcVtEkjMM
/EcXtyZrYK46THlg5y4q4g4zsvDreqGt7qCb5xczDkern2txtBd/N9xdHh4/Xq8lHHH3ttf7P0jf
gsmzBa76cbIUoRmzGXGvqlIYAxBn1dLJ+UPjWb8ZeJCYkZ7ZaK15C9N0I3vmHkAdbT+pTuwGlGLb
XsqAwjEm0PU4H3o9UpNbKZomC7cynpg3PBO2FlEp1AhzSvIveXjTWUAjvcj7bH/65oUX5sFacrW1
8wJSaZ6Dd7IP04tmqnnfFt1JdJDn5Cj4EDGQNpTGq/o/AQU+Pt8hdlei4Sh0P9yLesWzcT27WcZu
cSmvHLr/UwpgDNxENTt9VGD6hy3XbdYWqmUrGVu5s2xpzV/oPUPez9R3LctVMuMPc6UelMuV8IxS
gCT17r3Yq2NSmZWhfRKmFkVylgap1HJJjGzZwtVVxSU0evQLVlkGxyUDNhe86wHN/+bnu4tn86r8
I84EfP52eyH4OrqJLes8UVF1BUydGhihZMmh9J3oVH1BFrLcIaxoE7Lp30aEXTb+0I9bybqZAJf2
336twiASj8cwQUcv1FJgx3SOq+kitUIlF5MYWZ93dEmrcOMlQS6mwpR5QmQOziOnRWPihwXin1JF
xX7yAb/XCj+BogfgWlqUEoy8BUhSfGCeP7dMToRK3EsgXWFYI9kJaNnGL8QhvBdQzAaHfbnZnBig
rD4CxXpqnIqRlqFY0OkDYWKikRy8OxbR4xji6zDO5w7ywgScadbzj1pwrmbWKwsrAwKunqNXCXJ5
3ZFwDrY7auayy+v9SGb5V3q71/TaTsm6mwYzv6J2+B4FWvzLv3+rIYGJY2xqYrz/GjY+T4pIvzRD
TIWThNd7zlRvPbv5MMF9L5eFOrylDksIxlAXJNTqccm7IRx1UNSg4x/7t5jwckhoGSPw8hPelsP/
bwx7MIPgQwd5zJw8A2kLDsvZiLRIT7TX786TFrKSFZ4KFR3AspzJr6okAX/PsSsDeg/Cv6p6o81I
f/olZfKoStGJdgf4jHsFF0U7+ymTfawcFEJsaDmWsU1XWavMvrXspYZM8NR6QSeUlTaGb7WDPntt
NQK4qP0JNPKRpOeHjhPnJvSt1fcGQd9p6KuSllHESH2IdmZfjlrllqbBRC91ct77THHahWL7h+ya
pCTWv814cM5fKsTRTbAg7a06c1cENlMnhyX+v8/pgA3Ti5DQQFrCOrgFoE88QPZeWzSya6EvauGD
1x1mP4XoX+afnVdiZYIkCF6oOht99zg0X8YPxvYLGFxkKfOuUMqolbt17bvNSpetgeESNdLa8bl+
C4KrKo+GCVDd/9YyBLgJBU4Te7jgYfPUupEBjH8gc+5EkA4AunjTWbRY9XVzFsiJC02t8KRuD1oS
i1LChy4Kf16lp+IM8WVNLtvpIaZdCjLHzqsVPil58VK0P/EEZ6JwL2o8uAYNhwDc2bnLGXzAnMpd
ed9zYurnby8w+kTaKjyDZhRt1HnjiyHDvOwaisfWs9raI9LUrPSgAtjE2CPKUq/5lSA9ZC/jK+L8
UWpCR5qzqmKP7kmQ6EtYhA8lAff/ShlF/czFFGBQ+kvOz7AOMNkC7KFKq8VwxlX8BMvD7iDApaDT
4fvfb0rpsZ4dyoIUfm4p0rLSENqPAY2zuC0caLf6IJT4Z4jIJBXrRfhBwITdyPU6GiP0cSGwVKlA
VltCbfO5z8DTiFZcCqT1RbxnuRoRgboJB7TUxYwGzLezFghfcYcPYmTyQtCzKjK2XAvc1AWDtpOm
dhujXmwIQzpWg/ZVaji6e7ETbf3RK9YntNu4krwuPMcLeJ0cMpnF7j8kIS/mp1FdH3n8SnMLHA7n
hHaTWYfs0aMY9MQ9x7+i3crBzKFXo7WiI2eNiFlvugGiuaHZECMYa6bB0x0FbuKQnEUzip81wVU0
O3K2tNJ0cmyBsDHSOYH/1E03Fv7VpcI8B7ktrpool/jFrwCZpeigAKBuWXF8TGLo+Lqk6M2DJlx7
JqsoM2XpQK88IqjiNmHNuSlCLOLJw2biUilymr/rt/rcgoFcj3jq6kMQ3PhE35k4U1hIpP1XLQdZ
4YAHxENQp9sYUjlf36dLljWdc6gzhWtBLetnxMBRdm8m3T9R65+HFIO0haN1RE0K6WTZ95XFxPU9
XxcS80580XmteLXzditul9F5TZPghKWtxRPS+gxkdtRCJryvFwvQRdL7gESUIg0TEzNzy0zDJrx4
5dt0VPb5BsQrmn92M+KfAKra/utLIlPX8sRRY7VHd+eV3Pn4lY38zFP+y/UzTCeRcpwCOhr9lVvh
fSVtEs3XgcrKXbYF/LXMFM9gl7AzcGEC4j2zDDlhfb3MJLGLIRnWUDNUxArfeS7mSbr54ZG0YPK5
ca7lT/k0WZrYA743Rj7pKsD0rIeBrNjVOpepxHk7PcVSfjZlr+Iu1zFWaPmjBES7hXcqTjOkpJPT
uDrGOd41PniqFc7trHX7zhvTHfhtawi1RV816uBSLulT/9u0fE8XOt3mlX7OXyzjrOZhZ9Ff1jmZ
Bzjb3rAH86s21AWxUN9CleyEfkg+QQHLQtUSpdthRBSBpsTD+iP/aAUaJVHgo0+BiO0lj/9CQtzC
NniJP9NsWudJQO+Gn0cCKgjqU0ViAnDeek1gLzKVWY4So+arPRaLfzvmLDxfMvSGdwbwNWY4A35q
01cFJ0lNtwDrlQ9jND6jsNqWnbYxEMAMhiW35jDBFOVrmGSnfaaF6F/pkzWsVF1vjsd/1c0hXSKq
QuUAvUdhrRllzTEVxQb4Au0ZtjXOCOpQcfCcYkOcqTcoZaolejgMkZImJeh5Xy1XWeNYxb4cyzK0
yhzxZZvCoYv7mMhH3yoowUI2TuELEFysrS/+ro2Aneaqo9xbOZ6AgWZq3vFHzJxzqq/0NYRF7i65
kT7XudYUcOuzYZJ2+8OJ/ppcXS7JNThnEpFt7cVarrv1A1rrxdbCkma2pRzGeXDK10U4HbytzVr5
U41V0YuThE0J8wcdh7ZGB/ADsu82AbIz4ZiVCb/XBmzqrOk+3GX+5NuQ4NpTIZHLo6iPqc0/fYwR
6qvaV6Dtkz8SF9kipsEzkQ4fSseVi9zFNtpQSYcLOZZFkQ0atq3Az8d7c1eZRbwN7LnQQjsHvZNv
OyO3L4YFsduPweXTm4qXF3Yxog3I8e7skGU1jWvQbrB2P7uWwJMoq7+QKISrOtsYUOnpPp2g4eCg
A5ny/pZtOv5eGZZWOgbSHgvVhaoREiZEdt6vuDo9moITc1SWOmhCcrXBcTsNuJaBMCJfTBD7AB4j
ksJ8lDk1ve2XE0LBu7vJb/K4GqVbVGbsIsFYIHAU1UExITZ/jjjsUw23nfUgB1HgSq4GQ2SNNXGA
ILZrBrMZfSSz+KIV7b95GvUlOAeWd/ZOu3e+6V+IDTeX7uMNpp2p+HKQ5vRIIfYqtdR//LpCm4ki
OwQ9EtGn8Ex6JE6jK4qpGKWICcKXHyHPe/uBgqZAVRR2BBSlvo4NdzDEg374mkqlbSoKiSBAWiTX
VglH7mhl1GaTRDod6ZI8tMWvrjvK/od/y9Am5OuOXVocXVU0kUJ7wAhsQY0YGmrDoTSoQ9LpbsDq
t5z+4Ff+lXl68fArkVyGGubHLGAqV298RkintoUXQpuFX1yrLwlm3PLqAF9Y2xCux8uBmXML7JkH
TFswgYJxFEC1IH4OO1jMrFPrhjkvLY/FlbN/tRyxDKlBChDUJ87lJqX/m/3U4TWdKAw1XBLUuw8E
mmhhMfk8wCmTeC1T6JJ3KuONq8xc2NneU8d1ZN2SSIy5WAykkDUUGBaZEAZzCMu54l13DPckbRrk
JQjAnMH4oD/BkxswNf0+7ReBSxm76B532V1bzgt9sD5kqX+WwKDexoswSblPdEikt07h8oovpycY
c7ejdRVPgnZnR49CYIXKUEtjmktrK5aosDySajmyL1N3WRohh3h1Mvozbzs4zwrwTH7fweYZ6CbY
aVOBWJWYXIbupYH0d6hpcxl/D1U+7/UhZ34e6y+kD+rVipP+2xHKuWrsyzWvKsxp2DOupfXyueU3
efK3SXWbo0fNEIiHAPK4GwpQxVSTdLejD0dUSQAwlBhiU+5OaAKtfPi8hYyFrtLAw1szB+C2Qq66
1D/QkQ6Bt+kpRHupvLF2+4vMtOTMY5TtQLJ7tB82jd/LKF2Qp6XqC2enOuZF0MMliyOXpGYE92p8
n8Aww+3gYMqe07RB5qxTDP7QVkExzyjD/ROiAcr7bVOpOZ1Id+/lVu9QYDEG4NWnjxsrz9hyAfBf
hkEW5sk2kld7LFFXWut/iA6JOTLOwolUzxIhGSXZE3G/NTql0Y8WcHslURgHyxMfZximf+Oi8q0S
ysbn8sPak0TfMBbJyMInTlDGdmmrY2/Ru1TPcDLqrJDbBhYCk7zrPmz+96KR3GIbMa9VHWnXT3+g
RcmPd7zAu/BCq45BRk0kw3sIoyAe8BKa8NfZ71d71qiYq1yZxM2UHPU6qndbifyvKJruaYXUQmwo
wZLQYUhr/GuYhrnxEB7R3PyUfwwJQ/gg/oB9mjx1ROJ7ugaHBYDDHOmNOegYoKYDpqfOZS3fm1Bp
UUpFUHukinHwt6f2bzpLjabfi4O+Iu0mUGjry8GL0nl4bGoYZFGpo15vIEUPg7f1jIRCNXx7ytA/
o2Zbf8uN4D1MjxYt1ccZP1384sVN+R0b8djkHKWVwoeb2GL1OlYMqPWv5Lj4O7U/Bl5RhJBT1Jos
04NqzkcKwUnizvG0XaXUn9+3X1qLzRsmNIMC1amkxqkCivXzADRBYuOEG5T+cnIO/Ud/2pk7pFuf
bmre1l6H8QggDCcntcEf14s5GRoG/p49CLJFKFUN6usT/0Wap+67VDGp2v8GqVqiSUYd+DC+BuIN
gZzOfewqa+R5OKYkCWJdvOZvPrFDcaPj4ESXrjCghVsx4iXyafs75DFHDS7ajItIX9OE/JQbNqbB
/MNTZTXyoSDUWBZi2qFqUx5LMQpqVH1spAKAcdQNSZrxfX1wXI7DqQIC4iyHhHiPaXM4TEV9rvP5
ouruSfQtxfR7bcV3ueRABLe4hM7UMWyKWPQTDodfZRFLV4uAXXljTJkBhcj3EPPnTNYhf4X0bZVF
C3m+zg2eNr2LjS06ItQJSEfLklNfx1xUS53ZzNuMxYdRUVUZ6rbzM2bkz6tKXQav3Nv7UpmFMKJZ
tKdeerJwdBSlsZThfEx3ajifi77cSFAkVeYbVInUE8eMy+4sNscwOapubApUQuU+lZndSclo+yq8
03NxWeDpyQm73XgPMEsZvW4cxhQoCVVDMTUGS1fcD6BsYVfvNEdoAQ8cWSFAL/FsJ3VC4p2Ws1/r
1oQ+IFkIoLLH69VgRQrrlsaWh6FvEuzTz8NPB7y9p4hyjm5WXZSSHvvNihJOc2w/o8bMC2uGQwL4
jX2DENYWN/RU/xGgSW7FVzQfyEXTb61p4/KR90phR294YXCOtEp4JsVuz2ZeGbzg9Mi+3Y0vpeG3
eMAPphaVfDArkifh30o2dzFrSSCdSee8ucwypnvgZFud4RpAYtS/n/HPTNdl1Tc6+Tlxg9X3dnzq
w04IpJUptn4a2ysHtQJ7pmXevkhsmmyCEJvxMNO/LfD/0l2ruYrDbTIqS2xsozfHsSB7zIUY7p6T
XnlVo2pwD4C2mQyxGaPu0KQoS3UaLp3zawJXNPciJZIOfgsV4X18pMbQRpmuKe4f1HcEgczbJDTr
iFlpR4p2wOWzdm98JPiMVvZ+VW4P3YMsCbyxLP4XNywdehbC3DsxE3VrJOAoE4QRsSpunmYd7BsI
08HzHwtIVJ8uBtcKdpx9b7mpQCji9VGkWnQFjn/RPsR240U8WzSEolQyU0y0ItcFT9vrtTt9IMSM
HlAQOCHTSwelBu5miUQJqSjAIuU8JY2YH4XKmhHtyPt8lqZFnLqYxN06A2EdSzy4In4uZ8LeEe3t
bLAmORN+vJeW6rrkh0Ql2+TvwxXZP2xsmsOhEYFS2eWWm71eZmUJgAyW7yorfLpLe9abR5G7ID7K
lcv/9n+BzbckC50Lx/E6pZPdoCo0Hr2wRqWgJwUQ3C6dZnnaa2R07AViEqjnGlvATTj112FY0BDT
pvTNBELni4breX89vMeArFsPjEn1sAtBXVeY9ksyGX5Ha2ppzJ6nwYIVsIKJ1WCHWi10d/OIXpUN
KJdiGiPcsG6VZBYrATJKMDjQvCZpvEUwjONZyf5ETsc006fTpc9CTpVTDaAKt1qLu0JzhwaVYhWo
s7a2OWNNGJimvVS/mkC+Iohg6Z2mgzLmipo1dp2naVnPPm8xbswWfbTii9C953cKXpkwxOTuRgWv
8oVWW2XtuiwfZZglOc5k6JppUu4fuxcNk2NWfrsPqYotp1ZWQPoAqFalOc/vTADbJebQToPUtbZB
OqYwPTDxkpFiND6bC7EJu8godkTcHb2VjCr8Lj4+GnkIHzs7OshVjEtn4QiqR0+IEHShG/uKdHUE
lixmac6taKflxyNfme8VKp7kknZkN/J4RCKbTHSFnyRCoKQIOgTQ4+qDz4PNzFRBz/kUKaPMx/LD
mFi1nh2mm6ABxPiIHpLXntOwqeCP49jRY5IZ/ItFk8yJVgMgxDeA3peaNLpKYDpyd9Qbxmmx7bAT
jn61btFikODCzvf+TQRDhi1gKUBjiOhrACuSLGXmdMDywonSXSotrve5r447Uu2P1F8rRdszEvBZ
0myeZJoUZvwEKwAxODLGeCq6uEwj6Dmbq3Ni+OMhaCh0p54oD9srY7ZZLXMYBrj9dw30DQZQBXNQ
YA3ejkWbYk1PPzHXRhhsxGylAyQebxcIBZSlEbQ29QNBZ6BjkPlqjuemDXCRtt+m3wNw7DEMm0QT
zedfksOgTrssHwiWWW9soxKWdVXbbLXU6+vf2CFCbC8KVOFkDPFIRjfZCN+mFlS1YY7W2obUh55w
za21nhOWBs4bziPql1ZoX5I4pQ44YmCpLpfJ10XhsSshdkf6eRA4LlNvBGuOE0qcqXYxen+mwha5
jlcDTzr/79QcaS15Pke2eaeR1i1Cv9S8+2dxT905ip8eWx7P6LOt3gSimdDI64RxWAB22eiltYnC
7XgJGtpyrnwPDdKy1dNOEGzgdwmXqaF8QYar4YxUKqxYsy+CLkJA4oJF61bmVoxQ4ctrES4EGIyA
REsqp8hOZG8/DHzM47XmvELi2tOf0aaJ12bX1fxhGFgA/zMu6lO8cuXkyldU051Vc0690AC5iJCO
wiykMRWwXWlxLEiPPfmu6Ge/1YxNOeCHRas+r0yomrnt+wYa+ShO7fJE0xiaYBHdLbO2OITUW+/B
zF9/4QtNefMSvd5M9ytcJ3Mw8mxQD7KiIXVkilvMxJTsCPqjyRBtDIdrIfOelITwkMTRo7Ol0Xcj
gfZUKO0KwfMvwATalIZz2bkNBhl9RgSVxOVb4snUDOhskPR4JnjPg1QOC7yC4j+FJELvvy2mSznD
7D7zD/KU36Dc4DvxfeyVdZAS1rGW+I1ZnFT81jPRcrqpgR57WWWDq0l3emVbLhGxCGsnIjzJN5iK
ef7JZyTJWZhCuZcJ3r5K5HNrSIM1gJ826g+dmTWZqZ/xlus6NTklpi0cVv1RyZoS/m7qVCbtId5S
Dw0yKwD8g01761tSJ56SluDAATKEhNYJUXH746gDpYubcEFoSs9qQixeEQWf5yyHdGpYB+WIh32O
tpnTXKkJqknHCM1nuBaoP3hZmZOPnRRJJYPaH/KN515xapwv/AlKfXRYv7BkBStrvL68/+8ahZnJ
7rZolw6WmubkZ95wNcuhGaB6DySuBR1kD7Thm+4CGxfGZp6mE7xhKq1eryWOVFhefM+SnZILf/94
QJaK8vR9HAqtt44btAv/NTUMG7bHeZ+0KemPVMlLYSP2OkwyYyE/SuTr6pxcgAziSU/mzAYXqy4J
+o39TcFCL0RTvOVdf5Ney02IAQDL5pnuzohFVj/dU+UrlohKZt2WKHxTe5Eacw9peClOjXU+beYj
PmlffAhPGFcYKo5USBSBesYKM+BhuRQpCY0NrGyNO8URwSfNVJjkn/FQ+7E0THtdUOYoyYcNJ1D5
VCnaPThuE6r0HzhTQ2W2alX/knvfNaqIfwVjyxmpmCDxRkgimSDcxJR4uukWTaONv+UQqRtRrA80
djWtDoMNsQy9ngOXc/mOSRhv+F4KLrTTFL4SOQDjlbifX1sdbiNU/DadqipbuMQDzOlWP5eLOeM0
hbzjfQ1or4ngxezinfknAkhzaLLH1x2Nb0AODVRd8UArS3kQDYYH1Eau67tG7pscTgZFJV4Xa7q3
I0y2D+JdNqZ0rlEUJBN0GWwXlhRTpA16Qw7j/prMZGZMscy0Nsgs02dz/KxWmRwbruNkOymWZtxq
u0Y58eJGY3hYg+Xr4DNc3OSakLZnqsUEsypvp7tXRFWaDRkigUMK//99b0W/IqV/isOCrzdhpAYv
Ay+KvFNe3kMBPbIk1hh13hlu0f5WSPdz36jaz3OahCj+rTju3Vxe08tUWaFTIQVwToU/axi1sqeb
EXdXY3nPpZqYQExXkWqOz+av2XiGN7fgZ1NMgX+SyeY/bAjVWikCKnlHNx64gGYqcnW69mW8eYum
+tp/i3hZTvXmZ9b5bDi1e9fILjQ+Cd5yy25Mt0Iythuvmtm+OZxK9LZ4qFR1gLorC4srwUiwDM7k
ipCcMqHgE6s3wqqPAXsCgrdwZHMCxSo6MwkxUqIRocO+afQlDCr9MSwcuqvgB29UebK/BT5Zc3Ft
1n56g/KkJGibqsfQuMG9q88mEOJSyE84Q18kfgjuFLfD7kuYbTBOkbQ3kKUymGlhOJToYjyUp501
/sTnyWyZqCLJJ3a0v82ywi1YKpeIihmEkBQjb3wq5mbcsoTjNA/p2rMKfvnMqHaS+WXX33hYT2X+
Q91nOoXtZxDgbqUt9fl/PPac+lgQjAp42AftOgnHZNTlOzYgqNx2kft9OsmrjsnR30DpNIQ1YjQd
+6vE1tLYia5Bp8+t7A4FacJTxuglV0lZDHW+0cjQNX9vOjjsU/I29QMS/ZhuOewkdg9wAk262yDd
UFjLSB96EUkgbOj0HhuUhkFCXgSbXQHmHYpXvTUyrd9fnvF/wDNbh+840V0bXKkGl4RV+Ao3+3gy
vxh7PhUVjaRNkU8HVu0GCJ4k4F7ZLiBI8qUE9POBq9wzx+1yjxdXbknLaxBny3DrlqQzlTzV6WcH
0P0nJk6MG+HwLVMClqathovfrNRrLER34DCjDsLfC9ZHee5FMdhDX4QzAECBUj1Az5XcY+CNHj2W
L7AQ2Pw1s0XWR4xZudjgl+A0jIJhGI7aWIuVaH1GcyYClEVJsKnZz4DPhESRtXDNlA6ciawoKcoM
fb6iT0xLFRS7uMZH3l5JkU0GNz/bJig5vsnfkULdnNqBhZ3xoiIPx+7pdUAznAvDdwfVOcmYuCEG
DFvsZaBPgy3jQHUvvx6kvKfjqJ9heKu8yXk4Y4ywxCfcqhHnogQu5r/ZqlaCrfdVMYLmwMTmB4HE
aJGiPtwtJl7iQwD4ld7ePU3iUxl1xdA8I1pDbBru93u2APEMk54dfG+IWOvXKqrgJMYwAO9Q9bIx
MD/h/NSmkWVc/lqHjxBkDTuizg0E2RJUPOhlEUby2QYRNMPCAIlQdQ4Cbbhk01F0yeRJ8jo6NThi
4zExBbuherxTKeqdwU4eH6XsrVUXMoN/Y8E0nkm+Nh6cy37JBP6NTydLU4YLdfAYqOUaue/JowpP
nSsPlfTL2TwbBgix2cmaD5BBziBwK7OcCvVs5N1gfedez5ETwFYC1VZduUebvUL8FtSWs75ej9EG
b3p9pOLyLJQKV1/qVF06pvqjkruWsZ4ll0+p3ovjqT7empnEq1KAqfUZOwu8nob4ALUS5Tn/hLo6
OjVN1ULw+mxJ6UnNqvVwifnNIM870ZBxMshx2vSDrzte6+uPMpq0vRcptP7uYoWGGsHFBIOUfsKg
ydAJ7XfuRjGEF9As8vGpJZrFmVp1ejEK3gJfz6104dJKTUNOA8a1V5po0sEB7LqXuCukRkX6yrCZ
bHgKnMS7GIZd4Qs83kOeqzdtZWTVlrY0bAgVrxH1PpQot5aBb5B2n22uKyzdY0OD6HN2PAz56KPe
S8i5BWrVWQFwTpwnUuRLTbNtPWDLvsWq+aqOTFERJOLRz0lmYjgevk3OaarSMO1nxs0ZARhC6j7o
lSrxG98EnTP43/zN6DYNcWZ1rkGRB2ZUefFJHMSBFetf0A2Ak5zyYKM/op1fpFP1CnI1L/t8LSGC
dLAjU+YK9aa1lkHONDWeBAZNgPi3MUx30K7k7gtt1PLSM7AGaShQVG6gF9hZUVN3Md/Odr48wwJE
4a2Q5EHOCXJREzsef54nyXLMkB2RUaXiFIAzn9oN/JgyIALGXdjYasr4MdTJoAh6HBSaEUH17Wmc
zv81ZaWwfkIjkdtu/7hN6U+ZSSVgp2DzJ9Ah2qUkk/5v3Euix7s30Sr17zZYkL/nC3u+mPf/wWMe
djLyUQM2j8evwx3XQ7v0g70XN7ZQpzMDYTc4v9Qb1P0NwmrOX07H0KIxvxp0YOFB+BgPaUHz2D5B
YGA3UgFjK0FgHDIPWiRYv52vLlzlbEnK3W4mOnbRXtIrmzN9XHz02FEFby0P+Rk82KA3fK6sFa0r
P0akxvSVcXhLlaeCd4o1PKi9qWdcatFSTp21lJshrLMEA6v5Z5eR0D2n+C5KM+awm5AyseNVZujb
iDsLD0IK81sniKLPI4/EF4LfFqyG25iQfJ06rbtaOlOQMYej8lfa7DPmarIlcxSjeHpbQELAZmmK
P+pLEoZt7vtyt6fC2J4l62ywYneonJuGXaBNqGW5xsUFyUaYD2LGbAOKYeyZBtUl7ELsF3yUpZaU
RbnzCydEfaUlFFjnMgcWJYzJ4m6Bd2vovy2wjUzyg/kaQJr5T164sWaNaNijh8zbV3cst2PfRffA
enlsFI5tg6VGaL2TL0hpvUl9hkEDnlGUb1JAk3MyNqt/KETIeo+EP3eEyEPIDkE9XcelGkFx/h5d
PkiX1neNGUG/2cfJFPciHQMI4y9sblGrfOA+CQK+UlDg0QgcUzxATb9kR1SqvIiQ8N40MIS2SGXm
XQA5jpRsCNTozUJlnH0HN6HCYLpDUtTVgZIS4iXrBBorI3CBN7jGYGHCPK2o1K3zmZgbUmhbSagL
Y6QtGlRdli4AVdk4tnQwb32gS6JzlrEAKK8F/uU50fhaAJotCDqq1GrMd3JTvvKW+PuNPh69Nya2
fxYNrgY1KZhKpfqt2ph8AD75bjlIPhJZg21nuwdcojFm8BnwpV600x+Q9Uyet7vnpwTuCVUHRl2O
M52HXGIFfuadOVHXCyvOP9CC21voxZLwZQR0T/zrHR9NiBFW0Hd4EsjEh6TvF2yrDIwOcw2fow+x
6SZwzRoikPDk0/4iCiAlMDDzdqPFGyYvLkitQNy4vGu5pEguu6kvwrSY9NxG77EEdTcP+eortO6R
8ehzHdOM0KG/mEsbYAptNDOP83Rxr4Hlfw3968HrKyBaG+g6gWcXkxEkoKCDJddkO0QmreFNP4uk
uxT1w72z2v5ziLVo6ATPrMU0XSRat3faZUS6VrPBNI6TbGPgdDcedIpiQbuPIcE5HOCJ3K/HkNPB
7WjtTWsKAn7KuBWXbDBL6fpujbtEAEXLjOKeccDJKD5zo4Po7JqeuutuWbViMwvs6DLkNnSHc9Rs
hGbItWx3iswWGnZFPGY8afRXb4BB+ixPVzN6lQq7WpHSyndBfgfn8xQzzV5ZUHA8Vg2ojpnsfbkF
gBEQCiletwKlyiGO6ovi1BoT4m9jgbPxe3XqnShV5VO/LRpG4pXRFXtlg9qasdFYgG7LybqoP3FZ
O7NIkIVXqYVj1WbJjVqbjxtsOh7KeV3QstDO+a1wKizdXq9ief84f4j7YTgaHXbmUjO5A2Aw2NzL
oECG67Mn8LDJkhgh2A41o5UYqq0b0IxDn+RPUIo8DRuPW4YM2y1e9g+kLtUtHuXMUCFQOvwSV6YO
nkl7WHWNiHUx2UqCuTjybl1agKH6oyo+UKqTkYMUSpmiTfA2p/OZ3uS+fLqPKFjmXAxGSvmC2O2S
rPGJJXYElKevEnDCu/2uajgXzT0yALw7NyeFH1jTvOSc3o65Yzz6k9y9g0lF5Fb8XQACPMyUyfnw
B5j7CbM9rbZTC2BrziCyKEzB7JYh8Je15Lb9V6Uxp2dh/wIXDe9sBBVLA4WYhhXqKwjKGrw0lfYL
GiK5oZiGHvPo76dTWT76JqXvryKNofpShOZaNIz1RpLnRVCbC5ZpdxjRn9TAdfeLgr1HT3HZi2xj
ttYPwGJwWnQAO0dajjWB5/PMS+A660FXq0isIvmj5qLFFAHg7gWWwshMgvl2Vn28aA2zjQKzITRw
rkv78IdrE7+he942mWfNntwyD6OWA4xKtFmqd8ME92JG6UcEbH4edBKAyJTKs+zKuP48Z3UTYBA0
7ByH5IW0lEVOfQMfbsVKTAwjHJfegAEUHB8i9I8BPRWk2/RfifC1zzmPsY7Crt+8XPpkTLlL7DJi
uAhf5tyCh/jXJQSZ03ZhxeetBdQli1FEZ1CeVeffv1BTR6fNSJxMaqhZWFWq147Bx9BS6n0oXApa
bH/s96z0IayCKIC32AOwC1P+a3A4yeUpCx3105ZNJZm48y8ICjhPWkXGfGko3jLaS9PtcMz6+svn
Qa5RX+rQ2iW5HOyAyPVu719blLrWFKXdEljpGCYOQme7azPQCIoSpB95yekNBWhta2/iiFQFN3dN
gN5qI3YVpFdLHP/A8YHKAvTRjJ06jSRdlZUkRdw7ZLOG0f5wHfqs1U9Tg9jHBJGqHop9htqQ6ybn
FTsCdmNyratQ3JTihmk+lOyY6i5MFBm5FwBqFVq6//fHTXxbbVRtVJwuiCGS5E7F59KlmDFu3BkI
vtIh858SXQt1XSvaRI+kjeuojiYJXvNicXle7zii14YbvPDa/olZfHWsfqPoMEzsqUzDA1qkzb2q
Xw5sL8jJwqkccCZqO5UYnM7DevpcAY9qmYhwiEEi/UQrovdtJs+24a5SnNw0xA6vYtlW1z3QxC7U
LH3DnS5zAopVnEAkxIfFKsyo/bMZ1yDSGzTDkZJt/IHs54OkcqXHR/xbWmQFiUn7bFeHqlGkim9w
627hhaxvzjWCSIcBH8aUGdF5tJvEZR/SX85GY6gygm8XmOribk/nFRvdW6Lm+FkQuZLXnm2SPzkf
gUYVzDZbMCdvOB0Z8M8qwUNW13kg0zWr5M6pqapwpO/TtxEC99LrlQ6TRMIUN6ZdmH4vOslTCNtf
0oqXTn9JQh1+oYVibPyqrzCyC1otWEFfG4k/Cld6C+R/EX79prRuBbTK+3eiK8ICtwzW1Fwin76+
s1Bpe/ZoAei/sxkVFUbNsU72BXZc1/lnGo1wT6x2qUpXEfyP/WE/zJpF9VGxSoCL+IaMxB7UWaO4
qO+5MQA6qeaNGLnT+IuMzkiZzLNG+QqpyLb8nHmCMhTBjXuDbbRgSBNtpoRaxcw5t8qJcYcInLZp
AH+PerR940xwp/e+uLUuIny71Z1EAdj7D6J0w74FMSrXOLCcqvz1Tr164chtKmWEJTp/Wn4ushiW
gTsE6v3XchQGImxHRB1HbaAChM1KPSHLM1SUR6uVio3I5f0FWVZ1pGwKYxPfllrnNnuiKa9cSP5K
/kc7+zkJM5qRHY7r6z9KI8VNydETjX/QY/c9C4b8TU5g7LI3qblgqDnf4ev56nGDhKz5G7tcdY5X
A0DzPeiAaOHdw5t5Ey0NjGKa9CG78UV03jsNllh3SMXbEOviRIWPmE0Y1HtqwSlXyxzj+cF+pfVN
0XZowc4+TXYpFRzfqcRz3vfQh6+z0YQfZimrmHbkn+k/AoDs+garn9ow7mevTzsuopZ7nqtUGHbi
J1lXXTvvWTV4eVTr2FYM0dlyxc1o6zAVAft8j3qlJklS8zzu+FxPDDiHfUc8vbmrS4iEtlEZcXP9
FJ9XypC+ZIKpgsrB+oCLB49JCRXsdb+kFXGFVZXyGhCtn8agk9HSNDVfk7/TzxF3Rm2qY4pxzNLC
ixG3HK0ToCUFYRHGX5/iagKOL+lNV2+2UIWZmukAlyaoACAIryNdt3h0O+xhrDse0JlCb/PFdl7R
cVQSfTvXCg3Zm7dK86B5Dq93r5QnGDpS1WVWbszd60U0XCXJkhFMMYQThh65NPUL5IiQemvl/WuT
lDPWWBsKOIslK7NH6Sv4RU+O0vTHPVcNbhkFLITtITD0xrLa2Ucm3tyQl/jHgnpv8wIEwBWoid30
O1KYl5a5DhWF0MxXf2bhlsown2akxzVUoi5EgjjO6MXoFD0677c3vYB0I3+UNnvu9G7dSoCB0386
ajUlOflJtZwMry0LW0UQPVTQFQwFhbSIrP/xXTJxUuoAqJ012QaZ1VHPCsyCDuQx/1mic7uJxkkU
a9de+h35+5+89h1RoZBMso9D4bu4l3wNAl6S13DvfQiIdV1c3B5xVixOWBFDWn2Ia9WR1tTzgZga
3NGxbHI981VijNB77yTXH23501iMFY9rnkbnvO9D6kbxwb+3dKRl8PfxmuI/fPzYJ7OVNGgEQ/mE
J5VL76Z2VIVsU0WvFv0/Fqij/m3x+BC6sSldVvEicUFYFlpXM0o6w9+SZ6gPu3yqddfsybhNUbUS
XP0ig5LUB8jPHVQQiXmG+uJYMa3I8fJ1HZCKBZ2swl/lI4HUYjbCcjhYNntPLwr5nOdBArZRW/xQ
2AoWr21l9q9TeicieeK5sM5yec14LgP6c3bwDxUHMpM/++9C2Z1lGdKX/+PqSiHrpE8Dc7+ltopE
9HiKqQ6vSQ9SZWd2Qh793UohF7rSWKzNrZVfl1hRs4QUc/TLF3q6qPDXfnDPvGZx9g7YfpqLcf6E
+UGipbCHgKCsAYGCCQEdVCXA0X1gLAD+U5BE8a3Px+npyzrn87LXoqUwAGX/6eO1Ws/H2gDL2Rdo
nWRHhHVPShhXRjh5S5n6vj318QKvvxAxiz7xB562L0yNnmyT0RKVToa7vvKf2PR1vJ9McfLKJsfi
/Cz7FHY65hDrHnBMZyW/Z5g5hkJKlWNd3QnaCKKVr0//KGa24HSXtB9JrNZaqcRSXOaB+vRtopkb
N6SQNpur2pAwWeN+SvqEaiqxqRbO8oInX+VvU03NDBs6YSJ0HLlBswis41wXH0l4Ofm4JAlPY9Zh
bxyvFtB8mTlRkquegTv/MLkc6Ge5+UV2HAd2jzVBUqU6yjmlP+FInhoF3/yaLT6XbaC+nRxa0Lzt
aB3mWu/SjFtYBl3DRetybh1BMrm2T1USyK3/Gf6vcEFx5NgfHiGl8RSpRCHpzRJgLuxWh3hIomVx
pPEoibJlJ+iMNGCeCFVMxvB+ZokKkYrdeCBizF+pO66O0/2ra7sjsibYk0r0kh1LBLJDFT+7fFVa
RSDxtgphdoKXZBOPmbu54LOO7IZbNaVBZJka+beK+mesMF+IbYM6HPtj591/enb5GmdXktBtyorZ
mEz3qU0q5NXD1j/Jsd+zjyeYWLabgLqWpvQCnGreSPxnjryH+rh6tq4OBPg65Z6CjYRNdViKuKMe
pLXAwsv7aIc9JLdI/jBbPKJ6dfYnNB0oxQ7XgOTh9h/YtBjKfxOgDfN8v7/iX9h25DCXduufD+hC
45zymfm6YxqjBMNKGL8U+RnHq1uchRn1S5Bw2eODDCKFZIE1TOTLo5jVzxErKByxnXetD1u0NCt/
lnviAPjZXlbwgPkeeFlJLqPGJyCENKLrVXpwlUvcm33ULKnOV91tJV68jlLMKh6DDbSniRsf8ro3
BMZx/Rt46S4P+Tq7TOZelCizkJQ0ezPISta9NK7uyh10yHi9nqoSjVWKaTc1JAM90KoLc7gn22Vm
iBzPBObByWq3D4fStQH4k8AeWrIaz7Yo9Dnv4yKJju2ZOLIx+zok0AiGzQZ+Qotdkph9lUKrAByy
HmhCuVnAd55mVImyDRPnLz4Dbu0RuErPI8KWM6Cxe7ssl9TitcrWgiRZmnKTG+xQWFziKzfNlFtI
CdFOpMywMVlYSzDJmnStPg4WRmzlaej++L6Y+nfOndwHBkbPUMrH3TzHO0GCBwDoVoXfrYshAJ9U
IQMxkVENOu+VaxY6aESOOcgAGTz+eaV47ZfRoI72GRGyoIyDGmQude2XGditcbVkFEj9g1AmttAA
OeAhXoooQbZngIx+V+PCbntr51j8TPn5hbO0PZM8GJyr2SeOI/bJsUKdpXzP3AbGMIAGTpTNyMdZ
Cib2ZzJhu/W835I6F527riyKjv1lv6TyZ48zAWN8y5DhY6SDxk31jeLiQ5DPwEtJntOxtptisbZ1
faJVk9WH3Z3cTKnvIwYTX0R6Fr/IxcAAFgR957vuRvZBnbUNNgLFk/Qfi8nd2fx1285hZjS2Lvd8
JiPr1lFmt3thn/GtNAYOImtJ5O3UJySk56C+5jOFhKtvCoCpdyE2hgrVRG9gVL2yiR8vh4LQiYLo
Dv228k8qEqXHkzVHUk3Wd9/ViFBE4RoCMRQo8t9hX+rv+winkhyKVmQOayM1DNnQz+U0JYwhCnRm
ndoAaEXc9MVZ5KuSUAsvbOrgTK6lkyf6uI6EkTgivLztMvAqWbHviLuZJjuh6RdjxveJoa6bBO+G
wKdzTUI6RVpW98wx8shK2+GCBbXL3JuThC2SHS08hB9HQV2jlrlWHgxEM2U1+SAHH15xH/9FQsJL
CS7djmn6w+/frDFYE5hjVsQqsi4CXneXwKk5/Z6d6wtp4Y65rt8oK4UxZBNw/WLXCFBi7smH+3G0
gtTiVc/OblnblkPXNL1Vq9fSwMrwnQzweMB5mlT1klm3bxUII0yf9gDmIRqeDri77P2Vf3RFDpkG
c24JDckP+ky3iUwrJMHTylYdr+ithQtRQeG4u3WVrscty4gQGiiVOCk8Vya6Qkt7+65wsdp9frKz
LHyPx75K0fwZSyNyUeEy2t95YgFb+bVwTYZbsqEhXCxrUqBbf4wttx+lb9XKDvnwn0FTUKYd2XR6
4UJD7asfwWRBi2nPEhHHTtd2De15iepD+GvPlg7N1TZex/Vqg3o2xtkFhy61nzjlhZ8DLrOBkGd2
AFLQPp3V33EMO/D7LpNi1Nle+wkmjiGZZd3ai4k/pQfDfMKSry2qUidrpzu+qn9OPhYe2GXBBxCa
JZ2KGWNMhuDDZXvZEq1XkjihlXkSwAxnUBfVmfgvWNt2ryO5Bf8yHZ+tUzzOAWI+eQHdJDzkoVcH
NjbwquMh5UMeOhvmTaD5HdW0k7T/n0ewjtqthSC6blzqCMdFpXu3v/MKa46/C6Bws+5zHqwCOYuE
Mo+TSjF27lvRJPfuENlhuFBGR7nFa4yLo1RjZkgqkT77UVPeHdp976e5aGczAh9W9LSW8FtRzAYs
yup0Rf1MpCnsK6qpz/KRdksDgpZ4kDr7EorcGKEkWLIfYb1rQ+Gm0dF9E7ypBSOPe7PE2ROKKbkc
Q8IDZCs93pNfNQn1t82nC3JoYP6GUmYdsbh1jKz29nSI2koGvFKmq23aSIb3CsodLL6qe6MFZxhJ
q2cBw7RwCA8ApMXaaKPCsNN7hmdnow+rHCOE4tbh0q+G71CGbjO66QdDBIbuRKXOM5PBIHTHgGP+
LlFCGsFkxE1eFgRTpd/2KwYge9w4difa3coQn37QYvy610A1/53HjkBPmoMuScmZJw0mgi5wmosb
W8MUBEjiwbDEAMkGfqC6rtziMUYHVqRhqNesXaeDSuJ0ra4YWCl9e2E1bShGvWmUM9DTjpXMbR+6
q6iTqLxKwoBK05XYVsnBHpx2Qm0IVEZfyYo4ssriYbfaZrCftYsCQWGKlUkChJY3ITkGHlmnw511
+rnrBnG9R5sm9MycmNbpe8bpHw+glDSfl1zgn+ae4YygwIka4XgxYx0UHbDqmaixhcBCsrURnpGf
hA+xRs64zt48EwHmk9ggrRU3V9jaR+h35itSNTpPaAY7dMqalbswybCPHEp56SAUe90ytG8VX52I
DZUiXav027Ix0zofjLdwR737/1cbvEXPMfMjHPZbvA/ihDgy10Dh3QY5/GCXpSALkw4swShcr4wh
kP7BOc7Jb5FRw60w7xKc42sU/WNjxAJ+WiUnul3X9xlJnR52D6rPW7eMLo2FZIPUgWEucjc5g4YE
7rLj4dKqcAxwRQJlmBEarFDmLF9XjgW8a+CScBqNdCRikHmrKiVRxa8gw+wuWugrYH1sRHttCaIa
w0gco9wgdOAMN3sBgRU7TF27lc7ofOlYPn68p8YiEIlaLnKsRpvHIMrT0Lgj/V2SqID20CJ3r8JS
kuftvQ2mem+d6dP15J478jH/DfZfrzHf1dYhQfqKT+TYp41QR3BFtmw04rz+byISv02JkDR0dpJC
2MIcYMyjyuozVS8GtW4XkI70Ez+WwItSawQH4Esde+/PQOnwRIFP/9hXAJZW5Q7PHiDZqrCpEOP0
hyvkx6KljpAxM9MkvhyM3Igd6OJrZy35CKI62iu/wv++gaYBa5gUxE0Fz3qAOK36JiSkSoXiUHDq
MbyqRg6eCHk9Jfnd7E57LWBjie2P/8qg3j3Xbltju2A9jVELIq9/5/EEiq04YlwFWkzzykM8mYSq
PZuKbTL5emfKHT05nacYQbvOCQl2S1Q5qt1Y133XV38uV7aKkfL2+NDbdJ85oDVoaQN1tWyHaAPH
k8IBhAwr5EQcmJzgEc3zIPSRJasHm5Bmr1dkKZfDXSxCEj3VP0tpDC8eXWlhX6S7o6BJqzqJSn/W
Yl19rpup6OJlZoSEiKa6KkOTNCPCgFUK6/UDOYj8T8P4vrh94TPSoJkwmpS47heSep1MnZn2XKch
2YH16D3zc1aMdAbSAA1+rJNYEW0BpmztttzeIPVk57q3z9SFt0EqUPazTAWYN/ZOrhREPHAC3yBx
NCZ2PvOrHNRMX0Fa0+9nkilFtcCUJVuKmgu5rM6BiGTR2wFlKSR+PgpSAMTjL9fYnEgUX5SVmJm4
kIPlV+jQRx7UjCH06i1NVwxKAeNX72H0D2JjUqTKHlUogcki+c/l4MWnPRLWEYDengteLUNxQvWt
R4ZMVI91MxUAbnhZSM60i9gX77wBeYrda8J1pxM1Vxx15ib30oig7Ws4x3DJNTAQEQy4lnj4D+sd
++VjLFZ/DgHNEyCNnyEAtiM/5MyTdGe83xs1LOnfgPmcHlD8OJ2u13I+4XhQvH2ajgmwXesOVs/l
97iJmqbGxMJ98Edjv1fN4ruUFBZQaUhOZA/wbdWTeO8H0nk06tzdeOKnqCYirEnvlWTfmgrLWJIz
brDVDSfaMKuQGG1Xbav0eZCrxUun53zRsa4toz77pto1h4WQy/nORa6SQLl/TGtqR7ywreWdoCwP
dAB0UiZ0SvZl2j7Gcc6kBc+Qj/oOIn7Lh6A9RRgJBD0lgAO67QSQr2ZzqscdAD6kkFperEg2O50j
VcVXtCJfMZ4e40QjNJadl56eUHptBkzfBCH3FjXt1ZFkoTs/24ueCoAaMWTW0Bn8qkRJqG04raCY
wnhixNedxW4jatLNrJHmFshTD5PNkzMNaGoHGys/7qwsUHRGxAucXGFUpix0pcWYQisNG5eHcIjw
4/JY3gfBVkTUTCKe9mM4jpoly5kCIOkAl0Kvz/vu9KLNigzfp8Yf21/+aBLUTrG35sU0X31U+zjT
nTH7VnCFCKNv9Sjc984auSIxbwrFzPRIte4e0Ewog8+GHf6UnlQ4HZginsSl4BSsaNe0BsjnL6hk
+eVSQrVniNK/sD0YA79tcBHyBgow58SDkfE0fwC7Bz+oVr8jxzkYXIrh4sUC7BSuZq3mxBmYXvoa
npZg08LcB/M+li+a2y7l/svcpZlfe4GOsjOEt284VlRNGbQIRsjeYU6gQ/ZTKe8MnF3nGcVuRNNb
w4+IQV4lu0jk+suc/Zmimn+IPvUc9+zPJy2hmJjhuLJ9+XSFnmeFSptnEhWe7HZCb2FNxIvNtrfP
NAF75/kETK5aTLCLqjczJmzHJ4VLmE9yxxWAr4MwtLRC7wLDYlUk1B4ubH5cIfYd8BvPKjgUwEnp
Ubu79C3OqjiMdBdgAfJClODQ1TCpjBrRIeBIsSMCYbjLoVybJm45Slb2uxexkHJFJhIBjIH22nZ4
ih4jTLtj41XimlqafTSY/OBstXWxmOn86y6QD9tu8PqSrVGe3zikfpVH99F5eUhxi3yyVPukCBKV
zfUht+CJJZMgJTJQuqWqn8/WNJbPA4Q1Tz2xb3gjLn2nOyUp1oUFGQT+yzinvMmBIk6jJ5PqyWAS
Od7JpiXK4t7wUH0kdARMkjVFuzx4zKsAP9xKcxxZldHKg1on9ryhQ/8ph3WIaXM5umSGeSXucjw9
sw9DibnJqJGOa6WRkWdS8Rg9l2f3xndP/eEkWATdObEXMgR+jtE4GTQegLO0u1ZVQQzHemgs717y
kPqdZJ9HnCWoEDQzIO4zIoPrV+i/fu0VWNBPUWIXJAscUelocHnVBCRkkC6mAIBaTYiu5W8sNFF6
r40Dlwako1tlQRDFv42nGOoAdEKc90ntwDMN0TXzUDpLEdI2Wxgv8suTIsHM85mkM/uwaMzjt3M/
XkSdMXtLubd8UQO6QP3FF6OcwBYsJ1SaHZlhtRqsNFdeIypunUh4efgluiErB8sG3dZEj6eCec2/
K+oEwrD7nX6Fb0Mv8pdUtJ5XaSMJ2wWC5UbDOfAxSRH2JPrf+A5NPgMh4Qp6mZjT3+mQ9WqgLwqo
Lc2bZ0rga2N2i4OgeQtMVEnwi2P/TTBdNUFuJ5Fk17oLkCFNlutUzw8kl8VHJwaAzqP/O/78O9PG
Zyy7nV6wTWT96QuQoy2FFeSEXli2UU2ZasFrOe2DbdzNPHUhQQ8M5yUENMQ/NHdUBbCrVlC65hkC
WvjWsAUYEQWCAXhaNFzYXtjY1aHpzrQp9EANErdVoyhrsHxS13ydI6fTFJqJMRN9/Cr6WPNrKcDc
gQ5tGeQxNvD6o+XF0PR03VChbbNicTP1sLLBSo8fuAKZ5lV71mv2xlmHtyDFjm6X59Yzz2jX8t1W
UDAqTlHN/g+9j1ReZiituGgPc45E51MCIRJw91NLbkfI/9h9No4nTwtdkdiBV3T+jtelUQjY9Jv6
8Setnl4crTgAoxZMm+0y9iq82lDgxku6FzBz1EqqUJDNYk4ug2IVrTpIusfGmdhn1ejhncgT2g10
dDMShRUdMrNJjToSvH0e2ApvsHzjT+VOpzEg+Xm3NJUybWJy0eTWOPdlydAnNE7VWTz+H/c50Wwp
EpkvvQMITd5S1YxG5LXUTZxtg54SWh4SimSndS22jcsOpM3BBgMct3eC9e0BASETmBjmEb9DDyUB
bA7ITYFLpU5+OUyO9rM7OeD0PMkLeu6eviYqSD9eBgwUwKtnuym8W50mLKh9+01C1e+S00vzVOnd
bCzOFNNgZFz1bQzAwpOA5qZ29LCinU1MZ9/LSKqs2lYXH++D+FZu7Y8CGVYkjZGv/U1IDCWHsM9T
gbFF/1R/UYkieI4L80Ib3vJ1zkcYKHXVlPLAwq9zBErG5bvePPk+RM1loFIppfQkLzvbsKOEqmAU
2w6TVnHMAQCvHb2YRKDR+Ty29jmEURbmN74D6LaOUUDYtYrGNI56GetxXd6c6lvPpgOjFGKouT1w
sJ17rJRJaD2GiW2t04Q5m45bfz+coQCcU7ylnwVWeCGuI8q1oH3N0wC/67k/J/UrGGWluD0aIjzQ
ghOtia1znyuWEYxAJKzmmr9y2HY8JNG4K5f1m3BY46naq+XbanPx7moUYDkGYWMffg7rxuiiw9kX
vwaGMYnoVYMbv1VhLMjTYA2cQu9FpUKN0oPQKtCo67+6LsY96V47ysiAUQfcOsAKBwtAHNLt8xK1
wi1f/OenkVijo23Cn0d4pL1rCHY7qF7n5qrVcUH7vbhgnlyVmMQKmWG3MNuAm0WBkfC2ZTwjGCBA
I9s5MQoOBle2z76fqCaTrQZDlEbzIz+/F+ZZdHsOoovjXjqgio4iq5y2C/ggG0jnRPn2xscU3vrY
/6M2DTbOOV6nLqixZPAKiZtKMnCxtrwp1NZ5VoppVvN5AH6S9zBqezKuUNUCFg/6EKvkSPW50r6b
pIXmHPO6kJrMIlqmiq5mYPozyO58Tsyfo9J7ZKXsuNuWRYKCa4RUU6Vgj2SEoqj8xL93oj8G8tHo
S1vC0jgOE/ZJjNrdNceAfSWO322xB2YkE23dU2AUuLM9TgZ76uSpUXopQcTwe6LSIxze+1yX1+Xi
zW0zGR4wleEe5ABoDfMTTV8MpUr85HDmdOQuLhN71JFNIgJGo1J1oDhTJkjyHJ+BTfOhlYLJ8MzL
y3KUEO3qAUOM7eqXES+Dq/Hu/elasGAEyOlomEk9dI4koo2exmvnIvxpIFTR3dQAhV+2PoTSzNMQ
HwIly5S6nJ4lbKOTYN1L0jCo4c7oEzi0QcFZ2xSsTQyQzDyt7O5+5KEPgLrALBpWJ+meZym5R/Ay
+rTN1Fv+DHo6FXSsSGev/TxTrZN7vVPQLc/09QnFD2kqOpFH3ba6T3jY/nj9tUfRpaauqlYYTviF
x7i4whPliiOJfF6bsMbUMd9pb9A47QZCSPyeJGVdc054It0/N6XgXQQYYciKItVhr19LQVAwnm/+
nB1gS3js93uhbQJSLSV7v3A6WVXGpgPWM+txaZjDEfim2KbyHcVoXvmUIF8/tVc3hCy/yqMB/aHC
G78p5KC3z61xS8QyWOV7+cR9kes1z+BI4zuSWIDr4NZFbZ/yE0rkClzQeJGo0OLkORdSaMF6dHt9
UsrueJf+epCI1XShfgQBfPqrYRL4gGMstcHTYFURgcKZrbZ+s5055Zmsz6gDrOrjEv2+5zJYUTg0
iLiyAHG7nXTJi22LdkTqnIoOWZXd7R3h9RVXuJ3Itzn2eYXWXb8suM2axljzMkWF7oROQBPib3NJ
rSG4Hj89V/vM3WFkHitmVC9BdGlHfOx1J0WGRBF2JclHnKXWKv+HY1VuEvwyXDb64q/ewpgNjSpW
YexAXcyhPuQ0uy2erxNYsELp6iKmNILNtLL6q5A3aBi60LsUW/neLvh5xRekdvFs1iEnAyk1z2lj
QrjBOWUjfNOsi8okFkfScKmItoG5gYkO6QnbIFaJvf0ZXgYqb+zIrHizp2sGVcQt9JkSfYbcAk/D
8ePKl+Mx8hrxxPyYXqqtnyDGKIhUD1+zYudpa+tRtoHZMovQHM5SGpdkzCxK+C0TxSMdItM1YKGb
WKd7lr9rZjmgsg4GgnsgQECnx+NqUojXkS96Pi9Cy1AF+k6OvB+XKF4TfcGBrDMyQkcbFdh4RVGB
FyCAZKsNtMzZgg4LUvRHe2dStPYSQR49CFQXcDaDhixFRVavtAxT4poMH9l9yMFhY7/y84bzzH8u
tpn6NzTbnq8dI7KG0Wr4t1J/Cd53IyYK4QExV8lnnCu20UrCI7sO3wPTJ+CdTB2uJnYKhTQZHtOf
DrySWQfbU8H9Nufw1mFfjzLO94DmUMbgj9XLUExWMsPaLw8PmM6MJnd41risYDjtAxkdKYkbpkj2
g72Pa4XSsTnHVIe1GQI3sWcUOe5VztnkhWBNx15wealer9gJk8ajdoBNLJC4HtyNOVxdvLuNo7+p
F0p/gAta4S/luW16S7oOU2OVqVOkPKMYQjRLpxygMt8tyewc6LqaTX5+RpmUEk8MoFW4/K+02+w3
oZbW+YjH+RLqaIDJ+UGT/c2e2cyZ67uRGWYG4ifHUpgwHpwTl0rkBAtRktj6vzINKBW8XoccUdDU
Sz+Hup75h4Z0qyvuCs0f39zFpW1Nltdu9JmzCq5A8GA4KMCElPlB59x7taij2NNVwIiQ4x23h7Fd
E8KiQVzpV/viPg3QnZO4VAgx8ds9lCnO4mkmYjEfMPSMwwh1//FoyMc76knzqF0oHy0yO9JmL1A6
nOwTEsG4RtEYX4TB5iPeFrBjIxJDKKO2jLXCNeaTCRiqsy73HAU68jfLzE93Ix4nuYSyFBnH/GQQ
/Wh2OqlIKclw/ElkqXLiHPWM/jm51+8C8WLt+PwPbbysNm7ptVnMx/CGE0zzCFxck0Tve94Bn45n
bHZvePNZt/vOrekpO46pOKFMx3U4hRO8kDhmRkuOhsojMAXToR7SNjLdBRDSaVpLekC3YVhVmyFr
eeSbSFc34APy62Yg3W6XLmpxWJ2yDnzySA/jOMcO1rL+O6CXRWOTo5Xe0x0a3guIxwj5UBN4GYhT
EUByYq8DvmN3hyschqWXCJjbHo9LO+9V/uB/lQv6CPG5wPT32KvqrSJo31jRDDUxL5lMktPTOak9
q4L/cb9SteVvwCGxmA3B4tuMSNoCd5xzKWmJa5PNygJRpxbHkO0Egd4nbYh86hat7sRfRZYyob+e
ih+SXw0aNCQon+KduLWdi5No9OMWoT72Whr6NSZ3KrGKZPmKGbqAK/nPkOrH2fQj+UMgrxvYg8LY
KuVKBb+3O4NjkSZDj2yOid9BYcZRmVdvHhcyCUuuVVaOHQlJ2xZNfSjqT3qO5hiJZobq12gvgrY6
ldY2aiBwltFN6nqx/sVxO2H6UynXHYSfG4JI38tm7HnrjjWxpXLKT2pEJg9VEnDRoCw1eKLPokXI
GSwEmHoEW/AAgBmNrh0MxxQbsMV3x4IMimmTfz8RoU5wwg+pOUaTkqcIIDBblCK5kvwZ1p2goimI
wmvck4SniOnrk43N0NQHhKJ0VVvgM7bjWx1mW3rJnBynt87ME6iS10BCMH+edrnwa8RlGzef3nRX
OTPOI7LUKK7Dr07pU5pb3TqrcLTos+Oz8/dODHMZE70rHP/h0MzZ4btxbkYQhOOB9zHwAWyyZw7/
jMlibEjf7+ApTT5LR2ILL+OJxOZE9CCpgRKWuW6+WWX5yX9jsuO6y5hYfi3Qit2S8nPGE3tG+1LA
5ERBeIa0Zdio4lV4cOfswhGNsrfDpinm9Pyu2IWF2w5GMB8E/f+1SXV9unGylZiOi0VJS2ac1BDl
lv3LrppS61wl3jXExNuaJA1qO5vH+duwepXMvz8WKY3EbOfkOvARrhAvw2RrTXMfGnOY4YK+gM6E
CiZE3oDmys/h3tVJoRQZhqUln252G5yactk+F+grfXuvE2r53qHy1hDslLXrIEyqlUVIrmd2ckV+
Dvdj+kX21E3k78fIimrQDqRyoKiUbcyxQYNuNlZi6HDwFPCtCncfgkxkJWkujmzfz5e14Du81Sjf
4S0VzR5hUtk+YwJhohveGAxRcB0j9SJTmlOt55OuVmtjCsfPVno7r3Ca3D0Ivuhl/Y5FrgRwiWBy
HoIyysy5YaNaCfMEDM8dbw2ojFzfIUHLDghf3Q/iFld6wuvEbXdy8l9UhZ5f0YlOp9Gv5QEy1Z2H
egrd6/T+RUWLlUPgmuzm1lXuKI1zGBwEAEe7ewjAqhjnYko89lvbdPfENWzKsbQ9c/9px68hr1TE
ViV/u6leVXuumXBYKZD9XqZAqfKzwv7SdUIiQMf3mAr90iOzWRmWnU2qFSor33arftt+Llowaey/
gLHiBWLkmgSAtOJJLwy54akZrnh2Fz/QwkSOtXNhdYR9C4ThJ31jJ5Mzrk4nAWi82U6LC9wu5PbM
9Xg1dYCZfy9+pTJsBVlsLxTKjrUoVTrxBPKgjmncg++7pxrTN4T4YMygdepesXLTyPWe2PptSBtY
Tf727wtLdii0q5NuAt67+Opq00oSsByn48wrFrTAM7yttbS9/ObdvF462nzdaFTqMnNgAGXlcJo/
EMCPQs0TRcYlMfH6/ji1Ii/XBZJYOVqlJ0vSbfKOjnwvH0Q0skuqSiQW5lCr4vigShOlfAVSB469
EqSjOixTxPe9sZL9QUE+LpD18NOwMSgRXo0kjrEpfr25xTPFMJwjboA1mD/eVD/nFQUzKJhDddJE
4tXmqreW9vFFCdeTv1mRg7d6KBMbLZ2ncHZwHCsrgqwb35fqMkcLYnb8RDBYqBh+MFJrNKT5Nr4z
apQdPm5ey8XwwP6IDzs4v4zdA6NL322iUB39ggEg92CVd5RBP6WmidYhS8S1LweHjvnA2xRmhNjM
0FVsaoCUqBagN4aym3iIiE6WB0Q3aLHovLQW2uv9hibH6RFRmcq2okDJ0DgC+Ljfs8+Q65yoBSxp
WyLd/bOFA9+0MefQhc6FyaSZNErZsUo/iHsQEYvLQzoC2v5LylqzSCOd6EPdmVKBtGJj5s/f5Iaa
6CVm16+7y76xLVH1HF8F7aGTmrbcnkl+UFBWDAvBQnu0uFMLh4M4IkB6Wdq5N8fMDBcjFmZZ0sfj
KHLNrziPzizXJ6oju/ntR7eHo6hL1hzQsUBFjDB5u8iTPGeySfiQ2QPFThFOBF0nqy2xy6hEZm+J
cySBtVbm1WwfcP8KSbb8VhyyKPOv1PwtQ3n+AxmIspNkOMNLUha0HpmHuJcN8yJDbMLlFoR/Qlnv
u1pcZ0ON9uDTkrELxo+tajQdABzDDUn8LRmeMY74I6y25E9+7HTN1qqaJqYDzC+VeU3svIXXwvbR
Zy/QkbAtD2/r0gT9hJLJ3vV1bnxeVIXpVbrhfu6b5Tg6deLCB/SbOdXguLzXLtxbhF7YdbDi6Zyp
2udzNEj4hhjYWKqrobVIy2+7+YWnLgXZwFD0Oc9WKM8LxAeAcCgH1rU7VYpWFY784Wf96AHUYovV
uBPXPjmkIu0S1P1Uuv+mkrWE0fSzKYBoKJIo0iSoii6/ZhoUv9icrR4pqpxxZsZptWLJMvZekuaO
UNzfsaYQK1XOrMfZyM7MsjdO8GSn0K48tMpSm+5palRkJEPrvcKbXPutWVhY98Bro1RK8cJ4R4Tm
lLxLCSz+muXZFIJQ/GIBVhB7XL08k5OVr2qHQa0xY+EXRTPJzoVZxvkj/rdtwnQxflSqw/gYmXUH
Jg9HwLkR5gheMED12M5cYBB2DEAikGDRzt80hGE/B+4mb9M5WgDJZ1F1wtj/rFvueyszspTB7G0G
sRdMJIwtkBu3OImO28weYi4FVlDRcOlZiSITucxdrW7xYZWVRdyNiOiODNUjNh48V9SIVuSJP+sR
8FQ70nh+Gprf3/L3aKW5F3vYgxtBMxlSDfFpJpPm9imLkYEizAPTM/ZTSAXRV5QJS6uGVXWHAYbe
F3ZcsVQE8gS/omd2/D9FvgmOHrlW+7Tv1RniRlcoxHnxt66yTxVY76yutY5xPR+yatlHLV+zKsp1
zC5RMVknhpPxkZ1LMiNZnLEE7UKyODQl1Bj6ljjhuj+Ytlgm/wjSpKo6k4e1+qjSQg0s8rwGeOqD
k16fkR8b2ZdMYyGStL6WzxMm56ZcjczixO4AVt0kHgBV0adWgegOM4khAwVax+/FTA/MjsKYkFbF
3YkoBE1vd1+WWOJuQSmzT8D8xIPgHnhhHXY6yWsPvg53UYhpGpZyZUAcSTC8Z9C2FRRGh04SpKos
ylaqElMDzJVzlnBJutu9Job2G0z9m3Zyoqy99uQWo6Cb6ZMsKmO3lFUypVwblNsg9m8WFeDLTsqk
Ejlpz5CDSlmgl81MeJ9CDulrvZqFyCy3/wy+wzUTr7LW+tUafnPPNHyDpx0tdb1s1mm3hQncDWDU
aovPrv3g9TvkqFjpbhOFbnCOlCo+PD0U2lpZrvwgUq96sC6LFaMMZwm+nij2z/sNFRPMAlLLfU4Y
JzuxpbbdI3iQTXDZO59gl+pri9zfyavHIW7RalJNX9CQO6s1LsxmjvKZX5CuR1wJNDEdnC8HC71p
GhBJnSmPkIY99ZEsWsu2OalR5FWFULEh/kQoZQcXgNc5rv9O8rM24lEqCHmEGyoU+qOEB/Q6Cdle
Ouv2hRTFXeFz4m4U+kcHHBObPIl0wkImJDTi8ZYDxC7oOoD4J5I3DFYJmlftmU8v6iiO2llnaD4k
pl2wsjUCE501y1d2AwAZpMwWm/SSeIzDFiXb0l+cgJpiniMYykQk9/8Cz+8NWMX4BUkhIk6efvmw
heQVC6Cq90tY+5dATcpMWHkQoqoiEb4UUHvqzZBgmPguYqzjKNwHmasgpQnOXVL3CuIT7tuV8Grx
3b7LiGrZKuE3JoW8sswDjf5w34fKK+kipD0PsQQkS5ppwVEDf/WSHNKiqOyfacUWgEjRypGeC/t+
UqwR7oeJkz04R96VomBrlTIgMhovI+vaMCrHYUl2E2FLZgG/HOxRh61+VT/MV9PcylRqdSZvuPd8
dkVDtf8IwISoB07W9adfq4eiq1LYLuaYpb31J2bO+YLe6I3RhjeUhQ9J/nrP+MNq2u3fm+dlSWyY
316USR9h4MpaFrISFV8oae3ZlSAQIIn+nbNyHaBcIIupq+S2oKD5cyG5i8T2mt5PS7b2GskZ/gaa
Zmgjr+p93nItoe6k2mzbISnoOK2xynuNOXvPH1f2x74hKWFR9OmPUB7BT4s4RbjP6AgWlJgv9cvN
vCgS/iWGDK2188J0kQ89Fo7HeA9oqLh4OWIQ0PnWKaM2UmN5cjNq8Ms+i12rRTZd3puhGTcRftWi
FyxQ2BFQjjN2cG0OMmnBrMX5a1PQ3ClbLLX3UPJTlk8f5AyaM29j0xKs04S7YbJG+I49K7eac+VH
6IXgMbhilxX9tqGAGLL9koRDr96ry+azWNMo36zNZiUMe4X9F4zW7Y4AZbweLfZVVvhVejRWD/Jl
sNKYlVQJJv0/K1ZKK1IFRMQC9SKVT4h5RmtAEpAVaT9A5Lrww0bW9Jz5lr6DSH4kRSnaEQ6mI+IY
BCR9Gmr9JMn3yLELxMazL9qJ48r1cMR3U/vD5yRhfR+Pt8GM9vA4ggmjCug81SeqsooK5ePDGJCT
tHVPb3cMbr8nu80O0akzO5vsEUk9Lzz7hQVobwpKMVsorc/YRllRtKgYynxLcHDF69RQV1d/Uo7H
1GHw3R//xZYiU9tp52qF57cybGMz5V1Vg4I43nnC1wgJJEs57N+EUzIbF9qNpVgURhqymTn3/O+j
hIx40IvjeokSoTJTtkbvVDZHXXe2B5mz6sRmqF1Bm5a7yOziwg35CtHEsuif5jqqbtIDunvXa6tX
WvAsPCY/eECAWYZor9aG9zIZVxShf4yhoNnBKtFRvR4sm2mz0WGvkKL9aK8skpIEwTGzMbFNivmE
J6bcp01nanUS2a3z3w2kXWRRLu516F1VvX206OLgIDBCT0wQCKHE/0szjPJQDFoga679iKIlgKKY
G3hLQ+b+52vFR4sN02xngF6ELYn9XaGKGAcXil+qNLwd6uOuEvabY3s7b84KoM0ztW1TWWJrmjvo
O6JOYM1TrY2zyeqdktFhGyNhXfVCxSrt0jyOOQ5AEXKL3HFD5u6yA75Sb5PPOHpNY46uGgNmTpkv
dreeroYjq5rFt24kKZcykWT+Y11DDu/Djapv/h8t6L83EcNSDa0o92HtUr+y53jGHOWEps5Rb/1a
L0b0rrH+djs7gBJS2Xv4I4Gw0adjWrXOMaIMHq9xzQ+DGUA58TqyUtE7QeovTG8mdOZ1fKogRt0N
JfiQdJAqltrpbEreUbGgZqRErzkmU1ejPwQBVhai4A0uFH/5xV3TDX+FVxKXInjO91bNMszmjPbI
r+vBaY324UB1ny437I+0dNrkelhR/rJqF4aihAgxmIzTYQ2f2FateHtPx5l0bJ2PDf8Vxu01vD9/
OntLF8ZGO3gvS8w65hAajcVtpNEpcTpRN3n2ZfMyluJin6il1corrRpCKQpL0/Ar3cqWGLDFvSo/
+pKYo5BCcZ1LnlF/PMAnR2e9xDP+FHdbWz5vdVq8LKe5g/qs+eE76XZ9RGHGyhvlHOzwX3FOMICZ
OPZLv6aRQo+mEdpJcm09gW1H06vi36xeZt0ZmhufvYu7wcuwohN7CtEmVDGXaKfv8ZCtf9HXi3by
2ohWTNJVCiZyTEen3FZ1gEWvlSsJD9REJnZca/uYi6a5eIV6HeyhkPrBlCV2csVCdOt6MZ0u3Ljt
2N+KjrkYsL18/09GSmX4hImwn/piPXeDbWwIKqOvI3JZibyC6PJ8gnb4atRu+ck0L22CIgYoHsOn
g7VHFAiYvbG2ydY8evs4kEiT+rBTPgkEy0npNBbCb/oZubuRoSH7XAq16sgNaIq7DoDF8XIAnixv
u3RoJKaQESRlKvKTCY3lKB6MytbGyWXa8fmHhtPdZarvGNdSqCDBh231yzdNd9WFXM1/pL7HRZ1/
At7m20BTVlwcsIb7WNEQZ108Wg5h2J4An5iB+aE2SEXBYHQpa4TMqJO80sj4WFfW/w2T3DvmUC2V
LKimdswn/U6FbhctWjBmPEzT46LjTCBhbkL+Hn2/gJRDFQ3FuEV70g8N9a3DfdVpb5nheJetmF8i
uQiPwS+iakOE+R/rqvYl+2NqZlzKTYXa6eurA5n8fLqkFuXeiY7GNNG/f1zLhKRH4Y8c7eExH+rz
l1b+NkC7gKlt50d7YlxGWWEDN5wb9O4NpKxfQWYCfaqkm0rq+GX2QsB4/03eQ0jZmeaC3MvUq/df
iCenVQeBR+xZFAoFLKbr7s0+4Q4T8QENtKeHSSlk+sLzmsS9cu1G7hftFox9yBO29OiNtYi9RRZm
DlvLq5b4vNA83ZlVqJv1mvwW+Z6QvN6gZpwzb52alNBq8rtXx9cmY3/edBd0ZzFiq5337LJi6Igm
oAzkw9jE1lMGmNY/rT74WaerXFMh4FkqvwpEH0oXsfDGdv+SIrI8aJbl2o2q4Ae6bBlj/GeT1Lox
+O90BboSSffJLloGNqN/4cTtVLO62ahx6nwphEzk+LopYTjew2HF+ovnroCAJ4+eqBRDLvoBUPgB
vU2q87Db4DHgORd++5JMorAtfZapTK4Fk+L+6/oYTzNejwDO0l8Xkn0fLMS4VkLtPFhy1kUBAdLL
WYem7CCUWD4dsOLQZE8BP0vO/6XnRkn17/IINVKQSXvZPI5A9HzuLI8PckhE6/UhsNIrcB3OlUpj
3uW/naAZezB/KIpSNG9j+pfenH/8G3qgfYH/Y0WJAV1ZVs8QFYAm1sHBVjmVEoA0Xvle1QeH+aEi
/CifmHZgrSfu2vccUEse6yvgF/YDAXXeTdgxJDjRXgSu6h5t8e19nIIZl/0UOXopFawgiostIDtX
hrJnUJMel8yAghdwm/XHWa855KTNKJRlCBtqM4bPtMm2GH4XY9d6Bb09u7hjvUy+aSWWDVqorOmm
9iYZnJERr8Ruouc09790zOKPNyWFilyx6SNwIeiNiUkuyVIZTtb4HZTda3njTLsvIgwghTLDkcPF
bgp3Lfi11+StfSqGTp7hO9wJ7GCiQE2WW7sIzO0My41m0sXzjCr9ZCMH17NPqBajwJj8zP+P/iw1
4VqI28DuugQkzP0WzC2hDRYm7Etko5DPWq/yrAj20YK//uMhdpzx1IVhFWkTOJYvgMwA26BBd5wH
ykF9BfgFuJgbVQZ0L+FhU0cZwnA+KBHPwAObdVBDUfjcMQpgNwGXbZOtfJp9kUvlGJnjqLK2LrPU
+bXF3YeUV7fyvlP0SwqtRt4c3AnL9GY1d7VNFLfWxllngIK8KodrRsPPgF2rcyiPWsRNgPrTRcmy
G+vyqiDdj5blWnzwaFA8iWY8tYsWZPruN91ZDnmLEi5O748sn+tK2L6SDYx95eW4GiDeJt/2PmUq
pOYlDqqNVCWBBE+1yf3v+mLWBXxIW63QlgLu/jCEXfuTxdKrpWjI1EL2MTdHh4Ykur+XZ5Wn7Z0u
2kUFTT5WMqa4eZK7cKyaiNTZCQ8YdN+ZciSw6ctDM806lgbiB/r8z0TT8r+FZVEfbPo4MU0I687+
flt03NEkNXD9PPtvs3zLFV12dbEcvksEGDwjQtCGil3J5KN9SlSFPNrDmcVVkPfSsf3MlGvR1lXT
cdUj9BB3SrWJCE7T18yLmapnfP2V+Wb2vuyVsDTTx9baqEBCqgnjExJl4ubO+i0oc0Fy/LYlu/Q4
mCL4+KE0RmQriBzEZ67u44D0mRceI2K11A2OYiElBdIQiKprhmJ8zALvDnE8x7Bl1n8kC6Z/BANi
jLN1a9XE6NUgg23H18IcTN3F6FY3MCHtmGYBOl1eJlaj+FUdEB6IyFjIGKSSeYtcV75+UI2G9TYt
xYjOqsht8R5xiEvH5uz8PdP81aBfs7WenB+HC+BRqgpwRKge48I2mDZkUBHXHnIS3XafxP/568Ak
kZrfwPdMRuZMKTWnu7UH68NSu8743ngleXMwV1zqmMZFUsvucfmoshK8fpIpBq9VSTZ7l0PxWfN6
wcP1NRPpRLj/tTInJCSR2DJK8RK3DkN3RhTk5NxutAuyz1Xe1vCQnTC04JAQF5lFS00YhqBO3zay
A0Ep+EAGajQvGf2jmPaixw2dsQTWA2nvaW09XcdB0EQy1v36OViBCDul83GuA/HoZYz0jwfR53Tl
8ocefVnjaac5AheTN+5pWk9Z7ZmtyVYd17tI+jR13xgKbohje4DcVssxUiroMoOYsO6I8/ZpzdQp
pUSock1+ukkWl9kG+rT6YdjtJvWjvEj8bfStUsFWubkqlu+UlOuE0LI23zKvKuH2ifZ+2/ebi6nb
cauToD7qjrsDUL2wTUeDON49ZjGdeuoYxxFOkG2DixtC80rDal9ZOFj/jYL6065bmmtjbyyaPgeO
w6BX8MxMGJcMIf3ZjxjsMwAAyaBduzi1JmB1NydSMs7utrYqdN8GDF18qhaSZNt+15CBYHqc5H77
MqMtTBRc/M48UguiMnSNr7LDA8SM79BTWVFUUK+7IjsMyU8YBfaYuC8tW9k945A5ZUQFhrtIk+wq
AmuDnpAPY5KhyEUdBqffOSAoRmD/30MCkRwNnV7X2LKsqNEv3eLDBbU3O4n2ML1R7DPDI5wFooxn
64xD5th8zTqm+/TO9e/QW9VgkJGAYLvyVT14U18i9+Ap5pJsr2nID9BxICKMcYIv8NhBHZzNK7+x
arlPHQlyZ9IETPp66/VTxJz9VRFt7b2WKKQD7EbMfy/Mn9/D8KeZo05T+b/WxCsw0Pru47Om0PtE
HfnwKcjfFxW81WQLBI7tmCcYdnxW6fkl3z53DzZTsJCNd2/kiforLf852KpR1n5sRW/cUxiTaI1J
tPy2ID8jsEB/1ULKdhAboQ5W7/YFTmIqFUiUWgwz1qy/abK/0EwJeffEqMTaalFB4VtHKemzD8/F
lriKiZGqjWuL0nQ7ZqEq/lqax0tjvk1XgE04QlhR7LoFiQeHSqkGDToftoBcpiqQkwZU8BjFuUIA
rgLA8Jy0kuULu51/WtgeGCz9AcON4M+c7lzCEWghot22Nqg9404UYe6RWkWLj2mk1dZruxJcrzJN
d7kdbbmaL1Mo8lXQwnlwBj7JchH0w/xoCBX/bLmVrNJ5oApi03Uo6JHvSW7iwjp2veHhepJqXNJI
wfrQkoE1gZSGG0+owiDWAbtFnq1F4XWoQHokFOlbJ9rVzqJFNcfHUeAzr2FRw6l65D1JHFRgdzz/
q1gNnTjedG/VenGtKGgI8ysFJYe0Puzece7hOwyaooCxSN/1elsDd5rXC/ns+6GnqcKHXc0faNql
zD2BJVfzXBhSatiqmfp+/B6xQRXk2yU+/kOoDfHkyjmdhuirXrn0huaBFtg5iUcKQDka91OgGDjj
slLuFXH8mUlPvi5hnVx7Q2O95iEfNXSGiFHAngIRWZH8L2JTbWrd/Egcb/S9dfFnBO2cKXGKbNdf
5TcEbNiyp3nIt22GANY8KlNX7zjVcb1+EcniZDL8SB7A+iSS3DYbss9nceAaCh5o9ZZXrZXxnKcS
amklAJz31MURdKW0ldgSnApzZg8XwsRK+r0XHbhlV2BfNr4m33OJoa8ymGigYnOLHZQTAyza5qjn
ebhlgf9aW+K8wD8jO1bSuSOGJwtsFU4b2HdNNkPDrmstBZg0FWPpx+gd5LevHuOgPj0/yoR/ORlL
14BXTpMQ0QfVOwLCM28b1Pfil1OBttqlzvdWedFMe/u5K3jhG/Xmx1rlPCx7YwyOwzbQYv+Q5BMI
WvyEoF8/HreU2QB30Ly1ldkWSJ622b8bwQxc4vSKiMh5wB9PNKdztr/2NkCOjqiC8KFrU4Ane9Gu
69B3725JwCzguvDzTBgvZEc5JA9/zuZqDHVcDZmwO0VWMuIIDQhrvgKciRywbLf62cpXWGDJNB9j
PTs0aMgPjq/f2bdeyqHhKkFj5qlBChtCxGQSMGQIja+f41OhbxaQUy9TjCvXYNE1/bCSFa0FWYKG
7SfH7t1CWLnduagxS1/Czn7bUzU2oMfmFoiFhqVtaYPwNAd2rKb61NBESSU/pp/+OC6zi61Rr33i
fMaIZqcHYA4YgrLERl4MA8U8cclgOaFUBqtekaHW09ORHnhqjphcSlFtR2aF6h0KQtA5UCOTAX13
1+6vr1a9/ogyrwIOuht6rKmksiImXnlxrmPRhzjbOzTG1+/Z2rpK9Zbz1OWRqrJ4lr1VXGEd3i2m
1BaHBDcc38bb27YBhGeF6bn8VjXn+zUlDBSB4VfQ/+1OksOrQSTVQS6OF2aH/UofFxO3D58bLrfs
/3WaneD/XqQCHWTsktTiO/778chccHWB0mexyE9P7IqN6yfYkckge6SOq//RFXBQZoBAjuu8jOOa
fpne9NFqPdTjLl5WwBDvHLl+K7AfXYpwOw/LvSfuG0AWORYSR/CDyphDen35prpyfNO8KRxIHiEL
ESuzHO5FSUOE6EkWkGVmWa2R32KZ3UzS8xORj/8EuNwW8Cic93onCMOhRYXK6W38gCAst0j2gcd2
RvuuVVp/7HPhH+iouTopDSEZYSjMirLmFMjrinOBx0MhhFHi/1u5eF3Wu1fdADe2nwNpmROQcWcx
yk3i0KD8j/o84Lddoe4w9V4yHDZHnOk4gLtvsVpD2CTLD/OCa/mZnTm7cpSxaQEHQM0HLbom9jai
xWACsQketjuybX3bnaayrRdw8D6KvnK6GlLK16uUf47wj+cgQgRM/RSvmpTcGDCjch8qLojJ7MBX
9V/QaSE1+xmYW5ypspBgI0p+VfyJ0Sr3y1nAQkVK+KFG13FkpXYG6D3gigm1dFxN1bo5plJOA/4J
krWffOfjM5DrPYFyVFqkkyGgniVVqGuuDteQFUigWPjK88nC5V+97+u8OUX5Q3hXBFOJpccdewls
nrNLMe87YzcM6FojVv4AgPXu1us7YP2GnMdRrcQ5vYT+VQTKGfeNb2W6Y9x57yuUv6UBHgA1v1YU
vrUbLTxWCeiQRcRq8tIJxK3upqank7skqOuCOIVDho2mOKWQHMHv7v3dITYu8DPh/8EpqlTfN6zs
gI6WM9hS6z3xWOSGjPv14EKzyX2Zj/k1kcfNih3etiB3yp4C+eUe5GF7Wt0/cOtfl5HcMOqtT7eo
1J4KjSFiHB57qoJS4ea2GypQCm3uDrPkOtmF8E3Jkyl2xpfmMd4kTp07BbwRTJjDBMFYd+h2i+91
zQ95NovljYYheElMiv31RBS4jttaXNYg7dPy4IgyT1XnWLkDbjFGtkVTcCSnOn7gWraCT83dbPAn
NUoptX75/PTWI5lywDGUNZe0CpIaL/GBTV6vXVVPEm3JmRVL/IGOFK8KBMppYrHp9R3VccX+AMhN
kTn+Ze5II6JC/MZVGqWZsTm5pJMLIUvBEQqQOob19y51Lvo037QSjLIGc3LXMtMzn8gpu5xf2BMG
tGViLNa0SxVk7aUnmle3QdnI8O/sku/XzgGYIaslpDG6aPXj8vie/5lZ2jV7o7sf9EQtwNr26gWe
NXX8053nsnllMf3FJkcm3GX5vO6DsEBM2TgimJyZvCMJqC/OahDpzuKHxk0OTYABYFKZWoS7yvMz
MrkLnX5r6Sp6RhqyvWkl2BpSUP6z25EQ6PgxILv6GaZ13D/iHQoIGlJ5btCNyn/4eRCHdQGsWLas
WNGL/nUzkkqrHyP395wxy4m7YAg1pHERY85JgHA8Ho04U17irPGBpWzEJBLHLUUmms0QaEVwiVTz
erOF0ATwFRvOsejScZyX0g7G6razKcrWdt+DDobk6SuisQdX56f0ik0XSNzs0TeyfDPepcdf61cX
33gjfFnnevmv5Wh8CMAfOp9pTD9NVnIHbL/x5P8wKWAZZuJNXLb/boWi6pbIZ82BKAZDxJq8pBGz
88WbNYs7fv8JAtrWPTj7+S5SFKwBaef5uGxB1gR2jxwFH2tSkAF0sX3Qy4O6dTApcRx9DEuyXyIm
SMKFb3VIHcyyt4KzGyAc0AwWwda+QUODgGHt68FVM4DfP4eMEComFNG2xyqkac48SMkWPvhOixJm
161JyBv88W60eDzx3lS7hAQaOW2392qU2DROFT5TVJ07EvSX+hkkDXzn6T9Qlz7CUn+jT5f/njxH
s6u8Egggr9Me210RJoaWHMLIc0ZdHtf8YQahUTvSza5DF2qNopfaUi0MJmTwK+Dpwq2DmszA6taY
653bymSBr0c6X9auIE+Fj9EyY7DyU3lpo3uqWlsGXkrew/mSQM/nIO1yMhEM4iMAdBwP/TWgPpTN
HwnUd3zH3sfZTG//2Jum0TzsAbs9dcEi7I3vihB8G2O8lF0YO6OYPbCexACzH0Crybf++o2LiGZ+
FmLlB9Faeve7tT8SsL+P+0o/cgcgnHkHKvANvBpLwL3C7TsC87W/9wSYo8ha15POD1fbLsFwSVOQ
FMNOIoYAVtkBAhMJ3lJEw8MGQV8Frlo5HohJ1U77iB5zV0qmzQk4PsIbvEAEbGQ4YWIGhqm8rgHb
14Yl3NeLXhR+0NUG4b33r+aPoC8pYbMgH6NMXU/zwlyFWRi0BuKxqOQn40Gf5+sA/QLgxnVaEKrf
tpQyW/NfNOeJlbqs92MASDEgOySIQcqGvT0hEAXaLEagZKfWkf3HLToP0i0s4NQBqfyPX3zgrenn
8IV68KfwCnxdkE5xA5W0zskcnFhnOwDf7b5m++r3mrtM6kLupKdjQpxwl7cmBMJWbEyiNEPs4WxA
3sNaY+WjuJfFVR219I7nRRPZiXLULimLPUfuLvUaIKkDBVMZUKq3juSs08CPSTKcXC+JUmGexGUW
4CZWWoS3vQy5RvJTAhzNx9/2SDNKgAgMaCXGNjTJ+ckfGGz/UgOdNRbn3Dx2X3awyQXF3dc/nPVt
01KFFx1gEMYCDd19K53rGmvfTpL7RSaX1gO09NnoL8MK6w5gTykGu71DOUGUN7JzLAV05W41yAK/
KwTDLQlHmk9634N9VTmE6EW4jpcEoxi7LuIF86cSCxl/Hm1jN7G2xFA81b1OI38EfTRgxf/VUYXG
tABCtQQXqwJ8mi+PVx//6swtv4G6aft7I+sA6AZ2qB06ycmNgXrDcT1Sg0loby247JzyOO7SLg9j
QRWe9LbavlVHVbfejh6FTBIIxngdNYAwLirGY1aR7SDVHpqIH/cCxJ+3y0vzdZOCMGwRyJUaS74z
aE/gOQgDJJJj/n65W5msSdWIGfaenLhdhy99R1XEarAUes10GIzn8h+3fy5qIK//ZhLJylrwIqD3
sGjvfUGplQsOdO7fhrLwp2S1XT4fCpKDghkPkVdhKXP+/hT/zYN09/Msp6X67H8tWprEij3jgGjH
3jMxwBarXS4PYpxIdjtGOsxKYcjhlfA9DCK1OkVxuIvuetOwmqeZYUYIjnjrymcnI7n/mj6UuC6w
xQghlL35K9nPHPZccqnJc9EMDhy686AiFTOHw7TUO9ge686uhXhM9gake7EqaoNTIm8VvwWq/AAu
vwHQy/AfIrc8aorFcWZZ1XptIwh1cf/2j8kzvYe6RQgr52NsjP6qUGgzJcvaqUpnGPww6cmMeksY
lWO/S/2hSn9yv1hoyQlP3Xt/83EItGK4Z/vQT5dnDzRFBogfp8qDYS15LlbBl7ww7kCqjrxyJlKb
Q8KWaJTywBCkbV6d5yZpI4s7PI8HZmS1YQ7f8E4V7kEt5SpW6w1XtCmgvpHQyHbHE/+qTIraHMUw
DXKqJlL0kjNfa1WQ2J+3ZyRCWw4dCdaxPK/uaG3tW0rTiXJMQNbsBamw0JmOz+mYXnDtTkdFgKCg
ISPpp/2lnXJNG043tkYRbpgqXn20YZHTUfiCnp82SZ/ws6ExunSTBhMFuPhCBTyNbVM5EsLhVNE9
0MgOdZDWcSlUyRhg4uFeaDYpBMMDKy9/aQ+L7Eg783yABPJcjKHkOe0GJYELVkONCFI9xFrRGcc9
eDkrN65osMYIjBU0XCM7t9YhzjPV6FVzlSINsd1bRIs4LzBKADh1ttF4lA0Jp2puCmFa9P/OT5uW
TC9DYSly8kvY6pz4LMsLmb4o7vdNp9ECy4Itk9J6NNWn4mFJSCsqcazk8ds62JoKwPLA/ti+8Si2
EjxS3Owi+tEjVvYEkAavQZUj4J4/FQMt59Xwg4z5TooPKL2yZeLngxRsa+X+yjPqoBL9LiXBzlzQ
4FthIewD1ZEn1754OpIlQzzdV55iDpNIny3AwY7hcJo5+q5p2waEomMXAMN4BGSi3qrc1C2t1WXg
uu9J6JIxA6pnjHSwlPBA7FO/TShl/fknbPGgzF/zVV6dQnvZDTGtvjKQnlwfW3KFf4jFwGMC1sWM
lHztEhQOu8nRAKD8NYQh5Dvg6/q3cyc6Nv1mS/tnfpMVPVLDgGJZXsHfX+kOunCG7JrjVP8B9ek5
uEIiW+WoE5S6JITod2Fj/c95D4b9+Xx/3AZf0wO4RuZTvq9OT7n8lDqwv2GPInmTe+tiZSiHTc1t
LMSzEa92DrGkwG+yjDgN24YMvGsbism3jHKlAY3V76kq6vSJdMy3Jh/y3BmSupIm49xQ3mQW1xns
WIY759CiETS4ynwYimL+gZ7pXGi3uFIMfkwd6UiBRwe4aUlsIW9j970aEbquh4otDiNhyDY95KyA
85OZkYzu0N/ESPooRzFxMknIrCPz3WxN6d+wL7QXl6Bst2udqpKA1ACwJ4JwQhDdypArkhWW6Iza
Sh2WBBxKcm1JZ1EaN4C2x2+rqY3aZMqbXdDiMkdetwUpVTxngS1HuQrquoOO94wHo3wH/GI9Aro2
zDkKV+FKZ9ojsuF123oBHvmBqnDbQ0ASB8NxE0EAJfyau1amsyq9Kj5KyOFz3LEzTE4nJawksxTQ
mphhhvfJAhtJEpAJSNAKE08mUuxC6Vi5qbgyfKHeBi/W5Mab7Uk0R6pTHrGiOTo4pX/qjMsckRSR
8wTuA+ck88Ui9Yg2gzQX5UbQWNcrRH8rXrWtybnl9Qq6Z4fhuCkmdFLoYmAD/ul5U3rraT0MkX6h
/Ra51zGoLIlkcHP/b2BmgVh9hKM1fhjzRW1OM/9kVnGzK5YM1oQ5p2Kuv8ueQ2v1ZH8l8WadCZIe
EfHOQnG1oa2e+/Oob+0RNFFjBzKQVm8DaZfuNyGeZj99n8xk8N/oaL4UwFk+fvdb2uowHcYLDp7T
NLiijo+JjQ1+OPed2ra7R7xLs0Z9LYBiRw0qQD+8CDDxRy7pqi+Q0E8TmBatAcEFG2HzjsFqOOek
iimwdm1lWwYwR0LkGt4Sbt0A94bllJLIleEkWcQJNPp58Apn7+Tm2/v5JtbclXPP5NVzHn4eHNrn
wg0DwwaoKtB/zOZ/FQJMc29KWpItoxYoJUQQvdWlweCZi/45JHX0W/bV+Z68vm9n0EF69QpYCSyx
GDqC6TR2LwVaJbuXIPsvW7aSrINtp1EMx37gSXU0vhrhYJwRIrWt8wVp55GVVP31SYrgWSdiMkZv
PwifO1GZzL4gnbGsOW6WxhPT1Q6kztEoeWooEds8Bqkk/LAfFsTn06l9EtHV6EC5H1q1I7UAqGrf
oLRKxZCj9B03jLi/gZC4KY13aaEj6hzgkp3ruu8CxCi4clCVJDtj/q/ENcwbCU/DJf7k4/7i3IoB
Q7a7baN1i2rvUxnQ7ZOq37suG/KHQukTPc0KhaPVg6CPWNS6kur9VmLephn2K8ttDbW0dQVYo/2m
n+8FwR/t+DjlQWhvy28C3pZ9T3hevIZPaHdMmuGZXSFGhx60j4bYUK0zN5hupkrRh07rnoMHSb6G
JvWX4CWrfSzbw0HDTKO7LXy1TjwEoyF6g3W7XUOe4sCLGnV7yBZLrqVHckRXzboVDdN0mREUwkrm
PmQGT/DJU3tcnl5+bLDlTlPnlpjlQWuXKCz2wwzAF43t/m55eLVTCyNdGTfIdPho2A96Q0qoYeHC
nDENBcFLcG856GBSVG0z1ZwQr54uGTwpwVXEp+Y6PehF/cyB50ism/gV97mDrMoUByBgFdLd7qxs
0QQ5fccODZBOX12SBjJZ97IyMbVPknmbxVAhphP8/TZy+DtuInkRuaNrlQBXK4aZGP9yo7krcIdG
wFutsMOjAr3m3Dq/cOMtTkARr2BgwpdZPIdIr46gC8asWcXQbMV+ooliurY62g2ZdLgFrz4bFguI
6TF8MPWzoyKF+bbb+oAj5/CDcBNv+vIFyrlgveq5g82dbmOx72QvOxgPdRKKmnKT/jkdUF1rm3Q9
Zj0mwX9+qc7SaZNBegNw8uIlF9jn0sdCSxBLenOrNefM+L7h7HmVGMLuqafCGEKvTTv4P7BiSTLB
oHRBegRTnMOMlLo1pfjsYXS1iUhRcIdDEJpLsq6tmjFTYfyk4KfRn9Ci3KzmcrpmniV3UVEF/u6Z
9OZm2bxip+pOS1D4VGFVBgxZm2+SGlSsXX5IOrikkYCKOGxrC7LobuSrk/IxP8ww6ri0QdhytWJr
/Tso4/fH5vLgv0pnXO5q9aSlsvLqIC79spyGZqpxp+oNPVT0q066aLa4hquiFuZLQh4NVhttGzco
/Dkw7bCt1PxTs5w+HI9XAmvTGYxUzDk0jtEHhSlE36rXz3ZkWh+pwTP8C0DGcSmqKLmmk2C03ogD
4s6emjZxfaSPmgOttqN5DRUifh5o/lseRYZAyI13ip/TTdiNW05g/l+z70bO+ThJL+BhIi7AdXrV
spBpt2kJHg25VGikrNPBDKcx+SPX5TKlBFYd4Ev8qJ6UBmX8YI3avVjBFBe8WVoGMA17X1uHj06z
bLWl/by8W03MU1Ra29A3cig5lQRIBZTOdVu7rKceAK9QFqAnx5DzPlnBdWgrbXznJwnwHwG0SZml
s+iQ/H1AWbbDs673V3LqaiETMvsoMF44R3KikXVp+X2EDmVzH/UXEoYVByjTLmd5rkQjBVEAStBV
7n0IYk6rMkPnY6AVUalpJA3NYKCETBf+TE8X3eewxbTxo++JYEDPZF6jqkDGl/hz0n1KDGAV+Jw8
dCOfszh35fuzkDdLRZMFjDk20oA+rc8m1ldWcKKGuj2P6ebiLRQv7epsz4fdwYvZ5K6AoSLSk/xO
IJnmERH72kgd45lKU3fOEp0NhSpXR8p/oIBrEqFC5rEkypAOwbobQa7s4G4KSeNPsex+hS5R29bf
P07QQeHGd+YMs+3IubOvoyYFwOUa0wQ5g6QzfueaiHDSaGyxG9xvkaPkG3Ennb5F3df0BcKVSeQy
F8KyCEFVRkyiN6h01NJEfIljLUOOdUkitTO3FwdZwMbbKSl9PD4Hu54NDXEN4IEVYMI2deNHqZ33
DD7lIkcKPbyLi3QVuLl5l55y0lvsfgNFoUwgaAnXts4rbsBkGrIMDR4Nhn0vdPMeuphG36bC2/jh
VfVp3SZV9WTKQavJU0b9tTnLaDBWA2TQonZ3dErYJpXZgRUS5pkEoTPyPIzy2PpZqlD5huZpBzJe
sxnqOLcE9FQzjoy8ljq1/u0qOhLFCfh71E/mnrWcB2mNxLaLkkcJ4On+cAcRynJpEZDXJ6CNLk9q
r8CeG8cR288XgMQr4RcxbR34Zf0HZVfDdZlCRmDAfAfP73xbbZYCWMuyztdYVVJS/asC6b1aHhL8
HQ8D2QDNI6r30zOprMpAi1vaGyx5vjNzttR1bSFtCWUuW95nK13bjfVgsg0NfylapmU4gulDX0Vm
Zwl2ihn797pja3OSHP6K4EzvATOylDihJgLx8Lak5Ev6U3559lL3ndlrygxGA9qpUqWIjRwgWRfl
vP/21vd7p6/w55/OQdgSBQXqbOsMbWT6fsFLBlOF1/eg2/0JlE/lKtiMJh8aoWlnVGc411GdxVrv
SaF6J2zlX5GKbDhUrmJNVNtLcNGQMUjBxrWCnYjw3y8dSlRNw22wKnYEeqJORVcy//IFDvwizwQt
HCgQ/0TSTl/1fE5b/R9X9/qkzCy5AWdNLxMQ/Gct8IXvpzzlCIKkqcHpO4B+O0ZMGuz5rHZc9Puo
tymDrlStu4Fbp/un70as8qyz/aXuheoIXZcyRzSV+9HpyKIQ9lrYvzIOlSDqpEVj59cljUx8aEeS
lBjxRMEZxFWbbRDpwy5AXJUPtklnabr78ndJM0QIxGgGRAhlTkZlKgkgvm6sg59f5pFU/6VPio56
EFlYcCRLdxeBPaYmUeM6J2Cz396E28BIrg/Ttz/nDY2xiNmPtrvMWAVfmOlg0V+8phOsDgaxoGxC
0xTcsHCm1ldjcUe3HcH79b3WmwvEv+ZuUhyUR12pFu+tvk4/EeA0vDZY7znkyM2n9GZCO6rHrBs+
91npwbkHAcGCx4nnmt+q6iLCGeha+RnhwA2j2zT8tlwqH+jrtUp+1+QKGBiSrFfTSma6qSSuoUyL
pvC8f/h2qbsITfqvw2+0uprxBlIF7jbgUmFH6E8iBM9Mty11GIMFwFH6X4mnboPLifuQuL1B/6WW
LgReEgAzdwNsJn1mpMezYwbWfhgs9C3FoEMyrFAkt1CGsRuXdh7PNu14huOJOjxaRapHfVHdFRrc
S5/PEzPBvMUq4iPEIJyCWoYhUc7PLclkvxtq7Ibpof02KLpEiAw/53UrdmcqwuoEoibYTR0aXnj9
ykxhUuQZU1TroMw1Yj2PEhtwENX1sP42D4cGRD1f/AIvfpfi1toq7AhFrMrYHq9KoA3li9uCYXQ6
zE2+SvR90Hth1+t1YyTaH1JvFHMkQrrmSMGZ9oHGlzlDCC21291Iw2QkRO1e2lzp/pXODTVzgTc9
3oAmw23TrgWAxNcHnsYXl/3fSNsFdg6Hx0eGlKeKku91L/tnVhrm+8bl7QilGueworWbXw8ovtgA
76nmOLHHtkBe82GN8Y4WiOoSphnLbqM4IiapWEH5rusSiyni6LbHjpouRkUvkcITLJw4d9HVsJ12
qqdPHx9Fk9sfG9M97yLiADzRMaZjzA7NH6Zeyjna6qZrM4hSAoAh11oHc2osZYKw+TojxdAqekh7
as4iRr903A/hOd611gqFTsBACehw2FHybL1275DrqF+ozYCgGi6br1OQ5issdC1qPXFUBgnC3Eug
Q3a8eQZ2Fj5jHbXWiGPuMNVN5+y1rtKcoh0QFXWGCkOVCh/9RjrWR91tYJUm7EbPmT0SGePFYSqD
qR+PvhbR3I/nUBL69NPFyyhb+oTbM7jxoQG5fUN3i4bO/hgdhimiVd212Tay/6W3jcbd/8WKBE/n
R1exauD1aKPFIoIc/KBQ8B3uBslG1XL7U4yVM6WKNrLJiGqeB8BxkvKv2Stf5IvTxZEtzZDcXwWX
ksWOKs0FE8MXLIofBguFFOg8VGKzknr3RI3xdWDI937o2lFFCW4jJWr3mBmRxkQCz/MI3ftAIRg2
dCVrQqPf+/QPwktzlMWE/ofgysHVCb9qa7sqHuU8GprU6NKO06eaF9yY5iBMG4OzbnaNsvMtkwLz
4iZtpmNAOhQHVEBIzfNQN6mIaF0wh0UhKcbr32OuhUDqSMCaWnYCX3GTjIOZXpeqX4iJwniUCopi
B5upuJjpkQ1u+0rTRY1YTgYXHqLTWLR6RCcUeM+sprSiNuTXB/LWSnwb+Xm9xGtmWqJ8NZjCD8Jd
7WIw7duGaSDyos/nD0xmt1tRUl8947b5KzKIb+xpvCV0M3VpV8nFjr70rEKjVkO54S0IPdIL8DME
gPMnMO5hZXCiYyIEM5fYRu6rBjYavAX+UyfXd3QGhDYnEIVjO1Ls0XRAAr1LB8u32hh3WLWLFCie
PJOREU9zbJIDT/ZwgHfKc9itdxYtNcR0DDqfUfZjIWXpFdB5PtGvOPxxFldpGqmlXGS2UpMLUBHN
SZxG1BLdI30N0dfxj9ns48G9MqA/+l4oilz99HYLMjK9UpAcXPXzTL52RrLtqd/Z2Fuur/nhQjd7
968dc4nA1ZNqX0bkHQdGjr+3po0TmbXGIZIJ6tqZwwPGU5hr2gSQGqSNX5bd/c3OKjJQyAVxofPK
t9FJU8IFIbspbfFTpNvqZRivEF/I28XbT3V55+NN6ZnmdxrvuEjyzjNyaTyGQt8mFU1Ja71ZEEIO
Ce0ZV0pjeylzz9mHt9CfD0wjw6gS3KTvF3pKcKUB/RHEcy6zwoCxsxPtrVmig9KrwLk1q/8kFFKw
u9NMzSg0flgSZTil2b8wszlFxQFYRHer6hE88u81W+IzhB1D2Arpk2XYG9TbOuChTskyaBvirW2s
1/OmDwWRl5JLPb4rZLMTCnujzN5VpnMC0U8EgI2fBxKmeOFhA1SDPdwGLtGRlD1MJIgcKAcDFJaD
ehLU34adzTemeQV3X95eakgH8K0xB2g9LQbqbMsn5ddzXKRiH3CQ2vEQT9UOp+iIwPkReMynfIRw
y03VeWiKMl4SQJ4rlXTEo1S7oUPh9fE6QNcWGAjujhPhvRvkJw1ADf3UfOjDq587BZXTAwmcB2JG
FhJi2wqeewGF3MUKztYIGEYOJ2bSx7q0GRZhEBsqIqFjRSE0nTlQ+8cQnmYl2tPKlNhJ09oT1n4b
4ohJWuA2wNXf4R7G/4MgX3VyL1BrN537W6g8j3fijk0pHceoMl4MqfdMyqp0sPthjt2Mbijf089I
0RaGee/9PIymQTqw2msKJs1vt2hNPoVYHoJh77IC1ZAJWIVqXr4JBdBi41gS9JfjjxduqgIKaVNu
EeNv6Rcp2iPU8JS8oS9x8QMuVrRBcUVEZEOR5y0o7IRGLQP2NNO8iga3vtk2gup4KcYBFA90dlkj
6CXwT23QIn0ChAqAC3YWnSe4giPIxh7XKb8Pr6TiMkKvzTKfycpQzoRLaOL5J8gFf3EMCYN4SAF9
OEv6kRp89yCsAmprYVd9Dr+mizx6V5CDHkqlmOINmMo09Uww1be3cSvkR1Pitlq7mbZpiDHj82N0
/q3ECS1Kce5Xt6TLqg0SwusdLTM51B1CD4NWlO1CijVIO+9/OBnyUMX3gyVO4pA0WaR8XqXJc2MU
5Bl7O8BQwUqTfcrLR90lu6bzai+7vdo40O5ljp4grVxHuiLwn9mqi7SqEP5kSo5Rr0A2679IBNnE
+InA2TzFd+ZTTOO7H7kEF5gc9XukhtJrJmKAEcXReFGX18jR0ymSAR7W/5vrJeMIge8rrZSKPMA4
rNrPHEDE2xqF8VA5BXGUqgjhpKayL1uyUlaBwyWPIhiyiwx5B15L4ivxVv+esQskpDA4u/ILwP2f
HxOfT1mna4pQDyP3wAeRtBPvMnpypkHEC7YRRntZmf2ySH4KYVIcCEqXzb70IaOyv9NV7Ajol69L
xCnrI2UqN5ao9FbHv/sD24GCNbfPKkBht7iFdOn6dJUnlijbNGjjjh43OxmBbkUpnYRqNRgUK6uy
rzLfNXeadf1F072tmJ2PEd6/qRD1hDCjKokJqtlOcuXY+d8YcJZsuFo+KrDpCRNih35Dsot6Ps36
Zxrw5ka8vevUjnyPPVU0Ah9OtIqscyWOct1U6odn/kygkpRfJtE972hYl9HjCRrccj5Ixp/k9hxP
SBCDeOXxTwUaY2+ZSsKv0HsHuqYdEpJNDQrRMpFDRHz5XXKpdr5nO6Rp5Oi3p7KsrKk86jKtVEZP
YrU9RqMaUjl0Eju+blxHfkxCO4QDPGOGvBjM4ZzljQILsUksJV7KNDgBLkTuRfnqDssrLaRwJe9o
VQkI9DlMzySgrOOhMYl9TTawkuVJ/3mLEOnj+UEIe2TWKJYpULVuDS1/8J9qhYO/fiFFhnaeEksY
C4tVtyhmtJGdt5EB026H+paLKiQDyq/Aentmk4dh9OBCC55pnOOBqm5KgldMJ06BPOlqwb4HIqPf
dGIi8xkBwVF2JSITJOBdocOy99jt+mJNn6+oh7x+WIRMXgk9rb3bZCk0Y5GSKCmGtbxzxkHuCI13
WiPxLvZMljU3I2X2v7IWJlb6vRK7LKaUaNsq/yuOIG8Rn6JRPvBXD8WvUUF3rn+iuFiy/fRpoACX
AAjZ66gaA9gv701I9OKzkSYx3tmLmId0pHSA0kUlfHpI/Qx3sBQO1T6wQQ8QXDDPfm+xj9HwGLrw
RKojDKeg0sFB3UXA8KYxvYag0FsEJ5D/vtOUEdjtPVuhmMWF5cHoP8d4KDZySdV01G1lvyMTp6Am
B4ruJA2IWPax7PaiWBRa58sigCz56pQ4K2dS1DEKsuMABL9TCWD6HROdWWhuVehBi28vWv8LkrHQ
bP9LXces2uQAO3pHkS2W0tKXjrjIT6FQSWKFHQ3Bq8ipdfgss4qxdGPJDLF41ftt5InrS7pX5z3E
LeZfzkrOG/7JgluE7d+LgdfDU4fsVkh78gymGrCnBDZDIxvnByWnPoKKlMzp+6eZizbraq8Z3Z2e
PXpAi3aNL3NdbmRXxBnR1TbTdJS9TWq3xpbUs9IQ2auht9ExhWCwb5X4jPfQaBxWnSbWr6Zmazrc
b/jQja7teR29irtj5rwAP9Ni8Lu0hoCtlLNT+so1KzEPEmQwxGMJrJNzDnk8tY5G1y5vOwvMv3IS
uG9C0ma9/vRRFYpL5wCUaqtrwm0qB22Lh7Mso+UlhpSbrcMclUwm8YeYfu1bzmseWN3HwGvc4V8i
hWHWZpyAFhPFhwFuVWx72vWlfA+56ImCI2Cskm95wjcvbR7xmacwsxxduHMmvE0D92NfKhMkQZZQ
w3X8c1qNhy6D5Ye+E95xkel6ywYlLsl/NlHvIRR4ApP89Qkze6PlyxxgNH3+Bg0hlUPktwQobDZ8
MzFsKNPyHA8H609QGSUVIwNkQyJGOuioGqSmkb9G/jGeG4L6anHrIlsGgMKrO+15Nw/8m1ZN/Epk
+668qod2Hh5eZ2+hafRBiJ16ZzcrlnfF/3aA5da/bdRuk+Y8cIEDTMzE5OoopnB7eBphiGrCxk3t
jZFc+6BvCBecHMNXUE6iFFyX7kJ85wmCk3v9QHT8k3pt53gYHdTrRWNZhoTpWPyic98bcadw1+KQ
y8eK+C0hhzgnpen/PlmCSh1yLhEUKfoHhb/Du+MJHI05s1wV7bg2SZfdE2jQZI7+9wW2amAjz0O9
RpEpSfHU8hhEfVtYsO4PWlPOOuU0sPb06lD6mB/Pc/DWCqY1RA1SI5S25I0w10ge/yr9vBN8Jcyq
a3lvqEn6YMbr/1+l/emWPZgGsiMv6fw9oOnZC1Zju/YLWs0nH5v3ddnMrqWnzllGiKw2AWYxF4Yh
DsHpO/w91hbzNctQNGr+X9CucdnGoswDtLWT9kRL8nXC83+1b4xLOYNV/kzM6ug5JanadCChp1Xv
9LTyeRH+lDSYfguPFZgl4rtF97ms53ViA1kFl4qQkeINyCfFsekbTBegZ6KvXza6t2M9Gcd0ebmh
lxgDQC4ZPzZXqFDnVksFEnq2a7Z1ZerPWUm6hXfRFu3a2yEdSjoszwQDGZoeO+ZTCmYKIDfbcpr3
tAuO7ZyKvJ/Yl2PZdCLbrXWTEz+s1XXu3KM58Vj1KG+zvbSnkd+te3EgQE0VZdMUBrLXWIuMxf4R
cBI7PKTtoIwDI+bO5pw0Ya+mG5l4FCSBYbMb6d9M7gRB5biJ7LSPci0cjWADg0peBZvNbj60cPoc
apVNH4FNtLnB9T1LG+qxej2uMe+1kXUD9fKwO7DyXPFt2ORqi7lRwqLeEZMJryvt9KvbVGd7UDAN
mANj5oX8JLnRuWkDjl80hGyJmjS4LDB9tbTWZoG8/hNgUoJE7kN+kvxf0T5UpkcPz8WJBTT0wkcz
Mp7nwL01Z+XyPnnsYw3aysl0UAbVTY1kpbqXetu1KXSdyRoRR5UQ3H7XAQwERS+uiwka07cQF61N
+qSOsnWsQsNmM/i3vlDt925I18UFo4z8GNwTsJdZQTT/GiMtf98VzOocgYT3vBm9NvBWIthO63xu
z49NT8/mG/CfCXAQE2WZWjGbtDGlQdDwTJAYGQVpd2WUtXHlqmeXhS1udxQMqnAGjgouat4RcsJr
0U2FK7tt6/+HYIFEq7a1Ietc48qUPTjQ6o12oN5VIIxXFOgATw1zVUukeYNDdPQ0RijFO0DdjOqr
hsFEOT6wrm98+O1yNEgzjPcx4GhJ6Gt+dejGpLipTIJ4qZThvYp7j2vQXPrXu2gWpUujJm92jwNC
HnNXVD4mrh1ReUMmEcIOp5Wbk1GSKBTxa3PBVHiz4JdVONSbXLxS0NepXpwbaUb5uV2jgtPL9HII
rPCgclcYirBo2J1IQUHC3aNl0YtgSyWe1Dso7mKRIlqn6wnDfkNF1Am7tFJWgOR4+THfGfyzsnU2
Ct+Bb9Df7oF+TAPmiLfvS9Ttoszw3CCL+RoTS/xJwC+DnsEI4tH0hpqmqb7/tib0OFR3Zx6o9+8O
/FjhQu0m9MltNG6jr14H0idBhVVl2KDIHlYcYac9yyjvV7ThI4GOHuQyvaDBqnWdCpcJd0myUskb
clL920SDuljPynqRo/t3d37nnyGbCyBNJJuy3irapIvRcK4DTHV8e6DiwsXOblcb3lEwUNvtphWQ
MBhHBE13yiv9WSL9VYJCwlW0ObiFml66zwEU/iH6UkgaH3CPeDMwRhmUfNq/XoG0G5AP7Gf9PNoX
XmkBxwjSw0Hmz2P33XX2pnZdAYt9/sikpieHAmMkkegCEztIoq9Sc3DjV9Q3IDdzCzRnYYMxRZNr
mmaAc4ojPemNX6B7/CBcK2czc5nISCmRdETXixxeswcSAeA3Wckxow0yzJuBekv5B84sTE/Gj9fe
xmDmI66xuIGaN/wEFMhRWV2QqyY1IT9j/yfgWeN+heT8fNJDz2fzpjBAm6Nh9TrlM6oQMjrSTFrq
z46hhRIEXy+iVolgpvF3uc9GhwS69YYkK5DnTWN+gANZ9ACyW5I4HhzbJExgR5CdVS6E9/OzRtBv
ZZSmHxKir+vUy7KN3qEGfryqFazNTw/g1BAOTL88KLLPxhdqWJvBFj2phS1wUu9Nqex0bbXL20EG
288wHw28JYzWxkUYasRazNB8hfYq0fiXzNGesjnlS+L3Scf4QeJ5MDsm8QoBi0ZPmbr3osJ8Q/zn
hGvGb1JzTgeu814CMgvZrTF/VtGQWYR7D173iSEpf89zhwi4Fs4sD+ddGVpnZMpSRAJbq9XDzJup
WEwW7hmBQZzGMWfDVFYPhliQ1ctJ7oBPU0z5lzoHJYxd08MAdpF5TzUd5pa5xcwBzD4hLPwwodp5
JyHld58fZiVOJ6Yx1cudlaBZrRzdqP6GMsnYEjRhfSAWhFQfBzr/yR1U9/zNwER3lPsCW9WZFYYf
W7dI89PjLTWPL8KEH0XhGMMG9Q66fRJK3j+9LR20nQW/QApcmfJssckkmxBUD0GB283mNuGKkh+x
lVrcBBEug4Wzm9JbgcQYf3gM0ZYPg8u2wx63unopIuuEGeRyjHideOYi1lKfj+8G3Fge9Jcwzi6E
2HPu4AxpmLcDmc9EqCoBu6YjnEn0fBzscXpeN51HegsGk7KGLp1Mxsx/zE/3LwCr5cg/3RKmJY42
G4IBPlFnQTk4mqaX2tIorh4yFzwJMw+ZqLKJHcwFubi5SkQQlEzA3CYnc15b86n3RD6OXmFU+DJE
yMibnkdt+EMcGrpycq7iObasTao0DtDhrWNCHVP+UvuAl4neR+TcCGS1Jxp0gycMROlpmMH+SeeF
t3j+/l3lJ5i0Uvz7ErJz2NfzkJhX/jXZjPPhD5PRkIc4L4rFNPpvXeqibp8VOm8lEO5dmrBvE3D2
xqH6kkrp1wU94rKUODrdeUPhk83+bO0S5QW0tZgU4RvmwK83qUQtfITXfOUbZE+mJw/BziXGfXNF
zYnC5VZfgERX3g81slvO8yZ1Bd7vmc/SXKTWBJqffgbcUmpp8thTm5CMHFP4D2uydCTZIRJeW2ZO
OjjN/M2jzhbUsQs/OKDjG9vSpVuEXQYfe1cDnrfqkinzAKliVGkpuktvPWOoxcIOw3Bp8rTTTDHs
qllWjG6PNefsWOF3m3LNTKyYzYqIBhqEiN/o3poGTEMVYgjsxh42i0JT32A/+t+WtM5QMAeTF2i4
m96N8UTrs+YW+MsViwZ4clE+3BVQy2JfIqkpWFSz6zt7Vi69Unr+uwTBaA1PyBqOvOpQrlb53c9c
RXRGK19QUvOwZd85zTRGF/gVAeyoaysbAziIggblMnhfIzjDV56Lxb1ZucW7nThLIqDZo+4GFKLG
N2ihYAeJ0ZDmOV6HUuoNjyi4MacGqFt/BwEurGaX9/TNKTvk1ppLp0ZrbjrbFmJqnUfERAAxAivR
XdF3edlxzxRe/ECO9FuRU9OxLhFvVsS34NG3AtcQMklAHJtkL54Y3xoGwj6Qy8eoyLZ0sJ34tx4N
JM99jLqv3uWKGcVTPbDiBZRLqHmKGdLiCiV0Hka/dpMhm5hO1LHfFIU0kHkSwK2y4Ls9Q/D7Ijvr
Er6grnvOotSqRBa0725jc2vxeRGx1zWU66Yiv5L4QVE9hQE6Ffl21fZ+WHvPPfYE7IB+HtHhvqTK
RRxah/9ufzeq0ggdMGwFSWWqJP8ZzzJQPulKBZE2kmkdDCRHP6BF5SFCbiP0uiJbXKaeHTJ+C7wQ
zrjMqFGDomS0XjmvQwpzuNu7eg1kx6dBQJ8bOASwiH1f2Iy5JOBdEgMby/bPPXPl5DXlpG3gC2Qq
s/plj1ER+Ee0JuihKBdpu6U0Z0y0/v5FEUdsek0AwrXkSoNNmqsWrA1jYFGhiA8RnGdOIPpVYMxK
rFkGhvlXT8DwnszPfh8z/GVbL4SIzz1gkigp3SI+TlW8dRsHP3FgnDBgMtmThZ+1iDEZIygt6U3I
L/oHSla9324xS0Ni5KyeQmiBLtvnB7IRFtOU3ESV49A68baO/nda/+wBR31bs8x99h3E6r0hKGAy
mNVwe30+d946AAgklKQATtvC2rNWIXF11P7gX8buek8HiD82ZAPyX9/VKLe6gmDRagS10jkucVBL
HkMffc8hy0OB6/1Frzu5Zb5Xnpg6YE21H8vS0nvWFNwHXTB1twl8NmVxPbAadfaW+mp/FVaMoytt
xIr44pLMrMZi/UvwOFTCJWWbEC8vxsDJfU/pO2aTv2VKat225On7XvveUo3GCo2/sC+jXDb/s1lj
YEZgES9W272LuPOF/S4+QiXBVofSeJI8Purmy39m6ByQCN7bBvwUoI2ByswFgdppRNjIlW3d/noV
mMavRbeQMhy+63ixS22dhW/SC7EkplSJaJ0MuXrfTNqBGx4cdUUlaV0XuufXsavyfLQP6Zv2arRx
1DPzF9cjqRd3BHz3K78st5F4zYWthEzl2zdagTZDqS9bTYLjrE3rMlrAFe/TUhcjb5GJWj3N2ZWR
wccvQSai+9rn3HbdLdWp4rDBlAvS26fqrSGkz8IlAKt22mEMeyoCesn0ASI8VZGTMg2GtfBvBdsv
GvQgQxRcjqFEa1VkJHHJj3ruebZ/QDOlojqtlSEq8QHhYptegiyvYZ1eVrhReQh7f3HMG6nThgWg
y8mzo2s7qgaknJm22uR+Llz2xl5vJyX0GQ9IeWT55qptJ/QZitSWq3jqLkqqEgOtHg5oLOSjl+SI
7hiJLn/RUUzUelolA8g+ZC8140hr8qAG8GwYPp0VnH8xEy7qzCg7Rz89aMtImzJbEuZaHMGkqcKj
qEm8d2lNDCPri9Ov1Qy1ZO89r4UDjKMgNX3VAx1abqkBdTZk+FqE43DKO4n4prbxDQF5b78qllh/
5DkSi0F264Fu8QINl2o5s1PHqkdbDP2LYR2RiIAb3hltOI+lOwWAA+mz4aR16dqLd5OaXBtrZsFy
KECHTIHLR3aV1HGUTwZf01UlzpxjqJO3EeknBnH2KwdDN8N5PP3t0603uiNQsKvXjPCcSH5hkL2O
pIOKpW2lHvcKKBxXxnCnRvt81pNFBq44YQzuZIRR4kQwiTtFOh7ftjQjeY90dqhEAzUkmUhDgmtS
cr0/b8AIWyWrWodBlPosmOOa3GT+BD8Do7P8cU+kXwU2kiG5y4+TsK85XVLUDKfL9N/Vs06obJBd
NOAWKd0FyRiZSSe9xruel1kbJYrUtYcTPBKQMoH9UU/ajnajq69I/t//wA8AoUSzvbB4tsSaVQqd
hr/JJNHEI/2cWeOFcGLnuHxaNveZsPTBB+Z2VfnwAFQ/IXTEiu4n9GyhNMwvom83Jh7XpKkC1jm8
PI5pea6/1KUYQRzvWGY88uJlYRHvBmQ/wka3FUYzX8aNSF5Go9RjMnpkjoXriQ41Ymanpee/pYJV
uVeZum+6MUs1vmkK+OUYlziwqeRw1Rbb1HLZMpkv7/NZKe3lGRi7Z6HsstNbb5iyoThKDsXzr9pd
soKjz6HrmcY4aXX8J2gMjHcJpbgX4d0p1FnIErQgWyFXsDSy8UpfgcU4R4xrDJl+S+3N8vULmQjT
RRujXgI2AA8gO+mXOH/U2Tf1lwt8CcB5wM1xG/0igHpgKZ8kXov80IZ/uzXW1MveQv+JGdx1Cz2a
pM5Q+RwKss/0LykiqUKqGKuux53qEZhb67IOFHwFX4NQN57u9oNbBUbjLzo3+M8kvxsQ1S2z+yBE
sxnRR7qnfiemowiDD7ey36eCmLfeY8t/pSN/ZNTGsoArk6r2J0hGm/UUbOOAxGxrU6wgxdCEaSqC
YftI7PdEC+c7/HsJVI22/xl88I02L1dH24GTH8mC4er4SuoDFx/70udl2h2brWfYlA2/ZLjWNGnx
4QkdY54V2YZXCpSQXpgEMCxOW8cRDrNoA9Cra6Icj5EV5GjyMOrUAuSBH1gBgTUczA5kwb0t+LSB
RZB6ic+NQzV8ozN+3BCJp0je+7TbT+gWJGwZGFNePcji8Gqz8D1xBPmpR+HBNo9nm9Ez1BMnrpSb
92NX+LjmkI/ooMa4KRhBDsLZM6YQ2FOub6KqfYX2zouFve6nMXRBbWO7YewSVj7UY5cyiNSGKTYn
iVlpNEmmTFrE16J/6gO4h1pBMyGgp6raKMhJdXnT+DgUrH4zGYaTN9zRfOe1oJGsjRICCPGg3m5e
9I0rB4DHveLbiltXPbjvab3gpgIoN2MZSGcvkh+Y6ns5z2oiNmRQFYYPT/zULQqSb4hZYEV4aAdF
ZXoNspIQTYjUeJRfCZ5OurRi4OnxuiYO8KrCUk3Uyi/9I8bdakQnJYnoWYPFtxhfiit+YyQt+x1O
R0e4slJlvtVtIUBXqRg/dG2SwniL4KUfdHKV7nUijsznseaiaPYzOe8WC0PV61DQET1eOMtrUUJO
UU88Yqmtzv9p8wKGeNP93gUQcXMURMTJsMxzTGNXowkSxXksTdjDkxNVVtrLJ3CuMgIqtW/Iovzy
z5Y/opH1rt3ytVf3n8Nb0Tto6BWJ9/9/A7wTSAT72uAxOEFDjDRaLOKCYiH1iiyiSU6eVj3ad5py
FglawF8ZB0VNC/UJx9vDkbCwOtvB3h1TTAOrCGbDf1ArmYt0Zzp6Oa1aWELzAxLquMQ/T/HCogyE
AGB+ZfKmsTS0LhOUe3LzcZGvsafqmzTivXjZWf8jVq3vxDTXHORQTfcEqBQ/mAqS+0n1IQX/DiJ8
7b5zR4EvsITpjzQbvgANEHU8uG1yVHA7uueihgnDt2xSL3x+0oMUUhz709bXMfSgQD75rE5kTjuh
UJq1Xbd01eHQmBvUiETncQkIiv6wHqmmj0p7cHxRd2tyJt+AYUuzNfb9AalrM2ayI2jzAhV667eH
+ZciXTgWKHvDXYbS8sx5p3iY+YQtTe2C7E3q/g048sE3BjMLspVOFYgIWg7Y6AgfTsg1TNynx4EF
e92MdX/Fs3mVlitj8msi2MtfuEGv6bjLLuHs845p28fxVCgKxlHtr+Eu/cgJmSLQvKgvNPA0xt5n
RXmzcx3/xwpVwVAuVirGvfVNwvVYaCZByvYe20dz0wie8pPTgJmEiSU2NvkTBE7EcFwvgBTAfqat
ElcwAO7LSuRG9vd14X8p/B1sLklxrc/gCnnP1h+0oTDzMm/AhMjOuzlYli9kkWy9XX58O/b7eLYR
9yhu5acYMySyn3tZwFti59cJa8cQ9PRQd8GJRe5B8Oizx0uioBORSSCWa3IdCLGuS3uV3i8fV5Ki
9txpZJCM8AyAOP/SJDZt8m7Ic71we8VPnSUocYA80dqWsY2e+zrFAxKimJG2h9gzS/1Wp1UdvJ2B
HACHTlviUwQ9HvAcxpWV4V1hlhOH6lRGU5MP98fLnO+Z/yriE8M+Ej0xYUeqwJnDx+KeVSN9c13f
rw/gfVYxc0r7o36D201It4VjT32EekSFdzc0WgQp8sm92IyNc96M/DfOT5uLOHy1KvVuawDlzr4c
JG+vyXTyOvHEiJqEIs999fHQ0QHxNQyI9GMoTQEnVEI4CGJQphpuAxq5np92i3Lt7CMvm0Sx39aI
mZViFzhCCwetGuMpRbyio4MCHkZolN+R/7B1wJ9ABkUWccEl6alQUhFU9NPRZJIJPGzlCj3r9xfW
yScRmxaXb8EZVMuvQN3NY2YyYCV2cs4liNHAO/rfRKXkWIAmwJpKZ7XCzcLxXOd1sysjWqTkKY2b
8plnrODPKNpAdYwu0f6+Oyg91fXdQ1dwL7ehjlaActoqGH6CqM56xGwWYpeTs0qES4OWDDA4qDy+
O1P36IfktqoeaWD1C40HPAvMuJXvnJyod7iW3EEZyQZ8+UyBWWBhFz4l9hS0d092WAMfbV8oxtOz
NhNbGjacuoXJcjL1IogWVxnCjLcwjebGEtKBsLjBrbOEeUQFD0otys3NEwmeM9ISIHeKvozb5UcI
nOWQnBMB1XjRIgGwvQqrR83QPScQfWaav7iZO3okZC5tcaQvYBvcp4Ic/7K36/6sQAGr4ydcYkGw
t931QoMfLq7HJfgaQkO0tAG8U972FZ96Plv5qk+qRvb1SuvEWXYidTHxtGzd75BHnHf20Os+CRKf
obbJ3Dl2stKA2GKZA2PbFiNaAJV69Oz1la34iP0V8uqFz8xhaO7mgfB+xb6fVif1XhHBaZ52lRCk
7/5VN8sgWD67SI6T1I4OSfPun0AFwc59byCPSaUZAfBQcGx+9cG4UUKNxOk3O/dwhM2b3vp8Qfsr
M4X9UCYcfG2QDv34v4j95RrbAcqiEypQo1tZFf8Pc3QgAjkxv5YCGDuKPKVXbf7pQxRzO9dTmbBG
mulunJ9qOh3cNbun/ms6CLFk9Qvd0iNW0WRTy+iqtmzLnpjqud+c1AwzUDNo9Lfgk0ZSOagRA4fv
NrYdTxWVh5ca2NPrhiYWNbT4H4gMViBxJ92QnCIR/+fWBIbBPW+XDHgnzMASGv1s/E714Mw0zvCG
VubdlV5S9D6BwdvWKQkXnB4x++vMZQvqlrVe7HJZsvXNDXGtT5qsMEUFICOxbufyMR9L62eMsEB0
5B3TM+DjKiFLtenCOEnblGzk/7QrDRnOeCvnqsPwTYonQMXhll9vbZ8C4dQNklbQLmddbWQGcoB1
AiTvRvWLE9C5dkeDMA83g0m6ONXDHmHlCGQaAPDt6ln3HW2+Rs/RmmWmtOIbXo3lDHIcNEvq6wV/
RJVpr6ZCSRtDkPN6Sw/IackRGM7suZZS6pWnhIWzhxf05WZOROR65s4T6OFtZVNqcIAxK5VUD5FY
c2hA7tVh9AKJm5Y6cH/Lc+5lxHRPtyKZIrJT5jrTxONy7VKWxMuvDEqjrtwD2d0YL9axPmZUx9nc
9nEFpJKQz5b5/5WW7TZFhFdGmnA3/ol6TIEcKdeg2b2C6cjD9PMzdRWOjI60vxATb82ic6i40PRU
GgoWYv0SRUzSx/jhDl11O8/oo2zpag6hNKhiXnlGj2k2aDb0/VTBbQeDjuga6G6z8xYipcYYt9y0
gzV1VxHeQRxmP/5q2CBYzzPyw8m7+3fP5eVgAVeOIFX94oRIwigMwMi8oQSQZEwqaKetYEs5vAg+
5+HrMfFPavcOPtF6E0ZKH2teJqg78bMU2xs6YFXekRNZJCa7VIzq8HRSqGtvwdRipc5rxoI/DxAu
UEZfl3dERzq6FIfjupLxecr1ABzGdKiPCkFfqYF22RfNaSBD2gIlGB1uTUdfKMMWnEPJDTG4qMyW
83EWWMhFi9GkhzyzVtUCqQgTiDrrp/JAsT0YEtDcwEpHRQp80XL1oSkw+bntzXzEE1RtpWQpZHyh
qg/Y3z7wqbmjZg0K7p8LfsoYeBJnuLsGqGSMdb17/KijSOShsgA939evK5KAypee2iE2VAxEvn9n
J0u/0GC+mtDILMIpWYn1zRp9a+EbPjbIeWmUBdQYKhJsFv8BcFUiEqBBpmhux6LBn9pqT+bat39T
iHzJXfA9c3db5JNpaFbI4YTRqebaxJan5X9z67GkfhK5RyApESDfQ4uI+4l2u41xvAK5Evc4lIrX
EzBrYtLD+8ntQYErVDmWgHqWVx4v0kczYlTbBOh1hNCEnSaGphEn4tBrbd2j+niNsG+zvXhfl67O
fdKvCITwGkeOF1GgED+OcuFO/386E+pAb9t3TWw76ERCh+HPWMH1SB+b1iZTU7AtbwdFwA6TukKq
rKd8b41HUoruXguGj/H6JYAt0tto/ewefu3rHs7nYn8fNuT9GU8d6Nozl1lym6kp2eHWButY0Qb7
f4UhOXQ4GpjP6OK+LxmxxiIfpMRDQQEP6mHw7IoDAbcCRyWSHw4EQe3ccZjHKO0KTi6gvT5wv5zj
FWHggRvR14dUB3PlzbD4GmTk5Xyq2uvp0Fk5BQ9gvI0QzfISqvMFL9lpiq5XhABWmk7YkXys2fR/
g7awVh8rPc8qPsKI6iE4iqsJPJJckelG31hiMfd4/apITlRcf6kpOlRU9qWFwIIsetgOViOAMYy3
rEbBjQJEZKdkh3NDWXWQAOwluEJZkTZuvMD+wlBAE5DEkjGypDURzPrD0mdXYaHEfWZjTjyIxUfd
EOfa48ne3uCpUavz+GQVcD0kOFFKwPAuGOjPX+6OwYz0rEGlCxngtO0QVpO0SSWp8hb7JCQwmb6K
6CUX/zxrNcqAEuPkdTtzJARFVZ6cSsnp1iCWONpGDexLEGFK0nR8EEKfGV2LXLKQ1Y/bnzVhbOsM
3M2XuY8FY7CrGijb9tCyBXvjGEjpcP0MRHVkCr+zScExwqHkcfXYOhFjn0h8EFuZ2hr2f1ZhKSvt
TlhqBKiO/PfJzFPVPOTvpE6RCu8g+MpsAOjUpRUL1ooyofRleVGS/GgVlyGgAJ2cvlsuzIAupwG9
pnd5zi3Sb5SfixWyhIiCTzPi/NUKvDHQtgg9YHJkxF/y7YxTnCDpUulEeF919G2Dfw93//XPowDN
k5AvCP2XSKytYdq690VpHlnehJ2vwI8siZ1hhYwyQzlpklvyp5AeYRsN/OJ7evcIwD09kCNW3mG2
eFeofrBPbKpHXhfZixTQE7rJJNf22OJVsdWVlgPhSNCIac/Dt+VsOQQCxYFG+VwQ55n6gJ+PCBA8
7FfDJAMWRAMGbcPyne3LeMJM9Yk3AlRji68mpr7YzCXUv0t5ivX9bvXnaRiDXp1HYGLMPy4IyTJa
w49UlQhvlNvbVGQeHiUxcM0oAy7ral8AAwWPoEgqpKG8q7R/imZ4lU3XwG3g6wZssWwcU4KSa0BW
7IccIFj+Ux+NQfJDfrSjzCIjCUvjb1+efz+ndRKAFMJqDC572Wp4Ddk8ILbf4ZKXol17v35SB5Jw
PaP25r2zRXTXXkuleCLCJGDEigsNJZhut0LdSIUXTwadtoE1wV3xnD3iqOrrfjRlcJAz586tjYbV
lAw4Tya77wKj5D9TaEBV7OUcmqA6UDlJYF4syTHFM/5Z2clcZxLv9r3KGnTjspvGPv6U7AJb30+I
V3CskVm9qqXmQPA9W5hYtM8ordj3ihpjmVPv0RfueDL0RvoDrK49NlOvHxygJG9Evt3wQqqhy/vF
cYplHtXvC5VeVNbLPa0f/nuOqV9HR/ZNhGClnEMTYI8QplZkhI//0Z9MXZefPY2OzaG3nVsq8L+N
iFFJfIpCpn9tsGR5XyoC7dihTQIhlBgCLQIXinsCfAz3xd6NuJ4LVMzMJT+0ruEzAuUX107g2KdW
FNIvzpRLy7hS2JZRmATmEId8F9qzgt0kVjXjhrgZYMLw9SQrKMSoafOIJjS9bW6O7YCGg6VMrfZy
k3/KfSc/QQ5pdRt4ft423IwlcKNkMEZHM4neeq1W4y0UQAyxsK5x75nvhErZ9fuBCqvimNQnDj68
DsDxiVhl2oTZQzu5OrCRczGO1soyV79kcB1kjzdlLY4wqBdIAX7B8NralLdwGEVfOPUn4MZSQv0F
mTy9IKT6btXtYGgdtv3S1hnBHDX11KgTsEPmQWDEH6GegjUtjURkZx+XN5Zbjx4oDvys9N/L5JI2
IiUAqRcAMGOY0GmxZgkvfwN4kRWQ2AznFc+1V333oDkozHgHojRUSfE1HfJPBIiG9VvlK/gdRCU1
2Uka5xAcYpEGny/OcFxKLe+komg1ZyBz4reUrHQi5fMwi8aczN+rEBxy+3pAoxVRLOgDuIQxPa2z
Y6o+HffzdZyuo8IaLHgCF7ixYyK2J82cI14q3cbV/BduBIRT8qcBfm1WBMri0Wnn5QJP5gsDOSQI
0rT1G51LmCfDoCT+EdSYYCveotqFmwrsR0eXj6sT9IyYMMkk2ULB9EZ0KbQ/S/G77jR10qA98wlQ
QiS9wjBcGFf3hEnUu0vaffn7w2HzbRK1ja8PaO3y5ZA9CfOz2SDKTtQ1cW+h90nWoRa8acbJw2xB
xYaGzElph1wB/zz2+7YDGVWovrgf0WBGL9oTzyD0fxrNHqQFm6LTm0v+2E7jSA85cbanuWLzQpw+
ZM0KFAf10n82/x3pqfR0BJ3F1CBoF6V/UM0vAfvsOak3tAXeXUDmTaE9ccrwJ9YDEUWZXNLn9rid
s3egCynKQfzbv52MD67Xucvorgglfe7xkGZxvvocfHMYtjIbbne1ZhavKsDtYlVn6lrfTm0k9rqu
QxbgwYQneLpLK7qa2ywKt0LFo7Bs7qSSO/REaTQcqXq8Q+LVwHJ+zv7R82+xdQm5kBD03LEn4gJI
+yZ4FxgQs+bzqDvsJvRTHycaAvyjTRaP/YsxXa282y7lShpz7KHv/6VANq3HQX/GlcHU5XEm/CqA
mS6Dk5QsO/C8do48nuNINdEy+E8cn+zvROhm+eYXHA27aTfQp6H+t3BBXqbwQ5hbXg2z97cSxA9q
z/0RX/RfSOv/1B6/S1FQPDb+glN8TRCTspJY6qgwwJ9hrZWZnN+5ARZjayL6WE83xII7bBdssSH6
/BlF3hpYzzCcknupCr27AN6UFfYiguFNMVxme89FBgDKN8HBA9czNLDK/LQBWuU4tYLYIlDZxaN7
IpymqmDEF4O2aLIcIlzC7Pw5PU5veJTEz8UVE9g0urjKhco+OdttFNSluLaCrB0jdHPw3m+kiMbx
gEY0zJ5aAgehAejLSg/K+3vrAUwOk5th2q5tr25E8LWgTp8RdKOdWfPLil1FaZClCKWVd7O4otRE
LW48YOYy0e14ojgbYdVIsySbvc1WAqAKIt1wS+8GYUXVXkfKiIi6QCBC5N88ZnXY8cOFPz95gUIe
L9iHqLpyqMTBBjNU6lJhFN34dqnoCnEcytaYN3CzkIaisc8BvPZbciQy9W/CnI+9/UhZJcatTsEQ
bRB5gyiKffpAOFOH87gl6BrFqjPpiPCtsqAEozIvcELs1nBKAC0itYlS7FjShnLlWNcR0BvQNovB
E/hiFmomO3qXNuemmgltQ2P2hZeAIjkCxSc9YSznYPDwXHAvcO+taAwqGSGpYLiHo8NX/aOhKd4P
jVnQsgyzJbdPPix5V1MuJVKKvzr9gIEs9+HOiXTQK4kcKfuEnr1IndYVVIyG6dmNq2R5/RMLYZGO
Ib2r2Ke9Q5bqxB94W3PpEZWvm9wD9pdAOD6hkcBkPj/oTjqFOq04IwBK3GlAvnxUKBd6mRcjhb5H
W3SPfjC2z4Wcfrri7OFAuYMEKFSR4ud4b//8Ci39Ys3cuuSBa5ZzK16bJVs3gErGf/GyOjO28b9R
Y5DnEiwiakoaxK0ULMEnVAMRqW84fk2ymCiebF/7VBIYh878qYRfgO4owfwMNWQG6xltHUzNF92x
RaTKLwv7n2qMG5iUz4adotT/tPuSCdf2Rax/xCCtQ1Ky64Ld+4H8njmEKuyf9D4XSR4O574S9usX
UnTYKLqFm7txvkRN3j4gjHChFBeAftqek4OADSd1naUkJOd2Q9g+1asNjy3Xx82OfBIruN+0ftqW
k6vukj4bqdg80FJjsIaRc33KS0Hhg8XQ6y5lUHDfMetKbwfJ2jl40l9uK8oYwceu5lx3HsIt3Xsg
gV50B7Qjf0QkVErA8LDGQ3u99cpFF7aIoHsdDNm11mrd79EPNCLyQe56mCB1yKgi1PgoC5J7Rfiy
k+m84sK4M6RIP+0Za1Ztk3mxsMKNoT/OjKQnX6bgWrYiaWPuCcZBgXSeiibJVx8g2ZJcE8WhB/sy
74YpjvVE6EGjCmI9MqDdnPM6yuar2tdYfITwK+4IV5k+GMldqKT8/hf+8bAdGU/keraN1qTVyhJl
+hU055a/CWeq1F/Ide+pmXWpvmHsw/2erQ7JxoWUZgZAQkJrdS1Pc9ptJNzIBF6xqPqKFW7gZf0S
gNVMdQ96+VzJLLFsYOJoXEB6TtnTIBEWI/LhH1IGDnXazTtOuKwaYk8ZB1mx9Dk/onavX/rXzbQM
SIETWV2I79OYkaoBImx6vZoo+MJ/lbb3pDWczvJ1ntoIjG2dVUwiIvdZByYFrk1QT8cpsNKYqV/z
VsWBz2YcnWgrKemdoe1gVbfzlpXLOobN8CWNcnCx12CNC64WBkD74/LwNgIVmONHhzU2zybFuKlZ
lC5ANksWAk2reNevoEJafA7DpoJmvpZ4fBNHBO65Kyxi85vsxT46TUYtGjGevUvdBb8OwykxK0co
oxmplQVm9XlPLmX8rcfXWk63LKvPjucKr2jjsPXA2TNQs36GPWlwhbERFXioWws1H6/rDkdfWKtx
5HU3wNYjg7itwySLfNt/wT2M5vmo64GBYZVR2M5mCYopiO8BQVkjfn5b6IJlQ404LRJP5S6d2JKN
Nz0A+IU+H7BuCLsKNPdKiZ4Aie6j2UljVbgcNGD5GDWOmNzDIIrGq9Ys2dgDMtBVbWe7wsCB6u6F
/NH4g9MMRlNG5dcRMk9oYozfhLrudvcR67k+PVyrcDAgGUVs9Xoi/62Kgdv0mZG3CRmEi6ng57Og
eAX8HlYAkbiFquYcFSJM0g6tXRUjm5a/fDsFaaqS6KntOf5/mNqVDxs+WT9FK8EtwKH97f0fBXdI
0f7/Pf88wo5Beuo8O7CM53XOs+h+UOiJ5yFx6fpFX66IyBVb2HwYbmdsvmjAdD7Rkg8JslcAyjWc
/dZFjE8GH/N4cA0vToANHhY1uoyML03YeX653m8Y2I+MEixw1fn5iCdIe6+I6fRBExBij9QXHyLG
79lkWkSuqF79455SI4HCicSlDBOHFk/7YLZo3O89GKobQtBqdcynyr5ytpdJIFy9XAAH8jAJx8Wa
u/fW4rem8VrrGtNtUUw8GfK5eP5k/k9OOWK+2sW+kdoe6tNls3DwI6UBjIR1xhvOwaazBT1wkZOF
uDnrQFC8V1/OmUwKbUa6gGmp/QyssX7+0nGJ07hkeylT0exm/vQXW5ITbF0HohZV10pKZyS/HYC9
VF7SD76VVdcUlKJaiRH9l3cNhv87a+0pDBnDSQPairPjbUhg8sgUwMifaQonUTVCO2CgF4FbcIqq
3sTqTr7uYicVmCPWLlOSPhGjakzgyA6Wmh21sQBp1ZcwEbzhwhTIHNIOtxqkM/2o2Z3y+I0DX76Y
g7+ZsY8tUtuLqliAP0qfVbKpJpFcbwaG0FWKm04elB+Nwr7dDkjiUlL5zA0Y9IvYjso5ivRk9A0+
S7/AXjV6jNj76w9ea4qZ5vpbWw12psndeccewjFhz8OSsLcS3Vn7hEj0pnBGxUb4YMy97aA6S5Fi
+UrLmsGf5VbvN8QeWYwl4S7af9Y8h6f3WpttnOT3/X/7ikwUfxQksYY35ptXzb6jybdK9wZYDxxu
QKNZCJFhQN+VjNDO3+C0h4p71URbvZv6dPuf3Y0Ny9AcR/xsD/MPaj3IvOJd2SFTpzteTblHeOLM
bwHJtmiAtBh4oQ+YUeVctVbs7tKFXJ21GtQEaEpxqZZFmjXwuz7DF8N1NrgZxPvwCTbMRT1adJhj
QCCTvyL4W3Bd3i9RsGo2VEfBBoQEbnGT5uoqecsLj98tIEVnNpLwLvTOL2CCrgPwp0jyawS8mpT5
B8LbWlbNB5mPjpBb3h+fE4IaEQIaU+kolWIqy0cCa2isZMp/j3XitkajnASE3LKzFvfqor4Yt4tc
3ufu7mZp9DiAcGGyX0bfqG20vLUTNXWa/P7LqoO1+h4V1+ByZk6Y4ig2M1g3/9PimVEiCEDA/cLD
3evRvtxWGPjRCnSx7o1mku1EXvUO0SaFxQcKXELx2Jy7O3nuRXElSReS5FDSIhmxjqYkrA+IARdr
EJCmMpzdQqJ/YLMavdlxdwCMm8NK3e4zuOOEJdUlGanuwxl2syAya8AzLX95EHRmNU4lHWpfRSU2
ga5A3PHi0Bat1ncdARU5d1Bm0VRoe7AKtvnDCHe0cd5xST487YtJsxHk1N3SnJd30iEMqVNT6ac0
vQ2ZwBZC4LuHnhixcxIYVGBANqUBytw7wfRM+1zbbYL3YplwV7dNi86Ge34fvsRz1MZDNC7aLW1k
b6VgoH5+ihUyLXQUtJot8wAHX8oLE5bSCEmzbRFUc9XeLxRnQr4XeQIIT93qZZkFQNm3aKycLhRv
J6g24xdCaBHzSkhol1fiXfYURG9hh/VVfaE1UhRkuyvp5BB/1TvjxX0ByTysQHons3bM2ImYPJ6M
ttR8X/VbmqkJHcLQZH3fr0hggL2qx7BkfcgHWaDLFxIiwGxg0vpe6ztDZr5tc7o5GYbIQrybY+o5
KiorZUHay1YQSYaDL06C0TZUSN3/EFs7MpZuKuQhA3+8NmLQazHm0nMnqMjFR5NrnVirWp5LeuMB
DJK2epuJHhqeSBaCJjdBfrgA/lJs62d/nGM5oMtx0dw+rOldzc+tu4in0IC9O8RSVLOzpz2Gpmyq
A1TrUSuyorrGmxfRIm9kg/jGjjvLjgcrhVXY/9fQ1SuXlso8hOW8PzYKNZjpJ7ftpknchXMY3ouX
qrd+sV3PXOSeWwjs8d1M31BPW39sSh20aTPtqmh8MuSKiBiW5q7YuxGC3bBfA/vITKBOdgdj1w3n
Hipgrp+86PwxsNvj2TunIiVuQjnAhMbJJLXtFD7PbVLVGTey8s6qa27JLy4SQxthe6Fxcv8pFIax
wO2Lf4LcPTl1pqUJ6wm5ziEHu/YnfB05C6Pl/+716xqAAVV+XOJfvaHLSngEEa4d8E/vkaqdiota
4uNfJOYAMuY1GuEngbbKowqtyBIOpp1IuhnUzw9qoD2eyWHLGXeZn2lmxmgJvXnfZO/N0SpUpbQY
rVWkg/V51bHkKaQXmEn9fWwXxh5gc5TeL+UBkE36whKmxMq7q3+RlnyEoIRPyev+D0ZYDVuuAl7C
mBpP/9jFFIM6/NDVfeGvpKeRVDlK0/tYUsir0uoAv47j3as2XqWJQ3Am5jf1Fu5880mu7nh0nICL
XaUOU1VNje99p1uePwpzeLNq8uZ4ePjg+DWvcoPCBhb1WlltN5wnuGE6eVtsNyNLbteV4tQ5DQkK
QMuwC4hoN93naMpnlQRsy7HPRYY5YzxgtTJv1JvW53vJYgfLrQUgt+ALWxXR+5fzLp5+iov7rL5F
QJnt+90h8MhOw4NQ79cGGu/GO4FUAeidg8ft3e3g9hVN7hvD5gnUMbPydEshsAZqzQGFhhLEbm3g
HBZG7ASQ1LkJXuHgO4+9xWd9GbbkCML45bkmPvT8IguGnExmNPHdR71TAvD251+UN8qEM1VOdrm2
EYPbFIyfOQ5T5JUXzU6NyzosLugDqwDrkVQSubVKIjqNpXJSb5FNq/nhH0bI0iq6AtTtpLRnbwFZ
cBgQdKJoRH48x2GmOwUgX5+syU0HJDtdG0y7RVaZ8mvLOvU79HxpXprN1Ov5cT2sUZajOGsfP8iW
TXCubr2buId68rIGUPnDKUcNBiVxuPEZdp7+2/nkm6O+vdPqXKY3GrWHPUDFfelL2fNypjS/K6ky
kAbJzcFRV4xEjTa7FUrEFCLA8jeaPjTUvu1LltMejgYXzjtCbCwYeZOBNvwtHOir8J0RwI/g71/k
8n1GdLmOsIfM0w+DPAVbZmHpYZQtItPe1f3pnkM/D+5iESAgpdnzXF8TevJsBKuueO10Z4118nmH
k50Owoiyo4r9dxmbOVO9ovVbPB/WEipdx1VaB8Upinl+0EIjJtm9uDf2DaNJK6WTClBRYNX0A9OC
8kT4ZlMv9st+pCW3ae/jV2RffdSzKgNLvUbVpv0MaSURyba4zVDTypjb2DocELYyR4B9p9S1m7Zr
4w5zoDxq6fPtXrJGWcofHHgDVK6fQgCzQaohNg1TeMkvi45mK9Yuc3qZFmJKaoiIYs6stUDyX3sI
oorO11hojN0WVs5SRtqFV78zbk4hXBoaRmU8VvUMpGbSFHyeuKBKEyPf3p0FfKDOjCxooRydyeI9
HFucYcya9J0hwKl+FG7qy2TX7pmUNmWFfksfL40mdbOpLsPazdabeoASUKECHRO4qDoWcaUYapmV
o+KLLKsbaE6xMtR/mI+FFQW1D7WGvXSAGhqBxXUbFh8qBTxkLOvmiL7pkLYcOOGvOnNTWiiWg3pH
u0UmazG4q4VHpsZqXAdyFCpxid4RA9Dh1mnpBQofc6gxJYINsbFFaGNomHtNKT1FkOESTU77eBcG
+Oj5NWkYydwjCONgQP62T8Ofim0mS2E5WPRlw3VYAsl/qbPEe1/az7ttnOFDUcpKxh0ttAVvrSCa
V30ykehR7yk2EHnLvJ3JpwdgExQkAg+IY5HwmQ1PHcPKuTRT1LYjZARlmO8uqGEiz36Xgy5SbMhg
a/e+HhpAAo1NXgLgKqCPoD4XPYOyza2+VYkOyMRtCir8A+sLOlyty+EP+ab9mFZrbi4dyHLmwQuk
hJD5SGmXKGjplNjZ1PlEunPqnANjnsXmvae5kcZnZmVyAItwENXFwLyGlyE3PET3153thxaNlEXF
wynPY3N8fCJLN1rquggJFLwCqoQhDB2iicgV0BIdqqYUZASaZV7eMyDVyT2AUPzRd7+B26Nch4pG
dqzSQMoFgmAMpdSfq3m0x77DjH6/98Eoa3mNjq2+uCDObHj6QDlECwsyzw686OuJTp5Fmzd6Zefb
4aUmBaXD0kIlUBAeC6c9rfy3ZgIGTLefokmzrbistQ9FQLcy/aif//IiYeSKoM5D2acNycumUaC2
cCvH68cFxr0v7MOut/LRS0W5g8jFTbBm6IFEf2n2T9o9vu+KqBCl2tJBoFmpCHrCmb2e+4pePxyW
qLe2uDKwo/I6G7PmZiwFvK4BUFZeYYFWelkfElFKq2iTPnF21UGHKH2dBLozOeR4Wxec4BFcxEiX
aVegINOSZE+n3/qV3mJS73a7QVdN53zHF8o6tFEzDf2WJTbx9gXc7MMdqWd913C8/Q1ejpX39Ogz
6fqwCfmXe7tM3Nfbb8yG0TGcLgIck7dzjKM9vSgR4Pho6/rSw1C67wAFpPl3PaViOkSy9wB94rmG
8CQBnf6ZL//b/GoAHBA5yaHa/TPUM9eRU+0HIRiTpwN6v6s/s3lxUwqL5TfClxizuTiYpBvTzdVu
oFU5bcYMP05Ne8vldq3KMSWGoyVT9jj69iAf7hWzqF80fPFEeSd7ICnnJHdGJQM1NzH1Xv3XrVqo
oZ04csUwhthLdl4/dn5qMajW1HG6E8zf/c8Ji0rjBL4JI7A7mPUiLPov9ikAQvn+oa+oHwvogIo4
EAhY8ORJBlkxNjs0gC3u7wIEENO5x90U9AIJ9RYE/pc4t3x/t2tKoVyA7i6QyJMXTXqH8EPPjRxV
DzO+H66XlQLHyvzQN/hefO8p22yQR2Cl8vViJONBlaHZZ3LYnk47vuxbXNlIseSzXxblafrns+V3
nqG/d1m17YhnBN7X4XOKqnn8pUr9yCCMc4nRZLPff3TYP1xQIRzG6qiqY2lySdxSWe+arTyo/Ata
fXOFp4bXt5VECBxLJ9mGNtaeuCjI6j3tFrpjAt1P6Fdk58XEoZHNm6jsYKJGha5p0uUYxyN70Vdm
0KRGAqSZ9RFuxXmlwQ5A1syF0apPgL1i92kC7CGPjeL4H+1OzKjl0NGy1EkdxZinSPeCRT3Z+Z5j
Ek+eR0KY8hwNEb/l6hRFnropAYtKglX4f9ZFafIKWEp5fgOXoAgpaW0L39XGPmlIY2VkSDmJgvVE
GG8CXLrAYEh1QI+r5XJ64f1YDHDrOfdtACBamcQLefbWPG6X66eZW+TiJb15uYReoDMNazD3i22A
iZ6APgcaGbNoJtU8sR3xuhLG88X7/kJQj9iF7X5FU83ebffxSVHK4gUmVOo4jmKMxtCnsGEHh4ky
PHCRPq3JbR+f944Ncb884igmAySQK93dQ3vjKGjyZek5o6qlVCXbJ2IMAb3q8Md6XJuND6jFf21h
a/48hjMojbF3/3rvXytmL87RAbsl7T32jDRW3DnwrD9RYjr7U+W+9yWd2mnGhQaIFq9M9z7k4x1K
7FxRTlc2yg0gXcxBf+h+p6gUYK6V5SyV4Kfv586emvulN6/xOg5LprY217LBSH1WURsAZN3qq1rO
0JfZtjLwmMSRX4qna4T2gLQFTAg39U8BNpGK/STYy7+yvlPPWwe+z1iBnKVGgCDjks4X9zt1uC/w
Z/zuqWF2AI7DA2CD3FGKA6GaFq5rp0uKQwo0JhTD0HNcZmqL/WKERh68D9J4tKlBXeNG1sl+QegD
4IqE8tj0w3XcgoA+1T/C+nnXewASegQCoMnZ/EH1DGc23eXfHSYZfo4pVB4ui60l8S4QzVN5gBzD
fTXg4n0maj4ZdkYOvzCF3U2w8kauJ1v+Qm/jgKD7Ee1U/autu5P9voD3bL6VooHA3TYokFUJbBig
ta/VBNX15JA/MkSm8ImzwtjZp94+mNezTDxOqYP3RpX0Cpz5/1lx9LdQ+k8QdePite3zfZxehcFz
QxVRRf82haWuk5GTRNVbFRkM+NaQHQR4OW6VZqMniBwIw3JDiFGcbef7nJ/urwA2XsQnNiF9UZwl
bSYLFiUh6TysDACf6i3UzWrhLwG65Grxz36fuToRWOlDS77QvhPxc9mNXxwpUOV5RU5N/+DnXtcG
m0Y8DzMWbfrJx2TKfXijjbcL+CEXmcLQBBdisxc9QZvRAxGo3G94seMlC8r2Ni7fYBjxXZxRDOIl
ZJiMcse6wdqmBJ3aJO2qV/ALumPyj7hUtuFqsmgyVNX3VLtoQ4GALZ/yWKJ6YNa0qrafUqfFeRrU
TVzYOFWqsTsDG8Rjf2PdZsXS0qRoA6zb35wCKqX/mTSPtprhUqv9ooD+DD39+aELw9CyW/+dpMJb
WUdVNf5x3oVrUllYthbCZWP5v++Yb/Ru6c5m37KCK/f41juGVGArbWPYV1/NwqivlRu/F0wGK3Df
BjK7SN2jjjizIM5wif0NE3wreDx8UvwnPLMa1ZRXUgY1tj2dWKKWf0cqzD9u2SkzIYQ/3x90YmGs
iEJQ7pweI78eHoITGlcaxyHyz2mz/RBwcdD1bYggVpw6tMgkbHLBO6USB9+Osz+LSL7+IKjzM18y
lQQKR4Fyan0IUo+RgV3r9kBW8D5QCs3JsyVlufZhzrxWpA5wghqC3CtV+9mD32hZj5gosD2bCG6F
y7veAfXnbUr0M5MM5Y0HxNpfTHGZO5w2poQOd6PR4SwQZpK/QWVcIfIoqHJEJ8p1U1g6SF2iIUzx
hVxDTcvI0jd9QNmvEcvlKg6SRvJQGbFExUfH6tKhtbEKjjkvlUYlVQNV4HrhZEdHcM1A6X/TA5/G
Vq0ql/G1PO+qnkAp9UVjIACgy8frdk9Xcnd16HKGKNgA8zOIWiB0gcnUCcB538lAgQ8A94I26BoX
6/qEtNP2WdSOXA9V/IThzg1YO/K/iHLC7qzK5mhoP4C9jhW6rKQm1X4iHFClNWrGK/M5op5mQ5By
uqTCckpB4XKGVUO6T9JWmiYUCPvB96limIXFo50nVw4//llGHnPnyeSmQcYgw3wimn1ZWoekZRh5
t5CXzS1hH7wpAS9lPEJ8ZxLnoNZ3vaevzF4AbRbMr42vsV8oBSfzbEsAcDHMSABUSitHn9+Zkp86
8V82iZL8P4JtAfPFtjz9dfAvSWtsyU4QaYDY/+8CYFODK2vyjGZvNKBw1kB2NjuvlFwVCUnEjB+X
RqK316wHKtxlB/O6vZOwts67fnj9DLtiZSZ5krwcWuxWiU8zjkYFUD6ViFK/dFmZm04p1YoT9zku
8ZEQoTBtXwBLqUdjkSgoloo9+Doi9/Lbv5cL7VMbr4RDag0zvHjjP5d6XJi5peR7cdlnKlvnZ4nZ
h20AQOqtSx7YqCblJVnSqFsYtKqq2J7CoZ4rTdUpx8uBJHMGsq4tJ9hvjgLZQ6JAR+O+5WDuj1ZN
Q1n/g65Lu8nAiaSs5h1UuYsFNPP8H8SuxRorLajevukxzaHRz/5D/EUSk9iM/2sJ9fPrqLgwsBNI
hW8ObIDULucbTorF7QM2CUIM1mo08gxRP5ZGHHmvR0PLlaZVS9xxaf2Xy+4g8ZOJi+mIs41skT/E
13qmeu3ainSuLjWWeFkEPW9rCQelcwzOKm5/0OymarVxdix/D/6qeBvvvN3BdYSlvMbky7A1FqKW
ENDWxXDlBK2+52ptAGFbFaeNF9dlKWAmdsxf1mkVC3pOi2QUaJoB99RueR7IPz4eJYjnQIIVoGIS
E8X0BHs0CVNgC+vB+0QjZ778I3POOOLjxWU4ynQ460vM6fat7WTXrQZPVXJHX7JND0aG9NWSfJdn
i6As75GQAzMLzcwtJxTx8ixSG1X/nZ5GV23TEM4gOt6ucWiriZ5iYvTqJ6ABgL257HoQMV883x0n
3IovW2FefjHA+KXVVye6nFzESbKcjBtDNapmOrd4vpMqaHlu43o7R81Z6NoHnvLBOL7/Rouerqm+
LkJtNIjA+9qHt0IV2UzOZEGTgnK7pUSrWbnk0WD65Vz5ZvQy1lVm6StlTJ4HPZQsBK9+kyz6VJ6w
fb4G+1iFIYN4moRqzd5GzfjDsJrkybY9wqfdWbI4HFHTMpjG6WRgWFoqVLgmBbi/QLNdsU7CVI5x
fFxV1v1ewpGZzOIyAl+Tr6Z7c8EoOQPpSehdKj9YfnGen023Y1fSBSjKPJwvFnOYAn619exlxnpH
4dDtaVNLWN9MnVNATlAowp6WIdPg+B34rUU4OokDtIC54/pHY9aABCRGW8YvTBlJ+oiWLH3edD1U
1pYoRlz/cvZmFAlhwjEGEgPosaSJcqJNBrF2WfUQ04f+9ZdjpmRcYuIsIByRFdOcsXaEd4zSwqqL
KiQL3A2fL//++zyCMmzTxakLdPVbROVAyj1jYFFYppHr5ND1lDSDZkFcLgtg0jnbNeYWsblbvI/B
buOM+KkFrHsYIxML3+9gZuq164N5BUr9YbI4hlxuPArBPJNffzeNrhABe+IP1yQ1Xrp0rQuS/N1C
rQT2gpnx0XYxIW8uy1jVsH09TR6V0CqfBpHX8DRYVefHm08VSHI9KrbsOK2aE9d2S6ppaMzkVXmP
e1o2Re+E/plGnFWhNHUcaJdi8kpReihgvnp3ptX/gJlDMDnGMuGvuJVgWUhjd7acIrLAqYUJnUg5
OmG6Cl6TwzMho30AkuD2B57a4ZWhLhVQIRdHRz70MbnwPufLw0kLk2WvPdwsIWyn8jzXzrAHOQnX
7vmO76MRa4b7ezNSAG35DmokrKrU8MK9okHboADaEpkDyXeCCJ8xI1vPsCriFsZW71DbF0sSgn6M
CRu4wRGr3MOUglVsANWwfTjfi0c1oe3ca+br5st5z2CK/O2YwFk2XVMVjung9FTwWyVyoG2HCHr8
YsI1vlbSXLSKuKHW27zZQGLfkRhybR3CRi19nNFCdal/rnOUTOxXDaavrDuypF6q+NORZD97YyaL
0S+tsKWP9eyMJWJCy6XqDWiyLWIlORIpaw0ULnM2wdvoeD6AdnEqB3hkyenAnRIhhKM+syarPGVk
4ICBpSkA1Yo6cQws5i+9OLMij0yHW/Al8j0GX/BuiouVvP7kDPcvILF3tTgvfutMpFtp/tTroJF9
6y/Vc0X9BPUoO5gD2CHne6+qnhZmIs5n41xWTX2VvALyhprOnwfw4tfpK6aSQMemam6bvvnQQ4/2
RBukLAhTILLo/fGVzBgVgrjyBRZ9tZu2BjSSfRdi8ZZqOlSI76UdtXQKweoBwjDYP/Qm5ZneIp7g
GW9kRE194xWQG9Xg8CL1LTrbHp6kt5sVzliHKdPzJUJVk6sLr3QXMeBts7Ialt6/I30Z78lyLC5V
/fFn7rj1cMg87i02jw4C6S8nROOYsc0cAqkEwcXRLSOcVxutHp6ds1aEM/TmjRmQIz4eKAi+Fio2
eQUbedB8NPuJ7a57vrwdpg4abpZYuG3wv2SwE/8KOSt6BhXiJ4oCiADnxq3etkULjjB/dzzexC2Y
a8rZNBhXGdtqRkAHvivdquN3ILdO1DYTg8+BiAW0QBz6pKS8IScgzriCeCsTmGQ/PTY92tZ/akt2
mdW5GsDAekGIndiVlL271TFu5XZG0GrAkRn+ri1T6LBXoRpEdgy9McPlAft0o+11RJMgXS7sSFQX
+zv3QYq2MLvh/I+I2Ae87vP1zsExTCSWguFPHKVqNCVl0ohaKzQEpaU66mmBKM2tFuSDaAGBlM48
jQV5uQIS9pLu2uI2+84hCZ7XJNRXM/jTFeEPGV5UVJjoSESZmTGrBnLVp0xqYtxhRt3hhysIUFe0
tiNmXKV9ldzR4c3hbo9DQsmaqwVdZFYo0Rdck5SU70/OeVnf+TDuNI8WvjfDUZB1LAdzU3ng174z
UkTHwkbHo9H7IZk2kjBxssoLVHcrRy46+asEnbTcuOTQH0DvpMJFrEtgUlyuiL+Gtc/0u3JgeSWa
iaivdVUkoz7fjfxc1RPu3hzfPO0r+SlFs3tGngzGzbCPh8W3fmmMUlWCCPpS2IzJf2S7RhuK/HI/
TYEM8dsU/m2d3HgM01OJkpn17WzCZ9qfi+lQgbZ12oXItpO3udKCpS2eCMKMlpYSIOBpK64evTFQ
GPWXAa+un369yWLVg7LyOKEEcuaPnwMfRc0LrI4FvWq+nc07u3f3+QAKfj6z6L62t1H/bvlRHsvn
I5E+iVlmN5TvvuOmVugVXpUU+fa7+kgJp5FOpXwwU9Hz3hYhllVVxhq3Cb7sgUD2uw+OudNfSkyl
/DyvUfe+itLE4gZl8xEzElkgOHub+MCGqTY0P7H4jCB+VWv/W9RVzzOaPY8bUAl9mmvzEncGlD7d
x/t883v3MnQJYmt26pJOwPnSNjqTWJImb/gXJN62vZgDtFU0wIgD7MCZZNAu+VEwcG6KF5TNbmY0
9vPyZqmo66G8dA7/5Y5Tl63ypKQX4OBatC5lPUYsR+gmL61DAjaI4psF2Z8qqg1y2JvalR1EG80R
rw81dqQUhJa1zzjQe+c2tpSlNlExc7OwTlSwbl5afNaCz3AyACQpVY1ZeBB52G9zogLJ3oI8vsP1
DikhzXfhE0qe2A218s7l9ULoLeGYIwxMy8hxvYBDoRt1PO8z4ggQ+V6wC3W35CNl23P5AQtdqqRJ
bp/x32zB383cQFZJNrBUtJaOtZyw7gBQnBopt3gIxIuLtAvpGIc9+1BiEkJwtUTneyvcP/vJn4wl
FeHaMmKxHWUbPy25rm0khTi+nxDH5vcEXwtqvpiPcNsZwPG4+JKxdXqPoLInKt5frfEigV7pqs0j
Bk2NGkRE9cjhIzdsBlLPyeEdjddAu8ArEoUAaIEtD+LEBG+bQm1rL6/IxBy6feI2b/BxT/KHlMEQ
HoVlDceQfdCcNil446lD9GZVDDbQUxRj4GZ/6ZkWZyJdoEGsQq55Na/GoAVw7zmG/jikJrY0A8vN
CGSC+m8iQHY2clVPrIWvXaPurkMXF7b1SRPXMPJXDtYTsz+W8ZjMBxBq2ZcYuBxPLu7ejkvgjuoJ
HiFzxlsB6vSs281TVlVobLjpa/tVC/MirXK/Jaa7sncUhxXGMdukohSgeeEzrl1FD8rXVPy603gQ
MdKP5D60mZBrEGIWHPx/tfRFNL67GjwKBTuA12vWsYst2hzsGCV+HSAuhgpY5Dmt+ayfThzCxUGV
5OfZCnkeSWDjSf+Jz6JFAWMILneHH81ZUQVJQhs0pQD81j8xysIg1flSIKerXeQnl9UlP4hmsyqs
twKBWG2HCZq04GiwciqaId0E7Pjw20YqmVbxCNEyhL8YqOIF5RqOWpM1VCiRELSoZCqbtcDxxQXH
BwMvsFg0b1p6xL6egmnCfG5CnClR3EnSPGZy7BlY+YbN1NqTkYyGnV02rpDc0jbABrMm/bLHdfPf
0rWgs5riWN2WH7lUqTijs7XN2D9H/eBKbEqnVKiuKU4nz+vlEirW7uQ/N9O6Ba0AiVThxxlFdsqW
eAswqRpTWCV9DaQU+UyOg9ihQ0FUK21N4IeLYluTJHMUUnU9t++isXgJCIcD+O67pMsGbZBufJnC
htMHu8QPUXguBgAaUjQpEKodZLpp+dYXXQjbwMlNPw56cN1zsBSbFXvBifUKT2cRT7VA+/S7tPDg
tHV7+1OJli0Mxg+ea7oa4bUEVurUB3TdZNsolytMczYkkAJ/T1k1H75J5lXIGRgu/BmtuOdWS/cv
3zDO+jx8JspNgHRgglI0Bw2xeRxOStSM6XDWO3Xs5e3v2WTBu1cB+UwBkOlEidTcZEyt0P49UGoo
ojw+mz7WVanhEBEMeH2V2iXAdkLk5anTAipobWD+f7P8aaTGaF/mUqYqlLHZt1T7lu8sI7ijRKn9
kzf4+H0594/wq2PIfSxBSPIiaxcJcoeqdxPB6b9PYrnBMAz26fYvRbativ4oX2r11u4lA6YMg7N/
Lh/FzBVjP9roLnQ9Q6gp64R8k3STeWvRwQpSs5KJZuDAPPivoSriiVsD5PEWKYUknY9J+s5++s+x
DhJenyFG9YMfZ5AJBB/xteXuOFg3E8mhsiKTYTDFJTK5+H3EzMExn+zW2pJVrI+GvHmWRcEoeQLH
CaDlpSPKtE750Svb2QGCnegaELo1eLP9cvF1mUID7tDVmkRbBCHMxF5+Z343RiBi0/g4Y3YlLaWq
ggwLwxKT3BU9ozkmmMzcG2cfLwUQEVfUuiLUAGkqE/3JCBM/OIb1oj4lD2/QaTpZnx4HsOwph9W/
/6PF09DKHsEN0/Wd/GRWdBHassOrE97Ngkw00R3cLKbYDUiA1Iv4L49X3Oshag2N30rBtftPo8NP
fkVH2aQTCzDecywkjLwwrCmvvgGChucRacSNEgKgvXbAbvlL4PuhTmr8u5XstDTYsIl/A7BwwHAG
Mby2nOfEQ5hd5U6Bd+4RzPsd1EZZEVoyAXYkl5p6VeA/eAQc5+Mo/9khzKUFGTBWKsEZVFyh5fHF
UTFfVsPqg22YE1s6j+LZ7M2gH2RZNcTDGSrlqo21FYVVOYB3C1iknae6DVqCrIwA8U/o1DYm6j8l
tTSkBswviBCggN8ptMHlSt/NnhgIaAM+vo/MKVRQa5VyJhep0BUYwiYEV7noqn8c4bi8Bopu6uvu
hGLXrojlbb094lI7L9RTWUt8tL/jT11Tjxz+IGTk19vO/Wk5Bi2BL3Sn93CCnsShFawOy7LeWzZF
2DHaw1emD+jKNXfduoRgnWhMSof22F8ap5L1IBKcEFnS85jGB3oMlC+9PMfJk9Y2xZWVWgcVEmuy
hX/HRZgp/xeJ3t6rEVmO9p+D+wZHEPX8wRGff0MhqXyqgFoPv08vjIxqMrzWa13MLWbk+YNRMfab
TIG7qTGwsLAj1MLvi/ZsOMBU5IJuuemvwnldQ31sc+S3n5YaIbCGxCxfxnInILHC4+bO/JLx6nTM
LpPsBpHLrFD03/c+uRh7wYhaEJk+1jKrwx0jxstuvhQgHM0GhqNWkO9/u8xZBP2Tly+d48U7wgh1
/1ty6iI2CD69WeKOdZypi9aQIbLeGxw913QMyaCAb8+KrB93wUxzLYJBwRx+gkZv4O14ypu+BzhU
ZnICH5ruCOvaZuLwN5VvAcubdwRVLZJ0kDm1zVtSgpTZVcRFanfMzmYpycIScfF/AUBJmHx2cBSb
J9vhe7hRLoRcc8mAGfUwuDfX+U8A2mOgEzaUxT69CVTyxUD1DWzzW1nzcSA7Fgg1CIIoOgIL9Gfj
GpvErWHIHAB6exXWnBtcWY+8R0zXdfsYVZdU5z9YTrbcFr689Gl9aDRpglG0e+eCrp8ScOnzvI1I
wtjl+X9HxAPuQcC9ZbFMpiCfLp0w+p6+lDxga5o4dNyuBZ8mOn3nRaiVlu1CGdsv2s2E3rRR8QBa
71ZHCWfJqKEqC51DIyE3NEwOyJbDunkSK6GC7c+9P50PwDmHFEWx/vdp+IdV7e1c2/rhAWbnD8ss
BgY7hXEqfVJ4OD4PWLxxFz9ov1xPIvur5yplsaoXH/2lHmggnKPj7TBvkLM2mxO306kjTFuO8eXY
pJivvOIGNIUm5fAwnK5yqWatsYUtZx/9725hu2CrDh2S9cV5FEyAn5fDl4bWo2e5Od3j7j/OgeAc
57SCplYK/uk4/rxQuRNIT+MyIStJHcdCwgrCyAGNW+bLcGNd3sRfR2vqIB+hSHO7uJ2PtCK3ck6G
nNUe6KTJ4NFCD5cyN1NFgKifks7jr3cLfAh2VJQ+5Z0i84zvCyCMXHujXoZojWd7Zn5rPrb8NWT0
ahcUskEslQwu3PoGx+l/i03zOBXmfwI2cJ/EIxgVfzMmAytdxH3poL0W+3+IsGcrIyu1GsT8Pjqr
XPGejEGdmUFXa74oW01yuzJCkdXxhEovATzx+s8AwSm2u96bKiHfnuyt/eQFLGwoGV3iq8FI/gBP
vetHfdd2HXc7mikQifbUlnOh9sbL4Vyc/x9KgwECgpzZCIQV0O1D3Am23QlqTvk3NvLEGQQcoebF
tfLjS+J80Y9e3vSWNsC9MnZgSG3dUkq6OwcHd3ZtXXEBV1dxkv6sZEBunao8vU0Box/NzY0dEVGO
D/XRYPHFAAxPvwYYL9OsMgXduziAR5ABoqtIjfEbYQl6C6MqdD5XKImZNIAeDaHC8zYHqogrhADf
PrmfLYH1WbKZnVKbkOOLqrM+pR1o/wLCC4Zzfh6uIhjrGfSGnGudHXxbo9l4WDiWX+oHpejUatBM
rVkHo0aNdyoN3DGDCCsK7PnfcaJuF6l9XiOLc6ZuJ7u3iw4eNbYUyIP+9/udQmSTea8O2IMzaeeL
Xqb4Dk6T0HtinA3orWzA628kF9CzwOLEx+ZrVuUiIPoYWkjx6B1PrHqg8X67IDUKk3guuHlATJs3
+KBTvW258oox/Z3gDNk/lQaBLh5oMLbIOUFqtFdqY2lmwjmcaRNVG7AaFRu6GT3zQdPorSzpYBSo
aT1nJmgKnBOo1G9UonBCkYhyMN6fAaytEcUHPK86hDBMhf4IITgXQELH6Cd9vPyMF5VUNMCAYGcR
tJ+AAZlMavw59MWd1p2WFWUC0RvRtJHWA4M0Q41RzFThpMl8o8v/ClLHvHe+uOink+rblTWouwey
aw20V3SBNfLVDxYe6TwP/eQFhaHFVz83uv1jUpr74vU16ccclMjx8kqQOLi3QOPkQ2oru5fP6kEs
4/5nPFSDhlgoBGER0Yidabj8CpvuwIoVMUpvA2trtT+KjRFB87Y49WK8lHmkoa7F3NMMOGT2GBka
b1+DkHuZ/EjUrLhNJC7oEJEA7jiV0sz14M2PwjIsxlD1/BDtBGOS/IDU80E7eqI820JKwUhJ9KmE
V/KUmr/1TrhtaY+yfWF6Gv3jkwb6ONjr/foxpurzG7zk0nvxInkebCNs9BcyWsdLLExqsbCAWjmT
tG2vdeMwiZDmJXd0fd9rciD9EZrFTQDywUpreB8CMKaHscpJ45kQur/AwL/7ImByiWzoGYRzu43S
gdq/LZpf3p+y/xgHkLYE9md9jF8Ho/SOsQPjsDUdR2+pFnsGH/E+VPPeNKHZvW+kBgbSviN/i3BK
VfOtABt9bj/i5QDkVveXNTApwSYyTqDbe7ydJkjpQFjrBjQcXl7kSYUL/KHlWkzxCFTgT1GicrjY
96I9/86O4CA96VyP1cy1sOB6D5NXu/MP+BETAJtSNCtpS3PpI9NwBopA8H9VTglZxMZDialKiEfP
M+WvWY3eHb/ahzwEPSQctgVsbtV0I9yixeY2QANCAX89SB0RyFSq6V9aQnImNc4gJfSsRQrItxav
4HfzcwgJ6y/Im2Q4xA4D6mBmBeIM121gtlaiU9jALQvayxWXuUk8bfHSUG9ieGVtlOEHYmd+ac8Q
PRQUaLbsOtUE+iJ+Pq/ryxJk3bdY05pHQNuOt+dGzWZPRz9lq4xGGQNxXf0+xjcNsQ9FPjN2IMlY
rYyLwITB1IKdk7tdk14Lnd/BByHVyikt4e/rT+EWAGJaWuosH8YeatWfeKgGjGhHIN4QFDQxPtjM
Pq2LqnwaSmOjmS6Icur3yYFuXCwV8FioQ44acFJBR58nMKfV2nXZP1fsrALOFiDRecHmDlUBEevz
0vatw7zG7lAEqpMWLKkooU1iwj5hQRnNo+TmuJafABp4rfBTLNFCzPCA75Ll2mSrOSyXmrWOlrrX
QqM8p5OOoFbnlNLgbk2+5FQVNFpiqKmZhIP3G6lRun13q5WZy1mOygC/bDnQ2L4y2zU71X4tPh1Z
cJiTXZ9TIysTJ6Wqau6tq8oC0tr/mtiCm2RE8ru7TBj/NuMnxeMfn6FIyZ8qSMfnWmjGT8J6lO1q
o+cUaxhH9Umy0w0rRKbbam5dQ+G0/bs4ghjgFk/e8j8OfA3d0ePXR7751GZAKyqkQmgZStVSyv9d
QZ4qYDQah1exiqjGtgTX+9xdTYbyO6aZZ8p/0ULlL9bXROynoEHGrrPxebRnNqtQEnt3/9PcdiJs
Yh21GuAVNtUVaHaHgCztmJsW6Cmjv2GHKkBcAXEU3WZvZNFTlhXce2S2ngBwIr3X33y934Tjp4IO
Cdtxen2chDtXpesue/MG+zRrQMu5kGOmgjkxyqGdjmW/vdaC33ghgdzuoSajj0OlhQehIsayxERn
J+MhBV4Gi0Vm1tUslL3QiqqL0VpqfAEqkSRauKQYCbXWmim+5hXYvSUk/ERXVHwupMCj4fkrh/2Y
Bxvh/citXaPypgnyuM1ch3v5yd7m4Nmu5veBQBr8ou7GDoaCayTjJJU/eNrDqH3/YIvpgTeBjpd7
hLLgOT53pVnmvnGht6WkW8Hy4VpokCnFdqx25Pu10VwspOnIfu1qATKlCnTQjCWN8iyXpF2tooWF
wmIBon0FTla6INQ5tW0hT980exhnvbfUZ7SFAkOxFUKLz8ZAR1OItQYCK/Rv1ZsZK/yRKLL+ORMX
TeX9eSG7i4/DLeEEpYgq47gu796m0PVF1PTF+kXBYv7ucf53KafhIDLXcVSUZYdxEhnDtfjLOaDL
8zp9MHBFHCU61wyzMxgakdYqG+f2fejTbUAIP5Z/8aK99j5DprhqjC+VS3WdpoPM8w6ZL6B6nO7W
IQ3CHN+KtAQtEA9ZBDnQi9iRBMnF4uYZZnRsm13Z2fmsGuTJ7hXr5OT+BpeMsbypcBCGLi3YpyKU
oNbw8p1NV88mcs9IXwNmbO6QqFBn+KYCP9te+OwZ+A52ULPxgthz+OhV51KADgShlcWhU6abAGWo
J+kxLvHwsi8Qr2ciJt+AHVt3WAmV9bP4euI72emk2AiF0NLCs3LI8aBu1VSc3MYhwiY5syIOYwkY
6mjzmrzJc2uDFKbeyXuU4GqTNVRo0tvc8ypSCQcyScd/j/iil1tMrUcKGagGQ+36SiavVUiqkkOV
aZgHMcq+nrNfpJiozuPuzjcCJpnf2bSb7/PCylScJRrxiiUuMhb7P3ABiYQI0cFwkwxrBcELvMyN
y0RWYKhYi8aXj7tXMeiwbRrAv9JFQKLu1V3Q75HERfRWqkF+UZrjsKBhOdtqDNP/4psYqSK3yqfL
dDtCpZsbVFJOLV/MnoozOKVAvAGgLQLZC1W+jjZ3Dr8XT7Y8Tdo+Fumd2Wbub7FIHwr4BWUvdRPe
LEIJwKM0Nl6vnQXOh8x13sYSYMmQBYbDKG5P3mIfp60K8qFFLlfQC9DWYOz5SIA5WEfYY/HMu8Ko
pNZKVZZfsgUKZqZv8zirkxUDyjl9V+8darsOoRfaHuWp0fbLeh3yc5a1VvmNeEu/vy+zmQaK6SBn
4/D/hMK+NkPegB5wXV8ZK+ucWv20iz2oagtlWJUflpQpmOrBw+Xk/Oa2nyvSguxwpH0XwRcu9ARU
gmPL5O5VdJaxJv3ay8Fl+v/o94jnh6TzPQq6jB/rTKevo0yMsvNzAPI2n+WZ0dmOfXDSrmu677lw
AMyIDFGWHcQXKvUeI2NqQEQ3L5MoHmDICOBxiU8uU6lZReWKQUbweGuutoUVKs7GPejDVb6tGlpz
/k3tO4FBr9vZzE7lzv778uoQVXYmsiRXpXu0FcXKsdh6q65MNvE118hzgocLK07CvtvG4uGrQy0P
6rXLPb1pWbRg39MLSXuoamgZrdMyfd1Re7zcnLSfk1r2Cpowe95S15/KXSJ4KLKdxvHvmiX5Qqt2
W6wfBcAUPl5wsuq+/CLlWv2lLXOrol/scOMrwS24t/YKZBG3++skOJAq1lftPeMnFqilFmictO8w
TZ8HQg8KmXKV1+WsHbBwlNXQghqGJlGO1qxQhHetYUf153+bRWyFtSnf6d1mILJ89H1WAUb2dZFu
pEwXT7fNqeSIesO/0184YQIi043oD7hfD+rUoSuixHjRRC1lBsyAfXAhN4eYkt07zC96ZTKMLi4J
elz2Nk0a5yfE6aaAABmc2PRBrPcHYveKefsLRP2oyKK84zbze7v9AQDOmh7/IWAfq8uD8b08+wFG
/JvvKyZ4UPtM3CcoC9uzJU3/Gh4zbhubrRSeOBB/CXlBfVgUGxSmxtb6MuwLN5QKnp/QGL4+DsSI
hcNHyUqd+bjmVWqp+d/cgI973IdQ+Kw0vpZWDEt+OKI+pqCulc4QuBl7XD+YoRpRqWAuImfukPJe
AaAgunqPSaW7xEEQvmhAEmkXPkphNFO1jco3DhhwvAzCGQYvmbjomOyp5o+/kOkrnUwb+RfwMTnV
Hil6c9Ddx8B8s2+iJuAKHnbvX2EhpAL+WnfywPJdldikFCrKFS9fHfMZg+Camh8L2OM5BUEqcLgC
Rhi+7bOly+2m93JJnLwiw5qs3HYXasT7acbMoYKOnzpw9CV9qakAlk2bDGhL1C3Z9jKRUNyvOT0X
gUSqKwNZ+feQ44yS+QvFFiiumNOwMcWZA+g4MgakY32EB0PJEriCzV06Hit9I0bs28gizFMOgBWi
3t487A/upninjC6xAQ/aEAG34QYVypL4lfscASs9d8fZC+sQLC0Pwieor4hYOj4eikwox03eZZZH
E4ccsmldNVXEjZf1u7HtuDjh7Ubm96PXVGQ56wnGu2WS3QcdbosgYypXzNP5c8GBcVevbIOJdPLz
Vwv9neT+IIqgbNXfxbLBzCcf0DS6NzH+eMwi2Dpj/RUlhyNgD4fwAyW96eYINf3nkSrpuF2RqRyT
K1VN5ktV9J4pgJbqWTVn81Lau63oW6F2nm4qcwUkPE8rjfaiEPbYvJocrpotBOZzL4Gu4rmgvOA/
DloUZRRxsL/dZ7Vuzk9h96NVsvDyj8l1itV1P0PdT/Lf14F8J3VPtHF7R8tqG14ZgnLbt6wN78mV
LY8NtSQeIFOYkCNA2euDYBGNI49yXJuQE3QSDn3X0LVNzoK08gjQFXjvamBc8s5ucGtZFrKToRbN
8Ad8RXboKE+hqi0KZTeXVKLMHVjLwE2SmIxYpLz1q+qot06uWqioHXrjzoWODOsThHPWIYDmQ5Jq
WHnJRg5lxDn9pZq6rss5HWBW3vhGTFYv6YiftRWl181p3gXuev//5aQOlzHV2mtCx1GcGt7lud7r
k0/WrPOFgYfIa+bfLfhfDS+aZfpjZJ4T3wzL1OyacMKEuHFHOwV9+zW2e1OtKlEiInl+CzqGuWjE
9Chp2qHCyQ9+fsxXE8DW/hNwGaAWbxuB9L1Nnyk/mbJ4xrHsuPWszfiVOpCwlu+pAORIjrFLzyQN
vhtPCOjoV8oOpW8GaERSfnOjo8dqVZCd+xDb6t+boNPAUgXLEdJAL9trwMre/kZEmKqGlAzTmkU4
q72V3+c+lfJZvQau/xWVqCRJlVFTuaxZs3uZuUg328LLmLKU+VWg+dA0WJCilQU81t7/EF/fgjXc
89j5UI60Ebrf+JfwTUIu4sCFAMb3dLdjQxINfIHnFAfGEU/bTWTF0IgqEZz0ad3PcK0haxc/QjUc
bTgqT6dVAHtu3dN54KDkgyfIvcZkuxomMJHI0UpAy1mi4yIuQ26SoXsjMvx2fDFz8GMVkIVg/uvJ
jVTXDR0CM00wUonx8YEaAzwQG0tQOWX9ZrUJArg1fqrDTyp0+xx8uUGVCgPYXFki+AwE1NoGKPX5
/BaZ0yyeUb/pWCy18+SyqyVywRc69QjYWwnIHIqrEmzII2I4Aigqqa2RtOR+ItUareKIJQTr3kvh
+AqsKe3KBW4nG6m4+OsZ544AByh4Mn7sTW5hlgY7XmEMmcEt9XybqUXotPGzaSFSPPGHP1InvTk2
grCLLk7C4ySccbqTRKOq2s6IkRzgff9jFE/rgl1KbPMs84mceVcFqxaRdHm1hyamw7/cfiA86aot
KFs9Q3sl3uEy6zSDUwnflmTgLNa8DTcABj1D1RHO2N6lNqxX7A55qsf/94yiDTB/kasduFJW+syi
4I/Oi6z4PVOcZ4Etegq75EEI9PnVPu4NZQJL4Yp4ADKNlQMP3ucaUVoj3Tv9lygVnO8bETWkC9Vn
W5ibi3BwWQf6EdSJFxT9aOkeaFQXiS2X1a06UrZwkVuURDZKnBXETWTQZYok3xp1kZjrEO496B1T
+ARgiCv8LzxvtsnIwN9kN3gCDFSVi7IZ/KoNRs5CWS4k3T5l1az5pfvcB75gogQxtqa1cdT/J/Ba
NNiez559a5tz6wzBrMbf8gCxkEtzrC3eWUykUGR0ETISwg6ZoqIzxqK+JvxXAViXqUrbkGV2kK1j
apRTlSGPLaymzPhYABQO0rMmT9w/SSPUObpGkijSK7sw+/SbDdSXucs9gSZkE+Nmxj/UVa/csBrT
caeGWqWBbRxd7S/ORSuSVRh9/UXF6MRJVFqgGVC6g6MUZV3QxkwimvLoI3l1xSvWmjYL4TBslLoL
2J19RLpLNYUXuR0oUqJhqueulvOqf2i6shgBEHft04woyRBequa2QSEFJEP8g9YLyyrWcaRMYS1Q
WjNT0eKIo53FTDkLKxLqv0R5Bo9uem0EkFk/qq8/rAVC1IzeIbl/l0tVRsxBSpGKCaQdd/ava3nZ
KKnYrDLZuWekv9AyQJXrrBC1yVXE77ypAhPMFqSfd9zRA6X147WUrJvaZ+cBFpqdlKePtXVHfAwE
i3csypC+5VK6O3b4VpNKaPdU17mBY8JCxiSQxjOZcE3WUi/iDAfjvOaShlCR8z/ijv4XLHddFvcQ
m6iY3th5RZFHBYHt03Lvk7GOFQEG5+YfM1p42sLrnIJX6uRJ0IU4ZeIoWV8JfqyHs1y0o8Vk/6/M
Ki4ff5j0tyhoZAbDmGkc3ZCH+NyzLNexUOjThtmg7/JXegxyN97stjPno+UoRtanKcCrCs7JsLNw
lCKwfqq5GPbNTPvjl9sBi+HHOu/8J/z/E+gOxbe/vRJJPoLRgPjD/Z4rl0ltbM6WZQ3UexpoXVlW
IQaSbXYRc5qUpPfVKo0fYsc7u5FzRUEr66Gv5lHK4ewJVi9yhB2ukcZ965DdDDwOz4ync8j5W5FA
ruk+Jd4UzIp7uUfOjbEEj2SZkNqoXUmYgwSiNs4TM9s6VI4EazzRl2Y3M0QgBjQ2CW7FTnZD5my4
vQxNR393dWMfr+N0UxmqKq4EiXkVosJMYB96PkHx47hQysl0/qv0ZKpVS8++p0B9rNnU28w1D/Mz
7KGa5h3R8CeL4ll3OU/9764mv3rw9Llc78F9zSV3uCSbukbLrNwmoIgNwyX7p8MEItZjfQbpL0o6
aitSmaBJOeyTRsIksTaWD1LJ2LvPO+uGm74eJMtqZIuhfD/RxBAvGN0jPlwffSDD8yqiWyjBO0wX
TfaHb6gsTX3SYNIhsF/vBLX07OWGeAMccHMvM9sq34wKNUoqgJN1zR2kEND4ZNJ2v9AWQXrGgAx5
vG+mBnOYJVgUmvwJ4MRFfPGpKY0WWrc5xYjBacOAetGvktHpjJK2sT92FxqGydWn3b8os5i93fLs
TwjK0A2o31TM17gvnqn+rLsSefyW4JiwqEyRfBA/1W7DYYnhAMsV7Uwvr07hLeLWCq7XgsAWfKuD
3u+YOhcBCyFCMkBrQkyzkWmMOMySZOAJLZYCGtrY2tHCxaX0ZMOUzLkmCtn2T6ZE30bXFS322DCT
zE19e6pa4S1xiaOpOdxi6rN6xHvljhR3SmabfShAcLyezjif8VShkvHhDCdobABvBEYMm79YHfXr
X0h6dVmSQJDk3PoR7FRiaX5WCZz7N6L1r8BEUxRAh9kK47udvLygO3XB8lf6R5BHsb6OIcWlZkx0
UzR3R7XQOnTRuQB8Sn4xGikrlH6R/nskzcJF4wMhv4eP7KVn23KmG2wmTF6+L2fcuuOHIe7FuAwv
G8ZeijTnOavuHNY1BgvQ6VzJckq3Y2i/dBmrpof6+RQOY+vXWItp5X9joNM0nGspcBM5xKhJWhxT
9G1UovGTul9UBOS5GPxY1iA6qxzgxoJ0T0CggEpkYDnw627hHdj1pI5LYoC5Hx4ezubAnNEvvLDF
gU8lcfldV0s8H5/lmoOR82JHPOsvK/fCRQRNetXq26a2+j7fcH45FirR1nHRSLUngHzHUjwDdEG3
d81tik3KfTYmQ6AZcEbkgWc2RbbRfsJvl5pa43blea7ru158lULxZqcQHjrfEiK5fmoHdf9NlDGF
vcBq5qpJz66/L2Su8GzhzoJ4UsZtyqDeXVVRf2iHdIki4XjQKiyBqj9+GHoJGClV8yeHvYbzVTwK
p7yBGuzQ9LQu2oP5TUho71vRgtUkkEwvlTA4muxnEDm7+RXMNSuTFP+/0xxLZyLxPgKvFIJGOBU/
u/fop07erCJ5l6ULdj1rkvMTXzdxJ2HC1B2ee/9YBxt0NA/C26oMaW9gYn9CyVHAxXb3afzPDH7E
WCdjYOhlUoHSuGWCdyK7xmBXWI5sX9Qm0HtBqXvNUZap4QVGFmHhQq3J6UOcksdhCoIQS3DuNE3u
zEgVoHjWr2Mx8Wyk4vhHdMceqmUzq9ZHVnysSkirj+jp9HxZiDqI0ZKa9zU6FLkS5y+5s6S+pOBb
mRayeCi3yYAaHQjTvGgIfvETW3ebgcGNSi+JPihlvFyD2iKrxUhM+9PXePLwxTetN2UzcSQ5DKYK
+Ge7v7YIbpMU0AZQ03ImRGTP/gqKz4lWHb1a18gMXVP99ttKRPTQ7yp91rBUd3EljeVGyZ7/OqN1
UYSxT58Ax6xPF+sKiO7lQKz+REJgzLW9HPC59Zsl1k2fPrZuWNUq4jT+twBlKWmbJtpdTdCKa0tn
rB7+GxUlWSnS9Xwpo+SX5dEuvdin8QnlYLE0AzbVXJ1fX4e3MzEXpBYslISFYobR/fjWKblUJq3A
Pevu6x+Dq79JtCZLcwo/KNo04ZAH1a+VRu/Hc3JaOhgyI8V07twa9mJ5e879ByvrKMz30AuNCiDw
oEeW1M6cxmhrrVY3LdpL/xaxU/yspbJH+ybUWvRNtN8JKVbcpSeoddq91p5LHMRMUCeKZm8xcBgo
CjKNibcfJN9+5vmdKUIcC5Vg35jW5w7cMFot3MtEIviTlI5A7g5RUELxEjyiDIPXnOflAGUMSICp
kvnGY+uDBAf8kRT7G+mfFESis1GhPrFQk9a2eY8Fpu0owqz+rg7eop/f/neJDGnxgr1l75/GrX4T
K4Om7PLlrE5t4THSYrLrEmvYYBboH/8ZFt8MAfx0ZRzcSR0QGItjoy53Gqxr2CcvDzyLJ5HM9kfl
oLtbqSvueE4m1EHedlD4YElsXBUJK/wEHBibOBq3fJ3RcHySMtPA7lUvVaG3arHcXmz1+z05T8D3
CGpNWGgqX6TYVBpEhoNUB/Oun+pdMUIka21C7kMk6NpJA4wiu3Ej3i+2i78Wv3lHzlxcaRJnAFZU
bEFJzCZuY0C3Ks1a2uJeC7za6URiUYBCfsDHIq9KboEKZ8hhKZuxbii1PXMjTjIN0JnJnG6NjYYt
P+cUldK3LkHz23KM2T603kYMLCRoUCHo/N2hAymFldpgw/EuClkRZus0+WNdXMhteQI4ulFRFBXC
VFHzYXL8QydbIqAsqN/E3C6eqd2BQRrnPG0c6hs8ub+yCHoRSNDu2eqSRZVT5JugAqqJWSpbKcwg
O2krbbTLW2B23mEnlcQmM8IS8SsP39yjTzzO0L450HrhFVyvftpR8sJyuPt+dicaFr3Asl3IABKT
B6Hq5zNNAF6UiEvufXlxWCKIkNyAcqFLKSMkwO+oe1pZU5OVq8RalE+RnFUO+ywb40b2Q8aF03eL
herr4GHT7KZK7mHnPbY8TxfC6rtt0MJnKA8OUdWhG44D/KTRzFvRf0rBXaCz25Yr3jgoEk00SiyB
KFkKblga8A8Yj5LjpWMh+JJb8F9kcm77fgccWOGc3HCr6KQbzqftn9yaORyC5myNUsD0GhxDnBZ6
a4HbVZQ8r2VJZwgZRb4iRmeg+GDe7SzlJzDWgzaNlclymV6FEI/faPUCDdBtONYTWQAubPA07aiq
Z486lpKxhf6NbojNBxF/s2NSjpcKkjAS+uqNOwmn85Rrbt+9S5QoSNHDnIycAjNK60ob3g4mwkAF
qyRJuaL4lyTXNBSU7wZ5PJJ0s5PprB26KGuduyMle+3Zncat3+IED4UGytMDwxMuEQa5aPRTdfyd
oA4zY5AEcv95Q9wroTBl7F3STVeEE5krtzbpG//kvlh4ZY2tBVbDRknKkKp+8vFk3GiiWu4kMz7P
e+TA4OnPh6HVsZmfJeRFJg668u7l2LZhUD6skyptKhL5HDYG9tDc4rlOWORoxhp5u9It/tVsO5/L
O4Hgqu39JUVII7yTYHb9tx+R2CQZZItY42jY4jdArBj6L+W+QENGzdXlvnmSH9tz7XET95DKMIVT
DQ81MGotkWispwwNAm8XjSYulgFipm4Nnpv+G+8wnGKK46M9pp/n34VnhZmqzlLOfSMa2CWrw8bu
SLXUznRb+a90lSTg/6ucpCdoUVnTKmg8U0+N1vj0Zw3U1YrcltaL3rpttCc8k4PHIdgkhRcgTZCR
OD6F3M3hFac6qAheQA1O33Kx+wN0jVokIylbVur8dsSk4/1GgqOoLY/6s9m4Zj4Xi8EIjN14xSBX
ElNdNlgPZ0YBV6qoUPIqNzD78vYSmL8Mo08evSGwpyV+TUkMC2g4J1jRLWaM2tXJLYndldZVBoHf
ET6u1/hQTokh0f39kpaRSEM0/bayJNT3HHiI9Cgo2h5sTK2xb/wCC4DRSBtQFb8AcMUDeVpREa5H
WvidPeuYJtWCDNQL4iZ98YD2pAGCLK3UDzsA3LthcS4Me0dnSAk4zUrPvaw1xdaL2Fb9mAhpVDl3
aPWIDuOvycP0hbp+2I3WfTkXvT9Jmu2Ry03etqZN6ZCaW2Q2HdKTXBNicnwuDJpxJD28f8Gf4cyD
dqhxn7G3eoYGGxltilEA6Rdko2rK7rT+4ERNRc9DjCtwRjIBdbIKq33f5NMllWqoK6oB9VQ7jROj
lmgTerf5RIchI7jsFxl1vJblAietLqk9+8ZQ8598J7t4cZ4FnlnsfHlINlIjRW5yQktNNFn6dsXG
WdIw8k1pGMNIlKd6VSqOw5ZGd9/Uqhek0Of9IasBf3Y0VOL1vLHF1ysLTCTJJ+EDkrAfSAaVLVsy
CYczp0+GV11+0Mp82svbb+wLlLBjkQTTH7KZGeosOHdJ5TlPg1b5M5P4abdjWySG+bSf2Zad24Sq
h4lBo+dStRX3dMvPKRAroiZRB/lmwBC4PKinx8CW3/aQ+77M3RI78Zc2M2uI/ON6ntN0Im5AQONi
qmJWdVSef1mwFntRmv+fXrm7v7ujSHdfvB6af/AjdThisudlRwHtWkoPAICSSarIfghrtBqNFI/B
rsgdsRlJUG/CAfKJlkhqZ4/EYEvS5AEoJv9Xov4rQmvkMh5DE9cN2zVO54EFZVDOSqY96zTYPijK
SfdgkYRPuKNryGR/XE9nBiHJ/Z57FKhuHqBvESeuP+IyCPTpPr9JLE/XhEr5/+4ysqThIF2XyHJf
wf0kDBwBxBzQWKXvUdOuGL3KviwapXqPyVcGoA+BJdK2Ut4pAq3wAHBOXLYSQ+1czmbvz28MccyY
9I+wOvId03RNxeVhke4O/I918pjlPZwVwrPsGZ0uBDn2s+y5SicnpGKq6QFx5U48cSR6nN5Rjezf
9TCtowtKtKyTGI/ofpS0R3DH60LIMvym8tRSzzEq0iVMQYg8MixOKZXlPbDjrS1KdYV2DvsYpH/1
+qyAjParxr5VtUNWq7NHncyHs9GlmuhN6mrNitL1MMg4nGMtHt5GqRg+FiNoUizkD3idRLe8CkLK
3hDmSWc2b3d+5LyhgBBb4lp9ar1cjhNn5Egiyy26wFiiuTnKY5KokQSZ3nwAF0sccpi5pgKqFnhn
ayjnbXy8DHZ8aDKATnVdT+EIBdZd56XgrBkCJt5gPt9uoPBZSH7dgyFHlAX726/TxufGwNxB2/O9
kSsq94GDDUvqIzMrmrnU38+06F17V1mR4xmco3naWAxTuKiWf77dMsXUAFwS551Vv0bu+ercBvte
p75HNvbiPFlBiQsTqwXinbHhSnxBHl/c4ru9RuiIm16k8ICoW7xcAPGdt3qclqQVWqrDV1Mq2NuO
9OuJZDrE4ZB8fC/b81zWaKFTCH8pdSv/ffzG9Lh6fiH08exTEfTwdO8lN5psTo74+4eFOuHAb3Kv
byA9Pmr7Hs8bbuDQ0K43+IbHnwpzGJhtqpTOJ+91sA13O1Mo1gUzoQXTCESh3mOmcJFhs6Ss4xud
9CbW01efhiAbjlNECAiCK3LJH27YywFrNsV8VMXLTutTewshmDWc3KWfl6srFbxhYbjB61DxLPIf
9Ed2s4mL5bSvvkPZj3tpP/z4FRMVUF6KBa81Jlse6OXDs4Hl2LZ34BD0a/ICE/7MFE/bqY4lKSlc
KkxwsS33ua+AzZOI79sG7oYT8xwXMpCIidHZ8wXeB4poPb9G8GOOSIH/L3TvwV7ER/Y1Si5AH0RE
/14XfKB8C4/4N7UNySSXbHlXgbFRi3rOop4SY4e/xHrYgZH1uYvTbiU7hSvB3Mu2NsoGND4TlngZ
JlBSRKA/a3/MqMC/jzHX5qdwZNuaefqvCxdltoqH1d18QIbWeF2D7w7OitJnxdRq9NSFiWW1SA9p
IromwlAuJQezplvQ9zt1hut7bNmBOTaAgpgv/IWyIpPMXuuIoyzMz+wsZdBY2trIaeqNsCTrjOdk
peYWeDSHVuQXwPSlZIyOrYlwFFIxRsc7gGW6NqnaKPvMPz1zCzu0lvBP3vaxdGmJ4cEb3Uro+JZG
ibx8YvyoHkdwaizF726wqHvkJ5IpzC2Olelp9MljdkDdvsBDbG0H4f/GTTu18MWivQhadHmOSs+/
aaUYM0EueK/A/a3aX7TCSjsVVCIsCCqq9AqzBC1MJ7eWc/TmLOHA+ylnaxD9kWgzzn12J6dyD/D8
4gVBHep/Ag9BtPOywotkSVLugxjGjydHiA9dxxwfw+RGp+2uKhqmAo4YbREY+VItE4TWD+J0jJzz
qT78gov106KNUYDYre18aZ/GA84khsv9824Ur2Z8Io6yzZ+1xGvpmTASD9RbsdVDa8pURH2gZw6P
CUSAo8PTrut+tU0vxD9xzprsx++8lFvsufqNk9Ed/ubUd2Uxf+hLFZwPC69qm6OucwUHjDDIbq90
qQZaKH/ebg1g5gZIjiue112QZNzLjOmPGWRYvuIfvKSZ0EmAEUWE368loQJO2bWmG29Vurz0CfDV
Tjd/JgEMMdJaiQ9CTEVr5V/+TKXiVR9xTVQGPeehGZ/d3qaMTbBD39I3EXz7KztHCG5dttRhgxrn
W7FRmS0+IEZWX9AOp5jU8+N2JMAf0sPHSxT5NVmVCD84q7inRka6piyeeAxK9lO5kNrGiM14s0VQ
iyrJZ1RwVsJi5XPzRLNEVCdJEqncpgNnEeqVTbnLD9GJnLssjKzlg7Sz1pS8y6djYxu+Ayz0fw/z
aYyIdpVc5RmD+rU5pfurSjjNb14hDsIfrnwz+ooku1vml3DWTKcmY2W5lbs7lOYyrCPAOSFJvJaU
8q7iqx12U8f6O7UxyZL6k7jiLLqHjX7m99NnOL5/9SSFppW4/36yltyeWty5UvfTTEELWKVa1B6h
lviYRZBFcOzQR9VWlmgiNwYOFt1dk6MQ9KYOuPAOpaQ9HLidTf4xYPc6c7A2GvNvsLBD+sxK2oFy
704evf7SEHlejQV0OKlTJicgUAk5cL8X3WPJSo9wQ9j9rIN9yZwmRP5UA9KWaq8gM49qWLyUI3tO
1LH2BIW8xI8HG2Woo8s2MGLpgEwc2Ams1YZSGDP1J0mfRC0fxeXVfAF/90Jn0MNFwEsfetgAzRzy
GKdcDNmPfYeKi/wJ3kbKr9Q3GygMwqtf5EJ1plTSUA4M0UP5IYTROlSnwvHL9temycyXE/f2Qi0U
4cnb7R8qGM73o57Ee+lGrO7LfPfrH9k+CFHh4/uBuRwDGXDe9CeClOZlRJ091X4tJuvO0QZOB01s
OIGD7Ny7bzrqXn90IhMOJpUxjZFVZIsMHud63eM+dbXy2HJ3VZ5zxCtNcS1hJ5VkaT3y/fsynimh
DGfLl/RKYbILn1MblQ3h+2PpUvKKcxnMEkuyp8KYq7bu6WlP7KeJdYJ9mlO38dlobxG+rAz6Jc5f
K2/VxwNfEYw11I/8tJTjGkerD9P9ksKHYrwICXAQeW8yh10e/JJ/qnPFfFL5OaFDejDkTuoqsYRm
KdTkRmFxvlptWhiwzti6iet46IE2fu6kvTiy+qroJzAJ6unTeXQKr8/D1QVa1R7OG1SNoDoVk24k
rXqJqIXjeylkqCR3bZluiaJ6VzhFdQVCaQmtOM3K0MMHkjyxOz5GNXZVbobhXwZOTdLeWfAi1OZS
W/J7lzHCOxFxlIQ9VG/rYRgQTYJYb0mpL7z5KCnr62hP4HefWlw9LHL2EC2bWL1ahRIf511xQHC5
0TMlXhdPlkQNvJvgBQFNksgHExk6limEopBJlSwhAhTEs+AbyUr24oTYSGCBDzH7MpnpR51qVMFg
mzhtysxnTzZYqCJO1Gy2ODF4t0az9HrIUJja4qKYGKqhtFSWewz2aJ6qmtPO0ipOUelrpSXN+N7y
mQD+14rZTB61UobWk24KMtu84UCE/2vl2Rm2JcmjVEX+0Y5n7TxhsOg5+0wZqVJoxKhdYa62mD8K
OYGS0V44gosG/g09DJykbSJWKRVHYxuPJT+zIx+8LagPXgA+y2+o9b3kIizR6ITIfc1pmNL/pJ/I
BJmv+/NO+EmDLRtAXVcu5yIzR+Zle6Cst6hrzfs2rL5/qBb21xL0giI0xQmF3H6xxYz1VFcNds2B
Ui/uajjmCV3wJ7ZVGI93FP3+VO/Qy/20aMUSKPjPMcWZFJuamozUe5ax4pLXZw3I2WFUUSVyhTHA
XCazgcjkZ1SVf1OxBkn5S2wCcH8e5LTSuTetgQXbgJlnhEVL0NzgoE2vrKsQD1nnyVze+gBt9Irl
mYcwNtkLFEI9o2rOLvG1JTvf9eE8Vx+GipAHuPZfbeDluz/r9LEmEUSeV56j+vGiRLenXDQB1Hwt
CzfpG7pCn8SRNrZfBNbfwf5JZj+Mz16TckHLci0vW9j2IkFr80XbgAz5cNIPlgq8Hn7lpzglwh7H
3nL1/P9slFOC6nNj0bV8cbUSuqiFXrWNWk+FQ7TEnakKm0u8epMgSHT52VyLFLnRiaoQBbG0UdAC
W33sMYHhyIlkGadvCKvtPiLhlsIflffWpPxse3zmkUlDvexyT4JgBd2QgFkD+uzGkJEQ1oSWddC0
NFMtUUtmpueIG3+AqwcqlP7GXhFtrm7XXhZJ6ZupOB85X0d2izwZGH6vwp9zypHqEqkDevFrPtaP
WV2umsJLaTJCei//0srmNZo8r+kYZPvj8ER8A0yJnCQjlBNE2DZ73+hB63GHyTAk8KKhhl7p+TKu
qYK5Vw4nrHEE93Qp3QCv14jV+HjElx1uLEuWxP+Nfy+GOu151sgNqLGYU9hGFSbpM0Qa3bp9phkT
pN0zXAKIvvWBU0WzGIXA9/D7WxZzMh3w1Pa3ZXSYvFOP1XXf69fpbn6WOgz0Ro0ESf2Fp1d1iJBp
+V+PzuqDBQMnwrsHI2mNe33JvoI6BMUc2iz1lk11wy5Ingte+TFxtg1pOuw4UXYeNyeSfcySp0Al
Jy60gSfCrshbQUIJLMHe+FNZTBfgyfBcZOuCZHn3HqEW363XS2hNhPVXJZP8d7u27BHwEUJwP0IC
iLUPv6peO0QpqlSh4p0pOlBD4of1gmZRGExFi4UeRzvJtMVwfnULGJE3QMR5GkmnoXTTugS4Ozj1
d/NmrCpu6nU8eyeOeyIqY7Nwit5v1mrmgxMok8fRGs9+eYEyi6g6/yZo3dziZWw3AlhCDEDrj0e9
Vbs/jioGazR/dulBxd3GmMA2JbsZm0oDG6mLGcTtXaO+OZAeqWjz+NJ6ffjkaJ5uAeLf/Zf+FFQD
HsFDTtfye1gE4pqC2jCpvEAviCx32qPXUIba90QAjUYYyGCQpWXQNzBgNpOfoSOYmvyHLr5Eb83/
MTfDnHXR51/dukA75Uxut5Er/mBaONTQLLAH4ea/wQ2r2QxTYwZcIdX6mMNQ3BBd2cLPhPm2Nh6n
DC6gHI5OAQO+/HEn1R93cTqOLZswG4fGL+xfFLH1G6xWNg2+S/k169G4xPnWQ8w2Yju1xNUloNjI
HaBt+mUIPiEGLNAfRKFKKynQ/H1vQMN42cketxIrAMXf1BQKAf5RTY0Cd1MSbwVGLtTSy9s0FZUd
p/eeH3FVYS34+/oFaiWoFXK6IdQQxSS/cmykWKLxOBkA2DTqY0oM1p7ZIkKw2E2sUd0Fhj6vebGT
CclqSFfft//wv7ZLC7itEWf/hcJhlp7aNyLs5BKz6MfpLLBLGZgsf/7aanIcIAIpKgAzyWviEn8q
WdmiZ3/7ZECsYKbJQ2zar6xiJZw0iiEOd6fHhfPHfPqx3vPijDgmRmZmjBP3+aFuBAqy83dB3eXb
Je587FEYYiKow1gFpuG2KDOdOkMErGEE7LNs+ojbGDGd9ZZj5JbNa7fO1tNf5k++NU8wIalqcJNw
UtQMv5Alc3C59gyT9wLWvcHMMq4qGa9cmCz/tBgJ9b4k+JYTqeRKwtT7XVdlL9GnPjMTXZFEXSco
emxONPxgcz4dcsXGIPRyT/hZEKZ7216QaTLNEXvB96nrZ3w7T/WwMowqrw9BUTvQ4oJ/llrlerBD
Fl2pza5sjdW0gv9aULdNREi53/XSHTqVXPJEhl6kpE+6Sjh7fo7nZK+zrYUOxqYwZoZXdFFIvOuk
SpesAXBZQd9ix6d6zycSpvXlqSsvU69OomTl2Abcxth3CK63tZCmNE0Qt1Py6OUdiRdIsQjexKab
8h5fdvtJ4Bwv2LCszm6+SlreXF2ampSC+FEswTYCoj5LG/8zlgMarXvRUvHvqdCt4pPmRupFSVxl
cSoSZGHMG/MGMHq67QnanLh8lCn+LfOwyYAla8lV8EYjUdlcoypnU3DT2iuhD42YZNPakqTmnbJ7
u6hhVqmF9MChh91gt/c7i950oIkkez9bm0kG2JpsM7AWrJdukjAVljAr+Vikxt/vYNEvJTnw9h/8
a9HEnkjIraYtpjKKcswAshDih1LEIq6Us1zms9iEmbgjCBpNgXAzEST7C3FqpueTJOnCbSNkq6R/
f1htQW7OvzI2uODu6QJBpiilVXCrgBaT3ErQJ6rPyJmjr++mO3oRpLzdrmqkciLqLj2J7Na1pisJ
SK3ANi09ee+ZhVmY7UCZOtZdY6qOqH8UFOViEn4cWM0QOChFz+gU6qdpm4ABmXDVXt5cqsYApkQ4
5oPYd23NI0UEuIIvqAHD5zl3DsWQOp9IHbfmHRlzNxXC/YEnqWGI4hH/lrC4i5Xg9kSQtlcpVFmU
L7G72fjV13YloYdSWUdlK/Eqz6sAPHRFpgbR7Urvh2vM7gb6Y2xVskgVoUm8/Xg0D9pUa7CsgYYI
Sc8CzaQwvL4h20O+whVgHqy5lQnZFgZ1I5o4Y0vlp/CG4eTT86DR3thbj3y8z045Wip+qAPFYlsv
0msHykUroFhJrSM8RCRL9xTeZrw1MgDDkup8BMfIVjHgp2RZAeSyR5V2XQsHIbQLkUIMcFpwOolb
zMgpjyKGyY+VQ8zr0/pOAg2BM1Z/yctZsD1kYxXvA9ynjay7BCVYx/TvPszpiPobiF7Q4sJa9Dgy
0aHSbeAdf+71rpC0nj256ztgQ+hRWCKNjwB4bW8RfJReZXYnaA3NLtd6qfrionMLi/axa18ytS8b
8U4zPYtpLnSCikdsO5neRG9Bgwg8q8kiblj54G0eZPQB6esjMNKFRD552h1rt6J/dSOcRXj5Ow5h
OtoSRn25asP57hC5Zkl/4IWoXPGvZGGyZqkRh5uML8q3EgrsisRjtTHJByyiGBMUTt1GyDYNE8hX
eGy/xrG3x3AcCJxRVLAUETyBIXLTHJepRAt8tTn8RxiwPpnXlWnNuR7CiTOla19xFAvufxk+S4MF
7AvVESgMoTC4P827uguX5jN1So8c4JbtjK0fUm5y9DZaBbbKjy0mzJt/1aCPP1v8CxPFon35sXLs
91/ROVP7JPV2Hk7qE51dPW+JyLhO67n/mePzu8IAWc+eF8+VK0VLdxhIiRWusvDgYuL84ivr5jwI
tla/7cdf14pI7mG0Tga2M9Gb8ANFPRH482MQRJKApos/u2aEjzsHBpdLaBhhpbTR7PbTFMfW5OIA
jN7G1azymBnTv/169uChK0ve7Pb2TaKJyIW1QOd8wWivUbkqsKQyB178p3PS+2MJbj/ihlnYujze
xh8+2WThxlTAY6d4H9kXYm72AOXI0CUHuvDCyrBz6pPIWG3bMozTmjma750yVrnfW0CgsWgzPQzV
QcSLpHHeO2uGCL1c+XTEgryKeuln606TqUdyPrA5+crZww9Ft8yNfZMmtUXi6IS16vqXwnzk1rzv
+qOQdldg3sKhkVF2TPcx1ZvAb37MrFTSwSjx7/i6mGLXjAUjWL1nRqrbUIJx20v1ObvMv1GsgiSt
8wIdfXvgMRAp1Is/MtPEmnqU+bZd8Y51uOajP2ex28F8/7k1rQpjc1crADgTkqf6MkMg6DYhfe+0
s62yRuKstAzCYy4IIIACQm9/USPQWZUteniKrqdhCjEYnw5v232JE50B0i3eKAVeKOIY4JT1NRo+
mZmXbiUN1raMLWftFGGWRVVn6r7/1SlNJrKE6On7oEWet+az+IRrGnm2EeWyGNAJQQ8TmZMCrXu2
QR1yVtb3vFm3BROw1HTTMCL3BN00pI/4aNcicJBQZpZBnlALWfv8mXiEleSR34SIoivBfCPZiDJV
CLREzqbk2qhlRnBqqQQiz6rLdmzeMUnYTJAjiklKiaU1MSRI+6ZI779fdRdWs3fiXkZKNhF9l4z3
vEaJFUzBmf9uvk1LECJY37JyfuTqL5fYs5Bsdh+2yng2cnUMa/OLPRm+SeyXhzdchMuDDn2YMNYP
S1/YDwPfmOGztFgZMzldkyE+ENZYg0AS4m+lAnko7tnX9PoX1YVI+wnSsB8jhq1kBoKo+F1Pqjmx
ucZCiQw3goLAlQW4k7XVc8ceOj1teQ3QlwpJQ/lY6d7uCWpWmhVV6bcNL2xZ3en34PgmXtyK/Zp9
jXG0ahmOEVNu4L/ORMJdz+QR7gk1tXbkWUjsGEph4qQmoxU714EDn2mGq61w4pWfMKGh824fexFK
NpUrK+ujwf9uP+IRXxH5ZnRV4qiciw6ZmdACaEf5ToXFBSavzSSSRpBi0M5vHWv7rbeWhMSWs7Mm
wxsWck1ujb7NDe3tmChoKE2qQnO55IMFTZxQ40KnXS7LZPABq9z/0P7mVLcDsHjixTVpLl9EBd1K
u29OjFDWaEQfJ+4oin3fJpge73DlftJZ0i7Zihrf6UNalqQE19ytTWMc4oBQp0Yi0Gu0Wd1bjcAb
QjVfXYaanlcIawNjKEqZQ6d5hXRzsbTOj9LaUopD9bOJAArExzLkIjRG/qRPEHEuoJOlGPicwVPq
LdSxZqrbfKJKzG6VfH3pvOfRwglh1qxwxmJu6wzQg0unQBX6xtfWl579sFKIEzy9OjH0UJgmmNzK
7YqcVlFS7k6XXoRnBrjBHfMbK9NsOPYkspLTtdjXFmUUpgpQ2HgyGeZICKMRjMGWdue/2e+NUKe4
RakHY9HD5p/o4sYUFezlVqS8Kn4ojMp3pwKc9urRCa8O+6V1oMMOJ+PsxdCvtGbwfUehy0DYc5cZ
czFFArbiSYr+uk2LQW9ZZJApQ+CZLeP8dwTJzBiNZ1kNoJ6mfHuKqcOw9bqkIi0LSAuyYFIzVbWs
ble1kldRmev4IRzItcy+tLd1BztguWVptlf8l0DvIsYiwXdSXxrClTWJMLvYLrR9LrUB0T4ey6as
lwznjSo+WPtGXDwUnbRZyVl9Xb+cdkICKwkVQIh7wlqRZW4C3eHHED2jnV5STivg+04ns3rNGCp0
hqZZHBMHNdrXtgZ0hV4d2oJJ1cRVgiqPCWX3PV82Xu3j7Vihqg3l978occ9H2scPHPv7eBpm0///
dfYH+FF6P9uarkHDUWo0IFk0ThbrifcvGEnH1r6oWiLrEYf3JA+CjAFOs0QLU+zKfucSlUoLuZYJ
3GURLzL6X9+fGznBNJ2wt7vVw+9Z/wU/PivFzFc6R27Au42ZC8DrqZo3XlGqeax+xIzItHGfYlZJ
MuLmTAcV9dBxj7bJOXeVHGnn7MCiPq7eEPK06C78oaNXWy6tBkBN1SfK5o8F1kJyQ/Unmpf+/ciY
u1YRiIx1KgA4rgIbxSXnP3XEGBypzrtsQLo4el6/m9QxUERX1X730zbxGkFHz713O92e39PXy2s4
0WFRNA8IMuFGZLGFYhHw/2qqemFwVpc6BwBRjMzCYe5MSxEj49+9YaMaaGP1pmXOXoMxZ3Vqdq6J
2C1tnmUu08DUY2M1bKo3HL/qTcY9DaThTfYhYnn1u839EqlN2U4hy7MgadTS6QiiLrpp/uyATA2s
pSDUjI7beyI1WvKIrCwLaFb8148pSqBPSYUF3KtfW4Hlk5SIpG3G+8FqLYnUtYD6W05myk9ta94l
k5gow21bdaYy9CJghw5Lz6usrqDaRB7tosJavGqmskXAQ+Xv4rJ8quyG0t79kP2iRlrbh2GTmNP8
YXfdieTxS4rEY1WA18F8gm3eVcHFSLQI/iUPIKMm9YvGiQlr0r8s31lHtLCcn9xoQRzIjR6aL0kx
rYMGLiFGaeh5eUJtpTadJvUdg2lkfbOJjUpmJxpJ6Q+mPFsblDmDQF6N8V9qnmTwEQkCyLB1Jkap
2mExyMy6bjEwunaOmPry0dTE44JBpXIXj717p4ruwSEcL+DDTiMH+dg9K9hYsHyWGT6RZg2ERhpl
Jk0JUVMfE61xbQPHA1PkXfYOkscFWLSh2E3vMq+qI4LmuV0libOEUdMLzDfCZx61P3NzcO0D8nwA
TJ12M/QpIWqtu+LfkJYc9asAVFUg2yBHgqSvsG+8shxSHU+/RsQ0DuRC4h6UldXx7PTUK3hMCf1k
WWGwxG7U6u2GvTphQFhXVbS2bpp0ZnkeDvEv+QCBq++7uRNzkji9JV0OHH4YhOE8ZRYfAA4zqg+a
GTNaUwDFxnTDbtNE0LRAayoEtlz30kZNAo96PC/xE+SsN1eKqntpgzLNBHy1quoVdyJpDAt5vyRS
F/W7DXyJMQphWIfDE7PIqCxOkp3E8qkWQrcqhyQ+UpAIhxWAtUILPZahbCBllN2wN/4aWYRqA693
NJRF4WTQWUS8rs05ZjEU+wwW7BWn+oSffi4PW3lrghA8Dcd4WMxgEOjogxmKv9/8w0VbgnyclQ89
fDOqxkQpSa4UVUiMFYPIOuPhI2Hl3ArIAnsMjxRwakZv3dDmLCuDtcc2iINdQsFsKLA5dZdYS72H
V0duntNr2fLIhbI6s6TQtjMiKycieXMLDd45yr00elG7Yfg4LTiRjY1qBFXMQ+PDAOKB7O2mk5Mj
7I8pTOYL4uWjtNtKx/NwHd9d3iGpdTAslge/DKvigG2z+DgMk0Nr0Ct2WOtPW8j2hiOcFS9w2ZbI
kbo0ndccLjy/tZqTBAkg84Llo+I2GoAA4vtXR1ElPrBEf79Xrfye0+LWGyRd9GOlgJvSXvfiJuPF
lGYHYnmPnnJys5rZjcz0nEVNqwYvtJ8APamq7C4XEeInqfX/Dx91J3BYTdvHtHXoBUVzT9hM7EKN
b+Rv7B58WTjFUDH2/5/9BcOzvb3Mi50WIYM32xgrqpU6E73X+VqhqU2mhv0bTV9qW6rHAfi4SOOe
XyO0SaX+8Yc/0RF0B2SIuFiPDi9RrDB9vab3l/OF0KEkC2HDDb2ANfqfObPDwu2EXV0f4Hhb1VeL
gXu2x7nKFpVSjFqIEtxsx/bq/2G3NSDbIagxwPFZO2vwsP82Gfamy+7ESZxTcZlMOmIenRN/+7vh
6HrzvsgLTQMjzGVtEqPIXt3CmRckai65GoDCmnP9zKU3MKciFP52DYpuSjtudDoZv8RtIyj9qRQ4
d1XZh0h7826GkPSoOZbkeRd7Ce7lWy0lE4bhwJFGo6teL2nbWsTngboyZobUITTNuplu1e2xxusH
c6gjBk975aXpqx2WCY/0Gy+ywu9oE1GLBOXvvwrbc36yECN5bj5M21xq92EjYqJ6X5C4KHt+y6SR
NBTFVDWDWiHf53g/hUYYbHdie2HDZ6BQ6LaxAGQRneIhQd+hH61GD5T80GkZ4QpLNpqKwc6ni6yZ
ACoClCMqD0NY5rYFlRqJ1v/34JT8qaBKZ0cHvRmPOBGwXeDqAb6DcT2SPEbZxPwnzyRflt4n0L4u
+VRBLgwTa9PCOjwx8UUfs2Szaf18zxU5BPyXN3Pr1N5RrTiJkLZE9ydZAxDOvUJtb08c5sOkZiPA
OUigQwrZigNB4IEO/CHz6hLB+neIDw+eBcXz7mUjNcrUyc4j39nE0vmI0lQprqjpujboTnPMkqyW
0nKrgMf+IC8CzJvEn8YSK3KD9dbk03+swtL1/SGYGChTfL5NOI4iUDhjMwk4BVjP/qczcyaJXhwY
PLPHc+JIc5M1Br6DqjO0K9z2XMCVMmAnrZdm//GqEIeAVVayY4J3dGmIMFwNGQwWqSUy8G2F5x06
270QwO3G2kPDleZub0J8kc0IT1rauLkRhIUo1Pq6FaKxdc9elXbX8KZ7SFvoUVBVZdbcusM9WZK+
mMttRdamcMPSzaR1q9ApL1agDandq0hOVvfrTB78QJWtmzef1T8lj1ptCXPGjLy40Pp7b4bYp+2l
1tHc5HbQLecQu8a1UH5RVsIGiH1w6brPy7tNcNzddWT6yWqiIvO/ZI6S6SD5VikNUd5pp9mNHsez
7O+JrzdtiCrRgjhpRbo9KVf5s4acVryGhQAVFWlBhn0HdLrxaaTwdAq44X5VnXDkA4LZAB+a8x7V
y7QIjhTi05sMut+WRqAFw5828mWfEYbWlZa4frs5YNQP+I3sEeK2vGA7xJ4ZKr6TV0/vQsYZrvRt
1ZKVT3i4gQrJbaLOOv0nts8GKwhzSXVa0RwM9ByVC39NKKAqzLOXaBnQhcd2ud4K0rxNw0mnW939
ww+qu+bUFW2nk2tk9Tgk00zd22XZKy1f/2NGUWJ52ot7BZ0wV9vfnTv8+RLW/9B0kiZsixSF+GQZ
LwHyGiguj/TVLrnB/xROla4IyN8B6xMlxa1Hwzz5Zd42OPlwQB+WtxOUIX5ung4wyJNXqO+WPiJC
AZKM9CqcHDgPJ2qE3xOFGCgElFbmVUQQPhal2xXWLzdeGrDF4Eclrm7IoaA3xX5hNN/Wrm0+YSmH
eNY35Wwl29ox0DDqNvyi/H9atj4OCJitfQqlfwYn5sEJTY46CQw+7lzxo66hWDzn92QQsgdCJwhz
yrRIny4SBX8Errt+0xYRNHgd1mc0lCrB5f2TPJw2SIUpJSZZ6dYBdGAyLVEuB0MmqYa5pAGZNItR
hfy6scjCxXB+yzFfhhebJDFyrcT0XCM14BRDr9zGuz9XhN03fEU0ahWQHun4Gjoai2BcKWyuSE9V
WBTEbAmT1K4nPgoxfHREqRSzqzONZdvzUQkOa75viypJJkrvDCPKQBXjaYH3hOrOuyyxJu91rIBB
iS+ObFZ+H3wU6SBUwjxAAGD1gTB59VGQf4am6b+qrIA8N8PRGyhn/HtlEEGIMEsg1LynUBdRk0KM
4Ng/dY6kugarblt1kKEaTsTKjA50eCfu3N4KE7iCmt70QC2UDMnBU2Hw7PqK7/l2VPK24h6Jtmjo
+gm3OWWKMnldggqeQ//KX+HP6DOJSAbAEoIg6CmF+uTbwLHIBeKeCuZ88JQslw6CpdRObZEwtr4T
oYGU65u0oAKWbTEVGI4ONq8wNeqYjTlES977/j7svVFBUNG+qZhsFlEtNLfxZmxuC3VC2TUlMyqf
T/QDdSklE0HHmk9I1uKZgBAwuI+QjfJjHhEBymAFnWgk3mqeH0GL9oVEjxTfXBm9z7eFM6asGDzj
SHapy6NhAdKtMvwAZ0zaZInm7Vx1SD3P4diS5CYlWeedPGwcc+GtDn+uffegoD4R4NSW0BdzWRY6
P3eGRi53iAzxDBPZkgn1D4jktutiqzuRvfYPTlQLsaodrn88eVg6BkpVe9NDGWeGqlxeyjErd2qm
ZuWJ/CE7MKuKzLszyHCzsYN+TS7jSn10aUTcFrAGeohPoczlyDaApEZIdOZ7h4aAiiFtHZqiq/FK
kNzQY5z8m0eNTU4zR87lDlQWx+CJdKjIC2NX6tWOnXXi1D0B/m6H0eVXBd3FEO9jp8BxlgOEbLto
MEMyNRpUo+IMkSTb/Z6F6JsHY0o8TC2CiZslHraJePQ6tzQh+6xFO71bAceDFSQvih9XtaezXZ21
DxrKkbud7cf59dGD6j4bKdDdlCzVPAM98eAcYZHxaHDouTqmx8M6WB8AM6U7aEOge/8eSMW9d7dV
jNhZmWn6rPbT0agnRBCtYRboveQ5OSnObTynx/KYczAF+h5Y9zDhm5AhyFruzKHVFDipJGNBe+ms
ZTsIHJG48EavZa6FPRgE8+STKgSq1qkTxfMV0KFDJpzvD36yaT2m/9Kbr3tPxrfTaYhvlAoCpcVX
prNkUVQsW+DkvvppyQR7pjHz3YBx2RUG8JVueNK20kgszZn2H2s0QDExhLIGFRMJKruLr9VDbN9T
J9lFVrQK0qejsegXgtlxBkfnXAhh8K1KeYpF6HGvEy/Nt/Tpy681/VHoAUdnP4lJa/riqVoHY85F
ft8kh2oGEPaFzsZxdj/dESAGvNRGXqPnnjCzKgtUddfZHtBWEhxpLZct3A9ASLL2q1o3Vqd2yAHO
dgRkrsnX6TDXQ4WJedj2ERe5tpRlcAdmEqkoLEgtRWbeZWFHJw7mzx7B2lteoEBWLKfFuKpWJkdw
jheq+DMnYkOf+Tmkj63kW9M1461oIWWIXkpTE3+sNFbWuUMQHJCDeA4cVWoMYyzVwzlvKkb+NriH
ERT4HDG3eGtMYewM9CogVTGhUJaXs+xncRCD6pVjMW2aAp5A90JKOVQj7qAdyli/orSZKc/k2aaI
i5jgpHcK3xo0eIXbxtAmClzmxWS5x/I4gimU5cVQRWlplsXLhjRTn8+n9L6q1vlCLz+O2Y/DzvrE
tdwVrQEPDbIyPJg9utSha5YXLqVTukJi7fQhr6OHMOK2VX/VCM06ZIYaMyAtyNfLi5IXhYbwyYl6
D/skQPVQjAFgWjzCRBZvOSBA2Tns6G+kIhQJgxTT8CfHuTW5/xPVyHNzmJc74O+jEqZxP9chXfBM
gaA6uKRnimHHcMwrUOZrMvDEq1KH6hXEfkciTUej9AkfCouPjsC2gvUDnKa+I+ee0XgVK07RMp+L
2HxTE8JePm7PkPeLzrKpVS33ZMSgYvcdTTdUR+GgI0GCbg6csPwmlzmkJNVJi725BOqpSFEmTOCr
W30nqP9nqy+iPQ1qxX1B5CL83EfAZBGtIm9sTtv0Cdlz4GBEtheMOGKVQe1u281wrDRfc2o3KGkm
oSUkDNN+o2dwXDVvjUYQoljlkBtdgUnJjL60wr8lgMvAQ9tlIKP/JLiiwcvTs8W1w2fOOUeN8pqI
nsNWdVDvaozy8jwufL24ZiSBAxTj6UdPK+STYXz18sYDUnS+DEp81IBdLpM8wtF1MGhLaQn7j5Wy
RiqLP+7egwW9aVKdZb6LOzf4sDdHykrKWrP+ge5i91jztR66GC9K4EqPyY0ZMdKwAdelKeGu9aIa
jAlCYV0j2jjLJh4D1TBO7hM625uvBlv0mSuYnfHnGQspdElIxQJw7ylfExz/CB3GM5Sd2i6Cu32m
bWmJ6GDrySc9cFU0NuPI8b9P9w/Qa7kXzjjL6usET8M+oPWhJwNBgX9l7bxKM2cXBDHeCwVrUlMi
QuGYvYjTr0BsQ9agxGwdd1ffwBBpJ9N7nA9T+yeurZXF93BfQQTRAMTxNVedrGdWV49pRRJSnmKX
2/PBaxi1ROsCbNEk+r1zYqf3XIX632hujoyfK01Qo/xCywNDzY1HCYjfuQtePe5kxfEwI5MzZNyO
5snNVripfP5QPGvBYBK+PAFyKFakFtGUr56Y0NGmqEnJNFCPsduYnLgzMh4PNO2cmleipqMHvDw5
1jglahToSDwcjdE2sU3+A5cbxXTb7iw5a/7/tRDsL1Vx+ZPNGBJP7QZ7qIiVRw54Hf7nHY7HX+Qh
iZmNdKHEPlmyqsSJjsHP+a+vsn4GzVedBrV4TynesMZJCOQ4cQ5uMO0T5ClFg7+2x/Hg46/r4G6V
RIwKrbM3AbR+ZsJRB21TurGuX9xcjp7nWYx7QIlygVfNFMh8R7U2CDCiiX4El7Myis2LdY5alnOf
lkBbTGw2s1RVd/dJLJDiEELmpO8KI5GieGVJGq/XaM4L1vOa7CThFd7sqXTGSpdF3sQEJ3VMW1r0
XQRg+QNHleOAw3pbA8EQ2QRNumdZJxjoEQEBwXX9Iib2sfnX8oSzEIqg4GHA0b7GH25PqxaaCVEI
J3RGmAFOION3qblxzI0T50FFO3nXHEiPtchvGMKo4txjmygPZ//YyncuGUbi0XafL+XwDir07cSa
0IKY7q6oawBW4mPd4/CG/XX3/70ucAV2gzuu+JvXhAtmmGu7u5GyzVDJRaGoo05SfbJD3F491jA3
5BG/K+2PuouXXc/CoZSAh2KJHZ5rDNOUt2/2HzQoAusfey1PHaiITgg2hkEeqbvU7tXcvn6MYA15
s5Aqx5MHeREbX8iykNxASzfw3E+2sUY8JxkpkkK8X2slEIkiouxOxaC5HKmPtQwop9vKNUfMDayN
qd9vxhPXI0tK4C7jEvUBHLltUph+DbiW6NDOcn5yvatFCzAmQhP8gbkfjrBoBHyz15hV3fvbAlkU
HzP+pkW7w2Bc3va1d7BE8GX0IaaJmjvMosWakxQOJyIfEjYVNjwkwveH2VN0cIvG0QRbZFFU8BuT
GbilQWcMqLtG8rY9AqLQw6pS2g9m9jXRGkzreukXieW9XC3cRNwBLa8d3Jk1sOch1UtwbTD57RYE
Sxw4FHTP/flAjWUxBBjEFwFR2NadMcW6mbRbrq+48YLb/HO6lf8lDarh5UHrh+PvnISsm3fGlCrE
NrwlGD1/Hmx+eY53YTkEk99nILdFJEBf4rpIlBl+BzsKf+k9gr38+jF14j4OP/YiEZgs7EkkRGLs
hJYEqJnzuQ2NBERivy7GC63M0R+vJvJRXqnp5pQ4lfNNufYwhCFS412pyLp8bFLGGQMcuTRk06lp
lihdxSeTvSPwJO/hyLMxbWafDRH2aGehx6ePVifMaC/bb7c2zUzlCMop0Q4WHrqFgBLNqhDF/PS4
AYeGXUu+AIi9FEL/rP+vulTFWi09dJuIlmHqZ14dy9Uw8WjhaalSXFYPtD6srsrjFm2MnKwugvzF
d9zVNw78yDq5GE/hn0i37B5rE/C0bDoJHaplLCtNnYLU2W4JtBbk+uvju+13qmWaOvOIiejIhFm5
KCV/jRIgbPX0vt0FvxIJfxkFLVlv06aJMbA8d44ZPthEhVlY4hsIs1C1/ASU/ZByyCNQm4Tj8Fg5
bln63hFIr+r+yFvGRIMZkMKFHoNqjjAu08iBBZLHj/KWkPDsvfAgSWKf2k/N7uCHhWNQuZcjoPYJ
ykNS2ANmjaM1a1ixRoYUNvCGYT2kfsHNGthCktGCtTOtzbmfRGp3wzKk582KfgBvJOBhi6jQyzGW
OT4qUPaI3x0PeAE8cJgW5p63G75U1BAm8Y3L55INv8vLwiW8vLQ7Stq9h4wOx1mcEZBz15BI4YA3
UYb48Dqlm5FfMNPBwias+MvH7gcQcCHW/ODOuQREDWecS5yxmih5TQWLyMwezdaDnco+EsY6k1Me
wHGPdJSyrYZQxF6GEVt29/irI+TwvnTv5j4naK938efH2mg4GMs/Tox+pwd2slBn8AhUXfEqQQli
rJUqdSIcw6lD6hxzLWmp+OJm+dlTLRItdfPUFzPCLb5Z2mwHtEGWEAQgdz/BEMufxnFZVQF4V7Fd
2T1f0fbSBZhd/sU+lImbTBT3XXx325zGWFNRckO3muyspGsvg8YB/TTDIMYKPw1QB6uoROqyrEW4
wb3X3XXpcuWQeVqqoh6mH0DiTOc9dhpW0aSOCLbY+VqmeOBqmmUtfxo+x4IFfFr+gl/+qEti9Lqf
DSH7tFTQ+VkMstHVnBBjxQfQjbnQgw4PqlW+m5yB+HTcgcpGS/YBmEPuqZVm5NPBudmL+6ur5goD
ygGDgY8N8HeI0IFHENd/kWd4FXZgziSiO47K9IalcUve86QnCeqqT+fDV3yI6kFusuAcL3mTyi39
xDK1ORqGmK/8Gm0rkWL3R+QSLUxOGbmS0PlV1POpfyj3igJioL5A8GIdOLogI9s9mz7Pr3ZXTUQA
WYjd7ibd2bfdXAccRpv1z5VLDGP67Z/Iv7GHOlKrbZ6aTe2hqr/6OW8/5t1t8SSXcj22nisOIgSx
a9xJnmfCpPb2PcABRQN9dPoiO6hTAZvVX7fCecaDR6/FEpcLVFtaV/0wCdOYwooruSdvnoTOd/bG
reFoSlS/6LuX1R8cJvp/1DGj7y7WATZBHSenbpLA0XGBSmECWRZkgnakmDcNd5+SffUxwMyvLxyp
KPu/EkA9Mohc58mSh88DDX4Ohrs9LhiUvaiBuJUOjkK4EKejHM03D8dj5+uLsNi503umgziSFlzS
86pM1hBOQmbQeuVF5H4FZZi+fz/A4D+ESU185Z+DRaTgr1wthOKjilLC4TTAltHYW7yNoXA3tlkd
Or6oHO8ayZh6iAPFsXxHHusSso+dB33YxKnt9GW4qclpGr8YLWxTCYZ2YWJrjm0N124IVRPtnw8l
a3xmLxHYpks6wW/gW3ak52GAtPzyUNZr270U/dCT7h0EDdZ/4NQYE8bPx+tgIsr5wOqplUbRcEGV
q3nTvIXUMdx0bqMQIM6/Gd41idvXqLF+/NXFobV1B/45Tdd4ETqfHsofQ8cZgMNf26TYaw7+NAkj
O7vRWD7HR2DlB459pEYVcEw/a+M6bYu3SllYVqIrfye7ByjTVFpEZX+4XNixUVaJV3dqAwb5mkEm
0dgbA2pJg80rrELVM68PpmG3Pp8I/8V0D8/Xifck+93pMb6H5tsxj4qT2U30m5DfLOMc644Awls1
MYmy7kySEi0qlo3wuynkZb/o7YZ09dbFtwVV3V0IDldqOToa29kQFoDyD/aB4c80xq0DrqGc/9UT
w081nj58fuv8ZFbySXaUYyHNNkJmQQRbLR+dJt09wKYZvSOJmkLeV3qnON182rp9e6TR61+Aah2S
la7fxUgnjd4oH7k1YNakBWdrEzMIIkY3bVxDghW42pyp1/mRNqkSfbVhvTBCaodm0Ls1KcOy9oAS
mjnC3gGs9jBzOIFNl3LTd97Bqxp7sZgLYooXiZYgMt9HdLa4IYW/pfF7MdIEIKvFBOs9Ru4OImHR
bKyS0tSQ54UJjaRGTdXGrlCWFZU8Uh1SrR0o1AzoS0LstpqHUW9faGy+lI8KbPr9DEZcp7uTxRV4
pWLUgAaynBhVNMVySzgONSx85Z9g+aakUk3TvbNyz6RFLZrXZtFU0AkAqAT7j1+PcdFHVZf0t1uK
MvLNmb4Tf8mbZBBhhgnTpkcgvX7sBXH+e2w7uIQMunn8z4LZZ4FT/3DtiWqFWAl+RqZn1BM0fBao
YgcDAuDAPMExkTS1iRdS2t4eQnOYL9QIFqaLzSjaLTx6CQPZZM4Fh3NlfP9G4ix5O/h65vEWefVe
Sw537iJLel9SFx8R89sLIn8Uhh8ezbEyM1h0+WjD5wmG6KKzxaQdSFq4G5Ug6ReTQGA0Wzc6HDPM
ZvCewTVm8AnnIr9J0gISS/akhsotfvg4B2kkxT/5U5tvuySt7UJTH/rQ46SaRP0kPRjKS+3i/UtH
vvL20wFSHkR9fJuATHEN7SezAwFWA6g/jZq2YbzevVkSOxucGyTJr0QEJjhJQpNwvV0NjF7gda6Z
xuCmJai5w9Zja8yhnYND8NGYLczrGC6GqX9pUl/91mPiSLFsf0BDGvUKlCocfd+H5PCs229a4z4N
X90NRGa141c870mBV8jI8J0raL3QwrLJmijymzmBaX9ESBZScEWdBNd99o8NgK+wGwfxasavnPd9
9x2TC6y/B4vPRUhkdDmNPsPtJUPfDUxWVS9xIAHmDIueLfgBR7LXOWEK8reoUFeBs7Z7KlzduInN
fG8Pc0GEQCKL16fWxfqWi2mw9//VjtG3oXoS3AeyPT75saz8L3SlFiw8EZ+06Yaio3/t42AstWr7
dZCzAYGMRbxNi0SlR3S51oJnyghboGnRZ4SYcVGSV4tl9UP0F552wGadKCsZuWq06a9g+xzPS0hN
jKHgiQYqQxI5jYBN7G0o/LrQ/M05158p7AdDFeTDhQNPK8p2Kqd3uAUluqx/6rzQ2uP9qqlf+a8L
+/nYeyPQwNQEbJmM2iN5SzT5c7UpCl+PRUr+OgSUBtT0Gq6dgL1+M/rnOCTP5Wg4iCB8f6cTGCJF
Btyf94Y6eE2zBX14+2Z8HzlLVrXEYcvNYvb0EqAxxOPdCoX1ibLUvHaNt4XrYxfpvW+uLht+iIfi
Y9nn4OuIcM/0TWgZX6DJHW9VFC3rRotO0paP8QD5hO8Cc2m45qSMEhFJ1ci+NipJZMTicUenRTJo
qJfqXj+iNAyv0+p9Av6Yr5s1jhjE48LDAYKHvDTICvk98T0n0n1yrfCMmugtWrEXsuNtHcsLudt8
zgyP+DpMdhHuQ+Dx5DyUewDKWFUmaz4Qavbyk0CAGToutj4I8A0ztCPRbZ5Q0fZ59qUaN02axXsz
nP2/8C1GdNMXgK4hElcHb/E0bw6pzr1+xFJXRXYRNdhFyI68c92fhVCh5zIbsFGj2OCMJLrmyb51
JmH0o6axgEXaw+2LyZIT7K/otSfDfGgTCFY4dlVIHSoyE5DAXOoD9pN0LlU2Q++Km8Z6AZV1YDpM
XOWjk7ON/Y1JLx2eAjYayO7RfZiFcyOA+DbV96BcwNBJ/w3KghxhMEMjAM7IcNLHjp0k5yPCOyB2
IypJ2qbWiInLfVNg/E8F2zlMM4M0Z/m3kK8pg4IWWwR+sxGaqu2/7StBYy0tLU/suvYwP02gtVmj
2P/fzN48/sLi2AoqcQMOh8VDeqYe8eLWcGa+3a4gah36tZkcEAjbnF7ARSqPzplP52+igYBQrecb
JHOzgVQumscDXPZH7bKxiyY2G0DArTXK3V9gYJSgrfsHJuUlH1NwbRQxYeIkUwoAmibwrARQpHC6
Dm2pumow3A+kZhpabUkhGxsvndktw2tfG5MTxfNswRnjP3twDiKwVKb/lcDasC5KVI6wrmTOrzKR
41Rf3pmOx4xzKyH5YBs3zpGcv8xjt/SbcVbPbb3Q8rdUWDdYqnl6utT7AF+qWMN/X2ffT33wFbOr
kA5PLs2/oQp+TiEnr4GADnIxvkEsvTJpxciTJzez93pRe7ykxGH091paqqBGZFDsyBpLI82RJigv
JRCIZS76SacJA/YckRcQ7kA5X1h5jW0JDkZ6eXWOVwEbYurwqskVfsYeu10nvyqxatLNe8P13GQr
xF1b2DcEIOkYo7beKxbPUvLNcWAD9sb6WbbAPAfL1QpD8RWFEH7w9VLmfZbECcSNvl8ES/8GFXLS
+ngD3OkMaASybeRmA/E6PaV3jWaxxNRHhjAKOzPGZk6fBiogPt/OMgu7e9dJcv03qDPssQZ1NXAg
ODmxlSfkGCBwTKIk/1Vea2EE+IUBoCu9RFZ/hEXkzLz2IQYy5jDPe2C++fNbAMENYRJ0HK6r5v74
4uyLrJoBrGMBCf9ZCLIDtP2x0H5QqZ7FDhsvIcgdMYg/o4UlWmWlU7NXi31/VyckGkYiBsnb1OmB
CZ9Kb7n4OaVxuOd7u4VmCtrY5SK0LQqhGjLu7AmG48vqoaaEJDU2XAxzar8P1wE37UX4u4Y60nqz
xNqWlR3JYobGdO270byHutc6UoTeSp/JOJoW+Q3tQNS5lKmkkBXeDOJgCNRSBr2pXFHXm8gK0viU
Pkl8tO9ZAwAtZ3Pe+KmxUkclF5GixuNf8j/ZAXlD43gL8/bqV9ZFwUXUKzuXyE9jqCX9PD7au50o
rkPcjEO71I+/Rc8KAYB9JRBUhybPU46ZMiz/Ggozbt21wqBK5wM/YMgQ3UYtTGZmMdERayqVjbYE
gCiBe7PTkfS2K5SsPLCPQnRoqHAv9Lmzc6Q6Ye3FxqZDNKZ6INLwLGxT/FDJf4WULg0WbZqGthwh
Wgj7apluVwBb5KVNBR+kKb49b4D3rhw50ZAxSWT7YN5TezgS2wbMPXsPVxEP885f3SNxWykqg9yq
pWXgMXP0pKyVeGYDGd0EwSCqwsXILAyYL+pJpw4mvpITY8bAW6JafTCKq19cIppTXn4WygeXJevM
nMPDo+GBJUjXC2mTWyCo6MiNBYDgTKKB9C/5U9oxh7QHH/q/88vq4s/U6h8pSr34VztfX1waU9kr
fUZyMRZa0smVp6O3wLGGpXbV88AANDsG6/UA/0w4MbhrUh3X099huYxythd6zuodU28IDFJMGRd3
BzKsuwoiH3ZqnVJ5QA/mpVK28PuFdLeu6wEl6ifed0hLj3rXrbYZYKO/TEItVkysHKKFQPmndhWE
1BNpVHTJIDmnSSWIiFXjcOV+anF2qIFpLeC/KNrh5jKGzhgpAco+/BHh/F8hCd4AjQkeyKm2Bg+d
rwMgieq1XV5vg5x+01trguP6fb5GIv+5EbtELl0SAd5B7aPGPdG9qHQuj0ZACp4dsTg304jiuLQ8
0oGCizm/qd8QSlgpFPPnedb1vHzwxjCLVQ5lRjHqSpS0nnbnH3li6IrLJmPaje1D+7GOwdi9uJ1F
2pj7ioZP5Wh6cGkpkPJYx4cN6phLAm3J6UdbxKDcMSS9CFQ4QGZzrcmsdqexl8fC6VOLtfqOQSEB
GWzjPupyxVgfuhPKNh6tf4GZ80SnQrtARIjjGwpzYgkh1TnjBhpqPfVJzbjYXZEXh+MpnDeJPUQZ
Ud3VCSPvfTHOIilDAEl1BezDbq0vI/+cRzXW7nAfVZw9rQ461pHQHeBpC8TlQkgtklRj7Zz8lMXB
zjO0ZoF8bdf5dtvk2XmVOqyos5eGsY73+vyyajDILQkeQy0lRE5782AfpdB7BGYbFqK1rAMVc/GE
4NstyxtlHobGcQHYTavOnCUr6sAedxolDoD/gYER53zuGOTH4LSi5kV+KqIu6MK20rv4KIy2WVsX
yO4taIyPKgTQ94xwm2ePASRH9KbDIPFKk4q75sfaVv5GeOSpcf3qqbJ8gm2YFmL1x6VNx1gEY7Cr
GeGhacCryHl/I8NgEn7vZLoCZqdsEydb8PyWmf3qMIcCJJm2IFj7QOB9gUdLFaMaM+Q/r+Y8Yq3g
Zh92Z8saKgPamj4ZT8I4T4bhpwLxpjgI2k9yuLCsG1yf71kDBGgYUwqQcHso54I0+eeo9UL5w3FL
pojxZwOu+P4OfOAaE2JjJPaw8Z2JBqQrgVehlznP3iiqvIeewBd8tFCHNoPVaOcUVd7Pe3/27aKV
nPXz/TrKU4luv1984nYx9mSS8QpEHUuFoCwhdAWpMdR3LlRATvpJRnrzj69Mf6MeNoxtRrJEKCX6
n7gUj3RRsgA9gsZ6X70LoG6IHFlJWtie/eNHoW6dKCy9NPGfeyDaq7Q4rycTQUUUE4DSX6CdRc6v
RLc01XRSjYKmzDDiqsQ+PK/qHBchCg3rKwnAI1RMOdXcY3oWIJ5OZJYTUWdzrtziHSc4Ed7P6zS0
wQMZNyHr2GkAmA7icptW0RsUe+LuAyw9N9J8GlHMiFIGMzVDhlsn3JeoqDwdZlKr+UN8626dBeho
uVW0dAcnrGzfcPcmcC1UUKbkidhTDEDkhgwD/lczBNd5CPCW7diRptZOwLQtvj1U0fx/O9aOhdPo
qYWzsIMBf1Wo4T3WOTVb5vYx9Tvubw7pRDFbVVm09rDho9lz2KmQWi9HC+nPZ0qs8rHQ6F1lVu1+
Lqd/BFpHZDLeLhiNOOnvJUDpTsUbQIzfaGTfjh189Enz44Bd3ju0VNCFwLbPBCz6BgT3YPvm0VR4
MdUuga3tG1ytdD0+XgKwAJrSQ+EaAhQsxVKBUoIzX6S0LyNSwopIsTEuu7jsf4cyhyAroZNGDt7+
XwXEhFKZM6hNmfWZEw3C5/u20zt6jcqwQxSuwUT1eNTyd00KZ03fZHYcPZvhC/0eZoGySdU6Jey5
Wgb6lFvQYUNz0aomZk6dpnw5PHtEQgnDgkkm+2sS/6b3xZiXtUGbIGtSLDn3K3nUmB7lK00qAiU0
OEsa8eSlz2KMIAQOCI4kHo/Z1LSmREjaoQBT8t468CgJ6u8oI/s7x5jr2CoQqx5nF9e+z5u5Q07f
xUY2oHcuqWJ3mLTxuOQx+6ZnxY2PlPVgJbADGMnApXS0gK9j8SHfYL3DgF83t8HwK6uMlOQeHPCc
lDWWvIVCIc0FK0gMByHpgf51GudD/htYQCL2qi0dV1CeKombXqys+YOamcIknjMR3hnKtYMzRE6I
1UOamghEmtaUwg+8dg9cK2aDSGURXoFysaB1rsIJB6hD6pjf4hSx5cqD3PxICD7FdPpv4WATk/VQ
jOMUuz6AoGmq3/I72gC3RmKahmp0tUC39U/5ukJC5pMFy3luVlVmqAVZovXTXByB/WLJ2jLZAzi5
TdAoIYuZsFWizsIsye7x6dLjDstkUNmGkyOGg5/5nseFL+ns231mhcTcTV7qmcGAbR/irwe72FtJ
3SWFexIt3b6SPS8puWH9vWcmrKH4l2H7zHRKlTQITBrCmC6uLU/zcC+PN3/wNBsrdONSXKLawIQE
OcB4C3b76Aa00pX5LlynwJeGKj15+4GnasHU2Qfa6KuBB8FusaUy3PomzqGqJ3/YhqahyaGX0i7A
U5jM0cX/GCqKj4T7pGm3w8fbck1pfnjvfp5ZJOt2gj4lOqPSQuh6Kl7oNrXoSY+H5k6mzrmGh2gR
T6zMJVk5XcE5uY56iyx87FEbsQtYXLG+qvte2+DnXUFaEYG3C08xyh+U8uq0O+MJ1LBoZxguxsnt
pYQUWgJj1GgxG6dHTZydrBkvpFz9wQLPqyAO7SJybTSUWlhoCrrwkkjTlN0qf5nSkzyJ/smJWrpZ
TW/qSDIITB5rVcVgWo+trNYz7k4DSFw0DcmUlL1vo4oOd0wMSxgptxi63ZxwJC4h+rOiLZWxblsG
uMqAilQeEYzgnV61TnySzyl1Tux3IzM34FxfGzN0f5WQ+PGFPGQC/I/WHPpigd7RuTHtCOtBIgrt
s3CbcbdEnxpgj4FCwwl4j7lVXzk8FBa5tmhInkRrdmHCcXaB9sIm5Yu8Q9jh69FFJAnJfPypee5B
BFbQ4tw3A9Nd3OIz8k87h86q6CJafNMQFYthfOHQ2BZKdfi/LhLOc8UwAkdOHc2IuNT0n42uS2Mi
4WjogeZ7tpAHilI9tJCAY5+X8ZNRY8bSmT8EhDxvMw3HPR1zKDZSCBjysIeWyp2Fi7j4u2MlHj3V
LwfJ19jOF9V0Azwh+e1NSVXwZ/NvfTCAuW8psz/N+Jqxf9wAenBsSNR1U0CqsGF82R9Ix5pPyEYr
KiHAZFznkvBDYxxrijRs6pJGyZiXPajpFqjuvTq9GS8ST34IuBPMgYK4/bM6JC5QIL/IR+3UpvMo
BdhWfGbdYR0vJH04+8TiMPuYyX/zEF5P713CCJNau8tBvfFPnq66HtBE8Dr8EuQr7boLLqCKndYZ
ZwO1DQ5o+Izr0gm2aiXGKpyuu4EJo3N+YPT0ApBvu9BoX8yLFl0yLH8/wy1mxPtNxRgu6merKEXc
Oy4/KN/hfeBi30jgXaEESjaEnzkGsiYd/ESif+qpL0gVGGcFlpTxcNkPgbdYdR3e7K9ExmsQMtc/
4a+4M2/kKFnYfIEl/Nr+Nlb9w+ujtimYdls4jl5N9F71g4Xt4kvv5hhFyApbdHeF9JnIcUQgu3u1
X/dwmuV5xYpP/LQoDdWMKVJbnLUDW6lAJe6hUkztLX+neg08QFrQO0lfxKdPqQyMUT3lK4UzLMxl
m9VIMs42V+WGav8e3s1A1HoOqTpQs8zNFzfNJsmvZ9UiMgNjibKobjF+nxqh0ZywbKlhV4KD/YnX
3NQtvBdnssr9ak512AtIunH4xa8VIvfN7QSPIT/5Ob6YaUoY7KyyZ1j4yLyHl0sqG12NujbnWB6r
RxBPafdulMATdpCWwWMnlLrz1Ee116llHqhsHgWljSrPfmOCIid/OiDkDZ0AqR8hgsSdqQBcVyOh
AcPkPvzriNxPo8XpTgx6n1+EcaN85b87TgRr2OgpCJic+nzW+CK9WGnR2fHOSkcIqPuvNEcF0tso
3oCpkxpwx7fPGde1ITzg3xmxi6MCQGMdfBD1FqI4rTw0eTQOFbhEo7C2DTIhB6CIpH7m0xEsFAWv
tdwSABohKzpeU8YGE2CwuQ3okzXinfOwKBnFyi+BAgVU2GMgKwuplLf/Z5IbvO6uwFOIjAH72pVD
Bif81x7J/Xki5Uuo6kS9RGQDfGPQtOaO41FuVo4qJrHFhTyYFwZ9BCrehh3WQZXM0zP2NqIgZEp2
ndiotOQg0sicoCu+GXgBNsWXJ6PdDJfpUddpmUJx52bURJchSN4DYNWOQ3FRoIch4SlszhZ5tDtg
QRm58F/qlqCVr0Gbw4lhEcYo/kCx6uDV9U4KE/eg7RbHZjHa6vrtWUvivux+TMvFTmUEzrBeALoB
rRGDSyHlenBkpz6RTU4XeARINN6/qxjnQrR5WMlF4s6BDvwPOC6cfQYZzz5V/IaWUJpOrFNj8LBf
HgcF5yGcncHqDn+eokrAa3oT694idnRf9SwDTRFtLzVz8tt2FBP5eintrPcTn8Mi1lHe9oNHCIGY
Omszp4Q/IIvVwaMeCz/uaV17e+53LDcMgtr1J6l7gDy8PWq4xtcdX80ZysSZK0SLAK1G5bOxtER+
E9bpUhtGefeR00MsbehIMBGJM0Y2/7Q/xgZcJIJO8QfS/KIMq65D1xNJMwLneQOYvBdwsiPeanp+
SPEFXg0yUc07vh+OoRppXmDrrmQu/WagDvzXfi2XoOC8H3uab3d5qPkKZ90Z29eqNv4q8MCbE97C
KMsPac7RXBNqSk73Dftc8/7dKsVr/0/Jx8T1HQpvop2WN4mYmKnUW+Lw5Jp89ofkc4d+1AfuDAGk
UxKhG559HtA4f31DwpcP1a4PhLlcrfK5NERv46YP8E8TerFT2OkJ6ugSFgUC5c/44PlMdMTNKD00
cti0Ca4o0x4A+O1xU5lVg6EWJDMhwQ+ZmVNKvdII/F7tKKUeZrG0XFYZ4J7RaejRGZLzreHOjLnm
9Du5kwBo4ggEJ1BRlsW0ceRLdezopklWTeIRSS6ZMGkCEHVDoMyJ3+17Op92TDuDe7RkUkC7hhI9
Bl7EYRxyhUWmaY3d31ZGbxNcErH9SMj0PgRmFefByOWlBNKYQ4g9/95dsnKM2yPa9yITF9odgiDi
Ko63vcPKtGRKw1zCUG4ASOhw57HVD/902RtsBpcl6BxrYFvxfmuu6jgatA/FqYbYvj3X+DtThU7G
q2vE4fLTUmMJ1+sxbBf6i82CWFHDZomTom65DD57EeF4+tBc0/7I3kzBJMH6OPkGniF/seaPmUcy
tRna04SRdfIqJTL5qNmUNhDU8MXFc9bIQZ7azTPQ6CKXKYye+Fj0Cpez9zK/Gz6OSwPFIDuQkspZ
VK3Yb1UyxCvLIZoN16HCWb9AsgW23ycvardURqSmw3o1wpa/fVDeOeiq2IPqYICzKeBW8RTw4Y6c
JMRdrDV0anbHPJ3mnbLlnXFXFIfyN4MOoDAs7CrnnXWLn6VfvSCOyymba687LAijFTguJ50WZiLl
pBO2UmMG05P+16tOpTSACU5Xo0ZEMSLUHelEuy3YHkFtBUyH3K41oyNSz7t+CtVrkirmro4/IDKJ
a34elpd0dG9tnJpQa7GyMNmKAFmV0EftU9K3fM8nbr+YZT1srEMhN4DriPG0p/WbBfu9grYvwF4p
QSQR8lzR8VOie4eZiaZg6eki/Cv0QEw0+ZETRXHr7+C4e/55aS1XzJmBiQXJMr3D3qDHxGh5y674
M/TVYd6UHGpFe6xdDGk5u4BXXAVy3tY8zgQITkku9K7ObgXcaiW8k7EQDLJS1Iof4VftssLN1Bcp
2+RDp1wo2QjK4fYQ2OssMI7DC4w524XbSNQro72ZhVrB9JgiHWscCQqUKhCkHH/xOUbYAIL3+IB1
OcRkTzbepI0LnBDle7wska14UeVcL1A/M8ECh9Lu18y+wlFwCBfUibtOiEnf+oESrW7czfwE3Fvh
LIzGwp0lca+AwH+nrE0g2baNx1AWlSYCEhESwKpBT04gAqcxAK6nbDCk1Y0iDkXdHkaK5NHRCpIb
yNMsBbEkxMhazwL0BjYNhF83HMTtLQz9azKlw0p5iqxWtXWpSwnujG71Y98tDq8Y0JXYD+yKsNKK
2iuhHgwApQS368vYqWgtFEbhPY+zUjxttUxYZKQlVkyBbdic6cZmAtSO8Ss3+lDAVEdZXf6Yr4p3
gvKZ17hvR7KlJu+ZhDCotnTctqq5fqyTRsWddHH9htvgO/1g37ndoHiKfLrUvFzWqLGMbRlHDhQt
BNwcti2jfAz9FaBftrQG3fx2SYdwdbY6A4uyn66s9Am+ndBBt32VhEJG/wjVZ1bUO1CkZKjiQ9F8
i2RTJO5Emqj8Y/AqCOVKLmJn9/xd8qxazfr4h7OqmLfZJh/IvCOmS4OINt4/JDpp6X79jCdFkf0Z
GMWYe1SO9i9Y1oXyRmBbpCglvI9fprj0AFEWZG3q/SboZh7lJg+HM52VVInZZ3rBqMUjzOsRezue
uT+upi8sO+jgJOiEGK4ycF5cQpg5KElo0l7jqNfIUPQ9SkgJ9H1XApM4BBe8HEk29N7oM6uS1EWQ
P1YmQOawt1fEkcWPEPA/uYx1rrs48ktr9fCPMf7+WyevxbeyyGz3KPl5aiPk7pXLr5umdrL+Iy2Q
Q4RD/Xe3JoARakF72VdKUnZVmyqpixY3L1nNmSFQRIeNPd9C3Iq+3tddW3Kb1jHVdskgXlLWD0Tl
iwDAt4DcdiHAkt+gb/JVE2k+ipdI1+ej+b0RM0Gr1PjlmP4cYSLX+G+OCmuQXLnZLBrNuAZOMhOR
A1tVe5dqi3KPtjXPQ9H5l50NRba1kL6F39pYutZWd2fnCWSCpar0HzzFB4Ivb3rF97ALAqxgVnqB
V12o1HJM4fCn2kU4mjETBVJpxdD5POlakPI0T5zD88qqUmr5ZOsIMAPP1S8WPaQhR1VwZ6SomDqs
y1vafNutufXJNnCzdlugYaRwb9O10Bh13BvA6Ri+r1UkVtTuIjoF81g2ohPiM6q9G40Qc43D6gli
K3qzQkjnlhVuWweyWRTJ39p72TUdcHeVbrFhCG3kVfQnfD1pLktl8D8Fy68pEmHMLCNPOoN03WU2
tF4rUMDXs45zP/EDMssSpUtGkn2UJcJZbZgAdWQzMsDCw55dFReH6PwykVUC28hTVgVyt7vHiKOg
n4ibMmrybI+Hv4Zf4fwOSrO6SYC3+2j3CVaZ6mVaEjkZzDOCvXrKx6uDGxUdwxVH9B3Vg8y4DDEM
M+GGD8Xnqgd64/AvbcrNrB0NMMnqt75zJdFn9mfHyCotcfFYjGWh6P85N3ZBW1YAdU3rAwEKJOkH
e0DDVPfaGNCNpfTdbgA3pP1LaKf8tFLzGiS7ZDsaa47fHqGC8tHftO7l//Ausjl4kX8vVzileWQh
bZYBvGeF9r8BYhJp3LLFKVbqo7oqHxjTQf3BW1SAYEYeHARj1hjgK5+jb+CiWG7hy1sZwu1QvfOz
zykObCa/3Uqn2MwmAmdW7TqWX0fE6r0bODmHdHZ0zRTiJWMvv3SMKwWeKzfKg9xtu48etQjlt0rU
WT9Inzp7y0huCV0Hg74ET/7ZpbSKD9ZLALniBhcc7KXF6pWAGX/CTgsvWx/CofmYupr05CM5la0R
ZTN12S36usuhzsooyW1nGRTdbH8VnsbtD7WrtSboWAjqfyFMsi7vJ5AqYH/qRCZZI309N8bIxnrG
b8B9Us5SgzowGiZNrH88uXrhBNkt5HnfmumPDlZYP7Lyw60/nJTZNiS8/KQYtASd/3dQddSWs1jK
HBZt8V4WJE8zkZH64OD/yQeE837D9P3rjsRqTzG/GQJhRSkDMkDvdHaqwtgJO3DXAC6+R9k2g+4L
jpj59FuGhXAdK0/L5nOts0KrpoqR8TYd91iweY1dgqzJrn+HEjSRKFj1hbwEGCiZoxu6B99e8e8U
cWIlh2h0WjhqGulkjV/NXeKLip74VXy6zoa0VOBQgQahf9Z2DQJnMMidC1SsITvB5M3zQ0xlrp/U
qMsF9r6vfVGQ7ULS5+Z0H/mDxcthgY9AnT/pfvUnxu3qY2/NfxezCa3QIN86xSxqNmdkXSprhb9P
sioDsD0ExqBSGxMghu+YnLgFVs0XMm700ahcvZkzrGFk3NIdNZfmXmAJlpGUDv7K3G6FrPNqyyjy
3C+7dS9+40b4S+684RBcClGkZoUSB1TpGPCRqbHangSi1vS3JJ+WMLXr8+DKb59X5O5KYMKSrmZi
6YFyokWLGWVCRuFzqniCI7cxtyCF+fyyQnPUB/d5jovsKEq5gQf6RLtXpPgS8ZE8k2nFy9Q3QKP7
6EnnLzjGipEpxPcbJZASFzDPD5hTmPCRof1KDkAn2SDBDnThO9UDwJe2wFeZ9ZxurJjTH2h/bynQ
Sq4K0umkem53bJo8eOGfnqLmjCl+5SuMgLj8jSzEvVuYQrVmXEuu8r9faVYHjO6jPEzwr9Y3SZiz
wJXt7B3dZNP1Gbc8W3kyhSl/mWu/EZY/xdbihIE2CjWqQw0xZa7TmXy3TaWbKHYjuq8bqeDwvJtC
tiqwwvrA3KUXekprMwtpQvE6cGpe119GFArn/kR0DMIaTzw1PZpVM5LCgqwJq5cg55A5RuwyMUJZ
kwqgq6LNKI3nFj1cU/Gw8YHqQfa0cVcC+H7mfTWYZ8p9fZUNGpbo6qen4CoCBjNwoYhPcbvN5rAv
jD5dwkqyHaxsv+yp8R9v7YWAgM8YdvNq8Se7cvT6IVW99MXft+xwos1gDwj2+6tplrreivPnAq+m
z2CunpsX4HVzV/hsDQKMRifc9MfxeTdpN7VR8SylTEORCZ5ZQo1KDs9lDMH+P2VJaVn50B2w3+TL
D5lrs6QF2WtjlumUExVSQiY5KYgXERyVsbZfHM7HiygMv7/YADUK+nlUr9kSHND85zAhcJ//5zxJ
iGjBfg0+9MSkETjE5evD3RakjJMd1oujAe7YUaYyJJ0jye7OSrodzcdPhyPYmdr+4vyAHF+xgbtz
JHIWk+TZFckdhMcMahdp0mJwEV4iYaPKVregrvtWC9xhSM4U/YT6VpJZ9r85m0JjkUxeJst3USdZ
nynWbk73vefbWGs42InOAIyYGXLc50qE0xoZQief5GgQcN6jx/mf7EvHGxvFkODg4UCbWgqElV1L
I1qX4n84ETd9z1/5zXMCOf29COJWdIMERgaOYfvpGKKSyiGCo4TidWUqQx6vlgqEp918icTO0k6c
HAvkBzhMqWi4p+r4YOvmC8ObsGzxMhabIKFz9ETFUUnClhzQLmxr/L5PTgC6xiXUkaXqAZ2Dwdbf
u+C6S65O90lVfQ5aChzUB6JKejxDSHURzXD7mn1a/3IhcTx1y3Q+9LAqiod+bbwAtTEO1Ves2wDU
r1ph2Vd6QvNIVqfeH44GaOwgaV/TzQy94gvgQpO/sHWgJBZaBdsH+/pQXIeVt5D+E2VRS/QqDdmj
FwUVYjh0jT19vmNPUQQiKlsHUbYzqXXlHjPrGp4qXIelXW1q5Nlkx44t/moeMeqyEYrcQnT3ZL5C
/MdZtTX5+/SY3tqCOiioaN2OMUK8VC1te+f9q/ztyScfPBEQ1mJJt6Uuy5Zq4Q+EVrt/LXNJly/h
PdwybM/TKTfXDtcESoa+nvEZNBdWs1VwXaTTKHi1AXl5Wlqxy4Z6R1k5BA51b/ySw3SJZfbfWUx5
CxWPqKkoydWMaZ7ajGCIrXIfWD+BNNQNGsx5aJd0gsSzAJCw/8paWXFsadAuaylR0aF/bU8ikKWH
zFjDrEDPL/bF9jCj2HxtRRq0wrUhghQvl4gkFX6zBJRxh75NSrVmtdAISqkO4ZYYdpccAzUM5fpY
Uhanqm3mqjORZcrkOJjhesmGhclSz2Ixbn1+U+02Qw77EvJD2VIcOgeXRn+WOe5QcVkvQQe3ygwa
OWb0uuy+MhEk12ucnupgPNovh8K4YEspyRAjsIOMOT5UyHcq6j0/R5EabmLnLNNIMn+8hHIJqUtt
c1ookT+hOdWGubAKiIvC/Xgx0y8w7Tn6FGqeDemBKFdLdxjsG2/3vzQpu/GKt58xWLWeE0xZv1LV
GxyDbDwQC/sytlSrdQhUodoPOQ9eYyPHuttbN67bdL7+JZoQQPakE3tcDHsIFjdFsptB1rjxsCxr
oFNBxbk203IMzihVVGiXKyw4/sORFJxk31r7eG+78pMA4rK1ix09NFNgJ64XOVIN0zx0nKfkMpZY
LJUN8HNwnxiZWSkI7xJ8NrT037a3NA+VqfpkuXwLbHnF6snJMBfL0nnL4G2ikl3Ss0Fte5ze+JEn
+0qQKZxRNS3H8/Pq6Rg//ve/o5qpBOgRY1YQzMWNQ2vVI0OlMSSWKmqSoq+DULiM2vxPXahu3Ct4
ox3cuAywEYTro1lcwls7QQE4VVZG1PhRUsiBWbB6YvYs1E7QKVsCx5nqz2kB1gA2g6m2VKdYFQBR
kpG7v5IvCJUjxmETU8kB6Y9YR9qx8+F6P5MhnRV/uoxKiQLSbUhanwctwvUAnjCF/OSKRfVnUbUK
hn3vU8UvDkdbEmgHdAH4v7k7Y4VeO3h3IYJquzG1VDmjRxbmK2mtElJrDTBXvCsH6w3RmNUaUu0c
hfOX5Ku3V857Qd0hRvf/pC1bGGLDNs1edWS4mMa/UtCFMSsbAPuXDG/T5djcBnm1RiCcaOeGsyL+
PrsjxCcka8nHvXI4xc2oQvf18P76sfq9hgpdjzk6q+aYckFes/SM0YnxsfLVhv9+tT08hN0WTBtZ
l/owoljOII56YFfCT71Fz2xLVSBCd8Z0HThTTaS6L98xVsMYn5es2YKAzNR6q0wZH+aG1o4CaAG2
IIGqJhuKxgEEW1DrRJptJRt6qCSGPAKvoloG76dvSAPQT2TdxTyfH3swfBYPqheQHSJqmdwCb40V
T5pAUePwvtlgmDkhGj6ujWU/393FkKcAEYPF//aBYBOe+xCVi6fsWRTxMW3c4h/Er65QE0HkFIfa
gy4D3j81WMHw0CQLhT9g8p+3ewtF+w88D8SWo0cd0j/TVJvZKFYVSUKP4oXeA/+jr53lVInfoboW
ut+X53EFAMyDiHJxHlfoyR6ZFQmiicx/n2qDzV8Tc0QHa0jbGZaHcEHokcSLn4e0CqlhbWWduPJA
s983LVylz5Lc0kP5lSl1jZfHqVNSCIzgsITEEqlWPS+uLChkJDJSYI7MaK6IJh2/mdCLcaXu2AQZ
Ls1r2H9AI+yVijoYu5Eac1G8HAgMmQcJ4YhKwTmAQhsVHOt4aVEPdDwrF9Zt/CAJlWl+vcN0f++V
m9b6Z2O6BXsnzX9Xm90Oc9Ed3botth84FOhtU2k+j0NsUkNxtEc1wHTNzxWytJA1CVOQPmTp8fjX
tM7iYJMAQJPXAyH9Bn5gWoe2CELjStokHKEELbcdq5iDqB+mCefKN9STcV3NwFmSRESyLiNMeXBs
IpbY1b3zBq83fAOnAI3OtzFBNampFopweRu273qp5gTYCPhcAv4DF4ZxeZbz8fHXvW9UKNETXTVG
OdDlR2ZlOm+4qpQFZZ6gWAx0LYkWPauekZp938Nv7o3ncUBWMkcuD4GS5QEP+jZe2jq68SBcuJj7
M0c1axejPV7fh3/rY1BnU4ao5X12cL8RVclhPPddcoN/x9oIRB4nS8AKiquA3wzVW9w+WxMXb6qG
BR1bqKOROTw1vrpV5It2udny7+tMfUPG9zsLA0jy38iOk8LNVUGlb0GoGgnYUQY32OLJjBG1rms5
MxfH5Vi8cnZ2eYWehyeWOYiXD7MweQeFQhfCPzjSGf2lDN9qG7a+zG+UFhm06rIem3shOfORL18a
EqUPACBflnXjL1W+pkSigAL3TEVIkaCbK+XW36lGtyYNaKbf0vw4UgPDXghYjtZq7AlGtJSeBpXp
eFJJy5UdR4IoQs3GkNUHuIhyFzcXKtq+6NCLvJGD4ha3JhfMw1LbBUQtL2WSdJBSH++L2U0Mavdq
MLVlKduNK6OvSr5Mu5m3erKdYFbriAJOZXyzfuKYm3//vS3+Kj/NstaVv1Q3C07so02FuDI8cLOD
AJfLRa3216e11T6ifdkUINhGJLQJv915GJXuH5Deq8RSXMRxm0/RJwwhtCdanFRhXHPmyD1zeNRB
blQrUiiBivo1ukm//sffaSjv7V0wmthaI/8+ywY2zdIMdVvueurwL01OY448f236j9H63gOTIpmC
t5gHdQ2e4qwzSb3o3gEUKZX6KHycnLs5BniDpeEpdI2F0IzQVBMZlPzB6tLz74QE30SuqB5NODh2
PbphKP2PQCPozsRQ9A2F2qFVM6LAy7iHhZkOJ83yyaTd/H91AuZ75xweRyV/ybfhw8xybCUGu/W4
pY/aQO6TZTs/JbpPEOlAv5lzikTjuien2CRXH7N+HXlJ8Ro1d53yRlbP3GMC0ln3wGe8bZqBauZ5
dnjymLtQGuidrky0GSG9qtovJnuvDS8qudY8fLIf58W9MygkWBGlYcKZKUb5OlBxFHtbbEBndjWf
teNv49cKfm8vyTRTbLBTAz/VZn/3AP0mzVfhWf2UfFocLRvXl/lvhLmDb+cKNtwZO0pd9QyYCKFD
sa0XQndkx/dA9tmCXXDwi/YzJjcrfp3/RLCGre3sNXteQw1vYO+250s6qx3sAo2a85O1uvS5H3Pl
VDnB8+vI0gwqOL1CZC47jSQbAE7RJpQ0AwSDTyRJTaVmZfuqgmXWLD8POUInQM0LHh8N4o1Ou6n4
xtsijh4KAA7YyCGtJbe9hZhtr5g3/W6+8s5gAP+7EtoTeoJjKx85GwOmhdLdqc3oOdDcxKJOGbIk
5PiO6pvfkiqm9i28IJP0x65cevaNuBXZuFtr3JDkEbOhsfT5PWnetqQl2muzqakqIH8b+NQo+0kH
oS1B4648aFMTb6Stj4nrKPU2WxljL8MM46jKwmSF0UesedRKDmRhQ45RaxlOD1J8n2BmToK2xrsw
1pNyL4JQcA+rBCCP9lQZZgLUxImpntrAvkWo1Vf44t1A6nzAVNFI3IZAFG53D0bOPOHdS+I0OsL5
OvNq0eZzqUXOd+S53CCCxkQ9JJXvHY4BVwo+ZTO7pTVpzhtvHvxYxyhhQS/03bauszPfOdV/b8LX
lKyg+jasXzVSqIg6/9BHUASoN7IVbrietr+pqrgXDHS27wwrwJFnZpYxybwkXNVOen4eYwCZ27+i
weG5PVOC2BQS4ysujv6egG8A8eu3wlIb36MdX3idFx3A/vqf5Hd4l42ZfSN8okdR6cMchJyG64jR
uFTnFktKGkv2VIhyfa6HPHXb9w+Qy28M5cmXIX+eDzH7pJ3l9XeVzIJkeN9efu82u57ETm0oRhkI
sH7QM9Mldm8v1mf27SpzzXj3Xy5NfekLIplhRNFBy8xyG8bvdxijteNsjZQofH9BxPM7o2v/LvGO
Lhvz/N1qB07Hu250gK8XQQ0iTRxGnCes1BsxpMrudeSCtdw9ouW/6Jmft/kOrJS7cw0Qy+YFO8Dm
L3IHkf+TxHONOeQ4vMnKhnspymGqOv0/4rh7ANByyTLuyosigs4GMS4aAmuZeRIHdFsGXUzif4aI
9ol/DBXIxuEd6BmfOxP/vyVz2rLEa6m5cobgA0UhnggdB6M1o6jp+LeYKVAqWB12e7mKG0uVjD/w
RG+AXwz/rccM9qG+6kWmUbWrQxg6bnlOa7IHeV23Jd2r3XNnlmMMlISFCtjkxYshuKSc7YpXwiVB
tMYG8npdmZatCDYYX2pcDLPqDcRKaNUdsaijjvAyoSSjhxW5ckqpmEN5nuhoyWSzFr8vrL6RIkwg
4rIzfvqCT7dr7YnpgXImo9uBaaILQcofUgyGxjEXrj07nbBwjxT641KDh6zU4j3V/T9WoJdFfPE8
+n5GcpHxGcbdbSvMVIn51FXUQBnPxeQGUhm86b1BP4t+/8yx3ShrOCMXJHa9RqPLwaJNjKH/JrT4
bY4eRyd7SY3QdfEibBDm+oj7u9IDAANyoifjO1NWKVSnRZhua5u+YMBpclttjDDX40y4gCU68Tjs
ehcZ9SgevBshchaX/fOaGO53A2/Ut05P5jYSWZVpLV+L2cv8GElJT1wwhuFExzguAC5nDDc2gjrf
t1ygSMz2ydYqj7afu387UWBPG3UTX0Lbep53x2hYub45OGDkRZow8P1aZksqzJ7tGZuGcpK1wI/K
4NdF23wFRTG5Ixh0pKRX2UIcAsxkfKzVmn8ZspjAIU1pJXhnLz+hrBTx1SVTHKfrf6J0Vgre1bIN
BGMVm9PO16A0ADIii7uHeLHb1wJzNDVteXVHsY7/pFLtaa3uGVH+4APorCSXKjxKJ6zzdhSCqGPl
RG0DndQb7M0/e/P+Vydz12PmRz1FoiAnGEp8g+0kE9GyHcdEzGXxZzPWkhWC0DjdSFOOY0lcimmm
N8J0hU/H5eC5J17iakmYfPsn02nDcnCljaEv9h2HJ8t9ZJOHc5rQFo5rEntCPFGA5v8fa9ruplmE
EHQ4AEaL2DEtJ/W0/k0kywo1yIIuXw07BNAdnjTmD52Pdo8HDSHSqlP4IZsxAC7LV1w8bQQ2KjHW
pnYPBVhbqct7YmO8tIAxfAPDOLLI/daz25R2AgD2dZStYThZyDbWkJs3C5e2LTW49prbWrlVRCc6
F5Q4OORxMN2nwzE+c6IwZBM2+A1dYfq+M9rQOuPFJMpOyaC//aigUoIc/Ce05dFVZSGQsijazF5i
5Qq+NmHprQjOGrU/VyWuemr8/snKrZGrT8Ob+ZGuj4gJ5e2awzVqyO+Dak844JqFBYKM8YwY45PX
9F5HGfpvr556rjTI5VSeJNivl43uL6cCfRpCYkwEb8+BdPciFuqf//JWb0xlVdOSlMH0LIqefCaK
ySe6bPRCY4szQaTXmfCgKPBoyuf2FuAeg7RTAzpPQX3aW0KV+MBSYWevZZyRox9V2YWZifTKqL8H
iUHKckjRdfcyAbZCvwU8eJeHOInoy7qZe5PmEeyYsVL7BFYEeQXfJcM2gtk7uYJA/qauIdrgTCjW
YTMUaSWtdFVHdqEy9LQaryWuyMuiMkzA6h4/+D8/RyZwjqz4x7k3S/mGSRXuHODmNC6O3ByFbnFa
1tB3NN2qOigLam1RNOjgcdZw9XS0cJvEOX1jKGrdb2cQZcOi/ZpiTVmu5HAz9y66hjMSo8G01J/E
DMDTXnZYfjhARJv8C/Lp9Pw6VMel/SruDNwOg519z6SgX9mhvwkO7EgBp8i+WzSp1+euAHbPj4Gj
NNLPkAQl3bR/RcKP6orbo82CtvE1dpb6Hb4sNWRG7WmNThxoJwmFce+bQ3J2GRNiVc+yrp+skJ4j
vkv9+AcygZmlJ5XKCXoZBCgChIKVxJPo93HP653kJroNoP2Xhh0VWWEwHGneNbvBfAsTc72K3ygH
kI4SGwh69QBaolDCQJjLi1AD2gWIkkVou7obZS9mtOmpmP5t9nd/OmZlBpAZ5Gsc/HTx+yNjQcg1
BbznriIL48edvpR+uVk1nw7ZiDfDhenmac4d8HYWfaOZLeoHSWrZgUZF6lPgLpVwJXJgGy54/Uds
8JCwBxL/rRVLnB4pX15yFvGRx4d8HadIJrkDezixnG7Kgks+BQVGHg9I5TLOQJ2LSamTpsP1C0Qc
L5++49mbMBNphgac8QcYQ2IyzF7RYD2Ns+dolJUldx8b+hmZNyn5IUIk+QiGDnhRbAGF6erOtSIg
cGA+nTzJQ6To73gtCSscGmANRldRDxKMUGCvD75o7hLuBW5/5kSZwnY/ZDUtyAF33OEg9FvRNUJA
4dWhvWLtHZeimwp9aN08uatlehEa3VrRN4eb2jdiAjGWw7Mopgv+gmIJrMri8+vOY57AVw3ZLn97
LPAXrsUeAZhop8ZO24LCgMYJB+/yQq0r6E2hPNZSLbmLfZQRmYJw6XJqXUjSw93+dcyr76ygEZvq
VblmId+BlVvqo/6Kmr1YT6uZ6Zx8MD+V0HIrSaWqzZCD2+SeXDhjGyQ8kuLeAGNEVDktAvwwzEyE
v+4FgYvisbPbPFXCKCH1EvS8q+7dx2Rkt4Ka9OZDePKqVhT8ilv0tuCwp+mTkFlH2zvUVKL2uOXs
Y/IpntQG0w2ec21LS8VMx8+JCsaUZNals8jpaeLRTnTwGZVMB0T+KviImgeY6T7pNGN6JjJ+L2M0
ckmo6VRU3IVRsUEVUhsJx00GvPeztO1oNt8ltDBWsUnx6M5mAMgGxF5E93TCfQMrnFLFXy4Fawzp
RQ5ZmjChL9mep6uun6RfgCmRV2acRsClZfHmC7Ukibr12T3BniM5/UvRjh7VsT+TJ8KH1CtBPfwB
lJfN2GsXPFvBVTxBtxY/ap94UWzA5j8ZdRUC1OOLAQkI2eOZIdt2pD3KfYDWS1+H9GWuBrarPwvR
jiHBZP/LUprkfdvWuyAe9p2RmjTiWv7JB7ljL6Nmf+PFyLVRSM4qermOduon6bQK6hFNGEyzjjOh
hSpKzdY7GbjRbs5drT6Dx3rjoFiZ4q1R+/zSaafEnyr0SC5nAdrcI/Z52Em7inzjZTjzol41xGn4
BzAuiLpBFSTwsqlY3l3YCxn/S+IybL1TB0whB4saHpIdeBf+KJ71q+hhfBaAFqK/l9VwIq+zK0IW
Atla+5RDoZ7qMWtCnPc9qBD2U1tXXMyaBPFXr8sfsAj2rOUKYVmZRfgrMVs/WRXHXQ3C0uvNpYPA
e8i1l60XRL7nZfWVpYgCzcnQTYSRdbf4pkSd01NUT8UtBRa5St1iQs9Ba9+pHI+n+mcaUoPj5BV9
etl8jYa5Trx1Z68pyPKzpFj8f/V+90ObnZiuhr9GUY0Vq6PDjpckXZJdnSGRgiW/7FSWxtP4cWHH
rUVSq3WRtEFNwYXEyJyNRFNHvSEYRgdxBnFoi630OTurHHmt1rd9c6koo8WZXXrYLtiLYfHHWIWh
slSUbSxj4d/N11DGWBODJxGxBrdDFnAGAADDUMtoOQEtKoaIA2WDnySpRDIeKtHnlbzqq8j2KGff
4A4dCSbSIn9m7KsvreiQ/niO/iKxC0PvyWRKJXVTZMwk/MAs2Ww698ILAeBekkPro7lqtm61RDzr
fLdLT/1PuK7s+N8YBvLOvAJDZWygsZau9ay0+2xE+mfQbpjSJotGhEpDIEGZar4QI/f/2GDuzXQl
R/fuQAe/TJN9hnsGG36CaD44E5Vdxi9LaQcFwvE5Ycd6x7ASWlo2XwAmDfFejk+T89s5nHYxa779
IgSQGGDQVGSdoAaZ4KfDv+WJg5b5DdRSfky3NgnNuxZgxPLgq8tT+TBSIImiRSsoDbb/QZ6sdnAj
9VLDES5eIyGE/HCzeikiBcvFV16D5lCnRBwYLlXMTyZXyFAIcbUh9JEF6tZepCw1PtNUkVt3vdGr
QzqpvPH3ikV9Q5wHIt6uiON6m43Jm6VKopXwGUVhgWiv0Q9aqngRXy+wvQE2XGxmTTuVBygwNWKj
elIywXCjq4qTf81z3gr/nDfpFcmIPWbWtDAig62JYQaZnBg41Nr0yjZV6ItWET2bciIGaCon5h6L
upY8D/su5lqoVwCLBWbRNZ/1SXZEkNsnB9DVYANkb5vj+Yl+txcNptix7nWD2mA9MGjig1kTCV9+
XsNWVHO0NyW2FAIHhc68D1VERI5dQ0ydXLSdaedtg/6bZ+OmrC5WYnE3VveOFLbvcQFn5ojmm24D
QGx+9+APMCllZ6qxYo/S+WvzBHwQseNL1m6R/wm62+GUPG8+fa9TciJJOsKsQbw0T2HTNnc/LbAg
aYC3DPTDLKpqsu3mqpLLfo48pbXvX2q87xApOIqMmmj+Umq9/uvZdDaCpQ1RBYIXOFF5RZtrHpuN
o5ToOHoEJBIs88wrJBcOza7LjlP0bMyj+uUxe2u7mVX4Z9bk6qOwB4aqUb/XnAwn/U/t/9LCLTAj
tqRvRdSrIsZfjjn9AzxUKfINxA7jc8QSGzdUXJ50+0HRAfiHzFu/TuaR3WCzZcwk+qMgLiRmRq5K
RbLq0QpSmwYDioGT/dvrpkhoDgwgn7tCPb/Q1GnyW2HUejHR2Rmu5KQaiqmD8NlKGdetuwumBWq1
SDZmeRiaM4WwQXohyQOrG3rnMMHxzAVD2D6jKngKwGTntKnRRxPhqBZ0S5bl5sPDztzAAzaUjfPi
vT5FPRSVerlmT1Y08C+pgjnZ9OYp1XHH9siIaStScsc7RlSmJmyM2CGcKGuJRAxmIBcFLkvdde6P
W3easJ/mfcJ+7yBCxzaP/sWqmnH28Sb6ws+Aw5x6MpMKahW8FA5jZbIiMKArlKSdPPVHsr5BfT65
x4Ww5535GYMxEzKN9pg6xp4tQdylHHM/HUqja/mJHgzyxLgGcMcmKdh6b22ZZyvP6lOWpkSgRlTJ
TyehTddD6pUFlVp3wXl5uWA3P1kCxtFpVjUCbwEj8rMVlaVefeJ4cSmM7kPEee/Tjt9HtG4NVET8
3wqc9XasbZb2J1NnDKNN549Gslm/bhHlvqHT0FaewORLflAOD7rikPHgG68QL6kbE4tGCciWb369
NMEzo/g68HqqnNmUWLrIbadCz9BfZeNLOOHExAxtHbujryg4SMUagERT6hZMU0EmbJxDKnLXdZX5
pVZ3KsRXyP6MxMAK9YeXIZUJ4FzUVzCkxJ500eoiYmQQmP8NgCV9/eKb2un7BXK5AHyBzcloEX8S
qjpKok1yt/2cDhqr04O7m3OkSW6U3F5uBxapll5Za7hbMPHtVHkJtoGgGHLwJA67WCj18Bu3t7JD
1VTtGPT5LvRX+snxcVs8iOlo5kiB4d2aHyxsxnonD118gvGLLUSDvlHVePWQ6O8AoFXjOETttQKZ
wCDORgO9znO/jKpzHfFAFLrXS8cvO9l60ZUbIS71uQxjnSCXPI1L7VizsbKLm1f8+/mZRFNbFfm1
63SgOu6uSBM+yb4bQDhoUIiJd3XfRGC/X4EmY75p/DOBW6AbE5/tMOSIhWqd+ynb7fv+arXBipml
Za/B5pEQnvm6/cvBAIU13jwSNlT8gkcfhiu9nWV3SJ6+jq3gpScRGVtiWFxWh6/LQYuvoLr6ujrG
C9i2uZl816W+jHxJG/ETw0w65kMh/a37XW543lEryCLK0pnhIl4MMoQ/QDKQlc9eNVLP41qw8Vu3
Yl7kp7bWEif2CB4GTR4llQ2BEw9Ctt0qRkqs175G4eimps8BJGZOJgG6Fh6gABu/97bDlIVpV8Ky
knc8Tv07TGhz0ktKn4Rc7lDD4PeE+lCzzpN8+BM8kXtGlAOneN9h4NBsDeOql9uE56HdcdtZ6qA7
HhbWdainsHTRFJzO3CmuF1XdZGc6UFdQBMIz/kFakdVzH/qmrn+nora4JvxssdCQcPwghwsk9DOt
dgohaLGgDGK/vylHRM5PZFhD9oZ0S3QJWHUfgIemhuJ7T5HBx3JUhagS5uioarHExRhEza+Cghos
WAY4vCseOGChXZCdpLpBUQ5fNX0HWh9/GVqyq74xaa3A65N8uFPebT5K8f7CuOFsMUTdBkrohkXO
/oorM9lZPurrMjjkf0afq2Wrj0G5GW98jS3+Sb/hILcD9tRlwdmUpWNhcOhKTt7AY0kbluQYsDbH
vcH4YW/QKF4DznIXYyZTaKCFfCJvnkVXkLdkq23pTC+C3XxVuEj7MVdLaNYvr0icec5myxRGs4yw
uWxyKo/+VQ5qzBVnoVB6veaCJvUJK8dTuMghZLE9W8pP3KCefim9MY/XGrRYUKws+Et4ZUO1gR6N
BX/f4A9XoefO3yvnS5pAY31qoW33NrSEDP0FjKg9eDaMpGkXfOJkuvwFdDGRHe5EJeR468N4PUNO
xQ/ehbvwY9aDtfR8lkNbXA2tLu56zfDALevqw9OatoJaHZDHpxI3tT//qUX/v+WUaWQKCwV+JRbH
GJ1f0VpmOvndI9Mtj0ouV0H4l65s8w0yFrh8/d5rwOStEcV2HWGsc78F24/1KxH5C30eR+SoG4st
cEVD95l63AjNqyz50A7UltAEsC28FlaGLxojNEWfo7bV/ZY36PLrCZcPXaQ6SfmPKUQuWBDoGjMN
/FC38S1zym1OVmxapsPKUlp1OD4NyCfJVOa1W9ETwfvYsPIPp3pzqgmEw8DPfPZTnjTJNh+9tytN
u737TP8Zvf0OzPNkU2N/kYdmMzNegag5lQYTJbdiR6nW643RFYGYbuen3pz5K+wPqObFq8ew69sb
JO56hDemEHqtzf85oPv2OMrExVxs26mPaCgisunkt3rWgGDooKy2UJhPPgcRdDqvxQ1iUm4ZDHtT
fkGfDt+JJ75+389R8ADh/IwuD2zaLQrjMpQw7jllhYOPJdkMLp8GQicGd08fiQRRbc8d/b9z4b05
2SKrv9lgcjSOmaVxitZ7ohizNZbM3Xkq85f189wpEANzWsuio6z1VjaO8qXbmDlbwc1GiCQZA6Q7
MtbxFIfxEY9YA2RbdMmNxZf/b12JaFyFezdAtxVewQqujBVbL5HS7DLTKCI5wzjZdx/041UmPq9H
gqqJFXOw9dsXX2u+1VZf4M6X96t1ZCh8DPrVYDBGsRDil3+7mtSIM8/f2Otrkgqqz+jouZIDUs4g
zww/aY6NcaOJob6e68wwA/bo7hS/SZOThrMd3we6MKUlu21icqJvzJp6s6XqAZK36UiGFSGDrOOY
6k4h71ccqOT6NJSBbkyL1y7TgSbhNpOR44DzcddoRYM5AEgwooUxMnWApnZqeRNDUqqLYG1zpAgj
nE+o7b64hUblQrhlkdWmnK4aO3b3DboVSTs+GIT6ysx8cOKSzNXO56YVh8hNoz6Q/80d/DYxpfhb
zx7S1LvthLVW1bI6yJTaakrYpbp1lK7RURYjurrsMVj+I7JAEoYkfJN8cIk9UTJICmE4ozDl2Ap1
Vkc8f9a9L/+IzIRxf3u0J8BYuqhz8xPo3lJkt5Pf0wirXUqs53im1GhNE6W2R2kSTSUQdwgryxQ6
BrgLS/q2oLZApxMsnqFign+lyAnnu8Fly4cT8Xg5BdkBcs865NtG46lVQ7IQyLrekoaMGxqtiC5/
+TsXpNkNdmDP3A5jD2UhJmWlicjoRFA7PosftdF0UrZSdD2h6YGqMMO08ZCj7DoOLqix3PWWIG5G
g8IwdawGgQMgPjqbHIKj5JWIuTHc3s3DCZtU+L2DMQsyI4sBSn2AsEBpCZiu61UgQuf4xJo7n2fm
sMspROE2Q/kHU1ws3Pk978DWCiveQ4JuKbRSA/HotbsX3E+Sm4lq1NORDB12FM7Y6zKMvwlgXC8v
INWK9cMU2bwdwfDrx68AVFJSZCFli+fopM4nahTpua8VdDGFF4hGz+9IFw4+3LQGQG3wrx5pIg4M
c++rneJ/DOhS1JFbx9b8/2DTo0Sf1SQNVvD5f6lEvzwsS3qh4zaBas7oa8KE9bGXeKudDIOgbyNI
X+q4J3sYmc+o0rCuvebiHiAtBlRcOXrStA5pgK/qb8NJp/s+p048+0fEHJQKoDFiVMvN1jjyevGb
KISgRQenx36KDFW41uloQTWjVmdICf71OEpZlSsRGvT2w8d0yS7AvZA0/59vVWcYxZeGoANQhZ4u
eCueOMRkBMQdgkIF82F3rGNjtoEeV06UGBiuJtLfjldE49XCx3zekqrJj2zftj3KAABj9IntUhr+
Flwvp99U4spb+83+QsT6MWYMKt8v/sslmaSyffeXhkNChEjg9z8UdMSUqR1m12k9++08rfAfgPOR
Ot6EvHPAcZSOEEXTF/UzVyh2kCNN4MvwR67ySa9Atoa1VI9B1S5QiXquuXJdUQYGQYef2pxGTsPi
4kiDF2Ze2c3UoMnnpxnwxD8WJqZ9lGcZLlCWnXW4uA8KE6Xd5cLU5vWeBZpXnJEtHbWSOVI8uM8v
o8xXZQ/Ki5BDlajeybcQyMnwfn3aEYW88GZWna+5MCpR1mlkWkozdfnfPs6vmKWcTrZCFcQdY/gV
e9C2ffgJL+hBjDKpYgRveqH8m9+uW/6cDCxHMw2LlD6spXVvRZp4OHLnx3665+XehN1HsUiBqsv6
Jh827lRWQw8Xs4xsnd6cv7jvC+InoROG/uI3Zwldnudf8FcDK9OLXpQTwV8+kxcD+Sh5zg/BhT3N
sIY4mz2JUHGLSRpvUX+SQPpCBQ+QC+B8jBuhls2l2xPuShOAOfX8TYCMM8cknFFhCjUrS4eNcUuC
qJbJ+63cA/dk0Bx9JZjKGDN0fFxCiWzsAoZfNWVqy/OlVkV+XN1fPp0pb9cmZYIbOqGicjt/Kfex
Mz6ID7wZPeNgmmu/mmkpJB8sJdbFK6b9UF0o9Xm9LnggbNAw5DHru9yzdeJNV82zl7iQTKukP9i4
zqoDYPs5jwAJU1jOe/dzv4SjCpbl0qHlEWzsVJaG9vH9iUIavaNSPk5jLt1Yw+AA8i/b67K63hlw
tutLPlZWEO8rYyJ9HDZfTGFFH8Z0iYnOHqdicgcAFgTAj23GiLwxgJvtYUnc2FUBpNYqlimFPDOB
ESpnuxf3BQsTs+AAeDvJu/nTQ8tO4HVJgQ/mpWOo5Alzs+THzeLRdfZidm+km4mMXfKDdglkD+X+
AXRF/7OnPf0nHkNCf2VbqnZG9ntTqIkVDTgVgkpD0eUceGYSnFbjIIMy58lfmu84lUODrPcbO2Qj
YO3ekW7sNoMEHgtXsaNtQL3k32XoCmBrZI84C7V39lu3z1ezR6CkD9HVFE52fkkAvbjJ0btQBX1c
no8HF8NzCcRDbIAzxrGR+gq2vpZ7diiBbAiOaZJu6ycN2F/clGwFrZGxgdaq8uwHAtKVifuprAC5
7eYkFfiQLooSLsWzurMw9T2zo/W8tL2kV+sp82+/KjcS2UnjtcZqIDRBHYP8PZCCBv/mRt5C4Br0
Snykvoe172Ft/+d4M3VaLwNwvFeXPkGuKDwQNuX2iPVwYG7inNcJJIvOMfUf5d4qId7/tHRfGlXd
o+c7Btc7h4PJaS+taBEcgAtIpVwBNwBC9CJwyQsmUBRi23GNZT/O64Mj5iqYc0JUoEog9UIUcgnS
2rY4iMz5hm52xosI0puBvJ+TNc5JFoUuCrX6gceX3WiPniW4cG5M02wfB+Jnqg/gtN3R/hCdr0Yu
9ts8dGG6ec8ZWXHBjDvdKGm2Q4xxI5SWbXl69UHMfUQiykxmaANaxYa+5e7r/h8//37FcnoFp8UO
+KdbMX8WQ3EH7sZFGNlwh4ySFjvzIfWE1hA9chBDhdXDJpm0BTnlNe0Yxh6tMYKW74nSVqBNF6mG
j8+M9doSAcBmcyDtNwR2RysE9D28McgUreXVbzfeZdikZ9R5vbH12g16I3N93Nv5koElSVMVnA/k
emTwVaJkM4toiSgLq88+9/ka8E2xKhLr/61eJacpT3cD/y1BHilSEd10ZdgLzWjmO0STfAaQTch3
1Syq9YGcVo3MhEXh27eryK5NE9i3sfhcocl8F3sP1R/m9BVsPjg4XBMQJwMYn0Yya1xCLN6eWlT7
mkdk4spWP1HGpST8nCBBCR1DPsHYXtH9ikcrWVrAuDF4YA6xCVsoQsH+5sFvuq6wOJ/LK+ElMvxK
U7u3rvwRg+vYD3NswW8NN8TmRpK+yKZyzbbjTBaI2qIG14HJelWImPbHlBSLyUN+NrodXm3vA+hE
1DzxSDqQ3B/T30cc7nhzeDwqjREZTNutuZTNrUlA7T6AfVlh7ZXAesppkt+hrscxFviW3C1VLy+J
39oAitF8u69qcDvyjZWBKAG7zSuKWbIQ1ZUZI3Zk2fxqsvn29Fp7l4mAXU+TWUTinUYu0+266ov5
bnm9pL1KyDcBKfB6uRu7+NU0yxzs3xg/vJamDJyXIvObIx4EkC3OlgFcbb7AI67L90b3KJICHJP2
L777iXvrJv5CeADZpXz3xLaTqX7VCJkAo/O/JGRBOeDNWVpZtcOLUepQ7eD6WyfINAa9IEx3xK7U
Xbli8zHlu6Z9ecLPopnvfw3eYGLudZprvyb/ve4NZa1NwWY0z85Re0JRp+Dq9QwTyO+aSyskDkHb
519bTnHNxzUxopuhwRWMcQEgAx31+kciK9XPTqJnJE3918jVSKdSPGAF9hbad1mP2DcK6a93/XXx
fZZ5n2/UQwJgbx2N3AF+xFtpg45e2zqofvt45ov8e6yvn/7bQhiRSjTb99BhlRuky9DXsscDItll
7oulnnB1p8OD7wR0lfGAo4ExMGc3Qyymmm2NCfFnZPj2aXtEK7WNqnqc0KF+3wtfLZCnyG2X0rCu
XApwm6DIcWCAzIqSJOwJq46sNKiEyVaLp5i4PMZv4F6aKbVrug12gNmFzy5QzWHYmXggwIJCaqVM
RaGx3d5cca971+jI+hDNzhpIjA4yj9nF+UVqgFNpZmVtXCSR/hcilx1U+mEqbObVsfWrFdJRMxA8
JW9c2UXi5kIcylepinZrntKu8YxBnysUwDMWUyiDgQ8Vh/dlQCPapZpmfGA86H27DNkfHtesTDqc
miIVx+uvXKtSnN4EmJxaKBQIg06ysfTttlWbgPZW3/vLmn99nDqW0MaEomMiBflU16t0uNm/Z3PA
WDdDeXIxMuwIohDZ3zmkqqoiyMWSzakK+puoySqdU1ldz/2YBavyVvFuHb514G0gHt1R68KgOLAn
FJjgEZWU3GwQ/3xrBfNy4sed5lcjI2R3Ioq/3d9zhERTB9602EU1l9WQe2qYqBMTgrkqzS8X3sgQ
hK9sIGFd1q2wW5X9vcdIsxxKNgHnQppXI1MEwi8HqIulfguThAlJGD24aJJ3aVETf0W+PxUAgeZ/
YjNqDy+zw2FJhmvKGNtBZhqk0kkoKnAf5vfxUYeZvhA4x6UHlBmT/ztp2oie2iP/YK8wME/VGm54
3Jk5maMI0qTjspyxrht9ASN029irz2EH5+5HiYgGlnxC/G5RzWV9w4fGEpX08PWwULCyP/W9cM3e
x8XozAx5L19fe945vE4y6zocGLM6BiG2tLkng8kANnN+Fk8awaQP2NE6jdJFy5Ay5aJbuemZSRwG
zFeVdX+E9Xj0moqmDugxYQeMLPDQr92IFE2q63lqwHBk7YDzKe/2/I0lyIEaDcdRqCRNflQj+z28
iJZub1oiYlo1xXqQMmHj5B9C9fDbk5U9PsqnNw3f9relqG5i0qI6gvRqxpq3myFJgOiz7bAdN9Jh
mAoaL0UZPl0NH0G0GkU0aTOsdI2uc1+d+hlds5mP6v52ePApDo9tO6ryJvacTTTpTn8SLN8GNN0p
tMqSg9mpWPkHeSfu/+/3VTHDDn9jRYSJ1MxU1MPjfGeHmylmPvvzl8tUFNy/7DrHihhTV7MEhyuB
cxo5ERtH7Ux7Js7ilAltHN0ZIkRy4RwF0j6A6DcoGwXY+i9GOUBiIooqj9a9O21P2dnrI4LO6H44
WUVL/m0nznmktVP0gZAn6VLpHwUNSZSl/Kxe4kkBysGmr7eaEhiPp2LyLqZSkzeVIhyUP2HZbbx5
WeYzaYkrpr9WW972YqzsyMzMRrPpqyg0bsUCXZmsjL3TuTK1emY/q4m9CvNbqQU3KBmUnS6I5259
fEfAJiHArnvZ3JUD+mlW2X9nITjDIhk7j3XYg/CMcj7+0BMTs3dvxAhnUXcEqtlwK/i8wYUh2TVp
caXkwMkYACxGPgFfLmUH8OFY6HKj8hqe2hJweiTkcFjO1kSNhq3zfD3mbCfeS8wUPIU8IQ+jKvFc
p4pg5IbZqUrAuL/QcM/I5a0/b1ydX7ftX8NBsfS8FgouOShf4b1QGFd//qEKFMsP2ihLOw5xdy+/
qOZGlsdrLjZgZLKZEJQM0scB3+omTSnazMyyHmF+D0zjIspbegWe/FXiDkXI5As9V1WAACakL0e2
GYkNE2xAF5vAaRw202vF51INlu5BPd7+FZFuW7RXI9hV6DCbcUUSLu7qPaMFOskjoq9Oy3HqR2ci
FRgtAKW0W41r4Bkxknw/sI5HXhVcGA8jwGWtrNK7PY5YVciBQxsbNIaCqiH8MO1Zft73Vp4j6ZP3
Ct3v2R/s7QENAK1UGniNjz1yvBgjQUgTKRFs7o9hLqcbAwlO3PRf0hfHVONgxXdSgnLihmsIJOsF
11mlHLIaFt96PLo+qQ1492fEf7h/YP+QnkFPquYTwey1vxkc7+M9zv/6AGQR4PcTVbCW5ELh4K8D
hGIpNoQorxloZr8ALh/rj4NG3b8m2yuOkLTLJjHjHN3MkzEPqDOVYMiyRGjIga9oEv0VPjNPb0NX
QCOeWTAKbBAnzY27o0klvj9H5sBgatBcRD7nxYvMwiVgA8Qw4tSPUc3YKKhveKYJg95amF/UX22L
bd/gYHL6SmIdgPMZ9Ze+wxPPduxx6JOrU6N92XaBs/mWFsdevTv121B/M3pOdegq07RSiWTR09C2
4lhJGqMUO7nvfOMVM1spRRjV/3LqG5IOS5MVS130eQgJuEXlzzbFDZjwJhLr+3GwjF8iYgN7aqFc
gSCEEyBeDC5qd/0piPMQMsruwK79wNXB2EXcbY3lNult09JCnuOcoFtiUjRwYGLM0Z09ucC92lr2
70xtV1wWOEc4ezKuCbCRAPC0Mg5+wr00uXWN+pOMiu88RgzglQzV+/cXCDevW7OV4sRMr31BXBhk
fptE/6ZyRt2FmE0R6q4XaHP36JCmeEDm49LrG1J6xNHWjYfEuRLawQGFke1PutTDMTSpPu4EIU5F
1Z7gT5k0V1hUjXif71ztDRG8MJwx9i8atu/VuH4K+D58cWBtCm01EyZJWbY90R0IUQYCXIG2ypKi
Gy1SCMmMIDjXt8U/RK1m+jbnOvr4NkM7atGHSsfsutG8V/Tqw08U3Nv5+/kje8WYXE3MZ9jurwZz
wcJPJwdh00iEI0bd3+6MpgZxSN+Gn2q1xKy9oKFFxp5q5jsGA+gqg1m8lQgRzMAsJADMk5rXClYh
KRXZlN0zzwN36F0X1MWdQoqjpXxj5EVSM84p9Nywhoib//bYxJBgrmSl0HK06l9qU0l07x2588t3
byVkG4+QyukXC/duvQZvhaUcUxiRDKd5xWUhBRhthXpwithFQyEgv4WzLU2ZF4RID8duoSYxIf0j
xwMKPW3bjFVNx3EpRA5cgNfZS9UnTFQ3N1Ax/BVsyog/hogeVApuf1teTEutwleOHSshbNgCy5Gz
wnTonpB1KG7+tibSNVh0pps2vu/mfanAOJtDgnGDdKpuntNjmWaG1YpthumNtDZCP6IUnb65qe2z
6HtdDhNwuMMe63tjd3Q3tjceFRPA8cPhpS/KHmmO06zlP7TWMPqPEw68CaAP8y6dGG2H7E3wK99r
PRFoN+TzaCpRPjJzczAyp0sULOHhvBUdEKzf9eh2e56Dy0Kv3q9zHo6Wk3TaTJQEBjdL2w09Tu+B
s5KFez/Y6+lI9ojPxZrj378h8EfYaPd0QVO46TcsKtuU1vQNenaHtQ7GKiwNyXqxshxYU3tMTfDG
/8vJOLWVTe6KGzaGXtf6e0VZ67Q9AiwcSOKsYOLr3tzS+5ujmc0eoXqFHprc2pq2T9RKcr5N/WkF
LFvufMWQrgsDghW2cLwF66kKcbsD38zFXOoX7CVnhsx6SC/PtE5rajplP3mB3mLTcnwkiWvCAFHG
sHh0/sKhz3JPOR+yd8f84XKa+KUBu5qh8OWGw600PP2Oc401GTjOxnz6smPheoVUPmlnsC0+EsdG
IAFaeRGBXg83RZ2Aupv0/mWqQiB6bUu4ZrApPQmAf22tC44IUL4cltHyQV+tHdY1M6ZWHh8VxU3q
x7BFBB9dlhcPa6S9oJe700FoaCM8hXXWCd12oqn3Z40mmY7l0AarGx+KvfR/4O95WxgQvNO/Xpwe
3Yz2K4f4RHDI9JmpqPRN8M27hkaRtOd1TLXdvnMgXLaqavaOXZxshJhuC0T0EwsEuiFKnqmVPBn/
nR79b3ZdelTfdV/YlFzkI1b1oyfITK6s9n4ygNiJ1RFv9klnbq8zlsRK8Ipj1SUE9Hta3i2wlVEG
RvE3oJmCZsV98twyKbC3PoavBHYa/0/321V2a77rZr0TtGv5ufSPusOmBa2ODsnphroS647tfsIN
xN7/0FO88QF13GlSc42fqUbQdmBWmSRe1UD9jUFDeD3s0a+7SIXwANOwndwdxbYDyWogVhp5Ukdk
z5el2W+UmorqJi+CxYO+L2hwopW8a3JtBloQFgGAMS/YtqEFJ0mXBKiwSOXTssSIG7mqFvRy9Fty
L1SZbUE0lr7sHpIkBrkQ4B3DZ76ABmxh0LiouxbIKOFK046E2VKTnrCQvXNMLb41r1oW37enWXYW
iTrKmp2kbpniWolbzRvzOMBfWpASkDnUbTcqOutboRbiXcSWwtxiwwl9FHO+Ib2dPHeZNVqXwvqR
PJjhgL6tJx/syRXn1gRDP1h1rMvowB81g3Vcet6Cp5WkfXiCoviScki2MT7Snf99P/aue+Fq/LCo
7V/gEBiqDaDIsAit4/RvhxBvNw5Iwf3SyrTQSMj1DQgHcAhiBaymkdpN2tahPvM+3dSqcOIRwmzN
+XX+Ip25e0NhQoMad7O8mlb5wj7yD28g8Rn9sy53bN0i2aOM8TvDyapn96twp65IkiMxtlLHd2Ti
eRTCQoMVuEDMLTp+q3fqUSMzfE8htiaqdF6WT/GPW++m8os58n/6ohAyBH8Wiy9gtMDCQ3/PLtQr
oBxKboFvq/Ef1y1n++Kf1Y06PkzUrAJ/xfMUeuon/7eIdE26xv6xEUyzLORIFvhKsN1zIPNtX/zY
TyQtgH4MfnVuViOE3NsD1HS2bsuCIWTjf1Il57vi9bSVQdAkPpzVvJePORzSwKh+wu/hDnOU2RFG
tePV9PxgEPwCQIo3UMPEA282pw33b+ywaZG5ypk/0bDORHQBMj7w2yYA6oqx/8/0wjE3/4xVG1L5
YugjF6XjnkYZIh8IMYELcAKuOgJwU4/gBDb/vVSo1sGNxY4Jxj9CmTxBhDc64YrWkoroQJnh1bHL
irYziAyPjdBLquvzt0w6YIX/rb96veXpCZm7uVCv0urLmiaZdG6QyoNkfBf4mr/lze8WdOkpyv+Y
gfMMyv3A2x/toW9cQSihrYUr8x9CNYaqg+iV+U0Mf+fRtGYUWv0i/RgyezP28gDy62Yg181rjRM2
t7YqTXT4EC3kuLkD/nQggzE1mmArPPUkFlyphoCevfDV+KgEyt4eNoLjbaMuCVwBetkNROcbVHAY
VlXf6ZaM934W82ZAr9xx6Ubn4r0uD9qb7nR/IRkGsC9ssOO7aCzBklxWOHNcBo7DdOu01fuLvuXu
SczA57JOm7D+1jeQ8LFnpcX/GRbu2lSfWmHrJOky2+XC5TG7MYOEK1p0K+JY+wWA8kYwqeBJ+5aw
pBOcI8L07lnwX0fUxngiB1KV/D5aRNA/c/jfHSuSPOCv0iTRxC5y7WsTZvjn7QLx3H92+vvOPBYI
ZuMkuIHi5GHgvfPGC5iM8Ah191B/CDjv/jTiURu28OQ9rDUzu+z/k8TzpdZg+mBJm8Go9Mko8fjI
MW/RYkV0hxzl2369FC19mg1bLRYf7uaiWaTJaP/OTgKRfAhyapO6XQJnRRCNPOuH6314pzAa3ywt
q8VAnaJuThKH4mXVOWOkB+6O7LHPPoraK3hOBmMvp1gd7KqSN/jOSNFZrmFLj0ISoQ7pOgdzwFbK
+wM5fUXbfqEpm/zhSansoMGicQYJgUcqGQQYL1MI295aRivz6oUn3GXCkZLyHivoxBc8ACEblX5D
CSnltNZyre/iFkP5AuOMemPj4XFIS60qaRQOebqRNgHcNXGqQSfWYCrb/uZhhQNejnPYCw+MAtaR
p5Ew3psAj2I36KN5aNoFyHN0Dx5rF8yI6DKMvbZRJG3RVWjxaYMx9NsVCoQWGysxXVxi4xyZkre4
xNmM744UgY2sY7VAvGSGE2Zp0X/msVwfQ02DvWCNvZubWGBNwaSsEbfEZ8KZZZOB3rbUJgzIrQAg
cHsHexDp5pqbUtanLCMzmC5J1rBe3o0Pz1tufRSe8+mwVwt2hBKjVG1eqAm6W9l0ehc0teUoS2dx
oa96SAbaEsgwZU55eKOCd0WI/D1RgoqW+PZMa7KXNQXgCuKGG5kxwhd3nG4SnmoqnA8xlrVIboVE
48BYBMAJVQDTTHWBPHmM/nCLgUQY1ir7ojMGUVzur00sB1StOflWpGyyenCvKs7CiFWx0RutjxIf
Cwsbff5IwLXXDlwh37sqJlI+Bl/kD75UOrTDqC2WYpvZ7IengSXyC0q2PXdXB7C6xHaFQA5QsmE5
mUdUQrZn+OpQVU0rFkHDMOQmbKejOIqr/4EF/AfMBOs8lcgGeIi8hOkWs4A8N1mp5vM+05MjeHGE
bL1SGDrm94SGwu8yxNbUYnCISgacOkTcf80DIC0kYe09vx6Lu00y71j2V+ypOAnY6qEfpRsYSyAi
5wf1U60aC5YvzNH15ok77QBYiPOF4onZMEbKne+tFLWBQ093MbgwkhzpV0OA/Vj8A73jQAL6Z6Sx
Scl39LbXjHZM1c3DBiIw4vXVqm2Ro7TY5+xhn1flpWryxC+1yRD910lu+VLyg6u1bbJiKyRAvA/S
Ch9HuI+F+/3x91cbzek4q4rDe6CwZ02kTGiTKdXFXevdY3PYQQRi915AFsCyXhP6bpdc2Nq1/WoO
3XtQvd/2jqfbR305nB7ra7pNk8lXUXdxQrE3JhFSeQz7aBseRG61+c8qMQ0G4V09euXsTEmri/1R
hhK9YL2QY4/FW91vjLXIJAmF2+XPV+zkeAwogg8FibYMq3kxWYT+LTXL1mhjSeqv9ss+vlDl47Ty
fwDfLWUZmprY978P7eLI44B6nJ6P83QQpMMCvNLHtBW+iUDaXM1z46+4kBum4NgwbXlbnEz9fUTN
84A40izE7d6dQIBYhIEA4p7I9f+a21xAYKxMHB3kVMSsHb+tnn13M52smpE3cveUAn+bF+27Lv0X
y0AtXX6aKyRBMYyE4jX9tF1biVtSDyBO62ExDHiL7hmzV82MzN6xeaTZSbouJXbr78LY3ckLglRM
zw0HzCD61aorcYpbqZoNcVGK/G+UmGg7xFNv7S8UliGzRsDdzf44hRU8GSOCFHWxLEimvHd9x+UY
tic8MzBDO7bwRFGDoWC2x0sLbCeEgdhYlLM31ExNVgMWe7Ue1jKJl/mLDa23j538FqPnvgfi4rmL
F3zhFkWSBOhrbg5NB1Cf8vrm0RS0X926pOAvdpBiNBxFJUohEii2zjIUvB9K//SU4izNKcD12eDY
ThtD6pcq82LYDSmgH2O5JNkMTNs4urrNfAbhD0GWHJuHGD2eQNvjPQaC6J8MieuCGAW6xjixeCCp
AwrDp/rVZL+Cm0/oQ0s53QUCW8nSUJop11DKU+pFod6rfD4Joiq/9PxIBH8xdtoYamtbQ8mLsoks
mAj7xEIJOR8xvP7b679Gcw/7BY+rIbtLlnecd6EiisFWOxZuEu1Qu/3gfSgOXi5y3R3DZpY7dWKJ
y2A244/QQ76lj8NLSOaoC+VdtWuWAiiip1WrmPE1mBcpQn22PGjMhWaP+1AUYMW7UIlv35fqM5Tz
6YESd6B7jDboYv2WZXtCpy/g+xmMZvhLiYfpy7CRx9E3XaV4KtJVOW5MjItDdyaARLSDJ34yHxYx
M/Mfg0IDvMvSL8AOSeZQyv3AZDQ5Mz5FZe7q1fctoCpEUd+YA3s89/Nr8B5UgRt2BxCWaOCIo2nD
AXpCSpwIHa3pC8BuL7FLNrqLMwJMgINr1K/P+RaqE2266KG+nBknnOWdawjVW5o8Gg1HutuBtoCE
B587ydmHmErkF9UpFAhP33i9l5s1glBD6lNzkZCKYPcdnGtJJciPyud7GLUkTBODXGNNn8MkJA04
m4oemxmCuRwAbemqElQWj9KtJV4Fjxd8nqHiyT4Yhnj8La6F5+2vTbiJNvQBQXxjCU64bpQucuG+
6dXlKUUvYytCkLeazQnYzjVu6BChG2nGTWGU3Q3AkA9l8qYstcEApLqWKQx1QW/EIrwU1UZOCGFC
capRSQUQP+3/QHb54Ze3HCDOdX5JLOcwTYHMZ+5TsAAAvWS3zzXrMDdVR7l8F5BwPw/zOVRgiaOI
C1zHv0wnHVY4Qix6TRRpC/MhLJlr1pVGMLyvTeTmF39TNQ0CuvGC3KoafN6JOoSD4cjgghn0nc6V
R+gichTAqOiZSF3qElno7ywsIG1D9/EqxdorS2acIGW65fyLG11BstBNqk0Q1XK7BedpQM54JGcE
Qd9lwwvnyIhvnpBUUYDyxmhDAe8m9XDGgKeJA2efFbe2Luffal3ZvZmvfi/Nlo95nwzEAt6uScTk
pB1+LfdCnrfuQaMn94rRDpw48HPq+TrUwqmnJmnynd3hl2a7GRzOmSl3LzuLf9WJvjNBMrAtUl09
X1ZLn/rJtpDVFxRuw2MlGeOcp8v0rfMDtvhw6yc88SE3v6LwwxSjtnG+mFBaYIEaBMXFQtgLVC4G
EANke2T8SMB7KDLV1uujgxOyQP7LDUuWtCM30Rvx4Frz+KN1kpg+a3T+rrlnldah0bJ9JBf6yhkQ
LPgfPvQFBr3UFfahMe7YF1IxQY+yudCC+yNCYjMJxy0aLE5D7E9ak5M5G6NPsYGk03z2ZrLXZDYm
sZsmDuhOg+MO+CeFK7njt6TRDTW7mPELxx56StVaitddW7YH7ROb7WrNWZvCEe3z5HkfFiNvJplq
ZvlBrgI7kGXdHRum1I8nRDIdDIWkXDrCynBSOUWs7yptKUmtku7e42U4cuAviYDVF4CckvUrodOL
Th7hojEBWYJfRZsYu/O4qquinhbaSeWvGH404UjLtKvR8E1Rno7F/ebReeNgvwBQTXwRSNahOeJz
2w5sgIYG8xV8RfumqGnOZFGdgdr2gOn0NsUUjUg2y4jNV+Ilbz6Z6hxID1WxbYCQdK+TwNc019Vu
1VgxF+ClwigSpkQg0/6bOO69PV1f1ogGfWd47RrRc59FqeoqCr9BPjhgcXwbTIG4mxK/7ZgVDkYV
BFgAbeMHqVyiqnijO8JEbNjenF28LUW4ZDxhBmvIoFhFwiHLva6++xNBAZtF1QRl5d4IOAmJYwkc
3Z8rM6o4WXrpY9TFzRC5og/KW//oAWW8ZeOBy/Ab0Tu2sldI33FCWejpWUWy4OkcCWyeUjDG2n1b
gZhT2O5ClWNGGseroP2rW6h86gxumUeE6+qaQ/qQ0llv2UmN3Jll2acoC3DWjDy1GM7ofHvDoQmQ
D5l1nvgN0KeWLlJxKRHV97kOBShhQnVx7KJeSQIY2OVH/8OincywoL9A7Ck8/YMX6AP/s5nWbUCa
Lyx3OEuPbaacD9CUnVndrpYFqLOrOICa4u0gUnDqLY8/LtAicPeHJIPBtGMQHeMR4+e8ycfKWd29
JzYWwYE3GhZK1cPxZjFoQlWjZtWPkIQGRcuVWu2OMSdnsraMbVqVVhQphy6/iywDLIWmegnPI1ra
I4R4dJBy+vB08sNtL9JwkaXuDiONUrQRDUGPW0jbV/oLm1eMCZ9wTxJVNpZ0JgJZDX3QjACvY1Mb
UtZnlpgY9ZrZGnhMJhH9GWCLag7lvXGRHzmZO4dIIq+NAkahiYhUBewVKoE7pr5pyysacTqLij5G
mMmAI0z++Jl3pKws9nzPTKeP7PaL6olFqN1B4Md/z5kJPx1iKxl6wq85ssB26+qYzfm3pPWbv06M
/vYtg61ok0GjIR4S366UTp6jvm7dZfADeSFh8IXLJXOabTPdBTgqvfToNrb7oOJRGTQPOqhKL7rb
5qsWpugh6c4tzexOQBpLs2rQDEz1xESzV/y/7XOFB7HNwdFe+PPu/leReUc5ovnDZjdJ44bOMprd
do4cuPxVeVEctzHL7zypGI2iojYDXiIce10pG6XRm/dhObBuxCXFUhg93SuoYMzWDfHt3rI6n9rG
PFqYwOsXyOjrVOjotCBVW3lZRoGxwD57dAizcDC/gwXgpnqRhC3nu30RfnKFzOZq/boixOytKdKE
YcPbrm4zov7PoXdNyCj127EZn68Ll1pNR4RPTyQmMWE4v187joo79ykhHTwXd92YVqJ261Qt+vnu
ky2RvT+gqGTdy8nbB4vkuUKXVp6vHvZxAZrJwd1EnKcv6fgfCqSm9OSszsEU9qzoc+8jKCg0tKlC
lIfJlodRM93U8nq++xHn3rHPiR5x2T5yesFMwCIqEjwy0h6+8FeokBqCFJdPPIb+1QOYNUVBOuYN
xNS5UwIn6s6UubVal6yDfqoclzp1yzXj6LmWVoiWliaQLw1I31M609MSwiefucWXjYQKQBjDqpS+
Lx3pwyxfoZSeq8kIxD3P4Il4l2b4/I5O+gEp+j4Ed8N9UO43IHdjvwFhWquj33unN5gmX+b4JeB3
wJlFRSSrttEjejkt+nhZiwTWo034w3f2geHdxccP9xVqIqEHDKIOLt849BalcOlMy496sl/Efh7R
PhjwMyDx5+obK8EeoyUxDCjgCAefYxKB7pa0tkr7dpSZPs0H6lo4/qeCvUeh1C7/flhwMRKaDoWb
gsHMZi0+gbtIsTZXjJJrigGD4R+tpk/arJ5y6RCxXcW1OMxIOrF0MebAUWSI5/N6wReGoyv2KP2T
vsyhNcsQvYac9EtiDIajRWKab35bMj90tQnGfz7NrxR1C+XJ7hHsczng/as42EySEhIBn+rkAihp
tZ/6KtK+95dHVcfyaJTJBfjGEmpyEdlj6PVMGBvZeyiadN4MPuyhMLXlAgxxkAmbr5k25V2i2R2v
l4DGeqyPmGflrvghDP6JtOzjDUQNrkGSFu5vFJEyWmXkWtXvIPQeB6H5vgSD9votHbmylkErVgrT
ueoW1LIFd2qpTtXOpHx6MDkI46FA3suwj/SGn9+6ypTioAhID05TENhxD8GaGaUQQOowhKL8DigZ
Pk4eGsPGQR7XZRRQC/JZ+vf2W1eGJXlFrFaJWRwdTmb+JUtWAHrevKn98REL3IZMhg1VaZYkxv9Z
plo4XAPCZFmU1lkVJVpjSb2iw/M28pvR8rCxIO+mos7WkmHTzCNsn2pzAbF6KC0idpIWcuOnbBd6
hCD4FZTqclMPGxjPCGC7fgRRPHCx5v2tq1guIjBn9+KAMBFZdg7QNFoupIM5f0Ns9wbQPHKjC8uY
PCnYKxCJJTkk1K9IqvEuhwR1+9Q5S7iGOnBgsNUuvfX9wYA4CuEJta4T49eQPo3SX3V+G2uFHecd
EMqglpkSi0R9xbYL5MEYOayj37xa6Gha3bfe+MVC6ODqku2Edc+ViWPIiGkQpgw9dIsH6h2D+pBR
ERtpOVZlvMg3sMcbQUSoKpJ3yysWJOBjrhnsx7NDqXLmkCyMqKM8j8PRFpvlTWGSpP7YNsm+mtqW
xSk6RtmAUs3qracmEmNP1HTptpIlHS7mWmSqCgPEksVE+QEcUZWG9rLBM7p2zLePN3MQzhQ76eHN
br/96q7rtVpJiDbm4LoagxxOvtEAu7EWb7zFNqsm2E8nV4StUIjQW74zPJhrLpvoZUyc7zw5gjTI
7MFlVZFGwJtjjqqtf0A6GJgBqyNfOHb1YaKWJBCghHaOQCr6u1nlu9dPa+ChZXuYQw3WXEuxrn7b
1xpjLoTePY1g4JyxCflj6py2j6SUVIJYaK0QwuupPIhoyaIN2fzUynYVMLsoeXhidieuSEyJLPma
vAwNzwU94RHLSNW6P89YeQsA5Oc4jc8hcf+8e9yPDnuOxxQduuIe7sNyM73pf60DJYWQfnAz/jO6
0NSerPlKz9PUhitx/BNXi3iiWrtKj+ZHNousl+LGeiiMVkYqycQItW4H7HVHekdfD/HS0im9uPpc
zRWldPW1/zBOAEZJlwoRBQN6aapequCrRLKlgjlxQiXUl655ve6rlJ+3FM5DdzgZFOlSggQHu2+R
MHPL109JGIlURp0R4RMKr162JkCo9HxcOmjhy/ka01GYvFxn/93q9y8e5ah0xLUnnPxik4R0Pfzq
2u8KLzzGzdAq8vT0FmPjPHkMpOizOsBK1Wk66dHqFPUYTHjvhCwDLxJwMLMqRR6fgognpcpckkrP
bagyMBtmB1okBUX+u/0zdgAJHNnnPH/nhvlAya/r+uTaMiUV//RWaQQCkWJBpWtS3bSFbhgB2T3O
tVvipl5VT1f6cy0WbjfN2ZMGnHg33gIYvT2CqTHaIYW+ft4/K5KgO2A4QvfAzeCQSjG7XoBE7Khl
Ep5SantLaYOMSfdiXj6hECsvk1lBsZlk69czVh63//VfOoRLILTV3A1HunkkWuTPkmY1dmUSJLVb
NgpaUiNb/tgM4gEXH0RZxqJi5MSCIzdFa8TGjPAQNJ2/PP2NxtAgbynhxbhH6vjPpYg8lTLFlmA6
kKX5vhuBLH7BZIPFdOW/AkUvPP1qcPgFa5dUnGs/qo6G3QceVjHf9BnwidpNlAbwoWJOfv77kUOu
dtx08VcLITNKQXfIlZJ3TGCcB0hfM9BvKkA5B5adza1Q3JbgPx84FwqdW8mABkKCZ8MPJiVD7wQ3
IZRU4QUJ15QWVDnjMV7uMQpzFEiCmBJSz36qn+ZpJ4PPoZeQGiMujPkaQc2XMlnCzUI012QKODah
j9nx2PY3xGcrpqOSFegblMNXA/vHIiJ5ZW3Y8V4QzDHx9FsH30UI3bTSpPppwtzD1+db6/yEb8nA
jenqwPIoBThYC/xtmDgJxCT1VQojQvOVpGXY03KiIEdx7eYn5XdHJNPoFQsKWCv5xGs7qshvYY3i
RC/XOjO1VA2vvM4JTwgNFl7YmeVFnWhbiHw8YQJaY5oqAqJQyuY4anRNln9/1RXT/e45DnLJ8S9u
nIsBVOYyFrK7ur5cxkSwr3f+e91tRvQJh+0Fya0O6T/M78hL2nxTt/SKpmbp3cSyZsGMUFJ+jbYb
Ki2cCeAbIkKQlr1yQ3YK3NhORwAT04PTmR9rEqUPdVo4uNrBFykWgSNongoHpJuXRE8/lpAn2zTw
aLhTBGy/P/nlCEBwshqhk6OQL46bVyBKtlgey0VH1HP+Z91m3bjnzbk7PYgS3t0qeFbrd2faKdva
gh0RbHF0+mkfOHAroJRSz/i7siW51TwtAAFZ37xYAQeiNj+VHMw3LFb3KA7YY3kjhUinQPMC8E6y
QUdAYcfpG//2+ZvkLmidXVXQ7IPdpCMbENaOI1AsUIQWXv9MStupOHfATHM23tKTc5mwWcxcGMGo
pUp9kR4jZAc0lS7EeQnTdMIl3hvpD8DvqIboPMtxR3la3ynK7d0jX2XUkAn6L1BOCdBKwwiB6e5j
RwQbHp/79LYAqb0xUnVsss0BCPRsn9SeTINeI/2Uu4jvDTaZTS4BpkW6oHNIu1QNAeS+0futYWhF
0o1GS4xmt2t3gQVwTz4cgyMW/Hxd0qBjm7U79UqSZ+2eIIsgjJkzNFQFlOKsq9RIgfyW6oH3veBB
Qbj3EuhFLgpATd7Z8XWyGlxXAc8YLO6bG/0Va0tWX56U1NovkmPaNzqOuvx3o/FeUVRI8Z4N6G/T
Fe/fJIdBVKDRavlH/yk4TfgkG1BFd2vvXUVcOqZe98obT8cxFKJs3rYSCBHxXobwUVbsJv8cTQQP
lh987OIuT+bo7f3CcQgxo/ab2zB1w7vcEmmN0HsRaKRXcVq9txPN5/0zo7FtB0xjJeN+h5x0bPcu
O2i7/2d62JJro0XaS6ERsUCEeX1s2v93aayikovYvaEYo3sf+MjsxNlXmr8GmC1nmTdl0/Ig+5NA
1wVUk2yD7mhWJpDFPNhCBS7pGX5ngEE8TlT8dTCUGwkleyKaj570njbffTr1Xx5nR+Syx1wsljpw
+6MaMtO3Aw/JWfJ3KtQgI8GJjDEWGAu9aoDgxTKb+ansHB2W8FN3IhXhdQd5T85Fh9P/q66Rn0pu
d1C04ORbPNGVE7tDeXvMb4Y9kMQInHZz4aIjQuaFDE5xkArEuwgsPmruXdj1Dg0tduzIOvNPRW/m
1QBq3t7X7NXxeohCcurA3HTu3IczcXx5VmYxK9JcyMunO/q0l7setRPgshYYPR+YqHMVzeT4jr1p
5PPmJjy6/Nstz7luUEAU+vbOwZh38fKv2g8jcxuSFIEvUST4Cx3di/KmREQhsZ82poT3Lh1sb144
Zjjx/fU33hoskG7L+K3NnzfxhfdAyXKH/iKJOVvB0sslnY67YybupQ1Ju6x8b7cgwiG1OL92rX/w
C01lz80wDqkvl8Yw7MIfWpfdCQAmJvJzEnpacYTfixa8IFSgMb4ZtQFC+4cufXL2lzMedM18jACY
dSCMPGtpkeU54OkUGP7kmmojXb978QZNPPi4+L5ZqCi0OQONJIvMT9cCyGvE2rTsrmHE5EQh70A5
BaV/DRKs7IYjLId70JWFr+UPKcfPXh2HfR8ASixLJr1tHkfux0/2DXUD1G1nRg4eqIWbjISYUM2V
mrPytZvSfT9JYiZs05zd3v9hTOdFS2cpG8e0gXEMkd069y3GyeFd9+NrDtGrpIA1NJNAMOqmfEpH
YY2ExdPu2KotgNbGAUraDu5lRFoaeESMSwfhNKs9f0NsB5hLquHYKFWnYBVLkTxEyPHNi4N5GHow
TgZrskoxeKik9dePkasIf7cMuVEM+e3P93F3yH8QKdl2y6bVS8X62e4Tvd4O36X4pO7WNC2jI6ne
9heLSrbSSotTb0i8Tsvd4vWlNbCewElyiwcNWe1RUoEojz5ErXpsuhHzWfgdUz4OTP66/SFwTznZ
t4u3ehd+M7Ga4nsNlPlI6jKerFzcydOmkAx71dNvPQd4P5ap51Pdk8OnvPKR4RMwNmLXARJ6GtDU
kn/pLS1r3I1o+plOHTXWU4vFvjVyf2ap9vGGk6Ebai7WSRR6RI39UswcJre9qLOSXjaNyOPFUDLl
NgOmEXHGEZ22IZz2ynpf/oX8/rK1oXIpCalDVDD0T945ya8zcpyVZDBso54EruLEo8jf1trB9p/W
JCMXV4/aFDEw3/ukf23IKfggjOfDOjFDj9gkg5EZ8OHeFUzvZBPDy76CeB0ujG8kutXXQXmAXN5D
qfz8Cg+PgtGNLwBkdzXhMzotV2pm3j0gyKeEc7AMP32cD7GyUagzJXQXmhIe1BCqLfjqGx5ffkAg
ho3MVtUd8G4DyPev35LE2Ji+GgwcKUnPj3Gcsh5hBYaB9x1/3yqfVkAjr6W/lqJElcPaeTKlDiAS
oBfBKiUPStpDAlrvSHlqr5F2W07xC9J0JG1XJtnpW9zO6NojIvHu8YdrLAfeBVCEsifTNeCGIbGD
v8shclunORD7jhJxfqjUD3n7YF/eJaZMUz3IhERS9MaCRlNolKySMhV31vnMcFc8GZlYSW7LBzUF
CdZRfCdvN4Ispw/wL94aI00lqN1/xTbrF5wlM4lofQRzzcz7FbNbr1vMcuKgNLpYHP1f+FYgI98m
5MMLDoGKX5cpnhd0YM4NN6cGv5ZSg8Hvu9/FiLwtV1q9qiUE3bgDXvbIIXYlBTHeHpS4gOENLZlE
4KJ1kYDLtJk+5FTVzyJWZjcapk8huEG93cgBwSJQwVLRMR/AVrmVrEv5nSVI+9B9OM3SzVTFsMbI
I3XP/7a0f0CyJhBo0kw4oqISvXPjvK68ElT7eyXgJpFJDcYG3Z5OqvaJEAOO/ZSWpcqCs+5XQEin
v4lZ2CkQ80aMkZg+uHyEqDciJ9PwypefT6RO1ZS/9k2kPe+RVuJR5z7+LtRnpfwf2sxb+hM5+54x
jWvClpDqLO3ou1OyFXWf00Dc1g9LXrnsxlz5LRHRBrXdzR6JPMuvMTqFJ6n6NC6ktj5hP3aMQ3Yz
w/g57jmLen2gG8M5H+P5HCKSX7SCtjcHTh0o4ztDmMqryri0l3c3J24dcw99LBPyduboRhkVkR9+
zhWLdA/MasUmHXrY0Gd3m0hzdtCPWgFqrS2SLPl8Nk4hxO/AbWjwwl5ytyqISpLmKTxXMQpWaIPN
8EVtiOOcQio2z6ejozyHe0oLB3GQfP06QI/B93FZkZINHpamsQuk0xnSHsJDYZiCwzZbcgh+84GY
nTyh+mE+fqf+Ki6Tyw4m/5h9dotHwcQ5XpPp6ckGG5pRfDd6JihV0/n3HEo4031aTE7CZMB5UMTz
HBSpkGPdvN5MdQHrYfyn5C69bqySAEnnZsmjhpAouy4it9GhcqjSf0KlglJj7ZJb+oEubiOwQDO2
qDdGE5SgjEwpdhjnNFf75wi3aeRATRyuc9uK7z/pt2bR/DoBfM+1sD8sbYzz4jDvAs6sfCf0FpTt
+WcxeSc44Z1v0rM20FspO1D5FEiDsiKleIq7HMLfb3fhfmhK6guc2i39fxGNuDoXwsUz6ovtGdYT
jQRhBTIvQn2ik5mcGR7vfWKFiu6uKnxK74UENLgXap8/ucq19VG9Fpkn119ZwLfY85UPfxzGh/ux
aK7w7Ycwqf9rT8cejxhwXc6KTOHXumfT9R7pLBKAQVeGejx8bjiuycF0yP/D36oVSSKYarZPoDYM
c7jrfnFeP8GxQ7o2WMS6dRRe96E78L0Q1Md5x/x/bHmx0c5I62aQoPQKqmdwd/mFKmATzjGphxFr
jUM7a+wcKF3FQbhrjykbb/EBp8kCJlr/+jPPBnG40DyxhjhP9sAR9DQXczDD0/a2GTn/Av71kjAL
tvx7P5JQXdzqLvYWGzUv9f+pMFHdILo9Os4cFWXhPqNbm7QP88VOe2YIyYD9612/XQJLjJg3A/ds
ymXFi8BP4SwQtpNe7AH51zdqZV3/uk8+uOUN+qSECcvLyn1lkI3Ic14Fc1NHLe73JrWAwOBIMrAE
lDwEdG1alGKICKwlQIjclD8barvDYcuAj1SDhgG0JXUa3e45vaR3KEgNBPMFRldNbGm9X3jA5/re
YODfH/gX4jso4eHGNSQo7dam9UlLFmX82BHhhte2fW6PTx+msofTfFhAmQWMm1sfjXtC8EJ+LBZF
GTixTfiZEtB6oACUcAl6GgPoHTa0tqvoirrj0spNolhE/hzHpuMyXvt7kFn03Bag/9Dqm8qCDekL
B2B4FwNwqAQghOnaCmm+bzQD6skPUFG/2daLr1o4akbiqLAVoNisPEBqbjbkPvcQ87T1jSkqFtHw
l73fvSMuQmFUpf0xJTwydEmS/5EAuZhHkSoqMg9vgguDgHSbSYaRUjZRXSqYZgSB/cOl7mI+IyDo
PPxAKOrJy7OHOJV4xueaQIGZGgXvvjtWXHEfxIQqJNa3b6nRPrkfZZhVRccEy5iss1ZDdb0+gO9j
x0FppELwILc47uw4YHsHwBTxDJo3FAa5iNKbiTkvKxg+TbsWrWYcOajy2B4gEfXuJtlITWAW0l07
x6FoqkxnfzqIq4tXFJWiZhd+C5JzISfnt3FRLElb4vOcV+101sl/hmIlw4MWhuuKQnvo6GSIUq+Q
gKEXbGaHcNFl00r+0K7kTOHnVq5cACJV9v7S9XSDFklLaAsgxj12JzLiTP9bSpeoYCkrly8OEmpj
GBVP9FYS2UBtcZYoZAROqY52RmUeLmK3d59MpaWC72NJ4Sns7OLYuQuneFB5+OOvYMriFiXCRymn
Ui3zUyp6nKSjfZT8LOS6xmqxpW9l54Pj3Xpp9FleIpOsf0+xgFmMQsPMryiL/dxSeUkjqrtDscns
9eLl9jCnJ5zmhKk/lM7Ik+WzjFXJajXCVJ/AHumu8WnEOCog+0Z07V1sca90+J0hrHSrNaWxpzuk
4LkzacW54xhaN3ruNmn8IETxUZy0gx6CfcDkD/ehbXMIaP4b01QkRNWr1DszliO64S+w3C4ZWcty
APaW3lidZZwRgbssmobkqoOJCIvAxE88AdgGr2rVkkmDpEQ5WsRirZNe5bwcq/ZcJvganXZAlnGY
HkXuoPW7KbtFIzL/eylYMuvwu0sr3FaWmyAHNa149zKQ2WWXyfF8/hMKPfVDwgZ/+wnRM6SRinDF
p4c+CfJmf139wyqohYeOB3xWIRnSrkYODgycybxBET9RmRnI2Ka3nNc8SLhHk7+wDWoG1gbcuMKI
Oci+nTEiH71M6xGK/qDXoGODkXvwKHeJ6Osza0EU+xnlVuqshlAdYwGArFotZGBAmZZW4RK6/Gd9
a/alTKdcbx6ASW+Cw6cH2sTe4UiU8sXT0wmqq5LJmHS3aMmM9OJP2BzPqSqg+40cEk7VOu8RxIso
a+ev1K8mVniGRYajVEL6HGs9oHjviWAdB+C7Cae8qR8B8Vzw52/8vALKrA6xQ7AuQJ9cqg+4W0A1
bp82TywcAkKKFbMUP844FRQZb+esyrPm+CPK+UD/0izwBcbKtDxT539Z/OzGMf7einp5lkqEOIf4
BXYIm57c7e7ZhcuZaBNCJDV5U1jjK0I15SkGSEXWSst2cbveAuuKFNm0l9QZN0AoRefyhmgnGCHa
eN5SQK3s5KVNI0WBNaXySuz64vfpEhObKyoD1SNIMX3YY++5oc5+g24OGuyjpWLyoeNcpSQ/FJ/Q
Idgflj5UsremHOKsZxr89qu+mUa6pmvixRIVkF9Soe5+5ma/oa/OQZh1FRO5TW9JKrwMqvHxryoG
HhxfPHMJvKaDtPOL7+AaiQhSkEjjUDDbbK8n2NAPoJ/HUvR/bOd8mOdYQZsgET5DICIrloG5pDh8
ICGUs/WcwJeAdaT/RgLgl5IQGtBi5jbtgxVwVcYjHwo8ObBDMuC3MV1u+apHrZaA5oM9pUKXVbqi
2aziw5KRCd7Eya21DZO4LgTo5ycakWQ7oMDKJopVLCY2fUr5WqCtLxAn6jYyBajNQGmPlwWAB6Tf
M0BxpV5mRg+iK7/AEJ0O93tVf+28T27bT6rcdSkHyDJw+2hW2upl8QcAnsdYHM9gtTlCf7HCHnvo
QESXmfwBAJbskkGeQ4AKi8KhrFZC0dDTghSMFfMvlvC3WLPIUb9+ZEMndHb5PkhuAOu3+l2zD7zD
42lC8I3zu1jkiww2/gAb39+umne2nKrUiOHikFNp04S4C5EHDpWjGDiGoKUtdLd7M8tuEhhDm1ay
Tk4yPolG11g6RjIpMpeB77MCGpu8Ixa2uh/peXW2HCSsofjV/DqE0ctYMZPNl+2AJ61vFvkChuVD
BDeJVuLH6e5q4zMW4krdPlVkG6Q1s9f4wZr5xHsFroPlO6ra0EAmmT25MAuyIzhLzlTlsfeGbM1H
NR+eIiuHvMxryvtX6ZEGopU5WzOx+d8ucFEuM+SchlDpbLs/Tw2UNAo5PPdYnNiM91qAhplPO0ry
WPBTiHp3sAnfxNuWnXflH9apH8FYNGR/hYEV8yvJSfyQCENMyzmw9mKMXsdPhLTlXSqru0132Jb+
zuhZiAmDlB9lPUQ4ZuR7MDXAzJBPHT+U1vj5VzS6PVWzBnNQiLOvt+T4yqbu0izCx6UpS2zYXs/X
U8j0XsCtvufGoU4tYtf9FfPmQalZxKsMp6NgpxR3mBuw6o95WscyRN0mpjjDO+RNReQmHj7m7EKD
KobHYvtKi0bN8hOcXpRiEC0hQgl0ZOndQMcEqT8agzUTQSf0L4wMcXWPR9yBRasnU3TekAgUMsYX
GymALMHgy4epYoHCp5ynuroaUwQP2YQ0nnaLis54sfDwo6wOyfTcr25/PCjLHOYZaLitFmxdjVvk
ljpzpfO+Tfh6sH2q4I/UXingTpiVmf5BNBAWUZvODLeQG7fCjclmEM9fALi8kiTjYXyMTv+KCV/8
acAVH7gBLon4SdLtQKSQrlUrk+0rbpY0vuxRqA4vgL4gXgSG46AYwK7YTZdlUj5LO3TbZQDQLP0B
POt5VHedZdPkw/Sh8RsIKXhWzcYLNKxbP0T2c56ptaYYqY8Ut9wJ5fRCuodqySwtK9KRVHWqww1+
6W9C/Rb85uT/l9KpS8KxSy/wjtgx/6ZD8JaD3DXnk4VbrH+azUWUk1831zzswRA4cIImt3THpxtQ
uMkuxgvjzqzg2+02lyDu84jkxYr2NsxjOrqOueTIgN857ZYrfe0CtD8LIsY0uZWRnutaqQb7PoTZ
ZcOoY6oEuj1svjSZUhY26wDmuGwSnOOf29qlmTzEQJfe0NFfopFWBW2YKxya9Roatw8N2IyoizO0
Btbi7DCov5d7YLNz+ISGciQ7hYHx/c3Daewwo2nzZXXUPiSFPtUnGBM80FtPltfTBNcjiKHdwgdl
AJUc9eTcGBExrLdxH14SUTcgJrPMNxEfyNDcwQUf3IBJJDXuQDAvOembmmkYEj0+wiAcZcKlqtkq
MtuNiivNuj9T3781+yNTOxathu8hbxHXB2ov7MXyrNZZLFTBE27Fmbecw+YJGxn8RwbL1+YrGkUp
qpG56dMDfZqXlBfyoZePqHCJESa/7s9d6+ncJnAxf9fFFK4ZnhqPW52bndNhfg3BTXsc869X5aS6
52th8I9IAkgrCr23tbVtKNmMa153nArsHTZy41aDMA5tPymGeYmw/u642K8Ov7DsDHFz2Dug5lMU
+CD+q4wA/bJ1oGUg6p7+ECIj6B/oe15wz/Q8rsARipvBcqirwS1vyOMec58f7+PNREe6dEvb77jk
3sBD6lOsjC72o0/VSZWimAZPJNPCiIrJK595O9zn4eJAroWvAaN6EWMWQa8WOmvA1vCPa55zTbWU
8WM3fPS3eASxbgWeeuqiQ7WCe0JQNaJqnMyEyrb4iD6ve3/+E2P7Wie9EmtmOzV50PZSETDNPkZT
Cd9L/gPb+Ryejov+VyGzCvBZ+ohLp36tlGofpUyEvF6KKRXXRGssC1ZdGPp5tTIXsAfQHXm+8u6b
Qh2yWzWnWkq7wkKrDYEWXxhPbVZRHu6LGgErP5/O6spYuzjdPXmJaSFPiFIuuyikTjueRhw+x9LK
nifhqjh+AW6K6s/w2jX6Hg1wNZIk54mOEerKNcS3JjqvtR0GlaKPMOx7A0/5lCT5tdRrTm+9D6ds
mdUrgoVMcHgV7TP/s+IqEIjv7Ooi4v35bciO4g3vkz8E3G8v3eDr6g8KiPZIvsN7ujVbDLgJyuIp
ugDcYHX9r0oEB8NlTliMvSa7h97YiEjD+wh2SNQtRzWRiBMp+ezlhxS/20092McI+u8oifvVS/7A
7RG/acghJavVFreym7XdkUH+0DcaYkAn+Gq6LAgeSGNxavvxhJynhvwBDD9mwKzeGEun/XIxVJ+X
7hUUeiHVqjK31XE2d9BS0Umg6I43JsEs4bdDmZg083X1R228P55yHBzTDbzC7//s0SY9/iK224KR
aSxIe58LdraOem71TR1nEGR6Pt9y+++sbor5kLhRdQCbtbLZ+GbnJ2adjrs5bmjbpiB9JFW9GLAB
PlljfGQK9W+6PbOX1KCkHFTfpRxpG2cQrT7WsRXJl815t/+0WPjkZqh/9MNdIXPNb/Sgw/AzwOXu
E0qILWtx3ZVvq3WENe5zJU4nnOzO71SJW6IQQRnB17ju18XBro2PV3JN/SB16GUeUcZFOPVseTT7
EQAspcyQ6Rkdu11mZCag1ZCrBo63tdFUCKbMOrfLV0RWyjCjAK9MeXLCQIAmU60MOJplKPuvw7mj
XDT+nE5ueLXd3CQ+ncvb4/RdUC5FqFsnc7gjh0mzpiTO1W+kA1mfJMkQa6OihVXtjqwSgfADnBHO
k9ieqHSPXfD7ex3oN3Q1BicJP/imi7puIU98TrGW7lrWdSSDuYhZGcD7a8xaezSAP8PQbRWFOEGr
KL4DegE+1a4CNTgCnoFjp9JBzWjgMXK/FPoWqN3vpknJ3xbDtMn6FICwu2Jo3R8Vf8DUauiyoLem
TekkgvylPlO2x8xKK/xn5CyEpSFjCcnqMMsqwPqefwR9Rm/dWiC/9LcECoGcLofCmSeL/ANlE3fI
k8yEtR9miNf+zfwbdU5MaEZANYDVGVZgfMpXznVLifYh/2IG93IDHCD98YiLmaj4Io9XxdxPy49h
0EdkEV+L0zGjHtc4yqcbh8mHEE2FFYL0CCQmsIlOm4094Rh2QNwdDU7olZzzIRTEBMC20EBmE37Q
BOZjOPVOtVz2oznjYOqSoW9Ul5gBwrRHSFLkb6BoAZef+BRnsKZSCueid0V95MhUjwCwAHD/YOdu
3Qu+l0M5hTT4doZlx6WJqqD0OmuMWrom0QZNSzO49ox87LN0RPTCq5lWLKBowc7lT1UvxaOqVHRx
JPzaH20Sp8ERAzjzvxfBeDi7A2C45c3dijd5Rt8Gb8nrjm9cNdgjCJPPxc/lbTqqLSmWZjsQkYr2
0YKwqfGToEZdE2fPFwEum0gkKwHw479pMe8ct1QTjKVMlhYNcEZt8uJvN91WYfxnU3c3EDy0xSyG
sR+zYKJxFPfjFvxc2/MEYoHlRhg4IwbSwqpvTL5duiSpauCm+BTeXdyMi7MG8Y336vBgnDFG/Ir7
DxtNgqVpsZGo6fwPbvFWs68+y9zqhjduoPHwKT/d3DAWV5eqRPwIds8j2I2no8iyLIuplRZSYCgg
MO6dO6dApWEvmf6oi4oXzhFIXsgRAWks1BQijyPFrX3oDi6C5P06vUW5/S+oBG4F9lh/fCwlu+IN
BQY/JNDVt88zFnbnuRQf1KHi5MaDftJ/INIFzbTvrvDXmbu0GmvTv+I1i4v1Bev8SdiS8qbP3mmu
C/5W6eVrTtprbJNx1cgPNLqt4VmKe8Bq5prTA3pdUc0vF5GEjlGbEejfRgZj5QNePk6089jsEMpv
1JiJQCwss0Vog4Ko7JPJo3Wisza1W1CEPPSQhfjHkepVXRLGsdn5MHG3GCx4keIwlp3TQb0oZzvc
pmnb4oGOGRqHnUAzm5GeWmjPERVszP2iquwJ3PSvVkUxK8fskLEo5Lw58E/fn/VkYMsVT7W8tnRv
pJOAfBdhrzGIci1xF5Lr4knHCoi9X8r2rOWn53lYQ9G5GbW44m8My6n25jBGHVCPlR6lMYkFDw5I
F7Y1sZxL1+WQhT1jhfBJPfzrpk7L8jVDak2FhYlNokA2sByg0ij9k4h+A5R736nGOEgzda2GwXDz
HoKilPbPtVEQg1xB8Ue6F+QoGsF6ifIZN9dMbdUrq0qmOBlxc45gxxLY988JhKbiQp1q9WH1hn0w
RFLDtk+P8ds4aJ5TrQ4Xa6w9xwDRXmBUeSmoCCOQZGgxXizq5svHF7PacPfdnRh9yz8ft/nFwzQr
YvpY1dSPLqDd9uQ7L7xXA0k2iN9nFlNyIBz35Iy5N98ozluTRLe4q2XYUnDPALyhntWzU8/sBDXm
pqgoI8zl2BpRWBUndGpJmQu904nXpfLRO/sWm+fHqdf4SgHnwvrqi0OMplFKTn73UUEoZOhufpji
Os+YZY+LExtsKWeWTUsgBWsdVqed0SEkD+eFDuAepi2WCIWRKOrH1c1HUsfvK27er9cYdCc2qHct
QCcdN50KNTx1U3/udNXSWzLcru7vH8GDQfnj4ZT/f+sS1DwDRZZDhFi2t2QlSS3xTYr3ppYLWSYw
1qFST9lX6SXQNVczofTzylfFZoJZRV3ovUlwaZuzu9QYr4xBjZW3Q4VxDLVr/2HPW7S8rrupi2I/
L86oaMGjzamLoc2sIRSbporvFjWoU4pgDObqsldHKzdb+4L3HIkLz7jDi2eVad1A1r+El45B1+Mk
UaPOb1WAw4rYzf2GHcrbT1Zhfwog27g5PFsizm1MtsPDvYczv7/5gAuQrBCbGkZ/Du0m4k/40af5
9aHsDNNS9INwDFviu8mJx5HrdssH5i66Je3BmT8BpbdEWA+U4ZE4/MMedOTFauW2FPHXk0mpu3Js
5/YGZFrXgQ2T2pXomRhfYHTtyf0Xsng3kicrRmKcbm6w4Ocf4SPm+Q6Pehv7hCjr5I7ER/RLrNg0
mR4qPp8UuIxFlNvPhHtxY5jiHgMZaVs7pzVvsUhjv1rgrXL8+Rb6LVg3dTJWYACP+s9B8Aji5H6d
VqOdIPn2k0kiEUsQBI/2Ik0aguNrRg7qd+K6BCGmGddWmZvQiMHPnCtLPJv22gt0C+P3dleMBSwm
C3arWH+oxhtTKjhhx4Ekl9qP3yYbAQ+RiNRpncXXtVgGmVv9x9ciSusmU3zfnIJ4eYgMM0RmN3wz
79CiW+4v7+NZXOw0B8L4du4D7x3RRZGfUnGsCJEdzVCkmtS5yFkQoMjhH2KDRWfLhEkOJZI2Yooq
4FOu47EiyF5uV2DBcu21//dNiFF2wmGIMVr7dfqFdDhDXi4PWjxsrCVBWhNSE5YwsEYzcQ8HeHuy
DO+pJHSpndZ+EOAFUXjdn3NwAWE6tUCXj4+eDXAhNZRS4bNCEaOA3YWlwnCzRvn3mGT4tlCMHwzO
DjzslaD7I+bdrg05xTyN++zeUezwa1SKNGngEIAtDoPAiRrM744HE0EswJEOj82Qc/2LMsUhzilt
Ouc4TnqTzse8j7Y/w2cjhh40gwA7HYv5rD5sIOGldED62gb9/pM4j8OkUwx37OBoDin9u5F3pGx9
cEY68pswErxxja3mlVI0MGBoS6uSIsH0eyyykZDPmxl3P2XYeKBklr05deMuEIjCjwE1+ZgtjP8Y
Zrhn17i4rYNEXbmh3nrhBOzXMM6hvZruBN2Rk664JsYrTu1VN86J8HZMygwBWXL2ooPpl/542SEL
ZG92ozsNl4udFwGlaIlSpcVF4nu0uqUQipP8m/l+RC7VtQWN+he/QNhAA1Tu2Upvwn+7a63XP7b4
jsyZtxmdFAQ01CK9axZmyntg4oFeXev8SuRs+Mcned9U5TnzOLaSafjaHZqjXEk0ZrJjCfLV/Abu
ODSCygQMuWgNcjxVFsAoFn0P+OqCh5jllhJ59lXuHOeZThUh/Pndhe/AUqn+Tgm95K67ks8DkEiY
x+BpI6Ajt7RUBLRFiQlHVjipaU91vKLw8cGoU/NCZ+4hI7NORTnCoV22WLWtDI7FbktKdW2kivkX
Lhc7LhTJwEV58dwkkRuI3SlcokxLoSom3Ek/v3GS9dZuB8UpfuaoAjXAGrdKnPsyAWQE8aPsVGCI
Ge3lfrQiS9YhaOzN9PkuNJBwrmFfZX5BCdxRoG9eJXuXqbu6OjS/1eBTuRuKQi1cJ5rGbpDqF9I6
8XVLG+EIyckFCcDp8KBzLPho6lDHbSGFIRvvRpn+gFxzvynglI2ImTB4x/jebu/w4RHL21+2fYgL
YtJ0EXFeAI8uMvJTV27Xa6a6A2+qYgqa6bxKhvaSK8MpHXLSogAY7D0uxkUFGIL2sr/EO8zZbv6U
02+Fe3f13d0g0hME0Hxd9aV1fz1AktTObadY2Hc+c7RrCMhK6EfDQpQr2U1NDX9lpe+HetTzmFJx
J9Ye8JJB4O6oPn02xrjbqiM/hKTDytJkM3YtXVvEEUn5BVNE36Hx/ne8gqT6DXpoD3gagHzRG4ni
jj9lMw/d8ypFHiDM/t5+aEjx267j7SRKQjeK68I/6Xa/fhl1ho3Ja94oZPpgYtynHS0ClLs71nBu
I11tDbgNfw+YIYPMqeUaBTIYkhljCQV94/MP3ObqF9Mu21EvjBfxpqYXxwRFmPkoU+M72wwGp8va
A7ObJxMH+CrKsukVwqSn2zDguVtLzpWdBBLAiM4n3jFoqEj51jaGDXgMZNmSTgSISaCLGG2khdAW
Qna3Szk81sjn6xvUYJ2WIhxWkfSOHfEhcGobla24up/z9E78g4m5Y65vQVDX/f+X9qNzOKilND/y
vfRgcmzE/Y0fHCFegf+s2w5iLoTb3Qi3xzB5NjOfZmP3HZlDifxsl3Jk3gP93ljEu16dW8pcjzsO
OsW4XRRIQfm17beet9j4NPTzdFWcu9ihBpV62o4W4GfIloIPtNRdhB+0oYD/m2Nl4nwlioMpNLqO
yljYa3hma+8Lr/7vFUviCgC5O3DIKCuzUvInQX3mp+RwJ3ebnx1ewDCbSCLQ5pzIe9IACWOAs2pL
THcusQZ6waARS/POM1hmhzQ6obi017R/OQw2z6pbj4lPiN7hWGi96EJOv/maCYEdgfmio8gaAlSB
FG0u2PGrwUrDxpDU0aoedKbQaGpuZe6l4u4AVF7KpShuZGMn0mk39a8wDs8Ppo3msmRmAkSO0ipp
euarYLR4Pq4/vrnZ0UGpe4hsFYc+Dh6c1Rz1r6NxHhdGRTqJytkukkslL8lxO9RX7r06hKfajsmW
5H2xLGWU2EyTrNBe0Wex2O13VWvo0sgQihQegf4ykUlvSkZ2f5e69vQyEuMq1yvZM3PcVAzn7Ybq
qIOusG5I2r59TvwEMgUpMqLadKMX+WVRIadudsc4Qy39fhywA+oQhU3dXF4LNfiCZ1Q+PZjNdUU1
DTBQ5r3JXUZ4IV2M6CQriRw1zxtVdgt11hgj8iKjjEMwgvyL5h0O9p2nhaNTQsPUZM2e+Chp8e7t
heRt/ZMQD+WOXOVBvCCkHrKuYajIlZVrAN+UHqgDpX+j7PQHt7t8PJHWhp2Wd5KOdW9cbczIbWzH
VTpkSu6e9IfuV71qlS7wX/70F2fLOSsd+6JSiB2789K29yvUhSQ4MfAr2SdhcRWTeptmn0tfnYPV
6QNTjBWcW6woabPAR/Z+LsUlCr65wjj23H1HfUZUu6qec+stEl0RvyyewzSt3nz3K8iGtKYtTUry
eD4GixzSI+x2ZXmB0hVg/DJQpl6MSTqdJbEsovnzjAIfp1Zb+d1Yj2bnMwWRFashgI3eRRAikD/c
3qgC7tonR8yFGUCE70bdcZszwZ7qsGSa11DE7GMmyBHIjgq+y7b83N2D0cVfumKszqPNVZ1BnAME
mTuPaJ30ScgXthwExZQrAm4H5C8d++lX39eWwsf2X4Kk2tvqeRgP+ufw1uMzvZKBpwAMtS/foakz
g4hhZK+trn3X4V8m3tphDjAynZEIR2Jtl73yAFwK7WdGd4hIlQlI7fm9aIsc6YUBMn80j/BWi++9
mUyHApoHiny3kvm47+a1YCeeUkctiVbKJrOovSKR3f0FL/RN1UBRenUx+43ZZrePm5vjnpZM6v6d
P4HQhSt5NEgfRqABFxjCinHns2S3/X5Bd4996tO1A52COxi+fstEroZl4YTPY/T/71bWJWrmxRsi
AYgIhGJiGghlwuCBLopfr9ETG+xQ03ONcH1boWrchf5FxrDdZVMtChco0O5iJ+4r91FyfCDsRc1W
oUQOgTD1zeLc/hfI94Iwf2MSa1j451Xf76ZNpdpvm92pG0yWa6Zz/jOOawYm0HT9pHN9riAvMZKr
lzxwgNcPvipDmKDEBup+5E7bKLAvqiYo9CtYv+q3AZMZ8D0PdGvN23+zVUZSkIqG1y+iEyPno2W8
djsYly8NZD91Z5JXe02JBPdYyG2yHyXJ8HpLcYrPE6KwWU5S5NIDKJqDd9Zo1yiEE628NyBQ5cWO
hzyWcu3lFrroI+g3j3M5smn12401ANVByp71r4Lbw1jOszY8g8Mrwab5brC6gTLij1a8Xq9xkWoI
k07Ms7V57AQEr1bCtaD/2skFe8StGAUztx/hIapiPRFd38L+xSFxUO3rc43NuwUYRAX3smOUNFkG
p4d4u53zTuAuDBBHeYYJvhzvF8oT/xHDX14QXzNfxsbZInq/vhg02npWS+nSlOT40q4aZ957rAs2
TGcrInZR2/ewtECEN+MuW9TRZuPM6lepuCvx7bZ95Cm9MZGcFZuhgEDrt/DFqTUVzUpa1Yt3xA0F
PHHq1qBzo2xKnkzEpcq2C7dAte1dl72uZO9styIDmj01PdWR3dvUhKepMEPE1peQBIBABP3e0tiM
PugdCzwWI1Wr+PLj3j9bJ0Ys7czPgWN5tPq4LVFlfqR+S9qJ0Xy6Z6q6zKlLDWTvoVx6q9YmmBRS
i4ZfbUvo0xLg3nP5Bp9ugeXJ0cUoGSryOypq4gTvjnXBbIuo/Q5aSAjgnOoeCRFprPTZj2TU0Ckr
2vO2MdeawQByNBodCTvc0zBxL7AiKfqwA0RACo9+zas8MA7dBOjRgaZImIdFHNH0MSj4LTtTjAeC
VherF2l16yYoNRo9YTFNDAZVMjfSYFHyYHO/K3YlRgruFfR0Rf/beKZwLDTvXMHismbOZwhITrrY
ZB98qq8+QT5PXtbYAxbCiP8yHSeDoUI4APyx5cnyBbQHzW8xE7qULVDrbKm5gZ+FiMIcD/jq532o
sExB9Kl/Dgksc578NO1Cy/pyXp5eCF/Yfnr360AJGeU6tdW1x1BC0g3L6xkApHY1mYj97BCbD3vL
2IWDlwSrtpBVmbXNPwRLdDfK9LXYUtAGtZ3xt8S7ZSOEIuaeb97NnQ/wT2xRPTkdFOdIiuo26D7Q
uB7QlSvPG6EnainOZIiud20KNSQtYzon2IFtwFN5niWkMLnF3K0wI1/fr589AX9NuIf4tb+fNlBA
ceUMwGjvVatrVnpMIVEBqYHjMeYVN43lKit57FlHho92Esx+G4h7RCOwX58dkWz3C01bpDBqW6/3
QzAzleXmtD7S39q8cuidVTH1Z/Ax8LhpW9cc97lU96uWf+KuuIZVAivOSQrtSmUZ6CiYygj1TU8U
H7bzAXSsVgNrl+uLDsL4qkFr0IWTbQgNM2UPdgflJCJz4YGJFwCVhzm8l+X3FJrsfrZWfFL2x29B
w4p1PjwcS1YKiuq3qZKe2nGTyFqeac4p80g/h2M7wSAWtOkONAr5SXB8DweFrLx6WPkponVsSV7i
B+HiV3473stQFLZ4YKVBcPLkCTt1kHU4op+CizFVzwbPiNWOvn3dC74zIpDnNj7T9NjWPdTkoQ0r
Zy2qAqIGz8+bk3fH7osSqVfXpjo16iJ2wGSYImWxxzFxKxhGwqV6s5q50ATYf5FicCH6Em7IFvq/
MAVYMsSEtJkCBq75EACsVUopcaceN0Sv//zuSJnmd53xnFxfMF1J9TXsCkLDT9RpNsZfIRrndpWP
Q09CrTcLzF2/LXrW0mjXEJ9DdG60gbjlCftp9z06JtRGZh/s6V6hlQaR6VHB6XT7TlHDSeX+C2RN
v78gMy4WFadTkgpthzO7cadfeaARx8k6knJ8b39TQXv545rP7F9Py0GU+D8drBsWXyM5x0KihjSL
hxj17l4+maLTeN5SZAb+s5ErPOm2fxCC8tnU3zUPxQMxhVaioX+kz67Edb+YKSNZOCCpQ3/zebVr
ap0ivAdzVFm0mfWo9BqGJoVY7Sx74rTR+AoXW/oPNUyZSaUN3RTnOzUp6xZj3MOGOXDSDHzpAeTT
y+zTpN9P/V1CTQQ3JY8MIV1PBe2I8j3I+Zwi6Qi8qczyyJjXsJtqk/2veIh/JAPlU/YY2JToaGbr
wVWXbU11gAlS3ECJ12bo9gIUjqj16tAO704V2WPEgy++m25E4EUpYz1V/UURMFh4pEC/bch/M4C+
cA8h9TGpL3DTzK9UfHBKeOsmixRXDErvo5JylFAQLYC65JnLbO0oBEDredtkp5x1fphV/ozMEo8T
cJ2Yzp9nFamUul4CHlWNEqcihb2GOX7UPB5Xr7upoquSmOC0KOQ+ilVXhtkFl70GAuy2p88lwMo3
EU7V/75+wDfuZCpSTGGULdqmSuDJ+S6hr4pWW0WVEAY5GWgidYl8kHXnIUIQWQrm0uav601IC2DG
ivJ2waqfmcL1iu+OblRH1NKvMCn6Ne568AzwAYSU2trC5SltJL9SVrsy/SO9V3qv/Wwl46MOtNpM
hwS/NLK0J8hqfjWlTLQybvhKs3CMmiZVqpQ2qZoVEpqDzIjVDq5fmV0F5KAvNXlxnz+/Jouf7sLM
L8p66PpODuPjN3o1J4DyUOzyuE8kFVtNwrpWf/apkZxZlcc7faIhKEyOdOkSboy3JPIKY62F2bOK
bSOPIBKuaTfFuITedWUW0eiqUhcHxbKmxMLWRGenoV6wt1Dtu2q8mX1QnRG6YyTMEfOq8E9XpEuG
lEs8Y5ufgTG6Z7saDL1uDscbyo1fsyU5puXP42612AxzoK/y+cSGT0bR2XQhxOnpu6MLFX6Be6gL
lJo4D+gYNVWr2YFwVNeJRTkzXeSqsWfxcRcwxAycYeeb+OnAfx5PplwfHJIhR1BYoMICOHrf4uv7
ekTR4lhV4wAU4ikruph2KURsWWWMB+PjjUsMIMDnSaFE0tRHs/3IN54vu7MgKWj8tieOqTtvPFF1
sUw/wKRFr08fgRE+phBgJeoJ+3drWjzRTyRseqVFq6dZyc4EeKNFKVQTcnlI4Ie1Mb7IqmgvCXSA
Va6oWcMD9FxN6a9WYDnguzyK9+m7B9wJedRmmuizt8L3GNR8cfHLOVOn+dsZTahjSve/J5CeQvZw
Cm51CVqWLWJi4ABwNlBfBeorNvKMQgVXsNvoJIPpHg5iZtLtKnwjki3BKnYprMarWSd5zw5D1FBt
MRSEkl/1FztJqITnxhoQyo5W+Zk5jrCquRKkGudfmauRQCKqjQAtaiUxjbKZNG1FXM7mIm0QOHOj
q7hgE0SvZlsxg4LNuBHwFMZ5PBaV3K/cDhYhF9pWzFqbhh0UQ8yw8s/bPkmGY9F1aoBo10ACUNbr
U294pD5wMuS2vjBHenZiGswI8WMgFuG8bOnEBW5nVD0NF7l5HFE/EeRDy94StJYHF+vnNA03npDx
yRklY75PQrG0MAwgyzR3PH24kE5/eifwF1c8wwi6x/TRy773FLCC44BBsM3DfVQkQXqTVCcdZDcw
dOjFfcdPOrpi+6utKYV2I2+oOPEKGxBB5LrQbfqBQA8/lp3/CuGG4skMNhDyBrkzrtScHb5umRHR
UoEghEHE0nmT2YG1Knu+CQOvaEN1fWO7Vkgoeg9SMI5RtWtWKzqRW0YtfjR1+oGe+jnq4YtGJJO7
9qFnJ3Rah+dkTLONPxyscEJDma2Czc9Ya1bj2nd3anKvbRGncug3uZ4DKNv6Wtx8UJnnMMEmdxrj
rq81x2HWPFPzHj4tr5n6a5j/7i6EpyVxySYk9YNGTFCr2z2+pOzVQ2mKV8IXeVNoBTGxpJdLTFt7
ksiVmsHHDDnaSYBoK98fHqDFAeC9ATqJOCaNpwFKu4o35RtzSeUfRriv6TX/nlS3zS4wx50WAXYK
C557Wfw9D6hP4ZUxZoluz+LTR1ZJFOzQfWxAa+bQZZME7F2DBtQL1xvpmblS71wmDOUI8QWS0ATX
vqdBw8tYuSwmEFAVNTp0x/7uJwZqETVWE4Fcg+yCi8rmSj0SxESQ5VwBa+xAUlnNG9oXHlQ/EvCK
2lTFuudKrCYkaNGFiyQSN7Yme7EUzQt+CB2qwg5uanqd1KmXQ1ujL0fn3pw8VWQ+u12w0StHH3UU
fIfHed6BivGXaAgPuKVSJ6/2OEcX6dt+u9C18IbFIsxEdgqZChGr0wnrxsdC0OMcaQvZS3lzjT7L
bMUMGqntLq7saDCaKEvruTf8f9U/nHiBKB3dP4jOspykYa0O6pXxqEG9w7PfjKWgpyoBApYZz0CD
1UJmumYt4ZBevLDV6hWYSD6L+7BOeFSKzeFJbQjIKkUaKVxeAByGMEYh94UPSKqYCbEJHbuuAWYE
AfUYP1EP68K+mGZTP9VwC5mNGjXA077yMQq1R58UN+cqNkQfnk/xXhWKvyK3Qvqvv/koSA6FW4As
AYi9ku8zCn0L+KZy9HGvOJip1ZwXd+BHl+2Lcb8tG3KRjiQ5aygOD9LYRZF1YyVPxdZTnVJxRipL
X1e4YBGnPO9h+CWdfzUPvRCH6AeIERUfyxSRUjuA+fHQLHEYRvbUXn2nmsHHAsjLd2FBQks1Ioz+
wC12EkYW6on7GFgJiemivrY9Q5u/4zJ+S5Y0EYKs9tP/Dnd7z3DK0o19Z1l/qrbqcRN9lYLuD+Wf
UxJULE2nfGTwXoscbDqaQjruG61+0QOx948/nK64NSGAal0mNDTG+SPSYLrV0t+78Z3xTg19l+GP
qdlrKnLYcTd1LF4wPswO67DwX0H4VCWUiRRNF1WQ85uQDYurZ+agKL+2c1+W7VuHnJQ76uhbnm55
b/r5bm0QFUk04QDjZS1VMj81bDVU/uhSDkAUO/UI8DPhB2ufOVKItfJqb2nj/UJWebtxs8cyKYfF
uYGwfL5Fq3D8y5z2CTSR2avlVszITl5GzuUM/jhsHUieijfWjPrmZUQDnatZ4WSY0v6hgl2VGO1G
NGbqGYDSd36vtx/I1+dvHQ9bkhGsUgtQCrpTUitgR1FRzKNoa79p3sWJz4t7IWErUCIcgKqjtC2G
46vY68+YJB5s2ANHVKTyDQr66/SJJqWQMFDFO2L8Nu/hfw5hS/L7ALMOG2WLcjC7U+irR6gZSq2g
McZ06vdUkWIe/h6tITR0imaqZqcBaFBMF7jcT5g86I2ksoNf5j/Ns8+cNl3NXI0r1YicQtHvMB63
F/dLBp4JIazthTZuiBJ1oyJTkVvJTIygcvkoH3Eao5IZ1YqVg6ZkQIDocsI8SV1/CbfyHPmRH9Sv
K0nH6vfGaVBahmSJ57JjDgQXDBV8/u8wXGbZwxXnlooqbOAXkaS+SZHg+McQK7bA+wlx/mxU7rKH
ZNVozmPvp9T3Q6E18R9X1CcXDchzUYuIvtSKF0TlDlNQ5k8jRCgbXFd7mndwXK/2tkEbfrMOcA+h
TPE+ccBvdFUgC6s0om4sArbrF7whTis8Hki8LaJ+1tD5EH3zLKjMaN7xlNogMtv4Iwyqq3WuuibB
Ic95reYoWXqOWyqBltzjTzY4N8yrVyLu4k3REvhid5rwPKaRTtSnT28a+BBzOZrDU49OGJzb38eE
+Tz4AZfxLQJCsI/SuZGxfAMTayHvqi3L/nNVjZJgPENV7AzlzhUCxtuiko7KFDYl9bMZ/S8rhfLe
QtxcL4T5aVTEXlfmePZ6awEj4bEhCK2Y5APajxc3BqHpWTSibu9MiMFzm7hzXoUyninAj74Oc96d
lFxOewShodJ+0wi6qQVtwyu8JwPIPAYV1y6t80QHEpv2jOpgjhqzIFDPaFOYmSldvEmAKX2wtVXv
XQEYScKE8Jkgp8eNXxgCLwdeU3dF3f2mcshazS7HRr5gJNVaHCUOABi/m4h9RjQNJHKJyn+bCryK
cVkwqWvc9B0tlHO89Of3rewyznnFjndjv5eIPASETgDPq040nZHBmLAqZ2OXsllu4HuLCmDA0/R3
5V4PJUokLdexj/9ObKYm7aDvMh0dKHDvLMWS9fbGNfMh291SFVxq7lVgzzhVIwmWFlXYy4cxgSDf
HenXoPG0KoodZ61wMgp2TDrT1LPRAEuyTJUfuBGnEoJ2PEiEi+AWlsxEPRAXmPjS3j9UfekQuXo0
lYUYAW/NoJ4TDBFvhK8ySZN7Y4adAeFwP07zzUSq6dftWim0P5sdsIyKkwkLLLuHnR6ePMb3fSGb
aRMlrdWw6GX3N3t9Tvv12Xcqtcc+CirWBwytyS2en3vVcsRA9TTq4GLnuUPot1+vO4Kjn7z13dkv
cW5t+o4aURSdXOVYU9JZlxeb5aM3uka9YWYaFhjmuHt7mlSke3FqkVls0EavNDDTVr0RZWge8GOL
LeS9Xq0n7YLbURICdKPrRRnfEy1Egj/nU9pK5HsWxjTBFIX4zwa2LypiNRCt3bf0f8qMkgD5nj12
kvKFrnInGJqBnIufFsWIN0Iz/z4qKLE2YFwIw67g5/obV8ZTBYxSFKmuZnhR64ZChZ2V4omYhV1P
DObV2iIZIjUDFZBYz5tnoXZBZxIn+/Ko2XsVrMV5M91FSQW1W/ACGR+QLtmS4PfQWc3awYjuGT6r
WjkJntMdePhl6iXj0nlTud7B8Hg7ZQof9FtzAhTpvW/zI3sPFdDh0X1XaLg9iwO610Ej6FmQoFa0
h+jOhDZkqEMTudGpcr57p1HfPdpphJPUahOSU/0CvyQeZEzM2ZlG2gj/iy1x9eMNbJrLrPP3lhu0
yYGWnL+XSXJz4B/17BITcJBCbOKYv7dyz5wGEJ5p9iBl1GlMHHPe9xPX2VP8gmNeJLqUkRt135bd
fnfBq0HXV0jrKWnbC759u95nEU81pt1y3Ha72gfwbBRVZe6pTk5mR9hQVqwheW+yN4fuplcMwQcq
uKDCS357NFaZSea42t/t2HazViU0i+jLLQ9qjNecNvdiIuQ96z7ZCtApxi1mqPuUcSYx9VrhdOfG
+B9yoCGSyM+HatVMjLG47Ue6rXCgpKX1bgk6qqNnOZxUrOShzOI7Degi2sadxvsWNN0i8puHoA3P
i6Xjunvkn5Oc6bhGT5hXixf5lWYYYWxb94geYsjvSDO32QS/XeXr+cdZsnUdVj4ENOyT5IBc9/Q1
wa+Bli6VpiONsP+NY3V9tGyPegF5xRmVbkGC0rGdvezcxohoRWNK38oVpcm/9jAP1mAm/M0IP8cq
YyP5vDalwjwwIzWvUPrdVOg8qHSbQ32yVBRqrexrwT6vMQDo22FwUJ3StGkhjo4OBXZT4ckB4YZl
LpV2MJl7HwhJfYrpmgDf1ZnJ7qK4jxQFzpRfLJVpsMZ89UyjF7bEgCquKS1OQddGkOMbF9NkB/Bp
JMRst+qoPJsBsUQMe0btV9cQuzAIehwQxx02xj9uY/VnGzQe/LB65VoOX1Yp1YUIxqt4zJHNTx9L
f7ZvueSQa8eN2l4Ro0S2z74QQ5CDAm/30Ejs/gmDntgSNuXoP6H7W+4hIgJEAikzFIxQTin1WK7J
6m2DWJB3HJsCFhF3dCDMxfFndlkZEl3OxG5fVNtnObYlvNx/Kh0TF52EpJeq2D0aHKccm9ZTwxrd
R054+RUz88XDf9XGPQagk0mUqFfovd34fnzR/ryxU+IOSUDSdLo8w3Qxo6kV8pB2qXzPMb6vOqiE
Urq+i2nTYxkpGBNWuAi5f3RlqCWoba/ONFh+4VGD3jNGMsMSNPoLhknkQ+qQA0K2F7oLsH0MS1lC
nTJ7JLwCRl+yH9RbvSHH0O38tbme5SVlHVTe26OCrX9uK7+e3U5UEueK8+XMsm5sb6LHGHixKr2L
9IFYePOGYN95Ou6UHlQdGPQcS0mNDOR3LROB0BlqyPzXDsUGmLBL4XHX1fbLT8tsh9rptAlQn0Lz
0x+Hh3CbwyDnhCvfZ0HaNidOkSGJnatqjg08cZAOqKBJ+lGFAb5jP8D/YODNKy0J82l8/8hElIak
FNNj9Ey0FI0ZvtBobO3fo8zh7uMXera1527U6IK2P2KZaMc0+Aw+G85ZzseahkzvomPgMIEr7w8s
w2NjLjL35uV7vP2IQBT21YcxiHk3oLBJRZ/K+0jOiJ/DOGTtLxy23w1oqGQfHNpV37WcfScVvxBj
/MGvd4PW4wg3y6Xizj17I6MMNTPbx/d1zmVsG7Kup/cwZpJU8KoofivNdN60ah77Z89iUqe0vSBu
Vv7RvkScohimuRRIMNEO6QFk4BRVmzTYY6Ks5MrCvsbycwEmhWtx/X9tfho5SKHDvc9dt9rxXs6E
6ZIk8cKermpQ7sle6Ykoc550rls6FpGV5DBaxhlmocKWbyzR7mRMQstjXFmbzuaSnTpoZ8MaML8I
Uz1CgZeq0RNAzYzA0cZd6uSu8mv6g/o7jVEODLqnMYvPC8VRGq+jhj4Me+DftyGc5GfRhcHn2exb
+HeynNYpo5JuzIWSvMBZtnWkk8QEs/c/BnD1yvkxeoewf1saY7PkS7Z5DbpRFy1zfoR4mvhxUArB
mw7b8N1lYUFzpustUa9sCVRaIp3eA7NN7Ydj8DJvDCG38COWAcoueb+x2N+irIem8AV/+FqlDUJx
ORgy1Q8avMRLao35VEyxrZHSiVCMewc13pP6qFlPb/+877eRox5qsUlWMquXAKO7na5+SuLPncii
3LrrukANzf/lcVMVvpQm0Iww/FEmHJ4MB3Ei9LZl4as2r3p5XVQxLWmYQ1U3cNnT6As1Ui//gY//
xPHHjJZhauAOkrb1T0sZ+JBX+VHcfMwq/qh7Uj6MFnIDkcDiTUZTQ3QJc1dZEp1Ret5V6rxYrf66
kzA/sF+ZMuY9/8x6wx0edWaJT6JAVb0+063m62tJBCwIIh8a0WVLGSf05Kc19y2ZDS1W7rKkVj6J
4NOfm5vdcGyk7HzfSJSzO4IFAH5Nz19ZPWNsHpenoJevKxr71hst4FxwTm4LId8tMDDoZScKPjNH
q9dKTw5LrbAlbD7N1ILTK9uESC3U1tkbGQ3ipzOVX7HLaWtMORReNP++wUj+sY4/bopCmPvZLdz0
WHYrAgr8gJkYt3QVVaN0dvA+nv1JXaNOt2VkE73YSTRLmqu9wbO3kg31Hvtm1bfIi4P+1Ks6swkf
7zVvoJa4WKd9jlGXd9dpWOQtIeI/DCq2O8iPr0VhvKnybmM3uMlBCyWzy68ok7wyFTO9eLQyB4Zr
XVHReTVDkB4oXP6fCwQ5/3dRWwdHyNRfE4xZ+CmpNQEo1I2JgoxlxNi6CQBQ4x3ExBk38/I6DiRI
YK+4aWyg5YaAGi8IP5QPWGX40zB/cJwAXNFyuybLHG51i+wlxPQj1YC17V+erUvISmV5Qzdf4gam
+UO+kLtiT8S1JHMFLTOTEO4Ad428Ke1hHphkGXPfds1N9wlfqvghl+gJOEgz5DedsTU/oa2P35C1
P3JS1qtQEmdrE2oA3mX9wCdpYQ8f9sK9GE/5ocfnNQ0ggqQNd+NS4hiwoILDGSMaIBJxrSo28We1
r4iWF1HwgikA6/8j4gszdXyX1gSvk0ld7U+9D3iDiFRB+/O+WLpzm8j+gVDRtO15h6C1uxiIxLs7
daHrqYBmfZIrvGvJ1fiKCPhrLtkC38vHFRzKSYN00y9s6aHnFM9njR4UqplXff26cJpwvkKKtK6j
PQ4BlKdTOzSvYA/mHUf5rGTeZo416dmg2iYVpgzQYS5F20VRGJBd6cMZ4IRg8ZU5EvxLqT2r5d1Z
4ljJTfmXwuTpD5NMT00YvM6gxkEweZz1DKUBBs2n9ilDvzsoE0PgEN3ZxIqW64giXuc1nk8Hdmn6
6ZFyLmZsXba0jMSlIiCHWQb8PWKkKtALe7vAUpwqtWRnuWj9uJtwx+J8jKlBgHG9uZa6rSasR+SL
Lji6aGnge6XxrEbNcx1XO8wDPMLruwZ9x4h/Zj2S9A0NG+fAFRNUDDm2vRPn7m3mDuwfaIsruKNn
XGIzjX8jB7sygV0BG6O6YPPjZXdjRr8d5AQMaMRfASEvhOilU+jrRy5za10hdJFty3GIlK+0o8o/
iNEqJUgPXlinqGWBV00T0EiiRUlsAv8+gVYU8iZEbMpDOqsjrT+1jKi+NWtquSdnD47BeLpu5/XK
IPePQUwo5s67MyDx+jO2lbJ1VbxtcqanAPKNrp5L3FtUldTwaGgs4JVpi612gEtOmRIxcdbDimyg
QK3hSECSEd25dmeVTMFLv6FrJRPV+UsY8I6b8Hq2Sytm1cuS/to0YaLeqVlmfB4TSgkbIr3ZHN52
aNZCOSrYgQnAxOQ8/GeGiLM/6PcAhMoOOCv6h3K6ELCdUsT1nr12d223ZBgcGCfunIedNVOF2dwf
xv1z7Sdr7p3oSoOvwrQxuvBKomKQE5ngBdmpQOTQEFpnVNwGw5f8VCvn7cHmPi7zjnfA3xcm+ayh
g8ZzfjGa2Sb0Myg3b7sAWYL9lqIE+Jh6mdgG3EdnMamtpNZgpTI8ycwFAkPIp2bo22ag3zecGMtB
q/rV0bvTXBRIeJ5eA79XuL38WjyKxXjGQjHysHzwxf7V8hXmNm+f1iOgEXFD9JJPBwSnYGB8rjbI
FxkmVJ6lWB98dz60OMlRdUiegZp9epSIcGy+Fr9fESWl31g1rNrY019jgJBMcyQE+2l/e3/N7gux
6Cei1auHP5XlispAOfqfkqOi5DkD/ckOWlXVmHbWsqslZ373EH5F45gKEcGvBr8zTutJRYrWg75y
u1B4JF6f4GoJB18oXN+JSXrwG5SqkHh/WBvq01V4mNDmRN2EAsmsoHr1ldntdB/cIXLdS/tHoK8M
8XWCXxUGSWVFLHchiiUUmMUmRLXMzbeRoo8ou4Klqy21+ay+/IHAknpRGsvawWNJNcXwugOO0z/M
ht/OMOHMT2HVdf4n2K2/lQFiGK2uzQYt5SIHY8sxhheAkwKOxFSy4uXu2Vjn/RSeqvjcTh7TgBEZ
UloEvsajtuR9cn0MngLUN6ndWkqyV0PsfW8m6hODLcsU++Qr1XSWGTRrmevhd1/toxt6ka+f2VuH
sjZM9xN6uH40QwClOEg26sC7ZoetDbOhwJPmaR/tE+C0HIZE4g4RQ4FumHJGujCCJnqW9qNEIHcD
CvOc6BruxCRV9c6IKmTVYK9VnX4fUAAXIp7xd25B5DbS9lzbBH5yGOgkXugSGh7zy8BjycdNEwtK
18sHh7782R9jadLjwmcMxOK52y4srcNOF2BrW0hC/4vdJjGvEkmosEbSr+4l2azTdxapJvMkhSxP
kqwmyHtPuJM01LxoLq8dAUN73MTUmwpWMo/3G6U+1+l7aBW1ceY2eUsfjMj7iGCXBQ2yuwAh+aQn
2rtniQ8uWMDbBi9JPjMSS9oF9imj7WRlj4BinHswAVk+AdEmPw+CkrR6CRyjg5HpxOjk/QB8mYac
VwlbrRq9erzMaDY7e8rAlx1HM/LDV92D3xUlj2JvZvvDNkk7X5GebrUwRsDIHvC70Yrl6J8u18Br
xlUViUxfp3lQZsiBmGsP9KV0TjPhYnPz5KIyeSB9vPtMmhLZN9F8J/jpFloiCVMxPgwIpymlN7vJ
zsgS2wdDP6X49Kh4xe6XABxUVe9110BKAR8X+siW1QqqiWLRapaC61OvfXHyviP6X2lDwP7PJ++6
OoZw+N765pvB+bz3mWMu2peBWsUuR7vjORG98WNbjz/aAWivg/BgPvPBAWXU0ZVN6Z/ZF57HLGlM
W/0a6DziEG8VDCWbICe7WooyrPY58nvuhjhW5/efiUkR03wnH8zVLXpo5zHjyuVAtooRw2aCGLIa
YRjeXAKbpYrxbYKWwcqLEpyqjg168Bxw++f9KjSCGYGemE4TJB3EKzyI4x2m6zdHgx7mLsTon89j
92I/2RhRIG3oGavbQiXbjEGOEFAkG9yK2QwY1L9fMZiyF8wG4lEAP+ZILTU0heeSy9PID1PjsA84
vF0rF2GpRh4mn5iAg8u5/PTjT9tFXy5l7EPdRG/IY6RIiUZFmJwsA4lx7yTQfqJq4m/yvJM5kLeB
hCg14s8m7TEKRg+pWPTZMyYKLve8rjQeCAIZcMRb+sY+vTmwBKI7DP5vuE6yI+/Lf1OkGy4eaR4c
4IHk0viMA+rhWPdkrCqcGJ8jM26C8d+rwapROb0z/1MBC1j4WErIYUp3ltCjpcTdeHl63Ps8EhXz
9zAJeInUagv5jGPHXr9d4g/H0CqmVl/VdAAY9DiN1W24pRc0NQpqvhSh2r0zNNckHQRfmmcfxx7W
Ynm3/a7GgjokpPjuxW8ftorGekE6ZqSZK5NSvoKYpQqiCvEp6VebuBR3Pj67Ltqtn7oLNLjEfGya
MS0Kvcu6ndxFSM3OSXHY5CqLI27JURt89QyMBQPJzWpCl2UwNiQ2THl+KrigkzBDdLwrgiATIqSz
b2qHJCNaQsf24UZ2H7OmYbUfOKQDtoaWoRwJGq/Gz4vvCpMbyMKGQ2e3YHvGtQyEfBsVN99EwljW
W6oYrTjbnL4mMe5Ux1+9d4EtBMwiX4J0/NikwY30pqb4gMWLhUAo8dSPPWXAml2GBM8avqtrI3AJ
RT5KgLCPatCzqFDVas56y+ajnxlx438AyjofMgyoAWFl4frbsBb+qcKHrecGLfbzqVmxegMPXgOl
Ikih8ehNG0OmmIp5VCEjHEQh/2WeQ5DQqmhoX/eR3E96WZaV+1XXF6NxDeyFbmbnYcjJt3C/870I
RWeBgHFjxgr6ubKT9z6PA4XnCJkEmrkw65sycobp2GA6FgLnurppzDK4bHgc9elhJB47NPJR2i5K
CqqkW+qZsDc1O9ytrUc4iryVI/52G71Fa7x6Kq1ZeI8auNMVWSbiuAmOWa3hcQZAkmYIdj5Iut/k
SMcesK7LjS7lsfXQNQZkb1hZnLphyMojAGxc0LwMxhXXNrO7Ko0GcDkPEfJRQ+5bM8FX4+hcW2Dz
ZS4R++2xtCdoGplpAYGNb4C/uzShFOGjwNt/ccs3iGWj9CREofMN8liBm3tN8eKLsS+qQHps0m2Z
tTXqpH/CK/fMngIB9NMqMlInjKRJgapjAWB7yzEzqxODdKvEgoDwPthj7MFzSr3phxuT/gvdMeGC
ZDbu0rbZwwiUkryXAWzkcySuQaNMiUUiYsOMBUQR9QL/OEZB2M11gbYStHpTK4cpu4jqoK2jkTM/
Emygo+ToerWhYDiQZeIXtlqbJWVM/RK/aeHpt6hI3q2WJoSlqqk2ksbmfCwvNlNIi27yOYEktLNf
e4gT2UmwZtYqR6YGQjzvBZogAMp5yfa3bm0134L7sUFAH+s1ehPDjdv6LH8SpHs6OH4Pbb/qR0Tr
I+g18yrL/2p/KMj66fseGQJEWMdyqE7Sb0sm1DQhZO9Bo1GRs3v3g3DszUtdQFfj7O74RdaQ6ixf
VXI4Hqbu0fJup74zWyuuBUpVKzjSpyKk27+Rx866Vyze9EGVNhmWvtmItgR0c6gZuAPYuTZ/ikdr
TjxZF1laD5KMeF8quPbC2ZMk1nRsKg4DNaTK3TZQITnrhSJHUMSuBQqGvNpuRh3+TLqnk2nQIunA
MaMlZqQRdlXBJYOdR6mbaehnD06wWv+Pk/J5VI4t/1T4chTnN+scpMjju2VasuQgT6Co5xRjHpmI
R3616weIxA6zAP/Ym2yrH8Covx+oQu9RRBdImkkU5Dk3QVEE/lWZyNPZcXEVhNBEH9pTivcb66vZ
AhT3Xk+u9GYjpnz3GjwJ+ErbBFgcLg5WDI2Urvp7diK34ItWnf4yBn+FbM8B897XNStxZww6Hi6/
mH+t3s5RQ8FXjajPHLx+dTob5xlLWvWlVuRC20ucTgWlU+5CLaEt7fx3Co9YB/pPXwwXWXcIV6C0
xwVryvpEBRPGm46S8XY8DGmfr+0/SRruzSO2Cj/PdAI0p1tjvZ3WKlKPHJvS0NxXnKqJ2cTP0AVl
9/nop9vFjDkEhvD9kZHs2IOtNNNaKQyfN3cSAktU1Jr+tyui2+iBkqhR9OASR/D49+Mlu5invMB2
/tt5QdghtW9ZFpef8vo6Lw9vHNiwRhI7dAUXFbKc9hE6rfataJEt1YidvGbxVQ5H0gbZbDKQDUzk
ljYNzhZ5yddDC5oRqufr215VoyiOSEORvnquD/sgvL3wFFzQQnXfgTrm5o8h6A4n5VlVWhNJqzZX
rA7JXm3KCRlVxqHYwuo3E5RgNyKdzsgIBQvEbxbUFNT/3Xv3UcKfMSnzs94uq55LC0HPxD2VuH9D
FkuC0cANdNR3YbUCmCsl0j80g6MpFQHcyQBRpiZ0k55kEJvwMIuIiKrtyM8ACAsyP08I/P/jPXgk
SUjUrpoBVPu4HTL3YG4vcA5mh84ymnc03T1U5oxiPsD8ULkTEBzrXisyqC99iMpYaYwAWdsLpNgc
7slXsNqxmEnBmGuOp7p5z5WSLBzAhfMnNOUo4Unjd0XmAavt+F9IpfsyESX/LEd01qI0JNtaeXZn
TP6M4ynFrAoKntH0GyAD71jp0rY/pilmC5roPdUOvh3G8i7g42l0Om0Q94N7nC5BkbOi7DzHWRw0
kjxQ5WXB5AvBwmqj4SzF+syJ3CPVvuSKESadtqS0TeyoIZHZomAqIeoXifmYTZh7qND+5+JUyZ5z
sbx8hxFS4qDcJiMSZYu1TTCRpqHYu7kFcR6+f67//2XCGEbhEzxemSDV/qMBDQ8/8ecByZIg/0XO
Ka039mqDJXt20ZTjIbJ8kazAZXBGy2NQ9gHbd4C+d3j9f/bc+4Zd3r+dmhPCEBEIielVWpl8tCQX
KP+aW2wR1KCUQHZYfxq99dLnPVk3oh2qbhioA+Fo5ZYYLTMjJheuudkekGWkpenBFYmKw+hKHUve
tFyuRHWr9pZfC5XjQCJj5e0lWp86lLBye7+tAQpGT/w/VOrGEYzVUZX24Aus7Dq/9Nt/vppsbgI9
iCQ2Jm/8R8pPG3wGvPDIib5ZQvVi42aQJ961pbH24k6wzibhGLbjtgv4XLkz321l1kJCFMzuL8Lz
olu579bWKeIkYdpKOC6hCdWfEyQ793dBznHDJwzsNTEr56ZG8j9Ysv7TpIke/Oh1EuDvNPpqG2tX
IWdxnADnQGPn8hhdruPrDlgid+MhLID4AzCnrtaoxetVgnTcEhb0JWMYn2A8yhCaKAX2Fw5wF2A0
k6btgozbOPaULyg8rV2d09XGJbhsGWONTxKm4WhyMU4ieaml8qF2ixqPikLLhMlnUq83u3JUqUqd
M3+K9aoV1H11PrsHFrDWnN/dCvR7RBO9LLJP2n2RjjqdfZ5AQfyUHsYYSIcGyyjERp23mAmN3oeO
tGeI8acB8gv3Utu4r0ra/CGVpA1y8YG+ugz7jJbTxlcnWtx8g4/9zqxedkb+cnmrpd690qdctr4O
U1dxbThBeQiMStm3bW9fpWc1oPKIuv2P0giDpg9WeYKgppYNa4GUIF62sQKZhrobHSldsa92HNuJ
LWRnnZ4mZYleVIJCtonAduHUvaxV63/1E8awK2MHS0NPxjNObQNPzkxx7hSiIz9CcKlgaBMkpMzK
/i4I7ibpTZ9mxtPcsTKg/iFd618YdN4Y9uK/7pu8l6oz6sSlmmthtnlQcm3O1w3lDfmPSv59vavH
NowTQFgPiy1F5srul9otW477TjUiB7G3DwXzQsU+cUhiQ73s0tnCQ20qo6cuMOZeaRW+YVzDyWht
TTZkPSdI/qVENzX740YfcYo4H5oRkSx/3TC7/2k42t0iDZQGc08S+5JeBIm4wqdG5hbIHHEauU0K
Ef3zW6WIO/XPe4HrAghaJNKmekOsyUuHZ1BJpXyM+AICmdagcCR5z7S/oB5271CVVvq8PrAggYkZ
4w67SZARrhAbaZS/phsVQXtVnGGu5PtmZZ6pe07VELL0GhIrwo7LoK67TT88j6YmdewVJQLnjJVr
Y47fgfhk87brU38K8wDNtHYM0Qi60+lNTSYGJhSM4WEWSzu2Ez4umSoJOXMCJP9kYpS/O1j2UsTZ
tj1WIEBSaUqBWgza8SMytjL396X7qr0bRiok1coNOWoptnSSWkfPtqkGRpxDssJjOHhx9EwBqpZY
feFVx/Y4j8ewsBLWIKuCX98U3CUdW02gxF0e+5oo6GktSbKjfzPF2X5XJR1OZlrZPH2wxMgqF3e0
Pt9PbuIXVDhrwcKj3ZIvSPOXLRsOzJnsk8aOsuBdoDOXQzCZ01qN4jFvrXHQ0NRzXxWFxgRDLvvW
zfBUuMw9MLy6m1IuSUdhG/mYKzwny5XXFuBIFBDWHHpyzU8bLCGP+ak9YgEjcp9D1wTzOfTrt03T
BvAXw3HMqb1ii+iatiL2QQCghzQytchC/gkrUWXYbQV6w3lgWCDqQZBlBVp1+lM071Wyr/SaXBpo
8BQpfoKs/6iXFO8uK6rwUzU7Y4ej+upcPJ6SDTbM24vrjZpHp/x6xrq9epLGzCU5GNJ81eYAjRiK
sBYC7oJzv2p1d277/cjUcs55eEpKGy1XJ5C70n6zI7Ar8LjCGH55dUfRLmIdU1LxaV/re9Ena3jq
k5tVn/uQXCfPZ9COsO/QSwRx9+gixdHrX725sLfQTo2RyXjZzvZw+ymsIcomBRHksPGDt5rf0+Jk
P14m3MVIVEDvfj5ITznuds87FVPKhGd17T/udZLLkGzICMzTm9RMTSeanbqlsq6qzAReigmFN4QP
olYuL7g4AZhXhLchIAU5MO6I0hyjbqCHyyOUNEfWk0d/Kfjpxbykf7/Q/4QH6T8uu2nnzaXwHxDu
I3sJpUWjQZGHH4GMWlVXP+NHj6TcRQk+qvY0pJwhhn+bPSTw64RDLZRNVaXpXKuoiBVlXjY+sZNa
wdb1FE4P8vkHBXiLXPdtGsQMqjeRK2W/6KHODmH02rzQ94ApgPo7IG57x4FvleEbg2UpA5IcxoU5
Syh74ZjXO/Ed2O1zEBSIVJBHj2w3pFzVPifcBMd7WCEylfvjy1YbOcR6xvqMpf0I9vKkPVVQv0Iv
V9TQKP/TZZ/O3Ey/k6C+3hTDy8I+XWqqF923qMdWVcHXnOhuetZknBSedBKzGmovNoCE27SHe2o6
qzsg54mdqdQp59RfFwTyJEiXsd/vQnjgClAx2m4oQvq94B0+YpmDi3qrTBlX80nSwaKghx1kaX7s
2igd/fkOCyCpIeHv5Oa7Pw9iQDY4MjuWLlmCOB/u9JtaatXC1i5zDa6Bq++qPW2LMhDtk1YDWqaU
nDkbDbJhGCh24YaGWmyNO2hxnTf0YS6h7bLqu+22PNQajqpUFQivobgj+tmgz7yVl2hyIn/F9Os1
m+ig73ahzOmkb+v3LDyjRW6RiWLCtYTmp1zasRArWnwwDIRZ0LS0Z7LUqNgtLk5LtlYCKqcdgexN
1Vpxks3DCFkTdNWrxlXCafr2NzCj5XNoAx3Rjfst3qhMUr0bhwykR0wIw3c2iMHJGiVjkXirdVNf
v3Rm9KvKOCAx1x4chJEr0/GgaEW2ioqucvGcHalrQuRf7B7pMy1yev7pWPMZg9mk8zePVqQmvz0G
WKv3XCnkFwbD4mM2iiPWKp471BOpy/JUg3MQKKWu4L1uzlGjRM0D2/GKq6zTUb2YrWaKMpZsh6d8
MmxRG08y6Hnhl7Bk0tdP7DUmtTjfLMWX5fbFmt8Hbct/rHGQRcGftJU+vmI8YgZEXEg8n6sU6BmD
ghxODuD5vg/NvXjrdBHvr/rpPeHRkGFJqDZ+TfNTadQdKat+99feIzUh4fABX/RzMIz6NYgTqYSH
khJAOzfkU5DY6goA1U0Lglx/4dgig4kMe+4ECvp7aic5OhewHF2KB0t43vSsX0WehcxoUojoKFOa
9JjKti4R+p0mYmPqwOa40twtu1r3A1OSxhp6t3jtOpA9Bkio5Qdc3+Xm3OV3UbcugaaCJ/mglXVS
3rytgySUfZ44pJv2big1J4t40ez7VoxVRSNTCg18mh+AiH3IlngVY2PLu3vnBFiqzSVVVYseh3eA
gJu/aomMBOxO8s7PPgb0VJ9tb80+vdv+tcZrWAoB3NRidwQw1Oh0LBIm9cqw5CUVB5gNZkY9ooRq
lzoWMpkGsAt4NsWH4thXoI36foJmDrORL4oYtuIfNnkVwcGUeLP7wLBdpcGtqBOfEoGmfhHPMk2X
LHJrzmdYrhWwLQDfh60Pw3PX0iYzkwGsrMRkazaG2XNSO8wl/vXZQs3c4uTj5tBBbAW/MwPq1u+2
sFDzH7KNhqB5PbNAObJsDCUP+mx/xbdA3DmNwQvknJJ3XYElQu9h0ewxZJFpIHBD2R4JYa95u7en
mnzXRen0yguCJC8QoZntZOkPIk2o8fR0I8zhw4N1HB778P64Pk6BYi7KLjRAQ04MGKDzx7q2Zhbk
WUV30QwqbgjR83NcqS63uIiD9XSNq+QugvJKqreti588SONN7r+AzA7mTKx80xVMT1R6hFvSKTrI
h0bWmCTe0NLlMNL4K3IK0ntIkedGNm1vojH9KDmg5aXuacRjf3v8CaZkf1lRX35nz8SmYIbm4Kba
CxNsgaWT3JErykRzjvwE9Qo2U/1bll/KCpZzlhNlGpTMcTZyv6VOz6+K/MRawj7NYlxn/QUuXb7S
2ytSO2pjFE+bZGIqqDRJE2IcP99H9v7Tjr/AxrhB8LksJJ46FlFmRsdGpDLYB5/+F9tgY4Tpm2Kt
h/v++hE5D+cfjCRzw8L/HkPeOqQQvvyBPnvAW8/tHlgazPwBfSYLHWsZc/i2PZvobPcEKfDmNcLK
V9AYHHzLw6cURgrCIjLP6B950Qy0BqUt2TbLHVD2O5geZFkGeUFTXoIhBF7lwteMDB3kok0Ms5+l
ij2YzFGbm0d54LhYYqC+4YdGnRmkZIH/WcKyOrW6vK3AKAHI6HYBwd3Ycq1LynP++OUl9SpZXmQ1
Ytg9uudB1pDVEp7fzqwO6K0j9o3/NwY8SGnjysxcQeQh70UABqEDcwq2W/6CylzNmxo5c1CbvYOj
mPac52tSqrVMUiLq6GdMsqLgOSsdvzbpCvOl9I0bt3VEu+PX7wTYhGOutDghtCNxAtxTRw5m1elo
DX4n1JXiP0IIfD/iS+xzVRhn2Qk4Vuw7YnCBMHy3RnBFxqkJ+I6rfOLRupAvomttgXf9oNpi7afe
ggujuEwfuC5s0s8GfUYNhvyskPJ5A6pRuQQnXtiqiFQSNvrVNciAwGVqpYyvXE9172/GZ7VPfxLX
n2I3rfBGeODa6DtmYjsDesGGEGuASkruC+lWyHZIKf/16kvaWG9NdxW2H1MQAYos1FnDrg7H3bne
xn6xYMCkqE4HaCygBchqqJUVWQy8Ad3uuVWF/TA6ZzmIsDtsUMuUAD3d7o/KftVrsedWw61T6S1d
+pAtJ4/TSjk2FF2qMwfnbAhz5OZD/gLRavG+bPZjEQWQAc7YMRTloCRQzBh/Id6dT8zPal6744tZ
i9NmXoNTYUsDY8wqO6S8Z7Clre/NIzKxKgyq8BLDOQKW2qNEsLUGQU0/hePUF0FbdgrBF5Lal08P
s1Hq5EjRe537RB7FUfI/cYrqX+S15UTxz+9LjfNG4j+eOVMKymH1GCBHhzHOeBPgy/yHm4mSK2f4
fW3VIDk1LEQoRb2pvqPFIfkUjciTZnHoCcKybQK27ZyrvScIB2XjrMFI6jJ5o8f6Iczh3D5tQq5s
QCBro4tHN9JTwJ6wyIvsv8ld6ZGcThhImA6USIdso+DM1wYU7+4q9eq5ydTjMMLR90Vw0sUwxfGP
HrWWPi1BFxvkB4U737/G3y0lxkOZg+s6HYBVGMDfW6iygMBQ07Xret63dtR3ILO8U7qZx7tHFgQD
wkIHuTzhhmnX9udsEGwI7YxiKFWqwEk0+bQOtBiqEHhAE/d8/ByQ5WRh8O43DYJSZnV64vj814/n
9bw2xjzrIPK/7TO8iWpJ17MDI2R66hE3B+AUAhgyesdotjP/PJAX88bA90Q643iR22yIkNUw5c9G
eDu529rppuucPX05Kkn6rpEQNjSTgB5kB8D+BnfV4mMAeBX4MwPPwqKVNSkMYVA1xNJbt/aADm0X
c1BbFhQJp79tSau4RqNUJ5OIWeGdbZ7eJmU8MY4elFG4kJ/bJiAgKy8qqufMLJ72AaZ8EMpm1TEA
18soruFJo+V5PMbyoNKknD0MdN9aVczlobm01YsXfaldl8MdNgV4BpTySNVXv0uTvAy6Mq7v3pkc
3oQpeVgjI4C+D+U44Jq97+RgT5cMhXGJh1mEE26s4SscQsfKc3UQfmD3v+AgwPoUUUQRtQBInJGI
5JrApfLrwXarkqiTx99UQ6g/G3xcSc5dMER58gNx/mMZY7FOrG2mgNSBtPuozr5qnitVQwL1JSAJ
wbJBkyKti/AFeFPAlYlyn1LzH3HDcku18EBuJuPUjDPupmg44uwLfNLhOmVjF93vCCEB/h72OwBR
ktfbBLuPVBeJIdBvac1myKKz7mN9qQG0prbL1lXS9JQhOaytuduNNoS6DeBswtMAgAYF6S+OT7xk
Y/Z89sMFs7drBus86nmML9++G/5JYjHyqyGwBLTd43LZZgs2JwX40EceaGxYCHh1rggEH7CFAn1C
RhSAuev8ltcscJQ67nUttqLm6AAkIcfemil/ESOX6Qt168FVhKts4N4mBd2S4MYxlhpO0Bnvqx0a
lS7AP9QVBMA2FVghZUuERaJV48hkHgbxPvEFJjDN1qco+2Jsr3tgJv/t2UJsr2Ns1aPn04sTqJfs
yJRqOS2m004vsqKKOxWCA8F8bXexFsCd9PZkQ+n1+HLL+vHcEJjgxZTGCGH5+cWgDfbcyS8PmfoG
sefCKO5Zuw6Cs4TYQ36OtjpbNUWVA4bvEudvQfpmI6jo5avZAUZUoF1rQlHHNSctSD+T59+uvw8P
k/KUPWVprMNeeFB8OsrCoUQTeRzASZ695m6kF1dz+SVz/KDTezFoNNX+U6dH39MTh6cGJTanvUDb
PLpdT2dSmwMpW7Q+ExaP8BRAsGCXJP6I6Na1hOkisKi89CNEzo65YYsym5Ic0o758Hzbux6Ydzml
AuxjO3RCwUrF3hXFKvB+vgA3NpMDf9bD6BCysfgA67GTr1Mm98Ml1njMITwcIk6Yj6Qcs4nRm6ck
iGNDciunF6dr4fYgpheoHX+aa6ivI3MJd/vZ871oucbyN5K6zxyv45NEEW1oWn0sOEmI5etnvAW+
dez7l5PLGnhCZiDXoynxgFI3wDHx30f1S4DjmKO0cW0p6tvKCY5qNk1TDpSY4Du5tu8MF4ERvvIa
056r2JPOg7VUJPxGHEBcXuZarCtkUtbALQzROn6EnOG06hJM8Jo7rU8rV1A7I9gT1q2Nuvg03cCN
MEZHUMatBG0EIlYTm9mgt1d1WNpKX1c3ymDJKh3IBg098EulTrvg0Yg/QzI44tFI5jDdWKyjELOP
3MjT0/4vENqL/SYyq1VRplnFqJd9rN4hBWkj1NQXx6nD6auBlsSVobIanqmPjVSPMjvBiGBJZi6A
nFovF/KxcZ58Vc7g19cKPkicAwiUMmvtBg5iRFKzzfFf4a9o6z3BQOmiX+JLRDaE80r8GQnP5ReW
Bl8pLMlHUoCYoaCcC0mzkORwp+uikemUcap8tVjxmSC0Ka4yJHaEfqBbGN81egmFVVHL40Jmokrp
4e/MikHcmuFCd8MJXaUJQgGsTK6Zd2xoMWR2QBC0arjB/odssFfC1QSXUlr9f3QPHh5okOogRfQ4
xQ+i4HarI27vhAeSGb7485dnWl5vC7MC4taVqfFL21gcXS00PCZ2TzMXDUthFvbfXv4nBu0uuwJa
2fw33E73+7M3CQaI68CQTH0/KgKik+CeydkGxYlAmTwhkv1GSHiTshdUBoaG7T1jpekdf99OdsR0
YqhIq/PIRYvngYK0Wg4hlh8XL+o1k2P7X7rd3HlW0mgomTphpOADQmYpK/2t9rHkJNH58YZBXjjk
vO6sZvKqCC7tHa8GiTDrq/6Pdh7Dyk5PnYTd2dFrWkpDhdYXFVAoYCit3Nny5W+fqC+LyDATeg6f
Q+PVOm+Cp6Xa1k8TRsnswECnQk1muNWtYxQD7TVvvfSFOakkPPK4j43gyc2S3CTi7teUigTxLt1r
NYciZPhXquSANy6+A5Hnwh0YCzSiZXNHlDnSON1O6G4a20ki9pLQw8GSacjn7+S0uYAJEa4OLin0
eSvFJdATPBd2kzgHbE5v+seCn+UFYvh01NfK1FTjqX3J1hegysr77604e6Ye8sulV237PURIdqq+
hBBQcI7bSQ8j1i7xsAEaBPqg1j7sFJfHe8hXH/+nrrMMzSBchY4XFEDMc5yD0jBcm26YD01dDAor
cvaor3kINaX9YunjPco+BreaiGpd2ueJ7WmYnd0Xji6Rh/E+ZzQBCuyrrT/ZWLAF9iFfZxvX6lgT
Sc5rXWAkmNiw1Gr+shnvszgJDn2UkASXZQuepl+Qg7Wje5qxV9gAFcdev6bRzxiKC4QEk1FnhnoJ
VddEuLZdLi2OaSePTfeVx6zlT61rjnZwK7+l/WWhcR+Bxrh9IL7KKR1Byr2uDJqcya8KB8/DJdaN
h6x1h2xGk7vu+kQ7FqW/UMgTFqixAg70f8rhNNHBh+zWd+prXAXrD+immHoCycHacOKpyolt1UNE
2m463MoLgb9QUOdZ/wyUFHQC1g9C5G4jR582+7dpLxKuqgIv0OdnOTrkLNMqcm5sFWSVB7c31K9+
p6it1LgMEN0IpeuL7ClmW255w76tO5tX6V9kXkNiB5+52KlWxAprOm+zVqsDTtWQVxRm7M82Ft2v
oIa9RiXpaLolSokE6IO950WYbAqrsIKPMhwdCoJDI/QsUooalPZd446PnPq9Lhea8tu4GBFscASd
Acj3A4ltkI2BcEIOKGgUceuKtFj4eSOiOtKN+EkgX3NwCYe6Mf/h1BjMJpIkwV7HLNh/NZRt8iQk
ZGF2J74QmIVcBLJYJ7E9u65zcGPVwTJrlcK9Y6ch2BCXsO9Mf16l/6kWHWr5clZw1uRtQfNlx+UX
FY7xNoGpoz/etQEQdH3IMnFvm87GexIMpRo2Q+bifPjayo9DCU/1agSfxa0hmnGdjZiKlCYOAPIS
7+RQacCLYA3dWmCN7HU3wRpcgugrQgylkXGwAqVfKM2VZf4YmFOz/terAzkn9VtsdEoe5pzSWbLE
b8jUfaY7HB+b/gJJDomx50EwgvBAf93svFIw1TR34Dth19zUdMI6PnmEns+RR5ZOG0ZW6z8YWSvM
MuF4btLR4WbQti7n+rYHJn/Hd4i9/E+VBCxKdK5WEy2ssb7CgIdF78fH6D62yt+ChNNH8RJnADjv
ig322b26C4r2ZFtK6WrCGEQOKIgtRWfK97rp6FZOpo80yWT/h5cMlJqEk+BjOYuzQRywshYkaAmg
G7Agd38n3XWBAzACzbMCk2gkX43gQoEorBTUbAdD7Kq1hXARFgc09u1VpFuAyjS2I927DdX9Enfw
YIQQKxMhbREb2167RWTrjCVmBjF/ib70gth9GvK1hX1kZzv6Et+suG1H5TMQ3r08u9OmBKO9pTIp
GewDe279kScFkpDBZJqODLbLaQ6x2EyOQ9miI5GbcLXtXEzC6tXi2ONqMbnH5dy0BpVQLYEdb6kc
ZXGv8ROnx5NrZrE6uzjxEcIJXTGGDIGGowwiU7dP5V7gVSnY0i4frm0BBINpY/pUSjBQtWEWMg/W
wRHqp5ycQc8PQDTqa0MCc9cd51/0edepFH7l/uz/o8ChNCZpWr6P6Tcqorpc0tqrx9XeEsUt+01a
XkrS26Oz/28taANhKKn5a+CzttAyFybMv53hWSo6BY/9m8US5op34V+uFlKMG37PNsf+5aXlZys0
xxIFUe8y+8sh7dxXTYWp9UCNajwoIm0U0ZJKVh+HrmAX6DUdrnE1VjcApFNalcpHoGxo/iYSKI6O
v4jrS+IbdLzY36lIf6sxiQEwcW90yvrAW9Sb2AeqsIwPzFj8aL4NdKnsHyLJP4djV9FHimhPvBnj
VTY4RO9N7LpITDlcch1k77AoVUsmLwmeMZj0joCHe3D+9GVl5RnoPQ7ukCrM9mR35dtTmFBerPhe
iWtlnwVLqKyQZGj9yUMs5QIJo/V89wa4Iv+nP1gDbzYoD8YO7QFIQR4heTHoshfJTp0CwT9VMDkA
s4GC1fqxf5H47lODi/vvJnG6GaqpOwDUcvk4xF8qv67glAahIEmHryMT0o32A30GTSYoeXwhQ6jW
ZRTKrT2g14VxfhdgIpxF89buI7fjFlIw99Hg4wxxEdR4eVffhFdKtIGFAHIL4Vyg3V7bfh1xtiOU
w4ZKbUaYRNAGbefrmqw7VG4RpqvUawQsQvIunJoyKPwv6IMIg4Fhj/ZV+xlFxjIdndfF+vyVAx45
gf1xjzBhmVgk7fCWShCYXxes+sJ/KN28lLDZy6RqwWtMEzC9310/46Q02yGtfUe0D2AzKNkAFaBP
9axXjxt7ky1FZobgDyOCN4+yFhcZduqTlTk3wxkRPfhuTGMjcnyGz3OuqTl40KY/OaW8nGX59iit
gcgESkXGhHHAZ/rLDNgEwRqoXnHxqx90uMl9LNVMTA6lmvbnReEx7iLPIqfdAfZda4g7WvntvXT8
+SGibWHAfKyZ+p3rJ4yMXTZJLo3wi0HhUZCJi87OJZkGl6xfQV8hIwPZ6SYPU8VS1xIASw0xQU//
F6A6PB8wON70Y+Dkn1sLQDRtZrarwTcnVQqi1ZE3zTsOG+2UoLrgbkKC/4xwWTF5SW5w42oTsmyM
hh/MFYBTeeJbtOXyrH/GktbF2+dkfA4LN4SgwVtqk4sDUDDZTRpQz4tZ9TX3V9976Onj4QHnyIVx
7BNjvUhqyiutCo3GWEd+W/jP3tBllACmbxW4IdNekl/Xg4D6uvIGWbiDy+lvYXp6QwQfVzq3ByXz
xRV2uQLuUxNWmglU+hUWKaaE8nNa1EeFz6djGoClMxd2oTb5aRhaWQHUpKyy502QK1XvHL9ycQ5f
40FsRqPTOkx0GCijUb82bzBCeylCofeBpxUUtnkXWqJ6b54chftKxwe/aAc9OYPS8qHnTM/Qhc6n
MLj87odAMBIMbinLPzvoVIhDg/ezm233nMa4DffgKNcSUbqd8CMhmxY/vfGdLgMK6+Hr5ZLMenQX
bqdt51rGdU4a7kIpUDN8kX9DYQMYRnrL52sOM6bUJWLlJQJSJPVIs31jKcZGIBy/sW+SobqTeFvz
Zip/e7Ku5+PIDe22HEcVdHc8G+/9Ngg8iG9U+CHsklR6aOtGKfULi7fn+l/ffWnoaBJQoxSzJfIY
7rmx7zwRl2kRxvYOWnto1vAOMyx2E+XrwGD59fzkTHe9afbOa5ZP01Ue6kA0Q22QtGKUC5Lh4EiD
Dj80Rel6708BeDROrmmVeNpKUF65ERnz8w1flu2r/l/wcLNz/uV5VCPK7Yyg+DCh9vFRuaJW+Weh
yOPsWopwHk5jKKSS9fUfteHcEraUvxUSl+E55zhdGdXwdVHzDYv8PoLsq3v5EAqlUMr2iawusWP2
zeMWs7wOJELJ74SLoclHZfjhTF18LuPO3WVSIisK4nNamWGywOSVE6+X3qHS1fq7gAZebAFea10e
bnh4XS18oV0LhnN6fwZQGc6EXXj8OYD3iA9W5mbBZHA8mhgYN9ovlzzp3mbdKsk238Z7Aw8dLgaz
hc5KQm1tDQ8fwJaGJwzDa3gC+1rnIVCbK7i/5sU8Pyr9LYM8XIk5YFs/aQdzmOMAw7w53SpSoByD
AlBtIELHaMAH9uu/CrokVxESQGZwt5pBq5Hb31yVgBcIy+tp/wy/ONan6lbPnQFI/AXc1azrCUQ7
qfFp29QG4/nQ/WikTxsb9JtqCk2vigcdgMyBtmDjQByu+zC0dCP51E0wv74nMorrw0Ex/rFUlvOS
PgJoiOWq1jhUGEklTpu1fDDZzZaGi8PI5ifgOYG7eeOZHFEBZIY7VYtWffmsc2vfH4yThFfhFxGW
oGLOYGk8KB4HRar0spXlKuxE4IpfYAYQ+XyKEwyxh9NqnKCt00VVsczgA7VOGW0p5BmIjre5dBVa
fGRuezL3Ywc5iuz1y85y4ruXV4YzHMbSLMWeu4KdjrGzkSoQDhtsHjdk3Oz4w+z3gwwzs4PjQTvt
2j3tTogSdk6WG3yE14wh57sHiaSQji+Fvhf2k8iuC0eQ0iJCDbWOX9HC3FuvNhb0TFcfY+wkZ9ew
z46Zo4WqXJCQ77GuCSTZCNE4cLvfhFO/Jd+ry4ud25vAeR1hQujt96IddclZJ4u3BxvQA1pkxQIV
v3kyPAIS88HXRI7+und3m1KcnawoweDcQQi8UzKMcsdrXNnvhRxOvh299M4/NDXPD/pxGqDEVOU+
NNaIflOxxsqRIVWzKeEHYYC6sfuVFgSK7JeIUBcyCwVxBfY0LmETojN5HJhLOG0YNoKcbwfY2GTF
CykzEftB+o5QMWvXxa5sPS6NgE8KlrFHxK+jD6PQiqcLt4wVgwOMvAAFudnOoHG44XBx3qw3XSb3
xHpMsPLDIsCFYVbQw8OD6vqLITHmDqYX1S4X/BZ0Idg3+haiLtdjKjpM8wjMdYVm30k72kJmA8di
+oo6VyI+SuCU21449qXvElVnA9nVtumMiHiJkNdzYf3jTPBbwpAayl9xeGiOp2Lr6Nre0AtXO/HR
2c7y/+zyZVweAJAMLEftVtp/tYflvB6qWYqW8hgv6/0tmzHIyQf7PUKWNwggKAkoFQm3l9uQVG5c
VK0XXRxQh8NWhU7T8tzi2yeAv5shPiBd2WsIDQ8kFxpG3MrcG4ebj5/kkMYCI8tvrlYTLZZS0r/j
HiBKKkah4Z3LiO7nErOf4sAqBXfbTD+6NOjhig30fX7VY9YQQi9McQkppHCxDtkmisB+yAcIjbar
4VecI/qSnG3QBBFP0hT2EH9KbskgD7DlN8M9lqvcLZW5Hli+FbSoGtQrM/7eXbGZ/4yaW8mSVrhG
do8o+esV+dBylb9hWhB+0ZHZtYTXIUz2jQUiJk2GMIuv2Wt2TxI1UpcpYYE4PGrmDRIyP9a81D5A
QBMjTbK+x7RxbY/LvWywHF5HhMOpBxMHVzEh3r+sJ0v/SkecBSv6KcA7ZtPepT3wbJlLOswxrcxn
130I+WUWCL2EIBje78DLiEUx40BZSEEKj0pjlGWsVUQZojIVzCRS0IibDyAJx5sauq4LUoDdQsyN
iBY1EjQBhHqsNI9q2Ir7Z1+GxDKzAoptBAoMpvSN1pbwo8qOUzL19BmI4fJn4SHm7J7cI4Q2lgiN
tR5AG3cwt2cySbdlLGAp9Kmqfhf6q5gm2hNa5feDbWmtGlCT2fJshjS99k54NiQSGRF60ca4bpiE
+H/SiLq/hk10Ppfes1fVmcOd0R6yJvGhe5i0IvcmLfO2DNjiOmf8wqb+XyR1khNHR+VHBrpqU8Jl
CLJAaa+5iF1lPyB97iYMKI2qZE2xpby5gSMKNHhA+tSSZct4FUtYqWceSc22Z5W9ensL02t3YKQV
v90Dvuwh13S/6Yco1JN4t95kJZDvQlZCOM/CLOleiapBzezxHF9CM1pR7SS4rbjoSdak9pMUzmCz
joslb48hFMYq7v60eCt0ebOAC+jGke3jSM44pi+LdJdShyP8rCHmcAVhPWKXPbT+KpUNBPOZ3/Wx
LJr6hq2tgqD0GKbdl+AGEcrHEvxZ/S9OqjHZYWQ6JEP3Y4SKJPOh3ZdFladTXA8QpUr7QvHrUT95
FYXYzxl+DCtA++Sic6+n+3LaG7jfy1lv6LYgIJGR1uHAynftT4UYAYiNdsV/MEOE/1T7HdzVdEAe
OcEQlM1OLTk3rHpfE2q7/1cO4CsEnzqt7B55Z32By+4QmphYZPbjDR7CD/iOhGW9TTyMtW5s+Yay
Q68z7QcCCftN0rqd3t0rUY7eM33UoQQ4f9DJVj0oMxMpjmpkkvi4vKlnGTEhytUDYrbsYfwFa6+V
2g4WMDaRrNo6w2DPxmW5WlChZlM6v67p52zXB/SlT6GNH0G1gox952mpeyijPwaPjcP9QCpfqAIY
IeUyLXmiKdV46sbrA2Qfk3roFM/kykZZOSTkRBx6WMeohULmO/NzviuOpGg8H040/20rf0ONJLvI
X9nncVl4FtW/KwUC0YW/FB0KbWNp2BL7rXU6+WpZytBSZE/fCWs0OHB4bVcEdjjSDmXZ1AwphyNN
bjVfDXm6h1z6G0VYrj8otOGsJ31x37n8lVHN4yUHtNrimJhvi1j+dv+fTCZInF3buA49YeoMC77C
BXnMRkygK72R4Acwe8HNgwhc1AqpYrvbL4NTqcputy5YOCIyHB1vPiq3fI/uc3OvBS0yBb3fqG7G
dMGi2t9DoQXRTjGHacsN8AuZVJgMWHMKkpVaA6x8YJVQkxnATAEe+GsJT4AdWF6SDhAEMyqz+aFS
/CYO+8fUVbBX0UFxnP/kXp4WQcGi0M7Jii1RUcD3gTHAR8uQlEV2TtpVOhEFkisy7IghRlWpBOlG
eOHAXzgVdPk5LMoObdE5Fx0uX5p8S1UN5yFNQd6G4mQDcnGTIxRGc4uclumTFDCYBRwRJcY3UjbI
zgqlrGwXAn8scfmI5lZ6OP9PZgRW9PSRTcz9idY/d9pBUsr0S8erkE4tjD3pLJc0XVwPUOevSEhj
hY7O8PEe2BQhlpFRV/RZvUGo54GapIZT2p6zr7JL2RsqjCVLhLLmqpuX+6N6cr8dulbkdNe0Md9L
VTACz470OjEVb9giTKOP2hfbqS7L4JYEuwiJFhatHuaZxqY6U4OUGGzjLOK/nRHXAntCkMgdLWf7
P8fZ+w2rsnsusFwJCm0F4e6fSayr5Uyg9xzDhGWRZMHFOVOjdZbMhF5Wvfyw5npiSYLaZmbZViu5
exEIbMIrjUrB/hboIAiPw4vKr2DNH21BkzMswgINqRnl1R3i2XWo+Kci7GsRGKEK4xh9xYFtwp2v
yq53uaB6tEsJemqfx6N/wHlDAvsm45z+QqPwh2bxKX81QRXH2bbMO5iwHhDoBtPcv9HGzrZLJHut
AXRzat1+AfXYNsF/xOnPBHWPk4nfh5ieMYyWoxWN81IV+OBxQEkYZ53vRT/Kl/5l3JP/mORYlT/D
m6BL7soop3xOYQVQNWFpO1/FH4VRs1I2HKnmHkTwGD3yyMxLTckj1RJLyUFnhVZJ4WoL+7Mpkl+y
t8/7ic+51tqNfdjIITCmK+/crKBz+TJ9aiewrdI2Mw8XzGpSfhzoaxE7C/97T7jx3U/2oEOFbAEN
iB+4wzK+njrsEYeW2/Q89EanBL8cErfcDI1noxjJu65879EmkT3pCUgzLxwb9UH9+xWeLx+ejmRd
sGMlL9SLVyO1nKsaqExAOT7h+UJHPrb9JJEOm+Ngp0Z6o6NHhGT/d/grM/nozXDlXd/XOVsSPR4S
+xZIEqM53TivtaVnY37GauRJMf946KGVWiQJTKLOVC8u/sUJheyQ9YPfEKa1dhbvZ5cVfuUrLgy6
6epBVYrlNQT5vzPCWNEzZaiI1JgDQfWIENOG9lWn/vNFlMmYGfKR4QR8dz+24KJf6P9tYoObhIIn
8/nkfB6S7hOQC78aT1ChlH12HtWS5ZVDaF6gsLAtVg/ooj4AdHh6TjLAdDXk/56RCY7yDqCXO+Vy
hOMB6ADhyE3I8cfhut8/lHDWpimpV8/lR5Njny32HQwsSqufatr6IGOZHCLnkdrzXYYDXuquAlKD
9G8Lf5hZNJ+WpZqT+YNuNiNHhd/AOKovzT299LQEaVRe+qxDAtEbIPwH9xgRovc/DNr0wLdeM+aa
QxXOneow9ipS/Ua74thBAG6Pq+AHBRTGTkCHxBWtNo9jid5te3yrAbftgDJfpApFf8i/Pztu7oHG
UzHYMb0R2c4U26brdDA1AFZhtWwHJEzIKKf9ZemYsuPWKmaDLCzcLQ62g3fWx1W4HgchfYTmfRoe
OIWF5gh6I2+wCoJvpiiBXdhvmJ7UPBPMI4q3ICV1Wrcdzjc466A7DAdnA4T7CIYbHnTv27g4A7ya
48KgHs+/bXMhoDD9J0HYS0Mb4h7FVYjA4ZGyxu6BW1Oc/tyKQLw/RNSPTHDO82bKGxWaKhX/rKuo
N1LtKMx3ZSS4/j/UPX5BCPPFdrsWAEqTrfniya2hBdglngDL5iSvkjTfEWdZFW4VUBudYOK7Ku0J
t8H8QNjKbYrReZwU3ckLs2me99whG+JVzoAwfzvpYBnC20rKJZCQ/TXNuaiBRDYYUpeqGzCgsVq1
fyDxqhgOQUOsDRS2rhOQaPpskcPAz7abHdRw3z9L152DAnNFrXRTDR+Bw7C7QgBvGHAfS4nSmMiv
FFu8wwsJe1WCabXPHqROpjenFUVlK2i5+n44Fa8gRg9AGw/UihE+I5kB0/ytte3w09IIk5kExNDy
JRrE/G0JYb29B9Jn3CAn/r9WHRa+hrRCBEX69G+0JfYC8ZCEsTWLRXQ5usOUQXnPR+DN8kCZUdF3
lWjXCaXITwl07lxtGb7A6BJRydUid4faHA8IzZthkvX0G8HfX3HxEmAJGbfXVsX5TitG9sV896CX
/GnfRvu4NemB9nJcsDu8AAF7JgIAUv5N7CIQpjK3yzB0RNYhlh7r9KrzuqY0vc+pVsmHsQUV4BSV
37PfUNagVy0KuXVvWWswLm95Z5yOHVncuKXvUKVUSFUuJLyG6GqpRiY2/W+pwMxKn84aRrdnMW4W
cVXVS4itIL0JR4CqMaHIFtMYYfmqxbJjQuDCpEgGveVjPW4cDOLvwJgAI3aIDeWmA1q4Bi+u6vb6
AZdrgkBoQC1RDLbgV3jhXodzDHf8a5t3ymSFeplhL6t5tXJS4e4yQJ/F/hi5g1t1KZDSULfrpINm
KdDuNcCmRrXSzrf5iMR6iwrburWQW22Z7JcGEm2///t49nS0mQqlZkQBmS67HJzHyRpFb0WLJjyS
8M0nqG3fr3HNR+PFP+xXDUP5t2kbxVVWlbCYXyAVQgQiDcu8NwSqx2/DCFGmj8VlZYzSOXBScfKh
fnMB8PDeALLU0ml6MPFMiHJiWDwa3+i9TN3sXM6/kABR008vW4//zUkpIQ6Vp33+l3YsLg3NZV2y
QyNe7gMQ5AMOP5RZTn0pBXGjR7QDbTmSUodghAkLtIKUINB3pBfJAgTopb4er53XSg1yKYv8eOXq
cR4SgtmvsRsOjg88drTKlCnXdxOjn75ljIco8RaxtLShP62ZQ0NYXlNLLETVLs26oubAnWmwpdAX
XNHPsXPQ0QFImAxQsM/U82ZMhbjZZ/y8bwT7Yx1aiaanz6n9UrI6UOWq5TdHLcvjL342jNiTZqZi
vJQh+GV0posfWdzPdg89EkQEySsq2QQHj4BnSQs+IOHn4aI+IGjcJeFIUk2bRMPaIJB5V/kZEUXv
shm9fBrW6x/WUEkDDsBCAjzLoL1sdl02OhOE/mvx+ZokJ73On4qE/2mPsCVfQYc8WzsmQdvGhV02
HSATikjkd0VgtC8DnFTcEjYLU+5rtaDYEIhKLScHiCRfYw2OHRet3hIhltnfGTeiOPcO0wN14BZx
gMA++u+g+cVDI/hrTMmJf7z2z0Hash3WuOfYrd+KOIQ7JmV4ZTZqx1fmYrL22BKKSbZOY1/mNZvg
6quAqUq1zJbMEA6gQZTg7KiTDVYqgWoklrJ6yQhTUDMjmIwYxqrmomaLhkI9e1xHYGokQ7wbOCsx
UvfLgTtcX+IeCYmfj7nLSDSpdQj/zTo/Qah9ObxAkCVKAxebNJn85BX5NAR5D4/BRYk+5UmoL+km
OTBjJkk3r2UrwAeWHwqZ1S2s71yEYJrI2+FmtoicqcJj+gVr7ggAiisK3Ey8ErNO/gufZDHfNrvI
9kGxi0+X2Hajb+uMhX7F5a6aLwQrCa+TFei2YoazEeQXlhhBm5SxUzpSZKpMhqoj5VBxUctjPnF7
vcGDpWTb7A6XU/eM5q2b5/cfdHA5W8I9SybUIjqZ+YHb6EVS75UuMNETqYMhn9dir4A5xM8tPpgW
mxaP3tBiW4zHA+i9IBkoAhTGSaXfwxB8RkePE8D6XeXiav2PRV+SZ+tGVByH7XRhzDYdh+g83n6d
Zib/r6IIvUkkbsHNIfgjgUK+Zni/Au2NJi4XSM6iBBpTbF811aWp62bCzRR9WstPQ27wIhRjFH0y
TYQF7zdt40J0zAzm21HVCB6jjvtetnDaCLs+foJL1XzWiUpqoDVpzPjnyvMkJxXzCZzf9VR5Rlf7
a1fRM30iG4c8dAStDmlDyZYLW0Ak8qcLBj6F7HnXjaQbHi/OZJ66oZJhpgK3Z5atkj+82wW6uNIC
UXAFgPaB8v5kfl77ZxE9ZcTZvCA/STwy6NRbZoCGb7kUeVIuvd7zKx1oUFGbce8nrAXE7NIigWRx
xkdxmFPWOhA0yj0TVEUf8gZOT9MDHbV3zSbmCjkv8KLyQo3XmjqAaRv8eAlz/2DuvKyrdUq5YO2K
FI/PaUuCZ2I2yGENb9v0q8vR1xLt9RGcyBeKHKOLTqy17bP1t9S3aKgXCqGLcD/DhkAcOPTsyiDi
LOBrXOf52dwqNmiO1MvNwB2uy38T793Z2eU+CK4dEEKO9FtVnLBTaN4C1PlbwDoRj30BD/xhAuNf
7RGhgk0VUHNOJP+WqeW/CvrKW7N8les6zgplA8VVoC6j4m8hQih4FKCcgkyrFNhNzoxcPXzw5r3+
5sP4YNpvCMfjwTHYABWP8ZxAWgp1wO3YeDy8h5RCQxX30DAMq+l8JZcHfXy/6/U5vEyUcr1aKkZX
oLC+w73yEsjADsWLqmI8xjyLLpwF+6Myqt4zWkwl5NK5Upr3Y2zIEX7xdX5ZHXGcfpLYkbKH86IV
/hA3/HkJFnXE3WcMGcM1RV/OPrQAM/96s4L8BaJtksdNy5GhdY+umzaguJIs7TzaV+cWXyqeNTWK
Ytg2VMR9i0sP3BlTQ3yg5cYTmfhTz48X2ohCWrIloz4U+Q1seSv0bxORhqWj14SoD8GyFRRt1R5L
OobFitePS+AJrm+hLpdyfsabwYZsJZcqnD6CebyCRsKmvkh6ogHFfuLbXYEIHx/88Sb+8VGvh8J/
y5/3/aSZIDzS0gVcYo390OxEfcG4/Hnm4UeBaVA+SlEk8RJ13bLY5eS/tEecGO0iR6ajJgsJ5vlq
tlYak/xhgNKa3SlATrvCW32FH0hSGcVpxkmrUkZXA6ZAu3eBVYICBbJ2uyiISJjXzOg6xguPJ44R
D0qDw4pBoASbd7FwTsRIShomOryAn7rwCGWuSlEaydkD/mqmI4YhGYOrnNZYqbc53n1wbreHUEUu
CF0ibRYpgHSVzxSzdSH7yUrDVzFr76O1/jwOoCSTZ4nPBi3BHtliuZIt7TW5RwW7E4Rhkehdbkgn
PE9wPbtTys//U/yV7qkvkKjsuZCflkyHVK1RcRbxVZ2sfsy2jcZsOZsL8V0pqdhq0FJhhHStyFac
F0FAi7kdUiHJSU0SpNaHkhsbR8rTRvUzxwURPItRkCjN8t3ey3iO/L+g7jEYph2gGXGTFKgcoDGr
DdWIy488qCtlkt7tc9Qab1EzHi70lKD/tgbgSP7OlR+fUHo5oAkjtTGMxyGacXEVpSP6qhhHkNkM
9mzHvTi1LMKE7B0BiTZW58RT/AXfI++wrVi6TeTBa/poDgqVjZ+Jdt30gXNjE2r6/1ZdkZK/BNvz
03ImtewLP6rA5O4RwkxvN2izcY1WDn/AOnonj/wXyI7bZBeoie5S0+TpePf6haIRrWXeOXLDQ3uA
gfLAKQ5w+CBcMo/x11fqt3m7k7WayQCLgSwrxPDED9/gu9+NbWJ/rPlXdcN8wP6UybTKMZizSRTI
SEqjdBEtYciwMvz5y1ma7KNLeniTVaNt1ea6rduDfOptx7uCia0nMT72YT5woybwGmTioOebAsk6
KDYk0FcFyQtl4a3dNpUzSkdXD3w1aOXua4iF71GcGqbNjqP2JYUB8IU4XO07JdDVb0wQQKOne4lj
k8iyimr4qsMBNi8IPQN8aF+pCYa4/GD3GjojqkOFpPj3McnG2mTlN3MKmg2C3/1vPF2H0WN6r/LH
tKQy7QLzpUV9MyMRShiVcFiCTwUQVjYThqvnteC5jj6gYmbLjyaWRxWZL2Be3K+wne1FKMfrTofO
X6IEyWBmu0JzMTcmQmaWkgVeZ/EkdRrU+0j0C5mJARljUHC1OnHyi9P9QtYlI3fsx0dLbbMP7cF2
OPxKddlaHfkDyQfhUeyiMELP1FqYk0F3y6GoC5Gt6+/3nmfglzh8XY+2k5YI2QhW7C6Sg8wrOfyr
ddWY054EthQiIeYF0bG1U1VRaDI85l7XNn95Wlc/s9xwcCk/3TY3kYeSWkXqFqkW9EiOd6E4vbaY
AhHbFjKv1ftOxXnR55Y9Ez3E88agTW9k1RLq6kDqmtiee0uZx+7CIhjfMhQymYGw5oEEnd4we9si
5Yf0cwLPpfQrQD0VbvUPwoL5rcw5cDZXoOAinq7SRlmPFGHbVC8IRhfRM6fmVrhvNLRdBzBhH9CY
1ASHqXrrYA13Y4WjgAdnHh9tACZMamOlsKSRLDFwR0pfZq95h6+DqzlhcH6DkgRApcneyStApuzp
9Uvf4jwRGmu011Mj1jlcB/hXKkdJjv4yxRXL2rp6hGbjgCPyegix4VTmAudflTvvarmbgbUAkDVS
xvrqhmAnA52wED4fyURLr3wk4XeGtIlS02W5jdzWE+DE0VubbEth/T27z+a/Dn2XSfPvrwvuuQ++
hnRAnvgK+ZiCBuMinmo9PqtDdnFr8KQJbEnmi6kv+zTzTCpUdQC0dcHUbGxOlWReniLwf4885mBB
hUhahEf9xNiPJfWnUgjQa7BzRTou2cDKN8Wa44s+U8ajysY8e1P1It70NKCmf4jj4+MraKCmPN50
5ur0uN2TBLObAosj5s2TAhTPyJKEs1HpZ5ba0dN5ncjdiywBkTXK5lGjeP7q8IxO2iIV0WlbTrX0
I9zn495xsooj6H4NZtiO57y6Samw0vnWyPHqNU6FjhzCsp4M2Kgh8/WjYUF73MQlDDfKiQnBzmNr
PpAaG3VY8VNQL6G6KyoM/qeb9jLEyyfmMsDyqQcQTmqkSUsYiPX5n/2HNAifYjGmlcyRir0NxCEP
iNZh1dE4hzwZSgopbAS5Niym0KLL1XKfUWAHZr+1fo0WLnMyWX5RjOzakQw67n60/pORhBv1lfA1
sF6zDLpv2R+upU5svR0yfvCkXojUx2KfXk5B5tZMGcdjoJErtXCLI1Vi+Yc5ekcxeoSeYOw+/0DF
sBG5oqRjmp05m87636sH6g2T8OW4szM+Fu5zc04/Z8jsd6IEnrTkFJ4bfVm36ERRapSfQP1JTv9k
/g0Cc5uAxVJ1W9R08elEacJPO73No7cCdkfIARvzHdwsFivldg9bYjCLKIzm8fIf4PqZ04fzndNm
ZkRY7ZiepozIe/qsMkmsD7Qkon33OTmdQGNlcm/lEkb95gv2cW9YIb8AZAhyr5az8w+q1hZSinL5
9ELaVCdqYMOIfthQxikx6pShmfuTGUdEdvpWS3qwTk32AUn0Pw8NUGKMzwLQs1XDd/kgdrkJ1U8g
1AJsImJPLCXwHAoNmns6tct0TsfGBXHoR+9iDDEyCl++mTgD7CSb7n2NJ+M41+KEAMBIOIC8GvwF
hWFsbr45MAgbbwR09Pcar9FrMz6+9ox0CvcSjyA9eJq1psKPBmcc6hjegJ1LUXaVVJb2WAIv7/M8
9j+MxtU+gzHLCC7ztrLK2MqQYsBwvRc7WH857SIUFaEa2N8LF/5DeGdaDusqrAp/rej3Ms5ySWEO
FIrYMu2VBb/Pd68hdzvElBX5RUZ+dSAn/1ZdK0iZMl6OwbI5TgnmqjM7Tuyo58w8lFTF0QhyyR6K
Ljsc5uPeYEu9dgOtDrh5yRcUqQNFXaROxsQu+nSg9O75v3XbZCUJU/wmPOGnB99+HjwEEli9iL1w
ju9Yf/XxuLvs9SLKMQYYHh0RpGtiss/nXZL6SjlGhU404VJC5QmCpE+dujffodgdJT2uoDFisgzs
dU42SnjWv5WfthRK75Zed74YM5snMLA/wtRVkBUeaTCVKFaYhDy96M5yyC9tjCJxLEmFDnN4OTqA
LFnK+NX1emDzH92gN7yfGqVK2vBnmeapN9wizSR3Tkf7DSBPQ+wjNey05dScreuUQ3FXsQfFesce
VonZoHKwo6Q6iRypZgA6MULUwS1vd0xapTfqu1VICUDf5hnB931Bf+ZGQtNrudHTqWgOy/uD8aZb
IKduB3k82kdQX0uUlFIm8j0ibefT0Rbuv/9ChjJc2aGSHTHA3QGBBGCJOwYyuL9JT70OD7sO1h+c
HlFwwgGrR+SE7z2nFvPCaLSeM9dUVM/ftzw0wxop8a5kd25AxqIreexsZKf3cQOkIxAnAKc1Ncxc
4JQM5+8FyRxQG8Sf1TB46XhPDCtOK8POXKNb+t5JtM+JCAAxM9YHrkw21V87xRlQiWU20MUhMLIA
ENNBDFpW9yDMrQpP9GtmDIFNnJRv6/PUHK4CRBodsPHbnAFeH+EUOmKh6NCiDQLP2H6COTHSmmuU
WY5i+a9bPJN3LwLtWKKzKieX245DRN5EZqYEXn/ohz0lJU4xcj/lPmXr5ZvgH0AT3DtA1PAuJhKx
meCfNaFEH9QMrJjTWbT949NskJT57npReHAn1rCRG8Prr6YGOjfDlMFBV8OzqQWMoq63YC+iJ6ha
BDqdQAFeyBV0YZ0voUVLZIdrPevaK88/vg46+QIg5GhXKF7pdJhhKOdIHwLns/+8gigkYZRSESH9
h7+46zLzjbZiZh+Kgdj+FLUWy/S0g5Pi29Bvz6IcIrZ+v3rp5mLLVv0xpW4W3Fl5dp3oEATOGQ1c
oiHB5asYaQQ6/l8TYFRfqA5qAl2zT0RjaOwlNBsn85xOCH2GoqiNRES0wHC/dXAdgESaKvQ8sI9X
+xZq2bCspabupIrXwCyDMK05lmklbNHIeyL7Y9TkP4TUNiYySJbzCRYMfVFySxxoDqCQLsnXg9N0
27DYRTm4NKQn2hW41wfosiz2Jq1JH0ldbcGS79FRhfxG9NYkxqqR4rQlvkH6u7x/YinoPkESLWfp
4UNbIb3gjpTa0hGBCWIIMAUJRwN2Bncv8VOBmcS2a2gFjjIDHuivZqWf3bQE7/kW8YR84Tlx+s57
S7710nCmWo5OuuWHyXYxWbnYnm9manx+KFQjjpHyYkCr++7G4SH6v2ULx2AyN+t/BFXQvVlLySh4
MLUQ5WqpePrbHR01bnTZa9JR0TyWFKDWBPesaDRv5Jn241+6zJP+ERups4kVL106p0OYCJg6eTd8
HTxdZ+T5VGZ7qHr0p0XR5rTMSZR5vfujW4C+/ohPA9rfIR8g+y98DFAMqoKbu9cqS9bxAFgT1We7
RPWkA2ZRuC2jKSRiccQOhukZZ9QqfvG10V6vN1a1E4ce2UBd5zdKX0LaCClyzVOT7LWP4ZVCTdVB
JgmjdV6wVvVCDb7y6667iKL9xkyLKTmJkjVRaNll5+IDgf/p5Pjz+8KihGEw9RIPQBIx6hq+pqdS
DrAf1G9aohogQ8XNKPIPhS95JcCpWEEpHBFN84v4NOpATBzZFli8ChVhSRTzV3bvUp2162rk7dBX
WqtGTAgmzbVAp9uNgQ+kvAGZZ3NQhqwJz0JWZwCPjuMobWOVlzSMYJPMJsr9/xEKFP+eb36K+76O
KGz5+4UO7iZqzMh2Xgw7+qxwRZQQ8otUuLFpjY8C5aYte7EPX2+431Lwd24WbepeRc7mm42jHhRS
fnfGoxFUi+788ijvjFATZfZuxS08aqLJ/lo5/CPEjYYPZOC0C4CR5bZtTeDuhwz380pgZ6nJimhT
TGYFWe0NU9CU62GlOAZtgperzKB1pluFhKG+DxnNcSLWbV7aIdmdD3SwSOr3v5CUr1qsDTN+6sO7
kmEcCaJWAS/5ohD5cyyyg3XzbhMOuyMGYNthUKHUt2h7+JHE8QVDCmVzfosglwmYAiDK9mXkY9B+
GWmEfPPVFVmWNsNIz7/KelKWBKy0+18YFpySaoW/fzHF4iz/DExfvjrFxLVt6+mGCT37uXCTuWhh
X2lQ7FyCxk+Ow+h5chA5/Q5oCPsq25gey2q0+zPx6R+LkCoyexUOabrSBhNecbjVKSfZDWOmYjd3
WaTBXZNkEOrvyMqptHjuDMYgdOBXAKb4VN3STDgXrRTwdWTl1yy0fWa8plqafY54izCANbvcsvEc
93qixqSEJxmoBH6aZPVoP/HsvuvbBsg7bP2fAnKj5huIp9LCSXJFhOH88PJmrnb/Tot1MZKLbxrJ
1eEMlFrIhNO/7xU2aPJcC3zXuQ+RFpBDkOJ1OGST2mvB7ZVE4lks05wnGCqcu2+Juvuvh4PbcJ5O
mZ71fiHjOXrspvI7MXo3R+t5cvStNEzAYarXTlJrvLRtnVqAzjSv/8Eqi30srELcQIo9z/ildREa
Vh9rqlaYclRFW1i4kpy3MuVs+hqjdI9p6+i7jEgs66ncZvEgVhU5PH+gxJD46Fu1zsJG1qvRT0HG
ya0YHdINy7fVFsDo4zM7MOGuTq6WftyR9vx4YSlnfjn4gXXWSsw2EzR8mW55DgAEhfQt9LHx+fYN
5e3v9nW5dgghlWxl+D6P1x329JwBDH6RGlkl6v3Yb4Ul44yyzr2mqEJAC28+sK/l3uQ3fZ01nzGf
h/GGo+E4pCKctX5ucdRMo049yNHuxCGfp/IeTwdsbTi+OMbrCmBiIUpRWsWcEkZKM4YhQijkk48m
loQPOj34Z0tLxl63fWQ/W9Fmh3I3su5RmQfXNYLXStZbq8nb4PuNJpLa2XmYupdvaDPDh0sls8rr
zRUaprpYhiDCX2V/+hLTmtOrhjzfNkJYiyd03uwhoX3fmlPkdmsbUD9EZh/pBDo2wRlxrrO0c8TU
ODaqgqahhV3upIzUTXNb9XYo3qfXqCbyCt/FlHA4S3+ODffNnls86T0CWPsqBK1e6S3sBgWebs3b
SlZ1XBgBpaBVTHffgmdF2yqYeqECm7iBPR25UwVu0abTcbRAGHBGw1IRgGCDo28S4WnIUahoe9FK
W4+dVUVjHTTPHAukjCTXAJi/wpzi45pYp+P3xd0Fnpplk4uH6K1B5+lYtd8vD+IDp/zzwEYbD7a/
CVs27SQNvAti84gccp1ngngojReecMFgzXF3UXhI8yJwMuangxiN5C5LHGQmWI+qGg6RN7R4Y/0Y
H6bg8l0wqxBF3l1GfxhZjS2NaNokQkZaE0lqi5LYzVpf+ATZ3DPuuyNU5ptGrRGehu0U4Q2UNXPF
1lzqkl20pcRpvsTkEjhbIbYW76yXdUigiAA4aG/LCl3u3iVO5ZTFcE6jbXAiA8M36hrnlV/EK+ef
2sF+yVemptKT1csAobIfxsELLL/F8XpVwdJeTxcHI18TRAZDQv7hgrks3wIlwpUmnSyy8astpdJn
DyoZ1vNCO0r7UILchnbJpN5sllQedw1QFJMsXVmfTY1kCOswtwrffJ+waFbhgfL4knw5ORUMtz7N
/R8SsyhWdXC/YdUYkfH7tBwp2dcfO4CW/aw59q2+jeoKb2YGkkBWegJ0+lhtPZwQBqpv/yIkgDk5
T4Ku/KFE4jDF+6ajBnh3fehUk2qimFTquZnWSEuhh+FaYj8dB0g1PEqUI/TsePg1OG6BkLrdWmwW
N3RiT4LeP0m45Zi+Cg3ushrxRLgwTLFN7dI0yTt6JkozmvCw+B/6qEJ+AKTHuUjpZARtL8cBgJ8M
RbQY29EY7kKiwuq/tieibtZ4RfVU3+6wEH1ViWK1X0EuzeXdB1sh6S0sdS8I26wLGbuCZn8oyT3B
l+Za3NFZ/7ULbwGPDkE8ztQSl7Z7WR6df8LtTyt9Fonlq+ikBFMAo/eOGNSgrEhps1fDT1IlzrU6
jlJQZQhkqolG19QAFyj7THO8AeP0ta4HfY6ccb+uFABB257iE82IwfiyvpdbQo81/v2nUIedyos+
WQH2slzgDWNZ2qvIOBsEKHGWzZlfJj3XBPbelDP3xPv7uDVtsV6++7qIL4yLVnMaHuIgPlpbRVqK
geQCcxK9Rpq5o/nkvqt56TjBjZSa4pv6h2zw5YHQhoXKvhjsqGrz03umx0APsFj/A6PAHvEfnuNp
e6F0ejvWEkNcMggAEVBmgWWG1UzTGlQpYg1KdZZ6vTKBO518lNIGCQDoHZBn2SxzaOZmyBiSXDwG
Pt9HBdhvEa2ks+V4W/DAjf/CvYMdmRFRgXUwN3nUFFflk06wX/dr7+mtIX2Z2+kSf5CqvqaL2fdH
f8f/4VInRZNzC+zjUacB56PZulry+/2UrMGa2ynkl2602NKYX3hJCh62DTIn/8kSduM7I6txuY5r
RrMyBy5NkPRKNMxqUXnKnBe2q70hfiPOG8Eb8l2Ae9uU2zHb9BbdFDQ47S94+DwTkLIG9dZ6pseR
lPeiswNVSzk8xAAgfv29zNEI6Qzvkeek6h69KuG/xUpJqOsfFElsQ+hoHTfePNvKZ2UQm45cSUDP
pCPUaU9tJhZwRXbX0ebqaSD6uY/XIcTauARzTj9AJ2dzvJVYit2xx2HC/rxYiOl98PQ60fOoxX02
PBrebx/tdGosNkdG9lSkAiU+we7vQCbl717GCyFq9wZYrMGj8rfW9XcyO2RQ3451yiiZePZ4foKZ
SF3yx6ACh6UgB5T2hMv0aMmBm+9Br2DNz1snkZBG+D0Ly0pvC/+bfaF1GYYh+mdcY6/nwfcE+axh
Eigr2/JI3wX/OUQwiLrV3bPNtp3jeu1MIzQvcToRyvx9XABVOJeJCBKaU0PmhI11iUJKYSLCnOdR
CxjWuqkBNWvat1nM4iv+ZPFYJuC2CK4zBTYSp3dxbH2pk6hTLn5QhXt3ZOLzc/Rfv55JnUMCHo3O
4tkO67eS2yIkXLmcOQZNT14P2CPhQlm3hMMKioZLtP6S90AvkgCrBJ0kUON8+s1Ay5feeIckrsnV
bCxDu34UqFUvfqpops+WScUBxIVgtfhE7nSgfb8IPsmRArxMKR4ulrNuG92GjiSJdMWrliRBlGDy
qFUzBDGtltLWJ8zrMi2A4QTDq6SodglnMTLIM+pHl1AqkfEySM+uMEHZaDBvDf3nTdLE12xJRRCs
2m4QWUHfY4QWQ9Q/2PQEsEORgi02X1rANQ9yPXnZPfeazF9xRtRW9EQa3MsETqd79kofa5+SmkUi
YKbTjSOjJCvqhiw1/Cnc31pem8XAS/wZiEKhu2rGPp+a+XhVxnlhu6ULUbWPbxWqzIC4ZYy9hcMO
sCElC/vP1XXwEzsC2oK1Ibdp6CqfGJRr2S1z5J316wNyGim7oTyHwe9lOUywdAtWqCAN3rD1an3V
ARTUuBVkuuUywKyxCvmJEK0+zomgOhyPD6yhYtoSY4AQWELEeQh/Ie5A5gPB9A8m7IoN1i47Jj0A
eyIIdc2rROM0hZ0qVPXEZi9RPWsggXBA9rBN1MtzN7e0nKD7+QkhNiLQPdzTluo51MKiaTIpcJxF
WWXKP3PjlLkVpgZ4a9pbIz9IIHi9B2o3+StRxFhvh0mnAeZSL6d6vxM037SUUgpd++JgMMZZvYcd
rxTsJY0aSmz4q2p4wNN78NOROR42vkTXoImIyNUJg/EGlpwdwRAT8RKSp8wzKgVsKVVTRxfTLeN3
gcI0S8PhQ6k6VuScA0IE2y5/cY35LMKciSo5hJuLnm9DCFa1mb+jjS25rdgyNuyiTGz4Xqwoyxkz
Gv1mdK2IG4Xa1/2wEE7ZbimKYFiZgz68kVULuMv2BNoV2XvLdgnLUp1SDO/5VUUWuIOxuV3t6zH8
Kq7TPFsw7NZ8DzgaxzFL866nTWsh4TeeAYrHMp6E01oTdWiHIU5S0+mY0OOc294l70VBv1WJ1Lyp
VqI9eZM8Fu4jCn521rwuDpnGs7xgue0Q0ShLgjiYWnJ0k4sW7W3Iw1FuVTW2AFi9makfvrFRHvwe
n45wIuQdCaZ3ag0EbQXmOwlPJL+bO3+n/jnXpWNVnvTTI8Ibvuf1WK/TIupLwJbmPZgONsVtfHUs
iw2I+tQNuePHbaC6nfQkmUTQQif1+M8uT9p9SpZtRvzzk2rr7F4Lb5fvdkpSpTyIa4Xw1GK5igdW
HCKnI0W2qY7c2Q6xE1cqnblF5F9AJyPCpNa48kzz8POrmmm2MUY2Gx3YRnV7l1Amcmg8zZRPAdXO
DgS2RTw0szQUt6qkXUT9m3RRgLruCiVG84QmdBuycllYncxFbtgkHVgxiAkErUpI8/+7kGnjzRqt
g/7v9KoTjI6kKc8EjLGstesYeggasrC28r2Ody8nFUqm/7+OrLuUgOEemRIqzCuawlY3rdatdZPz
A6gVVd9Bqs9pd/0jfknMIriD82q/wdgB9bQWIwEqQiFdfQ2r47orhZLuOSCtvK508jdCKUr/aJ+4
U7nLhHLmQUCH6xS5ccuyFqt97uEpteGXBXRRkiFHrbv15WjW99Y/qX8U9BZEjV1377noZP1Yh+Fb
d4wARCVmroQCjvzOsNBhNjQzgFftG4lyS/RRgmOJzCnhwVdV55cg8HFACO29GZVBNnzuhSh3KWA9
CD60gitJCUL0v5b2fshfYODqoLm7qhc8e7r4OVBvMhfMGcHGMPK118BbvlZhnE+MmKvv8mh2ZobZ
X3vIHrF786lLoJ0BJ5/BhpahLlimkhHF0sFFUwMsXdglVVvaVail0oQQlaqxWh1jNhN7asacMUo7
Jm860I1+pKhz8YlQZeOpOssO9CHNJIhGaXEHjn6qWSFsEEKHbUTJfa+mWZPOqat52gz8dXoNxFyx
Nooeh1vd+g+yajWD1/hEND9X83qy7LVF0stea98H2Y0UMEuJgAJScIJBbEeA8iMjAtG9YupOQ+t4
ERFRMGCui3BMrcNovwNRnUrJZx170HAtMtAIlbO4KtcaYQ8oNrA+JufHz4BANWmYdlk50v/2j5z6
4/jBMXv/UR+hoCEHcc2mzSp7A10e2Fv1cGXwREJkreBszwHJC7/V4ScaEJBEdJJX+RuiA/Sr7XFf
VPJLgvPBH+YXeND/Ni1gB0CGRRRWrDOoc6StrgVOUXLl57GNBuLDfTIq+njmNvOdFI1Mfs0zc3bC
kC3Kuf/+QC6C1SxAj+ZK0poXdj8t2QwjT7G++i1YtgyVnWrkoFBWhos0gXDc/iURObclfYO8unlh
1TXuPepsGNm3ww9fDhnazi/cpuaYZK09zKE674MJFiXq1XMIw25l+8frr6fAoEKP+2b+6F/RM4Yx
wEzoXr2FigqxXU1NAJnlZ7jUwLzqVAAetXBrEGCdN9t5b8bu3VuyLLjzP6zAzPPdz5gUIKRRutPA
UZZTVVQrYxQTUX8a6/rSkb6s05xo+8gH69cNP5iRbwAkmO/uCV8GUvQeDYR+SiBMIGCA1nzfC7O7
ARUjbaqe6AXDOCCWPhP042U3Oy08st5wPfq7hxHm+vtj0nss5wGSlQT7+wKX/IOA1oUWM9qXrx9A
UrDCpyIojCwcv5Vs6k/mAD7IltHhbrtV92YQOLWRHi3NQXWUfWn5VzrN2Eu3eACXpr21Ng96DLq/
RDp/7mhZUzu3yD96aQZ2UTusFJrZLT7UL5a3LnSPcAKqq3BjkBheHoz2ad1TQeFclAuYsSwv+oX6
aCWuWrloYTSzR2MtGgO4hVAC9Wavlisl8pyUKiXWNzMnAw9kA1sxD7HJVGuEed5Ze/n1QGX3Nsoh
G+t/WJsOm2AgZAXLnUT6GCSwXDyV2E8bROMUyFZvO6epiRmBW8lughIGQ4xrVlCyRDWRoRpqxcy2
GZWbY1xtRI5bz41l8e4lR1ZCzbHHHM+FMVJqTfYvFKSc0pI9Ngp8VqXsQewjiw2rLQ82kmlcOo8s
XAhQgVX9DmM1BPoe6UM2DdB8m4NeeZp61IYx+8vWERpz74kzgAnqzVnpICf/4ovvKD/PrTyEmZEN
KeceU/1ZVboqIL1aKmkY0UyDNvoBwXBaMUm8xlYF5selT2hgAAcG0Ot4xuJ6tbuVfu8/xHkd08ek
1kZklfjNUVdLCGttDaqsZ6riVWM0TzLv4ykuucE4dAnsDO9FKAoOr5BIVSXwNZQuw5KgjmkoIjEb
mAiMlvADPyJjjFz6ZQaXAjGZUrZzbnGxOdOqj+aoZ4qNzbrcg41OBnytDDHefupK7Deqjjff5nPc
N9obVsJQI6UfDIqAdBUPp02AOdWqf2J2mdqzIL5CmzJPYkXvc1uzgWw4ca6j2f6Yh6WPMWyrN2gG
NbeXbUsvpyJBLKZu9dkzQl3KRSMNLs98x8sVd+x1owPSMLSb4J4+3Yheq3VwQJtXLM0TfMBcnssb
sTkTT2iDC/SvXXdxi7mF5soRKmoI7XUDLago+b5JLZITp7uy1MGOME2Tya4lETVgFzLCjiMqzH7a
nWuIMXFeZydrg9mHZCX9UTPDB37cxE0/dh7mN5NUu7nxkiZOwDAt+jK2kCUgGDs85j2AOqZ59Vwg
F6V9ewT28Du3B4vP/AS4S9sIuL3+m1S65vL1mWX1f6p4MczqY5vVhu+4CSDOOHUEOSEm5b3JJcMg
WUfLdHjSPS+NnhFV2E0sumASydRyJivKGgZ/wrwTUjBDyyrYHRkqAwiTDlKtJjsXpQfh7yMoKPF4
OroW8+qzQDkdtGL317XJ9U5Stbtrv/cyn1kZ5F/FlzBiBiLmaWiBETxMTW2np4ER+ckKFMDKLDwo
ca9n8vbfYV/U/y2tnO1ZIM6fzOrkXaefoga38R04nDxhuRuCa5xM1G1Ou/NPOOllvLAYSdcVjDT1
XjXFfHHM2S3Og67QR2PDdwZGeoATJepewnw23NkcCVd10t/4rU+nnZrZvUkh/w2yDjiHCBiGSDAv
Aq09EinnWT5q7UNOc81GR9ZhXKjOQk+Wa4SSyfp0Np5dVdat/xJfO+RvzF9BifGDS12zD12dHLwe
X9OUi1rDMNQklSXpqDsN67qWP0SSgt91axUBC/q+NpJjGOtfZ/uvL5ABjltEn/DW1nPWedTfSJ+h
59vTzdWaTihdBLPAOKr50P6ZVWuMEmgpOcpvLLP15Q+tOvZE+yX7MCSvpjJt7iehc8dXJtCfBBg3
MW8VyB+4NsoyGbO1w59epotIMnrRHYnAAt6MfQ0iBF9Vf3WYtUnIK9JB9z5ICAkMTvcnpFKCupPr
P7ALk9WwhHw7uFG6v7ZFb+woo/OdyXpvgWMKcyslNUR90fAMntlJPLrMkeA2vAYxA9vz1lnKY/nC
ph0AizgGcH1TAmDMWFXIebphyLiygyZ+OipLeZQx0hZl+BBg6PNj7OVBvzc7TZfQOaezwvB4OCRg
JG2Vm1JSCTBvghYPNWvql7gZIR51ldC5Q7lC+WESUmIux0iJB6z27Vd6A4wzuf5nqHdvSA7e0zCL
AHmqLYBCLVD9/LK6FvtgtbSgSJCXojelxbHmqPn0B19bIBu+NO4F98EEt3eV+EoHAvGVMMVK9Mt9
zOvBW7F/fPTIpi75i5jAZMJ6k2jZOhv+o+VTGywqLxFKs3tCj0zZhkhw0b/d2fUGO6kQ3fJzeJ3S
iy0p4zIazpU41vxstM2GMM/S0I5bZBR45vkN44E97oWjccyZeMETXEAkEXh6Y3YViVUJz+cvv6TW
OSI4IfmQ2vDCaC/SWbLs60nHDNpgzfEMQyscG+rJspq3TkaqaNwNTVRa9xiSWkz5STw7tcrbCob2
ICLHeZ73u1NTiRBfa4ZhpnQtAramAl5N8Gi2XrfR1ZkFrwn8lfbH4An6xSRZDLEtOQXF9jJcIC18
iZlYz9m6z5BApks71W0eVJl8ihGh7wIm8/Uhb6nHYfGOFVxaBowYt2Yv5o+bwBnF+YEuK3pLHsoD
a5kTfOpwd084ylUduFq1pAHfOlai1qJuVw1UBjYLdLF0UEnSaJjsTyI7xLPdfEiel+KUHazM01RJ
QbehLnHjDqtlah4Vcxjx3WTMAug4upetSC1bMQ3fpESSDmTyuaXS6ZAo+RFpWhasWCAdjrWdUJ/K
d4WvL13HUdwVZV0YWl684PoKm1PJdHm9p8r5hothmIx6MwQqmAlLftT8DOcREYUOPqWFheMEX09x
JafNR/v9C4T2hiSykfltsV8KMLqU5mzaN63weZDJQyEHvCIvKWtYSjjemsLgh55l9cbxI54PbASS
y13OXUiQ7uXE2VyZWQaRjUNkvlhQ6VVMRjvFTBF8lJiAF+jCPa8xaiNNHACSeFqKfWZQ22ehj0hI
XoupndsWJgUmrQKiDCR6JkjwpseYVI5x6fhp2v1awL4/Vn2t7sSf1CE58CHGzDN0rz6jdEIJ8WZN
K/kzKKqqcAaSlXcE2ui3NAQM3eUD+YM72DpkDOg6r3gdDEphtCuE0jqR2elLNNpXxe+ocw9Fo5kq
TzTmndnzuX4BeHSpHdgNhF1A+5NS2/UsryuhQxW+Zp97Al7ljG40Ozea9kQ0Z9+TKsf0hjrs577i
vaDC6aYlREBIJo2lAcQYzsVtOLrZUtiUCTX1J/0E0OF27kgL1OWQi01RnhF8IY5PHpRBZ9XhcbtO
v4Ngd4wxlfZms/a+p8D+QoqN6USYj80d8vkbYc/MbYsrg7K91LgChka+e5MIcAHCuLlYjUvFNBey
nNs8C1RJPrgfZaEpFW17Cb2m2JDQl5+Y+xVCcBQEXO2AGJH4v3GX1ey6S54M3ZVSwTdVZVrJTnF5
ukNH2DrhYD85jBWycVq+HM4qmM3sdnb46g84FRNGFgcIGgp6eFwGFQAqzCCLvovF0R3WLDkUEbv8
Ex7duZj/1bwjrTEOqHpHc/ynAMb0edIzmZZE/uFYWiLvAMMwdUZhXsLvLl4V6DPk/sNAykScrecj
qr9aESJDdsp8UbqzKJlTUmiU0K4H4YyjnVlj2iF+ZrlD4cnDj6BuGWjvi0eLfBu45L+sp78JZKOD
67NpvCxA+yRDPkfsEd2hBJS48nxtzvp7xsm7QwtbgaBwzW+qIN4ClhAA8I8K5y7k3ZXqyyjIH4Ty
6r0EcCzziMr9KAOEA+KwUCSPqs67AeHF4A8jUUsIF7kese8JYQNrMD7RSR9gzNXLpWx5fVUEwLEZ
pDNthrSs6E/1qWVH0AnZX5kliIezkYrQzRNsCaZnlr2HbQbj3dbXwwpWI4AKkUstPx6Fv6fRITGm
AEEGexnptiDfO7TNiDUrQpUQ4dfTqJ9vdRQNNvxkOEJsZUGRTKFHmtRRh7jhv50yMYh2Nmg2Ys5G
Vbu8v62gdMWA+RDlnzvpmcEcG6kF1yWlXpnqfSGZ5+6lS+uIG8Z4sKexTDRtHX8LyQZMU7tXv+Cb
5mg6n+SaAhEIb0J86oN4wqm93xeFsLmXnjzY6T3nDH2efHRkA3IVJlCBwuBGWi4bvtSwhO+Kpv23
CZ2SXWT9n7VaG5uVaFsUWdU4gqPQovygBB/pdtE0jO7pnccF1KZSOKxxPOAG5fML6tGPIAdvDZ/K
ffFdIoA8GsK7G6ZS34q+NFhkhJomB56gM+QuImZMd/+PU2EfaNbKUkWdgOFgYGA3z6Ynb5KodBpc
v3bq2MYGAmeH+CIbF6t/I48g61qQ6UU4CcjXECtlVLcWQ+Qb726G0H9CraRbKXUWMgBSVI91h8cU
QANRs17YxNG+vUX34+5NjgM8BR2qimQtG6b7pjYjmxRkzV44qopG2Zv34tSlT5j7xvcLndxwa/o1
QvkNX61oxb2oEnX5WGOqQ/V6bPllM/Vh7+KZnktJMS3cXlTgg81IM5ed+xkEvUPjuuy5cTeWQp+J
pQUFSOZeXjIg4Nj9Q8FX46BnXzuxlI/4WVnQjVr0bM8euITjANxmQ8LN9udQUbue/6v8Llnrx9a6
p0NkxQsFqYminJYDIvz07dNWj8Pqc2kJE4hFdr85TI5VoGKyuewZHlv9r0++8CvEPEf/X/40HMa1
O8yzrdg6pgEM96zfqoRP5MF7y/Bgi/QJAmtE9uBeUPLNoIzK1JDUD8OCMKbMe98hR+iiPhtYwy9y
A4WsmRR9GMxfi+GbrRN93Grfw1c12rKpzYUSYotq+NdARq9cRbblVcdcEOHqvSgY3AUuELDecyYX
4lkwhmqxEvD4puayC7x+dKth91MT7FZLGdjsNvZP3J62hPY4z3zq9lnuz0HhQxPbqrsxK90TNQpH
c3b1FoZj54MC9AtUPzakbVRQRCTH9O1LJwDDkNVhoyTKlywZzpZ96avS7UJJsMMEQaay7KnxHDSa
sJ7AMnAab1O/3kyaZMguOzxT085Y2Ab8ywZyY8EYtTKpx6PrnqRR1QfM6Yk1O3wpUlkrj4FU9/28
q5uY4xx078HjmqUHx+xSwZ/zSxpMuJo2TZInX75L4fFqZvjqkyL0lIP7eg06rbpLHdIyA2XDI3C4
sKgF/YQE90XU+YIoxNlthTHVGpJkcNwKZ20knSlkEsqW24sI7uRkX+okjRCyvqPjgzjaYKqcZX7y
XnlvugzV24a6GsxGQyNI4O6S914blMHrlJvirO96+GsRdRL/VnExS0LnbmqrkDL7+Bq1yUGPCiE9
TX8WPIGnq0btPo54rb80M4bzFiT5DaYaYtCfd8mE3+htEqhUAjxIXUyfxqF6BhQVDIMh2Ofd4vD/
2ZdhhZkETRmSsjfIhTWdk8xIa/FNnT7VTwaKWca8SjVD9ZcLUvGXyr4l6okDrM3PdqPTKovNEH6a
DSjbIUOZXU1acCDppirz1dS0rSp9iZYfVIRBKr+53gorTVtdzCw0kYRJkBqLm7sk50XqKIPCmWJK
nOlJbyqoM5oglz53yQd5tm5RxxVX4P37TY97Y3OeKeHSSlvU7t4O9stDdGRfyxtmgAkK8aJjba7C
PRdXOlsQaBYLP9ocy8e6dtUoiPl1MR9FwcRAa4E5tOArnb8mqN9YSBrWxaQpsavribrhEU8hzCvU
7Wvxu32XEpgPqgCOTvJfhqrPRIS0P7nE/Gi1sBUnhfo3lXX+uqg/PbgiwicEP22lbXCE+F+MwX2J
gNUClq9JUA9bNmcOvGgJidn4n30oGTnuXyONoCk1ZObc72OwvvMCLOdPs47tZ/dZZRXFBtWYYMto
WFuKK9OF2rwv06d+5RCflf23NeBNG1uoGbbZGrb4rmjTg7z/oqevXc2YW08ducLSr45vese5/vuV
cn4s/xTbhAqlAqg4G4/xQRDab52WDkFn11jX6qvS2C1ZdXxqSPBYmaixctWrv/BlgCJ/j9qwzFAQ
CdcRy4ntlxNUs9EqFHS6M3THQ0rr4DB8D/kiZ0vSsQSTQ+P562uK6DxG5eMcGD7dAEAkMo54QtAR
KIKQmsoG4hQcK8T4c3LEtNBvfQ0zKrFsvbgKHAIlnnlI6341qL0K7LQcD83Y9PvNXNGKSA8+vEL3
BQfP8RYXiekaVY/Wg8oSCQ3OjQnLiCgRn0yQ2cx9GOPVqNpQqAvG9hl85WRndPJOC82FcGyLIfCj
RtYcgljcfxoE6beJRy/NKsUARcN/r6X6Dv6b4dHIr70/nXOMj7A15q5C+BHLQv5bZ61YXSNfewgl
bUP8obPGLMMZdYaOdzhXBtzHr/vR2MTqiUvZZK7ev6Vf9LVRvYpI3kOHm3U0SvOeUOqsxOSp1/tK
5+IQHuLm8BI+4rxuqlxQkjXjNpvS1xtQ3RGBR03TLDlIFSB/K3i9RW3ahGt8KrVWDQTJRhxNxrcA
H4hOP8zdLiA8aIrBx4ohGY1LhSV8dTLyWoRimG7zXFdBsPMsUsS7JwHJj7ymX7JT5FRjbShRlzKi
PjO1xXWSh6NMGI8GgjhSa9MH2o2rHhZfiVhT683puc8Ji7AGpynXgTDSmsO5RjuR3fXX8h8Zd46F
kIANVUxeqnHsjG1iY1wn13qdZmjzzPNmOsmL1KSqBDStSd/YuWa7kKtaxYW5zNWunbeUbKdLzJhY
X7/U7ph4o95T5kL8q8Qn2leIubxW3iG8XEni0BZ+X74Vg+j6LpZNbUun5XRdzH8XUlQzNXEwNuX4
SgaW8COOj4/nOOBD0THwkKKkphd7oHMfCb+MeX1V3KhQ8Zr3HwjRm61UWFFb6erC/5tYAW+o3swq
mQDadnF+VW6kXqIZPucAsPBIM9Womu9c/5kb+iqukYXt4Kz6nZvhvUaBsvPvHdggy2gwJfFaxam9
ii5RjtiZ6zEo4JC2REEBryA6xZJuNmIsTFTvtPuJ1K/n9h6MZ2EKoRz54NX8hKVEPDifwiH6ol2x
fCCa44w9GGH3RdFb98Vp1H8de85IQkUl8pRbhEwAdylnYyW5FuQY6VnIZFa31rYRgm8OG5Ili0zu
SijageR7Xd7J2SA3TrOlM6lQy0KzU4KCWxmc5ML8qHfNHiqIbXosKiVPypAR8z4OLHqRJ/G9F0/i
B5/fDCpckDcsJkrm0ESE9Jm4arlo36jyM97LH+0EPCquJWMnBXkO63D1T55kyTiwz8wuOMQVk0vo
QnRMdMzHzqyxOICT1/E3H3tGoLJb38WinDxTh8MZUGnmgIjoyffB0yveHbcrvuWoX8wsbrNT0HpZ
43RkwUkzcKqrr2YWgKmVv8BmcG+l3jGL4YwfjwCUv4SaNnTx3Y7UPiyzT9jdaQXVatfj48z/CXi6
ICaPo0hJszp+x87q1LP39eieUPxl/z7m4jUoJQFSrUehg7TbcYZikMKjrRXoDDP+rfl3CGz8x2F9
6kuZlSs0HtKh9Dt7EZXE59kPxPUP8k0MxU5czRbGVPET2nXAJrDnxKkRZY95iUzI6Xo7t9odbTiC
kBmdzLo2pRaJeegao32RRazOCIAR4fSwZ/J8sdeqD13KUEcDnABLIvnijwQYLsxnb8DvEwhd7JSQ
U5KPXHdCaYJ5mUScx5vn5n0oNwGNntgLU47hAbyBBm7VpmDu/PveieNWkNEQxqBiqk2dPguGjJ/f
FHVXcdSWMjCBHnkFWZZWQY3gzh2MxiJgZjRVu2kAYtnxJLVQSCXPteHtZg94nvTmHAPWmYVmEYfj
VBLF/P/77qqegj2nFMa96EDrqS3ojDMRapHwBKV2ZRyH/JT9O9+Qa9YVSPzzOwxBBOBJIfGetEw9
9Yac9fFm6pxKxgPwtGDSZhAc3CS/yiYYp3/37tj66z65GMi78Qn4Y3CgQBVXT2ji5NeVJySMNyso
xSTSyY2sikVTN+ppIJFruZwwPHTZAmjjFn1DLyLLCtogjg4p1LHvS2lM67qIpSrFYS/4vUQrWU3H
FWPW7Gs4RBg44M7aKVWQv1RMFxn3JQqQor11kAlO1RsX9h/skZHMg3LlqaXMbg8Susnbr72OWpuW
Zg8FO5YDYqadm5bTqLooy7BhGwrXfLUjIz9Ay41haRJGHsU4WNpGrcme3RSCjLaybcnYHpYH/tGD
QAzeQ617VacqzYzmi4XDc376JuxsaSsCuAYV4tFhvVehym64s6VGICaPeBqHU1qPyhoKW1d1qdZy
LdwWr4YL3Qea6FNQIVQ3K2GvPuQItwiM+fNuFb7ScEtCb3SXlIPsnNG9USMiOIQlLCfnj+hIy+uO
LRlLtm2tOyO8wQKztYsA9xDunLcO0693/LmBvnqVljzvjbXfctJBM5adyT0B/qon57/c0dN/wwYu
n0csB7WYXFO9RUvxXq6U3Hga91kQj5sfmJhqV8JW0ueP53WM9/BKOFKiQN9lgHHS6S3261SfN3zU
Z5vkyCA9UOfBNLrRB4fZKfjhieW9VkUcGYmucQTDEKfbYzqKHVJK0sOLGv5hPqfYzYIieeJpDXpp
gJdbSlIIasJOR/X/1MqTpylEcucaHGCNJFY18w+KWqXLmVkvDOAx7EdZ+Ckg69VDuKlV6UWO2XyH
GtxctjBsCH7POn2XEnSwxUM6rBnuBlTVZigu2lq44bByAvSeMUtj9+K1x4oKG0Prct7CBKeIOZlW
YUX/F14BJi8L/OBrmR6c/7BreUCMeia9M8Zc/MMCtAj0I+Zu7BtBh9GiyweBIVtwhtLpaTWkDNgm
lLTG6QFZjH+pNHDAdquBrp1u4FwXudYf05wKIXW45M9mc0ZVF69JMKIAfQGoMsnnoYooAnZsneqW
HhUPKx2+q8xWz0xvIG2+RVnxn5pPFxBpTSDDtsq7XArt1gkL8T3Xo0SxsnwI/s/J4KuWVnCEDgEp
u7OYo0/mkrwrCAJyhCVfWQoXT8ww9UqZOZfh8lWOPMiuUU2NZAyMoqi/DMHUw9VHZCRochIBoEQp
TRTAqun1eLMHcCH7Xr+ZmcTnHXtlmj+u/F63i1jkcEyFtKg7785UKQJqW1yHMTbHdk0gKbFVCLk2
HwNvyDAxJksIkW9NqdevfJzn1O3rXIs1ntsu1+q20sE5pZsZjtwjB5M1NPLAjBUKtUm3sn2dgXvZ
ZOCTiSlpvPaFMGnJzao4WUPiZ3B2CFcEptW6oAy4hnou6BFOrXj5uSl9vGoqf/tLPzyrJQykQIiv
qqwCvsIhi+3ofCmaHUVDLDGfeFKPk/hFvfE+j4p7GgB0shd3/bx7cb2tVM4TfYZhL4ALjfxtJXkj
3xKxugapQAboWomDLRnagQ8lMMAQEckqTMjNcx8FG+Jy0AmQxUJXBYURTXCHa1uaKkjLfvmuAvzg
jd3ndBX8s+VrGUbpBdIrrSa0QCFb8hi6k2wtFvLhg9SpO9+XbWQzK0k+DJjnHbMjCAduQJKEgeyO
46uR7a323cm+Wi6mVIRboSNgnToLjCozQ62eXydTGAuUAbWyG2HH0VTSsR2tQmFPTjdUjzImUg5B
35gI9ZFoVyxZvt6Ya0yYGyrDSw148on7t6QflGKqVhT1s5T/OmE1+hnybl5FtOaZHkCBeAleN211
vomiprWkaXB8Vu3TkUk4NgG5t8PLULGKa3//u2wL/Tafy/0sm5ez5DBLKi7QeX69rXnLeWIcsexd
hc7SefWzWW/Ar9OaY9wWiqk+Md0Of5LB9Un31ovUvv/ugr6b8kD63CWliUBJjYETTJ2kFTapQykx
SZ/Noh7aJpOXhKzvIWTzn6Bv23zC0hPc+012pD+b+NT4xOMXz8k/73PiVfaTDWf/xz98Xugo6eIz
76DLVwmuAkYRhG3TfiRt402QEeuEZqCsshG5LQZYQeV4iUMJCh7TXv4YK/YMId4s/sfRnu71+Gfl
fWbvdi/nYL23TbhIOlvHKKBktAvNUysdfmniXBoy6zDE+hXreg+kP9JFoW/hZMsF0sknsPf8rh8x
sLkRKNZJvPfxsf3vxxPAL9JX5H+1PX4bFBck4CI+TyMmEjEFQfJQPIjKy1Liky91PDUKWdoSr+An
/sWelB1FOAblFLNEaCNkc2BAFqnUv0tMro65rp17N9bJp5QGrwDBT9ehV0HZHsw41QEp7VNLhJL9
Zw4IvoggOsipP6Xpe23UbV0E6e/pAEODLdttcxqL4kNSS6+hjerQmePI7z1gvEMpl6DUzxs38EQX
oBawk1vPLo0mGpOLcpoIPDhI8OI+A+GX6+KRJcZamDOpoiVyqs69uy94HCcdxR9M4NVkLHHIPSVa
5zWN4VuNN4SnSzSRbMpZbmwUEqujOdpsMd7JqjMZhwVkeKtSGm+SQjc154JrSWjwlhE3o0yA9HLI
16OZYblIOoVEjonWsTDcSuHI1FvU5iUTO8ha5BTu9yiYBXwJix3Lh7LSETeW0EY+JmLk4h/I51Cd
GPGmbEvhcslFxCpnhxWw6L5FZaufIH6PNeC2SXKu4I6dGzZjge1f10ZRMe/iSaCzKMuWGypxYjZH
yKz/f+4Uhj7V78+oJchud31PmdL2ZLzs01WZ4yndfUX5gfeHcMS85g1MMbWFRu9fctQ1CXq94RUg
ummMRsPiL+6rqqje6hawHDZUGTRTMhKttjgIDnM0oAr+5OO2ehPwMzwa2y1iv80mHr4biC1PFMZ6
y6LlOrpQA2vHBBaXxS1RrxHaG5IZbH/oW7c7fM2yLwSsvy+h0AByhweXgaP2apWgIvwXfLw6cn2A
bgQ6n/3zW1Ywwd4E7/y2CEsqyukoKI1CF1BlbeZoCO0s8Xq4xDB8TMmFhSv8SnyzXUaUaK0lmjst
Y9Gk5wN6SZ932y4YcBtGDtdu8H/o/Kl/+CPs3S2dZc2Xrsh9bX3ctFskATr6HfTGcj0+GmGph683
tGfU3vy3S+wXpoSUQIhTphUcC4eBVfi6Ns4wjoEhzC0jFAkuFgFzu8a/GwmP26Q7ME3EDKS7Kcjl
Z/ZFxNNUzUoby0uX+jpSQpxYO/2S5IpzzipcTqcpditDX+cxZ/iUmsTLw6fgS+HRs9PWpuWGLb92
R1RJd8vQ8vYFkWLJeP1woCvdUQ4Zv6/u3Yu8UMvGWFBlVmqFxBexa+CADtm+uezyYRpb9ndZzAbr
+eJ8Ahag3VKrON+Rg7i5ENEfT+l34c03lUBqcDOSH4jF44bg69ftv/l5wIYDx210ZhjvjIb6LJ/U
DBm6MGvWNYbPdxoisGY8vtIS3ySvpJztjqdggflUoFZwg6Db+bLPkxHQhZXwF8GhOxRf35EfbbFK
yqptY24RXptEG71hbdVVPGVuspq/po0e+gI1LDD9fW9Q4PQ7cQCpQ6p41eays7s8zixNTQIYzD2J
pL1qqdPIeTvtOxKSKzbFzQcLyXGbEvBFbbyUToAxnA2OUDnq9dndiWWUa3kd8PRNhk67hZQJW1fv
MV7oa4IrXMVURAK8sbo0BodRLfBXkjV/CFzGyCD6Xtxk4tjueLMNYDmHRS+Ki4lYKwDYbULl+s8s
R0UGimSjTPbmkOLv8rV+1MtvxdVd/NJZQaNcQ5JvBMGfrwkglFxA2Wx93Z9Bw5hUWtx3bAizQUGv
Wy9j45gu81etpTneJNDE1AuywD8qyfmMMjRwOYyhoU2ngoUaWlB9bD7X0G0d+dfpJt+4+/mskxhd
IzXFR4lLIzZ5nfNfNpgeJ6seyUsWlPLwgwI/qt82IFuvpBCvcUdVAlAM770n85aWdkvNkHUIlIyi
+53xnzRctxYIE2veCwBI4Cea2xwjg0EwI4JeeQgpLUlOF0IazO5pWxfYrlANOvKadjOHhUgAlgDP
566MetcU2btBB2NLD6sspH1is9K7SJtE9LuN4oDkhl0w0wp1LFDAowzevEkcKzqSpNetyhXU/Pxl
XhqYkKjPiOQpGohkJj8l8enF0EJ44NdG4xw0qzWj/O4xNGBHTcWPpeVGqMpALzbnt/hqcqYUcXA9
zkRz2Ox+EM2xid46A++BxxQNHAWaHpPOGxIKJXq+f8BKLPEc42N+E+F8VRiKw+8EW3glKW6uZG8R
Dsdt7TiFkYgqsb2E8vhGlVBjFzVepWglEEazmGW2F+ZnMMuKOA8M0+hrVH9a/8ZircLQSadktyqN
+t8ReEF0ZL+gttqMPWcGg2FtAMTSELSJTo4iR9C2L0pzzpNRGNs06zAyj/DV3zrapr1L1myde6wT
wOKfmd1CG+CSk81NDIFllgFMYpGBiJOeX5S7CP7m5iX/SavaED/uljmjOhj8ZHa86jauMSPvrxUd
vU3YMytdHytULxdaePcrbHsHEG6Bm9pqX4q/aha9Z+oHWaQGskbgYBtKGp4y8kv+nT2pEw3KcuCl
RAoEeaDUZFd4wzrs610rWPStZE21v/CQ3TqwKjDIfBCATUh39dBjcP7rpAMRSxr4xXXZUiRpt75e
0RpCUTK8uXaPU5NMQvSHkXloVDXZxsMZNUbg+KVjclrNkq4qVnwtKReuBbpF7KYoHU4JY5C15YTa
znfFHzo9/PcndmPZYHfgdB8s0Dmv8q+8/Mdpvu9yCDB4GhaGxB/Cr563U2X8iXHDXozcJfEg43H9
vRCn/mlnGBjIxD69H8HTiTYPhCS7PVVXQ/zcIxVxVPiT8Jw2Mcx5Djg3gYQJirr/cw15UGOuywqd
g4MUkXHt/rKvm7uVdDND+gX5qRHimoxmEskyeu8HaZRXHKISlBa+a9O7YEnzaAXTJbemXpCc/Ty8
cDeQcDGM7KU1NXGb/RIE4xdZ4RiN6aj0quE8y1Ujju8i0Qgov7neEuFWdVwaCPv/xxaS4J/jumgw
JflELxbA1wsaWfPK8DkyiAAnGA7wIB4tkxI2u9ZWSOTFUEIgwnJGGJHDH4B/MGEBAXAFtId8cTsf
pkzZtbixPTD2CX9GchZ0UL2kQHXren1Ag+D5RmZe8JERG/+4zgeWboxxPUd3sie50kvh09RDNXk1
OvRyI04VVu4vp+L5AXOvM08MM6llTb0xCCqExAHVM6U/6eX9Uuy4itXJX4+uFu+ItlV9/KQHUs8J
aHZbT06SOxyEjqkGxUIhlkOWdYF1wOuTEwxW40lyky6t2FmdqvfMrdoCejN3QRFemnnFtPdE5CtJ
FePo/E9n3vMy1c8PFc9Vd8Y4Wc/YFEo87l3ypCNwOG09BpgfaM1NTNzcdZDSdIn6U9NmBF+RIEj7
bt/2XD2jChzUHMtgqP4NVE+wzQILcef2sS1k8acLBGcJlBx3acHuaHdPXIzBYat4deHjvjUKrfKA
aKao6KKELVR8ufaOpPQ/8kqfqxofFGJnBjqhmglYFTI8o20ZsV9odkf048pEoGXCpEULTR6zQBV7
jxuneuPhYpsP+UeWQ+Q6dVVaoF6aY0D+Ld+U4S1V0CYkWERV28886V002iyJ30I0fJ8RUndp4IJF
tJF4BMWhMSlIo9KE2eMqoK65wdoSXO1Qf87aE94C/m4y73AvzAQMIEz5L6nlBMC72HyvGYKi9TY8
6wDNNtQBJzW8RXTiXmyKF5hS0buMRZPv5WEABfl54uxOE7mjRxyl4nYYkAWKwScZ5RjbbIj+vu6e
L067xeKRHjgVZeA2bRshHpwCP4TZHLCMZ8khAeB/VcMHXieH+qR5TNHauvvsFH88nap+1XejOXtx
DTDCrQ2TID5Dd/7ssjKarOBYJqstSRZ9FV9zRHn41GdiClMxbyrBHhGK5kCxFXXPW/4Ba1H7zcUD
DrSV5LU6bDmS4CHf1WT5ZoAzfXgs7xf39x94JnfrZSYQy44IRNHotFn7q6pukQfYaVWAvDt5mTCW
HWZBe7bDg9UWXYVorxcIwRxNxCg/DRNo4wZEZnHITsEbz1x4DwqrsLEA3vllkPkYMI5wjtX+wWzA
BnOZ2lVqCc3OVRnvJ4vSSWbRrlbSr9lyYVeR+oWcC+KOmoa2Tvvvstl+YSgGJhJ3pr2GyJhz0JlI
McRa92cP1DvOAZWMlO6YY58X4WztA/dx7F51o2OTQSGh+RV95pVaquceEbBk5aKIrttQ2ems5OdG
YmBVO34v142jEGmRKQz4537szeyjnci4ghSzIM107OnV/EOXCaM1+EQwkNNXku4GbSjJ65XwYvPm
uHgoM+dIXDTQZo0mqsa5rU7TAwc9vZGvFwjQ7iqwFmNGe3zWnphs5Y5jFAZg58LxmSorISvRxVm6
vaJPacEDFriVSdXFe5yUn+Siom/BsGa+1iZiQqupmcoKzsjcFx2ZCz+r1pURmsPo8JJ/PuA6WNFS
ofNki/dRnDq9mw4VvR5b59NHfQWWHPraAEvIFQHnE1p6fzxrktESXA9hTnmkrHhacI1DdwVBBht8
DGKWZyQ+q+5qPlJeVGFPgu7RFO7sfuXapySlKAgNlylu7dFY7lSb00l3g/umJZTckEox/8ywFQV9
7bJ+GtjZrMc6wmugRjbP4t8B/Vi80xcKDUOaI3c07klTO9K7FLrQWLX0sU2XyOxO8rROagH7gH/s
BhY8D0r6cSQnxYMgYl8ST59x0HLWKg25KhRCOOwCOEGY4/D6c2vS74qF1pg7PKpd6jl2NW4fx0hh
2fNfkvFsCap3uthvv1F1EU6r0HZwoINq9zaeeNUBK3J6F1pElCnrBBxHFy7LBvdUZ8N/CizaKfWq
CCKdFuBW3YzvTtfPI+BdSMaMyngjOeEZWa8LIFbuWS54pKGlz9CMgU2lWTH3f/Ewvmm1WNu0GVRO
JhivTmYNc4VdqwMTsqaRUglZWnoh3vkG5PzctpFt4h0tqR1RVPVMlnPBTy5/dKsm5JnYhjiHSj6o
dA7zl+ti3kaGKIsVNQjgvOY8AiluoVE6w8wokm/rjEIyPm2nWB5vG1FYfOfgwaK2ds9zSbFEDnec
y8eI6Blq1iBw8gzlMl1DNAsIv8+adCWA9xqyrVMJ7FLcYOD+xI7+V+tJjwkPDavaW+E8eBC3mnn9
fkig35YdxvDUdx6oR9rg8CxEPyx9/ilU4uaXJNLXFumOXOv6/mTnRBqXfEnl0v70AKQoCff0flHZ
CJYp/ggvyj5S7f1FS4ks7RHKtrm+ZJWB4rnb2xTi82h1CtVAzzeg6NeypNYwcpNh0ddDIxs74f9j
HLXh5AEneH3L4JRTTviqP0Ot4ayykGMsVQdpsFG+O1tY/S9udmdzmpSfLLXUTBzRk9+WQl0B11I9
pL2YwruGURVNF3NnWLT8WFPL6qqYWNFA1jjeDmPI33eBmO0EYUi2SbtimoOVi+dhjPjJkShrdPkU
Iau2+kS/0OgvAquzyb7doVIT6SVvTQNu5I6EM2gTW55Shxv1EiouHH8l3nAtXruX7HGCnx7OguXl
Uq1Pi+jAKmuwe/cozS0DfK65AM0k0RnGRL5FNZ7bZ9I9GC2AORceJs+KT08arf3+BS7U5/H1SJkw
auEgSsLna02hjOQ53mDWGJHtQW23Ri3SMJTRLr8i42HFt2iXwrT5b02jAIx6MtoYEBYWHlrE1wBr
kXeHUWbCMXOm/xd3RKVJWYWnn+YVHWlFOz2u2Wwl4sp99mhOIe8na3mY+obMTqW2vSdGtVg+MaRC
hISwasasG7lLLLsbgYZ9VrpoRbzdlAevgBB8n7yqFbLleqvJBn1nwN5xS3B28zo1pDnVq4De3ezg
d0vPLBfJQkSU+2KjtDRbegFv4piJSjX99XF0O61kHo9XHU+35ybwcyJzju3IFTUmn3RFCDBHgV/C
KW3ftC5PITKEfSSv0k5EY87eVi24Se5oeUgF/B3y1O4PhEmykTNHlhPgPG9yzDXJ5E7uRuqoI8ii
UHw4XGSZnze6eMuyhpayFmhmu7eQma0II1euh7Cr7y7jkvNxj4F039xqN070Q0n/jKs+5PSizduh
KwPHOIBw0vp3dqu4G5E7af+KFG33TiZr7usYFj/OG5MUHHQsX4En0Ykpw5DBIoA5gk0vGIl9hpJe
D5KGbK+W5r+Gq/bZAywR070KD+/Zie8DpdM/EFKMCsZTmJeK/YpfmXZ4gvgi/IwH2Er5iGTm5GJM
Byg7DCDZsuvfLFIOiFvxD2lBkSsqYX6p/s75ebawlOyCKPir4UQLaBfTXUpkTQBqUNXh/IM7EuV1
yfKfoWTkIJUh6hJZDRuAtWhNMBPAo2hLTnP0X/OEsSjvXjVfMOoWYWUXXI/Lv6IJZlhKhtUEBcKa
0wP8UYpq2RC/lzVcYE1d9k2et72jkYOJjjh0bWBQSUOROjH6qFC3BjEHMEGnH0toVsPuaFKr2Tas
Sxf/MFgv97fkKS6nN413ebKmJEd0C0q+ZfrbAUa8LHSNXR3zhEn0gnKu1ziPg/oEXhdq7hnhXA8V
PF4V88ESvpLJYLyx/IeJlFdnV1vZfqi1Qz64zXdMVRvjUuWz1+nL6PU+tA420bhWSp5zokzZ4z49
X1FG5PYi5rVWqKiTx6WV69IeAM0l8LgcqSltDkcepBEElk22RU1BdYKGJHj/LjEOegCchCj6cBeh
5pmgGv6lRzd2DOgJuVBfJjzmNiqCfXLo6DJxek+p2nqltM1gFJ0odjcCu2zVZQ7akxW9QDWTkN3+
vRhzWyFwuSpmLckWneaHKpoY6XBuVNGm9A8/6BTceFwaWqkVIScJHJQxO3HwybhYgV6SydZSTsXo
5PIeMB0dhJPh3E3vITUm2zjZXElQPGmWhvbIEgTihd+uzUbwvXnPvM8UeE7DQt9hXI2Ow212hIxY
ew1a6GFppHMCKcl1EQ91CMIaGd91JvqM75DlHyFvm3jXbVAN54S97gNbNbfzrOGKKkJjnMyNMIoQ
zUU2yTojBMhBElYy0y0y4o7JjZfyXF6mJQI3GzifzLtrqcg3r6XKn8LgYgyy5I1uR1Ial9zUhqpT
xEMHP74HBZQOW6vgfCasNtvBJw7PBb/74b7HxtulvQF45zZzJm0ZIPox+sEApyTv59MT8dnVujEF
TJ3X4x8n2eZBsMze/5tp8mHEPcSeFodsoCfav7FovkC75m3GOPESHezMcSH2JwglkmeJxDzEkW5G
XcjnwBv+qRva+FUAu9lm9h0T/bKPL9zUjUgLGFd74YDl1i5h/Lg84EXf9bu3yTo47zpSmPUmBRBi
jhh2C2n38PK7slEyEZf8NRyXXbwQJWXNDffsTR1SQvP+AeHZzUNA5gDOdicbBf3z+QJt0c4joR8O
tKFiquFoU+0lyw4RWgXQZna5cClQ9I75tgn2Pq9Q8/VfTQkUgyN9Y0frgYMrzer16RLq70mbIk2s
cprqzF4un1+XlWdN3LZeZPGN2rB6i/xmW6r/DzhnfoETu1qJYZJqB5dGebDUyIlLFcPRF4mEfO8n
S34TXsQ+sRKC1ovquNW2yKNvO6kU40msLcsRje29h1LHC/S2LgzuBGfziL2hKs3DtannurZE4UA+
0YZ0cW1wzGVRLNsskAFlzyxN1VrjVQtTJ205CZY2+qY1I088s8Iqg3tDFcDvWGQ96uDLJTWmxPeA
afGVgo9k+tt80l5kd+mlImM23muVIPcPNPOjO9iNOQgwlJPTqgWawBhfK0pAQNrnpwu0A6Otiesz
nQTybMhw2APAjEDorhOCzzZt+REnXEhxCHq2U68Gr7hCHjGIey59kHUc1Biwe5If43gkOQBdM+mA
PtC2KPAZkUdhXA6j+3HELEoYXeEZCv9EI0BQQZ2uH/vOHa6wxGqmhIG5qX1lNpn/r7MdKmJz99fX
fYf7kA4DjkNU4abIe+puCR1YkrUY6/A+U0L+ka3w1zSygnKRTK5nuja/8FsGrP6wwaAoBdxFuZh/
Vx++5n+/mgYEjJhdiTIPLeQdff0GmNQFo3qPfgRNqrZgA+dCWUVAuumSRtKpnCvF3p4uwUuUCuQr
s5iI/XmP9yF58AYZys23n6+Gb4B+H2tngjn0Ur7Im4L2FvKL6wiKuQB37+NAH8TJ5ZpArwZKtfn5
zwW5YGMtcERbT/r2ODMiuzBQbvZOcNPXiwy+MqwZUzaiYUU6AzBS78IIeS6C12m/vw/oDRgS+Gwr
2eJ/4Neq6Zvat/Tn0SVDH62cxDypjrqTTAvH2v6AhCBcke4+1gWsWBQdtzDBp0FrU5zMhUUCziBc
owU296N3qajIAD7DXigqb51+DIF1ouPJ62CbgpP9PttQEFCoLzSkGVl7gr8gE0UaxeXkpsCSeZL6
jUUz1HKuPRxfmYBsI8PnZPlKxM9byyBJaLM9cIKg4xcJX0ktb4KfvtFHJHbEDoEp3EHhY3Tw7zaK
vvwEQrQQ+3hvThoTU1eYrcSfcYjrxUXK8x2jDNdJml5aNxEOP9/0iIhRFs1iSG28MJ3CGLm+caIw
hessw86wBwvaFM2W+O0Pii6okJ4ilbPif+K1fYAgYkKQxZjqdoXpGZSR12RlhRyw3PYBaFiVHuBK
T/5Q/pz/eaVUA/EnngIgQ0w6F6Wvc8ZukppTHLkbPIaYw/fm1uROKBcf7dgeHYyqfovp6SCqMvqf
k/+d41MN2UyLXTSKYSTdozLYAfOVLJRiRQt/oAlnHoAyEcZMlg9AGSRmPLSW2L1b5uWnj/9pTW5x
yvlQS8EFTzHy2TgumvkERZbBqmgl/zG4U2wMb518YmfyzzbYiaxIMvk0Rcd5UhxX0eTDSAuFd07Z
XzN8VTyvxXMxAUvtZR2M20JMIr5ktVQk2RtIq7ClUuj9MXeMEnt/rtvea9NJnhBQkKKc8QAxglkj
xyekKnGNQgRiAS44KN1LiIfmpsB63AMplI4XN6UkGR9cSbIwkuBnyiwuqdcGfK/K1mDNm7gzoo4j
jo7GNnCF020PhoCEBK/ZkFiOAqS8HBY5ln+KUcrzhT28W4QpshD4xhw6MP/O3UZKw5ja32+dcKBq
Crdo95+eJToI/jf3KKCPzjT+3+NmJvRSuqOLEDDgRe3fiUan398bH4JlGT47AOQbDSP68NcLUrov
zRHYNIQ3VT91xXuRwqi27Shx09G6fhmxkESgzNHIf/UtVnMzML0euXLPHfa8NM8rADkAIDs5HxB5
W6qeihUyjA3nMEJqJ+pFbEmmi1rUyf9KAFkgUSuwaw6Z2boGY37MYgEtgKHSAxefJXfhP5mDWmuO
0SA6X1kCZFbZwmMyaEZKCOZzWAgANVCG3I1Eiyyp+welevfQoee2wAurLm+3lAjTsPlEPTg7tCln
9ZVb5BVvE6GzV5/4lMwPml/mdFEZQDcYJC4YgswETACze93aT0cK0I8YIwXtbNQEWhlPRb4OGXFq
E12OavJwktnYLtLywlh3JWTtfbHtJwhVmECWkpBydbfs7D353DwUxRqFSiMcfWeNmKNaN13taRN4
Vom4hkMOmFna6Zugc9jpgniusDWJCbzf1k4m+IoyamVpcCyedmAiWB+HV+l4ngUXFl8QaQ88wGsw
p5xO9h62tEj0wfcEgcCGotBy48pYo008WOievTCheoDpGj/PwxqY7jbG04c7YUhS3GMN3atPOu07
HQWsMBR7ShATLamT/uBTkBl16YLdP1kY1jHrGc1GAQgn6UK2hq8ziv9n3uXMhIEhAwMvW2t0Mz96
QmEvufD84z3P/DgPV3lc/XXag93CvGOsIN2RVEvpZgD2aJGMoAV5VRyqEoiXS8UgpaeT1YC1X6zq
0WGr9axGwW4Em/L4nVQSWDPHelvM8sIVD41mXhv7MjM8n7JIx8ghEwLzFI23GzMhGa+cKjpZfslN
XIE0XYU6tEZj54XNlayzh+rJED3f3IETjU+EcXC8LcS96XVc/5KqKISl8MDd0J+GyjwS0/X1t9Tg
3r4M9jLh7wNO4APL8fiX9d3Tqu2+3/Eg9PTJj7jnhcn9lrFWaM5MRgaKYAO2LPGPnqhEhiFgUtof
KVJGSH1/dbvv3lQZTRNazqZBvE7oY8ThpCE88s6YSVEfQXYC/ZFuF9jby7ysEmdIracuwsNVP9o+
MrpjTKJ5zJyN+3zDZQuUoTJj4Ltsnv0fHIbaQz44PcsElPN+d3M390oqLVsj01d6MDB2j+/Z0/6h
ZyRiGDrSA4au9Cqt0EqFOw1dEmUyrjIdAti80n0i4tcmgVrN9oj2VpcT4OuJ0vAN8JIjvj4dfvtg
ZZfFBImaGloYaBBMNgLris6vW3cdAjlvSWwSzimef0ZsZQ8DpFpteJAezxgy73mY9lXlnUF1htaM
LkrYZKwhYiz4O4SqssQGzeK3CG5uRh/zHKB3UvRhNwjVSefTTRj4u/DXDhTRxmenbKVO43fUUFQr
embMRvZiLzrofy3oiAEfYN//48Q2J70n7Pt9OjqWVuCVfrjxy6OAkALwOiK+t2BjujBBesmC3Pt2
eDnzXGWfsEPVH/BooizRY3QdcPSlDctzchIPPovUMARkH/IAwIQ/VJlVVpMQjbarwnUMil++am2d
tnSfme3oPLJUBc0ZQDI+bWLIv3KFyCyDZGXRXLizS1MhHBwOuFjC21j/ykq40HetwoDMTlAtBuNY
TlqgdD9rDmvEvhz3LJuO0OlcLObDsZE5Bpx3T28n4BQ9bpezv1YoHzrzry2i/Enqki3ZqZjN9Dzw
ZDKowCQaVxlvwtUEAZuPD3wRTp/HWkXXBBGN7bohQDF+mGiUoWORt1/S3P7CxLyNDd2VFSorkpYa
LfCZVYYp2EBDrGU5YL95Ol77QK5w1geapcrDvEn7tt5JtZ+49JZ22wEYCo6XMxtph2zoGBd9xQsE
42TKb+XGzWJTxUB6SXSQcotWJCPekyuGxn3oM0mgBUPbojisB+EJoqnXV9uCQblQ6j37EMHr5cOu
FUKoJr/rDfidJWCB23mphY9/VrnfHg0fHfj+4DoGOdJECgX36ETvfJkppdVVeUh9uLGrA+zpgsG2
1dAydaWZnYzs/K9VFEeJQykdM13DsY1qdnbqpVME2NZIpFug5NxGkTlQkf1ao5OmEoEemPOAwl8G
XBRfS227y6xvVcAOROWDtDa3QGtwhldNpLkjukPIT8dcArbJsSq/4ecrOaHkF2vfppa7FpiCits8
k76CgWE+IgYg/kg41hkCnPTNInNq2DKZnQuPB6If2Z6kPfcx5Rin7R1HZAo6QmWbZITmtoGI6rUE
g81bZ7bIdnTQa/6ySLQT/fx/+EnMBxuN/1yh3TZ/1SXS6JtzGCSLkqebbbRx4pgZUv1m0GdZCi7/
N+RVk+U/yoZBacnatVC7TGb9BKah5u1VvVPsPLcjXfN+kOvYmaXhAz5wStaVJmXbaB6V7bVhCuxG
3ZZaMSVSqKzDLhSq0PALQmO9z+KoRQJYIkQrH8qmDd1oKST7CoZX5sbQCckbu0RlCSOfWLdQ34wO
kmrAqWJh/LJ5suzNTrdhHLqkJEsQV6Zrpym7uvlrHTy+dHEnTWdnhXKe5RCFKb4JLo7FksznYAo5
B9C4NzXWgUQCo9Bv6vdDhZ2tks++bXLenw6AJ8c5YNfswsOOemmqGwD6HAHKgmZihqTB7A5qhaNo
6t5fmuQ1WJWKXBQ3vU9OnZDHeQkgwaELMrBZhhobabA9u1f/0cj6Dei67fgdJ1TU5nUpDr4RNcKW
0+cj3WxVIk57QLX7LbC244L25bziwIyP3TI23DAaldt84yo+15LZ3dx7N2N7TJO4+fEAVHZM22yw
BxLWEFtW5zP8/KZDInmlU8MWXpotGa4nybN2krnChJdeux47x2wTHp+7KPHHtJ9rPe6YnJDTKUOY
KEwSvTWrpfFjxhFakZvwEbI+rgOUSIrLyVWY0Wd+Wnyosx+Je41bofO0R4kvkmpH2eW7yheBahi2
zRjn+uS0XRIaSuDRSwYitd7gs9r0E3aBJlIw/iayebaaTcl5WsPDyiFyMPzy7XZwOkg1ulDYDLSD
VI5W/eXPnjCaFk03YImBlyfgpDe81eimPs2VaKdaSKhrRH6n6eGZDoH51uK7vh5VDSALC0WR/M1R
T5Syi+1QtDsVRFb9Cf/+KZY+cyrTj4eZ3DYKeH/N8JkkFRL81Wjc4/R2a42ABzHI9XRkzynH3UN9
ofZ+7puoRiCN09dESFrCcD7zwbE/9GD/6qhs/5NHIhAzBVnGdp6yDkX5YD9FjrRpgLxxuy4r/M1v
ds5ytp2Qj9FeUJaWdgd5C3j0MBcengyXuYWF+NBZpOjFmIQleiy7PWuwV8ozOj+vmLMzWEm0/Llr
SUkcKYXSE5Fg/suwdobXM8aoXl71INo/wuJI+TaBEBgTfPstaQtqyR1jk07HCTxyp/wfEsQjAW0s
ZF9S/uHEzxekuCzrXHzbkqY5vBFMqgji/PS2v3UjGaNgcNdrtgiu+0YxvgL6roCcf/5qw+56YAkQ
sfLKIcPgdo0xoAy2u1AM4iB2Oc51Yaw/CC7mf+KCGGXdnGy2onHsJCkDsC/zcS3BVGvYVry7kH0G
kAXHsBHzsiw/JyezOnpScuQG9GKDEfTb1PKM4lIVt+gxlhOQLBQyhgOgMeA0myPT0KARsxTPJKFo
jwfpFmkxJtN0AVw6nfk4YQz9WGmZ8fcuXc+qT7T/6KhKeLsh/uVbv0k2qbGm0cM8sIpoRbgjNfvM
1rR1coEqfZoZ0MqVFVq8LwXMtrp8KpsqahCJUbMynm4v/M9lzpPAc1o+mJNEEKA24q4lZCelOMqU
T0fFR1afDG/6DB0b0i3ApLnlgVf3bD67PEIHylXKn4a11KP0d3Bz14Et7WSN/DFyij6/pONWcJ2d
NTzgTpB0uSejU12pOLAeil4T6DIP2OSRwp8ohYsLhK6ktRKSIPSoPoo2W++VxEeFUtlFHuLv6uok
cQORTYKb6FSFdEaIV1spl/p1eTVCOAu5mAS41xY00DcR/PvAi7NpFF3zMcLCZ/TH4gT2iDbFzJys
2qn+oJqe5RJYmVxFV1T8lffhIplSdObU02Kso37adUpNBn3CcaiFQV0LXMiT4xPH/Wg45LHeEPWF
JFyca26SvhB1Qm/8mftT5P40Xji7qS01cojz4vK6jr5cFJZTYSaDlOkFFE7Hsl+Pmgpxj9IzbeJV
j3T1OPw0xO+oFxklfAZXLTSsLf9PuME/St06kBxXiLTXElNH8m9CyOTr/SQLmXstbBvUARbu3Lxi
FIhAjial48yAuxnsVAHbqpSjL+ocVyvNJJvlLO04SbRFf4Is+rADQaaGJ+n6Lj1/750RJef1eLUz
PMv2iqXD3jrKZX7QYplvxLo0IS4sWT98VlOwHchqtYkfhNXbVZ5kGHlbbLPPcYolGX3s+qMQD9A6
JOPVI8e241mUvxJ6xTTvx+oE8XA7P47aKq5NK/5rO+WMG0qW9U8ks9amV0DsAnVtpBBeqYwIWEuK
QC+b1/fR/A4/TdTNAz/W97VUpALErv5/cM6E9S9rcmA6aJnLH0MqwuepqavjaUPZPDIa+ketWFjp
08KbTUJ0dU9ShY4gFrQn6JgpzUnSH1J0bIZgoLS4SMZtcc6qBk+61w50Ys7xvt33NE/o7FO7ADTD
w1EgxjI6bzyHXRbIsMbDLt4V/ru4MkygmYOkKLd3Wfn3EfeiK9i5/E+bG4OsCg1k8Og6+wzhgWV0
pUHnRu+DzDkHojxrZdPWLapmoDmEnC6Zo/6pacnQRJYr024GtzcAjhYNcEfiV6LkH8+/sAEkx1S6
uz/F2wI0g9xOAk+PVswjAiFfEz/g2fMjEgPWh15y5B12Af9DcgvyA5GiBIoquCkpIemeVAaCLkBV
Y6PRay4IL9t+w2YjdMD6txhjb0daLBsrRgsF/4sGDz4eGoP6TBM6+tOEulpu9Wza7OPVsx4w0X37
UmQifyiqheU4sTW8vQbt/m5Ug3WO/HNT+168x+o310abNJTFLYrw1gaSoyFKIiVlQeHWdkh2MDho
v86nMunSaADpemAzuXAiOdl3aF74h2JQwfDiHS3jzXS1KQHK+t4G7XvVHHXwku4NZd8o4eq1gSu4
tbuSDl712vjcNnGeSEBGR8nv+k/NOfm04x5Nnk7mQsYjhTgfL7ihNvdjm1LnuVch5dLI+V65OjBc
yrkKZqFxerz7Tisd/wnOfdDYIltZblNl9aBzGfcu2VVZHg3256bpcusfa54jQnghcg8yjovSwuA/
EL5nSKFb5tsmAOlm/J1eB1baIfK1FeoMWZWQoVGH4hSHaCzm2EMudY31oe1ba0T7Exy5j1dDYxmi
vCJx7dHRLlyLs72dXSdmwt5Okw73NT5UAySTS9Pk4cGPpPsqlWahRK2OHUYVy5WvKIEefZproqF9
XI8APU3g38gD2u6qR2r86ia057442RS8GdlfFPJ8pfDJwAx+Fd4LfNaXV5KwRtYPwfmWgmGWF7xt
M1jFL6JLpnrQpDLLFuv+e/+APncMKW/A6cd76pryfSS45zdDYHAUz1o7KuZPPNLbz9z/H7OjKO3o
YYtxkhiAjd+uumcqhxtG9SeZFayXp2ovZZNjxtv23/jdTouwvS5lMvq8i6jiT70Hj7f5HFUEE71W
4tqdw0BGGLgPKksICfolYlaps3wLPzkXG87CsKbL+KgpSe3KBVFC/OD3ivC+iV602jOsfj7C5Rij
VYc92vo2QLNvdS8HSCJFullAk6ixpxCu1dOy92xQOzHgoluqZPUCgVrpknGmPOv9NqJsc7igx7Oa
y2Md4YmbABGmxzvCS01BGKAqWW1ysoRjSZIdb7Z70IEY4FB8wW1SjuE49izqb2Jocg2xiU1FY1qa
cHZ4I7wrKhHrr1PjWGU0azG/FAgiO0472fp6DySympJGNfaIWpz/QNveYd0wUU/bzPs/ujh8Q23P
livpOWrl8+N/+FNIXON0EKRqVD25tSk2alz2G6+eMvVm5JnZlvv1N/5HlHUhVlr0dq90/zresFIB
MyzZ/K67PtQ8XKsx/9WZm4Wa1BgjNkQkgKCs1v9oaBpe4Yh6orBSHsnsaASYuaLbm8eazHmzm0bZ
xsXmlRFHJAx09dLngu+v7pFmERAOs/a1ATmx4kdhdY2K5BWljYN3GPVtenC+EvTo7dhe6D5C43k1
iq7LxzKNTWVQ87TpL80GQ5vPW6F5a3aNo3SzeN58ZGnnx+1cbtxnt9/U80zVsy7+XcHAej+DwToJ
uBsbvO2QuBQwCpR3tWD8VCEzFIciBBrYJINZHaT0oWn8Wm5upGyqc/UQfJ0Pn3mCtCGXLB+TLzC0
/cflFuKNZt9CZUocIki8a6i3MUeJBjR/sRb7lXLitYlwzdVewh3p+7ejycjvQ9t7V08U+MKbTcTk
HL9vsne4qIgDwShEl5P8y9RSSaqoNbbFIBnrFD0kpZc9u/24OOKhd3zvpLjP/Q8qc8z795nDv0MV
mc+BpXclgW5r6D88Q5lyFyAzmlfb2ddJEY/6AAdbXvA7l1zxCIPrPUXF/edTE57unEQ+DpL0L3bb
IxXHF/HbmjlRWv2KIw1K7lGHLMqumO+HeETuHWrI9/O825pAPGzUTbC1AXBKk+tcrGwsXKyMKGbV
EjziDma1/d2K78ATKT3n4alxAIQiBDjFcKRd+EZiK3Fp31Qjf72BwJNLMZ9Lq9081P+0MOr1xcbk
BWR3PFLaw8KAdz2Aj7dh6EOyPhu7lE2Sa1vg1GJw/ST5GppBSNCQCzxmiRMH5ftAHwQhZy9cbQ71
08HbI16eSRKhg57qmoTQjrSZOozUpzKvdzbW8JyDmxe6COjvZt87PoM67+trEhqq1toF8zDz8TTL
PQnEPUAB38fLTg63u3MLrshC/mnbzaaYd6yTtACuoGjhR1ImFoHL1C7EyvsM9eJgsUosqr/+PucT
1cZaZI1d8KUP0ZJPTzKvOcnUoGZDWCMEiYsTMAU0zBGY5yl+eUg1tCDsMKHq+6URXFsz/I5VIY13
DuIbDxpTaMI72bSn2xroKQmNZ/4ZfaKcpITtZG9lmQCqahIAFMogdFGr30+xKvwrOfB6CUo4AjVe
FVfV4kZOxHh6YoxtSjZ2Q12iNeTghD1hq2Pihy38PAtlYvVy/6gX5A1HPJTGRpnRXKpwiA5qYxSC
ifA/70Wx7c+Y5+qHA8mNTzl8Mhk/qSI5XC90pZ2QiBwhh0c8WQrGGPGrWOSicbNZ853LKTHYKp2m
B+I+prMmUNR/WZz7hZXIwmjVEtnQYCYQ3eTEksop94DprQCE8M1V+/KWIFyz8enwL6eCVX83zp1x
NCzz6/cbK/wXoMH+aBTZYS6uNgfyuHYOLxxq565joei9hbz+tRPyPwYSVUodsKN+doyL8NeRjYUX
AraigG3FEj507xnUwF8z2dlmiurwca5Qr/zic7pHhTsWO5Ozur/T6GgybgLfNqgx5Z5pPy9gGJDU
UEjx1ZhO+fNDx/rlqx6OD6T1yww7ARzsXsoM66eCsK7qJd3hlpsNM6lpO4jN+Rw6FbGfqjzfY1Ck
cKZZl1fWciF45clpvjOQGvjfl3sRiKbSc+3LZPBceDXcmhk1okggvYZPG17fb/AlKTaqPyUjcwIW
oyD8yPWq3/ydEp25tj8NJhGMBDMUDWt+zvNjE1kNvhEX6cbF4Qx6tJHNNQC4ltpXAZfHgFPCkNsD
Fi1o0F2QyVhzRrGvRQ+twJHHp3VwN3ng0C25DoxygkQlf8sivPQxPJ/iRIRGJC0g1WHaG9cBy3D0
A7QxSNqsPDQzaAA1Tv1m9rU/yVeJAAir9YJU4NGfLm9QErymCld5jQj11KtQqMYcRSkKPahakvpn
JvbLlW7aCIY9nucuyljv7FI3oOMxupXt+p/1Cwt7M3If18gvarXym78jibV7aki7p0D9/KYpdmCG
mm2NUF4WyXQGGfZMX5Np+kMxYhOFSWRpJBek5uFk+sYjwpB11iNxWTSLF6l147Eb0EdxKe7IbY+i
X57nYsDywio9sOa7eDJh63bWSgjO2GmqK0EsYmGSVPNklpZK5yZOD9XDUlLqTsAnFJFCxS3oEz9E
HrhX+nvAeK/a8qW9HsFgvYdW9RpVMQTE+lA2Q/jStWV3reAU9YAhbpa15NsKfXwDZDVEQsKqy0JA
bhRLFyJQUSFlkt17ib7e1ccf72nhRTQHyoQQr9h76nbz3Vo0xhEORpL5lLsG4aHUZWbnoFRfYcpB
f1ZBsK6Qtg6LR4xSCJZkxEQv2gcEcxP1K8GHCWJ2ilHBnQkHwgvuAOTmSUBYcXuqM5ecfoKsd3dZ
nb0CLFce9Vu62vjblf0gxl7431m8q6p6MbDDWF06yRQfQNhVHmmVmtVY2xHaooqvVN6eBtnmO3z8
qRxktXWc8359sz5GYoyeSB3NuLGACLdWFv7nPE/1HV2Ng6iaLK/2/+C2xI9Uqenlp/SEPqYTf6o5
NKitV+BSGF1a2x8rfRm5Ax6g6AsqDilMbf569UB7W8+TdB0DrCwBHkBzhFUH8+LNYxzLMa/OKVbr
3lYCpMPrWIGQWuzhs/iBGF75F61/LIqcVMqN25X1iMOWTS1Qc86lCI+/w2dMg5/wh7k7YAdSyMsx
e1gSoakEDlS5RO8PVTK7TXXzNrRcJ9Lb82A1oV8VKePivWyuBqVByjgPuLbXAXvoG+As5HO/NUsw
T/9hi3P6JrXL39HkuPwAwjewQuDmwCw/pL6f7uqfMYvLjwNKFAYZgUf+y0QRZc2mkLVVwRNyCGVi
HdGl0XQtlujQGDo2MIFZDI3omO5dswOegXn9qNxJwvi1qH5ZI4Na+eMH3JbtvljwYWFqmQS8te54
RSqH/3vK3yJYcg1HCRcosb5aUwLAPbrwooY4R0HE3Cr1piAWvKh8sGtB6oln7i61TqU6ZCElVIwC
HWlGvRVlVOJUZl/dGpsWcpasjH6nW2lu5tITB24a/CtwfKYYL2A1MAWjZtiwhE46BJWa5yOnJnEx
BJHAAGENSTJTqZC9o9RUsIZlzw8lxx2yf8vMyj/B0iz6lc73iGlgOavAQ8T4/oAn8vF1z6EsKaUg
V293DnXQ71veITp5QNurqQ0RIFpBl2YQ+bbYGv1qjwNi+oLhrvq/LVCKRdRojqStPbz1l4d/WZUE
l5mOI6Zi66Yp1BSzFfymOmjknsuLSN5MeQVmBiNfLqWdXFGXCKyusmYdJNJsL2LigyTmcddtUyNK
qXNSwz6zP31FebN9Ju1HxUFws/MoSV2nJejpm8+3svzjOX2nuiLhrPFLwYqOmTH1AVWFnPu4B1ZU
j+Dksy8/ifaC+a0cm0IRicyDhWntFy+NI+DN2TD72paQeNiBbmboiUYlfX6S3zZExGrefr7f8cuS
Cgcj4UBFaXle8uvARd4n/6cjv3MvzuygH0J12NdbJsEPiyQ1EVDLiGNXtC8xGsiJRqXO00FTg5lg
fa4Z8NIwKoDAKtT/pbDqXO0l6H68r7kizf0Y2tb6bNRSFz0HwL57+TbJu31Gl+Bm+rXpei2z6jEV
9Pd6FAR6zxyzV3rOPtnjNafGysA/UDI7UYjBMeQwGhXgJ+iZAF/+FhTEBXnJ/SSBUZt4miHhO4Oy
Uwjp50BganzdEyWAF9ByrBNL+ZaL0ZVDWxYVtdci/x+TamY35Es7+TNbrSG3kaTqK2nafvwmQizE
7tPlE+kHSpzdmvH5aQ3S8WBWjGEZ3pJcXfSwrHolofqO0Vx0MV5v7yBHqN6ieojQ7wdZpYk980Wh
sp+3rwCrPJgLrU6hIiU8CIKc85ZvniEB9v0LSnl1iJH9K7iD9H2dm52FQ/BH3r/45mfli9LXdwcP
VQkekHh0zp0yonnV08SY933ZoG0P8U4eu0CR2jtxxkDW49pQya4LW3s2Ht6IqX90hdNX8w0JqpXK
RU4yDqbSyjjXhGZskF9eagKIAWU5U3IMEdu15NXKAheL0cGG/AEGPqhe4argVCr9bD4Ic4pBUCXu
JoKhbnm6HcVqXudVXhfnKuSIJar8eoZz4uqo0f/HljF/fuhDIVfm15JFVPiBdhQW69dfNTYq6Ifb
F/EIviYJ9uoY5r++2Bx8NKW7vxwmvRnVj5poa9j2fQsw+35WyJx8dHBJxKpPU76Y5gAflqlwg5au
tlrKqTyHbAhpLxz49nXDJ4+wbltq+J/qEeOqw8MUOEQb90IaHTSDIJqzz+Jhlueqb5SNgwYL0Xn8
RZ5WG9G/67cLi7w0hw/x3OfsFlqr9KdiWz4pGG31kaxYnuj5MgNUxqnK0cGfDw0LOdVdLlPs0eev
v37c5YPuqV4DcnQRURtg101/U6dtXOFV8VEWT+owxXNVtSdHJr0hvkWGT1v21JEO5BdHAW/ow38n
e7Nk3JpGP1qGiz+YThF3x168N0kVOgtpvRRkbIxiaTNzpYit+oa/yEBId9f3y1Zs8bQRpK9H6Y6T
RtNk9N+xkt8/LIJ/JYii2r6mUh9r7PuiDR7lrMYvOxdXdOuTtbDwB4vL0A7P3/K1v3g0SBReErDo
k+ogrzvznX3ReyQ/HGG3YOgWget6GmjvTIbJWykgQjNY1agBj1a93HZODfEZvQ0GAzwVRCsT2VzR
t1iT2PfE4R7A07yjn2mnS+y8FumpFqdcdGQKmq84lOtOUY38orxicxJL1tFezP65t20T76ZxT7c1
fzoS0HcuZWlxSnb3FCm+T9itX7yOJqXfIL9wIbe5Q9688xnjwwRL/erpc+b69aHHMoIwqS4QYAX6
2zL7PGyZkFLj3HPUbJw7jmj7ln0pq/O4vFdSM8X3h977Yq59Ve/JahM2v1hdeUc8Ip01apyYl3r7
J1tgbCeRjroEM3p3zgkuI6FlxhmdWn2u+afwven09t/i4fHv0+p1235buAkVKftWlgLFoczoNEQa
m2gYt95cOXQwb8V4I7fIqJOjWXdqOIhn3tWBy8hMQt0s6+P2HWXnj1nAiWhSg8By7t+hAcDVX/E0
vjU+cr5pEu0UrVfHPjaRqBfyAgHOuLQ4KQ/mfMNu5tMAHNWr/HmkY0jZ9aAkqtBzuKznBC2wCG98
DUKMOHEIrkAcG/x3iAFst/VKTJFwzUzk2v7XeGv3Zu9I+Wvq2vxNdnZgHQ3d/bL9VLBUP8oqEsJK
HGLQtCP2BfUmnTp1oyTIE+Af8PAF6RgX8nxCFaTv8MI/y9hwwHjZXp64CABLbeSzIBvplxBxEX9X
/0fWLpktX2HHDpmyzjs04naxNzxgpOXcgVk5q+cEWwfpRgeMqGFIK6orDtepYWenzLvttOoTxUj3
+sXI7JSufdgvBI4q1cXRelWx0ELNIZ3xloRh8KXK98EiW3lbknEcgK+y1GXeQxJb+pelW/PnKYb4
9H8+p/ljf9IX8b5vtOdmRt5XBZaWo7drQwz38loE0xgPrmqhirJ3NEsFMzbz/vpdHQnccqxuNAbe
zEtf3UwIb2bKaNs8A4uIL+onCgD/nuHMWhygp5f0CcO2zA0H6yVcQjndPwzNujs5lKm/5neiIiwk
EKuIRqQfCuW68G9HuuNvL+VbqgqaXGgQtFq5JmYg5ocf6CEbB5BML6+3N+Uq2BcYTMKbW5pSNQEn
ztsLVr2DCNbYM9MjIUda/xZYxmZfBdi4VHJNgTnsiNUF6xszhm6M/R/Eq3apYgOv0t3H2M1mOruD
tp++mS5VVolG5Dzz5Ok+6NwuR21GiaruYbkjVK322W5ZWGqi61seAZPIQcE08g7cjH8ivj/HDbDj
degJWTO+LuNYmJYBjTcmVw0qScAR2DRt6YFZfsgL6pgLmnHthkn9OjDKAJaP9yY/b4CG7aZFRZvQ
hDafyZXAsIa2EjG7wdtqIfY4OUrnPUz9J/ecHvSqm23NcWGwum2jdSB0QePerjFJuvNYNQgjAzOQ
fXhvpS7mURq+iQavf6aK2c+G4PzX3Bw0pgf7bM8tFm7SPaFoyYyOPPDCQKjQxPTX0cioI/g3MpFi
XZZJYfFw3EHYDmosGTM0WMcaKfFGQkeuDYunP+WYsALGlu7HZa4cUwj/6hEpe2GyowduYJRHWMfC
m8w3gzxypmMZpMHpALW7IfKX6ZHzlC0LpUENp5zpYuJVkADNmOsd6LIxj4/Ne+angz7Y54gFS2Gx
5UgLsNZPTCWVZj6sKEypxVHF7yHaYXsuTcJHM1/gMbo62HdlVSgkeEisMDd3lFv1A0Z+Bqx8O1by
S5yMGmA8LfL857kLxUr8/1BsBeeQEiZbwoLIyx5fvsJ2d7Z9BzYoR7lDG86VcDHlLKQsD7/gkGVE
vCS0DoAYqqqqZaIR0kgBfWTy48hHD4V9Fwi01IHQSYoofn1sr9T7J3HXIAePzIJmPpay+SptDw2L
l1pXKbK2eljIpdkTf6w3gS/IhksP1KFTx43NypkGp+CEdTsvftYp/hsuc0kTzBqr58vKDg205Qeu
ZCAftdMDZ6t04/s5vlM+WltIJiOia/D0RLLhRezDYw+omycSH0xJw1Wf9B3JqAMq4gC3IuYVcIGr
gkg2SpdFDsdR4L/YTlk45veGXdl2Cr5teTL9JEwzJ8NV6h+eibzWlPJUSTf/0HQ9w4jIcY8fVGI3
Aujv8WNAH6Cnye14Trr3cN3rzdOTmrb1Qt9aF2fp0QpGUXSCcr4gscr5JazXYFK/ZpH7aLFSjBkL
gOVvW2+KzsaqMlOD2ikaHR3g5C/tuvMHNs2GUFakOr2KQeqWq9uVZhTOabf9jkq7kq/THoHn20BO
Zl4WSscM2cqvuQ9V0yeDYG2SYIQ6/+BSW0NyDKr9ypTo/IPCgg+pucL6OdEyZMynN8gw5BQO9Dhs
5ACKgc9c1WKzLJoaKk5GnucNI0vf3SB3QdYKKv/hHYrqarwl0nmsrzyPRU0QFGEBZqZL4TuHjWgt
WqGB1BsspwSJVfN+/IXLQ+u3Wg3yhmspcLq31anWD3mcPmYhlaldD0rSd99yP/ZOLepky4s654sK
ZhFBGnjSn6mwmNG3pl0c3ugzZlIQK4/xftp5BsJ8H9sGcPluQmeWHRibP+kThJ1pRWlmT3s4ch60
5C/OSvJpZRb/VcxntHYvK1ZvXkGoFn+9JqUp+rGJlOK7kMIdjt4PEIJDfCGKutnQMbM/yZm7lXV/
yEbLNe1Q9peqogXLjpMKujMmOW614HkVFN3AgYQ6UgUClwVJ0lfacc5RHcFnkrWjLnTofxdE7rSH
p7bzeUUjwZXy1w8tAQyGRXEjrvZx2Z1HY2PhGHfKQGHdymcg1pbD1eW9frgfo/d7HLyOSFz8a2lb
IaLKItHsnNBu4Yrwq46P1+R6kH/X/E0VGPfmZGe8I1DdZb6HmcI9Mu7+sXI2PByUzxyM6gOvF/6g
m0u7uDl5tSMIwcQvjTJKftNVX/IDj5szTFknV/E2Uf0x3sn205gf+CByzK1tlthrfvB5HBQwwR7T
qV/g4m0b4dCKUmOT+OqUGDLFlpJokABtVYy6DLFkaRYuu7mUgtPCC555zE4itF8QV058YuADR5ZA
4+4hrYj0LMse7HrmqaYpcD55xSexTD9Rw0zR18pL2/7K8KFNFwx4P6Wg/kK/HJBfcM+cem486qqN
rWMw2USyyb2l6ybuTEYo5HN8jByVBDmwMNv9xEBvO+L/wL9I8Gt9+E0OyRjYcGnPVb57F0uM09bq
KgYEUy2D7oWpLKDx5t1I8QFQzdhixlpeizHl2NOtGc+RZsnHOo01K/+DV6lCSk4dewiw8KQcLQyb
hIdXvCPgMbp+Tin8wsAKfj7WCoiu64gjz9EbrerleCrekyv8mZ8agnCYf8ts8Z21RDgM1UduPcnO
RzXbMQPnOIoKBI42BF32MwhbfA7cCWXv7ulm3JgUC+IzVGihMHaJ6D6ggbqE1Ow3/RywZR0P+4xl
/C4VHTnySfd9Wbztd8USlrSuNWbmxzcJ6a+AiVxBryZXRjwTR4/FTtP09DNxXn2303i+/jM0FdKK
ErQF+gc60QZ3b0pkUaa23hXRpDF4tzVlHvGVYgz1SN5aNg9bJXJ0KfyxUHuyoTo7pucOWhl0omyC
yMbI76eUzEb5EwOBqnrikeAlaWto0lKM99r1mWwq8wNPbENLXVgMHFEFCMMPBeRcYW0GYgJcgbDI
DW12/IWryYsVQC1CmYPFnn8OKr0cWKxJhOHOaCDhrZGNvFxB3sOTEj82pf6EivRQLCZlaCCiZrL3
SQKMblrpH0ZjXF8BkQe2jX6gOLAAOM73O8mbQhcfFJjrofv1AeHClwFxu7qfrghmrvidJneFq/va
jHQYTTy2va2iyECD19TwEuFwUcH88Nkq4qniBAkGJs1RRfA9Vwp+IL7xWX6JnKEi5IfotIOYTIYy
MmJAEtwd4p9I57O1SM6YV1ZSrf92eHVGoxQf4o4HV8O2JaeXSaVxbAbu/DXqqEFQxamfPQvGcQAo
kLAonAx8LqJGAjTUf5VAsxffv77sDq85PLokw121LVrgSaIPdj7iuzo6sGE3w8hbiJssKZL3w9rb
1FvOQqzzv3Zunk6TTs1OwY7F8cekZpelbytJaATehJ/W0IiHEVrl8sKNiUWcLAx6MTguGzxiorLS
Lq+iAYdQHtGto18c8uHo5SgajY+cc5/KIvCoSkf6aYP2fQyuMnHPbn0xsda0dr9d89s6hwHKhj/9
bb1ImDLBBzwVUrDjOPup4Sai6jjbwvVyeUjbCKChJ6bJZAkYEEs1jK3X6iuvu0Zb3F9IA/nnya77
cEgG/Fi5d4uENHOhKyTF+BxYwAOVWb5hddpN2bjPUrIMeEQalS8cxB3VlPYzNiT5bxawt+fYyLy8
2hiLABG87OS/Nno7ZOQEf/gzfGC80bk7KbJlvnGGqntp1Td4ZQOar48BKYHaV5U7A9Ddx5/3kZw3
iCSdeKYFWU78ezJM3ENisjhZvZk8cDF2IOVXqj4SwJ7oACF0T3QVxGFsUJZFp9HoH3l3O6ezUdOu
1qdnOjy5LZY9ZcBeldGhny/VhHDBgvyMur+NrPcMn/lJN6gH86tSXZkLXvW/M57QZ1YPXJdXDo5a
DZeEqu2v7pI0cYdQmTBEvl99c9LlwlVB5zN0McZvncQMdLeR1snDkwWanzAvwc2oB9enE+wYxSfQ
+or9NSKkyVETE6pjE8HgBsBLLv1plqaNHsCWRZDKovZlX0Izer1+qa7AEXpbraB4RjQkB9QxPD8w
5RQ5ebiLE2+5w6Phn1OiPiUiLGyqLeAJvYO2yb4y9VMd2EVY29NMv2OUuZWOJCfkHRcaKIJ35tFC
G4Foue4fBLJ3VQ1E348hGAP0i/+BzKkulo45FIhnTpeBSNsVISdcM5yrEJscQeaD4DNuKw26Bnsf
bEBt5GeHx4PO2LLClPjcXu1ole+ty+XYzrp2ZsV7Yzm+BvuO77o2t4rHDqPmoj7WhDzar9WEqlKb
BBZ7HygRJzvegLKetceN1sDgq9dNoeU2lZXc40V5MDLkQ1OrO7aT+wvvAHQVw0o5NWmlh9mfxiZS
5ZD4ACawMbhZC92y1w5VGtSiYqrxUmUCGTE/mi1k9MYSpTgLlPwvNDbcER8yyc3OK3JDslob+Jo2
Eb5n9g7k2fZnRYxG+cCsOQh9Oo3H4EkVNz1zJjYdTROCSiNKTbHw5MWO5RXn62LO8bEMyRIFeUPo
gxzvgO8do9GfQEiAZQlEw8xb5Ho6c3J4LuUQZ7xdkBVLpAnfmrDus7ujqrZ1J9ZeggbxKErqzTue
02M23qbtbV+OEn4V2hbZqlWZ6VjmY9nTzyvZN0XUJNJLCsmS3RPq6U8R4rWoV5/UbguGUxv/PvK1
yg70djK+WjUesh6BwqNbCa8QCA1qkTS8w3KibVx4ZOP9/gukRF/MjebJFNpHhFGIhTwbIEAgCTnM
AKahzsnjME/9L3jrQwZrlwT6d4t7T2x9oi0VFKNLdOp2GF2RZiY2jQ57LN1zJRJPhlcEDOi4y+tM
54IzTPAunMP3CKSAzLsOA53eErztXm89HL1ZowlSvpTpeP+a/3tLrddStkixSbg6rELDScsowQca
flNO0G+mzq/9hKZT9usTAyJjhSCMWGjeohU4eaDpDEsDVTVxgZZQ9rW7CWxJw9SoXo+27EnLNHTn
Ry5sJ4qgKYkjY/ZpQoYUb1bJHCSn/QTySl7BufdfhbBWYhoADmaXQiB0X1TXyNG6zT4alky9ouOI
RN2dzsFLMiChIscAtgta/MeQSLMsJAkCapeelU5zCz1vHyjdyu8mkOSi8fsMMEQ+PyGUVEBleky3
GUKBPpFKjpHCCdQPwkXA4mQFm2KYKlmu77mlBqun30HcBhnl1zdhWom8r9WJzFat7/ZBQVV1USCa
MQU4QqsmLCWeOrnplSwzVamDvVX1b7s9QYo/8+TH80+t8i3CFEhvStWLOIw1TYFKQd513KvfNbsK
cGXJrdeKyrePxEkRw4p91dFlaiRkYWkcdLhgmaOeStk0Af4YD1S20rd3lVWiRveDO676UzGK12/o
XySE82Lr2OlpIX0wT4px4+XYq4BVjnFshZXrzb196TqwRqJ+dM0uXVF7GEIqOztkn1858o/GuQIW
L3Dtcf4w2oKjh8W9843wePagIMuTwoNCZ7Fwpa2D404kkg2+MAodVagfv1T9J5y/w0aGz4YYbLQI
cRI2xDmIO3hcxDf/hLKE9LUjxGgdBibq4coPYy0NWa2lzJOxeSf+bRr2K1LYeaHgtJwsFdm/s1A3
GLzBZwK10U9MJTZGaFKYX5Vf+fcKzeQEMbxrZydhbHlTAChrMx3WoB396/9NCChFO98DV8YtgJz1
AYKuZxqx6DOwyC15N8uzgDGWxk67wjq/X39v2R2a8Ikq9+qKIFVyeyFUGJVqM7l0fLbPRyNmi6xg
Cztpy0MITwpIxERBrkkkkTjwhBTyzqjEq6nZw6EbJCsEIvwupdkxrxMBZ7r7Y91hq9YfXHVnwgYZ
ibOpaPQQtJ71UwrWbs45RbnyBQsiawqcNeUTMKBCfbTk7z6lAywGJ4PuaItMQWWwDC/0fcAfzssh
ydJjzyWfqJ/w9/n77ZAJz8SNpatYfuQDdQ1XrWT/Cjv+nUVXQFFmh01EdtUHMEexGpiNG/i4sEMJ
2aTt5IovXAAoZI/uTXu5QQUFInMqdN5fMwapyrNnDCaZmVRy6MiDa1VEFfoo7y86iE6hpU5tSHLY
t+KMiElyoRcGJf4/6E96j4aWl1FfaG0jitweA6iefeJBXL99FWrjw7L/6vZCpZOtFyzVf+aSlf8t
iWb6gxq5TF7BUAlDoygtjr32JNcX96e/xEq/qpRmJjT+JJJleytpo35rRznQNcrNj5oLk7FpLLuC
hTS5WYN96YlYYfcFFtbJKQCtSZqpmXbwYvycnaaY+zH4WSFMyJSUs6o/riORl8DdYBTMaJ8wcYDd
1g6P7NFS3wVjAjZCj001Gkoqr0TD+oQrD6Z3hOl8iW2HvLt5IEZ7NDNfNkuGjsY1y8TP/y/B/iAU
QmVq23CsaaSpk0BacGoWTA4awA9yArVNxlk+vcIEKguBSh25/b2J4hHj5NhsbRuQCASFR53D142V
3R2FAgyUWuNPBIwuz8E66AjYNk7wbM4CNoQ6NDJPKGdVT2aLJC6jCNNKBJbd6oOYnU/XwZ1JFvRx
gFQ6kDu6jEpRUWaL9H0wuuTm2C4xHAZAy3cRP1Fc3admZrSNFSixTiM1kH7Ue6bRG1HLNAF+JmkJ
JEw4h6xNIuxGWVw7odAgrrBk3OlGqP/q8qUb0SkpmYwIF50bawFH53/EqVR0079hPdb9kBj0TXs6
lYLa8e2ClPUltCHx3Ef4P+qT32bgXz/xyfo2dUSqsMjHqOWVx4SblkgPnMuKban+w6d4aqRw58r6
KQmTDCBV57DchmVmV+Xa+2wmGkFjlPJrMTNZHBnm74/xgD9OSXtc0/+hpXqXUkURzS1xVENqxw9B
cHkJ18qrIGg94chpa/u9BIyYFFs/q6vLyRHBfENw0OvLmoMMq2iLqtVNAXA7LarRKJCaZfH4TLAY
KH0LwBrpQQKj/uLy6UrfM3LWVsoMRPgBO33/6lVsjjBCA70iDNHiUgpkuiV56fdXTIvMMXOJeg/4
J3+N9e5FAXRtF3nxx+82B5UvkjzTpyJSH97OOspUgkSmYRSskocOw02E1MLz995rvjuuhCE5aeVD
t+OwrYd/tsR3254zipb/rEdZEDm+7mdWFXLrGo2lZxVNaM5H9v07DQEebWv5ZmqWDppzHTxnqDhH
z53gNthWjUhjYp143Vt43drelaHJozXTfwIj3pDkoP6n83H+0aFzEhEgkSYEhIAB4xQt9ux4LFkZ
CBwK2LkPKN3i1Vn/KDlko/nscZKGXld5p3WxEp/kciOm1CH6nHzNuQn50KTVWSUc4dc6/5oXZKAq
ZRPyyNQYy89ASwZPGKCvmeO4n+GfhhQ4jqMEEUWvbe1RcTfwrNMY1+VLO/JF7lj1M1/MEvYjQ8uO
7s3OWt4yMh374KTr/iXEz/s2e8qLtBSU5Ezf3gCdv75j7c5YcfgNOAykS50hq/ljrcEbdQuiDBg5
i3SAxNv4bicvDRqqyB9mqytHLrLP5u54MxCd2kDTpwpS45XqV15oZmR7k6ehaOtETDpptpxeCqor
jZuZ/sJgijcdSUhI1ZIVpfOiGAuyKFkv40SWgzplHm4fQQrYE1Djs9YzTxua6kIKXXSiDE3vEkiV
xV842wuOuWynPlvRejVaKgKxfOVTtElgIZbszZl0elTU16Yj89MRw6edF18OpQqfipRgPHwHV/w7
IX7FTSXSWJrqMneXNMgkjzqgk9B5n+BmBgW1ZmApBDWYaTeJVUmha8nE62AoWgBQAWULX+NUCXFL
6PPcPV7f5obWQcvKjK+ItFHBQT3mCBeoJ3FkPF91sxx+QVIIWwAN00bwkz+5t8P6NxlTbvms04jB
hurUnd3et7b0ZDFvwkWOfczsJVQ1xIL6SC5lEnY6VxNsImYgOg57M6I9usom1tF6f7ncM0wS4uYG
tVk+NYG4qH92XVa9nZ/IflTEWTyASm2DPp8Qw2EnRXc7AmpP4d7t/329FFLfLYvZcS8YfPIAIeNr
PKObdx4ZxHVxNTOTjCN0a8NFc/Ep9Fl/5Kdc8d2vkOs6pFR5Oq2YP3/BZRAS3X726whR8eRr3GqT
TtuVxcGGeXHzgQQ9Y2rvRQ9ZYjK1Ukzw4fKJkQvZvR/kjOwnF6QgL8mCHF4b8ALU+c7glp6GM0F7
hsEfne4MsK0Rkh5iCbd6tytoV+wRsl2+q8DAG7LL4HdP0kH7ZUvblKctSzGh50pUf0h/MWjA2D+K
l22gnl7J1+kOGndeyXJ50MzOMShHYt7FzJt1uFVb86besxRe4tBe2xYu129OLCJYtc6HtT7MffQA
3SC7hKTCN4q8d7ZbO1ccAnzIQEt3cql5Yazh7WW1BIqpUvbVRVlQAxadzrPyscvh/beLQqsayphI
qLNPhMhiEogRuzKy/kr1KGUxv1+nJ6ivqJpPZRBeJSRO5GdIDvHsWP+4Lq8P5W0sKUxjyOIDaAIT
aRURMhgQ9GGR46ow9YX4OgSnlXK0caW0rmYwkR80iGe4DizVVIGo5hS6OUmdEaYKvJl/LF4oytYP
eYTo1lrL8TSqmsociWdgTkYKuII575psz/LPLVAfp0eu2SFPrNwSiyLMyNXoPcWHGn/jypEi4WjD
hq3NH9d/NcPbHAP/vk1XZUBRU7D5n0kkQlMFvgPZU+wzGmVndb0qjg7jRRlVJpXnOKFfCHCVEqRb
xobKXzyAbJjRgXAYeHpF4RBZa07sDCKyZxo47psnDkRYbVIV+AGNwktrsFr7saYTnBKRwL+syw3y
Im56c3bf13wXoGb8U3jOmDnZVm2q0zxXUtwBBWLdnVNKQjh8U3CmXYROnai6hY0GaMq6iGiZBjtH
cuwHwFbEHCybC5BGynXs1iYw+hLzsZIx8VibRaJhWt88LjEuFV7OZbsCbq5qtRD41s8x5Tm37DBE
TQK5K30PfWbXZuFrwMGYQ6iiQ+E2hifroGtLawm8NUonul2sYpz1RePqAlUSUXaB4YzFquKFFOTx
E0vQ3B5MvsOMm2/Ur6ea/MHC0lCqQYNqV88OSEMLwUz2dDINqXkcKNAKgXhnwmaUEP0WhITJv++L
F24vh9l+dXsKmz2GhW7+zTDwI/Kyl+j+FD9KDfpLjS+vg/ej4qb7aipVKWGT7pQDMPdQkrpAt9c5
dgcHry0BjY/PMlN/+ek6R8upXHQ+2SprfR7B3dgzd9N/6y3Whl9LatP2Yh3u8LT9ziHFyAjA8M6v
ipwo+aLr3/zQCRcpwVrPjW77P4VnUsV9X4ae7y8krzxAyHSgFIy8kCe/sClPe/DubGJd8gzmFatj
PG6Y1Uo6wF70rOoBzsGYt7EXpsC0OBFrhn4VoPsqiUBF8kEH65tJ4YWG+w2ebGHoys4PNkOyX7oP
i1GD5TaUNzSZLHGxKDJae/C+Qeo4hIf8rV19ADojqgHz8Ng8EfzBRj/EhhmyzKo9QIYN3ZJE6dvm
LoWKOWhSE1txORJeMIgfIseFvr0aM6gKbsw3IsnykfhHxXebwuorWEFPGlvQUeGF4mb8EcZ5idLG
+7KaE+ivCQuUYviyR779gZ92i3q5kD8WcsclvXVC/F99xVjrx8xfTeZivNCozvvmmsPgRgarxIaU
ZnPSOPnr2HhxQNhScwuq5f+7VSTLtiHtpadqMrVdlsWWK4E0zILJ7i6hoLpjQ7IyARJBfwDWpNyw
vhoCW9PtEi0DimaGSPhJwaqZigHcbLrhGtxbKY6lsXQWxqvj9ce5H5Wdq6VKMXTWr2fDLlbZArI7
/+Wwbm56EN2vfgTrKa0WPwNeUr+T6rxhcAQpP3xhpTp/tc+n8ibKyWmSiASuy/8eZv3heg20m8Y9
cHGynzz95dB7RbiVE8zdaiU2z3zMYKEv803NUmC8KTcoJB3lFNm39r4kbljIfwUlS3k4PyL4GkZ/
+hamVzqoSwRwoJBh5cOgUYu3WDthGKIgbGNUhz5IycSAfu03M/OOSKzWDd19shSBedPu9b+bD9PG
PUebzRjuNmSorMdG0DfwCVMPEohjdLTg2XuNIMgWlvcMCAg+iEmzyHRn9upPhptDFSz+jPPN0vNX
/R1/NbqKhcVZwUPqBcyZuq8rQ+f7HXCiE2RpAKWcFMyHvlLAQcH6dYVNXQR/KZwTeqFUt8bhbvnP
ox3erdyFDdUp/9FOvJC/1aSdTtKp7jPCfsyZe3gdOyYH4kMONA5rRhoG/Tnde7Y5cyFb1eOd+0ZD
8NFsJTvbT5cBm43G6OAugEYGmUR8Nubtaa6gnl0rixd0PrDwYQt87vu30hagsOKA7feAvANPpJ9b
kusjU9ZicpU6FKoX7EOod4GgDd1GdKrdME+0PziWqus04Io2QCj8sSbvqsyk7cJlibLtI0hJIf4E
UTjii8qHKBCpxgfJHhLGAxu38A7nG2gkDNKuzHygzucQ7JE6dTwXBs2uZDxDtG8MwSMmQqGSh8Bb
21fsTv5ALkUOXq9EQu1aaJMsE9jxFWEkM3f5P6VVMDdIS1ZspJWpIXnCcCOjg7cINnrp9g44MFmo
I7Bwaqw+d9KJo2U4CLAZj1XmYnDDZ+S7dEeF+mUMGgEpXatpseO8toBu97O+dT0AWT27De6GzHZs
gouk3gjtH4CSduYrigwb5onncxYaXmq7PUU+LaAPxpRm/PUFCJIDJyu1HwRkmIdVoF7KZtiCKRvL
PonyWZoC2bpE7HfxcxZ2e/r9dtpg68O5wWA+4pYvQTd7Bga1BE+E9oeaSTUEV9hfDAsNwajpnrIn
T+gHvIGR+zMVkqEkJkHslOiDbSxUmtUTdhknAcTr+hXC4+V5st6L8InYC2ooUi6zkZlPTM9+C212
7iVON/yMbwv4oNDQJlLB771w0SkCgyF5pQQWbjK6SyDMJ9UepJ2H/fta/ivEAVpy0uRB2ysd+q9g
BhvvYU/oxYZZiYMGFf/zjIp1XVeB3RSL1PMhrIr3YmX++9vbGLJ93ZXo1GtDTEsUsTCKt7Nvwwfr
3jBYLD95V+0hADEum9vD3HgvrXN2f0xb3q95nQGkxYkdc0Yp5Oe49kAYb90g6v3QQwuntct+S8e/
vq0lV6sgGukCMn3+cHPI5/G4SSfsMr7hsJeIk2c1RSnjMDuFyKpR4/4YZJCKoVemnpxSgpyGfNW+
ToJ/nyLK+lbwlfIBQLZ1/uxNDn0jfrhDeQ2jUTMtcIOrP07Ndwbf2tg/QIxajUCiOOmAoxGDpz2r
9e4lyuyP6rsn+ijGv8xk+VaRzRGF75d50f5VaDvqd7SqEJW87juEuv/eFgUrhAKY6D/bpjpAirew
2rMICGDEUNHOqzOm+xhHgh1WC0ENe8oH76O/bumRffy8TeqecLvxVutiuotBbe5ZMmGdcYLwGkhb
d0vCtAeyd5kTaBTfi0aMYa6BktAA7GNk7FdVbcNmmJUdIuABmXptU/rCk3jjy+bxy/ZI+9V/t2wx
yUAp3WWqeankbTjbozqYZdNI2AWwV9XK5y0hAvJcCrPYCexHpfP3auwTbyQ1jBZaDIxsYJwJVRqF
LqWqcJ5moyrn5CHaDE3jp4iZnvNMDDKFoMExmCmUjUzdnVm0tf2LD7ifKMDz5Irf2+5expYWMpFl
YF2nXLU2kF1Z5k+ylZcU0VUsWd0aSuPrR1UxuqSmoznlicqvc+8g6vC+7aoNtsx5slj5lMY8/Nlc
OXtq0m+Yy2NvyZ5KcYzgPwx/9Dkw45KNgYy4ZCNM/m9+41VEiw2gx1RB9iv13DpZlF/RwogeuDVM
pKXooSNo+BaW6CD7iiwTSw7ENZ27B6z0dPRecnWbQDK/iBNZ8o3V70gAzN8qrJmmhqbVGtXSBPzA
DG1McxaGevWY22NGvERG38OEHv6jk3EHdmVe6sVpt9x8pvcpQnBKS2pzSOsTODg865XCn6uT4IZF
EI3icF1Tz/gikC3aMZ4zrCHzSW07ltkKVbyX3AjG4N7/OtiEtuEsRLjNcr5J6T+yXMv/0TxQYD1E
NPG2An3NQtEKqV0ExmxCkm80dC/g7I4DrqHJZ5i322++0hGTXmTdMesQfI9GiNU/Hs/T2vyAyHG9
UQVBr8wCWL/WjZurgrcrnxivckbL83AALLRABZQhGRaMFlDiQgUiIPpYVP+EMj1n0KMtsyRN9PoA
p22Qk3B7HC74v3ZRtPx4FcWgMDpDmT1v1BcDBT1upuqPqGJZUaFMiFTu9VxR1vypQSg6W4OgDZFA
18ILx6FfR+BwoV65NK8+6HeOhgIPSL8/gbRuMwi93FLUponO/Fj1EO9jN0gAljmeqye3Otb4pfxD
7QmoNB6nqrpXLABmA/jLIoRP/KiK+dAW23zWbUFt3ZcL9J1JUl3H7Ivhf2R4ZVX3m/pVVyLvhVJw
XW9ox9M1QMQHzCJMS4NEZbbb9qVXnO5waToVvijiwuydMiBuVzPj0llKoZsPPBWPQfZob3dwF9T3
O9Ezn94FxLuy/Ct9xJWnQpbRPN0YXfTOOu98GefbP5R4PlKR7o3fJkC3SyveEcTGG/+dqGUPH6g2
nqfAVhJnBpVs0sZF171ulYUfYb21icGgypYGBZb+kfi6fHMkT9pL5NXVLemQUjuRCQdPnzfr9QwD
TQ0V0ODVDP0ebasNsmnJib5voaOKAxKeFLZ6KTP5TAVNn0LYyjX7R4lY80qSAR39wDn2924EDn8i
wC0L4eCjVolzCh5TVnJsrUcc7ndaJM5rcdFznLYt/Q4WcWoinHf/D4+cRCQa8W62JdbiY4l0q2M4
9V1OX89WB4ujAr+pAoEkDLF37TgaJ+8BJ6/b9DcoYJKeTEjvcqQsNZpv9IKqAouYh/uzcI5bWw1A
+CG9gkYzAA5aEHFApMQKRFNp5BxdhQ72o2nThhY5PpywQOw8UAz/sY2sEUPwZSetimNYZahk+05h
V/QThosQyZapPb3UBKOhp82Y0BA1qiSGwxRTBssWJIO7h5dlCCS3wZw2SuOzbkr3TJaWUq9HZL3s
IwnUkfWNpRtNzJmL6V2xTZsH1tl/PTvuw7MjivG9w2JCyN9GXRhR4zfXwiv7BfqwyJCQu3h6Qa4R
Yqg6S52FYMmJZoBKLkrkcWimN6pyl+rDixItjcctdwa1b27I7M74ZVdzkD4bGqp7NSgNCKwdn6am
O6AWvQgcPEgBe5tHUl8n+PNGNj2n7jlnnReP0uBQpVG1w5rws773LuPBzDAn37HphnM1gWYuBcj4
RUYgPMqQpJamf3RGupIV7Nn3OfTbgDqiNpZLiiqOMiWpvL2KRYpipmx9v6tmck2MPeMK/3q08mox
J2AW7UheeGHU/F9fONZ/AWPgNvAgD2ieIjuZmNBaTYSNjHmP2NoHmfpAWn88pWgT1JLqEAGFALUc
X1FcsHESOcZ2urf3oImJQPuGar1OdIwMwbp+SBssTf55+gaIniJUHXjNHfCnNuHUKfOiKPpX69fb
WvV7+0tSvFriMudouClk5DPIAPtmm6NL4AuVFQ9xuC0Cw8tUNQy0GP2H2IOpsbvX/TMS506tN4Jg
IlzY+kF07n79UdXIHwIxnellc+uNKYUkh+YYiyZsLLlsnUmP4ko30kdAZooQ5xHRs95/E6Ud13t1
/BIfR/2rWCax9jKDPrp5H5HpIWYrJZo0eReOS058prIw+IJ8OKjNcNQdO+OADJ9YFC9QdSb/oZ/z
njBEsethN8G4iK3aunutMRBgi16YkBTYQ1AOOrn0QmABV6kd2UsWkQ9QGhiDzZVjETV+dSZwcFut
ouCHFlIT56qyaz1hl9adVw0pi1d/nYrobcq8tW6To/BSLBuheBFjxsLvc1LpEbDwJaZ+j/pqjfbq
kvCXyFB/o+1ZlqVP348g8V2rAkRSkZQoaom82JP7JxjL0d+cpKFW6spN6EFCE8BAFyrcpxUGPAT5
mN93I9tCP5z/QNSI7WPf889jjhW+6+myvH2g6gPiN4TEcGU5a3zr1h+xBK+JbUIhX+Hx+h1rteLQ
QsjpGGGf+0wCLfzOaUHnBsOWJFaZcpF+ggRCERmPdpDruDmc6PHHt4GPvUqOkO0RznkLmRmdnYEm
jaqlP9CUzMEYaSLvTCaFosJDWEefXOClowx7nO/9JKyY+Bz3Bb+Ioh410XVE08zYx1WF+KVArPfo
UNEjRCyLZkefKfJnAQsMZNCtECg24hpTWnqSMsQLooWeCrR30eAlI1Pm2HqNRcn2CJlc3ggJfLs5
ndyjKjJqKU2Y5KmJaiAaW8njhB/ykPr+uMMXlVgX7vsiSUUVzLsvUfJKBg3/3mejtDqvMZ3kng/C
Z+Pz0ap89dQfff/Tyvdw1lwHePfx2am4AR6Jkn/Q7fbTWti9t9hZqWkgEp8+N6d1blrD0MD7mv2E
BKnXlHzjutUcXQEXL1jjSRoAEw0T3AYI8kRW7z1/yOZ0n1WCZh+iYJhZcPA7ZqzGM2uKSt6olSPP
zj0hMtR9YdK6pUw1ONyT7mAqFRgOEIRJV0rU6BlgDY8lzvbf32zrCk1Fjh0WMt+2bfu8PWpXRJQ8
c+tfAhADVmTVtfKrJtwUi4PoxR6prnZ8iOnBUcnppa1OVEF2J5HI94OGB9QUihXPJu98eVsWhoVe
PPAPhfH76RO8dfA7DpMV+85UoeVcbydcmw8JZ+PJnZjjTbgvgswX8fq6JeMoVE/uY/IO+6Dl7jkU
wxYOMFE5xAFUA2NvSoN9iNbGsq9/7IYwbI6lmnW6Z5FGc8DjYjWid85Ihiv4vrcJbPdErm2O/iRI
7NhOMTlzh8lL7oNf9Ot8qSnBMS8le5eWcayZMG9nWDME7Ivq1vgur1sIiM5MLDf+TS5a3fSIm7fh
ydrJzzl+yR4PVI/OhXBd/6060PD5kTIDhcdwCpHXHXPRDg4w6U3Tpc1Vt1D5cNnVvyc21/sd48f3
xPLZ0wr3ivCipAShkhtrMZ5OjSYTAKeCdRydf871FTKW7soHF6muT2SPlOJZ1sGFjF9H6ZtAkbGY
/wnfj3KEvkjfvjcyf+43XzDx4244qmV1ElZUqPj7IZVyzbi0hJZVVMD7aN730rkAA4pu0UGsIoms
LUwJNE5Jb3+pxyI0O46JrmGpzekRHCPM/CL2u0+2cyLm6plKzVHmUgwR3pk6iKqMzsdIX+plKYLK
G/Q9gax64ZhMhSEZ127IBvoZjLz4ESim40c4mwdk+EL6PXhoojlPahE6NF39LdpzEPWdIetuFDat
BKL4/OIIWbD5p1B6qIxE8RtybOxGDuAy6h0APf7NGLQ2Zk/4Bc7F8KJNGMre2J3dSCqjZ8QPL3mg
mJG0RSmA9/BC4uRpcq6pRbLfs/fkx2QQprg4TiCXifjkWAXzDOvRhYtF5q8Qkc7EMzYJXVG8pe44
LIeKQkpRGLRjZx/yGi58TIkScu29XfpPHvpsUMOKdTPLxs9REeU3eyfLSaE1cYlqMdR+CxysBFNY
RdASmjJQI7rQDW/wx/oJzhS0sapEnSTAsA+Xlv+gLHu6BnKQrpD1f4N9jqs3pjVFbrk1L6BaRezr
BRHDsPq1j8W4y+y7f4uUfiB9YGojswLiw7/FprbMgitRtHwp8CoBjjsKK+BpmMAnjiWVfazrDI+q
41lilBG2JTSxOdeGYLBhM6qPccyKIPmq3RFBF39nU1nU15pSa9ZEUeeodclphA9V9YBp8BFFZ6YM
qDFfsXH1c4cKBFUbuVO6Ndm2D7ppWN3zeKWV3hLjFNa40YhhKDfizbkctrmqegGiAZeAJCm/8lmD
o27J7is+q74mF2mkTqnCf/ZHcMlpwDw8O/3li5yNkIog8A7tMmVsgV8guZ1Jazi2RHRAyhC7X+hS
oZBnx/s9yYitDeOV9QtFtQU4bNcJxKLMbAkUmktx99rf6JzSFLasKhEJXncBtIOkyHBlpw/0hHfm
mswd+quFSQjH98S6kDFK9dA6c3XWfg7GwJM0NIU2cJDZ3YW86/8PA7bjAo/KPw9S8IpZTpY5Om4+
PqnJZYe4xeoBCNjABMJXLnIXAbpOoBrwb07CG8T3ZLec3lzVpYG8gpSHp/hNxUCGw8R2HTvK3Z0Q
Tul5OKD4RSFMCeJbswIO7RDg7sFulC8mbDUXb/t6ElEHfKvPWnQ0pzevDm2EQ0Vox9CfFY/n1+lh
FuCVWqdSajLDD0hHnENVYMkbCOHBoA3ntjO9HiPMMOEcy/kUxhWm6r1kYdEM0TVTY/DXAQ4racEU
ij/Er98j41B+etUspGM4gJwn6xO2qa6DLp5bGN5+twh8zmph3bzwy3eFex7dBNy1p9o+Gcy51n85
wqp8Mgx/GTcisX1HLadiTCE5yOXHb4QK0w14TUi5OlmzV9Wq0Y8T2XvlMmtfJoyrSNQu2d4MWWbj
VCTudGzfXZRWLkD5xpBoIYGeJJOUJEsW8TpFJn0mk2Hz8i0iSPJzjVXIzHeabqLpeJDyvY20SdLa
/0jTdKwtH3zMYA1oybdfmfws3hFDz88VggGkBViUXKA4W9BzgubHEGEDJVKz2Nqh6GqGJ+Aj0YrQ
A3ojAZwTXl9FLjOeJ9EgV/p2BMTWkX+iuKBx68M1RvwxvuLt7eNpxRxi+Z0waTBldnzXWBjafz8a
DFsXQ0x01FRJtU5/cBfXfA2F4vkydh3u5E42GAo6H5fL6BcCHojdIiHh+xXBFuLcj6dlAEpfkeIt
oFwvoijyvMhCJ3TYjQNqWc8NLRFirl7/j9yMFnjcWi4jqgweoogZFYg25I9A0zJQ5z5LRnkhFv/C
pS0OzUIB2Dd0Is6J3qqG/VDt0sPYBic4UdoNgP5QP4hZLb0u8oQTCz52RbnfBkUARHyYUBbMHdf5
1iq7fQFCEwEsfH5yRYQ+2aaZnwOosZ8lkbEbYzzZ3Tza14xfx+peDqJgZl5KCVBGSw6UwaXy2U5/
7gu7MpJvcK8b26HZC/qEyFtTQ5DOPal07sYOe9WIJQCzklWmeyvPGpkKPeoUrNppscKisU1NNnAv
YHJAS07j1JK4d8U13MvtFiqggOv7Rqea2D6lD46A1aoDcXuA/JZToN71hOGtfzpRRfOJoiOUH0+N
CEUPM4SyJcdTjevafmymD8Dg3rEYZTe33untDWJGTkoKKyvWekeXWDX/X1WNtqkojkoTMrt4RrDU
WhMTJkNWtIYx6VAmydzW/Fvy2SppKjyv4LfJNEWq/fsr3+ix/IfiJ+0nxanArWRGvkjkjZeiD7dT
u/I9xl/VYozrzka3AuylEfeGLxV4x715wYY9EvYHoQjW7nOXs43EAajRReqET/X4Q/ywxYTRa8h1
/v0Z4x1KWpHg7HxevmZs3XSPSkFjEv6DOxVLqTX3KhsRNRzUSIroC9GudeQSvso0uoplNtQ+sCfQ
Q0MzK2Qdg0xtx/QEVIhlv1wbRrZp/EHqyb7QQ2DPzG1NHJGyBWR0tfv+RHF54VwzquVJT4cH06lM
0WsbnT735rr7m+ax/J2qZRKtrlXXh5cNWHJ12K8NQLc60XJG/O/qw71wYKiutd/g1/ctobxngciE
Gn3vUmMI7eSENjRTnf1+r2LLw2G3S6CpZGILgemt/QvbNrbXHf7+KMT0DPp6593LRbn7qYXg8/hw
txerq5ZdHCXeCpTeqdPsCLVqVba/VQj5/+TMIy+DwW4fB/JXwG7PX5vXSnkhmznWIaPXUiD67jP5
TEaF4TljImrCeCxN0/czFkJ2xVuODjV3/lIxM+Ph7+nyZeg1UWtLRMpDAEVrALhlRPu42KX6Pcxz
KfrIMuXNa5mda68mahxRE0HQJufRZVMnsIGByPbqIfdNCN0EhyjXc1yt/K3ieYQun60CYosE2vXd
emQZj3SFKYYygt+Qpg22tsu+3oYsTDjr/J2NigaY82BYiFwPycoJgVRI5wau9lGsQA9nikC+4fG/
s+WNHRlQmjJiFXcPDJGpDbCk7q2PpQDS5+grNhHoPjBtxUd3XGuOzWHN16OsTI+UYG7P0IccZWD7
IefXMqX+M/k+zHzQcwhHp208f9FS5/uWc/6L5blK9EtP4+JtiSYgouSwRGJ5lMd8NztnWk1NVMu4
rPgDFRDPpJyEV7rct8/FPWUD3FYRTfULxoP0WINAbJlqoIDof1OzxzNsUXFSe+xGytjQz55zQYAi
A8Zy4xbUkdsxOm8pAW40yjo0dgF0M1YKR0L4BPeCilBAeGkkLpOMR1p80sCJ83mWw8/0hOCE/dbj
tUcSO6SdbV55+iDBfmydMCxjLV+e0KPSujqhp18GNN6MwFhnCUqraLOju2S0fYHfnAf2Eho8R7ny
BIFdA3ogx5rs69w54QhFbyoFY4Jtp6Uf7wmcCSPUukVQRz5DWAearbds53//95h54EUHG/afT9Bi
WrddnVAHWDOHACxlXV57RAHy2eXtMYp29gK8UHXXsdKs821UCrZf9ARSB+WM594ipBZJ8z0iW/hK
GvAGWhZAhEAI4E8lF8n43uwrKy52Xdo6IWR33sTaurZuGhxuPQuy8p+t35U1Rh/cPpZnBv7/wPKt
bgiXFiRFDjhWN0CdjrFWZWfTUkZi0W5lEWs88kMlFq7m8v82AN63R/I3DVwLkJp00f9Bw6URodyK
Iqk1MeOMq7uN7nswAXRDdlxZUmasqG4giRsA/rWL2YgggdHUg1wHVQ7S+m2IHyPy3600uU3V06bz
5g9WYR5xhUMyU9LiRtMtX6B8bDRodIBtuOw3Y25WnxssUsPjpPqWiRmslrRIxHhOXfjPh/2b+Ylj
3bCGkvTTTQRWgFpFz1katZKkcbAVFfMiuGiMF2GfIzT4c8QQD7awXbsR6cuGZpDss35fjXQH+Ai8
p4O54nyDH7b9Im0GpxDwUoiqPFS56SIpL33EK7vvfrBEpWjPsmOlhYUe8xBj6bP9eSfwIUekER9R
jjwEE5gWYH/GkMmfvsqHwq11Rwxds4VRswkab5pdF4YIzcBiWvFfxP+CNBfU2oX6aw16TwtS/fTZ
tm1NZBv3wwoqiP7qptpgOr9CXHhQ5d7r+CsPRAYEX10BnRM3KOrLMX7pQNkOXkJ1LoARw5PsB/OT
0cZwxBXpSnYIGwLcHyUtl9cMMw7ur+p2daRxrBjF5DFaJfmED6QbNkbX80gUlicKi/eSDLTEGY73
WMPKCoNUGzGjFFQniU5hxmboGOK/cTsRqH6YwmKl7kZ8LbGXccElTVzOZ13M4PkELeq/yT4kntXS
g1Kr9MUoXNpBz0mItS4XBzZxibXvmvvKXaSroOFsnAF2aXcBUH282T2PgqnSr1X+f0QPBsiUMxGQ
2oE420eBgdOe9je53y+l+6+Y3DMt0eMRcJmhd9W81khPQNlYmTwlYofn6IZnVsyre6QNb5ZEiXjj
lJ0BryBty5JVsmjRUX90bQcNh0VLi3Sru37z/RKydM2J52SCjL2a6Zg6rPl/R9OxTeG5fr3eXak0
1q3pdgFdC4A4dUalVpwovyVvaXHUTfMWC4kGeNhiI0ayvVmJeAytQVigpIBTpKMxLgfyLIFvbls9
V/kSeqr2LB0ytOi0CW+kMBr7XkrBczUjz8DsARBEGPvAi7165wH2aC3DCsrx6zYm6q+61aPYg15z
EMtB3BO4HEbRtO7IFNl9XI80YIpZRaxtIiAclNDWNlIEnhX/HS265KeRZt55t6uyoMtFq9Pz0usu
SXeqRXBD5BASPHCtakeGeiX2cS1m2a4pWjVYIC9xzeItP8zUah07FnTDqEjbS9EI+GT+hlXfRuoN
1vzu26gXp7otUmX0VfptZyxQ2OxTFVWQTZ//jA50g8T8VYWMII2TbSZ7nzQReFgLTUFWojOSJTeY
/ut8PQpGUuawI3X2hEcQ8geGr4HXtqIfc/sL7uFE5mRC0yPMaJWeSoauKEDGBrE/altrW+JbJL52
zA2XzuAYzxJIOv7JwCtu6ohQevOE0cWZdKvyJ4LAL0pT5VS/4vEf7al2hZZNXqoXFKLmZowNigzg
klzTzOLfbNOc77ooKlzVP5HuKhjG9WoaNwV0S0kbk9C8EI/oto4PVDLehmKasMkftzPMfPBur2Aj
KmjcQ2VFCrYU527068IfvWpqugSdlSZzmt4QvbmfAFJtX7RMRpZzVk3ynyrTRiSG+xGXWKiZjQGY
cu3GueJUJrnWEhqcB8Cpusj8Y47tFetbEL34Vfw9SChFIz6WXFznuOAk6WzKpxwkDSJjQPWCAawY
Tm3q4TjdG7VmTv1XezA1IZxk/PJnDHoMRQ7jr4m/sJFudCj+w/BF/NmO4UAIFR3zh1jdvPeOCBkA
VahoO7kHG5SnOWYwwazMPvQRjPDjaFxxHYFUd51FThbaqLr6R8MZnkn7WdHB41C83v6co/YzZAli
/8ZIVnGDYk3gGipQwF0rpeayP6RDfaGDcndJrngdK4FJkiiwNh6LHV5/3AHlY7XRODcufJV79Zze
oibgHArXCPy7i5Ioj2RCyRBuDxpOmcOyAOdnJZMtNbL7H+WVB2pAOUOXOqqCvM9TQ419CFPXapuA
DjPS+rU6Upx0F+0tvWC+iWp3TALmMyeRPKYVIKLZ+U+znO3sOP+gzlhfi0MqwC15H7voctIP9nha
Z5LVUdt3Pd0pND5MwCBMgqKjrqmn3YjDBu6WA2rHZ2NgiUSZwhQfej1L9JzCKiTpHPffzHShzNCP
sXCLRTNRPwUJEG1KYA5daQDPLV88I5X10hQ54zudPCUpt+TuffaKsLY1aZK8CwcDdqpQxioSF61I
I5XWEUAjerwrgyExs8ys4HLRewXJopAj3crgMo8o0WBCeCQiuL6kF3Oau0D+3mycERMANtQLuBnJ
REQjSmM7X2DZ48+rRs0nvAUJUiC3InoOZ9Sje5x7QLe75dFbSz7036mCQjZfx4uUaA96ph7+XeIG
ya9zerqRqiV1JkQkRc6Jfk2JURnW4EyHU+0K7pvfkPxJufZvyVSOwRPGN0AfxOcerL02NCLcafLi
bozf43nNSFOkNOtOJhNsWNeuOrfzN7JpcdHE+HOLXWgR+eAs/JjlMRcwMyqBMN51KZrvldlXiMSw
bupAZ/lECVvjAYRgjOog74e1+wKiLbwM68D8BZajGfsrM9zWPbqjtkHdhZoOzsJUIKQ1ZBmHNRQH
hb6tK2Qng7SlNEYJsQTaao6oIetD5oX5yB57i+7qLWI90BEd1TFwOlrF9PDyhZ4kBNIXblAOdPvC
X01E9FlT8ZOzxpPfkIXOSq7fsToJQbNRtBV+/ttuQsbrPthpyrClw9n9bInGqaAUr/p62fLBaqkH
70Xpa+c3q2U0cNgI0NA4zp1XTsPPuLOd8k8VDEHtD6Fu7kT3GJSUwbnzP8Yo02veJaqaQD4rkwJ8
Q6CCG16EFHcif2ZLa/hcc1g9Gz5qKsr5qQP+R2q48+2Aok0gnsfK4Lcs4+4Y1bwjyxkw2QIKghVA
+0dd3mw+42WNoYN8Nc3cfFPW+UT9p95foWVEdZ8bl4SBxgeD9MxvfZZeXqA0AVT79zBDeyS1ybVy
4bIgUNqV892nDQ/H/AOvfsizmLIsPjfbp2l8z/VG/va9L4dzg/goP9TiffvJR5/J6xGk5DDTKa1A
/ycmWrGqUUZ9pB/xWDDtVssKvHg0eyes/JVvogzFIfSxNqCdY+CCQt61bXkJ1xmIfNMOJ6uYWmEs
VjXYeqSwq8OTa2zjiMmAoDgAWf+oqzCciVIsUR8smoy+DfZKGpDRWv2XJgkWXp4cTM17lWFhRA+h
YprujHTHSr1OjkjLEWvI05cjx9JflGVo/oLoLKCuhG2qQHqFD/ANXy5JYVdpRXI6aE8RGQKGHr+l
lL1/QR8BaUHX7IuV1H03etM7Lvj/RN/7WE4DCz397Q5BIifm2jzEblYTrakZajL3zVN6AKwJCneL
Tf3h4xwcLCEP+/vR/bZ2J0bH7EO/42+Hkte7P5SFMTw+uNmzeEGbdn+/S7yUUczBNTnbHvRB5jQY
v36jjdEpqVmOz8cQKecWcX8sGrz3jJqCZet19bxisWp5BaNXhxvg+lR63CwzxCClvmEnGIAKkO0B
uW7aS7pcj/hBcMi6DsWu2Osvyo4hV9FBgkiQSrzkJVmSMg3cxZXTG4vGxbrbE7iNEfhjYEEojcwR
KGH1goAiqU4xMfnVANc1oIHt1Y7eUx3eYuUm7heBbyzPq/YrwMHyPZhA/O4J+WgRMHrkRIZ0ExFg
MeYcJ2MfEKqxfe7g1F/i4j5mKVvdqwOSimTTUpwk4dkKcGPkO8N2q39kfoR0eZBjhKVQ0/Qt3QOM
g24R7v1RtQjtYRo0IBDxNk+rh+rIuTcKks8z/q0mx0+dFjyaT26LVSbyX6i+48f+X8E4m4YVPKzY
rqpH49lKJer3avrGa9BNGMc5GhO5U+o3sHkC/Xm4hSLQGORY/7vno4kH3BfNN2qoXZOKkV4O2kxS
19tJXjvLuBqhKXSm8qwKE0b015PJzBTRomMzbq/nqZBNlNPUfKrolKumI5353oPR+vRHZUleJ0QX
7+CXkoha7al9ZQ2/YSS/hWNHB8W5ne3ooq2NrKtc4RLMoFOdbE2oI1lZT0iP6/FHZqCoN+tuo1mf
1QsTW+D9FGWM31NaL8Wk3STjM4P7ij3izSYH2mgqUrmbei72EBOx9w078YXGfn70psVDDtSzHJ3u
T5IEhBUUwywvQSe6x6dw9GzxV2bz2Y3zrUn479L7OHR6OOa00pre5hdmt97uJ2XSQowb/N5sEYe4
/dzcKAGocmUwqWohkAR9i9/CtDklx8SaN/Tmq+25H4pvDat7gx8fIaSN5MlcLkNhkL9oXLx0LoNk
6o+aKNjMoIWu3misjV690DnLPqFlqs5KIwtmymG35/rnznj9MZTVwQgIZu+cSXYi/yrwpsFEKLX+
cpGojfop86o9Zs5kUVdhF4LqI1RCz6Aq9YWDWeFp65Eq0fxA7IB/9bMVYb8+A7PgbzW8rDgN/XYz
1j+lKuWF3Tx6ZrmQm9OsK7afKn1QutSvdNgysCSLrS9Y6etET+JONPUJscg66c1y7Qk03EWr4Zht
e+dCdav8AmwUQq8hbQQ9ZPmpFZprobGrYLfIJN8y4fLvvqDUdkyY+9GXWQpKlwLP0y9oPYTdqBQ6
jcn2Cx2trI9bT72/cr8kPMQS3mWBvYID4rcxbM3k25fMQQs9rbZnI8QRo4lDcfeKyuMy9awkf6sx
DYXSnkmXCf3LFkzV8fGagaZdUwlK3Ta+fSKRhS1I9oxmo0plZWlV8KL2erq0/9K+kBoNf3qfDD1a
1tUzpdQJ5lJ2KQpCNwpWeEKbYeTpAg9pz/5+RmGXACJsEY18lqru34Nsh7NhsRgYshhP5l/7rs3v
lSk2fptPYj/DTQBZSdw7PP57D7aCh/opPZ5nxIma8lO7CFc1I3/pD1WilaGjS9JmkdnVOFTDsYKO
cxb9CPkv1o2G1b9W59r02wArbBK3RYSaFaNUO/qM71nnnjA1tr8T7iBkM2FzcyrwjC1NPeI3eKqI
aWKTP9Xmi+ePlQMB4nWqB59jnVAVj36iGumxPmdiVyQkXF1P2ROsHF/ZzqTqfYDNxUrwhr84Eu8K
rfnnRrE5eVhpPD3CqZtMlhHaS8FEOxtGDLLhxySUJtxeWPbjbr6JGgAWMoRDObQYl0/3zmHMNyGb
ohRZEwNNOgX8an2odLDAyviqhvrCIqUvPugxySBiTRupl75G25X4qaYjE7auwsBgnMwoQbcXdMZu
XtL1yuCortvn0Wb4GRc4hiR0/uqREcdSPAaCwCUfym9nIiNlwtQ8XOlFmM9DEwyP/LnWlIUx6vQ1
4PKHjDpOsh9fzjaBTC5gDKJ9XNM6iaxRyANkT+r87rYhPRMCz2lObNqVggsYZ8IiZpjFYW1jrknP
m/Wk05mhjAOPgZVnohNlWw75fWp7vsMmH7f9AYl0SfvndAqE7WcShsuIiDLrkv0tbYex20URxxmF
rEUTqGSKV1eicazmmDjBs83aO0zSb4wFEA9cR5+/KlaZelDXTgVqquFDgCAGkFvUnFnXzkYujzKM
K7hwsJhv/032JUBgTXtI8MVk/uqVc+LkaAVmMaTsueUqV7NC/trkfp83c05elSydgqP0eGUdnDew
6pnH1RC9vFJvEHWpPgYRAMqd5gGLmN2RRHqbaZEN+eOg70QpnQO70BZxlt1elsOsk16HTHYgvmNz
Cs/3Ro+3+LjrM7omAiLb7EdXGqbiIeW4qK6hkD6klAIK7+7FIS91smpreoB4swf4/s05V1N7dxWb
fDlt0fFMjHwOTJCmRxvikYRgHTQgmdJanf26CiIi68eMiU+qM/3ZBCxVPBr0NAEDTeSmsZ1i7Ts0
jSxmm/z/JRvCk06mAdPpcwtaIcJhcmIQbnF805QvNr7MScAuHXfWjrC6QEscWfMpO8rQlqRqU1MP
0CeO+Ck8MjhRtHcIFMC6YlETN/zM84a409d8mMx58DkiwtqDC+4tptjTv3+SXwhwGfKuOTkLBVOE
VxROKth/16wD+t805O3MbyL8/dakTXZ1k3kZ9hJ1KdnMLGqz2V5VYCzZYLdP//+D9DXCpjf1H8k2
xQ2tq/19fLVbBs1eaMhtq8A/qD0+k07aj5xuZuernF1gFo3+ZCx/EDQ5AzjLWIRMsBnwY+A6jeo/
9IQfcRxT7DXvKsOzjrb5adEPl64TAihqyFQi+tIH+x3EfdzGeXGFd31htZR7IhE8KyhVH7t/TQhP
BwS7sMtu2DDd9775rob8QNDOP2LUo7CYJGwycJ5ZSb7p0LyD8OmpCxMNYugHel5UdJ/plNtfm2yq
4K6Bey6Nj/1BTj/0SkEb0Wi0NB5H65oMxMb57/tM4ofD6UGjD643zgPRVPZ1udWx9b2yHgW/qKRj
Q9zVCJV+VLLN/nOD9ME9YyPZxf/XRAzWue89aTb/TcvM0yQfT+rurSGvIE8x9PVM6yShDqIsRmD8
Dw1sARDEgM4Ogj8475lFRlHGPUM70AM2yi/xnM7M1+EXnsIVl+QgnQBkHSUufwM799QokOUzuMT2
aWjemThfoHYGHoMheMIq+c94cp0LKScwkVDhbOza1U+LUi8oWC/J4RAWJBi8f13szMq94rSiDP1B
YMRYCMLHTJHx2pm0SVOM6gUrD3aOEtVtRWzpkuRsclUMJS53CIoUZHLbDNJhrmK/jobQm+NDRDr5
1FsjxmBnQT7gO8nv5U2gVgmQLCRJiGFYl11SWqYPgRPj9Txi9czVydYqNnZ33n1MvJM8hGeWx+DY
e+yyCn4OFoA9Hsu2uiQHO8RuulMe7JFBy0FfwD7RQrw/QlT6W9qGLXVmkX0dmFgj0uTJuoXCyPGr
bvu5KwytJFskBmsJk4fLwv0Vxj8q3eSH9Si9p7MzHoDzzy18z/PiyzNUJA2yujUKcM0GgNJyLE10
GH5FeaVoaq3C4eudvKuDPBflNHdK6VI/sUh3DaiLm2gDvickkICkicbE26syB1Y16N1vArS/0th4
uhzbZjktqoc7pnpnIqWYIBWOW0xnysad6O8StgPtAv7sfQ6E8YdyMGD+meKfPb+YOVetiOTcVIFV
bH86rmp0qrUzEUlNiqBnv2O2/eH2FLo7F8/BN5SUYbGKX86r5GHmcc+c/MvQvZb5vqupYgopbOWj
v1JoSY+OFvsjNKg0R0KqVeFOpogl1aXT+MakPR+SPxMPugpbVO65TAA2PPgOoklXjHfHCzTfh7Yp
UUPcY3prxA0v8leMn0npXI2sXo/RBvjm+EdJu0W8ave3PhM8s8xZMns2pUexPQ5nr7wv3azxoUx0
m0IC6npXpVS6UmhWXFkGXXn63DLDjTSTphH1layEoBYcwwOSHhSew87v7KYtRxE8Igg2uWZsT6Vs
OehI3lMZmIFgch67n7V28LXfA3UNd53TcyRCUWoshHVhU3IenhIcoXKXmCcOUkJOp8ig9rV5weuH
fCCZt/7V7WX9AtLErHWKKQX4Yc2KMtQ5VhZv4es6HxjS+9QeJh6IfydA3gLnyndQzoSoOI+Fazsg
+1l2fBn18iCKdLfKbsWALg/wo6LeKyfY3vFeJSQTrjQ3eRxgNKEp+/+ZCIPXL4nmy7caAam/BFW2
r/7PVpIEyCGgYGMI4BIyFwBenvxCAiad65RzrrpcqHpjnmXOuvKjV9F/2BdTDskXDj2YeR8HM73b
1sTa6fz+SJimqcUdwRaLI7TANsGZHogKVDGN4ywT7Roitxwp7vV99so6raHfEmA9mwSCwy4jXCq4
pVuuopvnZpgMxdcbxqGCpbjHunhHzERp8b/NwCYlKFBDpOdbRFJO2qKBKXzJU7/tK8jMnjD6AuuK
Bq3ZRx0MLIuNCIeBFgnFdJewaiWycRwbKSwQ5SD1kn2FR4Ov2bzP8oAQdaiX/149YtKr/7BBGntj
vO/VEWuv2u6+/Sk0rpDCCc6hYSzq/fF+6YdRak9sL/FVSwU3AQpCoBxV3GxQwZg14EMq1vcuZiO+
4ybGQanz6Qfqk91Ic5Fh01rv2kynBCqINpQkz+oA/jkVmyL/1Vo8YJTpZPJCK4lE3NZWIhD7naO+
RE5t+stIZvfph615jHUaP/sHh0ncYgQj4ctA7YoPGnjBdu3JHN3mq0tNbKedlEoOu1kAHM7CphxD
RmNDg5ZHhpo/Xay3F99sXl5BHlgtsmj+ddQmcEyRi5BxS9YPZhIIswOFQgdV4ce+NUp0fLyYn0Ks
YJC0Xn+Um9Z8vc22iX4dZ3uw4f+4WdWiMvdgBAnzHCB3mUoaysTXL89dca7WjO2oQwh8b4rfdywo
XbVXypaRbzLF5gNKlIujFIo5OKrcK04reYvplrloIx1dAp3bb8v7jywFrxcl4lde3K2rHXMbtL+L
k4+8zNLvGnEJDNPRpQfXAHmKqLIONQjSHCc621HLT+TYsSs1Usu5fDp8n+B3mZvzS3pzaiCjfNvY
v2AE9znSAmOTBRbQYiS6W2+39YJol43JITPT53X0oj8c6OliuJKh1uvB8G1Jh5hDQd4vPoSpkzse
0OCnkBX5zSYxljX27s9naOV8wM3wgZjoSnzTFRBafZ4I85mA7muo7NmsK/M8DU6cAY8/cOWeoCh9
lTUK7noSk3rDhP1+LJx8YMmqNRUy2sk+/kgxiYJgXv0SCxLiBqiN0u6iotO40tUvfWS/DWW/JI5B
45V47dTqe0QyS2ViF7/rCETNJeHjU0tToRXcSp9sOxmlNF2uBC6Qbkfo5HgH5U4tlQeMjUF0nl6+
bALbb+qSsuawzQjv6mtJn9SKutxdtYlt0XVB5wCP3LdzhrHwx2KxsKkhWOAEynbANlJnGZSAsQ4Y
Iw0s7qvLzqHAhf1gAADt1Hml8EBsERfKXas27TpotzJfL+IKnbLCdGRd/9l8H4StTrBxw0mWAFyr
XoKIVAhjurrYc9T7Ci7q0jKKoFw9PnhsAKE235n1lY5SDSk2cL//x8dopPj4eLvzaIOIE0yadzZi
iHPA3rg5BVLR8DiHqWmrPJdWd0KGfTAzxV9wTQFEdhjRwuC6hrO0MMwVjxMkjFelHHVKcwfjc1/b
Gk3NkCPFTMJKsv/jikJ4mOIMveBQF9w9iUissmF6x7A9/P+vrTkl8BZb1169SFtp9RzqUos5P8YD
0uckG8vD7eZtgVFS20CXvdeM+YDNKFybMabl6xp5GyKiy98zktWJVganYL8w3NiRbNT+guRd92iG
lu+RZTg0pYYOsAHsmQx/B8V6WWRw2XDPir71sMOHVCNfjKpfCy01KH7Da+Qjo3Pt0udUnoNvWNpI
INyfPugM+sUsO69FzHr3KdkLd3AuatQTE+7rlJ9UB/3TJknFk1OE3pssjd051wi/vwtIaUIe52u5
qd3ystViYpd7jQNaVCBTIMCTWTStwGU+KUB+k2wh5hFEwelC0ArgmagNmQbmy3cHBtXt5yg0MMbf
wjRkeyHiOykzytSZmK/F149nojc/Pqke8ZGsahhIkqJ93AKHYFtEI6g1zk2BlnmKua71BysQHo8M
reBQZF2I0sF4QAUAzLJceyXoCv8ZJ7TNnjMtKTAf/ZHR7gNSucRus/jIY+hT0xKku7Hnha8jBVTt
HFFAAbfOqf1134tI7/3ClbXh6y2HWQ5EKRVcqFJdfGQ5FBjA9vqmwCh1xNWImno0X8Mvr2HT1APB
uuakPEmVz0buQwAQTCXdnsGyQAHH8AojEpT36UmHR7jxKrwSOGwMsU44b9/QdXr+N1z1ADz/wQE2
mA2M+athdhxrz0IypCPkSBdyIcIlH2xUrSPWvbGnI2zkmm9RsP19eTPvdB3PY9hsiP1upJH/F/QV
WAfjYH5TKPvjK1/lM6CAXaVb5Cs+O5M28L+Ck1UaLLdG8iAXyiTOPB0pOfLpCypsTdGF+ac5wTbS
U1nEnwavJyU3UTalpGiAlYs1qMhSYOR1A895AsfzqgphkM3wIM9qCqls/eiPDWBmQB2hpZOT/yBR
IsCpNJ1193K6CwX1JUDZOmUz2CX35o7ZmlS/pAii+nJoYcvj/FqaDqawWZE67Ar5M8abS93hniLx
MpMWCwUGFXT6AGe5AHG9urTqQ1aNc/0BFMeAxhAFlLOp2grL4nQM69Si+GiCnx5k2nrxzfGBZJ+B
eZPkHpeeQ+tRtSItGcmVubt6fJLwusOMLXZvBWIDlnz6vB+kmtPMRcLE6X6m+yUzvNhTnGreX9g0
k2Y54ph3vl6PUtppHWOR/OCisxfz67oWM7dfl3/Heu5fc8eELjwaffkQeKpptUYi+5KwahYLgC2J
YOVokBeD5DRRp3SBWGVifCINKYz46OL+ey16eBtjQMzcJ5lKKnsx8CXe/XL2i8y3E5o82YTO/u5D
24UBp3GTiJ2hXzQtAWrTA7FIITtZLlYEXvCwcEr66KkuBFLceOOLiWq8lfq84BGiqkWAjD+MhY52
LpDhamKBvPEg8g85/ku0fjKS5pMiY6trGcjdQFDQYICVGPKR9jGSTcPAqmC295mzcZeAMeSYI8DY
OPnL0WZ7ZfeWmqMuJa0QY1WJx0EDMfcfC0weBzTapDrl2ZI32BK4KPc3ZuLq7Sfy+lGfhoLYUdA9
kvtwSKxkfzGvfIrAF8T20ueigHi9T+x51mhWkHf3zV3O7zR2kNvS67Tj2cwEwP0TkQzKa/JLSFxq
WbQA98rSp9XUW0IeGcs3CPLaZe/gcYXYe94V1Z+eCOE29Tij6wQaunE//DSe73OrfXK4zEMHnfYp
Xoih/bDFYfv/zvzN+cy6VTHMtoHB209dp1S16ZHEY1SzPckSEbji7jBphPf3FBvzMq6hETDG5gzr
YHlEO6oolbA+N6hwA047WO0i0TbYGtZWOj/THBMjDsIHO50M1/+79q1lCK86ry5kCMvjft6Nfryj
u1trbtFkp4Az1tr7dWzovNDWWS2C6rVCexwMCMIONNlGqdND7wij0LLrDno9O4zpzcYbx4bnIeb8
YxQLl8/Mi1OePA4j78i5z49LkLJ37wLMXCnpCcyQtBlM9SNSnqEYqmDSRu/wcWKkHrD1FWiSgFx8
UhdKN1gZDQBJjnqnhFsgFS1jlpvEX9fWXl/hGyWLXmfSjC5o4onXxndJEd3hV+EuMURuzPaXdUUk
V+lSqBuPDurKN9rRnGxjPJCAE3JqvcFjnL+xwy0ptKGf0W2iFOJ9PbGzy/7iI4FAcU1fNdV74CJj
Ft9ezCw9ZJ/3YIH6Ma5V1Z65Hy1fVud3PPBnWpvK8s8mYY8Qcwz+QdvJCcWK9WtmqFoaZ7Wuxy48
F0XVK+IWjqJG2vyI8jjCbj5SOcWRNqz+AbZ6agYJXkTJJjQ9gMKbUCaKbpd2T64jNhy8uJz0Jz+e
FKcuHlPQtCqrttT391Cu3TfJb0qSgyBl/CJb4xozJCyp1yK3YOz9Jowv3MaLS7E/EdovSXcyPSw6
+me2Rmytj1X57DpIOyDBS6IVSt2F4DdjexMXJhbDrjP7Ou1Yh1iFOM4GWBBfxXNM4E50ncRtpzTg
+wK5/mJFzkNVKFBto83BO2e8UhJSIxL3dZ6MMJfYQ5D6w2fg8XpfgqK6llaaJ87qBMYghVBqUvF3
Nk2OmdGuXwR4GUQsPKDDUqTkXlzKoltl8Q+vMhwDnBm8RND2nx8VdcVug/pKfxJ/vynYvGHpFBGC
KDyyZmwJNa0taP/HlPdQ9uS1xMktdbD4hiUVW6W0M0BoTJLrDo0F47ADeWWu8adT8axzLeEu4uHn
BueVPXdvVAiVIHk7Ca9V8IxitGsPeAyjSdcXULn3cwXJCvZ4N7ItOQJx2DGFEqYPGIz+CCeQ9MjV
voZTAFTjMAJkUufztimrMZ5DwVFSZPVsU8O2fF51qWZKko0UGNpuOWsRqyYtPndeN6iyFi+AXZDf
B7Hd5vAjyO8gqMZVbLGGyhgli72nuPHYuApwcJxnMd6grRl6gZrsutjkNlBJZEV2iyJI18PpqAXd
PpcOUS68CsJH//B2hNs4QNXsuknVZXDrj5iXr9q35kDz8L2ZSuGOvaaE6AaztmFoN4H89VZW+FLa
C0Be+Zl+IJTGyVrUVFdl3n/eQHRiTn+oI0yuX29nXv81FWo+SR3wbbcNUvUOAWiAnfGDa593uPbx
mzPRdaPNn5jFOBjNyNMdU/Ps57m2eSOqc09fdEUMmhAjrRXwGsQH+Jxu2n1WmS8b86WzesgVKWXS
aBhsho4E0kWDmG+CVHkbWWfonbr3H7fcVOzQVXkl5uZqINNIW5jkjtotdbbur84kXS4q+PFXErRv
KPFpn3ucPaipO7Ils5aPStOAje+D18ZhG+dIu3Ahg8tLOOHw4KTSVF1SAPCiVtluDwu8tjcBjazk
OiRFQB2APyi5JiNn9LxO9WV/oKtEKh4pyriVIA+vQ4y6ZYrBsnZvjSvi6cw9zNpuc8/sT70Od+jV
fG6X68YNS5rH60OYYmu5P69bUvDbTSXQ2wE/6Y8a/2eCHSqUrET+8PtGAxVOUyGRdYJFwH1YKXzq
iurk7uhTSCIv1l1ecBAG75eB/Nyfv4/N9Rffb4AeN85bvR3X6VHYm4H4qeccOb62vYkqQHAOAkKo
0q5rJJVLMd9BEmUtlM5JJ0JRIPsTbCkk+zMa7Vp/79295UG7QbQJbL/0A7pryzrrkdeHCZmBI2lB
UJ0Vyiix06xXcy2IiMAVoVfLDqK8zwVx+8ldTbQDVy85QhDQy5NlF0EkwjBgV2znVxu7Y6on8kXX
kcHY+NtVXjYDDfdZJtIcUBavkibtpv2yBwDhIBwYwBdRX91eededcXxM+KfEKfKtidGbnquinlew
ncMsNJmbdhnUznGB5l4Ant7F84I1wJDMP4Uq7wlUaKVle8UnKonYUaMM1rblFWyfcWFCQKIBY8Le
6rwusC4SP6VStXJ4TiBzN7Zb2VJ8sDdV59beWSt5u18a5qheHqrZNOYM42pYkyk93J634vXIj0bv
vFF9HZBWEGAWrSdu4YKGtf26q9Fvhu0exKdUdfEQuKWKDDVOU7n6u9G5ux7ojjz51gm22GJF4ah1
p0xIqSbEMFIVA0txy2R5/JT2YK42zbeAWaDKnzTpQvEeK5fpPBmlnBDWcL1wdLCk/Pl/ZwtFhMRm
MLbX4a6Zdwdr/uxt8tqW+oSn8W5yXIbyb93ReJvmCP6TFHZwLAEeulXvu7RaMTtXC1G17H2b/uuP
Ayy6v5wfHl8tLvDdyE22jzhQohDO93ty8eim9QPg6gv/3TxHR1l5g9rlRWOaghBB1XzxbxXpyTd1
JeKUTmeB/3x5IAY+TfdpKxleQAoRN/hXbCjKXM5SbWxIo8XIs1WmVbMReSuAeFtzYIDAH/HhMDM8
PuASl/wP02JXMLyG8kkjTcMeBKR0yPh89GOleDPU+MKWKiTKfs953dUyiGbhNkpexfYpiPLhDVHw
bZD/jBvpaBK86GBNFrmuDk1xJL/y5CIdnWJGRlejwIIrKjg+qOrTqboXCBWWl55Y+2Sv9JPqBr3k
IB91BaJtG4XH4fxfnRWElK4Q6p6qoMRz2jlhV2ojgt4h/FQCsgOnIzYSPyMDIVBg0Lz32NYa/Nkd
m0Iafkp1CJhawon3NjAVajwa5yKkK4pqnDtTAspefuIkEbfibCbf2VS5LcUN2pwJhac8gKb4NQdP
Ty2pMYTEHRsIhXR01ph7dTHS1jswAMWmh1rZKwjSWK+x8Jlx7HsTPVsuh47+FxpZgQBEuupCNk1t
paIyn96CuGw7fuW67B0T25miqFfFmJ8QqnY7KbzhZnCaOUXLXf+nQQHWCrFICguRSv5v8vmLFK2p
FIhbfLIgjhokQi62OREPIxetLZTH0KYYAm8piEuJXrMo8P0BQxnJJ0fdwJgGUZsV5yHq10f+sfYZ
Yn8SZ7y+7fFAlBLuLMaPTGqGYjyyLqiIAoiHbxCXFoubJoyD5/Om96jgkeyFf1o3p10ozwaV9yt+
BRx3s6MrtTaYwwZNTl6uWria02HQ3vuNUedaWtlLt3SpQsqSLuljcd2fk4L5kWiwd8H6+zDrG8uD
ErDkKgZDPsuzDwCIBvQCAQvss9AuIr+DWIGlfDjCO6jZsJD6D3Voiosb6aTbuoKYUAnd+9J4hpU+
+pGv1Zhto6s5r1Nx+DTcqHhfnHuUFJ4gdYpRTp0gJAIVAmk8F3gXWfxlPLczVvSeZVytItrHnx8N
VhTPCH7Wnd8w2uDVP1QWNxV7v6GKOpGfiWEesJ7vt7bkEFHeIUTceZBhnCzTTO00DT2OC1fZOr8z
cl0W3F6xX6tziXrg6jJ6GcrWzLQDlYHOE7omlWtGwkD4pZTjtWRx4eD0b0x74DujfLFJL848gIMn
m4L953MlF93lAzir6vGpKz0a9L8A/UfnVIkDwCmd9YxdLULA3/Z2jlZ35oXYpOSSXIb0K+/AcZ92
AXzT+PCDL0OkQ+8vgyEDksQA/P+Ivnw2PZHdj1dNssukFFNvTUknLcCnKHK3MlacA5y/Ev/myCI1
wtgVZf0eXx3prrkFxe+uIrs+LvA27p9YE23p0tPD7uVBegmYi3BcmAcEZi/D2QPX8jVVe0FXNI1F
BeY7BEINKLKabhf1WSzIaNOLUrKpooevQNrc4y1Z5Dxonk5pTE1EwR53rN9JCWAIMRyNCBXV5jLX
d2fSPETYLwNtUcgsf6/FUm2487Ye+K+RmcgoZxeZxtnytQSfcZHlA9tiEbJzP8WJVwqHvEn+wY+8
x6mAFJNh3pmUy52wiCmhRbMapitH7b3YBvztQTS8JWFw7PQKZe7f2N2o+F9C1ljyo+vXZ9OTD62K
f5v9zqZEd/bc1QGAaoeCvYtZQBDUSeIwEYyLcQZY25FX+4TH4WlEXrJF7MmlID5ExrD/2Z4bTEP7
qmrXxd0EV5bzAjhteittcE1v0ATydthnyH74kr0w5XiSAGacZhbtCrT8Eo+8MYXeq8jKHZq0Z7oy
8cRYndxyC/GoN7peA6JnYWEniDYrHn9s7hDCY4IRZxpiErpABM+aOWuKXD1f5mIq7Qjj9CQF+NzR
6MG37LIMJpwyj/4Jd1TKpidtVRGeU4YBEm9JctvUYKQK5+dws/ovyrWY+wsQ8HjLs/CzOP5L0fYM
b872LypBtrNltHqTlx52Ah+kbR1WZjD9bFJvybdwiKdw0IhmuTby29h2Tbdcwou98KiRBzAC+yay
S4o2/WbAGuMVJmVZEWfyzixfxUvl3f784Tc5JzzkighfTPo7ZA+9pos4ZQH/Ro4W/2Bstbn5o9Qt
ksKyibfHzl/E2jeyS3VkXtVRczNkd/3J4KCpzuaLCCsExtiyJ1FDnJEvTOmRqXnmUo2CsP7E2bh5
Y2y0ctT1mZ1U8EuvPFJF7HQV/+xl8pdwmcSAa+B24yYKEl/Izofmly+MWAmd/07jNvoLrDbRzvVi
LPcZrFYBU6lJcjrHpPmY3jiDuyn7X+vTKt69n9oaiZKJmuP4KPEt/+ln+AwV++jpmTTKiXeqVcKE
pHQERcDp4QrJilcYkHR4Wm79WCtiEsbgL73zxdpRaMrtTjKpPEFsBm6/fo7fFGKvzyo8NzqpRdqt
ObXwa/e5o9ihW7leP9B3/z3VSeW+SF7JA4pwAlOd5Sds8UfPPGevEWkAq2k5sx9tWYk+IlkNFK6s
HmDxmvhb81j/vf9CnkWiaBAAHS1iBdZRklWUccCKP+9AmvN/UgdZYf7tBDef18rZFrLCEPwND/hC
djcnS8aFzaB0Eges5Rznu7N/q5vG1z7qS2CX3rJf4HC8nPnC8kJ8oYp0w/28b17jhsrO1mOC3qtm
BaXwy7gZ2ltquMOZ7TX5b3WCm5QQuSGhHl3NPQziaZhJ0HDMnJClgNiEImuJczdjy0m6Rkim8KmO
fRxzLj2CDdG1TLEN4pTSuVi1wFBgXHmJ/xeWJ2fL05nnnijzBiHjXs9S22hRZbSfn5V2vNMCreAq
ip/KE0G4H6EplNLqx9rgWzjnOwMcyMaMzqQZOCIHNFaek/OTPmTZKCvSCfpIG8BlxRqj/BRLORMq
9ulRCGfyP1YpKFPI9BIb+CKFge2Gmk9BdMfAsEp9+8kBu5uxn3n11msL9ZEOzBfdMj71DqV7jO0A
dIzgbRtWiXjrXFaqESRrpkQPrYtpnnjhmoHu5qIQwamFWgk2FJq1lUtXKqM7PZ51H5p2rkQsla0Y
o9vXt7fxdbnSigahY7xp6aYboZBiDopaCQe9Di9tRfwUIqtQ9mBnUwwyZyf2VIsn7pwkg6uSI9Ij
1RYTJSZm7kwNsVMyL+Fq7rqafju8uEmFlDphr9GmvbmdauwFrxcI3IYn51xJ/ki0kXwgNzII/qKi
7oCkJbNfkmL8wERjPop6S00l1UNpghA5026eLP319+OzvQaXsWJb6U8GhYugFMz2r4WVBFlmGCes
ybYYg6/WOTKxdNfTbsWIg0pthI9GqXkZvr5kbm6M9IZuwgVSCcXWcKI5F3ga6i74euCe60++/3tT
3JPz9eVY9P4FEJm9sGhhxQPNCpHuQrtczqTdv+HksHypv41RvsHNoseW7HjKafV821K0MSSFI+cS
NorKhr/PFEriRyzBEf/mQc8PuClwTgcaxIsojuBq2+k4MVYTBkedHh0IbBmiNS6gbORKzep6YnYl
wopLF6EzslmRr/a4SIwoMY+4sVaU6NMEj3Mr63YFygqOFHmTNEf31EHo8q5N9BRR6STc0ttGzZFB
AVxrVSagzRjEMTdLiTyQroWOBq5/wdUbKQZ5DoNzwrYs9PcjOdkzqz+LueZq4OIKp7zR/7Y1OuRW
FSm4jPm18RrQ2c0ilUPPyubpL63gGr6/jYWZeaxFsOVLZ4EImp1U0ItZRpWHUgSyRf1z7ttyBgl8
R2JObaPXowpUEIlBNde1MOr6X3GStVN90TOv0PNV+rvNMKcL4jEQJ+lPZNZ/BDaqtn3UwnpDVLZ7
Ngb16rJ7EhWmOepiV1rRYpleQIW+vyubViB9YJJyUppe7mWE69Dh8zL8TPwYAHBvScjAJwn2b/al
qtQ/P15+/kZdZSNknDBmcEsvSLF2RDRHjvK4ePgFzXt8CsputXnvK8HHRnRWngib6aZerDgYMgaC
wjfvkSxFkLb7FYT9ONYHYCKMojEh758A6AC91JTjwVGb56+wW6M+STej3FoofzBiVbzoInDWCxFP
o7Oh9/4b+8ojd2STzfH4TPMqy3iZ/csVH/sy78sTGdYJesiWmmTyHrcbEiHUdi4xAQEParedmbMh
vW9U8j6JqJG5aCYMBeqDATCRfesc3dmqU9qNmFyuNI75NsUcrDX5Sl/ipl7a2Ba8MxBNadDaX2CM
XSkeHBvX9BEHsdhks625yUY5YFiHmTz81rqJ/PVX3f2NypNwjypEt0r5Nm8jd0LLqnXtPWZb1gf7
VP7V59r5NdkiDirYRsyYhrYidaOUSp3fOBvBVYZ0R9gK6+nLnbZmTKKlhnpvav2PH0BAJiqMaNFR
a5UBxsFaOd/A8Pv0+YA8HdICVhT/N07ybGku7fGSd3GsS/cvrXEzPMhWENQ4YAer9yjCeXFqQx1Q
Uz7MOsYoU5crkcwZI2Ryyy4JSVL0OMskGMmWcTiW0jSnFYvBVlLuSP4Wrfg5yX2b4KOM+ObKyKPu
sbUtk64dlwyKeTw3fSirSLZ20bEqwF3jcaWduhuoqDEJgopgSig9LKk11/+K6s++Xblhq70Qga8i
0WvbHxSCDkUtiTv9aPXFcwIChUla5i298hjge5HQR5zXqnE5qNJVMPxCH2wceQ9XwBjTQnWhUY8G
xHFvlv0uQIvx5K08M3As7W9Wjdg6VW955cj21vW1nIzuEMJtVqdxFUWENuf6CgzrbY2WTMa6M2wu
hj3E/SYvkHojG4ijXf5Bxu9ZnUqjr0WpvZJcV0gb8H1xpqPTWYn3Aw8pm8cBfSa9i7rIOWVdM3fk
AzmNbrTLvrk4+JcDO+gYnBh1mQC28urc+pOWh8iM9cqYZvSawGJYGNWEaamnqFvxEo4Ov4j6AWYK
pZspg3lsHa+m16kzLgLoaLIEL8pj5KZSWmYop6cjQHoEXQrsiAW+wQiiEQrVOaf08B7FhYBIuDU9
1ZunbROCn0ytuyRp9gM4Qlpt0LGntR4drOL8YMTiTyzzP3wQwCt5j8DUXiTzLVd+RkJL50/iw1Gf
KwvGKMaTXaTIHbZ2atHHO5MBRBZLR/v5Oeh+buTOx65S870VZ9NxX0XpLSgtMulZjfP/ZTrMD4DV
UuMGMmsnsJdaGfrYHp8fbSxYyhEBq5Bn+OJx82I0jOk3r5vPjXhmvRmf/RtilHRpj05gOHs6Rdq/
DpIjXhIZglFhtQLO+v/owEiCu3Lctj3QF2/GuWbghX3NMSrnv5rSpd+fDWsxRrFFPkjQNO4b32cX
7nfqvQqW2Hrsp9IDbx2cdTsD8fuC/+QBSpu2Th/HXN4b1cM/AHoqMyyx5jIB9pORLsizoKn0Ssgk
I5gbFwb8C/gtNyp/R2h1wXRrvMwhbDE0Z84/nxN9/RgQpzW6XxOXVjo78tm714jlE0MH9R7UFIth
zneqLdpaa/JVsU6+TadlCCqHeYRL6jX+zwn1i7fBQJtLl9YX6GpjGSYZEWwlvKtDNBOhM5wv0iRs
dCfJLhrPVJEeewWtE55BcDPXUta8w8wAMG8bUbi7iCRcV/bCvUS49JByC1OEMI/dky15XpPCsMCb
iygod0m57F7A6ZyJqpWIlRPg0Tolk1njnSCKYr+P2/w+LzAwiArOFYwujKwO75NWsuUKQwbyrCd9
iMUVFBnHsgpg4JuWvdGh7qf4FYVzzS1g2HSBlEazmGmGgS7NGgBSBxG9V6onKHlebBYStyYXL9vL
IISII5b/aPjIzLP2BS5jIA6ta1pSXEsyNsm/omK9he8TqKq3+TTucQfgL41x1aWQcPgIo5A3y+4H
kxCozTH7N6STqWfHktB2ugWz/AcckRxaEvPczhrdordefAgH/VqgKs11WxnEPMc3HXunR+VeHewe
Bn40vo167VfuAVKZXmOKTxTrXpGBb4XT4G+XWc/R8sdGXjLWAWWtjF37u+cjzwcqlWq+35gg6zYo
tmr/FoxLy8CF2cU32NKDj6GgcpO1i9qEL4jt2MVVvgoQ4Wa8zOJYSktxsLdd2wq6/U+0GyORG3/A
uCchOwDW8ccqu5B3G+FDB2+a7a/UlnQlPcAaGzdlDcZvbZLLvaWUtpTuQ9aLch0XC8zANxcFZxz3
S09oITLi8dRUtYiDdnCGQCQT9eoH7ZcGpEQVSCkIM8aFah8L0VI7cx7tjlkUEYVHC8t/vCSuiK3E
mVom4ABL+VLMz3dWY3K2SBzn2Ft9VaTat7pwcZQ+XOyoAPIK9qsMoLz6SU9boyYdyL85sZtnIzCZ
PfSQBRgspb16cwt/Ph9e959oM18jpyawn4LEaYjHzb9WFj+JtB5wub46+ehJEV8wAw8EWcwTvkH3
48NVCInsCiWFrFo+rQa6VQMUpgdUBd6074OOc9a7ZC030A4OQoT4OM1gA4g9MscN6OEcgCe7J1K9
GgSS2sw4+whC5dMbMDlKxrPV6lDdk7wiB3eIhHQmOPkUQdON/JLxBTrMwql/HpdIYg7n/42MY8eQ
NUWSfM5VUgOo69681OpbSu9bmlhNAtbzVpKT32Q5eFIqaT8HDGB5BCkFS+jCzg5r5ZyZhMADQbmK
kqYN2oM/BQT3KkTq+c/Ps8E1701scxIQtp17Fi2aVCN8v2D/RfV2fmmAk1f9EQJXG61s/GxDHdmk
TTBVQGGrorDcDYowTWVvEbinWsKK1WBytabcqiL6MVrRXPAZQzmfDDk8AmgWcaG43zKYIn2rkhRa
jhN4A1uThLzPoFNhWn8EfkHzC6/x1yuP2XYqALqbPWBVjNykV2BEqTgY6d+ehkaLz2CT0Y+K/iGB
MgrEOs1Mbj3ywyfmvTCMf1dnoQr9JTmuN9fft8yTmHEkXAovZNgVjEXUxzzDIplREWuwf3CK0Dru
WTrURdS7QeitwN7J//u9bkJr8Da0MsGScqZzZRMUth/2jVdIMMGPlyex7aa0nnhynl8+U8YQlnIL
sLk+yo2ddL2KgIp18djq/88zV67uDYB3DgY1HmvuHSSFXBzrD9LKnmJbUQPk4+uv1MpAypDPDgaz
/uimEKpmF5t4+MxV+ScFTDwcbZKZWZ09uGx9U4MOI1TlPPWpqA5te55BQQlU02uy7ldT02moukbY
2C3FZni+hdBN+6p4BLU9Um7owGVNZqjvhe8z8WUiwu+R8OHUEbf50mDCF0PDdjkSuoIU1VCn+Tp3
sRT0kjgGCxjK7fwaSz8wvrp/+fCvC2Q9sN2Tm1TGfwOYq07yidqpNzOw3JOObAWwZMjHMNJR61g6
WuTJ5/HNdinGji3poHSCQ/66uYYfrOMEmhCCjr4BlvizYrXqXwYKbejivO7tVNnb++Uqh5PQU7Pe
BRaOJM2JcECRhdgGlybwe42jVwppbkt6zSyHsKqbsZjnKeo/WE2A4o/nQ+3nDURBv1DPBUMCyy47
fVEsU0uq+nmhmRVWXWo1v1WNBehtDtvHjcf+SXHgV+pMmC00GVRZFjCYsjS56XG740pHVsZYh9yh
aCl30bA7BeXAufe2N638hrJuyX1o1j+JE+U6EAo51cGjGbArhe+5Oe06zsSIFm0p4lPe99vSpNLm
rpOL2KuOn08jKpK6cANXi+Wsi+VCRBQ/DPng1ocN/BPEZK3Oh5/pgdCjv4gBGyTv7kAZRYg5QY9l
fqbxNNiYAfeDYm2eGCDOsATJQtx1tByFRU3H0Yum5J5AB5GljzNDqnq2iuSNVQtb3vzI1BI92hKv
vMyFRsAEqp465pnbfZM+X5Iprrwfrbe6HnF5pN5n1FKcO+Is4rxyca7n977Dh9Fu1+9VK/HmyF06
YkwmbdfWAVltPma4XzMaOmOEv++QDmNlR5kuzwI7LymmrtCk63AOUm4Ey04dz8fo0vHFT4IMQS5h
d3LUnsTH3wxL8u+VVFTT4ab1dsJMYUexMrMBeWs8CHGcNRY6fWaurw+LlnunqFpDeeIIsPeH2ikH
IzLmZuFhH8IVzn2BzGHp+ECz9ZlVdl3IzTHYLRFQALmEDvCNjCOHcKon5W+KVT/psB9FBi0tLKSZ
vqPRyL/JyKWpY4cMVYBVuMQ1vB6dg0zSY8b6vZO8QmMOuKi/dJbGMIws8r8oT2MiiAiYWlyN3/OB
Fbig6nCXOiOAWb1Zm/WJ1zvNV4PrSaErwi6SNYL0sGT2NwM01p2D96qejt0I/kdj29mTh05L/f24
EQesJafTh33sQIlJIK61o6kIfnqR12lc0mFMm6S6LVfYQIHNaozF3nJ0wxqw32ii+bpAtbQjIm2h
oYEHUwhj5cT7TVFm9ciR4qS/pd8bPThm/FTAx6FR15Z/9uEaRjFFr70Wvq46aESZ/3Z+aZ/YdlG9
np1XlgqFTYVWNZSeA/ihsUda4wSuNohl2NLO+cnLm9LeAQT1P0R/fCeSBLtwSoNhNq/+iZV2Qmeg
4zFZWUcj3uVfc/aA5Zh6vodAxBrqbvq/m8BoCEi8LjitN0A9vA7VGkHcDMhh4PRkk5QS2SyAMs30
4AuZm1F1pVpjif5+2djzrvf7suEu2Q7oenPvWOgZ31Qa7dk7F4mJ8fWx1BlrbVVrpfZgwqU0i9Ux
OP3YG123ENsVB4snk4R3R8K/EGF94F/5E2zc6j9gm3EaLISQOpAp/KyQqJuuLHOTu4OgtecANvLv
nvYEquKSRrL+V7AVF7KUqDjMJUYPpjkg9cQAtemKnj5myqv9y9fHdCy+L9OD48DZIvaFKfdKAzvy
Rjg0wP9eVkwMepRqPIcmGJ/Z1Y1s2dPDFyL5AUSQpT4BY+Jl8tW5UGZ93wcEM1o6wzi4MDfwIHKY
nry3Cw443jmaiIr39mzZp5AYk/9kzrbaxknalPAMzl3m/EDVYz3YLc8YkGMEVJsxZrj8P838AMLy
+BfmKq+dUHs+kK0szS94Gp4RJ2Wcls0Ocm3WFU5babo0DYu/e0ld/w3Ml6OzMg+EodBEoLoJk2tg
UOwJwIlstGvAxWe1WXmAmU+ONdL1ky8Hm37sGOdDcSbHeMEmP8OLB1dLw1UL4BqjA2rT0M0i4vyr
Tfvqv4yIoxwpPWpYE1ji6eREc1HvWfX03bxFRqruAMqecaGtj2XtgZtdV7CZUfOrTjB6BU2hUAe8
9CbbaO8dMpLH57ArulVPVcISHNCZg2dBMCRKwl+4rqRD0jHBPkAdiV04uFCf/6jy+HFLerWiklYw
YCBkSLXlBjoVh/EuzN6j4yG5tEBmeq/OJvQJbW3NQK/AfpMWrI/wr42CBgPTtexQALQLA9ZhNT2S
gyToWA9t8qdfuAwTRT08peEcJ22D2lFJeZRsaMD/ykBiIrPI8MpVXgG+mDWMEQhS+E1BKjB0iLQt
XTviQT9ZbsF7O4ndip0pMsEVhQ5xKrlZe+AohuZ/CU/5LBuVFAVPGNbc8sTwf1/OPdCBoIyozdME
634aELoiVv06DJEuhGRPYNjVh7qVxe5TkwENs5jqSaZwD9H94w6H5qA+01ar1KacVxllFaOZGhI6
IAkBOpIvAg1kDHkRKKQ6Rni+JTn4pRkjc5w2DkYNpdGEUPYKVa0SdSv+GvDv5+IKnkuKw92Uymqa
CRLHgXTQxeLuojgo7opgJmRol7XkQ6Kl5M0U25DNJAIQWgpCX8E/jHkys+I5zqothXMEpUStRB5K
WSjRfn5Eu4Ym5E7M58jvnGmHaP15WXoQ/GbdIkVQes5et8yKU2Nqjatm1GaY0H1smJCrPtgWQrGk
LtxdylI6GeI7b1smxJ65TYjH4Wj+IpWKSiKPbM3/45nF0+CKK9Bt/jNIRBfxAVAnbFzGpbWz9mVX
/rscTBsohPa7lqvvuPoaAqfyZafHpsO8d3PEKJWp6KTPVzuF/sPavPUh/8nRun+MPqhpRf+Ej27y
U794pDqLF0D6+NQT5NfZILyaAeQoaeVxN9MU58J1Z9ge7o5q2oNBGaX5z9FZvlfT40bW75JNMFlC
CMwCDe56iiVXWZivRRhfFdMY9soI6KDUorL/l9sPQ2v6OZz9OEf8lTjOKk8x60XX63xM962CC/+Z
x2zCOj4okfmzyhyC9iiry/iHlXr5l/PWlCbjpfV6h2jQH+5/5CIv7gP/QCLoHfqh3nD1Ovjp7uKN
wynM5+it+vUPghZkOYKX/KMpy9otWQKgBYNqeRMjix9XW0KeUoWbmRgyd2VDskocrEBR0KHw4pnS
irZETiwai45wsrPf7UAbnOfYbVj2bU/5EeIx5XH3Jbwxzdxnb66Hxe+ew5jzarxyi7SZ9X+Mv9x/
GFsCnSNZT97x4KGIYt3LtCUaNLA7ytb+6EsnZiwhgDHf9ZtXnQRc02UJtykhHh4ci83VcY+n7shu
c7NEFgVjx4fC9Xr13TUnTqGwWvEWjCbNPGaymYr4JEwYEOGAt4wgCn8Q7O6tG2HJX5e+mPHmMPIB
/Tstt5os94yKGMzPHgWXaTRqYepqWeyfEsJF/dDcWZTKXX+SkYSeSePQ3Mc+8B20nYEVUqApt3lq
Av3dsX3nM6h1Gza9jbedBufe6tDWsJCmBGkE3YaN8Xz6urgZ2GDW+5QEzzeEXcORDdwhWNPWlVf8
+4UDnzVF/iroyOt5cH7F5PxaUz0GuJ5txVBcl4X/TZNBGwdu44COseMPWDya0F8DVDQo+877Klnx
YniSuXbpuRTaLiAcearcFvWlhIERimJtGIoC7D14NMD2aHzj6fnoM9dsRtBRh07au+AJE7sT72kJ
/umpTZ83CAylIuywTJwbB00XeCTdQNMPHwDToQrucHtSmCyMhb86H5lFfFSPue/iE+3Z2uU5dayL
/32LcoO/SCAjMIAxp5VKIv25gdAeAH9zUThHtfFn+KXzcsnOph6xzHBuL/x0fYZYNV3RKX5i7Qn4
uNK7vUy7vS4orFncaO7uJyKjkHwWuhjKF7fbNjevbxZPi4noB+jAlo1KYn/C9wl/04h0qPAwJXi6
WcuKldqN6pemAO2PCm4+wPh7dFcQbcAN20V1ub3PdYX/BYq1E17l/GPTHN5Bz03/oOu/KokMdchb
yK/igprCtqxG8uAtifVVqs656m5Qv6VmDm8oyuWsWtW+2R1514SKg0b/OFDw5rycQgXFnaRg7ubw
CSUegTAKovEDv9xsdIp4NcK8q8VikcryeT+8odxA2/7Zy4mtxlOZY+I+mjy4W/FQALNoDInraiDF
yX9Rhno8+d7AjIUPX7Qn9CCT8wFJIM7kCcMJVSsbKWhx3p9XChei6Sswg6s8ei5x7C1UdFnRjj9D
ppcdVWwcQsLMtv1bg0ynO/B98y9db8Ppz6hLz+PUExLrjEPSh+B2lTtb1uItYRatKrawVB6Mte2r
hu7xAE2tBrM2NkX9BIjGhi4hh79jBWfmCsMHTT/pf4Dt9OFO+xHASKO6Batp2rBxZIZ7CjIEx4JS
8dEyBvO+kr6c0Wu+vD80ajb5ap5UPKFlYf2xu5g3Ef24d69o5cJraawpM+eFdORsEiWfN1Mc+PZ2
wnn0qn3ZBJMyKvcfdB9NtRDAHV05BliXTmTtiRFdEzC+QzGTWSY1kff5shkJ8MSc1rs8pU5ZX8wf
d0+5GFexdhnz1X5edID7oUQt2wCxxA6wPwMTb+JqnvILvhxfHOHeoz59deynCLvvsbJ9oOVipuPi
HjCyQdBX/oTmsJmzHzMQwPOUekvPlGHVLh1mQ6QnWOhg6G2jBjMNqxTCDXuKHBi6gAl1wEP0IJub
ViEa9voq5Dm8613V2aX52u/mWs4vY+vrqUuDTtGbbbvOM2o8lwKRCoOHOQCSonAteboYG5DLqvzF
BUYqoA4qYIALFIT48SllFDq7tGOdEzs8MIp7pCOAiAbeVAZ8CC0UPfuRxlI+dUeQC0ehK2GxTMA8
MMoNQMpHyuhY9xbrs4OG+uWTa27EF3c7srrgukOp/+d07j+4ZimOYAC1m58Sz/twVkUWOqR0JQJ/
rMDO0UJJpFA3kWEx3Avy9/fy2tZUVFR/s5H/zrlSeZQtsjmbRnInbl4ZgGmqWUOhdT0ECodKZC3k
ZOtFtavqMcMrgBZ+Z0RLwqNMsl/j174kqrBy4ntTP2GUu6gSBNBFDoAgu52Na06FKpNi1f71xFsl
p+51pEu3a1BGDLWLYet6oVPdvYExxnrPmTBYtosfYWOJch98efyHbuQDVCmqNBc4NPngswUC0zjd
mvkc4+uwiRwb3uyY4zSBo/8Wj+rZDq3arRzODOTFwVAG0QfcncJmCFymg9qYp2KzC9NO51enP5s3
h6dgI0B6TeBQqBL/6L/dfT7T1xwndtkNqyNDFc3KF/4kVNxO1zF26i8/PdyNJSCP+PSCfvceJal+
raoLqgf+VkOOltwB7GnbW3qlv5v63o6i4at7UhvhousbOp9NurN8ECnRcH6qR16UrMajBdtueIig
bGHLmOB3QoT0BmWRQP5uEWziCyIJrNxATSSfb1KNJrK43gkVU4oWrbQ5zmnrXMLr9FIaTuNZjMXu
Xqz3i+azyyT5vxhdvztoYLdXkQqKlvX0suCckPEi5LTsviVYZHyOP5fRwtSjpLjdDq1MtSKzitP6
d0s8qE+DUxDJghtVJG6CzIjAquTEYUS+Kdx3LLRwVXzikgbYCyFdwTJIMokEywp0KVgIie4cdpcm
HkgWrw8hnFowoQWQt4N/FdFDd44gpoaP2Jc6WQAUXHEpPHJVRKiFaSc3zIwB03kKgtF8i5buEVC3
LNZ0gbSsXxdFc72TDPvKXrNItVIBpHN+Zwj3UinCm18aBxhbRlmcl3B+5Tf/Rfu67Jt5k2f0+dTd
RGi3DBio0RFsD8RMbxUB3YWkjihKgRTMIy8vrYxydIKeGjAL/5H9MBLWfDVRBOyzSBrV5/oWJiU/
0xGfWtmLAz3PQMRbq0OrAyLSf9oZuOFVC5Fyp6+QUUGgsYgFN3SHd6lY0DLrptcmT8KRtGOW4nh/
Ymm8MHOVRNvc9xvcHK1WSAGP+5TkVSwOPST2SboWusPaj8LK3IaxZ4fSySl1A/KAiaIA4PRkluuM
l0XKa1bFhq1AqBzlFabBbeUFryD9Y4ukmAL+/bcQLIEhr889OQJHCoBVDw3CY8ViAMYY+4o4kBnB
czFlE5m5ZRynVwG0xtjR2kx9ryxGGPvPr+z0cVhR12hcEnhX2OHo8Hq5KUdJpxURgxyH1uVUKShZ
UsuDQKBrz75YbXaw3MMkVFLGOuk3M0oT37KSQy9IGCfrUN5M/82g0czbA0YnNucVi1QzaFhwTVVU
EN5FWH/sQCH7bv8T+JkcMulD9S/2eOj1rkqMlnodRnZ4Z9NED2sE8f85CPk1ufsXaS6n8X4K4c5d
jczz34ZZN6nJtFzao3oV/A3+uk05AjLrNxY2oDa+rDr7zRUoHVjSP/zAVDvh7R97bQWXPUY4rDX7
rPbiutOa9UM0/Pp36T+ERTDkujmFP+zpA8Czop7YR++icxBP/6yIrPrJkEEQzQbjySCurFxuGX9Y
Z50aOpaaEyIPGku3NYCHbX/2BrT+2F8sa4ogX12Dto2B/pAcHDFdYBQwo5cTqJnBglQ88m1iNljs
dosYKZ6wE5FiC6WbAUroqiqLEFcLsd2HMlAuY5KTsaOiZXBvDohZhrc/+wH3ik4wY/oM61ytlKVt
zF8WAVFFa7t2doS1Hh52/DvcfNTq01rEqZuHwLS5JC1dR/EpcPjpvdGr78EQf7QG9PPDcVX2sxmX
/iNSD1flASaF+RKBk+Joe5y2vHbmxO8YGXww0uQyb4A5VTTQ3VV+0Uz/r/tk2kExgzOaUnaZXLHb
xhL8g7G9NVir8smie+zdWDAP3EjRZdbbLCK4HFxreGp+bK2NofmyKZq1ByYvanPLdsWalfrBQb9b
cJNFtH2GjR/4sqvQFZWMsMrBvf6ZZ3fStdyqjYDCebnL7egZWxGoc2nq/tMWHf8Gk4KHd62fGw8b
ADaIL3Stcx+KcYpjxhtBAjts20XXkJeG/lPCjLFWtuYKMM3c23XSFZ83mmtmrkk8/FlzaWLxZEOv
Qs3lYV0yBlMg1jXJIy8HZs2U3rY/rnVFlBHIZarg88XdUyVE7zl4FunsF7zoIE4468rUJKaE5HeY
vvZDvTOobjsafN+/FvwEbHqDSXNykst7xda+VFb0K0iANQ3wXRR4mDmtknQNlr21pEhvyQEd2+IA
jph+NjEuISUusm7By58FLw6foqR1HldI5bSnj8kdxgXmErZMX5n1e0xK/5VhHaaDsxhZyo/ZpBP6
8bmPqL9dkmnY8v3srapvzv2mHebGI7V0as0mcqfOPv3gm7oBLnbzTpovq0WXuV0owCkj5UghJi8X
Pz0aEyeY67q15+nuyB+HbtpvuL/Mi+4E6qwyrnUR261lwwk6Y6N9HMq/bf27sWSDdz5wjpVdzJr6
bompu/MKSTkVfImBRJJhCgreapIe1VcCZFA3pkXmZj9XCxpSXxV9Ar/u3U7wON57lWpHj/7fQGPf
22d1li05EemclZAjRzrBWiIUo9jHj9Y+o430A7iSFgis18QQz7k0xzv+BR57xYfrDrXtqg6R7H5T
DjA4GxVmdR3BYXG2o/4fTlEvXgee469Q2SYmJF+Sgilsc1wnatvFbrFISDwe2Yotrp/egk2TFmiy
OV2L2f4XD8n0BmrcdyKtl73a6Kaf8UwYB4bJOeXj0fL0TsTF7R0OzKFPBDQ5oCaWVojdwd5E0A5j
vtMs7iMZWZDPyIDxIusKyAY1Gpf/omIdUeKncdqT80g90+mVps7IUS/esyLGyjy0sVL8tTnPHehQ
ngIJcgeyR9uWKndnfgw4NjJOgPEjJuuFGtvWNpcFca1F2fbWQ9FXJN6sa8a9Qc5vJnoWgh9q71UE
lnXHb5ozen+SNrlN7fwKOoiD/UrgSPcVPijIxyYa40X8OpAw+P5q8CHBVeJ4jlMv6tIgcTxXeug7
pyVe0yXNjsEu5RPZq0/55dHLoEyd6OoB36kFkaYqkxGtzqWZkpnwwfCIFPjiBX2RfmHfsDKCwSO4
6k17Ga4kgsNvd5PjBNrJdvwTmNE+/0Oq4GHi8OBkVjn6vxWNV437lNomOFHjTW/+GKgy9ls2u2+3
SURko00yI5g75QW14IpboqKjadoIAbVHUUuFN53UARL3QZQRft4VmahkeMsqfPchqKEYHMCk4a8t
slok37lIftFLiRgZHC4dO8WVRBzZDlPa0Y73/SEsaPDGg2L5X/XRz7wSUGhEzGCWvI4wcuu+2Cqj
GtD9sC/eR10bgQC/CSZ0CaTGQFUsztv6otwpAiB//t8jy9B4iqCuSZYGfZ3Q6uz3GPrW3QSjCFpE
Q6dPReWBsODvf8lP0htyybq2P1dbG7A/XUWJGbcPvZAHadLbTe4Imr6EdqP1pWWU8dXrN3cm4bUF
TfgMkkBLtli8zmqJ6Imyz9YYtz1ZHb+8hwVbJGGtPttQooy7p24b2JogLQnWf1bUxfssR9uCakMy
Up82JdrGEZagQiu3CYBpfTMqV70ysQ0Nn8Aar3lMlXwXV+xhpRKs+pOxSjTHRmf7T9SXNyyRReXR
vtAD6uwuR/jbHeCstG4L1h0BF6tqWGGHuD4cL9ACIyatOijZRp56wR1iQXowZl2bjAifP1fDMMYm
kOvuVhD0HftSWg9OIorycdoVpLo5XUivrsdun3cHqXEQujheMQ+vJTwCuibTwFwlWwwBwWCSdjsq
fR/P2rnfBAbuyvc6aD8Rlr0XviW/Yz0o/i6tZ3Ey3Lu4TlWcWb6syghKyqONoYlw2gLtOlHQookR
qtAWYHGryvAn5QVdK+nbdb7eF4CZZJhd+5Zr7s/D68KJd/nv34RulIavw82yUXcrovKVbd8Txz1q
Our24xYIB0lloENK1ZzFYeDxwtTtB+3SiC27Fng70HztXjdv+OG8ob746aigXiTP3Tq/2Ury4Qja
4rOFf5iket+kJ4KhmAw9tu9E5cVwNtUCcjiS0EfcDbks4HMTT182ZdPaXGOI9zfsG/lm12ZIan+M
5si1mMaal6OrmFm79pMZ4BLfBCmIuneWL7yvJw7212gWE/cHlJlj1A7/1BNolRyuBedSAGXNU0y9
KJH/fWtJmWai4fbBgaruB2iROYlVwIxxRqqun+Zz7Hf6SmPpLEoYhzbX+D7E1B5PAfSis6j6cryL
DmH8HIALwUM+3qjzUqS/5B4CHLOrUg2V8EnbFP4II3k0Fi+CAYxS4bXzkLXgNs8ZYQliHBiezBlr
sQ7oVYrW/NZCm82qBWpOG6WqqVaSj1ZWX6rnODeIUqvG1SIb3t0xIVOB3qzpRUPXo1TQm2sA/34F
7kuTlIG7bml5xzaKpq0cINLcp9OoN7k7Hof4hpbIuGQnVHOV2CbVwFTIE5DHl5pnsJ9GOmgz5Zsj
SEuTIppT1DkMvxhhiZ7hYILl0f2DMBktbhTmDuoAVA/C46pJyHMQE7ZQ7XIL4RSs60QzynP7eGOj
84Eufft6ELa/gTwKlhyHfX83yarvRQl95aZg97odEaeiHyuKDvfhwB3CeLoR6XIE3cQ8Nu90988u
m1CPS0aVqBAlXW27d2EHdYl5ZPXcjHU02xa8E2tLB7y6EWUwBCtchUmUvc2PiBuNlxLr8DSbPydR
9ZmwOM5gcneZz7JL6ndOMyGVs4jl5gxfk18ajDLb49Gi3QBS2bUG4D99DgoFvGGDWmoa5/xfXzKY
V9C0u4zRNRjrdnuVh3yrJcHxlZLnnjYXLi42MsxTOim61qUDC3DDcaFQlD1BCS+tOV3X71K9U991
k/sNw5Y/lE04vrIVuLC8Ab6sCa2JMmdz9epvlauBmf8XqhsmuINCEzH9ceuBJIhUdZ95IZISrrxs
4SW7N8DTH/0SC1LdjOgZ0aZX7Ik3GlfhjH0llfYfTcRU8LLaXXTDdAsCqkjimzqkyCuaWy8ehIwA
qXWbovECMERUS3ArZm4AgoxmENmTztx6xm7YuyDzsS71iyk2DNP/mQiRBuwSVL5CKbo04rzAF//I
u754O3+VtcAaew4vweO/DhcY5JIRMY8cBuUGH24d+vNoDpeSAO+FOMxFckedLLjODrpjZqw9QKdM
Dq74B7euRD0RWXrUR3Cygf1OA2aB8ChE9aBhLqm28b3ui/XAXxZnBS5Qg6NTEB5i5kCfuz3AOEp5
6ffQrl2Qlg/0hmqRUCxWRhmbtTzxTnb0b7Q4sutbM1D8DDt5M2nc//duLEWlqq1l/8keRbWvAOBh
EOlhuQMK1IoMbew/vp6mpF6xSxbJLH/Do5rL2rD1SWW89NWTbpZTeIdSuxMo8bC7P+KM9cYJgngW
PQdo+GCPAlgnb0qfuKEYNILJkFLx/jAQQ9jQOYEo//AeVO4B/fD+ZKCXwwQPUxuRxeX6Pk+x85E2
sysNSo0x7demQqHlzelRCMatGFR2DoPxa53ualx9DQOFQaCJAlIaIfFKQ+B3zdntiQkBKh5lT06y
UK2KMpVgqMmjLTlIZ251JutAnbz4Jmmp/Y0idM+9MvWX78weOzoaz/NkiPd6OPAbxCfCmtPA58bx
eGRsuvZnx4F+v/Gxb4LsXl1xap40XssyM2DfcIltRDDFXheCBmPk7tcDkqDW8lHGN8JSDyQVdxVn
rLzthyLPUOnFhK0CvsjhPFeIxEd07Bt/jJVtneQXpUk/+ow04045S0iiSIZfQlMnLUY87OTD7C1p
1i+oRnZ+3sVxfFKQ5uEtuibJV1wEQ58IU+Uim5AFUZE7KiflEP1BQXLRG7QWYffPGtK2eVk2V2PL
KQYyhKwjlVxC5eDWwo2vOkYlWG4Ls0JBcFRESsAfsxIDY05ljKtgEnxVin4QyVUd0QlftnLOmTON
a5vpsIe6EqTZ71YpKAgu6z3911Y6ZY+Bqbx14GwbkzR8VS37dTLRX/WVxI+/X7BO/NiYnaTGa2qh
MWAvxI9Db5FCw20M1V123lAuK25AFQoFXnlbu4J7+hB28I+haQD9C8pKYufpERDOoG+mtRlafYdw
1dLLdFbxpha3unVuOnzfHMAyhAn80WRoDwFepMntYcu5HCgSGRRkDB4/l4MjNfYegDF1Oem7x+sf
AmchwMCJqofAyugxrmaOZo/8sWYqhpgVoqWznqJ/XUtrme/x2qxxH2t59XMt2wh4tFA7Mpj8aYcH
OY8sV5wq6lOUTYEJCDMGgSWrRiC0TMSciG5pZyR42yl+XtTHlDW5xzFi7q7O6wdPURUCNzFdMPrR
XRwzBROdVKAszQ3ZNjOGk1pZ43WxEfWFacYIUw/vIj4gCkGYilSQZlXJPTVnzsJ1tPLf2TeSYz5r
Rdd5iKvEp7Nc+Y7UscwKbaX5uZtUYhn5PrBQSDIJ7KaP5423A5b2eL0JMs2wQpnyCIuzByoivh/d
3SmDtaeWjK/ALicC2M8amHS49gCPXN6S6n4aQ+aj4rgzPcfEPYq1NaTCQKfX+3JdbUpncE6a+0he
2I/YqO1PHqhPTgFlKKGmmJxHvfWo4U5n5Pg2fU/QhC5Fy8JITNfqVqxGnJDeczawdbj0Z1B5QPiJ
CwKyAV+lhRf00ffyTDgX8PWHCxf5O6UrKQ/AsZdjEJ4e09+BOlZ4Ceh/BoDSs94etgUsnIV9WdPz
KWwUlE6vEfJX3E1B3R1G/EvyIY5LCkvbl6prr2in9aslX7uG77l5WjyC2Dwpc8ExdE/XRoz+f6sd
ddqABmCdGhT7cuNJ4beyV5pz9jWR6HZu93mkbfHXyxCqEknRbBR3ekeGB4O4aRjVwahio+guiMZC
h1JCLrjfFghC0shH7HGCTXy+Ste9UO6HuSdQ6W1iwbVZumJTicI18DqE6VkMMxXjeGMYbXhMoHd0
bcp8DyH+eyMsxgQFbHDDWSz70xXZKxY9KewZmw870kioZLTieAnXJsxF//4wQn0bYCw7kaf17w2Z
3XXpOE7LatwneDVHfjxH2HKKFxJKcuZwkI/1BMN5TdAIoKolsdl40ZlaJWCYoqa7d+9FUJoYbenC
FGOnQ8sbcEfndC6p0UrwqDJJyxoS+C5DpAr60XDw0VcjxbHlaFQRNBsVx1ndalKUlmp6T79VX3j9
1Ub3DSHsOcAqqLFtoqBbS14u013BlRfDLKloKRaMqgXMW+3KpSAdjskGjI6PPLnKPwqYUyNhnURb
2/7qpZuLIrhtiHqRrVakkFLQVkw83Tl3cLv3wo/jLVFvT4Yb0bzZPTR3yKrNmOR6muywXhQMUd//
iHRXmgcx+em2hisf23ZzCNkFDSLaiwwpz3nB3lprLuoOMIqsl3QRz24UEAjF+B9aP2xN0Krl7rBg
ybynDhysba60wCphW40RxJjqY1AZNfWVvrFaLxgIwm7NRydtPuRNPGiV6AH6zkNmgzDJSLkagbNN
IBJE6OJnq5Run6ShWAsZXhZ6FMn0JvLrJ3qPpBohL84pp1bYNhCTzM4GbkDQcj3AKTUFeorTP0BI
he5tosG8T6UvyqF3v1Tsu0VID9u8xAfRs86OCiBU6uaGx1+BgC9iL07bnCbYr0kUNSk5Zah9cPqm
ApbU5l4xzwSFoFpfI0Tej0aCV6ONfeHaLiQcZMjgG4HMYxWi9IAlMrEnEzPFKUmV0qcT/J+iEJyk
JJztmEdex2AjTH5dIyykjiKU7IlGfnIXkCXNpdKvgOm7iBopLKgrD/Ehou+++fqOoHn4zXQsMrkj
8spLx8NGWCBwXbkiwa4mGCl7xte+SHIZSAH4P6PwmnjimYBO+4j8eUlZVorc4tK41aJdWFMxOQUs
+5sV3CY5NRYl74QjALa4M3Zy4u3ZlOSH08RjHqLMT+I/wiaVEW0JtOQj0XZ2rHzBwYuv4C7JTMtL
8WD89n7HYafl+v/bEKWFwS66TsTgtv6LlWAyrW2YwlQALNndFTyOvu13e13CPoMBfhNXB7qbZEOM
/P6gRhLWQm/GpBsmLfsrnue1OlhqJMlRkpjw70pcy3LoYUXzvV3PlRlqJnnE5ljHVc0H9wFIhLPF
//ZkfBiAHBM8GuP5IYixXqhUUORwm3JkN0yk7nyGNUMnyBfrh9TW+KHSyVx7W3iXQ6Yq5OVWybI4
TpUc9QWG3x7Zryc/FO+mK8QFQ7jok9hASX3Df0dGxo2E35Aaw3nTbf1qgD+lKc5LzqewLqvdumGB
jfX6CRGP6FdS2UBKEPoFm+rUphF7J2U/o5CgzqetZfcpC9X4Xc+d9tWwwobUlGm8amNkLRUooBqA
kfUnJqyypw0y4VTb+PH0RPjigxxUDRflVlSJXE+XvGnvZFubxajZ3QxQ1fDYjRwq92zV2LBHfWps
HgcSnWeZpQ65Ni8xLvv+AZGK4k/BVNqPdgiB+KxzeTXCFep8NUmTTtWhP+BOofPlgJWudimVCy8M
rqgTe5NKLBem4WaqzgVQ7TtXgK4qtgiADRoXkFJEAnQUtkzq8xOSzFXTndrm6f3logLzJ6p19biS
iTtkMGq31cxi7zwUgb40zX4526YCbZWylob8vJl2ED5x7fJ78Q8Pjg/l/s5yc07VuTNQyvZoZGtY
Apn2O0+xxfHIf9BLcRH2LCMhdlOCn9WLwbuxFznGJftBYT8bJsiHw7dGWQ4tMiwtzSvBo+A/emow
3hVcobusgmOC4cygSp3RzN0640jUpvwsRUuavANLbM34bGUucQUanLVkRi/i67rkhUCnfBp7NQXw
zvMlZLcOi4BwNvIcRcJGFER24KGHSP/n4JrJkd9/n5OrELLKc+ivWvUGweWrNKCPD4+7PC/wwWfL
G4OV7wiYSwcksogK/mfU3fJKko1UvDlnawd9oKfzfi5icF0GDh5sH2oxWDqOM+GIiIDvvnNzSENN
uRq7XPVagxjpr8ZTHcKO+G4aSSsvsXOmQ2mtO+2L+X8+V/fZ12BZC+TuQ2pSFARHa4y2NLc2m/Ur
3khs2OHkuXveaUz1XVeq/b5dIXln9KUL/DbBYEaYyadG42hGWseT3AI2UhEd4QJo6g0hDbLyY8Oo
lMCbl9iqgEQDs84OXWbvmmKKvoKH+5kbjpymsSxuTVQHBV2a7THtg1QYEiJy7/UBrIsHlLnFcdgF
DvoHSNm71BRtSwHbjJL1BXvmp70h3IH5MoJkDxag3xhlBZtrS706T8tUOdR4t9Xl+mM0ePbmnphz
jtwGLqMjoTFvQhuCWtKpXvHGX3uo99M8X+VfrM9BtazXV9Os6MCkXekXlJRRxCwpo23rES0QN/ey
DEU15+DX2BkTBsuqMSifutfI29K4yCzsNQI9HHnJ+VujB80/Eg/pHd7UwdVBT9W+bFcsD9nxFYkO
wl7E7XAyK+IGASp12RecGGwHfi6u01ZHeOI+/VNgdogw68SinhizeKjkIwM4qanIalmhHJu3BUT7
sOQBm95T47XE7y+FiaixHnvWWCqN1BLtjItu0oGlilRHpKdSVbYHcrUPJA87seHQJ9GRdpaAHDWQ
rFRH2khIXjvaGYLDbT44IVykruvYUiRO9UTeN8ylK8bk7pm9rEhXcH64TixoJ0G9kVfyimxKQMAJ
YihJBArEPN7nPvgboL83q6ylWcLFwBzwg38xN+YoImeisgge8sOGDXcFlAekdq5XYh71z2lVswmw
MbqicpE7WtQ+xQ1B6X+8vrI6i+/qOQeL5l97BQ8dkWvVgiKOgY11Ako5jZiOwTGyIX1KgMWbDR04
5Oq07KsTBOE0TTkuUHPy5T187G8zrUm/79cATW704mTVCxr48lIaLmBYQs2M7+Kj24l4ZokLsCIX
t5a6jayLm5NVdsDBE/VZIHeBwl8Vsd4Vr/ACDl/VUV3t5yApqp6zemT33+2mYUehWsnS/OQtelIG
KoGrsLbO0W3ljCtZHpok7P1bjjemcq2KhDOipmGjJFD0elL39SL9LXisPwPTyafnqFH1GzJxLmMc
DWmirSfWr3wcWkbP8PtXfBcHWj+05V3H49eF07Bx0Mo01AViTvOK6wnrz46FMahoDhnxWbmHwN0o
rG1s1oXLC+n3QVc0k8EPje7V+m24BayHXhzwEkynXpUGrI326YTGc0yv9rgaiK4Jd7BzMNMfpiQc
7Fmlc1kkx8vwWC+wiCWkC2uYrxwGZjn75AL8bK/gW2K6Ll5brBTPw/xhZu7GaO/0XscTqFroKtyL
a3XtGWWrdAN5/KMsOuUqT+6bIMGBO36/U+oAx/OYdzHbQMnmTXZ9yCsZGF8ROkb4XuPP8e4E9nBo
yh35t/zj3XA46favpqp75PPNlnIO7303nlA4tOJoExRRQOzNF/DSJvudSE6cubJuL0CVCdRYfR39
d7HlItVbg2LlAjvhTcX7NsvsKvG3Yd47g4SyXzVh/1zXWSCNyQe+DggvMUma58AzxRMFLHx86Y0E
pIgEugD/Bm1bt/stYXVO7bxqmFxwjeAWZBaLqneYDBp0z3Cne3H8tJddAkiPvxD4o9ZD5l99WPNq
zZfwwGFlK9+/cMp1aXRNUf6/YVTHX3iQt4EV734iNiuFHRHxGRC/GoH0aSIo/Fl/uUlq+zc1i7HP
E28WHdTo004CIwJul1DeOb6nKBDgYRpbCbAvHLL4wHIjYF9ZzOvgFUfFc22BhoO/Fd8KUxoNHocZ
qYvYLah+PUnvZnC0yyh/82tsFFR1EZsR5Kt/EjxP3A/wb0+7hhx5Szd9a7gM05Tub75i7Nbzmw7o
GGnOYkxZSVJX2ljgoTp7qjOJtx2B2BYCa9huvwQ0RL1feL987cyDXXWCMERkUW2wkpnILh+FVgeH
FCCmMPKluEYcIl7n296/QUlTl0MFXvoLgVQ+OAzmTHsIzgN4P6nxtL3UJOw1bveTgKWE49xjPBLR
R21CXqUrNGHQCjRuoyYuGOc8ISexiZMlEtUbRDehpZTHzHmzTx44O4e2Gv4QN9N2mEUljoOFfnk7
dRYCyT/mNkwHjCGto3fhalsomBZCFGlbKR9hGIGBfM5yXiBLkHMwFP9LhepPHEA5vr17netL7JZD
kSzLCBPn2w43aNC/mmGjk3xnGyDeN6JOv6MNZnwyFUsZE68GENznLLwJqbMluD/Oxy1+G7qfDfCN
9HPt1WuLkmEKmEgfxf94diNtWsnxOjUpbIzy9WhNmOJ2rHYZu0GA0ypmPkhNpiyeTFISVl6caM1I
fDf4jVgO77rtJbufdsg/BGvbFH2T8F7HX6kZT+YRrnwMCMZpTo19SaTkwrhgZ+bPlvEt5YEp2zS6
SB0blGju+hhxhB+8TQJf1VGJ4VEA7k44e5VYKP8LoMz1DgonaDf1p4Pp6tGzQdUTqOWhrJv61sMa
pkHU9//amnF3WMem9OYzlq17lJ0mD6KEqYsdR2L2obskYHFvatDQG1Y3EHEr7uUnAe0k41VLce/n
ev6RhoAQs43Gjeid+d48XL24Uw9DlxY/uOYNCmUeYNszaxx+oGsHm/GMjiuR9CSBFlh3SUGaDyar
tMcFqHQ5UDxbzvsnb3EDeCmbBX+MtoFAA0xqgW/x3UHRqKFkEiltdW8Td8tlmv4KaXW3s1V7dpl5
yPnaElaY9jPE5X7PNQKAqm0RDJJ1JOG29p9u+EdCvWyEIhVyyXUUFofVbqJB/mxj0oKJu7CldzY1
TLmCMMUL0Lp/mXUkHnyWMswENmPQaScb+C689BCFOqDldqpKpudtn/vark3dqNXagQIUyX6vDMxE
377f8w7QdNBZzx7+YyS07DGDToEqMpPkwZYDEYpszuydUn/YIHlwcvqUwjz4GUR5N6eO3a8O53r0
Wd0rd3lervrB/4JhUkVWG+tKwmq4dPDixJ1973mAcgBaFeZjqnQIp6Wzvfg3F8iGY4j6sXksgKaU
Z2Yh0jOT+ywOY34oYWpsWq6CRRqhkczJIeOO55+8jbn7xI8itPxwfhR+GUsuXkHGpvOk13j7+fBt
nlKPgCENCfdrlF8pYwA/w817pIhlKOug0Iza9tmOsDhSJ6Pz50swmelnu7XCVOBpqEyvzoQ9BUrE
OUVXDr+BIiN8HyYGmDlLwo8baPcMnN533pl225iPDWTct+5w0XxxMVIzB76vQt0El1nzNAhF6+gm
FG4DNOJ6IZ+qmR2/Nv4QJ1QBXCxqvq0lZbRpLKrEgJo1876Q5uW3A6pEokMLLjK3G9xyZxGUNne/
iRM/NxR4UdQIRQHfHvlVoYkVyDuDwwcEDoNjeOZNqtHytb+qUndovKq7Pue9UHaKxYUUHRLjceXC
WXLKZ9nJ38iVxyTXTe7DM16hGiqJ7dnIdq2v3QZX0x2LeoqvoTKbE24y1Dgs6PUtnIzHIRvL4IoO
6EzQ7Rpx9nBtKke0cM7KUWqyPuCsqjuaFBGRINTLJPUguPToY2oNlIv8xWi8hoI6EBLg5WLMkJkb
It6VCXlorJs7QSI136jSWf+Wry5TSg6t8V684Lwux4rOaEbXGyiu82dTDcXpg+4HNmPmLw++siZ7
bqwOVBAtgBHnCT8FF+y+mfJmhl7nAHCBKDxxoS8POj0lD3ifJXgb3r1qWuk8yM57WM/Cgj8JXSLV
v8+ubGDT6E1QB/nz4UfZ9YAi5mMplF0R++RCvsOxfa6pNkOKZl31jPRns0UVs/vumJ55EryyxkOC
uwqv3vDLq4PjrP+os8pf/NFLoZZxMa+1sinHBtrc5ib8Y3ZHd/3K3790GSVu9A1u8kVWptw8ABcn
CrttC0hWPryyiguCFqSNY72+O+RAkBSwd7ljKU3ms8JGZkKoHe/Y8fGhyVZ9V+notBFWnRFAV2g4
f1u8Bti/iMznZvE5IUDvbKaa0jLh58oAOx6AmmXTNisjKx+D8jD6mfkc1XjsLvOOKuGNbiJc2DpT
+tTuXHnTt/dBF0XvTt0W+zuoIkpBG93auPsC0zMnaN0vxU4UfnmSmqjlLx6JEThe3Nwt2ayaHAND
742WWU3xEXtA+5t/ObiipSr23HcZAd4YfpFMdkyLK6UroIIpSgIr7P464vmF53cRuJB6JsrKoC4p
MUhhhGNnzag4nnYEiQnM3lRG5J2FeIOwWGVHMCUAEv/Dr+4pZzz/qGQMvimTAKDfVlcB+TJ/SSju
owO+eNQIbh4/hFqTpYbGF+pNMqT2OoLmKYdD7KkdTjO8EFO+nqxe6jnvgUynOZZlaemmNrpnsF7R
pv3ckJgaW4NueWWW4cZtxZPIepNnwuPrq65JXomBWk22Ip0PXMmLpo0V7f/IUi/4nFdVGQ5BDLaX
gaCLkZaOlV7T3h1M1xkhaDkAhWZ2xc2j7DyS2rW507/8n5t+eUeZh2pim2/UI12LHC+2rBN7qrXl
m4eVZVbhTmuXQdUxoiP3XijY428DOoTXWgDhHye9iaC+udN/fQyCI5YOZMhwsoKk6WkvhkzkrYsx
yJg4W/NeBDZC+JFOHt62SsLNw/z9KncQzQuXGKGTeNiCMhS4j2JRceCq4QgVOwNgurq45LNj7h3N
EiIplEaKpSuzViBg/6a1x+Fpej+ChoVDLCNuqOkme8zkkORG2dcAlTB05bUNm5yrBxgXgFwSysHt
kwEMptsaaBgk4vgHfyjIEw8ODhPgHj28FAi18tWvE5UOlq/i5rcOcmyp610wnlph2oybJd06569K
0CpzWdkoAu1UUbvqOc/kvbZBkzYxRwzH7OPycdHjz22HwGyqGE6TMMJPz/zW4iwGlFtU5Zjx3ftK
86ghiFe8/e/bdmi68ym2axnXmH5CkeuqDkFg+uhoctG1nI9bPEth0jvRTY0R+03qNcb90ordcqlT
tVRoJsrCfXKHLVu+3/i7Ro2l2tghzoNWFiqSZJRhH1uGD8qOurxp/KjTK4XY0Ocv1CSKnuquWBWh
BjWIxAi6ZDvebFSTfZWS+KZsXyhhuPqh0QaFU6pCFQiCcE2hPaPVxG24owWLAUmeZQJ3STLvZss8
CKv+z81mznMiWL46md0Uf5+D327PlerfIKkU4CDpusx/9a0/3PAEVgzdI2/wFYsgJibcrpu6ptXK
aIGq58T3m2Y7SnjORJu5AYCqFG61/YM2S9WGfOCWqrDwug5FmZWnyjnH3btULKXdrRGuj75KXiyc
14uaj8JKCYGRR5A7L7mnxsntzVhWUZzynVTUK+nu5wIzCjyMQGNtNS/h1Ayip6SDM75QwAisZOGM
eHpF4J7xDCkhi7Cj2OOEbta5o7ZWLLTNT9hi8azoiJO5021zeSVO3h05dKL94V4An4WUQe9QvdxM
+GdAZwNGQWBJhroQiipl8HKuh5rrHSYMK5yee9yVoaP57kMIGCbA0f/8A9Dhkkxzw9a8UQwHvZdu
7fPLjceWuutIqRyCszzPqlW2hPxD5zPUGbm8iVBuV53I14oW19e9XZiftGV9V1p3UepAK15J/RdX
TK7kjBetTSypXqgOLjDd0yigC/yRW9epWjnlB+GhGmtuqPpjotqE6m4yQf1U1TA2E9fxJ3IjE0Z/
knU6h9120wAJzlnvx09nTLVpBkrdn3primZ+9RWGnBUwg/whNQCYyrX59TUPnCUiAYWX5tmpWymE
2y/WFrlpon2J2W1k2nbKNDmIfPGSj1WlNj6RVFXfsLCL2AYYDWIdRh0ae4qIwKuiH9zvycROLYeJ
e2rbkvLN2SSIDWfaCFXW3KHo/bkxha1Ub2uytg8HWATRLT7f+OXT2KOGwOHBMWDZB+Xp+JzKp226
YEuydWIuwVGAopa+kkfoeQ1hggpVaJl21zJ2dV3Q5SCk1Iu5KG0Zdtb7lUYCNuQ79zs7Odzyx8YG
21nSgBwZI8EosZw2uw50RgiESY7GaznAs3nd6jBOCUGCKpxvdNvWTT+SaBv6axv6cXbGAcTuVCPw
9Pd2prvEVp1iBOEAQGfKZsZ/u4t3W/zWfxYIvavFzkcMGnLaSw+lousLEJnzPPGycKOdQc3cDIy4
1p2I9domANqfrFpnZIXMzKFaKsf26V/hj1ViqLboP+tkKR6axHyyOeOTUOBg6R55yoaw2GWcB+F+
TkVD4V3QljWRJBArw2e/+q1zbUQ3IdFl9I0J9IWYDLdGKDdF/c0qLNBWUEVtb+HZs8EppCIjIx5E
Z8i0fiqIVFIngkDDsuc4KDDj6rCu5XQuGxDpZ73YssrnZw3PDGQgtI3Pa1DaIrIX38g8zXzJX7lM
+i6KbYzZ07GRVekv7pSUGFXZNZgSEIvBSDYu+6V7j6GOtWf+ufmLEWahb4FYc7MShc6xoQs7GcTv
4mPUJo6hvkjNJGbvfKk1/n+BTAPsq8PfDN4W5r911Rlx0eALc1s/JP5lKfe4xUuYJX/tJ6OfLc93
JlDeKTHfto1/p23Ym7X0sqTgBjnpiMB5Inym0o/EklNQKejDEyBL+rKa/Zd4hBewDWf+Mi/6ag3d
4vqs5hXwP/aK9pb1Q03EixXnKsTP7BRtRY6onAv1XAAZ6vtsRvR2HB/hmtki0uKGM5CW7HdiYMoz
snGEzuBfdgQifMEG3hHT1khLZbMQRgQI9En5GJKkD2wVquDQSIYfAK9PadCr6oum4XD4qtXU0PbS
xwRZ1yu75++QWTKwCJXp4Um+RiMBHtOED5tLelE1dzrsz/AtOEaOHvunIw6y690PIdEDXsRKVxXr
gNmxYhC+ONIYb6YHxd/VwHndzwqxYcY9k3wI0ki50y/B67TNyVyP2oCSekeBIQmGOfOFrJcBqQ03
5bycK/x878dujnpi00Wbtur9hbdQfYvlc2iVb7zPR3GPvg9OP0+7sCYW8iEhx8c+LUsQuS/F/9Ot
//g28HadloBapLaQ3p9c/hRWtnbG2cO9c2j+84FVOVKc3OdWLZysFtqGcXkHc3xumfTdpkMBgs5G
bLBr6zm7MvS1GFtuAPtk4EH1Hg3T4VUNh8mG49T4P0W92+h8bT3skVoPaGe2qRU/ae741QY32Wjk
KyLa7xYtavQvH7NAF3llRYKMSXrQNluxY3sysvOKbCJoGmoD5W85o7kXdn5tTjM6B7Ado5UTq0q+
/YkxypK+hL/aIl4eu69Od+A0xQ+QwcJsUxx1vTUDvWS1ohh3v9F1nPgKwJFUzOswK+FrRoEV0OTW
SJGeNKzvNH0OmcPQS7WXdybXUN3IfhIhVywSSuFmW73dSnyNzS60Ov1Oo+Cbhh7cJpudzvGPc//X
9vn330ZwOcFPWEZSU7TGKPVy3VPhSSuc6BiV4yyFiPgblg4Be2OHZQmDdR2+dRNmTpOYEn5Bcj22
qCUu3cyKqlfG7RApjFTAoODZTQlKWGMUkm/ScjX1+qFWrtA2uLPkHnfLyRLyfhgtAiBf6saMhCud
yW49yNQbNM+oihpvCAD671Pe+U6hKZCmskogQmxiYjIPi5VBlgXCUOiEeHqHwnbMhghF53QWGBiL
4+E7MJvC5CdZce4+JwbsxNwn/5Q/f7MdreVRRXdLvTc/buqEBiWILbFawh4kdSlPx4MUhX9tqFkw
qrerF0QHm6GaSbR8Rn9Ht/qPDrLnmemsOytUhyiGLTPZG/vgV+8sqTcOpyo7sLAWfiY2OrJeyOwH
GvOgWD/wSFsDSLjHeW5QDJTA1a/S/OZs7bj2Q4Le09SZojdy36Cwc4aVEiyJ60YamO7jbcYoORXz
c146qkWmmOiDjB9uV7PG2U5PbSPpudhRX0ivdMXAQs8QmSxvIaRmOnUxpcKmE/08Wk67B5RH0KVb
WZ0f/hljFOWCxflKUwt6QMEr5/teBUjERwqMg/iyUR9WUFiRCdfTxq8Em/UUFUjgQmUJet7JG146
Yn3CS6MucElm/soCCMimpjUHydCmr/h1lpnv7DPShnqemtkgslbY5ZRil1xKK9wUUc3HwhzSbxNm
JORfOUwTRGJ5nLEuwKz+NA8pJNhfUvUoQJVNwi6fmwrjikpRSaqTO+CgjxRDVuQNUF4YScOixcrW
rSt/eixEZhh6cUO6lQxkoMX0JbgzlwdIhYJM3wpqqIUotrzrumovWcNGwyT5NTK7SVXT/RDZJdBS
py+RNrfl3PiPzgLHmLW64gg/12BPmwIDgNV100+acyzQu8QmL2dEYWb1mI+LPpflOnRiMhsqS0JM
0dKD0mqirJ4ensjATCjoNCR2W0U0jQ9rS2KVhijJmqUCQcNI+2lmVcUdDRDpoSmbDOKeR1TCDUzQ
szUwuljwtVlQWaeHKQ/SQkdOhannNTGsTDLERyyXun1VgauB5zQ1nNhfE+arHnBEe+oisbz5opIt
dO6D+ZwLk5JufPTKLv3Bv//3G0aZF9P/P6p07gIPvb/VnzkYA0LIxzG0I3d/6a6dcSuebYtr3OiE
l151X+gsFLzrWeo9hjYeKmKDCHDwhth9c7ktJ+Rsw/xRhTSaOb+o/vfhSUglnvmsHbnhwTb99kJs
YWufDL0hHJO+Xvp/oIgOKvPDZCzp0hpJw5Qs0GVeuPXAiYi7EvogAD6cofuaVszLHyDL8b6x5xC4
V2PqgoMHPbDG0WkbhWyHwufbczp1DVqW6BgPUN1sfF36sF7Gi/gIGzWdKlTsut3pcu+L7r1eSXeU
xdlIm7tMqQlOqw7agr0p6ozxfLID+GpoYUDpBS/1napAmUKTwyJlXFdmwtWQ0iYxUnRINVAGWbgA
WSUogg92eFq0HmRdTOHgKZ3H8RsxYgGZGW1PaodZvSPkn5iynKsG1AUcejmPTSb0ZPHKrF2+O4cp
4C/3B/v4b3HOO3EaZ2MAy8/00D+CJEecn5lpUfEbTH/Zqh+9PAVktsT4QbYII5vOpysofx6WIX+M
xcrGhlqDjzv+zHJPV2jv/fpLafwoaT5X9+D0xInqTr1Fhkgc8y/cbJI6/zywJnbxo4B/hdIwncHi
Vo8Xtp4RdTAJntj20WFUVh/HNY8q0MPJQuNPa1CW9KXzPD+Rw0FZXRUduzNgEE820F1V70ycpFoN
K/1qu/wJkWd1P5CmhCJD2j5Sbri8S6W28YLXZbpVZfnmu3Ihi+aFhveF98XFVBtM8/1DjzgcIQuA
XApG/zubHO0H8ODECX77HxLF0cf15ciUAsLaUkkQViiRkTi+nZqgxiUIEk7L0JW85NvXa/BjYLno
jTBMm+EMA7Wp5ag/fAOmKkxKtvXkiaiE+mseLoGp0zCmQZOC1SDX9GGih5KnCvYyy6RAC9QXYdvp
6gMWNi9NVpBMx2XaGSZ3z3pUCvfRFHKzAo1xh4pLiOM4KHvdPl4+Bf+EWNtDZDBpZlFdvHGyaJ0S
N+sfSWferJGNtNTE+s/EuFcMKRjxDpZwlwrKL96EfVp1IstVdLVBCZhAkHGVQLMEryRo5zk0Gn8J
c9QUbpYhla45+xLlY9nTiaSJPAHHn+Q++Pkh0M1vs6mHLQW95THUYIzS62hPXREuaadguPIqa60J
wvWBRhXXgP1s/nFMcvuZdbVoyEzO0T2nShz2zzfWmNJ+gp3UTnuIPH1+qe10dBiHk8bJzG925DtW
XyGEbTL+orM9nirWUUlwzd0PE8HOKR+d2oNrfuL7xAsKra3kNySWSSudsdWuaE27SMLBsVYtupBd
5CcxnK7fwKkDVMP1Kzz9+ulQTRiLBqOrWe4HJjHTI7c3IHhviS0mNwX12wbxIPthZiNHzwznSM+C
5ngpSYNzx4hbuz5WFqUS1vOSZqgNvNIN6vQnDAqcYJbp4gDb0ZcF1J26wqdiDxQ/0TmcXUBcfKK/
jO6+raUngvj9ZpPjxPiLViVTKDIzgtuf/mxI1UXC05dMTYXIRY7ggjFD/OT4dg1r3HNpcHoIli4v
tHhsfvEas8/BDaqBETtmaR8sHt1uqUM4pkrag3nzj2joT2SjMrzOzOEADFbexLwTBEAzYUo80Vj/
mp0U7m6Hw6W1C7rJ+xLMidPlJ04n0G3uS1RXEB6NzSqGcv91kOLOSU00/MhPZBo0NSrRDovph5X0
cvjL7lYK4epXXg0wQgiITsczuP2ff5XsgccJAd7yV6ckpUHeAvwfL9U89wvwRCeT615OvG3D/vYV
5f6vqEZkx6hBtliwf7lseskWn0hkg5EraD2ZZieIWfk2t6YfuRZMAIX09fC5eIPQFDGjBSXSDcxK
oGktdeQzXjMi9MZRFhJZlgnHSckmKZ33sMTTPSCuPIbPZ3VINfVyPTONT6J2AIA2U936te4DYKuK
OzQgy7c78b7IL9A5a/aiebFEIDMyyK6KuLvlUEMgn6KnKe9IHoxa+A0oGVl7+aoUq2KxOvMSb2sW
FyknhePPS3kRNRXtegpbQHtcYtmiDN/zFdry6Ql+/IaIZkBM0CoZquCHoi8LpESk6OvlimUU+f4r
geScYUkBRG7CohLG9dA6BwZmpaTAl4tvb7x8ulAF9RDjFwm9C7Q47+ohsExojosZNdlXCSCixVAe
qdkJRr18A91rSbAMYq9dOKWZCtyCjH1irbXY3lcExc4MlKlZjmNWG95KewS4Rb/iPJhddfDBJisT
e/xCzXQrL2EL0b4pKbv6fjUDRjN72pIHJMgHdubFoFE0qqdVyLdi65Q4NU86Zmz0+4HjWvHNiwHn
jQCXGy5tXwMPVOPllrCz2mfBC/0ZIEGbwvWax2VK3dyyBhVslNnq7bJqPiv1GlLwKavth6hgvW3j
vmf14h2Rj9uAR+/6WtCfI+N+leITuYcgDnXTJWbR+scarvMB2mEKSIS3GE6GE+28X9CdZ1P/XiFI
/w3lYvI9jI9uqfM0G0IJrU7s6TjusKplLwCfefFufBcArGrafH/aUrhf7J/Q+GlBRyIuy3UXHZfq
XM2gHWOhUr6J2lHdgJlAwdwXdezFTAWA5u51zs5HnFcfR1ofmIT0jrNk6fmPBZQ2BPvFidpQzihk
tw48828pcka3WgBwDtKG7fCR7f1lwNtocy4+s8ZnJR0avKHegKkY3LuaP9miFCJaNILKita7NBRi
B+ohYHWzz9qd3svhaBoz7AqhZ36U0KOeIWDFzeR+BMVi4lss0RqQRTYHLAY7hggxNfKkWgs29z7s
5vA1YzGzGuvxPlSHJKih/2hTMlpGrWBruQJSGXaNp6a8vDd3vhIPrzF3JSBRHN9kGQnteAr36xMo
vgiDeXmksKdbxnOeq0fJlcAlZLXNI8Pztvpw2IDUdq0hBs4ZnAwvo2udBKviIx5HrqjKTpmLoCsf
fUqJPXRbCalCpfzK6DWAdbqVRsJ09vTzoqOepgsVBEbmLxyGIVIdvNczJHERrpJm+RjLQ1n4/yZT
NRCDjugZMwS+g4YycY8uxyJ3LKRJ3zibZo1YDTNUP67KM6nBcAx6OsO/C4pMhmzUaHwv0AARDdcO
m42LvAiaO30hAfTJD9Gt1rWrEjGz1fLxihEVim9AwVAvYMrHYjZ1yDVQWoNzFXnAG+uW4562kFcf
SezJatzdsSdpubBP2lhQnl5IGOnX/IODLQKcMhcIiu7S6gKVjIpOQJDkXlJb8K+niPSDrgkbzSWD
fTZo6J3GSUhYEFEvYDaotO9P4rE4rFd5FYDj5NSiyC3956LNZ751maeb1qoJn2TueiwPRVqmmn4F
9z8pEiofqP/Smd8NFb+8IgZG2CTy8T16mIZC5J7S3WYh8GoumSIlYynRkBR+EzsKXdWDMVEW3T2c
cspU/1V6jS0AzD6ahcupmOmqguamURZnyCBfulxH1Bx7W3C6RfSagVzLEBqFAJaGR1DOLT5Hecph
RK1Ocynd4y+0+6IAHM2W2I8pNiG1hnh7cGUO8JLpNGsVDHYDgPPb3cts4x2Oez6CAvHVavnLhURa
laQcDeldJjC0ihM/hBz5tJQq18qw/DZodPrC0zyKYZ0oTlqtVnCDx+1+Dc35PQlBTZRjQyDE2k4B
lP3GM0BsLLu1VoFy4XvqRnbx+4p5nRNTiwwsC70a902Pr4h6+qUloYwBWZf7HbCoVnVR9dAOVrTz
cQtTOZVmxwMo3qYA2/Z5CEND/jzAzXiLYwovJrh8Nht899t6G7q/Eroh8aB9W/s8d/Dd0SvT1ZU4
qrkNBixzgpikeX54DaPHS3Ii/nHcCtwccjpcBPDteKnl8be2AnP0xGQ1r9B8zC1HoOQpt5BmtVaU
5DL1ZZeUE8PEVscMhvZQQdRGvIA/kUQJR61XraGXEHJhm4lI6GQeESaf0ILcUpqoNXkHMbl/46Ag
LvhDZBIQKEwkCCDeOV53/OsntdF8bN5rTQxCbV0aiRXqps4Z2+7wYC2YLDWH7r4StXGzjjJ8lQ3v
UrpdU4lBrkYw3omrazH1/yDMo4/989HKU3eixxSdZ9lchfSnibwguvRIb+vXmdipkeGb5P/3SmDx
tMIhpC5yTymU8nh6/mDddldvRECfB3Va248A5pAdAPtuIKYuAehiwR2N50Ck+eb0bknlhezrhtmn
wcQbuRQv9lqfan8q6vR4niE0bCmfPGz7RiLgR2KtKtbnSA7HlTF0ireRX0BLMiMWeWcBRmRVuKfy
6nDv/uH9hoczt1qt+xjk1wi55FDqkMq516lwnjXOqKlw+FxQ7pq/uafVW082OAeQJwynOHgB977v
ChhvPh/LMcMBF0GPocnWvmSXiGe2dwo+TjD6b1ucLCPCZ+jPaGKIQuipETxo9mQ7Lja254aE9od2
HiLXTHi3/xPUR4KJa8ckm41J+sniw8gZSwXx6lNqSInztD5I7E4JXgVy3Y3aD4DgKI2NVAF0CPSv
bTIm743AlwC4G5rNmrX8WN4Uh97/NL2XPpOX3H1ErPaZnjmezOcwYch+BaJNrj+M2FJoWPHWMvUm
2qPN4FQib+HiBZPEk+/IhYPMhWGi/+B0XODlrctK3oMZEJrTvFIrPO3pjLifis5VkErN+ChN3I6v
2nMsFnpx4VHujus/WXiZ3RfjRw/fJIMXvkZsFN0VoMmnccrwYbRt7CqqZAjZRwgr8ZKOnsQdqf61
PPBKyaa8Oj4tE1roc7AQIfmEAL9PX3uvFgLnw5SOZv4XGqJSj8Dt6SZbv2OY7cwq7NDnxA5Ugyow
0hHCXliQmnuRYWio1jXixfpT6eCxKP8IBSWLQ3xQdUBfTmVAe/wN52Vl5rq9pa1A0r1BL72m8HKx
ZqSOJMUKaJylZChI6aXyfIhU+kMxHyVpGHEHsKWrC6USZpBrpaeFWVDH9CKZyG7rSlB89Io8AGtV
1j8WXvwl8ESpIdvJH4K0k8WjmxgO33b9ixq/vhdiM0U4l9RO2A42YsTJBJkV+6ksm5ZDwYG/ZC0w
axyK5trW0VbcDVT9h2OXbCYsP0ZpObeTqUDi275L8EiKz7HNcz63QRWkvxklig2trNKA7+fVNmO5
ZFlH5PXtdCIhL+nJc9madsdP7NTfgg9H6ONpvqPzj9qPjog9ba77b4+pfF31drGcWijuC2KBimAI
6sjLeztDsdR47Lrg7zcI/oK1rbO7USm2gLLuhFpSbaFdQkRKS2WO3MJXZ8l0yGaZPr8HfHby3HH5
soxwfhrjxPyVJrWX9F4B8ytKLjcOrY9Kng2Iq2hVEA26wzZfN+dLxrk3j/CGcxkbgk+682mEylhD
PMqTWPoSuNL8JQVe8oztXzha+sRiB9sxScU7gc6MLsQmjM9jty/40qppRW5ANr+YZM7UempDcQZZ
CKYxxJS3pDMAf/81b1OFyF0lVkcVblXjQf1n6OPLuI8is55xXBLraKyPkpB/uKpeftpee3j6PsKU
6Uwhdb/XS4xGe4ZAnfEIEcW/eN5kIhKzCKV0cSyKcUmTDV5KvqwPY4U1QNHu0btipv9YGbLLDJAJ
9Yo/3IuRkjiZDNuvq2bgvtYJkX2EO6Hy2E+iLRU9Y10wW/qZTg9EupEb4FK8HIbT8lP3Px1YRSUt
sQ8MGnG/z/yxy2v4FfgiBcRw/dGMIr2P1eeE0jISE3XAHYfG+ytz5WcTuLa8PGx2Liop9ln09oYr
g3FB04LfHLnDsySUFmSYLnx63isnAamRp7s/EjMOFRHr/jqHmazbua85ia4e3yieG1LeaKXdt6Sa
XwMR0yV0z2AiESSTQRj1hnTryTbs5y/oyR2ixIeEbew8gRxO+mWfURzxVDkp3RrQmCYZ8AtK1DYh
+NE3lnqrZGwvYAT7Eiw2+t7hq7EtQPGJZFvuMssJk+QE0IgS8ble5vLc+uUaVyNqK9D0hkyHWJHd
mR23bhUUrLHvJZszTHGhwtkIGsySDY4m1dErmQRL7NTGeqo5NKld6jo9g8cG46Vr78huzrMUWwJt
fSg+pmPciVht4uByE4FWzbfsE+WDgOknZ1GiF5HqKahI7UBKvOwFhSSnohFC1GvDzUPqG075Bo7p
aZajFex0bFgWBjdqTDj7i84zhfVgT/Y0FaHrYijbNNaP66zNqsF0XsHlZR/9A8Cs4+nKzGIruJZ8
NgInul/ODP4TVGIJBw4qeD4pqwCVYZE5aNZpF3R6KO2+48UwL4fETeYB/Z0jDBTo7ON3cR4ZKoQP
qwBUPxnInrE4W0kwkmfh9/0xloMFse5nj4DBTgN9NwvyJb2lyjx76zJYqEatNdqf682jl9RC/ntm
Gm9DgI0SQubF3NpXTn9rqtteAfzcqNBQjKSw9VN1DiNgUstQysBKSgNR2YQ9wq/SlMOQZu1pqyPU
v2pVNm0mEVFac/EJrj+BCMJ9sEAwHVnVUbAM1cvElWKZdoxl40oa/q+LliC4nZ1IE5YXngdTWirP
L7asLFOYZMSAfLNif1lIefDehqa+JoDpNMmKbqFpki11xCm6bjga/bdajsvUbWo0uOHE9iUuI4KI
/XdqhkUu6NOPPhU3j5kI5tvj2pjnbSlNMVcj4vdEjRzHkbEuvUpm0Ez1hdtEyMbFcuEWa1h35Pgz
hlW84imzXVY08R2Rc0Q4un3fEPkFn7E6SYbQ1P1gIqDDhdMqim19yuwsyJRYUTIbPTAF5Gm+FpUq
TqActXJ0IQYmIkvO4+Z1zgAMfCtMU3LrDqqu7vXaOimpMruriBpalFY04eQThbqFwdlOO7ldJs7Z
EyVs0MRvpoaSZlqyoTQn+oX6aRzdqFnKySIOFsMmvQKTzlnhWTn+YpUOsM2BURxcDtNnF+h4FeLT
Fy+V0RbGSqHVafRt44IDlORXsy37tMRDUS/4o1yeALYBmkLAXwAPjvxTFUIyuxUmm1tPVusX3wy2
E1Xj1uzxzSnCq5o5OtO5KhhAT4U4wqy21ZSXMTxYeRw6OYciOv5QC+2E2RM3yQL7uTBTccYLw75W
g2NJWiILbkslLFWU3AOUpouf6rcuu8FUC+8F3uq4IgIbr7HjOm1lGQztof/TI4uTj6a2E+ATdTWE
2lNMJTebO+plF0xjYYWtnVdF5v6C1yuyog04/yLPvCJr3TJHP/nByhlbf/yhTabMwk77Wf4Q845L
VaZQguJ0yORK5TfgzwQgGPaCdrh0bAkV7fFq3Gi+CucB8TVuZ6K8P0AyFb5CT1q1TVKkwUAhfljl
A0vZ0hOq5w7ZZXpI2W9Lh7cGUPwkXnLsG2eEx3fjeoaxbP0CmhbHaLAdNfNaYtY49VFaNgp3CVXB
zTQCq7ifU0MP727I7hM8DNxWYVlrb2oVgXJrXb0wLKJYo3gfv5K/tnxuv59fBVUoat0QFFCqnSmY
IR2kVUz5DPQwPZWI0L0efhE9s4enIzQTs4zvZnJiOsD7hWbb5nWt/I5Gh/wtRM5KIP1wq+Lb8xKE
VzUhb7pLaRGpK7HwXuXIvLYJLbx1kZpjwh0zbUgXHByPjlFcBqMl9kJU1v1k8WG+aiyHlrnHeEUT
ouU7H9HQBMgovzovLlw5FaDnhMBFR6+X4ohD22k4HYrSKVzT7zHnRPtxAGSEX+T3j/Zqktc7sdUT
G3TEHqhtaLJgUYJqqDXIzgjiTQoI9PWNT/4vPFwDY9qBM04sqrW4QEUFNNODmtLelKaYnl9+Q9QM
oW6X5INeQKc5c9Dw0TGkpijSpLmsv0oYs4j/sGeyb8HqFBNCWNjONY3Vim9U0l83kV1hSYa6wIVr
QqxZVSwJZGtwKlnbKJdIGOqSvDyo7zMHGApp65V91uSMWfQPrgsQzGSO8NjD12ZA6dwQEDkr2aSH
TV5Qi246V40IS6msbZ/QnjnvYT2JNVwq09UFy8PIHat9GAeCzs1ziX11WsN1Q9c26ZI7YXjGyeDP
p+M6T77ZmFWW3FFAR9YMIhY6V+IzLEVXzKVtmyzCsCF7uJp6iqAyNpeZXVR/ewMepGRwZNBzJeZ/
Il2ZeFYTB8ctODdr61zC43EcNUWK67cK9yglf2F9QvBPqbQbTDK4whNcjirmh6kAyaGyqc+O3wOU
IPXhAKBvirM25hoIE4mqt3pVa80x63feoV9t2TTzNl5/NIxc6aXfjD1K8o3e5zTMRPutHOYVscON
xiBIoRR9pCHPPMNgfiom5tI14czrSnyATDPgmEG7y7RxZfFFmnW/KC6+9Fe2e/E1SARRywocFEGa
ri2mwE9mxLMger+OWf34p3tE0LYL/bJpofVkTBKd28djKuktf3rDLdqBm2lqiYiIPamNW3dTd+zW
Eu5nnTizh3HAja3fhdel6zmir2daC8EFZbhu4pRu+fKvxZqzQGjHqCNafMrAGB2bW1wLIJA28Dvh
dZ82/NXNrM87Pnw6ObEPPBH+rzlgz+WAqUIufkFOM4D+5aLtNRBuGsLBJNLbIsFR5PGc1Q6121mb
lgeNiNO2yVXtXuZk3C+0dq/AVz0v1BHujASATbZdQlRfnU8YKin30i60w1Y7dPhSga/POEUROkel
jlUvkaQlPEjAjzjCSv/JYX27kXunLsJYij3jzHBB6Mv8aTIU5Ot0nsDoKsZh9sHadAC+MehH63/J
HtU9xqDzgPC+66RA1pCNVM/nLb/uEa2Z+ukgk2ndYCS4fgZcmfG00WfPOF8rn7t/+ihc0+iFcT7R
t98ld7DC6x0vkaJO5d/aOBS7DTKQrkzR64/irDXl4Crg+v7Foau+d0ySDnbH4Bn5XwCwRKpUbs2q
VUuUfaERBXCKCuBG3WUlJ+1K8V6R4Gms9fQ2mLLwciQfBJki117PTePZCLu4HyeYu7EFl4CNUtqv
PAls5MWwl0jLBR3adSoZQMpGqUSIGR7dKLdxV9HAIXEzaxMgQWG9ct2sxIB6GxhBSErp/9mli2nl
AaBdWr9o4YhNCVHLexMwqpBx59CuvejGWRaFMWrGgf6zYp4Lj6nJIigxXhjFCBLpuxm+6JidHhco
EPQJ6agU6/z5utOGow5nSCsJ7uyMy5ag3/b9N0cc2qArbLAHKsUGkgLPvcz6RAaqGiNVMZ0Z7gBz
EIbnkQd3ROACLjOj8+2jMT5XlkZnSjc/9EcR7HZS2PjLv68gs1cYpYS6XbzctMNzxchIBsn6Uk/p
6ymGvnSnMoQsI2B+PaszJjmiIOc6oii4LOC6c7gwRMQIsy7jCKKfWIEr4ImSz5E9k0UDj3AAQ5w9
toaaAye/uPuPgvMY0R8b0UKDXkO6g10sDT53aORVNXvmepcW21Y53ttlEevvXQ6rgZLa52hInIA1
7O+Bf01zAGDTphryUtLPewjmfWJKSuuZx+kvt5SFicPgge+HPTJeS47DH4tGQ7fZMNgAfy6OpgUe
sZeTe7IAo72T/xJwGzNDEfflbNz6crQUWNuxUp1a+fYyFfSEZYMgrjvkV5P9cFWYG6Kozm8jwVji
KM4OechNLeKjyTcd7u23TTTLbGKVqUiy/9YPvVYHF9UM5RESl+GuajSPvVlxwk4p19+4MvAJbQZW
aSu9KhnvU8f3VyYzltMS6s2iJrisvHOcnckPzm6Nc5lrefjIcT8P0PTd6Vg4QQyzykftVfTmZ20/
siHU70fCSxLrBCL92fN9Qe9O3WdOfgMYHszKYOXx+izMS+HY3IMy+aW2nZqO78BUBpeH2z7NiPrs
moEIvqGGIipO2apR0/6tkdmDdqh0Jg3P8AzCvr2kOppq6UTyRU/WWdNZ3kxALnqJKg92xkA55rDx
4NgO3tI4rFRAZvfOObVYb8Aj1IWwE4LsgTiJNqYKhcEQ2SxuIGpxzhB1nQx65M0cs7ystPK0wP11
jz5Q76kt5TKsmNcwWe2RfdufkbC0HeKG4GY7YSH7ZER4YtkbiUvGAIQsJMCpMDphOo0wk/D25Z7B
nAY2M2KoQbIcxsZAPxdgnlXxq4jeIeiBxb1nabwfhCm4QhwalaFscJJ34R9eW47zl8//koVY3Fbc
+Ri+2GZgip3KSCZF5urBDcBjtf09w3ApackdRV4rc0mIX5FYynRUGlF1T5WHxygIv2vPT+VYMvLg
S21b+rn2aK8lUibXX3MHAcGiCH7A+N47Qt8xmSenIyJ7smk07SB37NZ/3Uifu2tOPjTKZpDiy+Vk
ytpcUp86KmzAsub38msBz4TZ0C6AUl6gAe2dBrLGWpaK9M5XXiqaU9/uRi0F7LZ3lx83fvsNLNTL
ENR/7aFG5J7qT/6gN955cLuL/RpkJhY8vAm50I9hrDP/6bdPsFM6RzcQu33R1jWDi0cMInSQrYgO
hP3pEVHh4kSXt8jOcp0lLSQFSNIZd6Bk78C0wCX7h4PNBvdfZ0SkQ5ObNRQemVvQmbA0g9K2G+2r
VNtUZ7yKGMWNWQ+vxLlvmfGVolMtucOHO7XvXftzVb+tsoEoafTzqWKZgwyzrU0L3IoJHkDuo2P7
kc5phcjxEFPUCCfu9DPVE95bBFI6LnBP4pnzhVj+qtCkZtBA4rRNVQWTlZ9q9EoadzWvOczpod+I
2Rsj7xzlbat/eQG4AWh6TLS+MQVV0lwuVVs05/kgPPZo2uw7J2/QQJEqQNo8fzjlc+Ku+3tnJQ0C
ZXBvMhCgVUMhtD0Rb/hBEiOKWSjS5BjP1lHCnZhA/Eq3FCWHXXt5AAc6j8WrMNCuu1EcL9AszSqZ
QMChLl1klAvbgI3b0bFNVaHgqwdUlp/v1SB4NOUbyUvIOdLEi1aDSMSssRr8v7LFoLkv1v1iOzm1
4JMEWod8KqiMwGHYBHaOYuTbNS83d9s6bAncsJYHyEXRmMdf6ld90TGNrM1zfLyKW9N6UK7DfUt2
3uGoO7XyQqk0qQdfYPM73dz9bvYAWKrnkSZRQByF2MHGFbJGMbUZsoOoGMoyoRjLJL4WFwkuz+ux
VNsE2L2Aq9OgmHL2nhaOiGRJROS7QYBI8hYhO+G7jhXBB0HpEO/IzBeubS1lrxOLKR3aVa7fCAyF
03vB5gHqx7RWGnf/pWT/pzd8K1BYUebHXhyWbmO8BzrRWQmxiDs3OBR/cB6dObSgjhldYeL8J8k7
EkatCfoSEAHS+5X9tBhcZNG/+luR3yN/ODlBevC9vLfT56UMY8HFMkHmcy7I97r5c8pr4YKV0NpT
VpJcClPkrL1MQpnfXz2shIGCTmaU8Fvo+oDZqbPTs6tEpfPZ/qt+5Zkg1WF3cDRuEnJ6eam7YAGu
W21oKqKw2SieQ2IdCuu6hCFTK2nNmvl0f5G62GQDTLi79M0fI3iukzOzZKQreQfRLwaCHqg4Ncej
OpO888y4kPxUsHNmMInr0QX6YaT3eebngWWMyhELV/1Knnfj7eYY93laRpP+Ihwhd5eVywsW/SZw
LRwh4aP1bpkLAw7RkWOg6S9N/+l+JIrcX6e+hDdiCAZfzocvq4zMt0wCJz6HnjN9yoOnULU5WIYY
RM6gcS5EsGloNnNumltvMFNiY1q40O+nIqkyX7J56xyDnUEiV/w0HzjXtaOi+Lqv7rq85NXZ4V2P
igpBJ7lmagWIW+ai1R8Aqdv6QlwUxeljKEoHJWmVrnOIyOZ+LW4hx8UX/24FBGfCvEoj39nef8mz
FhQ/S9IGcukLVdLUatfA0UEXv8Tr7tplZRL5qBvlJ8jv6Y8DCHNpXieeOll/kXFGDkl6M52OI/Yu
Dh/TINJ3S+9uHiyQiygfAnjChGMgfB9G/WZ2perO9Z1cDb+TmnIE/iTvlcacbE/xWR+Zq/M66xXw
P84CCONUGUrs1Y4qqEGoi7WPHrXsSjdrZI3H2vILuzNEE6ylLLXPOzSfZbIE7B8aWOFJZxZXPJW7
5A8II0+Vltzv61rhfk7DkItEFjeAvXcmpjkkRdzIE5i3LlOlf3NLw6mehPklITHRBIGQLijU/bZM
1MkrBPwzTvHVARrKaUBWuIUH5SIo1couekQSftI13eyf/t4icViT+22hxORCRWyPb19frCyQTYfq
aYGErldTAMLP1c9MbcEPVlWCu/jIGSPNUoz4fGTkHD1rkO1zGlo+lF2NHawzIjkGx/Ssc/YOuhYK
LZMZjdk1qe+3k7lnJUjdeAO7+rfL1nNdFo8AiMJ3EUdrt2C3ldLQcDCzIKkEer5VXl/vEkceG2Ax
8JjHflzp/NNPoIm/sdzAOH4C2FX2P9WYihrjHGJ+Ljn2b7aeH96wyelHLQwiXUQwK/YWxQHpY5m3
Rvtz3Kf/aHPrb3bbEQDLK29HtJEc+E0tD2C2KmmRr3d6s3pdLFxU8ZgcZPiYQfclSPibB/RHm/qD
FS3aZcaN/OEeONxPLx2xdAtSOx1iV/bKMsP90ydRIaX4p2SI9Qo4tCVGi+NS1+k6+wyrP6K6MeWd
iXahzeFmOiduxWL15q03eNS3gPWZftR1JYR/X/p37wDmxmr/wUgIlUt2Ob4di6h3LgfMytU5ZA7R
8M36YL4h98Q2jqoad6VINWkf5D0idtLsw+4KZZTM5Jq9y0F15HwEWqu9J393U5T5y7AfwGNZJQ7E
qAzqgrnGQX15MpHN9k2jhDjl96+BQBiQB6I1IHSyNRcjvtdLA0M9CRIWZ65iBaCG2OKkc5YNS3Im
bZkiKwiYqpBdriPq/0cgaJMOA0Dk9LHN1BIDPSj2mlyw+VSbppAIGw3gBa8suyC3FOu9kYAQq0zR
XMNiZMI0nFE7mFG2gDiu5E2VYBLZjSAvBeg5B325E5UoQRqJFYagv2JX/KvT3UKWxt/PQIfuNget
OhYSS5JlfLxEqKvLkO9nplLSCbZZbqXptiaJ6z/+Y7FY1rodQrGsuKJ+ZT3xwMqp+FGX4WATaqmb
7CiiKJ66QYcxgu4vxh178D4MM4l82gTjhplbCNdmL8HeI55CvGUcjz3KFaHHKHU0UR7Gu55+wlAh
enl7F/8spR9nakKv2+YfASctWvDZCmAnrxw2re4fKTtI3OCJV8FMD4pYq+wGDfHIsGk6vlgQGm+B
AUGKC3QTZ95S+er5+9kLEQWtnicnray6cEMd3DhfFOC1WaQIydVztjZ8KSedMTEFZKfIvicbkiAT
G3YE7Kn6+zribhN3nTpg+aS0ZgCKD+Jxs1ytiy8ZY4pzjHcjLFvUVxkJxxuhqDqvcLq+qPzyXGHS
iCBKNigeXEIN4HHDDiwyvN81WIOGdnMDksFg3eQ7PSEgqjLcXoFJ1wW4uEbMDRx7HVLvPOS42MCY
k89djGMepA2I5KFfhtqCRTRPpfFbm1trceuI0KuZ26qkocboPao+nUD9nfKkZvGio8EtHU0Cmk4M
DyHr/gUrk82CLetZ7MsMegkUi8Or22n2gZkjdw/8+IY7+YI/JUjo+yJ61IKPqOMDZVRmfWwETtq7
QeDlKZx6s3QNrCHs6zvxwAJUS3YUCfffGAPQkcJGNR3BmjwTlOeHKQUuGDJDOPfzxWgJbhBEHKt0
roAXyH/o7EZ1lgw4SwV0M8Fb7m+37C3Tqajt/xOHjyKZM+y2jfoIBpcPBaYPUan/YlXy9Jja9iEq
JG7fhqA9IlDfMMinRQqEtm7vx8OdRTt0DAU4T/3f7wTkHEqcahx4JwFzF8BO3otTDoOZvlsvWXGw
+Fd5bS7D+1FuxDxuaGVrzefi6PhEa25WMijYlcnPtWhZWtUNhGi1X3Wa4jYEzID4DqLOzH/nRtgc
756+knL0I0c4foCzA1Wo53pnX7gN2eRpDridZXWdutsaxS/xMUSrGCTdBZMPOOKxgK2LU89lyzQz
RHr8pzCQ8Iuqi5nx3cBOMbfpjPxNSZ4NCpoG0Aa0UQ/Vm7lXewmDgVcUZg/J9dQSl62ws5daBjLq
saCVwUQeLJdYYUgK2mt8ES9H6BwZhPFHOxbKRl7N7PGsXpqtFhOMmOB1sWfPyKVp+Uw7iI0NaDvy
3b1yhU7cXtV3SvkZIl58rMKulQKkWMZiCZ8kdgsAsR1cUfEiaNTjej431xFWO2mwWOlTGmOg7EX7
pl8hSMlLJCQTJyr8jSqcgStmk/cMDx0B6C/cs3AhI2cat8fa/CkRYjEYXKr5aVSNekUmLEikalc0
qNSi9uCm4IhBepheFvukaDoFSuNy87qr0boaPzkUJXamAtS85704p8xfbUPMfk45grCKjqZAJ0Zw
zmUT6rJTqBjLXtdswsI0jMPFpEZkXrh8fIYjgE2KZCPievUbGkiRf55hUHQbKUCfDrKqQ7SOCoo+
C2Fq5HAEQR25wFZR3m9dxNLQQ8JhkAsVFaM2i7gNfknrf33iZQqf94U7IbR/cA+SjmwjguZf8vpT
mHgx9n/6qNkwUY8ulTgfor9W0HXmFHh00Nz4tzmPTzZ1qUR5BtlMHn5eoTJviyLcAOZtL8n62/28
3S7JhLrGxaZgLbfYaDSSldUGh31dnUq/vfSbNCPRy+l/+cRUwnu1uTo8CaH3Wqt25v9OFCCIYiKI
5NxFJFkOlAkuuNTvkT4GDpVuxqefmqagp9bRFKn2kNN13pEoTQm1Vy0A0mprYXtoXIBVULz630Dn
dTixuzesvmHdjAfW3rBlwl+uT7xESwHlqZzJyDQn/cjAlRRdFFyScS/jPMGh+Seu8eOSKNpFJAVl
eqYps2kpoTf7nH1r+cbuZrNFZFyNJPs7NqKPljWasiinGuT8D3N1eoaGR/ClzFhD4TsTuTNv5NQq
MRPuVXjMemcx8vh/7YXttiXuHz3i5MKCFUZ+9GYdW+6FJ9eODC/YMdDaQT+aGEqtjCW4zoumG8Jb
9AwkDQmLMqMofd2SXMsa7D08kPVnp6+abBaa//YA1QJRvb0CAYzWNdbBwPhzj/Yv9T193SAO1BLV
IObWBAC40cbP3UKGR5WAv8K+w4kP4oIN1elo0DlZg538R3D/iH/zTPOs1SCbTY4YapnujHvUBBcc
y58zj1oRx19p5ryZyE8msVMjf56RrMEeMli9Y6MbO7hIk1w7CVk86oMd02uGU/uZcIkruat3u2fh
/LrU6E2WDUAdmK8mwac0w/kUDUTToWqbQQtMxKfyCj/UWuSw5Hcv5iFWVEBWwoFfMIRPku2sEZiU
s4YEqFl6GlFe5W1/ndpm9/13MkSgdsQvKya4KQOedTqNjU1+s1sj9fEj4jYWN3wEu6evdsxko2Jl
RiQM6XeeEhzenPybXr2fPJwdu/N1Q6ESmPlQUPKhKhwizTUwlupJkd+Fv849uq/UELTTmVJTYzYm
giJXzfPGfJFS7uQsCqTBPEmXg8+w/zmdUhCWHNRwpTl0ax0mSAYTD9QuPmnZOkYLfIxWSf8MbLnB
Gdb1TyNERu6Ck+kqWiIv5CeqTtXSArObgXz2gVhoIEJqff46+Z0Mo5s5MRK+omNTyUNvrf52MNpr
iiOBTrFAHedIwqF9RexsibHEmbUw67qhmi17qaxdJAKlaA2fIw0J/6nlV0dTrJ6elVWdz9hsMSfl
1Y3N0vAjr89r4KHmSBuydH/0oAmf9o8KHy+7enZVp4XWEJvdLPCOhZH9bDiJmWNDDA0t6HBCu6qI
fKuFzin991sxXre66c4L5lyBtslvX9EtXU0mUwEDiUi7l20DT4WaFsTapAVIS2ROha25LCyWqZkB
viEcJarzpZF0JiPoRfho70xA1qFe12vHu6YrgfimaPlpUVuS3HhEC47lT5jSVHf+LGUhPrkcGCsX
3voURM/oMol1RlpLoy9ZVzhYShUwaNgSRacUeJUrQTf2pLp7vT788izu8kocD4hV56i+DpVoeeEn
+SF0z9TY8MYAtW9XLyrbyGV05LDTsV5wXnuCSyA3TPlCpRkTDGpw1PQQXrISIp3+ozTizVWWKwa4
A6+unLjIbDWQY28+bECLZr6fepoaP3qGmeASx4ktWxCUb0PE7bgQhXQjC6oi017cQzGnOpx9n4V8
xPlXvDpNBW0y6UsQQjPwifidw7jAVnNi6iG4mkadG3B7hVFC+JgTiKZ0vquUnTEGzNF2GbnfzI+r
4cd2s0bfq8zWCZGwE3uDFGFc9NeEl0QPQSLs1WA8WzsstmejnyrWIyhtlVGcB5KGp4asSqV9f2dD
n0ojziplpJUJP3hciCaXVg3K0JCk/504wTHAwF7bRyUoW/R9CXfEYId9LKQ6JFOZ1TocRf+HYfSx
yPrbNSRH3lJcuchF2QrFXbRZjP1f3/hBoybPdhXe/IuZBeI+TXOSy4P9gdYywb6gzO0Z3r32RWly
f3GzrkP8s7Zu8ElTcYe4B7Q4uQ7+3OU76vLhSIf2Xm0eadIpvNpxnfAmODJg9h2IrnIuZ+Kh9gTc
mIwmygSxrlKdtYCysx6s/v/KMLOd5G46XUHD8p8p65Vvh4ey7t4Ut2Tf1urAFh2q3F5dbTbrqFzA
Cv7qB+6g5CM6+7KnK78cX6LX6xI9xUhWqmQGcmi8KhnGSQDdLTWGKaNrYOanJuhQMOQ52XezvHtQ
Gd0+nSwEiLa9XwuMXoRcrGBtZUM21bUBCxryInzhymEwr8ujOCM7vJRJRFVlmatWZKuUMxxtb+4d
ZhjKQKs8OSkZCwBRRr9V0SIjWPfksRXjlTWPpGe0kQCLOGvoitdKYqHYix5N9XxXBQ66hB/yHe/Z
XGrsMYbzV27l7bp9UPoCM25KTpInyP9hbiBjfqjkMrZ+e7I8qk3uPsw8EQZbZl5UUJQ8o6yj3UNT
rdELJAwEiCxS5PNLVIMFt59iMe25TFRxYMFqofibBo+UKOlbkDiUplnmeLZ/w7mmIu9x1Jpmm22d
uHjnvvrlGNFn7y93C1fkqhZ6l2aTHwfXtDrGpWA29uPFgca0kA6OtQ72C/DCmdjHV2OXWIRhnO/t
2P22oJmvSg4QBLAtpYHL59+A1GeQYH0asegOW0IhFjFowCaswK+RzerATgIayDnouGtHmTPTYudV
3ecnpgIPPk0xgMn0JkKAPsm6CWtVwrFOJeuleaNagjGM2r6yHSHAE1S60rMnQ1nqwuUOidkH/oXl
GxJd+/jzDkwBtwlux4XtEUtCm62vQCoMFgBPmEKo6EYyJ33KoU75NEyYsGAcX8zbohpoL8fHXmIQ
q1zjJ+H92zXTQJQVUnWwksJSAJ7e+jPMiPDtWdZeBYEa0kBayIVPsWgCaLUyboKOXf45NbnQbUeU
0F9u5Gi9+glVwrxUUi1Rd+j9aIA9QNFULThlEHAudeLi4i6oDf83V5/b9AnJHGLx/6dCHplJoY8v
3H4fj4dnuHJbi9/+stnDoma/8h+bnreTEzySPLPRgcNg9vrsdY+LSmvWEAhV9t4fLKL5u6BuzxeE
UaMWEaN984AzkPlsMvFor4tQwNkBzm6juknUStuhHFDs0YAm+uhcP+EKdZVzMdSoHkh2134DF4dP
OX7CfNpxrypWvXNyXiJnFUVbpEq50GocTs0PcTV6h2dczyO4B5jrKLDtk96bQywI9h7zVF7b50U3
hUNcVfdD5UdbEHla+bbkiVpZifYlX2y3XKs7KJMkAus9gH7lZWYPrupmHq9yZne8w9sGAa81hh6z
2nO5Se+XBnrxTNd25qJz7TQpIeZuglqr4uN7DDGX54mwtQevVhH60Hm101fCyYux7kr1G7oUa7FI
/zdMKHyUd+3zdVcOWpRpykxpBuNKxHyBfXtoCsFniiKWhrBcUExJh5NJRTJvM3fu+KXtziHoa4S8
sHVZIb7FqJfnaghEPexiz8eZIecLMHTenxlwAOLEvR599WFPctpPItFmirBWc1IAMxeRPhgo+m8t
T4G+gtBZRzO0uJQl3RSmD9L3YMkYRdAv8YeAhGIxbM4Oo2Jm/pCo8REJyBH/19Sww3u1O2LJvJxw
TWbrF3rVUI5ZjBOcDoc5rGoOm+rq7oL7MvXkx5AoIGGZGST1x5UqtyZhzx5xm/q008tin0z7BIrT
bdfrldV4iKaXoQfyvnSjI0Yez6K6bvntWl/ta+vqIw/c6CeoGZE95+Fqc+rxBM4OFpN34LtZbJky
ca1fFU00bzG6jiU8STKo9pLZlsPzwh/X+/i9pedQzwzcoPDMbUHeUNtGQjWUhGP2VQ/qSy/mIWM9
0KM6CPWs6nTNT68gmRMQSPW7jfE29Wj6CUJaEVkFD/YtEtb7vZSh3bQpNDTVEskkUAFau1mi0V08
dmF3KTgKMrvdpz5oVXkYs2+X3/KkvI+JlAOsEkHS7N53947mquftLlY2aecAT0X8vXb283v7ZyYm
Va4cIP1TgKB42sCvittNqOg4VTvlcT584Su360FWb/4bM8toFhJ7mDfAj6KiAb0fzM/aK3uhtU+5
fK3DiUIniO1QTuR5j7aZhnnUI8Ht3yBWET4vdPg49Sn+p9rW4bcGbdyZ1MoltaF1GTyE61zT/M/l
FVOaDsk1aCBuAAaW5/SqA6hHWHikcbeoRYJgylS6HXzwKa1K3kAja1B8zQ9xU50Rc06Odmg4z8MH
WDfZg1GJb1pV2BavwehfbEVjaL+SqNDiAexAy7K7FYVhLWAgRiSa7lGB7CeUUbB7YDCrv3XIkVcw
yaBIROQ/DN4+a3mJYovg02aahT+LGxUTWdJ1MuCscTEHPhLxq6q1Vz1k4sAnEG45LHwGqxR75EV6
hFSqo711tc9rmcQmBzB58vJIiMpAr0fXy7HiYlQ+jfn8zmznp3oihFoDzjuRAVdA4byQ+Qx8B8+Z
8bmfPzFGmKneTgPgaj4EreMnPEtqA7msj/BYZuSBvXLN3XuZo0SUxmWPl45H/pjNzrzooaPlIf58
nQEXK2HJr/RR45A3uIKt/SPT0EBaESbI95Y1r8MNlAE6C/utFxup/ihbKXkGEb+CqnFKYsk01AeB
Kc/6riDis+H2gMORLgOhIYf2hD3T0pOZKezH2jztsACa1qIqjjO34MGM7Aj911RWJt5wCNJ0PC7D
J4QEpMl1S2iGCr0fmjY8LiAwd9lc3WClAmECkX5TnZ3OYTNpxmqomcwt4tnjsFPNLjFT5y4lzIFq
v0P5WmqWjxtFwMO2R9XPZG/hKl9KQuR6sqdJz33nkBr3JHc6r75Bhgzx7LWceBsHoc71U1+ebake
4/UnARyPtNe3EgvhjSBatcH1hIEqg0AQHhXe+TzrNEWJOEnqF8QYETgOBaZOMur+JyLSDbiHrEZI
UR8Fmnkkcn9SclsXnv8MpNL9zU/VQSbubH5S/CgOO9Ja11f+Ujpa2PlITv/qR+0/+5D+0OroyWkU
4nPYMwNg2Qs4bVXeesxtGMCyryVVNff3ZGhSRsDpHMoZQszswBWrdk6yYfiOMYAR/j1vZ+oVVPd4
z/8CVj202+kKI96u1w/ayl4iEgtYuqIgOc6TBoxncdng1lbrVMFpAD/VrE2h2kwFXd+e0GQyatec
oPd1U0J3fjekx0AB8lSkghzOX/4mkW3bTV1e5ZfJFIHGi3/PznWsOTFp1j2FYrZ6zzRcM2lU2Ll+
6ZKwy4o6UEnW2sJKIi3ogrimpU22Qx+tIZumpnrngISo4xhCOJRMwqj2uavHN8oJDrz2urXnCjlU
r65X5nKteHlPXGhar+FVz7sHJW9X3ay+hD3/Mw0/P5tQ6wSTGU73J3RtjFPVIjnn9jicrauuRypn
5anjFveTHRwoogaYlGeDbTUfYxagyTwbYKKFD7/5pNWPl44dxZcwKCIOiSww+seFcgKp2IxtL0Y4
yFiGvgJM7EJ32J2tzkjpo+5BrROxhee7kRNrHvjSh+2kaQyvzV1Kqn1fQJV1meAfW87wUM/GUZ0l
kJpTHXZIvtjyXBD+u9SpNA7jSdFEJ/JMD0MIGYv6LchaHm4fvvyhz1iTw4/k5Du4Ny3BSeqeZOzd
+FkQfoGyKKZdHu69eezCNBv0A6nj8RKBg3Cv3tVP+DhpgXkFtfHelM7NpBCCZrcMArXXlTynSk3G
nbiDZc+Cplm5dp7axB3bRQIZm3rnBpbVERCT4hETPLlNbUgE5RbDRbQFiQPyvu/jlLJzhHsKIcPY
0pWEVs/nKzF1Ez+H6ITEJvLM64W728nRlhwOD5ll/60joEM+EU4ayXto3YvlMnIEC8sCvU7WBYH1
CG7em9bbrEOTwWuB/x/+UBauKGTFlUYkcmzbh+egOHtD4KoSN4GkliNIEfogikg0ASedrJqWOKi0
ogchGTXVQJrRurklMY9aQi3HRDNcUbPMbSpIu4CyKv6/p/SThZ3nsd1pESjjmvxIA2V3oxp9QxCw
pM9pKYNqtNwJOugNAjVEcM5pWLQSRACKegr7dSt00cxtzOe7jEpG85fwt6HS9FXe4FV/wcRVU8sx
uD+pRJen5P4zrrHTGv9PevVfAeqHd4NWxGu2XBV3wl0g0co8B1rKnGaIf3gOeLKJwc8t+4MazfEG
Ib0uKBoPfD9pVn64kERVa0sV/NyxTspbWahRMTzmAiVd0mu9fbFxXxy4ODwFTxNvUVlw63Uex9p9
Ug5ij1Tj5aLWsywouhTss8TES+yJW5+pusSrxxTfgzEppZxQ9Yu8rMsU8xkY1eOeDZOdPKEH2EC9
M3eSXhyS+fewb5PaToXbiDtEJ6+0wVhV00OCPJdOm1PXwXT0imLqkpXcMWaE9vulcyiLCoFrdPVG
yDM9ZjTPXizMhAkIao6k0bScWmUvOSgQVfY6kubY9Ubf1mhwUEW1WLhgo0OAM6s70F1hv+Ow0EPo
/9iItxNeTcFR8lyGjU0WyeFqWLVIWzWGqD2z1PQMXHxqeyTIcnpR6lmcTY2UJ6D1VnbViiGcmtow
tYngoav85iPNSWqFhhNhDolDTjbVKQzz3Kxb3zozVuuT0rMFIMCkyymaOxuZVvUcmBDoSjC6pCbj
W4mgOlmOSI/zuuyweJZvWlI/hOJs1kpwNFSST8XTOy+cimpfCKutcfH0HcKU+EzHlvNgZypP+SAR
yhimEsiX7TNcmZxpO6mjldu+PmmWClgXiys6W2RJv/3iurH1XkxYnUWfGp7nhd3X+oZhtcWmqvji
DrfgwCgJUK88rD9UEUcVzPI4G+O57xab/XVAax6anwFQ0UWMT3xBuSiOF+nIkVrVPq7bg6W8G7pR
wssMxEBSkYJiIcTKw6CtQsyT0AQugMkhQgynigkOoBt/R7MNVR2H4eX1oTiVU9zjsmjjHzsZPaMv
pI6m4gnETKB9B740jOyJhGFfmOxzxQkW/C2keOthGq9I10XzVwJTJT7Qu3K17OL0XkoM7SUvE5zy
sIjPGElQCc1G7kFvh5zLC0WKWrrX+oVlSNQ1riuO+aC4BvYi+rDwPdoOcZiexIETnj+PyRqJkotL
ZNW1awhOh+3JtuoIju9aA3IHtc5J6HM5EbrGIeG1ihr5mx59RM5NnDau6Y19sjtgu85vKdE1kWqk
z70qg0MjJGuMl7AIFWl1LBPN9LeHm1yECqx3cL3LC173SCjwayOI2mK46d6RQs9Vc3W3V8/afjI0
9sy9mZdFyCKbJOL+SLV58bWjuhMcaplF3Z7NXjTc7E6gx/6LL8taQqeOlNVvpPXSNSV6cY30MJua
VFjU+fq5perDfrwnQC+Ln1cYA3D/kjrMLrQJJUSNXk/altiD9i8sZ1emqqzaAqvqVQ06CWF+C+i3
rLWDJwen4WEcYRkTjUrGtRTE9THJH6kZ7XfoKxetsgy7c/hMeAGgdKeZaifamLOfECWNPo3U3Yh9
i060TYJNuM8oLsPnU/5ID9AAm9G7JXFWrW5Ud5vOa4tO+KURzVesoaUlaeImWEb9ca9wx7fvE4DI
mqAikmuHdAIGVmjbBsdzxvISOkAjti0q0UIZBUqkwe3eOMS+8xSa0D8vvTwudsNiHT6ZsR/gVi2o
qHKCYZVBLxOdTPPmIPG/nooKtYh8t+tm4YtCFOLSufBjfwsy2oinEJZ1fKmyKwStZvT7Z5orUKJe
kbZeD8dO42cv55LCyKjVHkxS931UQ53sM6SvOR/JNjXG6sT+ljrJMtLUF0lG3zoFWohHDQgK5PIp
nPOBYxWFrNMxg6VAQYAIR1+DxP1ZPJIfu5UuUgBAChtSPXeduAoAp28RHkJzCIeWFRHHhHvPYcSU
289ppz5QAva4D9QCR7cPGdNZUYGM2f23kQB0Y1if469ZIlXpLM/8vY/m1GAuM9H81iHkiRNCNyKd
p6ZOqPq9kHkb+sHpT5sD4UzgpbldHb73qGAtZo2NqAZUgOj0fesWOMQ5eOKALRlO+impJ1K3CLv5
sF+rvTHklPOPR8iNfTQbfGLIFhaS0yHZADyETsCVa4UZUr/aTvMZ59FD/Domvq4OkWl4mvDHRWL4
OgoyWJ4QkvHKl2PsLMkwNoRqclB5NsnOW818G32uDlFQ1UPiOpMoX+/ZuYlI4JMPiJF7pBXolOvO
IdG7EhwVkrY3YAYysfQPdXa+++4hTjCCcSOiclwKmCWmYKvRVd1hMN+/xZAhuI3dbxueCeHO9FXY
D/CIaCgLRSifZNEkXGGvIvTKuaSUtpk/JKm5KA42lHeaSWZqwLq8XVS0r8yNgh+il5sZ/wZITG6b
56fKVMVhrdXC4+0ghX6/0bncElT7Y+b/2bJXCqS48opa16Idm/GHKjS+ED47YDb9bnmCeFKLJuBR
F1MUdbeOflnY1iHwGr9Jtgae/Abt4ZoYZRSnUdp+44OefZJY/C9rm82pcStKEpHDA+N54ftLX1eD
x8kwM8imlvyiY2cV19UpvBmn3C2QRFPDhFBoAuP0HJwhC8+j0/+hjbAz8V7TKWh5zSJ2F1W4ecYa
xhhsSo9tR0jAXqHrOCk4Ll0sblTx75WEaT4VpK60pm3M7WDFZcrPs7zRLjX/tBTtfdSU5YHxIGlh
DXEgc0/x91Frz2LRuwENUCV9tjmp6eZlGJMr7z9xTPWumxM42JNhSlsC8tRJiqnIUEBkl5Ln2Hb9
cy1lOYqTTdGXSbESe2itonQY/Gd35LVCodMtOPj/tPe0GDb40qO/FyEHw01NIlKtPrfZqr6Gv653
6ayfP5SAEyYam3NGeDpl0lccVKmfeNAo/ptZ9R1SlybXdeeQYQm7V8RwKEL2n2OxqADaQWujU4AV
nBpEUpqSg4mBOtpJ+5j/AKTbADwZ7lEfhTs8brAQBZJnNq/GpojYG1TIl3LVlctNu9G1qIROIr/a
9i5a8fh2AMheM+7g6Ojr/m1j1VYfHqt0GDwaS+pjrFR3pCQfkKnhLSDyjLlIGPhsrrpCMzHpmNe2
ZjY4VDkeKq8vcwLESMj0pkzEbDWAKA3eVvSumAr4nuQav0wo4wcdfxpJShut2SCDvT+B0Ngqq6gG
SZDBSKgdaMNSnHRdkpMzDou33xn1H/nLsJa5NQya9bI6Duy6bASP/vIbOsD5qUoasIWrQi+gk63L
38m5wKgEbK9FcefL16qWgu4AUztVkZI0CpcpNi5OflA6YZ0sqEtOPr4CBJXhTWWFP9+7PTzC+PXM
i0Mb+fdKvuZ+86Q5YSjildz1Iawpj1hmc5sHaCiynxo01jXH1RWlwcwbw/MTZfVMzwCKJFjOQIrk
qLKgM35UopU+KmfnfLMeW3RKzpkEEIGofZt++Htcb7MTZY53+HL7R8kQwEakmjulGxOrikZZ1B6n
IRF+jJbjWkneQ4bduUPnXAWBXBKHIk/8HkexA1ASvwUAHgQCzYDPTb0B6aD/jFcIVE4ZN/4ssIpQ
RQpc298wvnmf8mC7A28dILlecEbcHlFnpvNnoQLNTYYkbOJ8y/HnSxELGR67IX46QA9xChknLuP9
dN1cNXHuO2R4z8sb4tBjRGohAl7NLqzPJBRiVFP1NFqg0hQP4FSvC0ke7lnYEHxujiyOjFkadRbb
ceIT1bs9t9sXG/x9+qON65JqRGhF+kp+ymsapt0CO3p4oRxZ2uWPjFx4D017eOZ3waYnrDYsL9rL
d9qykq8g6q3eqdJ9YztNivpBl0D28n2Bw82QgovB9Ss6UQcmBeDOAEZIkgOfZr26JLShs0wQrzfv
hV9iI4XBbZO0qpWCLbhwW3uWVTvPN9r0xYwgaav8o1UA6xbEY+gJeIsJwIrvnyNMuiSDAdlRNfuC
hxuT/AI7dwKaICZV5+84H1el78YK67DGhJ61EU1HN6KoY8NnxMlggTnH8ORUmWeckAWZrDZUwJJp
9e24pBRYNcizKRft47Nn/xB24URwnJRCkH4d8DE6iye+vg2LQUTdrUnWFa57HTCaeeOt0Hh7eAL8
vkyDNvknay6yHyihM0EmZoJwHeKla/H6zjcHG6K8/8Owr3voc1mN0N5l59jA+FPMmtAGQIG7NEK0
3X2jMWD4O2o+TW/C4wiq0yvAq1rU9IIEk5oDsAazJaXeTv56xuO2Od6MnxC+BPvpbIYwelZDfyYd
OgtDs0r7AqG3DgctPTXUj2TZBoe2U/uCnZGhZQj8nhxp0oWjIRXAkrzOfzSLoOR207IO84kF/AKV
uZQFL4rDk/rVXRhgQKRGeYIRVLoI6YFkCHFcx6hgxnAa19xCut+KeNrKRto4lWMMUv5if4qZ2SDg
b+QxCI9rCQSOjLJGDlkey5ZUKPqIoTrk/oNekONhyPUUUmXtjt18wgfC6OtMKyTXMe3KQwQa+1lq
OebKElivSzfyT9YtVR3y44d6NtOZHcOKi7jWxFPOiTTbXIoZPEXlDDHTYZ9WZk83cLGB+2IDrBzA
Xhf620LE73RHfmspdHnUn6cTZs8HE5H110bjWqK3zz5hvMBpM1bE6eh3bDanLdk+puZbvzGr4maT
dZOEL3cYE3pqUyJXy8hIHfjsNF7HlzcioAdz/juVu0z4eDaX0f+QBtH8pUWvpJTx+vkRtYbFBmv+
Q5TR68jlv3WFdXmqDfh/ZU+qeHCtEtVbPdmVrOfMpdmO8dTqfWEh6BhHNqot6ez4UntDtm8UAUox
GVAVDly7QZfKs/OKmZ7g03T/L77aEXrFlg9H39BiHd9WTyz59zPg0bxTts52vVR5JhNHMWCppYRF
7hRuxLsZl6q9Y4IKKB7ipQPeSnvWMQz2R3g4j4AI7ecBtCvAGT0lVX+gJF7yMM3ZpGyLUE+GI7yG
XdRFKMrWOCmCG+IvR9rhRVTvwsA7zVmnFWJ3cXYefcfEkh6CYvgdKfbYLw7vwDo7+C1hclQVEPnb
oUeGvlnifWUB++P3oplF3lRTs4fAQBtJXgg/pEeIZgfz46bStkafDD6Y/oXWiSgvHY4ovj7LWK6R
mpos1Sm4u8F4TyvaO+XSVpfGMN86w/EYBOcDUqGMIZ9lxF1M7p36PxeGCX5dqnzT4QvpwncfytoL
ec11kNtzg891of4Scw1Dq1lI5u+G9WTcXn6MHwfW60LITL3aPgKuyGvsKDRXIYnwe02uXRJ+omzd
2Fb1j4uGDFaE29ruaz/t0aCBzhG42t6DK0JNXVrrqj3gj0nLzRwdNPDP1aeGK82zh085scrvLvIp
Uaz+CwbGzMZmE4kM10TRwuVGIT0rkwzD82wIk+s28GyyBDF0HfSk676P/AcvDNTc4NgP5iI3i9Je
dKeEX8+/IDcWqTwy6jaEiV5Y5mpj/o0sB6S9z0ocCRRF7p+HY+MW2xJPbBgZ6LB5SjWwJanm/suW
u03pg2MT6sb2KB8OlyVi/JiQFnC9xUsqdEDMU4wZifNg/rIQLMFOtpYZ/P4IcZs7bY3UcmtnUbZn
YU/T5m6DS4TCtaUZm6k+1FkAHpygbFHzP0z4QcyCrkPufU3wXW3K+VDjB+x5ehbUdpl/OgHgO5sG
+knMs0t1fjcTG99IqcQR54XCh4aRc8TeiesGXIwOJUrUsOCrcKDNxnXI3SCj6YARpMaxNDG7Frxx
N5pm46SoE6R5M9nuDJ4bd/b5NjDSfdQ+zObZMAyFCOO4ha5eBHDP6JXe8ilXhu9vwB7tpl6rHms5
QLP7qcLxGubJrOptdxb5KFisbkDsaFMlj8BXmY7TWiySXXwY0+qc2RW0C4/QIz4/klkMK1oeHMKQ
AHDBb/94eJIg9eSQE/6o77JAIXBralfNJB5AZ3zmFo+yBlIDfIj5vX2C6NsXityDWYxr55h/gM1Q
1J4o909xgyy2svGGd6XfdW2i4LkadZwK7oVQeyHx9MGrXXytczh0e3Y76V+K8XQQ8COIoK8mYqag
hhGvTUv0wdu0qT7KPSzUte4cEqQieLI+hadW3BoRDtsenGsuJCa3klyJ/sVu4k35oGuVNvgYmMlh
24gcddZtlvvw/UGyCH2LMmxJnOsthsB0I+2QX1B4tme7V2+nYVWSviQhrwVniUTpMNq54GI8yOBL
V29lBW5NRW1sj4kZkay3QnyZBYdTdh2h3rKWD+McN30DOnXFxiuqOiIG2NaV0qBbQwrQFVSUYqeR
0FL8XxJ9RsE/CpTgGvCOd/aK2GCGLVhBSwltmT5m4ICHsHJLL37bQvBoJxPwNRFM5ABuXGl6qADD
YbCqF2RvZABszFLJGNI//yBiTe1SEupvAMpQP43D+RbYVE2TOLgzoj+IDBkv9pXa3YIG3iIQEh3O
Mequ7GfNLBkodLZLP5f4EyoLVM04YCxCLzNDIPe4YkL7PoGtafHHw0h6jTdKrlx3znhWWJdFk8tf
28uYoNbYyawtWa6r6m++aCeVXDeQyNQRz81U7cSdnOdIZnvL+JM7IKICKeKwToPE5U6m/ZOvMD+3
qqEfmETacz7dIKq6NpuMAeg+gbmI/FJDlV6pCl5enrCecv3Vqis+0WusRFNHDM602PgDyrO5zT5C
5AipnBPsi1Z132lssqSJMv4oMzCY7fVJxuytJ5caNcLqK/eg5KuzxtoiB/BGmFTiL31kC7hlEu4E
G98q6UqrO/3BYiMkNcWWXBKHiA8BVL1gJ5CV/HYt6wVTVIDqQJTysszexuOlE5BNFVEcfGSoMXCz
WqQJLDJwC+1NISYu/5oFIISTVicZqfDCkoUDvAnBZGHNUZe9n7qbjfQcuoX36OWs3Clc81Csw6eM
ia1hPnpXvzaN/7aymNKCMiChkd/a1gnxaF4xpm2DZEz9QoXW7KaFYgTsSyNb11OsmYlB7y6KEgBo
zVHwN56v+dHwXugPqPiqFPHC5tlkH0yrClxWsPh5pW2x4KfEOKVBdh78l+WT94yzCBzPmeu6rjuY
ERdUWImAj5NAFizgG4mtATe34dUYiZ/t0bR4Uc5oM7yjgsfR0i57eM7k5VbCT7jq+RWVt970aaoi
PQUfqR4ZBZMo8FifRDXqktVxTzl0ubWuglfUDvHwOSX1CKIA5GBaepj0OV2FWr7Z+OQd6BhZmYT+
vnfNT7x2IdDEZfj6Tqx/gPwsMPEhfFAR0HNebAdqAwg/GkuBHAtEO1KB8nG+j7pbdR7sgCK8Rf0F
NIRFe2IbfUeXEuYr8NjWSLGbSONiDuS5ZFNrgzYf1wY7mjIekjQOIqMOyHFeGPsoPcROJa0PWL7R
wWG6JtKg5edFeEu9OcDUc9TMjO6LAuL7hAUG81fIl45YA8p7pONCgjow2oymGZYpfydVJCbFIJGV
PbSla8jpbFz/+LX/M+euoNOa4fAI3K3WtOMJXEntrhKdbPy93a2lx8+VVjO5f0zb5cZqVB6uWVaP
AkXvOdM6BLJpyojfobamDQpL5W6R/9mx/CcSM/H/dtDBuKA8dVghpyypbtm+biH0bIvD21GdcdEg
RwmaUQHVoXgTIJJNlRWmTGsrGtWxlIwD9gjvPWhFCYnzGvuA6A4JQ+pesdBuekoC0UYi8BmxKIGy
eiZd6K+ksYEWpw+6EyMmdH1SwDR5+Jt7KthzqhpW9RwIiZlpSizJBtrxmiZQniN6YRcjZGKCqqru
trxo1LDArWN5jRKM1nMO6FnR3ScEJ17Q4ejO2YzADMTUV1NezZbFUxH1H6GUTgyDesyIRdmFVRzc
7paLwjKagM7vSlC6NFjQgkzyCbnh1wtMm1+PIeqcfz5N6ofI/oHY0PntjHyyE5gtxIva3xlK5mhg
Yfc1fewJ0HfnqK4+4Rs1Q7IaFrBVifRbbx5bf7WHTGqRveAVVsVYJ+y6XqJyBxv6DFGOZG7T4wZV
Qmdb6fnCHtg+FNiXwjzkkd2qjQdamwoze7O7VSVLjWmp781RaUrakeVe7V+9fSXmskeHDgJt5Z7o
9NGVLSdAwj95jS/fOJJVmJ9+3P7MiQm+4dzuGMhAOUm7rOS2fdri+cql9a2W0R86RGh2m81uYomg
Vm1ErCKj9fBUwXcA2u0UvJmgiNQkrmxDXWSTYD4gJIUYV7RUk3sfDnuaVprLyXOUjKqll/MSvNeD
t5ysTgbOw0xCQW0Ed5W1xaoWZNzvVT89g/uuwtI0eNC1uAB22pqogHzlPe6d8JJUiICAt2gBo55j
oTQMBIu6iMsezUF9m0fesY8MiTGtwJ3mlt/MMw8UnA0fb7eTdnAjZqdDTADVWn6T7K139/hpflwI
Bhvj+RYPSw4pDkCjGhVtgbCVVLIGPomaE9gax+RWZsoC8982dWywitPM/AIqcjwljOedA5w3W9xu
ygryDvcxE5WdUiPcUYmD28/X4M0E1Odo/W/RB4PY5JPDPSkklKq4Zijt/SO0HS0vVRdtF5O2IbY1
4lBlAR4BFrDRhohY8UKfygbmVEyJ9rSBVbrLO4l9Q//9pLuXfPIJkwvNIzPKCns4zUrDcU7/r225
88q78Jj4T4Cja7CdP1VuXS26q0YNwvMDcWF9DRuPjlpSBG7PmtRCoaFJG+vL269uZTA/01K/Mr6e
0lUuaSBaolZmGrvgEpK2zpojoST1U6r1QOHkNV3lJxjDCEeWuHwKfN/+iQqMfRpJFMg/ueeNqdRt
4+QytCUmqjfVDEurv1yFmTdOISk3GO/fdqe7PRWmJfo/7kP45NJ7vLDcAiaGtH+Qx+kKN/ktiU5V
s7udSmPvlr/d36e1j5MMqUu44DL9wao9K//7LpCD15B6aI59ybjSY7YxamSYEPl/Y4mOb/fZUFP5
+qIjme5A9qLkGPpy7mY04+3X1gKgbsCdXQ2IOBHjS2AYmj8eaAmsiersdWkci44JQdeALb5kVZ38
jKk1j2IEnWMjB1v9iqEY8fiZpZ3pfgmJQmAeR66bUF3Jk5oaTU5XfitX/sY2fCQenVX8qf/nwRFb
g2sFihm2Wnqs/d3nit4hUct0NTscwNqqL8HatQ66TunZyl/KYKTCm0EWwGL6LePMvKLpekADhGgr
GW7cA7Uac+PyQW2O1DL+ZWaZU+vKpnh+ZR0kUUDJEqpMPM6xJtTitm3U+0et+j2n7dp5/j3UVRoY
AntIJByVVMT9ryqECl7l3cdJjlXyVMo8UgnsAfepav16co2xzgvEilrbk12CCTxSRCxiLyyWHBqQ
dZXGHRBYZIp/tZS+aFRD7ULRRaf0R9qqlwqgSxtjm3P82XFcscJA9Qj7abWd64VfgE4qCEMch/02
vJCl9G+Nhk/z3Uxa8CtIlQdmeHrPOjddbhAfeoA9rHM8jxcev9lGp6rSLWH7YBQJ7bOv6YWZIdFe
YAm2pixKgsjp/TM3C7zXnvsWxe13Rjo6KLS733eMvwSpyQRqbcAW8vdzuhoOcd6XvWdRo8wSfNqw
KmeaPZCksOQUhuPz7TnYadTJmjpd7MX6k7QS72XVB23So+ph9Uf5XqrcMnrgVDO0KjfCRqeaXiep
cysTR3DKOXJFqP11M5vKP+wtM1DHZqqeblzVu5mxJxAjSIaoz9Jv0vQiDVZjgy8ukQAKrEMko/73
JqW//NcfUx9Wa69urBO10ruO9MC9GHyKmaTRvhR2zhxFiEdpHQITQkOz1TJqPIjOlIqIqVGW5MlJ
/Pw2yi5VCVzoHaqmml6b4MADSOJJgL0oqm451l5OizZxQVlYfmpQLu5AjdWO8fvbfLdiGCFhuQGg
pCx7xn/7IHx+2hvCdQXPplDV98PY5X6cZDG6ullys+7efkK0/TnT9nSweH9isYVFYsbk7u1mBFMR
Mki2lmFdxehBY8+UwucKRVOoLcF6GNnedtuTBk2sxQL8a6pAK76npFf1MtnHBDrwsq/QsDAs1N3D
BIlp1Me8o5QmeN+IMABd8r12npusdJyepJWb8y1eQ73tc2Qphu4XAJwztLl5pZMUTYsmX07RYrcE
4LXaE7x3/xEvoFG8s2EURPAp8B6tuKqW3KsWOt56ozpkrC45IYRYy78XPDASQFRmh7mI8JO30hc+
DLIVB4c46xf86hS0jFOtFKtjwmWGDvzYDceFGiEMKIa6qXJizuffzzTSGA3ttbfifAdyFNCqfdGr
P0/2Ko74w7Uj6LEKeaRA7UZ588C6OcrWdxClJ+24cqex1oQHnfgIkxmTr9Wwd2XOAXyQn3G+j9m2
VKmSykIk8DfI3vMs2N09I1APophsLCPurxjio1JXWrVl9T08lrUJCB62zSvLxYbqhQmM/BiPNkeT
4bEW+EWkwDIWTjzIz1jxeUbCRm/3ZAiDYoQmdF0fcM1Jh5HDeC81Ymbe+ZOXidbqqTvRL2MkQYHG
ambRVEoNTjDScTxdKbzGFJwJSmc0VJUthp1/aABnFfrY9ZijgAuW9OwKlrdhGMS/mbifIk2xzxeB
6UkeIgUaafu8a8IJWGCXDL3qkfjWS4oNuF8g+mmQIMRbkH7Oz7wY9CEuyts7tlWHG8Yr89bqRrN1
KZDTZmCsaHMbiO1fN8ZTA6h/zurC5m06EgFRIfDO566QUyEEJ1UhbfwhBOveyhbGTQVgSDqYx5HS
TqKl5hK8Sv+PZqIDLyj/kaXYmwYaIA6hCTgei3UDCllHb3b7FM20V45mQ5u1wzM+K33hWXqo7vMQ
qeq72f26r3UL9RLCFfBd1AQxEWkoR3Z3VzMrw8EOpKDplLaCTtG232h+4hGBI3Wni6mJcxosAnsf
losAb0zsxYDGYNiKLjZAJM0ET5KRDypbBb37RJFm5ke1m/ZIzgiBJSG60g/yvtDof/21nJ3iJFF7
e6oNKBPGkYpI7O3MQ1sJhrE6D7XD6uOr+waeK66xZqwgzEZPk/8qOg5h+93fKiqgHT0VrpFlrRFl
mAuV41d0mP+hGmpuibeHmedKjcCPoAVmCluRC7D/fmYEjf7A8myrOhLqL2H4ox2SgkJWe4quQC/c
jrWlnV7opfYIJrqJUo/mSJs4VtrFL3Cf1aFFq0Og8wMfJBZSqW7NaXcvkShZDKDRlM6LxSZv/Eb0
7rXh6/h3BfH5q/7of0rTVL1tTzAtaQz/T+fHRKF4/lnls1TGz1Ds1saRi+tdTmA8JsrtYMK3IEpw
ZT7jlVZF9CffTi386ogFx82JTtShYD6+EQCuN2JJGjKuHCPrYE4B9TUWwcTigUBoT7eEut5e5cSp
QRybHYMIlVNxQyxIfzOCtbGwl81rZYhbkJP5ATe2H/5ObSLLTdSg8TwYSAme4qzU9PEzSVKP3a/g
h4VKqboSDWueWLC6NJSu14vmWNnN7Qiv9tW4BG94oZOvoypAPvSRivTVyvfSSPOcZiD+A5hl+oh4
bl6ov9u6HrSQ1gIE7asys6pP0BHtajQMnTiKsDTLnP1xym6JaSxu5WZvq61GclX90jVW7x1Sa4oN
mzZ4M3+INbK4XMdaxkFABg2Xt6hY5l+shPZpvYmj3/bePewwCGIFor/KcZN/CUGBglOYis9ARGXQ
mZJ0dz6knlVJpnPOI8XRoaR/x4UhxHRWcC1KLQFzAx2yH/VbGQdvbCNjzK5perYlxqXBXxoPt9wg
TkdIn+iIme6hiyy14lxUhmVoj5WeiCbGT6QKjVfiA+qLAhYTPY6S8TLhiDTlbENU3XowgmUyN+qP
FFLf1gXYXYKEhC7BC/6MZPFhbLyHaucZGSfT4/UnLwC9Tl3b0s2NASVz8Y2/R87wWD5t3CLHEuIA
6ORaYZohypwsv4hM/mAKHxUZIBc7QBaTArD/lurHpE6/8nJ8a8Q5llS/4syQgYA8S2cFWHzxcAnT
bdHIJyH/96SdYECnhEf9A5ouuBwjMCKkCOlw10cIq1brzwW0kAfTWl6Y1TfnAgrRNcs+OVj7oP2/
/zZIo2/nxtE1EUPYJRQeIIhn9ihx8nK7gaT2USjZUwr0JRgaFTXaH4EihkgfuapzrIBo/k8mKEc7
r3W/dcNprfd9UhTs0tMrO0q6UHyuBhJ8XSLdaQdFrX78+/QpMBmUiKXLtXcxcDiDSp/WnLCpemEg
2VYpJ/LYmudBvBSXda74Jf+LICWazxJXdkEEOdG8GHp74KfPHdFuvphNBDVMqAZMdj7dqJCaeKI4
96YZlq2um1Qbg8WilQP9Lcm1QV8FW3ugJcPWKNzgtxQjPc+SrlLDplElREMxrrybvAHEGARqzwbg
ovqh3vWHjGKhMGaeJovR/gbzm7FVJsJqP954pD582VWcQJ+C3HK89Go6UpT6COHv5NKy+lhv7NTi
16o/sfR53fjeWfmcM1jIoh9JHhgTA09aHN4XtRmqN6tiKC8w9JVu9pyav8S9eItJrF8SlRgr/P+w
zY4ULg7qQxoGr1tewxUk4AZxbMUXsb0I6BhOz0TFKiYl1Lv6lH4IaKk7lcBb8FPdtciiRIkNpvu8
1BAgA4Bq6TQ1lruD/ii/NIsRW3vrmywxe5eB8iXgtritabAGEtkfsRQS1EdGuatHMGPTJKAMKq+0
2XA+YKQiMNpCBWgowAxVBrI9lSSUn1KLQ6UNE+6LCbwHcy0sK656Z6JNdbrkWVZjf1miiVGMd1St
SnmabdeuNToX/bJkTS51g5KxR2fxAJwvpzrxfuj0bOoQyLvFqO9STtDCwaDzBVq7WnhuRpi8bjhE
PQ46xyuog/RLOO36BKo6J7n997TafMMDmhJLBCMfjrlF98kTxjg7V0c8XO9IsjtVuE+eqOukzr7A
TW+L8h3JCUlhPM7EshPQugrU7N/CBQUOuuwWpYnbgLVgg/MDHy4ePnN+DgdPrmGVIivYxjt7hjAn
XrHLRCYCiFXlc/6TTyQGRmGgGpiiriC1RHKZqzlzTH1WdE7XSvovhfZGE36L6xb5qsgG9+yYEeDc
nlSDLlxkvvpU7k5gFFTTVPjGPZHeTnt34uEB43Si7kDpifuQgkVEnNzk4kb3/+oLPbA0Leko5nM5
IOYpONEZmDe8eeZWf4VafZWQYuei3Llp490Z3P9ZzkUUQFOfD+I6EI/UBfAuiS7IlGaEiocYEwtG
t5/+s0WnFEVUiGSxWp6kHZNXKedDmNz2zH8eTj2GAx7qrhn9sjY9Ohub27cYBIxEtKoMdrtERZpI
qDliGdamCYv/8h2XhG7p+UsQ8MGFPjNFUOexqO/gc72Rav0htgS70GPeleXPu+laMtMoO/Fwikcx
jWM3Yx6CFeb9yfiSyRNWhor9I8mPRy0g99t8Rhf4fM2zKWuuKj79B0oIQjdpIbeg3c5x6WXIS1wM
FF0CvQekwDh4W12NVTNCVRwA6u8rA4g4MBp9hefTqA95VewJiN0U5fnoctj0h1kHaFA4CEnYYe4w
AUcL7qiH+NK/yEds7i1mRiP7NnfO8Ct7hD8dTdCzXQ+nxzDdAHizCf3ousEdi9wkSmPQY9UeGBCL
kRmMefYfR5Q4di7i5xfqlE3ZZdvT/eeIj89nYCiR3SccrJ0hCVTcbtSl23yVFWqQnWUaO/thzfDb
+7Btjs8/sHuI40rSlmiXr9CspUMBz0c30D2n7n1uJZFgbjhnY4r4f6PPZ+zsFj8XLd0ONUBlWP9G
jG8Raof5hveJ1TzPb28XqPTz5ou5OlDXyfSPNsqct26xWDvYDG/H6ZEntzJu2+7+b5q/J6x1T/am
rlcK56aBWyhH7TmkfWsG45rCNABNwsIaIcl0rO8JGUM/c5ZSHlPNKO3g+MHnQIxSVRD/pegVR7oN
7er72AtMNlu0j16j5WUydLFwASctYQKSGzB9FFOCUB4scJVU7iTqaAM0i3UEG/sraE5nYfMt5jCD
S5Bk4Y13knmS1dHrOrGAphzyhzpHIcj6z/IpcrBEJ1QjBQls/FiQ/1MtXHryn6U2ONn6K2kshUjp
buvUNSrtisuq4JyCpyC/krV7haYNncRcPgljHo70D4PUxl3ROx+prFGTfn8DgAjJMHkbVIOceOUD
dfhtLt2w+7qOEbRgcBEPNPjbQA4duA7LOj8qHZv+gjXsphnslsweGyeiah1VTmLr5STNqtoUX/Yl
J1MC+lw92uEc/HgN4YikpxPy8f3EOjCHFPeoDbsAfomj8ovrco+FE8kG4sgx4j1mU4YTXI6/f7E1
IKpGDmDt83hfkqlI74fUT2sH6m0ZT+aBJPy4xuDtaaSuqTm/wd4+eVDFrBTX23m8VcT8dOsAYXnx
ELx5TjJY6JLo9C94N6vLO5IGI+f817nj/6FrAymcWaBJKMLVtj/BFgtg0UtazgTCzq7qmt9lQ/HY
no73H5SIUb8pAoOJairDzN7N1RP7Cgh1VbKA+ddWARuhqSXw198CHWbyUBfShdtMsy1QsFyAgdZ6
ph7cX89wrUSkvZ9A5obnMnlzxNf/9wYtJblCxWD3elLTK8Tc9tpSA/2Vob1wXiuJ78Y6R2KNuOLC
9wfgtPhrHC+esHGyAUgUAJcqv/D5v4r+4bEsLKUVWHvXmNCa9oKGId0dwzpH7ddgPSs+aZcuTD/D
/Clko9Yoon1NBgIP+a5SgJUNoKheOQGlXI9mNr8x5BffMZDbhBCWhzou9Mws9uzDqzBDWMPkwqQZ
nti09ONNvkHyQ52dGDXKijkhx64vlyuBCRz62Q6EQv+vr/2mq91n+2co5eo1HQhPeKAHLlpo8jus
gzQsZQcdxuV1e7UWBrikfOoiRk8sodnCcEJW0NYHXgdK/tZUrT80YAnESQVDuktMZiIzpE75shpT
4mfbpbKpNixfWEyaVR1GTuxr22mbVeTxCX7sGNJxnqmEUYEO/hqaGVDlG4om5lEVQtomfYqdgB5w
C28ZJcRFTMVnGYbC7b6pd1hJfvv0a5p6W+6yG+6TH+w9YllTqYR90aJuSqhEQkMhmKY2s+ZMNDIt
t9ehFmd9VyLRcYsQTpmeQVhNfTxbSwJdbz/bJwpos8hgauuxNVK3n6AIgHdNAXZVDuJEwViPYeOY
RSexOCUcA9WiFCbYuuZkNwfTCzgQT/p2nbj7Pn9vO9+NMjZhS/GtE0n+YcvONAE+rYbCDhur9tek
Xim/iNxYFYuZemcre2Oobqr00l2Y3/j/48qGijHOueW7xBAAQ93cZVlXJMNyrzDeH29TNd8Hro06
li1ZYOrWastI9zn5NLBaFWJL9zhrf8b2JkBb28OtVnBEbJva7H4rHU5Po4kjHpSTJ5T/QOq9sVny
cBxRI7O1KWGvvUrgUb43+RofUuzJilZ2sOiU4ag6ZJecTukutBwb+KdLsyl6Su+ngimqy3L0+3Vt
3BwmLxB0wdKPOBZy0hYzsfITR//V6Vb3z8I+nuNWTjWXy1Dg8UU7NXH6mTc0G7TWoqhoOUAyLq8A
PL9yLh6os11KqV7R7CXR/9ArrDLwgKN/aIWVmUohaDuZqWCIzskmHOIjFEQzqIGa0Pm7bGcFFftH
KAzXGG6fCSwsTWlNuLYaiiKt7cgJcsigoGv+W/CbaSAnjkq7bMqG9w78sGm7hEtGRy+TklDrWac1
Tny+g2WuhXqHmrK720WSyFxVNHp1QhKTq0Wcg/pPT9hIDYD7jiF19EaZ3TKBQpG7ceoFgMk05Qz2
FEvPx+l1xuD584Hze9TRqf5orTcrli7WddvE98fn3jYd099grgDWyiuzXWpTrg+5WFhbPpWGin/c
pPTy3kbWXOQ3VyNoQGmNXKL1hUZbdRY4+oPpk+caZ9WFfnMIffEVlWoFsFhu8jmj14m1/fNdKhJw
is1NFWgRGD9wImRo70VDnqIwXIE5d3tflRl35uxcWWlCOGLk2DqBWtNIChIK/oQMfzn2bKIt3Y3A
jEl5FacrJoWxh2b60kKiwHB0FNF85zD1Nw+V8DjOKz48HTi6jTTZduXvezgWaGzxzPlCSxgin9Yi
if5bcZzkcUQtGATkvnW9mLwAakHxaJ4LGQxd0K+S54sCTm1THrRMBlkU4EelMXjVEL3zdkyWOWrs
yB6FlIg3SZqRY3QKH55ouSXInEt4mkvVg9oevL/Ce7lweQKzQ52Mcp2acV/03Wk9gX0kDKa7gp3F
tCZDM2UupwD7+fHShE8zyD7qRZOmShip35ujmiFbv4Yh85gNYKf3TG4ERoB/VKhCtnhI50WOOCP/
IF0AV2/m74e7cC9N2ncNS431YcpTouFF8biVZhAzrXNDOqoRspJeF2L7s+bRMg2P2SjnKnXMTW6P
RBYL2ESiOZSQvjUMfMZ1cf+oGs1pnSQNHT2RUipXEBuDYH6tVbqyE5T5WRwYEMh4CxROMmCX1JOB
ik/O+EvhWhKKgkLmowskTVUAKjg6RQyDz39iTSVROHpl5GaQ1trWtqqS2sP5dZRVZiEU0zkZm5w6
kDszL9V7lQnpLD156M/qF8wnIYnzNFOYXm06kneUimAgbdlWWFvbYQ5JJdCYxY8PME+1Cjc85Ri/
wYF1bkcqn3ajuMMnmKQVt9G8fITlQy7fCkhFOGkByuO0/Z4eySfrZEvZZPA1RoDL2lY50fN0y7Xr
XjzqA5uCfWruaAWiQ2TIDwBfCXYefk2JynM5mdpn1ndjqAqezdfodZgmUK+CMI7WoMayLHKF5S04
h8mROxc+c10JrJM1nc8UV0BO+77GmMkcvMxDwEC/QBxnBVyPQ/6hU8hNPs+g1q44N3B++TQ5qshT
3NMtPbpYdT3+K5xNcu+0SubK8YI4ScG+8xnjC8ZzD06W9WO3n9kNrWkhnklOH58GPN2QQjKUY8/U
lH46aqvB36LCGAng7nZzZE4qDEg/rqtCXzs7YFR22OXtq5MFWYgP8pNezaw/IjVpnQ8gahQ3iZrs
J28rDe/Af+Bbufr4PuWSIPR4Xuu1ESxOFrXWfs5R4UdgYXoaWIz8xbASsFReH8fIvlOqKvMAMJhj
BYjlvS4znGUZYKGPJyd1k1ULKIiuHmdfxx3FPPBeyT7thHD4mZwki3HIrbJMNsbpsMY5ScnWcb1Z
lA7WVPuXzbE3QfSzbjd57Bm2O9Fobv4XZ3ZkQ7+AjYf+tJPMFaGtLskxllBQbCuliOd1sqOqLCDY
eyffJsIpjb95n9UXMUZeS1qC11vKdQA7cUDM/N15yEMKCaYC1Evn7s9nOD5fSIWwBLg+tNYvpvSG
PRXlaw2SWXl3uYIGdjTamPCZ6Q0bLesvZMEnnNOr8xW8gvGDHHPtnjgwFzpbJnhd9Ubb0CD10ap+
M/EFzSDdcpUM/CCQXRjdq3IhVlDHcRn9waV3NVXIwVbNDE6KLHI31L3yG726dH48BAI5x/3cAT4H
NaPXK5R8dSNG9GC7K+kSBG0DLkxbergZinrec2QerCLAHLRu+r3H4cvArmJT6r9qCUJu99Dce2E5
DWoL27OJXREc4Fw/bLInATF4eLE3tX8KjG6rh/Ry/BiPYN+26+8qAyIV4L3eTjynkgZpGuQtlXni
qoLrscqX2gGwbFPexnW1RkDowu4G4cD1Xa2rKUB/uNCMTCVKe/MnGjcdzcRSPmDTn7ixgPQK2PxC
ZzIBm1jHZz99Bc2cmOgg2DDAYStS+TpxYba3h59IRp6+FXHGhjThBTygyVTFepnBHpbAxnkm2lkS
COGGFcsVJQPa3jI4Gjq+ZCp5FtC9LrIDhYfjwxsn+c5TjhVLxg4mIKXflc16dGkOLyKJsRkA1loD
hr7oCw5onL5jN+4EGNvx57T6t9gVTEfH0pkQB7ZTEj9FbyRn7YICL2H4AVjkSZxLOLc/4ogXZZbk
8ECxp6k88T8Zx9NxbNeShUqLAB70TqIpY2BaSCXIXGEPnSN9xDQtr12LOJOXZsdQR+8v8GWS63po
dHbWr/B9WswpStt//APUA/zl0wgZXn1uwnXg7BxuginMUyjHpMmu+PBd0rKqshABlUgkm0JHY+Xr
RedhXNZF7KTRPnt40YLH/6Z1tLyFaEyk/x6baG7UigWhSFdaXtHZDq1RS8Zm3kMaSVy4W7rAbZFl
ujmSvtV6eXX5UVIJ+kOvUYZXWh3QsnfWVlNUPbVXpNfxoNwbGrGWwZAKIqV3eyeZDSKNGJMN3lWG
fEREtJ9STpPWI3RUl0MreDkO8eB9mukPlEwlU690TsQfyi7sWpqeiuBp5Due/tIgsrC+l6Ydu53p
FStPyygcdE2agKDIAiDvu0CtMM4W1MELwBtEJo3O58mLz3wP+L4i5bSrpJ1/icOB0jvV7N+4c5+H
+qSJYTd1QT6g3GWoShbSMa1QUpqPLxEI7aR7OZZhd+eypfEUjEIAYCNMbYfGyhGuZ+XbAPQugKs2
6Nq0nLz7Z2SI6B3g90oU+p/4WqYS3GnvB8LnxFOXgMqp/7U+9EYRp9Mzm8rf/20ykXq04w+cwl4f
XfEKi4s7KDZop5jyIwaQNpCN57UVpFT3CLm2qLZwIzTahNOgGzEGpjB1mcGkJ1n82uv3SLNShx2q
t9KFEwpS61qrAqtPLcMRTv/EhhN4adu/Nu5mLN61jCcAC4lnF2R+SWWXJSOBeT2hFRt+LxSuqJtt
YSLspt5mBKJeKReEH6ggKQYZhVqRappaDLZWO5wung0LClEDdgXgmvC/ozZ2eUU3xshplZ2ZHbCV
8Vg6fNZBjDVxbmRBRNWxO+28RVdCt4Y6H1QwSpjxfUdLgrYLBhPY+yfegnDlGrtA8fyGV2uinA+Y
FVMMnIZvwCUlA1oG0/g/oNsvS2BMa5WPcKCjfNgXRNU3xtyNd1OgnUtwMYf/Hc1YtQDrS24vdylw
nsu0FZHc4tZU5R2+aADDCTEicU3tJdZPetkLklnf3MbyzHDIfftn7KDGwndIMmDcxmoCsHS0R7x1
iXj9jKXSo+XtFmDE2F05a1MYqbW+bmAu5pZI62ZMHUQD5BpFLqUgZuvxQd5cJn0ooLYVkJvEWZU1
q0qRkF4Q5feCk/KOlm1a4oxCNrXD3Vmdgpxi2Axg9O+nQ+hQN6r5te/kj4FNDzn4NOhZvhyXcBBp
HhjoHZPMTmiLxuStmie/FgZxJtDDrD3YqkU9vTp3eped6saNLEFfvpBclIbBmyW6FMfs+NgYpo9s
HQK2LE2YitseLRI7e51Yn6GqUoQHEoBZtaWgQ3FmEpkMRUB0+Rg13wkFRyLzxkF0EnuQr2vPZMpc
S8ewueJIsRpZdeYaQ9BWBxe/fAnoEWr+tWWSSQsovUAi9VmZqaRG1FCmss6KJXQn7n71XwPO23Qm
xypZbg3h2Q5aOdhOkkqtAbqdFpKarzXjw4ey5OKRBlE2t5F6GIbtyYWYq4W5e8Q2JbdsEX6WRcJS
GO8RUpCyFr/oLP320QELbpNfDv67AxITel+vCvoQWCLfHgffQ63eL7ZWhrCUVhOGSgQPIWa4IAbI
ijXrqIM4zhv/Id7XL7xk+oOuEo494nHD1JYkOMjcOFtf2kQ7TEkKxaHHP1d0tksh4/ehdNzJeBYt
zkaTDaihnPxKsiRgV0SqJZmcSZ9VVnmluZwURFigX4TaQTImp+5YBpHIejuppPxzX01sBbOuO4b0
Xtr6DQl4sECb7oaeafOTEONKY8Lb5C1dIhKow+BIrfyGZRhsM19qIi88kxMox0SRKnh7ik/S+k2V
p1A48T1sDK+FEPDcPtSN2EwgH9Jxsf+yLiRNXsmDJZaY+sF/njIPtOwGv4PFUeI6mriWSD0ag6oZ
fweM/Fm3zY6AolzGcCm7vRVYUO5faeGneqIbY6mrj4qU+z55ndVUE3Sk1k8Fr5e7CcreOrW44rzM
qe79/7n/06grji/xffZAVDV1/xo47LG/PMlcuC+OW5ApzD2ae5I0cOkC503tEflbOOZRC8rghHLM
bGxeCzqO+G7ki2XOUaMEm+gzmId3bK8nculpG0y0TQTa55X4gqM4bPvsRC54FASB3g+TdXc+OBhw
hn0qMCaDXUvPScu9Uolb0/X1Kns63AdzlV7+q/evBNR6Ol7IWMJ3bYg7mbq6YGULw0uAcO2WiDgk
E3cfuvkaPqZfFq9iMfehyUSaLLqzIywgUPj4wgswuBxy/+1PxJfrBc1ToGI7aaZ28oj100/YVL7E
FwPV19OW2rnOOBEwbc2UrxHkoKXk9i6scvZ4j9ynmdj12ekILv60zxQctU6yZUXnWfOadKcIJOXp
V89iQUDgqgaIz7PBZIJ82mihP5vcAd/23BBftKifpdieWrPapHu11S8/j2ch9A8ZN8y2sUatJYSk
aVurvY8eZJfUorQ4BTIm7Ae7m2IJAuVs4zcCgopvF8b0EE0py75qdzjzLbkia3/sc/YLr1EVNgmh
otzo7ppvue5CR72JFXmwWzJkf6XPeGfg4FjWBuhE2sFZja3WvBghtnzV9y+WbfMJ/fr8kW8q6yU6
ohg0glwFuRFX81rJF7b4DgTryf74k1bobRxzKoSrOFQ1mkYgHBjODsybF3kcPDUW9Gz3Q2K45pYh
u8Xdbhmdn+aeld0k/URlWJNyt0M505kJjcbrSky7/0vERUjU76g1CVxGYC/MZ9OdqJe65dafEhB4
P0LClzW9F+FdfUrS/WimFo5/ICtFmV/cB45NmUxKb5PVq5EgdjaRvvUtscBUZzsdOvobou/7/imL
3b0zKLNDkfs8AB20vXTD2lo6/mO+xE9VqZzYLhIPE+QrudpXVcYCW8otiaySWdIw1lV6+/oMayb7
deImfpWB7fwjVh1kd0ECKkj96mrSTjmV4IYopHY8VFrOuk07OcM0voMM5xDWzftWh7IpR3qARLqr
NBewV+z4lHKQXkj7y6IonfAFM3Rf7dWdOmiOjuss0lbAZ+aQVtdQjGc8xuAyKRoaW4Kq30+TFL4Z
zf4ruCTK4poXzi+dbbvqWO27CCpvwq8Chdyq1A+gKVW4HRYZhbDqwXt/JV+crAmG8AybwRzMQtSJ
ayAMy1NZndSsrMIe7G18L3HH1yDzB6b0zVX9uQSFPciE88jEMxzAVSBo286JvG/USEOlOj6iaVpi
Kv5Qf9UAKP+5xNxr0pX9GETY/VaDRNs2LchLrBVdPh+7HXLUp+8nCR1OItIKkr6wvFT93GV7fTQB
/pTRN6ALoyl07We0qy9WugJxsKQzrXzXXuDGyO7AG1CIz77LMFIamqJ6f8I1lzBDgXm2b2zUFvmU
5kmoDB86PicS3GOH02FQJdqY8c1dDKXf2yAai3eumtOMd0eOfzH94VMTAE39lSW0JJ1k0UJZGE9H
xQqeqXGwDtXFSol0R2cXMy2oqbGlBngqfCODtV3GE9NS9P6wv0/br4bicKdhjB7dpMna1cM625ce
biWCukjFZaDKF9XyP80q+Hclu7hmaQLF38m9ah0P5iFW/0/VihsS4Kk5sZNsRz/UO8+zTyynDPxf
sJH7LYu3+D3FviTRew3qIBk9e6ZUg4vX0VysYXOtRkajVabjD9lpgMg7wHoDyavVcWBDs4wRIu+q
OEvIIgFLaUR3Wrx5O9RL35+B/2MT4MZPUHsHd+eW3uu4XFyEf0s9hnkf8QnHFkU93+1G46qnKBaK
huVRQstmZE3tS/9M9mgHaJAgeeFv5KvQA8CDPk5X9opWHYbpRTwrCuCAnhpxHw7tP67JUx6QghEh
Y1eqep2dEiak344jIBXE00/oyIVlPokQLtTo3Iw/Y20yEYXtgHegWicAPM6Bovt2lCKqxypHm1Ze
gG/t6l0CJoHnwqYR9/c3wQN0qax5DGqF0oBhkShokn8t3FqwmYu+x435GER/uXVvvn0F5tMmV5Nz
aQWZmmWp/pZTYjqIN06xUYohe31lEWo8MOSFGnl1yYBSUJYnaYoP1auQYAKYW1fHg9btXfabB85B
AHqY0UEyRNutlsEmBSwtj5xpuKJe7BXfRmPKjr/TkgexHn3B/mz3atMDsc6W0xSUStCLY/rIhVG7
++fnoTvF/c+1iKCjB86ilBoc2aLed7xT4X9enskB1Yk7c5pgTKL3ALKZ7jjjqO9wcuv9/er7mctQ
qiCx5HHEzx4A1KIIbMEg6oktk6L1n3WQOEDEGajOP/UxShLhmWlb7lEm65bMsIQ0bI2UiKm9mfM0
pLVrBxA+TXmVZ+paCdqiE1Aeb5jrH4z+VGAVJPeK4mRyQuJ5qg1h5TroXkPBUVkxz+Wg1pn1GfsW
aTkkzIECZpUYCfI3wQTnvd3L+yb61RWgdJYl3UmPWGO+o94uwQVwP8+kDUXQt8zUGm0ESihkpY9l
vRz1mArd+3ZIXszAHTBHGvzp9ntFwdq07YHH7R/9Mut7VKkSpbtNS9hL9g8ZLrJ/gKzfUMa0+5G7
0jZKtyPpYaGuAoWby/XXEK+8g0YUM9gM1ZE+vmpKTdTwzpSAFu88t2ryNJC37nH+kONyDJAgvST8
PuN0nAmmUjnXr2h4aUY8kastAv5mc7omeb/KYCLEacV2i9fGVnQQ1izD37Y/q95/L9Q4vh8V6cng
lNzM0YTOEocjLfUJQNLFbdmDr8gTXnsVKzHF5002oBiemJWYfHFPeetaet33EI23TfRTF4pEjNtQ
F9aEjDdtpF2DrJcO6G+YxZ/qeY+Mw2xvMSR6xUvBefkrts4c4K0iR6X5ufqAM+zKdgzVd/CpGtY7
8LUi/rp23peP0LVO0XsmLLn6sCisTn5LyACJlNcrBeoe3rJLoXlfHyOwfE67Br7qs9ekVctRSpwE
cd6gvdC113rqlI7YmF1O9Ldf6SEnoTeoIgqQudE+kpo4WIWyJY1OOW7zroiYbjWu7xL906/geWFt
lsqCiL3h7NLa8KTTcFIgTymZ49QM49O505Dz3XkCKiRn5mhc45QZ272AqgWSSzn0byQl0/lgT3JZ
/R7EUPDuS9Z2zSEFxGCIz2/n+v4ouLMBDYpKgVsb6BW7b4hi6gr8xHbnadxc/r3CWuLNSf5J8uf1
33OmOD7OIt4+7JTKcPuNyDDTpSuWTNv/xVI+q6QBM5kZkZnGtIzcehreVHjrq8bChpTvpcCAsq6R
HoG6bGbvxHg6Wf6J9gwkfsal9306JRTU32WXT+dpkevHKEoPXapfr4RmiZZuh0INiJz5FXVYFZV0
O8cHDjr2qjY66SWOw/AmimTdn2+xPCCr/W9vHQnybgtSDv85Hv7n30xBwr42JL0G9SesL7cezTMv
dZer5gYyZuqZgGo8X5/lKhMgwur3VzVR0dwRB/IBh7Xf6DcGNBuV14ZPFniDPsmX+oUR+kE2/Jy0
JGoy1BanMiCJIX/rOvISh5/71s7q1sPX4CJ7NixYdnC5wPGNbSefkK/IZXLaxkVjZIh0OM/ZTlBK
CKvxn8mSoFjzi70Im4ZCt03QPQ6od428o+/YlrAfLhdvPg15CZNFJv7q6oEPhOHbZxArrnwdwPBB
Hvmo7bMHO6iozGrZq34ozuG54TAHcnAJM5UTbChQmFHRZBGiPBLeUVX9Y8WOZlfM4Z+cJ3xHmcFV
J+WA2Mg+kSlCn7+j6v2j8BLeqKJB6x13TxqEZYrfCFr5PPmxWl2KjNVTQpFcjhLLCXI+hN3rUCUP
WVYuG89abm7WJ4xiY2LO3BDZkzZ2vZoHXIopto7Dy7IXbBrEwGgn31bL3k5yUFnvOTflNAwB+nQV
e85aAYkkkMEhTXWBpkZRWOwMj8OTu4a93C2Z6xFFCnv8bXXvMR9VZpqvkZMPXIqbdeknDNslbnzI
7Adiwnw6r2FPVUSIUJTZQoS4QIoyYhZAsQ/7BTtZJCnCrDaxGpfF+FHng86VWR+ukd3wd08MLN8g
qnSrZblo7PrFeHnzpHUKytt2xebJ6HIi4y3Y7V82Q68wFl46CswJRoCeRdTf1K7mNMCZsYrX2YSJ
rKF63HpEqse2Xg55QhmeTYpEJTy39uvTMZl35ESo0ZEKoLZ8b1iDQpmWvMqV8zrk6z0x7WDEippJ
+Q0uMtz4Jnt9Nlsbef5dbfieXY6Br8I0nfWY+5AUWYTpqbRs0gusdcmPZ+6V0Lx50gVglnKOTxpS
1DAfF1ZwfaJQYIru+CydqQm5Ii/Hhv6yhdfKUPW7Rnrs5gVt9F3xjKej1X+UDbdNpgSPH/vQ64+p
zVTm0KBzZ4EiXnrdVq2Zia8jQHAIjKFnOae+7n3L0tklVGHYqZ7IU9v0jq1bQ9MmmYTbMW/kXjFL
jnl76i581vSXHybEibDeYxrTY/iCWdToE+JUTxhW0w8dDkDWqIYkcYlF3g4/ck8ZpewBO3z6Xq6P
0+9o3EEvwy51GW4LNxvSWW/0l7SUP91MeUKoW3blw/GOSV+z2DxlofcEDp0OkvQDb4njN0VvR7bH
8zaW97jUxCFP6MfvzhVSGChsExq5Lps9dQdfFucNYJ9IL3+ILzW+9bH7xQg051I48frTUW28bSO9
dQw4yDKkHT5//GhyLYVMiJvVlwd62lzPv/kRUpCx+4NYsL9ji1fZ4abhGbta4Zks8DIxOtLihAYB
xgW01ZWi6OWgqv1kByeATKM2LUOA6DjQBvy5a6gQ24IexzOUh/8B958J+ZE7aVRrSNrT067zJNXv
scGSMx5uFSZqWxlxr+2zFB2DrFr3/kj/SvTIbpnryUgw/xRBEJBB5x0dD/CCVGiP8JLrIs8WiLAP
H8gZFOwfWLnPZ8RvjZOMvFjU12APIaGkRB77WBSAqnRTK/BsWOP6yYIxB88aERNcmMfHwUMqZEPQ
CJXns+xB6I1GycK4P8MZcmoa6ba66sivEM+dlJjqhkXNl9STJy6z0QqsP1dn0AdD86EvfApHPgN4
GcHzDJTbokOmvIgWCd6MfbBFbMc4cAqOTdHdRNXt/2ZwJhptPqH3ZOlq/URFPTGjrAziOVK3KnbT
ZZhI2P45f27imdVp0hL22F9RxcuxT4nbtbbjFV4cXTmSqROgj74rXh9U1vowvR+QH2m36Te1BLcy
hx241PbOZjpXrD2PTwngYyoLtotR1Yku1eDIyIY8erkZQ4T/SzLMTuUczniPzj1EQM5hG61ovciN
jldzkerpzkZUXquVhijSY7vnhHDZu5G306M88bh6i7SvU+fFZKHumRWeaQWYnHSBB/auiVGv8TEj
o6a7bkD8sDimtbYhEU9x78ae9SRrOeQXBwcCPMZ+cwfI6xoWJcPRUAAqMjKava+9ngDFcwt+HfPk
H2l+i3Watcmkc8rEqT3iJVODfTm1ChfTSpPChddI3sL/4Te/Nw/aYyuyrLWANQH955NRlFdqi2J4
wJ8QmrYpSlXzp/bLmf3j7rHqkOxQeJJAzV2vOSQ/zfr71TSHeDXr28E0JsW5WU4pewaxypjkpBAG
/VKLuv9oX/OIacezlpw2cn1sRQ5dWZ5ZD849Pdj3KSQerZhl0zRC/aKz7uW/E+eKMMO1rpQKead1
3R7POWFQoMqvmdg0Y8cqqeQ6E/KjsRpjY10Co3JjYD3Sy9dElLjUUt0EidIGP8Eaz5MXcb81LpjJ
ExjytOe6rsVr65HVu2YZuJ5E+zEP0Nx0xwaDrvJba7G9sWVy/muLuSVfcLywp9GbdPVzrq6dmPsm
WKau5AlK/Zmmdluvs5vCMdIUyS/XGxDHzeumNGLPVMrGeJsV7vU5a4nS/N8NkbzFiISu6CEh+a5R
hMD/yckxJ47capko4DWNr2YvUvOYtAsbng3Ur13+v3tma+hER68EtglpoI43OsTlatULeStpffAx
Mx+YQL12CzwnwytKvVU4b+SNOMuPEYcY++owWtzJ7ZVOlYo5eJQrLi0OupNnU2cdlTU/53XLi4/E
mXEg1Rt+1/6twWb+DEFgmyugXlp/D7gzpOSE62pfDIy1Ae5pIqF51Hkk7VAmjsDeHdaV1tVBBZcb
aSfy+HXSZge1FKfIWtSskLknsL8mY4wV1lKPpwKk8c1rKTVjy4xYzVFzZMu/b+ClWYPcEhFdiCtn
CqWs7Pf8D/dCQVQeo4dZKVcqaY3Rap1FI+D+VTW84hRKTt98QQXvG0PqaOkzwGab+kLakhXfmBOZ
EoC+u/ajn63fM323bgXVr8K1Zxu1NAn5HtQ09baPfdVixXf1N12bu5aviI/P3JtW3SeSXsiL8h8a
Gz0w+ITp13hn9VOOAGK9Y4MwB3+cNdwwSCWK70yHfloCU7E9ZMleEozDpYNltdFy2OIV34xWwk6H
q1gFuPrkeA+r5Of1JQRNKWbNWNllAWBe6Zud9v0Bax8BQqzvKTKZVe3paCtt0OmS9+eNrtxTd4Rc
Fq8hxkRIth0D3tdvftfmQiDuI8gJjGlU0WJHJWSmFKKanKhmccU0mA242PwU/nwzYPZpO4jgVb17
CaC0KIINuepYnf41BhrtMtbjC+xApYCMRBh6HLIUxFBg0veU5VPeOsmbbFYkOCf8BBPnjs0JkHSR
YxDOWtFt8vaRdhkl355jOxfOmneYp0L4VUxMj3AX1Kz1dZIpTy4cW1RBXOrkr8HlClntDdOUzx19
mCq5Y2sTa60Lx+4jGoESvH9xtZnO7h/NkuJlsfPDorwuWa0ICZuiejKLj1xkPXGIi5H0IcXbUuB6
MKdSr1pR8i3SF5j4yGEGSKiQuqhRl8fPONlLnw7EQAKLLDsnFJqXogbiWf6DBv2xwN7D3bSzF9Vo
jFFwKR0t9GuLx3Qa9gYZhYj9fg8nXU+HEX+8OetnHPy9zYmju9m8yQAD1CowfYNCz83qRp4hXj5M
/kfK34t+c/Yj4BoiVifY5AmpRhVzGFYSP++jrrW/kBQUjc1vfEkAvzMkysBjYdrFWWM16HDpqCR6
hr7bOMHaSMlDnlHKyH0r0dA258uNhJDQBwKa0Ky3LliAIdEf5asWi0AqItFAy6oUnbhZelxYWGfY
ZnkacmEFkFtGLS5aEFW/v5xn6XDz5kdRvDE96F7Y8rXNbTaUXapMPtYXKr8a147m43hE5rWb9ZSp
fno5UQXweB9+SEMFGSF9+1I288KzF47/g0pJAPDgoDoO2uawkFIlkc4jRk/BPKo8B717gIGNaW8/
xgko3Owo8i/VuwTCZwmkAXq+HpHVZfmAYdzeof1RXsc3+ur82Mty/DPrDpwpWlxUqhSaGGttAnc9
bqj6GV1oDFLe7EQniIY25A59ezn+sqMfVgRkbycjHTlc+KXeFKhCt+zd+QkIkjW78DeEnyBWHr3T
ajKC31Dse5FPHSIDQKjqC2y6u/08qLYIcQgFn7eO80O3II+3X+2CPNnno0qhxzkT3p80rqmluUN4
yvtufjuM6VO1dV52MR2U9dVQlo/CCfH0aKk4NLcSkUknqJO1ALCx3GkHOTazhKZ8jFPb95WHNBp9
Pe4ugsqJc4gNLA0eEt7EG/QmSwWoS/6HBFu5P8aQ8KYY1fFg9uXzsJORk7pet1nj89uBkcGbshot
hqMTy89AvR90u/HmpLR7V4gWNI8ODSpfzH0HNP47wi6GyccMCTEGU26Vs9dIsTpAhSDcWX14bDns
KH/3BfYblqzZfTnbLZwO8z/of8FwYz0hRSHbMfhwJ4Yc7isya+NkJtEajLGVFuEKwe75TUI7BZlR
zpGqnAX3XmiVQUV1M21uOTXeYMKVCvpNXcQAmv7oWAO3qXkjUecQZK1saPigZhGto8a1zzEpN0DF
Yj6rDmfuudzwUTKzT9h7ibIUFoooM/eMgGK7CZfVkscmA91P7nEfxxw3x4lf4j388iYGrTTKt+PZ
0TgLNGphNbmxI3wIRFfOs13015+TmfTgdbinx0GcQJUvIaJwMRfgZYnvzOh9SUrK6113pECmWL19
aXSeY1BURIQ52pbNjIgWU142eEQPrNkDjp0hERS8Qnrjh4mohPatuvyzwkfobLqfdgb1CBsvLA97
8WMUCjGSvQh6QvudOQavIovU48v9fGl/zQ7i8EOtGtzrbEswx3T10efRygsuRwAlZ1jDqHnVieVu
zn8gIuN/RcltPBO9XWqTneNfJC08kzHZTxH3Meo2KXKvJI3VYPU5+UTmCtESFMLEpsPzvg9TwJKY
HxpjRSkJHzKa+dHhtcim2oPnGmzhuB36uoTqapjz9CPakTxZAjuHi8YgyvlKg7dpKcJ/+E5w/J1f
CxVcTTisWj+70FLXKa+yClh/+vhzlTG6BUMRy0i9AHmCbxIAwRKzsbMCXSNL7Ho58zkPn9+xlIQi
CnPI3wSauGhbBrj3gltTnDn9f6URheDYi8kFO/Wyg2j36dxqeziFfzuxYE/b5I3/3NPYj2su9MHn
XHt2fqvyMCuEMnJjZ4Dr0juEL5Ce4qRGETBn8LWXiBeLQoyTuXz7lLrRb0XQ5bRDmfdrMrYvjuZo
0UwsJDcudbHftx2RR/vpfqeTAnd8hy46EbMH/ryYfP/KsZZrELVp8B2dqI7+wznV2XeeuVS+xKBt
C/kWzOlPtwz8UhgIhep+vx3KOTJxn3eGKSCCdjD+jjyuL/iFLkSWuIcW1VVTI551hpLir+GjZA4K
krGbsgVEeMCfIj/dTtULghbfLqsR3WT9njhjhiM1y+bIFwciRIxeOmDnX/DgnZEwaPNGe2RptWwL
ooX7M3ljrV4BMgAJ2wA3AxwaqA378bWucIz99Uif0tIwTnvz9fLlxCNADO2yLYxpmMvJTBidtqNy
NyY3HD/q91tevWTKuhhYhMIRDM0uJSkog/n+N6TfJKjYJAGMyewf8ktw//Lm6PrP5JWqDPKGzQog
jB78EnWul4Vdw36ZjEo827ZC2Yr/OT05Ig63W3n3ywctVrHuItu93DJrUEOw1rggBZY4NBDVy1Rf
99u9rYMFuUzEYD9BP27uJ+IJg1BXk5bAFEV4UxALdXSnaqdrto6iHPMMIDTgF6qXTWtJgY6cqUIY
i+MzgVumuqMF1M80K7pMD7eHihdoL5mIV0HCUULVyFKRo72Il0gYskyDR6QK/5rYXLpB5lJ4HoA6
cJ+lC+UlrANkna5daQ0sepcpGx8Y0fb4TJzO3QCtjOCSMCdPyfwPZvyod/SkSXBgzPl4d9C/QXoK
KQ2C1//0YB/A3cP5cUbMLk5JgbyqRH5YCVSBOHMbD0ghR7YXKOcnFli1F1mIIa4gKF8POdEBROYX
UeXiwYSQ14nG2jalTJpudQk3VWp0AyIkiMDG7HVPYDfVeTicVXDoidOfaqpPrDBqtCApmfO5t8ny
1HHdV8HJ1OvyUVU4/hCHVklR6d9zwdl4i+LvVzBPUHbg/jzFMO0+UPhVmfeXkLIyo3OrkWwdaP7q
7OtZ5NBSKO7beftxF4HvL+BLn4TVghiIOHZl5bSIBn12YCzuQUobw5G8LCyYKOcWYGSTwRv/GUen
Pmz/nTGlIMt23d3eKsYKOgnn31RsIfqHBwVEpoyyhIhN+Mf8pA/sMj9eVEAPub/frDObEQyY7P+1
O8eG01VDebAWQHQDBr7Q53qEWBLNTLZAM0zO4JGUzG3AUaTuo11tTQmbVDeYhv+YCwI3PGfyYlNP
10W1mDhoiq3KX2gN63RTR5Vg2EXs/JAoECeNgH/ZxzXpJv7DMujx+DG1UzS1sQBpq/ezCUOMfpSD
1ZpHI7NuvXdXPgDMMJNX9Cg0g7phH3BqEGULX8Cm+04QwIHgQhZLVkS2fJ2a6edCAgbYHAeUuG5f
bYsIRg2jVSsQl0d4KQWbXhcOv/4bLvX8CwxxOBjNSbE/n1OZRgM8XPkYi/otiBF9uEMmBAGCtgOd
upcwYwMcJtBDACWGcjGgovmNmrNU5fezPkuSq2HeM7u82/e1vkFwa4wF9hJdqYWDTn2v4/G1n4Cb
F4ISWsZa5tV5lZefV0Q31IxJeLJnAdetp+KjTawTU8Nq2ZwohA2cIRQxQkYFIFy1M0Gr9OCELUHD
SYTQNa5+1lntEmqLN/9fCtTLO8aJMbiMef3qNeNqwjUycQC/kR7B3gBbp7gctt/JXFVk5Sj7sEok
WX+oLXB7cfqmQ+QWx77LK/qhHbFyGMTjixhES+A2PbsL0mjJYE81tqoWQEL5a55PsJtf25KUnrff
EOcsXCABSmQTz40OxI5GxFF+u44gDz90VMsbKPzFyR6O5wxTG9dxzzhf1TBWuFLyFB86Wk5n014i
q4a6v1mI5tjwtwsXbLTUah9di9we+y+QoVwBLO8QEoZD3NB5blOWYmRzks+u3d4XNcIazn9Yb5F6
79swAzA9JfHb2FoJrTdX7RyJl6/WmS6v9psMoEUKk/kuquI64CXTkBnasvY9BKEpoBvlVJjbQQUi
1DrSG6Fjr+UQKvYELRzUGtZuxRTo8ixGYschNac1bMPEaNXslPaYhmybm9oaErelSEWb0D7dEbT4
Q3ObLl1j8H90NJgB+tO/94GEi96yAcpOvfV1TO/NjzxlwehBrO3nNzcZUhAKUdDP1p37/+VYrOwj
j4MwEE1S0dj0x+sS2sNUScrmb5xDYQcIV9BZ4bnH+bIpsuK3yLzNplTkIn0Sar6I6Z06hKAnGb/2
6P+Qvbs0wfA+SO9MoxuGo/F6tYSSzvEVC6UViOCATw+S/NIa02lxbivi5ewCFv2DDVUEksHwzFEB
QJejUf3LJOxwatRg84kz895E837n1p7omwATVZPuIH2Oag+tvIktiR6450y+aUC0CkNZWgv6Xh11
Df+DowYM4U98IV3Z4bE1qB+e1kBih0vQaZelvN5TSZAIpbye2t++1fFysGC8CcWAsEvuasoXdjNI
MHZwCXKdjblmmKWl2TIllleGFwRS8EL92KFSlsRWdaiskhuN+12TwjdAV67TRvaDBUzYzkSTkO0a
3reqrZsMOlCBDmW84O8hoplzg6NdpfIjh8AXLXuGb2yveq6gPm88rSQg5G1vscmSSft1NP5VrSwM
Ly1KfP/AzDAsCpl23r07UHvIFNzekF3pCAn3o9LQirJLg1848n1coapLb09tXiqK52NVhYhPoMF4
8OwcloWfyM90gkBsHAAJDI91ZqY+8TiGc+Ddp2Ay+l8gp3e7jOSe8POof+jyY5+xavkrDRqGLPFz
0YdWkkjOnUNTtXMJVUPMeqO+vfomchLy1PYscCJsE7OpHJ78uRkw6SmeeMPtn8h+8Hi+f52ej7UZ
O9U03xxRAkGx0ew3uajnFJ2YHXzOkR7rvCgyPAz6SLb/nddJtq9zK1OIMMnlhFk4K3lgWEB7cLkL
SxVWXB9Gc0ii5qlfvVFpqqOAuFtkFY1b2jXDaPHqmGjsdjDHdeUIuhfTEXdLLiGjP8RmiyrgYzwG
Qw5hz7rmMeWc3h5+2IdDRb1AQtWF3uGdVWUyn2egD+U4KEF7Fqzlp7dZcP0NHu+VPDTlrxXabEi5
0uhAP/ep60JTqHBJS5WXgahzpqXI+ihJ2qWytaYmXh4VN4UKRVHOs9DGu8eXKW3QRlwJld9QLIZA
wwAQ6uzp+yHUCawEXxEP6mtjojDpdzWTzXX8bkRzloK7ltBbpxbraQh0qsONqLC3DKJUv02jy5dy
IoTMeUVf9tHIKWFCJLt/6kNwg9sBeG5uLJ136NwcAL7W1yAouNaGvv7suNnMeEYKUgCqiKBwZvDb
oToqjegGBzfzSCLWIK5i3lAkQkeXO/4MtnjNvvF5ErLcGWwjOwoD3Dsfbs0MjJPOcJpuCX1+yPwL
WrGHOXuTaWxYcFJpzEqTCX0HlvDuY8t60F+9WXQnBC3koZ4PtrNNU+wRi8AgJTzpSheE1Xi9OCjU
C33d3h4jTfD+L8ZYMNkO22bWD6NRuwKznUX6j9eUKlZ3FxMNVXiJ72zL+3AGd6JMDViPJu+oXZrn
8pJ5eiaPmYozLleGvDhD9T9kBnZTfjcUTvecVGjZ2mZJHGRgNwFFLcq6OdQQ1vMFSuXnerBvejUp
wVztBzsPZNMhwSFjEIrJK/YE+GNiBPAn/J+l8xbids6r9sSGZ8w6qjEZ3Mb9QZdrqUxOWPIush0v
5IbHNjyALAb+OIEINmPAWUpG5jfL/hhXxVDV786GJ7MfG+17UhX+iUY/ymXQgXKedrItSZWglLd5
PDF6w1Xx3nQN738oOfQXiUPWSrWUe4SWVCyYR/0qRlX9owKweaQtwR0ghOK6MMqdlbxACnACFrn7
bLU3BRgdF0Rehmi1VNAR/B030LhLmEZMj+8zQEfaJBHlQ/U/DqL0aU6lgFBKonUO7Ba8f6mOrYxV
Kbgh7xCtWIWFsLuPh/kwPXfO2lwUUHxT9Iynss3zQW1oa2y+yZnmHyGEosQC9OOfjcoYNboyw7f1
fY32T64yfgUKfQ9LZqzGfiqoYrXLmlDNe28oGe8GJAG/3kK9DvDOP0nxfGd1UEFTpF7hDdGGK9nS
cU0KqX79IDTn90cUDDBvoWRam5O3i5zPl0bPgSNkeFvebzrdnagx2gVwotoGWRSXsDeo2WlBFz4w
WYYXRJWolXfEH4i03kO3Kh0J3f0ImxLm8BsSd32gVwQ84BVAiUrey+aKL8YY1JqQpmSB+AEYjsUP
vYe375M17dF18VlX5sGhJuDr0VqAHhfAVrHH4/8HxAldi6X3/A8pKO9MTYZDhc3mM/E+QV72dV9t
IXIVZk2d/PDWR7IdVWgPjOviCnqFw6ifAUTeuGGuN9ne7wyZi82Yu26RnnFWzL1geB0JAcVY5tz4
/98OkD45dL1uxr2KSEQOx6Cw5YGh2ScpRny/GHHPQQ6dfciQOYYTLwsIUaQSaiReBbfhzIba0BYX
R8xoVkfCVHDUf8tLzvuGKJwT+bV1WwmHXWH5N/tDL3EraRCh1Lt/w+8x5d1OooBJYPfBBt6er0EI
XtRDGfzPhYJaOhMfRngfjneFz3hBE89kXutie1v/ulGXywZkaS5pvfdgOQ2Xy2peLs5i9wrIYFGb
Fuwl7DF4EN4C1teJ//LE3CNO0+deyjbOQuyiJWs6st+DyZ+hgYSC++x375BlvIEJvHj/1MH6IUFg
Ng3ZCAb3PMvSGS8h/5+Z7ApRBMI7FRAL2aLcCBu4vK8x2MbCV8xr1+j/9OuB7M5Pi6LOZL3U/U9U
3ELMBXo82Rp4z+gRC1FTIkCTzdvAPiWAD9Hkm5aFloba7Bfjfxml4LjLDDawMrsfHgpN1h8AbuPp
IeOjA1oOpjD9cbGnje5SrJx8Or7M+VIYB3l8xLncYbMZmPyA6UsP3QovvOmcgMbJzB/vTjEDzOkO
epTMYTEMpwtMjyyyiqJcDdcz31yEI2ZghcgYaL0i2HPks99+L+vDuLKwJhGqp1T7NEyst9dpcHeG
Wg9Ummzxl7OlOAIAGpUNqTJ2SMjHiCWESMdeb3RyvLfFKWD0a1PWxV6cb6Bql5xJx/aTk9zw9UrL
r9QLRSrq67dHIp9r0NjRgi/U8o20dSfwG5tXF2vFIXWqBR2GYN4EVvlAZVzAey4scUisVuwpwIor
QOjRT4ZjoaGipLOHrQVf4eDu18B0FxJ0PZBIskc0cH/6TQZRuBgpRz8GSPRpOOzZIuTvp73m15Mu
0GfgKtkLk/mkF1OivV0mCTWnrRD6laAIEA8mMOy+r8FBhLpE2UyYICMP61jZDEx29tsG0rIGUsuQ
yNzGgRTCFH87YyBvFexA8CPhaYxO4Ezf49R0svnmaZiEtxkh55mFBQlpNcaaCnbFgLvbVWhe/Q01
KEwGCrhxyZedkTcsDbztFMYiwyh/lAw/c92QvStVq55Vn7Jkdt9eEdF0lJcVHhrUOJto5asmXRYw
msLNtHGOVZDUoMRAraa05+n5TCOKwb9rKm1sUWfg3fUEIXqj+Z7yPPyx6xnh+bb89KT/dCT1RVWy
6q375Spe8GJFD9hTAEtNWOMzCSEF8SVeHnj8U7Awj35Aw8mH3yxXfAkVXWUJPIUC8OLro7cScmS8
fNdltHDdn5nG0sOmVtXq3mLuC7QOll2w9uUwLABCS2s3AfUTr/vfzVQy8vLlO1dRRGuMQ07Gmn8Y
W5IVGTXHb6GzdrDRcACkiRY+vmPARagYtnM7HMmnJ3lfuNq39e/2Y9H2+V6ymlqrydftS1MhDA9L
F7WFTDDrrX2cpr8g8oTnycui3ZC2zWh2HjWjgMTSFiHNEH4DjlgUqMv2vKRcNq51iB6HpCPKAEsI
En3rLN+ta/FcnaEUsCpapO9uB9sxQuTRb5Wgd2UwNpLTnjQP+2OY4SGYdzbadGzG+uGWWoQJNAIQ
5Utkadf7/AAlmZgF295A+O7+hCoocBLN03mlpzHgKl7JGwCUuNgc1OQ8YvvQFay6nDFWvzrrw6mV
w/QbnCgGI+o1f0f80mu8jOqPmwEMYh9rnyR2r+fbVX/FnSlUrFS9MttUSCIrdzFj76Z3DjHeOtjq
z51wO6WeFqaJGMYPs51CzkJ1v3NoGX9r7ySjRa89GqhKlRzNEJeLnr2aL2yFxeEpKoFL9cg/GlBH
NvVVeENItdSdL4ZwCik3MSq29A54MAG7jqdSU/llf9k5WRHEz1mInvErBi7dKPZqP39/4rWR0IL6
zv5RUILqpZWm2V2LTowMs5zR6T5Jm/OLxoBf5A5edlryCUqW4wg5aJzQHWhI/FKyHIPs9SaHdDts
kqhNJpgS9uNhayT85T2cp0crasTd3LUJuk8c39FCZ3jK3v29B1uzNUYNlT5p30SxBnLplKS6otJZ
Xz0u8S8/ZiWzj3wpG3qmPFKWKjgyRRQBaZ7PcfEkQgjR7iJUj2OXKO1bs0sTCSgwxCOIpt/HWjbQ
mvyh+0nuMgkxWYd7zdrt76opsVxnm+E2hSKg3URw7IRioa+/TYEAE2CXrwcNCMTm5zcLG9YPMrGG
uf89DewPTnsd84SdB1JO8YjG11wE/4/8HBO4AMVVzZJ0j670m3XF5i1hZMd7z963CjLucJJMtBQ/
96A3FSGRx2Pe9KVDpPEv3plX8cq+Fjp28X3tGFjEzuBA/Kc6f4Fo46dEtOLEOQvVqF/FXhuYrXfX
xa+APwx3ovlharwc0TYPWgWiEPsw6PMrG2w2JdnoNqr+4DmVU/mnZv6GZyazd+TD86A5QkuPhWCa
W5DhddHb5s5otlUi3NDkCrnd2pLKc5i20ZP5Nxk/1zRPja3LoTbWPjJcJJyUS4h7QqKavL8pljTu
UYw3jGaDDkBrSEeBsJSzCQ8uDgWSDmYzHZ0+MCyrRro80KTje5fuuRWo6JpfbZW3D8OU+KQdXc6x
bf8VNTgpYxMuyuUCFfyGm2Yi4sys8NEOhRbOsB5qrAeQZqwVn0b+zxn5hFdkY1Fntj7tQ/eShPc7
fDyfBywcGlWtAUzTD1jPm3v0LrX1lvspb/+6AiO+WJduQNmGBPI0ttmiwedJSi9VKvzc9Am0s0AY
S9M0maY/rj0pmybsEiXRfkztdcTmBKmksJDVX32fiBG75BOYvTXYAAPFyv6bCJp7E8znrnl1R5ca
2ALyIVeOMTusrAWm2/obZ9jddPmPHcuG131QZe+O+9khHhJZpjnt5tkzfVnoQbY0qicy3nV89sdY
vjX7CO67yekuO7tbhMoRC4Xa0x4bdF4Ixls72iZEsd5jZ/1AqrZXFXjZgSG2KIdfB9KyVDPs6Hvk
wm3PNNdP/kKMuZDpSnk0ijenLQaTYyLtsunGZ5rCWzEithGWvpx3GTxnpTa2qV7awNRqj7zx+/YX
uISsSmd3pUCTmWDasZYwa0pCT3Von4eZs5yL5YFBoZ8XJx7vEJ+9if69Yq9exIR3YlC6Qf8w7HLI
EiULTg5CHQPFjAtRzB/uCEMCw51jIOpUO2bt1IXVExGSTWL7voAqGqGdoU6MLAFIzsPO7FaBcmA6
tEqwhZ8a+Z2vFI9FtoFZoEaGH1s2anYBRAABZ0CBhW/LhPB3dctv7tcvGE4T44KBEuxabxnpIUWp
Z3ErnpDqqjCHP+nmgr2qCGcnSJllGPAxXqhMQwusvICPyDFU+eTNbYBxE0qbm/UFDb6dIDNpCvHa
TpBF4TG3z8svXffDjNCvmR8iCMMKMP0oPthOb9oFZR7IubTHn0eBQGWV2IdD7dElR1U39KKdfKPl
7T5jho/FtHduPvva2uDRo0dVY9QCPFqL4atytRXUA7CeO80qAH/TxiadyGauCNbC51ihSYTSXl1Q
VUE4EJ2gZZE9cVS4wSYqmObaZkSlV2bKcBVZhlKhZWHcn10sTfdAIzcn/maJjaXMCiqH0wJK95oi
+ALOWHeRiRuLqkgKJb1QjhaKA8b2+pYVx7PfKX27eWRmxJq/NTakcfStxeoh8yAR1cpFR5Bslt+/
IP1GXLXxbvbvApPwe5s5wqDaBUVwwjnWZ2UcAKFoNBswyrLYBFZMoDxp8ZKRFWsQgiSBrf3YIZsa
jPTwG1G/J4tOeUPu6uhEsPYWsl2j8yHWMLsvjS2ik1XjPZ3H8ywgeLezFRf/Hp6udHfSYGLTNarH
aAtGY7mSu6F1HhqaLOrbXHXcyGCLRWGFwd3RBteIuWRQrzZm7P1hvFVED2diCq4OCf5nKUlx97m4
YAFhvThaOmC772IaZeFuG/cT1jLTvqmER0gmbUuLgHmDbndzmy2X8nypSQhobgw0K2HzzYPdnWc5
AYAetN6asBFWd4TvUp7zJd8MeS7IiBxv9We5HhYnQ5sorSkwnxl0+WLr9rniV2cXiaD0WBaF2OyP
nGabhyDUdTYf6zyJgA0t37vQz0qNC8TG/npeQHiM69YHrJD84XWuMqSJexcb0Sittnswn5mjFBvD
R3k+VfVH4bKfT52M8jZcThUh2+Iog72Fr6D1RCzKb5kCVXixFoQ2ciHFifMcAoQ5l+vqTvtOvxYO
bsHGeQgf7RDKFxdQmWRcmhWv+F3fJXxJmDiR3CHDPHN42F2b++Av8gLM2EAlhflHqnttSpQdx0WK
wKtLryiJkAjN+hx/Rm4DiSI+GcuGg+Q394z0BnbKW5A0zdBcrya0VKiIL5DqeebsSy10pfoQGxbn
vS8RkB0LpRCdvqU24UU1e5FPAT8qrkMa8NJd/MDXHa5HsYKdo3v4ebRvqTToL3x3yEXqBo8B4QKM
ABOkoglIQ8FBA2rdxr3G+S46nZeY1Ep5M/yFNJYxZ6nsowMZHGXSFbMP+Km83I45lLRW/6KP9+Dl
sbEVSqFP/hMtljdDSKRg0ThmueGx1ksqr/KZ2e8hcE/BJZIjClN+luY8Sx6VbSu/eZpxXzKw/fHW
ROjTEukYL6md//dwH6wUsXGiRWYEIhC+KKymBsLs3PqPY8RVYBtf9LKqLAs0Lacx6LQ8Emlsx5BU
Ra/ycI+O1mkEiAvjk4NfQl5nJbTFFJPywcKYKyzkoIv6wm8TH4DuceI1zCIZfGimagFg7qb6VMRU
tFvSgVdxO12yDSqoOetXMPokt5SjktoVtzT4RErwkccmqj/dhy12R+rFulccLje+q+A6HmXif7/e
voIU16m5ZaQuwGvh58m23g14GuKi2ojaMKqlNArx/xh3E8AYUa348km4pbtgfNXVqL/Dg/qdTa+I
7+jnICXlD6VJ9KSNNLos/o8BnFLGXHAWl/7gWT/BoSTap9tq5glgAL/J6xLBZnWVy8YIL3Y/R2Cr
Z4sxHvi8s1mWVFXiABzhAwq8blpGR44c6Y1vg49g8E7RJ+F8cPysbAml71MX8mPzDdYDRJBFQpXn
N+LgeFzIMHqvUugfYxgaNWqpiCmCqN8N4TJleSVRiH38iIGKyNBQ9MK+HqAoe7ystcBjKG5OYSLJ
B5zMKm+RyPY6alf3AtFXxDjT5L5kcnJ13Oy7WgPlsPwpS9b0qjmXORQEETmQ4n2o3YX8iTv2YGmd
9Rf5ZOwQTF+mAWWrhMg1p9my1oEize/6qK3H2fo9SBv7vnyYAjqfKRJyr2MCm1B1sSgJRUtdT44u
7K4Ab0lDMcp809JMPTTq71fjkrPXJtSbpBjoTfPsKwRJdjdkLhsYw0m3L0vdlFMU1+FYR00RyjUY
UUeIs1mwPtuE0jlWBN1PzF49Xzb5um1kM8dpS/7vTz9fNWN+31H0j1Fi7EBH9vTnozX3l9Dw10IG
VWz2mWYeIbef1P+igT673LCIfcN1E0tMhndsvhlf3eoQ2KFlatcCdrDU4KWqCBsGZVR6M94X1dru
W+8nS3Qh00cCxkH9MxaqrggjIz7U3X409CjXMAWVnwm3H0eqQIetsvgtD2+xFd9Ia+dvhts3pAkx
n9ENyMx0p9Mln51dwWAt2GII4lXqzB+ykgM+xuSUf83YgrpXKA+JzEk02bESZRLEQ/z7NXCfjqfd
kzElsPv40F5TEdEHEx8rNd4RhtESijK64Z+cC2OiFc2bD+RHzLakWKTJPN2l2PYSxRqCoTrGtjw4
hxsijeAuCTIo7UqgHk6dQyFnCtQnaJbwIB9csJ60HQS0PDmxwDZ+pjdojq79qV7b1xZZrI4gNUBY
qIbCVEVcbZCTirHgToNvhTRBR3o6x4AuG15tDi+an+Yc2qYFfmii9encLnh3MGDM/G0pjgL+nH5J
m/eMKDhL04oLzdEdqsjHPmKr4CnVevfhsCReL94uabvXUV0KgwJhFSn2M9KHNPvB6uiSe+q6CbGV
8xBvaw9LxbeDJPY8+XsawJbssFgLzh2SAQokWoXQyrhS9t/IQF36CkV63uknHSLIn7iTAN+3gaF7
gBqiwnNQ3hSc5D8K6vT5KOpSUHiIwNRWnGkXuYIatIwdSenux0TSfJULgcIUGZsy++87q9am/1fu
egaZX4CjRfhMDH8v0FCcFeARUe3foWoDFcBwHlsip460BhDZUJos9HFXEQLewWoPo9ITRzNrY1K1
OAvTpu3qqApcq2FaXQVZZAevA9Dz6S0GwfX0Fc7BSwsxn05Ss2GQoj9YcMIDeXIOkaTWJ0fE6RWf
jplN3QOypWOzTcmfa/9XMwxq47z+fibEfwzexTMNAOupG5BUIF/v2bl7FBVk3xqULeIedGFlTbas
KuDyqzX5QBMjQ6yZ2c5+v7Y50yjtpVYyLLP/0VquNPYl7bHjvq76+yI4cnOCSC/AtCgUoptJQuyh
1XXsXPgSYE0pl0KsP/g9Hos1v8vSIORHGxKFFm8x4+sG4a90cdmWsHrgXkXHSxRuWUWeMT0LCqGR
9htgSSrGAci0es6ScXuG6MKWy7UGAiwcwJNjFhWyF5cJZ/6ZqFxfw9INPzm1I+V9ZAGzdx6xTEFz
0OSfvSvotOm86R0iCqU/j5vtyKWvOZvCMdjd/ckGkyxqvXRGmrWW+DCNLdgE3YEp4gq0AkDs/XAm
lqSa9n8SK4iB8kjQpAtk7/XrpO2rNfcm4eS9JPgRPcZ+9141vi8Nitl2sbcDJGjk8kXfDeAFOSUv
mNQ3r+T/jbyVkU+AuzPw1MKbRWzK/9KlDz7fmiQR12PqXgFQcGpPDS2NP4gVJecry3WFH3bOO0vA
diF+AIUIWqzgxioibfo6xMHUeqmAQd36YjRfvmcI4lUxGwKMiIeBR2zJk5C7StWaK01F7OZtYMMB
ld6MKwfG8x0YtC0xcSg905fEs9ZFUkaMcnZqBRC/GjiNLM7ThVuBfTo2r6+cZx3spPkq9Pyiqk85
oh1e/7wjIq01ewtQEBhEmQAqgyF9YKvtDyShnitI24D+FtizcR7fvDHA1oUz9YZTIUK1a/4UFfg6
BofqSCyFZUlNjhETW1sjkkVsYczgsACxs9UcxBE4jjIGkDpv45ZsdcUGhgQBlrz1A/j5YH2IcNBT
UsQnnwsOl39/HjN/BTqzZNDcY+mb36+yN9odHrw//WE3TIEkEEvswbrAO7zU3yUKJQsJqfPj7OMX
M4Zdgw3WwEzNGdM5z9I89Pc0egOEKYJqoEj9BsebvVRRScYHQw/kqzsn+KLLw1B4pp2itfjg6J/u
LpYdHqVLSiJcpA2IZAhBBxegBvhO5jcOivRCnHXV1hOSMF4XdysbrQXqLzWrOttX3o7lOP4aFAa/
+fGI78wftB1BTxw+YYd5NdmHiY5Uw97Ld5b1xwR/SwRIvxbRhB6Ic70QxcPJxZAdyre7LfFDTgSG
Ys2oC3yYP2xtEnehS+9fb86ftaU25DSvVhz1E79Nb85JvbG3q2yb3zVJo/O1jGh3bN+Czclp8sdc
z/ZJhH4GwnBYq+sGhX6iOg0qJMTDDu9pjfOkigYwZg1TqgoW1PrwBn7j8JFIOng/fZltVhupSk0u
F6TvXhKx1fxAGLwS64sHa5GyJ7i3kGA1ekp32iSWfbBcrVNn+W6tEB3JbWSVOeHUU7SCgb3bcFpj
kZDhk9i7t/Lrtoq7E+2F4wJ/NEnyQvGr+zE+JCSRjaWyGYzezeQkWrZZYmhrn8JLY4ysbpkbjllY
nQ36vzkzhdXzRfKHgDHEaPiYdD52mHkDt6lwKigYm+YpnYruXdaP9Dlb9B8OndMsdMgZMW2cXTy0
D32WKWFqLGRzZeoIhQJFbhgIz84VbuwDMZuZr72r7QyHfJ+mVAduw2aTVtvnHm9pIS7UoYe35bP1
sxuRbVswDMYzylLp2uiIYvuf7gin9yC6n6HvL/eoiVVc4BIlxlUN+WEJYrbIAxEJnnuTBWwLzh98
xwC70rt480Ksi/8li9pjszsnw+gOjUElMaz5GwWP2EW0y25c3EcKd0A20h/Fwuw8QiMayq97aqzn
9Wj5kLlstraE3y9lW0EFgIsQw47PIBKE8jRDYZH0Hkf3gO3aGonfoJXvwhdBh3DryHGOCFbdsyGI
DJ4486uch37N/FHOxAtH9oauXPcZKir8/oa2s5KMDB14q3a9zoD3AL4iWjZKpdVmrpMRJ9dG0EJx
xPbszeCfNtCb5CEjP7ASOKnq9dgbk1eagMRe5j2DRFDCE5R9Zw3nOihSKBEea2PgvS9ZUtJ7OOeA
5qVztousH73BaMvE2DhpqL7amD3wKWirtGicInHtB78kLvy7R2kbiG7sYLT3rfWO2ZwZocn5mRQ4
AFduEy+at+7LLQbOm9MVpAu9CHEhFrxGPTfre9fqwECHhWgxix+BfHbINXPten7ehyjpNmANiafm
0Mt1NOtGat9yu/qQYXIQxQoEW/3YgjWZkPtrpsUoBcf9kDuCE4EVMpKuhueLq42Jq2bpPtWfLqQB
XM2ti8J7k0d9JwYWVbPJMaU4aNUwQAxf3taAqCVVWcqy/myb/AIMAP14n3JgWxDhNRk+6RDQOIeC
BFHOyQSi1oZJ5kLJT3TwCybXlq/0zDRSvcJlwwT+rG0stIrH7qFg+E5gRN4EFSzfod2NTknu9yUy
yeIgKHfuhc3Dl7yuO3xw8ynArl2h/eSQmQN8qHC0F9pi+JamMe5WBxB+oEnji0RR4Sw666W2iF0I
VOkANms07H1t269eTTAbkp/upJRa0G0nQt5ZAIs6z9UxqLK6d6z/bqZy5oCU30K2GsJ4M28wLiDm
8AQw3gndp6F1v+bpiFoXLUh9AyqHVNzo1QRH42oXkpYRqD/aNtDaSfzyL7KajhWa2Zu1z4wvGYU9
i0a2fIdOZoksFYDr3vowG5GlZ9+ORc2n38fAfAai6+oVsPS8SMRAoKDlXy+dSdREwDIDVUENiXMI
y95cWfDsxFWwB2uxQqvkWIXl541fJ4IbyabsFiYATIB/itWbDh05+tOtxv2hWuvjBuA8wSj7v2Sa
iQsbLtPaka+OhezZGpcrSNUAfZ3yx9l7s/uejoGmg6zRsMOTdkh0sO6lM9l46Y9y+65WHp0pvi0g
y/+oK4XOWenwd9os8SBUrx9t37A94MSuqvk1jNJdN3hiaGDy2fnI+3WqIsqD7hpQiODSyaslM/pS
rGcjYbDljVkjwXHT4e0Z/e9yOR5ubNrouv2tHR30uwCsOIj9woy4FV6EyeCu4qAcdpc1uWKMVDQf
jGji6YRMwPMs7SJni01aC6enOXLll1SAcJ6K5oCxjNE7VIyZy5ltiZbBBf39YwJ1mH2XdeKJpYlZ
lmSJU8KB9yKx9o6625SM7W8NjHESUidwTreqTXgAlfDosZcNtMrhB4KO6HeMQlgd7jHXast/L/E/
P4fqCZcuRdXXhU1gTWldyvI7w3c0Pd6iNBZzDVY/0/8zw5nVKMHvEhacClgfIHHHRRfn+Gi2RsUl
rrY0/B4E1IzubTLGB2KtTOGVCUv959a3ZJxVzUhTTyUtS85B0yxVYn1FOrCDawrDWqH7S/L+830B
atCOUTH1UgkJsDELKzsTMeyQyLf0ea/mX1NZT1oLVkmL6oBKAB5gBeI74ZHtJU4qnQ9ebbhDKV6j
YHQGQ8kU1u3GnRowNPL5IbfqPYSn+8fk/mPWUVbxq0+f2M9e/coZT7Ft1afxj3rvKGb1l2ky67/A
nfQvjL3ehyRlWZRJIw5vIUd5kfP34Zwc8wgvzaE8ZP5JMEBEhB3G6DVLUC9M0ilrYh7+0N3ZfDFg
ST2P281DD+INQhT9gGA4y4y0We9IOqjYhIgC7IToPbZzRcwwolJFhwMI64edi8V+g+cfrAA46Xim
8XXCiy4BQ8SOHq7XpIW5CgjEXak2wGNjrLvm0injtiJK9Dc8i6PYZthadsMFYh8p+GyhVCfGkBEF
eF+13zZlg9sg6bixp7rCiI054s1LjlPqmkkc9lFV5Z7Y1+FKdX1E536/eHz26+EAXfraseaxIu95
Ye/0wAkomRygZ1A6NUEkmZgMP09K9/4U7l7WRev2yq1WREv7PfSoNcWvTWdaDBkk5WnKp3xFYJLy
m7hq+8z8n70BVOwmR1xbrDubyA5sHhwMeYqUcSOCvrlgnCb16xhI5cqAxcjVweUh8K0pjMhfnU2A
sRoT8X6PP7KY/d1xkraLD94hF9W9Rtax5hv8ybNbX7jVmHqZWRkj45YAoVSzEao7xnLxA6roZEoQ
BQrt843Z+31uR0seqP0JJ6HStVpKScX4JO21R21f1CSDxzc6N27R0du1yyq8iJSzeI69jotnejeU
wv7W5m8RUj5BOsIcvX82YngxPW/myYYqKZaJt+MAT1TObQ3uCsNlZd6A3WJvQwwbgf5cfI/9UsuA
8L5DPTdnSb5cTyZSFgt14K/X3TMcBBfMXky2P4X/1JnE4FxyOZxP1RsUmFoNJJJ7gyhTShnWZ1Do
mqDQ9oigApcR7HAewr6Leq5j+TP3gz+n4II7yqSIAcb7SlYwZpVRUGoSWCtHV+o66woE0ZVwv7eL
uIhosHD8jsw53YY+EMC5W0XaoM2crTvVqmyeRG4jev3fSCv7CJKsrhTZlcV+rTBZsNrLIJJI6rEc
qUW94F/OYd12ptMRMoUeKBYJZmRrKTUYVBeowOrr8VHLLQAsuOyw7hgXVG21eG3VJ3uiCTVZNDWD
PZuPrbLVjLcyavAYu8O5muR+M73zIplhyHSZ45JAs+BI0otS3yCkIBGT7+eT3UFGyd0lwD4YAM9L
rY7qvDHn7/oN8t7TwQqTUqPe+fBNrMc8O+GpZHcbcBqmOrulUchuI3hZyB4DlJKa4IjI2F74Hdpt
b/rHEJUUZf03eKvLcuAj2eHjV+E/VGDaBZIRVF06+sluECPQslJNm1+7lzqx4Q3msrTOcJtWOmjM
Ca1lMM0mK0ie0m4CYQ19/Bkfo/DupCmQ6E18qd6K+WKZxjXUbh5y/Q1853AF+0cHcl2Kjz16nxIF
flyeTF2RjPo5xAznz2XTeuPIujkwjh4mCgCU/TuSMw4PPHzJTaOEox4b63ZbMJ+ziFs4F7snPCCn
XL8rosSQd/Lg0REjvkSd/PxmnEVX93XrCEPhVRBepZ/A/3fu4u6JvcAt70m5O/zD9JbbNFSxZAaZ
6hnkUhhXLadelYbFNgk65o3gSzHD7GebusMufAFrWUJVG4Ry5fTOqgJ1Ziu0fVWdGtkOIa7mwAu8
zDBzP70g/9yjX9mqezTrh2TumP8sDZEXa0pNfxX9n1DVvtb5IwMiKx/ErRwV6lS+PdENcHrQFysB
FkwCfne1ZVPMLATritlbUEq21B9OQeOiL7BB7c871UdhRgAiRChmqMFHxGnhCPU9Gjxp+YTG8GOa
T1a4ZMqwbIxGlxf1BSG8Sv1wpB3oI4LhkYKok2oEZ0XIMMFNo6G9CxqzB9X4Y/i92TKGbyU9TcFn
iodqzqPj9hoYfqjurRag6v5UQhwa4EPXhd3oTGspbHxMmIC4ZA0ZOq0z2X2vN8B2bd3KMQQGllKx
P2FEpfRPsv6cB5Rt5nxQU1oHwBfU0RN6seCGyRX1F8DVFKcBHJUPzY2f8TusH+fyXlIN50x9qIFI
kmCd3ffVky8E25/c+/uxkS2K+60aAjgOV0LlD01Dcuj4ivOSRJlg9QwgvhsuftTapRvLphLliFMn
dYQ83HnSb80Rfoqvah2/zgNe1wn/xiLu/YVq35XKZeHneiSagzPWqPABEyJn4+A0yzGotLlgdkiQ
/PRurKW2buECtUu3ZK2wyXd6o+3/gPNYzCPwK4junhkqXdDO7xkmYftzMm8gexA1014K/4iSErcY
8aTaxHPQuiy0MQAI4fx+K8q8myVGksYeQwBlBVkVQ5zOK2SrIe9FcWUgIwPpJg0+zuxmN+c7iBJd
gXmYxzmjzIxtDinh1cOlywLW2+sZszW7MY4LvinBim4crUi8apTRLeggx9ptkZJYAUTn+SA4kgT+
kSo4eKH27S+wwYHThFBf0Rlxg3KI9s3+v5ckotvvh8mv9+n0hkPGWh/8B1NcDraDBWgxxU5KELxh
LeR6QYwxFUcaHNSpTLUjjFDS7w4H+9RWO5ogU5Iod9k5YlS3xuxFiEq/6f+03inhtLTmWW0xbrkF
uK78M4FqUfex2jw8/Ls7T1ATcstUroe+Z1wRs3Qkml3nV9YqynqWDNvd5qPrajTgvlxx8yZa29Hj
XWSChz+Q9eXaFWVN0Ba2Pt6VFAVdEwBcRiNnTUUe9p0A8GBniArizOdtR8m+2pk2XkbSf7Hjdf8R
4j/DjuNiS9crqgOIYWqxN/giWtstYFSa6/t+yXWNJZyYSVntqPtsXW6Et3V8W1km7zkFnq4oC0rb
k0OaC4J8/Jw3a2cu7zi9sW6JzJmj29wdgHIoNHndm8fpo8AhycuOEUaRE0dtoKHs2IobNDeLCsIX
csVTgkvGcbiUocmDg1M9yraN/uQXyM2aZwEcaDSqZr6iv+4JYmwSykzk1ruYLHSceq7nqeCswvLn
nJF+LsNmOJ2FQgoXH2Q0J5/QEkTBSoHbcAN5rs2701EMCleKP4kEe3dxlqKaslqMjETKGE2m0vLC
waJjYol7yMuLnHImVYWEsL9GuZBE+AC5flFMLHfMoMhljCKNPobo5pr23Pf/83jNlTFyGpP6RM90
qzRT9K1iDtMggkK4zLkmyEB2IGGAN7jjU9RGknnZhktzfCT5p/l1CH+WkdLPcxWZXw4kOTBNmep4
O8kppq2Yz5mC3d5hW99LHbpHDwTnpJmphzUcLEcuwI5CVir250hOI4NqtisH0CYXt/VbRSb8hymt
IGWz9PEGnaanExnrBPULdMp7QVuhgkSQGMA0+pr08uZYkN2gk663TABvQqH3TjVaIN836//CaoFQ
en3//IwNDgmijsXWGpi3oZMWv1dIFnzZcPXPgccD7zH1/dnmOo+Tptkg3edR8lKeA7Yats1QsFWM
txJ/npNLZ2yw2V5gmM5CkNGjZeXLpY8+0b/4UBwsmSs49tx7vawgH3XlFIszmcGu/w+MxAjQ/4Oh
+oKczfgUthvhxub549Ma1kW6HZEiBKMOaAg5l2Ti1ER+iP3hB85lr2yamZOzfs1y9cFU7pamL/kw
QTD659khhXaX4MVypa2/lihXyOcm89xPnLF5SvBlKJaZ8s0Nt4ioT3Ow4AUaSSU1HrX+VBnJoscs
fmLAxd71x5hb05fLGMN9GwUfad4CZKlLzJHQX1A3Ygxa9mC+fLvYB6pIO4EHGkF3Jv+LAlHDPtKX
48uR2DwHsPfTNl8BDp+r2XJSWQ7O2TuDZkpHqqHwgXGRRCnTzYScRwMVTSyDpPEWxPmRKpJinl0q
zGyWp/NNkSXMpLJF+XEPiF46iotNScndhftFkRhEEWLPUiR2UUAav5tNtyWrqkBV/qJaqU0hfY1y
zdG1SGh1Dv33HnBxwpnXN7zarOgSwznvZmbTBfGM/fpxUuFji/E1M0YyqG94MgcCsqUrqpqwA5c3
0a1+FIzLwc/vZUoRIDiGKu429bMc/fLhnCpTZ3I6HGj2IcJa0rpnU5YtYrkP7BrI4N/5C8xKXxxf
kfmdHuqWyi/5Y628WJEDjAlfjsAgYImJc3j+77sgJeAxjlgRgsGOLBGCKACTxIkv7d8b2ilVw43p
VjxlEEzoTE2idCENRkZlKsRWePcZp0s9TTq9ST5OiX5Bke75QeTOnW3ShGqWAGX+8pr/KIg6YqH1
kbpKWz1m3HXM0IoqUX6SMrnV/ayus7x8ukibDZ39uoDtSRtSQk1teU1o8fBemjFWT5Yor7gM2f8L
Q3diUEoubxMZSULDqcBCBUggIf8SwchVioNssUWS4zor1sPMcn8P6dGh33G3nmfv4gA1rQ6XbB94
OBrUkMhMHfVmTXeTCJ4/Mm5+O3mDwISYtyp7WMkQXYVSkHOhyn08PqNWTGIp+IACOV8ShT/TNR1J
BUl1aesg6WeorxvqCoRBSCcxjtc3LO9Z2QNXc8XOtqwgXjgGBvd+/c6uuXbjNbYYpjuVc7NlQhBB
0PMLcv7g4zwmSCTmMi1Wg9OHjPrreCf/M1Vp497M2FmR1jXK4Eq9dyZVpJjhF1m2ZqVprSqzFuvx
RErWtGLHB4v2opyiOnGv0HXDcP9Qxj7mIizlaISqa42s2OT9AKE1sPdWKSg3xj374z6ghHhCD112
PjK8tl/LI+Uv0veIE6xs46ABJ8n8S+ScYEoDJ+/UkL5kiIetvDOvNhx5gZPfcIa/gL1AImXoFA1U
1QY+8ZK7xoioOuwKawvheLjyFH+6v0i9lHYdCxySlod0vT9TzKwVoL/aRylWc3b3AjPGzwA6t5vK
DGVfkrLgpNF+Yum+dblDsVU6Md4ZUvK0Ap/wTpk4msFxAAoihfXka3PG+P29WnaWC2wDUZnBpBqn
NvYwU2CMkI5+u7Hyl+z15D3Sao5j+aL72wMEPM1u1kZwcVXVmyHcTKdsF3ePJ+/lW4yR72vNmZlH
u1KLfzXvcrGvFpFTp7AIqdU0Mr5XVN1fadElJj4jn+uzqnGltyilzQfLHK+MmuPbH5S9F+gCIgWi
GdS6ADvkTK6vPVPojRJQ3dGDKID/nrzh2m2+GUU+8RMaOhQfW9Fd6xIYbbCdiGXy4qonSV7Qnr+b
wgF4Y9/ZEbxOXSZ1zq0uUUFd68l0ezlwiOPmKdK3rvnBCsn7Tli91MepfoR+/j+CX2V/QY+6dkoI
o8T86c7meqWKIUsnCZGvZUdJNcHBy6mu94v/e4++I0FLjo/3IAe4lhaA/gqf7XAjEeA1COrLBxen
duN57uLwAWZuvKQWrzK+aMfPXq4g73a4ugs2Q45uxnm9SEkP2QL0quSSa/amE08KSXubBvc+IpVv
Ete+PuG8kcHO9nHPWLSW3fZd9JIpKiJfVd5EngxrroLRw07E8WxA2R3qxQme1bCElIs8TIQIrUwv
HG39Fbnyod+KOubT5ye+s8VIqbvwd20r5fg9nJy9uddkSAi2jCI82PYWjE39O/8IF/v9AG51nxbO
GAMN3n/xzLC9UVNjopHDPjipZv+oN19guiBvoD+kF9dtwvrG6WFCTuO6AConmKV3v4w6LLsnBB7K
cu8mSvdneAbh0zFUEwetrWazPtntvMDfdHxeKy0t8bUOPcy994S9+NPCwpQrNBnwJiq1UQOThXmK
N00oDE97LGpsHPG72HP3cDXvuoDn1iJLfBFNe9n5hiEajHKdirfzmhz73767gZRdNq1LyuoMT/9a
VqO1ZC+KITekLXlOqSrNj2gxrYCSW7k1UrS8GvL7JjQAaHSiojor7Sh8RXDlJn/99LAXo4RhiH/h
bgfuB5zT5N9eo6w+CDU/uR9woRDnNK2z6NZ34tEfPOZwfKeRNCWXtYlIm0MrqtPCRbsfOJoPPjI0
Kv494HLQJ3czFtw11qCyAINzuhXpWEAyox3koT8sW5qC3PDzP1c26b5zCaeuF2nwk+v5uiaom94i
C8vcdcLum5tIMRNDLW9M+YGf58AZWSjRfxVJ0PTKhRfGCqwpsX51YxZjzUzmAQ4YXHFIkhTc+m+l
w+AYYa74OxtH9CNeGBSIQBBYU2PTZvMJSX22ILucf5f0wZpmuAMrpFiP4QtE2TziGYEgnyzNZ4Dv
drjJm8dcdwI1+1VYftRXcl/ngeXPOcEO+tb0vYteoDlH3RhcZsMLpyKuArrUaxGeBMYpd3zH9BcI
Eqftz0sEulnZMoH+EAIE5FidQbgaozwcfZ4708VZZBo1ngr1RwOfHBiU5zgGT1ikXyTB0lEkvOYW
h4EP0MjEwhabDOQiiQU/dHQvqM2Q9XpkNvOsru21bLP9H/buElofzjEbyPqQV6J0Nn4ctwRKjCZV
MbTz99G/AyJN3L6RdcxrRRn/rULstdfQjFOu9Q0GLPtuO584LAx2Vw4W95vpAmU35gFcbVVHUxad
+qeTWm5APtjHZN1ZaXLJU0VCLEJ0TToW+gr81fK9HdVtCaaUUcxLoQWXwkoCYw32tfk5zA0gHMqu
tm/TesvRct3ewa9G/p5OmfWXtdwzm0bZQ1BHtSPoFVQhFvbMUhQFHtBrSAzW1qKaXyuOYUY5OoHY
gpO+kuthyVF9uLGEfdcB6ja6d0UhhQVPwyZRopp5C2yfaOKjeQe0MpMPIl59z5O7Dr++63B/tZkV
01kL5cEPS3YaIq8kJ3ueMcV2dOqOfJH+BhW+j68VN9EWdcVDpQvoV0Kp8vza2B0l+RJNuQk63erR
a4X9fwr/BEVBzVfd53gMu14SPmMI7urFNdMhLxaryeIlZVNSO7QmQKKrwBHsQtkJ7LgLK8joczWg
H7Lg6IKnMKbPrQKXiAVlcggrt6okjcMcpKdjFP+QXNcqIDYUxB9Skha/PzCw9EB108oWLjbzOF7K
h3KiXh27ekc1rXBX0pQVYwf99S1UvcxEUFBRzoHtflxGQOoeE46gileskMXHC6sEFqst7ZuYguLf
oGg1zuT0dJ0mB4cIkj7yMpdJINdHQVH4H6AT4z6+BWKaacB5TUjYE/1Jg6XpnIOqICOJwLAG1KeS
3D674qKqrQ0D4GTPjH1IZRvC2rcgHoh/u3gVgYggxWPXZ1hiwlqZ2QlADOgrOGzgEvAmgj8qNsgy
Q//W5fLRNQlwHTKHak4epnnY+3X0ITfZepe2W96wwERuR9OhN/q9YNRQpdQWyVX2MQMnEZqjr/Zk
g42ykbCP6mARs4m8apPoQU86a198JIp5TC4+I0Jzgzd2pqlOmm+hCSZiBpklrIwrHpNEvSdtkng2
d9w079+H/YqOQzBMvQto2lR6Kjmuj97+cBsRpmEGnWAyTKakhMBm8Vk5HyTbH2RKVKcSnn4I0VSX
ykD2ab5hRkVcLMvf5RRCg5WZqVAeKyz7myAJUDxEP+onjv52OJT13wQh9tQ4ay8Zc+KuKRTZS3cG
dShTfsSrMiyV6wTZKkbwGjz7GmNJL+hqfwntbW43rLm/vh6wmvTgY3gStGcvxbxl9NKul+0BPMt6
HsT3UcKrtOO0JQsav7HkgjcfNgju8CfwCFSBDalzKP2LpppB0lW8z6g/vcApwIPDLDDrPAZoIryf
D0MZFEeDC+COaFB3ERhMcHVUJPHagd6J5WhXmvTPBkXZHZKce6V4rIiDKxto2Sm6/peuLdxbzbTP
tpDfuIKFaQLzoUdjWtJe7mq4hcWd33iwM0OsV+E5eNPNg3uMv6UZBX2IYYOtPd0OmiIkdYNgXhs3
3k+0ZatkzHq8vmsAt8s1rkAVg5PzljEsfVF1WPl4EO7vYS5qmOv9kEr/LpCNv6s6CCuyxRdqC9uM
o2f7Cq5vibZuu3jLgDmXEBepEJyIvegB0R+CRddY3eMvU46a6HhOeQyR19aL4pbYJhdeRJ2tq+fN
/BW33/CSjl7ylI/7ZXHoTa0zZ5F7buiAp0tYMlA+X1bb+37J1Siss3HyHfjqWwTun4Y9D/TwkXGd
7EV1m9PBtMx4MtlIJSKl7z0x9QVMTuNNyZ3rVKrMiO+XXLNpTDarIBCyvT+ICZJH3BdbDH4zqwKt
nki/UOw1BsQ3OePXf7D/w1QUiexR5Mw3lKD3VAozPkjnr+8qr8CfNh3aAgljP+4difVwGluXf5p1
T7PYhEPBy7EBneH3G6DNRcRloCpQkIsl92RxZNjZ3g/fiAyZWedhFmlDUAUxwFeFT8Q88lTWJDMx
1wAHaptZz8KXH22RYCq8/b5fZgjr9b0qt13IdK7yA+TGNy0sVKUhK0P42M3XVosLRWMev5Zvs/er
cu+hmCF/1jvcNV9BEkfy8lLGgdLPqOME6tZ1kQunmDHm7dmXs+QRRXLMIDBps7L0LBAVbA3sQJ1d
u//fFiFcyZuDXD/hTG3EnLBGCYRBgbc78dhI2H/GqKCLn35Z1mc6cdJTOk8NIoqcAaamt206V2Qo
aFoa5d1xw+zGcnNFsV1R5WR0INC4NeTaIDcjMgZDcBYt1PLkJe5MKXxEoia39JyKL+MnrmUfiI4M
KEHXqfy6nq/Mr+hxRPtxfL5tu6REY69wRSm8+wZk9wGtjMp1ecX9xWaLxjFamOJjtv8XkQX81l5y
Whcbrn1ytkdIyzI1u5mo4SQPDQloDJCC6y7+Fefs20BnnQLW80eJ4/1ABb/JfKam11/IG4JYQE9Y
YstBPpbxZiNigdhusRsttktXDNGEmS5t5oO5GBzGEhvmMs+us0Aujpx4TnDkTNb8b8lwYWNqetzm
fb6fUCeEmTuEuTXXkEsq+eXIdHWAztjUxj/qJpI/FufNqHmhEN6ce40t9kV9Uf03MZvdpcrt23Ql
XLWj7cYLhaIzdcl7aNWjU7+iO2NGIKWpq2/MZWfJXzfBnf0fuL7ITBpvkYTkpqBKlff5AJHpgbXW
ooylGAikXykLwgiBKIrCxfO9CWE7FVXmsx7WfAJ5xUmxA95YR6iqbUsaHs/8ar3LXxK4W0iVM+qR
V7HkJug18xQMGKTVA+eQlzHQa889H0c8ClQolrEJB7CvqB+A+SL0opQlQIcl6JFdvsBUz9hXyO+Z
yxkecvLlWYGAWofWf19NO5ea7YQw+yFGDV34yrzhHd/uEQIxExdFOuQVLQBgAAD4dvz9rPVxv1cD
8D+iP+MPmdWY1Vk51Z4vqWKDjeRMQkQoYEar5cSAEduur4tOFyflI1XU6CKNjl0/Rp7p9F5tWVft
uyUw7+pQzt0PmLfWx8/Pp+TB3LqwgcRfksfANVcgNrkKn74+E9FCVNQhDcQXP7rT3nveIflc1L8v
hdxPCq8u3KvVNEs7QM24Gu6iqCvVfT77KqkmAIYwaBEgg41KyBwdU4TQxyQPhp5grcxhbUN/LAiH
qMDYmCqtauGNr1v7QvgA1h93StwHxDX2jnXYnsO4XrComm2gOP7PWAjbLkGJI64YxdqVhIxVppA5
FnkNnomlz3vI352r0Chp6XVhqqeSgJM4JvhW0Fx9ipgX7uffWegCTCAsN6c6y9woZmxnO7wL+QZ4
9ur31LuBQUkBorcHeka5FumLQXWZl4oDVazB6XOFyc0vs4yAPdBHkqjmLeDJXxid6hRfdwe0SWrU
lse8MmUChhqK8E+8O9YwzemDo5gTdIil7XghrhachtrGZXDOkHacd2yjR8Vx/PbQQRnfFnnCEVki
slW0JztidHBMmVfzmbCC3w4+VnEzzi1F79RCxzZxyV1EbnlQYtOZl7goAHfp1mKGdvmNTTQNtau6
qZ8BIzJmWk1EFaxm3ZyypCMvAQKUxFG9REjGZ2MWAi3Nbqpaaiyee35ZAKGfE4dANsWDYKyfP5AD
E36vMg9DUOmFxzDyuyrfMzHyp+bXNCz5ej+NpU4xn3QJ/wPkGPPE6saWEFeul/3UlggnGrAxIPz1
7PJdf6cUIRDmOHZpPd5yNBveAk8gf1CDMToBVCdlFeoQgow8PF+6QUiRrB9d/iKD9T7epSa60Ex/
TQFLTX01mMD6I+exDddKJAM1fDA2vGLRkE5TjcX81nSgQ5NUmPl4pnldS2h/FNU3xZ3cUDtB7Urv
klOEsgkAz4QSeTroJmL2d4XeaOxgGdxn/FFYiKMKf3ZO8N9OdIFuZMtCCb0Ne2g1Rizni+1JokNy
bLOHm4QTBrGYJiv4FxGoPu3OiMrEsouzlFfhTXLt8iiMlzMLAAIgQ8aNE2vC1kZUbtsqgizYMJFA
l+hVOvjy8WA6hNGNwnWpLtvmR9vYWAJGyZDVBf6Tyf9DyyIdR5hEoomDj3dKPNnrCM4Y6daUk+RY
3Inoy+JNyT+Eie0Qgd/3s5NCXvROyGISJvnMd72xuyaVJieHVj/UBSISeGwcAqCYebLi/WF2g0/Y
l7mAuAuYVIe9Ie9TJbOtzIbmoAZdTvVHd/Q/2PSaJOP7z7iwcconBRTZmNjJqoAglBzz6KipMVav
p1z1eC/SbULrocZ1oKmvRwgIkv3l6iOyWs94KwoTmMHJAxQeueklAdSNzpo/R99THHJj/rQ/U0Yd
bW+/wIL9GDv/5btdYiOEDz8E5xdFaBl+eG8QOBJF/J8d8zyiNWzXtUquZyDesleFkr1ZulXyw4ZI
YRHmBpCzadKVTH7q9iy2y6KRwhS/yLkvN/1AWpSXJ7Q/0ZR15B7xrGBDcZdF8UahfsUdjqknGWmP
HYPn0yAbrYIzX4XYbE1AO6xnd9iR5PBLiSG9e1dpWx5BkQMnZodOmsEKYwUDUMQQ6DUnMMbXKgvA
UgcwhdtftuD13PEzDdXGDueSpLXklPU+//Rr275AVjHTT4ldZFUf5LDist3FUcO0PE2ywnp56aN4
uT2KQsDFNNPB1zEyO01baCowyVaGvXAOxEulCWluRTTFyKcwDj+qeCxFJEi2AZI/7EEAn4ve6+4u
3Iw0he2Oyec4KX7z+c4CgOgrp76Wl5zkAD6gtrkV35U2sZgUAeyhi9GHl9Cc2mn7mR+r5lpCSEUP
3Ys22lHhCh6fPbkSOGcin+8YKuztrsrBOSJfVk3CXqz4eHDJZZwLGAPV4mxpRTSUYmmHviNeCuhj
pwftQk+cLe78PWcbcMFK8k4Fua+iMgBOoeDlx97zkQax7ACaDt3FrDgN/CgBA8gPZdL0UU+VM2i/
S1DyluSAlPbB1aYoxDkyiQ83U1h0xz5n1+8bjvhewy+4t/i1jHe3zISg8Q8qTJFBCjeyHSgHbv2+
jwBMZP68YrCwVh/Vx/DYOuoAnBeKaOSH+VXGr3QfmT9G/PFC0v4oHi+4cM7/zloNJcVOS8DOPfcT
dO4KpbxjKw+Lo2klHX46jMqVmfXv/8geGoUvQ5lUNR6XdZKDwM9aUVDCFoNSQy51lE4tAAItLwDr
ts3JCshgRQSZmggFRcXh8Hi34B/zLDjrt/9+uaTr+KQvZ+2S/az87XsTLyigOTrbd+WQowV4hKjP
ymdcaFekgvOiriEtR5iBt9drvnJ769uCAk7fnFvkkzTCzve1RQCg08eg/ZHYXOcm5jRhSxonawlR
uPFGH1ZunA56jImZsV1+7FIPVxr5qAfZb4n3tIHzOTxIZ29fpl5FjO9tVeKQpDZWu21ovtbSaFCZ
3Vbys2FYRQ30Nz1zZTg/CcSju54r6jZy/b+yPne9rqOf81TP5Ll0WXCdsyiCnZXFeCJHcLhHPenE
+/36E8d/LMuvB0jRpvIVl/WLarRsIK2ilVLLRjrmbEQAYFUbIHmSO/w/ssXLe7AhlKQVBCpVvf+U
REQD21+R5OaOAB/RP3uwZsJ5v3h6LkwqZftN8zdaFhKbrPcB6TG7dL0tUSqtaniTIkwnU/2CvAWO
unEhOAtuQmoVyibi3kdrJK6dxivec9GolXF7zaFZbOhmLIjQ5yMR6YL2jHBc2HC1YVhr5AjT5c9y
oQbnwtOwqjE01WsRaBLIhoiPKeNzeRFRM0hOOV+RF27bTcGJu7Z9HgXmJY/wbztGk4FzYws1wRJF
20YnSv8i/uDYRImN3PPEfHOdaz3V12PUIS9yf4zH7ZZnJhAZLhYujrXww7uU3G0FGQXqxxpEgTBP
t8JPInwMhBIpTZOl78iAtoTJKqo1mL+fKEQshuGyMvYfuUjejGc8WnYDGGKPBB+8sV8CG8sxywnx
kx74Rk+cjfAtnGSoclJM7qTKhlG+qpuYjGDSbCnFa0gEIq+x9oed/3NW3UWKOfNG0J2IxPShqgZ/
6LRrK6SU7HYOUtw+YJ5hn/urNxFEFJ+Hjw8ngmo9jADTqP72ulHI+1W9gwI9a7k4fA7mlML8WGCX
VUYXf9xb/dd+CRFm3PDCzcDM3toOz+Ty6fWlsI5FSXV3DUO6PgbdURHzjSakEHbvshOyDqrSNol6
AJJNhQmEXzsQ1EoHYEUg8u6H2Meb0HSTBkRwmt0silBR2IwcBhmSeqag1ND7pnjClpdPlCtKTPf0
RyyHkbOSdMmt9JuyXv151X6pb0mq+w5OX4iW0oHY6qYCpm57bUM2WxaukUdXwFW8v7CEV2oOJQlj
pz8TIfeFuEm3GKVDz3MdY6xbTLvmhH9A6pA2txyRv2sQ+ZETw+vpOL9Qz9WkqUVUszpRPVDUaJX9
CsqagwO4sNXeYq1kpO/A5OjSeJB6ENXXX+RvG2EnoZ75R047SXAlAptdJESXbsya8v5NL58VpWkr
wsa00c3SU3/pufT+KtgeEDaxkxZB8n08+7Y+RWVZlbCzX3NDBK3PdLOWVvNlFkiR5SgsnfTewsJY
HH6WP4bVWVCcU9kNseAdHnUgOIjCIj5zphin2xmxLnZtUMDAO5lrXScBEs3I5XINZ5Aaqcps/dXL
/qbE1UMCPXXR7cVUSL5mAvGNDSiU0oNOZGuj8G4mzL9DmN4isBIpzqnHdc4zepCxcivmz2Myslk6
bZl7CyF3VVDtRFXLTBvITsmbBQgaye5gv0jToC65GdoP6S/AVNJM5QIn/8JmkxoHLLc0CvOsYIpH
B0V6zK0Esjo/NAPV+sTRfFKcD2zoXDgKePwaUMDM10AF6zCzqgyYfbwZEv5GGeIEGb4vbhRuaBlE
thK2D8u8kfR3e43K5QfdSTzFdqJAZRHbAIPUtpuRRb1i0N+1aDvtp7P53vWclyK5JeuHlCmGWM67
pUoenahlVmKqQzx6aHN0wPhgCLX+EQUaKv5OAOj+n9KBFRj3ngaK9EihVHCXA1CxoLCsFKDV/Cu7
oV7/dKfl9tWKzmWqdzB/0nrdtpgSg7LP3ARvj3OoWBpRWco+dgCkEMyOWpKFOau6ekOSOXAPOYQB
gsxil6trSPytBwn2KuPQuAklE806N/i9BW74YVwvGpcn6/CuTp7iRzOmAkIiuQ6psExNijDweKEv
Qvx60w2iTKMdEnfkCgWsOyTqfynHcr6pkzskVlvXXl4m9F18YZ6K9Xk6xHoCberRlwfDGPqQt0oZ
XD3OVBmBVhlPaq67TOaEny5hD03RLOk2pLhaY23y2MEoa5nHYrfpfoDNscMC7deyREhkTTT8JOGX
xjRt3tKeyShRH02StvjOIeBUvYXcLT+amNDyqyTKAqkW7YnleAp0cZzGgZ0Kbp0omJfsHt0BQXoD
kOUpojSr4Rx/34wyI3ZGtp0fkNMOmETfnuGGt/2tRua7uMobhHlZWbduRpRg0RRdLtacP82e905L
ENRqE8ABAw4hb7hE3gmF//I6LxJAYVdD/p5CeZfX1dO34N9hQ+JYDdy26Nzsiv1Mu/ZVF4uF/CtO
UPZzrYHjt8ajGcvNewfppA3jJa5VNhBO6mPe/duKe/UHLs1UpGBfIf/PHUIk4pebdDJX5sJ6zJKT
Zgk5zQUavcFUCMxOWhFSaovruZ0kLoyKxBphEKY7L1AKstngjNTLPWuJ24pCAQ3V5rg6h+jYXiLv
L5xTdOrBq+EvNWAoA8AHzSLvb5Ooebak9y7QQXfZBQ5qdIyBIe/EMm0wc1E2HdiXdZxUjY9Mu9O4
YCpssbE2bEsN11/yU4SujqcH8yXKjJ+/RhpmtkzPDfGAUSKKHojiKhgNP5bAVxcm+abYUsQ4Epvt
iF9Ejfvcm4FvveWGG7XKyq3sSdc+QnaBiHxHSlkXSzOZTArEvvmnN1O25JxoufolOriNySuwqQH7
kompypo8flquzBtIoMAG+eMyZaciqHAdE/BYHAOhaxX66jVwJPDDT3LQdMMAiAfLY2raMaB/8gqq
l2pWVXlZ+jz9NxlN6Ba4B+vR0cM8EAr+hpaFG+CwPAZQ1b0fvYimI7lbK7ONAMrtVZBZnKSngQUT
Rh5N3il2x0ydazAk3C44VD2xX2pEtokR2RTVGfTgMweOu1uXXATBsLQsDUFidp6pvFCB5vkonh9t
Iewv1LX558Mq7rGeebk/EXjYQVyQ3sDaAv22FcCOZdoDlP6UGzx27f/kbEaxaC8hZucgqpEO7G+1
goRVW9JBGQgg1c3C9dZtz1Oo2vcFV6ZmmQDRL5ehqoMSxVpAIpKyiqP9K/q7hQODIGSUIMqAfnf3
PUp8n9iIH3XoGssI5gEMQxn3r4qVsL8q1/cs8JRiN4MDLO0kO3aWWt+vR4eDZYYhxKdYuFGpE8CE
sgB8frtZOrWmp06sw5t0OJbSfuX7+Yy6CxcBShghAbfqtvRxk40JfmAE4K6icNiKaB7ZLqeL8YcI
crTXnIHL2hhdCWzfMqw7nRZxZtb0ldh9j+hsDVsUkLxAXorsWL7j5Zcea3dJX4z7s5yX6tDcSV2s
x5u7PearCk0rfEZxhH8GnkeoFLKfWowoNlkGxZiz5D8bdo0d3+f53xcQLbyhZd85OfnhIAQsxRqN
RikKO3/ZLXo3HyLgzEFw/NaNmg2uIibcTri0EslYtVCb4GoKdJ2ZeoDlbYVNu0VJQjhcGN2r/QKV
EZttuNsHLgQ3XUcKQhtjgJPuKrH7kuwLD0R1RYRKXIb+pFej0jK14wHTRPqiC8CIPbiD3TRNIfLq
G1oza9bdfIHrm/gXkx08ck6lYOSGCT2nKqssliStJJVwRQ11iFe2WBu/RlsKnEZzCnmSN1XsZq/6
dyPqEuq4g9zkOkBtnRJc2Z1TcRtKj1LCZwRXT9AUR1Rw/hI66JcvhhIF+FXcHTNWSwsxHRgqRtZc
trI3o0jY/ZFF4IySEigtHs/XTv8kpgKLvRoDTYiUdLZNJmP5jIrEBmtk/gs8fnz9GUOII9HasTdJ
bXnULfLbz0Zpa1Gq1AI7zMM+uaoHnAPC5D6YnuDo1FYlnchZm5Bi+B4A49uXedvC+UD77Zli82ty
XstZtzR7TmjrdrtxfysB5fo9H9DFZYZu6t+T7BdE0p1OjPtY4B3HpSEAiZnXD9nfKYCrrtttgcIo
EiD2ND0wHAax7vE0DqLRQQ7AfxPNdk/s5DeLSh+mXGKTovJvWbw6a3pczIuRF5xYQWQCB5if3TSx
o4KTGM/m2u5qkv5jM2BGeGjpl3ukR+ZwVQKDRMR91YqqLLOeWMrplIFczDuO+tOSZU/yxoc3X72H
xYxJ08ZYrKUSWr5sglEyVu/yB4jmfm3Lh8CT9zkXeJiHid3ULEYewyKAXcBAWgN2e/yx9p8TDtnV
5rEcb16iGBWXEYBK8JslTqi2dSbJg3v8LSt8C8zQurD6yuKV4W4N2Zpxn4yly/JDJSO7ZirPvNk+
nxM1iBeo9PB7ibajmg5OBXPpWjjFYWjx1wNFKdUfPrAtV63M8D2R9n926SZwsNZ6N3ZGXAMeIy74
QR+FN3pMYt6w1AJwZEK0cWbS9hJxlGUvpg5aXuwaTAgHVXpJoXyeCNmmM5pSsf8Ul88z1A0rXzYl
EYkfDAU4tVlqaRG29qPuWTxAdB0lueHhPmmE3of6YzX1jiIyt0vlCbUGS7fIzstjwu4NjP1XO6TU
Jorf6UD2f/3tUNkCfG8b/6nO/i+SEMZ9ZGii6zgs3B5HZfY2zzMeoqDu3xwHO79LuiugtZ/Q9C2Z
Z1UVekDk3VWB8lfr6towNFMeY0JDsX4DnP22wsZqqM1bg8YcNa5yVZ8j7PcSdzxWx6mj0YiMSsld
yRfYzvFo+0UL2bvBefOYLQRE+pD6j71X7IeesDvOfq4rF0TOa8x9B9wjPFxbbdh1lCbq+52Be5Dt
x07Yo5O9Lsp9EthHo56q/rSh5Hx9ixj9XIkiqCay7B6gGUnwvdCTe99dqOb7bjwPZhVZk3SF53ls
+Z6SBbll5PgH2BOFvyvvM8a8qRsCx3N6CUhVVbiGqvR7Ey7hIiEOPljazjxo/4Kor0PGDEXkVQ+z
TCtHksuXoGyY9/WmrgnlSg4h5bvhznNVEPn3jWMakljJ+t9qaO44bQZfcAAiEgDS3X/ShAQZ7Lzr
YG9r9OXLtU+TUKQmy+j7IuHvWb0RgP+QdrUgPiDRtHR8S43RQ6PoiY3Su33cvyIa4/gXRJsmENRj
/GgXeJyqXRqfPWNO58mIIhgPDL9c3Pj8usBqlJeaIdtpKBGjxrR3jOWjOnn6dyrVeW8KYLTxSwct
MRbkhgfnqXTpxiEjdWbFe4xCIudL8KCLBFVX2UB5H6TP9cYavyPyV2tdzKGm27m0oMVsLI9d/dCL
iUhXDaA9A6+4uIVk/s3+Q5K8hXUn0wlvyqP0nGT63kfqocDN8bd+phmcUAVPIIBgPrHyIJUazMGe
mjyv3/XXFEDOhArHcNBlmiPsNYClBDPY3TcsK2SlR6YETh3Jg7atBBV/ps5owx8HkGIXzEJ2Q2EK
uo5mVG3UgEJD+zoZ1xykW7bllSF+5m4DXRTgkG+hks8upaapIILopFCo1fFZKRyyZLSwfT1J/ri8
RxhUjlcD3mhzjwAtybjBmRXl6oaU1zloJFz1rvLxTTfptB+WJYH6McB4oJeaicsO4qamKCjf8ty9
caWa/iLNYKWLENtb1V1OWBoHch7PSFd/karIMy5hVBfWqX3GmanMe+otY1gKvZxKJs3NCtA9aBHF
WMkTEq/clwy5D6sqeni2uXokejHs+YuDo1YmC3xMhLgwrvhgtn6oTQdRRPburmlTjKllBXNu8PFl
ffnTlDOTt+3AUx7Bvf0LoerUPfdy5KclJh522zFZ8UtgpG0lFB7zpWJ3380D8vgMqH55iQGkd0Qe
2dHMu/gV+8RbrtM5bvtF+VImSfAGY6xK8O1i2Wiw7CZQrpxfLI1WZ1J0aZVRiI+dnFsMvXxi5141
5nhrAJZ4ZbF8UbUCdgTKOIMHK3K7jCXOLfco3UigyWkN7g4kUt1oC6ck922NKUwh/0x+SDbANaYi
GJKHm3C9Vs9xPFUu08JeDrIiuL8FYIytSHj+4PzwUtcnRKkpaTqqULVLfIM4VIVVEojWtxG66rtl
c1IrpLR6Z2u8RehoHukyejrwS2d/pER7EkULUt3+kjRFD0+LDFXIkQy8TAnwoxMY9KTRRanTGKsY
TDRnrgt2kuvljOX9Mgj1/no9bU86kauRbd+mkeskzrBOKOajQCpAiXTnfBOAEmiq1rhc77aKxi58
jvjPvYfLWMekgSG4mJAirHM9OuS8CZaqYNp9gG9zUBSMnHhMqMsY3/xG/bF9Fkf9GTFpmJb7ThXI
vAs5wDyKlT9wjCw+f9u/oTbXpqfNpFlYgvuYdEBjWjg79MD7knvo0WKTRP1qlZK6R0VVofbu71LR
kPWZkX2LfTTc4rZ5OKddLJWhmXbYbE2/515+ZVV0Um73BB3hbKAkj+VqA4rMZH82Ni/pDhUmN74L
t6o7nAULSMGxmFFImLdnRVbzqK8of65OPQ9jGOtwWsn7NciAt1rr5fXcfVPVCw0AIp35jQG47LHL
KS2nYIHl8ogBcncCCHIR+4jBCo+HMEXHWl3DcFip46pZfIKF8Np7fo7+1D+MESRvPDwj2CuXxQiv
VITbYnaUY3I4TbauyQHqEH1foxcFkebUXH5lJ4Pj3r/FUUCqlmAWmVN3gYPWq8+arGYyteoEfimd
CqLMw+3ZBIUoswaAMnnecYyImltcqEb4CXJQxyjieLpRq6T5YkhK6GyBhbtPP30M9Rewm94HKsX0
IUPFllZnolFYV8dEQHq2IABsNXlbzpbEs269B3wKBUcHiicG0didgvzYl4KUr0/IZJSBR3C+d+xk
pqpO9mCoH3zemLW8dMxi5Gf8d2//XRTVOQO12rp2ki64aVQpSR/GscQFJQnuJat6WmJJOh3fkKo9
ezdHHXZXpUMV9THNtt2S+KSt6/35oCVZpDp0w4POMgOKlT++w/xRr+Ig65POSTl/Ymz/zdFQbI6u
PBIEAbGXPcQvSLv+kPJ4AQcAY747W6jL9NQk7tZfIwaJ7P5CiJYZfHvHjv6gBFK94UafbOU+Wdq8
cYn1/KFsBYb84jT07564mJhzl47FmvZLg815Q/2wkpco/b1/25o6JnrjNX6/FFiOQUl1gy9/BZvF
W5fZM84GaMY8SsNGCEOcfptJWmG7JSrjD1WcJs4PwZZhaOoD5972N/aOLnCbU0cXqZxRVhMaHIJG
1nLRbIots82ZgZePMJdIFi64tpQc6prHxWfUmY1/ycP4ZIHRzqMWNDxJOy8bg+fP+rEpPcre614V
AqUCLa9ktDztdLqWvKsJoyjbUXnZIEM76icSkiT1tAvHKZqM+D5zldENOTgRTaG9J/je4YFbq0Ur
GYzbooCfNC6CoTc5M0AKF0r166BqQO6ZIHRZdCRfgaLRvYPfctG9aj+fjj1hal7IMbbW1KBpYj/h
GUV+a4L1KcC1wubbINGHPfGnkwboQSZDoeu2wFump9vtuqEsAlR9glWnAT78g9ucH+GPSXaCdh8z
/N0O4tt9j5FQrsR1mpaYIzOBu/tGtFtBwy+BMR8T60+b3SNQJ21+eDmLlM/eJShwr9JLYjQy0qN8
NL3yG8yHEXRq+DP5F3+ohvgWG2oHg0UPQJwH+FjN1FlFModr1fr9cxf1vkOxk8HL/aJllPVNOEZW
wiDH5RMOWYfoJ3KiyitM1yRm4A2Zxk63+4nC8q794gLCZ7Wu5mFYI7746F5rT7cUx+3M9LUOsV8g
BEPNE7PgbXLjUiB6wJxcoZIzyhR0sMFn2gUwDPqmrDP4tbOHAotgW2zcOob/G38mk8WywA/lB2EO
+ziZmKz5dLFDiH79k9oSy5zYun1Wll3r8jyYRr9y1TyQrUkIs4z5pia3rc0dv0axH+Xz3edbLXZ+
z9ce4+vbgoFhcPYVWJHqPN0bDqzVT2IhDR8a9TeToaFWQinVW8iWqlC2jJKuDkkpELouYuBYLurj
EtX/q06rRrEywYDSaV/X/ZYmujlqCMrvMEmqy4M4hwcertcsOlZcwa7gyfAARZ5ubj8fRczfcKG/
IgYzMABlvpN/FTznl/eBy8a8pNPqpkMzXWKDxovfRepORlnEglY83CUc8/cJzMqBNF8CENb3pY/O
+LcTCTIl+9/TS4uV+Uaa+2839tKb6rS/aa1DIYDprcxOAlGuELcvnlZs9P7ck0g6RqEx8Sh6fh7Y
KU5QlF0SMqhK866lDzLKaaXtOS6+YWOLnLaVu4+OTvWVVLZkqs+eYNvHwVmRb1S2DG+rxSh8PWFP
PsIGYTpOfUw40mrgBz39E1T8zv6QBap2OMQTNS0YFFWUJAY73Rpd5iXS/2pOmc67/Rw34MwLBUpb
hjTkB1mJUYMVm46uqDOKxypkr9kCOKOkHus/wIkHMdU8Og3Ry7xNxq9sQESfMCO9BQ4yBa3ePmmh
tx0LDuU7OVPP2QRwE5kFsZj+9RsI2+n4ZAU/6rDSGXPt/s5o6PoJaUGKroGEaW7yqj2K3q1SHEZ9
3OPHpK/yJd5NH/38Y3i5wxt1LMYW24OrVXIYL4Wplxz0sxg/gSLAeXgbUhOF+JGk/yUzuG/uyJVR
vEwsaELjtvaclqqLRd/1WRasWaKVg0aBSFhNU5BJVN2ft+CV3/8tILbk/Wu0jKwqq6eFWuBMx8Wu
ZAmccI/0frwba3zDdwPmWMyBNgX09Xjz1uw7ZB7o8+CExdcBhF44VeIgp5yEBE9UQ9kX4C30YUVS
Ob6im2O+z6waMI8uM40DaXtd1MUMqJRJjgaus6IQ79EWOb8KWV51dr/DVgwD/avWet5N1ZBX93lA
/QHDD6qhE4aMCyBZQwdkZN41EG+1DPAtz3+5OW9ULn18kBqPFMQFC7HXWFVrOG3NF5HIbwuII+lX
S/lvKt+hYVRtlNVIWZ+E6qdQHZ3wc/RforkvlT3KCYy3qCO8Grja/XKVmwAaA2HzrMw1w8uCsIIZ
OxW+o2yxXr2CSERoF2s65X47mt858dr2Z/I7eEqY7caf3NJjdhySTMbKJGtX+GwBJU/2njeYTLhR
gv15puEq1Acygn8xPVtIcha3Pf/0Sr+mLTFlwdM5Y5SxW/Lc+/bKxoas17d1UoPag/e+OxNsN9PV
918JYvCJ7+B7JlN7YpeFj/yL7lRv1EqAx8o3B90tPir6kCapGxM6A78R3CxnFNyBMPMNwjjEmDks
Z/Aqk74mSVScecu3s3JLyeRSfKLhd+zbNdsvKWZCbJg+rrf/5P11fMhzSe66xto7QE9VeP45m2fz
4/+eCZVkRAqwuyN0HV4OyfVWhOGllGx6h0L+uPl/pHMX2slKpCR70GOvGygDQGlRlVxa62dK1HTU
lfOob/CKBir3uHuHQc0sXnfqxnGQ4hGc9HpwXx7tp6wnZQprZkhktxE9g5n3dlchy/mf7LGXufb4
aXls+QTmwXYwJcy8Y7U1OXflPVt4gpqYGam+gZODZMy7MxOd8RgRGluXQFy3IYCe1pFii9C9EqFd
tSnCAcaYhxMehxKwFwPBaEhGEWuHKyVSrtazpUrbFDwiWpHYnztniD/tcJtbQfLMYnqhJq3heZQ2
GwERtW93tcm/zKujLTJeUuCpJKvjCsfFHp3DjSsvLKn3uzW06VByDwLaNZCMQlvIdCvjG5ZPUZ4i
WMHc57v0T+Z3+dGtEJEti87dBW7r/dhuTlp3Ir1AdQH/ac7WCvT9nAvITrvC/aeTfLNAJs2sJiuQ
JafKEk6wMOp+nwQPefIK/1djxjuKyagJ8IC6w/6P3YQHSE6ixd80VisGR1vD5Nx5El6pocHhoc6y
RAI3vpocu/jtNdvBO2+P7ZK4ZMX6T6z0P5CVFkZ2WUy19mb3M63D0Gmq7n66ZW01SRYBsCuuHyiA
0Bu/hc5GAk2O+IliOszMB4G8OLOAwlYk+Z/NuySBXa1A3xcp1GUar+Uz3x/6UtMMCmTQaLdv9xLd
FBWdykXEPLs15eAt0ArVyBErz177Gnr5qnkLAGr3GMvz2jNAayMWvT9Sn1u6hh+3iE7kJQ3ZG+BI
YDtsGHduYKTjiKERJ4QOfFA8usocva9gTblxx+7gtggMs+3GTtTNSjnwGZj68u23sJ5FwxcKJaT5
6dIukbdkS1tJI3huJt7/48UJETMQeE0ukgRrSu8RkV2Mr1RZeoejzC23y/IcYiuZCP4KVtgW39lD
5YIRzM+hgQE56+53d1rtuTcGoXMDkIhR7OKCpD9p6OSKBBsxYtl2fbVqgtuk/k5gajscdAo5s5jS
TxhqB/nflO5Lw5rNpAkT7ArrzmLQ9mftUK+xdaY7fOz9/kfBkXTarfZXBxGm4nHIrQYkAtjWt7EQ
+CJNqhMmKdlKIdU5AnaH6Qv96VBIfBVlXqbfvJtJ+I7m7mHeKIzEp0CuVAyr1bAspuZ3MRFbKJzu
oflk+4jJnXwU3r68yrLF6QL9Ds7gQMLibsASuA7EMz9B8KEb0kX4xsLIWOMKuSLUkV2tfTFV93/M
KTt6yJpk6v6elDlQCetPyY3zn1K3S1CPiLw4Pfi7b+qO47OOCpCBNWzrssDE4Ws2knDaqo4RSwWK
7Dfx9XqIKrw9L1GFXANOrl9Kt6E7HTsx4nyXeCgoxiea+jku2n/fAIVV8EhCwtna/bQWsE2kNK4j
CxgcRDUwjAnyq0WyJYK1fvXyT3UQ5/VPV077ykqI7lZCh1ZZe2d03afFVCpc+qHKVAF/xG9aRpsb
YWJZeFGi3MPHZatsOrlj3kwu1IuW5B+PmX//Wn/TMmDwqPaeko/RvNEKM0G7D0DwwrprQr/zTo8b
2x0lXCGIAyMkhhxHCRwiI7HpUpmBmVSpmTXJulzHJrjg8j0RqXZxC3gqmZscKuwsYBNoidZED72f
1BxOTOpFn9UJNFv0FzzZpMmVHwesphnG1ZC5vMg9/SbOS0qKobrAmapJY4zXNyDK57WR9oo5pPog
pCUmxbOENtpSMR6d7o6aj1iQnYek7L2KX/NUgik8zmI9sIpBmjchv6GDYj9gGzdvsP9nPalhr66X
/n1Gfp9oKkfOrAOBqTFbGZ20UAWlJ2NWFSC+F9bvHzKNYZYFkyIzEIG+opamQ/Ib8UP8PQdzwrG1
RFRA9AHDMgZ5sY9iiS9sZLBdoIqElPmYI9E6S41+dJ2KNQW7Earvc/wPnTCFHc/gf5JzkJ4BYa47
sq5euNm663OgFpDrxoGzTm/cE4IpHOh/Qy3TwyWde71fzlRcBaHmY636u/aEXeDzKa/T2VzEuDZz
aWPYKbjQ0b1e1eZivMbR0kJlF8SHxB9xlFPARuOAGp4mn5ynyzpLDxGOLzQMXMbJSBA4aNieaJRC
qbq8pq2XYr97jlOcq5A3SkBxiZ8IOg+YxcP3HDb2DGnZ8AzJgcuzMg6pKtDbKFqsHjMhnbnOPQgL
YZe8B+gU/5ulXb1/3cVo0Oc8Kfu+ympNiyHY5ZGFSANZ+fD6vNS+6SFCyBLaNCtoV1/5eTH11+DZ
sAbiL5XK3fXTmymf0YxMtsrhjt7JqIFSAK+4xcYadfxbobDKaQ43mSTgtxj05tnq1z2w/KjY1+Ai
fM2i8lCRbP++Wl0uSUUsAWvm1eOiKSnnWZyPdFBTG5oYE7H+kb7DYPrSsnP/cRnFtOvjDfW+hJy5
PtHqx8oCYDhbrBPiVFjCzf+uF5tjKpaHNeklE5lBY6/74QU9AOWJ9aeVys1nvTDm5D3+twKTGT3c
X9agYJ3vtsMBvXHb8hCa24j2+9YxeD+0L/LBP0pUS7bh7fzi4iDZl89FbwqKhq0hNU6oXihCk0Mt
9XFSdYwLuCUKjMFfsOWn/nmDAfdA7qr/It03vwF+hWu6108mKYwDbtFM++kfBfsrHkYZeaaD4mbG
QUXv0zJ99wtbGOTQGVJZNdsaOIBhUEwZ2MAzGkcYsGCAfJCzX0I8riW41sd7RXcoIBt6H5my0Q2V
2kRoMEwxxHz+OYpJt3q2JZ5iaM9geHuWu3KLySx/2U6c3Dgbr4VUWglN9hqa/4E6jxSx9/JSXezF
nG0ww594ixG9SG4bAEJuCEBI8D4oRCVfPvmQsoNig12W6SIHF7Jfotka4y24pY8WBnC0F0rRLsut
ZfJOFuq5AGFxoA3zHYM1zZy49HppNbBEwKglIczZPwu4SOhzeFaNqmqXb2g0eLt2DrIfmy+IYL7/
5RWmOnZQRBOpLR2K3cCR5/lquvh8srvoCz8tY9VHN9P/xBWtIpe3fhBrAee7l8r5nQsyJDK85oTB
3hg5kwYozXiNjExxwArqtWNjirxyNphWdPs39nZGZJ91rL+GY2yMdyYCk9sbeSDWeRaB3lk/kbul
bW7swOe3LcOqW9PmRV2pYlARtGuq+TQu6vAMVa2hQIww0wyLe0B9zigjqhCJRk/nr4mDCIANVr/u
Y39v/CmpOq/GAlFSjs/itDFOxpjKnnA31OGzmmbw+t788T+ie8tLaDw0Ssb9RzcMcbhXVfwlK0wn
Mpp6mBk0Q0vt0JmadXv2r6yp46GTVeXx6evPCgH3IdMHbfa8q/65w8zwR3+Kdttz0wXtoPk93NUX
yGMuDnvxVCcEapaO+gYsbf23I5BDgnytgwj0ivNCfHxW4Qu/mgBLMJJ/ivXMT2u3unisu2GzNFWw
5ARItIjsKMqGnBI1Ri1gizZ55gT4TEOaftQESYUxaqG5kuAExJORRo90RMzZ8O+WqZ1YD9+ZqmUS
qEVmnJaNNaRz4FRVpN4M+rkvUd0rV5SRCLKTHbqC/zv6iFZM9Sv41zHAWJmVE3/VxJ5EfNoNVOC/
0lyvjgpkRtyBpdqTK84biwPxjeO0c1NGaXn0KLyk8NtlBMNukegoaPIAke/Di9JNRMr0Sb2z7vkM
Y6OurLkg0XaX2tSHY9dnm+Mbj3u8n5n0F6CJDx64E8OOE4i9Pw+pQfj+oN6hxyzlTsZUSAE6ZUGp
+M7pOSK1+b48o5yD0or2O0/FUk339R5+f2/cpspO9xgqOO6Fer0G5ruxwd2XTefUl/wfK4DO0bS8
8AYT9gOUulhwR07LnlrM++UswtlDJg/jbp5bIoroREvt5wgYrqATwQijQyhYv8x1PoZXS4MktdkJ
3gSATqqegrPCSRHq6Pwl+R8C+nmNj9lUL8E5djArdmonqW4JzUOt1k1Cyj5AdhFk8rhj8JxVYuI2
P1jXqCFbqxZVAasxXApAX0jtcxce2wnSb2N1gwxo4cwmntl8+o9ehSNYIWGKHxmsMpqXPpwFcqUx
i7smygze/M6kC80RjArmZo5kGPQ9fNEXLwm0ye7VsAI9vJEJvVui7ognIpWQO526RYIX8grofApf
cEN+eYBj8k8ZUukUKSTyllK4Ci7IoetCSeIsm+vneAgC4dNnlkOQ8yZNkdhh2N3Ir955VPgIHb4K
KUgnwj913iwCkcCWYL4Qj9XlQKYqmmOooZz2xMVTy534RVtDRJFHyNL5+BpDi0Av85U78y5EqEVz
whInFeOFzwOIgL7Okq2N2uBkl0V/3PU4r0KKpE5CBcvpTI388XvSCn2VWDiPTb1TbqsM32BcGN6e
cVEUxedyV9BDcH1TyERSaggbOfIzWolT+AGJhX9gHMPAPNpk7GfcUUECS5DkxkgfnO7OxhdUWb46
sHFbkzCElnvr2AsY/WZ9dqGO4Wok1tHn/8Frh90YQ3oK9APLlrfg0izQqH/dgpSYor5jWNsIYTil
UNDe2vu6L0itg9BPanXakinCCjpraBk+E3p7rxvyOPAGcEftUnjDdpd72MrMEMJ6Hdpd4PtuBwSx
wlw8NYRKFIXzNC7XxMi8JBkD+E0pSLGE3YNoEPRx5sB6kftRbBK2G9/+EiWFaEnGaWK9MuL2T+yn
Vzpfhw1LDNVHUnq9zmmLd7lbYP8hsnHhta+B3lWf+TZqkCZXDZKB2lf1qqso/J4R/3UTy7MEF90m
7JSKLqcAjEAMi2WjcmUrxIhIHLNZnzr7eqoFQ/hOaBshmo5HZ7YcqZknp8juE1CDo+z9G55Q9Sb1
fH7tImrJUmk9S+XAb8jWmDOzKAxw5BcQ32FSbnkxcqiFyE9Cr0xVlqCcmidkI9KgvqFJfzLyv2QA
XuvwRfc7M0gYCak7MnknJ/cuHdBtuG/xQlmSO251KATnLwAo913M0AwncHtg4vY7qvBfwz/ohE1O
TYI5tY8dFYtSTS6j63XVsaSyYxuMYg9gOnVJ1SYzS17cfnLNVbFga3CboL3Xsdb+QsRdnaogt/X/
SpAr74R6/9X2wjUiNquMJuf3TRdFcodDmD9a8QwN4kqFyShaXIzzMzIEIqK8BkLVk4Ma2VJL1Mve
kEB4dnIiZ3z+pTgnwSUZoXEZqKkjQmsD5ewY5ItRiXFnnqAV6OvvJHU2xA02QS96biEuP4xAX8MW
Rqm+ADsOMOKlGegpi6ACgOoCvibdoPx2cb4HiyTnW5w2oPCr3pVdQl3+mzv1nLQQPsOqXe0nKzEi
bDYisy+JNiNzQki9fVL45HJxPrERpssThUBPR3N5oMKajasZ9MEROnwVM18qZKepf6ipEiGdV9Wq
dwo8doXKKLdgyHaZRTqhsm51HaRqNSP1zV5IwgLVtmwyzpMIhC6dyKG861QJSpTJJW79DSxrd410
WlQE9Tav2OlNDtdge1MGHenb2fFGp25x+/WiK6c4dYVICAmO34VHMQuaKWy2p+/cDNK8w3LMaNn2
WohK4V8gQ2dl2o9D2bqGe57AbeY20Bvcx5GnObORPxE/6TOQIZJyYkCzKSlkcd9VIodABNYK4JEK
YP6Z876ytQ2WdduN6uSlBGDWZv977VheBajmaAuI/ghqieHBls4Cqn9gUcx4Xo51tE/E5P0pRSU7
Xqnyqeh6yHq5ofraIiuMGEL1zv48Jj1b4QTfGJJD8JQhuZOJ8QgVRltGTTg6xQtjb9Znyf240Omb
MLFJDPevQvc7q/7PqdjKOU6BHeZ04DcSdKYKVl+iMPX12XPVFHuQAV7mAtjmX/DnCGjIcNATfNEt
WfjQD3Dr4PMTlQDHxjoOZPtJ67itMHvyOD1B39moh/raTDHTK3UML7jkddP4EEeADThfrHJllDQl
Xvm/1RoRSRFy2otdXPH9N+gOTIBcQcfumKggZ4lWrdiBSs0MvB5nCbNm1i8lXs7U/7rTInoivII0
7n407vWacYvze2vZEnekKS944r+GS0oq28WHXPeLOL6ZlYSDK7+fCuDshkHfx/IZ4aIwsyuD7v39
NXlAtGJ8kNu0KX6SjrWTEfFhr9CqTxOQdMzCUAtf6H7jsOzgBLBsf8i1fvqC5bNaT6KqcfLZ0PZ8
m9HsmMWps6tIHCjVbEmeiATFyopxJm6iNqMP/sFauM+ypRvMkBG3nehCzSpfc6Jvy/aLh2XFvQPa
Vh7UpAJKGiMdBcVTBCbIScaNM5AQTiOMUbY1mA7+F+TojyzoV1iiyD5e0SO0YVimF+KMeEZvOsg8
T5SQPcTVJUyrcIqgX7h4w337NgE3/TxGJevvTDuh+vNLW1sU4lLiwPCk1yMZhgfRRCfgXEHGea39
D3B9SN7eZ6r9w0QYvFqXNeA/9ICRCWK6WXH1azIoK7tpHS+MKiXcAqoxCF3e0MoS2poi6dLdbIJi
sJTJsVq2L8nSNmL5oYlEvnKVLpih2F79bxJAjUJZobNmY4WtY+LDfm5ZQ1PPxB2VbxvJaNED8Ep4
DYveaY6Hz4YO16vL9QAbG1ngnQgQ1EwHbnDFdokzlxscIZ4sjaR182jvXURhQemmyXm/Lw/HcoDG
MqbgTTSlCY64d2jR+MAeepj7l31cyU6nEh2s2iIKfcuOS4csmA6CfZUQzo2OAHCKStXqBUMPYA4B
iyel9YbIquoG2t+4pzEsvT0sTOZnplASnjOLPqWenFVDXM/BITrqj4ZK1mqa2V+sbqOK+B8ItEJA
m0XchgvH4Uf4f513L/nRlCYJFaHayBHXw9APmu43fJS4Ysj8GX4yNspuLViA9X7e4vFY1mVyrEZE
uLdiYznnLj9uALe7jRgM/vOTRVEyUeo18S6H/v8DWE7rhzXAM31Ur6kajeZLVjWlibLEyjGKH0kC
86Kc6cx2LGcDMgJb9maE4nKR7xNrd85gY7ByQnGt605SR+QB8Y06XhE5gDAkC3zmumv+M/nT+Ajp
XbT+dozJ8cNv7aO6CKjgCTEuZLXBAqjHmnlW/70IkhqejnxorOGmEaM1rEwh9u7JMTFzHHxjdlzU
z9FZ7sofBaAYwCrQfb+yi4WkNKhmwCsUkO+lhRiFQRb14RomZMsdk7BMg/3Pby9xsQYAsrEGJmbw
wLAF973vNi7ar59/Z4KMS+gIW9UQudtwCW3781I2hiBGLjTP/QyETgYiIFkKY0WZpxQ3fN9NTn61
Yp5QQJWBFiPgfnK4maKfmz12q240v3YoK01pTOI+r/LWnxepdMjXpFVCGhFkAzKTI9uBfzNbjime
AigAYVBIyGPGAng/2BqRFjupeJwyua1qPaMwgv2PsmBYO0SF7O0W3KnWlwqnH3rGsAxrCd5IhlJh
60gT083dcrIZ0QMhCltXV7oENu0ELLpBfxMPcoWz1QbDeeXfsRltvAuJQuTVXwVtluVhxJHsKl3w
3Yvj1K+ePXRsjdsKXRTabZUzwdRCcEBMQeMsZJJhzzDh9fUIGdUJZYuE2Jtc7nBzJPHawZCrWCjN
2W9oikEK/UFnEwkTof2+g7k14pXsecE36Gd/u9HLcTnjiFMfR3BqAd4koM3b1rzS43gRxFxcsPVr
NTuvQ0CGgoQdGLiJNzBEPlYNi1HSr1HSM/fT7Exq5iiHlAxQirnxKsK6vXW0MzZh+R4Rti6F9lAi
HLHt7fCCLNqLbhVl5F8MKnzO3WpXlSWEcsxgv1B0lkQX4Q3J/TVtkdXW+L8rHxEr+Skr6jttNRjz
QaGu/E+1ERUkzgNFnKTxojM7Q1+9vizmqxE2P6mrrFKybEoVo12wQW5eMRf3XPCIIxs+/WqT3hQ4
wCuzh2v2w2SWvD0A+irYsFjilAygFB+ExNYPXCLFtVhYZnoFrRFvtCOnbtn0gm/sdhRxM09QwtGV
R+zZ5coZNIJCmQlxQd6dIPuyX0FkpJG5ixoRM017Ek66mI13Po5s640hcEHP+X4I5aAcCr4Lm2Wu
mDNBOCccafTV9DIVinKCXIAnwDazvJ/mmd+1mrY0DeBKDcYbpaoENG7UxnwfCfftZGn5WYNWpeEq
WjbEQrhnXjPubOVc5F7KAojEMKroQhLmlIm7mZh+QxHLHEuihXCPeIzui6KpGE77hipBPDkCH8t5
CLwrU42MaJVT+SzgjTRY6NR19iFHVnh6L7HRmXghRensso+I1/zvc8rT0YV/uSZU2xJliXnErX56
mkzwoDZ4GOHMsc9utfmrsxfGTosJXX+jXrjWn12kmvLLLOHVMA1AC4DHpF7PBUxE7JR2d+sXuq6Z
DeysOQ1MG9x8+tarosWgkmINvvpz4lwHjwNK5o5za2ILr8FVG66nLDOvnG+eJxUXDHviyRvCz+wE
Jf8ToX9l1xkqJkr27aPrcgJ/PQm+buaH51e1ElWWu8jnc/BFf+RlYfV3WS1CYP8svDM5vV3PHbdp
OwtDj5cUjW7XceTA+pjV2cnYWZnBVASUB9UtblgmG4AQgJEqcPf+C7CMYTkCAQOHoBJMUMmojiMv
POd2g0abT73PdxvtiinJS/Li1itr4SIYnzWEhcaJL3bnH345REA6RH7SDzsch868/Se2Jgp9mUoj
iswLaSQ55vJJLwo2beCZBAD4eLftQpLcf8Pc8DpwdPCLcAgN37uavpHGhdCX9Wt6LR8QZJFa92QZ
jDH53yiHmfzRepl0iTwUyDTTZUmutWIqlGFN/OLcXfGwP1gBTucRo14em7l3qxobGd1gtGkk9IbV
k27vOLoCk6eXPlB39G/4DObuvGdfU/FM4WulpOEi1aINmfpjjzTFHnFQmUOuH8VLOT+CWK5bs6r6
dNIkkqI3nsqyQUApRd1kPqzetubVlJrR5mndxo6E92nPekEgPhc0sXII34VnyCPHLqpUrKqhBvtI
F0lS7TdO17a6KeBAKrROOWM2AJcROophptSPUmkmcDkiqBxfW9VMOanboeE4q+heMSFBRMEodktE
R6r7fQ6JdgMRhoFeaPSewRKJUzdMq2/9Uhu/1TZHmu483HCzF6LFgw64EJw3lDgeTKoH/sV9r2xy
LVtMMg6T9EKTN1oLMwmr/tXRw94ODIZUw5cerG+A62iY0I1tAPN6PE2mggB1pckTwSCFM2WKQUkL
jf/evbZNyCSfZ7ZHyts3Or8M6YpkxpRUhbvnZ0wSq1RQhDkkwSC+0y4rVygSSpM49OTijtlvLCZ8
L1VrCClHqdEm5mrp9Fj1fBNKgrvF7RmKhJJg0R79D0e8SFIlE21zJtz2LALzZVlgfpUtFPUO65Ql
CdxAnWrBUh/KkYT0I2uBkyJcg6SGAcnjXMT/m26q2qadnfwQfN93c7Gb0fi7bGh4yXNUN+hPvPOS
RFrLJGlbDh6ofUYZw6kUPv5vlPQoUN/Bt7G1GKqaS4SYYnCp6peKoBOiKvivLl5JfXpCG9j+iu6K
MObbz4xLKNne1YVqDEpWq+uh/Yg49eS9e+0deDNGr5E6+jmsOy7SFumslc9P2FeMymrRVcApcMtj
YgwtNj1v21V1uiqfNUq605cUIwRUC7rcr2BkImXoyI0gQrODbyTjYPtLzufYWJqwP2E1oZ9FyI9D
cBraxMWaLN+1amXNFWeTcmCN70eBEhEwLrKHayRVJp6+KDNArRO1656JxyhWyY2BwP94EJ0rJzcE
mA+J78S2YD17GehCRO7m3csEKRMv+bo5z6plgeECugXg75ffgNNShl761KB2dzqP+R+6gh7LyuRS
bftTKBxLVfzotIC5MlcCu9KyTwtb9TJYDMpE/STIU4BD1TkgJrtLLE0Eiv69Zt6F3J1sHWJWZI5Y
jxY/9iCgIq/Da5u55vq3/ipZpktgGzJnyl1Au8k43q/Dc8WhLGcXoDx9fAoiUcJ3PwmZ/USpLe31
FTFmM7xNpQ2r72P9kv3pl+lTPP+KOVzvV6H1/pxZ2H4BJFL+tzhpb8pxiqyjbCCa4v2/bf9CQtM4
GGa0xZIzGQV7wAZoRhSrHQ6MsdfDccJVKE+wAOfyyGj82t4Y5l/EkjrFjf915o/Apm4Hhe0hhuV3
yw/SeZY9oB2Q8YB/AQGge/svFoopFr84MmIoDdQcLDhPC5jriLw6JODtM9fvz1YD6bF9JM4iEIWe
3amGVbrjHv7ISVNpDcpi3iqx5QxjXxbwNXl1dtiv/rARsZn+Pb5Wu1f+OSiPlAkJZhXnHHwaaLWM
HHOhxfznUA4ZwlqDEDrZ8bqD9dXVhPUK2y99YsTafKqaENF07zBdIuwWUb3S/L0ztM58URsNc1OM
YXsMxp1IILWrmevwqxK1kixjdEoUr7qP/dYJqYkFqVdxz3OYfoB/lyidPwePUbqbP3btOz6pp997
YoAESiyvn27RVkbBL7imkyqYVGjGNWZdsKoko7/3aQtFnzw/Z2NH9pgMGeT19FFwEZL72VoQfTil
CWt+/hoKYK2qe+Vtozg9Go9Zf3RCREYXu6yYKPnrboNIdIwqBAowEjoxrbpnz/waOpHsWSd8Ijbn
9n9n4/R83jQLgZVpsbJtew4ikvU9DKs9QiVhX9LjGt7EL8GglOfurfoaZQQeQvXH3vfWKaskrl+H
4pN47diI8q35NVthlxRDGHmuAcddmypaO8bBIQGVbSn2q38iU9N8fwvoUlB8NqBDYjVWI39/NMI7
p8VV8VtN4SR93xxawWwUWI1tO1kmpQsk6mRrGnF0Tv5t7thdS3IkzV1i8jnLOApcZzqecd7c1ELn
2S8yn7QBqZpS0SVbA/321R7MV974UCsyOi7qCdDn/F9RHc9j3g5iiqWO7bMzBQ/22LWYXh+QYTlG
jbeve/Ur1cVn2jv2CRt2GMvdp47cQ8JwnfvX3i4KHYzAf6v5DurM0mDMg+u99K1d7BUCufrL19ly
2svlkmokzquT9UPe+U3n22URVTtgQN2dB/j11RkGs4UgsUjLlMiJCNKTEAgcgNAMaVHjzcfRDHe5
Efr3xcChplhEoPn6pHIXu4O6jZRYdX7W1rX7V7OXRaLQzFGDak7Lcz8+nibFRGcdmHwFt9WY8gth
ATWFzXKfBpQIWjZQPMXDkRMsrVR1WsyDthejuqgOO4pnAIfh3o/x/c5ZaofJwODzCaIXkLngOph0
lTwjgxxB8ylxhM92qTNnL4fIgIE0c8x1lg4yUcRsvl8kWMoNaxwZLNC995dWYMOtrxSG8du2qUMn
GHuH8bf7d92uDY8q75aVWq5MA8pzXzaz8kNYMV35uRKFPFLZAuw4Bh2KTj2HyliIHWWj8qEsHC/m
eJNfaseZnLskAv1xa4EQjbCMVzA0LOsjBEGqovwKy21M9HG/YBCuA1aIHzXLZwDgUFf1olEfhiez
FXN1YylmqHvsz1n5bTkmoXzK+1mwgS9Y3fHL8H2EqdZ7bUlt7S/rrLFFEpmrqxsLixRVMt9AEMZF
4IEShup7y+IOBK+2XIvZV1piBMtjYeZop+RPQ84vP9U96Es4Ogl9yqfYUa/eQ/nPhd+xScZlKOK6
5uFaHReEWyrt29oyBVvqdN2Aa4JFJP41KwFsbBhT7//5mkGnCZOh3JpK7cwUmp9iPoNCudK4mfSf
kaE5FCWDMbV98UsjJyBqevy5JMwiwvDofIPes5mCKQW4XPslVPM3SH+4T1Y/bJjUlXBlvXoa/jjX
/o/bYIgJ6MNwp91FZa+aNJcsWMwtmjk31JXtWQPi5AeruZHZRBw++TlVNMhu0VIFeNVOoYDex7yO
YnkqNyR+j2PRJCy6LUNcyIP1Y1DBGWy4eEK1D73HHGzC92nzeZnkjN0sI4fuPGgYnWzT0+g9JCSx
+JfvWvPKrew4BsokxQmQvIc0wcC/gFVzQ+fVmxu8MHwGbIZRU1y9LSFJVWVbqsi08iPLXiGFMVCq
JwZEwV4jx9axeiNsQziWRNueV7eYDB1ZNTV9qH9j1csvfNghs0xy1HBTPXCgjz5sbr4nwl/tSjIf
yxtmCB/HP/Gfz43JraDeNIJJxanImeHwEnN3KoqO7ZIvazU//DlgtSBM/i2SMFhTnO9kETRCIGYT
PYK0njcXuteOSrHBw5xpctrmtdQOR1dSjpOtbPdBme6Kf5lnR8H5f608IjA3ONcsjvbOOYe8YCOY
KkcLTgCdFjQbeYmWfy15362dibdCiuTX5vJDa0fGKaw5VkxvNtAd4AUuEO16Vo8DXHA35G9bMIGS
aqir89SJS4f72q2MZHpOMUaufPw88C2tXNbPskutHLDjZLFLBAEHgFCbSvBrthq5P/2QvQjgf2M/
nYAEq0HqJOp9Cv/JRI883SWA86Ryx5d7eOrd/BrVuBfmFA46uwnT02/UdF8JOtfgZhQogxokMq8O
mOa4yy1HHM4oiYGE6TfnbMNBonY75VIKcnE57tk41wWlBAuOqwUeXKA1LDbL2mFkBcllivcmdrBq
pIebwFxXmab/6dY7lkbYpyAP4EQid11YLHpFciIksxYFvbIzLto5VBK+f+cg33X9hpeiTDCV5/6n
4m0WEPxdrbWeKcNor9AIS3tOGounE/vHYY8yHbmk0Wsk+2mCiPP8morXAHE4bNYNPDR4r4chnwiB
87KC/EEOU7+iNDzIoDotbbLnKMoAdlmFbvWgrSt4ufmipQv3HD79VvfPa6LSwLkgdhjsMSFXEPTi
qNFxvuJOQuE3oiD5KjI7nxNXlmggjoA/SpZNwlKopJ+llGm/weHPhzuY8LrZg734WiWgzmDL04W8
8mM724kOsRCIPwe0T/EWvAnZKqGMc/owkwGsaivGG0/Mt9uYK8S7ZUGMycZsRwUBVPm/9Ky/Gf3a
UlyQpLVomDXJ4vml3bB1GUuID6K+FEGpYN3514qZ2WjBqDoLdWMf6fLatGxalFxADsX88G8c2StL
mlPzywmSYmpXUqqZ1aNZq1MUSnLRkjY4B6PXpUN0MQmCJF+Z9iBVGguB42awLkMPa11dtTW9SMdy
bf9lo80q0CqF9rBDVZkST8sECWlYpMzCXR9lxUYyPw6aiGOl7uliR4mDu3fC2yxhNHtg5svhEX4I
KMCVNIfZaT8nx8E88YyfdS990h0S+CdVgdx8W2VWR0ngMkYjXRDarZyeNQDIsGurM0LiAGdOT1H5
H3kIEr61J704q6/S5CWlJyfI8ZxcEjaLIzcrLtOr0D84EQhEivuW4GmwdSjY8ewrSpusGNaUFzoE
VQQ9Cbvllua3VIV43MW2JOJufUxG52aasxBECwxwWYqQ3VT+2mt3iaZjrgy65MCQS9Z2rxFG3FCw
O6E8r2u8nbfCxMS2HSru1Ov56Hat03w9YpGWvNl/geioI8bQIc3Vw4GoBwF9+CevJMOyN8WEh8e5
F3ss/ndezZ6Ltvs3LohdGRI7PtHeqmQsmWv+zVj5ffiPv3kO8/llWXGH5dhaaxKouNPJs1QhUWl3
ZAlpA/2ch5km58d6SgJbEuOCE3uPOeokxLxja3wK6f57B1jH6xiFvj2GPMDZ/6HKoMWFgVcn5ijO
4ryPS6pDf/Xt54H33j9oE6t6WXJc+uCUaMb2/q5YQlU2CQfwCWYUTUAx26L4iHy9VrLeTSUQwk62
0kU/pylYHmgF3OdvdJcsK5NgbrWhpiHT/MzVI6sXZv08C2nyqTp5yOU0X8scu2AeEzbJ1cieXMng
/47Rq49Tq+yP1HPjHUETRaUHPpVZbgh4v/MHORFyXBDAigm5dqKdfZ0UjS8RRxKyxv+CI+Kp8VGI
NUSNPM4xBbswgLIdC0eqZOMYp5dNWv832sVP6+nhKDZArQB7WnIgJVFFjsEENugh/iv2oF0OIZVq
zIUzzsJhkc/HmsBuIdzBk9pE46k3FOX+4aN2iXQV7rHiq+SEYLsPXxvL87EvsSkZ6lc9qj93Tzx2
+WqIlZ4xKwk9AmnxulXLnUaSvRpik/GAGDmAEX8py7D+NaoglC30L1ckIAIiLWHh3vlvdcLmu8mi
Dyl2dOrk6BFmUdP+xXHUHQVBcXQF1DFHnSwSccT60RPkUAcyPO5pVXGHQc9xMeGHNo/9ngmK6uNa
y85Ya99bUM28hshtq/uf/NOZCC8QTiKEIaZBJxVDIOtmWOqdgkMpKtQQdPGrS00zQYisWpIhj7mk
LlWmoiQ6ijEuuLeppJLIDgMRJX0iAxhAXUxgUIEFvJT9pVSxTNFdoRiuFe4n47JCRLOX8aR/0B5k
5y9qsvcYaQ8YdgCKoPHVZaXPk/2rdrjXlB/lnGVIvgh+xKV37rMHsjC2BF5Jyntn7CnVyzNlMZm8
jq8B5lOakeSkgmvjmSVDcT1b8UI5u6t6SlaJ1vNQ+/T2cSUJNYWuhVuyMlg2hTJETjjqO7H8uvid
0tRku4rBSgdx0vqhzk24WBFtLDDxcLYwtMtC5HLR1T3vMcqn7ZCWKiQPVYBcPMzMfpbl+R4AjzJ1
fSqpAvntynhqfl/wQZdooMULvI2GjzlMMH9Ou5OtbRfLR8D3tDDXWHqQgiLjyjnLbavFZH39D7pF
99QcNRQWytFAidMqq7Wm7awPrstp2rlaML8lRAvCrXn4V/4SWUegXDfmljnVNgEyIasalPHh74FH
hDYx0BYab7KehTIA5saVLt5f4MIM3HkAva/Zs60k/dMPXeC3ZE8StWa8FwnNvxrK5uQ42BRB6lgg
o/G5IEHXX0xxsCm7O9+2FN9xd2Q4ShS+GusBU2xOK9ekdJ78xeZXxVWSaBm0RFPeM3YK7hjdkZT4
Wh+d+UOBQYuJqhDDUdvyqRCG9e3P8Ost79Qb2c+ZMnyVxKYlyxiZbSfAXP9azrgDYWi4AnmALuOn
3VMTHXk10ebae+ODbZqljggQag0ysVWCV6D83maQggS7V2nFKnOWxQOu1k/S4hEz3NIfyQC9KNT6
Q6aMS1V7ho8l8CHPhOGs1eoZEDN3djCcXveyMjGlxIrGQnNwGRRwczsayLxqQW3Ka49SFf1yoqf9
wdywluHhtF7ISPK8gUz+Gm3ih1f527UGc2kRNbNAui26ULC/Ct6Yxhac6u/s1tRSFknPbqHK20u+
CqYvRTt9sAFnE9jonQVj7JGNH9/nScd4EeaIJm2Ow98/8hjRNwsMbAUpldwkcstBsknOnvIkB7CH
hZZL9orvqDsb5Hl31nUJ76UrgKReEuEyilYORxU6hu1DT/QUZLNAJtfNMEOtnO0f1HT0sGrAJHI8
Gm1cWEIghi6rZt3tJgFFNHdxieRuPqEAP/H0EKhJpzNGzH1Kn/FgbVThyw9l66UWksSa7EFTgtPE
/XG3ZGFFe+UWIrOu1gd20W+d2mUTE4A2sK7FTG+nw1KULXXrev8vRU9W2++4v20Vnjt63upGWZgE
VDH/F2hAt1F+tDwyVnkHPPgFmciWXZ51hzqzpXzcAJpto9VrQYX24wo6DxXtrtph5RQTIeuOAOTk
LWZ9qXstNWmBrPx3cohWLcsnT+DXuVXjhDYTdzCV3z+5e1XY/otPaysXCeTb/M8m5SrbBIpqMBoi
aK9Oj4OhCV157mawy9fPxfcO77ULHa8RC1jvYAw7l9f/G+LGvzpU41TFCmFYs3Hvcmxpy/AFE5fc
Xs2Up3mTqcBOddBOscNADZXDGLqDl7k2jtJ30Q154mTm9/uuEmTrrG9qAhwYKzpmwagKqMelHgdA
+DdSEShvDHNMbrilSAEV1cOS/xgPw59oJtYimT34CdNPGxHG0AV4nquxn3D671+Hc7NdjLy6J1h8
UBQ9JT3cg1toixbHnpRyd9O5mQ1aKFQoYDew2NOyqN+suM8FGHRnfaJjY/biW6xrOZZ0LxnOWRA0
nzrfv3vjaC68tlDKqe0kJ4XmJeD0SlwVjUewQNclLnVtE4bHSfU4TRfp52auBI24ggMAiTBUesAp
J5H8woiPO9KQEuu3DBmC3paB72gzUxG3kzyA1fUlQ6MMOr+eYHm1Xxw0tt0EruuiX3IZOTjTOIJr
NY2R1k2Z9/77YzEisXveiajyLtVv9e1aHjV5bFaPlAd/0kDICq0D4+V/8Guw+VDVHRJTJRC8gUJV
mdh0BjZSx4UY0dkhCiXfg9tVw+L817hRuwVSwfCC3xby3yhYynLFE7SJAJ36rb6o2bc/oWuFYHVB
Aj+7Sc+j56qOaOdXKZWUwhxRY6H4X7CymV0X/5oxZ0SsbucWnQ+/nJ+4X99b+hfXooCOUFOifutH
pa5URekfWwQzamLNW/IyY54Pr6OUcE4GrXEP6K7aSgxOoy2xj5tGvcRGragRvAFJa074FZfzhirf
U6EUl/D8U2CHIIKPbEIDw3Tgee+KJFpUS37YiG4FmaiQ0ONDRNLIjAy/M0t4Z2I443kpYK6YnVio
4OhtIhn+H5XnjBLVdfEioTzmwx7hJgVNdd0hvNYh8jgXJRt+BwdLl0nOrzdm9f06t8dXBAFhrMD0
edE2IdRgmUPHb2zPZPxqcGaj+VsBcFlCAZfMhAXE+FSB6ajw8SPjClmQtd0ak45l+r2DT1wzbcv+
X4L1fFg3RaHgPR1GtgGP+R9rAGvpm8AYfvq3UwrTw5rBhxypa19j4lgTa/dTXlQnKVbCdHS+t38c
fpnnw/NK6CDrRmYSmOwgmEbv7z8RmkDYRN1ZH5YreooDwuaFDbIsSR5aTEFQy/fQKv0UOvPO8tNw
mOqWXMSC0cxMkbAHmr5mPeaS6yOQXD0+aWrjrkXg4QW0oTASkHcISkM/2krBZ5P5VSxSphReR/Mh
G6J93MZ6/oNSkjPCsDDFQBzUnYyjLpwuZa7Oj8ag9XSA1xcCV9mmT9kMmvETCEiKpLExLnbUGpXd
jyjH2zEf4yYEibpcsbcK8JBPk6xyeMevUPsef6i2wqnoKMbJbUyXzfqXgKryZFhxqsDpmrI5uZxx
PmvNi4ihY+5X/gTpeRzBkOy01M3w1wYa9v3JOXweaui+7Fu6iEHoclnyAVG544IRJfH8rdNEqM6o
zMMMmKUs/6P04EIHYDn1U62/7HyOamAW5LrjG8safsLrES8EM2DTt/RJPaEsq+AXGpL45GtUGS3v
AfC4nqigKrqipKJjJLrbI0L4Fp+r6KHZbmjfPbiSANwKUvuyLh0PeLA35GRMzdaY3sExmauiIbCT
RUsLtJONq7BNagmmL4IsipjKdjzs3oeWcBWQv9EVJ0wsDof5dHlmMLuW8ViynekbGf2qLwuf0MI8
VI0eC0H2TCzt+Ch4GWdfrlfKQkaCYAXUFALUXJ53/Ap5tzOyUZ8TCjBPHUD1BGpxdbILnDwHxW2F
JNV8C3a35Ex7ijtkOX0Euk8Bb0+l8WEv2ZPzutQEo52d0LStScS3x1eOol6qb3KUx94sPQn4Mas3
/38yKrFUq+rVR1mpEBi3Z4WOLPkJ0cnYp7sFajtN19X5HOio+zs3aW8my9wmDDQh9p6B1MgFmRfx
cYdTiKRrGPFPovO0yU2ezYNdiX0HAmiTSf8PBe5wMOoe6bulxQ4a+mBdd6ZW0T0+PFpzi+nZ644h
EGXmrd9jrkpcRG/2as9oe+qHhGf7FGRXu8f/7LVIPhb7k0msT1sGsU7pgd5z6UVIaaOhyqHxVEmQ
9cof5+JILJcWsP1JkgQcThu1i5a+GlYv/5E3rbz1k2TAPbCWpPi0gj97mYnH0Ddvti0k1oxuZrf3
JIfWUhBwrxly0YGipMJto+hG5YFZcms79f6N9LwVQWrI2Dp3nQe8kt5TPYNMHJu51y6XNMTnuPa2
WUYHwxEgKbxli3iESYZF9ZodgIhQiatKtS0AUI8Km2PQiD5at9dWYD3qdJGwAl3zh/968nlW3FbH
xsjKOcE1aASz7+wvESVoPkSuqRMlqfXK9C3ZJ+9oHCGt86I7W+ktyQD9Csmzl71Rpc+jAIviK3Mt
I5ZYUQcNPd15HjDJuANInQdgC7MVfsSe0h3hz6+Gl9KBPeCdEDoKBkE8f7+H6Oy4/nz0vqUq1ijj
c96AXJHVapr9BdpkKZr3FSB1QY4FGWT8upjuU8yUaBRgOMeVZI/MjsLabE0TG8xJJc2u5yjDIwMe
HxPOy55S2oWVkiVqfGHbmcpLAwS8sPc69O6mWtVMkrgVTkkJY9TVpC/B11BbUGBcU0cEpZUhLK0I
nByrc0RbrWoN5c27wxbRqScNSSP05BRsxC16Obox6Y3moXpIYOYkuZEKg2mdla1anU5uL15xggd5
m767N/tMZ2WWfp365J7147qhOHXGuZrUBwvINK/fTiPlOCYer6TRuKNSs7/v2O/tFBFo7L8XFczg
Eh1180Xq1Rt7ACdwRkXaP4mcl2KNXN7mfkPBtV9nogYISLkJb+600do90EGgKbsFwCwdZAMZ5fTJ
T0UvssXbjOWr+MRAjMMEJqT6FnGJMVIu3yISgJjqAMbpweUwLhpFx91kEQggnGbEhp+lddQ92cIj
mD1beQhg3pZZrCqrxI7P7uSZNC2Uaxq6EzvA+WEgsd/Iq5emYozZZQWy2eV+HsgKXqQBcmYQX1V9
l3+TtzCgn1mPcVs3VZDt42JiFeqCyuW8gv49340HtDcKUoCERvvUDqZYrVo0Kc8PP+f48gjLEQqR
EUx8+6+k2kjcVEw2CXM1xncRJxLr3mEFByISgDiBpCCRHVB8xvmICnYDemG6JLKsiQe/uPNzoJfX
enY8kDWPwzDZPTTji7vVPTHsiS6DaYNoSFNUwVREsnD6tsGMmSkNr08bFx70b/9yFEFkaicpOSop
42KpQcFUNFgcUeZWq3LaEJIVyzMMDdXXTndqH6cE5y1kpszPXo882KwG95vy0ODC98a9oy48Jx3h
PU/VJgl+F+uDSgAAO9cm3WQwhbYqH5LoAq8fjWv/gHhBQe5CnY0dHqDlhB7mPjryHJYNSeBA3V35
qJneYDlkdH1gBlZskpFCEc6mn0b9bk7QWBnTDt4N+CufE4dG9+w7fCYqdM+5hG95EzMc2ol/dQH8
gHLbC+YtJsGK4z1cVEKVFRm8BEuSYDC1oe5pu+gQPW+30Pl9dZvoI+xMy/jn6JbmLtyC8GI8+ts/
oymbEcWX/lNk8n10+Cd6gv4ZsVBl/VkfAZwTAH/cL4iGRDHHEPoGtDW1sjNrTZe8KCNjTLrqfPzR
XqQNyJScIqdsNOaEgvVhlXdJSYh1TFxJFgsuR9ktPXez9kPT99rY1QhKyyhQ4dVr6OTLQg5ipYwO
KQXcnoTxtIU7fQzVNm+09zhvNdDX7XY51Txjxy7o77JyJ2gX3DBAE637zgFfIN78kr9VKshhaPjk
ObuVkeUQs/9NzrAVzJuG1TOawc2Czn9DyZwhBKOqgb2BHhSUI3eXxPd3jZJh2Zxjkr2p2vXBTmMM
ys64PtmiZJW0l4j4xNUGtbB/mZ4TVMHDIzKMr6Y9ez5q5SxKEpUGz6eODjz++1KuvkMuQLm1DX0R
G7GDbBeQBHxcCQIg6JnbbEUUXurqLvvzWZ1CJnOSnoRT0HaXnH82bmdiHX3aLY85JPafZBpHVAy4
/l/NKNEFWF22oPC5h0cnrfPD/THBnT2PmycGWOWG+2lIrxL1g/GKsAjnkMPwAm89Usi7bkwIuKyV
558dC9eFFLZKHznga5uCgu0OgFyzdAxh62i+rrSc24cZoqdKDMeVQsdEvkxIosxuDyVk/LX9VRlp
E1JtLE2RorBiFxpmjow6sFlfiklVVrw2Hs0qwrmHo0CiU3hbUXKWJRWCWljB5pbkm06D5SwYFWWw
7e3v7MsA9CL8/N0CiawejmjPfwgDwPKTMQ9Gsu7Sob7BoyDW4qrrQm2bcaOu2yoBO+SVIpLugM0B
a5+DUg6unJCOEfZRQgEKAVH1xfk3Ulkw4zWhelS71OAe/3ep3VhOds2tdSV8ugd99nsKYcFexQO+
o13WWVZZEfeYruicExO+4GnKTQ06Y2LKnIAyo5ossZcHCdzBKTwoe4HhTjj7G3ZPibmwKh90HKuZ
FLiJvm7aT+ln1kGxRENTBtZr1s7fg84tOuOB9ndkMkPI3Ib0nId11otu6Fm3vAa8WaXihhY/5p8q
S7HYKmRCvcX9IOoh5e8S3exW/p6gIjLU92w1wWtGXSjJbe/18Gp9qslYVhs66YWeZBldhIbrh9M6
CZg8pZcHUYMwnRDBYLZrWJm7lSDkVwCd6Xmxl2uhOBGjNupbYVE/jPk+hrrKTGTpn7WJ65wiHiGU
XIBiczzKrnkepHBx5SCNLTGV+kG7Gc5pIN9y1Pm2Zvgum2n8DQ0dINO/lxUC9bVyOWD2t+oRI7Vn
VnWABwNcMYiUMcqhSc1I0fBbKvlNV1SH2fzAR5NbeUxqVJT3WJT+9u5LDh3WNtnSXDr/9d3Z6n24
165FI/Rph+4gyMc3LWZbpyC8znkurSJ6QgJsTcbrOMYBKmaJ19p/X+aWbk4Bzf3mW4nmpWl2kbSg
JYC4VO5LnbrQ/YJDlRgV3NGGDmYgb67fJcluqWROJlbmHna+l59X6mbPvLj29F8OqYghl8+PKPuR
WNs4+VcEyhOJjjlciYmRrsg26J3pWsHe0eSGDg2DoFRWhxb5I0x4zF0VAKDhSqO4vpQDNSDOtFwl
pb1EyfLkGpm2SmFcrvcragkP495BfVLsUj2rXQZvTp0crgGfZu/iygcAQxgJ9wa9u7Xzp9ddYyNi
VDDuqv1xgmbmaf84xGydswIFCpKQ0NelTBrP66YeU5AuMI50oiP4aNwfVplwmeLf2Dl0/NbkQ5g5
LXGf4d76nRQf2ve2lnkgJrQPRyLb2fzTekrsxokG16ZjWt3gNwVfL6yVdQsYSEWK1Hc4u0WdDvth
9lar/Xim85lG/UpB3DEsqCyH/gXgA/6rWQG6oqVLoDHd81UieZzhY/vn00mNFxQJpkRtTrhXv/G9
WkOb5p63nCyL9b5tbSH+Sr/npMFYvBqkwL47bRuSAb3HcX52VSSn9RUpcYKhPPmfKdYs+kMgrRPt
irafHgBMEBTJhtJt6kAIxk/3SCDuYsBiZKE7+xRA+0RXFtHKrCRE5R7HJ/nlHLqxfkHU/BLlPElp
GWc2e4O5yofBNYB0sfbg9e+Pz2RHHimUyKQqZWhRWUp8AxsjSp88uYxESK76PqSgP/a2nx6AFJDk
1gsT6+UKvZhWVVKsbqANEvhYmPJeVA6uQ1bCmfwWVVm98lIQW2RzpkwTKwPUz8GcUS098Bz2hYW2
5fsevwa1VmbtXReAW6DVuww4rSTap3NCelnfmC1xkJPNxoHXSPEN0wMnsRowSSU5Yn7P2k2FfnfS
35MLnAjmhliAdgZ8E+30GhbwW5fK1ocWxeb2wW9qBrjIz5tKNjH4whIKltTLoOMn5u9fIVYTqs6m
CW1g0l0KHU/aadqpnwXoeddlcmwGm3qw9RZZBkqMdRn+vJqByt+N1sayr6+gV6Mtg9x9oovREs4k
wcYm65oM6p8j/m9rYf0V/g7PymOAaSktHwcx81w71+Hgvphf/Z+/tR1WBJE8bIyRxUoWV6xWtqh2
ZYngZG2gdZHhjT28rjdm26bgW7aXN6PRrcCo2b2aD8j2ZJEutl1vkBnSUss/dnLa3uSqAodt6vAa
qZ6RpeQM5wSALy/dhwEB0kC7BFYyjVRV0LPVMhPRri25rN01eXGTUUQIBnaA/jl4Ta4YFR1O9k/C
Y1U4Z+FxGFsSHrmdwQ/pyPb0tYyW+/U0laHyoctBY9pA4FWe2z3SAz3zRMmS+oAEUWsNENq3rZUJ
U0h7UPUBchUSFbU99tr80fe186r4QR+vaowTVJNT18Wwxlkfadw2hpKz8xAqPYMDmdzP9WzIAO9H
EQQ6ptMtFG5Wa0qUloa+jYGocnMj0Iw33bMyLSveYvWi01CWZstkzoAV9+BJwbqijGR/lnQ+1Kuf
URL1mALPiqFKZOrpJNhkmoTnXa8QWa/OlkjQlVlZ/OEFXpblVapvTRHwPZN3JSUy3SaBZqIgK0Fc
CDxKaSJigiEIYHXgkZc3bXSDMWaKpPlwVA3LDbUGh358DEbpd4+ayg+JLRuyuBmBEPHTxUw3rD41
F57vWdzVrql0E8Z967zAkRFNrKxwn4P6FFFB7sQ/9z/eSo6FWHYJmyoSAzR56HrkL65dvYBjV9lz
IawOuOVPwkYCKMqPU6KAhGCMujt6krfh5wrKPMGhaHtj1/VXjfXkRX0vJZIp+el7FpPpx0pnKft/
d82mpHPHa3PfLzJUA6oRWBXyYfss66LGVRKLGvq8ZMN3tEvWHRtBlBgy6LkIR5HDfA3EG5yqYzmR
UH3iCQ+nO765aq78u41yspirvZRptJzebhdaD03265VNeaViDnSxwdBhSePS7tAG6rNOavgdpEhL
kUAXxLjv8krTeQfsBFiZPFX5u7DTXEwK+BbH7qhUfvwcA7m8LHUzW8paVBHA2B7VF435/bqKYImz
2RUjYLe62S9O+LmzK3XI9/VhBzQ79YUgp9bikKrlYK7MSGFUEXZ8k6B489xAIEgIpEyNEs4QDUrS
hff80wDFmsHPPJA2aca1pZfk1QvKnyf5TisqR5nyhI9/LpBC/OvKfvabmbHGECmCDndRIdhZ/Hjl
1bkavppzqy5DzNYsdgwqLCLk12z4VcM6+aKzeEjKy8tLjAs2xeud2121QaO2mxlViU34HsUzYn7p
4l8jJuGHXtUo9xNHRDXOm5dNlcLqeChZQAfgCvMSApKam0JYVEjH/36bEm0XCzV2CygX71qiFHRV
CdIfNiGsMlI+pDXRIn6bHKu9Oaf6wDe3oDKfG2CcsAJKPkzgOq02WXPg9YXxhWO4EJcG45ts04KO
aP4aa5eBSUczlTZ3BQmIYlw/6/QCo+i0vsrXzynOiko/J5UvtIn5Si7RDLT/nalrnTqllVfRzizE
WTXzA0jA7lIOb3Kr3a2rbuIaMr1liOZrkyM7cjPeHPxbCwLZWF9sB991RRL+yVJbpfqx1LcQP2+t
5ZJrMtVztl2cDfU74aftnNq7giPYjLERc8UU38qrB4uNE0HTgKH1Vyk1k0kF0k5QNxrSrv3kbQhw
UoIR9oQZh7IsUqzJJFucVDdriUMBHX1S5afl0CILK8ZhHljAGf2ExA+Hl93aXrT+qZVnq3+YYkCD
42SD3+wy/Kkospo4dLgQ7A506/zVmmJgQBXkff+TTQOccBIfIqf/JC9809GeP6UfrhtUvdkf6jex
lKym8JvfRlTooURbhnHI/o5OX2Do3oH4Qdo+f+iupeIgK+Ey5N1lB9oeeMVUgarMv8kWgFgmb3m1
oZERxPXRYByvVGNq0qxqCeGkcLkx9sGMRy3SMmflAQbGJSD/3NPEq/PpaCqbqNf81qM1Ukpq5TuW
kLme+KY6eLgkGFzGdjJilmZ3tO4qCz0nU4JLBoxSo4XLSjvh92Y2SUpWrKeJE0Wlin0HyVbFOT8P
kDmVRgbln6B+0ptMCK3EK+4N0wrpHID6XiVu6LZONxfLATcZjD5NS9AJp2G+iEFudFKqNWsxt78/
/qCvix/D9N62KZZZtl3QPRSaibo1xBInb9StVO0QOXoO0u8oXsj7kuWbAsTm4wfLucOXfCMOgzk1
jbRtr5Y8Kzj36hbq55djcKlrtNRuDFNFLwZwRv3pmYMG0GCiwnIKapQkAqArFZ78wXxyBKidPUHA
pp1MA4JX/8E6TEMjeROb3RSgR4POr/YDEiQmu094XMYGq101Y6Oih1xqOgorvZ6z+suSojtMb78b
b45navEcyNefsOlAKYdcUM0zRY/NOwjS93w5+fOU8+74bmiE5zCbgyiW/pz0JEFnKqWOyh0+NP1X
rkSlk9qCF6Y5cI+2kZ6oaKk6mTHSBEHu0dF8sTolQFgiYbhx86sbtNtKG7qFHnFqkwK31M5803R3
g6MgslqCKuw8aopILeS7PDP6HW7SFrCJw0xPEryaIZQcklXhvbBABYnudAmY3CHltEwXUyC73PBa
UfroeU+Rdk+IPS2YBl67n8rFsnIlhj76lXTa/PkkqTZD0LO1+6pmjoosM5YlhjFnh8IGepwnUs8H
JllOwiAiuCYDK/Zdp1YlbP5k4iyjU5LzwZRsVP9Ahl6Er128CMxBdfGQqtykzTY43ik7r5NIox32
f/PKHyWFoz61Pb8CcMMZJw5QveNki4t9wQ3ucdjzqAq1L0Xsgi7zZeovvOki/WtWdqoOWMRfIHfO
EzbAfWbsYLc8Lrf6LTyWoWSTJhltq7EK/Xn4UWFzvJrlCzlF7Sfskgi01qMYKii0Ilc4XDeHsKgX
UqI8YHFo/5gYkBJhZrGYFsYZyvN7C7IMwCkJsp6RBQ4+gyuQWcjOLyOpn/6xjkzPf6fq7uQlL1u0
GOIJC+HleKUE8FGUZFpAqJ7chKf9Rooefn/vlpN1q2HV2zNLx+22TO67yTt0ZexTR93PTUEUBo3v
bsX4bszXw0i1xPnatAaX71fMH/eJoFKFQG1FltgTf2Q1NmHBvupLq4Z6TDmDi+Z6tyHSekv6zjpq
FvFy39MtwnrmKFxptRl/eo8yiPmyP7FbnHpwVvzVQxxSDnRNZu72DiHWmUM0K2tf7n46psuzKZAK
kXMkWd0w7keQKcn1IgOsAmPBjtpUvgKryCMdFg0dlsTLLOeAhJkJO84gia3Rkno7neMwfkaaf1yk
OcqU2O7klZvGh9s9ehOQI5gOzcjjadMBuMaNp+EMv4fnYh6BqQ0JQyDlwgq8Qcd7JFpu/dVyPCjv
ETaifTQau8kGbvEVA9HOMh2kR17aD5TnfTdp1BUCx3Lq6yI2Aiv6HUdahDivnijJRQU7WdmdIMvh
SW/eyJPeLxiuJGDNQB4562MbnFfEosSc0BLtyZn/qlaKnXAXnRFMqzk746aXP5OHhw6j+LnBUZOG
77pW3ivkwtcVFQp8GZciCt3+X+PSbw97mEdM5jJHyTxEIC+HxRRw2GzK3+qx2ZgM3ZonBQM6QDAM
l9g6TqB9XANoXGovrJ4fXIjnl4OnvDgfCaLeKUG4UCEKeA43yg3IlGfg3PWUORVfLBG/rVBbomWx
eILf0csmrjrTzEPkRLvDY+Fcq8OGCJNU6Nc6fj8L9uPdXc/2RNKmTlmcRHEG4MdrLqS8dr5y8R07
IuINPSxk4k22yN16Enr3Xt3ijm/2YeHlQSkUUt5Uyufn+1Wx7NbMuMij9y/848GQck1OExEO0g8h
r8KN7RLnnW801PVGNJaFRNXAqSH2wO+sBCWq4RtbYvXRHSfeWQiw+q5WPebX609S6P/digbHqktW
ApwNY4cbi1RSxhLCGisEPDpQVO5r99rQGMc7GSJ9i5IpuUqSgXcMwSxzYUjZ746ZHTHDu+BCQ7El
GD3LRTOIqKW5S1XTZzCvovw60PejUG+PM7AwQpKUL+nbDPe94FI3jb52jy5nswZ4ZB0AtRf5VSaT
QKaMYg2W1fBaUw4/QH0JBAsa5Z8Xi5w1BviQKMgpSrI6+oX3XQckpEYDHso8uCNwpTLyYhr1MHeX
sE1VhA7qdFKdKbr4VhbW3WV3CFq7Gaj1Ag1phN53sgckHJPCLTefiy8S/utp3F49L/tWh4lPiU4S
scNz+1sKzGxe1gGITuInI7LMG/nrbxKyn6csk0nuqUzKDE3DbKABYoVQXAIFb4WNAu1ahtLXI50S
DFeWMkHl7z/DN2OQvwCxNIbt35qbpr1cPAqaS58+BkHBIVqiU/12u5cVE4I92HFO/KTeDeiI7iDi
3OZ810xfu7pUjHwggsSj1rCYTSbPJdRUkMCzl2hmDo6q6w8RLnr2FBQr4gOt9Q74CwNUEH8w7A/X
fflr3GnqnzxfKOguWsQtqFMkhbYBDfhig4thUztuHwu3kckABezzxhXglPMOUyO9SyzO20oxxumb
802Nqa4iyP19yVsz+rJXCCKFsYS/wWEO4j+gN5qST8GhrjnPY0G7+wDXJcJLzFY2LBNteAENpMkm
Z4fpU3YdV8Q5f6JQNBzz/k6GU1REe44XfsU0bE5xc2x131tOwuYC0QB/Mm3MJugZApvogyZO1jUQ
sFQwoNrXd2JoWrumAQJt+5c3Y4dyyYxCy+FTRHKzIeBl3NwHjjBX2uYk/BXx4i5WP6ejrr8KOb/8
QmcBoq5Xlc1AWsElBIDOg9QaVVgc2ydsFjaC5kqguX1fN3Gsf4VSpIEPqLDzjQd5iMO2050JLN0p
0k5cbWB+M7N63QConrkIoBjT1MhW583IbzTk7YJn5R/d/PMtPpHAfvRCCV0pYwsDfdf7wL7u77ys
qG5zH1ui9H57IYfQLayv1fG5jmh8d8STwsZ9J/m08Xnrq1ou/hcChCG3J0EP/tqZvJD/31KqJdY4
SWHDEhoGAnMoXGTwzoRIDyDHt3U7pdp2s9qoq3eKxumLdpsRUbnq1/uW4wYYbtEfWkQHtP/qH0Au
AfV6O81P0hj5WO8SgbXjp5yO1C3qiPcEu5S3IG5N56ucRDNBLWFn9/wYtUpqnaQrCtDHhFQG95hJ
154sMmSYTltAJyHgZo/PzqS6efDLNhubu+zoONlbcFD7/dweSS9JpjEJC0UJ4PhzHvtidcqjELL3
nGPZT9lcK2vIgOX67VRCh1w0Zx0YUBOzPg45fSKzmPzFg/CZ0W7vDFQLSjb5lcQFtB04ssxGW0EB
izvua0WgytUk+wcznzJAU38d2KxeniGkN06raamDHniV89NA539U+htcwY+38zYGjI1tZmx+4U5l
iviftqbMPosfkQ+cpC4OLKM4Z81+wQJtkInncRjYVxfp1rnvh6/CEf7ZxCt+jxpfzdfxXA6BxgSZ
6f+43NjT87w1SgkuAXR8yUomXdo74uHvCMT3PEosSt5J/njOhl68BAA5LfQ+icwNvzkgEeJVo6EC
9xszFWJzIBwpw3qzWkbbRcWyGPffZED5VZ2p70pWWKDJyij2e3ogLxyRrhJrj+JofEpdHT1S//wA
5PvByB47wckEFExV4i98FxZFGSEBuT1wSQopBJ5mhJN0TjtdRyKmyoyxzgPZ6jwJRtOPnJYqeYTy
780SVBI8fnBM32QnJWHkbgLBcJCx/ggkUuZBP68TZNJsNLAyp6janUJ1KKBB9enjXXmfDth1AV8E
axzVhgXUbBVDoi/qQ1phzmkLz+BS5ldktxwT9Fw4U7V6tfiIN+rIkYpynet3SzUad+HCfn8r/B3Z
u9nTkuQ3DPWXXvXgk9AGuEOuw7QQKUX3xdbavBEfGvEUrvYHupYmKBkX2uGyTw0MGJvLMxvyDWx9
8nWusUnWQx1BlZH37IbxZ8yh9hbUk8kh2D6C0SGy0/8YfsN8voGsITAxbTCQs9+naOlKHeT9sx79
OJxY9pinC/cDtNHTXYCUNm3xTkFhmgmY5/rsWcTPOFIwETk3dXOJRe/aWKhCVxqRWK1Lt7/oWcjs
JjJcCKpuOdNE7AJK3FE8fKGT3fMkhV3M94raxOg4q0zb4M0Jyw6inAtv1enzFrRlyMsEFwg1Hau0
hPCRkIZBu/aOAWHGElh3/xez+ZjVSgdcUmsIuaVZTnVPg3Fb/bg9slEe7c2h7YO47OQxC/lY6j0Y
DBEi3uZTJ0gmfLayDe2V31hNV523MhjSIdVaQCQ3iPK/+gnXx4wMGTkUv/NP7cDPAOfomdbwnc3p
N1HNAkGScZKSPmp+p1KjTFw3oHIX+oGwc2XRP4z/utEC+/HproM0gOirdLmhuAZB4iFcnkI/4nXX
tt4S5WvyjFGKPgyfJOaXVyzvSmUlHiGwF6a6YWMfW9iz3CrsXQIjnHGRot6Xmql8qe9ih7Gn9nfj
8D5xKVhxj3LxH00InVggAoqu5MqNHaMr5Y6L/FkIdYF7dFtQLijAbFiNL4HjU6w+S9d4QAUBdRUv
gkZfPzoqA3v85nqkuM5Rsn8qeJ9ZglnCicqflmnAKApWAKJ9PAeTg+w3gv4gmbfuylrk/xzIkkhl
BCUKV9jWeafeQa8TKDOpp02QJwa9AXbQZaiZp9AN2N9X3CrhvyeKk4g9lAymQr3+A8o5tbTH6t/q
q8WbzKo9iSU1F8c+7JJ7HbEx8BqCjgL/NyG7jrBNRqJFuiC8vu1LfgbK/tK57NLcLR/uEtIxf8vv
yhzSX5cTZHROmwkNgNN0ANmgq5nARGE0gCuF/819lc3RYt7OxOzlO6s57JeJci/0VbFvDlBt9RBP
2bfx2+umS3ZN/r8fJWyLiLaUV+o5EcyVbb/bM8VKAe51X51m4DNRr7JwplpPC0RGDbWILEfTTnAs
bEdx3nWCkTjSeas+bYVqsV76RoErU1VnoSXgVdnxfr50tqIUG2VbA+RlpBBxNMwL976Rehi9pUVH
QSoAkJy4y88hjgmBJ4PoXQMRfj+7wZ+SGWSHLXS04dacs/iZGSc1GokGHTANJwS8LP9OHyedf+Ia
IF/ruXblS2I485u1+zHBgJkWVQPVgi0mibzT7VqrAxzuLkboPnin3JECYrQeEbyWp7cNkZ39XDTe
TvN5+r8l3J9tFGaup9h3WbaSDcbrVmP+g3jLrX6jf2xsSXCspow4Kec77a0b7LIctI3MPXkr4rLW
670ltvJrFREWSfFPNYx0Hrfgob8fF53nhC1IeJj0ZAMg2bY+kmumYscvuKPfQl8aUaXVzrlUsYxg
s1Wn7Z/JN9aNXbxynorJ6DKSXNgX7Muh/Am++0FFpQPUkJdrRo2uJqvqrTdiOYH1KKNF2e36RlHm
O2Lr/NhQnyMPSaA6HSt/hVD7vrXskRvy4O3KI+CZ4Pniavt/ZAaRKiMl3YPLEOlZiFcjwJ6kEw2Q
UTIrj92exw8ZXt5XzlEJ8Me1f884nTP/dQ2CifvxKNknQaPfClaxxUIcASwHA8h9WlmSwjTZYUPm
x9hnhl03VMxw1WxycRsAWGgsLY/vbfNubRSKBkHqzma2vK2/csRBCVqzM4mCihfHNKHR+nkAF7fQ
5JXdQGYVhLZQG59mDohxxlWlaEOO2SkGlZy1fHuW2NnqMasmHpkCzHP1IOXe7sE3U9qQ+LMv08nv
8Qji2VvRE2EP9YPHv4ICYnaT3NIMggc+xxHFq3JXQnbpsoCIWseZ5WzG5kKsV7UMAiwcW8U/D36R
idWlNLh4wpW1Y8jHzBFgr8YdNB1VNPv0zWnnE3N/pqp955u+WF6yOr/ddJGivRb3GiZEL0J/a6pf
P+spgNPbpK/bJhbzV4FS6YqC49KXd/Tp+Zn2XlKrr7r460DovGdyJp0gmJDM6QIGJQ2Oq881jejC
fCg44KnEM0Cb15J3Zc4VzcnqL1J1K42w8Bd4qmLzN9eBq/v6MU2JPykUUrRwfU8JAVFfFe9pjwqH
1dHb3AGD7zm4ohbAiNYyL1mv6p6Y4+4+m5o3+jp191WnAkmYjt9bAcL5MToNW+BOqSbPh7YCV+kZ
DY65itc/GMgGXC3iVUTIEjQUGSqGInJYrmuGI1PvVDyR9PxCOniJv595P3YOs8zWzhDFKSZ2AzmI
c5MWbM9VbxUEVNWlDX2Csu/JGEOdQwdLhRUBgMkqPZzKCs/CC4I8RdcHeAxFQO63N07pdQTcSwiu
zrY9+mSVtsv3FnSDmj8/FRDbD0F5lewJdeikLxVg4xiYTZ8wrrrkaWnI8Tu/tZND/p2QZr3zC+on
rd8XlrHifq6xBCQhRv2JXCeiFlwJ9fEhNCy48GMYyks4b/rr9QMeGxzqjF+MIxdN0a/HWpTikf9Z
SMaJAct+0B+QnpgwHmb3x9DxAl6Uvkh0Ii7N0c8ckh39X3PI0ueuAVp3cdsX8/CzycHylGsCT9r4
BjXAHHXSUSvFa/o1Af3iVAUQ2GHhe4xU2uVamOshMlA+F0z8Ki+gbHw/XM/Y0QkFvJETu+CrVbWN
C8f9iyTI6AYqrq22++xc1ZDA8VbzFC01andjF4aEtOc/JkFB9WWv/4x2LVctn5qsTLS0zwwXQ7zE
3+UK1mEE2n7C8AxNaw8O3w+U+TM/Q61H9z25yo99i8u8RH/9/BBjD/WbbTcR8uBpvZBJ2lPvUC9n
DeFwHVKkddQPSayZoCTIcx7X58zDFbMIkJ47fhz7OrNucdudZi2+mEVe+ysoiGtE6wP2SqYZTD2K
WlDcoaPLtB/kDxnyvjMKkNaCTOJPAFzGW58BU1e8kRpeyuq0ngtsNl60SJuTISXTk4TAgP0A5vKB
OTAoDcFqsvfHyaHPS1Tw0cNBLMCd5gNC13CfY/CpsrGqo/v4K+ebykQ/65hMfgLUv/Borld8LImR
5sqStCEke22YsLkH84WG9gAOU4TZYY0QZBtCcTT2rXVfRqLV1eb4QupHcWMk2XlZCwFSKBEEMDtp
8axcWAO9x+XLeoM23O9Wv5AGJMuhmJRikuV9wYZLtqz0Ux/e3HPkvgy+d4aOCQNyqcdVK4GeZejg
mQpccWMiMsOsCeqEtaWDTlgo4edkG4z7cGVCV/EzYXEa918uQQG8ZJinDdjinByzXckNqTkaqrqn
CmjijzX3FlUj1i7Z8Vfyp5QySDfmkNXplV1JGiVyYjU62ZTEFcqsQ8vz2yNnm+XMtCRr9VXJbsYc
H+a0Jb3nEjaGuBVWpY3ifEH3uMw+jSKmf5dnuOD3uOeFDA07Q8puLt6KMTcxYoFqJyZXuvtddvWN
xfQmN5/GMFq8ex77vMU0bjDb69EKyPbh1/mHD039bo7F67gCtKb2k8T9/ohFyPqHJJ/Iz4K6omKo
HlRfVoKXjhy8DTolfTqj1tSMuQgjLkNJBSCQX7InCLy6IP6mxJue3adiUuy+7YSH1o2iOnlopkF5
Cfx3VdgBzPso59rqjCtGN7hn6bWbt2RyRtUtNuQk1m50otf7PjM4uSKqnCc9AEU/VVSrCt0Ki1Wj
REHGxBPbfEOKs2mvGsOBbz2EjMk+mOWnye5TspweHMNTetrDoC9fQqMIkbIyd67GU39vn2ybuSK8
Zp70n8D4YhewXhN/wcO/Jce5XDt3qTvddjXaEDijwRs5OJTq4tCLFDLs36fak95HxTDshmsdW1yd
mbY7Uc9/8a4/TFSxSW2Zxgc85b1eJm7b0JIFE0AH7UIUIvIZvpnFRT78s5CL9S7W8IXAZXnQR5Xa
OQTORhoLjDsD16jOHKarx8zIM0cgS2JkNTgeoWphgRd5VmK5TlHR5XFnLw4S00RZmDG8sR8z72fu
fIReVFXClYWKi8Ewf450b0b69bdUReUDoBV6SmcpJ+8WtonqjaniJxc1vXBUZHuEIwEaed21HZPv
x8ayE93hRCzvqVRy40zat+dDaSF7zZOPpofYcIEr8x6mRTeZINy9Bagmz3zs8WJvBT5tvZD56exm
t1lmo2ct+gIkaVcKqY3M3pPPmHP1MqScu7ppvRx0QgEitJW22IOH1wUlxmzDhVnsugYfGylYVqyw
jSzOVQ8hWDqaZXHN91QQMt3FmhqhcA5QjAvS+tUDl7T9WdPfTcTmUJ5Zy445SdJ2VKoiLUMXv+Ak
KqpD2lJUnvcJ8VD0cdJUmQWqQoIQ/xXerTIwv/8KbGH6V3CrWSaOarhPbyY0/rsmS8Av3+PvjlIj
LAJhP3VHqfXSwqvXy8iN8xhE1nCavQxo4PT51pY9il1FN/UGh568mUf25URhlr6ME9cz3Hz+hq4X
DqVvDVSBCpRq5FQEXNnXjGpxIGpcL8YSCeKKdzNAoE7Hss0I6/YF0pFfcgPmtT/cT3M/xSYz3b/K
3lSIUtQOD2LMnZNmqMp8ZGndDh7QXOomQbvAUBxbBooPEI/ho+ODYQQ5Z14lGg1rLNwbyfFVc1sH
KejtU8AUV3RdXNJyHPRRF5+9czxsCDAXxXHcj532EU8q8+VfLIbllpx5slrJu7NiyrJQEBTdRlWy
YgtagdcVQn+OQdA5fkBTUzkh+e/Ztvu5sOLaoB11wWJMgdhaWSAkzrkOBIbjNsZ0Q12HpWaw/NwK
wCi8ToAuDTx1wxHVQDATy2Dk5qjczxmHJHzx9YCYfO5EpqZ136hkQi627abTXiVz0ayWLdztKR1+
XaAnAD/fO3N2tYaUtzdvZ+3Jt4imaGoobKK0k0/5TLD9vE14HZnOp5w6aX5DfAI6p9TZ+xBzt3xv
3HprERZZueopkrPpij1sHhp9fNXTuJzOjJzWuBOIEUzERXX+FEOlFHqRU0Az+Hr6/uTKsJ+TtQcE
6vfFWnJPiWryfmsPSa5vGKfdLbP/YwPac8PQRW6TIxskDgGiBwnGR5Jq89kr24MTujgFek84unJV
yi7n2uzEoKcYO4eNlNTyLYkr1tc7Djr8Sl/4HN4xahUeusyT6BYx5dExgNP10v+VbXFeIkVLtmmY
fDHMNpYCgS6v4u9DiL3cnn40NxArjwh/apifPRI6Qyw8iscMUSPoQbxoqoqYQgQvLF+J/3XJK1Rl
xJDAAz0zGY2QltjgwFAbS/ByEwPEdAfuqmd3qh77MK+miX3cODXc+x3sDiAQFPJmO2Ga9wQGPvjh
DED9/KAsMVkDmvVZGZ4omWDdgSJ5T3NO14vJMGAlgtZejNFWN0+MnMnu2W07CNjxTjfPd/mkT4l0
PFnvN8zG8DDyJc/WSRqxtKgk7/D3Dco8M1UJGNdla4a+D0NtCA1ykLpc0Hg2Mb865rK67BpGYE25
YHxX0HhAVxspGRIlG2J4mv8ZAoP6MTMAXRLvyGNX/C88EUcizucqYWkzIHOtuxNFn0Hyfb7QK2uC
jhzRR542pwW27BISiVPNrhMEyqlgjcTgn4/81jKzMz4za9YtpFDtfdtncxV00t1UmqO1p88BGl/p
7+V2YGZnXw3GiJiQMt/CToJSrP00ZOmQHG7bLK7vkI02x+SryKZOoUg97CclV0U5cpkEVReljXwh
xLs8w2OkQtRt9xT8JrOKYM91SLO6u2a5+S6vBNBthr7B1BG6GhejmvkNSX9Tz96WthNEPL/7kLMU
HdzaPPm++Jx30RywMJh7+QVyBncqLN4wx0rSufeGhGTAM8TNYu+4iq4FsiyRMMXWpY2RizzEwhuj
yrjAbiz/GBvvL+NdhVqh4AdCrj/kE5LzNGC3APVjiCVpxJZFAZVepboZVNt+LUvoKIuRJCYT5TRd
XBNuA+8jSuhKf5mCPXXZ2Q7yQX+6+traljxK72rEWujjjqP/HpaeOteUKrVlmsul+JEfaaSASlj5
ky8KflEJWSUyoYCm3vTXwoPkza1aZacnDRTtJoBq8QHV3TTBQtmO9/mobRJUlLFO5aiJ0LSc0Xw1
l9eJAQFRUnXRI/xyr5bl9RZ1ZqP2UEgknWnmHd51yC6u+0k+/VBJsfktSFbxEQz9vXCz2+fyEyPQ
MstHQQPdVEEGWmIl+edSgg64jJpo3QIy1CBuiPBIZ1noMhp7EswwW7csUomsV3w8Xcvbgdyu1fvA
0DzvfXCfoK/q5dlDOiA8iYNZLaPG0aO7MnSKPeRW0cZQEfpNSNarxmW2TeyMA6XOXhK3rW/YjqyZ
TgwQhpn5WybGb/Gxt58zAdxZ9mGEWZ86nE5spIjCxIlAkjEyd1Hn6xt9Ab0PGiO1lJAVCQHarU4K
AVfKCMkqMOCiNNPmIbM9NjUlKxnWVfgWsGO0EjHbUyR+agZJR4yeQ1DV40Ybty4B2BlWIgmI8HSi
aCWyDJma0LMZIYsYAWWGyiZvMWOvpAFITGflZbH6qixafdw3rdUFQpeC8AdaAB0y5y1R498yALqd
Rcr/7X8pd7ECRPgQezXWWi4Dt8GPS6dA9ksoT0CpeNpexBArL+LZD92Au+x4BbPxllTzooQdHSh8
AUCBPXZzi0XKcHmhny/aBY2uaZAmc4AzHdCyNNdf1MepollSVAPtFtRCUz6RqEdrUpGhRNfaLYFn
0x4Q61KCuEMGiytsUwRG5lU2O6G04jAXuq4ugVgUuN9AIX4eOd6fP6C/XiX3sZsNFj5ovo6rid6e
MImaOl3OG3IdscVEYt8+d+MDRdPEBTZkAZqwe6Bwo15xbakZMN0g+Vx+Hr/jSeFGgLmElreAaiez
in+w4UyXeA+5IpnOnPM9KJ4C5WwHP4+9T3hFjB1Ho0UpiXSjqWywkZBo0e5J7dexWstTzoHD5OzI
KwAV7QCbxBC+2cWvWX+G7wA0+FptnMtvMARZv3rvlmWFR9SY3M4I9tNE3hFNoGAVk2BUDmeeHoWt
MB8Cefgk9Cs9VP9k2ua8qN8uDomX1XdEWAcW3i78pjAAN+D4SdvxY6MWNLTpg8Sl24fyx2p0NDe2
vBG+7D6lR8yTo0PqtcWmqfEyNWdcG56dA7WTYUp5Xird8qZ098DwJe0hfbA4nUyNxy35kGKLCiq0
VOyji5/5vsuNRwUseARG/2vzZu6h/jzmZbphSokeamw2v4UzC4+xJtgJU7zdkzO/H+URvR74ElJc
ezJ7cwNQ4hL1G+RKxHFQs/2QZRV7Ccr7eNmSUB/jwjYiu0ppkKSoh+nINnkAGr+OjhHZhxsl0Ocz
6eVYogsy18TMkvFYG0Rr5ijyiy7qenE2iTxOoxaMGumA1G+d1IeymM8kQBPDZMBo9O86CmTxiOCD
gPOUbHdp5IN2ioyhr/ldSevXdLNACzDrjvYFM77CVOocDKPlKOfm/RDezj5ARwTVTFV6eHmWwaYA
vS6KlVl8HDkY+ZxtMT6zttdFPl1Qpe4z8OESXyKSzcFBK1P1IaBQqPdMepYVB+ykQ6SkpqRzrSMb
V7jIR1SS/GfOZwPubQEntelOWQZbr15BTqPCa7Y1v9DFKPsS9NYyYkrb8a6aGYMa5FLboz55H+Iw
UvkYUxneKbp0Xqs4ertQQIdOqc8WXYBGeXXM2BNmLnqkGalkYZ+6pUAOEKfEU9I0wXDYK6NNvw8V
KrbiSx2pfXDTgkpMPy952iVp6TgNd/89TJzQoDO3vCCZkDiGItyiqEkPHAPHhhdrAwac3I89B7pZ
kT6B1WLiKy1E9w8oUFvr/2Eyn4cf4xagcZXJLjvFNDuv3QY+mDda+WSpUBcOfFUjXglWJvra1Lts
2f3VfSUt91V6tLC55Wo4/1bFyqy9LdV0Eg9fCT0VqAOZCs2U5CsdTc7DxGSgDBcOGJfOynk/Azbz
LpEiLAi4NnhIJieM50IlgKiQQzGRy+r0w9heIIL/Fyjz3A732pyHFn3X5wfJaASuSpjcxg9JLIWh
sSBsmQttpI/NFHgXpGpz8c/vc9m1YuDnGpNveWSMfET+j+Gz892drWWQUXlEz9ICLH74ufQcxsv6
Id5wkUWO6vAtoKc6QGc4gHp805rdmoDZw7LZSc9Tn4PDKHeTgwB1taoQOGrhEiEO6ZSaQepjcwRw
SQ1/+LJAY2f/IgtiaBaqh433IYL8JcwOVzBX8oiQvM28EOs9Dx1ZlSwjqelAjksESWNrQdhYLoAT
m8rnxBKg6+p/6LW3k+ac/aR+tLTgh3sYezk+lOqb9+9TeoA9ekhJceCO5hpZ09OM9Zff2U3DWq2D
T+r0tv23zXIm7OJCUa82zEqIHwhqbb9IHkG4IPya11xM8slk5wKgHbUoOlgSF8nmcanGz3yRH5/0
QY80lMtvQT/4qpgWdsS43f9QzQuVSCEHt69aNwOKMXIV9hjuDhma1VWiGcHSvs3TZvgdwviNNC+x
/aoqBuZ72E3DHa77N74BhvBA51NbQCMA+C8ZSPoZC8tDc1qSVXSsPO8W0GGTY0gnRPQMuoiHbJXC
DGtyOf22XpSXXdZyEYy5oFzWMVGzXKLqoXVkW1PM/3yQ2joZKhUfsZraT1Nql1sKqAU5K87Zn/rw
ozzE5Pq461ww3mf3LusmkcLR/xq4Qnz6K5752/CQF8PinT4B/bdty4zntQM2LEtBkvY+j9XqTXo5
zWWPsLRdaRZS7MiDHUzUGlszPqSjQotlN8Pq3B2YThmdMsHyrrQ+KpjtzCG6Ax981NegVm713kla
8XxvGENXZPD54ecVx0rA+OE3Uawvb+d58BGRbIOvEiVOjkVnHXD5EBlYgss+/s/yca3MJrNybETR
EgP9cXB9l1QgrupDh6O0FFzlQ2suBqdOrIVvxnuFuIU3/8qR4YDgehyVKl36B/0E3TQ0UJDyPcyq
adkSqpQLVKcnls7VbX0QyUbjzSvS2Ir6fPoUEoC2Csqj5IRIu8uEcI0BNd0zfKTHwSsKtfpwyP13
C3sO+/ewbk8YJhdNA4szqFV/OqrEypJDBGxwfvitKjD+hNoJIk80WrXNwyXkkm/gnQgy2/2wQqGQ
fjOG8H1yKwpuCVAJ1vBQbqEg0bgIZHkvRH791XBirys0TPbZ8o22Mvq9ZpkrqWcRQuRwJv0DlmqY
twtLz+SOZ24po0aSffHmclcxY8rwSDH0aL5pcdVcS3ibPtMwDBCJNjr1NsqxxuEGwbI71C/BKT77
wtKhP3ng2kvSaKdSd6Iv+VHiyqmDFFoeEhWqnkGpDe1TC+mTWa3uP7UH9bKWwuHfhAZ7VcshshbC
au3YxmTDkMfr4T/zxWenTZIdMEmOn15DJqo0datfvHid8Jng142opiKqEVHaCD21xEyEwes2AcqH
6H/63ewy7uYAZCDJUwVk4JFbTE5uGF7vtWRnqCngGR1NbxU2cyrMsjL5PPt8uM/GpHu+HupCzksO
SP7A3sD4AG7h/xhmx/udOAAmyixeW1GBzjwKDBNWPnP7nvZK4yLglB9/RQ2tvFSY5s34W3cM/lhQ
aI5q+07uXBtYNU3GPjegzEvq9CTtGVbhGY+LEjlejO6s7QvNRELEe8rKGqn6N4ow8XiIpWVKWhW5
t1xdFjTIMmCyBnOF/509ebHWDankJYlbLHrkSnMRBn7I02NLzrq/xl0Kk4qhkuaQwhg5qoudjHoi
HqcEBwH+dtrQlFfWwAiQnc+OZOtHxZ2dojI4w8EsUB5U7W7tN94bYuXLdTBdTlM/R9EZBvIcXpPs
9Wj25Iov+8dG+jofNeyzG0os3vHBIExVCRXnV97lQcCThPYmLrTe+SKHAMyFs/SgDT6wt8OOrYkO
fTQ/uvNouRlP/gfU0Zwr3J+7D/DEFjIo2LhO2ycSCYtHi0oJz9CQQzbBrLhSrKnircQTtV0xd2q+
1sMLhpaYbqtJ97/1BohP7FwgIz1EwFEJWmGzcftXfAVbtpsdT1J0je/UKWnwyouXHIdFZC26aMY3
FjUZRkD4cAE709Tg3YOlK6KjRXSGd6EDzCDka/7snVAYYXRb0qlYBnk20k/MO5XHXsk0slqRUXhE
ATld9TXn/NUPQoTxcljDwDvBI/7HAriZtvHxQOvXB4Tmtv+zmZ+JXPPa+Fhvyt9NPmmr3knPuSq9
zrKmAT5w4W8DxLWaZMC6XhVMsUOoDVTxJnQhLc4lKXgoNzoNhHBJ4vId/LvE1tewI33HTQOOBu1n
+K5fi2sGuu2Riudf/Anxs7DXUnst0gVnW6DgYK5F1+YzCIKv/YA2YV+lEUNnJRkMKTRLj2vT7BZg
pZkbQdiPNRDVk9L9WEpldXcLoGIGf84OqdX9zFFBuLXUr9L0LIg4JGZ7kwbB75zx55rbLkkKrN7F
2CN7WovKsmtTaHxWNLVOuHTEezD83AJGgIYees7fAg0GhBMBDSf/faBlCTja/yuNT6sBFtaBGaMV
SgLQKDNQTqA89BfhT4ogfZLqL+Mose5HL7KXrhd0emX5xMHVG39aB7ldC0d15wjTbpZ3su2UpwHG
mfHpR+TAPqlFCRZEM40P5dfLDnmcAyUiftfCGZLtZ45ce6LH/zQzN5CZXmewoXfzn2umUEL0tEGj
oAGocsrupKERotA/Gm5DGKoQWYLRUJ2e3aZCOoTYNIhafhBB2qwybxSKnAOqJKOJCvD9y6e+u0nX
wD6iWRSyfhNwKu0tp32K/kkSFAcD2NK70m6g/Bjkio8GmzbtBtqNqq80bX/C1upkU/eg3+2UdilT
DUQMG24xgY0lU2Tftsfn/iIRiS/hciWBPIrApl5qxXtGSWr8Lbx9jBwzy9yZ7356YUaQjiUkCcsF
Ze4+i+/g8xPUxyQSsslJbQ/wgXxEUlawLO1qa5mNbh1aq4zXGhu8nFv2ANGC4xc21mX14oRC+Wg/
aqtt5w+XtkMlfCw4VazKpXRnnDNjL05Qgt1R8rwCPSLHM6s1Gf7s80G3tysjvTQrVvXxpCCna6PF
6hEMPVMTYFExxaUtDDOFOt6eJcn5wLTbELGY/iA4y6FlMAoCWcluT7c3SPwxHCA/ahwb30SNmIzk
1SRrsZX1gvtKQBmGc8Vqppz/iGCIDeM+H27LPcPDJ+A6R8/fSrxoqWfCzU2PxExaNH54TIhgwhyb
SSD2ihI9t9iRxW0cpgKvfR+oBEjOvGJbD5YpiLZdQodeqEbthzMksnUYoZ7L7OXd82vcDik7MSSY
7iGeamrhe2nRfCQMfdUKjI6W8Wqm1hbjE+b0bE3NeIlEIMoFTfaVrrMe+QzThyp65RyxyXksPoX3
z21wTp7wcfQdpC6OD9kEghWMbhQYd1PY78OlKtJJe3rwCk1telvsdfI5p68r+PKNHtoxVjQGk2Id
vqDBC9vMOXvwBKp1rnNWXsmXe2mvbMSOdEBMicGBThEfNM5m5YyLJj1R2/vfBakxYLA7H31bLZI8
FjxETywh4srmTIGrRi8paBTeA930ONqLR5P6CjXzxf5S5Gim1dy60MohcNBnuSuunLQL9Q9mlwT6
CwJGFCK8hPYCHcY8v9MIKZFXGmcuuQfIOWkxY6sXzuFXinaU277GsuMVk+7QnBbVI0CRl55wObIl
qnHQDSfN9OIHHlCqQaNFXNGHHzeuT0KGbVmRWVznEO1BiNZvg51Md2ejslA5aaPR1EY7994Pxd7G
O93e1MrW5WJvW4fsB6RSz0J50j1N71cjaB5qWCGQQ3Tajk9+qOoWq3mMua/GFgdv+69vJMlcfdnj
wQE0KVzKp5xzcfsLOLYZgsx9HOsfJF7pPdGPOxOnueXwyoxUWST2ncbicmmedH4zVpmyM6l/WclA
b98yyAe0Oa7zZixL8yxgPKha/S9X5kbEoFbe/tzalVMei1FDCdBpbMAgf/WdJXBK3MZIBYdgWPrt
tVly7cTl772Mn3L8+SUvK4ayUW7PzIdS23QN8HnovlRs9rqXyb55WlHc+9OhPpT5JMwIIRtZbDrn
tfmqi74eQB6eaV9hoStzpzG6QwmpMHjhMsgjuU+tVPtAjTBmlT3sTNv0SAJ2oDFttwm5er1iEdNj
/iypHRiLI66h6kZude/gWiBokd5E+7475PlqEbHvOTi613x+4xbQfUp57gxsAv5fEDXqfrECYxvF
CDNC3HkOVDAfQSYywyrpxFroDl+2ECEXfI/1xI1u50Wr+xyPqA+TRp7A2K/JHUX8alzgO3aTJ5en
3g2kSZzm9eXCdJ7pVIWycPMjC4SM19Mg56xn4iDITs3yDSdkZ/5LSLz0furBZDUM9AEMf0GZFQE6
Xd6HQH07fK9MgIANFM1lN9zUaBtD8upgXAk+VHVtb/neEQl/HcZlS2TinjIFWfZDGnoINMpR/p5c
cx46b2LLIaPFptotop1haiWRFELybafrf9jQbtyeTXVchj0Nl6yJWLUhZUibOTORt5JZT/EpXsOQ
cvGKuE6Z03YFOIx6N/RGwAVCAJ4APTTF3SI4aw8XcQTLH60xOykLpzhlNwTSQ95E0x7dM6o2fZkG
0Z4YGl9bjDNyt8X8+xiiKEGwVTqYR4lY9R247EhLsfg/MoTexFP98cepTJCsdg1XZ4FgSGUidHNG
5UoxFLPEISR7JlqiEnJh7s+Dce3sfkZM0h40E3Fi9oR45trROr/LFGcLUtgf9FfOz44dc3Lf5FHC
aat/v8vC9AgOCE2ysJv9rhQF+7lLalLoKKiFjupXH/ck9Goo4AkRHgLc/MthFpqH5OFz2BWVLlbB
Jn502yxcDqRbDykfUboJCHQ3XNpR7HCEj3v5bK7Gj3ETQ8ZuJ2EOE6eIbT6lbgUp23rHBu2wpTEl
sMfDnAmuEio3VyZjKLkyFKGCq+72+/T7I4iroSJxr+C5FLp5O9i7mh2UAw/2PWgVP17OvtxZbJdy
/Mt4TLFaBpc7LIAVJMikabypMpqgaDve8UwTxSr3KZQig6ON3tzGURjZ7FhbqfnBj7dr9YWtDwFe
3lfy12Pl2TMYZecZRmlJpp+YNNvYBvM+w8XdHt7iSGek86nUkv7I8cqDS+ybfIEryAsCrE3HuITk
ZdAv1II5nur9UoTDOfrRy/G1nxuBPCWWZIS3XYToXCsiORG8a6W76l1OSfUk2pzCMsdmwXq62Dq3
OGcbm5Yyfmt3OraI/1V82jhkvi8In7EvycXk2xgBNoHxB3R9WXV4C+gy1jl0ptL2PIQYN2r4NG6h
fZkqbelF1pfTJoCPq6HMMan6d+ChLbW0/0BWDgZQDNvMJv+waYD2o/+WFttQ0zBh0UYzv5R3pydo
JfnBT3hEen9Ovqt7QSn/CKV2DhNYXhS4ih2FKNQYJ91mVdL0PKgn30SFxJA6glBP5+iiTuWpAOZ0
W4dgDU5K6eNdlNeottGJT4uJUZjrHwB/s+AqKxz9DtDg8MjqzZHliaBWTVYnytr3nsBkukCR3lEP
a56xxpO7af0FQj3QUEafWE3blQ9CHhI3OY2B0GFjscJ/L7XuVSMzj1OYBOqqR5NkP43IsNCntP83
SDzodvbjQp51R1vkhU3aEXGl/G7ZFvBFPSBkbBcUD1dziTcsjGrMGhDcNStL/cpqvRk3Na1AUaM6
60WH4yFRDYdLQ1oeV17ychYs93RE+UzZOPnVwn0uQJgwou7REAJlqcOK5cMkgFbyFurV6FIEjzG7
iWqZzZVShWteUge0R0VNlVq+U34vvfi9o8f3ssPXzXLBg6l90WO7btbgYiVSWwim5G7c+p0cRagY
zdw6YDGjoTNfgoOJzRgPYeKqZUwtFbz1XHuqkCNqvulIDp0HdmDgJx5spaL9Q/T2TYHYLVdzzNfA
w+gs3sQ5RSZfxcZzwLOlg5hCLpPSPAPucy2GW/Acp+FUQOt7sHunUj99fRXu9xZZ4GD32PYfopaY
qJaN96Zk3C2bsqBnpox5O/aHia97XKpY1BYcF+gPfJdEUHmimL1172WTZgaM13M707C725ZiDw4m
xiRqFJQVACZ7VUaEE4WZC9uUwgXwcKQ9/lU3Z9csw7+bxXd6bfTYZSlvnE6/aTZtBX6gPbTPV4Lr
482n+joLGX2Q4r3/l2VU/PV8Jbyc9LcicGNA/P0WtuFI/do3Rm5I9geE3wGZRH6s5Gt9YateJ3z3
6ZkSL5VGOmf7QtmD9rZYCq9hwgm5aKVoxrWLcoFhvLLWhCmpI/cBk4zGo8QiIKG3X39u5fLKfxc4
IG2ovh9T8vrfkFMFZ6pUG7bZ7dZkiQU1jnW8yKA/4cOs8M6Ta1fkwnTWQaYuRap19jfT2G/NC2Hu
wGtHqulatz3hwuGwYVTpWtt3EVLw3IqTKoCIyuhajSkz3vUr1PlmSgF6IfAVKfMsre42ompWjh1R
OrdmiBoxCsonQEkAPxnn3i/3Qw/ylRNwnDwuYL5fe25M10kyIB0ULIYtsirUl+htwwBFkUQydiWi
ya1cYY0iqPdRyh7Qqp7LryqmPRsHTsAkiyHUvCp43X1yiOXhuDyaY6UN0isE6eArLJ5Hp/ATlx2y
rBnWj/vIAIGgys3Y56tSRcG7RrJ2NPf3a8P6ijvZhL6c9Z/z0un6KqCI4L+hTlT+rEN/63r/s9yD
E99TZbcfiYSUWkH/DCiciy8sy5tzSipFDy+3M7v4AfQzVrx+2CnlseTAxIvNHGoOxQyT4uYK1pkS
Tul+InlH/NZJTCzcKAYe+C8H7lF2ZuFDago4O03nJZRcmtKH8qfuTVn1QTnAZfcOoy1bJe64Eia5
eda4+8q2n1oJgCCNPyrnwLGKtPFOxYsCFdAyyefa8Tpgfktha4PIPGKanRtsXomcHRLSPne2nNNF
sVMkBrXlO2cn2Fkid8O85fgWZ8t0FvrMM5p1dubWQZT3C7HJPw6xf3TdJnqj2CPMiBxHk5t8xbDk
uwe011Qe5RhhCIuJYJ2qXhn4SxIBcOTFdXTlmUWiJOvG8AwFkocB9ACN8x5RJ6FACF4cORAGZviQ
ttONvlErKGiCFQfj1qY6FwFNacbyn7VJqIUGIOfClJu8uGDh2JYaKSp9mPcf6BX3gy84TksrR2Ie
22bsr0jqa3Ni8ooaqp6cBx/kpM12FFrHJ+NIzIPh9Lx9oh8F72qtQdMWZiYjbsrQvQwpOmSkST0k
GisD6aP9+jUC/UruxtOCXJ+koCeI39txLFMJc6pyY6h9nCYgSZVIuSvE+rdS1h9PPHMnJI/xRaly
xlFR1s631OZ+7EAv2alWvTcCGWkRXk8G5Ii1nSgLRhf5xwFnZLmzO3wE4qLEkZROaexnjZ1XALnm
CWt64CIadJHC2PucXE3le2e7bIhw66tQ4deDKDMMl7qHaS+V81PLAZ3ZeNbomVIExl7mFeprDa2I
T/5hwsp4IlZJzn29FlFI5xKOC3mCM9Q6eQ1pG2YsUORB4pNUnQVn+U34myZL2hRNc19vJ7G7ejay
XlWAAd+kv8J+WT6vN+C9zR5I5qVgkKlOHohuwPSNWFVQyRL9Log5VrxRBKb3eUKri+t7sRkeoTp4
TYD9pLaVWD989i4t48onioqTK2zUaDKts9B9UV/npzujjSSa7Pw6fNZcA1gcmOeah9IrN+OlNkuP
1kOCH7aLzKsxt6MSRwuoiiZ2Uue3MmzeroY3WC0rR3FxAxZyxK/R0RGGNBjuRX8FWQoy+NeAZ+AX
3xuDwPh+uWImvrh1InrfBaPhIIu8f9+ijJF0WtZFOr38sJnUz2lTgJaOm9ZysJyD/lSZyx/MAeG4
R6q8l+JAxYXSVuWDsqRCBAB76NZgCY3c1ysrq3rDG53L01j/iDyykJ/HP8H5JlXWFAxZrUDzE735
bWhjAVmTFZjz+DpB8DfxfvHP0bx/1J7cwMZqmWUK6vMMCerC4oE8cgJem16pESan4UBDFyKOYdBO
Pd9Jcyu39++AO/T/c+o1rTC9qUP6T77PlPmTkJQiI6nXB7KsslpfzBbPmMqvF4K/YL/b8J36lDLs
Hp7IUChLceRWvDATOZhlr9z28r8kdiyBFgvNEYDrphb1Cr5Kxax7UsprBYgTijlM3bKUo0pWjXJj
qqcayMm28eum2Nnz+3z9LVqb8gs53dOzRco7xGIy3NtHfxkj8Iz2Hyr1l6oHMdsCCriseH+WzrlU
XSY/buHoVs6lTj9rVunk/68NJlwcOZvHo0I1/nKaCMN6IDgkVX+0k6z6rrKzBdEIT/dHFAIRLLPR
TDFFHMB51AKCP7T/DqOijTZFxpv10YYq7jFGUpIIOB1X5I03rBpm0FkgFqRtbYdT9Rfo+CcRr1ak
fp+XLSZUk4iz3VQlp2OtKprd+wPQiXefzGj4ByXV+7Ntd116/rfgvIYMPQ5VehIprxdzt0dWPrjE
e7B8edhoQHuuN+EWJjCFvLGzpQJG4rOhG6K3c5Mw7B+BCKZvrgroq9oPT9Yfwk/jgSMthrteREnB
uFTUe1Jx1Iu8GqLO1C5v5E3sDXW/HRwbAd37IF1wcWN8hp2bGH6cNFopmIrCS1jCzvrOl79xsQb8
NCP5Vn/XwzcW7rqOvZpjaKidmVWYpeUC5pKavzMMEyP65E0OJbR/ZLgE31gr/1FT7KKmE9a6uxfs
eNAvMbrnLkYLYAITOgabebb2nQ2FKqt8EiD+4uTXuo4W90ePRMWbR17k/YjDznZKYUno9M7ITlR2
cTYajQEWiiktR1zLx5cmV+Iz4d20gDN+k2evHSELAPJ9K4Ug/jjIEhsydzUZpHWMk7+x/Bd8fopd
x2QgW2bn+EyKuMayq9vYyti5jTZhPHv4GzeQjck4KZ0j8iMlE9sFMegz1K87H+TJbR7cIoTr8zmH
kNPuK8xFgzF7k5y9WhQSPcpVFCdVOkvlCY6SgiPhnZ7Kprq6cj0i2/vsUCJHBAToBFwO8F1yJ6Yx
vl1eFF+UC7abKtZE4H8jTYk/UUKiumnJR1FvZGkCXH8bzb1lS6rGTdZGADQN4dbaRG4NkEy3sE2M
7kkAq75dhxYnlxFx06QO5n4Ehd6zqeF+vT+nnHtZgjoaqGv9ShZAccU643ZEQeWJkG4qOAbYYgXF
i9T4vfT/QpPZEZR/oUPKaAxVMJTNtpFHzyMGy8MsO1Co/ffpcZVtFg4X4/ZREygcjtcYfDvh8bg1
J2WfYIyBwRIq8ta7HRIARA9Q9YCAzjI6MAeS6Pu0fLt/GwbdRdDN/ySSmKeiXq5UvvCskKTGpSeD
cazDbfYfqmupoR1fGMaXV1+N8CIXOmcXTF2hBd5L/KfWLY4pqicThLyMsT6yT/vN1lL7jjsapBh7
mruuQ310cJky11e7ZPF+ltKji1NX+GH6NY91FAIaYTH8n8tRz+luJNIWh7BLc+mDiBf67pPh8KJi
RBSPSgZOvksdgFmqUqmmeq6Wf9ZnR1gZugJFObgycgjmpDzWxy2bBZmN/AYGBACEW3BtAfMpugbj
crRbxKa8lHYONckzzkE4eTKQ8Y29CjGoHL5U99kWKTWhJ8LGM7/CkpZfxul7ZieLnKrl/mD7vRfa
wapmH42APcao2CyhzLCEDU9zF6XPA2iQR3A+oYYtYnihw4cPn0by1oWr6TBja0ANcTw268EyaPYu
KZkaetctOynCh2pvGiV8sdtvjNu5hqojII7kKFcus+a/Fu8ff0bbYKV+jl4TBpXEHHzbOfqyqnxu
xnGZ5FHesD17b1QOzjoqncM1BXaxdCva0k/sV+HtLjeGS3sz647Ov0q0wS2CpgGEBW7yyNCP2Quw
cxn6af8HzNN1npTlLIs7VNPU2bfmGfQS66yZO9J47YyfQ29LvCIfX2sxDCJT/JSomdjs9eL9pZUZ
4NBYZ4JSlWKuFRMs9FoFdMJqkL4ko1C5SvDM3RGx6ovHqcro/HEKOZykoM//235ubjXcLat37zfQ
ZR2Lp6upCw0T4TS++w7bSZsp2irKJ9h85NDnSIXOos1wLiLQNA97C/WElSx/9xvK5J/fHgnnq/zX
6GBI2Qh/GLlTp/g45/T52liVmERyBVvX53NoOQZYhB3t5lp/JgUHuiqJtSp2zIfX8hfyiHCOWKt8
f9Of2gvjH/Skw1w/qlJp4WE36vaC5V8t85hKeQBsNdceke1lMIumRIyTSewMFJewDsT9LNYm6gSX
aMnhgYweOSQ+YD/P/2YbzWBa+5UQOFyb7AttnXiblZQNVmf1kxOrVoAEJ0MTyp7kupfyT2f8COJm
VF/MjfOMmO1Med3/pylex0yIxczFYeAySK2TGzGdHl4ZZ6YtS1GbnVE6QnSMVc6sur47N1Wo4zCJ
dZbvNy2YofBNJWS8y9p7OKv6+Up9ILh8dtC10pbYHG13LZK5Q5vN9BNKvKaEY5QQuTUq4y4xj4cn
3GKJ7tKrfyQzdf77GHr136id6b335L0WovXu4gNLCS1VOTNf7WhdlFdKmwoxcblDYEKBZRiSl2sO
SPATaKU5Im5Q6X2PHvk3cwy1fZ0vFJmmetXCJhmvps7BbzlFciT8NM6xOaj8Oy4UMcFGX3npIyFX
mIzVOkYzsaUTiztqYiNk8NbCEfv1jMsDxXqv7TRazoC2+U/X5GcuNX29gXspCpG2rhD5DQ3khr6S
PKSJp7EcIh/TAJoI9UJssmhzry/V19HLSjJS16Z9voF/6bAegylM5fX21DpIoPKI2hWFDFLjZPFb
8riFBp7ImlcC09ioQ4RfXKYn6H4cvEdQzo7SZU3vR5/4JxUpNSKr1FSBX4cRnyPzM53cUs5VVkbo
49pfK2WbdwbqqlQkrXLjhLgbehS+R1jyoANvI15MUhVfn8RoNyKePQOnzeshRPYIfZmHnDjMNn6d
ZP488uLHNNYUNw5e2QcHMYORD9ZlF/F3i/NCWSvcmrjdZLH0dX/8JFBV1eKyEqhTn+UzVg1oVS9k
soCXXYCrekBBs6gOXVVKmnTxU9JjZDwP28Z5ui9eiwIPz7sflmoxpAEq0+aINqsyMtGGX6+EDV6j
yLegIMxd9255Og8azc4cqOhd3l5PfsGqLCG/NYW1gHqjhI2PeRMcoFudoQhwt0dIBFwnODRqFqIF
oURvT1C0LCVb4xnZD+mdBNz8TKXkkBPP1HCyHCuijIs7Md/awRwUtCCNefW/2rnI8YuIdYXOaCRz
IXlbrSdXIf2imkapnfFjcaPi3I2lwkz13FYQro8Q0y06FJux8xyJn2/aahIo+44nhchySWZUD+d2
vNB5aIbGOdeoRcp8w39VQv1FoXnPcsQdQ3RejInLMJAUkgDMcvhitOr09hsIDCkjEghqNUCQErd5
mEggGUzULH7kQshr86iGJBuCTO3VhD52dN5BcmElqsZSaSf4xjmu2eJE1MO2aUwmVQ8wJ22FjZOG
Mab5pttP6rScrSTLecT0+BTP0XSKjpAbi2oyNphpAbhHaBfIuDtwyolIXUyZ4q1vQvasO27VPdg2
NFHLWAn4Ppm8T/3V+JnPTNsXkWw61lfjvYFh0qIYHN5GKQ8ukSo0ZMSPOYnCo9464xuYinecn1oY
T5FUpZJNjEtZVSef96acTX/rDD5Jmv6fdLhyBaVPIO5lL2R+cpt5tTLBFrEIqROKkUSvQF8qYvqb
bkZr2DZkrPEUNUZHWFayPFfEs2NLMCJbtU2JdBNbqEdAgDKPt5vXucj550OwzY9e5V97tqXToEup
WzH5tWG23MTuS1GE9PppQOvw43jbNbAmjxhoAkvWTinBpNiVAlLGhL0Pmdnh9Zg+PJbyjyx7Q4CG
MlNyiAzQmvftld1oG4BfJPErlCtJX6n2HwzLKnY4WB2+0veBS+/I1HM4VipPz6rR2gsNo8+htxIa
tK2mcK6o4qlfq9H0DPiQjVU6Mjt4QasXNtAwhSq5RyamZjZM7XVGTh6MjA3hLOMmzilQ0q5H85F1
mr0xFEBvjy7rY1xlKpOZA1wDYAAcaGMxNZDGgIG1/IoDKm2E41dtA8dm3mFICNmTTPG80xtLV89/
FCePqdMTR154y8RUF0kQnU76+V+lJCA7ND6O1VeZSgmJzpCBHfbHmSOnoPxDenuc/vojPbMa3hXo
gfys/QPKJ3VG3twg7fkeVmWPuSY1sEm0U4OsFSzTQsuNAN3C1EtBPOLg8cxi2E/yRVdIb2RWIcPd
CBV6HgVQGE7gPyeiyvB12zAzcIvl6i6NiIw/x2TxtTJCYzTncND8JNko3IY764jwgz8FtoMBTOKT
QpoLzs1S7mcx3TH/+hJjwBxu+zdLwQ4dIy0Q3af2+KQwA7UMSrkD4qtnJprtAIYRJfQ+Mvtzocd8
BZHYRxqD7w05zi5TmJ1MaHZCPDedEWg+Oz/9uipXhwcLR8MgzeUyFNj3Nz4iH+H3S5HXFGXZ3Xyo
yrRHQMsYlhIwMu0i4EqMIzwpTOy4v3m1AkIUjmoQ3rd/gOVraw9TffI/HUS3e50cBDqAx46FHuAJ
wycxrOCBwN67/FJDH0fUCGDHASiNwF9JLAV/dFW5Nr6mKxQB4R794nJUaKiVUmQkFeREuaqSX2sp
wlJ4IEC3oehuiSAc3Wqk5nC/qTdLsnACTcHFtpxTe4TVvr+f5WbDKZL4w7EdZnadZGJp9GxcDp+s
0U972v8Z5cLokF/Et4UwUZBxXszG1aySTSgqyytia8PQ8Pa9iJGsqYZX+uM0YLbijqBwIPHTuhV1
qPv28qj8qk1GJG0qmy201qcBJHEMaCt7Iy1qRe9fNaqCuEMaDFum7SyjY/HuePiU50HFWzGItjzK
6lwY6LX9lNn9e2JG9I2Bfz1xiCUAYjEXJwILHiD9Jobhd1kMigTbimEkpyVp62oDphoPjZPCAunA
RvHt4r0NylkoFQsBMNVP8yqjmN4UwiiY9l1XgzR3Bp1LCbhUeTmjqIUk4qBer5E0M0LEd+xExeM6
bPf+IU7k+RhSaL4p1sXQjxRPGcKk4yC8WOdS/1pwykuH1Pii4gz6hzU7T5pP3l4QG3geu9rNqCxn
CMeD/CBbTXpHFl1UYvRwCZAyXl0zUxSfnu+Y2CQQK+6I0ME6thKIofuI5LZSKAvOS0miZ2imDfz3
cq7Kq9gT+GOwsCLwQl39FYGd8CnZH9obLGsD/I4Q68/kpVf3lGPZQYszCs6oVOarrdF7jKmyEYry
RNjzY3f9caQ74D+kBpAixiGwH+utkXSYWIGOP1szwhdFMLf9H9RUM6uTkT1djmfQChpledG5q+KP
O6oZB6x46h6743BEroxRPN7agZXCOG33dL92hH5/94nCAXXX47QKu+EUHMI/MtFYOBjC+pMbLasq
5mzT2eK0T2U54M9ZEim595hd+wKMDm+/tuegYu/a71PYQ+FvB3O6DMKFN+qval260g0augW46LPl
ffmOalzRol0MiIOJgYdkI1nK5Cjt5Itee/QmVFlEetH7IUVnx1Q10V7xGjcf9Hg2JXExcIP2aLk+
7ZqwvDns17ypPYMYpKfLLaP5oMLFp+IRa94TY9Gl6NsejoWgKVAtut8Ufg7pCJXyYMDKOfxVPeUc
/8uWwF8oZupR+DbcabvRi6nEfADgl9fVY+5GD+TSz2VNSsiE0wMEwEkLFyihjslfr4Q+TThzlfeg
RJjH0Rnyp8mYvXdBF1Ts9UKDc1nLQzDINabeCNA6scDfAfTiFxHXnstKRHbCtLRc1wSdqbl+aVRp
xSGGQ61tcmhh7UrgEGI9c/AHXfftXVSonTUMHK7nvCAeHMYsBCffmUgpLglgdfKTcB6k538R9xXZ
i9Vk020Yo2nZz9oIq2i99TVKhd4SzYwpKSq68nnlrZg2G2L5l2HcG/Ro3EdzPXpJze5N3xkuUrj3
SqsAfbKakSWZpQcXoK/oQXqQ6afEHXndr0fe+SETHCCsz6F9nF1/HDiqIpnIHZZ1u5tPG1ik3iPQ
juXJBlivmDrbjoRedr7L9QQRbbZUjXU1TbRpXhySS91EKwydPDeOL1M0aqiBwc61HrS6uwPMTR2A
ISEWk5+rgWi0epwcg5aeXXTfn/M8d5nPPKkM9DejiyEHUYbTlSDAb4ede3oUNPmVZ4T4BqVsPzco
fbVGYHdpPJrvogT1pPTe1MUeejZ7bnukvDWAPSKwCyOpDwnFkADf4dtGoEXi6O+dyNFlJQ72AU11
aKByg30kzeiklamCKufL+Ju7Pas0Yy1Uj0kQWevIEhLhfq3iYzlPlA/ifEUMSgHJ5yzMSpUk/9Js
5C+CQ2QAhuUqXQwAyFpq/ody3m+gUZuw1zAWpeLUzgazeae2JFa3S52z8pLayQygMYGjrenZ1QS2
XzVDO0ufoIsJ/1fzchFDpqQHoyZPwZZ8wMIE5+v5+oqqDdqmOQ+dYavUP3jqHIfDonYwniy5Bp0z
/Xf6AnTZH/hseqV/TGiR3SUG+1yCVgxU0dmJh5Xu5VA6dyL2lFd9ebduUSWVicSQkMs4NJF220uR
gKm70eHsTm8cEj3KfFSiztlcxSkZlNLY+uPpQz2LbYcm+pZ/cqt6a8QWKtI8td36MdMmJBkN3Yoz
ziOZQiCqprquMCkdZgPNEo+aG7i1J1n31vYp4OyL81tY9IDvTl7uYRCdxAXCANHkwTCGra97PYmp
E+r9lnNuqNgGHMIELKjqg2Uv4b1X2bWsVzn/5Fd85wiqBCosdzOXK6vjpto6LC0Jz9wgcETHgCNW
h0V+v9/IH4DSdu2EobDuSNgcFyRQrHNgyVE5PP0EoKaVk7ctUACT8cEWidlayJyBL+iAiGmXx5xS
2fCgX01BMzs0zwSmXjDpNLcJYjllGg6YtGISooug0zyxe6etJeSWQt7X9LgEdQCinqnfgkdXIMdS
IkrKHbNTmqiG9QImv56SW0hPhImb65ji0NE1Ux6/c90Qal/YsIyPQ7nkQco/6MzMebgX3yc4a+dE
odhMRW/J51GiPGMvX2N0W2Js0zIpqwFJ8eFRAfYNVPbHiF00e0rBytx/89MrA8G3dTyeNi7oTWj0
mcumyWrSiAu+c/SycJRFHNx7wQo7dJG/eSNqt3OFMNRpjgiJ9L92kAfvEv3TQLJwkNbfps2DIbxu
baa+6bWxWhmLoGl/FFNOkQ37bU7HwK8UrWbdef2lACjdasculQSaclQOjvWIr3mwm4nMwzBJZIrK
cZBhVZaUnbWWigADkE3pcIxwLrrEqUGPgV5IiKeN5u9RwW8EGQYJvVJ9GS3CKI+NZdwaPJf3txqP
KeghEuxuCYvypzBaj8xXPQc4LUIGBYlO5WSHg0vqCKmc8Uh21kzOebyz50raRSiZ63xq4r04PMPj
HAGmrFfHyR3eDbcmXiipH+NFGjWq1zAO0cMk5qKf8ckIAU9tznGDJrathRLvTHQbMKHQBWVUWlQi
j/f3aLx4kq/5sTk/GLeM1dvqsLtJBWA//o5uwSSmkCxkmqDNnVokU/zTuAx9XRMz0xJ66G8PSYid
X6RiFEVAOP3vj4bZlxW2G3ssYKP0j7z+8z2ILehXCafjGVggWnQawQqi+BoaWVd7BCEGFdqAzJgw
NYNnohjYoqZrWOhKQtaYU/4YWWgisbKQ/WJZ5sXYEiAhSAgaT4dPcWxT9+ljZXP9ox0f+mrKTA38
vzTxnS2ixSSMrDB3LlPb+SitY+9EnPxMjAzTJB8pLbQc72ieEdeQSLuqmxaG+mWHbhuRwEADcbEa
IdRQhCH32KZKmqpiroyB6uRicx7hkN/SXjrJLXFqLwSmXAp4CupFTBNybqv7fUcRmb4S5W0D2hrg
ylOnfFQ3VqF1lyqSjsoVgQtBDHJCCCje1QgGbuP2TG3dtOkhkrV6xuT53fWtBf5eYcCyLujYVrZk
w2Ms9algVR/8hjoGCrp/c8lG02ZGue0wRJ4t50XCdn9/GWQ7+U9DVHHDrtsJrAUn5WXWV4qhHW2d
mco/RoSCeve+cxWZsaN2/W/810eMB/D30lttDs9SeO/7zY7Au5RjCiR5OntXX4QNumPdnq5SECZ2
VY+K7RDzZGukW2tJV3a9Y1JA7rLP2Mahb5X0F5lTufvgz+W8zlBjucecrDnXcn0e2dXmudFDuf9f
1gdzwsuNmZRyyb4KwjAljRiYrGcMfJowBs5s/e00+pO2jWeNHiG6D6i199JVdmw9/85vKNA0SDYG
W71VErHdqE+fXxkjFOkWwqpKmBrP+GPwhWr5Dh4Bx542jjfj8/L+kQTAid8oAzNmWeRB7RTYyByo
jO2mbupAjPtFsfYu96WJV/Y7HZXcziJzuGqLThV5UgF8JurW0DsrzP5P3ADZCioohkZxqQ9450em
CwtQtMD/NLi6cMy7u8EJSf9Td/Fpolx/mQ9Uu9Qi7WsT+qQozb2yaBUia3+MecNKL46kdyZyiuK3
lPoSxOzGgzAL/HhfBzRAI5YOGDOk+J+evD3kFDm16DCC2NYHwemfFjerJTgFCJQgFRqPOo6SPRN5
ZMfbWFj4bh52UDQHMP84pZhTzRor87izgyBQpTgSiS1+b3PvEj/XLccHJ8d42oZvvWCBH0t3S5Z3
kpDBGA0LvO81B2/zklQFcccohkDvInHwmYrd01BXDjjHsdLO62zYDV1NJsx9xV45NLfC6p68JLWn
3ifcTQPZcTTtMmELGoXlCcQS5uGL0ajO9bQTld/Ebu6NW7ixfQY441SDLYS0AlhFOIUueLAg2kxc
NWR8q9HOQHG0t7Vg4d77pas/JKnfeA0XFlBKxwJmYfN9m0B45Jy6VCc/her+hxCBXVlVQ647e1U+
0kAX/P+3PbnglxIOR+FExhhbRuFfmyJkjM7QwlROQuDGs3tabKUHC22zK7bZhZqSm4nLBkbkLw0r
O/yOI1b3DVPkb4Ut42QAhSn2+ZgZX/JU/DDBzMp6r1rsV5bvTqMLjdjoRUxI3xL0fv3aUer5nJvz
l0x3DSFKAMZ7nXRU4qukO8+nGbkU6i0la/OSguJW/Zk20/XP67zc3bKnb7eJl+V5+tVeWcLrZi+o
7+SOUKICklq2wqRHJs/UGVdkEgHyYbQRExyWxLXEMl0l+z6ejlA1QwgH5elai8xEQapfPmeHvwNp
+iZYTmBk4fed15YYSJ84yfm29NsOggZgTIXiZANzIi3lirdMvz9dAt050uzeR1495KXogpYWrkeX
N76m4pftTla13QGarjtq9JnMC+dZ+IV+OJzjU2uACtvmZLxd5s+qGrPQQB5hLV+kiwIMmfpsChWd
tX5oAaBtXGnmTiN9Ennx6ltXsi9We3IiOd0yR2a6jD9zr1ZunAsAkC1soYdqKRPvIZEyNAc0pyGr
z86j2wdj4If9rORydRfdUmICUqR/8zR8bEmaEgaCHJHg/t0SgXNVHhI+uhy7yVrzQloUfwfvBZnq
Ax545GGR6TWQ02WGO/v1dOQ4A8kCQukwm/TnpdbEtyBGUBvGrksj3bDYMQV2nSv7o4xMoo9qZrqS
nwLTcjffrN5MqtG3ux0W+ouDLeub/AyO/8vZRSGdK2Z/R3nML2WLojukFpM4n8LSUabrQEc5YT9i
GsMGmwZPbpMc56rqOPTsfS86RFHMl8NdgN8jlCHynuakGyWyGjTaF/k/u0xH66X5p+O1Di/Eimiv
kF+5jBnOVWuqmond8YxgNSVuhHcaYjfcyCtD6Q7DUrsiizHteHXqWgVxookVi27a1ghPVzwUyeKh
mQrf2Ij8ziGr1kUEY03AiagOMfoLeFiTTvDmdIYiSRp0qir+KjaKdycIPTpyEqXgZeTtF+/wY+mA
n3i2AgJNq4SIT9oAkzSOYEK2Lj+jRhjfr/tGSFPFzk1oOuG76RIyENMEcMxoX/yn3FAer05dhAUV
BLUCgvVvG4sZryEv64OjQsSiU+OzDKrhHBqM0UP/Rshmd1ltkTe3+zGxNzgMb+TkdEELaZukkG20
IbJ1zcAxoyy/3HlOhXrdO+VY5Gm12gDZnm/+CF0HmjmpZkKwaT72smEe4Nt66vR2KaebtMH0qx8x
oVgGsOfGBBg5J59n81IJsWu6KU/rfJ4sWeEgZK/j90RD6AFXEs6wC06DZR1Vvtm1FaJsTCHv+kGg
HZJagfslxRAyThLaGLr3Vk3oIpRJ4PS0H4crzuMhehaK+Or/YV39UnpmxeMt+hmyDCjAaFIq/W4E
9an3FgqxG50wLckaNnMPfHmnVRp9hJpcEYxt9ys1VtCmd2vgOIJ9QNabOOr2FcTiwvH+9GyDBfcX
AZia2r+yL6NnS3/8t2P1dPoTnbU87nztmgTXJyO5A2aL63t+2xI3zvOQlNzWAQvFlOcxmmXlol+Z
AdqomCb6yKwvV7jkLV5jwedR2EXhCQqJ2AoJluks46sUBZNou7ya91oAIYytyZU1259tDl9nMoK4
QhMTIcM8/Y8xn52PkUclPHmokTUCnpw9x45SFcQf2tbXt4CRTMulk4xFPJbj0Ws6b3rvMg9yJQBq
IoDy3hAsL7BPzj4L9eUkTDcqCkOA8U5KdXUq/xe4NOJ5KN8VfBSmZB+TvpCmSiZOHa1SP/BzSoRa
DNCUrwKSYkg/CYu8Wpk9CpDLmSzodNnEgVEhLinbKeEjU+cEqpaWWujUu+0TBUj7M/MOkYf7Dexr
Y7KKINaLZtpyhaq6EobkAiysHHy4b+eXL1tOJPjSTpkW5yZS5bxK6J8oeurCPbmDoKK2CsqiTH2d
hfTLT8IxqxWDQD35iLAi6tbDDyH5I3PRRty2RTQuvOU8E2AgF87Bz4rhd23+L4O9D2Q7k5w8VMRG
UDwGIg4WhDLxnMhQZiwZvTucOXa3szEeTopbkOgMjG1YR5P1I5zhHaItWide5AVf5mJH0MfOWQU7
DPtXuzvafq1HRoMf9tKR05DmnUtqAA0L22YTlcB7QOSB7AjrL+7hl0ejdh/GNDLndKZqzQ//JtaS
sAdOzjLBrA15VG48FkaPe0GpYm0IYxt2VCtLuT0wdILBKI2R6jEOl1DrXdCYRNFK2ckMoXHqPTmG
mB/Ta19FKrg6iDinDEXY+12IW38uLZuOH1QIErj/0b5prRE5IGvicYvOcuYz8j0BBpd1bVDsZyh1
0tBDv1+3I+2vu5qjNb18a8KYu8mKVLOvKmTy9sLUXFGaDWxGEsYcOSjjJAiympHHuYqWme+GSowu
8vRFnLHmO4fkbyg3SUkBXaeIMM1Znon68heord6pzgevuP2l40DMr54rSkWOm1xMX9l2lGn+T4XY
bl4EVf9Rqv9k1E6bd80BwNhuGixg/L06lKC1mG34B6HC1iBbM917TfNL0QocH1PCQ0OIrPoeXrPI
eAFmdL/kamnAJ1HaT935OhjnKCWHgSxsCBbrEvP0or5QtuHXpYnwZwXmANLtrZA+0RWtHM0q8gZb
VxVMn2lD1bTcaVi/bKGYBK2rri2Y/HjclH8cW5nm2hpi7E+0hQnDufiQhxMjrpzHxBCYUW3/i1vh
KMyn7bjdrJ9uROzKfBSRlR5dLUshZFRI9mPREP02OD3GsSoDVPeS7XcfyoSIUBkK93lFPIUwxU12
Id6mzSrOmFKyowYhl/vyrYCKVkPQGwrhOfNB9c7zWqX45e0IrOMUp2WpFE0IeW5KoO1AJOCv0qEN
uJ4QCRrD3KcLj0Inki/IxvzkR0yLrf1SPVkpuTdS6gjArT5dY8hrN0e1UppLYQMkePEdau482EcJ
F7Q2h+7fUA9p+i40je/rNgJul1ywqJR8IdI5DnHGNkyBBtkOAPptdgxE+RKWwV7g+YYhP1Lw9mo2
+XpTOFPMDM/L+S+FeODdLQ9h512oZm98yR/Y2nW7/q+APyW2+Oio1ahDNjIVZxNbQ7ls21Oi/0YZ
niq2z+ps211QJjAdZKhlNEW3dAOgCsbbskJc4apMcjbuQVBifB1mg59XBoQOBmoRi4KMmen5KebJ
BdpnqsRacHgwEHnAiZmsSRum6JcXN48olng/mIbuosZlpfY3ZLPtINxM/W9cEhtNsFsA/1VzMAH0
F9AxJIdBnGgo9SNVc+JTF8qUE0ugHpnCnUW+M9MUttTu0z4GYx+IaHc3d8Tf4CHnFCf0vnXVLRc0
ZBoKg9vgmXcK1aX0qNC2Rhai5S6pJMfKNgqDgGVI1yVFGuH/d4xBP8D5enWjpprFtNziThgkXQS/
ZsTLHAOmy4Jjv0zyepxiaQXWhfkKafdQ6hAXXJn4CO4WZ6kBkKGP97fly/p5lVidoHaZfNUymsz9
x09CZf8urGgReZlXquBe/aW8vaa1vWMjM9wEavUDSYEaNbEq6Szt3VUlq08Tu8Wb8uzBg+e2392+
XFD3NaZjpN3SY2oJrWUs9cpSj3Soyt1wbcofIeuFRvuU3jn3jxRrtlMk4u+5PsKPLF2t6JjY/Pvf
qXq1YH7wKDYCfSns1eh3koNHe0RceXOHm5HJeJmawF5hPFSseRIsvCfYd2vCTlVp72jYsc6oJSEF
FQ1EE+txVnDZpW6cbP7lUFSv1NhVFrVKwvjSgFm6Pamm5RAEeVTV1ITzIeULkGlA02CIvCRuyVTJ
dE9T6CEC1JqopH6NQrKFhiGoZaZfMavcu89Op3zlDExVZi2iN0fCdaMuU0W75lrkqYAVhsxV0DgN
L/uaR63Q382JEe/p2Spup+ZeHSqB+82aaGD5NBbfimts7DLlPrHMk0tC20fUgDeBLVW1mjJvSFb2
St/7Jn7W4a7sLt1xBJIDeD+/LE8o2RemoFdZ0tsAsuC0CVzQwu2+pgrrSCh7DhFRDCvXAZ/sIOM4
hgaVz+pAeKZonaKoBfw33hTn8lLmkcepigmECfOe0gWoY+sMy8UW4AZhNdwtzkdBgOpBJ2j5w+gr
9vGk3b/UhMakrVBOqhC8XeSrM1b8obFALWnT9q5RONmOp5hzYre6iB+MXzbH/Ff3mgaSUlPhAczj
pDU/JPctitOuR8BcKONvaPfQDBm7/reDYHdgdLNen4sGg4NMw9cOx5UPEPqc8V6PTrVpbB2G45Kn
vnBXzo45QBXn7EUbL9uOHTjyhen1eb76H4Gu5ADKv5P18fl8XCJtPTpOdTdzY2xR4pn+xUZd1eq5
8Zd4dHO9V9wQphr/AKkGqDqLqcSLufYrQyRq99eW1T8UJ64jpml5BfR4EmwqfJeM/PCiVGVKz26Q
3MS3JVMk0MfWJHMMhsR3P0LPYgJJ4H7sHzeGfxs28TNnqQa9C3Bc6AP4GwSLSgElsrzlqvu2cLRC
Wxi5Q92+Gg9Mf5DH9yWdZb2YL92NKPHco6UO3dUpXbTuj3gStqRLyXpjhyiIsXWGBgaKXraf9q5S
p8Z+VU26Wy58fc9hSasP7AWHmsx/opQWbd1Lu3KhGFiw1dU0MFQdp6A4T2qkWangQJ5y8402G7II
dsAnjLXUv5E4jKqfvAtVpX8qjzJbEzDXF5xwPypgBMitwy+MdOtV6leI1txQpPnYef3jwe1rFFsp
C5TrsBsCDzxXrjdVi5I7Co/XXXVubzgqlIFfOxe0m1s96lmH8foJCwlQCcfYuBAKfIEUTmGt2R79
iGz38wG3sElyLdISa88SoUHB32xb6ALwauPZxY+wWBXbGWLVh31zkOtp2tUMsYY8Jcp6evvPiyiy
w8gMhV+mGsGU43w134tr/ldUErZoHYOhk/tDkT4Qv9XKAKbnUM85YlI95KIlt5OQthfeugytvmJr
n49e2k6YhNcQew52khQjEZkN03dyaO6zPOCnx1y+S85RxCmun+apnAZB9lDECokB90UVrc2+g2W5
yCujPYbuYzG7EZ3y6USVr7CJMFr+TRQazhb9U7PS1u2D/dWmfIvZbE9j6LsFZX9MJjh8yunlJhA6
2COCjDRbeLzaMqOagU8q5HG6WlAs0X0nVrOw3/jWTGN/TbHqzN99+H5DN+b1dy7pUEjQOnJN3zaD
KdicRMRysxWqUfMpBdM+ySX9uZGtklXQPB9nUFtp3JdE074giTXeG/W1Rt1gPi4z60GxKHjJZHsf
zfGWSAk35aWn4tmL9D4D0bwIox+CZ7gN4RDZb1w8TTQuKmz5Yf+kcCUdb1o/iphU6HtMjuYPhBe/
l0r1sU4PI1LA4jcttjqjav5krpSFrqjhp0qIQx86c7HWCeM9dAmXDyrvfRQ2N3dNZ6rWzMT1RVZ4
MVhME5IyRG8Ddxavlso8CdtfdKQEhob2nR06JdTs3AUxAiFafeg5geVzpN+Gl1rsZpJK4W6PtpLD
m9EkVW3jhzWu2X9RhuSZ6oVvi0ythEFPRMk6sqlZMyg2SS/I3Zj1pkqQhpwi/fhgPUywwMSdwzL+
ttow28702jo7/gC6mpN730mWgcoZ8h49AYmlCI3qmqRO7Sz8kRIpyXjrigIdUr8GWD79FVhRPB7e
eKhM/r31hgrbg+csTh+WijjlYXCDIwwWUmdLYE0GAKoNh6T9TK9QxD9AXoOfECZyrSqs4RQHs6DX
P0eiGWfwqHvOdxJoa/mgkBGFMFJXKQyDqVQrD+ychlTV1wRwUxMSUK1OxtsS+YIaozNFXIe1hGfd
tTs2D2Q8rkuhh51p81mjmf+1MmyZT7zlNXKVVxgfImonZR2Eg7Whx28sedJxHJjo/hUV6Z4V4nGd
9xA+HwsFE2L9qPMIiV2C6VEyJcsG9DhtpRbjXlzfwh3XYXzwEk05fNUbUQ1XGCJe/YDq23m17K5U
S0KXbQZExjYsTlVIbIZ23sRvp1u/ovrtrAidyt3yJ4luj+EIR7lwu9cT2hMpyRtClR8UNkd7d8sk
BFhwBCZ6chA0oVThUM+eb17rjD9ivKLzzA8Y7+4uPS7Nu7NUfXDTykv5I4Sq4+hfAefXALFWarbU
G+/p4ICF7vDwxpentDLsSq1T5vzhFS4mYymUG/lJGQZbu2GwHACbIDMneIcVmE04+SQTqpxkADY5
QsjWLZd2U+V9DKnfMamngDsQIzClJpyStFSKROBJQEXORQB7nDtcXYHEBYTU42lRe54SrczyQ3Pp
nGSNSGy6KWTcwiAiFlJgZBsYXBs4vchRADBTUPYI4JtuCKm6JUWM5484itLYMXxD81AptCFzWFp1
ZbgS8M0YixxWBd83BsF2kPfDn3tmhhx4+OblFkDXSlKwjnohdI8aYKHN/AZQq9bbzx+jNsE7vTRL
boQka55tavWPfa0Gq+q0jAsyxHJzHFkymEwwLbFp6HlW9u8OFq8sJYoZLIKV/C6N8pnRA45HLCXR
r0mU7eLERO5E49vRWl87n/9f4QUMUF6mUQ1qhNM5HzTpbvukA+G8oI7IHkV5nfp0l2RHlU74D1RG
HXv4b7HaMcNcbYE5jfaos12MmTH671jYTxeUj9n8i+JAzeCsHi0zsHkabI5uuSYqS53+HPsPfBxB
+BERMg/8bHwSuk0o/rAmjL9QOTdNUAsW8UNulgiwX+YEafGARGb0tDzurFp/jS1wyTL91pKPYTj8
98u1x4GCaBHsYjnEEICWhHlppcwKZx7mFfq7M0bHrviIgCrQqoqUDQKnivcCc1A1EcBh8ZUEkbgr
krGP8SmikDICigCMRK/FKb+MEsdtRwgrnH/Y/X6jCCigPt+s+0aNA4XlSllDi22de/BXtfdXS3yg
ldBxvvNdK0w9FDZhCK4BC20Ss/5RRIeLPZ3am1fVO8JbsrKDxUMUAyBHx54GTC/zIqt7Sl6xz6HD
9ZFkcKGgtAsTEl5oF8Sw7g3PiEIoqLGvy08jFpLpTSesdmijIQs0rNh34fV8wjb0NitiJZt6FFN4
+rAgouIUzcuvi4/4sEsl0Vtb2tSZ851nVjE17vhOBBFlYwxV4+iIXR/cXUvpeATZrA+DNenZ/mUw
fNnwOncFll/glwNSG5BMRTM0vpFd9fTP5uQoogKEl4m6tnmkzMECWuipL2p1jPbYbQ2Nm1zSDS60
eUYmNuCOOX+YFH4Yapl+07haxPPeXX3EPdMOw/PEhhaPyQm9OJTGEyngUrgHNpoBoWQibRn51PTK
5ydWaOFJF5tnh9GHCbruqggriQ0JsHhtv4KNKmcbW1qNu/HfO9imHVMMayEgCERSHXiEJnnBV7Im
eHTMnGOPGJPI5L2YPIrYfj7e1Utg2nfEgR6YjkzP256Ncat5QW/mAKWAZiqCey/4eAE3exf3ahDF
0An3DxxlloyMSw1uLhAzusemXKObAjVNCmy7dBIIIFKk3UveMeEUhtmU1LdwIo3JBccvzKbN0isy
rtIxKB2LfqQHhWtiOff7E6+YO2U9qPFGt8sSInZpZbtaomy6R1BJ/bx3Cqurcrc1RIgae6/ZdDUm
GDDfKmhDYeqmnUo6Nekto2FvRsdVm4gi5xSGWPDrdc+zbe6+M47BryxBSKrrpRDERrsab0XIoQr1
NMkKNiX9qa50JI5p8qcThwt/V75ctmHgcLOQhgsno74pwoZ9oLccHKOjO18mQK3Roawc0wPGtly+
xfAYF3YU+ZWaSuT8XVer+ndj0CIT6x4fsknQW1zDvrIl+nTXUvQU3iuOc0CGpyiZlVMmiq8hu5vi
2VvWPVaUF/HK/salEZCqhsysFG44Tc2TfEOPrI/3XETmgZ3Vu7DdKch75ncFWhgbxnF4C8iQiRyz
TbnPt5T+E7yAK7eDqOSAtcZHkcE9vHkoHCBSJ46KzukpEfxcxlkmbOrvd4Ar2+oFCUasUI1YFhng
yRd2wUXqg14OYjX56QFdjKWzBZzPDOlRagln1xRSm6XW1QmzFOWHsmeLBhV2U1U62rjbJbbjJo9a
BXCuOdpfD92z1/wL6yhbn/R+UEgnnU8XMNHNySMUNHd9PaiC2MvevIiWz+lJ6SoXYkzmmC5C+lxI
rz0FQVTMPiYKXIXHSqPi3rBGLNvFO3R42GDEIivf9OlZSbxCErRzAplKGyTdj974KW5eXPyGlhXY
TcjTgkuDmSJ3MrZ1XLWdGanffpelvNYus+cHttHzvzkpIGFVN1Ev1NG21DB1++oqsccvszYrRK6F
bH9r0aE+6vRKJYDOFwruXKA8zBN/0LCAignSMNPS7uT45LiC9Hnb0juFjbcZ/1tNh/uIBQcIGRSd
8rbSKSfe8G0qYOTUKWftMZw0DWCglc6y8nJ1rKb8N9hRQRYjdPoUdSQZVzmjINq19psNNdEWc2ud
vKD0+yIVtRJB6G3ORVNZGGAYJrMKTlwr1gNLWQfIXyW6ro6bPbP2tZgiZvp5QH+q0CZ5chKs0/xh
Cp49dLUI5LcSMaqbQ1lFVsBC8MepQRniYGAPtAyqqzxEhJVw0tr9n58DMH9pLOD+4UndBxO3/qaC
2b8lpfmPRdWXWm/5lLpWe2+kh9VdGiSF70/3kg/iWmHL1Pt0tq88Djav80zEj+RDwwd87+Q0WlD7
KALvILBAfsBbHfzxqqEF69gqW8KzR3zCOnc9G1O/Mie/ATJVFnFfedrINqHWVDGsvciZ41ANCjr2
2P7Ik15H+zCVtBB1B01MuTOJY+ckDABc+PS1984Wz8hHbWBb/c8SeNFEci9bqCq01PFnaS4tIcsR
6lpqmtagXHtAB7FuI/ateH7u8m2smVOjeA7v67K6Xa52bkMOaFRfo3ls2QnsYK0Lgux/JCP4dq8h
5PK1websh/BYNLNesrTEmLb2Kjdp5brtrp+UrbnpOJ+uY4ZRTYpR/qcvl+wIQpVvknYAXLXxLMhc
XYo/xDtVmra/2E1l37qA4X7YWIRSZQqj+17VfRbu8+EO+AZfthtcbxO7LSpMpVZbwXPfX8cLi79F
JQjyTji/phqd2UIeN+92XvL4s0e3+lZ5Vl/ZDidqUWmkCJMS7/dYcrjDIVmJaZ962+1Gpa8jPHZU
0f0PCHS4p3v6Ad0EpPveXAjfTjZL3g6QHvAUIm5JREmiXBPkDn/PGBSWSvbeNV1S6oJeHoB+6X88
fWOlWziRf94wCGe+7ENy2x8gm/wNucksU34o/zxN4vcBDK5oayo8MuvyK2LzW71qZS1FkC5Qv2aI
XLQVGSAYt+di0vQ593RNB2LgxwPQVhatbNucFYhzadvE5L0Nf6yY+Vw7nnke3mEpJjgWWPN3/eke
2kR0qMuIVQRAoyBBOhhNxeMgRtMCefDxYD0Ah6cGbl3EkMBAEdRaTAryPyqX18z7MlrebrNM/pow
kHHE4xoyQ9ikIWLU45gkiHv4u3FHHYZsUbBG/NgHhNpd3l55nKUaswF56HW1vTOAVuSlc6eT/CsN
Y73Z6GpL4Th6tnOFBqqax3xZ5PEhpzuCP+jzTCaiDe1e4I0cOXJbC3aM7NhRFrTEFwbgP4qc8BRc
UVO/1M29MhN7y76vULGHigXCAbHOIw02550IGgEX4GXoxP534oTY3oqFoLa8r1QkpJJIdcLNWU9h
3ffTsPOYx/yW4/67i/hzzpZ55805jWd1Sn3HLONY9SJDQBg0r3oBmlxIDHD2YeI242tk+ZpqcoJq
ru7zNftoddlDvPBttc+4fWPq3LKhZjLo/e45NqR53qYi3EnfqPoG00vRQAJmxqCoXg2Rgdg3tn3h
ZjmIRI4lfiCkyMJIZ9fF16GaI1jwWnqhICwoxvLzmI8U3knkaJHVCZAEetN8urOZK4nxmaNEaOMc
8xJBel6tXAJ8pmCIuyj8htkr3uuxpcXUxh67AFEvOGs1W5qwPPcjmUkdvwXBR1TrMCWYD8aPN2Su
Afivzf5Cq3mwb1QSRSXSy8hOdxcSjg2w3fH2K/9aXzG/+3czO/a0DDdcjN1ua7+UQKDoS8GrAiTN
pNr3GNSuEoc4/nw9ss5zrlb9Y7Iy1/LbeAFiaEk9/pnmH+UUbhM/1dykaNFdS0Z2nYBcem/7wTts
EVqEMx4mf03PoIeYDsPIWssSkCAK+tAwCXIutAjt6DEYNB9/Gbn508XFESlU33VO98sv0KC/eTiG
RA29z0MQhBcJs2TZewqWBwI33tUUt7+akQ2qoLlbwSGAkJqGcbzPZPNQX65AdOLbVXoMyrO5eHQv
Mpab/EWTtywKWrLyKDUSmH7cJdavGbe430vFrkK+lW7FpHDl4JDxhisG2/enl0/5VI7aCaSfoLP5
idr6kW0683Eja3iMUirBCvWOxi6F7bBnMYeogtxNgqbVnGal6kF5xbzxKp+xIM139yq/R1ri6CTI
rAvStRkeAiCfNM/S5CrShgmA+e41F1HviPUmBv2dlkuSYNLHBDAHUSl4H96plDLQDc0lpN42qd18
6Kw2ZIWERVHdmdfS0K9+y+tI6l9XkNxngOULi3rWOqkFFVfrWX34pPxpWT36oV+fukGgLw5kOuS+
vyUcOVn3S8uNF/ywtsnWFbSUAINLMtPdIhQvR8UhGw13v3VENY7n3+7hoLXLytOxtJaoCHIRuALZ
CF28APtYNvX4oTy9ERYDzOvEEM4xdQcceFM+9Epyb3g2sh47+XG6XIGofRFqAX66pdBRpdHl6jex
QhQ8VzVMij8oWXDF2hg1J+2zy7u0x1K+ntcDRskwxEM2uE+jXuauz0Rx1e8X28blSUD5md1orue2
pP7B7tjgR/ZfRnO9LjiD7HQ0O3lMkhZjnPF5hk8hd+/Rk2laq6zl7c+VMF7gGFt4qRZdAnDz1T1V
rsYlx5Ej2B3BnxOEZRQE0eJFTRrEtz6cDlHNiLuabhj5cFtqF82QrJ58MqDxyzQoX7qheJyh683A
xPEa7MP8MGOsMfRNIzcw8FPi3cUl6lnYgl3dU+Hfv0rdG6SZDixLm1wpSMIJedf47gg0CpdDQSKm
g3MyrKz9gckdQbpzZnE2hyMSDOeuIDrSishaVgFvU//HRqa3gmeBKSlcIw31CpN+LQKh2WU2UcmG
RgCPHMKCsU54wh31/loTVSLRpDFLeSTgErEI65UP+0EWQh+HuRjpjv4CCUxKyjvVcMXpNA+UvQ3r
sYZwFpB33PtKodPhny7TPsuODVlJzm+QVK4Hg4qH4+XZoiLBTcYnZZ0/WV9QUlr8WuRPVlZuoA2H
hbe7w7VtmOXsosCWg72X8bdsVDmKOf8ntQSfi7bhFnlHjxO7WUqexdWGZbfXjstqrpvQw9fCv+qh
zQopVeQPsf6WtvG2+d3tPSmu3JHyQpgUCfaEaPR7vs5v1TRGzAaOhmds71RcI0CJnbu7OEJqfL6/
MGaHb5UCRONI2nKT76AtkSyEUGnIo5LHMGbJsP39xB0BbptLqtV8oJDwIz1Egrrk1ConXUetqfHO
oqQDhlCrPwZkpAwsun6Li7taaTtFMo4NuaYerX0UFsMSTJeoj+kVDBC2579DKPDL/vg0P7Z41OsH
DtzCmC/UkEFmSkY2n6C5pBSzyozIR+8p7AWxFYyc7SoUb/eGpBF4ptMMf092lC5j0TCLKI/20wGT
+3hl4SZKLLzTF75rP7SZIkVNKy9i+XgoOQrHGVTX4Tgt/0YJYiocmAMqd5kRw5UbjUpi92zitRn8
NnFRim+yVQ/0HdIQ7x3le6SshqSVZWyrrnKURl3wnK7pXWhp3XF/Te279WwJZfzAUMCl43K6OVHi
kyat4UCyS7/hZUzZH+0s+Z41GVAPCnf4Q+vauajoq8HAsbjKOEBlHElLwC0kBhcbuglTqyG5jLds
0a39cBTSxu84ASBmqpsf9j8/M88QK3Ajk0W6Q1y1QAQgr/P1zItcTQBmVsL09BXNQiqnVVoNL7YW
u8ywKOzRLLZYn/JsLs/9f4l6TOioZp8yLYxrLVIzmruoZONupyWjrGNaETQ/wEmphLkJBBFblXpZ
+4NcLSJ1UJVKE4rBAfRKL5Gd/lFymXrxd8lkULLcax3ryU0worvI+c36P9OhZsk2/C7/MSiIGaw9
sia7paV1/Pafi5Zpn8DoXeiS02Ydm4jan+gdS03dG9hCfhboQ+tPe3uB5RKHXT2gq1SSKsSRpoW7
zUQTE6vtlwRj88NJAlPanMBz0B9QmlygLW2J54y87S6putsvhzz9xz1S6IxC6Zn1nWhZa/Ci8lw9
J8a7hzQ3JYG7CHC7xky52P7Sfaqy8hUKGXajQKVFPdZTbXTyKNekhikMmMA3IL3ttfH6Xco+j7l/
r46R8LSqJRa6H7lP8jZb+5aGG8507QJnviVE8VhPyE3aFCqOStx41hgLfgDWdoGTNl2i+iWBPbS2
FrLBcNAeqlDM+6+H+c7r7wCEOOrwQ1RI2B76nYgr13jcxP1CAkiVzo1jSUzt7KxOEfUAVpCqtOcJ
XFrgIL1tbldFFdM+4xnGGn+8hKmjZZhuQlzESCqz7bRMDWvMVdnwQj6JpodV0B3m3/QZapbF+tBg
dTKO8wriMLeHeAF+FS//ipV32YR2bat+5OcSjGCHJUnA2ddjYr9h8d1ckh5WNzdY+RYV5WDYI/Oq
Z0dr6oo+b0eXgSHYbH49znZv+/m9hRxppYUyBJ4Shnb9z3xT8HeF1DotRvX45QFZox/9ej6OPZiY
vJgXNVnfch1EnVHBfKtZFsvJrO3MhxSD8p/Un3PMMm3VBBKXx8a2PeNYSDPTSt1qzWa0qoE3JeIz
ZIFBLnHQSIsipzPtFxOd7W+/LAWEugPe0P+utXIJL20ujPmZ7Fg0B1ozfrz1QSq+3Q+rFP+QyVyP
gcm/sOZpwcyj1l39iGrEvZOwVI03KzLCNEJrj5BhYIvm/H/qQQjzfAbALPLuPWXgzFbmVzKW6p0u
LEhU2qtKQMyx1+HhV3PisYV5DyBCvEN4SPuVZbGen3shDLzqxytJJH0flfcHffjbaUOKlPxqyA99
v81AhJy6iBOdzaq000PPmwD40SikISbs/HzDR3U/hArVNWpcYBQuND2qKYv56fXs4Wk2fSvYd3JF
iFgL5Or6+PSbib1Kg6JFEIUh7owOr2OSQ+Z7EpJZL7gusNNSa6avgX+odkHdtvdob81JPSjfxta/
eFWLVtY3Lg46eCDBnQC8ZwO25m834mT85oNaoctw0xaPUvv2muBpQ/GhcDl5xDildW/G0VY/PVGU
WlYSCbwkEjHGMmIQcwFG4w+z8PqHe126wkRpX0jYhFOJsYuq7RpxiPeg0coFBc4PxL+7dCLgoA5I
Suuz75XJ5PQCz4tB93OmvrtwF7xuIOcyN7DNw480oTD0g3APujK9hcrNplsbrtEHRnbawXJAn7Hu
6jHAyV87wQLKCxGyTLre+dkkoFKfvKRx6kkcsCh8gEZzPYBW1VUNwQP6krug6Kv0a6PoRUVHYmjy
D0lq5tuCeI2qxDOntQS6QPN4rkfGaQqHpKAE1ukbvbp2L10NAhtzq86M0Eohj5ycQbuXpHtFg4B6
3RqzCs4xnp7l7Qh4Weoou8j0lXO8DDWkWJmsBGsbhAK4/Y4Y9Ph03HyXy0b5AxBBU4D/8LvwxfSr
xFKxymMnrLRvj5G2/s4VWwSFux/lS8mXp0EZ7/akHWHvMWbiKDzhgsgJWa+zdh3TH+TNAoDswQkS
4w04ZFPNp2W4u0JS3NQU9f6vSsv97uD3EP3Waj/AmdULli+Hob9BGubL2lt1iHVOmFclzXcsdWLy
fk8uWmG8tYCadGUDNnpyH0SrfjUxqXg//IJEo8B7Fzk+sg6PKSlRS0x+Jzq+pBTmhoqyp3fehgbL
++G6RY5ItJc0sPEGW1imDxXDOO6cgpoEhUXA7f85o3abbQXhcV+oCpWRcOGF7BJRy6n8CVNSQlB4
FIa3lKaoFlAP+LX2F1yoEjk3jPTU45ZVXEw/BGOoaSnOjn7+K6dCS3bkMxwxLffpU9yGkmEK8Se2
NKGRC00P2hTX7oCBYKxvn6G4KLCeM+wkfWdqqm0zM6UH+kAzFGJBL/qaw5k2pVpTE2CehqrfToEJ
ydvVxTq6oRZ9D90sJpSAJ49KfgyFXJ0+xYtTjU/1KbETj+wH60YOvxx1ngq+wjdRuc1AM7th7VqK
jab8GT9PsxFTnBsZ6bnik6W6EOng2/rtguoiYr/CFH6Mb/218wIxtWGWfbEOc5j8PxeHcObPRT8r
ToxQoI9UxOkNDgU81fV6l7Tvu4Lle6I2ueCO0Fmn2ufmQFiLhUuF8S46ebEod8xRl64WJnX5T9uW
JAmffcfnvwn/aKNIIKgoqcPddCX+x1gTqW+sbj8qEAD/aUv31HnNlDauCH+PLo4k1Qa0rW4CcsYK
f/D2B8n8IDmeVFJuw9EGLrLUOIES5chfOM0d0kP4qrnfIuqLtusbwHiMQK5GPe3FL8xJLaFy0/wy
jHseAsf7MebiJylEIFEge/Mx/WgApDbpyQh53juAzGh31iXBMyizTqPluGKWrczjitmmgcbp7G8O
XOXFxrmCeOiKYPSxIBkz5qmKoBWtTGSLgJMr8WlECrZRHobIpJ0nydoRksD8Cf9FsgEbMNHTWizP
RNKkcR/EXDjlEkvidsm58znIVBiX2BUbKnfJpdrhmWKbO4QynSsMoEjqVcSDOdIZz7NNG+Jsdoit
RNB6rdVb+T/Y6nSuBr289CAUk2hiYCZhH4KOGZdUYr4kF6N3R2xw1myTkBvD2BfB6O+UL/R7wnbc
HVQ6W+0I/uQISalBoffRbXnRDa8fEH0gcaayoXFzh+VI+32BQu8fpF8wqEVThxGeunVf1BRucwtV
4X3rzqo8wIPL5/7dfu3m9x3EQe9J8DXSTl9wdi8qssmP9ZR7m5aBXM2A/iTxZGuA2gxCTeFHoPKu
HYaiqg5rJcvFrnPFGj+h1oaNbr0HTtbDFBnXjKiLHlcAA8poSDIJ43I85mBaj/JVTp5eyWQCY8sN
C450CtbYudpgRP3Eb9w2G05AGOlDN/pmV2UcB+KF9ZAj2cFt5cdg6olOsf7A8JRcrFEWS0Nszu0Z
vDXZvloO7HcsunAIIKDmxvQ79/NvMeVDw2CYWPD85NRTOutO0GfWjpUpU/dm86+k1yfGnZTOup0E
OTyHDZEr8oEwnuJiSrqdOOG6vPt7QXgzqk07Em2QDwt8CS+EpV8f9D4vWo4/6tLQK0ReN1RPhHa0
j7e/Qv3R4OVqUlR8Ao8+1FBtfxFq4s9Rxc5nQBAtOV2c3u51xgaww1hNjtbBITN2DmronG84rXNH
GcUMcfeVQ62MddXKfO2DhSxJOO+Y3GXrm5b83WKvKJNB5s1oBINw3AvmOKLdKi+SpBPe2RBraaKu
8C4HQePRyYJZUfWWzrS6gLkZ5UzuWV9ouQno1q1OPRwi0Kn5K9jyZ8dXbqDiUrbrMbrPptrByrD9
/VDDVBqTk60LAOazCUzm5m8Fy42d8Uj8F5hl1eVFe7/Zu/BuHvsRVo+lp3rF8YGK/r7V6le1z5IM
kBuDNtZWARUwbFosVaWVbLhtyY7b5hd4tV6Jh+KEzMOD/VUFoP/ILDjiNcGR1ghP4YCIY2RTqctF
EqgjAtV24S4qKcId2ocB/GXUZG884MKvwjdd1aAMxx1eJbLYCbIV4Uem3rDM3JSeSnP5IxA691KX
y4q0csx8KG8H65Y0ShP/p8IbnL3CfgSx4Tg7u/Iv1F3FVa9V2Xb5LeWet1HcJLxElnXps8R1Ao8u
Urxf9hLi3FILnQKbuCjyjpYw2OFEoSZYJCkb8PkIbllHA0K8wfb+8TkoHCs49LLoTBK53sYhwKns
V2DR6m69cQ1m8khTlqCsQQbz90D922FVE1G410pztHA1Ko10DDsHBOoI406un47ymM9pEhXmoVRJ
Vpitz2NBD4WsfjzV5RU5CNmpxdRRQNGtxKoVaMe/oZ/aqh3UzrtAmWnWbppTcrnrzv6HRKzoYU39
RMvFl/5Ib3FW2pA3yU4JJZ8aVUbUQmbWYKtk+1McAB6iF2CflKVTRhJH1KgrWHqUnMP1PZ45z+aG
QOJUz+DGh5xEIhBrPqdJLsPdWW2QfaA25L2xwEXtmWdWGFRGxuK7WtDplxsck/z1sB3g/GpzgcNE
w84r6ZwQs8IVEdDHSsOWjmzDTwVBkPcJmWX/oFmY/+/MdJ5zh4i6gi6w8cfCBo4GhVJ80ckUC2gR
8Ei5rpHK4g6A53PxlSOUh3DhG6RJ/d6z5KunwhW/zdxAbyWr2xoPer6eEX3o/7Nx36OAIAI9knyB
TTQ1FtWJhNAoA0vuaSTQXmZAA2kIePnSsNAvObzIBtqBcvMszS3KGWcjwCihKrHXCd5dPdkk000/
+WP+yw1celEB3Nh247Hrh/PWYoAg9+DA1FZg9yZusAvhxEHrcJExSGk2v4O9mG0ecESEN85vIs9r
TAeckr0uYfbcmEg/Bvinb310Yt5GJor59ZoYeBgbwz02mV5Y1eUzppFlXEhRv6i4v3kYV25yFH/w
ogpNAjCti9cZ/EN8ppJ4Ec1z/oLIuV1ZXmSM4222BUzHoGJ1TAqGRVs+I9bAfO+CB+X2AJS/PZr8
H+/QOEAOwVjaLCtPfv61qsPJXlPx1bcK48DP8KcO/jAxZbtwYqxbCVabbrTcWUhVZ3sCwJzrQOzF
iulKQvjPAq8jAIlUSjHUlvki0WA3PxjmEabh3hXGjzzNE4joqWViUfpciNhXQKjLsQ7QCPdjeQRP
vR5vJjzzOSCg12zgaFAleC+60aNTPR4+1aJxQLjr69zdChK49sh7b+L4QeiWSqxs8Gp5q2dnPQHH
Z3wFzJIi3UWHLc0YxRYvoeVu+yWhFsFquUWzhVQc4mqONMyx9+c7Z8c8R81erFscFmak6LWmxyIB
zjRuC0p1GmuO5Ye6s28zg/B5pnYe4RrQDRrUaFUDgxkRZjFLcrd8abwWr85zIflJ6JrSWfuo2ocv
Da4/y8mHpJ1JXxrvqXP4iUdBpsIaQ42AQsz38GhXuIAylb+lYzPPmya4sMts7+UUalcJZMhV/1IE
rjTkSXvOX3McTh7cNoNaqAzCX8Oa7zGBCCH/CcnTuDPEbH0WrpS16dzakp0wn8Gvss7l1cJaBjct
3EgaMCzJQejAjim0koS6r+wDFfpl37lbn3UciGxU7lRWjEw+LosZvTU3vwnt6Ib3yU23tb88idVW
rBVk1nrI9RNPBOgdr1Oszz6VyxwC9KSWjWn8ZVS84SjbUhSRy0VVF9LA80khI6YgZ4174U8KJ4XG
7m1AddECRaG0YWUs4ATVmlcd2DT2edovBkuUIArP9TIInVFzijIgR9BVAHhqIBjRFpqmZ0LnXsDm
g3WTrydv+kpDXQkB5K/jJPoReBgjBBja67eUAVLpRthQGh+8jYcoyhdlccHcIuYPgvIXCeY8RZxM
JkPEpoUPQxjemYT1WCURHInw+nacgh3hVvlDh4s2bycuN2CD7TTlw3BsyW0kWuW78o3Makwqds1U
S1aM4oVPXbaSW0FLlPObh3ff2+9lY1lJsopfc6tKTxqtR4gKYytZR93Rzs0+Fs6wVuaMSVX7R2gy
kyKdSNmIh5uSrwwCEEDxkKvxKFUJl4KVBeLZV3T+v7+eBGwcc/aFbFBn6UOuCxQmEe1WwXJq6PKz
zB4RzzvYlz0LD2TIFfWpiB9fLrJRfugl+GgHhoFFdwBerK/YzgXG5wH/DXSLciIOsXCmXNXHIvpl
7axxnecSzk/QMd6hCtKJ+M7pgjqMhLvvgdTDhi0dbNas0XK5Uut3Sf+dpY59BscYtur8tc6Q8DTF
BKZLfTTH3OYrR2joj7Igc2yctlsp7mImi7cgELoKsl6lsLx0VSebf045FcwKxboZnQaXhb3Bw+i/
Ji3l/rc5RWUWOb4+WnoAAS8kUdzBFYzqtRQG3s+BxLgqeDCyfFmgI44BSaADsZqH3qpi4FIuYwkI
/cJY8pCLOegZUoMdrwQOHE1F/VlUtxJP1adlF9N3C+zTo4mYmM2TXOpunZiypHKrfS9doWOCd4pL
YrqMkN+QifDeg94KGRySlYg6MaS9VdtFBdPC9N8q95eVRxzP38rB10bK9fFAlzzGoDkrUoLNH3cO
2zdb2wrjG45+dIgK5MsPMYyQIGmJK6I+IAeauprZN5Arc6O88gl9jv4rtDHrAT7KynXDorcyMLUo
YeJOz+VNHN12VuMUXtxR/iDGpi44R5C+QPyT6oWIXqchbpo8LQJEjxqwZVnfjS9WvmPQAKYXhKHS
e3dpbzbqBXyk6PoFHko6UvXQzSFIjT9aHBQW5K7pb/MmYvYA4SaMzEfs92B5RcY7pxcKF3LR6eo3
J2IPRTOUhdbdozzzci0L1YHR/JRQTcx8jjQQbFceAsPPiOcjOCGvotbse7qqI723e1qrXkyeH0gi
MUSGf256g/BWLl2L8dVVKZSq5Ctv6q/+PahTsq7SQ+qQYMgT/7dYgVPDXmj+lzvRMQe4C6EXtamE
pmCIA+Gmb0MsYusM54XcM7h99d0pp/yWVPnkfDB5M4mijWGHMwlpKBoV+dkiKC7RgAaX/Vu+kUIG
SpGOnprKqYaJ7LIYGtjaYrA1+EkJO2L+aQf/20171YLBbxIii2lPTdZ5Zu3ZKpwyR5lN6CTjL6OY
IG7iWb3ioEJlsQJ9SuNRt3vWqFvZpbsJIT+r2NbCuikfPdMFF2R0GX0XJ5wLZaz28HyswUFatHtQ
5REBCDndDMrwvkORUf2OK6MGv7tK+EbTdeI/to1FSijNht7fWDykCY3TctTq0f1gJZLViw9DuoUM
00iOdBVovRqVWRQPSzSMU8JqHnFtPmWbhE86XUgjwanObrcdF7o0QpZXKWWRtjaogXhYhkcYYCUI
gfd86dBsg2CeSIHJHK33pY61sINmabX15NZme1+kQkqMR3A97sJfU5CqpzyM/G5qayg3TTP5AYHu
WH84bkD4QDV6Ch2naTjeg51TiHVJune2OO0skdsc7u51wrO42bHWMeQs8XP0REji/WdoE1Ta1hGo
uH9+IAm67W5UA0eR733eViq19SNaG4rYo1YNJSHCfaM4En9BR9kP97h52U84RmzRvteXP6vcwBbD
OEH2hIIKdmQGFp/2eFTyfllcPmm9G6KyBpreLBr2TlvixQ3bUzKNOASyvaAmp57+sxbzQyTMOq9d
IQa4ltYbFp7W6cfi73IB3NiUthYvcYcLnR6Bp+d43BpeFRcTZ29p3GybONUMNdsRfwsoSrNz3yvM
jgcS4ALyOf6jvn2JLrQxRvnLjY70FpuKqRQDbb7a+0W4d3Tk0olS+m3WZr1CnTqgD95l8xhadN7m
vMtMvrfd7OtjbzZGIGm660HBjLZriJ0xs5X+GbUUaWi/Yb6NfI7fccyuNc5pOZhJrldyBzOXuull
Fp/DLVH5x0JF61X+DkNQE/U7H8f1lxs80nt7tB1hdhQWR8RRKGGq6g4u7j5y5GUiC5nCAde/5q8Y
b1riE9g7FfphBYJQWQUla1dxEXegYV8b1DpQHJ+NLzjl9CkltzVqxSeEZWZS2Nu+aL98mji63VIm
dq2V57VIhuoi6C3oaD6ZDkmXa2EWdM+VPCuIKx+pAQWrthmH/sNNtFRH//8Guw7DW8+TFAQBfw7a
3TfKea3OoJ/zahDNuuSJN+AeIor09gyyWIY6OjicM9KJtxFrRADMu6Gwqrcb/dRcC94fic2PjcGN
loCZIlO1Frj1LQixFp/Ntf8zqzfmD7ax3/jzgrcqWJroYmA7bHOEHrI7JK0FvqlF/KN8LvrGlvtI
PcwvodsyiMfJps/23wtVspvC7X8ywSRCABwj7iTEhEt1Jd9AUf85IAcdMhk6gfBAUcznc4z3i4tH
upHQNVIfNNiht5Y9xbFFfJxXtFBQTfOr+ajn14UrLs0Ql1XooPScwV26x8cEAM3Y04koaAbuX19V
wacP6Xs80tlJy9bSu+473N7apiosVFmrK18NdLoLwFeIaWYQdVOhL7lirb0U3949hfR46x0eNVv0
+PpYegxLvDRYo6ta3zooFyhM6HEJkxJu1jz/X+GOza4VGOAejq2rspY3avdRLFaLZfEtdZc+ogUr
zNdTY67ErAfZfPnIzL/rvYYqkmx2m/Lanj54prxvkWduMe19UsmaYg4nL2pWkbPX2iS0bPwk/hAT
BHDrrVt3XdMzbWG/bgmENVN1fKyx/UagYh68NnOqAXNhBAy4sgD6L6UY3Gsn9cihp/9nuExzxyPi
N40igen+WpAbjVTUZKEJqpROykWTXkm21TiwFmKiknQhnbMH2ou6keLtvR+6mABiYx7/YKez8NIg
7wyjPbQwnuzcbQfGtkTRO/AKWR89NGzVRAVLK0g6xj1+VRTLrZXtYkgRRN/oXJ9i0SpIe4yP4ZxG
JG6JiqcFNB1Yf690MYrePW53n06v6YqT2iWyewy/JIbnoWHktY5oLDbSiKaUMQJv4JvAqur6DY1y
qfniUXjSUzdkX9nLcHGrkUafdKPdxhabdRzL1w5F/YZDG1MZ+Sw5nPnay6mP7grI+fkCbbCL59Jf
eTFZjVSY8e/E6tjoEem9VYTiXI7ADk0npzRUJqnq0l1nsJr4yUyO66nYvHt3ka+teE8JwBIjNaUo
vtAeScUTZDH7Wdl+NXsRdA8+d73DHQnErFQWBXYWthlT9QtaysjtI0VjMSJr/wp0M/wfrwwHt6ys
gHFYcoSou4O6sQsB+YHuFNOqeiLf/a3gVAiyKGPGucTnMe3XZOSncHtWch2ewJ7reJNSdeR3yddS
Qbt326TZv86/XUmQJqdLM8mCpMMBBMXFrYS/pfSPpmyiHdcnLrApTWu5VVskzMgD+5xdjXjILV3C
zlTsIn2cRk3Tib6UfSi9NT3cBIcgoL3yiNooe+Q7rRQmh6Vn7EwaP+vek6DYY5pcTYPRYymNjkq9
8yIssVKcFvbWpp/ahN1PFnB/BxcWpGETAhmmc7DmElQYpx2vnARnDH5OheSzFojLV5ybmkY5XCtX
eUYFyYiw2LMNRgk8kZh418FgHr9DHO9T22dUv/p73TEBbAsjxbIg5dXYdRWD6almHkKeVqYIgc0e
EafXwTqbj4gf8+YNs3C3PMfKx07Bv//vJZB/6kHCQuvwfwewhk7IAWB06I/BnBAjnWlKk/97H489
bTR+a3bKvYxKUib+qqb531cEdivUCgghKt744eu9xe1eA6woOUvXjuz8pjKDlfEGdzu618kTkLnR
0sc6/P8cz/DiAV7j75pY+1ZpoElwDTD9VgU6d6mu5xzK05o933iOG5yaHt8jR9coi/aTw6WUWLRD
Tjrj8elJO2zlDhk/mLXjVMQxbkou93b38JcJmaENsKN7jYjeODUjEX3kbN4NK/C/azUJGgeqGPgo
wgxYyiQiFC0xkH/fzabwUlH7oGAymC/F/WHd2OhXlb40hfVcTtCR8/2jgvu/YtkrfxevydXui+y8
82Lw0ngUHe6YyXDI5KqD3xRC6pSLKdNChYVueNtWkyDOmvepSvbgI0mWCLSBxhxN62VVL1xTm3T/
dyVPLx+DbGt41P1cAMwr9LpxkNl1feDP2FXMDUUeTiToE959cDqaAMSoGq47OFojr5/h0QOJkCBo
G/hLUMFo2CzdO/lUCAplYD9FTt8sqPyCvlAE96f2pwEfUL1d+ay040WrYZTwwsH0sKjXi14lcRrK
8DmWPHgEqTrI5bNLksc/Jv7CPAOX6BxWlIktbM4CC0nAavxqOQ5Ht/89hHpHPEJu9r60jJbbDQ1I
tYNYjlHdEJzaHVLXZQ76FFDYcFiAaGb4ZbnzN4SRZPjaXd0tyP9kNYJfugtkl2aGxM/gvNotQdHs
hvqP3aifGNg5TV0+dwfG705YSwQsvW1GEkMzswtVNrMT/JkjxciN5oMIUZguqr4gUXoJXwsJkODj
JxACL1gQ2eeSH3eau8rOG+OgY34IoMTbGeE013BDaeoKWICIREtelmG6a2E4+tzMSlfDOYP6ahIO
sDPI8BjNusj0EnrVdt9ghYTFBRMXtA3PxMfVfoltJZQ1IEpopQxIq/mq1bgQdWFDhBgUuQxNDBkW
SmZJJdv0PQiFb+MGF6R8EiIktUyDZJuRK0sTajIW9PKgisDwO2nZs6Wd5j3U+AOnMboZEv3kGkeu
+G8GVZ68U1DsNKbjmWC/AsPEqmiN2S1YvI56iB48HY7grItP7m2UMBFieIUYphafqzSN91tFXA33
Fx5j2K5eI/E/N+D4kdcOrNUgN8ucLDuJ9NgytnPiQyrvhw26156OYNHP0fjAMLkSL5zJZ6SDqgkE
DFGnEvYYRcYZYYffCusrFwjmf2AmkuZVtVDGQDuC9+gWscBvXm38pQ+Qx+2S5sfJfJuEAt9o4oGZ
9gbTiwL+wfOBIXQzdi7XOPuc2LIk03Jiw0MFc6CwVej+7Xn1Wml/kONGOtcIhRF8OpP7NDNvq6NB
sOqqQm1iAF147uqaF6eczAsiqgEXK8H/TY7P3fzC3qrBf5a30QxlISHGxfr94mOjqzE/Vms2ox8u
tRFtwPCyKOxwJxnYekxrkQ0j4gRXuvx1NIDpCoosMY3tBgkse41VNFX3lSWKDSDzre4vx0X9Zctk
GHtslFK5q3YKc03R53+h+3lib24E2OcMcOUOudSTHvTONXvFWY8NmVXwT0HXk4rEWfkpbNnQwIQ9
u1uE1cw2KjDTvXb3bSr2fVcX7FqAG751hv+mdBCVBqIB2An3Tpkc0/OFS3vuo+FUtzjQifnxgplr
K9WUBxbO8M/fiI4LdPARbSlz4X/vlJNFynsAS5ALiHRC5iY2DicQFuMWqN0naVWollXdRvmGTlBj
8hP+mKvKFalKzwQvmStP3PAJdZWQeEy0DG1w56qbTRkiT6JPKrmrP67wqMxFIV2hXLrmtuh22KfN
lAGhF1sOOAQYLgLAB00mcB+E3pS0IdyvlRF42r8eq45xuSfX+qY1wuhBD/ybYEszZk3Gr7Qb/vSb
3sZ8dehDHcYrR9j4TJrPVNVC7XHsyn3inO38APvSb8wvy920IUPP1RMZAzhx3XPbrXDyE8AUDOkT
gL2vU0n3qBaxzL25BYu1M55ChYVNcAOQtx2pPCQEdi/PlUCsJjowID56E5lQ97lcJ5nmHHbZKfnd
bLz9lbg7MnXL5kaMAZbLUtwQmjnGP2AabtKiaMSN5m5vTihUmylKmyVVwivWEseT/T8cig9hhMUK
r4Gt76c1eFiWAUmAxHz3qUH+sKr/D+Dpe4w3j2pOpwMRxCe8IjUvKtnZ6dxi9GJTeJpH82hLtOkJ
7mKi4rxran/itIKwJkKGtdToRomHHR8HSlG3g41zc0n0PNvUVURXU/YnrIAuX5ABHJZoiB1pxbht
0AFouFbBPv0flr+xw1mMYjuyw3gGheS4kZZGU5ovYqhiD2AzBhd1Nar35ahf9NNA/Jd81JxihFcr
icYsjbCLrowMdi620eEuSTpUba0ww0qTFf30lAegssLn9ymd5Mi6L6qu49fuNx2pDQSAEltI0vbr
EVbCv12bS23UgPmZOdjIZ9JJGYVo4GceR2gTjuO/7ku/pYEDkyKIcqY2RHiRmAYVp+XVjDuUaUzU
5oY5cgA32a3WtlCAEDf5blz6Q/vXuLMk3S17RceWOTukzs74tX5ZAhzBJK/xXNM5XSI7RowiyIMZ
Vo53NsYwTkd9qP2vQurlDX5PIYVYTYO2s7zbOsaWJMvw/v8PcJFw6ehmkg8M2eFv5LevxZr+1FrY
r9fqvOdoUpoMC0kzReKpnWeMbz/EHHM/q4o+HFfufVs43ZplJ2tmCG7qg6mivF+2eyw5ncyMIttw
j12KFhRj0YATKNO/SOpUkzvGVZqdc+tOI6x9U0aDkXJP62LhKba/eJ3yNew5dhrjhjZ27mObNjBB
iKjz3eOW2wG6oQ0zY95Jy3EYCvDH4AMwgG9Yb21NkYGJ7eHaN3GN6wRY3epe3i5f6kdQLkeUGOxJ
cK0rwtmx0kz1SPSZu2Xv2t4q+3rcoHYu6nBLtWp6z9XmTsEef0IHAp+NysCRCYXYvtjWiTl+A1GE
IPjSrKrC+VJrmB3m1OAtY5yN7YJmkvVG6JvPrIPdJ5V8BnF/dxfGOnepqz82WMFK6uHhGT4LNQQx
5nnqGx5z0tnDZ/QFt/dRY3jxWh4IwSsj+Qm4AII817ZqFy7pOOguebpMqgzXn1s+9nbwOfdI7xW9
1Jh3yV/FptxiUj6ruCK+mEgoJIbL85+fdfD9lLRli+wGMF74MDrziIm4nOojGzbIQr732gadhAzA
+m3hXKPalJpzzRwwkDUINX4TczrDtUjrDcDim16rpW8uo3V8XEqgS2jZXii3Y2fdht0H5T0wg3Xe
rvRLXDp9jym/pFsSizD2oBv7GDjuMpfMjjORcbOBrgPFjwxZDXp2tkkUMkiNemm9Rv7PBQ/zHYYs
VraVWjuPA1qsH5bIjKsIJupokEOUGzp7BQw356BkPsiPU5mI2qaobWfpybWGXe1ZqSEQ/d7o2+Im
2/rHdHVMxpOtKg0SIMIAg52lv8981/O9L/MyCNEm6B40nNPZz5/Q88MJINayLZzTav23vh/st2Kg
ic+kh6Sg9BGxV6LDeHNQowG0s4khKvCDT/fE1xT+G6T5H3PIIKZiLh9eo+BQNZtnaDLWxuVOdNSu
G2itlNXh3f/D/4U7dBYShuDfin5SAlHHzBKAxwfko0kMiP3YqScRytHdm8/N8uGhsaTOgWF7uy5y
nJVQe6KQpkFtMJQmS+JHiVN3qdRwxlXV+6WVRv+1SRRj0gEoldBE6kddk2VBv0YgcNY3CO1UIdj0
cQTbbOewo6oAAn/zSLqW+pZ2eeoJ5Zz3pWon4ZTOQaMztB0zbUZQ+r1SG0JbBVTXItet/mtoTqve
LmpLTnAhcbLDIpBRKkoKlqv2hZoqyNvm8O1Qukmiq78OoItaQxcFZpTbYxVexT4UVaBsXEb6qteY
d7QTN3jHre6+z2SAeCT+hh93JHIUuL/IYlhJwgYMRaC2Lc9PW3lFOJSyVNTHHcQXY/RjAU1YPSiJ
5ui8abAh1Bf67DIAr0dmos16gcTnODNa+CSgNCcXQ0/nWw+9HwahUdF31odYhiJmWhs26cOAb9W2
ZAuBp6rDD81/mSsiLbzQ4cpjMrRxAtu57cbPI2DNZQn218r5FIbhXEKI/S654y4AD5dYXBvJ//OK
pfHSF/q9icTTIrNj4B2XBaWbqb65nV49JoPJrQ2bJduZjfFrvGjMUbgP4NwZn5epPXLO0mIWpSj4
CFScYEMAjZEB5rZqQ6WpRXibGg3heUJ8bCUKDKsqd+1sxxKEu+3USVnnn/QryqvMPHlNlc2M279X
7JqXpRmbPVdGHp6VoJDswHwfQZEIS6w/8jggJX5eyjZQVsZBXfMTZ7qWBh4lY2jZ/lTx6ZMzkeb8
qL5l3tQGeWewUrWEK83yIY8WT5ASMj5KDcucdjYrnGpFaUqPqW0hkcQCJxpGcfBFQixWpZ4ELvn8
UHKJsHn8E7Qz32o8HUo3jx3Eenan/SlIcWHYPwvJBi+9RzLkACeGymrx7MNv+lWvGGB3X5Vb/5VU
U7muuPIkXYLzBWPnSwEdxpUcaa3yWxGwgLKFIWEIORPq2A2Z3FVL8TJUULskdN08qkSsC6J/3ePq
F9xaPfEdRu7TkStZ/xHS4xQkL9NV9Na8pq3aMVL3aALd57QBt3iydinX00IZUJWV9exsyDCTVLqV
O3jHAl0NNv6Y7eVT4jViQ90K6LAN579PNndVHRnxXc8lLuLERnuu8K3JpfaY99PYK43QGHZg5qJ+
rnHlWTECBZTSBWRWVFtVaBhQTcU4UEv/wqEF6JYZrYJfja1PESdecbuSi9dQvM4NKlbvQdtQcXSM
ifnOSoORU8K0JRMSz0zqr3Qad1i6tg/5IAd5lDr18uUcufHbIYhwaPuBFDwXvmNWz8H5IEIDkBEi
cjPc04bpI5o8fj167bjTw4qc2u3gXJfD3c6LCcbYicObi85rlc1OaAOoIh+UpmxBtcKH1bV8QQp8
LmkXJsdWjSOkRwdjBb3gqxUEWCJh0xO1tXtTdqtMwWciSFutcrWtFdgUumHMziyAwPZu329rw4qy
s4JwCIbGx5l+h3DqYndWtR5TzhdjWyWOJH7hTtvuBAKR0KP6OO5729J6PPkGoK0HYiyhYSNf4qiv
8rxpvY3cO3bz86cMUeZXRyeycKyHl7i3/lYuIkCJcCQkWy16DSCTBEl9lmNlPxZ6rbYRjTYKnAO3
yWL5dNyDoqaO+2Ur5ATWs2peycHZruI+DE4KP/G9cGVoVMECU+9rGJQwZ6xhDemM+Q1ihPRxFT6/
bErRWCuqsENyTL722OdZAa14rgo30Q2OZGVf7g8tSnQLy5PcUK4kiZWC2q1k/S4F1qUufwjm60vI
BmhGBhRnT0Da0c5kfWKxXtFP/sEmgLrhFGm1SXkmvR/FF093eIX7mo7PWnWtVCZJLDGbIINxfz9s
/mPqzU6jDpvji1Cy02e0b4cfDJx1FRQH/uliAe+f0qYz1kwl3OH6I+gbul1hfyJtJ25BMaUT4fzk
R3GkaWg33tW+1KyyHMERStdFA1yoHaLJzMhaf9/m4AELqOwxuigLwM4QKdFcBN5jRtvls5zi/DsD
kY7GpznrdNquKjuR/fkXGdU256+ZIEIKa/0Oy/WO2W9rPc4fWJ/jJlee44Ys+drHEoLftBSlyDtn
3jyf5qs33fv5Rnc+1KC5CxZTdDfXvi04MIx7TLT41v5vUctO4kAcWxjGeDBtA/LV3Z0YQp3HcGpH
epFmoN/TCFe1VP/YmKWtyzegU5x+ehho0k313oX2poZpVTWArVWmn+1py5Jn1KtY+QYqMOY+KsQo
jstu9WMb5pfqbN17yWWX7dONNrEFS7q4K+s9h8/sbaG7PCFCFrv7BWXK9xNd/OWwCDQg45vziEna
9DgWGUk9wUDwp4wnqs88mhmVynowbZF/qdUV1GA6UnpM82rhVXeh3fE6BINdNXwdLVvQe7vnQEzZ
wbVVRM8Zhh2bMZ9wWkJD2YIKJEnWpUsJl0v2ju+JKWiuO7mr+co2n9AtaVsKt26M65Zt31XqiiTF
kEEruFy7epuVbjIj8MkDKukFowNWiIu5NYgIpeDrlOziZS5mX918394EEWIlpqGGsCz/Al4RmUrw
pqxhMvdyq8K0Ogj8syKDTLbI8+yoNg7t24H+XF0bDDRxgyVu5wXvfzlVb2PTZac6S0rtNDtOlAhT
0ZzlasVu+pprQW2tUm1+1CFQn+SE97ttqBqHhvYKfUb8GjbYC8CgaEwBTtOtCHiUzN/eVl5USE5X
6PfHHxvs1vkE15L53YwgsnKaVwvRpuX0AZpAJcg0Rl6l94b4fK/L8aEtP6BqThE6FsBs/I/vmyyE
1obziGo7hgshlw5AkXWZW+okvM7LyVl+sm9nOPwAdrW83frpsvBCWa3pjjm+Xc8GJ7CsraEBVzVK
bnmgsjHRQrPtPYQE8GCA1TkkYW5eBCfvzrdNu3bOBR+JkhWAPh7UhhWrL2CNqXdMf32+ixWt4boM
5NUKqXaLe4qOve9ht4aPcGMKcc2+di7N1ZxjSPU/YCf8qOzFmyZSkeChyWlIugksPbee+bOyae+2
87gARZFK02TvcoKyMfkEG8DIN5LAuBWeHKa7A5qg70bYTgIj8g6JZf/u2t305oQ3BpqmQoLCQapf
Bww92IXPma17wifrbhtTQ8mC1UG+GuiQiZmHUveOcsdWXc2YjcAWhLddw2DnA071EbCOipsOvSbS
/gRCpTZT5vCHB/25X2LoNjBalCnex5CZCtSQL9llrRFpL0ypJeHzuTThusI7QdFovGM/6jWDXa8H
28beF+js1riFTI2qXdd0UumwM4j+gloXZaHGnmdFwBgEH7D7RN0KlYPkjLXFJI0X8ZvhQGYmtZ07
WevinmxnowuGMyju+3UeBBa8IZbXR7gbfOzb+k+83p+XAy/PxX5ILCq4SOoGgDTuK3wcaoG6sYQN
TyKQSiqSOZXFYKAQ5zmS0VOK+tl1EO7tVUPyLguvBbFTv+5++UGRL4k9JiVqZarCTDfyjB5GZvh6
EpNqBmxAHbpYLy5ikvNJsNyQqGMx/0bkuKboDNmGdVdrDmL6DHFT1NcbJg2uqWrDroH1UjImYlnt
OZGzjkV77M1XawBvh0RFJvKIEuAuGMC655HZoIv6N0S8z2M4bjZKd3H+XkRtOH08eCXpNkqKWL3e
/WBGRYQBQhd/+fwfMCySYLoWyMJXuIM1NLV7PDkhkftYPuB12e4ScOTbihOdR4bhcZ+kx3OVdca/
Avru27huDwWn3sD4w0owfn9PWbE1UmxkkrvTEctP+QS4oc95d5fSsHd5+H4jmG5z6+jVIRsP9ttd
U4k+BYfub+H7ogcUN0q6WXQT9gM8QLzUvsAFwohLwG5UqDFSZoRXQz5Zv4MsXiRhZ05uLGyAdlpQ
uvGpBr0luXNAYiFDnnD/CDNrf7YRV9ocLPcNbV/sZE4ViLYZx6Diqh7KiQ44NN2rfQO8l5rQZ3sq
G3rmLY48QxaTieMWcMx8fzAUj7X32Yk964iamu7FrZnUtFJU5QiEZJ28oorxzAUZeBspR2AyJ8az
Y87D4asHM8NGEZUthXSJ0i1H5mPIWEpcz9w3EiNFFuEMXkTnqJPji+ljTFP+wGZMDz3+bEQnFy+S
StJ2tfnWQkFSOQuSKVWirfYoF9KbgpVLI1zPBqQOnZM0jJ/yDTSMCv34JaWjZji6lwrD44ubSSMY
zHieROf3c2xK5nzhbTG1N1J554DqUqlpUw98B+vm1JZq4Y7dDLYCK64mYHzvs6Uacs40WiM36WNi
pZmseedWsTCcRKLrc3f9U64iKZCSDT2sIWMHuA5LBHBBPwvOqWjf5zN/5EkDuJEoKYqpDpFTEX2M
GmoH5nHbtzSugct67Lqvmb6ro73YISAShKaWCvyszKEXowsmSkAkHFP3FJvmcmi6oKXZUuDqpQ6+
jHWAQgfYogFlN/Gadwn1hJAaOneiI9c+dnNAbX/z8CXTGTcOx7ji6y8yyQKSD34S2EQ9hDEzmCke
3RGwayNJNKhi471oC2HtfEN17iuFRKzkCById+cleUT7TimlXrJSB6kh52It1BcK5Hwxq91dJ1e5
0l5IJSFpdrtPxBSnaBYosmH/nqQ+AbR6iljUu/gWJ5cgDIlPUIhTOHldP//lEZxOZO3neTXmBW3m
El3Vt10UFbvbGKHYeYx2W0zB3d5J0/79JxdzU2Sp2ym6m8dS5seXYK28CVSQDxYDr1jrL36dTYw2
BsYUyL5Let8E7bcrfXK6eOujPPUddZcw5500lQE0xY62jX2cMsvnOOhjhgX3KsBC+VNB+bo0GGjS
PfF2iK+ub9GzwL+6pS3jGUU8BwHdkdd0dGefB2ph7xgWL+Lm6oXTCRKHKxWHj0H68XiZ1h+5HIOM
jofqK9qo27eaMlXUL4pBksonJW9H5D/iZvXIPbwZEDI3xh7OdWTtjNi1lNrO45tipSMLwtiBX8yW
yxXPpCHEZoxkY54RbOm07zKmlqBnTPg3MlU3+dYQWRAxQ8eigS1e8Pi6vRZQELvYNeVG5yGLY20o
CuZn8NhaZSbDTp2hx7w72wdMEbIN6tNpr/UZTvLato40XHaTPA07OUENv3O8D/qJKIcMFNP2fGIW
vooJ0GNPqEVSro403L5Ie5cFK7FdYVyisjWf14Og85zvIMJq9Nisp8GNVFbU2PqNJ+ntQcB6W/Z5
JuArrLSDNPO+12aycr7HR4M7bMaFqdOXZFIf2WSCpEd4AXcJxtstKa1WfEpUL5DcxTX/M6JukisE
/YpYXL+0dD65ZPnEao3FWx5JxZLMcYdVX1URsrGMmR+hAKW1pU9Rimbs4uANoUoriH4E0Z7DZeN3
sQ9sMerh9AC8YwMiSTa2kbJUUSWfLImg4InQEfpasBHxuStDEh4HiczzyqqzrJV21fTbrEb872jB
MaAp4d6Txx8xjpuBnheFFtYc6RDPh/dCze1In5c8iyX7P9TeNlAZGg0Q3ozRybziLzzh3gqQQCdp
kfaCM0J2hE/77pwTnDKmPMypFCe/8125mTBHxxxOhq7yS0FnFctUgZpJsxXqq57MosqWN1+IZgTh
Ge8F8Q96pPegc+KfEsnzfsJyCV4nprKpDDNc1Z33nSY0ADRVA0jQahcZYSqxCxL3kziqziluEfI/
nOZZsJx9jm73GDMGjeErSJDzZgyrGb3ZuaN6kMfI0FGy3E4a1izE7h87vlVPPyf79nHNlknCw6OO
h9cai2XMZRFDUzWA2bl65MSXEEI+WPLai/SogLQj+X+bdSHvzAJeXj4dwPa8DchaayQyWw5rq1lh
UMmWp/iqkvWgmZfxzNW4m+KhZnSkkEld0zyI83e7o6VSrqTiwM6itvEhMDu+3ZzqC/EVaS2IaVeE
YXi/D05MpJ/d7bVpookyWsfOcE+SaMHveGu02u5/rMUq9VTfbzERdLDdCki3l0z3pTVAjcWGfu1Z
ZwRfY+w94ipBs/lI3DPwIQWH2GsH/t533m+gpRx4jF32n5x8Ajnh4NDt0sSienngbkmaXYSaiFRS
RmsIRhRvx2UGRQ3YG+NNI1Lp5Q0BlPh+w04hIdWuxhnJQJR0LxBbjXbsuDO9IBo3QEMTKCWzHy/y
UPu3kmP52FZ3mfQdwIfBi3iU1W1eIVSG3HyEUDswGhqdnzhTLNoQravfKAcXjv7RrW8b9vXD6AMv
saqIsK0yprPpVhpGwkokRzpxmBvXWC6jxfElUf4vKofTwTVXzC9jgW7jm0Crks6vnnIPF+EWa1Bx
a0E39GI+nZMK29WmVJ7TdffZd7/yTN2koZWriKHQyqhByuk2D66C272877c0jd8fxwLFAY9JCQS2
DvuByTxKB+XqJiCcmIBPsTgW323wRbZxMmLmEZDWEwMWoHxloeQ3a4NrNPk7FUVKkrUH8Ufad0Lm
uPj6asxW2NZvShg46lSDpqdnWzMkiWywXa9dzsROVvuTgeA0ouukLGJNqtPLqnT251u7RocFQY5f
W5FFZidlX2CCyxJUVejuiNDr4ZiA8aTuFwVOtwu2sy7fg0tADc5yAbMl/FvuklfTOJE4mmhfgiQZ
D4Bxrbd08OeKOTmAcJzBy5vSFhkiLjck1HTwFzDtAtNjP8XFD5p/2oBpvR4aNHPfCM3R6us4SYwv
c8wJDpFgc0vkn2w6tQEcLELYz5LDvQ7ORY8RqX4V8mWkeJvJa6Krx1WXCdewMgmNeHRf4ugOt+jn
C/w8Jeh6pa15zBzGRwGbRyUV/ml+qBmQCm7qa2pHe++Jh38/JHurbgdGyfPHvAB+jccyPDj4n7aq
VD/O4khpt1V8QI824tiq5i4Ez70A4NkRt8mgkGCgel+zROnfaztoNWUL6Pze+hkFqur3DR1uuWa3
qspcFxDZrU+9LYAckQLEZOYc01XpUocjqk/mCbELjZrRmVn58TikYriaRBvWuJQgtOYCxUacddl2
liZPctNTTKF36RVX1hulYoUSV769iT4sJfw62bORxmbpc3jekKkDOCaIkMCkHLCLaEMcqrYq4998
Rdl97kh7k9Wf6RGfQftYFVx+CF3yHF10IZ4mhuXsJD7d0Jk4eCxv0GpE9er/wl4+mhgfZ7lUFzKL
AjAYJ8Mp8mG7qkNg1DSjMAea1j+Ah/C3IudM4K7WG2WLQBMSqmHLVQdOYWW/pKcFxEjJwhRl8I8e
lp61G5vFtW02i1/2SsDcFLgRvKDVkVLeHJzUKQEzyXr6x9uhXUdpEkkx9rH2LL1uvl0MFymbXd1R
CgTDTOjXCqMaH/+TwsYtT883REFEfWHaHqAfIUOgZ7z+9LkjZ4WgetfZ6D5lRWsY/MsLL+Lne9uk
y17BXvba0gvYiIdbrQ/jzHFX6ydzRTsfuUPVwq1Su0VytD+oHc6RuEBHBV5AjK0OkE9/CNfnunVg
Dt0Wii3yYCtpotdW62ZF8enM2jtcy+VLtRjvtV1ye3uwoWvXXdgSG0lN40mmV3vIsIGsL12zsd9y
+SINzIN4A0MnIq63/4h3oInPYNEMxlggfn3/RNPSQnLUHhm7IeOig+wucH4Ke/1bO1Y1lms7usOL
by72QX9QfmCanPQJiBi/m/iyAaY3JUkcB5YL/r+zl2NG+AbZP/0cha99ipzJQHlVTA79MFoI+Tjc
3FNrnmpb4XHX1hBZYFuqjbx1laLYsg5KSjcF3XIuYC604tX2WlnX+42Y4OaI9+i9bAO0XmW+TEd4
zx45KGjsA8G+OQ8zOUTynlbfSBUQ6JoaCA7rLdXuRwpMYD0l78BpP65w0khc5HKy8Bt/Lts2rEAh
yl7J53mOua5f+tshk7cvgrnuAvTQuB3v7ve9MrHJzBYMA2WVW0gC7kS/rl/3h7ADBA93n5P5jfzN
s+KcEbTlhc02OHdOubL4w2IF//G0TTSSCPPAct2ufBvWm9ntsN4ipW1iTs6OEm68Qy0ATjGbxAfz
gAnzAL3mF1hwzC5gwZjdj9Dsq9h9HPYP+7V/AVow4ap/HWqGJfttULFN7ei4aCl36TB9h9ZpCzNw
meyo1Zjol4EWYJ1cZW1M830X2nfVUraKFo9oMIlbCB78BpSwwzqiEXWeKXNqAuZ+5GTZyNy52qK7
cTlDRO0jrYLJrJwcROCpbcAZoSx+DFAzoJThZHZKikUqdetOE1iseCklzkQoJp/Yr+9wbuiw6Uxc
tpMuGsgUum3dxT8jo0wZBuNs6WHah4MPVk+5WD8wg7MWafp4wAEyTL5/MtnnamiQsGJtE2keQLA5
1rMYB45VhRLKrhmtOhJd5F9M10ceR09t6r0I0Mza140S5pdsupXxJS85Xh+Pru/GpSPdRbYPU3RI
ZtxEKmH0Ht3hEJxg7vYhjQgZ8AwULhUVPEoH3ZpdnZrPvdqyC2cYWrBQEDYBFNZEAx/NDqBSOZL4
zDylSsiFXwkjaqlASP6crzT7n9DzNGDhOcGUmZ6d1wgvlYO9tvQXeviTfFlh7iZt0XOGTxffWnb1
iFzMlWZGjXxKp7i7kkftBJmgQQ6APdWDhg1lbisLJxNW1bR3xSZp+cq3M/T5A+tlneihN1rRJKiB
4QIeKw5rz9hAp4ZF0oXQs7RRogCYOJDQWTF/7shkTsiVLQPFCxDeYxU1yySg8UJH2x6t4hbg1L1i
i/a0HgBeIacmXh9O0N69hLQ6UzksvJ9uCJ3KlPOL4QtdZ/g6YGme8+PZNTYqBqt1acYEAwr40qBj
2cqcykCOPHaYSV1z5SWQ4zFgCIV+4wJlkUwuGdh//NJ3378HgOTwZqNVzvKNPOC4UoawmCewRzr9
KAria1aImdsA/NPoT6Y7Sl9imS98l0t69CPlnPYizGZSIcFL1MB/E+rRlTkxPc7kwnik0hInkrRr
YIKZA77TIGMxe7u49Qi9nWVHvKM1XX+vKymYSCWqQfUl59EFWdW4DwUsM5TLT6cyVk8gWLkUfONe
h0wqE9ZH0UfDI2Mn7xZzi9cde3UP16//kQHBU3wrXd177CZaGeba9rxVonPGhsAX8A53EqRykI18
8Klt8kY6gcham0wsbSfqyCqUXUDbAdDebLKbKQH58bHoF4BEWPvSEfB2mf1hFWvnGl1kUdZPPaX/
1kzD9L7HCaYLUfo50cXvy3LPxKRHewIBlEsxNZZnj9ELESrsVXNJxFhh6x1/aRJkm3iPuQdKmswE
3Sa8KXGdNJBftwskKRtujGibWuonc3lhlhokZzOJCAm7PKU2gOPOiTmlEQys5OwiuK7aXELfeXTI
xINl34jea7M6mjRbiRvRb1yQTvu+EuIUYZuz10gnlA+Rc/DAcB4TuQuT3YIofQ8J6TNKD2pOtGlV
0HsTqRO09iUfyqdh4jm6+XK+npmypl22xmr4IBhSy94nSMFsAcLhGU0yCM/luhGeQKcaI5DXQ7Xo
zztoXL62ZMTovD5U2mKOLE5lPOHafubvNVReNORzpgpks2EjrcWLaCpwC7i1Za+IuB/i6ctoG8aa
B0HJk9TgAJvnPuAF2xbLKgcsGf0sxZ7urvfM4XXREOPh95SZ00ebMnla4ormHZN9vzosscT69/00
JiiBEVrhecz+p1vmlCIxmHucVhhmpQtA8x8rbVcQstdc3p1zDfwgGG8AhIRyemA0wYtP3a1oOyjk
lhaxfr01O/zsCqjwPlPVMq3CWsCwrlIqtafvVnM9hxLTccvNnvPuMeZJy7SBNuO2w2pC5YJpNJYd
fYss81vkcZzEy3cmzzRAoBnwdJ6nc99XjFQFFaTRL1593L8ZbvnOJ5Ko1AIQ+POLhFxo/pzTS+w9
KhpVla7bVxRxkp6v6BPFKGR0AK/tCfeIHL4H9ou/smCdG9uLn2o/zG3Dkp/gU9DTBPY/UePk5Zax
iAATmA3AlH6oMteFimxxaC76s8lmIdu7nPupVV5IjBZnDWbaj1xRN3PUd/zcLTo//8j6LfMVexKq
AUndTmT9GP+Y8EwNcljHsey7uQM9j1dRu24FkQgXUPuB210pp7ZM0wKsQ7oJF+F/rHNWQ8FkrNnx
LDY8RUF/7nQSQtktcpDlM+W5pvun24X0hnNCPONUFpQB2q3GgntTnDRE7T1z2Zu0LfhJoQCYQlJy
U+bwEIiuGcJ8X0FglF0EAbGUXlH/AngmAR/TT5Zp5V4MifddNrBui7FPlYfAHYrpYSlzEdYwujFj
vAHS46otXLcbcBph4CFcDKGh6LzdUtZ31n26J4kNjKhVfAscn5tcnBC7KdslnQ4w9mMZ7Z+spwsZ
SWfMmdXcd6V+oQvDw8mLFJZ15vBapPdxeZNz+xpnmp+aPIwweD5qHz9Vg8ahdRYWl6ARJrg1C0c9
cplg6xRLZoVbCmM0+4zTLder8+ZAKdi2wgDI6zvJ1h/SZ/m3JZhH+wlCZIcSE8qKdvZaAgrSkSMI
qA+rhBJBVaRmpUDTlnsZexvC/SqTr0T1jpAUJuWj/XfyLkCLeAnzega7LPFZO+af79Bl13n71m6d
hbSVMgfscNZ9QPOTYXxK28A+IAmcuZOW21t12xBN8MV0jV6NEtKsZWV82eDeYFFPLvb8PFYVsprW
xuQq7f7wI4fbpp1/yRMD4unnbQBKloSgfcc6N46bGFtVdyXUVC16Sp+1I/PsGrOivQ0ik9F+fcsv
zNMEaCDCHYMtAsttxyrfIv528gHuXIsQh/21HU4/hIYSQ2Bt2Y39Kn4iff/HDOmbF9L+ZJZ3LzXw
1Lbdmaoyv2Vf13UdRY2Dqa6FpTsPnbsIMD4I9OT9ScgSCyhj9cKBh+3QhpUTOBpc7mSUhlh44UFg
ukGkvycU17Doz7ga5UhEIaYSZTZXXvWYy722iMEksLMljSpHCTqIKjtilNy+GlhH0Rnw5NiT0bCX
thOAG6oba1Riorpgc6qrwKoSNfiTWKYIvLJlNJsWHFjuhEI5mW441WMFnPwRs1xELNykdNp3B519
6BUbmsjoQc2hZ/+fXhrUCJ6aziFOB9q1b4YHCTa3ZrkfFkMRx8ixE80a5wca98+d4sxKFCMhObuE
1Qv6mwVacyGsn/PbYfei49jbjErW64gMfapUIUS/YKhKY7pwTSoTJ0sje80PtB4Pk4Os2VEbZkUC
ADr1JMNUg+sHjVM5pWG/VT/kIYxVq9ShiiHyUtb5CkQKruawptulF5ft4LJVqFOR1KeG/Jp1WCJ+
Ay1s7oo3Fay0GsnUYvIHsDzSRaHPT89AGpiyzh9dz87+EbfMolNcvhjleWZ4AEZQdvR+BCGo/8MB
N1cckTaE3SJc8ZnhQ8GLax+CiO++0i+Us7pYCkGIGQ1/TQ+ChzcqzKKRWcgnYqw90y4blXAKgbAC
hk6Qx37PDzIKspPtuyA3ssYOKouGKWRh6sYBA1bTOczcTiwdSnwb9Ru+k8sG6uQUHClUu//cBf+2
zZ2uXjclRjpczFF7Ill4DDukGphX/DtiJa6n6wOnOA/u5CtKboBcO96nKiIQgacVE6ZZbBtknoRh
cbjxUCCaT7eA9yLimSSdugKCUuDGDDkIOqXYd8oUKXvviRnlrHqnwTyYHpyc9D3QCGafYvXk8OrL
O/w/SZK9glw7i5Vefa1LnOdsYBy2l5NhF1AgoYKwrKPMkzUPvO37dnqb6r3rW2ZLjfcYTODmWiwf
hPskhJEHU1IxioddSwzr4pEbRmGefH2bJR77XXMO4TSiisJrn5jgs3caAOg575SxvjTjbSQTT5sd
PfPy/mWIr8ayFvhHNtK1TYTAKDdoIzgr+56gHRcoaSjzVW149XJV2OlsOEFgpO5Aem4Y/UeE7++0
0BgBD5mbH6IVMCv8AOkUtaaGWhWU2S0N96rd+mJnPmKNs0FgeGy/Q7kL3FRQJh4m1oEp831cbqlN
sd2VHVMMkGnS18f6BHT1wLmRZj+/g4ki5Ao1cAENVlJji7rDGRCh5Rln49mQuzA97+SeUFihAVzU
N2RBqQ2V7XFDw0NkgzjFEEYZFwhBJCbpSOE76YJOagVMCsLAhT91T6mIjeU5lKpnZtxBDyoZV2LI
mAp9m9M8XfkbaSaN9o+ieghdaQ9xRAZVoesewRiKgOw/2O7zsgWs2XCxdEmtnzQfQhk774jiK/Ly
7Cl+00fLWm79iZJqo2RTD1j39tOvIb35x2sLl3PpUb2czj7ldQa7C7xtfVpOzrisJBrRz7zq0SYx
YMz3gXgdgVh+7OZNeua3VrHVZqQ3yX5yn1SaxZU3kMl75ScZEZTqnNkz2ZjTRRGXNBVzEsoCWOCP
teHhF804+OcXE4f+/WshZmN4ul0fxoK9IhnxZZCHfU45EpqV8gAYcwLXTE22NN1J2oVzg9hkwh6f
z34ljtfmPCDFx2Ptxbbnw5PGMsfY2s0JBTvaZ01fuYx8rXpI47FkQT6H0c01qWtZYiuc4NaAc2AC
5YTugVe0uuK4ht3WdPMId+2wJxC4nri9TP7+Qp3cse1DPcUMa5ppAjWlp5q37uUBr/NMyRLHnvwA
7w6osy0ovXVTp/cg5ksCNPeiNiGK9LtPKMazXJN1PJMqTtip5JTVj5TpDaaVJIHVmCJV+3MjH2Z9
5S3dj2I4Pd+Q/lYaArJH/g6nkPFHiKA0vOI/it+6p6mMLjq9ri3JAuh0fRLxtWKbxYbsetQLJ+8N
gwp7Nv/q1K5DgyFzFMtfgTej/mS2lsAQU8a969YShKAt2gD+9Ctd0BxMyzOV4VRA28yJVrbNBidT
9wDLzMA0NdF0c2fCp0qa0pitLdicfBbumyAIUcG+oHoW8G5nLoHHi2ZaesL8Y8hwpdIibnuxWfU6
tgdXRTwGGXMb5tuMIWLXCRpdvqT2/qEY3WeOY4JcFlprWVeK1VvEk+dyqyUHWd63f0/WNrrTqhxe
Lmy2Bu/k77Qd9CQb0Akq+Cu51uc87tGEzOhNpmTDCUXIBswRJjl5EtIcBPXHvOSQbRWw/WEDo1uD
NlfK8uAAd3nQryfUDaQ8PU0HKZljhAmzGd2Rel05Fljy733tUmrYnumOo7oZYLXBhwUSQZq0cfQH
FNr9cAsw3shtSBcfz4L7tf6c7AVPQ7pFxQCAJ7kb/SZPpGk0wREJwmMMz4R198hgcAILxOMRzyqN
ckZIG8dJU2bM3HUxm2BpV1sNkvT6SHEXLA6pxs+aChRyIv9hOrMKNE28xaqQUTuA+Ewd+RX6Gswc
rmYcdS7eJb1tOJAsLrQZ0IY4h58bdqzLckLRxPneIWR9GqDLi51+8xkthfb4m61J06V6gZ8/wEzf
uupjprYjNQmMFAsX2cJioxo+UKdQyVYye6KfZO5Zp2xjjFdUxqnxQn46MNNX60jQrkKWfXaZcmPv
v83zxG6jJHfnIL+z4tJ/yAygFRJ7tjJEyuG8iKj5pWKTCBybdk2pbS65sbuuBU4PnA8VYaBuZiFl
ALoLFYkshZlLIgtT6OwciJmtFuVvjnQO2jZtBeKr595Bj7N8pL2rnzuI4Ivrp9GZ6u4JQzr6TeLH
7XLfxJmRJIpOZ/BK2ufs6GUTmpNirTpCmgAUix32pFY7I1p0fTp7LpNwlbxqPOhGQQH0N8LBiXiD
6CtVpnFeaSuyvFi0iwx5CDqACX0k7w4JRX118Dd7WWwRqBoIKsU454p82WWfPjjtw9thiIWJmKCD
oM7uvDs56y65rqnSDqzNxgbLItF85mlDU9wH8hYNN/Nt8iIKXvqD8AJ+oo66vXeiGEdSpQ178waF
Gmx14hKGIqq84ms2UojiRVp7949C/OQiC1cjsvcJTU/AN9HUxZUAlxCULQBN5GmIDEEc1i9e2Cix
nm+PkglXbJHUdfZpKqOVswRYP5cK+6BBAy7Fz//MhkFLSDAwMF79mde2Uf9IM8s3phJpagH+bzEo
jvWcJPiWCKfpj55Nl97ekBpq8oiC8prFcsv6XxqOQdv9oil4tbhz0Z56WJXK6b7HiWzDSoNmPXQ6
J3cbSf7xm/Pkw056QHqbUMSFCbTyZSMI6IVTKMRDWdccm0uzVTqD6BqNlQpfXkcLP+8XAK6Jtlhd
3PnDIbYxpMAdRbqfC0eymCNmCBvXscoM1XYWKZdgJEE7R42RK6nP3rBbh1CfnKx59CxaFdNFraTd
sBlIeX3fqlm3tNNB/Ob+pUjiKZwAs/HdjJJxPZ6iU/0enlXRMHTEUKHIMR+U+zah5W1UibY7BPJD
JbjWBV97zMyXCmJlzkOXTaZ7ohC/MsEpfFZSK9xSniWXU1NZ6kztLd3dbExmvzV/IQ9Hw+BMfaAs
Z0IiSBhkKMZ2/1dicmrBRpXTmDLo+jZxvxkvJ8lGAzXdPNoEbxwRWXM2UHFNoDaKF8iqGb8AsASl
EvCDGrDDieqnDhDtpFC8E2ksfUjM9F+mkkY3NC26LzALx7cqNhVjM5a24dl/JJyL6kZWoDsX7oy6
CrcKSdlHqaSWWhiQBQQ9P84SurQMXN0dSrZ+b//oJ8I1CNrfSMREpig9HYpCJOUZpNicqSM6imPI
1/g6lkVKTx5RlWGi/cFis4L56aIQFb5zhHN9RNwZLZiNJ4XRJxxvGScQnWqZ0GhH1FIJ7X5qiUVB
DwNg66i7lNMh3MCaYWj6ela4v+TFVYgZvSp+V81dW8lZVDZBQkQ4UEt6BsufaqWiR/8Ziq4+KAXO
zwSnRaXJJO4lL7/yJrkPqkpWojpUFw4sJtN1rhQzSHEPmWl5yVqGSwYlZ8POwCeDTytp9QtzLlrW
93Gz/tbv5AkOaW9vaUylVb/wj1typOznBiCjnO3/AnDMfyhh5mfqw3HcglkCSc5y5tKe57ef59IR
8pUSfRhvIs3lVs3RWT7KUGx7DB6IsflsUSnf/b5y/lPrHZozOme5JCJPfdWaGp6PxEKiMsEm0r5T
sasRQk1rDTSclcLP0q22XLrYf7jbeldEr67/JbgWefhBbBewE/7U2sukTDft6l9jOYs7nLHwODtC
i1Mc9BtwXLAxEFDrpnzjYiOeyGDqhfOZAplACn/BsRSR3y/1GKzJeaqKta/DQc4tC+uu3tFc2nd2
NoluuYl/QfFHORKYaV5Jn/EbCOHRG+hwI8MYp/q1B8JQbt5sxIQA1YSftNsviZKN8d/AJGGlkfLp
Ky0UVDkVe4ePrPs8CwyfTHldGZq/u+tWHAhKHJsNwCZztXkoG4IaTV0NmWfui74M+17eL6jYc9tZ
UQztvYd12hNhN2nNm+YyipuhSLO1h9nq+5xrH4n2W/zdHjdnSxbOQPXlz1mR4Ai5md95Rjf71t6x
uiOXyliqtKL36ljSpjedqB1E+4O1n6bFWhEFLMsE7OloTKMwcIgQBUe2OBgINYW0Z4Zb537G36sc
S9ATthYr65DGAIk2OV5m/BbHJPJNwEwcE9feOURStV3NFkZRWH2iEBBq/3D87gGxhRoB68CARioI
NWVLmezD7FLatEVSR3q3G3wCbKlMMPwbX200OyhJYCV7I6WxbgZqhBrPyUhbSMk+Y0dTdd3gQDb0
xgXuo3sUa4ZTTFSIX5W7Xz9mc7LEVI1X8N4hYTpzdkZFauD5csz6HDMQ+x+hbiE4iLcJVTMw/1LC
F8FuPiJKjukMdgd1lRcv9AgGkIpNsY4bk4u0iRRy+f+9nWY+wW3/45XGM5X48Z7iF88wOKA/aVnz
o/u+NaacbcAFNDD/gxb11alB7m27YXr4ocdhf1DsAGjkHv+09OBwfkmJv8lfRuxdAzXOFCP2fgs7
F+YqVOcxyp0ecuMioOFyXQdt2EZzCeeMm0V5bvbc4A5BxbppTv9ZymbQl1JDVGbiVLmKzYGssIMl
otCGf5WkywJo05GSZUJZxA/m6rgNolTvckb/Lgo05jdiTCxWUN3xLaRZKgDDgGj1tPc7orjaslbR
/dwTA0iy1SN4zGw3CL7FRHG5n4IvOioLa/wHp0JEqomNyLuDo+knAuRbS1Zebt+1iyTHmxSW8VHQ
Jd7J68N9OcP3at1La1sGc5ErTI9BGyA1XtHalfiPS7j/1VCd5XTj9y4wrqINQMPNpaZxjdkSAFmt
kL7P19iC5cOkP2DNh3nIo+p/R1WHZm4UP9+zKzdhSdV5JA34Nsqpr+6igoy/pKS2N8rTw+CCmn3G
HR6w1hC/Tl/qKCDduZi2uXwPLXgWeLljeex4NI9ldXDLoj9PVrie6wtcYQVd1mHOC090hyNvkmdF
6piscgGDmYl1zzeuFqHapH+s8tVdKf8pK0OhEayqahxB0lmiWZqUF3QZeIbQ2VC3p98krrNgRtix
fy8u4SjUx9720UHl4+sN2aZMJv9Q+XEfWcvNbrHxpvNcI4IBWz2ZGjrB4Oysx1waEBsAZQawTQMq
XTn3zRoWkiOCCCsRS6AontTf4aPHZs1jk3KpeFiqYIEEoh29xeYgpjoRdFdDcJJEDzxjpwGDnsoR
cFaL5++vaB1Rz/r3bc3g2qQckVyVu89H4D4MtNGTurWjjzw7zk8NYrmarQxt/qFIeu1zdqu4L+ui
DIZx9bLgl2VwfQWY5OIOm2APvw9IMmTPBK6nfu/ar18KBJLwHTDFxn6Pv7DkHqIoiRqs2B+WBkQT
kX/AU1caNOeNbQ/lDUBd/I8rsxR+fUDfLNJhTQ9xmhMqln+FXkHlSOZqNpiEflnpWtFyp+Nc0nrg
UE3weAgZ0awBV7T4hfHExbXE42W99WlZdlbv5RQ0QdgQKIxn8Ua0NzUevaH1YkvKlx5C61g9UwuF
RKxBWr75pUCwxelg5U0cWddXetWc3o6pGLTPmSvMrrVJgbnpfKQpef6CdcZcP2Yg1GHHim/7rrhw
dDTcAP+YtVHnBxMbiwIaTHdKJNjgVxVfcqmk8yLBK0EIsSvZNgCXnrDAE5uZBWzJIx/iNIgeKan9
uZZ9LgAYCAsiNX+d6tQp2FmItK/Hg/midlzLqr8+P13Io8Y5RkAXpUTnHP0UM6zMqI1QzM6E7IXK
OwqH/rm7b5+lR72cdlyeUHlbWOcN4VFR0+tJlAQ8QsWwyv4sN3C4amShFBjfM/FdIETJPhfCJifr
Mnju672wZB2FZa4n0sOfkdEj4r5AT1qGnWjnwhkzc5ewHYqih9/suTgBXKFrVSwLYd9SZyoG+O8a
QLi/CmqJR8S7hAQ7zMqqWm1O77UQRqC19e31mLEuQli2XwaUAGWpreOcsJPkOsk2mJcqSRYoL3nZ
NT/gpzTy+692sPVGVrCG4m14vG0awR2+YI9n6+hU9ZS6BkfdYBk0KqgtWpaFDpt+qCxXOqziQh+l
ktOdnHp8IEl0jv3iyNYuuD3+2n+UDTAPZiQW6fRN8uPFbBsYSK6jKv7Wrw+ttGK8p3deU3+NIdbu
/4/sVPLbN7JAMqj3xFopYF6rrfTsDnEzySAILBjcXjT47wdtV9NEL3PuOjlVLIWh7H3gmIfSP4Nq
2kct/NDpECNReI3wXWFjYf5PftZT1oTSAoQMwjZujyKHSiuZVpgUBjSxowQTql1OyckesOWBn+Hq
anwzJ9C2ooXXqvOQ7+Lx4I5Ud81RGAYGPSFtkFyAV47FHDB8wigx5HKnWtJ3+KePEVHfC9oIwavG
IWOH7mY9ne8a/Byvh+YSqjRf+h6OJIaMNOIM3kbeW4/GiZcYkR98YHk8BfWrCWDbnXfjYe18j9YU
Ynn51Yih8C7atOJhCsBYpiindYtqcN75Sd47jR5bEwkThezSGTTTNSiGSLD0c3sPcrOUi/Q6YJ46
IILFpZDET7pF6W5oLHZJib2/iMhY1V/spfkkIN8RBZUvsdHmG+48YauDWv0Z6G3CBVUDK8+0D06m
GXoVvjB/gfNNcyN9gy8udEecYLi86O1TKVcLSW/coIE400GOEn94lAfxHwSHvAU7losWGShw3h+l
OHLjQ4GzHOdb53Pvix7N6++ZgQAc6nyV1Kal0sFMKijEmykmtla85KDT7hCztMEbyoz11q/jts/8
Ph9JReI4IjCXBDMkpTORar+2QAMsQjQjMpt2bjgM8ACgAiedhd+MUGcEl7f6fS4ZJJ/wG+YCugVJ
g6WBXVmjA+oD9cjJ8dZFtxG5vKxWfPOhf8fVG7K6ENpXbs+UB7ZLYkA4Ip/F10za4DvBbOUVhdvW
zCEYy8MqqFqRXekKnFe6QMSHLok6JQwiIJCU90L3t9RfSPxFDO1a0I5zUrmfnuN2Im8gq16WmMRx
49XWeGHiVALD+YPCUlR8fOkspkg48oEh7BCbMLQaSW3iPU16EMGERVXczzi2dm0J9ui4WIgcqG01
wMyTstIdpJsW/sOVNZdqQBkjBI6ORcbBkr/1ffysfl3Zb+XH+NywWbFzRejD72WUwvP0UljrOHQI
sHIEnKnobTKmvRHIR8jr/tJnk597SJOTgc6WmL5ZyNCZW3MHqLT/0AkyNCCBdW4JyeIoMjMM+4AO
RX+orQdGM5dH7K11H9VmTExQsJBqhFbwju5RrldRRiqjFO0JAHBwbSXpPEDkIzWHK9czkQILi/H7
nr2iHJ7aAi9hZB39PH6ScCX+AM12hjijHsZVTseCiHLZVYpqYIxNTaOdgKI6T9Dg1a0QCuNCmw96
D0ei/PKsuyj55No5jU8dTtS+76X3MmWEOH3eOc5la+yMD24EACfZ104kW6JLrKQ30d8pV2eBF2O/
wci7/KHewoiqruPHjJIh5OOqGzDQxp5wJflJd2AwAiHFiU9Uvd3phyDebERVlvWKx4f6GcE219Qr
AaLNtsrl2UcVW/dyLJcQDe/wB8JJ0rlVhIHOjb3njXrqDmQ+EHww97ScAYnl8ut54T7mBG/hTYcE
Bt3cfmw7vavSmGvR10K5r8lpCzjYvaKEnvaxfnHw6XbgsJJRmHs0EWzM/Qdd5nssDmcdJC0A4+os
Q+gqFi1BQ9ACgb1q9Tghfdua6vMcVfFGOwf4xdYeWPG+quTd4A3z5KGEoQYcVwNaOUye15vql2/y
BMtwXyrsiJ257xG//jlGvSVYWX64uFuNXO/LtYzft394d9yfZcEJOL1hflmKYmrHucYujkGDhWGm
xHyj1Cw0rIYyPxdtdZuWEkk4g15YgJJ6h1iDOji497X3ftpzSC1O3ejUeCtLInadQed3eFguwG+W
9ucw5RxaALTtLSWBaN8vHftshxpz6jdvU6y/0RZprOfWOZK55L8ePq7RGeT39lfs7kD8kFbIhWPl
Ja9US5Q2sDNm1Y7RnMvTMLsk1JjnMqJlRhG6bjl15I7enEdlt59imYbpxDuNzXXoUBvOwyhxVbnX
Xox1O7mVrGYdWx9sg6WEkJ7YvF0wUE6LIL78nNQQOB8yN53Ww6i+u+zC1qBJJtpRolXNW6rUQLiz
Rcb0no+WSClFLGhYBzU8CK5Wn25Wk+zDPhnwuLPWMummwq5UMruFH1L+O+dmb6Z+0zbmS+xe5ud/
nZ6jFtLdv7qCEpdp0bL/ZjdGDYpi+ogJSYt7JcyxnZwp8Oz1cihxzUexOS+vBWXvc+0N/r/K9Zs1
PyWaMnsHB5nJIRD22wSnUarlppzsjnAKApyEw2WX1wOarmzJcSULuy7s22ybYi4JOGDtVjDAgQMa
kOhLMARqDgShjUJYyy7WMUHj2KyQo4Vka/mOm4ACgd/vOjRX2xSp2pwckR213rNJV30woGHY570o
TqejgzA1zkkXkSHH9ASMSZ7bX9EJ+6oSxG1m9/jRTXb7qJ9pg0YSvrAxKEr6KMw/5Tr+aqbPG8uq
NFUAh7tOrHL5/ElswRLsTd69gLgnCFDwvywGEhgQ8QV3+86i8dUr6dcoLbqxbHFgfnrO7nSSN6rK
bnqd57ph10j9Y5wBh6XSGoGiPvjoKG7KA/5bag4g+EOKWmtzGt/C5BQyb6qFQZRvHDzQ3ISkpKzv
WAaugntltNpxAyFV56474opKcIEu0fpp09u0ZTM9CYCM8COMZGrwutXAyzSzQ0rjsIC5MMasqDN+
P8sVxP5DdgHq4Zpw9IwSCNBo+gq0q82yyZMHTDsgzBiD6c/fucxXrQ4Ln5wtVyT42uCoHITjhjsf
9rDc4jCs8VB7nnVGFhCQJV61mbutUQQOGKnd7G07OAfv6Te+xJ7kJOWF8Rfb/t5zRiIfN3W+g5my
C7eAqG/17MhggPyAjeyIvJnZvYorAbU0Net7Ne1U4zS4zVI4Frovx5OvVgyiCp0XHFmDsBj4tyg8
uqVmh/67THBcUR/HXHGvxMmjWeUfh9wygOHSUWkCLHoDV7UoCz8x/lZCVMxnbbXtIxvL03c1W05e
i66EDe4VEpRLQbI80ezHm4xNM/JdU+8pYbo4nlDnF6K1PbXSAlGmvdWNdbm+pEf8qlKJKYurfcCU
QtTXQZPKTNCHIK8h6xQ1j6Z5QvZvl+eXCeBM000OM1F8/g6LrxFgTBAF75emGi+K57In6vtfWVeO
72/Pvgvu6XmVCd+CtHUbYA1mrTsK0VMXbuwVH4cayPGZXaJwFjoYqViPHWI2zTeM4Eq3lboL2RKo
azl/htsQrZCXpgNmMxp75cV12zZPigIWb7tOJYVQQh2o/lmCMRom17LsNXDBLePdB6ao7IuZrXeW
+Euog1kbgXOW5MVKOH4d7HKWE6SyY/UAAcGIVgnfAZu8bFTUgK4XaYPPS48f5GV4ndFkK8hZRmOe
Gw1PHsj4LqVVbTXDZmRrfYmbLpCSbQdYfV3Y8BJ2dUP6FPSbBtUoGABazZ7WM6/kfH0jCyvBrvik
s8SiK+utkctclq31VKRKArHZij1hiF4r4ExnmZeXO57heP1kik0hZcEwWBQ0uo9adDKK9gPny/Js
KwnQLTaRArDgOSX7xeeKtYm16E0uJRU99oCijsasTIhgelCU3wAXCEw8yoVxMN6RVaLtnNDfyIkg
+uw5JESzzWBvApBbjWMSstdMZiZ2KVROwlt9AxqdpCeigVqIurZ7U/6hhg7stlr8E5RLNVpyDttc
eXpkRnLLd5bggrniZkdQFqDTkwYRf5ZF1tIgmA/o9sRRLb32ZVdcGqa49JGNlFGUmRS85/bSbJCB
XbUhSLiJNDAot1V0UIglL028AhtGRgcZpK1msWNB/SJORiRuGPleZAwisi6H8BhFlBcKuVZbU+CK
0Fw0LgIP5QEPrObUJrpiQsZA7TS6C7S+U9O6s9ScLCrJ127qzXFmYNYJWhbHDc73QenSRFZVp5Ed
RJ6QClR76xV2E2AlhGC+FOZYFMtEIZ67s43h/GCO1Xs9O+UwTblM3s50HH0uhJPNnPqcioUd7J56
z5sJS9LEUT5/EPlIvZ0kbGmggvQdRFrx88wLrkjqpupiOybnwOGZxaGDGx6uNKT2fzlZhLaj+/nW
CFnZ2c7F7SVpxuzAWQmBHs6zEt+Zl83TGU5AIvwZeP/F6brnqyylC5zuDrGWrdHzAO7/xOEYF2it
JxbgBrMzYVP6uMZDhK/vxe2D8BrsV2waLh02oz4ubq0n8YMBHVmq04eGnGdV+oR7Z3BnLXVzU0nW
ztpH1ba6yb0dMZ5yRe/LPEgO03vcczq7zTU2pKcszK73cMFnLjrxC/06cdP2EOUbqVeuS9P4ZiHP
RUP+24Xcob+v+66iazyECbWBlzgsUschOiA5YFz+ItyKT8ADfbx6ai12P1xlKucQMaxP8e968stA
knrWY9beRuppSnhUPiZYfw5MVSjiM0EhO/HB2zh1XAeSVZNH0tgIsdPBR0qlm6CSDVQm+B9t26j1
kQTDgNBPOL4uvOm6w64w9ErDxz6oGhb2Dp9b37edQuw9OFOmGVgi43jubwUW4bLXhFaH/zvrjcJ4
CTyomrl7kvxOkaaWlrTu1aV4NEJEEaDAxk34EuHdQ6+aC3WbtnGQHpaulXghrdFJPgAUIQonsKpv
pkY8qPTCztJKzm3X8BMEjGqSrad8KZchRHTLyq88WNqRHoosb+rqN+sOnFqkkvBUAr9q40J2O/lI
W2o7DAljgJQ4sPgmLCzJN3WaBYvNQjtJkMDi3qhauOYO5CoRmita4I41KPd6asRyVccL6yBQ0hOT
D9k2EzpQu3pF73s6L04GY86dCmBqSOwTC14DlSXnksxZJNNmDEn1aCUsW+NceBtFEoTcRPZ1sFyB
ZdfxSa1GdiyOOiENHEFTp6/Jd5+LXfeAAsXEB1fQs887B+SbUDdvHfyV2LWJnAryO7ZpJNPHN769
mlqj/4Q3fQfDQE+T4vw7bjOlDOmAGmRCZqv/+Ecs2NokPx8c/oj9VK2UPjRSPyegU8kUxbfR2KW5
noTDTa4w3UtlkfhD8KSSgnjG+CFm0BVkDTvLcRe8yBgricH0Ajrtl+HOnoPvYfzoYpbVFrN3aNyu
yImL0Dc0cqy2PC8SkvR0C0z6WvqKXYBYC+NW64NKZOVuz/vDzdsJ4NAWth7RLu2dCKXxJIVIRppa
qGTWC0cBJgqoLmfcBlO7j96FoyHtKu9RrGp3NRKfOTvnzqe2JXP3qXGIhYh4cF9mAMZLNcw+A+09
OS4/TLsu9nOjjmd0fz7vDH79+YP0a1/5mHhr0nDtkKZPnHT/aDkfnSREUOiY2JuH+1Kqs4SDf1J2
IpFdJKadT34z1wnm1EaNtyVu0cilJI6Z5cZ0/VA4/x6co/MxlNhaoI7G9sYomXu6OY1V62fQqGnz
07M2FUDPbR3lCjmiyEF8BF/YpX5dtQe7662ilhbH4cQ2n/GytKR9cMgPYLtyfroRriEtx/mcH4Jb
nL2wNK+RaY/kEsBCG1FRhw7s4SODzAF2ueplA4DlM/l3jA8l61RPxMIsZEE/atw+jMs8gVDehQ7P
inSrTtRseL28QEiCilJdY0tZ3VJfLx9v0tLlP3Uem1Nw+S4hZhL7OAqSYSpUA+eweLclI4e3CG76
DanOeE4EpIuoGmpX6lBa+APMYtUIw8HhtYN6Wl1U1ozDirflRAGAwYZjT/zjXzLKLN+kSUeUB6V5
1DvAB7X8MsCSu8Y4k+DkLtHBLHO96kLptlaR1bvn+ADmwMd6WjwV/N4eVV2IQ3GuyOn6lgN4YtfB
j3eJ5kZZseewGNPGSYtCBVZQzzCY1IVbYV8GBL96BDkc2vuQiDy2ThrPLw73NX/ynG58Q8Za53bJ
yEupOY0FRX65eVeR79BtsYwOaFgqx/XLN1gMGhVkPvrfhLVA7F7CJL7Sw4+TKXwK83vQ+BDUL6JV
br/HuxzHYCrzY6W5aNDlzRNioao5Xn0pTNPIyO9MZsryoI1aIxWKnAZJGX5JpmHS36R7yMwS41uE
vZ67HTQ0i8IjvLNmagFxowYicDSlm15MM8KVIieaqMEO8DF5+yH7h5zh9NI4CP4TH4DAe/CHfCjL
SanM8/fJ12iSb86j9faqR41UHyoS7VnG13HDOQ/4TVmmtVHZnwB43JYfFg3llpvrQkXbS5XZkS6b
KxoAX3A67OToEJpqXyJ6Zir/E7Ii5bwyGLrVZIcfG6R0CzpcOZdR8D6cN0lvBJIujLwTrRNCiUNf
6hXlrW5Kr1NB49cI5Yc4iCzYrL90mQ99l8hNQWw1f3OJ2KHcr7Qw0POJrO6F3u42bMNkNBlOuya6
g8FoqMUQiYCUgbEbfVtv1QcXqokVrLQ5JVfXqzLd3g5Cq9+QiqPJs4I/LpdRoerrCSrAv5uffD8u
M/vRoJZ8ftBXesUkEAVf0vA9slqVgU5GbI0Z+yYfmfIRGzUksj1ym+EKDdcd+r747oLE3+Os9Gne
H3fpJXbY4skbMdAvLs5r448ZGNZ1LnfhE9dALeDyXFZh31xe9QkbgXBm5DZk7/3afKUxm4L6tmr5
d8HmoMH48B22TCkPf6Osx+Er1hdZtICB2/adh5JUiK1c08UvBEx5jRXXFw5bp0SrrfTUGSeE9fzg
UROLiYe8rDnBOEEmJDaYkNschmd03gKvgC+CJg7KMHc5kbT+xfP0Npjcp4/MfNvSr2i0tFXjN4f2
IllxhbAdvNkBB8wrzTH4WCq8zWP56PhzFOS5yyNe4JYPDVeY3gwQm5ogkm7Mi0v97BkRLgvt0kFp
BR66QbtaLTIhZA77yt0gaQY20Mi5lOfW8Ddp+nSAP8I8yufl9izCN5G3Cje0fenYa1v77rI/gafG
aWoR2gpR48FQbhuIPbUjUO8XSM0MiHTBsKf0zrP1MTclo5ipn5/jYRwr01pccGSP09Mr6sP7MazE
xWgJfB/v2W8YlCGh7ZlIXHJfR7OLwIOrGJlc1MW74mrukCCx8eB1OrhRyMfRVIauwMBeK4Bqvzwh
54nHZaXTlYfKidVdVVElQL591Re0lFRqqXMGW3vcsDVXKF/LBs1RYXRZacIdmCP9PQqG3NUab/a/
u8iisXzg8ND4yFwHOjOjkgy+HjQdDjWv5bKJA3nN3YwDK0envHEZOGpgozIBVzFO6Jj7Ye/VObZ3
tyXXZRDHseiJfrUGJa4Uuv/jh44kG7VUCtzMo0E+msPY/6IG7MlKSUsoeGOHP3ZL1dP2k17WuRkr
utb3OANcV1RkCBOTQBbZWnMQdTlSqaGxAtWzy9Atmya+bNzplWgCGjGDK1yGQvgPJwUofwrYAiNA
lorfQXLSkS9jGTNW+9lgdU619YqQgqOqp402w/xRXiTf3Hesk4RZ1SwtBQo/4YxD0fh/b13Bxzvx
VpXpTQ4RBQn77R1HxLBNvo6NE2tzaE6k/DfdRJrt9vcwmPezAz0dxqCWY4iHqOnvP28b3s8x1wDM
BQKc/NBwVZ53UzDgoAzRHYodZh8WEjxxFu91MUZbfLn/jZyR/sGsVLWSxTWy4AMwyfhdyk1Xux8w
mRBuhryjtG1+/sONTUn0ZDGJQcmbMaV/vH7OI5ANuAVCmEJdPlo8qgBJngrWSeyjykd/+DG07jZV
CZ29Hw7bYSQW3OitrilCg4s8LA6h2qCvMpwXDdLaCLAEz87B5hRJ1JytKDRTHgCJ22371EDjNblr
2WyvaswwYECgKEbvb4tfsuz+/WgmTQxNH5vQy8772ec7uLb98Q4dbeGlqVFPpiHevRQWTApAFz0Q
HHdUMI47W7FFH2J7sAoAgiwPcJavyW+w5u0eGCYYtxjbTz2vBNpkrZb3hwla+Fa6U4zHsPJZPxPJ
c46VxM3vyWGvNUyTCbDa7T8bJQAVMK00XpKvN+XOw8tEyyFH8NhNWWS4b/lmYuRI2QEr1nXXkUg8
OGArm/Xc5wRcAk9z8/JIG+TBZVYMcGWYGPCjnAMai0yiNbskbIqqOkt2/9YZ8T/K8R26b2wk6iAJ
OVgs4BL7B3HR30Lnc2tBe4zHH/n2ZPLupJJmSFvNmE6iAgbisTjSBh+Kudaxrs0WQWxHiP7pI5Lc
scOz5D+2ENJE5sL8UYneW99aaZGgmUOlME5nvNeJAhTefpHKeDrM4aB71+nk8s2+QrFGkJ/79aaE
g4Kt0M3ij+lAdq0YjjuNg76W25l1Eos75+rfrYl8MVVQWV0m9X0hKvpQYq051IK2p4rL72fizSQ/
Ue8yPjXL/XKo9M5Rvbrk+qZkmnpFMg/Sa+rNOgBqm2nsK+eDL/BE6ADibRXNjd4r3eBrXUhWH1Gj
YIbXZsJPu9LA65x8Zs3dk6HhF2ilo1rgJHDWr04+FUR+B2I3j8EnqsNEgV4qlMUpyZQYELwgjDx5
rjk8lV1inczbdjLzMH86swegA1xAXR/TJZftRSYBRM/fnUPgjYXVoxY3KjbcgzOGytKiBap6gzBW
sZcejbJTcpoQfi1Wuu9O1Qp4iZKaBA39N1PLPh96eLCcfgzEqMI66IfbnlnpEaMMk+hQ9UxATyL2
GOU6wx1xS8GwJ5gpH7LvvwGCSPlbm+gv1adg4AauUqLFP3PN/Q/dX5o/YeEEHMbuaX7iis7Az4CL
FkSXBBFgfMmwlhxzVwMqtML9Ld1MtVNRSl3N6jmGqP4lM3Bb/2nAxO7wqag8OJwFp/thQqL3U1nP
Fha6yeaI/p+htMEhGq8H1VAgCeOxkCzqMwf9qVXlXoq1hO4zY7Cgzqrh1Ykd0jeaGvvTO+93jecJ
ShmsQ1/5R086MhRkDNQaKMvuJBV/hEGbhQjbbhY8MqnhyMjroYyzo1d6++kPAvPMxO1QAcoQhwXG
siUgFjiByBvirhBXzGXE+gjX/ouq5KdwIaVn35jFQEArs1VxbeNl33+aKcCnELhwLFNKSP1NyWE2
0gKO/6U3wK0+VkHRVkBgrIrt81oxH3KcikMtwH6dZkNzM3TqMHWXLBh6NaMxj103XezdYD5dalt2
n6UUljYxPDwv7+0MI++9/4W9TyvbhMVNKQSrp8g8QjAUz/LhtQpq4LiWfBj7ehjdRJoEHxToCSYy
z0KRFUQoRdpkw/ZADAiWHmHSW2kZ7EiSA9RbmkRP4qHuArgECVs4TnIJy1p/VTOplTSRtrBsI2m7
aCct/E2Zg0MpuYTOqRny1lDsbhOuCfERT3PQA3y4unzxyxE3qtkGFp1Hc2GIjExMIVl7Hk6NiT6Z
spFiYkUfVXR8Jt580GQoV+04mlLUHt3GshSpE5P2G+YF1MokE+7rGB3HYkgKnJrMVct5L/HKL9iQ
h3igWb3vrpa5a1/c42mkLuyx/ge3Y6TVvQjsE7AUK5envNMDxIJH0/8HOic2NT46D/Rnog3wmcX2
xT8Z/Fdpoj5J4iaaQN9eAgLBDQeOIzO7lqm3Yi+yaBkPXJKwflfg6hqpqgmnuVVDZLAS46cNuCiD
gwptNpqbCkXCR8xeXoG58NwQHUBpZ8SdLwj/RR3jznBLiyPfkKO7MruVKnL2Ey0/sJiQ49I/XbJy
SX459Vl8F7sYwBbKJxmybN/29GTJ0Qh3qzVPON3NVzZ0vx4iFYBZZbVfwmIrLWMerewnFsPozidO
ni5Ch4LPpeXnQ/U7JALEBB0lQ+I1CZ5WYMq8WteTIbMp0Y3YAKsnzR3cE1pTlwOe/tIg3bqFBK54
ELrnYYw0dRWcebbdweloRVY3lexXpJ+0UJPVDtb5FlgN8lp5xNDcAt63Y9LEv8JvWmAAu+t30ncU
mpUbPzND7i71y60bqolCtNHPhh2lqzI4StBKYT5yBiSuB/77UByRN4SXJEU/k1TPqIW11hCENGq5
IXf3ghpEw7C6Y91CHUtqV1LdDQsKo6y7puv7TIeK18zVBFr7Jc5RqpD1AA4Jp4sGV/MTEyDA/C9X
XOoBYkw5n0t8+kprwhz6IENo8AOsqHcXaOqzww3LFB/SkhxTvxdxHmbn5xPRlEV6sSyXwxCyj+nw
aKWOIpTt2ZtZf2TCjBaJF6KwEOzBbaU8GTqXhf2h9jK39+gRLtlnESNAKmaHLijvl7Y9nzbMkNul
Xb8N6eJvoz0SUrt1HtzRIcTDcoRmmb85UKyoHw+McNNO5SJLutoqH3qZnaHK55lp8CcfDs5KTvEi
W+3ASODoOD5NC3FzlZFrHTzMuy6MJxLWNDSoPocBdQgmqTnMzK1OKatvMHofo3cSUyVC9ZzvipeD
crlT5EM5FyAD0les8Dh2lUxa279Z45HO2eSQ7h34xAbArlyF9Twyx2xDbDlrWE9KX/S7Gz0tNixb
BqGocazury5anr/7qHUYDk49S+I/CiskYXO2/rpKGy33wkoE/b+OfK5WqhTgbuSd0H40iBb430Vo
QaJjeX+IsSn7VsUMLY5p7pm7v2pap+VVZs4fXKTxZnVO3xOJurs5nxtvWNrhRDWa7GCsgj7r14Ug
IPo3X2AuwRtdua7VZMEfrPtGDB0RcFk1wQTrcP+831Em3yyKBX2FCZJ7BwMHDzYJuMuUZ5p8tp02
n51WfMd/fvr8Egmnmr6kj/r7lVBNWezTCAyJE16AZtNU9uYYMJPAiTHcS4ms3rfO+mTMjorxBk7c
bS6Fg0zE59ckDN3TS7T89ckouKr3R3CCYz9CuR8nFpB+YqNWjJUnac+mLfYVSzcdNNyCKGCYDBev
AiuqJd82uvgQw5k6VVeV26qGqHJm90DqmNQmIPxH2TtNi+1P/FA9jz6gqwkeBLjV88KuOVFtgxOE
bGrC8kf9FTK07X9CnS2i5ToIpNC/ggOjw5Bwqxn7MoppEepbL7tmmN07U/uJaCp2Q7T7zHPfskHv
xnR3kAaO6JpVehJduQNZW0lyMxLhS/f3hwBLLBUI75iVfrcZWQOnVK4Ie6j6wx2KAQhZ4tHW3sHk
ySOnxJshKyQKdXJo2iKCBjfZfl/4BcUGr70+4bdvynK95RlKOIIeL2F9q69FsRCHyrfBFRxQNPBb
2D2ngyxklUM01Qh38I5hIr1oe/M+YA7Jw5hBdbhBHOQGJ5vvCP0GvfGMlrB/y+AtoSgpuzrU9tNx
NW6hcuPfskeFOXd+No6fZmQv86bwZskq7zXOPtBy8NGQQT74eQ2nUlXi8jWw1grZO1bjnbZIowa2
GPiYwfiUXpDXWOmXDJ18Ya96N9Qyex+vN+jguJWMhkqru/emNJE8QyMB13sphh6gOShHFXZ3ATow
ZRHJ4q88bVBDAoaDzF6zCeCw6IWhhfN5lkQWFOgAqFU6f8R64Gp3gFrHDHaucdCFDp4RqWtS5jse
YWqZM0axP/6tpNiFUhLynh4xIqf+QK8QCa0u+aHzqJVcD8o12X8HOH86l8jLUOplzPIyrn5EiqtB
TR9+tpkXvblQsyX0BmETxYUy5XMisOLkBLP9DX4IKHJvOIsgCcNLZ2hoOX8cN8fvl5Bu38FrwV60
va4I6CZcw8cULZRWhGXpt9fklzS5z75+9s033acJRhAGIxtz0WuTd9vOw4eSjLL2iGuQ02C9kxd5
xaJ4ruhE6FeTcp4aUIhQxqb+I0UHJfAwZ2ioB/k+5yLLWUzkpkRkZIdW8/Kl6EBvGyd/+tXJek/r
n/vkqF1FfVBBF+dSSxJcchOK5/+p0IU6uJnQhgqrbS6vvfsahaxOcW4ZUhGdU9cmF9lmVBJP2cJM
Co9dRTOUlrAVfjhHvrSf6apWORcVgbqAuHnwkpaFjmnJxav3UalnHLaHblJtMkYra/ExcGTkyEKf
gCl+aVsJm2DAmXGGRDn6MAt2PM5TvSgLr/CSMvSg2uevh9sWemftqRX27727Mw26CP/5XTmKFQtf
AXUa7/kzUmzJhlTpHhtrB4yM99/wM5MM7Ll6e9XvPccw20O9SDxTlatvgcWt8LT1JKhqPJyE3Rpm
0moGDIMTUZ7SchUfuBD4iNNUwTYjlFRp/72z0TXt7/o0+WYZzFC/RBP/D5OQAcBoqGAYVzLWSTMW
TE/GbxuLoibZVOsu7qVq/S/1FxNBhvpfmm/Y/f/esHOoatG6hdTSjQye4Dd7KdTWZwGhNmRXFWrK
a8S3VoMRfguFiDOdDIkqHzHq2hlYXAJhGJjz1KpukIdYPb3gMNtuDQc/yfdkEmCJ/EJuh2kELaGa
S5O8f2PY6T+sf2lkdI3wcVTh0gYvCSUk2Q0LvHJOZQ1B8xmI1ipD5pYW7teNB8LHqHCvtZ8ibJB2
AZR6mG92HOarvEEGpn11b/3Uv5uxY+p4Ci8WEdpJPW64QbKSPbD7L3RJGyWo/wRH+XosOWPJZMka
0J5Io5mPZNStMPjDYWsogukgQPdKibcpBDMx4FhoeRRwyMMUERXBymSj50CyRJLq6IiU6A7D1GBU
49jdiY+FLdWY3OOpaJjNVElTHG9tlR8Vj8egF3WIj+41jg1rUVsuStxbYAWWM8EF0VqoA2x1pLQ6
UpHcFQ6ymyIPAFu8UDOYQW0ujeqqCumUGh+AJsSfsZjCMMOeOI6jRXtNWcIvO/62SYyT57KRCfcY
aQ0vuRBujRvkbVLfRWXGcdjpqfIYM8Oipkw0itKVEu/BFxaUljbm5yRQUHnve7kUuVdC6a068va7
WEO6wspR5G8bRQdH8WySeYI4Vu5ChSOC16scqP8vtGIw/IMRW07I/xAe13bQyG1n+/LU0R0FQSpF
HYolejckfosrxM2jsw1LZEuVZ9nOjY67Q0+OJ/CeKHq9uoUxmN6oINYahSqM0pcfQ6Wns+kw0g2I
9XlrFKKyMD4PZ/u9n4KIlifSbNRK7vhQfpUw9Op5IBa+0vvDjJVjTY/bFct8YLWVrpwA6C/oWtMm
KGjj+zzrgk2iTFkiWBF6Q4gw6BMSJGwj2DmtghIsEFOt56+y5LsfVFUM+6sUBiWoxwq8aAenpO9t
m251Ss5hR1VfPZuPue3WPnxRmnCW5UvTf5vpVQdmQnKcXPsX+mjVc3n7GTHyaAqLgpnVXCIurqDR
r9S7DdAYjA0VT7Q2ZyJf3LFtulbkpxNK1+d7lx4XIp5dC6olxfaSOOwzYwRSN7IqemBvNPGeZ+Km
/BAiIkVVVe0+IgK8L0oXy05zvgt03RJaM/4AGiRUSnbAM5pgrkqvR6ZVDrh+0+bRcV3b8gkfVlqS
2zfdNIXP6xqY3ed7A6sGLwa/gDTgPDSmbxaf7LCE1RtqsXCWbgmbilDxjCuG50oCdVYrCxbA7Q8+
NSlwg4wu/t6nXKlKAfuZ9JMy/6sR/LZYYTUnaX18gi9RbTB4g5Eb0Du/lOIodHZ+HOWlRR0S3ICB
ogu6PsOxxEg+FzPJPVSfEoQCSo13WctsvfC/cWM5Y2swKGOS/BK89wI1EdatNCtkyzEfrSIoVAPr
VMzXTobqCx7LFKA58upnTetXbRB0k5cnp011O8E2ltQ0PCXMU3z/6vkizq3zNdsQE+qFctgqPl1u
i7Gwoum4caLb16nOiMfw0wkXgSXEaLN2vkvVg/T6luZ2irwqH0b2GcJF4pxXdXZpCcpklA4rODJK
ZlB+yQ4ES5ulrYifiHDLH+BSozN+jkV3eLZExIDjgmIf5YqQptqFWYI6euslQm05yigP6t0eCYWY
X9C1A3o5rPa1JXfg1kWCbLQf4/9DtMYSMnbK3KiJpJYU9YphjO1y+zLduMLRRFS+MA9JgshKFKpm
8Ftqkn9qOXnabLx75xzay+F/aqNwe0slZUpU7yMGCJ0NVkxMEoW3cMJXqGDlJxQo+CIEzpXf+tNk
stah3W6UdNjXlkHEVk8wbJLvf8UJZRhHgZ/qrMgvHA3vaMJqPGd9fV0z5F4s0CpXgfr7REAibN+f
j51EMzPyKoA6nbj6PW97FiAW4eSxKBROB5s+ETg//fHtyzp6ETT1wBcQ51OX0nApBi4/WAmV7rTs
QcICdyALqfamGKs5pu3fC7jEQt+6aRZGiN04KMyKAa87G4B3Kj7Zshc+IK8jvmnzFVuEZs9yFkNb
VUTcS3OyJE+5mBcR2tHK1JBpC/yh//nmVaeFUwsacbgQ9qx2DesUXhHe7jDKcsZASMEDO2l3Ahxc
++qdz725u3UxdI2PViWqLK2sgdqqfb3w5WhLKkTINFRnbHSHSb7fqnmAmp+7udR+/gLrxzG9mwm+
9xFzZyxXaCqz16MMOftxq7KpAD1AblCoCj05cH3p10H16JGYo/Z9NoDIC7Nc2WcrdvOeE0omT0Ll
naENjTcboKnTPIM+WqIcbTQNYIWGq4rmQHJN38zH/Q4TGiBEdG/fDerw5y+P68RovGADAOAsWnJi
efkw4jWVC/fxR+k+MiOJj7d6bfzxvXOouzziGg0h+A3U1R6vKbM6Z/j0ID76eNxL0eAYDOMBPXNm
r0gLsNoGiTXiyfyVPdFV1w16Zy5DjXTPlUCLmqVRWIvGYRAZP0m1F0hSaCodEpmL7wM2bDBjsnmS
rIgTIyY+NE5c5UpOa2xLH7n+z6X9paRZIkdJZX1YgaS2JLGxZA86aWLfNMa5wyl3KX4DUfEir40N
mHs70F4pDdV3N1Nq9NxtpKeVA5VGeJiHVQR4frOojL98Uf4D9mBYRo/QxCbzP5QiH3LLzLbiTS4T
MIO1u0XsS5DqwrmznD5fopDMklF9kGdEM+QMBkMAs6Y+d5NtlLvIYCxcT2qnKDeaVEaGxcIi9MsN
oRAPlGDfF95ow1kYeNW8QJS7EhLQ/HrdG0+0JuXs2GLcC2CIC0Dug39KLfa2lPUW3uTpzv7ppYIo
tzuxlvFt2nighIY6/1Ko1NEPTXrdNUEDHG/dsxNsypN0o6v9uHJzr5Req8uQoQR7fW8VMBtfZ7Z6
HHtiO3B6JCYXPS6uKGTxFOCtMehKDFuDJfEU1oBmjxTzh5FCTpnAjL8FbaaZz28FsAn/8gwMgAeg
6RoJKkpf3gQLGxs1lo4SkW4eIIozWmV7vXlyE28O/1MfbA5HFMjLNJGdJfMy5ld85hnh+q8qmUJd
4iX59BhqGolcwaCST8hiW6Lp/FyR4c9LvrtYmnbvil5M4f2JRNeS2l5H2F9vr8e+9GVN39FMPkbo
Ja29OMZ+q11CZ6f5PhCgmF/Ip5dk87YEi8ta1/nRGLAS1SGJnzMX2enKq7k922Ykeddq0atrEDbi
1DFDBHfhJ0ZZVMcwkH8edtuR6ejgKXPKTAhTGMZGHksEmNRkdz0NcGPT/7dzTHZCO9Lgziq24k0w
ZzPBrqQrVXl5Ul9t3OPq1BLV9aqrOgUFAdzp15Z0B3pHwgbeyhkH44vPX7J32bhEMx0H9kxSkOe0
oynng/XWKzur8962ijZagHFI+IUnLWnZ/lY+QXtnNZ4NdkDU64/Y9He/TH+9wO+1uL/QhtHh3n8Y
Xcre6eY12nrQBbCIaaPV5b0v248au2nQHLnaAuZGUT+sRfS8RAEAl8mB/lsX8MTGU0DqJ1ZqF8nI
6cIyRaO76aXt5i/Ctah8ZruNCfsc40Fmgd+0Gsq4B2TjoUs4j15goS9ypJs9aIxoFOSHHTT3HTCK
XgL2AJZcjNVd01G53MzWiyPZnOiIaBuekqlfZNyS3YIgyC25dyZVX37fqbU8p1XRse04FNE/oXn+
uyvxnE6lcCUJyCx8+JtbD9esvoj9CD6RZw/XzPCGLQxdQatwEhzirv8TeqCfUhJBQzi2sX4IMa1h
d6HvXmkAPYgeHAsVCS8dbp0Qxj5vnrVt2YrXsYCEhem9u0YjsZoVIO04qln18GZbxQ6t3oT7gyf/
WPEiTH6JxJvBXPaht6Qnt3WzvIOx/XGxBrep0uPQKaGisEJpCkA8ERqgOv1CD1bVgwTsSBFAtsSG
N8qI36oRLGgYiFypshATyeiv3dN3LEeSP5LpCpp/BV7EBigydQaWSkPCmTqCaZjvXNQ58M+L7Ise
Si4n8YwKRhNxcWmN9pln+0WaBPZw7SwHN53XYFV+DCc0kNldgMzc0ElB3kP40wQfO9gCOjDTA/aY
G2q/39r+mbz9YqdihdGp8HRadc90jkvVaQjiydi298o1g29RgBDqyBLxbm5sUFlIXcELXiPoQAXH
wbABUxgQz4cB9u181lO8PbvyMTnr4Vg4AgCZuQ9aH+XKa/WDgbfMqStDmPPVTtGzOBCtQFLlPOwT
fm9X2Rb2VwN/rQouVNL5GojhbH1ELfYcABYb5zqY+9URytnvY+ASPjhcBNNV0hRSxccIOJQlsltl
yIDFZZTGibqsoy7i/Dun6PEhKl8gg7HTV6IHRExmjvPgils/+8Kr0oXqhhRUUUZry3bcmlc6Lv2g
uDr3dVc7jgu/eNSNI9fxkO86XYNIOSUBKNtvrx2OeKugUEIhq020fE1IHeIgnZUNKuWHG+8GoGZF
3haSGtCeP22CjgUvLEY/dW9HnacZSugFPiufSbuac1hibZ16N1r1n6ZH0Zpop7lBrERwzLTnTmg7
ZSxFM00B3cKOZ8mNmUr5qst9wbY4zChIeMgucnyQddvO5oCWUgAVLblM2mzsmNIwqJYumh0ROI4v
xyWccTAuV/lPRjR8gB0o0tXPOHlJSiy2OFe+1DPSV8z/xKAo/dVtu4+BBShG7USSJW0wgnvJ6K6y
cmQTCQfr9scDAvASJ/gZwyN8bd7rz8AkyM2CB0Df99/pXVKMEunH64ernmYaKaTxr+eq4/EOkCCg
hhyKHXSbs6dHEErrzBJFZPA0T1mUIDfaLAji3m0FQsP8W1jKJL8cT/iLaxT9/96uOHwzIoLTayx9
yEw0dyiJPlbMz0tIQZ1rOg9xh2PBlPEbk879bF7GEW05JzgcYbcB8LoeTZIw1/o93mtTmPQ7xjIQ
GMaHzvoKspZY+VIIIZ4G/eoTVo/Im44pZQl8k6Dcwcabl6phSR86Ae2Lc6X984in4q0LFQ43oR1w
89rs7VLaiHpflr8AR0CvICSTyjiy6HoD9MpXeVKQO64+U8KGZwMc00bUbv/+VV+f2QOCt63iBnOv
s6PuXSlPaMCDIrM93dce5slkFIioZ7NCudb/fnGx+7axCUtqkOsBc0HkRiz2IjAqYKyXG5QoQas1
zk3elj5rCgECefDZfaGcXsxm3grv8OineYQ5aRbkU/qZwwBP1H20wAvF/m2sWk8NyzQ7Ezkryszx
Mqqi1x/STeoHfHIAsoeqIOsf49N62Fv80XrylDd1hNFn+iGdBVco91zOHSX0bC9oHm9jkaWXZ3Af
jaDjF9E5mP6QjJPLK9p19uO9sAuNoSUPLPX8AchGNW+Y31lLQJTzXRjjIKay1sAJHmPjuf+tL5t8
GRW3bqZNbUNLJqcg/DFK6JX/ciZ2nxy8bfs3UsatckY1KlAC8XQbJ3weuNH9xybnF2l0knyPw/+3
D9fCFItcAU8VbZ00xyUs35vdTFtjO8BoYWYG3ZSDFieeSJxeiQ30RIbaqW6vFNg+zZOv5SduEdCV
LVGrU6evqrMe3LJbXgpUxys2y5RQNDcDLY3qJgLyrGmlGM8GEgptStnK9OgCTtMRujOaoqIwLamF
5OYnCfpEHVwfT7DT4vV22nIWtIc3u84PxEq6jhxSY3XnMQd+leHrStYmleV3RtdPpWxGpXrCx/3f
Yv5G7BdGRTdYtk3TMeJD458tVJnfOob1aKd+OogQaJMCDFScK9N+iPsdqMLDEgffzLq0i2f5C/Fc
j4181SdK1RkyjHSCWIQ4130jxPbpKYpAmSnboSW8I2/HmZP/fqSGP2snwHBA6nmz1O5q6aRJhSkV
34NRwiypQNsWENwdf5DRuWWWnmutb5WxT2rC2NxD/M9LiUdRKXK8n2h1gJn5Of28ZkDGDA/NbxlX
f+5BVNb10ZezolORDRQ17VVJp9JWYvSb1hOeeW1fhkm17hXxhTNAXzdVP9PyIBJRI4t8iWRy45ry
mcRnoc+G+fmtl05fmxSUsVaP5lIq9FtpGoqPPKFdTKvrt775USe3n3Ok30KwlYeAuswjcFJaHlJz
K3cxzjMxskIZT39XRO8cJd+Dgo9a0R23pka4BTelCwz43aFOvhla31TBqZUQjC+Jd+h55NHQt3fQ
beH+GjayZpKdGho1jEk0ITc63pOikpPTD3eTmiYC3CESv+htTE/AqkyV5IoqLbNUcT3IWrNqdkzu
LbEea9hgFXQFPtXoEYgA+Hks+LJf1oI4aKY88O+7bON0kxJYAU5Q6wr4YBREtcXFhCFWT+AFV41n
D/fX3z5xIKBsL36BjmUGFoPL00fEJ866i3aFssBPRpZJarFYx3s/BWTtYHtqYfweAmRt509vFw1X
z+5CStHAU5+8YKIpOMgJpE4KNLAeE5p3yDH1QWfXnZ8CDwPatG0TzUl5UKjK6G6ORG5oc0C+n3Mb
0fNo+nPQkiptsO92sa/rZsNse5noNufPVXnkX0sQxD7bZ3UNVln0YHuzTykfji7DCjR1h3m43oLk
GxmknMaKAr8Gst4H5iop94RTanWhfK+uu9Kq3y6h/p1bGcvifWLO123NUYWdGSCrwBT4a+PQH7p+
6+N2lffaOyRaglpyn+OMfWvDt9t9tbJExFnFZaC+o5aexGIrYc+xvhQqoHbJKIzkQaS/qIUPgQiM
FbM/c1xVjbvx56o6lQli5WBYlpOHm/8Cn4UxSDpOE3zUCp872ZfUV5XFZ9OU5nB6Cw3lcO/hp2cG
HUho5X+blHRyn8RJqiu1ospWjvaO55w/4G6lLCP+9UUlqQxBdAZcAtQn9oL1zrXFz0Chd+TmHfuB
gQHdXGLfwWM0Es/AM/J1hJR/sb8A1FNFm9/47AV0bImq3kSjtwr/SOoaEh9u58GFfIr7QWpgAWOX
JRy0Yl3vv+Wk/ur5l7mv1Uw3Rvpiw2i9lmFJPeoE6m9PTNGMDKntLQ7vAfiabLpf7bJi1dCJWJtV
0klHMwLn0xY0ZFhs9GZJXwsxfp0uWh840nSsSTK8wuaJB1PY32QtA4AN2gYkk60xrWoZ3JjvjW5X
Wdm8NfGvdu7QsrlT2xdUvbYQjbJQ71IHWToptJ9WwajpHTG/JmYNs3UUBGvwzas5tP5M7NInZebl
+o7/P7hSljx/8WuT56zm2RUOEilwD2+44jMjafft/G+ZUKx/ekvofIV6x69AQENFqYv1oO1rtqVc
FXojPi3kSt732VxcqZmOH1osBEIfpJenTJLJy4Cl2bEWzQz3nRxRVMlk1/5nJYhb/HgNXyzxZL1E
lrm92SrE2ekfQs6tMOy59NdIb9LydlT5sb2Ddg5k5Xyi+HaCdKBh9m2bE7mY2Ic0XyXrCYFQ/+e1
GFnv37JXUC4wM9KolbrwaVNl3znWKpRXtZOHedovZE2ql1sXyXq7NbapnacHvUJYNGLyA1ZyHiA6
dDDG4qWItKl1yDe864aHcGtjnrFx8dMTi7DWg3ZLTXhbdUc2ymtxkcKmQYxyq/La8euI1AQDcrDs
lyJjPcYimWHRxMbgZBMTmBspdrMUqclEQ21j9Yr3vt7YzLT6vBWS2DJSawsAjdwnly8bDEVfDlSh
+W4uhQdhcG30zo8rGyxDYDKqBofiiON32LGXDB+uygut2RviqSu8ycJzO8ObMYSM3llaJWW3TzMC
47tN2PyCxmz3teHNweqidwvnmFly9BjEppeK8iqBK1xmP6AnfQRguWktBk1ma5pTR309C5LJ6D1u
c2djnFqDnjjtlifsiCFXrw5hspUu8rFY6mjz/2CD6dV+j6SQZcZPvTOD1lppgtmdhOlN0GwgULHU
m0dSdlnhL9T6wy+sjrEI8rTzMYUOWZ0Oaxy7BlgtdveXjcJNboMn9nJ0Pqfdq+u4b5kFAgLOTsgU
1fq2muugmMG5pS7oocS80gKJwvE9CdDMvY1clG/vFgeWSuaSQTjIJtvKRqk9WKWEWCYLgUHJ9Okt
YMMPjbHYDR0z55Rffu6f8PEO1QWK3eRPAJH6kaytU64Yy/uAEzd1v6iNbJs4mkUnzodxftbw+Hhw
YgPVfxG9XKlMnRvPs3gjf1obfKQOW5SCHcmvq5J/OTafpadkOp8byEp3r81oYo0ZJVJ2JlRK41ml
VT9xymKngP870YX58Jp/+sZQ3ewmSx8CUpZ81l920iKr9LxuLqxZRqr3P0pZ+oc2l6Yv/DCjoiT8
IMjWRqItg228FMxAly9j21z45pynRMAGP4R5O86uYbE9O0vAyAKPmsPC/sDH70drDYhwYoFsqI+u
TLW6Ah3Py/KnPieum16Aky1svVPRmg6kAVe4BykNCoeyI2P2EFUHb32Lfl00pSPVkXA0wXy5WeZE
FlmHb40pA0OnLxNwaARnDEP+ZC16p+y+GlxGqAIrxc31Ep8yJon8RwxSXk+u0cQIvSL/HrsFSwkl
ZQFfm/HSEkB7HXsNr084J6kJJdMf+M4m0P36JjogZD4mGo7zKVajMFFOPfyH5POn3A6dJuGNBK+K
0M4t57AGQzl+GuMJOtj1mPSdTfMUuXT+TtpY3Xa3jAi2V/bHwccfSMkw9ZmhYhRT5AOhIvNRhsSg
5pbW9XK4askiQm4DK8QQlWsmWN8bueZG6TdSxZGzUNPhy2jKBioluYz1Kmg5ySjEKRIgbPa+5IzW
w9nJ7CO7z/AYEqudkNZK/oWwYR+nE2Lzy09A0O56KCkFSw4HxgzsGqDCEpiI77rn+yRoPOJo1DmX
tH25VjUR8PO/4IpjjqvMjdmnqDW9hmqCwPw/Oj8HeG5oRXuUBd+hTtfhJ1CWHxvAFwdd3tbMKgyy
Y2ECUxc1dnTX90ollyRLf4Gvgqb+FUy7HnrSWbsL+6BaTRai6kq6n0lcmuVp/W9T05isSGxIgwQx
nCGEkygfBj0B6ZgBws9y7hwFM9/WO/d1NLYwYf7PE89Ualfh93gyD6WqyystOnL4DcVD8oD9ReHW
qBw4CA+MUgwqnqAuOfZRi+UTKduD9Rs1EQAsg6yco6HYWj2mE4Thzn0GZmYu693HHgfWPiSPkgpK
aFoUeEUsL9645JXhi7rMlORzHhuA72DN1cw+TufptKBP5BjJNHM6HIASHC86jJR3peQQWHwft+Lq
Vm8nA5M9v/r9SDavgheKow1/L9YiSqdCx1HM5qGuKUaQH3kJGRRVStdJICC9BLvCQDPXXMk5tEIR
yLqjFCbeXWVlo9mrDj917GwFCHXwnP4dl4KSAv1TeQlN5bBccUi63c6QlYtIg4N7vBOTdvHyg/1O
EiFmdFrP5bXgKIYRaWGD372rbMqIg7BE5kzsbv82yyf/g0w/RVcf/iXxUUKGT1pXXzfBszzQIZa6
r2xG7LGzNhsY5PsuAZQLOQonDwvHsolUGmBkVpN+E6+Mm+go+pHWG0I0H6QCBIvlHe4JS3ZqGE11
go4k1HcL//1l2vMgdtCpOQjuQSaWOafaMEXX6YeUl9eCJGf0JWk9ncmW1HSW0/qOCCPgL5AS1OsU
ESa9Egu+5v2v9NOe7glF3ufA43xub1RHIeZxTQH8PqwOZrfn/Rn8nqH7EUXUSQDW/CFEdSPui27B
SPpDwjzbI19cnnt7hb7tTzh8sW7JwPNup/EjUoq3bjRd2klj7DlczqCTd4elb2zS9t2hGPsTftso
Z0CI6cIcVsnBjIn+nje9cEDaiSqgB5cdCOay2Pd2FrCFYqrTNprn0/SgVh6rVtJUqHfkseeuyFmo
gG8Wn75u+R2nYaD8Upycb6UnEYD4L9WjfXfGxYez1ahBmlH7LaDRSUpexLP1Nr/excibJR8nxEhx
JfRofHVAfoczi55SuU0AKtPWRaTt+w9523AwY8yw67cqKx6kM8OKNf/2ZR0Wpr8ELRpoz2EaA5hX
uCiOrtNakZpzrF269u7SWqRZOOX/aia8HE17tAhx24gxrEBIYT9D3kczJ4rjEjnciZWWTbeFbiZe
qV9Ugz9qxDbNcupKImVY5eX5lvJcLKjhG1gZE8NdoYzpUDXy+Za6KO7TK50wS8JPsJLDveb0gYTO
Zl/0RT0fKVvm8QYYOXiassL7F2WzMzQ2C80RO/qM16TUtJzMA6UBc/rj2qc1NB1kgayLivOXhLms
kwIjQjzXF9aJhCBV7CO90ekWeeQjNtKpPVnIAmXyV72N52ziVXce461WfHN0cKolAQsGFJFnDlye
CeCmfiBeuyS/yBA5L3a7q/wT3Y3+a8mTRkLeoLlZ4udk2N4NR5i8UdJDQ3lmH/wplP6aVXIORCVG
gdiUoO7+SN8uyf5dyW1aswRokX0aIvY+WPJSGnXPTCTYbvJMkNYqyg1qCtUWnHLgLNOTBFp/abf1
xWIOvy+YgVlZX9JIT4axeSuzXdM03867IQHxcpoXEgRmksrPDtuVHQpzgsQTbG6nfHyTpo/Vlb4a
o2n4dkhfgdkw129W+jWT2TAflz+K3FmY+2iUxTpH+mO0Q1wAInqMnHZ+kBKDx3H0RBDc1sR1dSWb
A4dt8TCxZGEGsH2e5zKdLn88zzm6xhjrc259FsLjR2zbUaZYfo8w3kATn3X28Ph2vI57hkTaIBnc
xgw+xk1+8cQOeBaza8LalXoAg02IZVlH8m5FwKMUX/OLIWvBAqBAT25osnUH7Z1UHi9hCW2Mr0Fn
1AM1Kf97StsGI+1YMNic4O2J3RAdWJXJSPuV29Q0dfwqbaI+nNiAGdPanv0mXtj7x4F9JfImMkx1
Sq8B9uy5Lj6Vskl6JeUBnNsqlhzzj33OvTGVBlED6KqMYoWEgNdiNwsO+NJxN6ACXQRl63+izerF
2Lq364cqlN/6qI1uA5gp/zrWDkrtsKBcTMpSBUaxdeGZF55amlP23fu+4TSIVAaq0iUKDUn/r5B6
KjIHZv0gA/ByW/6ktWDlhYQlkZZSO03L9BFczGo465vN8q/26Wn3Xusg1OIcQBG7vjxwoXJb5gQG
SQq7g9Uense8rKgfr0gpjKQg93U/X3plHxZd0KEyVWZrM07t+UTjH02b58YcoPzr/CZEZD5QNsMl
NE0Eu6dEJnPYYouZ4PkotRgJb1rBKoNPfXdYVFpZmGgV95u47xfXqppuhAe/VHcSKV+hjBgqXBx0
D6ICokC+Orqswtrt5svxix/10xW+RVYWiz+DVKm2f+fwjxSm4DYKS30UmoP9rQxdBolGzvU5fNhg
irRT6MeF6R9TOMAiV/fxBcO8oW8pBq6nRNFLD+hVOZbAfcbfcr4Mu34Otvq+kqw8ok3jDK8r3qod
gmG99PSQ6CTP9vmkGVGHztwK4q6D6/uIjJ7FVz85owDwmdfri+5Tidtmm5iK1DQPTgIDMT7K747L
zmUyHsZ+47XAHoAd8KR0H1TACtsbY7Z7bNwJtPGl0nZfA//VX8zAvoMsyZKHJe0KXK1GDBzD3deC
r0KDE651X9mqCTiXu6f/yGVOKe2ttC3NCJjvK2xegHymtjo+RrCEYzm6lZgAjLpDy2nRWhrJR3My
tUcQolm2rT6oMFhnn2tHQZWkkp3OrhkGeXcmvYQx198q1gZJ2aUc1XVrVndmqxipUOm5K6qkBTES
zYWFgbUD2cbkTaXNsWcSg9viishP+TBXxQ3ZXMVAoqdvFBUGS8JDsOR5t88IGO7JBleCU6DyAIQw
4Sv+/IP13dobtgIxtutEWd/Vmkst23L/wl75ZjrTyy3AY/Mw3tVMOaa8guzFnH2DhchDnd0Jhldp
7ojsysfGmUrp1YtfRMvbJqV5yl0/VsQAuQDr2kWDSHhta7ipG1BoI6Jq/F8K6PQx//7VMFEKVnkr
TRKKLuXaDT0/fwc1rWAyWMItzNujNvJNqWDtpaI6hEOPEa6+sLPB1YYMlb6Xdi4t/iLfOknQI40q
bZVCm1T2L7HRG6OdLqngNVs+9MkO2TP2iCpJygAFg4GWAzjFjofajwhbwM0STx6NtzCbpOmJHQq+
txAoHkq0Ti/FXMRu0Nf/wTWgpGGjCvS5FDRO2pDv8WkRShVA6uI1F94nzK6u/XOf2AQWKcKlA5jP
Dqm7kbQrI/ieLT42pVEduDHI9V7HKE5NQbZDfp2Obu+AhGe5h8DFgKAlDj+ujn0tbwCVyJYGGaU+
ElIuxLoqkxWPbGdZREh6Wri672bEl2LpmTjnmI2srQfYPyKIR/hooRU8SYTLrTlYu8OMB65T4Srh
xg2E6aGbEenK2GYpohgC6gxb4WDktV4HepjWrOJ2zKwS7fwjcktkmcsYEYLt9VfXq1Ir98KF1Isb
22xC1u8CrO8IE2lbFE12P/ncQ+zim+3G1wGzl6iO+AeK8I/2ZqbqPJgBzMZZ7LlZZ7W2nDD+wKm5
DydNw0tcKML3B4HYPCpDtxNl5RZmdEwL6UeludoN4Ocf/VbRcl/iykSMXeTeI9BonoEq2x7rsBnB
9b0+h2vXckrr/2SQDryhIM5JciXpO1E/KblqX1G6twKUTl+tm4tftZhL64oAas4tvvaOuc4jfRuJ
0YrivQb8bHTUs8KE9vncbnM8Ryb0SqblHPPGVsZpWRgePr/3xSr/hpXkRfom8qkeKW7BXnIIGdcM
Favip21dsGWuUXaTh+CnFx8SYmfeTWIzIOJsrr+z380/wQCtYo9icjMo1ogG+HWngRuRVrJqpi6M
qYQCHmBv78VRZtGhhDDWSIvOpKeO5i8+2Bf3WFIS/oRz3KdQ7m6gYjSnT82VteZCOSJLq6SOFmA5
RqQr9J3f4H1gb3tynGr/pi2C9/UYgB1lu2pEqb85KTAjjdkz6eywhuShzySIISwKI9lSWeKciOdu
twC5sz0GpGfySsbSfBZ9ZqY9dzL/7xaeTbKjYWF/sv+L+p3kM2QRzpxOUFIEbWszKa5estqiAhLq
ycGluaxoz4ORnowptHosWa9p7M+AAawQ+HbtciU7ptiVNDbbkZ/MzLmU0XsPuSQzez5TRt5wOESr
v/EnHLv1pT2Z9EgB2DBgZqKXlaqQssBHEfwGphFBGUt5YrvDYCURIhXQGwNP5Nilt7Ed8S/g9DXU
gcBSaasdx+0ziFGFC+T9POUELROdDQWt9hEnJGzmBL4VBRza3dO9xJiQfSySC20BxNDcsHS1lP1J
tC6Qw6TUuFZKKx2m23dGOxuekm9lSbjsnnU6Qd1oVAzVPlun5+8MHH8ub8hcd5XofbrOvTtXBot7
cJGY3aHLsL+16B5i6sb8ytQ57qylwcQJzbNwxmHREP0w8/TpZAvNZ9VzXWDaJTCNyf8HmdWugPJz
bdissJnFKBWe5yRJ2tQUEoDapfNTQT6lfwHPgOPxdcN9/RBVz/9try/+2QrILKcsklctjnL3eGdu
ATa7vV1WNFmOWTRNTW93BeEq5DW3PGM46xllXinT8i1MyyvFAtt9L7MHeS2zIGgbxpB4jK5y2lAe
BmIQILk8B0h69l+myGdcpv2ojMYN7CLwOt0gqqG9YYU/Q5YIMLxPG/v5MS2qmT8+M8gcil/OBG4b
lVMbDnN5isuH/dHmoKQSg5N7s8VivylT5Ljc1PbhBLD8s+GA7GlPqqji4cFaeS4geWQ6g1D+htz+
FogVRUVRQXusoZsUoy80CGZr5cGLepuQVCqDD9Gl4lEeDe9RZgPtg1EtDbcpz8JPWtxUkhFfulqu
VQcG37cZoH1ILDXiqCUZP/mJcfykMtSWsW8QWiwb5+8CI8MKT7Gi4qfNk7EdHq4VQa8rlIkwNxwV
prT5ZJtzUdTez/HsKtKNRFmLItXxVZb/srflrv+Hev8exa+hecxKZfIK+8HSc1Y0+HD0qz3g/0vn
WklSbjEsViKCWz0/yoe5926iGpwXNTZtGcIPgENZlL9B6yVq16ct28G+dqrHTSpG6Y3teKkFhAp9
003Jc3l7sRcuNrfQO3Hw/xuhKxMi0cMLIgdfxltfidgHIRTgDM1eyozXUr+0orNTFYdRnfOoBpzx
MmlZxtn4AsK6rb2z/j0fDDzIUgNNkAlRXUtwaNh55iWNW9MYKvNhM0ORwF5hMUusUowAn0ItmA4/
iPT09QIBWiOJQFiyFV7PsNP/f1Mnioy3nP0gNS14yaub2TJITdDMFqu3D76m4DRB7sIlDkpsUyUM
uBBQSf7peuzDG+IdcfEJ/CVRLjIVDER2UVZoHlRACd89cWH7pDA+5XuM+yHYcEtfoLiocRwJLx2w
8tZdZwLyjHrudZUMIsN/G2onyJd9Y0NkbMnyXTxfZ55xpfkoVmGo1dVGHA4SiqNioO2TukVXDBSt
0K//LA2OycDCfrWw1dnNdTq2aaqcWbw4TNjYFpQ6Bv+nT+TZ11ue9pHs5cEUerTXtdJ9iya3ZMbf
JL0eaqo2fY3IHvr/3QclJRGLXYjtGwznighp9Pnp8OpcmuywI29bDNrj6EIQD3S7rUy9qRaeQfnU
W8dGn4/3rN3lwjLEGx554UfWvd6sU85382pyDKFGV30SmcOdyxMc6JkWN8ajg9L24iu4frVRuIJn
BwRdH5Kwh2l9RUpHxPLqlJK8Zj2BFxb2wSCubMham5ZNhx2fKmcIz3t5RoKsK04xzYL1e9aOrD8F
gMyZtFLR/yxkg7AktbCflHR43X/sggQnv2OKJ4eNw+Y0VovdT4kiaKfwsH+ZOMv/xW1p2W09YQod
3VPxoQE2+jbDFzlaHopfzsbpqxrUPSqilj5OF01wZBbxz573/qlW5nszr4CdJlp7CVlSJzvl4QcB
9yKhbJHJNy9533O67Rlkh+s8QqxmMqXMizvgjwdb3iDRPqkKl6aItE9MyEopOYG+JzdC5OvLQKnn
MfsbvETPtpzaW9qS2xXM6vvrTkSwlwYYGNEcZiTV/a7hwjqTVx8U2P1duKFjEI7RSjJqQPhkPFY0
KMU8YPuWe8sNaD2GXjpp+JLPXr7HiKJttAv4nGSfU3xN5WA/XiKq5EApbWEZ3ot5Rvr0rZ5eOjc4
3G4nQsrU3CxBYnEcH7dW8fw9KyotSX6YoBaLnFYRo+wPidlet1U5LuyXFr8AspeiO9GneDfYWeiW
+Gs3IxY4RtJXBWbYxO3NIELaajy0khMXpC4XLRXSNh6vJnmJGcJG2/keFlCLUPXV9MbJAMVkWH2n
9+vfvZuKkWDIHkdGmn22ML3smyrknZRGkgaENmbA9Ax+gAMxF02xr9WBircIEDMeyLkhshxrZcmd
t9y+1YKbNR6GYaUu7g5GTT4NtFlj9pce2cTR0+XCqglxSKV0GmUN/8ofVntQSVW3ArLbERHw853d
J8MkrvuGysHvgJrfF7cL1zVL7oofS8S0FQJRi4yc2YOu3xDoyxKEb8ikhVRTFAKxDswf9aajn2iY
jo8pxN6sE2mcHtmBKj5WgfxiFgh4kc9xTaSQN44IVFXRFofF8Xi8THEBLFKH4/TcABomcKfFYlEA
pbGz1uMCJy8l7nSbwCuusqdSq8tl8QWZ5HymOCA0EXU45QEXpvBLLPtwkmY6qvVLycxiT2k+19aH
0CwU8IqLDL3+d1EXUMFYBbRlcpdjg/VoWlLLcpWcfQNgAQungCICQv5WsaE3wC19OVkJQLKpu9rd
8SLdR1nM1EqVw3fe+cZseC1r4FfV90nJlL6qYUldBbqKKzT1HBRUtaLWRS9fO82Cv+zWZbzO/Slk
mpF1ikupl9JstvqLCNg6c5OqtMVjiilZ6GWrXMnLd6+eYPnm2rkAIVortPRh77ZaRzd5/liI5OlX
imQKf8MJREho7vOWAj/xKVOvjFVTxNnJFna69kaVIpJo3VTX0MzTBKjJvwY/rDJS2g8ZwDIjg2Pu
pKgu51necWt2eg7j6ZY23G0caHPWQwjkfOU0Ntkr2t34T3OypnV5QdVYw9xyHs70rKR68rXkoizq
6oETY4tdOtRHignGWS/+Zsx+3xejC76FoLUH5u69A0oQ0uzv4sLknTJqZfLwzbmjqaMKDxiCKY0S
X1bFflmFk/+igvpDJQ+SA0bB7bMX4i5jvBJdJvOIdgZs1rYRfRhIUofUo1aaegG7ViGwDCIdUSF6
qEm64+QTeJOxlr99mefpKNlptGYUZ4hTOoe0/SQeqisPT+qA9v94tk5tf/P0JjbLScwRFMBB/22Z
YAVBE5BzbI/5sZDT3leUD90AcQ8XTZuD6eSUgQrne/vRTfXm69kOMHDTXhd7bYho+xQXDGSTZ+yy
Q8tVZfsiq1Z+9Ozg+j6Tmk9K0tojhi2s2tpIUmmd+XLuOFr7M67RPbNDENZwHCqfdeD0avr2zRhD
q7SFcOISOU1Fmq7MQW2a8brQ+gQ26ocAtfxiHlqE878g61tUCEefkp/pqY3W5w8Rcyn8F6xlC4kF
P+dGrf63A2b05Tcx1rEECAPHhbXuYRnkXrKGiAf5vyXI40Stag9rtuqMoAhE80IIm3T1yYb0KfPA
zm3pF8TlehA2ZsVopwFzZyfdj6OLNIit15poiSPCS7vfG4K7oNQiVTO+smXRE1m5Uik/yraZRqwx
EUfFt3sFnP8mIjxv6cZZb6elHqa/Fc4YaXsa+PCM2GZYgcKpPXfBxHy7LoP+K4B7JBFmMgveRP4u
LteMppr9P9PGLzLuWrFBX8peiK5vujV4jTFAlXhaDJuKK4jnLAVUrDoW/iXSH/H897hOhOczYrpl
uC9odj5prRmtgwoYjLJ9pDjU7J6LIPk5PkRDTZ7ijl4DfubdmjaOk2od3JlW2018jdNd1+D7rZBa
A4wQaoBjpu6+VcdKrov6EEGxZULrG9x2k5hBQsjUI8crOlKUTfbl4pFXpKihoYux/5WW0mBfYrVr
ElfE9ZyKaBlh5bDuXzQ7fNZuxTz0K+lnaeTlA3a94x71+RsVTlZa5OCujcMvfZ6btx5ArBm8JMMf
rOMKVa8Y8obXFBgPiKkuoQ8fqKhh02dItsgOWNf+BIDIEBK8VK7CGmioAZVrW+4szYwtlNS5wsk0
Qucmi0E44hLZQfYQpQn8aomZLYXGtl20Up2bxPnmm1yihYa9jnpMq1RuDCrEcAmvX871GDHMY05G
XsUO05t5axkLa9ZL9G85n8OvBBqtBdbeUH5+nr1KOrHmOAz7OG0zgTdFdnuNfBRMnh0/IngWQuc8
opILqzBdmuUs+MintKa+r0wFKfRKxysr+l5PteY94mhbCWlq/m+1p6wOI0LiQaK8hNP7bRRE52c8
e6plOY6kPFOZd0KH/K/M1vo6Pt8UVvySIQ2CHXPGk3sVNTRzBf2e3nsPML6a9HMISomJWAZ4b5TH
Ru5jJdNl6oOIN68ikylDfdjHt75q1Gt3EK9E40l5EoAVlUsNS7xRWElJp7goUZ67u0yZuG8vxSuv
HAS2e0wJst4pypYDhuoGNK7GdDCUa6Fm6xhbcvCJtZJvjU9p9xJklw8loXiYv7J99aNn1mo7+/vm
c1gl+xI2Guu/M6snr3TZ7O5dyN84r4zAszI9WqqOOuVBV9uo0WqsT38+k8E8RQDx+FB258FWDJSn
s1LVqjk0NBj6QK6o5Pn590VuT0HV2SCLGkuVKCn/rwRZJPkorAQum6ni6E8NXftQONF0F0DV+gkt
5ssWX0grgWHjT2mh+IZp8l13zWpJUAw2PjKUnadxmsSoKjt1Bb1l3+xbzprieKSY8Jt4oJxE15MO
aDXuYaEBLGVFf1EPPJz8e/FcnNdvTzceznwMdFpaOOb/ZruVvYAzN3C9kcM4gF0GSMRgoqvUqGtA
2PDMWgioJdkyFDLS+xM8i93YQllzosYF7Y2RNuNHt/MaY9iqUfUXdxgwnItqqS4YlKZGa7NNnX+u
fSE1esRNB0rk0aPdXdSBPM+Rn6L+c7Knmgfjgimx3GIKjGlXxYi697DDrVSSEF5eFer1vqnmdqQO
0H/thR2pszTg7WuuN7r3kU61GQ8CxvGsS92ZVxRYz0BBK47gXNGxR2SMOTj9uieN22lrgM551dsH
Eo/CLthaZyqNx4qnub07ROg0eHul0EQNDdwe8XcE5XouKjET+g74BRpTCpqWnxf1uCWISX/64eZI
U1lau8Wpnu9PvBfOvuqNGjBxTmATnpN2TqeCDpvVz7YqNwze3kEKSZDWu0k5hBfM8jnQSqFnqaLS
P4TLC9Q9KJBUsgTlejy3Mu3vToQbflMqmdD+rA6X5s8kJCfUVN7eB7riDFXW8mz+ftQOTVA7tQI1
j1bAu6dDpZN2KsCDC4ZUKBSN9bzcnroaWe3zFUM6dn9atc1V5YblOt0y7VHxFzWXTZSB8UUUUvPh
VbZSKbf72vejWBxw0vLXVBM53UhDF9W9Y6ee8gezyIyW+JsZcJbn3QP6ds74YtQg0YbfeHT10aUv
3KUVbCBFAY4/Y6ZGNQx3joBwNLyzYad62nj3y50TdE4e+0+urqFRs96p0JrcA3TUQaCVos3agPrS
QsRgVIocZgVEPoav1qj6sRrXK/iyeWNrpieedtbUDCoXekhUSYSa7n5hw2w574k5pP8ZfmSoPW/n
LJf/IVd7lY7fBRhVrvG8blpDU6snSLA/J0piaYYrbPDJXWxF0kWe9M6uCnQk/d1N92ShF0MZe/GQ
a+4iGNY+YicHBsO9Zl7tDQBqB7jQ4udXm0JZmY1dYisnOtZ6Po1ON5DrgWQM+qyKojYujOHmYsW2
GYlRC7aOG8vAL93GYyf6B+5+QuX0+RvD5pMnTC+tZqQuvD28bNoFbipYe/5jNCPR3e2SVOgS8hh0
GesRclNHI3V/jvuxQoNc4XycBBvN+UklXqbr1wCod+Ix+jkQ47soVqz3rmJIeHpMwDCo8qo0g+Wk
FNFlxixJ/+3DHoImYdZ5ISRE1c7kriStNGuexd+CO1TV+QrUOrXZTc97p58+1ky66xu73dQyQRtu
Bsc3GVtLlpZVE5C8VZanwxfDojJj/5q5qdxFbjTBRx1aAuTEyB2GjIuiZTuSWBQkIYNB1Gixqzu2
cUjTuQC6qhkeriX51DknGeyMsrbLwTrTetA08we0/+07HWipZUCVQ0yFt8QyqU2ooA6bMvhYJeco
xZkiHntc6LO2FTjhQVzfQdc0JUMVUYh3Cd8lcQmEVa4gOgrF6BWssZp4IdjQWgc9H5g48QEulvSD
ua1G9QnQ5MwpaNg6v44Dc9Eio2j6b3aj1AQ3qpKgmkKCDx/2BxKo3O5pyxci8qhAwSRKW7dEwXk6
QJFZ398FZKnAWe9oljYg+CcKlTXvII9d6d7mCmOyI888hqTJ+swWGKMvY0KOuNo4/V/n5TzqPXjO
MCc/v2NFC+jqcqvazK5e/+snpBKnnrztX6WxQfUzpKw1z0VQ2H204z81zMXCchoCL5COvfVcL4l5
u/tfRND6TW68fvIPFMIewLwD3wjG+1IDjlJim/dA8TBgc4seTFoIuQI5QLqJ6c+tnvL7fMOEsik7
9R5QYGHJB7Fb2XoWypeKpcA5KsKZThNVzfCKvfktqre/6YAn3Ze95WRBznUhk6nrAKRxbgSupsJv
UOXrhDleuGvnrbh222S2Ap7ydsKlBL7mb+ermunjRLr9sPlbHpgbPpTupABoTLMdioTi3CEmvgS8
yXPZMdHRSlk8xQUj0d2Dz2OCLjTo+G5iZHLhNhaAr0XLA7tjiIwXNsYUl0cJmdeWjsErkqi1JAw3
SwjiHh/2ioYeytlkYfhOvK2Gc6WIocBetHSKfWn6rYBizuQM+Kn5s+nyNzITQE7Z/y8fAUUpU4Hp
na4Iheq8qzBk+XLr94WuYiwrX/qeXCtJKXiYETO3hri6UbPR1C26R+AsbtJSYCNS/jTfU6Pi9jQo
neHcMKjiQ9HlJNnAK6XbS0++iENTvZLZsKfbqI1H/b4v+bt8Htd7QE4Q9Z6zzW1dzD91mJWBgwpT
PyOFCXsyHE3QSJnHY7jS/AEXD/eDrzbokR/GkAalKos4fXTEk2rKAhzc6+hFkS4jyyah51k0Hd93
ClY2DqhqIDPQ8otRKv7SDOyAJJF12vuYQbY0PJrzhNO5H2L+in3KeAWZ974w5TNnR3qKBP72oxCi
X0FmOKDb54Y1doe+S2wzioCbal5vVw74eEcSaoDbYUAf7EB3myA6xkapUUHDnWEObzxXtQjttEYF
gO9AYv/Q4c2Fc2bx+Rv0jmKv2fZEFfuzIgevINKiMc/fswXNYIJnqYpV2AogghepnhOtWd4fL4sX
EoaJS7rQ0s3G/v1QjrwXD372m07R//GCLlmROcoCrye/jo1ww1Oywg4SiEuE+IcaYVpku9wN/bGZ
7ILA7lIA3uvS1d1s30XTemrNMca2YzDBqcSG+tvpjAE4g0fSZfPEvcb3jvyPaYD3b88RGJ5K8YPB
FTbMNfTSi6QJH4bJ/+UOhORd9AFNfPJeX0yUC/0eY3v6VZvV/slypgE0yKmCFK/g6O0yjIJk/YKe
Dakc6kK8NvTq3GekfSDWQ6N0F20IBDWSP3IcUNAhM0gonE7aOjT6qtGy0jkk+9PvFqdeHOUkNF8i
nbpUlnETuxGxjD/VrmQCfSaJXuN/aJNFOjOaWq8koL+AIt4lneYjk2gsJY+kyfIdbaKb/EMyHxbz
JRseZsHZB+jzJo5Bo33Sz0OMmSstos3tyvVHBLukEUcKMZhBe4DnMoq8s8H/tDJA7WY64Zdbc3k8
jrAfW73zpNlHaqjtvVFYSC1hnUI8FpfELKKFtU9/pS8cCYdB2IhY52BlayUV3RZ414PhM/GZl7FL
fWqqASA6oYPipy8c92byXoByAtJtRr94icecDGucVTD/LYbM2UvUj3jRls6Rer0Nsbn0YkVA2Sto
ZB/HxW4iOdjjMMUeuYSjtztU0UyMGD207iu2JoIpSBopxw1drKfi+jCfxIboxfqkOqKqir+BkkjA
KL8ZVJjXp5nWRkqyvCZ0y118GVJ5h0ctirDaoPsioI2yVF65z1grfYoP91EadKwYo21SfffreHJz
gltSPXocUOsk8JiWxPmFFZeeoShSDiFEw1wohE9WNeuYnxbMhG0gwaVvsUmoGM+8NS6DXLYR2s/0
bw4o43gBh3mtmZKRgnqJYU6UEeeh9iLj1a1cMCHSY8xy0n+KtlXoHF/t5v/JXgJ+sNnA+IojIYPm
WKEothU9WJY16TmTHy9IcpbhJyaSNGrFvYwivlow2LOkKZQb2aDyr6/TAxsoEEG3YeHYMVb18kqF
5t+yJz764sQFgSMT3tOYFy6HQbpu0Szj8UQpNdBo1SysB1L3ZfdaXNfKKgle0QW9Z8P03qj7k25n
w9h2UMtXO+ukhF1lu82znFDpNZWttb5jfBXUv0N6ECbmg83YkHGr0jcWfC2qZuHRzp4eqAXzT08w
/zpygyj5HVpjbvYti5q/bStd49GlTq37am62fPSHnWeunb8LFqKYP818cpeiU8H/Hdkl5Va6nFc6
lGZmGb5syPxTnaYi1jrySBJCnGVKgNecn27S7R5XU5aDRcfD28QTyzuxVE+h2GunXEklh72ddgBs
btMxwWo6k4K9mRYz2cdaTbIH1vSYj3fBD0cciyaHdj+K1+RYNgX+0LqjT6pYqgLkpXXhZevyQ1er
ID+guAyShsMastOclusnV0870IIpL4U4hJitiH51xjzrcm++8j2qCUI+pIGxfMRqjo4QYENs0KkN
1w5dvmIjLfhEg3kHn12CRF5fq0ZNjXCtUtfJPrjvunx6DGqP5GJTxzTKIvaYTfzP8Z3RsS0820on
xm5P/zfsxGsTcdthRQ+CI7gtkVIBmSfWyA/YtEASa8J8nPuGb6GxdWl2bZo5dxmjjULaVKkiSIu6
kvTX2N7K6Cfv7DRiizLPbFX/eGWhT63h1hM7IcEg53EJO+AbVT+/6yLuB11yi5HAksBd5IKmMp7g
/OTpA3zHCXThKTqlTB9Ri5o/dDUO37KTwRnRHWlD1KDuQ2hFQ+15eS3hICbgU7ErTen0OcgvayWP
KxiLA+D99tb+liFW36CpS106NEmS6m0Vr0JB/b1YQBM0rrQIEvMY5IOZynUEGtTSFjh7oSyCG3Ad
zIX47cZKR/lGzUmhEMOdL4cKNuyiP2eEVsXSypTAW0h/q1A7D4W2tt8nZE7ajJ9dGql+ctHcmgLq
R+sdd/3/nH21E6vKemJJSkYpPvs6eSMMIZPNdckQjkVzsLust0E8H+SCnTYW/y53NGRnojMcIdVf
QAY493PFfS7PEMfqFaR/xCKiy7mG/FR7N1BDftDwemoz/2es3Mcd2rJggRjtxFklSR7ErfKJx4BN
X+K/r7WfOMD0lLhZnutROU91L/0EoZxQBWG3R85EH4DRdONhcoB7ZV05xPkT7C+ltKcTDGkLt60D
1QAkrE/1Ihiqbu2xbWYzw+my9kG+qnKzCAE1p+8Ml8RUB+iyTi/VFNzIm7Js1LX8pbvhdba7sP4l
LZQwD1Nev0uzQYbSjRzejrfILB+qZ8G+XeHA5jk3CIvRNkLedUjR3K0+RDKk9WcmC43xSqyhnIoW
JzTxBqFMccuCCRz+yliL5eg7mu7f/VKPKPJbyG/kKZxDAeh15eR06webNFbia9yFBKgHvCJ8n13i
9YU5TCRERlIrELiZ6Hb0qqtX4oT5KDTBRhBzqL+tJ9UJwuxlFRo7aUDSdk9Kox7FAOk/3OLgGd8N
v1yZFaS3jcgPSqXqDuRnS/nHX9p4ckJZkS8rUOZ7c91CXldZCjpoiVbIs0IyQ4Grm6wE90nvJ+b7
e7zmcGpzYCCdgVwlD6q5l1eghWVys3J/RLRltiv7TShIGpgTl50mdIWH8E+f+rtsDqfm1hknKsmt
NbfJSWZO08I0nrVqAx5AMb0mLaO+xnf8OZ7i5K+PFjcbe7lBrkMaGSn5hZIdtqH+Xdn7z7D1uiuP
HWdodxT57ooGgy8x4IOT/XFmrPV1f1AV5Z10RxvmYZqfEPrv3f8rz5oWx6Z6LHtp51OShVe2dDjB
Q+KSCO6OkfndZk7xRB9ct9teVCCU6a9LjDxl9lTCtdysRHQvRDpqZmn42DT14MLKXLE1farBqnWY
7b+dza14nx6b4VCcw6uzsrqKaUlMUZH8Ssnbyx4uqiFEvH/MbYxoN0YQgGm8Bkrx2s44t7j+srZx
HK2l9jaTZ21yiIVCWdILMedB2Y1sXxwKTl/lzSGM75QVGDFBZgd8khxnVVb4WP/yRJCZ+CdbsGdD
glwJ0uUF9Kq5zgrIGDHtETSrTx8xp4Wcv6sQWW9R/zuobrxCRb9gzp/RF4EI21I9bGuKm5lRWuI5
YR8xEJvHgRppurqGgyJIXXm6KC6ojqNch2NrE1zW/ucfV6kb5UZiMosAAgJnlWwYlAqh6oXnigEf
zctmAPuDwpjjq2oT68Br5y5pHSKYt8YSU7cM6LurtlwbrlOs0xuoV8bimcrvPzI/MZGnJlqtPNHv
fiiYWZ6lAmwLVvvEkD75CMXCRU9m/EKfK6Mhe+NPPZML8GeVTb0/2ueK7BQIRumZj29b+r2t5BjA
X8LRWnxDLvrWo7cu3ITYGWF/amrVrFi8Pd0rQBAHDo0H1Nqj7uzIBnyaFadGlvWC+kA6li/C3/xu
kzo+pses9kMr4GZwqwF/0Vb8tH8vWSdR/6ok+fSGVGrCO3pzxvhOWLrQdhUTun9EK/cMikPFtAuk
rp1u0/APGlqpR8THBzVpSOYZOoBEsm3emi8wNMbp8vkNj/Nbf+UtrKRUrFtUe08x5M2Gy/Fp2hie
wVt76ZPHvZFO0R5aM3fTq0t9tRJVmJAIa+T11h6mhIjR4BNv9/rMBDnRbUuboiVmKrXHJEuKytC6
hZliOBaRBb9qhkIOX8qMbW8f/mRomsq+/2ShCliGQCZcnesYT820YE2WWcKOM0w9NPvjLTys8lLD
he0D7E6UTuKSV4l4zKhOE8MpAhPGGLNJX3Z8vj2NQxf9p1kgMcciNTj62lUA1LvPJwvyT3PRXQ64
sLsHdz1nVsPTyv/YkHBzcwrzvpG33Q6fPzxbB03OhqrMeIlqDH5YCqtgfi4ZMqLODn7eh936ZAfo
38yPJUFff697cey3UD+EZMkjnZHPOJR0XeeAk7xBmskoRzxcmukOS+qqu92F9wqCucexi3Tlj/tt
UB31Eq/AilS+1onFR5uli9khmxVUhKmLkMSnAROvkBN4LChcpuZGGhUZovYGF5uWxA8poNCtEsOv
dl5aYOoJ+rWwunxa51ptmLBV0zuDXhwXgFqqBOviKKCCU7rCW8/Lmj97YhiNyaNJWjytjaJoUHVC
JkoloWzNMeDSnT34D6OOpEGRTo3FxA3jupKKDkBgAEZms4J9xkxZVCuFkuqgzYzpX1rH17u0CinH
GOqgJltQzySE/6q+JMbKOfMNIlz7acK3mkLGUFNEtyynpmuWDj/vbegna9aAiXcg3psN/yLPTsv4
h9kOiYa8CnguMEUv2buVsGNdOSx9VMouxOHJktMDGgR2DyKT1B2MOe7ihcXhuWR30fBh/KTSJcZj
aRayQL87TGvqVqVFNMp56m64Ghrpfx17pIHn2jopdKBQBPscLPqiuvh/BY9ZIYwbeNGpUifCy3wt
W5vq8rFBJolwviH3GYoBZRaumj0S6Ub7F88sLARmoLbRNwedLFYNmWClBDQ6xwH7eeltecGFHxZf
Ppc52kaFSJiS7SHCKhjgsYZPq+rhuYLLgabzvI7jJr7FSilefnYh0hnSajtTf+Vv4mj6dertPi9L
Ye9Phcn54BhTT8xnWIWnLCTxsCu+NT/+0z737zp5sZx42rcLJkNIdaAI7XDAgFJjtJvDXdthNhE0
3PJ5tplGtAnSxd3P+Sa2Pog8jg90dk5HOHC+4/td/kb3+Ty0WLOqfuEBDakSaRSoboQrX+qkgEbE
954t+snCyVkXw2TobvDes0fYc/GwvlGBFrnAt1IDdRyL/wJvEs8wqIAtdIuzbTusRGXu+u8d0jbp
n0QPCkLNwDNRpTlOKVFSFdeWkC5CRKShrgHSw/0/lQvG4tSCl1pxuCI5hLjjsXwrsb3nSvGq8EAL
77CXFklDNjwmlbpgCYMrhD9hJwTlefG9xHuPLj7zBhRACQn2KSmSD0GW5P9Bw5iQAA7xl5CfgGPu
r1JBsPKvjjVKqSF9WseCeRr24ll3sF6HK6bdtb6HMhHQyhxtGlDrH6ZBSqD7x5dLcqQ8v8OziOq1
8O9H4T8qEv//ewqlwySDYT6YJX1ASxXXqcxP9EyaGmzX3dCQJt+E/WfJ1ic12+uAIMSHwp5HKIvH
amISayORhGM9Q/qEBihYY8pPSL42HGCo0Io8hIr1nVDCd+yCZ7ukna3Y5TqtKVYoi/xA65RnVAdr
NVrUilczEtsxuP0b4Kag1JmZCUY0BkdtzgRZ1dybdLN5lcNkrZvQg1g0OQ55P0ahedgkPLx9949n
cnDrgz51XW/lYir2t9TzMigxTGGw2ZHbB79KvCmCu13rq5rzBXKN9Pm6yOUqKSymUZ8I0Jwfj6NY
IKLBsAWQb4zBVk8aHMw/tFRouDq+iQKNKtSGPzlsvvOnY3nGY5Q80hyLvjqtltfRmMPIX0AODrqV
x5s4oMNzNHAqqaBqMpnPmvUH5XWp8BbAs++5rdwJMlnzhAssE4RN94MThWljHWz/yKPhdMphQ9k7
GiCzHMWvVM949DTGaihu8FALTUU8lnBiVlIUGVy1lqBE5DIYVpmjs60BjOQvlQTnVlFK33dCOEpe
grHL/bmIvcJ8q84WmKaEu77QAgitklrGXlctGAfi7WdA4DnxE+kvN5PFwBaunfGZUiQhoXslpjmY
tlfI2gE2ZegveNppcmCGnhszlbzCzBHloe0QV0JiHhTlfbbhRGx0hvIkk4VAgQ3tLn9ZD5ltO9Ki
GgeEFoDzhyve7sBapxtSTfJzJrnQ9dju25SDIUeHpmKhtZwsODpLKTEmW6qU5wAVtQO12hHoq+ps
FUbmc5ugCJ8zG2sz6rkLcmM8X1s6iAJmENNNlXqSGVvgeU3e3gD9lCuGShyW2H5/5m/FLabJm9T0
GR+uKNf85yz7EGzFqEEOOZtXumKKctGp9pySnoqquBauCgnP4Vq5HR+X+M/fzPOe6JBKeUqB7LVm
m7cQjbsm5bhWpN+Arin16WuHN4wkeGI4VkPoaBbJh8k/ylKojq5Lqnk8anJnUq5yjWvJSQOy+CWg
wNUN0cYjlAY3f4fZ6OV7pP0HsbiGVuAw8NzxBge2ogyAUSvCx3g3HyaRLjsqQY6r6MBZFhPKx+kC
C/aCv7pMG7FFb2ie+wuan1hmRR6BV4ODyEKGBkCYMIiSq447Ij9pl9VtEQ3IL04KFeyB+d6zN9TL
jEeNu/wD5O2rGCmGvnyi4zvZqZM/t2P7AdLDm0lwf0ianpCbxHKNsXVAaodfI4+SJtvz/vTBYGqW
NU3FYsY6AKgRrWG7VNNi+IJHtSxze97F1ImpZNyguSmjrhn5DnjbIkM19ijN1qQGNOArNAawm/CY
AymLBivdRJ3vIZK+S4PRoVI6BU+AGiUgGsBxKibLLobBbtG8EnZ7mtupJWZZTtHVgzsRiaVzI/3g
KAuu0TwmA8I4LUlNXITXgbAPBZZHUNLoqYn5W4ZBC0+KoO05y1st6ObIvnbiYD70Y/qiOybygfDE
DzFEAq+ZyC5KTKrD87i9nVrdtR+WhsvXHgyzkQGAGSKvSnr8opXkWQSjAMDCxLSl86MwIRXocj9A
2QGblwxWe/efUCkrmXb8mH6qEp21qW9wCc3JUrJsJIz0Up82JYIt4gHCL3+iky4qgpsvKSNMIEdx
CWWAEaTBkXqz/KXn6Ff4mgTKUNMTa4u9OBR+QqklZI9UQCPwDhFGt+Y5uStgGkwJXVb8lA+F40bv
2pkiI6DzQp+8FXxgNpga/W1ilbM/EGHQbu5EAdjUVXZZRSDC+jHLp6u5pPZBvdH96xnzVkwY9P6N
Nu6PEpbQcCqPecndB/FYnkh+ZkfMfyPWwkNqd0yaRGaf+/KVP4NSkQh9pxPQWRKgHyMNm2I328DV
se7QfZzCV/usS4X3D5LfHmd6M7uo5SzIEzOXXV1bmxZha4WMB/0w8lFpEbntyfiFECJ13z1Cl2fE
f+Ecw0XvunfAdJAHiI5U03afJhdpqDnALL9nSkMwIOHmjF5Din/YsW1ZwfTTbiBPnIhMxy8vhTVy
FPjzHlLGoJLAbshs9tCVnyiH5IKVLJJCA1JZQYot21YI0g46jj02HwLNn2XzHYy5RjxRXaxllEiO
xwzK5wJltunXwzTp5GjF85UbtUhJ6cr1neD3Tz8G0ep1zC12hlJIa8OBseAPcve+SJIoXrqhjB5G
R6fmvjHzMwnOBvNuuEOn+Mpzh0HDxtJwEXBJsB7ADo50kLuzEKf/K3zTs+s8rfioycaL0N003/QU
tgyS6GnyAqTQu93gZV5aMQwoJ4SsUXLlI8Ixl0Ns/ITamOwBnIqdR+1xeN03GfzFoN2JZk76u5tN
hu1K4IxQVz8gNmLBDl+hnjOK+vlvhJCpuwap/SLLeVV0THMC+2ULlJvlm33c4Geib57Gtkhm+Ao0
0SAWyOe/A4cr7TBuLNhLBYoR3YDdscCE4X1sypXIZKeDDUEpO0mnxzIMMJHyGNLvNlmVy49PWJWX
OJBeZ5g4b4ctGfQ02ohj1mxc2VvgebE7uJFngX3fFDzZNT7ThCzvkPfI5N9PBt9ZeOX+osjI7rLm
cyZf8MKqTm2egWOtiVBBK/qo55d8UoArw/NGIFBFUM5/qNmyFZnmxFP8tpN8I09daxUdXrGm0KgN
hZLqiE/EOWzV0nGd+Q1tLWprNj9W4UFhFLKsxqqd5vuPi+gZlMNIWRiWWFShSLsMaT/hqaO0VuSj
1dcj3YYdzYv+NJYbcBYS4kBZTKu9rg9bM+DurKJSkPjQg356hv5wNQTUjDXvc+zudK83KPq6CMjh
EVQWpaxO93oblPcx5VHPCjCicJ84odWM4Jb31sNjEDQbY4OIlUukCSKsvIqPy94z10oRkRPHmhzw
3GhQ+vg3PIp4glmYIDRcY98xzfdRRIiVROc86yEXbNevH+tgyVaalEpQCdbGm3yxhzNiPh3Z+d+6
LURYCiC80qHbXai16FyOooMBIEXAiAa4LfNVRr886xfrKiLvo2B1WyWA+ladAG272uaRnL8glUmS
BJHZKlmtzHeXSclYQCzJtPCZCew7zwRzaWJqC9zPM/sgY0Bvql556eLbQN5Ghdjb9RXyBoc6MYo1
YBsSRKoP57bP4mq/P4vGJG2/Jbpzxo6Rl9E5yIgXXxXrw86ZE5ch/NifitsPXZs3UPTTXdn4aynJ
nRwkwIEZh/1BbhDqmP0y0CnEvgpmRnu9U8u/fDbLH/ZfNqhdCctbIshXFPgMIDofju569Uo4bR5k
wuWQsOCx9wXHBNoM1D6jz6sapdvFiqpoz1rdXemfLOx/eIe4fwBMreP9527jlTxeKLPIenE2qWQB
ADV10yLW8C1dim0XDviR2FEF4d7o3NMKTxRiuggPRLnLDgLn6A+BWV8lWCBHIXN9bXTWnC0VsjVs
Ctx8Jq6lEP94XazWt+ZSelRmp2Tor4i42IS6hBOfbPUNIU3g8v6/RJnwK48uWoKDbJLTWQImtRT/
mQjWJkiGRsR5tyByM/XxnEWsKBzGqpoDX+rEIztacfxUL0k6+HbtWzapnpjUj1IEoR5thyeqxbt6
itCDPGkzYK0LgLLNQOYVjeuyZ+aEtUmDlk7fvyWraCV6bjvVEB+ZPxJZ+wO63LWwmllgNysspACT
US0j98Yg1RVi++nOnfG6mgiPCjXxPEM/ayPc7qszZsV7NV7PZ/d0t5uJ4uoftuJ798vaGjy3n1wA
zIVVhZIMLdKDEeB15Rsdz2amyCa5wKyIad2tz8xGKyjqnFIT35n5zXVNTpv5aTnDaGPWfDMSYIlD
c0RS48Zk4ApPy4DNFYnuDJjW/ZycGYRAWyi5az0nk9atbAlmogwfcPAKJ5vpDaDhzMLryfO+tAZJ
kqAfaRyOU0ab9+nh7XR/Nwb9xhahgnC5TIcGCSDlQBlIanb9yCV5MGxLqSzLVMx5L2OOdKunwnWz
RUne8sUYS+zkEz2KhDcXFFSsUVdl+GdhywvNnC5Za9CmjMleF2qW3HliGm1Go/R3mdh0w/wijzzN
4IzCdto0I4/eR+XxyszCPUokDEWta1vJti/+lf78kK/JYcEmZ1WZWitv8uUrZxZMi5Ek90A39TDG
Xs14Pug5zQMyhbaNu4sTXcvEdK/s+NPrgA6jy5GNBg363xoSjYMqdpBE8g9idWixKlJNQcUNso5u
1LH2O7cCf3k/kSDsCbEQ0xe1wh6fLZO5+exzu1+ZLpdnjuu1kszZm2chrdBuOUYsBVkHkPw9E0Xw
qJax9nF5odsnBoPn3Z4lBZ0pIioU9zJJThtdmcmpsPWBhFpHhYdP1o0k6f9bKX9tdraE0qEw2H4+
c7kaTwOSvxKc+odfkGBO5A5xFE2j3AeGHdju8JYtJAw/Q/HVM7NYfzgQ/Cb9b9jeq+h7SfwKS0ay
9535ShwuVjTRjQS3ihuke85OyMlkO3Z5ll9OWwNc0KmTg5S6+/WVgAyABcNGMgBi8Mrsx1qKocv1
9fW2Tt6rZPPxKmHOTenWlRMDy59NSdNwBbYEpDhTTmbV5TKlmpYIkKt8W5lkS3ZMY3hUsT/mQXSt
K2gum/dsi2xOGFuKW2+5N5+9DaVU8J7IwwBa2H362SwSlxWdHNiH3MOTtnFax6f4DzRllaxdQtAZ
Y8dVeOtrAOKFjPD9XPcbI6j710TTVlSeXzTxC430qUMY1Y2SIZiQV9xBQ93+k9trHzHAIEupumFy
NAM4fSMJW4oa9e3/s7aB3KreNAcUtp61i9ZODml23AUJaOo6bQ6WppaMkt3Yma76mhN406MhL4Ff
yhC7z9y7ly628Mk6bjSMftQtBiMypCZBTHVQHwTIfu51Im5hShKDKELVGTO9ywQFFWM4wANapS4i
J08eYUcurckNnwaQNBM+MvQwcg18RS9DxgJf0C5vYz/XjxbOB7fgEKqzlm8N/chKURJl1LOrQfQ4
TRh8Ukgmfe3KMshow9mb0ChJKLudT4xtgQc0V7VADUuA2Vkk91O44uxCfOfinG1olSz+K0YXVNoh
UrPR4cxvdLwNn3oa/QfsVdjzLqnMsiLtdxBcmWFT2mEJeDVi/6nfDkpZsq/EMLxy+shjNf+ir/ss
N/zO36qWM37qfjn6NKDJ6TwdOo37nbcr6s6FCPDF1sH05CcujIPRTeP79ftoL12fsB2Hy9Y/Ip8i
DeTSrZnJ07QFpekHOx2c+d4alqEFW7trucky2KvBysP9WIB9EYg8ukR0G6lgyPpSaUcng+hUP2es
g8o/G0P+X2+DTRr1ZN93DaojdemVlEWO0hi1wcAwVdFhKhkUqF5OfA3f4qTi0p42HpB7VTnovBxI
7WjtzbchDtzlmdYs7Oq/FmLn+V1QTGNZjyTME0wS/IpulQn7EM91M8Zx1SN3e5scQQa4NhQBzQDV
UnRyEKbx33cFEsjBWgIcSuim7L/Pfri+f/eZ2pkuF/OispGqpfjxDU5BJ7k174/T6qFKFB7xKpwj
Gp4LMTtGoMKNcu6FboSFpDVG0nXfVwsdGT59k7xT5igLm82mEn6XiwTBLsdqQwS69W4n3xwBA6Nr
w6b2mR50gdh6lRxCtRwolqPyJ00aGO4PF1hmSSsMNWJDYG+wqIBSdXpbrRffmZ45dah93n6fKVRE
2bTMwvsChv0fLgb6UINySQzEtJXfjgdpuYKL7Sl9WglN2xldbkLvy5uMeWGMVREZh3Yoll9pAVcM
nBq9ek2coXDcoq8j9ue6d6+CzZdVSedO4/3QBqlrVJ7WS4UvscNxSbbFmF6hSjpJ7yt+1f7196sT
LC67L4Cmk6nU2iawjD+hwknEsPeED5rQRC/ZfaYikC1MnwAIg+1XolrBx/YpTP8p2zV66XdpI93m
skf2Lcw2A+ltaK0z+Upf5p8LDS+GlPVtxFoGx7+nKMufnBZNPPBelAoamya5juBfWXNLBiwpsKa3
oMXNCyMsn4XZbm82+y+N4BAtDjoLdrxO2LLpSLLMQZAfiwwZEHZL/0D+dIwRl8tIucAVvd8WX34T
JOOxQIuG0+NxrHQzaV8rbmhznAwHjgzOVZ5iF+J6XlEr1ml/nlPDkcN/Or22dnzFrdLGzDwRtm3s
dN/yN0ZT64wbmEYdt2WK9ZlVlTorJJfMvors+gvcjm3RbTke7XNfg851pkBP8pvPGBB8F3ztooEz
rsbGv9GDHXCppZiGY+0iLHQacuPZ6hIVenCfVKxJ7QIXa2UIwjULR9Z2teryGRzIGGGFD8nTjhZe
6du8LsqjKVOtF+qD1epQ73faxI8Ra91NE4ACWC0Qh2oPazW8ib5Wd4lZptxUu/hoasY8IIyVm6sU
PJjCxaEkMFTH8fBcbZjFnitq/AtFeS4cAyywGGEPKhoxAVehjM02o1ZcBRefB9qXb4iLY+3aXerI
k/utS7KcHuWlJERZu9w7ezx3h4WT6Fbr0QI/Bxkf3Ur+AaDc3NX+uYNJNefaTxjE32i/ffPbfnx2
sYyBY5dATpCl3+i/0XjgxeqV9/oBQjfc48MNc3LLAAyMKHw2f44YXRnXrAhsiOAqChYELLvp9oG0
WRVAT2N0Y3az/hRAWlEVouXDRNkFX/tgnThl8k7r0/t+pYFSB0XlXgc/p2d8w62dtDFgqIKl4QrU
is7C75V0T42rvtIj+Dsn+eZxI8AFK6NZHlkx2JJ9IfMtN6EcG2LOFMdZpaSZ2pwNqunX7BiiVPSE
+eqFGOnu83wekhwb0AuvVI4r6yqhhncGSZB66tH7um+O1H1GdeRUvB0Lfy+YjOD9Hg+ncmT2mwn8
jn8hZmEzDv5mK+uxCxlZzZGYvEUDazrVjembzgP6IW0YVDeX6HTd2Sob3VA/K0yTHiz0nX7//t2f
lOmNptMsHRRq/iktDDjnSNYk4Ro26dDAfIhG0gEAwxEwZOv06esWCB+Bf7B0uoKb9nHPgaVITnG/
07b4nrM3grlUny4VjKWj9DOL/qAj1v6b3BvV5Ls+7Zxd6KfbHSOXqGXzQzEjKL2bGYirDgRvZeN0
Dqhbwa5i0wTMcUKpPu+lCi2K+m3WtlPH9oSknmkGzhRpE01SYgdzj6VoCj5JOtQ1l3GMQF5TnIFS
QvmE92dtY4TVtOweypdxXILlUNxLX5McCdWq5IDiWugfBRUQnMV4QoYiLrCEW8t7U+AmJ+YH1660
legUHM1CZFRvlWzmoulFbZwPLOmqGAZZICH/ljPhRPcB+txlMD/A0JXaIAD35InmB4j9kSlcuXPX
YLzx7V/7Essc6Y0+27gBatfqn+tIgSxjX9FAhG1elsETTnNKHhPExOoADcwrxYZnY3eNRhO4eDHY
eH7tZzF3W1+7ZMi1ChMdbLhmj9P5q0L0Z3Igmr1XeYXHsYuK4MeaTmJww70hHHuuDL4IUp3hB4Tc
DWozuKEpZUQjAcWuTozVveiccrXT1576oY+5n1vI95ZsNL4sXrIAYI2DPWkgVsbp1RIb4oRrEatA
9CpI3+RQp8zjVDlMrU/yuGHB+F2Rw4KMEHWBnYSw3mRPYzDkF0KdMM3E8aTMJl3VnrttitFbcb5G
EFspO23lgVhCAOIpDKdgj72WvIyIVMp3kHfZegq3yNSm3PDGokcQl4fG0ZKGnmc6TXpHufAk+7NM
X92LeKw5jk8j6rAeUYGZqIyBL+flWoXJu3PDTszNIxW5+cQHz70CSyDbFYc1WaLHOVG8Li46Wt+o
TRgasrfMkyZsZ/kfylt8a2vVCEl6oNbQux1xKozM0FWXKmHYCpEp4vVrmEGzR1bz2lbCtOsY9mUJ
fdnBM3Sa77WhByBu2uvuTwBgCqO9POLfqN4KEzqagGBN7KMvsdLwsWbkKNY7k7Iafp4Wb4fFrQO+
5STelod9IWQMSSgyrBRf0x8KK/yz6AL0FdQWu+TdhUEHPc2Lv2gREWcqD/gRE7znrO7VdcN8GxYI
dxMYKy36DfeQwitlIaBe7U2PPrrxKhnGKw0ybwUV2CFJM2dD5AUbccNZwQPpIsLouHmyz/8DrBfw
tVs+wvoe2BSXsO2ZqYyuRzLnl5txeu/aloKsNWtS1N3+u+UmLyS7pCk1sBuhJQNeZKw5wEv7K153
UUmGvg+Nzhhvvry6w8MgUb195wzV5EtJegXcky9zHmu5iJKicgWCrsCm2P9dOs4d7M6QcRuewICL
TzYkq3yA0BM46FQrGoQdMNMoRxtjMYbHadSzCeEgkJSV6sXWayNuz+odPn49LQ/iZ7PKMIAJgM80
nJXqXkDQCNkGY1RLZrD2SMpc+eyzYMPW5Lm8i0qckwBCLWbL4T+C17RBWEfOKL4nbTK0E0pnytFD
CfejMInDTqU3XAKddeLeFB7ZIb/p27llwh4I3vyxDlW3003NDkDDUN8KE6UlUTVpkCU8b3zJoRpG
MStgSzB/XxGmh+hBmr6ztGcM2cpSGdiR2uqZTIJa1/kClCdGB+4a8CWir/YykvAhsxbzkXkgTHSc
pLgPPOL9Sj+PEmBpMihJz4Sx4WFWxVgvc11ogJl48BVrbo0a/Gj2ALGpzepWLuQ2Ha+Uxmo/0enI
9j5up8BdtH+rLoO271epDA4bWaepI9G/gNRTZOc+4sUDBpbeKGDixjryyX6ve7nVhXVOHV4nTQSa
Aru0VW8TiU7q5/LAZWUFFg3i7Vm74bXQ8kwBIQSY0zoxmQSJKcgy3Hjiv2RlBPd3/EnhpuLCUkQH
ge8wD1seIcFYPJDpe5c0/gw020NFM6lHd7HwvE3VsfzZOf4k4Rdyf8s1lvmvyTadP4VfrpIqOQE9
7zz5HfQx0ugJAGgVeDn7RUz7Xd3CHKpWZK0CVzDXs1mefwjreocTUYohjUrFQskJn61LhkWKmOSc
YUCRZGm+IfuUfLa53Qvpd2fWK1dE21vYgchM+z4MeEkvnBwBT96WzlbHaxeBywU1apv4w8k0tZ/H
uy1mnzh8pVKXpbKiJ6rIrVs1H3qqlzXl6DkILUs/fdxHGoK//LUUHKwt8nowuGTCH9SkFWuqzPAW
WYNw6Kdo3fBEi/SaYs7OzLt2WSHpH8qK7jpgeoWhOX9cG8kAFr9voe6+pM1res1btf98cIfQ70Ip
uTzkiNViqsYHyfmxWj7zGD/mpnjNfNKrSs0bKXPpyqMA4VqxlKSxzH4ezuXS18l0yCI33VWrK5tx
6KS+u1v0YSuEK4Of99lHTpq5NYU6K0a6a6qCWTOIQXe6H46AhMGdJZ8+57uyI22o+84VJDzHjPX1
NAG1V5n4WhbRBGrCcdKrpDz519MJUDsz7am95OsZO/H5KMmTwUhaBHGVijmmPBl2PzMLgnnHSv1a
QQqFI6NHMNaAngfYlsYsk1KnRIP+JRib4oHzfm7gHnoqj/2mnB4mSo2IaTtVZdX62v/v8oWhVFVm
1rNZdanneF8ICeNKEiDOIq3IeSGI0a8nbr0xfOEka7965hh6gApJmBuufBJpV/m4iO2Eqy21/S3c
uSw9ZYg9d78mtFjzdBwO0ouC9HAUgJ+wiXAnPocBueorcAd0cXtXrnRZrONRXQvQPudc+OvGnas+
861domECLfAl9I97RjHRX9OKbpTXqOwOgQlCpljUnxk1ThnWMm83hFI2PTUEoSddhf3pQ0U2hvah
YevA3URHMsm7G8PIagCdsIz5O5FAibaRCj1y41XeaQzlieVN94QKOVIYbruoQeb/4IV+hq1BKvKl
T0O1Q7d9jtGHCcG25nso2+TvNNylICp4kDm3/lhLj9PNvS46KogOvarT+J6qWXVoQwWPkF0AyHK3
cueYnUSyiokOuHvtDVp1+/BOr/X1EEIED7anYoMCBbsgYcSOJgmzwq6MSSZzOMcQSPMSftD+1Yzx
pyET+e//BzvA5uBpHdxm8wrMwYx9K9aoFTF8kdJqzhR8Ifi0UgyFfU/ly8JcoE5uAX5eHiI/9JhH
bLE7O2sfxJ0iraZzTbSkixXTBkUAYmB6dpb6adLQ3Aej3TeDMs04OXyyK1DOVK51Ven5T+UX+qpC
Ae6Run7vVShcodFW2iKm//t+Y0nCYUyV7VwWReYfvZCYL4EN1kB7UDUmDKcfMdBA0T3S+pOKObQ5
BA1jToPHg80yMuqpiaONZ/Dfivbnl6U90LCR9I+x/HO4kJEJ8kY6jRM1gzOTIn2lzFBZRYo6blHW
YpN7hrcwQ92KHXIAw/6TZD91njU5X3Jzh6STNteoyOGjQ0McWp70+G3401HVhu/ZeNTsAIORLzo7
L25bU++UjN9PulqPOYjtw0KGK8Y4u3Ja/aqcpuX4wmkryWtet0rBxXqPTqeKG5sdsJsbS65cmGsd
zMBn4hNClcm1DCiIf+K3JcChVQTxuuc9JTHQql9H31poUGyEVDtpo0W+Yv+wRvpmKQEluiUGzU9k
QoLyR5Nug+f2VBwidnBJAs66lNz61y4P5FKtc/HfjaTOY0sPvGVA1fhZwIX4FNmHd6geIUZ61Zd6
JD91FFVvqi4mFVAv+n91Hmu2Wm5yjifgKiQvHXHwZIHH1vfVWWJ4zniybrupfG93h5WFZ/6oWIWK
gNpddvUTHDH3d3Nzc+jtkcJ9SSV5qseVqJe7mf61PZB0Rv/UQLkL/XjAz5XBeoDxLRKST2KGs1HP
Kj5hKW5nQ8Jf1v2d1hTYSLRzB5SV3vHQOq1Ep9Sb9nu9HgDRnGkTpM8BLs35m9yCUled6r38tA5G
CvqvQQMRsBoq669GNMuNxN+kefXMLAeepAwedIcKYx9Z59+yreEI6Q0zh2xkDstSTvKTlmpGCzFf
w4a7ciPnED0ZG5yHaQMWgKJLqJqcn4nHAVsFBFlnyVNw+8PXTS33NI7ovoNuUYYGz7kJqEK7Nwc3
yGMA19dz870VtdheFeQxxJgrLVdUGXo2iN+k8ipNeJNU9GtlrsUFcaQovl597OxTS6i1F/XXRoWm
P+Xv9wJ3SvhyfG4SQ/BqK+e9Bm21O6AaQm2SG9qmImdgRgVWk36tK4aen+PAGVES7vECNi1nTDJq
dlAuF0NQMcrUKqXuldootcAg68K8XvC0zYO4OkW+30auDm+A+6kpZkIa/79Ka8jlwLJllm7fLPpr
7uRADTbWANklMzB+52TdQplIGW3nUrUar+wKpX/RnjPUtyPgivuAEr07gyIXKxvQFQT/qm/7wUCl
GsTTbxZYd5P4Nc3b827u487Iu8kjrFBpn/MSA6wHxLUhGmldg/gmkFKL1DYYYzB7Z5aZ/EPJ9ILV
6hfD/keLd89pLkegRhxWj7KfjfQ3MrJpCa+/IuL9kuG9zqMuDp4JjIUhBRFbQzrQ2IuMgg9pXtVT
0iBg8MKp1COrW9U22NNkh3RHT7nQCMmg40XCdMf+VDWLg42dRdPFuk3ar0Az+SE3qTFcd6VBUNOo
Ve20MYxU97pDVWjcxio8uHt73/weIbe8wGt7QD35RyiHm3naK8HEFPEDRcDyOvT7Ydi0LU2khw/p
RqlgOaUVZBkRoakn07gQL/7wZ0rJUD4EgSf6Dylu+nehkscIJDnUolhgAHJAYISJLaJLjHLbJkOZ
itoY9RTPVBWD900ruqOfRa7oup1f5FL7Cp1+Rc4KMpKyYnm0+bf3rYcXSBjIU0rxuX2UQjP8xRG6
D6d8YFZb1AIjsbHuNylmWJ5d1E41+28/UgbhHhAdkiQZz7LdDFD+ipBUeOVwUY35e+DPPc+RRCux
V6SIyK3+rEZW7jzPBLuTRnymutMm/gwURcLdL7x+Xm2rGM1kK9s14xiZYWBXIVx5NS8O6GjvQMRf
dXtI4RmM48yB6Q2R+iVaFMnS6x/WvqQQSW6YFtB8BFsbJauBTC7AREq93boXDVv15YZSIcKEYDbx
X9ylb6HGwU1keBAUVXZ70hWVmpUHAVXT8qa71Mq9TJvoi8xxdPngr0B3IZMZu7uqsFN18yOoU41j
QfJP+0D+Rlc1FaeFBUBCFgNBCRBBsvinoS7KglwKgMR3M2aZph7lv3DkwlYNzPBz+NSOCb89aZoZ
OutYWshbCOoxgN3+n3jVS0cSdSOmbKMJ7w8X/8aZY7rQ2iTJq/bfZQIjwUvB10QKnpOug3jInDfL
opajDKXUJkkhatgjd4+oh+qWeajh63yKnyHGRdVtDIFK/GeqrgnOpfk7SEDWHnVTp3KmRFvBbH6+
4O1sAPRpHq+3pRXXvBD1SUBc7X7D0Re3bG2yWXpgzr4oQlPi8COck+T4DiXOCelvW4Q6VKiXCa+u
LviGdY2MNursKzOwLFZjukQg5xyM/pafNkRxFEaClaWFDuPDo+0oB57tusUB/eA8RamU9+/0T/xY
vQqxS0wtV3TFJTbTcflai4uUGVwG+xJSlwHyv4Lp7MUXN9ZzcvWLcz59XSh7sTc7l6qT09X0Opad
EBS1bmdbvmg6G9XIhUSa4w4M08O6xVIcokKTCqyDqJZM/auEc256Mh4eJzUnLe3l+O3C09GeaF6t
tP2aJQGAS2Tu9uEBgPFH0LwE3PxL5xRyVA9tzgGGETeYFPp/F3Hh0UYbFsojddL1L830/KeRfnL8
lz3hN1tA2QG+YXyhaoT2QwERyOFzRCltX8qqm6oXKjqBmfMFAaoQ4MZ7bETn78XiuEDVhg9pbE9w
2wnzEAO2XIi0YZ1HmK/poy4X5ysObRY+0urBvBhLCMxm+KUDJ+EkAsQtQcI5aqNMWH4VK7GCj4b9
Fv+k9B/DIhDks0Uq3NYICbUEqWYl6UATRbbDkwXuSIFljy+H4RFAwaL+hh9E6wSnyE7SEpXuSBwb
Mno2yo+JrkxKV79LwxS+C1SQyPMpx9EdqgOhRmjjFYyA/jxhprY0PHvyBgB3f7I6sXDhIJw82S3r
X0G3dxrUrzML9C91zTZfX2c4snGc78OiSFLv7JJA7+2JwYD5udsXhVx6tDMDgh3ZYdoy4U+2QRka
13NrYWh3aJEMmgmsTbTtJQsi+gF+9i4aVGXWGT/rPyy/MLqrCvS2h1Z/UfuHjMSTO1xLiNOnE0uS
o4ACw26uMpFcbXkNrxzyZLOCn7T/bsN+x8Q3ClMDZLZF9H+VM1zUQrTCPTE0fY+Nvy4JuDB5KtkI
0+WtHfd2YcMryVOXMkorV0WcZrCF5J/JJ5T49DBuf7kIrLbd1EJBioQt1nMGZNmkVAR8+jhqcSj8
Li7OpVFeMX93bv+PDagRL5lSsQ+Su8sI08O5Qbdo8aGUI0I5c+S9S5FnFXY+UNQ7aaOvCk6SxqEK
gWjSNlUId2XXgAIQAMzDbPEZhHQW5rI+3Vgoq3knSnhtHY2zuFSHIBbXaN0twDy+xgK9+F4egWTv
HlSFUZgRvk/Q87OEuXyXyrgP4DInSGXoWzcVIPhfMkcRhk5vK/38ehYmnKoEZ166pHjUPBtJS2a/
ZbK/cOps6sApk1Pr9xbdkOEkmu242uptznsf6BEX1BSRPEu3jBtmSuS5X31066QVEf5fopQhxZsY
W4V/pdP4ybB24EmRjteUgywLZxTXiB6GDB2RxU5yCCtv1VSxbhXXHIJxsb+5lBliKxV27Aw7Xdez
D2dbd0ACxDyJ0ekbmdcCs2vnLb+uuYWOxZWEgVr5jy5MfJiDL+jBWEFc3lkDJ8vssh4nKJkhyHkl
XRHlZhddg4kW4PCY6DGGF2sPGFSFjx1h5USK1vgRiBfvQXm9/xSk2GM/7mVEsM5l7xKeoklM7e7r
i+z3wftngrDbO8tHAkK7pvGrGRYA9u/7B7l3IKDK9+TKdOHYXWorT2OMSyZT/lDDCOCoZoCNFI04
zni1cIHTs+pv42jbe75bDEzkJEEHyKUoZ+cIBta33TtWF5gSOnsKdUjt88+OAhmVw2pCajDEylNF
/zz0Cfv9w4iXm/wjsBdtaxaZJ3+Ud3I8gZKkTZCIbvak3hUsRit+o3iIf9LSG8W3yvdKbnroHwjv
AbjKWb4yKouNVhmOkt1AK38tJunyVlOVdFxqymBMhOs5Ico9IN5ANgAzuO0r8SbpWAxeP49b9KUI
2GutN1g8Nskjsfh0IITH1h9uxhhqUFXM8TmwgpwwtYblklanN4rBIkdsvgSHf2XzRhuwdt29NDuc
e0Ol4bS9BLH7n0eG9dHV1LUEekK8HuW+jLsat0/OJhNtzC4gw213pu/L8zjVRtQV7mOua40sI5z/
OgUVjbIkte1ya6BBjVCqPH2+7WkmaOA6OzlGPfBsOHkSHsWKfoQ9vFeGbHl9oMjVTKeRtJ+XcFCt
l95GIMcAMaahwgUxfmtiydKSea0KP6Q3f7T2XVNCoyTcDDYzXha+zq3XKDv5TjYei2EgJ/3ihuzU
3R1OM/LWe0NvfMN0bUAGya11FCCajOmSvh32tux/mBuFnQytpTANzRJjXPlMmhjo9BA6vn1Ow7h3
5M/xncZ5jhjtwvlpqENBt7YaHSSMj+d0eEduZDa07SbL753R1rst7QpbRWTeVniDmnDSPsA6BqaV
S2+OHTrRPbPy0p6EkWDn9HI0tTEekrsw3d2fM5WtLi9rCgkPgZrsi6DJMBQgQNb7PLTCfD1MhFK7
0LJbbY3NnkH/VDbt5BH9ZMEIkPiWTGSCl9AllT51Tst56VTwCshNn+iGpgEsTr3aBFFyo+F+F26l
pamGLQ30uJi/YMaL21SANG64jDNESfr6wsJPtPyXYkSXyrQtFjWl3H4wlUger33QefX8JhkWFH37
4KJUIDU4VQIsL1H5xIwZLJ7ch1TNo3U6lzh2JigSGOHAWo4Ly809DyM02Bt30c7qRG6WGpHMkmw2
UQ6twDfVbcTOGxMqoubI8O2fMK+Z+xiNfUb38xCDY68wcVdcbbD8hQjk96esndRtpYTrq10FtkAD
KZbV1BeJZqW5HJpktcuwvP9kIR+2j0A06OL8Ao5rf4CmKcWXX1abcuHONEa4VCSi+8dUMGuQvMrd
PhHRYt7rmGC+2Hn1uR5dg8wZew+l+qdWBboVAujAgWJawgmoCCjR+AiKxrURj7IWdXMznhK9SEYi
d1f0SzI3JaJ9unXYT/Rs3LDy2KfRb5gy2SUsoeMfDfAazDKyWiiYdV3DdMRyVufLIbieUekKK69E
3U1W/Ycm6pnxnXSWZWoWU8x2ZNvq/aUYnSjvjbHeIptChPsA9q3iLORx4JoX89wQAAU+xlXvomV9
ySy1eRjaLlXuzZJQCbKnGCzaEeM6YKuoTyS/InspRBPiiCa/gAdv675ao/cFilwePt9EtOkuioLF
neGQFDG04bfoB4uJIRfC9szPSrXS1ZX3UaYvnT+GAiCXgfdw9c6BJsHIgqFaoz/kqQccl0Vg+VmV
CXcpd4DNFu0PQkXq0lAv6IB5/qJIRkeK00fKI6TT3MLFkadrJPJNBzEkqf5WQ0y+3qL5JF4817wC
VGqS/wpPab7URoEyGcLYNT7GEnciQufgn3q+Pci4H9TlprlclupjQc47UcAk2+N9SavCLst8ccxY
gqSn7wN7SV4tzwtbpSi9AV7zBZsUQoZcaNzNUBKTgWZfs+Yyg0jRxiJBB+wigqpUrGq6DxhOUn1K
vxOeuivvtaIUw9GhFNe3/1TTHpWPols5+wByRTEK7Zoibcv4GJjAvJafjCeDIxFzG9/VnAGdwZ12
QrpqcFERlR1IYAo7Vq9uMIl5ZYazjBb8AKSyEFzdAZLx89ZC+h1zC9cWhXnoF9rckyAUfP1QExBa
fzasxZR8mNW6PLut3/iGSLOMYE0aoIxyiNhxxSGz5m6fJI/v6cDjvafXlrKoG2T5OoyCcgIe++l3
n2N/i4Rgo3JVUCdzif/5Qnd1qrx69j2XlTn3479kRQd5rBt1XibEg9o3zEsNJyW4MF5COfwkMbEB
tnwr5TXCvVtZlWmUN4peiSh8gX9BNAijIRV+3Qm9n5NoudEf6qmB97t9L+Asa1cp/Y6PjdGqR5JX
HTE+0DwkP7zy3wgQ6X8tfHBwN1Uw386M87jpuZ6RIOZ07rT1bi/n5LSGjgHWdZ0DA1wpYRknuqRn
XMgi2MhjN/eQ1jtapXBcg75xPuebHGkivJe9CIFoiNNxP9cGOaEWiRecsokcKISeZ/TX/ExYjuUE
6KNa3DHGxcdWTHtb7GFPlqfvLL8hTcDFlWl0Sb/8anPTiOJBzxLo+v0U22/RqtZbJTKfYrJg7t+P
t60gl6OibYs2rp/S9OR5AO1GRmQAwpGB9xZ8pBHNlQc4hTBCKPTarffz2Io9x3GY4KJCoDZegnjt
8jgfsEcIGzfunIdbPSOw6d4OBUS3c9kBtXvfdtR2ZWe1GuKtJCl8OIT6/7Cfg7I9jDS4yYn/57fH
Z5k7hmbp19NgMi3ytKNtKhWt4adwhL+ptLH33Vb2tL/X+idngU6j3HAmHP3qT2l5mEp3lDcZgNwf
kuTrwP7DVIcfPz5fwlyNPwLxWFwOW9kKlOWtLb8e2Lop/DGRYRDpZpK8rVrJ5zKkp6SyyS+P+6Ef
WWO4VTbOOYbLqYFsKtHeBRwiNemssL+iRpZ+ny2sPEQCA1CtlBrzKDxeQ4DmojHrysGMn1Xi4vco
NKLNqOFU7FuuRL+KH8JVFM3/VYiGr74IqbMOVgnbOCWDhiK+BK1LiED4yYIwkiNl3w1bNwRpdwLn
DgcmtBmrr/dYIV+3liRYIsdBsyUvMNkAugSm9Sz+lzc38+F4Z+hivwfJRXF3oJy31YuegaFo4uJt
Y2KJpRLPaE+FLqAplpsXj8FtiVKpaxmCgoEUaBUp2Kio91o/xpZ32vNIF7eV/JbANObjaL1DZeWe
pqtb+4QSCS2DGRHbeAmbVujNGuUklOHYIi639Fj75II+/4Nw8X7IGg4Iic+e2/QkteHmSTpE1dhb
FBbgptlsgazBHkYJ5OUbjLps+fHs7oejvMy5Ztntt7tdLk+mP+aFh72iXCgyDHfjr7QTOkbzLLd7
xOSPybZS2zGxVeYQmCn7IiJeMu4fbf9ShAV+j6bH9IuTEjFYGgVzFgwvS69aJSEjNi+jWQCcsO1V
6rMzKh66WVjNlzqVbAjS4x6UrfdpCRnX/4gEKrCyEPGuN4g8vE+5MB9bjXIYgJEJ6NuytZ7ym4AP
UkswCGOtLrddniNExwDq7xi9WnhZt7Ln+d/cME7gHYej7xKC5zsN8/vuEyXiVJseMxWbQN4PPff/
N5HluONItR+yvK0UE9osLrAefEj7UM/VcHLGV3QsXvQUUkgDtHGtACqNaW83P23Hj9PYTptcDERE
k0RZsd45w/SlLDrJSIOKxeHNK+NmZPBIt/IkaVuvkkexHBKiVYofALCe148ssx13m0m063o6nfiw
GUgFhHxQsHk+vk9Afuibgeq6LXjb1v/2Wydni8yL0g3aEOrZSNby12RMLUYywQbkF9ZJgxSOcT8w
4GzulSrP83vO5lUzbUsw4EUMOco5gWzcKs5WkMeaAxLz09r1hSJE+Og81wIX2LUgbQDYfmgiXzWm
hpmcGdOGdCeIjMnmpATR9asbAGt4ATnCmvw4D5i+zsC5j9frC5bhIG7EaB2/8b0+Q1olK38pMcPP
i87X2wPoLxPXrU3as3oCNuTIo3YS4IDDXk6R5RbSiquEIxMnYB7KJyNq3uXuHz4lCqqsS5g5XDQz
U8Igy9cNSOUmAhdNReEYa8vXeDHSYH/DruWq+j8PeWmMSKAOjHmveC0ZR0vwZwjgyW55zs6LRy8d
Kg3VhXarx6HGo1r2Fzh7K/XpqFVLyM0Ykb08pwfIH3riW/3duJchngOABdWeecJVdNbGqfkLRHFE
SJ6rcY35oFPMmqfSZSElkOk7Q70hzwrCkrMlv6oD5Zpwi08Q5NnFlIQoaFh3QTDIqfCm1NPSDVjX
UnP0HLuic9GNl2x+JMPSxGlkaXhDZX9bVgt4EDTeZxsrtv/ol+e8R7T4oxABfN6uSTN6a51x/hc1
6R8ua/v6ErHPSR59124G+03f2iYinuNq45zfmct3pIao/DydqTJnu1B4L3qhHCZvqCnDf/Pd7iiV
4j27niKnF/wqZv2yYKot35TvYJmMX8Ga6bXd8wKscON5zdylV8Kv84raJa5ZxJD0+711dYwcWXWJ
eOZnn87DyYSyfesWSAunuIzYbD5Pf9bFLy7DAsl59xao7M0t4LssmGMGb6hHOudFQO00gH9SbXqP
Znw2KzNI5U4VANBGyq3oKgsvGUmGwVJ9DRuq4uQmgAxTMhxVuqqdSOZJrmOmO4E3HDQ2j72uRZn8
T6a5mo2LMaab+gQL5QfDW+9FOdzt+EcKQfSdUtI9E0OLnTLRBS2bmwNMv8MJNN7C8yjv1fuqlCDN
orEHThnjJJ1ISUESYTwRnmDSnCKqcWH+Nw64tEZFGkKIGghKaM42lDXV0PkQ8LjWrD+rXL2J/J9y
g7Ik/gYUHnQ/nNuVCs6hMVq4A4f1cNpselmnI3zaCdYs24CVobHdJohx3jfLQjF0uYG4K2SRRc4J
4bgy+ldXJg7GlATt8gw+6dmZP6ABEfbr6I5yfHQM8GdKxwBbVqfWvuEHpwEl//wfQdLSiX1WE51H
DGpN3a9mE4zyTkdfvoOlJE5zLlgDJdHPArHLh74ov3PKnRZedUqBbsxVMyIxnhrP3GxJqjKQx1qa
kYzOgzn7WFjUtUrMO/ByBJ094TzPXCWg0OGEWI5PDJa8iHCc87+7BTEoPtaVDwNY/1hapHpOFbUw
12zTR7cU+Bd7lali7zYkWR73h8qvI50HGA43OGFkc+8ZNTDza/dMzaePeLB8PYXJqY4smTTnqQMO
YWba9kRJ/8OoiZ0K7Bkm9yLzhMGqizu2yGQzggnv5e9umNt+cR0DJ87DNM1c8X059yke15mOFEo/
Qa3Zt3yFErlceCQ3jHP+JuwrzsvP7Cb2Nrmi1EjbA7dwu6C0TDLBy7BO6bvsnSU+f6UVvxwSSJ+U
rdssPeppqwO7Ew5/aLYkwtSCcvqELZAeeuajkVOR7qKra03PIfVnIdCg/FYXn33+AAKJzVq1zd7G
2DVh2Klz0zkSFHY9BAYxT+OPRCLlakUcaJYzzw0MMrXGbOQOJtZXenlJedZfBk7Ky6MuUPNI7Uh7
E+z1f/VKv295UATaSx3Pp6KywNKIEskzvWnvyeqoYj3g/gb9MUSLJ94hSweCquzNNGgBd57z4+da
2lzxUbZxgNXa/ZsVqZ58G91Lypv+Bg6PTXGuSFnMF884elYLBesx3vS98JeIyKqWtDebmifXZzrn
2wrXAjpAq15XVse/QYIV8zG6CCx4lYRvXnHPAAhstk55VzTqVOtO3Ey519wLNBAH24bw599olRQH
/H3InHjdRDF1W3ZEqgaLKMjlu8pyv26w43jiX3SQLeVY+oExSYPyuZjRGhmiONJ0v9hGcd1wgi6+
0nOcIUkjQj2Y2CHSJo1YI2uCyogHn4jszovy1i6GXhzzMmk/xFfv6drQHB3nt9ZCmu4nlHkl4uWj
+dl8qCo37WuUdM2Om/XnnqDIy8rfFifUzYkjrHvCjpY9OnQPLCVfVYtKpQim/AjjN1cfo8CkyqZv
WRd87F3Cak7k4yHZ64PVhQhxoLI+gZp4Oe746a5An6iQOl6J2yqsihdW5DG+qLSo/Y1UbX2ljQpK
nwevniEYhPh6/WAfGMGKifUVOM73YS5mDxR/uFXmJBcHVTrIQEc3GBmOIY0IWZuJLjRsFjGQcTS+
QIuBrDTlawR+xHtMw/zN1Ra2erlGmc0rAkgxDkKZHVKJIhM+9DgQ923LoT04VPF7yxFQ7FTXviqD
KpJr9NemYklLFTcLH5FmzlU2D4LvOGI15gHwjm9RxnwAjExiU3z+hYkMEXifCAhUiRDpHQ8Qn8Zw
Jkt02MUH98NX13WomEWAeslW5UEWcpGf9iukz182Za1utfbKS0Ebn/R1YobnE4ICFfhUnLtBPuL0
6RSkMfDhE9HSi8+sqcyyfq72rmQGB0ln8GM+392MfYFDr+1q1UVYtU18L+kscw3Y6Q2ruPLDd7IC
+Mp3lxwVSYthS19i4QX1lTvxfxNM2hEO9mE45lD4xPYf4f6FPSDfSEMCID6sXXPpvlsE70YNncfb
GHT/90uTlC3YTtGa4/NRWECk7fAkwEPygOifRmMaZS2OWAF2i0gTeOcd6DruVzDblaEK0TsNrVox
aT9iVH9HIcjzdyJnY9/LAC38o8/gPzTiw8ZV3EuvfGHvGermiyVJZHyXv1LCZrfuv1BXTrq6uHMp
nppoCEOJq3HZmWsHKv5xmJOAA0KH1Vb0cdZ/O+/rkDI0b/GgHkfrStukciiRcsN9mzpwb5TXTz1h
gt2vfgLg0sFJOvmARhO48jDyVfLyxqkwc34wFfTjmugONuG6hluZbW2+K0rUORl5QKUUBMx0Kyjg
QQmJWIXAP6b6Z0bC2j8uN0JKY4waDeoCs64QBqhNyp0dVTF5RWdHQqY4XiuieW9llrPj+OBBvYwj
kDbmyhwJjgjTT9aUe+aN2vZO5XU93jUv8BtehBw5E1Y7WGqO1cv/aAhNQdOaetj2nILmke+xZQbD
ftUrWlKj0If905Yiedx3M1N8W7oWQVWdql3tIvcYVzQaxWd5HLR1gTpuw1zTadc2RkwGCvlN50UU
M/uGqLkok0gLKbecrPqUAXO45vlC0F1A+ukPYEZGUHyL80B7q9WT9q54WbhoqAfBdJKAE6aggrJN
JVSSNaVvOHL/SqNKkfC4LGFrh3AbfPEcxAlFpx9Jo1D0zjhLPoNGUxufm7SJ8YCg69xX1mlONIN7
SD8BhdlNVl9hVopg9dK3L3TdISyZOs6/VpyXTi3OsKQCQZcHCzLZx80ru45eYLCeORgNtsO0mDy4
/EakU7mNDJWzPwm1bKK8B7y7BSUwz87dRf6Gvy1VMO2Q+RNfH7N2oCX0urOfIKWojCHU/FiZXs0d
lx61EG2X2DEaBw3FNx6l4QJg7eFciuZ8uJM1/PCkPf2nvQMmwhfRnUxVHACzUG0mpl6heVppKvAH
HDsLmL/65GapxhAUd1uSNDE2nfKjYXJuMXSvr1Uu9N/f/SAKYTIH8PmqSFJroIQvwKRip+h7YUWh
bwA4TkmHxTmcq25A5fezi3KL7+NHLMIfmVMGHxHCGXzaIxcSYfjRLLfAMwGSPTohpOUWN3QlrPG6
235LPEl4CC/zXUi6pgVxQKXFfsunUaVLIaW5R1fQw1vYVbQPqi6tzt8U8dfs0hygLiHbfWcz9yQO
34EJePC6kL7M1MCigQd7usZxHbjM9fXXf90E/w2JCNTUhYVW75QrGJGyrVkxEfA0eCzetUozT16r
IBKER+RuLDd6vP9zOKxnDJojjeNlvjVCCmYDXwhoGRvI5nFBdJKbrE/uuRKFP9yLihLJsQI7f7G4
qV2iI4VBzg0yQfLVIBUiOlZgJHgKxfp9CAlc7O6bAq9+feD499ooPXMp+58T3hn14paRqJHTHm6Z
PkVnN3ehEXtDCAFEVLcMZ7b7amJVSuI65JSY0U8W8nidTHq4jafJrXQVZ1dB+oLCZd0Dj7igUNvM
FfLyGcnPHi+xvCrG2/Vmh5ybmJTsr1yYvAbY9jb9a6x+6FCHtlWvxsqc/iTCGS4Xa+BoxYSjFwZ8
KAmtlzJ8UMiRHNSfIQNRywwrO9Cp3xxXj+9SRKFOYz48OeXTa3paux2eAQ/DmO1ucmZxOT88Rgac
ovfYbSRXbLG9UFIM+c+iH/jU3CGt3ul641JESa09MFx8fWQXu6k6gd3Eto9YIvQb4phcjBqmZ9aS
FGrtLg27LpwbFYldfld3mQnrmtwwIIwo9GUMn5bfusi5eAWkzos2Ip0sVE3Qs8UMck16CxVemX82
Arz3iyIZyR+VFEEQQv73ljwT6c9TdbKz3L9Df+B0NShoIs3yE4qA5Ed9uC/6jPk5Cm7fVPnC4sDV
vCFyF5VHFbrWcOvKXv/u/iuxviWsRZ6wPaN6JPZov6jaS+qAKJZZlMcw+TYH5hHgh0NbFUPcoW+S
n9ohGAvsHqpmUeVakPmwVQflICi+Q4CwdUrflU8vQ4/4GgyoeHdl5Tx569wVMdrcs0bE3Ua5wfAP
p3Q7glehqVHKQeRERMa+ci1ublkCveMa27LghGB0Yx5gJa/5SSO2AU+7UMKksfr3O6I5njA3/Y7K
E8U6P2kV2thd8R3wq5C8t7TizFhH4u2M3G6HvRvvQpo9GZeJL1rzfUa5zgJO4L3sIrTK6Cx0r6w1
JaQjonbyPvCPSz7LYXtfo8heKQMiUoCm1Hk8RCAvHcRBGT+/tJuwNfDb7eh+YnKyg09ts6raeyRN
z/9IHYSDZlFLt25lxxPIWjHQHqhLD5AIqXf0SBAiMlk5WQOyOl+X2Aa84eov3TI6MPZEykKYE97Q
mbFvwei6MRI3inUc5GFkIUCz70bhUAlti4jgXi92jmNCj2kjj2qipLdetyonyGAZ7QjFJd/2qBxh
oNWiKgiRkCdudIc4+4RCwJkJ5ZCbr0W+otYrWu0VAHJS3e/gUdooQj7ghOoHqqBJpOe/8QZXaq/+
29RK76q00uGs96pDko0SYAmvwgur3x1sSYeLZz2ZD+2N2i5qpRlL7AEk2qXxZBbijCaUFXOJuoiY
FY9YZhkHEixl+3ogyb8Dpr3fo7YQKz9UuSAOc8vmz+S4/V8B9L/Dm+KVKhuWMa0Onm9c2SKK3VWv
QjV5isNEwkwRqBDgtl/xUICxew+yyhk3Q3wqxlpRguy4W3BlzroxLNJDrnBROK2fLez7Yk5V+nhF
qvZTf8iQ91PiAvDQPdx1ekqhKf4rI1jdAzSKlbwkCmq6wRi5eDsU1gZYDTaz8uO2dCdkFww1xGTA
WTLvTq0fVMBHsZtkl0hLO4L4/7gReDPVutu/0cZ/TJwv9014sFTk4lM6E9rKDW2o42/082N1WIyw
USsqm27j40cEJcIRRT9PwtFd8gvnXbtdF11/z4sG5Mb3zaMAJfi1SKXfg+yoNsD5LIcbyonfUPyk
4GMjBUKwvMYK9w9XOZnb9EnvVaZTKsW3XO2r63L2XSIT/LuN1Pcxlr885UUsPns5x+bZmN1VfIt3
R5LLTw5yCrZdh92gaAEAIRvRQN8Rdx950OZNy/WxBIIw8BGSv+aCoj+exMDE6DMj2WGxGkA6UJ6T
BZ3OlT5X1k6uRs8tX5H+KxCkC1fRYvQWwM7s/0TvrVVfBjBWrtdQuqwYi+TQC4TlLKBaL5S9qlIm
7HtZXIBXLKNzuK8HezJHxf8Li+UQ/7EbooiYVpo6DEsfrM4UL2Mac0vNDBtJAOsbt33ScORxq3vJ
GwXDT9g+9GWQJctoduSLoctvcaUQE0YVYCqY643eoPLEkLQSO/4xLK3Q1MJRZV9ljWy1foxVbg+J
kxGSiKa13yyLGkCt2B/FJqNpye/oxkB+lldpJQITo3Kfoc2ONPNLsLo8r+/WpdCPBkuwDBr4kbDi
N+J6ZOEbS5WMZASFw6Nj84en2pHDX80l6nN5nR8zp6HjHi64JImuI+TrP5UCgefaSX04ZQ8TOsnB
9fLQzvprGXKKQvZZk/oMWdAnxWgbg5ZVSdqft98Dm4Xwq15g8p7A0TOudrr6rpI1hQGGDHXyTj7L
T6W4nv39VOHzs9LbjYItErygBl/De26WAczJSakFFsbumDZEtJ3mMyNjKtz4UK05AaXRmLbKwTJR
+xXEZADV4D3fuiao5608f+viKEttXeF0WpDClEeciUU1q1SR4EOBAsrkFAfI89UuMjQw9ORTVLvq
G+I8+naexRiUbXl0IptOvFjM77xseJpodS+yMACR6Z3atXjmZ8hqj56X0aC9R9Txns84BIEWvD/0
XxcadXnQP5VqXHQBRn+VFeQMVO4XaKkbfap7ayCvddm7XRlgiuZK6l58grQ9D0OEytu/LoDggzEA
zETMNcm53OlyZ5IIRmgZZk3ERXwQkvSWophB4mAlEayFwc9wKL2mieAsUk0bc9wZool5W/M+TV4P
ZoR+L8ZJ0xfWM6S2K/he8C03GP8ZbCwwF0K5Ckc7tU7/xHDzwk3uv2RztSO0pw3SD+TR/zDIy2db
tQ/s08gHhjyHjKdGepZM980mHaKJAenNt9WQo8Sw0p3zaajSZnIYZQ8NgjtbfJehgytSH9m2/zrX
cufyrPVq0jRFpNmfeMms/RQ1ZSLSqEWJOnDzvqiADotCxrx5mCP6jQmfk6pgVgGnlFE5tkQQe0wZ
hRnj0DRjGg6bCyXthHBp8yYzQNYKQjKGdJPbtAebZcB7lCgLldIiVyDCfqR0gYZwqhuVLXe4Qdwu
lRgg3C6gn7pSkzX9SXdyWxAajR6PyzQV5z6oT4JXIxHt/fl3oKEDG+rKUwCB07Vc4fU2D435VNTg
k8SpxwxWzRR5UZ45eXxnp+WO1sE12GRX8x6ztA6izF0/N+lgqjFldGG1tx5AIwfGuBQQ7m+5kpDC
skSS87GjeKZGG850TIm6SjIl+Ham7hmEQVe1jAWo0Q/NYUrG9hhIJfSR2wL65TeR3PpbTUg/w07P
VnNTIQ44eQxPOttrfpj9kO2HFWyJCoEV1oih/E0sm08T0kI/KsCXCA3om+8zVsX8s2p92b/B9PKb
b8CaqSPhXrsVo0NVeHaB7mBHrd0G4PFkqVlpe5UI+kL8+3Lb5tc05cvoPF3Oh/6jjukNJgWm7qUJ
QKjWonNm9RKnSI3bMQIjSKrIpx46SNzqkzq6a+gfPtFIQFpVLpiYKF+ytIviD5c/uq8Jkx6qBkkI
kKVmM8PJXQkfAF1aYq9WcXeYZMEFkyX0OWoJ/jfc+c4zrIT73ZBQowEXiIJC4H3OFgL/T0ekxzYR
aW7TSdqwv/EmRVM4ROpCqcrV3sX5pykwZv1OrOIio51qXLazQEJa8yFYqTFyeUWA+SxoJEn1c1Gn
7wCgvDGqyNFbM0PpKPlG3NTS+pgaXwTn3cdYLqNXNFBro2XVvsVPDkbKx083hB2cF5gr94QV2cL3
e1eO92XiX3Kj8uTsdNoqoz1UHcd9nyjYD/22Kk7wx4a66m6sGJXdJ8tJeFzontUrV6EC42B4pnLt
rtVQ36YLCRVE7wCTAQYIGewMKxCUKHNrA8mSiC2v9zH7IwGD6uu4b5Tta/4SdrCJbOzFFDtHEpzf
xley30HVS3W4gK9PtONXmNDgx0zHh+hOfuPYVcuXIGKkowk9NIMqQ5Bm182JseV0DQrAFbflbyK9
idpyrgXCmLpVDDODCCrD4pfw7ens5dK2VNXi5oAK1O+mEvxDn3gXvGqYhYZvrPUb6GSCf+6c5jkp
qJ3GybS1W+9KxAfsnyT5/lTHs552Gx4g8QETZ1Oi+BEq/TlnO8k4HONnURF+bw4geDkZBREf2VDp
O1i3f84jZ9m0ph7uIC/jsQZE1yuOSiR+t7k+5zXqcQnanQaIdCqyEwP69WX1GXl09MmEddifN0sB
V76S8RDcnvBPwb9Q9U1+gAgGJgsyLegY+HpBVL34C9EH29FM0cBLX84yQJVtNCrwq+FV/Udt86HU
HgqHKxipBEYWWK7o6VIz4LBfT3czecr8w5dCv3qqGu/UNyJWGkvCm7y8THBUbGGIS23sdSTvAiH7
Gj2yqdW75ingZQsrZWrnu8n5TI5pZ+rrfOLrRPX+bachbAKs5YmQB/X/CbKCWGC+Rdi8RNuq+rR8
r8UeBruPIlW1+NSIQrI9zdTFqCo8lGQKymAGXDIa1RhUGK4OPdthut70DDQfz/bfZvMDj35lgY6N
oTBtSjldOHjHOY758fG+TaIrr1gHcmtF6r1RgAoCxAKI4VN3wfcCOX77Y1sQwgh/tz0Wc4SqwAPB
nBT+XkGxYtt28igRYPckl2vYxEsNTH6ZGBLbNGPdS4a6gKuQxJ60dQYy+pGBaqIhDeA8krvCmHJf
5w6f/lR4ozTaVr6M8g720sMZeXOiM9uUZGi3YbtbTYHgOXqacWfAR8eVH3MEqFJ3PZQBOPHQx9Rd
cRG9l1qRyQfOhnSf1yf6FLH8dPkFwdmCD84974xCIZfrOe2Q1D9Jy3vJcVG/PV5lnrf5pUWz1kAS
KIKwCF5o2xjGqDuFa4oHV8L0qOVtchFH1uekdYfGkAUFWM9CcL3dAJ+EOk5x+ONxBFqit2uM9R9V
ua4utPQZqby7N7YafoUEUckCxwR+FoKQkFvPGc6er+ChpsSUtCrJygs83BIzboOgeFdKSlv1jeBC
/7JngbPftXl66+nn4rkndrLxunImOQzcz9uxbHBI+vFSd5ZdOCP6STa8YSURsYeMbSFhRcwdVfkc
mJSUH+mHx1XgbntTOV67gzVSFEcBmcZfUYmmkzLi584H6AbpUaQhtoAC6seHnWb9e63hmBOeGtGu
R6svtr6EpqK2A4GSDiVQty7eHQmwswsLEJsQ9qlPd5FQ6YkndRlE94bM+UorpxavsvvHNgsOhkIC
QrcJxaYEkHOYvCNA3n0YXFd54HLAMu49cBv8x/jf8nhBXa+n3h0/OHDfnF5xXIRd9yXxwxuSK4R0
G7aAA/JJc6RxqOGUhVRKDJhFsntqOI4ITR4swr/rc44CrR79fEVQi59yxe4uwsuCWXpDShgm1/AX
WmkiPIS0XLKqb5GCoiCC3hB8row1ILaL2hsxT89T1dVU+5Y4uuRS8yvO2UvzvlBmUG2UJ7otaIoj
c8HRuanBatCm4Cefb7zoD0OJ99dCEW4G9ac+fFHB3O7aWHC3U6Bec+7yF8X9xObOIQR3zqdzsz5n
u8lUI0TNcZmnbjZajie+jJ05dUOqAmMaYk/TSFJbxcjECp5FqyUJLt9CjmhgRDOLHG+xb38CdHyS
JfzRgaAHv0qj2ofAGWZ9oU8U82DcOu/fCbqOu7Al4t+jKd5cheTpRpKEgHF7yb0vcMWnCcCXT7AR
cl4eqPwJkJx8Bi9qZJPCEZ0DrNEGU0Due+cZUJNJWCuguOFRIAawlQMUzHwbMUqtMoa3ozcmpBJa
6FfGLQJr2VVfFlBW85/wUlRAdHmjKmyS/lbsLBsaOib+rBme6OLzksEDdd6dgGMdjcJMp2FoIMC9
87h2fZu/2Rw4BfD606wqaXdSLvIsJE37rq1UHfthpTVkS11YMPE88iPJ4e7Osc8+EWnaoOfBMhP5
OzUtTRH5aEARG2jP1skj3/ou0/j06Q87lE2NmSKMEAuHu53cCd7Zin3PWAs7XS8XoaUcYcbwjrb+
OoYRjIKPVEpGYnJ53uikqjqiTXiu9ErPRJ9GJyATxKpIZngY7bIhEwAVk2FwUov4O2oCWFwTs7xS
7JDVBPvcxWZ1IRtIjVvhXKnevBxQ5rtACLVkisCrOUcQZ3h5BFfGP3gEm2aZd7TboIBv5XUTsOE9
6XPQr9V7yfqjUtTZGTv/1WNz8qcHdqaJgKCWBkYs6plp0WPfhrSJ6zCKL7ie8IUcLkYhGxqslx3I
R89tKxsXpgQNOQln3B4FNaHD2vDSMmEhdhQ9YvU/bc+tndFbNjyeQ7CpCPxRHaZJy4e9TC7nT7z+
whlW08ki9SwhM+bJ42YROrYJ4DOGEefw3h+LdkUvRIunbqeyuJ+aW6yRRwFnNlo62fCEJ2aUevrl
bMQYCRFkzmOd7xGymKfcDyYtXTXW1y35cbBkKwHNMFo1Bosn1PVh9Dgzf3ODr21UTzRbcIoZmACe
XiKX5dTZTrqW6XXdomHTAKcpcFSuY5eT4KVYr3XgUqFjScePERTu+VxPKShZ26HQJElA5gKgRZAS
kustaKNyTrMiSYSRe3XRrXCgDGRWNJA/3mHPjZur4oVdD9crfqlD1y71xt3KVih7kN0BPZbpfJHj
JxSCeYRvfwBxuuBNVa43B2yYRz9r4L44wOxAshfcNizInbVFJ/ievIE1o423+mjLaEhZ1U8Hx4l5
apcz2VK2iffgu14/tQMQosKlTXmYpI4nKmF1tt9D74LKZHTbQTn8X/1l+fd8ms0phykQhbTOANhU
7cv2vtmEvfb+9DIfrFnNhPO4uBbDsQgemBjWUmm3uNCAUIDs1G5fKBDpLb7FL6YV7KPATX4v/r9t
sJUJ8UilaSaucCo67S3lc3E7PNmkWxO/AUUkxPqs2aX+F+cIB/52p77hR1OsAOoBZlwYp647ZVsW
zqXk1x0SWKviZCQ1df35FKk18S4vWvd9om57vDvfc2IFAFbpiDy5Nqne7BOvxmgAxtnsKlKMJLXq
XsLeB+c8hyKHL0UXqBAqsU2oSEd+Q1gqr2QQhc3PSv+v52uEka3gvrEKvX6WIw90T/JMDp/kHWc/
isP2OM8DdjFfYZjZwUblqFgU1Vxp1vwAl4FqPOpCfiKn0F++3p3tNpoUo+MgYvCeOx//p6nZK7fw
ubijwD56BqCGDXeHWCfF2YV2ON/1+0qPzyBEhufKPkE/dh0gB4jG1OKXvj5XL9sVs6yKQ2KUDNqt
9ixA/KEa0xcGQVTUsJAEJJaa3TuoahKhmDOZGvfbA0Xn2wcEx7SO8PsfQ+zU2+Jac+vPpjOFb0xu
k1DXxA3chzjBO8HYSS0lJSkxww8sQAlisP63gz9fCNzMkW1+g0ulFQ5l0ZEiKq5M6axRC47s7NH4
RpkqX4H84cc8kMysFjlAN0Hr75rYhbovxA+nW9If8CqQK4f0LoHKxuRwk+T1SbDRqVNuNYn+42vB
HtvF0MWBZMFvADNA5c733XlvOy75LUDxsEYElzN72L5Vh3wFPHl68SzjV0CpEwwOwPtUmu82encG
p9e3Divw6lt+MNiOhwekc+ybDWqRsTR1bkB73WrXRFghE+1gDxxjIH5h14ezskvL5K/rpUhecShR
NXZnP7Q7ADisqCWWxLdDAxcP28emfQaIZPsBOsCji5CsB+Dbk8obtkmHZSfms84mkj+3OXru5C0o
FWOMAf6vMQmm+n4sitSiEIXCxjeoZpWhH08yokivRpQzkUmbF60ATikJtOsHmPxYxTNDcd7y+Tlk
a52m6DCEzruBuPBraIA9Hg59VNSxvGlU4m6bII7cSjBtJiCp2grlMxvtuzYOJIrHRu75qVPoFaS7
d6IImATSDfRU6dOFtOnzRhfIDb7P2c/uyYu7oqFrc9b7qKtYNxPwREZwUVKPV894LBL4+Xd2bL1v
82+iB3rST03IYANCJibyNA3iDZQKKY1lEt/uah0YUYlMln21D19sIE1DOMrQFrjRBfz+6uYbVEli
1gPiQ3sRPZBXP+RRo6rv+1/pzrCirlncez0+BV7m55tUqzlkFHeJtqW8wEVbl31nMoNBXqQl0LPr
ilp/KW3jEUUg0cXKRuRT20R8sX6MJJM7WXzpF2bJ6i8MP3CqMoWXvn/jFJiT/FzCHI9V6FOBbvi+
jP2fjFmhkTbCiPZ5QCIt3jt10GW9Wcy5uM1+MRBdH5aevVgvgF8uMKpBZMZjAdEA5vDG4tzTpt/5
nIbKjq6D/4D87MwxaymMjyljku7nzsDN4nQgG0o5r/zKPgWcdGgOCh2ynkDS2UwwLiTTBLDfN0k8
fFJ7v1oPUVwusoxW4VlM3JoKDaWCKwALZAR5c014ZRjH9+x+2VYPVj0lm/IQ3CBkWoXpVrjRMrQ3
2TkTMFgcw4WoQjum5F1PTrDuauGHm4PNbP+gr/aCZC9diHvqQooRpbSxOoAwpuujLDG1PcDLLsJd
vjQSeEtoDRqa10SGRy1PROCnGYD+UwSv19jQpIQgP0a54OXDCJLbd9tLntHklHnT3LvVQACG8PuQ
Rj3RfqmmwM2GZFZLwL7faZhGvNXmScT7kN8YH4x/ZTGfYsWWJJjiLZv+gHjDucC7qezA647p0sxs
wCB082CE20WVwtMHJFM5DSWCnQomNiMgFxNQtRzup8AVzLhtmZMrsYJ3/pxi02PjjRKfVK6+uVwq
SSszjatGUzyhNmolQnki4ufxip5mDwU1Poun0nKyYTjSx6GKEJMef0/atCMLsIBqwaKH+Crf37iP
IW9lximBXPSvfKjdQMx0JliUrh/U80B0QBEjRlqWe6aJX2a4SUjLAD8s/kcO3q07uTUfGTYnELFq
QTFeE55OJd5P4OyBPLMcwTW2UWtuhYs6K2Ss8WuRlIM0iyK2CwNBiCvAQxJuw73wGy9Y8DaqL78q
Xy50FsgNzwIg8fbY47IJ2Ns2OKGkZ41XgMvPRwx+UANxr4LhHexNJfbU8n7aAxVf1y6HWqtQWPo1
20OmDwCrb0sabUPjv8/JrO8HJLuiZyJTZ7M50K+1MkCJS7XYBJGe066N4G54z889jnZDajyI+GJl
Hh+nJluhlP+95neWk+mgAJIfBWkWJGnCCOT4ZMny8yqOj8oVjCtpU+bleScjKhQXntxk2cwBhDVZ
8mI4Mq7vuId+Qt3s5s+5j9U1sQm1KQTz5GhsgSis/IRPFCFHRllpdHvkjMC9l9A5yVypEITDC++P
K5v/cdEeaaMXC6cD2PbmOykmLDjRMBL6ouqxCo5GWCF/SOgBt7vy5fqO1K9/PaDWQM7OWx4aWq4r
Wdb5sWEE7JMBvjQ3ay5bxfvA245jG9Jquk25xWg60SLehOqSY4YkzcmT+Ag363S7mOPYFPbPdQtJ
NbvkPv6b2ZYpd/pgrWUD0vPq682KZPjP/VivbAkD+h/FeC4RI4lnk2BeF39qbOhMtjs8DGEP/eyx
XeXaMG1KY1hjlE8wLXS9v7E6P9TJO9swqb3Em+eHqS2fpaX/gatZUivZiiCH+60/PRxNEHqipnMk
zy6ExeG6HQkkI1yNS/vDdpXSxiKkMw1Q6Pao4HZIi8T9blYDh7rPqXili5Ufsxo/1eSTWewUWxnG
INiH37sC+pT/nxDSDQPA105kW9MdHjLBf7qAJuDqMLlFbNjflAKSETC5YvRKdWiMg+CKf/BgnrG0
2RyOTYpy2VWxA7AMmncd+l8Y25W+7TzInEQBnkRBPNkI4veUjSXSxdvlVecxYoiOfw9sdZGTWVb6
cGbCY25K4QDwg9MNNng8r0RGEYHIQ/97vFzYRCMHShw4UDYU142zLVcJ8BOj3PodAbL2nkA62VI3
lxHtqXTad4RxTfFJwCx3vXGoydxyqG1c/0xSQk+pd+KdDPvhHKgewicHzbxBGuILbBABUx79wq1b
jSn/cCrQPHFoDeu+ZHtfo8lbZ1lEhXpAVtdVjv1kHtv+RJ7pBZx2OXIN6TwY4+XipyKWJlCitxZH
AICGS9x4pJRgQcoagQN7s+L4fTgsnfk2QG0FW4kbvVqQGvjCqMlbAGxMM87TugQ4SqxdVJDLKNc9
mNwefN09HszewlG4s+yKe3+S9knWNj/HnnP6vhZQG2r/tSY15YxqSVFt9er24OvG1W3THDyNR363
+hkdaH/sfE3s12pIh7g5dS7pkt3gY3R0CRL8e/qQ+/Le8MP/khZbsIvWqs3qHClQf/urOeTvLgur
MGocdLk79B0xanePam9waNN37v6u1drOeuFfzDc7akWLeUhVKmuQBUBPpmRBhqD1XuS2grr5SFHt
dzglv1Gmx4OJ2fiCDbTnZ1hUY/qi6/fybRPCA0Bd7IdnyYFcv2EynXzQ6+XPhbz3ty9mdlF0TMp7
fRR3QmnT+9POpfeiQfthGxPZA9L9Hez0nTq8of6qXyoJy3AU0odpjQca58pyXNwJb6LdAmJWcKbT
tpoPZoM8lLJNnBgMDuqqO7AyfALUKvjvsf6IeD7Nmv065lTmc4j7ruaqVb1bisYpKN21I/XOqC1A
NKMx0KGab0zBaIc0otSta6cvlED4tYxLcvnes73DpVYk7rL6dHcdYhNkQkFVprmd3p1UzeUouSvh
SVewABy45T2xtwos8bIEFXGbb+WFl0z0DP/7ZkNBPlM58/cQIDwYQparKI5AJQPDBPStLTMBa5Hr
pkfgR/mYDowXVDWwHnONJmXLBnC3gnsH3EWREnnrELT03hbZ7+isdWwPyCspw7CCAsUsCnnVU5ad
nSpfZJpZ8NyBXBdx0HCYnoOEaeyiq6KxtUe5kzChBUv772jpipOX5e6gRoTfAKf3SNgnM7ly/3uC
UdU/4rXpL+kJhGvmcxxwyRUfSqARlcoSOHkVW0ksS5i2Nad8/VYcxtdRvKAk4gicyTS5YxBXaSqw
hLPIUqU7iDXvR/kNKXksQvGBwTSoQ1XcA8QG/tWyofjsPQldzP4lMQ5ELe4V/NtY+bru2ZALjs5s
hIe2izkbZlvrwiIye5RACOhbiS9YIM885mGt7T+ECSTfxHcHOlUs4aiHDZdZllF8yOp0vGQowhFu
LtB0ye7VTTy/zR/502Xb5xtS2YShkS2P7BuLZpf8YiiSr2WoVJeTz9DQ6u+ZL2hZk4njH0VvHyD1
SyXfoUQeXS0XVzZU9w1qFDW57AEa4IRjjgyJL9+DInfPFWEJ/A+b39UT/HJm90wghw2MsH7igI8G
yYRRO1E+5012k+dG6XlZPxk6KwjgW/ZdTy2LX3kN7rTK1XmOoZSy/JIMJIV/WxD7Od2Vjj1EvhLZ
KvM9OdHq8Cd199ElOszQ2bm3nK4XL7hD029qshxOjFt76pLYqw9fmlCWAjDEegVL/i10xxRQvgNB
4/2H7gFO74chSSRe1sj9m57CuSjNzE2zzfwPF9Fav+rfKqiF8edQRZ8sr2m7uci9v7gWsZ0YY724
lShgmIhf7V0cgAe7WL7Ct3r7BHQzch5m5EYOuUcBxucnj+gu/34zHgzfok+ZQJysdd6IOcGJQk9b
azZ5zH3JNMpzBAAkDjD0Cr+Xl/998C5/QshMtPIhFfPOaZWBbZkmuJFI60Hn3QyPpU5e4beSKGzp
bXNzWmVYn98KDbXCLcl9Xspmib4KPkugMLoFxG97ISuE6K6lRlpwovzwr2Xv3UWLB45iNsrdbkG+
58Czb4BKFfD+W2kw3MU8F6395q4yvLihAtz/9fL1M4s4CQ89YOYCCErPQ/H+lsKfssS5HgGTJbJA
DFqpPN1uKSxZ1Q2G0pvasTqKaXDG8ddRl/IOaow/say/dYrg/itukHRqkpgNWnIdNsoV6MB+scto
lWgJvCUXPQg71Xugas5lpygxyyo12sEHP/Uh6jdmkvU0fXXqed8hkG5L2q9fwnV+b95rECFSbwO4
CJELPwzZITd32bubcgNwkrcZtt5/Hnod1ircRcYjpl/n0PH7D8Svu63kkj7wC791HYA186NebC2i
2Aush7JpkNk5iEm4Jtcx0iwOsBJA+pBNms97uOXsxMRz0AblECkBkDNGyaqwniupLugZiXQAUxly
FBv0l8/DaZFJg9tjqisT8IwqRt19XPNCa3krg7+Cu/oqUVaseCLGEK269CgGI+K5Oc74xUAaDFbq
ro9lLWtqrQNbnYAs0QtSmgsH3WwVpfh+s8xTIfg9lA0b9XFaVjq3dWcEfEiT6uJ7jEikM5Bc43si
R/J/Dr/MmLx7QXb3kcDN/g6rLVFfgzAsvbADHUx3ZwguqS5gTlcz0+g3YRFwM5Ax/zmrtQyQlNxZ
XBOB9kvlb4SX0DFCZFwjPqC2orlD9oCB3R9OZFtty2szWdyzCQ9ZOEIAQt+CPLd6bsK0eoEY3s4p
X/jA2246oN5dT66Uf2frn5M1Li+XvGKGKsm/VnitNfC/Y8KQFgOZcZXhaLoLEGx7rsVivF9Ng7A9
zLbS3yD18nqIu0nXsJhVaQwyKOiCS56ZGN1i13BTbYYw0ahqIfyyfzZh/pnOeVETUfawSW5G7bM5
Vn2xNAI29PcUmGlH7F8JXNMp7NYi7Ql7FoalZLZDPEL6YFroHT4PVJ4L6n6DnQotxF+fNN4/JwzC
I8PYE9PMwRlYeXEnbduVaUidluBQJYgfpGnb/axZIJildRMkG2wldIWE4FOTNMZN/sLLeS/8No7L
MWddOoi17A8leq/vXCzwXYAIkbADf9ySgDweh4fyzmmOYSUGc0THsWZ6Q5h2fGh6DTXR28HDVZp7
V2JuTpHR7Ux7i8vk153oenPeMJptRLimWlaeWysiDVxRO2uTHY0TaH0OI2VosjbDIsUYCEsW/43s
px/OsiPvmkMBjKgfWDuU3/lO9LPGv0bxXXu6siiDJmHRMtVDj7u/c4A7D2uC0afURPMd3Qrh3QSx
C2skDd1FhGZenkflM+0CCmmQBiqim3O+XMiHAZ3L5nkbpCooqppUpYcig61dkXsqXFq9iyo97NxD
nWjcJLMxynf94uc0eS8QKmTDQKsjsa6MR8/OoEzc61d9xbbGwpkeXu/1NsNsZ99ULCpJA/Apzf6L
R3MS905wG18sQqpK4DcKcR/tLhtuEmPwPBq/z1hw7/wsNj2RX5eHPlOhAiamymNXQ6M7q+nYzzhU
CM3jQtcye1LXg6R8d4SD2DcxL0/TU9CI+6aMVn6wc8bco9r0QLpnplvKqb15r7pAY9btErtp7ndN
dAwJrKpKUqtlkSlWSKS71M0f6AVL1ZxsQUGD2rzw/KFQ7/WGG6vI3XmvYQIEssduazGiMEtq/QGp
gMrf+E9b1V6JWb50ALVJ67wjL4f86M9TCH1ub189TYqbA/2x3qml2mFYZUFGeQIwyaF1derxyRi2
WXhD/pKyAS5vBZWzQJr5Y3YWIuP4siBOPOEzPOTAKKPMKVqfp7AOSlkJgWmZiGJZa1IxvV8na90Z
qOtrdNmV0iuDyTD3og8DIxypQb/7Hhb+KeoQ8KOo7iXpZEkUoVHGSwLKmIwF9H2xM9TEFTt06xIt
X+8hNQHPA1VvKc0Mts8x8sMT/usBJalIZFbn4KhxXkcTuKYoiXY6hTgh1AEEEoSpqqgxatubBhRD
J/v96TH7SgoTPSzpe1Y6YgCy5FVvqhxcCXqxfV0rm8VE4eSnBGZJHgSrEof7yKwvSk6D+KB7yRvj
VBBb9cLzXHsaHGAMy26Uw/DjFtrQtJDA87bi3ApuuP9uvSsZjprbZyvRYYHMin84Cm48e8k/wBbs
9o9OzY6KWUes25PUp04FWWaHMpvZ7N0rRWs41KCOKPS/lKRI68LjZj+T7HMh8bdBkpOKLG3kc9iR
FpOoM3wOEwLTJvKtBaeGBHuo8Y7pQDHpuIFPG44OQXc+3v3xWNbJtvv8/oeQ7voTqq584bohr2/t
7JTPBOjlCoKqPIFfCbeiRVR3QItrx9H+TFJ89KpuC9RcZHV4OYxb/CA0MdB6XMW8jdGC9OblXqAo
nmZ1bQrGyNfe0bUiGH26j6bWD+ekRHlnS1HOaT919ZwaL42WzyTRm15QXnWc4cjQg//BtFQ9zCgv
za+I9YoMqMHklju5r0xbyWmP/b6mVhXKbOH3H6VwzHd1sLk8N7lxdOrQHyblJoINbmftaIl2+KO6
2W7A0bLeFqAIDBzucdjP4b2k/vjmv4PPuv25EjcVyfaokG44WqCrVsQ1lhd67JsVQccpHT9WCYD9
2FY9hLNNvfiPwi/5xCmGrqqHVxyfCMBas2qmGsGpHuvBg0TD/bkScyNc8pErrJZ0gR/1V2wUVth/
y4se9IswBesLLwvRTfsM7gi5Q1YdunfCnr/+UVSWf0StKoFHqOsydLxDjWYoQQzO6iY6UHp9NH4G
cuUwOeHwvNPjUNn2vZ9jH6SDCbuPSxxCo2GXe5kpPpL1/JHvXZGgI2F9cudxJsrAB6jEbOQOS4i7
l0wF004NaTtCMMbDi4+sRnLfM1s33P0NDoX71XRJzyNWpZFmfG9anqsV/vumxHGzr838a53rgHE1
Ai6MR7DQn4mvwYCV5TBM+D2ngmD3/s9w08pLRvbhcpzp61kL7k1cE58N2n3UhHT9uIpqydE0AN6O
2PpIMrDP6026EY0JSb8NKmH4YLoA91LefcWR6wg298NBnQkNPgxeAv8e6iGsg3GUaxmR489jB580
+5+d7tqPKwSBCwcb8A2B0/K5nRlkx75CdVJpNbQdkMzsSEbrgmqfp7zEhnYKe2qxUzKMqZcHFn5V
05+nPCQOOak13ssbCqtIV2AEwPUpdzdGgcPqujb3kB9MfvElby8X0nUoqW52/Id4IAzS3HH3+MLb
2Ga/MBK+251s/aXSHUExuMCxI+QFkqSJBqac76KF9B/i366w6FgWM6QuLnGgXvi1T2rPJrPtiuSr
x+E0pfsqY96J88ettgVoGmZaC+Gq9zxNnICRSQtDAywHkiryaI0R9Qh8QY8nqM3T+PGfdr/hLWFj
6o2jyOv4SVta99KDoOYpGDrA3nvKlea6l0Tih/ewpEMWsImRCYRhVHozAqEvoX+4rw86ye/gF0tU
toDn8VvU39eAcl4myoT/LTeg7cYIq4pF7SUTJDZnMRAVMqL1VvkCNF/LSnk2QACvkMjTe4Wlbumk
DwQuxNwCeXF6KkIvo02f8D3Ifu7WYT5IvPG7Ney9rMJn+zmkQa8kNOrrN192LjcQ8a4/beAx/hsS
k2YKffvoSlJ2cHFnbP+mt2cRVIlYtAZrTdU4LEwMSHk+Awtj8dmMcQ/59JZ1JDf+pibIas1LAMSY
X1hZXo3v1o6QRA+gmX8UR9iSl7QsNA4tDdLHO27DvPzs0DBVC+tn4++cy5JaAoOjtnuNKcvWHQ0Q
ACiqqyWbIzp9Z11TL95gD188gU7pJyUMnO5Vz0BDmjDk/ERcIYE2EOU7N7wWNTEUyWgUki/5JTii
INKssUsNEMdOTgOlsKZVyTDINqHLlTC3dr9AbDxEElq3rLbxbxe4475JfCSivdoDuzfq2lh+sCq2
nnh6K8GZXuGbfn2auXAlqBPgRujqp1I7Y/ZT3zs4l0LHw2EYiFYrSo1ts7URdFBieKxcgmjXCAhw
J+O8l72xbDf62Kdpo5DEihj0rBGqErWYcaRtCtqp2eKQDVJmeEnvYzKIG7xtUZeDnbl64iUQaooa
z4m+eRieShrCFzBM7Pe4rs49JnZFcDZrCpP8IFa28ZmbPd0wf98ThoorGKoKdyc6Xj4jtE+uk5JC
cKLknRo6afW8kV1sTq4c7De/fDzOw14e2ixTeMbm8ARxkOPKNiNY0vVZDjoXLnalrZ2ItirbHDBG
UNL7cNUROnRhsAKozKGbBxWolUqjMJmJSOsHk7c3jFVOndNkbMkXa/wlnu0lAij1rLtxZUMK70PU
D9uS6x88qOpJYuqdOnJVgdCgTm6nDGsWpc+vdox1sVs3cfvShDYuH1bbYfTI8t3AChHyFKSd+rQw
7w7+XWIndcIT/dF3Tmu4dCCrd3eNhK+kb6wEcYL8pC0uX8sArE7wd3pE7au7g9VE/iKLkVn4nHF6
QV04wAfrSZDfvNmOgBG6TkshfbhhCAGETwiSu+SP+PD0SNMEMDL5yB75LaJTm/xRcka3TK7nr6+5
sLB2/x3EwXKcPEw8/n/Y/qoMhjr4xRC1GvcEBmzr93dt9uG59s1VRZW0niQ+X1tjfjwEWuB+MSn2
NPjDRZJEuZXpOwWVYPAujohF4/ssi9KZy8ywsj7WX/hnyae9eKHZcUXT388ahh93Zy4y+X0ub9Oi
2RoelOiud5n8ew4dMUSKWvzc2R7IoeiZigJ1sQ0itWyyEaVcl4PPG8lVQNTQdXEvMK0OFAI0Ia+O
Omy/oEsUQqHLjs4K0M/C9As3LWZUZRUaoq6eME3+gzkLaV42UxjuRhQ04zem7ibpf7341d2JN55t
KkLnUGwfsCDFQSqaz6s1FWQTmFMwIzaLVdTO4aw179KRVQzRrwi6Ei/yxA16I3me8F6pcBLlBt2c
qDYwENcIYJnQPjfXlMn3DXhSjQXhuFSZybMsihy37UYBezTqrrvpX/ZqChyLLls2bHmDPVX9gowi
EoRipMCz7b2LD9CNfjeAKtu4tcqeaCOw4960YM137FHIlQgdqewQ8yrb/cbty9DHDdCD6JcNnN/k
phFSNZzjYCgb/2O1IIlsDcwf2tQoit2WkipucnR9AvULDoIMuWYdXjFKnhq7UUZks40Nty/RboEL
r9bHenftosb79TPI4gmk7wyFN6Ub9bTDfkEJCtGqeEoGcZKwZL1WHjAlm62TmnDrEUunP/tMWg14
mD+6jLMzAwP+CYC0kOcGjKU59tUsGgZxE/ByiLHCrnei3pZ//J6H17RvmpaPEyhPsoCtIFuRX1Qp
VUw01fkMk0Q0HxD7ROVtFPF4AeUX650r7uS5uDmK/iZtvPgpyyG7lY1eoTS+R020nJ9oEGVqsS1I
XtPNa6dOwMRjX3jpULDolXN4mruYFiPp4LK8B4pFxzLfW//vg8Y+FlSBjxwBHQD71ZWsR/CU06wC
7ws8GAdYEPYd5fMNh5i/isuPwTTwf+a9cmMy/MqYmI/VQtUI4gigSnrWN3Ev6ruZ8KmYrTBtRZ8B
NxXv1ZHmwM987lXIXcQKNxU566PuqHzwTN1p+zrmuEMMPz1s4MO2zNZ7mWk0PbWwN93mGQrboo8x
YGvlKi6KE79m3wgavusaC2AqXdVsTqlb7X5PNwZRCN4p2kViDJefWzhYQdd1KZ+xcygRM0EhXKRL
JGAX6McEQz1mWE5y8aU5Vcow8v69MsO4IM9/E2kzv7yUSTdEfQfltWVJ6age/8aZjqqwT5P4jr+0
6dF6J8k0PaniUXJEBEyHWcg4ZuIQLq27KYg+xEUAohNTRsdoQ24VjQ7JBefTLGbEqlqa/dAgQ/z4
v5ZWQy4AV2LLVSjp0qXY8S4hDvLCtXHVIAQSPWRX/guoAT8eKkJghN/RCW7JxPAORBNDrP+t1LJC
xTn9YQFgULGVoy+mf6Uh/ross7WziX6gcsZFP9ms2v2HHIVcevzgpHun89qDe3a9cdYWEPa5H+Zu
l//XfhW6Nh42E5qEV/YFvpfEdHihVH6E/l40YDYgT2cmA+gwgjX6VeIw6VksMHbjBieQkOYff5DJ
YzwFq3DCocMW/5c19BHCrmDPIvFlIrGqNmnVNuV4NOcZXEwMh771+aeMg7UxU3Kbx2Jd8JdXREO8
WJLEdSDwedPv/KChErvnxE7u9Xiyfz4sqG+agYQFZIC+6hMZJUf5XiFxL4xFiq17NHUVjMAS2hpw
/+ObikYkd6Pb02kPMB3DyV5Z5zRhWjjGfJHQsyyWXomHEMSjo1qQDl+/ERnev9WeDsbyjii124LW
1/LUmbCSIXQOJcdCLTXkFuJWGCXVpV/DD/89z8EeNW3ylE4iNG5A1xyY8gT4FZIKKBMv1NCkSgco
AK7WJVEh3qTNFpmidjpabVCFoSaBDdznGtXFbwE4T4CRFmx0nXG7ox044TrDjOjqLU9AmIz74SAp
RXD3roz/X6E3BfxdZya9X3T+6yhCRxr6Y1kgE8oNq/4PDkDRsPvxvDGdclw3NQALN9qmQpbsGETi
N3iV1Gz4fj4Ou1gQzSJq36MZ5hUFpkbdzXM+mDCtqyK0aH8soyDbYs1SnQzUTfTs9ryE/ruW2cBZ
M+J28AEI+85qF4uD0iomvNiG4XvANnCOsC4mMA57zylZTY18USJnbwEUP2xaMP2BVhuypvos7UgV
MwaYr3i6Heb8dh29SXsnGzyac004MUAFKvx+QCtLQyQKq8as87tB91Q4URpazuvWdRbL2rc0JuPa
jI1Acf+a8mwkRPVCWIBidWnavX2WcO1egaFa8q/Es6cReZt/tdgubseYCF4TS6D+2WUHyzZfoRPR
cjq7SNHfRA59CipZZeGccSQtI5gjtdgZws1Xm/ed7x0MXC/rtNu03P8R2clA/zkwXatTRJ8+xBQ6
qG2eEWs2yI9ziTz+ufjmOQMwAtmdx4XmMnVG10xOeZI745lrSugPEzQr3Q0e5KHVut45DntKrVFS
z5Pd9ReBzmDbLrdUtDllCjVYU+6RwpINb9Qu060r5Nakb2H9NLabulsflRX6e/PnVxBwG6GXrHT6
F9P9UDbMrfvQ9GKVCg4NfyTn4VjRDvWSoXxyU5R+FKSq3FYnH5jG+wgyvlpZOt9l40Mio4XwN9hU
vO02vaLDE4L3yM8ft5ebzyyfqRWvvXUPdXMgTRjsMCT8nxyNOQw/yZTwuJn2Bx3+j8HqkB++gzCW
xGzCDgWTGhrSfvBr9sc1djCQkriOX9rCF/5Rk0kjE4/YVwiQoChAG6Qx7K3jnM78gzt6u6aqbooq
bUPI6ZqXtLJhVcjnmixxPrbz9VDT+x020HCTT4B6KtI8xKu4nAnRp6t4oEoAWtMRfRSHtfl8zIAk
wJUXu9ohHa8QOJAsRz/GcAMHPniaFlUEi3oTQtGtU/SApSxJDlqswBdcTGn2V9rMXHEz/P2hPI7q
PDi07V2Mo6R/RJQMiK2MF73TJ7Y0cWpDQLS5ElwrAKb78WGSihw/OU6NBjABc2n6YLxEQzcrHZG3
ZMWckEzHQilzZ2XAac5YybABJqvbe3Uj5Vd2RGkEc6QE1tMKAu+6EGLIwFXzAU4MSHlXkdCWVx4H
rQrmfoVdb42wu+ASAM8+8hmMoxqLKQzPgmHzWTB2KFsGO9AIgMS4b6DU21W+FrqX1G6ilvvtIbjN
7t4tUg63ojUFo/zjhoMxI7UtJqO4kWJYBq7npOYJyFA1GOC8qo4JNNRliwCR6y7BgzZFBw6K6uBS
SVmRTsujNK9xpchLxFZE5ZAbgdSHWEPBBKjX1vHhMwB9g/9vfbP66pGcvvBjbm9DttN9YZ4d00LZ
5yHYPjeY0Fk+PulzqoTRVUoKPO0wcnmL1tUKFiBWXNuU6wIC+EelU8UqRbxw1NSNRlvQ/xXkHPI9
CKuWPw+Q0O7UhsWnljOf5gz0pH/EAp4FtYN5jySE6vhAoSOMEjW8uKuhRnqOOKZT2B84Uig27/Oe
YTpc/wpM2DTNqJnzG2F52AUzsuzG2bu84oEiJ9x+xQB2Y7gc22y+lg3EDqM4tElKxAzzT8sC9CpW
xsfQDMHrIpBzCjoT7HJ1fHu3wQORmHJvDuF71w5np5e72r+Du8e17zSGYJDhP2QKuIn7nk6Bx05x
fI9M4Zqf4LmPFG3wXFbunkPzqRIut8YUwITVPLHksr8nIlTf7x3f6SLm04zGVCBuTIRyeoFHINqk
Np1rWu8KUO2bsnZzZ/kdI1ALpJpRuZ/lefgSlFlAqEAJ1gOVSL+f1EF50QJvaXQq0N7mUy7/+G52
O05/92bwFTuURYVlsQ+M6RLhSMvP7cpsBGn/7wznE21KzE/LTPUAdwHbBy2CL68xch7zfAm6rLNR
VBqNJNb00b8ht0omtG4VZTsfGB1Vt4a/cIOaTNPk7WPSvNBJN+h6X9gx7PZ/qbtSEsDy/kdTMme8
+LRr4s/ehc1t62foNiycgg5HKHHhAVsiN+IlUiz5gznlvx2DBcmRSf0AcbFWu3AdCh/DcIR3ZLtW
4oJ8LV90Navfv0qAe56j5VG/yn1jG/Jslb9v+x7RrwkQVyCFccUk3EqJUcT7p3Zaf9THBCPQkVJB
QGZRXZGka82cQpUHQmMs7DJtyL61EOAy4H0b+tD8UeZVuwNDOOoXvScMitVLC/12PmP4eQ+SZ/dj
u6WrJ9ZIly2IHi0DYGMrDu+RF9x5jCOKmDdfQBDKmtVcMdXjZm2Bzf+Tnhs3TP5RsoaYbmtDLHKm
k8KBn3nGTHA4EyZnGT5onhtf1kzhOd+yHdbtunawl2oCoiomsIAHBZNrbbMhHeHqQnAOzZDNJWlY
Y1hPtyE7Qwn0szuADFYEAAvH1A4x9Z7SOUJA4ke58MzPXGNGfrG/qMKgYLKCXOctp8oSfptW8jnu
ZXu5/MP4qRLATmkaQBhx6cYMYFK5EMR/YMkZ72+fhyh87qOOIeJcivcGWzKoCe/aiuOCzbNmWknH
i8bWSxeYij/2VEUphV0hW6BCZs4Hds31oySVG5H8b/2wvnt9puuy6JaPiSNgBeYjeuHIxQKXPmVV
eAlrycCbAZvb9F13xAnBseGa74RzhDEU+qKnYrcoXWpiN/QiQAT3QpRG7eVPWJLQRQaX5BO4xQih
Q4Y1Y8A0yhE4MQG88SaIc2bhEMFn1wLwUIwPaQK3nlcudyFgZ22ZqkXnlquTpq8QszePWqGBPex1
GtROHKInejWHYwCqgPag4z/lAKZSbntoIZF94+wX/i1klWKysSjCDGtsFmgwcjEnWDWUEyOnmPam
fEDf/wu+8v30Ox5T7pdchE4clE2ykJHRY3pamnwVP+ISjjE36uuSSOxmdpa2NQAAJ5aCY4MzEZ/i
HrMLbjDP6zbkOc5FStn8OBYTh8v3l/OB4KQJx6hdn7r/L8Jj2HUT5ZNdfjriStZLJ0qDei4DJLMW
c5TUEHJNT1Y2srtAYgsZAdJJH1pExyKch7HbkfWcwvmFtMXqz8pZ+vLBF5Bc5+2yPgFNZoR1o9LJ
x/2H6aemRPLn4dQK2pDFLfzE/USMH5wj9ps2QvZ5TKSTZaCGoYuiOJiCOA80LDbc7AKbrYkaCmpQ
SxcatjWxjtRM03LCqx/uyMjWlw0WdJaop2GLaRLoi+OCBwhuivqhUcTniZ6A5lj0P97hWOmy0eFy
xToQcWiRnwDU914lmjSBcMHndn4qkpCB0sSdsZ0qRVUKJ1D5Isms8qf7zxd9t4GU4dptHZijFT+y
dijbW8dpPbjOAfIU5vcnyp0OADeT2zKd8JpnQW4CrozVXjdVtNXExNZewVCgmcvyzDXhkYZbyZ/u
TKCbhqP0li1q75JJsX6+lr+yJVI44LIXWrBj8e8WklVLqRDLFIy4J7KzYZPdUsmLK4c1MtV4YJxR
8oI7FFb1fyOinM44l8he0QxJNc+fQjam+osb6m+FB0kTYHii/P6ol8dANVQxPU5vlSAEsG8ddhzJ
Mb/cBLfGQ95WCbY2WfmrUfFMjJl4nNPjHnf+YQaAuA8SI2GO3k+UvdA+t3Q1dkGgO6xbdmvFdze3
bfk/Z11S4a447SfZz/4pseqq48C7DI/44q9K2Sl3un1hQt1tIvh0mI+rsONbX3cAsDpntrE2EFg+
p13zbFwNdo9h3Fp63Cl4/DPY8Zr1U2Wr8l4WCtZ2rRs1kksj2EBa7PejDMbDKFMCoQ63ksGNXKRi
HeQJWybhSi5tgMChsUGZGEtAs3/m3geV3eP94HJGgIZh1jtW+bCBm9HA/hsKvNc5VsFsg8CmN1ta
NXuTHvh3Kq+KWBja8YE/gGLENSGONIcNAXe7+nnU5rU3Xf1TrPrniV2yyRNQM2DdKAciN1iHWobV
CljDui/8mMTCzmrs4I0LqQ0TStR/i3wf4f3WZabDWGqktVU/oMRkP4f+ZUv46hZZX/k/3s0i6C9l
2sJ7jHtTOAHE/soqIR9F1Gp+B+uNLNGkOA+UdAOmb6YmyM72ki9P4XPZbi1gK4PzRutzZyyW38aF
oSYtJM8UA66lntkEyTg90Vjhn7X9Buwzqfoo78/m52SM5MlgkSWUkSv+DlQ16Z4C4ARfZNMLWiYB
WCePP09hytJdCQ5hjyi8n+VJwbUNYjridJMYUSXrr555ErdzLGlSN6eFuKe2aGqQzQppdcmi2npe
GmfN6+uQh9pbpBSYwLTcuLpSyoX2psv5/swB3CBqMUuFMMm8EZ4yEIarFiPQnxgKLqFD0hJo9/hy
0mOf7FR2VwWvdF/E2mB5K4m017YzrHq88CEpWMKDd4Ubbxckgi8EHglYMLnKf1CiO9Bv+vauecV1
cIwkVx4+AgOj7pIsOtFXOiL08VT3Z+4tqzih/Jk7v3xG07RMDZS3Pfp7JEqIwyBbBiKlpr+irACQ
vb+tB7sXRRw1oAwkXf6dYa5DexiJEgT4YmGZryXMlAd822yL/mtKTCsmVwLK1/bUyuAXpOg/UpN4
ICcFjtHrESrUgxfrPjn8nslrZzQp+pEwCnm9yVplKSU6iJXu2NJOHHRQmZLZnqxmJRdxw07omTtn
wwFC1Z1OlLHM1eXT06qJdat6RUB79WKqVSEIl9+cGCup1yiL8vj1Kdezee6Tetg0rt/BJ86ck2MP
Ivh5ItIZQtT17Evg2avkSddUGlgbUQPodl1+FHuaiqKzFGGlMYJ9ZIfv9iF/bdSgSyUvKJ+/8fve
M9wY5Jzc2JRAIWhi4AQZXRGVtYdHju9hX9xp/iK6FZVDfr6mj5CBewEW94LHHP9C7n11gU5BxS27
RdTL+B/muuGfCbaS+RMXXKvgOrboF3QfsRykNwg20+7K+Bi7J/POlfzlyAC8pwKFnlPXy+mirOXL
ztT6srDKONOf4Btt7wCzikWm77Md0PYOMHSiiMMs0wt3UF8sQHqnz3vtixkHyPnVLCtAS3cgw1z4
Blg9NbEDIbPZyxDCDAEy/SY5vKPiQJobxNfnXii4a81BOu2qo9lcVGLg1AEkjl0k8B513rVXiQHt
fvh28lcqgsB6JQeFh3AbAg1QmqoilgEx7swClUc2KPq0ftYZBr4q0BcwQtsuvYxubgKP7fScit2A
PxzMBzcQNyHD/XW512nvvJl1HpjTsSHpaX+k9/kw1OgH5PDw9a4RySx02gBFi604yE6JIjzVNJIv
HDijx9f6N8/9d+WvUBM3H6aLCqgmXVdZxtiS0fBL5nfB3XQX1vaPpkBdmUSSSYhb8qccDevjfAW1
vaaq4BKzMHbli349xyin+qEIGooB8RjceAwcXfpY37UW8zTIs1STJbAFgypy9i4KcwZYQi0bUd5r
kweY9rbp1Uhgh20NwxiPFpCk5pRdgBl7YWGDLpJsxWd8FQMiS70Q3PvsyKFCU8guccpvswdEwZ18
JgySndTvVVLRPkD9ChmAWNJ0CHbdpZ4pH7I/dfE2LGiuivKVz5YRdinxM6M+Eoc3accKUsGeY1GR
sJv0MvdGyk7OCZIEvr7TVGgPKqDem9jV22OlZyIKbCw9EhzG5Nb/XO7vyC37oYKXzJhXJO5vd7B2
x2wdi29bhtWDsN4HpZKQwsePUsNplc3STiffM2okgKM1ceSnxJjXgw+HHU4ZEJ9VgJUYz4Wmh8d2
KjyFJT+3o+vjDnrGGoXdbsMc4IDXNR5HIOYdjsJ3hv1qlc0pvETl0bWEGDe91ng6yB1lgxEV1q/A
yaNnaFCjtKGvFei2JB7vCEhdZ0qiMGhj7PbaaSBKtLtg/RYVliRHXyTAJtOKjE3mhEb0lsJmhPar
zsBzHt36KwZFF6fJXRMXawaFIEtJkme9VUQJSp3Bg83wYuTqWLCyMx+XJuyq+N6UAkSgexNYm+ju
UM5tKGjtJ66bzNfb3s+TFyBTYEClRANXsh3u0Q9am++J593q0d4h6+4axNr4wsGfuC9RPTiZFbSp
csQDiOL9EYLVWI3Jxtniw0mCBdTIq1IJgL6FuzWIihJAM6enhG4bpjc93h71o/fpYLTuGfnt5Ve4
ZsVBBexhAClkBjpotIkYJ4LDs6vEdFfGsEsLLoWOZCTHq5o+mieeuP15v2REPTG5BMhcE8lx9vhm
fGZo5o6vXSjqgHAyGgryto+nWfhrYGZBlrs8CXM1Kw/5yCAIi7deym7zT19wdWqCPhedQ3F5U18s
D5SDmreGuB08pldME5BudfqMrXFV41dp82Ttpd7k3v9wvSqQwqnhjVdJXwIpYX6j1cMHFHN4oWqy
7eDIr++1lPv9c9FAmna3du7DVNRUc89ziM20hrXiq8DAxETyS5QFGucGtPHnDs5in7FMh06ng0xU
Lg8HBhSoO9BJNJXB4/RclUBg79SdaUeY3KZXjXDP1IiSd0yYloIHVbgqXCGRImlsHGHDZMR+BXzM
+0plpgKeSdrvz4yjv7hk7KrT84U6HKzUTf/2pTRvj2zBzvZdlGdkaKyvApZWMTgV32VX7oOc/OYw
uTcov3BWlkiM07B7LOTql3ujoKxaSwUoMAjPNtQLnKL2DIWbbTr0VzNWTduJpZ3JEj0HgT6MDzdH
IIeLSM0cX5cd09+8wu/nxwY/2Y9RmG1xo1tXhnFslzvDsuBsaWHG3SkG47/FHmSl3/++J94MiCFk
/K4JPUaEf+d6Q116YKRSIRQSLjxfpuoKya5p/PqSevMBRmJUsKmyETbOjTBakSGlDHgKn3uhTfqX
KsBx63HLBXyhMttP0kE+satPeeP+dXFKC4d3mhJRCTD+RikxBnjmlkS+gF6Buml/TACg85hYozXg
nO0klpCURSPEDIRxnsycvOyLMRl5m7LjkvpRPRz1ysfool1V+/yJk79AoLVk03R4uW3ckFl32nLC
jPk+4+p0BWRnvvigAgw+bYBrALhCZ+D8N9gVm+8MeEDpVKOhL2eHQS74SvfYKgQ2jwt1Lk6U+qn8
fySXomIRx16SfiHfW2id63WEn8rxzrxtbMSCQ8Yrsv1Y58FnrusMztVOoCYNadZC1TlI51dmUkuw
Oh8Th1/dSaqvdG5aCTt6QZV3owrd9T8sRMTR769SJ1Cn0s83nIo073OnKJL8iUYslVVo/3GW7TXh
dBIUMYKhFswEe0b7QfAvVdyJCTSGuRqO5jX+gQc6EE0wMUkhUe4MPWL6+2AxrXRZgGHbt/LgogY+
fKnN2ImV10YOwCdwK87bFgz5e18DpXNGlx+vEZws0PIpKcRgIpwWndWQVyvz+IyRV9EGVnJmrqlK
QPes72WhoH22lO3cw0SVDhk3HPD47YhrpxGrxCzA2CtQ7ROjEW9N1tV4q+JfyAVklYznQn4johVn
twjJNUq/lLjpiNqa1Y8ay21E52Toa93IN18WQn0vY1v/CaUexli4nqnU9OjcXJw2Ek3nMWv4qSEu
9/wSjuks8BnGkowii20LrPeclH7iC6O1FbUdNPZfScEJi7zfF3TCS6sayRO9IltqOqMnPqWiivgl
ra8UEoqj4AIXQoY1vCY+TMRFH4UWrpdT8OuZDS2HXHDAFoNK4fyPwu2TYFxeX6V8itH1Wx9iC4hW
mn5/x3owwLcsU8xC+C7Z1JgI9QzjGvfaZj/VJb0sLX/rSLCv6wh5js2WO6XpLelVaXj8BCB0q2Ji
/qnXwETI180FH4byOvIbPdN06oY76iululS8oemKYTwnUDI/UtIf2FfWroBrpSeyyzPE2Gbjw6eA
Ilhlps7OECMXTGqC3LkgJVnLN6HKA+se4M+B9AEhL4oxw+Qcx7piIQrAVABF2ztht7QWZp6pRUoN
Bp3SfRub6FTipn6qVMsCMZmcA6s+hCAlGamucKURFTYkr23rU7XWdQSPkKe36ar3AbfB4TnDnDu6
Kxgz5Qbf+frdokYMVtzkYpkPRRgihEiOQDJtNI6IU7E8xXm4wjcQOeF7mNRVLQyH4zqERMJVYGzg
Y0pZOHxUM4y+Gf+1+EtsY9NRWnPaKAFcIY9e7tjVvOIA8xpN004c60kPt5ZVHgT0yoT9tdexibBZ
M8ejU390zFTHo+ZISbvQZyvlJSorVF5b7sOm0xsmC7uMgYd4fKJwkbjEKHkPvPSa7tFlLerbDiUh
IzzzOf/u1JJwWrEy2Il3W1gJ5d2jOSIKGsLCanIjvuKI1RbIgxL/ylyFoD0s5PFQhc7oFwSSsXsk
Qk6OpaTEDEp+50nSAIUhQZtP9PyZwvaMFHWS8uc/XtN4+ZEeSXUvsETXeGN8tZBrRyjIrGLl1suo
BnnUa0+/fEFixhzQqmAQFl26msFmzquMOJI6xN89yoEIF3nPiPdiw2jjQ48zFiBq0cCB609CFskv
U7ORFjsHx84zP7zIk65/5xEbYKEGOasK5E6lmdm0EIwpW1w+wjvuhCAM3a9sQM4TkN5fAgcN0u1T
kkHbRrld5AGQfZ5OK+G9hDLQTMDHp0qb7mUR04p8XYRKoxxxBSTkmyulOlXDnw/+nLx/8rSw40GL
hSt2aKVtPKUn7fvMruUDUBW6DgyCWGfyimqGkBrwuFYBcot/jNsGNUUKwblwc6yQ7mcTzI4zuVN5
+Mp4V7lUrYhk4MrgF8+0GEoSMceeFepwSm+pAAeSwuLoFTp4eqEDbX2DQ98ckxD1rGkLqgXlHcHq
Ae0Y23bxEp+/CxwOolCFgaLvRqd7o2yeY2UFghAfrzjWGYIuiPsLu8VtdEL4FUtIHFxxBS7OFV3k
zffwhIDGcI0oiCpuk1XoKrRcI8kM38XKENrlmDdmgQKJ7X0PXEtibXwMK/EPWl3sAOlM6cwhVZiZ
unyws5t3LVSRo4j7JUwsdyn8xKHh8tFM+uaDOdE1Nt/lzd08gUc0D/Yo9cQXPDuh5glIpcb+2mJm
+l8QXHyoHo4VTDA41CR3fdl5gVXwB5gz1p/oAo9hxMngieDgc1sEZeomJHw5exA4yhUxTXX1egx2
UWsoClcEibNIz+eD87jlohWkQi+Y6Ava1sp9K6cXJUp7aWlyvCOHYsWpt7IhlVv/F9T25YgHlzYs
nlPeP7iUry27b/qqOHI5nox/eHH8JKSMMoVj9dgtjfvIaun94Efttj98qkKri+Vo1hwVrS2wCCnq
11ZIDeEwEFWAP2o6cnmWuIzc7aqitIJOFasJDhgWdfY8KFv1iIxKbpnUkh+kbnTXaVLfex5jtQjg
LbV5DlIBFbUcdHPHDkBD9+rygpgYK5nQ4SdYGh5r3ooQd2tkZHqvOGmNMZdiZs0MRRUpFYtf9WAD
kI2+9aM7XVQ4T3Xf/r7tcMGE5RrhCKske2FCL706H0vEVqWNGqQkLWAivc7GcmPRFa0azhARDr8B
j/SRqRSZJ3fD31FzWjThJ1aalKrZpvfDOjjowPQMn5Jz9DrH3FsM/FajNnnVH5mX0oX9O8jddXlw
GHHkxUW9VlqRCsbSH49EyBOxup7yvmb7y8B/BdlC9rQA9QIs9m5L8H3Wqr96YUc4h8zN/DBHjOsp
3OxAKfipTox3QpG76ul1jhmmFiT4WDwujN7TVHFGJtdMvZC8V+i2pvdwFFsXBWUfQ7nmbt7epBYi
7t7cPvl5ciBLbQgDlDQJnj0BmZ+vS3BsrRND93Wu0jwkLJDE9wjATjquapJw7CZJ/oHeQO5If7MJ
MGY7+vWJEyy28ejx3yw509b0QcOoy6VZ+YPqQVtK+a2G+by7B5L7EV6wjBlRd+RsXDzf3OoZWglc
SMNX/4rDVgDZ+PWu04qA7Idfrwl+9LfCsFUiuljlTk2ZJuMLsi5r9KtWFHdRhuqvKPN9qtE/qcNq
pv31MNb8X1mah3T4Dta3jmW1WoWvpEN4GteDIXOHy/t8kwq4igqFRxje3bI/1kX2G+1ckvFI91aQ
UCHJ1pk3szbUvi4945UQkJRZt7/KimoVaqo4gwDyI2vQImZeji7Zmz2K+NwP++PvlsD3co0LV4gS
efm+ppuzw8Uvy12ctmY9bbmiPJ8x/nDpzg6/bGzZGGxJ890jFK08PB5AtkV7inlaMItg8LPtzhRk
ugjcuwA0RPbc7PT0pgNBU+3bKg5hgP+7Zr9SeJ5HqjtGARfa7babRASQYqm0dRC8CmAwnHOGLdSb
p6NMM111wtfT3WHwZQQKz69GDjSwec94lQbwJyAOIPogpQqVI6/W+Rey6nF22deen7yV6bz6MrlC
HBLVe5sG20y6dh7GkS+SnUD4HVkvIb6gzXBtio0SY0tH0vvSVNJUZsKK76i7Q3t5q55kW7BdIiIR
T0WHX8P9oQcQHR3gTt+adTY8zncbr+ru88O8W+903vN3VRVvUS9xWmyhVhUGbDR+6GaaG1iabYKD
6jVQuk8ljcjYqF2Zh6ZUeTSHhm0kmiuFykFEK3+aMGPKCZAOT7lskk43UxiGp/H2T35WaGyagz7e
A4EMbRvIOl7i+vy+EgF/8P4RWsKGbUNNJKtDpDRmVVXveFdOWnfCZxBh8cpYQBqg+RVcKD/SfTMN
tk80YxTdOtth/LgGtGkI6dbhszMAmEivtptxZghkcZpczM0+O9VjB3CEKb6ISlO6EKkgnuXqGabN
I3fqsj4Lq+KPzqI/fpowl02L9PSj8ILMuo+dnVrg+P394j1mYyoSV4dvf72SliTk54JDO096DEVZ
e60om1/qDc2d4NGURMGzPXPuOgws4MIOsXTm45x1R/B9vg31dYBKr6L4gx3c0aIR4MQaoEI1R5Hp
T7g+IfcDCnraB6QisK0eDMA0CmgPkhjy+dwoFBHS8CmVRq255GJ7ZfBxayuf7W+nVST5v4BrSJvs
Ql0fSxlZctNVTXErV/ktNe82IdQ6637vya0GA+LS0SPf8YewY25EHcBLx6aF3REIyGtC7x5kxKHL
aotFJ4DGNsTBDgh1VXuyo5hq5UPyqRsBSWcXBODtiBS5bW4+qg/6BTL3wVMB9VkSfGus4I0+9KG6
aMrQhfj74QWOSdFkAC3TDpDDtxduSMr3lb/uY7E4NRFRkE3R8ZRjsBNYU5NQdFogWzuUN5TqswwL
Ut1nnMSMUh/Xx5rd3kbyYEcfYl4tQGCWFZqQGoD63ZUk9tNjKtRmcXOVjR2gRlUL4HjJjCSgxyc+
owoM88GLYXoUNJio5i4dlW0X8saSMKK2UCWsVOQhw1H2DNAKkuoNMk+JP6vlAjtQtr+uxH2bm31W
zQr0ORBXL3VDMdtfcfBMi5DYR67ESk/5A/do6bL7+BovHfS1BqMde305MDlo+CWNe1my23MczPcM
gsDQARDJ3qLboX2oc9n9SPR/t8kc7Mj8q2SRV2vmnn6wmkFO5lr6Pb9QLjmtNwqckWqxSiuEpmaw
GNjTi0n8OytchWDOa2Lvr9cZxIOs9wb8tJ3m1GLS1yJqkoNfnC/JAwHjGWl4nbWynC3c/TPqoteG
phNmHsNdvFfajOJkJgYiFL6aEtIzFDHu0bWwi7QqFfTnQPX3GyQYh6CJadnSqsT1RGumQa4a0KVP
JNVHCHxj0ON0/ybsSuA/+8Q8IYXVsEQOb3p23k+ukmc3Fy9vz77LYeFZQqBWgw6892ycvAiVgfkr
ZwbKa/hWDbj3OGD/G+PGwvCSX+fmTcaNu8/fq2HLMs5pi6jRAm/bQtzWMpfvOBOV9SFjYUQaNnaN
8sZj4A+vThJswKa2JWzwpwfzPK848nuVVXXkb26pek6adL5Qu2tWFoRJ2Ir9TVVfha4Inzy/4a5O
akTQYOZFy3LV6XH0M5W+sQLh4e23MvpZExQhfA0qgr/G0tedVIg4+1zDcyKca1wXwJmO4paYPbS6
EWURA9Cjrf5E4moTGm2j4RZIs2nyYb1B7+7bb+1vuPS7wZ247aHoqI9+lo4uDI7qK9qOLvtUyYnl
guak23xtCOrPkErK7x762KiL9fk5K7Twq1uy+kJI3XIZjzbIojRmYONFVQEcdgBcxkORoz5loP8W
l24PIR8Ni8F9OICev9+uf8K9s0pmkOV+VY59NxImMBDOPIhFh5CHW0YyAV/tzRbwQfQwDDqjr6fH
W8qvkBrW64iHG8wvAf/LjbXmzWjtyEba7h06wCjRw/WtpAX3ORpr1eqrI7jbVR/9gEiMxwOFCkAt
EKkmRGPb9eaQMHmS4r4f7YKF9+Ut/X8xxu3kY34q3z5BYb926089USgMXpF3hwT73yuBBOSUonZC
OoxDXnSdjphxTiFvLpiI8i4kShVQr/GLM7ZfGX48mqH/4YFeB1TpKEbgmwfDuAnPOibsuHX3HdDH
NS8oSG4guChbH+n+MsYw/0XMs85nK063iKZpi5k91ao2jdJDOKkfgoOPhE+I13yx+pkr1wqq7cdB
UR+U2al8q28VQZ+AK0u8wVOOHOyrR7tafsVlQ7OkTyBv8qAqPfoff1ysg3wUmZXS/Vlo+6lcv/85
R2bdJmS9/VtbA5HtxWhDNgxB11ix9gbRq74Z27KweSpOGQTKhoFRrLiz2JAE56CEuTt++5qZvCNy
z4d2h0aCG97gzIg2fre/S39PY4g9l7AUQB4AxT7ZDh+EVCS/PgGuWlo2qrtEDSHJ70NwTUBtBbQA
m6SBrLfGvgRJcHKPDoCN73uJC6ngRoyFANSfha9T3XfcQHFcuRxdXwlB9S4rTeJf2L2PVUHxV0fB
D8M3LhTwju7ya2odpKwOu0ixevaU1tQi3PBd3PBhK33daNI2Dyis7mcPedIqU3doSrki0biJI+lK
Sgfwndq/G6p9F1htUyBYGnb+pmZQLlbS3+r7tg0iWXyAxBgnOdKC59llEbj/IkA6R6hnlmjOWDBT
ypi6zfAlRWKOXuFH9Se5CkpOX8uB8phzDWF/dLzakQp87G0QRWpqdxrcXBA10RtS9dl/FFXJBpOC
csNBE0Je/uv2VDqUS0uqLR3v2wMiHQCMqpPa0luLC8wcSmtWylqw5EJbZGeIKYOe9d3HKVlDh0pH
l7EPyGk3i3P4sMXYvOgIy7uT93G3hXvfZGmE4SAuadk3ginLdKKgyg230jitCGaM86IoSVdptvaC
YMKpn54/8o7Lc9C6qlwE11KxK+XuM2b/PI775tMZEQ9DThCK3LQiujk1NeYR40fjQ/KdQIfUCWxK
mqaK7exhMT7+r4tJczgVkwZb/nUHEzYEL9nUvKsAaiT7yuH9FLGF4eh+MI3sMTqnyeZ+vPiJirED
yUnkbuf3ZTYJDAWfNjcUUS8GWwZBb05q3eDhSL9ferjTWhyFy+B/d08SjBEfrzP1oNbyNX6fWpFl
ZEBH2Bj3OV6eAsixWh6SE39FpyrICh8ceQacfEtBoQzD61ko6xFBA6anmGSi20EEwOi+ytXrB1qg
BmZ1i6WEi1H0DxXhdeWDHSI2zreM192CwST/MXSPXT/hNL+y7jGtmXsObeQgGgcccc9FIgMtlSMu
YPLXfdVaa2Gh6WX9if6Rb92ZGXPgV2oLuSCqxn0qYZID8qWT/QjMpczSldO3QIj+zwQCzNXgZzPy
XkNAaQ8MTK/LaRUXzsg/pTsNFNvNxJsaNW5BvXGINHBGVtaMRJcFDyJ2pFBvEOQ61lZlF6/utUB8
trzVnoTriUu1aItaWWIJgqm5CYIEXSCtzlAQnLh5hY3ECBvYx1etb2GMZ0FFrhf1b0Dl5XcQq8ky
V2+/mXngdC/Iykt6OkVXsP269cbgUeL173iuXW2FwIHbYbHpAsHogrOxfGifcaK/Y1+ysG+HZdfo
xLBKSPUPCvMpIp+1a65TQBvyTelaTFt9L6k8LgZfgaJdFM+OI/37d45pOKGLIAFX3E3useZ3gbO2
XL+EwhdvwWuRUUwi2a6PBaxI7526UpVvrJPAgc9MBxjA/2EMYJ6DffLcfundp8UCkmlMoxM/SFIb
EWpZW2fP4AOByZt4YdDfeBdmpE1T0sjl+z5PF4dwQNjnhZecI1XUtHuj84Ge1J+y6ZQKGqxCGADb
LnOtq5fLE2jH9QWjlMS03ntNZnO++N7FX5OpJLtWyk98E0ivpuBcLbGum+aZmI2lToYkqfUxmYPA
/gtsQp7NIjlKLlxjoEflaDJZ2/B67FCl4l9cyfupVCTRl/qaTz2GW3s8ICyimTPWNI0a8Xlr1H7G
uSQ0hS+upi2ReB/UVt41Ouomhe2Dg0mltz0uk2AzS2Mop0yB/x0qtkiRFomi9JZdp9gOFwy8UpUD
GxD/Dk6e8ENRwn9iYzC2YSLzUX+vqKYKxuvBCkULYx//9r0JbF5OG32RfgEy6ztPpw7k9bZNAVgT
gu6A6QaaUicItVEWQ96tBcj9yz8JU6ldQZ9fqgMtZ1lRPdNbJDa8vLvfVT5exKyCtnVSEf3MiAE6
Fx/Kn6NaXJyfZc/ua9uIWgipfuBlpG5ZDbLWKTZ/aTXxV8BwXNZ8XTPSl0TlvAKq5Lixh1lM0J8j
KaS+FyceJx7/QjdAtIa9RwxZ9ycQiTifPVppLDCbyDZ2DBGVhfoCgb00nt0xGi1w8EpzctWvCm98
+R3YeSoFSIJ6K/34LD0OZNpwE0hgXFV8hRB+DH8DR4edgva4+acRqp8e3kKajLklmmmpUe4Oiyv0
2M0g3IL/aE4KDaSAEQoHSboTPcbX2HV2axtHxTrRaX0uyAkKNntiiFBRzcRdLjzmigdu0YBk+thx
4RNiJ4l3IjCBqVmJWlujOE1uE3uL4FxdeDDmR0f+pfxw9PbLNrr88jDmZmabawl0pIRYEFENom2O
k7DwCmDlGhRyJLD80p/KG/B1ZdAJ0r9vWq6278I3+OHYZHPVh0IUQteTkknOdys9NmKnicAdeoKV
F9kaIfvNkJTQIlgSBkX2yrrBh+1Ev7Y/FZk8A8ewzokw7y6Og5mkSNBKjM8/oOFX9g1stsoOa18g
Z4KFa5AEcEgNKMmGd7hATnRMmkHCu0yAgea7RU4OIdAt614aLR3+NrBIjJptWdVn/uroC4YAkJCX
vyhOABT1PaCMcgTsQlpaqHEfX8QBieiNbMur6LBgCMQMPRGAmweJOT8cFtkoL+KyF7+jOIs/hZ9B
/b3O2ZA5/9z8DVA+HIqCEeIuXfdTSYyXGwtr0jLmESoSa8WA8VK7xTBeW/JCwXdBgNjgQ2LEUQjp
l40wyK/3a8hRx6uyKj1HW9JuhdLEYJw+PDGnWPCF4EuUDbZLL9dg9qPI0EY3zTo+TX+l1d3Paq+b
lkne4sA+Y5ko4cjg1hsgjuSBfk1Pf6z/qCqqB8I1wtHF0RHwPUCtZlnR+78yiA7UIFQlYVX2PpdL
iVZTsSg/LLw+CoDWkIZxKpOsLxDniAiY4ofP2Rv8f4uTtT778DxIcPIJNtq7CxFYmamCStBGKefJ
K60m+Xsi5QIfDJw08AKl/4gHA235BDEEI9wE8ycf6Y6A40d4AwgeQKrg0n+mGiugE8UtwCX2JmVh
7wI01HiKZrvMW6hzKtZs4M79VnrK2vgzoQc5VPAFITWsXffWEj+nOn4E3m3RYiEFNw8HYkw8u8kJ
fLNDslXohUFOaokZwiJS5a3ErmpHrsuAtUHglBvRxt3bhh+NlcPimuF4KukhoPNMmdDr5/WAcG2A
stHnjyN18lmK3WNzSJbogI8aXRd9tDAZxVFsVKQ3tKmkh1mUBI8/RqTIhIjps2MVbxIfS+2NXWcK
Y/JvQY0mP6t7FiioJpyYCl5BPEM+Gc/Scg+TFsDAge7RXhJ7//UZawOhr7XfV8gf1p0H3FsVlOuv
4FicNxmeQScMci9Jmss0Z+g1KwzHEhrCHYNL7kUYgsPVwR1U4GyiV7UKu8UJ1lSctmKthpsxYVO6
1Fl947XL3Jjshe6QDpNFr+Kk9srvWsPNfMrVnJj6i7EUUG280WZb6cEXj1Y9OxzIgeopP6dVa9p0
SoOH44rCOrD2tUCi6UGPp/VTNxj+Yr1RcWuThkjUR2KgFo/5pACBVeK/DULQY1/kV4VJWFGPdnyL
QO59tkxsxdCGta8bc1QEVHltAcdeOLJtqAO/V8cWEXwMBYBPW+KR+kn3/lsV5G6hMm1P1G/DAOc8
rtpj+QWohJybOS0bK1Iz+g5TEMCBxdy1JkI//VfoEy9fdgmYM7L1QlXkqJBZEM7s0VcnAIrY2XNl
rhtMokCTMhObrv56KZ0Nv1VXO0s1NISSIbODq6E5BvMpm0dVZaorTwOZ8+N8V2E/D++r/yofFIMt
WqG5AcYe+qe9tz0vxerad/vn3Et0m3Jd+PavdQAo9+SjFpOlFp2u6ln4bRfN4ybHJzOXrsGKx4xG
FU8xILaRoO8Ct+avSmJvwBzWyIOqbL7QNaWEcuOS9svhmBCVf6RDZbIQjQmoCZyqsiHg8P4m55Fn
NC4XeasnpbKRf2BaVPxFmJzSpwVpEUwZfWCcldsrr4bv8VwEka663M4snBT9dYSwznoh3el0cdvb
s7QKMeHlvRj9i+H9yslvvmd8TbCpYhxB/BWcX6boHY3uGwZTr4Zi6/uepOifGtOKlqFGaAScEi7B
5T5NDwRdUlkZLv/b6kAhdL0aRSSzCJha/SsUCiOW5EyjAUdc811Zg+NzPeY8Z/99c13vlcpm2Nv2
9DoXvPra6qTfmGUyKJTxRNXnILQY46F3PUb0Tk9b60GkAb/L/CYI0waJ2j0inpuPmjjmuN47UR4D
5PYZYPMSEuT8c0wTKzLowNSJPz2vmnlY4I3WrNOL6myZS+3N+jrcGDW2whihoiEM4ebAxQnvAjHU
V237MJ9biQnyG6ajwbeI3TlKDlx225VN9zeEFLWSwzQX6SSRN1Lc348d7l5u8dDnsoBi9y1B07xt
ekMsSmC+fpSXLWgnWWGtu95UkVrZUfG0VrsJy2iNg1FlSZpGDBVWSzAKtFgJmfFcO2ANks797S0s
d22N/mF+DVBc/8n3/ox29ghJG9G7NhBOMZfcilPflnpJoVboYvBCUdSrviU/wgEiVZ+r7Y7d2Tb7
8gF4cxVb+mS11RvwL1hgw977AG9r+hlhcWh5A62Ajujqn+vTDHbbBd4atTBhK61DigRGycGnraoX
PnkKjONPhVqqN/ShewQ63U7ZZ3FexiZV77jT2SKMuI+KpWz4gQlobHDCqhaJezBIpfX/AXq9ZL5K
Yo6pi5qzxZjfPaB82tq/vSD8sOXmjYHWOguTpei7aoXQ/80RbPTAgjKeG1NbQf/WsbzIBxrqmrt+
eHm5/+cSnVED3oURAjyA0bjFhcSGKp7TpvZ0wJd7EjSOePtH5G7axFpB09Ot8IsGeKVcr1aGmNKR
+fF36VV7GoOlKP/SVXy1tlRwcX7UBWRIA3zDnh3abC721qCwrrg0/zS0q7RSQczuiDdO8+MB3tvb
VeAby71tB/jakhJPgLdGbV5WybPU59Vio9N4GHXy7jkhQS0e5DJkIz30BuiA8H+GKFZK0oiDaIt7
VTh030lBqtR7EJ+3e0t9addozFA2mCOZPk+azcdK8+t/Hl0jWGfymt3hZHJKI+9SyVgrY6odCPKD
zCrN8L6FwkjC57bTf7/hDA7s+fUktkhVJ+e8UItXXVOaH1QWgo2fJmB5PoIW0tlaBLv9uEHbelAZ
klougdn2NL3RShas0IANLplUZS3AufUU7qXwVLdfixwywuwpYpO+1WUsqe+6GvQG+KIP4vFr+5HF
nHkYkPzwpjdoOz0AtSiMZpkqNG8j3vMpyF6IzYowhoAIBetnmZwitgs7z3SSixvYzCa+Gwg6Ockq
DZ9fP0+ubpLMGL5kI9rJPa9HmAKNZz+85/b9+JYIFjwVM96pwu+FGPF3wYCMgi7mEPCbKDrDJ0UR
mrA+tEr6MHxX83ZusZlK3lnPgRlvKxznkLFf6/x4i5QWUw8ElxvIcs3D2t90any5tx+2vWWliZ/l
gcMIIA3a2JB+A/XAkp0YAzoBDlLU89/i7Q03PTtEJwOOejQkXpkauo3CkJx5EfLLLQ1q3O2MiCYg
gzi9+kRrtOGiZmt0fefSSS8F1OenNk31sAORlHattomPMJyZP8ZJVfnBTps5awX0s9iuhhbnICjS
W/1YS6nrwvz3lDhNw1xmyXkkYUAQXedSn3Vo6py3yIMFt5ZU68Yl0uLNQ7IWomZiARwbrjSqPPRX
15gqQj9zrD0U6qJhob8SQIqLGZsGlXuZq3ag4BPCh1CJP8Cdi/MTXlH1+cIY3r64QOmcSfHBySkq
ZOD2IU89sLJVIB7AHUiq8g1rJVK47sg2spTbBp+IO+XSmUA4cajC2qi7kn9D6CNeaWdhzFNLdZPi
G/nOTV5a8FRu1RmiwqixL2fWL0F+tXFfYEkGXVUHhOFzQFA2nqUdoWGHU4bIkmcXiPDHSdmEe7js
IpeEqzx4rQeumMFXsSmWMMfniv/BZtR6gaTSELbdUH6SEJeEY4Ty8obo+RC4NRuC692rUfQezFgJ
d6g7ksJkEfi6HGFFvSGYDnlBcAqFwJnZR/kBJsfqzwsxFATFf+nc7MjlErRsxuEGC0Fh5JQwdpuW
SmMauGvEJne04KDxOqVkXjG24vLLWRF8dGMOEEUwC5e2Kn/zMDJwItYdAc+V5QZRAqg34H64loo7
1e60E4FioUdAiFffQO/EdjH/zmiFTNKVVsq1+LzGbTPY+MByn/Fux9cLRa40nCg4j9CJ7dvBSGw/
r9zW2jK4nofyQF3Xmop4AeR986CR4AmrzY0pz0MxaLaf8Dg6u87tCjsrHtkRl/aQVVHqt8pR89zs
EsBjUWNWZQkm7e8r0lTdTaXD9+Jp0XJk6hJU6ff58i21EemSw95fG+j3rzzEB8ORjf4OdOs0yz0Z
Qv5AMeQqH2DL7EZ1Rzzry0WHq+DhROvMRX5B8Cdfn0RUV5TpS2fIWiEx2khu2rZ9/S75P8xLh3HT
1FAGSPNE362i1KS7klFV1lToJRWZtAcBuwZd+MKfYV/RdWaAWC09rSck7RVcg5dGQJBSEjHcNeeM
brXA7Be/Oh+ALWDLBeTuIT1fpJiIemdS9g10660uTxAcg38XGo9Gi6oFfgjSiX9YiTAXgTLHXJGK
yxCgwY/3wWPl9JKgqGfUqnt1c6P2RTc8e+5CEJa4hhRs5UqAuf0aaX+wXH10AipsOQrzXUtn05Gc
+YmQvvCuFQgDV3YhkdfaepvJgvt11lCzHpJAVCjly5Ja/8xPiZ04QFw6XYRGc9/jyuW323NirLUZ
2vPBZWREQBgYJC3WEevv3dVuS7xuS3GEAQxpUkvBU96sKagPxv+AtKO1TzfZOXUjehDSDxGzigFn
CEnDdlV2DaR9cCEnVQis2B8FA+hSofHLyTFD8Mt+pa6lLQBdCFKwXZZeurtc7zTPBddgCfXW8JkI
Iq4YqYvhcz2vAXbHAjWZjuWqEeg6V/sVoI4A+RIcagXDowaRuErKafQkjDC8Yw6raj4UOFZKDFBx
m3nhH9FDZ6E8vUI7xr2X0YqgsCei0rUbnOfkqxZavrOknWpv0sShwSH1JEHOMy8PaRYlQZMi9dmC
LMIAQjKgBMpf/dF+GexEGbWv3XheSyC0pIIBpTv/2zB9e41LFNSdOdt2lpVkCV7BHG9JI+gpcTcl
BmFb/2/I+9TfayDUwXJLXmh2iUiqBinjXcVGJ2F1e83v8vXP2I8OhpbnKTpjcDdRkWak8RcwXouY
DaDEzlX2/d+2CyHFIPA5cpEqm60WolvlWPdoEhWO3M/l4qBN5A/JvWbmLFBfCBd2Pi+sMJLDoybi
INxGlasuPhkEnVSGKwCKE7bOqNw8ib7yP3RnB+Teq2tNLpf8VGNFPUEzz+YbjLX37UCNOEKAXUsn
eCgdXlM4KupKI4wKSG/wfMXqsyX/CKqur0F5RTXUvMLnirUYmnhIfJ1igppcgAbVyTJuSlnR5fJZ
hto6XZX8+Q1pTw8zS6E9lJaOuXS90Kg2SWRdV1ilkwPF2vk8y+gmip+1+xlAuzvgo0PPtI08HuS6
YjvTzAUqJkta6BqQ6kPcspecNadkQtacL6Y2Tfmedu6OZz/x2+Ba0ym1ST20t6vcInWTF0r6jOMx
3wGhcC0q2+lYP7+OHgoQ5irn8/y2KtLQzNbAq7qUM9weHqrdOSPxNQmVih2fXL0yH8iPPS3/GAam
pojq9sXS7vYFhRPxGNTmYwKEqH7FrnBJfboQS08YRU5dihtLAp8yDcag7D8DA4VpoNb2spWsYx68
5cJ1NtTFW06pZPNrPZIfYaZPlayIDhu6/VkLJ5/xdNcbXvV+Xv8vmrjt3vos85bhEMrn8lKHQ5sf
1tt3SlDf0ADk2Pee0zllA9CrvSIe1klGjcCK+NJgykJlvvUHzzgBYIwieREX4YNeZ5Yv6RW1S7xl
UwoZKt/PgWED7O6XCiWimaSphB/JdYEwo9t+SJbxnQ78usgNEcmGkUUWIqfeNw1047ecwLqjB9VQ
OlC1b0vukoVMbKQy0RvlvOB0IYXHYlUWv0O7Sm2Tq4cXmulGQ2003wf7/CtXaqciv5zp2YUyIuzw
M5KQ8PKV6EBxVdQwXGTEIVDuz957piAuQIpb1asP7AitJWh6q6HL24q4VlB2LjJQvck1gvbbjB1T
gKYccz75MzVRPwqMbURdhXyBsJn7JErJ2tUR2EWgF8Q85d1DBnzqzp7XmvoUB2HMCREczxJCGJRC
cRUQYb/Z1rjMStdUB4QXyYa3eixgz7/H9MqvWBPkVNEhRpqPmPRgkpem3D4Pof7et1ByzQPmv7HF
bu1KKAewfHNhq39CCx9zf0MyOuGHhY6tdhRfUTU/vM5VD6OSvCKH0cCKQtJu8/sQRUVv7WKU3Z2J
5hmxc9JvWFMs1ocqZqtwVhWdq/KDphf5nQAYDxJbvqj8RVA1dN02RXA1dNwDVukPA1n/NP+NVOMG
HBwtdIudLKz7jTAg1Y3W0Kzt+27kBCJ/kln20EAEqam25EOmffhwo9uxp6a76iRsj3Rp4nWsSKIh
pNzEG/ibbB8QYPu7ZA/KY56vLDbMgsuTpuP15JaGvlrjjNZWpbPM2wQNaQjLh60vB36CzbcTonGV
R7Jp618VcodWbAKSHf5QMoNKl+hL/uQ2Pr7mgtAjvrxQ3Ahp39Loa2u2FynxOSIKmthpsgULUQGv
bvLURKZxVJscu666HGWedH8FYye6NRMDeus9DfGaUkzXPcERTRx0dLpKur49d+Cl/x8U63Zxcdiv
+TVvUVZjYy//NCI2Fr4LmvljEr7gMFlFVnVgWIQGtxDK5jPJoDXbBlLrFOE1TSgmgd89aYka+D1w
FoTH1dTB9+DYdtmnaSc+KOzttJbD/kqLxJA9amUIT2B/qOLAqA4NMXz1I+QqG+M1B2ZyWQE5+TR6
skqqJrYocY0DLJFfjAeEY8uyb0gF7sEG6V5U/UK1M6Y1gQylnHGFDTHnXe7PsHcg12yfctD2b4YE
gHIeDLQpqqOd3Zsizw5qeEL+OkJiiUe7eO+qE/mOQwP8WfC4FUqCjTVpE8vPRgeeGzBFZtZ3oEKd
5XOB/2XLoBfwwOqrQ+qdrRseAqHhfysMWgdRIIPHgK3m+PqB7fx6POkWx789OE1FBHWMX8b7wiFl
cDvPCxdf3cqjVvJjkzp9u3LY75h3h93QPogmoU19lxbgj6mAsI5jRGWrQhYSBYMbpS8buLQN6vmw
TxN7kaaUX+GUjDEQrAwvc+o+Q/zHvdlm49cIyohBZb4o6mwVTlrI9zJhx5L06DZr5CxQ+xR+s1BY
w6eUBVFbPf84FPJ0yDYQQhskVBcJtiHuW5YXj7ksDu2csrg2nliuvwFSSLwxXazkYRXStuQQMLZy
q0yDEnGc/l/X7WWJFL5TndsbbMxYgetN6SU1q923flWbRMsPsOzpHzVq3cKSJ112FMFOD2X+Yw3s
Zzg8D1WZK4txXX4EUdp0iGmv7i6pD7IQ7OU2Bj760cSElW3XG2vDb7X/DksQv5GV6bOc//rb/q9N
jRAheFZjw0zmMPbrhNDlL3n43LNOkQ5F5RJoCnzruL9tP4JhWG8upWs8wSBvO1DUxtIciLdiA1JR
xYranwEceLvRUW0ojoAd4OPqGG6YOmZPbm2iyi4txfeBcpzluIaziPwypZOQlMqpcLqz60xe6XN+
log+sScleDlQIWYgtngvDcpDffpohdoRe2bHr18da8m9PMIsJ+nvXo8WFDl9xu3K/locgLYyl7ex
XaTdWVATMSOrpvAa0V4tOT4OmND47VdFXdbFcEQf9VctGj73P8Xm/ry0Mb9eogTh4FXUC/VMrL/x
a8JEobbeUKM/XrHL6jCS/Sd2+AePUuo7/+trJv+qVOhZVXggl4r46GrEPWpTCf8cQrixJPvMh8eZ
w1Bz5aCjXfqyfNmzBK4NaF5+KX4W/cjFwiJ/XZaljVFxH1iNN0tsTMfiuNh5NnfZAkkPAZDGc89V
uTY1WutCZh0TsbYkEtqHKDZ6BBcT6FyUsylu50aIZepb2k9nimIwrVaPcW/Mq8MTS4ivwvsoT/Nh
2Ug5wLO5Ia+OqBXZtRfdMWqqfqKCK0kdwkhaAkXD6Ypv9V5uz2AoLm3/waMHSmBrQ5i1IX9gIRsW
DeTrsmP747YG7yOeBnnPlcFWQhuC3NrHI8hfYgqjn9ZefIqlyMJlHN064pU76vUWj4UK0s0cGtSR
i915Tx5lp/AoneB4S+kaPvCbl6jbzwMzLpoZv9z/t3a/cwsC7b9m/QvaVCl96CjmNn3tJqNjOd6P
s8uOLu6pTedlX5q4mO6aAjmAT6nIaLLk0q2RXqKi9rgWM8KjzhUTzf+15rqPwaHEovaKTpcG8HtG
QV1Y7P5uWCJ87mwoJkKzKHfqQ2czBBF3pXjm3LPyZl/r/jSXP91cAGwty0GrSz8r+X1Ntz6Y8JRK
8jNZBj02MMrSvmm1NCl0wWj/0yn+y258qdMhFfR2L/1SAkDh4gXC8VHV0mjnSpBULjEi7rDrwl/8
NHdb7EjVOezRJKVAt5gXnlJrGVHC5+edggbeQopshNAlLthQk15FYjPwLKig1aaqsr4TI+SihmvC
ZwQbdOq7JIeeJz4sDP6is9Qwc465wx4cUJteZJCpYP6eJFmgAAZINNTfWPwCGpSNcVyffTa8XFuG
DiGZUs6WbL/S/P8q1sNQErspU2dAQsCrIGnvjW4JTOYCGG5+Qth1XddS5Yu6uHTuJizUeHxdzM2V
nhSq9kvVC+8/R/+djVMJvsoobmtAv4LcSO5Xbz/kCxywOPz1oxX7ebzGPzFJ8wJH80clYoMTHk4m
AkJc0SvqTOfN8WtEm83TqypMXjlLasB1Yxw3p+YcF9chhZDPwWYt4D+U28rNHyvq9RyAQ0b+o6Cx
4dpW5Q3gKmU0Tv1nMH+UIASW+NlMJ4MgUQ8WtE4ZVIuq4qBAOHWcgVjWIuO1kR34Ufs/FgOWtZEf
Ll//aJ/cuF12fcC43PTtxy2km7meXr09Jq87qIWaLCX/wp2xttfLocei8LBU6ULziK9+SA8SZ8cQ
hFXU6sLOUXuF6x8x3aH93wKt7AEpPaHyTtdKRAnBj1P0vPT4yLpMBqmvDpNg6sldXLsljW6LQnLo
t+v5+HGKqDNxC87Ldr550fKdnkOsv5wxjZcH+PwG/aQT09DAGXuC8lKpvTGxgCmZV9SAe6H2uNHx
eUgOGAdJQCgBUnR6IiVeOGWZumZY1vXsLsHwAedtvAIS0f9rI7x5a12MPNmgBOsxs1haJBDJXxm8
GrM0eC3VZ1FNcxvTrmDB6vt3pLDOhkGrOfWKsxM5hN6d/GNvtS7+WF4aApDdmRtuN1LUwTYBdMKn
hSjwyJjlx7fWUaS+KHqn+gNwDUI8ihUxns7DzUD+2H1+mtvjN7+iQChxsEVZqxmozOnUnudLDQlW
f7k1zSGggSpwxWrWikoaxiTn5p+XF2vtFFOzxjMd2l6ErkdLy+0jeuNq/WXj/eu7r5hQ721FyP3h
qWxjTgtE5SmhCvMRD7Q9HkDHMCfBqsc1cfkQGiWQOq4GAfdI3ZA9cfsEeRjz3tDyNuPkN0NRapNK
KJG/ALs+ww5A6jdIhyH7EBNA+IPMXEnAGXxzkyNrSJ1l2NRJouGhLbS2w6ynq9kx8JkaM7hTqpTC
vC+cS6zu8v3r5VvdxzLQ6CSqbgzZ7o3esrXeNu2sOmdlMxHvIPFSNR8nsnSU2zroMshGBvifDSNg
KTCdBxkcr6UT3hWhDSdmorEnkurp6wB5escBzp5nOlsEt7NItUGU3glxZbMx9N4kgV4ydy37OY7q
XaUQCwinsESM8A6BGstvLZYd/K1AeBJrgMLnDXHSwIiSuKT4RufRWM5f/6Oomf7UwTl6lR2tSwEf
4bDANHerlgPbJcT4B/OK1iXq5yPgQqZc0f1t58kr8ht5TqD+Qhcm/2/OAVC7eAGGfzeQM0WzDjBo
V+F01dr5M2wB59oWjGATb1P4m6eZ1GfhkWxrpUrdg6zxqeZ0l4PX7IfgYS14n3UWhB7frt1dtl1L
deGrGegKYhXBrxFoZ06V/7E9wEUMJvnRq/LbMlRYWm5eGleWLwVzDni7Fo8bs+z9ChD2e4ZCvFRa
/uojPzmp8KeMNNVGqt40fi6RBwlN1rE/80oJ4hJOd0d8iGTSJyRTfv4dckOO5NuKMW8PN9XHPfi2
nSzVl61TgTmdR95p2KLj7TqREPvwp6qx+UpC68r/kiUg6RSTIRgjSyr/tO+Ma3o8NUt7wfsXcGuZ
4C5kcx5sTcy5v4BiPb8JixQxs66kliGc3hQLaotJVpRWH6JCsUbfPtWQIIpWNXwjKR08LSg9Aa6i
7svmgPiAiNL6EgJIurudVZcBzB2Wgfgp/2xa46UCtxuOwpjG9njD8iBlePYAFpP9eAEkU30AYlda
Alb8KUU1T1/kQPXlOcrXZ5PsNFBRNIrpbmyQQAQ9nc5UqIKwn9Rd+wwPdDerlaLlv1M7EJhePj8E
yogRpw8Kj6kz25exiy47kF786Zu3oVoXIQ4gLJ6S7pAebWHd1DVAiFjS1qIwLNm6NvdWqsjhav29
Pz4GqmqEN2r8ICbLfuLBVpPlaNueIqOIFNFIoJ8CYWmV6jbnkRWBtNeTnOJAy77JUd+3uTZ+GVjz
t7iZk1UdW1U1pnAeLe4MvBQhDrTJnIoa43AxTvhK1W1oAuS9pRLvExPcYFfUUTNfTl1PTRMXi87/
WH5G7Qyo10ExWgtnnEw4f2L2bC43ecvNPK+2LUaf4fGSWBGcWrBytrgHc+MuyVpT07KyBgvIsaxC
aULRyvPrbeqQ8F5oeZdbKchdVNWsRjT2iRsFh0DvRzPyy6Q5x4bvpZFszYKghaS8MwYbXLNGhr2h
LQMPOxLM87kaZ+GLgFZJJkBKysCJXtNnwncSL8jifZnGGdO4pjxgAinSmueYtGgVbB/ORrK+sJHu
e/BS6ek1FUmZsXymLTXSuJJTXUdRqclveazsRyqAwhYCR/GL9AIS9mbKFy6SQD9vrJXqM2p/8QGi
VPCKyLYZ5ZdWUPTgkVfDwjZsicmj8kgSdbxe+LDFe2fFocFp+rDhLRz5i3BVFF8Dm9mmf+FtujSh
DeMVy7wimskaIcXWW8nK2xvkb2pONkIFapOPbySwiRtF84PywhJnB1SXQKk7jmKPX7FcsrLj1shs
bzrXeEoWoZSPoxv/lFEPCWe9nG6UJcSgRAb0IVP6HuhxEUx//BCgRfTYuwj+ndLXfHQGgHz9kZFH
8sa1DjgZUsBPtIb+lzedvRymH1x+dUXGmY8zMQ5ncX4B2pyvt6JAKyruGWS9NCUNtYUaWE2M8tKd
/guVSSDO4gEeAWNvY431GtPNFXn6iE/kZpXHZj/5/zem8lKKKFRYy9U1lQ5eFvVmjUuft69blYN4
E5XoTTCYiGjI9fFdctMvx/8nJjutqXVSta2UsWJOrKtwuRZ4nwBPimZq1AizAmE4xAcsxbxCPRz2
olcE+VFTvM7jglgH0EwRHm+8KZS8u3/nFg8h8eTVBzaEJXwW/GPn606YNZgY2+KyGeYYub8NzK0F
uZ8UQwvjkRCD8Y+5NEbd7CCRRvjsnR4iqxQUgGuQzp3I0fjvvieIdpRLNRsjx05qutoArA/Xn+Qt
pLzlyFpSb7T+BYGZa6+6cQJKHQ0vZIqCQhBUU/YvlryBa/cx6Hfq5AvN7wdWz9MeijF/7/1jpNIt
WMgGkvv5vIybaZb0Dm+rlB7GvOr6HFPicvVNFjz96kRIRZONPKtaAgdGH+q+XplWeR0JAAattY5N
X5dKm1wxrrjWM4VPRjpA5cBSIxRmxaNDJY+2arLXKIerW9b5dZkjSVi5GH0h1njkYQFj8GizJzrL
2Owr5s/L/hiGMO5DuDK7oJ8pLWGuPAszM+rYLUea4lDwKZrgSnWviLtlbCMOmJ6GKQggnP9bdxxe
b8XEFlQ8r5Ck9Mkb9fVdSULutQ9qwVsWS231vwrfMtkbf7SrxZVMeo4OYp00lUnk3oIX8I/saV4Z
r7T9tfc1E/v0skeijsHC581/XJ4wYuyKVS11A8kORli0P2pxhkUf3pyDZEh9BYf4Y70tPgDKjoGz
tfxB+VV717k9SxXEcND1GVxpM0cpU9YQeRYci22dTnayoO37OsV4Kw3Y97aTe5bMFMNKOooDiWhX
2iCZjDZU+TrLttDrHb4xxvXBV4SH8haIPuW1D8+8UeTEcYriicenybJAl7TLe9gCDbHAieglE22d
KQaZPI2/0Xm4ezXU6YN1tUYpqZWxG/oJu6MeskE7NZeaF97WY+6KhtL4aVkunUT3/HjITm1cFbBk
Gys4kJD7U9jLtOAY40nZ5XbcKFoa13x4bNL4XjXx5WjlfF/qNEQ2IRdPf2Izt/UqyrribOpn4fFf
EoMq7SHdxmMynEYMREFM27kDtc3m9LXOhYkwpHWKPfDP01QcRuD/mg84lH/fPviQ1R2rSIb3wT7G
JhSz51t4PE+TsqsckNSk+EM7/BnTFwfKPU/Po7uu6orPUH1KnpTgNa27s18TYYCgV/U2HLIb1oiv
eySPFFzhRwRq0TC7zqYtSCgfhG53vUUyq0D8j1ldT1yzQU2H3+JgAEzqnEeyAiGrzwydMNEWvIco
SGgCyR+EBlHa+YSos5aPPUlCFp6XuF+7xLUzvXHPneiJuOd44OQunZJb+fbLKQLJkyxNqIpGBHlk
mfylVFMQJ+EtcW+DWTFvVBejXtnSATZz+Ds6H0LsSO360qRsh4HNSmRXoY4RR9hxuz2ck2Gss/RQ
rLE05GzPEfgEWZC9aSVJ0BReio6P97hsQQFVIWIsQgL+LkAfY5J5AHTU3sfySgFnfu21mFNywok0
/G9XqXmC/MqwrgnHBiXeMIm/l0VyLk0lrxIz2g4hYYw7BPyxKUkFtn76bAPtKVgoaka3nk/pXp4S
eyT4ewMfGQwfAX8I2pN7Vv/lfxBtMFUimq0I3J/zbqy72sAdCgq0ToCKWrsN7K3OdsjhZdBZXpZS
aula1bBSSn0X/S4fgkPT/9nvYYsA2cDppCODhxr1abXodtNaqHpjgDWOaxEafOnfvRv4A9Urupxl
VrVkgbynhZIyFkIeNzMWm9CfPSI/oDgz3INXnppuQMWGJrJPwdQx4wQIKoK9CMN1drEU5iFw8jHO
CrF9Chun5+qsU2f6fdl8um+VlRnlAd+4Bk72m/pcjukn53+j5GTa5uvMVyNI+SUvVC4MtTNjUujC
IhtV19qiAcWyDWUTYTVQo7TsuPglTcMmzdMk8VFm1fLMcPwLV+yEx2ZhPMzK6MgXpUSF9oVTIzhS
T5ooW1eC7Yne2S4SZxBpZ0hfjkOFszPb13ij1yrQ9MtHly0yBESlHUFMbru05gN32tvB0unNfWWB
wo8J5j3hITZMglZC8XTNPWCGhLQSsx9xaqnZv31gycFLNwC2tHztTW5xg665cFWznUgkFU00V6Xr
RfGZ+PihqTHSIk60ZuAlMtPcgPY2dK585uIkvErwFp9c5G7f4VA2eG1gLv3H8eHf/SsbeMKXvqPx
QyFLVsXpBCyKsyfP4wIfYaicSK89Pnf7SAnaohedCucVh7ieQrRTmsZvHAAsyWWEmxo3LWyYGDkP
iGGaEP4urjJ0bNuXH6woGZNJnqEPwD5xlZIcGiH8A46pJBgFut3t08M+IhUe7FevztbM9bf3a5/G
YV6OFzKaWEToov40hH/G0bqFLY9bxj+n1vaqRyPZ9BEbTyV8LHTZvUdJT+LO/MRLdXwSE9meqxrF
7fM35Z3/dXJDpYQ9WS0fyRIRsS1wtUe2ZEDQD8L0vg7134K/iW/DMDf8y4SpYFDp9e+jBrfb+uZl
M8+Mx3/hNm+fbBv+he6T09jPn4apYm5GjKAsxvmuOv8xgr1wU7BVA9dglyCa91qZnh2UkqF5uIqS
63X+1w4HEwQu++3tYLeMzGZUX0Rk/29EAzOCkNfNpBhNGpd6GvY966MShYNbHojQF6Dq2VxOcteG
iam+9j+APICddaomoZYlbRsrA/p/AspurPCj5ZOzwzZR5qTohP9TrcJ9C8SgE8UX2moQiB24Q1HT
mOCdz2YGW3kvkp6fUO+NhLze4L3Ny3FGsCLXNfnw0FRn2swbbGOZmoXKmCjgmjQI7UUS/7Mu+Mha
NQh/2jW832/Qm5rDr+ukEufq8g/7mqwpFU8KK3B4Ct1HMIWEe5UI0AxIr4onbkn3uy8EykIoVcVV
d7TJ2Xa54dhdzBs6uSSnmEiWVPeC9VGSJKwYnyKOO+KSdWSpvpLLF3sk7p44lGmbcFt85YF3i9IC
lieJlYFNQKYq7V5TBZc92QYdX8Ix8CY8OYXist7I7lBFA1A1EF2vkPoAtfU45OU7RM5A76YXv8rC
kfroK5/SoDfAYbewF0Z1YW+f4BP8aJ6kCROhk/7jjXEOZiv2ufvSJ3Ky42xKDYwr3Op0vePABm6U
ITqJVzrtvMPbo+cdoP8aECF2XJ2i8nRAOO73gKlLxOd2Wz0HgL+ULqEWRC6S7Atg7r3X17CTCoHe
mR7oiFECdYQM3qvsmWD9FelMaynYXWBLkk1NiTGBdEZp3gdCjyaE9lVEgslMoqWnn3/YkHdilQxi
Te1XbU53s10kGEdg4HSXKc8TP8iq0ctF6pp51BggMycxN/ug7472ZM4d8gSyY5l8PB6NqDJ2M1zs
MIYkH6XqRWY1BOtBe1B6a5NkYa+FgZ7jqGlnmjbAHIx54DMCMZ9wvRbWACSwfCD2K42LAmZ+CxbM
20b3oK2eJ49g04g2+k6xqmqFWPFrh8qvteU+LJ51FX92U1ngpv2+yQDXNb/fpfWoCQW017V8VJDw
E4Zj3DYW69QocvOJra70DlnFl2W2C8gS4FAXOkqg0/17BfRXPK7PfCzn4j5/G/I7ooEm2DK97bnt
ze3r/2HtLjDFXY729ggXfZtLVk7xLMxWLJmU4HHUwXyPPYzRg9mlYQUFHkUvKgTC2N4O2LnSInAv
N1wYweu9jLzXKEJHqVyeCbuzbN+7Rgdkn/eboQ05D2jxmFs494e7iWyz2p8WMr1cO0TSoGWxiCEF
8GpDPOvvFhzBuTebuvfv8FV+NQFvpqsgnj1haPew73qrgtdoRdpqjraqPzX5w1DvW++rMk9FSh5A
MHCNVLsl/0LAgwOE0rmNRQMav36v9ghH0x9iLI+JIG2T4Y4EzNUgvRcokP3qRqhz59pJfwa2k58n
oYAKTGjGpDu6NxSrfNWIXhrAlCTd+CnnvAiwRSyBnx2KjZEikvL+WmuSBJoYjttawH+PM0rD3fYL
/xTGOsjcRZ85uuKqrq7aYeVCL0ZVP4yjFKSZtShpZWliWDRbAwGKjQo05WdG6M1MRIEm+eyBJa9s
UIqjQ0veV1QkkZgS4TXCGDx0XHHaCeL3SOqT/CbHFoY/KqbLLBgDmbAmNbF6cK1HcOoVmN81SX45
Q+Wc+cG2XveFHFWrzGS5Td4xAY7bdaFGLu5qChja+EaTBy4cAU47KYEq3jqoA2J9EO1MwU70vZev
2D0cateionstbZLUXukBvlJ9pVvV/4fJnWBya/dnx9s+vh+CIQka/bc95DB4hkOuRQKsKBgUuAGJ
k8dCq7UfoNYqNoQMEDIpBh1tFn71/b17w6+EfpzARKbdAHCLmCfzwtcgCxhCI65WqWfonO9+95NV
xjVwZSW6Zmj63V39NRFGoqOt7EOTpg+A4JNfVAl4oV763SWWoaeag+yRZ0Hu/Wd+TNXHJZZgptan
kVWOj7Hu69Q0RrhU+udXZyE4NwGSK8gIuY5lY5Dz9yAxt9PTi1/MkMoHhgk6tZkQ8J6ypD5WsI1h
0Cy1Uc8mYDvpJKrUnrAG/RdT1/1ZzUNhFe7WBnNpEqvUwqF7QlK4nkT+R6xLSgIV/JNPGwDVFjjF
nhTm0PvDJ/zgSxYl0esyI7qMThczvScIvYfOvF97INP9EjY3aH39KehWG1eV8F6iOuHDjfoCH4bg
rNlj4H2uPC0PvTYX+3FKB3RFAQL7soq5gjh/jDSavAaFo3zG5L7SGHFx4PUBoKBdwCfg5UiCNACK
+u/xXAFFXqT1gelq0elqtSVKiD524YRzMLxt+6plcSo6jADebO9LKlqd0MZA8Ysdb/B4SO+u8SwT
WrZsNNTIS5w7YHBXIkjQi53EOjbYmy2fS77m49SHZSy00nPKSKyCTSR2S9zT324egJzSiuzUBJdi
gD9SKF7YvNP2mNXvIHRYBgHhK8YFNOamm/eXB5yY8vivgvIMeUuVkWsFOi7xUNmOFf9QC+2cnV0A
XFinB07M8MHyOReOHeX7dz8WgPoJq+GKsoBkPGbh1zN70MwZBA5kap3YbYlw6c8hMTpkZylv7CRU
wJNrRIcG4itXAO4OWMxb/2wbgr+mCQm+vIBMqOD/w526FVaPtvJhLTcoy1yT5yQ2X3bmuPemNmaX
0GADrFTx33Rvx+9/OsGz01bm99TlBe0RJtn3Nbf4jnn6isA+jAWfC27ielN8jNIKKVBmhvu9L60b
1LF9euW8ObIz7+5HzibxRPme27SA8pfR9AxTIlXEiU3wW7TqhfBVuo++ZVEcomBjjn02kDYxmvty
AcR1Fm56KypWlQMQ1UHXIzaJErmsOX1k9MuVmAiIi8VkCd9bKYDtq7b5xdIgRPXg/2touByu6Cs0
Ej+BNUyRiymVFGv4jvXJeQowFzmOnTVxzCW1kE1yKYruImwIFUjPr4ELlsGrX5AUvqOScxW8UtCD
Rce2yAbSdDW8xRElV0JSiURobRI5gJaUGvIq7KbMJ9saRqIRquP54A6NH2ldEjP0sF0uWBz9N/IJ
iEiNKcTWq0f6LvyRfjPLZoBuJnbVAWd+Xk5sh8VancG2HHPbH3Y5gDq5/KTdoeNlhg6g61xrcpvL
nkX/r1tcrY4314X61h0l+KMj/UeZiFScUEUVVgU+mgZQO+f6AxAApAt/0OeV7k/PQeYqAuyqW8Ns
N6tha6nZc463kN3HlikoZKuZXNoaAjdC/QBRiRaoX3UBPP0/07brIMO6ypcJjC/7MCcj9sf3Zz3k
GaY56u+rkiax6ks1HYAONEfucFLLJ7YwW4OxY9hnRkz1osTBU4/sVlUaBjKnWVmSw95MLE9yNgTE
GZmQsstAStXagwLa+gs0udNDRFJ6TSddLrxdf/IeWfZIL9tgLqKj4xsUsrQpoTpFBcdjmFjORnID
iu1mg1qtD6TYRTHGrra4r6701sH25024Hq30ixT0QQkHYR/bpo02R4qDckVwGC8psAjB5S0L9n4i
OkPC0ZycEDlP5pnNbyhF6JNd0Y2WAUyNsqjWotpJmHtEQj1+9aq7n3eTP27Fs118PdXITJKl3NrB
B8lM+rXNgq0SKdVHKC28uP3LIRH61QWoJiG2YUtqIu6Mn79GnM1DtQpjw8nfCEjUUj0z7V+wbFCr
E65jW88Bd4txprezx39F74vfHkK4oFjgyK+jhlobNj9BCeldexh4qfMWmwsFQsYGDYpPOvkADmNJ
+tBjriaxWh8Cq2EcvMo2df6N2gultF9khad+xQOnXWcIEvCF/STOMczJRuQU12nMc0s79xZNh2j+
XyOi52LWuJ7ZhQvzkWUdvoH631loVyDWy6uylCNFC1Unj9AD3lE80iFJNuIR+8RNX70pA0PLlwjS
eX4MJJDDO9DEYuI8LcvdQQXq0Uf/cOWbB0xXoHJBZhbUkkTxZYje5nGBGZDJmRyU5D6CnqTC0M/z
yrYUJrRzUnyvSNnBWMnc9DUM0lG/eCHGqteNPydtwYCSrh9MtyDhph7PlP2ME/8BikKoJiqnlRbq
ffWMRc1gxA52OVQkREheXHTFpSJznQtxQ/w5rRw8pzkfnFrDGSixycBsHlskGRqYh7c5ICb9RYrD
nVbjVZFsQRr7Ibv2Wt5UVLqxC+L9Cz3Tmo71lV0EEMOGH/xxvewHkRZAoAXI9rXddKMT+3UdSDD6
0jDo5y/kpsvd8x/O4O6UfRPSMhOISMK4U/R4brkuyMDYfrcETDSozqoOwFTeQ5uIlYXuY8vDi06Z
dj/qFlFN4j0yX0I/NQAZQqaiuNyUzJNJj9QREFzK5U/5NpQaQTVTmn/T2jpm4VH5EzpTXA4aJILI
qN+79ME2K+FN+Uza+e2OEZC8Izyi4FEg6pPRjIVXXmqtA0riQprs+Cmo7F3CSPnWWKknoHUmuQoz
xVww+9WRVd7Rf8xPhSzead2/q+RN6SPySGC5WOviqBQRxBZj2tJWozHyG6xW8Br0OIYd9TuGHlE0
MoWHwPmfZBwpYgad3i9Dpx/8mfFaddHu/IorF7SMCJp7lVQ3nCkWDYO7/wL2dFD26kXehMb/CqEt
zLLVX9dNXNETbrhnB99sVdFQEJxswRQix1rG1SP8uJN0OZEbNL9I1wzy6hpOmJArDlgWmkwjPv13
phqRHe2sh2YqmO9Ixv18vkNCeEyVLHeOkn4IeNYC+pkMukefZHXpdr3+QUGk/DfS53xYTPOOdEtL
1sEKOXN5xXqOqI1Xo8b3SOjTW3aFlovf/JeQWVXQZdniSPiRSatnf3sqYj4Yx9zS/mYMGDT/dz58
fSALkiHAmgzRlFPb0sgNUlGgW0B0gn1rJ7/xDycmLIKIF1hi87gQ5N95fhnhoAwiL9TPIMDTHDXB
E6pkVnt7P5rf0e3CArF8pwjkGl4dV9V+iB7vAJgZUqiqXviPzXQa1zFT+u6hzv5WfY5E9YDMEDqH
AFclyhOz+6alfZtGSsPKA1emPHT3VAOPTcNdpM2hL//hMM3tTfsNcQRyXhkjzwJR6THG3oWvq89x
f1TRHjRCqJbgtegi7PZBWs+W8zpTFwQkBtZwffvPKj0NEaATr6F7DiLyegVARUfRmmercchv3BFm
e76XBXoyAncECAucbzr64bzanBIvBz0465O9x7VupmSTsfLn9GCYhNBphEp2sOdriEm3r8Dv7IPE
5Rs5lfzeiDuwiqNCIM0wzfB3tYEFpcyovIM4kBj0IzO9FNDmUVUL3xDbO+GHDIm1ZnvZz5ZOzAiv
tCT8Ddr8AZk9Dkd3knvvs1QNi6fI9orO68IBe/EQSbBjIr9muO3mY0q1Ni+C9ox12bUITvcAcJe+
o7cveQYBufDUzbov+XX8p5vmAjrpSKjofybEFESUh1s5cQbYu4c4y/4MFzS/myPqbttjR/zlciOV
jl0kNSoH5ttXvqv6g1/zFD0Pr6HTJl3KPzjOab/hsupeTmiCqSkg1TE+T3uXJNcHTks+LVk5oof1
Gu+cbjjb02PfUXAxcytzbm4edIJgU+JQR9BqUvHHPTtxpeLaKtewiu2jk+1Z4ujq//uNjUbiwc9o
dSeLnEBhMCMbSJ2dywXPnDHAJLDHwtjSE7UxmPnNlYHIHq4IE5M6hu/nkRPe3vByXPIl8lg9C8nR
afXgavVHrLqknxyDp67zBx5oxj1Ryx1l+jRh4ShDPj7FabJFfPIkAN8xmOw189xo5dZrrQJWq82s
o/oBHSaUMDtK5BKlKu3CysSKfuBIsunY3wVMIuywqn58UskF+cqf3DoaEL3+YlCbD7f3CE9vpzKe
BBSz+S7aZo8WX+hHes4IYC/Gj+xYUv/YQbWmDrbzV2/0ptQ2IXj0wrgDHIhI7Xpdgxb7N+luFdDW
HCW65hXr7BO8XTYH+iWfKNFK1hTQcsKYS5NkziY1yAE59gRf5SeXbphab6W6+33nVuV0sfThNaoN
WX1qmd+hZb02Q+SLsAt4ibjHuzMXlux3zyUAWSe5FLNK/0/JhLK8qmD9uRzzbH8ApltosXMMa0Cp
EZqbaM9o371RTjCCsdR1hvi6ZZXIWmtzB2tGjeSys8lIEQxKXBH/JCpJJt8tvDakj6afLEC1/3NA
cd8gMEPLvCCAmrfm+RWCbJ5ohPwnx3wNmkReQyHhJH6Ds2GGx3Gmb7mNrXptINaTY1dlawoQzl0X
FEMpRv3qKSxkj4tP4WuAvEu4zhgrBxfKmxWHB7ofPeITwL+V+TfyV3TJkNLLv8FVsDmYf6I32mUr
mrriG/bEZ+MzjDtClaav5ymQ+8xKu7sE65gtysa5ujujPTt5haDaVsgcTFS4jeUOUr9JqUq1z15a
UxvL0KS3Ie47GjgU2lu2sYumiL1Twnj1GAbrexhXkKWODAB2l07IlUI+WSqasLRq5e0t/H7vhgkq
f377sI1yvn0DMYLE0xbDaInycDAoTwnPg3eh/9S+InGrZV+0fjv8MuPSn5kkVPkIXSdorTSsWPnk
gqat0PQlQm74/SkROuh3EqvqFMwKDo+JFLUTLshMuOMHHLKeTuE+IRqV5QvCLZpR+Hs8aYMWqQ8Y
/tqSuZBRFitgiSWa67FC0oKcFmLLFne0t149okkKdFaiRpQg/k2TMSYCByfJ8BB0PUGFC8yLkwNj
VbJkxVdzrUOZYGQE/QAMpMDdHJ2+rMirT5pCcmfWZXB3jXHY6/Bnvs+iYe7wnpy3MWvOD0J9nDzG
vshNNbAf6sEXEMYHAolSoR/Mun2SN7iNVonLw2kSqF/vv5664s7zGEEnoXWJoASyWJMR1vHCXXkr
XyG9Bo1cl3WoXcK4hGkn+ObDWyzHyU3MBHcWsASQ/rUGYOjUtz/8pxNFMi/S2gbuRPwpR1dDQ4Xu
wz4D/zjLIAfY7dcV5qUSj/xAmfZS9T1M2QfXwHUyqwZD7M0Z41yTz9bPtpRMcW6dcfrfBfXMSZR6
UB8NOTuF1pxK3zEbvyU8x9uetrsOw2EYxxwqmVfwhZRGRESO9D6GCMnHsmHr3Mct/dxx4MOiW1HM
wKNYcsZtarRAGfoyNjZR8iSFoFmAWJRk9SdTbgpnmelup+tQbvH2j8eK5FCob7apqoexh2+M9Ony
bxEk7mRnMnDtFMBkPrRVuUwtM/Iui/kp3s3D17Wl1KMdNWbfh9agrtPFXu78OAh/QIy6+sM+jLbX
RTdRcbqBUvuD5Em2AgK77j6mjUY6YQuPmTvTqdYxRy0OEE7EU4oYXghVFkAFJEKLm7j8ftfK/5l5
647TCglt1NZUwnyfdjT2WUuoQiLI4q9bMNnKWl62e7Q/L8F/WsIdU7FfZd6R8O4TcyhmRlgKy2u7
PN8HVeROZS9S4fk+jhuvJWOrXknwpIQvvCWex22xnSIeUK4qd3xnB66nfv1XfEDt7UJyXCg8oHxW
/yEVO7B0h3MRcqhz+62760gRGe3Fh5fJd/EqWASVd9vMEyEjd6q+VgNmE28+Y5wCxw4AySIi22rb
hlFfcNeC9qJvMvmtAMXS4GDiiTlHt4kWQczTNl5rUiPI8HTfQuHdmRUIuRrQeLB5wpQnnAGCJAqJ
FMIu2ycPn01XK43tY5D5xLyESLD5I2CxUYz/jakU1gwaOdJn5fL4mUMKYhsWhImsj7NsHg2+eJof
UkBTrCoW1rN9HCkJHzxKJcOy53CypvLYDBdOP2hoGGkN3Q+R8SzwUAK7nIVFIpVNv3LQCyteCYGT
OwE5KilbcWkFQAinAF+xdeQ/BBtrFrDMz8+1KLtfQGg4mVg0vvC0CnzF4XbOD57ItRUIAx4D4QB6
jFM5Qxh2OC6L5W8fA3fwOjllxzDODJkiTrqpV0C4BeDfxyBUfHiGinUhCGKiLAcYE/ahgEqEYPjI
fu87/dBtWe4D/UFY+TryQuYmSFzDwDEaz5NcAyqkCBbtb2g7bRHPgivvIwa/zhLDjyKsB8KG/fU5
3s8+EcBwsKFd/8q2cOBwR4RbSoQRfJEZCYTSSuIgX7C4/dHbuHmYllhRNs5CxOzTQbJBGaOsop32
cIbaaoJsHj6KxGApGxVDzGUf1rIJg1PyDr2wtp4Hw2ZNRivaCli4zPMtBQfQwwzXTm3ipWFNc+Ks
Ofe9Jb+hP5i7Thdux3O8tPovmlW+xrTw4sh9dzQgzVkU76bYhp2IACQVc2VRxHsPw4Qxi0ROUsQZ
rqgfA15dRdCR2Sr6Loc8WNy692y3qAc7fG64Hy3mCWdtegMkqLGrSUSTvlg0AYhxiLL+4LkPv920
YoMoH0gDgsqB9z76xPunozwI6bW9DQJZgkVJbqXXnsiTskC4+c2gBFAe1j6UAOr9mm/QL0HHhJDp
IbWS41e9lTzMDewBqOjRGbhg+BGmvQq7CI2V74jGFTTxopEfjzW9AKvy7Wgxxkab317iaYwrZhs7
rkz+aceUImP2yHW/0M8AOy6JTjOmcNG5O5oGt+GUviYS3Fa3OHrBqOCsyQ7IZ9KnujIjZXPepKDn
rp0KLXYYIjTamNQWqFcmxLV4GolbNKpty3loZ1VnULSqImZe4XRGPDoRYz/dohmcFBr/bbFgtUM8
xFrIRrii/73rc6iGZ+mjhP9byBDLiGkbuGTk997/YmlZ8UBUvMyVVbndYorwgSk3Fec16KFa1tKx
akAA24FsqWzkynal21OHy36aAiD5Xzg9XrBq5Koxp4AjStMEoAxX2pN35SURiHOXpNZPXNSiQ+ER
XmNoNjG/+vxpwXO8PeQijrX3xNuVkEg4Bhp89Y/6t5WJWEkTWOr28eys6IH2ptVeBXxlXCDdXpzq
9rXQS1vU+Rsg1Dp7gl0eLvr0tqFdrj7c5f0jEbf5nicPExU4Si2dqWYYYG77xRfstY8fFHMJh/Rb
xf4nlbrU6mHH6G0giBqDeXeU+9Pvuvv8dVUKUnPbk3g+iOF3EPFfSSmXXIrMJDpdUBOl1a3HZvnS
o2oRm8kpb1kYZvcZ9WtVX3tkSqxQvsYFuh/tTjA98ic+VpgyjvknHUGdMibGrZv/a0KU+dJZdghu
i3uzrEZjZJwo34N8huWdP6CHA5IY69mpowlE87YuMFVL81O5F3E2KhRtkg8R9b2sAECiuNnE9pVW
NllEzahRJU194L5KOureDcBgjnQjEBmzqNX87lpwhboT36tD00ul/J4fkQaNyvbmZuBCI/Ccds37
D//Xoi/YqaCPVByFWlHkufjXmjZx171dGwnGVdZ29IEyjlcX3h0l9WSFdzCOUlXsT7YOKUUYb+nK
tXviFT6yxbIUeE0endmrSx8vmROrmlnB4mb8XYhrdTd7n+csrpCDV7kYVA0XBTVHAahWb6LI6JBe
qYSEMwRNBHJID2xv9fk8rKhM8sdt+bqExKSK+OmiP7Wps1PAo82cLiu5SD7CkHRB5SmigLO3EaG0
UWuMGyhzzUx5wfgs7uNUSVCFw4lw1KjeN2h2mffmUiK88M8LWAXbZPpwFXefj4mbMJA6IsbDjyZy
o/hbIi2+ecpHSFHwicm9+R/kqI6sSR6j6560oFv14Z2VfOuR2cu8n6mhBQqgJy9g0Ywd1A5ATdeQ
bivSh6qRQEoZvxAkmDxwI+NgOnd4xCKI2UdxYRacN7qguzLvdIUMVyhdoPJDT9BJd9J/m2dsN67t
OB/1png+wxtjagOHBl8aSQi/tdCuETPeALPr8LNntpLsvXA4+qEZYHysy63yi2QrOSsMll37TNcj
UTfPf8wifF4/DRIj2ZcOe4e/VMz40SBgKHKUloZmg/XqH8JGZAsJEAxQMX5w+tXJXh3aGo4+ucUK
pezSKoXgREydRcif3e5EzPg8ZY1T/OI8YWS8qk2RxV0KfUSY282ExMJpHzIKju/gigCV2DwwbmF+
LGMrPxNSKxn48MttXtZijYKpeFLrE/UHDEDncxASfw+a4QVoUCjx8zySn1rFj5qlgmdcewP4hFoW
LGX3+ApPCZ7CRgzkN/Ex8uHYJxvbKgN0AQh4Y9dKOYjOS+ZAadpx2B/K2u6eq9zjQiYn1RUjxgtQ
owVdGAiBHi1qn4hBLKCeABzICcj6/DxHf2wbJh3M6Sxpsmwj0pVnKOfMsOXaiRefhRfVGefTdVgJ
pMzvrIDZjBCg1CB1s6NXZOMpFfXStQNOy5IWTD3KBiGb27z1zy3wmzn6sFqje6RY96wdJw6oYQNv
CZ6WHoZmQ6+LEfu2axU8Iq35ng5ItsNdvV4fzeT0u6mDuxn4qbaJ0FrPBGqvX2nTRRcHFxU/Rq4H
mDoxCoTosjJFkTEGvhTM6CzqCJZrKVYXGyc4QXtAsT3hOjiXDz07DNftFRwB2Ry6wqy5tycZvgmv
hCF9RcN7hqcht883XvaCtO5OFpwlnhXvxYv84AiePyolF83s+k4Br2DtnpUW3lX2FahHUkCK/WhF
NLrSPwnFlx7VtgRQEeaD3A2jsoXxiJ4k1xdWwepfw2Yfqv4H7wfmdB7leBUjQ0TjOHyxVw8KgRbU
20stnRYExJ6Rdudi4OCUg0U4qPCngB0853P7Qis6A8FPoIQjHjGZR4fxpKqHHJmYjj8FoSrHD9Nq
N6a+ZIaqgB5F2k2XGEJBag21aquP41B3Nc9F5CBcAqTKvXLaaRbX2vK+WzJzSTFqMj5tq1O9A8rJ
vBYppVsGwCsGebrY16Al/+/r27K9Wcd7aRi+7ou4W+1GDIv77Av60pIcvg45AwI/OX2JTnHBhKcj
q8fAuYHbOuFjWYmMB29ZEfxTTyReExG4rDOfNFyWXXYam+8H/pYr3ljy1SbqzJt0MLqlpKYqTh8w
sS6UE4uB94N4vHime5TUMVvZgykKF19zueT5iU2WbgHt1AzqpuJGB7TU4hwKxVnwHePMF3wUHRb1
1x9mtIXbDyt0SfAAYFs4bmuipfJMm9f/IhHGiu17XKhvhiNREl4BDWOsVNwBfElfB7x1D5Z3Y5lf
iCK2f5fI2/L+YEXudvW726EA1KaV4iowd8G+oHBiZJJFOHCz581obAJI2/CIdHeSQJ3W5gSrauP3
6oeEjLDCAI7jz1bl+YRiF9kkF6cJ5HPmlCJmdcGJMOS911S0J25bCSYFFr7/3oeYv123j3JiiRoK
6mfozRmHAlEBqwx5Y3g0qvuO82H0mAthJO7sPfXYhm2SEyjNKmXcHN8MoYODEHEU3faCgCr2ccSl
SXbeXTWerqPkmnKPSOvsn2UUHuHPC2hy6UBdgEdHNfypvMCXe+JaXz2s9nmh+xNyadLFxBaD4iH1
ds6ogG+8YO0QH/WrsdY7lGl5NSD0DHMKUZSz0TOATxIDHR6oBv06uEXkx8VOvF7qtmKlj3z7JQo/
QwYeEG0iJyNx1XhfmXEUzJluXzccS6BKRLVj1yeeug/qdkuN53neq0JOPqnaAsUFXczxiW7rLTPL
xKHGdJfVMWxQTDmRYzpzw1HGj1s6OoXLkIyVN3kHSI1B+X83+IkNoJc2Fnx8NEYBxa1fYizxLZk5
0flTQdI1tOxOwHjm6LChfdlcdbAcJR8qm8uiaZI2RItUYlLkOl58q+XgKdox6KOUToWIt/rmHhfS
AX26D3bZ/RdJ0nFwOwtH/0ybocsWAohgTBJVmJBKqjyA7memZY6AkxjwOWWnWQKB+/RqU8JzQyTJ
/JQFhKRPCNQZAe8vc/psUA6uQpG3hLOuMSuuVWurHEtYMJA5dzFQ7QGE7T9BX4K2y8HOQLItTC9n
xBoggiYfoq/DnyqeJNF8C4dzvbeOn63ZI1SFuwqHqq3xZDxVvZe/5SbQlGFn5XtgcOF3LOht2IR+
qzgBSyfM+ePoRmfXmLMve6dfe5T9f+KtkD8PYjZFZ3Tv09RV3rA5kvt/wA/iFXcj7+18i5P7HbXo
g2OcAQ6zAzReozQ4pLvWnL07wWb0yu5wbSFNhZmHUFBc8FNQCvBhQ1mgNtHlWqr+oT0HIVEP1qqI
4iViGOVZUWpjsmkjFp+GcqLkKaZ4g5I2BlEGUUpIrZ1X/uqiGcXh/DZ1quQPKuJdy3FOtgMBym9n
gvnpgsoydMvI2FZBmfZ9GtWN4knAMYgDv2Dd1n5OmyC8VS3z2x2Qa7s/DA5olfj4JJ6s9ZAqAldB
0p+fM8Y1JvdmAGOV9XP48LJci637XBM6keyUI4knznTmyGL+E1bdl87n3Kc7qN/uvbhblP5BiQr1
XdgaHHPkX8areoA3QPNc7uZd5ZkA1tJJcA5ERD7uf34wGYTo0Gqi5qs/bRWaQYC+AFiL94hHIUlL
8Hp4U+9TKHaraaV5gHAGUkCOcIZBZWDAMHpCqT6avgK/zirhZQYP+C2swsCq1sRkWQY8rMbxfEoF
0Ij8A3/+LjEQSOIizonoc2EfzA0f64UiNX4jPFarsHQH4iUw10eVJndFy9yk9iZqT7E9SVf6VFzh
qxeodo3RPasfCi+11BQzA9oX/EIJ560jfRp+kHHlTjHY+UXFIWvf7rPqLmU71QM2NS/ptbRwzy2H
55LQHdiJks87paUzXk9n4rSq7j2AvAJJFMte++dBG0wo/2Ro+epXs7cRQU0KdCnSm7xPOJ+5/2rd
FDpGbcU+zfsNJr1/umCoePttvr0CfCLR5sqLNs1UQEgFMY4f/urig2U8QZX8LucQvXhf6Ejn9aHN
gtf0go3EXNhlF9iFlxNASvzmbhzUxo4SUDFcAg65GOKqQG+wxuUMjOlk+fSZvYGvcD5XoAijtFEU
daXqFe7gOlWoymg1dVLnlsgJG/tKIhjqktEsdlKTlAyZ2rV7e0lILiSQHuTzdMHlx9/s36GgmbpI
lKOuxgrRHZ03x5bxBlZYIaV2f8XJKrAHdYiEdwyNQ4d2NKqoFScUY0/fqeiSGLgaz3B07VHd+CH7
MiQB7ZpcfdDk3Bsy+P5mFMgOjz+ubjqzNn1u9/EAyzQv7t+ahKDfVLMA9YUV8l3wB1RzmNj+qD8V
dr3lox1ePyBr+mrWbIPf3TlYahbX3PFFiHwAFYqvLkbcswjrU1vSf7LMGBv/CGwjjT/OYvxzakiP
h+qF6t0R3VEeRVK63J8GVE6OVtf9dItDP1vbF7c4FR6ocFDe5PH7sQJtK67BWO7YbAFu/ZPhdwS9
+HB2Z6g19b4/8AEVSyYyGkvo9NYPDL5FM1QGMuPzGJXKq/lRloNmUvhw+6a7GHv5+XGNtZSw/E9E
RbYv4k9OSwRFGRy0VQRt8fcpKDoIstP4x+ZA4lsqtAM8R5nbx5U7BuNDF0lwo9ttxvJ2Ff6Uu2UU
GnyDIZzv3Qz+C5At40p6XV/IdOiCrlhjVWWenvb2eJH0Y2lPQ7JeyqX197VOwn6C4qdbceGjnPRe
5GYbn5Q806zedyDgfFMV91NitfqLFufCGMB86mjXG/m2u9dab5uJpAjN9sq2LgsAjVFT5na14gFP
DxrvTBGQNV0Dg92OULeiTbLR9ZcX0niThS2QfqOSDcRJa7roY8m7DGKTRrGYm2xDdvke0tNJFNTd
qtcAe5WG/prBSct06jU642I58F3aVJwoW+sTiZonl84/nMXkS67SlMhTOvDq1aoeOOFKO7DCSx74
MIN54yXODYMALy2/JAddG/1Jaz+Uw8ntVnwkHYcneCCem2trsYebGjDb+yVqRVgYSDTFdQVzQz69
5zfErXhZ3giNhWp0BY1dOh+aeHeh4FpIFqoVODOHNmKl8l6GWW9Pv2/GU5+YkUXosbw0C/PbkoJT
bc3cXboj87/++9YSrK4bsVwCSmAGcQrPjow0ag6dn8zVf9DoBlZCfsdts5UvgRsXRE0xQj16jeSo
l3WN0M7Tm6F4UBNmZ0c/nKbo19rbkn/5sFcYHiNVU1kXsEBW+qJ2K75L/2d0yl4dpEPv6OMt5fC0
nohxxm5eXCSm6cy5Cl26zgBdmkeWcO6Hb+qpNtWhjjqtJx5HR6LnSiA9W+kORsQV2v/LnutEKJGC
9V80lydFWeTpX2pkmFMA62Xr8gYENdA6s/aRn/7Zf6EUfOUUOWGmdHvmTAL7pfn+Js0d88tjfa0k
rYqJIpsId6+Yqpb8LVFNO9Xy4R1XZjea/+g6vUn3kNq9MaRwG7NrUhG9UBJ5Kx4WYGzm2/jT3h4a
BaAYE03icUgtjLQYDrBZrRFEZFZIosywCWcPb6Y+6qtqb0lxd+u54nFXnBmP4tqsd1oluTBc5/3S
hKKeSXz1qZHayFaBmTBV8h2FFSAtimXgc/mw8Cq06quUKhK6Z4+u6tSs5/b8oFbhh8zx/PY2ODmI
1wjctBM/rZMxtVRtbm4gtuzRnYPW/AI6AOudzGx+FHoexZoGCSTcrzmbqfhuWgbaKxRx0sr8q0NV
fX8YeLvpCHojIz/tmNzHkBunxaFDWYYcmkE9pjM6n7IuqSEDuylM3G3aOVErmabMnt1DqOs9FeWo
HmBuAf+HRduSwaHeL3m+jIZXC58gC+Sm3YruDsz4LxUgfUKJqmWA0Ejac+5mkLQ2PCM3g48DUdLy
VZ7XqhCmhTl8NGeDhFSWejhbKkGyDCWZJHd7kK/AfHNoGO4Ukni/v4s1FuE6BH45AiZ9aWvK40nq
MsJtoKtK7hXtMR5SLPLAxjm7LPThUFalLW7QFeCyt6M0l+2O77Kk7kOBuZ4wlBwEK6EpJaBt8Av9
Qz7SiWt+vAY12wjDlCeqPZalGmuJ40MlR5GEJc13eoAO8Tn5M1usGG+VOgp8882VTw/INcuSnnMu
jwUE7y3eipMP5ZHrjdTHYrrbyQ11QNu/jVfhfpSdL8iLzYyvMo2QVA68Z4XAAOfcntbtCADeYyb6
OkfBhwNeQaxjTha0WKmQ+MDhVLqD6JFU/63O+Q0oyr9KVtowImu4GONi3jlD1bCJeflnBogx2TRI
NmkMgcV4tlWO0tauTSyjHm19btupcsTX4h7Rcez5Z4rw6Wz6KVSbMIsHUSbIfgnAEnCtfZI0bLTZ
wRdl8d1TSoKi01Do5m20J8flF8BnIDnozpKt2fz0ftBSEVw/tbVftJzT6GinOJpoiqg/c6Gzunme
2KB6z8abTnnChaGBYRJs3zEWVr5wOXuAjRaJF84Kivvkot4V9022n5n+ff5iDfupom9MbLFsXVZF
i0zNzZqRGE+IENnWc1IlG0B/FDRJb9YAg+GZ87CZIpS9dgFzZld/rj+ZEKY5q+mLHXeQatgwlWG6
Rx18D6wRIQx2Bf6LS1PxZbiSj7xQP5CXuWrp8G4cSV9FORLmv2TJnFvxkbNZfZ677/0A6LlPEku4
qfvuWOvDjzp9+aZKP384PFUIiqbxKDlQGJIFMW69LzVgm+SDFum9aBdXt2pM2D17hFgvOSdZFOWE
VDyj8gYrgLmn07b/EPAggtSe5yPV3da8oDirStupTRjvO2iz77Ic2S7JYG7dX40oZqY5nLSh9WBa
pMd4w6juhSg2FAL3gqg+OC91syW2RjcPGd2OX9D/xtgTOQTK3qNGdDcE6Ri8F/Kg6C7hsoBVhcao
OmxkFaHRgsxpp3LyaFv+ki6MdQ0/s1TRkynUS51towqCo5G9EF5zZpSi1Gp1FSqM7TtecY09K7sg
h8FI++ddsibwigLmv/4M6hxJwWi65PaA1pA6Vtfc2Q/bNevGMu6vpU4yRz67KMKLPhdRRbcF5i69
dx7CDvoOdxG6U0ehbKyJTvyY9LOdeTLf8QGTLRrBxUC1k4c6p5ZFTwFoal4SWks1ObhffQtF/9mR
N8KQERCliKOgo0yM9tKztp8HyHrAt2teAZoOZzwugr/gMTeK5WCmt6t7WDuqiR1PluUVH3WYQWhq
fgV+NRRdu3bfkSiHSu/WCzsU9yZUUEa2TSIAwm79d6SBbr+E8JmEPZTKksJipkP6pTW6RzpO3Kmt
E+De2PAulFsdB1qb5xg+0P3Yab5jaIMkQhZBJb0BevGLiTAHF1rgZLyd5CMppcXDm296xN/qz4Be
m4alq4nfpn/olnMTBoE+5Cv8zyrAYdn3IXrpAV4CfFYenW5VEOA0198z+sZEc3G+8D0L0ebBVqKX
NdCo/3iSds49t6yTUAsaqp9kpLabsBIW2RsINHZdrouyyjsvVDyvYdh8T+MMurNVnjFvxJtA6c77
TskppVkSGk01/v1sRRmbifGr0qei8qD9uN2MMX+Nwr8zSbIlIN4uQ2xFoUbTBo2VkI/sDBFbCrUi
ZO6lyM99YehNIRO0v+kIunCfHI06p5q1xgRjZQvvPdNjhsik/8sRSNsoCR/sR73TcUh/NX3Yb8Ok
5bxvUIKpgHxwV4Un3PCcx56roexsIlUzpmSyYBDqQyq93y7PEgobDwOEY9GbEA4zRzAQpIhoL1o5
A37eCmABpKVIUGQAoR+DY3h01r/7FvX72NBxjLnVtZZWqOhyuPHCBMkPXR/Q06riqtv1ma8M2cHh
1ktgp5mUSBvlw/k5FDrMLzbw8MUjV0acxO5CoTLJRYNT30jWUBW25kGATROAMwk8gR1rBK/3bMmk
mpMk4mkEKB/uqnY7D+Kr0C4vTkiRvlKarMwiOQekXvOBm3LLjt7qKP+HjzfnbFMId0L69doa2BJC
saBZUD86NkcDt/nNSXMly+LMk6g/OA1iR5/rmSTMn4FiNMNKoaLU1IbFJVWrTDCqMDys1Gc+u7c4
02rg/s49YxZsa2hUpAhbDtFOHG0e/jkMQW7dvjGSF34OLyRAmX0rAePzZaxq/xmcSSQ/Dcp7t99V
0r6tSjsGZIunl9t4MHCAtiU+mc9qI2AhAZq6bcd0tvY46QPH8iOPxxsvoC663DGUkYoHD6IHo7cO
BT8vD7EkSByukoFNPp+T0AgxSv+C8xUh/TnVXNB0Efl5UMqrcz15mCEjc/L9Ufe/kccpTmB5xEnh
q/So0R71Zh7agvQ7G5WMca9mxbwLWuQlMmqiUr/aaOaL5/LWWRYJmsuSYEFs+Ph/KASyAtcCgyqh
/jZLQyFTiyN87QKOpBo29WIn2ZVyWTQJXYBW/1J9RpYW+bhkEt9JJVw9jfn/1Q9bgbPYG26kJUnD
mTw0S80cFbVf7Ye4eK3t37gV30aIuCe532t2SAe+av5gomnrpBQzgUmpNymqvjWKDuqRZRRBRNt0
J1L463G+96Vu8KpHASeZ1RiDp7LJQdTWgp4epjQdshZHV228cneZJFqg7UB1RD4jYRMSDic/K5/H
tPcdBpiUEHavHYmKeGWI21IcPlUdA0E7xwwrD5STO6UNZnmjri88z5M6scUam0YTuUbOG9krHAj0
mIo7tRE7NgdypCer3cLlOGky53ii9ngo4lu/mIJ7xleyRinLKtuNKlYu19miRBnLqC7PAQLu0ulc
goT65jx//xsniN8ldQSTIgpKi8pdA1ljBsuKBsrouFlNOOWFWCI2vGmfTPelmJWRdI1iaQft5IUO
QfUwLQVurnPPL6vpIVugE9KvO9VaZFhQxlZg4Lhc66boZqU0huz+sP1JsrOYfUd+pj0N0XRB1o6Z
vfVJoWgisRrJ48jzOEfxxnIBo94xl9Y1mNqKL6RDg8pnp2unzVpz1yzGurw6RTpQ/SJQxMwQFPv+
pixZvK4n4H/RxB/RRn87MPH1GaK570NR9p9A2cnM58j+2snMB/TZFaqbijIxnuOnKz2SQu12G8l/
QentjxZhdFn4jLx0IRYsh1hEvIapwXowNs0QxcuOI0WkWYo3b3tfy4B5Kysas9WRyLqGZbWbOxaZ
eUNgx7SsMg2CC9oA8JpBgOoHIkJbW7hQ3f1xIc62NYjaaSH1J9duzTw2lcPx2QzBKwK54eEt2wj2
/9zQ1SiIU9AEB/X+0fcW8yg6vYHFiFk+x3Z6UIY9mb8OUZPVE46zwJdLV+1+tKUnT151dcyOcOUY
P6HLdJDMnAvCwjYZ7IskxsPx7htx9ntyHWG+ud6O3O9znacnyH0Q/yHrw2WRBT6ZiMI9R6beo389
mVWNtwjEkx8eaK74227DY/C1HkmqBQWRWpQF4oTFfNd+edQNHhpcdrCPpY5jN3qCpdj8yUWty3JV
iNLoF0prumFtm+jHKyAvhPyenpCriYBYVwR7Ex1y2s9FCOqYwwtTQO65Pd2gGSjXKlhsWA0M9fcB
Oq/ri4VTIF3lVUTyD5N0cU2UzBgE29T2EykKzJaNIX/IOPrFv8m2OsDgj1k//sedsbOYS8KCWq/W
PaeWMZWv491TlHuwlP9F6GEek2PWXMWE6d2JTkpWsFgB4O2rfxpJ5hafdzxiFxQESewfTi/GvGmF
xk4rNUnjP9K9SNc3+R2hO6UjGK9NC+A0JsYKYweWJRboLyAPx3Tv9EvqeqbirdNMqQr8tmvTyid/
5ZgxNwIt2hBTYXgS2EWpyOYWihtn2wDTyho0ovw3QmLyzPaaCEgleW/LxZHqMdBYEZXve/DsGZHe
wXUC5fb5OFZJBl4XkY0ce2wn/rsbra1cBh7fdFvGKLcnxHd1zRhsUfELA3eSpBgpPzrtMB5Iqz91
ym8zEMuksjx++makW3aOQRwIBGN4auzzcXX0lscAknqyPjnCBkD59LbmiyP+3Y419sWgjdcjJl3s
AJtwUfPIOSmjcQsUu+iC0XaZL6VsbqGAsqCd0HeP+ZJooUQMzBstU2oH8rozEqZ+0frjVyiUoBah
Swy54KmwpRy/vGPi54+abkQV/ksm3Aqgym+eipFYOPP+scLaOkKu6e1PJtIY6XTLuN/kZ9AOBwWU
U0aYhGD3JmupfRLGlZJhEETOM/oi9hWTXKkiPTnw3GKe9E/R3NKq34ps/vNSRlFWK5xSh5xjF5NM
gx9oMa2s3Q6DSYqmHw+b+Ut/5O+5FOQvcF1JIMtPlOsqCDrexOFir/vwRCd3yuS0Vaj/JY6CoOOG
S39U88AgsbmXgiPpUZKLD5pGRni8MpZCbC22Yp8da97oyazPAOOeWaCLi/LYR1I/p70DdVkogKxr
oybU5Gdu7C92KiFSupmV4EBFM8tzOa59LLd5lwQfyXWJ7a2snk9lMsLoCr47K+YGw5tRetdTxUfZ
PSH6vCF4YcjQCQ6mbnH9TuUaYTqMWl9YCjNcsoR4Wm/c+xDWhrOFmE+vDYztuObTu9tASZN06CRW
V1+QVbsc6LoBlxeHKtNfnpLvpw9niKxn8y9pmyNBwcMvbW33iGstGAglhQoRuuvdauWDsl1wHwXL
8gmrvV+M9kIhPW8Ycov2Czvi8GshaMQD2fQKr2OLDt2lkmtDtubX9StCLUlzf7c612qaQmeUPVOw
rlNB58lFRjGo/gV7N6eMR3EVOQGp/B7Hmi/BETRbwFKuUvUCgcglPiOESgRh9wKir7Nal7loCLrE
aAtmjuufIF/KbBLnWP8BaQ7LcXfgCkQNWgf4tjmjdZPoeAIaUIGrv1ZLbd9vHlCHLCjTOeG7ZG1h
mkxpDirxaSts3P6mcZN0gnPqcEwxGPCpMEiGUGB32M8V3jz8cW2oTLUOOoG+JuG32alFgqmVdECz
jgxhjb3jbuD04CpivhzMCHVpQc0L1jSrtD89hE943s8HV44P/utHMhF2O9QCZUbBwP1MkUkwdknp
rlsaM4K7am+LLZenYoNEe5LYPT72LqqlGFJ7MJTujYLCkIkJHQ9GVkRoyKhw35KA7RCUdCmNHvHR
IVIe/sewF5BD3tqGEAZnew2MAAJZghivyssuJM9phqvH3eLVvSx44e+fk1LIWkG3kBnhxvJvaWAI
GRZtca3XmdQ/uWHhrUFQmbkAiSjsoPZ5FrUhU8c+RrVRoFiBN0sCyTt2/DLnSkpND0Bj4rpbqZMu
w06YyIrnvSKG23eX/HVmJHst7CVfelOdlLRZS2d5sCNSEd16AQKZtcYDsvrSY/rNmTNIwTuYydQi
3dc6Yl7BbBKcm1qDzGS3qIP5JOd0zYx24FPHIan7rq07g7NLnC0Dp1jBpfEomt0m4o5jHeQ+9CRM
xN/MEfWHgOEk5t6vetkOIpiBtRm3B4lwzr2J/wS0QlvwOgX72BzCWq/uUGd/hzPEoSlNNoRqT1MG
4GMl8pmtICljOF9arfWI1GKu0RURBwfgzJe4uzsmALRwkmCKTCwT+hjWNtFeauTsD7YcnPVmR5Ux
bdX0Iw0wNMgo3TqQ5tcAMpjj4N5W2ub3/78Had7RmWxXdyymyVFI6S1/apIX67VA1yNsGgRBuXzX
RetcqaTNk2Vl58f1u5MxoDzmzl6/NWyMxqsArpZFkh/uPzusMw6YUv++HD9wB39rvYnZxWpT9DYG
CfUsUM057XTnzC9kw+/7ND1eORZyEVbds3oV4OGaO8X+S3w7mpgSIrwOB13mckkOd3rQvX7R/1sc
ky9Y/2UIRm4LccqF45tVozLz3+iFGy4TmE6pZRwQGx3LIK2nMNLUzNDoIQ8+yzFaVQaZQ3nHcUpq
AgbjVHaCvnOL4KIiY9224sOQXSWAaLb96dihXbT/AQmVfYAkClgylo9OlJCXbY0YpRK1KqizVRAa
Dnrh6Ys3gCgzesYze8MCBQvTMNOP8R2f9Uuyn6/CoX2IeMw7hYECgl15HswF6Jwu5/7ZlqzBG7bf
u0U9PJfJUC/S1RuMlLo4HcTfPxUF3OKpHelpagj7MbjOKRvoCKE7K3F23IKiOc3h7nLAwbATiB0V
pQb9k/gfcJp7iY2dFFJx/Ohacyqx7tdYh6FYaQzYqfDXp/QP/G69/SS1AFm5Ay2mydkcIdpNWG6t
u2/pXmbIJ841WLCJ9wvrNa6WgAHfaQv8LfFgA3o+dzXzzVV1RbpeiRbxdAsxRRqc4DSK2Saw70eo
5a+IXyiuwKTeYrZV7mkp5q+zyyQgxc48foGHGJYFj5q008O1rNtPnpxcabDEpR26a/nL1pviMYQl
b4ytSmWa2DVMfE6X8xfp/3Mkiw5vZmKf1ntWox5gt5YThmD0BK6xuNyVYLvdbNFGJ5/FiehwV5bH
LycW+SFAJdm64M5GfQ172Y8WsmluP6MSp48n1BZ9F7Oi0eZNVD/zULcvr/vzPR0qiGmp4GhH+UW0
EYT25t47yrNMXVbadiwYstpRKu3XdeoUeqeeuIagUQPv4D1+bPtzI4k8DgZbP3pQcasm/DUDiy0M
ZzLRS0Jq7iOuwhMtvcZoZagOrXg/wKjgFSDM+SyNzNpdQY3HF6JJ/mdjA5O0/FAYbX2//SRcZv+q
ss3Kd/FmLggchmc7zPOvAHO8mbr+QdeOKtS/vyeUG7UCoCiJbDZz8WpNdPmQmETBnjpIqLsF7QhU
PpVYZHOiTqIhOdG3uzg5jsSxyZc1ZQ48n/L0amHnQyGsAxBQNqQXZ7qB0HVLkEkO/p9K7qvzswLe
jWsmuAyg28xqGoAUxPuGXn2VGmAH91M56Ra+BCSU9xg2vPKkqwfMvUtk45687qPJF1N9dV8VH7s+
RuQrL1FdK6p62CzJ3vMLlTbykPmtbj0OTnYJ50JP+Ye+Dv3F97MGIi1vExsi2/cO86UTi/GCcuIp
sX2PrJFpAJoZQS2z2GQmVoUJy/qIpa6sh83hIJd5zAGrWYHS/1VF/5LwabZfYIF35h+XX+cpe9mh
Hs76OWJIV6AS9d84YAEHNlYA4cZuCBtcnBGZyGZUtGcJm+TynZw7CfEc3E1eSdnhujrCIHUyV+td
7BaWVFZ96We2KVQEDzvfOoMdLu6taS4Blso93CwkoAEQx9RBcUeQSyMM+ss2bLcna4b4PExgSMTL
V1gk9OWtvWNp6hdqJEU4882TF4FKt1ul7fZPvWztqJHa1u4pzZ1GHX5QRyFOH3D3eRXSBzap/QjA
VB6E2jZnwIjf76RwJf/sDvwGRDA+i4DPdm+9WGaTUFat9L4msNFmbK4pzxXIUXcd7dSawJG0TclG
lXWcGJNGdeuYSItaTsUtmhmHl6PzZRJKNW/o8Jn34DlwIS57hnZmyxJlVR9ghSAb9JzB0wEpIT/c
yVQ2++V6tpwRoTa0GxqDuNkgiO4u5NFC2RPbIyKZPM/1VwRGYYGXmDCS9Q+QYB3KVJq/ayy/Y05b
KZtk/T1jzufNpmMuiCpzHdPXu2XOaJ4hjYVRkjP82nPPQ0YU4/sBXqJ6L7ufnTOA/dKHEGOUihFv
801HmE8t46D3jV/ZGwE9dso1p33XwIuGsx54WM/oiElYCkDdoJo1rCOXwR41082kRhwPuQcT/0kY
kyOmy7gn/CC9VHxHKB66Ay+3WHwHInmbiK/LQhcuz4hrsN+XqcObF8RQnHvW35n5hZ1/Y9GFUvi5
G0rIZ6uuzSBRntr4CI3zY9kpXuqQ3iQRaKXRCgajZ0pS8Ojrkrv99AMi1zL8BWAsL5QT8iqdbTCm
RJlcQuUbQ/Xmpl+QlDRWjHQSgc254TZy8NBLkv/k4gj3Z4IGa8V8OLH3dU+gfzDDs3REudWJFx1d
quUe8ZKUWC+jsNgaBaJkdGJamq/Zp/G9Ts+nHHWAgLPINin/7WUfmvDvguxgrlvs8+nNmt1PEgk2
+nS5hmGk4t/xMBGpLN6gykXUr8dONdvAsb8MY9WLfnLd/V18D3y3DT4btPa/taZA2WDLlGk0TPm/
zm318zmWhSA3INi/2qMlEz6snIFc3dxvjQtZxBiRafuz6tsTBxsBRkV0gbBZhLBIPpnVS1YAbTKH
Suf8jc2/DmM73nD/z2OMmfA9Y3vTnnPY2QvukgKEHYw/3UHB43wgTgL3yGZvtbUNwo0x4qTdXTmz
3vwV3fOTF/2aLFqM3E3FaE51NU5mWFQxym7P/rioslXdeR9+FRLDomytDPnaNrY/HuqMiI9JqiZ9
EeWcT4E9vNv5+MYDj/2AAzwtQIDFPmqro7P07C903O0uO+XnLIhOl4xi1Z6hmZ4LTB4kCCu/GF9e
2+5MVwFYL3xa/lqsPJB4cr5jfiVMeLREZgZykVEJaJAUkiDrhrhclX7LYWEq+uJ8WlOnictqrPhi
bmcPgbEmHW9Yg/1ezpzhdHwEOYP/zyXZiK3jSttCAL1wn7ADflbsRpEzQMqdtFnMNiGP8IzhCbCS
BF/J6e2IgE7NFnjxkbLbQ6bfRrOfHn1aUWm+UqZpfv6am3W3yr4GIQNc4HAq0PZBUt5aif1RzhgM
mSABIVcqITofZ3uK2s6I0cLueLsZoP/laGZCiE1GOJuCQ4um/AysYW0MUtOhzb0P/xT0gVEN21w+
67dUirgOvFZg7UsUBrQCR2GqZKhZ0yaCJkzAMjPQbtllT2kdxp1AlJBuq0lgfUEJE0UNy3Ihl59v
NRtmWHllqRDdl76yGp0QKxd1FxKU6eoNGaijn6XCUTsKgB/CUmozUg8kbd27ZP1uvBeiUDSqjb2I
dJwlOIs6t/pZVKlMObJ3mDzfSBX6wOFLzooQ4hW+qDAMu5PKfmLcGOlpzDkKzLQH0N/Ul838J8RW
fclKvW5YYSyOOU3G8CzxTaNkj0F1JoC6SUFyZfC8Xqu/hrX9mu3J4z4+K5uAazTaeNnfe3kteNne
aXucg9w6cYYevVFvOQ9TKkbpehKaRIyHfcWKJ87UwKdci1ZFnV+tX8LNjgKG3BjpuW8QvzjROPu+
8kkoTjxz3pqY910YumlyPZGHC0iPh+H2nCin6/+F0vrganOOaKBSondGDWlad98QwiPBfHfAY18T
bx7rZKBzltr9dFOBrsvMpx5quwcv5D6NWr+Au1IKt6X+VNgrDWqf/0wItjDxvyOzvMqEmzTGpT/L
O9VqZzbn9huOf8/Winuvt2oBf14tNZLW0YYU/ugeUqBakYgehvYiky3bLKUfEYx3/9n1Pf7y678I
7v8U74l7mMFz7LINUD0I8PC55MgCZKvZfJ25thN9/VxMii8jGTZ7vuJqgmVLuTswyu5PbR0CwV0Y
ME3K2wAjffWTqXLlvt8d1VgANQsAyxH2krJYDglSD3P+heYW+rExpA3JGVfyTOIckjuXdGm19xVQ
hJIAWyMEn+JOm9VEjXAq01qXDddm8cCTPC0eKMN1Zv7zShQpVvmc7lZbcpz4aQJCuF+G144J/saj
Mr+DwssZ6kWEYqHeFp6KXpTXIqTZP1PW0mr/49J+gQk4Jph72u6E3lPyOxAO+5r1Umde8eCCk0YU
Yd67YeIhX74ngIyzNAD3Q2q6Ar42soEXEORJlyscJcuVRnJ8M9solJWcgWNRq60tHTDqpDhPHx0o
6dmBWAS9Mo+wW9VD+mXWuFiiijRJam+UMT5XItjf+IKIQKIfMLW4KZmxPrUNP1BbMMvHm9GgMJ46
qgiqbXlvxadgqt0TEuRtVYUsxE9wYQIRILJUu3WBNlsiUU3GV0bOZ/JsVWzccK43/G9yuRNf/xXG
ePOzkPMr/3T3NGUv/JZfRr8f1hPs5SGjNXwGqt+v3Ik6k3jdJEBccoyAm0kaVVE3/CD5ibUpFRI6
AYK2bg3NMuDa6E2raT7OjYSLaONaoG6aNlET0G4psyeumIb2wVl6k3f3yzpGB5DL9mhtjwCLPGJ5
/quCtQ8OhwqZ4iLfkK7V5A8XG+tkFJXjnzrv3w0937X+mlaJWkxtTXxeNrL+gDXwfYQdSqJrjZHc
cnLzdy/wmQDEW858PNm+B2YoDIGcbCglu0DKWU+lN3oGMuGSPcTb1ip+wt878sLZGwDWHkaw/SKk
sE3M+QmD3bKe57/217/i0tE8ZJdCuMmhCg4YGTGp+GcZtEyBHFA+cE5TvcaZCfVvqAD4NhkXOy4Y
qy7X9PPdb/e2H+LsXDxa7QXPjttsb5AtZxzYmuMt93loiSiGQkoR7KEIKOt0N84wOJ1VjT3Wl4K6
MzuUG/bdfH+KqiHPoBjTv6TMXKj4LWB1I61XzaOFctH7bmzHWvqoBaNNJdScga6KdpclKDZddXTG
OuotvAfsFE6f7L+O7qqpWdsesAfBfCQAmkwCdeNyyImfhygwKALY+sz8DFw3P+7fIlbccuupiTAC
CXQ9DWrTJzw9G7RK1VVlmKsknvLx9EsFaWS5cTWeDaCdEijhFgv2jQywbdvNWVgjgfQ9tQXE0rQ4
psx/u8M5qRgcrPvhmZaPl8lkVR4Y2Qb0HXnAU7WO+aQGSGBUz49Zk2HCVuS6pMGgj99XdgQ4BnNf
D/VuRv1ypdBk2VGZSmUXdSMMlB7HhfLqHd5k6jk+EoK5vsu4qS7sg69ATdCeKxpgDx1AFHgSOLk5
1UaPml5Cm7Z94h2/ujF2LpOL/OtakKmrwj4dKB8HXtsx9OtWgAgeMly2s8pk4I2cztuzNB9j+TK/
FH/YqQBlV4PL/FQuy5xbUGHtF94GfP4EwpI45JnELepfTTzhTFbIq39dS3eAIZVuLz+9CFiqJJN5
bJNtV/gcvQfSSHg3inEjMz+mY8NNmoX11T8e532rzwNT/5U/vMKlny314Q69JdQfjPawLhoWd8Sq
JD+Y2yV1uN+6OAvTsi5nu9afioIRnjGKxbSdeCUReEj92kAs2ubL5Ftfz2oc0wkw+YJRUhGdn+z+
E+vWiBMmsLRB8QNye5QMIjQlh8emZfLsEFtKn3IBSoU3uvTSdvxQrZfLG0lZBaFxidsfo28Boykk
CfKuxphkAgZwCN8A31DoGcRRCQ2c3xWXg3owNpkyQ7yyoFLPvKAbHK3CwwKnQTVk9NpZsqq/mcBT
SC3+0nMXRCE0+ReC4vwXDlg/lZ/vfNdOmbrfxtKU0IofoWj080CzP8MM8CfiadTQfIwLBqi7sMR1
hFgdjkl463kooYWKgPmFxLVHB2CltvOHQ0Ei9NrMTb9BPiIkyWqtQgaKswja/VHbjG3wf9AC+boB
YM6f/g9IManTHQRlU7N7Rlbl24QcOC3Gpv0YnenDKv5N4mjaQ6SnI8LqcZUkOB8eCaeAIRbeWinc
zGGV2fCUGkcr3yTY8s93LZoZUfNQIwuBIdUmfZoD2jzSCEOaVtebPuLMz+TOErqgScHCVWymb1I/
7USil9iD/+yyGqw53V7BdS3JR3dZ9MDE58qZYQ3UjkQE4BuCjx8HkG4QCiEOkGpCD7/rLQAoH7EN
vBZIQolYUzlYB1TLnULUKDk+ybY1ItWknDnNONDUcEtdkXPorCUsWHhKnqzcx0EPLR3h7fjR5Y6a
N99/6dscUx5LgNfxmDnxf0cHVRq3NezQjKB3g0BrXj+QZaELrKtm5w1sB7cTZNRNqOEo+zC/byBC
88IaHOVjDvflFPVAj9xsCowV9sc/RlK5pUcy0BYaVH6QGPfuLoqo9Tumv5JuzD1TzxpIlhWZ7r2m
xwEHFAqenNdgZxik9Xma8s+d+QotprsbH3ay2ypxVVqkZ1ZabAYo5zZmC/sYnTPPocXaWmzsmLui
UMY9ek8kqbEf1lwCrcUmF65k9S5gRY21w0UBQJKY4EWs+UEdfUk2mwcmy0UQ3Ecw7n5IFyecEtXf
/vVUBLZ6ydSoS0UoyB9gC1PJfgh02cnbkLiuQK5l08TEKOBMib9vd5bJCIGtKLWJtWGY7F7wnxjN
H0feCUGsi/bipaBsWBgiJX69oJtfuWlKfosTwh9BuPXsm5ZjpnxnWZJqQgIzfpmOxEztn9IvoX5G
23MFnQadfYS+Si/V/aNHNno9BrITbdpq+4HWnB7+E9M2GBSDDMi6vnn0VwqpzeXUIfR/oYHFr9iQ
qXGoi6TGnb9oVTKlWquxyB7kB02V/Cyc7v7SDSIx2sa2MssKh1z3gJeCouz5UC8VX5jZ4PgLUkCG
mI216NMD2vOWZGbpHPYPUR0XfAgG8P7tKch1us1EItVdrdpxNLMQ2D4kJgeX9D9gTq2BPJpX3d2D
S39ziJxGZhcXrUED2NfP19o5BJfzf2IkFmEA9uqJfALB5caN0o1pFJ2MnXEVkVIkoSEi6avnsYbG
ndFsqVeIrZjuTVsJuMKrdmzmBhi7RWNoc6xMGoncvijmeaERyMUbLJbeJ7gS5mpwEx4Pg1Y8LLtf
bp9+DOweFAMmNOfF/C+OOW28Hl8ugLnOty2MVkyrwKk/EdWPPjYGbaGr42U6MWVtW4Ad3/Fq49+f
RxJiy9tnMUNvmc7utKwK/SL7hLT3k0R80VjWZ6nXsviEjYCetFgVfkSNtO/wDO8q4kF1WsD31Pcg
yAzGUNzw6wLmS/6hJzmnWdwOiooY6Y0B8CPGJCLZ9W55eOlekwqN1c/+hSUqgNVk2dAkEA7UeG8U
NqkUiPumzB4Jh9klLvwAloXl6nQsdL7a5y2cIaDk0BvYUUqEpET0Yo8SxrjkoRy11SpDugojHnWV
XF25NysZgune6Gkgg6yEJvLVYbt1+8YmUGmMpAdGcZV7xqJknQJ7jISY9jiwLeYNMHN+9kvMXk7M
HC1hhquY8tKfbo6+WTcqvvuJgkdsug41LbqOlc0ZFvkV+coh2q2pruWCy61vY2n9Uy3A7avC3Po2
g46z3e9/YWwfsArKJqhTQp1I3nehxpnfKIvldeD6H8rkmPNfUjd/prjoXqjDckFv7wari5OJccy7
9clqUz2ZSYeuMDYMNqya2BTjqVxU2QxOVvRi/tiHjNl6PpD6v7PByNYK7JXJHyLRoHowWPmHy/gL
hqgkJRQZA9/bZCUuFfpcAFkp/tmO2sLBKc9LrC2DankC2HSUkuA1cFa5w3Kbqsj5FAO8a/FYUICv
C8gDrH99HJTFP4cVN9AdkTVRD8bwOzmc1+qNLlfygpUOiLEHyUeb2LxAQBhxeJemECgxsGC3obvQ
p7e9XSdnoEi2OyeMQYQ4KfFPOfc1wPXwZxw9Nv2wBbLlqYN4qjPTUS/Qx4FtmOyI8pqNF2QL5x55
5dDcn1HBbavRX43PaUCVelclcTguepEfWYb101LhnXoRhZcgZ9l2IwhNxnaBl+lJOQi+mPmuvzPE
DaVrIordS/Gu/URPuXbnOQfTVC/sVU/X9KTzSc8/I0qxgLjHsbC+gvAlTOZOF88q0fkhpgELEljz
jTlYRnlWpsG5r5u02dEWbRFx0J/NGX2ubuykECHVRk2PdTVVKJ81B04LTAiv7795JFMi/ZoNUxmv
BA6K6idTqOis7riMDvA55aCJZEigFhr7EzG40DvNv89j9u2YHYQFz297MNrAHxVniyL+QFNEhVVs
4WX4DXtQZAO7q1+VBn5kkDHJxonDIR2zDAV8QoYkUizpHilgE0AtSyzjiZjNmwVoqA+WII/YkJUT
OP2sbpui0eDtIxjqIhQ9dt0BIe/TDUbDuVFCiuy3d82Im44X34pd5iIqbrNlqKIgl8UOi7TYnQNT
OJlaAZCBLTk+B/zYQfvnkNSrazQBrZJFbTiyedFhZMMANcFNeomh2k78RSleoEBi7A0SWYcC4ru4
d5N+XPKcvwi6NZBy3fH1KXnuxxmYmxzR8UqIJ/+7NLLCEzBTQYQmUUiXT/IXUk/d/+Pe2IOi+uXv
AfaLxyJx35Vi7IC3qxkKbwdWsciEZCq5zyKIxL6CtKSNhlSskXA6N7CeCxkrewcouU05KiLOpk+b
giwwMpp99NFD4UIbL/uaQyNH9OYZYAuu8tTwunPRFzNCxi71N7RtnEqtcxb3RdnlRi0nj2c0UDz/
hiW5gYI/Di+7xZAcUl/Kq5ul6DRHsGOVmSGQ1Cj/yCz0MIo4eTRActpLZvIROUpEOpBTGnB2oVS3
gmf0v8AL+quXOnRpxM9DkWh4qKeaNZgc94NpUBKCPORpW/OhAcIJzCmUTCTAh3AETXm+wNCbyClA
B05ZmxNZ1i/KRhkFhrkqMyTU5hAXXXSxyYWydb7rKu9KjT8NUPes6ursl7MRMrXyaXxm2pWgds4t
YGTY+9X1qX6AZ6T+c5JQspGIHeAbJRfR5u0XQxOubXHRd15QY5dgDV66KfqkzplKx0VTiR4yVMhx
J0CPgG611kJbKg7N3+f9DRqWhfrqkSSjWlv0DXJwMclbW2CCGVwe97ERe/twb/WhjVAJrDI7+XXX
exqSjmDXH0wHLlwMGlmYJgWIS8s/F9whdd0qn1Bxw92eAmGJY+1QnRs1BL9mSr8n2VGELAFsw3XV
iKxI5P1CisBJpfN51efFaabEQpzgNGVjVmSe2EWTvDFqB3awCipHK+bYFVqWKLSyX+cgel0qIY2j
YReA09vjnOFyQHtALxcmQReW5ulZXBOFkQrbSQ8XPnM5je/amuYoLyboeQ/pgdEJPJrRLCrnMaJH
5s5UL8war+uJTG7QN0+0P5wx3lDSU6ueLkKoyNIgxQ3sj5iu2cL2WF3bMj7vqnmteDGnQIa0PvYh
OIG+dFy8X4IIDnt0TFULzhfpnGz1ztjUMo/9uS4t4P2bMqfnMpZctRCutuOm7Sm2Glb864bIOfar
Q2HM5opvlQ/cqVZOt6CrvXtakuDUxja9NSQcXD6yeE3lLz3yxjEtXKzGtVZwO5tvffw4brKDt7It
GqM5t7jzRp4pUd/X3FkOTXs6ZpTBnA4BtdcREHFtiRMlT3W8gTWe/H9rnbWRXw8u9ELVCNcg5Sfp
SWrUO7MOgdY3Y+RbqIffM/PZEgln8OovXq8rsw11N4NXJddRD2ZEZKlkGmp2iQWKZx4+oAYUYPt3
SEH0LuDwCHbQ325pilCHpYIdeicmUdCMc4He4xUuavE8VRLTO/XT+PbE2MNRK/00hmqHiDoRBrPv
C2sK4KhSnZQeoW2SQzIQ/p+jOL4vV+xa1LwRfh3y3I8iR6p64oeoiRn3cMB3PaAShdM1ANFJgbzm
0FqvWb+Q4waR2L3K6k6H7hOKq74qq2DHJUeGIgRs7W1HqSkXDqULi+InTku3VTys/RrWEAdPI6O2
fDg/ivF//VypQ8gk6+n6jULfzY5tJjn3RXvCzqyVwrO+KZIHPK5fhDlSXL/8hevVt5HgoQCsP6bR
1//cLTMzTBPLP+nGjgMCo3OEn/x+5NCcASOpqot/5eyxzcwxyarB76wUY9/sPIQIidd8zEWFcsQ2
LWYDOkH98oq+fXGbZ9YlbQMN0n1A5tkeT0nkrjeIzw8x6zhpfst5R/BDN1RyNglVzAnxP4gL1L/l
li8TqnWQmGOJu5w28T67YgyJe8dnxixyY4VMyDFhZdPFOlkOdOAm1UlSuOsHZLI7BO6G8hMKBW6M
TvlskbCByi990XpsX3nqKc+iYL3c3Ngq+vBoMpNCHNp9x6BJl+dReSXbwJeuOeFFUnV4WNQ7qi4S
Vc1DkVJ8y39QCiG8WdO0RsX/c2ERCsih56pXH6Sb8XEyl4VWAMKzwBJgkiGo8S1mUOh8CAGTk2mp
mshzTBlEIQJKz7eZwBfsFM+T0yWgChUzPF4DIWamCPeNsH+7vA8IFwjYJbuScqGr6aLoX0aDf7VU
swwqDnQ1m5v4FHRiAZsECEvGDowaCZ1LQAVmHS9e13WTEAE2WYE2hou3VKb1N9vLMg4aoHtIS9ha
L0ciPi3hImuJEmXijgaV7X09i0eODu/d1VJMrCHmqAWhQZ5PqqOZGACbzfvWHJWOd7nKy83pBts4
49ai2b3diRgn/gPYJD51J9plECyfHWxfWlxkdu1g2sdtsatJEtVC0w9UIE6jQ+8c+j3QdrpTK5lt
+sB1hxACcEyg3s8pnwxLo87qNCUMyMp5tGshbD5ouwsC9kj3/ysdXUZ/OdXJByqANqGVHasVupEt
pn07vPuGRBznAPvJxKJHrP6pxpo0hVWMVdDLt/DQP8BLZEFSg1jaac7ARIJH82zZk5awTFYp81WH
SKEp/1+JYUcJZsJfzSAYv1iLGPN/xdBwcqIJk+e1EqCOCmyM/I25Q8KzjFzXzlJeXEL9uaIPc13K
SQHTkl/LnfsgfPJSwR6gRuw0+qXiXoA0MVqByX65g9Ix9THq7xlAsYh2qhRhcIb5orWtFo7Vf32Q
8AW3sl6ilmJU16KTXcv0UFRBvKXUfnQokI9sPn+geLjHEPIiuwpVJCFhUn7AaD8KnOWA2ki+hLPd
ZvfvSPiOdU6F5Xm1afmQLE2jzxK7GhxnPBodkbCf1J5xYb+oleW+JhB7skkNPKhzdFUNOKGoiRoG
O9sd5/xKN3Rpq9BjFb2aNrHYcwMtetBs4epy3qagD4ea8Jw86VL+mPv0HHvif6QOzkdYagH1EqFC
4bx0gztthATJgtY1iSdZDWtvnseyDP0SFntPcRWa1RjbFIyuBpIPJ27JagSRq42njPqaiBV7sVFR
oiqr0UudX1f3FAvofAMcGYGnAlgpVT8beWoV9l4JkYGm7y+bcLUnKi0XBLxw+xqaZ9zJK5hDtbj8
iJQfbkxFrsnwpkxrbUL78iZqfYRxu+myf2CkoythsKNil8g3Sg+46i57I2ZDGmwx8BJW67iIvgxF
qA9+njx5EYp3/BqbprUxSl/0CUv9Xzx6HEwDkFrxTp3w0H5kfTQVGxEgbhasbzIZJzpcOhRRn6H4
dwVvxra+V+bfBhZGra1zCDtWB/ylQaJTR3STceseu14BJRxhpVPccnOQ9v9pnwepgve9JsGtmmDD
Aij+0/1k8DHuztX2F7KSlW4dlL5g4c2Jn5ggo/Fzes7YX4ZHVKFmkv4K8IS3gzr7Eky1Zdyghob2
GPm9jH+SEnPZZkvRGi9OOeSyfrEwXVvXHN4z0z6e46jvl4FoKktDsgQ80aj6ZWANlS1BgK8+0yRb
hRB7lwRFDuf/sPtvZtlUVI2hd2SzbJi9yE3+BoVeU4VVY+ZLzB3akeAnl94Y9UtOkcGqxLE/fI7N
aHKORG4QLVuO6ZrtBHmEahVdzcCFHNyGeMfddEikzW+EYs1V3eN2LBWwQK8KlkGbgs+pvLt2jCof
6s5KFv3PfYvaizOwqqJTiG1X/jnt2t4jdVGCeMer/JPXgRXXvO7iLDqQlI5xLUGafQ0IlUFd3w0H
xEEAvk7OoFEioyC3qnT2z/kgtH/CrInPgZgjn/hneJn3Kguva3jT0Nhq3wquAKYX4MQAMqOmi7va
esLvOEh/luj6DhEx/r+m7rkZcn/nJGbI7RqueZo2lQRfttx198hOxZmhG1gJlFmQqH2kyYvZzDHW
xRkQoqXckPVqGwRGEZi/VWuVGW6rJhi62tazL8+uKdHTqGyqbwZkuTbduJ2kwVc2M3qcAKMaAFUA
MZntm8sKcmhDr5JZl2bi2tkViXn7MFkljtWzLa5dXgSQm5Z3xewiUEoTsEUS0g0yf0rrS+w/BOay
g4ItZUV9hoKqOi/yV9UcHyOaNfkEUBn0QYtQJsrxtTEQmgs53OtPdPkFfIM0x8QHhwtz8HzXxh1A
sgX2yKUJcElq+mVb9TRr+53sR3ctILkmCLyXtGWYBioYLU+aKLXN5OcLTPaLAbZXrqpcMI6mmCeT
Ory7uRxvgFpZXcZ52F/gTML/x+Jd1WwhuHydg+5mwDUUJp7ZxiUbMvbVGj4Ir0cXjnAJL2cBdo6u
A4Pj717WVkWioU2aOQ4ncPdrpavoBGAOzxxCarOnZLCFODMO4O0QSyDntQu2+3XH9Si7DxVFQkHj
nWwcCEt39Nb6UDxH0Qn4Ci4oHoaLHf7JOmgfadCHC25m2Lj8ce3mhWGBIMAEONZfAk/m392qE6SM
kx3uEmu2RdfOjuuYNm0Gaayzvy8gYiLygo+atVgY2LnZKPhd+a3kRrsOly//ZqSqxeB+CqHyD9gf
wPoh17N3yQtjFGm8Zrw5cGCa7seqzCu9yrup73Pf0/8AuHofhqfZSib+pLloUnlbs8lGAoq2isyN
pO+k81Kcm8I1F93Ak0hkU9QS0N4VFwZBDHZivzwNSS+z4ap/ApfV7jTL95r/uQiTaL+zMvjwRnml
9X43S4Wc1YIVnYfzMzzKfUgeu8owdT9MT/BmPE86VRfZNw+VhQ+JxhB82CUE14yAL9J4mriRNN6s
smrMTdwWnEvvbqKrWz41YgVvogP1h8sWtbA/IcKGCu8FpUZVYjdfM+bSIHCmVc6Z96t6lwkbmiJU
Toq+uioF9nWxsKaShzpmuc5gibbqQO1xEhmdN9QfGEmqEOOtUxa7jJJiRGJvi0XjaMp+uL4laZWK
W0YSg2OBN/5HlVITkdfAmmZV+dF+jB3tm2QQnvKx7m56RX01lfYMytNO/X/hzQ6vVLGhFrVrhMWY
HlwakM5T0nECgMlCY3gefHsDDFDSpKcXq64k98YtQJdhqrjpO/1FW1xN1SHPrChrE2RSdjC87IhN
20hcqj28YkdUv0GTVrn+s+6wCJYxnqANTOd5b2wIl4+F70ycyH7ETRBt1tWcmN6rNsrZeRpKrCgC
Q8lmT7whG8a6W2l0VHyCi9BT8hd7nxma52Uxj2dnL+niShWJ8vU5VlmFOgbhfBdAxvtH/2nl9j4x
2AcFRkSWmuQyrgkiJ9NsBPwB2ArCG5f+2MknWH1emNdcKjmp6U5huf+7qcBZP3purzOhydjQAgq+
tSFrnmltuR+IQDkjjDYn5e83fQOThT+PP+Neuk9bRSRKQMuJwtL55IrUw1b6wwTKyS8n0NOmm67q
4jaRuuYhNVp0fkpeCaXkUP6qEijggpRPE0XshYDeaItYzL588gE9OUN78UtKhOxXrqAADbCSHINA
VpOqNG2abKu97RWc6oVAL9+nVnP05D0kHDT1ntfqaSLGgBmFBX3j/PkNy5kV8RTuyLY2gXQC1uoD
DSklmDvdQhBVD/kiUaxHJBEP1/KW8MfpZgk+MSoO6Ko6WM0/2IeEXU2cXLjui9FqoKFc5dYAQWRy
3mBpsB/FP9Wlh26twZUsLgYUuxA5LJ61hxxmhFoMswVpbFHxtsmfdoyrjo/zeArxCILIKyfeDMys
UgKmXVXH0OX3TBTcJYu1wgHUgeNasjX2B0fS4u+lc2qJGtTXJYiDPNwUrLthSuTe59qlEGJMqJw4
U5KGzaquOVAjNXJM/GY7fiMJh4hS9vEdG5R2p4wX/AZICSOnwpjPboGl4w37iEq1vZr0CT9p0Qf3
Uu8OzpELZPCFkjy/fwTHNILTIa4jv3nDQx2iGxPEzJFNsdX/SuIDMEOk0mw4iYKhmpJT6bMN+F6I
0hIxXfq3t4/6e78XpzpIVOZYWFITclJ9A3BJRH5ToBsEC/mMy4Lruld2yIYhAwO717xi9t2CBn6p
Yq6bMVPj5jKyDfeaRuSCt4TGQjZ5O2bfN4rrbNmrWOz3YFJSq54CpyUV3FlvtJvvhq+E0zqLF3WS
LmQpuUVUkPd0iPTX/haTb5hHFtYtZztoyXAbcACkfitH2UkUlhHaL2bXw8/pRwDBz0+hYzr5PuIc
MjuidRJtb732zrxq0hv0iGSoVWC03P+A9Im+nD9SjyMgErBi1kHoeJ04XgPUDLEkSy+9oVhAAySe
CNTZMCQ1o3Yus4YA6059R/RfQQRWLEKmmaRtlCAX+OXHNhDsjXPv5ZvGysD6PwC0cUt1ycAQ7OpE
9flj+U+FByiG7bRxg+sfY7yUILlxYPC8kEQ5JKgWwuHWUBN91bi9mlz8KU2NKmkDDlkdne4DYjPZ
oUU5ElVSsjWukXwtiMQpTUNphKl0I/aUl/nTc8y+tG5HHGN8UUYKI0Ntp8RCzz2ErCnh35nqxO6a
55FD1nMXW37BS1J9GDkz1zrPJXAK9hwQRHUONoKqY5cDchEi+yuieboPKePqDroqV+IUpaLIZk64
wslrQ4+9kiM2hpe91orNcoCvrY20yJt/kntQ9qMtjvOltGjpFNCDk/60BvrI98FYGwmNFITkgYuh
lhlN0VZFlPyrLilnHDhzcEs3ugnYuTw3yfb6e7EK/PI7/N6S2GQhi/YRN43RDtoe/EmK8bcymn7S
l4y5j/yT4+Rj4qC8l9diXdb8bwKKxwhszf1p7NK+bQFkujgF8TwjJX1dU02Yj8ymQ3GJpnGSTbBp
E7KOICpHFLl51gA/M7e1QyfR61EiSzO1aZHJVtAJPq/MlKbhotoWy2XC49c7D8ktp3/mWKc0gO2y
xyAZpPLyVYGxSa1csyoPocMdpV7Do+mQXyCz60rVvK8oetPsxE+H+eGymm47aN48ZtEC0rK/o+Ox
GHpIFcTzvMj6WXJBaD4bAN5ssd2w0G/eVZIDdlxWlog9tXdFDRpFwQlDzXSG4FYflq0JH0XnXrZk
YDrw4KI+x81v1FeVOoKUpfEq+q/rEjst4Zer5b8siXi4K+gi2Fu80v/nHR2EEcxsNEE+buyOp4CI
AQTvXBWM1CkBXbSwVQFSWBxd19SmZEyEhqhNHPc/BxiUN8BDVn2/iajiVXZWlnXcisNd54G1w2id
rJeXOPenscuBQQ5MnWKJWVB6i9NbMav/KD1OSUDYoE5BTD7CghcIE7eU373X5vKUdiP+I8x+iKTc
RQ/j3T6jInv2yPdNXE9DOU/b+zDdv8EHq5Az2xk7mZYqNbibyktlTeQt7mQ4oOqy9iAap06WJ7sl
wl34y+aAP6ueXmL3kdTnGftyP+hJlik1jUMoqh1QnEsRSUukk+aez3pXwV/Xb3c8LufqxljGGFSB
nSpF8ho4f+UdPcyQdQrS80vftvJj6HkNFeH2yJ+NiFKsaBqdarDXb+1dQLE2HOIym9imo31nbVjE
fHN4/VDDePrT8guC0PPZ/5e1b4USTu69nyB0nMJFVubXmu6erFAW2ptDpu3BQLOHEtMKRDBrcZr3
zZDHXx3r+UVXoF/9Hcfyeo7tosI/PYK5tJh72XPDualRN8yN7q+r3FOPPOWWg+x2GWITVQPaaTDK
7C3JqL1g48gmsuxF8+Er6jKkU4ZNYbQHiQzXBc34pknsyB1S/ZcuYeO74aG38PmCpvrl/CXm1k0C
k0Q73RQjaXVvzY2qQWL+2ReaEgJUv51SEyzOtGbxsNtqp2KrAn370HmPge53iZROD47jYOL0KGug
1j+bI57eI5h/VGTP7IdSEqnQiTq4TKxMOnqsKxXXSo/Kv+qx41sOyghVOG6XcjjmpfTE4T2xMYfE
vqBNQ86JA+WWmJskku/X0aHqbI5pG1Ala1XdjlWNA/rQ9bmx9OnHadguTiyMGdfcnCKWEchj7JK8
L00ZqjZzzz0ayIhyBDe13a0aq5DCnb1DIMx3PJK1Tyh+9lrBMZPwKPnxfRi+Z1g84ySoDRDvQLKx
unyVafkxLYSFkXhhuv74enfEro87eyUXZLE2f26rRtZjTVTfh9erszE6lzxrb8I2d1gvTpM/0KQ4
AxU3dT6d0Akyi9+8P1hiJjGreV8rGcdcfcawO3eRdt6aitKW2xCxeYrHkhVj2awntzi/g8VGjJwd
Wb3tLfKR9X40ok6XosDWnMX6rCGRidCPXj6uB7RlzzrMSSyWAJ86Qh7Tq/scxB3jt7/JZfwIqjiL
+Hx59c4PO4/HGW3TRVPAcwyIC3WyDRuZAnBMtQ4RkBbuNGLQQ4YQdYqT9ZP68VDFGvRNDDS7k+1K
erdQ3xVU8qKOZ2/Jke/DENrqJ3nV3a+LLjH2u6tBterHQXcbkCbfeuWx/04dKsUiQBm0wSu62CJ7
jGS0NP6kiAMqBMcOwEE0Cd/BXf2slKwWYg8CsZW1sw19QYtU4QDA6+ydDu6QATiSzSJn8shls3W6
NrxMKxUJ5ECvz5TsXzaHgOzrmugPiwviVbk94bAmNi6RLpYpCYCfNcasvlxAnK6eUwQlWkG99fmY
cyIicRrBCz3KjBAr2s5/4KOR3WjkqNO8ST5gh0bn/sXYIICWqQ7LO37EvGyWS+McpytHpWJAlqcq
fqRUjyjNts1/e+pj04q+CsvU+T6b/mpdnYKEwdsdlPpU5r8kQ2QhYGji1mpwtu9jWwpTauJAytYF
vAtVwBJSasgPk2qaWpezaAs9+3lG9U8287cohWkryueyPTpZnl5FbJqTyTuO8SnMxhfb/wHEHy5S
MnHjPuXy0PZ4tpbuexgd4bSQ9xH0aewQJuMBEVv2euhVlaz4/8ZMKmJ7GKWsjSEded/R/9t36h3Y
YLpgIYq8JOW4hLOXH/XW1vtRvLLYyvEWOSjLKjRjDBvxnUX0RqfP9cKRXyZoFMW6RZ6O0JQDmyH6
anmnZpQw6QmE/tdueNGHKz8xq5l+QcsUmLgyhSO7jSTruDWArDgB7CT28RS4bd0CG9JXJ1RiEz6G
RsvkSzBMzIjwLoqGrPJGb468a0XI2hyMWAHO0aH5AUNaFYW0sDHdWpMfOW/DW++PboHiiaUKB6mY
cCxMD7xptC3uEoS4scUrRJKVzAe/8K2nScuETyCyF0nr1Q6Xi5FPo1Nn53C8rSsFCOEZU7s6Mrq4
smRY90XjbKQqtF/eoEztUBxjtiqAAA8ZJaCgLLid4kv+CiuXqB2YtMqeZ4GAKVZIMAaBsYaAZK59
+cNn2aVGpARurjHpdVqEM5IOJ4VAVSRtvKGm+FrZwa7wGa/VJLoQYqgavQsJjaqpIHusKGbcByMK
jk+ORLZAVWY8wm/SsNJ1qpEQva6Seycm3bJaCg1KSe+LfN0qcPMyapLZsoeQ8qJMYFr52tJ9TgIJ
1t99Xe9B2l6ndTIG98i+1j9cnoYkkoic2PAxgJRu9Re4ZOeT1+7KnuwyR3wziifubUHNuOsc7B44
cwS1JJXUdDGC1NnU4EdkZ7etPMl/2dmjPAl3qMNzE7HIcH52TqlHUqEdQGMv6bMzR5vCSyVIlhsb
IHemxZG+7Bv0q0861jon1M/kKzxFRfPJaTisHz09rfwGCBEr0XAkjheLTWwyfJDGSu07bXGqdKnX
apeZA9ZolRsX0PYUpSOeZoGhj2f5wQI4lNbTodwlz7qVG2SrHC6llLeel0OJ/wRrlSGrz5vC3qYE
KqCOBu85DPcFE/asUDW+gtNbjWXJjqnRok2Tq3JhikGx7vtp36nE2JucH/Fm+5mhLHThOALQ6FqF
f3R6B864xXq/B1xj6VU4WYagO/pQlNGgf4lr9MSE4jMjvSdqU70WbRHm8TY+f/ZHmNERmabwuvd2
b8hkTzasGu3qbezn+vSG11kYJ972pgaKZ0vVcgxfSb55vwD9GLeLGTDgMuddsQ+K24FtNqH4tYhe
7rpH/lAc2putm+JDGG0aQ3HRaOEREUwa6YfNM/4XsHr1iR3r8UH5LGNF5w7d72Hl5wZHUNruwx7m
jPbNqX2GDg0xwCD9R/QxYFq+wclr+PwX70bgvV6sunw+RbgD4r1VuW6V8uVuqymFt0pO6TPhC3kE
ryiqMTp4xNEKwUwtonXwalqBhXEI3Mwq2a5SvoWm8Xn+Olumw65XRVc/iyQJ2UU8Ifge31HlFGIT
Bo84zIc5yQrZ6flfjrhjZXLEfcRxUuDcpqBTJ1najBIn+v+sPP0keMqV99sGSJV0AqwCkVf8ixwD
WL4FB0LdNtDar3jRdh23biIwblz1aFGaZxT6sB55zbdYCGSXNRZUcS4mQLfVEw85lxgdEPjlij0Q
DA9lAEzakKPPHeFRbBSsSHV9kRWdDDUtHT3vk+hiNe5p96wV/hElf1YHTKsAt0zemCmNhrTbRiPO
v4QCX3QJmaPvMS7w9NbnBBX4Xkbzz9Xpl22qCmNILYoDbiKREhLiho9hKFc+Nvc3SU0A2GMnENNO
yfFmRJB7NlXVOKLMPCBmaM1cw92AIwaS+tFqedUYhcmYX/0jBh613ULchRpyG+fy0e54K87eLqbi
aoDSZO9UYDMIMT1jQX+z7NB9ro61nXspku412+kXWnrVcz2Mps6vBccBharzCxNoVpsbck6hO7JD
Sl896sdTrxfKnwF84PlAro5oYBCC47CiviZ5eGOFRKLmDGonUUbQqPDVBDFP3+2A3pmt5TOnxwqv
XwOTunTbMmUKLG7RdYRppRq1K1lx+QXDYsnEhQXmQysW0mIADrAceEbLX+rouTJFRMGNk4nmUVod
HWsk86mOlPtH+ZFJXK5tSgWT6OUqrUOlTdsoFkdNy7qojRvsAQYN0eKGMZJ1tdXMMkxvTcEjtnnD
NEdW0XoxmQYP/K2aEGmbP7YEHUqZfKHmPveK6zlmwKw4LVWQkGqHQ0P258OUBtn+T1ANcqQSDRih
FrENcA6TGm7W+VKDeKRoh7lTgLP6X8QoLBeeWEYznmllknrUOK8yNCSp34VnsWygu0gE97YyR+R7
MJ/t+l7b4DidCqjBVq+LH73TX0n49A5sJjR8o6OrHqwLKBsvB5PT+aO510v0ryT5URBW9RyRscNL
SeDv3Uq8uXx2bKzQR+ZjzSSllkGxukcSghaF8JJoCZAK51z8DB6EYcKl9v7QW/nS3PIQyyysOIg1
J7UOhkVrRt7yz9hMk3pRqX/6zfnXlE0Gn1+8e7+BTDuq/vR5N8guEo1NN785SFrki8nVKtfg0oau
8QxTQQ0fueL+SQ93lAR1ExJF0yIVdL6iNBq9bFfFobkQyiSATP9fOmajaElTpUYHK4wP7knzJQtG
gbJkQ9xA3+2SMlzD6qIWOwV+ZG+5qj8ra9P6k8VFxLgng3PJTLmoXIQcj25AmNeVs8xt2QJMI9G8
BgpTIZtf3yzWGPhg3fQR8VFYvQg7IfQgKg9h6QUUsLVW21Vg8lpjH4awJZJ0hzvqVGN01J4hUpJw
VRONzhGZagdHtIFcup3ZbPed5rZe8ybXHpYZKzj8HZn7jAITvlk918XPbwfc2fZaxvt3hbZZG0wF
zz9wEhHZE26V6FSF2Zb5b5TsibAXMSvs5TjAJdpcL9NEJN4Ra/8WR0d5Xxihy3NcAMY+IOXKqV8b
MA1QhQ8wb8naJKEIWHPYfuumG5vv6+QD8m9dEmEUdwD2at0jhzEzvVGprndTB4NOf3rdsszLL3Sh
IBFgaGNAAgoDgsSVknN2OMHWpaPZ56hOqBEIvVjlo/HVuxNmzVTrzBG1aN7SuumsksWR8xg8JKeM
YkGVKB1zlhxr7OBhQdHTOJVHv4t31vqzwk9bz2+PGOqLJDvLfb9C4VybxZ0Lw8iwAvBqn3TdhIzE
3x+yqTKN+GhVBBKwlK3qC0AntAOQG1E0H5yeES11U1AHkbI+IS/omBMqHfa1qdXNUSTUsghh0uKU
adMHe2U/CUSgFQGfFSqnOjMGoP3quZQzY8C7JPTWC6Y288b+W3vr+lPbIbg79FNDV/rinCF74EPM
+CFxVO/Aw+pTdUJGLKJKXhUPCWymKLEoLHvsH13weh+NSTNO3umb+EGgKPTPwBD5QcolE1hRYOf3
EchqoJFXps/gJObTsdDSUFZtml12YhL/2NA8pF3oGPvURAY9r/vzUQDs7Ijz09oUOCqaHcFrK1+4
TiA4sxqEhHDkSlev6f+/FUUoVbb2ne8lebCA3W32kzq2OJn+sntGz2/PvacR3zxTjXR6imKOJlmg
icrb/ac1lFGefKTv/GHs9kuPlEKVonmv+ez/+sxJ3UBhuaxBHhxRYx/1HH+au/a7TeEf2d72lxQG
PocwgwPAFNaGtns5vFDMzQMLriR03ODeLvqZHHcS/k5TwDF9ZCD7lKASE2N5p+53u9NZeCZt/WNT
jmMs4ebozmX0brlLnoRLDsuNh94BhMsLWzNK/1UEOPf3M9C1Z4ug76QppzBlb3qJRh9OUb9y44HP
WIdys+L5Q/v6RaWUDKFx+fpOWw39FBYZ13+zZpReipLDikdqxAR1BnN6O8tCeWqn/ViXIVur9zDD
vcZPl3XMkQzKb7QrCv2npBRSYCp+0RejC6nE5UwN2jBMVolWyBrKm70tgJkA+dT/tpSuuHVOyJyg
j5eH8aN133PB6PBjpofkiYesd7dsY7tI+jWl+Rt2+XIe/77xCltuDQVZ73ccBnWFEG0n4Es507X2
pGpkZgF9EMpWPFNZqc5J8ppGEIkYrh92FZ9c6PZqW69VOpywnBBr5xRKDL3Fc3UR/ToMH7mJiN8c
wnoTa6kpCqL2yqTsu5h0o4VouiGNdgILrceXGql1XojJXGvLUdePZqAn9j6Xp7ZYOlWNaPsN+2zU
Daf3NLaV2XnMI7Uk6TxAq1ZTkxQodZyKEwhx9CZ9N40bNhdDQJ+VCs05dvb9Fk6Js2ML7DliQwaC
nWTd/fe9eYWmsnCfsOOk7A1TITQEKLXWIVKCg8buL4OzHhfdJWoo4ttn4qi4BFLALj0i/Z5s6RMJ
Jk21OHN7nOddr2ejPwosVuEknbxKHVE3rhRS5dePGz7AYjjSKLIBgY9BPp6sLcYsI1hEeMOgRqPb
iet+OzCoH+h3gqTpKnZt782jMfD6//PbuQNP9M+EugPDu8tjFf2YH8u1i3+OpcXUf6XXTyArVI2A
NQ+D7rtyVMGaxrRVwonaGnVJ2IwS/dKWVSag38P8TUzVFNSUKkQkjL0kQWWplRSue/fTN3vNmNyh
aNsUfVncIm4A5sEJKN7OOXWL5M/CTdkDIsKeIk+tLljUIMCiEa/uK3EvnlIHHTERt4HhgJ8iK5kA
cheaDYyC0SSmMPzouqyj78yoIJjPuQBRzLlJHBGlXPA+Wlqmw+XJBEdfVj2PY7i1WVTPJLbqBeWM
myS2EVX+LMGoy8njTIRhKmgfiF6aQj1HNOq5cgLl7dL1B/Rt95fhY8IobnRZu+QKvEst6PMiZ+2v
CwkpTbEMFMi2S83LjzGcPZScxlwhUch3xcXDZzNnrZnf5xJKTaA1CKfulk2GF4f8SQRy87wNMEQ7
7cIg+laJHVrYIL9tdTdhF9USNV7GKn15az5NdLhbFLTwCAKiG471Gy/LORp8uE54zhZ9xJNFHr7H
X5l+N6H0NccvqeW1vbNf+26WspIINrr9GbTOLWNXAfENpTwsEeSzoI00RPM9fjkqNEO7/xj/WLal
JBkk1J5/6tMhoib4fG1IcIQjY7bUMAdtk4ITpGYOEHzfh9bbmOqA4pTKPgLo5alL5hmOMNmzC3zm
L3238kBqg0Fgo9w/KAZdsTQTgkEGO0smSIvdR4E/OS4xoy6tX9EL5Cxi4zeze1V5Cw4kG81pwnHI
7snhaWcrmVICWfl+P/pv6nRqbQSMkg5cusashTqMlikpqCwZeFhkOmh+Gd+FTlRPE0BX+n/e1WH0
MHKb1s0s+xCA3PuMlv3GbEDDWaZjn6E88guSpNXvhBGdsovAh+3iTnY95if1W6Xr28FzBBMxfEiZ
kG2+mfyZk5aOxPE6kuqqlRjFyRisirndsI2jwF3rdOM73RqdNmWPsLbVZ4m1/231BGGGxL4JmeEh
Ne6LlhK7fZZD7czM3TWPwenimlAOo4dHM1sGvPFzCnGIMFIDcQhtYhKpi7RpGl1duhOCnB95EpF8
foOdsT6Wz50lTfkVv230MqP1/zgrREiWNKrCHR2zVFMDRpVXgdDFV7hbKev3crN3HzGkUOYhn+5I
25hYXlrhJEg6BQWf4UvoBL0xppR1wVFvskge5rdguWqLRW0r1y+9VSBKYZlwfvaWAyd2WIWjdzFL
vaC9mtL9aIVuupH1zlnvnhc4L7GLx3BWtVAveRs0XgbQfCadorT9fXSc5kq/tj0yMcMHu0IG5Rxd
xx+Mct4UPjjKypgkanySaLgaD/9IvZkz2QNfd2tYaxS1s9sfBq4TZLrOVIhoEpnNKNBpW2Kbs3sO
jj3E009AsIrVvGG+S71MVoEFgvOCYu6tetfgiBVpQV/C7iZpeAzY70DfzoEjoKaoD4O/kOF23crb
SQqYsXVPrW1fn8bSF8uWYy6ICVoDwjdXihYTTpcPAVxv9moPWQjGK888ihN7utYgS6qTHqG4CCW6
eGI4dISWzr+wjAgTgWUcBDZGhBz3ktuAOkUD+fZqseSp6u7FLTcbhlf6NSAiL5euL3a60mni4YBk
9wa+Qelcnl15mggmSdrAcRCoGpeyjRt2Oy8gtz4IUGjwwlODd5dujxf7CQuR/41gkI9sQHcyRHDI
tSIxHj8aKhqlntfNqF4Nn13fo62We0P82Grw32lKDJSaPI6yXDmkvw1T5W6dMhNNg9dIO9G22dBI
wPyxKDb0YIklo4Qqqz0dJ6LnSRgPHODuEHVHLKdSNz9lw9IVgKBYey/i7tEbJ4GWbTcMNHv0y0H2
NoG9VW1Tcrd8bKu5R2YO8syFkovtl94k2wn1b+sMeLv1hbnRfil7OqeF+FRlP6l803xKeKzxrBsI
uEdft+ShozZ+KV3mtcx4oTD7+v8SDmXKJ1denXgBSPunVmvHobyXf+WhGo9etl45iLGoY57R7coT
fjhRbsHdnx2NO7J4h8V++igk+pmuRALP5+4AHp6PafdP+fLraqf8FJzuc9o0kw74uLISxtuvws8D
Sw/or3r5scHUzHhqv9tO5zOdMo71bUSwmFGaPFafT/ZXHJ4AncFJvoF5TZdGrPGbOpAU7ZK8Qa7P
uhZ7hraz2l2u/xvyqIDzHHbXLZYzFB1+Dl7UNZvuXWIAW0BMsV5rdRAkamoHvThpU9cuavsmIIsF
CjWFy30NQPfhY5yEb0xTbRmn4CANV8WRIocaVIiBdGXNAsMmjMqBfN0axAyWeCnIaTkNgM+kS2/c
BDFQnpyD/SJzgKSsIcQjGCyrmw36D86wS4/xwwhU43rW6tsYPa3gaKps53Vrqs3WD/YLblmGMEv+
CE76mgeMEYrHv8mOz9IXI9Z6W1KG+gzqNvSrBnoNojfD2q5VyBiFUL961G5SnC2qsDTmpECzwUqx
FAQ/NHpIv2Q5Iv9VVA75Rw75nvlS7v/GzVObz5HV3v2AHEpZDAvMZkkf8VeecsBVryYnJtr0RG+3
LpssoJWrDzKrTSfDYOMVbLCYhJ21wrLgMhGd0I/2mewRBTOcsIAvk2f0U2+lcg+CzZl0XIbd5Kiu
j7FKEvtSolMMrhvbmQVGe9RgEyiveX0zPTA/41TWOKCd8qQ6cm6ra1AjEOcYuKUHUcbVuiRY9TAg
3puQJxsCfVLTsBSj5B+pXf2fc/y0lg4PtcJzGLC57qfEeQoM7nzeik28BKKzwNHTPpybJ6z5HIVA
iRUPXP9ckOac+IRfuJXswc8YjnoBP/sCsoqiJLzWFUmaTPaQMZPvziE86A4cy1au3UC2AnTJwDA0
sbWJ/dGFvRzcGIYsU6BBcs4Vn9i79EyTZrygC2tfEG6kgvvSR++SmtEWiWlgZjhIAQJTbqrIQNuG
jl9v43rrlO3Q5p2A54O1OFy7JSjVl5etg8ji4DPUpK7r66M08fYSsFQ+QeyYqowiRnp4g/wK9njj
J1ddjI2ynepuVb35izY0NwW9I4aO9A6ilexY2ksqCjSFAKQkEY1qzDowUBF8usO0PEVin5c5F7gI
YwQfWHbdSpN/wLZcArGjYeDuK7YJfEy0Gc4TEfc3Kcj3kaVR7gXXcJ7zoV/eAUWia3HC3cqYT+R8
iymqaN1Xii8FmF522QixcJgonBPF45WPQjahK8d63X+mW/2CEmq4ZVORpeOoq84O3r5Y+ON8h6ul
YjylmRyvmQh865/WLSz6jCfD7ktMrlmKOdSddeL0jDuzDltfYO9H+aqmxkh508Zt16H8+i+qB0jL
CnltaL04s6p8RzbbonbhGxLoAM3iqGLyUnAdLL4/nMzMVwQA5idqNqyf/ZQacMR2JMOpHL8wKq4U
3FKuWXsryFqoHSXzRqPrcNmsmayYk6Ez6hdk3lDphJjW9deANTQ5VAUkF6swhVZRB57QrMf3Di9z
DYO4otuYBwQ7KQSKxqyHeddLoqfuhdJM3O3V32nsY9KZJLVf+4H++C5tYyhstMfMI8Q9R+V5JuoB
DlNVwM94QP8UM8pucEM741XG5rcTiRxslhAm9RFmcqs9RejUJRqCVwxx1FZJU8jYYVMIldSIrVGf
ioNyW9vguj+RWLT2iDWkyQSR1XTLay8aZryBsfOAddX6Xd6RZSClBJtDYNlWYiCXvjx8LijIxBNa
AzLsTZLqiO33oOfqKFU/8CQmUaE9+OZgr7w7WbpcW2AnF9zzB2BhuVjHXZb6Q2qPLEQFer/pIF1k
6HQEwAircKx2juACKegLa0ZbLGiGdj4pNBQSspyVEwp8wIFDUhwg0v6doJg19pJWRQamQHkac5ED
lm1k3QLWRGRbZ5OKR/R3MzqKh/GqRyvBZRML1U3oGFctFaCXMokz1mEfIscOlMHEAjd8y4P7EVmD
csiEp6Pl499OHDyuZeIvP2dny8NzitVx78nmiXjB3mHTsL7VoYj9q/EMbXdYuVpRLlhcHokJgHj2
vSf+m/YxptrzSGVPSwaFjshz30PUMCIV6xnw0dtEC245TVykLIt44JA2OR1IiPLr/kdMgU77UM8f
3/W0IDVBIB+O10lUfWYWT6aqincOHIVFHanFSVVihonq5iTuXzCKRmEu/G3Qj0V3JrMFedvFDT6a
camj1VAJy/nhuoQhGT91Y04DgGmPkhtatF3kx7egIAtDjckO1Zoh4T3inqFdXf9JNTrYHJUDFeIZ
wGAEAe2FJ4ZMe/3kTZkI/Nna6pKlabfgKlzVq4M1fn73CCl9KbGvA64u5gJcRkwLYTTv/wj4uW9h
fUJ9ZonLhAg/2iQRzOjXAPH6Hha9zRvDhIB+o0QABRZ0db4inn9dGuRiMi7fWQxtMQzPleV4nPRm
k0m+oGd7rx1hVwK/5rdKxPWXiSSyZrzgcj84r3W6NDyUFlArJfmH55fCFbN2E+yDWU3eSyFZVBh0
FUX3UPbwtEmy1BUGaMNOhamU3tKIV1SCFhzuyFqdcj3TeMVwg71XVfUzRAmx1OkB1Wevbq7Q6iEh
AsaXK0CcwRB37XGy5hXFnetBN0OyeC4bp4m/wH7wZyT+cjtFVl98PtjwDuDgT6tTgM/o5LHf8tAy
ged34Q5kZNkNd1sOWT/m9y0KfwHaTRiviIDb3yWEVN3u5SLG6ABRJSq9SO+w2rRMMIzNYunV2WV8
4MI6zzvYdiQVWSywFA8Ir7xcDcVajBdMIrzrFCfCIWeLPQFDA9VB5Fb9P7uFhf4moe9ssnUVbkfr
1pkcOjHg4ZUSviG8kv1plC3uIXFlfJNPFctkukSKFRkFZEgipDm5Mx18TsgIV+Om/m8gcH5buUWk
jmE1ERxLwbE18HIF3vgdv4PAySRv69Ok1EMcKCOqTC4zFxei+G5Mpig0l1v56tywDJSakF2N3EQg
r6JDQO45SmqgiVZRfAyi9KyaomXHe3f3EpitLRmmXJxTxaYpLbHEXP1X5xEs85qR5NgeJb6MxjdM
wbnlMLSRa0b63GWzUtH3m+BwMzziy9xySnk0uk68LLRmZ5k6ZkPbM1Io1/ymTw7helqnR2XSAHkY
jh7ZUKVN2/nzBwpsgbesHomB8aIWfdXz1Bc+sBdj60se2jmlic8YnSqSJsjrG4lEfP1QqNAz6Me2
T/tyVmQ2bBqZ70Hzflj6hhd2S2oeEIfeOi4KXW+svhD8cIsz/k9iPB2UQoUWBo1VzibLr1tjqek1
HG4s78xi6n+73yi6YrAL2Rz+NlmJbNr+Vk4QchomrinqfLP00oWAzZPqye481NUsEDpDDG7x0jpI
AbduXGLbCKntXMiM4CdpbO9WF4j/L9+CDSFxxHk6yfSUHucaHDU6he6znDZnC9832HHRbK7/cYDQ
OFCYUYAb/O9gqKY4yuNotHqvVulxREjIWCWyPsNbOLtuY8r0YCUziHeAtrPvolw/sPY58cJdW6cz
LQwZMQZYiLlyOoOJ037UnGJvWrTcRGiznba3Z54FjIY0zGBJBa3hxV+qckv2wDkQ1w3PuNgK/KS1
AsC8MrbxBFMhJ37BRuUYREp1PnZBeA4FNulBuJY37h2cP/1THsD7Pjj//fCJ7+GUhT8RVTxwoR5p
x2CBj/oKE/o68Xcm2wpSJM46OpdPsbJH/do4brzs26KootPdcHGnYfWPavkRD4sfTZvOxsgv0jaT
w6gAYh2iAX8/nydTaZ0m2ps5umAcTEcPQIzpgFDl2gU6hFLELkKZhiauWmpg3jp1c0+fxtuSnhy/
328WJJkId7RThEwmPJkfkfsf1cavnqbxKAngL1FcKLpZDYJAEElJCD3rx/kAM1gdzi99AxFrdlLX
h7lrS927vpcx95ycxViEPpgD7Dwj8DawqEesThA2ggzr2LcNafWHqtcNPkdN7DEhtiSdPBGgsz2D
xt1IHpJDJQPd/FVHLhETThfJYCe4B0brR/8sf2ERyqc1dG2qSGf4Qw8PO5BlKwW7pxngkYJ/0YBU
2HlsAlYLsoWr4xHJsw+LTqWqqA1NVJt4tB7Eg2ApHcr3BmFQKXMApSFfJrQU5OEO2hRuBDmnOGvV
kQnXLYvBrzLD3zZfAQ+unjlpn5iN1saDC4fY2lvScIte1Jbsq7ap+1Xk82jqfT1DEl0C+nn/kiBk
gtUKfgkwJ88RncDKkGHCqNWvaVK//MhMD7ISnlbdV5qFy8pbo15lsvqx8zoPfuTN3NWXNCy3nzRg
UoTn2HG5ZQHJxJ3hN1gfS4ZuQcseYL0IqCMRwju4X5H6iEZskxhr0yq81HFPH3uL64gsG6/EGWtz
CQlhl22OLEyUaCyHqIqHSk4LyILkxyrd9yPZGrpuT+sBt6jyuj1mTvNvxg0DpKr1xu4mL2xUDkIf
L/4RsuPgUMlhytXZEn/75ar7r2Ees4nh/LDDNOhkSkcbrouqwjcf6wAVvON/MMlZUfbOedPfAWeG
Fx0LVBrRM4VNApUQG9rdTiTa7fkN5qDMXsrJJef8HMW96Zhue05qVedVR2KRLO1CafBNZg4Y1C2P
RC3W5vAap1vN8eh9FbejTnzzaBw6ebTP/r0M/ds7AJN5x1ZuNOdWamj2iEFFz/DM2WsaoB1A5h1m
U1ZD1NLaXxSsVCyXr4RcaU1wt0FR/WpESDSNd9vNCA9KqLJYY65GDO0LcsJ9iKtv0cqWW2vDy6ty
ktRw5WFbZt5eDvhinlH2+3v4r+9FlnU+ANeVmPg9+aqmj1d4RM7XG3dcRNwdVvec54OyIfbYvbM0
9EroPeOAK3HbpKRlvUgaepzm7Ptp1BX9RKXZwMgxXyEUksuxgL21JeFuqQtRdMbriYltL0NIZBtR
/E5okDk0xuwBL7A8cGEiXQl5yTacjzL/KRDtjHPyaUBe3MmSM6p7swOcY9phDd3G7vmC+QNVC7KB
nL5jP9GydJ2PfFA3l9JBDb9y7KT63grt5spMrUoPf0yCL3dMcBVpvMlcVyjbUwMmDYz91XqrPaB+
YA1m6c2C0zt6Igf5bBWabJ0GWQw/21ilJkEowpTBwxSgxld9Cd6bsl0mOKnwOh1vow2UishSwkZs
1sL81k7MlDzC7tGRd2T7xiR5OB+O0g+8x3k8fna6za45kHZzIqHaKJYU+J43Dm23kSri7NvZyzcu
HVSBEW9OQH/u2zjj4Mn7bb6fCtIitjNm+zkwNtaB/52+Zm4+7bbrc4xFdL0I4Z10B0gpOWeEmael
I/EiLy5wVR9eitaaBAlP2EFg3Ra7GfDy1bb/m4CaYOmFvGtXLRh6865YK59ejYXHF5bMuws++OWe
PP4zkMOrTvt01QMEzdQlWJdQt51jPJfhxu7x9yFLyxFUTfhZJZuteL4Cy/agU8mJ05FYcHmWVfj5
v/eQ7gGyp2hCgTvY3+KeGabJ8qmCrFwGGNVsYfx3izX8mDuiSwKWRIP2PdSU8NX9Acy77KeRKz45
iucW0l575l/Mr3+hqHRUYpRxsvyUil3deza7TbVFJOfV4gwalKvXgHr9d7wz6QXNKCu/Uv7Ejjs4
ZP5YpE+2q6b1GioRpZj5pWL7M9VPPywnHV/yGiKUOSM40KbM5kmSb1McTg6cEedYK9o1HbSiDpnA
cIVSTuZL1vCS3bcqhYOFRjHAl0gNZ+EfeJa/+4oeRkt3NeetBkDO+kdVtjAVceKKEXaDEurO0cY+
l4VhpvIglgROyMbnrd9a18lCe2vR8G2SiQRjwMn1RmNoegVRxuDTGRLXysBNTILh9Ii9bqemfcjY
Q4+8dtR0kXuHXdTxfKTw8hjNKnO0HZQw5G5bupq4rXOBuWQw2lRHzaGZFLURspAuL2jXdAxzNRH4
VLBI8E2Y5c9Z2lUrnVQE+iWt9ncwNM2RFj5eGRl8kzV4Do5I0LLCoJXLb4uUyaQ/nLDKFFILaq8G
Pn2N9AEbsQEv6/s//ZMvPNUEe3qGJUwP3Hc6sKuzgDm46I0UFdTsM1dulBEVZRfEfADnJ0qFhhUn
TnbBxjvyDatIUxRzkS4f73M0ytjGNVvlN1wmiU8a37fJNttnXxK9hIDak67FW5I/t0ki9s/DoLcB
1H96UUG054hwiWgWUr39JSdUZoHz459fruOaZzjh6ucCAV03LOaC/wpelaMK93H+sEloKLZohSau
YwUucw9M/aey05Tf1OcOgbf5KnIPxLNxAJeVs737XnXv+Jdpcau5Kgx8BJUw/8BnycSCC/rnmsbU
HjJmiAlQVmtENabJXwKRiAFvsSzondJ3QIb8oGfV9rG+LQjVl7R8oYHNM1ZGbs+FFg4EJCVRWKxx
xsDfouj7g++JCGKC6BhZz4P+a0PfzdpTeava2R60siE/b5eNWcQ4xA6HrkFY+V7AJlGmKGhBr9rY
ynKsLptqx2h+PIP7vk0kDiA3X/75RNyD8tKbtXra/s+D2IpB318Vj4bYLNHgrK1BLPiD9Up582Pb
x5Tspp38hxAFceGSifqDk70Tn1EtMzZUxP6ybTQnRf2KBXCtAntPxSXers/BjdM/nNyBo9C6OhcU
o6oSdyXpZykXMy4XV1CE6iRHt4Y9+HccHkRIlS907bmuQYNMN0F+TSftwqQTI97Ou2iN5jL0eAWP
lsei/7/Y9eaSaV2WFmxiYw82jprGICQTycW5l3U6rFJR9QtjM0dH5naxDj4CTHAASb3SGAsqnlTg
Fw0wuIQu9mbA+DrexYp0yFZVNlOzXizWr0IW5nA0euAjuHXLjBg/3AhNU63mosAEWEOpQIuEPueG
ejlMewkroZnWiCzpvtzx4hjlUacY1wx9YwdjpmmjehOIgsLKttg+8xp/W3dI2gOOymEGHxKaOt0Q
V8yyc69EDWN/BdPkSxNAmywy3+P98h6B0gMcb/+ZtxTym8cgOf65iesL5GMuGWo62uqkJtK5qcuu
iF7RF+LLnc7KE2PQhh5+UKXw1l8trYOXYoB6nMS0aUvXiavKdqzGp865KBNEwVNzMt+RGxkmnvsk
at5q2BA22dQqMxIzxeM87aMxOMRSoiEgmHZAYGPgkYD+a8UafCHLUtm5hAwX1HTzhFwJ+mfV0H7l
wPsRfYfcyHisP9a50P5VpCUn9TDZ9QtpBtGY80fTNqdvtP7ap7yjicJuGxZ4n+LOy4TnLLQCDbZL
mKSPwbuodG81d0WWztEgcke7J/YAJWRP36NBUuoE/cLJ56JRW2jwbrYZYZqZhpbyKDbqlGscY1MC
Zglj5YH2yg270UfOSGIf0nqtFLiiXDvUAy55NHnXqkea6Tq4LFUJ3zQx708khODNtDjqwzc2wGK/
ClyYizJN9sYvuS5pphoxcSlQsVd26FVNGw1LBP38UPLoAo3ogFCM80gkTAnrqy1LOmvP92HMsGh/
hgjVvO2uUJaqfEGWRonNiLvt7laXHhsnAFY8YIHKjcq8/aqkvOtianj21gbBEQI/XIu9lFvQ6Eq+
VF2Oml/Jq79t7vyW04WUBIDvG5mzZhFgEK6RSwva/m5td/YZFNZ1eHEqAbzn4LAMkBd+lwyVhe+W
rficgufycz96hVaPrLxPXXA+fKsbhbuK0iNM19XOvnIsHr+J6b1bZg4FK8YPM9V/qVqoBA741MR6
1LoT3PIm4LhVenRrm9CcB49DFi8K7W1s5+ReWTpHlAvp4oPjQ+2cItYM5+hjjBPHVRAnpO3nLh7V
SyRYdxQCY+iwEQw2ku3XPObl4cNGZEyFCYfZJ+INpBzYij7sw9721IcDvRBNyYGBqANSXoEvEtGQ
wHuxsuCvOdPEDcnegKCY0QexOK3hMHyGpgC0aHFxStSPlcdl7vGfPjH3T0uUGF902DQwfhLM9i7b
JaZCcNmFxeKY/O9zFCXHrdIXofAxtvZMSKT+4aKA+nnnZMiGeUDICLNIHgiuU31oyf7NlV1q0mZS
An2AORBOivC5KdB0i322UjOr4e0QM2/P05mi0RpTV/ZNVuIyl9d9W8qBmkMDFHj6dRBP+9UNpaPZ
MMhN9pl1j7sEcIM7a5FOfQqIxZqFjlOv2A9jsN64PCdMVDzYjjndeLMfJeaYi9eIIdiD6Tm59vCi
VwmR4kxPeM98XbeRJeNOyBRjqrltMFhBLQ7vcPB8l1ES60cLiJzVhlCTEZMKG82xNiTxGozweZU/
ahAIPgIIa5SjbqzrqFDNr7XV8zRQ9GQ6c3TWZxtugYWNOtHGSo2m6Bt/DxLKCGPl1lPgKGdcMeg6
lx+pqVx54Scb7THX26unyok6n1Jfph8M+lBHDuWIWXIzNHgB0hj2gKFUexANWZenvYTecMO1vGCw
zcBXSIpZWFna3s/FVKt+3QPfvz2WKXrW/76YDLCIaKZ+4/sgTp5t8Ak+VYh+7XJr2WA0jdvK/Zos
XE9GrwXsEIxWgr7EigyOE35FSupOfeEZ6xc0EI6DMzF+QlDQG/0kxZluq1bA5TLtNFat2Km8lAZs
Fihv122SoJQpA93aEaHYCVFrgwsRSsuWDbIAIRzySAGTTRyhTnGVgg7E9Wrljo33HRN2oRoTjgrD
HNxiN4ZuCWodtGcLLMW676tPe8Rw8C9b8gkcShv1GCMNnFef5zXqov0Kq2Tu8d+ucDp5g98q1ZkQ
Is8/N+cDyvpehUXv91MJ+coMNJ1JsABOghj/Y0WHC/R57FAdueT0dHvpwKy79LcT+gsaMh39ByH0
+5rc3IpAil2hoMt6exdgdiO71gZgrrKMbmKyn1zAzbETy3NeKl8eYrsgA4XSCZk8rtxWQIVK0/33
ii12vpfTErWsZTxTXnzJHPcaIETWtdBUdrPqoQ2d0Uo/pjAdAik8ghQKosUHWSK0Tg/vFa1+yjWw
iTxVGOzky2yxiLrfG9SY3KK0asfLlZnyOoCo8DutQUV8l4CVgSyvkfH+cxXCeFG7WTVZusdMbCO5
2/iWM3dzBtS7QMMrhU8njt5niew6oxztmGj1xJ9ULB5r8XcAkw5koHbvszbgfq28HUlyneg7h0jW
Gpe5dptlcs+6S65aTLaJF4miCDtMxRZy2fO0HYDs3NVZEbRPxNQRxcRM+DIpU3eoNCW+1lbCk7QJ
gxtfvdfrctBZDGPgifSzob+ddwlcDz/8umr4QoDSNeEWz3diZeFrhvN9a4oddESoQ72VVLnVR4+y
Y952QzPmnH0rUWZsURz+sLCnXkSKG9EtBNoSoSVbHSEI8zlWEcUxOGt0cdxrj4uJpv6Dtp4k0tD5
GuCg4H54kod8GI+JH4OXviz5Vh8FVw+wuGeSHbUOPlQEXB9amjb7kPm7vAIah8BAeCg+tx5Dl3Zk
+9MXkbqGw0L6Zgh3HWyZ80T7zI3pIHSLrQXBO3e5ul+Igx2jZ8fhFrTvIeFU+z6zxr5BMPXqIQGP
xZJwBKhiT4bxqmUlGjha/QeSqQLz3Xjcafs83bmDUHGs60gIztMcRaQ9VFbsYH3YWpmZIkarW5WJ
HYvx2tUuPgsXKVtgcZcy2272mPrEPjA41O96BAdDXLO65/aAGe29WuMZhhWh4zE8w3d7tIMp+4W2
+tOwudXolY/AbCdoCs9azy51i6U/ZU00QyR6pz/eMhOn5Sx/CKB5avOSyIHkcimuQmsluanpA4zC
sCLFGoYvmI3/Nhxwkrgmeh5drTBKLP+T1qe8Zee8EDvUoW2egEbl8pe6ARDjvc/j+rHKvjOpwGLc
3K146cwI5fpbxbgi86WXNTfZ974sLkodR+itUj3CK1nrMSmIFa+TtMDug1H8jPUliMp3DTaIFMHS
620YKAceIJc1p9FGL60UC1b9sOBthQ8vlMltAeIPihBTObi4DPoRoZ4Af4gTPZK3xgMJhNFs4NJh
8HpZAegkpa8CDdXD65GKenYToHi0z+2ZiH6OkgSLSU4L1aqQxShuBBGJm9jo9r2nogzQhimOlw9b
ePMjO4Yjb6TxYs630v/WelDjXc+RM+CJ65Z3+C5IG6dAulKmhhanPJfz48qsjoO4kiKaSrVtTeLW
JlCmubF1GjPoAAMwgFdVNAowLF1XgS1kSAmS2/uXijvj9UOXMP2Iyu707P0+ivoM//hutFGONChB
nEZqAFGDi46Bh2kusDHXaXvFQZehcX+EaS2WvsUyLRhMb01Pd8UGxz7VpxPN6thjFxaSjGL7uCq0
lqD8bdZDjar5chE9gpjmHWzmWrDP/mGJOUZ1JAFv3EbFCRkYecQpoOPqyhEjzNH+R9wolm2+BqQX
3M6VnG79yMmqrtDMLwIOB0Dt3vPWVdSGqIQeKG5WaEzLKwkAelrQ520y5dBWKrBZ8q8mD5J9xQ3g
z/xkjwMfZE+l8Hh68FkWFo7UqyBqcbTDG+YDt9VWTsYhM9E0pa6xoY6EcIYaEM/dCDplIEy9TNQG
MrP0uX1FlVq5acauUoMOHNQZQFBVTHrLNx/2uIyO2uNlIx1EKjqeoXePBqFMSrjGy0zGxhuplLSq
1J+rkAlhAlnbSIdsT2fzGstRvVRfiSSMcTvkw+A3tt4+Sbyz5Hrv6zzPCJj065nSCU9bsIyLXKhm
UtTNe4rWMO31tkh0cgUOGqq2BJg7/lUqE4cslrIa6lgyid3j0Vo/BiZMclfsvD49ElTIdmtc0pZT
GKLo8OJcBamzef+85+NGOlAVjMQ/CCRJykRuDIn/4RQrX/6dVLUICh8b/yPlW+k0wi2w1R69j6Ca
xwsujsT7yTmkNhWwTcfPPU/MYswkJXoNfdgbwwG+3WEAcfEeWE5KWrZNpKD4eaojPTSSiJWmZQmk
ViFmOU98cSuPYOoC8Pd264J2x9w8mLpQ0d+Wkfvk4xtETVtYDbiDwQxu5qcu9EU9GNXqeBfHdAK2
6y6E4USea55iVMFPAf4xmeV7nxu+bvy2MHVT5EWuVW3Q7Bi/sBBgsvWA1rHbgngnrM5IjgxLUfpJ
DKmuwOqmR2CuP+4MEqammH0k1pnc5UT8HGp+l5qxRlrnn5sdE8GgtQ34PnSg4NMW7sYfjbNdoepO
mNIojdJcJ/ICBzYN+UZCo5fmHRo3Y0jkv3KkAZgy2FqeMJZFe0TnF1gckP6QFzrgZrDviN/1umHh
90KoI7lXN6wuqMZ5sVU2rupBNa5i2nu27Mz+1WdYjhs47RxYCOlBqLe+ti+AI+GFrBSQ5uQM7iRp
w097UZB65+SpkQMLDW4peZ2mMByS8AADxSa6f0cTCRtqBkDPVSUnCGAUcDSiT5QEAGak1wV2LkFr
Lc3eZ/vO3N9W6p+pmyVaZwINy3G856engQK2e7RvxOcef8u3yPlYafUpiHn45DelPFn3Dhuf9uMw
vzZbQ33R0Cs4rNeOTUmdRHfIISeAFcYF/5Ny8SwtWuxMbuxvblftAB0M8Hxs16Zaj5NKIiojx0Nx
w+FLTQTVFgHnJTphA41EkvJ/ssy74vx9MF/cdRq7wARRYAlYkVlaRNA9Qo+2okAUu5/nFPUknTLZ
vbul9gViEivngbPBuyOhPwS4ip/vk34D68E0n/MQLrc/LznLPOVwPswDuQ7Hq3tAAmxXYx+FK3hT
1g0rmYmqLiKP93x+g/cgG+CB3U0PotSuTNJBK75vqQie4x3wAW6ETqpXGfdt45ql5LW6FMXxOFb+
P3Gx+xLC4XjfvYawlm5yNP9w6cfr8wT0hlXoFbGb7gl27E0X5TJHQMy+9qeEKBUr9bu+pt3h4uAd
w13Jtq2C4z9eUJoT0FgBZVlu2Psr/EeQptGRFNEDTq5yKlq4juxYQkwpw6sli5ObGVCcCGRQ0mVL
/2p5MpuWoianVrdfZMbYuEu3R3cjEan17pRSLFfE6vR79jwyi4UDXHpRvp5yqGtff9zvsiglNbqD
0BIH+14wC9vvHyhgVz/tW5R/SJmbgc5zQ+QS/WjJqQyCrZVYRaBucv9e9jIp6Sr9ft/dG0FdhGgj
cP/JdEd+a2jE7Ci1yfsJ0bJJjonSp/Un3sxv7hqzQyP787yDQBHB9AQdknmGFlt7AL7gpeCyerFV
kCwTOE/7FsnatqDoFKl3R/XvmLFIxlmPSnK9hFHxp3YRtuiZ636uRX1ZNmvcGwhyf8SX3B7bvXCG
fTVrynAzcUIgv9zfnbKlnrofFDBf2Lc4sUb/jestoJ4zS+F5kEKNoIT7GP0xfarkmB0hxv9nGspI
i1dniAGQEcgyOl7OVwtIdNIMS6dxaNe0F9C9meoG1A+Oj0GjyJ5jQevhjcGomu+BmY8S0JDJPTav
em3YniKriJ+/qC3wZuUlColl0HBofjvDqJtqw4MJswLeWG4iBzlYtlvBirJeust2zRfxrXdU3ZZy
5smGGZ9kGYqPLrZIRAnkMoVOAxz0BHq67ky/PgetWq/UDRpmDDcbOiwTk5iDdOm7JR6WBYuBajsX
M8UGMCDkoFBnnrwCgLTatZAt9QnHjaKPx8eVd+htlRILLBfgbsXF02Q5XNjf5w5Gc9d5/PhZxGjt
1Gmsxr7Y/rbx3TG/xyx1PQ+jp+TL4lr88fGIR6ATYHfCB1WgcCBDYHReQLqRhJIks/UQaLCPwMmv
p7NEq082zgq+1M+4mLgWjr4etffMViJMkQgQuZ3OOe0J7UgsncEOrG7f7od5VuBRtK3fUcW46xY6
XTsUx3FbNbnVah5kGIdj3+voGsNMyvYSa2i7kdzMZgK8QAlCfPbJ8hOsat29BsYkL1Bnka3qX+uJ
lgicUIzVBTZ06jrvIHAe9khLNbGKcxkACxnYQWwq9EFAENDA1QUJtlaO9WkRcOd+lvcCs+R5ZBsD
JIzF2T9EGJchdp7c87RNfOVni2gVQ3P0DklNuvs/M7lg8VvrRmAINMPD0GBhUjtreCVXBSci2TEY
KuCqwqXWxZpO/lwu22rbRrU8QplgpfVNvBo8J8k7XUAObtqsG/pfc+fO0jwA0sEVkb8wMcUODIyo
sIPxztZehjWWmZ/IRvHNkhYS0lur55gv2r8n14A788y3M5FKHl3qqGhcw7N07jwlfsAHeDtDgltB
PEMiJGdzjnj0tfebNQqoTk91oRtzCJDaLVC8O8no7mVMGoIoHLzzw50pSBX2PyOcyhtpcz2VntDn
1Rh1+TY3Io+aYhHyNMiS0jukfYcFuOd1RYe/RPeP1UB+n6I6SE17RL7gNOJMGyOHnEOv4/FTuEzi
DA4mgqMx0ycxiHeK99GNHEflLGsVTa6y0M30/lHodzMbXk/GxWlVt2gNwyndTis+1ynlz/WFL83Q
YycLAE3AU2cN+eHS+UOs+OwJg5ntHSfP0R4ayLK0X6on2RPW49S9b+7XILzbkSAj+tEgXe69NjNa
abUdgWZRJ5Pi7HOkipD0Kwr3RAO8ojTH87JoeItZojAj5IaueITLVeg/l6Ln9HLhw68kFcS57cGS
xbebLoff5uMLHEfd41bNTIVh0Bxpxqe9UVy33ae/kl3K5sfOARqPQI1tCEQ3C8vDbJ9+fuE180Nz
2jouj300V9JzhVyRcc4ioxQUMyTMs+pEKbMns1o+tUlHSIlAnFYGgl2MNaLVriiNcX7VxTND/FdR
DP8a7IrEdLF6VGg8/CZeUSWQOrcBZd68Vv3ZxDm+KBDD7EkLFL0ZXtGSChTGWV2qgOIoeXWVUBlB
3WTXXHJZIB9RkmdCqOxN4V+XEKfXVfr48AEZfF0ftc+9+KtC1nP4ysG0ErXJIOxdX6gOVI5XVM73
k1JaX87a/TdLkqEE5sAXWldbx4Wav+rmyNb3nxPN6nWLTlka+U5U1+mhPm6hq0ht4FxUnQud5ono
OnICEfjSJMmqT0rJx2ncUwRYG7Gqt7ZOLfdOIZQjs5tM7rmBrxIEg6QJqcozfuutNraU8y+29nqt
WMiS0mihCtuKINNkYBzTYbLDtpKziUlV6MTKeVbsg+5DcCa1n3DuLU2jejDZJLHKliV/xT88Pc7K
0hc44DZVIFksz4nsKV6h2H4gmTfV0i17Nte38+/lXIorp2m/4ySsmOmTXMYD6ZrhREmHmu7oYv56
6IVVKIDJTsKpQ3evfkqZ0YzVoOoPdcJx9cdZIo3sf5lJnPThJfPjN+1tdo4lP65VpTvzS8ojGbct
Yz+ioRs7Aonvz4oozFBJ5iaidw+p81kao2s4DG/jdhClIJtqLAwOHNPD7WmPB+SZzW9DR8tPYdUd
U9RF7BJg3ugQD0K8SbXKyD2s6JhjDyKfmwXPfPuzrj0CgCOIwTp7x5vStnG1GSCI3plWuFORi+qy
3xDmsPZcCM3/H0RrCVWwXyDT7W5hXLNnlU/J4Y48gf98tY2iGHIJvafxDqEuvfijDfgPVR2wyWAD
Xz7u3s/R6sWqYc9303zFfvpAFC0avemOYgIbSsLyZEJ06zCbaAwTMjsDxVkzg7BE+2STe9RXxOcx
wFvCMXHOMiFZo644makyfafNgySvkyS5P8ajXim5PJ2yMf0BBdGvLivWHK9sA4nJq9s74BHOlH8/
/GAte8YqsgG0LR57rfeQxlSRaye6fNEMAwiAFxNSlREp64WXCXk3iyTk5rL+7IIh8pOufDeXaP2i
dzzSxDKICCVVQojkpRDHafWyIbILSzHblUpk8D9ZK8JXUBVLGKjHufqjn9Gpud6ChICkibtFVfpl
Z8SCmGHBXyuzZy6iioZBq/xXF1eU89sXdCLuUVnFQ9qKybPeXYxgmcsFMM9SpOBQb8QhwVEu2/4j
uwPtmdR8pLztfOXGBHPot2ymEJZRxz7BA2Fz1+zhp5qcERLIUTTFFEG5Xhu60rznO4IvMrp4dNpm
ibNYkCQsBkAQnVsUZ8urxUy5wRLBqt1Yd/Oh8zA5ypi5kPQEROy7HzjJl8n7710O0FmokAGdPiHN
0aj+llSyU+dmWiFII30NqLysneEi11Lb3c9NmYn8jJViOgVi8Ya3teN/tFybWRW3jzfwc2pCxQ+T
sEkQ2cbHJi4Qxi9OlNLg1zYnps0sSgCh6ZBmsVPMX7ltGYm2GHTEnLQ4v09LxCA5IXiNbmXGID2Z
mS2/wpPUn6LVzmeY5wjGvqJTyv3zP6Ve1vOjxJFxRW5ebjVqaDNsM5I2B6Fo820Hvuo053Vn0nrt
NmAhA0VT2hehll7Q1OiT2nDUOjuSQf6NQYic6utt9gFiwO75cp/tfugs2KU4HM5XarEdHs/yFZ6w
/h9z3wbHe04pWkcsKaG/qWrR1ttMEoNXwh38vZ6fOe8P+8mLI6puEUFrYHA9DurHUWUSS4xqA8Fj
/YR1kzYp9U5jetjvz+PwJXLTdg+lh/XVjzhOn6EHeEH5cdTYHsk2z+/Qwt7zqxySQCEVEeP2NRQI
rhLqxZkSOsFcWdSvBoN8Fhbfuu+f+HHYLNAI2FHDrqm7RfaVkD0xdSFifDa+J+fpWqp2sPacKi+/
vdfZOCizyBsIuUR3Iq8UWwrsygCY36fxaLOe7jPB6z7rMbeDxselLhaVxoz/AAXjsFUoXVnT9Nze
ZoR+58It1il3HLuw/5nkzHQ63771wiGSAIhN8lamqDROP5PnIydBmv1qj+kXcDofrpnxIteAzwxz
oZw7c1RXpOx0sqwPdU+WL5oGB/6zRwAiPf6NXA2t/rdz5NGeQiCK/cHPlpVG4tW06E9Q4eEjK4oZ
4x2mg4HoCqJoSPL0ZbOinWI0luaRagjVjSMCn5vKBMKq+IVQRMHAI78lM7+7p+zuCjiOHz3ajz3+
a/W7WC+XZCvaAMCVHrXsPPegu+mKVUIxaGPVqpG+t52A/Dm6egrU7CGcm5KRK+CgEwDOGSa3tdMy
B/of8Ri9WDokhiMR+sJB5gVg55pQVCKIINfvgT95JYOtyxYI3dgb2uF4beXTWHNWfYO/wCkNJt/s
JZzt7PdJJHSReb3j7UzfAifCkvDpxXnxyqdw0DuAwMLBQNFCVLSCmxI+qzGAzQOJYkLk+Vef3of1
1Ty4Cdidtb8RhdJPl/X/kP1ZFMWK8vbkflk2xifSNNOIAvSt4RatSuqCu2lbhUSVoxc79048nLcD
/44xmBP7Q9jSV5YvTrFSDY8NuOGS1OriMmnlyT/qywNt759Y9Yape/R0dni6cv5yKNTB9uf9aIBf
J3lArefsCQ4DZsnjUYoO3Rp3PQSTDi7qvq5bv2C3wKvVKQh0ODDq6K1G4HHJbws0PMvZ5tT/Nad8
q1vRJ3FvTSelbrfJJvlaskmkFGoDCu6Yh3bzslMevbhRwyfcBij6whEaomzA0sTsRliPUkOkj5sM
UB++ibDGs1+wFrJgKHHT0k+JoD4EIbzf/AvScy8LsZpBh0zZfIGLp8BwIsL0jilKYTq/Pg3DplrU
mof53CgsnRKM+LpYMqNtuUVgLOn4bx3uszjlaFqFPyafyDskQJJxC3LCVE/OsIwcNW8ym8rAgyMO
xDkAps/QN/rpy8nj0c0J9Lk3Dzk+oTes0M1g0ILoeMTg2erRxDkl/ZQQ2bYps2KUP40NV4y9pc5Y
/Pt8yrtS+cDN6SNXhcKLPjEvpI/u3e+cXcBX31nhKzH17CQB+lfhasBTEqNuBbm9XFl8KrQcDa9g
/MGxjxhW79ZLqh/ScnhtwpMyxf1QaQh3X828BZEYABkFTGGcN+dUsIyaqs/eAUJxt4QgWVYxf6ZT
HQM1WeaBsczQfAZotSVb4IWy/6+WHhlPE/v+bCH01KTOwkxXDNvuMeL8WthRurIdSAmbxBxMg2uO
LSZ6Ho7abG11ZI86Nsvi1bpFeNqY7zGTB2oWuVsOMNCfXYuoliPKPhATK3CfO5XnEUS7nSVO7GfJ
EqoA/Weg7WBuQx37DznFHcJar9aRGAnUg19ltm3VD/PbZdJw7f9l3hl3hsjLlMLV2LHt45V6eqjH
D8siDZHnPcJzXeKhWJpUv5EL1v9NnTIIAh0FjlTcLxB9ZJxiVqPsCm/4uSncnxu4AgrMbiwsO/3R
FE+b5lAfyxn0F5FHtcTbWrmf8lBo5UTNsECz7V45cZGe+fU8+QCHUCJXtaJFSm7TbOKPNw7ONQ2C
6USu9FUFVZH85JJdWZ/O1sst0vr6H7FxrXQll0JmblL5fOtWbPHyYxWT1DePi02UHUZBy3YpHKyD
X3JiJDtUfqPWngT3iHuzmE3/kIixkpT4EYdE58iwJYxZEZWUZhbUBcU9fUI1JrALA30WPdUKQNgx
HwtgG8zEhR+K1sQ8CubMHJUq2TJewK7dVwhoAPra6NmFFfL8ddyMkG6flsS99y1GcqEgggR3enK3
PBecHt/E7sCT+6V/DBVaTIxqJwOKs+O9cYEanVdy2J8gH+66nU94lQqDP7ExHBwR2qOAsatcNWYk
6vJJfkzj+IjMchOyLPH7C1cRYSq53g8YtkXyvgsJvo1tuyzYRcSPOCyzBPEerRc51C6g4NajIWfV
0CNqXEIgQffeblPjs7Am3WeWiICUlR8rk1UQs5g2KG9B9GYfK+tQv5G/gSmrqBFHSqenyJN+TxkJ
wXDny4CGNgYgastj8+dtL4bHfKFBP6Svs0v99O3QOvED+dhje97MApJIcv/vYrcqfvrbfDIlAQ9M
pr91EaTB6iN3OJ/9nE6EKvKRNsZFoifJ2kiMGY23M6HQ8qLXVGXi+gjLGwtR+LaBYy3MvD00mIn2
jAxPXtmXQkgDZE05pdCXEjdYszdTLR+C9/SojPgcFPH5VnlIoonC3Iea6/TkBUCBzlaqjRrp3sim
g2RRLU89a2DHki8l1zUYxVIVazBsNVMvZXmrzbnCZWU6Vx+wBCNhQlx/aYuH7gKFwQ20UILY+DZx
ODEAWQ/x19kh73piXgvtomKrfsrp1tKMweKoweTuNoqwu7090xZfk/klbgIlI5HXKb3Iq17F2GLz
+I/9+2XnKVEh0TO3qTzL1YPPGVmnn1dBYk3eiDvJKqlUC5yx/if7elpSoJ6EdI8ljeC//VV+y4Vt
ozmk+gt8Lz6rpxrvEYPamD/wruGRRnqRGIPBGwlNGrlpgrkiWPy8yrkSmaHTj4187ShZnxoKahAl
Gbrxi0i5QGGLbDH6gqp2hv2MnWjOlifPUJfF76Z9RkcRx71NVrSW6pNU30+qMAUzoo+bBdem41WP
JFPEjxG52zL1HmrJpUSpWq93FGEAA3xg5niUwmzymdMn42GYXlr5/1BKAq9gQVEEzAjUYcwid5SH
Icoh7hgiGBUXm8dcoCJx1rxq2xXONO62K0UFNV/KPIitAjg8JUMz5CsQ6zRtEL9ddUUCgnPwgW5V
zGDW4W4C0gtQAhOPtRfKzze87r71VEVeaOFXHTMdtqs64d2eC4R1x9id+oZSOJ5ydfcS0KKjWfsC
/4thHMadazq8mk6OOPGEI6lt9gvjr25FmcDQtrDVPCJ+BCmWJ4+ZuwatK2t/7ptLxqI085EdojHk
PuIdE8HVgPRqdr+AbJvbSb7TBm584kq4hyKkgksMTrox7i+/D8Yq+1UKhP6DvefYeGoPvH44XiUO
hf5lpYwruR0EH0W9zZ2IeapwrfDP1ETQgvJShO1a+0e5L1+lFiJ2eTfxPaLDNCf5uSv013zQA6FY
UpVIV0CwjeVSVfsq+qyRXpjUVHKZWzbEY9ND7NoVU5Exb2AcvcInRvd0UmNG98gGQTBBfTljNgZx
iSZdTGwCV7f4Z0b+3VnYIdXeq6I5ct9pukaDRPWNrxt4UKtx12I2tJo+tvpkNm94QmQRhjs2AszI
wofLPOmP8LeL48UWtcyj6qUNOeBeQW/c32Xwd/Gs28ftH3kKLWlJJRhmFhXpt3gYLTE14igELWEg
SJS2vge156qX7JZ6TIISpQaC1NbGEnr0Ufn5DiIbcTteoIovDDsA1zes9w2CH53MhZm8N/GOUr7Q
lwVCtxOq+VadTJoJJhOEK8+oBIV0Q+3VS5uVZ6HLC9VhXDfq1TPVnQBs5hkoUTPbvHXh97mylFdd
RtgA4mfgNz7eV0pHRAjYE4nKts8LMqjiV+0fPjMOMV14Ia7i34+uxmAmxiDM5+DdrF/66aHkw/BU
tJduX9jPsx4Mcl9raPgJlMZlcIfxmb7k+16ZkH/2JyxWrGIFygLVrFg14hfFM9xJgdlqW3gjhoi8
ZC7rJKE8SCYbixIutN0z3fOSXdGSpKEU1W/bp/9rlBZQ4wMQFbCH/+/7i6Lpah44wEABtk4y+OJl
JXVB59cuP/kXfLAAwzNkPk0p3uU1kO2O5kAjTDhzLHUYHeuuSGvtkv0d39EuzdFX1VGCOxpd49Sg
/inDymjmiq3DZYuaynCD28IVXfr0vZApcLA7YKHxws/wKPAxd96jy1Ix9Oc7RwhSkVanNFgDeMAe
cA9Qp8J9QTCOs4ca6LgLff2xr/r9oUJAursp+WEfJyJm3mitEpwAm11gFy7RIZTVDJioE+UdgwqT
3lUP/yq+gIR6r1+8kySfP4kTiODiiQ48YGgLpcdc/sGdXGTu1T3T4bpFZCweBgNOC9ybR9vBjqQm
TbjMBzl88qZQmfu2tQqlmkt9sie64YYpwKC7FQuw2F8wbvdL6iYOJUErgGrvAHT6wK0c/EiXhvXm
iEN2g9IJcH86JmSasG4rBqryFG4JzuswYM9mkloVAxFIJVUy9oWCASpYT8whwdzgk9KUYSPOO19q
e9hQK38je4EqSKBnMXMi7tz79xmHBIuBIj8PYH07WHruJjV21OZ6SeR5U1mlZbl1S+yMXDeTltOD
bFQqnet9KwH5WxjWsi+YYzRdXfs8aJLD1WFENhPzdACjbDpKUq0kbTVd6nnuopbscK6nj02qZ09h
q6hqGNYayvz8OT6CFTGNIfqUL/c0mGbfyBjAZIGg9kLI0EmWjTNlwLfduMcro2UaRQGn3FluAx1a
iU3cr0Aqw/Si06q5gx2imBqmEMgac+ehEHZRpOS8YqAg4DN8cbXXsoSvVPFRzP3rGsgDa96huzLg
YwvLZlVYUFbz5vYJF21eWG4CFFi6iLCW5+vZzfsee/+rKOvPo0M0Co/8wYjBx7Ns/Ky6FZ5VDoWb
0VhPWDQin+VFR2pFb9pUR3hWoFgw0JDEnmEzbKF5wsUdd+S0LrFNQ4/wY6OdUGrl0Yf3QmYNF60X
nlHIeDKtVVNITXplHw5Tq+vb94PSIX0FFsiCSoSmjzyHEN0jsvIfXO0d+hg7PPVdKYxmsQ0luOHs
UYMq8i6/na6F9Gyz71JekmY4qTWNn0EtDc2BXAqG8icXSu7wYb21o3rC/Axa9lnTEmipx49u3k7x
UPP+b2d/Y/ERH4KvPyfgPXWBznQHkR9cezL5ly3O3U31Y7WueSOFJ7hqY9gb4qt0UbEquK1VFBqp
EvwugUDEjuenQdye2wFydM9rqlrIVmj7N5sHLCBUsziLNWWqeBUiJhLwtnev7ZRnGYkzdpmdCLxJ
h4IcvYlEB3g4IUwyQoMvfU5AbepMX28YDngOBLD3vTpqNhujciXCEO6Kyp0kc6KTzgOUvj/EntUd
sQtVD+sXvzWcAOVJz7cVi86RX6RhEuTNZILlhm5/H2uib8nj8czGlklUG+/NmTBMPUqRU/VZG3rL
rXp7S+VxL2qiT+hv9BpxR5y6k4zdiXu5t4lpPEl0a1ty7AlyVd1UhGJpp4TZ7tBQao3k9W6pHIDp
wJjnOUOQl98J+QM8dct1F7U5k5G3B5dfxykIsoIUNXFdOsVrTGCpNHZtjBynQgvdbYWfLKo/gRpB
Qf9DY5rMJnKzginr/kJS7AZnN+dEm9Xgymmkd5gpjRtUlqlL49q5/EFX+tqgNWzw9Dt08enjMcxh
OLDjrBDuVrw/07jHoBQG7qWVO28+du4b956U44XYwfI2KlJOiigb3yLPQslRJsZEjBergWwPBXtt
65gPMRvwBYpBZx/HCIiK7hfbEoyNlL69T7wCWcXM3Co7KD6YDMtLCBlvhcmU2R5XexsWiKXvv2+Y
wrrFpbfGW0OkEGorZk3w82TfPGFLkV0Wyqy5GlZVTy5+F86gL/GO82XB1KOUYZDtORykXEju1SvI
Qi6Dvp4Jb77SyAYK/bvIRDRBIFvHlnp8ht2D4VRs1E8e5vRwLhshJj6MUdfh9rti5Y7vY6+RMEey
qoQ32BkMobz1G1Klzxnt4CrKQuxG8zgIab9MPYyCqZG4DzFjaoAzDuv0poIS5Sa0cBLuwB1lKYRe
9FOh8usQvwKrA2bL1N1ZTvHMrTJSkuOHBUBZfVUY/FAmgIzJGs3HWAW2Zwz9cX24PFfptvP+NTdW
wmmo8EQlGN6peWJmbcQY5prAWzpzM6y0HoGLCmqh+M3zZtWlT0XGd1Qjd+sV1fi0j6zIfPZrmJPB
KCXzBZ8xtgmtK+OQb62/cHD5PcsPeX+k2OjqU19ATIxobMtoh8TldVPqikoPX5xmehMqlZVqwx9Z
zazma0T6l/07wbxMjWTfLQcz7ZmjeDgVd7alxMjFUNdX5BcyzHJ5NOXcF2ZMHgC5AQ82Ji/vn8AK
Il3b//0/tX5GkkaQFwOkvuKXQy0hbIFZ/ePmcdrrbWFF0CJWzyy8mFe/NFviyWaYW/7MY9drtTAg
34DKOOO25fzytNZfIBaMH8DF07FSJDe8Zz7lBKXIOp1ffJPSYNzLxUozLDFPLgz8lG6P1/ZWPtmt
ffv2SyKLl0NYdrpYEfhOob7aNYkdQ7y8aAt3LJcDzVpJkn/+NkNmoJlTY3ooccbVTxadrsKlHxq/
mCvzeAlim7gx/22LVFUXj+XG/N+0gLJEB+qy4KYEPbpHivQAN4qD+oiwDh/dgqHO7Ce+vYbwyaak
dL9M/MhXtEdBy9N4IehLlMKlETqFms8zSZ6TF4dsg+AF5n/xBg/jx8Sjd+hDggqDC0GpsIq2fx7P
MlmlFRmrCrTQZqUtD08A1YTP7xACJtHvsF2zfUBhO94QvPE2QyuTZja2SsOxQRX7KWHzUTbSL42f
oLi2A/VJIUuJ2JJgmYJVp53ejvKT5e1Iz5Y++n2wDzEZxfNFmhTh+xPUKbFEbcFEyTC8nvnOSSfW
M7TeHTXYe3Tv1iUmkR6ONp1jIwJWHsp6YGrvUaiXEqH3H5dYqBkSbjg5Mjvpe1cXPXHiaxCAcA6i
gutuN++A1n74WgzWNQxJiU6NPRfWfLzjFiRKMevpwV+KqZ01AfoKF+dqELR97UsHdydCdsE75Mq/
BbFC99Pp5eUylgWH5ltvPckwXgFHCVkGn0fHHN/MLt/7PmSDiRh8Gvte56ZrtRF+rkSpV8D78px7
u0qWRACTqWU7E7qnW5kuCHEI0iYLpgelKRgBFBzaHwcnm7XrVOcFKUS76HyAt4OgcmZUFYEl+oSM
TXwMakPt4/6tPewwXofeGX+YWinaGyvOcZO8Qef1wzkSK/0scvV6lL5mO6UGFNUJi324AzzcLpLh
7acSqP9XSfbq9Va9NGaxqtTojau98TsciLKBMKmUqCbeTiBD2A9fC8J0KhRlGQkwZdjk3NOj1TN8
UKcL3QTmCl4vhLt5liuANvc+gcTggdcLNYapUeli/CqmX6U5DKntz/Az33/cElnFaMaCit1pl+It
n2Tt+kTcJC2QVtmp1TPnDEIECM9SjLazHEGtkednLXKKSLVrT9JfreCw2fCFxcGxwd64yYK52nqx
5Iy50ZyrJdS7vAw22CjPxT6jBhUs6tV54xJNMmPhrcFnH+GwwR6k2K4Uff+i6YM/nc/mSUOG95kg
I5EUbd9nz0VMBMTKbNrt3iQrtUTWZPUiEdrrXZ1G3YRBR7fHvd9Emr+z0Z+wqSUdbAB32ayir4du
l0lCD4VbDZH5okdU6/IEtBidNOy8ikz2S6UKmyOCPhbwcqqbJygzF/ViC5oQJbM5hb7e2BM4Sv58
g7BiDTFvo56Yh+0HBtq7SoctZcr7W7Pjqu25f62xSPhcJ477tzOM9j9Bh/xJgdAezbaJC7pdj3/G
ScdFJCksLbtQ88Il6HiGsMtjZK7npD/FKvj/Nd8zzdUfna/kQ6N2ZRaN8EHe++NmOSv62G9/P90t
9ahQSbagTEAv1LNmiKXf7BFt1tWRET+qkN6CatIsOWFCy80wXkckYYtoQiGkob82ZAEAMRVI5x/2
kY+yxy1kXWvvse828dXjp2QttPESC+6iz52F1h2VDfI/8xBnSttgWM3fvclbtVuaoSIX7MBRzOzm
TOedBYXeSxLU9Ll7kd0cVPhGlmSYF7XHufQ4eHkiXM0Ntyz2TT8Fxppju1du4LxWzOIQmF3IwKJd
mGMYBRbjrFl3aYv+38bgZ6gyHt49+j4QfN23Sb7H2NevRlZ+DKR9AhMAB1FwlSc5/xgD8l84aV/x
C3rA2SyU8tX+rGLa4yhXX+MaFVBB5Q7pYMaXs2xCwBsakB3OPF34RH/cru4AiWkT3+VU2oY0e0kB
ArGuyovTgCRcgCRYXCscgjofv8IKFVEU+xCc2dfvmMWiiAvJRikMvNmgT+F9wWV/ne1r//C/Pz8D
rbOujf2yCmHqoLcgt9LR0JC9XR0C2UgBqkQwtA7vqkt2VBpgl+o9atnm9RqBt8XIuNgbyBIaWYkJ
YXEIRZCuEFHuWjsguAyLm0ICddhmfgOL0Gba9dwQv8GF1dmUjEyQsdK0piFqJ6JCcW7ezpkqzLIK
qn99Nct00BR4DVPJFIdz66dpf7aZUy3JgH53uz65m/TYLzRHWNN4rQw5eSaMgRlmojZCvTpTStKa
09lxFZ1Syis3l8GtIy1UKO6zzLR7iY6vEULQoaxR93cWfTHFrz1ZITPln8z9ZFSI+c8kmz88CrTA
JQN9L3RkHOIPaRoZdn/32fDIcjZuuwpzC9dU6P4PZMRHExRMXK9LKb3aflykavY82MAZ24E6ZnPf
TaKVXN4Ht86qwTQUI1pUp/L5kgk8wOW/bw1JM9YpSxbFvQ90NA+j9OTsh5Iz5CYVnYBpEHy9ixkD
t6Vl+ORWGtvH51Jymn0o0DdnqWisIfHfUBClB0lEd4+ao9hVGK5jgcsifr4DDilMVUPSlOpv+9II
OLObeMgmFGXLSRZszJyx4m78OUSfI/73ZecN+Ksxw5qjMPGii80iVIqmknBLw7nDcQIhLSDrs96K
H7QBSNSb0GweuXTDElZ6z3RRtexKe4HyUVTiWfBqZtIeSfZ55J8hPkwel4cMrPK8NkjGjujveZ/h
IGFfdX1qvUEV9111ZqYaVZdWKQbEhUh5/BchysoSzECkes5/Eejs/K3MJJ75ElDi9DUQny6LWs/7
ANe0+/4Zt96qJz35a5ukEDsdilLt4q2cEBwMGbD+Q+vvFvRgQUBs/iva+LmslQUnuDxYbY/sYSpV
gdtZohdYb33MlEb5VLJzC9bNUNa+kE1shPYzzFo8Ybg0K8MDvCSSnjLXG7ucdtidX6HSsF3UoYUZ
617/UzyiCEliTFHBZqR2FiYEcpHQM10rKHZr53emiGsoEMm0B3JiQSpMe44b4pRiadLsRizaUXOr
/y5qlbvgu6Qesksj7XDvhiUzSbHIsJ8nSc15Z2N1xWWuN8aqeQBP3137FWtSrFXEaOV7Z5rr7R49
1Ni/E+O7lE+t8zG2pH4HSS1UuETEljfnsBTradrPgPk9ou8sVyGmolGGQZsKhC4UXWWumodEAXTQ
he7GM3Xg+uYHQLZcBE6exaIntFze/mqRqP2MPkwZGt+PhYWKmWM3seRR/BQQaLCxH8nuBScmlOUS
okprKwpqRWjZ1dyzxOah+C7/eo+eIRl4gAdTC7bYeawBLRl5OpOFlLecHIBH4ACQNOw3zL6+XC3h
8AK1NNzmPyWjPTca9sSFz+VglgM3rl31xVo/V18TLcgQrA5owc+BnhhyP22Z9QmcUamg1tSx3oHU
l9RIYqg3UbZdxWvvs+C6lMBiwlSSjpkBaY5ES9tEanBui7FaT7rwkr0AHhDrThwuRcT8kuaCvFGa
X8P1DeS1EYJI85lq2ghYsl9oeiaN2YJoLKwFIw+cMk7pEuUr5c/rCF6ti/pzJrRDyut5vNj1pxkO
fighhzUt5jVDgC27YUUvahKalmMgaRhyPZwAyCMQg2TkGkE6Esh7VjXmYydeTYYdjHXP6dVeApm8
Ay0RDdUFTDqO2Kb7FTI2K9Fm04DvOhJEzq1R2MXFJc0JUWpfZ/JCNt+v7PfVa/mNb87JS2biA0Hw
IGs4QbA4k+ZQl8da0nO2XRtueh09UvUmswoSIfiuy9mcElURRnzwpjolsUUkbiZHrI6TLe9/JaDC
2n+uC+oTuK1S3GtvFbmMlITE8sydVdbuy8iyyzcXAyzT8dJz6AYyNhOyoLgA+9zcIfLT4OLkNpt3
54XBwXEwu7LlQ5KZ4OtCDj60PTkDt0sIa+XK/xoGTEdooSN5lHGAc6xZMP0Za918j75Ro0bNFU+h
5CiMOnl7/r+tK8SwWp2HQYDM+Ho3WPnFdMFoy/m6hZbxS/qNu6MZfwgs2VaOOv88cWkIUZuKmG7Y
avMb7DuldAG117rjDas03cG7zI33cZbOznsn/SwhVv4/mzqt/9f2sDmRt35ng2CDrklKZzlmCJE4
r+bGAZNKKZnygSPeuTGmI2R/4rfhDfm6BgYuZQi5Gqa2bH1wN7bmZbaWgJu0HMaiv+Cb2ksdpmoh
3x60gggbWnDmGSVW9+3eTy5mfykIKPykZdWmQWOL/vVTCt8CBQxyeqO+ROUFveHEGc+pthHx6itX
DNCcYIW3ziFgMls1tbPyC0skb/CT3rvGITsuvrZ+UpWy5rluP5GyNrqz/WDryluvl4BL1gpmuiwM
9e/TA1LvfViMF+UOYbz+0JVaxLqZUvuN6HXCJJGKYU4+sUfv9v2Mfd9T0Fyrm7OaK/tHceSbeoFv
Gk05syj0em14DpCKoDmTbB9Cik/j4LsgWysEQ0vmNwmCCZnBDBMvxr5ZXJQQn4W51RGDsWHU8Fo4
ik7kpIEhIIUYA1R4fkoR/h/a8mxbIuPFuM4I61Wu+XwBpP1RyTj5rEwPy2NSREzBLCgB8oNxIC+h
qewM2F0YBki4+SQVofPRZzYRQw919jTQ4kIOkX/jxo+skYwn0j1mKXegrdLoATYTIV/58qgqXccU
5eio3UyWc0FP82T1xlw9pdiNFCtQt9422e/CG/BJ7NBIlSiaVMgG1rBf8mcu8jvbjoDxRMZVjs7x
Q/rco2fIX2Jvo4jYFDOdhzI1HNb78xeZNfLuKbisyNcO54u1wMZVk2yV5yJf1u00Zjjy0cu0wSSr
89BF7hJjezMjii23/FCMd7j8+gI4vGtizAxsj8vQQ6cp27RPiAe0Oj7NhnMO3IAtkjH41sdblhy2
rvNw43V+PvVIhcrPGi4mjyoAlB3sEHfonAAw7BivDod3vn52y7/UhF8VWhRec7HXVo0aPSSuSKmU
yRBtLUY6bWmwRmG7L1RTSgIC2V5guoe6tDnDPPTkPOsFebyJjJ9jXqOo5LDDc/P58H4UGTLCn4Mq
KfYlm5kiF7ezVbyW6USLt2Q5shVjM3mYQvxesL3Q2taLTHCmm/DmPkXjKR+QIksMF3gF+SrdqBGp
xme9WWSi8McY72lP8X14T6tj/NTSDeMjs0yluQSJxPuZVGItOjT8EKjdvVTc4nOFxOYISC4zBoUf
WUkbbalD+aWHt9ZrCMAo+bjJBqZ0w3BbjnrYbX8T9dhNwfOnRq/MSRZz/FphxPibQPTnLLRPoLea
EB1YiEIA572iBTRc2pMl8NyYKUnNPPAaqKDgi6eNWvX2oTQEJktmxDRPPpcBz3eEK/rjQVAcDX+3
mGcU1WPCyW6HpndzwHQAlymZse9CH3Dataq32CXvaBa9N/UxPQVa13s6i9f4rXf+zf2GlArAkh05
UTULdO3eHXkOXdojNfHmvZ7q4gex73HBeHiZ6xyZRDAY68NL82vrw9sSmoP+92NHLcaND1WHe9sQ
bvP1GzDjWFRJwWbp+YGxHTa9x1DnXnuOs0V3UDOzWhcY7lGhjNcIc65NJgGYwr4hQatj/6NT8M/L
pagHQWI3vsf9UnnIcwTcMjolc5+B4q369kauGxFox3fn6SCy36lGAU9GE7X9MDCpgP34hgiZLQiw
1dGzXJ0j0Rbcaz0AtRjyFqpAhySpQhKY+seUtTVf+GYSmYcLf0YxEUKq/RGko9PwwbrcFVElHDkT
djIaBoT6vcvnWXVhG6UimfgmTJAX+cJIEi6hdZLSSnio/BleFlBG/jCkchbivKgXW6OMmf6p9gA3
hnD0iWVTtTAHP7TpTgukfhMO0cW2ASeLdQC4ukdjyaS1lXfgpWushuSdQ9N6ZlvahRC6VIPlC/L8
nt2TWyI4CSTz14rfFVtEGdhNOEpn0lsJxEX37ZI2QBBskVI3ALUvZ2cH0s9PH9ZgixWG/w35lgMk
7OdpGPCp47LF/wwm24j2Fsd0DI118n5iv0wrcKarKQv6M1Fmcyb6DnHmz2sG2U7D9Q9atigIPDW1
JgClV78+QehEGEDuu9IsRG9yPzd3DQOsZHbjasio7yiKulUZUI8V5uLlXlSa98ZSB3Ud4PlrneDU
YH544bIdJD4XS2ULfveQRaL2MIdBIfWPoT9ykyJdOFRNpQ+HXTNlLm67JWs708mJkvR8gKS9Sj4n
knQWBf4XUv+d6T6RyPOqr5kX7keIYv4NBREDCZYONiOF3XbLpN0xr4tuf5mruAynQwWD7/2UN1V3
N4UzIq0fHEqzGHCCr1ItCevTOszHcTbuLiQ50QwUrsKu4c+1/FazkuYh0uEnwV9B9hXCg7qPaNgm
lVJmbLpxEg7m/4SrkoMqHIZTO6577MCIDEe3gWg+lMLp76I9NAz+U91nwsCNlZiFoMmvoWDqLACN
c7e0UF7SoEBL2ZWXowxiksCx/YLgsLo2MEc1Mf+4/XfUCsIPH3Be3tK6a0QdKkcPGSwOq4XmHGDd
oP/Ybh1bqQBPxjAMIyLlFU4xV55GpbM1Gvdgke4UH1evsaiC6dQ36mmdHOQMIBxriYbxOIraVRXg
F4TJECeY+5pM/T05efKeMP/jNbeoK+QCAIxd5R4CzizmxD5d9AbkaJxjg3rLbdmp0DcEce/aXtM8
pkCQY0fD10VcBfZPxqgsRkvk23p8IVK8zQS/qpmc8buP+IzQuIKkMZ7ivW0stFG8Wu+kdD2uquik
olyWl+rwTUHuuiB7ZtJ3jQ+SI1cTcuZ5QKBFPifDDG9svnobwAn4hG40Pp6VuPdiZ37b18Yk9IZP
BqRKGzuLN0sL4cANWqxlUjsXCfob/WpjxFnrYRZqDtl7coo9rsIkDqpTJxGNsbP52mJFPX5c3cDD
ftd34B0hGKqJDyS6Mg0nBmsdQpasA9+y0o/QJqc72RlXSRuytrvrdcEJqG5ysRHPTZ38bcCskaaD
H4E6atSRcteYbnkOhP0owAB+JMK/Jo2TL+fJxP2JxeSrvlFJsCoiqc0wsvuR2DwXbwv2A1XlZWwo
gQ0Pv+eL2hKxIrOCjbIv++HytYjKGn+tmTOhhJN5Qw7Yk72/Y/FNMInV5FWyoyKtsDwHUUADrHFM
ml9shjo3c0HbTCwYKhgZJL6fWhGrL7GNRVECbk1TaLMfeX+3zM0zlFfGFXNW8nPEZG+Cgm+KRISr
d/FMHRa69VGWusU/kZpwY+kY4y0I5H2BRLXfHAk+vWXOtt6klp3EB6z713jJ/F4XDZiUfRVe3p+c
ujFe98UNFXce+LqqdBQ05gTiMIWrx0JELKCGIC21cTrZiiCt8oh25pR/zYa+jSCmbHzFOFDQcE3z
vkeXQ1sPISIt8kZCPoCtEHe/y/rye5RMRTwznjpLk5UZ5klN5+BWdwnDGCj+bd0/2esDzCKKTGXU
iEQRW+stN7oGiyLGZImV9eL28b6osV/fzvRZypfoVeXyLLl6YREldFNwJU4cynsoY/Hj2sEUfJ3H
nmyZNde+w8VAuC/ZsJIlORGOb/GY2UZlR0zrLtM9ezLEZPGHYMdgzM2XI4Q501t4+4PVidZohgyx
vRzRnCNvmZZ8wK3XWVjFrMEdn/RBuwkllOokDUnDieIDSPnQtA319y8L5C4Hyn81Gk1iZIkCEb9I
Z08pZ1hCGPwLyBy8M5hdr/E6Fomflwc6a9MD8K4A8p6MR0RkUZ0Y+MTgXNe7Vg/kD6jo60U75CLl
Jcsv4i29L5dnr77us+flTPfFKFDEnuBr1rWktZL1evljLhYOVS91TGk4vd1arQFM30AHKePoQJyA
XpygB6hXX3J7DAE6p7XIGvhWpQADSxwnquCAdBdg4snCYimjvOw9SA9gq7gPkw27lKMrZABW1LjN
xBDTuBK/U48vldO24TjCyV6eQVVM4jc9NwEtW/hzht1gjkn2h0KvD3s82avR/v7Hwdeg8gDq+lgv
HXwPCVHfTdjIChfcn2yBejofiWIS+g3yeuqJNtsSapICG/NEaDeEl6DjZA8SA0osvei+wP2Mdycf
Y/8bGpU6P2OtYctuwiZYAtk2lFWnrIz8Rpi9aX2FC45VKxW7q5udl1e8QFf0i9V+whLlBYEhMaxF
gTt9AD1K0NoeFfO+onpqJq3JRZo/fjnszm+AT8eBeU34Kqfo7NKepgKIGahqLe/igu/xrkNompy3
h5qz/00VrASCHt/lylIfbpxMtruc1EuIKj15b2oOZWPwuOo6cQY1GRhq68l+4hH0uED4PVy6I0H6
Uxn4MZw/+QV7Nbx235N0dQ3aTLCCLG2IwTUn8/enLGhjUHTKOcuvb+ZgJnxaZSlofZz0T5vHlwJD
51Teh7SxqbqD+Y4fjVqP69wAbPeHCsyaYmOIQgJgLAGrhfqn5juyjeaFaHBqyAoa9qYu3KvANFAi
NezsMmbxXkJBaHeyNs+Sh8l6bDZrUq4w2ucKcwn/yENzLf8nv5leWD8AK1WCPKQDmZT8alHRtsNX
+LGAG7I2g/NAl5QrnkCf0x6l3WFydmw07r5fUMFSZ50ES4xhC2LKBg/tXfo7LkA5JZlv8IKtYnd9
ksewVTbNoEZABv+0QqEe4a+Kv0Pw8qR4gpTZrPK39W4QBZV5ZG3VbmNkLyQcJHjFinH62UbjlQew
DGUHRHJDo8LmJENa2gMjbfLrMsCpHJx1P414dSgsuiIBI+ss72VvtObGqQfDWzhNh6gRXGkXUToK
LDwXBwsX3ZmJO/XHWbtW9oog/PqNwjkvzVdyllRknwnjLItbE76wLRrMjry1my1qXsHlFlB5v0NW
8lSet9zP2SammfKNzO84QeTtn20aYdSwgcDdlGPZq+afr7yBgJTRizYCvemvRCPRtHvRkvrw75r1
BYYCaNTd01tXsmwHoxa6zjGs9yIwbxebfT6pecA379dJifIP9GP2LltOD5X2Qw4ok1qlLuMBSA0b
yax7JBvxNrNxxN7NRQCdVTRIaXyXoRSytLel+ZRIRTbaVCYY59+daoX5MtqL9PDXDbj0jtrrSpgv
LQxggpqkz5qR4epKF9ExlKlBesxJbIzZzD5IE8VZAryujXv1muE8NB4KTrpnSNmg0YHsh2ey+Vkx
e5mriuAmrAYsfKwzX7BDujNYcWEpsf+o6eACMIKPSylOIAWzqkY/clb9yCdoz5Hy1k1OJFmGcNP3
j+kZibRuSdPx71wilKsiwxXgvI/MeOF9JTn8tFN7qgl0FTYRFxW8V+g6u0KyZJwDSyB2wywNxQev
7UG61uJEz3YbkNH7GF5Wi8kaFqdkJpDSyyd+1I9VERxGHGbY8eg2W4cn83tGIH0HMaayQZwJTFaR
H1tczysq5QjNRxkKKGFJperfaGQwLPevDJCqIxJ6mzC/ylE8RGOBdt2DGu8VkS5H1LOZYi7whZbo
J0Yh5GlSEXLEl1UiEId0DGzgf5Ll4JzHgrAy8Ps0biKwlLKV8npGj/B7OL63ju42KTShR+qL1T/t
ct6kwmVOrxZrfV8y/iNUh539MQYuLkT9koRyLFqwkTsn5gzsdWVzJjrjaB/1UxDb8K29p0XLrlxo
b0Qp8hL4bcXkjv6iarRNrZQShN1ADEw0Cgeecl5JGZBXAruuB4016+ZLE3zHPzQyV1qY2cEgs9VE
g5+TrbIUpHWM/hkPPY+6KpwBUUKxor3isMiEDGx0lsMKbZlQEjRGtbIIBG0sd2Wlx2SVHm0Ilusi
HwrLuDR3qZ2pEJ/NtxvhgsenyPqpfGaRMDDiMazRsIuQl8r/F8iBQf5L8JUz/TZm9xXI884BHbfh
COeDisMJVO67jkQ35yy0K4BEWJLJ4Rtvs6ehTbsf4/z9GArw0jKwqwB3kj1mbLY4MBN3y36Wcv/C
ubG+bOYPu7TjUlye/RSOKYcYIKhQnnBD0NsV8qdUWZAycvJ8ilF2/Ilq+CgdoujG7oxt9INvqcog
cwMi4z+aIy13ke/lGVFql16WZjAGC6G+ne/IxC1jcqfuQsb5VHrI3910HblSRze8JUGZzOoQjjjZ
VtVepxM6nigtnjdKXLyjwplg8HskftBWxAx1CENLUKgwGvOdVYIOtUBmf0bBcjxNTWOrjkWz03Ml
jByfkcGHpzSJIlkdUTpz/agSqjGdUF0csKUpH/qgozXcbJwfVlhfQaAUpZDIVC9d9Qsbj6ftlp/p
wQdVPPtaA7Kef3zyXw2VcsndRy4L6zrXoh1rGZG76GUZY2fiMaOYXwJhmL8aNUaRgdmJp/qyCBbn
OJf5ik9AoQmbH5nYevRh6lLmqB5QlOjdZiK26IrY15FvQA/5h7wZsdZLb9n4MQi5mrIDP15VnwMM
O7xZ7iN8wWVcukIieVe+Xwx+hJHHCgmSKGqalaO9Hi64+JkF9GLCQwLHb1h8ZLZ+NRLDcrKpp369
Q702zQ1SD9g7XtF6Iu+DoGdyZRJDQOusFAlShO5cWfs42giP8cW53KlunC9SsPb+oaDYPS2yJ3kt
0ZEHnXlcemSgt/pKKFkqVAOtEFj4iLNoSlJoSZfGsYcIJjXATI4lUC1U1cF0Xlwc7DdvRNQo9ETN
Mf/qmw2ReFNXqEMqDE1h10MJIIY6k6/IpN1bX3oKo8ZgsvcIZ/r4f5Ob1RGTSwzCuZrNLdw4siY3
ape8+HgqxJU609NIqfLXmLJpCM4pAYyex54i/1nbGfVSrlZa5jTfuaauOjxcJR6sojb0NvSV8ktY
oGzu2SMPMglON4Da2bWfIyCzJVj5iKnextY3qOTjcOdmGtdjqa1tSdQetTTL7f3CuoTS5UpnOrpe
JvAbto9xWmg6/BDWyyDGimJaY6JSn5MKvdXtKRA8hlQCpP7f4JeYtKGBvpRmtD7aAdal7Ph3QH5E
/D9Kh/4n4Z2vXZevdlvPD7kNIOedpW9AHHUJIciYovLl338HsslxX79cqP4BaTgQBgOWJf5BK9oJ
Ve77df0LjjrNFJjxbGy2mwknZDh30r13X/Y7dqqhoXXtHxLiaQWF+rsjjh7YKrBVxEweP8QbfmLl
sgX+hI++tZqOKzMK0MtExgbqGvdHh6/J+3NbhoPj9Y26ZuMSqrDRpz6Z/d59RuYgzih8w8AEllKB
RLV15jkTltiwUDeFVcn9IDK70dpYhb5K4G2lqJDA9BVwf4VvHUdsVfaONE0v9+fTZ9g0c88QJPbL
8DG2bSTD2rTuf+GxynRLiCEjw9ZTd2HA8jRYVPhcLhq3m/76W5m6mLHw7Yc47Kf6Pe+XUfMjXTG5
t1zeKBF3zR2hkcIZR/yNNN1vCnWrXpLxUtHUaA/AGKeQtun1g6s+QnFoP/BMvgH+v/t2rdUYUAQD
753v3dgUcNKTBvdRw4GuAVXVpzcx14Tx0jxv18Udw0y2oxqe97QhEjIYu4LYOSN/06dAoKSUKPKp
Uxnl8v9JD2kXe3fDQb64TFDWb85PID2fvnBIxeoN8ekLDEAizKto3HCmmUugeZsz93TZB5Pgt/8U
+tLEndywVszBHPKE2JNMBMtILplVXUqjOQX+stggEgdJWKuzaMSf13xQSp3Uld7Z1FWJqsC2EAyr
K0khe46r0QT3u5Yu4YXJu9xLWWYrnAjMe3bvxPszjStLIzq213CuNj+20hoA74pKJ02CQ2yKgptD
zCEELMxHFaRxtM+vTONALBHXa8xMyD2f8b4+BHniy9twCSUFcJ6jfiB4aiXF6oipttOF/Lo45kzL
YTz3mPZkDHZGpqwvwsdEtgrR7yIzQYdo+9g36r/qZRt+SQGbIcYstPtYpHQsMxvVIu9WLXPKsqMe
DPzU97YWlIRVsUhT11R3wELmWAmBN1UXSSMdYF6ypqHWbYsHT0wcMiXGP/8RrznboJSVjDwjtZe9
doP4RXdvCa70QuuPX2DRqZRFa+j8t+Try5+qv47TJbI1grfvDRCjOKV6Brk8eEsZKULTa3lyLYoy
Q3nyJmpnKh+to4TvQCTvT18J+iVVJLLyXAkDggTJKuJKksHX2UcrFWXqPFSFho+kNz535JDI15//
dbCYFsvwS3+ql8z+0i+uP+mN+8De0aabQig5orEhHfEtlmIzXZ4rSM949ojC5GDUR3YHqXUl4yQS
FWHhBIRwMe9pYpGD9UWcxv+G4i2FZsAnJmPEv7/tOI/EM4OK31DXsU1fhFr2L8jlmJ0j9GATmbg1
YsF124V2xRvxikgwmb/zBPkgyoMIbniItkcjHxpHfwZxT2b8jHCzpj6MKkQBCPkom0MhxW9vQ0tz
mkKTd+ey+1r1FnBxXIwUcEVlbu8+AovgseGBHMrZ2d8/XVnsAYSyBtF/H/IcUbRltUrkTxHl1PJ0
zJoKBF5OsSulz2JwSFuP/9/QCbb0TyaNKH8ZYmKF28+0ODi0PLv4v1HoZkkyZRO1j2mXmvYltLU9
xPfmXKXRD8SugpIZ5oGlCHU10XxfuERBBrVxA2BArBUi0LzcmLQnXuRw7acyAtUB1tdDIHQZRqsY
KZZrO4Kv+catGwjthLcqQ88BNflcm0vcftw5Uah/QvJt56OAD0y5+zFSmX37QZHhJSyu1nmmU7+M
6l+K3RshXMtPnVZKNd5M6XOZUZehZikGcgl6WVfeNh9h6AVHjUt9OEggJ/3f59gCnNHtL3MuBfNm
DPyLNbh5vCTdaGNhDxZrZsSfl69i64ewcIhtokPoSh87Hv1JnyncctcWMB4R16lO82F6Y/kWq6Jq
XbxcLp7AYKLeVurrnHuTNe4Xx35WQ+Ok2ihmVPXtBk5fanJ98sikfjEwQqsPnXy+tiLL/wQY2Wqx
4Fe41LWrs0SC7HrlPkc92IlG93Xx9QI3bqnI3iHkHQALc5wY/DEN930C+hVjXGpDw8SgY1nbcGDv
8jt9V45g6yJ48oGWYD34eHi9EP+P5JCVjABA00/ewEYYsvVPDI49obULc5WSQzvIsNd9vrKh4fPv
kNxmPXIzOcHRInkcEtGEAf9Kd9NXOOIjMnocKP49w1197TZVeTeNJHUMYJ1qNY1E2akb6jtkilJZ
UTopNi8E87YpKtyuXTlNTFdwSq9zxoDF9n6n1smuPUKnNH3x/hbOYzSS6Chyt4TW9l34soClUoPi
I1V3bQR1zYi4C4Y3AWSIX5Il++XVWr17CnTNcWfRv8DbLXn37Kpuq533hwSAb9gTVe8M+GiAiH8T
gtzJadGovRAN7TdlJU9q2/JwUbVhLzNQEGCoSwL9TpVCQ5AiwFe4grg6CSsUzWZ8UC1joOc11fsb
SB6Eqrj4o5wvwA+rC1a+xuIIUnvXZ+/vEQnob9Lc7Os+Pq4laAinMgVDdCK9frW4fgq6c/e6vhg+
YiilbaU4xNRHLxsGB9aesGoZhOeirDzvD1GreTum23PYhAT7a9MiM3UdLPKs8SuOkLrd4394p5Vz
CrZfH2TXbNrBXlBFEk16gK5oWPdShLxSwgz1PgKjCp0RKgRZqpjuL24dVGdSu4wF3hfE4ABcQSDQ
Yl520pAuGMZxRYz6+OAA2TqSPJwkD6H217L5p8Xf3ykyTrsRdR1dXf3TvkT5cdJd8wYNWOqdZsDa
KDTleHL2MLqZ5wtK2FQdE2LMIiCIDMt12DT12tEK4EnDzJKuHSUh/SFp/ylq3kIE6/EDBJ1aAs2b
8/ZlMDkge7teW1jPIcUd7hc120lSZExgodkp3m/GdhgqZGi25+buh7rS26R2qz58y7uVcoQIXkhS
khipo1XYufmKRdsMStAhPFudlbNHdCHOYj6d3UpNUZlaLf6IXo+aRGQS0y7K4jiIIVscEGxgzbVI
BYeKA8/Yhyn0q7i8yvF6JBXefFNhNGkqYLE2n81obhtIHkg8R7tZ70MsPHA2w8Xyc72lWc8Ozl6y
ESnjobp8i2PVCE1G/j/wF8cNPA+9la7Rvvmh7bcYbIcvQ3+OcA1azVsld7L+htlKjpkcMpIbys9X
8DXwFqJts18r5ZksX13Csqzt430ue66cb09Ug3LUnTH3d58AXMYG/+9V4Ug9686NfQ692AXd2H6z
JGTVnd8oQZmM56GeqBRsTMM4LkS9c8YV8S4eoneeqG9xN11MielJV4Q3c8xeXdzZDdFn/NxV7f8g
luhBv9+ASPm/Qu2rwYyxrfFQKyJr1+54fToakBOVAimfkk6p9vAZVD5ybXkxOk0SW9yZ6WHh0LPP
RsB8/JD7zCGWZ+H050SM4xxKw8Dfq8lEDpLQE+2X+evgTKYzrQaYXT8ZETBcRe24JtHrSkPYlmmc
VXF2nedAKLhfSlDZrD0CGrUDbA6RIVpxpkYntXkBpmrpoow2A4DKrqxXTXIyBJadw/e1inidkAFa
8mUgL8XI0TmcMd174OlRxhPC03tQMPVWc8aXFIhWLPfOm7uNMB5UhVZ6XuB8Q6XkrsWByUm3dptH
6+V+3uGfX23SB1l+jB/DLW0skIoW5ju56X7MwoccmiIYWODxZFrXIp8nWuyhT1e+xQIurClQwBVw
gA7XUAmwL2UzqaPZM9S9Cst+Ksgwr3pQJf1RDsW1jznwsf9wYUjG0j2w0eZGnzUWbXqRblHIFhD3
/0wFiVrqkPK5NFqWM5B7lXHbrdRYWsmCmRs8P7N69pywB7S7NQQzkX0FCvqWZPzaxj3+k5W55WLu
QtyfQskU9YLwGuVWE9+tB40jnxFRAwRww3ZBB/S8yrRTEpg7CSUoRliDhJoDtRfEtf724lm6aOdP
5h3cHyuorj3jWxU1r45t/VPpgmAn1knBD0OTSBV6MPDOQfN1R5w2gOVzE5G1PGZYuZsP2j1TRzQn
ek502AkbAWyfjBdI2FxxDue4xvj0zTBzVrzAKm8PmtAT7gHR1UlUgc137AK7Qz9gAvHhE+U+ZLMJ
rsWDKnLjubxdKwuNu6gslAGekmrrfoOy2EVnN2h7cyBrml7qVCxRGgodXVI0YqhlJH6F8aR6MIzz
nPeBIHgLcCyoEKJOjUTncbxJk4XF6ztkBvLhXjElvWMX2XfzUVzZtyvyW5IDA2DY8Brz9HmuT43+
D7w9u2G3Liozv4FNvRLYgHL7iMlecxzawfnazZ0+rpGPt8H64b3XQSe8U8eaNyfWfQ3o4qmnPBBY
oxohO9x58viy5yhzcXx44K/PJxvlc/TAZY9KnifZvghF1l2I7aSjf1Jyc1xxXmySDZDSrcuThWe4
P6wZBuW2uVoz87rG2VugQlb35XyvptI5Xa7k+KyUAjpyu5TColfUzsGk0JCGYwu+43HXp8eIofUl
KP9PwTeInY3Ul76pXvEuMTcgyW/whqjvreLySOeCsnKS0joeywgEI+Ag0xuhGMHiioWL9S0Y1nSI
BsRgRUyuT+SyLMl2F58jrSf1fPYrzVo+VFU/CjuV+GozAuwjONw64zQN069Ibx9wkwzGQmwEgGEm
X9XNgkb4jy8blY7qmMm51eitWiV1At+UQb+7/kC3X2LOzGb9RQEbgNxnlFf2Y4QfJu5iMcct+RBy
9uVfp4kH9fjB5hAG3r4PCrFp0v/VCDTtIrGKD08A3OMPgL+Xme7gzJFAgPTNtVNbkCSZBovxSBo9
TC6uWad3LO0R7jlzI6Xmv81xf8JsqcWIjG4RSbE6JxEj2aqJS9WCAtDwV0M0SykWSJNlRk2B9hYA
ckRA4pBYw2R11J8pGPZWdJvKrUvfnKxFuy9bYOunRsYbmkJifzHwPxcyxsv7tNoMtv+mCE7ui9iq
Wozm3j/AvoqkF6vXgVHWS+1Mg3svTQW1UVEriJGS/YzTt0WAXHhB9vSFbewjlutYZXkv8+XlWTx8
1BhIjK9/MAWIKMyXbkZxKNCBV4AVeJJnS4fYGGyOMG+f3DCtpY8BmR+m+gRK3PGWFhhyHrBYZQDI
PUazqOgZUHUdwVfW/saNBLfwxpBEFH6uwOKj6FO50uOV3IOD5mwYkTdhJLA6WrR16GCqjr99SdFz
vfdEiwzrjhSsn425pdmP2dyEMX04QYs5/Y2H24xdQEYm3kMoVyj5ahOCtipFrdXhTF35yA+JHPU1
oGlgjNjkmjMdjbZJ/iRRtuUYffyssJls38HJuz+ypHRL7APkXXfDTfaH7n6sUfotbAkOG1kuCk9+
YF8+YDYROrrdqspCJFbMHXGAkmwlB4eaxo7qYTLbYm94ez93guY3ptslWKwV683OsHWDaWoNciEq
YdgJnJM+DEfYtpHT7DMXq45L/28yf6n4rYbWv65xI5slasp2Stzey5bvM7xRxI/I9Izu2IYN+TtL
vSmLCp9qWD57SCFqBndBotzi3TqZ9EXG09o0znqtgYoipUABZJTH3BcZk7Py8PnBLQNU5ZX18ah7
NCbKaGZLmzfBDMJg0cbLdTkcF3rIJbNOfwf1h1qobd9a/25OFELjoCpXcyLoOD6teICdKpZ2wOiY
6F8CzyQnVv7QY37tIWYPpWI4SlMQO9qu6uNse4KZO2OeFzs9oUMIV2RzeQPBS/vIzucxQQC2V3tJ
jPJtRGi2ecW3+9Ue8F+GvpwRsvCS1TSTymtpa1Qu1pm3Ph4+hhYFvlDi0kPHxrKkgTAi/3xC/zxx
HvhLXhGmg50MwPg6wWEosraSDcAuU0yFV8qFZV76uNAaz3SNbPEVuM17oZgzFzqbV0fWRvbKP3Wf
vHO37rYQvnI7+SXkGdvKvxA0ql8nEI7CSBrCLBv3j9vsbjq06PwPjm81ju3tHpf7kMAS3UkF31/8
caYPAqnwM9IIX/t/SJPhV+2uKxf44FO3to3tDZ/ui+oI/hLtIGTMoj9dvmBHFmahl21JA+pBdhVI
ycfOBk2s8tQeq5Fv7gT7FbWz/d0r8+QHzjELwzEQ0dhyKzr3o+oSUvO8rZUEttEGuzvT1Ml5jpNk
e0P7gek2uqGxQFN/zgSXByF7ZGOxY5rDsDI2hbZ9suzvwpeUs9MfGG+pA5zch0D8idDJBy/xAloj
O5xki0EQmMR4wBor7ailc+r443eweRUFbGVp5asY8qJl+0FVHgr/NuAylXD7HMMtOIhT1jINgk7M
k70HFAtJUoGYJj1PKPXIlvZIyfbfLhDRXYGd7bNhdzf5Z8+rAFR9UzICIaoXonuKLqSsQdPAJKbw
feX7TsUNWuTGty+sCsOT6m7e+1QKJzT5Ij6yr75ta2CAkqdJ13S28lFfl46NJNcg3jeF9rca1BWo
uksGUkSwieE7uDtf0DUh3+kEHlwO47ReqaJkSDFr46B/+eJMSNZP5xRt4NpPZ8/CISdrAuy3USL0
hQgEL2/uVBsmsHobcAm8ydcob8hgvwxnVtsJosNJqVglGt6ThNxRo0YrmyBOK75u7ZFzeXStSuXM
5YyzCvVSqiIcDXel/USUVHOHT++GAU6a+Ywg3GWPA+jM+Y7FK9TGeF/g/tjfpTSNwxzyt60kasTp
W9B9Fwr6lArkqE/CEAhJfpdBR2Hr/PlvyUp6s772Wj37MFn3ckCXJ1128q6IanmTKvHinxEQAxg8
2xf288j+wIjf8n2kSEvn3ZM3cR1g5OG19TYIyCD9QluZPGR32iZkTWIzEKOUP10/crLZceZ35BDG
8LA7gFK3ngFIQlTFXK2vn7ZbqZPYHCYcSiiweJNsKLRmXDeZwOW940ES5DoO7NLRBx1remaox+s+
p3EkmEDQJzvJzMqGrrIldO83+X6YWOWFKRZaKPynEc9qO2Q6zy62A0Usk4gEhI43glCcWiBQA/Xb
uPy3G40t0/7NetxfNhq7QgJnsd1r96x/weFmCnMhyE7m9dE5iJ4IFN+bdvHGpKz0mOcZjhli6t+p
F6m2tuYyBVZWqbue8uNW1y2IXdGTh6Y2/Y8ToF7HyXYIj3l3ymlBOxPGfWZTRVXDK2cL+TJv3YdA
FX02S2wcLez5AjM0stvb0nzTv/Ia/DXScdgiehcooJHhBgWx2HM4jV2q23NlMwMd3NgY990RmlZj
UZMUdDwNn/u8C/TE7IgnDpE4TTxtT+7bFmVXk/8gmHA4XZ6yBQ7NyuRP9STq3gJlzGXiCCqFZo21
0PJH2dtI5W92TaHaF/DSPjPhsxZOdPNSWtBV3Ugedeo/zQvLLV8NYmZR1xBwLS6liz45/IOzI5RT
U14jtYVg5th4gCt8beVYByMiJ7lhCDAo7bbIHyMJZZw8k2zHaTxqFZ7Y6IM7a6NNiJRLYmTlXSBq
ELqGuM8ziuEH474HUuLSJZjiF0CGdtywm0F5dyj4ZFRDD9tDnAocwArjdyUebqc/qlQn3eff/hjM
SH3NmDQONpnw4JTAWNqfSB6MpNe8/TKpGS4iBNk+EAgrRrm/mWGGIEhncq08dbiOdewxZZXYtk7P
u3uEWOP+UeVuy3n2DDhRO6yw+ZNmgM56nih9W9GpsKad5jXLKUzWBYmO10bnGNR2LCYnxzlGrHbB
pQdDTSVEJFOWjBEW2f7xuO9eThtfCh/F3rp3hnhZ9iTWqe/IkDikOZSudJJ7p4vA4ZoAVVZvUpXh
K1mGg/8n0jAf3z36m2cBHxODQ+xnZ2WlgqFt+xDAnGL7JraEElQZSTtiAtk4jzQHUaoqAq//2mtl
7ofG7gl8N7KJseDN+oXF1nZMf4gSQSz2zR4PEhcM0omEYdIfJAg7Zg5PCyiDOHzbeO2MKJI7FoNd
FzDSM2PzsWkl3jXktKGB+2eFXmduOOhuZU7O9iVkxLzEYVUzcJTEsEUoHBZS17ZZjAcgsQrQ4ctQ
2WM/c98PEnIX7jC3zh4b0F4qETNua85eCF6+9oNGlJI3Anao1Q2iKNdg5sofC+9trHHqiZiocrAd
3BC1vi2IziGyFxJEiS/KY3ou+m09M0t6rZ9DskqHgdnhjL2V6zr7RIAtp4ttviuVpAAqDUNTiDKL
c0woQnFMUq9vwqMB746luO82GzcPokv1IyUq7OuGd07Sx1+2edkkgT6zr36WJDyOOxKgh9T6riIi
/Zg6bvwEwyWclZXgHO3qH8ezOnnwzccRqqF/ogEKxdaCHWi4r6V2B/VLGWQ8yC85VEUORtxmtjos
iSZ/soOoBwpplkdnhPxsXffxbckBfIXv98og4DthYWydzhlm2oFC8h3mkd/3IdIuC9EEkEiCZCv3
s+HiMWSE7CkwyBLqHa4zLcrsTgoBur5Tr5IEGxDN5XiLdI8d4QDgbDpU9TXmg0PBTGYx6stlELq5
yurwmjWW5fgS7hC2zQspE7XrjlTaH1CbH+adiGesoPa8+j9k84vBiDN/ceVmYcoQzOdr2+ilfOZ0
fK1ZzW4lFJcMPzMwL4oR09CwDG1+1oHd5v1nB1PKq44UzOZVD5T2F913hNt6Jtkqs6KbsHUqEXx/
ATnQmmdi3dASVHbfq8/WkkbGWGD1M57DStmRLvAxpiKFsWlVW9p8UHe6/oQeX7SZxFRtSY7DosF5
rP35/vaxLI64QitBD0oEa/hzyIrW/3pU+iqqvnYlJNTi/DsdEZRfYqOtefa/wFGtg2L4nVvPhqoG
vYlP1GP0zPDjYqVN5Pt5pPcO/0i9+hz7UqYuSPBdAA33Rz6Gty4cEQiQ6ZhW2f4HXk1asZg9EMlv
veELZEwyauz6e4/Xle05dcaYZNZvg4doo5stkCmLhP3Y+0VPsBXZcr+hTMdg8PtpQkpFS+h2rczU
gysC7y9PQ9wBTZRwZRs71ak01HgcA5BKAmeQk7TtN5BBpnuPBxIDBcXHgyeV98JWzDC+O/3LFfg6
loq1VrXe6531LeIoORpDh0lM7Qd6ueYs2OesDWu2gBT3GmmXkEc2KnijX406SLmZpU0C/hddfliY
brvAUr3vRygPhzI4ICortwF4f/HdoI4VPQUvPDMQ9JxOrKKZuWb/LEURyEUMcS1XM5dJXcUk9WN9
uZ7JVkkM77nOi+as4zr7OFp344u3my2VPv4sl8oXn7BfUqXmfajRr16YcyxWT0GgivNbcwkSP7BI
+lzshodCynb9lFP8XCDSy9zDvBfTfFUMaJaITGMI/SqVYajwA99aoiBDrKD7sNXRFE9F8DW7FVFj
IXIgx5vUbesdCpg15Z4ZdiKCKp+ZfYzGSd9BiegluN/jQt6+ZRTR89r54dzny7COtX8MKijh0IMF
brqHyKnypRfdyodXrft0wmiN31Ik5V34hR7ne12bp2yCRWdRFytuM57q6yae4qdMgKND95gVvECT
j+eqcPaP08xbL6/47QOZ2TaAYjBARPu18sQHSiy+Mp8ShigPuwml62qmge27fhtprQpEuBq0V4ZR
qty1sxJRS+SroecT5en0MQrLfT2AIH8MeQkgs2zD5iUbDvT4Bni23epeLMChTPDa1MbQekhzuY40
x6kw9YeKTbYxs5khGivjkT0hY+jCv4O/IjH7NtU3MWryvfgM0jbCc710miO1uKfSuNbuJ9oRQ34L
hQvcifgD72tdTHrwllU9gho8NjG/6u50Ru7eT/4vqdiDID1L/uUaUMdfEzBp3ehEqpfD3r72G61K
msxgdK77KFtli/0ZY2F3j4I2d+AGvxX+iiJjDx9wsdMHVW2GxwGnmHBDXwzaWhitdzrWnouGawoq
1MzP3bHg/bjnY31nnMZYsvv/j6ZclbvpVUwS/FvyTvCjPLrQynm15stsGx9Y5V4L/YEPqYKzcZMw
EkKSsEbadg6Sx2KDHVm+1Of5gyEw0HgYbvpkcXFHTjTO69TfdxSpqjriQb6gg1l6HAI62vsHmK/v
DI4ill8lHzCBIVjuyusthxPT7Nz097W9oTbrgMzvVb3UChmWTWYdf0hDn4A1tA+yfTtsk+RSO5tJ
5cLzAFvaG8XQX41O2EojfRgHe4CfO3DNhaNR58aoZ5QrYubepnTB6h38C2jX4sNnGYQALd5nsvs7
sYXoT322ZvVbUbAQAwQb9DDxxaInOfTgzalMSp/00zxSAUJJ2ilflUxqUwFG+7CzOi6QhEZPhQEd
qpZWSDY/4VuB4xEnw6jmI3CA7MWlmhmsVspfjwuutqk+ZIun0RN4k3dHbnfxUy2EAeP/JK6y2EMF
BZci9dDZY0GgAHlI4auAobQds8El7k1ivMW5NPb4kwLwAIFDZLrtSaAkJ7K/zD1pmBVVrftR197i
njMzxpmZLGicytdfR/re9ihJ4Q6ETxQHKDe6i/NFTuI5E69niJgF4fmv8ubWdJyViiuIQFBmKHiC
Bsv8DrDWpQBPPottIFEcAnMsRVq4qIRgSa2YpAjWM4mYdaPZUXxRaJnwo+L5STKCLvGMX5vlu/HT
j4SPONdj2p5zcF/rOxyB9sT0CFrj/EGFfKOlsDrjJVDYxZb89HONi/GcGhiriMgQtqxFAYZpF2Bk
CNbP5teVRCFTA4iS2X7yuBJUEtle5XWme53NpIqO1H0IsvR8sJUeF18fcQFa6lRL2vWx8EwlmhhT
2naHxfcPtMVx10FWA2ftEQ5wOtGv9oroxnNKLRv7kaUFlj7aO+XftqxkqCp3HelOyMdFkhO+j4At
OOh/auDsW2n77l00nrqrd5QCvv05qKzImYRvJqKNmqK418IzcsolkNWh09qRAr2reyvl9FocxHnV
azCMEnA5So9r3wGz82TLATZRAlZo0udRGyCeBo67dAQ2XaC8oS9XZVBLm+UEQgFdb5/C4t1Jt79x
mDgg10b1HCioXLwsnP2KJOoEPsi2l7ZM0jdjPzEjFX+teK0A7/+5m32xb3p6bDbNQwN97DnjfgFK
OzhKLK+IAjEHxjmodNZ5xzZDtzaz/mCKivmSb5hHr42Kjny2HjoOdQdB/yKnRP91ljc8/gGjs1DO
r9MEaZLrUAb1UlPJuYjsrIv0rR29B8+4GTY/n5drZkwiKUmh5Jv7E+s7gIzQ0/dlNWotEvRj626T
h2Nrk9wK5+O3wib93q8HNcHOzszHTqFcZQrXC6LhRN/lNSxPqIN25Pox75u1QrU+yOrLupYpbv+G
wyAaf3/aFDlP4FX8eoOtoQR3qGwyK96K57DZjbW3V4KEE3LX6ejN4jV6hp7/LEuYDIR0K6LL5ou7
wSeVqECNQTZ51wUK1vUcZX9jpR4MG1wCB3U9WRGpZcYs3jEFgOl27iUkvt2hGax716/kBrsUo7tN
tqrpEeJUfNitrq8RcVM/8WySbtyp3Dp4F+HnLx2IZglCVD0chXV/LNh6D4b5axXBTUMU54S6v5j+
f4JKyggBbXsK0LL2d7sOutj+GGtpWtURxmMcO7nd0J9AQETkJ5ZF8qVXx4URdgditvIP/F5W1ClM
Lq3X4wCL5Cmhqs29ZqwR5QvnXRsSVRoK2iDTRBt9JZ5v7oyntyX5Qia9j6idSRz1qHrtJnV8GjY3
05HmXrPT5FZhPT+v7XqHIPs6Vy5imrDYcbpdDbk0o38g7Jcy2cuvdRxAoR4CdsKuqN1iV6olxAxB
fsaUe4w6WmwsFSWvC7+PA92stUm1pVF2wq2wMI/TbJXta2I35fhMiplJw0Xl5LxY1+MDTO4xV603
L2J2YyoMqN1bOjF4DbaiJvRlAlsaMl4X8HMnTFfrjXJ8qEaqWDbFpS8vkKuR7/sayYwlu39yKTq8
qLKCJI0skQS91pKO4xnxpD4tIJVKQhT8Tu8JRqzJjrt7guya982RDsEHm2r1O79IUeGwvUH6yJzV
CvInTRal2cAJvqrZWvrJG1ZjLgxgDbM9D1sVZYLX0nmkU26n55kPuz2WkWkgMov3wDZatlG8RbcV
Z5LNChaFAoHQ1/Fqjh83KDMC+7c9xbaUXImnqUSdpvN3tj9YraeY8cy0lPPAAePb+vushHGp0UFy
wHAZZrMBMAGNdptDvK5YCSCjBMvug5qGKLe729xpScv50Q7qCvJPua/tYTOcY9aJ7FjKxtRZODo/
QFRBA12UN/Gr3xaOMidj8y4LGe++cACIycA17iHKYhMBkgOGuUcOpGAaMMdWD1Eos+1+ojNXalNA
Qcm7tWqCJsBKFgICgk7gN0ZnQhAqaNi4ZHWz6kwTNJhZpdJJVg/PkequB0U6aDbvg8kQa70w9oKi
y2Fws+KidSUKElz4Req0SPhv8qjTWchwqXWskC+ySH/dwhN1+h92mEapQ5mHgwrhuksqjTC4Xf5R
L/pXJ9PS7SQ7eRPT530wAHbjRP5JHcSPNvDjAQ/BlRHElEb6Rx7azOYXofVLap1qMy4vXf60Yekt
8vAMUVPqpjRyM2zbl3SGCDT1uKy17bhEWvLRPplMj9xbX8iC5h0Eo2zjFvAyBbs4SzRqeKHR7RDB
ACPcy/ZmpebFpcXcc464nzHloCRra4AxSQz7UBrcQqmF5QlRfpdYh5DbjXhhJbouW+WsSx9/3jsC
nd8Oe3aXWCYyQ984N2PypADhidua5MdsM6IJdEjwNYRawUUuOS5d+NSpmnM1lBO9twDAjSBMhNwV
vR7bRD9qxhtyIIXx1OUM1rObx0JgO7CZI6g1F62YQlAIvGA7zUu+BaOTNaHHp5ekZiKGp8+e/cZ+
9qX5d9CU84+1DqxHD9pa9NGvLQGOiYc6BPzJhlY2JIVEEDOb59MV7AJ7js3c74clUbkEkbwbKyB1
kjMilPDL2S7v9KWOkXA/EGHCxFWSoN9z52yWj19qYx5yZBu81mSkyyNPWVvKk7pUnzGV/NRkKf8e
AWB1aRQiLgRy0rkanInhjxmbtPQjSFllgnEj3lVfXMTSAweKybyspPuJFjZQfN0KbEtDqRgZWAgH
IyNsixxqdxZDJOSFVuyLzecgdMy7ROFSfaKPLSvbsRpDZ29bfGJy4itC5OwwLQCMWAqtXlsYIF1m
dGeuYnEyof9R9nF45Ivybz3hNEG1uYf8hBiygvlJyc2TuMY6XufdsYOwZ1a6SCJwEODFWHpuhRPP
wr3ZCmdpZ48wLbgxRkTdWCtixlIyfzp6I4N1E0jGsd+Z8wwFbniPX0W6hlrZHTQ886m/djP3JICA
Tr96um17ope2nciv4kzIFmM2WjkKTsDf+rgsGqGaqDyerqGi/hsfPwheCq9nYsRgJDXamFoiIVsY
jGlGKWETYOyuuj9TG+He4X0FZuwWjKaV1DSeZOkXz0EwUefX8ZFWURnOyYpCtkRfGFp4L8B3qhZl
boIK0Jw/QroX30KloIJBr4GhjKajuT03CTLohBPs8pRAxzS2nUNXmrtmVlb4HG/r1qgbEFrW44NL
9BDqVc0aAWsrpgXi/9tI0gsLwCWX0PrsZEsanz0jKTMqstQhtdpOSt7xfYejqrcQke0lM6VYzx+Y
uoMHogT2mBJPEpxJZCOsrqgPOllNIM7apVYmfYTOtUR/FXfM5hE2Teu+Ee8O7hjYq5OZOt7y1Sjp
VD5HY0UnW0RRmmcGfKP5AEGCxjC9M6SYtSr7O05Ia5xokKCsMDNC4jsXxl/yEv4O0fYDbW4h0920
3VirEXjcYLQAE6wZUY3lLyBrsHkz28fmFoRRv6yUbxiC2ovAWHFT0WKR8f1FAEAPXGFcaJc20As1
ekt4o5J+7BQmysZkVvtWxj4gpFOXFAViDyR7eZInBBBadmH4IVBemsaWhDDEetefKI/e8XXmL4BK
uEm4kE2rjT5zthq14YUMEKZjUjHurw7JmhQna2nGj28C4I4eeqbRjnoSs4/fguOWAxcxzurba+71
0wSwPcVuU5KLPfvlGg9Qg8AHXaipFIYKZlvcB7bdwWtfAOTYFgb/XYKRAJ1acVKzXRP4Ua6awGs7
Yn9ZSMIkCwVwjjNVn9IwZxD/3ESDF/Mrzp89kFzSEuKuT1KQSwerOpixY9OMItQUxiYilJBBvLeX
KIyZseiNUUL+ipzsSJGA42dXaPqPr2JDdpci41bmPUgbrLlqKSBqqX3Ub8JthxIntYmmkuuLZ52y
VO4XSayHrhRHsaDeV91AIJaGdYardc8YXhqFRz0PNpQgePx7e1Opl8fbGcW1JES+sGvl34zix6yt
5/HuCTU4qHONm0fX6Q1QCRw5AX4o1z/nyNvcgiYU4wTt7qHcBnEN3k+PIsQt1+pDS3zWNXMjhBOg
V9XxMhliZkoTBtcWCdLCLkpjbCQOYQw+6WyisTRvMquXtr22aDDDDBJIq3li7523Fjaoht8SjlCZ
lw3C58dEhWJsaiqrGVG+J1R+I+OG+aYYehszrlICV2b6hP8YQ38mX9ZOLS8D4Ie1FE+glwDA3qlt
8gUUrTw2kbBr0qKBDfsxmqsKRrFw2g/lYj1vmC/TRDCXlmXUMUpIya0H5lGy0onJvkaB1/1EJT77
X9pIDPs4NEKamvzM1CrMgf6mjbMRbTunWseOFWOQ4GHFNnH96spSUJKwfZDfpcnWhxYS9UWECaSI
mxbWrxBupy3ZBlofA6odFZWYDTOMo3976TzRMKiCwTbk1XUL/64gex0Q4xsKq5ALUl4ffOj3TLYd
l45Q+RljJeg6PeEDHMqSIfc1s5fkYiMl0xvHFBMOFRXMQPLTzqcswrjWAz0wjhZO444NQJrTSAvM
dLoxHp1hJuCi+5BZpjT1M+0TrSLefag2nzzAPwfgu1AhIsQfVPcZBcgTVQaVZDme99yKoROuofkB
mDmdm0koyeK10p8Ip9H8bIHJZR/qKBAKPuc3pMh1ecMNjcE6CY0NKSQF2eTmxf5fjy9IbLj+0ZOY
BXmg6q1VIlMOoJsRYpIIMFVJyKlpFo9y8FLrXgv8TZ887fF3uXPZ0HO8V4GnmZ772+lZPGUCHScH
dvOTHzI9NQc7rf1+xrSzoywGcFtdY+6K1wuQuxX9UVJHaHQmBxnL4P48uoty5cOvGubL1TTjtfn/
5AHsOIxmgWgrF/XuirCZ77UbJm8sye2pxNsiNE1LsKR6p2WgHV+XiwDErn/jUqEPlMCljhXOJbgQ
V3ddKloPnaHeiBXBSWQ7fu3nnDvPtLOvZjtQuDMNJnqQIT1OzQodLQItoSMhCWhksjYp1wfGFKQO
x5ms6C1vpWjWKTg3h+HF22FR9QrMo/AImSVqwVBwjU/dvW64FSwkrmvcNYaR25U1GW9VK/23AgmI
Ljj2zbNaEXHPvVcpsvfd4B+8z9PQf5PP9gx1gAPqgEk4B+y8YwLk9cjW+tYxJX1PD3zIwRiTKxxD
7zg/nTdsqR8MsnZp1siWaLyAW82e89p+kYXfDslCiG/JYsOluKuK/WQ5KpEvLpHd9O45R0ByD3rb
IfYD6T0WJjq1xCsPNG50cMme/CNV49xYo4gbDhF2gBrL/dyPllgplrjfN58M1RUnEuCIUou3fwws
hsbcyYMpHYehFyamyg7i/ql1Ziv0C5iollJhmvFtuP+oNd38roKKn3RN0HiV3/rVsig1t23XQmd2
BC3p+0VOnzsxpTPDm8cQ5gQlomLHseKxDVi0zKwjs0yO7oqsfCPJjbEYR8S7RTBSUHWyvEzSQ8GF
ToAeUt2a4LKkgxbAKeX+7iHtT/GOLqi+9U2v4+YkABQ3hnrTJ0P0VNLrQ7dpPAhcX3eeWOHx75GN
4DHSj8TswMhJPhpLBukb2DhTRGNu4l7fuFe2WQ8zDtXb+9JbVUafm/moIMXN3L3O6QIbMQNh17qg
F56DvdIYzdeJF871cfw3s8aGqnYbLR2yVzIskJWBUlWQ3mDapx3BRT6Zwjdmp9OQ2WUGZk/z06Xx
Anhe4NAM+cYxFfhzJubKq//E+m53ccSKaa1L/MFUYHxw6NdesQWHUd1XBhumM/PyNnzey099xP+K
10YLQ3LqtKhA9OHr3QqlEQlvzke+kL0XrsF8KpLMusSHKMIE8e2zlPjbhShH5txkQI6wH0AqM1Sn
es0ky5DUKQQ2w9jLaSAceauY6AK0JLGssOSxPa8yxrQm6Pg7pmDjwUipYLp3qT1Ujjaiwivjr16k
Sx6wLnQorZZnpmSQMwlc9HCbCfc/Z9ZkA3Lv55fxTbcmLNCbeGaHUAN/S1V/iXpy0vUHxrWAkBlO
XAXA8CgR8TLBC6zh+SkNIRbz5LI1zB1AU0WQmW4FwBQPLIwidz3DvqRxTtJJDAeISVpjUTatojLu
c083o1WI6blE2Ol08j2OtIv3kWCOj+wHZdlgRqb+Ryaa5R6rrU5fx4Lv0lR/8bORvNFcWJzYjPH7
rtk7njRPIYRfK5bffn7bf7H8fZZRbAbA9gPyZSiF/U+yh95kOn8HKW8QvxO6mrX/V5ArFp0u3CXN
sPeT03SWTv9Zlt8yIhSjbIDT+UhnBnRnAKmMBU1hkFwodwVqmm37FLjIqEqVs4s1QJXxl8mt9LDZ
6ozQqNrINuWzue34oqvnlVcMEwj4fcFqLzB8ACauOaLZDsUVYkYJEmQQI+O4qPfgd5TvQUNMX4tW
Fszh6xf4//6jSXxL4mroepkibSQyAKEJAyY7chBLjDUBIMQ/DEuD6mb02ZYNnehpaVC3QhHc85Q4
YpMVa0r6QDuDJP5D+LApn27y7CdNOXenOkOB0TKo/+p+1WTsEUcw52nCfyfu4O/9hxs8w5EIoPsr
aotpIkWkxW5qfRqJKq3VFaw9jUbSoGkRQxCvb/p6qkBkq4P84bnVfx9VDXG5/dLhLRH7FfStCgdf
E4Jr5zsGKzSU8dTHXBytU+i0XTZdNqYVeJDrBERXCP3Z4VF4ue9KSZTGtaNOoqU+RQVq4vmMXMF1
TWrJlY08PkitoXNJLm0Zdin0mU4MNKRQHq3KhHecCJUf1fhANHBAvJz345WbidlzMcCIlZGzSpsE
LSG/CXri9DlePqnlAITX2Q8Lj1y58qcWwCfHJAiszoqP0z4zo0sdbc4FrpOvzb5ceTrnbNjYskkV
/bdDDRjn5yhtVEe/SOKs5071QTD7vhxRBBwkUAkUGryDxTWXgeZpHSGOmbCkNZKQxRHm4ADWFLgX
1ZmtJcFkmxdq0MyTZYffNB4tS24EOm4lJBRnokqzx1J3ca4JoQK3AdwSXn7/X1UsuaCsKE7FHv7P
+/fKs6n0GY0xPfWrR0YIw37J8jVXiOu/IkW8c8pYXX0OPOFjvau+4LG38HDILBEZkzAh8l7vG9op
AQ8JtUvxkTSstbOXrm00bBYtos17OOeQP5mZ4Wal8GJghsZysajrEsO/zGdUoTIt/c0cokseizpT
8iz+gg/hCg2WCTLFIx+WHzG32pJrl6KEkrpbVGYgzOdto6gYvL99QpdmY1tQxxn2NSz5JjaLLF9M
qBZLlca419IK2HnvEuixjpWSPTGBdBu44LE0/OOvsFBusJrSv/HOl2JFowgZnvUemmgEbCBEYrEJ
4DQ60/+2gJdHdr74VzVIRBYg6Oq8LeGtVGSfgeyYADyLwP3/+RQyWR3lZIf+KqBOIi9gkp7h7XEi
AgAfaJiUdLrogBeNGzXZikRJ0UvXsLw1c+OG9zc2bEHeTShdR7L1UJ6/Eve5SbrbnaR8tfq5NC5n
lRWXKwPr52+DPN3c1OXRJer+uOnn6qyNXYZF/S1jk8YZl7S/fOwolnzcakF4AQ3OM6pZZpLcRDzX
D14l0LEPVPK7XNXq5w7PA/9jR8GQnuzbYe50ifQ/aa2tCwW2Pf+K3XFa4YjC/gUFpyXA88i3S4Ky
0VV1NvRgXWhKaYb0LPAi6ZARi5M5cZ62I8IWVqab+udoSeLxa1QGacLlOdvoRdTXWcevX4mBg1GV
bZtve7+TugMUZ9oCB9PF33LlhgIPMgMAgdp1iOe2Mka3KdUNTQrsrX07afajdhExt3KkDTrafmc2
0czVgCqBaUKLhsB15YeRPaYUpnUbActTvyLj6EMNfMjywhlm+oF1Ymu/Z/yxUEnDzHwG93Nbjeqc
5u6Sae1nCfp8OWsctQ59Q/XIw1y3/VCMxAUNmIUwL5xWKpezHaM/ypuPH2udcPjel5VrH5V1+8Wu
WffCiriiXkjEg+2EIGnmjrd13zT3RtjEjZzGrajKpUcD/AmJ8buKsjlZ88rsbH4bcHlL9/Aa7DCP
aBp4+Go3OwasTZ35t6nr53e/KqcbpdCvtGd5EOLRQtU/8DBG5u7zqFukT1c47cGRu8N4Wp8f5OAz
0dO8PLoL8HcsVm7ajw6gMaOBHGYcWhcB49cFg88kHlJ3vBnFsWxWdIkRHyS1HQqMXkd9WkGyRNjV
/qW9Ogo5/JoatOVOI8uyueY7UJd97hh0LP+X/cHFqZiantf+NTNH8Oi22c8fitvy5WohtDoUVqaY
7KLWT/CeEx4H/heY4nqpSBC+Q2DwS83k9nd4LzJiGRLlajPUErdzNkIFtxskR/Gh+mQzPAyh7PHm
9ga75+x+iZRBW5C0Ek0ZZznggGgktbOzrPd5fZheAnkOJUEU++Nxim7NL1GI0lIoW96s5lUOj0hb
oh3YiIUCaOFOoxGxKmNRBxaaRfGBEmbOnoeEus+vs56EnMOav47fz9BSXRULBw5O4ECr9wJnZv3a
LnaaJBvfYMVtkQtfWmDDycg7ul6bpxUugtkg0lovSPNdODz4nzXhC8lcdF7YuXBREfI0siC+rFNL
BLw5m2shRVYPxMbJN84r/Izen0p1NyInPeRmNedwRNyEMPF8Ezsg9R17pgqyeve2Vad6K+Ia4Kh/
kI3EjBX0UeI5nKMJrrJCeaJFwDCciOvdOrN1X11TCKfSB6eWm/OmIutmHZkZ3/cGM7v0xnFMqlQt
CZeyfknuMLeLWu5Nus2Kj4ogHk51Ta7scwK0wRN6aejOHEpWhVv8LatNytOpsy0cBl584v+0K7Fg
iw2RIU9lCvaBghczqS8fqcsWt9YC9gOXT+gn/P23TUAZSTzkfPyF0HZb0320xb1C4FYaTV6sgDfd
6YJIxtuzru/vrFw+gMqUC1EYjySipHcGcBKGrrOGE/nlWtOeVCojMsbItrkEV0Hd4CeNXvNAYcdm
M9lGOpbu6vCKTDtrkiTPhR0Y+Jbtzm8hL+vSoIVTedAfUv225g6FdAilgh9wvzf5qaJb6CviATsO
+60/kZDOJkatxJtf/3uH63ipYyCQrWAnV2/+fyDFMg6rn2b2lY9HVab8DnaadXql6oQvjdy+dTxD
1Tgk//uSPhKZubw6F0fa13wxl8jZe99TE7r26C9ErSYyQ5s+q1MM/dEEIVzgUvoa59wO9UIg+d3u
4/LCJmnBav575dFAsE8qrW+xULWRcDCGqbxOQHwbBoTjvu0f9H9iEom9WF1bXwgtZklI3fSP52sV
AVMfOqIBi2PeNhYdY3qSattznw4qVOHw0+DRC7gMmLHLmV+C9/XiY37a//NdfD/nMoMVNrcmTzKg
xHporEk6tgjMI/vX21cDizzOU8XvDulj5rUBVT/VoDpur4emT9NKYevvHb9bz8GdOMP6M1dAyATY
hpjVERsgHwbuX+F9zITT615GKVemxIDsvxtUiG2BSxXQjpMw9MeSxprnySTdV8OCznEO+8iLkKhG
yfCyNdfFEM4YfksWQlENSQW6CSYP6HQJukjQBJIEQF6S/hhlSlL8/Fx8F9ASwpCPIsn4jptqC926
wBS9Kk1SIavPigRaGMhR+oSpEWg+CPP6Ema70f72Komzz3ZCM2COzu1GxU7NkSRJxOz3GeBTNw/N
y7trOGhnvO2zCBz1j7rFqiYyBcaZBg+V1PZpQVgNeGNXDB6qdE+K3VSdvitmqFd8lhwvqD7Oz6IY
R/MXVTTZ+UzbeWBLK3b9b+YRR/JdtOgFHpEm9LJJOMeDgsy5barz9yHntpa6LezjlO5AbAi88bpo
AWBEZ11LO9QxBS/iRcDPCB0O+bVFP0p6u3dYWRv/7V1jb05BM75dCmpFbMGJsVH/CCkh2PGhNSW+
K26IR2O1iO9iNEuDFQzv0VgoNi/uCjzt/9Z09Ro9p97s5odWrqD+35n/pJsNGwlAsg/vid2fwS2r
V/P179xNj8NZ9qc4SMH3dlGH3UEEW6sjuNNU+Uz1m5Z2zINyrhxq89z1v71qmhDMMK12N93vQ4nE
q8vWBBxSuwvJy2M6U0bc577YPNJyffpZytn6cWp7LdYYdMNdAeOIKlIERfschQTRYPKbZqgXntqS
EtWsC4oWxeDM5ZS0Xoy6aLg3VTP/xJfwImMTsze/GGK76dYg260K7BW39dKUvdcpV9rpZresVZZp
NecsT0HLxv6bkGTorcRzvowLtGu0HAg4XjbPrMlM6dzmOYOpwJMaCNW6YCEmPkrmQD8Mh2vrl8Qt
E6S3Ex6mWeK+55W5kD3/GC/soNoPVr9Qo5SZwTOPKuLPOulCKSSMEz6/WfmG1HTi135Y7yCl/ysA
kiE3EFg5fcPAIdvEXHcSMM9boF51a60CzLO9R4MlVqilcVf5SCnqEzUyRpghmlRiGDmtJLqq+HC/
HLpSzuBH1/lCfR1Lcbc+ExwGeF8bskz3VSxAZ/ZBTbZw2O8WHG4U5GYNb1LQNicYg7ETWKthXhko
RTHxYkzlWtKN7GtAgY/+zkOs1DZuHAFbp6FOfyDTWJ+18zbNZi/ApzkUzS1fA5CZy4jBp3t7QN7p
SXVqF44X2BMSkzElN/Yx+7kIgU3+YnqR6iH+p9SMWgTvcZd1xg7lqx/35SZrQZxdvG9AIv55Cw1x
YUawtgC0y66epz9CPAGgBQ/YNowXuOIZN6Zw7KkJNywoo+yuiitBabwQRpI/wZgWxuwk/DfNFgfp
9jfsPfGOedjk4GswwRujUlA1L9Go+YqHId0RKcIqDRRbFTla4F6CJ8uJVxc/JSbeuCVlsS9DteT+
twXOgbBFtOEDhjbYwxBeLoymoXYl7WADwTU/mhWL7kqRKTiWYuDqUB6a/pU41vGj/Svm4olyrmT+
nsM/X+c11G+iv+j9i7IaXLy6VWTt2Ii4cV82v8aqo4b5dBc6flCtqKe2/S/lzbMp7mN3TfY0gj6p
ucj1mEFexn1IBXgRWKjmzxBvCwomJ4FALDiv6BNiFBce7KWmWGUERzxCQqJfLULv36ll+LVkeJn7
EgeyjiK59Ivs6CcUqhqe5dfaRBaUVPReJ6MFU+xZMbhRplc6TtnfESn/yQvbofLFYHVUSHVYzas0
r6/y6UmANa9s1k/8+FMaQtHMJmjsZwpZFh5FxRll7ZquZ2Fpufewi8ZM35si90ebtD8+lnUi50Ut
0OboBUpLX2ALpf8tOojz/vIry+suqcT6O5WX75GC00qEMhgyX7ZZhv9SABqO7/qP3mI6OCebBf9h
BuIaJL2GR7urvprbGrGgb5/o/7nAlq3M6RPDcWm1ATOX7giA5MIxKeUgC8/YUCq6PChyNQoawfI3
cwITnqSq5eb43PiO0O5mHSHB96RDfIQcWs9s0GYf5M/zNywraYWE3hlhG769bRq9FjWwo0k4UIHr
YLxNHFPj0Gtpz+Tj3ZsQtHrvhLK7SdPwbct3MOSNnjeNM6xVf3MCt5Xuw11F34grPkBiKk6waWBg
WvUoViwP4q5/1wQjYQ+zt0cerAtaCL7pqD/IdIdwDeLuB2qSKhtyWnajrCra+Y3i6vC07BeicGLN
v+XCRKt9FHwxH6+7z2Xt/itriz8/50eCVURCsnMmHRppmr5QL3PwDIbZxFBslwkP/LVh6DCtFhNS
Y0d1+xL7crotIW8htogLA18WFD1PaA0IxC4h943fGCUFnFgKab8z1UpBr4bZeLujBn7FHemnzYBk
W97Dy8HWQQ8NbQgRftDA+sCZ2iOQvIoNuZSXLv4CEuzQYZvgY4ZPR/2c/CRc0K+6TgnFVuXBuoM7
8ZRn6CTpGHlLOFalqzXLxy9PhQFI4SsmUSZZlXseeY3uJ46OHr9h030KFZpvXLLmoSgDQssqlFg/
wHgFYtAjmE29WG8WvdGbw92OVmjAZgw5e6Dadujyk+uwhb2o/bAJD7gDvJkn50eqvrBotAFMtG4+
8/qeLfYL/+5bLlcty8ScFqsP7DHTLGvE/kCOhdgUT1AbUhC7qumq0m16w5LtXVW+wBci+3OzcfSm
6/66MEI20BSN9hSYKd2ip8cXzNDE6xTJ3bpK+Z+o8U2LjeF0asw4H5/nSNdlE4JUB/nSqLELR9rb
QZY4VMaUQIbAy2XfjjOP6UjnIIlFuzuce3NsyXX4yeD0hLQgy1cwoYd12eqSjbc8LU292kV2Z4Ic
2uS40YuNJP4hoxyIJEjEkGT6cW+PN/OoAEM5nfYoQbGpI4p2XJv2yBp0fIB7VC9jlMio4l7z8FTe
wToJM3JQjvjMreE50gB54Z5MeotQ6mmYddgUbicSTW9EVOCvnLdcI6qmChMyo50MLTUbgLIv6uHQ
46NkLfnFr10ebXbDBUKZbirwHCAJFrn6nfGKLrb3yaWe4CLSZZaDx/yZS/Jwx7nACyRmNiBZU9Xy
ACqC8QuGnxEMw776KQNOr9mGXH5gEq1WzsvmTlft8GRa50i44pCoJm9rOGa06aZOveubdDhDX6lX
UfF5Mq86uc297Pq4I0AEgHqR5O0Wn141mHWMCJVI9SPaePv9I0OTRW3l6fWLta0MWjLobyU3nUz1
ajIwVaMzY60LPIA/fQ0aFCsOJXISIvUPRtRo1ZeVYta7m575ivtvM8b/V4O6ZKbLNzYl04WeRNHy
VYME6V3Ag71HCZ8vvkCtesHoXGmRfTynpWWSOs2KPgSOtQmP1q5VBKO/WOTa0rieXrjUfGsUHAMl
oxTmt+S653QRYP2TV9Y9iTxejOriKuv0n16eB4SQgkVV7oGKABcqowdg/lPpdaaR1TMbXFQcIC/f
8/G1edbTF1LnXm3NeXcRk2DiTsgfv/cp/z8I8P0+3kVf4VoWJ/TzkFSRAzHzFeXlxNiDuW0O3nh5
NUh/GspAcEQ+5FgVj8/EYtSDkYXkoRrRBljDHfTvfQLU+HO35KWml6U5bBAn9sCaiKlt+X7nqjK9
Ubbq6Ggoh2W0veUBxu1aPHYaj9J4/xZDMqXzlj4uRCvIq6i79vDT1cYC7TExp5TXw7dwq49z5MLj
i427TMFNAj5MZefZSob8ATXLqBz7pFMqx/tPA2jHTewSGMz5VzsgUtlwcCnoHuxUEqcN1BEe4ysE
e7OHoSBFs7M9vcLpZr4FVSQR5Il6dOuChy8KjeLxvfMqqPScOt2wGpRW84dea71F6LWNgasJVLl8
tlrVG/cPVUAzzchNEqsatze/DvSSJJZU9POt+sEen+7nENOXed1nu7LS6PEF1i5YUOuEGKB3IWmq
f2BCWEZtBw/nTHC8ZIBN19+EaVaRZhChdJFtZI2k+wekf+fcUXehexOPWlLwORGyj4wu7VFZXQ8K
9yZS9xrQ8iI6xpP+zvN8+ARaekXK0irnKl3e+/z8eg4ZAzypLXAR60ocGQ11Yr5xJ8coJXaRktYG
UGFJO+/6D3b+UTllYEtrwWCMhXHMZUs7sySyhuVneodRpN4q/mZ0C9tBuLOfqfLoY4Qxf7kDJaR/
kcqvsLDRqFg+L/qMiS0/dgWwgnBFrIbGxJ3uLV0NbQbCHlHUKOUE5uDQG1w5QX/vJ+0k7MbewtPu
hOZsRhjlLIkCMQQ/Tr8j9nqtG8QK8bVQ5DRHsrezlCwAl9SGojVe8aekjl+dwlsods4eweWN4gCx
iJTSJL+vlq32aRQtKTNSd4Vj1bmD88aqvBcN+bhHdmZevC/ceMFeDQO3V0ftLSUaAJxrjASdY7jw
BjkJm/fgQooxLZoEvjWOXTiZSNRncivz8JpikChO9I7RN5iSC4xStQfdo5COnZzgRZf+v0tQ7ACf
Z/Csc1z+hZS88zxSrIVNhHCQCO3ZnAen0lKc38mAs0ZWMtwTcv0l2qP23oKV9NbXE333OfuMmaPI
VJ2bbShkUl6e3jvbo0erbO/kyNCYIY0zPAxM1cb9yBS/oOJoGfxCPZm/kg1w22AoYMHgKyPsHPsb
GvIC9zle6Fa4Pz3QcO0BNnkhi1UtprCl2VivjF24Lag/T9+yl1mV1Md/gFpHc8P4vJaLMPEjpoko
pAYrAPaZUwfjKcleYYePqCsJL7i51/jDZsNsVjzxn6P/WUIXlgA82FpfF9IlcX1Eqe7eU6CkngHA
hGcPC7U5uWWOz//zQwLpV3p73Y4Zmau+w9srMvOy2c5cPUKRxE+GDFEE2/v5xPGgcCTz1uSSBW1o
ykw5OD3B+W88DXI9hVteWhc91a4DVmE4TdimntZSIsg8+BFtrLJ8r76xzwOCTFqwmOpNHmlQ2TUD
Ph1Lph3D2QGaS8ZO2fi11F/jRwEnzH7/szVcbgmvdO/dW8yWekDxzmOFU2rjGFdak/dLwVjr69KK
JgeToEPgHew2x7l/JnEcEBkPftKXPVVeGYTdPf8vNOQY7AQu5Ro5vXjm1hw90tRAuV7gCRtqnRKy
A612wnTswIktC0Yll0mPqFmo9a9k49/x+ytAJy5n0AUSoLKfu5OHNffNkjHaR/H07SmQNMa/v0DI
FzCMnN63fROLrU3PhH1S38cBOt3PpXapZ+KuilBXk9qEyMJkRk5piP83WBbrtZyhSdQLgU36ySa1
WyiMkiGR7HS9iXvwBZfK5gD0ujbDqFLc8i2/p+C2LwRxUDXoFQxfbsbtvInJQ5D7Lpx94ezDZBg7
yHirU6S7Y1ETd5ru6Tmaet8wNTSI7a+BlSITP2gSS6GM8//tOcLhq1hkmO1f0xOj8Ji3UQku3E9y
/z0MHcBghrgY4cS0rugpspZheNPJ+hUV3WbCYonTi88jI9RvMIOhMLRf++DZmPcUS9m/Ox3qrrVZ
BDGTRMZ7RrV+RRpiwyBQrVwYvW0TajWbT/Ef0ErJMEIXnOkurOGsWXXmeRayjfD1IImABG7aCvNm
c2xPm3dWoqwP07unKdJOF9xEPQlLj8xZ9r7K/NRouEWHy2R+mlZQ44MZDhCbCoRKC5vC6NpuTFbw
quu4QHVbKX5mwjmt4+4xz0g4CdBwHn4Xy5tS9oEnkj+FOEooDvsusy83edO/cToGnY17TMrBCU+f
w/kIK1qZE/dfltv76d4m2ohtRL4TmvDpFdUIrKrocP5yEuqyEhbEO7b9sK5yItoe8Uq88nTZP8vg
b+YYCnHWZ500KDA4aBHW8QGtP9mq5p8HWpBzQGL4LrO/ENst/2OJuMm1UzKhBhdNOx42b1VMFtMV
5R8LbMGpEhPEvbdgsxfRGRC3mI4Jnn2TIPY10SOcMQdXCL9+mtWOP787yJqDYzDG857EzP7TBwNi
U2ScFtIaq+UFXxsvBxCDKfooyPFnu8tAclmFh4gHDcBJseRuD1eKoXnHOunSDtYNnv/wEhZOIlnr
GcQqFL/BJrfk5YGyFP/QX+dpHUJd3BswvH6O/UuCK/k8bLpu1U431Z7sCkBviO7/Nefs+ZMsBq1j
zn4mJ5Z9GEgppvXegpYqsR08qCkssuzE212nWgT/1KENQnUWjegdiHmWiglOxU1XFFcPtugH5jaN
SFx4nswl/XRttSuXRrcVCtdrcrR4Rs4zBWyKjgEujyMFKSKg8OVWXKPNX+UQlabACQAAy+q84wcd
eff29zTLEp/L3scBUgNUz5Gfy7Bo8YnWNOyX+LtgBSzfheRgqRQR2dYecS7kb4LrSrxn1+6Ih082
nmrDrG5wnhHHT1KSgK2IdtAA5a7NMBN6dkz0u5N3CuZKgIAyt3WDsACxJtGGbUT6A500xO91gXD6
uZskxm9vPuAJkuBOU7aigoEPYwG2NikJdWGH/HXkYxw8Z2DAJ0cxmHr0hRWskUcG3+XiUHosOI1u
2cRBoBHvTNv208gh6Xfl6k2nXnmp9JX52vW1t05qkR2MFZLTnXMFYx6M6/UKx/Acm0fUNQxuEmbb
6d68jW6t+5/e6kPtryu/r7RZcNedhJOY/kS567BZKO1yQcdYaY74CxrHmYcHKERWdhLv+t1NMTH4
J17nzZ3+KjD+BBS4Wtlmf16o/U9+cWhPY2wkksrK2U8yZhKWhHMB6HUYlP1afNwWGUg12h0HN/2F
oT18pVEHj+Bq3GoGwPKHv/5yFcEmq0byGp8o9gXqMuWS0SWRPHIxA4GLOIIPPAHRsbeRX+9FHPQR
FTit47gD9VNrIcbeJfruKAcfleKaSj62crth+2vSwyUJzz23gRf5DlTHe4brm0vNH3DRL5W5vBCY
KpREQI0dgPLRs4Mhm3XeQTr6ekrTHbMtCBZLiOp0SIlTNp3CAvKlj8LSXok0XWrtxaWH3OTqui08
BF9eQ075tXkL3RgqHEIpr1oTOWdSxs3I8w/hR+wqzXpNtypa9EXv3FlVojCQJqEXWMwhznbW0Fur
L2nMiV2um1mpOQV2pape2uazujgJIpEdh41fp0XytHD5Jphb7+yh6bONCsEjfnLMW3qD1Qj3zJir
gW5peM5blzIkvGnaOZ77iCQtSSzarLxPvpTHitBDiz5R7amSmO3NQ5ZdwPKSXDlrDuMfCv3fpEep
4Yt85cIK7vquapZo/TjU/C4ZiKQQGU/6o8nKZ7BBr+GwuMKUTWpGlMRPxL/D4PLnrg7f3dJoGpg5
duUv4iwfDL7JtY6PyAkIFpS9nWXGopFoD7LW3HwQ5VU9t2KJt2upSYUIXG3SI+Q2icx3PMaj4YQ0
LQJE3GZVnRRzlSMGZVf7gtDs4Ytv4weje8dkIgWRIct2nvLQqj7fhF5wcU41WcxaVl33Wz/pSoui
yirAOnDNuxZE/0NxOwcDftA1gQMdx9uIbivzeHryF4CTjQ6LejXV4Jd0SM0PdmdyM00/FxfLpWAQ
1UnUb0J+YOMJm0xlSTUnUrUZk/Ty9pf6L2kpt0FuIcDw2hvUQ+GB5Gck7UMFap0LvaqfzSXV0E17
1QRfEECMRd1XMLZDcIUT9Z+VyGIcu9AUk0AdS+EUmklT3pJnc1pOysDzcNitJMHv1F+GS0C72erm
C8Py5ou+Gr7FZFo9dPctxad70XdJsoibpD2o1tb8cDzcP+IF7gwK9HOBKE7ZjHfEnPzoSWkPrQ2Z
BxPLC0N/jDg9PG/++fCQEbLecZ9G5ZDDHRzJnCbSI3ic/00vHkEp3FE6KLA2kaQ/yA5GYAgbFpx1
CUdCyPwpxcCDmv/cLXb6yX4hOEBFUwH5L93wN0/3625R3Ia2wOQuHecVXQNeSCQZOTVfy5qXXPcO
DqS0lGlpo5LcYRfj4fCpwo+VLGzAYhxMviYa/LgV2H6SO8VcTzQhWLgRT35KOQjHgRe3TJu0k/xb
qSrPDV2hnQfnMb0wED6uscIzFJL5g9aox97xqg+1Tlc8vp4bWfFX1q604XLmxWXTcSHLTvoViNwt
akcBH85RUJ+3oT13fc0tuPFnJw1578d0plrXUcx1TjC2seigCsWk5El2Vcd7D+bdYoJ55eQRsVnj
Gk+yw0k2KXr7wG5t1ZT8ngmkvrVOSnA3TgxP9CGEWLN0JHZoXxedOipYDd01pPYsL0XiQHD4OzrL
mKLswc7Prq4LYy+fVVIVNzT2AI79Z/QqV77ljohlCOPLELorhdWWBRvvkXQTJvelZmaxnfrycB9A
G6CnSPWXPZDam6OLONF8mawKKNb3FXqyKJqDD5b3J9RU14dKEgKy4R2699amOVPAqJcIlv2R17N1
S3J9lPrmHO4VUKVDwPyT466ae2JOvya/FXN1GrAPHQSDbL7DjST32rGuVkLGS5TE5xqX7+uiE+Bh
eHPXDtpPwanqYOR6EzmtR62jBTioudhZrmO2Xl60Lx2/A3Xog1lUGPIlxOou4JZI5jfkLpoKwkGz
KnkKNUrBWJEgeKdDP+nVmLbAhKmWQJP/tMW49lN6spMWIPS7/X9PlkfeE3gCDyZ5x3XjUdf0XZma
FmKo52NY4+s18hdWgdM/TAu0mFmZq96CcT0325CL9ZZi7vR935JSLFCa1SFQe0G2S5OpcTn0Ceb5
o5Tekk4fYzjnEPWJ6aES+hiRQM2cdfMxreNOzbR2GFTOFlRu8QEcGRHKcoouKv6Qvgn3O7/c+Vg6
Kue65W7QjGzA+dFEzdHZXqlhZeX+qqMeIxLbnotkT1sm4tQKuUQnF92IyYKDuuGp/QTeh4MAoE0z
rCk08PSRL8Xilc9sYm9EsgV281e1gmbavZGEtAs2PhwW1cFBimPNl7y4dMvSf0Sr9lP656iwTqYL
W3HWIbvTJTaw+dHB4Xb6Wr/pYquexlrl93xvViuOGgjIo0DQC4iPXmVAjcflcVh82NgqK7KWrYbw
e6xXUhVvhBInik5HEV3pkiqN4nSaBV9QHYnhYuppINvsTi7+wxsQHFEQLQevWV/G5vB3Z6h4nIJ4
V2Cnu+ddt/wujTHlj2wzxVU4ZwSonKopCLXsDAUeMZGgLZnByajkHfQXEkwRiXIt5pkLvaHW5VsU
cpFrfD8ZlxsQKrlvvoZCncO5EpDbeElmOTukBY+qaXQJBXb8yib7YZY1F54aboNjw8RMT3LMStcK
Hx/tDzYtlne8XEy7SCQyCSBopW1igXuIzq67iac3Wubf6SsHhQQ8/IJ5i0o4vzr5ANAA+PKAHawT
c+1onYUYfw2CqFoNUdG8HxZY5wvHDevFKQkJiSyI+VvRXDRw4qxHtR2CB5X1NuZdPrq96q11I38L
HerTDu1VYLQpw80BPG2BhCcNijGOkHcCAWYH7CDVsChV4oNKC7h5ToFbPd/7WF2LGoYXKLnMOByg
IxFHwfhLxjd3Z94SpIyJVc1eNke557H7PnhLFy3j9FLJa4pRUd8Q/XAbcWV8Ff2olbk1nuIiCYJO
6NzghsytSlmQoX/O99S5afAoBMBT10QbX+5PJf90XC3rnw0j8n+t5KwXEAWKLRjGbiSAlNN35SNh
cGRTNANW+I8eJa4ehJ2OvSWf4wyI7TkkwZ95MftNwfCEMRbmivhcDa4ad51s42x5JH6wKuH7RRCF
YFTXD/pSZccgey/m9e2k3L0zDMgaoUHdbIxkky/aR0RXVFIRsbtejqQPasBuvU966ON2VuOU8Hh3
cM1KKSZ+yKV1hxWeBfVZ8mo9VvIEnfzTdNt//wPPy3ezM+9/29wUScWumAATOkmtf56yAnQ79LUY
swkXAgBOojggtzvOU6aCrz3efVSIm99BlvqTCbJ6Xlshlcj0HgHi/+CfpFgmVH2mXbRriDnREXcn
6dnQ2Cby0pWSRKtByqaZyfSsM5GZIT/JXUR1XDGlPIo09A9+89PWjFpAwrZsh2XH5hLLaC/4Rx2P
IYCVJyt5BX9s0gqYbFhmsjVyz2ucTWKy1M8uox+T3TGUcYqSSRO6mI7OtB6ME6xcEdtuhVt4GKnG
IfOpILmZ2vekFjiesZaDbksbcEI0H7tqdbJvFq+cXoq9+HQ/MmDIWsezUxat78HxN3r5FMlNQEz7
jCt9xroax9XFbcvGrcFelZlfZKgv+CAGhy9Z3MxEzFFv4KrBQ7WtCBYZHgdFRTNdJwJWQAG4tpaq
dh3yRk4zMeTb48mAnXbWyY74+DWg6Yy7jSN3k61+DsheURntfP0/qEPoHio7Qm3SDr8WEM0SWn1I
spQFYqxNTAppzWeJU71HMLPjzGJY89M0YfWztshTkGTO/CFwB/BgWR+LOGDw19tseWp5fmMT697O
B8GIg4p5nzVsALBcaAevSf7Y2rc9Pa2x4DWP/xLczrZPVs867/lxiCNoeW7uMtSKXEeOoMbeZlzr
gfDGKcWdqjVKl1/paf8AHaflCqi/d1B7VCTt22zgQ5UqomOtYGgOT70T5VQ9A+eRiKrmVda2huAD
oXcOtZ+d0kCgv86+aqUA6nbN5FUtV7ilrEg4F3sagYjf3FusC7plWRMETg+1oG/nHKl+fMpLKu4Z
bMTk3JLhyCa+epDXaDqxBHqeYBSqVN2zhidzJJ1tHMTAJ5ajijyBLMvOd3lqVdr15KvvXrPkZcUf
+N9l/wH0sc7XKiIWtXsMb9vt5vVC0pYQSw2sp69UA5b8X+FTFTDFoGMbihv/85RNhrbwkNdwb2+i
6cRRN9vB4lDrqh6C8teigW0aiTA4xWIBtwhadGjqyZRvxBk+xfTwYd+2BN52r69iHk6SKhB6A2YK
47zakpZwOxjd2CQbcP6zAkLdzKJHCq9SFH0SGHFDhgMrQhfGTYdtKOYgZdcsnLla9UMMF0i/8LMb
d2DmW0T+9ErSzU7FhRS5Bb3VFOrp5GGWLRKNLe9tg3VkAS6xy9G6zNGuSiW84uAFmYfAH7rBgK7D
jMAIZZF1/ffJA/hTFLl1hQu9/3dvOmIY0Y0mqqsCamRiDqPfDVUMWb1UyhdGggxGtRLaxxcn2WBg
Uz5GxwJqRjloTYfd8t3wkn8RS+ZHPxyvkgMcvrI7mZtZ2nUXRYu7kN+0vyZkYVuIsBwVC+Mi8hxS
f73ODOwRARKEc55PXs9/WUTP0loF2nq5EK+KqomqK91C4nd4aK5lD4YnuBkjUSuqFCjDpfTtNfI+
zq9ARvqcpqUZtVIsKMIgu37wbkK0Aud95O3GDro8W4lRmaBPXtKg2mLzmV41uyUsHN6peQ3jN8JY
66TaswzeaiyCRvxgSffxazN8+/d9NpXby+XohxialVeAER0ZTz/mcScOf2KDZL2Wi9HVx1y1L2HZ
HPR+kcbZG+2gJ/gtHQTVcoVh+tpbW4RoQMGVzN9K5cfoHAPsAql0aM1taQFKmbjhOtKKSW5UMvoG
VT1cLS7pz1EFCWS7CCBkM/yE/gqscRbQ5n2mOiFM28iT4aaSHuI5wh3HsuiGpLfNfon4qTD3pFQ0
NcgX91E22O5hfVp2vgap0FggrihI5jb+CJV/BsCudUDz69qw64rKax9lGTVknE2C5ozmn6Bf4kyW
Mopg1JkKJFKpNupI7p7OLLAvYUTpaNEB9VrPJBK6BdvS/Avjsr3cdZMDEPUE960qoc2zvNRIeSks
wEv2t285DQSyG0170jLdxs6uj2+XBWld+n62psSYJciAiuYKMqW/XuJroM+nv+acnbALGVqBjKH4
rs+NylFmPL/eH8mAKZaNMTu62PiQaBR0BRLOyqfiOE9/KspPmM37Mi+XaVUbIu00Dks3JJ+nneJl
mVp9nJvM9TeZVzW8fdOJhh/cJ6/Z+vxWaFeVO9UqDl1SRdQyuV27eJzVLvi0h3ohhmtTVpBvfda/
BPtuTwszcAHzBgbCuFu6WvprcA8g9uiGcAJbZ4Iccb7CKFtOi9jlcWxC3Ua6ocJfsdRt5k3wmfpU
40FBccGUa3dQNSq3U3d37+BD1ErahjAcVR/KmxQ03oKxvU/krNgGZK7MWY/zonSFjQ/ieP06iWel
xKCZMet3aSoWX8eZLSOxxFR+KTdgwewCFqZddP/5wHetSxrkcC5Uypvemuvu183dIokIIwEy9B0g
seArGhTNd/1F5aQhZggobPIgMg38NlHgSgF02WpzS+I/CDt5PtpriOGu1rLMCOcA+vlNw1vMzY9Q
YPR/SLBazR90NqTykml23OMZzkEaxngMHPLkKCiGyVAREc7hp0tDoPjBDg0PE83OJ073/MC/vjDU
cJdY37AIBwWeZIaYlvZNiHKOLwG1yjobJ8zTjp9prYFO9nY9Hh4wyPDVXGdLFqpZclc1rK2DVjHQ
K8TpuDBJwPhiOpPb2w7/dXLTfUq65UAJYuV52pmlVvrlITVr5e1lDsMIVvxwkfP9JXLBbZykp0Eq
oTU4G6Chxqy6UbB5DB9QbNP4dig3H+hBAxOHnGDfZEHouCp5rWNCOFUrpozwz9lR1ZzXbJcXMxqT
5RcAyRxXyjDCMOuzbngkGuLe/U/Ui0SMEGBHBcLBmd+EbB14LC2sv4SuUFGb2Freb03aKPIzhYmH
iK/QrydewfLz9/k08NfRBunsJQEhIqRzoRb2pksQvZ+ztemGfHHcfAixLCl4joXoOf0CdmxP1Gf2
UdCoMpMABrwkhkPs+CbLPxAc/ANeq7z/bzHthzKmJW/RN4Dpfi3vh9ASBr5pU7KqcYZVkdm3WFvW
9/qm6uym1ZkSNqEBXCDCarCsbtCpkKaGkt0lo8P+l+wQkzq4RggOLtLxgkGCCozPM/qWgw3UHXMC
ZSNT4Mmk0nh7pc7iRk2IevVsBzT+NXXNmqplVqmMdV6XN9aHGtHz3wuc7UhAowOIiMHEL1+HClU+
TIvnFrXn3Snagerp9HkMj3Pe/n5LXu/NlHBVfQ9jcAoMkjranBeJjEUf56UkxLbP3o6V9vbhAmid
+BH+dIqkmZRliUQ+PeHySY0WLGx8BNSNOZydy1zQSiLCi9sRDC7aKs7ZUrGMkDRKGLJuHZFhyam6
zpctMfIWq151ZoK9FjVWjJouAeEubBK1o5q6UVy61FWStQemqVxdgjFm4BtOxw6VZ+z2rcuLqk+S
E6KyA9JqCLqsN45vyEm9ybXsY7kr7lDhaA2g5LVPH5fU5LkAU3+drqhCxKuup/ZwtmMNIZ1hp1Jc
RoJpF0thzZoFfJKac0MvQoBbXfyUqqmgZkhDTeFrSZ8rqmbjhbjEawE1Qit+gpRgLc+eD63RFCWu
htbJ3pLz0e/XDVRjqXyjh3j4gDVbh6JrFHEWfTBhdmozP4hGbRHPHIg6g66kImqiF0q3ERFfbER0
LZuQaY3UhUgyB92pyU8ZyD71jKnUgADzgP/01z5mTSrQylbnFY2pDTi4XHLkFT/GUQVYr2wsJSan
sZzADYQMm4uvhSasVN4CfUcdHA5T12Cqt8FvEQDYAaoe24nLRNyjSz62ElhOOLflDSiQe/NHsixs
rkIMkpOfP3RwaT+OXrHHpmkISnRnMMqUwL2QXtn4gdDDINBL/RquBY5VZva5KaTFi6mDh6ae2Ccc
2xvnJoc7M55uW6ADxNWSrHH9CzdC8gofSLEOa5vQyl3ctLrwhlhRfXy+XOAqmwp9/dlBfjWxl/DG
N12c+ua3kfr86VW91fmnv61z8VAT6ThKEoIsWCZQXNRAZTxOnBAOPAXSL3dDVAQWbFjMMQWCo7fk
LWhipS9Ytg8423dfioQDXW0rjoLDjmbZkW9tonXc0i/Mpxagigsaglyt0f1ynV5Z2wa7N0MUmo5e
YjO1K6Co12n3SlWVbKaFQmLWybaYp0tHOMJ692N8Ajfw9IPJI81SAJrmT0oLpl07T3zZEDv0OUxD
rtAXhRyefJET+2ZjhdsmeXriX4xy0SkzhqXgc4kZ/IGBPmYg7C9giNDb3o7UD0O9JWSaJArezZIf
kqIiW+bSkTXSqxQFGXB0N/D7LaJa24Okk142eyg9/heUxWtPC+evHFCBHgUH5HOV6sMAonRYiWDf
lXM0yq7B/l0LbWCUltx8oYQ0AnpceBbj4pHt94bYUB+kMP21Fr+JRCqTdkuqYWo7Ywi2pf9NaA+u
N9LuaUQa8Is1eW+0TQrSxTSj7Jdo49iqhNl93OQug18k9OBjXDYzL67nUqz1eZ4WauAEWA/jgl7r
h64QTz6fm4nOWxfMaRAPvZpMNjeQy/Vwm8dV8z3p1gD8GdEIrCWAUqe6EZvKNQ+AtFdH+ZVdXxug
GBx9C4ohhNejyBAbXIMlYhqocG0oPJ1JyCEGgR+eJ41qNNG3pgjuG2CEt4nhUETr+iv4bt2TdNrd
VxmxC1G4hwwZ2P5nxIqqHj5Y7pZDAyr0PdzhurqF1whUZMLfIDp+mh3cp87mJWDruSOgtxa8HDyq
v8p/33w9W4HlsnHI1m6q2n7tv1DDfFmf8F5S2GvYrySngPQf38Pe6Qi6l5k5Uk8weJpBfZOsI5gk
vRNTKPThZ761tqUk5u1yVOh2STrM7Oz4H0vhaioBdxIFffTuAmhT1LsGoYs/Qsw4JTep5Vp9BtlP
lHoWcgYLVOIxRG8LF3tuSe9PbGdnipdsM9/3BkfmuFo+SYbE4HbCQhSzERm6prCjOocdEj9s7uok
DwMijW/PLfWt2+OLFVls4uA5cV+d8o1+UpbU3ZG2ICibifZDbgDF9mfJibS/HoKe2lNbZRCFDUJl
IoytObQG3lY9cDych0zSTdF/oL9tpr/XjAdfX7jeT/sYqbUKFTMg4A8bwnNp+L1ulVAPHHalhhdi
Mp7/BAt4MK372YsTxca/aN3LkrIOy13AwMOGs2J2+OaAlEve3NJ+A9ia7xy4bU9nRrkgfhzfljgb
p/mGyjRRlzFDaACVnwVSTNsS+m5aeTDPmPIsB5BNyWQv1dg0wqDX21gy9UXbwt1qXKl1LUzkrdW1
nVDuFywH/cn06NXXnFyc1pNiS8fcAIHbnJuoRRgyGEw39aeGCQfqHlOSBXlLPBBe1cdoT6+4xjUH
VPV+9txj1Coesk/H6UXNcIP/QyB1FIN/zwcSLpMyjaktw04g4RIwEcGXMdw6FNIOHG6siTyH/Bof
cLEpRvB1GUowv4y+eFOxAsFInHu3o6h+aRoLq01dRwtXSHAZXmWJidCkKDG4SA9tNkITgjbcSZfB
zNiS4+X6ZLbjaRHYLNCdtrL18/wek0vSKzP4OgbCH3ZyJwOmqVC5PNzCVzEuoXgOgC2u8neguPYr
ZF8QczePvP3E6pG3u88Vim+9FMVct7gVS9jTs0sAYcdr8ju81ygTO/9/42Bv+0e5z3Pt4jEBFDUa
cR0D50Z1tmqbvOKaNZfv9v8WdDS67jedz+QAU/sSfsOUbeakbv2r013Altbf/hXGLlLRF3U2WQSf
aJ27lQmhXLltRUn+zJsCzHsDhywgL8e+aH3ISGGXhgSmkAM+qJOlOMNautgYYXbVZP9eElwat/EA
MhKZ6DZlaIRn8o2AGDkS6wJK+n2DrKSEljEnTa6QLQW9CbLMP1grudQim0ZtrsqApI8xm98z6ZPP
F7TzROMOXe2BawsIqOCBKZ/z1bV38c5qcEH+EhksBVrpFohKKEJpfJhn4yLd/iKp0MqlQr45j8AL
dwM1vEDfEiZV8G2EehAITWLRVgUxl/w/uT63UzXLlBoj6eQHUwGZD8zqqzDLNlw8JI4rTkhq0Y5p
HP0mF9+cksxcjxuyVpDjAXNhl49qnEt5HJpW4l+GJqNAkmQMDgI/1R33vn97osmWKWUd+8yO8Kwu
ChCobBKpqdJ1I76G0SKYKRk1Wk1dqCu1nymwDIsq0h2jyDN1Vssig7S84/83Io8CEP+lhoofkzsS
RES65CQSid6CgMv6uEm2YkkdUGaIxZu/xPJTuU4S9mGOCGuqobtYkC+r8sm4HGksqJB0HRHHGpUf
teQPHO4FnjZYH/apbAGRpdIxINZ4xHwPVw5J/c3wLa3bb8nqY8FXrJzNqk1GCj2KPe889bJmDpeZ
wrkBSAwFWjdGGuNsRrZnwCgkbzoQh3CUHzWqJ9lLovipc67H9yyrkKdLnvGMj+849sZs6KAk4CkC
SJlrov7uc0OfqVJ1XAQn2jXBfydubfpFfSGQmvrmUf+QrqQvfABHsdE4+Iha6/4OgqN59NKVCDpT
LxqLPAzXxsaz5VhxT3g6fG9nnfqiKLsIkmSchGvqotDBzZc8yBm9h2ySVMvkPGCB7hF5VF3bw0Ey
JlXi+j2Vmm6JQA813AKwRKBjZoj3IlCWv4YuZ9ZQauXnnSvFMK+h6oElI/B5XvC6zHNz7eI6seUE
h+6ufyVCcR4UoQMj2AEWJD0iBEuU96fsNN3GoH4kmy8RU+HyjYPC2Te34FmtnABamengP+SoaEUi
ykCc/DQfyn5jICl5221Gtah1g8SzcSc/ujSc5icsmKytAfycF8ptCSo1CggzzgCoEujgiZuT8Ub3
7bxiQ2KFhhkLRJ84jeonBwQ4ao23PQc0EaB56eMUnOuXAj9QM9A07vj1rA8AZc8emiY8nUT5vBJd
I4Hp2sKFGms67QMztQineECNm3dI4SHQ7B6Vqk/RgOCAJw6kRh4g7S+WR6JgN7pcqOLhdPGuUg1Y
TN/Z/u/vy2fDn0u9vdYUuD7s3GtR+yBG15RDdkvmCVeYmrglOH+ow1fP9TIhi6PkZlf5ZF7hy+KM
i3s4Rcnmn6EwbmseEvfYJCETXH1mbyKdUDSuawAc6NzxnhkCHMQRKAI06KGbtpB738g6X4dl4j2f
dmX0Zhp2MeKHDsxk+oDgy1JjY2CPdrNSiZRgTcS+zUVaysDlFNKcFN07gJLK3NzMhTgAyf/Iw/wJ
3Qndz38ShUDNbtPCmQro9MhnJj9ikv+nD+vs0H3f1ROXnm1wz9M2oL0JJDvftcO9uqBbDoeFMDiT
xtraEvHraOfHKyFMlIK1Gld4q6CelWR/kBGBy9K9JyNlxFHOxSImY+UAjikQnM020xyGW6EuyhiD
AheoDVUDnThzwLBuccMIgKaKdzYVlrRIGV309KhzKntIQ2doDxG2Ip9iIlAji06mgTq+yYdbSvzl
LjfoX/feAnN+GC8nEi/gfOAPNUAEcLl+Gfj77FzQ3Jov1/2KlQVmWJXjbuOqFBX4aWwgY2SBuUEu
IrKBm735KQdFd4s4lSDGJNu5sP7vNQ94YGLUwPmbWOszB4nD73+vUR9pAgSTthuCk8m8HCelFZ/B
qp5wR67zYkN17JVY4KHe11T2sGVZekPL88P69sM6tqMLpvmBhU0nGK5gpdLg0/ppDa76txdyUmtG
fdAEAVP2oy7gX6hTA6f8fL5MxGGrlcYL122oAWovU4OhDqEfZdxYde0cHb6WmSEpQ3/3wZPZeY3m
QMIpZVcGWSgL4p/ffWK04GCJXoWuQripk7VfEa+nf6W/GxUYsBCt4+hSiQYGwJLm2W34P3pWziDN
8ax1YCJRah4l+6ODP0+gBsmYS3i60/8P9PWbRVMeUtg/isrnlSZPXQMxFqMs6sRFsv9rIxRkUXdc
eBM6GevNpVbEdhirvxDuAOLvnquYhS7BlyN14fJVRrFmM1v+XywtS/tk9KqK28hcxkcV0B5aKsV8
jJ2N1ZPVS5J1xYzYfAyGgB/9ifWHybRU9/mxNHWuB+/zIpLLCCgJNPqi1ND1N617oTbML7ab59Dj
pPVvTAJJVnD77hQ34O4iDeOsP60vRJVvUWjltpLiipGWTjCLKlQq/CYKADCSGCnx5WaekvWkGSDs
FzZsrQKUqu7vKpqVaehmX2UJ4POhBxIzRLjATiE0gUaSVmqFkuY0WbOlEMyKhTZXcyesvSfnuR8/
zFM98IFo6FBvCRo/OZJTQ2yIeimTd7d4JVCSesUKCW0yniQR65kwdP5cfl0L9WsIiNT5wK+f20Rv
nqwGcCd8E11AIcxXdDymN7LuGIG2dhk1jKJSOZujVnrbo0JSnKfv65PWjHJitu64Le8ofZ7/ZdSz
blXRzt4ZWd6GR+K4BVa/RwTA9vhyKKjsay4pqo5FI0jWqQsD/lXqNSQPVpMnrJHerh/vTXFmb3y6
030FWZFOKO6nQfS7X18kYOaROgbOwGCcslAjEmxbcGALZywsZSDbx0jy/oa9/lWYC4sk9f/kG+7z
ss6ILP4vKcItFKtpMoHTcpaCqWNwX/biz9WHspbRa4+/IzNz5fokLHD+BteBCBKSUC1gHErCHOIj
ESPA8Vr48Qkz2rcQ8pwAAps0m/xd6WJg4mVK4YZYUhFj8H02WuT1MXlk5hvCvJ43Mqygj36xe/iE
NulYgpehqjnllgMMNI2oNG39R84lAaaC5VhaEv3h+FCGZ5jFoYOwn8pXYkNwVve11uR0nj146Ueq
YIOU0xKvQSoD/P6KM23gnDJ3RLTRgo86pYBOJFxAmXArwm5eU0Fz43Fzzd4C1bxfYqXKqpn33wYr
gtLdzcWQwd2Prjofcujta24Bo2ecCi2Q7sC38nUYc1suzwrubGzkV/DvNVo7L0yBWc/J//n3mGXV
4VL8m2W/g9g7oRFcryiPUJ/aQsxDYG+HLJ55bNsgLx4wIYszblmyhSYgH8YdGLMGQ52Hnn/Mrn3S
2d9B++CaHtGrbS+AWX6/hkVnkNl38sDCMefnTedQDZ5MznRhzbg8+EkpVKtrGUyG2psylWZhgk5Z
HYycwXBFA5zM5ou227yRMx/bwjoKY3ZxsWzyVPZz8bSBLiCwbJsfRV1+dAtVChB+3yeowEtsauBt
uQFJrlY2NJRzldPTREsWAYCUbJi77acF206jP22rZFYPl6HDHSdk4u3DA4e95vXWkHo/pUpvxjGl
Zls41mDoOmgpwao2fgN4wp4pH2MKvYbDUBwN8kOch4XYX8E/n9Vvaf/vLsElSkny7E5QccuY4niD
CY+gJh48W2bwKjjwOSG9Gsx9HdEOrAhve7KkB2uoUuBop/CbgUHJN3aWteTd7dO0eikAaCxjw6eZ
74RK8bty8shISf3JtT9TmS7LNKLruLv6u56rxOnrUwUloMRW9ThDQmwkHKtcm+1jNJ2znbbFARLh
vQ3NBQjv1tMpxJQpH20uA5KG0Ck0smIxvUVtwZAdNvnngMUF9YrpdMBSG8wLFl8gXqSwawlIfOEj
AAQxfeTqRsmCvuZbyqxsD+P9wNB7yel5+UabtScXfgIhxDyB5779ROjsJzPq2DgZB/UKdk3UpQs1
+gYg5g7tSTbZQflKn7Ha3zBu1J6iA7wejF/Bt3D4SuQAeE4VtQfn3fhJMwX1SDIkawLrqV7l2W5m
3c5BdneAASsvJXwgL2Jsi8sykriVfI5XZr3Uch9NZhJ4gcv/AgZsUM8LVL+g+IGZagRNJKrSRAwl
aO30U89O/IgLK1w576GJhZcaVr6cpoMfNtnWg4L5ir2LfmrakmsFMMve8MOhb2uEm0lVINgOYQ5E
LBt1NaiTP4lcFhUV5p9UA7RcPK+pszyhxjzg4qUYtHIoFFeu8K+gN+DW/yvXBsoCSmN9+X0M1fhZ
NbjmCsmSV8gXTwbx2Nh6J5nJkZQEk0FXRIPPncNChQVLFFqKEShjFzs0W/Ba5mZJZ2E3NZAKl5oJ
+KIKGYFxdVzAt9xuePJeVVjFQ1On3+VGbjGI3V8VFV5oMKOQWUPzzrRU5SLH0tmcx0VUujsOpP9N
jgv1BxCrZqXSfObUkuVvY6E29Gm3PS77ODd1qUEWFfbq6B2G6s1fuoh0h4yngs8pJYtqdfBo9aBP
xGsDSCSaZZMMmzupB2mKJTh2u6w4I+/vCXwuoFXp4K5cS1hlZjbZVOh1+6sgppP0GnhFKWCmXJZP
kJZCm22GZDEeGOfrL4JKAYAtPWFbsr1nKp2VnwfYcXeg8EhLXNSmG9HCDPD9JT2mujn/74euglo/
RE9vBjS3j5uTcQ3U9JZWF6Qn8reQFCetOKjXNMan7wLfP8vxs0GzPOuiR0KoP05joBtR/+FWAClC
wdjdXIswK1vXkI3663095Ti4pHgAquKJUe9luRYtgD2o3ejLkdNxLIaTuUiJXDjsljQ37xDshOLR
aKNsbqaMwj596Ub+m6hMr5QAmgC6/J9hdPM+xXqaLk4Mg5RZRQ/afjKEk/r5sbro2yuu9TWC1fwU
E5vmBuOGIsuvhS6GN0z624NPiZ9SHut+/9KgtQfh6eyqvuvU4iEKYIvJIOxxC/dowFi5grwMQScK
3PMN7gmHaeJkxUOhK9rxmKgoJnqnxp2tkiJBeoM1BaLouCHLmyLpnOhhnymFZeLH8r0dxfRApRfG
gHqUEtlh6gclqQ0XRiwCkIhxl41+hSAn0Ntgf1Is6gHMe5hU0xHE4C3Z2/1i3KEgXmfe1aD5WbGd
fOAodQQ9UDBl57KThrpgodFuxtemR1myGmuEL7kjrs2x+x/OP4IVM5tdGMdjMs2OKT0wIpdiBaEa
RnEJ6vC6/k3qo2Hq9nQiLz3MfWJBLdT9iHR4LXKkNNZKp8scWgm2AJgPH7ahRL0L4qw4YEG+EDbw
GoAWqWJcGMks/Exxw6Ma1Hf1rdO8n3rO4PX1rHGh2+mG7x7JnfQf4sIi+qBZSqLPu4xIPQgOc3VR
2Yu63xeDLGZh0a5VMJq4YJSIdINKppItyQmeuVwO1hJwt2oglDYMw9uXWCiwoRTV8IQfiXDHEo9o
qiQC3HkJmUSuqeUYFKZehwi37655vgUkb5pdgfIiQq2MoUJReO1RWPj3EwKLbMR4njgLCL+Eiw8+
fLCgEZUYbXWN7DJBWzu2c7vORMUrZtLVEWoi1qvat6Q/mjZ7xsiQI7WQUKWoQ6d6t/W1xAZ35LZ7
eVTxJ6S1ecWm9kPWz6DNFiBqIpSEpKTDZ2l2sXJi8t37zoBoiVLV7yUaiJG+h0P8tFvP2HeeuJyD
zYhemnpY1xTN89aeHRc5Y9k3Xr8N90sQiNa2+7YWuMmr39HJiplbGY0KZE+AtwnmkdL92XO1uhWZ
jTNLO5CSbdqqui4FLFYWObMhzUvNmFqGhNhjKACRA5hIbVgmZ7vt2QIDLeWr2B3PzWRiGcRD8277
gGKlU5jzEG48odXd+a8EBb2mNijSPUtCSk+8JKZ4x1I365Ru8VrkAg1zMI7ndybmtsyNa6tgL9/G
QDBzym7ASq9K5nJHnzMOMpDqkqN9GFvRAfoZ31VHL4QYG06aYF+X2EJ70cijPRL0adGpnoNbFuJu
nqP7H+9y+3zTwRRkC4l7W0NlaItyPSspQWuQ1iGzAW6oKm3txB8dEh9IwBFMV9+/KZ4ile4WbPN4
xiRch5DqYYDv1n/+OhldnxM9jpHrdAQe49gjc7Sqmkaegf8nk5YFcq/G9TSm00vzhlmcn/iIccKh
s9WRo6QXLV20l0Rn2q0+9vWwVRsAlop4jj6tXjevMJN6jPgUbE3XGxKWjqvG24C+B+ei+O2m6iq4
oHb1VEu3VHq/s5Tng4/nTKCsfR4OAwiJjBMPlh4lHTOGj00Tr+S1m03aoUXdivCn1GNglhKDG719
bZXGgvBzELx/e94DGh07b8OVNeZqzh3qR4R2RhRUG6LO6ss+791U9BdWTdmSAmrveVuuHnA9yXis
6T8+TFDY3QM10TMmYjyb/E7XaY/Uldp/cpyvM5Br1h/3aXILqTfDtUF/25JX/HPg4T4qgXAeawB3
KdPvYKWRuKU7Kg2eTk9edKvK4OhsrME4b7uXlA983o0JMRKUVJKW1ukugRYXxal9CAvWPSzVxa5Z
j2BoEd+N6YxqoHEVekj6ynEBFuMqqKym63JNJA9e64bC3LAQFULPTy68xkToY/Y80hCbQsivOAek
klGQUCnKT8HSJwUGSYUCi+cL552e+6v+W0ynvyNguEWi3D6iITygK+7zF+mAJyJygoNq3EUkVDyV
LIWbnSmpXEUBeiRfjaWAmaDgmlQBdWGySHaIu7+x0WoMIfHnyw6//dMnRb49/jeqV66H0WxCrFxu
4sIGQUdxK5PGpm7Xo+pKzCX4OJoxX3LfNNqa3pqS9fO0T1txDXbCfxHBjNC55rG/vzZgIDDf1De0
kyVwDbPGR1gP3orc4a01VMeyjc4KJAFzcVdpddo1LcQY6o8OPlkDo1ZjppBmWrZQTA6CENRmAU8F
4RciEsEfrcCLt9/ELTq+n+YXFZVe2PviQdkVybVAmcJOUhzRS4dKnBPzmcZMZNP3xSkmz2xqI3VE
Vvz9nuhbp2rXjkLOD017QsyyipASPL3egbLBQaSurMDZRB6/TeWMo7T8PIzwKmM4wg0iTF5JvzmS
rsaCzrH0S5f7N5INidbuKjJQKAUMrZ6ilTlJ8NzoHkczQrv4eYHpiiDjdvKaIxmTmkcrFDy5m9WI
lpnPc3ihLLWKx6nx9NESAIZArBt8XO+w9BeDPZ5/EBxwbzjNj6JTyAydtGL+d7keLS4Jie77yczs
0xptgd0+uNN9QiDq1uA/KeTWOZBnaGQ6GtN+64tDgCkZUIuDLngNHnVn6N8aUyUN7f8Nd5sahAbL
qMlayX9hGIaAaymopiSHaxzUIx57bNncfdg9wl/SLnty8auGflRV36PYYOb9sTwJ1iXUTj5ZkFWF
rPcduIMv4L+hkpY/G8IMnVgUScpfW9OMaU8pqlWoED755dOrya29c2CrbppNkR5JBMN8+rm9EJ0t
n+ip3mqK4NMfywUvYjQmY0qqafBMLzTHNgBDGmtXp7fo5YzXB0SaMroANHUT1n1lT9WYPldWrdYD
XseifVSeZipLqKED7GA4MRS3b481Rpd2h9tO5iBjz2ZYwsEJc4s1An8bwl5CsUTOInIqvPx53NVi
y9LBChgmvRp3JDLjDx0ee2k+A3jrCGtlTpNILfovij4Fk3wGH8BPAS8/+lk1MywQS9evW7cRPYgl
TG82kEisOcH5l7iNcl0QqTkYSxg0kafV9/siWkeyBh34Q9KINoNaVqRIjYSsfVkBE7jvcp3sb0V8
Q8om9TYZe3uIqV+X0bbp6/n314DEFHNl/A1Dvk3IfYwj0khM66LSehj8dlHzJPn8nVttNg6D6v47
Eru3V8hqXH8u2G3L2ShZviepyexLCo2SSHflzqCAWYEFLElV7p3gHHkpz4RDnyjbKmkgrqrOJXA2
A0DkvJT0n5yo89dbkSHy8KwSDiMa3Vgn6Xqxz+Vwj7D2GY2XsxOZsizeeCpzCqBHstCnOOBmmBPE
Nul73aG0Z8VDI36wzZh4vUGcfsRa1Xbv6ZjufSMXSW2W8aSiMvDKk45ceCXSXtPiLHzEpQ6ly/bF
k+XxMRqn3Prbkal/UaRacxCFNf0TYfNUCe6gX7dyVMapwgIwod8ZKucRDfRzkM+KcPFjfXsAHvpI
an1D3o+I1fiHjToU3WTRgS38DDyN9i2Xyd0ghLPbyjHgC4DKDz8PPORcYMDyZ/8/l4vPD0tFu1Dz
ev2e0lFClz5hCB7nJ9epkgTIxVn2NPesrQq4quDk1L1PwI5xlkpwTPafB6xUE74puBRSNjhrLMK4
bUJuhKK6KLHeCMfWWAlPnPCsOYdd64hVhxnR1cTGS5GWHSwAAjpm4lrI0aLaquRoWMnvPHGP+XbO
8xACeo9FX4j5Ox342UZT52AE4vbIojrzKhSJXIN+ye9VDmZD2GJLMIJ3pwikpI5p1GwrWEvanL4m
GXn83IEC0Vpvpum8+nrkXU/gye2K9p0e/N0hd3mv5W7wlOIibDhHKeJKyrOc9yyZYU+IXfkrrHbv
1986caXjRTXrdX+wB1Q8KF03E+maiB2Y1d8Bao9pvkAdMBEha/8Gjlatt/5p6+kzCKuKi/OI9+GI
mOawwluzLotIO4HVymIXdzvT0x/XMHrgkjAs6ZmJ+8NbhGs8EGT8j0CVygddfEnnrraqxg5Yx3wI
wgoS1X+CCJmXCzLdKyP/TOgyCIpznNdO4Xf4UF8+85JnXopBPfq9GG+4sIXTa+cmwcxYEZ78hcyc
r/47fIMya4zM8GCemUY69VoyC4TN3PXf6fw5yLon1VZi+Wdq+ruj0Tq5vRd6GfsqpxBqDrM/PmZ/
kGJKNOZpq+spVnysdOU7/n9IRu6nV/+lTB2Fd7GdAkiVmdMm422OcZgEQDghxCSo2Ib6fGf0UmMg
Km7vwb4Jnz7/us0L4Iu6xQjNl310vxrEzTj5pssaRkNEdq0REBZUaYAkQS7HcMUGlCHQT1ELWaXQ
EppYy4bAmKG77+RPmYjtw4UxkWa7N93zDIpQCV1G4ym1Mjd+bztM5hN+HpX6YB8rErqPgIohmZWX
AToWhHTu00StuxBTWvPietat/czIYoJ2SwZiJWWP7PjJt0PFLk2T4lCA0CLW6zWPlIOz31JOQUFN
x0Gc+0JjRn4kopxJ1zok4iS6oXMpQ6RBKtyMT1e+R+Efu8Es5DUz1zyyFiQ3XjG4INntFC+wglXe
aauggcK/76NvwFS4isrs1MQLFeXKIWtI6BF0+OMAPX+9mIn/6+K6Z/P6jkyBY726pHxMjpr4cGcj
0tqYE3rp1hYIU3/+5HifMJ9AkzLXEDFNJ2VX1BHTv9TC3qZ0e0FYRpCyGS1lOphlAN6y609a0ykF
jMXYO6qA5YN6T8w8Qcg/Umphdt65FTCblThbser2ayYmVsisrGdU1CL5tte7r3luRQbeLl2jB1EX
K1fbi7riz86iPL5Q78pVyFNyR2zUdcIcgdp81i4m979uBdnDwFeEoqaAsLDaFitfcd5KYl2Z87xh
lC77DvIc0wBHpF52AIUBlHoWtP+t0KlrK+r89z5C8wjH7jMvY8NDbjMRsBU62Hy3MVHfg4rqTBBH
ybExR8qAgdL9epq3qCElqNC57Movsey84b2Tk528Al1+xoskSLn/gNPPr1zTNibQmiNlWo3CeoCm
yvjd2IlRzB/+SC/LvosY+S68hx++8q7ovhf5+KF5DM9SC83t7Ufb9MFeG7+0NeQygDc/CzjU1Ei3
Be4o+IQJ1vQNonP5KRZRg97uT+oymo1Qqh8SCsdG7F2ctxYbbckmJykBTFuwsuEk3QkL2mFxtP0h
KMroLQwxPMEFMPGe4Tde/qf3z7Lg2dBb39jtOh2dtO4os1zj54e/G7knxSu7rW1QMXGTu/cZRVDq
oX7+r6oeA0nOgCeZw3fRlF4PLq0UnNi5un8jkBKMz2rni0+S90/PSS9Bi1zr0mwICCW4IUlOxaas
ga5NP8kODYrRR3XqJ+aqDffaPj7ruGPNM/LIBD+xbAETjMDDKMyJqMOi5b6PoquqnKyX5NFEM39z
YtEnEbHRUTuzVvYGDUh+A+yL1Qs9kOUkmU+CZJBbcpG1d+iR3ojRUTKiOYCkONkHhQIWR9AC0kJ8
VBVnQY/MqAzS/dZgsoGdf9+MVydN6ZsQ22Pcv6Ly+/zY2ZxoSP1ofNaF5ptnzbzAJOCq3dUy+EMK
IILXsAFvUbT8BhMk7Lo26fjmPJ0s3+2hEQfz8UGIuQR3Cphv+rUNYf/TzF2GbYhyjisVFVJQSdqZ
vvA3GRK3CpSXcaeB1znNFf3k9wg30lScSjNWctzMU5t0O8lYtDmVhhXeenabFMl9IXp0M02Qgm9H
GFUNxAtQUh3TdVmdx+VQsO3cGwX0DAtDReCQy3Oc2PvHrWVclOa1+63m4ndLYIxT81s93gAV2szE
KUtmIBlDAhzDLhldkKKoXLWL7lRXORyp5Lr5XoWu+niqrXqL9KR344CeQ6RA8nsSyWGY9GQq1b3H
XCBX4LjxSZbpfPucWlCGfN3Atu09+Jgub2p+MBK5Uf96s3vu9jTmvRgzsSOF4tnbVR/jiT0h5kaY
ut0gAc17cIzsAFBRZprtxyybtUDSjCX3p17tOpY2QpZ1VeHHhdKSDP5I/YLcV9hh84Ky8IJxhFqr
j3eD0Z0kRyCs0LBU/9RPCmje+hQcyOXSPcVYmYg7Kd9envrNjLbx5SLV5E2SilAp2jrFWXTAO0Ev
a7SSHsxbnv6mrdYhuh2ViC+eh2LIzgbivFQeE0cIMPAyDaIIMknO6rBOGVU0ZGf4b5/C8rcAnkdu
DoTd444pK+bPXioUD/DZugDYfABsshQ0DCGM4LamMZVB/fLodRDGuSZ/cSaNbMlcGhJBnqMrj6cg
S+oaHl0PC6r3bvfl+yAOoryTpJFHChFsVgyx9807p+5phTMPWnkkAN4YLM5eb4ufhaVPXCFojrll
rovNDOcGP/sU4W+HsS3GkzDE5aYU8nL0pdtgU+lR3fmx0IIrDAfeH9ZonIeKB3IcFV/fXaL/iGsu
zCHmNVErKD1QQtxjUZonQN9B+prNV93sKX5tK2GLzpdvwnnPK/OKq0CtMgdstKKT53RqSxYddhxS
c/0mPMqv+mKchg35L3ZGbTd2cUfVx/oD1ZvBYUNr8AlSAmBePuf/rmksuqmvOCLpqnvBG24fCmzP
2JZlaMqYu/7BKT2D1ss6CF/PVCjpcACW/rvU9lIdjH8Nvw7rBc15PvtTMPVeU6MGgHW+PQGWctxd
y+gPN3abdNgiLVRrRVX54UFD9Yfy0CnW9DrtPAVB4yfYFoKu1EECkg7UlSpZCJmWwbl8XKhAk4C3
2CVVdHtBEsp7v/+r4DtDWhdFr+5Z4EcQAslWAOegXZIFXsrSI0SdWDQjayUVoCOjuQtFEqtctfL1
yOu4QggFeXJCYlTBu1gl2W/GYXslszoQ002bC/x1na3UKLLoEyggP9EaXVT3VfrX2HFn1eaPtcH9
uIgcdvlQn7OK5UodXcWv6UI199oovK7blTPPXZEg/t7V8iDWMTYI5BjWlQOVfYyRAUSGIFpHyNrl
Le+QEMDl3CJPqunyLvWWeIylyDpfQJgrrvK2Dlyt1XiwvEHn9c+gXw+LEid3Fg+Gi3UXUQJNYk8d
K0tlNEeYCwohMtXmaq9aLYr/7PhkSou10Mb1vZMaf+mcvVIFkwZ+OGxpc+bjC/mfxwoUV3C/v5vg
kbOqzLv8liJ+1odtMar831o4sK8Vlx9dpG4WA8bBgyOcs6agGkN07tS3RB/o2IUVSkQlMCHemmzf
r1KMN6Uniz9c7t3PIMYUnHlgn8WeUJcl5yvePm8SkePyutyuo/B27N4CBTX3ilbDo1rIh00F7IoC
XhrcCgZTjX7s7++iwcT2zFwR5JOacx/NYyk1e2O8L7nkwi1WlpRrHKjlu9OR8wK0E3Mf2zZAfr8R
XvJpBhGg+ByT1ZYLtL0/4LvXTQdsJJ4Gth9X4ONFgO4G8SP/PL1UjF68GXtbiF65hdwFITN7M3XH
WwA/fD7wmhUe9aH4c4BLg2ts8Bz7IQF9fDgHFQOWDcXO4kRiP36z2pBCr44PMvqpy++EKJGygi8g
5llXpbWRDeEX1mfQIZ/1HZcplo6xIGb079TgvGRq9I87WQ+UsMqFy59xiDkWYkDSL2plHsMZoruO
of1QUOKfE4r4NVtGIt/E43tS6KSZijQcC4QAvoH3eEJwqAtH7d8si74tWfFGDh/hi+AWa5+jZKJg
plMYlE3u5PT42W/AqRi/9OjNVzogG9QqszfZ9BPAu26QTBcu1rkXvkWb9sRTOqS6DNI/pwRxT/Qi
DHzioe0f7u15e04lTDkLX7DKz5VfwmLdRBavzAg07R1KtPCBO53I0KhmfSnm8QCMupj3uiF9kj09
N6vf9gcD31bLGpOpANa/arBG3h3iRPlIhyKbb6wZzB+SUbDvyg/0cYXsenfLtRDrcir4PW0h16vL
/sVSv+sGeYOShgSp/oM0dlh865D+bOKWQWe6gQoWaazE5Uzgy9oIyMp4i+R+Mm0I3lfOTtqXPJS2
Qz3ZsWN9nFj1ZtbPf2U3WdXDvJ4RgIB2g5X83ueMZlyMUlcL6o99axVb5uB8ia225YdfTSK1lMWn
piKjYO6gi2pMqE16FNsrumXFln3R6cAZDZrT3W9Y6/mOEnhdHDhq8Cn2TK22Kswrbpjv//XTQNH0
UlqyPzlEV7vIrG1fEorUdVAgpiuGiEjygPkh2DEvJ3+QtmahNn/4NdaeuANJ1kcwFsUnbFcKr0X6
lPpM01xg30zAVrUCkRvsBMao8odn64HdwsCjX8pe/D4mOLZVHrMjWi1++XVhz1bpzxAD19c1RfW7
aw+7oa7MazQC0Bt06qBsYAqyUx4VUlsC99pRTAOGEWX2Mf1P0rsxlOcTfEFwrhZhkhqNBSvFeL5L
C/LQA7Yz1Ak2z4ArhhfMTNbaJQPwqJdxReqteyCGGpyJs1iiS3NCXmkjXWqANU/UZv76aBZ8jb2c
eLSMBeSTO4DH+uto51R5g2ef3j06MyiE4Yo2dTH8TcUXxD4j5apQ1GJwDu/FEbikUPrX/M+Ur0IS
m8xMKfTFkp6lvdPDYJwHZnPGA0kJrgM6JPAgFvd0nSVNjfZ5DwblNvLbL1uFdEsgMZ57wJEnZfEr
umgz38g2n3rZHlyfBp9ktnU3ScRKablxUGtztlp7VtNl9czPh39YRL+GBOwu0npMMq1iR9w2VXUe
jYSxlCREssVlIMa+pXUZCUEyGJXioQ/ZCUfqx/Q1ot9XNTOFbJV3Spf30j+lF4X5SGgHtdsn1CUc
6a2mpg/F7A9Kb/7XGVMjSf4ZxjA+2oJfyq+ctVewBvsWcHXHMfocquO9Dd5QzwNngFDJI0mhXbWY
JMPybHv8ls+KqaBWpfNf9iu5nFVudNF5XazVKj9/ZH+eB/9AoMnQEE1xGgpS8ccX7fnAjYGNletQ
X37wvUBJ4dvsA9crZiC7Q/94cIxVgphB1tdQkqAny4hfmOpG8gWzJI5OTgQZO6sx7pf9RNwp71wG
A1jmhzfLL5xP/pJ/3kmUEaDQIpZWK/QV/OWf6NKXs4i9hJlLz5gC64GmcKbEG0JX1+YTgwpCM0Wh
Tvo1iA/8BcHqx3FBGlvY22m1b95zu5kvuT1lhmeLpAxj5Fs0B+mjAVt5bgV4Ac7EoFGzlV+qYua2
tPo/thNFKMtqiwLEDyRufIqMgGTpfcWk7tqdKmYYyMZEIitFUeYoe20ViN/+rF4ZMDstLPGTlEVm
6puddTPYJV3BLhkMjszIQFHE3wLRP2zj1BYUgowm3PH7KVrZ15lRwrz2v68gFDLslB5gSkiZNYeV
ce87gJ4fjHcTXKwqxDyhW1l/yGUpWvl5/fFg4oegiZRwDm3F6CqO8IkMVPShN5oFut5f4eSp8xsl
MPwxyl63gB3G7bBJxkmu2LRtvqSUyvW/zBmWJI+6nlUTMfLUnleMhWlSHmQKPCGeMzQkVOFCAkog
izyZwO7pxzpziPPy4WTysgCR1ISx/ySpTGJMLLjEMaeYplLEtKQ1MJaEUckxHEC3nCjyHJUhZquw
qW44Ke/PdbQjH83XXQ0vYJ0bF351+jU375ql3zYs8c15gw4WmHmAD3g5vJi7U8LDRakblrpfXW93
k3mk1PBWW8jePsf2ES5SaphP3NIV9N1uVW1iM+ix73zoPV094mKQbV6ktKlVkUX2XBvl/SGPJ+pm
lK/i+pn9f5ZgJYplWPz3AV/hLMVggnXwVPMcw/Zk67JKUxVUTjSQeAsyCweFAXSShHmZpfcyOoY+
9lms1RKzJDh2Tqz6xoU6h3GTQJ1kx/IEDHo4HrmFRHq91Qo/1Wz98aPA5tQP+SBYFevuBuPfTwOd
qyRcVsUATOA11vjB/QMAuZMJTDU4xdS0cg9evbpcf47hkpg/OiIml7OmGKXvmhin35oXAfpjuRWZ
P+EnGCAdUjr6qg4FgRCLjK2ymK4MYBdOe9jrXG21UKzNPQWsUGsl68ZICSioc/37wnurgnP3k3Z7
Du/kH9xffv/E5Ir9Uk95toQZilc7K2N6ovUtOW2XHD3308vjOgv+SiCcEmMj9efJ8bfNfEdIApb5
qBOnosEVgKCwjdT1qBYPmRBJkf7ECcitq2D1Hvli6w9UK7yRQcuiIF1olryxvxRsT1+k94zc6o0p
EKBtWV1ML7lqgE6g/JtBEOzDso7fUWgbXiFnEScXuperJguTsoBHSzsSmvDsPJuzTWvATzGDku/W
K78TnSeHtA6lF0P/BBs6iEr8MiYidZSyKHk2Ckflw+8JVzYiwG8XCYJGMwmskkzgAw2flkzeszvB
x55Eb0gOwxj9gA3L3nfDlTeR9/Cag204FnPW9ssn14/X8ZpwiVZEBTe//SQCjkdWNwrCu3m1UWHW
A9ppXyzm/PkwrsWykz0t7DOSyPyyTjGyAXP9c2GvmEhGzDr9YXZUVTH+487BFznSI98iuSnCxzw7
Oo8hEHZuI0KT4OpU81f9MRTucjnPkr7iNoDv0OqXP5b3CUsfpndO3eK/9M0a443uoARuLuCtUwiS
CQcyJ+PSMa5iI9hP2XLOXnsR//giImv06dAAd/B4ha0nWOu66amkziTVeSvwd3UIEnuMV6pxA3JZ
kSIPCStVtNN2kxGhoyW10qMU/9TTMcV1PVDGvEUEnhoq9bC2X9+byXyzHTLuCMN7oVRFMaoAQHEd
/bTvd7akPrcIepmI+XZRamlPJWBbV0HkfjZRBemnL1i+l8zc0bE8fKECexsyND6sJUSFnzCrGnWp
zhICutbHvLDGtUjEivpnh3rZu5aVsRJNHcij6o8P/pd/TIPk/6FQ89A820IypEUpTdYyzp3S4KNA
XtoP16hGlUf2aAKPG3zxZeWwcdWCRKurOomEQnXldm+E2sxAEMKKoNEbXUTCCCAIpyQxRsOIr7bx
3iik5hcEoc0VnG6jWLXWGOOFMvLyhojLRLoaUnhjV7eRSw3s6yTjMwMM+NOUMHu2nI4iXQFF7bBu
iqoyPcdrTajYFZNQzzOIJe6QvdzXina+WWww3J+5LYKBOGLqZYQ0dK1Clh3lxk9l3lDJoMg+Z0cK
wttfqwSrPVqGCr46k1PUGqMRWRuE94KrfoUfJhZoMZRFZ4j5VzVzaV3KFyWyQY1A0b/H7lRTG/dx
Ytq8tG6Kkpt4/Tszx8krIT508SPcrJ4LVYyEeTrgOzWw+DpT8oQRMVNPKKqxQW1qjMTJAxQroQBk
4SQKcEybwHIUhdSkJLiDZFxlfF6E//hJhVki7/TwvX3r7Yq/9kziecBIupQPbF3AEPXMOMFUfkXq
2BPl2Vx5RHNEBVVTo46FDaI71Nbh9g3rxcfCUaIcMuO8iijEInGT7NvrbXZALHwd9H6juGjIk7zO
OdqDcr9PxaAbeLvya9UAN5G3DxLPxFzrMr/j9J1+5EVKjWVhhK6lrdRV6bQSfKxPQHtqFQ+q7Ijs
T8GHzZBlnVJM8jAt8MAxmPdtLdsAF7NK+l+M4SmivPfTJOYVbNajSohc356gdDyvrcN9hMaiILEm
2oGEbB8Ri3SnL8bq+ZOVFafjlBxYQhk6J43hHJQrRsKRhc0y0r05hKJwpl18k98TjUXtNlUD/wiU
2kJFnzA4BSFikhxUPokvlt0BBLrSeb1mA7nOhBXKjAWC+fUwcKeJRX5Lkbmbtt9UgP9HS7RWFxQF
CwO6EGmWlZkZpkznPH+tI1oZIqTCr8Yd7K0SIxifc/IJrJSs3bD/osM+x+Wz/YgPcssVxIlUnYd8
s+YWwYyNrPblpbIxKS05eH1FTEbc2Ao3uY1sC/E9ApEW2c/n6KJZEEqQmSjAHnE5oueTiKN1SD8T
R9vGXZspUgRSKCo9yvgIdDDWOlJHbZZDRpX5i87eVH9nc2HFTIbBVXRXpTcB0Wb8lT+JxgxvNPV6
49tTh9C75nQRQKulXDhXT9fhOXGT0ne7DsD5Np+A2H/oNblqfpXX03aaJ4QhI9nOm/UjwZ5tglSx
QWkmPgJ4D/OzQGW8ZWu2/9C/Gi3gW380GQENlklZX2fzFcFutQpSjwwih1roKHXxv3TLCC4/BB0i
1mNkAPAy81JmPLu8SNcY9CU471b/lD65AMumniz47bx4HFTA0WgiV7pScL3FwT+TVMHV5dwH5brW
6pwl53EEeTZJCNTMaDj8gv7lcRkbzD0enOOLp+Qau3K0tZNc5OrL/1Bmu0n5lyL7logzBQyazA/a
rgdx7j6MysnV4z3ODCzmVVhQ6hNF09LFxwALo3hJkeDdOy03lYoRfvD8RFY9rXJGumkYdAoEbMuA
0N96N4H/nRAiYo15u9Kl9Ymb3P+qL8wveMluQJSWYTKQWsKGdSXP6fa+t3cUnA5C3Nh8u/5mirLv
0dElUbu2/Bk+y2vYYdwkjv14Kd+p+uKcWGj9g5My/xWMsulbfuOivHcY3At/Rxq09UF96Y9aEaAC
mQSTfPaxpETpQX0YwKdi0+KCYtayClhHliKqdJ8D7y6pbK5WvY+TJRbJC1CROAOdvQJYYcukU2CP
iEAvuHSdfyHcueujg0jIs5lSmlVZgDFMdgcgp4xEXJMEj1aAAg8//sGRAR16vQDofhIigDSs7qyk
U3OGxH+biIAf17yWW6C+Xnoahp9kGadXWKx519k5z70W1NKgBhGxvEZur/zVJKiTvFJdQfuyEmw4
IjjPkT5aoam0r7TeXhmk352PJJRpJM2veKkhedw26NCMeafgXGR+JtsSjDxaNtDug3z2ZbIsUG4k
NSSHcffjETHBhsu+PocgCMaDSZCXKz+VwdUM9xTnv1Vz1Eyk8oh6/WIIqCIJG9aFRCa+YMFGiKNn
gFxy1P6JBUkL8L3l3jBMZtDilK+pcJD1i3JaobcLpn7KfMFOfoxm1/E0P2Pm/KXOUhjMCrzIS+/j
lPLEnnYA+/TqYF0AkVGqmbNhaAd9tY8YjtnMsNhNcn940afMTDrCxtTnXWX4mNabCOJfZB+PYnjK
5BGAKSYZq6adU88cUtD54o9I7MnhXnGp9tSnWtK9djyyPxpO/m/owzfd1MTcnnL/hee5RvReA69G
8j0uLOFIHOuQcuNpwUGcl9zyxE97Y20Rb9+vjnAPyjJBEqAgcY7kzEsiJXQtUHhziNmXlWY2j6b7
YIFtbv94G53E9+z1DRLt9Tu+o8Jcv3C7H70n5NCmVHdtXqAH15vWO3VfKYOGzGZ0S8LYnSzv2rx4
+gW7YuzZoRNCpuGxnKa5MB5CbB9oH5q9mTu5j15C+RJt0pLFnLxaW+5uj/LM+xu8/ThfOd2zk/r1
fRnNArKVr6X8cJJy3QKBFtvWvc74Bsk9LaOvzOyiXhTSG0MfF2bD/q3/llfTZPv3LuIKwOOc/iW3
wxrmeEiva+YtHGW82/SEOHj+bDkwzDli6mQLxxJLWjEEC7QSx+CP+nEKSrhc5JLV7sJz9OHnCOOu
s0t9Xgw56E+7gqPyqrXyYnnE6FWwLvO5WgSiYSfkh52W/kAAYqLatDXIyxE7TGcdFGnocbbkP/mj
Q8xat9oxk2XLx5DkDzL6p3LRQh1GazvzTUyH4vAwSFBx+c+FF9LDGKPgy5MIX2esr1o8uenaGksH
aCC6ObitEu6LOBeJGYC2V1VQ9SeeCiCnlSziLpFquSZPdBUL04Cu9BlLcMYBgget79HWhJGJM5hu
Cpmb+m81fAlwbC3HnohnYElZgZumBZq75/8GDHPGrhzBa/142TEiSuJ5fQ63z74Pd708hIuUeMz6
E2J4bdOG/UZHm/8R4hAA5MXxb/0HCNdjQLY7gY//HbORNs4c2wz4NyoaJXHTYcKI3yYKCJbA47gC
7rPOuoXkUjlj2zCQXqTdJlt5SpcqxNqJfIeWOUHnW3V+xxGg9vX6Fq7cQeNhKPoZupcrKjjGTxv2
T8Meaehlcd5zITlKWpEVAK6oUTq3IWMOOPrrrZBSK+XEoLi8Bce4rjp0h1M15Q9VkHnNk5YIsuPe
1oO7+wgwCUNCCzFbWZ89jkIdrbRBptgrfNKnv1n8OeY9HpR0toLMaAq5q+SBH4zKId80GZsihJ7y
JHQDeXatSeE6v/nY2qYKINfKtZTwvlo3Ax8GdG1ivGdW9upVA+B/u4/U4/rFN8h5Y1IKweNQj0PO
h/PiaUEN4XcDMGrkJ44lvVKdKZUsDBq9CJQzVRYkytTTE9IKbepQqiXPI2DmmxMG594JDkybOxrR
WD49z2TzECxTXXK8UXEO3uiqDoHIU4JrCZZSoyEwwFJNthtNJWjVlw4dPrW4oQGYcB0p21CCBO/8
3Wx/s1kebJGy2+DEP8IJAsqgcHDLAeld2g/72GXxc5hs5XEwpm29Dfua2csRjy2c7SQZfc4n/2Vs
QK30O/w5sEZHjYTHPRi0wji/V8CitLyI/piIdcCiR/93XotJLFru8YjdMIJD8nov/EXjOt//xoTF
A87A4BcVF1xms36RPwhXtyi3ooGLmGQByMcSGjzn3O7o1EjQMXdI9B4sGnPVFDKbQtfKVcMItw9b
uQvIOxOAUrp03mGLkic8Kd7+oAEWoFvgDDdO06Tpr+ZUxNph0zXXAM4SQQNVt1v0+KgXkMfj3Bkl
AZanc4VLjDqbnn8dwRgwL9BE4MzgRHhPT5t0p4P0Nt1j6fBcor8dKRthgi8Dpm4lFzjyKqXVXGUF
yMQmB7UEj8Vt04t4fcymMWQd2RxBRB4UKXZcL5JocAbOr3eLS99fCBXeno9XuZZPNEVatXk6QUqe
hOOsIFcjawSNxvklt+3QfoNOFiXEGAo2lryI6b9G0BwkKalKN593q17msQHk1lmMFzAoJ3PCSfBU
TaNM8YvYDozBmN21E6pilQAMv1fFIZkM1jkFUn+aWPHiAhBsafntBcBXkriPWfuttAj66pXXEsVR
iv1D+aFMERkTVCj8fBmkyP11GWrffwYej5Q+NYnLQbnILCGfC+8J+fit4sdXuKine0p5ZyqHl6i0
s0w66+jZJ4kl7ArQ2/0LWyTITjc+H1D9US0l8pJGG717fDmnN0Mwld/v4oDLT4OHcugtWLmy9Xvo
EC3xh+5rD/aIl86zQfhAIUIJNf6WPlXqZ8WdsZr766/9ljroMxz9CFCIfMaGVvhHb2VS5a7jjoy5
bB04EcWCdtYOOxz2mppx6xcSNSiZFaweqm9McZw2LiY8td1h/dj2c5HTAMcYp1W+vfNc5RiHAXsz
SKMzvRc2b8ukBylpVsxYHD20VcG2L5l/26Z5urLz5/y5rchBr06mJZZaZvnl7gIimlqfO5bIYF2g
eGvUVdF0MtD0MkiPrDegcOt/2tFJHyv2tfZAIYb0IeR/xUEPvacaMvH4rBymNeOqT1nI9bXpYWnd
zJjoo/0TkBE8nhTth/bJS1LHiiwAYajpDHRXPee79OH/g1VZOcE9iEUAupFY/D6nJiIJIFusTBDe
TEf0wS7TEpQCpZmTQ9wEavH2xLdnh2CI3XPTiDMbnPI/nwCEZsjUBISGNXWpKXVuTAcmxCFZKX+j
ABrTwae1Zc5Z9cfqHjakWbVgJUcwLJTghnAVUQ1i/0+K7a7zN92g+IciKVtCy8yM7qd8yIcHe9XY
vz/32Rp6VlrlCVKDU5vt8AkeQEb/+Bj4peWpvQT/DkFmN26CQTZHtVEF++EEnfsfL/s+PNGBaoY8
mh/qQZ75aKb6R6ZYEirwQPQdCIq/7d7JlJ9tMaM0Z1rlee4bNvgHn9GvpQQ2m/EiHoulOEmTBEyn
s7sbt5ZjXU3GrswvPhbokdMmRbMowzQ9F3Zl2zyGhRT3Dlv4I0LxwIDVyKcIU1XRDsOsflEPAgjC
UInyg2z1DC/1ciN70VdkMrJLIiPva2nKJHCOqrHBPLc5SpI2oqnY4IYpo93Att/WWC13k4UjRMZA
QC8uSk2rldk0CqT5Ji9xfiCL2A5oy44Zj42GfeqkFE12mw75z24TZQFRvmtisEazCiJs7R4SLrde
F5CaaL0EQv3fCbO0TGQwRW/RH/RQtz/W6PR4lWJmWM6r935HSM99abeIB/1cgCQfZalHeJxrSjnu
j73GB1ajvjbWlwAxnSb+/HoMiyV7Yw/QYmLY0LEjV9K8ottQaer6O4D+16Si6Mtetyk7LOEaoP8F
yNs8QHusyTZNycmn+ab3VpeNnTAkfLuEMniykmBkWY/86KI3X1HZm1FlK2Dlnzp8SuEqIpaOgAog
5CtnV3pTXPPhhn5uVUSJXUYBMTOuONqcd+xBL6yu4BSbHul861lTyDHBjVHcVFF4OqC+K9kMuCD8
V1RNredsCcVFV/w1/ret4ANEVtxOHUJmyx1T8VR0i+hYw2CgOPjT2fTQCU5/1gbv15DdGrHk7PTR
0/YwBWMDCcFqGhWoDxO44srwpDIxuZY4TUow+rxuKDmTBlzl3sKXO07uB5cR6JHTgfOW4okh8Q8d
6HNExgQlX6CVcPRmqEtd+n9INXbJZU58kKgV1TalcEmCPBaqFV2NiKn7HI/I61ADAUWYyzYWGFv9
IJqFic9I1PnDIOf3/D+qw4CO6yvlIHlxzSa24QZ6wes1sTjUR9zT5Mqb2kookEmGUKDaqmFUk9eX
ooHoK4AzJZuTaU6rFkVMievl+bgD1spDmq2J9bFTu7M7XgSpxlA4Ppves6BI3E3Z61RwNjAlMnJv
Jne6aKcEr6ZSZ2SG3vxl1tWqYqfUpGbMvnP/KiX86/nwFHmZYYngcceeg7xajRqI+GYNseM75Prc
Xou1Zp+MrbRXG0tb0k2UYOAwRRYaeOS/bQifFwBgv3+JvTmRYpJP+YmnWiEzRvitrtZY41pSa0Jr
yF9Eg+mAgMaSEpTcvp5UJO/uZnbm4PCCswHaK5zSlgZJDafoGqV0UGQe7DUsjXe5dR13wjRqNFBk
Pf2dUpFWLFmXEAevyFrXZ/xAv2UbFNEg9cuz/6ZrlHVpR3J+maJxeXfRFeRVjZC9+MayqqEdZ9ww
EkvIg26JBrcgdQqRI6SqxTcttcjbWLyvL5Ofbb8LW23vhmkMkX2osaDLywj9qZVai5J5uvuVWT85
1lovlGfdjKkgkpv8s+74cNAO4BwuHs/Yy5l+mJLenCESgGSOww7rxajpgp6ZWAAFVQv+1/ogKo0f
6t1RVxtdT4r1DXEPPjcv8dV1gG4sFRPfgUjNY6bqZdUIBczjVta/po1qJj3a/waVgJbxsMG5S0cL
9XXhjffikCQdCYjsUPHjaKpqEgBjLUmLu4NnPf53G+sGqaZTLU//lX6fA/X/ltQK7XJja+L3ugyW
TQX85agv9M9fe4fEiSv9rQdGJWYvRaCo7TTtJYM2T7LT65SeL+iyvsuXTmT7j1TgpSmnQ6Hvnefu
8Ouy394Gnbiq9uVJ34bVGdML2ggdu7o5KoSwAwidzUlOU0TJOjN11/YP0m5WyriCQqmQpoziixXr
ifW3A9MAPAIDh86chqIjOMnHWFoZId3KuYer6zUt6B6PPLUz/F2SMls+UYO4Qt6ekppXWN3yDgni
g6CZuD3DnDLQ6fHzJRdfQAFDgd1aNbXHupwCGy0M7JprqMcrXx2PcNhVz/h9fcuwTCJqldcwz8AQ
y5P168FQOHKxZjwA/tII9PYJTo2niXDeYVWYd3kOa9l9LN0lcDG6alJbu7Zv50ra12TIEfGoPTp1
hHL2XHZSdMyFjw+nRsoIT6j8+RP7iWiHKkVSGo6z9C1jFno0SgqRnEIMF5r1LGTVfbQ1pUg0hhtB
sTlh9iT+mDv1Zr0j0Roz2qR89BYbfK2HM8UGmk7zRRhWaVz67+l9uRwwb/jwT2qsA4r8NPaqRpLd
rOd3O29Ev7kXyijiJtRYBmhBGMdBlqtAl19E96bXFvaGJuPEy899R7o7jO+wcNRUqcytWklm9/4l
TInOXR+cY/G459kFNhFJAIgRL5o7sACcLhoscAHqJvVkW0rp6pftxYSScopcECpEpUWqggFzBawI
uykpYJyhraxTeIXlzKkvty184B5rVCOQtIxJICnjGBTDv4KpuhdtP8eEUJUn/qaFQ7J96KkZhZCE
lsX9LS2RGx2mIX3BLteuli+8f3t+5U1il31kqlxMNHJxAxIvX+rDsg4POjTNEfvLmmV12JASpERX
wjJk8xCSdk9NCqIPFLsgCF6GxkrO/CwZiBZwnEWEIKvMZ9QfK73zi6//lRhep5Q7QG6lGmh19Mlc
tZVq0ujtZU1BVI3Ljje8mJB5njYSAvo1z3jr6dVeSpXkQq23boZGY8+MCEKD36xGoToHvx+uvDNv
qODCLB0I+TDM3KPaV35iPeaR0NvbVK9En++vydvcRqi+A+hz64OWnE1alURqxQbHkibX+uTdhsaf
DCIvaSkl+U/iEWYFvYceGmOZHebE/RQqxhH+lcCem4OEvJgXCWhUfa+ndveyMHtYEIghqSamPAjP
I2D3SzARqJ383k2PzYW7r3g24VHCxeaRDCx2XRVH+nmWJacvUQpwz88z45Si+6kRJMtRAWZ8j+jL
B4X2lvltn7zJWbmCEa55FrpSI+RCzDj+pqDwc2EuH1xHpSwMG+sUMUuCkPZEX4CvdWVIPEbop4Eb
v9ET1rdqO1vBGVf5oKdNYz+2joE2EPo6QWNNS6PPlcLuRHilrj/UHC0m91JwHRUiQKrMvS8HoGrF
iz2Cf0Q/FrDqqoyKyuO0EO5W/Qk5lkpZ1pXpQdnsTz0JxeTFQM24y88I7VLWn/+ieDxDa+eyV/9e
trp20aJ8h4Vtsi7abbUkZ4FbZ7l2FK9UyN+eZwfDQhBUcCNhiSWz0JlmBnuDDw7x2h0YHo+8mnvu
/8tQsxSudqXHbnKZxLg+XR+4n8zD10ouO6TjAG6Tp1GjJyES5j+UR//XV7SQ2Ic1K17mbKfFSe4M
P27tJ6DhNUqmBkRZqyYS2MxwLDVssbBMUxQmcexhHewTv09L83PeJeAdjnpKiuJlDpJZPCQf9K6g
u4uqK+6zabbW7QpC97oJJrmHx7ooMM6vKbdNZ1x1X4LQP+y8nH+8pijXjuEEpT06ME/soT5dSu1r
lnpiMRFL8eT6YK0ppFu8mHJoCZDBjhh5NNSSvJIAs2W8cq7e4W9rrV30RwiP22CVUpElYIV2ff8Z
DkdOdEIQMq/g7QV6Kmr3pWLFhWk3t9MKvEDUVqmiyNQ6wXj6QkRJNyKLm9RTaHL+tlamGVHNiC4C
Q1auv4WrQWBxFYShIYuRF1iTAXlpq+92gCjh99/F3tnlTEYeauBUphTb6n9CCrOX8yyGHPlUItVp
JXzRzRKlqV4y7ZXV4XuLxwLMv9f/6ROS9MRYxXaRtL7ziHUHWac3mpIiOSv6XQe5CIVHPxEIFUvk
0/Jrab2Js/SIT/4vDUvqQK00oMHGX/cTMNz1QLUmDTfymyCQ5cpksAfF0MKANHa6nuwJgjzuAuzT
Vyn0OYrVbb/rX9KXl2yiDiKh0uyABnA5ME22e3NEQGNdjpImjL9XCAiC21zJfMhazltUW1DSoAOK
bCRj9PMyiX5E98+3C1L/FVtnbbNusBG1fUWyE6b/3qN5N2KnBg0YEHZyGzSjrcIBPfD59z24luBg
XuoLLGC+Cq+R2fJKugPQEkkoUpop/I4UX2GWsK0bkEEsgXTIFeH/9U4hebG4tlo4kGCNveeo+HYw
fGWNHVZpI/q1ZE5s9KUCej0XeQdHpr0F53q32y0DXnjvm1M0bN/PEjigYLnVo+d0/un0IvoERcf3
DfNyjjIlZNG1qJeK7DcpTMqooINqAgtIc3Qz9Fs5rHfsY5fGJyQT0IWSD5ynztThpBKjJpwHDZbV
COCf+v6s3RqGZ4DdfBGEyIw+UfyxAI11ZMvmNFixW2YCfypVE5neDbJdZX7yUIRbUMQcRs0Pt9Rc
QCdGjni3sQvnC7kZ4U4jRHN0bB4OLsKhgXlzG0tyXqOx0/MUbq3Z8JrXP/uDyXkEXdpqpbwK2lui
JE7htEN7/R6/dD7TamxLvJRj/t6MNIal3VlokVLpBycRCVvp1aw7fOgJ712gpuYD5FAL17xn0hgv
CAO61NTSFZjMWzdF9C5T6f/EDWd4rH0TWzmcpfRdpesry36+geHawJgHDoZmlJlISgDyH/Snciwg
8HlW5exw32xdJXbuD5adN6hbvBSgg2uVs+HRexFwbmwh/ZE8c/YxMPdJxeCWof7t2OSR/Wwgot3o
6j7mVI066Wt8qBr3aY9GSTLgfs2W6zd6EjGybZurjgRnow5ETyRQEMhlDo0Hu5St3NUk5td/x0Pu
O7dyVJj4e+SvSPn/rWAXoXophOBnaIg0sTtNPt3GCCjoD/5aFOMR4tW9KZbxMGzrRwr42o8oUSeG
j8mGwklyMfhrEdbaBrvrIcMPaJ2+epU0jVuBsY6CQybr75iK+Hqg97fjH0YoQRbVecR4sVNhtire
LI/+uleePxIqgyYR7iRgeK9GTYqf91dT7VGZaoU9q0taTEhm+KGaM7k3C4PCqYxmIAu8zdq7g6pX
frOkVDCP2p1wI9YjbcxBpPhux/3Qzq2O+DdzMd4Rs8bzi+IUb1+BJ8lNHBVon1QwoSDEEWsLx5hU
MGMiDGTH4kYvcj0XoJtvP80yJi947kmDdQVfoyii6WwvqrmVa8nKY+a5zO18rEz3y4VdMwRV1hDt
O8ogkxJRdIpeN1Z2f0hpalJPQHD1I2rnXRLfCEt1XbzxhDTT2NznTisMfgCajWeF1o7o/RQ3NK5K
T8DSV7Z8knd77PPah5ZuNwm1XFRa2CE6r8EdrAjUjX1CfYeY7FgQTJThGbZ+VwADjQZyAEu4OXln
j3+bOI+XvxHAbsSQMWZx8GjflTKp3ebxEyXtjdDaME6tagChM3K3aNhlD6efNJp7M0IEgNGbh4FV
a3lu6j6HwdvEPh1xALAzESRRa96bDzKoK2gL+i8Qk5wEgrNdrorJLf4hIh6CtLUxswRTw/mXtXBP
cn/EMmbvXmXB12HRAciJmjX0Qjd02ul3Xj5zOZeqmYgTIqZV969SZyfk2iZdL2LkfCNgmv1MKmaD
2Ie0gRhZebHrYDt3qeCVDnU5tuBg3LQPt4ta/fJPMG2sVtboty5aZwCBoz0qfaqy6fOnWjwPE9tX
K8BG+VTY9sAlaqVhtsbDqbjhIToQpIJVOW4y8iInDPFkj6SHh59OdSK3YsiFslYlRvUr2DzCHJv8
46/abqySIDv6o+vHXUafq9IX2qCxLfcDp9hhNYVpxwyfvyWZwiciBCo5A4QI99ZNlfjrXoTJGGrX
1dmmtFca8Fg7knFmiHL5LPZSyiE0il/2WjWgLRBLhEGyn2rXZQwG/8E3omlNQ3rEQi8yCWvwP3Hf
xCopNXNLqv6PWgS0Ej/XG0CTwBaPPsDGJRQYPFAKGIxrcWcqC/m2nmlptiCym/q2VLpSk6P3DImB
nWgCIFnr/Bw8nVGVGLWqxt2MSndxceTPEJsv5PhtwPkm+qfzUhWnJxYzgizRtEFFACuakCT7YS+E
Alo5Lbula8z8KKaTQJSdXpjs/LZWuGaANFeYUyvZWKkrYNxY7lR08XS5IoHApYpE/cLNZteyz38m
Y/KDmyUyALdZrpWsxOHJ7c9Jt1Wu1CkGFzuvIR934X/IKlrqm8jjX8qpqHcy+NHwjTpcnlyS4P6K
THFpPMNDORbQ1rApT9uwax9bKqsT4VI9S56cH4z9XX+svM4adtWIppBNrb/DjAn+khLPr/r53dgh
dxfn6epqSDQlH8U6q4HPesWAaTKSjQkGpM+pmj4FKrsKOLrXf43ArNZ/GEMcL/R1DY1z1KBGr1hf
bj24ph+iUqWw7T/fhVb3HrnMtPNiU+kMpCRQ7ZfgsB6SfMM5CbD/BLz/JJu/TSOQM9XlbbCuBCWO
0Mi/SOj7L1kcCkM3kCgxKLB5b29sTq3dGhvKQaMcZii98C1IqFNGki802/tT0lOeJa2lNw9Far3X
0ikHnrOigDdy2SVIne5Arb0+o2uva8T1vB9x5Ql/BNWt/0yf3S0BMZZ6EJGbYW/Dt+6+hZ6jNTVZ
j9cOiIDsEg3MYLvBNCqBFHdnEVv5GsLwqr/eddbaIZzHwpu7N9PyWG++j2MZSy4kzMr7DD2gHOAV
J99CbTlywo7PsIZ7qClES/fXneDpzAzd6Q9IdCTHJEyZ3hcRHrLDaEuq+bybk4khEb9tl7EeGUPU
AI2BbSIX7d1E5iqCSORIjUbSNUbNrLlDxM1neHliCCGbuamZaxCryY5XS1ZDbaLkydeJoHGS2xlg
sBwMILkM/FhuMZ6cPcJ3rgNyfug4IG9I7OZ0ImiucHWY/3VMGFY9xQFCKvcB0K3VI+OYIcGIFvUZ
a+OK+iGTcZx2TVEvOl/IsiYeRvKX+JxEoqYCfG+wNP5pWqTjGPjdpycKzmEUBwfFLIDIM29J198P
ZTCG4jtaM8SxigTWwAZtD+yIo4V8KehLCfdq9nb1yCU/oQLcj9SGEUA5ZxIfjQtrXzVXtQOlWUvp
2zzBhNhck+hEoo7/qO7HD027QBFW2BidGv/mVkqiTCximh9aPg1Oq8XjPjuTbg6GrGkGT4LbW1Np
bkZCRp59Z8qX6NZ8b7sNvQbquPgLn47Fbp96kvwcwuIMSGA1aYSRkBQOUAAJHg/3T8IU/9Ou9RQ3
A3ytdPQXotEj9rIzzsKU6iwWVu/M1tQ9muL5crcv0riObs3s4SSJe4KoseejCE4EHP/x5pgXn1uW
H6NI+jPaHq97EzRsVvuzl8yK+Hi7uBNhOBPNWzxSqgFBiOhEiaD8IoFLkJBVryUZy7F77g8q4Onn
DcTwqVjP1agN35sRHd7+Hqj8gP2WXhDI1VQcYeB0kz8q2nx14MPFbH4Nh6ZE82uECwVN4DtdhwdA
+FNrZ4p6QH32T370n6FM1dQm6nysTWE/rtxSN6+Ap8vSlbZkHBHoo5L3AYyfEkgwjM0C0lRkma4+
M+Mnib+H1TG5q74CLTZy0SfUyLjRvCTcRDObOBoraIEyoRaLbRSQfLlW7cv5RpKieiPjENeOlEsR
vDbq9lqxCwDj0Ufq5setejXzw9oAUgbjl2B4xhcFRhX/TohfxrbkNbnrUq76ISEzjnueE2p4TcFv
2hy6Xl++QErOiV266p1RohM0cEQofzc3GO09GR4+wD3QdnqWtkbI9kG+HAT2yy8onTkhu3QIPULD
sq8jSJ9M40o2wYyIxgeXDvpgPabfZfJyYu0LGvrVc5q1Q7TT3D8pETA40gzSU1WfJi/Jex302/kv
KJJ07ekxMuQASO4JwmF12kLE2Tu1E3mzrM6BJaEyZFZncYvINgy933jhFvdBIbynrVDxXfM0Jq6a
hIj2UfP5LViYsNbLRqpou8H3g4Cc5YWRIuYL5FoaZQXBP5mkRyQcHE1OCdvnncnNEm3h0v7MkfUR
vDrN8gym0WISEIEWntmoVz9O5D/TCqZgb+E8GowWl5BjhoIsnHYSTe0RroYp0Qt8ck3MJl3/5gme
OfhG/hnf/eC6F+5bpR34e7F+2FPOjHg+CTw/ju+1bV3obLTNbdLgmXx5wq7vA2BmMR8N5qcSU1Py
33wY0T0RmgxygrUP1D5BbiRJf4UzRwsYC/wX9oC6bSesN3PEOOR76DfctDj1hMh51pKVQBcxjsVn
b96Khmxsl1/0BmXeMxYT9NxbRnJQdN9VcYTxXXCt8xe+Qdm2q3bNXSR67oq0rpk8Ff+pRiI49OEI
ydaSOKPh0wjqYNCYo3iR0736KroZAQrx0htJ5SEsAmow7tZfJNPYACltDXj2HEr69yhUv7U7FE5L
+Nqv57qp9epIyN4UUEH6AocMc4y1hly1GgM4cf4qrmX4PtpM41crjPYJmbzQH/SY20HxKmiYmS0D
U7aJcJ7WMVL+SeGwXQK0z2CsMuZo8aY5MeYWjTryF+zAI8J+VYJ7HB2vBUtbONWQLJz87siZ4M+6
Dk/OmvP+5UOvUMxbT3TGGpkXrUyQhJEUDK9gqrrQcBPPAEG9l8cRb7m0GXDlVvqdduXoj4bUJf0Y
2rToxyeKI+/HQE4wZKZVl+LMZLO6zs63DMXGO4n1FoGC0jG65DqlRnOquML5aF6TT9kxd814P5I7
29SMT26yu02Ddd9LpEigrlXLchzOhoyBl2bejVq07ULfgW1CZRNf873VdgoN4Jk3QkRoR3C/Wfet
yfITvtTbFGnWN0i/Va2BhHGCXLDJuvuS+q5P6Qulx7eLR7JoUgp67ADBS0CDkmTD4lxAxWpfcZz5
Z6kmUREL3BiQCmvvu+RabvtK0Ri88ymnqgQv/5w4xWymNouqI+pGl/6MNcdiBbFDcVnbPMCGGxDN
sHF911BZPy+kkgxOTmHQg2WUnOFM9fS+R2E26w9FgxkvBBKOixB6kUgzElzUHogHMaXa3NILSyHr
IBhI65UCGhTrLRuPN/tn4FjeECcF9lAmUW4A0rFlzOi6qwhyeOoMJ/zmX5iFuTiWnyQm21oMVt2S
pGVBH1fDbSzSi+fCWRP3lo7opOCGNQWqWZbKDHx8JizHe3riORhAjOuC+fRlK1SM8h83qtimHUVT
HKs3Me3wfxUtwl+L7kUKHKmGNjd7ys2OiWr3FfUJRkMyAhT18yFqW9nG9+knO006nKCDGPJOXul/
bqwwABom79OJDSjnFNLJPjpjwe7/TChK+rC2jWQW4evKEm48TnGVziSxjY+etGOlSdjy2XaXEMce
+M9jEVTvIZk5S3/12TH18i2GSBk52L7amZeQ1aUn/tENLknutl7hPswAUq8CTmHQFrjk8lH7yrbY
UPSuBDjYJJdIZvhsaykMgGFR7HsSkogT/bxrMwU7872jM1E7qGn8LLffsc8KGgK4k4cjnpOWMq57
jqFlJW8PvwJeA2OCrqD2iO8MXcxFUA3mToGT0dQR45YZudQt5WwJw5FbcUihWOqfFo/XEKOTxaf1
om602+K0rwkqRWeYsmG5znrYBHvZHPTs92b5yNlD7SFiag7Nt6xPkGry0vz/kEEWRuwdMCBTCt0e
E14nd1+NAh6iVEHwmx0O8bhYi0iH5/mAhphO2W4KqWsXFA00t/uGwlNbwKRAiDy1qk+hIajNSzwN
CVxF6vp62heFYPhTWzzlgazT8yasK2qDophJmybbD+vG2UINhh9EUw2rJEYcQk9enfapB4lGXr4B
OL0pgVXocPn/Uqj0tp7+mf0QCdZJ/HEUUJX526lJvUWTepUjDdp9MASdCwcqfsaDlyDk/Jqci57b
47sL1sF2WzAWPvx+6NvWbIiJ56CQCHo/biaQ71/Dw+q1T82yVbDRqQvDmjsx9WD0IOUa1xoHvMsq
3WzIrYgB8g3bkuQp6f/wlBdw1cNOGuXiDjOvQTugC/jO9LohoJRcx9s6+a7bfXQ+amD/Yg3BbHHo
cSrqsdxylzqA9Zi0kzO77tyocghgcqFSlW6AcTNFmdS88i7vZBR/Rf2k/yda8vcw4khkN6ZY8mL7
BbMyFlBRugLc4Wr2oIzr55u+MBsLB9cHoeETe/hCVBnrtv3bU9I0vYV4PCdWVbK2KFT+mD1+swCU
U1bPgSVwKxRBmAhGxyN48sHbsJJr/nQSob/3P2AOrmPYf4sTPZcfCG5THTvjNCYR+JMORKTAJmmR
tcfui4gPb5mIMLPHiwdF7+qzfoMy88mQBP/I08spnoIaB/0XEGbJGjxGcadoirEEQBIufrdU1DFd
UcubqMX6UdaRKmcwPYaTqcIiTT7nTbkk+XsxVu+zz/9m6NhNPTcbMzlXuZ67ZGnx5rE0JNPPXMTR
fCAk5Lz6Vxn/UgT5YraiIYEJDuwiYQrGTeuPoJlJj60N5NJoqHx/PoRICvcIQ5DZo3hUXeK3ylta
V8WC88kn6hnJ/snu0sjivTgxZicQVfcwNTKbcdWQFRGYDoV2KOjh2i6cobIDBL9Bz9fr2yx2JVmK
RoihpqCxUEgL4c0cvmGLkVLo85vjlP24LqJ5+H30MDEoIKO8sBPt+CbreMI3hE5xMB9hDxzhNN76
kE8iHaTNt1/UUHao6a2n/nNStNtARNne1bjjvuEZkderQkVLu009dL+D+t0BvA5V3Ak6bkLfxXoR
kR6UzC+75SFbwzqzG3tzm6qo89accQiOyFVW0FlGhYLkMt6fMm9LEg7uEHqRxLcfX8i0xfCi9xwx
CdKx3C+vS9Z+QB+eEMNkvtzKk8fSAw3E0ssoqwfMmzEOnMd0VsKVfIvHVvr2Qi0eSdEgTIIK5SOP
tp9JSeILStjgqO/YgtKyH4bjw5WIh0PY/QBlDuj4jqtuuHBT4UVHZ3C+bH17CbW8rZ6/dDax0sQV
OZcmrIi9FlYCKPKu868HKNMEUjOInOBLD2ZIEZ5is3eHS+ABqL84BFoa6qsZLMSFlLitCejprf2L
5M89baDY5Z3Xrv8Nso0exgM1fpLxo+ASAbRqxx2FFtq32sV0OzPAMR6rw5TaFbCTdq21yNL17i+y
SIfznFQwmB55nK0c+KcW9ryVOATI9hCmNMSckYwuRFegk5ySGVMB2JXlFqMUrlhYNJmLbm1r/y5A
YYak2FMR7syyyCTb/dKh1BiEdZsvHYMGRweh/8o3wMSaghsdJ18RA9dPtIEOxo0oKO7IXDjwlyhw
BwEsGWkjp3mW0darp09pqPbAFo0HKk+bOslYSII2db+nu/ZpHrQPbqfHG7R4gdLa3d8jxeDdO90N
etx6zDdpAub7W4FFygns3fnLlrUvPOeEvmpNM3+LAhIesJ/q8QJOlICzGinW+UOc2kxN7WGp5ESG
cSvMuK7J5uGJgAnIzxa9hmGiq+ynFQ9d8RfXF8X33g2ICcQF25UYJ/QLtvuOyh8g3Cr6QvJhkbBy
6i/Hv8/WOt6L+Bc6IN4Artr0qExm4ryAS7Em0k92kavSEz3qnY7faPOHpZYJnXngxUOv88fqQfnp
A3WufbLOfddebqA0glvvMLgEJGH+c/GrSMzM6RXpUZuaBszjCrTo6Jd0KUR41VD2buAKm9TR/bJh
AUrLgjnA+UrdfE8v/ufcIVHdoys9y9UEcT7p70t8onFMN0AuukPAl2RtYycJq4pI50QxGYRsaeUQ
i6Sxfkz3auH4L+dPIisFu2/OLsL5Bi4Wu+XdjaD1kGuI8sKZq311yUaAkpjpHVZzuWKjHZn9DE8d
4UdD4SWnFpl9JiIyTgGN9d9F9w3Cz8WjR1zPK6Z6U76ecuKO5cFIM9ORWGoCeboIFt1e1aMGYZZE
Y77jlLb8fSx2pP9IZ/JldCwh0oNgOws4p0a5zgL5YMnIkL+HGGdz45Jd7zO96zYunNaBDUNB6PMX
ZhAD+2fDpkEj4k1LXQD7SaeSWmn2npkBei75gkFJkPzMAZFwmcTlvvQFrES90gJEgdnmiVkwfMIb
Lb1oiA4ADPMlF7PYr/aXMGmekQvDFgWzHsDKvsMkB/uoI34HH2l2Kl6SaRYVWI/SM/3ESpcPgCrQ
A52qwYn2duJgqIdDH93yR3RClnQtxyGpK9dzBq2f0TN2Fp+IRI5TOJYYpvsu646r+tYQxAAiVgAo
mzfUANs9lq8ckaoSNWWbuFWk4JisSJIRe4kAEPy5hOkDMlhxLx2AbYX5AuR/ms5o+znN8GTUwQBs
v55KWVoOIXErZ0qzsfdrOomhvIFoWvWJQsiv/IwiCEsDhvrFAeLaz1jPR/M7BBMQ7d1jRWGbAYsE
qGyDC7AIZgOljKs7Nox3Bae4weP7p91R1ZcROmpsGURsnKBUOWLWcizyrYrwR1s983wMLxcj/AW/
p3CmeWGZEFkGuvyoS4rti0qgSHN4d9r3wMRIaGmRy+853dWoL9LKpMCLv53OlD1nAp7UhFf7lutg
W8Xz5DxbbHSxvLIzFoPilsWe4UxGlQdS3g3s5SJLkyP0rIby+dwMNXrFZz1kxh8IRRrjE6gfevT5
ozER+BWRypF1b2iUDtcqdKH6ShiKlfG5lV0iS9iu02KX3XlsNYia+uTcjhWWNolAcjlampV/NK3y
O3ZhvybPI1/aGBUCHZemkvFWAW2sFgq5STW3TmTK1xp0wbuBGHB5Kkex82KxUhM6tm9g2/ss01pW
DY3NkkcLLi1iyAA69budiV3A2qxdjuyMozifFLmPWfvciUINbls7PcedN/aa7+/TD8L1Iyz4fZZT
bcuhc51Mrk7/sBq7lOHTZ/xXNKPt74ZB7u9iDgSFhgnQI1/7YQFcJ5bpTg776yVA2Fgofhb1ekPI
7l3nC3FoMk3bVUQFVcNHj42bn/wdgOd2xX5Bx5bNQA4IRTsbbkNb1pVEI7hEgjvamo/GBQMSNMGJ
oWuRf5vgbcOfSsE9ImKmxkFg/7+rt2cxZ4WcmSLbKmG1bZExEyOKYgxt6S5Ms+d9LLOMmzDfGf0p
IBvsLBBm072pZNEosHJ0kKfro724oxgT7RuR9NDg8ettbC6Gm6LmEh4PjgGIy7gXiZMMklFVOmdt
r9kGDXuho0uYIN1xHLAp84HTXjoaEBqbMRd9dVFZgOBmRgVAbjNhafOQRiSAyYmP8stFKsw/YpIE
mGyDYoUATYrb5OH5h32A4weRJduTAze4kEEae5p8XZhBF0dOTQa8b1tcbJJKz7u40qUkKk+FBVjD
siKO9R8HAVd6T7d/+vQ+xer7gSEsIRbqS+BKr3pj6pfzYkhgzTK0d+LDfENzFJOU6tD3mGJrcbP5
wiKpSi8CRrRf5Dshq9uzS2H99DBt7FhDp5vHtydMbJt5JGq19OArdYM8hKEZwMFXHhA6hmIV2QRR
IvIKQMZmnWqsaC5H+HgnSMgAEK5MMiGtSXlCaXD5yRalS4S7oBaj1DMOrD+HXAA4nG1uYirfNN+4
di4s1F/uR00CuYfT4zigORZrUS+OExwlgt2qFYH9jeWOCaEy35E+RilFQFhaI88LeicPb2c/TT4U
/i/Xog7l6p+jHbCQTVFALIZF5cpEuY9VfOlFYI5oIviuhfl6ccN7Jomns23P+vrU2S5GVe1CDRG8
hHNHzCvmM5KQTyqjix4MZyqQMiRiLXG8DcmlmPR40uN/Qgfk6u87U+Gw5+Ce26Afs5DbswDc8QUl
aUMX/oVp1eWKTpEc2NzXmluG+YlfapA2GNbOdl76lejcgEEUFFzjlxHyu3s4izGseeTfbr4cZAyw
tmaFde8MemfdpUJ+no2dPamXJS0hp+vHAri0TJ0e5Hna3sMnZKgCr6HbQeOdTrxfTY+d5rZG8p+w
iaAF+BVXXSc1a91KLAjI7isemZ25aO0278GeKt0i0roTS01Jego8+geIuto7vu/TQcOrIfrDxEZA
70ayPPm8+IuL+/ewcN+ppffugkrf7dNOn0ymR6JzcNuzIRx1ciW0plmVY9k529IZVFg2ArysbbYQ
qaa/6dKP8R8tH+3QkwgpjNfgMcVtin4a3Ze/fdbwi8xML0ANnPom8Om6WoLuunE4ppov+BW2R+TD
WbJAKvWpf6uLuNf9zgDPvlF5i9tcxijMoD4MvvVIFACcr1t0N/beTM0exNSNcRjZgBZOsGeP+7Fc
ajDOPgSNbEF91oAIRhVuVVrTRAD4OsRZax2Cq4DyofkxfVdiLsX92PHQD8ekmM2RrgoOmQ++gz5Y
j8I0LJxwqs9co5Kuudeqpdq2BfFIbBNPrLScSSSc2zIBDHY1EtIUQtZXF35WwrN9rVkFOiBxdbrk
Pe4lbRXlib++1X0qcrMNIu226kcXIQyLX42KaJ8GmSz2+FTol+iAbRiuu6nuzcWyvLSkB540hlTF
zbOKgeLzt8sa9YVnJNf3TUDd/VwAfqVNFrzVL2ziRgv4D0XMEiwaXrlOl7aN0AdJUxWwATUQIJxW
dujGbFAMnunMOr2aili/+FqySNLnZlYVaaWTuigDPLh46Y2vtq/rCJjy+w1x/EMpL3g9BrM7LVeX
88rWndWRGLiiri3BZrw7sZQlaYLoAHXXpnBFHpbomYXPEKCY/Sa4FwqwIepSwJwIN15lcGXzD5gA
M0l/xAk7v3rVdcHYbrfj8J0ldLqidp96/sdnNz22ToGbfPyH3cdVTAJWqrDyoS4kQr81cgQOj3Mg
iXAeSZBrtfzFjTUH0D2ap9a9uTpSJSQh4qjiCJcOuefKhph1PWeEE3IzrOSlFpI6uuNmnPSyhUin
kdEBvIpbd2PYNbocN/J4FpCpx2GUvuc/hdpbpO10eS+KJGMVSF2UDM2UFcrKvU1g5F32IaNV3ciD
aLAhl2/nmBAb1dqn5rj9a6eQFla8NwsnUDeigFcAlt4cNIkpw/xWXUTHUHcyZcXYcKIj8BJO30p0
2D8GVn2GV0P7KThAf86BZuJluTIdmnqIykuy3i7mQYPhMJgC1lznCHt+XwFAMFQ17MGvbimSuoC7
ydz/Bi3kE0HzHfmxRi1Skqgc5PypNX20H/N3MMOZzL5qEBqWMBgS5YT1djoyejuLarS62qYCm9Jq
UnfDjp+4+3INsKEoenO+FLtl9S2OgI1jfQxPQvrzmvLV5EYSHW7SY6QwHAVaKs7iVjOLe6TBTy0A
hpn9m3KhQK6BC/LX8WvhvP0cVlAmqZmakqxcHp2U2TWbUssadOZnKyjV+KN62LbWorLZBYSb/ZU7
e54WqbZnyWdAg0sm4GIlqw31KUvqxnnhEi9BSXP5xU20jQynebkpuSrZl7WAUlJH3b23feF6e2Ka
vVcHEbeb+81xhIq4E7/sqLAboKYuPyYxtldbjWxpONELMXmbMVmCWHCi+O8VqBZEykOjX0iz/0w4
GkX4WH44bAKY4PDXW6vRRoHnKuuUXDPKmVd7bdqF5VymeSDOWaJAZrBqqpBuaQ55prNJXUh4y59b
/nLAcSxmJp7c7T+WiORrgHLGdLpf5z+/UaSYwRCUhBFp5HP4UOKPQGAlSFR8BkbawJYt8UT2mV28
fvgJmNy/kvekVTgksuxddR/7SMtImfVorWtnqcVv/8L8OLGHp8eXWR5T033Mim6j5reusuoRfDre
KaPEAR9hHNT4TY/SGJsby4eeRmS/4NggmGkOqD9xuSRfH6i/nPqlzwzxCHMQBZR/MfvUm6jN1Kw+
J1KTu+0gZe4+VXX0xwTAm9xTuDqwCIidDBMFIrkc2Y250w1XbjxNU3OvE0wiWLntaG+eB/eFtnbO
UgF7k+AowPxi4izFi+tZ8JPtoTX2AzvcUYEaIreF9pgNOuT0c8YwfG1hll6RGU7M4NAUrQoWe+5s
BzRGNjjSryssLR5Y2KCo2EUJBSSVaTq82Wlmn/EiDZs4naq5eOVPu5XOHSAqaSIjJBgPHnkidO3K
zGeHX6X8ZE9R4Wev36sLA0CBE41UEvcCs2Rqp8UPe8BFIuHRyAU/GAzvB8/NjQBFkGvXC4t3Z4ua
xpi6q29/HfFiP/JTaIZHv0OmzWDQ3EcQHIVeQB+w+gu7HrFHArz4EkVS/hJLiPToiFkSwtdotE4V
KctcbobVBAy3ObCFOuwOlm7VzNpHVd44+q8C6AkJ0CR8KovnrF1JadmyTkaYqhGttTrq/DVK0Y6R
qD3zHYGAYyCocvlAK1amX8fUZbEKo2rqYmgycuS/CuP670fx2F9Apg5GPOXkIIPVCS5N8g4NH3EX
j0DHG0SuwM5+W3W6iAJFDxSaD7lhlEroeU9hqkXpjN7tK0TPWbKROXz8TSFVRgNtxXjONqYSmaey
ytLEQ79fy62e0w8su91kDkBxx+QbKGRTW+0jKKS+O87AsCnk9zNgW23pGbMz9zqhNzrVhlFLOW20
e3x4kGSUb1wCxX02gVW2mHBrYGk5A7CMlqSI0UDRIK1dcFKQ2u+Wd3u1Mqs1E3Ju1yno73ar4DRk
MNPa1kXlAI9ssxP8uxY79Y+XD5GcbgBImH0wpWw0XD9Mpe6paArOHHw6pynR99uIVYY5ywHUrMHo
SvNwunAgVIi971/r+dpyz8Mn9Rxx6KYnwQ8YuLqMqmXiT1nTFTmSZKE8p9+fyr3j4EjqHPu6MF4J
TcwXxxsVaAO2QQJm3FLUxCuho5oa+oc8xFgudKWuH5XGrqtCGE1tcCV2p66Dkpw4RzSQbgUMXyKX
yD2ClGvAg8lz7iNODzVxSijz+6az9vXkTlQ/L2bppk9IqjojQaUzaxtMoDbIXQVfO390qkvZozvd
oxIpSK14Y1nJU79DAr+GtQskxbFBMKydDS+vs9jmTDHVGIGlAu0TCuMrxeoLDcNbLb2ALrkZP1Uo
xVesMvo3/gsDYHTAlvG6tRK6zASxTUtXra58JvgN9xe+IsW/5tL9GrJKipg6Sco7NicPTlnpYpn9
8R7OSMmfie3Ao0HK6A1k7UsaaXrYDC7Onv+6I7zXxXavnIo2Yb/p3tEZ0zWmo/MjSxEp/+jS73fs
YN2+ZlrjmlPMyAtrJdmyGFSTzcSlllLKfBGCDY3X5WE6oBddSxIjUZAMPBjnfljUF7RIIXO3mAND
jKRJk8J/KGFeP9okehh0UcQcNr4Yl5p+YhtUso3XMh9ngTpzhaJbQ8JapGhlINaSGz9BZ1/MlyKr
8Dz3UJR6EcjohYTJIE8pUkVM0kO8lPNT3QL1CkgLR6vMCddF8wyW2YFY1Bn+JDFM9MNj3AjeK562
TZu7nLbGg/dEu5ZH2NjNM42JsHawI/Jrg6F3b37Yd4XzkPmv+VYdUOM/KeCxbrZUUwPzWcl/Kuz7
mAzLLM3mB638/T5wcbfVIqO82FhgRfJyLcRQpOEZyV0AEcy/QsSTQyxkcttH4jf9hMkTm16Qy3sK
1ERfEtLUYxJMyWIYv3iy2lsMZlb1X4ygqAYXSemk5yAlw3JHMLeNt2w67EeTKAlnVhSoqwCgByP6
s1QEbwkgUNRdNhMaBMU+VwjdBHgDGRKfJGVcxLniggPUDULmv/Q61KJsVSm15vrFgbPz57IxBav2
1Tvay3JfzbZfV5IpwmnD8X6834WnF5noI/apIGTvvOT6tDtYCkx5DpdmZvJhLcSY1LZMIzdLzhZf
2ej7yhgM6bXfKaB2HLLuVYzoiSzGjYGtKOr0spssONZJPAYJGuuoxxvQ4ZyUScXUvxzJFrLgZxes
RxGKD6ST6EpS5gu0kdxlGXKGQs3rZtKbytG6UQCzax59WWeFjrRIl2iXDRo0jNMIkh9vI8P81gqC
vaBmXbasmAeaRvoPRJMGRS0OmyfYDjO/HHkjzCTjMLkQ/4i7dYzhKzjfNno1rmmjZbBz11EWaOp1
aJ4cgyvGcvoYBeUwaHF26zK9Lzgp7ypVXu3Kq5hyOUOPPXKlOaDgwMn3AAYXJBazUjDdNxPu/ybm
YbhOP8OYi8ZGE5xixjJ3WizJyIGZOkyVQgsEu4IZErbp+oSazvAr//AAQqMYEH0i4n9xImoSZ9gP
F2mWc3bNaFXcqijm2nvwAPK8CUX6jsVybjGbs7xWroi0ahp2tRXBGjIbFA2JZNj+vyZ8dn2iqANQ
YDS+HKsB81lxvKjSdc9oIyhX30H2jnmPuzWMMYGDyBxc0mjqMFZWz9izC8jhzb0XTplMAeMrxsmR
+c/i8yCS2NHsaf7yF5ER9Qh367VO9XNL8H5dOh0C73oW3cmfOTaYW/PFflbkCbkbAaKOnIrjBUmi
j7ClFmKICXqHn24QpL27LezXkqt3rklaHSUMS8bZDN9bGXHeHztD8ypX+wC8AGnP7ZZUkJ8LjBmF
adbaDJYmeds33e5nPPKKTz0aI7CK+bhwNHicld0la4VSC3aRNgyt06POk2fz/X59SmNTVIyM7RKs
FGkzEbaB0fRG814Hf/U2moh6AZl1hxP9GNwHIlur7Rh7ai7ZNmozA/JHXqmEp1Q9R4dzS71WLcLH
sD98mcc5dYzZDp7wEYrYr/hEcU1VQ+y51s0uWOtCj2T6KFkr2MYr0wbyjjFnCS8FPutNZLDn9+MB
sFKpjMb1if9zMwy6DpLhT1a7ODLg7yba8oScfO8DceBuvZI3igEQxVLtYygDM1kHRNJwGSn/9k1F
OnPRTZcjkrroPZhMvQ6fHohTGilYmjBisUQXfDrpYwV1KnW4bOtvBiDlqdUjzjdTeAFdQgFYAj1Q
8a3epQqZQg9Gc00RG5HkeBZH2UkUEWWUwhpUxwTtz7520dbbd/D25VgRGgplw8mcUykHwGNf6F6e
2alAjG/u1Ui48C0QGlR2UJmzNepClZM9gCyr42WwsyqGdk2ApoDdP5nVNrNxsDHV3lWNoSA0dAhT
qrS09W2lcdIprDWHQfaAQ+cYrI4lAcB8no89xq7L5obAWnAybFljRzITbBxkc9qc35V0do4Q01MS
QcnbsoVwjzpgP6FLWZ3w3oob+bkCoVtLmUUBEZbUWx4namEDE3fHV9unJGAqwMNRsiN77Lirz8fy
yIzcvfLFL7CdJ5qi0uz7fcVImGQOFHJXz/+lrebsQtndBM58LLPaZScMsc2+m0cHH7GN+q0AAJvF
qL5cPKkHfwJJA6+cma5I/ZDeUohSxS9I57HhoUbuxtTGXNLCExLVeHfKkbPbiBdnICYiJoYnjD7M
MGYKAigutIQvL+jEvIc/C73xa+6jLLfxm3N1scUxJf26Yx49E+gajaPaPG9mkkN4nwh3mac/uRgq
1XDNUXoPM+ihOevIRW7lpZkkSgsYge11jtrpwQUw/46CFa4Ptc4xkT2AnzY4uWRQVdW4lUdPue3a
cp2ooZNdCrvLO8y2JRAxsm9Bl3PlUuBxz5ps6kbmXOq2avyz0pEG6AjMIer4snS+9ZaytS69IF/G
dnN7ntrLfz23H1ZXX+jHJok0tjx1vmMOsdQXLHyMJNlaCum/TN+gffRtj86JtbaqMObhDO4GO8Ev
xen5PRNQCJEwL2/y0gKiETaZ93ien/M4Pt4MwqkKmcGRifx+pGaW1JOPwHQU9nSy1Bgvnvofzzy+
2G6UFFUUd9Jz0hpM9C0ycdmyWc7EKvQA/2q5pipuJrOmhJ4GzqD9yq0+shq6XQedUZkcE2RxC9eq
6CLo8zDqLx0rQaLXukQ6mDtAagaXZI55ufvmaDjImLn0ijHgPprBHG4dYdCDHi2wGnl+lKfndSda
XTRQammJYLoFAE2lmO9jF5e3sR0NCH5m4vhorE3Q+/Rkl3pDHBCX/kOlyomOQlniBSfsUkqLK8ZE
1W7eEpXlEs6vKQiE7mX04fodaJN9zfYenuLuOgvBlC/06pZLDFtOHiRnINI8waO4Y4nwwUHnAuFV
Ae/GY/ZTHdV8p1AJn0NGCS9qgllEZ0WDJprBu6QPeUpr24Gf5ovFZX+nLhl1ZRf/1fKI8+TJtkea
4wQZ/3bxlb/ks268ULeFb2qmt+f5k4dNj5Yjicwx2QOcaALJCp+ktIFZWgnpQpRVWmL+xeq/gim8
kMWY+tqQFT4bLY3bkvbQs5Bs/Uh9hfPM5WsiaPIv47cDJ2GGzEwerhJ7Mg7V/fMLK0KEHkk4flBv
rcJNfi/2CFU+yuRUo8WNEazgCw5muR24xKIf+Le1nE/T8YNlyS+tkYhjRDE2iEHRppI6kMt0BvM0
42Qc3ZzDcfWE4JE8TiWGpp2mOX8gzqh9ykUFV0koNcGEsxFZLl4nj47I+tl8C6tfIWp4diRXqywf
fUYT5vutK/LbJNSEKOonqvx3B+m7qo4lqri8L8EUVEwkc6p5NUsMoZCGpyAML0Jbq8zQ6754FPPi
WukxLnxAefy5h06klldWDDetGu4WSthvtUtjV+9WrrwcuC2xYGOHg93TQcnyg53N8JhEhYG1X1z5
lTanXQAI6VGeiB07RSQjfaqcuTEL/YjlY9x5gYagQHqr3cS3YVlve+RUKjqHe0FyxQpAPTzHexDp
nd3CY4KPTjg1alNvBoEvYbOYawAN7LXNc7mi7kfAiaBT1/5hzUndI7O48ngOxiIWSPfY9U4TY4KA
us/DtdE1JnnmF308/dkCCNAhIqm8pDLCOaGEmnFoPVeZrOZhhCCQqCAbbP6kBvAMO8WhgoUEs6ze
ZI6DM0UHUzU6w6xykmX+9T6Oi5KVOEjK16Qpbh80co/LcmYFBCLqDhl1MN49x4605tzUWYZW0AGj
alzaAayMODWPMjbiEu/WyjSB5gOA3R0OuDhckAFv+QQf+X/cw7KvyGUrLQ8Q8sl324nGEMOeGHaj
vMp45GUz8FcT1vWcvowsZ3x8xV+ZBvjniojfngnWWPhaAuef3r+WfcII7y9MVrHDgeTpPiD3ZfZv
P5u8DOyxNyWzKb2evpSX8D0M4YeGLAMa3oYzYawVfiu5ANtNWMaT+3ZSnr6dKv0CLz9mrSLXgQo5
Wba7mHVTJl1pPgEZ7NHij21kEawp1ATftUqYOBXvXv2WQJJ78MoO1uGUrfa9PQy5/J1OsXK7PzJq
F6lLN63ENXIrrdRjCKRIzi1rNOu9InpNwN/9lYkV0SK2ZmIx7yUdtrabEuWbZRmbl0ju/NC0OD2P
SEDBAOtsrqwb/eC70g2BXURNgESEwOL0chbi1l8GfjyHib0KSnQ5u6CvVEmUJv1wMnRI+zeJX1Rl
tF8BicXcs0TaPBmJqgjMdhvvVy0Nf7KjKbKVQzGWiibTHbenBAjxZ9PzcMfRTXb7N7zcMuuJxbta
AwyxfY1FGUxlIEZUcwFnNvAJn8EHrvDWRU7BTOzMdCHQaZyTWleHLI4/Xn4wehiYTOIL7QIEmxTi
VuhjfL1y+epLXV4DJFgn2fzPBbXF/eLof/1SBcE2ahxgPnmux0G1FZeXVDbw0FdA1mzT5q9fr/Qv
cz7Tf+ub0DnkcamctrUkJwe5UxuwnxevndjLsU/X/qVnt9J22IZu+DyALuWcwuHM//IF7UGHPrzn
JfFOvxkoE8GIe6h+MuWkzu+Ypdxbqu4ddP4gua1hp1al/mZ81wf2hWWjaovOablcxVel9EA85AlN
cj2VTU+jenBWc1fGqdJjdDUwlRLPQtr9meYWjNA9j7aRv9n1eC06X4e+8xLBPUNxcWe4e1EjE8di
DwdmwzEeAyj/OLOCFiMgR9TTxXXYbIVNvv4GFgLagfhbIOuo4eol0beVrRAYIS4I/wxEQG4X8f+i
O+fThv3+i4+n/ffqlIcNRa33NLv/Kn3rsMQHMxDTNTBfWcQJHArZYA5jovfJjFAQ1quPTyrxa8Io
X+G73GxPTj0nMzwbdNVT2wxuIlmZPm7rhaasYUMttiuhwfz8TVBT3Q5UDSwOQ8VGKeKtHl+9LhiY
D/yYo2gytpQvKFKWT1CXgbD0i6kNbZIlZddCSJNJ8LrASOo6XrtqzrN6bEIUEjCU6oRJ1ynZl1zB
2gRjMR8g8C/lN7J5QBEn8ypXMyYIEOO6kosCOctRZV/wJPNQ2F+/n4vcGZxeZTsvCVDySvN2OcbV
dl5CdDEoN25ti+dvfZLqQFDYSwXu0dZc9bTQbzkZ4wmHkGru66/1VFukiUj7QtsuY4nC5KFf0ApP
9zj6aTttKV5uarvKAMAlfZUa4lkHYD4LCaWNgHqt1uWNM0vt21EK3bq3Qct6uazN7b8POXlPR0Rn
TH14tD8r3sAt+hV7dm2L0aDhuvtm5XczpzW31lwMjBMQxqUqE/7p7BVkT1WTIK2PdETdMzXB7Gd5
ijm5IGhQTuP1rMg6NbaxA6mw7fzbcpN5fw0XH6bLD+/P+XmrbuApbtdwyjQwqUZTblcAeQrzrVmx
1JXRCwv5lq1IoqnF3sTf3bwzDROvyH2JRzrorEda/spuxRya0wP7fdZ3aOz7TW6JD21WXs7i2bdA
/WhtGb2MfJpcIFa8E4t4zOQjHBWWgYF7Rnqyr2cO6TRg4pP/gzuHL6kZcQjvf9DFpOUYRlJsQjp/
qs8rRtM9f6AS62W3BUzwo84xHIUVnwV/lOW2xgLHoEhCGvHT7Q/T4zq2GUHwohMrNMIKOnGXDxjJ
b/w6M8sxaheYTLFa9oJGdysB16H1JmPyRdwJd8+7O0FWofaqMgVVDcYEZ3o2q6Mh5NYYVMLzesV9
mDqau3MPlBFkIQ7VLeOl0TuIuLFFQ3wOrh9tcArDNC0+Av5KLuzb9hei5+Qk0Gxpd93/ev9eGYfD
LZz3NildCqfhkKfRuNh0WHgUNS1qoXkXxacuRmMvNGObBwlnW02ieopgroSyh5iMzAQxJqgszBAZ
7e0H4Ud2CtN1TC5XoCJl63vu+rUciXPS8vLHcY8LyoRHoltmK5NqQivjQuL+C+/37XMV/DWmZdeT
o3BHwI+FSuwF4yb+65P4toQ7Vl8+Xw/jj5GoW1igOlNRnvZ79mxlAB4n4e5OSCIinUHBHc9furyB
s2hyq+rqeERJpMZuhW/iBaSR5J9htIa0FEcWdwQTn+rt3Di9jrhjBwRGFMyIzXHhSEw3URmg+p9N
w/BTVgBvI9sggAFhV75uJvKyk6pDa4NBBcR4x8u3KU0IYhk7zw5tmmfzBnBj+9OGMWPLHwTkRdWU
HFSugIZ80hiL2csUPTSxgBZdTW+m9dAlPqmchiCShhEZwzOCZ3WDyndwzFVZdpQIDRvIaRXPKzjD
DjYMbvpKn4k8YTKma3WzeMp4eBVOw4CcsmKkmVV6KOfI78KNz9++ZUc7GwvCj1OdrUj36lPoxYfP
3jaeBW934roOx41mlAs+vdQ6Y9zx3Ji88+GJ3Rp4zxtNqbe2tBCFc5OCTwHBjm2sVoDEIMUx3tvq
/HHyYhEISrkA5FA+zG3gsN3S+fbikNsZrS6MDTD5K9+VTkNquEE957w+SMwFMjLbpA3B9SXKBjKu
URvqlTQux/DeLqbuSLIw9cI88igX4dSbJQtd3Y73aM+IgDXeqLPPvIrwrmTD/mKuQZe4L3E/TSzh
0RDjUymGtzKK6GkX9H2u979J9wQC2XuqsJKWIJxPrHoV0Bn/ilZHo9GTtA2LtXCN1biyOOak9OVo
ts4PerXlz5wUm+ZAc5GdW8ziwq3IYE4OlRUdOMeto+cz/f0d8Gh+HpeRLm+4zPKRemV9CVE4iZUA
EqtAglPOW1UGOszoH5q0aOb2oJUTjesCc74tjLvStSrBHlbA/DPpQt3FrFtFbNz70TMIeRTG5/UZ
Kwh+5ftoqp9vnRJloqZPKOVUFpyuX5KxGa/jQ1ouW85qrSt9bdxlYknqB1loeZVB2i6A0o/y9TSH
9fAUoTA4IuSMzEtwu+8Z/OJu94IONc+v6dAxb3Mg2NGI76MWFNdoyBDOAHOxLKlJ8QRb/N+MyykP
BV3eKhr8kPBADWb84dLjvHXD5mMRHbLfb7s8zWUNfksH0HYiuqmdrUaycoX5Dp9B6bpaERtFhCM3
FVvTCzq9bUR/SpOQq8Cnog1mQoeKIWpHSb/XEBJVBC4D47kcaSVildzL7q6kRY7ZlSJtsPKZSVen
UMO189/eX5QR/jRlLenFtJ2p7kCV4mqwnWMKJiswDJoMS8yD4Se8fjYCSrTf5UqBUhyN78fv0jmu
niApWdXiUh9bH0RJ0IQq6MJNrY3MGFh1+tDK1Z2mn3NTFVv22IQCisBVuxM5kafc5XHFXjfnQIZO
FDmKSpF4r1WAk+dPPcxbf3OPTo/QhYKASW96y3T/NQuodSDuBY8cEd9drhspaKrSHKluhgtT1fPc
dXya+Q+4mh4BoYaNo63Q7xhmaHO8jcr2uB7lYcLos35mc0OcO712TD20MNmLYsyiMK6s0GNzKom+
GqduaD+DvQQZLYDvVMNOvvtPBuHFojEJeL/4eVRgKpiJc3arZOqT5d31SQ68yY98SKBXzmpQEyOf
od6kh5NFWxIJg0RllqUeECauf2Hl935LzjlzDMaUDACKECgNA6TcIDI5c7+daNzal+TPQJBFgfKp
6d8nwXcDV2ncqThT6YOTiXygORIEDjE3nbSlTimd/6gBQpzRPOcWVDSwmwOAA/FtXjp6FSUglEXo
QRNeWTD/bJJshfT6YCaQlFdKzFqZUEeQ6Ai1DLmJ00GXYo9rokxne4H9X81ZuMsRKwbTi4jqqPfZ
PZgOdy8D9FAYgaR2s/iqMJ9hQv6Ww3SoG0dYQJEcr8fC6J+5wxOPq6iz/2RZp+MwJJACmwI+f88e
UGExhowvUaxbmUWuyhiQ4tirc/APieZHzq92lxbDCD908wMtJ5K1Rr7U/11DCXL9C0VhofkM1lYb
WiN3dXhFAOFsvrdbeWSQ96GEdt5ddXbGLV2UWYZhbA60mLyMWnMAdxG0yd/82NX84Z9s1/A7MxLk
jZ20DlH/M7o3UXCfsHzTl5xGCYGA3QFvA/FEFdG5H2OTMFzRu3rUjO6Yu3vU0t5fi6W6997fpqza
GB7wiN8WPSf9aT7PpTNTE7dD4QFgqoIORnSJB0KLBbcoF8yOyMHqkuMc8iM0kK4WqsbCw694tf8V
6FcEOiRKi8B9vhhkvFmKbsN8HBO24Y9iX7vuDnauNDuwBc4g/HOW1oaFVlyQYn/Q96aaJ5V3DY+z
ipPk/Tojf8qV7ul0C65y9RCx8uCOKQAkCqfZ5SYKesQxfH5m5M9H6lnNwbYDQkfO/17BaIGsLMQK
U1Oz/kxVJScfAqBuZD+wXPLBzUJouZgh+YWd0CH0aV9z1mdkTIHM00gCL6kkhRkGwnKJyWFHE294
itKQYyOPCl4wQoNVBSGmRXtXsm3OFcvQZcx5edwCC1xWxlIUI6Hr/YXE6SfKyrHCZ4SE8k3bwiuh
23kIazQpg4OTyIGJxKYKL4KqwlcBasH/onCe88aT+OhMXhkNuSXZf16PtGab3QeUqh3Gm7mkXYXD
xcr/FnoB0WmCSmFoF4htGqlyWTYEjVstSSJUq+7Rr+bsCeFg8wYqm4KXWCl/htDhM0MyhbTz43QI
2fPkhl1CeFu/VnhaPp93ntni+bz2k8ehM5IOnupSjh1OCA6saJcQnHEKgpsUmrQSG+Bz739kwj/c
Vs5ggA5exUq4gwh0Q5pn8q5ja3a0OVcAv6C39MDHmll12wfeu1T6z80IJSSLjcqiIh2KdD1CbYt+
lun3lAeJxo0gxw1WNOG8rF45vrLxyPg5nshL4AxDXZWvkbIuYbh7CWRI5DvRT+8toM5QiNB14xQJ
iySu8SwEC68yaRNTC9Vtxqa4ZVHX7Idu58343ECkDfPtY9+MdWR1fa4cPWuoQKdZmsb7sAcEvxmf
4OJTfWaqXl0uDgjpl3sV90213sCPj4kpO2UPSonRZsD6AFkcDsYs+Ny5YERckWlHXbGBfY4whHET
CMqne+Uf5HZJT2QbqlIjHOSz5txWstQUatBcjOQICj29EUafQdEVvmHT3IrleQo38W8OHTWq3ME3
9Oz7GlBGJ/cYOabqBWqCRKUh9HqkPHpwLe498n227W7G9SlPFw4aKQ0luM6RDRiZUdoGD80hSWma
dyaxgiuBjBWJMF35Xn2pNL3yXhtTr0bsuE/3nGWjlurtI9vvAmhx3ateHwfrNnS2Mc1Ueudg6jEz
BbNDvVc9gLPr56/0ZeK/wHKULOSyGe+Iy7fcMdGDf0kF8SLNIEWCGL88BCVOB4M+WYPykhYXsCit
BOeZjdkxku4MEntbsgLGWon12BZ0sOvcvtxMhyplJux3oTOgKELDJpEIdPml0p6lh1cctHFWgcK/
K4PIuVw3gtyrMn4WPVMUIKTCKx40y7ZMDHIMMRf1fLR6tqOZ90WJ/RSues+EJhXvgLVduyyEeFkK
EX+qcWJs4NQsRLuw1lMKxnOS/7AIZI6t+M5rMIBWQJTViiObQhNcjb5boXYdtbH+kny5xk4MZzl2
ZzORhv+wA/ZNMm9tjy7V3Z7whLESvSgpJ2DfML3WLQTRQFAONNs8Qm4R/cu8dzCpdcvEJZGEh5+v
jyemXYt5HD2FyUK3vkYjy0RL0DB97s5dwe7Jreypb7v8sGirPFj78Y3FX/ubxHmdor5Jn69247aa
CZ4K8RbScpxXsF4VMI+kgnjrpkCsB2JXtrgqdF/aRlR8j76MLlnDDtIweTP9rmbaM6MtGMFnFKsd
pizJHDzhDqDoUCgDz7QPnn/+u1LuSRiuvC62VAWxxEGx41TDZTvTTExEvCOFhz3b1Z6IJIi4UWOD
UjIlnNXrUBn3ThUIACL+GH7BsYy8tg9/NUKVzW2bTdE472TnVphl21mH/3FUYHdHbNbTHiKdbE0C
d0KJ3AUjqUVXE8ZyhqG53IhBM+tScfZ+G3rv/aDS3zvXPlXKPyofwwi3vJdCEwgspzdW6ZY9r8MG
oGYq4LtsILn6nQbjT86yn8RreGVJLW1s1dNdRRAA4FPCKvKqP25Sk8rrtczcJQeB8YES5Lw42yAO
eFndHTBZ+WPUxnKxbrrxWnXVyETELi3cwgtqreslOTwms1KIHI0Gor6lTvy2xsNSvdeoppixeYrM
oWOWloKQogto3SkvYUDqAJPXm6nvAQtxVCJCh2WPC+FO1HIwvAMrDSK0b/a2UY0XICO8w+8m+i4B
2yZjd6yYHdZF008INkOFc14O2tGu1EXLXZyJ6VnSEHpncc8VaJvLr4BoTndgCHD2TmBc57GkcdCd
JS8Lc6MDZjYgO3JKgt+cGan83wtpWuexQApqZFjqI+gb0FxHjLQ/8eLhsbMv6hpBHHRN0/ERqgsr
pGHsoEIiCcA7YmnO71+R0Et9AQndmOe3MpVR5myBKK4up077Ou8P+ehmxxZz8vsQpbzUzUsM5wxQ
4DilGmRpqiMxCTGciwhit8EuKDtpe2G3qiCM1NqLpWh9+n3AMWRMEVllwex6tfOuCxJQJhAoRlWc
jId8QJW/qjggaUP9nCkqAGmHn0BT/3Ul6NjvV3ADVdQbQRlX2eR1rRpn5RUj7FbRuKxXconcXvra
bsly2CkkTiZPldGLem3bZylVCwqEWpLWGYvM8NugGV9/yHmmYewOeeckMhVMLV2bpy8G1jhe2C5M
Og6uEPIu/3Us2GMGv+hbsSDvnU7Ek+I3hlCwSb9mGdMmlO/7xe3S5YZszFcS7F4X2jt3LZD1AMW9
iF7rkDdj7ifwYmjDGJ45wfUCxXwFy5pOPDU5Tnunvp/PFedkt4yrq/yTZHK5d8EloMZnfrx+Vh7H
FdXcDkQ9bMYfA49VzE+iSSfKCYpdQH9tTLLWYgfMakUvfj2QmIR0fTBB0o2JAVYn2i+RdehYap0b
q3i9zuPycT/pg9ULcZe2G929gCGY0/WI0yTAFdYDKa+9dsAKMuAoISdyGxMdi07Mgdzgz0k6gSyf
6Dc/FIwNCdrRy5H17btPhifRN9w1CMxkD3Tl53qKMBFp07Da4lIOTzzaYIQyj4ORLDGECsI8Km8S
6tNMJx2k1gX2YvRcf2/r5j0VaGDBOKv0NcWtRK7PjUhBuyqBRyButKnUZFfAC39PWYvGI7jrySyl
UuA8AmeHs4CBaO5vJ9m4eQWdBHYgaj9j6qW6JJTnp4q7wW/S5t1uJwMfa7bVaxTMy0RdrFN9V/sm
qob13z2hPz41i2M3hAwpKyvzCJ7rwFY0O5OtNKSCRi6M9t+SrnzTGLgwzJg0IPxanBi9EwzazXYk
66boCjtTJTDNNAvkVC5EkUV4tfVqAaU5cmFiHJWbE+VKGWGa1YjLAVezgJLpnKTkEMZEZ75YdyUm
fpUdvbEmpaULUHPMPagE/BLkYZ/vR7t7vzDY6KR529Y3iRcXcSu0Eo1cBG0hQxCiDEINn+sGkufq
d+J3azj0JTEuVlooz+XLew4V7NwzyXLYd+FEwOjuZvzN9A90EkYTr06smHSs2O7izcH0+B6yHZ+/
wKwTJyf43AMRHFamj2WELSypd43Socc1J/VRu3w4f+7Swrm5oJWb2I5GZZu8i/iehfITKszBihTp
bnR4weRfE6yAaPhfYIm+EL3rPtLtXgJlbH38KzsCykFtiraaSKCYDRTuX7C1rVIQAkodEStL02SI
FpHJXcH81fOYbGf0/QM1bxS1b9MNaAMzk3LmQC6G24Dq0uslcuMuribRnCzuwk/HgkWuQfX1ksrq
ie2CziZzY4PGo+FnXnDmbLmRyh5G0I/l/HygkX4M8PiojmmFBPZuH60gOEhv/X9SyDaXbFsBgdfC
LFlwOTX0aP1qh4zELqGQxk/L6PnHkBICNAgd8uUyXk9ehiYoFakMPj/b9Ulu3v+JjNIxhCBFlw03
TxfmX43viamadSez5AiyxfNT9T1a063ZVycIVZCnEmgDTrtkiWiQ3JwRPn6XPI0JVYVXJIeTxg01
DTNw77Ux8ClYXHdtrvzipfeOmgbFPUHZbNZFkVEKyVtlcvNroPTc3T7cIZ0p344z/OwypgHbnT9f
2Ebo0mnUDm08qugb7r1/tdJguX53N2wgHaBTUGJjkBglu5bvKdEAMcmdY2w+JHE58JauPmYordoZ
HUd8LUau1OxScqx+zZqFz89MOC0QoN2FBQS8sHGrGQjc9zpWsc+hFccjwVMojwWw6eEraMRJor38
pMh3ERSmz+D4oXSzVRXXnLx84WCSWviP9hCkUhGxtsOOWX5XXMEvcseSaXrxBJb1i7r9kKqTjzi0
RQdqA9MlTxx7bHHpDuEc52wiA/2339pVBPijAB70JWxkqb3gFpn75s094ECOIJTPu2O1Rrwe3tow
GfZQKYhWCVqWYeEI4IkSl3uOqq0VZujReZoa/MZcnEm+GESYEJgaXs7O/DeyjjaF+y6uoJNSMju6
DzwBen+/rO4RT1Fwr5vSggonHc/N0sVbTeawiQgr9+70NOA0r06e1+dadjDYm+4W5TANIMHNtBms
FlqipAqgvyO2T8/jlBH7Wu7B8DagY4+6fmTLxRLp02ZagNxt9dFh8MCTT6wRt22WA0jYCnC7i7sD
kwYjmMjknzo3kVcQs1bUiI71/+szg3dJMMr1eaIi5b9QLPMY+J2jgnHkerkfPQUGrdIkEq6U7RBx
iFxsVIkaFt4YykrVuOmyINsO9kKv+tCxqmVgQXXDTq0PexaBTznvklKNWfd5VvwVwsL8KKsYo1Ji
hICAHAp7mCgdpWSp32iA2/miCcMMw8mwo63A8CMKrzwZPEDxIXnNoyrQe0qEk8wNkqOw9gGa645C
t0BlqiOhXzez12TSeJJQc3PlPJVKqAUpWfgF/ywMPfFl1diEmImrHkLtifI90LDIJCyHGue75ujj
1GpsjJ0HJin09ZMgEzZ06bxWpcZTa7Mhz2uXRbc4m44WMxGwhL+Y5Gm3mL+Zs5WBsFD8ZjIH0F4w
cNzhXTkh/yCRqds9XbgeF6NYQirAL00E28wH04Na0ANxDWwVPayh2y5r0dhHli3B0eMeBiUJO3Fd
upHSpsX6uUVl0ztLdnmBBPHzsqy8Efel5t26nNjyB9DtnADPDx8ZdlilqKLS9B4bkIAy3jVLeUtI
x0H4+omxCOwkXKAmEy3mm5fujLcrg4ydIIvOKrApJaxkzLlMnB67ILXOmHzTco3bP4Il0d1js/1b
SL/9jsvgJ87TSmd1d+q/aJKGYTc34IerRoPrcknnFP919XwTgzJw1NtNGtGMLKE3Up/hGMbayE4J
DUOvROrUR7nBg38J95jZZXN/2oODjIMSZIg2+rclOliM34hTpoELOCsXN6EkIVxut1kQhvlX6kJX
g82sE3Fug3NxjuppHdQASO+f+rE4A5D2xBoto2mGKmow36cJ8B3TjOAtqsNUGiPpVCIg/d3v8XtA
BNuQt2bEMEx9ig4PREFXSk2JQxk4T0yLD9VfXKin+nmw+LrKfLpazF9Q6sPifluuwARfCdlu/GkU
7XEr9Yueyd1X0PnY/H3xrWNrC6jtNMtLU1GYpyHp6s/Q4vEKBKErgnr/XXqp2c7bfuBGaI2JDLYr
OpHL2H11sCWFWA3nGA22+ov+TodCnjMESf4gkaZhFOdqcLntfQYHRKcruDi0kEBa/t2GWd/2N+w+
enaWqiu/MF/8WQEiMt/S8MyGljaZDjj4Zey5b9xkPL4zNlF2Dca6Wo73x1smGiIF49ngfKKHOuTm
O5LOE4knQZBbLLidCf3KqUUgeLjJOfziJlQ5a94faJgqdmNSmZny8ywr5X9iPAop6S6w3bczYn64
ChgCVAkN3ehsaxmSS9NDXjMr7eemyDvZjbM0gx+LZMXZATEckkiE+0b9SAY2dQyBlSNa7RpfEmGH
bT/lypDNDqeWuAhxlPb/os6R027MOVpvq2DdZ1YZp2Kw3tDqfso0qcIRw9vjTOhBLm76rNsYZEB6
k4vHhwa0Ixp7mJS2cIpfnTanI0rTlYO9zQ+3R5OlUwFaPpC6JlfrvN2l/op3KE8gGtvS+M07DZxF
GahO0nQRGJBPhy+l+WxgEUD9Iq75ehQ6uq/qOWYdrnPlDzdvC1/xava4hpGP3lFe3ZxWgSTd4JjY
WqFwTLS9eiPcmtkfH0FRgbORQ+1iwKMOwyeqHSctBAiz2wn4ilbZxczsVQhf7GyNqQDNpgtqkIlA
iqw4sUjPVhYqKbsM5JlFc9BlOdKe0cvL0+9R4ohednEzUh1LNG6pePIKWqa40/QsljXpv4QuTwjZ
MsBrK3Zf2RfgvDQaOzYlf9X3kE+PGf73dqKgKscX1aL7zZospFYG42y27AxNAKBRJIEA/lAZkkjD
fjYczE2BvlRhlR077PA5+rllvHDHyJT1iMjTq1M4V25Nk98hB0uL3Owc/XAd1XO3ego4hszTW46H
/yu/7C/jwJWUoeIqpWhv7+nI+xb4Q2gI4tOuuhLR2aDuBuTyKJ7KP/T6pyRlqJqWDHemK9pslD6z
IiHSGMqgxmZrUfM6e54qvPOAflkHXamzw7W5w0TpiOG0wK397FTP+9qrOaI6mtj5A/5Z0WaJU3r1
pLH4JB8J61Nns7ihWF2mSB72Fc3g01SPDOXhkqLf0Kv6d70qft1llG3qt3f5kI566fn8Q+uQlTFL
OqrgwNFZy3OMufqTLTt27vuWv4RMd5Yq9+eAf5jEHHE7W776Rop2iW2dtKRjK1QokK8Aw7KxiJYI
dyerRVp08l6+iwuybNxaDobXYQCcM3ymASkUwvQQTxD5coemMM/sO2lmuMTStFraPFF9ZfUjVDzq
qSx8h/IyaVMjmjgOkkMyyyVDWEFmmULiMhVkE7AOxun1iDsAROWgYA8DS+joU7INgQ7nunjlEitG
xiGXoZWqKsRCoiWgPFa5ASE5p+25qcaP2/MM8qr+nVk3NYGd6gwkSP3ARom9IzB7JY73e4G9tgmH
5MPT8xG3u/ODBIuYIPLea588b8QhvVXb1W+APy6OkGHw5AofYKZvpWf3IleW8EsDoJu8PKIqTVVW
1BzxD7Jjlpl50VasZ9KfId2XNxC+emkw3RV4+ZReRJ5fUlbTo5VOnnkDtssN7g+D2cFYbL7GQkih
1YaCIowlrCeX4my0jnbe72wcHdC1jPK68e/XoJjG5tR/kX+wNAYij2OC7vXUNB2i9gDg6U0FFgjH
uvLD+z/1mbKOtGkjbmAcOHzkvJm4bPmCmWpxXRLkP1l/MS09IebDGGGoU3usjl7yzE43Gn4z7DT5
soanR1Na3cxgLELzP3HIr2q4nVpD5FiWfBJf0IGHDqf42SU66/5ekDOJtF5YUjMThClm7CY3YqtQ
T8TF1iFB5Vi+waqd+29jdMlzCZG968xy5eLRMyUI7H0bXTC054nVjgxMaONNEJiJG/YzzcWYVWwl
4mMLW4+8XoKtlhK+r0VO0HG8Q+z3jdYFl0wnRAyCZMFFLhNMGN4DW0XEA+PaOJAKGL7ICV4m0KIu
fQ+smwFkRuOwb/JF5kYastv9zpO4fulzMSLQH5KXlCe7smJPlPwiWkVObVneAELTslG0CM27KpEz
6nccx6RW8YUSoATRORUJinkMj0lQ5BrDyc78S/a84rkCpRS6UZRAtAqf3rxpjzCPUhFHpyif/1Zu
7GcgZIPsu+EwlIFz81q18jkupLSKHuJqhTBDQ1btRkFLqV55skQyF2Mvsti8xJ2SMisDvWpbH2/e
Zkk1aLAsK+S8/SnB9syXVdKuFXC//JvtDuGkpMmWqex5h8yVuLl0pxiOeA6HRslYq2jILp3DnqRw
+bOvnpDXYgR/ucelrRuWCVg664lEA3nskUW7Jg5DGKFAq/i6TrPxxI7fgWuk5w7CiIk3X6S0qAfO
TjltyL5o4U9bHotCprnkgPDHrAquH+BQlWy9k7J75hP+F7KieD/L6/Ub0eQ6uTcq9tcFuHCy4jpc
R6jaHsgi+BmyPbz2l1NQTED2ewAmlxJ6NrdZ2Zyqht2satrbuytIdZIfCVBEfXiX69ZPjx3LlNYx
u97t3sD6Fu9Hqo+kBVLfZCNXb+7d4A1hmqbHyADBr5i/gfE/Gi9dubeo5VipkzQummx6bwmtefB5
5Vz7e2Pd9fisZJCb486Tz2O4vn2JqY2pLT71Y1yfgH2C4KaZbr7s9/JsK+pvJlq9c5JLO1kVHDqR
HIdW7TxawcO7YJVJz+WgoOwgBQu5GUxWiyoNscHMFFVaJLoIDUyi4U7KxhzdBUwhSNUeJV4dUptN
964Z2mXKRZUga8FNlXN77cBcl5z2leG+bk4u1Lkw86ObkqDdj4R5Ba6ybJxOOS0mJuc7mUoWDRFP
UQJIvg2pO0aetjFoYxtJRtX1lEfNd/gIl4X/Q6GAG8ERqUli2DHoYrime9pdYS4HAMz8BjMzSPqZ
Wa9I3qVddEXGYShOrG97pNNxPb0OzZsL6bo1R2Lt45Nn4I4zycw+1cq554wAy5KRlIdg9DFXqrGT
8ACTILMGhQ1v3kUT7v4CWoXOCgS8LZ/ULyvxMlfmYQ8h2jpkSDjZaky8YjaNrec5xBM6qP8cDITX
pQwPZkgZyWk5nWlWtJRHeZIsgKAcLqkDmB3Ir5I3PN7ny/wkSEdEMPdCnrF1FydJq8yInJ/8waGv
9XEZYMogdAP83vzNEN97Qd0otJRHeS33JpGNscY1Ow2AT9vzsKtduDgNYxXiDfFPbIyOBI2pSIyK
mmeoiyturn9BnEGP9TCByz7WW9gh/Vu9KRtdjna88VQ+sHWFzZ97WyOCMoA2b4pCkRhmh8+VIscK
eSi7YBeIfyPY26XMfvvd/ju4SR7FNUC06evWWOV39k4PORyxJF+VZ66/V7Cx2sXzUVrkw254vIan
Gur+uS7tqMoq77MxpITvu2UcTq4pDA5yr8KXF3Gmow644hHKoanjfp1A9b0W7cs1epCNLYKz44gu
cJX6eO8DSK9IQWAjs2b/6k//L8th89h07LAh37scEWzUgueyP1XWrI5y1wBGtTjM3DvgpVrC9S2y
Z2nFX4EtMRfI1QpXdGi0XotrYuIgmzLa7ck0Wvw3Enog/JqXmzSZClib4ibjhoUnSGmp40KEMbFu
OtNhiu9V050Tk/O8CqnI33K7IWtC9byeQ5EN+AAyJAIRDGDeI6Ln3Ro2MVcZnaoV5Cww749nWVnA
dIg3u6QVgQTQZ8DN8Jq+dG/1HzOoDP5IMESwEyEZ17SnuLHGeQ11CvQSvdncwusg/9gaCJ2XFV0Y
4WHzamVBJJPApP++pcB8Wp96DiC/KOKsZfZv5S/ZbtNIijAmuOgifWROvcqEga1WECugWjiLAccQ
ifh0+P7vp+FisSpHpUdybzFhYldEjqYa2hPvv+1EEgV3WYZvgFW3DDGSy1qWCaVJM0qJVk+kOzsJ
/Z8p6GOEOQqNwOcTSxuT0jdHrilhRWOUMWKRiAXeqKH/Wyip1R7suEnfF2J6hUFCMpZR2097Uejd
ed2Lqr+Ue+hAJ9LxPBWruyjqD5hb0PhjOWRoCt+ZFWJrQ5yFSV38qKER/RAlCjbH/P2ZFvjJ3a/H
yMt9DVGML0PfFbVjqrxs9mEDuBQTr9+TiqyKnVLgWp67ZDz6iikJhHMCRBefByl61GWLk8bBH6Dz
E4mU7TF0+UjL53w5nDbY1h/FXWfsyJ8tqIN5ctJMPH0GYZMgBlhuhqGmArfWv2OV1WuE90PaMXkQ
oTLLX0JGVjTMz3RH/dZAfNXmrM1EijZ7rqnrKhgJ0mildkJ2GuKgQmpVkg1dANd9hZGq6xC+gyel
f8BvAZfx71V5I6wyo7tP1Fa+n5YmtzI/hQvPJxb1hgmqPPanCdRqrfbpz+VUPY/2Us5y404tOnTb
OLqv2cAl/xQ1YPqiLpykmbAOkYwaHMhco/VEWhxtbHns3jZSWfmpWftG2Ufhcjz1zOTa2UYtAZMZ
IxyFYMzwZ+dwtAmQJM8vLiOzlxEOZZbZ4hOt8vFoZ3o67hca14xUEOejqHFWW/3yngsm2ndB3dnU
ov95xKbtENsv3MpEguzCe5b5JrEkujg5cOWtj4rZ3w5NqgSBuaGLeq9EX7R9ykiBEDXoDpZqNqTj
czNowhm3l4tvuHLQbmiGXLD/rhIDWfmyKxRnnaBgI3ltscoGyOp5D3Q2Up6HvvEqb6ypo8HV39vH
kfhCHj8VtCIvnFbSX7nzXPQ8bPC2RnpQeAC2zGzHskW0sOVJGpz822821xcqV6Ufs7VnhaU6jbR0
QRtB2y5f7XK5SeW7sIc8EB2igVFXueG9lvlDbAhq03Ii4VYcdAUTmrEJB8FEmsm9F/pzWfF2UiHp
IH5Zu/kKCoSRSJk1JZTEpmjvRI928winy1F+aa0Li1iAYeWklPuXO0AalLmO4hzOstYUMrcWpE+8
er5WroAwbZNPCB7GF/FTcP2h2EDj/4tLSNMKwE95gO530/u9YO2IEZ7Z17uF2JD1mHWj1EtFqVa5
rS1mIPIwVHN5XDDZdU1AbmzizhLWt6xdbsdkicWTuLX3zLAx1PPXwGJ9aVHWu3UIif14ifXapiAY
GKgu2Lj3tNLMbcgM5j9c6R2D19Z9sA6nVjsFLFnwIh+qHIIDaEh6iwhyOoq81GTED5eYFgN43NeN
XpAsnsFNkRfMFnctk2wW2RZYSJ+PKsSJ4mt6b7hQpCP96qhJMLXeOX6rHAfDADUJNsUfmk2kdGSA
oCEiz6LoAn3I5kmOir3qJhfzjccLSUdbWEMs4mUtwOo4jTFWVj3ooe2/2BNfkbunH08bjWqJ0XkQ
JuAH/yjkLZu0ksQ430fNsBQgEOUBryjglrgESm3v5+ICv0X5yzUNfc3rXaF+FIdjoahDlP2uvhCT
ORaf2yOyz7gENWQ5lnC7gYJmNDw6a/K3k0mt5X+Oc2zHSMLrYW5E8zuKXb1Fc2ha5wBSU3cuosV2
KEewc7g1YAo5nW+WAad/Ubg8bEu96eWGouog7TVKUXTZwH1dJsexWkVaMwfFcG5WQ0WvaSZX1z16
e0bYTISwBceQJu+63kQW7vxDsWaToLf1JSpIiY6idmbLbek4CFDXInfV1OMYIJKdZwmKHxogUh36
fL48JH2GcGKvNTKBkgPP1XIwq3VcH4mTcSSNPX7tGUYcmX83LYKpDxXP9SlNoJfl30Zx5u4KyJWP
gynlax5wEsihMujb6v1lHyceM5Q5ZQqmSs0tOOCt8Ih+QQeu2fsWx/JZL96hSdzRVuF4/IWP7Iqz
na+W3ic3QGyPKBcKPfOPuIHmhyIkxgkZ4JXyW8iq7XPqFjdvqtyNlUBIZqY7W1/hRZ9ESqw5WgNu
P0mV5MY+dEZ2YlgwAP/fJ2heaGWMkBYd9FImLqQUKy1Afq3HpbXIjOqLLrdYSBXu+ZURTBrkA0c0
nE67c9Pln3ogGAgJnebiwwWaCi7bLa5QIoKukjF76icMhH1VO0GU9vrBKlay+EsziiZFR1R7uedH
QdjAn2DtC0+Ynpr3EviHJz46FKUf6HGujQjiZDcs+Ck9ATTTrcBP50omUV/pxjQlj8QosfnAs8X/
rX7Tji1jlANKHWvTzQ2hXuEFLPyUztx9mTGQzLaPKzSJI30usMFG2Iwo58NFXk3KGkmg65ZXuWqD
smPz1hz2vNjCs8wEDTgbuoaTmpK/yJn38T/z+Lk+g9EmbP+rIkVK2AZk4L8NsKFEs0rOVMRaVhvl
bts5LARXHv/t0+5Z7QZ83Tur28RG+Y87TX7qMvl3Gr8ukewTBFHst6nPqGA9lXqa+JRuVAWqRG8/
b+f6bEhaDlIh2GhHIVp+PF3SzqQ6xPDs/MhjKXQS9D6WhnBxjqoXhfbjOOxTlmWXcpVnVqJE3+nf
UITyfPRqJj3PCD/3orcZKQJxkZ98x3bsZAEARNNsdhS+nTWUVWpY+7Xb/V3qDeGFxwqJYIway/62
uvwwsJkz0rUArK85AcccN6krcBkhCu3p0WVfFmzeolmeL/BmIeIZ2PDBluySw4Jw6UlLhSPYNGaM
c+140toaP2X6Nxu4ncE0do7XIppr703f1vvEYAIEjKt0KA5cAJyekRmujRdUJTsv8OnFVeOqpQhP
vLI40C66LlKQJ3LxetdhdhLMrV6aGkTYF4G7jsWJYnJ8LRBbPjcPPL+2gSf83ISjNATEAk45XaJL
XlERL55OxNaa33r/7j96LmqfifKUQDTA9InE/C3j+UVK7E4BZ+/sI/1efa3pX49uJIAZYrg31A+D
4ZBUBhRG0uPOZLbggEcXheGj7bH/nUmW1mWDGX/qAEhIK9Uj5f+kFZSFEfqGUkjMJjQ57y2b8bIz
OaQvVVpox+Ef7RyhuvkdzUTu7KMQpecjVbYUox5iuQ/ObhrC+6JrSUFOVjE1Ah3yF88M8YzLIHmS
emUDLvmFRO0v9kLEifWvX8vqFIn+B3d/u1FBH2ODUJ4fVWK6vemCWZ9qes/zwMcuTEqt/Fl0mlUT
NHaeIdeZaoK1oWmzk2KYy+k7gbvFk57cANgZASjRe0zeQRZovcd8VCpqf6NW5v5KLvnKPTALM/eu
UwFi9eTayFRJO3BYeMB6AW616oHwyrX42ZnxUejtYIwtSe7H8nQ5s5iMdoL7aLZglKE3dD6o6nP5
AcaIMbYbZoFwQZEvd8bOygrObzCCXOn7VgySnLQ6IL084MckUZlJ5phDsDnk66ZChY6X6X6USFju
vpAFmPQbWbklH8IoCLziLxcTYnS+yTgzJs68COU1iG6H+TkDbQKubzp8N16PfSrZi3IG4pIy7Oct
paDONFxlFFUll/isHiAB5DxwRedz5owCShb+S2Yl8C8Oadk+IoYOoq08r/EM4U2Lea9SxGSB7S9e
K8ynufFqUeR5xsFug5ggxcLL0UBM/zeLVPCM6ld26CjQm2+HIsmg73DdVKg+nryrEvOxcMMLzPr3
8WnKSYG033mRpm9nGwUUtzm8x5j35XeH3y06hYmDaRxQhD2ZlIv7Jr39PybxYp3vpw9P5k01+eRt
OQoAxuAojJu63PNKYmmQIVMXCpy4jbZkhisRXJqhXDB9/2/d8qFCtYVQoC1atjTuCSRp9CyiHO+j
gOFoCP5VHNAz9+PAxbgAGVQPOHZhmTy3dxC/kopHbVB65gNiDYVSgC6ryuJiLi3rtccEpwScQBoz
WpW0la4aO5hJo2s+wJui4DSKGpbmEWUImJsv4od8FloW5EozMHdjPRiKXbM8v5VJEOfO3gNeaQGL
JtPOF1jIHEoS/otpu0UP/exk+W5/jfxXeoPLN8FrDVmCb3k/LW8V/gyNcyXHZKRruyUUpVJorDR7
Z2flOsi7ZVvAhfvMxlHFmrRbtViab1MUq12j1N2ms2qIWGE9JC5oeXJxx5fvpfPhlKQNQR4a++nd
1FaiDp2bX2QSLYbLZ26vE9Z5kLlKoJ0NeKWHf8eQtfLsS90UzjcOKxVUFKzUrDzgdwERsQyQz3F8
MLBOVOJwKYKyU8x+jswTfnK7h4FSYlkU8AyJgTk2u/ngRbmEeCGW06ikcR8pQrshWxsAotW1UrU8
Z8Pwswyig453axvTmkxrca7zDyR5TA8bSgiypshpm4B0wohKcxuoNvTFwwCihhqz5Z/yXl3H+OXr
0Ju2HlMKwKw9zcHOlnFWS3x0BXTXFTWIl81gMHkmv+aBA1RZMaLI7pTKnHlbvtFHEdGLPJDV7M2c
AYXezUMaXNH9nZrTvfZn7ixBHBzFlWKMYhOldfqhMql0flMbeinETx8GHS9c/XRktUhHSROgIcey
stZlHulvtV4fhXORNeep/7osWYAqbXFejHPsJvUPUOuSTsMmZLNvlH8MQh5TlijN9fRlBc0rOSpt
CrB3jD5acTZ6TUiPbQLVpx+tum6gy0MQgrrsjYjTZHYAvS1seAFP5qeywnRYI9ukfzuIW2vHTHFI
jkiBD5dS70pbH521gh6Uxk3N8TMNmnxC1q5jBwDDAFjccwxCDTx501HMj+F1I0fJhxIKnajtOMO8
amGDH8q7uPf18dAtzBJDjzQBx/88boSS6Ok0SxzQ/JWA4TXFlY2IBffEtp+Y4uI53oZy2JM+JGqY
rS0QXGDhyH6c7M6+u26FRCq1VeAXyO/1kJL7OaNQa8WJOHNzXHIA+uXGo1A/WsInp5u2XPkqnhee
kjwOGlfQzE6l5demLrbN3mrv+eGYShTbF/vKjypPQ+brQ9qUPf3ytpJXRb36s9x3UECQwT+WTegv
sHtlZQ7txkneiakomhuhZ8ZI6Mi2gcVL23lfHB/N56fjL6Wr4XVPDGYXRQqKPpZTmBCPTM3ZzNE5
hw7Aeyu0fbrjq1qVOPUB+wnu29rkxSCqsls1siqSZsN6KhP/WtjZ36p6Iga0u6pP3cC4QHEkcmu/
lNYB9YM+2GQOuEFD9384Xf4+IesZGmH5g2NRV5+0JIPhXrJxIJCIq1ZAOj2CyDT2OerM2pciREFl
P8HEsAjy+lZqZBUVjEvQ69Z0GShmORF1f/O48CVkGAUJcz8Qnid2nqPrFyv+meU8q9T8WgLA3ZPH
yBRv/T7Q4BoI1hPak++thRB3oB728y1Tro3YkZnNIJBgBGeEZV2iMQFZrrRdD69/iQ1XlaK8WzD5
7om/XiaY6rpAKXei9sdcSZuqr23Izy23+J7QfGo99txkIM/5CE5SdG8WMMNeShakgOQeRwAHeb6g
gKs9e3tI7hCq4EhxYUMB/nl61MGtb0tnhK+xZOwNhkrbFfvgEg4T81f4NfQ7twd00MZoCF9tiktS
Ml9JFjCmDwwbjeYcjxU8YNf2T2KeugwJrJ0KI8b47CC6/l38lvhhURA2+ccA4sfG4JhG2Oq7OQWs
qb6UPxzJ9IZRQpFyYrn9fH1Ag9LEGl7n/W2UeOuHEy2K9xrgrp1VM1e26MVwrflviKLs15UrlL9R
ZVCoyyEC5v+yyAtbAl7XDwYlDMsycYSjmamx3nMJlxr9+5lvsOGq6ZYLwP7t62KxgDFS+QYMzUqD
VjY0HIdigNpvBHoyfeBFeNYfrAqokMQsYl8IuHTkzmb22P47NitBqwWo7xXXL/Rz9NB2yrPSI4Hf
W7KlVN8R34c8o8hRHxR98i5nkOJs6aEP7ocAErvPPNcdtpZKfZLPABKGGmG5RtfUVVzdx5jFqXqb
OuMOaRAViklXmwJiJDpQKtdXY8IGwdgU3ExLb8eJjFrNYdqrpuH0dTwzQxy5+gnzcXSE/TH9/n1n
DSWz7GtgMjKsdgQq7Kunwmed8orlNIx5TDum4Smx8W6WaCEXFQhz/ZoXcbxf9clm4pAtguMqBOyD
hnX4K4hM/00EGchkhkcH0UA/aCtjtRFsllG6j1IpuJDuq54+JqF2ouSZEH6KG49JwLX3Qjc3TciA
A/P+Vys5AzP+CpRnMyVfd+Z8/iYJ+urT246ZsHlxW3dOWieRV6j29WKElhv64Z5xvxgHvazdfiAJ
dsc50QIDQ4gelQf43/m2PVhQfsI0IhLh/mI8kUsjWYZ7V1jPmNx2Y7WMG5d+o6VFS90RdTKUKmpk
sy6ugQCgPW1fPsLRJap8DdtXmQhKDnYstOp6texZHlKxrS7+yQR2Mv8cFvuUlNApguYSKbDDjMiN
16nI2TRo5KNwyuUvixacLlk5Xsqi//7Pz9SKREg3/xtixudPjOGX7Q8ymB7O+v67OWjNF+vJ5jrJ
ZSdKZwtLnd0mdDtwYeJ6BmZjlK5vKnOZ5+AILzF4YcxE69Bkia0vFExFrPF1JbI8tC7nwTJlYkSv
IqYughDfL7EuRRYI3u/hVwayuUbsrqkFyCAj+CHn3jhK31WgXPpsB5O0LFNsW/neCMGeFkaTsZnl
PRBDawUIsoJdB19cpCOapGfYf34jQZ+PVxqeKyIpq9NadX+Tjtt9ToAMZwmjoUO4zvjSARisYzOM
glTOSCSdK+slBQUmPT4rjHp03ATCSPePymvOoHRVqfDWlEeV9Fyz0bBiIdV7qaTbn9B8HUQpMI0d
VA/klP/vNqrmmOFC77q/xx8N+zOoKgdBfGwYMtdGVDUHLT4oWU8vEaxQ8eRlU/iDN8/QOmYg5jzx
ksb9vKbGXDhSVK+/b066Q1F4d9D2H7Sbbzlj8yLJojnPOWkXBUscMciNywRMGgDlEQdSgSHZjEQT
LpX8b6mH/tCBWqIQhfMDWHbJ8Wk2fcrWrj9elcHf0OEL9ecmf2tkQC0k3TzzcAYd6k167C6GjUtJ
YOA5bC0h+PJX5wNUPMPus05/jYyDIkJ7tH5uYw0IxDJrI9Owk7jkIVkVD4t3MMR9uWtMJlbcFnBU
MGZVxU8sEIV6U9ApWbxIqqnbPq7TQwRphHESvoKQCmJd7sHkaMpk/w7SzHY622gQ8TZPMVzha4/6
OhIleszDYepO7KZ3FUdZwGdImU3d0xlDv+pmDJS1h7B+J/jrtAqPYBmGO3UTRn2r1ll7N1/3R4x2
uNIWeZ58Uu14PfT9GlXwnyEELG7eoSjmnhjEAhFXzxozqTaetwqillS9oK0r6zgpfBsbgo1tzAMp
isZJZ3bvvrEyJf8pQwIN6PD+/k/cPNzQp50GmAkQLdThlhaTkHQTg/y6KnP0Qm9ztr6pky2Y+bx6
GXu7ZUzkJm1JKzvZZrCIBf79AEv0AEovCHOkMrcbANyd/SI9b87Jqd19vSEx+YXnOLvZxfpY6LUp
3wzYDkfRGQhyIJ/vDNiG05qYFozJIuhtiXkiV+yBpuDOd9BAM2vwa3RlzEgYA/oZeBAjZpusuJcp
fF8GTZNOqhhaL5PwPs5+Apl4lxzNYvOSh3x3XEIgNYUVaInuRcKDkYLZWSLp2yx3ZsoTGrZ9/Tbh
InzbGbYza4pFudztwZFLFwW+YGr4TuXDivR3KwOeAjeFLHZjvqGHBfcRZG1v/Me7JpPi7UIVtYAp
N9TV/tzYZ05/+Sc9Pj6BxiSGgdUlx5Nim5wF7k13WcWWOcenW1SPwouKTaWmUVfd/pjSxgOn4/XM
8WKJIqA7/rASSKfD61WKxw4K/sP4+1OeFVod5bksdxpoXKggrHSz7IYOPtHARYe//InlEoD/bxI9
6BceFyHdvhXKqXO1igtWCYIP/UPFyTW+5wceZVKaTu5JB+t1SpkHTtzCmXcH171A5F06OnvvcjnI
9zFQtVDPue1u5It+hrB1IZUFFCYu/0S0HMybhcLhTfHS5OoSCN1QgT/VPJaSUQpv4mtBFbYk3Q2s
S089hpO/gxljdP+a5BSell8LnJc5SbowgqL2mP5Jh0NNYB4JbvQH03R5FgJvq6x3ktSIfWJLBRpp
5m/tk6jljE7liItCbDpMuYsI7LEzLJrjVqlb3u24QyjaszBykJ1h80KXfdqn/lMke10wiVzcxMhQ
vBK/LnbrrTAUXfTGiawuKJrhMOhM0EjWFhy7j4lem3VRnOwCaJqYVGEm7l9G3tLYouLWZdB57yTq
fKobMLnCLKGUi0E9sS7DrUP7Fqr9c0xd1AA7Hyyf/ola8zhZkjYIpGXLwfBSFUbaFysYjpUZQtnt
yzPDjesfdqI6s92hVxFaVv+sCpNYKrDHHX2TZ/9Q9cfEqPfrQSZ3rpTFLvxrfsxzhWSg3v0/vG3i
q987bQSMRLuF1VYF3UuFlgU+MLPzLWQ+kgqxcGFEfJmtU9Q6TyZ2XWcxz3/9VmHvER7rbQIwnqns
npk9j7CArM3d4fuMswVg39xy2q1W+DWb1UaOXStE1w2wv1geIJTEkwRQvK7qL++aKrxcdAmK3F0n
f2ggvHdRws6p/XJ5FPx6qeinSeRtKf48SZOViAIicdQm0kPc2UISZGXRY4J1sDd7lKANL68MfEUx
ozy2IvuIQ9/sLFuyiLFnuxH/N1QeXAmcB5Nh7s5RB3k25E15Mtzd//r+pVSaVQFdkGWT5Sa+h+0q
q7x6Ip20CpBRcWcfS75obFuvefmalobVYNr6krH5OMyWqLZMicMWFynIaNaQcCwhYmE0stV+BIpQ
MlK6ytK/GRf2BEo+I176oGooAezqzJIxTtpjDCMmOhxkwdVYIFWLb/GOa9dbDZPnV2wJ81PK2kzB
wXJHDbLE6glInLlIy8EzP2wTbVIZHhNT8TixHkGV83tHb988LP79FE2L/1xNyKf35xnqrUdCM/LL
oLzOmx+8JwUB8nJPvJebNARDKS5ADyoPl1jGGV1Sb5T6nerUirxFnybnxy1opbf9B+WJgpNmnEPu
s11QW0MW8/gZ5xsdB7qwgiOe18eP+3Q9R9CR2yrunvFMZZxx7f+lkzVXPMS6sQqfW4jtsKJroAJa
HrpNlQ+HQNi1OXG3eOtKODxZawiHobptn514yNqnFrKQFOhlVG48mgXeDG21svjhzjbSooSiTRBK
hHx+899ZwNfOy02ncV/JibuaexhNuKH+WOvwXkSsytJ6jaUWWMafZstZocNmSBDVcCAuoLMQyz/d
YzWEdFRIrJn4vMs/Q9kT+u4c/Ss+Hxw8tPIHg+1R7tLu+RrKWp+/TVJQChYrfSCnydwYX6LqOuhf
un7/Sp8P033vQqWkXrQ7ZTLYy3vQmiSR2KbQhuXzprTKImbznqx5Ln8EM9A87xnPb7UM8x3cRywO
ka06Ykt/PL9aLEF9J1BCaFrscVIkBKVILLgvLp+/k84JTF5vw7Rv+7XW+5LNXLr9KD+AVTVZQjqt
mxiRJ+RRh4uAiR5VX9eqgx2yh2ia3ulv74Hdl5G5JGCVNJ9nqey6ng+dKeha8PUJqTS742q8B6CC
bu9kUI+41GKAi+tBYW6PDAEfLlEm2nU6aRWQVrD1ptcAKFCNGC3LsQSsJMxp5lUqZTKE1p0aZ7ns
l0QyGc94NAuFpIMiSdCFu5Y2rKK5gVb11C/StcGYutZ/pBNLyRHOKu3Wd8HEXSacwt2+EKMhbFTQ
gBvYprP4UAsT5jnCeWWx83+4PCyGgWgjRNspUgLXIU/JO4GIH1mGXU5fwFZMaNYHzpj6rfj1jKQZ
B39VWcZ5AlMpFb6zxzPVfNJ24+FWWUmA6VbETQo+z5Q2wIDwulI064dUVIDO2fVffXQw82XRpC6Z
ZAeMcCAKLa6YEdsFcGNngq3jsvlPyQKgZOjtO6zmAE/DMYJgWyyJnleSE793cvwwovWTSCCPNASM
hhu7l9BbYRi9chUUrSaVZ7W2aF7uwi4PDYNVFIredoqK2IGyg9z6YvQyh76b3SWCCZxaszDI7jE3
uPBKqYjX2IX5szyz5cnQb9izz6jIlPGM/sdm6cpfN8Litxv7XKAi7IDbIl7E5o3RZ5SGYAZ5g4hT
XWnMvOYNCN7T8NWwz4CL2P1e4Gh8zW5DlXo2CTs0/2jKG0JsY0xLASuQ/Og87vfUw5PgN/yNpb48
qvFV7MOwc6M/BcPbNy1c7BkEjKNOylkV8I5XTO91D4WjqLfl2t20ZtXtAh4ZagX8yg/dS6vtW2vJ
T1aR+qdhGZwEJUj/Bw/xj7jkoGT3JOSk6TskwjLJ8k61j2BvSQEuJ3+TUzj6qfP8lb93fvJDlvYs
AiZHUkoyfnNjM75j2UhF6bkmLWoDgB/UnoGrKQ2wpI2DIoUtt3B6BY/ejccCUPdvxVvj6g256+Kc
7vdzAh9m4jV0mTI9hquCv+oReU35up0yvB9woJLWmvOmTEc/euveKxylZ2FZBX55fL9VjmGRc0zh
9c3xdsljzDtiql8L0T5al2PHiNE994o/Qmc9vFFHOiuJ49ACsyolxoip873ov1/sFzb8GM9DHkLE
ebHm31xfybQFkLyCskvVbrQhSSFLXW0CTNXbgfjWxZXU9gMW0dHJJwiLxNrrfQ34W55NMR9EmtXZ
kpwVjB9tJMeks45T0TJuDTRLB7zp+37BB2s+wln//h1rUBx4JF9/rroPL0iVKlgE0iVt+XlC1oRm
z5QUOVbYcHfk2zwgZV+LSXP0YebUybXivCyqsMFIP10TpRAb9QnJmPLoCc9MhBQmacYhcTYtM52a
/SaCKzkHXOgJ8fCM+LTYfRScU8C0qYlJWxUgqBiQkONFR8ch73dIklfC0yPJfZOuD5zmY1KNODFf
28Gc7k8N7dVjgib7P3f8hI1YS0Ug/HymlhL9CFSvqiZLXGBb2DNI6VDtCpc0Fy2O4jiPzksMI6Jj
hX/usccOABJQjszxYTuOQa3Hl/o4cgoQ3UDvK5mtLKfSt9qpx76dH5U30LUzuP+YzWKFsTu8ttGp
ZqtugBO2hQqvg+NBzArfOl8aXsIACxy1q1CSjSkKJ40jmCMaoeSmcUyWFe/NN3tlmK9+iZhjkOft
Fz1PS/wv7QGo46mya615jVZIMOzEjhjRkM9XnL+bdTqmEjZWRdB+iqrKAYYCuGlryWrxSn1+dwfs
8pFMZ6bhGGYCAftCOBp8Jyy59Xj/g14y1F+Cb3+Pvz/snYE0ndMYmULQorS8CcnZcDLWFOErNcDV
VmNzqe4qF2pWHFhNdmGvLkqyuCAfD7M7lVoweQX0kSvBpORimfs+2lAax+Ng801+D4ksDIFCOrij
zd/q4EasIyIFk+jKCiDcuNh7Nvi9Q1NPCHc/Xew5TsbgvMZBGm2VL7OulfVaaCbS+4tIC2dHhw9o
7XKltvduwCZ6rHKhgZb0OxKklGf/UvOwJ7f7h5IxgVQWWGbIbcaSwubO4ZmTTpfOkDkDAczc4LrO
Mlr5KPzP1nQFPvcJ7I6r6iX/JFnBuTfDaAR/GMQFP732hZvY2S4+gYFKE+sayJXfxpmk912nvCwY
QPY8RkxUwNmby+BW8jv3FUm6UAyailrIDfgjLVyLiSzY/rjtPbc/TN4DUvKrqQ0SzmO0Xycbc/El
IXu1jmND/RN+Pefx3gU61JtRRavKQsNFIsRcG8ZRgVHl5BFF6izeJn4Iyoa4CaTVkYfM8Nai5CIF
/zjvDXeTgh4+CvNIl70dGkQLEluQZBAsoW9vUQZ1iO8qHf3fecgfuE1aPwIaBucXZSJgWI4CfpJ1
o/FItEWs06lZfquu64Bh0D6ZDjBJSa4c/gJFVF89uowWSbrNefpUNkRdS5PhhFsshnHsIezD+8X2
lnfl18U75GDEogp6wWb/0rNKZr8EawZLmpUYILo9JmebEBoRqItWhV6IfhPdYq9W9xKrRiyzJPjC
vfbcOLT+pwogQLMQ31EoJVkVLKHHGs8rhpQILZTyPNbEfhMRQknDmzD441G0V3DvBJYOf6d6CF5Q
HiM+gxVUZ0Ijw4ok59Zj8O35NpBLyW2g5aLS3w2To9zDAswTyZA27fYozX3Y92604BwySZMDx5fq
U590JlCxI/Z0rs3rgYM2H1bK0JUb+sjzk/io0ac38eLZXIBeK2gQ/wr532XESbF2fXBmptV87qe8
HUWtpWGAtpMgudxX7M85iaU/CY96pc/kYZokGYiRkiuYeEYCsPtIpLbj8XZ2ZN9wX+RhvdMH03yy
o54Yc6x/Be8SV+ueNz5+GJIsoyu5Uurh0/K41WEddwv+nAEva5+F/XSyNFb2q7UdGRdu3+WlQ2d+
L8XgRQNL4Tfs2FMebK3B+sQyvXs5s0eS6zuMbBAerJOB9TuwvuReYtrhu4bqSViOZal7QcM8s8qo
Kf/qjQdA+XnJ8ApBS9JvtkhGXAzv0kG8vxFr77ej1JCkFMj4EonJMfCHSBdW57UADbzjuITh/Rel
n4ZGf5LrS6bqEVzXC4ezB6uvJHZ79XTLa1vyHsaPt1QOsE7hfDtoSp6cyozKLL9qEVaOGVXiySla
umBQ5LWcCqycSiF2hjFo3kMfXxu6QvOSf7RHXWiuDMVjhEZQwOmeB6DrOz1xQjKsHulbY81sN4wS
pN1fQY6cV3i7eIT/LE9ycB5D7yHFEjlDzIK0WFVbZLnUiDA2/PCvHltHkMrBwWAD6t5kso2ur+xV
IH5VLe3sWbjAIk/FxJ1guN1MD/zC1akEsz/vWNkZEtvV2FxDmtXgWWjJCQF8ICd04Ck1wuhK/5uq
HwoK6n2cOZawPp/6PI6040+KbIZyx2HEUXW0uUqSq9Skg8Ku/iQBMmxOYfjEg+25hg1mThUOkiyy
hHh71NSpJslm+8n4ZzCHDh9MhQwc13FYIJfrFhaIusse25iPyWdc/7pByCZ3MPO3aHN/dEx15bUS
97LeP3YLACRbzqubr8aABxto/kJ3oA8EGusFGxmqilIVOpthGTd9eL6rpf31WOBo66St4kuV0Kw0
D25LLcEZYMwKYrJKZg4VyhrpkJDTKz2yGFEezKtLgvR33u0sF7Xua0IxhXOSUDNXXVEDaiP3nOsd
Pihcpe0C6Nu5e+jKthxcbccA7zfgLdfa3fyiS7amOmQip6DMz7sMCke2GeP5R9dZ4bt5i/ebHyIT
EKkq1FAGm/W5+3m8gEKFxfaRWnmVUzV7oM9/QxjxB6xmGFbgR69EmjPsNjDuyJvG+Pnx9HIP/c5h
KuE0mllPYwzTg+Y1kOQNmtfVXhufB9N00NH/c4vYZOgsnz2EC69JnmUZm4LmNrqKLl3guabOCvuU
XWABDfer+0ZLV+fnHzND7SB0dsXssxmf7t5gWfL0TABCPs1/rc2nCj5xOnwJ2vJbwldeVMqAJyk2
shaMaUxUK+W+m2zNvqfrJPUrA/FMQoR3VKd8lVPJsljttmJ7GlUTTFiQmt3wKGHmR5hpmfr+EM+z
SF07JhxZ3AFS3bzf0Z2GizjsVSKdZWAh5dNmoa2tAXS4NMIFsXHHWH73TKfF2YcAs8pVZQ+qYCPh
xce1rwxx4Ee5GRmsE6HTQ9pjiZMV4Kw+m/dXcjf22L4gfsB+xHNNQqTN6YRaWwz2VoDVwVvLUIdZ
kK6Kg22CN2QAKtqj+A13s8gEI4ZOPl6bUJeIHHEiL7zXycRfMEGWML4RF/eR474fWgeMtu0aviYj
/4JTrq0Vh/MLL346IAIORfzzvFkcQH6zo1g1OOC1P81yEp8aYVyYRc7NsZqm1BtVPktpiNd/KAb+
8YArnivfGaHylcOKvLnfC53+90gIFhS77i6KKPr1BUYEbzjzxf6orf0Ga2U3UqSdmdgMDrjhW4co
ZneGivnkw4Fhu+r1sL+/CAmXgJlO7kNk7XU+ufwb1szecsZg06CEDk22qhiaEMr41wAa2lq4p9aS
96wpUicDdTWJ9iTYhbDhyz5Dfp0wY9317G3LX9LVQ3pMoaNr4xESNfAhN4V3EGbZioU9Fz3t2/L7
he0A97YXVfxCF8UDGvi//inMeK71p88oEmhaXyRMoMdWGboxamDOpSBd0wVlh1Ec4b8IK9/+wci6
WnofAq0PJCWr5RpJG6L4Q5oCwEiVYIuHBScrNj4ozZli5E0E0F/5bdF5RJkO/9URqLTONa+rCgUB
NjiQXPWXuTcBmYBxKVMMXTxY42vjv9/xsr0l0iSX0yGjQ//RmowvnyYSx6sQqpeqFo/yBvMLfbil
AKqNpWhDuhUco/iPjNE6QpDk1CkAE9C7CCp2Lb7PEdrdStMTEJ+LzzOHdWpLxhP1jEjGHVqxhR0p
GDOUv+biuteGUh22FXpO9oIYeDWhEVxInQKdzYiu4NGmb1ppr5oaEV2CrkScF+HQSSWf8AXdDCiF
szEsAxIisB60aegGpUW0GXzDM8dOgFtqM8Hv/CbWW7lv+uvMS2BFaJeMPa5nUFo1EHc3fwgCBNif
lsRy/otTagIgs9WIsmAX6/2LX0fauYx/Jscjl69LlPD9RbJ6sZiOgWxtM7yTFmI7c5iN9tjCOHC2
EUuIqhJiseP+PcbhMmB9NV/7LOCbrcHCJuDRYA9Z3DpN9FEcSSk8HUWwaOzwUsPqcIznKUdf4rOE
gBTON/YfcyPSvI5zOMo4/sZclO8loAuzir5PtfKQx5bNyjJr/0gcWJSVjSl/ZOSgziticyJmK5O4
EQk6h/rGy066uTIKw7FbKl4LIa3C2o10bHEWXzrghotDVIBcLDkB6T5p1oYFxob4lqqdF2UhY1Yk
TrSQhJKCndAa0NObKGFqOvExzHlxCk9ZGpYYnE3cPzWvDp9AS07fqjWHRydY9GkI3bRn1t+6WYH9
ZJU18pox085OrgHfFqdP2tX0/yy8E7ozE6kVQbNuRogEFtt1w2J67kSwCQMxdvUBFtVYRe+TjR1v
Dfc4PQ5ja87LOEcwUmTO/m75CpcS9T7BYmjT/ma2MiJz2bv7ishs8FpfSDo/kvnmsTIJkTVqVjq+
0eqnQRFQXL/PwuuMTlBTRb4/RJQcwmGnk6feq9lLq09VPt/Ek+y4kI5fZhsAQj6CRd9ie8k6ZL1g
gnCVDXWegDwifku+ogRNFKXuh6YATK1q9JvpgjiMjOiMN+7kkuoPpnQQ6/f3u2D4cAnfc/onjMYZ
qCT3vuuNxqAe96qJpYNDYoWWMn6KH744F9Fzpi4f0sIL8KHl/pCjhQFJyY+uzuj1wBHnixZ9Pak6
iMZ7ADLZGWg5tQJlXI6QDX/1dWeRPKY3JiCDLn3fSKLSK3yQb8A3i4XAdV/48DucWRsO0ZzAUIuf
tmK0AqsLEnZYmOY6xhzR0CwAo/i1Xhdvn5qKhhaJb0D51ZmUs/zxrqGC9ztgnUdWi1EEhkWEYOCB
gUCd5jkcqExD9lxIdLYNAe6N32udxwAB2cYhnq3Eo2aUPUUcv2mJnD9kwuAh+z4H5OTpulYxBWf8
AY1FuChvWZi7JtAqlYNAcLviprMUlhgpBleATQTVpW1QyRMeC3SH1J3luHzQsFW+Y4nBoaZbDN42
N5ES6x43yD+iacpLWv/It3RoqjPs3Pi8mCHNiQGq0WCpDFN0sYtBeHmjkaNXOhw6M5dDz/pJzIbN
ovoPKa8nLy0jgNzAxBtArkk83oks6hWU4mdRJ1k/32eTtNBJIHK3ZFxS+YLor9/5WsjbcfHVJpjb
bhbJupJFMNbtLXtAclBaOL7mNVSp4LL580gXrO6mST/bBy72aCsZkErNeb8LfCMrygkYAkVIFtzK
LOSMkUqJFOu/z1SE+16Z5W8AC/57V86OrXpQHU6vxm8iyUhd6s506UwyIJLrpR/HFOTlycPvv2sJ
HKV9Ry5mgwchbGcUiQtztr6obwdMSTVX/Ikvv5cRy+THywfpzUo2n/2qGi8fVKHOfEQw6Z9cXeQ3
OZeQe0A6OmgiKCzJt8chLLQb8eSEwjgDcFI4jXwqOqR4MCTPTU4wg1Y9Hup2WhaZvAkgNO8MPU69
4KE3pzyua/Ji7/CSP8jLt3OJmbuNc/FQeSa0ciKDcZmCGrvNuO+tAxDdGxDzc7IltsQ2pp5STM3h
pCKjwNiOhyJTtHWW9KaXBpeuyGJyFjjQAaMQgVwVQycS6isL+Gk76VwBb0t4/e7CCzIzdg/c7yyi
285eX51g+wbFixLEaoNiVRRw+b+09GEe/xtXcvYbG4BVNQyincg3I5X9OaCTdJe0UK/7MpxEpXMm
kvF2zJwnhWMtTqd0dJ3YpPhZBJ+K1TPT9vBVSjVqPtci3yS9aBSi2FwdRiQxrUHzpUt4wBSbZJld
IPAHKzmkSjD53vracuKivVxH7/d4IjK18dBeLLbTZLB5QKA2QJ9+lmWqLLsekk6462PbOqK0V88r
mLc4eQT1dYQFLPkg+/s2aOabpME7gk8dzlMWwxSwcR03WFjOVyk7toJiCwAelKPUXnOSs70uvcBm
Bv45xf2FUhlwyVEK/1xZ1o44fKfYNcwuPRRva2Wmm66laEGF+dfuVmsZ09852erAdbjTKIv9cvQn
ce/MYfLwnA5ndpv9L/STjJWp8dcHzjdxoQM4WpZA5b2QCGj/qwoxVK9qzuJ5ZGhGCw+XPIra0YkQ
Ooq01bvv049jP55nz6L1uc6atlzw+KpjV8kN9WkRnGT6TkM6fLnCPKxIdJbhor6rAlC+3BXTDwDM
exkGqm1fLJSbNhY4NFOKQpvsy7+SA5PxOjlVykwW+TKc1X4yLGr6TGqtqeB/MgWXx7IHhGyShCJ7
Ikf83TKxfV9zro6bZM0T+ILf6Nu5NEC2gJI3d66fVZODX/+W8K9Lc+N35szD9sZ/wcuUVm1oKX1I
XnrEnkUpgTOgk8Y8X9jmFmjMnAFjk0SI3ji/Ui/0RoNARwT4Bngm6V1aBUAMI4dyLCaxXwei38x9
zHZr8jF7IVvlPiN840YNDFSUPUCvcrterXA31y4K3Q5ihPAPoRNyMEhgmZvMToDMjlERG2DIkHVB
VSrcz7IpQlfMygaOBjae8zoTprSV8T5276PADpz/UQHwhXPSLvNwN9PrVCiXcUIQRkx3eKmR243/
TfpAnDzF1S5dCTIuWKwBGwdyNmv9TFvurymF3Q+ioYSf/8K0kCzMCVoF15RhSwUw8LXQVwMtRd25
L1W3Q5EwELr1kTEeuAR/+wkmMOALvdWZ2SMAud/5Sbd96KTFzWA/Pqn4qaweZ1B8BJyFAPgqgNz8
TCWbLfpDFH44xS2hdnvLdhbyKvncZnU3JZ1ZwO0f70VjdSeyb/uDgi2S1SPMVAZ8iMCGhZ+et7yU
+SokUn3CEgUd5yO5GHUp9hUwGtV7KiFKhgrUT3C8qEyqQtEbmJqr/6OgthMVbtPf7Im+YHuCZ5Vh
4V6K5Y9awtsVTKm6sR1aORSolIKxBkgnTpQYwTSW2fAYU3M55mX/tB30uGWLxfZJb6xPeR1MtHFp
PXFmm0GbCHXwEVR1/cqFSjFogU8BNlfUmQT1VDjJ02u3mPyh3RN5ZG/GmseBc3uXaryYrvXohQIv
iQfHjlWGyWER1x1RglIo98ADM0wKdF3uE3Oeq3Ua3KBa8IrpJQlwrxzehfzRr1+yquhAt44uYi8H
iGn2InYUpJ+PkscVVd8htJgscrJNuGvZ9NqBXtOoD9ZTInytZoQIZiE0Yg/qy035D0B6ToqCKuZQ
MZJUKYpeE+lMJ8kEUcByQGN2VWCnTM0SK8lpy91sJldTkAh35lGa5XnjucLDMxft5l9CxBe5dmds
5RmZY8z5wfvoUdcQ6BOyyO+t3akes/q3IaeBGDwmxcE910MxjuUBE/8SzG4sydwNAHAAnwLX6oEo
S93EjebN2Oj/VYLyQtzGjdRfbybxy/pRwLJUQRxXRHjipwPs7MLdqYdnwFxKJdYLgqeJfdXkt7MS
LrwLX+1GTI54PEMtrP39rlReleFKaIpDiluI/heHElxU3Th6Mo7kIEjEV+t8GfbAK5JJrEAEtDfw
L045SeVjG722hUIgYZHbv7R+szriD01kLNyG/2C2fF06TIJQQrJg8NAitMBVD/VPaO2x79Hdk8SY
2ANVSi6y2ouUmK9lrcM9ITlVmxuAk/vbidlUcYxbdghpTKgM0gYl1yZTw+sYtEbl8KeVNKCmV4sH
BuAALI9IuOd1ky8lvXJjYON6/gMGhHfYoXXStcwtNwUrTMSqaWW879GeGkkEPf6q+Hcz6jb6eH79
ad6ZE3Rr1JDUujxuaUAF3uoMFVCx+V+GBsLxTfLWm+NTTaUFOrFI36SnvyVq584qUYLDgt20mOJj
jPZVGQWysenB3C03YStnHdqEJoDgtE6q2csqQgGw3mKiKrRgiJVFaappyRU7e2eh+TI88NMfFD9P
REhD05yWnSgr6AII+xJECLf/bcM3wMb2Ep+G25XCzWUcwnnAedCgUokusVuzDpHiQ3B8qrFtzDPM
7vb6UP3jZjAEmEM9jbHXE5VU3Doo6Kok7G8HsZzq9JNvhpo9Awx7JrXc1RfH38pBOa7xLf1Hm9wJ
KY73jv5jN0dP/KMVXpeaI3clAB9n1BMJYMR2QtCe43TGmsPu2FYqAOxJEkvTPueYnGz+n+791yZp
gIDZbMax/w17h+9mAODTggqxS3rmpg5ZvOcmnnjgxX9Vc0sz1WIHC2+XgQ16vNTtzMXU2TnLh8uo
n4WPnRuAu+UdraMj8023hmyIJicaWqjMFzcR1ZZ4calrDpdGKycJ7PSErrJRliQPKLpVAvdOoS9c
9ZOpvzlVEyGEAtIz9ujMInBa4xsv+LueHT/VkbfRoCvuNCgr3VvPxqRLOI9DoXzkboPcAMRHpZRG
RDJ9UNxlzAQF6Xk4emm5x/AwI412FYu831roTKIMaDN9T//hh1zo2YHMSSs2ITG5h2zaqTlq29sN
TV104Y/fxEh3fC/NO5Ap6bYZZvxB6emjCVOK2sP8XPNq+ZvKzJkuAp31y3Y1mreubkSt4ifVsC23
GAPDWvVZaxg46uFiOacx+3S4y2uxd4USHNXwikTm6SRd55acEKmc7gZ8EUg66qW2C/BImJ3fzojh
ASDgCvcW3bXCdt8my8EyKo2g2pqKU53nf/yKDTpfXVtL2Y4HJGbiz6kj5ZYKAMV5AVUa8aLDEFR6
kMEmIA6HeqIZuCKqXLGsWveiXBs3cEdJtRhhnUHF5llDBhFwH+jJ2JqScVdaVMLaRZGX2yp1fyD5
tarVwoYK5VUlSXlGOxDrpZVH+sfBygnMEyB58AJHdTOhPMRZBq0KIJJS7Qgh3oLX9iVjDA4wjuqB
rpWbNRcWxwpYOQQghFNpFcWLGGaYrYYDXknsPObFuBmOUb8uMP0Yl0SR/jZlaQySPcKdTvL4/zer
Z9g8ROIMVEfHXp3geJS3bCivSIvGgDeKwCuTFQ4MjKg2r974zaUTn+w4BdCrbWorVyF6E+rUQUsB
Hcwro+dESajglGXKAalABqFXl70Z9UMC0PFLmWfi8n21eqNZJ0rJhNYGpW45D1aRjqSdnj6aGXK4
gzjPE7Ey4nyiw9lTMLDkXtw3HtVOuX21hOjerDMRIcLzhHCYo34xsUCTsi82yTidaWUyfZsgXjga
v9P8yPC20o0xFygk0BrYYhhHuYI/NENXkjCdelAgZ0yrP//3TEsK3tfTqzIZsvxBmw6+Y7b1AEj7
7l+BXvJ2HQT4asyZT5Q8dgS6eUMYeS7OH4QZrZSihTOHyVFV3JTX5t4vFWEDYQjCAQDh2QWGbW3y
AamMEXpqxLyqz2R4xhkoY6gS91DnhIpQf1a2671MXLQZzKT62RjHzj65w35NixIg0du6/JMVuypA
DxTwyYVAsCRl6FhV+2vx+7cINucxFQyKPw+HdoktUVgR56lmvUsZi/MHfWEckRXwgtgSpl4xO186
xBjqKXTCVCOQGb8liwSpBHUKH8/n6xDlm5ldavC6oWIzdIp92esIW4HHmlrHlflkf0emyleNlmhC
QmBh5mbD7e9miTYsASWp6zuAUdMfLqo9ZyR1Y2gWYKjsXEIsNCby7MrYoKRclowMN2GybFnbd/Q+
8J8YsaGk9C6X6ocXuKaOHwXR9czFq9iDiqAXGUiKU0veRoqSk8ZwBN5LQzt4ejEi7BB2c9PtaE1V
xnYctyYUExmgNGiStNc8aYXOjihIjcE/WDPasRjmMFgUslmN2BQfyoYFlOTE1EaoTOr6ku6xV0ep
0bEXGk13q9v6OMXGZ1+KAphmtXsG8l5pvxgb7+uIemG1g/TtMlfINEhDtCuya3Bs3vGwqhlRrTvU
KsCIhQwm228Cx9V+WQfVxL6zNUkJ8aBqtr0bTGiRPpLvUWUj6YHW+CnhzuPjGRp/Q+vTRf9kGdHD
LCEn3rNnsl/+kfjhg80rlmUUbUtRWYb/mLuouQB9zL6MJ/KqBO/z3YtsTi6BKkqd49tPZwfYXuKn
Grt6pXKxdBGU0aDKKV0NXHPvzF3eO2N5Mhfho2+3mZ4Q2PoxalURY69Z5BMXeyO4iKdSZTRohDWx
Sv8H1AqHtkMyA7lsm4l/u+yqXIssieD3ZuYs9hnbQdEcApO3i2nWy+RJFoFEgimtmfyUTHZ/OYYV
lKMR/kii+qyjOp6MKCfHJ09MuhHfLIbGNlcDAt9q4C1jGJDvfBBDYMFeKJ2754AHEB90yjzeZgoT
z4t2b6eARZ70bWLTerYzhq1pbGEjzAEq8x3I69nXDHkTHaI2WO550Z6y+z+C0Ss+EGc9/gAni8Ti
P+XIHqV4+jJvCOOvRQPTM0egdK6iO6CImLfWSZfNiIZrXjf6iFlKf6r290fLR6lFzE1ZahDwvGnc
b0wsOv/utMffDmM1A443CtiJaCIlTRq2gQgRp+uhJ+Gxej5jgtw5ch6WdSqbTeyfPmJ6IGc4YcNR
yz5VdqXFtgEMcGgAsRnMOmEyo1J3Rc09o9+/Eyy/ddoxwy5Ffpz/nTZXOWmj2/uJS+FvMtnKvBxF
4quKs4j8MKRbJ9dRHJvf3JcAdDu0FeON+R0l5bNJX8rqZlp8tGyRDqys3X/PDm/78LlyC/wnEMcE
1v6A1fiVgZ6O7ZlnmbGhXXbbuNVhaa6/y1A4Zwabd6W1IjPp0fQ4ZmZcocnhsprTmGMNMrL25usp
99vHAIOBuZAsiCkTkcVwhUgK7ODT35R82J0Xos6Kgry2js3m9MYJI30/hJJgtTSoKjpAvMvlhVOy
BMrwKr8C2MtQD1jge2lfp1gMWBectSFP7TbCqkvs07ohHvsIH2f4tYJvqA7aOxyY9kLbRVLqWktp
IXzl20zR04Ptc2tNJGxR54VTxXayRPPUw0xcuXFy372CCvh6CcvZRdgejCPIvXmRtAUEhog7UvHI
7jyNFN/kmN3JvpwyqfDtrA5eAD35uqEQrzrsqaDCH0OiTjmPEvRUhup6zh5PyBj1fJYGB5NXbhzV
vZPL5rGGP7FIRULq5gXzSRFwny77xiG9fzB+qJpAETCOEPHWS4JILw8yBQV++z5y0nqTCjM1l8+/
zA8v24WbufwcY8ZdTrnIu9pbFz1bWaSsAbdmSX7q97AmL0G+7IgzUCAGXKnp5MgnRpu1EqhLRIIz
LfV3Wcj69s5qpRnkwT/wWLANjHZMmHP7Xm6yU2MO1Z7k9k42LO8aGP0pgrHlGrbSYsoNMQsF29Lv
f/JDZdA1KzbylyjaH0VNKT71baygWUelS6t4os0F8C8lynEwNcWzEHj3o2bHd5XbpF4ZzCAiDUAb
lQDGEPQfl8kxZHNsOkNBmK8L3HSaWnifA68Oj2KhhRFBpvFm+P1KNAR5RlFBl8rBZesKUrrfvRc+
SkZkzCKJAWDowALI83FP16/zKv6zESjuQ8/8gT1N0n6XwKvJnMw1KFyIRZp21xiNBjD+srj3cOXp
4a3bxhhT4lQD4QmVFVjejh8lfyzokGCjleWxCoCgeS/oMrckl3Qqy46d4qLae9+/VBD5cyCg52QG
l2ecivZdFiaK+Hu7seSE0Kqpv1vV/w1Z6/E6OTT+5YhSCtMABQfVO5bBjGyYQsEnwD9grmJjBouB
kc7/ijMKEpCJwAjhAvCafugXnXa1rAY2InnvYqbcRGCdNTqWkzqehamHRctwUANjisl44HNcSjAg
ZCRPc7Ws9w5PcjwELQf9tv3BkhFrfZkaae7Ba7gInsNahJKhgreGPxh0XXIMiOZOBGoItvDyUuAU
OPAAPBE7UdN6S1JysVwNxrMfFd3xiQDzqrCEZQ4VEDzPJAyXddAamfhHR/qj9VlY5iM3yIbpyWlP
lcNCz4YVwivCzbthabJDHx9KoB5fvYiF+FzqwH1oR71j/3wM7EX1gIo+jezITNVCxIxahL7bZdWk
o4WSt0hfjuYNbbh8cE1AKtXGIBLJ1Zamx0YVLw67Y5ZJcg9Ou9brZwgCU5UmK1omkXIgM9wHo43v
RHWNayUnvhFAKTFZM87XyGX0q0iFYO8J0wjOZjme7gV4r9P8A8zlxUGKCmEabMnPkWk72QonNm4B
WlH5YRBk2J1CZiEN6xe1mneT14ZQuvyriyjrsjoAKe/OCSB/Q/dVMATqtUp7i/qUs9bAvon6tP3b
8Zsu2GA/UMrgyLjqFftqyjgkH2Vxs7Vl3xKVtSLxNFKHNLTEq5+aPb91FvN/mrUaW5GlA9HTyrnX
U3J483pDNQMubdtfEvqLfylLJgU94Dnd5o6Fk9Kc8jYbr6QPy5HiSL1XSi61BufN/urNtRjTWPl4
H6TSi/xebXgjqk+7fuRBJ+Zqoua9Vsgnmkqh/elB2+lh2D8AD4sC+IWxkQyVItTBXwDTxXuiDFZE
0miACVBlZIauN8IA/aOx9nAWrcaYhzeJVntGdV6JhkNInE0+h5kYpPRVPN2PgE9fLo1ag91lELZj
u0iZFYKXCkqmW70hofcleARiz4yDVX49M/ZgUCErxjhcc7JSil3XXPYrTYYBM671tGH5tHBGbUSe
qvsPZuh3THxWv/EQefBgFgy/J0ymksargzMVJiGVXR/gFfAUKlU8ypj51jhZQMna8TgZzPbb34L1
ZkVtVorJPYggYd1dNTJ0+QVW+ArFpsS4XLT5QVVBOBNfvTIL+pgmVPWkNmZVcZi4ZvymL5JIJerv
0P/ykY1P0DaH7L17s0Dm7FnR8BiA23GqP1l4OzKqvszltxCIafS1Vsh69W80gWNpWOx+w0vUnOKW
yGrM034SB6q3dba9sgCEOK8KLHaNpp8eUjTuXa6OpDniWybuGCKp/kikEI6bR9R8CRsC/JRZYQx2
GLseVlCsiKcWB9cqh2E5AyDAu+caURaJm+4+L1S6I0Q/C/sDx51oeNNmy/DgedggkHC7rJhV2TOe
koM7tSaJXWNtqTyvNBFZRhiAPkamVA5vTNu2juBpRS2jQzpnksbk8as/vDOAdZBuVpdEFmXvnBHo
nm0zUSR4YTPFjVBMePKQfVB5IYiVs1ARUF2hpM3ICp07ES+NTqh53UK7YLsGh8zLoLuRIW7dRrD/
Dw0ka4pGCh28VxuijI9VKfbsKWPRayxzo8o8IJxSfW91Z5R3R02T2xtVjAgAUxsNltwcss+0cRjj
txydSf4EkF7rVcCr/IMmk1wWriAgRIoPvupl3nHgDUYCPLp8APbgavfVDpMJhMLoWQOEcIxRXwtj
VokrwBXyiHrDS4sM7iVLesZE0xBa7J/vLBiLczsGhzlp3Kptepk64pqCGucbZjfMbzwmVKK0hPpi
rQKsB+rXU7iTzyZQAu2Hj+JVVPT7TzICWwWUWzSC8dQ/B0Bz8Z+FnF/kgIiKkUvbskc4t5auCkcp
V+t6G785UkXr5+hlWWQ2arWk24wxu5dtJa2XDHpghaPNeBPCFN8h8sPqejJUztCJybNHCpvKQ/QG
i5RcCyNej1NP9VgMsOYqmK47FPzjwhuVdGBbmjxOu6nPTn44XuzvgmQgP10bZuO7kZOH3zt4y20X
ZgCWyrfJ5vd2x5BJ8/s0eyFYnJOkCCYYPJEM13dQDepO6voW+1B+CIP2RZwHZrQd3WEGsakfoJg1
CSTunmCZbULtyzLHu+P9JDh0xkfIeQ2IuttfqqK6+5uXKElO35x4q+f1wMfO3cP7pfP7ULcCJLul
s43u5hB1DV9WpVlCUrO922+n0jVLcMazADpdBdyxuEqi1/3XfoLJpS5ZXK62pJ3ixM0JcrXsEaBr
fo2mF8ZsndGDpeCJq9VMvoYdT5Pcq6EauOTknUdmKIxWXYIna4VWhJDBwkkPx5u4MAs4QT4fSv1C
c8DMI6jehHyElaaFFoDB92ysZrqIuyXH7g/71TdlwlZXl5wBdL4ju6yO6J+HGJ0VkOWi/YLrlvQv
o8R4EpvYD5ypCeZ06YfDeanh2CvQhyMnLElDWV4Oj08LM2pzTib3t7MfagjK2VX6T9MpcZ7k3QIM
9iCiSPMJiKkrZckwV+JMQjjf80xEm5w9gm90xyaxgc7wusO85kp8d3ps2Y2y320eQRLdismcoLM1
yu8wU46lGNRd1ppdbn2JktagFMJr2X6sG8FzgcLEijFh6B7jGqmJYySB9hni25FnweX1NfFHqH4L
mL1gbwf2tVBr6Uv9g9e9KqgRY8ure2tNXWpxUsIML/eKi8jmO0f0Q0mJDZdvTnrEI662Ctky0Xlw
UYMqKa7s0znkLskXUMJwdH4RMn+XTTVQOATsKopkzkGjt5fG5O8dzy7oKHdQRjKkpFyETnqLB8B0
HdzgB+o1viGxk4zq5YfMwdWbKQa1vxyVXsUIPnES+PZNaWZ3l+hvHn6va/VdwCe6Jfh8IIg3u5se
65AC+LiNaOYenO3Thhx2LGMElfeyPUhJDDjhNF+OXIsVjpUukDGI5eTkpSW3VvId1ydwLz7ZjweY
3X6CAbtkPF9EIG3KKLsyH4BA9L3euuZ7xNKM7xH9TGqa8O8UqkKXjFx2Ao5T9tZUJDo2tkobmmK6
TRhdJEZUzwTGyoe6T8QpYVWMOjxRfMtixLbseQNqQHCnMpxq9B+48O5PuNdux1z3Flm12G37kUAW
Us3yMXJuGrYH2efq4/RIPe1AAOVxPLlpqx85vHSkPbk3DRdc3JALivnNatAPNl/FYMUOy5VMmABm
8cJ+dcZCfDQBOxdpIU8o3wGg2AcHhVcfKmobdSnd0tKbhQ3rZ4achEV7kDZWxbubfsVz0zriqcc/
39ONTOEywJQ0FaPEcMVX9eMEBmzx+Tci0X0c+32IE4Sv/cCVEaobzzc3V7XNIHu8zaBqP+6IUHw0
fYB+uYWxDjYiJKryJCkqVenS2P0+m6GXfTrMK4EXRfJa8wSqxW2iAY9fuFIjwDx32htMr3TpUFeA
Kox5eBkMMVAwjpotv4u4RWlkFqQ8LqP9BwUpvUgt1iRSTMUNFeIloSkl+W0KoSNZ1zBKgeAXjhd9
TVd0h1e+G7wiqkcCZ+Hpt1M31prfor1qUa0Dx6UmGoT30FCcvgyNHUJNQ0XPM5bken4WRVwyY3aG
CtT8kb7aU3X2u7y0eFIVv5sSlXo0SFYj7FN2ImtJ38jQsuv+BvAutDpN9Tk9Z7dKZq/+0irN7Wje
uqBLrBz0bnNhncvYHdPXHekmCRh+3aGbqHY6vyzCR+lzBGG9WX/G5PIuAbOYQkYK/jTpmp2Vm4og
Wh8MD9QySr4nc3qQQSdSzJ6siu0X0XDIqTFDOe/QBX5br6giM44ut16F8wfGBQMLFNVpTWmsXvAP
74zdkdArYovDafdWWi8Vsd1jWM2Be8FsZdtPRX8MxpqYaHG7y9iXdMdUlF159lJagEy8HHRCRx1S
QF9XCO31GQUbC8CssCBlxQExejlKxcLyQmQ3eBCrz22nMK23SFyEZZxN0jN+vK28/oQjPO3dG0O8
7yuRgLgN1tn6eq6a+g2yDbp6HG1PqI8q5UQbrnjoJYQUXM+WWwumpSbHe7jFfvkW08ICXmKIUSA8
Ot6UvSmOjBM1I2KMHbVDPnIa0VbcX5Zx9LsVbBNsJxNVqxBt4CpDPaYe67FwDYBoegHEAYDG0K+z
N2gtVYPXtAhsSVUd4jjwp9xIU/2cjEOHPdexPLIVwc8qzS52M/ek07arfPhffc+sLCGJQdoEafjQ
KHq0u/BgKKAtCVsDFiXwG4phPxkKQj1sBSGI1WlMBv7wSeo2uIucXGqvyc1Ue5gVYwAOvXdNSJxW
MLKiCuVDrssJO547rLk5rQYIDQ414pS+ssYr3OF3RalFCwuFAG5pqI/ncFZ6rg1gGDtWp10ZrqdJ
xpS0P4eo9nt7XOW+8snTiXm7XtbS3qjVyd0uRJRcTFptUhNe8C7k5UHH/TN+SezSOhMsaj/hpq2g
wZZfTdoEZJxL3Q3ibT3y55YzOV8bb9Gpv+yb8DnzSWa8f2l5bF1p2M6ROpz9vVdnt+3UTQpLYe4E
ycmAB5XMVZk0T8LOq3pgZD0p3z0cUvAHaNN3Y8Vi2b+qMbMoGNlqZR1H1Pa2HWFQXIB4T4Xli8Ok
kvpoFt3HYDmB60lyPEvnm9PLueCfAhHf7g5WcMGhJ7VHQ8qNDt6A3AJYMQJctusNy8POdcrY6XJZ
WcCFjf3hCok8j3TZUNiZHH0T/D+Xo9EEy44UX5eZ5w6h9DiPiGhqTsJXC5UY6SQfF6lPgfwuY0Eq
w+p124RxlWtaiz3Lqjb6X6iAuEWuOuYnzgn1qVqEodkqUSN+t5BCbSolVfVVTVVtvIZ9x/w+qONm
07LEuFtiTq3g6dOYCGu5n0P0iMNo5X0DcCal6UbFF9hJxEjI3crFlcqKLz7yJ3uTJWsG9uPvqioo
nfsELCQ7bwSbN69tRry1NGxa5rmnAuefQEVDZXKtiGpd+G7ogDR5RQ0NAQ7arIpFgNVJ90N8o8X7
JoRLZooxRWaUuPYD7/hkdbmGxVeE5lclOMjfsrASIsLJbaWCBc7MPDMskfgkKyfkWBCVTaPbNzG1
c9uskJ+wFG/fA5P9lzmS7JjtxIz3YaIMdZuy1+38gmkFhAkn4W1FNLGtLAs/j+ON5I62aT2n+a/L
cep5yxJJXjp7B1Vf5tqfBrHyuch/SVOEV3aUG5qxLkrpAw5NX5ZEZ37+wiCuYtvZYVf53fFFGvmR
065lPHrYxyNBvDxZe19B6R8muxzQYEhLzPlpypy3yVD+4S3shDBBJ46A/pksg4jpq5E4HSzz9QDR
4+OoqpZa2sTyJX+Z7lamY8ukMFydIhuX5sjldJ8otcgA1r+MWOm2xnqC+ZaUmK87H3pMhZvm9RmT
t/GtyA3hPKJWTckbhwNFZUX+cIthkFbJQVsVJ7WMVL0IgAoVxXyY45Q5d1Zgct80tXlpNWrcHXZf
oPUAnqGSgzv+2uymk+t0XQPcr7UgmKCNVmJLvVxDPAA+ZCo/40CdHlT1ZCeDEjBLD4Z5G1dU+OTY
rIa7Eo1s72volTlRzcbLHZQLeelKn98gkluTSizCB0oWu9QzKJ4qx7EGJFpNsoOpnnLEpn0c33Xq
Ktdm7ZoXvCAOzcdRf+2EbwEqBfMIkUcSFOM0QTghVXVU1BFtVqEihro13nwLQHNOeP+z0an9WsPZ
A3iirjZLK6xomr6SMlUneXYltz4xflU/Z7ouThz3ewiW3N8Ps8j07cWuGNNr1Oj/ej5dqgl4ODdj
7fFbVJPaEjN63xJaA9ug9zC8Faxx/5WMJYNG1jCj1ZXv8Ea9+VP/TsiZ4DRfgUcGkH/ZSHCOA+mq
iJtde1ZiV6M3G4p1EPLq1x7C9LkF+YXW1GJ3wMr+Ze1F/YlHHL0bz2yqdLiZH+ll4kX+nmEJoIsz
uMfT6pkprFuYDrziKE9mTjH2T4hstDgpDNVo2ZwGu9mYz2e1wuj/9FhZcs8EdkrKxsEpB9t0wewb
L1V3oGFQM/EtNDBteasoXlZJR/hjVYcFr1eQJnTJZdRTg4F/1yZobnCJ0T/+KdzF58zlCYZH4eUF
G3Gx6wQZVLUXjixL6828l5PPnDAXzvECPpbdqd5wBmHHLfHG/1CW/0ujisiWBbe7TLSRS5WWMLMy
yxHVAPDwRwDGZ7TdRxl29tilqntC6/IBfHL+oV13b1O4FJhFK4fUBvD0cbyENbBGgVZjyX2vk6W+
MGYnkfFOMBSAba/VcPDMWFL/WohmjkEYriFuJk4S0+7BwKKs7EFIhTTUi9YHlrLLTPMZIjQWCCoO
2YzLQIyHZNUsgILf1ZRHi2EXZLfD28RQ8fav38+856JpLMP8suohcXOctG2J5Ivjv6U0E+dGT9k6
G9h0v54n+UMMwlnSiJwE3JLy0IkANycdCjQv6WO6hvV5pCEaVRWV45tc2IcjclTjCP3UCkPWBfNW
58rBaWfT6Uil56RZoqU8lkOMHvwcdZEjeNdcqOkT7UOpUZ6KzLH/wp421JU7RUhizL+O4AQ3KlQ7
2gckYgNZFkikDIHNVD954c9IAM7fv6mooPNgI0EhT1M3LckR6VFvXofLuulKvcTDwTge8Ep+k72/
W3m4L7J8b1Xb2BrfA1YP6TiED2+0vredf0L+f4I1L5/UneZDPTSBSSLUqLQbUMFmR1K/QFFD0ypk
sRnY60yijXLljpZYl3zxlmURVbFkmw/KWmBhfh+Fs7V2RncneFyLZjMlZnUXFkyn3+tJNhasOPJw
8UnzSxy7wxCMQw8ckZbWupFC2+hnruaj7fIhcIwoi+6I/1h4LIYDrTnmNVcbgd80e6ROL+UTMx/y
omYU6Ikk+3s2IZOguvxXLnQj7BEXGqegafElQ4uI+B104v68mov4R1Ov0ZxKUoM6DVLRNN3keLYZ
dKBEPK5ZsePiBCtvDoAWOsHNFj5buooK/MNpJi3/wDnz2/LyEKa5dIA79sMHRrat+0XD5x0xY94M
yEf+8R3zaRf3bDgk6M5DXo6goasZkxoq5PLCXFeWB81RjYc59MY3bZnBKjUtbw/WTUfxspy/H+yz
Tx4uh0li6WW9p7KHTYg6+X/Cd1q8N5YcRBSpLUpnOe9esXvFEQE5Knyl/Cqw3qR83MpsrthcUCEZ
6LJWDERjsBqJOkFvaKkWuf6RjTjRSoSdrc3mhz6CD5xtvTVY8XvoBDQDFlvQvRzT6WO1vjtaH5SQ
2lqkMQHdkWorf85U2xQ+M+J/snjnCRfgap8qa4SwBvdDmoaoN252xVHpGDvqqYjsVlfElxaJ63yg
gDZJASf8Dy8T+h9CidSLnZZvnepDhXua3tBkShtTkFbyi82K86jXPB5AzurRSkl1bDgoclWvpp0n
8FzDreebglIXviUfzLmalgzs7F7cg4EoxFps39I6ospnyaLEy7G0jGzeYmuuv/iJpHpeiiu9w6fz
WozkHru1wOHQ4gXw4kGmfI903XxknZj2nGPraaJ9MFUiuZs0yUhy9TA9fqJfDoDqIGYLA8bvwzKZ
lHPtN5HRLhbWdBJBqBjrq6p56HzTj/PPIHWDYRImp77OUnlRLcddwSV5U41LbQrUZxBXY+1gY0Df
7vYm2quk5xxYnR+q43+93S09/8PchizxQlrDwMFXpggjWx2QK18lYKYJvHsQuG4+LL3zqGB9hDOM
0rqkCBnBfAmDXpJ6LE92xgFlFVSOj/BTViI4tftJ1K5UQFQjhjpHHRNTzd8hajYNZHyb7xPFZckP
36JIRq4FQWCIiIaRJdl56Ygr2Rf/2J/tTpl5/e2cet/q1Br57lK99sGXkHpvCII/Va7ITEe+th2r
lP7BXHMUiCxduC6YGA4hYvsZ2BarRNtgB+0Ns+dJUzZMEHr1phtDcpHwztffYuMm1hscyT8xp5vU
Qo3GdPzztFvb0gWqurgAQ8qJXivw5jCFvoY/GCEdkWQOxHqPWfmAOr2siTHI/p2kG8Dsb3c0ll35
A2vWwikTbLXhgU56qyOtnBXNkSWug7uKrcm35Vkf66WMupkhdtd8qJP+t7zIYqxneIThxHlCF+1h
rWJVNPuSCwlmTftD/69IR1wlaIL7BbbkNGOxiWivzw7aGCviokIxmplB/pcrv6xiyoGxfw6fFfw5
2jwEp78SCy6cvnX3tjw1kBA/O/1LtukAu+eJ8Y/IIkwAqYok+2BEXdPiqynjKp0AHCLq2gIeZQjz
fE+YSdMC33YIiZDuTsTQrniRW0q4BwRlCllgpD44SKvQWXpfpUF90OxzBC1rC/HENhXpLrPzmOie
tn1/aDe2VSXfR4Gyal5+mVq0U0P7FGXe04yL8BoWzoSp6qc5e5HRBlnIRluKu7PZX5fdnfDY+33z
jG/uSmJA5NK6Lyh0IJD+CZoIc54E0ZdAl04RfHvNqr2+Qr1SZejcaHjBMMOMIk6jEErLxsBAAmFO
jj7zuJ+xfD56UfScypUNkY/FU6kE5bTpwRS9Wanh0zF96XHPHzdduJEUvmYL9Vki8OSnZEE6ik1e
VgkD3g80WxYgvGSf3ZABaocEsn6oMwDpUacwaAX7s56KKpTsap2xoA9Znx+51SDXC6Bzd+WKLJVp
6v6X5ObJplSB9/We7OUIjxxFUa9AFO7x1SlC1xjpXXBK6n7SMiHuRc0rXDb4fCH+Nx+w3alDDwMF
cT82OHmMa/MB3poIhUg/p54AeRyAm4kbDT7K6zca9TVQKQXu4nus6hu9X0KF7hWs79Jb2RLJKuYd
wCwRPrhhGC2Ej9ODDaYAIAZrfLwhN6gdG4pWXr4st0AyTiSnTVP38x9ss7yjag553dIgWR6icxQe
yTs7TmFHhSpAHOgdHps31DUwIYxXyXFKiDRnJFOMVI/0zU/eUzc1hKm5lqU811x7JdgjhoDly6Lr
ddI/rRtDvP1nliBGtlCiunJBK8X0UQ/s8getU5TMOBig5U176EFYaeRIxip70KfoYLy7nsSZzQC9
M+7CDhduQh4h/yOp+oVjRl5CsZeTeiGB2c1xOrVD4hAI3v7pBEan66BYYKmrwFAioiDRBb4xxk+i
o4dcrD4IBiGRHDbrjJUQHocRZrNo1mFFqiOUWLyIk3/OZYCPA0AKBTahaTdSvxapyc4ObzBThkwP
UPOhZUjNtrS2Vg1w+CBdg+UnTZfiwM8SobE5W/jYxafgoMVm4hH37xlK1F33LCZwgk1AjfKWlkwL
5IGelAcX2MxmcpkDKGDwfNiGSg69CQ9moPC2+nvIW0d9Aqq3z3OhGKmqM3OapyHoSZ8dwnMTc8Rr
ZVVCSzNFZTZa8pmcPvZFP9gGVzS0guf4EcpVW88lLnxwROEBi6v1Npg0Ber8FLvmDwpLJgug7pEC
kTTeIZ2iLkCzmNkEyZrt2bKvLp4RihOQ1ZFezCuKDnzdJvucYnFkNmmEZKPWp3cXtU9jG57ogz3H
qUCdo9IPBa9jllYE7Luc53Nca4BDl5mzOMLSEphwVP4adR0WbjV6Rb/jHaH/5EVZU19gwloZfO+F
d6pR7WxNeNDcPo6X0M47R8/SMOHqfK4Wgp5p8u3Ur+0QO/A5HeO0CXo+Elfmrn5gzTK66Jxc6/A8
Fixc8TVNnzs0krqVPSmVVf1ji/AWeOa4Zvti5end9te5Uaj462eg309KELEI8Bi8S9N8zv2rW6f1
ZoPfTyW59Rct0P29/a6L/jSfrjFCAQMjyPBAcjKZnhvjC/VeaqPExXo3LUSzeRo43oelo5ciiQsS
3nZtdV0YDeVT3C5Ld0qnCtcL77PjbgC01CV2baG2d6GR+hmWcR4ip1U6MAHcwQpq1JMoMZx+WC98
hEI8sf3unBPo7byQAbtKQ0j6K3jJFxhLLgYx54tfaKel+6NVhyFQARddK9TRFT1Nl5CmTYggrQa6
38fLxLtAcbqLrXquWqylj9KfBgpCFS+M6rfEIz33rR3AcskAytjvMCjOLo96ZBa8d69ZLWbAn9GZ
KiwzKhWURLa/JlJQZlY1lXJQ/RCnSxfgX9LVgB6rpTkXsS+fyy/qglJ4t9zoQRBG21kJQdF/lu9K
GHNCEjWwhIoHXE2jwrExZNp7Urv/sY4LEhlfyjdiFAEvh8t1RDPTpzYFWBllCHlbTH1jgmJhEpys
5nuZA9CLMrO2U8prUYo7R8nfIrkTtCNkR44NXRQ3qzBho7vLaHBHfRVAvO9sTXPXC8cBGdweM3Pa
nrV8sS8pt18bB5XofFkQg0bacgrRfANimFdWg7BePtl1R48vZRNvnctIx5pfWzQkDdH/wGcpmRnx
Vn7hly4jBTr5e0uH9Y0NTuk/P8+0zUXfmf1rPkXgWmnQMf7qq7HGAXVHK9VfvQ4IucfR9s0wIPFJ
7gI48X019uyffotXxqlPDIZ/KZZ1g/JbAs4GvgcTcPovcyuIsb6ZwkySJkUcHg9HVdEoP/6P8++1
oNSuCsMYMsL2jkzyebdzEs5X5+SRQhcmTxc8osfMDGFigxy8B57BNEG3K4YbkQfu3OX5KpvhgXEZ
Xiy5qSv9sMtvpfEyt3MKJCLG1q0ptiAfgU26uyPtyc4ZfllW4CIckLBiiUlrrGpvNksYU2oGJOQH
bnyvY3JInZCIV75jb0JXuj1aMNX7e2+DfjGS8aOmcriPNWTfpTSfkzkKphQoEi1GF5gPcv7GGV76
G2k6CPBcsAQMgFfGAc2BM0w+w9SSHYdcfpPkP5T465BwiC9KK8yAJEzfEhzG9x7fR9EUNa+OOHAw
i+wdaToYgos00Uzza++iGhlosdIDQkJ4zDhtCsGglf0ScvchyfFtzmd9zOP0XDTo30D9UzyyM+wC
CqMytc8K/yPy+L4/41+A6FAm27vCqhH8AQ80dAiXWbEjZHRoQxb2m2cpVrKzOHTQOwZhFjxl5NL3
RayVZerOhUaZkalV52PMvneZKKs5jhWT8wS9VmSwEGlvOSqGe+KsZAX8rkfRl5X/B68xY/0ghqzp
/+Efzj5q/EwHZEt6Q/lR7EqC9L1xJ7mUN48635BZbVeCS0b2kSV13mcXczYI5xflwJ5m4kc9yRP4
f7YEYLEDIhUtXmmFVTaYBu6zAbdAb6LP6RBkDZdbo66gTB9wu5qm3/QcedqvCjWvvBw7l3Kq3EX+
Cm2PzCQDpdk8qqJ+spYdzokzwSmCyYdZEzVY66B2Qq0R9LgMhTtSMjP+qQ5Mylxxt33eDM6Bnhw9
2TmBaSKyLqlrH42LiO7AXP07H9ImxsOImKSO8/SNxXYVVzPlOHtOX3/KjRThXe4tv8gqqN7RU2IJ
0L5Wlon7JzovsTN454WPwnvrQJXmmi9k0zIbDNhHeKbrzXyezRT0d21QgjeTVp9NYROSck4vyMzo
THiYdGbwB3s3FhUXLqA8YqZP8ypgCrqCsYRpsTlyDkKFnYqBuxqMHGb/r09K2UOXLdgWkUJim2zU
lod51Ve3o8rbFOuxyKTk6770dLvTPJfi4ot3g1gEjSB9fkR212w1wKFXzoBku4PW3AMGvSMTNJNp
BSU6B1Ryp8QDvo9RiC3FTzcIYogqVXG4HnaWcO3iXMRPgrRFISAsUPKNoLFzGyzIP+E2jh7cAoqp
qzFuyaOlKB/anM0SZKw9XTaaTt0qxKtFyoXbjNeL53uJCaGTdCHULJHSUqbgUwjvFwgVpw2J+d8X
JInpjEsAzxBCnKF5ZSytHad5QzH+2xDUWT1wN0rea2/q/miASP0nirxeGX5gPBi+9UaF6tb5aFMk
sjoJMiuqI9TllF/9jSTdRmmLwv3pNL7lq0EUx/kfWPrY6INyRXu8Q44LRnHaHAz1aIBnJv5PlVcQ
Vm9KNdUbOPgX/LplIhR0JTMBBF2+zbwO+tTWJp/LZnCbvDZOm498cpLTtoXG5bumfA15sE4rDDPJ
pg7BWK6/8OLFlKmsZvCL6wMBSQh6Z4QYRW71gX+h5Zi+f42joToYYy2SwEfNvCK0YVK65pxoSZdZ
gcm1P3kz66BeC085c0csQ6FQb1j80FSQSGEubXDhNcKhoBuCKV4uBTlxU6wV3J5/YhOHC60TZan0
Q11stZSbY/rCPEi2EZcR1zpTxxa9V3aF1yP23erfWj7xG5GY4iPtZ8teBfEpKsapBEjUDjmzEyCv
P7yq7kScDhlr2GmNdJmglh+Yw2+/JW56xMLUSoYpDTlYpvVOZGX8upYV/cZCh3Jq3aCRIPi154OH
PZQ3ZirxeMXZ2+Han2pqd0DnNybmqAtPCbB8qoKH0hKi3wOjE63A2Qs9Fll71mcV058xeisTIvfb
I1sCVeIw/j2iJimKfA6v+0xm92J/J9MJnh/OZLugoLDtoRxmRP181y9ZVzRA3T/jegTEtr8dJvTY
EiN3cZ4uihRtEwfEhKpsgQem+b8FnK1s0JcYtfP8WJ01omBl5Cvkb37uscqQZuo4Cxy0BUaln7S2
+gabZfbVoq2K2L/863cP/egTRei8lGuYjALbe0mGfXBxxk8chYuiuoxPthBRlJ0E/7LXUNGWxBGd
RWVYWqnScNGR2vAYh34dqtURWyJeXJeUgSM7ONczTnAyVmk3okhDTZZom7v7qR3IwxAaFXgwemFP
bPphgF6bTbGpRihh9rQ+oM69zVjrhFhhTkJqdbjhd8VRQCGYrqiT1vOohqvRXo5HRGn6E389nnpl
+AwNfFPb8nWcYMehRCVJU6Gcrg5l9a+RdC7MGFlC2B+hh61Xj5LBiAJK8jfMUe2AUjRemFvHqsu8
JC6U4LGMQs3uEp6dRb474VPKFhRTfooK4NsU3n4+7bNvjKtco/pXBTEX1iRIFt1aq30GYrUGZYt/
U+YPJzGnoxhXsOKDLOhxRpYPedVzhEkNj+DIaCukXPTJBA0ylL0eItjCDBzkf1TmKx+9HR0mT78u
yXrTV8S2Nidbixa6hqhWOqEFYrw380beZzo6oQeu1naO1sx85zp2hKZDI2vhduixok7672o9Rwm1
AkDu7XGIOWjnFxRZSdbqK9djMsGZBtYaE6bwSNZ2VGyev1z1u/tevUl8KQDwNcsKz0CP4E/FbZCO
Rmc/jDA/XqSDJFbNRxILobzHiM5KfqZYzjF0eaX4Eg4k4aBkiTKU3Ig+owLGncdL6bXbC1mfVI9C
PiQg+jXvJu8chJsN732JKt+HlhzTh52Tp7ohtjwlg2Agi+5FjityWo9l9l4SKIgtYJ2raxE42rRp
m5j3gJ1eDH2xBTrWneKEb6pX3V3qRtk01uI++Oo/dBI4HYMsG9DgfaVd5GXFjpFlWDCIQ7U3AG4J
x9Dw362D+xJsP0IMHKKZFICiToe9UjKgWyIzEs2VnOdXdJukwzo3NtdbPvdhR3xkYj9+RYJfLBIj
oQZWkEjx+XOQDM4Sl0yHe9a5HsN/6GXpvAqzro7VrAh71GvHQaEGaa1twgR8hWVa32EcJnASGw/D
ga3jLBH4t79U07Crf8P1iVboiDe/UXpTUeO0kgZDTv6bf/jWUSc6eMDV4qdn8oLw7p6laZUDtzTT
y9/f26KUpQW1KnuMAZuHt0Ze0EoxLvUBqv80EzabuysGrSBs7sRmDZJ0AOl1Mg/fzZ4n0SrToVIA
tzX7THBfprr248EtAU4EbKxQ4TErqGV8nnPiDa82kTnxFZ2wLLVMuOj4FDT8at+a8uL2WqLatd+a
saWM49DEsnRRZ8p65Kaw2XJPIPJt3QopNYrDaajZq1Rxrq+Xc2neqHTIDvuaY4mAKdnM8tB6jxFw
6XjfDJsEDSVYz1X/BzwrpLtC+D1onY0aWx4grD/RN588+abz7vyqS+gwQdrTMf8ZpqOZJqnkHYdf
9sb17ZLzCvbQhfv9D0a6uAzUukW4R2ibr+57COAw/EmkblMO9WB61zho7vDxth8TYfQ6HVdFc+CD
WbrE5T0eXqencXGkmm7Neo5bus/JyiG7Al4nfBkI9bzKNh90catMUslabcP3CgHWhuU0RI2aplI0
7AXDcwOhrCciWXIUSf7sShuYInSnii/fmD1oo8kDJmmWsFcF8FZ5ZzfIBV4Xo9t6RTHckvh4jwGa
r3PpZq+ag0XF80MgCiVfp7L7PNiEHdkshSqIkRVDvMZa9sEESbfvwW/Csx0HcdIeW9J39ijpVV4g
CDLA/XOAfnxvk2Q/k/+QHxbDOLh7+S+KXIsH/ujJ/Q98ZZtgJbm1SgCt7ysRiCfY1OS766bUikmf
vBvlXf8UpTyRd4IpIGwtwUNlXt8dBKNGUkT3n8mlOTaz78MGG10n8eEtlOtVcT0emjkNbr6Xc5U2
u5k+AmjlXS1RFl7ZlE7+GJ9tbaXLyA+SdIQEJopG1nqoPkP7emYAA7/mNfSvObkan1Cjin3sEPn2
qsOZkQL5nVwRzuBsW5sPVnPdTG0Ks1RQDGDJ4Xzf3hS2HisEKGopEfQ/jyX1S2jvGxpqxSVQcMJ3
NKDFuLDSTtSXabPtVcOZzWvQTUIzKqrqZRPPmV+z+HCnoq+42+wOVOHfHnuCt0gZSoWgGt5+xDZM
Ob4gY0Ahi3RN0mtyLH1Whxpig0woWrLRH6A/LZ3nf2FjCIZUc4vo06LSs899Dz3eYcPYGh1MtmXQ
XvjWDgCVEpM6hFNYlx97VKWdCFoSys1613eI+qVXnTvKV1oKIpTjzJUAWTfh3oMVATNF8AxJpc0m
eoSWtZ+LHZG/tVlp0f4z/3JvjhqSj5DR5YsYjFTL0IW8voRVRgqPfuFwudGDHnCAsAVmFWDYP14X
SrigH71neN4Z+cEJdwGparnHH7Ldv6eixpktWhYV5sxH+A6gO29GVDT3kPKdanq/urPW5P14eQIl
pPYL5Je+KlgxMiiWMgByP6ik0Pkq876OjvXCuVtCQC5Z+nTiLNxdOtJdj4dIQxSTFwz/V6w8Fgi3
bz5OIRPyVNj4btlqidPUW3kyAAZ/kBA4lgsreoV89FRb/1HW6kTY977uIsgv+moSkUFxHh41hMUy
oLzwGAjqIfQSHch0qZ7KPWliTwtgmh1BvDYAuHjOF6NA24MX1jLUc/IKqgRUv4kosv7oTCwWnr7h
6y4n7HtLaRUFbd9AmBFzHoNeE+593H3eeCcmtnJCuHQTWKpnTaBTP+bsanqJXO8HLtNBF+3l1OPk
MJ97cJuhhiFiMUTMLRfcJTuVLYElHacLz0MefeYB0GgrmIwTcNIXGXHjLfndfAHfWaNcrE6tbKpR
4a7cjHcnMOu3DnYlIle3/wJSiKbx9hlDwMBcONX3dcw2NQ9xLaGWkUkIqeol+HiAAI8JBdYIre8y
xIe8bqHoTjDJwgUjauUX3BAvsSjZN5+KEXT2AQ8QIwCO50pn/rT6RNg65G5jfSVNO2fcVeYp6FJi
4RIjRqrhPG7xgaa/z+8Q521WsD7yTN96MLTQtUQ+qR1VFBijYM5IOJa9vgmhVDi+TRAoW6zQXlAp
O7tQy0LtnufKhjp1OXA0NuS6eeH+KkgsCwdTshm+DUWkfYHKNvBCdTJF+0FUyciRHsCxdZHs//eS
D+zhElbbYiOhR+/xlMuKb9/DTadq6RPOkqFwZGURzsu3Ju+RToiZxX6sj2SHLY0YRLcED5JEpU++
NX9yd2WPRQQPqb2wCmXbZAkCdbLNVzb1qyzwgZSP/dBWDpdqIewrrMMzhe7QIKU0yn3VxgpgGs0n
zHrpIMTA4AHjlLwE3RTaLgg9xLd3nLVvWfB0NrTBRXJIk+CDzW+1ljbhaMQZRsjWUQetIEx7aCUP
Gn7QtYM2WFFS8dqIlfIuJmhiuzVEg1hBev1LBIzquBPut+FIblXz5rv7H0r7PFmFqDFmj1o1FQE1
lCcMItkLMHGkaHkkNfkRLGz+jlN2WwZj2sxI+nwxdXErK1xY4EktJIpo02YIDZbgrepjeA7vUJtI
WWzUnZKFHphoJ1cUNJEqkTSvRpzcF7ggMgoSHwMIGvivPAMjKnT/fxDHZ8XT9J3Vy8nV+WLtbk2h
UTADL8U5FBRkS49DWcDwQiFMR4q+BcoTRUwyhployeEi2EEi5wWsBLbqHEAEyk+iLotQkSv5AGfR
BEqUEu1AX5dxdNx6uYFmCxygh5m83bkOeNHz3ARsES2sGfOeCB4yK7sxopnZ3sGkhCjkST1myMuJ
V4zyFJ/5oKw9JAV82SbLfEtmaRPnpNaNN5JDiaK5TNmxWfijAdUDMODauOuNxuEDB7KvqPiKxIkw
k8eyKmVK2Vd3k/yi4xisqWZ7cAVnQqC13g+WTIM39/wc0wj/cU3w0maNCFyvjVSfXtcz9ltUcOhI
SQJ8zu1B8e4e9tJLD2Xw83t9ppjpuh/04/iMpt/5gC9LdBxlz4xodOr5MCS5liH/sWZOk1o3tVz0
a8pEohQcAP41kQG/4GKX6VUnFexAya1WmaZA8puT87XsQenXI+bqaS7adyzXLPw+qQ7HKLqQEpVa
6HDacicNIvetYOrP3p0Ts+M2SF/+jsc/XoV8Uo8lpFY7NZJVB4YI/LpBnWjyvJuqVifCDdiPsOwA
DhJczcN6ZH44LImEPGwU+dgi/5hFSH0P7qMtDXomEFVH6TPBw/rpP1xVhpGRuNQQxrmRvwipZN4t
ZevecS3l1vAoH3eqM6YwTbeQPDfut2MQ8UUR7oDUkIjhok/uvoEofIDC6hsa7n2JfP8tWPjJ2m+7
LVcbg9sypBlj+cMepcOJjA4Yh2gUGgcigvVQQ4VexG9Q7dxnQMEGQwON0G4+AMOHi+WHP8HjhnPh
LmIV+XE8THjTJmDZCZqD+8KJFw1LujQFAY4z0+U1yvak4LMmfGvlgi+6pzwu+8zNNLcxS2UdeBqp
TfvEDx9eZPTRfwSkLMXSqiVaIqRuOv+WmkSHrREhzyyLZYNgN/92/W8r7DbmxXd+cj+RX6PeK2sg
apNSKfUX/ajDgL3rB7msTGaC7vo5S1ZrwAWb3I8PBaHUbByv0nYrrVZoi6a6lM7MC6UY0ehHOreM
QjRC2LI7aIYcV68cyiI/7RiqDezgU6L4jXUjhM/6cyXalcMupcj5w6gs3PAz5sSfIJkMxFS6YaNP
acvdd7L4+w2eKtf9jmviTvJbcKo8weMAz2GuvZQAzAftpJPu70H88Vu3dv0RupsLOwmZ+5uAkLZs
Gexy5wop3IwSqh1+xlHVkCowo8am1bTeBAJxMGO7/fqd4AX+i0ed1SV38Lah1ie46ABTSCQngcOe
MUSePZvnasdSCkZ0A3nKfP/xOA387BLYGBeDrlBSWwnGFVBVZFOYDMaGdX5VT9EMh/sMXuqlhDXK
7ViaB2IX98cqArrhZpfW6qSaBzOM5t/y/bhegkbLAjaqLPAOrNBFy+tjyUFsPpfvf6AMRxbO+X6w
nqzu8Ro8F4sGYE0LiREtcnqvznmocIz1eBShLL67P3vNuV4orBQE0w4hJUXL9H+ne4JIml1UmjmN
F7oqx0hiQkcakUoHn6gqQt4DRc5QlkZcD+q7nuNmQyF1nZTDTFcNakZOLTuldyPBzIKzFMNa44Ya
Zqs/clR7+VrWApIpvK/EZ/GS8Tz/mektUy5cZg/gUoYHGqHkEHfX+dnO6yt8T2ANI6ik6714qLVe
FkJsM3PYzObrICFCBsX7Yr4lTDmYA6SuqBnlZJBTCZXO68juuPLA4oTFT2vtSXl8izp0RteeJGRm
0T3CV0Ohi+6hmxd72mW+kM4rfZ7m0XbgcvS1uikLz/eRQ84Jd+kbVCi9fhJUfQwX+Knijb6F+NrA
R6Z4ghZZV61Lhgn/NKynY0gQNjSf7nB4DORENWRTrz48Fi+A0BZpfNXYqbDoTN/8AVZZIcxwFOhg
UK0qB2H+b59DtuKzT4aukiUW67T6Jy1AkAhU+xxlDgyE8fynzGPOXsmb6jc/4PEjsTm33eAGQ0ny
cGPSEOLxvBqeggiNLwi84Yl4dSmpH/+AI6gOeY3VE/TfD73cM02mLP4mnq+KUYR0naBKUonS6LG8
b8M9BTansFOoVRr3+tFo4ak0Cue+FnPzPTlJP1p4gwOqU/sn2ht2oe6heugfU7dXLrxrOxUgrVbQ
CW0J2+zylHTbm9ElUIvs2Ixf4kGfYFmakK6aeOKI2iCqUZf6lf4QBntUQOnclpwvrfZLqFjF3DXz
7pPHetM1FTfTM9Ap4b9s38GNTOB48gibl4VJ+035/fjOAOMO1FA95R7VdTELwYk+sPTLmN2mF7vQ
ixeuxhd6BeLIEsviEktaUHT3R8oI0hBQG+ZmNGTSdGSD9tRchBbP2ywZvxiOa2fSqgiDzF/ZusKh
1stED4RlARD/ssdKdWu1AHTgWaxvl6cv3rXCCRqlwmQAr0FE2s37DqTcSmAp4fs7iDzin5rGp+sN
L48hggz6ouhGytE/GHn2rsZgj5afQG33Y1vABenscCrvxLBHq/SSTy9xutCXUrNrg3YrOL4SPbtH
LUN7OzKrfCOLAs5YZmpvfIAAsnYbBNlYUdETzf7lJUS43pWmjaBBT47Dp78H1w97lOrzoshpQbip
VJXiOxtI6pffmaQ/VLvl7RHbvjxS6Mt6a8yL4yYytin36spVFP4/uDLglGfp1xOGzAH7Tr9/HlF7
vz57qNDYS2860PoSGAm0qcYDWnoxTjRbzBnBovJfA2JxYukEfpV/iUu5E5W7V5FMBmZXQM0fVW4r
FWKENUEq8qf/q65yJ19jnXKlF6GRPFTMhqgdFQ5mE8bUqoUXNgPwkIOE6KAUXsZnOTKhkvsFCL1D
BiPF7Etbb3LV07kGEx0xjgnKFtd1enjHVV6AuN0NAG2XA3eNhtN3fqvc6DfPBLuoolYf8vB3yf77
FBX1J1/n9LD+o9iBhMN3t62MT7c7TEqqdz5Gdf3e1f6/WUjtK2p5VOzm0IlkuJYgP5V+0sV3a5++
DuSJ5wg/TvstiZlUU80iU7Z2eOnjlbxmmbDcyagrOVxKg1kktKm2Pvinr7MEmmOFlkcsH9RQV9f3
wwZ8JYGp4aOxOd+LO4BI0EBk7rkosCDWYLp5lXLvifaPLSkG7l0XVzWgOAzgaRtzu7HwHsuxTa4S
N90fqasbQI4Fict4i9ZhqA0ST0uD6OIwm4nW2DId60joYWvxGAUYLDHeplJO99Sa/P9HG/b1GG17
Q6x+iD9OVFqM1wwtF1tvhMgIIkehNT/cQIwDQ0NpPObTg/lgHREspXKNxG/anydntmeYwYehFeZX
tkiAdDVOZ88Nel+wV3lBUHCBk+Il7htrPdvi9kj77DAl8Afy+yuD354DSlbTiMHfukD8rk0UlW5k
NLRfrO5mg4tlL0va6yoCojQ8GOwg/TjiMxxzf6ppAYjZmKhpUXwuBSGZ1AS3iA9w04V5pqLYd6DI
Vic+oF0fA/xZjbBL2yNRXg+baoCLSStpy8rsiA7fGD1zfQy+MOTwxI/3ztLZJsWdZLLSXed6KZBM
pvXaidHFYUlGTdgjd/l5BzOcMMi6TZFfUA0mUdC4l0+jJvGpomquz4gcCjsWVoafjetFXsOYkylb
7JqT1IoxxRTcflMmQn76Zrn+wHOnA71CdHpDND09iVYWjWjbRM0KvFaqz6GC0TZx5lqd8V4xWLaa
+kpBvM0ys0GUdgxYU4Eb772Q2h+d8w24GgzKpgAIzAo4XdU9BS8qEc5J56nfimGu33MecFIAPWA2
Tir6jXoa5bHEifPXe5nDX1wqwB3b/rMn3OJ3TpzmLVxOf/RlyBF0pdLS50UzYKlqa4/5UpbRAgnK
N/guAj0ExIBg6ydBMUlfWHhj+nI2Q5x5OoqfFKhz+lJLSCR551kwAYOXVc0AHHfwNRYGHLf3UJn/
M9sBirCLlRhsQKHRMY1LT4bTik+3TjWgVHZKBSRngFj9v/aLbUWaNLh/hMGtCpzYA4UTNJqyRIAy
XSRqswayxDIMzTPLvvB4u03NNsoCN+vWP4xgWEQRH3b/ZQNQojFd7haXWsS+CxttN0T+yzSRoCL4
/2OpqvE29wWay1ipeaaPT21gW23TD7/lEaOH223e4XhRpm80FKLKWPLnKZKGeA7rD/iWef0CvDn8
1ErXEWgrNx8gTHEKo2s4NXfgCof599xJKcPlJDz+PcDV2kiiooPSMg+ml1QtQnRzKFbO7k4HPllW
+TCEmpPfaKfkWKINV9sp/S6VA5nOulxvocv4HQYSz+EF+op7c43RNUmY2yNI90VYWgKKoNUyFRuj
nU8bKzYb5Ls54ugsjCSGV4TEGqpbDr/659ECk9dp7aatNwSJ+zsVdqqDy86Y2rzeSCYU5YZ6xuPO
5GJiEYHvezdOGC0Y2Q3dJTRqdBYC+d+V9KpE7atYXI27P4kd9xK381i1ua0R3O1FO2kFk/8TCszV
wors9RV6+Vr59Elc9E6PeA4LE5CQxiR12PnK6k/S1Ve9OPwBwl8O6ua8FohnAfXAa1Ia7QXxhRVe
Ufz5bSlOATt51A2S5WRVj7KMpBKJx9e5ot0HW5YG87zxgwIGS0xxmlllVCPo+jSbSgUPdDuqF8hv
rwFQ5oZc98CY/NPDb1YJkuWs5HhQos9DVzd39NV1kSG5dEOr8B5dEyQAkqYvqKb0Pc2u18jyl3PF
pK+EMr2Ry1GIcI43KFm0Hi/2ZbHvrK1FGk0Yr64CiMGsBYCFKKgols94lASWGYX3iAGZWYEp/5hb
5bNUONQ9w8oZwY5om2u8plmGLwo9gtLZhWOHgHmJsF+mztQGYhFbSceOdRbyg4JEyJUVpmbPO1o5
OmoruI/tDhl1R5yzjuZC6xUSAR9aaCrO1vSKUTTuCpyAsVbIcJxFzZ2DijSrZ6THstxrVFc8XaFm
FAqgDRUZq2GTD+16VIvMSnjW6x7wHjFIEYElCjRK4liYSvJAmdv+6qh35iV3Rlx2uTNiKeS4Q0xE
UFTewX1310EYRQDDf9fWd6Z/FZ0d0Wlzmn/SAE71DK3v5IDEt6ncYDdtnj+FSUIyraK0UAkU27RR
FykgsJmUzhXWk4LsGqUsmSezJTjAxd8TbO6D9mJi3X7NsJvXp2+g5ZfHbuwLvl9WY/Mrp2QMS0WL
g3rB9PhVLXxg2B5hMb8TsH5Wn7enG5y36GovdBfx8FqKf147w3Ec56+NOJa4e+/YtRF/+K66giBo
KTOKAhw7YsXMkasv/bIcCTorR4MoF3m9LFlgaQ+3gN4nagsWetShd2rwgzNmDTpkNTWE/XjESEje
4u3Pm3ksqUEtF1fjosJ3HLOzW6j76U2g3pz1m7u8DD2Tz9hzm67+6jxQP5UAnL/IIKERGd+uGsUg
TUkWRglyjkF/20dT6icj1qpENM+zk8SL/jW4SpE1GvlZDs9pAt2mj7ky+pxL1hKf72G3Koky1PN8
SwwCo3vMazNaxWOJlfQay56jDUUiDTdLKzouBhtHTVxzNzM2h0hAfPWhtSARuaiLRmoLWw0Z3V1S
CbzF5qgptCZmenwnONp12ILIljmRgZHNnuKraFACxQiqN2VfhzJqzVqoG2U7tQCShBhwBIQ6rzqP
yN1R03ux8wLoDEWvkG4P4cv1LaIjNobmdKZgBwVwob+0bu2B2Wd8JggH1gLrKo9eX/H46seSvJ0q
47bUB07blSASIXsJnf65hv/HupN5JXotnI/eNVQ2GOLiBd9AY4leNuPN4u13CWxH4/Pl/1Q/emPo
DFfRsoug98k0wKTYDxYSTPeGouW0uVoPrBXzY1EK3fjFFAOZVFB8cKAyhel/THgqYMYJlot6LIhU
ywHHfvgHQ2kxSID4zsT84kwz+XJbTgVtoIQc8KnEFumffU5Cy70gZWK2hMmJvF6SfA11MpUCcCAi
P+pJUq+hbH5QbajEgLe6jHJBxGZmO9fDA4J2BczlBV70S6W9zx5PtWh/1bSxZqJ7+FvGy/BV3T6y
5M0ONxP8BVRjF2d6C+oBp38/2WwWDfvZ7u9vR+Zui1YWR3b5ojwYyX4UXk+hAIOTASkgnzYifW4b
2y3Ps1//1kyK0Uf360whmlPFNIKJ4N6yBeUxnFHqzIfgXn/6Py4aK3mtJECNjPHXxy9+GeNYi7gL
34tPuXk141mHAIqwTAnBitEWEPG5ST7HgB7oJl4tyZnBQQVHkOGdh3gtiY5qv2JM5flFfxhpFzRR
uT5Fh12g7cvDBwaOAm4SsnmR5mPdVkhxkMSv52xGUd+qpAbunWkm5m8ni8+A0Rg8GzStKvunjpLr
9wXwXR0igJ6oBY+Xw6h/ZhE5tDp1L1KxxS6P2O1RWyiNULmWa0zGz18g7U2g1g9NNjvecJAXyeFJ
oykXCIW5fjhdJMDvJqo3kPT7vAxHQTmrrR65LEHWfi2TGVQbAMKt+ukd9/loPMhSd26/tDoG8FPf
lni3rofr9LAzSQQumuVDuD4dalqVCOXty/jFqJkBZzgrHGbpDtTMuNyBl4InCwP0gfQrwdjIRy/x
Tj0ZMJHtataPUCnJyeboJRFYSKDMWmUjg6J+T4Wuw43I1nha6xXFag9deC0XqBnMOEmSAD7QciLj
hp8emSiDxhcjy7A2i5BQLMESc5JgrA2DA8tIXDHBmw9f0NxwdhZ7I9dxOd9JAAj1wdvDmlnsYRQv
y5IjfWJ4SN4gXjykItmilysHarldaBK4HGe4ljfJh6HXGIXF9PFl/ApWHo0duXYsHWe+rHiVLycU
Va1XuoGpmL0xOT9P18k/rz+g384tjz4tYXBYRVwzt1DWW/8mP2HrpEvp3f3A9ITGPxOOAwKkXaXl
3eMuoEd0hMqeWEolHBSO15BtFz58S+FOK0Wh2SD0U8jmlJRt9mm0PysaNCTrNZix8e78k3CRBgPR
UTJ1oQXqZCgrbw7pplN8Bz0yGTCMQE8IbStw4xeYmtGBR6qITdanK4Gtk58vH6CKMEVW57CtzqGZ
oaqlu5QXk/TKni3Pdt5wFZecvei8J7BPTKGyaTxZJyaiI1HPP1/UBrG4aa0pyU4RmMhcdaWmX5M3
bZsfeikj9dBWyy/wnkmOY9btqxgzj7YvbEoEMK8aZAHB7a8QBrNbQqmRi8KjWTtF0JLeq5niudSE
XwfuVi6V+2D43BlmbPecL5FLRm8xeBqmgz5zNLrf9jXhQp2WnopALavCG1m6vDIsRKkvpeJntClG
/uP9+DXX0cTtg8D9XOrdstLJIAyRMpFzaw9aUPcW8Xv7TAlIwnwcwmoYHFtLDQr7o9pG8OmRRqGE
bmMeQBQxYQ2WNNfh4m21Y4WO73e0thrGkgK+b6UFMLG+fkCLpWQxjbzp1jJ/+VdzAmEVwsgJKXdK
NvdyHsRSgf3y/09PKUryVgrDE5IYxmwGPB6U4B3GTFaWWwxRFFiCe+3nmadpbj8an3NdgU+/D0Ce
AQ9Zro4s50HxgebEaTmS05sEnry9DWdzPlivWh/bGQggCoHMGCtzkZxJVikD8eeBeLZDRANLxwWa
xATijUXxYV+YW8lJn9x68LTXRfDG9oYpH4bwjfFaHTSOajdP6KzbJThpAXDA/ar0+ofFP6wsQe8d
LtEvKKeg/jZKADl/SQ9atS8Ymq0Ho2ViAjl5W8/DN8LSJHnm5oNs0wlWIwZdF0+Km2MG3+ML6cnq
Ve11QY3o5K4QxpZbGFuiPN8xtecbRH+tdXOVvd5Tf9+0uh6WumGjdk/to+rwggGTgKrsKtpCmfnf
qTyAQ4msTbwQLFvresexvBeZz2CIjhTWm/7edIv2pu7sJSf5prXWLJk1kzZz2OdBWTuaTyy6We79
ywrkbLPI6qsQMcDFrkl6/8HGALWdfN2MoNZSBKqnXcuvlpIQyvWBYhUl/X6DeAcPLKsJwz9Chjaw
2L5gcbzoju3dDFBCUyo+oLKbjU4NQpnhpJIOY71+tECYkCEO9QUVbmzLtwzVaozYwcZvxDJwCHxz
unFYXAcEpt8OyYGAjhGT/QdXFnAa/P4OhUTzPu6gSrdipHKOCv2FCu3oZqLxoNxEPGkQhhn8nQ05
mes2YY7NANsfVFfuRNDX4tGHlIeEe2NzazPxNAUcyHyiYKhOSF5toK8kaSE3pFEZC1FyRQi0qLIj
AKQZwURRX9f8XP6q/OsUP/5Vza8o8s3oHkVz5wWParRtFiBU+U+o6GV+h+oqycmE7S+ZpHRpG/cv
q19Pw3z+N5l/PyuAJVvfRtl+RL1qwQDwwJIfb45hqQ+PqtBE18EgCqpeBKj2Iox9B+RPryiTM8nh
nozvPGIZ8cJxPnxXHP5g1rVkh+MZeAOXnSuczFQUXYsvJNKNXW9iFqPzx2UmX9hlOunIoOcYcRK2
uxms1kfuj3JagWmAYTJGOUuvOHz7Tb53muBjArGh/yoATcHnj9zJ+6OndMy/TJ+SzPJz8S2IXAEq
x36ym10WcAqP292YwwGGvSnJcUK4KXMFJYx0hwcQjpHxTuF2nk5mdgq14XPLY8FaS28UFjB7Q4lr
cCr3uxCvyx/BxVIrlot15ouxSwjPtAPEWM2ieNMLzF8H6Q1LOk4xCuYhNBOODCOn7WXRFooU+udi
JnYESDASLaJknnR9ViJQxJslfxE0Yu14n7jRz0tXYvlE/xg5Py6U8FLb08YnB0od081kF0z8DoII
Th5m5c1PYYA7tTGFaU2jWkuZIJ7sQErcbRP1VFg+hqC801+qAF2Ed+mL8hsuw5wK3C/8jOLkc9HP
EXo24RmXv4HkGDtTmH7qLXPG5kkUBGC44nEuvuVyulvXhTTaKQMXz6iCmx0ShKBTWToddGCq95o4
pplw9ng1G449Np8L+SVxQI4/avggG4PGHXCbwrS+b+6VrkUdP9s9Hnaat4TgL6AOaTr/ePvwBCBN
v7/ltedclvQbgLfBGsXmQsRRA90O92dAdboaoHV01gwaXetWHS91FNVvQNo98yI3gougEQqzaFyQ
lveYI1iO/KozqUmbJes+oNPx0AwNuy3H0yZRWHOWO57tzp0CsIHSAsWcRsYbxXM89nK2pWlJukPD
klh6EvSUgID0Zsj1UK4qMxsKWyHofEaK/dWBBBaBmulOxMQrXkWHvZqjYg4mcz/aPQ0GNzx5Js/j
ZZq/rHx7mqNbeYyBlrOI60LUvQwgiZGlR30r8qLCWh0Fx1PwHt9OJqLYcJhpLCngy9AGQuAEgSrR
wYNF4/a6XgQq552d88KzrzS3JKuN5L6gwUZ2abVfJAAslPTASOApJe/xdpY1tz6EQU0wfr7lItav
6EtgPxCBZCjhi/VsDyN4SwWdo0Nj4PPOGkmxBtW450TjLlQMifOblV7Sa88HIi7RWeiOyzJZyeiF
d9K+hiZLxgp2EZNofSvGHrkpZmKTqymWz9bZ3/RWxSJSYytkP54kzJvSGWKj/NbK2UfKirQQBqtx
JlDq72HNx0GsAxJLj5KWXRyq8Awr1x8akaiw+89PjlcvgsAn/uzANMAECZ9SwQCECNSLalrc3644
BHXh3VXt7zOk3FerR6mUROsJLJLkU28Amhwvkd7gILm9cj2i+D3/d+nocjX/oQFMPzgKtylv/dTW
pveUYy1bT6Uyz65PcVrWJXMbP+eJjToyhYt5mSjcxaoxsw+usLNsN+0YRfTQKXWTUOK12QM3EdxU
sDX/K1P+NucKM/Cz5eTMr7MarWKs4ZY8LM+0qpb0E1yyJ2v86FcdqFzwsBb1AwtmVtCZd4VHUAel
qkXC9ccY8+T/fRJ8GAWPmqHH1BQFc302Hr3zRuGL6nahsjUBEQid7z/Xoi3EtT1Gp49i8yp54Zlx
ESh12iw0aNAjZUqHpS833Axcmrfir1Hegl1gnVyyaq3pW9HGyyDQDGoi3UJFXcT8XOEHQ1xv5hG/
ZqAb+q8pyjkUbI8NGT5bsy5gaI7ivcU5oV5SXiR8y7fr4nH9T093vWTtoSGrJwoBWivx0Y4PV/Zf
yvEIvfsl+z7lAdYEiG8+HQI5NqukANrx6qILAmVME3+PpJhNDlyYnYcl+JVXv/Z1N5R871GQiLLp
J6UmjQtj89/ii0RqgFt4RWeG7pqDnDSlowa1/sIOalrLBncEI55NG9CwiHT6mBg/F6121oC4q61H
hp1zoNeO4Q9Miylhv79dg8FxUIi9S2Atmjnyu5wTfTLZihKO5V/RK2eKrZd4xGzBwJkuip0mwgBw
lMlx+ebGR0JuJZLJA4nfhxNqHjmHjVawl2zEgsWD8QMz08P+vzy9Ua9AzMXkN7Awy0yn+48wRad6
mxrQjRA7utQDRHf1EwvAQrw/61sL7a6mfwCe1IrmcTGYMtOWE1Awuu27qfc1GiF+5Bdv82AY5WOk
JeJWQKliAE7bcy2azd3WsTEglR7onbCBGaS8LYyVF6YyO1OV+EDm60KiTQ48HBvIEfUuQ/ND2uNJ
KunUXePAs0I812X6ykoJqLeIoI7KvHffBt3TYa5HmJdgN9g+2uNXP9KvgIdOVUwbPCj6/pM9Jiq7
73U+xq5GgiuRw2Y78u6u/XhRBASay1y+0T455FRbN5BNAW2P18YKMRTx1NF8cENautNuRsLvaP1g
lkTh5Nrt2oQezSZsQtkm0RrlZuk1Z9uO21k8zum8PuHgPdICoGGcY9z3X1H11wBt+0UxhX9L6pH8
F6YvxQjQd2CWAd4Eat2gTgbZjYYWhSQxiS5sEQ0AAHPrRRrBZoNwnhbJsu4diGSU46kF32j6MFXA
HNTS/o7HCMwcXUKPoa5Yvc06aFZJYZy9/G9pjneWKtnWzuc9inSbP/qtVyoc4nMF3XLkaMiGIoPQ
PghiNeqJ9CZWiL2ix6UWCVnHiXSQHM3HajseHCKzP3m5cwXSJtDG7DGNShzcVoDVcy93Fu0hBY80
6zTEL6yhvJBvXlh3egQ0/m3MUCbWFUq7CJasDRLklFWgUHNS+1uEd1SSkV11PcPx6Lxpf5rs7R6p
HnumtUye/8DTFmmTnvEha0bDUXjywQhI4lBMYtpREsaDMgT2RZmFe1pUG+y58hnofV3zra9X2fXU
ek1Sss6I27UUO6JV9Q8T62SZGLvnJzp8IXsuRLpL2laxzl7BRageMC2KkiNiLb+805qBJF1TQKIY
Vdi8JIhQa5AtxdDDxC2xSFS4iXRl0LwlbnmRkYD5wqAtMdrUBbsx+2EH1sznzUBE/fUrSlZPXTr5
MbyShfDTsgpXXXtn1350u29lJ+8RxzpAEhG5iAN91SWlmo2+aKMLtYvBdcmahCKFUC4orAMTbHLB
F0eBmQyh87ka2/La+Qgc9NKg31MyYC9QsIvDvF3lCsrJc/OOPUKU4yaa8eRSrDoO2kXkuX2YBugq
OLSy4WJ30EjND8xFrByWXZlptNUGNr1JsJtbHLTIKuz+/txS73llqW4uIdaWYKcKWaSaZv+krTck
LRZfcsjXbUDMuv7RyrymlAZLkgS5ezj9ETy1IN0awaiBAjJztqCjzlVOkC7pOKbW0adXnBJvpP1K
MDJoWWwPb3IOOlr2Q+wVy1P0hPaCr4iDL+ImpjVu6bY4sEzpK48ORCfvfVrOHHaueWuaenvtnssX
C43Lff6r9959tRJHi2w3Etv79NuhJVQTUYwL5DHqp9xROSHIdTyj0ocWxaMZnc1mmakXfEicl4jD
/yUi78VqUIwMVIV7y1aposput24fPZSIOqpKQ9qRn70ev5g0ME5gn5pl51cOziPKjwQpD8OTOeXT
P1rcEPBRB+kdCgsw7vRiCQiEYxQksi3Nxopb6aFf16KbZ+cKjFugt//a0bHDlMLy56e6ziMNKLK4
ZCE3aU63y77GzEH8ZH7keJLWb0b5qw/eWXB5bDJzADMVB1XSo40X3WaNu1aafr+vK/Mw37fIpk3h
SQwt1PGnzkmsrWK5SAXvf/VtbzS6xJdl8muALb3Q2QcSU61jAWp+PG1gValB1aZlD5uI/n5gynZm
AC6+2zkTMV0/1OZ2fVcki0NQM9Jm2FNfPmSqevOUqopXxaKnHe2mofiaA4bdJLe+VMGPa4qbXXfp
jCjursWIJRA0ZUyiOy7s8cMdh6G5qfM1V8HwaxAqhiT03fE4WS+Y9b8yzZQYRzjEZTG3XD4DxD5R
Fn6fAKRqmh2TOe45sP3m3fNUXYEvd4m69ZNCgm48qHVDPzRHcQIqZhGVM8I35zb5j04UquCqfAEJ
Zx6ScgA92lIlP7qGwDv9d/MNhfAY6dx+5hZ2J60fWxPKuSpW6D3rKXqXEuv0RqQre/C79HmqSbmu
RJi/dyA2gnf/SP0jW3J+AZMeO6QMjxrRu0f8mukwARezJ+GGohE+T1ULcsjhRZ4hT6t90pNnp6On
mGL6swpViWQQ/XNw5C1OYd0jHo2a+fwVqLKmCg9UX510X0R6AZOc17XeAuvsUWWE1xD7wQtZeP+u
t5S5QA1czHAtqhK/5yI0Hg9Ysmt+wWjRct5DvG1VrpRxJf8m8decO9r5jxuok1EpPuyB3QtbMupP
bQ0dVZAIRl+78WTi4ngv6w25DvjDl2YUBCmcUfUfBD08cttdQZ4mKRQ0FtPNN7SKS4TQc4fPX7aM
ymFs90NuOzq5bFxMb26bwktCOIRkKQsJx1hn/eCsMi/FHZmsvhSD4DYl5YVNKW7vvwa12nhazIT+
n2TGdbjZbr9AKCThDXypFrTXGKo/NGEDBlfTClB9WiyG68KJYcl+XDS1odMDs9UVUHDNxMFZ2XhK
/zpr+DwrYnok7LS5pEZnPITv9HO+sCezOOg1+J1tmv/L1i3BXJ0VIQz6cBIHw7q4YIM4+PVuBhgo
xAJRSOiILyg/bVqI4vLiM8nskBAoD+xLAMkp8TUl+AhWljQjQR2GD412nkJnL7DFNJqLVa5A/EFM
fhCwRcKWqYn06RANs33E9fmSjiBE2fUa3shI7hNdt4b4VPKDOMUEW+b+H56y9kBkmHc6TDhie1ch
LUywjWCtb5mbWqQtX160fSwGKAeIBJijMKD7nJKBU0qHCQPjdKzxfCCQlC7GSla4nsqlJrgLCOm7
GN824Kd7iwsieAlF79+k3orna3mWN5/6WGnTqsOl/eIoHuPUi+vmQZUZPHmT1bODcc9bMzSLbhmD
4yChMusfCF9PerMdJSJEAVK2/KMTdEQseYiXn8jNGqYh2xFH2PHwAKfV2dnHLEXPOfe/TSx1G4mO
8IdE9LwHwjFUXCs/7r6VaTGJSdbexuvbggdNbY1n9Ln2pqccp5gH8PsW+5XCMs2Hhg2+GMjq0ZHG
j3+WIDflnporm1YgDeSy/uaJz2AX5+k7SeAQBkBpunjnDOQLWrocEpJ+ixS9d6nR6IZC0z8J48Jr
fYXQzNhACzgp9ZkRm0ybKBK8h7PlABTtY90R462t+JSBoXvvy8rzwSvh1GQf8hdPuJCrHLrhn7pR
RHn20vCJv+JYJEgNHUngNmBY5vG0ZHKdiQ0HcmCtXH2uuUfarz+sG5gtoyHN08HflrBT6ceWo5Vw
pcQQLMFCevvsh//RNuIIyf801jx+aCni2AJnEP6n4TriJTuzA2u+MaykhO7O88yi3ugMIGIWhU/o
ImZQEI5nkD6x6eMUtS7bdGlO5w0SehSIL3LGZ+2gomP3DlRazNpUjCbpShMDdp0FbfbPCChAEBPT
j6jNgIay+Jsn2gIo5MoufWISyTcrzPx2DojFpFdrY2SRSlGOBV8AwnxwinZJ5HYKO9AcWfpvXtL/
j+6iEXqy/mX2BIagqgj3JBNTHfx46MZ93vDth+2Wt1tUqxSK0ygjA3GC2F0oih0ZkwVbzfmQsRPO
hAG8W01ekm7DB7pNJmg/eHC/dqZE4UlW5DgsRZ7SiYuFGYEJQMZseDYNzudpc8rIbWphKGDhuYEk
sWDvd+weg62ojjqdDBYCuUCWl6JfS/C5NKsfWWhFvKtLbqXC8UHYaNK4e/4k2Mu4awIX2cJfHtXs
KVgRRYdeB0aHxOd4o+8Q9WN0XXJZzZ4k3RMv/no6ALqG4rcgUHA49oouxey9vGoWovsAnseRJLb3
OQbzEtDJ6haNVhEngkNX3lAGXMj4b9K1GMLCp5W6wISDOd10VHuhKGTmK3Q2dgz0WhlEqbGmF+37
hXbsJ2GGoFhmF4jOilrrhHqAhRLB0i5QJhwARqXT81NunjDzRnWqDYpzy8pvv2+eccA+YdViw2iV
gnYsxC9QDCx49PEi+XjPRnaAeRNU9kAmsYwXSJD6HL8rCzNnQCMA5I59qEER3kHnbFtizJ8pgbha
6cDd6/8xru5VFNTuw4V04xyL+P64G1OdFSUZDsO04Qb/NeLAbX4WQduq+yhC2uhVolpNRUrEeWbb
i/r8vM4QxcQPfJjYnzUCLsRRZ890O1FhPjkTu42yP1y62JdrPP8M/eCt7XaKtXcQcYbQ4XPaEHyx
uK/Pv3q4XVMnXNocgnZkKyR58+vmPOJErf0TbKhAhscWw/w8URAYddYGshSFKHbfozRoQKSQRvmY
F8HY5mjD+Oa1RRPzC/uFqIM/K+ji2hE9KKgFdwMkiqImmmh2cWzJzPwGqTSETo+VsV9pxpuPkMhY
e6xxrKFGKIVS0uztLA37rBjOjI3JVgsnQEzv9pGsNfvEfgqf8eIOFwB8HsvlM/x1shfMfNDf0jpc
I60I6W0Pxfn3/u1KmSBIU4lf/4HBQIFuhhxpiJP7K7olG/iqaJ0npS3BKHX0k/p6R+0ldUV0Pxig
/2DKPv/HcB8HeJXYQH7uyb9J8S2DJNbTX4vHCJh1BSb5mXYnzGOjEiE6oLIEfMnm634rdrKm6Sbd
jg2O4McDz0XI9sIC4cD15dyx4qUW+GDain+STeEsUs6dlK2XIoyOc68DnCWjG4+xXkGmPo0M6uYs
O7L0s+J1rTTsU/IPecRd+s1boVuD7kEk6P/sHVETm0LdvoJzxCP/7PMCb6ZnEN0usbv4gJx3XzLd
PhUl4ZsSyvYmCs7AhkMW6/f/nBbKu5ZhOuFtFETJ1JHNskhThZ/Nf/yOI1de1GwEjRmZ33Ir1GC2
VXJB/o509T/lbwey1JSBjs3M395JK6SwGW6h1jcw5SYBRe2IOTNYbZJRtp0X8RIsCulKBTKgHTSq
KU2OttaThmlYZm8R1KRDbakGrNpUZq7wIB/a7pXmicQMAo1vslScNlgS6Nt6e2XEWI7Ib0TNm7vw
BnzeHxUWqImqgzmEPDVqaMFk2gx+6YgUqd2ubIzqnesMifGdHuwl+jhhfUaMwAtO/M16VM1V5l/u
pgWYVeEtd2bWowRaGLHYcx8/tbEla+cn4PAxBkh1UcPXZcxsBQyM6jpr5zt86aE/rcv9Nf1BBH3i
AWWDt1J3746M5bEAdRLPfgdrRmQ35KctJuZQTNs0k1Xh3M65VTrH7Y+9LPsljBkT23z5s9c1cFKg
wtevTaJxmFud9Rr9EHJ0PlHIVmjdQZY4DBBRrbFooJiELggoIGtELYYnjRUjP5lASoW4MzfqFOrg
ni54HUG0y0sKfHw1NiYkXvW4O2Tgrgjdo7laUfL4GSh1VsZBDsOPgC9FZE+DroFiuxEKrKfVAvP9
aGebhu8faZdpaOVGNa0dxKSpvRvSuERFDEbzlWJiOssgmUUfnCLBnbNJ/mY7FFY5mSr2EdupKK89
aewQ6aD2XWNsv67xYP2qWqOqFffOC9CgPCzjKzewFNufruD2nY/xRAjliTIoUz5mXbonwGMJAK+R
5OUO6FsDP4yLmp08Fh5c4MkcNK3lX25ZuMGOD66CafbS5qwy1HPtHYlC51pb+sNXucN8UFMpPgut
ddZK+QB3jdruEOGtSdHWDd+/US+M9byTEr8l2qTdx9qi+Cj0bey8b7fHPEwjzzjkCmIg/mtYWpLY
8irayz0IEpaNXCzabjur7ffoHEUVo5F8vXSaKAjPxiabGmkRNVpmeQX6hK0+i4Tfl73kLiOkwMH/
jDeZwLunldA1N+sN7LQGLkeBRvMfBY+JFXxzbLLnjXm7CuBwdJh0m101vRDol2tjWcL4BdAZ83Lj
4oUUytN9Q2bwUoMKpRxy6eXuYAJZNpcypw6j6osZ4DYBuU+o6c0vzy0E9ExzP+s2aXJsQ171bZqs
BalEo6xphLVy7HI/I09CThtDbTdzdKTnAgjmwLYTrAWdfKWMNE27JAIQpdwq4pgcFhWnxMvhp2RB
/IYs5ZTyOep/kqy6hnwrpzCMT5SfWyw6M1VUeE0Jz7+nzf9CEQlapBdztwzmaq+QnNVLIbZX0+fg
+r1glPU8c5RYuOxs1d02MVIKFqecaMTXBJBxpdu9lGa+J+8tv7ajF8/M0ZPB9avMqHzkir2Ap21L
5QFIh57IL4bS/+Dl9+6L5QvWlbzmf+syT6Yq6v8iBXt/xyAVGxVV6ypmjKvNZRmWCppLplmI6mnQ
GrBsgzt3tIGDwCsdSRtjiYjrTiFRcLJlpAPDXjg0lrB9umM6s84rPEegJcufATnDRWxDEtBiJeW0
9ab3qdNZkKeanyYNqQ4PQhFWyUMsvl8OAZxtzyi5Agmwpz3CrUQZnAHbjGAosoSC3bVRVyFsfoOS
sB4IyfDsDEIF7kxqEGYftx7LaE9OytOh7b5C1TbLhTTtHxuPEjABefNW+VnQt6/qCPQjLSefL5zX
tousD+A9ODueRSsZi3Db3rjzdulCbYTQEx2LhXIJRGEV4UYJ7CmRyIGyV2D5bqG6f2q6Sw6X9s6a
11pQIHGi2TNEWiFftzZd/EFjj8KiCZslWi0QX7KEe6T8e5jeoZvJ9rSMVmFUuumJLn0j9BHFuRJU
QdlSREdvp4gxE1h96u1IuWrYVjc77vSWb530Vm3F4WUPCBmRni7BKg5GDQeqmlH9zt6ApdcjSJ68
gJGUAws73NH31ipO25Q7RvQCpYkHRwNwj5GrmBGbgVHOm6G/f6YLoia+2jT/KHRsVgMzx0VZz/Lh
jPx4g/1QJZkWHnXtDFQP6XvUFGFZKx7h8l8hHmwJdJ6jHb4LFq3y+ogp/1SsA+vbcHVZsJOxxZnX
F6+2VUNt3ZlPL68k3iIwiPpDxl50CqIyG6Q3XUUexoVJLWBVIEU95vOlsSvQC6lU84pvix+o1P38
vhD+YqVhd6WjdYg/DhfnEWOMb94djr/Kfc+17bZqoqrqztHydU2N6nDQbCeK7wwwLYM5QEN8sFm5
KLtCGmR2Qf3O0JlXn8k4gSAB+ULHiGdId+GMHy820OSuJpH4aDYNSCIdMNq4e/DhPoGvPZK4vI22
v7n0x2Fnu0+shGDcGuYQidOA9GwDzbV+q2UMKRiKmE+hp0iAon+IOaQden0SZVVeNoobq4T1q8gX
jN7JLP2rZ6X3i7SXd0rmQ45w1Ay8HDdQ6LYvRFClkGoToNH0ER/Ct5uYFrKFak3V+VlOIRyaiBDW
EZo0Vu7DCdurmV8qiyP3mwn4U23S9GBbzUVZ9PsCPh8N6mugBL0xrDpUvYt4IarjkPg9PdVR2GJx
G9bRc9PWufxzyd4llgB/GU2WrC8fBT1cRDD7Q3WELHEPtIJPF+CNkKmUyBZy650rQroYc2v+KUBN
yjMqqq7hWwh5+p1XA+Z7y2ufbKfZt9i9BbEMRNAwJnFPyaS90GWFp63GEjJZMmS0pRIZ+jlc6VVx
nYuAVPmVR8ai43ghU+0EpUJ3X5Oe00Y2erJpq/lbmS2+PYnjDGNXhlDkYTHMbPveS3ySEiJtiIxq
yh4JKC/auqooiN0zT4HA5kQjHuS+yy1YIN1C3RaopUDfymqLAiQqBH5i7oJ68fMjdp9ghqpwPBM0
WcbewBQLsyZtuohAJXUg8El1oxKc9TBpp1WdrutTBJ/I9AIcgMni+GmmGLCqQA0UwqqH37cBof1Q
aYws7B2EeRkKasPggC3P1AkcRtxURnisjHEczaUk0E+L4RfytFlp3UYOFLMVp9lgSjA656WHsTCP
4JuToUFzhoiDQ50nddzJqutCxzDN///Rhcz0JUMWaJ3Na1/kjUwXcPyhlbFJ+ozKVvB9O54ssoBA
a7PrdMixNfcxeQDevaxSHO9Xn8U01XY4p1k8ZQ3ZmmHEB3bYI6gU5w89GgoVYt+qRmuTs+anLiod
AorDrItq2CYdTKMU88XRL8AHqimx2tuJkreb4H0mO80cFJkiMjpa25qDTF7SfwvPZekloFvnKChQ
UFttsBRIQUJLGMVVpXoxz9mzHyzlEqNwDg4utrlKsGcLuXpqc/WuStEFZWuGuxGLWWOnqzB96MsO
hJ1MwZgVkwApRAhBy5yiInElX+nzHVfG0/TWEsFBqsT+awbE49jPj9olEqxRH8IXbvPl8zVlSbYt
PxsQu0/m0/9qryfhMVrgYAvle/co/YkzqxRbbLOz4BpneEaEQ+zmhXr23sh/0PofOwhi2krALtnt
0VCMkSaaCeB+U8fF4VthgzkabRRHHLV1+2sNM9BQmXcO9S7yKcKriSuQRQ9PRVeZP+wZ9Hugk1Hu
ZjfvU/w0Phv8ro2N34Rxm8nNmAgcN9AsJt0bipUfrwwfX6lKvLogmMKXot7KXiVq5Sj6f70F4nUy
RngDkOAda6EVpmgqFyPyPPsThOqUb6kHyUN3FcFSiXS33Kunj5gXRhnaY9InEJ81FkLraCVWKLqA
ExiKoQvjOnkJFJEQrI12Yi++sSRS3/0eMSBibIyvN2NVgpydZkb0Ssq6YaJTkRaY28xhi8PksHdU
+WoADwdr6bIa/DYn7UttJ3Wi7TT/GFt/Ml3fUKRp7hocyFrp6bYUUBagrc0DEu0uWFfgSdu119tA
uWWHTSmgIcDuf7pEKZoM5TL7ASV0LWiXrNq3GziJT2nm+nLtobsKT0EPGC+S330CWqyAkkumDrUW
hbwRNvitoOlJuEI/ruK8WCcoXrhE0bOGyiOG+CTLuCAIj6u3JvL6B77xIL0JdsBARpMdkRJr169x
YzoB0ZrxR/4OuFOKDalnu+UZBtBmPbqkVbAz/7KnR7x4DLMT4pr/izFeDvU+iE1nuRedwY2Cm7OY
j8U5uGPbdIJjhSOlr1PF8Q0CnfeJ7BSJBm20OGVsB1IWjAKFTgfz0ZqYU998m4B5qb6m3uyA1GL/
Z3zawAqnJQ0BmRO/FZ9hIszPEPxAEsk/nMowU/TdyZcg0t5nf0rqsfSny4jAqb1mWx0ZLm6sEthB
LHR05E1ZOZXZlCfcu2PB9csODMZvljq8pkC2pSBwMn7Ttad/Kl0mOJdjioxlBte5sBGrUpixXJdp
GHfQ5qlce9Pmjwlc7Wqi8kKtdyEbA2R7G8V3zTWQO5l07y4635sAPLoJ6LE7doxzYKbRpZeQBLDV
KTAoZXovsKvS7fBzWFSY7bUhx823MfW+PtLX3OrqNq+1cZDd0GN5qm9tK8jUV6MawXelmrdWYi18
ZcJu0daRpyhs44fUvipm0ygoa3ThASdQEskfQxGI/+I1ItJnngRZ2p1NHpQMEFdy2F97jxTlcQXT
nA7KcolalX+f1G6MSdxwq9Kr91uu5Df3WIpPVD31YXC+wGb0NlNA99k/zyAByAqROttXlITQcHJg
rpgnkmB0bKip6lAb0NHc4rC9jmvoX0G6YPOD775nD6dfcOCZMiEZ5zV7r4XfiJbUYinFFRjXmVfk
MoJlezWnWRP+Xof02IFV5vQSDap2zUvfEj+5HLHAdVYrtwCpUqHkm++DbHnKYKNbqdxHoauvfizM
OO6oTE7y+RJ0FGUjnqALit3MBstwlYN/yQME+jwR/HpwND5y7M3G/gzQMAxZ7qvg++1iUHgxwlmL
9uzMqQbfXBosFgx06By+F4BJDT+JhO3RvqzvJAiHq7CRQT2o+2veUp1vqZEhLLbVcGxZ7NhlIe8b
gOhIxbdL3ZCdcun4CzKRAJyJQAHXXwRFKHmAFIfjz+80pywVIXPRjkfVzWXxJ5Jdo7m9mzpbbYl6
Z1KOROlOY6Mkd68y3uIxV+/65LbkBpP8fmpQP06B/Z2Su3N2JRR5P2Ww5ph3+k/wcNBXjaHtornF
m4drR0E4b80wO8KoxTNTVYY7+dqWUKkWywiKIEwqkP/dA+3uSPmueO04PenB4ZvxbJqh8fb9OwVj
+ODSxsXeNOErWBwTkcdVH5UsXy8cIvfj3Fh44tzF2pEacGUZWn5IofxVqF4PCJ4dRF2oCyTO8REH
fLOzIt1/wuYWf/xNTcD9/SQDI8ZGW5Iqdh4fVbvIuDsjHOAX3bupWgnVahKvtTKm1tTM2ZkE2Kvw
zut4J9cHK3YJ6zINgyHhr4fC0rTSwXtRgHCVSHYRCcroHIiwsJpGvjbZcjGDhoqW3O04YndiJoz6
sXXyqBHzmrLdfVhMI9669pGyZCkxsxUGR3aC3EUDTZTZ6FPRXKrWix03CgKATlFy2toolDuXijMn
ejnz3KDpNUth9CZbLtoPxPZ7Io/Vt1XhJon/JNIgaO/MrZk0MjOIr1ESCvXcC1f98KSnjXaYzhqB
/WDRrXrLBAI2cH0MVQ4PVv1tOqC0e+T9i9nAqd0CZ0wphMx0MwaxeAwecXAf4/2ysFWFgxr2GGGI
QGwJpxI6X7/ZXuQAuwrC25NWhQw2kZQFUT15Yhto/F24RDn48EXq/gm4bZ/tq0axkgZkurAkregy
cBqKCiBvKGekvGMbdmN/McGvgEJwALeZ/Ya0N/MwE448owUt8wpCzCXznVAvwqNPPmAEYQIY7OvI
egANhP/8KONwFZEA3Szv5TDXGrQjHQqwdn7/SR8OPu9GszRRv9wP+K/knAd+0XZC8lCekCLVfhWJ
s2DfKjyVeiO1mnqiRb1WmKdHiNn4Axj1AvLKXct6KqHHZ0+qINrMVnAmU0hfk53msr5c3BiPZsup
8KmSh2zeFMsKL+beELq/ZpssF+wA9xb6oJ2hxdkMTRd4kGTex8Te+kr/ALM2lw+pXLHyqCCYgE1Z
OnpsD55ljyTx4dgWaLS27X7XBpCbDBlS39mWyowUxCOPNkO3zPJpMlmtetr1q7fZyesbU3iw/L5r
oEqfazqI30LGMETkh8nwYzXakWKKhDaWkPBOAcsBh7qWlEsyPHi9Wn/hSgtybfwCbj3wbThUbhFL
grZj7UwJQzpFThQxIG93/Ad/lz47J3LChNCqzPwKiY/v92jegDNGAV16HZpG49tT4+ILTOJ3AkO1
9Tkygw5LMtR9Adgclqrm7BqkqyB3t12omPX1psp4QuUUYoxnGOeJC+ymNloHtvRGACqd65s8RSyv
w5LKFJVhCsG8lewEaNekWDRWGxVUf6MTrDIPNuP8/nWWjU6DCYhi7roQFudsrR0E8WNu8D30mghw
Re62l4Xqh2TtXwmJHmJNRUh/lbiS1jOIyqifiOHosk/mgEp5oJEkbqkmSnHHvCUw7hrcFc47yrj8
RZ2vyMAKBrORLGdHevYvEvJ4jE1U7Ubrb95vZmtBlY45EU6nwOTZDemp4fJX5aQNvr1MbkJNjZoS
IDOyvPKYZoXnAYPWKFLQg5HSRNoiBmJnHHQuW4GP8rqxsf4B8O+uDENQPramPNgZ2G6gCkzZwMYV
1g97jcHELO15qCF5gqtD/mvsxfzMHfCFaDVaZy/CQ+zGmMpwvfNJ8yygbzfSSE7+GgbQGP7Yd+du
uth+bnrf1FeCjKPYokTqdtLA/uK0wDj8CWIhmot21yzb2UhxAK1xXVcfRGRM+2Cq8JFbinQEDesl
8ViFwzM5WKW1wEnROAtXUWIZbCdlMvQLxVm+XZiXTsPn/HTwzdSCEI2w8yE0XKyaABziQqe1ZocA
qmAmJOoV7+xB+hkRxi7yUj7PKToNazBVPmfY5FpiNN2vK16+fB3r9V9Wvmc3A9AcMBpoU7A6CTFc
0+r81KK+1qY0UBCjckgBFVilHuJPqFKin5VU7P2YApBIaFdKmnueG4An9461TT0LO8uQB0/IdEqW
EOk2BNBwrZIQjadmnHh+R+GgiAQVjM52p1+bP7/hFW7foJ7hb7mKE0NnS0CtexTBOg+3SdC3TjkF
VhmH5+A+4fPyinb9OUUxKh40mdRZqgk8g/es1YVz0vaBYe9KkyK0GtT68HCrT9AsqsP5i7U+/u4O
5TK1386/iDtoeCUtViEYewDBaGOEc/YlnF1Sm6uQNP+BA0BPaTQHDat16rJeSwR73ZK0Ze8lMd1F
4a1d6FGbSxoy1qXiarYXhDhwLbFNNSB49UFMRxHasGfnLhxwyAHof//FfAXtfUuqtYmk98EBWfUc
ijdtd9+wVIAhb2h7ylkZvpuT+pi+3EgySwwfXadC7vDjyLFEnlJw3cho8JonbHe+HYAKYD8mrASk
RKYx38fK969WI2q6lWU1A+4ShSiu64E/V4+c7ri025hUNfsO1ZJZw6LtugNACHCvlqmHQhLsOekA
vv47+8G10Myhpx03+Iqy0e76gXcpj6Hg4JWbe/3YIgfRwu02TJ9BHu0YaARoAOtJdDKZaoQIzZ3d
TXhH/GDrF8ZlTLGVFuL9lbsDEKT5MyeMMN5MJacxFtae1a5kbTZBZqdnH7Sh8GEFDyJCBCgJsoQl
hwH/3e/GA0ekWb/mztWpIYmgisz2zL22drFKgf6mBQJQ1GFBf5mtO4wnNXu0Kp1qKO8KDDVH0J34
ZQPTokUWdnIYORh9BpAH+blp3E3BHZmBYDTMpb9gEPEwHUDZmsW99dLbK1uOv6m0bDuMzpuABJtL
TuxfQyQ1UTf79jSN/reEx8Dwd/Mtl+KQeWCCKl8VzNJqEeMuKadZ3cEtGvtWlSQv2xYXen5j7Fwq
NbmeAIFyLMFjuKnwvmxlGaFSH05WPcvrNgxLCnX2SdaKsf8VvvOVfN9kr37eCwhPVw9KgG9MlWe1
QptmdvNIGTI47N6lvfs3pMHh0wy8vhZpfjIYD1aulJLk2FMa653iB5W93K1jS8ACszpIjOOJHDBk
ZYOKhMLo2CCSWIg/R6ybFt5lIEI/JMrdk3VzitDAEwUq+zcebaX7eGiKpEhtQm/A13n98b4cZp+x
tyVYjSSIm2sonXJNbLT1zijp3DoVC37WQ83y4lPCq398TEs90wxZ+d95g3MpAg8sAOyOFXmMZHz1
iucj5UCmiDvdLc2Tuc2yhu4TIowxQYQqxrOaa0Xsyu+oqK42ekFiJZOnjOH3jqzk6FS4Inb0Rz+j
I+VsauuJa8Cnx0uF60OIPc4tTMqBY5VHZr0vSRIREfhmRLt5ULtGw97o7QiY8nkMi7tT0qpxMMeu
KjOlNnMEzAZr3QBDSTEhIiCR9GnloaESrbJLkC4F6pkRnoByqjTKy+NDcO2FB6OAufL3zPsbGXf9
PDCITvF74slcQta5t+ID2ZHrXtbc+MQRvIU871FAWe2rf8Qgt34U1lUMYtSlh2WZH8qXcA4dGyzM
1PiybkxeTwBeeDfoZ6lkrUFzV+ZhfnlWb5pUGNuLoqZR8pXBABGNMgFBS0ScjBGtsxHISWXJeRj+
mgyezu3iycFj2UWcQFSHV5Mvo33B6Ogv07q7mK9fixK88EdSvIE9g7mEKl1nbDe0hS4DwuHyB7J6
/j8bYGo4T5Bnzu07rGHXCbFkTK1KPXFCN4D+RWHjGW1v598j4O35FheHJ7ISKAJXX1rMFNyVtlDC
nJ1GcyfGQ+rihf6oxiyaLvQ6c4TMPd/tCoP9xc//pJZRjR7QKG4cPEdqx/+qINMBHsAUstJHdPiB
2/E4AzCCALgSE1m0CHEesTNJKV7QK1FBsix23ymdFK3ksw2eXXuZSPVBQ66sIUjYAcYYDvQN641N
k5w8IrIVVSok/5ARgHucnVWP9Snqp5h0OhLjUgg5YY15yrqW8dfgDTTE2sbeDxUS4cI5LCBHXk4U
cUJ2NKPDo9idTqUXM78CyR5FBk7VYY/UGh9tKBbFqud6bn3s1/Yz+UgGOr0fq54bPnCUkSC24IHL
mq7FvthX1/b4i11Zecezzx5aFv0LHx+uMLRc7O4PktPA4PgLX9SDkeUP2OSjzUhEum/iYyHy8gUh
gs7BKQJmmL4Oe4l4r5bVcqLXiC5J5tH1VtSQmMeTVAlZgWNZuwdktyjGuydJcvn0YW5BBDwIpcdj
+mkHDFDRviZULKYbZPKxNwJ/d7BGv1ssYvgXMD0HMnwr171oOODLRINVsOozFgGrnyX0qCtlS/9H
n4vfKdbn+tnUi+mMhDdBXV+ofOEzHojYYkKFw2BOKZK6EyR4AbiSmrCYC2Vmk7AXbjOpUybcmVx9
7FB9S8AO3HkJyKiEePtmbJYP/v5hAhQ+FAZXOxqHkMfGdZzSszDhMDfx1Bcf/d65VoPqGe7Zg8yZ
z8jtug16QLxRjZ+D7VmpGk1x2aIvZd9lY6FvgVYVy+e9awXTRaoD1cYAT05Dz8H9IGWi3H4C+YX7
lDWvT9DfcbQH4VIDDBDnUqajv4pw2QxKSZJUFKF3rRiayCuvfGHJTqEnixOpTRQPDO/+KWCRaDNc
cLM7dvPeNi4iZd4HgxZAVaNcnMuPD8muPybBrnZ3kTNTgWqLhD3Olby7dkCBjcYKt/fPTpruhrB9
VTQSX7GxuPffyNOdYXOxKba2oUnTGakdjn6p4BFGLP4Z55Apm9NfEoytgRkYRtKhd3pAuSo5IqfM
8BYYdKlBQt+yeV6oFKDZ0EWB6an26vi3Nk0FMAh2HCjWsuN2Ab6fPvUmUArIpfOosqm3Z5GyXJyC
GK7i9O/sE7TZhcmhTFI6kc88iFu1hgjLnF4SuRz4BN0J91a7TFM2d6J7lSdAZPIyN00ZbjqDx0xb
POLL01WARd1q5TpSw07c1KGAnTD4fQmrFSdHBRHT+goqjAy4ChSsMtP9pMJ8jCeKXdaq6ykEI1/e
d7m0xafIVbEW5nEHicqQhWG05SdW249ZUL1Ae7D0VBznIcUcd5SQryDjurdQNfhq+i1EHh1SCYdz
IXPHns+RESU41IaChlnKOU/I2dXGhQkGZnzJ1v+YYRwYdCPft2YZxOmJn+E0FhPF2/Wwb3I/9B99
a6TIeMFDVUZWf+EscGCwjD3FjSx06FDdbIPikTL6g9cZwyKtYRIy5hmovugpFKXkeoXhA8Lgm8wq
ZRZBDK9EDoC0fWNHqOpu79cvt/YoSp8wageu8AF6Iax6WCUwAOZXpaoGR4G7PNelsC88h2tYcX6I
EoMtsPUSFPVaP0wnCcSJAuvcNd4hJmhem2CUruLsJ+gBTiEmVACSRB0c/9U0g2Y7PMBEC5bR+Buj
w2z3U6UE6pUwsScXLNmMyvbdcETIEpocoUNfYZrQEPhWFTLs5S/fkFzUT1skb5mrD4LXjVyZ/Wda
zYCONZs/ksdJh8LBqeGArP1hyx/XqxLcBCeYH+y6qJoM/13iZ3q4G8rkpAwooQeCV9rH+OgztyaA
hf2qaKRwUr7mMH08OrzpvOHjQajPNq8FmcZQgbOSIY5G/C9mSPgna58YYMKcOze3F7+qqIz00FkO
9vS0YA9SBMdDmmm36J0xcTsMAn+4PpzeRwz68HS2c2qvr9oCn0RlA5QJy9UeQgf0UPcS/S/kAFNK
QI7+sCcN5dTHQTmei26+aoq/Lk5+dubeeB3aUSFbYDU5HbvmXVse4FSNYF/M1V0VmmkVg3pcrzsU
zu5UElI8CnrxTOkOV4av07bjYZ4XjYEFw02vEzVGxnJcIOOi26gxWg779dC8jI8ECQEp3OpCBEoG
OFAvTCGL7OCAYPWnnE1HGTUvijqcCVnuoN4T0Ixha4gMkNIAVr92ek6cDUN7jWqKeVQOB7h4xTnO
eI1AfwWOrSfnoJL4BdT00pki+aXVsX35aPEhFBwnhcUUWuu3pIGzIppy6Paq3UAR/ndBTcHtfZKj
PgXMLC9L1HQd7hnq6WrwXj5ipVMWoB3Egva1lNeCRFVVMYuRWKaomMI/+jk7cPDrL7/NO95iLwLr
546DsWbTUSbgfuR3OC3HHn9ct/CiXIuOpG9RzKzwD6+poRNp+vnns6chPC9A4bAmYuJfrsjYPDxB
kmMRmEb+wWE0vb/akQjBVeuEqICuyIbVVy01p58269MZ94HJICf0ixL2zt/EDBxRh2Rs8g+9l7KB
DVnYiCnmDxj6FPdZS9/fCyrzlYpqr0JA5Py44Vaj8bbljM43PLKE8cTi4KT9Uyn+P6F7zVAsnPMW
IlBGwTr7IlZvA+k06aXiFxDuei7zvHu2jC7eD42D7B3GGVoJvCtwAo+vyWk0NaPL3cmYOwEGGGmu
rMSNa8/rwvp6B3vrpXlOpiCumtcdzxwEH609HmUTFVseHG3mSn1mq/wHGjBwgXPjfkrtB+/kTPAx
C764e45qujHKOleO7yMl3ogwCs8tNkgYg/n2OTXZTuyjBNEvOGD7T6Tg9iEU6gYJR8VYxsdM7UIT
qqd8/jeWCGYgLBUYAlAVrJS4K95hAWBTc5NKwjxOje2u0KLg4fZdXJ7zSc7YaJI0bReGyB6IdQm1
8C1E9LvEB/fLWV5dmpi15VUQyHMCFusuHuTkBhaldCUae9v5socxuMEVyvtWzDte9m1bTxv1/M8h
fCueiy2HPpR5mCU0BJMQLb9PnKNMvRE+0Vx9sVXSg3ubCQWGAmtT5UMuxIUVVyUKTFK/yxa45Scf
78uzxG3u6dzL5j1bYz/d/FoJmuYAFHLyjcwjxv2BJp5dhwcx81y3toulE4rAegQABxkGMUzuNFjl
fux994Vrp1oyn3rwIsbH7eCB0UD285LOHgGYZmOfLzpri9PrVnmD+rlmormBuIKV4WV1WuvEtSO8
1gs4AJSGWY3QkDa+zq5Yx3Y7dIsw5Ra/f6IodHmEuYfnmLj2/zLTNUVQYsk6RTXLZwjSsDg/w3Cn
R/Q4et10qIqRN47yt3OLB0ToaF/bPcxiwfE+rQ8JXh0LLWW0qlMGFpKIwmjrMJ0iOgSx6cEG1z6d
HglweAw0YNmb8lry+eHiGKHTpzatWIJQ4obCTM/oFrp39//eW3yEihvygEUqiccE00njJ2d5VqZe
ABXfeyplSoXpVGx3/LwPpqJH5rzx0+ki2F0AQEwwTnhJMvbW3UNZuKEQa5BzAEcoQn1EAI7yXEc4
whbDXIyYeKGg6LidMLPC33GbWjXz7Mp/6IgGl7jBnmAN0gSAKnHGSNTcY5RtVIP9D3l0CjUOGrID
TIDkeZj53TXhlEZ6u0glJICmxHtkyTPnM29KJMXJ+BZyLZPy+kl4IHdXiQ8vDNaJD0632k0GxN3r
eA/Zoeuys4I+PorTELRSxrUHlT1RUfbJOBjOJDTBxZq5B26nFMxlKoROYrFocF+JwkRWIoZdkBD9
89emZWfDXnCNIfela+XMQgWzg7hqBiH5/3r0fi3rTF7dHMwxyaaWh2l6eQowt/1M/iI6jONdFxzB
PVFGkTIQAhgU2DmP9TqE1dcM9VTEdKqO6PQvdRQMETMmoFBzzINu3fvV2yBhdp4y895fPBBcO9AK
cbdzbqkCflhDmcK138HnvHsIUGCj3rjqh3B0ggKGWSc1FrvTC1fQ9elomg8g/B01FMajllISXQQs
E66tFPiqXfchtTSWeBIQ4CVa+IZYHYJVrCL+Pc6GoeDqxAKfPhEyluJTPk/am6hkATLqCqWpcLWN
qoiL6LP+5jPj6vSr93vbNJP82hY1mqELqjsTuNpiZBVJfQ8we1p+jh6b8PsK1+e6mt1obE+QvzlQ
rze0PI0ehu/e68wipTbvx47xD1J1s7jpqkHYnOkwawJ5kemtmQBDNWLlBVUSZz72Ei6l82/N2UgM
iv81qfn4mjL2wrWWDukup9zeityPLOzrenZHErmkXh6wn5vWGXYyZYNzCWN2D/XUyI2N+muq6i4e
Gskrm2apnvz7Rlf+LG08Wgbvb/0Pk+aiOm05pcxDgxxtHH/vZpNXkVl6ZITG0OvBRZtGza6yYYGo
BLKEM2MnxllbkfyJxfIsA2OjlkKQmuxOBA8v53L/DjBfJ3bF/m+U1HxK0Fvr/edlB48HcYDOffXn
5zCTIjqvTCe0rC+QinTfBTzc+o97LOThCKdGcli9bOAkol+H+gqnH8H0NGLYYmhOdeU2mJMx6BZL
zhEeLJoiJvgn2mlTu+1aoFtFDjmagbLSEEbXYAOq7RrsdsdMKBl65Z+iVekEb9BcPdXsgXYKtKDZ
2TOweOWuveXP1CQ3G3jHdtRz2ZOySP2tLJwxxEEVl+snlb5qq9rN0+Cr5/2j/yaw/jf/gXlVBJ6R
iOwmqe8+zbYqRcAA1kjQ+ZrrMUSyzE0xd9WYqWRPp3XduTfqkSutxri/1P/ip0kq9xD0wZciLlx4
GFTWRC83ZXKHo8rBzcD2rPvxQB0FyVfl+Qx+Sxp+SoalsL3aPXltbVsLOp9+BsuQCbMrcBrKyupk
V0wd2BOoZighSjpUfYWg2cxm8fyrrXGVuH97CNLyIuiRBgGrKuAGK1Ppj1HSHKNkHB9nsWSADU0+
O42RvzpaG8sY2VbxfWvVv+dz0LMIBOnjvOR2KoPY6NzyAnKqATtIKWreSTuH8bdTuj27PNj9mxbr
U5aqz6F/Suj9Mx6yAJhF5Rr7THCKJpXsA/yUpyUYlxkRG+unp/yK4IwxAK2g1QCpDj0lB3ORy4Qh
JPXDGGJzTicnwNzkkPI/LTuEG+0WJhdaMs15+O3tb93EduR9fc/a5hX1QunvjPgs9qORaLUgWlAH
0pPwanW02YY6Vk/btqXQLZIw1sfCtvhfHZGFEw+jKBHTMJDgtDKn2s248V/OmwnzJsW+SPEIjqEp
qsAUaOS83XVAyHIPaE5yVhUu2/zlHtGl2U4MLHTvH8S1y/b4A4oyEynQb6nvLXs2mABa5WUW3d78
LI4rS/0ajirkBVS9g5P1Kw81/hCLvi7ZlHO5nbZzeeqKoGUsWmA66qVhS65AgFK9bs09Aszy65gr
RAoQSLsXMG+ma5des6Pjj/XfViVTM/sWo0d0SjGRDarFcuU5xaxMhaEyL3CIeAp5FBX/j7Iqja7i
SbL5JShhIDS42Vw/PqPCUzJXXJX5L09XMU6T640f6pWFXZp+zEEie2378a7kyngNVLdoAaUgUS3Z
FERDNBacxG9NMYGjzX253HHSJERGsKMwIbE7gMJT8s/9vzkoHGDFFtv1jrG1mT4aBSijk9F0fPqE
QO2BoDFU84/wnXRKuKlgepdGhCcddNtgfIPqCTjj5Nlie69OaeJ56vqIDkRpQnTei6LFhhT6gHby
mXsFguecp8cWKBawNQQM8+bFFTxCDMU/YQPaDFSiPOEG6zGHJowifBjAq+w4lOhH9X02hYjGRyX8
73mxFWuAgRkMOChEDtq1XcIBfpJwcQjOSpHq0CDjWHyWqXYV33/h7uJFoXB4jYIr5wUKpcCdHDrX
2QGP+IyvdBY3Ik8wxy3qkR83vnajzK41XDBoSJMrvIqeC0DbMTu1szj1HRx92TIMJc4Ka+5B8BYp
Ft5bvKUw7JMvrZ3mtN+3N4s0rrcCjgzvvZ5h4NQLVV+dWxmv47Qa91xPzLCmkPSxCba1BQqBXHsV
ofFrCB9Xn9OzXHWqt9hVF2I4ejQ/UvEg5n0ui7IbxM1Qo06eI7uPcBTSmALRBMUiJLdhC/AnT0qM
pdsxz43QpN6FBR0Srl290c+MvzXqylkHEZpDW5wf6Fj2eScyOkGANyy103zkCgLgS0ksn23/MTe2
CEu7g7Z6tKPM4/y5OzFpBVHzzjdTzHZwEP4+MDSm4NlmuL7FmV72boEqbuIPvpA+Fv7TLKc1V7X8
1V3h2INCeoncJpUu8EqVR4VYppVCjol+PSx9Xpvfpl826iVY3nXbFaqzk2quhF82MLN15YRHkI4R
c1kiRa5i3yCKzibsH+YXaUgN/lznVUt6Ya6oeehC+CoKrQd1qmVkCBog2Hlel21k7TAPG38+V0Je
W4poyMU5c5I75elQnl2Y/ljF7AAiHJeffJw4q7K7S5D5VYoNkjr9g/SyJrJArS6j7gjhewbHAQ8a
K0ap7hqMkucwd2apOVtzHMA/PKDSn6rbFtYdc1P+wwdSPFARBraNeP7cz+HU9FjuhiiQrYaE4drs
SM13UiOjnXEYoQNnb1WMAdEJZjYQKNpI14MncDSzhTLUYgfUYLH05jh3yAMmBIUMWs6qhKjJ7Xhu
9aD3tMUbsIY3xmpTVPGs9FiR2QteCZXUJzEwR2skXJWh58qyzpN4H+eGUQK6EkNGxibGS0Vcvwmd
17rTzTwuGXSznTrI4tfRwcwrKSzJGUiZxgyv3uPK64kYPvmwzHmG9QasBYagdqqmnrf893plG8/C
V06Zns1HKZtMaQTvcRuwy8fDXZzU/bpLfA6ikpzDpbzXWYR6TTy+03CJSFuIfa7ugKqLRsAsN8uA
uMDxaWL6nFiYDsk6dCCHbVbVVWQN/pcrTF25O+Y2U79aX/9KBKHF+8lEgj9njCCdKNiKmYOF3qf4
Jy/k5ak6TqGdj9ZvIuFQ42eDltL4TdHqrVpKEBqBs9iY6Ej+gubfyu9ga6c3ZSoMnm2RNcv9ACNH
qdJ6qLDINqOfom6tppYcff27Rt/7SfPGSdYjRizwMW/cF6LanAhUeiCujsW78NIT6MaFVty6hwt/
nxXihLL09TLj6fz97uzGpHqquwdTppbMx+86fiByTbDeOejN8IHTOL7crD5H7eXyXtHga0ooCk+c
xpabaM4a9wlPnu5jy6jaKaBOC5txtDLuDLiKouiSwyFvSclUASwSrtlnENlXSsUn50BTDJKcUVvI
xC4s+nK/ZtFblYuJ1AF955Ennk9upy16wInc/0b1uZcicvGPcwITA738vTBiDSRnD4FN3y3G6LMV
ZlgjghaAkn50xcWeuEOuqSJ9N5gT2Bj431ELquXefdj0tHwjniE1C/egyqLOpgVe7yNB48EAQfUL
ly/wEdAxcxdhRUjQZj3TU52Vn6zobT8OgpudZe/owTNXBMxsi26GDIfHbEoWKB70DNfvMeyd+7oe
JWAr7276sCvmFUSrUSdYuQ7FoSeubk8ca5kMOt+tz/De785uZmfq6+mZ/JnlRv/+Da4S55nuGbrM
xT6cWCtdeW2pm9m5BawHFmA+mjm4QlYfqUyallxuPhm5Zxft9TtiQaD+oU6Ncxp4GWVNSAeTXmTL
HlxtWxD44u4fMEFe8EdZ3VovoJpMYeffEgzlDjqqdvpFfS6R1g8jB2eUAbFQSENDLqzEIaYt+VhY
pWEJCbKtNOc8LKgicrWd2Ux0/jDZPBAUXCKrImuJe4BOanrHEDfXRg9BbQRosS8kvhZ5cM9A1MMa
nbkK/NygS1A1Y8m5FKLWzj6VfdVbYaoUR2gJGC1pSxdpakHDroYCIx18BqD8XsXmhbjHd2AviXpS
PMqMlh1IgMtUcKoWPGMjpOox9M1ZCYd1p/D20KUh3BPomU+DQFdwBJGWmg82TZkSPetzEuplCqA7
Ctrn9hzhPHCbLiQebhG5RBjJdKV25YKBO90E6SEkMQjU5lnlnVQPR3kUUD1z/85y8pFPQ2vWTLjl
oPhLib5CpBQCaP9XTl7wHx9vb6HuI3+qt4h8nMNLIO6C/XvhFjjO5xBw1HlRYGva6kN3YXw/k9Sd
lOp3k/xMu962KbV82XI5BHsn29eshRk0tgxMPm+eB4//3T+iJJ7NdZwObyf84R8jh4eCGMdeN05h
KrJVIrBSOY0V6u+NlsJrUmrS64xf/DZkbmhYE1Y6yKPFNtzgDqB/MX0I/NBzRrzyhGKE2M+QmxgW
wXpIvxKu2IpTlgW2sgVEecSwg8USegAnLQz9EDW7LxwHNxzYn0WaVzqXZsRkQza2cR0UtpLtEReX
s2CUJ+PKayNqOVB6IwDKPcC7d1w0VNl1gwsd7yKtjlmW/fyKep/zpsBrJ6vgvGGOaOgjOKsFs6gh
6nIT9PqiAExRFVjGkgj1k4U3GypnWb2WFy1pcXzvgac0QWj7ku3E1gdIaU+PNfzodhCD4WZir7Uo
oGlb9s3220C+CJmD+RzXKAWtT+nHFnhYAgLb/AkijZwmB2zN1mcw9b/UQ6wea4qb4auCRn1RVqrS
vTQYTpV2UA4gqorJPsTSOVdhmevFmkMG/eGu3Ds/hyl/QkTbj33VjZ9WFCSFaLBk8hzq7tXhGSkj
DadL8Z65aLHeeIQ5HC1x1yL6/XUkGltwdBtrGKSeSB49ia1drUZ+Cyx7fLJ4EJZYcVBbeTsfRNAB
KPlw5NMPp0nvdqSSpemyAbNUdRvfP9vXIClyLyoEDHcyWELV7tDADjWGvgVftCtekKLhR5aD3h3P
/sq0dxzOZAcwlWEYe3eMJb4CJgsEymR7/K2Bw9xIgECacpZj+KoABMynaEvXJJdB02l2mMU5JwoY
YuVpd1qNlpwgiCib4Y2Ci+BdC8VxaFaXwedxsQYDEE3GJvD48DuQND4I09aZZYiS3YVTg8V5VpkW
Wc0lna1TDamBBJ5XcQpKsEvh87tlAfoR9ZlutEZyCQNpU5uHqq1CE+ovsNjqFa5LHlmQ11+eP9GQ
6jW4rPkkV+iBYAjWfNpqToQiMrPoUULHn85awGnnpxQEv7/pT4w44IFUYiPFzVTkXswZkXDsO3h9
junoyLWthXZNe8wvv6ZBXvuSJK7WOQI221/dIi8DIZyys8cEeUIG0hMthgddyv6r586ooadBVEzK
9TSvUEP1TpiZxosKFnKXek8M9O7S/0iMTV3lpI990ZnptHpcA7+zaC6Pj/dJ3n2xtph5y2T9P2Jy
rrMBvGONBp7z47jQYzffuWWsriPiTCT8plLPapGiRFi1nrgMW60ghX1++mv155YAsoLO6asScCZ6
l2pTtTCj0BmaQtdhyuwbZ1PsOWTokvdRzUtIFUx51Jif9LveDaNgeT7O/mbzapGmjcbt/+3pO9m8
h6AEshPpgfqWBEQKjdUG0qNIoCXXjxSXQ+6e4YMseMaZZ4O5/bfJmnBf33GNVOsSrFjH0UT3Man8
DDxdp9TBKz9tPQAw795fF7DSIL9TAdhX72zgo7RfkY4tHwdaGKr/mdxId8I9l+xS37bvY+YhdUZP
8/4RehYiUhiUc055ug1M/pGTCc4RUvFy/vs+W+x3VhzaeQUReoIS7ES9JyVWogCtr8jR/xTpu+cB
dGdqDLgfoxlmgcWcZa9BgyixeiQGCoUnAojaUMfvB5Af1VAlQVer5fidBexuJiAVzcrWvzqNfXKU
0BZZbk5egM1p2Pt0L+nH9F2mrIzzMQBS1a7ffgWt6KX0eQOGDbdUXYvRI3LsltKXf1lhCAQqhZa7
sCSxkrvCMdjwOJwiYMwuem/qst3yrLCRaBtn6xewrFoCRaD0eg0UOSXtRNgOqpG1TeKTKMizImqO
HH0l5aPI3vowMlrGpWafo4WiBYyq/hYZIBC3FDnAIpayEi3rPUmolfK/+xExcjuga50hzLZwEExX
3QFawVAE+c/f81mCGWKjSo14FHkQ7qOpweF9fZZJFZpGHEhASBAzNPjc4rXt9Ib2egOEDh/4DWJd
1Hsr2SHmRFCnklqPCb7PA3ABhCLR9VnpWB2F0EN9ZybeUIMYFyQo5KrCH1kc5+dLlobWhfk1whw7
ha6ixNQX3l1bIBuTi0aFOyvVo5FHWQ14JWQ1ogWjgMDWYlIqkCjiaF4ai4t4LRaas8sA5Z/5a5k/
Kuh+MWzkccrYN+fbaRhS/if/YE2RxSz7izdTsN8DDoTKrgCi7JVv8cbmuQzgfP4KkZ9DTZddMw7B
PrkKt6GIkZga5YYeQsdZQ0IC9iwckW+9ZYde0TsVrk81s/NXKG2ieahLD6v+KeO37YI1ZwaInR9Y
CfJah1cjwu6Vx61PPyZUikAHf9dk8AdN8QhH49qOI+Tw2TLmLCXPr24EUYH5QYoYhHU0v3NL+0rS
OFQY+TIpGGKp2V2L64NMgJjivEiUNaclnaJBtAzatThblJayzcC3RYcEI//ro35xvdNWIs2FPfho
LRnbXW8xjHv+2NuOntCdgXdr9h5mcqanP2Nze3NayBpuj2TU21AVWdXkvtAVM35gxX05+wYVjPqD
X/xg3Qjj3EK5cuZ5Zv/I2/ddSCvE1O7/jkm9LkquGVObcxIrXCMK3q52JASJAmfxgKjtFFYpe2HC
+/dFHehOSEvqjGr19lAb7ZH8KxQguNeevTmWDADwfiPd2vOamWG0+ElUPs0Q8zeL7sjvUDwE0r9H
IdQKSw2xknEbzZT2Hi4yzN3eyPU9uCxUx5OVM+3aTs70PQtw2qMa8zQl/nHiMbktP4y5QyxP7e9T
HZ68BG+xp1E2qRmDPPrp1vE8TQlzi8YSOgOaG9WPFjzmB2KUYj87PYyJn7G6tIJQAVph9aMP3XTG
7R3AfMjEGVTyVCsupHU7agopDinQ43lCr48GDvLJ5QXsgoNXShkMA/tBEXlxUHKj1+lhVQLh7K0K
5upV5Y6z0hlxh5bSM1idWValG1xE+VK5I0SzgA996RvYONCF7okFkpKBYaCNtDD9HH5UvSPJbSpY
mpyyGJOIvYXX/H2uFVLpIYqYRuoZ62w+70WI7gxYxIhPA09xvGN943162eYOIEhdKz4Lq3rAUPV4
Y69GKLRo/EWj+IxaH2NX6E9xqfgQxyXwv0V8RB7qG0qik8HhBmOisWrtj7cLlJyiTOV6CHqqv9YC
SyOHh8YgKc9jOP4k/8llR4+I4F3+El6JfJgzF0L81g0BUVfShj95HcaRFvPfW0jopL+kITMokzno
GX7RMVh6meK+X7tRu7ztFr9ko5iyuLFhjttxUeMez/XLkhHE86n+lU2oTrhOtHWLqQzbDb2IEuWX
yHkltH9ofdLoO2q7bvHuiHB1cY//lv4XYg5mAIBERCJF3CVxGFK82G9igWMY8OTTVbuKG2SiBJdc
48eouYv70nsK7Muq3sKulKmU3tMggr0IDASP25DkCW5f581Es71eIChQsZaeOWDF9zPACkr+iynA
9NUrQ82JUa1OQJN9r1LqgnV695z5QA82AUwdRWFuChmmrtKaElqZruzmBWkYOOzeZhPt9D5vS/cq
e55AwifbeXhrXYQMr2WBoE6rReYLnE3dAgOod+GqiksWM4vRzM92H6OafmEz3ijzYMEMNEsIAOHE
Rt8wltwSUCfjdIp4+Rk1epNqWgRT5mrKlFzS1qaKAUI6bxm3L9e0P6SpfDLyavE3vJTwFI53zwJE
xcE9JNjhfipGk0p322M9+RQ3LFsXeygU4zF6OmaDvACCKhY13DihFhWCXhn1BDG+EJAfvx6/akqh
xsO3QAGXUMWSg0WCQ02yG6mVUVEv0kREs2zU3/cIxe2L428UURlPHwuKAangR/rDUG9aGD3zHOgL
DUtgeKSip7EU/HOqn0b9jtAM5Jr81Kh4TmMOZbSu0xxuMl/Wftr3R79FF51BT/7ocRZqY5MaOPRl
LtMhKvGIxgkcFtgq5Lup3gLnSeAGRWYe2cEFoL8lc2Z9vbLp18Bkypm+k8Jgj5OF6cUe/IQBqTlo
fA8HjUpjFAgx8LauxtCHgJOCt3hdZX9wo3NJQOw4wa4u5QEHXMZ7PsorZ+6j6ARrMzEdKlLL5dNX
ocsbDzE5nfeT1zGBdbQJjaB6bjBjNLBrhYONYxUeqo32vqwc60qsaYIElCNQbDuYmY+HU+R6F5y9
kIG1Wu2ocSUda/84uw0s/jKhKLgqztSoYEyHuBa5106iGzyjVCjgZVmv9PsBgmijp3D8tYJlkIdN
rbNGrowvZGGQQfIe4ISLoLKDCsAu6a29OPHHB9neAPutbizMlqS8hd/0sDbS3sZjLAZ2jVSVxkZO
UlSmUOhigXTGuzotLsUVQmO9es62ZVBu75P+ub4xufe2xsVvLnvmxAgRA/pCerVLbYZY6lg4AwFB
b8oWoSzmFEfU6ZHgHZ0C08VY1TEdc4wmDHeSCmVCMOywFKYW3OtNo0lXgDcFmBFHIG2ne3KNrBgs
aLZyNBxWpmiLzIFxuLJrT3GQUfdKnhBTuJfdTNQiwuoZUcmKPB0Vhpfa4ZPHgCNiGxBxVQqmxFU/
+XbBnD6I1/0nQhZi6sCapb8X4aKfhlkz3nrRx6LNgEeE/XVpyQG/eTtQ79YoYbzEtKKOaTt3NnMM
11xyTeOikhAKMXlkq7djnMKE80DekPKPDFYC9IupWC2o1X/vluI8R3km77WuV+IpD6vUsurmXep4
DTZbqloO0DmO6Zmke7eNTZGWRFvki7bmyeRPzwsPDA6vn7TNqmCPwnB23gKSOy2cJUKjeXtMc9j2
FZ9eB0FFGd6WeZTzklrgJlxGGmGMzn6acszgj+3+mrmW5JeFqv6li33lnSgZu35bh9aFt5ZR0f5j
fivQzqpZlcCNgqPpnmFOoMAIZRO4pVyQLpE2pMfhkE4fHszqNXHXgChk9xyOw+WxnyBhPEq1l0dj
isR2RKzUf5QPmDySnWDzEZ/v0QyzrQp9MQtfelyCN19kXk23pjcSZlUAFLXqmAY0jSA4qvANv/8f
3tsYg9Kk8jJYtYj3Uw+O79/ljuZs5BgQ2euNn3w1s9/5yYokzw96Ld3HZpkHKeDScQdIyza+YA2H
E9VctA3KAkEECSZ8fdXI7AptoLZqzWNccVeVSvpmXFRKS+dB9BLgAyBrej7McV6g9TMBZkFP+Nxm
61A2W6IH+BlxNfuwERAwLBSb5YU40+6PKfHxXluwmfTlIcYlIUD0+b0fHnmn1SPiBlmW1wdecAWm
roblIVp4AZjcsThL4fdyYCrP4trG5QGHE9KC8qRplmKRyPkH09zOnwY7Z69CGKwXTRDAnkeCxIM8
p6acRMq3IyEoWMmCNgltr+KaaOqMMsKD3R6mykegBLRjtWG7icK8eA+4+OtfRXBwuyEX6fU3v+3A
uCGU+UHt7C4rCJEx9oYh3cw/toUBYHjXJnOVh8uZKJOzxG4aQaq5SDIAjU49abdilWXMrw6lrun4
uyWTTY36E4LyD7NIvMtludfwVPBvYDYgRDT81r3xrI00OgYQyEVQT1/qj8cUefn0/qJWZ/Qi+hv+
vrwSbG9WW2yaRlLjErkSTjD2P2ARkBEUfqtApgl7b3AheOpS8GvP3e89hPs1MnzqFCg8KS+k7tIn
CrANAyMszGvDXAUA9ZnS0o+WggaawMe7IOEvWx4ORlqgzONhw93dmAYW216jBuJW4hK+NHsnM8DI
9/ws2Y/n/n9HYjHLWZHAmgSe6wGmBraz2EGX4s4AVeZGVstuUD4KabG4inQIwuaIbk0ClOoNgxXd
3B/0vxnEYLfFnEtF6i+TLaeOOyd1KQ+P8uP2j1wDYz1hOAoe5ICb3WXci+kTdCl+RPcfprFh7+m1
L1QVpgOVD/RPMHL0zfnH62w/2jiuA5fmv5jaGeCthbHUKJ0pkV6bEI4YIGJqGB+n4ffaNjgtS8jo
L2tcpPeajN1epeUS1IiMupqE8mxgFrKE11rnLiZnLzeMujVE327x/pGwDbOeqk0JvWbkwqRtlSbm
0opfF9Jri9cA3aC9zCTTFPW+vsbvOe4BPewYKv6Wk9zaIiflC39jlEcjOHSSzQV6GjcDVr8wilpr
Fs0uUZj9tt5KMindd21ucew4t6xQDt3KPVe1zs4+o+w44C8wPumb8JbGFlJgNE+r6Yj38NOsYZsJ
1E3XdFWoIGKNf0fFeksv8By8HgeDORzs34Fg2kGa8Vc/OEsZYBXATdnOYR7Htcrb8puzXSBP8wH8
az8vG6U+3nORFox7UgeR5jnVY5j+mKK/6cU2MfK6ekAqoAhOKwMxJ4uAcyeU1Ufww3yivQ/lSdtM
vy8EmstESDqyJS3A5JjEbS1o6AFC3ij9+uZB6Adc6/4mvFGBqaO24k9bpcIujbjscXp/mrBXpNbj
caMbe2b9rVgZDeGTVaHMEiWCMt23VLFzvVCUnFpq4STjm1BqopdlTMx41tg2IUJVsK6Xx7Kxurlt
+hHshzuG2eDudx9lFTEAfTQ6jV1Vqe+B/DPpVMZdgn2dZpBy6pLfE3jdWR+RbJmKVHMsyjwBBaSW
uSoL4adPgbtJMXf+fRPOKYCDSBboSq3cSb5qpQxmSoIkASlha0WMzDu4PkycW8tDkbkZp47g7gT3
BHaoKGmN2mWlVkCDbfpxv8kEBmN0s9cdXbzdnMr/xbQ8ol64F1PNrUtoXrQiKrfmFqnw/AwH6QgH
0kM7BnR/QN0Z28x0aZTsjFh2wp30O1Z3VXfab9DqSEYL/nI4f4MbylPzBZyDKJDELyQHbtd0MKl2
ouWXkg9vj6A60n1dFvRBCz+ZdudK6setZgvSXpigB1aeCczE6zonqJjZBNi8i+wTC92pFsFMGzLo
z+NTmnv7V8qG8Q2AS63zt+xUW5bHXQs7cgsb4RKm2g9TN/xUixgeqQM12STatRYRdOtZFcP0Wt5C
ab+RalZq0bdYzOHDZpChuR51zkpMgaC+Obd+FMpLdkVDgLyCNgWVnbo9lFbL9/UR5kUff1LZjUXw
6Qfb1t3rVle6BYTTUKfRD3zIQ0dHfcVJDQHk8yKdhO0JWJ+r/llIkQxEZZZi3AVbX0igwPZK81nh
CxJEytzKIdZCYcElDgTSV3VAwHI+080SOr5YaWuAqZw+10rGHTH1RyJvpdgBrlNeTFIJp1zEU51v
dt9R6ooiNtyY6nxuG9Dsztp52nJrmIVCMpNyJCbiMFHbbOTyJDrYhxPrkPWbtmGmkyz75ixz8Xcb
xQOjDXyFumW3o1ywV9Vb/QrFv1YDLwEp7YcxGX3htvB7WgUeiyjtGCaL2R9f5vF7zC4liBIVvQcp
TG3DSa3mJgomrzkCVmQjO3tczv2VO7ZgiLgxA4Io808l3gae5PjudA9VVVcs5ieirZIaRq0kRb+4
4dgkQEgt6QOoa4tN+8BMWsSeCX/nsSYJW5XTSJFcBWl3kzboD0CBZ8KLMuF4bLiBUBSUUP273Omc
6wrs1d472srtNCUK9dgeaSJFjYjm5lZOYFNmiUGA5B9CzBYobCTnj/VxJSr0RWmyugh9FLGX59Da
6YOqdhHt8t7cfuWKRLMj/mjwgioSVFHKze/r0boU4636/QZCnJ6pc0NrdY7ffeaJ5IYwd+94DbMW
1/BzXzyoX23b9c03KcDwAuOK4O0NWiYDhz0jL3Kgaak7Z1CpEmUWSc4tVWXSTCHw1dhdrro55+bD
pGt75kDe4rhSVKRjZwSdzwJnCH/WS0reBrVC1tBMlx2UKr7I3meoY7O6yJNjhiBStCn6jUCnKXYm
SII7mm/FF/m0plVWpSYJioKPIiApBE1Xz7mut+NcXCoWL6zXJH8KDru/NolYhUHokiWsgbgLXPRA
cGton0ks1ccKnAbsZcxdDP/2Lm9Hph/jH+wUCYDCUeILzveLuRn1DlGikbnc6UCBvK9capn7wNGZ
PnXBT3oiYZrSHF+BegbY2iTbGx5wjjEAsALP2K/eOHguvyp+kMor5R6hSRnT9aBthEzpx//rmwdx
QKtPB70MqQqsYO3/1fp84aMO6sOLwGQChqyXXRsLMdX9jel+IHhMBdvktu8lk0rYDcPEtwkE07rk
Rc0Xy8CuO1gc/fyp1JgsbPQ4AyojRgaJUzqYEMOFRY056q++fYVImorI+MezXtEcGf7XsxAXUAYo
mmGrKx6O5cirv28bCk8X5e8a8v4xnIkZzIMcgH9yaKNpd48j4KF4GhLqj/CiHTONSyGpmRYY9H4R
HME8oAVB62mhLveQiNbTWP1/9H9pHPFiQW6eQBYxzymMIWiPq+EO7YsB3air0I12xWsRHAakIeIZ
GeUgCoMGg9UFnpfukT5hQ5rVBPj9rDIQUQmlg8p4oH4wKwbApt9IOnn8LA08oIxKps1Fm2/6QsiY
F54PPjpFe7GQXL6R7J5XCOi/34ADz6vyS59+/oWQqjOLJADwfruCpKYZ5wgUwgNBTDxeIRQRgWhS
u2X4/8xBMaist1Dyqvg59OBeU+OIVfSW5zG+cOWcZ7ikZUiszcJg3SdfGaYT0qt/htTZMOc6yowo
5hHS2vCW0EUGSVQ9219CLyN6Vvo+7ns5X2ae5AApB6qusVmtKF8z4uxD29b0cjGEz4Xq8W6s9GWn
zDh5X6FP9D9/cIv3OFojfAPw+AAK5d4Zh+JMRzQs+UPBlDthBnsJLaaTBWcy3UwINf/uFXFG20Jj
mHLb0tIj1kGGNovOjV7BL1EOfTyqsaQqWAM1VHvf8v2E5hcdYQ2LtLH+CM6tuEMBhJgNYU6cPGCx
J6tBLrNVtzGMMznnLdElnQ4u3h56XADM6iZGpXnQMKknHLTEZFLaH+aGaj25hR4fPI80Uzr7PMsZ
Xu2MFhfPU9chiw/qtiEg3WKfvOVjjjmQtkRX2Mg9OOZA1I0huGa5gHOxnX1cpfO6lr3Drm+mQ2QY
wWTyJhbqhrwCNyVwQNvE5GFWDxCHbF1sTt+J2JLEocazW9TZExUnLY+BRmuuG7y8Zt0aAZ+wsXcf
lGDwtevOevg48mgJYx5IHPd3uf2J3zLjMFBW3s4YhW0H8tLdLDaXFdxFvyy6dNeSaOL1Klozi0BS
gnqJoneOTINdivWhwp4vtPFGXCbDIJAwzuYuja1KZHjPxtZIAD2monnYPcMpnKYBXWZoQL9r/XzI
1AlS21I6MW3VyMlkjqa2TDPuh865CltlWCdvu83RBBfnBsN85UXi7YCAz+TZAzHp3L8kPRNj9gA8
4DZBlpLj+fGJdMMz9VW4ZrOdqr0AGGIdThh8AbL7mfP6idgKOLekdKTXsmAcGgY9mUKIbTRkyf+c
xJYKOQ/jm6Ag39ngk13FxY3qY/ucNNW/fF3GktZT9xUX6IAI4RdTYYdibq0IveG/a+bt1Nyu7yZC
PboUJrVZgDlWt5hIMDGSSzP4+KWqmzHz9LFWZBrVz5Mmj6Z/Yjtqg5+JbvXEqs2Wf8knfySu0EpQ
rzSu2pCD/BsrpBmUUQkIBEcVdoED21Z1neEvAUJTWCNqzvzcJ+iwEYJln/WV15LTiIznoi5OHEb1
RHZ81kVqy6k6e5KfRL0/y5Q2qdN0HyxHhVqhGjLdBmewdgCbXzS71ogl+uOAnlLYirOpTDvi2/YM
zZ9EAW1rhO2ZQWn4ceTAZjMhhWfuNtLG/Stpnsk/cY+Bh/IM+2SH9LR0kLkYTwmmslq2/dhljoV6
wdIp219dJF3OOdjxQxF0TmenCzjDBALhwypebGrh1JHNc8iOXpcdtkHdb4J74O65bx2oeODudiJp
j4MGh4TAdER6tVOo4PU8BoP4OHqGf2MRCDJjGfHuOBHgptJXREFoih45P0IsUOeyg+NVpEQ0Zneq
i1if/lBdMK0yus7+XRtkwKXickVU7/irGueWlA8MZE1HJks5v2tybs91ATM+k+ZC6y/pef0thcQ4
A2IPmyVHPZS8AurVNN+7tnJbgFCVIeam7xBSCqRhBVcLmFU/mitJerkH9BJlGUSCzq7CpGmHOm6H
nP8mAcoMvmhoDNgzhA4QQZngeEgaKYcQb2V+4orTJEWUS5bznQu4OKoB6boZZr+iYN9tMQHDtZuB
+8ubSopcseWNgwAoe43iVBn2jwrwzJb7blh85PLAhUqTxg/mO9vE9RIU2Wl4KIO6fhoKRHLV+ESc
ZBJwB23Aohfi4uBT2Mw0aZzXi4bFPbawXl0K74UrrvdqcT8UdcA3i11YqdkRpuovfBpfx1aGxzMk
A0DCHZ1RW4r690KknXDXWxgoqIUKOKmN7Rwvk83LA70aM+uJw0sqVXKZnBbPo0kX45xxmbCxH0/C
0ZW8UQgNFJUfNVfvBs/kAVLtKxe7rb7ctkRwoZ0O818SOk8lDIMPSM6ou9TkBd5oEb0yGX/wg7k4
IUq1kFXjGl0fb21wz2t0ZjDVOEVMDrZk9Fa5fvNkDWQz7g2AXfgWbcTCSTYLNUygKYZGq9vcHJm7
YpsVwNz8XE6EkC7BmIWUt3GvXDHAicZsoVV6z0qTI7PPC6xymBoBBrirGQw9/o0m1mZYcMWXkZA+
Q3Brr4BZsXMyGpczbeRAhvJdc1VzgRIoImtndaS91AWdXB7EVcwzc36xeBTikmUFvRgASiKa5TmM
KDHfDdtZPyYvmEk6yvhRlE/GjR+mgEsb6TNVH0NXmq3hY/HDnUOh2unT20652pC84V5fhQV9LRtR
5T6o4Ojx66aAJPvzOvziemL7hJG8X5Zf6ubrkhIEoEemdHDfXg2zH3E9FBcxWRH80oNWVTa+h7X6
fSxd7Aw+R+/GoxPur/gQV1A6D4ACwNVabOlZxlz7O1/XRocJv344PJlGignsKmbuIEN+SjZoBerf
blAwgERUD4j1Bp9fkoa4QtlOu4FJyK1/7nqjApMhQuuey9neAAufVmR+3BWPXV/s0Ts5K7j3TQLN
Zm7vz/MAcnTmg9I7d3P/nj+U6tJ+qo3h4qbbFvISw8pTD5BpJqzA2BvHEf/rjcpwv8ZaDe1hGoGS
i5wqOaFKUyWWuMfwvS++NORcwGP2Cdt9Iit1LzZ07yIZxYzu/U2bkG9xu95P99rBPJ3+4egsKJKO
q+vyT1KIbiFgbr88kX79YDD6gITN33uyQkB7e6Q1v7CxbchD6BRYpa4kRXIcwCPm4pA7lhHq2+ua
gIiSB9ARgonHrdWxDt1e40QMelKpNliu6/WWxHnc6tH9UUAKSJ4AuoMUHXbeAPdKrhd0DBFGHq+R
vcFV2T1CNMOC2ZHvE1Pgf+5AFmTtZppZ2pL+Y/NTYYeCx5A3p5UTMP/kCSbSV7e+4ORSIE1A1ebu
ICm9a3SUMCmQ7mn9EhLBvRS62zFv6uWL5Kxz4XtgdjIezY5LCH9f4EhLhmCMd0Rn7nsrK5rFl1SO
6QGxfYuzPaE/IKUk6IShK92uCn02AGNewcg/u2ajwpmSy+D1mAlb3vZPUNuHUH73mQClTGLFBCEm
yCkQ1wIpT2+s05kaaQ2IdQ/M0c3jDgeWlbm3b/rMWr8AZGGAQWa324FcromLSt4BiA/XFpMvBJu/
0izHRmm6cR1VDvWxTnIq4acThtDWb6DnvnbQLK0lRKSOrNm04J2IigpROiurHI8LFQ5897ZiZyNW
BM8C4NLaZ05czgdJfrj4lWJTB+pbNbWwexw9UemaL5RE6aTMUfxzubN8mneKnnBZ4snXtpmkJ+JO
PdiOuchCieStQUJGyU5s9rDVDNYKwOeW4Sxv2uXCQk16wTipk8gYtTc4E3Lr8hF1U5Rqueh5j/Ts
u2vhZxr11EvQGlYuCr2/LY/KmyW1+2bFgZwZtQiUen9jEuxjL6LTNpWLJkQaVjA+tuiNgtjavqbf
VDHS9iZ5CFhdoQeDlgKO7NvVY5ipQTv85Hr+yJwQSkqEPMd5wClnho/C0KDrBcNtM2cIxtpcHLPN
dtj53Yabmq9i7OQ6thTpBrXJCMn//vo+t0hx41aeAi9oSUuVcGMgKSMtzXpkdg0S+qcxnKRCdSno
CMyUNSLLaaClxwxlQdirRM9X44lE6oOqR52k3d3C/Gro0aH/inuQCrQtulgAgwkMna784vZOSjXy
i92UC1bdCymDRFJ2LRpvDtqPOFLfdyT8gQPJVJguZnQ1wZobLnKJMiManKHHXceKwKl9L/tIYBSt
Wo1zMczObC/kiyfWfBD+9aZfTr1G6GZFaqTLh1nv4dTFShwF2evS18/7WiPB87Hy2O3KSvBETib/
TrF0TqHE++v8+dHexT4rpsZidF2tEWYg7IVwrJn4sHpywVOunni04FVWkTfhHQfVeBRcpGUvYfvb
1xNcSZBhoDv7c1k5ClqyLlh9F5s4ixUIBCBOYNdGot8jQovB1eHbSpxJ5tdkWLtaEVSdxUSSD1zb
Kp6s8riWZbmDUdBlAVVKZyJ540a0TeJJ6yxMGaZGpk/5xdhIffPts21IzytMLaW5dDrVCyGHSZP1
JFpHuJrExNmxZ3pq9Swn7nvhyF0cWg7QQoQyqKxbXCcNov7VMElo2tsM4mJbcDjeT7O1IwACKht8
r892KBSMsnC3/VcJqq6N4mT51Eqo0eHHCE6BoQfu65ZwUW9G8jBDuX6FooIvNmrobXNIRMFyRYFA
Db/I9Zg9owoSVPopoKi/nkxJNTtHKidLj2v20+PzRggQGU5GBtfpfZ8pcXcb9oddOPAcBgFzfMGU
niJsp/N5JveHLWvYMMstOCaJ333e5uqyzfoExWCSw3gkO4GH6wM5n+6faeuqO9TrgXhSAy0r1PHS
mIWBCXeqT/VsnYOaskBkSAWo0MbKzbTG5k0EWWpOS5muw34WCKLoaGAghIqj2XU+/lAWQQBDyULY
FyO+VAH0+aD3mBfX/Ko9avWmAuwYOEBxVsSUkZzNcfQ+jGEgkrgqhtgSjD8r03qqpFp/5i9fJ2we
XFrG6JhsAKfASYvbVIY5smrqOXGZ7N9HmiTsSelVbjPsxquHsxD8mzbdlrW2Kx2IpvVgt8M5fu/K
iLUPp+GfPYzH4SgjpmxJINpK/rKDvzjJd+pbDyUBeo0UfpNmLHSDhT3m4iVf+xeLf0CE0C02YIo8
NOrsrOjhJecn26xoDAydpCpvy4fbfMAsDaYO1LDFaa59DF+O2OiPd0YHA8C1pioDx/ApEYUdpXgC
n97J8Z7J/0Ei5mn5LU7y7K4SY83eOqDfeZ/Zp7PFSRnaRxNE4IBzciYxXWAhGa47U+kfrdb/yJmG
75h1hBlza+vvyLgHGKtpHEibrlsgtqd0C+C+qTUNrxcoY4uBD4LQHhyO08r//GY2ds+l7vphuz3N
n5i1N3le+yxIDT8r/C+Mg350aE67hQwrRwgMKEBRJ+ncSShi4diC3iEq3UyzynGM7lKyMb1q96Y2
HnjX+mG3DfAiJvXhmnY7k41PkC4GN3sUL2rDjtOZ0MyrDkw/s1L3G0dd2u6VjPJ2d6OkqC9d34CN
FOGQGTQa+oMOJnDlRI1U6qzNImKMEZcp5J+ZsTOJU87x4wCtl+6lPuhjPDPXcclRUeemcQHfXRbO
uX/HoNZnv6q9Q3RAi7N6c+9sNf351QrVxpgwOIKmnfOh8BP+ExiyI0jpt60tUc/1CBEKUcGpBRsV
mVhUwwzEKht8wnd4W6KYRPcfaWgo0evuosz3/qDIqvflhA9bPZxGsS1NFz4wDt5q7pjt8/S+nG5c
+03Ft6LKn2Dqfr7YHs0mQCqZLHD68f0qIrG1Or1Cicp1gBaGifa0V7ek9pMoPpNtNXRhods5GAz/
WCMTJq272LeJWOhv87W03zl/x45qBTAU/3X4wl60WDfi+nRNr/0rHYH5pK5uSB2CRNMwpxIZiTUB
29yjO0YMdL7nWk6LbdOG37zq4nIvzf44/R90+gXRaHfFvNuRdP4rPehIRM2bPkvjhJNS+MAeSre6
deV11auFPCPp/4Nj2JuK95OpeB5rxjOI2LsC3aI51GULDrqK+/1bSSrC4ATl0dfBgTZHEtVINScx
nLhGHveC6BuM730tZrKfjPZpIHrVr2PdVnLecXMe4lQJayEKN2JHVm/Bj4LrqL17zW0dxtkxzV+S
lZIaT1NRQb6rBHNHk6LzUxqATY6yqBIPhUT37MGoorDAkQX1DOKQZmzEfHVFGJUd2rNAK49wcAZ6
awJSYDlO+TGqHDVOpZ2SQsgxuoKiQgkR1uZZU2PazV6pzoP4Ld/YtP+BkENZ3dzGParD3GOejjAP
FH9PakTxKhwuKbxz/8PlwYyg6wIB1Dqxn0LdU2xmux5SKOro1KM++bRcXz/3Dto+7/6lsY4oHQxI
D0FoEu1xW5idjAkp34gQPdvCu7DtjnrErKzLcpDH5DNVeTr1AZvUenCx2PcNfAVLMpLodZ1u4Us8
ExquMF7n0RkIso/vf4P8CmFfBbIV+Z1VoJt0Epf5Wj2oGspBkEKwpLxmi4GA0oDK26JfZMo1ZlkJ
Gg87ir3lPhLVN2u18QFPweFJnmflJZcuFWTynRL2cpYKrkQSHF97X5qqFJjEH+0+AsxX7QGsMV3K
pYW307qLuesafI/rDbRokIza/dgdF5FKb8LoBDw334EUyhonF34nEfNKxnxRVncZJjqYQeevglLT
+CngaJr5u5HzFKfjgphPy0IKqFLSh/nBpujPFLodE7L7Hw0yRp6GdlbRuzriOm2dJYKbUzZrxZip
TNngfIC6G73+GHm50QDqHi3N9hbGO/EuKIVUvdQ8zncHG56JGk6LBrt7aS4HeDdNmRDAIKcawz23
wZZ9+n2blrdL0aL+alRcALjcFsF6qiYrsFd1OppSURoeQquktVOjkJATZdCDVl2x3JfKiwUJ8BmM
N2XAsSwj1/tEYYKxi0SZE55+GvArqJ/Bq8QsrYHmvkP4JDgDglhQO6UkzgNitX6/R1mt1IbVAmEH
8nn2ej/oJ3Aoe8+I9hOWdHNTiSKHEFpEB5aidYBVIhezBDnxikRZ+sV9OXri197aiJ/ouquTV+CU
mNmIj7gCCOzkaRE1JdNbHyD1qEQvj6Aa5EnMBzSt9ZiRYYM4EJ7EO4W2qsG9YfI+NrYgtG/xhkcI
xUX6bECZanVUPvAnhCDM/Y4VXTbh+PNWU7WDzC5ZofffANdkxgC+KdNl2eocLwhm7hRai9Q5CWDc
Ef5SmraVfyhYUAiPLDsihJFaboO+7ZPOMm7ZUqty7TDNzMGz3jr7THWWFfdIP/qQkP/kWKGZMPNW
h7bjgn+M+MRyeTwg2w3aPkuh6ASFwbn59HSTfeOUK84VKr7cp1br77V+UfZhjst0YSNUOdko94r6
OXUQej18byv5liNFOrBkrdiXNLxL8m+bnv9jQLRAS8Qb8q+QTDzYYBX+h1JzoOnt8UzjvJh2kxdO
E38pxeRXRJtZhi1uETrzmQ4UFu2Tt9Axth1qM3csyGuypXqAO/pXNOidhyLRxlQhgrWeisrZwz4n
cPfYdsw/gQZYMnAy+PU1oVfQ/OT+PRKry7aDqgMNteU7kmJaUmQo3ykKGWONnBnWVDxAzZiE1pG1
eRRyaIO2K1aLotji/UZgSlb8vc2/YppDFv3m6uTg4Qy1WHy1QDkUDHTEvTVZMc/vEPFcSSUtEqS5
6hk9U64H1qUqj+CcXSMwccqmEVEinRhx6emmyQJVXU/S8kHcD2rfiwkohd8Fz0RazCdurGV6PYyS
oN9lGE0MHtdtR+hfTSawHntZdZN+5bP/zToWEEuz+BpVXA3+/byT3EqCVrbWfccApD7HveIiLuV7
DhNnXamYhQnVaGUVjV7vLouCFl8ZdfnHwfnWjLChrudpOARC7KW9KYH++nipDLIq5ORTWLWTFIku
8X/M4jvmdAApW7WvMWwxvtCyPOnfRfrJ73BxmDX7sXN8Yw33eQA0SXr3htxbhX8qguNOZHHIoF8q
e5S0iKEL2NjH9zKirYj29tFwCbv+Vj4zJH80ZrPLuvrMX+LujvTq6/QmokWbg83vZcyVIyzsgQtt
p3iK7vbL75MsLUMFI4kPfXLWAJgRLCexROHw5vaDwrtfItpHuccJz5KT0RH+6TZKCEB34Sh0L9zE
p8HYTV60ths4m73usc/jwXcF8v+Fm4Uq6hgWTNkIBRlUS2GT7LnKqfcuWK9OBTjpsCO8DOzLxmGB
hGtnhYXsOEpQZtEhTY8iVFVhEC5AokEkkiGMQYa84EbenLGUjeWWyps+sQCecVnzQrp73Aug0NOU
gRrPOZ40XnMx2rxrlPR90E+Jgfm30yy3kAUYtqt6YEY4PuKvC+d5V2uaFhAerZvImsoKGqPwboP0
y7dNz9X2u+wSod2K1Nnelpv4OIt9iNKr0Kp/Wkfeqa4sijw8pBDeE3Ro/5su4szf+Uank4RSbf71
jBAL0g26z6XdCzOJIq+rz6mWQlGlZ+9Md/STj2u3NicSnU+1rMMEl1OJKZFekwHKxpp9V/XSyK4K
l02NGnB1xyw21aTxPM3hxqQi/EyMgps8WLiKzcXFdZiZ0RsvZuugqEhlqwUR1ZUW94MK0t+wOfzC
xJ6ds5+gG2RIcShJeeR680l+iaLb0xjC1COhmHTRBTapeIQmUK3mGzdtmMoLRhQJbFY2PE/bRbDJ
8RabBbtl0aonD5jh/xhrf7SriuibbI4Uhi7FGNdFAa4pe8u6Gy5H5vhkHFMG6Gdu+Po6BOq+nRv2
mlkQCnNu8mnK4x2quWBWqS7/W/GP7qgw+UAXdmY3LMM5ih6AZwjs/Z1oRhzcpwuo3O5jv91Xx001
WVKdJE5pqtGP+zNA9fp0UBCUUFkvDyjgERGcG4Hcz5Mzs+vFWcVU1FaCGxWXI2nDObap4Oiv4ubl
D+6K+jSM71zlVpMHTPkNe0u3qlWzXaNNNYZeRoaq/O5yoW8/36QplNWvkduHI/I3WwLqfGFwIwQK
2sLMD4nkz00PkXCI+tDGCCZ7lywv3gBB7T3cF9iDj4SHi/UF3O7lswOXwF2NhzDEXl3PBkzIXzB5
VDyrMwJ0yydSn5jtTA8d72BQ5jyD5SNa9H+1cg5p0Vku3uZQEWBpt1gSNhNXldrQrYjstckKhUWl
Y8U6nmiJLP2oISXVwo0sG/+p+xK6C+7WGqwlQzV/BKkrM0EQ9c9drrl2xxxEalQPxEyyW4e9xygs
rf1hWqxmmDMSmER60SXq75lBJ/T1aemnMJFx86muhdLJuTXRWF/93vwNa4GZPXWMy3aHTiVd7Atr
omKLWyymgkmy9X+cZdH3mzMVX0zYjMYri9zZrR58nJ9hzP0MwVFLy+wz1T4Z+QwlEer8oGWWK8ud
dnfc9tP3/phUhPCzvJG8Og2yK2dYDA5MY29p8WjHppKLV5mcsKlnkU3Oj4kJtjzuOj1w9SugroB+
mQJriwQePxmapVayIJz2YTCG9Urk7/brc2mi2V7tNJZeDjLXuKVkWctTxtjt2oaKSz2cDshUuRfl
x1cbavg+8AeniauUYvLX5/er11aXOWqejcogIA72J146FxBkX/1f0e2OHHob7xi0Xw2crc5sVJ+k
wrLwrrYnrW+fRbGx81rXH1R6SQQ3g309yNrI4wq/yXkoeEQXHml3Smil81b4mCCtMDunBICIK2DX
UCqnaw+tyQ1NTSi7qV7PWcxnRoLGXfTAtcFp6HKoK5tiANLwmoTOgBn88/jCOKWfLVvIIjZPZZye
/gSLNfRyY9KxoiaHfl/lMAbGCoRaGEwlEY8uFobkS8AJ9WkDYXeYpafjcRqJrXlTdhuDmV+XBv7G
gVN17FJuWYY6iCSf1d1hgrat57xgKJEIXAvd28cy+om8lMJgh5S0DPVTP681uVlC1K7LFRRMsTqz
9Ir37FhZmgpBk9PIv6RrHkPAPFQ3B9WVo+jzqwLxTi/UXwEfyanDJOSa3cloc1KxdGj6L50fiQV0
jY7awrdLnMCOOv2auCxH/459kTmj4D2xryAo9Tn3b5CWAyTcybx12tbXVir3p9aigKcylJW1pNuU
5KN4i21Hxd1U8Tk2niiO/lXVvdQ6c2atWxqLQWQdmJd2X76k7nG9K+oFvfmIclW2ExkC7RdhiCLu
tfPyOpN2iUUZ80T6A2/xW+n5W1hZeju9gPZzxeiwYs9xPpooCzzIdxXAXLghrA+Ae7pJOJKhkHR0
iWCGkvr1iFBm15AeGbf2bsI1mykpo/jbV8tw6BBLROJ2TW65xjq8KpobFVNTOIie7vs2Vm0RQQbf
3SebOlznqKbXVYPXFZorClVisMJO1a6K7cLiB3+9sDTVRPZv6tqT5suRDx12bfiDa9mXeKUbTPE7
yRSaaV/DPAVSnIsrVZz4BnBa+C1uMKBpwXkSsVH+RL0ruigBHsJJZ1YnqVIl/H2KBaRxSoJcO/0v
bV1ESiT+q1zQkjYWC9YTX04CyQEFPWYIak0d3YxbO/SybkSZqUwgUlmP/qXIC9WIzOMAbfrAbK1R
ojtyTn+PaikCkrfTzxT9e0fpYff/6Q/yD0yze4789SW8nNpJN9DFV6WRhtJjcUAN2JaN7ibQwpZn
cqInil0Ra1pFBHdyZwRKlvrqRgt/RniGKZTNjxvcdDZ3fYUTmsNrP6oXnHVabgZJYASBwfb8YLZU
iuXAig/xDgxqtJ5e3OZdXIyM6UaNfbZU4uqg6X1wHc5hKZZ98VLET36LANtP+JjfnM2/fpFFhsP4
94cI8eczymJIKsb85kmo9PWSTGErvZSPuxQrLk3vCINUKJv21pusaDoV1oJXph62m2bpI4E/5mXa
ZWKYmEHn3Iop7d6d1U5vZfCKn8hbxhj2uU5sOoxPprlijrSKPKyxM1aD/TWmMtMEm9HfZeCc9Dsl
peQzRbiGcr4JiPuOwBvMJEoPAqBeXY6KSVfojntQyIGgwXMkVRVJkL3d2XWS9ss+vW8UgNCBNBWN
g/rTjmL0Qy4In+D1fXtvnPcNV4GSAXnaqAK9qCKQaDFGKIxQionQmrMhea/gVocjTPosaYf79oYL
0bPyT/D+q/EgIMmimVMCWTEdzgX74Bwuy5M+w/8nvTw/ZUciFPNynsCNg6M/99jPgnSjAQbIB8JI
2QT7U9v1LGCBS8eyov8b2QemWAwlsyxpf/V7zFR/KVZr6mUPTlhktRjHdACbr9khv/R4JzCUglHa
LbOltLpao25JsO1wlcyoTkCWqlLs4RkZP7aUPRWPmUEltX37IE5i/rxgSNfThPsuztpY5b86zcn7
8I9rk3PxdzYW4rL+X4El7BxxMRNSePgCiaUy3eKcrb8ymV0uq01vYOtsrez/ZE5R5horrkRLg/FK
wXyD8Nryhm0CT8P1G3zdVyF0XtDWvUycjvOWUAsLyKRZOGbw5g+vGdaUAG9IxLs8EXWL6w88TfOg
8MJtuV2j8fAcXHqnNuNxBr1F8I4vieZUZhyxGmnOSTd6uxZIaWS82QdBtOGZ1iFbrIYWfHeIxoYK
Cjhh1yR9oPdPBSARwNMX2CtKAQJU/E2vPmrKQy4tcCPcH7Dj8AVu6ofgcJa8uekq+1NUWQ33AhHj
PByYQTPM5ePdMoZffwvF910u15BlTYRDyFHaeT01C34w+1kTubU088U1FK9SDdVtv9axsNdF2N5/
ZZrDb3lR6M9h8xOuTq5bop8mRg48pyqmcvhrHXjK8XikABz2Ayns/vb0VQYsucL8t5Nt+r93vKK2
lrz4ZQLz2y/hozSPP1gh3wHYNJDRNlHu1fn9tD5vKF9QcOSdfw0v4PddxASkoenzn2BgXve7XjSA
aSGdw+B1M2jQRrOSjt7WZSRpZNyqtB6/vwrI+dBvV6KPjpIz9TIj4FN8CxYhw2mY/0oyLnKRROQL
+nkLlx71qRTc7QWyY7WWdmTzvdZcc74tHx33BoEv6QAFf8cjISiBtwFA7+jgMD1kuW3BVAhqYWDs
9A2c2K+jj2Qv4bgpkqM/3VATKfxT8uvcgsqfK04FScMPOPhd7hSMFjCb3SKmK6rc0Zm9iZTAoy5Q
2a+LSBqUH9U0cnK+kHh5ysKabNeQSKXNvOeVDth6+vZ7X/80kbIXcvBQ6oDa9k12ShumC7hKwZkA
PZImWphKfEVvrEy3k2DjglRojaYHbsfLN0vYWBejB4j14PIFuks6qLrvDftgEawBXOMSe2mKng5a
Td8U9zT6o+LFReIJQvLh6TCXQzT5AxPya4ircM9NDIQ4T9+rlUUnnV8b4Y6jgFHTyTZ058tHEfCX
UzLR++Y2/iNSykNjscz5fpI1XSql372RQyEDpKKPyykOTKaT8gCwRP2L1e2dtM9NXoig51qm5b8O
k30P7i/1QGo/Ct+MCqrS0L0PU457YhJoYPO3ukrbnV0WC6YaVx4YJrjJT55tg+u/mQDr2uPc1rkn
rTfi/WeQxjZOaSChsyjKZ/lanX9FrDZDp+XgzA3D39mGPmDxsrI3JEQC961jL911KqvZxPBh5PK8
4R8G6Gfgu/1od8wWBwBM9BiZemDr5RuKBE/DL0Ma5Ci+NLzcktxumhAFf+0jnquxVctT2M68Eejk
vfkZgOEM+74zqHEcRLDs6rqKeUGYy4oQANxcwonTOAp5W6r1wAmgH5do7+d25N1Hjneia5xdH6je
O5+4XhcM7LTDQ2dzRbY/ryULR75yCcWw4Vb/kX/IxYZxOADiOsnNcHerXyOVj7yHdJKs0kafmxyn
tky6IzJbi5H6CnMw++7StFijvV9yJQPnKIM2lDAf2XwIqOkxvEYlMgXO5U9KDfV5RnTbAcLAeeiM
fEzXwYuDBE6wQaL6cz0lARWmufv0yxaeELU+7PzZNzgasn2jU5lqEGZbUGKTE1Pc82n7jp1P0Nan
0CwwFLwc2hIOWj29s429jNEOkRMUOvp/nwxZGanyvaboQFNobf3E5oQJFf0Twu9C6YcuJ2kB28Ep
M4DkgxLfHVS8ikPdTd9nHBDUQR3SeUSUImrACK0tvg3Dxmi9jXsn0Wj7AOuwErg3eNgCfUCJMxpo
w59An4VaEXJzmTL6EemQbqmSSuUhu1G9syQnRyKIlCoGkyOVl/RUp5tgkQGPK/sVimSJDNIsnu1E
6zlG9TSIMpGOQMN/exNsHnScl3wx8TeP0mT3G52do/KNg4x5ICvrwpbL8HrCrubBFpYG4Zgp1HkT
hQi1sEc/z6TQTEPOor3yyNUL5osXs6OzllIo1mbnbLfgcCtlwE1AwUHZ39p/cexPv0zZyz/Pxp85
L0+Keo9mFQ0Lz0LNgVOY7F20bbiMyaPrnScSbpQU4zVlNXKwZm7kMy3YswuEyK+fuc/AI9VBqJHC
sKSUOnvfoCZkaEs2IJYZCaF8bxTwmKecT2Cfb4Rp7Jk1hYAtxqHjPuWE43uL+jj/g9Xfj83v8OcR
O5Bk3s05pTimKmGxahKdRyy2rgaiXCqVacFPDO2qU1pOceA9CvnTJUbj2Go0+oCQlGrCbR5/GFou
VcUUIwzDe91h5bim2TrOTWERYzMbsa3IntiSnaG6QYDlbR+/dsBpdnTnNy6zSPrLlyYcVW5Y8rym
bdWZh0z4tA8CffWcb6iwXeROJQtG5PIv9gNYgYPD2NzoQH4vKMZRVKKwd4LCU2UVIC4/+x/TE6WD
bwzrbqXP0srb+JWGS3/X6I5/M9xGkqDJmVn2XSs/GOpwYtFAFf0FU7pOwJeNMCwQPTS0PVkI9aBo
tFlxzIutnnAmZvzW9GWeMcOiHHyq//Wp0O71fg9Xq2tmgCtz1PK50EXiaTukoh3C82l51FqSBtt0
H0az9PseXap3ItQh9aTwfgHZSZrLG+ZuxD+hlfpAYyNk0KT1j5uMZIl9EwSDXZTR32PlIkE1GabX
TYYLQmUrwMFUqyRenqlCrJedcxXofBPdXId3jIMj0DAuHm7GLHaQoYsHJVUW6jrjA6mWCe2cazIR
Tf9aD6qBan/hUqX6AI7ByQ/JnMMtVCETHZwbmYf10vNa7l0CqoJlHhHdCCcIdA09VdHfcvwrpiBw
aJoDxLIw2ag0CXM+QDQIZL4BNPArkPGojtusU2Mrb8+EkDD2i72BrBgGxYO+JrIF3GDZEWGP610o
zfcR0NLEzbSDbBBhzNrMiz0eC8a1HOlNGTxwZpFiOKcvAgGFA9fRPLvCZOeGSpJRuZn1/UE2wzeB
IsqTU0+FrVNnjYh5FKZ0B1MoaaZhmfuxY+gRUnahJ/qNhXF3m1vJH5xCW4+fWe/CK5j2fgZL1yAC
73Q6fHFtJT/eV44Jpye0aKiUJwHknfaIjAHOcG90el1EGVmyJLMyls2pKc0HprhXdTtUrqTJDKre
OzVKykrEC7+xB5GRG9jLqw+kG5qIbFm/i99amZ4GKw2ZqIh/a5Rj5mevNYzYOpWDny9o+zbbpY1x
zhQa7pe0oFmEAbMq5KieO49FOztqJzS6KHyBvlSzH+frG9WtmrBpDT04E3Ohni9K5yIqoDwJd2jv
V9SPyMFfnofUZ00PH6w9ZvkU4b95rnW65So7O1LHK0JwVtlTKSDFka+AEFDr5cCs3pDokqAQSRys
+ZstQ5NQTds0FUUsPupKyB5b7q8UQBAc7BkS5pyKWrxs1TezOACcwjn5M5oYzvY6H5YbCP5BH4k6
8PWme9TmOwkAe3hJSX2oUnNzIoFwMLWYxz7yKfQRPGsPO/NvpXfjTH2rZqYY1PYmCE1WMPed79xw
+ngSBE6W6dtFZDDilKAP8QMh2iOcbRzxNEsjQmA/t8VdTcjpivW+Ud90Uqok84i9ahC1eYQcau1r
WqFQB4fxh4lH+TbZ3zKD1EIl1/gFOJZJ9+ppXKSEYHwEUhy2BPu7ZAcZ6K33kE2A+EcLlva7OBhM
kYbzTYsfUM8k3yTVT7Qf91gQ2AGo/NsyzWLvxLGFLfXgNv+wEEHTJsf/r2b4LQb3s6BI/cq39g7R
T9Lkjwg6EJCSTuCeYElVkJl0LH8VYHNGlt44iC7okEunjA1V7xnMGC4Oqve0OXyEaNcLkUQXBJ8R
9kJvicY6x+9Bp+6Fd19NddUfHv7bZnBh3NWCkk9K5wmBa5V0UGy/Vo1Oz2/xFGcQxBf3x6gGpv5j
l9EtfX009LFeoJ28ySBF702KqiheR0+HvBn2lsuJvDOTVSY8QtYpEjUBIPBJ4mkLlbfW2C2mRPdm
TJvtUu7yhwpj8giN9RN1jkt9x/9BvgR4DfVb2UQY0J54W2D3kpvz/W1B1oodRrr1M9UQaMUxmHPZ
YxQD4hF3hE0f2IvP8ffRWFcAsZEHYzQV9On8DitpP5NqDgvHpHlWdUQ3n/NdGBCGSfeyYwann+Gw
fDWSONIt69eIRYLmziV8cH43vp1ZsQO6zAPEURSLJl9AclNOxUTYSvdXy7kybnS+AxdePBNqBmwO
LnySkg6leyrfRfzuCirDU29B5KJAij2/G+KNGXQ0tuM/VzFC3XOajbx4FDdmEuTjkvd5oF8JtWsg
0QKw32sGQ7p7mwBjMjzgHsX2Y9Xg6rlston0v2W90TF+2N4g5vUIWdCb9A4nn5HQzNbKi4rTa0uA
g8BGuebngBA/RPvUG8fo86wAz5GpcNpKvSFTTrtrjEjCfVjxktRan2YBtDMM9b+yABQ/fYSnH+bW
1QY+FpZw5f8B224qr5mrhWrW+cygTRjjrNq0zqd8FgAKLLl8/HFLpGHQomG4RZlF/NYqrNXevcQb
blRD049xClY/TQLX2yuFcAcOrR140jrhAw6HlcvINyrwcrTOf2T96paqmZlm5jzenhArVuVYotCk
sE8gHhmThHHlVp5lh+YbpaPjRbEygOCaWwsslZmLh0zlyGwPTH7scWwkitE7YuvVi5hjsOVkiehB
oDWOzg5tszagmZy+oylnizZGG2/kQGi6klIzU31A1zqPPyN1sH8tOsVe3okk+OAzx0qAxxDUKQPq
KqO7bqRAJKnqTWlvAFjZ2KxUkRWx6P75G9en7I1whnLn5OO4HJLNkPAPUI91K+5+7fTR60Ag00qH
XZXnKDKA5ow0eGwl2fiWY8z8io6L4HkcuJx0UHhZmVpBHAmxpF3B9FYAvmzZYvfFVVA75NGpo+zv
OMqplOopCKmCFw8anSZi6UCBg56WGCUeBYynWUKnIuwGNwHfw3jH5ODp/MUSW8hGSU46UNTR/h4Y
EueHr09vijcd5N8FkO5TUjX6VT+ZLDBMfxq6JaWj7u6IRZe00l1u7B/PNYmsHdko2xCZ73n0VDWd
f5KWYRDNq5VsMvsW5O37VvMr9InSW+9DK/LygNv1kvAyP2b55BG+V4zFNq2yB2k/4mCakRunkN6U
WToweLXZQWvOcRo92BMDY88Cbe6RrXJGLcVDTLEJnu3jZzGI7lCH/P8HEihSIGWZV4103xpXtjlY
pbyOqnHd5WHmpfe4D9p7XQiY6jQNi0duxYZs4lTgmwyBzD7kLKb6oGzmZf70v290IR6E0xeEdzHq
xiInZ97nurkYexSOXLWQONEhTs3MeXf0l9b1rtoT+UyrSirjEmCPgXmxxVATPrjtwe9pYLYFQIo8
U+DonkiHyu5ojaZoeshf+FLljiNXCrGVYfWJVnSV9KSH7b8sxGxmsq8tB5AMuPwrS0wdm287nR/w
MePbtuU8NHD/Otxraxces5XoX0/651U8h42wqEP3sl9FGGqkuO4NBLgBC393HwruKdFv2th2oow1
Glh1lc9KsIFHexd7ARsEn5TTdyjireDlSpZ47qUzCiHmHQOuvXUz6eup6aMpf3CCXq9D4ufC04+S
FVCiCS0OoF0YX8kl337i039LAw9rKvKNKWku7Oq1Alx3+5E5+F5vvM/iKqckl1Ca6Ez1a5A50GzW
VNIWP5J8Q1kJT9EBospkWv4DgTdWI22sVLo+m48eWuUAZEJ96jy00Rj/S7nkTGKSbnEBhiqrFqEz
bMOAPu62BbPV5+3ayUO4muRm6mySgbsHhXkVgZXsYh/Umm3eQ0R7vhn8gyO7cNJ7mFrbwcFXI7hk
0e+9MMe/eRo5EO1kyZ+LGuulXeOmLQha2dKjkfar+vBlZIguWSu0OBM8fdZIeVQz0mN57Lsuoj6Z
LHLW8TSe0ynHrKSvQgyqTbH1OePMaJfWrazlCwMuvVdtTGzS89T46ypnPtP0MFX2LvenVbHwbxz/
FQL0LcP7e+jZ/LugzaDkAugIPrkulXJkwG2+gQmF4tgaZrnsS9xyO4cEFHmjc6DcpniKtb0RZD6s
Kb6/yUg155uF0InlWWTBxmmqCyhBikj0Z3C5fnY5S4B+Zmzm12kQBJ3DJaM16Ay5QwmpzRLO1qJa
GazC34hmhqN1W7vCY3lMA82mk/pq8rf4RophsgR+jbUq/hWleM9U+9QToYpQxbD/FPEjCUkGDVkE
9Z/MWfFgcJweFEpsj2WUpVJgr+Hbhk4OzxziFBWRaIb2fuex4dpGuP4NdcDuovpZ9h8/zOn1S0MF
G8yVaTT4e9oadgk+sI7rLjMBODb+vKNal7voxFZavnjCr/zLsi45wdHShCPpklShMQ3oo6LY2S3J
AKtKcwWPYzm5FjhWDzhNyxUbdIf6hbeoZ6VRxzveWle8yC3qUP4zASeHKCb9w9NAZen3zMXq+VsK
GBkbsah9KTUBNTMWv7WGNQNOFsCq1JiAxQdwg4+vpA4goxRauA5JIkqn7zqmW3Mj6z0Xxmnyjh0K
jlDZaFV1D+xS72sm6Rwzx0BX0SLiMKx9HTRa2h764aZVAHPtx15nbkG9vg+XAwrVthH1JmDhH8rT
BD1G5E6KQ31X67TaYPgrkfh3O3TWUtyoYsNzrJFJbvTIgg5CapIP7GAARrkgfFTu/Vm+m4WWuv80
R0YbKeaSz9I7ny5/RxiZKbOUawjv3kWr0/AXcG9hmL0jOF03GHUvEY9qz3BADBPtlTJouMOJCd/b
xyGEfkx7NlimFdbb2Sbql9SMENh6XRrxYJ8RnYhhKZBq7PHIrSr5GW8PDsDkShkfs8M4mqCPBaFf
ZKJtbFA33b/YFcJgbJMPY+j3DjHsAOwn0GIR/ouuTWF1tLbDhrUnbFW01S9S4tCZXiU6yJtH4Kb6
rZqZJ9CK61Mz4HQCS0mSIKAA7ogw+1Nv2/sBWWdxTrdzYUjm1KeBX4NcjTQxxi17hs6QaiaM4JQk
/xi1u16g9DeFRvMUceRavFyr5IHRgWcU+abeiPCIE4cxAvvZwdoWykLZilwKFcvbhJmgZT2Socup
/b0s+y2JOJLH0MYe4O4vwhm/g4c+km7IUBQhnUaa75GQqPrI4kednaDMhffhEUADxGLiWGYmtEf7
gX4cEfP8vdAbDUcN6KT3S8LjxhwcQnjjZR4bKPfr5vGDOJ07gt8howl7USGBqBKndgDp7WvOslmW
4SBQhXGjYqmhxOqz5Xu4N2q40hV4l3XUMTtJ2DtMte4wpDib9WG+HwdNlfA7y02xkC7MfkbcJp3n
no+C0XRtzPHUrg0o4N7XxddxdhzQcPHGz17TQNRNHQjoP2lNAJqF+X1i+TLqA379v8nRNPtIFWv1
yQN/wnZVpwwbeRKsrPr2tnkvpTdlw32YKHTHA1byetDmQGgr32Bmx8SS6i3sopvrAMYCU8OXstiW
NJyHOREzGHkuQRjqrXOxr/bQmmlgsH8u0Gs69YE/Yb1IJArQdhnbRvslL8pqIv+apblp5xi9jvMr
fsoYJs+y5VV22uuzbMuHm3/2i1KrrEp9rF5t08Od2IKd/KtVA2BAnGkKNcjRos7CgP+p1XYMTUQz
319+iTu04TXHcQzyBe9xKa6HvAJ/sEw1Fnuk28sQH7sjKhWmjdNUC7N+oEo4edbsQjkyQ6OR2QWi
1ogiiIkbX8y0tSqnyywRfqzEr78zVF3Zk7kjia9n1sVPSwR5xXsOtzI14cVVIfQRCpZ7UyrhV7SF
wI9HCSakwvQkOhudByZeL17cdKkz4dspFY72p5zvap9VCtR+vT4bM+6JEZasvAaB60G2twA/E/E3
qRS/EC0ejrr7URCy0JaloRcuo0ryD33oErma4cYlgFQzUzi8CBv+AQseT6cJsXvDNGvPH94HC/99
B8p9jcPgVO5kkXD9IsFWZcvvXfU1OZDcq+iTRdkYaQMq8kzhhHqYr3+s5XOfhEQlD+jKiU/B62L+
U3Abb9NTcPf60Fby5UulImjx4K+BP6ELSoGwzrdr1SksfIia90HnSmr4L7vbaRJ8R70Pc/EjO9Dh
a8I9A+KdXS+2e2WDLNkYbMk+l3oyqn+qUC/2JxWi8KIOoBuB5G1ywQyDQefvwbIGhgGis0DBf+Pv
BHupzJbzLI2M+BfHQJ8SRD0zrzKMd7/wnALyQCy1Bl1H8xbXSo7XtZluJJQPRpRO43hpxyLv/wMz
uTeojtNq3LZ3Bh3wRcgivq6CuZE59QjikGjqvK5fGzbXoYPn5YWIaIkKBThnodB+muzv4IKTLW1b
HHv69/kLTqVtQWHSTqzRj4otdbucDMn36fOJiyTgMXrJytbqwdyS5EE8+fdsKPIQ+OgutewTZCEQ
odGuy4w8KIu9NPUrVN6cyLFreVD9GHMmw3G2ss4dwNrGrfZzE3NSKry2/XxQ+BQ33uNUSvtCrNBX
gKpyrB91Pk6jX66m+tg+MBeej9aGzO0/D/ygW7ak+XdrngWweEbA3R4kZ6yusQ2PLPokIeY9GFGb
6MTlxMpIVd2ywS15HZAHBSh6xuLdwLKRke/jn6b2TKRQqSUrP5Ah0fNj/M8zE0WqBokFJrVjo5wv
BgPfHnET2EjFm+pwbgoCusB8gqWtpaSUmfhsE8OOherrg7x/9N0o3zUAve08D6ivMRg+OJqI6ZY+
+IctRJcfyIkp3Kjr/6aR0c/++Z8DmdaG47X4I6nwGAR78vcqTEv+ojML21xMUVCuWs+apYPUSL4u
JVlwTSYimnEidlX2CunPNk7B0egLHfao1Z7Px5zvTP9QALjQcah/LCS1krVhm1g3Iap2pT59wEKW
5+pdYNdoj+Li6T52WOdHs9vGzQNWMwWVI6wgogwudlaWNMccjUxB61EzQPFWlOFmbFebznr1OaZA
O4EzmkJVqhhqSYHotolAoK9Otizxx2NXNN2FPBlCkwx4F5LgB1sMzo7WZooI3ZNLqWmJn+OOvOHm
kUGuHexbYoNYyzgoEnkNeZOXlKFqimyzVUO/N/TA5iYQc5c77uN0D6bG7jFm+UIozTb66xLc6uAn
J721WtSH1i5Rk4tcpSPaPwac8aIF9QFf70dqZ3pRton8VYwjD4US23ZBlAhA/O4+xLf06wIrIrEt
BKJGU4HOjQgp/5J52B327a/bi6Pytj68SIfzyX62ndamUT7czhd6qqW+zRUr/VYQrCL+Co4MAPto
GISZ+OS4IPlT/y0KvTrz+nB8Ohq4QFBieYdI16wqA62PHFj88hJKskGV3SnUC3HpZN65msKqsV0v
OM52kn8yWxPBKPMegSIC6AK/MUOuIFjKxQtAPVt4zkmTusUvfMlc599rsdHyP4xRBT5OCiX03nR7
nnLMr+mFU2JkphKAolxZF9VPf4hVJOOWHdb/85YnGkXdyQK3yy8Z1/GPJo5DfW4VFFWMR8cPTQZQ
uw5mfNKmp33IsKt4KfyinHmvxR0jF+O1+47vCQqqCb/2SYkaZXpDFabV5dD05eLgNHE8ZdBLGV8l
kF55N5+PDh6nOaWxgOuQcXQbC9FVBCcElFdI/K6tT77C+wA+EEx6tJpWneWraMKwUxC5tCrD/AHQ
kJkEbF4jRSMyT4sVDbdyBHWqBtaaz5jRNDPsMvo9CNm/2L2SkpUBqCy05ijL9f4t03SZrvCnS5jG
NIaTo0gHlrSr9pnDHyoKmpiWBD4KEk7jeU+N/Wc931IafrIzRyJkfmtAmi0SEghprjnT19bcqQo0
/UJM4RPnVwB04JHVK5zmq4VzhHdFOVU7Fjx0XFfJsgTbqy8tCfrry5nwnlrj0OzFDNn1jsAxFNd6
98SfIzQz3KeI2hOpxPMLurqURs2iHoXZUk5k9H7zwtGsYYPkGu9/YwiOu5iwXyxQ0/Uu/sbRtMW9
eI3TiOHlquImOb6D9OsMpyqXlfY5AoqMgMljsSlcNf6UL8IJxtSW4a/uJbYXhRIBURxFJhz7UdA5
BfoRiMLHipPUPgje24sVko7Hp0p8k7u7gZZTFt3g9k5TPgjKdhzPVSR7SzFM2VDXAsG0xmVC7xDO
1c2rUuwkCROorATlca3jVwjXZkTWY0qpUNNkbK/sORPqh3DL9cnkMvVCvZYooRFRE5UZv2hv5tQd
Nz5H0FV9WAN+sP1t1dRCS6f0XZ1dTygzIf2++vNcxeL25KfURHA//C6DoJYYiK3oqhWMRkBTwzg/
PDylqM+7w3eDvyMcPoqK9xIAt1qq2ZdDO+2Hn6I4jX6sOrdxWMBu1sq25n896KkLV2fx7CrMnd4F
yqkmsse/mkEk8DXjf5KMR02q9kBDz8ImFh2RaaheVUWjRuGojkRBeRRtyuJBCCCd4dizAi5qPLKH
e6FycnJwyQ0GB5kJ57Ftqbcb8r2XlF54Ae0jjiyubsYhtlq+c3C1gpjDA9X22+iFmBD4QVsWMWxZ
89nHePBvXQPOTHcqPuO2RVYpaZL6pP+HE5/ba/oMrBIjCtmPvpb+cxKjxS4UObMpVq9CxxQs7qjo
NiLUYTl3bGit7h+YSZn08nv4em4mPLL5IdBCco+cN7g0pU9W1lCanpYvTvvSvx9XrOItygB00CFD
r9TUMny4aCzKPjqdUZJMpIcRiCcK/MnZkaZ9v00zYy9eP0dZ9oaKsLvwEUbwDwzDISouiNJpvOm0
MX/7Fe0UJkXzl2NhjokRA9u4TlJJJBXYIJEpqCCx3jg7cslhtsgfQIPW+hX7EQO8xyzcLgrJ+TCV
WIsI4KC/rtrv0h1i4qZ5lhGJblnq6vq5IPPt33/D+Ry+5f/5SBrymD62utWCrHa+BxW0MbB+o/tH
kb53T8JUcfPp2aMZIlf7FVu6INdvVkpdCcuvt0/ZaKOm70HPJd3ptOL3Md5mlnQEkyHbFr+xypgI
fiG+FYfCLlJKhtF0n3U0fky/9SUsxvgssmaD0OOrVDIV2UPaMfYz35vk5suy2PkS5tZb6mprRXKh
wOBy9EbPNLtOiN9FETj1feZLB2mucsU6kjXksYxDl280Z4kWJDu/uj33ymaX64imd1jDbncFduXW
vMNfkiOva7V2swDxJ5+NNfT0wwZWXIAe1fYFud9l2rznPepmWthnsWY6zUmmDzu5vwoLoxg9ZHCN
iytdP9opT7YGQT8+36c659tOOsqhlv3Umjx9JBsS1kKZrnEjV4WXJboI/+bLYfQrg/RaEUhXX5iQ
vOq4EzDGAWSuh4lIZNbfjm+23sWYqqAGxGXaaDXEwzRg1y3qyDPD7Aa1cyv/NFKfNH4MqbCZlboH
Np+kJhOXW6HJlVPSZYQz5QnDs/cCtWNLP4gz58GsMitWUnS3fLUSucn5GNGO0++f1AK7kjs2uqB1
rJljufJCRI6jAC25wt5zcQDJ6t5oTT+4LemORykjSy2uruc9CPPWzw9B9qNw5mtUoNTF7szgtYBj
iZkEwUqBSpPR7BbaxMXoOynnTdRP7n/QQgCvbWlWbMalz/JFP4rdW3U/kqRthKOTw1OELgE6dmWU
fhln+T/AxAaT+D5wwClFznSPsrKYFcN/blP6dGtyFG+vWZscVMOM2wSFhsAasc8QfpP63vqapOLn
mHBjdVgDHHrXYi/bBn/uKRS5W9+GKi9W+jItiUcG1sj4Tzr9xs/V3V8Z8Raiswso/OaeKJbqBRcJ
9wvrDPZzbSkqthEHGj8Oi2f7cffO59oWZZfnxd/4D1TZcncW7DXDcqvc6hZBYoY+L8k6S5O3NERK
yJKM08FXwJOl3RTDReqqvlZBQL0S1GfGvhmZiE6oGd6C6IUBBG3FEZkxwZE3NoNohlH64EO3H070
GMY69yNlCNe6rYlQm6pBAalrsZBmIY3WyFKqm+jb0GRIua1DrU1bCdHt6+8lltLNzP/jLinl1h1D
AtNCuIzKbe6V/PuXl4O64drO0w2n0YUSHk3upx9OugVEW1Jg3A6dpmuZXvnxTQ+CtEb/UVERPNFF
VOXwyOLcl3ckHt1Z6dkUYxQa8JKw/HoSjSkb+A/jjlr37R/CGchdMUj5OGCqkU7YpPssdn1ka/EG
hOLvkqnr+hedl0jFzs4iUyfqSbOlH9kak7eKWJMHN1BRKjQfEZXc/brjzSM50dTIZyxo/0On4RWL
iOPL8lMH5Y9K5YI/ILQoZw/1oqvLjK6CBNHnT1HWxUONn5bv8OatIgLK1OICs9fPhFDXE7Y8UaZn
+1oS2742yO5hbMq4nT7WY+2q3uqShMLVowxGal3iaZ4YqnWrT1ANtAOzCWbWJ0KEpNSHPDEvksG5
AualHgHGPL6EWOheQeP5xb3JPK5S6Qfdj10pWlJtk6+j9SXJh8hcJX1cTVMBZj3J3cseBCwWLjqn
ot4HMt0GjL9yeR5WDClk7t9WI6oHBsm1ZRsNGtE17Dv2ZGythqN+Yo+tXp7bumO0cLaDpdmE1S2x
QqTHSKmOL2LXWiiw1T5QkgwMFva3enqiToCuNUwXsK+U+zbggfOKHjwpgY5n449qjrRioYgNASnC
FKn//i+yxRpTOpKBveCuXa1w4bXWyKnTkd1hct7IqVvE5zRmnQYEZMeAk+0qPqX/M6Y/zxWPjJ8M
Tmc5Yfvxg+5oC17QgI4Ri6Hamo4Hho07q5nAj3HjYPa0Zbgd377CzvH+szZrzKr6C/+IPkSd/Cff
/cB61n2Wx0SbXCWhQ6lSyqkXY0kNd3MrhXfTqQOwN7o5lEq132SKd+s8u8ULSTqKGw75hTtdrr1a
YkDTba8lG+M7okqgOiNKaxBScqNXRN/Cm93uaisZwdSkq20yiFdM1OL8rT2xcp6JEOHslFVNT2gB
6YgWIecEhBLjsY7vWbyCxMq3JxWrq2SGu2bDMW5IQX8SyiOOcxDZOSVldQXuxGO/67f8QPgOUPwH
jKsEdTLG5JKdXjRTSAz3Vdi8tq5Kv1klNVtYP56vfZ7NfPI1haudCFCcZT+mdt1Qy086c73Wxkv8
ql5USVBApZe2vSDaCv8vsXqMEMoeTWzYn9rBMyblnmbJ07Gsy+W18HvGK/9dplElV5WcTU4Kmm3A
eUCceBzdOKc5aSayoapLZGKYiTQl8VEOBYkmeyK+Lu+jSdGEKMLPM4VSWm4jGw4mzERh4og4lmEX
rTSbE2S7tE1WhdGnid7S/JilhKcKTu8GUIuU0pz+a3QoHd2BTeV7ACYTEp1SRdsh1Pl5ng2A+B6V
vt70KBcy5OU7V2LNT7Q6rRYQIjJX3MjyFaXrC/BglCd5PZb9fNL7t9R78bhbeGH8qpkJYOPI3uDU
XY2zbjgJVMPC90csUUpg/Qa1/pVxiXr0cxOjLg7xnTSoOQ4MhD1zn5pb90+BSSB1rhY6qNelKWl9
b8LR1gwk0o9zKsyGhock0HhXfQms1m0P2d3INgl7V0GYOk53XSdSOIm8ap6Ft+R81VV3AaLqJ7M6
lN6IGLmjTECcvnHLHKEOth3dJvZ88nSXbmgogW6E1q7tItNzBqNH/ZxHgBwCefccRn7nM3k6TB86
wtHYSHMm0uF7p8SysjhS7bn3p2kuHDQ9HGJqpB8xQSdK7mvmQUVlXNPKse5VdLGZnzm+R6a3yXri
eABK141hpq3a2Np7LdV6JgJVP0KXUdOHgUIenpYiVzlFpDHemTKEo+yb9jkMptRp1P/ujw94OJBZ
+0NpjIMsdh6LG9AyGbZJOoJYkiGT0lxwdsiF2ZLPZN4WxrrB4ITXf+S2ceoI0qeklrAoF8sUiD52
ePJZKyl99UzJ8K7HuOlMV1EiuM+IwbDDjwZ6PKcDdRTnR4Equ5XeTajfi6dWVBT/3gXxOveli1M1
hgQJw2dJT40hRnPQN6NQqXicTE9dNkpXDTgsdIn1kLpwb95uIiRTDR455e7nlSm+EskKdb54DYrT
6or8bHdNtAPQ9LVFPt2hY19aJnfv2Fk3tC6cQc7Fq1BCeojqBUVtlS31fkuDJMAmltIVXL92TfOY
gAyLKjBmpveX1xUy6Ha1hJHd8VPFTaTCZucCHHdxvS3vYAlxoEeX0mtg1EGYxBtu9uFsIWilJ+Hl
p0QEbmpmc5yryiNc83CUyTQg06gpzZqBT2urewqRtgreqtVfDtPaP1eRRb0+DETic6LB4BzgrYpl
pm8SGEIY0+xPUz/jKxD4uQl4W9QiXahgjeCome03gDaBKCv1XId4ruk38TjCNeXUrdpux15Z5Dcp
+RFTNX4R5X5pSFfJbG3x0WWXbqFAapGXKEq3fjPgL7izONDdbLsu2ZK2q68aYig1IOR7iUjzS2m6
uR+Rzj3MTQWm8d58dOL4OtqUuwa4wFZPfeI03abwiAGJcQzelVOQX6rmRZB3cwRlq98VvxsrgqKi
rCAAIxwCjFlac4SrUe9cOXOPd80/2atOFj6wUt57qMvHG3oSIdYHpUDxbPOJo/zrkT1aTW/PqzDL
lppxuoKbomtoWXYIchSJduATP7vWHCX+PYYysENY3lOPX1VqtKxo7RITB2qTm6/adS0X/31wR3+G
6wUqyihydDVN9I1grYcTE+6n1OrpyAF0pgIeVQp07O6UGNdMGV603bsj++rYsB4uasCsYBsjM4YK
+zRQnPu8Qqhqj3b7hN+mvZfkvHUPEhN7/cXHCY6aaDzJYT92Nj9wysN0Q25rjq0Bs8DKAtunFivP
tvfyZ99gPRifPM8ld3gUGgb0ZhNFayEK2V2QCGSOcpgoHdfxyInfg/4ZNsH5avi4yRiPLRAtcaAF
JAEIehZRUFFO+PHUsktb2KEXFVXj3pQXpyf3xiSuxLfsznb9N56GuOCoaEaXZQdAo0mJDu3OpDht
yn+yUcB3lNNDjU4fuL8QpdUW+cVt5rU0P3S8CKajmXg8mzr4B8sKcL8BfktyRImaZRm6ma210+p8
cDxO44uaitAkSjgtkPgpj9j+tD3BvOoehJH04GcHmsSlrRJQ3PjKEwwMl3tdGKP7f9Z/Bsg9O0+8
LoJpkIAUAIlVZJ9eGcIRvCJBdYcrSlHzNMxj6rW3y2eHMjAC13Y3H3yi5MjGScCpDy8SK03UFhIY
220CkweOc3QXevaqPXkCcLsOe4SGLAMb0SO7eREinjLdoQnckPsVICR7wtyc0kULdjiwC/4s2nLX
p407sM//PLBQ4qeTJuzqTin0q0IEnLsc3H/C9ibFSddWa0D64HYPWWPxfXPKXK2aVnKZ63HHzCYO
Uu+ZZbbjUQM4e4VixNUs1EPRSN4WVCz8RJwKwdcmwrjZmJY9hGW3TaHqlSIe+uhtjrZS4EenPjQF
ZLAkGflMI0poYuM8uYv2h3iyjs/xM14rqsCnrAxF8hDEuq4fi0lts3Vdz00I6nfpbXhvoZtRBHzB
zYer47T3VdjrslAqFDWSGzmhT1aHOcQHjiZORRnkzwL/TgLloazDjog5AkkjpmcVVweVL8Jyv3xB
HAUUcLSmK1M+KKYIZvKUfubAsevr65lXWGsKjso5raNqOlcH0OMAkx39eYyyEqfJIuv1cjHCDwSu
3AllT0Lkk+9blyjIOoAZk2ESx8gA/XyoIBGjR9bOLHynW8ekTeFWI4ktSJAwTyll45kotRuswR+r
vJWON0FSgoA78jmXRdhiZflHyrFMDm2NV9kQbg0LRiKiw6qP53JG6unetnE5Hlol/V9GdmPyxhgy
6qOc6DUgkV81oB27DNkRNtQIfG0JxfkUqUF89P0ynaYUrpCqSNBh1hqvVin9Lk0glTGpjY4CtfwH
8oDNHlrhY8nYURIdgY8gWwnyRC6p7/oTWdTxK3IlvyNjpv8zy4vv73SpXLh+GuQHlWQ4GB6lYgAU
U17XvIzflMEvWeZSOY4ZlcK61Y13gFfWjhTt7vJqrgdkLtxrWMU/esZO4p20obL8caIUkpp670z7
dWMoExM1ZIB6kENbzqeT1KEnY7pqu8uzyj10RSSk/0A73Ddwok9Nm7Br9bfE4edlySeFTK3tG/I6
hVCyxoCBDcRnKxNC28unErK/ykpi0uy2JOwJeNCH0Y8CGO4zfoO4CNX7bz7g5oUuD+yi8aHVomO/
Z5bRQVj5tj4Fv2wt8b5rbpqEIboe+dzdugEdYQCfQkxeOA8fd1cYNS1jIBr+659Z/BQIwsFUg2WU
yoml8Y7eW+7x6Jlj5UQ71z9Af56mu5nNOqzbg4SXjBMZ3feqjS2yrOyi4QSsaeE2Q6x9n0gHPIgM
Qe5+kPK6QX6dHZN5Xj/mkBWnI1aVfgcS4Vu3RLDhn0GGp8XdOD4poxaSCup/vwxkAYfUbpvI92IG
Y9kXy0PrRxHIzAucLAXqETbsJ4V5MThpV+nKxc/Xqjw6oocJkyk/4XAw2IalARwRM+iAulJU2bia
JmtgAw53L7bxiRULfWIqab8r2Acldxz81fDjJiYMX1PBk8Zm4tDu88uHSf2AbDqtppgOFVUfYvzZ
tNpyA7N+nF6Gh5c4/obspGCtYYPncYnpXooXCCdNBYg/QXEnHtQMh8Nqpq4lMvl7+II6cpNrwurc
xazI7U3a0fBbRMF09ZBO69CfFRKG0gT4pz088jB61UX/3cMf7THYZZfCCvu3hve0mOHzu5h9Bm8V
Ryl6oEiqvUM9GaAgKxA88ONPQW2K4mS/nemuZjLTHWeXXUPckluD92i9Ksg5O7KOjby3mdQNMnQq
2Av6B+UL0L8QF2gLEa0NcVS9pVx2fhCw2DKtsOh3fVbkO5S9mugMisrzLJPiPEeHYwSKVeZmueKq
y5remPppqYi/CXgBq4bSvCwOdgl7U8e/CeYmT5gt86izJVdzC7Dtxptg9iq6V3QaDTiLWMrpBFjT
7MhblLoexmG1Vuj54Vm6aIWWlJPpCYJbFsOK0Tu5q/lWNDSRkJNDmuHx1xJtEYhvCv0dP/7MhgIl
5Sbv8OVM8u2a7vB6sbPF8T96m06HctPfMaQFnKzR9QBsYZGR5/2IdoKdgWC6hAzkgVqpB+tEdQAA
8hbI16GVnWmE0QvLKCJEM4LvGDB7Q0zP05jx5xFVDgGP7JYy1ZNoVYcfmSibfaosIyUGcEVZGyov
sZDTOIeyQ6IYF411IkZHXieGbOk/6WFSIy5GWycKTDvi17N5yyBlRLC209it0ynSGUEt6UwQcLtI
WFaVIZmf3m+EzklaQwUCRLuc5j8dk9LByUv8SQs6DhnUDotgxVBbqI2SixBVvmkn0siPLTHcU90w
Mc5prHOusWe9ZKr23urdbbrUwkudArhdiVsoVPRkl8m1wUfMFha6MJvE+cJ2qssoFnpp9xPgJbXc
py7qaFJ0wykJZyK6++R2tSKEpjSxIklCaty/4pcVtJEQlGQ+Mm1SRntsb+PAj4Y79tZbp323o/Q0
NjRRJ6opVxfTQL1Aqb0lyy0AZX6AKt9YEpyKT2+MtMoq5GR0nQ7oyoDGhPItcHhmAnTWek/3d8c9
QasJnyGfzDenWLx68Ui6wgRNCF5q22dgUxVz5nvpmVb0vuFycowMS7EUNMbH7o/MQ9I5PYeArQLr
+VavzcyvXq5ZKW+jXBMonJi2uPXcBViOkyiptiYrq3CGgDkDWDTGCEEAyibPfvQtKS2gs0rH9cuh
+TdKkf/Ki25ytn48lwR9N0VZUqNPY+DAd9VAr6vuxqPix5ZbFs4LAKYTmq0vOcYH9dAIr7t12mw0
Qo0AJVr82HbaFBl6eiH0r4L+tVJ+J1DmjjpcWeu7oxF2Nisf5ic4bqrfdTbHWXLBWR1XvJYp5Z7/
J3ZIkklJFQmzz1mK4y1jueK7xmUYYf4aD+I9rwsglfxXQDfNLOyWvlA6vbt5XGkvu/IGHS3KLAjG
aeVo8pJy3DUioBnEZzTo/WiPD86WG2OmAOitqhuFkTJRd1qRl9ekweJwb7ZE453FvGFZ+ivuWmu3
zuBCb5MV6V4APa7y4k4ntmkWNpfbjKo26+/9M2g4C+gQ91ySoJR6XroMacVwhg/w0131juzbBrQh
nitd8vhGsDklGp7IrBRD/4E8/EGSol02ngXh3/DtYBtelZnobtbxTIoe1x3TY/voGllRebNfpEgB
Cm91N4M3cyYN220uoAyO6SXfbyGa0y6sRNAjAIoEb1/LNW1r+gt952C3yH08tuweFkk3nmXE43Rc
kN29hNEGwOxrRuu17ZxtTA+YGQriEE0xlHK+b5jO7kx1KB9J8ZDJ6ri8tJ8KQnWuSOx29SlcboJo
zycK8NdL4IBL8Eyoh7NnNqbwRGYbQqZjJMZmYp4kjKFAjlyXVbXbRRrxkBo5GCnKKrO4eisci5Pu
qOj4MLz2UL3x9+CzNXaRozYvBcOuN/BZAmvXkz5ysiYAPaIPsnbphmqSwZ8Az+Ys6WV5GoxHjyzx
zB0kHkIT7TlkDtHb6BBk+3WUdf0U5epKKvQSRPpE5s+LVEm+iycHl2XVvC3M4cVedUCizHGBk/jf
WoSCpRZiUcncjGM4CPGT/MLx6Kx5owDM4kJ+ALdErpX1EOYp7R2RGQ7hmCV759/8CZnODHnV6Uou
VX7FbzJ9RF64mm8NLsrzPtZ5iumscVgm6XeQSl/U3WtD+1FtBzWwVirhNJZ2kPTZ69D5LCznk6PD
PPqmiDEii7WlJ4OaWYVZN3ADtswZBlAnSfvSfHZD5xBL7IZ9qZa6/4uQWY6Ea67ZD7Rwk09JrgL8
Ay+aIrUeSd8KJdP2bOlKQAvneh69bu1ApCiQLfL74XFZ6BxqlRwZCkLwuWra+PrtuTCUdl9L6DU/
VAEwmGQDXyCXhXS6SyBuA0PuWZuLCeAgwZy7ForxKlaP6yrQEkUu1V+JUsxJfBTxz65H3WbnU0VO
DQ/MDb8yvTHO7s78pM2PHdTLleDC015kRhTPkAEK7pVcusrTk228L+qLwpkWnaYABX53axjL36pM
PSAjFImgKQjXR1OBeq+mDJiCfLtRo1bktE3tvQyMEMbpg0v6CUhmkjTyWvdbT/+U+9WWzQPwyY9H
TyjyGkrHnOVN4JLh0i6LFrUs4vdbDQJXt5ijI2bUT9HXGHLSAopjexdImx/d1sA+qKL8Asmnw6J5
XoYx+2CP7bgTcPAS2+hfaY53zdkFA6QpUphkcikLzYRvHGp03m1+5GYkFipGAJHFP36Hd6oOv+mH
EMTD9ZlDhlGS9iq6YHw3dG/9mcjJIPHG0g1ElEUdDDYECyQyqy2fmqE3szqfdgS93oSzjYjnliGN
ul1KlypRufsV/uGcGNcFM6WSoBEIhgClT2uOoWa/OSp2uwoqOW/glKjGRv0jrh40fAIPEmRcVx5M
Mz+h70AxHuscSnzdWNV0k0cJF6rUyYjQrlcPaYmJM8LdrvDHOhZmMil8ZxYKPJAZuOD5+9gtsZyw
lIuz6jd8ruxAEdd0cbAKGdDUZ7rVPyMBa29RJcpndf7DM9osuban+D9c979NYZDlk1s8Yg6vZDdY
3NR16+zxYmPZtoVyqX5rpbrjdNKGxTS9TiyXD6y3PdAdRAJikYG4PMCm8gbmpwAJQidMJ2fYg19E
yGMgRxhay48yIBmAZYVh8/Uniqor6ZWYXv0bufW4in3EAIQs98VJovicZFN+bxYB5wcXW2V6eDZn
rXd1tjkmWS4RlBVPOQyerkhwI+a4uLODvcycE5ls4WAhgWD1s47sE/LywYztBRTFf8YRUSvHwEdI
oFQv94gkjhdBRY8FMZ+VKudlZA5dzE5n0MNxuuusrAy7z3d96RiAFd1L8ZQFyl7rYBauf8mwDTw7
fXY2NV0G1MOAozTqrGXQ4n5JPU51/LzJSt9S2lS02TzdfESViUyoN90Di0IeeEWPpz7qgORcrZv5
bzk7SN8YEcBbGoJpnfWnTvqlV1APuUaSWnC8W6ywmNjbOiaQuG0+vURzFRhsJNxFVHmeszABnkvy
b7YhscvjaG4gLdhLW1LJc/5rJfQu4RikRRRyS1FJuHPiidDhY4adkjoUbPI8GWiwyQleoNoYmnUG
Q+e5rn22IdMygl1IkkFr3iSW3+JXdvqjzEAEh7yxUQc/3O4WqWIjovccguxchNge4uLsZcmMofq0
sS0JZFOPYDhp4eQ9G2f1iShLtlR1SAGqeUw0LmlM7odF4Ze1gCDqrynZjq+Auqq8GStqjI28YMlj
4R2pYwEpxxET2Kl/rSzVg3QUfywOJkie1Btm6gZJDqaAV5o/lL91sMF4Dl6YuSApz6lx8ZNtMj4L
HmW4rPbSphibPlYb6cQWZaK1RaGTOcYSdKbBRKiph9F4NBA9GQNYnFB9nJm5kVMHH4+ykAXIJR/z
XFFpp1EPCMiAvbH34Jl3Ka2TAtVqDFg0dpTzxAqVmDlCdzijf5CsmagLHi0jk7lNBzujV459RCsz
WbriVVGSjv46q3sbsnIFsA7f51mdnHsFcJtLsFhhNvL1FWAtilos0jOerHVOoMNBxWv80IgQxJcy
k6igr58EP8jpGNJs6fsRn22XRLxolhia3HsPcYX61lea9CrM+2+uDfcD8zNylAfyJ2bfT+v0d58p
G8sBiXWr5PoMXiKE/qA2INPhx3whPvpn1AbRqsSd8MN0wAoAtrMRGKU9Lpmo//yzucbL62Z/M+TP
fhQ134EfsIBr5NoqXvSh213wBzqGo3K6A/RR11n/yu6t+HF51WnjxtP+WMAWDbNm3ftkUqQ9s6bk
ofEO80Q5WPtBh83UwH1HUZLFMMlRipJ31NqH2uL8/DUfez4rAI+g7LmfXOQCGViMd+HwPJG4zsXw
6oOOQObDW+8LqxPLztugjo+ziSSTA6J2gwriOcRoml2AFYjODQHN2QUHs3hNf5fmUHjGWjxpP+dy
GQ1n43PPoBHK2PLRuw2WrMj6+Y0/KEdQYAzRoFvUQdnRu/IhnDwpMIOueWOBrzpIyEbTYLLjXCWv
X2Z9s1PYFNnYL7bdNSuLWcfIErayLfzNjyBpawkxfMKbjyyPGlEawU979w1fIo4vjMN3+YZ1cVUL
UxBSUlv6OxVHpgVS5zKG8GkjQpyHeNtEchfRz7hH06rMOUwyYMkBnzj8X7bq4FJmbLj9fgKTYyf9
SdWystAZ//w9JD0YA4mIhq+0YNSsMijc8ASAwDwoEyONUHom9Qu7UW4RtzstHMQIMBEEDBnAVQSW
DjvqjSfnhc3w5NYmTUPfomwq9smC4p3Fw7FruGnfndgThj7MRJDgIOlcnYjWh3lhFMv4wH8kvRMA
l3JiiKFKzUdKBOCySrnVB9uq0DmUirrTX/NMB3m8ccdWCMWN/Iy+d3FEzLpBKH4Eb+rx3oQ1YbV2
mEzSBdtqtTcaySzmwDpPyofN84wkhc2CXwUpS4miy1q6kr/6hkIGnFW4gnLE9XBgAFhFVQy2ns2Y
/He9uKsfsP3dskBvyk1jWDdvMz1p4Vsa1fxfIT0O+C7HVD8FQG0aibZkxM1U9pQZilc2Z/mNRIhw
NgydcTURUipl307tBg1DLki77moaPnzvOSoPX6qA0A0itJD233ZCEkNNVsbcccOUE894DL9/gSXG
gmPprO/nrRguDJNQ2yHCabch+NgPhnREEd0DSG42XEPon5bJZEr/1kR6wFctqCvpUrZWGd7B8G2L
w3M4SvgCAi/8kQeY88uoX/wxz+vZYxow2vlnYguz5x+i3S1JRaXY0wGtUCE9pLaKGHS6k0dS6w/2
EjV+eJDKCL69adDdL7diIlP1hyfPjpvCApp9hOUSnQSucpRQpOlcnB+S4oQRWE2Fm5ZnFMAYR5K/
/RbSi7PmPCeavCttWPJWlwh6KNRIEn/LE4LGr5BkDnp9wjV0WZBvJzETtw3SBv+BqhINmJTYvdzS
qRoixbr8zC2fC3XKc3MlcdfwpkRVy4tJCWHpjEht4hb8s3Dslebv36nMkkhyxW+EnALH/AmTSMQE
NvxWB96XVTk3hp4wbIvADqF4IHYLefP056d0dMvG2+sB1hdk9GwkiHMBJ7f8iFpP1FKexuCZmVVL
FZ8pZ5k8sWDsWcTAdTwRqW6z5vMkebSeFBnlCliF3QKhTD2uzl7RdO3k9WJMsvEwmlNzv2aTLrm8
UKJ44WtLeNitSMqH70gspMWqaA93Q6ItW3DKZUZ+Npswyt/W18nE4dpzh/knF+IHyf49tw5YEh3k
YZygvFsOxgg274k68QKC/U9gvq0s298+9ak8VFuMGiK4wy6lwCbxgV5u+XMmmXPRgIjAGOx/+kgH
1pvpdszTrvj0DnjWP3Rx32yVPyh7Gr1WSLqztYn7+CdjPB5gVmH2NtqosoqcogsigVhxDSD20jwL
eZj5RYzxa9CaSt87aRPgz0/upqcM5JZLvGIf5LZGK1YbZqTl/NWz1EoGGnnLJRCGhJujfAjWJEWG
N5zPhNQdDCSWaa44ky5nCBHZorYx8ecAO88rxs31cuzqwHbFn83VTYM7vwZg+VBqj3PuA2y2cpg3
GdqfMHM75glrr4wrhZoT3fnzHpf34M6cYcmZ0YR+WIYQgtHiRe9livqPWhtBpzMnvUSQb/kVCYxK
qAhP75vCkOsNgXe6ZQB7yA7CkQeZUVauWwp6qFJ59bRLDRdRru3LW+9PK/4qX+59u56b4+jS+LRV
jlSSHaKaLM3g6wPUH97ArHn/+ZXbc0m+37/tAeD0lXyar8ZlVGgXmxAiueI4Hjq+22jXneCI2eqo
qBCiQNET9zxUlvw/QkxOLzTco4qjgV/bacmlNR7O+5bqC6sj7gWZVEK9uVeq028vqTK1Qk2lJEOI
8IxCzp6Oflj1OZ27QqwEuVl7vZuZPCFxwD0Ov19QTLKBoz/jKF0Ab2JHfdOkFRP5Pe0/EonduQ8u
JMBciWwgrj6COj8rW1nTTAxixMfPrrIDv9CxSM4P9iR/Zcdpw5OdSSphniVLQVs8StIbVhTWn/A5
vvdK07fcaiIfRfT4DvONFS8dzKY0RVNq0mwU0iYRIwvwLaIsfNkWyjC2gdPXXlp+nz7+sdeXtQJq
bIDDlWKimVi5guqYG/4u2QMS8jNVm1sDWLinQxYC2K0u3piJLcHcJWkLR5z3BgF1ldO4BfCCsp9Q
jdIM/TGLridiAgajKNK0pxxWvf9BeyzxwROnJsNqIE8m/eZaVYYZSUiyX+VzZIeoMVvdu9EsHFpt
nElteslaCgKDDDJa/8vLVRHqUvWkgXib+8tEECPO2ixMgYeUh/LP8ST9Ihu6vM0+e3+GLTUOp2EN
HETi0/Cz+ykuKKHvQG3uhGJ6Qmyi7bOGJ0xTFHVoXDWXh3g1Ig9Z/xBFH6UnIKkB06b8PujJ9EyJ
0slsLP/as+DuNELXu3FNtiWPWGJI4dbAggQU7xX4HjcVA5kHfD4lHAOsphpoprcICGAF0K75z7Y0
trnBXhqrKf9M/+N3SWIHDSbx8c0EShRvDDmRtMbzl2scmdP8fURdbKSZA7fLhRBqo2GCmUFsb3Z4
AM+nj/fA4wr9pr5gY+tZi0mfCG6UEFdhaL3k55RtxjEkTvDK3SeYyk+/m8xGivxDwEejRju2WLEj
vDQXM4fktNTq2MPv0qFB15Xlt5SKVfSoO3r6UMAMpJowwNccK5XHRlLMK1EK6XbQDSZpenKI9Y4u
MHGvy1DPK0CWVozcExqK9RXOAgWyvqmZEpBJfl1yZnA7OAzdfRHvi3fL9kKhTio90iEguh42LZmp
fTbeunW+sZLb0+OisPUdzGwMUJqEIgIqQbKLygRC5h9yCZMQnRHcmvipS1FcEmInSdMj83+ebU/p
hb38lpPZuLZMGjeABRPMFq79cDTmPV6/5Si8DIQgwTljP1y+i78uvnW9demeP7sUmxre2YsdKWZt
usdwHDrutXoGxHGgq5hKlwgvA0efc4tM7qrDNP3RQ6zX3HPmQBe4+nzdkLW7427aDz5C0F/WreZL
9kTk2Q0diMP5zratHbKmyfaYXWTtIyoassCsGAMBEpX/KXTcvBn+30DdCI39zvMoCVU/3NGcWCJw
epXaY67MrEA2YvZrLMG2IBo01CJo1fpdzEfVHPgMs9uObyBmjVUs3ZDFSBCZt0Hh5tPRA6hu7Xnv
74gjHdkyqo9h88xbO/G8mbQ4gZzHlZYQo47uer1b4Yn14zuP62QJfouxz4IC1pNZlzb3kvz9fhaa
GzkpRmlcHuWI5NLQWkvIvQifoNfZF/JcKjFK3hXyVGiOIe3UxyPchhdPLz8+nLSvCEHUGnC07Hr1
kiORfIuP0Lxw9XD+A9gy3Tj6EBINaWXArruHNehrlTiJb5aT8SUiENKy8ip9DKRn5wNonOSo0PEZ
W56qcBRZCKKDQ+rioq77PW03YIkOUCNa7iyvru4QlJFlEm98lbU4AnUnyoI7/4lEma/Epy5pKStL
l6Mp5UYUG+AXCufkhq/NTxcVll004VhbdIP9XkRouBlPFNp/L/4kQuqrnSWITTqIaAnFMMiA8Ws/
Xm8uWjVdcyG1m+HfoMUgMIS4cNEjcCBYoh5TyoSUOhzYPq6Zh0CFRxDUCLuEG8UVmjw1vELSb9/x
dSLphjTn15r+RRw/hFP5Thua1C3qGfTcjVxJxPBdddZ+nyZjd4Yf8eFA7n9rb1r4c3dXnf9QfmXb
HhcbiPTldU7Cw1Wzv70jQasXO5wk3E6UF9+xdYm5xAQSI5MYUGIlb8NozUBOJqCF7WGke2/UPCxg
CW8zgfar8B+XrbPt+CxNMZ7CBx2gKm7WIIwm6dDPlL6bokHcCpTU592mbp/s4Tsa2HGrfVolhy1u
K78zybxNuBevgZ7Bn1BRoJSeKXq9nUcc3xPDDHe9aNXfXpBDbMYoKpe5QUQOHjS+qZUjTPhkHJHC
JAMxOJ/Uv0fyapKil6EshTkyZt5ne7yu90YcjJfAXA1m7Z5ElzRQtOrLXnCFSDFo+fbfYkTYS7Vi
JWcmMddp1DktHkhX+eaMtwarnz+4zPvs2t6vie4RIbBNCgBsehatpzBVBgroCN8yYLpFuqo46ju5
iarTEk4jZFw3WOTqyHnZy9QAKBf1YB/5M+Jgkhv2Lp2GQKFrKx6/WqyAGZJHwUTEKBGUjV4StbHE
RRuSsYq2G3/HZMgkWurREiSW9NZzFYh5Qn/FMFWWsyWZz/QlH82+GLxPZftogZyVpSKvXGUQBGEo
3n0xnGCr9Skwl1k2PyADa+rdLR13EWNIdCnXLZCqYMb2TgfsFEldXjvPpPBOj0iFyWsAXKBd6pPN
BU+fsNjg/xidiCl3OemMitZMqUiOZ7cZaj/G+dZ2JkJKgy9IGxV2KIZZEw66Nsa1X84AHQDMll9a
pMFsaEBQ5637JRnWSsN3a3qK8hHCUNAS03EVPiesJk6ZU1mAAsxbsba7O0pRqDziS0T+tZs58nKs
HwQE1QqQKlcGsrTBUcz/9LrQIm5XyCyBnZh9GT/rKum2rWlkwixCGsX2lOoV8ph+MY7GtLWtB7WE
j26U42E1cXIHPUWZmvYZrXu4gKYNFY6zUXZm7dAyCKsxs3WQo8LR0QUl5t9Imcb6b0EyVHqwhNQI
HQNcHQLzOjsMfrPG1GWc/L/PTgUGS8EFTfpTBK1ekMhFx08KcjjbLJO2j4ncwTDgBMh/u9Mhk2G/
W9Wll2VGS4ch6OEw2oACVO0IJm4NurrsbJcGfdk5CA5OH9Y3jgkBH/TMODoo1WnvG7Ye+IgpAT87
Hqo1ynaRHt8sx2uAaRRex5yrlhDDV9OaxrI2jjKUtU6nNXEdnN6ZPYIJfo30PD542trY2eSL9snZ
nlbAdCoy3khWw/9yofjNQ/EkZzf81FzV9i6kvQ0uhtjAw1/XSIFPlDNnu3G7bpO/E62SyPpi/unZ
ld/MOPp5jPygW/0TRZhfCDitXbxIhgR0b6FsnLSGBhMU+SzHxcvJH6R42u0QCWosvtl+Sbsnfr6P
m7f6yUHVJn3dyjJIstOB77qZ6W2iBwYgweWS2l4degrz7FySrQB0SBkb4pWXDovtV1Sz4dqECnCD
qp4RLmETi5m5nLAR7ofKixZW4pxkBcRnue0Ez7Yw3fHpSIbvHw+pfhgRaD/XTpRDix8UKa2ECmYg
QKa/xd4p6vT28z0Pcld0tHXrvuooTcxPgpxx+NXqV3cru+TnT9d6GxnTNYjZxBgtUBDXA/fgjktw
MRR/trh50jisNROweRAjKmcfOAbXcd01JQpdLGTRv1rlrrM2stmE87Qpth4UHo3dyO1/7aJa6hTk
EVHKYQI44N22w0S23Wj00BW6y/w9Jcnd8lijEhJgyp1hFjjD2vM4NAmoO8l4t4ywObrpOFQDldu+
TGz20jMvHvY+WPBqnomSWoQ9oJeec6vw/IBMYzDZz2IftQu3NiDT5U9lLjSKp/xZz7+OE56z7W1R
MUMxf05ROhB51jXxVLMLmwLBvl3gxpVs3I3egZ3I64U5afNG5KLjIIrECl8xNaND7VYADJQkjJ1S
O33m6tzwXRVFvcX6HsajHqJNPOiz0BTpKFnFQ+wsnYA3zz9PAhuU480DKSDZSwNwvUfvh3Si2sB5
x3VP8j6ytlfi94gmk7dkiH7hxqI2fXcAvrgcJy8mOohrT1S8BxtpHqnbnASFI9VpOz5lu6qrXXVM
9lL/7xf/BzT8wQSYGktT73phVTOPwY2pV9Qfk32K/TIaLfTxRIx1i3gQ5ZSsCMLBQoru/TXhVK0C
S8yJ6BsZ+osx6o9K6w7Pwc17mAnmz+0cfRnXCWTvPATStp/0Popq8IDyTuCbYM/mZf5rqzP/OcqX
Wg29870+UgYlT4bbUtTSClh8Pt9+EJW2I70iCqI6cNELj2ZTqgBMFwk73UOEpo6VLnN+mJTF3R8D
+1RTV4YZnATUXocksyMajv+3qvqT0NbOKsHlDXBGYFGTVo/qC+0wjqtQFvX7u+4vWDAt9XhP2NSG
lG2uOZKXx3/9LIoUkjNroEAwpO1CgSQGQijW3kGzNTV4tIG86BN6uBKZE+PqKWYt8wxD0Cnvv7Fb
0eWZ1WNy8458iqMKf0bLF23V5s3eTfCV1ejGafYGGdiG8e7THe7hAIeo9jfe/h3NITGZntgPZ3dN
4NkQPsCCbCfPn2yFeQc3gD92TdFe7d0RCl0jkFAR38yMaGL7ZxqMP7fOWRWmHQobGC3cwr/QGyfI
yltGIJCZ8lpd2YMbpUkYaUBN8KTBxYpAqiPiCe+A9Re+WKvNpI4ACC5ZKbgNbmyCdrMdwxrA+ffJ
dc59Ff7SHGlKsnzNRPlYy6e9YUDPLKahHCRgn6ng42St0U9ds4Gr/6NZ7lQSk0GhCio7WDsEVghX
ExEMUvvHxL8gtqJwGMHrX+Wp3LTrAxcWazu2mTTY+ZYA0J6wE5v2XZsgAwfbBnBbVN8WxfjOfXFF
olP1FhLXXaG1Jn1u0LsOCJUQ1jV/U0wFjQFAipU8oBH8fdgSSV2ckUTw8j9uImqYNBa89C8kvaE4
zAs6vlsqhc3FL1XPSUb8brPuwkMfPruLgsvk7TieZFcgHx5S56OMYV04tP6NpfO1WBmtXMAmZ0ZT
+lzZeY9oUCb2snaIijOppX+CjYH+756vL6JCMrvVLfEabGutWNVe+5Yo54ZZqJTp8fDhCEU5ob6k
Vqar180FNHVMkCfvbNCAsYDJAm9AIXfmTt3wCuYxZf5LNx/10BUkKPz0Mjh7rLhUIUhQK+19GB9X
VB+tfSkwli3BoCMZI3+KOx+YpHsmXki1JWe3tgBPRFYXZzFpz2tBmRJX/Qk12pPSR/FXAKHyqlkO
k+OTTaCcULOyWF6fJwDCRfGa4B6MGnBU+yC+TAA5Ixt40IMxNN0+mDiJXv1kGnU9hoYaAd0AUJSX
ZdcMH+48ETyGM7VHgytAwrmO9GtPiiLvkvYKpbkGdkmjg119OD5L/F6tElJv/FFn0w6F/sC4Hko3
ZbpRVaz/nFpQygGJEZW3aD4XJU2OKkld1znfCpjBfj7s/oHIbGrlIUy6XQ7K/JjHu/blSZA801NS
JMb04WwgDQN+hK5PXNczNrqOZVakVW/z4wOjZTjvwgMKGKjRBGqPDjId9PnnxeHCzhFOoTtUMuoK
b+YFUmYQyq6kTq93F78Vh5d/7P+vtaNIYACdcu4XmamZymUX6liGbaZvMifvmi5P5L3dclPYCX+C
hXlbPEr5ep3q0itFyPVdQueDkEMZVGcP8UIQeDiNiOn0k8ownOk//LNYzEo0v8sMyzi+N2YYsXG6
aWp89NzJkyHUCr+jx9r6dYJdAOc5rzVW9hpk5aMgZAEPayNXUvp5vwrU/3M5vuOS0nD+adN234jF
YzrpkgytqYcgGsCKiqnpOHx3OGBrlddWprsmQJr+nvlD9JrmQiPNcjCBoH/LxTr4eqPCgl+XVJ98
zBErd070iokEvCw/lqBI0pKwA0uuImbdFA0LvOOmuXFsBBfsurdOn/ADA0dfHJr69ItdsvDDmFdg
HV0qSxH6CJeZRpbEm74ctNiCZZdluTkAUXlMFL6vJnXwAE2dBO7iaFyGu53FHDQAr3ANz6vzly8P
2cxLyRYgXkx8FPu6+duLpYytAw4Y3e3f24bCiz0WMVCEuQVoxzEGs2J5JgxU+AYzlrVj61aPyUzm
6Ciki7rjILIftUUiUr7tHoL6k2gvDP/0WhZN6kARHxu9ZXZfq2wf/DmXglcqSmftQYr/wfOtu5Ua
wbdpGtPwZzEF3LlM+1hX2Vf8OGkdFyC48amDSEIiivA26JaMnRSgDBi/4ySmt2mgz+1FfcOaYpdb
nGvku9noJYxaNUhxRTzI0TAfXqTle6EPY/WpfQ4C33xKp6kFjAblvLWpjFboZ6ixv/uEi6OfmSwD
a84/o2zGV3E4YeIbvqe3zZXM7niZ9ehIcKslmIBA/N8mirNRagkKZ3BT15qCpI2JZIlg+RigO0tO
p5qthnkDBpgiUzh6RczovJZtmVrj38T548QLYzjOT72mNvysVAkgkISMuxzgXuEvhhapyvA6g8Wo
l3U5smsYEzlej6Z438BsCbhqygOp9aHWUf7A6c9SUi0aGYuOqGtgfNIZsV/+jgD0hbyvpHgTc2uo
itDk7hgG1GMU1NlzfXNzIdZgL4A1VjGdRVlijFbHavfWCLCqVKoeHlD/Tm5Wwp4L4sibUGDiNUhJ
V7IqQimuilVyeWUFRApqtbuK2mAJFo1XLmrIIR/SbPjC2fVo+hunIRiC+e0s62pph8+a7jUaSIAk
mLsBp/sVIVvLnZQQGw4p8BuFjwuWnu2rTMEreQgXMXbgdW1O53W4SkMmshCE/u2FuvFZUZ1yY35R
j2IUy3dIwRHZCsZ0l+g9hdQNbwG/peWyUAfruPYGU+M7H/bfCgrIipX4uKJvOuw8sHyPFvk5flQH
uEeBtMDS3cHUCvK+VgXDYKCrDKbPDA5pmyiqVwaQfMu33LZjbu4FVwW36+6fNhHv9noujT3nhw15
cjYD4RNb0lKZ2mk8Lm0gbyVGN1QUoRCqqQZQtotRnnaoERp+btkN8Pim9nsilE1edwexs6GigDci
M+1KQHmU6cqVErt2zcinChSKEvmSOutA5aegfxq2KtlH2O2+pn5EqOKlQw3S8YkBi0vYAAseG1G4
xHf0WFNPeED/dlQSaVQMzS6pJKA1eor55ME7ZXUgCr+jK57aqYyAzb+m2FrS/twWD8cHwKP9Yfm4
mDbaOLwleSXQ2SM93OXcdGIyZ+/prKsEDRYnfPB0cK9Dc0cinBwkbiYyiuReSQ9H8fcfWR6e++Rz
xGJyqYraPY4aFitRNTCAWq2KcRVv18Af73j0y/dh5lx1xBPSkG+SSeHDhoHA+sYwZCUVVEWLF9N9
WHDb6t1SSOcJiw2XQkTKykA6ore/7ocbstGpC4D+j+9frd3sJfNoRCWkK9O98vLle8YHvx5P88aq
u9GBAjTFxx6t4AyLwMjC8IXfXxlLWH7sl4J8qWOGKEI/WnVFkjdjk0HgRUBHVLxtYxMcjJLY8Uw6
P6GhmY4hjNuPLrIyA+gkeK8XkPat8gbpIR4Kh6CPGRwuv/OCV46lF1FhzgRI77oB/gEZxO4iCxCG
d1qOmGhMdU35u/IUgT4pyzLfhu638yfA1IjN+JEs8HbVvrFdlZ2XpHCInfuu7I56lIJFn+3shEgi
9OebkduOZA5FYE2SiVXAzBmgNOolkJ/8RpPqdkpbXM/gWpF9Omb9/0HrkIeybCKq4tx57iGDq61R
A594j6C6dcwoaokwmLsJgZLV1TlzZh5M4z3M1tl53HNl4GtlZtPgVwv0kUYd729NzAu0dTvLKWra
PDEZh40TLlBzNOJkXMj8n14PBJW2W3iPo+ArTAj5iAEVVIBqljTwZQvne8AwqojMz5kp5oDWp8SA
2l98zXv0kClNhet2z9iWYU31EJU+9TWUEYfmldIR44Bnl6InUbqLSswefdhe3o9s+sisGUr4Rf1q
E/sMMd0gFTIBjFyq1aay5L8uKnhi2vDrf7bR85HwnppTRP7H3xScdqWpAWBpUfdE4DiYGf+g6OyH
yddWFqorR6rATmNG2OwBK/k0ifVAhgWw9D68NClNEuo0Lf6Ri7Zq7QEeRaefb1jlvPT177YtAkPl
V3TSHtSAuKEdyqY91EwcH/3iTqyElziuDOQmBxnAylbxZYs95+gEoKFZbERg/iFOS4vzY4GHvfGw
5DkCslJ2G/U671Nen7QHt+AdS1sFaCAnaS1gMgGPxuqghx64sNS8F8++FIt4OW7GhMh3duBo8669
hH2o4l4nCLMUuwplUzP62MpMT7FLk1o/OJu+MkWYVTuRcfidpOF/SMwMjEX5fCAqA1B1yOo9hR5g
jRKEvLPyoyd4udIP3S6EXW4EfYxK5QAZShtNJ+grLDZtlppyhxCxpdjZydUSjEBxy7/k2xII091t
y+ulEJUoonfeRrwSiBTQPjw3iPikHuVeqoyLIsUsUEM2u9PSlEjr1K+gyCuANhd9Mw0nfpwwRAH8
X0Flv+8QpvbDYxeElZAiEENygwSQeb7c3fe9sjj/acQ38odUFRqKgYCCoVwGEtNaAxj7cl9JrNhW
6TwPKkBqF2RF8JL6Go2EZlP7k/f7qWprQQFHhKrYAWAcogn9SAuK7y5yBj3jdvdHRbhDeToVVsNI
MN+jGX6kiHhwnmWxc3bFtuz6l/AzrDbkm7bJH2DC23aGfDVz3dt7wZEbWDClEL8GhPkUF21TID31
RSzuYjSYFUPyByGrsJaHPZIeYG3XTdrRSmW9gWM8h8OCoK2Zjw0VMXxDUWaTU0q1XDCAeOHz4A0w
dupLw2c99GmysDfIVSOEOofruT5vzzhnVfRH/am7vaEn9oFGwZoGvU0CiTUjSiyXdDr0ZlDiQ3az
8aQv+UcsG5F1tVpQfUVEJD8zy0jt1/AmcY4NT6KFVn1Ia0q4CwzU++uc8n8IPANAthcu6AehxRKu
PMM21tlUMQ2P6tY0pDkgaJbtroOohr8uG8xoIVOB+ocMfQ3h+5RmvJ2ZOAbEF5MpqB6xwlfUvduW
jWKv3/aOe9CIeFP1EOrUAw7zYcdqkRzJTLOdP6po+fgWejnX3H04/svI73ckVcu1fCe0iVbhje9R
47Qv3OcoEj6X+aZRoJ9NqZNjQoNCAGVJyaWq8/HJ9hh884XWt599OWzdrIB6k5EnQ08mhXq5hhDD
JL7r0aLi2ko8lX9ztdp/9QQdID+lAd49rqRsD3O+hosSM9O/v5gNX89rfcrIViUYEH63hb/aBMQ8
cwoKiPuA19zg5nIPE7lKKi6qjfaFu2xD3EtrZaa5dWOwW5eXXJHCc8eBLMw2p5rc3acj1XSaIjyP
+H4YVZbvH8P86tiko1CoSMNvzXP7+PtIcsS4uK/rZxFq8PIM11V4r9F7GbKkkzjpGzQufllO1PZV
vAYbaZdW0eBRJeRPdlgHCiZ3po6YvvaeUDSXCFvMyydMmPwRpP/0NMuD3AoViHI2OJ7ZILkU8BOb
sv0FoVH9iBYs0fKmfiHJN43E0B+Sz2QITCHDH5b/lniwkGRPkZu2UiTTH3eLoRa1bzdSMm6WjSvY
JVsghL0k1+LlJM/I7/CD8ItU9O1aVCQbvnHJzC36ZHk9CtODxxn3Bx12eFe84Cl/lec+g1ucPa+y
BAXNvTj51Ew/aLeakA5aaUZgj3QFq8yUv37OXDTgKJkKoPLbz+loKLOSGXUFMQW+x/jpwiaL0zrK
PoLRL9KQRsIS2maziGboEc1fK7em8+nQArkZ3+CIoXt3lHnFnLtrd/hYXGOUCLDiIgNM6K48dFSb
/HtieqAUoDBOryldRe0j93vPp1tQc8pCK/YzXnmYcN6ETXHwhmUV4NsgwC5svvzuou+USKt435ud
lXFVbbzGUGiStShjeP92fOsZOx03mrObLXYqPf8j11HnFZ9JaIu2ec0rZeR9SsgNRX0kgoO4Qcrw
5NlUO0t8SDEpW0w0VkGf5yfZEPA6lRaK0gmqjWjr0CZB6JGExv6gjE3dZD9XTek3YRJcdPenZUDu
dqEPe7Y5iZqEv4UGLkEmCNSBW40DPHFQ7EO5PE1og4o8Irzk9RynqOtb16uvA/B+D7tnOGSMkdfh
trRtwXB7Qup1XcoxLdVPkXx1f6VIIrMuNvifBGrfnARwRQPJ0fxNV44nJqefbNwU+dSmlN0Z8iQ9
e+FohuxyWHmAGh0qY10Ohax02pl/2UNKILz1xmpViA6q1XEP+I/dfmUM1RxJPoUGQpVIS0DS2yc4
twmxiZrdPEJKo2qQj+5RfPM8RVPL7s70V7KHh8DAVlni/nkVFbjwUGGj57w3t5d2DfM9/Fn3Kjaf
ahlmEcjyFAEYPaJTA8HTnjPdyFL5ZVUelxoJ4qBTEPa2NiTskrvfSl4J/SQIxZB3nObSVYI6BN8A
UaagBgf5ruaxA58EJ/Ie49JNLX0MLKCjPqODAxS2tOQEGkw+KM32Q45pjzIt8d8HBBar7JmhZD7a
u1flXmYbC70aqPNGTT4YcrQYnWShu/iy3mabZwTogKa1TBwCW8teNOZqT/8HeNVRJw8EemPNKYpG
CJmD9Y36fYjB+Vq7CyRfDfoWs1ppz8+NnnbB2SqN89oWqlnuwRDc5BA+2dJICZhKepzH9nqf+Mx1
nSORHYt3LeX2gJbKZnz+Q6sEna6rA8f4tZgMhkGpYYrRaPVor2GD75bZtobVbkZ9JXmwBcXWr4X4
Hzkhc3kT8qzKH91bRiSqdW/DEWZRf3BIiVBUhyI3RHGj70kfj5H+482UC3FJQkj/rRlPuHHG2buZ
YOSUjeLqoaAiRYnIEgYUXqx0mapWF3za4IF7LVNTBBfCnmePZE1gmHJekYaPWiQ9STFKR/XHs6al
cNwKJrHgIErCTfJSJaiLone0fkOIVfthc1y2fJI6qbVrMmJNb1/D2SPxDhgRPd+XH7HiHlQdeDex
Piaftjs3SuIENm/RCuGyoIFo/7HOhWocC+jWl68XUrcRR+KTPOpU4OtlL88zpwjCs4sJPzgLLQ3C
ScPOIbBNJVvrhQmoQFynnw9OryrEDtAj61DZ/08T1lGMYREWpOaFJM42C9EM9Eosh5VE7J3zMAXj
O1ohpO3LZjbE8ShB87MO164t7wSRT01yVaafy4LmAB4b8l+sYy5uaCiwku5J88HeeG0hqrgn0u5b
4b6o1Fc2qFZGyPg1F0zAdePLaTa40Mbjn/85nckS6/aWPQNEyDjy4GPOcPgOxY38xzDNaxBP28zM
ZlGGOGskDkidRMtkD67OPBzCl9nnNGHQb+o/6OwnA36vA9Z97Bcg0fG/8W1fYtbCBYpDPzdhF7fm
U5DZLbXMsrptVM026Q5FXjyQRjk5wtgF+eRmzj4CZEk9x04rUAV7HwANk78NOqne58MjQR7D73ni
blx132z3fObGTrjiQDGwanwakzxssDSebr988IdMjxpwKSPQ6E2kd7ynMtGs4tD6Al6puWMaKbCV
OOadDIccnkHcibdLYOY+4Bwd1EZRqT0v9v+MKTulLaP0NDH4cSl6zigK5niZwlbg5ZFQQa47E+WO
MClGUt67+lCOMpxlDRpDOIJja4rBn3BitQNzbuGm01myD53xjD21n0irqVn1AkWWkuYT/UBRZBhV
91ywGlkwa4mB1Rbn4n1d4xkjCQTyswQo7eYbmvfq/ME5mLDXPLzoMmlsfLvgxcFSbS7YVGzEHBj7
NyUMPG2yxD0Qxj2JcQCof2T6MvooEQlw4BbqSm3JBpaQnPgPErZ3onPOM4YV4uwI5utx89rxldhI
POwKfEKNLJYmNwjT6945m8SAHEcW8KWoXR0w3cU8POwp8+LYmLtivrABrNHVWGD+WW9Z7LorIyrV
2GHiEe30T+BiAbQ9wPlEhDEqmvGUHS7p4l+7MYJ7sG3p9DNRiM+Wh3DpMvcru7F3IzEQ0Nr+BvVb
Ca4vrGqdjriXybHp9hI3o0b5wKqwQ2J9MO2S1cO9CFcv2nhEexvRepnNzjI0tnCEiEazKQ7sh9do
Ttiyw7oi1yB+5PgDSfgKT3OpoWsfXfehpIAygmLRMVnXdlizksVPgjfHn9u7uEr1AXyG+CHTM0HU
7IZn964BtLY+C0szNRIbh4piaczmbTsOAjKeu6205ddzA85fF+4PteA+d8HpIMxiVq9znh315eVb
9bKaT5YTHA0IUOfAooiK8/Y0UZ5hdGg2bYH4JfS6D6lnswE1qGR1fp0SvqjhevAUXB1M9cQ125E1
z1u2uSgP6TMrPHCXVU+jVIBBZ43lqr33g7uPUM14+nRYX3X/rdNdMSGy+CVMaWoOI+YGgQ5nG53M
iUCYHjsrHJW7eY0Q9YTN+xhkz1R6eiBU8jiwQ3pzynpUfrIt8VLqSFRkr2c5UL8raTyHXT8WuEkm
UBHgsmOnFB881izul/w53iSNirQunx4onL4Ql3nS0bZ3iO0hBdIBRlU+fbJRc/eGwgBgJkyJToaF
WhcQGyX7T2iwh/886Oa1r/AV13fM/AsvQKdp+3UeBkJ7Sy+4cxqeyNeCREdnx/AOWzzwcdJ/UQDb
3gVkCGNORKShYz6x9+N0S6QaNhM6PErZ/2nxQ0VN+Zlt5RTZ2apoEymrPtKrPOBUgYW0jQhk9e86
TvfiBBxdlUI+rOoyMrr+ZDm5QUuICpRIgd4J9PoM5JCs2AYYOzQpmCk0Kn/tpRCYVrpLbDB+Zi0W
5lRW3h/q5TAUo62awPof/VmGg8FKviyY/ntXY3KFLWE2POrd3tOzsz3cjnJ4h5+w4962CujmHQUP
kTsrscwISZZWyFDFKvbdkUw4fpVTcuUE8ETOtIT3oO1PWJwI1pykaPFRZD+FHbQwhsLro3g6o4+B
Q7va39+r82ujPwmiMRyMOFnxzbpGoGxNxs3ZCltGJCVBm6zA6fbScsQsrP0MNKLYQ9QCbx8mKQrs
copue6NY8vGG99iAXtZYnADTfVuBgUG22LKVKO9RmhZ1vE1Y3yrcih1wlrb5+Or4fu2S/Nu8MtDs
djStooOm0nIGAy0PA/vTyE4v80mgq0R+QUCZ8nuF1+H+wcuUt1aCNfnignVXYDS1V4RhTcKZ+62t
+SoOgGZ34n6lazSC6ivbKIi7WTJ1bpmj44xYKu78keVcumNfjTFseA0AeIJ6obtzzEEjeBXM2loj
YVmhfOhjckCLRCxREgsLIXeZXUnWPVJ7uRhOAe8Li1lIujOMDAKOO4BSdS2PXjB8Uqiq3rpxbSSj
dmAdkFPFnq3b24cSkXEa5g1GLaAUPmpGZxRSaDsLekxh5AcIcTU0HifiV0oy8v0XNBo5ztrzahHa
3RhwRC2rZLAYXQeHEu5JljYcR9h6667OMRJ9M2FGKiWBaNz020i6nFvxy9GXb1Wn5k132/4+pjB0
BUb7za/aAgfryLRj2pwYcjqiQpUnEhUeJ2c5mMGVzas16JIVoYNbzvdLFSzVGB3th6zhC66VNQNS
6owwg/SncB+WCC2+MjkKcBU9qzh9WzEVHcsbKSOo1rfYqKxooKSh8i7NF6yNH3vFvNTbVjIDEoxr
lwdm5rRLxMuNQeAqdYS+9sWYhqh8s55EOXC776AhyghK+3QPChHr3NehgC4mhwzxJmdF33tekJOI
fieY9Mj9G7zJzofO0+Nzmf1AHn6KfEvNbld3NGHkf0lu99vZqnWrdycZujORdp/K9g94bQsDyjiW
W9AjxhHF8NnWGKbkwXP9p4tOiMAiCEgaVnq5fVRk/mLhkw4jpy3uOwy7n+svF3+RpC9vmCByopEu
e+oeTNyAsBrhbgGYxlYtCZZVetgTw9+MO7+ZXHCInwwe1MsuNP2rh4XSmoXcZ+7Twuq+jWqjSiID
kb5aGQpJK9i9IWyGNo6i0VI/ZXo4RTfTWgzvOXZ65hAtp+ooww01h0CT2BSIoAyzQJv2Yy9z5hYo
xjyasxaXcjf3v4/kTlF8sTAUDwvVASpPStmpIPSvWSynEFZn5uic5CwQSXrpQdUiWR/ER/2/4RE0
DY9QcZIiBVYhC0XI+RQZCLhXyO5pcdkKj0IgU6+aP8smVNArM46GXteG2vXHkbdYXU4PT989fmWe
i/M51QFoZs4nJyheWk1B6y3tZf0/OKnCMSp5Do6Y96lC+CS4txB0aB/RfMXrKcve5IX+kaNwHwRZ
2WAX4fNs0XeC7mWVBaUKCxXhHnPyeFQ3mtM7EZhn9lD4EWjiqg7eOZcYShcxwZrdUmz5mwxOQvOr
Ju8N7FQtRn2XZFvoC3abY3e6nHT6ITcCsm9y9h2TT58WMTXLqrp1AxixJWKpoae6DEZRoh4VcvG4
60Uf9rgTSU10B8MWjXXVRMieOwgcTvYN41Zl/coDOoAZneniGW6/hbI+Sv89KeS1ZWxoXR54dN7x
W35+xobPCAmnWhaXp8cn2GivVpiOikS66ldY48J5tNkA8cGu3Rb+aO38J1jyDNZdMECTXJ/qtwAw
gPiR5ggol4TPHi+D4RtHYqsNSbScx/iihkAz7MdbmkuCkMvB3mrTTczZHqLFbaPqEK4rC2objJlw
QU36D/zyc4d40jkQekdjXTi6M0y6r73+saR8iMiaafp7zb9n8NqosiMVtrh55586If0o157mmHj/
cMZ6SkZMbtEm4q0nLFjLJvZ0/HdeNM721aytUW98tInCvMsJU58hh0QXXJf6z5QKH0Ajt5sjN64b
OAW7B8jX0zOBRx8xTCP4yrZlihsCLUyzFmacv8Da93G3BDsDNHtidyXrMOF1Ky5+Xa7aKZaLYjOk
/jTuEyAi5z/yWWhTczT/tpFBY25C2rfdNne1LE7DNSmlP9ztTnV2BzPK+xlDPZrvJeBZd5Ckmivr
P+yOR9ndBJam75KBoNH1jHtzFpMVzxU94mN+QUkQd/wI2VBvuIdoCKJ0/8/REYAE8FDRcoL4eX8D
1P5XyBHxhuwsY6r4GmipiGRFJJiBIJ5LJdedFqHESkesUO3sggb1VV3uK4M7Mg8/MljultsPzKhR
dYeLu73/GvSgEB3e1ecVDCgNNeqqKsWd92Jhy6PA8H3sRS0Yr7Zg/KC5+i/4eRYKJFO2iReFvDZm
Q4gDKB/AsYeXacBIVJwhI0u5uAWc03wwlPGc7haTO+KFg4ACKAcG+EzcUw4rmHDtkO7t5ulKQehD
anwzdRLAqFHCqjcmnBmsjhGRudBglPm0GHZhPfM2z+vxvWmI/6NNpBTPGJue58GTPOQeeeh1cmqY
KuwBIka9Q/HkgzY+t7jB8V4efok8pa1U2KaKaQ6s1/W2VH74FIEE35MSf68TYb5/6gFLxjNSYACF
q51vHo93dfXg0HYGhSCCpZId3YFeTU+EUzkJ6Vs7+e6Nw59o4u3yfgbDPgYx/GCqKfxV9+kSlpGy
eugKpZoE8zCh5exyxlTmKxjFy9QQIA71ZeW1kHEBfol1fwTnSvKyP9OrYSDF6lzyrF3yO17tERn6
dcp/QfSZ3v4bpNHhguSF7TKb0c+ml7SbUVMR9kgnvnxaVQxjVUnDO+CdPcXpWN9hPyd5lAE7ej2Z
GZFjslvUlzPQ7EqqMGuSDv97B4uAkzLXaPKsxjvkelanxThizA8e/niGznn0V2DqXWiU5XltNH2k
jgM/l0FjraX/v3CwTBXp13700KL+Jkipb0uOpblXcrs8XRl2BVLCinoLCUZt4M99ErVSbVNL8JIS
PfnhmMlteTJ3ArxfrDn2hTNw3Mei3sGs2uAA1+Q89rh8IbOKDwFerkrN45rrL80wWBE3TcwGfQwn
iD3Aemb6RdSnY7gmeP7mXXuApebwFOJqty/g3sD+cvsyBYZrCHT+96BeRCCqyPaqosvzhS3KFq6J
UApHtiY0IFM1Yo6HIuz85KIKqYWdRodNGDpRI8BsxJp6/+hmePRaC05zhBaoCgPV4YQ6lB4OuaTb
73eCsMiUkiU2rXaFgitsWz1a2n2VeS4igojtn0FeSwwyENkFBk2Fhp/rF9eHSqClJcDpGY+co/XK
LjDOSAtdlJ8aTAsgRRGqoZgYfKwkeLgykZGqkMtwmYW1I9FyKrPbrrY7MZrP4dIEEsTIMfPy/Wkf
TpGZ02mAzSDyvSXsHlwnXlxHWpuEy7FR5uc0nyfAsJ0za0OSeIK0VwNdRmAkI0sXBMdd6z7KehSZ
n4bPgG3rRWiqX2wPw/gI5P5S0tvgOpRcveZkl6Z4P0CltfdqbqpkPNz4146qT6zzor65xsXE9d4K
z+xUroCOJnDOV2a3wNr+yMPpfHuhNeoW1VTLD4M+NTOfg1prVv+089E+jNVeKSu3+jkQ0lla6TPk
2BTmggHiISztmCxf0SKGrttBj2Jz7+UKH5luJyGNcG1KaSW6nmqB+Bx4T5aQl07MwjIwhf1wDPsF
ayfGZ9tDE5pa3J5cnTvmgj8RiSHfVxR8XbNuYmHuyCBoO2WDrAgESxy8rDy0o2/zF+kTNIxOtJ47
kRKgLVR1bHfjaPjyV2fYCUpN0iHxC92LVay1ECZuS9smvZiAF2qkaq6oK4gUGXOlWfio6XavOUBH
EDnDPJgQSLo/eu5mTp6vRTUtvM2RxcX6EEWqpNzJE73eSz13Td0xctIUXm9bGACoUovjRdy74wgy
5yryBvG6SXZUbaeFIApX3Mz8Pabs5k8f+f+axUq1L8q1nsVSkLPxihSul40OY6ISdo6BxxgaCkGR
yRjYsWEaxdtPTq+AqKD5iczjV2NaiNERzWniwHeWpfW5myaRoO4pQL/vuWS9aCUSDxMhz+TUjqhw
1+kGpAMcEKAhAba7tUDjvq9A+6GQdqY43ZqUN5mTFAganCfMAwFRyTZh1X1KvC2KMP8orRPPCliU
JkZnegVtZQSEsUCziLvLoIV0+I3P9YhrGd0sMlyDrAndWINYO02mqtqEiUSb2Ood7ZgHsppO5Itq
uR/La4Vx06fhFeIFGkh8TPoXvnlE3WpTwGzpcHwiyQqPfeXCMUX/argoEoH3dGtwgguXgVN1iJCu
cefiZq60xn040F0ZLF3OR0tVMViUyVhbsqJ1LpYLkytTUKLAD4mHbvBgAALSqXyKyJsp05tvVT8O
8LNQ0i13yVWOhrSUoARYKG4i5reuNKL9VhxD4DfUgVvsaEC+Lx90dSZ8BR+7dW/PMEQIjLqx/TvL
r7Hf5VO0Lil6TAQJDM15v9H7EqkqmSVkRozrI1YeNVXA4IaD3WWnQMY/7y4dzdCZ+AP0k2rLtAOj
1H78gMPhsf902csxgKEW5ebdyR6cItk0tO1adQd4D4rCmAxK8ogxY9YMhW/imAQIhrRWe7nhtAz+
oQS79qc2LPoT9hrpKhyrhtyrCtB50tyc2bOxV5miLMWukb+xm0N9NQnupGLhhStBvTNVGY1wyCbS
7D1mBaY0g8I1x8iKNjj9i3F753k36XUWBRVW6XBu0kDUX3ru73DSP4Db/ychlWhTV4/QETeY2YY2
1LUrhZQbc+KfPYfms1VicraNNeS4SFRLVlMgk1xgrQgHEgEKQShpY/EFggRcn3mYbzBouruFFDye
lWprM7cPMGxe+oDyI6NOPZAifcG6pH7vVUd6LkZ6O0K8rzuLx8/aXUI4TP15pyZRIWB0pTVYzPPr
XD/PGYUaiOd7oaOdRJezMyNDcFja6X25Cd7bZrRq1rA2LKrhDEbk+DR1lKCl7FI5MvxCJ/4EQOIS
KF4G9ABDMeBvS9kbOED4R9iRHsJa0cIsEZRG2xa941yJKDD+Q7sbI5QOZClwVsgSRnytlxs7KbH7
5wNaErJeC4ZxdbbhMed8vTrh9mUpnbY+2W9YwA43cpzLVZRnvlRmRsJ8QxVuJmHwAD1WhMN/XuNR
HyOrPegZS03qRmLnk6W80fyat56pWXcPFSlOOhllnZM8lGvVonpTgypuEfT+2Kb6BmAbnmPFiW3e
ydUwr2i9+rJEZm4XvyWw0EQXPXqiucC9yQQ+f6okZt785zv5M0UqBO8QTr7lVqgdlMubT7kRA/Qz
N+uz4PxYY9yQW023wRZ7QqekNsdWh6JIgCiS5otptyDMUkkrEMY/CEq5BgbD/FGppItsP7b+i4Nf
OI01wJ3Y0+GaxsGoP4bRB9vNgYTMi0SBIDgoavfGHp4r6xIOB11ttM7/LFeQE3KXXXIjb1X/tC3B
3mFbvthy7ZdTwA7wjTETeKJyon/E7bev/xYhAQbk8YDUNIrgpsw7C4kv2SGn9HDxwv7F1T9/lykY
yjFSiH2FBr5yATWwHgpm3mW40VRO/sXI6SQW7zrUmv1Z9QwaPn4Sa7BVkBvWMaHbhBEojPAuJSm2
OLD8CyOXdbWgt8esjORdC7Z3EYfjECXVyW1KazF1sfA023RC4Mju8NOP82wf63yL8Q6VN+bedsNI
FF1T8EhIw65EUoQfgb+Vfksm7YtPqut2QSiAY7ujIUUs8mRQ0SGdZvbwC203Y7qvnTy2LqCGP/zS
FXFhjiRoBJrQTsKK5/6SPGDitjYHvBi4ip840QarPNUHp2Ssx9rTWZgoJUZ3CkfMcfAWYw4BNvez
Ulk5juOWCCEpawr/RhcKlD9AjntgdgUaNMefh5jAlGxhcp0moRBcLI7tF3cqsCwUYvBG6VTkgisO
lXHiuWZId6FmBI+GV1mFXoeqUIgQnrl0vQYV87l9W9zY3ajAiVpLIUU/L/sWltErez9viQNdj0pV
gvi5nzHmqLnVRD87N3K37CWkBNBDOrpLJCwWFtQYX8UY6uxg23kDxmTWUkurZR1ygvNTmBbzsh57
yCXxpZF700Jzr8xZA8SnwDJLcz4CsjcNPKJkbor2nOZ5dNcnIypmclDhZ99obYlSlJHKo0tr7V3Y
NSQvkN0Ea8DTgSK0JUEboCBIVFdJDYeGdaPKivlkBenkGlcS2XYB+eQjYLhhswJLILbDYfp8Diz4
OQ6GJjHzifXArUg/xNr5I6d3KjT+reFosIfiKZhOSeu81yIsyVLdSXxceXZHBuL0fV0sp+u8NSWZ
hSGh3rkwEutKQOZ/tdDEYNssCVuBNeaMRjgGuPCxHOzr+mt7fHL4+t2iRSItvhMymWzOaSMj1b2n
9eqsxtshpcDanzE8DGsdj0R358uiZu38vntjeAa21xA7hGqlJlhirFXPeOK7sXm+gj+b2dtgKgQU
JvSlzbT0F4IbNsDrG/Uq9e/LZTSVLnIfRN7vRco84XMqZgwWvIl5sCm/h0SNui9LFwbCZdW4mw3o
pYh1fLoMuQbErWHCyqhM+3Y/6dLJhd+Ej/fl2/7htSfgZlm2YiMdXJijigfrfOP/8Tojir1wFxW7
gdx1Eobp45uIZ+2MberpX8keyXvva4je+wpLX0dbaEDRlGafaKfn1aKty8tj8R/ZxfqIkpW8K5wv
ujebfgS8iAVRz8FCbaEnaP7gg0F4u20QWKZ0cvVxiME5d7YLbmmgePrtGIe4L6ET+kJyVZPhuPYD
4yLK5TRovGStyuh0GgCvU28w1MqdjfeK7LIvSoTcdLIJn4guu7gWLLZSVw2XmsCRCOLnUGNscHlr
i6wNG4wcAiuwZ5miZ1Pxw1B5VC54cIcW0K8XzrBuJBtKGp6PXfq8MphdUK4DgE8pis/cRWD8raXf
KjogmFP3Wsets77AO9FLjRFQopbFT+IZBXN8Uf+HfUX9f5XomJ3WcCLauVvfjSuYzMsjENzqTQ3w
9leeao72YmfNxbP7yJdRoaKkf6L4taEdf4134ekdkY10Wbo9trvqSGq5vn1sq7lV7TwjHVuXpdMJ
b/UV3g30J8k8LN1sdkSCHWNH2KOVB0ES9UK3gl4Eby7V8JpJ+mdDB/qY2zCAH5qbR1RX4tXh8Yrn
t1HlLAGXj3/zZ5VJJGYbJjMLpFVX3O5unV18Vj6PasQiyeCQH9wf2iGW5uFayLIEgBM169ExUnHb
Zr5NUntS7Zli1EmA0tkcxHSAaklR4/5S1RfvIwDA+A3r92Fgd6rhumRimc/D/7bN1RsQ+UZLRZxz
T+RdpL2YaBQspfZwCfoZCcKloLGb84oRC6ez0bbZlndRonUfT6Bd1g1wuE1GuEwlsMy+EExqfxje
KCKyyWmt3CwJn03nSngQKmTFD1PxdUvd0t4yr5i7JQwzSx0F31Cyq8gq8MgPVWKE+6ZB/Dbeq9fA
OuvFqdToO9DebEBXZ0un/zsYvi7Cgo47KChsf5OERoGiESfT8CVolqe57RZUVclbAjG0+/8FMIDv
78p75dwZlk7VvZ31reXrP3tHi7MOlNCp+hU15Bcl8zdqJ0s+ausx554xhasZ/9TI0OI00uveMJyb
bVrO4fs+slBRFJDj0S2dXUNSN1kXQTWsUFCuvK1ziWiNZ1iNZo0YDQzPk3OuU4uRD/dt1TEyXr4N
0qW7E/gfVB5NmhQBzoFU1SEJtHi+ctcc+w8NwMUUNnLr8MP16vBFUBYtb9VmZAftPIkzTQkU9ahi
8ZOeWhci5bOgWeZuvwrW8Mwcdcj8OwS3xOO0BCH0vgACbwOH1iXLhaUFXDiQKT4lxv4Vm5XVW71C
Tad14SkqPVH8feuNnZaAzSkNvyMmxh8FnnRQqtSBzuSLlrpHgyIl3gTYc+5JRSTJLiShir6uUmJC
rDDqA52nintWhDw1qKFq/A/RwlM8qr+oP9nStOGJwo71TaMk2cTU5s5Nh3KC8AM+laIqAzFtYYi8
igNc3Jlm2cJMBT/bO3hI8skbnTpnBmfXEHlXRW4K9b1FNiA7FKiQsmQ/WuXxFyfDXOothRZAJg69
3U8kVJTh48m//NVxAKWQHiVovADxBvbFOgwAq+ggGTWI8Ov1nF4p0a23yp97UKLttl4a4OKl8o9a
qerNxmIi9usfr9HapX1dIdwscmBIX8HX18RUipjyDqydUOsSaFX6FA3b72pp2WBIyXmxIiHXaCbR
KKKSa2EeM1IcbZUqpjVDAYPnMZCaqcoCX/7g9RXU+kP6MhO4BAXSDAfLltd8uiSFZOk0BsTjnwNL
7iuW8hruTxJZxOy+tsfze61ScKx0SmjJn+mdCD5GibvsMN1CkKr807hWfkRK7iYlR6aiSlpnLtGK
/Ub/l0iP7R2cbU9oBTW/FpeiXyDwvERo3dgGsI1PX3cb6K+MxbZycgHDbXsfpGkD/Y9Hl2iUOW/U
3I98+hLAtwrfubnCSTZXN/U0XldMGf9B3T9ioY2NxaSLJaFbDU/5yAawTeuj8Fv3xJ4VyGLv5Ygi
DC6FqoaiPaA/QHHWmkFRF1ZeOf7oyPLE/rX1m8R6sPLVkcaraVhWpwFhMCXIOKlzhtqRg3breSo8
DyyCNfNRWixVngp4F6Wp84oCJJ61exfXWjJoWeTI5EETMR0v/wmo2GWrnv1HZ2TpUKQMwfuCAoQs
tGdYNWZHqUyxVoXSo+ylzK/ClbaYC3VsX1lEErjo4wdK07Evml+//46tlhNKExT8YDFJIWbU/Jjs
6XNUlBPMBTWuHKov0w3tzGCwwxv0lELCosG/dNvZ53bs3lAaJbV7LSSc4rK8zc6d7sKavLRMUKrN
/HNrTH1z/Ex+YhYoGSGlbo8W7hy+9ousya646BWe5q0nyZNABqIkkT4FrVKqWuD5MNBvrL0IOwGP
IHZ6OoGmpICT2wnRxoMb/hltdvYwwH8z8V78E48ToYkUcffh9k+Ed/2zoXTr0ML7/1DQRwJfrF/8
rvufgNoDfC9g3obexmYFTLEVz2Fguyo6UfQMnsnJX6wnpcev3ay2BoFsJLAr8F1LGqUqMoKE1ymX
+los+eTFQU2YYowoMKJL0O89ZE3XEr9yUWMgTuhT106nkUuo53zh/hFgIqlMmUau+HWDEHu8rqa4
fD7r7CvHIel8CLBguYQxWnNYoO+WVxZP1PmWVLblXZ43PeXCCNY66+RTcluiMbTSh0eYeV+W+61g
ajEMBt9fN+vB50b+W7s08fUJHiyGDUaLfPj1Mvuca8H/2sDLvKV9J2sXG6OgdLymeXf1KUhNjfUa
ITO7HFCjlUpiHtAIeBwXxIrhdCSzRQ7k/a9AZvjnF8aJoVKrkjzmzbFOJxSkJ///RJZL0UDJWcsz
h5hurAIoqxNmdwRnd5hGguAB1pX/JVd464WmMSbWIbq+LWqTnl9wk2p0rG4wJsVWynMZu3mBn950
lEGZfwHylh/TaWBr0OpKG9RojSsy8SnXGM4Y3LBQPpMNBy4znTOSLurAAX5ihnerhwRmNLRd9/qg
RpcjwWBRNg4WsTrlQv5/Ln8b8E2yiD0T8cNmFRXlsmtgARDvKjJwfEPm8bDWc/lJvSR4Pz5AH3aK
xVCP96f8Xx8G5pe/l9d0KjP7rMGtqpXIM83Dj2U9hmu9irwNHYnJb1/yJm3xDVTKqsNxI2E8Bl2d
++FyssOvaynVsXPII8hq9s3skXxvPzPd+jZh5Wey0EUN75Myr+ZGuYdOI9mS+DQMjBv24k9IzSow
NM9q5Rc7OuZzE3o8EBaZAz4zMuaAgdnh6RYexRGoHX5Tyy/XIMCGQmiCOinaWyGFYQVfC7NGcsFe
PVDKULU2KFKxEFwlhCumtcZQyOL8BZSB6ECIsj8LWSbNEniDY/9kVxVcn7Ly6e1jU+pheoTBFsoU
idRUqypIh7Q0060hO9XY3SAT9nCa0hBDlK2g//GZzFxPwQqOucfpTRygFKpGyvAjC2o0CbZTgp1E
zguAg1D4bwdS1Jw8EdQwJgAs/7Erfjzq9c2ydGQaJslGqwfsRkaAYkMC3y4Yf0Szo63eWSFRHt9r
3qNBiJQtzF5dRdMT27GpXu3M0FF3M9iulrwBOVADmfrAsMMBCShJiVZeQJ/yoRnMNbTumoZdiAoZ
mIDMTTS5iwXseWluf94mvxPXfXNLsFILD3D7SpcVFyH6UoI4lFs4AF9tI4vRMgRI1pgzBxgSfBFX
/SpxTcnVYTSFERt1nUiew2YCSH8d1ftbHBZcsS3nLC9ERqRm/UV2Qk/7uqs7+RH7rldfWKSmQt8D
FhxrnTkC+j8BrC2L8KUWGYgbys4fUczbUeULwdaNLHLogOaqlVEEq/nXrvNzilqYi74KntAcbt5S
zELq9SbsR8xe0wgSzMvErawZ5iPfR0nv0+BC9L48SnmTAUt3SrxKVTwaP1bTkP0TGuKCa+jxA/VH
d/JC3uGyynG0W5SRl44QOwUQe4AIV/wx3nyldC0IXLV3yGh3XhloJTz+0pv4otAsubGRrOy2nFjG
KalbhAzM93UTYwDx91PjoDUVSK1IKSE6c4U/jRccX2Exf9mFlPE3LcLWpIYLHSHixVyEUdNrMdWU
UREFIrhSnCjWFqokjZl6T+Q5N3QCa+qi9IzYgWwCyVStOFBd9fpTPbIe/SCBTH045Duqpwy+k5bG
Uplt04S7oaVi8XpZJueeAz2H6WdszFKsDw/oHzAw74UfVoV+usi+RQ5ojYaJATI9onWfvL5+y2RS
7QuVsjUx0GLP0N9xlhNlZhDYkdKqCWdwL/7LMV80w5Z3hZTTXq4+vJWSG+olOECIZQvdjSLGTvuw
8viXdj5cUWrgJwmJe7WXPAgYZfbL2ZX+WFDeekUo9tMHAPSJAoloA7E09o0AK+5dE98wZiPDUDe6
t2rgdeMrBudUfMG5xPEzxTqR+x3BJCICltnvsIBgNIi34C2YFYrr4untvLVUfvbyIJAL6x+PpBJr
0ZZ+748+gvmqaRjeD10UIXQ2aYXby28mHZ9jF946vb7NcUhSX9FAZ9P9Xn3XNn917Vxzlr5cMIpb
HTMNA47mYJQ5uhoLExOF2smmuvD7hDBSoBlbzd2f+2JKrNgGad8uu2Dvo6VMsghiV8Ktlw0KnDZM
st5ODupdqL6JNznE4piIUTMo5IPVOIqQSGYbhv2lQNYjBil+AOZLebY69Dqj9No2wjq2G+FOGqWa
4EL43zXkh3uJ5E6LX7oERLwFW87dvE5Yi47ocO4rxBCVlO37itkEVJhvdX2u1PtXTdYNG4Tc6+tt
N0H8sjoy90xoRn/Eft/0Cij38VtWdPZFadYE0XUqtgGDopE6hQZFz95OhXE5V4iIl5wRx01KD+eo
ZMHDI0HdHCZZc8tGccZQf3Fmst1lczi3GA1YCDO8Xp5ivocnOla4xdcSnDv3H4aVqMhZWx5nlIb9
Uo3dKGdZ7lnrj4yG8MBo4284B9OL6LoS9DS3dlc1Ob4g5zcEY25NmUJVNLVwNLDzUjdwRTSULNtG
6tg4JfwnWNBnTKjemjgNJlr+m3+Mo+I7dLjafQBnQ3WtpfNff6yNYPhDA18rHSG9aGtfbRgYFMg+
6zytDj1SxxbdONZhfbxK7jnH5FVliWtP5+YYKCErzeRaqc7+2zYpqcDZO/wwUBT70dt0hksIcRT6
co0HkNTxCwl4mDDcd8qN91a5avTs7vKMLOMPPJznBPM7qEP44w05i6Ermod6kH5xNLfLaAw7MCDZ
5CbaHatpu6mhfAavrVTmrh+/Xb8+Qa6apKaQejmpFQ6BGcrRykDLvY5m8MaY9EtM4kAk3GDVNHiv
BB+BE43QkqdwyJDgNyGhxgDKJyM2zI+enOoAJ/36UrVG3hFJTu09RGsTjO3aobC+rnPZe/ZTUnrB
vxHsFvVgGECWgeMQAJf6/ZPmMcvFk51GvMm3IJMK2eRFm+80Ykk8/CmDL/7rSilYEi7qK6ArmMJq
dg07jqpPaQcjCg9OPRrzMZk9sA9hKjYtwCLoglmGDiW8tIf7vrNaUdg52jkOnGWkea4JYgjeTI/Q
qJKZN8LUju6JHWrHLOkWbQDbo4ZWLGdyp/K1VUMvdIQ8uMud8k9jk8DWE7Q+JgVbnNqrNGDkHMs5
zpClW2cKeKua2PrFd9PkZLw6GFRtugQJY9BECbPCew7JH63KfNVbQlR0Uo6D7Onn0qemS2Wn5Jqo
qUhbTiO5Lk8U/+2IDEdWejwlGJN3hI0nWpprsUZc/2k8Byk+yovGKxWPuwBl6Pgz6/t1BbuS0sce
m8jM4DoJcSh+2ogOv96ccI0UlmYtvjQ4OBnCkkMNL2uJ98+FNk6hbwcdGyLew5Q2wqGZUaoTXfyD
KG8573RRRvDtqQw3/nzd/sMH30wjHUSnU/DNbhyeI+G0A1S6iadCXuEeyMttCxNe8zMU99/2TMMY
STfSgyjzCQaZ4Zsa7UY4jIdqkkzk1P1XuLE2FUq6Y6RqX9DwiyktHP7zlJoV6xPVXJukxU42k/eq
eyHoFaIBs9eDga0y6PJONXf0anzxBjJwcSd6ky8U+aQ73x3BeCmWqtX0O7dtu6VTGv/ev+rQIIsC
RVE5TwbA+kyUC37XuEUuawCcns1/Sng1ANkgPYDd7xhzH39hLPlOg+AYOnXdHPg2hW1zC42y+xfy
hlOmsVaYuOm+7Y/yc+Hr4hWfOtSRauKVT+ZTVTP9aA8eqP1+WmWjrRnPQPu0mN8yKdg49JMJfnTm
m/PuNMyj/vrZfPRuKP1aaakQmuCZ4dq49LjXyTQV4DnoZgI+lieAbvm4s3R7UYr1yp7uJE+WBOmF
6IUIbVfCRcOTt9mnXTZ5kuNob6VhURXBeFqYgNplR6xGIFHtqAshfXF9UHXNACD7ORl3jDRAJb8R
p3ic1P7Ycio/XyuXxlKiAzwIq631y9kOcCILvoAAMf0c7xZNbhTQFWVnVjBK8vIQ2OUMcxTCMNBN
sh+0ZAzcD2X2K2bwCXj83vQwcHtn493lpeZsKuc+NpaxoIyRr63mnzMQSb4sG77nEmE7q6JLz5as
oI1wLZdFgx6maXIcReP5B8T44yryyeuw3qk7MeVfj/bHYn4w8DNg3YggiGi3cL8LSeUfF8hxyRAY
Jqj9vZgu8XEP+sLn8MQy6CrZBiF1MELgaHTNfo6MrkFH7t8Rj6tuieREuMfKtbfTWnRa3/skkxKJ
WlaLRamfUqQujVy9IJqJTNMwMP2vK53wZhByxOD4BUd99FvNJknR4idncfK7NGji6rcD6zy6ym+w
CmOQwE3kdX7RZMo99psuCuLG/8KZBoyLGIMHSCqRGSXU3oFVuoIphBA6Yd2o8IFVQsY0ZQ01X/rw
gWidbX1C787dxrf6BqTvtKWEcharp/T6oPI4mX+aVJLCUFsqJynYx8RrDmhTU4kldLaMbTkwgsZj
0ncy0+Q+Mp6M2ZR/MXxAibErHJQpuIvFv+X4Ze7bA0mIyy/D78TnqhfuGSHWUB2D19jqhun02w2x
TvOKtK+FKiOdu0ON6vBOkMc0j+4UU3xmZQj3mfoPBrcigkXmsHTVuhWLUlQJxJ6z+8i6wU/iTWlp
t4bs18YW/bpZdX1rJK+tiiSN+tyPzLoMZQBlIH229wELnNQSn1Whqqb2KJWgoHVHLS1CV7pTG7Xg
0aefuwZzUb7P0x2IH+yqv+wrXdLEekAy/ow6LHZBn/p0if8aOwISQu2G8APB7Sd8haAylpWztvXU
QkChzSplHVltszzj8wrqit2RUGjUUGAO8Gbn5HcEhWQEsukXDRExP9N5F32K0Lxb7L2D6C7BM40W
A3vyYCWrfSy9EXfOyXXG1ENSwMogrfjkJwPQiu0hUxDc3+VBpT4AkDtrZPktRISXvyijHGFfyB1i
wecWIK2OZz/IqUT0l9Ft6jEzLaq0B3gbvThNrpPERqVd6a+XWWtdnUeECQC2zTnzWmrsXpyDPa4N
V+yWEvauLGERKh6kKCfALRtOsIXCzsvwq/uRsfnYrD7DpOhWT3HlycolCjEDkAEr/eN1MphzDImc
sLu/kPVAloiziZ9ImhdhOP9tgi8HM642XlaQf8Op735n4oqi+rQdD+eyE7QYzLUWbstYDU1d7WXQ
h57tw81Qu6id+BGwnshOXNIP4rOYSQgxtA92sk3383RP8wDgPZD9uVbrpXdVNrhjtuMX/SjVNiFc
Q3tw7W6vhGaT5ab3+tOLi6B/eoxE4qY9MpIztjIwfZkXQZd5I2kFaOdfEhjsGPACVHsHJ5z+4pkc
33FXT4yc7PWbE34nQ2fG8j4A/4vVU7gWl/BO8Xpg+LWUEwhKdicuOeR2i5QulGKhpWOogQ3EcKMa
Cn4bGZiAfGHVF+eocnmjXrnYve//+S8iYw8H3/n9pxmwrwK0HgFq58wOq9KyrCxbDfL9IUCHaj8p
0Rp/lNiyUaQIMTSljVOWNBdkIJSRfFkQiDupcTsouuBU5BWAynefpGgXzPJQPixmWM5Ske/hV+L7
xtS6U1AN9377TqS+FdM6eZJJ0Vv/qJGW0/sR/7TRs0qj+lAUyWxbGPDWtROXCKDQ0hsiYgKBE9bq
jBTnhyy3DLd/gFWS/DZSVr3gT3regXVemYXVR+7I8Wc2cj3NkIeh7pomW1pkqGr3B5xKmqwYR7uv
jLi+pesihpiTvo/NhckRgO7RLb8qHTZYapy43ClYRAFlae9RLGgsHi5X9N119buCGQmRc6pUgfSh
LYqLl/Ev9r3rYQr31IaV3y8kVXYW0AQQqLMgnUGzZEsx6phic3i8tTbIdRdzDmMJf7M0jt4G5v4Z
SqKMKTKOBVH79e/7sijdx5OkuOwHYhOcrJFLgECcWLryS8tfFAlC6fdwS8RbH6sE4OvCfGWceY2E
fPpevg88x3/RBO6TjfbRS/I5mLScVUKUqSpH8bDuvr6vmqWuu69K7Eh2fTbXArKK2FDouCjorb3g
wxDR4BelkbBShnbRvEwn1Qc6wu696BRBJoMGUdqGyS6LZ6ldjseqP4Zf49PNJwjiebS/pG09++/w
EwGKIhJe/VrhzeXx9nsCK1d8SHq+jwdodEG/jZ6FSnosFtRiBPKbXtJQz79+6kABTagwzJofDAXz
oUH+OPtS8iu1BPCM7/1vGAb1zKpH9u8GGQ8XHRXo4JfYgW3CqZ80oBNfaxN6klgPJ353HBhCf1pB
Y6yMWO9M6d0r9FTLRhMg4Q7sFv9vyMRYMgDHtOvg50Ou3GAnSakOepSnC+hIomxR2P+13rlF1YSU
YvYwKkQLzn8xgBGxDj2dLHxeENA9WMws8BGS2pzadUoO3OzSH5LsO/ILetx0f/DkO0SJNc/N7YTp
pkbsCRDOr0A1evGuHG/riaWiE4Fr5x+h/WGH3vhTT+Wg4QA/QshXoKyvegRJTpb4KQcqeAHX4b2l
NVJXPQ4nNFDJNmW5si4ZIhth3npEf9AuLptV90iFk7DIGhNtZ6qUbl5jzrfP1Q5ObWd2/nlbmfPi
0xWn2oCRWwnqpO5O1XctnlBZP+AJuBve6Aw5cfnofMo31FxMU+N+ryJRcBkLCPCizrr19usMRvXQ
QD/Jlws3z0r0jrGQSNj5ZV1NRu9aG4OWNm1m9x+zZqM+CxqNQPDHRTYMnWK6rzEKGa0FpIeEhZ/M
4O4cBhROwffmIXLXy67c2iD+X8GQ8qTP8+hyD+THn8kmp2STa/42wWLulrzqkWlKxJeF209yJK+D
GTmNWr4CNBR15GHybkt4ybsd8wLm4ZEAuKYDWkrOYXGWhMiVwy+MoMGGRVXWsZX7/LJZ1Hm7iJF3
qvBUBdvmGuI9O91FYFXBCwOXD/8yhsiedvvE3+n7+TMpeEsgy0f6Yyg+t2555rijhJ7Epuos7InN
jw0o2tKqTij3Nsjl93V0ivP9h2MSXhACSuiqGy9axdbhny1uz75fH9JrT399TCCqz9YD02melCfD
Mo8+unsAR5OafLX4djxjaWJK+QHSCIqQfC7igh5v7PqHEd3PTz6mTr3O6N5O3b2QikRcnH4vXP+9
4EHLKsJNV+5Eb+HkopOPAoX9X6AwbsG/EIMnEkLRJRKhYyjJGnPNHBQakY5E6DbUMnqmt9Ry44d4
NmuWSHxtk5pg04A0ZOnIkN72bZdbIXhH91WT7ReQNwMweedrhVZym7yq125AKo4XfVOr4DrPf33U
+AcGd2ZtEqPLQiez9VEyMy8Amf08onBqxcOXSfcGEilg4Nma23lHNj+2T6TVLNQIV8nFvG74Sv4j
GwB4kP/WMP1+VOMNOID3IHjT+/ueDCbnIAYojqaYjZoNA28qAbqZ04sS1eNt8cmXuARCZfUNmK3S
rY0dI8OG/AHTEEIKDoabjEVl/xzYE4gonsVZ0n8G56nfnTVp4OQMLhrYuKiegR1H05VbEqyNsgZW
gkAxHxUWC5pR94hDRTE6xo1FaDU0keKtTYW9odAzwEzvQy6Bja2jzCV5HP3JkWbW9ASOvW4KpBjO
/eUmhyg2rX9CsZzkM/Balu4UferA7IE8JX7ICK5/oQQQ7R2d0KSwlXFjtVFehmybuiXREvG7tJFD
iEkn5CTxZUgFfBq+UlqlLI75ErPkcq+M+VTX75yxpW4ArHx1fioB3SfQ1ks4Pk4qrro2lK4PEVbv
fDuCeJjUhrqwRrtofB6Wy5ikPl6o1hKsr+be/hbXTWUEAmzB73WBjE0D1ZlP+Y0CfLCBEulANRXX
Qwk34OzbsvahUMMjl9fN/rics7JmMkV5TzYgsl9pGQbzlc+n7swjKefRlFM6DbZo3JI4aUt7IbDQ
aFuadApz6PJ8NcRLkqh+s+EriC05M9V/Bh6yuLhDOG9YeO8Pp+DqDl9PxkIDCfWwYaGbp9sUj8gp
HeswJWFMgP3+RSTY2/IYcRQyUtyQDHzolGx3w9fEFEYKFcw0lZ/z8ITn4SwKii8rWf9w74lWsqO2
+zNduPy5wRW2nX1d7zGj+ACKAexRI62dQYQFi6MzTCAH+fPtEdvLWt5tLffuRzdW66nvsJxuuzjP
JN+IiHHm3GaLNDVF3GX404uNxmBAl2eTHjOu7uTbvIOplf/e2E8eiwlpmTKLmpx3u/6/n2I3B10P
Gwc6e7jGmKiBCdp5FGRajlNt3LzZeUNi0AYH3OOQiVwIXUkGkJI0U00wBgCGx09vq7/BYxiSfhuK
G7FoyQUfdyUzPekvRV8BnkeBeBnEYdRX6VPz+6BzOY063LOUAMQjbGLhHctQabIRDlQ3MCM4pccL
noEJMH4AN3/UjmeLbMi4kNYih7ZH0IraXLyHn8Bw5fNAy0nOIuklT+e50h4KZNSTFvHTQ8QlMQfh
s1hTNWTQi/J2fEAcE7wcKCn589lWKFQsIL6VeAIDk6DGI+P4OWuBeP9ITBfek68mxiNHB2s+dL7u
sZbkhmrSMdRXdyav3gnj45uqALYgoErj32G6mPFPIeUqaTUDzkG7VscZpTgevqkiUAYzSSpMkUxk
IjzugRjMCt0nIgTuKP2lHkyHn3DUqm5Uj+zd/2uIqJdO8veimxjyklGcpj5EqOZILDuo2q7zho5T
C0V/3OPan2C+KCrVOT6s+UfREog9f5ArSrxAzX0gBDSknJMi1s0B/kCV9xOyp0wUxzFJb+0nvfA2
q5P9VMSp1mUPvfupXXQolKNh/WasrJD508vChTE4zu4j4j4mNXwNZr1VpXXuubeGH0aKRXgvn5U/
PBtOJrynAoNxfiLTawIM8HkzdLg5iMuNd3lyKg9C5LsNPqsbGpajlvL9lyjv9J+0H2/O6UQF/0Vo
vbgGdD5/Ky4XCUvxjYG6SNvJIj5ugiU1irWFyTjA4EkWrXc3lY9gjeBHGJ1/2bi1LRAf/lS6mARz
x2IZkyjF6/uVZyWD1YmclLnwwG3mSvaNAFyDfKdHW4nt3PTXTE+LOIbuAR2s6p3K528JECvXNJzy
xzQXUskskbx0uCF7xrmXZT3CzKSdO1q0/PDD27FbtvdzLWSw/hjaxLacteFA6BEFjfPCSFKJDKmG
EnXYp3KwjyCrnETRycvmYEgr0iwS0wXbyAGjNi+2Yu2tL7+eIDsADeNWV3q490ZQAHgWj4f7328j
gzKhmlgRZxhIkwMeS49lfmDmk1w1GRnAWu5CITov6Yt5deFHjN3pDU7EYk+mkIfBxr/XtnVHxz2/
AhbUw+8z5Nr+igeyfiBmix5vKsjMC9q4gf4FDG79rNrDMxNlajgEb03FjicO0c/jms2lAu+xZ6rW
6uI1Sawuqgqn7AVC++1TMSRAH14fa+LI+i2G2fKfAtFyiT+dM0O0YC/r8hkSpjBduPUTDfo9IEi2
oA0dmvxSmBUtQdfwKdowHsuxxQa2IGJMr7UR+UdRXr6RpY0roD1JcRS9HzBpgr4ZPhs/816hWzyF
r1T0S8VHN6IT7j49HXyfzOQXsteksjYqsfiThetWfWUMuPprp7yHThJe24Y8axRul2vDP+xHcUf7
l9CjAwUeko8+y/DBu5rLqR22hZMWQDIk7lz6tA/UaioWlJnIpHPZ5jGtwTDfOFp/OZ72N3QDtWFP
gSlFJ3e6JbHzYh48gIGKK3Q73BQ1LDuPfi/WO7HzsGtD04EoaWZx/1IzbG5aWokOjK3/+yqwi0oi
mj04mCfFSL4IbJyo6x6BJ2Wb6eP0uTN59c4MBYVxKQrmdLad13rPA5IsWH1FbWR4Wg19e750qinP
5D6vfWaS5DFOBnXWNY+yPmEYgHElvJG56O6qMqSaSoLt9QA3N8JdX3yvEzXOiM1RKoIghqyICtBq
hI0yvrbwSBJpgCxQrjS9vLVbSfMDQr4mSK/55KjPSPBwdzutjaI5qruZrpld9IFGpSMNaCCwgSvu
puWDrFj4cnQoKDN6ocZFF3DzlIj2soXTHPJwxKcUNajulWW5lN/yyv5flK7xi7Jf9Hjb1pc3IoBO
/624sR4m5pyFDSPyiewo08qX3KOPQUvgwwd/wOSh51Cly9yaoZ55ZBPVcm5T9OEclVig8mbwlix+
qW3kQFS+2s6U1QXWlfZtNOut2obBYeyIeHyLezWRMBBVELxdTuRL8Jw9cpspMkj4ATMyMcPfe2uL
ASEetfi7meR9+1EMmnxT9x9MkrogilIDznPbAAZ1MT0j4CKtTgoQZMvdTYVUzxyPFRc+9IFtzVOx
5EI5TEVyjWsQRNVvGHPJjDQHJmOhx3p4DTv15aneNDjQIUL9IELZLIq54yLyHdFae3TZ2rogtRHB
uEtmSPb0WfkbOOxIiBGppOPBPgIs63JDBWdmavv+RbHsZZtRwRvXs+g5/hY2yfQw5mRQVH9TiYzO
Wlu/+4I+Q6NYxNC5XnPklKgk00wiFASwz7YoEMpsjE4ojc/1Efmesn/goUf170DB3wEfTdveUa3N
7SiIEM/L7TIl3l2mKbepSpXfTc0zQTMTiTfkHb4RtfF4M4kLecz6kdEH8ElzR3mFGfxIL7nR2etL
HVIFZIVqzgYATS8a97Px6ilUxAD94iKUaSI14qgBhFziYnkotV07XIQEgFwZ638FIJjAY+4Ru6u2
CQzPIapDMXNPApdOjieDwQSZxQ79su6h1Bafw5kpIrXBTcxE5OPKb9em5RQ73W54vCqRRLc/tvLH
ELpP1yeD5EVOynMl1uuKILMlCuAK5Fs/+ayN7Y08oq2Yt/AOWV9jxmd4JJiPmYMwTY/lHyeNtomV
FZOpr+ozUcfdW+1cGtMhI58JLZ/+75zn8b5gBSWs6QGJib3cUhTpTEdEQuMaigJijCddPFdgLpVb
9TXY3frLROvV300L7c2iTC6yyBMvx1ffFFofVYGdCAR4p2pkQ/QN/bF0RBR4cRzllD2VjzBWaRtx
hDkbBsNA9D/gqOLQDIoFqZRRQHV/oBt+PSbgVFTT4SgXRQxb7eyQT1LlJFqU87HNgt9ibnTmjPmB
fisdV8wjviCi4RHNDGoyIUfr0TPgxhxRplS6rf88PC5oERyvC6QWyJJVFwrVhIoeN50TmrK/mLYS
LorpBiF9mZz5T/0OjUCkVZr6K3NXH9Kj3AhCnSyM5Fmp2iX4KyB3BesUnpBcGE+1JNWKtScPgpHv
mKHy7zzFFRgCXcQHqYNcWpaz72O6gdla+dnoZixVo16ePVsqLS0BP2tQQqSVGyF7Dqc/4qlM1Wz6
Fo7j6cVo4meLGQ5C0fzSTGwYjHHADRmgr00sFQq9+AG1xhx8iflJ9XiSrmVmrals+4K3Q8hrqerW
qtNnQ4HfvEhLw7Z370ze/iRFGm54Hyg9DCv60565qgqH6LTGyCCh9fxq3YU/sg1xFSJzEWf3P44M
F7N13k6XbOaMjtK5zotDSgzRQSeI31xCg08yb+kaPtS4JJbjsTJp/arfihYN9vZOdx0oXVYC1wp/
9lpwZ+RX9SYGOicwpgb3+rTs6z8InKw/e2QOGmKvJV02vWxtoV0LXX2Y6sNiMasOQePRWcWLYI31
TGXxVHWHMAnWAaPX5yZItMFNLY/4QbgZH3k04cgmCnDYpLvdNZUFmgPeZdtu/DkG8LmrRoFxqLZs
VAV2Y+76E42jCyvu2ZsJlrMQEfGbLg6uvNh65Xyehn2oHTWRqGldzDvJSvblOYsuADcPa+Ug6pBk
ujTic5AHftpfuO5xkzuqbJW5LRbum4MIAP7FMcm2jel3wIunuPskNGRRqE6JpJbPmf+IZmEm37rn
8zSYmWPcOA143OZU/b4xz+6EJ3WeiMliRzV1nBLTgZoo1rns0EDvHGTfpGiPU5hn3aotGJShYgTZ
zBo6APR5dB5SvEX4fAh0XsNpzLZwMsTqh6LXWVWxOc5XAPMYZlJgYWxeryS8HmLyDQfKFMu++THn
d/KDHMGdlFguk9LLRrYKnogBA9+OlflRn/W97k7YLiAwf3RFIl42UvEIQmx/xkJuCAy1C6CWnEAt
+sXYwe47ehI8d2EuO+neFu2G3Z4+/C3LNrUcxL3feE7WkWNBGP2ZtgDWhAtJgNFX0lP+i9bqMhzu
6Drel2BW0VpYMN4sz53XNly0+loyLS28xW27Sldvsr/j1BFqpigXIiCHo3/mFF4m9JLnrxrpbRq5
+C5lGOPlXT4qaPZEIyTIWOXEtnPlFahSlt8zhmRIErGg5/AO5Oja4JqMHURoIN8urKnge7Ftxsjv
7LdVvnNWWFtpsnXlumQG4vQ5qyE8HShjhknSNZwNaRscT2zAQK86Ab7l0GvqHu7H+E9LUsoVVg07
1ixplVtIXHikdvDjDDK5bCu4yJIdmx4mPwj9OxBMgcShJljyUwd4hAn6QFrWjMO6XssfSqlKdDkG
jWbfki2Yl1XeEiIgg9B1sPsf8fKQNN3l4G+oyD7N97AjLcGd8sB9LbHA04apMlMUguJgx4hp15tK
GfRJAGocnjEJpeTujIPelgwvGxU1UuFf5Q4HjsvtCeiZbJdRHr0TU9+gis7TryRt5z47gohrIpJ0
L4Tv/rYz9KiHGA08NKrbda8oFuUbI8Y3Zxz3WKO59Q4jspdV6LoDOk8Hp1S+AICdjuM2llQr7ou7
589Cw4hg5riLyOX4XfYqMP7Rs+IDB8kElh1wcVEyYqpquWVGAGs3rCnAecFDmqHsakf7IIp+xwGf
wNOW2xC8G0dLgQApVnhebldQf8VzS4T20L6otWNjwxM7+Vfnzl26oslBjxzFGjySuLLwnghxkpIo
s9PI1563flLGpi41aLaDzmxkxIz1yUre7Ev6D524KagsdycYIKdS4Sc1a9/+EgmLMTGHexXkbt5Q
zIrI/xfkFuQjpAb4bKKXjATBK7mc8WwAB+8TCV00S6JvCMxWk290WL3IogbdDrjLAsZHpZwL10tv
kr7FXZneo8+mlhlh8NGGuhr8SQYFFxbo6ouBgUn7XdXWHYvBxM6HJhhHtpXZdvgDA/br6BF7r7Ds
cl9QiJuc+a16o4g4iv2UCidp1/dDJbQfDF8zCbs3PeAk2A+/ht595eHB7NGwp8lb7FQkwKJf0o+F
WQNJKmZPfJ9oizy18dCC/rwl7GERgbtwfoyKJ/LdV9c5B4YiUYb3CUMPCXfnQMG4IAJavFJLyupf
6atJ5ApnTIkhJ8TmxjSIE/HzB9sVgr/4DFfoUvoZkmyGAih3RVCtI9a3+Ds6lcgOt29gftDFPwWi
f55FbGJZncZSQLXKYtmcsAfQMi2wkDtMNbzWql4Qel9Lo1qrrMI1w0KgpUgseq7OcteF1GKEFwuG
eQ2hGXHXYoJIREE2VrNpGTP25YD1nH3cKNKOB6q2tDaNgyfddoYPRhKAJR834luaPD1zxsH8UXL+
Gg9Mu2Ce33rk+rSmqYigghmmcCi4jARAvdUO4w6UiI2Ih0fBHc8QiLV3TDCW2mrnRpua1jG+t7+t
4hX4ONF/SbxdWP8ytCPa0VsAsnf5KcUvZi57JmXm+CaMBQ0Zql+jZaOZYh8c7pBt8ml0JS/k8iP7
ehMISUMhf+GrgMgb3b+PmU7QBOQ1EIHRdxHeZPdM9MBPJFRmoFghEOpFIgHdmySyxmdxkJ6rnfDJ
+g5Fjf7+d+wOi6SRKOMhzWFqhx6DoaAdYjkAtqt9Hg1GWNn319Q/wIIpaPPjxBjixEQmJSE5llsd
ifgyz1UgSdlCfouA5nugQNTwUioz7RB9/svLH3kLUYn+xg8gzwXaKfZXB234E1nC5v0VQBZL6NN2
CWpzPlu3Ih8hs6AJBZDzeKJ9Cf4S74ac2iPY0L4CNRyhlLK35kvB320Oj4504hlv//dXlK49iiS4
Vflmlhzf0eMKgKxE/7O1cQJ6hRki09v7ZGXCjOZew9+Xw4fGBkLAVM1uutANF9Ptvq0MdMWx9UYs
6O2K0N1yLrEDJFsfnxR/liQGywEplu79nBKx9Pbn5jj0fWw5fsabR3k2LpOKi9KfihSr8bsFvb/Y
Jg4QYTL2SHgEp3UZFmH/HCg1aypp7zdY8n1Dl1jc1H9bsDQUOGWLXvMdTezT2Rksfya211QwmrOe
1C+KxEFWdeVM95S+wcroRa8bKW7oU8G+JzcgsbfHAwpIfaQWkU0/wc9NT2gZCLCJnfc5FtPTLdAk
7HVMb8g37Py3oZhAhR3/X+T+jyjrfigNeS0jyPIdHAsxKloBvVukj9v3AbtCpaHjOHRVDJ+DN6IB
I/d92EXXur9Jlrqa9wLBM76QYQDM1JueMWX71Qa7nQjhumo4AlRUL9KsgJLxSa7uCe+Epy7Jo2xO
PSnaZzX+nBlXgMl7PtD6eEpYcjbOd3EO+9oDCE3ozvn+xyetsUBdGoxb1xl37vG2n1kYJblj2Cle
dyMYmUdJmzCaPOlm0eEPcrb4SojaCaFsGDfdMbkmTVZmB1z72hUx7s2b6IbBz72MtnO8izsR81G7
0iKCygcGPWLiyzvOZnNzm2NaqhsbGuNVFJYWmKUlUIj+aKq7GIGaEcZIG7E04rufvf37kjmEFRtP
vkq0uapl9MJFEfLSdZkyJ8C8jh5F3lrscJ5N0VA1tOzu4D78XNUA+9ztSWmDmGAdj1fAlT3/BKDo
i/6nIE4YaM+fiIW/OhMAjKbQ7bT+kI4A0ZIVR0bTI25/VdkIGmbQjozY2uWcwPWut68/GX7KbH9g
cCilsse9lhcX4iTONy9NG/7LZ6yVfe9zwuQnHAG4hRd8vpEP3lwTBSeb8SO3wckrZFnDLEL8WT/Z
ZFBk9gqz/5pOj600w0Z6sKV4QJmxcdsU+YrxLEdCES1tq9GqyEp/dhMw7XveWF6szHwchAPTucJS
1q0gWKyC50k0i1vuJE9YmcGDFDo42I+XvadNxzntgOWr84zPZ6nHGrJd9uJOL46ycAnIMSasKzQu
RWHaBYPPgi2bfrGVinb+BOyzNNya4GMVU548kmCb3gJUqwXMvUkmmEkptzI6phpL35OYbAZU8EXd
GXBUs/lndL29orchXZxwxx7QUaCBL4ptJn/6Rxv4iRRfemINPyQpEFsqDY/Nli2tn1piHAjfcMoE
o9RBtVmRWACrUIXY2whi8XUd2FmuEyBiSy7V4DTMQ2jpI/7nWy1VB51XtvZilfzCiRg5nvM0Kys2
iIe+r5p29SuFMxuGJH5ioRgv1Rgyb+V/IlBzo5jzX2IZHtEP1CLB10bELYk+vZP911DmWQiTHVYk
kuQLDstZePVR7YT6nBgh6GLab7k9EwYyk1GIA/bHhWdD/EbrMY5QO3PQP88SlXxXcA8I+jrp3fRq
z4e9DbOmPfdFnP9yPqwLOiZE+9UOV+ighz7hcjK+6P0n0hiEbUFwQGKOL4VJQczIezrP2rNtLrd1
wPl2pMVCEDjgLJCI/NzUqNkXf1etb7kMnoD6ILjKNVVm3+cA3kk2AEgNH7IjAlSd8SXq5Qcy28BH
+cYEJQX2MJzDbAgmPYLRxHh50Qt4NrT1yjpP2n7rbHUieUzT9ggfDlne0JeRZ2ANUQ3VXsa1iRpO
zvy/G1xl/5EHb+zUlgX+1NsxlKL2V3zXSDvE28UKnWie+yWbcOBXEMSXk+9W3EIiG9qavDUXpHpW
KVm9Xlu3DQXkt4+C37CXx83J0WKxfI8FYLKWdyOoMDc3LueFdiKRMYVZ9lghekAyHOCVufuW884U
VN9+kefZTwmLPdgPMab1/uP4WCAWRS0XJyeY1Xj6+MWoPCL6lhAoVcaHTKTvHXsrDHcwOKGpHT/q
i7sGSazOFZ0l+O2fCzZAtR5x34LYQSwAgRXMdEuiCagjQzd1fh8iJF9kgFXAEh5TcrmAMkEvRu5e
HVlXL4mL5+MstDwo2dXIphdjmOliAze710i3Ij/tB90/k5xvHucKGTpP38ZioLyHQPFe7oqWnFbZ
YxUQxIuRyCRJVqqXnQBn9PMpEZePHGfviVguO4npdvxHPo1WBSfOSRNZJjm0cTZfGUcwuB15oGwn
3hVER/em0m4kWJWH2keKrXb+A+/znnafEuvypaTQMuUwgHBGuZVF21EKnuv5829Kz39B293uutBK
iAinfJneKcpzNLvBrNLP+Jm2ua2MhdFmH3xN+F9vJN9pfS5GeyyMdajw2K37CtCEmgIgWgpxNODl
Zkz7JV6eaWETduOeN5MSi2fGXFsuVurjlI4U1hRECjzzBVQO/F49/aXbQ9WbfJN10kBDcvsf4/ku
iPwmkIgwbVFZVOaaFd7Y9M6CQWfP3o6BF8u5M3chOoAsaeBmx20jJSjUqVE32c//0W/V7+i4i9aG
yh9fY8LGUdkJchQkpBE9hWLwZHlGxEbSYn2ExGdvbDj7ttZj/JNmzTZ7/i2fSrb8jiCTEFHQ4GOp
T/mHBswrsDjlD1SdiRbxrWfJKxhBwBoY1Nym/oqM9w8mv7mCfc3PnOh95yiKITsgivM+2eGPFbDI
rzLVIkM67C2zQan4sq0wlG+5HS4uyGBtnWEjTwxbfRpQpaDm8/NblVOiEi4GfyIuH4yVCmsaQm6B
hhbFlkeqdfBnI1cgf6B+ZkH8aW72EFgrRb/B5UIn3PD86cuXmPP554lIn1Ztd+VQXLOtBcbKZJpD
45Uz839GVx0oi1tOMhpr2MxBOrtizldiK7vRnX6lWEZnCC8PLVYBKjD+iMUc1BrZ4SEOKmkfMJR5
A4WhN+ednaQFLJKRkz7Gkt7d3hd/e9RprjJtQqqvzwJcCyfs8qEu8+ZkEXVgEJJVqSh0DbwNKjQI
mPGUIYpOwJ7+jG+oNsdfvDhgGYTaxs4Z14jabJqAbqtkNSlBFuGOFll8k/fsyTxxlV9sahINntwp
epgIGKTeMS3aia6FHKpS+9I5bnnriLjMo52t8Af459hvhlUm2S3VMrebk0bdd2Xt5SQd/PI8J6ru
Bh2ndOvFTFv3fRb7U601yyAGUylODL+gTEkXRh+kB5H4scd/0t1hpAZUulsNf4vd6vdYw8PWWJQ0
wA2XT3zBgIcdFP6HQADIQdQ8jFhvrovmwNsH5PDmYWEhOHUWc+GTrEgZp5ps1L2dSvE6yv4MY9zy
Bv+5k9akoWRVUzTA4W9PJND6L1v9ieM4BGMBb5Kz7H/BH3jUJ7eaOdxd1xeetf7mhNxfYRxIX7m+
frv4yz8ImUhYF37jzvyo81n62x4TWy8QG7DXty7fcr7Cl5jKKmhzpYByTs84c+pwNpE83aKef+oO
KeGPzorOg82itvbp2P3ADpj+EvQcjhAhqZ8pf3tI0UWwCWJaiLmHhrlcjyupwjyiFm9tqBbmCiv2
BicJVJEqN9FdDTAUUr/YCeboccbtv3Bc++1C7hC1usXqGR2j447CucQ43y7Ma8/43Cw2DKDNysyb
X70vaS7rf6V1mgoA9vl8BtN0HJvbwQSkO1cazI/h9yiih/dkcBAjq+OmA/Zu6ENd0ZD8Zj66aeGW
nwX6ixx5KrzzA59A+diAaeJJgzw4SVw2tmuYnek/vAFxf3SVoi/jRBxU/M3hR5UMkhicLsa8YLN5
/YPoYO6/ABG6rdnVWkB2c7qDlsMAmyjh5IEexs59n/Dx+tO+6X9hyLXPmIfZ0kIXZfxlvggG65qU
rfO7bQcUXcuB5KhQ1N+84UqRQfKQTshL22BP3ms/oNEd0x49Grwyiz0mLJ8JXK0ApqrFdNpx9sgF
JgyT1Hh02N9P7fMbWuU+s3IvrXrYdKjCqxeZDprgOOvwyO2oH1TpAiqQgu1pTWxecUyB/uuMWT5S
0pUrox/YDUvm9IWcQCjTf3ARBA+c8skNvMRuuRMpTtnKM3HaW6B8IkXZqbhJih07mJzEvGwKyCgD
8Bk8p5N2VtG0g4HASN7EmWJxRy46qSVzRzsosBsDGvdLfQgysIkAAZrB4b/b/CuLJwzEiJ6MbAYk
iixcBufcmPM4LRERbRi7O0XplFp7mEUTrqPNeRVuoAUylYBUi8k220qcaFahtqdV8UJIy1y3m57t
QtOSF9RXVS42vQbqw2iEJpsSuvx9h/tLXTV4h3EN1QRc1FnzTZICEBrFjBVjNrLrnxKaFJ6sRrl7
WUSV1xLHWfIzx/0rODiw1l3pj8YZTH7upZS8BoPEsQFJIUrzHXuRIt0BfeMz1ggk33qUlN8b473b
FZEE9UsO9Ezbc7KlPGQD/9QCZuTs6uySI9E0PFTCmZmaAmIq7lMx1hzsRyeKuGgHrWQpzdki4/cu
AlOZLGjbLlHQcl3VafBuFy8LMnPJgntuJUSjLc/o4ipm5KR130F4+/YQXRXKNenxeMW3o+uDa6qB
lQX8wsslFIR1AC/99HKt4h8aVFGAzB+UnUBN4WSPGtpWdvJtyN1kgXjfFJ75gQ9slHIbW4Nx0woR
WpTPm11/vYBJt2KwAIeHMbrbxmDUmrBS2ItBHO06xnlbWztCcu+PmAi8JXRNNyZkxQj8mkNPZBsB
UKLkVokneaifsMEFhLvazuQKS8JAsM1YUu37uECZSQQ7igmN9jZzxzw3euO/sTP6A6F8VnY2BG/s
ezdH7nikHGKSZZyahQR0Dfd2Vw6RfyEr4bX+ibVj1HlRqV8A6zB6fJ7aNdnr1ItKiKGQBaR4xZOQ
GDSd/+4Dt9egNYht/u1713M6aTEWj8StbDPmS01BqakgPCC/nyVkrhNVrAXECvYLoQRABbQOVSrx
3O7m8OxixUHOZ68HpwjZ5G1DxKmgBidgi69dRouqLg0NJwLNVsn0SGDr6ogPd2u4cQYxI8oAghvk
XDSi5nmkS/LAlAE5kXqokaJLhTtfgT02xOVYEe7XL7+VoTUo1SHgBQTdttnTehkuPfAM3UfQF/Jv
YHZlWJXF2rg2meTYJl3R6iN97el+Xf/hRCofsIrPZ9cRbgdJ4tCt4pJfCHiZ1kVG0bhMiH1kUlHq
xgbjihZ+Y+pS5xrbzQRFbgIvB2vVnSWu5ewC20qCa/pA+7cuJM7Nf+nfbFVCtu7Spt+5+iw7gce4
kbT5GjB56VOU2ksS+GV+0OO4DsgH7DWPcC3s/SYMUk9X+3F6AjYCxYUlttSxN5JNuwMqPx+U9w58
s+AlmnNToAEEmchWhmRqnuAjMi2GgfIXnGKnZyKnL0l1fDrpV7dA+jqnbcmpESbGtFRcphf7RVxr
TdTrD9B6zqKedTLR7pSkNsny5dpaZXiKxspSlVc6U5h29m+MM2LZJzRhXnZO8/rGCY7jzoYwAz5D
NOSF01M2h1E3O4rZKhqYKQGMPjGjj3h7laEPRUIrn9xk3LHbNMIUV2lRhiIfV0Kl/a1kVGkDMscK
6/ga7HwjTCP2sfFSz14trTfXwj/KJvNATg1LibljqtAVQpZoz8bh7ANnfuOPdLbFZ2VLOav2FTr8
iv/8tjQy3j2raH9qqXIwlg090BIyvGndrClF5loQr4gS6nWjwLTdrGwud+qu/g2BPXzmws4A1VVw
pvNhvdVSBihE62KY84qVQ7yxs8yGW3HayaUa5bmJmzhl3k34L3o6eC8wNINm9ZoG8oPPRLs/PlRG
Y3SRSHexABLt0mKzt9kCm2sgn8X0VxScy+f1woPXu78ysJZ8Qw0dq8JzOEk1Jv9dcFgNrigT1+7Y
nlb+Ncy2jvTMlajCpcXybwsiBy7LBymQTJR7ttE4K5uwFHYf1rb4XTaNmVwMk8UtSWwzaK+vU7qx
qOShsSdYmD2+ncw2V6UnU1RLhq7oO5w1WD2gBRAvilEjcebmcG5BRrN+fppgzIc6c2WRwkYqButE
+kkAYpvDHBB6s3V4TTyksRAEgQ7lNZJy6d0esg78Xy+19hLRX05QOVzMm/8bHjowg5lHYX2LHmVX
C54ZIPGyD2rmIMp9YtJeDJ8WYEKU4XwFutBGZyo2hi19kOFzfu+4sEo0pSAWycHsThJWC+MJCXKZ
Y/FN+IR2TeH1ORJBVY2nSfjiFtIlO+9Ph+HTU+WWZs4g7OygvJOa5EtUD+KyFrP6y56dJ7rjg5B9
Fw6QAxX9EQ/8QYEdrl3mFEqch5lpoLDfikdversAs0ZDKkh7TR0ZqPEdOpxitrHB00r0YF3VqgZl
4UNzY/FA4chZ4DgTB12pS+uTUMfGiaqfELEYRS4yTlhyjiBn+FZMMLHxB/11yLEk6RgBXD8SXRZ4
ZE7fu7IEOQ6FDUcAupp9IdM7FBluB7QzhrZJdLMZPHx4a/AdDZKSzeKTycCKO1vQi2g0iOm8ZvLj
D/SJQNe6p8wc10rY6Cd0pDUqbSanT3YSgNqQCi//lpWikCBUu55TRsYy8cBBCK+ppX8qlaCb1rIN
V8QYBnEpePGlyFoOYBP85ofHNsAJn4hdzhwj61VR4I956pJmWrRfwT/toS2gs/ryUXcnSE7FHqPG
Xr9mmxD/GJmN9IWFis9vUveJLgWvJx5JYsm+LZmxIjbB6m0NYZ8bDPZN7VUvPKqvCAVrynRJhaui
0MhL+D/PZMVT5TXR9mvTRvEDlM6BorAsgL3990+wXeadd9jQUZh6eFuvp28z4wl2Q+YGe604fTQe
XMB3sL0AkCshX225SQSR9o7x7MQcBbTSximP46T09jMuErQBunBVJmF+YwqG9V/2ViYyPTbYUnTV
kG90PkOrOor63ZZEbtDxaH9DXmr6imlsHHm8yOlhvpM7J5C6LQTJGdGef4CfScipZGjFTtK6yl6H
9TrJo8b+AlDbinbAj40mnlG2kDQn4deMH8LsM82tsJ/4hQJk3LVextlFjAJ1AXKmmhW5UCeqacPR
Wc9x7vkb/t1j5yv2ZAtDxJdLsO3d4ynjV1CmcK+vdcQ8A52IgXsQFi/R/p6wkO/al3WkMbyDML3W
mFgtU0O/ZAbRgKO8ieG+oE3efTWKOCN0oGGsUTKz+04FBfusS+esHCvR92ja618nwPWdMx7Ps5tL
dPZemaG2BVEo8fmE1o2XQf3fAffAUp9y3XpnDMQeoLbEGb9To8oraawk4wLGTr/N5ItR5F8tI+tt
lbdq15h+92KqqU4Lf/n7shNcm8omr5+gCzscliTc1ivUTNIEglJbE4POg7jSIw9y5b/47J+aKRfi
5/IlAek7+jEhtBfu5gaohiPPbr3yGUdnsS+zJ3ODopSG3AjprC3IyCfvduKzqLjkeZlPkb6OqFdY
hJrMzhTQFY7c+BM2dX6sCEXTKYu1T21vv40IOOyBtfiNDf6kb/GailvBKJzw6nsr+lBO1OTRmQPl
KSqJsF1Vvz+iPYo5aGUwH7qi36/sZ6leOy5kA1oWvKalVViee8qOJRsHZmGCAqY051rQPBkchLDI
EKYUkUl3Q0y95AArIHmzOhoTjF7F/R0Mv3hLwyiw7Alb9DfkkAqVG7iq4qRKXo6aGdWbD/vOfOSq
GY5RgIWbr1S19iY/F4+v0fU0pq/wHgdkg3nlTJ8kmYORujuah7bIBn/JpUVjIAgDi80vcEsccebb
18547xdgyCRJIEvHKjT4xCxkCk6CatD0cEPcqM5aGJAYymqytksuiqmB4jr1CEuklObiZP7T7Ds0
dPmwGfU1gPPfVfggTPXRUpeiCvNh4Gt098drISF8rLZMilCApnyHTDALG6/d6AukEZ+DCFhU+Ai/
dhcTnbjyQqwvVPqgZUyJ+FioII6XpTkQ3q2lH5kZENemZUxBV4JLxivh6Y2kYO4PKYrF8dk1rr+7
95lqrSGmzNyuKiTiOwwoesfSGsIifhcIoXZ1DuIOhTmNrXUawiAmj7yqpZNDWAOm9BcFlGqOqLW2
j+akUIT/7kLiXeddnyuh6+opw/jm1Yi3z/4mO9vkNCRA+zOMd6H8euHksgcD1FqSeJbI7KRX2ksu
RnaAvQN22ISSo85AuXirbLgGPLCrNtAY2xqi72MJv8CuHOSU9gwYajXtvtg7+s4pY+6f692OIEca
8+EvejqR3s1U8cbmiMT2C7X7SbMGxSl0hV0/41e2Xei3BLE4r1j6V6AghzQTsqo5BJAZ6HVOSsQF
hvMmpALG4pibobj2PGasJbInGSuca3jefB4+RdJm1F3sJk3jWXECU5Z0wGFuM2lYju3wYGPZxAB3
ArIQ82ykmx6sEzxb2wOeTTbLmicQFcBJ7SawOzWaau2xIl6CFktBNSxqXdjywSbyk6xFl00O7j2f
XNtEO52YWqCDdsIoLB4A/LDKg2kPlGtYkvFmV1+UflzojTVmyS5yAy9cLlESUqxBan0susxvVK75
keon6vcxTy0KAi2KhL6/x1SwH4RzWxdm1PAGGFkBu3G+aRQlMkqwIryP7KwsCkBn8tcpUUTDh1HO
frjKPZpthgwD6NxjF6mrOkHgBwpEUftbgzSgeCM2aE5PqEY5bj00qblQYQ2q7UWv8Muj4M4jLFu1
h3PRFkUhQtwKBZ0O+JzUMd/AD2mZrzBDj+26bSdt3MDndwxEUMPsb2YRCft/7oOz60YNM2RyIAK0
qtPzI3k+oNnpuUgk5bb3O4PxLN8e+7hZ2r1u41l3caMrucpykLJItm7JS5CEWbnAhXYcDftHFGYK
Olujo9XSfKcf8FrZM84LnHVYN7uxkKxYdtVGmLSudcuLRsbx3v3XMXHAWnvWghxgbBhe+PSNTzW4
3OAtwQjyt6m+/YHLKZ0/KIbhYA5po3/K76vVvOSSYePK8sVlYHJxF3kxp/9Nh1SXn4d44wfeLLj2
ezeWKH+lFUzSTCrfyr9PkD/MFeYWSoYLwG+lVLsrWHiNTERAtbv5/j0r71WbM0wFyNa2lXGdRsG6
qQm6dM7HTvaG0AzJwKx7c/F3k13Ghy/ayJsmS7L0jafcyneMmo1X8Bt9/XC1sugqBZsbip3Aq2ws
08THorx+OsC/V/xWbVMJsu8ZhiC/B6VYlYIvjdY0DgiCZLYb5b+m1VdYtu9fe1ZqDQN6IYxu7MmS
GnB2q7KBRnlRryCSjszd1GDUGqRMoTRQuETRmJ2fobeOqNdXRvYbNO24Fom9tNSGm3qzJc/uB1pC
RlYr1qg5VNUYTU1TqD5NYHNGtB1XPLV7T02NjUbuLendYu4kJ6PegZANoYfbnZ+xT9r4wt2wkISD
p2NNc6exuhkcbO4lULHNwYTSdpeWWAoYApQsH+5Nrw7RVpe34Gf8s612uPblAHNO9wR815UhtV6j
e3njcZwCU3m/49mpUQXjXkv3jJfO+gacSF6WV/XIdjnfQkRM7KDgyZMTplidNqMFhudiq4XGf/j8
nz/2MEE3nshP0rjlYRlRPNy6wea8aP7+ypkworUI45t2JL3bPmyk2yl6w33PSmcosrliryEpE1JN
DS+D0JqkKc2J273HKzUbUozXKGV9xXeUTjYieb/V72vzoTHe4vBK7cEvo6hEVjyBzeFc7P6eKK6V
a2c2mFvSE0EnUqYnQF3oaGynBhyzI3SkDnWEZOcmlQWF0yMY68/HkwUp+egaauwDjNYoVXTyKPEf
FE0TNAWBO4Lz/sDyFTjKtMCS1le+xnKW+YHKEdRoI2cB1dxnydeF4/scFmgPPHhxjdjnjgBqxpzJ
w7XJwwUSZjmar54CECr3o2bj8yKwdf6D+pjStaqhYm7LQdDv5pu0UXFdOr/KdenagdrklAIN1tho
OZn2FwAJ7GR45C3GTMKGtJJrBaAa4pgsZ0rkveCx/nv4H6IMxxs1HoSLYa+pwhwdTS4owsolPNvp
+zjoBp5HvJ/fbA/HDH7Qfo+G/kETGoe+SmImMdVzwtTrbi/bhJyTrLQ5r1AP69nbyeikfCyBNePL
cdzgto3wpgcQZymdQLOpDxjw+Vsc08ZMSwV5SBPA5yiSVrTASxwI7Zw7Ig5QkTpJ/wpztt3XSEpH
Vnl8Fiwkt2N4bVHIPT0qUBV+GqoOTaii07ask5P0JbOjq/IazXD9CVvN1sPYNkD+NfoWj/5LqH6X
4JFdzKeWQ9rdiNEv80Q+kmeRp8j1HVIGdXgcELsqZctB+0PWXeJ+1rQgCypSNV9SyjlX+HDezjlw
Wbu8GiAQMJxmenbpxPuslNIYU4PUMvc9qTiFqFsT7t3VU9d/5Lc2xuaqMBRDIuHCvykxdScHccSl
0Q42/ZV8+/LPGCceMWVAUyT7BfVsHWOgDv7lj9a4rgvNS0zhio8R/YumG/4mHqKjXdKmWNRlOy71
i5x2ESkO9RRMG7eCu1DeTEPbWFEFb58KsLqF0NBUU0r8VnRwmo+/NwXWRWQUfw8mX7TlcKNl1fWu
vZXagg72CjkvMWIOxm6dgxfyCShw3iQsQ/sQA3onB2VFiVQZ+u9xnphWN6o8cC9AG7/yNfcuuPnb
4tqLM6apV1v9uKcpAC2uVkTXpCr2EVF2ZE1LfOw0cwP/OJgEtz63nLa/zT82+YZd5c54jrXQ+GpQ
fuwhGSy277XtsLyGEwac+6x7ugAI3kpbUesEtOiRVlQdrN6HdfTW/viwOKJoUahsx3ppKXEeo45D
UTQYVmyNh0PaRvdzBOB//VuKe4eKjCXX3MXyPtLskVCIU7UZUrEpJ1QrEYaZospDRUNix/SioUTM
5PSg18ncCKITHlTq+bXFEXTpepgowvJ1jBZKmEcFsa7L5NkuxwcrcMb6KN8RMnXrfpIB+auAeg+o
o9CXkkcQQlst9VhhEF3ZicW750ECIFYW15t5CqBjxpilLf95wU4/4TLnClNctszln6AKeFillh9H
GaJUv56IouzKG+HrKYLevkLu3PIyIE/BJQyBwgbRmzhIFVb0YE2FjQH8eaI3GfMJEHaUe2+mY2OE
VTE5zcnWrPb4RAMBJTu3oKmGiZ/HrO7c1jtUX6aWBIE7YoPxOvbbmIvvFqpXKU0MT7nZgJ1fSoLU
X9TYgK3Zvc8evniLFYy5k7as62l7QK97BENEXM4GbiyBOQ56OkRrzdY+0jomVonAvGaeAV054Jgc
5AlFgKQQREjdiuDXmiCgZwF5XZZP+dzxgrBpVwHR77lCjt29rqGJ2BoWIhnOeylzGdW0EZSQ6rfm
jcPcIveSoaIfXQ9KkpCPCxSmQZE5V6sADa8DZFG8zbeSZNZ4NlxQhxjVa1vxNv6LzASbxMjukhfF
tH4kPvHXWY6rJPbz24VdUSzCLTSZWnrEL02wa14maZf+whM3o1vXRgipBsizrr0T22duR/nIxz1d
EDgsysrBCL6OF+PTus9L/AkHEfByRMiaXRuXp0RuR0zVhHxi4lv4CyG117niHYUZ+Boc9cuGoEOO
rCVAeatobQymDWA75oD4gc0gB3daq5OMKcQUXxraaxJV6lUXeB6uvvTdUpgZ1Rt8/iOVGGuxAeM4
oNCNvyQhHY2fTk9WEenaoLdCJAwJGh+PqN+c/h026DtqB0/hXM82YXX+Ky7ywS1j/FMndbEYFsdG
wjSDyLN6s2ui/lEHYiusjG3j3UwrhJm5Qtib+khRzYb6Jgh84soNn0x3r5IO9Hn7Ck8xgujImy/U
8U5tUgOzurWxSnaA85R6zycl6cNDRQ4+mKmvoIoMw9QftlqT6qhewXa6rNIt5RiuGW/8WHSSVIun
V+r8/Wd9Hbq0AHKEZij0F1EPMl6NeMQmas8CiG9BgMjdNVOac/WKvZcehqzxHzFJBW1JaVOB9GAZ
4TN3WzpfS1/0wZ6kDpvzecsroqA0UTwZF12FKtm5OcuIWGaR8Y8KfJ0hHFUOSn/6HUVgzH3V3gmz
Leka9FlM26Hyhd8jHISnwPXRQ1aMBCgB4Dt+g37jPQyIs5TfPFnNhJHsr97Vux0/nU4euyCUu3Sp
JcyXMl6rFb7IUwXoBNWMfk8oE+xOz/FFTkrhPjDXej7hlZgr6N9qcRiuHMuT+ai+Zdxr23luBm9o
eJTs6lSENNYAVMcQKPx+2atsQzfffNnE8SY+FWRLVAPztGAcItG3LVPY/8lRKT6QhlmYfPSNEbOG
tytjCf38lCzDzKDYvf0PpEV/CYWwT+emGMUHX3MH5eJ3w2EE+jRv/jM49z4gsFyYWDMGcKGRS8Ah
s+kpA5PX4xntsATVpCIQ9JxuZDpjjHbmIhjebHx27NnQqiXCzu13C3J4EQQvdxhsl4dsvFgUv/fU
pS0+qdIdP6Cg7kXjOt3oZXqBMa2Lhxx+Qbni8HBknvvnxnQGWi007MypP0W79HCaECDUukvqRsSx
gGHh3KjG+ujmqRtPNiinjq3yVrgQstpYJLwrChd4iGZPGmD69SAx7WAy+r6I5pUDBb+qK3ZWPcFl
Q6VpVyJvI00CqZfel0N9kw5d8G7DKXEGecIaZCu4jOBO72M3lW9mNXLH7mLL5fVazhGmN1H/7vWD
kJLp2vszrRZJwTRdaK1Z2CxWbzct2DcWYClZYT5X/PgPRWCiCmAxUfKktJuo++DrIS8yukVUee2e
Wmq4uKzTQpTzlphdnFxqU3Egm5zMYw4pVHqxXk9eZJayk/dNgiGvea8vYOfk1DmFKxbdfvGkBePw
3Oo5AojDjH2X2E+LbyK4E3stnyYb4GM7mhgqn+PIPLWlATwmVUkc6dT97DtudaT2C1q/ywgAsOA4
fYVKgeq3qStdEI804V5V7UkwqsslsrGLtBp7LMO00WkCi5E58icwtqeamibjcYQ0QuftObM3ICvw
PXG+5mi3EayOV1KjzPSp/jGawmF5p+boY3nTn5774N/3E5b99iIF9GlVL7KGHcp5JjLgMHUUZphB
L4iDODqtEoFs6MPUH5lCpTY12ZXPTQsPfM/OPwEVCLeYtG1aPO2KWbcZ64epDkXRMqDrbUmw5MFY
/vQB1Q/RLbzJNuF1V36CeOlFeHZmJ1mKhpxlE0PFidkFku5kpPY859QxhusKXolJjMjUGrmuhqAw
AaWxOmSKndxdE3mkla+t5ruC2p8/xOlc/XwpZJ9PkwFdI0SxdOplncm5Bn5vWwkLqwyxpo92imNi
IplEbYy7Swk5ETSHGbKfUjZoSfwz6hVeaZLgckJT7SvEhzysmTS3tUmoytkESnWrmT95KWI15yII
VOmlQ9ADqEEDT+Z5oyezmtiJb+p+L3TkvkliYZyXkV2gXpqmcM/YA7vmH/K9X7uDqfvH0MqM+Inn
6+s+LQ5S9oAI71eF8YKx7vcK4E35HFSBiXFYdkXpfjhdpUBoq6RF0O+BtcR5kC12pwK3Q+mcXWCU
AzqAY62WI64Hq5ZKY4z9ALTfCOkWSEx9m2TSgFnuR6ONJ1A1CCna5/RSkkUQYxl6LnGchdN8sgrk
Un+QiSSvs7M2oXpNwxD4/S4MpNjlYCPESh56rl8amziJH2A03/rEgQpgE7pX5SH9KGYe36udCaaq
i7nM/BfDIUlTtZvOrUIxhWWohsVimDQnrC6w8swxUvw3XtXzAGcWgtpuNQyo/WGeP59QaNd2pWDS
PZBulgs8wpFR5iW6gSr/Lce7Mt7u+tc6AM4/qIz6i4Mi/HtfM7zCVGBeeLWaTUg/G+OvoOvSwven
GcSR7kJrT94gFn+oLH9ou/b/FyuyhvO+gRogz1tyhLQ5/i9Zw81vcEei0zsU09bqLGW+nrPJgGOj
MHvwlyyojdqgikZn55OV7ChYrxeMWEYTlSEqr2BAgkcnHocrtMsH1Xqr7S6vLvA3CSWUfMMNTYYZ
5sL7c+uST1Lx4qnoEbnQaHxhrI23yCuKL+HGXlLAhDDC0OdNMudSs/zqZqHcxK36NNxCLCU+v7Oa
xaL/oASGXmxJ3ZkLabDov7/U3lY9QmzjRuT6LgmytEfFW2J+ZHTsGEgH7e8G9ei58BRw+IeHpqd9
qwAW2GmpgLCdsi6db0xtdcX40TeEZw0p7hrW74mZmQBWWkAsaW/S5fPOI3xcF8UjtMttyagHaYJe
m5JQG1eh1uFjj0LdZZUxGpIASyPAZ+9G6CccypP5608LoPrP4URlkZEMnjiBlgwlyBqvI92fvzeW
FQ40kr+j7fSAaFZYwg12c1MYf+hM+ELDOmBpT05i9X9b/IsUFK8cvj7q8jcbinzHgPDJ27IS+KVb
2JcB9JIHRHE7eSjqxZ4+lfPmM7925h2JoiBBCU9wyprmAFRIRY5C25iGWQ0LzozZn3mogl/BpXgy
/8Zej7+6dqNA/KVk4poUFUuRDLHRdQEm0E0XnRCIkU3eK2gaD5FvIsbjtk75ly6B5YHjOpxIOfvz
MVsgd/yRPmORQr+qYGJW4qWf6fWBzoJ/hP/EbVAblceUAumbP5F8J/LTXzR2JtgrmT23Q4duW4SQ
bNaVfOHv5LhqvbZkLh0z1TrfoabcSjhVdTPTFP8+i5sGwHx0ZySGKq8bSdJ0SsYzPGK3+VBvMHbb
mSlq0l531H33tnlzcFJDlhfJZvcXDd8WvCGh8rUoaZWy5eTlDqewFX9oQ2cXROwvASXRW2RGZjId
rnqBCfJucwgBi5H/vkqzo72JOWcz0GU7+gPoETJ1reiTRzaHhlKwUnY0dGLm2y+cFZgLcP8/z9MG
cHMP/rKvd1SehXkGjQ2vROF4+CRy0eD/zKe/e10aZPRfPdcu13feblFXgHTVFBuIvKiXpKUzeA/v
uOTUXroHLIzgeRbkI14h0MXRfO2vGZ4puS7I/AWfJ5s1CGUgIMMQ2/tMEaX36HtKPXpUWYB0wdld
CKnQUJ9fnp8e9PigYrd8WSV5m1xtTm3oAyOiQ7BRQLNa+N5EtJr1RaqLFX3bbzFF3DVQPq/+ikAo
TZqldj3VdTGr9GSPcpsZvwaMKglCw3aCuRGWD7Zr2jCvGJ9oifZB0NIWoMhFnRh++g8zYt0982x6
YiaRF5vyyGXMH/KZdQDmhwVxOr/0TwdYMu6Z8XnD0TQoPmn217xN5hlUvd65e9axdaHnhX8/TlDD
X8kWHDa489s7+uKFhFXCis1HisPG/Q30UgYm3m7OQhq2+5GxZsP+7mIsiaZXKEAhaz4ztf9c9hjl
IQ6f+4nVinp0nkjJzGQ523yuB0KyZHA61tJ0Vqh4X8uc7lqgSPbVLwrewYFgJ9wuP/rlLwZkfdFo
bhqUAMYAx7/qpQRmlSf8rzX7lVFFlHXrnr7sRyGyyGpuV4f+oaMK3uGl2SgO9l6Lg583/PQ9iRja
mNN+v4ecc+/qYk/d/WeizAhPUSfXQEusuF3Rwd/fWIlRoEHHTuIrnv3QNCdpXac6Fc+so9JhxLbP
y6yeEXY7CoW8n48cqR7LDkONuIt4n/dW6eGff6clnTUK26/U/8pn67AqoydpBW/RTX6h5UF3vQEm
mOG+XXA059Plegsq9TpaYDfRNM82qrcURgl1RrxR2t5UYZxprrYTO6HqMBpgdLebbhetNWHg8sKF
m0MORkBmUMBONqa5dp5EzeQRTskkj4WXYtP4wVU+YfWoI4MZKfIEC5xY3BSAWeWBcXWOcIOmvJsY
KYLXaYnpKWdeQff2DMXRCbYLl8NzzK+d2ZlHZrZTugp7qjQSEAU+ZuFX2u+D+U1PLRUB/b4Qn9bG
jEtDg+w49pm99/4ZQwTLAZSmMXRdnrbkDrxGiOP/Lurg0XyCQRcftSdIgEHCtaHTGtsJMbsFM5CY
aRPujCvhD2sbPMOvDxB/wlQGNAvofkrCOG+ndPzjXpkgdEOuYocah9RL3f4or2K7zDth1QHSJI2j
eEPfaV+1/7V90KddHn5cJRqxUppAHCPiSpH48D57snLBYvzm49dsYCa+5bL7K31Vn+UTTiuvkNIx
GhW1xFpBDRijTNYIptv6XZZbmQzAPBlglt207TVx3Ukv1Ft2RyUCrM53WHqxyK0xAHQBliBm6/wM
/xBZ3FlpNhjFLhKauDr5q68caab+jIJyssbA2SBHesupyHZNAHZD0kTHr4AE8BBg3IYeLIfWraS4
CJfBlwJ0WhkHHITlDPT1wc92qgb+mslKLhQynMJwxs3h/ltbhsjwCLC5mPuVEUHQhNp1tb6Q7qBx
hq4ailWAxzAHc50iUR4jdmdZ1n4UVmTA+OlMhejrK6xty8FwXBCJ7qp8K2wcXG0D20lUzZh49VZN
jUOvzmsuOep6gC42rnDN+Ywy9GD5tAN8/vfzdEJh+Xj42XrvJ97+QFxFQaO635mjYcoVro9q5baW
AaCyEyLNwZPI9SanMA770kWThmWlGq1ezSZHjkj6lPzXkwPIl1mYbtPgC9yePKP9O0C4Q4Ur8jY4
bLmLzGCPewRt+uIyZp4XTXyKbk6HnAFfHfslcTh5ZJBfkOEHIYp9iST4z3mRRdA1Lw9QiCVlI6vQ
QWT+unmsAa3Br1wvWszapg6pkSOZ7sm8PzFxxVoBdnagKCVyLupZhyIS8q81S81ZJB1/hjbDzdcU
mqZF+atnsQLGhwq5AIVaZYF8F4oF+nLqh6nGJPggGa3TafdLALaGDlZg6mvewjMNNLxzbQRoFZ1C
qlf8gDr+NW7WoMN9YUKeTuu8AzqfUwKIzN4nxyDN5rJG+1Xsc0SuyT42v7EiBpBZZUlusrI8aWZ1
et8Csl/zihABDuBlCPjkXjtMPbnqXLhcaMzijWWKgX9cF7FtiW9Su0YWIcDVCfBH1NZooFAu+xuw
AdTm6XtBPx4b0XoN/2Fo382A4jR3Jx6Ux/SrEYrfZsVtEDnxaMI5iLVMJi7ZddtvJOdiBXiMZPgb
226ax1KGx2uXdHbTeToVQkf1RWQVN8c3Hg2GPfXLFl4tsexqo/Wu+i20aQ2PMVSD0KkL5s4HNP6G
nYRHDYwYJ/j6ljhtbih3NBAntG8GcnoHrohEuxxKGE1loVheT9D2NfyBGgYOuayTm5q+zE1q5jJZ
19MULp3X3CWctCcjw99Jxe+SxXM6QV8sOZQkcm/NG/w5JCzfBZsvZBJ5F+mSAOwq/J3pl37jJiA8
NKfNMLQZi5GYgzIQCCo2rNWdGb4SDxnpKErWuEOcNPwVGyoOlK45Dl+6f9LYbGo3NzO1i+wFNNQP
2UtuneaDb5aAlfu7FK+4GY3gnI9Z9qouOHNtJbM9pFVS7Mr8XgYoN7TU1v0spjkXDLxqHcyM1GNw
PVL2tgz1R2YO7jjdXJWJeorluwLhy1xyRedDyAQouEe0evuNNfRcl2t+wnTGoA3K3tRK+RPb5OEv
U0qi88CcIVLWFZXMYN0htXztcpre2+vZFS0Cro6r+LnwY+c/hjMla5plpK+pjzc+C32lsgEUOQ6w
VnFXEgZ8sb09aGDDF5RvSOA/U9WvNd1aCraOcyKfiZbBDSt5wynzjf9FnjB0YagxaJvg0l+ZGFZR
lCjPmCzOrn3VUcfyVNP692qhvKoS1bide9MkezQ9oDdlhozrSa7AaO6CKzHH3MLL4IhMoC5eTTFw
xeu4P0y0Gs4AwrBnMteIw7NHMrKIE7cBOR3tDHx3aJ7Zmkf+mtqjmUH1/RMSxH8akQ0RSa3xEK9z
af9JMwbaU5I/j9CHMj0K1mwaZ4nbzpUD9CRUPXTaCnKNLBZoHTa3hUjdOM4WAi0osXtAuPWwmbyq
fd0aB9iW6OQFPjj27mT3Wi75frVl4jY0YneEfBd9CgyfFjv+xNgEXXL2+CCFxbVp5yK0AfbAzAgm
n2kCDtgGawMYRBJY1/GlIy/92FEA0XHwgPshk+BZhY8nmYfCRNujEYNvgMJG04hNC7w0YToSdfT6
PeKj6xk73e4vfHdMwJsb5m5CJzRogZLsbZ8uUFqdy3rDVFmBXWIU14YlO9tGsTpCZ/IyUxrwoRiI
gL/zhZ/kiGvtme0ygIlQDm8tGeSLqbx6y/94t52Mp8HMCsUudDlnhpCJs1NM0nEJ/G9ZWRQbobCe
fniAeF2Jk1lsy1y4FsNVoLY5o3J16IC/ETE8xTTAkZPll+HowL9Ug3a/8dOXvjrZ9al57KBugsIf
SNB/P0lT+rnE5bjWEOXvVbnHv0+kO678BbzSTtCgPqnoHymC5QkKmk+zyxJEkW9F+NSD9MC6Xu+V
KHYqbt7CnSJazvMdyDQQo40ZloWzMsBXJ3uuoLMyPThqHK3ufuQWnbNPZgkWfAvuZx8Aj1J7ray6
y0AzJ8jhyP0cxiilOXZKxrVOAQZgVV5dDuBFzK19ih0vJiUTqPfEHslzxhKYYujdIktBKoWxM4H4
+y+dn0rnpzNlW5LZo89/m1TCunXdFrVBauXjGPH+I0w21ABsVAaygV7jTFQ5hg9EoLJgZiILUYFf
bpeY9Os9nceggNSyI76IffYXZV12Jm4KbQcUmG11J46qmNbjyPvRcqdfywmtmuGF4pvWtvskReRr
dH/fd/DZ1/sykW7BjKQfzRfU6A4o2qFe+viccIQ3NY0pr3PStUjFhtG1JuPX+QFxyJP8x2ywR4Pb
h+WhyePtbdrPoKVAp2dNbBFwB72pYUud5bfKzCF6a/yyFWRD+q2qF6jru2TeldJCPOsORN9k6CaD
9eRl39QA/ogiOfZrVqHgQpMOAb3TKJ6cMLZimGk8agHpQdfci/Ml98nJRkvw2XSplSFHb5CqDBL0
Ln8+aaO3WVI1NEHqN7tuq4bcA+a2dk8iGc2/956suj4UC959FG10NZHEuf2C/IlJAvpCfeN3VxFy
D9chuIYC4LZvyiVUscXwgxDCjnZlrC+F6a6M3ulkKUEcXo8s+PWcjn4tokJz0jpun7uPTiu/plDN
hI7G1HU/uTAv+nuLtSvxrHRkkJu38XtbfnBGECsx5bYFM4DkzA/bd0wBsICdirjaq1b32tM8lgbV
eWCQ7TWZv1KBDVfzWEvc0VvV+/mvQscMiZuVSAnRgbysNjlLuNMaUrfiY+p0lLV35sETX/FjoMGj
BRsNHAcL+w9dMRXRuihHON41CrDHBNsqgGuLCUITPySz4v2Hc3TJoKWKLqBLwm/MC0C0I+Qg0ROY
giTlvCGqfxPvcGaJVM/0vBYBMnjE78URZrSt31BuTFt3EYKQxcenmLtdql/xakdLWyrHDbvw7ebc
9VKkjxucNpC0ZKckPoshWgyuBh3d6rAqexZ3aep2icKNBsiQLwTwYOhLNfLErSaEQHuxJsexNzyA
9G+ZjGYvHAZWAOjeIYWqqvot87ogRq7UKwx/WGcThHyTa0xyzzwxwhIaOhpgGCNJHb5G5GTgnE5T
WrP30zgee2xOvtO9hVZgLZHRlJ2tVOVTcqGU6plHwR2LXg9MO2Vn3xIud6zH9jC7EAvBSZHffzdN
JG/M3gkSQC4669hrUgGKeNFn/VA2nGf9FBoAdJIFLxwJkDi8QYXoafAj7NxzVKnQMvWhP9O7QR3O
pBaTNVEz80fZlITlCAbuTiU85vQ7q5K6z1LvwyDrGSJ9CitaZnQByOGFZhZ1XlnyAQ+YY0PxGnKe
yVpTcsTXeZrBgOQfXf7h3CvRMSPQupOid8JIudRbbdVVl2KwQVj6TSphHXx+jrKz85idtDwisPGw
8p7D96LGRcC+wr2PAELRyCL0Ryv8Cwb9aCnGbPKwYfXTEPXdG7KoMzG18H45NmzMziUyrMUBTttM
byNbBDjU/cp7RrzPCUD30ln/04zWu92ZAEo5dvVYJDnOXdQR1bC/2eMrBKfx3c2gwChWWVY6GYzP
ErqP56cgh4iz5ip5TDnfokxHF0JQWnqGQBM/lCcDOyAsrqaggkEr96L+yj+X1Pkv0EFTQwimjdUo
moYXbRsrbGafwzvrAnKK59Ur7XOQbUJFFzAs6PKjO6V0br7BaRA1iPLvD9cdDoCT8VVnq3D5u90P
1opR2GGHU55Gq3OyuF5ip2mIkoJ1xTNSGQY/bvcoKMv2PXDgsu33fwAf5Ya7257J9X/puhF5dL9K
d7Gd7TRvRKdK8Tmnb/gTW6YJHKj0jnTl8RnFXoMsnnGTuv9C4Sjgn+PcoluonZf41JL8NbPe5UeR
Rj+lO8DRCmN3Wv7gKUOobZaTBFfYFTx5YaI0yEK7r+/OW8WUFBXF5juYnPUuTkN8B7lGuglswJ1U
qtFK+UO9X4KXAitKNH/IetnPGmHUtfeohwaqsBl2UeKF4KbTy1vzkcDLmXRXSD92p2uD3dSNQb7n
1oW3wKejvs13r7Y6DLy94kOja64PnGgcFnjHs740VLPtC8yvS2OADeEYBrZb0dd/gu65q9kyDvKa
cKWa+y1DourR2SWvavdy3B8izXbu3wwSBcpeqUCUtGFqg7dHBPWvk8W+3fOK8i3diRrfhQkPsK4/
Dh2uFe5izOgPUhdxeQPyUCJ/HEx3QEC2T85+bWBeDA05Vx3v+vxII7rJ/KfHY1bh2v0D8SxEy3WA
1A3MUHfg/HY3VsEkbsudgtP/Z9N8gJaDGfGxvPROFan14UGAWRJkFiH2aMb1c2P7KFduQReQH6qZ
JsQGCVTov39ZYaxNpRKui26qEkW/u46BByLQ5z4NY0VcSLnRaADRDY5PbpNFFp55KAuHZR+/Gb54
S8liF9SCcnnfjq8+CUpYKh7GxlTAAHaBYFzNVvjxnn4vuPC4bUvaF4bobpTSMfL8vdie5ke/OZgp
KguJKqk/8vusiSoMKyxQFwHkOZFTQyS+X7h2jOCJDtwgUid+P4LrUkn6hJlnqnO2xX0lwXeiAvvi
+kSsDQ9uSQugBJzzzGcBEBc5eHZrdDMh6GlZ3JUWgQ4Ax4mSwfaziuYW91HZzUqwaGJaehjD0YqB
btulN70z1PkYJ8Igtw29h4on0oRKMzcI2H6JFRORgi5AlTSTSStOWAd/H+TwPYNAz+NLFT7EQxnC
OmPtuH9kXxR5mI7sBBtELQ2a5M18vuyDNTv36lOrzH/XSIKF2GMQm0ctzhofhy8WpoFaDwQNVXNg
ukJzWv5yGeAHR5D3PZpRq6eWSlzkfuYBs8lFFicWGWJTdq/D+vC4jpsTPT+Y4ORSJ5qA6Oz8ScaU
buq8Q2uss2enCYQLEB9KEMd5M75clXNpPEC9dNDhheoUK7tpgxNvTBmaDB5bVWU/Mzlenwu5Y71C
4OzgOchtFhHLUljvyNhxlBW/BZkAaziGVQcVvkrH4MfE1KuemJMrggnRIqMTUmwPyWvS52Ev+rx1
oW2sHI87ExKRfupsqwYRavQ5eZdbpvAu52aDSEBATs2/HgnaBbzE+3wSi/99ihW92GU0h3j7hmhd
1u+M0nvdH5v6uklkpumsIzEEBHwGE/uhaqd3G9YbeDUzsB2ib0l8syqZEjtUDDNJR0sEDybNgQqp
nX0pHH6bsmhqjg6XEi7hyYwkqUjWApnZOgdBVXg/DGeunNgW7+0pdEBPQXqagWYNt++gzS7qSmSa
ZyXJwHno9+NR2Cp+ZnF+e19O0xpSvf4R5k4OtnusZRgCP2iNjBfNBqtq9vpAURa83FcwMb8YBNFX
AVtAlgwZ9Ifjm6Xjn5DoHXg6/DD3aSaumanIhxvYQU36PHEDT4yRNhvGZ9Jp9YHtDXZ5F5N9GTZi
t13MMSyN07tSr9puxuHtAUKFjgFfZxKElJcVQRGtgzq/VhRyFcpc7etO/vuiZ0bxsWAvwBcFIvfP
+Y5F+/y/bTaCMvdndQyAs3lNiSnqIMeoxLH1zHbNAtgz/XUAXMV5M5uLpwf07Q6nwMeKEwuek83O
Y35vQUio0xzNsJryDZVSYGR63HBfsaposErez8WFOaqYSxQtqbh6PxGTKYXY/1bJu4U66AxVSUkq
eR+w7v9a2fibJXXWlqB+/aTfLF1j47DDKpmynizSNsOfiVvMKGmZfn/lKg5S6MAN9LO0HtysCdZY
5BRGWWJwGBpNK1uL7VGJDrhZ8hOgQI8CLFP2iKDEJyV5y+ZBg/m85EmfN9MroI7IOLmcKzcW63iT
IlN5mnt0v69HcyiqXvWmM7Epl6qJ9EMdGiY2b2KyPj4cT+/fq3vYfv6oW8AKHz6AvBSDygclYl9Z
QsbEMozQwh2UrjML5BsMRiJqfYO8p0DWXyksr5aHp5XPjVLeJ5SlZJFKauPooa0owNYgYm9i1odC
0v1wZZBH3mH02kj2yJ3uf9euAOqhoPGjDFcub2SY4PSErSbbcNsRlfi4hHA501vUBsaTWJTDcqmu
xJ5+N9QDc5FFVF7TM0vbiVwBf/oy8BzcWzyCuErcfTmDMTZ4o2NWk8S1BWHWY9kRza0UilMSnZPa
2E2nOMFh8I2Tw+h+kbnQsicai/15FBbBgX/Y05VrYSEEh3xgup3pVEQNaHeuzGDQX3O2mQivN9k8
3I0RT7QOLBhjTXxXow1lgUlaIDNiZOI6YYT8KnRTDrctDwvoD4bxPrSgDJwPy5ZjGPWViA0hXyrC
7+SDX/DVlb/Xdh7J9Pycupep68TIpbDzSJ1LRjHtz8vmPbHxA5VZUOY1ITk+DUalpIhlqq7cKpEF
SB2vDo7LDWTWiGSnCuBp5Y19llayVm4xprKOmkj78TeFAp4h//hktGOL8TqzFJP9eyNxhyOtgi1e
N4XblmaLcjYKe/39Tp9bbyngdHDc4bmIPGCqtrsFSIsJ3egOgLgjoyg9MUXN0ALPWZzw3pBTIKX2
6Utrar0HEqx+Sqz002Oo7c16T4hIlwCFhKL/IXZX1SgBrW0Pb10mrtvlyyeClgHH7yi0pxjokY7J
500VhoFlpj0vUW8dDU/jnmbbAcUw1oo8gX/3N8/O69LshGQwkp/IVnAf0U9fd3DMstcbSWdcoYAb
8OZfdWNAX3azWrdWd4lNJr3yfnc2TScipoGS06DvVtME8M7dHvfNFyKcP+/kQgQPwZq1B7MEddmc
T8jspFnaPIfGRZpihYmKgyMervHtIgjfKNI5WaKA/keo1hAMc9rcK+PGOI2uKUefHgxZD1C9eMIO
EvIQd+zXdfiCrvJUSuUVU5Sxk6tB6zuvBRHhXiuV2V4mF1xr76D79+C6yB/nDulIgSDajymHCzII
3HbC/+NCAQJGoNkRP+g+38FnzUUqxMD1ymvqlxk0S1Q6zu7/Pm3iUO46Y0OdIFd8CT6Xs1Y4z7Vh
sOTi78y0+DHY+KGI0h1vRxmqPjRjtZCKEC/z33NAQKmK0/5GC/GndLhKm4X5I3BNTluOSalZh8Qv
WhAVf/vFSshH04qUGYDFKaqA18CbN2XdqK1F02Et3/zVoqHEzUYl39bx0ghyoLUeolNHmlYzDqsD
CfknP4kUbo0aa1yIWoJ/iyF0yvWeNjvmYZ7IPJ5r+eh5LKQURM/aFPW5SiZkya4pIpGpWhl7l3kY
HZhDRazt+WRGLArmDAiIRND82UgctHGG+04RVcfhKjYJK7Hdh2cRyVSt8+jCvF788CwOkBL28fCZ
kMMknAnfrOCctSmr0Pe9oyQ+yVgTE9wG9TH5ZkWAARVIb7CtEne2Bf3yTO2kysQ6jjXtajyvIaq8
krMg5Q4x1ipbp63KqIQsVZkVMUARjIKVcfqLm1OPY0uqFtyVZok6Y5E7LdcR04D1udfnLq0VrPzV
MXzmbtBJUqs9VXA52kEQkiLb/waj94TzwHQVoApmTo+ZGbCm/hQyNzU+xwva3CR11gJKq0GFItSV
0Y1TQ/9rgJomUhx3J+y7GXqFsmzoaSoO6VaYsQ+UBs09ibgjcd9cfpOO2sbGmSGD0GJxb8zbj2ux
U2iEv//O15Xb8ZKoukxCbH+Wr3chTve0hDZcZ8YVko/zt4gE2h8LthC4Etsxd4KzbBFuKexxKlHz
ujMyqGdQJLo7cd6ht0Gz84B4HnvcMj8qz1hBoBS63q1qm9XztqfSGzIL+hztqteggTexddbUbJof
Wscuipn6Y2vQ7WLxNSu6RjqLPAcgxwCnOKGZLsahUzrfyGOoMA7SivK88NeN05+RCYJI6WRkRzXE
9d7iF9USqBBd1ycr14aLOPF2kxqJImdo8vFpFQnTcfQMYSaf9yVwz1XGIrsk4NExJgXm3G3teZVQ
+3pQLVR0EpOVTcvnLNv8/6RYO0OUy8n6AvSb+grjQ+7nHCsB90VKNmzVVwIwcUDAZ0Uz4CaZRXO5
8wZqPKKOXh7WA7nRrZG8mA6x+zlS5Yic5rC0dye39CpnpG7qMKTkdvO3jJEt3B0BJbZjH/S2UC/W
CPXN3D7ZiNPBl0/FlrOC1uQdtPf7XU0MEonVAjb/FTf7PufzhAk7CLaDyd3O1LXDOKP4btEA/F8T
hW8l08cVkTJZvXuLe8mNUVI1lBIFoe+MAYRvfH5lgAxhaCNSk/5kHAFLVduoDx/YTE8NemVJ70y4
rstcllqPNXMFQlyTUZUwRVgt5/XHCzosv1BoaExTgc9fudaYfdl+2AEzz49l9dbm37Xf396jVDJJ
h5oU10OkJGnJETAqhjs4uEfC31EBOhaWGJp9DPRBbYaQqKZyaZdBxXTdg91RUy3z10ehw8Z0V59q
GkQEOOwC+bFpnlJ/Kt1n3blBPCXcdJ9o66D6wtPjDyz90xu1ty1NqmAOPqZD3ee7SQ+Q/pDHZQVE
WVF5wJRNBz+OuPJHSSYXKtH4lBV6dfHqkNIdLETjV3OZNcjM2vZS/K6jgKaq4a7TuFBxeyFzDVOS
LMzZnZsIC+8KZ89QhZDYDwZNSExQZTRTfQ+KFPOoPpo9K9O3G5S/FiaGgpxWBhy4xp2xL8TJiGeT
yNBnbzCBot+36WGlHylZt13/1qQxF/jPx6qaAYdLMD/g38w9B1Hg1KCaCGZ4KyOz/fpHJ68CiZv1
jqhqWM7jbmvTjX+3twXFICXnbDJP3B8ylXeXnS3moBc3J6qkGFBcTePtTnrZar+H/S3qKQZmx/xL
l7GHHeqoLB6DE3jVDxDeISlIdkmsLtTI3qXfhxYCcjJD7m6LlODN3QcHHbCwlNYG3YvjjCS+BsBD
vyxpxfXeu3A9R2v9PNyC/j2MyowKO1MBEEAiwOmtlqAq64DXRiQkUi2sye2S3z0kMWswrFquArdn
Oy+mYsWBlD1wyFI998IUOzE+Haa0sn70VizPww7ywjQoEh+MM2IEiS0A/eT7LWoHbblvVGSc7fPN
BtJRqIU9XzK29XnrIfssci+YrbY4rojB8kcf/DbwbDYbnxwApMUcJiHa7YJfm/nKv24xktPHzh6A
mfVaucFP+yZoP0uC71QU2vtl4VTLxxD35PqA/g+2ZxYe5Of95CIQvkmyuShNbf/+piWzJm/sgjcX
4jPaHWFsRwWFPMH91tpWVDBhgjhl5CpDP5D0znyV8Itw24QxQfMgGiSSX+b6OfXquZrlErZJW9S0
8RPJ9RdLuSN6bvp9mOxIarVMvgo9CStPenhExhzYm6BsYcne466GSff7hyTWYVigIG3nA2nkYY7r
WgzBDoY1+6MIEjzQAzLh1JQi4tyeD8LBMeFy+Je9FgWqlp91G41q5qHhW5UZ94QiTdXWAJVcL7cm
GRwbTFBjAr/B+FhFlMQv02vAMSyenLsbRzcU9SjmYawnnq/RwO4D1oeIhqFzsARKjeUxdFDxgQmp
P5L/uS/6X8fnLhb4zvMr7D80RBhjManDpRM+4335tcxt06yHSeJKjcRP86dlpZFIaf4csYkBuix9
8g3nUBAD1y4c7fUAyvweHyQJISDur6dczaZxBRsNzviKINDyVGK0vRuZc9VdQ21QWaecZj9qlf67
o9FZ3KmIS2sPeZTSbsw6Q6nKZgsYcx75918/iL1q9dlLrctcEqC01zc/YQ5WNlT4PhtSS+z6s3po
SxAu/PnxK3qOYX4A7zmIXAB31WvxOW8SMdqXltC4foT1ewiLdeIvAFxP6pod9xEq/YwHlH4MARW2
eT3SmD05I2d/WlsfRbP+GsNA22aLIgaWlT9aNgjanMCAvbnClQhMWxYBiW41KWvd4E9anjiOBHf4
AIjpTfI9YdfFb9uRkiuTsjDF2RVTbH6vnFi48jtSdkEJgZVlQBMsrKOXlb1P05OtQ9KVri8+r5He
4wkiRqLQb2bon4KmXcD8oDpP6hAkjNmjF6xjp53pwzANFPHmmsL/AzY/95cDYBeBQRSt3ceJxQrG
drKqtzw6NyULE7YueNEs4upHjSCBPaSYxYZDi9kOVb1JaF4ZMfRbF5EVg7K1Aqg2BEFQwKQb1BHz
K6D8iGbSQPBKHkaUtocUrntz+YxKdao8ks4zauNBQv2MflHFkMPKEpOk+/lOZvlsZ2F9lcFegY83
zzvMmg9nhynB49GCDXWvJImBArkQJWmYCaBzZA0MFvTeoRVf1OfJmv1Y/Uq2/GSQ9It9phYJHgYc
Ki5JnKUYk96jfeU08Lxelq8JUWZCtZgCB2PVidLJufIh5Twb2wY23wmbmwbYZ8gy7cwCz0ZNgctF
+Knze8CnYewD+R8WYr14uRjDWFXI0JVZadnm/G8x/FDZbtVPwfF3gOo09LszxSaFm1ar3g7xLhcF
kcs7U9b9CZqggf79bOUhGPOsJ1/FHA7Hot1Ne/H+6spwmoAYaT5iPENHUnl+RkHrmG+G8at8JIT1
qWl5/uIR5WvceBn+GudgpTcwwEkf67yjI4IRgjXG4UFRiqyLNgosIGiJbYH0Q9XtvIKAuhecVVmG
IBlhzSkANnwOwb+kdf0TG9IQNq4MQzKgp4LDpjprvxmk+mq9l+ZFL/JgyQnRYe5pRTRac9cWeHre
1W5myziiltRf/V9nF4Z/jXvJD2DD9gunQXZc+uFHCTs6+sFee8GOFFKanSlIAxGucD5sE3sJOX94
Pk5iROyDx0do+turOtjzv1rmdSCDftLuCCxrur7CcS8yfxYLJu8CX/HpeN1Z7xiahpurEi8odUno
LDWPafh1hPjKFPJI0glRcCrKX3VVP/3BxzGUCFlhy0O+urv/5FbIWHos4lLNLQZCA4fnk/kwRJYR
kJRJq7lNI33wDzdMsTFRwOBbM54RWAbTqHiOcW8qO6C9XQMyUuWTCjXhEU2xOYErTdwt+695AerY
F/m3T3+HGMxr9VdQgMNbpegkkYHtfSMb1CWUjYyg8f89Q37rCrqK5UOWMq1Av1aA5hzBi0Sp//7D
BGeChsouyw2gnfXkI3F4Gb43mXuVeBQAmyU9hbbqCQVAusYfSgwnbi6WJwHj5g/7K+sJUC4fqiw9
6aD8jE/FetcVvELR7xCHKf47ldG389hRwmxQtBqpfIXFV+xOVpF+iucAJc4hRfEdNOpgMkAH5l/i
kM7m2eRciYQcgGfRseVsCOg6jPh2G+iK9uQ1uylooXR5x8joFDfEf2Bw4ZoKnLPeYoPfgTJ3pg99
YVWIppnkpmv3cNdBZ4QiHKtd2jDviLwaLi+i44PTIghRvFZJ7D1GqvRVLe5SWGj15ceGJYvTVL9r
P5Zy2DMSaNWhGjh5S/fBVqadZkmvh155Ycn6GZr1FdhdzrwQgHXNIyGljjc6i7b0toncexlTH6H5
Mk2nk9iaE/TxHWtjFfc7R99Po0Fkc+u/Dx0Jnd8/od+o12GMYyCDQD29CuuefUlCPCFu4ezesZ/s
fXKHttNP5oICmZR4T7svXslfCeW8y7Yp6NT9ve2KCZF81BWcSEanqo3O2uNoRXskRrRnx9Y3WMea
FPgI/qKOOB9FHiQ+sbX4eZq4r497NK3/2cda47dOwiUaGbmhRZeoqvKAcYFqMHWeaK25cxcPlhaj
P8nzmuX6DRoeUAdxvOY4IZLe7oePDlBBJFbckYGf+OFiHJbVBhyYhAh2n/H1SiJMnHms/2SRXct+
cNSkv8tCTCviLd27VOB4bswSTEfCEcCW0tiyvkUAD77ZgRKnm7wZVQ8lTnkVUkXVCJjgr6X+mdCP
pZJ/vHLUS+YJrJwq7CHAPp6EHyCCap2xxTZapsU0iccPoyt/xF8cDwlJVmZ5dhyLpRT1y3L9rf/Q
L2cugrOdvwjWh+aqTtGFrdzpWykaky4ysSrfdbVCW8Yr5XzQSoBcAkPQ1nX6Oh/TTzpYgMCvTTti
AypQEKX52Uj8CYaYV1wLCyPz1HI2G8mjEubhmtH9teatuuOlYzCYyDwfkeYUOwQtUkCw+35Xob7d
1Vz65wfDWAKwkjsXKiyTuDCAXS0Pd9qTGtMYutEKbdQ+AE+oQChCTgD4cw4o+ClQ6XfxoJXLzshI
oMR/A6/lpcoLyMSmGzSXyA76nTHJWKTKoBKZ7VxjUjZlaH2mn/lNLZmpw62HBGkxjKRIMuZQMCr9
fUL/c82Y7s7tWMyjJiVDBuY5Q1ld837D6xuKIi7MqYc1Xw8tOCJDAPNzGxD/9xIdjC1wjHvLiwts
Y7LYPp/3wFsONk81rpjeohNcB8T8xogY/s7XsQE6ysCTo3UYsEtKaDPLmLFTueliiiMeAGYs6unI
0NXMW7iFbV+nMV8DqMOTdFhnZokq0sRQw4XlSJRadXmP4ouXjmDpArxIwb0M2mgiBHNarWPGgL+/
E47PCa3AgB8UsHHngAWvtSe0tgK5usdMyG3olGDuTTN17Va1ABMBm1+8lGwc9YKpGrCUn3OQ1pSu
bOFwDW3d4KGFRFTnSNri2605MPxzlpNRNUoSfmZfRnMeq7eBkmibvZ8iCCehCtdeYBQxXSnUTBvz
T+epproKXDi9OTlNkVqd1odmz5+L3FznecAYFfLL62D2YNZ2oGo5gMVUsa9V4RmD+5zplS5u6xTw
TV1F+8eSdkGuvB/FOkssN2HWI1+D4DUhn7AyFW3xFoyex0sVWjmDA6stBN4iQpKdtPYXfESSKa42
PMJnLlic2O1w0FKvr7QnGUiTqS99zmyGUvZ5kzJ+9BDO5EmaNhNMz90LiZ7txFu4NXJjiytrOSpc
5C0QR5IymamwDTT21It3tFzsTnAy4jKEszd9ZNMWF8HjAQvm1h5jWpvABR6+1OLHKJsVz/Rg16OJ
NFRswY4OIN2kRcYCoZHGd0sYMlJTcbuQNSheniC3Mm/XYycHZhC3/Lb4+VYX3MOymYOaWsKvz9CA
B+DHCtA8wL6pj8y6xGvOgfbBBMlykHvdBFHkm7SRvaU91+fKMdzy3+2AcEuhEKq/oD/Gm/caPlGK
MTpsC5gLzp/bM+jx5B55KNeHXgjfwQJWGCjsnkAF846HufJDGA0R+1Q8gwFPeySMLEF0VEV8BIYb
7+MiNVhr86wxWLpXOKz37r1o8UBfZZPwuIaQAwh4P/GagPw6khmLX/+Q1ejU89s0uPj9T3Ue2SOm
f65k+lWeXkpFYHi0MMHGwJWU+Zq/jKsFmQZN7YHJSYDCY5ANwM30/5TKg4OP4O39bXWAmlu9nkMD
abH8xHB58Gz8oEuYEpbdwiE+NKZi/as2lrknKoea8VL6+98k6CqRzmQ9Ws7PZgP1SoFLo6cZHsbt
T3t5b9bZ/cpLPC29FlpZ2D4IdD0k9nZerNDDmd9Gr385zbr3h3sNV/alkdCpbAsj2IYP+GP65IFS
0cNNT5gHEj+MtfkdLqCiGJN9U2gg72Z+/u7VagIW96EAcyToN+69KAOBVK98Eg7ka+TIaffcyeaw
wogpvpo+kbogRPQ73q1jrO4GrsoruPTzAMjXTSpySkN0QEV+KJwvCr8IT33f2/5e7RyAcltqYxDc
Dz5nU8htEmwhFCLUyetJGNZghjINs/C6/RMMXgURDrUY9W2VMXCDJ42kRT3Wwy9J74n8VlRDhqSs
Pjc80QN+6PcNbNJt0W8HTXhk1HOC6ibbq9v+z2KbWNardSRw2CujUu4VrCyxaAwdYPUDix86QTIJ
3kagDAHSU8MI31j+3x6wrdfpbVd8CWbrSuIcG5b2drUL1ypVvXAohulOvcXQmWOnMtTj0YOeb4K8
rnxH/V96aJD9LZIU+cADYGwK6N1PgW+f9MJHpigRNRe1vXUfagSMioav3t3XK9JUTBYzx9TOfNJr
IIit0cDp5qKfAUoWdXAKA9PTmQl+DjIdCOqmLC1wFwB7ghZmwRouTmLgBpFrmdQkYKUY9B2cAGU5
+JP3RWyIeDYgX6+HfD7DIBuDen8C51xYC8JcDKOyci1bOrCXbgippE5sibGkPM0+wOH+jOvhml/B
m9sHtHl64MpejWYE0ZfejU3UlHv738z2WrYrN5Lo6mVuvnZ/qdd8LU/2j1lclT6Nw4HjjjwhIsfD
NbbTwAjCryunY8YIMcRp2A3kuwOVdx4ocxnSWs8pklV8tPKO6BeltYwqFQE3KbUwxajqrPRie/07
KwhupThiuQsWxaHJxVnPpp/mgrkiTJh6fYTK3zpfZs+NziFD2/qmWz2aHo/hOEBHB/iJJ5KPQ9yO
w+CV00YHV17/TI4Yvk8t29ZyKq8q9bO6aLEjHJih9k1Pzjf+g07vaFTT/c/zLN4dbeB8t62V0mmE
VDXCRRfIw9tEFQJ/diMcDLpWFrQWY9hIQ45yq+DZsttznqDQcj+yCIMB2APOhOXSs0n6r6xgn2pm
L1EQsMqQvL9U4k5VLmD0MMmiLSWaRUZbRyzxd88zZvA0zrkvXnsr9R2lVt8qgsj8oBD+xYsIRRNi
LvFAkv866IEXozS/Dfz2WYIHEdqpFQbKTuP08PdKEJSylomxcpALNw27TBLlq8sANIHTUjZ2c3Lw
C+5dWwtFMZX2P+HMoyymC26fqDwah5DCRJR09gliig6xFuSSIClhKvvEHjZHg/8Lv/uNl8jtDQw1
XUyhX0gA0vAqZTLZ3u6DImR2dx1csFAil5xSwdlCd3ZyTyAZoVARRP5cq31hmdtG+NwYovLLG3OR
KsHV6+pdggZSWiVa7SWWZGIU0N30S+sun1Mdd2o2TfEBNAwHXlLUHHS8diqv6A4FHmpzdnmFbHek
j0Z97SoPFDe94pnjYix+wPRqG4K4TnNi7Z3l+AifTUSXc3VGPXfVVsNtV8H/HdLckg6Cucm0Ahgh
9k+XHhFadr9DjrASPJPsDYyE9SRpvXtt0HA7PWGAS9YOom1VGzv5doaiz+6Awdn8LzvgNHq+upc9
IrEza3rOaNMCMU3WHqGhc7iJPM2dl9U20cwQgnJM5KZZB9uke0DslbsOBklxiNLeUxwIsRRQqjff
lMSRP99r3pTBigtWWKLT7ezJeH4FTDCpz8aEgb3eBpgIQazVcDBMALGBvmRW32jKF9/qIpaPWekN
Gz5B5Jtc7XKGqJOSN2QJl8OmCjcecH0jHP+EawESHC88vC2c8hPG4fP5aD8CvSdz6GLaylj18EdY
sFdV9YcQG8re/gDOwlh9XS/cagLDz0rJLhjarThD/Zu/c3zrONa/hHjuw/gcdev74ZtV+w9XUlF4
qCOCL7kAHg86KuSvSkKLFoQTNFEcqJXDPI7r3Cl2WAmr89PogV5xRHPkRRITgQKlQRM8VFPa78dq
JOzga62x60YodU2Fs/aCIcd/MouXpJejHhK4mdJ1vugDxfUkhbxMzekqttNVmr53Z/qjsGmKd9Ue
SX5XUhi1t9pRqsRx4MAiGmgQvlraM/cZUdHDnYEaBZFKjwtLANU8bbuMinKzA7cjTSzlyYAhsWI+
yL1zlbSlx5P4lRldvvg59MF9lou19yenkENwdjfrns8QpiSxDiEoCrCddFnj7Ie8aRMbeCzy6+nY
ALRlSHpYGqOfTV6BignX4YWKK6bleAvNW8susC6QVKbVYfJDuzOuiGvNDiSyf2YNp8d+x5REOYt4
qJacbh7KAG21mdFYAhbiAkeYRXX/IW1eJekxSb7MYiG8ByUNWPIYBqmcbo/qvL9y9A1HO4f4rpTS
J2l29GnB7406G5lz+6xCm8AvPz1cmp2pyAoLl7iABenZFEwM4g5849rnakxjCDYpvfa4MI6HMpIg
9bL7KbEbjPG+kzBF7lYfh9HsoxhddbED+jQH4w7aT0bH23cx3hK8+M6l+m1LAMKNNrn2eklFSmiH
xB2Ja/wTa/gmXyec5CxaMIEkL47reBacFXUljRSrgwsCcIhPolPsXEBa0sixsq0lJs2Wa+ecrol8
pY9SbtTQC7ia4QkKmMd0tCViWuaacVNdyXF2vJAholZyxIbDe/WAqvXBWJxYXZYbiAasGGIUbVg9
HIsX8yEgSMqNvj6MjZyLcFm6GIv8/HBAtscDIjq3zZADSn057GMWcS2woCjv3OzoKOVMVMiD9dhv
LmiEccGHErgFOxFio+6pDUcRF8Sgku9M6Bti03rzCOmr9yLO+6hZBHri+cy8Kv/eAZ6vGNIZTwZf
XTYBma5pIE/23hMoS5YIeVFsfkpDMMl1PFmX8kid7WKdyx+6kmkNR+NuXUyZxHq7FTyE07qbZfkW
1ZQIN+TO2dNQ1F+qTl/wmm3210FJGd6TGz+RtLHQHbI4Jmm+VTWeI/gvMEoHVNjnGnuVFJ91s2Aa
Z2h2xytHX9MOBkjsYCGClICZV/SEGDBkXWwDb67p4XxVAt9pcE/eDjkxBOtYgk3ujiISxEabWWBX
Qh6czetFKVHhENNGNoTtICXhwOCNxdsum6y1HZYUKnvdRcUbkL4C0WWjWx7oU8IoBj4KiHBpN4nw
DCDI5SaaDG5o9iYJ4ExJDXBP3KjlNB2y4Pw1BxOvcYw4VfKU2qUiv+5XbYb4ZSWjWlHouvN8N6Af
3ht/ZoKK0SboIuhh0HBWq/zqwsPjsDQv/jdprEozTHza+k2WMg+4GSeb0TliUXrQhqsHf7KcZ6xJ
1tFD5Sr2XvD4yK7ZM2zQHT48GNhX8G32VEm4LOnPUlmY9pJzPSTKDPAl8q72eWEkToKR2DH7JBWB
/oNh6lM86uV+ffTPEuuVPC/U+bA3YrFE0N3uRGhiHzljGGMdHpmw/SwEtgbGYLxP9da2vvXdOHUm
77afvWzjqgkT9kqS33SzyxJDClJAcgSFDdPwZTsD+ZSKrIB47o/IazG03HhpLwglzzwrpYONZuFL
dFz1gg9pdRxA498VYMEyHFVspxlBP204fWA9Kp6alhAZXIuw0be7wCuCBpoXlUUFTbRWOwIDBqk1
3TIgMJYBoI2m3kfEYmQcb5tny0PdFmdkKUBB/DfBMxvpfeLaMl/SnXKyCgASqysosHQNjbmtptNc
TXYnq6rXDqONfJ71+D/+3+FYdC49qX4zq/IJ516S9qtO9FvIWlqF5XoxgtHDbJ0X9EA3LEGD530W
eiKeDl3BTQei6FTPEuTA8e3eVLDragq6tBVvN+PR7XC4bdkbxlz2Ct8/EJhHvWoRL22LzbngzCsz
4QqxmHTx9G1ZACHI+yiP64dVHtrErdeMorNDFS4JSCXQN2zLcHYL6pDN9Le2g8/r7fGh81iA4Cqq
Ycdk6RX/SQ8mCgQliXSFFcXs51BwaPjV6DI1tNvCqP3faDb9jSO2Z85R0zSUCCYUBHJF2H53Aiiz
jopt0fugo3EVWB0PokBUMkRvfGFV8+DcxGgnLjbgYoNcCnM5oEr2UdBuo+NaFzb2ik13S6iZ/R3N
BrBYgn16Pbm1MOxdX1ILjlREbbVxhCNod6Th1Dzwps6d+SXOUcpyMvOcdA8PzZQlSoid3UIU6kdO
I0uwW00XDZPs6cPVrtDOcNbBY/cucJqI/MORa96xqPXNcN2fH/RuwsEBljYnOPbrEwJLd5TTrvcZ
I9sH8NWy1jLC45/bECe7YqGZ43wrzwlSCG04tk9CkO6noQq6W+swnhzDwYRzFK3PBQmw4iN0pLTb
Lq4QEvGBcFqyrvMZR2bpYdRb0U+8qMSHDxbtaOdT7f33Q7E5ull1zzeJCVu7iVMFevsCb/HEbL1p
nRaMm8FlqLq/p55R7FmVNMNkm93helSK0cgBuzmaP2AWNp9I9GuZEtJS4h4rgfG0lxgNNKUBpzCa
JdkgM12q47VNFfVpBdimSaMDQSIiy1SJnyb/lEMbq2qbTyCmN89Xk6CjriOedm+THELcSCIZmHzc
nuxJzFU1uCyv1YPyb1aAEyzEtRwKI1uUi3ss/07kUhJ89HkoaU7n1Q5Z6yMUbdTF7VxfyZOKrCJ8
SO7y896SWfkEEP2fLbMXmebuRIjkKbihE2/Ky03U8EpKP0ItJkvJOk5GUZZRH8QNp7fQtgavoDi3
736yAAXIsaMoLeRAVpg7Q8zH5HgammYbEvjfm9HSOpvb+CErTvDBdoiklo0l8rh3K9gVLTmLM61g
/RPoDh4fFudPYjK56cYpK+okPw0Z3xMN1ecZwjFZuORzU0cPHFpcBbPyStHMshdJ3Ge80tx/ZN/1
dxvfYxAeCeSLKZ1AxGZE0c6RCwOpJe6072rabeV9+UrwuPBvXHEUpC64F5qbMYDc6dheQptoTyUp
ShHYexwaN9AuC7swojKGJQdXlllQsIUCwV9wsaDIHv4Q+3Ss56IrEE1U8plJWIjfKAVkaEWkBGVa
NaMdk1VVR6JuzYc3cfyiXo/VRQ3OXEp8ySzJg9YwhM6XyfExMxnmw70DmSrMr0JLumn48028gppp
JIfvACTXscDTnE5jIXp6mXh2kwmm1YKoI71VxJzczIN0ZAdrZXAZU57MrnMWHkwNUJyyELAQJRLi
qVWqa+CB75G28acr0v4vwtZjJKG3QRumCCAauAnUJ+qyqqolAbUqq6cxH4E59WM33mE0FxZIzG5t
wlDFLJnstF/bxJGrs6X8yloLh362v7EV+KNCJLFyvFjecESI761G3DhePNSzYV30YFzopFahx9J8
6F+9+c7U4I8lpinFZSnuS5iX+qqBPr/P94iJUi+CO70lFHXwbnaTqgzoOCVkwGy/V2o2FFkgsYSy
1vL8YUf+jif/Jwi3vwMQgJIBeTkLLGQS10Ab769/9LVZdbA81+nlC3g/SA1l5DmK/21F5iabeFqK
kW2UVd3AXTO2rrSi8ilAIh6UUX+vebn7AktCBA+kT9enGb+l0hi+eQYI/GZzURZmleT7Kr1czGdU
n6PgyhdNwh+mglk5/x0FjSBDyIyeM+uxXOzka3lNJqsYK2CdLpO8vN4ajPBVl4xr0I63TQbLS8Hf
ZXadTTlYlGKgny8YW+lMzlQW6op82Qqcejxv1Dz/9XxYI1UWlZZg5jRKjCSmz0ONCiUvE6eFJu7D
EaxJLgb2uZTbRCYR3YS7nzrhcrahQ44j5hBlWJHRwYGy7zD3yWsvnzdqB+pwg81KZPrEi42mBzza
am2mfXBjfOEgHfxJRrA9BE7j3fwlgUJ9b2O+AodRlqi2V0Cg+xlPn1SOc//y+sH638h2LEoYZUGo
BZjlLatVXiFA0zUQWXvQNcngY0uX02NHK3yL80TAj6ez4mDePyWQOnfbfhC64u+alMK+FYERWb9e
DNE+0rNKq2hlgf+qR2rTK73uH4HXm1oFL/B0FeuOkDLVzxwS2hopo0PB4QufOLYViAnHoNVp+tMq
/SxwF77Y9OJim0pEd0K2pqjKEmgX3865RLrcedBXZEjW0SP3TbvHfzXByXpdS+CdVZXonTls8eJb
QyKjqx+Bq/RPLX+s+BRYsrj4tpGKyPQO9bC4bRC/IRovc1xXuLiiCCIf6KHB4905CqSvVmUUJ7Qd
D6z8JLhlPtw1z+nPG5PxP1+7uPnONSVAX+hwRqycPfDWbZfcbrmwZqdwxczCI5gafRsfi151QJ6m
iyRMzKsaNGoZlBwgUXLCyJWsjm9l5MPcTg8YN1iSANAWXi+6UI4jHNA6LobAMPEWVhmjUCxYqrPu
z8twPITsz1OqEJ48RlDlS+5CZvbKgDy8K64c8YWg5eOHCLXyRdz0/Hbt9Wu6tXqdK+xavWnYUtW9
m9l0tL2aRO77avlBwrSRBIv+gDA2JvbtBicAZi4hz6dxK0chyMn691RSdC/tUprTnM60kuepvdjn
zkmctnfCM1D86eXjSy0slblksr6zQusIhM668WWzdzaT7suAC29FW0SbBsDe0h6a+JqS/cXK4LrR
QYCEQ93OjsGWVzf4PNP3jv4SpGLWU+EjnFi60N+oz6XYYUe1X8k7Ck3/++rkFeFTdOKb4asXSvSO
z7a1d7fIDKlk+zP72e8QweojyZfKveaTww81f48cA2llgavwD0itSTUGAhiUwS6OP660njtVJM/f
Vq4D04q3XAgy4PoAUVICsYfuFfKSppCPioCxxrS963DGCsRvxuuBjl3DhuQQ3tIcYj7X5w58DM8G
7YJ2cseFik7LAjkf8DyQNXSIy4Y5cmXWqEjBFPqJYurybGbOB0z7g87FyOd5+w4luDVt2wLrc145
IO7lqn+F4omb23RBEdOMb6pLucKljaJGlqsnOmkR7zZYlPoQ/32dodE4VUK4etMjaEiLJ0H+/xtD
UbF//2hNLhV7aJbq/TeWVAnid08YKM5SAT2rINsew1fd/KixH2GwPcfjPNCHS7fEZo1+kg1Le+Nb
//nrq7YL0tAHgg1SOGz65u27t8EIHcjiY6yqHUIjDyGw6iFBgt2QsmhgKu30X+IqFQBRW0ep4g/B
teQzWe4kGZzil9llX+qlvgR127U8XxS43K8S32Z0kQ2ZpNq4iW8qBIZcAVs4BCQMBjqKP3u0pyEg
KusX7gqBzeYNW8Ua1/0g9+yDTdyQkKzBwhtH1fQX+FsrdCDRCB6QR7zs033Yse3kgv9q73vfnLus
naTfbEiRy3M4Tc8SW8VvfmfM8WOjqUOnxdRbLqM9MGCSv7cDo+OiB66jAxNNXXK/7QSw1+uI0LzF
bCeL9M/aZacNw+c5mYiLKCWCNN+HBtvbw5GLxqwoPZrQxQpMHDYqCn3StPSbMNkBkJI31EPIrXZ6
ENG4ooT/uEh9Rrz1bb8OTZutoVm8XWTY7fP65jYvWr4cxzZmxmHqdSX9zkvNAK7IEFX9snTrX7tZ
dKilcw/ZxJHjOstgQFdqbwh7yzeeReUBUHzHuGQhbHyb5A92pG0XDl78QAgzwcMw9BwSBstdZ6DO
kIMP3AuYM+23ojnji1Hqx7QtRNg8vkbMtT/PjGn2AD8UvU7V9lOko9HgnDvzS6zQEOxDLVHU4l0A
rNxvJ3ZNgcqWfzMgBrpUWHEWeCRvGlWidf1iadiDweD6aCX2qOOobm/RtIb5Qgl/8J2mt2jSyW/2
snlAuhAmrDAqxEcT2S251sCog0IT03CU6527kfDPG9nldsPFJQbe1ly5k7OeDaFi5nV8MZZOElJ9
rC+vVE5vYvR38lYqsY5ffxUpQY60Iq9i5gzNm5e3Fo6whg+z2NIeEHDlRf4wy/YtEgmUUHhTrEzi
c2lopxfKRoeHGmGXveiScxL0Hjma8H19InCqPDS4+z2t49IIqjeMDqw3kvvzMtxe4be1JxIvMCDU
hnHozDv83otkuiAPBPcm+KPe2yzJ6P+nrjxUW+HoY+3bk5wdq5JQTyjkzK6/jgUtGqep7X1UtPKc
Ax/etXw2Gjd81w09Fa4KsiVNcvtxjkj6aBXG1U4vgnuNE0gdB9Sqz8KhGDeX2Vt6I5ejM+ETuujN
YgKWNMyJKsKU0TfhanG9p4Yjvj8g5TkgSTptbXTYQuiC6JV+hYtWrSZNFBjmp9fYejiYlRsbVYPm
D3hHFw4hNShCyEi2SJNcZNlNbSHboK82e3ierQqDkS1DP4oONCA1sOfIfG9LAR/a/qNmA8C9u3SA
9iDEH61Fr2unXRin1zps5uLZdgYo/MBk0df8wHdabWz25kfGkX4Y8roKz4n+S6M29yfl2vQr4xAV
aNMqikk+rB2hKUCtLhs3GUFcMtKv7IAepO2nkF0lYqVjXcx3di/LqDX3GZgCccKP9g7u0rQHQQ6A
NCFB5jtAzeckD757k0Ws+RDBTF8N8+vx12uK3yR1OqEKCCtf8mymu6fE2kwxgVLsGWCmKQrd0k5v
ADUyN0TPH5rBDearJdSjbqInFCluZ4A3ONJNw1OZ4R3GjjbBYWRmNT7n7EmxJ3Z2dIeZF4LYnKLN
m3sykzcqAZQDdvqiUtN4+ZjkIJ5VRS0mBH5zTa7xIVUKLEzum1w9lmavN5liGz/T1tMVQLYpoWEm
XImBr/2jikWOboPVRlTzlSYj6M0KOtHM+/c+2ea0/dPxG/RgFBn0bRAGedczqv845qzpcJWU83Cq
OUsA8AWrAgbwAmPBWXMi1FBMy3AGyei0vsk8q81mpq0MsXTMy5mU5unkV5Svg47tNdnepL81BYgH
4l1VPWYE10A9/zjX7VDdesInRcn8Hpg2DQDJO44kDlrn7v+aCxPme+kIhqCa/rNBj/DjDUYYUZVj
j80F+ZZxJAxM1ZTQ7mBVshX4nn3g2Jdss0PPEueAIczV/2haRjAUOMXwR7vC+jDpK/qg7iqkGWnU
Ax/Mau0v2XeX8DqGz3cMw8wlJhn3DN5E1LJrP9JhvzJT218dOpA2VCzjtfHU/ef47fgNZCXbOLyO
rhys85HBdEm2JTXFyxu9NgbcOLJpuLHcTzGzi6cf5gXpJfalEMYw8wT+BfOQz4JX5pOlJ6mCWLj3
ABqL8hKbrulaw0/HDUwScnmwURG7qat9mQxEWtVuVGjedyL9MZF1UmpfiG3H7EmqKj5qBXQwo60i
YwOzlETqM1hhEr6intxFL6uBcxVwzzt6UmkN0whkCDcr5yN7jKo3qmI1QVZ/mLZU0JGDx9gIYfcJ
4U8+9dlTAaGlRyWqZRMey8Txf249wbJ7n09yDzoRo6WzE/MEz15GyPzyAjFXSBWlQIuHjwkZuuTA
tig+RAgEOhfrGIH332qNbhPW7au0kzsib6gnZRNrwoPFrj+KVMYgXUJd9rjPQXuGyxUfnbq+iQGP
Xg/bmaKBtCse/xCdW0JPemccKE9fA2QvARQpPN3F5wgcfmk4ckhh0DTBoTuz7ki5jLn6T4us+3co
PmdS56IAr/E6PlxnLTQLdNL5PbLsX+ykR8wwXBOeCAl2p0ljFv4ARRYXnnCfm6gqw0v7xbY8iv9Z
s3/pHtydKRA3i3l9mylGPX8gyKQtlaRKoRv/AE3BKPNlq0r32Xh6SgOl+S89RAu4jku2LRuKfVli
zTlrm4re3+9a/wcRqZJ/7uZomdp/81Gajw0LcnDJ/XbCsekCieg4TULFUza7mbh+LwxufvlykM2P
EHrNX4I6Yl0np7zijh9BaPd5rDVIPzpibHc0sHDeAydiuPpUoqWKvS5c7dMi6apJ5dXqTa3mIw8l
Hgia4p4MHNx6EJ843s6U3RWAHGOlvEWP9vJAyf7q7n6LUbCwhD/a9Oy8HqugQDKqMpThUVuWrNBP
aJLh8I7ggkUgoC5/74hPfNc4iN9VrgbVsmbUBYG+ll0Z6dSIsGde1bea0F+ONngy7+NFjjqJUIV2
ltuvqwk/l5cfWQwtrrxsqn/1vRgtZH7CIKiUeK3PhgS5IyY3uLhE5IMHFLxkLz7hduQZDtMo+c9P
FKxfe2pDjqq7++EZbI7AihXIUf+dnltOW3HRFBschSenM7ARdTkfgP+x8myCw4QyjAZSR6361FYp
Bat/WD7WEZsi27O5DOQYKKBxRhJJJFBpP+PQpZ8minmZ4MlubSlNwQuGipxqzx2V6IhPISmrkjUd
50u4QBk4cciv/UScqLOXE9vDGCnfqfLLutT6ecb8Jn1DMrZybIG6Wb5RC0rLWQV4q5S3uB8zWELV
noIruTPfZ1P4sJse56NRKYVMUe8FpsLVfdqW1uqyaBT3CMFG6csuoaCmhrTlE52WSRRLV3NftAdD
O4daKb18ug3lsbkb2jspnsbecKiODZgTiGHfDoz+YmHNzt+k2+I+pt7Ovz8lrnue9/dlEAp7zFro
JCkrEs4KpR1cOsIqD7jGWZ5Hi8anBAKJgNkcRzCuBwGhXCwi08WPT1ifvlP17+9Fm/E8Xr0zVS+9
TpDUQ3r6jTLU1gZiy/uQDmBTR/Pjses8H/p0X8A0rMGL6nKue1J3qKH/aYsWgXe9arDb9gwFDK8U
SaGgHv6mqzfZknfwg4W2OGpJWX/Pv8240g0AuHnar3Wm3O1Qf3GBw1XMyAKmsw7ykI7g4HFIHiEN
megwWJcGnXw0lHGJ/Wz1HldctxnZOsnQmltlF5nLnRxN+AJ0c0ZNXu6BE1VwCBco7gdmPbZHOB/9
GEZkHyMpf+0zk5muJc0Yn9XCDcro5ngSv0NezRtCzLbhmERb/8VNhN863Emk2Nc6U+297yBu3DLj
jS0vRwFNAArmUaNiwh9wII4INgrhg+M3YLLIRd1PmCwLCrlH/lenlBP0pcNLjFlSo4nlct2UnwxU
k/D+CEUYlhj1ErIi+rHJDxklmk4BpPHULE6Crl+fFLXSCzyVwNpDDLUJxNS+QMQG+UU19B22Fgx6
m+42LcQLQEYjbYnnLrhfM9ILeTgvoXHJiiFhSPVdMyZO2IImuS5nfU46hmM5pfOpNtNV72UchqOl
D9TF37Z/0EqGLgAniTfJzgmDfkal/PachbGmncEtuaLs/jxvilCQ4LcWSkJVhHFYVFLT3SKo5hr4
/4qGe6LaufzQdl7sEg2RZ8t31K75jrQYf0EaNtH2gmc7zF0ga5rtKTstXiqp9M7yu2E1Ue54wo/z
ppJuUZ/c2TxsIOHwb9e6Q4VzjnMhmafDjaVURW1plKIsKZPL8jx1VxHy7ghANg9aSkbZoM8C7Wir
a0EHk4n/jHy/8ojWhe3MsJn/rApIHPUxGKAlOM8fiRkpdwS8Wuvr+mWMKsU1g5zl11raQOkpOnrT
z9UP2nxmVU4C+3XggP8NL6Mn+FBkEfCzHF9xSV/PaPggtKL4+kEudnmoFl7HjBD8qbZu+mmIATMS
fH38FFG57yfsEaRVTllLBjgsfChKRdYRRTi+jN2A6KyRdCQJmHI4BhUf8CK+zAZfPNeytNk1DE9y
cadVhZiqSgbLjJrvnCCAneSyBNtlhPtAuX5L6mL+hg1+yvJOY+8DttzgqFL/JZH2FedMlH2h1P58
jbw57R8mYLp4W9GV4V88UckdLh4xZfrHM43aenYoI1tRE+SftgphhRookwAh0p8T439L6Tm09Od5
eoPcTu6uU15J+XBqlo2FAO2xZTY13sl9S3c0ENJQMODhsJb5rxb5v+rRSHgkCtXJ+ucncgiamUPo
u6jZlE5bgJwHc/VEgGc5/JZdshiYwEKVIeaRp/6HY/orTZAwJOlHjFsMW8fDfUFhBer8nh3hz8Mq
IMv/VEZRokLISKvn7Nvc3VsCi0Pb9rwQVIV4ivq8coAIzoNT7nQNYwE576aSyaR3aiWluLELbvJI
CsTP168xQpmB35/B3y1YCkSIEOJA0yc61ZUjqNZmH8juUmZ7GZBNMuPSBF9q9LmR0gYydWBh9zH5
5rQN9ulyf1nvfMClMTn3GolNka6tLcPAC5vEc5vpsAKA/f+UaranGwouqa2xyQYfTM4xHT9Di4JE
VQ06wSAVh/U8a6ItJrqSPjBQzOD7UTPNXWJcUaoYdiG7lha2dEJA6tWT6zzzbyDdXIL1i2RUhR8d
w0z1jg8exmaZdDXw6OmmJdx26EUw+7XJWeKMyXcz4YOCnKQHNjSN4OVmAOTX7Rz4p2WSEEtJ3OwN
UGrdrrSme+iHSA842pMiD99skYxYQ8jGJbg/506YJsSevAuwP4Ow6mzzMU/Jjc+X/wcdhyYiuu53
/Ru7PuFvtWJS0bIaUipKDfDId3Bf8zl6GDgahS5Ln2LBKVwLjB+A+TWFj47DumlwK+ENUoNgkBZ5
ykM+d99f/UZ7aHJQhirjX7Cr3xg97TX2WILmk5tPbFfR4RVFZT3O7tPpi5RiIjgM+ilNG3EzeThX
L8pGa4VGo0deUz5+xMTSwXp3OBuO3BfCYRisT3V8wu/r1xbvSIxMtd6OxM7jZWqo+xHmCrqCLr7m
+LOcoxBb6/E9Pd7xGpKp+0Lo5iNdHvPGzVVotwjDZDweFRB7+MPfrt6n641ga+4JdMA/C6smv7mU
eJAoMfHsVltSwXMCPBuUnDV/MarVgxf5xCaeCi/wYvThtaABWcEqFfGCBnZcGLnEz+5WeNLKNkXK
SzmRkAupQ3ilCvjJTVUUUUCsfC56T4uAvTuEbm6v4XFe8ivivJSNKUXcRF51j0j3/kY7+lMiCSdW
iMh2f//0w/oZA7YcyGHks6jdyeNfFhLx/h3jc9d4JA0DYkc52VO7pOdUgp+s98RgImcKlYSK9HXX
LCV17e7HXPn5WKojESsOWtVUAsHA6dGdHzY1jm0bUBq9TTQYF+QwtFRr8ALM5cVHhdlx3+1IBLFU
ax7oe0okjuTQaaJgAUcF1Txw0Mbvg9mJJF3Nb3RVdchKPNV3m5fzGgO2Z3FvjdK6yhQZmdl/IgK0
TbPk3JlPdJOtd6JpioGymYzv8EW4HFcMwXOKwDU3ohdaHBY+nsdylN4lFDXsj2rE39RLN4zmfO+t
UOsN3mUpm7pINMEvHhvPeUwkZYS15RvkhFkLx/UW+FnADm4E6WZeAeFtRdDRINn4ApPxzIl9C/x9
nyjFI9rfzOonoeuJQ6q60PY9BCLPFQBDcj2pUjm51qbYaLWkE8Gnx4ikKEaOKuXJ67IfMKUc7Awo
UVTnbhf7zC5PlB7ZhDT4cqHxJYdL6RJOUZq6T5u9Lfurt3G5j9u/hEf7F4V8cXwMqXp/4BRwa61F
Qft+0ChecXEZPaB7hPOClewEu2LjwVpMnM8IXgsy6Ng0cxLcSmRrhUPTQYDnKZ/symdRGWaKreFw
3R0bDZprAowveWlVUi8qwMJGYxRE5zXvFMSLhsK3tbiRQ7Z2l3EI5Bp+yUHA4KKcMzYRwXlJToea
wr8gw3KxfwBUmo7Vt5NKoBN7dzki9G+916MlYUlXULSZ2Ngk+snLzhjG1JrjMrJpLEEqrDZp0H0z
vxIVX5rF9s+30k7ZhEWsK3pV7dhYzYWMeaC0V+HY3h3J6pLYJTWDOAWH3z6Y2MJi8SeSjav12zcA
91f0bXb/puIlN1eIYQMZQG3xrM5yl/e0DVnrKTgy5DnAojWYy3iETUs+AmmcWhkRwwWLE6mz0o5a
D9JcDEC+6ILZLjAN44841F+W4sWvmcoo8vpylufmy/sIz54x03BwSo5dOgwYK7pUyJF3ln2V/tjo
abiL0971y3nlxG9nzanA7fV1S2eL9ARdwMO3lXfpsNLRHMHk4m9d2OzbvxI5BEYkLwKs1uSy2LQu
ctlEeEQ8AgfVlwgIB3dt1AIHqqHU3YSEQ9Xn88HaavT+Tm+HWbiFtSB0ppQXeu8xg1G6XykOP9Pu
gn79O+eHCA+R6FwZDqsxm75VObL5V4hACQ5LRxB0pV7uTs7zNAljpyk+tiSWVv7p5eH9Wl/EUDlP
AqqKEpw7SmnQQRtoZdw2TCBasjCIOK5BVrBkm0hpoN9MAF5XqfqeaVckzDFxH5t7mqF3yOBp0X62
+tkstZemEDy0uGfDN26jBn3C1JXjzAvbTUBgqpefUa3dEBtbM0MJhLRiO+/42vsi6dqr4W4bN18p
S3U61L837PICS3wc4XqU8SOdh/j2UW9hnX2BjerQB9zccDdjDauiUTMSFYwUVAlVSOY9RjujJkNj
Q1CKZmaXw/z7jHB7QAuCzjhoe+9lI9Fn3Ga/DxJ4yCtCsEH0p6NKGpVkwOgx56q6E4aJlhLwv5lE
WyCxJf0qTllHWnnWZpQa9YJXf3WcOic90EFYwoEPCNNTZOokClLvGFS0hsYyjOFRWjw/p6wXEcGj
TcNSqzoFXiJJocfQeNSI2oHXeFJ0JzeD1pFzqx4EXhx/KOg04BvgcgJIiDO2SOTVvPcHDrEN+3YH
ukWtBd8B1KtsHUzp7ZGmsNMjnz9Pc7pIN4HLJQgOI/TM/1WCWnOw2OsvnInRL9cWJ6+MK8SKlZNo
AXE/eCtGG3O/YrUPC4GJSPcaHqHNYQFnc+kaSHV3NYgdwLZFZREXNx0pK1LmFRQKCgFZVAwdw2VT
CP/8E7TzagfKgU1SDr6l64qUTnHGVFIgtAzO0UVk8whY0bs78rkcQR5WzZmOSZrg5ygUBz7dSE8s
CCaLwMkdgk5q43M8mcQQTAI2ortmL66K3vkLTPhscjGbDV6bT3kYBzy6/kWX3o77qHQ5t54N3d/d
lvLadB1V1fiA7h6lWNcjWk0C0nwC2izTyjRSCNkb6FYaCMWiI9AFcm9rc+xoonGsc3b+dGAt2Alb
28bm5kBFalWtB0qNju8kYNzIh+zs+4J9+8HT56MG4dk01wJ2i5Sx2WvkOWbyT8+363NtuaGtcoiZ
t0FOIesKdUKTMh+8dBCwPsy+KyHJMDc/LGcsNby7Uh5wNhh0p/arnOC8v95sw34GaWu5m1XCEdX/
L+Qxk4kvYDUdgkdJcOaNOqnZZTHhj+p+1P06FVW5WC12v9VlGBS6mxAC5zinbiR06av/0pEZK3E1
1xlh6vX+OqBg/H5yj1n3JUrhWR3RAgPeBfE3dBibqVYLxY8ssFpZpC0bg/3XutE9UZf92/+Jjirq
3b9HhkjGydFJt3A/2LxjxIn6rSxRcLFFS6jVlrLdYH2k+thm2hvw8Pfm1wuCb02j++EWeE1bUCHV
utDkPVK5eAWnO7+VkErN8W3+2oef32hgW81Wp1Vzn4/ePLwJawl3r6ql71nFCBXp1KtJfIE/kNO3
ou+fvkwcss3KmbOUkjlntdGiTC+NcgzVdkrWq+7C98FBkUxMN1VuMD73pYmdjAoYIdFj8PKCsvrG
dODE5vzYdETJguEa7y7ECIQPjQCLV1m5MzrqeALvvDEutAQgWGFgS4KGKtDz4U1G8Ul3UURGzrxO
3dGCXZAJNSiPUaizZaBIaujZt3eDu4x6zFBLcLUfnUOPMjMMerBbPFEtZkLrUCoDRv5RVe3XPkz7
tVenM0SFDBKtVdL7J63SOeaN/2x02R8DEBYKNfoG/yF9aV4OcjDmw1BJXU7TxCXreDR29Bu++So3
fElLq59mNwJSZFQvTijBDCwsuBFIdU/WVoaWFWHM15xKmeI640e/WxZ8CMV1E0HuHOgciv46QtbR
EC6GOTyKCJshcbyGFUSyDFbxyYo+iub8iAtEzvGS2r98Sy/cAe0J63zNQIrvWTxgqfLBBWkj/wS3
C60rHmmcngp3UE86Eg/XaAEidzKUFtisKHzpJViDQdqR52jsifcTFX99aUSZcdICoiYWZUTFJKKf
L/T8Z7Nho7uP57jzHDD9iiHvlhNXMaosnSRNR528XFFTg1bME82pFsOoCAhSlfoLON4Ncip2Naal
aBesVg0OKep8NWtqyeNc8KA8bHKnoNQqYwHTqo7zAc6JY3pQRg7dxooAhnw9esHwZLqWePLvtL3+
xwWZV8dErQwLOcJYgOcfJQoCNmvy//0ovDjZObRIJ1b4n/XdyyZB40sDIRo1QhkpwMXbzNupxh5Z
XaNq1c6WG0tXIupeh0ybaQ3GvSEMywg1Hc1SRxwmQdGUtJVN2oMB12a6pKJPBOgQWvXb7Aha2x5r
VglymcjTpuBGHF8Gst7SWUOAzMtUxcbM7iZwJfAW6CLeXr/W/0QVtXcgjv97twuo4IFIT6mpiR41
IIcFGLXxB61tepqSNtEmp6m6dFpsIhsVkBszCOSkuGS6XmZZOLWXCO/s/tYfkCHTsnpToKfzrK0b
qcU9G1WOeZHLbuSk4Fs3BmMf/DRv/5ezKYqJWSQkxHB8ZqRnkiwBVcPBqcvKm77RTJv/g6l/yLDr
PvAo3iR5JvgTa7kM19rFJEHoQXEGaIajkVY1TxpjZQabRyxHrgorOawzV/pna9a2xs7oJ4Zo5jkD
Pwzw1rtn65g6SdZA12UgKaNJ/hiDRuZAlQAutkYghkyspcJ1OtXY9ZEHcJRJx54g+zPdiRPpI7VP
m5MyBVtr1hRN5YY/Aobw5HOezn0+SyXk6huDTOEGY8tON/SN8e3CdGTa1IT5l9XwFbfew7lZ3A+H
hB+j8+C6Ak97ZsrQ1C6kUKEKWXeOm13IBeDmlx3uQNXD2CagDffnX+Xk1Z2H1pBFtJz+1AcYS6EQ
bfEFRt9+1V5QYysWV4OuRP4WxHcNsPzLfuIu6SC3zacB9stARbS4Iu1ForStScRTaHyzkMLIoNIU
ZF6HPFH5cQvrth3tCTynPtXQfOeJKPTE8a7Yk/EF8c+BhAKLIMA/KX+Kw7zF0CzguIaZwbAKPdJ4
GvpiVysncGPafKovyARIGZQUS1BnIouu0tfv4ceCqVmi68MNOb/KRw1C3L1f+cJcy6yX1nmFY6No
adr1UhmR3u7xgrN058lsLZOSGRVJhaxBBHJPkW+oyZjPQwvPV801LzDVqKL9HYBVZrYysMTMokf2
OrGk7Xb1pT5YFlSG6/ibW2YCwMPyU2J8qiKoZmOw/b8jcGoIm0PpIzliLWcVPLGsnER7oM0rHcQ4
oEWOZX+o/sSFyRn3ksY78CR7+4lsZZaCeOenhUcyQ1pktOaOMUcs2qsy0odPAC8hAOOpw2FAQOMt
83/CEUN/k3V3a+CNueeKt7aycE1dCltACQ3zBhItoyeftGjE0HyOw5I/jiSqytYnWmyshnQa9W45
c9k5KUvjzsRw9rNlNhyQDcwsgw3NeUGpzPAIyTp0AFcF7aAYwkx8R9GhVooCjaGy9LDFQKn6A+tt
amQECaDVAhP6LZ1Td3QgZFMJg2Gv69cvoLF+WPJ1Y0Ya/AdnmuEmtDlnmLIHeEBjTPL28NpgUHZ8
nAdIqJ+hCRl37TmTxx3lETJuh2Tu0VZd0yqz8PP54/NWULJZTiBleUiBG+PJN24+/sVpW1szGHZF
PPqYkiATAu78+AZ3CMm0LugTqL7FSM4PZbYkCdpSIEi6VG66G6DZsA7Te6sDTQLMSTmpT/SiI7yg
vvqn8wkGrilYkjjcb5oNkc4p2xLEksGzCKWygf2eqHg68B+zC20Q8NRgVD9AY9DaOyUcDDsoKu7j
E0u1GNjWcWv37h+B8VKSvS29vQ64sPz4j7RNarVj0QYHB088uZBXMjuckXGqYKjStVE0MYFwvjmN
k5Hv9Ybj3Nf2kLryQqQ2dg9wAfp6zMPNRbb+R+FvEP43na1f5obIwgPzovB0bV34oBrAPs0/ksJ3
Pp+xsfVwrm2uEQR5hUwpv78wXIms04nCEfsO0ecl7BmMF0S88qCAEULpPGBdptAF0p+in6YVBQTr
tQ5eA4pH/6ZShyOZ+K7Di2fhNSdWXzAFNb3Q2+3ucf8OLvgkntB72RsMApIUGgiRLNyvfDsB7SaJ
37KZa5LZkwDBQ0EBdNwClnHFxy19vWTyNiU+D5a4iPBDgENZzfwhBw4/51YgvMSDCKM51OXTkvhW
zodbP5RlYe2CziKeLbP9thN2g6Ix7kbud81DSCzvJXYDQTTf5JY1qTapVmv0K4MBQyPDfQf2lMW7
46zgF5ajhP00kCMzyiAdJBbxta1vIgvq4puu7FeXCPhaV0FLMTET8KkDMXMUifKD5wWOP1nYPNnu
oGfvy2uYhJc0Hn0XyviM1uGD5LcwdyTddyAPOQ4XfMWdOO9rqeaFOgarW8dAwCKZSc+zfuJ2nSVQ
8l7AQeFA8sY8TQXslV/PxHNfbRbv0PLwigMCuj0oSE7kMwmNO0reNQEmt8/yQd18TDh8ANuog/8c
Plj8X3z1QTucOhdaYdfNAA+D/G3UvpglajvfxzuG4LCV+9gXuyifkrRgfWPLB7JJb9ocMgwkReTB
2FwFuKLoS+FvvEgm3FeDf8C/9LV3uJ8zYvdJu3Eps7mGwrmV7aGC/q6dMNCw/ve91co75pSoEPxc
kA+xLA0LpGQcVx6pD9921G90r4Siam+uyecjO9BrKOtJNnqtxaIAvu61W8v7THL8krgO7qlPpiNo
HtHRQ8/goDneCDv5cd35hhZbcqH+i3lxmMGS1zW1wfBB/6j51bdZFkMLD2rr8QfrGg1RG0DJYBy8
BHgXTyke1fLYv869t4MwLdQnbt2IOR70CWwZipNdWoxZQNpdG3tMurPt22b2rX4pXGFgpQqFABu3
82cHRPgR4EGMERMHkEWOO5FlEFYxaJBQDb0LmmHQDPRslFyEBlrfzFaHhSs5BpymRqrxdmXIbfYL
tRoX5KN85hXVJdOOtmGGslV0zJ8dspy8Vp4EBPgq7ID+qLON+xvEPnAYn9n2YsxbsiT5CO47EkXQ
9Ue3CQ1yy2ZuZQVCZlxAwxl+ZcZaejbONCgy8sA0Mprrzjrgo/vPbHigeDwRV5RPO0bmc4nl76IT
qPlieU0L60mKs/bZPU3kPnpEsxVxpafzLr58Gp1tbfo38LAD6jrtFXtbJQb1Zb8Un3f0YrVPxp/E
tFeMbzQRad/j3rFdJ9MPo1iaItqNsNoxaTLHNLiXBM/WjGufVuPoqMYIvTAsi014vc5Mnhu0RqNR
DkYumTyqB6qGU1de2D13zJr+5aki5ZLwNLEnWCy4PWzmHuvHcqfxZvPxX1cdCJ32+/SkLOniIPqe
Wg7WwuZpN+zFaslqHXiUUQ4xexJsqTORAL+3AfyiPauQbbqTOOVBMH1STg3YfHw6hqMVQtDMQXwk
zzV5iiB7rCTbySWe00IBQ5sFoKmRo+od4pYJW1er/9eU0gLQdMJRJSy3nWkoYPc/vm656V9hASSp
X5Osk6Jm5sbpGGr7Pr8S8WNvY9l2yQ79T5uOA9vySu3Fwg1qDxQ8UmoI4Gc104/PpD96l2EJIglY
nOWPuV2WEvdNXTTxf33N8hDZX5xmFhpnLAio0HsXz3akjfNJcmNFJUZYPxbd9PNtCoC7UtaHTVAj
Khei/4LkZZQhjhlyMg/g65DTkotBYicKbJw8s67Xyp7/WRfMZt4A7POcrQhd5k8oAHAcbFZXf8R8
jmZ6nom1NGHfjUSt9MWqp1sag6wATR96KSvCUYto4L7NGe8WZqVrIx9xtjp8YBw8oNSu7Up3C2sk
9JrbtYuFWxUxLpv8w8qfKovkzXjmerV1HAdh6Gw440M9cH204qQllwExQn0mb+Pj9kBoSi9nnikQ
KRtC6KfXPjdHDwTV3GCULomwEW0387dy+T8BzBqUAHpYX+4rpiuWs+EKXLI9X0+NSQTk7HNAdzrV
68I/ba8rZyVSnYWBklJAAkTtxOkg7mdophfZ3idbf4mbQgEwaTQxovT8+Wfk3DnuwBRQeeJHQQ9j
UQDC6oXjTOS0ySP0I77lm8pkwqnzwNAxVpwPiYi7NzbaSuLYJadbeMy/CBAXT+/xBbXLS4IwY5Lt
MGNMTzWNrEm73HATWUUrrYkmsF4TKMUPB50jCxxKTzYVToEJZqs9BAVFUL0swkWB1zOKh/9QiPkM
kiSFOnb8AqJLQEvS/pE4HgZdWMwY4cAlLAtV03ZhEbBL7P2UV13Xo0czPHGoFRJoNCVYAuXcvxRS
SUVaZPm6KgngziqU/JcZZxqLZXtmuvgLHLQpVenLlYWwlUcDLU3tSmv5MDkVPiG5vWUb6ypioLi/
ENdo2bpOXdW4BOk/mkeu/cNYnFe/E8b9xYs49iwXVzmT6DPHeZwrWPsIEKSMG6DAZGVlj3WjkI34
MJbIONB0uBX02zR+9uDdmTD2nKrsK6OGR1x7quOmbabEOBCH1Y735iQ6MMTCQEgMs8eZosXrsLZx
SW7Bh4F6FgUdEl0rMw4l2nKzFlYWpshCELE9MB0UoEDQd0uZlA/faL84DdlNeep9L800m3Gm/H5L
3Wxpuk1mfpCrCXWvFqQhUNfULy+Anta5N1qTVeVdOulZ3qYGMiovNxQ4mknEE6lNSHCz44ab4hE+
TLiMCNCSweoZAeAtWKHqQHQ5FDLdPO/vqHXlDFOR2t2SaiQAD9zOHgwavnnfY1AjbNJCKDBQ8CMx
QZ6Y0JOOx6QXMssRrmIfLm78jETvh+Eo2wniTMNaX1J0FvhmgH/tVXsOctlfDrgarF+M74BjzVeE
sI1rQVOt/jaFdC0MdQUQ91H1XgtZzqsvH5QtuxIWvgjMuczxfULy/WvzJrR46j5dMZanj1gUMHzO
PYGDOGglW4cC1/Yj5C448MRJzWgMv7eWeZVGdbImVEDVKkOcn02SYm97uOrzLMOXISi/n29nLepE
/Ou39CI0DVpHIj8xp3uT5+VM/BmiJA+TzQEJglIZjVvx5Gio7w09iCrgSTR1O57NY+A7DVojw4eP
eh+HfKxjAVP72+myHfcr6HYvBVwyUkkjoSl1LytDGsjQawEBvBY4of0vGp1OLUiqwjBicmPCtyWM
N4vWJc7qvS89SOBDB/+epnqMhKA7zmwOneRwwAnguNbMhCjjFkP6zBfe//35uneU1cl0jbonW9Rs
lGm3kIWlWtPq5GiNrW8/coeSsr8N2pNG2Nb0GKwLv7czH+lMfYIDhIr6LVOHwFvhEXOUO6N4wXOq
Y1fmiA7nI7Y9hEHjkjgyQWJ7dPsuDNfw884B3AItzwKhxE7fKZrSZgb4f/r480YlbkHJrIRhI4i2
B8NXwVRz9M2rY+3Td286evpBpXpW4Fwx+Y+1mKMQPrhf/CMc1CEqUINe572gO5ImFHob9OOiq4nf
CtgKPpWRqZG2SCpFv9pYx+kZtGjnXKlgryoMcOQB+zJxXulU8I+OSAY1Jzf6FoGdUqG8T+y/eeza
ZwWavj/4+777Vxxgu4R/junTF0vLZ1gNMrc188FJ4Wg1YG9tYKQrbR/kO1M7vOs3GtSi+iNKZPvm
X6uNW7FtzEF3NYPF22YfFSXO6QVa0e4c3lJ2wUd5YjuuWPuntOWfyj6rEmPpMvIOzBmuFagJS0nw
iVQUsuMOo7eIKGIFlD3GSHYx4E3E07UdChgSGjQaI7tYM70v+nGQseTeUlj8WMMDkdjEB0JkYDBQ
W7OfvzJksO+uWpv+dpxIBFJ3YaUuF6sLcRmkbmQotQKudL5Nb+gC2ODOA8Gbv/OaPBOpqlzrQECM
rNsM/NkxkeVf5GzcTeLDFoXPUhjX4GOjGer0IVEh0LHrmPNoG1TBvkTg23hQUPKcwNbOds5Djvza
A1iZmeDZ/F4lIxHvTwhTnqgPAFhERS7p9867z8e6/vdFl3y52SyGW4TVPfvjRe/ou6w/vF9V2YDF
NCMzwhLWdV5XYC/SvIZ4vRBetJqUcOlSxe7bVKC7vS7Z4vAHFNzmlgrJU/8ALRMZ8NeM/a0giIIl
BOaV8l5EQtzWNG3m1sZ1mcs+lU7KVKtnSRZrPLmch+uY5sqNG43sy7tJMQ5BLW1q06NPaOBYDi8b
wNGY/iSCFgYtsUz57rLpRq14SRjmFafqKnIE+MkiyzqVxqfMt+OL+YyEPDS+weuXgTQyWJf3zjTy
ZowuJ4SU0xb0xdH9+CWO5qK5hUBTxJa/u5gigdsu3JqOWTylla/3/AmeWdk04SmmQ3lMc02Vgl/b
Mc+FvgGcTRqkjsoR2PyKOuZvyoQpNXoHt0TFaFNpXera22T90dzIHLq4WxnJmqf529crn0vluDfq
kSqQz8WPcpfFQVTd/2mCTPrLeralkBi/Y9xy/vjuSegxlSR20uGyePwHHbgtgKGfwF/Bhsd4D4fw
YM/NwTrs+mEwQB9V5fXO8eA44xZUkBZm0axqMWriOkxtC7LtSk5SwcoE68esIx3sRdZ3/TTtYmN6
2UYio9NMOwiv3Xbu3NZtpx87AE0KwZ0O4Jh6ZQgtcQwA9HFt8myu164QBxiHRAHKyT9PWg+2KjN7
b2UCaj3+MPanERvSV+ofPQPYebMDLOE96Bg/b3Qr8rJAvmqcbcP+/9BTdix+Vc5JFNhKXvZjOj5j
sre2IInhbHT5RIUB1y7i6wUdQbNLauwQ6gyolmMxfR672ArMSweH6dtmUuqJ5FbdzslFEz7Cxn9G
L/dt96Vz3prytxJmUHVjnNynWHRtS5BJlluk4IrsuaCdBwJpFiJxfocu6IlAoLv2l5V2IMex0eGD
c9tOTkQ+wGuIexOCRbiO6Wwa2ercm9fd8G024t9KerXy0XP5fmzodHF8DQngLraWcMO2sWIVGEAI
VvR0kzOjSmrAgHMFluJeQeGIixYTr/Wy1sEtDw8H9h4MCNsS+507P/sXsQ5ZG/P/JoDGD645CIx8
OZ2YD6cUYe9hR6O5c411Um8iPb2AUl40EfIUKM3dGdIPgh3SxU9+d3sZrIv2ZVu/XL1mk3xWr99d
ebdkFLR9JRy2H919S1sZ9M3b6AIDwy43BPWLXCs53mKp5hMY7HKuBJnjMDTXUIXO9EPn6vH44n8M
qVSIWGW0WOCVl0AQZRL64bZ8mvClqdksbSUmPsrI5n7N8wPujP9jTlk/0MhYsYnqleD/1szcVZrp
mwVSL4Ghl44hlv5eneLrxQuw4Q0SwUagtwKCGPG0elXGDUlVae7UCv/tRbVLkGk2qGcbIWKMiVkd
JQpHJpU8n6UOkAVs9+ReAqxA6Rjix8E8S3DRa7nwAbJyb7QeDfnKWISrdP7Jw1jRKYEXGxjxQFD+
3+6bkQCVcUC5N5ZZkF4Ig9bbS1Ldm24QgIKUDkB9JOHtzwmJzjFG7ntQ6q7vbKZJyOvJ/vd5xiRY
6PLmeQQrSJzRGkrNAQdabEgULfEMl8GLLx3YEAxz6UpvbRpBsa6NOQ51W2GaIlnudXPT2QtdtUMn
Ssr/yYvF+9kXEz7gOIc9k+nQ0M5H7ynse+zEArm3HS96vtH1i9+9iiuOsmP4kBZsTuPuMbLSwNo1
4w0qIffXJtC9yqO42NvQDMsmzy5SbiUvKOeHkr0/T0p2TF1CGvo6bUM6z39ZVZlHIWsqy1pHYm+2
26n6yD/WjrLWicchYCNKPdscShClS/5SBZSs+LeU2TsObHdVXaXH9WN1K6/FeqrYCm/peXuW9I50
9/Ea5+W69QIIuLtNiCYP0VGXkTtxwrjKQ+by8JGR7PfiZ2WiAMU7wNW7RukzitJ1GNleaaKXQZ+s
lYdlz+veBUgB8yWf3q4u408Y+oFNVw13G7w0+LAM1qh+yqe1hzkxijTc29wrsPTzNIqC6ERcC/9A
PqPaOZukvvFdIMcgxGVJCjczudv7TmyhL4hb03gHOSFKyL29qzztsCxxF42w0H/yH0BkgDY2HIpJ
bxFj97T1mR0sS32q2ZvPrOvjmO6jk4XZrIBlcKSDmCmTJgcFxTQJHSUcPJYeJgtSapGuq9GDcsuC
1CgGR165FlxOyLXViCFxSJP7Ado8ZQzTqRZoNuC0NcZGMYvJEdMbPIzqJ81vpoATE2ZUOutq2KMw
KfKvsiiyhzc6Pa9d6xW3CU7wz4D8743H3BsBAdfm3npWlhF5NYCj/0/pQ1RWsjI/QyxrknX5SbJy
Wjb9O/3qf+PTtc9I+dvltLllJw5mu8N4AeV/HRFqyKNn6L10a77NrG23bkOxsixgPLTm53y4Stxq
b5DuVBrc+MPmrqZhjrVGdLp093f8GUrXJzp/79RH2sclJswHVEedZ8AQw0hr1tSe0OGQX9C9Dynh
mMKUFh6AJ2Fesvg59keaLbt8Ow57sqXyGys/dWH+mTx9hwz6v8D90ovhu8HGlskKY98G5dINfSUx
+fVxQUNtgduDGTUVP7roRiRwsW+1OkkOekZDR7D0eI/yntyAiodyN473w+8gdtBF/GcomIxEohCr
tD8yubfIBXQdTOOSPAwEnoI2qnBjttWMh6q0Y6sLw858ehOZAN/c0AOHkV7vStWU7qh9TXzfHQs8
RXhKTxiN7gPEisl2OROA5YzRgFJ52sM5EBIT0w38BqDiqrciMLOwd5CQTZj/drwJpG0USZq6hH/t
Xx85VobEXz1BinqEPEcOYMHMAEYi8S1YauSE6XTo5xCONM3F2s0fX4ZSm/Y/gJeZjdjuWy322otu
sf2VE4qPcasqFUjlZK1zsAYWjWbFXKE+wELtjD4oV71hYNTfK8EAzC7V77iSPYMMJ8J/RRo63Ifq
T0YKDfugqjB/kjZX6Nym/T/cjSVTJbQUBkaCCAtezo9S4Yk1MBeyF7CvuLxcOKufGfKNXlEEp3CK
p1j6KaDunARPTGKYcj33Y0Y7ftOU5tfUCSANJhrcYgdWbmEEI11BB3GZuwvO0tVj5O6FsQIP5Yne
pv5OwWi90URETTg7sLLdUgnezpNmKRMm7tpPBFRVqb5a65Qd/PWwOjVxff3USbcN0NlRHGu62Noe
cecrGFiDlsu660HFWLvj0OuFpALW9jdlK1iwXxqCVMrClWf2M9gPf+KDpbGccbrUN3gEGA3kc7Ph
JypAKh3L92xM22DXl9ocHYVny51IOlvmodz81OcorB2tTkKYA+9aB5fGvX+e2MSy4J/bI2xDRHDR
hQy7YNI5c7CG8d/R3HtDiLtYwNIMXYCppB+JlfaWQlGrZ3CIQcqLQaUpI+J8uC7dvOjiENLUtbFI
6DnvImglQyMUNdG/wJrnI8g4QbR1ZMXDnq5Yj7bqwXcbXoZtxarkLskI83vbEp15xzo5jcrG5mLx
1VBDQIB0hmxjnu7TVKbhJKjP4WC52R4RPwb3cZ0lJxdFRjAUmUgRZ3lHK8cTWbNCZfJTRl6kNNdX
FGuLUm9jqulntgVC2pTbrn2tXRYfYN9IgXtkhHIVUe6zk/JGe9BELqc5S4uHl910gttasAZzm1Rx
lNmmUf57sXXsMRlz2qS5cajHvnE2HtbjU1IfNm/ylnVBBO5ncprZfms4VIB3KTgDqFKUvUO1xd1u
iYPBgC/jU43MKdGP2KQ4hZBmbjGx+gzpfoIPzX6cxmq72zZOJOrY1dLFCckMK7+R+gtY7YmQNEVx
Mq8501SpB2UAuP1OHPdVMwJFWQqor2ur94DPPe9qTZFEOzaO4Dtt/8zAcjDYJcd3NT3XzQrCSajt
9zrDJ+CyIuGdWUEaw9bFdpZuKbVKy/RO/JK09BU69fSYJ+oU+p4H/XXBVrLgNsLGHGU4sKX6ny0K
vb7P4ZGSrMvexwRapeb/och8+CSnVJqNydjS3+OYkqcv7FECF++piYv0EtdYWoJzvLvI7hGLEG1b
2wU53H+5MjGT7aDDrp7frA9tzCPWDC4J2wcugstuALsk3/YXXJZ8NSUSA+6UjtK8MgXxfHi5S8VK
06jEkJXWdaGIyXuvhB54Aka7FdG4Uhs7ysUjeoW7WxAv1byCzKm6Des6cWOy7TiYpH5KjNHNfdRk
G3BsnLIoIDeAdi8Mrq26rC3bT7Cl93Q0IxlZA+dh/yoe+7Nasw42Kcg29oHI/bYBERqWXX/xkI9P
VAePq3sOsJnAxRcD1CAuHlJzq1jAN9yD2Wkp8kAmPnBkuE+qqSt35h43Ri5+kD0vnzudrktoQxnL
2x6aoElsiTR5x9IdBkCATGYGf5EReJxyjvIw0DSgqqLRrK8cDh5ycyQbjGbWlnx7yAhxWBdrEogT
aDVWuZM3E14Ei7qf1jKlYcRiG8Rpce+DQrItSnoJz2F4ZtCESmLr0DfyOumDbtPsunm96JHKu4Bo
84UbBZGoh3rJA+oNgfwF9yovATkjXhgqaxgeNManZ7pztUOvJjz8c/7C/sP6iNJrPayYnZM83lWi
TVEuEqedVAtzhkEAhW2HAR9kISkXuzTE36cyKk00zogn5p2fTMhyQKUd/sxxhJw16dsObd87hG/2
Z/yqgaZdXjVT5HZVv4Ss4K6P1gpGTEH93UvLLo6Iqx9hpnVl0bXTDMdtriFZ2xBD/nOeKAK6pP5I
TNNmKGk6rObYCj3qmCTGJjyJtEgmazco8+4S9jjax5TMj57y9E1ZxGZd7AGIVjHczCAx+N2pPU5H
JOpwW/INKRKWZpdL00ocQLuAYsGiyI7KGuz6HauI4mwyJ9DLsii1nbV5SO76UQZbRrYulNTRbKVg
tYigUktNEL75vW5CPgu8h14nq64wRIrcPP0/lQJNecbRpVPi24O/I6KUge0G3bnfuvTVNMjqfBDl
Wp/lyua0Lf2VzRQX+7JQlf7gUvN7vgJxanW6dJtPOZyUjnrqSBAaOMs7wwV072t58cMtEwovpBze
VUZqj8J1vQHk1dr8y5oTKk+ot2NgYuJM/hwQAvD4adpawdvDFEOzzh/qsOLLY4cGsEQCicLsNXyz
fBxLjPx47ZLRE1Y60o7Ec25+DwN31gH6CT37tvK0hkCdQXc3/itbnFWn5IqAZCntQkrSky/QVlmR
Q4jKLKciQ6AWuaXeYbAW2DVt+wxMlZ8ZWzbR4DF/A2jBM5mryBuSsFFhiz6+3fOi48Qn2Brcxwwf
taAs+TktxwdTLu/q5BlctmAMyW4a0JZmSror2/loANOteGUzSRmYm5Ez/CjX78K81tC8/jfvjXGZ
/6dXKaxAnjJVU72jwTGSdFAUn/709tok2oC3eODkKmCRAut2QASSMtsjVUkSvhqkCQf9PeLHn2oJ
BQYVocJMcExtUJIOnr6J+qG251pXybkJdfVoh40q8ce6g2qe62gz7fNoRwfCFDZ26F1rf70wYYUN
I8xdDTKkhE70RZL/EGdEerXyrEBg1sGVOlQ4pKNDvGYvCBP/YyJ0JmC1RmffJQtMcgNmAwnkoU1b
d3KJxvKYbPNZ97K9jBv8YwBM6DEmb3o27JhGPl4ptUWLTwvt2BNYFQg+e+AcAgpzzC/LNQNQkMfD
bAz7Uz3GwquL1sPujm3fOMuRrWJRjA7u6b41wROi4R+ehE5fMadW6j418Oe6n6euRrzb1mo5NIrU
kAEZZB218j2MKPsQUw9r9mgHD23KHROm5S4aXKoR1qDY3U3irlPGDOZ772tk7DhqdM80kPnsXwV+
sxYi/mV7S5R/6nHkK1kFIXU2NNE1dP6R7V7JGoOYYYX88PrdxOWNQ/k0osIpI+Hq9tuyhSZd02ZA
PVGwamzGNGx11OPsHX0LgrLt1LQXKNWUyOR2Jx5/yCYJGgfISYy2ON0HWyEMX4yUFR/+5OK4O6IR
NNZBd3y8a1tQFms6sMA4v1/olCa7urylGWHNtsZzEzGc3QX4+INpkaUaqZ4erIKl19VD6ZjUL1w+
huJTTYv4YK/Mh2L35+OfQbqNgJwy2FwebTtpEZKC1SABl0tfpwB7kCoMbqqdCgsOPZY/EySlps7w
Ze5+JhuM6uA+HJLfNiJJjzR53JA7G0fVTr5kJaFhqU5UT+yIBPLFe4D7hcAL1Zaslx5yf6VHqIsq
n7K2++7dJvt1uKEnva+WWI9JnUl8ZJs5hxceLqRgLCgyI5+kcw7wupruCIxBUANfrMXuz0f01MeU
dlkriAmvtEBz1Tzf3hG+StDUbAb+oYyD0vcyI9722fwfuQoJcxTy/1RBWqPISUJ5R6VrgEF+7t4w
/CwB2+7DJS3YZhGLz3jbHjRQQ3ADyd11yQQWBqxYj64G0JVeGl40MpQhl36Tk5Xc+uswfuMTe25j
YaxHPaz83CRdm0J9LSeCoe+84lWFqHja4qI+WuV8HsGmLqgcHcfB91AtPyHZi3ObDBp1V34mKHxJ
jqiXiF0RPV28xT5erODb3rESyE8eV7VQnmi2uEL60Ae30L36xbWZbjQCOkmrjRPZHbSpJ+lVP0kf
Hw7rMsk3DbVcCfV6ZIrgBoIjdWfUSGfeHgxT3MkA2xCjtMA15vxQ1vyCOlN2PG+PpmzMJhsEvnkW
F7mebvXxpowctfW1rXRj2rKR40Cg67tssdWXGoNO815WfNPHLZVtWNhqkRltgp4T7oaZzSNTxkmL
6MPlliMdlgIXAvJIzT1iKXbe8nXvy0NTH8kJstNypD9ViEnjj4KLXDaD0KTOW40RbUapjni5g6tV
8Ei49GFQwVGaOnblKbTKtqD3JqRVnW2UOZdRC6u2WWmHR82NYzd9ewPjEKJsBg8HP6a7+Zyh/fCs
8bhrmA2QLPkZFQVhzaNJ3xSdFCPhx5MG90btYwKRsw3BRl0Udg8tKx5S1RCiFPIuuuQRiIs+NK3z
spyO+KQiOwlZHJ6ckeiaH+W5sCZcB5nY26cjGg/4c2hklYFVo31RVVOYg1DFzBga5MwzCPqPyV6r
bz7s4Gg+vqM4N21rxgAaBDtWC/IXsLlPGgyuLPPyhXdlfo7grziFpfWd9txTl4vSk142nBugPH62
Nv1FZobR/A0pGxokRtPJ0CqoyGzVGiDtCXTltAVBmJQRCKsqkeELliZeaUGcVTZOeNt5WMy+cDTl
AkP1nHtDD4klPlx3ko4xEtmepN0DXxWfWIcoYVEtGbV2wUTquZADpVCcXEO3AElw0cDXdxgDmYxS
fqIoiXRSbP35mUK+C3RpUAGJwaTs1wfgiJInpvfGQVevHCbO2Djnn4LR/CkZKSzWNWMso2ZaFO4k
Wo3A3Q0OMcVI6IuzhCmraziGMuuPmOt/AhxPFfOl1DfjaX5du8G3g6y7uFv3roDxw963HLD7iv5Y
Ld6ZX71L63E2TeBeENvgTS9miG/VXyDPEBXBixTJ5goUZJxX8wuYm2KRf+TphQgTY4qVXEA9QraM
/BEPKBk5Yll90erZ2QKjstdaCuo5BX3L8JwloknRltWPD/MP8qaFfRSbL6/5Y6ZGBkN9VgrOgkgI
rWKhAdyUuB1hdGCbRDpjeIOShk/mGs3pmAFcE+nSLW5J0porS2lOfVNm+VX9idpckvjFMwpGtAvb
b5J8yj9G7meKLsv4MgvK59/pYrbdb26mNScccYNfl99sJ6rfLFBkJ/CGP669MZeJfUNYEGzy+BNZ
L4TFyEqHn9YqTPcdxrzjAuxD5SQsU/tjeO1nsrYr8YWixSxpvZQY0G95QuODf4NzMxMb8eGf/7Hy
BQ0K2FdZJpqBmOntrPBEsDElrSzN/ZMEokMN1gEz7oW732GfRKee1PHrAfrqgQ562yB1YYWZusfG
cqleD35WxEiSppoOaXVAdRFyO/cRSzIHoQ/1jYPGuojLSocJeOFSHT9MOUtJyVokTady6cWFTwNK
q0QybhHkUJidbH6DFZ+OXzm4mDusE6tMK7yTYxGHnrq0u23E9qB7iUjffY77bEtWg5smhI9oyjAq
J3RhADmAT6Ibt7VmXRe5ObxU16UwxtKOigDq9/ggn5PX2wYkfVlNR2tMpxr4r0/ZbXAkaSi7eng/
oHiNmMQlRBaywuXw/fh2iRO8hSszkUI4i9ZaFjXO0TNfO9pFGzbHeevVRC+rbb3mFPHGMjaW8y6J
VNBS9Y0z/eSJisbZTaKhEyDt7wCmJVey2bf6vcosqy6Xj76XHXJ4vd5yuJd0IdD6RS99gXrPOaXp
fpMhkezu/YgwxiNqsDMFBP51Rru3+li4BfoSIOiPgs7bATlJ2QLmxOst8E4jChU2bwkugDie9Use
6AfOWRE/QzGKqK5yRnwYGpNnPEgov7qmH7SKJzpLe8M1L+CsFvzNbiKezwzInSTEdv/sWa8xIkTs
GeRpWlqZ7vH2RWJ/0NXFSYOlYqV1yxzca52tCbb6rpy+9j/UD2OBlMpsZrVEeb0LAGw8b9lcam05
kJ7zw2DTqfVDIETHO/D6Z1uHsmZM6rSn22rOz9gewz/4ORvOq/wNYYTuYx//MxX9XiBYEmQIjCru
hvRcEWwYELq6glURRcalDnf2a6r38E8bLcRDt7h724U7aN2IMD7EpygIGHtNlaC/O6Rsere0qo2A
NEgZBmWm5hRbWnvmzzeR/Ht5HM4hwiOSPhfpyH/269mlFKNfdRGFjx+uxDKth1jZW//4C6nNWrjk
1XfFrrUJy1Oihbz9OpUK9XE6Egm2e4fbL64nJgxnbehqfxAaX0gUgttCeBaCM2F5vgqcc0UcZQg4
SxaKWRjHNs7xRwNlLliPknBKGrOqBcM7CUyuoenOPGEUvvpQ4WUiyJJj0heW8DG7bDpXs58DDLXN
qY1VsbSRU705KCoQfmxD5OpBnJc+kAIjxEG+ug7iwEncIAaF5pAEF03WyNmogjQiY+qyrM33uSfj
3lbul9ZynOi8/3zzS20jMstnTD7Hx1akfjK0Wx2uNGQTQcnDNBggJt55hW1VRcXXgzoGBMxH9a1v
6QHNuOXbJvCkMLiNbtOKh1fdN3pE1Io3U3Pb+t/fdrqe4UmjmjvNJcrR1+dWuHLZztKu6vlKWpGb
mR84l9PNDL3dEnAprig6hPIdUVpNv3llkDvfH8tBu4new4o+zEz3J0neNWB1/kRUdsgFmQjKvjgh
ivjlje1NeGeomuzTbIUrEYeEJ27e5K0DhhVKAMX8t3SKVc7c8rYSXbS8Z1dBDzcEG6gvLgtXfFAN
gEF6x8fo9+VzYp+Y0/AIgRn/wTXl89ZSKWg/hHujHPFFNlPXP7W/29Sm8JPjr0j7n1PS7VEMCUJ3
09nUG5XZcma/4C067fBiTNcwmDCbKjOhQ3OXMwv5WqNP1KxcGctk14RS81UZE7NcHF3mXH3RRAbZ
wog9b+sI3Fc390By3AJd1pFH9o/JlGqGqX46qo5rO3db1uepMiHIbj0goQ9F2LVEg6yp1VyU/Sg9
TvtbHQ6YvsLALjG4Z/NRthqIwWl288+kfPp+aD+kkNy8KpwsoEl9BS/19BEwIX3Hl91kP5v5f2hk
mfQ60Rpl87OkET/sXMxEiaC4fJgH7SrW5XPQqjrQbQEnqeulbi8AnmjLt1zankyHOI3efRCdW6Qy
FkuHnEbzD/urQvthWja0xJMyG6t29n9FV9auAfgfnOiG4sQkRxI2WKMJdHNW2Bj7Pa4Ch+w3DUMt
a4mharxTzUzfoauyjp7g/om6EsHjjFp2tfZdL5eygidSlUUmoLxjKPqXsXLDufGzVR7reqDZrXWj
fAmaRrnUUazPSwPEXGtd5G2oV83pdu3Z3/n4GjQpZviclF14od+Xqyq2dv6XjxE+27ZY9TTEJQzS
ePX+PKulwEpRkBkH+y7oK8qnva0/fPjn6iP3tRXmribk36vmHWzlir0scafmUf9A/hdJpZybmbS8
MbZ+Qp0zlPbun+bQrKCtKXJEbDQPUhKpUVowrcGkDWKvdmcaBnDXIHD4dehDRqtHOS4Obg47WcEU
HNvGQanfQDlGxTstnwaX2VC5ezG1Zl+0YCul3eP7z6e8o+Ko/ouqJkeIUgq0wFycUgtfDKa5LSOf
poExEGIWH46MhlXrUQn7iGBEBcU/vnXC9rZlCuxL39r81SFcXtfX9tprnKUdLeD3LEMaDF1/nEla
vQxttOM11DoAwyTTuzCnSmk+buGb4oQV2/vOt7ZxIspDUHLzGemXcYXq50lwJUjm6s+h0L82/bJN
bVo4G+ZcjcqkC2QMWoIDTfyltZ0+U0biaaMHvbVPV9EIJ4BCVEL9rqPk6WszM7X3AcKqJfJRu1j7
UPv+NKtazNmHL4c2deW8lLRdYPEiv61Dn6fpge3Jjw2zELO2hAYSHV8VSMwiG5S8AIZxm+6Q5AFr
pxNtVeUPUS/Y7MKsos1qXeEvxwTo9sUU2n/kDvwu08JRTp5+CFZ2z82q97ykzKR/N72/BO9q95ml
l4pj3eTYRXe+aNCGvY/b+JMgy0i7hnFgVoilwDtpA/gLP/lruh+n9ZvGt+MnQc+AmOulO0Bla9Nl
rqL8D+g8II9mtizgbGmjXgQr5TJRNbpGXuEgSH1+AVSKY6cWUR7/ZwctsSfS0m3PA8Tu6Ysm/xX6
9CvzMxsk6A0T/sJjjIpYvfKG11tvzSy8VSA9GUY3D/hXinNyQ6ghv2gpXfjyu3B5pMn9KxxInOXx
I03xbxIo8oqpMH+83m0fliO+bRjudDtX9F7NJZiSMIu3BaXbWaPDQDMGwaUl6SkKz5hhTAtR6CWe
+yDfSuNb0qb4oez6emfScFn3dAvLWsx4drzf//Pwl9EN62m4oO3cPVrKofDuF7WWB9xuPwXT+ewt
AgA/a5rUqZCfeQce6JeBIVIWB5NWBU09osBUzqFHIsVu6c3RTtyTk48vVIj7mdTqcdkrtJckYEeI
4HRdqcFOOn8/SAVCLvXDe4cDhO/Ais7BuFVhlvekkVkSdqbn9huF7ytvMnSWuyh5yfHRVpSo9nGN
jh1tOZ6rAFLGhqaAU09KRS35SA7xw1W4lzQiScwKOWJ6ey6Nfn5q9WxkQrhGzlJZu1itQrFAU7R6
UVWizR8OfvPlvdRMYQ==
`protect end_protected

