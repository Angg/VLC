

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
DNkSCrKrSZZGZ7V5MEC0Sa+FIa8Gkzj+o/6NpxIyEzT1r0pebmEX5gzn4ZglnkddvJ8/1f149Df6
ndMlnzvmbA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
W3TEk2OoVAEcY9sACr8qvdTXcz4KMrr0wBUYfTJiYRXEKj2r9L+Frj5vlPoRfXyR8BXMuNIvntP/
hRtRCfRyewmxrXe1oHJIEkJM8D6eCjNM+zuIptS0mt/AsnOv+MMQLDkTVqLaJNUJXubQtL+dhzzd
RD9SIj/ZMKv/oOZJjHU=


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
2wWKJdgoqz3pSafJq9a67M/dd2FxPncTZHCUPF6InCTgFQ7MOQlzLhplRl102JxCos5KzhVt25al
HkjLSxu9PHw1ru871OGKgua1sS3EafdVjGCdT5iL+6+M9XT4bQzC8cVlky4YWr6qOy3G0Bl3zGGA
4U8j4LRDtMi3U1kOYa0=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Kxq1/5UngNEJdxzilglpkl2MQX9t6W7lRQYEeATFLTlsFzdBmcbPaM4E6/H6jb3hTjltHCzXXzJL
yu68g88g81H7vk+zIgG9p+bAH5mVTWnGpTcQ9Nq3V+BFNfatOquArwL5wvfxgYh4qmnz5LLzO8Vn
ZipCR6RyJHvmX3LECK4ZGhdOjgqLTbHPcqhN/bNhl+BKCVrOY8qTWY6WSJt2I/pR5hbR+Gxpp0v1
fzycz6IA1AnyF4dzdl4sorgs97DN/Rwyy5DX+iGMZoJWJSj+jKc0DU3coqqjuApwjmgaPZEOIkHt
fmd8I93zHpUVO+LU0o2VXdLy/rhhX4k5zyqLIQ==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
MMro34sbMT/dSBUUDKeWGj+AS/ioQgVbGWAXG3XMUY+tNHQekxt+oKRBWcwquBl3sw3SJLbR1Rnx
TjJ2MDDzEH5uCz1vX7jZaQbMCFAU3K7MBn40b87mRKYgK2nBkQ63tKhSjfklMsYEEkc5/qUdspSU
GIdrS3bVjN2jI60HeE4r8Ae7725zNCxoNO7hmmiicY8i9qwR3Jx3RLeEISc/SwYIBg0patrQcspa
o2nUblqCyHtuSc/DkaBV68tb1S3LDYROKbnkmBVtPajoK0FwTW/5ES6DuetOb0ujYKX5ZJWNoJr0
DsAiVxbKY23jSFr7uskYGQGx1K/crFks1SMEuQ==


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
DXzksdzpRyBvPJAO8RW4ZhlhoWO1yMLSwz3BzpxXSQKUFJz2DfYgIojvnKP+h4SEWOeOMQNr+agZ
sZh5CyJzK3n38AYVr+qSmIrSxy//25NZBDMRWM06jl3lxtySkqX1u9lRJvnZzDG3hVY4BI+zv+3m
Uys3/UlD6y6GV0iCZqSqOjNMRk77t+OnDh3CxzRxxv1qIqIA3AkY4LV1fP5qMWjFIYo2yfPwXZ31
leLLHOibckzEYHfpK61VUGsfYsK/Omf6e+sJIk4DfwW7z+qr59Fv/xjUYitqPxa99lpT0eMUcAbZ
NbV6OJqwWXo35ZdTdYOXEUb32x+tBF6ayvy+zg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10944)
`protect data_block
6+ZT5N3qKm2jjMRLDB8m3IOAjae3bOkPJKmi/b+b+SwI8QbTIHiI6XqKHlhul6E8da0sj4o1eTkY
2mKsKl0qWYrhm+uUrdXxWLavXGU56f9rRDN2jodob5VNnaDO8N+7NpmZEP2GTyrLHwUfuAaTd8hB
vAwwzMAxrqTN++gY7AirZz7b7+Q/QKZ4w54B2pBf1UqskBmWhPJdKYi7eNc9/ex86RYcduVAAa8z
Ek1ckTUOvq8l41j0J4MfUsmFKJORdpTcOCtMr06ye7As0N1/zr3p2K88zO9W9WUrCqulszZQpG8n
nwGdQaBPb5pjPwBIRvCZBxClBmqdkxRFpwGN+rZB6ahLYQ3y/VZ3iVCKXMf14VwvZJpkzs2j14Hf
flXtMSgzdhNdx730AH8BQuCb9O5/ZA2gXuhl7VHmYVfmwc016xJwd6duLKUOiI0+oua2N9rOZnPc
qvc0o+9Q8Q91KuZk+bWI+KLSXeB5XBi28wb6kvTz2TFc7MOgku250+mt9ph603gUxxGKq3ctbMb6
miDP31NnMAr0JSAWKmWW89JMsIcBJ+s065KGTPjUHrUZrIQp/elOnUe8kEOgGdDCbWsgyT5ufFgD
nX9ybJQjmvWil6BdVr5JDItGvWIGeUYVF8U8bTM1z/X9gTpvTSxIqhk/7IyQevLGL7nTl9m2mtlG
hFLlACOW8O+KDJFQacFkWRjeM6eQ4vkNKMC0q/ath+R6UHFwb8bDjWlO2T7p/NcF5uetMMoFz+4k
xeevhlaU4TUt3y/yc1swPTRP3F69iJyUT++aMWk3a6ZI1XfQosYEKQcAe0Am2KZQqOw0zZnS5v4p
EOAOqwM01aU8gHHlXXrtKIWMUrh/2XL/dS64Rav9QfHWSh0bpm6GAy0hfQRwzNo+gA0YCUsRmIHH
htxiMaPDxNJi9Pz7TVwruP0Am9+alQOF0Usg2swC+gwnVMsmkOuTghtU/UlQ/IKbaNt9OZ6CiOf1
+RpbenqXbpLSIQqDxBU+sQROR33eNVcP10a8XtCf+c7d2oopyfJOM1GFdI8bkOcozW8US7jM8nGX
dNBBmMS+ukVvEZInYH0KnbrsnTia1cdrgwO++kTXp1xznKCEsgUeiyfNTDYp4wu5guGXKqpVqabb
BFt6SXeAcCr1kMY0HoKBuP+yg0Ll5xzZyTaFZULcNAPA3TyZru7OwMEMyzh6JIfhZRU1LqKyqtJH
TMLZ2srEW+s8v1nr8x+e2xL2G0cFe9Ali/it5GY0LQ1w70HeblBbKnSfNMVt1Qnn9hb700aE+2G8
2NA4IpZIQedz0ai8Gt+vsTbint0GglSWGzy1hwWB5VsICe+dX9rkVjq0UcQSF6U7rCy105YerVjC
5gQ9Ov6bAzuJkol6Msw5TbYVRIhOFT27PoaoCcs0qcj7buaO7XzcPUdmzgmcjTYywyapUF3g1746
lqwgeL4MmB6pb2J3zm9CGsFZ7p8a2l2+FgGuRuTkrC+gH+QJ2OhQZ1s1fUJfmuWKZKKpCGtesBcu
Y5JxpEssXjxJmSZEy1O/se4xIRCc9FZrJ3yLdzPnMtWajOobTaoOM4rXrwLqY3evusAzed3EdaOs
r7bcSHuIfujTNGWnWnLmHtWC4b6fNcQDRGFhSh7SAUvmfn6/WgODiQV73JUwd1nYa0w7DaJOpFO3
JJ9SRMYVLXRbN3fckuqIiy+qBSnfbMrK4B3/epeBA0GMf5jRe7qFd91tP8mvjGC/b8tOWjEd6wJg
D8V+mNkTBc8WbD8nX51dgFlSJn2JbC62qkT6jAIO2H84B6R6gKWk6JLAbhhCCvM6INoHUAoX0lxD
pgWwFZp3AriuQdpqCF1NDRiZdnWqn0QNLZm9ygklrjZBtMxc9ej0xx7G9TS07GhAjY8r1WEWiIwA
HgJnABoJfuFQCHAQhBVT/AmvfcIKFwm4P9/fwgN/yUehD753FXZBEJ+C0vNvG6TCgC3dwbElsn+S
ga1PmrF5NPYkKmuIDqDgy2oaL7Cr1vNaV7WEtA0em9l34l2awAmdi5Q7lulxyRkBa51YG4tU1D6/
TJvAQ9IfBEHGeS+E6aJCM7W4ULJ+pzgY8KtwsElm1L7RQ16CAF6s2R9zV+uFdsPiBJ9qbcm/mPvN
GHmWPhwGA3EPVIc5nbR0VG+7CCQYWJc9YNazeSbhZ9q7eC3quqAYTTR2tKl/L64F9Ivy18b6uMff
M5gLX4ukr5aMd8OwzXuVeKm73hDoDb61cMGF20+6BS2WTLvocZ4BGfUZVzwAcGqX1H160VUEaqtV
zO/z+ElVrRAj2N36fWi1IAQdK447f8Ec7SYQ1/MhBEmlcUyvV4UytJA5/ATRiCWbktSN3oTayqXw
3fygI7pcVIQfc1gNwyg/RXyHjEVwIAkaKUaRGJu+3T1nz2i7+43CIYPz4Yd8HWQPulx9JZgoitjB
VbVsWWHXdd51pTO9cegvDaH7QIYVPz3N2481pLqMztDxCnfJmAuWOOxs/f+hTjxLSJoJGm12bTh9
mUgqKAxltKxUa8SiA28nNiDU8LAK2+rREyR0nzWidVH8YVow3BkO2W1pg9Fsu4yyF3C/p+GtJfIM
QwAyRcDv94UvxgI5AzQsdqp7ptvKu18Ov1K1UIads90+KLRn4b1O3lhTAcfXYl3h/HYawdCKvzYr
XsXbfmxKbBdu2MeRo/fp5radGA4gJN2rYGmlAOSMyBWVHXrcxh8wo6W2G1RQhx+vZ0XV7dWPQNnz
V01km9vkktLFPs3LagEVULTYA934suSAhGWsaAombRFZrmtTzLPPoFr1SV0JPeWTVYth+RJXTEPm
PI0LAGX+zKpulkMxh/KsIo7tEelEgwmox/R5vhXsyJfiiNVR10V01LsqC/0Cqa65/CVXU5jf5b6O
tsuyMweSRoY6EgpVGUluX9TqDiKV1cbwSxWBKPgXEC3N3d+AZrceUA63KwsvChLrapW4JBXzixOM
V5PffftOqdtTblCOQHgKdZu45PhQ8cBV8y/0g1NiPxBdtj5uBDbRBDWNMkHcwRV9xSWUay8Lo9cA
9PlzoXmeIy+M90CgGrF7SRhn5Sm1DdFShDCX9DhD/WfG7qnN64Y6sT6/8MK4sSkvaFBqsxq2pbCW
trhU60Kad+7zxcJIMnetSylUQazN2oX7Zn56xijK7tTIIk9QtJNI53E3Uwfmj6PdiHcrIsEvcZck
tFCbayquGdxBZqnQcj6Rw2FD6cOePS5cRUVFm0elnQQV3va/xmt2X4IKqN3AEm3Xs5VLgvhF5Evp
+m8KYwLd6kMeH4Lck4UrO896xGfRZ21dQXmUvZMNkSk441eWlBsLP1NL5znm09P1VCUFp4wmfALb
OGZAa9h7qtOrOKSfV7RaJ1IFK/p4RPmmaYZm60YMrM90AZSMfyoUYDokFUOSRWlSZUMGLL5BhdZL
T0vGxzOARKpeBFweKqUE0eer5LFRwgOO5tZdpcXm8Qn/EDCAMIor89Fp24nPsCBhBlALTesS/kSj
3Kgi59Xp6c3RbASFwEFJrLIR5oojh7j7FkJFUCoggEDMM73tpdABdNe0BQJRzvlaBLk2j6r+ipjs
4jNNyYYPJVx3lerl05lBaalFe3VvDyD5em2Vzr1Zih2ADaPLOXkcx3wI4Gxss746jJj5UMLjwCya
PciFOrsdBlW3Qjh8UNzAEpbcZa1Wbvnf5WBBnt8xyn6Ogx5JRleQATvTGAVnZvfFyXYIvL08kYiz
1EZmP+GyDxXC6pgP95xyNg55RTsjLRmDo1eTa9cdEYKwJeblsM5Z0oFo4MdbGhJWyd4mgVat7XI0
HM9vBUvwNxa1ji/Kv9tHnWuHVVcLnDq9Dnx7nXO5gWzOFbsAz5uoektQlrUrym5Aefwp+QR9ny24
VfDWxCvZWuVWpKO9WcNb3zLsyfhDCzNrPtxhmPZZPRu+LUVeZA5zQX6d8XOV52hybnTy9Zjse4eU
N7TU6sLUjV/z1wqc7BgucQzlgaekCLHI1mOe1h4XBLAnUsfhsrgbzQmQKNZqG/SJAXgmviycng28
VJZyrtBINa3rI+seeDnQXKycIJIazTwyKc/2kZhyAWHjcsMRUuP2OgKKWwt9BkjJ0bpxd5RHkWM0
lbcx1gu80Yq5ltwWm2NEYyXtlOnWdhvLZbiiekspUBdlvyaLojuUevkcfF2u7mR38OF58EadPK22
eu3gdErm69txstcp6GOKTcuL1o6LWpSosOxaJ/bnuEKPVdfikicaZ684EYz1Yq5D1wWKMP0U0acE
DB27jr7w83jqP1vLj5oSXXR8YbAKfVF3hNQTnkGyXHNe7p5SIfxx/yaIteXZ4/ypGRS+q1h79Lg5
se7kTfvh3HYrsJmvNo2aSf/8KwkOBRWpfw6IKV1PJlEq4m+oQP6cb3cnoqJ50NfmyUnG59w0AEiw
0RjPFIYlH60lSX+1ebDEvO2BfnS8srEQgAgOdRqi+JLKvB/in1m3X6Km5d6GDxdLrU7e8aUA56Mp
UZXW+V27oybF56Epyx5Hh4um6v1i2aCDoCzkFhrsOGJCZP08M0NXUR9+slqiVTkHAjOlEf92pOca
T+0FVIrUkyT164wmW98wNp0CmWYyWHnlW/VVDskCrAMOcJFLQd25NmBVG6BoRkqtoL2yusdosGGX
Hz/wQf6RSqE6et7rFFBJYVdRhoYe9NSnnATTNk7BzOqVr/kXO9CHaJYeEXvMNS0rQRvuKm+Xn2ot
vI/eMI15nfxwKzEWOoBQS/k9g+Vhahkwup5isf7gkZ35g85Scs9HiGa737T2iLcyg6kyEL+Zm4q3
OQfXZUlUcCATxQotpvS19z5HtrXNboshJ897NECzLYkszNoszOatuVwjpF3Y5HDuk79u6k+xbB67
QlKQUBtpyKk3vWcRQz0FkD+tkgTE7AOz7sPce5Cg0tB5gt8X3GMO+hZEmIKPKXFW7yOFLNQd1IkV
1RBgmj1t3E14XRKTXKyXwOzX7MCPXWN5oDdGd1xCUlH/EiGIG0t8cjsf9/LG+/W4E5g7PjHpisRO
d+XIHVd24ZCVlrm0l7TNiqZlGWrw8IZvcp73f41ruydSl3aTN2H+CLPWiHDny1iSQTcZXRGRga7t
+l2BJ7peNZCIzI1kVuIhZdHxyB3n+RXboeMu+yNbzVHdHrRhC5T7mZH5u/HQsR1mxWjGUpnyuphx
FgCcv1fW88m/GfEJcXOw9drl8OyQLnFRVDz/sU0Enzo6lLZ8D3Z24iOk7mUCLYoaHvCXWxZTee2k
6TFxGVUCVK+ePrlS+pfiiX+z/T/K6wAfsx8M533JQ0SHdiKJkZPMzLOMVia2ceIDw7o+rYs5403N
EWy+u/mQ6jsBKRy97mN7B1THmVIN2blqd0MmbaYduOVTg7pPGD7KemPuhVAPK0kDTYhtVQYPRvsp
Vl0gI46QWxHOro5I0CE7lwlg4oAX3ROi42SykOn15pEUnI4jt7GxybsCIk0Q9bYBjXumEkSVbuGJ
FbJtSJIzUlZYSCSLnEDgYxqcmo9SJIU0GUyHOajvAzzE0yREMyhF0nVroX2HoDMDjqh1V3Z1CFkt
Vcw88BeRUdO3OSYrWokKMuh+NsyiIarS8KxoNvc4LO74MXtzMh0gupn8ufj9Pmg/BKlOZc6OGX9g
o98GEgYBWiRfLA828VXTArGiH9jN0yQxBgrJ6hXjotUntpQUsYwLs2A5m2WO85Mo+ae7Oj/GvsQ0
8Bcns3GQyMFIKy1A+iWLzmnmNu1efwTJ1B/fFC8iM2AKQSAR82Lh0MGPl7inSsc12mr31Xo8/rU+
1xdRd7bD6w/MU0ukbaQiaHSm9W3xmHcue009vWM0X9fjZ+NwWXY8wNLIUNbbdM0wsI0yBMpCA1OK
H6TIBvzv4y/7JT5me2MRmOe7+Lkp1L84gxMrLN2YOSYxdSy0P2fiTomAkScfMPFotyWoGEd+ojli
bcHn7e18uOCrHnAvV5uZTkl13qNymwNoQClmCZXiC2gBAlNM9mQM6cftTsNTEJ9SEoAATQ4gI6KD
OqLXn7/IyqOxuxl1MHS2ejaHMkO4iFv+zxbWIS6eMf+gBfiYhhhMSghyygdfrtSuOHuRnKRC+bXx
lKKLKaFowcMecHU6lFQgh5yKhcEO7XSrnOLyVcIM/3RRZVG49hhrzqvy1ezMBICWnx0S2s0NyTrd
5wOB1xNN8Wf8dZ6r8SaQgMXcX35iFZgGpCawHXpC0ehqC0p+mBwtUsGzQdwojqDyBdAAWRSv2jkP
QTssuAdTZOoku1TF4DOHFhye8TZ3BJyacrDaVP/0ggHR+sFQQ3noYWwEAc6WNGrgvXp9POtzmG/e
YHdGv233SBYMVF31nZvSIzkqYz5K+z2M3XnnY3oqFIEFpAULG4Y1B5+eHInvKdWTJ2hyMH8matHO
A7NYM8pOsQ57AzkQga5ErCFJyfuEGCu2qWfe83to/x4Ny+WflBmb+wWehf1OvSBp6CPdOJTK0w3t
6Y1oEMLOAMdKKbLsBUiLVmc/GDluJ9+G/g2TiML2D1RLsH7u8pqc2aqI77hhjZ71iQ256H6/kBkW
UzRCVsIcjq78BfKJGJWl/pUd0LvPlFap/aQDu2aLx7dZpHwGoejZhRZyo3f1T+N0zQWNfwE9imds
dk78/6vuHJmJ9NZdI09whjS/mmAvA3KYYA5I7dtcla4/YFjWGt48L4h4W60DOdkJE4Aph15zr7VJ
Vo2RWkhGWLNWTsxDyxBat2WntMV27QR5aDlkCtfUgiIlZU/4LDGTzK1c1q1auV4z+jymRw2cwZ+1
Y0TJRvG5MRisjO3IoDwPN+b0Xri6T3cpC9sB0msu+pz1g1AABCMuOPQvk03/slCOHGQwIv1pa+mx
X+3jSvb51Vehq4W6W2LPLAH77necw2ouIxxwA8nyndkzrpqIStH71LDHgqWaq6OxzYQl+guKZ/jL
0zpAPnBczsWgfNcQ4ofDuYlHosJGEGUSEwCq7D9lIicG/UikvnwKRRW5bcER9mfVTKvTPyCeNWxR
nWgQdOJs2bv9uDKVarGyiFKepEyiXvhtT6uA8Hvl+gBjXOw9MJuDwJkb2rLilCagIfIb//87vPQ5
QCjuGKhq0M3QlzTXbX/D7uZa+9ODpVe9EmF/Wk524l4mVgazG3Z4AlAjHT3jxIBYpqo7RwONza8Q
lrI2NJSc4SThXjkhx2Luqw/A7u16P9oPCzGJkGHhrwrFVyH344OEK2NVReejEgOAKMtWYwfQ0HNX
lfsBR3q/6XNnl1w9tc1tsZCdVNtnKKCjGlS8qH3qzzUvE6K/T58DyPJo21URCNcwVEJyf160g6f9
VjVNlW3rBq8Iu5Ioj0CU8hSjRXo5eLf4J3NfGh0+bdlZgwFYwpIX/wIj+2fcnOvJWZ92fCf4oCo+
xJJ/utbHBoaHhRQOxkXkgCQcHBnsG4WZKOCfHlNhSKN8w+4CfG0RBPYi4zNlOLvwjEz03XMfCQPZ
ZRfi8WsysT89+SeRXaBGwwYssMiO2GVNq3jp2c1sy0hhQhOLz9LCTFSJi21T/2TahAwf3v5cGZKQ
4CdLIFMquC0hi2JVO59ERvXHkc61pUw1aah3MySdjxbnjClPybUy5C6FNqSWZwh7WfmM4rCCcWHe
8+UEGPEdXgq0rwR61buZKAKHImb3Qb/1oJDv9ohZfktl2djU6zLmlhmBDn3fsQJxXgU4d1JjwvmK
qhCyV/GMVz/bVroL+1edz5x0N0X5V+eEGLy42ulC2gaw6UkOdWjNWQiOTzOZ6qxDBeWakrx8eYRa
fqKeTIxHciQdRMZAVb5lwbQMVWU5qxnSLVtavwghSpL5DeYq80/6c0WA8xSs8SEaEydRS2E3g4Ex
iDSkY8fmBAzL0LuGe99z6AsiZ2geLRWf7GYO7haZDE4QocpgMKe6mxNhMBSs+uOumWg3Qj2bGoWd
RmING9Pr3dXShUbSl+kBWI6dWdDlADBeYBnL760Pd3/Z+S5sUUH3EnC4HB6pNhoIOcsi+6XvlVUB
7AQ8umNFgNKu2SULDiTx6VLdN4Az3JcMYdZxrOc3u0Gwew5ySUCijRaydwRgQ4/NRzhZYicDWZJX
R6l/UeEZGXZMuEh49rvahhYHeTgI5Ua0z5v0bcKHp1hhbrS760KAp/xmDCmAjSaSid+PHM6lru7D
1VRlwgQXgVWRPC+r1BQlCKekYQG/ZdsydwVp0CLxyBfNdsyV+l+8hxU/OXdZ946I/cKrmBuVjP35
5CwPqDoCHaPhnhTh0POew6ptNYRYt5a6XhtFCGAEUSGwUCHaXZfeHro8Gzek6Vxnsj5VgqWCMwBo
XC3qO8MvRGaEsG7fwhFFesbNHiYdSvZbFU4gaLJ9v82fd4r82qH7AvhFpwdJl4fk2072ofT3oO2t
0qXz9MtkElYyCogx9iltRV8o+1utVChxZV7X1RE1ArSUmCXiIFEpXmEivsIlrz24wh0vwkpr4d1P
JweLozgmTjOI2qG7rf5UjDl3T6IUWlyyhqLXYQT5aujt+o6C3cNx3eHa5uP3UPGEYyHWHhLSqZga
8rZdDOjc+RADkQ69h3pmZuNR9LD86GnE0+vinXxH4fhzgEeV8lJZoHHKP8GMn5RcjaCOaGJHB9eo
gWGDl+kgU9cZ6JlF/XJ8Ebe7k5xFagXIacxDBRXpRdfDu3HNG6iaJ85MUfvljCB1YyrYJ27unjeW
7W6OaiqaQNf+HRZWP7nS2ggEVLjBsmDmDNwuEAsiWqD8NSlM3/dfOuYwGW+REH17IRqnZFNXH7PB
gV/vyJZ5uj6mKeUnFPPAc8MdKmqytFJDMzQWZaumjeQXK/++SiKSQhGgmlL0yhoZ/Uc9+5VFEJ7N
hy0etfMTv9cN+rDanxOTZTXhO6C8oONwZdqYMwni1krwkrtpAm+6LjKrw+uAlSIkVvKZsmHZyH5U
jtdFbIOP/Stg6juPAzDnsl9MuQwA/xLZY8ACk4KQKNjugBhvarRWGNkUQ9XLEboCFjAqvp6zCL7r
ISkUmQrczvxNElWPCgqXx+bDTIUUOzWufaZ10U2in9Ttd25V0lmwO57GoVDVir9a+tbzYqy3b153
jfmkEt5QCHtAaFJAn6Kti2AeYoLbPBdC3j5YbXJDvMXqeI3C7HeIwYEA52GXOM+ioxh1QSCuC1pL
LQqshpFLw1myelMaql1QSB+hdsKMLIpjFn2Aht/sapOiiyFICNyYHFEL7h2rLq5rdlKwVV/s8gRo
+q0Vb8JBJ0JIPp2VW1t8e/7TKY8PSZEfYMozYQo54n/K24YYpWHrmDzuaKyueaWfDdBTU6IiOhEO
sH0T0hnWB06oJlXD0zX9VsXknvmZbWNSyceXZ10HpSECzTkJczQ2ubgUse+Z8kuiHVt4csWdj516
SRh4A4VY7cR+S+6hpvZlNBBWfxd+O0/09NJjhGP+LNSvFMqUjARxDvy3yeh8hoXh2HE3y4jmjhVr
HzJ/3MHP8kbn5y2CM/vnD6hjjKNxYzt6iQ08DSRFNFN2+VGul8eSa9hYN6It689rAenVHZDC3L5v
jhtlNfTZ+QIl0Gh5YJs/ZSow5ZpeXAs6frtIj3WOYLnCDfkKbgypRT0sh75OlGNbsf7Q7s5V89rP
H0SK3KnIQeJZ2cyfLWxSbUD0DQZphDfnH4cuLNn1E12XyMblULsAhj3xH2A/jKzfZ1KPK4UYEscU
FSeYKpDsAa18KzbFTMqwOhRDRHyHBfm9/VB8Kkl0whx+WgsJv4zZ9inoqZ8q+csuJefTREOiPRDP
3iCRvSSFY9pjG3OsEcbL1XBnUk5iHQvQeYdi4prsd4n8IXla0SwNzmgbm6jJT8UcUveUgF9mPbVz
+CpkhZhmotXJ9MF8U8I2LSp2gqnUGoJ/Mmf96tOsO0P1Yd7eaLPkFs6E78c+uOy/0ExpPvCFmfeM
CxNvlmPpjRz12eT843mVumzTTN/uqG7tVMMrER9LetjqtgJA0ocIQ40NOrloJ+V2LaXu04yw0b0T
5mmC6lSNYkQX0FORa/eyshuXBlk6ZjDO/gL0A04BoW9XYTIU8wuYaO46kevtvb/obYBZZZktS2Ni
ZWGwzdB1lQgB+XEmQpyCwwLS7qzBUmi4SB1zTdezWyK009Mzz6uJlElee2hwao9tHSerKKJCLMvR
wUaJZsmVXF4RsEIdUnHnc4brmC1zbJpgUU2sMEVyvHKu5SWUq63aLqeYqX3acTFit7cDNOoeEVos
7YLMcQiFuKtajYgSOVhEQGH2R+N+jwawpHeKvP9HCqPDS+7tpDYVK0P6gtDmZVacWUp3Nm1DQ2m5
iG8ri3maV1/xXKpKHnHXsLpXOIa/FjleNkijUtwUsFUW16ZMoqq/4SvfqJBNRu3QjCAVOb1IZmqG
HvQQpUhdUq8qX9U35sl6cjr1ypxO00D82Kr9/C5p2JB50Jyh1QjLQBjdw/Kess7UZQpHdVe3DOAz
iOzMSrPunsQPbGR0mZcahJpXIV9w4r8mpFBjcL81esE0i3I9/f72nsU9gCa3BgMBa9GcJRVXYf6l
uNkOdOkBKj/PYenVZ2nVTFyP4Npt0IeRDPLpjlqQ0luWirTjAPAzc9hnXZ12BCDXSWv5+hfbFtr9
XrsGG02xg8h4dZyJLbVlrY+QxT/NJYMfqQ+eJq6eKOvYcilnWMIP0PWdYYjVELE8GoanPzyhaNR+
Y/wU86Ee81r7O50xZSMBstbsmWL5yZpuG4i9q9TpmQf4rOWjnWFx9aWimAFPgyMIUMS6HohYRT6A
z9MdMa+XWzla920wUiIaGjEX20PXIJdcd9vZ8MjZQP1T6bTY6V2hubUOZaAZYtboCdDSiG4I2R6r
MRq5fF15vAZCi0NgWEFb15zzPVOarc/I0tgcSEiO76VQBGbCrREXsEF8P/knTQpwV8kEp2vF8cN0
O3PgbS1car3fOTz8+ufGABLL/kpUYrrUefvYA9DqZSljmhOVaKfASYUWsczKKCaWiM7OYmQZum/P
Cd+f9eniS3NM/8Xvs8NCs3EW0DKA71tIdckrdo+V0rUZlcX+esHuem/fGjWzBr7z2vC2mt7DsCuB
v7wLSjOpyAWRDmEomoHcwEFWWBVLftg1I2fXYFFrxmo4sslRN1/wZhfmgjfQIym525SJdMzEUTlu
96J5pThq8ytFnPT1T6BRYkogEKJRM69WEv13R34AhdeMytGvboA1Sd8jqbr7NIF06Hd3PfVPS91b
8DMDOWpLwYOuOjzKtxIUYzAIPjsTlb5rWIMpiBdfoUlpAeHJKdwndiDIhXo1GiKQ07/rs4NSSLxB
I3cIdBKMn5sy/GWtTbEtMPhicac5hwfhyJyGeH9O6R1Wd6oXfv1uhOEgfrQCiW8Hv7y2xtN8bkyo
Sh6O4B6SN8CrNWZRpYmjEoVlCGBVyXS1c1D0ZKoDE7TdcrXK4vo/uOpmxj2YQ9JJkKSAmeawx0GA
fNOt6c2p7wunecw5P5XqSsvCxXGVgbl0si9sUJ1zMUZUzVeRWf1bvovQfD/6zvJW74tWhuk12TzU
54oKvYicQIUxbxQx4PHu7DgOkHtRzvxkMCoEvhtA+9NBxUiI3qXot65j6kCti2Bs455u3jkHqHcf
n4MSHbYofLMgO1DZc+frqeSDyt/xb7U6IAN//Vh3BN5p0VBOalwtKpdZUXpXcsw0z3+6nCVfJXvV
5ZragYr/ZGFQXZ+D1799B3fnyeEmpGJ16bd0kpmpUoUvMOyA3QAW5ZPdxF2zEUsHjE46rEwz6N5Z
opP5EfDZBGsIdD7bPZUTsGT6KoGPsBKgZZDopcINHTpdl03uXT8vP4Zty+Y5L0fArbNupjjw31w+
0+1fS6mRUdj55chAOZ4Z9BFtCzAiHYo8z7egPjnf0JiA/Hj1/aG1IZRUfW6Kkr4+LyaRKs1XTC56
6e03KQdGo/ADoB+xENSU+CYIH5l/Qd6EoqY63s70ZtDTy1/3CLSfY1rG+OrTsJdAr7Am43Vqbj1V
oFPCkSmAKOhtCvYK5D8mnCXQpXrgwPn+bHhUUpMrQ8jMOL1rg+13J6cMKdx5JPHyBeHsuj/UUa1x
EzLQoEbw/JMLZasBsJ8p4HYacresyqRxVAJWtZIrvRNZKLfjmu7vl87ZlOc4kZFF1Xk7aikCr+S4
Agyhto3+iOD65eoOmPOMxDL6uMYP9Z6hkZX33BIS85yxa+F9V4X3I33jLx525ifwW2+G2nh+Tppi
K2AQjzWGDpBj+jt+qbhiaVm3lkSBhqshWr8eIjpIFsE+sEMRmNCmslAFlVqHR+XjITBJvX8VDSl5
LzkcU8laBEN07vzDyOgDB+HQQAio4rYKV7+7Q6boWqF4QvEDzR+fVn8hORmZQm4qZpjL1JQOVn3V
2G5su4eXTKX9MPGIpDJcZ53fCx7CbllTCOXWE6PtGcNywwBcFiPdz4jR13kuQ+XA8M3YK8KHZQNh
AGo+uh/9NjVSOs1ISk0zHijY8VQkMxqkLN6u9yIeiR44yAjXka7sEllppOhbN5QCl1fnM/eZ/p7E
HuTYDEERzjNhncoCdFZ27d67P6EKWR3VyX/r/U/HoNvi3BjuMUu02rmp5+vsqOD6WHXn3CU78HdX
sHGLFvvXuOf7FvhuDnqyW4CTNesp2ef+C4F8lgdovDtvT9dwqo5L4NL9XUOby/d2bmG4h6Yc+T3T
LN2P4cw6/Pz04xtS2D5psqXuDZ/mk+LOsVJaM3pZ0ASsmkHeA2asMHEPmlbhOdRNWq5DWhpEYp0x
K+602AxgQZzuk9GHnJ2Cjk7kWWaad7lYqMEuJg4dV2WpvTwWEFND7F1NtKFIiV/TXamFjaENUUdr
tFojd++AGWte3KSScNJlERFJdZZWezulJgZ+yI69lieE+KWYWTDI+No3CoBvhdYqMBNINYBzB1Bb
ViViIoi2eDM+kRXiycYzSTmnt0Z70nIcY535JfJBi/EB0uFIyASbPW5GlXVsIa5N+1AE7YMM3+xM
8VvWmBu+dwFtxvN6vzRDPT+DbNrEHXJhS1x0xyhBQWw6BmVTW+8bsYNRdL7wJGGVprnJ9vmVYK1Q
K98gpNH/lwlKj2C7ue8KuHEMAR42fwemzEAwyK4mTJnPMvMOsA4wpVH2WWNYiL2eTalZxPSTatSq
A84sLHkAuFkNwIFv2OsKdbmHIEe6EH0Eg3OCN1k6YAeztEC5M8SHBwLt8Tat3HeBF9VKDb2xR55c
UxD91bQb/mF2W9AhmcjyCy45vtib94vp7TDmoUZ8rrKctiiZwLVlmX6IrlXSBTRHmyFLF31xkXNU
nay/L5mNUKb1GsDU6XX7ARjMzzlkQdgLnEQY3YyLwd9h5yXTt0RksVCZ0bVZ2MDodf/oDEoVDbz8
UbsbYhVaNMuSUzSFcntjgblBdiZJg6kf2oD4+EFU6iw77vrhmHPXIXLXEyaaUorDpa3JBamaq8L+
2cBJniXzjBcPwqALKSd9T+fi/+bVO3lO+1+LvUIDxsbvBL5YR+gmoxElyIvfJKLvutSCXzeIgq1O
iKlP3XuUP/FXufF6A7tkIj2bkv4kKLTSEISvsA4rbujoduvbkBtNv2FwaKHtwVJ639T8sMLzBPJM
37CAYJkuBvERwW0nSR3HV71Do7iT5UyzsTHS0HReZLN5w9V5VXT9DWHvhAwFtDe0RnfW1X4LqZsO
RP//+GtOO/4QENnTWgPBbFceuxoK3LEC9Y5zB5p8wpSe8NlybNp+zMb8cuYOcWjmNP334q1CO8pB
bDWXUOtHj7/bs2KKGQa+hGlrpuOsICgZYUSuRq9m18vMAivcKm+FllduUS+9zGtFEzTcMF+9ZD8n
yKAbDy1lNaza6dW2eJzoj7PnyQoP841sPXeg2TXy1q7O/R6pRxWmBTB3x9jBMkMI3IYq3156PHQl
VXZVrARrFAjsB3HSJ3R+BGE1pYB2+ZbbPxjNshb/vohmbDw0heDXyuJF8uezkMrQ09yiEDj/M3pB
AzDqV8xPV/kZ/epVDlxB1EVR7zMgRF9178ki1kyW2j70Nngpa5PWGy7cVJEaqpA41cPmtM2xzwZ5
PnfxCPVyauqMmx/jsUT9CBS59Zl2lA3sGaHBuXF4TOZ3mujIp8HjB9ypxBzPKCZcD7zkz4aVeu7O
CCtPY4k8fK2613qiWwhWLBlUqBMULkaGr9AIlPS8RQrHQH2cVSbey/vUgPw4Rb3+cGFYf1hmAVBm
8kdAYj94nMjBHW/VF+scOKrUVEpoQvduNnS+sBNRUJ2rgdazuHFI9QEOyyWjbub2lQi7c4dBKfXO
GeVdn5YZIHyCRBKoDa+d/CBUQvmbYOIw9XOmRsCQcs5TBSI9G6w5A23wpf7x3vgWsSYSDc86u6i2
d4QYNCDidVh2cRWMcCuLEb1xKEHV0UWwIAa64zboevax82TVPtsffThA1GSHpE1ukhA/4d4Dlp4r
r9Ut6+aAfbSolBz7YDuhNorEZTPdd/in16PXhcNVDTImzZJSC4paN1iV/WVi06iivw8e0f6Pvd+p
YZ02DSZXTkHP3VXR5cQSBagvbccT495MN+nOPyaT+VPgMx7mqMixFyxbdluyPWtnbU/+hCKLgr8O
Lb2y+7WCZ99y0ha+kSRHPBWg7Ih5zEH2NEwzO6sFNzfKvHLATLsImSZonsZ86RhU/XuFCQNrCBB5
`protect end_protected

