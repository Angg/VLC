

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
lSrzbkVRez7TSrqtMj3fFBoVDIfcRk6Ys0Ryw08YT0xybeh4Imxhh4Xo5waHds9EoAp/p211hEtH
U6pvrX+agg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
icUbHhj5bYGT0RXX0Hkl3qTy8gXjmaBdYmbJdfGSlDqT36aBG1MHxVot4QdFfhzT4y4EGe95lWcG
bY7yIo2Z80wxkaYltPsUfmPKSryRYnC2RQpCalRwEyIV5kwyjLyH2PMI318/DGe2zOgfAhyaJa7F
upzBPe1dc9VfrYuArL0=


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
PxuYgPP9isSAWV6BDGFF7E4+ZyEAPJFkhVqMkmalejPpQU0gnnWwnBm+iezC17JL/Xa/VJE7sfaC
AKrBOUostq0vvu1xdTV/TiVQSkSuCL/ILd0KvrM7zY7byDcLHbE/HiK9qAiuHZ9X9afXOA3LUXa+
NeIijoXYNpcPKApFE7k=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
MiGbO+1/w2LzUP9w4vcJyQmRyNSWoFP9CtT7NIPM6EmL2LPHcWpvAOqX6yz7ntfA7Pj/Wid64Hgu
shoIM7ZLSfclvZdj2d/qq8ODrS3OvMB2omZlH7/9Hf8BNQx5cdlMGt2EQPapbaczdAOSVlqfQP11
66CJpcIpu9PYPqIPi7gr0sPciFBMJNEeJMdBTGrQns4LBfJmDRE5WdPDo1iDs7+I/XoFMkZhvL/0
Y91WipnQHvefAAlRLwBWNzObJ2omUnJDqA4fEy8FyO94l2UP+gXZJY6q7Ahrfb11AzhWCQy1/6kO
U8WeGtgOmdPeP2ApeGCjofaQkPasVPK93MY9gA==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
J0hRzoctT5uNrkbAOYhG/C1YYiqLYlvZtqfLxqcUZK7708gdRGZirVbjbqEBeXYlyHsw5AvqFtqw
52FoZUAEGkFlwIgKWxiJl46IuvZVYEef2NF6y5tgMHwEjkFVh359FztlWhDp38jj/NzWHKBOuK7b
WD+057fNTohIPJ/bd3naYCO9ZKinhXefS8bjBLsa/MNn2ksi+KfipLV2LY3t2pcBC1wui2dHqGvO
RvXXOCVCULpb1KAf8M0xySyzObSjDR2pgz7PdVOuusTxXaD7SgOSTCuvcYLUI/CgGUFhDdSfpo/T
KUE844cAUxLN5mN+SZcv8YXfgpboB0XGbtZjjg==


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qRYjS1MWZ9AEGoXk7XbPnWevWA7a0pAx3waQwdjQYrYZZwvwBmZMyfVb85xxDCsnqBfY/X+z1MGN
R6wP+/VkRwqWybLkCI2H+eY/JIxV8wnXukunleMgiWrZralQzn5HM8wFmhN51HFEHt8MehA+1v8V
GkbvyB+NWGe5V/g+PjZbUP7Rip9Ktc37bLfQ+BBs+LxyODu4QecoyoLN210+e2fQTtiawB4NhORz
sjQ8EkpqOIGx6NCgriSXgG0/5bBCy/0+EaWSre9yzV96ovJXPqneFAFAykHGk0lwBtE2N2jTlUmq
4YOLU9hzvqdkuVeyE1y7f4GZCgyIM0Ch4LciMA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64000)
`protect data_block
AAAAAAAAAAD30MuU/X8AAIWktoPPMDGdpPxgKllEE9xsrCxg21dhH/9rJbpkD4VW3vgDOqI1b2lL
IaN7ZEu/MTD8wqxzO7FL6gz4sN2pFrTSeWsihnGq4scBzvAIX+ohYky1Owm/5WGAgainECp2WOvK
hO6u+VTk14XcGY8Gh1tS3ZLhX4ds51FJQzhCkQI2bH4m/f18VyzM89Bqzl3Zss1w5+UbTkPIxHp3
JWuFvldJs0wDV2E/3j/RHRfBeiWu9hVRFsXeFtbNb2+JVxq24WXlVJ3vHkxDG4VfOXcatV+CewZh
hYJhu19kwkRIT25gv7IzmqIPM2JJRg2vbthGfRfN9Hg93FF/HIQ3sPHUKuTkB6YL+oAu4h9uDGiV
lwl+kF26GRv7d9+4vY8P1tV60wB51saY1lAa5rtYSg6svMRb5bOk7xan5D6zPsB5TMSZki4fhLsS
1RVz3AzmCBI+aBQCnuLjaKubXI9Qb+ElO3WSQDUjKQHzK/go+8qCmnondvHboQdvTDvOataG0Jvt
GX9K47/2bEqDDHQ7ZhFo8C+N4989S5qYtqC84K1nkSoV8xhMtfAj/jO6OjxdsTmeYY995RHRU6Wg
EfQsv68R7qM0PRkQIYOXQjR81t0k6Pr2B1dKGP+6R5htJ1239uoA99MJLpdhnEA9OT3teYhF6CjR
xnr/EJxBiLlzISYBIfipHHoIhoxoHP93lCh2NdJzABlbpUiioezoYUeUtXVz0zcBorqWnQesRkDK
i5ikg7Gz0mQa1F11VmvwinB5OkHIxoYMy3L9AODUo9CGBDC9xZkfzwiMg6b5z9QZXb2Iu0RXTcK/
3xKWYVNlGRvNLiawshrn2FMKFvM8oaxbXdLjSeun8IzlBZeMDww1roSuQFj2EsysWzkM2oJk9S0G
dS6MHgmXr3dV9NIHRG/hIxuRA54pJFt/FtqUSFa7/2+3Wu95shyVlzYEO65kptHlap7bVk4W0kG5
ATwNxjRZUtbgYvk2Q8WwMMJgGBhL6oTkBPQdkSd7AqlmbIcLPTw6w6QgOTf4BZHerDOFLO4gecsn
nqkEzxdOLwksd/g6YyQ6T31qYZoHQ8jb9fYG4ClzDtFS93wY/3Ao3nBgMWgvgqaV76kdyuaII11X
++mU9a+Lpth3/s7w1FznULD7yl40v6DUk0M3QQ168QO+aINm1RQlny3ZrTud+G88IbwYkZMrBmHY
LYh2JZq8N2GNenPw9T03JTx+ttzm5RjSRvEVKcojhn8XYd49BYc3ttv9Ecypefjq7bxjePN03KpA
G47fx9Ea/wHqdVNBCJ2UZas+BliTNtYijJExT4g5MpnfLHavEuQVg0ITsj98UpcXfBps2fTettKl
i6qnruWMYvTz2FXawxIPC/p4Gp/d156Cv7nMsfEVwjeh+gga0HeGkdh2bZSay47G379bx4rgokb+
yUcs5QUt9BTHbUoxGOIzwzLPJoXnlVpJiqI2LmYGLYqWeFC0XRTxrVg4WOVuMNq98nPCe2RKfGby
SAUs9FVX/JjsRKEhq5gPURZxPLYvraqJyv/AMEPaStRuT0UA9tb63VerEB2dKim9BB9HymdWx741
f/mPVtr1FPX8lnZqiCV+WvxITzxzluBkmq+mCFSAdLPFfAIEAd+OkSDKuP/zb62rjHC+40KR/8Gr
H7EP/MbijmQd+Hax0dQfzM8k7baOY7S7p+RRHvkFCZoy1bHrkaXkXAr85iv+7Jk9vBl+y9cF86oA
SHb0q0QFyvkyQVjlBv8m4ys4COrDnAqCMJ03g/UFj3KmIYjZWJWSY3MY95QjQ/8W9uaOCpz13+sT
xwwwRIMXKqWFPOuZJxMYPsxKqDWuH2D4QldVxSgjvtMr5Zwl42320MdkTFLke+UAcjw3cJTP9rtV
5Jyp/R8xZBsDNJLZEwFm6AngDGpRcBgWvNrBoHhhfHNxMt7jvwcbWOloHplyqfH7LO+VEOMxoM9n
l+EbEzFMU7Itnl02HAR+30P3LQP1gDBDWWQhc5lVfUqylbow3bq/laEwKHkQimYTTM1smGb1lBIP
RADJrarD4Y1AkRK2i6fq7duJweduq35GZ+UI3ft8x5fE/c40JRDyAqqoULY9ur4L3tgYAgGNtVX3
ZeMZq1HScwcK6o3+UxrCZteG0kvLsuakr/RT/Zp3T7tLVqitsyEB5daevj66WAn/Qh+ChONazZYw
m/JAeyludwD8GnA0+4VoS1zZep5KFrEMTqYfRMWXTZ0sOMEfNmhhBSH1VhNL9p9P6wW5FpTE49Yx
lATkPNbA5lY33KrrP3f/NycNFfb+uD45yzDKtbrSlNCgSXAh/wLu2T5turbP69LPdGDRxTLjC3Vm
MxaecHB9dJytXzyR7D3qTi6DGPfEtfkMixJ5bguFYLA+l9NwIqqBHyGZRnOq+xDjN219ELw+lh1j
BN/aVZQxDtpLjJ4nmjROsgrYPLIAxDd6EKNYkYcn97vGFoBZE7qhWA40EYfR91V2rSRr6su3wv58
GLQ4FXo13h6B+5XMSqPKO0rtKhPgHfZeqrRL8+dblXAcB+WApVM/D2NuyoXk+DkTyyMzcqeVg6wG
wm0A79782dICgTiFU/dG/XqJe30lROKGceZPhxIq/5nySJtgQsL9zzVF76AE7uO2RnsKqiO1Fvrq
hoPaPiNxUlirMjV7yUwucu0xZEaDyUb/X98WAfAPm6Hs5EYzlSEMeZT53Sn4NVpyUNVhGYHb42XI
GID3IukLqQXuHpuW4y2eNJhFon1otPSlFfVlZguEfbKXGg35Dc3w7Rc4V7JDYFtyHR1Hq47P6YQV
jydn/9zAASw3H+FaE7SkbwucoXwJ/08Ro90GsoHbGw2cUO089KWEa9JD2CMg67VNJxoRNbszZHDR
BCFi7JgRiSQrx3g0ciW5ZjJSoY/EhhqnBt3VYwgPVSi4CuzpVZdIoXxcyKgSZGIoriBjfn1/pXcJ
t7Y+QDho9Ct9py2IiXA55HUDxUw2j8SdA9aVSGwxmNlt4hayRFZUBluPdp2woZZSGxf1Kv6Jtr0B
S9kkI+Lc9ckfjCv9lzhGcj+hdrRsVaCjgM7wHq1AlBg1jHk8nKSD1In0GYTDT3TCkyi1NVb+oa7l
E2igSH22ibNmIx2iZZ+EgNibhYUm6byES8SVPujKplS67FtTf9SJ45KO2xv5LI41Vhx0nzbVLQsy
o02pIH+HAQGJ8b825vP39ig82td89q6YhE+Tz2EOue0wMcmrl4GTfHyxSln6ScnZwdsqxqDIK0TQ
hzXVX61x97cO6uRo6IIpJbxkq0gtir7giQQHaX6LySdbBDbYPMhO9Djow/WRKA29/iB9qdstKypj
fpJeH9yDi3VZohY0iaYKkTamIzDnbYQ7ovmLwr5st1oazpkqqOGzDbLxlY0bPK30G4ReD7cDbCQe
laUFDMWoefklsQMzSXcaNjsHxwOCsCRMerzzXRYy251FgCr1KUveZNERKlz0EwY5PJ0B/6Si3UwL
S9YceJNe3IbIHs/uiefZh7UXrFbp88AYrXlZDpG965m0v38Xc44pv5xhAeOn/kM5I2kgBDPf1TBa
Fct0XKAovu6Mf7EMiK9vINAKTj8uMqWhiSs8d8iUCLgcORGBi92Ph4SCqC6oIngN9BCW7Zd3J+aQ
Fz4i7vaSRa7Ak1zKHZk8D4p8nVA5dUBtaMKSndVlUQJ3xtSOtnj+VSMWtFa6uUnbXpvJyzMNyrTV
R2XlX5jGVkA/MLBkRM26Wju2OMSBND8uLwyjd5q8LCcTFzYuW5ojdH0bZhZxjpotHs2LBEpuEeKT
SLnYhmAmHCUMaumyBq7AvqvpTq0FmpFJdzVqzqpIhq85F95f3bQr7qVjJwG//UnEyYtMCCbHDDRH
kh427dXKtJAUKurlkOE/zF5toOWFuzix2NCLR0/DHVKMsIoFST/m7eWflslEQa24gUfv3xvm8cok
2aXg/a3KT2CLqk5vLwi1KMZSJA43cam226Ts1VSJMn49XToJk+Pg+RwdBiiZEPhY54jwWVXVNiN1
5tJzMt6HfS4HvKym33HwMyO8Yzq8neaD+rF2c091oDpuuNVPcr1Ix2zJpKrxe9SjY7qub89Wv70b
Do6sPf4w/Iz5G/Ly4LKjyw+qClURNeO6eMID+wvBLh+6njsLKkqRV5YK6Y4unPfhjrI1IcuiKhmB
kUJGdmJWWqwtrfne4liHUf3nWPcLRuLy2b6EwARlVT1/jNXio4CbsPkvTfjGhAhQp/EH/hKxuvp3
9f9Kitn0fyetVQKTxYBfPyTP1t7e6ZZOguHxRm3uxwrEBDA52nWrC5jnGFrhyS9hJ1tJ66mkkyKP
16wEER8mpxwgGMbfML/M/z8vg2XlPcOqAFJjeYt/Zd2Pt6F6VyJVgZV824fnX5vU7LF2r5ZeE/vn
wFDgIGJdEd/Q6l5rGOEwYtVVZQOglnr+ZNFLxuYWZpleEoCw+x9+uKaIOW2lnEunYJvfZGXqCl6p
Hg3auRDFOsmQ2y4gcURuZ0YRnDwDX+V/MevuhsUovVZofsPjgs59RWShi05I7IrUrysABhHjMhQW
wFAfTifQiQ6evQEMhsFKBZIQqszdqeaZBSW+4ORuwfK115IAyXq//wVUpHVI+7RwviPColpbAeyt
BKOCGHsnYKr+CTZchqG6qRVPQxrECQOXi/3NTR612vySSVOVKJTJWocRoBMMHRV4Apr8LqzumqyC
Bf7Hiu+SGDGv8EGTqvIzuQKUEdJ0XrUIgn0vZCgyhFHijHfou1PvKrS45yQk7vruHVg9ceRdH8bf
6MCDCJgXl8L1uwlTiL2hss34OeKQJx3FaV9TLuZB0vW5N3SEWB9M2RKL3pGbyyH+Wex80llhd1Dk
2sasGaiAhmTzX1BLQ9I22HMOssP4ZEw55LWMgcB5hkisgm2fTNxosbwLfE/94OdWTOmy4ndeIFUj
S93r1JQi/IrgF0Z3mKu32QbwmAX742ZeJjW4adaIPYcHcxzg2QEHM5z56GMeIIfPbZpPMkrGcf1C
wZUYV2fzMZ61NTG5hUQfzyDWFafeeqlt5212bfPL/tvKePyQ7u5yOZ45bxel6BGjlGC2B3Kr4nKR
J6KOF1KfAHLOIurE/y+rEMttbDgGawfUFCu2Aqnv6eavSG0gBYQg9Nj3tq8kkACVSgX4Xirhf1Kf
2K2W2XoRRzJpB8CG+4BiLhqfxVqedO29LiXCQhRkTdiWw59s5ZqCpo2mtyliufsZHVo/roCCe3IS
Rlmt4PBznjgFpOKIjSvPrWfl5HBQHOv37cfFqBkrwaXedXQ2wsQZFYzsLIejZqZqkGu48+0jIMFU
Wc9qIxDzJrG2ujo69vktJfx+O1XqdK6C8VBeiCC/m3CkYXI4HUtC1d9NEO/OXpPECHJ0h9xseppe
VmovIe+Dw7KbuV9lrXPI070C3aD52lCTAZncZpG0aEpHM2jP3FL+ifaIbJx33haNY0xxO4Mr+Qyv
ohWUJd0n38D/VZ7MFGuv5DW5/ZROcAXx/9a5hRZl2IDN2XP1xLDsPhr/522hCH6XGJIc3IJAOJkx
V6WsGTKjJNf8K33+3DHuRU5gsvwJQiDFJl1KdGJWzaiXrF9DARKcPHWhcOITo+BM1pBkXCpjqgPl
LvXQlZKxoPb5k8ihAfVpHnJ2goEuUUpMU1bL2sSEKIxLggrdcr3oX24/7JaqUdEB4CjIb+bLWhYB
ms5jex66e57czZrg6k9JfLMRaIpxlhE9xWH0ndVyk1fLsr5TeV+1iMdUx0zb7cN9AWD21qhsO7NF
FoOOuYy9UKHkW1ZO0QSziLXB9rA2VZNe6oGCRdq9ErxKsOleTL5l4kGxey8Hi+REaRuVso6dcQNh
8g5UzbqjCQaUPz7UZCMYzjfDYqALlxSrAwRPvcO57+KV2g0it082qVdzGVPvSHVdUWRrAwNH7LTU
wHHT0mSYUhJlozxCLeJ4YC4feZl3+rzXUjQM2c3cD1e1JQEJi1SQJvFZLK39MhLFzTCs7r9LUXVl
YeMad4KqGgHPV/xlb87wBFklQAtCS3wlug/kxGFHQ5Nmtv72gsw+CYDpXzjamDKmPImU7l3sTvhi
7AtWUqH4jR9d4iDl2HRBrttD/Sugzg6GCs7qNnOv5RVFv5NISKlSXigGpuo7raIKEQqKXSDYOQTu
52gxmY0jXIgP9F8b+9qoIrLiGNto3di2biIacRJTkhTCiXYEPJp0JdlKzHEbvlP/wsBtxbaIjd0N
Q3lRbSClNYt3b34zLw+HipwqJYjwGVUIpLcNh8O3GEtv2QsSKUlhMLC0ljNnrIMLeAd5c7x9x5vV
7sJVKjCjasjJOQA3RrewtjmW951uLywuF8f3YmjHjdJOmOPwC2+oIyRWmqINjjPcpNea5v7SP186
IUV5xPQOKICtxRk/84dCKXCa2DfB/9gsokj/s5DTQ7srgNLVf2tiAYyx+yGrSzjz2Tg+6sZ5XuAJ
1zVfR1hJhWRkFpuz8lFFZjYusjx+CAk2EhpZQ+lsQ0lGe5J9X3dbn2rdeXXtvNSzF7/0wYTx6KgY
5VCLF+H6cdEeHgmh+kG+8J4ApjyZYvqIj5U2VW+WPkOPvkq23ik0KiKjeRfsoRfx657qi9Y/JL81
Pjpzttyc8LLD4i6IsVjLh8cCoNdwF2qb3Vv59ycJJ4Bmtb3wnzwGSS0Glgx3goQ/lUH+uRTxtvxK
8Iz8YW4fJ8LnBbySi3GqHyhiv8NbE7f2Cv5uEcruWfxbkc/2kOAZzZjyYhRtf8asL3XoNIOhJG/G
l7zg2uHPQPvGQndl4MPd558Eqk+7wvMFhzixn3OODFIEv0nFolkUxsyW4EwkPmQCVfuDDJWBCFht
kDduJNeXztPKzUC1G3c72+C+Ni2/glqTdpH0NzgFajiVypkgNwIdcMsDPmd0Aagaz2NMuelOeYGx
orAj9bS6Zd1zT4QiJqXjrmaBZxhTB7UXiT+dzUTzdbeuyOj6mY70iza0wvDqxkPlwe3cHVHhtqDF
/xJbf6Iz2tCIc/fxrqkRrvWmMbo2CXWQZ6Kq/dXBExQR+MtGHld/thDnT/Grx9xZpSfmaY+2UCKM
eH35yiXLWJgpuRBKy4lWiPr9tVJJ1qSAFEZ9CZLTz107tyx7fj6K4SsIkj5iI+954DaIdEP/48ZB
Co9c+zU3P0aHKOX76xk0GXKBPmU1W1t+X6H+aAEsT9XNluj1qcvH3hPAUUyq4gYYDcIT0zgBcuZq
2V8p65l1h/JP8FgrpTwTkPOGF/HdWUcW/sYkRxzXjsLcs0ve6sH+FQsnL2cwk9cNhvrzWHnqqmo9
/7NUA3L08jvR9/0kY70aUPUSRFnh9LmQWr5g0KDNSBySxGvCcw3qVJLhLZHV5eO8IRWxg2NUZ7xI
8zlExB3dHTPfMte8KWx4bNr/YOqQ12D/2NJJ+Vqer7KVZkVi0nPexJZO92HkDAJU54/eJ7DO8vb2
aTxJgb2bXlrUmp6KyCgHYAho+xzkR8YS0x6ARGArwqaCipeB+wWRL7asmFQ1HRzURz1iFEr9lJbW
9YHjH1N+zK38dQxz+ZuQqBXk1tzpuAsBpNof/x6BWSYQegbJ0rpU0Y9AD9EhhSVWS5rC+owk2mMz
fqwLfVF+g3zl0TtErQdnagJTd/vrvloIt7Y1Lej3Svb8EE/QjrE1F1uMyzkVswjX6q+z4ytVBerE
1BeTKXMj6aQByk7oM2/sGZefw4QuTiql3lPvmqX9UAPbKUnI803h/hr5b875xRyZVDJVoLM5cOZp
JRCjr+TLIfVHbXcyeuWCJtnclRrXd33sOWEmBaI1fw8pv/DjGp+FpKHWVUoQLJXA52qZs6cofirI
htG1IG6OHjOyzY2uSBmTa/su9IgMyGqjBt6gsRBKA2wOUq008TTbeueYKhBtFk2S+IhOUsLkSPG7
Qi6i6/iUJ7hWf2jJFPhHxdWbGkeH3ZtZ6O5Ttwc+X03K6Jdb4CGmsZT15qYD+GMzGZIxZiItEbdo
ZYZ/ibUy9EWfjjJJzBD1Nr1uSMI7i4uAH+kAa5rp1RLfhUU9JK8TzWIc/Am5FsuRs1h2dGRmyJ68
qZw9cuXRVsg8BDfC/q1YwHYrCYFkovDrFO8TIMB35DBpaEtFh2sWP/86zBoe4pF0ZCfb5fqr9vUk
arqXMksB0/WDwvpM11k5Re0/srtVEEDc65fpDCMv6snYfCoUJEzt0F7acZvQBWyWobe7JtcMmILl
Rb7/VJe9x1P+xCGxLuW/hGF8vO+w+/lIhM6F7MBCY7Zg6qSr3O7o3qgwX/si5d05mJxGw4eI4fdx
baekgjqn/xMZ/dmEwy/05uPlf44tPkFM18Kmj5YYj9p3GPtba9zSGCJSqng+NTqCcwwGcSGqD2+d
T6D6gbGv0Ze//l2ACffhy+3FiZ03TIWngqdDOB2OuPnyEdkQanPB0hZexBJBIheZOxIIZI8WYX7K
1D1WWpQ/053UWr+3aU6Nxm2bjw9eSmSyTwSk6AQwJlFZbHvZi2QjEp2Tncc03TiaAYDnH++C8raY
G5VghWdMvgOt8XCqmoPJJOSnghA/XDaZkO164k40MZ3GL5rSMZWSkcibgPaeGynCfUviE7u4aGXA
3QD7oa/wligQgBBbH0Kto6eeTFrOGsMorv1sZNzCvwCnkBOIRiU97bpRutol0N9Fep9nwjoZU+Rm
WjddyeOw2OdrH0yc9lz4LBGQ4MCzMiEhkG39G401FJhI6c3dqH13PZAQ0a4BKF9fgTjaBuB7b34D
l8N47sTxME0z8iMO8uPaer+jpZ/aK2PjH787+O61Z6LGOHTXo7xs8igrtAMwJVbFIL0DFBZNvFIA
XOi0ehzdUkpEoYHemaAAiqaULAZ2ZtyQVCIv1k5n5WnHn2M5+m1LBmYlzYf7Casqk392K7vV2OcV
QbqAa6QTDJF/WEvJefOhLOwBAKx5z0wGrrCEF9gbxaRj+MMmGk59Ti75c6QC5EWo4y+Wgt6QEPsF
u1X/JTXOBe5g6UBM49TLCMeps21FL570cxBTL709EZ8PNT5DGkWXsuOBTbP+5YjT5bej7UYwxrwT
GFgd1vEkPD4uAD+qAMKaFRwz34YFiU62by+iIuV2EWkodLEFmaaD1H1e/PZrARoWKgKBnecByZXf
ocnEw+CZqeWz2jaAXbMclSlSc7mg/B9aE7if4ePgfgbaSXndXcv7hvV9E09dklEHX2apPj8bzTDh
qwVrdlrhsIjL/LT54PzOppfCOSFv3vC8L/mEiu0E68TYyS+NAspxLfOkr4E8o6Sv9jTRJyPxv7eR
lbarCR312H3r5GbqdIHJgUV3Fr2qnzz3fAVhpiEL8FdBo4vUE1m3oktEM8CBjNyacqWOqaxy1AUg
J+/AdxcZrQ8y9RHxyVNew7HxJKHTdHThl4tFW06xrJSUV3iCM/h/buHxBAWLt6Cz4YQ8YlZbpeUa
CjH9ED+b2PSIslliOgVc7t6hdvrHFRnGa+z+/4H/TEA9MKUFtLTI9azFF/vvWrqbsVzG7uaJ4ADG
GvY3Hl3fsmD+uS6MccoQmQKsuFoySV1sRNwvFt8t2oM+66X1lBAs4VyfYctTA5b+3UcQutzUu0Ln
EBsfuR+DteGV0ahpsEePJ6bSCaxlRQX9i3XaWmxemK4fMPRabqAVRzKjHizZAg5XLFSVvkgCop5g
a3Pow7kGGLuqOOLbbXITjD/K7bX4OdQ96sPwkyYRqbcLG9hrLVmATTAHKXI2DRnHRXe7Rsin7ekf
5BvRAMnJzccOBN3RDsMkS6631O5BGaQUfhQflisyt5N6ROYqxWc4Fy6YhIV+IxCdiunkRtZJOtOD
DnJe3HW8UI+68Vj8DOo2pzRGc79K0DT+zablEIGhSI+qvlnd1OLxmIuqwgBSQC4KCePvRSi6UD4H
FhZujCdLXQSxs3fQ83UWX/tgHrmYuNi9ZWMPBfTdIDiFkV66nfz0f7r9jyLP6Nb7nXB/hSjfK9yu
kCa3aHpjyGGSjPKliO3kYfmvzXztGzXmolc32qbaXPrJiyRTa/yjiCqH64JfRHQEAOIERVtb2YM1
2PmKT4q+X5pQDXaUw9rfs3rbd7rOSSznLqiTgLGy9nmjtSqEEAOjYUfTSA/xfulZxcqKeX1F77rg
e46tLeTH1lkhwvlvVoQC0DPnpYHT1pYSP/4JRhbD9bw1TLpa+Ohd1ErL2Td5ug9+foMlw6endCQ6
zfvLbMBnY+0usujx/po+xUPOiX9OSl4z8uSIudEgqsYwtvThmX7+rJ1VCVTbou2KjCy9qtkaheOz
2PbfGsrRev8/Nm2TazCJafxzVS2RpjdD7vEzaqBHx5obOlTP97PHuqgxb/ajapwArD5PYQs//kQv
YcB5HBxMrxvAPuReYaHM8yTKurCNsJ7ha8vJmNuBVwsXQvAKNhEwcGTuL+7S9eBXB4sXwGbr5D7u
oBs9w+t/9dafOghxMvxQrVmbOwTHBbxNu7sJNoyQ2AE4Iy+gtK9RcjizuCG9AxrVTxZjrir29rq3
P4jkoQibz5sPMhOZ2oXizf9xb0+8eHcz59gVm0CDZB3Uxmc0pkDyvsQ2zFCNjmnoZHSpYa0ktkku
4Ay3LIlQNrmEj1uZDL+X60WWaHiSMfC0DHN5DCl+MMnUcTUPpL7RturNGrEM9hd3tzQguP+hL9qV
CwDiYJ4m7z5iDZS9QJgN+nW6Afr1QFJ/6lngXXssX68cb9kEqjLDIBhYEzvdlRLueYGPgpnNpdRr
IE3RkldAEY2G8zsBnN4h56b/K0Kxep83hoZgd9J8fhyoAHb52azViZyzDVMG8HUQ08CPSVRNcqWz
6bVwGWlVfDqMViyhXfGoqu6q+WQEbwgfKXflAxKo7wICw274mBRhzPmi2vaDAULfnFLF42lFiaja
p8EnyUKMa7i8YmP4vbTePy33Bond+nqy8cnLyy3DnuacMS+Y/nID4xN4ShIobS0l0MbVJClJ2nxy
ptv1mmlbKjbnCnRS6rk9L4Z7bdvYprd9aMlLypGHkQCgWNi7S1NV6et3Piruy/Vudtl/z9B62R6C
L4VKOMjzZuRbuCvrc9AKhzVP9a8OUpQQ+d8I5Ee7bO1lXR2b0Pz19QoNe9DHyR1y2+v2uIKPy7L5
/OKEUWupNy/gYv0vxM8MdKSePA5ICx7JRXikf5o/qONI8oNg0tIdhEjQiuQCL1o5QTBdrbEekWA+
s6UfjkNuW4G46B/SCHJpBh3ykulhhi4g7rcbm/G5iFgulMQkv66xbcWscGrXjAAQFycMe8yVRCpn
neQk2lmsYJk4mQ0Eet9Dn/TxJPTASv79jaw8cZoMLkC7yO3r9QDpFDCiCZXEQmLeIqClp1qcBuOF
CmP3uMV1dn0Yo+6xElgrdPCp5LGuJwnW+7LtzHACOiD9f2oEk3DVRL8cxD0/OHJbV0dcACw7GOBk
giO7s+HhopMDqISlamf3q/LmypXp2r6wvGKvRTx6EC6HIISdm1YiIG62+DB1YwMK+br/3xTMAW01
VNAELsOYq36P+c1yz30mfM854B7R7svqfPGmFEtnMBrdOU2hB4kpQqWKf+T1VQOwjMmLQDkKeKmS
SByOY3AfkYOzl+pLpJfHNHrWTI/CDw0yFZktX7RoJEh9t9c0P8f5Ty1yEiBogD8XJnErW6UmhvQ9
LUsoZAoIVloRi+uEOiLndsySbIHn0iG8YyB+uLsXxXhAOlLhCAZ6baQK6YmPy4jPrtsgZO0SdWNr
7m2lmvKoMc843zgfsrukzUZ7FPYAf4OXJUGClvT3srdRP8ayrxx06XR52YQonadE4n7v5cogi8X6
XTGzJguJ5fz4H7bmXXJ1AnXEZnW4KOhTt3O21WkcOv4jxpUDygEInhQKYzDmT7QnY+ZASYINozTO
bG8JUqIMjsJn4timFOvY5WAf69/945b2uGkCIF3vWysU6szXcci6aVJ/5EVYj4ITHmdKkK4qjdIo
4eQzCT6ltyVPtQNZodKK7sAEbhGO+2dYzTnB4IDgyYUCZCjSiBSIL8b29nktpQq2ly3njmku8U1V
+aa7wMMBtPOmvv9jVxySJJ22Tcq1t70H5l9iHkS2kOeod1DEh6DZFWzMQd8sFSOGXw5Rew0E5u3R
vkxw7cATcxCRNrdW128DF7Jcv11y3U0I25wyfGtti3YYm6ILUxv8ALhUVGpNVGwB9L/GXu4ShS4y
3KDLWf9O5qjIZiRW1bdQKDqYJAVsyGtjjieen7bpgIMaVYFuMmORaqDtbAlQg+dMwIc2fwbJG6wc
ia2pPGJlB5jvwW2GGr9tX8YppL/QdFZB7Zqy0aeILHgkVn+z898+5/9cBDmahtI5kv8zLW5rh8rw
6LiJli2YagSRtqdd8VHpA/DNGVhTsGoQgSCKRbwj9l4IJnYJ4UTPmyyNPu4TDkMwsSoVX2hWxAe3
nEfsrcL0no8jVkFOKQ70ZTZ+5tgWnoE2cWv2FwnlQayHMn7M1w90H1/kHLWf3kEY36UTfwBjsAoe
hRhbnt/lcA2H3MKfaIsa9CGFnnD1IX2iCf5jb86U+hSN1Ny5gcj7Lr9no45dsJkG7b1XJ5v9sCH5
HaCCXqgB2fvJYzDZKtCvnCQYKvUn/rGigOmLI7IgfmrNnePr1kjLQiSO+62Y0BR5AmwC5+y/f1Rg
G0pXIBSO13UgUUlq2qDc6SRL463FCImdfH4LoQ4ERtjBEo3yu1/iGlhbzJumRztKis7iF3upOy1r
tcKRUbWzC8wmGAUGO2GCAS0ylIaSoxEv52mGqKHLoRvwmbfzmwXBGAFhzK3G3vU1QuCb1MeIErc+
MJLMN/2n6B8TBON/izlK1AnbPBcPlhwpCufb2RElDQybvFv+LAR1DPYHOuovl4krXIHOk2WbsDWz
Zrs7YWmJf+qkj9LkxyQIRsJSIGYpvjvDztrwSnQbAlJYin4EjI8ShETlqxrVzaKaatzytcn+3UT0
CY95K+hZwScSTQrzI/j13Tv4gM8Ila3hPilNac7xLCHmrOhPAPhWHKvdupsjg+W0NXsHFz4u8Kae
WHKUDQEg4Yd1DBMCpEuEDu56SEdwB9OP5fVTZgvUSKTloSaLcV7DcWrRgoKnkJpFl+lta7X9BckW
MD6n9bg74OGc9tKBAnRu9mTgYAXaPuvFGJXO7aqok8qQyRaN8FiXh77wvAniM0mrW/vBrDMkqZe8
LZn0EreafnqaYLwSLfP5UGA80fjD5trkpKgxzesMdN9da2dsrCxq1bnqJ6R4MucmLcXF+13VmHCr
jPlQH51NHkLJ9m0Zw3JAePn1IJApOH563JCWpLcnnavK+VT/1ykvggQvBFADKPUDBDmi5TO5vRca
pv6SFYZI9U/BHyMmFlrU1dN270z6qnkup7NkgGHcR580VIrWEPKUhmYMjZR8qf5ivgIpBQ/qMSKQ
JxftuRuGZHNPMvAEWCih73xmmYKwXpWa48aYe5erE/bzAthIymb93AMcUxbejJNYdCAM9lqlDC+5
AX3x6+QTcFo/hi9G4nSWxn8AF/X6t6CS5htCJwrRg9XWQ2BUb2CJOCNL70SBVIUbPCP6wex/vbOH
lp+u84AkeLo7MVtHU5Dk3iqakBy1xA/rKxqfOEhQfwmwGCMQPSJ7QuCtESxl/lgNYnFMLEvd40Hi
x7XpZ8Dc2W9rgpXwJtmqBpkLvmShpBt+MqnUYJjE4z8W1f0yUyv8UFvziw/lrAZ5fMN7F8INgQJP
pfFl6KHp8CcdtKjJCXZC6HL0lM7tRgVBCAUagk/pCsE7dDihjP/DVKo7ryLkkxOKCGfiLXiUGmvL
L/XDO+MIEhZO55PyIPdnoiSqPfKIUJGESH9y9z6rZwReU6YayZQR8S0aL3cGSd1nkXsJc0/mHFxC
A1NIkRWqvEYDvOWoMKFHl0jwOi9GuLo/VvvJt9OXV+5DM+2JKDei9K/QSduamN/VVN72E7zUpRnM
XK3eGbGqTg/eZUBFEgu6baVchl+T21tPBYx8rFgRsL5ja50FJBz6aC0YISkRY2c5YMC2sHTI9oUs
rxOGcE4T0u4cWXON7Ga9nMlYYRDQgSvBfwAVX8RR6gxXGlOvYNsKYdpeL14RzXKPGxKXjIAWHrbn
jqoqrMJNGzgZQiAqA5us4K/cDEHQ4GljsTsHIn0AQOurKoaLW2+LWDMfktWutOgXnaorz0wJ5Ch7
ayO75NCAGkah2g9rN3Nn22xO3JZzbmpz0ZOzErT7xF1/4S2ekEd1iN6jkz/DlLUCdpF2OnkwdDAm
YpdDjJeGMFSugT3fOoyKEwZbT33yL6Hi1SdP6BEbe6xCl3/UfEGNk6GU/3KEmux43zIAFT6L8CnG
pZ9x7j7WPdHhc64LC1mfxv8PNrKknB5XUK+2/DqZiV1yFthHST+iUqEhNhVC7bhtHVTjRken6di5
eyZJVapx0SbX0lDVQ0A10ljdhC7ltOn6rz7ZV1N6lTGyxUx6lZ5/Goj5pboJMqex2BIl9OPBlMWA
w9Kv8raCtWL4wtBFzLJspSuj7G9Kk+60j3oY4OUNV1e1iium9icpjzFZRubiSJW4i9Hhs2+oLvUL
lM+22ZHiYEjPePf49nJGpgd3JtaNuUCtAVPltwmOdIMWfF88NL6qWtKurLIlZk9DXcIZXVbmeOZO
hTh0Ae75xYGv8P6NEZb2cyJjgtDrDLzmdUucVqa0voD03LpYQYNzhRljU/5bm7fq7eoF8FNhg9xa
qZeenLMcg4fumF0pDQsjBf2zufXzlWFyy5Uz2Tn7bSu5vr3GnouXXLepdf0kH9ey4DJAJeSwbgbz
mhrIDRNf22iS3Gnen3kZ884wvNLorTvMXZT95msUo/a3wqJh7Ds5djwqB+QU24Hhir4riE5Ndrcy
Fw5f91QhVTy/CqpxMLrfulEQr5yVvx5t3eduAOz4xFzve5BSKY+/w3w1tko0JQkpJFDIiC7MCwbx
k+R7DjYZkglj8WTo5TjmbloUTB/LTqvSR+7IUup7z78i/wnDZ/PHrii7Jy46BxHU0xB3sNirDXWm
+H65yUi/tPoqfT9MBxxnQe4Mx8HVTSKLVRhqCMFwvNdLT8mC3lW7GREA33tGgaR90/6vW0JYRJTi
6NpTTToXEYWNfXSt9OsWElIx7wgfNgALC1X267Swtu2Cjm5mwEusssqru/iiU+aq1MGmc+F8VmkC
PFKVlgio7iWrXsodZ/yqc3RYAazqucBHmNbdjla6neJSvsk3sgfdM1CZyBLAAGNyAT316IlZB5sw
t3CU92mIKn9Fc+gD9XrnNB3SGxGiSRLgwNtyR+Mufvpza6qPeTyw9dYxwYHJWZGLeVLEBYypVPK3
7Mtq+FjVOM7gY24ZpALquz0kL5rvaSkCr6LKqNdXC72+Ufl1yvqLJ/5AjraqJNsiPV6pbtSu4Mjt
Y+vbm2UUulY780pZUKQG5f7/T6iiiENUsfYnFO/kj3BqZohl2EvAYckeQHpEdopLceERyw634jj+
pDf83RICtf6k3iL7116SG57pmx3dy72ACkmU8T1k0umBRSZUs8SGxrxIuqfv8dKvbNakhpFtvNA0
bCLjtlDXOM/0ua3I3rSMErr+5pbOt7wBRaP+AqeT7slbtOvNjvtJYVPFXOJc3DOrsoxvrf5gLjhY
iE+ejlMn0oxn86xwkvKI2lJvWE1jmuQw191kQNtpsGZfDnA2PEM8/dmsorOZFcIUP5TFanVa/hKH
0jWwncUcwXSyZNd7mP0qWPbWpoJZV4AnNbVHyzttrW8+pSmFzgecoXF0zIpfKV/IkEahqidvsfsP
g1mdqt2bFfluwc0RbUcggk3mBkYUE0tm7O6P/PAnALyhJWLlCgGoeFI5QH9ZXbsOJSR19YBNb6mH
w2FgA7tkFHTZyrKzZurlIRz1ItkiqmVjcHsZ2GeYMCEyj+BWTgT//hPItmTHnqSqdW0P7jsjb5en
m3a52KG5oysR0i1JS6xbL53aihz+WYoimW5o72PzIptaxnFCsoHSmyQuycYsBO+x69uJDbx7grST
NxSb6TAEcY8PJGfBMs7MAHd2E8if1fWgPkQ8hksLtEx3x0REDZONM+4NRH+Ol2EXE52EEY3fEUbG
6yTzfvpO7TPZvtKiZSgZzfYCCpbTJ5uF883SajFYV8YYJU/MjLbm7OiO+DtY7/uFpUrT1oRD5TCN
chnAILqBfyqrkEse6WXbK4iEoClCDtAiARNy4ZaYQ2ye1FBR7EsIm4aqghQgsnXEac6Bn5p++KyZ
aO6lzbZSBjhhXap0n4rfUp3Lty6L+uSPOhLEj8ZMjMFN9WTIkDW4rvk0Kibi03z1aab6Ia2Wwmie
FJDEU9jgOyqHZDoIlCAR81DkLfzAXvofy8jBuX8u47oZ3m8FhCa5MZd2N7DFNmBBagHFZw/LyXhY
fmCIa2WqIXA4z0eOqFrT226nyYk6tR9x7GQKrE/fc38xtjga07l3tcb2BoYDZdArr1Hsz93s0qaj
5ZdvEWpC0ScYmQaDOtGD3PQoOJbMXzxCNMvCKXkAEHZ8C2Ili8oOH02+c/zLkA/LZyoSAn5wuzC/
Kbmt95SxbBytYLGENlb32zLhsPb0XGWD73XRd17g808tVSsidrU/oeMHVypMLhVXYgn3m24VeIJh
hDDkPgtXM7CzBY+tejUPKcApJYH6w2GPJCfIITNlPo5XMbzmVpwfdAJuGmozyn2memiZ6m/4Y2a3
4DwIQXMvus1Z4byYegQLJZBokPmrASc5I1xXHzrPo/ACaWAOHekuB0PtFWw0TlzVMVDgG3nbWwOb
z/AwBFvHEfM/GFNHb4fFAAg0SURGfW4J7kh2wknYsm0qavU1WKWtLmktMdoPqUh04179KNZ1A6jK
c3p0BbwRnJE/V7gflodoESRQThe+9j+nUN3NbmuchzobBHAbML3o+SdUB9NgeXkWuq8IRwluzzbo
56vOAIgOSS5Iu6NIuHvwv75m5Fo4wu9I99IAcf8YRrH/vSTaq93hNQioYg9w9FfIcrntDzTP0e2N
xlB4gTanL5rDcIu3w7/isXmEc2yAn0ekk5ozwwMhYNw8Xsp5d4ciiMWYkVrX1D2zeJjCm0rs83AY
HbBpjwc+kIGaLDHpA1RlTgNAek7YY4c+AV9WgH11Rc+uHlMQwKep+qBoUOG9A6oYT6oU5Yq0bQRM
8rRwRsRINk/9hP6PRXATHPRLJwW3KXQvkcQgLZBvkZ886tmNuQgOJBLSRNuoHuRXII7LAxBnMG/G
409HUBFAqIw78AEv51GCBraOg4wwPWG04lLS/4pUgn9r1nzYiA9B/RHhNhotoVLs86dFEB4+6zAZ
zKtatz7BA1llR/5C2fb9tW6sfN9ZI4a/DiKAy5Anj//VyubYQ9hmh+ZdHARTtMw7YpeeJzCFZRqd
WN/AqqTxEzC2VuQap0aeallv7PIa+Mo795I5Utmln/pyMBCdoYn6xilDNhAEG7QHqeHjvJZGF1gV
VcqHlzUATuje5oD7JciNONZazHZOtzrtyIZD9abbXNNvIgO/R2dPF/v/kLwpPUzRozmzZ8YDcAdE
lqE0cOP1/sQt/7m9EQ21zo5u9WCx1jSX9Vm6Du6rBxFwtkToHaDPhhSZhhRqaj5XB3QODVCN/G14
qIYTaCkPxVAE4L8l+Gg4Z2o1AqhFVH21MsJULa+EKDPwE/GkdlEU67l/AHTldY7b8exMUWlcOPwQ
D4tEgd/TMA1UerV0VrVvcn+GoiQE8zFaqHwsSAugjtPNoRQ3+D/m6s9g2n6rvC5U0ngBKGXKae7/
C3OdOvh34ThsyrYZnVfQK82Tznr59K+9MEKjlVGV9g/gjGBLL2fHZuJZWQ2R63j9hJeOGgxAsPmp
NRSSFFOlZyxrCIIbzkPbfzG6jupQmY3o3HZMdJOmQV59kPMLB1K3ZXfC1qCFS3m9Wpmpt8/MmK0D
E3BS74HrzsUeLdU3JbDNckS0OHelrSjPukbyCVn4ZIhDaTHo7twNv5B8S2SeyOmO08cI9eWqtdf6
N2IyB0bh9/SszYbdTdTl3KyFeN7JwqVWMv2C56KZsurQhkCtjzV6xlaJ62Qa+G2L+22l+GAKTlRG
QS0AnGwhbBLueDwgNrXlNheZ2oJvWVoQ10kLVMIu2sNP+nfLqdUSf80wn6EcPoaVw+Ve7ssIOZIU
6KUkV0USLVP72OhMbSAHNPBJc/hBLKD1LWqm7hOvVUS9k+s1J35e0xu8d0SQpHNAnx5OKpMrXTgR
VtSHQUTqdFKVoCdr24AcfH+cWX2T6pTh3LZXPulciRyuvLQNvhWOhnkG3TkRfMTXfEwgF5jWAIOm
SSSaGJH4bifbz1WxnzfTRJdZL7vPz35XQ/VlaO3Hc3iG6f9HiMWNAZlGbAVJAXOutBDKZqDJ8wps
6yj9bGt4B3bYjcarvreD7ivDwspXHVe3E0mCROpmwCCDwDzXy21CBXUz7l5XD8zIm+ymY7CDrxl9
v+myPXJf3U1iIYMlNTWnM9mrIdA1s/3uOCUd+aWNF5zzMQmkuonvABmALg5UcRjl90Tny3Ds3I0w
2UI10FYrEMJHDwV9+xsH2KD8IP6yrTvxubt+J8z0RZL6JK7WDdZnowmr49M5Rkzllar8/t8lO+0M
P33socvpXoJd1zERqsKvG3kc1xHwDAYgD9L5m698RmiMzDvRl2nM2pO86OoXgMp/k0RNadyDFlGy
mk3qeXEpyIi6dMjDN2KhiCfmxGo2TLnMWyb49UNR6zOKMLu5ZwFuF6RwquuJRjDpJsBBcm0IQ+W/
eMXkWoa6+h8Gzk2Jm8hqtLvKcTz7pfSHpQCiMBxygx9LT/2VRakfbw8NGUEVQYRv+XG7PZqC+xdx
B/YurhTyyH0Lr4JxWAvvvp9yVY49OOpO79AjAO1LBvohaVOu15suBl+jxl1JyT/tjvrb+S2GkyFQ
KToHsCaqCZ6JkC9cE+/lX4J2H9BDmy5hQkI4ggAB2c64lwDPj6+OMbHDFbjFbHfqpaAlYHUh1Ghs
WJI7fJOU/2YmU1zOqdi1x+H+DuHC31dw49KF55PBA94MtDP0+ie0/44NF5PVkl4v9YuNXMFDwqEo
KmVBTokz4bXds2GjWMRM6bFBcxVhb3zYXu3IphR7wkK8CnCTuijZ8SCMx1WT8o+dGNkje4MN0yIp
tZ6piQu4exGbQ4VLGiTtJsIGtP9Dv1ZlExcMepW7H236pKFkKEKdgqJHJqpluhwDo9MJkUga99lu
9LWCk+k1IhAGUW1tiOAU4Hn9nhpQh+oPtvSlo4rm5h0aF8ws6vA41B1JnxUSrDL61SzuZ6GZJZaK
QTnk3s8WCKfBdajGoENpOWkvxGpxGB5oYVWIXQPhJZ6lYVJEB73ewgocCUnESmg3s0zhulTk88ZI
zc7zi1325vICLjiyCKeKaOvus3nofZp7Ow+oAFDZoqoAiMBVke92ciMIb5i/7gSWQtbhE/dNWOhA
oxGSyxi9veQJerygQVdDZrm/AF/S8Ag/XNKlGFtkXiBGezHQrlNY4srkGrGczl5TjJdyTJF2nJKN
ApN/J/DdffwOSPPHgHIOj1yJEzygyHZ0mOEkkvd5zq5WjlZyc82pEkdYeRbhxaN7B7SC8rMgWxNn
pYUKqOpwDJxY/Oek8s5Lz3SRfjND3yqmcARfM0bLlfepUYJYrU81HmKO8W4c1pVu88VYasb34STx
H79cmO9deYZiAnVnptqXTAieEDIaSeLc0P0/9ZnK+UZFLepiP5QuhhrU+ux89vsLPp7TclwhTVbB
qN3A+WSxQBGKe/arGV+K3GHOEouHS57CrX4leo0MA4xcV994y7ltQL6yz8zVpzYCCTlW8Untz8MD
MDQkT40O8ULZzEuBY5hcSdHzJDO8SvdW2fYtCbz3okFf+9bBM45A76zihIQwoek2iHwxd0Ozo97e
5LeOhKuOCPWz9A+iUyp0tHNepHIlXY/Txkrx6UB2s1cs4ICgjjDY+0ZE11khBjDi1YCitVhszdxI
1RJGgA4Xv6VZikVV/uja6RWaqWHv5hxd+n9/6YSNuXynQEc3ZrIicwjmUM8OeaEE0Zd2kbPAxF+c
hnYda/zJ/ng+iQQdxUnAdgOxmNFnjdgFehwfbBuBmF+v3hukfsDVeUkUZGYDS0HKlwrZH2Yh3SI4
L6ErLwFcPEt8srPmqjBWojDu2xdrwigU2eraBTf/6QNreBvaY/9Wb6yMEdrRTWzj9SrqQWIcpZ8F
9qH+YuBIgImG4OwvigK7q1sZLR7xrY6M4UBgqgASoVbaP/69lh8/qngquKvuJT8SkcVzCQU0uiiU
+cuKha4TT5EO38cP4lNHMfZf5byr6DC5uFclmrZwsGvQltSFC4/cQxHPmo/BRwLmCZUctxdlg6lh
2SFr7QDnVBKXCcVIFQr8nAVdWamYHH3cS6zkDTKELk0W2R1ijaG/g9AYStuYisAXHUSMA2NgbAzg
7CzEuInTHWV8PvQ/DqT3GS4qOXcMbnxagla5KfMayzLZSx9OcoC82kopYU1Li2HoStoy8awlO0mP
2S71/+g0aaHRs/mMgefOFCzi/dcXyfeVMtH1JSsD3bQ3puj5Q285kUKVGwQmRNBSsM/4iwZx+Wv8
LU0sq/5ANF+f91mM5cDoGvT5gnF5br4/hhzstT1EuCMOfDeyXXHuzD/oWxhkNECTn4kNtc3UW424
4Afrjun5yEtcfnZfXAqS43jpwRX7F4W8rFKzjajkkN6zLQQXOYCz05EQW/DqdP7Si1J9DKxer9PA
mWBMX1lzMUpnPmLW3BRPOJaJ5HzNlln9zjQ31i10JFMTu/FAtHCNMDTbN9gwaxP9W6OSphmtG3+L
OzqJ9R7yvTjtmA9bRVZYWmD0iPSDdBHli31Vhv8TRr4f9QxGImvEiTiEu6SRUO/j3RD+XmRK+ZnO
1fqE0IccvdZLt9upL5aVfFsT1XWzyaknu9L/U7o0IJ0UvkNE2VEbpBXkeViVzK0rHav5o/8KLLbv
2YyYrVeIPHoLmXHb3qBOoilCrIcjzUYChIJ5ghIjsKmPjMdtbnTMyq6kjcH4AbZl5qJ6pPzluDMa
MjluRjB2frHx5r1L1lCn4b66Do2yEVEXdJH5AiZm3h7YzaWpcKv/cYUzay0kYpXtGx9Rq2mcPoHj
GKSeqZhFSv4Vpe88+liTgvdOdYFiXUo9wINAXRXa5C3Pl4Qc5UUxBEt9qQaGx+FjOHwYVNfB1jIw
Uf6Q0dVAerHuey2WI4mmF7ftnjF0dJaCdUUbtcvDYq3jfiLh637evgq0QCK9pnD1iHFJwEzSSlUF
r6IYy0oyZrur4DUj005l6vSceTg0CtxyOJngUv64LOz/TEQSww4vB6lEtpaCrE3y/cEkLDwQc7Jq
Kl0NHuWZp1xH2NjbfKrW7F8k2SwK5FVnFPoHfcGQxKuA5b8o8bho0sE0FDCHS8K0G4g08kEZIPBv
xDXL70s4SnlxTeGZ6ZYB19vhoV8ipZERyyp3f46Dm/5Mgar5g1A5voZcJC91m84guzxJleosRjZi
tiM20DoDDp1Fs0VBlPWzXX77TGUD5KwO2BsLlMxXv+f8m/5DGH7+1qYAeGdA+JCuTEulCHKxLDi4
P3ZFyb2FB3Hun0FeBWFovhTCQhUkoA3wuPPanwyX3bNRvEGKkgqt2caIcBEfTu5TUH8fDDIuTzno
fOldNf36VOXwjurcuNdKkF3VEbhb4NOkltevQ2ILZ+W6aDe8/LOMM/i6xLGFy4CqBz32JxPp6QCt
NR3YGVambsilI77wE8dAJuL2oJvdh6BeHzOU9DGBZobFSdGiyCC2U8OrPYXxqVgbc1kxvZZBLylc
5KDY3KLs+9wI5ZO6kkiRt1cglBcwItrdHQfnejFLMEhH2Vfi6z0hj2dGiOw20oMYzEv4O+NgxElW
LJjHYTzAyK6yMq5SWHRKYYHHv8nAgMEE/dwmftLAW28pLJV89xXR0XHhZT9TiSXiSUUMMBE0LFK1
9uGpgCqQk/1coAckqRhexomBLLppONmTcALf05cPYep6ZnHI926W9MiKPgis+SNkUS6J704jcKsg
oRBTw8fnufZ9Zpkxi2zR398XJZ4Pm9IjnRBmCmnf6t2Wb54UqL6wqZ/MZuJcldH4IeI7dn4Pi9vT
akmahra5yoyv/KQkkJu4fYXX09l8l9OPwwdWx511ui3awNyp6sxfBRdiymwstKThIvtB7QcOR1d2
Cmq8rW+zhgCjUaHBaNXFsm1yI1+Q6e/QmSt+zwQpMWXasnEG3EF41fuCYOuHEbFQHRUzvBGAJ/iU
Kr9ampGmXIi9oEZmDkNbukMfR3wd7nHhMibfG0CBvpZn8mLljLASKF/zA+u1vafUa2Oww/SYhthL
0vP0VOdXUHIBCSwqeNXOXQMSpLGodcT0ebJT79+tg0wRVDx3RBDYBtHopEX9E0PgNqqdhIXbZFtV
EMMBDxO17VFUlkGH4UAJneZi3CcH7sRPaiiE77llVtmZd+r/uhvchqh/EEg6R60Do9oW4LcVj0K4
GmzP7IWv7oCEiFKWBqvHQ9k4HVrelr3JiZqhMBqaJYeGUIPx+o0W3G4JsGQ7ponTZnsrWkl6S3Io
SVWsbLRspQDkxJu5biLRlQs1lO95N4kNW4ve1pYpbX137Y0rUuyIyBqPWolaV+xyAJj+4ewFbb/w
3pjuX2PcZbF89oF2zY9P2Q83i9egt9dpvXOSN73vV1bsAN43iwqfj9+S9wIe+OOP+Paffv6njQ2t
r+p9zkmolt+Eu+rYlkeTnBXrVKVP82YvW9mhod+JRB3p5aExyqcjN1aMoPdjBwEOqNogGJf0C5F+
eCSXNATO8gnbrfku/IH/kDRUcLoq4jNbS2okZ3/jPDuf5mFFfHu3WDxBam4UUpCd+ZmDlUE7Tz2k
n0xQTYgyewlVY6OvLZf8DY/8ycQxGMLD7iaWA6hWMXyI4F/gY3TOrPmKa/WfV2gLfSWHG5Rc7PQP
Bzd1BWzajL6THwWzHSxoSYuhOyFTpGWTnXbEz66SgNETEjG7zTxfHSXUyLZynEt16gKPOX3m2pXI
HFyYFCEkpL/EXFZZrEHIwZ1kLzGd6zckfbe+vwd1P6uP95AV1GxOwn5Ho5HC6FIOtQ/FtbrKjgqw
EOzA4oDaqX85oJM1gCb44Qq4pNS3YyHM48WYnMgaw2QfqgEKUqQqWjtGi7iQUcBsjMchLkveX1jp
BFZujg/5n87yyRmyDv0k43mfcsYpazog0ArPzgAPXMsldGf5/vuxZiEoqrM5uRENO4kbISwr5cvY
cA1kBDBOwxtb6cEis9QxVuktPndpEXZXzpT55yx+OOygvs0SdejcxlCCbY+6Ig5juB+tLYx8yZKg
WLWsqAH6fa2VB4/UxhbqOuz1vGOhl15WX0Pn8BougDPw9/S44EDwpRgY60M5D5atalZnMGUTWRX2
AVr/q+weqbD+AkFIkbfTJ9xwFFA9rKlt1bk+vjQvnOXfWrAcKw7JtMNpsomDCZyeE4Peluh6HufO
nE7hP57rjP9xXmMw7MEfvvEwCrc23g5f3UADWHURn35IQr2LaTCtt7KtMp+1JK1uESNwbF8bG4wv
sy//VWT+HMnq+ngmM7/vovjf5918n2HgFdJWQ/6I5E/RyKMjSZYhcApx9dND/X+fV3PYqDUxD+mY
RkXk2HDiajtzkfqCwD6ufc4DTjP8feREA5h+9G235dJQVYZQxNEs02igY836jfb+qn1GssNRqmVZ
x/wIUAadl11xdkQt/MZieGZ3QWRtb+FY14ZhwDmaDxaKm66RGG3QUC2Z0QvUZyap7KPXHGyN43F4
BeYf+QSyz9guKK+kdSCedj6UVLz6tdIFyxvVmer0q7KFF53Rw27VRIxGwu/UX1rkDmoFdxyx1Yiw
3SZELDQqhrU92NMrc6fbk4SM2eLwjeuTVJVVYPlEeqYa5hSq6ODujcz+3PMKPl7ByFX1FU68vLGK
nNAOZEU8i/qjIqaK+wORdSfo0qwYGjq4NjNPFtANYnT+bN6Eae6plKN0y+USdjXpBIjlf5yetJ3M
sme/U40dgSEejbMJVlw3uWySIkzyFAYPalUxlvqWDM3m4Kq1KKdSZ0P5haSXlkjYWMMvp0qhwQkA
4t4yqkICalcFr8bRbe1TQGOtF3/Prwzkd7PRFIOkAv69ga7y+PY9EPAbN+8U12vcrsqZA1/T4eix
LLpZXOatkE18FM2zn3sFOyoilD6BnfEW3S08Y0ckpTECWv+x5YiWfGGKWbJrySaHmROcPnytCe4I
N1eOVGjaXhUpSAY13HSXmSji8+/WbJvxvD4s7C6rmacBojDOzR2Z/UM2EPbfccf1vI7Mzgs04NuM
MHoS0rWgBcn43Lenu0v8hiN+7dtEsLwMGWUjbXjFdG644buqo8ORiQhDPQHKRgVGexNXQ/5qn7ku
VvuGnykoLZ+K4g7zA3jSgXBs7SbdqEIFCfxOFlLndghNRw/DnzHZDmubpvWEWKWG7ZeK0ivVCJUi
/5Rey8kuRCC/Bl6K/UZobI8gjWYOJ08yhpt+66lLY9z6w36TFKqKLs2+jD4ifA8duQC5NzatCi/u
NhYmnPWO36QRNmDVAw7bmHozQwb8wDxB2GG9jSVtZZIWzc+y0m7mgL7uULniTfTkEmHPoVt9RE5a
dV/20w8kf8GKo+Zpnkcju0qf99aiYbV8Vk2y6CWvoz87ik4ktG4LBFj98u2t30/2LPsbhdYb+Qe9
sdWWDAC0Q1A17aEjDjeU6R0+7H5HeyvvnLKpNJR3IdqWOsBuxIkUL0Mipdd0mEHhQtErs4d+2DcP
U4tI8osP0fU30HBySUzIz/YL1F7vy0eb6mhZznwIL8GZWo9qCWKfXv//OrFx3csdrf3jOVqij7SH
7GNU0Lune9XsE+BilLYz/MJlCk4aQpdehm2yEyGB0lxgx9efGY2nCIA9qFNbmolGeWs3LvcxwmGk
e0OB+BCfSvdVVE5YkGV3+SkjNOkBScTJ7XYSboU9id0DlAIzrYx7BZeAj6ICkLwRgMvYSx5u5bjp
1eLyXz3wgZihNsqkAOCl/AvHOjg6cM8R4evsjZ/z5gltKRgDnol38cU6yKAxA5m6rR8AApb2wvt+
Zpp/JeIrt0FMveRhdNijVT2DCprIjX0gWEYFXiUR590aFfR5nV29m0Bc7/X6c0oIGJI4kc5Uulj3
0Gwj3VkrIV/RLjWMkHzzAsMLz15khTnkWfJp6LEbLLKg/2CjKGixo4tKHB4B1Efca+hG1MDh00RB
JsbwjRWykBi6afuwX01Q5JNxQnI70x4MvPPAvORt6ysmPjOy9tFcO6kAbRK7K/YR3ANwE0QJcwcU
LHe4vC3wU37KpL9KvROgb9yIV99PQO/4VkMgqnNa4HKPk6Z9KSi+jY1uk65IJuYrq7TlH5Q9O6Y2
yfBPJZjIZKEWVafUECEzA49P/X+y3gOPRUM1Lxyj4J9tLnRzGFS+DEsuj3BpOR1LWM0xHE9UOTMY
DdgHexzMHN5hTTOMZciMxW0OuqWK/ORVuLlyRAPE3OoHqJGJmTIFC5NWduUWUuq9FB9sD0DIzvB5
oKV7Gh5b3r8TTIzzmOVsWEtA1iBPCDsYItGkgiELtYAnPUoUbfS35BnMx/YEL9KnM6cEZUPlRfhg
J/dGxavb5xju3vPnvVeD2ViQp7Jh0FCmXWJgmNJj0ntjIr+fYi2OWLXndwxFCHaT49hJ8l2dt7lX
qzL9lRrRs7pumjq3VuQQG7K7OrZ2HVr4tP2fKTeO5PIIWkuMq251/Pa5PvmkoDSn15w5LA7tyTjk
HkTxcrgdZ6KpIkeigGLxd3VA1trNv6kWAspWA5v7/OR96UitUPHS8WWIWbXlgBhRRl7t6P6OjVNr
xkmlK8QHiBk9T6u+9uIHxdiLB5zmYEXY/Fq+qyy/or6d2Br4w3KU/27m/1bZZ84gD8Lwr7wJpEm8
C9CR/qsV3FT8j2s3bgJjqSytNi8Na6lcgURRrLn+tRRWEENY+FAM4JFIiu1eoeohtEjvpcZ33hB1
SJMWGzfmckUDLejelKKEcyF62HvFhNpX+Knf3tdqVveqUmNxFhuxZhJ3nzwMFS6C8x8K0z1RKB8u
x4gR3zQKvYuzFGbKnLym0vOdmEQnCZosGHWe5gVBeKtnNA8vg0DQpwPONw2T8njEl+6vSM+UllkN
Hqt2YMd5VhhNUxE5P0fdSxThLmYPXR70+Wi5/uuOYffSMB3J2kmKKO8iNu03s0jRweh9OZCJOZue
3EIDPDDa6BjQL3JXA29HCLW0gSDbNvQDiFfqw6GoCQoJZetP/O+evx2yU63ijJ7qHwge/eLXrhdV
dbotUIQEdRkGv0lQyHwcZKkJDt+IYpLRkeZRmTwMVp/vGLJY1mLCfOgQ3HJZ96kG5EAQY2qiEvW/
1emllMT5rDcSAKNi/zUA/zmM4BYW7i1ddwuESHcgl7sGKCzCzWeeX3w2+2RWMPglC0CkjnD+F7Ti
Ew4lFDzyQTUQgkuTRIv2km4wlaXJuKXlrOhq+uWe6cjUjrF/yTm/WoVLuhwQd+DSFtZMUYLamLqU
OsJTJ6Jkh6bFtvQNGlw7MZZRirqc+IBul0kD1CHvq3QoLyGlxFt7jU4w4XPF765SaBBeE7OmVrR3
HGYUdEhHrCGxMVLFJgTBhWVaGuYNAaBZlMiIsFEC++U+Vm5D8s5uFaE0G5xTP41Q2aKNPIMKyvuL
4emGlO0zve8zFDzPTUTN3IROOWY7IQvJQR3ikI2WLLuEnD9iozglVkZXXf6SOOTkob6HFDhLOcWG
zB63l/mrTvJpml2CXYVlb7R2zNlqZxYbJnTkkAFyh7zZGpRrZzkz3REyRcD7PcQDQqCW4kw8kein
nYWJ4ovvnA2/EYKZ/gfMqziNumQDKP8ift0VzLKtq4W8bsM9xGMaHkL2iSkx/eSeKmUChpewSge5
QiIvy+KrwtHMNuD3lYhlN1+C2FjNYUlMWm0uPC1CtKy/hiIRltJaRl0doURNOR8vSabXFJnKfJVM
pjuo0UwzCL66Tk83g1YgdKY/t8+KaGWtMYEwI+ZAKVgi7HcMzZW0IyefHVGw9hpldEUDhtvtLf3R
nK/EQXQZCBv8LuSVFE8yxR2eIXtD8kc+6FC5yMy4JBFzPyQ7RFmG8tSgJTewKchT4rgpfA3gJOGG
jfsns02vUGru5+h5Ihd8kEOJQWLCtG1DPB6g0gl2jWrmnjTMNv7LOwfLWacKeCZaM+9osN9FJgDq
NC9qnjD+Crol9w/40rgoFhK/TScybMfV9YbuP9YR9aYcFkwJcN1jAQ/1hItEF+6g2MynMyBYooNb
Wuu1dtYxE//IaB514B2vrbIFlBg4U6u5PceQYrP+iZyuXUYqnxBih9l3Zsq57JsoRq/KA5pcoVcA
daZP1L8U28lnJWMnJqJXs+COydEcq2+vHKdW3waHo2V4loo2VGF4N0DB/8fmMgTwOtPJG8zbEhhS
qkblVKu0tghRIHonzSpYk3hfoTVIePtgKURwOeKIzZ7HPIZc61EMRA0V3J/+WWpFAK5DowdnGPaL
ojIhulk6Dw2eZ/osKN7avKjqRm06W0Yxom+jnxVjnwAE6CUVWPjkw2YlBcIdYEZfqxoOr+ufuXBg
ddOf8gSelPgNwmXHYsl2Pw+LAHifrhU4BzfBL2vVDau0xymlvF1qdBk1IjCUPo/Zf2jY4FIRBCkO
5YUkBsw3Q1wMlb+LV6LGlRQn51ssyn278DJHXN9wVGADfsSCLq+lHB0XE5EzMtWkD9R9yAyhNcnR
Au2GpIqkvvojR9eAiEHKYpFESE3lZQSlopzOoDC1T6EpXhFG00IiSVaqMrhBc8c83Fu6U7ANATXN
rQIUOAAfKOCddC1m73vS82AYiHtIch7SoiQ9OrZeftLIlBtXMTJPdw/IL+GGNAVH62BHuw2EL8Iw
eDYTNBNWet2d6q+8gyQZ3EidRsKsWe6kBbjAP096jn4A5kGum3smesMpnABy4t9wHqzSqYzSJ4YY
ll2eBMYUVvcs6zP0lK/Ta0/tMdW4ysjbsoAvffMsEP/nhEA/ju7VsiGy268WG6zQ1plUhWqZX9+h
jdOU3OWRyH1fcKzJCvBdjP8cCeQLlHpXQ1jDkOIAJGNUN3EoZLU40MFGXFKwO6ht8K0NgiWG2MTN
ak7mb/uKMviKfKjv4EMDsRRqHBICcvh5ig/FNVGyxnZpCtUCtlqkoio42GoBX4I+BaY278VDIJBa
FpFDbvpbGDwIXAzarRMg70TAndqQGpt/Sb4uU0Ro1MaAndjjvfTcuS3Uz8NdPp+/gBFJLpYWhDdw
DEThRQDap+r8B5KuOcbTWdJbzZmUJ65VLj5SAEBMYFKyQ0yZko1xMbWAhIREprSx5KRJG9/u5OyB
pKdVlBY0nuOG6EB/tGApye5gj4R0A1oa6GkMxNnC4xUeTRjq3yLQgqM3ua1ixcVkS6TmyZ6FfXQ+
1a2O6SUqm6nl/5JbghXe5XIKQxKm/aQkAnXQ52MTdRL8A9FiUhO7dKXN36n/lLKwdqWhQALp+dbQ
BUru/7K+3wK7fPL3tMhbla/8hN/OtqrwGZx1mgQ8cs7420NLOqKlsn6Ff1S9zck8mzpdNl4dUN0T
wd3lVF6NvF0kSJe2dyRoZ0ox9YEYBmY7U8QZabH8zkNMtTkBJGHcnSf+RoH8QE6euFMgD0xBCzY/
aju19vjJhggPzP3M06tUnAWriAcb5nnEhngOQ7hgPmH6/5+MiA9H4q7cwpz8sk/58m9Kn3Mrlznm
r7VLjQ8H3zPC4tGOJd5v89eHVkBnqT8d25zoP5bqoClMtWgIkCfVJ/3q/j7/PDEHtdKI1rkv2+Z8
KnWtMukyJhR+ywHwvaXCKTnuW8T15r5gyn1WDTEv37aIVXfsJKPqdjNuKCxIg7SK4e3ZP6xhq7gM
hPMW+dmy7cXInoHPHanUm7RScWvkWSdypv/phWvopDyUNTEjVh4MVFbpjZzj5d7aV0htuQn71Epx
QvdIFzoJhThRF0V9R/VxOlZaAZTzim68NKMi8fYy0sjCbLN1v6T2H4HfUlvkMNCJyuQlGLvHyF7C
ZcEeDrI+o0Dvmk1Zyngy1TLnTvd6Ep6kaTKyn6iO3HUt75M7JtJ3QkpbtQir1T+rJ/NugDokGNV8
fczglpyu6uBC0wa+nYeiGZutsbWCVdSbziR5MaGeDOm8icecIAhAKZLTGTnNr8+tB/cNhPz614hK
pVFom0VZD1lBidUY5F09qDzzU5yVWOApx/C4LD4FXlOPV5AYmz9LACezc3qWGd4I2+hVysWWvLzt
qXAwzbOcH8zu5KEr+o7lJQeCinv+NO54ahY3tvjWV0bTNKXObGmuTfYJbYCYmkrZJxOfmdNJ2eQe
J9HYf7jKXHmkdLP9nQGM1zQmv5dbjWXuNpSALNeINnwRf4LEEabXUhd3i246mviSlE6e2QV6JQYl
+QV8ykZQHk0rDAYeerU1P4+eEGm3WuoRQhuY5CXnvM4OwGApj9tQAraOqAFGmdTCYKXOmyOeUUxM
YiHVxRlPriZGd4LId18KJRR17f6jInxeMzqa583l4I9Ey8QACmlzg9nncRdYRrJqBI3TFi0O2pms
SB8Apj+2yg9czfVGUYxmeYkpxw5LtLNOSFZIbMGmnd5K1Bidz/1hyZXdGoqTytcvhJ3y6henL5OL
n4zw7qneqlxHZH2hx9lfpY8NamkkJF8xXVpM6af5ILC4ZB/dyOnEH0UOZlWwynVoPQXb+lS7zmFO
me/xJNlUOha5NKsDvC4Hv9jd1CVAMZHuZqM9qFcBwVisd3HKMiEVMmGh92zXC5xirklDHihu1yCz
M7To7KdwTkZofiCJHyER+qTm3NT46kxxTPngqRUlnxkpb2Aj9P3JWHVTc2v2lz7/QLz0MAsTbLMI
buznMi1tT+Vo6c2UO3SAoqPWLOSXJqL/+BtE5iLmXQVWDePppa5eOQP58vieLkYyWfaApqq58jwM
8ffuztqdI+nmozIewBB3SgEQrQ72/bdnhRsq+hpemxK9IUmeaMRk9+b8U8opccB2uX2RDFqC0Ch1
8kEuZbA4mtCqQ899XQfCZDex1E3wtTZqizqDmC1f8LvvNErfly6VSL8IgfmxpP7sWV7I78fB9EN4
TMKJa4c0+zQqXcMyTJ4vWiomBHuhxx0biy8ydlACgmd8wXPrgVhGRDndet/QtZyJCehgcBWNju6T
EnmrZ8S0icX1NS9DVY1t+CQqZ8/XGcwj31mQdw8DM81VOW8elptZBPdCFbiW1hxk0cJ+mhid2hp9
rs/9Ky4KkVw1K47N90eLxpTr5ONYTaE0EyWh1okn0moqFWZ3sHps2ZbFWGMQilt5eLHwusdNCpkk
EqhkKrbcBkwYJoI3aO58uORp5TYML9r254w+2KLDLpi/YHHeLS0HHCuBwu8Ig05HSmXHEQVdoayH
ajKOEi0U0tErnZn9EYqPFILMuO1h7IZZ+6DGxIzD/s9KZw4xOr7rKTjrSzmcHJvBdGjMY5p3aSaF
/ww2W3FhlEn7cPDQO4zlEMAfN/UmVsw4KFywH6JWT8HF8h428m8uybE3C3GqWWmC5LJ8UT1Ebaui
X7KNms4+3NqKcg5TudpJw6w2MccAfNMQFWhg05RK4yClx7uEOw9+DK30McjukKkeNisFxZNHRexz
575LwSRQ2vpx7hU+QVupgjr/LPiDKvPucO6eH1oLoJxWaTZJC5P4oPYsQODLpx32JnLyHnW5X4c5
oum2HR62cCUAahsnb/TompAxB/9l1Z2WKhmvp/jRiqnK0opTHbri5rn5b0Fh1vjOt2CPYWB1SYbi
DUNqm7W8Fl67xXzGlxJEgpKpMoIAbOTbR/95vyZQHJGWUGJss5v5e3CKIqWZGwSlp56IgmGkfEkG
phpVNlZg+gF/dNXb75DwYxCyeC9jT5dBCwTYYvjaGqpoEJZ9g/RrLLTkRh+7jVZKxEIB7EEVrVRX
ELdiP/Jb61bam9DmVIDzhPMEAy+iBOaI6jN8fN1yS+Jxel4MTokeEsKDG8vpilYC4TQfikm+3YD8
A5k/lVlL5LV9i69zbDdEaHlD1pBCPFr31k7gD6lf8Qz+VWYdk6K2kuH6XrBaDbfwWbMWn3295SRE
U21Skh03sSz1oi3Ulf4kqFM5iUO374UxH8V1KDn+/nl/P1wu/h84HR2kXUP9qMYu1MIWitgpaHTH
U0aXG82nf3YkTCc912CvIVkO/LRP6P6Kq343/EqH8fbVY2XcbB6xQVPubxCdJc4l9XELwzm3GsuZ
hsdT2qLxRNG2DgpdPLSC56mLMwtVrAoKclqGwuQQtzK53yDFyZr7Y6lO/venUtGYeKj3f/6qvZhN
Su4TBBanpL3yEv+wfkmQlsAUbrCIabHxTtC3pjytJ9Afaurwg0iueR4+aZO3eI5QNPJbUMSWcPlo
2kGHx6+eX678gygssmRCp3ku5Ztf5d/KxOogSnd688vVUAIRVMXPHxfKXBVPI8wo1k0frKektTzs
iIRQxX0b6OZ8zLZ5ibLgXJ+lBWsgiV1q0Z1pA590vVGkUxkCfdi3KR0EDKZMzuN7hsFZrnWNdvpz
RoGf+CiE34ZvI769ylrAKKcAOJ5+weYxjjWx4lRNGFho4j8JTi5makNHEaJMrNHOmKdXYYmqhKZn
0Sf2nVji54z6wH5hwF73AmVDP/stz69yMbQimqyFO3GvgFb/9BWzAhrKbzdteK3T0jKmeAvBHGqd
zdheasPLoGJnz1ydkvscLD9LXmhCvgO87UAyqK4rO6G9yylLrVXlxn5KdO3S/ybu69seWrB0b5ws
ElurETLsC78FjXAy7tgL/1hjDJHAnWZpLnuxtnu5IYzEQ/ZaY2gMYUKeuJrWeFEdE2rJTlYEIbqD
pKETvtTe4K9zsATT83os7ymi2VpaxR7tzfYcS1h6QA8gelRrzzT/Z0kveY5+ml1DrgIJ4jzNiRyn
u7FNH/GpVNxq7ZHAUcqEO/b/gsjUybtTOZHpqBzsrXVxc6V8+wL1khwOxvUACOpP0n74rVP53sLc
Z/35dvXV9FMsXGWRWRPNUCPNxg48SDttK9uxSP8NU5kxfJptEXYs6k/VtjoyuS/lqeSe2MbAOC5a
GuFIPIaJQLGrXpcf/Rn66uBIrU78ejdw4mbM0/jhcTwmcylzBHzh5ww/c5pnHAkswGfJV8Slnynx
PL/VPPZUfb2ajkAIELAnN2K+3Z1oMIFWI00odE4OeWKHToO1C+eq5cOWPSWJ30iyEUADbxzNgJYJ
my0Cr02608Mb+/JT+K9ZfoAHH4XajsZ5k0bI6L1Kd1Cez4W92gHMXpie7ciqXT+tPHar+qQMDnNL
kL5wzRk/AV71uIIzPBXj2yegekmDKLtcbQQw0LmhXYZu3FECS+Ag5ntRuyzQyotHSnFV7oX3ebO7
mN0KoUygqUSQXxCka+YLN0Y1TSx2zIVffrnySWh6caCP4iYTqqg1M3lCw0rwy7wcrQWNVTQcIyOd
aAweIBLHJtq2LYS8kskXgjPviPHpH0xdWZMQSF6JIqkv4BP/V6ZWsNLywfWaRdeMqiAz7nl1mA/G
jyA5hpBLfZLeweeLqWnWTHilktRnPzfmrVS1HP19wcb1Cfe3+M7vpSlXx1EOPBzNha0XztTEa/Te
jON3xCKYOqArKaDKhTVpITCsrn/RIQff9AEp9UFFzCdEM7FmFBI89wjplwcInJbhoPxNZevWFiza
k+KU3L7eAuu7r1PzsHNxg4a03pF40CuO+9Txir6R9zQ51YUlN+1MEAbjWK66RHZ73vnO4LLUphO3
6IOMM+jWRAxkWVPTfQ4ONt8a7E8WGK7tPc1TghgIFVMTdviV6uiTM0Hpm/AqAPzJGmcwZGwVxAYl
ivjY42igElWBOiydMMw/nwNyFmbgbe/Dk0dhMtkpmA0NxAbO/EY/Y0B27bunxBWGUG7ky6mmMN+z
xjkaIRzEJkMFKb8RcwD2qBnNCIObOLJ+5KtPo8QAyTIEYvGvxU2rJa7OMDV32ci/77wk7x4BbZBT
hBaVhZqdiQMwaz31Y4IE8Zdczk+kQczHGeGKmWmNDQkkVPOp8jIWVxv6U3cl0h5f15O5xykipWHY
Xy+MMQ3j5Fb35fiozv3RRPKrA5QQoNpg59AmdSHnfCDeZcvQxbzl+MkTVSwdEGoUVwxTRWwZCyit
M5AkzvBSaFuZSvyjmwTjTozJWslKotHoxEru8of8Mqq7fbUG2zC2v1+W7qnPXKvOglZikPz/OFlA
ObYQeGxPjDEbu++v7W3YbojYJLAplzER6HfbPP1ZeKDJcBCL2yIcUv240LbMKxz96qrfZvmZaB3s
GpHKN8PIstZ01IYi74ow4LnersfljSsbYdxdZ+E45N3JP7icB8w3LCM/deB/BNviaA2Gwi//5JeV
/nkHoA48O4YlFdRE78at+pSuHnK7oiMFtidu+QQoUNkbaaIX7+9QLK6e58TQxEcSEAbIpFz2eJcJ
C/JL1PApPE1JX+ppwxDJ2XbJTVAKvSSE3GQ1+Fvnrjuz/Ueargt4PWFc4Kx9ObxFEc2IcEBq02EY
Hkv/DdvOFTcgGA8app9w62pe47AAnj6IpKEMsZaLMzsDWcD98RFc40Zan8DQ6RC9m85B8M+RQdiz
D1KyBlDRugapVwNThzswcFLIJWdV6j/bToufljD1RX68ZBQDMmy1pwo3EHh8TZOJWGwcNjG0X2ti
ga1ujl9hemgIGZc0AI3L9zMxw8sRSBU9UT9ARcMEiq1wKlRv+p3W1DVjBKDSkNAa6WEulrpMN/ne
2WR/2xckgHqORpplPklroVAr9Y1y16kdiUcIWjxzpQr79wIGZyQKHy7bo5q/FU6igRG1rD1+o5FA
8UDTLWhOmnUW6utHYSXlK/zuUdlGb2KQKvZa95cuwG+OdEbKvnh2d8AKXoD/NdhZINUp7lYtqKa/
IZhGdeeJaTSm1b47Y12BKK9qaNIj4PBKpOs2jKRAw+ElmHuaikNQisMrccVUVau6o1DhdaE2ED1w
IpoOdljXX3olaJSKvfUPFZ5mw6L/3e1QArSNr8wCspYNO/1FVqQdQuqEuRJKCOjTprp0L+rHsqR9
qwFZdP5KLJPzHztSSjuUBrlgGN8F2qa5Od8Ba4L00QTP+MmKmPjFQMn77+1izNfv2lK+610R0DHB
RLgxRWMwtyksOVGOy+Ai16BO8qoQJCAY421MvGya2VttcK7QssPj5IUVAzHlXLw1NNzjQYMzBhCu
8+xXrZ8CfbHhGE4gq4M8vwjQp8YdA8awwqc7nTMOIsWnzmUsfsPd+1DgNzYUngxMtC+UxkiZibtz
VwjM+tG1GXm/P7sb2Yvbv+gQkSZCsEmipgz6HxKMCUcnuPT/Z+RuT2FDOrRZIV47mdOsZin7EI/F
ohKsZSG+UZKoBV465V1ROeqtp2c4ndYnKknOINcZNiG2rKEALexmL94JQOwe356NIJXa/UlNPo/P
hUs3H35ijK95YWT/c6csBD3RipsBqJg0+YTMouJ5Efn47vNKJCVo6/wFXHKxHPetxhsYXz1y/VuZ
KQI9JD0TDaxfHwh1NFvJTGf9Osl+RJqtqbnjHWDbe7b3gV5ez2CwuaeYY4B4o34EHu2w3Qvmx6DB
bRFHG3cb30irYBdBWJ9sDfnBfFI0xGAtSjWGaGoBG7uedKnnNg/mkPwFTyw2Edzyu01XrvIxfxst
2YaHEbFDPGZ13097Cmu/d/Sb1AFkkE4Ksq/5RcjN62cJYvHOp9lOndPlKcrkCq6tIR5sPHyCXbDW
vThDL3n/+VZqCGHH3lgvNNAF+qKwh0Y082newc7V1sMU5uiOdqu5n66bGA2aPhjKfzzUW7K/pRbb
Bn5rfCTVgYt9CZ1ZCBHPfrS5d3xCGC3vk4P+6y18zBmg3vyhSrNfqf5T/LbD70TMb6Agpv7lfuVV
x0SUdEf2PuVnNtC23lepjTdXf/DFcWlS10Ir3njnyXiEegLpVfIRYHlHL4dClfv0RJnRHc54k2Up
KAMKCcoe6RD15gwFnd+FZdCBq1Epmi0/L58z3/GICbKA2TsiBi8KwWEXvarnhWNOCXjQCW1w/tAh
BgVhidHa2WVZUQSf6DsZAiYIg0KFK5Jj4at5PYSl76qCnlHRpumL0hGp53xplAiE5BVte81txYU5
4mo8hA602J4asoFkeuYLtOmgr9prrAMn2YIq6iF56reW9yt1NLlyz7loVEaFzMIk3MuiysFkWnVv
REcm8JxOcSXEb45+EkH9gZz7O04AtRIX7wkERkJTqgyEy6eycAcXxTNKT6kDj3T750CxrWU2RsWY
TNph6eHD4U7rzu3s8YaZQ95/A53JhVeRHxL3eRR8I+5pDNFVVa+8LEKrM2subcvZyoAoYcChnNRN
oKtCtVOOTciVKjohZMChCar04eU3bSiICTkWxpX+GRevEafcClfzX08+L3Kxdy1OAVrEtj5e06w6
rPro0bG6Hw74D41jq4p1wk4+S0jqKbZM+TVpgS60Lt6Gp3XcW2Be138VVq2sbym+iwZGNLuIxeAZ
8mTaB5sHbQXy4eQ6I1G35nAUyu7NXY3gOGwVM1VhZUV8bmPUCkos205aIJrzWmCxKb19nuEoH1Wo
IH1c468ePcGGaPoe1leq6cOGeFSRuYee+hCFTbbiqAx/0uL830IRSYOlaFL7P9zcpNgcvUpdvDP+
1nsawrAHr9chyHgX/eV7+VruiqgYzUdtJrRozc7xuznwW2NWcWy1nUBAAUskhRyS3F499fEH8a0s
KZhujkWMBbc8d9Q9cdJ6mMj0SrhViDQpaGLpKFZRC98gSGZAVR6ZWGL3tmrKVChkjSHLBT1AS3xx
7EhEw/k1NvIabcf5cejXm8HJgQMlsyLU2IPKHBeVmpda2LSTlgwhlAqwzeUW3RMwcxjgehSHGCWN
TO2FaeckDQZyp9noBtGuXAJOVyiNWUbhz9y9242RZ90IoJF2WLNlrZoUuo9p7zxTbap6brdyWSRb
zz1TJWRAiy6YIq+/tQe9zspCpi0Ag1M5xIIGqZWgkIJm9nvlK5qlX0j4kX8YneXzI39fX/cDX2Et
L4BglSdozimX3dmtDpMb+49yZnKNYIvOmsOahOBhfmZzzcczGDalPK99sSTIfzeK7zoRU3XgRMmq
sudjFojcat65KxoTf2SgTqQE1MH6HFH+krQT7VsfV+hX9QmMaSbM7b4CXYLu+Emjn+8z6gxaeuBw
7tMCZ0wg3aA0yG8T8pLtPhYcGyoa1swjyPv2LnN+mFt0E1n0FKcG504d7eHL+tMhx35YsbxFBbvf
GbGsK1CHpPDP7SxAiQlz6Ofrclo6arC1bvKfFvOrpjWLYTAkeornSeItMPOkyeUEFjPHuSp8zd0C
BT+etxoTFYRkrn6c9GuKzQzSDsUd+8s9e3pmRCsnbC7eAjcb5kIxKcNandb7e+41tTrzzA9ELzmX
hmDqnMvePOkIJAjx03voME6d4PwFkP5DNeirIvY6oGgIwsG3cOehQU6NcLxStT+pK8Y01KWIZO7a
UPuz+hn85R1BPgSjP9UfIbY1z3V/YGVQcejxny08FYmspmoF+v1Vv9ZSJP7eJtQgPTHMnYKULwRF
sMnuLbZA/tN2TMkuoRv3BZBdXdwNa6UVD5CLnJkxn6OWF+Mm4k8RP3VnsOjiSbsNVvpSmjXCTLWp
vDNbn6aEr5Umg+mXenvIR4e6UwXvEjMy8VHiIVt9x5bNJvY4Ue+AOCHYLAX+I1SYARnH7JgfftKK
J/2xAPdHIFNfUI8g5ui21bGB1YqvdZ32nVIVaLOD0R32pg56ZVN5HW6sFrGoHJb3WewohF8sVAnj
yWFJBgOTSyVqJ+Rf2STGKUWIKX9zLVgGb9giKP/besH6UdY/TJAY8VHoAm/FEKQBYrn1Mt7t3t/q
ii+brZXpVVu0Efy0hpPkShpof25K8Ceokwd2MzYUYXy4Lfxxdft1YbuzJyvZpADtH1Ev/OB8ukRs
88ln045yUvJIkKfPqFK/+JTm2/jqmjCRzqjOxm6BNvMluWaCWMAyyr7upoEDxYPp4diBCE1o3FrM
67G4nwiCNLxsRbmdZcveUTKw4yKudkD0tmR+OR+kkX9a49A0xYdaPGpsjExiT6EHAEbtY35FK7Yt
5nYPNj2M7pUNPwsLPZmgqcEB2Z76k/DTeItZ2mVMM24oZJmtUMetc0RUz6NrKWab7AYf8AuOFonE
/3DaK/InvX0/OCrtcBh2RrxfFqwr5kGB4v+Ft+eScKdfI5e8XMngbO03gVsJxKi0s8rOJpnGJKNk
OYZbpxP4bi2k6RKjVbDde0XMyGEKsiEk6QON/MJsl1TaBxou17hPHmbbOwdpxDQ5HKNy3MjSt9/i
Y+JE9KtNDiXkzmWJgd/n6ziScg14773M/+E3e/fM/JSckRCBiOzwGqSc21TaRSATc0lbkkEid3vO
18oG2lq/DRkvncr59R8UIYFRwLEpp0Q6WOfYSavVkPQ1mePY5zVho5B2HDSJkbJmjfDGL9Yrf6Zm
W8pgvOAdZsGuv6o0zkfgqPMTHN0iADF6RKkh+PQU61h5DvJcAUr1d4zD0ch9UmP4QvU1IzN7d3W+
D7RNHamsnrShCm6s46S+kZKejBfWRlS04omE7mlBzKtZdc4Q/0nhjbVl5Ogd0kz+sQZW5nL8MFUT
D5fOUmzlZAyP8cxNjmPIh052ifsY6TMtXgvoHyD+lAq7lO05Jt1KSDKEFNHQ2puDo2MbfFLipZlp
18rpjvS374SJyXMm5sGqIvwBdVQDugB6Y8pfaIaC6VtUjIuvD2K28Kkvh9D2r+nQ2aXEOB5Iw4/4
sxIQgRf6vVFA2TzMdl7K4rVtAfZLkES+sPI1eeA+MHGLaQR3qfYSijgEG/10dthdyE8IqPLQOw3i
rNedzHIjiwqQuEj/tuw8d0uWpOcd0S5lF6W6E//p43yOirrJ1WWI/g9bAtlaQgZlCcriNToKKBHN
uS/EUdTLmM74x/UOJfxG4+f45Q72zk+xFVZbobDeb//BCEV9/NcNtS24gdFeoZ5lfYXGMQdr4l/e
o8xDyqg2Foq4MAbYdmYHiCoWzrxK+Smu7G9Y2RD6UomsiyqHu4+8NDwT8YZE76PZbZIPJFq0cOec
8+HUtHx8xkGhFsfZpSiHhxZbhFbVFqj6De8pgJTvZd6wJ8ewihv8guJhhZN/AIhlGPPhgSLLXAj+
NalGtgPEJrJH2oT/HBGcMxgNC8dqyPVpb3a9QRomP613hR0SQwUX2YbOhGBtp5fqIvCljHK45RWs
LSi1OQ8Gn5xHGfIbwzSOFdraFKtFjcTkKfP+5jb1nBw0ri/aEW39H8OayEWDcnWfC1iHwT/iI0rX
9zBEt+UFgUa2DCPQvgEVE+ZM0+g8ToN/Mem1R4Hs8i6sjWfqDfKMHkpY9VMCWKhBkJ4eeSfLpZLP
22JB9zpRX1Tl1iH4f91oSUmiBEHKM6kRWca9f9qsiBN6xicHiS4+jjto+lhBIuiZnB8oKw25tSJu
V49GG21Tpr6uYl1Mok6+GknQuK878pJaQaDJrCV31XyZ2hnJCPzUIhL5ID5Ug88BNM3CgcibOjwY
QvpHHGNd7q3VksLnzZxZY2mG3gp2aEOddbwH9EPRmDy+Jfzd6qkk+Z7RK6x8yqDfgbjprlTQECpR
HWPyBu0nOQgbkgkAZztab+DBYtcyK0+jNu40VFoZIihIJSplQOjiznKo467TyNaYi+B7Xtf6spOa
4hXRSXS25EUtFJRTEHCiRVdhyIA8908gDYiEGs6lH2alodWmuKtwXcS1P+PzhozdZnKCu1BDNc4y
7y986kaNtkRKyPAm0y+rbLNSecEdx4lL+SGN+XydTiulY7foLHVmnyJmbbYDtvkLmJCITMc8R8Yo
4pR9ZSKn+c7g9orqvwE7LmXke++jltrckPD/poRcf4GywCbpNNXs0RdrJcEFN5b1W1gGXueUwFxa
Y6h4DVYhK9a5PPmpdvEkoqdcsOs2wqlp0qtjvXfIAv/FPBn6Q9oFDmjYmoT1FxyOoFsubR6P/YUk
3W0jtvcDXckdUNKLrGNaJYeAs/4ouXtQJxoyCKfB7hVrb83SObZP+eikR+4l0zwNEc67ZHgvUnAT
C8wf0yml04i1nwwYqHo0CGIVL00DI8jOIkuZSDRtde2+nOBXsz5QRXVFJOHTRDh0FDkfTqiceiA1
UOHgEOYarboBc+1LtzmPlU2TDapIhnP93vRmSLPJlt5GC69KmonqsfUNblwEzR1H8Le2Pj6hwepk
SeBOowlcz3mVg1xRWDS/h3Bd2n1Cmn1N1IZ/jUWXbknF19HETe5y3EE/AKquXVGJARBKWx0QrbqE
cQ2cl4UI313YW8nfXtu3gawnxAEi/WBHIPNjoalBwK36eVroBqbHXjxlWGbKF/+VLWrr7Mf5vUyL
0R/vlugP2vvmWTaieyrP8vyvp7akmm6fjBwXENj2LUS5+3Bm09ybe+MXWdzwRS6iHfpOUx5eRhsL
vpY3gpkwwQG7RmIe5iWrAYx0KXOmldekXI9k8bjfNYqcoTfRXCKsFakiOGdHeMyW5SuLquVyy456
YJBNFX7TS2FsmTyziwi7KfuOVzNRjGUFYaEGYiRjKG5jairsWyZ5nT9zvt0KVLygjMm56CdLJ2Ip
aK935TEQo0AI8dXh2MonFOZkkfoPwcvceJbYJ6JOB5bHMFNYvGQBMlX1qSlYzvjA1+qTWFqXmbZh
Au+jfveXUB4umkVg2oLKND1HWGI+mEIP1libzDz9AIIZZnJG28Ez6WqSkVYXnQGC9QKuT/b1azKI
WEza1jgCtBEbrohtnC0Fn/P9VrqleiZFS1mIt9qUMV7TgMIVAxsGarVrAOzVI+MSm9QB6KfXsOvd
fArMzMYQOH2vxbUXbyXDy202XV4iHy1w4wX3kWDZ8X3I1SuczaCrUIZAenGwtE1coYfAcgQhkHmn
bci5rF1QdWgD85ROb41qJ4d+xJzH1Dcrs7462lSFxYFEsmpqzlgrvHDn8e1KoQNVlHuNJZ0UDOtB
8vcYdd7shLn1MdEVq+KPu2P25JXmV2NYiDAQ3HTsGK21zuFNMEWcFm75DFrhcgIWGScr6+L3zf/s
ZGlmUYB0nQHe2PSCjK9ZTq5cNj/TgNgb8Y2jc80al3oJLMiTv49H2IshLjyyadUROT8s2L/wSV8y
FIxoq4/5xaUwAtR3augUA7RxGvGT6PNo19HH87MH75waoJAN5glg2HPyZhMBoanxs63Fj0FtkQiy
zlrnIV0OWQ/eAIEVlZf2Ci/yQWdJ4xvtvG3ImynCqhlUTkstocmNOQ4PqIUnWKmTTCvsytiv/1+1
0SIXVIY6CSAkWhV3K6l3CY7xn7PXOuKhsD5g5137wRXstc+EyRXC2RkoYTT9mMjzXM3Uazp68c1U
B6cd1m3A84PKqkYOI57/OuuPU92OB9gtqr4cYAl1ReaVZZQKGMyyIel/AR37n0bepJtNk2yYEwl/
s1AcT3qGzZqGO8qSYeMLutiVoZM4CX6aoH993itFxddjnfMBYFCN6dn01HCGwa7fgVbLKgpIggeZ
stnN41zCbK9CneRUbo8T42CsRTmt4UDv+3koK46ZMEQArVpSNS4WyGfvse2w9A3Bm36DZ79STlaU
4WsjH+Ynq7Ld0F2I7rF5AP1ep0UBiW/3e4Qu8WCDi+jZcTGr905ixqGTHKwJUrhHS0tKDQEQCFIa
6msMOXug5YyH34hODzCyJIAkuMXQEOD5S1gG1fwSnR4cZaBpKLn8TB8sgn/181b7fAKb3KyaSPas
J31suR/xMd212dGR3WIHeMhLA7bVgIwzUfCo6K908lG3oeX9lNfPMtonz6xoW2lME4mFc+l2wUbp
eDyEopGA29AujmbE69U9QipZcGd6q7vjosPodqo9gyGFqW2wK7eEd5yAuuE8ZHkuauTHV4IbSiUT
l2Nc42RUqrjm6MGjGQkXOepFTijCu8/cbbnAQJGiYpsS7gisBINUstKVC8bUDphXaEo6JJurYG1D
Quwc5pJVOe81H2xnTgqEa1WShgSzKvOjX2x6JIcXm5D2sJzLTCfLRZLX/6rVMhMrSpvqPX8jytwY
iLoI9oLF3Rgr7qaOlpusAHxBo28uz6eE7zWmj95K56dTN0I5DtALnjl+7m+8WlQdYTddMoAYLA9J
a9Linrxq5YGCMKS8qkt7ecAZ6Jf/RgsCS8tHk1TivltPE4v0vaYaqrXhckzwHJnCCCtrlEv0wtLO
YctMlVK3ry6kBpqOJkK0FIk2TYo9FAguaNIiDqZAodje1dbUvhKJKcWh5WmPCg0rVeoDNPerg/hH
GFLgGlP9XLjfpjZssJCrCrl6jsbVQhel2cFANoaTsB+xicCdD83tcjiIgo3/w4/GuptRyxv47UER
9t9Bw9Ku6sAgaSPpGl2ybN563SnHtTpCVk3f9uPRbVsqm/oawmAY4OBPKq45FnRlHpPQDsN69+5r
UMFmgMhCUE13tldbMzOGSNhWX3rnEkV4yJoSoSWOeyjGIhGm2SMQXqhsDDlMYlkDDp1SGzywbin3
Ouuna5gwCqXELsrtk6F0sl5GYLPAWEe7b4za+huc88GdcwO4jKZkOHHZ0moav9GlVf5bosT3PE0k
xOJWVd+6AXfMUaXodPt7IVZNK0eYortnP1GC+ENEaxj8wVl5kSSMCSqi5xtPdEZRzUiL2GxHghjH
Bhs2qEmNDZZ1vvWaZ6WdR8XXGI5op5uNdUkr7No96Sbm63xJW2VsMZ1PqW9d+5gkQnYXKfj2Frla
j975y7NWFzg9BpILehObZCP08Wc4KYu7nRgleCqlxasq9pDUGuXELboGx52/fidq44iVWVxMLAgU
j9hOF6jGQnf1ldfEGzrCNXzqfcJ3ldJ6yv57GGx2lsUFa0QO3HJYXPLdkQ4zxSaHJ5mqudmiNMJu
B3yjX/NvbELtVWAmBig7tSKFcWuGUdEFlOYAAnkHhPUgjwLlV1Ro64N8AObOo8bhTkCx+lk2Wta9
7owZ2Ztl+e7uRZ5WoTA+Rzz6JYufN+x0yxq2g4XSzPuuilujzAv3++GRdPh74oYXfSoDF6DbFdI7
vmJ5DbtDEGLNYHyl+CsrawwVl7DAdLEc1t9jsjfCSHVQnA6GaFfyCqfyVuJxWOvuoUtZrGmWR7Um
fJKtyzghuSSBRH/XLiu3C8cdKqe9jjt6UgKOrbxtZ4dLLRlGdi+4lzq4OkNsDrtH4xIz7gcUvMlK
8SmLPWdCNF0lx3QuFz5a7TiKHeddK350WcCl2AODJz+cwW16YIlu8N/DrBJirc6XoDBnjJO++WLW
SMFpB2elQTuJa62gnJmMLyZ6LEBte89UxNPaoH7XfKA2tamrDUK5eSWJu24lXXR8JBGU92ompE74
H3k5ijuLYzyA+G+aJC3lsszgK5qmLBdcvFImVxSsT4N/ETol6Qm0+tPwo0fJKAMWHiq0iKkuP1Cv
AZft4K3IluDc3o+ldLWSJX9ldhZ0R5Yx9MR8r7AjiiYH5hUd0TEJIJ+Lwx/LJcAtVbOkXWbcGFlw
1og6B6IzxAIAL69gIgYMHcCHmm+sFhvz4HpuoxXJoe+65u7GK+9XqxHZkgzdrb1Wx5rvVgQ4e7CI
2241MfPyZQmpeM8GkAIja5LbJZdQiINKf4brGlrIvH6cUV+M0NsYOCXBki3FNW/vUe0Kspfg8iK4
FWhIa3SwQ8suqUWXXEtU112jXSp40ndsLkVB9cu3hgQzY/WRT/0QlWv3qPkBFsYxAmZfYIFNCjrC
hRn6ZzMTSJDRjxRUGE1rTLtWcFiuC9aLowycXeF+4DzKCf5B30JKVMul4TBjYOs2ZW5/cJdQUfO1
e8G6BUOD6ir0niHXyjj08cyf70vUy1tT1CvqdgmxRaq5GKHC5+INRV4HI1De84z2I3yT0+YtnuO0
k+dR5yl7xQAxMO5adyb/C51RXCmLrDVB+VgIk/ZsV/g6tzrffx8LQxU1LN9ZZBA9MZVmrWCJClBA
POwrhn+LRJFmlyE0AF75qg4+H0Oxe3ZbvYnbN1oCEKlr1On7jEWWdly4hUOKgVV5mKV7FyPmPOUn
DChUN44uI8ViqIsh3nzu4HcOrmlHV/+bY8ahFOjBHWVGv8+NsaT45iAf3+1GW6vXD/1huuBXZp1H
zDo4ffXQde6ENixRfEmtv9P/g5SiTnfwW98Q2ucjj+zo4Vsln7V/Ma4+U4R2VAi/Ixf9t7Dpsn+Z
yuWRdCrHCYhN7X4jPhNEM9005Uh+klnDnDxM4WztW/RSATvIUsvFmWFvy/lKAqwe+QSEWb5m1xqB
uhghgZ3K90cvsULSk76vP8bLB22NeCrvQVx035qRqGP40ohj6RasM5SyodfOeV2j937JPgIENPJ0
sasBE39cdKi9PDONHCT4r1adaPcM3uEvbnHYBXeplpG3El7/rgFWifDBs7rtxrVpHslBvFcDo6I8
HK7q2B7KMkaF/exYIjB9aaw4WIi7BST1/z3lmNRf8FOHFXlFYK9IF8DT8G/guXCyjuMUBobX6F9J
CiJY4nu9gz3b6hlJZcFLDP812IHzhHurZ+sPqZaMde91phzdXwiDLeNt2zc488VvQC9Wh+/BL3mb
0oTJNu6KPEC523Epqxa5wiz8cfMm+727oOadt073blplVqYH38Z2mjGDkQhqz4YERtqIsD6LxIQP
CSNbkpikPRXPtxbYtIv4xGVtGATvq1GgkkTXIsA/T96T2tJDHTQYXH3p5glI5p4SiGxNXeONVups
mNhvdKzX00PwR8UZUXvUFzI4d1cQFYNHyc8Xs9LaRALgQ9/+AlU1uSfHhjm+jq4/TyXuQNOuGKmB
G3s4jnN0Vz4TOV1LPnPD/7aFy6AzsmhhmOZ74pk3ekOjMQDe/MiF58iMZlGBH+SLTbonPLCxZH5z
i5qn4EnckIA2aj8/T5GSEs2SDy6kzagmK9UgVwdoBH7hrOhvx6wb9XnRPbRPExcFi4gdIVqOlh3s
7l6zXd59DzCjopeI+Gp24uBWKJokuzDMJvuT9wIXVqydTsWWx3YhzljAOtod1Lx6IovNMt8cugUi
KT+9Sj/Qb5/9ZfZSowvqn41eiM2yeMoa7p4xfbvc0Oh2kASUChLRUSKxj1MC34IGnOSujKnWRnNx
BptQbbtYpOHbPmlQuZg15pim6YJ97vDaxVILDEEiZmjDrkEXzHinvJP6ybUX1d5YyBbpPz+G7LXw
6lrzsBHwgln4jovBXl5xut50RVyaTNjMUEAyhsjE6jAjUUC5XCVBZT2qiAMjV978QAu/sI+63U90
E7WH7EnO+vHyInF//ofQoLS0BB03CY0Q0fJViLPKRBcWcPXPLPtalI9+uPCkqd0AXSpPpcoMBZlI
AvM23g/VSqO87AVwNjUMMmzqXxvl8o01U1kJ8q4Xq2bEmYBzPxY0lFuxHqxK8JOEZpxt5IHTQpzf
0zFdHcfk/GfvlA7M5pjTtEp5VDKE/T/unl8V8iqsDDmWhbcbiNibXoP6TseMHdtiESchHgoeZD1J
+q3pZvcSdVrgL0yvUgHJ//FmUeRCbxZtuYJyBQLrVirYL7vQUtmuBPBwpDfHr5pe07O1bG9AkiHx
XUDb4/K5rWbXBX7a56jEidfFHj1TSX1mJqG3v9nYeG8X9yUcCSCuA7/fi9VrL7Gpwght2RWn+U80
G5l5MmWzUWa8mvO2g+SwIXFI5tBGJiwoSvHI1gTEYAU0Kx0O4SE1pvUrVGgT+KJMq5erNZ+a5jeJ
S5LVgMhbEmMhJ4KVyCwy5FDOI5kkRiqbUv4TWqRc8cWgT2kq4xfblHszlYCrHuZgj+/jgFtJtvbc
XJ0/t6uhRLny8gfgoCduWaBKl0lwiWrB09bKBHWOn+GU+4GLX7fHPPG+t03L4zKRHQe+0qxISsy1
wmU8snXYDxuUkGW2GQnddH1+eUtaWXfxkLR0r5HbkUCit4wIOJUcZwUB4FIjBxP0xyucCLH7NFsR
MXtrPQ6BSdJrdqldboufsC1Q4DC9xWbEf/+Hx+W21ycnBi1If7I9vba0/uM0Ww/oYk/PjnBPdlgJ
lrmVA0TW/m7maFj3XOUqpD3Oq6I7XY0Fft78+LWh6j+gNk8hozMC7dyyCGRtruQaParIt8rbymiA
Jl+i7PIl+b+0Yc0LVscYNLi5NknG/5QIWSWmVq9x8/Nt+qpb66/Dvcjg/2lmH6uHHBf+CTBuJqjQ
Z9hi1xhp6KKnC0hzSfA5XoTJoelFrpOCvAtE+mHkHwuYxXANSm0Fb9c3fsx6+Qy7zT2XS7pyfSXq
dwclm8Rwm4c9VirI0QVMmPwCRDNi7zcwdNLC7iC3rVE+Jto3gWszp9M25XWZ8fhRimpVSRKEaYZn
qTxuoWCAgLR7Sew7n24eci6bYR7z/Zpvj3vy28lGHIHs+j5YlhXnG9sCb3ZtAt2YElvku8Zpsaya
K0/vTNRs2EryieQZ9paxjpnTdAVLChFFBEBMDagQjj5JoCUQc18ew/r5VaYMr1FDPV32FoQcjU+P
6R0/Cb+K6CqH1/GAKMLdh5lK2TIAhLMRD5RzzDsMpHdOcjmj3R3gzJcEz1tHmJjsdFSx5NxzMA+b
UpPjxQvGvUqpvrLG0CSLOHBddG+SrKGuHRAZlih81VBRZiA/Hoi/roJQkk4H/OVJoT/sjCE4N+mD
kfQfJo4sugR35XpAFP6iPfmLvcg2r0Qzh5/a8oKKQ99IHsIOlTl3EpRefp5ZTvQ91fKRsco+kXPl
KA9l8XATjZ3qLjj6imWbvwlzLBmHyDvBktKlVaVioAC9TCDhX5KmLN1expPb5wo7ICOUbjZXd8LB
up9oASYvyOG9f4QePVTcB8yD2n9riBzLKSd+pkNgZ30rCnIlOuqEGcrAR2U485vy3uQBw9rmBCPg
pqQb529fIN7R4M7gSX8DnEp/ueXil9e1+HwL9wPuM1ORatA4PJBdhrcjMlmInDu0t6ygpcJF1PUw
0TaXTBNOhVZr07E0ae4QOOl2WAh8X1Kb//gWT68NVYhxzpR5/vPqa2hoyLS7iCaYwaz/9D4AGjHh
/cyH8CfBWSUmTwNIiYr/8H5CHxm5fYI+j7TNoa6CI2Dw9CRkV6rfLw742MCtzAGI2PecXcp/G7my
nBeIZ4Tq+gU1MUD6x0LZ9bC2DRS1E6F5QmcnUF61ACDIToPtANY8LZIE+y/2cAxv1GipeZlSTngW
3YwhgVC7/zaoaPRm0+mXTBIut+vLMQjcqYuIxRJ+HLnc1RFDPflU7QfTTR8lgO37X2s9xLyX75hv
0wLuzfv2/SJ4UIy5R+00/RkWRy8/mm5Z0OpV3Ege0/Q87ZAC7PW9J//Ifr1R49wv5K/wL6qnksVR
m/TA7FwBaZfngDXWHGtlll3xr0kQfhwhdQ5FbfY4MXcaUR2sb4Qyu0rLE4uB4wiZ93b9Lfl6bkhQ
1r1KH4yiCaBdQ5IKyHDCK0K2YzaCl+CzE3oUQD68tZiMFtKONrPXRrwXX6hG1n3iiioiKHyS9diF
EhGyG2FwCFfGkOTqxnFHeSEa88huSVG0zzJf3aPkUNFPFjR/c/Cu7VbnyOf8IOSU2wWWFr4ueSNN
6POEioJffdkPcLQb1BlngUXa5jsgLm3QURpG1tlfW3gSmAYR7DKwd2fTI7GhzyhjV0UBCal26hlN
MKS85EB5Kufh+t8bObYyEDiOmohlwMJ61eEzPF7pH/NVIPfSq1wHJTtoTwC5e+WwfnRQNYMRTBkc
jptkh6xGVIUZiBGc0FEAAd3tVT6Gx9EHF1XtLRb4Rt3+66+M/mCuXayHp1Oj4XPafT6Eg3XoMu5B
YVaX7cfp3N4BjPM/iiAWYzV9t2tcvVIHdA2vo2fT7wPxLyccz1jLHQQmU+AHSDhjgFOirUZozu2B
KHIHJGKXUYdAi1DkTvL5f8KA/t1TOTrR09jwi9Z2a0qUnmgZn64S5iSlpZyKQBTLoc8MxFT8iElT
jC9gmhHsgLbaEHlBUAxTimf8suISUuIpksk8z5Y0UfXAW30/d812QdTp/rt2dOqxO2ESL4Sz73Pw
UA00KODl+p3ECeWIDkO22epzKK06MEVoNDwWhmojzL9V68JnGOaSPNhVhPyX5hmxdCqdZXuQk+fy
5+iXCGX23DHtQPig0MR3aEgwX4jgyEbaVT6np2XcoTuLisojHPrHk6DjdY/JsOnqq3TKrD6iXVsH
t2DPvucLRfPCUQpusUhAH1l6rmGbdutoq0D3PR35z2DFdRa7fE5SNao4yJ5+DyLB8U9JFwClDidw
8HorJBQiix3KwC7VmIMC7//VNdtXZAy9B27eFSsJTgeyNIKEIOpvZVaGCCBGxcJoNxkDJ94JauXb
tMs8/MfbuNhnBCINbaYhVpbowA+hVsOWD0GtJGgbOgiaJO+KicRu1c/JdNPi20kUOMIHdb8zSYzD
PWkRjApoSAB6BGWvMKvHxKdl6RS9llvhRS5htfE2pl54B/QtjSjcRYKUErJW7IWiZ1pUyr7k2/NK
ugeIURP5nDOj6yV00bvGAi9FYpqg5/smXUubNjRRh0iiDP8jaqfeSZbVQV9ZWDEwx/BnbDXXtJQV
gFB0V3TvKkBcRHW09yTzhtF+XAsmVSZ2yBastnMtov2H6ZaXAJIZeM/pFqm0PHN/OUxD8oiCZL8M
EmkGZ81JU41XO4mUNOtgeoaKG0gPb6dizK7rtGhVNptb2zTaxES2JGYsei6yjkRFyG0yGYDyeJ3g
8xmMldXw+ymBJR1PNQeCZDDcgU/oHkRkJ0EIxWkf+zd1EPjTbu8yXBUIvXYWwnXt+uBiDhepUvNU
WQiI4aNlI7frqB10P2GtizB0v6Lwn9E36CmI4wPQWloXZP0zIx9q6gpS8xHjkQHDCTOOz4FK1xVd
IF1yBnUl4nYoq/p0HnY9w6vrkOCiM3SC7CzJfJuV5DZM/69F77olVowRMJFiaSEOXfhiMylGTXtT
s9Y0u5Vjzc8vQLyOuyMAEWUpXRfFJucE8KP+pTAd0iO1sLcsiIPuggu2+n4nVbBdQsMk8c+jAmTj
9AZYx8O37S6oHn4b79Dny7hsbKq3Pm4b68oL27JCseeropJ0Cp0Br9OnadRkrjkv7mIEvApUa5H5
my/k+QY413IkZzcvTjhKKB1jq5CuUY8BAuDDOImsKLfopik46TbvxMFYTpgeGqKWmlBHzjFkCfIQ
xpMYGI6qL7VYbAhnnmnAstA1WYp5DJPTU3rN6dfubPxaNm35B9uU8pkNsL9kebuttanxr6iucOnC
viG2G65VNGRXY0hnomrCPqKcLiv7ULvOBT4f+JxPr0bdcMOYWINKCbBuWc5lGLlaNzQs1LTxECEZ
e+ysFWFbnRhFKmKjJ4EEopGMiwRw2rhEMRz5v9XlRmg0QsGpTt3dqrQkwAFw7i7SKWOjPdHNcaXn
nPFN7MzeNMaWn0l47lIb+MTYON93KiFMYPC+XEOjcDSNIBiCNMn+wTjibUANUfJTLpTceuzyv0Rq
YhfO4/d8gFNn2p3dmBt+i9rjtTWvOCEA/rlmBwR0KkJmD1uNKhk32Y18NmT5DX7RLG6BIDBdgxLG
zaXXFvipNIhD3fJij+iL74Oljutp+4THGSPCHiLa0ey9xZJk3SKhHDw0BGTH3Mkj65e3tRd/jcdv
44Zd72yLpX9DTeqRvPQrYt1x/txpT/8i9ComZEjhF4CJNTzKAN79VGJ6R/45yOg8lCNwpdcUwmSt
9mONUO9edk1XZiXcagovc55pLeY8SDe2B1zSqg1DduEl/lE9JaEKdirkl1IyXttucuVTASaV5XHD
Q1wjGuagMMiBYJXexph8jhCeAVNn2MhhHth9hxuOsBvveTMLE0hX+W8oPH1Y7t0TDixNwGMhttAy
ncb9DCqFyUy3DuGeytA8gUhHJDF8hQEu5QqPF5U7Pwqg5BHStzVlaiXasQLk8f/u0fKLIC6+gsZP
2dH7M4RBJQ/VQfW9yxHXTTEpNPNvS2QKhKnhpBCVDZRl5w8bnqTUJdGYQ0ljgSx8+f3nT1looLzP
ddNeag2pTiSMYNT3yqoX9Wh4aDS57I4btrtfGEDIdi7T+/5SrfLa/payyOHnp6jHdmYCxk04Dqht
Yiz3PIEpGoXsdP8Rcczf2bIq1JzLkAX3xJjvjy+kxJ9j8GoDS4kBEWE/f/sdgsr4tC/V/0I7xCiV
+iHw1udLYKM7SbLenw+zhRTa2OJpU3S6VwG7gbg/W1Lt5auglX9vaSKzcLxb0ceHTBZzDTW1IKpA
MIyBMQXSebSL8WY9T8yiu1OxJI6MM2/4ebkRzcSG+F2E05Hl4KHWcdkCheUU2JIr4m21SNbWBsuz
kv61ucF+CJOsDZ2Qx9A5rXKVjJ3LOVeamAPMMBWirdMPM+JC0TS5p3E2azUo41i1mcnzvl7mridA
Hz+rtDWagmqqqDiF/qKsm+gNwYwTg5AZkwOJWdmHrbNJ7WSolTW6uDFqteO0phVowdKPR9rkMxoL
pwSCG8LrYxpeiGxUz5r7BTYX79MXZSRJk4L0jl8kLb5wwAdbdwn7vsCOnn+7cdCQ/B0MYPTIRUQc
f93dB3p2b72Py9bp2ApY/fKX/jL5rvceMCGV1CGj7NLFYeE0ZtA+isna+lUPWSFhv4WwB0M8LbCZ
F+6jwcu93H7LvyKSpT0tLKN31AG74lyPiBA2G1+6NNR/DNteIbCQ34vpaqgEqnSpMQpouXU38nre
5imZOExH+/hadW2/oN8A7dyPgojUTluUxjM5m8wwHAjuqidQ/ANb3CG6HtKjsKE/fUIKIw+eXNNZ
e2CTARjv5tY6u/S7f9L+D5oU3pZaV8BywEA/lPqVV6yl8n8ePG4dIIJa6hZ5YIr0pTE7e+tzLDEn
E960jehPs03aNf8k5LAP906/PxWw4If4OFPixi6AX2RjGjMIkJCwkC1/D8M6fKi0Ewyrd4e+bpU2
k6snyW+0zmZFTyFb2H12O3sc9Z5pOxln1l2IswcXUwjAnWS7HjUtIAUHr+21AaFn78w+/rOBCkvn
fUr9Wk/pQwasNbiHUw+mrK0Jcr+xXZQAjnXAqyFAg0/4h3J7YMZ8DbmfcZzYBE6n/lVYDd6ONjlk
UqMhQo8KLbWvnUYD0YSEhIjXgXyIF1AO7y+/OvPHBzNVhRyvP1soePIM6Ez5RYbalVv7XmmCT4Pt
eikxWNhkuuVT36/eC+PeB7SHALFM7yD8+nix8oRIODKNFu0zPGwv52uEh6ZaVowb/Y/4ib6cAzA7
BObDEeW8qp7mEioWSIPDW/M1CRAtwladuURaMHXhMB3S9tV/AzzrEHZAuCbQTghzzsQz9fBHMPIw
anCb5hhb8KNkZjNVW7Q0SiEhvrSr2B6Ml7WG3jiufD3VYlOrfMr18dm5Jg/QwtEiF0GoZFFm79b/
NxwMULPljQSfreLHuTQsowFK92RoLd24kROEqlmEMe1D1oPDenbLbIy8WeSlJ3eqaj8hyYtTdKSC
t7V+NUYS80n7P5mCCsBeUO1R4d8in3Lwzhk4uzcF1HJbQayQp9lhJAikmWdeHt0VPVtsTLKZj3mO
qSpVo84pgsMkRrVifu1sgjjNcdb5wSkkSr5HvTf/xW+xHldpVGewLzM3mu6m5khrgAuzTw2xEXWl
95RoVzLgG4TYZtR+sD3cIk7qoa2/arSiKyyYc7iK0n0dBfZiDFKq6AT1bFy7OFkjbuxNlRzkaaTn
PhJ4mNhOk65C9ubEn5peaF7cCTgIJOEaaU5nvvZh68RJjhjHdZyVBuPu1Wy6tL8YHqO8k2PWzkCF
pXy7AYFx6xoR7aJi0hA5DwyvRl8U7La8ehBVsQDdstG63LLOKYEXWLU5R8gr2UVbO5fT0cPQtTbr
0Bqj23yHQSdkoPmS9ZZQRwId36JHHxsXkhs/fm/ea+CzwzK0y0mP2t9FuyjHbBMTSFRg910u6JF6
5/t84HqHRIp/g3r2O3ClvMwMgCWEkcAl8SK4UFWuaruYunTyZ9WMB45XtoSgCWF+0Z+TBnDtLuGZ
R5JE+MAKGxg3LR9b1g1sA4+619UwUbnJfvFopvVHXoR/mpkp/fWU8bWilSJUgNXse4vj7OAKG3dl
rlRwHqkbQpVICUJDV1zKPM0uGtTWGVnnRbfaGb0UdEbx2nNfxRGvuG98AIuWnQobEmNROxPZk1y4
YMJqe/yym1KJEM4uQ/ItNxEanzKBfaZOZvz0GjJVp0Tv+peWJC+DNeDK032CYi2Q1n5ZLsJZy7u8
0PL9SBOym33fbriKHvPw8RkWKzTBBg4Bv47IskswTRHLQ0rgJTgHkQXl9GyvXYx8W422dx+Ejnv+
ikKYOjQ8fERpB+lfYISYoz0TArfIq6TXBHShuy+jEspUF3OCtTXsarRZuxYdPbouEH7brV1hHc+u
GFqZbetO515FqPz1bPIhU7mMT7POMw9DawA5aR2W4VWOq6XKpOUd2qpETjCa4X09cPhRGYI7ciKp
omMFX/j/xYqE/0I68rutSCyni/vi2dWrORWHmziAQsvGIB608TR0z2L9R8/ipLd3KRE12ZWEwNYm
kKQJBpweyot+GQm+UApg+9FWVdE8Td2g1optbD4IP/L/30oHVAeN2rkh4IyMGNHRyJEuuodhYJRm
ePnXvCyQZg1f/o2ily7F2MxjA11k5StBhYaKXX0Q5a/WX+59fBUg78DDX9Vndb664icP+V9+NDyn
T1AmCRTOV3LDgJF51bDkEEn5OH4KNIIDrALJUdSfZEYwkKSeqRza2yFPGhfn+/F9i29YB/tDF0Yv
D2jq+euCx1VoXpOAgW0Bh/NkEryqS3yD8quAOtbSAiaZBvboq+xLvHx36nmcP62thO9EZamhfIJw
TgzFt6GwIq5qoSY2bRV6swCCEqdj1efMm6NEig3Jj2MK7Fmmab2wJJPPuiL6W7y+0NM8AKnTHO48
2zwSaT/py+n4emI17dR449JxLtoyBDDJ+YmwSq0zNVWH4Y/va/Z8WFSlCjfu5NCT67dP04pwfvJ0
GD+lyNS/2nh75OFwIVIhXuqJkQf+OlI7CEqX2Qd0BoJXMybPzPx/0ZwYpoFGj6wLG0Iz/qGVvSQW
yA9FmFY4LznzTh7EDedGSgpQq87XAV7fsMXK9xD+AXNySifBC9FHE/RrqTNIEjqE86qf6QGaVgFC
wz1YzuX0c+yB0eK/q+J13KcxL/iSPhmN03kKnkpYUhqKrE+UDJ8G6a8XJgb7CziwbANBvPQ2Noxg
iTrPUdXHXuvIF7bEi8SxYY2lo4eVNZ7TvicbHSdzK9Kx57V0F/E/yXE3oKeql9S9Cb1yaMQfpb6M
WsJo+A2G0Qm7AB4+RwkzVwKknH/YMRgcoC7alDQL2J5o0TAm0/LlAk+IHcxfse2uriP9qdO7ZA9G
mXdAwgp6XmqIDPfJtiklmPkEY4Gyct8AOm8CGVP8vyWhKS5uBqNAQiEv+bbLsSVAqYXObrTe9mue
VCK+JI6oCZroLFj3KmKSgtPEBBiO7Vki3aA+8OTmx0e+X0PowdAsr9jnficFh8QeCqQB391twjsb
08U7aQxkzw7uc0+jW/UKRa9ns1QTjM2g84g74NLfbamhex/AuUl3SehOdcQpwTtzKGsLtD5cVr2W
u5T3zIi9tzrYMF59ial4FWiML1X/y33y1qeNFK1Z59066OWpWpScwVC0iDJnDneRnTIR1ZC3m/8m
TwfQhz6J0nS1nbvrFtefJ6vwZVMBGPeyOGodbp+I6mJvmksT2JERruNc/ie7lhrwglof4H5Ek28c
jNp4M43hUsAFxGWGtezPNW8N8aoXmOjmD3dOxKV5/1pdgxNlWAn/eGMaEXZmGcRXGpWpY90E/Gf3
R1f/f5d909GwGO6Qq6O/KTPXaKq14yJOaVUAxunPMxEqO1l9dHlzZSA3rn7nHGgZAhBJqTHN6BYC
Goaz64QgGFadnTCBNLlIp3dTdM5jsLm5AZUSMUiwRwxTjBaf4s0j3kL32wZgTpeZqg+0d/mgOu0C
Q13dt8Dvo0qCG6hma32KQ15IfSqCMqLSgSukyBYKFpEkCM5tCvYQYu+0Db+VfIDylJHtXLgIr+qJ
C25z7g0wOQC7GkFFk8WRXNiyn1SI8XhHouYsUD8dGqU87TErK+oyUOHebLIsCQrqeV9+PtsYI/Lt
pUPuvX21iQ5ASGGtAgDDeFC3QgTWi0MWfRuTVliEVFnzYA9ZQz/QRGrJFzeMh69ANb3xYA0QsyU1
bmO+zu2VChZFRBCfrv4MgS+6IMZEvshkx0KnRZf8EIuCD71AUIwiP+dPGSWqoxOz7ZtjqN/HLT0G
NdR8wSnRxj/9zv8II19Rl+OCX/K8EXOIxIZcLiPz4M1KIOb1nTJcd7bFfku6ozD5cOIh1Yf5qAHZ
4XNu1y+z2P4hqG1evvn5TuWg2nwmy4wfagVa0TW6L40CHDYHy4texUsh6WItI02Gz2Oob9oI+xky
bHQRDMk0+0AhiOm9KIfmFgLHYVPLP2XcaIz4xCMz+J0fDyqFzjsxe9Gk1LRrYelKYRFNxNG/DM5Q
CZDCu1yvKlmzjrNhD4LdUcQWenbjFq/btXpFf8huNebW03FQ1U8e3YYlJbu8ZI7uCBzRj2LvQ+U0
IGS0X1gwtVd2g42wcav4u/71odQRtLNGiH2pkVwvEoJwkp8BHfDoD6wTYZcp0OoJckDrc9smFPJ/
tT617paaBQ1E6Zigz3ijLSNDqR6tDOlTfo42A5/GrbVLExpyD+r3lNVMaEGwL9f0tdZxiFrFc3fd
wbJ/Xoivu4iwlez6ouJTjdnS97GLMeXNj7AtHhBLr3B12Mc4uE7FKkMOXqQ+4dtJx8XFxWz3U2GA
RahqpA/L5HEE4PUbCzPzSNSrzNZBBzX9u7jD1xDRQKNOlz81U/c2HMLzAbzfChf6uNJIUhsXXJ7w
PVmKNNn9elTEItw+rAeMPzgGu7G48Rrz4qqz5+f/SMBJnxcGy3Psa8CucqzAv9Qqs9W7SXPLb6SS
IX7wfM+qGE8qNW6n/AUsJt3IcwAlw5tkknFU0E2oKdKEbpoZATMEhwLxJRPWGcMBMQC/lJnrIB6x
kaQXOPgrGOfNTF/KCAeBEJrtzSNRD02Bp3xs4ks6EvEIESt8B8fYohrjLDHeisRH9vtSwU28w5BL
vH3cAAwkMjrVa/pDQgOUVunjsfsD+P/UnHM9eSZ5j6cAr0LcAFmL/kC5Y0a4NuEvLyIjRM+HlPtu
WDx7H8Qdz9k7ThxXFsWZlvH70NznsWuGJAHXC2ztk/cwbg4H9hek95aiQg0p1sr5l+vsFwHQIl0/
bmePhZBNLnMBL6Qk5eO5pdCzC6ED08NpZifCXRVoJrRUyQnMkvtz0+8fIMKv5WUtF8F8MOq22vKM
3QoEsQMt98ZyNQ7qRZGyUXxjdtZ1gxQKHGXDreeYau8+zUHZ1RspGVF1IfTT/SgPBCH/3J1QWyLU
bxMzf1x2KhT7O6AhaDR1/YEPOkQGOOUu5cgsmDy1or2K2CWGkzTZXMv7fqYFpPg1u/PY64+v7B8N
c7Iw2+1zbq8HxteyhWlJM40oJbilsE0tLpYOgBsb0ITwUtGGveZ2YqAlf39S89TpeBgvA8pwetSN
0oPXMdvPJkLLFnqV7Njqyi6Cp4WZyR+MhgrHjnBo3kb2/IVHYmIPYj8Dds8OdRDbCwjghESKFxjC
yKH7EoLb0qA4E9ATTR7egZH0UQgKft5ckIVaw3MbWaT9sa8SSavPTsVY0KM622nM+UHsUDwBBUAG
6g8uZS3kxfq7dagsRY9HhYiVAlcNA0NQu+iaAif8fcgGgGnCgI8nYsYWDtb5QOneC7XZcuCVC7S8
B+sCjHsPkJfZdTUPbDDkkYWMDDR+r1i/xhRdIkH6l9zW4yjjCKj5eYvgni2TZIX1UHWBJZbZd+o2
TxIiSmItksK6Vsqf7FWQONuBM5dvSHEa0+BvJk2biz7MqVeuJWOeErlHVe7o793e17QBrjAsUZ0E
rflUhV/gQDyTSPsex0ztiP9wUOO+KSB5UuKpz9evSX0t75VkflLKW8AEs/spy5QcURdnNH+OwoZH
k3FUe3z9QrVWb0aAoww2WORVGSeLbHn5kMhnnwHMwJDzng/YOM6E/HJNGRwO6bwr9xHv/tlx6Hsg
DdYQ6hssHliqpc8gYOtzFs4ShUEfL8nUjio/FBCfRnT1PaN42HalOso0SkNj0omcN4klT5gqgrUM
+4MMD4y3jBRVHsQtfoDFHH3k3/2yBB8y4QGUrwRENaltUQGuqEayqBn47w/geMOF2NuxR+GviZvh
p6H5qrUe5gqg5zxjnbkn7e6dEfQwewqY30QNI2oCmwDleYQ7QkPct8tNLj4+u+1HE6DwnPBDwWmN
sKq3eKNeWIyhfz8PmbBEq2yWo3wdawg4w6+2xSlGendpjfop59fJrzufHAsp3XwNAcNxVxw13dfu
zBO6VWb5bGq2OETIowze8ArEvxrdUgSdWFfQRLphxGt0k0kktCDLXHvx4Zp0My8GFYmW67t0zZBW
B54AWiUz+NBVnpeN69grdP0Ol5R7j6OLZvGsEAlxutaINfi/073ScbtHJ4DV3djLsPWYFnUWiKDt
VQmRKTuB0ae83uyw/uK3GHARqtPci1mPof8vWmq+4hIobRcPMaAm4tnrC/NyurIVSVEUU/w7K7+o
isnLWXt7DmOeIzg8NnVjq4YuH+IoOseacz04uigzU4X5ZHxC4NaKJT0J3mQUDBfiosw8jQXBtk9S
/+sNW9X1mjujeyTPFxSnAqdxbddrZKjx1EEfkvy4zGOP+SVevO+orgOJ/5/rcA9q8PXjxnZ1UJF/
+tzuC5k6s4fT8GnuM9bk4WyeaJlvVcgwjtTR4Nf+cJoernimldUfmdkgzDYNK6a1YoOXN/H3fPXy
v1timfZgVG57Tebq6Gg43eRNz2Ec0ofOw5572YgiTlNOZxlCSfusLsH2wk6eTQooxoMmdvyBA2QL
GnkiGMHCYqlDfrQUFpSDfE3T9a4THL5DRA23VO0uWiGZ85pZr9ex9YPv0FSMDlsmkgNCDx3ZnUFq
nRMV5YfxVGqFVBHp59FgpDBCn+D4m4bgYoHEyZ6PWGedPDQN/2gTZF6PRw8RDqOWXWuNe3byo0CA
pVg/u6xtsOB9YT0D9BYUkxDs/T/sskTAZAPLD511o9YovwqP7jLIQpsr65r06NgSrF7pRLQ8t0bs
3IbwAQmcCI7AT5Nr7Y7KIzlFU4BPJGMnsmQry3SZ4VCnSfoiaeM9kK8qelFFG6HtCxKr1POIoccP
aUj+tFB98/peBy8Qpzz45ntXVS/DSPRiHdzzlaeV95SlF/HV+pp03Kus7A7QOhyDjL4oqBuEVER0
8/OcXShto2ECTou3JN0SXfdDa4n2b+jeUD6f74weTigxqlctA50hcK2rxoumfeK2dmiVgE7Qr3kS
k/2b6L/IsYoss+jyU72ZarWnlDp4LfxCfcn6TnhblRZJTf96iE5dJqvWwbKYpmhnN6uETBjAQxln
x9c/611ntVGo9QZTufvO8yKV4z9flKT+JWdrf07x79LwQPOtHwq4Fq4jC5mVv7G0enYW8W9oVUlo
tzsc1ljqAlIoz8sDBEGot0IgYq/AvD57HVS6W7zxYv+JHDu5sSmA35f8Bol/L+kb6PofJ3TRODoY
01HUUXwPpspQqw2CVZV0OBmlR0de3aZAnmx25CtcOL/q3pOS6+5F/ftaLe+U3IG07+/3eUfyd2qm
2mvshsPn1csMFH3FfustoSOH82xf7Qv4JQxYOfUNdk9X0/YSYTgTb2CaWKV3OyYVAGoJqgGwmFM1
w73gY2Cy6SDO7SWZER09Hl2sxqYTL6nBxe/EhyY+75+pVGzWgk4OLUo/7WOu6eVVskp81bLBsTXH
ChWB8JVHqrO+PHmTC4u1pQsjAPjnMHAv7uPu7Ha6iafZNh132crjkx2vpHFtoQsjX0KGO2Zi8NIy
gLm+fObv5JmCK75J/qYIwMROfVCX9XxJFfZKpBR8IGTQ2ObtZHp57ZSYFPzdcEX5y59tHRTECsnG
bRouZYUSRlBoEmpR75dXoDy3DTJqyrPiH4LZPT47lbARODoPfOcN4sxJTh342YwBpjNI+OODo2pd
L/4UH8OB17yyl+XMeurWOh1kwk5P8HUxAlQwZUFlEL9pGUCw/A2Jsxmcr/MH796Y6skaXP89Hjca
qX6Qp5CwLb550qNoWiWeTbhlozMZjxbYYkI5x1Vb4saLmLwTLb3YLrr2VpN7zgXlF6PxfRvtf1Ye
kzASJWwSMbrBZ/OMwhNa4id/iSRHrj3PUpn3hwvERffn7i6btceD/OAQtqNgACdp2hlZ4THcMK+V
2hiUZmP/W1T3JCUPO/CYWGv7lmuPxpY609AWoIz7FOAndEsq8gJZXsy+i+7lYq+aK0IfiTdsLCS1
mD1/HMKbuZXsTiPTlSKYb2oB3aUUx6vtNFQDjuHzpSxxCU4RB4EAVLWT3tc857HruHnZv83ucQCh
FHz/O6dkhWIgCZV3mdMFMLkzC3gu9hF60jbbEuGjKxe0dSdyzfAhYTNdyNkuY4YOUVP3pe6fizIj
wG0tjgmY3bHKmm2EMfCAdjTv7423rGmKv6g4jKSbC07CBCVXTzeEaiAyP5FLmdQ9/rlU4nYVO3/K
kZg3QlJ0eSyE3QAz7dJocbmhMUAtA8bjgsCeg9vUDG6m32WGSZETTS9YZrxboT5k/+MpPrY3bQaz
sjzsgswcka0fMf4poEW4D+XiA5oTfY7TJ4P6v669vafCHnP4dp9V3G/Uac8L8lud6IJoQfKAZlTa
A4N0V+XfzlMK2ik5TbkjsUXN2pnKyA1uhJDHLN0KRMPyc8+rTflZ2mSB0F1bP7fFU3W7awdW2mEc
uCYqaLnlurrwOG7LtTKpT77nklvl3RlV5EFXcm5n7nV6tCfRMpe9YW0w3W/MRThWaVIW+IpbJFLt
+dI8GE1TtN8JCmVcYwcc35jc8ZxPKXrfHrlQkT0v8NWLPy09MqOSOTQgtUOBshpyzOEprXg1REhK
nNmMQuiwIj7WVyZV06JfnREYwsjRjps4IQkYp+x6jSf6t2RBDE/UmtNI+RLWiUdWABmPxELPr9Qt
nGaSmEf1uhU+rIMt3jAGsF96Ui9AxyPyVAnXbkl4L3jggewjBFCuGYNAqrqMqQqYX7hBnop1uN8k
CnBm0XH91WnqVWGVvskaf/JYQgHV6NJevYjbiZyz3XFXLrunblnKoupEd3isD0jaS7kupYi+Quaz
gaTk9MnlVJKvkAu+KHnL68TgG26VOxwM1k1x4HmbrieBpbmaVBkSeMHOta0nYig3089PbtrrhC3/
GWrO1/Gqhb+C5cOAXOUNMjnRpvMxuldeHxfY2auS/5Uz2eNP5oIhiad4WHK4vGOMsV59TXQ7FBrn
OE2M451ZyvlpB+PJCwDZuWw9VyLUlrMcj72YWEvRTBB5+tTNFkditFpyMmhFUI3kmgaAmfxB6OnY
S4cuCgr+LVbfggJ3YgDIDmOjfwCQlENYvNUrXcuRraJ3BoV3sncEOBr4BpFk0U9fGcC+pgrP75Ig
6wayCY+6Pjqqocq2rf4fNIKTzzR7AJmxKnqq41wcqDyTpaG5RgL3nH2cVPITDeh2wWkzI97N+9Qn
FiIS8Fl20gW5xyYHForLrPnEX4qf9OfhkHcD03kuTI8YzJS8VH154lKLoSdGP+6tMDsBRls3Q/cK
IysHRUgY/TPIJCeQ7r+4Fbw31h5dJXyTpjp88ZSd1728Ou68fK8Bh1y6klqWBlxG5Sw7tC+QHMiY
AlQM5gFV39/KBNS64qPHjvzS5ImhFfBtWOHml37foHzsQG9ucC8hRD2C/lT+U6J0Zhl5s1b7zYhx
YQIMHfZsiaXWEr9485x2Rd8L1I2gn6O0Eanv2zZVVdJnixJm+x9L/tXlOjF3b75QvA8jcZMszu1T
IoaFe7wuXi6AwuG5mk9NEWyJ1P7gOsUasSvxyZNOP1g153oRoy563Mt0WPwdQNftfBjSYDEG4iPk
//DzlWr/3PyGuXzSbSA1IIR2SDl453UtH/Ibo0SNdLB1FwNJ6WEP17XInnIEq5plbzIDsc1huaHE
9A7MqaRGO9SoFOajoL9j4g8AVq1qNvtYS3NNtJoJu+KlwN7QcFKNxwxcGORgg4Gp+HlO/iPIfZai
UGFPv88x6wqMT/A06qloDTWmccF7WfHqQy2bEcS4L94l1WiT9Va5KKiGCaBaVQAQkdXBDeR7f1Mf
YFtULC7MBM2/WLnARh3ImDUS26AxoQ1ZOSzlUuBfnNVRmA3P1fgP2SpItRpOqtO9n2zha76rreu3
ia9+Mnyau0GguLo+DgKP73CoNFB0fe4HfFCGCDV7L/qo0aXT2UbeaSk8DDOG6Rq21CF/HqswUF6R
d2qgkGcCSd2VFdfd729nXa0H9ariCZbbyISUPK1HGPUOdP2Rv+AJmDqVdZeFiQglZ42loppqjtNu
6RH1ZVPPfv13H1KhI4ngOfJ7gBMZNZ7GgI/dDVP8a26JgKlRejEE/fia836rWb1V2HFfsyMA1GyE
zB8gw/vXbP0wmP87E8aPW/OthiOgJdJ2gZp4hzV1TWHrKdaUN0u+5NfawK/yx6sGy+6fphv7tH7j
5K/AOOiYylY+BzX0SONbPyqZmROkrTffFphriSwp2xMKO3clMa/DpJbp6MtfS2033hqooRztSqxL
AcjDNNQ519iWGsrO/rqD8Y+gmDeBHSOVroN7RG8tKFUufT4+fRV2lHQ9JLpqzaFjw1J+Pe7nWoQw
erQxqB1o2f+kDFflLSW4AKCk8qslhb5Eh3ZEQNbWrsFsjA9VAsIIG159EFP7p3wbZf2/+maaxf9q
/TjvzS5RDbi/1uBU19eKXPjXv7ahg17b5Gw4pwncy9ZAjAZbPCTuNrM7Mvh3M7zC/niCV/I1YxRQ
SgnrBsi9Eu3Sc2pCDzeRwqEsdvA0q1eWnZ6ECP0ZiWl5QZDljZp7cj64n9ZzLiUqr/Uj8mhM74nY
OLOjkkl65euDhUVy2zEekIfxWN9pr75KnXRw382Bi4JK7a1MlzZN4F+fLTojwnuf6PCBuqHI/e1R
WdR10xnrWiXyawtPnY/s/YzZPEXeGuWGpGKTV5RNI6S020kOPInZdtNWnuu5OMHkkozzA7DOm70+
OVUDH0owB8BXfb77nugFPJ7HbW509uXya7GiMhVBLA8QOD6Lnr6+k70xeIVTx9oHzXN65ErP+hGv
iOgciheMhI1XjulEUskRUz1JefLCQ7eibHc2NFOCd/t9qhSDCl9CFgB9tajrTey+mrEnxaxe3FoQ
E6FOsOQOR+QcEA1Xolg7FYIfDOsrjJu9bPzCiZMjm4w4bILY6m7iFa/5FmmLJmyRtrSqllg0TwqQ
QoRNOqVdSW+8njDIKJKKpyuiOCRGvTMm/za0vMXOuMsDVhL9Q4MpgleDJ5Dsqc1UzkwAvcZnzekC
jMAnymi/iHjUoODJjtkfFF+paLyriGkcWuheuWirz6OsfdYIarn+jgebkDa9cms0+UWT8MsWkTaJ
6Twf2qE31WlCHKhnvoK3haP/GiB2gNTohRC5jBxidARmI0MoJHc7schgrpgc5cwq5OYoIINpBQsx
e7F2Ow7YxjCH2huCBYLS32CGHYSsdKAtC1zYXp3vOTHO3BlPcsPrzLkevur1pL2mNQJgZ/H+9oF5
rTaEGll2bsBj8EXOmxUM5o+HPkEJ4ii3vebbrVJ+yDoOdqdmTwJ1QR0Y7VeIFz43bQsBmjoZyCMP
Btn2FRXk1x9kUJqHDTMji/9kWVLP+jMoS27afiu51WNof+rnvxQYIcTwYt6RqWeGjrRHWhz5Ecq6
D0IvPHoHmUNekYjxnpb1XVFyCr3MCX1HFM3KCEyi5Wt1o2KKmdBXIal6l9eA+2wZKLgLi7O+g6UN
D/YtqzhV42M/CRVYMP4o4yNivFnzCCPH9EMm2x2BzSOuUQXh6MPsVR0BU5AhI3zVzvleR/YugdL+
uN2zw1L1+zu7U2KJUIx2ZIdeDz5EY2EWymSXMAQ0r3mgksfx+g7jNw2AIjugB4Ttx+7O8rvkbIUM
0/Myi6xKiErIqRM4Ur0RA9bvEGHrWnpf9xW354BY64m8H8u54mTNHxA152psV8j1HWK4P8MxJXvF
1EGt813feBadbgjJOqV+nrlMdQkqDivu04TiBpT346e1ZnuHoeYyUFjS19E2Kmcg/4sL8Yz9f6yL
0+IGqaXZIQ16UFxN/e+c4n4Z2fKCgpVjEEonVEEXbI8U8sx2ON4OzcY8C2lh0Dx+r5xC3QfKtqne
cPRpEK+J8faQzyE43goT9SA3iNShTquLdJXFyKDplyklPapsL237Y8ZNGYDEDsRQDT7bTeIFrE82
mtxtmzPOcoxRCXIAbkJnAbjkqm0UY5FcOOZnBxTYIyaKcKDLuKS+pnYCRABP5e9nC97uBC92PSjB
IB3xfSUiebDdypzph9MiOukvGSUMnTQL3enhBbbkIEOXTzfYRpzgeeDPYwXHrikNIUa0oP6L+ZFw
dimUSL1yomMpbzKTTaGBbdKb2tglGWyXmeboXVOTGGyLytW+NQUShlvRHkCvbSqX3RNIu++1KUxX
7eGfW0L3AZiOSoUNG7kr4R3kbVV9LokUqExsgYwyKy0nqjP/STsWwGhWbo1lzkWqSnfFS69x+hr4
45YJsXITfgf7nNtTqU0IkYfvnfmt74MATHP+udmm21NVsUiAqSTfGT1sbo1H5fMBnPdJbWmBHdlk
l9Luj0EWkOet3OXw3LXqHS27S+J1s//7rj1rPDjIL8JKfj1NXodjZvZ2mGbxsxk05DTdieTWmJYQ
xnY4i52MgzpIwkUfxjHlf+jhOXDDg27wrNPyMP9+fUpbXfJLcbVRZkDboVK1cLsXELAVZnpEkhqB
pkyqeOc0GUoyIIf+xU/UTxGCHcK7fjh7/RTEH+ffPMF3qXAR+dCO35FzASMt21mVmYFq2JYS3ea1
rXwJTMKiQ/CcNofds0LC7CSZHCwzin8rZZyPbRjiwnBUBiJGwFz6dyxw0IQVPZF3cjeoJeX7/18b
FbEinSkG4KbNGGo4Agt3DbQGnLWx8Hx5DWhDqZfmYH/3JDX1LMsKDQQ/MlQB23jJiQPFdZECFtzT
yt6ZklOPtJkWAER2g/Lca4oCDbBlsvNrMYyBab+U7xhftBNNTJn0yXxEK3jx9LaJuH+MGoB05CAG
mtISq7SyyX5HDHyZ6DYsXQyof0Dt/2Mxl/4RS5cEieFgRYQ5WGjaxp3vSwgyQbOHnEFH7/trdbeG
eOqkXO51FWjpbLkj54KKgXjPV4q8M6kcNrivtOfjmvrhc0vmCeNnifnSAjMwZX/FWRCmsmsULDkT
7+GR+T+leF12JAWQ3tIHXg+V4ZP8LtSa2huqJrJVwopiBt0PWPpQeM2eCumui5FSHjx+pRDwYGAI
xCq6yfq9KK0Id8VYCCOZZNxrIyQXkm3LyKyCxTfe52YBX12NLm8PqxXGhhbRWxJ8DevU3k2PI6U8
hNqaCLUg47opYxCPm+H+qoBgJxMDFaaraAdHhujdpQXPQjREnUmPKOSz/qp65Ob1dM5A8MNxeW3u
N3gJXUkv+e3+62kb7G7hES0CSgw+3243L5d6FJ2XdOH8loSHMFYJzLM6PWVvJRV6ce0vBLD2OEld
P2Pt/NedeH3enDMa1W9ovGs/sdyg2fk6/9NafUnkxZZh7CAH8vYm6KQPRXPK9aRMiiDP3jmtpVM0
SdG1fsLTYbHrObaXwD4K7JqsWahHkW/mEhZ/qTNyhWBPN9AijL0JFLpqAmS2pxqCtoIGT15pZutv
x4Q9DNsFo5Kg3O4hoMEkjEjbx9z71NsplV8ROvDZbKnGVepFKtkjDPReYuOEWxA0mInTGgdxMZ2k
IXyoF1yj3rs7LS9VPYosEYdj13yzqutMBPw8Hwk2ymC58Q2M7dcMJGy6CC4Mih/zu8HGQHE8fQYm
9rmHtg19hRdi3hmQ16BmlPiPYDJhcf/dt9abVd1YmePOKcXlx1Rxx4Da6kJrC64C40msI7V8pmMZ
9VbgmIRzGyuM33eaVU3dPYObH9hhNLFgajyGtH6Rse9KJ4wp9ATQXuXTwpieP8u3931pEeo8EhNY
X7fAxgUoryDLC+/vIg4yTijxc89BHIcrhU1N9PzKFvgl9IdMFRUY9YzUyWUGm1E9zuhxW0Umid2Q
Q/inkuHgqmngc99pJhQSJSmSOd4f1SK3Bh9DLj29VOU7e6xWC2Zov47fxt5+PYryqvK06wbwxcGg
nAx3Hs3qrGIsax+XMHvV+dtA2W0YK7OcVy2GffoNbl3JFuhd8cb38+D12Dxz9Bk7LPxZYRBQLZu9
r5DgoS7cig6aPxH+5pvQPutI1Ot+y12/F5/pKy1BXoEIGqikJXwpPehbSDwpBld7d6+VzHincv9P
yGjBwEqWpGLbvVjjgu9uf4afEhpWp0rT7ckipTbX0RWXbJgaZ0PjilTSMAB4PoQJSoiSJHd7lof6
1/8ioRXQLdSxG/PheXiqVEX0uKGsr2QTQWkN85NT1rUAGTmIT0lc637QMOANym857fyN6ZC9VoFO
Rdmfq+cXwtywxzuFFUZBK/VeaJaqWEwxXtvQ+U58sDHW3miZMGlfJtvRU4l9uSu6+Zatb2XE2lx3
o0LhZUEjjYQqSLDbM+3KsIj7ISN9iRDLnYkUi67Vdt7EmYNMogMXcNAvuUC4gUya8YcuPx9j5boA
lUW+tT/P8x48wFFSlfxr3C318dwvK+h4c6TuBAPydjWpZmouIEXQjfcyONUEEWNIm0Nxjg13KFyY
OSJnJ4FZNhKIzTXG4dMe2sSZ5LaZZmn+YpE9EQpYVrNS/DgsjMnshDC7GJ+HLplg7AOR63/HCfGK
fy6vCKL27NvUrc/+80VlCSmjfWTBRFcom0IdORs6d6D5h+efJzCnTIkm/af1YpYVhjbWKup1FQFV
fWKcrE8XUm/f0T9Q3lKcfYtNNJwZfvphlz6IDBTz0VB8J9QjCZMpBi3WjoRTZCmcxYaOnOqiNy+W
7vSkQUHV/AvkjrGHkGz2/0Hn6a0kG4FFDOHTuIxckPsTA8mUKjLAyvj/rW2z0U6pio/HwztyU7LV
6yz88cpvTPe6EBY9NGm0HNUtTr9/KGdhIhiJaqlBLDqggY8KduloPZkEgqE8xkxbowHcCKNqAZ13
FSkhqxBy1rXLtDBDHUrBFnw8EzUKJjs48BDG/A1JuJdI9AmRNcUc+qj9HQk+rFv0OUhqKOnj7pQx
pqYv2uqz1w7K3qGjTOcqeQ4kFJV/K8IqnAuHr40luPhHtuqrbp6B9FZo+cA6m0hWXqYmcrOe+j/n
PUcpSUtzGN6d14W+vh0sGBBpGo4qe7wJZN8xMY+UVaqATSqgGzO4M3497WAFT2/IpY9Myh68uida
uiZQvbfK6bJ58NSl/tJBvg4X06c47vubnDgvzjbvsEExb7V8AtJ0D9BjFUZNx7z591pWRwKrObad
2n8wViwoKeXlFK3rubwkEE/lBhMn64n+Ss9/A3TUF9hw+v9lfRygKy1fruCTvTQLLJ0Dh2WW6Ki2
5HG7vSwqKlbfWKq/OVsG3o9yZbFf6adjeMAcJhUzEYeXwISJKRo04BWGoUnrPRRDH8VnijGboolq
PvfLrDZlxujXeDtNjZplWpgEU5eubz2EssixU2W6pbkV2Wcluaex9uuJVbsF7KrnaijIpEsWMY+K
/De7yXw4A6CZ3+W+wBAurOwxf+hQLDYdimgw4bXWjERB1oeyjS3EJ6VifgFDoaPu24FuXZm+y0ry
alMxM2QWKFUeyYMTQmboUqKaSDLk9lFsgZuAARI440nbGXwz6k+T6+AFKU4TmbhHrrC/mhlX+UK8
5hNQXFMpEoFbQnMsTRST2695nY3sjtGLvnfhb0+yUrRdabDEPwdCyzYEJS/qBBAs7W5A+PgIv6So
Rlff8B1kUHMGLnW8IgfcVeVILqolzu4Mz+XJCjDcAexR6hJqfwBLwf0dQvi2b09iifPCTw2c7Sjr
vwZxGjY5w86UKwaVJHUxnaHz1XbAzAzNYeEyZKWbAjyu72q0HBTs/7N/X72/CnzxBUtgqoJy6/5Q
cOzkYapuWAUhi+NTMgRgRkiueInMIa/KzR14H1XsaqkbLG4Fl7Nfl+sEYpitib30rLBDj3LFrkct
1afgEi/OXfZTtyWbuprKfJJU+ASeoEiU+ySsbdZvFGgIUX1eeIbQZJwte+ivjpCFi/F/9wg+Asng
kK3l3ONeAXvIaD2PO+3MYrxa9dQnDIouLcb93xs1AeKopnP6nIgpgXkUtN/sNTbZ3dGnDEasawD0
DkSNWqOn5oYUJfaclA7zd7hT+1ybb/i1QZ1ayWImyyL0zNtsZhZEGHvZSGlA4Wsdig1x0dgeHkfV
UlmHekuSV0jAhqvT9ERJ1bGQxll90W8VHD/rB2RI3voT4WcfpS/XSAsZGOF7Y7COAgu60vQL+W5r
x6Rs6lUJDJIF6wd1qNCtXDsDtCBDn/DT95MiwRzsXwnTETlqbtFHZMRBCbT3GNM5kDC8HnzjLuBc
BDf9L+YSg5kRCb97O8Yl3FGBP6ODdj/ftM7SwBOx8TQr67Us/V6y4pO+bMxHFzzj8GstY0bQnAbQ
9bl9tFYS1Y/U4+bjkNpUiUicoCxIeSaqa6MnOU2rgolky/ie9ucY40WCJH7YLf6MpuEi+HvqEERk
lWfDC5dl3vQR+JxU0B5iJoWpXXeH2s22FYhnJe0ta6Fq9QaFsLYumPECRahjnwrJCQ/yUPhvDfBK
n9PIVTTZQtafu4Zvcj9B0d/LldHWn5AShS0iYX3/OIbwwHgNs3MgU24JQ0Qv4TYdkRImF9bNtoej
i89gmJwk0L9z6qcTiKuhZFk9oByrv2ooN5L36ALWeRKtEcVENnL8GbGgdp/UTIeI6urRhPac/eeh
hD2vJ+KkeVlI+bswi76dE7VL7fK7x7OokjXw5NpHiDb9aemX14/pGMqEjEGk/W23DMr7q+FB6e5y
N8H7jqxE+cGBMwqfyaaKQmdT3j3nUzEcISCpQNTiSUbVOy5/Juuz7yaCiDjeezNapPyD9RCkCX9k
h/UDUk8XDVi2QJ4A1AwH+ZzPH3dUzEEdbX+R9bAnaNlPYhhPvze5gB9pnTFZcHNrveCdadK45weY
Rmc1zblVyRe8/wZkP0I0FiduwqL7GP8IUtmhfYW+TUfvZjlZ1eZNBTh/5FukbnPEsrwULM47Otrp
zNyNfaF7s+zNla53kg1vEFZFlTCInFOUD2sTscB53U0BAeuDZ4U1sxG2y3WZ7IAkVi9xUnu0mq+A
VX97Mx3s7Oy1QHvBZu3rxaez7Lnm8tnIPgS9futzeFfTpTRvpbdD0grxIRkfFrHF9Zedx6tBysCP
xpBcuzHgmDO1k8D2EkAM7mGDZqKl3jGyOyvaEaTx2A10YlI2flAU+1zZCEZK7AYtKNP4CtHL3/AY
QfzfD57gtO00kHH1OFiy6MeXROtT7qu60AWJ9L6bmgbJ7krQ1BBJ+bhgSYyzfmxJYz6OOYaIi6BJ
/7v0hGyc3N+vXgqNEj8F41V86/rSg3JXpAjq4Y5vFfIp14uSC5N86s/nh4952otQv13i/gxyGtpV
z2V9vvAuEaGuAievm8DnvR0jIofApFvyetMlHvPZVeBwH6+EAy3uMoK/C/Zm75VsKhhx4Gs3Zd8u
0CvF9jg9j0+dNIGzTiq3mMRTm3NbchqviEurN2xaLQXxul268AgxnviDVMR4PdPmNMKQelH2gWvS
UN+jgBxuc/K+/oa0nwCxRq1v5nWptSp1yeBUK3NXO3u5t/12e2GKlEDGjFHqWX4RloB0WOXiyqXN
vb1GjLNyxhcYliIxV/vZBWm1+I4IzG/BcV5zbsmQcTy3l36WDrY2lMQZxkmJgutSSlqUmQOR9SWP
t9EF6mWkeJ4KeIHDwJ1Jn+QhbtRjIh9n6IWOwR+FRwypJUcAmUZEof//dlXCgSH348+P9bTd3+GT
ojXoDUdkOaX4h7sCfrE2FiDGIMtzkRlKbm/+s8I5yAgiD2Xn2GpXgTj4iqIDgfZb6dU+lU0fgM8e
MvLg/IKQbtCIy23oA87qVMZgRHoTfcmuhZDEF5vn9/5f45Odx5r+zgUXEFp6ns98hOblhw4ETwun
Ny3lGUDtNwwWewXHg1GLeMwv+3WDoUw6CXr7d6iSQ4Rui4I5gcOWMtndWL7fc1DIk1F8mqPDpXcE
knDTn+q0E0tLAOAsHqxXQCdRxveWzaMOrYOpt9T57ZhNlxgJLkpQ4w4bnjeeSSoFKmzith4QVuJr
UNLD+geo07Kyaesu7I2mnDwsr3419W6bSD0IaMt3buHnX/IZXe2dzJkfcCl9I2FThYFcMn9RcmHA
EoNIYudkxC7mt7ud6fs159nYyXsOgleGTJRlWu2opIf4mJZKBrrro2n1jBniY8pKVGYkK4OlqtUv
X/wZz+2ucgklQ0+jnLO+yIZfvvKNyQG5/i7l8rCczP6843yBaKuLMKLF2BiGGNbdcKOGssOsDwr+
YSjouM5R4TPjsy8lBW8wevfGvuTBcPHKClNM/iOcVofhFM4GQw2zFh+6s3bOkzJ/P/HEa7ty0KR4
UnDvbGRPW/kLcDgZvt5kG5767dRAoiDTXr0KzLcMPanJY9c3Qd9RTd++GEkwECd3dOWr0GIHuaWM
Tfl60U+LPxdpVCXTjwmTZ9wEAHHXzyjknILcFvWCidXYxL1y1PlFbL1c4wZfgsnYO6HaYzg/Xofu
FuD+62/GM5OAMb8NeoIz8xKvuuQeeeTVtVLZ7QnKCcRxR82YUua77JNHiuLE4KlRL2SFikPuZf2l
Jkzd6e0AnVs7NbDM8AfZWjCe0F6qDAKk64LLLX35l0bVS1JMIf4tHdy2JblPxBkHzTuEG/yWltPp
S5ZNohW+nfKR/oqL9GtL0GlNQfNaSLymAFOJgonmU3HVVqWbhkYAPYHofXBlIp6kK4hUmyRIJeZl
7ErIL6K+W2ArYW9J42jBuPm5xxJVfb1sVFt12CUar9kx3yb+G2hxEyiuWq41qqxlV8MplXSsBhrY
clYWsrtQBG3RTsMTnlBBFIzH6tT/Z9Lq9TOKzNoQSNa4kY5GvBWa/XwTKIcnahaEBaqLPcFvtC/x
Xt9bo4gg7iamPE3Kw43N8yKm1gnVE6QyqpNgS6+Jmm39L+bnhQO5OMEqvbm0Oj4T1xiSmpqPa4ae
5xQ+Ev4ig4W/GCi+/Spj2oisZHAs3jryS7aTkHds8Q33Zxv89hNpf9gHi7737wcQ/dqTNrn/ST3N
m+B6TldxRryUKQ8LSaZwKWToznRAniJAmmpFHj9Xl2G6WNMNv/qCELu6GWly/DNBp6ffajjmifuN
GbhHU036AnLO5CifUa3r1gtAIqnBjFuafuRws8syS7d8+T0knldC8J2UZSawJ7Fp4ZZBGs8MeWwT
2sGCzR+vQQwSl5wFi/18iuVtPNsR9104vHsMr9HB1hkw1PJ64Zgv0gTwvITb4aIFqB33gMgYaAKc
IADy3kReTAG+ym9OhJXFLAKGrRhe8ddC2f1VYMi8ZF3vMvd630cBkqVtL+erpSyygDOYb4HZ2sBd
ORGonw10Ri50wEw2Dq928W2qlWVAo6XXE1xTODK8ET/IvCVXeWSghONpDyAyXEKjUs9+jJ6oBy0I
JZF33H6g8KMYUyFe9b3fBVaoXFqx5/8LyJ68sWRNduU7nLo84DJGmDh39riiNnlWllIcH60EZlYr
aWjAJPGvhd5ViGU/RSxKPZ2PpQP1PjJEhnDUQphfyIgc9IygZmshwB+I+Yxxt+BpauEDJo/m3Yak
1t03j2iv5qAL2+4cDKzuHp2HWAiU9QI5UE2FhRs7rHna1pu8jkzCYTdLY9UP0CRIIe2BBuMWkkal
DRyOdmjngyzsoSrND2m0iRitqhehBEySzOsYWyCYLzitvFyMyKp+anfmJY/FSEeLBl/MCqip2enH
lJ9eLnHeKI5OPmrGBLuLoNLmI9aauCooeiFWd+mDMtO26iHYroKrbL+XD35SJ83EvYsF4/Qxm2ff
4nkHvrt6D5FOHbX1KWt2Muwl8JTNvP+BaVTD0ITh5hD8uUCc9M9jjA1mRq1qPXNdiFSrXXEhOWSa
EINZL1C+w3NnLVd795L9yybj1ZjCGiOJF0Le8/ioD+6cc+uEszNVM+tiNV7ZI/l58fas1cxbhJFJ
sHciS7I2wnlaDFhKpwZd6Z8V6AdCOZjZaOk7WGQ8ipn2Rx+KQm+e0Lf4YRutbIYAs5AmYl485MES
ngYk9SyJQLfMiWw2GHbM2zJhZU2S3P+qE2ZuwW+1Y+3necqOl5ESoaIECexrvOgj0RUYPc+4b8Ag
zGcHvVP1Csaxm2UKsBOrrJAVIgs9jrfJu6OEOlQza1WQUlpVhDuqc7U/aR4d9bp0xY+KOY6pWgh5
2l7ljLnqMPduGbAaEnC3IORQ0woOm9td/dW67y6aJw6thTQyJ2dlhIlqjC55fRmBuTjoWAffYhpp
4WUTPP464lxXoEmWEx+kJ3m2NHhncqmZ/KqBxopGQcHsr0NCfH5AGnKGGpZic70uCrR8lC0C5jCb
LOwOKAh/Agiaz0TEJ/h2ZtH1zA9HQNGZliK4wpDcW9IDpV7HRWfBvItpR2l/BsrgkEkamO4UFrbY
GqdEZo+0kcMHNe4mq2bD1ILHIOdE1E5WZzR6ih99PImmRyNd/ju6xKppNB05mw30av+TOnpv98kI
6koFEtip39V7vNRdqh7zYUrmtj54Mnc3GJk017HxlMHbzNtf0epLLUfkZwF95E4OittSoS7yGaHY
FBrdLqb97FBtzxTl0rULWmT/iBr0/ZogIagCcB/rFzvKSBKs1fcYwKzMhSHPT3vc4mNeac+Olkol
HJsK3g4gqe31y04nbvF/LfWX7s+bZZLeArMQ6GmkN+E9TqQPX8Z63gr6nrr5yI4VYg3VcRL7C2kD
TJFfSdabpQmQ/s8Mh+aq12vT7tElDqn/Wyz1bDIPEGs/MdzwryLKEkAtcPDVctnNjfisSUB2hG/Y
7ARHwRMNPyNCH32PGWCK/xtc7xwAt8uhsz/lnjUl8q94xHvCflgB0qEQeMHkQf63uPvP98YhtZjs
QW1c96lLpaISQ50WzkdRk6uv0vpe6oL46em0xpUpxBN0uIJvCQlhf6I3GAROfTYBnpg0YecDGTJ6
T45lhZUtaBA94g/7OsQXFtA94urPxaPAoCFiuOwVU/X1LKn/fw6L9BM0U4YCrtnlR2Yqc3vG9Zk6
LGgOWur7tqaCfWah+5P/vyIGrvlmE2EQjbYSA1GRbbMjuWmQv86UT5pdfdUZ84btSfwyESMDXJS+
Bdui6sZ8KSGmUThziYXWPTEzBD4BduCAwAVHl3/5fNjY3fawcoN+sTjYpJ+00GIAijBLIOJk0tAu
N11fkuVkmIab1QuKGV4i7PP/9PO1nyMPPuggLhJt2I/IiKgQfYtrDuVyZUzahmPdqvCV6SJcTHHT
iGWaX67oaC275btSSX9ZHZ7KkLbW7ahyLCO2U9ROb5nRgMEYPNHnr4IdD/1rSD0yl0vbv/s2vQWh
9epvII/e/T/WBorT+Ct3hdx9cSHY/agl03eZuAAi9qNMK7U4H1ZjcFuiDc2awYZ8/PZAFsYCuVuk
yWd8F2zHcIGalivZsZiZimBzDBHtLJMbkkxmDO7DAznWhepLZZuDZIzOo/xO+X7uNK/gFoDJopVa
r/HyjnFwgePwdoTRn2z9EKQwveRyG1g2lOjdacOoKJAEX1zv8heVqks37jQmQLpQncgN9V5wq+U9
xzDhduhvkhubbLJxzkO7hNHrB++GCzataZ5OqCHSNlFBdaPRAymeuEJDeajCyK6v/aUKljh7uzUc
v08zUKf3Uul8Z+mj4jV+ASDKG7qdCc7eNHd248Ljc/NsFwuP+acI+te2mhVvmH7n5YJrhES69R5N
od8aR+l66Lf3MFHCSuVJcUJV93Bfqii+Smftg9ORrFH2LCCdDQrB9/a8M2l8EwIgwCKMGSS1Kcjk
LpQs7GouNQy7ufPsyV31xp/qmkN8a5nO3AxPgx6/vwGEIO8e+6KHOa5GY/O5/OQ2EOuk2INil0YQ
VIMzy/AGmi+9ip/UW9npZXdUSFwOdUdEExzjP2PZhmtg/qE8LCeGBt/2PWMaDf/LazLLE8SzTRXp
78WBzg86OujQHQSRmShqilsy8sMpF91Qqy1RvKG6+HKbyUBGUz22icBndc6lpm7XcjL0WCE602pD
aMMS6tZ7qCtqZlhswDjhCQFY5q///rK/HqRiZOF5jgg30Kdpfpqri4yOgTMfPTz+LxpOkCrBxnOt
iaoRbVqfC2ElcgOXwSlCtk4glhCAfBZyDXB2LGU4HSucYHzuzWqjtdeVDlTM/PtkYGYRkIfrfk0J
mzpttcZdST/jYWX+grne1wFTize2guJFDpx/YCA2ABFjQ06R+AeKHlMM1zXVqSOCzPcjtHEsJU7g
rCFjC9yHJZg6MsimpjrKUh86KXfltZZVrrcPT4ZOhs0DT9SMn8eUXlEnfCI7V6LViNgSrFXZze2F
1Glbod5K8awfR7UefMSdcuqVAdm1DqQSS5Ge4WLysJtZsjoNMGEPN3t9mvNjJKI4YzydmfT+vVqy
BjpjPVkJt/qtcScBv/t4Xm0HG6oqJDizyMtKBfGHaHxuuv47Dm/iBAXx/jjwjNnYSLuI/wKD9Svm
i2k2zi6pXWYPWFP4PQikIyHCb0wBQbdl22mlGvYjeg4R2hRnvVaON3sGa/PmCgMYiR4oeuRY+6pg
AyTG+Ig4QJ3zRXkDI7dPDiEFvXigNxgLdwdiustEgq90IJ6f7qnRxArZUQKk3hfjj6o2ZP1paSuS
hr4tFOAI22i3TVHvZXh5YpMW4/q3lhM3u7hidNwSHKa1G0+lPnyYJsd7ef2aQCKjMl/yjfcBNraC
1dLQkZuvxcTs51fXLPNoqDcjXgMJBLkn2UrxUFDB4Mv69wzIWtXG1LvxdDfstfy6yFfYrvsOye4d
RD2RQZQS3DNCTchRv+nrb6vtPZ0E+jaZDvKmP+690spAck6OwdFOz23f/J1yU0gFyQkFcAQAZ+Wb
/cZz0LMigp9Apa3S0rgc7BjaATKBxPka826o5cki67wsbdM43zgO5VnuJE8U0SjwrkqIwJHHp868
RvmrpucUT4x0xZ9fw5CXlOZ4EyREPGSySbzdVtNKFnk+zY4fp8N9qJ+4TyexjX6Awysc5gOpqVHC
+vQ3Fdmgs6+QM4E4M35BHKEs+viLLqSXVf0pHuL/NMwY8meXBjdx76zj/csn0Z5rwBidLTyS3jn9
a6StC4iHZa7BMtSGMKAk5mx87GbCdtbeN+zS+k5g1iXL7GxHDUT8sUKFKX5quWLedLBdQHSz+Os2
jyW/ddeasOBG6Hq2gZI17Gxo7iNyT+kKhbqa0oY5yEOzzpZoYPocdNsOHz1977oZMyky+75nACYl
sas9n4rUKI2pv2Z/B4QOV3VgG+vgTH06NLiaFyTLiajx+NgaR42Umrs0aVIiSIfFG0pwnXU3p1Ej
l7mUxXHcrn/VI7oGH7G4GdltEvdq3SIqd89rkpxU0YwVQOJV2KjjwJ7wpBeaTR7EvqqBJFsEV8gT
wzeWFsnTPiWcogtXdPLWXEJ4GVkaZjm6AHCga01ofUBn5fMGLg3G07i6Nn/XaCB+INfzWT5pQFRV
bj7sYL1S/XXE6GbeF6aLtV5DJvrhD+ic/FZRE3vxvWRoROyT8GNcVHTwPrfazaHwQF+3KEvO3AJr
FU+7l2yebUtTuQUnhBek6ilZTjZCkyCkaDrVCPY9/52o1xlTQ91LicKH/Y6NZbbhtFnE6FFkLSFr
Ye3TcJR0cbfSrr1+8Rs6aFCVNffzKZTNgt3XMa4D7szBKgGoc7j5qApu2Nnt5KN/ee+67a+8k8Tg
L/XIT0aoCAA1C0x55G9WJTAD4jb/ypMjY2XoPfD/ZLYmOmIWx48UvXfkH+F8aPwkVPBOz8Vxvj1s
oCcYvXvnFLt2xM7B/HRiDcxraT53JTzrRSxCXOfuuzXTSQ532VbsBaLCbiBUqTYkKjTTJ8XDwVGm
FfOV20EwZY4bX4maR+wHE1f4LXD7c3OYbODu4riyXIemqoV3lUH398bJXAQTQ1vHrKe96YPS5a82
j5V+71S+1toYa/NeSwHKE5hGnLTET1Grpu+W497zlyzUmfrrqaEhXMG/+aeL4dDgrHOVTPdTCzAw
yV3PRPMY5sgPSIwMsIaw26Ulg4J/zYs1BtAmosdtIPmKVhaqA+qo2J9NAKBPUVlL6qB33Uhe/0Ba
XFo3Xkw+18+oqebzwlJLHUwm7NOWoFqQ3qPaig5RAP1OWhkNQ0+IwvjsUrf15dIXSK/wyM73VJwy
vVY6Oqp0giVj76yvzAMHuELU69v4+hUFoG9oAYjVfD2K50ZBmkGu9/BAUMas4ei9Rn+o1WFMctSl
wPDh09yeX5UdkALw/aH46ysJWkIH/B01digDIv6w78azALfU79WhPLvQvy59QPaf/BAdC0JqrZl6
fVuIrDmcq4lxIJb2409mP8Wsh+A6f5U1kSv2V54k03jaMB5YiP3F29R5CkQmNKhKzzGWK+5pDBgL
vlm7YqUE/NpRdQToe9IIxEx8Q/4DuLE7Z+rEr/bFT5UoMfJ5ts3mGmk+sCHJCjRhQ28Y8uvD7OsA
oNlifUTz1szcxZujzwb2o15UGn5jrCDyUNRq2uZvBbhfZxVS4xkSvjt5IvbjDAU5qJN9jOp9HolB
fn/qb+tbhhpeGmCn4Bk/wQ/tgK+6U3hsWhRzHV+a5dPLrnME0CqsKmDCZHOVE5QYd6E1qwMheFev
UmSGlQMmP6Gz4OrjlbNrcuKb0XNHvPiQ0CGRKej5VkZRDPVPdINLZe0+S+pggBlQHnM6WChOBF+e
cmpdqi+IGP4Z8A1v8xSexduQ4jx2iVOYmx22geLS8RWICJoeib8D0qfPdOhEaGrupd2De7kFBl+4
XT8PhqKacWv3n0HbfaOkivOFCiiTzo/0AvoUpYrFPEsdfdx9yNQB0VmTWyYZFrzi089oXrdVg70w
So48bN0ZKXRfUUGAwnqvRG1ecotoSmdZkQCg5vxaizxIOTU0n0E12dyYcwgsixJFKKZ5InuMgamX
rDoa0v51HQhS01DXOJQybOsS+g14JoAYcVcEh6eYFV2HlXf2OTBhqGOi5hg4Km5uPdX0HV3k5wuy
Oh/6RMF+9VsptZ2B6lBE24RD3R6fHiVKNPW2u/PN9WJfjUoWinfZI1FKeIbyG4VPnxRao3v6Sr2V
FjTqTzUr9kVIIIec8drdmUUqeJVhPAt/7F5TTEwcLh+nkNBIiE6NWXROZyMl09AHkIu92yAnWDbx
rBYheHzchXGg1wUkvq4AjrFiPsgufcZpFsPi3XAQtMvHFmad9Rv2D6gFWnsllLJV8MCkkDdP1PrX
B8AEvMDvLUv+jfhrlM3sJALe5Tx6R4bpF8EfEKAMUoxIGc70fAtZdP15Zy4BiwmYmet9em+gx9DG
Qnh4fotwqA2U7GJ+EuGonYIbXBM/s6PxAb8mtUc3lffJTYFfr0ll3K2Fr1+bAyKq4XsnNfI1hbVg
7AOlKd6Lr4t4oGocvDzfE0zzMIv1Ta4wYNBaWyVBOX06FTixJtOG7D6U2klNnMiT4/EtVX5a3GdK
dqUOlWOdd2p2JsUSpDayppRtcTCsft79ZZLVaQbNwKoLLEyWpSrmZs0bFKLpne9vZ75JyTK6j6+x
rOFutB0tq9ReXfyoJGVcMfLvFkNfyxx9czar/n8rVkcDpZlmePOycfzc+Z/Lztls/UxwMF4PjuzO
dk2ftnZ79wCWDsQraLkb2LvHwlDW2K4PHwEZrbBJcfSvTHsT0k80OEShzmBgUQx74FyELS/MnHKg
DeECfrGuiknj/ICRp+W5IQbLfvnt6cj6QlHZIRPOA786qfAenGB+kx/fJHK0KQuCIaWy4PY7ymaQ
S8bcPrneMgywwHGd9PUX4UYPqhL0TTbzDtyGql5MAki0En64OfH9SgSAA9Cv+Vw46D7ofOfgH9VF
xjykJze2yR4O6Yn66tl0tzymk9j6P6BsnFDxzC65vKpoFah1lsfxJ5mnqEjF2miIYJ+qO3W7IVN5
568sO1gTNJG76j8uSG+RUnw3iedpwVciXlpjj+yqTe8ncAyGryN9oo3oHelCVlE4aVYwC7zdhDT8
wZi0mG/uPiHCZ4N25DJrntbO52rBvMzpsZqgys5jxBeobHTlgqMbLX9Ytjh/o7/Xf+XQBd2FdFYn
iZcLGmjoPXBaTndbbGU7aRTzLpC7m4Mwkw4uEFGj821r4DVgAsYFXFvUG0yAUtGvi3uoYEeFUvTX
bKH5cfiqbAa4nPb05KtCoe5Z814K29FdwSEb+5mDgjLgx6xuKjDCbFW666kUhRoMauf7dg1pyVU1
bcvRIFoOKaNomIFgRGrwW5V2nqIWY6jTXHCLR8ZwSpcdU36OPNh+nB8eLIda5/o86rKl4TFD1wkY
eAgAs/5b+M0eNpalGuHNizN9XetHe0Ah7zifyU67UJk2QB1VtE+Cno90kXfXuUfgtUattsZsKcCb
q9qwNZ3DGLg+9WsjZWeUQNbw9kG79n7N+UHYLhI+oz/ds+lFf0wogWHiXzF1byppxhBCkHK3gmFc
X94sJ3rzBQhXTBmTS0UH84DS3cnRT0jKxqUB0HtS+2vb/vHIAH4AqioGd61ldubMRW/6KEXn+H1x
R6yGtKmrr4tMsM6byKJgOzaVB07MHDfdKjTyv1Ss4tdbo9udHl/NVVljSwiUPhSAvVDj8wzGn1Zo
wdOCiDF9+9S9Hece8wOuuEP5I4OpNAa6bjo1rL7rVvo3TMGuk7bMvQz8QkB00N99pU3li/kA6+tj
gtjq02AdW8Y9Xiywl6TJ+W5H7Oz37VTA8M3nb5dTGQ5vHjGIvgIxUY4Fm8bnDjpeo1cXE7aDzdye
XCun5eNlbbJhSUY/gaAUKtl59DA1ZTJPiJNyOP6SxB+fZrebvmArTi6s3UgdYRxS0JLZa4ZvWwu5
HDia0bFM7gNwdvhHDFVfugl9jbOS3x0p1sQG8ZJqNy+sgwkpDdXqhXXX5jlFXr6EUysK6zu9d6PU
nW3vt8Fl5mSkMkFpZDgRoHXo3lgHuZzNe0r794bhuE2Ff/4Oi07VoT+blm4Obk6w5PwBeW6zPwbA
tSvgVDF0CgwR/fSW0ymEQ9KOku83/e1uoR19R1lzF3rXUsBwcVbwoSa7iHVROYp62Jqjub0a03f6
5AFLEZIivX7xry81Ypne4jR5ODWbhe1knDPqo5wIBP/yMfra8egVsf9GIOna111Pm2i2lfgWiKrG
oIl5/cVhZnveNNapS+xPLNSkkq2XIzkRtvG6u9ClNxmRmbldKQN7XIoRxrR4+OQLT4CJyCkCxtQb
Gwl7iFBX5eoLaaJETnjXhl2y7+t9ohJr4+phrm2hH4plps510oYxIJFACDEyxTIwkz5aKiVA5vAx
4VQ7fdqr/rJHUIf0Y1k1LKKdNRRSN6K4AsTyFIJF3OE9UwN3dPowWIDsvVuW2YJE13Slw8WRomlC
1wPpNcBLFWsrXZE+M1VPdjkA4pjWz+PsKDQ3wURIBO+8/U/fH0lxIUFAkAMIARJjSdl9eFY6A1IC
iiZRlwt9MHvJuW+xFiC/3I8+c2WPUMZoMbJDYZUn5xy+uWNdrTGUyvfDHloltTaLfgPOza9GgvJM
XEaQmF08BO9hbKaxVACdbew5ZJDt8gN8X6Ety1eqTJKAeRf85OkURhwxl0SQwjoHLtbMqCkfmenZ
KFypwrF8gFOdN33wDf14w/beMLPK5XIas9zu1/o/+OKSfwK6T9PVKNSWkvLs6DH1fzKvNSz3TbTd
uLdlu6Xu1PnIQzytnu+eAfmiW6S3k8d4UTiqKqBqYVyO9Zw7uEYjd7qTgNYsIZk4jMHPYDCCoK+0
JF+VX4h9rvkJTGGlXRSvVMwzrWIJ0/Gq+QhVng/qB/BkWZaElnuITxhkwYJ941nmL6h2HoOTU81b
ceQzESVniZSNQMNwE65Y6MSKvsvlWhNWKc2vNIn3o8UgUErizuZFjAX6u9xwkLW9zy5skD125O0m
ubLX2kKsA/0lg4/XX0+b8q9AB/Ac7egFDZiCZ0O2W7KVoG8PytdTUhemUPwocgDhZOSHE7HTtjqC
FP641swKWR73tIsTJP2EeYmDpIp9+S19WVY5MEYg6PY51QCZmmYvjwUFTYF5RFrNoqHQHqeiOZ9b
MRbK95z0m6iadbnT/tkzN4gdnju0M50WZ8lviPXIGgGM0e0UszGh2nb1OAnRilje7oUbAN5R+O2Z
fZjRD524sJTJuYTmTMJttWYRKijIS1FDMG0QQ5U1zl6giIt0ADtrtpd2BnqMSXTPox6JXj2qGTEV
yT5OyR2uYECOi6qhToktfgNl4FHW4UiZQxk835TZd5n5Fnq6Y/sW/D0SyBfpiWel151OR0wfFm6Y
7bX+kI98a3v/E41MT1lbjtNh+Drf23SyHRBv/Lp9u0BDvnkRQ7XPjUKQtTXMnoX9Cc/Wvz+2Lszn
9xHAj7SmLiODwQK22wXpazavc0cBuVuvx0+U9ANVkGHO7ah4VagmaOTziM6aURXS4YglE2Wylv4u
dMWN3grxT9EWjK4uvilGm1B54GYYv8AJVp/zI/SGCd8JS4HrGnATF2zUKbcdxRnGaYTCDncWaSxt
W5fNoTiOoYvQ0zRaO0tBYG6qDklsN1espubfZcZEyQf2eMXM3B+Kv2uy5Osa+kzRi+3ksVzV95qc
EXNvD0qLh6ui9IsTloTRIVb0n7TUbcZ+t9VSiRFTVICzHRgKj49SFDrc3e3tVO5MdcJWoDdB0msQ
M8OiJlAMnMlzenHVu9lXRM58nDQvwoErkstgOWNo51k0fqlraeyD1ZOIJsPbHZPSVcpQj6U39cdN
xOTnN0p63Wg2BTOGJzAGkI1WsbAsEPwVNXMMRThg3/PBKhopfwTtfxbysmSbSo6D96BaqIh2Hb43
RCIVFkzhgOQ9L6D47CFx5X7GqH9AGy5HMPLBkp+sxZvkK8tGu78qbe326c40ryLJQRiRjpZJ/WBr
hYblSgaTFDOMYLLni5FPiPfa3X7cIrTZqOFUx7KZSQQuNNLc+jaDV77RdRcPi1Uk0WZlixXtvWZp
fVWSq+p5qd49G3h/w8ACE5cJlSznrOY74BVILD5qCbTEjsKjdfRgx6ZGAJn29pa4nBe+EJselH3u
Kf4WMBhb+QrvdZ6dZt5cLAqQITqcUnojLg+u1jMZvwkiEFl0LCg4CBmTshAmx+ei4O+Le+mSY44v
gf43/NWerk+Tzn81mzQFSdA0e9jtD+drZ3HhSSodRzmKS9Hw3w7vuhsAL1wj9PwKehmcJ0WhDQ+9
NZrDIQRDnvE5mUZ4BMU+Ehq5XVRAwYnKHP6XuIUHppiXewhm8dDYwYQ08+5RyNPFDaUBs4u0M7eS
OTB6jnfKEW0ZvtsO+rUMrklPZUJXq/R6nJRjFqYzbt+ZPCoKLwpvnqGy55RUwAozWLDGfGgvXigg
3jKfye7OROWO98Q5aoVbX9HTAWbsgDSpDtY/3Ak8pFklc4eiAzG1THg0o2CHpFkx0Jw6YFErmExJ
N+TEC+HftxlnYF9VN50BQngBKZ8RL7BG6NXTjOH+LbDNe5ZSWpoSlEHcZjN2THnbJzzJSkpSIRpS
6nG80+hgkwb/qTDKS3TUWIUsEuCP9DmSbitYCAoMcdD5HC2oHwiIvFQvKhP5qbpj+3JVQyL/pezj
hhLavhiR7xV5eBf/atf3yJTQwz1ixVNqBeXNFMdAH1mo5s/T8w1B1zZ1JE6Qd9AeHP6G+5fuaL4S
KWBAA2Oy6kn+8i62dC4BhJAAvJbtyL9WK6GkLWEu/qoITrjkgJqIQ+Ad9k5LF31Q/sjyGrcR+2/8
185IPr7vbSKrc82zzYx6sdwu5p/xOwNSWbJGYZGsISy6fvVmIht6KjD7V+RdRj2Rh/oK4bVKkYRv
yWAz5IzNvzvIQAQ7D/FgOujprP0g1e+M+EUBP0Z1B81JLiu9r25PqBS6GCQpDjZbgwL02y5oiMAR
9WgKQUSClU49PeDaNchNGjtzowujnVpIvlB5iFNUCMYQSiafI5AcBDB6Bn5qaghixj0fQPhK3Z0+
Y/VQrMXOt5ft+GVdw6dYRGNo9aigBp9lao5aF4DnRM6J4FytZsyGGjZPhAT9FAp/o7Y1EReIxqsC
yh80m13KzfX9VrHiwRl5e2M+lxyLlNhPwO9i9tl75U+4WGuP23jUDb/zEtTXwR8Ja34mh/qZkvKi
6HFwe5SR3f6sBXr5Us+rZoZp23tSU3dq4KrmUzvInrN2HYrqldUKU/n4WT4vUMYlJT3Rcuf8baGz
L0VygqLR6cJHYJUxQsYgzKJ/pjD7vxKN/KmtS6K3wR9SXRKcRo8T14nDozoXZB/gmyJS8nPu7R2d
dIdhQXdgL0vYEvyW6ENDHJEzWKmnnF1VrKC993i+uSrgOTN6js4ovomgnf0qECmpfw2TkPXgbtQM
eOkL1rDeujvQCk+6oDMGeXyGb3Cvl0MwbiiyVI+Dy7ihJLIzc1AdfEm+uRFxA4upcQW8JxdZFOhm
pKmxMKk9ai0Fe7lqCfsVSDXm4U6kfzP2K01vR0RZ10A6j4lQTrMJYiM8P1Fb2q7GbSlsiZMtQZke
pKJoBb3Z+q6SQl0ZJpgSZXqcOVD+BGtrVSG6kf2yozdBBMFNLYC7NeyM0+PHxGUQ3LwRgz55bbp7
Xmq2zDez8A/mw682DTrUs8vPHxtnmBI5aLYTExE6pWjfi3ifq7mqYTJ7B8WBdDgG3NFEs2in7hCv
GQUCiazFn67XDFLtzTF9B0EecKwZ0ovwXomA3CA2WGS4+zWScnAkkXhu8t8binvuqxmAAo/iTxRC
LQUY5Ou3DZQIqR/087GSa/EU3hpKLp96QJl/It1aCdtRImaxkPtC3X55W2vnJezAlB2cmHxbZQic
fragGaGI6do+xl8iFao+P7EDiRon5GDTaMrhP4e82wshn7PMoPI/00/0whX7zb4nZD8V5Z8ptp+s
M71iyHMYDo9d9KOCjvDFwzKJPHwz7zBf9FQQV258vrgNfcLl/aOw3FHIEwrbt+6d+pSIBcvLqr9Y
BvvNk+jilyfolYszNDZbKW2C9tjv1EDX9RButOoSJwKkTFA2X4P7yhdxsiqZvvL6HAKLXwAZn+Ag
Trgsdry2cta2qzKwEbvZ3iSuN7WKUpH961We+nbhOHUc8agNQZTsjl6joZAYzs1pkhivooJPsDOI
nXz3Gz7xjmh1XkOeP0SanYNmLlO7x6ZjuRr4mH3Y1bQTvMnpqDq0D38GYkMf65NgGjB7orClrbHP
K5Qw6ijU//VoEEJjC/98JFSUzi/OjdIA0xBsrVtJEFjHNfnhJH0etGp64J6JWjEw7N+YXmANuEbw
V40CQ12LPs3+YCNkvf31KZFSj7pc3C6caoG/8PCJV8i3nd/GHFwgLuy6Z7TepKKHqXBAjWTI7KEv
XBMHicsqZGyMde/76wNg5cAZ9bie1hov/B7rIR0IEC6FAvqsMj1dao1r4xricLOsyCnJn/ct9gwl
1xU/EkEmsCgtyRS3EdrcwlyxgxrR4/LygaNUaQXbPlLP9TcT6l00PPcRh+CG5jZ3NwlZ8nfgQFGG
I9c02uYZKtjUHlc+WekQzoXmpE1plm+V92uF3rzKg+CW6MgMywzMytmmRzJTKVYUAkjnqUx5ehbi
9jnzv8QlKqpwMQmnRawM3Ho+GUcHZphNfBDVTFmQnvKM3YaLRfr9lhLQdv6TCRupiGyQ7fr2Vwzq
adlasvyUs0KYFzFQ1bVjArK1Q5zJBaTCUldmBOEVK20G03iJgeX1PzcDso4NI1WeJyQUChtJh8bk
FK+8SZKypPHKJDFToETkPPOEu2VttJQAT3WXx60zJ8ksccRfrCzNus/E2JDyvQ/C0NA52lf6Bfgh
5g9lHiqJf1JrIwf/W6Hd/dWmpzh72Ms0SlBWiTOh8T5UtcTBemNIG1OlMLduPHtc4Z0nHXt2kgMm
qsqgv8gsrAsqHt5ZtKraWD90E96Unkt3YWyofuOlTshPDP6lHAAOVxxtDUsEd3iMTpqedsbDwjQN
aTj8cfBAtp9PR+cYfXWOvu6DqHJu2puvLsU7LIM+gheijX0IvtQ0ZLAwqhBEOizgTE3SEE1iVdHS
XNIGTxzHgN9XDs1ouBUUI1w2Aup6otBhH3lqbKXyjPPxSFEY/8oMf0sNeHJBoO62Usy/2R1zSfua
6Bz/MIzbB7IkP8RrUkdMw/FwWe65d1Y55lZf6zSJ8x5cXjeO0iRVKg6sKyyQfTMmelI67rtyLZpy
8/5+WdPi0eZz+YtujFHJQq4wkPa2MPtN4Chq8sKutOkxL/GypkqqquZCB7xc2H21tXDHdW+HSN3d
zXOkcyScKt8X42Y8HQpWMTvYfdYa5naYSEgY2IL0aKH+1uH7utwJFXs8WVelhoWuuPxno8Y48laC
vjEO6IDXZ7JGml05tLpiJ0jOHOeTRHpvxYWSQ7Izdbq3cbNLjbZnej8pwz826DLC0dThkzzCXNyR
9DyX+RCirVk368YBv+B9gUN6pgUB05M0hfcnijDjRhK6QnB270Z+KAq00sXSLd/kqAUqhnPAPH83
TevGd6OGcVj62AcfTw6rvhx4beLu0yN6l4Q28HEcuf33paepVEZFFW5h1xlt/b2Cr1En3BQ+MfA3
JDpd/WekRErRwAyR4W2F1fEonrskWG+KXgJLzGSvB8o0U9EOoj6PyhMHuZoX6HKgjdKDNZotinP6
7oGrexz6uqTbO65JQFnK/pvg3EhnaqJ/f9hq85j5DlVGZJu8E4m6Gm3q3SnjFXdfVZo8Wr4vnkZY
0Au5Yp6XjVtWJEFKy1rC0E2BhaqszmVoDVDfC8MciMBfKx+RA9aM9SbEgZqQbzF66Dv+s+A0M3Yj
AOxaZodh2L/NBl6XOaGsktUcFdaUQHotH9FjNzGG78uinzxyFE6AX06Hw1Ev6iJIY6vI1H2u4uPD
HGjaZfuTsGoav7XXmI4AGVZ/jMJZCJoLLhacQjqonjnmQ6Y7wiY+OwMEJLeFC2shEpRpHsqKkF1t
J/wVXKbBkH7LWjxU4HyY6cIk+R4+IC7bsRREm47AQZ4IQuPmXCzfOO7tUmtfPSvlNCDwm54+sTuk
Xk7xBG3mDN895p6SbLB4bDoM+epeWGNGsioqtkqvmBVZiaVrhM7UxmrFwn1u8sB57pJu+ZOGtn+L
XUZyzGdSr2x/mS+vM2Z9ajI6HiXerReMAluDXpBYs2yasnxBD/xZC5+XB9debr5ycpxgOmDII/pM
4zDczf2h20c+sYwcjXscx0wqSjhPoqZUEwVOlOWKkQcqI9qMFcfVgshzEfAbMpI998CqXBK50zg2
ZM+0S2ed/67Q4GAwY3qKgFdweeyTSPXXBCbWkdaucMyoOJENwghPzxS500XSce0SpbzD/LGDm93y
1u/aYFxurs1xf0lzQtK2D19bLmCcG6n077/uUO5CXYL122Ja8uzFlUUQuGfDjqEFcz0WSSBhoXct
3M9j4Cyo2b1YN88kkBBnpbApjmfKnFLbTQXeoCfznjx76VwdHTL1EgZ+NOiys+tLZgiXaz67O1ul
Ayb0ztKkORDt12zUSxSqtr0z65ch/Sk/gIz/5LQIKhjg+i47MwXigwk/t4edizwV8zFDjaUIg37a
dF/fEoJrsjSrAuaNuDnN90dJbQXb1W7Ds6OAHlpAavkFSIWq60Lnp6/Smx8P2niaQUSOaqZ4AL/e
B00UnQAOu7ozWcJHdEon7txec014NfxHMivG8qkm6TjVXp8WTjJxTAiGbBVvsoxB6ACvMCMwE6IG
3bwn2+qFWYNGOmuMmhDX8Ok0AFMd5ymm9wjj3bW1KqN+wLb9C7t92SnpZRjjZ8kK48g8hlOQfb/F
qz7Q0EYM8O1uOcpawO2OQg/A76hrkhdRSA0PXH9tWsx10i6ZtihNhgcfh4drLZ80yOJty8bFEXgj
6QLzwleRLqbKzpK1WGaS63rqyZJUXEbT9QVd91zQF6dr4gONG/YOvUMkVc9EVv7uO4T+z7BTR6d1
ytyzGnP72OeuArSEssFvOkOoAiGwcVp1Q3Vyx5Q3ZZCiOvmTOhuyh/uxutYgb8rLuuiTjCnCG158
nJEGf4XeAkdEQBnAb2UiGFHXTuhVHvvTvmS3Yu3RGecp7vhasix5lLGe6B0TIVsGPinWFOYr5dp7
svwTfclLA27MhbudaZSX7e/zUW45xScpEIeLady4mI8h8yrjh7Yz+W10jX+dgHCmeHuHsOICx2m5
k3zW8OIyNuxkVUXbYU0ehtKrdooS3nBMc70zr3Ije0EHlAib0452crny1Aos1Ck9aN2PfDVqGX/p
H6Wj9eT5g9OwBWxAqliOvBAK1ph+moyCnsjdwhT75I250hEzNRJc0phjr4muZaBHJAoe5o1PRldc
T0Z2cpQG60e3Lg0OLmcphLJPg/PMSc8rNvYpzqnJ8kuiH+G9q3Z9mBibgdf4CVsxQJyYAaCriM60
66Te3dvTz8oxWs14E6TMr9CxiCTl+1Rq/MABxBaMF3D0FABsKKVnAKhv04AijUsUSZ4NRg5zq6LT
lAkv7v6Mi3S/qONcQD12BwrK/hnodacouR5nCLdogfN6bFeWJ8Y+O7HZI5VpXQa1N7TJiNM+AtjD
oncgB8XdPNUJ9Mt4ya2DhiHOQlxu7wj1ot7Ld4zzSgxbOpE3phBeOVcZV2O2Ov2SDqQuQDn5fMw3
0NsQAQbzgPLsScWH19H7QoK/RPNIyVr5aJDXbJHca3GBf3bqeKo2SR8m9vMtttzhIz5QJ9zCeRPI
kI+RY1w8ofp4lAVoHVpe61LHVFmgx26A1qWaCaG9LRKkhZ0qL7aWgoB529DtYocLH/52g7ktLMD9
saRaXxnSOvexBJ+0dzJ+sE0enk2eaFliumPESsVx6bLGbLX3P9ZfAL1te+qtyVZQVQdWLvrb17G5
OaaLAOtnq4SIC6hQz0/93Mn4I/VLot3HbBygyBgrRVKVc3MDbWrAJd9lhL4sN80Zc3zja9E8f23p
EL/H5L1nD9i5BtYN4DmG5fFvGs1diWpBWOP3hXmr3vAYv5V0E9hAkirC4LiPeIUXyEPXVMeQH4Jx
ZZPQdCX49gXdT7EszETpOBI3CfoYqLQ3Eidkqjw2rr1+UhQG4GQjrf8cycg30sLAjf6lZSge0KnI
H/5b8fbMpFZQuTpO8fDqvowfS9ez229bUlbPdmvB/OOaoEpamzmWFre0/4/YfBrr1PHRo6tsb3Tl
bqnXuCs4MrCGecR34H3iLuN0cY8WyBDdTMIk1TOO3I5cV5bzNg7rcgNVhTnfXdELOaOi5FwjmRVA
IIZno6mLh+iA3Jn00Gi0kTmJOOs3kMr3E4NOJrvwcwjp7qDtYoj7pzxngGzOoBqy4rg/BI8K8ZVz
TJXLT+PbqPksNrexawY+sjaD1C3jd8PxhMjPEfrbBRmW63Mlq0gqWj0mQuCbgVmddLVGN/77KDvC
PN/NrVUFskIGWRaQjqLv9W2tC4OBqiQ3MOhx/lvBpcakzUG679iB8xq5ip+5fgFVpdGWRi7N8DLW
/BVm/RwhO6Bz9cNyaFBJL779xGXTYkTiZhaxZfPzhAoRR4FK5UQslVj6EAKL8KGyfFv4tJ/HVv7+
L3FWZULmGYg12IcOGv+vI9nLNW/JvbElE1cBGtfokb2EMHz+7NBfDcYtyTckUvZUQkp+CIErH8Rz
qC9pMYPJOk0nIPCCOsNEha/QeZo0bSDm+OF/2FdAquVMWGG7cx77cb3/EIs+4ag6ctcY3T/VZtMX
3MR8J/BHp6vwWkVn6kYvV9sCqbJhtPfu9+WOG8N7zN8wAxR19VaPphqpbhQTIx7kZ9ixNMd4533U
x++SpZMWMBo+/ezsJwkZl5/ajQyuy2DahBMxThjGDet7N/WNfbiqFOMl5HbCF/dOvQIJYFn4SZ4C
kdL+1agsXxxKH7Rsuq1PA+S3n/VZAwgs2Pwtd30MJ90V9wx4L0e7bAGPk6IZHnO2SU2hKIuM9Hk6
hAzYomgJTWwOqwbnuC0/5CoHK1lAhnL0cHDFaUO4G6sLtmLG8TYtH3bL9KN22x50RllljNJOzvxM
bLtEDNS4T/HfKyjKoiVjzbFaDsyLeFoaZpMtNA9KFgj4951A6oWbmnZP5Qo92XzEkjAXZfEkBkJd
YO9azSSCG9hUhVhe3D1O16WRv8HYyGwvP6/32zU2hFNTUOK/oC6Ytqa1UC1VQQbi9LeJCABkhEpo
f9/xVrxA9iNDFrQ3Hd/7x2AUkgCFLkU4gQeAHb9OFPdrnzZHu1w9kb16sEY/EPbxQMsJbFZWmJQA
gEpVIRQj+jvoEa85cwIdhI/A2J5a1Q4GpEXbOnxMWSuIL2Ng7SC79Upv4dQDCAfWZTbDteKAcE+i
jJGwKSE3eqs2OCYa8mHCr3F3nqRyVMTuMDqLhBwd3CXNrmBc005Yjub0j+wV+Q==
`protect end_protected

