`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
nwVS2CJXupErGPDoD8Ku4o1Zi+AYJi9tsbcPZPL/xRo6X8XC10paKNinYKLQl13EAkPXE6QL6ydM
lbzHjNTU2w==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
FkhL+cK0BtU+W+i3t7Ytk7Op0uCvIYyj8H/bRZnnNtxqo5u8IS/D9K5RShx7R7YRWNheaHMn6Ygv
fDj070P5zgsj8a1IJ5dI5LDna9WXkeMYzmuMalHydMJ1kudEmdOLJKq5WxEG1BRQsQ8k0lvVBfgM
yAAoO1x2DHNTgSLvZLM=

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
nLzdtZ3REDuTjhApuaykPnq3M52YDJo3801ryWYezzWQ1ygkRNQtz5E8uPdI0FLOp++xKvtemVgi
fpsd1/BGm2yq1zzsODcsA0zWeOEVUe7Kva8zwt3+QlNFRV985vvD4PADEGD+1Pg1mYbNGhKEz+Wr
J6fh1jXqY/tdPQg8ybk=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
SXLI3j9g38Qcx+QksDW8F+Y5+N+HgVxbkWGUtbeEa4XpHk0wAY4iMFbTv+HcN+rLS1JoEudk3H2C
21mMje1B3NXO8DeAIBW8MdVNYvUin4DNeufylRor7+Q9+T8l0TKYEjLntggmcDF9aBwMxPgXcYku
RdSlG0f0o+mSc4/alN4xOpAWw1p6czfQ7Bnq35E9wIclYfqCrWOKBuAljScCce4lHAkGi88+FzjK
g01jPDvOfPqK7J7gDmOV4VSR8BZsg4pBqTLQbnfmYGUwhsGr3Nj9GemdhadU5MmfYmDY3imY7ZeI
kPUIS3pjESpw9iA0OuTKr5fKJhJZ2cJ5CvwuzQ==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ftcg2N48NqCHefTwhpYrUPaMvMzpmuLqgqd3DtpYFLSd6DcixuBjwhWRln1WKGqWTyAm0n0iCabV
JiPhKbQAnTvEOylyW8uLjd6IH7B3qhSAy/BYI/1Bgnqd48An4sDXFIT9ou/WloM/6gVc+wY0BSk3
tSt3jTcfvZ5JIi1GjRXAUPYZjCQRrC1e1saS55grMZETTHa/hgk7xaDBhgmHlBHqrJeGKkNc7Tpj
OXQFfzDow7U3v49Kr2+5nFPJgGSKRUkg1X9xMzj2m0BoyzUNgYP7wZ92wQODUCegN8HM3JzCt4+V
1LvHyqIFm8cgkJZknu/d1XRyxL1tOTHlqvDQng==

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
UwEUSIba05kuRZ9C3VePFeG4phawLRcMXZ/OiI2pQEyda5H3pdyOO5c4P6VMWnOQK6zVjMlLJHME
a3HoxAS3EjReH2f/s9l+uJN1GOCXQFIX5mDFVCm9sBuDewxIsFZlz8PoKwVAXTjVVqKQJ7MZrTZv
CVU2unSpN7KHWfuHsfJJHMR7qoMfVxRHgpGUZmrnkbejh0Fx3rGZB53oWe81C0QkicrQDjK1MsQg
jug+MjAYVrdnlj07wJtTfleJYMiM6cBAjv8hDLe4hNRdVn8tG2btAMW12tt5GFrJEJqwWB7Ia7Eb
VxTM3bbsE2y8nRoy1mFThD95xJ9/8OzaVhSAAA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6704)
`protect data_block
Ex/npHjWRS8QPAlNeaCVNum0E7uwNWZ5gLPLfb0VHCuG2we2dOy8F2fomxoQ3cN/ftWSLe5X5UBJ
BjYlBiI9QoCyfurpE9nC/qcoIgB5dl6YxprwTtK0G4xk41xBL2vxFynYiQzWymnA2xz8f7R75hWJ
I7gvcKgyOEq14qE+jTLU2Qj3pcc9ucM3unUtCpZ+DNaCM7vr5ViBKefrQMQtGvkzNvKkDQBd4Nan
RmgaTb/y00kr/k5JQ/0odWxzCgKrM1Mnqc9D3EMOMuulxMm+exyutWYkAL64U2BW5+UaqnQo+rat
gS++wBklfHR2DLlOKE5WZT55uOUGxhqHG4AlyZK3tQxh6t0zFFGocaQdYrCY/2/zDdncfblfzf4e
6RsM04Xec0HKdf9xSWDvmamIFDbA/8CNS+ruAw0MPRXmzB5capDPuwGEDZQ/1godwf4Jg1zQd7hk
Y9qjC5nBQ7NfifyXFX/3ZroM/hBA1TT2HjOuMq/UdLMPFQGGMFQdZ/OVcmVhG6554vcWYMPtz6PF
SqizbO/eoFpG6pR2PC9bQ7jLOsbhPNnAjoiEYZn2k3+DrJ84mPTkdAtTX+PuG829IHvJCseBGlaT
QFT1du+crY/WhHDXzMBGeuu2+zFT/ZKc1zHYxHn+NGIyZOztV8CGacIYe05KGD1P7MFGbHaa8D7/
OTdOR3T4FROb7kWUW5D5AT1qPEmdwS7nhvljKx3YdoGDnIqHHJxQ8thehNUk4TbH2QIeoMfEv+Bl
CNJcy75heOi1r+3RVaUGV6bYovZ0H1kT7np7b/vtmNC1diXo5DcIt11T1ePAzMfRncU/faUSQekP
JHuPLaa7rQhOkR3ou0GB2MClGmN/vRDbP/NJkcd0+c4USf9VQf/huuKUNYGnLn8ig5x00wmcEml9
c4jHN++9m+1TlyeHUhVXat78/0UdxxcgAWJN+yIVPVHbWOWHOm5Bo49oQOm662N1tZq/FTJOrwax
p/lDCUUNtBobLJrJWtqyqKm6D4MJadWZem+HhIDQOm0ivej7fT8sN7gmkcAYhVBKQybAs4a8sBkH
ci6ZUyiuY6erIAja0cWuA7YNB6Cx+neQi7E7KgfR8COnNVUCI8tjzmcWNgZJ3ZC7DjmtzaQ+xNO+
XMcwdy80LDRiwPinMaes0uHy64cm3Ifq4jwlQPOWVaCjDceV/cJyErm/hY8Y1dFWNyfWWEPrpUP5
as+cpmlIsBh2GOATCAnlxYJrYFeXNCaPlCtfnouW6FXM87HYgpCS4UP4XqCEMpgn/jlAt5jFByiS
L2VQG7DSHVww4Sa53QfYEaZ3n5Dnn8hm94TF9FHUlnmOr2W+CxEejaAi4/uuTds7l/5NpAqBcl9Q
X5824bJngYzoXiVmnADzWbxsMUsauo9pwQSlsQADt4OLq93ZWC9MPOhY5UWWZs98634+sOWxd8Bx
OGKQ35ubZPgIKNikqgiXh1Vuiv6PRcPfQ8OMhStTzJoXvO1u8n7jobhUynLkbBY+q5bJjlyeqYbB
1krc3sulHNHiEHY7HiUbJjvCM37xjjx5JhEx2VYGumPne3s/lhaf4DnHtinG634NfiWipQzNvJhY
n1LqdbccW36tKsAwRzqNAQcIjCW1CLxEoWLxkX6vKseVPZTkJRLP8Sw3jhe5HXhEeiLTHT1DFErE
GSrhpigFQMoub3aV+4ie0yE4SIP3vW10eYKYsfRayMq/T71lIddEYIRi0JaQLCGkIJGrW18vJDO7
SCs7kqcKumXANgn66uGRP1+WtYcOgk5f6cN4IkZr77fKbZlqDD6lzimrOMOz2V3qHIfxwEFSkxZ2
7cbFKLzPT2igGsy3WHlvEiQt1d4oeZ7NK4AeTTlz3x6g5oXg3qJ4ClupNiVw7f//zL02zQ9e8xkd
LF6KtRXbcTgisBj8LSifL6LREW3BBsQg+d50IrdxmxtSb4w41yFj5gu6yUvmfOtv82/fNl6up5JY
8AWI8ckr672ksJxt4rApsOXhYuD3HHwrl9dOXk0uKBgMsAyy0dyOW6sN/3STdydT6NyCQFX6Nnfq
GNhuwi2DuPj2EbQjZRhsNJperV05Z1zfpqYG1FQYO4VqbM6aDvJNdBmx7AGQcHMbqDuPmLcfmu9L
CkoBym17trJEt+4qPN+RPM07hsXHZc0HxhWuP/wT4bz8miJsk90MegEbHE4X/kd6WW3LDyWqNZfK
GEgQ9oPwlkXpyEW2lGpU2Q/w/zUO14ohCVnzw6dKnp+OvSjmXAD5rWSCse2zVykcQWAEwXYGmOOM
qV4rlfFPB00yvDcipC8A6bbsCmrmyl+9x7p+rCv3gLNAe1ROkzVRNgajjE/G2KCMFpwSjdbojimg
S2uYk24q0+S82ysntRT0EOVIk38InEZUKLIYtbmvrzugWQ21XvYAnaHENplsTXMcxnNSmlP4l0zX
uwYZkucM8gCbnKzRQ+DVNJnhCLH8kgs1ovmtHExvDa96zoBr8J3SZ/nXXnoTOwkFf1CTpEPGhtid
WaCnaKKLcy66mZk6aKcbxFAs8BSkg5eIzVNL4f5IdPSwcDtc24pVuHGrz3EHkMt19+nXyspgJKo5
elrF3mVqq9JaGuf2AJZZHureqa+VE4w58ZoVY2pebrvBnn2VGiNHihYopEKQ4VxTn+urI62j5hI9
KK2Xl47DU5Yy/YGErGhQsJHtUAwGBd54vNi/i/6MqmdtNZJGnmxPsrMBuotRIvNcqKMLiONKO0EH
KPFuKIEbH7ssC7p9vdXi7qIhcZD65q4+DYijXH9GSAz1rctxiXpWpKtNcXl0TmtfmR0UZMyp+l+H
PLb47JOgutNoq3nWcBMCQpJIbt+XBjYJppn+3Z9Ox6izqKnW7j4SV5AnCYv0UjDSwF2cUj7qX2NX
YcVGdqME6tEDxv80uGN8F0gVqmRZidVv/J0ljmVHaiSCyKcydP6MyrrwyKEYG/IE/wf+QK1y/6y3
irDKi29G7A1gS8z1vfEQAwP9E7YNGFut4RxeenMIya5FlxbIXGb7Uuo4Lkg0mesjDK6A1ZwLWM52
1ZC+eByOFCRDxJgy1tNM6efX5TvDCUcSPmRMMTlpR5VSvtMoJDr33Xm8wjPUu5hRlBbz68zb4cXc
hEw63LbNLooM4MIQlY7zfyv2iAiM+x674AB6yMrFU2wI6/xQcQA6Wp2K3dMdFTX7Lh3Vg/DbJEaR
srJNHr5M0K7gCLooTsDqppsmNNb+j6GASt05y32Zp2YBHb0mnNnRcCNlP2hirK7NfT+W8EKuhuCy
HwomWaNaUFVS0IqdsIoS0o+WJVMOiuestwefNoLJKf5L2WWmYidydLljL5kDSeZGY5kl74pxDCgm
FjLC22pVl8ENG1tG9BwyvJ0wkOzN+WdUgVBj/5KKO0oYBQ7R0rZL5YYpZMt/Exu+GhWcPs/YUupf
AMIi4LbihMnqx9BbpTIDBTj3tb8TAq5lMBkALAN1xYDFFtJ8QBrk8bK+ztHuV50YEQEuusVrys1J
TbraWuhRvAd/Z8c27pOJQk9fNaYhKpkhBQK0XqhelOqTiz8K/SVAuSdpYdSGw6PE/TXot99dAH12
mqMGexBZ7a8c/TdLEsYYWsi/WHfTP2z0vJ8nI+ISsCJ57JmW47rMl8T5AQaXky8aPFq/Tz55uAh3
ojeZuCbPUVoybMm+4+DrihIMYwyUwWfvxAgtxVKDETpue1pW1UEExqHrp0HWPDNagJJS4NGXTPHd
7UTyZlTttWY59x3iGjYOfZu/XBJGEpG85Hz99747b6Mq+WcsVDVAmHsRTxFF9OQqeJrC27z7VAz2
rhRoSV1JUUKnVFfjc6aU1GW5ZxVo3EvrG3yRYHkZc1o4N1+7t9kcnXwYUxUMMLXJ5ifkdjFwkKgC
6E76TIzQXIbKgWBn9Ve58M77wTi8ffzcNi7kUzBMoqj6zpS4UhsUGM8iAnfmX45Ke9R21/OmKyQ2
FcHPUvaUno+pL54cd4iN6F1f8q1e2JWsbBZHcM7UvXVSaFUBb+Beh0l26ysdtHOZFvgOFYBjNEmy
OT94Yr6MpHFoYjy/XNnjyvvdr2O6s5CSLYSWCemDxWXlnW8QsviPx5VgkIpxWYz/xapWX2Bf9KuU
yCTrru6GIgmqIzlOpgD58Rab5c5E83C84Nesk4VC2bzMRaq4nzfG7Xf9/fFDpUweYNuigAfPWpMG
T4oTlrt7fbOO/lDkhFXSB7lUd5rDK9WZHEd2GQOWolGNRtBz8zYtJKIIAcwlB02ilyPaE/ocov/o
/xFxO9SizPQRp2V5DR+XDkzJNvktcgBLrb/8q4PBTi5JUZJA8dMqbD1Njr5dPIG3WtSqjxZIF3Ue
fTlU61uGg98C2i/EYfgJKLsFD37kr1+BaQ3FebQ3TvkhO3L4TYmRL1u6A9Ib3D1WfnCnm8Ux+hdZ
JFdjx0AjagRR9qwZI9nDLfBssv7Iaedzb7yELaWwVaaAQ+2c/MiN3B26NWldutpL2d2gDpv6ak1i
7UFBHiiO1chKZ1PEkJ7cIUAiJum90fbczuJ2ZmixYzv8Jks9yIr9cHDCvbe/uws2IYFM7Pks30lz
kZY6YFHWDUz5btJbi7fUqHVNsJkz7hebRxnKadNXL6Q6w+qdJcnSPzW+WXxjBaWK+outl165jvgw
SSZzDViOtxrBn8Bwk5EuhrD0e3rjg8JgnEE2EWESm6/3cAKYRv8v6SI1xBtBSov9+itbdw3p4Sgc
bgi7heYOBNP7S/yfUCdtEGIqi0/hjeCXJ+KgccqJWrTyaCZniayKutw9/8gQYjjsL/Z4aJC62/aj
g41e/tNcpg5lfyz+CELNNQWI5S8+UtutSXm0q0QlbkNAPZdYW6QD8Fg3VUxP0a/VuWC26xxEo+WD
O12amYJkLkNmDKyqMWYDta7a7RRTGHQ3U49BKyv7QISzKTQPYx3pwf5DHnhmRjR4BnnMKKsEc+NZ
9IEE13lfJBapwvYKCY5SkXN1HvL+foa3D6s2c4OtkOUn92zQCqDkm0TkMv18mvP+xcQzje7u+A6q
iyJn8H/xyHYH+4D/NhGwSIQLKE96QYIy2V6rlNnLE1b3/bMLoNHQtxOt7e8ngx5hpVPMZM0dJ+ZN
GQ6VM53PgcFhoWHFu7g6OLrdG47v/fokhA5FXUlSMZLc3mHDYEcNHyDHwOO0d0DrahpuYBary5p4
r8as6iWDPLKpVn22ejn0aZds5ilz8ZcqOAPsq0Z/7ZI4/eHdvETLplGUzyOqovYnyJK14paBprIQ
yMIzkyHRm9WOpA2HFjlBnATH9CN/RIvfK3UhA+MXZ03OE2/ERHy7TwAAjEGlM4u8jH+9O54O+xr4
mzyVTMUauPTGwY1AjD0ZYEtN2gfKOYQ1cCu1HS+GJ4qrnohuSdDU8HU5Y3NmP+x/xLXC7MCLGE9g
WhwDEm0vV4DlNIM8VpMvnXxJBIdTE15eqUmAfLH1HE7+jyFIA/4aARDVMZIz6D8daB7bB75Grnmy
tvzL0zpBYCrDOKlNq2U24AShvpbe4cNLwZQBaAO+DcHRvFQcu713m2ApUkZiDcMKdEyGfvEE37BN
HdQ+2XjWTZN910lht/EeiEiVpCrqteOm+FNC7eIgyNtMd/OIKgfSzYcnDyXTIUtYMiMONX1uSuC+
THnHMyXiZH7wvMgj+ER1lVqp6PJ5EXRxC4jD3vLbZRjYkmqbFyaNIVj8owjHC8nzS22P1Ddu1yxb
Gp3w6YcGH8jBRONBuzdlKhTI35xY7PXj3xaI0psn6jsApWYk1MZyXr0Up11CJy0lKsVRZ3A6YZdq
GwGii8I4eUx1XdYpzy7WKHSyCWg0BPI3j5jxvook7ADIqCLENplepFmvS19xbTqygvA8uVB/Pj7T
zSIMYS6nsh2tSRD/iTtOnstsxsyH5FxxGURUIGT/ojzfRN8G0qzghHVusTHMQlZHv1b4jt3bSAAk
cHaDMB56yc5vBb9+M8omli9susF1oyyoS0dr5XpzA9cIZ6TprxpdNOFhFvP+M5Gb4lLe89HzZCtF
vUGLs0HmLJn/CpZkPxA/TxknX9gVVKzi/D8OaboUmwPsfD8a+f0/5OZmfnwTc7MVJPu+y+IiP/Zb
VBlYj/5lZoRoTwGp9OoA2wywhZ/I9YN2vkd+sS0h8L8dC4Niw0aM7dh2mOQzGi9fUNhs8udmBVFl
Xqt43N8xi/Y/yVvhmtOCzNgh0BsvofsqBwcUzBWdVfqtidv4Uw5Q6y0FVQZjhtSiyXK/nGe+L4rb
HdWp1w8OSZDBd6EePk5n54Ws9FmIENMaaFEbLLO8De5hK2WENlbWmdANDWbU7UBk2O6VQlxevpJZ
Kjrhr5NIkx87gPoMXrl/p31h5DjLyZ2AtSdrYb678XVAJDFtyXDs7AiY+PBCD5OkH+7iLtHEIUdF
sSNhntgPIJ5ZgWj8yKYxt+yKMCzUVVEOCoEkdFAJG7C25VOOrVvOnfFFbrJt5X5T7Q8vsnpnI3tY
aXb+eOyogt8RhnFarvwyKt/lYzM3/NV/IzaPHO2zn+qHtuybN1e6hGoe1Gh5K8a0EknQc9TZJc2Z
O7OJvFiDCZJQ63hAOhezznRQTitXle+GLDg8Lrbp0J3nc9vXx9W2Eo7FtVj8MfDyYzs+NU3iRF6l
V7KnXHURRBuTmyAdPQh8JHaC2JZ0HX3KYcfAeCjDgT7NObK5rx/TCw4LmUAZ/9AfKLg12cmxVhws
0F9WkBANIcpu4XOtR0HvC79KtK57tgV2XQ9nbwR4uX0K9X+eqkgaLAFL8QR+CkhEKvnIJ/SGGs01
Qwy0+BEwek1+NCJmMJcSl8otwBZbblAo2dkL1MemDnWiL92hGVZlMSYBEFjXpumI2WvOu0i5KFw2
xrs1/RC+2EzHApt+4EOUzrkXh5VB8Lwk2djEnU/WIGdYf+xv4/5xp9lr0dRufpRTR/qzKdiTDIhP
sMbIsDdu3ihiDNKIe9gOUZzQIgqhM8tK+ssPOXfW1nJ9XiTO1ZVkTITnSj+35eLUuYAQh5HUqYGq
/eOh+c9y9gJoU9GPtGzwXHPRyRiIov2igXUABMj3J0S6sD/U0LH1nfiCrZ7LtdfwztYEyiIIsT5F
IHO1DUOHL728kiwqKgV8J/It3JBoSdegAkR8uidJcoZHhxyGYItJQrPfDLvJS7/9zgIYwozzd89z
pqKEgbPCIUAEY8D8jjfpq0QyODJPCMBrAkSKeW1BVae2rz9T2ayQrwjNO5R4zaKlZE0xn1IcnGe1
Kwy/lSCau8fz2/13odNmAupJlNZcKs8XDHqe1Wdiv4ltHXryxwroB70w5yPHntk96Qa+EbRQpDBt
LNUbiM4wL37s9/4g/rcLys45f0SU+cqkbFWxbutjJtZgtVxZxiNm/g6+/HlsbzO2pbR0kRZd7ftD
J92PdoepBbbMmn4qyJIEk7z6JcDpOmP5zh2z8k14xqm/DXyJWG6jaDNlPZU298EVkjUc8C/y/kde
PsW8swa0SNPudCVBnN5FRmBJG9xQUujPIGiak8SufkKq1y1HW7VrvhJM0BaQQCXPsJDsV/JbM7ks
e+RGUnaSlB+pLF2JZ9zIAKESz1pxZXiTfRoQ0wLqxJXM86GY4Kv9yWKKIqdLcsZ2JZfpkY+Fzest
fHCUeKIy7DWR9f5zWdUiKgB/hb9fmJrfoTKUv4ARnsZfl0ZWAE1RmZu+4K647AOtYLRHqGjh+VdL
9krV//w8TbZtLufEez1GBI1kNU2JWPDnlBO7YRxZd4VvWsFuM1i0kX8KyFbGO+7ZL3GVd9sU3b4i
c/OxGI6VHtcEtbCfp2Gn1PYrkn+I9oWYh7R+YTzwHFyWAOLdimEiw8f88bj4cF71p3lWFmh3S5BD
dlmnriNI74Tu8Xm8BlNTFQPt9kL6t1QO/jgQbgxEG9a+So201jEgVrSaN9cQ8U79qNPPr8R3MwAd
unkOIHKtcoT9RscNAMv6XYz9ftFtOHRPNtZ6Iry4nArLYMVXhnGngLkp44+ZFz3fHdRe1ef7I7EN
QD9ow3Ym4LeLm8cRx5VOFvyBAtGlBHfSCbguubm/iuHi4AbI1o0/SvZdoxi93Pq+ReNKfn57m19J
fSzwB5YRXqwswZpNgPhyhcYmv+YkqkRpbmnXEl2ZUtdiGNaRPut6OZJasExaLTtkQSaTCyhKqezd
8W2zrWRrS33RwsGGxNYYTpWpXcGMJPyGkrl34o8yHZTf9DY+AJr3bbkCwwY0jYtKKWmhWWTpCk+L
bNFI7IzgTjhat9T7ZLn+/5Fd5Fq0ukF7lKv/gL4hCxkkLi7ASH5biTG/NgbbK58P6RTievTFImIO
ZEPBeS+F01l50zM3Tke5zSRM+PlUOmtDpu7Wlld4e/RnjfMVVprMzdoEMDILKmOv9ymK/GTHYuKx
XOS4d1jDehUsTQMo7UlzFnFj/DUjcUN0WvQmWotZgg34RcpbVy6Kt9fgW0r9qq0NOzA3f2Ly/mA4
4mYeAH8bL9skFMtlw4jlR3kP9IMxnjYzOx2CG+lKJrMXUhDsrEnX6oPbnzCobCOLbCKz6QuIDuXS
aXah0YbnoGriuZBODOQSOZNT0BQBQEx519caSXF82TKIe0OuGhgHqIHQ8zWE7vpOaizAV0dc+0SL
baUtDU6j4RMs4aZXV7rMv+Fm28P4uoByD6otNy1fESD0sikXByNrHGqJHhyp77RxTTnWtD9xHM0a
aDim0dfKFPFYuA5bWl7LcJCgVdjAQq98Kg9WcSLxHxL6GkTgbZAJo8XENCF2I5g/su3tM8UxU5Fg
x8xQpMB3wGtSMBSTO43M9LW3XHMa0Ze94p6/0ilqt1hpH6nU4cIoYxvJLyFtuO7vvReidXDwHssv
iSQHTJaj41cOYY20tgGQVigrsZK1vcZfVkQhvXvBchrG2nYfi9d189vuioyc9sUu5d+H8CdFVJL/
C9DN64+8f5J91pnnjHQrXJfIfUUK+3xAxOfxveaDpZ31TY8=
`protect end_protected
