

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
DNkSCrKrSZZGZ7V5MEC0Sa+FIa8Gkzj+o/6NpxIyEzT1r0pebmEX5gzn4ZglnkddvJ8/1f149Df6
ndMlnzvmbA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
W3TEk2OoVAEcY9sACr8qvdTXcz4KMrr0wBUYfTJiYRXEKj2r9L+Frj5vlPoRfXyR8BXMuNIvntP/
hRtRCfRyewmxrXe1oHJIEkJM8D6eCjNM+zuIptS0mt/AsnOv+MMQLDkTVqLaJNUJXubQtL+dhzzd
RD9SIj/ZMKv/oOZJjHU=


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
2wWKJdgoqz3pSafJq9a67M/dd2FxPncTZHCUPF6InCTgFQ7MOQlzLhplRl102JxCos5KzhVt25al
HkjLSxu9PHw1ru871OGKgua1sS3EafdVjGCdT5iL+6+M9XT4bQzC8cVlky4YWr6qOy3G0Bl3zGGA
4U8j4LRDtMi3U1kOYa0=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Kxq1/5UngNEJdxzilglpkl2MQX9t6W7lRQYEeATFLTlsFzdBmcbPaM4E6/H6jb3hTjltHCzXXzJL
yu68g88g81H7vk+zIgG9p+bAH5mVTWnGpTcQ9Nq3V+BFNfatOquArwL5wvfxgYh4qmnz5LLzO8Vn
ZipCR6RyJHvmX3LECK4ZGhdOjgqLTbHPcqhN/bNhl+BKCVrOY8qTWY6WSJt2I/pR5hbR+Gxpp0v1
fzycz6IA1AnyF4dzdl4sorgs97DN/Rwyy5DX+iGMZoJWJSj+jKc0DU3coqqjuApwjmgaPZEOIkHt
fmd8I93zHpUVO+LU0o2VXdLy/rhhX4k5zyqLIQ==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
MMro34sbMT/dSBUUDKeWGj+AS/ioQgVbGWAXG3XMUY+tNHQekxt+oKRBWcwquBl3sw3SJLbR1Rnx
TjJ2MDDzEH5uCz1vX7jZaQbMCFAU3K7MBn40b87mRKYgK2nBkQ63tKhSjfklMsYEEkc5/qUdspSU
GIdrS3bVjN2jI60HeE4r8Ae7725zNCxoNO7hmmiicY8i9qwR3Jx3RLeEISc/SwYIBg0patrQcspa
o2nUblqCyHtuSc/DkaBV68tb1S3LDYROKbnkmBVtPajoK0FwTW/5ES6DuetOb0ujYKX5ZJWNoJr0
DsAiVxbKY23jSFr7uskYGQGx1K/crFks1SMEuQ==


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
DXzksdzpRyBvPJAO8RW4ZhlhoWO1yMLSwz3BzpxXSQKUFJz2DfYgIojvnKP+h4SEWOeOMQNr+agZ
sZh5CyJzK3n38AYVr+qSmIrSxy//25NZBDMRWM06jl3lxtySkqX1u9lRJvnZzDG3hVY4BI+zv+3m
Uys3/UlD6y6GV0iCZqSqOjNMRk77t+OnDh3CxzRxxv1qIqIA3AkY4LV1fP5qMWjFIYo2yfPwXZ31
leLLHOibckzEYHfpK61VUGsfYsK/Omf6e+sJIk4DfwW7z+qr59Fv/xjUYitqPxa99lpT0eMUcAbZ
NbV6OJqwWXo35ZdTdYOXEUb32x+tBF6ayvy+zg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10944)
`protect data_block
6U0SfWmc9tql6Mq4Hk31tAzaaPbY45ugwT2Pach75vxDHTmR3G2QVaMKt0ed/TtgLD4wsGow9GRV
IjEMaxnXFhXGzxWw5Hrvyr+qztfe8cH3vA5DaVGglTrrRax1rJzUVyccKNHmUOFTNCrTYGDC+55/
P9/ROfMPBwQEN+TrOWFq75wid5o1zfToI7VsbEXf4R5onsMs12kaShL4KSO46teG/iahE+WlLvXP
t6CwhT/blY8D4UmlTu2xI7LB3bqLNAbVfPzDOnMi2hkQs+FUCCs+pSaF73QaU6RnBNMTuNoeuxR6
2y42Vto1CFs6J0iakB9yq77mVtPRbSjEOVnmGaKMhMSUGLG7JRA58gsDWXZCLVxxnKAITXdSYKKn
39FLkRvRInFXNHdU4/jC/BDGNO4CYBRecRl4Oc0XNn+NX+wxQvws5bWLNaaJiSrvGZJH64KZiK9K
4ctTuBL4kgCADTUoYVYecJs3yAzFmY9gJ7AgfAcriXmwbGPDAx0BGdWoSyd/Uhe4fh082RutdYUi
BMizkLyaBGwdXaE4nr6C5OllNJhQHcVy6PAptYujd6MkqrmX+W0HorGbeumbVUBLlCUu4j2X7mNK
K49AGGVLyxx9xnBLb3+HZUfJdHbIdQpanTmZU1EAgLirtbOPU4NgELRi3lon/nUM9CWBTEPNv7m1
qVpsGokOQDD9c7tS7uqc2+kKbONRmlreTDgg3DEIfwjAFfz41n9jajS2s43G9kO7q6bINimkDSJ5
n8SrVbVtY1Mf8NNmipX07r0PTty7Yx+TDe2uZoquyKcyhOXk/JKDJxVg+inIyLZCEwCZyyQQNqln
OexZmXb4g+ZpippgAODJufTyHZf3weB48R8p9Q5awPfhtMIuG+GG3SWOHQO6okVZnZc2lA3a/Leq
0qZhRb3s1ZowlMOYJwXf5zbkioNY4X0HTZjjpTaplRJqFlHcPD68k9Mlk1AyuAa1B0lHLH2IchxK
FzgXNNO1YbM3VDWckd9iyB6gYN0ExcdFOxUNX7yBbtENzrb1Y3k8vbD0AH//qjwKMDmvZrzX2/3J
Mkza/2ZpMcQ/KPnmf6k/pvhxjoUBMCyzl41MJDe2xCajLucTos6pUQ3H+FMkJU7nTYAj7ugytyO9
bLqUu5/ipHCowUX0wSPlzcKwEru9CJNqDF3qKxvAZW4zMGRkA2ADoW7hNaeM1kkFlOwEZqyImzcc
h6DjKTrqTIQTFlazsAxqMinpaoF0mAu/P1zUInZQsRlB3I87R6COYqnLGikEe1G7GmPNxy1Ytmaw
N8Nvj8gv1q3z3Qd35dGYqxx+Dke2HXTQnn5kiC10HhVSgCN5404tJqUkXpOQk5irc5oN75CKFZyY
/zFqP5M0PzR+f4pdQl2fnboU+cdVRlX6CHnAFkagUz26GApRuU7TpFN/fZGbL5Gq4z9sRG6a1AUt
wyCSInLmyk4F6zRiBGT5hEQtX78pq/mQStCJJeJXoJ2mBlMkRLMpK5O33t7t2b/v1E6/mrzK6nOZ
ljJt8li690j4KokUvlfaxLKPgMzULaFRBD8mMzPfDBx6vLuP/NzR+Bp9W9PovAmRAPjdCWJm04mm
GwNDHYEu+tLVcpXniNf9EejT6LLCajZj8KE/tA3dnzBrMbRCBWbdW0BhqZ33aOcgkUnS68dm+jN+
bd1k6wuR9HCqeI4wOwrBN46C6rHGb1i3JNJHz0zKjFBID8NW2m8zrXvg50tTDNdNLlGxS4h7pPW1
TK35RsadHeis5b8Pg6c9iXkQdSgHxH0cq5qxyVJsRRIvYWsXjl87TpzJeG96w9oHJOw8udPR1v8i
U2gD8/Agko2ETyTxYLXgaBDdIpfTcKDAS9w/40JESEJvNtY2bUq06EFNQERddvghBwb3GM5geKjX
iAHtlvTgLKLETwO+fpIPp5xSh5sUv71f+SOcKQ8CoKhKYneEHmn5xFRvq78W0CcXTs9fMllpfxle
+NMoKGJlVWZAVj/hTPy1YL6y6ARSI+mF7i8YQ30speRAC4c/oR6YY+iyYly7MpX2tsPRpxTNhHkY
QcrHMXWUPKyhVSg/NQD8V9sHhX4+5hoWL70MtaSdWOqpPhovkgXWBwoS2LMdaGOS5e0ZZtX43ZdK
qvfWh2ejGB+fRTXJiOptH8hOA9sF9IsxcA7QPZW0pQD+Ez4YbGqzKSIyALnUiUXp6SYpIPf79DOT
lJC5PXNuIIOuj8iqeCnhtA2GvFHZl5jZvQcHjugcZZ82WY4p5lWRMKfvaCZl4O/K++DkXCvDibG/
igHdR9Pj2pJYyCqlLbFjtQpz+4/+gBQKD+9fcDWaCfEPp0R0/ETS+eUaQFNs3XxE/8S0YOPxckwh
d1cbHbIJYvppvgTgA0EbMtM9/9As3kg78ni7mwj9WSgeiIKnlpga3j6FextNKBwF1iXB68261q21
34+n/0v2g5/44nQ7YSx9CaagVE3CWlonYiNOjVuQX/WhgAfx0PpddikPDJKi80O41iKB+QbAt7n0
zCid7BTwlolT+YsTWbkJAkUW6RwC28c1wffK5/SiEGatCPp7xxPdtWkplFjm1v0/5+K/5kzlUdau
DmfFIhDzqas9wwWfAqNsylL/1e+cAh3hPq+sPaXDr+4NEUIjUQyUGRH16CbkUFEUAGiYX3Hi2Ipx
ysDvcDHADh7+l26Zyok3CKWNoIXdwJNH3GQLXuW/FmFo9o1Pghg4rUdZbrArw4dQuWlZM0thxzok
qVQswUo0d6Rdjh5E0e/mqQTJZjQSsRvXAhrLnK+/7/bBcwBiARyveod59KVDcvWZhmVCNTVutbel
42hzqtE3HIweAbMcNKmGNbKYekL34ifGm4GJvaZi7dB5y8kuiUXHh46RDoEvNJPnCn5uR8tw0CcE
GO81u0mr/XGor5ajbWqpOmcF39WT3hDjMbb5cQVjI74wZTZ7JLnREo/ee7vnUumCChlxKXeCSNCH
09ERHSRF9586M1t7xzkpBj6eQPUXA1ABGcAbhA6QtUakOuoqEWge+7m3VcN7/WhntgEFYlDiy5pK
D0nX8y498dMREHnSyA+eMSZ9oiIbKfickr/1C9z0Hw9Pgo8uXcXxySoEZU8WLl4Sjzn/QRdR6gWi
Fvwm5ORx35RUwJgArY5FwiCQqxJu2Xk1oZm5BwgPzLqEl4poDtZcL2zD2KPE1vBh73wZbhZyEgRC
zCywvEao1NVsyrr+WnMvxydU8WTkuhYiCuCyabu+y1bfIXx4MUne8Bb0a4UJrNFALtUXKnHjhEHX
Inryk7vyGxvOo2WeHKcUj+MgiXY2aRB9QKBELNx1HpEL2jhDGXYPHobNlXEPI8yff5HhWUqKQiqv
iTR8HpmSq8qcMXuFxBzaOo+V6owoXcs3QgOK2WbIwNhZwsDCC5GHKeHU0/UZrRm1oINEq7I/Kdrc
ZSooD4rw66Z8IRCK1scLV8BrZ1VvryfMq+4atesX7RKDsT8y/cVC8VvaFdQhINnIonBECcH7jLR9
DEK6faUlRTh0s6a5B+JmsTxJix81G/bPqigsuZg8ztW+GwEKTHxqoClBBkKtyftt6aAYclUV+nLQ
sBxN6a1qrm+Riz5F6y8cExFhcinv5Mpvtu25FtAChMk50xANXq6NrrTPbmGsN6FUdPXmWg3NnWdU
/5DUWZl+thAcx0ZTvQW8XId8b471J/plixzs3+Hc0XxeN3KGHG8E2ovZQbAB59a4AP0jKviJLSAY
l4pzihS5maxLC+V0tpdWJhDCGw+04henUAGTbkmWGvK30hOabZGVApWeRtBKAVE881IUYs3b63OR
H0fnFv3DNATlyGRlYpVMTnMRqAjt1BLKY08qZD2HygpdnHozypDWOavjY7Gyitp6GRb8bg4nCK5h
ip8491Tnkl3GiFJZTKa2cGMcg3xkA9bYohR+1gwijJLQEnVvStgneEp6DKrDponIE/MadbrIqMrI
AK/swEuwdTgezHIPoceE8OggXlB8pMkznTifZi7/q4co879NxeyxUukfCz4pbWXTIvSETA0r8qyj
XvLeGnIPLDT2Y1ybpDKwDFkJl9JKXEU58fls155LyhH4jq//nh/w2DJgQiF/dtdxWou6A8nlrrb3
WHYvzP87n+I/LoMi49crSHyAPgad/VOg3bScZT14ZL+mOWZAAip0OO3P6y+0vj5sU2RHP8WPMmz0
b6Jqxiv3UJN/HbvfkwSr46WHSdXjEA2adkHN6KI0caqORdFQx9qHFXFckncnYHUc2PeYIUAh8W5h
FvwAFuaxcLMnM7QRpWs3+lhe6jnVPltClFLewTOUz7y+mVLf6gicnMHcRLNtmXkwhlfWDzOBrnCt
4vcaztzIkEKCyYo9R+ggzeb+i7aF0wZOo8wlxNcz/iK5KLHXxLv4jexxqPZ+M4u5SgQNqRfFEZbl
70jmghZ4N3snSGolZ67ngw1fKGhsJpfzap2Z0MrJyNNQoewmzB+DlyUgW4qjOe+VXX/BDWWLpNul
VYOXITtfnS6K56XelqhXkRPAn3MHzqXckLr+1Ynqbq48IfhuCdm3LfmLYhcpkPM8TZjFS5b7PudK
BIvTCKfME5vNkbEA+jIaxBzyPuvOeiVIZciPAY2Pe9O7rszl4d9n8G5LGnDkA+ZwQEE7hmnzI06V
cHuenOVsiLXeWridrZ9aMzzipWEJmvB5KlzTI3q4rGVZbv8m+TMhubEvULvwJcpfSSFx7eJDwmrA
rnXtXmgSZkn4tkJJ9TBp3Icv/pEPNZleo88Xl7MnRH7frWg2acahnEychlRTqxIQ5zIejtjjHF6E
n/1uTNb9R5nP2B2oQxsUopEwnkCIJ55Y0YmxK5hzY1KpDi/0ahpg5ZAD6vTnxsqyB9Qor+xa3M3I
LgsZfBYROiJsyLFHh0bF+Yzbj0gLJERAi9xG7HY7S4/j9Pj2Uf7gfEi9kMz/5GkaoWoJGYZcm3sd
rX+AApeS950uNS/gSp84KmL18gQbiCb5a63nzUiO5lhanZe2QNhnTe8dJznaPJHoyCFx1Qr3FlAs
Q021tKlc4QTu1/5XrFtKWgu89f4ckopHajSKmCxFou629OK1kKHNlhzEFskUL5RBkyvur+w/PzlT
79K4ZK1RCU6Gwb43p20BLwKeP7dlSct+DOO8uQGv81ChaHtDPbC20bW14r2vI14z+xfgwJpzzcRH
yg276++U3DctYgyAkP1rz0rX/s/35zC7PGVWX9ocaKqyuoiV7Rr/fgidMsF9ySjPN9wNIstd1sGJ
3m599USMg8PUbdK0nUePo3rn9AHFurpiPXaPnUjkpGuOnHiAFlyeGDOwEjqCs6JoPIDj39NCU9tj
fDR6NQepP1Ycg+reZvVXELd3D7F13cPXjq7m8cYmBfMLNePS61a0yJEN92Vnnd0ZwKfD2tO2CqJj
JjNs4SSHZq9rukO8mWCPT3zi1+Ulp6Bf5s/bXo6Zmu5CWH8OEJSgr3Vl7dkear4z44JM3IDzKJ2T
mc9UcFv/E2tLJ4aILB0dH/H/ZAZc/eudMXK4t5hOn2SNA2wdmDfKh/hKdxXNSp+4FJw6NerBt8dN
2s36lRjzc7tWGfZN5gsYDItbfQx/L8OY9lE0KgjeIxqehVyePkNg1bynp2H4o05/CMCfrDBeqJG4
9szaVJwQrUgsQ/vcz26lC0oLVjY2gTPZ2PCaHooqgmAj6eHyqlw/SoN8dgA0bbh2tprPQIlvXU88
x3LsB01MB2DV0dB057NOY8iGRR2czQyQ3ERaTToKAPZqGt32TZ7qvb/bV1C8Vzhm98Ju+zC08tao
WQvr68vRZVk+JjrhK+LZ1oBriiWHxWYmhbjIZIBRsqMioURV9mIk7lBS0CbkAdseXsFEAZf0bji9
W8zpk3QFO7LE3/SYfDVO6FwEP5TVRHR7kQw8JL1nV80BGi2BawcAE7fxTQAmJpZQvYcJYmprDR7J
iL/383FLDjeB5rxCE8NrfDdCn3+mTxHOywWbTrZxJ7HS/RezZhTIhdwC9w8yOdHRXZHjGOcwdytX
KDmZyRWkh1vHV50RTlnzOVEajYx3qCpZEe3UhjxFblK0atXRD2x91r5FS8PwsIIYWwt5h5yxujL4
OvFZyY3x8fN492+odMgL7asD3WfFk2LB9oFHkNYRZpsq+tBnT2NGHgIDO82DpD/zjJZFleOfm9QU
IOCsBSH3bOnR5T3oAriN1wvWIIuClqwz924ldih5vp20OVPD5RLevQ/cS6YOVvld5wDHDmWkZkD8
hrFiQJaUnUJRpUPiZRyA+VKXPgBG7mI72o9TjByQA+PDlq3dWloVCVe9zqhPc88KfdTCpirP3YtJ
eNAd8z/LoTHKL0DgWKI4h5bfqkbO8VsTLjFPpXgXSTqOXIgmmUecqcyq/UBV1eBM1ZO/n6HY//rA
3j3PVB2cURqGy7WCnYJ3bymJ9q5QBfqwF16ed0JIjk3n5rrSg93CDGy0CWWOduSYfe15qssOCimT
kg/j7QD4igRhbz6niLNRqpEcxGlR8cG6a0Xn2MShvs5bLMfIuASzGME/1EWt3b5OMDMlhoE6VxqP
w6TFyID536D/NzkeOua0JkSLnTMCAgm0xabiiuRgni13GF1uyWN7VRAfZ9o8j011PvlYOPz2M56/
S+036dNqPTO2rZKouEA2yt6Wdc2RJH2LS679bJLWeEcgbNSG7vfVpYzjlw65TMRpbuRFHU4yYqSS
SZaLzCjIrqpKuMzUWlIkFXL4BAylH2EJ/3BTzZd1KEBh9x/+c2+D3X7lKgNhBz50+yHrQJs3AlQz
xHhWKSDQp5C1N/gmERyWbzT+rjWkwZKLmcEhKUObvEXjbgXUfdvyQ8HU/Kx82Cfl2b2a1+Dl6mCW
48r6qRTNwAHhAN/8ZiaUtZ7L2SZgmw6sdD9+Hb/ETOr+VdJ/6MYcLbGG/SqlGs8E2dHw/JHt6+Cx
/PnHWz0YY2GpW7aqqw8EpRI4fm7NeS2M/fcdsibCUcwTaV9iAE9eo8eBfYbpj6jhYmo2fHxXcgQO
yOgQBXNM1JP4Lx2thQfHaWWtcdgLp0BRFq5MzJgWJQF4Q1fX6TIkkzCdZS7y6rURN8PKKojcnmO/
ad5RtWt4KK3SyXB/xosY8T4uuBvB7J6AVmuntCkODsXaFhy5tsW38NJYuXI8R1MGnfI3Ph9nM+to
bdnqxM9ghoJ0hCNf/bEzrRjI5R1mPSQP/styV3XGyw80+0EGnpYBQrF0XH5xUw6eXl92d5T30ASx
g3XnSJigkk3H6wQj47Ja8httmq+yob0jY2bv32Ll0EsYXIsNW6HFlj5/9tF9g+EX60XCEf0Nv/tf
Rqf/woPjesvPF+Y3YQDLtTOJmZb1h6pfOsXDydjY+wFgkUAxtzYpZk1w8ckGM16Ojvh/kADCdTwM
Z4FFu7HNm8HZXjjRXXwONWJKSr5Ol782YrALccos++JhIjC+o7NO334687K1td8iBq7m6P4cArKo
BAbH2eI9YRNQ7lHXRdGvu8QpvFqoE9PLOHrFFW/qGyd7JXfK+P7+vJ8cfQ+21GKLJ0MUWCeVylWY
05YgTIG/dIHIjRp32jhHCOpLqDwB9CaI990bM9jjecdCD8qB/9FpAHfdyizARTFueV/6dV0/yZq5
bl8PdtMs4TDzTNSJNFUG/nDwRwF06bDH/sPyAtZmt0GbIsoKN6b6oOdYsBq3cHuHXmfVjEctByuu
1qUGGSvH374cdtWo7evIbMXv7YUAo2ClRJKqYcbKVqfqjf5IlAvWXtWC82OJfsVV8nZwz7+VwquX
/RKfU3ZulJA+KMO5gDbrOEyBIrf7Q0xSuLtNslJ/wHZQkaALc4Y9FYJKXK1RvVbVii8eMpCG5vDd
HXgEc7YV0ABpNKQAIFgnoN9IwnFzudVzaWCuW9POPljkp5PyJhN4Aw4h0MLjnXre0tZcnKUgIJrF
sNxvENqtfJ9GlRBz56Du+SjzBwlKTuxj9emNDOAreelEX6BKvN20LpCRauUV8J/sRM331tGe6KMJ
4obzULjnOgZYrn0e6+Cjbl0/vVeL7c6JDrChsnHT4GJUM3vXHdCzVU4YFXN5FqdvRt+9mmGAzbme
NVqFAMdfrbMD+dn581OfsJ9v0hpJv1o2ZFckLpFLg+BB4zxNoGCtBMDPxQjVlGJbJ/Wug2ZdwnJQ
yLTrqjLYEQwk+kpTYLeyTKa2tEudO/7YHUhR1zCBA2KB3o8cf+QRigPhSD/LWZOy5T/mZdK4RoSa
lf9Rplp7JwoKTx+7MAek1ODgnvldiVCP2GQoaNBc6qt0magTekR5TCb8tPNMNNV4gajpUFKRlVuB
ZdpsnnRWC7SQPbO2GmP3FKoD6vkOVqPthzP4YA1prx7HfduHDgaDEX1wZPO7xLxls7crxVWCcmCp
iIvE5PQDkEdOdVyxztiXk3TEGvZcAIQCmHyMHAzMHW1/Ph2Vh+uTxGvGxI4SQ/XZWHQjurwma6lb
UQc4Hsbd5ABmiXil/Zcw2aX6SbzYy0eaafvEHz6CspfC1FPz+EDGXpzYEc7dzcWAXNZHvOJf51h1
JNzQEJ3QpDQDJOW3OE9uAiU0mY7zHQyLVwlkAGmkH5Wz74rtUmTPmG+YbVnFpYdZGUtIZGJHWP5c
/iShmKyuQT87W2xwYDm8zf3ADvjZDbfTNXrqnv3e4DZp9zKztzdV6gBoBs/JI7E16OWqMWDbwqE6
6YG8pu6Um8X5uv3pLNAtw2xeHglAbZsZHyB68/duFn0KcoNv5KTdeDZKHrloWnQOM7Os5g/wepXD
smnlF+owdzlEPFTpzciD/u5jr9POClmVh2tYLP1ydH7G24u8Qmo6QISvYXp2B3BavRT+5Zmai+k/
x897R0TyIV1vq6MeeeryEe1+4rVTPgGYd+jmVws2LxokqDgRrombpFGvosAvRUnzZIiGb/5T1l3r
d+KXe5JobGzuGVgDe7BrqxqIT10r2um7lybwp3+/gTa6u895B2vKPoH0QwnFKDJOyzulAWxSflTL
eJ/G9F1ZtD1jEm+jKZmEoLfRLk8iA2JGGYshKm/RDRSqR3corNQ6K+eqNXl68JKD3g+0TW5RXrGz
7kMThLWTRA+GpB6WvQAztUuK+nmZRm8ow9/O4f8cIUxOJ6z0IVNa3M4uL0xIlVwleZ4AjyUnrTNY
rUVAJYx06PPnftElFB4aF/Co2ewOVbqjFLpn7IbMasuAsNErv8mBsgVnTZCYwGloUJMKJf4G8f2d
OkoAGXbnXvi0s8GVd5zBzmtywcT4uS0QXYFz6T3HkzqOIPzofmPsx0CO1zfl6mf55/glzA8yImRB
TdlXIVNj3rie96gMPc57jegRiO+/E933fk99NEx4obypmEjn12GTZ9Eovr4tOpkN1+uO5HnDmMq5
ttJlDsgvKeLeClcud+Qfcb+I+t65cnB7kghP4RDqHvMnqIbYWm/zT1e3R7IMs6o158TBFg5tBQfc
KrzSzuGpdquDXVQgNJcqVwP3ie/yz1NOf+kfaFvDqi+vD5wETjlFwq6TfDO5/0JrN2D+U6yi8yT3
HVzma2EFkVSLVeGBHjXBd52JlIhlG/+cpNjCrsbv/E74ajPyrrhV4Esh9EdAiQD0QyTfISEzD1sf
3IsLp4pOTrlAGiOkuRAe8/1b3ZUBiuEiOUq2Zd4/HsLmeakamV7Bcj5X31Ua+S8i5/wQnig6reiV
5xFwnqhQRlWcSo+Obj3YppESnkDveCIPfDRKNsDZchCy9CHNFkNfL8RQRyhWFnDTvOzIaxiz0/N4
VDHXLXpUkjn40e3cFm4zyqHzStDF0RxC+acmnn3sCJX3VeTHBVF/k25shJ5ZJ0Q28tVziY5PWxsb
F6Ovx6LOVx7FmIeUkw0hio1aLGZk+Okax2N44xUEpmZY/y/3pk0LVHqROgh3B19IfgsEAiteykL5
/aSb4e55UlI3GJPN2S19Y+5YtKGfAlQBxc/gINkgkEByzKsWYKjX4N4j6hLrZGW6HEgB9dZEiOv6
N0GnJzAVyzJxnKz8CQUw69O4sYvpl972Hyv6bkxWA4p4Ymsb1EP7HJxm2ykFjv8GS4UthLnkhZls
l2rFwtBCj7AXbmAnSAUv1O20JYKMCrBccCiS89gZ1h+BFSqTYkbW61tTnANq6Cvly28GJ+0KZ2jm
5pqJKlsGYbiqDJomp8SDx4zVCF1v9CVoH44DnUXaD1M8YEwn3MEkPsu3r2fKZ583cG0IkhcHpr9K
9Iyf35FdTlBSOqBjF3zhZpyJfOjiTMKxJXtqZsmxO8tjMiTrck09aYAQw5n6oxhPBZfu/UHwfASr
DMhwZ4CSnMgTQ+Zc7S8MSQpeHSpV4G7TxL8vxjc/Uh/4N3etcJU9xEI3TV42Tz/Raqa4Im4UBBFE
/+v/1f3WTmEf5zHgabjPRUBvBOgrcvmdEpoQb4WpjxdGahSO5jVR8WmfS2x2Krsp+oPd/AsYiq7R
eXYkOqDGwJ2MfTJoNpw2fUlR6mA+lXjhT5g4CxuB2Dufoy8cgkab/i7Mg77sbiEBnN6qDSpdkMN2
otrW2Hji0R5JvURnzljKnNMqnnKkjn1jk5L6ecZcHgBFipW6sOHUreaqcQle/Ctr7aQG+9pOUsj9
yqGzuPSK+266kTZqOa40pwfgC8x8SIeC8CV4aFf5uWrlzuD5jVXrMlgAF5WhLIdv9DSZFcQZ91Ot
b66VZ7b5OIbq9SVeA9pMWOWP/XpJnoMIrarI7VNVFbjcyMZorNLBm+dWXZ1AOMRxuS8ty8tuAr6y
/RH1WZdCL31txS12uNQu4hfSSe2NTXOvpa9JX7Jp2rXm4Y9AV2yQL2V/ihrha90A2OIjqpLot7jR
njZ8LKZh+Mb0PMqiSjyaU/J6jJwvBi8RYMsw/QVSLjU6dUeckmE1tOQ7KqbtKMSFyfXK9qep0Osy
LogUOLzC01Sk2KgaBDFS0Zxgp8arZa/h9h6AlYO8RdcUe8A1daOwODehw6sg0roN+4/FZ1h2Bp18
kbWf+3Rtq84oL52IJlH+rhb6m/bvn38G1WFOvAASdVE/GBEEJV8HFIhCXuVCIvaOX/EW3mqHZ1oY
EzWADo4UrR/FOYW0MBs1agl3pGmA+MjH3Yar3jtHNY9fhT4kGzz+UgdHvNZ84kuwgWAUDVYa+r2b
DvNu/70i4P0K7gxKAZCCRBXVvTjZKQelS6igU0nFgIZ3Pyd3TDBckGVcRwjn9Ggo+UeVxdTF429U
YVB9NL9i7y6WeEo+4DcFFjh6lM8PDGTjsd62hYxVN4LGzotOP2jHTa7HBI/faZZJ3A09+7+0dSGO
awJqKwR/loP7ImRTZOezEXe3B/px09BJzB3RCv5Ue73zZCqQoGH+co1AjsTIk7lR7mkusdg3IA5J
wkeTUzulRKdmY+Hwdb77lTMS2PUDYtzceSNdCUCcNpJYYOhrKtLOyVygrylmFu9CV1UeGEkYslqA
U+m97hrwcUmki+PlfYVQMHFzCeCWKIFxDg78pHFnJOuE3SqVH8Im8gbsgstu58c8zlCLKpRExkuC
fDAhKjuFASmErSL9ccy2ItoWgYSSg775uHvCF9ShkNNEvfyHIEe7YjG02AV3cq8ffyzlDLJNevuo
YISeL0s3WasC7zzo8xehhYG+iEwIavxw8sdWoQW+4+vkbbu+jpHQHPFbft3PEjlOUF5y+4L08xHn
5TN3ZgD4QHA0GGau+nvBgaJAx2ODEkCTIIGjjNvxXjAztTPDQnkM5LzBgHfFQyMRRBBUfCAuaKal
zAWOd8HaUn/I6i7Q2pyT4NL1jZQPgjzmRBm49YOATkoJ7oO4BoqnnT7KV4Og4UyiDjLcn2YSlg7s
mcl6VQiHrsXi7ghAVvRCKujds0PDlohqBJY8ni7h163ZY9CVcRQ1ETrxN7YwY2UJYA4as6916EW7
rSCKF7YARhEJXivCdQgG66lT/5nZXnTvtKx12tCYZe6Nd47c3prs+FLQuDSfTrZVbLwO/aV59QEf
sDL9QeTuYGeCLJNJ9FwYJwT6MyWbdSCx9IkqoxBWVg9YEnRUU4CeCo6A1+VRfANaeGXgPl8CleZ7
EsGZ61VjmheD1AaMDH9ufwKZM1tNqbwULEZ+2xow8eTFEesX2Zgz15gGslhcQNChXwTKa7J7Dk3B
YiMbtzO04lssgV51qadCWpCuMVuJ1C/CBL2jxRniDYWwSKQ6kaaS3I8Jr5NnReVl0udgjI4mswhD
0qUz3y5ZzfnHofSx/TS1tzfdJsTX5uXaDMIanv3ndMYpt4yMmgkj4dSb7FP9L74wPuea100fUoW7
G4e3T0gCctnn3fWrtvpVMe+L4JoPXYgLu5KWBnEQIeGpMhkXjp1KSpEa0LTb3vOC6tnzOWz3SwV9
hdpY5+GYupU3SLmYElIH9L0fdL9YhMTUYiiJISn8hGIoCRsLBXME+sTyAjhISaVtUMEjom7HUoG1
eKY/ZLXDyDxMMAiBdu9ypZIMeIEQ0TVGUl/3czzLDG9MMnVy/z5h6I8xSp7NK96zeviRnQXtryBW
SW58gcD7N9j3EGgLxj2RDgJ3K/0nOFFYnXTFf6/yk9rLRJqU79vedsauNh8+JhSwBZwh8u6ox3fy
EirXyYNvq1qIqvj7bCSP7kWex1F2KJNP3HMVp2A5AI8XdCZKRPY0NVXRKkqGcBp06duyfuTx5LgG
KFw1CLICskE4QRWH8bwIdD9qD24NOvhwtCahCwQ+eKCDsGeZiuZugvMex6LVC7BBf5i3ul/AN15U
0yyQ3Ub6zZJ3HXdvid/5OTAgqriV52E67p92NPZAjhS75JOYk38XqDN/9dZ1yFssNcgU4C++Dl5G
kwwNborB7AQ29iF8oqs0gQZNxW/09PplJMeHOQRM4kPEH93Tv4eAQgm0y43Rf8k8PucmQ0bitWO+
Hg/zwRC5uJDP0Fpfh7iCWNkByl1BEBEiwddW5beOCK+V2j1RGDLlvWsc/zUXtitTosLxImFRyDM3
WLcfvxleFEN5wfhMgMCL2YCzzCAzjkDcpnzSC6tbVezWVEoA045uWKWL4iPfccteCfEodRQG3pJy
/3nog700x5HIPNBtDlri3dt3J3gvFuw7i/EMEG9Yy6bW80DmfSaZmCOZe5Os6gQexcCPfwwOQgR+
9Rjbk+0E+EQqmZhoWLBXlXimvSg/lP9vGG4XcaSrs/SZCUWmpbpZNBnNmPNCqK8JQdxCngHooEZ2
YkanWRR85vWX6x036Lzh7ygEk/rLeELsSa9t72bthbKH9Of8o0MYTzAoaiERjLGHO6xjbhAcAWtJ
0HFlFZC2nq5M62IR63+UBQ9mPc279NgeTHSEPjp89jTpX+SKUD0jHvOX7yARnBw44UYpgmlJt6fN
d9vZGPqcM5ktpL/RzHEAQvTzOscn22cb2TJYZkoKIu+yJ4LkXwWjugvmYcFwow1VO7ev9qIxTzzP
ps7JYP89r5bH83jXPFBlKhU90cFnCmtsqLFWAzs5N+xV0C4KliTJofU/eaS2hvjmAG8qlSbSLnvS
atZMLAxgvb6MPk7hNchQYa2KFgOMs02nBC3EikOi04SKlhnbjUfrY6q2ueyuXBgv3Jo6NPvEl1TL
IDY1tdJNx+ICBvWSmujhQ4YaPJGIlAudl7gbmUMlkuQM67QI1J08+Sd6AxHShAYyCDPUS9NF+1YN
Buw9pO814APwbauhAkL5AG5L1TeA9hjWw1/QSbZWARA4iZ4e6ADrCT8sY5hseMfNK+01KF6x1ulg
EUZow/p2agTny+cvSP/EHf/2913y99K6uo0aq3sCQrp21oHE/mV3VyT5/83CT0zqUsabmX7h3vhZ
bt+4xzvVmHNxUiDdJ+Lc3FcRvk2kF3x374tOU8UAOYJX6STcttOirwpGnw7ebquqlOJwsy756RYM
1COGWVTG3coenXbG8kWNtMXcvh0J6DQVz055rHmsgXN6ecv3wkrPpIl0D0zC4tA4RIXzaZXDV0iE
Dvg6xDog9IC437vMELOmjApiXWxAXi/jrD+4Nu7ELqBlYzWNlrF22QZozNRkuZ9d87doI+A8g95+
gfZadryqXK/o9SdhhnX0t2ACcg1apYzk/DCak7+gutfmKwjzVoqt713aL13wBorA3/pBDNH/kU1O
QE4BNWqn2jZqtALMFsWFL8RO0NkgiaJuZ9K4bLks/Qu+TOfU3AiN/Wkz6rFusS670iMbiXczHEYl
4z7sLFTCEjFq/i8MryuaaK9BEi0KSllK5AePY4RUupMwTCrfVoCcwJXT/SiWJcJdW/cieuf9TuOP
XUS2r5VZVroiVr0jlEN3CPgn8hBDrr4iuhe1c3L/j1u5Vt35LbrQnbfTYqKlMSG2tlry5VVhKCmZ
VZ9YMqDPQR8jk3QtzUSgodtRHspljD1s6hnuF8RRuy/vtfehi/AJsaAn9/REI8F22LqLQHtK3JLo
/xLTKJdSyUy9UU9wmL/4j25WOViGDfqD+2oez93ISGndge0BGOL3OtKsO1zaiUWToR+j/mYKB1om
D7Wd8/cVZJplL/n0oZjn4CI3MnluJq5JB1nbsTbkRtIFIwAUZZbJyjZvUViHpYrYrXCjy819h+gv
k22aZYEONhX8MYQWsIKpLxjKy9FyZXy/Y9kgLGz3Z/KqhFwc6abO5Tr6RujV7eCSWBSs536whp/F
`protect end_protected

