

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
FEMO5gEygrepbyTIAb6bnTzXzKtTa7hkErwuF8UlttB0u+dyJHGgNZ7crkojw8pXdXDcfF1p7dA+
pQaP5/BGSQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BUAwVhxzmgAogQkTbbeTYgQQyI5Ea0fpFwP7NYo/fJYalzsEKCNo+mHLYdEEN5P2wAyI2jwL1Ldl
2cWWTvWw0FFDx6CAqyMZZ6MjBcXKMrbvZz5x1XnEF9Yq73tmyh83lBHL1QeXvwFWsV/MtPawWibr
DqrVdukNDMYsS1phrww=


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
S/0xh+8q5ei48mqpxhA9UHAZBmce/qaAZdB8DypuX8HuxWaop+hJCz7/amofM8Y/1RIn9ynwmPIG
lcSFISHwXxQw0TOGzhwmVeIUphOOW6Xj8efDxrEsgqjlN4uFDONpJWsykX0bjYlxDKh7V8VYmxsZ
W2QII8Eg9roJuKe/q5c=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
m4EIihJzHXIjlJlX/nPXOZoP0R5PF62b4QI6DPL+tjjKUW02RGUxgKdMgmE9mHps5NWzgwv1KD8/
U89gIWVIYKuI7AkCRzSIq4+7kF2eDJ/Rkcrj2wW4xn9mJfkpoCsS7AtOGt49NAv4zZwBC027t3wc
ufboERWDi1EvdAKPgGQm9PlsQcCafLmx2ptvdo46UvpFqzYZ1W6ZCuZOinFXuDbR5Dl2XITXUKEf
6Qit/856vn+C1AiQMPBPg5t84jX1T0muMNdiJagE6NH9TuIZh34Zh8xMpiJVMleWEJ5+ar5ZYsLd
r0bHpLmOwwOHnlbs80+gfl7gGs5ckUJar8uTrw==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Ugm/yKAo2KdQRz7pCWPXE6yTuk91zWS8vqvbp4N0Y0rRLeVjfYgYNsoxanpin9oKBWGqB/EwwFiI
OecyJhZzQraiaozD95T8G3Czi/CyjQfIuIxyZlOURLuKQG7CmONNSV0/exWSPuBfn3Pm6VM3OjmU
JLfuRDs2d4YDFd+q56oiiHQQ8vCWNnabDnJXcPKxlSBuxC2iBafhs1u9xdnlfbPeZ3KQYthd7ZgT
hC+BU1U9gXilj5HY81LPuP3oaZbJJceer+0o1dASuDQYfcDQjic35pfjZvrWfHg/SGJYnP9rBSDj
+CEsTamUhMcogvVE3I0C8I+NXEkM9BpD6lpS8g==


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
QZqM4wdZAFPtQs4YrlRwMrWNZIys0rSI0ZT1kN94aimnqT96e7hJXmu8OIn/cJHN+QLJpyX2bZsb
9aS/bO2EpwxEH9ivoPATAnDH84ywTGBY0z4TDTpMdmLig2F5x41qoVx7Xjt+NiM1WzZMdOXtb6+T
7rMRng3bWtMuYeGIO49nyrXfIsdW/BWSAUnc7REbccqnnz50wxmKOz8/Cxc0CzxowbVvovJtn85V
3ZbWUq3enzYLdYiG1rbSQDaPniVAqH2+PhUK2ZHB0HY/TJkgvwTPZwQdfAanCA/ekvY9LLeNdJeh
Tfdqj+WcsCML1NkALEeSJjr2A1ERcuQwgDCfyQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6000)
`protect data_block
i3e+u4mQuBrPzehuQoKgUqMxB2oUH30A+dqwqWwlaMoQP6Szr+IqCmnKZvBLQFZrM1rsukuc5vew
rXlaUOgNCZDZnTD2rWRQtQAFo4knvgqAAOPCRtNnyS9LcHtBQSdKxxEL5aajOUI0d8PgKBI+PTv+
MiFnv36/2Z1g9YiYfUVEZHzQ1YmULDXMM64KTRLs1ugd8463BefkRmfu5u2j1KT7ur5teGbu12Pp
ioiA2Gea6TqNy7su3rXAhuXkxwH2qOA3T/jDVNtS42T9AXli7J7G/1OHPiMNlnSpsUMIW0GQvg5m
pUb3hEBVd7P2ISjJAbJPGKG9hH/djo5iYfDY80kNb7edGHv867UXnzgoJj/o0T5H0a+YDM3pMpGK
YyhZG39YJIglDYlZ1+E681U0jdj8iMYa1nxq8XbGEaq1srucw/um7PCIqm+g2KUBGn3ylB1IPjAs
7tf5PEVX6+13/SP9hsFA4ICo0EgdwgGBnYOeH1pBP6CYK8fzfdO542KBLFGARN/gzKBwHzw9FF40
7EFkivhCeqFYq4Nn+w27l4g9r0H5wR8x3o6juHO7s9HXTsSkNp5tOviGSiu8OX4YoduzOxZmTkeS
vMAX79TGEPVR3RLwY9/WJ8Tr78hnNWKbqViT5e2l5rGKx+KSTSheu5vPIPIm0+wUve5iE5Sg27Gl
HU1NEXbJJYAF7Tteta5Gvs4sxubmj/q8NBvAmHSdSaSWwSacP0ygjdRGFpvyot3e9eAlqaJxd0sg
60vO4jDTbN/gGxzztcbeUBUvGxPsbQZshAASHnChiXw3zrub+OC6oJexEJoRiFlti+pEEdJVLmRK
98UU1hEtCrLgeHAtGPBAAz4bNNBhCoRgLP5Q1JUr3KR/HidAdlP4KhuyLEWhqVB1L+IQPIb6wC1n
fRnJBhSSiTliVMh4Wy+3A6qvruuZxQX8BV/AZtrNI/pCEnyz43L9PMRboKTt9FXZ4XdVcjbkRKYB
MMhbVfF+kBnUQszz7PKzaLz+3PdCT9CQXGN64oImoW1Sv0Fg2K8AiUw5ehwH84kpabVZoGw4heZc
IlG0vLSksSlBVV8keo6w98YWT9Bx3Pf2NaZ+2eUSVyav29hRhjH5CNN3bJHRqArjzImXWQyzOLbd
dpyqxBpzxlQ2InEk8h2Xy0QAOCDzN1ZOaYpd8QhcBSLqLsv9sOYYVkemHtj4Kbq5ZP4TeFh6l8Vw
sfhTiC3j03+pCZtXLHVytiMaS7dvxq2hKgBlMgO14oDiaoFXdatb9DeHuEu9JL5GD5XlnfiXJi9t
waf0VQxXbNC5NkirBbnxz5usNtdgeQppWW/p9oBsvir6JmfiitMarKKGPaLxYxONE2ZhBsSqUIi1
Q+b71OffVQ0ItaOAc6QDV2IGOPOaA28NdDJe7Ln9GgOq0a3xDx6Ef8BFWWyxLkLEg4AEZSUyYVLK
kkkjGEa4zkjPU+5bG/dl8dxJeV/lMSO2hFqpknqCTqNlSkF2ItpEYLHtUhJYrACiRn/8FgRjhM6V
KOKPS/nMZuMZK3YA7T09FBXCPy5inZZSUL6+edI7G7J6Px2SdPGpqmKxC5VUN41DLp6mhYvK4HMm
FDCj4X5X9+BqplxZ+86yzlcG77vyp3H9imovMzbW2sdCoY3tsuUcs7LE/SNsfAdHOsxXUaD9EwKu
ehUD1WI35dwlYrssWaeJdWXyDdH7JveNUTR9NVPQuuFleFF8jyW2FEfCIIzJ8KF7EsMMp9e6RssR
XDnH8BsMDW0Gj9yBiUiCfLu1w8gRTUFAQXKcXmRn1T0Yp70/PI3yaF4I0ayVu02OaXA+Bsr/bO+9
nlTgQpqdWC5fr4objzWdxYLisye6aVzYZlISPi4iRFPgt/7N8elgpuJjYGEk01n4SVxyIgoloybY
YwEpX/idp1tu1uy4Lfi7stRt6XdCRBvdsdxGJGHVl6qnS2hNjx6roDH+LfzsF4gAjW3KkUPCYhSK
DJgmvk9F+fO2grzSh9KGObV/bB59jPrCG1p+OWm33yjCqzwKmh6v6wzqx4f7tDXlQr9n2mUW/cMh
iulKFjEFwxlhoYGHYB5H1kOoFRDZQ/d3zrjVz3MlLpSpx/OU1E/Ut2LqLFU7aZspTElCaMJc5mjS
t2vWpFDQ4fxCrLTbnNfZnyBtn4lAgQ8oB/ZBXCfebTRQVmDKWFlmz7KMJ2d0C7Ioqo7+GWj3TXCg
WhO3RisgFUkdhtU0HzHTqlnJ/OGj/xAo6CrsK0PBjjce4GI2/XikzII3SrPh+U6PO+VFGA5j++aK
dJFzCFPYVzj3dJN+zWL6+0r9s/KC6h9sJgMFU6jNoWiVCHorz3Ycq52sPeIc7o35/hijjwz12rST
SpAGI4CWWNurxYRSJhx+XTqtu4SyhANo7h/SsvlCiir1yajDVjNIER2xIWy99p7CUZMjrUC73i8v
izEnKOj0cW6651LKg81VrBkry+bhMAOzT6xFDUPwPNOk7mjA/hNohU19FJ4iMGclPkdRk9GBbIt9
FnBcHMkojFbbrmFxaHf4p19vsOWBfy0pdLNzRuOmFoo/9FqN2EUuROB6oDGxMVe+qcjdnWtad3zQ
HnpLcTV7cAkk+xuuqnbjYGaS3YX2Y52Zhf8kSCO/YUd92kMlQFmlsryKFJp+5tssHsOgxrTa4r/q
GUjXrMEQaBpSjiyKe70ZW6Deo52DE9XzAEjVwPa1lQVWZxIu6Co5CWdAUaO9dVNPeFTQvWAOzf+X
oHz1cvuhK1M1zJqAk5ubzSHsxp1r1IGAkqlKrvCVaRijAgRLnLZbkI71YTt4BS0uDcuQjSzW/THR
fynrbQGVI6FS6y94yz280tsZQ3P5aCwOEX06Vyq/leZKIXAe+ihvJn2S5zfIqRdFrczbqnTVYwll
3KqKb4ZSXBd4Ub9+yPA9ObU1KErvrORSKVooGSQet7HUMvd9qaKX6871Hng/ChdpmPhfIxo1xY5m
tb/ehCmFbSqNJCHRKBte0yXhiFdQPHvV4783/4cckyeg9YAhn8yUjojVt8RhXb7CQiacglxwu/4k
EM/m4N3eplmXMJFDH/wEY2cqLFTnCAnjXl1s/mgyoZxl8fpBKk5unDMxTOZeZwbDnJF3m0kT4v1i
iuN+NV/pVRxbtsqxeWlAsGRe5npKcHRaOUVE1+aVXxGmf136zBxF/gcnPultcrPIe+3Gva/OOp9w
h8qq1VcVWCfZytlalAGwWtARuXYtVYJP3rmwGbtzX4BoNTtWlWnSDjxKcZcmOpemrMPMZvW0AJiz
yF+inZvIo+kKLGUKLuENxgh7nkGa/huz1lFZ1yqeE0nnKPRR3A7fYrqzgTTR/SAtXtPaKW8f8WsJ
z0k23DZj3DxKYMTTYgqjGuuYvxD8znxFrjrUnzcm790bVmw8sYPQ7ks4Y0RaJw1ar+SmBuGje7pO
i1gk0zWlVJuYKCWbZOBEc2uVjnSgSq7a8G9tvu+q6ig3thhI9ZCxsdTODmZ/Gmzi1cMrgNsdXfo2
MheECEwU98KmOPkQ/W82UANCSIeFe7E3VE/p+dKs8UtDOtjiC33AeY4f3WdxjjMPTshZ8v4N6io8
TfEtwMj0CzPTeTyhfsRNYnPFXpfIgkXlOrUM6ePQDdQ2g1Us/cfN9E1nFdszIZJoeNS29NehMsoO
0Ebt+npFwV0VNcjIqLxCFrb1E0PWKzBTL+F0DFKmPSc5bbmIQqYlM/hR3eCuQssIq//zAYh4Mqn6
nnJvVL+PDliKmxaVUFfuumuNoFalKMReLFwp5s6Gn3WHHtjEihybePYshuK/klLvITF4JwkQRXRQ
FhXA9J3GF59yQCE7dhaGls6QlKqjzHWD4V74mW8MQZsA79n7E2yymEee72MB2dzqRsL0a7gVxA5p
yX0CV8OP0XrjQsaX4UzhsxVif3I7tYDUjT9V8fE+XtRftYj89EPf1wfJXNnM3OBOVXx/zZ8u9o2H
4ML9A+ealrMKDUtgTczHJnCJ2vl9bAhagXUWkKwsuKyy/cbMcB5JDEGJPv2zk7Ykky8ow7EVmf/x
DdPYVgEx60B7+1C3cPyjBKTXVjA9Ry7/ydUF/nm4PBjCOfoKbLDIXq65hn4ukW1mR91VSwGqqufC
lHEnYUd6k8mnysKQnkPnkeJZdF/bSHjsLqqo5CuFHbI1cQ2rjtm+vM8vCJPQovhjm9N4l/ZAO8ir
0fSyRnJZhbdf0ve9RTwm+tidg1rANeSj7NkfwbYPN4VZpywNtK2A4R6M8ZqmBc1nhkBtQcPEpjq0
UW8Z2K4HptCZ01ZPyN342WbzkBHUsQpWfHCLAu2nGX7HYwLVKSHT9RlFatLSts/ENfcL2AhgCHyX
UK83pqVDBzv80mPVzPDEnzeNUi5n/1+ZTAzNBLFYQDrNOI7PjXgCBJgnzuw+9z0CM/+1HBXkYX73
In1xT6+gkBkBGfsrxVy5/Bm5OF/qf9wG+nqROzhvrrXznMQD92ho/2B3dzTT0tNtWj8pp9ToxPLU
p8AKMLL8nu+xU5tzaevEGWdIbuDJowhPztFAMe9bH08OQSVocvoLUSNUo3acY+MqloEUBat1/eFw
TJ0wUo/XF3iwWdGlixtMeWZ8Mh5CCvDY/gQ3tp0q7J3wFWnb39uxI5Dv2zm879cQc9YQsBONZ15P
AYJ45K7oOzxx6QK/zcgipsbXW8H+r34su5HJvly15dIMOSzorMHpPmS98qYXCR0WrE99j72cBd3s
iWWYPWVBAEMD1ciZgGzdBlckniJdU0RrEqr8yvM8YoT+Xqct75Fq95L+yazkElgUXSccLDwsTUyQ
0OlJRBKJn/8AcOSF4bPkJop8ppbpouUTHD68P0HNQZ5UG1YOy4CnEC49ga7Is1e84Mv5LxenZc31
aHM+zdOzBNgAqrXDDQoqQvkGaMFLT1UHaY/7vhAeEnDpGd+SQDpRs5kjWMGaWmcak2BHPa8xa6H/
/qxmRsMwap6aZatqmrquJOa8SRzKcGAL+ZfLRh3CLwtxLe0mjnZE6R0FVKBnqTJy5IV3Yblfa5iQ
889dZH3ML76ImPx5BK4hNeDpyKya1KPEHIEuB96wbXWI1+BdpEeB6RSFIPti1rzfeVrRvJVHbxC/
Qp0ylKRJbdoF847Tbgzeqokr8Cgh7pk/yLW7FHVc3epiygVSm34Iw/RUthJGi+ksOGdQWXDgk5LB
B476sKb8SYnWMLrhSM87Bg1XJvs85Yb49K38HpTMbf+1oL+C4FOMa/omeUwQlxvxFHHRRho7E+mw
YkKHVK3sFzM72nIp3+oPPtvD0Jla0sKTQ5SFtaUAv4FlcR7lQmYi+qklwZsYKoC/RnYPYzvdmiXC
Z1gkFZ2xNGqlmeyOeqO46U/dcp5SuoxL3063PduHGzusmoVJkRk97m+yUQkiWdt/cPK6afTCHADR
oClj0lyxTZ+FMTvlPMY8UlFCu1oWA0jxAXyIipp5+5Q19gIzxS5+8Nc6OPSVJua+opd1TpP5yxEX
v0tSm4R8qX+A7cDQ+GXqOJSY7Nl/p74tgn/bUpQ0el3jH+FSHjYsW1J/85PNCXDi9ojZz6CrM6wv
MM5vxrb2c6nKnMLdJHUOYHu8hpCQ+Cu/n2d5YkecOBS9zyafZZmN5lvSQuYaXt8/SdqweUSS87h/
UzcIta64JOg0fAkK5ZvMCjCHstBp8mjfsowRiRi47viGGKWCvkrdfRT64qyf564M6GZHuDLoypsh
cJmbXOe0/tnf+RUy9evndCc8d4D/DqGmUaI6wOzc2SSpLjiSYg8CF14tQgHeNnrXFYKEwh3cSyzo
PwhYw+4WWn/DMNhPIV/diXKRM2kl2C3vjYLocyfNLLSfQaJjKZAq9TaJyCelyrV/fGYSEk9Q1ybj
dJkSa9gbBS3KcXjZXC19GEyNsuhhFTOS+mYYeHkU7jQyGy3F7ACfrMVENGKhFPm68NXSH17Rv2Ot
fY0Ba11/AfEEtgB1gZqRG4oZs86sjIZSSv0CYlGzJXu620dn9+b/zzEbL1RMm6Fx+e8VhBYgDaNm
+6luRmWdmNVKoADY90vY1gbj/GLffW01Lr+OG3FO/UVtwuJNybeTxyStpPk8dCS/36cESoAZ1s2R
yeVjvcXLtSgma2prp1Nv92FZPK+CsO5E2e+CuuBx6iwnUXl27Cz5DicZ7UZwoQe8dIMV2xJEdIxX
uNWLpibJV3AhfdzqtDt5+gj9uCkpIYNtBi5NBc/3bgVmeD4Vmut0HR85ct9SnKFZzir4d8SIWJwv
gehRtpwHC7jkn0Jv7jU2Sgz2MAnsprys91dSEulvreQ3D/iCSMdWVcyTUaIojaocu9nBJYcW7g0y
mkYR824Rk+XNcC/mOdqqmWqpQRKlHYgMZ4xaZdtZWBc5lfehzyZJGyHwBDHwkhW7yD/JAX/V9fL0
yTpl2Z5xs8SdyGPigfPHCWggBGHWnUjwiRRcuGDIpmZYw1DzX6uWNFVZ0VybuTOBoBAYwWIZ+/s/
gvVbnroQRHcJicElk/vq/tb5N9yfZjUcc3jcZErHQBRFew9x5i+5vhlBad/XM+UoRbjTTCKv83s9
kjBeVkjJPy/Q0yreb8tSfMxYfxAYeMpHj3wdNsF/NoPLL/6hpa9n9x6TJRoZj3ObBCH6j+UZHvic
+TNiyJtaFjDdoRhuaVoLk091KUsy13rCp9WaaQPonu1FTI9/2OTqr/i4lkYXoAvGFKZVQKEXvCEJ
CWmelLP1xqLgm+8VAkAjOOQZxw4TEdALjNYt9bxS63nQPc0G6iwE7AsA2x/yciceBj2GFxWdhi7V
ovf4aJVme2aVv1shpq9bouxHhqMo4bPnUDIlAKy+6FuK3Zsv2bvnP9JGr3kc2M/XJqqPXqthrXIx
SaqDquYrzRRwrrdhlqmFK4zm8Vhlmux8qcTRtnHlkU1ken+Fm0hGvP/TJqP/E/FFrNGZbTHCB2pS
lIP/cDlwrXAxlPV/8d0C72Hx742Abb0TRbIRZksaN+idytdU172ZQOyj/njZTUpYaPSYIN5krE5h
fTrvM+TpZ+CjLwkpDJ7iZ9M26MGapsrS+Icun5azdXqN3rIlP9KXylt7dB4heTrXfHMYm5ZWqA+v
SIEcVIgJ0hW9iQVyx/Eca5/Rkmp6ohs/Z2nB5YVgn6Ij7v6GwcB2u1usdPvm4KL9Uq47yHu/DyaH
tHVpmuQhpUUJifb0B3CEF1zXc0QcUAJNPTGNkIE3BbzrrbCNjkSiRQEkGo+vuipNlS+orUDLDYAT
tYH/45g/e4PEqORxWBx+JZfAFCZacESdBwCz931RDLz27lsRAO+GuBStVE9YErXDYMWxXcOfjzaS
ur+LL3lqHCz3hCr4tTBQWNmaieGpKS2IXdGw7QuUiupW4Kcng9Lo0+aYCImoBjWaQfvLPZwsScUZ
l035nlFgzdqvCsLVRrIcemOFOIyZIfhRHRG0PQMKEVLP59/T+WJG3p7Co2jgGzqsP9lOUIpeoUIm
qn6/e/n/ZEgtDfEtbMjIidgJ3kxaTtJp4JL4U8X9xFxA3JYbpkei1x25Tfu6TwvvCQ/CvY+3O5hh
0jrxxqXRwBxFud91Wbk3NAIlh5sWh0uC6ZPsafPKfh7xbIiQBNEsUy48fA1acoXa08NCXij9kk9P
jS3sCox883xinUx9nQlRT8jeezCIECKHPvprlYWAnW8LGifKJAiF1/DotPVp17vitmeABf8PlUE9
Uc9w+92iqLRXls20PAV5wixoW1JcKdwvcBChHUd4nrNIjdqT/4NSsVX9kkTL+CgOCw18VQ8uhWIC
QQPyL6gOR0KcsYgSjZLEajCYGaTMsdAmTYdPgbLKgcfI9RLC+rG9KtL0Oxk5DwAMYNJFNUmE9Xq1
S7DubNjwdQ09yRaqnEA4TSxEl5YvR9pBygDHUNx4ua3JKHa0//Aa/eIj79LbDhhROeplGQ81pk79
N/5zL4bAyLGhzt92N1maqcOFzrXIQq2ZbEEzXdThGF+OA67o/UVP4Q/7vyMrHH+3saMohBd2EiH2
xf2dkaXYY/JRNmURUjq0
`protect end_protected

