

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
gD7l84kB+WAh1ATog3H36h0/cMgn9QL5jGe9p9PjvP7N+FJAVvGVlrxcgBw6dZaWDNZqNANQuRFv
ZSE8fsSCFg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
YQUcxim/tlzHeVlJ7otHN7u41KO3Yg5DFb1yF4GCsbXGLtUvWNlkFjY+UPIlgYImR4Zo4dTHJQ+j
3BaUNSUOqAVzT9CfyUelv2YD2ZTfAtzIe1Mboyb3+StKnuzxnZmIhVPiZlowdW5lQ1r7BjDPOsge
ztxOfUTbvYcTUE1ABIE=


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
eu4MFD/NMz3pssr62VCh1XDd9mthYydX9VaOq3lWUwHi5/7e5dl2SAWHtYwTnBgGPY+jCcMycJhy
WSlkhQxVj5BsMm2aAItwXFvH2mSbjlPggtI0/+DNGQ4x8LQSFLTDYnnQbBrHlJymsS+/asMkXACD
SJ2tF8LF5tMhAlMPZZ0=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rNAzbNlIFUMjdhvgzZ2FokzvR4AuFtV+1AHGDKa9QgeBsZ1e0Fom48uKbJ9iakvqUoUcKKAvRzeY
OBkbx9P7Imx0gvIgzFsgiVw23cBYWOhbhSqVb7mef9aKx8yeF8T48n7gKldUkwBHIPeqaayRI9/Q
HCZO+k2+HCjRZE6L/Gzd+IOdEVUFOg3NtWFPk2JFkfZkxs8X7Vg/xxtvH7uvp+/EbVyiMbnwDT/p
NSqOyA+rJwBJYD3xRIPTFDI83XJLCF+1i4E8hyu7Y0F9MtjKugqEHwAG+JK3jde00nzNNaeLVUQ1
OfFMZJpkk0Cg66d2cvJY/G11oPkmvTq/JZ4+5g==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
apuTRT8aJu0TR7Ciy6ONiGK4AT7TUEiokS4gFf1g+kDg6PdKk9VRun4HKszIadRtahjPQo0of9uS
yvu3GS4EQo+Y+T116wnAIXnZSa8EQaEsDkziOI+rCvXv8IgaPYN8Cq0aRlASFL7IHOWNI49V0c0A
FIG/+5U7ZyNQFCVwuE4gCgK/pA6apm5kY4FGJft/EdZ5YAbR/nCTzK4P53+XsKHrtGfw+/MthFWz
tI0OtloKqc7laKZWKOVFqWq8Qmq7UL6utFODtxEQqzczH+q+Gw4rkUyOosIY+cbB67hX+GlmXXEF
jMwvUcen9t6c+wiH6rmBDcUIiuUHHz6q+jCwJQ==


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dfDj35aI8y6zqcW/IHFxmCDw2mpyex25qQAUnsL+tIRxivv/85PqpCOrf3b7NWnwUKMrsxtw+JBY
mtlPsVxQKR1gn6VkaHwbEgwxXXxFe71Z+1nWQhfF8Nt55jGvq1joWKMrurSV7Mo+HkvHMSszXj3v
8ElD0S6sN91oml0nObejOhxzHf0ybK+sGag+CFA7aBr4k4rYglf7AzOYrPl3nNoCkyrFDQFa46/w
SXJm/os7zUHbsDI5GGUH3BU+NktHZV6GK3iyhtHTwrMgDtpGk6vKHMKULM1Gjv9g1/jp9Ao4cUhr
bCVOXM1v2e8A3564rmh3if78zTzCKamPRAB5Ig==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 962560)
`protect data_block
8aYWzANd6lzwkn5rzdbEEtfENNGg4sgJUdTFXrnaST5tT45+c77H9JD3ywRpDfxXnZYx3Jqmwi2P
mXjDkm5OSe95Lzvu10WkDrXWZWJ1WbbkBGVy9quvqVadZ4kcBtVKBHE17omOyrcOCYr9+zQ8KvFg
UQphyj1fQDhyFiY87HNT+DDPaC7oAxqNdBznbrbrS1DKdl9kLPgJIP9s2A5n1S8JaFa0dNLCUOl9
3POInjyMTzQi3Td0y0E4w/PYzWyVpTDOInuFcJS0u0d+nFdRKr3Wj1hZdCK2sDZnl8vGQExycehX
exxctPswZPq666xZPyZefh+AHWxoJhT1B8R+xS8MAvYAskCq4VTe7DbVKyOOtJYQdd82rZPMxCs4
gyL8P+g5Z6jkk4QEH2+g68LYLLHd5nSZvqBJu2yUjoc2+k+5A1CHmaUAUMLIhnyijzkX+TPRqLI9
JRGLeZk3vlzH7ntG1L91TjhRMZev0Vr7+5leUBVXhkPzWtVZ4B2XdfPoTkdVJQpOrJr5nglzs5vV
6aemaSIQPM+YBjlx3VAAPOei6T0tJIhwLGNWglKpM9+7u4h6LF33bzPoBBowwAbYTOMSQvN30Jr0
RqqwvflRxrqVQFwvSZx42rr33sOFZM75V/KTlSR7hqy6MG7txeZkFJZcBZlciaBKnpM5Gju6j25c
orWRi0wRe+roTnMOISC/8esyV6e+HXjGLPM/bVzDjIahCfFpDaf6ZG26FTwZX/Mpl5Gu4qlUWF8p
REtNVhlfmyjSGnSJB+zQtstgkO8XOWnh3/IQdtsdKVm989zS4td3kezLgwEr7tydHfUV3IBmF59f
Catdowfp0YD0kM1J2gi9m0Z/B7krtGQPm4ra/Xbv2mtjYxJHUoWqXENO4FR6NvZ/O6NVBywCAyXr
m9DozyrDwAG2QStXBZvqR9bRCBBor8WoGek7qgKUqgHIDoF4Ernv4VJTZcx45gcuXRvrXJAhXgBC
A/WwybqhT4kd8oVn+2b/hbcLnx7PDNeeT0Ijh+EX+twbYTBBdew6lmZV4F3VD0je6mLE1uAGLTy0
aZusb2iWUpnp/nwg1J2Vt8b7stVHMHBK82V+gpi1duWgVR1cC8SDbOdoUWBzJ7BYe5PnpH5UVZFH
GvJCA0fipvFBFF/6CaBU512whoX4UsG2InVuOUxMOPoSuJtxY1GYSsiGfR6u0GETMdBPUpqTvRfC
AzrHri/6mulSa+XnJ9CtVbLGiztd3LjJEZU49Uxy1hRIT3aObMqa6fx8601fQFQjDaVNc8zA5/Xj
bzYvjTzEzey5y1mY70bVsrTroTnAG0m0TtUzNdEc1MKqvHTxFhp2OQTDf/ZdDwffWVo+xKc2UWGH
Urtsw+qjozaLo9TGbVBzt4TQLJ2KuReGNY6fBMQE6zThirqWkYUXRAj0eY46Gk0FHpeQnKHPR3zZ
ErIZ1dDsq19lw54OrLP2rIa5TMao2Dn4724EmErdTj1066TGPeeTvT2sxe5Q6CwjI+l0Enle+6EP
CnFV1wLGOCWRZh+kT2On2DWeNRqtrmlM/yXXkrkYXVf46TR4lWqqh5NlCVklOgf4qjLv/crNipAn
1XodXmOZL4bHm6Gx4ZclbNnCazZDo/iPgJmjjnw4TL70CAyzWZStn6oxUzar+BhkOQyYBFz/7WIs
09m9Kk8rab3hpdJRsPysCIhzyzevMzX3orm8wsScbGXDMS05igEk5LOLPwFLF+PtNxYTzxai/s6M
rgi7azwhv05J+f+Ub78RG4SULYacfzwpwBAbGL4hJnDRw6ebgz30jhS+nqvHuAtrUozw9cctzd3v
Cwj2XkLhwp6dnPT29ODwUWukuohN6b3tSNgB1lRBdvJ4zrsrFvyJ4bUfsJ47wwdHTndH1rHeoeEM
rZ+7E7syUna95JA3ocqjEy0wDGFldgIs+t5aOVqkT5Z8ihYeoAoNHBNK0Si0rmveSRWzdiefeOTk
ZFCZffJcWtEJGPNH/LczX6ee8rkUkHkmWHMoW2Q9uhkHGvtcoNMHIEhLAvsmwYwbQUMDfZKXg26d
s1jBEm31qk6YxJNu3cS95Awkm7/MVI4QCjp6aM8mlKA5/xG29LJVclorDzCxn8lvaYwHlcHTmubM
xumq5BKVeC4ipTYg4Qu0MUaH/hAJ6f+DJzK4hkbIORf8oisFuNPvRRgvz33hYXHMTMfWpg3gluiJ
9hz1ZoxuCDsQS8u/KwOWRL/ma9siRxbBtfQoa1kUBft1mppQJcED+2vZLen2FAGIIITZ36h6SLl7
zAxTtBHtdr46eYVppIqIhDfUvELR/L7baA7/bu1Xiwh7vqa5Vpj1Giy89ajTQqKXeKpkqObMPj2A
ZOXFmcgTLRM+Zl3JeFVSEuKOrCJZUYNU4F5URnLKRdU5iz4vt3Yjybpm5HyJ6ogv0ujIutK1ki5T
/iC3kURmAk29QgWumThEpeVPfMIAVjE2fzV5CPc5n2QTmAoc4WeFc5qFnr8Es4qPbsexBEsX8UPk
dXIpNaxmne4L6M4Bkp7Y4r29rFAcKJGkwzDILpLJu28hju5O7ZbZdpBg1sXBO6GqRLcerkL4fSOK
PPVPnFU74/pKbvfYwJ6gRP4LWPl9nh/J92UpfNbT0bPL4Sg3j0i1WtENQA+zAW9vWfwCmAifIU+J
eMemJHsS3Bafk7EtK4w355znI+EplgyPY01i8VhIevwOuNaOp7wZ7wdMzLF0p9P8LCTBMdqzTZ7e
oWDoRZI/4GjyQzpVLnLCndEsikA0QT2a6B7inLLFJnAUPpVIAIe5Br7Axc+opA2z5lGuX8eK4/UC
cjrymZDAaXrzvNSqzra0tdn3nTERJttPOP++CDqa1u6IDWhZUZHm4wJHZ+XFBotk0JiCI8u0ICaU
TJRG4bu0Im5X3RWqXaGM3FkfeosYInp0P1p1BCwmr8tFHT/zrvMrJSWI5PW4t26qPiyFTdTc1Lcr
CVzyH1tZSAsd6hEX9lxTaQ+hyyCLmQV+5QjFNbp3p0xWNmBzcto3f4l56bqnQsJSn4yHFnX+S8va
rMVlfh5lhj84WlQe9W2Rrzx69chKHbfEiSJZjy3BRWF1exupGtour/IZoTHbaSh5BzwOgz+WRzLx
d+BVaCes7/5PtQqMix+ndPA0/F3gXCN8lPb9my8blxZdtFTxaex089RQylZefGQRCLm/3jO78a1C
DhUw15+vF7pDLGpSEnKqfvadbJg74QF/wvuvNrohz29jycIdDOjk2QRvEt6TU4WH6p5549nHyEF8
aXjQQtKAgxzi89UYawt/onEGEwBR/XJTiKaP3t/DYB+mTIgxn6ABbyEO148GIsvHv22c4RB2EUyP
nUOTQ8SKOl0wsMgOnCtJz8q6Gfv8FoH6G4M876g6+Z1nlxKI7/KGZfVitM/e9Z/9LlKW7wat2c1t
XofYcu2VToedTrBZF5XJ8cXf7kIpDp30F21fHYc/P8K60y6CiuXlVo+LLajgNCsL20kxS/iicSzO
DNhWAIbqlARKtidL4ver5SIKY49GChep68POYCQXWNszNku+PbThJTiIBLnW20Nr2guSkkkzlpO7
p5UpbWneFhc6ONGoBbNm0Ibi/KC5UZsnYpdKadae0N6dZxdE0J+5SLGndpkMO0G91RmgXJQYzXhr
RNat9naMNcRQcwZ5arlSQNHu+tknQN8F28naM+nc2fYqyH5t9o+0WtRderQIXJcDRCaWwfGCv3xo
eQ+asWlP5yv5M+Vm7XBZzPA/HToUdmYEsE942HaUMapVIUNij8MhHgY2HOi3GOzdao3yv/+6w102
XQfEjvJ649gQ1r536p2WuSpsusBZHbkfFclX2rRR0+VejSVSszwdJvg3yWf4LYD4Ywk8HlHBRJOW
khhgzP0QS+g5Vwe2kK+U+6IPtJV+kaeWvWUr91AmmSOtWb8AaMbpxbX8Eyn6KuQR4Wf25LGOAWwc
qYqlR6yozHpqgiTy8Kbq44JGoL6E3qw9HuB6BFPauCGpsom6iobn1gj4mhdXyLu3surG7baD9dSK
9LAlRNamtLrpD+OlnLsc0aw6jtqiqND+ujTXzjv2VzLC8Xp2bOeBqeKlmawQ8UWSi/jaMLB/znQI
zwlH/ZJbkow4ld7yTAdJZiqRObhJS3UUCiVzg4k+lz2ceHH5puq27KTQGC3MscHEWNnMagoET3BU
IYab3c1pxjSq4xMEMwSNjc7oNBKauyaL100g1q5s4fJA75CD2kM3k9q11fcoEbYb4fJ6ic4qHOjT
Akk+6+wdJrmKg7wrVpiz0BE7JUoYdQS+DVZxZb4tmD5nVWpMY80Wml9wVCe0lrmzz0eApwN8OhCU
PPPZAzTbmLGe3UGOanAN36KGZnIKK4Ry8tXJyCvje2lc+4HuD8USmfHvj60PxYG+pgTFGbm6sjKs
LynmYeh/2F8QERUs6pA14g+cgpiKHR6kk8QKeJFCV1XLteYjIGvaSTME2tLEdiWXzVVgT1u1vBEi
om0OUypsyhyMS0cB5Qh0Jjh+aimWSj8IYUWtb7Or3ADtwq6n9QOb/R9mGBE37+YrNvzxHMJzVDW5
pIs1ON7WmJQ/qRJ0s2diVriFkxL1uDXNZ8woZPELnr8/pYziHYo9e7XQ4bBhGaNJhoUKka8B5pKA
R2atrjzr1VxfC0yxvz1IqdWdkrgrCxUcngyHlJ2iS07D18c8U2tW1peUQBkghgBFLmytXtz76XAM
FLkz9OJG1k9iO9PxfDC89pKSkPUYnUzqWoWRtsmlRwsgqjlaM9PgiBQTLq26dtqAEJVMHtpx8oqO
/Pk4f+M/lEMnBPZcuZo8C2dI9gn7HJh9OM5C9zLlwEIY2cXIkmuPiu7rybELLaa5/TN67N0+qD39
5IB121i4nOTwImtTqBJ8Jg/PbzB8piaA2y9/pPUXR6u/9FCVHiWXYYhaj5d7GBPTTj+Vs6btNp6S
zgYJrpSJrUMBH2Ea9F4eWgPP2UgVs2UZQVg0Tn3m3cyqnMaDT0fjByQ3V8sJpFWW3zTeLnMSz1OG
9wOkwQIJu0Ue1l9laaSqapWk8mXMA6VDoIOSSrUolqYyVDJIZyQQSZFmL1H3mNM2/9pHeNt8q5/+
JzgGeH4BHuuMJ9pZjmN+XL/ExeLg+S88OscjjelUEmWeRwKLGblc6yWi9DQhM0JCV1/h1qkTisVA
Dn/K3MmVKRwAmG+PU2FTcUD7DYrdE3KZftQtvBBrJq3wPm9aVYaut+3TdQBenz0fH7JgYATHNF1Y
D/dagWoXtYfoy7GEi1sWcGH4aC6am/UmjipWhhPmDOSdLJHpFmvEJWQ7A2CUG2fWEXWWYWBt2JYf
zbiqvcTcMrlCu6G5sykw3go3pX64lGWQIuBMpcm3EDXeHYQ/wkH41HzGMM1UDWrvQFshyFcss9sq
80UjkpiF+llNhcBqZTX+QPw1ZAtp5kvPYTgKzVzX0sG/hPCnFyRWSTnKf99zIdkU/2+EXWPpNJE1
EfyiJOj+PX4lm4RafRwYzPZVsRfYaZfnU5SstRvfnh4aYIx0XH23szNh5QNCLqHY6Rgb8waW4xEV
MWo7Rw6prElpes85Lw7iR1uurRSJaMkBhS3wtWxiIDsNePhUtxLDt0yxT7aFQL9zNBdFhc4TlkPd
S4L00tLv3c4tsiJeclvgAtuX4mlDaSl6nw6kqAie0HdUpYH4l3rD/v0gk23fj6mvVaE1CKWjoKgJ
W1mOEAjUUhpoOCSX+c1xBa7z+1K8aieFxvDKO3iSrCM3aOwEH5aKxZnUJ/gIE4YM3GvpPRAoJ8Lb
Tsl/yh16s6tc5l3o+smcAnY95xuNrEYZc4RLnwKPuccDt+lBvm04dz9nYqK5+UK6aQYpDqim5Enk
T0Lq3iqv2mfgu7+TYGp1MyEPVXMOlef6nWLfdl3Hxm4EFCw3ofedjPxGDnge6GwJjX72JF/tHOW5
zEqT4qWRE1ML6nyz5n5c6os3T+VF35y4v0d1Ur2477bI4dQIvO+XYfbYc4scmP11GeFF403rmoPK
725+2tJXFCTerYDXs5woyJg8HjkDdv/+5xLmDY/VDn9oJSXxUOguzyG0Sjab62PF8EcXcvpoRXkJ
yTT510y/8f+nnhyvIlqR4pFBneQ4InTR5WDbEEzlv2agzggadBBJ6hG5RQK2Wxv73XtfhQ/kth60
xZPvS7y7cHti0kd7CCmUb/Qe1NqTQ0wwxaYqQ1FrSKgUfcV6ntsCm6EnpUGALjKvoWx3gdvrzzq2
GjOyf3qIGo8r4nV6sWOT+At8sIBxm1ROiU/6S4wEjys2rhpKvg5RZTNAeE2YhpjdP5sMkDlafw2j
MfAZdHHk/VaYTG8SfxLAmEPQSfLqa9nF9KGExpD2yeDAgi+8k44zVlKSVRmAqS6XbQfbss8B7zLg
t1GHa+iX/7T1OT0wTfUo2QnAClBrf15uqVM8LaPuETDwI1HdBFgLqYMNOo0HAsbJmkvXf3Caem23
zXihsoR5/+t6+lb0FbJMCT+6mQZvDH/vf4UpxmCHVjeb60FGHVgSKq+uOP0WOgzXMweu+3e2FEyE
HHoxVFz6yuhayNp+0uj10Bc4hY+l87oamuXR4Oc1qi6M34AmfaKHTnyFDMh4eIRl274JapTnQ5/6
6X/8HM0N3ZCFN0dMIUABsOroCfH587n7+tDl5v2J5WrqucBdoW+t5+NWNmpL6gHg0aDWHaiIj4N6
PUmlJqNsLuTjyNQnGIgoe8ZSkp3he8XKEcR/1Zbck6CrS24DbPygvDARaFlx88LVXSi84zHZiAAK
1zXTCWY+HFtYNSWLm9SQ1D9UI87p3mrU18Ymyls0fltwnwMUeER1lRrWmV8hNEZ+AVQYWXjELD1O
ioQ9NZdKJZo7Z67le44tpJ7i/IfnYZzC0TKSoruBnd8OQ8HfY1UPqTyiDVLa1wRUfeJ2n4vPR/9/
Uvtg+lImVfQAa1cphLPieBrDRMV2IhUNJkhlwCB9VVZiB2KXLGX1SN1tLLKn/k8q217WroGj2Js8
ugtoL0nTL1kjlJEK5xFEhF0tHXc7bJzWW7vkRexAOnnCQcDBvXxYYMqadF/5R1Ot1FTJaCSynSjn
GSX9w2+M8uhVrN9awTXYCwaRbrIPx7USq77eWDiwpSdiwBove0WX3nOpSQ35vHH5kgHoMf3h5YtS
0cWOmgbDbjdpNjGKlnEffhhP2Ik4WkDwNY2tR1DYSNmjTdD92R+GokooRjPRjIlj/twu/8/CsWrq
lzvV2kWageQl6EfmRc9b5f5WdmcJClFxABlKYRMKauvmkEYdVj2RnOPQLHxj14QodKidX9y58jic
ShTdczbDy9nRneqUy1r01utznLUil+iLrFFHjl9bJEfbQ/QCmUuFXtJNEw1+I6xDsJbZMUtoV3SK
dviRsXrmIqSBl0ck50nL0LXYY8KEtQTqhV+eP3Ik+sHLfrCQpY2+mQoao1xH0xUvWcHumG9/GGRp
C+h/5n4NZPj1KzD+IRkfTgRaFcYITEp779RoyVW6N9MxZ3cQ1jSDC7dQDgQHaisO2u+YPzm2Uo+e
LdNGsv/FoPNiK3ukTvq2viXKbHhjK8OBYzNqNrFd4HpdZ/WezobORtyeTlWJYq6Gc7Tj/pXUXKzb
4Ypew2yjH12hUrJjHHA5TjkHsT4vxMp1GXPdDt3dcjLNQMWUc5Yj/sWqW7qYWz4AqdqrsLoQjP8X
/xmGqYvqXGmT5CXJoKmNdY0he7cygR+dfKlhJsQvMDl5n8hCwY1fhi9CAajz9ExOJrebTcn/gIcb
hHYFvvTZiEczHdGnaXetK4hQEKHegR+Rx8Juvzol2zHs9reEKrOHvtygG/Hgl143ZnTXI5eLsZ1S
boD2cwAGa7J8GnAR5fNEY82/PWFY0LO5y+ehTMU2tD0DCgC7RfWRN52HBJA6BDt2sGX5QT2DFywL
GCLTpMdthXANCMyyniK4EfWW4DyctNYJT3Y4BsdGdPVlRgJv9tUf3al0AKfqU2eWoQkNUWLKVJzM
OAjo5HCAmr88T20hLaoZjiKmmPN8uni9S2rIvBgsgBgBXzYsog9LAdeDMNide+wTGdK44JFWB1ag
HwPSUlRYe9H3hO/MC8HvEfYi0lcQWADFN7eZPzD59pRR2ypGxhiCVCzewNW7/hfC+MwZf+Cp2iQi
F4l3gdZcRwUBjTGXYqKiFCwsrkmIGPaHYNX7PlgbLYjaqNaZZ0uaxA+L6yt4AwGbqff7gMiK3WvT
m46kOIo3tub0cO4oI0NyEff/jTRYQgHkyB3B35Y2v7bOOp4omX4o4fZz9ZfBeA36YZaNP575c3BQ
1xNYpM4zxB0vug3t+Z//21ydiQmV749+GC4FWLqi0/7cJ+KkCwgi8aEXKxZ1jjQJU/Ds3rG7ycog
JjWMSBs/kVw5tZkCRvLc5z8/OZjATPeQB6AS4HYHf6rnNMD5aSahFOCX9scF2QlcjVbp7rNQManb
zrZnjqxY4sPrh1qDllZWV7+FI88ykuJQJROCdKtgw8uiM3HrwdxASs/Mhad7fUptFx2FmZXwA83y
WpbNP3F//qy2W9sHDuzMuc+epHbrgMGSXPgE4K4N3W/NJ5jBti4BxJ3UEDVCTMQL5hKdisf+xc/z
Wzq/a+pjvAseR74FzceZDADL6FTp8cmK4m8QtjYcx82jR9WwSfW1VHyoMozwo5m3ToBCvPAaMlHf
v22o9X1U9LlLPG/3p4fBH5gUaoGpucy7RY4iL+uY3Ab4JfnuMHEqCq8BsnkDuuNt+0j90Q7cn7ZD
Cvq6xM2p7BsEoqybPInv9CP/1XIqiBK8c1y9YVhyZZ5j+b2WSzi+AAKyXT4DSeNsRITWFErfqIYJ
l1YQfpjRyUQcXKfyzr2gDvghC9EBXVscbeGnLC12pymZlI3eeJkzk8y4yQ/dU7gHSv0uc91taSuy
2tdCZLgDWmsfK/U1GhU/B27oqDwh4MH+xwevNQ3lIee0R/dK5SssSsHzEKHuP1SEUD7pOalA4q5K
EpmOdNG4I4FLF5u6yhnwuoIv5AwgtEbwOrx/JbBimtDZL5xOHL6EZygFOcNPPO4M0GJTWlson9wK
2YUeW1qXBGC7WPfhOK5+xIPCHADE+wz82O/jRIV0aS+hBsJdQph2aDkxGdu6l4p1S9Zc42s8sEUw
aDVbqIN5xkY2NNSmHGpeoGfK4/SPisk42P/81C3q2/y8o23Fya4VgMT1uSKFwev7uUbgDteZWq5b
L4Ieo6VLgclR14/9vdaTyGxJk2iwJ9dLEjR7StNMRGZZ+4D/SB5z7BH8KuKLM5iev/mLoq+/BxHe
1s+Okp02MRv3vXX4LsFhtLFE4czBFEJ2Ec8ZkqtqImHAU7zc/R6tgZUg2We9X0InwuPG/hxSTpMF
a5smnHkUEGbYZywSasYs56UCxD+bswE0YhlZ/N4ulDJ/kD4xkdvC4RN0vNPkdk4gkaLfuprqvIL1
C9SKMHiQGCZbjhHOz/CQ/4LKzCmfMXjbDz4K0POpdapcHNfWF2LVPlcih6B9o7lpsu7nDgeRZeiJ
BGXT+nb2jHLY9rTVyO3zSxx0zjG5VQKRwTLLSRzOK9yO9YsXSGJtD4BYl/stOwHNofj/S+dgnY5m
k8FDQ1IhtzbVqdL9Qkw4Jtm2px3LpIGL3/AlnqD8A51GOWxNfOQSGs75MBJB+n1gbsl0+AGXUY65
e1KK1clK8gynyHqo2GtaaiXvAGzd4KMPP+il4O+NcHg24WIjWYiIYfzrBRnfCA7w1zqwUGgf8Uev
vCKgm09vMxrTuIhW2AfGL45CAjsyJVfCdRQZR8DvipfKX2cA7kiK6hMc60dQhETvwzYkKzvPifjG
bI5Kezhd6bMTWFRcZEqTwV/eSjJbmGsGfH+NJoikNcFcv8fOWamVQ8kG17XBZee4OLbMqFp72tb1
gdLkVidEAEMsbZfNRJwHySs/4hxIjPwFesUoOZ0Jm40N5nfkO/73AIp0AEkgtoj0F8/LvSVgrw62
t/L7gOcgXYDHfd0ucxpWk0k40phlO1NtR2DxtpA9BrwNdIZt8nFQF5C8tsA/aHK2DU3K94ay1IfN
X32jqNa3VPPYa5UDm3SV9BYYctzMPl//mrXKGL92koUwe7epTBdoC+hOYCptJVwJV8DbZ/t8aQFs
MQ1vlcikoJnhYeW8anx5egShtNn6fiYiZ70JSk5kL3cphWc5QT8m1Gc5SGFIvk2x8Cwqc8Qg+IjG
ybeBrM3EjyOzoBijiQaxgUGuy3G3XuC28kGDkz2mPdSyY0OXEF2qBfjlO3HX0P6HGPJtYGlWlWj8
pGXOJIBsG0BrpLa7sUcWZ8MtoLLonJVpr0V+zOcYlWKCExyyaeKcdorZu2PFmMKcxHX98fhTMu28
22vpsqeTchBfi5rU+aruZbGLOcjdlivZLcq+hRzKHC3am0O7y9cDEgOvhrIssavWI9U+rQKZOU/F
glM7ZLP5YOuHgLlTWX+kCFpGGZSn4ImkoUQTZ1MJVo2f/osKV0wHbNMRvaiwLVvq7zgZz6pXB1DR
270n8Nip9xuWQ8mgLIKMmRJfNKmWl/uIw5OOwSn1OBdu5t7ld6m3Fd3C/+FR+pomeuc9xCpZ5NEl
OkX/LBmj5R/BbV7RtLf0oj5ypSZ1lFupg8sOX30E8WlvoF5S70yoP/QlgUWjujVaOQ2KRPo7TefI
o6HKu2ULY+s/X7o8Gu+XOLmaBldHecsFUDql0xmicnmRl8WJoCaBLEcD3pwGh1LnqQFh5nAJCVCg
G0daH295VY7VX3VV403sudbV0KFAcgGLJT/La44H2a6HD8n1oh+3yQ2UGOn1SRwHDyBQWru49XBJ
vJ2Fd1BOn0Np9pgxle1Z1Kpe5LL1gyoKcQCavzlGdtSwzC8ahq6np/T2HUwR7Mo/ypOctBSAoRH9
gGj5eprOAbJFIYcdplTdAlLrXNBUVa774SDj4w3l69I8JgUv6XB9VfV5hrXfxilDCsu+Lp1WQuJX
oBx7Tz0mqfHx1HnbseZb3CA4yW/r67CRw82O1U/DLJWUPMOwrSkFa629ABevX8DSy6ABqnaFhc0u
SSZQOMAX9EitVGEtpzHrxHUnvz6eV6tieSXPpQUgj4FbRfpGgmQTaO8Dr71Nykr1Yb5R42/+tfId
i98xW9HSTBlsO60BHE74rOpXlFTVwgmAR8HU/Cm8JrCkPzddNSrPR/MTYIxJZRjkU9tka6px8Lg0
MkwpUgzaOK6+ltz9QohqQ3XyF/9Zb1Rr+a+cz1UchM05Ac1YJd1TSIRDWzAXI1ybP6rCzuM1uwSX
F1ZMd4OC3t2hjAEkQa9A3JkUwlpy2slkoxqrh0AF2Qa+/OCdwe1Bb08RQpPeiXC2qP9iLnh0eQ5+
dyebCtITUR2nUwNXrUElgjwL4IC9+AZ4cYwodvAQMVI6+cx5pViwgzA1+yvxrm4bKvd6IIyAttYU
hlVr8Mw9rszSPks1MS0qDtgB3+6s+jkQuXC2a9IolRNo6jMdm3EbZ3muF5XYMVpb8dDbfHEnGGfS
je0J0MibsyyBYCxSewZTlNEwDf+LYLt8DmfAIWFSBnlvx/J4RU/vGogY0ub7UE/wZZyKo63Pkwua
tkQxZHaUV4+Sp5fSmz/drl0vqPYV5ycISlAb8fLirA87MeDaJErC7LWeykX9oazO8I7yxkohQHCS
E2fgLb7Lxz0Ya/4YJlXMqlI8D9bShDTvC/XGW3sDowbjxm1dLvGIZvb1X+9+7n39xcIeGPH8SJHX
qpKeyTID6FtjFWWcWajXFrtsHJHdSxm+CRpcFRxYte/5049KCrJPf+Y/ivCB1KBUb+xULew0Xhw2
5iPl01EvGAFE3VckOGwFcD1yj0K/mKjFsq6EagNDAx57NlQjNvEzfOdA2tw566JtNhTw/BNWaO8E
/pOKFJtfGbX1043MYFC9bgEYUX1A9vA6z1DG4jciSPN2080dHhD0XQJfnKa4SQNVDdUQsoW9qBIZ
z/sDuCkCvxdDwGZdQi3+sqvwY0tp+EM2bWEcyV23LjMTqLtd8MOLqukafrRMt3CQni7/59ayS0VY
R3zR/jAjGt6dSzrVE6QtXgAcWPcwx0r61+nNI2nzg/SRCMMvWyRxkix8G+bg6eU2qDGgwtQKzC8r
KLSQ/No87msWLTRdSUaFFPVwTszad3FDCWjqKo1RryIKEQ+xLtHcsEv8qyt5T+sWG9Wt/ZCOtIF/
l4KZq7fNcfZhczXssEO1GsuCdSjw6g4eD4Oapp7gKGc+Nh3apdHCdqSQEP84zl2oj2RszFDmZTE8
kM65kILloBa8PbjhEYJpmrbsMwPmCQex2JkErgqY7adLI+6w1MAmqgn6DUNpmvv/ZDXl2oqnczkT
l1AvWFIYE0duu5Xn/y1SepcEzhGyjop+o8gWeXAchCTuUKpD/EP3dSs5j8yo03ZsqJwehslqCwfh
vt9yTrKzDjjMS6EvTPdVZCV3KXsluhLe880HnuDS2iQO6Nv/fEaVc0ArqkUkRj3pxVjMY7kyy1Fa
iJKsu8c7rcjfL7szvYDGb4UBLi/TV1PnTVBCOZB9XcbHxETJw/lUGux2KJVwOLUNcm2lsarAMYP0
WLPxKWnfn9gft0sWw8/u02f+5ToScEupZF4lHzg53264ULVXlKpuYDglYY9Ce0nNY6dkGl8c62X1
W4kTA1e0OnFyaGv5rLCxwWS01VmNGq6vD6iZHxnEBn/peYcN3sOWbU9lyhbXImDF+idBGpwqbimy
Iwoh6SBPrJGnRbRBDtaEbpBU97qNhA2TGy7ggqY4y+KeEcb3o9gN5JlWt7QLKSXfcPW8nD9Fnrn8
SVTsIcbJ1IBeVVMacJm13xsP2sFvZQplRT9PiALG/xfXVgwCNWlpdH75YsEgx/khAWoihJEb94Qf
GgSKzivGTi7BeB8vXm1clUBtvZxpz8tlO9AwTgvTyj3H5ooSfTGzOvs/0SiZdUQs+ajCEGe4CKCO
i6ugt+R4FjBA/1mKFjAWW6KxfQhwawv7M88e5GDlMs9LdqT9qGkgSEXgk8Ln9QRNVXo52TW7mW9g
SEuLXwkbVfg1vb/pYU3KV1ByIcZUdKlpI///gg8lNZN9u4wOQRJjI8zHK/mWiAKfJNQcdEGHoTrF
EDEKXyxCBs6bNXC9EoNjDI5NKhR82im1COd32nFnzD7s84x0qe+uX+BNteJCdsjYD4GoN8LRCZIB
R9ZKRCjywbp2ETsp8PMuvbALU7fofHhtk1XsfZQgnX0PDblK8W5uqv7ITLwRvDYkmlV/zJXyojWS
0fMxoZuliUo/F4up2q9kXXPjguf4PJpadi6vZyqV8q1W5rnshM1mr7Rz/6xjfMvkkh8olmoXOy1d
QijHm6fdJ2o83xdtdNeoJp+Ed3W+EasRhnHRUN/EMRhCRP/bUAtWb8Lr67Af4+euGBj7U756rqc6
uBBHwPdEnOa/T8wc0NGcHbDtp+3pe8MxaWaMztg3Kg08Pe6ENP/xG8XHTkpLkgImpLJl4y8flBgM
oWGimpHnWQhVdJ8UOhvMMor40Q7+jvijvsXtV+0Q0UaiYiV/bw5zoWJ7GBVmVv7MZmappSdcA3Ib
76xT8dhasH0RV7xDk5uRHxlgjdqHy3kOW9urvPyB1tixXafETxC50znC/t6CVrp+a/N9jH4lx/oL
/P8EV3n3FismilFu3K6Gi8k91o+Y7hkHodgQ2FT04Qk6g6FclC8H71gLLgh0d1dhH6l2WPLErzep
wiTCZTwdefnNSK10WIhguThfc7TRR7QVhwhoXdiDTnAQ64o6U1D3bD3/TobsTwMMMIqC62z5RS6Z
8/8FKZ04siFGoyD32/Sp45Nz0VsdP3R/v1IqXcIMc1zwSG5tNMZfnWVInxs4+k60wOn7+vsN6fcZ
B5No+UFVaYi3o3Nw1Qk9p+lUALGbrrJPG6Uiha54tqL4U9gvwsKRnjClPTytLaBpTd9veeOby8oW
+o0JJStKoDlKJtQnuMTgI/BrVaxYd0MHFqAx6YJ3VQAeJPAPLu/tV2hQeUSwZvhilGb/9riobzfM
BTgDBSjZ0Bzt0h0EBf/ZrmN599Gd3qj+smTh+Svz5q2KbgXC/MEWc/iem8HXIq77EkEM4fEP/fq5
7hPlPEObGQwD4rPPVcrVp7EaJ9NBwqM+INDzCuIp6F0R043PibmKKglZHtzgY2pW/YBkRR1wVz37
G6PU7Ny76tkpGT9t1XWTPE360ZplQsskZMvkFA7jrrOiqpqoA7oM8HHLED3sHHELSsk8P3L6ccrB
wpbUmagTe122kGhIw6nUlPhy6B04C+fcO8KuBbgeolng8vmUFwetlPHumkMZ2yZDNfoa+Z0lCkfU
RJPRW7IXUMAEvgwlze1EuNkBsFwuWyTMY5IrrJBawlnVpSobLPcLAJcOuW23QdUEiDlpDDxIA+ri
aQ2uM3ZFH6s2q2btoEiAR2WX27Y44YsD6F3I/d8IVD8sspfvxhQoLXZ7HCzXINzfei3qgE6kvrUs
XmhA/4z4BcVL5MKxSkkhT7qRjRK9n4EBLqsoenxw8X8OciYugi86Sv/ugEIQDazp9pulxLgDLBxT
4BEVXBeu4hdmI8hWGC3Atls4IryUl6Wz9T4eVAH0PEVkZQtsYq85Kave+xMd+TZv6UJPleVULMkV
7lhQ/C/Vy+JGOWx4VHsa13WhlRBNancxHxQZNVee+qqCHOd/9/zUmRDopmuwV9hPb2u5IQcMfEaW
0M9n++L6OSrighY/vCUaOqjM6PwlY47txRUjCxJtH1CJdP8M1/IgBIkt82o9Q8KvE7Uj1ltY+hhg
FsX7NcLHjkRs8XFJy9CBC0FWCYRPmyGGcQZNCSzzruYbyrbqEzhatDZyjAqP5bb5N9lXsoaWp94E
H41C9zvAfT5+ib3F6tYuvfqQpugFWQfeC2K+QPFug9Swth5u2narDZHAg4JsWm7qFZ5bzdydAfMt
4chFSdd81iVtCRkW6LA8GKlloBi7zLG5U3gDBAC8zhL9UNWSCKP5cFG7hbWUEUleG28slB6MJBWt
ZvC4qV27dr+l3ix/Q07X8l2gbstrYHZxM3FpVOi5IBunBbWtzgiZwbJWKaOpbGjM+EWc04ed5Y3/
HAW11cwYCiTgm2fl8wuZtovWWLwKz9ygF99JF2lnF3L8AXR+J6Fk0KiyMU8jfAbVx1GwvhQYH5dC
DuAXM3oa/YXGQ6BysRyQ+mk8uOnDPvW35UdqEnC87W4G6yHLY9lvp3kXa/vFjU5w/4eQN7eRL6kW
hfOdWHQdVplQ5n+pBdbEO5uMt+PG8FTwwcT64SDFkfGE5YQkiAdRRhO6+PAEgm+Up8EHoRngA6gy
dVOULwPjAnFW2ld8Zh0lUqlEZRmIuvnfK/OMlr6PhKzjTKs46ZY22ofc1erBDJhNT2CiR+gHVhoS
ReZ2IWtqKMvrVJSWgLR7+//jkIx3rRogNTPXhDvPpeAQ4UZPVW0AlvTIvHs/kKsAbwTJPwnWY4z4
+XWGoGrDglLGijwqqim0pK2DQT656qR7fsEFZGlttFFMmK7TDvQQjKG9rRJT7pE5qVEK2PiWzaNL
Ii2e4CB94USb56D4oLjEmzJTOII26PPC6VLsa20eF1S1cnb3SceS/bwwA/V9ZTNKUZ/y2RP28vLK
acrJUMr3qsGgoprs2wcmpieieooaFjxW786qJRH/BUMfIuKkyHn//8Z+/KZYsaUGFf/DcVHHQTIg
iX/Hf6n5zXBcbPm7n3hCxlf2P/Xh2g0ju6KWPS1E304xja7fUIpW3CxuENqrON7z69+BwF/3PiMs
1zkpukN8sq6Wqd5DkHJhHW5FPFzYdYWFpBN0ZmPN8vQmm5JV2L80smynRn7XNzDshKzm8+NMsvs/
uVp0PWA5qXy3g+7mGG5WYkrB25ruZiGiekPQnv024i8I6DUlQhH3xrz0NyXwRyNroJwk9rVWggpI
HfUG2kEEDEL9ZECAJEeDf+DBqciR6gg7Ai97F4VE/Lij7zqojwlDgUTsHZ9vMsqKI35DqqlgZMWV
Rx+fG3owXtIVFDzznIiJoMBaj0FBuHRV4KYsjTU9UjXrvOomdGjeQoIQNwg2PM94Ay0C2QobI3O+
ig7jvshonZRATvpbgUWULeea3R3JQf0MwPwHw9F3u5VjB9lZQB7GRW3w0ieAk5u/60SPvAaC31cB
OKuWRGYEjnferXmfiGYC1ty360Nq0/MJmK9CcJ3IJbeuDVo1J1KnVOmMDDWop/Ja/o42sntz2lce
mfuQt5/eJdPt9KBK5ToA5H9zJGW5IYixQqxytRl5HAtUS4HidvngSamWH97Zi8olZkZm28SeQ8gg
/QkL09xhwP3CtErnfHdSmWWOeOFCkt6q9rzmiXTf58GqO9ePyqtVkoUbS4j048j+l4US3uETNG5X
LvHTtxgnneuTUVvaiVq7wlEOmbltYrihcpROVe/6kunYC6PvWfH3GX/RcKGXT+7jIH/YTsOpCXvC
7pWzjDREF4uPL5BrOI0vZdIt03xMF4O8YVbQEeAq9FPMnk9sOt2uEO8fIwVW7l1k9kbuJWgP1is6
NIJN40/+MwH4RllWz9ZhlVUyv3yJAdU1zrbbWRBYQ8kyk1E9Y35tAcyrknvGUwi0+tD4t+PqwnYu
XTknHG0kEhMc9aCjWkJhUT+7rxDziHez/hNcf++1rlPrtRfS1eWkGjimLi8I5AU8xzXbhq5WyQIW
AUFUzrRKEIMdcZzBJsMuGoZS6pa5xYmV2/2KvT8hdTlGnmZn+LxBPIfckOh1lTSui7FzbmlwZ6OW
7maKArvi7PTpby+Nb1I2rzCiuzCqNxGg40D5+5zrMhy3B6mdps8IH6AM4vwIpsF9G/sNG6A0z4bF
URDaxLscO5iYhqS/VAudtXtgTbirDRB6c1CKDej4JkA2ZuM/RwtS93m6uDFbMGs3DJWjkYZLXFiP
I+12JxRi0cvEyTPfCwFwoEz1pE/ChNxEP84BoYaYhMXe3GP1oYw2a/k12wIdRtwLVmEGuw1HB6PX
8h50MxWiX8ogWIleis/3qBRRPVXSAU3fvOt3rjck2YJMopEOrwYNbG4cjjg2C9GryQ+bXE3sGWn7
h8rB4XEGwFO+xLg3TC/+SaVuTkV8M4H8pPSmyJCRjWdEzSjE8TQDbQbAnvcbDRh4aXOzlhxZUsGa
aVAKLzD+yaW1Bj0FsPBNWQE0uvoUAMNIgehU3+/TmY4PnsnHZ31uUliq41lx/MlWw3aelAHuQFrI
yNf6s7ivOYxIIZjcS/Nopr5Y5Bd50sQfrdKRj1sbZ60t6IQcyKHmF3z9WdeLJ2TWqnv9gZWx3ccR
52+U7zlxDPdxtGqHt3U9JhIGE3HQIdsQLvIDtTJws5LtbAkjtGTduy0t2U7DHpSc4cxRwOwruyeT
HY6HLDSgs/WVt9bVUbBMC2flpffI6MOpI/L3ZCPqWkzGM8WMPJ2gVFtB9m/8vRLaXgvzmVcOQb1J
IHqVG1crzsK2Fnf7EAqJWY6QheGYxtptH05dkIF/+v6U3AiGl0Eiw6/38Pq3cH/QitlU9wjVNmDs
nTbzpX/ZYqi717VQpXD4F04zStdLcOgUqPgNHNDAM25IzpJ8ukadhYC5kfCeWG/5Kt0uOR3+p2uV
ohVT7vPnNt3VO/gHwJNvhrcQY1wHRCXSDFabIWfMoWud7NfXtg+nerVMn1DHcT1WsaK4WUdcEOP+
Nii5M++ug7TGF8lCbHvCilDX11i25/EUbkLLfT+TN2iyycYjcXVa9Ni4J7m5H5PhXrDLlzlCaOMJ
aUngI2Q+dx5HGlNlFtjxs5tc5M6+facy6RLAIKDv+dsGRNGc4557bUkzkjAMiE+r35AqM4s4sDJ/
xxTO0OnqtR1wcnuA3Cd/GCYzB82vm2MKPRWC9UMjNm9EcIIUk4wDy/34XbgBAd7l3i3PMz9VzYaK
hGMw4aRM8qSz028eOGt8ntkiMvPk9fg/FMjWrciHMC3bIlulEkyzBoF8VM7uM8jJIm09eGulHns6
t6L4EbXiFN4A2bfCBEqJPahBeynpEcgCloDuAS2iLv6Y63QvgLp9UnX32qA3JWeHME5BxNEkwixx
yJrFpN0llNEMU4vC5P3F1Y4C1Ym39GSoMZeGIUCzOyOGvi09QTLyAKrbOCgsur2VvzS4RMOJWFkZ
qgK1YelGoFFEcJW3ymMiYAO63TSZaEwdvLA0kIqTFwPTHShAuqdCC2YDWPT4v2Ew4gE5uD0gkV0o
8LflrzSuJiV+dWs4bRAHNUydSrzEAuy2vCrVW9TJp5ts95gyTQx7DWcpi8rwKDPvwnXHZIBP9sk1
ikAAu4qYDpAUpkh1quL7SkAC62DmM9lk0Q49CrxKKN0KwlewIqu1mANZUJ+3KR/J0QZNY6DsXJ8d
kVNFOQ7hcFiM6vJQ5QkIlsm/tKIm9CeXscIJPvU3w+jvl+UY2z2TLbEBMZvQLC+n9hhRG31oLwAa
g8pVRngKIcmDXhc8XoCuAiL85je/vGFO5ffXtQaaujQJucs6UmLrRuSLpcJ4jK2Kp7QLr3gID8Fw
2ei85z2kJPV78edW21WjaA+eSEgALnp2+RPAVytM0J+au0bZXWjBaGmw7wWmOeIKNT1DUJ4yy/Pz
rGS+dJNYyRWuDt7cLj7nfNtiJTGVAWH6ij81C29Hzzl2sJQu/I4TEkRzUEqmShw09qG8NSOiHJBv
wXbvzMhEgbqJyApD+XT3tv2kAIt5BFZSIzgTLYqtBNheT1/qGBLA+Yyg/McZ9f84V+iJ9+loyPMr
9ynorhbNCFnvlYRMw8FfboKCwV2RPl2nPaVixWqG6fBYKrad7gL7qePN70wp4SSeE4OKNG2GrK8B
9EL8q5OV1mTXJsoItHa2JTQ6qeiUff+txz4x+SaBoEXT3EeGUYoPfF8bJre10mv88XghwBE/3NkW
I5ZvI+9H4tUCOPOpYgUX09BT85/VoaaLwcc/093i7JRMyXrA+C7muKGthYmjHNZ2cYNYJdkRh0kw
rVTF8/pcgHNgpOCjrmy+vrFhRxPiTJropQaRGadcEXTG7bBlSFaFN1W876ta0Pxpe5DOIEWFKdJC
tvGUMW83Oa8QDSF7onKFgC5OY4KaV79Q1n9Gqjt1unDX5HAezfo3WKCUObzNN0Cf04zABTfU2iPL
rK0HzTx8dzJGDpn+4TxFGhGoMq8vhWJeG2iMOJKdeuIjGrwHNt0T5E49/prYKkbpChY1nJVy6J3/
klwGaFrwpDNySPS8LphMsL03TrpTpVkbL7mgn7XmpQUZlvQcftIo+Sb5WbiGU7F6/S/6QQFtNTS2
M1ODTn677R9ErsTmqQANTRRLH6pwA/OH1dqgWXHQRIWn3Jw1xypgeP68la06Xvyld40uJkpwWSRC
sFDWcQdux/sg0YQE+tIAvg5/zL5AQyVJ7UCg3QdvTksnQcqVx+drv0IhjGIuBOrci3oUgtRB0K/7
DCGAg8JMHLMiqUVDRh68FNSwc6JXDp5bb/8f8eBHyWieYN8UNL1Lv52WGlTJD2Y2VVmGyO2m5hOX
F32hMjQQ6zQ1Vbp3Noiaq6Vsvgq5Wa3ei8F+9gvYnW2qJa04YKVUumui0rsoMq7oFjYoFmelSgi8
ptM8gIe8N4GL1zaxhsh6VTiBb4zePNvbWSikW1jVB1FRZpR34oCJIlh6eo92AWXN+i4zGq622P6k
jNbtIFXSpVQ5k/VGIoqzmtpbOrQ1rQHzYiHBzKe7oYDATIfiQyrnU8ESvrizChzV0QKFpzOTLJ1P
MP7G56EFtQNwiUt32Mk1zxRu2/+cOIOvqCs6YL+PSd9jMBsUq3tIRMYPLN39am43xW2EJ2Tuysto
ZaKQE3aSpzTqBKtzLbi9OVbZzsKLeVFdPbG1AE3RPspoQTqOa5QGqRD84msg6E3GAPQm4D4NileM
uDChvCE0MdXSdjrIFySUC+6a+Q/6DqG9O9icv7y6v7uWiIBrZY5nmQjqjd2qttoWqCelaTb2iWQT
dbozGFHLRqEQ7OOk7N7E0gBy1Is5jMqx1MkNoZuB2tZ+/QfFMDOQJuW5c2+IWlDatGApysA/h2/f
Q1/PeqX4KDm3RCqO5h9R/2S+G0s5I2W9IlLEyh0covxy+W05uwD9r4KUzmvUswTJElSFmtkb59B5
kbQYRhZwFpkocXHpt8opnM4Aw3wrNW1I12o48t2RHsYVywABc4qJ/AAKdh6OfZGbx83QMOW1DZPC
3YgX8QUH5Pyfyr0pAO52Gcx9JLVlNR7SxHv1rLlG1EcZXhALDaTFXZG6NUoIT6qRBR2GLh9YXK/5
BxKXSsd9nYS2ojwYSZEjLmvX3iMBfePEwgSqLvqIO6YnX7+jmz8iQcqf8CFofi2VNyPOTzzj9yTp
mloI2bhZh8No3kqpAWhRhAY5XcQXlLq0U6iqW5fE7WMrRNtFMyEzJuE1sxWSauXVilddlxSx8cd6
i7tMucd5Y1RljjDdyJPbjui30lhVhZ84wys1ESDIZ2Z5h4y3BFsa4zCt52wef0ujSonkT68iAH6g
1T9CmiFr9HGPKujjJ8WpKpjAqhs2tVCRunMOkXXIXdtvhFtCmmtwDVHvIa0N1u1XPe1wfCBpITos
sEJ8MqSsrCTDHScb7m4VF1oQgoaQe2VvbOauIQhP+L/xojHLWVNz3r1cIZ4eXEq0tvtMTQWKrm8B
Qkj2gdQzrl7udI9XNUuHKVNLbVdVqP3ZcDU3IZEcg28A4rP8BZvhRDFG75GDLP+H53siWNAb0Juv
m0whXssbN5lvEo46umOvCdPD1/8pSORXVqwJmPzNwqwmoYYoFeLg2k/JNe+nbtmFWzgVZ2gdekeR
u7LUhP+c8PmjGhnzeqYIDClWSjkxWi3dfzKD+ohrawBaQVB3+02BJrguw8Y7khIUEpIuWwLBap0T
M1RjCisgo7KXHJDpi/LdrIIpnfnZyVtUrQDlTafhoASegiTC1NH/9mzdyLTHlSilDIA1fW6OeRBI
TAC8huNhmwL/3sjqfJbibt4NGb9brX7iMggKKa1HgJejgisCul32ecxZgu7AzbSeFN1+tXBk0JIK
W488DW84jEvGeMA8yBxngR2r3F6vk+P2zL5+i2/CoSHucESwwInlYX+yFg7TZ44z/6ZSNA0/7fUA
VI9HkwHcmnVS/24Kh7TGTRKfRRkXjozwVZvkriiHpfSJ6sL4jbyXCqyLg1wK1Jq+jg6p+sszrqA7
CecEK6urN7BXWofnkgKFcxHWr+Ug2iT26hW6NPahmXsq/HpalOkVCVwZeqRmCH9qT+jKvHsskELz
Yr0+Nmlv5M770hjnDYyu4ATGy0cnZN76XxoerYHChK8EE8giirAeinj0a4WOW8nAivfnsFd/KplJ
Ql2jQ+yoeM3dNEFiPJtUV5Z8DJ+1aSml2ezh1CQaPJbfYIXNiXJhO/6eTnCPNvgExWH9w74NXfZA
fK/aLhmf4a8VwQ5TIwc64Dz9hTDSSGdq8A5bfdovs2ll9As4dzIOU2uqCixNbLl4LnhzeOEh8Hqs
YVbEpUGZXafZBJq7+26FNVqqxKB/J0c69sfT2iSWuTpv2B5mdcqU/JrtsHFyW55iMphpRhmlW+UA
R4EaKQ5Re1SVF3ORUd6C6hx6XxmN9v3j6/4UbKJISihkbTIyX/F39ZHPBzb5iovGy8GrI7cNQ6I+
F/G9hAytLCgKTYIqC9zbm/jzLSw6SNg8kOydwjbYEagL2W8HU+yQaItlfXi5O5qP15EU6Tp3E1m+
uYnw+yIIay7uhq4cmBUo+IhzTiXStQ7bpDCMCN8dgrfizRymwE72wmMH/f1Hm2PQ07caaNoqDvXR
ecmqXwC/gQwHpf7h8atQUusfh/hDMxQ7tbN87FtyXTm64vCU4J34kjWfxBUlygKnwB7KepQ0Zp3i
TitnnC1yq3ebCTh/N0PQCDR5+K09lqFA4KJNF9UNpAi4YV3IB36BQtUkuFRbIqfn69/l72ZVomVZ
WmIEPWvArcK5Q9Ocd6mPF8nkZACoEdka9fbxObPJpE8mT6ryloKk6TPrhMxIaW7uUf++PqgSn5UE
teF0rk0HPV/cyn9Z5GNvHnsWm9xOP2GijiCjNmxCPS7GZ4B1cIMlYaQ+cxp1VNmfyHnurLX86Yj7
UxE2CzTu73QtSTMFwYIURqN12YUzbG4QpnTm1M5Qc3uwap2d10+XrPbrYl2pMDJs6vc8WG90kSMW
qsO+xLVUUUUSuFEjDCXMkDKZU9SnLxYUgBk9VQjW8sE/09YIhDTPdjZGE7FfEGPca2uIoFu2HRxJ
dL+3PZTzl78h20dOLY0VSQL2HX/tUhz50WQzlTuru8Dtkx24TmOflqpgbJmqc0mTcQFSEDfiiTap
1XxgVYg4yz9VEXo7Gb7zTyX17FHRKaDo9Dj8qPK0i8q/tIT/FGYZ0WFOs6HOcqtLy2m9V9Ygu9ux
upDh+1cSZGVa/RncFKCcpfMG8HfFGxOp1oQmYtVwO7r6GrN0ew6oS2QQqhTSdMuCqUYPDE9sI7ci
nrKz+C4IRWDAmSRIX9rK9QdfXQkzJUfYYkc3W+/beh/qwugDkkDbw7x7qEfnHlmiGB/256jaAZMV
bM+pcbhSFhSEsvnbo7bb4CmdTdhL1oX3l1H265fcW0kOS9xPV4MZ+KivP1TatPJvN2noqrr+XEhY
BF8TiDrZ3vSSQHtqROYf3XludYHZSC/9pxcdXQ5hzbSu1UtZyC1Bz66nmXxDz4TREhU+KXxSwVoj
ScflO+2gADWPLSAlTbokRO2NEeIP2qOSJjs2QDIiXEEJZLulvVDqLmnEYrHcj7AUwCwuIN/+Mctt
xayDspf6bEVGm3+gu9Cwbc7kn7wz7rLxOy/UM505J5B8hbApC8ILu7kejYdA1FmEFvzWIlyvJaY7
+CpBwntd34PzMldmZy6ks3zFSoHIAtx9b98qZTuNrXc0rmeitP1WVAWy4um0aZwnAaQcfB/5q5rb
bt36xjzA73As4QCEKs+dZ3sZBYiiJ8Lq+EsldpW4b/xjf7ZtIqev9Efkdyb8QnQrkY2LvFGh3GYh
NAWBvzVq7HFwuD2b7fSAggOOu+HSb4D3g2yZGfBp2LMAJsNzOa3OrU2CSDSiBvwnTSV1uNomiPAg
9SHrCvCUZ+ASArLU6EXzHtOTlQawthDnZ3VS8U4tCRgCoyZjLeAIkp5Yud4ou6Jq0FkDMCqk9RbZ
up4CFb/cXnK8BH5TK5MWEeyQar8FbNbdQ+92HCNn9Bmbn5weJmmfQ+vS9Hbgw97HL5i4JOQky8Fq
8FDwQtA2RIAQfCiMYRTEq0OOfzhykA49vi64MOacKVuJ7hSc2+eqgAxeN4oYzU3DB4NVD8c24Mvx
0+0yIBL+E906h3SvBjqZ6vBxyyRtlXKJiEksR7+0oO/F0O9DnO0f7kCUYPr+lH1PjJ1U8N9h8ocC
oZOqB2k3oHqXNwKuD90vFiW+f51A1z/O2Wqa0uivW2h5BS+46NKd45CPtzKTJE3tqABaO5IusjLc
0fME41GMGcAZH8/cs2czkusUttCj4E7URH4ydRDk1K85fmDvXqX7xPHMd0JDm2B0A39zWHIRFg5E
+4jegpgtjvsNTwBj+gJbh+YlYZUaboXBiX8640uTuHsJ86Nb722ct95cos8XgtAIsCu2wahcBvf/
x0DpF8tCWZn0IMpmeU6cd2VjXm0fjYDQVzl6Q42Rs6thWKJ0SJagy05l5dRDnFRI50/X/PVb+nqV
ZOHBThLpdHl7FntQokEKX18wammXhGzzoqXSYI33BWOLo8NmoMU6TdMyz4V+Jf/Dfnb9W108sAhS
cePIiXcdn+iYURvT+KrcnT352QKYsQ/P1moR2j94aVQ7lNQdhCGx+uusQLmtMAIqdDimeXGL7mAh
cYDebt39pP0SnhdbEpfMEefc8uTSXA7QCVU0z6lzu2Ac02UhBW3htHKhk5Url9UPKshxIEaSVYJN
8dV5UpfrAJ+uC599CTgnXoif38OQO8uERMpty4HNg5nutEaz102boCGJ5djZ/x4wziLoH6Zbx0xZ
/j32YxSPP4OE4RD0v2r1nc13tI8pk/7V3gk4bKTMo+RYzeLsywjOpKBUZKc/jwpsslbAqkDVibB6
5r+VQBlLx86NaabNqnWo4LZXnPQReWDHbgLt0ITpEM2a6BSDUj9kVJ45hnx1i/oyX5+kNL9XuxbF
hTN+jtGUXx3Hvo9npbYXRq95UuxIO+rfqFPsFiqp7A5gyaQmOTsIZkkt6m8aW1AtkWdLBJWP0ruv
VuDCyYcqE+0XIgnucnJBvhqjehQTnKoSLRnXfiyOn9M1UJRQDelz/f3xUwA7og0bTCHRc7vwzM3h
zF+mxhmlQ7UiqQGcG+F3o2f0SKtvUcdLhPkasacKUTBE9WkpEVRanl7iVdKW8CsCkXzagumUp+d1
RPIDL3joxpbjHzkIJZfDgtkqQKVzmaCb6KUfQsddQMXV1Hn3rQS5hcskoIl9IDFIDz+ybaFXhwOG
9kFRC5nP/HxiQZmXkBKZPXiPOIjcrJ4FnQfq7LyWJ8pF+JlVqBSx/iul0nY4LoOX6HMuxE599MIv
s5CxcdZ7hq8XqiSp5bqwiq126NIUd3r8VwKfO5UqlC7ivrBGGEMVlDyCVJtW6syLZ1vkh9l6U+KQ
3plnC16+yAtCzHaJ1K00SWC/0IKm6tSAo80yaoqqe5QkmZc83lofe7eFflwaOv96QAURRQX55vEg
KHWtyv513awAvoYK4dA5x0Ic1ZXV7RxcO6i0kiamlEFOwpNpFGx9rHoPy4ADr0K0UPcF5FHjNM8k
PCdYDZmFSt8wjTMUOdy6OspqotvqRHLPwVY4TCISgPrHGr51SZoLiwuDypVmvWF+a9BJ91TZe2XH
JCmusBP5tkgpUKOjHVKq2RuD4ojkBZIuZpxB6imbBh8ufivJauibuhMNPLej6BhYMX8YCU0DyVKo
0Bk11o5/HgH+NmnItwGEl3vegL/Xv3bDd5Z8uWoqlst1jP4jkZIbp9eCY3Uo40D/JtYXKB5J5YpN
GGSioMW4dWLSJ2trSdyKXXhNwz4CWs7K//9+/Te8+Vim34Dq/a07Qy+UlkLcxrOKGyYuuvyLLu/8
0eMO/J63mYyHVf6bmnmN/ZapKZS8heZAZVFdCFf45EwS13GNvNOD3MtK/9AHhCvDN66NUAajUgM9
BRVyArJAcIAKz+vkIR0bqb7ypTPIdmMmJErg5qJsc/Ib25aMXPtXuvPVIgh81T9jBurKtgJeekBO
I9uZPpniqmSh4g0nISzAYEuIL6y51DjFAQ7+zVRGTByLZ02nm6F1mLb4dcg3ms67uBXiGeF1uCzR
8TaMp40RcChhwTQrXWP2JjVKMoMvN7IYG0efja+Gh2JAHAJ/xayrDAKbNgcXe+WSrcSJTi9PGEQ5
BgfPpdclD83UKkOOlu086vyGAkOstMj973b5zq14nR3tx3ChNYyk9fN45dRSvjQrn3num0J8J2Jw
dxdJqxcyiPeGdRlvD/vFIUVlVSCWQbDAQSUEqJtXgwW7S57B8V1PYJByWJ6l45ss765TnsXRjxkF
3MixSvuX/yx4J9gyrSsrxAXnYvMTdDTj1Yz4nmudXCS+1lBlmOdF8fOpMPq2lbysnOFaCNxva/kp
77DB5BIFuecWylqg41fIngvGEGcH/SfuSCPIzImv96jz1P/lpBiEJzHU1FvISANfgMEEigKa1pvW
x8Hx6awkgJxxyuNan6k/lhEfQk5bGokMHcRZKvs1apK4wPuZhoKh9DkDAD2dUA2joW40IHBHcGr8
pb7c9kG6IAIP1S+1GMcit1UvPOxjK+D/TvuaVlWGe7+nBpxgi/wKqeKtbsw6fsKaHPMi36rxkpKt
+9Y6QlcQImnJBtYDL9iCzBy7IRF512MMOUkLmnEegs701tTNTjO2F8YOlToz3lbSEoezfvJ9rkgl
yGklv3UVUp3kg5Tt2rEWLdSSK8hper4AdNNCFWsp1m0pVj1hUjG4hrbqTPY9167SGriD7A9Cla13
keQCYIjW85T+5F9EbVf38FqD+0eOzSTbTTG7hG9p16kMSXFeQRzSO/Z5+PWXmX/tYC+AWSzB6PwK
DAw07NNfGbLpiTEedJ5ppftuZ2eFW64Q+qmq3n4cNNOcKRVyyhRhur9klmZXlCol5NPPi6qceul+
TTJT/4XhKMPRdryxsREBNrR79fxQLSE9jaWXUr7HjDo8bj7967yHLwxAGHqAUjLCJsXRfKlWKFwd
AVNjgR1inbyA78NXVouIYfvXczwVBAIrrSfEEhoOIRpaLOmxGtKrpx0sPgsXjrbhD8N1liq9v6BI
747TrV1WdpXQMawXlcycgDqm+rNn7J17t8FalPBvuqbAgwEToXebxHrUM5dnX2r+Fmyp+paYGqaP
Akwmc8sMq8S6sfFLhI7rDlMr6yPyOZjO3o/J3cu89FGMdL1wsZxYRc8w1ZbjK3G1affiM75lXuYE
G4+hGMNnuE6hY16MJZGYUnygx3Neh5igrGuYqxgHZ1SVCywbX3boa/jm98P/aV3xfMMT7H/17dTX
DLT6sMIuVFigdVE75y3myNXPAk2vPO6PfgN8hBJjOnubyoQYY5sds9pMRYLgrfEIKzC5+oEEujo1
nbzCb6BwGBFCRwv+rj+rou3wJnR75CaW/9CCVOwiOghf+UIjiMwaMhPVAsIzTgu7vHdIkdDCMz8F
s7sjzdBR7P8MyNA7y6J/osmNRAwZSsyyR874Ke4zagEwR+edtxrZR3hvLsgjDt1o9DBkSzRCNTMD
UfC3ReHB3qiivLlck/6GHFdqj9rH4JK8EqvVj/aVdRjvF0LgejQStQPrjX4e0CRLc+SU4TAB+Kv5
HVQGomgWUGQyeoh4uJgYxwQpMsUjPrg9z4UYda6qAR6gFOY0AUO1lb/fK5SrPGbJcTXMkP5L1+js
y2rsggVQkqlo6VZkiuSoXQgtlg1sjAfcvuhBvs6/iiHDo9EFhI2OeXse6dZ0hN6x87HHQMsXPclG
Y/1CVS2U0Za04M8RMvMAWk5c6HyRLJ/eBTb1d0SedTBsAoZFHNtE7Ehz1V7P7m4IwtpOfFNAVQ16
BEZdP7I6RHlFyHZ9DeAPmP/K1jWn/oDSQrdNcZwN7pUa4vaMkveE5/AV7fa1SM1sy7iQH+vOHXiS
2twVQvJSxXXZ4pyDMiC3Xpwb5bEGB1ZKSeNsh5Ld6Y+fsW5Z38JsJQwlTLx15o87SvIM0MWFChV/
6zuoVJjpEg6YyBDKANlB+TXsMiTQkXu2t89DnMrhdMdcTohCT9WmsZzIvNhAWnN085so5L5bLZv+
FNX6Unx+R3ZhJH9eYC2UBELSoQkudTccN8m50oK6Mf1NvUZ7F3JtjaU0w8JjPO834IouPZW3uE+m
sHHJVcImrj1nhMvYRaDnNcG2Gcb/J8+soBI8ONLHMFEp9+Zj+geXr1QbAhsYjxLoFEmmx0wFDB0r
cGVjabn99hrLljCliucpGWHNE90/obmKXpTbBjZtbxYwdYVxO0n0j3j5EtL7XNUG/VzQM2yfP5TI
qP4fBngdCtuZksy51/UBaXKf2hSR2Dht5lnFiWsPtzhPopQ5XgQN+oWYPMR758cCrCwDGguneH4W
JtCAXsR1bLKqPNbnwSTOTpq1x0bqPw6InQ47ZS1smk+3f3GD75IFmxZ6JzTwDciME3s5IDOVW0TZ
Eju9ftggNc/AEZ+v3u4pTL3Ezq1ylhhoQg50/NQb+rUbfejTSj/dPB31DrMspMkueZbusFJ4q9eI
IUhodHWHUtSjc2l7NNm5K0c09dKSbNUDY9Y08QjHjTslzVGHZaVKx2V6zlCyM8gNGkfe/Bn8K7Ru
9myl7TJ4Gom2EVNwQQdJvVFRup/0MDt1fgv//8k3RTVaihe6Xd7INSg45xfGDilLupNNUUbowvJY
80TIwZQb+mG6VVvCmky6fTXxQZKm5wihUWXcdJvZgRx+aDQiP8+YrXKQ3Ntz+myG1Gaz1s5soFba
OlzjqAPN6bVghXaEGb765/dwu2r7uvrn74knJnH/Xmesfg22SX+y+Spuk42S3x8GBSJQOjadg/dT
ObD1Ud7MAXTiZ0VtDLPSCN/d+/sZby1j6cEwYyN11YcwE2Ac2mP9zMsyTrvJz9LrNLgiNbPcH2dc
Mh2atxrzK/v/oNWx1rzWNlu4Owqq1d1WEJ6ucrrzPnx7obIi87xwq5DYSrJalhtMq8VREvqYz6Ej
RDy+g/1Gx3IkrhIt+jYX+6m5iCB2zDMyz5G8B0+xs3LmwTJWyPW4J+46qjx3NJuFD1ej0DsfyjLM
3aUmrG1ffbzXxf/mV72yAEuWOz4dA4LSxQvpqw8qyms21uQYkScFgtbaK0szEGDF/yJURgDVQ4W7
gZ35z4JtJDcZRVcHvN4709LQ10ec/lX+7eZj27OXgmXj+Rr3/llI8JmWAjlHCKvl/RQRJ3mUQ/dy
K9dKmrAWnDuhETd2/Aw6ICo420ux3CTzfQFcmBQ0PmPQApi5lc8jD+bq4u6KW0oLhlpOCWtbjlqV
NXVqxGACCmJ9+mWGB4wzVgwD76XyyYMAwrmVrVClzrpnOLvvywbw/rboJVmsZLXHPV8h4OPmM3bZ
iRN6rj+S6UHJF8BSMNN4XVljSK5cvFig+y2ueKrURkNiNJeUu6T0vi+wRtgc7PdI7AJgNlopp246
r4tXO3Os/0kiF7qhRBIZn47ZL/OepQTkaGggFhrMcdjdDMHwHIS59EPbQHlayy7HJWz46nX6n1Cy
1N05sdmfMAXTvnImfORyzPo1wG7NxdOQQBLkdooKBqsKhQquinzkPoScBaMEUx4zKLjrKZvl1o6n
0TfHjsAexQGk2KgqNLgEATaU/fBAHSzNBa9owk73y/OyYM8xL3Pa1cYNcAjo3jZm38K2f5pH4Cu2
70kFmTWTl2aIWgjyRC7ZOSx0eho9PeHSlcgyFnB5ohGjz1l2aOXAfUgqsaAqXemDTBj0nXeDE3J3
YSJA314xg2EeH3fXbhM05LyjUDZKU6+nDIQHuYuYNyDEreHKfnZ3m0nABIzbOLjhhfr0EqNb2pJQ
tHF8aqLHFjc13i7Crp7f5jrJB9Rvwpm/OgeNRyJ28InsAX8u5ZAWcH+MscwOGRbtKV8PcfwqGSPW
rbEoGp4DvwMdDSE9uKGM6/frrGnxN2Da1s59T1dlV4yJG5/lBbhCXQ+3BFvLt6lQd/6FAvJ1hmm4
9r6KPpDeNPDtDDZo51nKNdzmI3SZIqVfVMofybkBga3faRf18H9bShHdMiaSJxhyNQxEmvmbHFzJ
R9vjr7NKTLXySlc3M4YPTEE2n5dZkIOQ0t7GFrH+cu/rR9MqtOAdbDKinfMvd6PDf/dG/wH5YADb
kNBQMBT9DnH/vfDDPRaYBS9Zihpk2djiBhEEFxucb4d7zh37HhG8Yrb2Yxk9UleuzHKa4G6VLITX
rCdnK9mKydM70CPqsOB5HblaNS7IATp4mhdHottIiwshHpcFscRBwtYEpUHdk2yqiion3eOtBCoF
Lk1estHIQjOEGc2GE5PuRQr5jaqL7pWBm+zeiv0dkpLT67RXA9i9kccDuSp/AxTheS1PyyJy4Uoq
k3zT8DlZokFxii49+xMOTxUQfaIISOZMezE/5ugx2aVKxndm/PSSc/LRbxpLu1SOi2H/LU72dO7w
G1HQGfaEHPoUv/PEHm7xBXbjLU7jq+n3ResB04PrixmF9gXHk7EQB7rnI0goiVCvYrlYUpdBcWKR
APL+rI/zLxyYuxFfnNIZGd3s2gjq7v9FZvhcs0Rb/ilWvIuAuPMv6iYkwJdmDy8X8hZAD5YzQBng
sZ+4YzPRDHX6fK5wdB5EN6xcy1LTjdyer2/OTpeA5Nz8zN+BKZnbS9vYiwlO10EzOlwdaWJMzbkF
7PCwPC4zDKIHsyrr8BUJySuqIvxQU+zS6zA2eInlLt8A4eionxydtNzyJoiDU0ayFMr/6IYC4n4v
jrmnYpOnHp6ao8tgluHTpviZeNgEWD7+LF3fYG1sjgrnFc3mQwDBMyXLTWbQ6i8tJHLN9rEv17fl
Xf+b3qZnAEKdt0W+6y+GPkglJiSP3x6tXf5jjcpbAiAUHrWAF8r2jyw0EK0rOnixP+qx32sNRpc0
85m4zh8PbVuYvk4ZZiP71ZbTvEG6Id9/Z6K2cokfsxmR9wLPeKvCQmQQTEtF3ZBfLep5eKafBwVp
o+qCegFZND43l8b8L+QpW+yVWSRou+G18IEJLGmodsRNFEjeARYyEorUj7dmYCBgZC96rg4j8q24
Ppzs7x/9BIzcdCBNRZkW90qfnQxqb5HEq7PLK6rRFndlLdyWNKqLyccMNUDRUmSlJNoX2mYRJaEU
OztH9YVXrsJKOWLU4/V2FHJWlWQfO4ubp6I9CfrvBOIAf7uZJ8o41mOvLMfIsyfhJDkDfjGnAFhH
HB/p150WnCGfm/QKQfIMt4j60FR4I4nSe/66CE6v+ObAK7B/cARKP2GsJv9hjVdkwF81dpkGPotE
ns+JmB5NnrOPxLkskhJxbqVy+xCxrp/4gd59oihi0/iqBnWAqQBh97w6rQbGdvGpAv1GEVdeNKT3
IqpkgB9mBOkRZ9p/ujMnjcnA9iCjbPQyv2H6hlIRqz6XEs8Mkp9kgEGZsuF+TdR0BKUTgS1p9tji
TEQ7pPhWxhnzlRKVXKykgLRmfPMMT2zCxWrVUINZbC80a9Sm2zw0HBS4OBcutisFVLBGMVn97+Q6
7Fzto0uvbVcbktmBx8MOQ2mxJ1K49waPRDBqmzfGcJ+MSrDETww3i934qVaU9m7wx6wcxmEbEE0C
MT5YN1Ojk9uAL2pWfXgZk11fX0K+hxtP5oZnuoAlOH+x0up40FPu11yS7u0+e3SY3RSu9O+LgT/o
1M870DdRB+KN81R27unoSd3uvzVC40hw8N5cOObz8TvP1WSuf/CbWwuq+sChe5jIppSG1mq9IuYB
1OhIvL2CqeKNjQ/L8e1RwcjohYshcDjrcqUs8o5X0PD177xcXn/67OkuRZQPhaDoKUBQERzHpEyT
oeImKhAI6uZav7dDC/SqFPNIdS8I0YZcv1QSaJo80jF2jv5ZDerNiPrL1T0VEd2aNT2hyDXwXeJQ
5SwgtWjKmpUrZ27/e/rCS8IlRbxXOEA7g3U/29vSawLSJ+laIGh9lOQRsVWMsWm9E35Jph/j7Rrt
jJ+B+VHGQWJ0lEuOzQ6TT/iPg0NGv7ct8euUB2hrNZTyLDVzwZdHYbommkTlp1FqaN5Hlhaf5rt6
ngW56qEfnGGTQmo3wHgJeLS/whnoH1m8WcJtgzRyMOpqY31GeS2UQGJmug4LaksBZ+nKQNNRMAPG
fo8R5iOWzoe65s3GbHn3Q0IqdcYANyoGm4ClwpOk92Uh0vSTe2xyCyChOyfTZ4+HibHl6gs6v61P
+HpgRHOhgUEIqdrzxZA03yfKoJcV3oHzLNUUcgkEG9CMcp5XU8JuZHx3vrRzvNHyoZrZPdDXYtPR
Rv0P5XW4+06u6C4UBPtGVPWMs3R/7Tiv+IWJ+gpFMP8xwcXPb10crFG4MGpr2bU25viDha97Bcgg
b8M3Kml6cyAqSKwVWrP5QcDPqtOEqTKcrLpDzdpeb0bjhYLi+EVAMVNjGoDj0Uwow0kV4z8YoZLc
3fCZdBH8SWBen9JyEfMnfszbEwzn9B/UsraG6Sd461wAV2qHE9MWCfg896aLMMDVc2sd/seCj6Ne
NjyHOzFhPs6tUd5ebtGhAbC5Cj70Hg9M2tjxTQcwpeSnEjbIOVhVzOy4Qqt3sxBW7BOX9wwGVOoz
wkiXBKy6AjBHSrdt/FxbcutvP47ZGF7fDfxF+5rTFXKlXsEOC4O1W7ecKDEUvl1kSWBwuBfrimmv
mr30bDhtPUY0hKyqgyx32aPKt/ystwFYDUy7AclEKNzf3Lq5vWrZBBd7qfHuB2uF4pzKSmTPo1Nb
HguYCjfftbt8Zl8k3n2b2E/laF4yoTN74kV57H1pUCY8P30pLy5ifaZqDGvT+1SmQQwu9dSvIuQA
8HTmRdsS/haPD4AAaI2aMbqlCWDVgSEV3Eja+akN/OHnTltpi7DqTUBtCYHci4x/BFg4K2F+GDfM
TRjlN4d6o2UDsJUa3PodDGFX1LtWbrzH1XXAf7novmkHX0oLDSLgONzGqlOwZztb7iklYjte4b9l
7h+Lp4fdd3I7dyx4uhXj+tnnWA3ixchath0eNc1nh7JXK54y/JFDOS3BE4uWxQA4BvVlYjpw/vX/
HhWA9OQZC/drdHFdD9f+ZOta9P4JcqMXLXCogJdfQAGOn9iBkChGDw+dK9pj9WEyZ4TsaRhrYslJ
m4w1MHSPgCp1z/pk3/WIHem21aqDos6Hni/7Uj/uhcLYi8HhYyUsotmH3k/ls0RLA/pqBg796IlD
qWlI8kAXvkUnl71NODhaZ21YrFdsRBlm++/dg8/KASYdR1KL+YKlW1a60gT1B+btF4oAaKe6WRS7
fdoPCJ0VOhAFayIfetsYK07TENbkF+Z1H5JyVv1B7WHkqnfYyrgc+n7uAYaJ9B5O6TA5h0uJZnBu
HKjeWe8nfP5Vl4ve2anx9oWI9ubPVMBnnHs7vnfQWbHexxZa+5pJ1EJOPbz98zaHzHHu8qJKu+jX
sjQffEoYsmae53Y9A6W9eAnA19l/0G9hLS8mi4n+Ye7MJEZs7mSPwQxU5XOe3Ib5sxUJB3iYE4nm
3nAisPEJMmViSbjoIioEBNHXitefgaamN5qS50WE57gtSVwliyOuIEy1j15YLBfuXQ4hWfMfSQVF
0UmqWXFQXoKxQUSlGSi4/x+YTtdxl0ELPJwDRJ4TQMGhNmc+2UvcO5gx6V7d+jBkaO8jBsHOjNTw
QgZpss/m1A5KvU8BSA5ydWi0Wsb1DYZop2fZxtej2R4ZzDum8w1DgqhVbHg0aZh9aDwRstKDukIZ
10DX9Q9sENMnxTqApvS2LIpM6ZMl3f31RESHQbnZ6nVrSA+PdVJrD6HWjYy3NN0NwYr68tyEx8pt
o/xuhPhqIFFkAwA4zIflWdsOxl9DcCl+gtCnjnV0HTV0XNvf+Ky5MNhF9GAFIAkab4oASjC2hk5F
9otEcAppmtFY3YYeQuN5L7MVi2Wo2T1hhwykQJxV+kfojy3r9c/CabwKklQOZL3DkBz7HpYqWZKO
NGmXC57oqXMjUo6yKZlbA6AaC0fqwbEZNeTJXpvoIAUUwatASHKTAq/htg+pbWI3xdvZ3AsKueZy
xPaz1ReTyCGuHk6ZffdFRxDdrdvF6Vq0UEBJ8xvLJ8j8vUumTLaKGw6xqIG8JNA07XmiVP5pAP5U
bR+vCv4wWhTy4XjlmciFFkRPZXuSniwoVMWmZnsBHH96HpMgrEN0Onx/Q9D4Swm0VmAhfK5QbGD5
YmKltSwXqxi5i87ZbPXr9fLGs9388N0Mx1JwIkeHMcSUsFPa730yJekRzB8dOiRvMSE1ANOKaEuD
sWk9um6Yg2QynQHSpkutS21fsXXyWs4ytxmk2VpqXPpYY/P1MJwJuFCc8ydyYJ0Ac/XDcSGgueh4
D0mBNFBihOJkvBc+Ik2hVaXqZ+AXnCqb9NMV0p+ODzuylzKSn+1vo2w1G7bvhg8ChZHsyBq0K7fy
HTwAVHz42vLljcyEfjHS8sYpXEH9L4sXgNDNM1hrGPafzPMm8yzpv/WaLm6Q0wepAmzBSAWP0+nb
VaiH2LKdc1Bi2QTszsh5dFRo5xkFsYG0MgT3lccK7+ugzSXy7dUuduwf6F5BQYTuNg725vSbhJdA
A4aQn7GuKBly2OYRS5NsHKJVs1jcn5IPWDFO1+341zUGPBa8vxnz+gzBbjT96pnUIdjUxwCSIyDS
2DnYE3udNnaqv4TamhCu2j1fHlN6hua72PR0cE4gWN+LaSaBwXyr6jfYh0XX/AH62/ECwF7vYhOS
P6qg7/4gJqS6e02JQODWhS+GiRUzRoxAwRLhV6OhKeAm1+iRnOTZ7YIn8j4BiWCf5bxjh+OnHcst
5zERiCOFk0aWm5rop6P3BZzHvbiV8Gqiu1iArVjAq3nd9Mu0z2iTZD2ju9poyvX7JUPDk/VI7VIP
q9kVoOqBlL0hXZrLBTPSMq/5wScdXds0lrJnH7TdRHwLPsqqrKq7EFjymuRvMjX3zbglVZ09+8y1
sJ1DkjDLQMilGomBS2EKNK3F2A7a1F2jg/bjn+MdIvGS5K9akPnJhmfDB47qdMjiS1lzvgYxDnNR
KDdTyi9FKT9DK2WiBbR0HtgQ59uGMv1I2g34ntQetHTKlTktO8asz9B8Itbv6M4uE63V5lbsg0kT
c9riSsXqw2cj+Bb5os83vRVhhjLb+chikXcl779xpfrfBq1/ahu5a6oxd4m2nBSsutOMe5AUr1zc
dEIcpgRE7TO1Nochn0VWp8UIVvhV0iBmFY04npyCKkKJEDrMA3UJocyyR5UymUfBWQtWcYUV+7k2
OSd3VbdVuSDUh3yqofm/WU7N6d6RuzL213bKu8KgVlrpFX4NLQot66/VkNvuvo08k0lCLeIG1OHR
b8O5rhuBZHuvJEkICYqL8dXO6WGu/sH4rh92OY0pYuJaPzCQKGEsmfTet7p7N0C72QJ0GrU6R7WZ
TNslfwJTV1lMbniZZi9icy/108JEArhKchpNsku6GFopIDsDRRNNWIy5gw6h4c3feFTdFwP6FYlc
kV4+OyP4hCB4w//JfQv9pNnlIuWkHk9My68uJ//aA9fv/9FGhLRPRZv/HCTzO6e+n/9Kl/0XRzES
9De9+eTJEglWlxKTaXZb9jsDTu5sBsEKTgXQCp9Dg/FWSq1dzWAsDA6D4fkNmRqaeNraPQFitZdv
PxJXWh8cnIlO2lxA3c8pmn8r0tT1VsyqPGQHMHT+rHsIr+lCjm+yXmKi1wzEewRxuH6HSyFQHsi7
P0Z5Bd4KwPuxlIZc2pxKIeWxur+SOoxDZ0sVYLFbRF6A2OI0inEtzanNJFNG+qzeOHCniH6Hp4TH
ynkJApIu3T/RG2ugaGB+dbpnnHW4JmecAvnrGp0RU72g16KYgh0VlWLCW3QyYRJcGt5rlT5jb836
A4KhwL0wS99rQZiTvNB+sJ+syY0z/iCopBnR0fJW1w4vFVtYv9WfRUqgPMVteJzcJWhvPnbh6Fw6
iSgcCUp1rllWM9EPEbfUsuNYtInHeRMq9rEul2gFt1e/1aAO1TAxEA/uWCvwegf+U1Gg6iDqRe8x
C9wG8Bgi6orUzHL2TXYDrEh7hkciY72j4i2uevAPmODXYcbbB8gD80Jip182S9sgjO3oU07Zyl3i
tdh/0AjalRHRke2fvW3MsmK4MdSOlOoPbILp4XZ1jlES9bWHinzKbpZX8puO0GPtAftvTWyLWTdl
mobefJRbdwbQljm5vM1YoU0ImnVuxWVtyFKXwTK3AplJRhyrFlMhDTc9Tqkw/tvQYCkHb0FDMm/7
SwGXNv6XuQAe0qJrXex0hph/GthoAzphzNVDJsmgEwLrUSf7z9QsJYM4tluaK55rgheuvn06PA1U
mH1S8eRqNEyD7DZGR5+HctcW/9fu0fp0tAQZ1yPvQ69ztmzX3fnJHEOuM7avuV75sLQZuWfZ4Gxl
fKdRwPLAzxnAtqciybWAqujrfv/48PQEhLVCRnPAQpZXuNq8BrPmI5hM40kzmNQ++Mv+n+kZSyNm
bG4AT7NRNqQ3n2z9Rvinh7ykUxupi/iAS6QAG2lVORWeZoFzxT7STESl6yxjP+PRxMgQWMM7Wv1K
FyN3zFi7rkLzyUoKYQsyLiamg5u58d/aFPpXRbor5x5wN6Ty4V3ZZkiTy1JjsfA2hRCPmLWggjxQ
qf0HZFD4Cw9vQD4CB2/dDqJhOJs6bUs5sopGcZ3G4/qWf42jZ7bptSkQlXb7BZwWnZr4S0y84IvK
Y6XDag7oGrCvsUzqJ77Jt69se6/F8xlrUyWR9JT/HHuyztrRkrtbzowrahRKoOukDTTYuhZkWff3
LtI5JhiW8GSPXpASV7Y0P9j7/d4voK9hkDoJz3O7aaPUIMm7WVt8ZOxrv3nGSPBfwCeU2y1RNh0O
7qtu7kTzRH9UKf0aQ0hgVDGEaD89g3JQLx8ypsnWq8tiEemuvKBbiz7JO4A6vudjlywfTAQQCjH/
Hb/SZgm5XQwyltLimqlpVaB93Po4yaruJUqG8tKnhHR180m/dD5r/RidP2M95tGZn0//Ne+PGUM4
D799FwwYhrWH3YzHbq2BY8TVKuJzurhrbG68FKH7YuOLmhq42/MrMMBb/sMMgRFLcX5vx49qIH9B
R6IQwu1wXMcAzEC6OwOyog1iSuKwpTfvKAlBw0ENEnKdlSiGYu/lgIRgSvmUtYQe4+jxGsWjp9sC
FQrp47+CBCcA8sLmoLex3LGpEEc5shHeqwVNFb0incq7tMUFhIkysKbHUKfNrogTEkSRrFC1WA9g
lBt8C92HRbNODa7rGS+ufgNT4rAxzyBtIwpCHeoDRgGdvMpAbWioIpwRSTASFGVzMbRy5an+njWq
q9xIcfHq9beCfche0ZfeEMu3cqMWeeMdVDWsfdVGlO6rJnjpQ3Dq4Stt6wcY1qI5WbhvSiSIHvuW
Q2KA6/E6JPTy1Jl6KF/NHzu8H4u07PHJjdzILEcavruXgNuJqhC8Sx36e6GQzojB2Np6WKjCmAXl
07wnDpfSrUqSAkFQOtu1gz+msvXRa4CPhPhNdYeYxt1VKw4SGrgYVEuYEHylgomOWXCr2c+rUnvV
iMrdHZqsmhgrasO3yCcsLMsfdO+c7lDYJG66c8Ve4OvY+cLSDtfHn4LT4QYHlZdCJ7IzsMS3F5Ts
0hgO7g+aL9IMExXwAvnKIzZvmA5IPAkf65KWvN9FISjaiz8mc2V4frvtlcZKtSCOibOQ79/ADXcm
g7MaT8CCLbrIwdhbseIlZBEu7b6xcorlw3/r2uSPzHsB3Oay6fKr/K7mnYO4AcqhsNusC5o4TfU6
/mXKqZmPQRg2mv9A6fcc/bYWnodiFVWAmHIn94PpPmtGgCXj2ribuU/8LBpxL3Us8akA76XHyN7t
/+BErdA/8uKE5S1aIgK0lQCRlstAwHmTZLDUZ363OrpLE9dvl9rvuND5jd+gTzZCpkp/l3sVd5xp
C0uFv9R++zr4mwtELFeZGUgwSGb62biLWNgSZYZI89wyPkzT+KB1w2PgAr3ouWUj2B/0I4Wx3uGY
6DYsMdNpGWAKflv8GixeWgj3IlbNquRZDaWZxquz6Djag1cD6CnpugcwZj1PPxv/MNXaEkfWrs2n
XzBYuQIK84fU+Ohbq2QyA0RfQVjP6wFG+NTOHgL19JKMb7pjjLeoGsVeHJf+Lnb/l4H1j1SK20LR
qCf88AGVHJFfCgpP8TCBXr4miry64TMFi7qMdwJJLMLAcB7Wc4QZMCImSscxnVpoeO13Og8jPsY7
W8a7nQHujwqm7TMJwAzLWfpVeAv0tx0GE+70ihVJWC8U6XxUrDvU5tQu/cHpPnzd0rwR8Qs9Lc0n
5pfYCc9VgWdCZQXfiK/wDSgtIjzULWhbYrTtKKaA2r2uYPF4rFI9XzKiF10IW+7Wsu+UcVPByV0a
kKcqCoLmzWr+WYluzu0QCe3ZcQ+Gj7khQnCWvuD7FhWzXjSepvCQZprdtCuGvj+we5JX6i6IhBUw
DuQqdsO8/FhI1jrRLMbhGFoOzpPOfC1/606PPKzxEYX9bP3d/9lYrWinFcMYebUMa5TlczpY9hSy
eR0Twzkh3wAcKmvSdvJOiBKJvL+xnjy2HAz55YyvNl2yiMDWwEnt8s4crP4Tm1A94rCsaCQ04NYA
2YhiBNe6CquGWyA2AQkidh928DEvDjeybLOBkBs3M39c6hF3756p3Yl0qOCd4P2LAUHwCc1M27VU
DhG7U72AAxA0FS6ioR1Ud4MTQAr2BDn7dt2oLQjzPpzQEuU2z4Ko6WY+N26mVSBazlgTWzzTJje0
f+rMkdpSsO0+JMUvpVwM79vrBa4pFRP3k19vfBV+Y/TZKfQzxK+cCFMTncdQvLEwIE5M+iv2Q1be
sffrXbTgdwqlFL8vRlqpSoFrR8sDbbNicMyia3UGtTywJ1UIeoBn6wQC0eDevAijAo6baoBmL5U6
N9Hoa+GVfp+f1tAcNtpSokidgPIjfhb7nTkfUoVsU5hy5tWEf151diJVE89lxu/iJpV+mW/E+PQ9
f3zjQaAqtfRn0h2CZH4OcJZFXTrUVXZT8VXMCSfqMuVYi0gVEZ0glKas9gvDr03xD9akF6RuLeUH
mE/+vWs20eP9kC+Acgr0q4v7e90Y8gkpzR7FS1ZHa14BUzrB01CghSFEoNFLC9577vBDQJEddGqq
GGaxIvrfPrcDx69MhunluAfnntfSwLKwnCC/Yo74bPoWTWciMnO05ZBvW1oHY7NRDQtW2nb2L8NM
r4xqObNEPf+yZ8EuikK46Nd/A0G2QfHXDYLvD9p6WWvhTZ/ByXfXx7SSPUaJLLmem4ZrEYhqet6j
54I13uDSRImfUsgI9in42Fh7dj2AtpGfCRp6jwj1f0NAtweMRr9pRuHhrfvpa+YddpUCisthtNth
a/KVQEv+eXJczDH5iFUNHf5Eex5lOnAT/swcq7XBaQ7GgbCdHdcUY3ypLmvmXs4aR5+Qwf6yLnRD
DUtv0l/G6Tr34Q9QRPGxKFwEECzEw17xdzK/sn7QHuBqoGaEcv1/Ro3y1Ub65sTqTSC/8ZoqOuqW
5LGXDPWWLgArBDiKHtf9FkZoHJz7EZt7uEB55C01/DP44CWYaTRLeT1PBgx5Jx9cxIUYwQ3qQBMx
0hhjfBOxvWR7DqrSeGwljWoG9fN0VhoOcOqEvXWBwdqhe8/HH4r9nM6w1vCuxtuiM37JOuUyWGD/
VwhrpFBwcYMb3Jcxj7Po7At1x/gxnBYeiY3+2AypKIkwHNVeaoGOwPqCrXcfnCvFsH1NDrjubsg4
I2buFnzE3JOFNwYvxLCKIOS3XvQLqucapKsgaIBXRAm6nQBFkeIIknS/VPs5KK0wWtSffK0YbDof
Iy27umIjZO7+s4YdLLnOL4cWirdTVCGfBV010PGcJfD5swLMZeVedXKJ2Njlue93qwWntWpvRTFN
IOAtl8wR3WAMLGBqzHqmx7jKJ0/XzPv1czyH0AT0tBfxnKJn8SeyVhIAcAtjotP5AG3oL4vKxzQ4
Hsz3ns7VVe1mUWHLGMb3NINT0a0ERzkv4CL1aRGc5A0nXQ/pr63oGDyOeJpcsLaDQXxbjwaawaUQ
Vo9+McYORYzbisxk96Su7LUB2M8JkK8DN9j489CnnW70M5Q8IlVUiV+F/yMKdFOq3WaPuKu4ma3o
JVRyqonz3ES2Sj5u86Lk2yjF7dfj3hJh8CCs93tUnBvo7/YbHfp8p14r6OR2CKt9m0WP/eYHSD0j
0z5PrHJsQgElLM4S6yZk1RhEwWbTGy0DTmnm15owJpGOYcLV62qJVnblEamI1RiXwZ/8sWcE2z44
zrEKhLr3tsjjlhx7Ep4/geuhVEWEiOG1zEeW2qf6S3XEcVhjn9/+Z5HNjcI9SSt8abgYNs8/ACXF
H4F0GQU4zrMKEt1rWNqA4C2bjISUI+lqsJl0pKPMlpCvenO+/axR+26TVkxDAd3WKe3Efsbi7e9E
gaNyLhS5Trq7TWBknODQkZbH6G16tC9fa3q3TwdG8LWykCUbK99F3LRRdF+N8spANnhHgaW8/Feh
KkJ9z2DdQIX1xLPU9AVRHlVlSVp5ZVvwyJL++pX2rUYUs8i9wOoOCyVDnkxS4k1Ht1QyyqETXSZe
u20CCLMzG5mdTu9Im1B93fo5SqP1AVfgk0bGCGzxP6ZMqx8hPhoXvitWkkHaW7xQQe8PFcYnP2uz
26+x/e6hd8Q1pNMNwNhPkRN3IvnR9SIyTZoqHszy6Uedos1jssxAfkzsOXGWVXg38N68jtfBW0W+
vC40qBI+dFY2qGXZF9yXko39azvnXTRZVCTKn8nzCm/lZzobEXMsLYDwnFEkMyTwB3FZH6p/WtFa
sKwQ1VJaXR/+0+7JxFvzCAT//Cgxk05yxcPTHUiaBiBNzIK8jsW0i4assRqCxlGDhWG7cJC+lyQ4
MXbMGcUjYXFNPp8ozIJ2+zEwoxVrDCw4NDtJIKPYI6bAcOGJ+Vt26Had9aTMy6uhXHmxrq0qtPbP
8z/Kl1PCrSae3F/52sxHOzf7P3Tigu6fyVrgWjpqOqFlhCKMwnUYcHSM6Rgmal+PODusYHJ/Qf16
Zp+zEgI7kDGH6WVzIOMR3XS+yPQnwABb0vSV3Bb/CvM73ZhUBMUixjKZAeK8KM9IzThM1F+IvWIe
xrZZ7fcI+oSN3w7PoTUMfwMfjRBT2G/MZiQGNKkCgeF6f23vog4dCMvYOm7l0lwpYSVI3Dv4S5ay
ievEy6qmjKp84GlVFOhI+zhzdPRpGwzgYFFmLM8jnJg+GBt9jUcLhDtIkmQbtiQGwtgj3oL7lfVe
lfb4ztW70xHllzZXk3Rj8/kv1O4ryk+YP0wP9eRGa1T8ce42SFsLMp971ZPnucveav7BvEJV9BsL
LV8+3/oI80dBcUd4/MWvxExB28BmKPpbxIoJV/tNcbVOO/wa/Xk2rGuDng1E18Pr5W9qcNJVu2SY
C2ibfYSMcGe7Ve0KXp7P8iPJ9bKtlUOOJ3ytobQgCfU7c+AfqmC1+RjK2SwEBOl/faBBIvDSwCji
95ee4MyexUqdMog544gFPWuAOCIzdXg8n19QjTm4+m+2KPXW9dIT8FYeNWSEXPbIfWQeHK9TtWp1
kOVDYe2vabHzh2WtNfJo2XKOKwOSdd9vIAHF5WNv2gt6lwpVX/+JcJWzvkTyDn59DU03GLeTFXAX
KalQAsz8fyCFj5wYwMR6a0T13ggQVlc2YkIuPMzIUu2liDo6eiHVv5hyYxZmpvDEl/qlEV6FuTY9
/+qu+4eJkxKp8Ydu8V++NRh+IkeqXIIpVHSOk8fWK/EwkRQd0M2PX3TDY9iEPU1+o7/BTHWWbbti
oAgOI59ZVZfk6Q69G06fUpm9L0p5puts1IvCSeu/Dv2WAAos68wtg6Ie1kHf3j9o9d5n02EUGJf7
xI7XUJWimC5vwdS602/nxMo0kWM5dVzRfBRb9mO6PWChxAxRu6eXxzsIDVBdUyZ8Qo9l2O/9ueId
K+SaspJEbCf02z9jkH/5b0FvZl7hx0ke59BGA5Zyb2Vdv7KdmRWaTmiJjqg4pi80djgrkfJ9INGS
EshhstOUruNIr53Lxu0zoMVlfZPczYO730yNKNYAaynI/UTFxr7GX3c96U7ViZJ6XNh6zY76cjor
y+jstfhv79eUHHjyHSRpoj/b6QuQEa5HjoHL8XpZFtkPkp2ZJ6Wa3hbaRBcHwx6peuen9otYMxhd
MLY/KrdIHKXpBov+3VWy64kp27hE8emkfNleLQUEEU7dMLoFsE6g+2lP5/2e8gDQf11wnrt4ZYff
+kXbMyHT2mF8vkCl2htDG1ZHaQjzpmNjtFm9G/Ufsy9xBK/UZSkBRGfsId7hScplZQerjp3MLvWb
qRRIXoZNTptJYTNW5OOGdMSfeVXY0zuRWa3G4fQDhgZLM/4G8eF0WiJ8Ar8ojCXroVwkkHg40C3f
ttI+DhpSMoUwgTDyHBi4nXsaiUwQtNuYOps8/IJpqcbLa6PJllbuo0KX8CSKzB+CiSV1Wqu6U+R9
wSjkdN/OpuroO23x5Kfc8O/0NbYwv6ODzrxzuK1M5Kv0R1Pfd1m5FjffpsENMeSI1qXKrg1umJPD
wuQoisHQ4Iq/UF0NFNNirKXH0k1XZlPVpplPkL2AiknauyG07uqHgE7it9GnYiGMi9Ti/UcBDEMR
xafyDojq9jK0jdqL2e8zD6CijJ0aqH1n/kohi4/ZwatwCfR2Vup8dogcZeXpfZu2/kLZ0uo33f/8
7yIxCj/guZkCVq/em0ZxrudnBb8qf8yR7DGNMITnGoaL7W15xrMzLzEYFIEIrJf+GjxgHiQtjbQ4
6HBWjVKFmjt0R0CAn3RDuuUdYTBO2r7K5KWKFunzyWYxY/Gql5JTL/9K5nPNMdMb3C+gtgp82741
4E0N1QbKKRg1ppDSqNIuNYHvJcDspEytypPUnHb7vFELWaxuF4+fAMg+2BlzhyFwsW76eVDcVUC4
cq0LjeNsaFEE2kJ3/7QVFNC9gvC3LAC7tX7WYjQJvdWecPPk80DgpzS2mKFiXaLl8ZF7akHQ/7Kj
Z6srnfDlejMGlv8FXcxuJ/GmVePGKbeuudOfx5BPOH6J8LLdNNwwDGBzatnR9jnI41a/slnCn3PI
ElLk9n15NtX1M2aDr4nvzrTwRRKkGpDB6Gx9Mc4UK7jhE0arjY0JGL4qJr5ZXyuk9P29EgpplH30
FYUT0BAUfxP9z7kLYH8tIA+2K+2KfI8XvUbiv6ioPw8e597zc0aTmbUIBGJhLv0nrJx07tURhH/m
4wM2elfwbT07Itum5cC3TonvlbrpkPjfT4BriWL1wHWVGIx9toCnlQ4WQ+m0Xj2E/KW8urqtCIFe
kljwt76ilOANyVwCse2TyHXMEX1p7YTHXyyYL1YCMBs97RDLwXeptbaAeDebOFlrxcDLxlFGeYdc
mH1OjU9gUsbz5Gi09p1Td17GrKbpF0upFiuSNJ3nKXdPFvrsBlpNmWBklhXxZVLWo8ob8MHmXGGU
mw547oIF/uTIPJH7DkX74PsDTj4nEgxdBXJH1deFONCdMu34RNxH291wOzjLOtT7WEIvf7DboOJ9
7IjIM71vOJEPAq6BuE1F2OEz/D7k2ucBHC7F31aiKFW+fDfAeFMPLX8XlFO+1LBhupNaUGKyOzQo
X6qpF15LJfQXV2TvCuQWGcOd6TLMIswtSVoRB4yqD+Zx5PeFISLzTY5XGiUV+7kpCmGv5I6dS99T
rLO1WjnMHAZkcMKAXUdSfAdpAAeEA65VAw+i+h3QLglwn86EYBc6Usqb4BigPPr4OG03Bzd+2y0k
ziyxAmhW+0KItbt2PwJ74V474ZlGOej+psC3c/fFewSDTNnOJeExmGEOvJk2P50bMug1Kgx4Upd6
B8VFWBeP/vkFJOgz1GUdZYJkGmBCs+G2CAPn6JGveadGUUKZPc3Kw/Z1B/pOoP23mDDMBmTj4t3C
b65yob9GNWrw3VXdpZbgKiz63xPJ93NNMHVI5V19auybuaNjJ3IcsWbNVkiKT6CBA9P4UAXPCpwa
/6R7xtKBIn94upRtHol3CTdG0igoyYp04IAUW9FJ8gX8R3gtvEU1udNlz5d4DixBEFvnaY91ItRy
gMGn0zrDtGPTVzCgxYpQ1e1eTAhcgUHnsvdIljel4Ooxh4J145EQHLRUkRvIp/kLoXwLtbMiyzSO
sc0kxDcUtqkuNFogT6UEwPbwFgXBYuemLxxvhiCt2Q5hpb9ghITlgDkTKaYU+XtLDUG9WGlTfKiJ
cvyEzo4gIlIvuwYZ6fjnpFLgCLC5qZlf2dbGWmoxX8pmjGkYNsQuweIj+bNtChzyVWHTu2NSzwRl
L6b5N+9j53HbVuicH0faFQZVvCTgxpZmpdg1+QxXGGEUT44w0WRmoXBrMaNQwVXAM3YtA6w1W/JD
IGblbTblRNV4vl3fes/b50e6Zp5La+63FRj+jDG69MbNv6aAldqSVdUCjvZEBs8vKZOnq0g8rtWs
sCBNWzeddF3LcwE6jn5Ecq76gu3ymR/LKXQzIzq46nPwkZ//9iAc/CvyroPwoS0+qQV+AmoVagCl
hTKObsDCwFQCXDaTVtp1FPm0m1YXDGAVJiEmT+7IFgPmXBlgf79RacVTT/wNJA2xouhYN7qhAS5X
kiK7RsARPVT2P3Od6iCjkf2Zpy3gCleF8tnueiD46fq8lZVyGmSMEI1TuCtW3ZzcYmZ09YROouGA
n5WDBF2P6AmLcz/YChDLJOF9qJz+XJ3v0U+xTtnPPgoTd0vHXuC7RMrUd+Y0yqV6wpXWX/gYmHeA
3mQtS5hbpnDLvfKJOHiDS9sSJDa616ITe4OcWHt3CAAKT2L4VAXYzDG0ew0JrOcaHzrL1iNz91hA
FGaZYo42v+N8OcDRdW0MOHp7p/fP7JLb2TVX51Br3tOGD538n6nZK9PQvxAkTtMyvVgUNcEJT4lT
rFoZwecWqErZ8T2dATIZ+Y4DY5gUq77gt6aZBh3/jU+Qv94svWLPxKpBy4Ksd44blYJYgi7L9VYE
IwDaiB8p0W0X6X5PyJkG79une6O7BMqPQaUIR8NWmW5nv4arv/f9OgMq4IyY3KHZKu3irU1lWMHj
pGJKTXEoeUp9YCtVZHBh5qxOqOIbBRALpLnsRls93YxS2eyhE9BeqnFvbxfAlliZozWTdYgV5xZO
bWKenSbmXWkkF0HdspHpD68d4lxsAAc6Bu2bxp3xQbvZ+hID9ke7zSxximCS7u53FBMg0RaZXNXu
+6ZeIkiY0XUFN4v369OgxWdABmU7KxcRNz06Ekj0SsJXSfvGRMbxDRoMzbvzRdFtB0zhlr++CjLK
rPulIMuycqcM0z15agTXo3tlnhhA9FU3ADDUUc085+g9kZNBENgvEegq+1v6Bx3maXZ2bggtxtcn
Y3Fvq0vQoZzHU3HHiF79osW0A7YokMBhn6cC83/UP9got/DDrfPknA8HRaUEekPxG4xdIGDsR/sf
hWAiW9kFxKjgfmeM95APfXUxIZ/T42VXzzQaMlm9sxpgDPt7hNCQ43x2oQFA7v2vdWJltIZ4lc26
X5Dxp8XkN5EYsmeukjGQ2V3r6yEuKU/FdxgPRTQ3MIZqsUiEaA53O2+MIVarfk+Yw6VZER69rBO2
upCXagEwtuOpMKSwJsi5pEgef9n+wyPi4a48vy5nupaROOTxUoHRVVR8zADpwjorx8iAZq1SDEOo
kMD3jpykLP5oBNWk98W1N2RWH/6PtorHnEOZMI9wwyZeJHW3jdvfm07mmJMgwa+enAnO9524GKVh
AQ4NsiE/9kgPsJY8FO9pse6uvMuGEkFzV03F0fQFOvgTd2bqXUnjMWjt/KrNaSKqba8yfM9l7wdX
nOsuovSR2Q6fjBGaUcg19tsfYrFyYDIwni+qS6kCNcDLY/zQNFCqbXXawgb5gZTVZRWA4CNjIs+q
WegopCh+Goc2yji087spbaaLT844XEAiQBaxEPvBHyuIoSQkB9So9nvNo4nq0Djt349Bi3u1GOb1
of0Z40GKvx9eFeQ6qwodjlw6Cbrw4GwfnL8hsucTVXmR3B6OLm45Oi/tDjItAvMBo8xbc19t2Cnh
oIC27Dcay0AuUjOSjyFJdQppILBh+pnp9JvXJ/PxNu4AHtTJYMV0NlGyEaG9LGk3lJ/fRY4y8AVr
9MEODGw13CrOH36r+BR6cCoNdyPwmX/nosMzvSE4TtFaLiY46YhxNhCH+gVZmK9Fnf6jTJu/p0xQ
M4niGx4WxD0TUPT5E2VJJFj6mEFeFLxnxOvxbwg7HGM+gTpE89UqXJgBPQKvLevsCV2fcsNnf+m8
Vk+uyzrEJR0FD+fBx5/oy4kM/MlfG5TQM6Bt2Jf47PfDgnKe5CnZBTWV+R3BpQEgHSH1mTbSY6Vz
WiTtY2KszruMdNZu+ucsnawdUNw5YRIrma8dKxRzAoLzopvPtpRqT9RYqmCxSwobrvftrxQTXwH2
Otw93YAG6KzOHhFa7pHQb4945HK3YREVpj1559UhodSLH8mWi2N4hx3IwYhdSz+8IqR8WA6ljJc6
qS51Qf1fNydO6/gID6fVTA24pPq/5VrHGhvJInnthMwPWMgnNOX6nk1nvln5kgCjtox530F9JqcU
gh2QC0w3BgQRTBD/FE5GbVmywAs0dLsG2tCF2KPdTq0OvF+qsQDwWM0ubAQr5+cUqgTXQvwKx5ny
suXX3s3/cU1qdAtqqRRKJ4ZNcLxOpZ+tFc9cGwIbsDCUcMxMvC7a+dv9bFNlvrg+Jcu5k9l0SG44
NrH4f0PrGyzZz8p1ziXhpkky3Q2EMCVq/LfjQUO86n7XS97cB2AR/vGvL7ANXH0kVPsXRg+TZ5Jy
ceqsyMUn4KXk3nCyjE88K/OHl3+URcPoLhA9DgpQZwInnsCL6z6wtXzS3KQIJynLyRAh9OeTlA+x
Vt0yZu7VKzTzt9z64j5CeSO4d2u6kWrqZr0FAubOEp/Kc6ucVH2VD4Cw2E2xSZTLhXjqczCKR3ym
oN9S5NNR1O4+t8LTuGR4MbWy03DcBMcHvVBRfkFqf/XUvVOVmI34dw6TbGejYDY2lqYPOb33xyey
MuSq21sy2KaHEKt33yDSZr1w0KuhCAst6O7tDFNdrmnKy7fcPJ7taOIeO5EEkQMA3/CKLyRBJI5y
48Fw7pfmjl8eiNLCv0UFsMcougDW9do0xMIu/1A58ypJO2BIwgH6/qFlgXSvbkplt61JQPOCKLMG
qiV9PKA7WVdwvl1nkadl2wfrDQUugmO3WrG/tZJ/6o+gO8pTxTQy+3oxMLP39t8WpGTjV/UWjPKj
hCzb+q7yIhIecQIah+SMCn7li65EuxI1kuC9Et2x+/VLKnVANtkNCoZSMQjP2TagDVzVeJ5PIqUb
GbfG+9DxiDY6tf4x2H4/t1917cX/6t/u1Dp5BSpJbMOU7iCcIC+wgkpqjGDLZo9OpBHWBwtffOge
ZeyDD0Q+lOgVfNPDvqa1vOJM1XEVT6v9vapSaLAkgHPv1mDy7A/bCacY7WUBaOtU5cYrzrd075EB
KpM2aC3dia0EI+Vv86oP53de7kKpKsRgPzN7GBALjxsWWGPL68MLSYmQm+EVOQR3zgyBG04qdLYZ
nCcwiSFtW+v6CN9UJHBcwarkEIruiwmegbMK5sit3WbCk91fM7K97fEntfqd+xajmuIJJ9KbrSUJ
BuDJUaIMiSPRlRyASBeiDMMJOE5zmGRsVTp9Kj7+vQMoPiD4Yu99Zfy7i/V+xvRJrIqPKnKktHLC
oJp4ffAn1zGhsrr54/2R2irZ4xpb5kIiS/PHpCl+iDNr/LrwDBf8+sbhZDeH7D0SPbMcFR9F4OVx
mHxfRjLtAtLfGT/KoHdCoq/B87adKstcBLPMFRK4uqFYs1ZHdlcLPhu76/UOxocr44RPGh5BmPMH
MGE20ChSJiZLwNUWchYxEw6NdrZN9ATS6t/G7yiEzKh6wOzwY+zftt3c/91PmcGu5DS5CiGpIO6+
ny7vOX+943xSUuT1E0sODGpvrQOK4z91UrsBSx1leBuir/Ry0BcQwcs/FgpVA4nxQuRJDtpw68co
+lfg7OWlfP8gJUeovTH5OMFTednkBxNFKtSMKhgmoScLHrjeGJrYtnOQ/hHZjG4EP/jJfGkWgu8w
/ugId5GspQldzhiUW/3X9rJ1vQ3AgzpDdqHvzwZMYjft7v2a/eidDYDMwVnP18daCVfmkxeGHSvz
TmIRPKm6l9eI8FUQ0Ow5ooXDUV3Pra6YbqfrarRRfxgWAzgUVANsfNWo/Vx6LSb1NfzEIE8eOA4t
Mli45/V7HWorGZViFxkSrOzNa07nnt0wFXEl18wwFAc/fZnl+zFBA4Zy72ggJrozuWOz0DALehtG
luiFwQhbweYiYDWeBtNGW5ogtCGF21BUyXNgZgaBEwERVvvkQ3S2PRthOL128TpdakVse/i1TY2/
0IU5H0S5VpcBd5rWFy3p9NYv4i6boUBwbQ9tKkqzOASONy2jPsGX+g9kNlmzb6357MZwWSOIWSqE
a2ZhGFBzNK9UEAyKQL1i6zpVCJlwtsrh83W/iy2NieUvX8QymuILrXli+71pg7wxy3y0devrr5fR
2vapQuWKdDmJk+Ryon3M8d+ItjotszugjKjZbWVGnZDP+T15/hUiJ1MzQLg1YYHRcETcvNElMz5r
iHgkq29r/VxwwEsyOKKhNwu/Qr1um/eyWDn7t/sQcjSc2GYyAB934hg5eKaYTN9AWE7f3bGWB8J5
6G4X7MqjxjlfJ8Gn8na7a9t3ND80t51GhkWzeTnuZ3mZlrQBRg7hWj0BLA7xGgmDVaINxwvP9c0s
GpR3QO/ot1L5WI+fMWUeMUiPcAHrbiiKX/GvR4Hjfa9dGc94jqUEkwJr9y6YuSGeku2d4qSBYq1s
lWdBVMPZbaM1s5hNnyFfDv9UQZKJD1WmhagpFeWSimzx+awHQVz5/07dWYgiTyL+rFHjjHrjeFbN
s+JlKzTVIcY90nzps+DLr2njRcLQmgOy7lRAWRXRRQiFzPNVpX6gr3KyxbqkZEhYbUUopuSlBVaS
k/FLpf/0bhQOv9LjhgwM4JMWxFG8D1/Z0LbWmmhIbNAqs1plb+C/YXxLc0KvMkGo9V64EDiMrLYc
Nu8enCXQF/Paf2c3ZYSLrJKBcW+3OGXzy9h0JedBW3ma4lppah0b/CkmgQEKkyF/FKQFUu6bc+X4
ufjCJUrBKhNizdnnG8fo7tKjK3jtgTUHdL8uve4OePXgWlEzsiMYx2eZ2ge+uDhC5upCeGFNYmOn
fasQoRhlDBlE3kemTfFmlAbqbok7qhg61FjdBobSaJu6mkB/RXxDjGYetkqJVRWeEJ/KvX+uhiNT
eiFr1kFwXZMS+e0rg9inaSEcNPuGKbEw49kEcp9WCgDOQ9A+37HSS+/xmNlSfSkbbmUs1NRwbk0v
mHYy/gcuQEZZ980qPhG1VPE+Ig/DQFKdCJd0UwPatPdJNADFaqYJ0Sj2VbIf8c2aIdSbosclqlpA
lIBExnEMk7CScJIXgUu17f9fY4F9czJ7Y//tDyz8gesWJSjFY9Qhfi16NpUD4o8e/HIUvPrOzsLW
ZdjI2foAUf36eGWtAabzEWSvvSFG0wPAgJX0kRvr2U238otvkZ+Rpfvkbb0oJcwiZVPbgnRXFVuF
EajHXf6dRuMfvPj8OtAtjt/j8PUhzJhAqvI/1lBThbktcElUtr+SHmWP8jNXkXKzd4Cvsn+UIRBq
dRjh2sSnyiz9v/uQs3WOtedhySKYi7vmpUShUHsAryPSaS5HFusfeI991Nug3vNYkJj0GninaRnI
DXkCq480Ju3YfJP6Uxai9yCUKjN0X26GzJzHMNYQHYpSaQ9a26O6wbo7QbwFmn6eNKUiYXy5CPDw
Q4OWzmD5k1zlsYRBWxu7+g6csHw09cw65902Ofno8PHrviI+HBcFnFCApaZx2OmXCzzzUW0JfMv5
lI1lKt9uXfJL57eOlzcZsmJ1UoJOIxB5qJRQ+6zomlcPV6r+21ujHcUcwhfzQbN8/Bxr8N1o5mte
PImGyvSKOs6AsrJX6fwfYITnM914kFa3tDyJ0TKWVa8aGlddeifAlDUmPqTsJMpxJUlj/v2pBAAP
mPxdAd1LW3CiEUBEG0CFPA2ZqgWoU+7sqIIQ6/zLrtPsYT7jVvIYdUIFs8HCILYpzkIKvqXlQ2F1
J+P2DU+DCAOQPZI8kggNqSS4a84bksjtwc6Ef7rk/LlNU9gFa/ZB80u6mQQyoiy9ixBIxKlnPji8
fHplKdDihLQ/mHanT51UiIVMOH8iWPoyrX4wX1E9R9v2V5BT+GLykNgp54L7CpQnlPFaPKIiEU0r
5XMVg8s3PuDiLJzQSNWZj0EpDzk/iIgIdunrQOCEXhQlKwGiG863YPUPa/PtHN1fSfnBUxuVi5gj
woLTaP55VYHQR0B8KOy3TWrxyGBDxG/NVUpCI+jaixcqT/YbgrP5Wz6mOkk8Sd2OPl4IQ2scTu6e
8ymZuxNDSvHHN4uM9mwL8oREe3CpgFddqNqXUS/ibH7nPAJPqKI4cYjphv/QDQsH7spXXhN+g3QN
bjbxnr0KS6lCsxtyJwaLDcEycBDcTXQIGI0eEucfXtnyYm+o3z8IxVqRAf8UrBxq6kTYyqPIg12q
eCWusYSStroUtaPhUaG1CX4KLKO/3s06W2zXBJqH3FdNhQWwGYd4+i/s5UE7Jwmj+sri+zjSD0fT
kz78A0n6/Rm1/7w6pZVnutPJ5XQJ3Eoicn1IBd7bNbFw+rNygxK7hoEHjXUB5wwO2C5+It9AY6HP
CEW4AIe5MFeC1hHNsxmxmdr+3VjLVp0zIja0B96fNDYgsMKcBHn8jfoWKk6A4KVpGVD+uJj//3xo
1cv55kldLYpuHbOTn3YHLvh3uutZsQV28wdpMaMgXW/dFLDBYx5/WPpQYcc0+j7KA1b+hGH34vLf
tJzVBkAceVJCR2/9a+MsZ+o/5Ow7Hi24MjQeihO3NpBgJGFkGlq2VULHnevYZtyR7gnNPQ7PB+AC
we7jV5V11/qqQN5a1fa6bpWdMTsj8K2YXRhbuP7J7aR6P5j2FgekUR6MnG1jqg2D/toXYHp4KRWC
hp5+0mw7y2SJF2TMe6U4P8sCmyYOHiiCz05zqy7mllugkRlRGXNMjsKkgCwOQGdqSTbC4s7dq//g
TEtJJ78RQ2VzM3ZrxNVdNdrAnD94Sh50q5RgSSKzuH9Zaw8YYp6tf7mdvPtToIjmW5Lx9dOc4MYO
c9RWGA5ARV3Dpc+5O/vMC8ZFI5Ftxqqo/zuzEDJjMt8XLq6dir4MQIiwGwKXoA6HZK0RVrJqFuXZ
Q3henBT3XBJOFAUlaLRrXAOghZ1V1EabLSFJPyBRITguhdDfF2G24UgWxCCvAxAIFnMuIZCJeuff
IxiuNX3FUv15xPwyuXCt0gyr40cIgtX52J9yTjH+kucUoRf4+O+Zt7zUjTmngY7UU99VHO5Iza7k
T9NsHI73I50TVxu/RvSOFUVBy7KWRkDoFlkY37jZf8sekNNVjWDr+9h+rioIhWDaQtL49XGkPQDN
TlqyunBGXYigLhq0P+yzhxzBv0b4FVLirMT17U6+dxH3OQx+szNZFR77cxvN7USznJLT7tdv3bDF
PsfZuepXx+vIxuJ56GQtNcTWleBcbkRd66nbQOfxgSpwRCPkiuBaHj+nxmNtrDvi+0GRor57SY0U
xA08XkO2PaoiLrPyn93vWvP16loI9qDui0iYrri1kOHJ2zU3NYlqtnKmNyH9JEeRmrRJ2lOOLP+B
ydbpncAwnOTanR8QhQZL3A1rPR/iPLNf4ru1FnZLAHWTATw8qjp/5FZ3iCdX/ERcoe3BdxJ269kg
Sea0PAbfkw/oICXoB+Pc/DDrvSsKYkqFqWR1WI/JoDbxmruHAlIb7jUCAMF5G22Hr3N1v2xDu2kw
OPvFXm/VeZbs8vpwBOHfOQ6nqC70KNajUMVTebMoTI56NHeTEsxFFwGgzGK4YliTSiyGC/DGyVxq
h/zRCJXJq9XWinCwAjae+aySLmublrxqIaHibvqc9h5L41PXxzgXqgUxU8g8G2ZGmkcO1ZgVXdcb
rws3FCIbj72zLvaB3eVqK8ZqighPiOndmKgHVUY8+bwKOJfE5yfFMhuoIeAxcINK14Nk9LwXwQtX
DTeTuKtxwX5yhA2FtGJDGm0jU4AmS7MuZIDtV7IOJcvjShl5mKpy0s8pxUSQpwsw8L3CL/rrrcy2
sJmpf2qZe2o1xKlzky5d8CaXEoSpjxQ0a+25YKCrSuKknBVp880vnt6qC4zItnJBbCrc1xBruSVE
rZOa8bHmc4/EC31Vhk/uIyquo5+dIfKAek3AEpp2K9yAbjE4dlUsFHcdzTV/woeQLerp6v/RCDML
JZXvdZoIgTdjKdo2vXaZgTpDpazLouIAdT2F8EWxRcg0VR3FlCHnflstpmR48M0pA4oU/3CjD673
IjLDCGdBlTO12Uq4aOvqinysv7DAcxLkw5nx1ECCSU/XaCWpzoZLa5f2s8X+jELpRSkWUvNhjcZm
NkpWFTuC+EeoJz7EaMi+04R0Py4WUfgViywAQ24c6mIZhi09Yrpw52NWi43QPugwkh9L078jqDIP
cc16RVS4tOV9I2I0KXp2dnS2WgBIYXpDoRVuxnGU+1QB+4JJnWf2OXbdzFGUgdS/6db4cGNwABnt
eCSS8rWE4kPatld4ethSHMzLaP7xW9EJaOTrcSJZE6cFdlfPhbDYOLyy8p45sfq3kpfOBgDYnKCw
2AvrwRTiP6PYzT/9RbAhMhoi7FemxcMefoYFaY+9XFmkLnYToMbdE8yczMamAABfQ2SEahhHBTlM
z7WaKiC4TB0QTdMWSk1s6spIlBhmzpkRtx3U3N4XFVYCel39aLF/1VamtaC7syhAhbebKtG1NDHW
xBqZGxAkXmYC3pS6OFO1YORQvEM2kKM4zJrJFUOYLjbbyzNUQ4sho75D9vzaN0F+7W3KjaWEAjU/
nHV5SgIjsreLXR53cyoJTudosV+Zo1h4vsmZkrW92OgIikj5911b1CPkexk/Z1a8yqreIFS3xNPJ
XoOkxBJ2Vp4oM0JkOILZpys1mM8lI1qGGgRX4pBMaJcMWNhHj/su/lF4KxZDotPKFyU3SIIC8pZ9
aoL2ibZ19tKgrJswxV7PFuZm3E19LaQKMjQSi1wGU6H4HSbrUbgAMRLUbD+mQpUOwAA4VkNbnf3c
hCF8c7zxZvKxmmBrZk5ehAjSJ36DsrCTgFkK733tA0e1i9fe8fXFI4jfP69bBnR63OsvhuFEQLup
E5P+9cwSMzgzunMUhw3ot4FxKQLlB1jtpTdSH8bEq0O2SIGn9xrttTpvT0HUj4JTavXnJ66/1Qyu
x5zqEIukmpEACeOeCmGcQk6W2IpuSxwjT4Hy+c8/yugQ7OFbe7Pt4UIzJ5hncOySUwzIgVa/+WkE
2VIRZKKOn3JrCpLKe67ugkO5H6x6MNPNrfbIIla6l1djBaHZN5A/eLgGhyLbSTlj7VgKeaefxLaf
ZLtHIASPLy4MdGojfWw33hJXQX6uLBMGf11f4jm3pfOoc1LA8bbkiASrPelItdrvoRh1alOyOrn6
nFRLyfQyaDznZIVUJw3EY2n10bTSuIrkKCMP7qdWW7HQuvfVtQeuhvY56gmG4svgy4QiIMbQVozH
mcuodGrIiEMqrArnaxZl2ta5OKYyAFxcwzAVJau7OCQwd2iOgYsk/n8XxtxH+PPlRj3ZOpzeclNW
Ed5t7sHcfpmFFdX5OVix00vdjJ/hf5F9KfV9fPCfzJYoWBUak7lInahbOXCl+WeZDL1nGNe9OVHW
T6GpN9GdcvC/oXuNXbtqn9RAqCBRiCg0dH9I0kAKS4FgiJ2enXU4U86AsOJhnhFg0yEFy5iqQkNL
6Ja5K8ks0q84e5cQ0iiN1ZSY3uZh876KJuO190ZWXOf8pKIH+ZCSMwTGJCSTd0TxoSiuDnZHHlWF
zFy98K9eirFpqhsG0NRILfNzu/YSxH1cz06Lb/aVCVeG4ifU9zYY/26DXMyia9bUbUMmtMon7XcI
U2/pmAYT2psK5QFbDKbC/L86J5XShCeqMIYCKXc9bFQezboB+m93ibMg7eDA3EtHU4Tz5HFSj1Pf
swrozpks6+nUBqxp0Q3tr6dAOTKgtPgCxyfD5zkcvPDHh3iMP3loCXkGJbhQyVXLTdr8g5b2LyUl
d5QaJh2B7HT9QRbSD+hSqOfvEklOCEatkUH6OKl6Ydyw0xTuEWxdyW3l+P3K9mvF0X3fIEQ4ZhAZ
Lja3IbtVRny21fHq3KtUGgjtGBIuaoApj6zxR1jeGhyyBo4WxAyBPTSB9g2r4tgsMpJOxLYmoYYL
jnTqBHRpJPeEQCxqPichUe9AoFj8VsRdcvx9DyU4P9PcDwFV4cY9LgmVqAamy0LI17UE2WVcpi5F
MzmrEscVWKwDQa/Z0hNm0a3gI+Gc5kAGBVUt4RUT2Q0JmzmeFN+PHbJIA3RrceAyrCompGYk/3Bw
3Cx1I6rifKbN+cJZD/vZ61g3msdprj59hQGNwUawToge5IpUKvAnkWQ50RoJrkRpptcjMA5GqDcA
dx5riiCLuOlnXVhGjq3LjLZow5Amv3v8mkSp4iSSnz1Q53nYz3Gk5jzes57MmB1vViR0BkELQhFk
YdTfWQxQeSEUGH93en/CLy+DMEBm0nu87dmkPD+EmwE2E/nBUI5nVBEkgWe5m3j+OhUMrjkfWmUr
OTsxnDlV5fl/ALhU823C5XZh8fQMGm3HmlqBzcs9xfwvhvTKYzL7XgQiSpDPpBcRdWtAtGu4gSye
dLRAQTD4Opk4ONX9qfqZdJ2QOYH2v1bN/+b05+7Zp1Sl0qBMPXpyehxLbLl0OIdsi/EMox7+MtWK
Is6gfafeZ5sslKtYze7ktlAiBMHnnc6XJ7iGxD4W2TWDz9VPZ4bCdf4QJCkMzv9oKfw0nHrHKXYw
E+tJc5tHBhPFxqU34v8IJzlQV1XaQz/w7SCnE1utTip1jnNMyAAWJdAEwnM1JSdGkYu5ZdPX3TF/
zYyZEEwH6ZWt/K7gqF3RYPK+bBO/v7Seyen5p1GQc3arwlSOwdtG3tmX3SqmlboSjhplXiUNOrSJ
ddzWf9osLWynWBhWBSYtgs4MkN/zWGIw4EkhfN1Q6FZQ0YhYekRTVw3ZSY1p5KVNg4K7p628zJ3R
v6sXHCI7xREHo29LmTmwndjnm4zSYnlPfBK/uQcgySGh4XGAUVCEH1oCOvmBEY8IWrYoKRaSk6yf
aOPQKT9OLdSqKFU9ByVzEYd46eoDYNJ27Eb7VIFgPCWfzsWXS0QdUDHMaNUiPSkmOXGcz9MbiLDB
OAnFJXPOC+DJFpxjkfadSOg9NRtAhHbb1er1SMfNEXOQKC9UDhfZhlWV+0ePKrDM+Ix96kX0uwXZ
bfltuV/dkOSRh5/ggYDigvVv/8dUDqHBP2E99Ddeq8hmZ/B1yTey1mxE9CWEBbXVe4SIqUQukTrv
gpt2RAGUid1o/rT82NFtyY6nBVnzR6WBXnB6YlC4j3hCcnUDBYiVDXQXtmDMiYyBsqSxlxYF0D5n
qv9CkDOhI1jBvV9pPzPE31aQZmzpV+BoeI1pfJyhI7msch8ktE0QG+xm2cOWRZanHUZNlO+rj1qi
dHBG95EUfD0P6ULNRnyp9K66onzxoVWL9BYXlMS62nmLlzSP1TacByBmhcPEWw7o5OxgG0LhBCXT
pDa1EtIr42m7TFY6/G7CBje3XRNsiZGNNFuq+IrQYL63rZNeQyEwH5bYNgqn8DG2ROMuq8RilfUq
rWXBMJCDnx+unuu8oG6qmEPmd2HYWnUvSxgUIYAY2tw1SmQb/T6bQVuzuddQClHULLJLZYHpfP2I
2QsqoYj2Ae9QZJSD2eclvCcPRoxSlasGAktG6IORMiDG5y8GqexH0RESPd86LjwZXoHbDF8QqRDa
d8ubig6UDaf0azXPq2pIHMxJp0xu9VhI3hzooZhwkF1LjV+1cML1Kikj6B1+wBjB+qNY9CRRgh+Q
xTd0+TiDU3s3qt0mjS8WEfq39jqxieXA/GBI8zYh0yETn3LgnDpGtTfc3uqb69MzycINJ/z7Lg2h
S6OryxD10M9vD0F3q8gkADkg7pk0UAqATbJbG+g6V14Wa44Osa3zKkujHJJQ/S5nN/AqMhsVvC1/
vzM5jM++hyl2/9AFleUD3yBBLBtYpnONMVaH/4Ri7INeYCm1P7NZB/kdWUCgIrMhAn5OC4X1eiF6
3eyjlI5x1+hCqoU8LNxKylYVfHbOzQ4HTWaJzmYoK0kWOffD2Tt4D2aFt40fwlw+dMRTN0goT9Q6
FqUSJfmsAMNR/OArt6y0M7+a8uA4w7tJKEWX8kLFO7crTct3pSqwkPBFRKoM8bnvbMh3cy54Dr1Z
auJpDMOIBsaoQpwHcz5fH2Rl4UxZJK74Ki79sODHScPA2YcaEyXsCBQUvTYXiUKzTyCmiUPS43zv
vFWDo5Igyy1vU8mQVCrrTzMWftIw62O9he6/AFPIcwr8YqBeFr0RIaFRPxugpj/e5h3LOziGG4zf
WG0UWzZklUjZvro2L67uoyAwPJMGikXrBKqixFk+iyXZw6/Kj6PDYmKjtepYL+otPXsHkuIjE2hL
UshuojGioW5Ks3tcnBlJz6hIo8oDXN2RG1s2oGw2N7I3esvp0mF6w8JqfZ0uJn15j0zfn+nfnpU8
i84nhMwRIY+ZCjdrtn9S/ExDx/cXoFm4WB0fZV/Vrmoo6wd83gLEiIWHMGDLDP+hy1GuVDOi/J7P
MZAhQaFCdzmBfC0cMyLt/jx4uoqyM+3/qqX3QIkz4Ii6Ekrg/j4QLhI7kLoh/c8XnjHWrEYDx7r8
7zf5XVn89XjTMs+q0klMmuL2yCz5xyAwyKVzKilrHa/Pfg4l90NY37svao8TnRN3xXZOjRyeDLZH
rZfNcbbV3F489j1QFumkcqR2hkwvFkbK0dUKeGpAgpzq2wpFfGXhlgl1eayskyWURHvfwHo4P/pM
UfmsjTfIFg91+JdU0zWDDKUW4f4Uyp+MDzwj/EFWL4XhjYbQE7qAp+mA1UlQOQ68iwAwYxLakmr6
n7TLL+PIkrv1StlMoYV5Y5i7PYVbi+sSyrDXFIWF/UEVCt9qUBRXj3FTlBuhByqoHndG3BOnyEXM
uKuAJ1SZHGTwagFqikyU+K2iB2aIhEpyJChxLGa5aaQi7X4+5AGSIZDE+PigMxRs8UAEFyFreK1Y
k4B9XnLUm75lxnquw2geyDm1tqLkwwS65UCUjLpOjh3nY1hO13XRhP+GFQITdcAYZz9YtFeE2le/
m141l91AWSVhr6Z/oFX9CgJHVo/JZAYZqf05gWKwjhwdvHXD/bdB8MwR7RU2IVi2zsVog/Pe29Ps
hA7K2qlSH5vT/GWpgS5W8WqlfG6jK8HoQYvbm1+U1Wb6Qf6svHXbNF2l9aO8uGxLIrAB45P/5kdl
tl6EG0d1bhohepaD9xgG6HvezPB2f/QWXCQRfHksV2tIPpU8d3cpZNK9IN/94cIszNhpDZqvtqbV
3UNz+L2clWx7B74qm93PI4ID6iInm+aOyHeGWk4ZK7JMoGGEccMwHsin/3jDMQE5zg7W96ckathx
SuHpWVf860vvzBhZ2k8wYLGd8U0p1E5VcrTfjMh+dwT7BVjmfz0jBb471oi3Gm/M1KYbvvQHAOZ3
pjbDzOWfjQzP7Hq+VkDPeG+gu3ITS6Si+78hb48R2jAWYpC0v4Ediu/GDLDk4HoVnTxivAkcbAxU
Efx3ayB7hw0ELAkHa0vR+UMujKtLeFvK98MXbvbk+NVzzDgke82pHGPxRWdVaHmxhswnR9rAOuuh
/h0/4HbLhgZctonM3cVXgy7A6xIL1cfEOAgkGscLq6KVQcXbrJCpL+YOGbFJsgWhp1J1sG3uhEKu
FnKsyfJgWjzEwA8aCA5Iv96oJQpYaHB88EvtF/XhOv1zy5uD/RweYxpBnZUZyjgCTOVbNggwj8Di
WotKcPc9L6109ZREXQebK+66rZHPQaYUltq7bSUivk0o6CUuWsgVQkovOyTlUD484n4CMlYAXPa7
GZjoW2E+gt7J/MxU2YOWt6Vi5e6O/2HUHmFGRnstjPFAlOHrbdU0FDQzvnttqy4n7hGN4o6Or1KH
/iX1UbyjvrWEeOL3DIEQxV0pE44rNHKt3bPAOvTFHhElFe5oAdFSVNYQdsOSQNZENAL/DGbNfGS/
7suyXDqdlRyFd6YaUN8L74RWk5rU0cNzHM+oS4VScytjZT3RalFsyZ66K/Re0QLIejiTHGS6Gj2b
4qP04DhPgaX7C0uO2o5+gop2BhNl+oiq/8Y6d5VRYrHycady4slNLRgxcE7TQ7FJlIR7DQbK+A08
wNonngAjCgxDw22VZttJYzX2kkkE9LloNDZfyXPxK8QKYHJM0j7o0JKBDHtEltOnP6rlag5QeXyj
CLAFrIBQNqpJzDtwkQVReLA/B4EQGKn1t7xRz+qWS7kcST/nGnlXb0zNis5zEhihwjDwtL0VmVGS
HXVYHEO1ETXaDMNHZvVJluGM2b96/t5lbiJW2a9aJcGQNUFdmtZJ29DuRrXKMgbV9SpNLvOIyZ/6
pxWIYr3SUlLMs64SEZIug0aGaj5hwo0Jq4RedGYOpUI4pBzkHN08jOQ3lmpp2pFFA5kKYmusc3u7
HhKBI/UQVER4imRqI+C6kvQ/BiZHzIEX8mAT+4yqBiVX3cRYoEQKYiuwHawB6XYAsl6Exo6A3iRw
7QHo50fmf+2KYl9rOMn/e+xregt15cMlAUkNdZJ7mVYYWB/kugIPCM8m3RYJW+vVmmPx2QNqNgic
L3BF2vYRlwpOAAa/5Lx09FrTw4q5GIOBGsK1GgAjRa8w12h2MMVH4/X/Av1H4jSE/aVv1BvJ+s3Z
wIlyFYQHuaA4DCbxQtPXT3U5PLn9vq4Aqt8kzdY8/OpZe6DZU0r0mJJYuTCVrZixSo591lXhGETW
8hTu030/wGEU2IDjV+HvjFc+FMweF5UI/CyNn8hVm1YP7E68INsmYzIaDLibEjaDoQ/zhb1bG3B0
4zcq3oHJvqhOYMUtm8MiRcOOILTHnIKTrtjGQ6z5jlok9y1HmKckAHgFLwQNDMh/1HQrshfCsBvh
KN1uPx1wXR7tKIoz3NInMDXWsqWtypAaLIq2UTfzpBotpYYzley5bp1stOFOptbqZrnjSnoUfA7+
8o7w/hqFPxIuBQIjqywI1gWRpP/YXgjz1uBCOxwNA1N47Vw7VQDSO0HjckTOrIW0U10gcmGqSWTl
7YOL8LUDEa1Wc0mPkK1jF5B+CVz7Aiib/3fkKnBpKhYHj17MBegqEzytQVNS9QzmeMR1r6nubMsK
jCTCx7aHy6cAim/1bNFs/nQr1geW8bq9S6lNq3wC5zuz4J6FElH9jgi2/Z9hkNTcdG1X4E4fiTXC
+bEddXWF4x1M2S3qyaN87+VfV4lRnHzfVKB1bKk6TJIcgTliTDmf5+5DKKmCz4Za0NH8mmNi3SQe
oi0ojwlfeC+GtbBpgcyu1B/RhaS8viuRIjtEIfqQa7yV3tl8odz4viMZdsVSLLb/u7IJ57HJivPK
jj7jo4+3Jw+R3g4ANT4flkTlPE9dbybxGeicZgAApEbZTZqA56fBateA7rhvfua4pJ9YeSu/INji
wV5uTWXSGbDkJWeLU56H4vWfd8s/YRvZPlRh9kKaAO8ZHaIERKck3BMvP2WNRr7uwYNloRPPGwiz
pt0C0+33J6rNwPROof2DEhh/OqyYBxerXZmQs83qlOL5DnZmfKp+EqJt4mvJgcl2OCNahLI3r6ad
nfXmR5XKfxwvpRtPKusXS26ZnRRw1l6scotO2ZNoOpcOqpg8UYEweUqrMbqpX9zQj8e9HRoq5NlL
H1g5rqKKO73pJuQ87kYL507dgVVLn8ypfmpBcqcYpD0V8xbFibbnjBG1SZt7Pwhkow5ApVJ5dai2
qM8r8JwqjEzvLflHK7Q61osnV4YIbbFHyUBxQIHNcPpG2Vu8UsbsBT40ZOO8FxuhI3kqxvgWhdXf
tarEOSlmFF9fUb9HdhJEt+UGHU40kDslu+P2m5uFhKUEDoIK+p2rtWgWYnC9q+kZvnCZ64Nr5ECG
6NlaEAu4R8Amdd1p7Id6iHcOMuPsAUuC8PqFb9RixykB825g61nKKmZ6i4NL5Imxg+xeZiShAtbS
TeRcNVTeKYPsXNaUh+rUfXYZlb7MIcmTiGqa4cXOI2WkGjFv6F38TuADe5hv+CAjK8rLH88JcKLd
Vf0AlpU7EOQbdtMQ9Q4fUpXW4OBJz0ATXQUQrZ+QutGWCvrAmHa0ppKMHfGBKxHO13k1HcqGkLt8
t2Ophm0X2XZuSRMY69CqDnRoQ+s+vlzyVU218jtjiVqqxqaFURGTCrRA7YeONLEfXuGnSHtmztHy
wLZ6sfHzPGtuivR5jAZTmEoM2rRneuVzwmN7O6C4vi0QTdcQM1dwBMvefWKCestWSvTxixHQ282u
dTUmU0nOoyavLXJ6gqVC2XOliRVGKlixr674ayZ15fxb4a69mtdwoAHc5Hc2n0LafKlHlGxHDRU6
eq0qPctplymiNf1WnOoiDy9cW8vfUcbZV4iQn0/hD+Rsarz7qmlTRc3XKoZfbAJxgf+S325WPX1R
X6WaagTOuWcxz/XwlhZeFlC3LmYze/dQUMnYTuWzhgjpHMw88kTQUJ+oGQZmNrLT4t8X7nXIj2pl
bx1XGscTeDJ/MovHTFuZKno/zO1+lZWiasedwD1YoP06bdIlQ1lzkm+y5K/CqTHTiIT039WDa8is
nLUV5K+X+DocCe1TBq8VSNgKyfSPaqUthp1ZcpBQDl+sgnZ60IaDlyCYI6zlNeei3LwPIp9nqSn7
cBJmLylJh4dLIp3jLfDvTHvNqXq8ePIyHOnC5Vz4IWb9eu+NexCwe3Wlwl3G1QeiqRC40wyhzpSr
MzFwhztD0T5Ij5aSrg9VKOUIhqti/77KGNr8udnF48VGXrCw8vYZESX4R5axufQVpWRkAlQpPv6t
Vvd22Pqt62EeNor+DNvMhxnTAY9+SWbdf2XfW97fjrcEJnPNhasI1m6Vr1riTRSXZe5F7MIlta+L
FrFIk4xAC5G+Nbdhl12iDBU4UyR50cl8TedAqIIvSBjhuiP1uWN7NhAUSIz2IbTmjy8mYzhfHUro
LaLYwFAHiKDED9dlELn6An6xaU0cSHXBryEW6pijV98uoFyQmIWD8F90/gDr/zQN/Hh9U7Kf57xG
elaPmCFIHeN0+Ub69YvRZIEhJ44TS5PbprbDv1x4crsPvBARXXg6BeK3Hp5Vyfio3hWcfz2jUo5g
Us/rb/jsCsJI1kKUXc7o30gzjkkj41oxQxzZ7UKZaUfkepKdIWmr5WOEz784UpeYh58YEQsoOF/O
9k+9yfyoEXpIeQojCfyjO7Bnc2bcvWj2hPXMMIjD2/fACXazD37Ux8ST2AUaJzT24/i5w/aMpotd
6STxkT1/8prsDyLrcW+GQ9RJT6cr93TD42G9TTEmqRDUexKX/LsEFqllYk5QMIYXIsUbP+D1qv0w
zKIkXttJ4h4hPBscnDH7EIgOCZyOnatodKBH+Cst6JfYm2/oj8gPxRWeC8K00lE7s/PyghXhVhfb
a5Dau4IKp347bF+h60aXHbXQBZIcdmA3Sa3+uW2ODuT+h8upXZPmPs2U2XPHoz5YYQhbljtE2omN
HKsKq9z2suRjVJjs39Q4PKl1CY1w8oJQ1TeAIEMkMoB2VmL7P3QAVWBVIfvI1cdoxEdp0Iou/FvI
obvuHwzTwL0XeetEQlLLMEp2pvJ0v/HAEMsEAVuyoeFWQfjswZXYmlcxHCASLI/Gb1D7RrtmQmYr
Jg0CKf+ax+e5PDwLG3m5H+H6zylKZWzyGoZWgT0VftACgThyKgmYvpGKPW9f6BKtI8qHQaKesZZc
IrqsGpFN1fuTiYdlf0p73SRBQ6EdVGxDkFte4GjMZVif5oiHCcxPP+CLw95pNIGFeRIG9r/54qg+
xxlnYx+YvnmZ0PS97L2uHeQnveWIhfR6XeDjq+HXn5UoqOC8bAyFB42lYFU6Q49qmhAUQTHqq24N
XfRvUltVfr75KAp0jrA7q58L0AE5lj9nKx+9pf+dxjeuXqAgobjvVx6veuzZuz0q2VeZvNfJci35
dCiTC9X0hNwnAhI8gbL+9iSCIibXAkAHM8cLmuSJiZIWndGvdAz98zUYA1wdCfSBCURAzdBCUX6o
MwPzpuzbIIA1TWkHs3A3xTX4RVlg5UJrxNrBVnFoxKiafJPxM0W0khBAk52QcKcQTam4jeOhDhQg
ciViVl/sMOtD2cUqNb7A599DruyeHdfD9jLJUuYa1K5DQ4rIdB/rOoXQis3pS55S+7Zgg+XMstWR
CGpK86Z7EOHH2xUFNT+puKODuvAuVAgVuv8IHjLZoQQKQiV7IS+IDMqnMdosVp/tX5NDZ+IoFk1M
fWwEBv27rjrUBr41wrXO3TenPQ1JllMW9nazBZ5Q5f4aGeuHTI9dSp8tY/OoXT2XKEMXDpPGOk2k
NDb20/lAojFnwdk7JSt6A87TQX97EgFoIAxNvuhuJOj6VoEPb6aFXNU5RQvtQJeIGzp/nPvktGWm
fqBvsGaJzoGmdF0oV6Fow03OKMTztrP2a03JOatm1fdMNdqEo5bL9FAED4X6J2H7FkR+WxUsfSZ/
YUGW64FJ/RC31BhwemzkV9AyQ4AnhezF3cnGynd4Fm9z3vMpUn2wrry+JLbSgX4tAIK9MZPUI3dj
vPyK5WL/Y9iShTkN7Foo8zM4Lbmzn6sp/vcbMzOWncGLOiw8Dve4zm3U8mVKNQG2PGbKxGn04R+S
tPVLZZrdgZCs2kd83MV3j/HUCIiyLvVDo6dTznEYEpUnZxyhotLK6nAEJgbhlgEu6WiUs/OJpI+E
vHeoZM+GMQDy2SkAJe/CmRla83q3nNs6oq9z68LsP66wsFBYfVOEwAgTAggTxK1LHiFndx+TPBOJ
iXngT8DrH73aaoKwNEgQS2twZZdUTUYZTcAsAWTih/Xw+unBF6ACefJu/8UMKVi4rl9/rL8rLORV
bwBnmiBO6SGyoAsxvV6yyjBASvHbm+Zr9otFJconXdG/8ldYGpBM+881ZwbxloMrYW3Xa/rgK9fz
e8Etjy1gFE9LFJ3orspuSmXcwVVAzq88SiPHO64tSpOEEqoGPT1TtpufmTx0Gw4BLYRyWC0z5xky
x7AaFInBtVsUGj/c+z3Ek79BzGSd9m9ue1O95DIz9YLw4gtAyynKxVa+XKHmXaWNUy3NFPui1xw4
rpNOwRoGtKRGyEI8oe498np6rb8gNfJwHaL7nPE3jEYyTudGfBnt+ShNiTuuFDJM7jmB90vQZsGY
fJbeSzdGB5yIUQi7b88aAVgym/QiUcolaoxz2h/sfL0NgfXUSIt4Mepnwsd9l+dOnfupG14tq4qY
OE1Wx0H+RUhe/BespENo+lVN8cZZHExhTEbegAus33Hzup8T6UDlmfNuYESrgC02qFzvWP8wjhyV
j3WPEshUcn9kGosxxdbQn2Ch58Bt07drEFJOAEt+ZIMR0Ab3Tw+552UjdnUVUSgmFpOEBgA6ifzQ
IMAhFt+/8t95Il2q0kIVopKrVCo2IGeBK+NrLKBdm6Jiq3VNGa1aU/YaRVGOCXu7+Rjy0fWePFUN
WLAQHVG4y4nLflBmmy2VKShf+GojPtjKq9vilPhzzsdFNokGXViyn5+t6h6WQTxVghEKkQKAiHWh
Mj/DTegov+t0TZbo2at6L5h2Zx1B9AEhQUygmXrWilnFBbFy6Mb3LCsJc5U9Kl8kiGFEJW3hna3u
ZHuZbfmP1k9XYHN0Oj9+NtHvdwyzxfl0eRfqAh3Vx6Et47zj2gE6m5ghDrYNd9AT893B/W5h2jGO
y+zzTsGDscuLwyEPA92Ydqf2levyuHZlrAy5aHy8QqT2Yg6aVQMZ3Fj0iFBEmcuiTtU3QB/xhkfL
5KUSPWzhc+7JWmfV88TWFYBt/mf1bKJnGifxFQgfzavgikCEKFNLeGgd1cy7C+LZH4pyedK5ZER8
mu6S/r26SERLvZbPJ/MhZXvVzegQFqysHz7Vv9vGy3KajZ1LN1lQx4qhTmVbi8OZiDCu5ZityXtn
7sdLwLhTDP06yciaox+bd9oNncMZ5sokxlcsS7JJT9rdB3qiNxvzt6ECLU2N4O7xYfG0wH1V7DXu
8IJGru/11gC2d/MS3p27OymABLNhwRgXQCou0DoGQRju5uJC//DkucZfF6/MM+SJOq35PS6zwmg5
cFAYz5MeK/9iQS3hSP+qkkrojn8Nvoet/ymITHUlWK+4UxsGeVYAWZgrw1/k2J7Wgkcq9tHFkdDw
IAAErMkYNkB9i5Y4LzYhe0IhM6lpnwdSNJktpkyoPZqg/y1kcpHB/u9kO8EeTRi8hYs84NnuV+UM
V7fi7NmcTEDqRtNkRoH7r9VsRSy15Pe78p3Vj/FGlsNvt78ZE5X/sCckLegjWaUayd/o+fv+fv7h
COxgFiJBUkAo7+1OZ1vBYWX0u0PR+XjyDBoilw7tDrn0AM//xR012pmSU5qE4bPPYcMfir5tYhpG
S96AJZwNkssMFNw/GYCMm9EVXRtePGwFjdk28Ft+ji6vC2wiQCxuG1N4M57NYgkm7JSoazWjx1co
RvDXNPHljicGRGzj1WqsTY2yGgD387d36Ket7g5BBq1Odid6uml+cR1YsC1Y0TVz6UG4fJl5vKRm
jUkIN7D1dWmIdyC83ze9EOZlLP5MmCrJBo5telb4CAIbkC4U+fPfbAZ81ObmdLS4NIcrsY4ofUpJ
JKElE2NjOr3U7eQCFsBS7e+AKQCzsW79f0E5bBhrjSHM9qi/TpbC/dpobYP7Uvb0mI4UG/D/3qYz
AMKoTa1f0ap+VIf2pefbQVZNGK2EcU6LuLMrrdELQLC2YUx+1F1pVhnfnAWAO+tKN+U4dsn0uTAb
deXSjC/AjFuc/Sf0Bg+vtzjKRXcBRZWmyOdDDjZzgyi/dnDFQzuOZC0PMeMJ4UG+OvvzUgh3jtiG
GtVsvrHHEWy5nw1E7gX3BKD+PBSGyRG9ZCSxRXhi24Kwo8gy8etNp6uDyKsyQgNsy2OSSMsAv1Hu
0iff2zftlDaMCM0ZUrsOuZZj6QnYEHJaTetuQ3l1m9Kbdx4xwXP7WvL5Evi0zkN0LoVjbgejD9x5
ltdPUCLKXffT8QTsQDzt/BpTrgtoZ+y3YFoz/MI1aXjbHaaazNitrhkj465opFripEhloFzRJIo3
tlxtxFOExuXU2kv/lVI4eIRdUBQ+VacHziiXGVwInUtfbO+2SX6o4UF76M0egpuLymz1xvjD+7eq
CEjzXLWpJ4OxOB9N1cnXGUNrHC38ufGD+o6qXIXxq00jeGq5jkdyStTU8/y67uTEe7enJp5um6kp
nS8kvHcYy1AQb/RBcnGjJmdUr42sLSbAe41UjoYHqMFrEEKhvxoKMgr70g0uFT3YccV9z6/D8wwg
jM+lsWsESAfiYa4VC6+wmMmmW3Z2FVpqyelYMAt+qNCbY9ifrR2PaUlJinr47hj4Bl5CM4XOknAM
pLp54cWTF5pxvrmS0SrXCVkVrCrPj1lJE1/TvGrDu8odIv22hhgHM/ct1IVpfMe7FxjKOR+Hr23J
3ZbYNrl1x5weQWAjbCk4g+XTkfo3ayHkhjtoA6bG/5XkKKwKNOmx+tOowloAMx1NKWrkLIGoenyC
uE46K/3rnWviFe2j0lomthziqyrc/UsZMp0MbwTZuHqPQX4HrRiZ+jw9OwfuQ3cxlaqT0qfKzRR1
xtKfjwTp63hX9lwekLUB5nCV4jY52iL4s4BS5GyDdVsegzFXcOAwkHP/vUPLRaa18QGmDi7HmaKv
nDI+JlmaYwoa936Ioko0zF5E1sH7Pts7vjKcGoXQ1EFAPDqI0+IRSJHdEHWmkMJR+/TKzd27dQmn
2y7Lbjcsm30sEvK7KoXwvQU0BOdNsukQRT8WSVDv8kFsc2UZahhT+hreYPtUjQ24H7114mZFMcSl
Up8Imx9bjINLFsPTaXBlrPuHOPF8Uxu26WZamWFFxMK0PJr3BchhDloI/CWAqZczBwyiUzTcUroN
VNM8V5mCHQXxVCiTGtX1KlvU8EDD137rAFAefESHeCaSzPLD1dT6M/1ZpPUL2AxUzF+bSDtDbAL7
0uN6NJI3kKOmm3Vk6DB1rmH9jhuieXVna9z938132rB0UgxzkoifYfVXOe2XI4435sZOUjDfAw/H
Vnll4C2BZJhXDs7j/MtaaJOy3BfKxobQyaVs+BkIiv8GG0C25ic18OKky9/kkoqmtbinYmIslx8+
otDb3gxktxMkFOPqgVVJSYAJY8Mg4Ta3g8fdBbUiPknuwAioPK6rPLHQO3+K2/e+z8PXXghuX8Hs
G2+W+Z3qKqX7gyCabfeynVlqyNX8tYFJ2ZdVOxhce3i1tBR803EQFHZuEpprJ0Rqik27M5XmHe9u
Qm5POVZRV1q/nsqPQDk+38WVe9z6iOBnNZI0pGjFEIamRh7kvsTMdppoENIjnFx0APgJKVNFoBD+
aSPg3/AHvTlBPtEc5Wt9l2spCHh/MCNxGP9QxWeyshTl8QlsE9FQzvqJX5v+Ig+nE2/+qnhlkd9J
HuLEc1UlUiC8W2NeHUGev+oB11qU5l1nOLhM8/tZO73kVrdbTrQuYCk4Huc0qAGjaTnDqiJDPdYm
jQ+FtnS7HGr5qISyAtwUYNQpTDvCCAT3MJoyfSTQzp63jswMfR5BK4hmCJf+i53d1Q4X6Ver7Iqi
Fw1SFMymKNQRNpESl82Z6vnOQVR0TDTSNNasLRlLgpd0o6mCTmfPsR5NyLlb7YABhfMKRdCzcbz3
vE7yslKQbiV4zE5J/v8x4nnOk4Eppo29nz50PleCamdgDHTCM3CX7Y/PsrSG45FbOcdeXqALvhly
EsklQY9/BYKPwAdCPXtFWDTvqct8MDopZUyx35Im5HJB9k0pJ9iubFV7hqqWXHc2JDYqLeRUKBEq
WR9xHKN6HJHdinTUweQhRGfKq9zXcV/bUgyjr4mOoNtQacetkRsmMr8HW9fFSWDI73gArNlcq3IE
y8GxJOJkixLKHh+pVcYZrY2nrzxbxwRlydiGXq4yibfU1GW4j3FQ8j0fEs/C/bB5fk7/DdsAGqlI
LAQw4phefbjSprvvWP/ftP4caIwl3lFs1uRB51K3vxGaHj2dunepyFAolJNwC1gqwavUEIMvekRV
WHF1sin6vIa5uMO6b9AfVuZO5rmDEFyaltDebIehO8GtkdJAtzxvf9vx2kQiYA/c8SnZRcK5301f
xLj0w+o8jekq++zTYzWzDaZcuoUIeZcXwwgsEu1wZ1dHSbP/3Fn563OyVtxbLDKFeGUvX6T8rH0J
9scFydGhLRGewWNKxaXCkyeCjhHUFVfwW1SUidLrxG8lCNvDQgWuEZDq1Jb1xHSHY3bGeYcOyeJK
eQUUHkDY7mJzUOsmGLKf8ElaLAmmiVsHrj2jmoHCISdhlWwreGYZfI4WoRUmodwfF6yzdZlgzadY
0OKmfUXcdTJ4bInnK2Y/qIvJ0dd+4m9K+CP63XSGvnFRnTfr8mu8mwxO0xornxn43BJWdtUeLNtN
zyYjrqpcokrv/XS76dSDBM/XbURPD6tVJCQROSdmo2Kvj+ZJTiSwWsRZSY0xNminXIE4MAVwkzAI
8NnmcJn5DEjxD4ghjtvMlxOS2mV8WSYmPYWWfa6ULLVu6ipqdM/4/qNaVWDhbQk7V+9K42cKmV2h
D4gTyJUj+tJw9AY7eAXdVXfGv9sxno84E+I8XRTwAAT/SlGl8O5OYzrenfmFC4iqg2oaxztC1flE
EiQ53C3H1qFQ9Xu334mYmO+drQoQI96qcjpducIBIoURRAHkQhWnnbtyXThh/EoxYKhz4gFl3ao8
rS9IVAUUMW7+YoDI5diZEACOr7+/bxKag7BB9K61/ZLWr5El++pDrw89cWs9erGDXyaTF9p4sdU3
otQf18Ty+MX7K5wDbSxpl4Rd9aEUpwWJMSibxj4xBb4sNoDA6DdxD4+d0xna5kjcli/cZNmkXIBu
WYEXaGkYHwS2eCo79BU1jUIAaxVvCcfgUQMvi62vGvWeO/W70XyfGx4bJD3ii4GyqaovQtzcC/lx
vFoIZB+ZF7ulTV4M6d9sDa8pFzpsybYNj3sYTeOgfvbGghRj4RmiofLgnSEeDZLN9qnQGzB6HWmW
1Dtvi/wCPmLTHazUjo8/Ye1L36y8ejB267iBl1LDkVWRK04tvoCaROJpYWaXz5jAVlBBe5TDRaN1
BTrFigWAe1pfCUridmathMNXBzngMk8GR+jJ6KJbl1kvKV9TE9ha+l9LPb8+R7xwE3T0Y/xg/SPg
ZbQG8T0Z5NCulwbBAopqhyT5ouSokju17KrOtJKjlQOg3X9ybqSzsXCkmX/+q7rhB1KhwrHEmum/
FZOod2sYEqrTqZmB2+6jkvUTTyPdOsjrCMEab4fGs9Bxcqu/eCuOkX+h+Wnz7vdNGXvW1bLY3TFL
/pqmvZVDMsJgsmZJNmPkN+tHst7H9hOvXQt/PloL66RR92xdz6RNOlIVjcX15CuBYd1ObaeBLYmg
HqCkbrITnwAgmOHjY72Hj8X8D/zzy6Qxiw0M2FHccBQc7Gjb15njbIg7mRE6DbbNLrieeUpr/Ugi
pq79hXOUDgZlFJoO1otdzHI2VnW+RkoGkBNDO7Uf1/duhf4dM90o01UT+n6mlvXWFYA0zd2bO9pP
vfybo1ArqkDj+hQmDUsD03cjk9lNMcUFpaIdWMM+7JX2QfXy3R4dmIuq2xtcPV9eY6bxBQYzkYFX
CXP7OskKuOBIR6wa7/lQc+BWXbaOT+2Zc4nIQCt6bM1wBQ+6qMg5fWjHudw3FiWnfpW+Fzs1pTN2
x2TiaLxNABSaxHLbTgpUZd57Sndp2RhTvMsS08DZfAtVcnrWWPzY2FoBr55SOobZIW1u+odt6m89
kIrW7kyPNXa7VHWRs91lkl6TSuTh5xZ+89fUB0qxj0CAtO8gyrJb6c+AvHP+C+vUvSTuRizkWsl/
SbRDtwkcvCj0n7GSKFlWiUTUILIcC6FwqqzXGrg39W7lb6VqqMeYjCsxB9u7DK8OH8Zhbu1sQanS
mUBnm/HR59EvM4jvL7L6C+fW+XvEXvXl/TQCDzcnpbQUNMOBjz3MiiuEbbcZgFhRsvjHMGIgFYmu
wCIwaxVnfU0KOu5FlsFjluqk2Zega3la5EQUxQaIIDLX0G69zDn+pJh+TJvYnwSFLyt9VjAXQu67
zcKED3Zp8syOzVUd3CLoO8sVR7f6IBdWzMNkOQS11dKMRvIo3MoP0bQh18pMNiQICkuNsyTUC+At
2JL3wYhwaIvCLFiykTUyUtB+TzdeBkV7PhyOE9aWM2tw8+JueisZ2oVvx5bA7iTRADwuzbqlBc7L
rNcMeYxznECqgzODfogatt6nxwB7t6QAkiVlWnjrKz1KBIx2bLB2HtKBO1NbATZHqxCH+hHJohWD
zLSsZZBOJBGJNSHHOmY8ZbF6+qmxlfQh2DDTBbWm8cSwUnTjVDKSg+YX0LWYgykOU0TVcGyNvyGb
UvEEQMW8nTk8yRh//DvVZ4x9IjFQRrpU0LOiJ+qUvjiFf/ly9Jhl/aSx1Yt4xv+9nHe2G3cQcfVy
z5Ier4pVlbBl86mLYTotztLSeCHQPNxArtAwTV5S22VJNSqKvaidvq1HF8EE+ipJXhP3n7jCfhme
I+UdwL/8SlM91QLEbiRA8bhwuL5R9IXsdTB8sYNg5FC0jC9Dozv5kdJP6LHQZdlJ+xyF3yl4Kan7
kDNE69KtAwDW3puDh7pZF5clZiJoevOwQEdFn/amNeODbCatrB1svIPHBUryXlxK8PVS4uCb7vOG
Nt0s199D3wtNkHq7Eh1+Ur4wkNh8CDmxYVVGipsY5OWUgJbrz3PJQX2gq+bedELoGTeGFwmrFSrY
tVIq1WRUJDYSgK8QolApupetu2RrEaRJt/tr6x/fHUa6jmqLygCMVkGz7RH0hxoUNblDvWmVRRMT
Q7qOnlMsbWOV8cKhkP1TxDh5Ly4BQHZMj26eI55L6MW45N1lL355tyadYGXDKOCsihe9/ECsnqRH
qY37QPbdy2XCHYKyO7Re5x/r1gx+i0GvJOl1v1W5Glea5a9hniD1otfXG4M/Tgrb0Cwtlci9fmgq
ZWRoqVqXCKiHTXdXjFe3CXS1xGH0FyUNweNgCBcwSBGkKedaxm0SqLBoidDQktXGBI66DdV0dabY
DBRYycDDFTEr5N7Gw6EiyqSJrHhD7qtb1EYS8/AntKfzNx9RtunHJpaWOta2EJXWZuAqdif7RUYj
xwfT7zqEGxXfIuXE3R54QPPV1k54m+le+B4KMtoc69GDoZQvvIuvRbp7p33rVmcNKsF+pnC/efeR
g4yrbgx8iOzkjBVTNWwuoU1E6AovTGVcVmBjUn/qE2rW+LDgdGFCortEqT78FaGpfpdV3hXwH1vl
A41Tw76ypUa/o8+mfv+ig5W7LgWO0vRRHi1zy2qw09ShlkkZhjyorq19KHff9DoZI2f9gZwmdRg8
Xl3Coup4E9BTL8Gha7eQiYiSDl+ajex/uRvlQChYFRqi+vgAccJ/iYOeXyAUdgfx7rLeUZN1wKmc
wcZDz9j3Ea/Lq2oEuBuqkLImrCL0/wZnbbw5QjvL6MZan97qEyBV1K82qRcJFs/9x8biUKTWCYKr
XEwY6yTybpa+hiFmphqhMaNMDzk01Y0l3UlW1VT99mmSpbYYZSJuXXE2Gv2hxEVVQI9tV+VzWbGu
lRdJlhONrHzhjuD6JXfOyUEyUHEl5jYMYfZ56Ie/JRQw0S3iwFknpOwgDykVRkvEZsDVtMD8c+qK
YIQmoS+G5Pzvi61HSetNkorPG2/e8y9/46V5RxMZdYNbEa1vZ6X18+/K4EaQp+b1wDjrNqo13LUl
c3/udzugExHCdQwVn/DY+G5KtgIFuA+5k9MMpJjfm1LvScAWEW5FG+gYk2GeRM4Uz2bAfb5oRp9r
lGE09xDTcM6h0GIWEJJ3Qsx98O9maxP2qCcsN36n1hB5rq3k4w/8lzMj7CWlJfIr/Yc7uyKL4Qey
bl+4lc6UNYkLdCLL/J6c9mXvzFy1flYDidF4sPHGDxh7kg/iYi61s3VeZzJSQV/vPNjepPQTKZuz
KfEJbxq1pjGATSaKtF0MSEuNvDKy2p+bcN0k6wepfpk7IFEsmKjmB6w/QHqJfcmYJZQKmlcxrTmF
2wIc5nJu5Syn5lubwBiAA8iynktY0Xwp6j+7zXkvpHmGHdt3cpnPtsc9tUEqyVAfmkjvNbf2fbdb
jX9BfI9jQSbsJSR2NdKdQ2zf1kL3ItVG9pizcm0KRcK81xWTRXRY2L90SI7gI3Nov2MNm+rempm6
c3ebVM/NcDO/U4lKb+P64c/YRyRB8zExvZMvBPQyje3KKG27+Q31iQMUt7tX6JRujCWKRA4V5sSB
2txP/9zZnTat+93ZM7aC+a/hinEBGed2GJlsCudDevtV9Vu1hLeTgpSXDi0RC5x8uoMymPwlC2hN
2wgJg1Ikkvmn+L4Wn8rp6zbHasAA9cho+J3kiSqs9E629+4LXepwKFYWSgAUNMulUw7IuWu58EDe
e1RpbDsNnj9+jUxpLUoYbtNfHPAkj9WEQXwnoZD6AoHwgoGMioCTmP3lJW5Igb5Cmuair8dlYLQh
zhO3Lr8QKrX1Js/B79eosofdTVD+BKqTI4wUDGtLXijAj+n5chXJF/ICrBj5trMwoAYUX77VO6wa
JBkhg1cdikEIgd+QSeR+e6EeTrXqX1WbZiIxpzeR5GFhzcsJdAFwwWIKBXGv3I3thzlElp8za0x8
MtVfpK4JlTNffad8IJBEn5VIMB+zEiBuaTYXy8o0rCbRbsId/Q0RoMMnAK3I/5ykIBnjNNT2A9We
jRd1EofzyhL7ccZrxrCD1cxHbXKvcgp9ZqpACmJxamOEY9DE7uuAyIsv9yBND/wx2I3yh3YK1McM
EywHLgI2clTl9wTLOpsAMBqRDSgahbxrjyssQC/3Y8sXNTohK4NOG48wdBBB6jtl0snCREKIEOWD
HdL3jjevWMOuE3V/c7I0U0EGenK8VROV670eLDl4UdT8VKyRQQyveS1DEW/6eecKGTe0p5nHVU1X
0q1ZiYFas7gSSJhg8NGWar84JsW8+nPKebtCvz0aveCErxED9oe9jDQKNN+olWKGQRSvlmPgeyJA
wmw6L9gsYoiEuB9uenoZAcJsoQhPsqtNDJIHYhaXB988pC8jQuhhMfmB9GyDqxiTE0q7cL+Xnl/r
dh9XrA1tq+uw6Qc9J6ThnQlEX/e2Ce/XXiV5f+I8qNu77t3GuSHdELHpb1QYJMEoKRUEo2VtFIjr
+NUFiu26E1/MdgzUN9GG1o7ClWIxJPyo/WoSu1WMCEqv0gr1X+aIXfbOdLSRalRvDp4bqiBuXVGt
OpEkW3pbPJuSWE4HAXXaFZFon+fjL8pX6Y0gE8exhrM1u3GYwlLvIqmuiDGWTvjz/CulLG1d9lRF
IdUqzs769ArWHxDa0y2o1wH3j95325z8gBceGJvbCGn4PeQFUBXJdBIIvsXesA+vXNEJDzN6Zjuh
hkLgul/Fbnsp/zOW3BnXvLAk1Ni73Hg60FM5quLqrFYrH/fgGAs3+p9ClZ4d/GuKyXNFneBzmNk8
gd2kC7tPl7P2KKKB6knsJg6f7cJF78JqRsrIGNMHHZoes60I+jKvRQ6501VlYyXOGXfxE/jwJGrN
JGfj2IJd9qMhyQsh3/h6AyT6a/oXqDgD/miA7YytSNM+azZiVZU/rHvtBESgUX73Wv2oI3nJfLK8
Hxushn8Ma+alWn8sqJcSyRs0nvTNCbKclZoxb/MJQC4qNW1PS0wBPmfIU2JHgw4NriCQ1qFrOwWU
5qvrj3ibYUlKamLRedKL+tcBa77uIktX2sEioeGPRfTUAuUt2wpCFvTA6Gs+gvpiotEcprDPPToT
jmQNvj0koy5n6HARltQajJevgm1d6KDQgbBKFXLCEROhytjP6omX7lFjWxv7dlMqahw0+GHOY3oK
/32PmpDnrW0qEei7UGdMtPEbh1vs9k6+9WigKD4yHG2MDT0E+nfLFnb793ttsdjm1CL2pFre7E9M
jmpWjVeMf2StHgDKvr5kDWuaLR6ftrjEeiZCG9mgBR+aMz/lNemoEg31GZelihTd+3cStFDtqcWc
kVPFqusbNktxiwUjbLjJvbqAc8IMlzlkXyBttIyhfqw2wKnEtuuRVo03Bx8DxSOf1Qds/tVQx7wC
nlHKK/ZwJlF659xLOOTb9hq3G3VIz1nZp+M67wj42yQppTlerOn3PfUROXT33ArtxcUczbiWk67Q
RXUJ2lI84xhKCPr3M7gVqJFxmj+Ip3W0CowXX/Pc9VboshYsubvaDtS1lw9tNnpz6cgQYigr6AP+
yWIHMUF3gwxy+xz3eWD6rLNl7UhUi7OulZDwl79G5pnU2y6XfweMX/bTNCaqBtuq/UdQqbUUhTcz
KFLGlj0nbZGG3vCZ480KCjNiRilzW9hL3dwemTkwNEPNTCKSJm3LvMISyA6mQW4V9evP1tm1GnuI
4oUSl6dJihK84RzzfhkPN8PWHi1nzSL5sBZP/f6I0ykM+IICxHHuhYV4YHtGtQyidhu3YXW7PoXz
y1K22S6yQpUNQf4xvk7D8F5v7l2BixeFONeZAbJdGJLnLPKSndK5Pto5ApXMF4U8pcJhS7+E9+3i
ZvuHsLYxlYPnz6QsyFXdeeMPbiy95fPLj3Wk0v2j4NyChUgeD8IRMm1OFRo8sZOqmGTptfIhbntV
7huSFkkkalvDYj+JXAOwxdM+Mrvkopv6akATfZakdeTfQHiUnTFIdlwERzK3UTTbZUnPs35cPhJv
s7eZ+Tkn0Mv+ZQME61te8AAXSioND6ZGyDkJED33qqQwP0PKHuxO1KI4HByQiklNUYS4sx/CM470
zEfQkRyHf2p90Cd5LMKlF4KDOQd9TQgdNChQ1xRD6AJ2sC4vvFXQg0M4X2fmAT+NTmLX/bMpb+wy
z05Qtpm5Wl2XB+O3la3nlne5RyX3b7mpXw7TZh3fozT8lKBwOkI5gclHyTBOx569v7SYCx9VR2un
1ksYPdFEMlQrtmWr7Mhi682Hyj57ycLs4OP71mmavY5f+LTdx8DogdIEzktBBnNwBDqihsEhcDYZ
uEg7Z+zZRuEQVUbBidhOA0HN0TSGGPXkpHZYB7ZppKXXWitR+GcqGra59k1RABcJx+lGuEDbZcNf
leFwRvzRsL3mlnsB8gh+SGFn687OlfYOvCXik343T79yXOxnEWqT78Y8/dnufzZ9Y7A7dNIWbsre
nAkDZrb9LtEYMgbx6qRsW8wQKp94GXP56fJRE7u6bAdrZ9CZbiWtIdgMQCwFy/amHoND+JYSFziD
eYszFkgfmrhgrY9Vz6RexaoIJF5ZeDIlwQ2SuXn9bCexxkiDJZ2nj0P0A1gr3aWZ6qWNP+Sl9aG6
BL7zc6zm0baTaUJYkGrfOadybo9qEfdxAQTy82VWHy0Xn3iDlUNbOwVmjf/ORyQW9wm6/TU7YrSY
cGalJLD1qJ4fqR9UvbgAs11uxwItirTYj7beFoiirxv7V10qhCb8arpFnoPxTn5pKsUMeq8YT3eC
rk5j9YZf7WqXYUfrqxcm0+/439wMhhjc45BB6pZAuGLEKTKrkODe2YcJ7oYVwGdwNd6Bg/uGf8x1
lDh7FdYccDYcy1jXLAGMQDyxtDtM4pjsDrpJ4RBzw77/n1P2aGv9z+z7Kr5RsnkmW+IU/erjWsgB
Rv4WllNba9DNsobp/yeBNxaoRCIRPR6yev/PHdg6g9udxN0bBDytWvM4yNTHcScorXFlrXT280Xb
iMe4ALubFIn8l+DM2sayNeN86L5KyY0/u2mPMTcEhgB7TGUYm1C5Q7tr+2T4w9GcRgptAlKsUAFk
NKzy1lZKcoxUDxLstgIbeKwy9MFVJCsKKwsP/WGZGRI5uuCkzVdUTCqkoLMtTLBtxaXHDivTlsxK
1zXL2I7+c398TM+9DWEarl3bullv2mWrTcqBQVUx+Q3nfTQ+hvrXFVDupC9EsTN4Lt8SGBXNjgBM
BnuUCUT8h5pJYU3SGtPPPB75JORirPVba454Xovnvurj3oY0ZSWm64Hg2q4/p9av3KvShbC7GGlR
04xDMaBASa75WrLZn8RlWNA0zi2NJdCt86SlcUMKcP2UwF3181VRuivfAHQ+bqxj02NCmffkvkPt
r91BkufSvWn/jq0f+ahlzA1N6T77Ol5MQnE4PrugkB6+hxuZxb0Hr9k8ZxWiymBWEwsveFUB1m/H
gs+K2LB+IOKeQhBySmS9oGFPAQiL0q0UaJeLrVw8eKk5qKTxOVEoRLQCrRsKRIeEpwdItsh6Mos7
W78dpnHSd8ZQk8FUwiz0W32D2la0uMEOh/Kbw4v0iJIReOF/vhFcCQxdsEL76gw71t4v7HKz0Ppn
NKjGul3yfUmjVioSdheHG/gHuD+qCM+QOoPJWCG8LxVbOe0StDjhsbO2wDQHOOBagPKfwlIfjEGd
31l2PYHFHiWCC78uLstVm8vMgHDkdCOPE8zaM2KtT+dQMXKFpNwInKAh1JlX803eMm0kIgNbmWYD
0tgE9JmBOSlFilHOxDc5RvCHq/G+Jc+Ped4+LpcLQwi3ufJYS3J29C13p1oupukpoBBmGw4BnBJm
nEKO5iKrfgOqC5sC/JVO3YuXJ49yI/R89a8EaUqx+aeD0n6CUqHj/4ONrDTHh2dNY82s6lgpGgZA
z6+n1Qwf4wKbolSWfu29Olgqmk3bR3HjCPRq55ArRWhkwgzYfztaUeqMbiaV4xvwUV6xWahZJumn
mjrXWEN7vr3cCVwNpv7sng7oBMPKEAyI0R9d/WlUMVKUn7M9c47P/cIJPW0hRlUrUb0yDFJ1k19l
KJ1LvI1Kg7t/YMjvDP429sGSC7E/eRZ5q7LoAbsgTgwpGDwFziF4358w2DffhQxhrT19kg469AGO
otw44OXqd19PFrDmaTBmFUcIjvZ6KxOGttJE6lnG98PZfKca4p299CfZyAyCkHSIDqgV2bWERfRn
ehrlAAZjHT7sFIYcIYQsnYjPShxv52L3PXSLXSiy6Y4x0mbHg1Clc8HvmN3QzBxB067XvpXRhgfy
ap1IQln+D2hDDndXtmWq+TCQBHEO/ZagZhbHBEGIEr3myr0wIK6zO/9wrO/AsMU+vL58uqZoeEJ5
x8sejzeAGqSZ6Sl9PUB76ZmquOtFNtwphOJbxL2nQfBngsbAp+o26tKOyhqAOs4lJfAnTUmXR8qA
pqP3wyIQ7yiEgk23M2xRDZ0wz8lmlj3ZAy4iZkpDlyfsYOSeAyzI5paUTPBjsukCb3XKxtdqOijV
GyvqNvkFXuHMyf5CPA05YrCQQWWAUQMAitMJAJqErJTKQxBu8Byn2SUnz5FhbLv53zcfQACButwU
nv2IkgSIhi70TPg9e7c1Te7nnh9jdLx2+MbNJbCVxLUzjjxzslkMGdBWTJLkRWVulBSndyWrGABo
f5VXEPnIJTN3Wa2lv7WT7xaa5fSf+9weaP26/8GPYTacIyUNpKJKjLrN8z+GILlbmhDaIPaCDg/g
U3jWC71CiATar+73i3wE32W3nXipSET2V8BhOYcaYd5EtXIFblozFYbCmQYIxbWSzZJHphjlfBOd
N4Z8Ic5NpIb8NOVc21xqVr4E+deuJ7lULuQy45sQAk9R8QOPK+qLFQRCWpX30mSgNcQAB65Gt2bE
CGjxhV9/OCQXrULy+motMqR+ZwH5iroMhGzg26pldxJ3ZRT++i3m5LHFDLw7nv5NpYyOEL9z/2TN
jWX9q0stQDY26obRnh4uHVFrl5W/ZWA5IecaXQ4vynp0O6BwXo0XFPZuRYHsWPF/JR2ewKDN4DwL
/aC6JsUuCSjTHEK4VK3/FhLHxlR+1mWbbNJBisUv2HYF+NZa1MB13sD/rurs85LPrnju4WtceVrx
JOT7VyuSm8SpkssCkDhblzWFqYjF7ZExTI5nsOr67P/MqJFINjDpkEubHRJMWitX5UH9p5RzXz6H
FuhyWtAei0mSzBZPv8F+QE/55CGg0TxEj57odVVxCyvdh5r2/GdG3NedtBT7aNSD/cN0vbEHb/wW
4GG3t/Hz0Zg4Tt2VmrjVyqOHr9FqFiXKI682rwB7zRajheb7gkklpYyID6hwKw0dzw4JTJeEQHvj
RCqQA6tzBXkLS8HGiA/oJY8rpUxbPtOjpEQSjTdtWHMLeUQqhE6mpP/HIPfptptJ+Vj+OLKs2veM
jWx5lmAdaavA4qnsaSeSoI+kbwOSzP9xxD7/tjaj18cR55SVpA0tLPNA54TNAbT5LXQ19m5PzsFj
pYQVi4tQN3OQ0ofLbr+sBIhcFqPSdLW0Zu87ts7Ci7IheQY0ibEux1R1EZH+QGJinOWWDvssRi2a
2lud7Pg581Qd4a7xqj/Rw+p40DfhG060soZ5ivItm4MKN2mh6A3Bngwq2RYcc2c1GhzsiPDrzlCN
feLaoLNUDoqFt6MoLobkNJ9+m50QXbtLKgMxoAgZkfrpIEZqPJKVUjKGfO6PAhjuhGOM4sz5xdxx
l7IklQDpS8LKT7AdGT4sWNqxuhrAClJhcfwPUF6W1iHMWgS+2bmRMWwJcJy7h28Hgcw8mEkZ8icJ
pYxxdPiXx4FkYFbCPoo+HjdmBKnqKos544V2Ze+vbV8QX9Hoe9Qf3iKI5wtLWggkoOsJvSI7YVvM
7jxgiXEH2jnJse++UNIwd9pDJmQnDP4jQU96oq+aKhg/9eowpX7+CYLhUWCvS9F0Jkcye23IKfCj
RlAcd7o7NeXrktk+GiB4KnCIDe0cqvpImvem0Vqj1f9die7YocWrh6bks0NgAvibzNTNZP7Rshhf
x1bS0G6Hcc96BD0/hFHzF31A9Rla6AM214K0VQlsI6wbylhyVFCeh+V7VLImKfl9yeNT6vQO85Yb
NimFQHSoLpL69GEqlPkQl8m1oQJ0DkUm8jzB2M/1K9pNUscttmrp1eoMDyk7HcdnFj7k68YmOVeF
NIc1kkmbyqh+Pq5F3rbQVC4D62QH9pouDFM+YNO/DtyUEAWaA/ArLnyj9BCfHVNHmCzQuGXI+Zzi
PCTCl01FLsTvlKrVHReSrgi3xnaq0pPKAP38ZDPEhsO9dAfNPpQE9Bj7lMas3lIwHr+du+mOOUJ6
YuMswK31a5ddq04KoGlM+s1Fl1NFfIyAHF2AMYckvzlzStqSKnjNxdRW6OFHmkFHpDvm6sSj9ax6
tGPnNM9sPSpY7bow45dDG2c9rY/PWHfEIm2toq0oeINBqn+EktvLOEk2BsLzXBxvlZZWYSjJ51e6
gODNySRg/lL/VQ+31Y9emKw3Bto/mMyUEwr8pP9G0r9ab40z/0XwkFsNI7nLNhNSmgkmYPm75RIm
lHB8RyU1CLpdbZjv5DMmtQ+W7tgb5cInRCMEj8OlhkjVl7JQIMco5EerDAY/uKHOiqHaIq0Pfy+B
hoNPnhE1Y+Pgi8ZsM7m1OwndYC/Gfl5GDL8CAM2GDFGLhooOCeh8nmQwnbwlFBLkiTacPGpGpKZY
reL05a/XNkRsS446NvLxDm1YX8JTDXbwwjM4+j63pdkN3g8UNI7LDuqvSmJuEKzE6Jw/kFLqvHLI
mxL5gDQm2bs5vQ5ktHjVF1TCEHdh4uH4aoqGAmh8CptOSGd4jx9bpCP1IIVnCLOIZscD2aikiv0U
x54JuduY1NisZFo6SQxNqMuMw/BoK0atj73u/o+G48iwFSB5YqqOWwqdHnQfFAF2ev1WJnJXbyw1
BHIm2Ea6OigJtdBDCk1NpU966Z34XLQ07gvQUD2QaJ8nB4uM0oP/mSm5NvFF8xjjv8vePH6/Z5Pw
O/agWAhNFIRFKZbdlJJyDBkXoK4xKl6X47rNi0j00OFRIqN8KoB9r8uh0slCmDdPugvxdFTGyIFf
rTD7DjeNzgWxFn7uQEM81qndyzyvCZdBY1DRw//Lt62wHfAvK5WevZRfgBq6dqyfTm5/hKPGC0qH
XPf+Q2LzCSopWY7yMcvHwL4g7sMyzkPTgXAIwmrmZVIq6USIXNwoaGxQGRrroaxQ3aNM/oTOXFGc
BVROjIKv8ozdg8Unumk9HEaQ3TakoKkXoBNFDpUcu3T9wYr++nC3BAjHmFk9IGUHXAQ7DFy508mf
M21wZ2K4ZfxPGtbdC8LmlfU8BdtfBl8TY2G3wvNMtXQrfHUOeA+ILVIW0UoXm0YbfeRUPEZLhxtu
No1hiMyjEfim9j5aX9ouvbnMjzRD5fMhBawfDBEbU2sxuX7sy0ALyGZd1+Ksww+j7Y7Ffa25xNQW
5hIjkmAar/P68O8o6YM4lAV/zFi6ytyfqbVV9cnCjYLM30NkKh3A7vt+6BMMWfNjDyQ+eMo9XWqo
8hxb68/S4i4Sr6PEJyKtObluW5D6dB22yoy3J9biLnlisYl4oFnaGhAP+5jWkFxz4SDU2VK4JuHz
UiWdUHdAzSF6xX6q/KajUw5YbOjEU08QTkyNsyDQL4oJfsv/TUgBh4Vv7lR/o9GuwyMifqw5AGyb
1/21eTEqrMq2yrm3KLp0hYu4x/AvY/fVdb6T/FqQKm0PONH33v/LsEWXGqWNmRgJgfziMs9of/ft
GC3yn+YVwaFpWzHRBZxHms2x23OFaJ7c5OjI2QCJ/MnKl0Tf9uDTCV21d35q2LLNg2vsozbKx2va
hANe4OUctzctJNjze/ga8Kiflqq+1GIEIta0jGuXNYpOi7ZMBNplLViTRMPFg0l1L978BB6USdVs
ewecJDBSzMEuZHDnNWzWvHfPU0FLYhR/5s+/iwqFFTyIp5Ds2JuRnO7JuFu72Z3Ma31HNPqWX+wd
c41VnDEVQpXqdoQlh5xoSFgO6TChxk6t2y4FjFb5MCok4rQbx6eQjO1LPLFugOt11zOyJ8VuGNuv
SY/05JniITLtXQKl+gmLYuccZUWRsN+lTtnOhHcaG9RFsMQAWRvxJrVBbjC7h0roDgC7c9GLk9c7
DpLfLVokCvMUoODVwsCHH/dWyn0eJ5Cr7U86t+i5okF1loMU6x5hessGB+1xpqqyAC/fzvmKmvPM
BgnKW1WoSJB36lOmGRpxpWDjILVgVYagncLZ0cJzv6yXeJegnkrqGEJpf9FkAaZuCB/3OKOn1xpy
vxNoAf4bWY/mXtFHQ+DbqSvy9KgmrM4/+qra1W8wIInf2zTG9Z7bEAB0/IaNb3pVItD2KQTnc3+1
6y3H0VmlIf5QF4ViOrnqD/oAw/ZCjVzTzfPUF4m/YK57gdfxEiBj1staEfFN/CvBgbZKnEQIxStg
nzsYCB7+xC7hyxEvunLhvQwhMUNMrPMv7FyYUkxAoN+bnh5vFM4C5Uva6XDOG3GUGKIC2ka/WRRz
W5Q9R32ozlme+f5cy2XkwwFXKErrqN7Mkum5m48TjGFekdWq9cZB2SMUKNuaxiJYIUdrMUKuyKP4
VTebOOASgzz+xWUP7PT4Lh7QsLR2U82+KlDMf2t1ej+9bX0ELbDZOXP4d4GaFSQ4BCOht4b68iv8
Qp5OBQEmLNRKhCcjshe5WxM7AarnJ8KwdkRbIFIJqzL4FV/wfyuO8/fIE1tDGBNrxKnXo2IHZJp1
RrLRMNKzv3/9myFZuhBoNxm9PfeyjFgiLMteJPsE/1q6f7Nu3Gb5o+QNd4VeYKrGMiU+ehaJ5DWN
fXp29KHOjiUwyb4whJ21Kfxb5zTMJYFoUA7ElrUNRkae4hVq127a9G+R+UMDfjPWMl9E3YIBL9xR
KTlRk21OXXi24gbvoatDL95C6aFodyFA0RosFOgw1yg/ht6abosaTvpt7vOFC1bg1SpoCaZzSLW9
o99OxPLTnGvzlARmLNlapm77WcSSJxbgBRSXXFmq1VyHQ+1rftQsK4Dhl4drE/3aT5Oer14V5kfd
qPvppNXCobPby/F0xH3JVyOjz0iHcxsyxhjscnJ4l04SIHjoK4oO9oRTpGgtmYxropVqm8reAC5V
6Xxj4nYvtXVISr/tjskpyofW3BUbttSxMYeAfVw7VEjPxejvK+YaU+P/jEwGEVOAiO5KY6ve3IBN
fmqhAd0ls1WUXRO1PNdkXuSiBOsjkoXapJAHyydqm6HmviekDVhNB9buXgDS7/FiKOu02zx/iCZq
Bc3lAbhhHNG/+pCC8JMA1NHY3UvsFFxwbD/M93fGS4RS6ctbNc/agajVEe5faPLr8pInq2Uju1Jq
rqEkTSSgLX3hJ1wplbi4hpKHpXtwjfh69aAlG1PJkQYEOUt4sVg5Pch1D+2Au2XHpjs6m+NytYJW
CtxCLGZ6aB0qYG3twVyIVX3Qn2j1d52TIOUTGTP1aliXseJ6C6kCpcHplFpXjUrKhUiCYsDdAyrq
P0XyygWeZkt2HkOymXTa3aIEx98I6B5gtvu2Pnxxrxz0TXer3ekSt/KQO5ArGDu5lqTHhcsFsRfz
QNe+55iK/dHzKoht8zN3gVk7FsjH/F/2pBibzc7Z5Kt1/urUKaWY1SuHCobc+j8vMCShhyurdsUK
1GkAseO/rUXnSAgM7hGz+yTyvABguFLrX5tFW0RhtI0/eihiyseBEbuVBO21D9SVemTDUlupaPmR
hjQ5kJiAcbii4PRKy4lymSyn3kCrUd3D7XZ3VvB/J4AUcnC9oMtBvD+WA9ykVMx9PpDleD19VleA
eQ72eaI7JzCAJEtJXrc1ZsC8Ct28D/IIkxMQaYGoCGB38BUBJzNg7HL0v0ssSWe55/wjmLXCTi6L
1ggjg+/Litlej5AYy5WwNlnzewKUcNXtf0qHO3ZNAuYDSwoDaozQFaFcVhqOL0JxeKifk+XYOLsi
3+ZtcPa1VIGuMpzYE04/nzZ7oOJhszaCZwY4DRU9Yoi6aFaHSvwnwTSVis/x6RJTN7WKRuanyLU1
8F0kJzOZ9hUrLhV9xAkmH9gx8rG7CxTwbay71ZoWY8GudaITPq9FXQLQkw7zcPqG8nnU+uTmAiyQ
jpYXXRVxm0B2xlZ6gagBErQTTrkVc51Dbqn79KNSVARc+Tksa0FlXNMTXG9qtvZLcOygQyABOY1g
eYUBWiIi0mo7R40X7t8Q9aMpgL6NsUjQStjMfVTIkFSIaX9WPNQ3mEnLQX7IXhzwAtR6C63yjMKQ
URlQIbXyLSLPnu5DSAMffPqCtInpvcQtCR/5d8Np4SNoJq2G4TJkutIBNuxshT+Vw7LGgR8GHZWM
AdOo9ILpoxUMkaWH55gZ1HlA+gC9gZJxMPEtKm9VT5/1+2ZbTNLfkwyz12i9WPGgSoOz4+0se5BM
thsxGJ1bc1uLRBYhRY/Ane+Wx+mEVBVxHp4bl9NdvLtpWUKwFBJ0zTTcMMUHac+3v30dm/b8R3QW
fVyCrWmenL26m++cYandV6JigTIWshLRHlVjkhkuvUErWGhm/k3JvU0T8m0Qzuc49NztqBnFRyYN
BRCbMKtwZcTVuj78uMILS+3cbE1MmPUoZTElYPDoauUrTuMEhWro/rNes5CC5gKu5QzyOFIMvYIb
QtvirhkteOlQaNbX6RVKuI1PVcmGSFFndE9vmDCZVYoMJ62YKNADymGaeFnsBBvv7MhVYbNcKyo+
s1mpUxp6MySVYS1n5PfPWLhS841SHv+4EQG2ZXXC76CGx2TxViHbR1s+0MJ9nK6HgzfTQJpeCR2/
wvYoq9wtqKPKV+Hq65sG+aVO3fM0FKKTsWYjGIJOzGLTXRFhQnjnpQhbJ47dD1NpnhaznQ9GGCLb
6JmhOLko/dZpDurYJlkbWYNIwTrqw4VZ4NB9gnzTqfFQhjsAObiFgKQncfiySGF6rTU8Xl4JXTlt
onULcDjL4gEfHR4ry3Rbz/68hz4zpPKYvrFSdI2chk6q4LEAsqP/YVrZGRRw5+T2UegRx+yBgFTp
HgXMFlxYHSMg0PQkQ2SiwUDPxV8w76FaxiDyD1HgnKicuVg3BcDva2jGVEMSoJpKz6G/UzdEALs5
hkwOuwW5Dhj5620DqSpt+3iJqiY8NrnYsB/NOIMVYFjNeONbllwjqFocf37FNpmD26+lvMOeD/MB
J1ILM8PoVhQ9pFgskmA9lWUGg/zadYpDbbv9qvFE7aMDD2EaZiQj2hD60XDs1+DD7qpDXTuIhZhi
pkr2aMh/bFyTEQzBd0ECTfjI088oxCnfe5JmBkRSrPd50CHrB64GFPykwUuOGbCiNQ3A4TBQC305
Pxxt4DqQiBz1Mj2fir1a6Jwy98B1lsq2Vc+8Wt210IunfF9Hxh0UG5ScMjngOmfPVp8jNTDElSex
QP1RRrB3qbOs6qU3VxLWNxjBxbwc51X56/KIhurxM4e2EVqe/cI+jF6eUBh1KfXqeXhwvM97l42h
unlU7naAn7pmENUUS9ZqQoT82RvoWnBYScvgR0S447MuuP/t3BM1/swT5Ygp8+sTvZ8OYoGnEMmo
riG0bGEGwSGbP2K5TgNqKVY0XLEcBSVLrbpFUAfW/HV4uo4fOE5olDaKx5cmZYn4RnxotEJWPrl7
XTrhO3oM8fZ+kuMVtFttBGrrzpjBNn2ZHjsH65EPvDmGLTaAjTwBX0Sw4QNyHnNQznxbVvif/0YU
P/gwIytyzLQaMM52fHp7Z/jsSFOd1SEL0SDz7SfVa9TYnk9d+Y9/K7icXwf9lQyQKQhG9kRbzFfL
Dp6/4+ub0wxjG06BTFEbY2hch9a2YgIac5l9DYliUoslmsLG3SkpYN13JHRin0u8Ki6aXJWMeVek
flXcBU+O0u/nW74t/PL6BG1gEkthd1kIyskJ9Z34mZMgJ2sFKWIU/Sx+9NgtT5VzlM1lmYaa1orn
ULU4b/pZmqqje9IKRYpgelMe+H3qw9L8qrU//W/olbTfK/2nXzQG2wVF4xT+eqPaVDrW2Ts5rIzQ
DLdIuT6f8gnC9PevKfrBE5tUiF/rnMtVhVZPVR5XlgKWqELzZal9DuRcre3AxEebUtsI7Nlly0Ps
q7JVfL6l3IWKISyd9qRc3rAp9ezk9uRTMXI1nqhKH8IulMv/bFZG2VVuKWorDXqtm/MKRBLqrZyI
6u3eC8ya2RBw1KNlOkAUZGHVzrImZ1/hNh5jqczXalcPp3r38+yTym/TDVB6aJ2TQ/Oc4F9pCjTu
lgtLrN8Obw8wwLjpVOlnzoIN7WRcq2TXgqZsDkjNx1/5deKjkbh2yvCc0FM5Zf+Xw6RW3qYG8Dg1
tApB/2KgusPUWBxnKwaLm+rcqgFnfPVlQwwr+77BKk7h5vO4tkGKh1Z+6Y2FWSxrQTtbEXclo9tF
2tOLW/oRRqZCo1nBgDh6rBjU49NFIRgX1s/lFuAmc+azvd/nvmZXq5BCD4oXp1rN7PULGDM17Ksb
q3eD2t7K5HE2pgt1J1Tnf4jxsN9MfBnWuk3DtPPAm+m4XRM3OoQPHL2xILKm0P2ind/xriN9DKWd
5l/oz/KWOuDIFuDeIDi/TI8qpOBXgsjN1Acl/kYNQuGyRB598nxhPaMaWurG6fRib6J94Iba/5Mr
vHNOOIS8aJTFvfZMWsTxL1B7W70w6SoMADmE8IfeCSDtp2lhQPMeRofbb2049+iXqTkEhFcJ5Y1F
9L0ygEoDx430B8pjcmg3xjpIDWn8U4VZm6h5IUKhHyTdgDLfdQWSnXqzOX6SRt1Ck5WcJ8VwRPLX
0LDJGJk4aJPQyRR9AKKtZdlW0I819upo2db/4WtvAWuA6bqLu2h0rg+s62F98zqT2QAG4xSq9Xa7
xkTPtRSZIVhGx4PZSMQKodVj0yFBD+OZ9cc0tCAGDfqQ9yyutbb0M5FeJpUyY6an1P4KTdN2/+vL
dct0kiRWCMD78LU0IgI2/uQutdtCnbFg7uFcJZUFKK95U2pDFqtckzSKe7a1lEu9tgfordLmjInz
Nvq63IAzmYDoMt2U3I2hIXxA7ifQR++9BqLWXqaNBKsEQ2mRKXGMbcX8Gg00azUDOIUNS7oOJMKp
P9MoIFEgoK0MMZoajZ39a2buOzlMUD9lBbEsn8mPPGYlbJixzJ+SEONy1cqcn3EYLqiy0IriYX96
vqPQDNKIhRGcg5XPmwey4ZVPyRfccXN8bYSGTu2v3ALY1K83n7ZoNerphxVprzPWwU71O1JyIxVZ
Nry/laSG9m6I+v2hiLxh9T0gArG/P2mGk3d+hzQzV1zy2P5DfcMO/JYvq1F6jO4UeQ/Nnq92oLv+
22Xarkcul2ImlXXLHVA1Gia2N44CHAVC9DoUxuw8oltq/BYvpKyAEpEhcynRcejszJU2L2sj5Wz0
WZkeO5fUb6D8OMhF2uqje1ZCMzLXlsCN2XD3DGyA556rc6ipRB/1hH8IpjXiWoJUyCnASIypn9Ch
WlB+ax/1ideZJIihKiiLXhJV/aUJSiqG6+fsYNlic9+6Th4QYqMLs2V2fs/cMJM4U9Io2O7I6uBF
OhtqAbO2ptdYzn+yR0+OqId/8QNMmFcmTtc0zwyynz9fY0dOYSSIFG1QaLKlkJVoKQb3xtPKgBHR
trJ7PcuorfBffW99OAPR2V9WMKnTnaAIzPo6bRWkMuS3uaOOL0jOtWTFpJS0nanXv4CSuiCFsblA
TR4EaNnb07GOhv0ECbsS5Dl81RsOFVcIULO3YQb3lrLdIvysgakT/FBGvrTiOa7bYOpuFLN/dduc
3XXOgSVJk2v5Ex6WqlCFTL+P1VuYhNKqJKh4d2xuROlM7V7ciXvbLgzpq+9DNwEPGjkSq274VAZT
kvy+HjFlTvnKKu8y+4AsB0hnAnbDbTWW+R/TIoFKMamP3k3TNTFBCrxfTlp/Kzbeudt6AR4FYnU9
Bx3pm6L3d9DxGPriSG/nlhyrd/EXgxKVJx2zeB+wQdvvGUciL1TRBMhGaPvJM60o+qZdX7NcP1fz
cvmziCoN1c023GQJA+ybNDJSfOExyJ48IYe2JCsoELNIqxd6YO+BdjkrMWjUjqaUeZsp7X5RfxY5
M8zC85w8+0rAvZVVV0G0VnNiCbGdNglodN8mzPY+g72XBhyuScgIfBS61onu5wvrdlGzQV5iannJ
qkT9xUv1wPaxDccz3Qj3NgIvJtf12nZRx0DTgnXL+Onu3dZv4q8+wlqleUHxejmMyp/0VrWI/OLl
sovUYxsYHR4sCSmbq5p1qt5Y06WbLzCS+bHRC+OXNSAFiLoL+ivt0Q9nVe5SZlxq6hK7YmYNIpN0
SpOgj4v/yDc/ce9EHH4EWg5VoruLYqz2kyW/u94z3CF0aa3AZxBUitwvhJW0DVAFxR5GupD1h0Ts
wDEx9+CFZoRXuXJZ9sOOweg7wewOvrhHAqZoumHKEhQSFPcIaUGxo0OMhuKroqGltnX38SRoQYN4
zTeMiDg1jnYPBV4m5H+KswGg4cCGtoXqT3y9ZfsGPqYfjxxYMxSboNwLqCr7pkGsOp65yV0Q+xHU
35fEwBn+Jl4zKlyKli1pA15mXMI7sZa8nagjQejzbGsC+HNOWydEFjRKdpfTHjd/tPXP4ngn/Fve
2OxqcAoXVB5mz7om198JCryLKjLCwDsmGONArEdhKxOGtVvWypseLB/hNbBv+wc3wndhb3EFd72x
nEWBNkWqVJ2eQsmtJWN0k+iD+4haMfFfchOlN7cNuvm8JBJrX0d6hI1eZUhqiSDyEl0Zdjli6HTs
ZlYPnQSJBlITGS6f2p7i2vV1rRUYcMOU8Aq4W86Xde+qKXr9sLynDnKmGmf+SvR+vwoGTiYLqSTb
ffzd6h6i9Agq1FKz2F++EjjoemBS9A81zfwfhJVbPpduFdTcdA93e+BWbqbGKC2VfJr5lypqOjyM
QwD3q8v2KLuDSgQ0w4EU/+oWlSvhDk7swlpkE2BtFyS5vgh8uNZMpIftl/88Kv47jUUCxgh6ueL7
WyX5uOEz/qAG0pjZfqzSs5UQayNIT3QHaGnvpy22b8kreX1x1IY0e54vqOI4lIxQ6Jj/+0f8Rw2t
aYd8GB62chzhiYuqvFHSmKPKT3N2KLmqSS4nyj8gOPCKsYiI+axGMfjkLQNSdRy9Y0mLtg0dut77
ImZFgESsdxSUbZJQD/4X0ApZOLEMCsnRNoLH02eTiZZBr4FbYxgPmqAIYGVL5yEXidsE4sdgr8Ma
6/1UN4aoh3OcGdZ7lqjXUj3V5gyvqcauPO8dAWFz0wqbdMa5EtRtLIX1gWhbECN+ZmcoC+JCRhtC
HO5tB85c5GChh7zde4UifaYY43gkbo/tvL75Uwva/XXzHLQxB7Ttk+QF6G1i8yLZ0SGgyjc+naOe
i36fKsSCfwwXankjCC7TF8dqRODmdvOYqAfOtBKRkMtVVNHdgCwaP3cha7Qf+WFfprGPAx93a5+p
hzKcUuEXheq56pAR2L/RaXmHGXAOe74VhqNtu83CHAj/DR0azCFMUr71nnYU41wpD7x6Ahcq73J0
/XCHR4+epejYDwir4hDV0GWmGIkkOTJXpTGayUpXxVeBRAKmuwIDgnBJZdHZf1YW7Q49SjRjVGFC
p+o+U+yvKzcQy31yX1Ux4w4RHPLa+ENRGuJqTW2eE7u1xvDznzWf7+xT7ps8zYS3kg26JDrxSqL4
Y/Fthc5i4ZDzXZeELJBdyO1tSCGV5cCZFSsH6d9PFlAW2TFNJGxF8MxZSIQIHsOjybIXN6ZglljC
4QlhLJVJMYaMOOG4dsoqFF3r8RGq4H3nl/RHWTbEj4GlzIC93oDoXQB08Jf4QpaSWIpCS8SrEd+t
I4jg5BVCInMFcjHQ75tIwYpyDzp4EObynpg00e6T2XtEN9Nwv2GFgR2oUdIVtzywxvpBO6TrjJBL
ceEQ+VqIdgHvfTevg0K/iX2/8Di+E7K39X5vLlOAB6NZVC71iQw0qv6qA3poUgqrITLtPXN4R1or
4mN+RDF1w9niq4WUpJPFoJQKx893smp4qU/2IB80W7Wl4uvvN1POCXLeopc8DHX96WqzXSmOx9AU
PkjcWbtld2uwYzVmb37mr8x++opVGHWb3MKoKc4MUsYeFD/I9Y5REHiTYU0AGoWlYFl0D5R1Mdjg
EVXRzkx2dIEYULYe99viWynLfnDZYr6uNULC+TnXl1Afg807AJuWCOonpLOw6NY3CrBq7vLKkMzt
ZlqV1twFA0E8UC/WSxFLf0BBkNr+pfwOrK9JhuRPlFYdbJsAqDvvpTcrQmBUyKcwqIkheD2CFOxK
XbwXOVKCeevvHmgiXwgmy/MH01n4Ditess0vYUFB4NjeDVkcXk0g890l+efmLN08S6ZAU9zMbclm
HGFRLd+qSU95OhnAIRaZ5ABk1yF1lRIQ7l2obwQyC5qWg7RP8ei8Q9RqsNDH5j2lzdEnWZZkNPXC
g9dTwLdMUJvYIfvVxjLUoY8HYoMldbgGHLJ+9bY4Q4FQSmLvPUovgB/46Z7+hOO1wasJMCk4C0KZ
BYegqcIViJaj/PIhY34SDcD8cBE9F80x+ta6DZcF76IRL1dmG9ESr+OOEXZWsEu56pDS7Q9hVgEx
DmGCoLM8ecqCY7oGdXAWUtZiKVJkq66burz3HYNDjF2oMcZ5akHN8z86ck9+1udIuSj2TLN9QoDQ
5LcIgIuaheijZCMihPx49Jia8bbDqaA8s8wZwYp3ElYEgOgBO0F9YOsk/qeWxsAw5erGCMlMy5Hf
98grjD9pTm7erbbvcFqrnBFuJxaFzvvlLn5QiRdzeZ3C2XJtBaBlU+L7ne7g4ZDvMNO7dFnNmpOL
SuTheS7/jP9cahKQbZ4ZanT/Q+P2eEfnuvarjJXSiITZxZfLPXDTSBbXHlDEU+FnDh06Lq6wIhi5
mHeLqLrWbipovNAeSQtTzJ45cEr3p33Jlp3IDZlrSj9SaivMujo9t3FQ55pEEiutm7qrvbkdqx85
GJe12bfO35F6Q+yDWzsTtC6qglBtSKp95tjjzlhpsFhvIdeXfUJmjB7NN6y3EB8qZEsw12dpOw8Q
mzQkZypWCa58/EWdi+kx9TKmC10w57RH2FJriw5YopqSBjfDPqdZNfzI9ek9NkDoiuvqF+fqXj4W
TAQjqnb6PBJDdBKM4JO6u/0zGKT4wvcW5i/BcIdah79KeAfy/n2ioXLHJtEA+ZcCTBZTj0AYz0yP
4va3P/6hvWxAXehg5IFMI7+S5T6XiWT8S95kVXiq5SIBBJh5nNbxxrn3rmDhojVbO0EVbB7lU347
7Y1ux7vPEY8MazTxmMiCduQeeK3aw4D3NKJ/XB5HZ1bZs5UylyNEa+80HL/UDuIHW79vxVI7a5Jw
H/Jd7+9YuppzbyFEVou+2Z6Fso8mf+J0tPkWcP9rTf1q+IUeLYOEVqsxKCKwPmXxVW6XZbXmc2s0
2ZB4xFg1d1/2izu3n3rKJIgVcnnX/nlhP+LQxsUL7uF6V3zqGOi41uCpgbQXc6FyA6s0VRg6Mozj
r8ZVkXU7GEcW4nZMvNA94DJe1anuiGGQBh/+S7jnCT6J9/3P3jlj9ImS2d23pR8vI14q+WVH+hS8
2iqM6sE28k84D5IR9RdcUgTMi03w6fVUUVWHdCnkHr/aCW1s/sYY4KZ8d2amHo9PIGm7cfUIDlPJ
7sg4MDi2Yfzplq1dQQEsipnpgNS8N2C7dCQm/5qbpB9Usujjwz5/WFrICiDM9qF/GM8wupBs7CXF
vCgtAC/VNQJd6hFYz0G6B09STlnmEnWW0D1g5f17O+jNUSMz7qwDJLNZmvfXgBuyoSUrvaxBaQOF
1Z+nY9wvl3OJ9yjLaz731spUb/TBQmdfiVLDxzrJTWqBpYsknAwRqVvLOR3IVCDMbWEB1mnqG1lq
YXrX6+KcaILSJUiGVlhk47hxbM0fcvakjjd0NFZsypeXXRoQ4wUyL4f2LR9Hdd+uzXVdAHgoA5dV
XPJKcHUkJAdHdbnPWnrLm16Tt2i71i3VCra9HDtatRSB+/IvwKp6g9gTsKjk/xmaLyNiHDbvhkZh
fc6ESKIYhr5CwYTtLfbXkJZDQQ8UsH+S/fsq2cOtko4SEelaZM7L2JwQiBVU+2dYFOcv7VUaUi4q
UlPJ4wNbkM2A0BVGFh4BfULZN2UxoHERIk1PTuTTlrm25rxRHftGsTsJby+UONqURsf08LyfS2rd
S2q10ZyrnCP26UvVG1g5FWzqZgM+620jwfaZfL2F5wOwQrk1UxUbwUoszjMl4ch0vZy/6K6ldbFO
O/Wmr9cUrlugXnuXvUzJ2mFrshkg03N1l8pENsYt8wyqvPBpmbeOfJ2YeKcnAb2QHu+Kosq0rH+w
TUmEUCzD1PDIUljOf3g2NoeDBMQpZvxC9DUeit/DS3Jnx0HSfB6Gdcpp8Bk/2+YL532pyHpxHd1E
s0bpjD+i7OtJaGGbdz4d73gBHDhpEv8jENrhv6HkuMVTSY01R5P7WYCxkcfNWKMeFl3ptN9hxQxV
DN4iZGkiL9n4JNLUTchgYYT76Pwe3qhZmf5w1CPQfwImjCmij8wxukXELGdijeBXfMUB0Q3F5RiA
/SoZni6+SR+4QVhIemRu7kVIZvcqZ/sGmWJYw9vpZ0JhFz6o5WiApQ2dz/V0V02nK/uUyfpRhyQ8
Oe784WhwKuA+sCAzPHQwaGlcG7M0+i7FjIde72+vmYEa18z6SzrMdhQmhFaJgts149Iy75q8xDVZ
JYj9ext250H52ELu1FvrKqBv+gdVSgrmsYgJQPQVtNANYxqR+i1e2zSkobELDZXtbmLiGuyurp+3
9QqhWA+m72tmUYWKIOL0oKGIxSi3Vrp9zoYujPRj1F9W6j+0uOu6s6icDS14G0s8x1Svcdp7kcLU
oYNYDlBZRaYANuq/bxE/JHnJTlLYhlFJ/4/82voQRgAuacyDkVqtevYG7FLOKKZ21gHQaqVs6gJr
lOS2/8TrJEaj3hqwataCt9kzqghWnY+Z3NtlXwWup3T2ptN72axRoYxhhhWBtOcnZ9TW0PD6edM+
dVuP1LPu9GG5fYavnXmn4q7qAHclj/s5AqZXB7Cn6BZT9Nt8mLBF2EmwuTzJF+LjqpGGLA4Sr6x5
8Y8vlVNBRR4GGtN8q18bQ53dbsZ02Rd7eM9g34l4ewqEtkYLYvYbE6BHkoQ8KRK0vNU8Aco+tKpk
2oLyp3GC7TktB+RZ58KBMFTVHN6etZl3nNb3ZBNmrW5t3erc4V4muGPtIuKy5orR5ulKF/x8xWts
b6Jhg6oxO9By97LfkCjtGU7WxDCeJCF9eC/vSQeG2Z0OcNAnuZ3Xh0MwIChwyezPHqj7K4814odH
2BMelLYel2I2I+CnXgsNr2Q46t2UmBIFBcsCMNFzX/PcMbnDG4+oUOD4RbvMwNeNCmrQfY9aD0Fy
jHshDaLdOYrKSvihJIPxnIUT4inzDgyS+/oIyi3Bi32yVwSzkVIt3sTq499eYaXSiuJfhI8gKElv
Q44BYJqaPBO6FIT0QD36hzkRAQKEJ4eCOCJTV0/mKgZmgPhKisKboQ/zzIUgIU1Y+3WncXwFUbDa
qO6+WOQSgyDcCgOJJ9r3BazAKP4IgZ74GErBRY7CijNtEiuSm9zBZNGijOos7jovMct7hGT/WUzv
m8d+Pw4V1twiaAQGjJ2yYap/LJxVB+EXJ8peAEfkTrI66IK/3x3V1BeTSuUXxS/9nvsiSB/p7+nA
4FmJ/geFlT2wu0xwxMCghIYXVrrwUHHyw2srrB98HIEMNoFWGg7fIxJGxWHIIVQjAsu+VfALvEcJ
mAYBfO9t45cPZmNMUOzmUHiiRfiV2fY5o4U1xL/cPayF8H1Fe7abq2OVsilJ7t0BIJwEFserptv5
tjLbfJvXUMvmMNfDt2H0QFyMuaDVcweHyfY14+rRWK/bX+F1uGkylLORv/k8Wjf3SAUvb5NV4Gkc
dwIEalCxKHhOuzZ0q1t/6itLKSN9mMaDQN33avqNg8VzhAiUMKLfQbPqxI0C6MGuw36hcZRnDIa8
RlXm9iRe63sWwZOx9ybEVO81PZ0rT7qtVzpnpT1iEvuhUWuUk4aXCO14KhUcKLYmtH+vTS03ez9d
xE9T/OkBVO6+2NP7gVkVZ4v6yEljQ0cc6nDygz0leHvJ5Vh/4/ETGxn07RVq2v/FXhwEHNPTGDES
S0Aj5JBYehfNl2+pcFc+WQsDIgxfe3f5BvM6MxUzfJaasMOfBpy4dCQ5FQvBFwmUL4sn8oPXAclQ
TVdgO8GpbDivRmrYg1Jgw2LWnsdq9+V0vrSUmOIos3VwqM8r32nYJnrPYSqPFPBznsqyw+2QfUY8
MHuSUFK2OVHwFla6SxwHBu0Z3wi1OS0m2YPEvHmZDs4nw7ngAKXc7gc7hrlzxULyVZ7DNEcsEFj2
2PyK33pjuMzjEq916d945xKhewDJuNPAAUVXywXfFcgeHAcED5sqALmZ9BNCDCzmU6jvvS+OewRe
PgG1sOajlz7R1hEpZIOtfNhiT0lPNV0ioPepp1M82MZ4dZnnlk8rsSU24htuG7A0HV3f/UzjW8Qe
SbOtFm87YdkXaGNS/YT//RGDHPDYvprXrYMgcwJ3vG2oxUjvQK6KYmWCRMPfkj+Dyr5WzLcCzBy+
IqS+drvyTRFXkWi1vSEK8JUo2qTgl0ckWAKHtg6dL0Yys+Et0DGjLbpCl2n98UEfaFSdL1f4H8k3
1+XmGS66KvcdNaJEtmLk1reuaX9AmbHYWVtKeGV5FLUHozajveFI3tsmk+kj8H0E6+/NbLtkCZ+Q
4fRPI7jMtajHQlPrX0hXdBuGftBoEkTbQ99rI9RU/qFh/9sqa4Za1ZA7v9PHwFwkMWhU9T+E9O6f
OfZfnuHQQOsxDX7/UHNHTYZbo2Qsrb8DL7iXM7zLBVn7RrqPl9MBUzjYKn7EMnzmFlWqgEngP6aQ
7+O5SgixNPbSMewogc/9bAVL6xBQFDZ2nP5B1qYNRzB3ZYalrz667dT8aqT35tEMU47h/QMKxC2d
uDIYHRXfj3Gbf75CaJlwwc/xTgCnZwL1YYOK2nWs16gi4YHzfjCyvhbcdVMFoED2zKBVstS4pDKG
YneXVHvaSyGwweecgB/ijY7zNCLT3ZJijwEKvdXuqdNUJnXn/7P/7pKqz1XDBGcCaPgNoD42GYqI
h9uZzWuvqiFuvDvsdcYfJyeTNBujGz0IVM18zsfAM9gypWl0pGCiqVHJShZqHP2Abxr+Xyvwe+e5
YlRNT+4t+ysbhJaa4kLV1UDJ60KQJf7NkDkr/5k7Gy+DsccYUGISbHM622TWYPr6dd3omQ1pIdgo
Ul+bTakBqPERjUqUSlylQF/2CnznFCvEX4looktOpGctMqN8OungCOqsKcmSqwXnO9xUiXIt8G+G
giAvvH2pRVKhunPsIzvu+69Y+XTF2dUoh2Sv7jqJDFm+V1kHn34INCoyD2QIZwiYfNu3txfAayvf
CPpkiVm0xylx91MMmCpyWzj20KlMdeuY5dYdSf/rE2An/CKJYwdG9umcB5Tz12k1wDktSuGl65BL
ymRdeUklyDRD9dPF5WF2iRoVS8L2jFfqQPkdX+cW2nDZ86zrSQOXN5qOYVGw4eDc2TzNGI08K/k4
A5O2l3OpyVjG7ooU3Plke52U1038/vmExzw3Q9GVjwd0gM+YBz9fO1hlXTbh6lsEsm5Rep4S8PDK
dCkXn22JN975/v2IsPRy7Q/Qs7iMNpP2nA+O7yyPg7tujVWRS+YzitSiXKhwaRdcbsszvKwpybpG
byqGxwnibfTmoR8/0/KffxE0DUFx9aZ1MBZogRVAmH0OS8vQSI2Hk8GMJUEuxxmzy3LbeQirOeM7
aUgxH52TbNWAOnyMdKKRFJnfYG60ouKJ4BP4oanrg/ONzmVSy2klAMo4ZXJLl9n0w0Hpo81OqdSy
gbc5j3JXzMtI8Z2DhuZVjOmMoQd19VOpqen0oglxC+YK2dLzuSsEyg/SEFf9iGa8pOmsTKkUlDrL
1ntwSp2URnJnMvKDRqEKZFztMmwIlORKvOisvAltVCCpgbEzSzCWfg+ryGM4YNGI9/VeYEtdT8Js
rZ/TPgcbdGIfWDH3ksdW+YzwavHpvgouPS6liuyufZlU/tY4JRtpQti6lE007MXaqpIKYw8d9h/d
MGgB2hUdPazLOEYDkP4yAPeYaQIC4VcIUmEIF9P9TvJMa02RKwRt4WGWzpNuHo6oMwC8+C03H3wT
cdwOETCWugPbzlaQj/Yhv1ki+KFiSiBQzyq1i+eI2cy17eYacuwYTR81P/1jCguOJXVR3dNVwQzh
/OVucpCnAZwJZx992yT9ZHfpyKd5x5l5KGrsKNg7QK9ugmeCyxnDwFZAsGA20pxkYg7tM7PUNnwX
2e5GbVkbI0rdAq5mUkQhDOyjoIg/YCQN9BUvYBdHaw3ERZBJBN1SovagfdzfyaPcvPkpi8X3XVXO
oltiacVcIAFUtIa7s8qh4D7uiFRM2S3Cw2XRrmm6yOi8z0ClCNKjtAbOj1843EVwUMBRgHkDZADn
9h2VNUdib8whv0B6iXL3qPXZH4aW8b/0AxkQZ26P6fOtChxekFXTiDcQyemDgkR7izrOL22crbtl
iPTTZ1fKRh1/WW9T3lzB63Vh97LAt1CsgUmCU19agm3rRBQiOuwJlIYnWFeDmq1jDPDLmcPW5rSu
UUNq/gefFA3LII+s6nmjyrWtP40K+RbT6FgAa4HaYos2Ts9G2irNbpMOCBTs18vFuZqt5kZLMesF
Rete5oTwlSiXi8WPGqToxzune/LpuhUXrd8xGddnjbB3EEKD/XWbbojMqV5WwGgWYL6znKitib+2
EObEqNZMECmL2v0ZndXCxfdQ9Yj37cB2L3Tx+MyGoKw0/WXIOwYgvR/QiH/VcF1E37BshbPrkzV2
qMqAxHxMMt+CXp1QopnvdSj+kVrFl8jx9L8HA68lii3Ld52SaNQm5Wag3ooeikn/UydjFrzYonXQ
ZRRoXrg263fYvV76NVmSkHrt9mJAG9wUd6oF0d2x2ibsySDdtFIMvnTuptyfPjoIgYXgOcwcYkN9
8RJ84Wa4L5zkjvsOPJJlwfxR24J0OU1iijtjnIDa71NhhcDjH4YVljWkyfjSSXSR8b4V56V1/tMg
5WLbGkPy4HSZRBQZkJqB8szxPH3iHYAl1jOn5BxKUEPj56PCz9VuUQWZ7ZIlNZEoOm1Jb7hmuM12
uLMH8gJW6f4UDRQ6yEUoLRI322L6c29I9Oc076dAGaD0tPQfkbVrjHdSPoPuancxozETMvy0TWsX
U8C2F06aM+PnLbMe9Nh4P4aIrBnCIV0cg3AhiLUNqDSfYkMcYTyPO9sgKN2lLgDyeNj1ZgGUcJvd
viLNlS6f/m2vDAexSvsZYS4KbJWLmwvJi0O3ajIzAT2IxqfI9IunCINBPp5PwcAkUqZhKRrCpMQD
UdiHIBvuvH+dxfxacFcrJygVrzMyLU/uLY0012MzDB2Wz5bFp63Vl37/2N2j8/NJcgGvhzUkYITQ
dcJafRImQorhGtf294il+D3LwLrKJcUwbTxNMWylsLtB3oBdvT6OZf76uVV2+vbdBdmErBInOe2a
M3/Kd9/F7063z7arWR2j81gUTOSdL0aXtDb7EtmHZ2j1fSpWlh5tAfbXzGwxMXuDi8nSU1Hz5eAB
TAxYAdxnL+6bd/wk1PcTSKNHqQKQ3SCh1pyEpuMWGEEBoCnrdfGafi2jOaoQ6XR71niKNWUJvHL+
MtDSFAqCrOxKWNnw2DQf22bNkn3tweu6oaAspAbJpXJviIynFU4YUi6c7K9HN0hATM4CjmQRR8lN
if9XQUExe9G97Gic/pqmnILvzriziEf0toJY2Ic6y14WkvPZDsmBQj4KuvJPyWDVrdyO359iS3Ab
fMNNmdytzyZ7FP4rR1VRF98A3ynSIlyB39rGnhzxgDywAOhitp2s7QlPfpepq6D7lRYe9VHio74R
VwVoqDatYDxegdqk/pdAsa2prrVEaJxVqVfg9wG7FUQ8VPpKfBPkK4wyA6tZYId2UKQ7mVO8KzQt
vVS4kiM8jUJde3ijNGDgWJDYI00i7mOErT4A9MZFXwkKkuk1POs5NLgD+o33q3DneunxVJFjmDcN
7J3DMFcqryMHLLAQJ215vreCBcvc6+rGqryHBJnCPny9ti2ldyJ1A5ZvOOiL5tL/MGwi419753Jy
tpY1LoPqT2mG9SPdyG0a/jCk7iAbVd4LaU8G5s8p4s4Gej22+swLQDOaEWyC7ie//6rG2huwZ2D8
k3V2wczlhR6R+UI3cOds19OlRYehn6skMqG5g8aEeJX4DcAttbPvaqGDn7JKpfGlkurh/1f96IDV
ej+/+o8uqmJ5MZDMumNtzUtlh4boPLY7jlVFDyOoWEECullrpB52pnxfBKew1Ve1wQuFZEPaDCRp
07exo+YVhCNp85mc1BCsI0zxML2XV6H1h6cdr9BahF57jfQvAVUvqaqXIHiEjbHZHUty6PCK4gQI
rClhUx9kpLxLOktSXlh8y2S+K47Dq9IQmi18J6eHJUQjPCfw1iyJapo2MpQ1Szt9ac4Iy31qq0ZS
Z+S8tXK1TcnVoeiwfTe5HLqRgIICw8bwhpj9r1yjhZXpTQj2RcdOabng3Ym64PqJdrs819Ag9LsD
m5wjUIWyy13P37FJFse5FMBhg5XPqYFbng9GjGava4CL1qiDsBIpvmUu3FjgHAn9GE5ZAs/wPoww
GTjgHbGvn8awxV0Mo1u5i7BLyX2OQUmDEcCiOxls3SU7iUd5wfAfJbqPw7HYdxn3noD/rLT+EW0V
lco9QT8oww4JBjkAE9QKUqLZ1/ME0Y9ELpNpNXtr5pBx7N5yuE3q5YE6mIeDJLTPID++zkQI6MuY
VlcAdFJJDB0VSWb3r6KuEiuSDcE2Iv7m8+AzxcUOWgT9oYX8dhGaEAqWwIWG0ut/BLknOnMMSJhz
riBzrIOwj3nLm4IjBvARzh0ImSMzcooP3agd72R9mJYo+fpXAhJKIUYCSMz80VeyzQr6GFk8Bg18
EuZbqFMEcQwL0lSwDwLNO1UwdzMjLKNrbDEC5tT9PR693vBUENL43jFeZGj59ztWuamBOmw/rzaN
ALmBFJIEnc77RGpsA+00PyvPPq5+GVuThsk+OJXmjbbLd7OhVoF0hw/jaFXrUgk6Q0m6Pvsc4w32
PLSdjZpqY6n8GZayI09CdxIfxCWchhOkZzrgb50M6owdQjuincqdPNrylaF/kNKsCEueSz9w54MN
bn4ZSQZVYsqHDWgoV/MqyhBzP6QoU2Uu8Q90YeGgszMtP2jXK/bFUX4YkUPCbfWTrSEubkGM7si4
9FyPB57YsZ5K8a9LA37WNsOw2rY3qljgyq+glFA99Bjbm0T0PkxGhvJa9XQlF4jrBtbGA1/2J2r7
d5fQ3VK4tmhuEA+GyINmCmKN2PM35KQT+otoSQjva+ti3wAtV/cL056Bmb40kBC0LT6uiNGcXl1x
x9dTps7OW4mZWSMZPnS9+SRNgN/insUW1oMZTgM840xHDDGa6WIignufp7easB+jJZ0MfwRM9hRa
Pcz24oUpG2WU8o5V7h5DEeb59mMeMtZdQTeMDpLlOL+AAVMAletjx+J13a8b2AJI274FmcF+Ys3O
uMS7qs1EwFdFmlz+/adUBt3rLf6Qe/ec2P6QMdJs1qudkB5HggOXe8ZNTbftgH5B6y242PpB7/Mx
heo4ygOQAUcJWb/NvoA0M8XnD1tNQdYDOgO7HtrbWqJ+v+cIacddozFQTAlRMffm6p5vl3JNbxF4
nJwv560WFllZvBZpKWfW9p6A3UfzNHxWmrfGVGFkhbJ2zZ5YW9f+MwsfSYG0jM6c2sNkc5xoH/b9
XzgFgFq+I4YrNUuL8Pv/tAi5UjR8woNEdcCYEfDdxWkCtcIClVZeCU+Iu4bC4jYiiFnyGU4YyCEj
DFL+pissX7tZ7HOS84uDKx8hJm0lEehjZT00EZhwn80n9sP0iy6acmO9iABropUNNkEdnPx9tM+h
iQ819T3s8M5Ls7aNwWEO5/uZgqVgw0voUApHVgMC1vMPNX52HMaOi8icBEsb7lciZlfhP5+C8n43
3KXTeEiOUgTWhOQtUf61xzYzDUO2+sK9djtINZ5x7WKiAxehahdhZYGszZ+hyU49FjepI08a7TKe
HPWfsQlROdGINzUMQ3F7c5iL96xYDTjzjOS5T2INDW8MddPkY5FaKjlwNViZDx8lT4ULU3lI6WRV
HrqwJ2vur3PrY85f1BYvLkDpnByetnEk6CdlxYJeu/4N/HM/eYag1axUM/sQTzSECdUayiwHYuzi
EeJYF6rQ51D+dTqzAz2oanEUQ5crfoyNXsYvNukDXEnCt5swnCOUn+pJsmaH9lVDk0DKmauAyo5x
ap+nr7lQcdeOGsZXQaNmWBwcxXvZZUlPhA0FNTDgJKOWiBVxZBHULiOn8koEMmpw+Ao9rFiJk54Z
QhTOZhk6PqkUvt/Jdhojj0+EkyYBycyc7suorsqoZfS7vEn6v/Pc4i/mTE+BL6jGnpHy9IzuF+s/
BkvFb2qs+iyLAIfKFJxiKw/I+dguPSHsLfwnZvLy/BONpvmP8nMURhR3go68nSwjWFqmPGY+Vp1O
SZ8sfsQp1Td26FIilcl4Fr0viIapTzQ/3CyODa6/Gtpc2+Ikzm5uXDrewHHaesvLxQ0uQHAi5pXz
EQQ9pijLvX92xF5kWcmEwXexmy/XVaI9xzEUA6HeBNLye+bSh1Z8KP9x95G3ATmjY37wt/r6BKMD
T//CRc0wG1lz6X4NvPaeRzOJegg8U9qKGUmPKI2uA9uSux4192KF4zRKvMlxPm1qXnL4ihBXK0bY
6vfWV5n0QQedxo1zlJ19Q2/GjWntGQHmRAUyhVaI7xs4t9smSsQ8/HAAYQwioTt9L60ZWMAq8/MQ
GapPl2+/iFByabtz8Z+FQn4U3vjQxbLY+ygCUowinvfMz9JrAC4LyKqTEYdD9P7DXXnHKhWGkLP/
QL/WdWebpE/JAv4Qr1GmPWcG/VWM3G+m1YjqE0mR5TkZ7H4CBTYAmu8zOYLqYMXZz0h5b7GS0+eb
AUEO4FUXSPp+dQJucMfNN8y2NqSeOtRYF2WDuZunkI/oeUs4CnuGN35JZBSmxEt7KOpYBJ0DO97p
Ec+t6xdVEv4lwCiLzrAx3bIz7+V/D3jRDFlKR6c0rQVsU93MPmZN7AGbbZM8kwlc3XhmxEH5so66
3qWtSlqkGgNJDmD/02gWY+m6RAb3FfEf1ayu7uewgTbw8xuyXGuL6EuuHyDMGOL/++emMU3EmtEQ
RT4LOUBMp47pF9OgsclZcniRKA9BvGFix2UoGQbQQTRdfO1SyGj9eeGAOVz4WLlLn/ZTEkAiICR8
xXCmZnFyx+3b+Zb/foH+HX6laP0BVHQG6XxZgKZlg7oNy4g1OIy/XxAs5ciBj7TcuQ1MbeCmCdTf
diWDSQnHVbd7ectVtKDZMNoLo0q7vPkHVwFs6EXUhUM396tAJT177OgMMJrXrQbzcPM6onkk6hSb
q+DfGeKAjj3/0qsnfU6gpJbl2Gp9lqKZ8VQpiB5mc6B7J/9GS9lKVovAYTMJ3VBRp98Jk7F3Ce5H
yOPfVnuhQOYLN9AU2zIqyovyOvKq40xy4UsLPbr6HpmjsWHtQVgUJwDQAtx+Z58sXqaLXLE0PMH+
mfOowXSdQmEGNbPEbtqYlD9Pnrown9L2KzEohtXUpV3xvME8A6uBo3xorTsqQAyasAUoUDiw8mXv
+z3ERedxO9dw0q4ZzHJ6JPophh+uBqBx/rpmi5euusVUlBhra6Diza2mAhTGFJaChhoa4vJ6b0A4
aB+/yRmnXWJbsR6K4QvvvfM7kv+XNTX5yX7LJ6QX9Vo9PV3v0ncDBTtqjiv/P7rMd4QHuuMhbe5i
f66L/tbwP2wFrylS9oQy800S2lEFyOeAGxksptolHuZZBJ4oYIUrcf33/r/KFvHwUV23sbZrRSiR
nxlQKuBqCn54FLFw7cuJ9cdZxEK11RNhBkGJSriFYKHOibASaAiHS1Ndq0E+OU+zQHR+22z+hkDF
i8GvSbgsZPNgujddjhuoBLgTq6T8hl0rBRgJk+sVGL4tdwyubszbyiGZxl1q36XewIj3B3r5r/Up
NjTO1xDwFtdZZWdZwFpcfvbk7KI7VLMGkFYuk2EkPBeHK5JuLRyWTYiP1U8ElVsXE4sdJB5eNajN
iPiMKpbgtk/OWPkRFcPoGWB8EvPUesYb3sscsuA+N030MAPY9y1gK+9arTIf9KKIACr61dCpTuGP
XxYlTJ3gH9euxacqRVax+f+/b/nPe6hbR0ck5be0VgWO/2q0iK/RDMcRqAYwbTt4AYNn9s624hj6
k+q/8S01cY45CNIuGQWMlew3vGod5H9chtWaCqbd4XnmHDuBHTzMf04B7GdjYRRPlwuUsiKXVYs/
KoYUFrS5fkeOWiLgLqUOi1TE6zqPHzrxoXFLWiBhiH2OI6iEC8ojafweRtRncS+lsVcDje4i4DQh
hVLhpfZ+rzV/VukrOJ/LqAqkDmA4BFKN3Ya0c2wXHI4Aq/AjR4b+HplTaZjOniyNqxqvl/YoAqvj
mEUtQ/9I5gcvfEvCGX8s1aH8W4WNHRtEK6P0RIZCQkc5y5XavLG4ya6yUI6cmFNzJ2pVxIxtmnFe
WBuVGyC3x1Y8EGYwUKCjs45nGQZZ8Ij/bu25GEG4tMC4rme9PZ1IpqX3s4mc4nKeyfHIJhnikbmk
vjEzGD+1YEFYHGQDPHpPLaybI+6sYLHhApxA26At9SuJNpjgWv6sxP7jL6qmJwc5uZ14KGoilIE/
R6p2g0Hu+glmgO+g48VGA8ktq+Ote+FyAGj+231u68zC6jE14M+QNVAq2F4HPAW61p0L3wvK3PuD
5VISTvs70fogHCBQX0JMu94yJ2+oyRRGbT7hNRhxcaRrQwtCluzkXh5dl1aJOVUE/iiEpNuNROx0
096LeivhMi0fh6zXGl+OgyK6xq61sppOLQaFp+nHbNDnKJILqrGVibkKnlPD4drvt76YM2wrsUKr
mv0SWj3vx2JxmAjgFJxjedg+BhGQ8dVmbNV6FMcxSJMNsFTLhh5l8zO+B30Ah/K/DOPkUl6mUGf8
Ld+L9sV4uWp9v/FXOK+2iEXPQ3keR6V10Fvyw7TpJJv8JPR4eCSNwAd3hJloeea5edrsOaQijUPa
wIc+vpADWkxgnU42LVuGKjAAu73aSQKXlPwTXbnY2poedR+++b2WMXl10kLtscIPOj8UjlLrSv3Q
BqIy7fKTo9z+bl5Weh4T7CGHLtZl8jD1kn4M2GTNflfVU04EUXfC2OGGNwfnJ5wnAuKQ9FsTxXA6
4tVyjqHeOqglLmSa/8umn8tFHmWrkMGh8Qy2V2+MHsX7p5JtXEv7VD1U+dfUvngdjF9t2RyQrEM0
8ZFTq7adDdzIGfVsxkDM5Sut/kNvftQLSFY6dWcOXF8AWSygPXv0VdXZcHIhESOv1HZUQQF8a0e4
Gf86MX+gGEx17gg2vJfcqOOsJCzBATk3iAgkbQjSrlPipnlGUJw+lIwPY/4O1UaGpwb0E67pF5q2
NUCCs31yaESgXhXXvWlDqltAwCb0snMR1QmjbhMD6INz1A1dYfU3wbV2hA3u+8ygibQw19XOsxjB
6BcbVF/+7o3FI4l1h6by1qgBIYVX4hyz/CrZcu57TI4vMuqQuc07PIuP9d6ca0FXo/eF+5CpoHje
jcYPfzOOdl70hpuCnn5roDdE0V40cA/nfbS7hSuMqeMpGC1y/tCmZFQb10f3iocLzx+KHE3IDgKz
f83Nn9XdtTxG0brNW91P7Ihuoz+iRNMT4YSdnDJtiOsnzCNlD4LGnL69WcyjhLsH10Zs9N5Qlk7h
ZWxOSSKIUjizO0Z7iCE08wKt+YIDpRRQydHuRl3yIxRD/ssAhlHpK+F4+bnOQQ5bw7gaTbbsT7Hv
TR/Ylzun1X/ongX1smF8nkH+y8/ksFAWGFMMQ1B30Zc28udd0jlREupPeB3ooJBtM608cZR/gHPX
pyX1kY8Q37IpNe/zeysn87RA1XetSEVwzfQ86w0P3GNu21VUMpuUHHAcyqv+g+z00yqYxayqfykT
WBQcDyaL/7EFYQ+SWxAlf6dza1jUUYQjgCnoUXfjUxzIuoDFMiPXA8ROD6bT0mgdkZsvm1x0XlJN
Rl+VO1MCMTXvJtpU28D+BeuhAiHIQTNTWPubAsvWih0rZZqfB2sJomP39n7lNjdVknPBGPYW8viV
PiAsDKZm/EY+cx8ZBH4uAHlxAZzt1mtIgZtcHH8KegZQLLmHopLfrmAtAnUa4JXBKVh5IpLI+YZt
jzM2oN2OTIlD3xToq8rayn3G2bxv3h3OLnoaCIvY8DV/43vCI2R3I2OxBSjc0flnAStJLpcuK744
yF2nTmSxiw0PLDmq0TIptQPsD61TBKtAlBxe9p79yDka8Z/u1UL1cGiOTWoto9Em9umgAVB2WMOT
AGr7tbzqTPiVvazpc9e6L8k5O0KSP4day7orhhYeksFGHaEyUTm/oW0mxyuzQUsih1WonLGPeh/q
Hj5kSJx2ly2axyH3YI/79rXlIsH0gLSTl5hzbRJzb3kds2/AjtiYKmUjQ5Jl4vwnE6rUaLugSUFJ
ORnh957mey9nlRZFIgLduM7gvi3g8TYGuD7C/iu82juqS8M+D3EL/PxFIPb9qGF3hXi1rsHmVq+2
OF6Hxtok4DGzlOhP+cwkgJjvYbgmASzXUFnTh4bq2UJsYtJPENNsLlIhSczVDHekK0ROZOEyjDAV
o0NTHtlHx3T/ojQn32/iVkdIR9YvSj/9Hp6l4xPUtDDKyd8vPMc1vbYIGuMVm61sNIO16+o44e3z
KRP/vFgP1LMWtddO4A07pjHYZKf2FbWXr0qBMtafFkXOoIDRUqTNFWvjYGGcSPKkSkFkFOPFexmq
GY4zij198mTVYoav8IRPF32PFjqP00uyBkmFRfIT0wJZhfANj272+OglTEv3Pn/0CLvkR+a4i6Kl
FLk1yYFSPB8soLaZgLPN4Dly5wKMENq0Brti9uSYqQtH58dL87Gay9TCmIrNgv0CtRmA7jeVslUr
kIXRZaL3D7kt+sOYk6vLRqzBqBezQawnP8nE8hgnHCdTgXdWAwKsfTYP5ykuU6v+LlzbcwOOD0AF
m0gpdC8+zlZ42Iiq3I1O1QxvdecdOnfnTW+FveqBew/55TE9/yZV6Y3V1GMXK8bm1oTOl1bFzi7E
3uPbTs/hDsaVD3H0IfzT0Er+eVOPZWl36eYbzoXwNxcjijll0OsWB0UaH9kw9K5Lkxs7wk0o8c2Z
haqIDAXujOZEphxJrnAAkaUKOi6zE+rhyiVZssBMQYpAUFtBLhfuEiEmUlYeMePcjf4N/5LeZgoY
t77qR4YAHkfmpJFTEKKZh59aT27JvI6LiCd4kbTR7MeHD4yW0wmLOn6+Xb/6reRUqSijtCUl2wVc
lk1CyZNyb4PD1CjbPUqSuGjQaUfh1OgnYMVlHyMAlNnVqhdEdilAuk604nQ9piepLsKnUaqR7pr1
kSNDwBFnUIK9YTZgczRNAp7C1fUQArWzREjkdnCKuvCmV8FTevklisFgT3GDzR42VWQSrKdY6P72
Fjsjz0l8iRCZ3EBJz5C83e1aZonRj7RcjPXc9Uq85ExGjoVty+fmQ8+uw1z10eiHyLGIBQiGXJMP
/HgXV9Mxu8lIFFcC1L5ZpW/Ut/l1xydRZfKBPYT+d0JRqIBPGDAhuRcO6qIT5cZiZCWuwx+DwObm
kyvVwzcga8pbQa9LTgwZvIlfDEA4rB9BFrEpue1RguVomNaG58vK/XEFrOu/t/1L/Y7i/zMN/cvs
2pKaw8Avlxmi6290xzq5ejdLmvBwzqHlRmViix9NKkxMwI126VNoiuwO/3vot58R90+i8iD8bvIE
Yn72fSlx8qPRG6SOyvBFTJ/GeVKtV/6Qzasu/OniR5P5+W+abosBPNeYLJ523dHhlZN7SGG1rVne
FXxKV4BJ8iIMmW6+gHbgRKCulB4kco70lvyGjZrqP2DIAope93sPZPG1Ef8idpJ8XEyVOhnx2efO
M1fIaHSv1YA4RCIkkmE0vaRird/rzOMu8HFcF2YSoCdurS+9nWVC8/WW/onbtV2187w1FsKpIEh6
XIt/M6Wy7m4Iw/82MP7jUEF86WbApbgzxCVM7rXLuvxdhuoTqsmMG0LMMbO0PMSn3nLPb+tB8sTY
vOCRgltSl1ftOPnB3g3fvJAGtwi7PrPRle+T3d86bQkrbjKWDVMqqcgQVp8MD9bflCvLKeWQwDCl
VLR4McdwKyqoGjXIIQztwWJBHpG4Pmnh8aopFWyjzwed2LGlMJ7UYrmr7MCdarv6De6vYQoymKCy
EUAHJK24ILzbCe/SyuanVbaN6Wj0fkNObxqA+7VeNFuWMvEF5a+EvKzZ5du+Ik6dPfBFpbRBHHix
uKpKnHlxMjFTBnndDlDU1ZBORmurcU5LLuuiJVuz3qGrZN6rE8zsFgdJNxZazqk8TB/+m2fuJ4cj
TNBxfjRBmn28X8NkjsuPpv8C5LYF1w/HhWVqez5zeeBA6IQuCa3qEeTAEx1SScRnN0uuSd04CLM7
ZNcD7yKMS/rDKqTmHnnm4cktVmuWxVhOZ3J/uOu7lghxaT91wkPO8sGpbXTLJGxBF1HWtM5dnJuS
Zaxg+Yb5OuJE/61EdWST4JB66DxuBnxiNp5su9yPVgzp+eyxkJ5nkUnFdtfkUrStoKB6IP11zEv7
R0MDgcmogUkH2C89KgZHXnpg4WK43vLZWcp4BYqnsi+Eyc5a/R/GH7SZSPJ+7d8jmOYbeTdGCoqk
LGEMEdz3xGqXZ6IXAO24UthbZuqjXAsj7NjJwrIAXJLkzn5JfQbseEIWJ+HtjSPNC0ZfV6bVFcgq
hLavtamCx7TAZ/aemiVauq+5f840OHU+WYjKgLyToerKX9NlNUZVPLhMheowgSvqxXEZ3Pw/xq7+
P51cwfAeWS5hzh+uRlGkAtQFS/wUvJ5cT/kEnK4whGnziqFfnj535tVvl1AloEQj8wa6ObqVt058
G2n1QEEkY9aDxr9Ojv8GBxWjEgugvSteDtigOSKUDs1PvJjvsUCWkFrK8MhmMMKHB+oGV535vorh
SEbonwyGkKwFxYD8wTlUzPLGRwb00nQhLLenNt2cF8fSJ537EKc4EASWLBvogEn+oycKJ+aO3Y9E
DsGTLnozEpWw0QXl1g/cdqRvkNg1twHqRilxlsv0A/P/fl5u3DEH6FI62owi7z0YsPgf/M8YmmSD
SLhIuXJGsG+q5DlOMLj48DDkoCFa8AxCksgM4UmoVkPP6zGKk4fRLTv2vUJr790z2qlMscgPCX8v
hkSAgid5uiZYspn4ONAFAG4TpY6QtoPahOx72BJXajb1/8AJpfESHPnvjQpYz+MHm0DZCavSlm22
O3NbThf5q3hmKygADMWkZtJCwKK0ysSpzXxAyA5KcSWfyb2bWYya37xpHDExqitEoIQczScfd1R6
2U0Vngy3KI0sTrOTvuI8Dh79UpUm/Wfo0aLGOOhhImRp/norGqAv4xOpFk6QRGlXrJ07N5PGsJk1
9lKiKtSIRU94NhpB8pTnatpFRvChb5BUvZ3y802GX0a7qgzW3/Pph9YJqJn9xjxYvpUmJTxzSdhG
sBOawyr9L1S7Sr4Zqq1Cu93EhTNFJ2atbsOznU6xnGWLKJGeMydifQkocGVH8dQw3K2OdSxdQCOa
+oY+IF6ZAG5Du2gD+3b4oVoTPGfcNco1YhqfhVYO+bZFMXFoG9ngwjVc7e7k9/4gMUjV+NqX02Pk
hkV4J64k+3dJZfXBGsvjBZaf3xqnK4STm+y1UgFAXPGgnblvLTMVoU5t9l02WRrfCHRYeTzTiKPA
iJ1rV+J7R1XI/sxDHvJ4A2sYD9RjY61sX5HX+nkq4v6DgSnuyz97AxvJAPxO1l7/hYYs6UMiM1l9
IKa9vjcqjSnYmgtOXmPICx4Uby9ZTWKLw0spXfiRFKL706BOYkllB6Y/GCdz5Jtgp1yIYl4t8m+6
YV/LTrlHHpju1IVbFjviLi5xEh7HW7oeKS2AuuofsNL9TsCwogpE0B8U0ZHFF+HJbUWf6nJ/gQoz
WkuRoATaYSzSzC9XokXmoJSx+qAxgkY44djAtubYKKtSyOVk3SF6z0Tm4/Ke3/JDOI0lz90a/jNi
sVaj7C/LbJPKj0wMctseP3rCku5VjpDL8iZxcuA8t6R+4Dvw9k0MniXZf2TqeaPGTquMD24OoqD8
9oQZlB2BO1WiDPtNyh1HlMHuSKI11/X4WvlqN4/4wOg/+OcJtEz20q1jrxjwSwvdmg6J6doEvLWC
8P9xYvfcY3/GDvUQgiCQ3iQloqqQKkZfGphIlBGEo4YwdJQhRJWynV4LSD9FTw41kZk7/YxgAMo7
DP/HvrPcKSCmNNlqGupAYdgsQ/t4RHEP1c4CQ+JluEd1SZccWluyBI3LTAUnKCgWWVAouteWCDJP
65aaonKQt4cZWmsL0gACYr1l1MzMZGOzAoFPkwqvvJxILoYuFj/3eHsK3ll70dmWpYuvwR24xlO0
kQ21q53LQ9cWqnUFUWIHPsY/W8l324JByPYjIUqoYHR/a3gvCeXUF+XFDAJhGwwauG2+4oW8FNZy
I+/PWZ9cZ/xS78ubAnyY5j2LnccBT4q+/gpFU3v2ZzaVWmEHSeC/ye3ECSoJILHfp3AA6H6aHwzo
gp29Ly69UdjJsAG+Tm8zl6sgqeNiw+XVNLwha5sfd8fXlp815UnjI+S4X9dpeEaikUc3qLsfeO/v
lHTVCkjHA0vNGX6fk9HxbSMSmTiJVuumPmjQkPLkIXy0SN9cfSPKhcAG7GwOGw7JoCOUe1LvuaIt
Obu7dm0ueYBZVuUvTqKqOlzfv6r083IYaK/J1k4qufXJr3Oo5Q6OA/iEAa49feroOfJKJ+YIBTPt
FdBt5e+vGjaH/pfaHc6lB7b3YjczcxpQYdCeE+/gj+jV8dtj4mcjGI2N/w3ONVWDgfvR+34mft19
Wgf82lxSBFLp7yPfTrEPwZ2tOCHJk0+lVEvYdN0yT777GnRxnUv8IiGVPZn2XnINo9Ae+WxqxARB
3NKArq0vmOrx/JHj0lcLHNFl66sraUdAIZAYXwV0pUSgbfpS1YVSL9SNmQqWEcoUy44ryJ6n9Uok
iZM3fwIn/xokMroWpxsHrK4SZz657AsNlJFGYQgJ5zczHJWIzVv4hy3ljavHFeKjB89Mt+KNOFWQ
ezTNieow7U+uDwr6wZQpH6CE/ctjrTaQwTSwpSaT1mXFSCNhElbariKMsacHYzY062sFleCT6x/r
9skwcs69QwMeSx5QHjNCnLDntRjgwo+sgVUoe6hds4KatP4HTfpuCFoNsYjIc8KNeHMJHuDSn9n5
bgBr/8FonU8OxQH/RyaG+L2fzTzcXm68fwPaJYFtlkJvwJm7q1UKaB9/z830rOiMoz0lT36pkUi1
TMKaXZUgs185aKVjF1OqTNyDeWOwx9qXfbEKPSqfmFdKLVbPXA22G/1ic8uBgYXXNxKOFH9wCa1v
XjRi83Cp7qY349126cEIfDMBJQWqeLctrZmoEDGSsVtpcF6yBX1oXFwl5V5YtL/T8s5lMXMmp2P1
XkZTX8k0+GJ0cQdUgFl6L/m5Q4vkXBtsln+bqwmswJ5RlW0iVTeRLKVgd6kX3Ckq25uKTOmu4H2Q
0KPfxNNchtaUF0vmD0H60UXoq1zLqNFmlh9k178NMSkuz9PcLYE8U9uKWgCoWPa+Eums+ctoGJrY
pgyCLBQSewlrhH1fawPdxK2BjfpwVMi/rWPWtDx92LgowSrV7oI+uQX56AlGPThItEw2lECb6F0v
c6/95c35iTW12eslWO2V7dGiCQhSoloMoXtswyXAUclGScUo0y6jzy4m+g9ynmLl1QDH9DTeTMud
9+kdvOLS7kEyb9TLn5EJBEEsAF+xZy8DcTWurxT1IIJfvrIpCgGXLgOF7/CbYlZou83qs/4+dmf9
V3sNl8VXaSB3+lemytOdQj4Q9XSBTbp+3O0BavmXxinjDQoOfEcv6nvBx4pAE8xwb/E484vezL+7
UJgG01GkkE+HNO+x6SWZtajuIJ6JLk1aHN2zmmstkLR6N+1JxqDyDPmD12sFX726XuwUdRhb+9Td
tuEebaJEoF5DEDG6dHnSaeHsia7UxoIbsMmjNsWwsCHWNI5KbKu1f9ROlWBcfXWGgCVSIM2yrXzU
yGQOjLsB1UCENHkxnu0xaCjC8tcqgXlNwpAlYXRjBXV5o72KZWKm1HkQw+UUCNWnsX2lrMLECo3z
XmbCLtLkTS0tAmqc2kXZ57qKjhY7zYV9QO+o698czi6am2mjf35v6AaXurDUGORmbzasSfp6hp80
PyUIOz6clFqMftj2wX66VaLwKT222971pxtowPme69ojHQfPn8u0jdMNWs34L+pQIdShA+QPLMHn
1SjkFfc/DBOjTzO8vAgQSGAbyIQO/AfxjQIYWtJoaSIB+Hg0012HTdHD6i1xWzrUj4rHyC+A5GA8
jWnUOmput5jjIhMfzaKZ1nS5lujFwd/N1FqlLrcQCD5i1tp9eF3G+JBDfRCrSI0mIFlT/kccph6J
sB4vfO+UoqMR6PgOH/B9rJMSTLPc8eUB8Y6kn21fYLJUHjoEDBuXEFwTHP5Sm2hKYkjrpyT3NP7l
8IIjPuDk0MgVDuvI8BW/eivyXufQJfVLJL/B8yPRFNA3UAI18NEd3x5Qmq65f0SjjewnqsA9hW5H
cpVvfGC+Tx0bkCU3VIAWMZhSsuF+ROyHhy2vExq/iBEKoAV0ntRedNpV8GwTYCw546PxxW189HuG
TH3zyR4whVgZZEamIKtLTd/ulXNMn9jW026KmKSUVSf4AtWpCbydii21/tFsOXQYut8c1J2re6ca
J+jxtXOHrDgS4QVruFWbyjweKbLyTp1nHyaMp+voYXGQOu1sTF4bZSUFRmQHhCkzT6Rkjlf+3+lm
H2D2H3gBh6yeNBQGEzoFXSY/oY1sYb5sRP8SVO6sH2GY8eVy/HryR+l6oqh+Rs1syWWE+ou9mM3A
WkBcxyn89vokOCWfdQ8h9a9a+O/nlLBmaq3dmHTu0tQ7F5h27evtYSaEE4X02WQZID9SNvExinYi
+OzQtMtXYwAnrT+Pqb81qT6NYOd0E+S1084oy6nrB2c0wz8ZL1/SZvxcd4t7qMDOLwc1QzcWFykU
atVzn5aaro11hKuPm7ubHXC6xKmarIMA+9RhwT2zSFr+yXMsMD24lq7hb3PI0PqdkhzIbHjzRcis
XMmK4ovUcRDLxdrj0q5ml9Eqv4Yvf++ducIezo0JRG93sAR5/1Bux3+s0UzI88I0U1hUyGfwOYPn
lNlf2aS58aTk+wqkfIOBWTHEX5mN9ltUYlSGYKzQ7lnr3cxk1DlQhHJjKxz0XJsWnPLFC7SSmShp
sKC4JHrKMtEyjfzlWs8Va+Nm8PsRe8K0H0Hqyxm73OlaR3F/AKH1fs89zC2/mx1hb94CIjsTYwKA
nQRnk/wsBQ5q9TG2rJmQenJ3mEBB5ddQ2TeqKSN13+K/ODEtyfl2GtkPCRR6eJJ2zK0TSXIa7up/
bHo3bwcY+ikGlJOoImGK6YVL1uElMv87rwrzCIM+DJVsy18Qo/xXwqTl9Uj6Ss74m3Mmtv6VY3Cl
aHXad2A1UsqCXgxdrtcPhtd75/B7BBX1xIycWBeAhoKej98zRCL2fE/xpU0XHeKxJY8SRj+Yj3oD
FU4MzIV0FlejrR4h7Jdk0l1daxTc+j3N8/7bcr2lZRDd1rpc4hNkT7SJN/TIxuJB86ozlv9zNiVD
wlJX7vG5aMsFaf6eGqKh/zNdCRaiH1hAdxvIdC047475cIrbEGhuIIQBeGifbEyyBl2RuMZsLMit
x38VFYP6k+x8TQvWIY7z2/aBoEyBlntN/kYWGVjEe7PlRYHSDqJyLcAMV/RHEyVzccnWChiQBNFF
oo7SgYS6kn2NRs+qBozgUfUmyGSJZQPhF6SJfFbCetoY2R8AefXR+w5llcvmlRXLwahQfDxYG3z8
FDUXfQUcHdNXH1j/sDeXYYfLBQSvRjDBOKGwkkc9clWcOsYCGyavSrpXr6lyKArSmgnetrrzwvNn
3XKVAJ0TtRwJFNNJL3pz5nAjf2IVFYVCjDSkdbxssmdArhVUhYwrvCnerxYTje696/Hz6CqMTJUN
lXpMiz/nw+c8xDPpuH+jNf/Lo0CT/6Su/VRkz/MBXzNMSjQP887U14ISxmJto8aSQi1kPA7za6iS
Nm+1aGsL3w/sugEhV0FIv+S+VJj9uMhLWF4Gk0uH+nSaH1Ja8TsYklzTJDPNhAL2R959qSCCBuyB
cY0ImZWlxoCqr6BtqNBgqwdPi8wndBTtM2HTd9lFgA698BqFhYXQio8T2lERRmjw6kCunZmwqY1e
2Gt3GiNhGIFRl3YNmEq3Rkyyi3tSVM9hm8l9iq7ird1mhe+wLQ4nV706T4shIBTqTLyEAvg+nvmn
mUQEv9NFizeFmFoUi9hwiJLIBSWj8sBl2FWjkXqMOeliru7NXQxKFUJ4ISwf44f8uLzG4aHeHEm7
drgQqOd8C6YZuxreIxWLcK7awPsmfYPQhpTt7t+eKC37VyLlyy7vHZIVq34HVAXdGiUS7txgO/mR
PZuKuFcSyarH1SOo7INvH8/MPCtl15U2tp6m56QH2/DOk07YHSW2TUMGvuS42Moc2S75foQcTH06
fb/BIzizbPgu12i9ZA+6xYHceTnUMwCkCF86duUsyQmTwYbB0u25I0FAe0O9TVxQASv1t2+OQoZa
LUDvyGEqF2j2onQ4dTNIETCF6sToDJBK2SgRXXRvV3qV/PARwlaDPd5NYn5IN+CEp553I10BImst
fOVmzJhEtyuTwLOPxA6NoFUEtTcb6n4s12KIGKi+nm6wCUKMfxWuaGvg9raJQGHiTmN//Zro9uH8
6orAaBPx0krzudTgK4TZUgz+Z229hKJFyJXzZb0tWuCNkDMibFVdXB3xL7aHi2CbRxdI2Ljiiv7w
iIbhNK1HqbL//9Zo0Md6CycsvnuKloKZfIpY42oJGouDCzjN2h4pXbm8W14g/RSJgKwqOueVx1Wa
wI3VtVqLyxLfqvfK7L3eKsTxj3MxLeRPp4GPWyfqjVEMihkr1zaj1Jm+7zQIaEDApi3oKZl5htiq
XmIC7z3JediL7nhkPuG6I0sZDw9IJkX2dLewN2B99gH//rc6vTeOSL25b51MfnkBv2gqOU3D26bI
IjJIGD1ctraaHwV4JLjAVLLilON7KXX9dRWL3/6ArPXX6FbsYwayieqmwroUy5YbM2aah/jvxeDf
PBeMwWyv7LgrvsVghS6l1uQaNm3+yaqxJ+WJ1bcrnveMAFkntSYvOSc7eDAo4Lhlhj0oZzetw0iP
1g/oRoOwOL8S714w0ohGcd1taWraqNHF4wMxymVrQEYhEOVDZ+KtwTPcFqyOsGDTcEXm6Rp4ofVz
kcTmk5bSZo6teKyVjJRs6pDDqfbT32edXAaYFK8K3OCTSqkKcKcTfDfECuj1WI4Ci8ehg5+eRGMq
7YX1MHGeoeickBNjyrQIs5xLUebIpYbLUFwbmcLkxjtDjbjwavt1rFUiPCuTjxnsQ7tUPQr3kRbB
P3JsYGwHD9ZoAewoDgPqF7ljQzeGlKVpTdHnNV/sq/eDVWhBD+b3V6s1MZpWadZJBuWCHaKGzGDp
R5/CxWQL+2ExdiEkQOKJsp0tQqp81c/Eb9Y0Z/+M+zph9E2wjN9n4w57Rph374cglP/5LtZeIUSp
4d/WQZV2UrEKX+AwoCCvR0I6nXWXf4Q/YY8RgZFQU79fRmqlKPEHXQt/SFI7n50b9Ijw3t4Q+Mpa
hbdkDu7Vi+Cpw9IeifQrgIYXzV+5NaSR+MP7y+/sEjcakZTQd81GSRuPhNWIo2MLyEW5T2Q2pbZM
zlxAfn0NgZmvuyUHeXEc2W6qpXQLDGY6P5asrI66pWCwQV0vkGXkcZWV9nDb/uLf1sKQLn/8JS+9
0PQjsyPNz65nPITtJueOTU9pbrSiK4zToDMvLuS1IliAqlNMG3jcctcJl14U5XKPiKGhzosOwdLZ
S1P28T9PbfTgqrN5GgRspt17qcU6i4vinmcnX35FokQaihq/SJFzzhuyMXfW/mTzHKX/w7HM4s4O
oFwlhn5jnZnPGN+xRmeaUyF/Yh+Px92/fhwXf1BqJfV+aZy0sVx+3qDYvwlHaw0L+qrspjlJ0V8Y
afVeycdxG8ealHvHEyP2ltL7Y+xK5h8Rb+5zI2mazYs9vNmxv2qMAWJXrHxtRcrbpENSM0R67T6T
247dwH6Uj9+vFRsUvNKjrYtRWKSPa2SPjU3DIHwcYq4VDR281Z/z3OrZAHJkxP3gd5qjZ97PJN0X
Il+KRIsJ5KQtxx2d3ytxuw2tJEF4lJbMdtcwWVXV3I7ifF6hcPYUu5ftqFWxi/JM7EDS05W9VJkl
WAlK0hBlabRAlsP6zAYmvBNRRNB5Aq/IY7a/RCCkdOvF1llajnAJ8ln0wCXdF1b1efiQByjJ5+BP
R+I2onbjJmJnhv1oOt5ZxanDrePjrj9pEzzZ0Mz1/QiEpM7cI9dtMK/WTaI6q/1AKg3zfkq5kWRE
WRtVMR6Uy539aEKXaU5DRTaQpO8SkaQNOPjRQrYn4lA/mztha3Y6a7VMAfXBXx09FbZha8F2F6/p
Bq/QWcY94tqOpNCGPXei5GBjdJvDM/aOUhi211GaeQMJSfCn0teg17zrKkv+mSOUKTGBwiRMmHT2
TkyUh7145xgQBfv8dxFUdwjuIYJu6sVf4VWzm+6kh91UOVIFiKi1ExknpXeNV74HEmgekfRXV3WO
B1tXmIhZbVDND9qkJ20YHKPRHF4kwZONr9CNeg9h0pOCM+js67VLYEXfyfraSJNWkPNBhLvWCr6d
GrxCxeV0+jxjN8uJ4YmKH/POo5GwOY6ZrRikOPt8x/xUujuBzvpQ9w20uap8JyktKeQiV9JImaWs
3D/UDQEmW3MjqigK6mAcxkN+HLGO4dHG1wNSn/4SoF0KsOb/Wy5vcDFn2OdbgjglzigZYETZnNES
7Oj9errh3Itiaep1EczgifG5b4CavsA9paEjpBjYTc7jYuODA/nmls1XVo2qaYKzFhdgDXiYaO4Q
UdRFYL+YCPV6WP68fxXHZP/xpM7B+uxQMaGxq+0U63+A4VKCIaOGVvcqc5fhNfo12E4j8eptbQDt
Q3JoaBpsiKkYnXV0x8gFcNxLwfIyb9PjrTyx+9bXGiZoH8qqVMlu5QKQWZB1b5MT7POgLAjst2lK
61BVxDXcXFJf/FJle/ybd7Hbt0HSO4GlsBHXgkLEAoE6phaFeyG85isfwKv11iRgWvQ+CFtsxXPh
cQefDNwOCskD2XoYayTPVsGwywBW1fTXhlncFoTEuunSSIjb7Z0Es/BMaN+zPKxa7YV3CtftT5Xx
UQgCmqdWQf4wZgXafH21GolUoc0plRMk7sHAoPrYsAmAVRw1YAnDUsHa0CFM8S+qSSJqoPoZW/q2
5IBcZJTbu194ISaxbXPQtel1iLiuDoX/pDU8uPWBCmZOCPur8SbQEN3xn1ThCSxhgvT64ioBqkxE
2wKFLyC+Otym4HXwSAQQW0nB/zqdtIy8a+sJImibTKz+D/SOAFlYduZ79HNA8v65ftYehM5HJP3k
qkOjiS6vRNDMb1yjKvb5vNCO7YqsCORxWntIir49u50awyv0Tb8ypyuXTgy+sj9TehWdNxrRGm48
bKIT7U4fIgacBNM9rzIpre+Dvbt6QGeeft5ai2kcagW1qfvsxk4vQsA0s2mEozCwv7W2y/lwCFax
nPSRnkixR+vgSdGgEQE4NAMi/PAc0vHZWMg5+lBnaRkKsboz6Q1WtCarJVpTtLnamZxAY0Dx0JMm
YzBeKpncLXN+71jrg6C4zt340CoIRspUuDymyWbf089857NiSY5Jk98aWWUbGXHU06GSCdESahFc
zxZ3CcbSCWCIrxxoTVieVNvjiP09YF04zZoAB0tMk/LenDkwYbfdCzBZTa2PstvHrkAgpRyPrm+n
TNMFCvHOT0uiljUeJg/GXM8rO+mtcvUoZYA0GmTXiBO8GWR9HK6Po0Lyf5EZdFWo1qjtmsC7BrPH
/Zvw1mLxCnv5U5dXJAxsu5r203oJVzgL7UOxZlTqpJlyf3AnVx/Bj6UUJ4BrM8pg04qHbeG20xkw
HPTbqVCze1DcU3GFf/XD4wicqil6OpgV9U99JDdoR5cqJiNWRwqKIVYl9ixpdXbVckdPMSmIUQqy
05p7BLo6jaUTnOwCVTeHvnkRkvvPk+iU5oX2YXimulMs94VUermlUzoGzg+tdtkT2OOetvRVQQmq
kqxsBECF038whF4UdJCu/enoMaVr6rbDMG/LbX7PQvdQT9nUs+Jh/tfCF1hjS6O/Zi/G2t0ff9rH
kiBJ69Q3BDzqUPzPA2yoazYl+C0IPLz4vHOX3Oj7BiXwpi/ialcGv+qsTll57NWrzU88aNIvt7pz
hyu5r0sPtnkA8x8PoZTorIx2NQqR4MQc91zz/Qvc9XZouXK++eeGA0U67gcsLiPZjH8kib/OMoqZ
fiiRh32Ov+H+z89cKYpcxMOAOAcBHIQx2eZVdUtaONzYWPS5h/wycxDf2Yq1MvHTzG4qYThuLxat
ohxno/YICUHC8lRdVNMGrYvfhWtaN6368K/9Q1/suX0we7xIsYLhcZFGs6ebpAYUq983ulJBThRn
YIzMDeSHBLo1gnjuKIryiErQq9oNaO9T/s3tUZd1KP4lBoFM8fucpeOIQXMmubsXjYqSkQYY+AP3
A3f5J1+evfDQFnZgaqCIW/EW8ij2aihnbwGMUExizRyv0l2um9jKYBYO0aO7sAih/njAW/D4/BB6
stsS748kKdhuBw07W5iPuC0JuHfpcIoby9Z3/c22K1K2Etc2bT3d7oOvxsd2ec5+vkNTK+Sz//ps
fOe29h3jNT0B6qRe3Drc4WGNSv2LF+5eZqJjDrBeK5LlfL+Uwr5G/nx27Y1jlcA0Va31M91hYa5A
KQmpdauog3eMMbRtVU0eIFVWXw3hvnblbrqa5k5VqCF/kbdiyCxfGExqWJXY6KnCMh4rZyKiqYLS
ovyEpclywuDAukLvMY1ZqYe24Cz+DgKiy6T11N/2tn5snyV1ZjisbGwFl0wTugDmIYIiu583StRV
ASv255TXzKHeX9YSLQt5Hdef0J5zHEaxZcR3WfoMMGbQo4U0z/T775kzYjxy0lfsfE4Ke8WrAsoz
LzU3MIdGMkrOawviHKLd4AwT/5QtH7u4xfgbLDkz/5ochj1Otgc5TICbTre+DAbzJ/x2nDSS5ZN1
FrHzBx4xRUd9hw05TdGuHs+thGiH4qN8ti1/aTxdAnDQFfPRjMekPZ3yc+PBAPcoa39lfZ7BO4Es
AjiUkGJW3gfOZqibVv/yn9tT3k8kWpeRCBm4YVnoajnRGieMrR/RUd4LYYl2C2bX7xusKJVE0X90
n3FtgwMxt1F8THCiHJAXSjm7l+1PRjRB5ScjyimHGg+oR4aIi11zs7NpUDxJYCDZMqjgZ6/xbdau
W02oH6Men1btgrEowxGGkc35nwmCyNm91hT8yyRFhTb10mQlGBGr2BZB0tepg9Wf9e4RevJG6eks
/cwm3NMsOjZUSDyGD1+oiYmqfNBKZZsOMevCafWahdC3wzcj/sCnzgXQaZJ/iD+P3LDH4ozuL8my
3IwTIShz2gFNaP0dNw954fLTF3YKvOQy/TzdbkEpiTY1KNQJQ/l3rIc7/2hPbWXQvUgdmqo2VeY3
xaTMZtaBvr+rRM/BzqkUdYlNh4vnJ1UYx59FcHEEu+mf6R3NJmtXPLGa6Qw4wEm3Ce6Ybq5hLw9z
a4+06MY8jZAzQ0wgjN/6i3aR6EzfEp1iU2Hw6d+PkecGYHeVq5JN9JdlITQYYD378+QRuOyakO+G
ExNqmEjRfNH8roc3NFMPDP0wF6hpGTWxeTCFBA/YYROrJ4vN00mrnO9nAJycrxqFHmXNE8BOfkbY
IlQmcW2qPD8iYYjYT3Vs2lTtqT1jDaxbbIUEOnyOTDg2nXz1CiTxGgbd+21l6m1a0RHn1Rg1FSn6
JFYyfBlHt1NY7qtjDFj7JMMYltVSNpSWevoq5AeHNiGXxpxRudqZZl+Let0I9MiIKj09LhFpj5Dz
yu1C0GOxc31yD0ERe20XCE0NkyQkqHxPOoOwxPKDt/xe5qyM7Cgc8me+xfmJWlP3cmDf7/KeVjMo
SVkRPBdKOA0SpSqQDKB1B5jgQpRS+nAEc64OtJXxo7+pCiDiIBT2JF8ZvZxMzqch9xPVmORrJ63s
5Uwi6ioVjBZRzFvhfF6UCotEsyBIrczfCTHP8mod+0g4ZVXvBJj2QOPD/+AjtLLHItCfh6u/TbsU
XWiur5j9IcYb1OvE1gemqMH4CuUXn+R9Ibdxm40odz94fDgGHXnD6cxu+ftB4T0fTGOB+dypLwdr
vWNrrK6kNOQrh3Rhwd7ct3fyF2jIUPKupbbt74u3Al8hhF8UBkaBQretKXUJkzoGKzJFNq6zD0Y5
9t/h2L41QqDpiOtjevLLkfJywS1gTYYWGpOy/FmjsJ05D+2gNWBAkzULysE175FghqPDKLQQvx5b
bV1h2ySKipaTND8rGeWCCh8FE9EkWRl/p5n6AzvH9rJqWTTBeazLeBSxZjjd3TJGfdbiurJJ2Fux
agS9V9O5bd15o3tz1ogAcc8E0M6swg/F7dtk7dBGnEednhiLVuE57q+PV3PXDzcxY7eMmIBPRm7F
Usap9B0s2RqyOGnya+AAwVL4bJ0qsjlL/YZmPEDIojZ03CgbL+XG5l0kHN80wCC3HiMskfT1ilVL
26n2Xqm17fwz1JypzsWMFjpL4/C3RFUww619PfbgeA1dXAYGDEGdXMkTcucHMWFpeE5S8d2abQ+C
4fMPO+h0FatbQTUpDaemeKTL/RSTIM8TmVB/d0SFDyuiKvxt14BL1QKr8Gng1ejIMSAFxmU/K2uF
ymyc+A4SIgzz/PvglRlakVTJIYEWYw6wWWsKbr3rouHNs6ZeTJTY3PCeWfBFytXy0uqCpwiK6lMj
3AGDZt7pjDPBtIHAIxp0PhHRXMQZMxDsnqQnRXMD+Tftmeo4o5M2ZzrbCP4iMkyuLacoWXrBSXFQ
eRWgt3z0wSVywS+0NBKJfsmqmAJBGqZ0R6M6Omy2T+iA9NeJmoNnrzZxaXZ0pvGza4PVgTU1z/Cx
rRsE7sl0YepqWWkVG1q4O38aFV1OOKAH1CriKziVLc+AredWoDn3ANzmrQv5xdtpIM3lbjIBCCT4
qeZcY8prhSkNtdSlGOXkvhiJ4A0rr8b9/ucobin82x4V9974/h3QvP9H9rv6m1I9684yQJSaLIIy
jguByzSlzpGeHPHRHnNqFb/Yo+IYQwyYOjrPtRXMo64C8jMHZwGNPstvU6uI/JZsSKEQJ6TQA7Uz
GjkzGQC95VVTHIDP3uZnDYYDvKXwQjSo5rnwpfqDF+0LmMfvlRs9r4xd3uW3KeE6O5zpnvlIAI6k
BWKSphFXh4btjofK9mzxjnZrJ3iNV0D5g0SY4xxnDX2H5YtqYUq/svAHc1ATZMP50M3pT6UOctWn
Aa47d+Ssw5+XdaZXtqLVohpBtSjtIEecblS9WaeNkrt+/xpiLfau9oSMEnZ0oUEGmdGj8Tz4ev6j
E4um/7WwjHQ8dwPwJPnuJ7BNU74rXDES+OTmd7Th5cZoUjPjd+9qsefL5cmvGyKtkWq6C9QLneUS
OGbUiayivrKYtEjQv3O1dcEIEW5HtSdJOI2tpKn8ZAOffmHfq5zfHTc9dfrmgjjljtQPobwHInaM
POHi5K1BApamqkgtIeb2Q3klLsqfhkJfwa23h7CN10pLzcrJXXXa4VTS+spUlGo2ED6CuapEz31n
f481LJMPrILw1+f4qfOfrkdkaipdptzlbOgkuoIUyiPb+knYlir+Am4IprSdtCmfW2UiC1hB1e9w
vslcw4HNWYEJ1B5NyJWKz6sgyknoPBJYRtGnPmQpB5qfvnOQvAeYXNWDcK2n1AJ3StFuJr+Kjqd8
boPesi4HhF0YsWdX0CxmgyaoKcZ9lTAivBNcVjDg6ke/KD/UgIYgvy1SZp0FHpnR8C0I4wz4mPYV
EyfXTm8y+qPB7Yc4bm6BbT4BzykpnQDTNhFAG3T1O7KKbOcuSj9ywUsobMm5bg+7GOZjCI5YYzfl
5ZTRAV3nsGbqPRQT5YcLj3mY3SFmyUllrSFycXtgs1KvnoWoyFvjbMExa0FDfj60y6/DYMQ5wj6L
EJyXoDcQfR/IFnnZbJSGpxujYL+SKBfAx1akGIxV6FA4jog+55yfQinUcuIQcRUWO6sGbBqv0ybP
VAdpwpjnrl6srpFNIy9t3DZx0P8HXgTWLh1sSTbJxko8xViR/2FfZKytydqxdPVNgAE7W8lr9tqj
zAzk2M/xiv+VQGRLcBW4aUnteczqAEOvUpRFtHsvxfpIp/nDQuloc0lTtqa7NCWp6WApiymdu2JU
TYy8MQ3wAAOZIHgYM091RPlZq92E2j/6uhoYNf2h5BNhXYyYdEKScaD3iJhwPuwy5lBIaAtZavGW
aBDmIy+9cknCffOexGxxD7fvHFemgUPzBxDL3FKRgaVu92gqhkoyu60VpcnFe81xJG8dJ+FzFpoa
xNCut9B/m7C0tyL/BpmcI7w7pzKz1uC1lA6uPofjir1v6VmfTjLp7WygsmD4H/YbDGuAxjSC2zbV
nBOTsWX8eWVEKDqDj8IHK1hAuwgBJe9jA9mtMjWtK+V7ChdbKPmNFoQuUuyBLrKKoI2wIzz/kcei
oNQVaP5d4o4fZQqLKEUyHpLvJWZpltgwf4BWaoEaZBP/qwaWFGqMX0Er8mLcndzFIN++lAou49sZ
UWZ+dlYffn6JiUVOORrvROkR7cHqIiEEEu8GKgN6v6PXoCgsKwrgv5ZYdlOps5jjQOKqeqp1hbBi
YIERiFDKMZpRM+oh+HsNE63wbTaq33Hcj1Y6vNVDoGerUsBzUipspjj7juFUiO1090Md7ZNcqd/Z
nyMsFsCpyMC3obHT5iWHXC7R4QYq3r8KUR9EID2oxFnrr3cF+lOmuR8PVtwkUJzbVnPDYJw4Qtgk
6TcvpGyV3e5G5MogqzB1uerQ4Xz/fHTobwcflbJQuH2eSw97Ps8LZndUNneqBNJVqZH4IoBbWqrr
N21yQyQ81x/bzYWzFjOKYKqZryhuGL5ycO24kr5U9BqX6LS5cFDtH/3c7ZZO1WqC06Y3f4PAih+U
L82hOCci+brpSc+/NlmiW3hjgtNSbvMOe7mfqGYxHHcPz/JIVuz55ueflbkkecQv9Sct/6HV0RTS
nE1EiBW9o96dztCiK+YsIfgarVtDcSshpnwkg6GWnuXV0yTEEYJoubZNIzBN2YFJWiLOFrj3G4bw
RNMWChH5PHdSs/79NgTmTgi4cAIzGqzk37+FX2eSpXS9k8Oa4t30KOW3H6SuzSZRNnH38jSdlwxx
auGWVeuk8xDgwgGIafPe46fl5OpP4njM9lmtWZPgt1OVizqJIDTjsEpywX97nLk59aoJ/6cFlhMI
cPBQpmDqUjFoFNBYtF2A3RYWcvwVDWU4Q0fUkPIrOwomPbIl02tNDovoYNQpWW6JsEWjg3uhq7Ni
NBuZ9oTIvFlBSKfanuu3nkvc1LOPzdl7pODaZwyI1h7bOe8bPVQhk8qVfLuUalIxN6gl2Km82JLc
Y+szuVBOOIsIWLlSCdU3p2Om2oyKUp7y/LyS7GnLMljus9xuVgH57pv9zEUcTCDJmGkdCUT62xWE
wJbEDcpTS/reIShhcRdn0J+wtHlOnzrzaQCq5YnhlQI7K76fo5SgpdX45k8BLMJN9Ei6YWMy2V3Z
6Lug/fgxrVoDQCIm17mchBN/3BX6Tn7THz+opVEEQioXTwCnKWmFRdLWEcgS8xjRpe5m5n7ZxcZY
FguKB67nMvWGLQC9iWAZA4Abddr6SssXb+04MglYYtk6u69xI3MdC4wcvYFyJj4bp2ZFktbD329G
NQVdiJERHSvJ+Yuaqsw45XIZHJoTmzwLCTKCYPbgnsaEzatwMVZ1vKXqDVAlRcyDFUBc//VreKGX
pBE6NsQLT1h58Myz2ajEUg8ru7HiveDXuT5aTBB269vTiUziHOOokxq8b11KqPvD+opggDttm3js
ngwejT7afpCooP0wqZcWEmVFPD/zPoDhF1Ji16SELaZKJyWml4xHn9APwRwKFREVqipKvtBqUsFf
YleKc3izzEX715TBQWbvLgJswN2vZEadu0kpQoIYAxVLvTqMx5q0dtNf2sprOGq2N1SM5DG5+aSp
MOs2zHtDb04D6ceMgoEC1PAsPj2+T2DTp0EagAQHneJC+mBNX5VRbkrAohM/krBoNXCNCJopKctG
KXVB0zLmSdYr0cSrMiHul5GY8qfW/B6k7t3QKCzcBuXFaEo/nXzkegS+OVup9tUEVboP64Ki5gbP
Ns4MQpDBlVrXAaasKmP6oqY7TwaGPfzLEQRqii7cDcf0Ke0TL7zi2mI46xrtuxvYreNhwTPKxdRW
mBz5/jq4x09/tL7c32jrpQSz4eLSB4ERTWL4WlIStlDlj5q95ThbNjH9NcbAy6sPby5HbNEiX5XE
nEFxAR1ei2/L9THUHtwz5l+w3daM1M7xZLzzejYpUBeJ9wvW+VSJGXDN+4ksqWSqNpjBNBnphpbF
8KpXodBlIys2u9rdGOhBEWyuHVivIFh+QKxuYy5fiy6XL180k/f9DEQ8Dal95YNb272Q5LpFztFB
ZQBwCenFUw3a75s2AatJ1pZBYhwbjq9n541b54TmwD92zXrZRrKl4Chtg/YKgVhxxAKeTkb1dZHQ
dxdGirsJoXerSoZzqglCCrofNh2ho2gglPkge+opZ5y9ZOWbr7tXj/Cc6T7quGX/0m3FUfBsZb/0
y6JZHFdwh4o0ltwA/wwkMu+loGHfwQLuuKjN33Kz9d8Z2qFNarAMCr0NrzU+OkMSxdTzatT+sNwR
W1zcDHM3llO7v5Psk324DRNYXbSzFBpo/zjIF9+3isyp+2Ia8v65EIZuxU6Rx9ZGmele7n+u7cBT
UITq7oyOSw5z1C8O+6wjW82eS4H9QbK+g2T8m1mNYulodyrvA9uY2lVKqMe0t3gEdbvKyTABjWQA
TQD/4MazYBNJaZabpCRI8rnfKJRN9YT8lh9KQfZTsjxq1SaADMcZeNsjsxqj2WoKVZSqiPHqZF7q
wLSsu1RY8F2fgBNzEZRM1TDUXnj01v08/qrWs7A2iP/+XvtuKYFmc0Ychx+TPsuenzOmCaOjQ/h3
/fNequ1P0zleVtRjVhTYOCyxT7qAsQOVjiRVmKF4+dRVe/sOjIDLsSDu3W5ueQXUFl9ZQ+pHUMqv
FVUNXll6lQnx3Kv7hQDtS82oetUCIfSQG9txbNgbqOoPm/jg1Sxbv+4GtozGCPNuwbc7T3GgJ//u
4kYWAVd5e68p3NyFHWe9Ih1vHSfsT6yOy8UxptV0q+rw2ddX6sF+J9gwpcX7ETbWJDR1wlfDfFdM
IJurJiFbHyzedyPU+GvAOBffwuG4fR98htom/CcLG1Ysp/gjzixuOwBHuFQLTMlwguU6ZPg/gHB9
OKMYTgqbzWcpAOFRZe1SXUjBgWwYKtBI22RkTcDZ6iLmsckrFosuatYUCoY3M3qS4SJI/WUNYWmn
cgJl0HPP+kqBsWBx+BRqsIVgNrIHi1EbK1zNNlzlcZWu7HykBAEjfetnf7lggK0JBz4jPHBOm4TM
n/kJ12MGiDbpxSXAAwJUo74NtKpeKqhLcoV7z4hjXedKt7PQzrKEMYUw/hXmtpw7h8Hbv4oTWFFl
WMcQNQWaYkdRbCmJ1xQ0qBMc8ncFHd9S/r2mxJP/KT3cgEC/lYrXeO26TXQEllWt8Kaiv3BwwEve
pMWmPd8KgAIgPFSCzjXLIzxcC4K8IScT2ThKJxsUqcS3Lo0jX8gRpD0sIMnn0otzQWNmrMKBie9C
VfqbelhRit8v5n9Tulp62K9vPpu5XHKir8Y3ufvm8/gf24RrKvFBxF3IaBQxs0CAAS//0fZph+lh
MbajrEBwiX6yeGXfPdZQ1HeriEv6q9VUYG0kC7a5Tl9DWAsgwgYJ1CimwU91cE5ABW8T7xAxQ/ee
KYVJbbwFxGrP1h7BnhfhhrdwK37uQhkTt3OJeFxmh5JXG9couxyJYvjlSyUhbzFk1QkfGmrFDoD9
uQppWcKAAkPxXixz29jg0F9vf81vJjs7xUjN1W8TDNxWezGNYOM8TNrZ8IsBWe2y+n533umM692H
m23glXR4TfSobbIqChJ27BlzxL/Pa56Qf9rsebit0yRMSDUI3qU40TxqKQKifrmTuAUU+fkadpxj
xYhrab8pl72roM7gcgYv7lw59S9TZlNjNcjIztHRiaqX4bv9pBB7Oz8QIsiWG6lDWbk+9ZYwGDIX
HocS2dJMT5r7Lu5uiafr43UrV85yUVRPQeKwziTSELt7BFMW3Hrc3YNfguxzOQhaRK8cwr7TXdxE
kJhOZbh14PuvEVOt6nj9l+G36ykKUGIlSMDrm7J2UHmjZBHUrmXoWfNFyGg63UmAvpvdpqUbc+J4
fT2JHnI65DrRaqQ1YuY8kQEKDeXyxVTdQ7pQfH/4hNf3bKhG3CxsBjuIPv4eD1D2kO7UJvGdx/MN
mUkixOvUmLKcDHgNb+XVjGh3i1xF0GGZ7ALXq73saKnDfRGIlJk0AVigc8mc6AoF3fPkyRHGaMpQ
1bYfdWa+uVGq7zBVPfX9HhVedJPg6VL3hsbYUF9W+ZcNLBcW4JZeY3QE8HZtu36WmYp46C1eN4Sc
0sgZJtcsnWaZ/XgVyvh5KnBUv+krR3yUuGIUJjFtsnhE5zcCtSs5fmnNZ/LqQwFI3sBORaUnFnmW
Uwkt9m11e9YD/vfPG9sYcxApUBoyJo3FIk2dhAub3cpqSpQJVmim5icrg6QvydWFZKzcUXOR0/Rc
MroKQ+yfVcjwiTwME3cbl1Wrjygj0OqhBeed1vjb2lHpTKijus8ITvDKO6+f4SL3k+y1+56NM6EE
srDO2WvleDMuyIaxuIjMh2kUCJE4vLlXako+Vw24cS9e/HbjAbq8N+L5zODYRLd6coZZGLJRbZEH
/QHhEiOAy4CUw/Yvei7sgBnHSzue8CDo+k3OI0xESwM+Cu0s+Da6/TO+V/70f1H+3EoEjnvlo+Et
LOF/aAeZV4QSVSL+jVDwYxEalyjxlgqLDYi1M/XDY04Us6wjHiQ1LDBI3ueKdjXd4/R4utHN8RbE
nK+TbYpLr2SAqteR2P9rwFwm8uF/j6zOad1DXQIfv9LPgk8Et3Fi/NJ9Na+4hC3CSPUjWGWQfx0E
Luxko3O8rUOLP8T+ucTkbFulbfwyvDlNnV3fruGWi5wIiGCHIVfVdtcGjewr2pGF49VqAQ8Y7msF
quAT/ParITJWJS8/YX/CCLt9rU+ES48cmRXwcTg9fitPmqF1A5U0fcvrnod5nSYD/ObhgnK9/++7
ZtF1eAxB4VeAYdgM2/QEOrAd66C1LCYcHXXztMFY/xNd9rHHkN97mC4/vnC3KRb5daVuEHysLRlk
efc8qvDieo0THabiutYmck2/fn6iDGu8ZYUfqKR4bSgyW7uszwUnDLUuRWXZAxMrTPO/y5pa0Jue
7BWJlSW0T/EIJqVVnqmTlsZIhD3YjTdqMuus9BSLVYdb9hBTanHmC7wrHDNvurXPvtp4jwK97IfD
1QsBpYh/vQDu3Q1DM+vVKdmv/W6VmU8pX/OG9Df09Az24friHJlcxQ/pSCu37hJJtszy6pbFDbA1
iLb7AG9OoHdKWtF11cyIpkCmSDy4+4A7KArjWPg3Bmt6E56+TzPlLb/9RH6/G+tjP7d23IM9M7WN
uy4dVLhXCr2rz+s9oCRRfFY4m2xEmSUeIRiDbHbiGu7fs4GCfIl+IeFguN1sANf+MtZ5KQ++535i
vTnf/4+NjzHLcJMnpx/QJVGQXGkWYlw64v71ewibOHvuNROjF68r6JuawduLOQH7aHVwRYKSOYhI
Y0+0X7uY6Ox1zfHmKQFS/+0jPA26emnHbZmunnoE8uQyZGN9olm0RbnbNpg5stfJnY0WJP2sHhGz
rJTUQv/0xs2/absZhjRNslGMl84ooGycCxmvynv+ff6epmH7I6ONjslEUkWgM0WLY4OGT504cP9d
LxP4RTnejOxe6mzbsPjjv6FCoL7Nkotv25uVbR1VV96l+zW18Tuzz4BtnmfrXm2CbBS3V/I4es9H
YUlRI3bkXPqOn9OqOVVY83IfLMh6HEjH3zWIKsZRwg0CJAwwk8NkWIVQeq//VI/HbE5QtY7E5Fn9
8zLUeUJVogdxIS3Shl0BuLS7f5kv7NW6NfNud59rOiCzaPmnicqMfCFDcLwPlJBSA36zz+Yykcuo
El49COsCBkIH4/bitzqMyFui6/CqsHPWcpmJO+lEugU/LQQhADBHHJTlBiAONNkx7LRz23dWffV8
IPq8jU90SGNGoh5Llv96NQErvVbbn/3euKp56pcJDTzFgwuuiRdvG+UHJyI/ZmfaIPftiRay5LAx
+J4JzW1DNzdJzSlk6Qdev1jQgPr3HUFa59MZq9J1yzgKQvkFG42ooEaQUm8IoNbbnNV/vXSuY4WA
PH7p+S/RhkiA8+JEi1ftqcGqjzFINCY9EZTsHRFiyYeraZx3rxDSg8/OYsP9/Cs0Evx2x/il4dk1
DZxAkO8Dd1SNkjsMKi8lYRkY6jVpq2LbQScSMA2vIEc9Lc8HdM66Jh34SJnJRGAgHtqU8nZ5aCfe
fleAl3RGQZM0pEV2bfxTccMZN6wGjR85B9RG7KiiKKuHBmSJHArtB6HUQtJDs3ITxgd7oXUWhvvZ
NzniaD59J38+ComhE9mcRoeCRBeYVOyGQYDX9wIElqb19Zw605jxwTxzDLwXcFxHkRrSnU6+lEnb
jWbfsy9eAo7KyFx8iaJIvLOUL0KkE72huDHU/wA9S1xjO40Jwp/KKIK2apY7UJel/BNdVd9mxI1z
iKIUZTmJ8K6fzaH0De3ZZJRlD7PtBd8588S0TUyA/38/k8IIxLBhbLkgebAmTuXSOcOYO+SIhzER
D1Mc86Hx68F67mETK3GJHDWPkbDACQBgYkeLyfGz5oCGycLC5IE36MIgrNTEzKdZn6vd1iuLiBlo
aHG7D0+nzbWz14yqgnfXjiCkwLYTn5QwkxevWmIBed75BJqxMZ5LAubQvxt0JHl2C5CTYVfBnKra
sOJjewJlYdTBCjbSuQMFBcVQZhvmTnzYBV4c5TXerBOT882O2pJPEt14itlZPyyZTAQwLNO/GVoN
/e6BT2Z4h2hBfQv662SXq7LOLto+UOKL/Jd2sgXvWdxgYvAk0nJCnjM99nvqWH+tg/dGoXr3r2DV
QWXVv4CIbhrk4vx9RrBtbxO3W+kSvWIU+VGXLOSMpeJJ4TqZ6/s+J+BUqqmJhzIptD2kLFjZ32Fd
RUIC1tBrjYR9NBEXzbVY37qzcpcc+dYIDTDSUyQEg1V8rsi5zkr92WhO9wbLFKvomZNaHAh6nVtD
HK42YjKjz9a2jQYyNtoJnPa7nCPhBJU9SLVPwaAJHuch9AAU2nEm+OY5BL8dPym2QJCsrgV1wnS9
LRKrwS2RBvPi4b6ZU3NV5eOKHgoKK0BfaV56+D15As17WAkhacS2sdhRhqQqOAbtI1ALVkJabeSy
wun19qq2NdYii+7Ah+bafrdYukyQ1JjuxUKe9jwtpqNtBMzpZb8NtabG0pqMzf3R9MGdlFCm6TmJ
zFQR8Fuys6fH3qnEdJrQozzDTUgfH5pxCYqtWaAA8Z134Grb5O5wOdfdnTmo04d+D/d59Z5Yx/W2
OSpiwl5yGDkbPQJ5NGKZ9O8Iw0FKJuN3T3Bt/bmrnFAiCMaZ3LioBVVsIU1jz9hduBzDGhR/+JSO
IkV1zk+ToCD/dY72eEBKhyGiB0N82O6zfTh45FvZdEzLlmPRORUPo6xMNoNZONkwvBDOzqK6rQBM
xjlMI1Xlo2L1/5vH7pCVW2J4C/RGMGm0kV9SadhDi9KklQbCaQj4VVY6XCElGPW5tEcU3XHY/tCD
pqCVTvQhX0EPi8Ie8RPyLMkTPeuycPxnEnMvyw+wmNIdNd/xnTB6+R6mUUwNry/yOQkNr3NRRKFP
EkuXPpPN53YrAU8G6NMDF/M76R5iK06WYuNHW+7Jim9lRoxbdo7A71nmxc6E/CgEQGeKF2uaz/GP
WvaAQeKmPICxGb9JAY+9B1KubjqS7Ku9mKFhQVm5uTGG4kl8Ky9K8IlqAlm828ZEtgvPUsvXfi3I
jpi9ShxlBs/vE0/0IJ/FRgEW3J5+wPUT4tg8ABARDeynt2dK2exFkdZAXtH9n8tV7qa4iIc56ZjC
Qu9UFP0kjdKxu9L6w5fqtBCjiqeAReRVN9VDTvX4GdNzWQJS70tTQ3msOTpbiYpkFQpkJ1hI7HwH
5VZmMgu0Nj/3Eil5l3QyIH99qBHd+RRO9CZVT8RKtMs2UKfNpq6MKIPYAGTUxRMH+NQms63wcdxi
vFhVA6G5sdRxK9BgsZQ/hAlJ0PsmC6PTVTOBxMKkyoanAUZbVTVP/hr6Vgof4gk88ijeqC5xeXCc
PEa4z7O0givj5GNoeuKR8wgZL/5m6ZeYUGVL/f1G/i7FWSA299flNzjf0zNQwAaCtZFMXMPq0NGV
yZvob/Lv3O4iq1vAHG0Z2yCsdsmGHYegf/MHKQe6KUXKJd6Ks4u5GI/PvCQQZmNL8292rGGdkXmG
MnX40JzoiUwwVuGtnDMamTbcdGz64ueZ17/rWwABNErCZ841VyJptFiDCny6U11k3BePusX1XYTr
pmZT+rX2MReJgejZvmwH8T44A5dU2kftFV9iv/eLCzMwXPwleHuGo9VCkw+GM+Q/qHVNd8ISkS7F
TqUvKOThSKVKJLgh3BKkEL50EaCQyhCdI4iyl9IPbVjWKW4dFb1wAOEHzwNw3aMYI0MhkGlM5XYL
ciLxLAuXd9QHDRdJg+KDMrj9Fg8PhQJXVoWI+znhumPhCjLCVBeOT9TV0GHb4MtMp6BjVzRuwpG+
soXPnHuRNBwh3EVKsxFJz5Knxwef1q8U7lcYfbFsZubw7Jm9qg9HSmVgWt6Sv0L3inciqN0ECENc
DMlQ2n4Cyw6IGL49ry30U4tuWCp3THakEkgUJ6jdmTGflGwTNtVSVIc5wyBQk54Ho+LcLIhmXIek
5fEyI7NdShVzc4exAhtu9xm0VBUGSq9bCRYwFPGQcuL+/FexgK6vEgW2a9I+cDJHFS52qEYE9c+t
vH9lUUujBpuPbRKpR2fKjfEoq/ize9qvSG3QIt9n09Uo2c2uzgJ9MGAM0ivpI+jLHvLx3jevhI+T
2f0XHV3u3OrE32nG8Kw33hl/2XOKJjBNtyGekpYAVRFDp2E09NF2nqt+g3QLLhtOKDwOqRO1Sqh4
0/3PElKmfezrVCS+GunlBqmOTRoXzjT1fcxxmPGb1SQLuiqh3KnYd6bfQYRb2V6qbt9YNS7CTAKB
uCJqbd2+vXCWHNhZxhuV4itya8uzbAvMrfLhIk+A1zIU8bAeQoWH3IJsFbNsmBvio0VPSz/9SmhN
8qR9Axf5iK4uCP9EH8IGatPDcJiCbt4VWwXYDO5JdmWIh0mFRRdBNJVtmQkE73Vl9OBzFMqYTQVq
l9iv/Q4wb9n/XcZHFH6dSZTzQ37WyqWX5f/YCFCG6HmX898saWT3L0nxwKX3gWTfuGnEoyW/xa6E
s9NXDseTWcJUhMQven0zNqCPqF+t1TdkklRMtU0MO4rtjYiZuDvaD+Bnm1+xdEho26KyKab2DxHQ
r9jC0b5U9WPtfa2WqebIwnl4mr3jbgD0QDczMfC/Y9FY/VBS3d9s2NZ0OWmLrurbDvWcQkTMJ72t
V/0hRUouOse6+EpwhZhJdr8B0pOI8UZ78cjwPcj0i4bp9masGQUlMSTQcGk7KLvR2MeaZYQe59uz
PCaWe1f82oxlM8KYFQrDD5ojfBFiy0aoAN6oBXLulze9X5Dcv4me+m575uUsCUIRn4rSlgFtKgTr
PrwuNdLN24umyDGuBHoYOEy7wHdTduV6J3GFGg9JH/kj1DXsJei4n9fKMWMg5Kd1Y74PZNAT/jEa
E6LvNYVmCT4PmFU7RY/TckSKwYPL0l2LfV34SgPpRLrDMFk2vV9WimaNeCdJccjdB6xWoJr/O/iX
TrvSkPDkP2TJzKA7VCGrgmBUZL/w/EpuOXY1HlEf/Ne+ywScN851E3cMwaan9d8X2I4ETt6kKkve
S69c5TG0ff4xh3Pw5XUSsdqMVrgK567JUrI8X2hZ5NfDajWCUI1+MF2baPC4zsy39X+JSyZh7pn2
rBo6zU01loSuLDKXxIv5dqLjQgf2e+rSIhRFkEEAh3GYFBIWjszpyPku3VJUuPUYxTPW6QRDKbK4
LCtHkWYswF853eH9dIVhbE4gnsRJ0hRqvmxuXFBGrUTcBPLA0R7WbWcDjaZOa/3ebzEIFmWVSfbr
9BdB3u8q0y/rzGCvkt2nodKj7sIi3CBz65KPY1793nw4QCWYc8FzxqxkwBCwl9Gm5ftiwVANz01+
iiKp1Ql0v0EsX9uWUI49MOCy93fm34ApNBu/EoscAeWcpuujFPm3sBcGIhQGSnHrqlMCoQ68jIA7
5ICLclfX/3Y2pgjyDhqJllYDQSs0w+3mWeAHUIW4TY6i4JMULVPlgunuk9mIx6Xq0D8be9JNKW1y
VTE1n6FSepMJdTE6saGUBxNuzQQlnuQxVkcfO+/poRLdAMd4e0uRzPW/aYyDbhauQ/jet9XWn1lt
BQQD1lE0nqjxVx5FMD5sAP0rfxPe/We97hj1HN0NflWonCxrXaO75AefJ0rVWa9a/jWoq403p6Iq
X0wLIQ+TQw0hfPcSEKpFXovniOZ5hqzxx2UqN9YjP9gAdiNluEulk7drdlB+jNwCazNoNhv/nsY2
2T3u9cMoLjO5VIKLex4v61Y3Kt/cGjf41WcJjvFsfr5zISVUF8gCJa8bRgyjS+hK10+D2OBdHcDG
VnMaDuBj11kXQSKZtGvV+3hwR6NrjjLezEnipVuJxH712GPq8aTbpRFAgYe5toxCe+VbhR0YwjZ0
noKp68QuE4al3j6fjFGHs1UOIX7KVBkSvcSbeEbYtJ9RBpHllstoTGTADuz7q4/v1OngcV9srd1x
NAYfvB6CCGrm2vRBz5NUPqhXeeDrzp8RO8VHPO/q3IDoeBKBNx3a72eZfVU//Xv+JBSW+mHgc7Ox
R03QHHoA3shC6JciihdcPQupfjpo9lSzLSXqkpYUK30Af6zQQHQ9o6IWSfNYhpu4zlygHNeYmqgf
Zyk5S+BKTzfjHlwyFAZ+yTqE7UT4q/H3mPzOpJPGoGe5vpvPDI95jnvnBmbsJl6J+VsvYB2bPTsz
VHUjtPMBkhnH0/ViURTG535RIypawG/eYzVWJ2mVyBR1I07VzTiNkCAKjDcwTIunOPooVhFZXcXd
KIL++fSaRyFUfYL8Hyxjiv5UFUWASCgnybIN28m75adj01YOtkioAO2nFHRBrcWaIi9OayUrOO26
3v23FGADmw53OpujrvxUA5zTe0wGFjFtBe4GIvHn+mTLJg2REqU5lIKndgWy/RSncIkrJJnAf31z
iJSpx7udKvURcHtjDFUx9nbU8BIr54x/9W0E6JT5a+EMcXW/QsXV1BTxMmc/kRFesUwiX8n2ZljF
WufvfKXNnCvRb4CCM88kxMYR9bYbGcq+JngWZkXkj/5VJrXlet3un4xKMEN0UKtyWrfCa0AO41bg
gkUN7P5ZawfYI45OUNfWMRVI6IV0tJif1JAWs0AWRBkrLEUDF/2qK6Mr0ruegK6I0m1XHBEDAq5i
UZsR1wHCtfSY89hf+CJOGhlJHp7SQ3NAT7KxpU2ZALKleN9azXpK9Zi7DTAX5SI8+VgtEbcukW6c
nEsXy/SGu6l4LsE10+q/77Oc6Xbrukr0wcu25kYMGmDpw1gcNzHE5qJPakKyjyz7dCrRuiobrhmr
3s1U3eKVrm/hWL672Ye4m0WZ5Ql9PLiChQUcbMX/AA+IbxlwCyXWmo+rhE05GTv/gMdus0NLF7ex
AVKMRS9+dum7glozGIkC97LcK9vg2Y0/wI/rX9Fk0LDVhDS47hcIFrifTBywDXI7Lpt2EsJ4c9c7
OctLgVKzS1SMLyoqnWZdSonDBi2byW6cVp1aSd09rtcEuhH3IXAc+BTtLdPxiEdarenLREfgaAPg
QtZeBSAYmPMwihl+B8QcIyxd4BWqI3CgVGh1N2YE5r1aOlf66AyJfSxj9kB3GqfZodEnlGOE5Pmu
y9PGm/msxgbdNvzoJ9pqpMcAe0CFlfDDoPkmUslVqr31XRIx1glxVnkjklAiIU5vuFubGD00gSAf
koC2W2M8eJ/DMtQUoEHSErsUMSNqSWEowVZqYEtXl4+ajGC60hKHmrXl4KfXPlLb+2/D0uJyU5Ri
5HLorUM2MSXDlx7nP3CUPsVdfZJ1N4gGpcXAVZLJ05tE7dlOrJ659IrpnBtSFBwhdIfLN0i2bLzI
Fiuulrzyyedu3RCDINBOlba1+cOHkvNHSDtdp5aBe1LqK/nFRbJn92SD743tp4IuBlMIAkS/UMrX
R0zSkiQr8Ei0j1TEnFnbVbAUKIqFQBagnzZuAQj5a27aVLqjS3QjfgQo+J4m8DyUj+ElXid2HCAG
5xZmuihQAmgFZ9f5qO2vsjOabcrlCNk2VX62E0wrBHhfiB3e/P6MjIWC2ZKQyZdrN8inf8UwHiOb
HlEqn7BFlQNZ6DahzrGpHQuMxZk/Ltpx7VVMyC3v/b17caw042rZGisVRDoXgx355FaDchvTuxQl
OdgDMH4m8svfeUhvrhUDg+qE6MeupsqzTKxT8pGRMQwnfOY2eb0Z8fG7Ehzf4ROteO15Mkg8Qe9Q
5W2UeyVsil+DzjTSKuA/qfjV+jiHyBh3d/QUhOrgXZwMKZudDZ0JaGOqPskHZ6DUGqDOnoeakhrE
1Pk9Fk+j+KPX3FacWTwLQGRwl/DGldfDahy5oE+wl3NrfWQ1kJXdaHokCjgrakQaxoYpkVP5T1nn
RIBQiswxEoFy7V7J4wKxEkDAM1Rn9tvIlWIOOMTWWk4iR1ZYW+3Y//3M8joDGICKU+j1IbciYXui
47ef9adCNyaVIotPXwgPNcCPKwEG3WTuQKW81S5toybdpCNsd9xUutpxBuBnCF7SfVOmg0Wp2oZ3
q65fmjxZIgw6O3ZPTUEocBj3HAc+qlohbzAobG+rekFwpbfYoHH4uHl7HaA9QwY77NagYU05gLR2
/X0fM8Sk3Xi5vEddvgqGInbC9ajgf7uFUBBHHiJM9m6TAXPKeGcf0gp1m8aKNqEZflkb4s0nklg4
hvlAGGp50shirmd7s8heJa0RgaRIzkwwhH74EudeA9xx4fu8NJKdpw7mUtLUtRa8+0LyTjGxXHlg
vfjV+4frZa45489i1bMC/uFbt0HGqe1R5YGfbJBRrgVzX39UxrvvKkfQ/n30ws+lMzE6EMvg6918
8RmrHGbLL6blkwCWm6HB2xLSrE+a2XVoNxEZDrYuLk27xUYAsmCr8kqd0PKFDmPaMHG5ByfOIJwi
AaOqIDk16K6Ng/Uv95kpqhogmydMOB6n2SNnmFayeChQrSJd5obNDJWILV3shvF9cLlJaJov5yW+
8TQtgwzoA6VbttSzeAaTm0UGQJLARkhCikfiPeXrk+gRZC8fCX3z+Xq0T9FXwvW+pOrjdX5v/HC+
XfkCIr85snBWTTKXblhfwkZJ2hjDXlQqA6kjC2Ehx9GTnN39PQnSV6BJMXV8N1g4pMWLVbYCC9p4
RAdgQZv78K+pi4MY1FIQlIY+RnZuRk9iu/wP+eTkN6Xi1cYiZY+8iJuLibOKIOD1KjsdEaLWdthB
K7+SoZHbptfPwcxI6F4A9QyRsX+H23iofNI92VsPsSPeAinIvSgQGVrGXcbk+G6TF93JAv8uQxHw
3gN7PiNMSfVel62+7vgT3/RsKtv2Yz0sKSi4ht4mqz614yUDmHzWUDRuRG3FxiN2vkK7c2PJxmiS
TbCp9YEdmzlt18tMf3qup+ptFuCEqmyeFf/d8D+Bd7PNT7SJUVbvGSw/tckSqhTgDyt2lifmxtrm
1b/e4VRzVUDY4Eyh6P04T1H2r73Uu4sEN3iKkFpQk+oi+71TRudQwimBCUe7Mn8H97ty1+JhKUZZ
tqjebec3C6xmXbua8U4LvpXyHbtA9BvscM5qNZffD/c9kF+B84mJA7DdvzeKebyaDclpgv/zUt5U
NbrafKeYdSNeGnfAXbP0OMiHMEiEbF3s4l3tlr6/5pdyRuSvv04RHC3bzbF6c6VDC1nZi8CHTy6n
otfrCrxfdkzcgcOClKkK2bnLomvuIzegLJfvIvGs/vlkX2gW4rpaPsgmHFisJ5EyaeyKF3OMqPQS
Cpc8HUycLKAbfIxW+nONLVAn8zR8eFObpqBJsfZssu1B2LtV5O/Cz9VuFSAGwGoPK07kL7oiA1Bi
ZRIJmmc7NZPA9Mt0eanvtf/Na4asUrrnHkh+9W3zjsk5gm7c/cCiQ7pxgliK04NUnzNMoYiuc6rY
7FR8HpW48brTvOu5ePianENLEDU37r7Dff9fTDwefdmgDNwaa5ByZHyDYRFFJQgLehSUbq60vwo9
EgLhJd0ZTsm/BMxQvbA81uWrDTRpSn2W+giNv/LkhrWVm/EPc6eGR0GkJ+m0Vz8o5HccxfdorSne
Y/f7XMSer/p/NLihWFw2uWTMRQZH7XC/A0jL28EBwpGaHnmAo+P/hzC2uK37EEnOfm3dbL5rmC2n
gn/zB6PM1mMFNA4ej4BjJ0+AbfpsgLBKtuX5w9Cx6Jm7HpTw80x899qR5i8FcxgbrJmKWGzBMGxA
VXEX06LQ7oELBdgja/BU+aMhPahb8Rcq+tUEW4xsmAKYploPPJsKUC9oNM+NhTbwBr4Cn2qNpboX
O9oMwNp7xxKFHOe9/QbPym0XZFGR4010nksn3C++beqJQDN90qMfsrl3W+sya3zEstVNIDKMwd5a
ZGmaPS2nEvrshrkLflTyH+uzvyFH11f4EKcyMinFrinP6egghQrOtEkTMMUSZtZs6CZGtD+l/Ekn
NO6T5mKH+uvLwY4TIP0jp3R7w4pU2ACrrxbT0u9EDJcx69lRQAoqYZWRwTy1nMCsIdj0RDznECoa
E66hvkfU/ax3e4F324pwdnaDLVWN64Di3hMc8Ppu4yMPEHXJobEeA5Z/GvOoL6VqQsFaTL+BjYT5
dRDAOMg9MD6bcHU0/4T5mP5/gDFn1eM5aqRvSioJCBYDLmHUDqjg/DR9dbB+VSkyk5kgQ18u0s7D
pQ85j19v832aqsCW59VxmUXSS9Kwi3Behw0yD0qoNNf+9Py8gEhvQwRGbs/wz36/ghxoLWi55bGv
afPvoF6jTcxLsbImW9TqmIOIebfcojnK0KdENk+ci9wFhypULA0wSmbLcfWn7C039pjo6yjJWCCq
1Md3ydOGSzTsdtg8flyFc/Pv3PAZdfsHKpfFXxVWCkPs0OqvG3GyWI4w3vkrd+y5nlPjcz227QsH
4ulKs44FwnAstYmossMFSubxykgIA2icpfw5gtUsbm9rUpxQh6SMymO9lqTJsoitWgaloU/WOIf4
nx9FTAFLZdZsBpv22BP33FAttFsgTpLW8Rb+DCsfbf0cyK8QQWlevx0oclMPB+ajoXBZTwdKiSul
ixuCrEc+EUCGS+XT36+PNTc+l2r9KbF/13ddulPYhqBIYJGLEfYfyyZyIAVwMhFV5sLguWU1fWVY
rv2ERYBvrvEecE9DQ8s5AVIa791FoJku7BXQ/Bvb+gJjImVGLETaFOaRkIuLjd/VjPlzzXK3fxtu
VFINER8iJKKoemA53iO+tXZry/qp1LdtJVUbNP57+CjEJwBP6z9pJdppME6+xm3VqCzsi2z8Pdcw
4sSCRnVcc7Sqdt99JVgNKEduunRTd0anuWzWLYqMe9b48kL/kF2uzSGGL+opeTBD9lNa90DZDID0
QHINHiwv6wUQlQrWqGohBqjmgQQHZtkwapzbInbe3s8H6/mxMzVc+ZEq63Of5IHUz80lsMz1A3B9
xZFfvCC/aRlwgX6NbHhZAEHCmY7qp3n8DOn7DxA56jB9HAiCrTnJVagg8esepXvRsfIeWruLDJ1B
wzgPgHvxf8G966epVPDeO/nlR8jSbuglJybZAqS8h5HpDWl2J72TG5Zhyrb8g62CbI1vIgxUoT5e
kWXJFn1VVU/URfz46Rgk/wNQq5LOZvur2EqTZYHXfpoqyI+oC8hz3AibdmSTkgOBtoulwRH0dhEO
HndeOVSnHCGvISNiMuddOx21lMuc1h4ushWQduOSbIICIFpt5DdX9vBwkms3DTqKGpmc5kn9KQtJ
S4PjS8pGHBZOBlfe7sSVMBNalDyvb2Tn0RsNsaLq1bamnEEClTaYc9K4zW7fGsZk40KlEW9fERPL
gUtpGTdGfLBnjcz3ZVtR173ofoZsX5wzN3GBk9Ai7X+eFW6BCFezUTygLHK8+lG7ylWMaWuNbloX
/jGcXn0tJcgsdniOPf4/Q6LnDTamkj31EkiBX+cBApKuaj/jrq3kvOnolWVGeVu7IvHmOn6Gm7kH
Nqk6gfxU7ww7dgwllzkckMfCmFQ2Mch4Zv5Lg/8j4xxXqWEd2Uej2fsz5OapRunRnJ1v0fgJxWNj
6JjwRwVzG6yYUf/kifpT7Jt24SNkH8978HB926ZCaOq+CNZCbgbMyBvdF+abJRF4T2xFo5wLTeXX
w60Ml5rGsrlnS+VyCCpHsR3UfPdXRGpwrIShOZBh04e8fIknzDzEQh6lBQzkkCWjZpz53Ic7vBbM
bHvk/OgNg9sIzs8DQSPuRglREIx6NyKwj3mB8PqVQ634F97CsGCJagYesdqGxYvOuKWfbozD6E0t
DS6r6N5fxJZTwkQVv45A5KI6C5HQV2f6ObaVMnPzKBDg7F/xyHCAFEk5KccNoyN9oxeqe9514vXG
n4OqzzvNF+6MUTgLvGXmHlX0C1MahyctBBxo3V2KY6WRW75uLvCJ1XK9mk4huYJcgdAtFe2OyyAa
ITMjZHjXplUlPlsv8w6t4DaIpJYbiRMVlOKmnqTYdnDJUETo9ObyhODGCHeRXpCPU4aSYKrz7fX7
wG1sCDyHeSUjAbvgvIZpVW7YL4NnfDqUE9v8LN1SUn46G4O95xTw5fLvvL/qumQjQ73B6zE2LfiU
+0B7UodGqslHBDoYAnFFKojlags+kKIre3SwEX2sn90wBWq/hLYjQxenhL0d45yuVQzAuJYvo0CQ
9GaLUX9/TKnS8loqVhatdjEv74Xs4idHB9HxUNOj9UmWftEbgvCRsXFeXtel9MadrXAAKeGjo0wv
wdk6KsW/jmkLVj1+6dMWtR52IExBR+JA8MXHXjgA+r+G+sk203hVPYtzrh3ig9ChKNPiuMKxwonj
hp207BuJOR7e/RV8g13YhP6guDDMFIz5Zxf7OVYrjWtP3JTbWDi8J99qSWTbXaeILh3MOgPXWEfz
sGYhcxaajyrXCf15nQM3xkb/jdnbL5Ft33ZrJbLfzPOvWm5hUzHyjPLkqSujIiADInLmcPpemPTu
7gHhDOrEj4EolOcbvGXotjf1fanBP64r2w8MaEV2dVzfv2IAtDNlw+2Vd7Dd0Fz/8XsV4Bwlx23C
f/XybPaWLcf8I/0nNrtrg+TuDkk9VbBVGG3HLJH28d4ksdgR33CS9Q3oC0+pP0sr8nxchwH7R4vj
9ejkFZQpFcK+ScXGFSYf0UxMZwSv+FA6nxezGsLR0z+mAcq++sjfM5RpP4B7EO+G50VrY2G4vu+d
BLk/wfFMOp88rlzEMwZGVN4Z1byTSpSW/tc37mxXzJ3mTPwPULEDno+d5B4UHXh3qA1WB9SyrlzW
wzE2BQ/oRCzFzlKh8E9EVepF1M1z6t5MBhyABRmEcGtjeDVCrtragcHnRhCDfj1goiWvvegsolN/
vjSKZie/Gw5vwtIAcno9FktNKMqFLzJYOxwQ1eKfEdyx75A5n4zXIBJns3W16O8reZG7slkb1Y+U
axAhYgSBW3qrWdb8JZFawQaHQL8EYn/uUHOudbSNV3rUT8Fm87qHuEgNPVIbR48EFqF/V2+gHqFs
Tr0IPNjfeJ1UerEI8aaMumXS6Vgyalj3NuGrEDC8mNSs/jCOAFh+WTJjMFdCB3KobRYEN72d/STH
+hmm3hgGZ/KXoxPQpiWUYGGG08keVvFDodG7Sv+uWELj2mLFVdGcQWYwISUUN52C88FI+5DcSa3X
9navkYtOQRhYjqEX09uqBEs42NcDnrtAZ/cBwS4d71jCy0g0Xz11TfAjceF/OMTChIgb5HuHfJFW
JPAap+0Z8o3+GLgymJGZw7Wp2DvVxxnixxGszbn4ueqKNz0X9LbDPNPghR+il2EX/nTJ66X377+D
g92O9RnzOhhIiSG8kiKxADUjFkBeyXmjosoOg3x7yuhyI8Pf1jQfOdLaPcTp6LcZuxjYdRhm2mav
bxTms1eJ4irHiF2z76Zu4dnOy/GwEcfWJQoorKR4SCiEe73R63pVBfqbnwFjg/0IIVuVXrG4pmRN
ebWMTZukGYmPGEL5DmEPHx1brfWU3mKHcvom7rPwhmPNKSHyacBa6DF21m7C66ciGPObL6dDbd+Z
oiNQ1GBYQ3E24W+rmWRSy7a9WhEVD1dkjWcwikiFCeB+BVe3EsMqur5bJBh35TtsVKEQk5skgvl/
C7pDT4xp/pdUgplcZJ8lCizDEcLwu2wtPomD8Xxx6VdPOixwFHu3OjQB/JMIwHjCudYe1UjR1yg5
zrlCnSSJUOGcY0TvVBPSIK+8ph7vlkaDBeOjzs6TifW+TVrHO5VjICWlyIZk4+PINApO5ETb1mMx
8Fee+nsrOy763v36CK5M3D8pzIagLY5ANWwM5UwH8GKdall611BB0rAzVlwgLPbnIZ7Mzmv9dEnS
s62ajgGZdeCh7wJkAIhliDDXTa0sTEphNx0C5PcDOB+TWGog7SmZ1Q4zsECydSFxLQL95/dX2k1G
dORfw8dr52sFjnbOL1SEqEbzFEY72Ygat7E4EhWv82gZcFWltLRBctXp7eBgk7ro11CZXDepdx70
+B2vneV66oZyCxsn7phST1RETLjCxJWNkzYrH7IG/VR0u2Yd+SiwjkMo0a9E+b76SXp2ktKjUwa1
RBdEIJm25QJgcAuWOJ9fsB9gNCszTyS0Ql4ijU5WuAB3yUdQc7q0ImL8QH+EXZHMWoK4chTBtRJc
0zNYVYPBKMt/vznuCifwNdt+fcub0z2s2+AUfBTsh7XkuM3y2wKrgeaM3NZDmJToYe946h/ULJB/
zFgVXCEWk3zJbuhgRWD1Xq0cxNYPT6GQsWL35S11qBZZqvWTpKh3LNVPP+KwNdFPWK72zXZjYCZx
E8QAFpcyEr80cfB4wNiwaMcs13B4/8MQIhvRBdRcbociLE/+4Ypc4DII8eTIRpdyCQrRMJfndk+A
p2gs7Quq3xmHZZcqF9h3kMuQ94333vl9leg8k25CMXZTE5Fny8YvMzvWglZqRmkaxW1XPaBlHlNZ
tCZnpBIgkNuj48I4qMcUn3kmsrz0WZUiAwuHglaQUMh0E+diToV78FjHMC4hFUXKZOr9DSxe3vo6
19cL5onQSSDGAJ2Qn8UQFc8JGFIs/wM5Lf3nfOGr0ZEQxbLUcJxesAdjCrP0H3OFt8l53+X6mOqr
jKgJPs/rnm1+qUs1iTVGxUMbtMXfCV7Yt80T77Sgw4uMdGvDOaasdYFfPevnf/3y2SQURVF1RqUi
0tynxqkfs/LdmdaPWEUbEFdf7U+liEdubVQvTqBsP9izgeNEuRuPBS7MGyOFkE169ZYvYUFuUnrr
aJDk54mM3+A2xv3rAJImtZRdR1Gi9VX6ydmJGlbHHazX/Bw8/i0afY+pXT5iTrMmeHqbpNVPM+t0
bWyMngcJu5J37Bw1Mw7CTiSIfMyVdLQmey9wWw5BOn6O2HHB78DoVOshLqRhHZG5rQ+6dK8BvHRc
eeeUQ7MW04MAh7SBwEa1/xMc0dh75rgz90w9zQGEF6hBrzeKdDQKYBFxw5Kr7siqGpgeFNxj4CZg
YGx7aVEpLutjfLYfjBUYatqWLLLLTe9oghU/vB3gBJlmEafxtQPP0YiGq7N3j9cXKVRD1khCGScS
cqIC/WHcGkkHq6KqJpF0i0bT/HJCV+XDT29fVbn4m7akmIMJuO/TIYgq7PJQSBQAoBvr3FjEsvFd
xTJnv3qp1jxJaFYt0n1FscRQ6Plg9wHp5l3VXUBQzAi1ajSaF5AUEpgqLYUXcqGR2LIJ3lYdoKiy
OvdfnLsSPYZWn8o5Box+dmMB3HkpQpMYA0jP+5Jz8wwqaILHrzUXnKaMykX6glevX3Dndbxx25ti
c3rEsObHCFv1J2vn6jchfLmEAHaBfDOjTKIPfmVYDXf3Vh8OZP8ypLtboCF0GXIbReELv/r5pNaC
l+D+o+BEK8nf/3LkTpG8gdoSXwgmNhmGmQHTBmKa1fx9hUy9bXp2tBmOGOWGFh853iwoVkwx8AX3
XnCww8EF20PToGpVmGoVbQwrvYOqfDjaPCHxKlEmHWiPYY1nMKcQKPvivStu8QkiI7F15Nz6A0+3
aaXyPVC4OXjy1gBdRUEQbc9o/1vz95iFRdKz48WEIh0iOFOxaxlYZolCqMe3mhFUgJAFjZBhmNAe
Z/r2cj6QzhgI4IYyqKymdMwbm6OQR9UuDMOOMwOLPJbDlN/nier76diNkGEImtzZn+emNTl4lcOR
OfstpS96bf5umHNvAZEFoCGfw1Y/Aqll6asjrmtqCam9EgzOtYqQVhLlPdSrFfI2qnB3Qf6DdUZK
fW5WP5Xwnl/SzWghQRDrTJgZfNg0Ux8ebkfTn275YHoHDaAWmLRPNF6HtbPo89DjSTpg+9Cf2Kbt
bCeeDD8nk+LKz0QGSvUeektZzsUBlwXswtTjqBh7KWXPEgra6A4tlRd6zQsUyvJdMd6gKWSN5m/5
2U7JsMa53VJexAlA4sJXxp26oVhL1HtgD2rxhJRU9B/XRNQSo7PsL7Le9sPM8FNMcGV2gTlcf5Uc
RFDcGumz2X5Sizu6CoIMJNsKZlZFNxo9ap0ZFAiJwzbt7gBK7eMihIomfivyqhlPMnsvSqkz8AC1
QDm+M3RRKcp3qb1NOj2SS6e93RbiuBDrwhH/Hns47srNMI64CIaB41dXMaSf4T/sTejNQa9EXAy6
plLfjMEqlT/EFxe6wVC7p0boiZ9Hd7h8CHhT3h1p60P2bxMu1oyqTYnGu98/3puo1h57Bmo2XiBL
U6hhcdL5ZPWysxRAGeHFZkGEfiSOLd+Twtty2NQmhZF42B1btCUs4TF+EfWCvdJQvGseT4emrbXU
06oXl3xicO/1abq7tgFBWPSJi4GGLbdfwfPmeI3O7FeYk/4XM41OUAuw1sSigOpIB5FHjXYXe4Fw
J4Yv21KgY8w3mwACace25vM+3Vfg2TTY895TtXEpVtKwdi+duc4yqJYQkNWRTjyOQVrC5YTXnvqz
8pYlgf4s+WDlq/pXF2yuz8dMcPPYfCFojVuu4iOVZtGYCr29A8ZWPiFALF1SQx9xfi3uHcUJdCME
aWiBiAC9sfto8il3Pb9lfCYB2uc5JfJHLLqJaWapI8jA2HdGLiHPG0fzKVf2sJpHN/0pR/NM8EnK
TcJopKNiKDe1v+YUd8QZd/DYbgsW/fklzehwzSfApw20TQRTkAJlHn4Njj8oMrskA+Ut2NwuqJEv
Emf9zU+ZaFgtSpFIiA/SNUE6or3xJ4k1XNMo+cZ1KFsPpASi9qI2Kh9dfFygOHI877E0IUeDYJPU
uIysuLAsBp59Hp1pV2YnyGWII2syFlsGmFt31bycKcFOLoMi21/iNAuLlAkLnJVBNwRhj4wec3x0
10ymaN72n4T5fBloH3i6MURcwJIFekZ0bRHsy6yef2aWogAqTmpo9SDKAcuM/LDkL5YayUNsKO+Q
Dmo2Bpks21g2z1d8fUfxjhhgH65Fo5dT/GddlfIW/MR2K5g7vxsY3UDuh3zoBIpuMV+upnMMsDlp
cLMJ/WK7TWY7zgxpxLNk0CYff9n908JTTEia6/ivJXvQiA/lt5+MiQ8AMKTnXJdY2fQ/3+9AcJ/L
q+SCyhBjmIgjSHfvViLNQrbEabSkGT5cfpEgwDlMWFyvRgCaJap3d19tUHJjjpiNv6QOjfSi7B4Z
eQd41SPoI1VtVaciXr3qSR3hh6h3APQ7KP40M7IvwFjearJEeAFLdhXIOxQMcXTfdP6GkPDJSfYe
vB4gT26ajJOVc+eZe/RzP3ewiVya8EFKku8CNIYCgUQofpg+5Zq2Nocc+pd6mW8cw+To7IPRC6TY
stH+2OqflMyZ/8iEg3eDj6uFSeZ3Lbw0qEL1fp7V8RazKlQZQBT2SstxEbtbd6PW30L1+MNCZyFn
KKdGmEnBRLYMtdIkWQO8ppLuO41lIVASV9WJQa6msmQuh7kG+UnR1NyXE30V768h+k3Aa+fhGG9Y
8bMr/DFrhAcy6wHz0uJo8upaqsO9Bmk6Tz7goyb4bqlAZRdvok4PYbSFEvDwcDZg0+DnEgpBgl/F
2742huwwLlvQXPTrLGWLT8SnLsENPIsIthfpZ3cRN3n1cO04OR/nGlw8nr753TmOCS2LiO9cfhFY
ZqgRyk0y2NfcqR4PV70XlS+Qj79gpGRz3kl2uJatRc/f+iyaBv1CsptJmMllWqgUWs7cnuGGEUTG
UxTH4r5iYTm46wZgaLmpAy22mQ1TJMsufiGP/n8z3yLvFbU7S3OuzT9aaAGY2GOtmUCO7v+aIdnp
hiX+Qwk+9zmls87ws9A5hMLTaMJCWfh/gqYjhaACuhPyeINGlXt2HVRVp7l4B7lJgQFu25MKvqbr
KT7u/L6O1v9pEVSTRoPdAiBE7/bhCNEH/+58+oLkDkiYIhPrP8NWhTC1XCk6ODAUza60/TUrIz8I
FXAgly8Y8GjzEr39p4QCDzpXQ/MJzZCs348zM7FJH+5yGuojoipejibyM1ZulFKE9YEVFZ0tsWBy
rvKwLC1mIxWyGw1D2mA0/iR3UXOCdw+m0zpH1AAkBB+q6B7FEevJifYDPPy6jN91/mIfYZHQro2B
7DPGnD9e2ewr/dPbGpPuZjISUR9Tmfg3FGoCSXSU2pNhaRSznOqkw1TGr7q/heFmVfe3tSDmPIav
C9JfXQ9lhpZrhDZVux7p3mr8HNAfrbsjN4pHMloIKDahI4110uDFBs2tcT/zOU5FmdmcIJJl9kEw
82JWQZVrKYc90bHiITondVlpnfLxG0Y9EUy5C/JkxSmaW+yleGNONZktx98vuUsHFGTzSmFwpkdJ
eStH9EcKi77/j7KyGfFFmZYskqRgHJNWf2pVvesBF+COo5L2gs2pzPWeXol5lhrmr2CGXp6OZifm
/xLeIRofR2/eEhT6xT75r8cXwJiZ/9t2eWOSs6vzIXvaXLln39FYEEtTg1svtmtgyMkedsQSrZT6
drRFK/W8x7G69xAmDK7qmBaUHmBj4GY9N/+TEQ/6OEx44Cq5bd9y/NsPmKEaAjLAIEQLFicT7nC4
bDEJV0HHK243lGpNFGIhGYkG47Q/7d5T4b6e/+mAR0lKVqyVK7GEaV5xm3O5GnL1uacNfRYv+75S
72Uw6cgioWbHzNcOpvaZ68AR+q531zLPRzNvo//doDiw537GJNZALiDcHWOPsXZLSrSF2Vn4sEpL
609esqh/gwloDHKJZlDIvYXIIzEYU9IagAP43GpvxwBBXtjxI3kcK0Vry5CA2xjk5DvKJXDD/iK5
hx50b8ZNkTwIrqIwLcUkqseUn4huf6RqhimxHsYUN2IrQXR884JoN1qSTKcw40p6VJrt1wSp0Z7N
R8NXLA4jdE2qUJycuNOArVV96uCdJeSXcKSCLpJ40f+6yGrKCXGp5Qtxc67zJQTyimewIDnAQNNr
rAD2CgH8/ILcQjltLVWW4ffOoTcx4gy/wDSjQZu+yRumTDiIBRpBiEtT73CtdcKN9A2xCCr/s6Wz
wt8yCc95lQvgk3lqZx1gTUkGc9lF0YoJCNQkqPFg0J+rKCCL+I0WJ1PZCIoQ0u4mpLtfZzDQ0J4u
BOGcPj7jQ4u6kBePmltOmxDOYseHqeiWU1PXlyI68MfoFMSgNBSD08ZN3El24KA76rR65AUPf1E2
xzuNG3oYreu+/BeOt+huPfwBa6nGB7JCkFOOFOdSMGku6/UcRDbI29e9SqPxL4pgFqkVyC6QYwJg
dxDvtxL/KPMbSgvZ8woYz64/karKBUhKsyOmYDZCS+d3HZ8rfsRyJYn490zVe12ioQtvGVU5pq81
m2KaIRirRn+WdQsAR9Mwm7ODxpGrgJhv/3nYuCuAa7zTpXOkYybpO0cUw3oJ6rK6OfpEYOuyAUbY
Qtw1Kz2ajA8rxTskRb7sHunnecYHYNbEIcqvyn1zHAiAMIXbIPP2YGBK6Dkwb7LvLAuZS/XbXO0y
/+rDuW+BzMn4FpMYPScXzwvyY+hpdI30M8ED+Lx7nIzrKQBRseh968weOG0Y/Ck3ph9rC71tlZk1
uh4DtcJ6fT838DzHghpECvmYiLw/nO1kgf4/Tf7GPGBRw1K3C8rDKjYKR10P61UHMbEeGnqJyjQH
SGve9iQlUx0OnlOfmtcJ3XMwTIYDxbqSauA38oI7jzAWv1qdRAFEoL14mcokckcDyVi5Rbh1CMBk
ZrHEDOfWFZz9n3Dszs8VOCAtpwNDJONI1H0mGBCnyqCIj4ilb6tKYOTKeyoZYQAZLbNHnNGf0HTT
IBgEha9IoqT8JeHfrfnPQG/Oesg95J4m64rrjaNzjuNbyzHjhRzHmbu9pkpIFxRtT6jVYobleO9z
LdZhQao6Y2nUPg8N+JFOBeY4p/4GXUppNJ+30UWFE2m+569kcEb5EAhfeDgjKUGj+3iZQdia4UiS
Da3SqALn2FKnUjtAuG5V96E3/q7LTHSzH0FKcBhKQqkLCjdLJIm5xw0C6gt3a30fATuJnl/YbafD
lCLT7piB5JQottXrk07bApIRKDDRUurr+4SoZaqSgPEbh5Pnp/8xzSGArYZrlw7tp7INDmWXJpF5
Ffd8R3xN/NpdDU5zLpR2n2Mq2rDJ8jbBxwgb/WDncZt58PI0GECJROb0HXM8RX6OuVf5m+dBv700
iBG3dotE7JJ3n8igog60V6YVZRkYDT2aKUlAjCH0VVaTOPZzsI/Jv5ynT98XMTIvuDYwE+WLI21+
2k+RqOhpLRSmb8VS7j/yF8qbDCjOl+zr16iA0Anb0V9wkcLCusmYYRmi05OjWfTMdr324jJl9Faq
d7nS+xI73J7bBvyg18su3/xksEsylih+YcW3pFwFgux73dkOHWocjpYHqbLDyJLc0IiN5e/1lUwu
AcNfAJ0m0nvJtxVjhsiB9MSDMn2lARFx9GS3JIz6ixC9eQo/hE/B6nIEFG1AAW4/T0u4hcHbki1X
n5SHjjvPxclM8LpuLI2D4MULAoECKZXDoWCIGfB9yetliuJDYJIiuQWcxePkH+T9tZjuQVZKyFdy
1VcIhYQhSn7y7kVJ8jLNfdqtDTLG8BWoExPuGCZucuB7BgVPmwDcL+kWCSAGOD69I7AgECW6xNam
I0bqaxJx7x9GDXEdW34P8S3QyJeG5GtjA8tWwyc/iVd+C4xm7n/5wXEKwLlse8UkTFGOyDYrhKyD
MVBNGbtCTsdS2u7qGnKDIamVjTQ9PwyDNLJYUh2tByjT/czub73I49uoZlCOT2DoO8ojiDaqRwjd
ZxAcgnngX/XWHC3ybVV+e27Xv8mp7GWVxifz1dlm2eb3C0xkrvH62kkiqmyAWnsu1qewXsJPy3EJ
qyPBYp3U4hkmfzbvFyuv896q+tbtXhYrmZPYqLQAOJvdSisx7eUGOyHwg3n6erqo6pcKeiURq7sM
B/Q70hbt/+vHM5rEF9TswnjZiaHHa0nYYVYKHjAZUPPQ8VG2SVY2EziVinos+RxNZZSbjzCZDExZ
dG7rIqs8AgLwexFx8uGtxPaBTOxJbQwV0b22mYIHoVup+jYWbi+SHcd5Bo33MD/jlu8LwP+7Fv9C
rLXrX7b0Pzf+TtG35vTw61zosm2IDP25IdjYJoHWVw97bYk7ANZrrkx5oN+JEyDbGoG8EqPJ3JOL
Le7SIevX7YUtIhDFFUbNaHbA6yZIIOaXXvafQeEhLsmG/t20KxGTHzc+3XAtJYz6PxDPJkAaVVMT
WuzwehewblFMo0x2gsn22CpUy/b8RdTQjRY7leAZTlVZZXXPU5CWy+3gxNLKg4M5mRmBVZvxQA9S
YE57sb0jYtD2xGyDWv9xy+vKasW8mpzhRk4bzewho/2SgGdYxUrFidX8u5HYPhKXykJ+zKf8AHq1
Qvcqy5ZWZglPyLXynGszEXYU3i94kGmtMLaEvjid/hUn5G9qyoj5XXyKyeNsjhIBYt3ig1+RtmZZ
kmR57JrlQKwdNxybRTXa2SC1aVTY2njlula1BbM5ZfAm1zvvznFmdYsYgXSdfryJH2jJxz3Nxt8J
Df4buSKur1cJ5P/4fj7my9BtFk4ht+Ct7SUb6nNkoAxZcgmDpy4Z6TC4tBSnKJyzsc8qHkK3S9y5
wPi6X3iZpZ61KpNW3urAgawJFpt2LT8W23MmuD++Wa3A0Z2UQM54ohwNnKmRg0VSdPYzgSuSye0t
5X6IUSEvZUGyfhWcK//jW6lPw45BfIix7g8+aJHy63hnRJhUmMBc7KSHg0iXgd/OwVF4moMAB7Vx
SpEX8TfgDS4BWrbTtxdDZNeEnpFwts4++Ewyu3F0lRBoxUmY2YCVvIEfr6YiH5MmbjYrehJKXX79
yDC7gFViiZ0r/Ey7RtLWpE6uFGcJ2DyLtrjIlDmIFaGgSOeTMWBFSjaSAfQ5GnLeTonv/U7mCb4Q
oj24K3YWAC96LIJDmoJd9lyiz4ccbcdCjiOKx8Jw4vTUryiN4NEFM+neZ8CPMcQIut1PzcdcNU0q
1htCezv+WRSPkSkV1UxEZlyPf9duGg/j8l/owrpsQ2I5Zrm7JFRhWAF64IRGExWhVEcoefAfiGRz
cqgQIAVeBxxnCFFvLHt2sksLHWYWMYKZ/prf4x6AeR0bBYx93m1wIE4PpQCMf8w4w/9u3vIJv9Jz
65lRMoKezDq+v0YYrCF8MIRQvP5DxOv02AB80ADKRGiJTtSwAaNiRe8VAa6vAXkT5sntn6n0kbhk
r5ct1mCCYYnyDfpGFbImoeeXG57YRSewdHfG0AUWVRYlem3BWiSSBqjqcI61oW5oa5M0w+YhQ2iz
QU0dqGTZKPE59Zaxh8aJrr1CYa3mKwKbPODY3Lp3lvqWEnDwR/1Grp2Xjp77LpkLD/+uPyp7kFnJ
AyFF/nn+ZpDFSU5+fQVXRfdCOxTPpLC9372Ccz9wrPVptU/wR9hMMZEiEs2EOeeY80Xx94tvxzlM
dw0FyjS5nEeWTvP/40VDRmJjWILpDDDH64lfbKZYrqzb2XxyfKStJeQ3Xq4UlZvUFECWpC8jXHOK
6AbutPNmu9ILu+/3PAILfFYowIiMKR/ojINI96NFyaCYq1N1koJzbhGxcMsux1qdSnWFPuhapyIf
9tD4keVlNmKmGJ/DB9/VzfPheROsjsf1nNnLqGy+BsvkddqJ+0HP54Xwb6N5Pt752x4haM0m028k
B3G6ANyrpJdV8+VgsvFW0ywikiWu/AnwZkLlSV2aeyHiDgibLQMTtQVqImkY5Ghjreot9tQjfo9q
FqS8O08cutehLjN3zeedEDn5razYVBL++ljCOyLvsSungi9yxRgfFCkiXaqWqD5/hLQGfawBbKNQ
DmqwZztRMm/zpLKXwmNJZ1A+IOvAnS/joAlJxvusfrdTx8FUovUnMP9guTHFXHOeu1H2YuHsvU6K
OvUQSe6P2YEaBubHSCu8MSE46oRP3vLfJOcQfq8RWuh5Xos6Yv53Ya0k4qcFjzcpwXp918Fcvoy7
NNGA5K+ZM13BuINuXiHdYit3bUVTrFqnO2ZzPGnvbDKWEZg5W2glBHFu9FeE5SjA2dmFo86gFM+G
6CPBZ6sPe5XkvvDfIwlvjInyQ1yjqTjjdcaI/ohkjCQMt5vIqHCyxqyhLHLoV6iZw9/os3P22MCs
AHIJjPqPPf6ylmD/tWnBPQpUa1N5CPg6WQ/UboBhfUbhlbQhMLCgmFSxS06t1/2V4Mv8H+k8S1uq
MwKTUoY43+n/m1w/Z5yIQanOfVVPxsFpOG+J+3Vb6KbVgaxVOxipIeU7v4wVQke0UfIKy7/dREsT
knUEVKf0Q2un5eiiH+EGqqRqd5rfXPa6RkVj2ALbEzekGHogtN9b7Ak3rTSO25Tjs1DYjGwJw0qs
AaY6wmQXVMRyOfwgV13DhGyCI89jomFx2nxjhMfQ3llxqpu+jRpfWzdeLx1j++pswkJ2cTofy2eO
BHbAofuhylv6ABUybXS7ENxYW67+oNSYC7eBJCE2lGAWNHZF/HT1amnrF5ASmfVhXxs9jyNY3OQz
EITZSM+lPa3S+bYwijD2fs6MGPrLYFHzpGLYX38K7S3XTRyyZI7bpGibIiQV/stgyxbAUcf19Ib1
giS/+FOTidtqWciBhNnwh6httDJsT7Hrj/NyQwBerWfqHGLNMmMUNrSFenO3/KNJ4+i18nP4tref
5ihk6fIyzUpAtIYJwYjn5av658Jc6WB0KX731yUpvxDA38BW4nDawgk8EBwgSHhjYHDcis8xHODY
5zpqxjQ/kGa1Iv0dhsA4FemCUNoWXkCNw8oBrvCjzpZRlCR2eNKUYb788BPrlOuVfKOWZuwKvrLJ
MurFIy+KTLbi6iQBsIRQKOou2Jk+ZHZEaORGq2zrvJoxV28pdoFK57Kp+Av2oy5Oirdlij3BirHD
oM7M051/2h0HAlWVRWdppxI7hW7crm5kP7lfXHMz3co3Heb2YcqctQ+bjQ93iAP8AdvIh/7Ch1Qk
2dgCHwSzVBRrxzXjylvPNP6Vjae768TKdnyHDOjx74CRf+0gCteYG9OHwngb9+2xog4ZlzokQjRJ
espkfXbrgWNBoVpOVgyM97L31ZBu/YS1T1qt7A3bKwrlMSrpW3X2WPVPqxP1Je9G7dbsAN/CRF2B
XKYP8fee32dMqi4GXuHLsCsSBu4ZWwN8OM7wCB1Rfx9Pq7nyLDaRaKMsfKNlSJtUvNR+PfC61okT
Md0CRImeA6G5fdBgwSQIq64Pz+wPwlA1MigPoKzNVy3a3AyFonrOSfvCPJVsVsq9rwJ4h50gZwFE
XDlXFziNnN+gVm91jYLOarQTRSEGNHuEhU7KQjF1kJjvaeeE8S0sG+WgDzMc9mST5WljJBYTQQOC
cTULV200jfRuK8WfOllDNB1+S5duM8kTo7a+zpcqobgfv49izjIryFCWHThrHxHLk52CIB7VW3jA
+m6p5/SfVO5qI/mxEe/PY5fXsXvMebWI9nk36+G1VRA8akKaUpanRotSONDcllycT3w5QBicypFC
z97BS4IdoPKSDtS39qJ8Ch09+xqn1X4tNFhbMg4XgBT+uvHHDaIS9tzolP5/YH2gAjb9NDwNzfee
rOjh9J8xBpmSZppDPMPAA+wVEE6hUxnU2Eo6EFmSEOULZv08f09qHRZWH/VqvPewSDzvfUa3dF1Y
4A0BGzZIdGrktYNovZqb9EZbETZSyaqeyqV8c1xZZc0e+Ig2X51Mod7ceH5UB+tqY3ig6tWctdkA
elKfpDqCHd/QWQThvMc0DTX+G7Xr6OHenuYBifofQ4pu5yRrgFuV/dS3P7DnSY0gA2k1Ko08uR+u
TR5ZoupaHHMDVLTICjG2fGkvNvA65GY7H2R0cKyMSZcGc+HcLYXUusTQKFMyre4xHo0qcro5h/JA
4YUId8AhJcYO1qsijtYBeicoS1OkuDM0GMm/53MEdX1TPo0kIE3kGQi8UYNL2qeMU3RzfrAlEVUE
MHW21O4k9Rh1c5BJmWmfSoeCcFHYcxnOmKn+/ao7qnpchmAccYHuhBPR2p6Ke348F9ufCS2XWiH/
jehdwc/Lr6KoYKYC5Dplpng/Zi5iWmviQhK0lf+AmB1dmJbUcvMvnf038/hNrkM+FPY8IzFbSR29
kW7no7FNZSEI/g8ejQJQeXTkmJ+jX81qg2NW3jxs5XpD5YrpqDtqi+7KV87Z6UUyffS/pQ9SlccV
QIcOo/aI2k8rdsgBTqB4Twa3oiVwWnXADE/4cNeNm2DmwEPvrrCjeFyC19c3+ksgt9qaj/gYgAzC
UdQFkDl5bJEHmLEIJzqogHLwHODOoZ3YKOxfiIomsF92UY5IJNpahFPB3Tftm/LnVfTYAiK2wo/k
IrVqDr9opzmZbiDCMnxyKuMRjZw0ZvfBi1tvSNZu7QFFujnTrk5UKkKoQhvBvGozJcpNnxR4ndxi
3j2CJ0MU6fX8LavWiRXRhKXLHHwLTCqCvZWNUdFFXXsJiwvZlj4vNYreQxjOQyGQa6MVzfD/RpzX
zyrUio8ukeH0fNluAYo+oJJCIPZfkB9vy7MLX1V4xsi+aYpxgI4nNcZnF1v9K2T1LYcS9MZsKkjG
Oc8YEKvZ7LeSzbYOinehNahbTJ+bxVbVQ1Ebmu3gJ00EMJH7tvBuhEiQiDSPDntHkHR1IR7SY/E/
9y9HWkcTWEmLBOBJ5bMmQ8J4MWTr6vBpzXoFo/28jUqgsisZAlpLC1x7TT0Rvhm9l4P3As+7uGcL
hJgGT3J55/5sYcljCIWCwino7T29DfJAf9I+SZhQX8kt0a84GvwdSV92W1ArNeivJSaxQWpqEcYP
x5q9y3ca32rugjBFiXvbl7eK9vklg32+Amsu6E94/olenSqVwp8he9IBGYmk0LxjN4aVLoouvbWN
Vgi2O2vNcVQimnlbJnhjtPVzvNolQYNQIvarnTXR423wIJYS1QV0V8Pidczbymydy4xwCKKL3Pak
7SA1rg8DS3Z9IA0yTdd8DdEk2cLNx8tiIZw4LMaGizkoP6yNR+4drywLcqzyKkpAPzrhIBbHDkkM
vTJZRhewAi/kntU8KcMZrzqA+3xpoB0jq64iNEmDq9VQF8cJPacIxoQ/5ZJUHimYAZ5sNauRAyzx
wMPJ3VLBbZ1kMiPaIjHV08/lHZ1yYWn6ZxUx08VRPpC+oGLfu/6kBNkAJ2pgR2AQzjWB9CRdvTbb
NMSdv8IufNa+e9aSztuDALyR0P5p5DDu1jLN3uKcucyTqqjAouaXPt4U0PM+n+dGFuCyso3f6Btu
+UokzqDXwmicQkaRN0Uuj8ednCkqISrwrUOfQIQ3XqL47hF/Up0isL/6c1OEK3YuHRizRzB6zxFa
ezLbiy1q3F3EikGEcraQcW/dkFagsq7KQKgePPXAmtUKoL/1eAoED6QvYF13NXLtNj5d8zWpxLkH
ZW5q5T/Eh8A+n961BCfXBNTd3pA3jJ2rZKDAPZqBV9NN3U1CTW0eOdMc9w02+sna4XYP4kYAoD3/
mMCdAodWcCvSUXgy/N+c1eUVWh69UvRdTrWz7Vee4gfGvKbiXOfD6PU94elqgcNE80gr3j7zvhKu
ZwmsS6BgO0z+Mif41A+Y+36b6XxrDsqr8GnqKgo5LqMzXLtx+KLWI3/R9Qs1PblvhGJtCrPF3sHl
pqO0ZqZYHcLqBbltfl7t6vgb6nNPhQCmQoCMxxdE5w7Jo0gW0aOvmNQXhqCLPTO9GS+iRWkjHCHy
uX26SSF4IIttJZcwxtl/ddJIv2ExJQ2S2xKmbQOWFkyJ+wxokRsFAGmyMBtlWAeZ8NHel7gE3KXg
gXfBswOF03Pyara5WWekTRPK0MTaRiWqHkmzPM61+LKCSz+SILVPLXIBTo6UEY8EMw8PJFuLLkiv
NkFfY/IQvFXWs0hul1yUSEmRW6KT38kBBgLbOP2BAkmq7FI9C4tMHdd5lqv+MawfF76Y7gzYf1AT
HhQWe6OnQbqxRjA3WiRSmEOmGPd7BvilDqVsVQHOUcoSrZ7ckQCi/MBJc0QHgJOu4wvSwfnNKZ3V
/XrWs/h/ZgWw4ieeIZAHwAaYvlKHx+3BbXQeNwFIyylVKy0dteZqGrk8NHPOOB1Kojsl7Yha42Xn
Gjklvz7RWujc7nsGuEpf2+nl45bWW1NtoE2vvaIXuMNjfWSD9XxbiAci/KpVZJ99g2KZ74fYWfmn
zX5h/7H5ezEjSR072O3GTyv6yWJRFmwI9dBptGOY/sVJQqA/M8zJaGJ5/+fzVIV8XecRO91018Vo
ve1uoy/kwVYrb4cq6a018XzVVjSZjcAMRs5p/kLlX/2Z40FQocBkGnvKHWNQOy/xWFrNNJWSaB92
sgVt4EXYWzs1zveQKT98ldQG+4V/GL0Bg5Kns/Oj4v7ivuTVaG09e+leRgs/lsQiuIlDOboABk9u
qOmGsgNJEdopaN7e+EAQDi1f2Y1DwSEOEcyBt787eezkqSX0V4n0Y49ia6q/ovxeKMjYtOOW+Bx+
jQk22FI/Y12adk0iss9nZog8Q30YceoWddYbWb67b5mQF1W7JPaq0mY1EQAWKFLjT4yQ2wl89GyF
OEzjpQ6ITnTuZEMFZlAAoLurYYrQSD9ZAzSZTrtYkRe1IvSPC9dP/aqV+xyBpGfEfLT0+t8cpZTl
tXQmwlTW2fYjZsEU0KOQN9LfIQgRL/pwmWV4hQ3FPZFwJ8MYveKc3Vh7UrFX2OtuRGx8E5ujS2W6
1DudcwAyY0tP3G06vvEaj5D9sBnpZOY+OYh3mtVueHZxGLsPkEOq52NkzuhYURGJcbHTSe823m10
LLjpB4AK3k+XK8PyuTPxNCp5aZ+9utQHCs+3Nk1lZ3SYTA9Obl6TETmiQomb6sZnn0NCBdvoL2jW
3+TebbuzFMKReL4hZVp9RpamdyiIyEvD0BQQFPV26o4Vl9R6eEe0XF9g0cJB8QWKY7qO9w36YFue
TjIzGrLUyV4hzm7Tq6thBRWZKhvXQxChVBMcjg7Ozhi+s16LcId5gXVnBFcL3xUOJR2Kdk+USZcS
vDSXF81EOomcXwLp/0GOrZCiSWmtXU1RgtPjJvvW/DhsP7xKd75TdxHbldZ2MKhxltmU/kwqe/yT
WD7/4oLN+bFSkRm120U1AP8gTiUhy+mN/PUPoQYF7lv0ynImvpQ/8IIzMBG5RSPNxXas11QAkmrB
GKNUqaiUiAEMY/7QnaVVBjbZx2VkylsrSjnKbbssEIDygQqzXzQeqidCiltYVYIRWRS6XKVhm/vG
adyCqcTVvB89bOERyrlT0mO/LoZ3WtOnLZRu1CToDsS4GOibgruOyqVZR4+Fns5EICYeRBOH6K3e
n7CMlc/pxAOEb0qPUlzhy1K4lDg1tj4Ir0OPYdMDCxgiQ0N5ZMTyVgjxRyubJexq7NVfGbXUOY6W
JgFnPSx1OMsXdCm4pg4D0FOgLO0v0Q1X10gGUu3FPkDCQZwApfID12ETcghKJcSswrAgIgyMxmM8
LOmZW8p43/82dphNewRpJVypTaChHlpxj1fA2OSjKZgaLeJFmvC5JljC+cGN6IJxTCg8Itm8CrRh
iXpiLIvtX/na7Z3SN6De6/p3QjUys8xSsej/1xSQPHjlQe1Fvv1op4WWGwCTBuwvxSgm5y7AKd9b
27P7iLnstiljxNeYDi+2vIGOGUJBmN4cmFSLKSGnuA/z96FZx67YC3+Iuxz+nmjKHhiuol6IBk4E
P+TwITz8f5tcpNq/Edt+Q8YVRQdn2Hbv14mKL0PdvSOuz2b0tPjWJU2AF1WaBDFQs9KlSa960nCz
Bk6OboXMYEGpzMLX65rn6F8n1u+pFMv9kofJ0g5xjf2+4HKxWF2YBQna89NVsaydOpmMVM9nT6uB
dUyzD30qCkKuQ82sc0FY8zFlG9ZHBrYYeVR863zMARKrMG5c8kjPyqBebXymUAdFRFur1e9eIpyT
oNabzuLM9xdjquxyerEendTFjRxwWQfqZvMQxv8HbAN71LgQ7x3L7ltwF6AdNch66s/ASS/ZRwZC
PWDD3Y8P7L9AF8dY3xBHYdnMqtXSP7i5/orU4ZetTsE7Byp17Lh4v4L1zQUemGvZpiJP0Tt+W8S5
KD8Yo8/oLcZiMFSPsqCZGxU8uEuh/tUh1WmdXH6vUvt34UuYDte1BusIkYAWXwhHn4m8EJqOEnA+
AHckC8KC4Yz5ec920P8ecoGETthRKFZZPb2+mNl8FGRrzlzUESoIMiiSP/8ApymYB7Gmh9H1VLKY
nMgWbFLua4lxlzvszIxuO585hjqhhiT6eHhOw2f+GWAatGmOxDUubIELclTblHVMdlFaOAfUma2P
1qteOz95gjQtnhH76s38d2uxJV7Xj8Yzk2jP1XUc0rQu4fTTAWES+i7IAEZnn8voiPFsaGyUVmSr
RXWVns/oi9EiLk6NPTtJ1ZPwkU7Z6OAwQoSII8/zG9Smg1oqZtgLTNQtjXc3HiVH2Tk02MEE3oCw
9hVT4mnG9ExlWf93zYKCADP7WqqMb/6xYyOrPojEUG3ZYZ9eheypvwPVHFHGzl3sg3dvI6O24UzP
VUe+2acpDrWE7uq7ATVdA9hcX9Or8e0o3/YM4IN9NSK0EnaxkhXOk0nhWw08+oJtj9nd0Tuk7f7v
3KkeU0dL1jd/3OEYoeVlCPkJWwM6y39sivjILKTZ9szJzaD4Ih1Js0D8SyJ0x+QkgRYV4PLr8Zwl
kGYEz/qQt7ZJlGWY8XTn2AWZho57r7qhtgQnQ8fhu1xLPs2CK0NcTPyXArGVPSWR514KuPCjou5K
qk6leyqjj6DKyxpbLc2BP5eherhfFP9xzfmZB5Zn3cYUhXGpQ0n2o3k3rd0m4kIr8K7QMLikB8lw
4tNRc/D6e6wykmw9eUA2agEBLTpUcv06R+VfSzGSgdCrCf6oKC/yXapCnxrWR3yAlabDmxUyM7Ph
BT3NdRpvH7ta//ueREyBDiFvUN36gFu2aYPj9IhlSnYk7201F28jflvFrwiXTGK9BSRzeMSTp83O
Zf7nbveN+rZuA6ai565wbaN8gzU8404nbVG4iz4Y1nbEaAifvK9E1/ogkUrvLdq2jTwpWLOX77Se
hcs6pzjF+iwFVU7xVqe7Ervo6alknQ1JlhRa4ERQapVkEn242r/w4/TNkR2h/c4114Dz03XbgLDT
EcGkJF/+Lk0wFpSP6QCp2JvIfv8MIJOMr/wuJv2ZceTU9MVgg2CmC4YcP6rRtZTbNlKXhN1cnM6/
Uw8pJ5f654owDnMDejPDbxBjYWnsTeb1KppDAzHHXyhX4sbAVTCdU49SePqp15Rq+2TmFhyGNZlC
ZZ7KF3YvxN95VBMUpCSo9Dq7hCn35RA5rFK3SrMp6QGKd0PEcy1eUOb7f9ZFbnpQt4Wk8s/arY3X
/Aj+Uvyj0aKmzJiSR4Mk5FaoitBHZECcNfAf/quI6pJVSOkz41p2JVWsFG08M8IG8uriqj/QpiH9
ds7OesUNMRRLmj+3okclsTMtNivwJaow205ZcemR39uODenn/ztdlJpz8cbiJXz0Oe1cuFkyjefr
HQoJoABrUq5newAG/BjvD6q0LiueCrCo2pkEAJKFkqscZ/4l2qw/VQeTkv9SGFkJ2nhK+ve4AFpf
Z30mhlg9KNiN57RSy09jkRcvZLiz5EgcZKemjOmMQKcXZiVdd8zY+/yDOTTHOFW3nQZiC8hDJHj/
gH9Xyo4emFUcpEkCm9np/x9etiThaGb0n+epZwBrDLAQ0gw4BLPi/XdsO1unAzoIioOlFTTBRawY
NuqvlFdCg8tQ16p2ktIKbKBvVHXa+RwB/VNqj0r7CgbSIoc6CfYXItcCDovWtRCqAtoUuAgrZMTh
irHrSuCHovIvcttlvM6LjvEG2Gvv52EfZXEH2LNTLJr0zbsiL1O3bkp3ZzPSnDGDtqwBtxNPi7yY
l40yo/YSw0/1Kr9eUZkDFwqVlK2slkBwDjXz1LjS5e4BTnPnpZNA+fxgbP8RaPUVy+yDbrYJiQeB
DhW17PTcaHOWmkTCEBj5oYO4C+6wTBy6SMb46fC0YAM78c6RAMWnSsGbAfcPYgUVMdsEQaCoh13L
gRbDQoZRHG8m6TEye1SV+2oTqQOb/yNSLJPkEZz8XinWn00Y+6cLt0H2q3O4DdL+97aodti+csSq
UFh2BRnBf+MgfR0aQUkaC6FriXCUt00mbnJiCgnkUKi7/JEDswLmFokpfOaB5VjG4UAVi7hobZaT
LDQNnti0znb437dk0DplSkopkRkcXVMUwqLFKa+xjwcN7n5fpaT7M5cpSjsZK+y4MG/btsCEK3Mw
zBmNBVolUoaanQGeDxuIjKK2kUCHbon3cgz35LLgqmaBaPYf21c2ziqO5XQC5JCRvdWN4JxWlF+Q
5j7eavazv9kHgz2RJN9DhJaDNq7A8fE9rZ6Q3+vB1YyPJntIIfyXTBfdMixnTY0yM/KFpiPd5myD
A7inMgFesr2/ccPV6JsE8z86hmGdqT2gLy1Ib9QMltU9zVwf3V0WPnZ2e7b08tw5zjWZ+UAspnkj
Ddg2RGlbtprey19poq7ORLMf42thftcKO5wXXlUzFfHykTZbeIYCJxCX17IOGZ38Jcf0fTa4ry22
JcoE63dA756QsVlvqlT+D5ZzAhYGATaH3YLsLzkOX3GzBcxohFEBajbiMwEU21ThgJwuyZxJRiaK
uMJlXaHjooQysqm3mqGwC38ZQtoRenBbISb3cRzB4PoY5lLG27DkZGqOFN5hq+2MMSoZ41LgtpXa
MmDb5Vsn3+F4Z6lmrEAd2/QdB+MGkt+grz8rOJ9aEpAqCvC8rYvckZbPGDxr8ICnipcv43bXsAvq
sW/m4Penv9B8uRvHJsQzMfVXL/oIS4cvN2PvKiLoIWlegGSzG0qPGnwtQF0RkvCajJ+9gRwAyVaD
Wrtji4EUBqB0Xllq4AF/g8WYeyV3rVQhr8LdLTfunxxsDlkbnJu0y2OY4fDS6wlZUomrB7c56swx
0WfGvuTvkYA55QPIjIV37VJN0bchP6zh0Q+9z0WcbFregHnZNUggO5N76AijtcSPa4R3/U+xwkHP
qaJsR9HrxLN9J2JUGjZIM8PEvaEVhd6hVRZhlXpDRpdAgIqpvyoJkXG+eWex6D+XCUQoDW9u12Wd
XSnv/1UMifXfTXqoL144M0sF2seq+XWa5VOjf+j/39ZsgVcJ62KJ9YLLK2UgNPmIl5VbfBb/JLo5
cJbMF0pGxLG/tlHF8Xk0ZBMeydrzKS2Rh4Bx7YhqompzFa0vH9Kb9/BuUB29du88mSXzY1Xo7n6O
LOkRwNhpoMLOr8a7Qec7Z9m+tkg8VkAky87UdpgH/FpDd78Gi00/2RA4upDcNPwdrrMdhtVt1Et7
u27tqbSutOBOqTeF3DLRPdiKhYJ4YZKUtZVnDOeHJ84xuc0r3738XJtgETLUCYnpb6EqUug1HLDm
Mn7/l+xHjQhQlABsypHcfgEo8qvPP5lrvRIvogOhwceQ9lvULELjMz0oXkBzDAEjo5xBxHrR3Kt+
6vg85A5jIBXWCNDhVAcTAJ5Kr4YtfSE3V6TbzF/YRF3SR+jdpOba2N3GfmTxv/DaeYUYwMNmPjeL
FQGMb2C9EyOd/imJZzJx9GTcTuLvb9OhILV6Lp9eDEpOdiEW8/EIciih7HqHwDsBoTRntdvpWyQD
H8pA3KLjH/pMqkN7dQnNXiyJD0ft8GWaSas+6/mJS1TlmcgbH29Y37dhbq1wRdCzkJiewsucn428
nJ5+gOjmXcLJqlZJsZ5MmEXMHXwo5TFB25zQmOwCnO2TVwim05FWXQGQ/Yu21UHUebCcV7s7AhSH
Chiq5zfpWPOeh3cY69vQmsHtj+6MBsjBizNysiHBUGnE6uj33+ccBu6o2AmlkmEeJQReXN4tXwey
WbW4QOzgEzSIs2zf/MPdqQbMLoEcDG7nZJjEw7ZZ3vqzT3EycjMBArhuAd+ONYLDEhJ7jIyd82vt
P6Nclz1q3fOhN2Q/Rw4JrqzN4C4M0PEZRGL1Oe7cj1tmLjikrb4FZ/w4OBooap3oZWhBiIL8rUy8
rjkA1FYPCm2RN2RDAJ80Nowf/WyqrEHO+7bdsf82OqV8ySJig2i7kP8SsTzoRID3bCGt3i8C0Vn/
yjVUXE4I3Mz5mLM7X5rs9w/tagtJ4UA2bdK3Bzwd/atbtrOcIukrL/gLYbrM/0ZfjXQPkdPXolE7
iXlftwHgLHBK33w5FynKbpJP8M+c5ZVEhlTqZNL/a81ltSqUUtsZCGMlMWjWJwb7lwp/J140bM2T
iAGK8QnwJIINeuiPUd2pc+Zjfr3oDEbGozVd0HMCYSH1YhwxF6msm6UZDdoFdzKZaICNFAjc1YNH
h+qixBzQfEg41/bOq9Rp9MNr3Ext1k4PPi6hqWzOJuxXT4S9KV170eoJb16oZgK13SVSp5S1q7B8
hkba5M/NHADXCWEVWxUa+tJ0MI9Veq1Lkq7W1xn0ldO7SswkFwjEg380usjp670On9/JCR4uuuCJ
IQ0KeXbGcofrBUjPWrv4+8uqghD6svSIPK79izzlsO1PMM4Zqp4yptxH8zJc4BPXcudG8F80v8qv
uQj5d7+/VZce/QLO1YYP7aPNtSZryzhFN+msVWJz2QBJGP48YAcOE7ua97y9oBqdMf4ilL0On+vQ
BExjeXJkvk6GgTXMRQi8mbusiy5fFY8Dez6AqpiMZxDadncY9KbIejuK9frJ/FOv17u0KzltktLA
wCnvQMC8uruoI9sWF3QjHWOMARuGuZ9ZuxNgGV7s45sh8+uLEokqlAwmD2AZGraIy1RG9AdP5dz4
qMj1uoMCTqthfaQj7caRYKYsEFssFp/IjnMLw27g+9Wt4oP3B3dOyNqJSHZkzhMG1VsIdgFRRZcc
DzJJjsZxrxX7/e5BtyCIuEG7oqQVOYSqutqRD+EBojOR0g9q+pPEyhOOY187uLCMhXss9BAzDFh3
FfKNOem/ZxObs+5Eslks/HpPfeEFQyCdumjoElaH+oYCObyaytj4Ajey7bYIrnywQSlRBLs/Dgz8
Yt5SIV9YtYSvouHvd/HPtbVNKnQHIL8QCdh/BVLzennyMnOXerigXg2427rz49jCRrlLAltwauPn
CWgfIHP6bJGlhMvkGZKrLZotYfqNZ5uPeSS8B4LzHf9ros8NDBgi1FB+wTjYw6E0yaCq3OqhChC6
qpcWaOUMAo17X5JorkBeVJsGvLEJDznCC9LSgmAxbMc0b2+hdMfO7pOOS8kXIWYuNsVG8nfeQ44M
RixARO1VyioMrI9cwaZxZ031w5tkMq+Pt0JHrpqr/t8Lc+0TnTLu6+vbPEiaaFIKeTxEPI5Yyy+U
wuDyGrYwS9UXxFVKwsy7X3bR08O3lmZ5zz6LB0ORqKUQ8unHyTuHX/2c2MUyRM4DjQx/Z8rf500A
G8wwta7oY+bJ2lpl9XyLLVGdrDw/wE+knZjjEgDf3EZEXu2PTYl2bB8P3Ew3ilWw39IBREHmo8EU
yDADwhDHv6p9hS43q1dTHy5rifO6XRGJ3zRW++jO3/aualmjfjeCeCnKmesOBTFDYB7OcFhCQI2y
B+prd0qHGxLkdHHu4tTPh7FC2pwoEx56/4x4dw+7aIT3kn6GEHNRinS4moxYGu9ZxvABHuRoeqUd
DK03jATRkNaximXnguf3mqeM9/W+S8VsvtZZSrwgrvY+Tz99YgWGuPsRMTZxP5iXIm1D1LXxKemj
dM3j1i+du0Idp18+CirvwAzt98a++7mTCqUUm6pTIat/VjmLHZDUIFGvkPY1L24qF8OlUfFd5S+n
jChI1oGdiKnLw05Ltg589926To11nDtGH9CR5noPTRJcz9yW4wfZbOuhWWfky9IMkv5gNAcxvjr+
PmQhKADf9G1lSLZWZqimh/CW0x2rs/8hVMx16+os7iZ+5d1ZdaSIuVj9ELeQpOi20FGJ89GHTPWZ
RuvqCrJ9ENbFDrf4g2RLIGWIf0X9sIXux72+pT87Q55lmUxH5ymTBsU52kWQbAF3B+T7DhfUg+L/
pE1Qxxtqy/SoP7wJY4jeDmi/PIxxLpQx0YOrDMQz9FRUbsfbZJaPMQXkt0OIYY0P7oQb8QlXluXG
ftTJNzl/569TOk164sDn1lOosDx88xzdTk7g68gVasvcQ0l1pP+tq770N7gJ1M4uXds1W12YjKgd
jCE2Jh6StAAjBFwhAvkWCgiafpCfun3CKj4FXc98QATeAxfA34Q2LcnfQfoqvK0nQyg+jTxBpbWl
bb6J8u8oRTEu3EzXRH+zmB5SWRKSrCI8vA8EOFx4OBCP0cJmKjnN0n2RU4MkatSgM+FAYoEmNTQP
4+piYDjnnWrgJffXFLRqBJvNpFeH5V9vDGn4JX7g3bYOUfPmpvWlR37/TzokcWqQ0WtuBq1v9WRb
09R39YLFeTXDqAmhq7/IbdIw+qJrERiUnp3roO+5dzM9V+ha3LdUnfrqSRfhLPmVeTbNq4nN2xRa
JQ5mXFcNMz7MNR+AUlcK4tr2iUmm4Yvs/UKbiPUWd2GUYI+GmWhmKckO73dqvjJIR1Enm88/2vST
/q4mprDBbMqBiOOqbskJB9LDIkKIFVs4fPCBzN0buGb+9O5bCwTZFMWCDS/30o4Ww3ZGZH3hoPM/
n5nxjJ/MEoGheJixWfhB6IxWFNUzs2ZKnUZlHjlEK9658e+2Oux59L666u6DVOn4WzyIZo0nsK9O
IAgoslcs6cELcd/E2cB5mfJOV5IQgAyzay1WE+84mJWNF2SWY567bOS6YDCvO0mn4jjqDemK45sr
nWEzp8HAs/1wIwSS25R1xDJjONjFz1J09Hm1BDaMN7OI3DZSyQlyXlTljqetgKoTZy0Xrjm6bplx
VmkR2B0Pr49WWuUz01RxwcoC96WxCrZr+sp1F6ZMHTbu64m5/8KwhsZKltmHxdnauqsGOKCtp/NI
Ea7QMvITG+/5IOV4fay52Wygzcpvgsf+1v4+bxMgVFf4bhsWWpdLqXUagVYR7D+yiPgbnEALtTGw
aPSjq4awYg6CrEQfAiqLjw4dP5qVt/j3IaDuPpboH4wxCr5FOCxUCa3lEJfYCBH8ZnN6yqfHM/6/
g+PzINO/f0C/hopMCiisowR2EgHdiOENELs4LMr0EmCbMokWm9IQ2WOZt8561k8qK8g5az0yndAx
LSu9AnsbFgXQOsm8zt60wDYJeXxSp2nqjhUkrLQR+ZnlDIQt1XvuSHFpzDWctG05WvAGKZO0DMLh
jAprEqOx02RDlPsaPRcOqbkGf5L4nq5uBe5TxudoyCFbpWxETD3I4m8MomWS+VRdHhtu3DF0nnxb
0/lGCawbRdFjj0sxz8QLYvv+J2OBlZbFvTv6M6K6xdGLgiyfEEykkaZFVFZasN51M5yQNVCC5Hov
rlZesCuyTVk8FxsOCbkb5HxmJteb5KEY0S5/j4o2TxznsO8qomM/tySkxc+C2JEaiLcKlzQKHqVo
EzaxV5scQ3YjQ0/ZzYLoFCd+xABSXUCZN3fSuv4+pwiMtO5BRXmAgKbAtA/0ltnKqN6esHhcF4uM
TTJwY1qMHBPuRTwp9b1TeDlJLyApA7wzhUzC6LIaasCI502T17nxh09pzm3UbT+GQBxSavb6z/1W
AH9K86yBxfCur3pBS2ASb1C9vN0qimyM/yvHgA78uWLvS/WD788J7ttikY8jAik7CX2Uy40qcz1v
7qM3bvKPeDx93hDopLvn3PhtiUhCisKQGiU2YPbmPF7tW4s2hoMweg6TLWBMpTf8QR7le2vKYVm9
7hTRCD9X0geZhnJMYhMN19YHb6Lv1vnGJB9MOO/aSfxC8qKlQElqfLxbenVQ4+62lgxJYAoi0+JR
S+oDGhPTTc41lbVaw4DVinra0HAD7W9DExTRHFKjrAcxwxoVio/jtxMBaidwpFLWufmZ3MsCDUo2
0dfzEzf8AcW3d3wWEXBblNXOQJBZ+VtaR3NOajPfZzV9CFgn6JaSyaLR6YQjpBlq8y4FBP6Xfhj6
W/PeA9CQjq8S/27v2oAsem5KJQtgRjHFN+0Bd++QjWdH9SMlIuVCKGF9PwlsBENY0jo0xI2TfEnC
R/Oc5T8CCXv2yrRomGqja+nU0msvW9UTsFa0JJN27YIXIndUJFHyqA4KZaAAPigMsNUNEPDnEzPU
78qDOnEwOEBXN0fEMS3vjP+k1CrVNWZzW3Yen+xAfvHFOEd+eXHnnAia0D1zkX2pTXGIe9IRSVQL
SnK4mmnZ6XObKSyjVMhygz5PiBXUWsizn5fwThKuBcfbspsoQPwybK6kyEjsZtKUv6jmDrYrhsHt
jLi4kwuApBLY17Jr8ezzQiavJMtTfSFDE6nGLcX1Tpvl1Jxntd7fDeR3lltGecmIPqeZbIVLHJ24
dLuAzTtsbNzcHt2/J9m0jfHIB/gBZ0AxCmK6YkZjFJWm7rqC3y7er610TZ9Nhp4OAm1OWTrEEDw2
AQipxlRYSklIVkewDBQjSbUm30lCe3f6kkRy3/2VJktj9IMTT69+Sr5XmZ8O4YOhxhPO9aKaVj/h
iVvpQ7VZBilGaPQx2AVBasHrSXW8VZJCe+LXfGZWf+TjqkTKWQ+MGaE0Xpc66M593JeOKf6kOx2m
Ui+4UpEnVogeBvJKcuO0jotnhgE1r5yJLH8GmyUOh1AfTO4Q/aVw362h/EEltld+ViZsvvhtZTmr
uDSk9YikYIkzV77Z5ydAp92ybInAoCs743kDd78J4BXmgnbvtgOZE5rhtaypw7c7JWLvwTczjSzE
KTJ8pHYQpv/OvpfIp8VTDDLgM/asx3FIpO+Xq99pVGhZ7osPberKiBhSSQDRBDigh841xHDRMaBz
cJhnyTBRYn3xVgQYOTglndyj7Lz3oy6qUX3In1aOMSfa3w4ugVzrDNbcpyL8Y1fCXHRzGqNnuDy4
EHgvHwvaABsx7EGSD4QFgXGZAThaXaoUExCCRvOu25DR7QAnklYxeM4q4i+svxx6/kPxm90qUV/P
mSJ8ulrGCBoxHfna/hwM3RWt8thAoE1X6YDviIF9iPGopoDPyNT1fVt6DDfiXXhcWaK26PXCr3ib
cKKGNdKku/DX2/3yGeqKdZkShdSRHFOk88QmbxrczDD3m5j7Cs84wTrE21p/Lh/GdKb+Hxk7/Z6X
i1EWC/stffsmZEN2iNs9U6BEp5xI7ZZ143mI3U3PcH4SNj5ueh6rAGz5lS+P31hMIS58UBQmYePp
EVKO5eXWkkOLo893Z1An6dMxv/GKay3fybjWW5UXpwGQfKozEL/dWvcHkvcxKrDB/ssC9ICGA3xR
xtzpMm+i04bmLY0eVHjS4b8ZYgoibmTcZw6frGq5sCZXLYC05yeHx0YchpgEhXcKiweZTfpcurC/
eyDmt0ftF4VXd8UmXfujGTlMkYYw06QP+ouk8nnFY2lRHznPNcCWt3N/RoFVNPLCN7a3ty/yrp46
ft5GCmOh5J6MAYLx/ph0a/0XBF+6F1NsCoalE49lypQmXNi3htkDOyjJxeu/JorKgG28aPuN0RxY
ltoLHfezx8nscKt0K5rEgmC/Xu0wCvkxOYk7RRffzN2UqPE7LBztoOZOdnRA2RpepULde3EQvTgx
VpWkvY26DjDCC2RoSbxzTuiP6Eq8BUMYei6Cn0SiP4okTT5ThtTTjHjP2rdr7E/V5+sUYGhyOYhz
Io3GcaDO5rVsP8lvI6MnaTkfuONmMgvWM4iq2FbaUFWb93Nw65Yh/nskof+tBBNBM6tRrqXdW3Bt
zVMNs4X+L3YXxRXuPgysjO64A82dFMv2x5KVjKe4TxRDFuLHrDMWzX4u8SKCAPxmy1TJNV9M4k/E
8LrgYZsBRasL8ss9YgDxILOVP0KMDQydd7Sdhv2QZ1iAsEgDlBij10/4LBQQWPGbsmxH5nslBWzw
6sWBRAUu4004SoJ27wTF6BdfC2p16DPd8D2tkZMV/Qn0UZ63eD4NXBe5FiI1vbWgb8yO6gApObFJ
kzEV1BB2dxHUmJ4pQ5PlC7c+3EsEIfCO4gw3lIXwMuAv1/9xmt8C4aV1J8N2Pa32a4JLakdVMc1w
7OUgpB5ZwIVHMNP2mUGoHrKNyw1CuU5wLTs35O5OmDjlvWodDF79UCGdIq+o+1jaN8iY0mEK+mps
I8/BFy9GbnxPFDvKmSI73yA6Oy9dAff+YBVVONEQ4tQaks8fkxYA4ceKu+j/NGBCPdo13n9d0SY7
BPKx78Xf2Yt6K9TQlTxnjKBObVnW0XkKTS83wHrbbYilEPvINtVTJlDxnEAVAdVNMKW9CYHHYfe5
ZG1vfJSi09dX4eeEKDBv4O6kyEpMfvzYO7j0OPQ87uCO5XquOkse/6YzvG6KKiXfPdlbQ9ktdLZd
RN2/s7PtALN5YTnF5mLYAkbCYPKuX8xK9Oeve9Zb86+LQO9PcCXmQgP7lsFdC8kThP/0uR+bw8Ku
3UJ1v9jVGj/pQIyLP8xjzSLQdINiyZZrswsCZEoPcvH90PIM1QEbxnDX01q1Bg8ivCpnUcXZBzUp
7t1c6vg62xMQ2LXxQz8dw/bN0rdWtOeZ+Tn7a0HIceXKASfADkEWz3XYd9EM0MOKxMZCPsfUvK2K
dRyHD2H9nJxsod16I2idSnDrwxxcw0+oH1B1GYQHQVJXeL1wH7jVbn/0cNZg4XMHaDTTE/BKiw6M
15gdXyKA8yMh0neXWg76Nue60lKWTMFGxkU7K1xH09W4eGwgQyitXpgh8FnzAJcJdpDJ1yL6MzWZ
1Mm6QmlbON4m9pDdP/rMmW14oiFsGVvsme2aKZ+tyTe17HpEUPFEnmy+4YO4hm7M8NSSR4hi5ouq
WLX42AeaVKPeqH2TMgzqPCza3fpa7+wb/lG96II3MpMZ4fV5qfKgvVCa7dRLgzeprS5lf2d3DIES
akGHr/UEqE2UCD5Vzq74/O39mlj1vXnV8hmTrei2OOsCJZJMN56ce8KXCx3etjiUdQUKk1Pc3Zm5
nPSi38KqDNrbiAOID3InGrvfkQp01PiFTws4BySoG/+kRD7frn03D5Thm4VS0qghCC0VAnb99oTm
LakMKBGoQcIPG3jUrqkEkNRcH4/Qb9mrn8BoO8ZJax59xtDKM6hfV2Zw/xGrTmFNZO7COf8w0SoP
2PYDZuRQWir4s9s8x88GdyJPbK3PLb2Fh8rkN7NEhNRFg9wfCED5wmcw3eI4FYJxJNmKhWiaWNcg
dqAQuINwln99HiAX2ixogg0So9KPY9UOqIRy8jk2s0YE0UgzX93DeNwK2B7GlRsrSHN0RPGNJxgJ
exno/cXZn1DjL6PXptGgZ2mNdlJhtLq0GJOs3sBw7Am5glFDGBxWx1YN8GGz4rdeQ0QBvYcOTMHN
2IOHdi7aOtczTVc0f6Z92HMhIqYfU1ZFs0SpJQYi8ZAoJZX4C+iV6QRpAHunwAyRB/0itojGXLhM
NA+7N1RprfszAKiELYvxm8aXSBR2HskfVhE4nUJ15+LpnBCuiEGMgRDr5lplDmjEvk+jknt5b8qQ
5S8c9Znyiu9czoH9kfkB8gw2jOgGGwodirnn0/GC34DK+tYWt/1U6JelOBu8hDQOLf+51x17Tsl0
qKdIS+kEhNPIaijwcI3N6q6sTBF3fcYv0imkL24szOlryTweuOngRD0a4qY5oLEYDg2MnsX3Sbu1
A4H2912/js0EzQHBUbNlVWswNzKbty7thiOYMV44wQ7m16OVkhpyqy2RgUZ51IzByb/RKrD2x1ZM
lxZtK8FltX++hfFUJ/D+LtOETKU5Milv5nuO7Md1GZvjo4hkr4o5LIQpoj/wNvB40IJam1nSQtbz
Vecb9TfVizMQV6+CUaV9+/AVLNFmLlxSRNTjY5Mnx0EatnQFGaN67WDSa6lDExR8PBv5r1mr3Kkn
LqDNubaSioiosHWLg4L3rPqt2IAz28wpr0B3wKncpnBHJcl3FM8Cvza05HTi+8ZRmUlTEauuIj/e
/fwFYazVT+aWnZrvVFImz10CT5jP+anMgiuxV8vRClSd8V8H3AYJX6O5fyfMFrYVrD/z8bLv/9Kd
daJdkYpkfP6jsG39iFfULRkQncWHvWGnpKtKWgMkbuqtV9h5lSNz43eRsWHrvWAJq9ccDs4pPM0J
tuN+2c3UiwtdZ/dG7h9hlhrmOJY6lv3lKUudo+RaS7FPN0hWCMgUCIXKyG+xqt/Ol/AuTEeun3NX
rn/+7/iExpG7jb9Dqrf1MJBVtPMnu66F3UtrYP/yKHFOUSu0gtk0euPQWN5pw3n3djwQ273phgGe
bpSmMLKBvT7m2FKWzFXN3jmZkETfpVDo7doaloQvN1uC+1nRZb3V/QXE65lL2GoWHHRBmeXr06kn
xMIz7A/DU2rlQluW+41idwsd5dkb/9kiFTo0FQqa8Cdg8BZGm/CBXO7ROutg4hlURxm/CQKUAlCf
l51Sq6lQgctA/y9JNqLjU/GjmeOiGBS5KF7bOUD68frKO+ObwIllLD2RR4IWOHfOfWiSjb6T7S2w
51cEdOOPELBhSVcNxvvzOkYtrZU99J2gVooHu2+ELCDZSniyUlhtyGy3WfYHr9+x0AIoI57N8ThO
qmNxOkram94Yr01LITtkMyQI6y2fR+94FMHPO3ulDhp8tanAtZb9bQWOBh2nc6pOP67RuS6RpBf6
sFr53ZRIdd3nXQ/j49DWhYJDDDDd++GD73rnYL/lUABbMjAlI9LyaEFtrx88phG8HbuA9r0OLGAL
yLakDCeL2lq3ENeqiiH2UN0Jw4Dle95pu73wY01gzMJhf+pAW0ZYkOGn/0bct6b1LXLVWlVSJ/bg
kJHy60C/Y9p+Io+yzDRPZAFiiuzE54WhdktZQxTQMXTWxUcrdkA4N2MF3BGcwgLAHLJfx2HIzV/3
DP9u1ShP3m7T6KZeexaVnjpSnpCeJadnf8JgxNU/7evcklUYYPIAvHa6ZE9JxoTU/P4A5pZCKdzk
2pEEDPTnHIFPYeiuuO8qjdoZizDy+T40yU61RB9F8wVxtK/kmRyTPLfWwhIUJ/oI2dgq0/TWLmMT
QzHcX7Pe81cYDC7nBqdmbUnlevfQ+zi1r1M1fupjWuQrFQrmmIDsou/fS/bvrynC8HgNhELO4X0o
gv3RnoX3xYXLx6AoQtpnNOg8aTOrS2lvv2ivkIOsGvTiv6TcwdF2PRfTvYXtrkizXB7es8YXJQcl
E0s2VgBqzZmQVbb6Pqs/HQs+SEFGlo6K4jen0AdL0+r+pXwJIWQN6QUg7lREYbXfSa0MQwPgydx3
SgvTJvdC3KZs7OWYtRGxYhDVGyOc83A9Vun+broOMhASy+oQLgHZ1wiFHyV6F85kHY6lH2kkgDoR
4xJj0LJm0eOulnDDqbf0upPgoD6aIDml7Ulto/6eWobKXmwDT+9ilHwjZblDFCrR+/Ms5G3MsUSp
Vw7HadjyZtxmBbJJB1H4mazA46F1osiYo+iD/LN0asNnVl4pTx+71azzh45IEhJDGhcJacKKT55R
SLV7vlRf5jA8TVaOZhiiRsRKllGiy3P+LmMZGHZ/PfPfYJu44/0p6doU5q4nZIo7J+KVd6FwV9My
+OLtaeoCrUvVVJNDgwkGOFDC/NI9yolfFPHyAI7MsHgEjfboVHc3QQ+HVtYFS4KuBoMhuXycymfB
ds715tr6Xp1/uFWI0AFnji8pOhBxjkb1zpyC5xG8bHtHEPW/LYlJzns673FROpwPB9R9lFc+GI9M
JgoT4BTrN1w+s9z2dP6W5fBEYGPlrN4EMKJyTwaGHMU+OUsuNduorM8btOsKJw7cJ+KXdm3M6min
JQoYORY52MAwcvlGwRAMxQbh62Ckcu1tvuTV9ua36h0ZnamLod0QjoY9zXjcrj+KAGSFHN6XitV9
Eb93KQkq2biDsZCRZhaGdTF/EfhLnrplhMTTRsS8uQnj4pbIZH3bYIKzTQaufzKu5g4Y3BpxvO+J
ySpFpmo/Y3KbvFOfq/pwOfisAOuK3MhQgb/7z76aB9w4LdNhsMvQVqVzvFaWgl5gY9Kx7LraR8Yl
Px0clPJL4YmP9GIVqFLKi1eQZRA8BFmAg/Ha8zfVFGusFH7JmvnjggsMIgEGUcKiyy2AO1OLvF9q
QhpzJgyLWra8xt5nwId1K33VsgDpYIXCBNoFvz8CEeqOHOjK/DRREVshCuixVdLQAnOZOvvCMlUm
I9etFLcN41tH0S7T8ToK9eOUXeBhELfsuKTxsUeDiymDMR+UU1huzXI8ar1p3g8x+YLbZYbKMirS
luh5CGKBr/9tDmMDx5+j+Ydccah97KMbnbjA7OIqtMEmsMf448qEft1N9UUOgfxLPT2/RkG7bgGX
mKWf/PFfE3rD4lGxUvXljuiVNPk/0dGvn/59/iuN+BqlK8M4Sc2NoCe5SsNKEMWDZXVUpP6JMVl/
BmKSmi2pKOmqd5BMTKq4bzmd4IiW/beyayakztg1NkzDC1IzBF1x4fKNxBW7RPfCJkim2YpqmeWZ
dlNtOPsiRqAZmNUkDZrfNdoMRQP2yroFkJHO+upxRbCVA182jvyv1OcF+a81h038Ab83K7GSM3Lo
0A50zHhlgbjdUT9PU7/QsriyaL0grUd4LytFvaFdxRAKqJW0sDRYdNEDfu6U0vivIs8tJ/Hyf/u0
x5dO/hVxLGWsAuJHanc6UbAH8CYs2EDg+FomrZaTjWggAyqR2eJWiHfjzQ0JfiV0sJoAB1BDcqEf
OPchsQhYxdzLSXw9NIbEv8TX4Xctsfvr5yQpcALPkIbBWpets/VfK86kU6vmPf03OSQt7wA8K/LO
f4W82vchRA8R9czXVKC4hqgvHFKA0+GJbUdW9S9QN1BWLpLLoCtFftaabe5mkcfSbTe8SsZWqUL8
59vi2MeX/geEdAFewwNrwu4/VgdETOLQbDHMj8ZMXBP3chOAEwxBHlUXPOOE+8VXSj+/bmAqtlso
TYLfbxoyv5AslXLrctf4G1+4eWQq4cj1fip4oQZNtjIYu7BYqN3iAQoT3GNM/s3RGEhxQDgDRmlB
VpDK24dW7OZQeQ92PDPJ5ipp+ODtYP+ivuz7f9GKwiFqbMx++GBL2sCrXUQQF0AQo4TL0+neGvgp
1uVWlaMNXeUECig94ol+qox5dYWaGq2jPo7zjx+q5WSZdUwG3sQu64AxWT++w1HHP5p/PIDXBhuY
4yWS8X/gYce7Q+uT9azhlipqimgaFXWAhtcTYw19MUBl2Xr4EujWCUfMY3EQLRxrvLXVPSSdCWIO
LLA108uHcbkGABUwrHU9ZtBzWuhHIOBNTNIeNxXEj/smk8KMJmkj8zo0Bm79syyvbeOxXZSvaV/w
ofK2jxRYURGc/rAuWhp4cZFwEINltSXbk0105SSkwnre8GX8S2MtzcnWYYz6VaA9MNgRCR9ssytl
60wPMy1vLVme0kXZMiIuI+9Y7h8IG/1y2TV3ada61SKZFeB30Xwyp5IoOWbdkDFpZCmMDqiMuTAt
QtYxf7GWdJzPBdjlwvPb8bciQ/gDH+KPWsbO13cGIbluPz5HcCeSFsTVF4QVlnuSyLnVPVMKJUoh
LQlUyEs+Xq4bKNmOk9+nIF243C7Fgm3DQaFpD4Ngfi0FUr5XrUrfRZPKYZE6SMDRv8BNwDFXVt49
qUx4SS+qpNQ0sdSHP8znuubgtlK9f+qTtpCOe40vSjvgX8levy30CmGUmzwLntacxd2EyWE8mBjl
RvLdioLt6kuZHkQpXP0DFDI/sr6JUkilBFP7H1YlHB/mO30KYTuFCwTUOQZE4cUiC7Fq8DD4Exjf
/5UBtl/gk7347X3rhf+STf4H0tX9pc5iWmtgM4CNiWyGMD5mPu4OfY3KsV81LkCvTyDVy7c3Ye4S
Dhyj15JdS8mGoNxNj0NRfHe+PP0I4dRnnAYy1SCh0RO7z3xPRMRYpGSGqaE7B7Rq/dUxFSBkpmaE
0916GJTAPDXX3aThF4TNfxBumvKMpYoNH6dZxD4kBbb6WmFuGpueaXmiuUkQPk+j3+y1hfAD6Shi
sM4AAUGOm87H38Hy2j18Ae//wHg4GpFMROgyunBHtxqzSkmUlArLoWzB+wUWszAd3huWJ8LxjFeF
P2/iV2kA3X0c0vXRbItlmyqo0CurkqaAcIjIRiqmfS78pYR5BqSfbbfbeFqDrnIxfboOsRDGhCCU
LaPPJq+NbF2qyvnQTCWlCDFlJwHgj+GHtO6i6Ga6xjb1Y+8eUQ4MvnF8F1cbvbisbjFVwLvbTksb
KxPcVHP72MtO0PKfDm0VMFtv9bJ9XrMRnIDBAh1p2ed+A18DiyMYUsHKyBraQiHBkxAJ58hivxUI
/wZ7bmiXaM5D1FB9gNdq5LsZ0YVVPlHpGnq1iLABgEbJyoq22nSi9NslbxVy1uBMoHeRxOt0V2Bs
CQwlWk7XtvDChoueVVMmiFWZ4hEyDRvK0giBPCfP+ytZ5r6YaICbU0tWp1dpv/QHJ79B0c6xrccw
8bdcnGZdPXhQca4/W95IBRuBqFh+5xkAQT1koBgzH3I4+sr9XReXlOXcwqW4Ix72MMz4c3wXWEbA
N2pmuvhp1H6LTpSD4CXuudpQTpPoryUDSRKXZJqyCEtM+a1zOeYecB4ZpE6f3zBVzVGqGB3mBPt5
2kJgglGy+wuRitUGvFW0SpR4Z7pR2jf/THOylIiWQPc8RVz8MOw8U/9ZCfiy/43rW1nqpwYcNzoc
sB2qg1MDCZT6Pm/bQZppJ4+Ncf4WOyrGf5zof6PkKLZ7mBoY54rgemoUi3PtiHmq96cm/H+SCG2H
fRKZEp8wccXavb5esxmsBDgIMnFLKZXtsKiLZaZcVrHfHoW1L1+zJfzVhJsuMJ5jGQ3Qmsl/R7+n
Hig2097pVngpzPOIFjONjhNOStSzvgvFCyPL5GcJhcN6dzCN5Uq99OyNxl4gwmw5eChH89mOSNNq
RgXya4y8LKuWW/GnGLoqLPrSFEc9dADxCaYRn/RvjkyU/73MWQa2Z7/dZ1u4gMaRQgvp3qLrYIDW
kkKbbjoGuv0vYqFaXjYZCYJ+w7pGr7QE41+qc3WcAkpj6dZ95xIq0LJig3AJY6fnDQALfKtu9OC3
H0Qeeu8bFLAPOqYmoggqaVncBY2O/Ynfaw4PqUMqZWdk2wVimrTtw2fGtSIw36wkpOmOJv+BLEw7
oy5qc8h32wje3jdzJDbYi1QVvgFoTJBx+mYq/lMRoZGOmV/l/mNu97GlJpNee96fklets3HV3xl3
S/A5Xs8oFPxASnx9zC/3aFufpYaSHfi82nzDimp0093aIox3nx8LSicEEmSWAc0A3+mWPWE7fQIo
hhmXsB1K7ZQcyh9/Pr/ctZDv/TBd0vweSV1WNxYJmwEBITXA8N8P/R4xarKu3EzyXmdGhOb+HMY8
F9UK24mYrS539132shUFdkLoc5ikZzmvdD9Cc0F5Mfio/l/kHvSc2PRlsqzzDwmLOF2/+uweD+6k
9Jso5P72zuJSZSuDIBMUFG65sbViJo3/oH0bajsvUijeHXw0uwdPECZ0QnNZHyzQrVoDQniTCWFf
NDzcyUjTjI4/P/gNHi/J0pFS4RIATwDsUEWuErCeihLKJj84lyAnH7hfGxNDAIW+GhqxHcMkGp4e
LjqAB2rxZ+rfecV85UMWFneKBKmDoy+bwh2TsMM8kifvsQIiQSaQuB0owORKOAq/Tg+pf0GtS+jD
rm/AVQiQ1+Qu8YQkfbjBpgg9nQ78tn4gBhc4boGzu5XyPB2/JCcWhLimg3NtVj4o5FcJlHCAVYn9
XsOs5hi8Nk/do8QsrTnHZWKTd5aGUwCXt4N2TWcuaUI1fk6p5nMgpc9e7hot3gPyxoZyBYJKgn2X
v33XU83p5y3K3D7ymkcTRhKj+KWHp5bJGgNjZidGuSttqyKnh8Usa6ZytquG+2HcLnzCeW2z6nB1
Yup40YwFnL2+19vIJJuAcTqYhajoCYTsp3R38X6vUwo8rSL1fB8ckv/HCTKtbNn3b+f+JIeIryWT
oEQQnAfLPJ+gwydWq0HVnoIwoRavzsJkkafAhaq0JtIFb1F2ZX0Nc9fALBYozcxMr/YTADBUeKbq
5fg0D6G1MdRHJLT9zbZMG5r618u3noZAn52HgF7Ku8OxgrJuZKlzZF+A9LlUWHmg8DeVSEai9x7w
8KS6RTLO9VhGQXa9toJszCNtJx5+SNZvL05uxP25GL9m0+hZ8XWnTqpmqY4CkeCxXO5VwrNmJEcq
hmxdo5zf4br04MvKtOb2Hvb/XaGLhyCgx0dT6RNsbj00dnZwSAQUHe0/I4zl4/bb5Rm8V6QmZfHl
zVlDkt+095CfGSdYe6K0m6WBCSu9Cy1FBUSzHNllTnKy/OMkVm+vbYOkCilxPe7AV7IJDwgBvioq
BRgJvSfxAyOBvT3uKZWl8PxxJI11xHDKFtzMSXUY0vZ0fZrYmkt/Uv6OXMb5Ssrcwty1RVOtcpPq
VXsOTx0PGb8NXqETByQOfN+0fRR6hsKtkG4HG5MMHLgGVZauGKdaCRIKdL4UHJ7aLPOwtOq4I6B9
1RslkVweklcwGXDOwXt9Rd0DlLsfaScY0eJrErQ9lH0UE9ESsqq+BunFj9c2Tj4sxSJgMclpj5iI
tw2Km/iQP2JmcNNvngXe2eY1XWr28JmSRMnwHtvSCyc6Wp7kj1MsKieoyO65TnOEapaMwpYWS16J
PLRvSHx2GBHlPIkuQDPBfEIdEdu44/UPS0gGqMO0G8fdu/qZFQA+X98cKzKIWoAH8ciiUVIJ7EkH
zZyTAWrN/J7U4HGRBKJv9/tlAdKU6tJNyNeg3eYMJtmBuV3RfMTIzDsgEEC5i0vv/N43DCdG/Il3
+7sq1b53Bu72xpbct+Tf2A0GAMld1cDnCqKa0a4T1ezbvKG8OjXb1KMrIQkgKHonOeW4rpVqNcYs
6n5V2HPkhuHXCanEDSznCdQjJJCEhoIDKObZxDKgzTpBhSvWMOKdwgMHc5KGOmqLElJJdLBDrSZT
X9t476g+9fQVNg9ENPU7z751e5ILY7IdvZj+qBv7f7rMNWBIzneIX3l7N/723eYg0jjiIcX9r2fP
zfvjbqaql1yxtLzCwnMjSnpCS+OiUW2DUWYyJ8s+M8mssFe815djL6yc+VWZXyzzNpYwbyJfKC6i
PITh3Nz7XLocrRKVy6gKofN/7Ohenu751S67lgUaAhimeeP5b9OfZ6rsMysZuf89aBYksdWLPAn8
5ZePrGhNcJSkJHgRKAypalXh4J7nE/tehr3H3jc6fVAQlM1+UBKnyfIrNpTZiUl2/cL3FVzSlB2z
8IRUIB3q2LsMTIERqHJxLvb56sJHdeS17g3moz5UfTrsJkrRTjNBFgDveGkCWI46COp20fxYdiK3
2XSMvOLbxmdxS1Kk1qrpS3Tc68oM5aARAjPeQsCPgwH0099inTXin3JeBozWlJqJ4O+/Kuq4IBSQ
8g4UeYHoz0RVCJgprKAjvZn3fzKwmooqgEIzyq/galZOhbv8z7QpWByReqRTCjctBWBSHAzXvqp1
oGth0zWs+7sbMzMYniaNnIODHhC+jktl7mQr6WS344h0vPVkgHRgNey/0GBlkqXsUOow78vZo+ov
HEXsNzP8lQMsN3ffXnXX6tSqgmfJCKxlrwhSAs8DJ8sFytkkfQSx5SBm20HY+9R98sQ5yQ6zc4PB
Ng6bBRdz8RvJwZrfp1lM9B1YqNjP/IbOxCTrLHunQlceYBvEwpVuVRxY5e3QDJ50jrIiehzoSY73
ZWhbrPuhXbzgkRWDBDj1zhNqc+luTuBBWZB6Hbp0OT7qxxKHKhxIdfFKhwoRGLaG2yTjF+DQjtLB
7HJOUH83ZOxA82eLdp31WGjWjNClpcDlRi3fWQ9oazmsYEnyQON4rr7UbphjPuFSh9ZqL4/TLyu7
kOv8FeHSDRk9SpENGdky747Cb9sa2u5MG1lFvCGDHrzNbwdyKA4StvL2i3MKQkjsY3MUfG9nfiuy
G2DFC5+kQuG+4c7ZyI5SPbqFbE09Y1gv8f0SgKJGe0xG6JTuJYAKCrYj3RGfru1dM4DAV+hY8GI+
0vNVk+oXSiS71cNWTRwFmX+J1u9QFoIipWD5D5uo6Cd3ntOmWCnaJYrNby35yOtDih999319YFCA
BnAOFF9A11jpXKJGiE99xxeO3bCT5YNhgkYux+m8beYgr+1rEC7gfAtklZvzgqJsxkiX7MHs1NBk
6QiwN1PckEOJ8hLPKW82EB+PCCCHnb9+FWW/xEaiEw6FSlB/c3uPmjr6+yUmOlerCZ47+NDNTeRN
a5QtNTmwCEaSe7b8wojCnPGO3Pwo/YvSRkpXwN2D/R4f6iVM7BIUN4LY1Fd3arUmKWvniyTtl6x/
3Nb2oqxjW6+Q5yShl2oDAiPD0Ag3iFHNMGpl31sT3J95js2v+FXpmRB5oCCgKkJJhI9BTCetgvj7
2jM9tuMFslOtZa60y4GwjpvSt1qVWS3ee3N5TJrJKzFwDSFk6K685qXy7wzZppsHto1EAl2OdqRc
F89tQqpPMWU3V2Q6VyQotXvxxkrglGUuxzfZbNx8pELf2dErBOQHSNXZI9X+vN1OBiEM0Dufwcp/
Xiwe3ScPekaFW1hsYcxT1V3iUMh1lEKHfV3r/eCOY3tHnc/OXxotqha47U+NpV+wha9enl3Qq3p1
2JjQlryDmaOcYRADUO6Uicb3rFnoCEM6VkDVI/klp4sQpq0YecXhMHCzfkE+UEEqu8z2S6+FzYjE
7pugb7a7r4FVZtBUkE/wzYk97bGofXfiiinwx8HiEgPmH1/LsHNKmQPV3HDaNbo2TqKhlmd4qYkz
+gd6+aXpvPNahKmvtvW1kCxzE941Hxg7zFz3+k5/on65/fbFI4w0UjTVppa/XoUfKr//P9hbSEUI
nIQ3da2l2IGLgYIXYfIOO2ldzP31YYSnBPQFvF7zvz43sGM5i3lZGKla+G0PWvX3R41/0pHpsaZ+
460rvE4zwTiyQRgxgZQ5GoletFZNAQzrreHpcNiUU0lPejf2miIw4PSauytgukY3QwJyt3qVwJ1n
10XsBDceKJ4lbzKaeuLy+/wbrFHVjpBhCBcfE5sO0CANYqjbc19Po+Ts+3NczoZPr7vSW6mNpR+B
AcTrAV675ywnnpxY9cHJTFzWRirl8vLFihBp1quTr1J98E7EMCdtz/OLtIMAFAGV1NoI/Ny+LurV
A97hFmBvJDWU3Fq7Lvnb0VRF2QDOzv167YHOTLjrJ/HruwOp2rhon7iPjqZtuK2n671fM/x1Vuxo
5e/ZdXAIsC9CzQraqSe6B80CVEQWCe+bzJblXgN026ncQHu9D6INEfTNq0UJ9ETgeOg+xMvTxu6m
oi4brU+Pf0mSD0BeZRA5jNt529PWNqQ5yke80xeFKtUSq7VOY/sGYfg9IkWWQ2bQU60/xheL29py
BatB49xDidWivz/mczJm1Zxa5X/IxFclM+7q+IGEape+opeEXFc6KbX7/hpLFpV0MJFF2oPTpbHY
1zzS4hIbIl7tVyAtfyfHGtFGAKN9fw2EGJIQa9B7PVT9btCtZ43aecRcppXy7TLPda3a+V4YvPa6
p1b1IUmCfZDt/tTqnbakPB6p7/Bu5uXwm8CHah4BioRi1h86pJ9yQCmoSLFWtRM1PyO5/7eKKalA
0kDM2eVHKlQ4LY5HUYINdv3x+v2L+mrwbsADGSB38BvA0O1K8vCuuDwhKIlbVrfmYf35zSkxp7Wg
TNblbgLYp5LYxS1T3Sz6YoMe+l913B5W52I0P6iROQvfIIay9jq8tbz2PmwWcZO5AiwDFYJfyGlM
Po5xtXr3L6Cj9S/4/HRxxqJBSd0nEkXHrDlFGC6fZhOmpVWSBsUL1KUvU6S3/h5IBRr++VE5TfXy
IhhYrukzu9vio8Y7QdIkqXTWLzzjCVEWwJMIln79jKVVzKT0eOsGzXC87mJiOegZ3mWZGY1JbUOf
ig1zYlXFyb7n1BucNnmgPIXC7Jf5M127Pq6V8hlbPDDlvy73eJ7+UJOhC620ALsiMbHQNfVMg1LG
0zFGU1SP+HpuS6apPVjggeto7uSi3OQ5Yf6OEx0q+k07d0bRiWK57X0iO461SghtdITc11R5oj2q
2yOS3pauAne7j/9riTI5lRr9/CHpP1/wUDXH7/eF49ITPUtGmNPwiBxf7cAXKLALw0/PMaCXAIof
eqtVQAATqqgkOV5joFspEYE4hWHfg9Lksu7i93VO+eswDyS+VFhxicjApRT4vbW0K79ryjXRxX3Y
sqPIZ58H+dTu3aaACl9QqjYLESSAiHHmCGeRWNpxxCBm0Nw4yNlPsO+D68dt3SqKaL5quc9amji6
MkjMJ58GiSEJJTg0ykJUgdGa/ImpaLMWzJXEdXgS62sCCHtx+hlCEDLTlBRGM9w2HDZAkr4j82xu
hiLymZohv9w2hvXI6ixrDrsSWFjmtHc8aYWf5P3rlAh7L4pdOUGzYyopWgOp5CSqIJYCh+JiB9/k
OLAUPhMA7y/M4Zwx3Dn0pm1Kc4vjcl25Bj+bGgpFCsfruYdFBVjpJe9KzGUDaDWgg3y81DtUUALM
X02bkTRhq47LJOfZ0DfURxqJlakUyz0GaxTzbxe5W4pKm3iKRPRfHf+WH0mSuwCcLzI6OBrAcVJN
x8sqGG35WTScPNGKfCRXcmz1FHMAaG/NxsWvefyxnJLRKypjfojZdrVuFs8PUUW6XzxJ5E5UA6P9
PdxaIxnYfh0vA2BA9DiYP/+gvnyUv0OqAi0Qw66yLpHy/+luDddZhm1WqaaXte29acDkOB0rxpZQ
fF42Bd344zfEpxbwDQUvW9DedzmDu0EwXRxFXY9/umpNZdNlycOzSxsGenZbuZpU+LRVPzTXeXxy
xJjSdQxc0fhaMbNc/+E+6Js6suLNxckaUS1DZFEVv/pp8kITd7BArtPMLQ/NfbHi6R7ttfw4oOlX
2yaazP7P7pX9Yp9/HXnRf0kivRTGAcRAz8XC1wngGTiqzRsuekYsKUeq1bm5HTw8hYXjkJ5xwFe3
JCKAqEDAsg+G18PS1tO0xnP22g5RKypc4bZIC4YP9xTRBgLaABVZs2STsKXyuHeYLIxMO/XtbdYz
5iFaa0D979VV5mtrqi6mGHP7ah9vVHXqH7inUwv2XlNPr/hBR0GvNhY+03Ke13pYgwSl6N5ocB3D
H57nDnF0JKTmSNlFy1P5tmT4DlQGZCNKILLFJyW0T2ZIjb5ioWn7yCY2Qazg9CH4G+IxAaP57vop
BEm6s6vrDopJB1WBTE2ieSOIr+3od5Klhn84nTncDQrZbY7mGJx9VQazFeuRQIYgmheeog4vYeEo
dy/sIwX8gdyHAfdnnDSkbLwC8tC4zCnvBAaq/8YkNRaCALY3ESswHeXbLU4COHDh6aSQPzp5qYSL
4jySJghEqqzXdY9RS1L+qvb8/KDtIo7lkX41x9ozGzC1KgL8fklaL+WjEZw8CE1kKDfMIC17ZGyb
4kc0Np7HzY6enRwqcw/qdH91W11Qh/tlpwwJdAuVlI9QDoXJ/kam8C61wxEtNuMxqk31lxEyGdg4
qiDa6qfLCU2L35B+pbLIzQVDrcuklPj2Dmg7J//dMH2JlDhXaM6zw0InyUhXGiUXRg9DyhIcYGwa
LX/faMCNBUJQzWnmCgmltLWoqtkpdi8CJlG5F1czhmbil1lXJVhG7QmcHUbwYaQ7FmpPS0TNmcHG
sQUsGK8zbdKZEOCyEjkMtEtebBvcqd9mSvY8W5XLD6CAqwj6OK64A/+zcJ0Y6xsfYyD9m0lwJF0P
zamOxdTHqPNKo6r8/S14cc+HLU7qcEgj/M6vUX6D9gp8XbqfOGoI+SkMYrN8Q8y51eL9jtJ0EAPY
UfaY3e6FVAvoKf9Ywcf707FfedZsNg3T22K/ZyqRGllhT79M/kcNoh0xGydf5ANUgEfxb+bNUrPY
qUBlbd+VU2zSZ9CeElpopsRaVWRfJZP/CUzXHO29DTtFchszt+WpKUhLqRWZALjH53M1p5LANln1
EwYgJ3liV5p1nJ0MM/AC9iz8MPgCLJ/At+Fp1b3IvhD8Yy1+fXDkD5QXGqptame08Pcj0ZeFmVwB
COAh3LQ0+zk9FNBrD7yIhJKoMOLnPeLkSrYjIVYJAz4bcAMSR+2+GZ3TxrLcdJD3p6RxMhDQ8HoK
jZO2qM/x9p0/8VobPm0LbzV6IYg78ywWuUwuBCO4f9Ae6hn6sOOuJJoOPa1BWlHAWZ60ikcN66nJ
4AsJi3aC/5eeGcqA7ws+ewJueAEKMonozPAUq+NbgaID+ecJg9X6n4/84ipvPLI+AjeYLK6kKaUC
uaN0EKah1vWZLMJJbiaYRukkpX+204DheWDNfk1V5SDdXlFdYDXH253Vj4HwWoLlKiT55FGeBnY3
2ZVbRzXbq2i2WUSKo3p4zrZ2SFT6GZL3kOSbkUW5OlVHIat2LSG4A69yJP9Hd1MBO/UyyW7q12kM
CuPyVkI86aFkpvJvTNzVO/JdNV1DCcS2RadwD+U1F+cgSe8LChSldf4UtO5RH+yQGe0bbf6Pg75E
fI9oFvDDZUm+HVt6SRvvPCvRhG1OkcaxZ0zkLlJ1fD4PfTsdrG4/E8rw3e8pEoclPOJSyyESASO4
isCBmaSu4f0C6BU04LdAnbJxoUmbNZ/vIakApjuWdZZ14mX3fxNAkDXfs3qih39Nc6GymPxyq4B/
SaofxUezABDJYDtnkl8AcbfHpQgKVBxSDtTy6PbYJv3vZZB9G1Y5djlJJhTtaADK8Xjv1SVrz+hz
Y9PScXfjnvKRH2bV85Kn+e1sBSfOMeW3YpSrebPISg1ZjqTi5mUTYRUiCXzVdI9o30kmPtDWFgXM
ujm9EPtb1F/lkASewbQaSPFhJPxvUZZ5J+8x8dgqOyvCVJloUXWWbbsjNLL/YvMIsJ0c/23qCbuC
l3UoOS+IIQpSZPlVSwvJl9LuJyBpNztXo8Nx74lah8Y6u+r+yOKloCaiJQMVBJZxQ+yMdLo+Y46L
rsvyAD+9YARaot+Pw/omF2iMh3EieMdPXmaPiMzuzFM/4a5VjvTctOs+NAAWifNo+10z7eVjEdBU
0pC0qZ6YsoXDxI0ewUFAwfeN1kOgbkGh8PQuNJKpTuq6Zm4tInP7YSbkseAa2kUOihYnavNe+dN4
SkfdKruNSeh9Z38xUPI8yXykAm7onyPnQHuLmg3614gZUmEoh9bffjP9CwvS1YTxIlsRbjjo/Mz/
IGzW9PmtPuw3wcaa1rsSq3FNpOylcCbeR6mbPrzagJXNX/AOABHP/1s7wMh0yaWpeJ9MpaMcaRXp
jsBuBvNzkod/2CgoEPmvRuvMdr96Ikp2WkwvqA6OeMX7pWLYfb0P7pPQ+8ZLyiVTm65YeiYJiURf
XCavC5e0Aj5RxsQfKQn0bAitFqLtbcwNnpoEsx7sfzvcRzJGJUMMpV6oHiXpIRv1vbpwa+7Lmhwy
/Hz+XZ42/ic+Hqyatzv4tFk4DEGInpahJlxC5+2x1ZT3Yj7K+cYUYxM788DCzFyWbmJ2/55yFxw0
Iu1nAnZLX/E/VSntaFl18tGsyoL0b2D1zCqW98oM65VNMWO4fy5tjjJIj7BDRrvTIToyDQf7mwFv
7c9JjacyzOfJsY52uLFv1X1Odqyzk7JP+xd1QfIw4D3kH+96UIE2nM+krY9ZwVOUNWhQwkiCW1Ht
p/vO6j0J5l2iaC8OZMamSHYtN96SG2oQIsydYuONs+tRmwGYDaksfnbIKzu712wTbE30UGFkzBdL
vmHwos9G/IXwXK9Ajab+JYcdUrWbzTYMxYBu5sKnl0R2JzqxC4uvhfCwXdJ8sWZapyHn3kDbL+I+
PjA2xIA+0oJd/REx6Ufo3We49idxOsCO3T9v+tUHK9u8am+fXtl8bino/Ip4QaftdVEcyg9m7Zpp
mCzsOCQhMbDQnOj+EJxDODP2+oIPuk+kxUdQoODQaccllURRRNT6R/hWEyrkfo7mrgJxxbUfcW5y
/Y+yrbeXZPIZQzw9Fvlk4R10jtgMvBgj/1FYbY3psjEfVwz5R765vYOL+ni9qMwl5NHJSAahnV5b
0jvjsXh0bi9zvE5Kx36EiXmkixKc//pwpSHwDakwisfBUCTZwWXi1jtF8yDNU4Y4/slHMJmQF4Ui
E9WmfYUsRbmRPyRGSBxa7XH1MfAz51EDPQT1GVs7a9NBB/4+nuqgwKa3ILQ7X6cDgde9OStdXFPX
tuO+DHy5z9jyknTQvmzFtfBlv8jZer+xw8iCHYNmva/EwVkPg6j0LyvSJrhuNWl42DcM9eoQ0Z5Y
CrGl2h8GG/og2fRuIh+1PaHS3nebUG0UB6IO6aWeVe4eTvUZfjGecgFv6p2jw/cJTkCw69B684Oe
ieLKeJ33CXOBnStLlnbhzOs+PyHBdy8fr7KMOVj115SCLHieNja2FbDckzWBw/7pVLlzGzc6f1rU
r2Lhvsq+aWw43rYWLrnZLao0TKxNE9Q2edOKYbqss/keD9FYeKtkYwuczbP/cZIwAdiaHIjD64nZ
bbg6sAOTJUu/fi8YrZAAq8OMVFkpjupDC8AZplrG1jFxakmr0ITKDW/sKFH7RGvb69RspHX0rhCg
9fR3yXewbD+0WtptbI2Ko7UOrjbYFdvUr37YOxfBEyKUYRssImDHGQ3/bNAEpQi8VGwG1r6Qx/v5
1vU/jp0Lc/AjHyqsxJ0NN7WelxnL6pDiwcbCD/T8PxCPpjKZ2MRc2MZ6GpR/bpoa0p88OBI5H7DI
nFBhC18Mo5x8F4flVtO82CxvAsHPEcUpU3kNv1DYgNIinM/yOjTGMVA86LSPwSRuDFxc1BNlSxYA
5KWEpbkFk5omnklrGwcfOp+KF7zIXRbkCnvaucGJgPdnZ3G5GML6dUFftCZLD920+A9BL7EsIhkF
PYOnkewIC2KXkpRUhah6L7BXxql00oRyz5d09biziH76JEPBkPoeXtOF14UjaSH6ndIPjSQiWfTa
Dvi7C1l/ReqyKpFJYSTqvQFoTjcFLrhC32264L0oBUoyQhxbn13yCe4guoArmraMWqSFku1L/Y/k
odsGkbtobjQCVjuecVV0FWuY4eYgoa16MesyhIkL10SU0ayelvq/gBzA0jEscmiGEUANun4vwdY8
XFXJNQzrJ315SAO6MsQHK9osxIJm9U3Hw+3z5XjAGT3V9s1hMXPkCI98x/zFwffwg32/pVB5DrBj
uyCwvckHgu7dxynnkHuCKFw2K2Mt6STsPrupSVSx1m6KxrU2W8xjLesQS5BJ2Xme9V5vtRv6z2CV
A4xcrsC9c0OSAnfBmn4TjPAQccdQzke3IxeNo+jB3IpPM/DjTKSSyXH+sX1HFK2nP85+eC/XaVbN
KYY5IlykvrQZee1oouz9EsksMtN0LuHAZD1PU0vW6nYSPf5gcs9MFzPTmxpZLThttp8UVbx9k2vo
yXgEvAmgXdVx54CB3DoJhFd1jkisLufb8I7dcxWPK2cvyz19mmkyByOTScn1axrbQCrDHUqbqXpp
QReoVL52S3rjzfjPIucg1f34Ul8FATi0Uc7mahiLRsvXODYfETB4Ydh5S0GqcILA/GanOF+eTKGG
n1HW4a/5zmL9VicpLwFFrJ7ge+nJCx0Qj16R5bUFTmcOC8+JzS5vIbfpErwh04t0fe8E89Ew1osK
DrU6ilT5trAMrM2zk83iYun4eEh1OuLK8pVsj2l1hmRE1HoL9PododxuthD7tli5NRdV3A/8EVN2
92wm96nwxLv30fyRYSz0Dw/2F2cJtsi88SiTxw0bfn8Ia4jnCy5P6y5xrkDiEYIIsa7k6G+E9DOH
UU3PsLb5cvjYlIBHB9Hopbkf50cwNhfXoFgfoYgMSJ2BqdgulwvGSuz6/EyZs42GoU0dhgYLb4xr
rMcn34OYipcfjGwQRSmReadYvbkj5YtzBPMtAB2Ia/dmvgKKIG6emOrS2fm6Je1qAkoMi5XXERJ0
LtdmHLUPYshsx6od2uz+wl0YjQaKjoBE4ADZSQPT8Ad2FqOpg3BPwdHWc773y2D/WkFBxSmCBoL7
zE+QMMYdDEeMWgKUvExChQXGGMvGDxnPNmGA8t9zs1y4SzPYIRkhcgAo1n4tiOxcXfq5VvA+a44z
YzaG2E6RKoRO9blp6Xmf05G5jfIZexJSdk4Jtt4H4zZILEdlmZ5Fo/tBXmNU26W8j9ZfBWBHhr8t
BBJlxmq5WpqWnSQ5PEhjmmkH/uKR2Cc6DMXXC6D7AXYKWFIS9q1KX8vY1AjG2TwXcWtNymN0/Neg
YcZxEPPBc+j/iwLp8vwjse0/VSghXGQ7D5uE82sQvDTjLKbXv1Ov21Z1uX8/g5qS/DoqBuxz4F8f
WBVT1qQm0EulGZlFWljX+rSe/R9vvihJqAH5T0B+ZzdbHoZFqEW+i2rXviLDDPlpQHs0Whiloqnt
9XvHd2l4apkfZxlFRPh0fR37ZMWNnL9Xamo+3+3jXJg6PQtj02AroFzY6z5Ys2aiOv4tptLbXId+
1petAF59u6coxSbqvnRmstQOdQQlZXggrSfrNlrdmXeRgWmCT4AYiVNZDIUMnLhVhKFPtNJICDop
do54T4KLmQr2qsiDoclEFWklwGewe+MjNV3iAQuQRqUIY4juv05wSprEOU2rvXVfKSQlCDqvdXLE
L1yGKQs+cKCoz57ZXtriB5DHae4lq6b6uW/b2KcWi60qBboJ8h7enuKHek38IHuxSO5jKZDYm9gP
IlSBVF5pfDttb+3H1wyNupkTcnvOOW00chuPPzs8ajZoDAfDGKT+d48iT1qSjfS07v25folqRLR0
PknFdz5YFFEgBrVgEJksV5NlJHIo4b2ijcF9lCV7AGr+73RQu1DJgreoT5fKqeus2xBYmNk+rrPA
JbhgI205DpDQKKeDwdXQVkoc7TlGXJEn3ZSr5RnqHYI1+BwVgfRbvhAIXMR+tPaJuB3+wQsC7g8w
KvaygLTsJtKOxuMhis/4EzTT5JHIuwHl0GlKqlRznV5JjP/RFPXkr/MjAkex+cSnwWPoJY9kONwH
QLAGeGkcBfJug2DUfSNK6jupb9i1z6ddxqAgyWq3pUk0juA5ePlAunVGA+HmxKmyokHAVsY8EuO/
5VS1y1fn/biEMApKJWgBuzBfi6KCoA6NVBmmgl2l61fGJ5lskUUdObTV6FhhHtJs8oFDbYTuwn+j
3rz46ybl0O/fcb2VGY4dG61yy7MIu5vSMaKz0GuXWn2hAFKcCmpg99BtvjKS7puDTO3X5cOVvuKw
ONrtlgudxkEJkcdugrTL2RkI1H1g3+PNLblQ9u7lpD5J/9D70g2Ja6ocywUiayYL2rpCYdxsomO7
x4nphOa3hX35qP05hurEXJgH0qfJv2s6Eh6LbPMIVC/fPjBLEzGRqqiXCHQA1WqvIWTtjehcq/ED
4eQZj9eXKFm/R3V7xlhTN/43gis2uuGjcO7Ci8YDtX44++G2h4T32Y8lxcxIbwFU7hmAO3rSC6Px
mqkybsx/j9crhE+Qt3IgY8MYIZ2Gu6eS60VQW+O8m8d/r6anxzGYiUuB3MXd3jeZwhGlipD5W32y
SVN3fpYQ7szlBfwuO4x7oGFb0ZCJAkLZxl3QLrdSvw8uciDLoGuotD1Py6LkjJbuVZnocQFtQx7v
6SBCUytOkz9j9EJetKQevMpjg/vHn2/Q3a2m/TUgnGwRhJkWt1+nviXajw7fUxjDWHvXaD1ogck8
vfTBF9qz4xhaIjOaEHvvyHQKXkMlhwdwu9BjuD+nGJ4u5qr3aur0/DyF/IuT4ko0rwj3O1UdjzGp
DK2oinCPuZ027Gz/4jWdhlcWssi44WwOjU6wJ2B6FK2BwHDq2iq6Sb+cEC6Fdm1iAlIKLiq2dlp1
plT/pMNrh1Jg5Hv4L7UdLfq/LWODlBoN1qCzl3eP8QGAOVTUehOl0PQR215R6CR/dTpjEsJYANIT
O9pB+/saYqQpO2i4ZmBPv1J3WeBxXFuO2xlfpcBVUsJhmgtX8Rw/vpXF0mBBJgQkYG3AYYmMzcDY
OkLLSsyUIMEKJyfQZGoAJ7q7XWspSfHsRVARbb45jx5Cj9y7NKwvcHGae7jfX5YoS5uqphNZE7Mj
jdSLfvji49dEu0e0ql0fmDQNSBTjX1NdI1Qg+yAmkz8eyFVtJ4jdfyCmjDIdLFvkrQnQIZv0dxwI
WxzEw4tHVc+UMFjAbzh5/m8ZGGQm1xEETQilJrgrIs/dAWonmc7/SXEv0mn/uwxvdkT2vh9QRvkk
b2yqIIR4/hKCQikbrt/5JqcNH0cKAPSZEY/Xnjgu3YBF1XFUIpEmkeaLMyIEg6YYsMZXXBcualXL
yj6y/VcJeUJ5G9yWnPuSuVO2XfxU8FL7ZCmC33zt3r2uRDylRxYwTUXCm1liO0uV3W40mOlDnAOA
c/qzFq16AWqbDqxpm/m4Y6+APA/7ftFHd4MPN8bUjVQjWwRgMD+9jrNABUw8Hl4318sXyunbVG9G
TYEehTLwXbfK/aFM8Cjz5yWQkU6+UqPbXLVCL582J2gMtR+whq0FcBX3Z+1PZUQJy1prUUcX9w01
TxIkP8RO2AmUKm4l2gBn6vIyIsaCfBdjCGsPb5PwDaGdH7AkH3iX1Q3506flAhF4Bx4WI0AdbaTd
ZGqTGgdBh7P44hqBFQTdZaLJVMlpBP5UNRWG5YSQf2dR0WpEcmhJhvfIXF2GWM50Q8NX6SSvig/C
5i574Gi5sMTqrJ980dlhjEjG5tTSAJrI28KfOkN2JFTmL4EIUPX4j7HaFs6lKgaEl+M7Rqk0mxS9
GzUTxLY5d5PhQus2hg/H92eeeDWMp4BP9Ane/AC5OvHN04Ab6HOYS8xRkFfeWLDFsPNZyIkGVIRF
2ofts0it1N0gaLJwu/vh/pVaX8cb0I1D91YfZvWkod+PKY+NJ3rlzzVdMLkYPXBKjiTRYld++dGP
ZzTg/4EWquTRGWOCfrVGQI97T8e46Ch4fd7zg4tHu26PCFyHpgt7oNP894TrYH63oFej07nQ2TPO
uLa3UajZWqaw6inbld3Y7RBcKVoDei5cQuI1+9l/E6pUe4QLI5aHt7aFuSSP1azqDknI+miFXAti
OJWRlmru90sThUaON3MoIsmHo9VMid4OOemjKWIBqZl6lfBRzfB9V9flIrBm5HAb2b+tUJpERNXR
Mcwyvw+ByJCBW2E7qGX+m2kF3z+FIIvV5Es2WhpyjTUJYo6oWEmnGSVo/jxZQ7lZjWKQS7ATWjS9
jPOO92IZ1TdWbOvaBJby/znf+sc1dbEdBQQs7DdI9w3RYTAowl86U6HK4E1C29haz6/j+cNUemix
go7aZkkc8JycrYwvUqscvVo6lIXUuPjPr4LXzCKnr8DX2jXh0cCkQqqyzqH9Zahp50WDjTIbtiR+
uHmthKqikAHFW/SCtvmhWuKbZeu79UOjQVor9SOz61t4K2X7Rk2InHS1w6Oa+Zyt+RC/d1/lE/Zp
sBDe/1AegMJCq7wu3MQJcD2WaRkoagY3bcNG6TJxGP4c0aGHRLqIssqRMZe/C4Ce2Zy7g70+KSpm
zt3a5sKAJlVxlAqU0ToxlA2x2MYsiSNDPHWrFFgVg43ugj5BcDmQkfKZK3AlkShlW7P0AX31HAxm
7HbfWWzl30LKZQSr3ax44qKN1LMnxYryBUAPwQio30u6v6ZYVQW/pnfIF6kyZTZuNzsLENvA+RlM
MksCp8Dx4h0Erh219uszp94h97EQIlTYLXaxKwQdAGJiFCX3iBYBYBN754kmKmbEPOF5639mF61H
phn1gsrN6F20SVZEuZ38sAA24kziu8DN3nCGe8EYIS98JV3/TX0zrqXM5oCg2EQEXhAHUsUmo6h3
XC3ZzLKGjLoTooHNN7UFLhjQs2RlmdhMuLNNTdlQfflicb997J6F2Ze3hWwbPd+e7z0sVdqo4eJ6
QupZ+Gr96FGQljtX5wFRNPP7UauryPWREtib8F3e5SepFobrNgDLZq1n79M+oClMjncJrlIllgAb
vrsvC7YhgQutSLpkSrEtbP8MAJRnJaASvv2EAY1NwJuH91TbKD3y2jPhVlPXIxHAK6cCsuVacm3v
9o4AKGKzP+DaeOg2cNFci6DzdeBq+YEl4iYWtBzI0BCyM1cadcC6BcHtDFC8qBwqblcWq6l+tuYT
yZ/JyQey7llWFaVc2dwya1qflsIgJMfCEMNb0Wv0+TTTyrjzjspx6OTtDlufH0/Nl1jOQDS1RQed
TjDxPeWQdRtu65tqUxiZAv8IV1/tokTcaTJ0nMLET3fBgac6cyEfheyfzlmDQkAGRkjud4BtWpaE
JUi0qWMP190aST+fRtQKuNkSrrE5lY6Aj3RoyRWZrTSIq/63DQjQQgLF8eokNnvBtReT8fMn8dZX
eNNLvWrYdJHjw0Ner3PQsIRKGcW8p8iVro0V25uWMB2CXzk4SWjdPtpwNgbcSDCzC0gBOZmJbQ6S
c8gSgfiX2iTNPaem6L+VuC6BZc4Y62KuenqtAbZgZ/Hxi4e0IqCmVUo7A8BIHzlhNXKxFTViQYlk
rTGobPfeOgxO4BAGynTIaBwf3dpyr4hSIH7C7fSwFqe3nU73Lw1uher0R6Z/8PQPM1ROvhwt2sW/
Q2CFKfwLKN5RVjoIiMOrj54nCKNrWQVdwz+QuPiCs0CxX3iWJktLf+0RZZZysDfC8IdcD2xU5oWa
xocasmkRHFNRCZ0K9zisNGwKtBbw16mmVZOnTmMDLkQB0lnEZiMRiQN9DQnGe6WwbQceg5cNLxws
9Yl/Uy8AMLk8a/qt/OwJR6RS3HnPzswiUqacxZIeSHu5LVkwwCtP26dsRN5YDsX5MRnNCD2lBVGO
AdQptSd3Hy39A7fgRcV1LLSCpCa31duL9JFhub5BKRBH0VlVCeIMFkciX1rOeiNrYbvQDBQowbqF
lPxRIr/+dxHtHugbNME2/IdwHRC2AsA05howhr9ol0YdRP9ozSLbYs/wb6OctFK/899spmxOfmQB
FauZmKjoo1uWV0vCJGZsvEsctu9yTlji8dft7iC066KtZd0AyfaVIkF9/2mK5+0ogaWVqq8o0Zb1
qrbTP1DtgDTjtzk/xWjJAtSTmUzJpfJP054aG8th1A1vGF66IniynGg4t9erhXYyJic5E8GdIv98
4ccba4/thzqO8wjEn0hI8IFk46CljiQ6DllrJuR+N1MUAaqUVRnRNCZd+6JfhEzoNS/h3rpOYoVT
CrenjpUi6o+4FOP0J2zGCQu8RiA7/BfS0GKIyIsL4LkvMVKo9pt7tRTkD+XI3icxw7ro3GwEiS9Z
znCUSsnxb+Z6h+9bE5mQYlghwifWHELO4AzcppVgXJHP0QT/5GnHvIyJ9E/xo48+h3enyIpghOuL
ToX+842Et38k0VMvYInDiDMbzVfvGfeFE/Abq3hEJpwcfV/6E9GK9J8+uO3ab+4HDriPb3jaAZvL
ncawZf+1gLviQ5d2lHz/Mz+ZT3jcvETWfZ+b3j54qr0XYzGWApQQ5hF8lJJaTJT++pkJ7DVgHDb3
UFCqL3CF5zVwSuO9WfdyDhVfpnCVwVBtNVhR03wsxmsCz4FcBm3PgbJTga9ujIiNUtKtocXYm709
tRCT/I4scgCgd94uq+areKPTpE+iK1sAY5woIcf7+7oRQzEQ0+VFW4lIlhZQXVtDzXfxPzpaMPYn
PyWNhnERfANNC2Yy27lGW/s8szBuMFoAD+YYWQctdHbcfud2C1V9EdCcwx4kbjFX3l2makKrd89l
OolSg7Nmm7tGfk6mlm+4cBbrFyAPLZ3Y/xyjE/EcMhqLsMPNft9CytXPEhQzJFclOuH6mmLGWGj9
lzQ2JV5hGFTwenIhQRDtxE7WyBEl+HJEdX6G+vaqxlYbzafQQRdWAdx81eNHYf0jQoqspY/6a4XT
Cw5a/S4mKvZFO4rpAzAzvhRQLExvX5jj3d2dUHEsEExp/lIbojLeXi+ObkZF9nuk7k6HnuOJthKq
3Nrv39DLGQUJv5WsR/ZAspKisDao6W6dvdPV+7M2RXIUnGvoWuupuEnwS7EP0vLHx26Uoi5koAe0
wQfOAdItkzn8XY/deawHkJWOfF8VxZ4o3tLPwYe3mmSxZASTR8bXA+e+RwYumyjQDjrBHAnIKfwF
UZAsCznIIeGEpKZNotJ32jawQSZVxTJxbrZs5kYZbIX2TymDz+xzgyU+3fFN0ONmi+Q4CaFVG4Lx
F6lZxf4pHQPUlVYRHuEW6mOfB4E9iliXplbkzzouVheGyTumr9giK08q1IyKvQIyoitKb2U8aCqi
ZtvnHll/OWryshuWcsMB/Xbi9hzuoEtUdKqe753oEqHdzXl73Pg8pPhK9d41CpiWz3C/dBEWbulR
CBAND4MZFu76TRG6j5iP24VVxksfICHULpnfzIGW8LkpwleyVDnvzX2JUx+K+8+xX44Q/bBhsQ0J
nsMM3CFXOjOlZnNRkHEtmAz7ypqH+g8RZKe2mfkrKTwMZbQB1qZg8owKYqRnOifgTRD1fGPwfMwD
QYfJLl6en8cLs+S+y8H8rVZiG3CuSgFsucQAXN60GqGNG13NTq6ANFMKT6vX2GUMU4lFGQ4qWgzb
R0bqcI/NBAZxQXGSY6D2RcFR7iJ1YQHuGS91MYMQx0ruBTBefYjs/P7ZVRbrHjuwJNMjR0NuWEJA
Z9R8W8/oPf7eRKhymlKAyAhihhAnd59yXsSPLUkhRPc/SSzRW011+/2k5u9UquGqRb9kGZDqzDB0
00MIXvYOcu1zWsiXg9TXr6ZI3JBd7IstZizkIyBdJDLx7H6jGNaAiKhYDVJ7ZgpakAHbGDryeP1V
XeSu5H5/FyiXoC4IH05JfXWDyr8GHRrH4RALKA5chEFPvKx+UUbrjvPIe2wd3LzQfyFMxUHrALOd
wI6SD4Sdc+cXHWQ01HxiQl2MikN+H/l+XX5oJ/FWvfOoeRki8a3LQ4c7ZZswoBDtwxNTA7hbnEDJ
WyNEZTkiiCL++rVebOpFKOWuTIs385UOBD7Hl/DwHOIlehRArhshyqv7caIqdOmoTC2LhhylNgIg
l54aQHtbIL+09S1FzKfWloHHgaRLOEuFfGw2+07IwfotIB31jrlhLD9sSmUxPVYYuORhacCsxCPv
RupFulYf7u/do8rb0iyjqJuGEsD9SeDaHVlOrPUydagJ2SmfQ86IFA1o6DUOS8kEerSS1Wez0URo
NEDYQ+7itzSqTo8YHIyCyMDq/H/n9rhCzhseBqZ1tUUZjbmF8wMU1jV5Gyz1Zg/r+rTgNr8vtdUE
cPmclM99lEIpG+sOQh2RUo89ePUoHLDvQh7X1FVQJ1Aduk6XVCjsNoCcTAuF4Afm3DCYMziDAwSF
fGB86fyqwkjzTZwC3IXysUTrRSE5A2e0OVUPNhZO9sIZP9R3W6BsbCa160g8N8YyIpqGWfWjqnzT
Cgo9FX5Or7uWecsyPqhHEVDHMHENueDkQaCkMF4/dQL18hX6gLbFS3jKfuKIrtk1myQyvdbNpHVL
biXSL7ZUBWQaFAItU092vcI4OVCIVBcVxzlv8BHxWf5IjB4qOmjjvTs8sK/99kHN9ACzy5gDb6vJ
IJSVSAbdLIsDOgJeG4k3OhfskowR8TpzzDKrsHA3n5zDHDwcxe2XkhvIf9pHCXDPb45tvJchQLnR
J6ifLIwkOWM4iNAJCbECy3RaWHVzdpu8wLPo6neINuz4JabcgjgASc9s9FijE6hH2bKvONaaUtEG
GkoFta3EDnxmJAC+OpNMWolXp7hJY265IRAWU6gpp/mr+Wzaofs8ajIoH8GkvCMemMaO02UyQrV+
kS/c0c4Lwk/Qk9+zfCEwZ7UrWvg5ll+wjKA1l20yhu7MtGFM0FzDQ1w/t0qZC2KiASKgyZyqTbZR
FC1PhDxlN8eJMcYh/9P3yXOLLMsoWIAssI7i2EZGWuxo5q5fu1FYZd/fDE5YFb20NyV95OJG9GmY
Fd+9JsNdpXNgE2smcrj/U/1i76aHV6j/rZY72thCyhVGbc/Yu1BrXInyoBuapMCMctgtFjlzxomU
HjqqDke1E/H0fjWWoyPg43/bUmelT9kCU7tijsif6BHKlOzoIj2L8U3A9+4mezcKLe3pB+3qnIif
hGnl0AQ8hpSnQKA67Waa4iA5oFowZSuVFvsXg+gigwLDl01vV90zFz6ujp8wg4QtSb4TgUcksMi2
S5auXXBAQy4Ld1d6hqwrrBvZfJAYHaeWIdJDC2Ps85gXddKTTIye4cRPM7/FeKr2Lq+qRKJKJAH0
znAkZzWEh5XCcbD8o3CVCiOK7wRXrfoWTtSg/JHOXU1dHhe5Gm27lM/b4y8uXXCSgtEvNejBmXCP
wl8f1ElRMLKvJ0LBpzcH+Ez5MbMrjgVlslKSQCTJzUQIibHfBNUsCflGFgUbxbVj6Rzz2kIP3rfj
Gy7ewc2Nk4krXAoyLf0jBV8RvmaBVnqskINPemBM4aAfC1vlosVho9/wE4Kr0Q8ZIFTZDt5uk49U
puhWiHYpHMMzLlVBCLvzQ3PuB5s+wbyq47v2aKxBV4NRLQABpQOjEnXQhwU+Tml5u/OyxgdXO3+M
ZeWeJp+bFmmj0qNbi2SPNB2bU5WzSAMS32VvR0EfjvwhcrC66ZXCrBZcIrxU0p97z0nYsUWNJ+j0
GB9by6wD9s/ssDqQsXzKia9A/dnUByJ05g8GN+E4gKfWmQt8VUROGXeYpxQPhR9iiKKZmDRFfytY
wGZcgldJ+Fpx6hOlVXc/Y1C4P3nB3r/jkJuejVMcXfGxQs/uhQgPWX+2Ut492YjuGDglT3+wxDUL
GhT4xqaZVDUlzSR+DEMUwjjoD976I7u16Zkp3IOiXoj+JbDIHiiHjRMUSBaeucTOAEold0T7Y0oR
75X2PAr9A2aGkk2oAuEwCAq+B7+f6APy2HQKd+agVq3I/N3W/ZkvvleSoB44J2ubOJ5N3WZBw4GY
zDgpsZ1xDPuEJEAzz+CNBUSVTx+1ujJHXnD4k0bT0m3Lnn2he7IkcmxRP8e4cKor2xLoc8bwiP1d
JCoWN6DD1euZI1TaskZ7ueZkC77ccuO6OkIfndhZf40Io1FVD/kYwhLgZspLn+Iu5OPVc/c1sIsc
Uwj4SN9yWCn+dxr96z3mm5mgPL4xlotT2NT56cHmV7QVE3JuLi9IshEaqAw3yf4aWaXbnawSxiJT
BskmV5ZFXzgUO+50quWLtkEZug8dywA1FbThgZzJhV6MvPiznsx4XzmGKIRoczR91UQP/PIUPWtp
GJCz3fhTwCKCKsYO5BsZt/fcM6si6KtT6/chGbNzI018ptSo275fjVEpr71UoSxyQtEagpM7NVXI
WchkiuIR2opwCAi8foR7chl893RC0HFPUdV1yIk+s8vNwufhKbB/UHOm7tHXdX9UFlDWxidxhKsD
mANVBTn2mbu0bGh7wothLOnFrUs5ocjlcGsXgyLnYPhRqrdim75utIwE79Bp9D1ajrXCUolXm9qL
wZCLDRpvEC0hGJuJMdz4h8ysZ7oKxlZb2MRtcoZnekL7YKX2LIG4LB4gO3gEekmnT6sR6DbZrRPa
CsMFtnH2ZiQngf38WN0MwGq+5mjPIAX64ULWESqhzYns00k5RsNVEQFSE98LzCcjH/YZy1yDUoCx
ItiMzqEDtXGEefiR966gfVILLqifj3W497uyML9+ENYZF4V9QGQAy2/KTINxCvFXWAzGxIast3io
DrCTTHOSuqLOwx/o+5uaYNlie/zVfArq3Gz7TOvH5Mn3xe2sGsnnlgtatT3gr4qMagCc118hmH3c
wbDkYII2vEijahjAq+tVN9117GL9Q+X8OpyjXLvg7EtSgU0gX+s9yvcYag8CFNytgbXaH2OsR6oz
FVlyg47iXb7MzpeHxOofVwX/1WUJLFKDs0QNIU34j9Ho/qn3RnDw5b3SgR5K8/MlP3PJ9lVccDNw
9ufmCXWeFoZ9sDvcYY7CSwiSw1Th36yw2SAvBLGXVbRrkwn5Gi/3YH+3GINrtvB6AaJXwf85HzT9
mHJZHzPcL0s0C7Hx5mqYdZYZdqHDEHAPr7agKywelAZAkWUIkD9bN1uZteZtDd5+Q+mS9deDpYim
ED5GRXeMEJ1YgRJ/qEGFl2X21JHXKDpW7iK8DdBqC+DGkdbvCeOwYoJm+Q/csuPZ3xIw2y+9mu1s
Za1UrSvEOpkWgxoQAFeHUPZ97aa61/v2d+h+MNwqJeVb0JzHp5T06wv1a9W6HBUgGWid9CAGUKYQ
VUR4swbkjw1rX1yExHSuFNufCHuhR5DtTLg669K8cjm4HQAmrbfEm2/zxI68a0oThOISW3g0/nVj
ZBrfN3bMyqveWtsyEIZEIv/nB1v5lQpSE8PP/85QCbJpExgDaP8wSQXbxIxfcGBqIPse4pYpMFLd
GWCaPXnDZEHQjcQcg0B7S1qII6eJBA+SkXqYRA/q25ueS+4lxbzjTWgs/RJNAOi9eabXTz2BmDHE
XPT8UZWdNbKo1RccvlF6wcdyAtbVihNA4oDA5hQuC2SbZmpeO+/3/PrdooQrQzS9qXQU88zAF1z4
YaYwhIePstkjEm6W+BFtU7r0oI2IHU251sgqgXWgg1kNSiQDfileTG6tNES/ZA6uqSjJWHfiAvPl
m8SrrxCiVKgBDjwgOWUpt0c61cXXRmplc6JXbWlG7OmGXPs0bG6MJYtcJdUYClUS+FQBMHZfY3Mw
6XYQ9pFuwmVhcNTv4eF0tnN5ftaREhVFS2Ou6LJT9bhMXnX3lS8aSXUhNbv/P2DIal1VNGCOE8Sm
+sVf57GGr7ZyCMYMI69x8G5M4Cf8lFHoqKEsVQyQyfG3FelmBbfmXyKgUjic9acCuIU8V0W+rWsO
A8pHem8ateyveSED7B9AsDutyExXo3hz/+ZCINkKxxzIKhKt/i9UjgziM8vYUlSW7wZqzhAvbsx6
Ur60zzEoNo79G2OHjA3b43NsrOzugufH85Ov76ZpkxzRYgOTAqVecqQUrlM1fbSdNWdebAc3tLVC
iVyAf/vI7TKXX9WnVy4pvk8CqhG7Ybvve9c9W8ijRc77W5n+2cmYOTp4lssjFlj0mwiUuNjd3vqZ
K8qOGr5J5Evm+Ax6LNbQ+0keUwywsU4xRVWbEUfMMOagxzaTOLgDU9L2Ea10J5GBg0xuelgmc33K
NC0ogxblp5yhBBjGqD9shx55nInqwJF0AvzZvk1TeuyAPTSF1ZEAAQJYFBznGFcjOufKxdavWY2l
qtjFOeR/E6DV5rBCzUhFwBCKsOFC+diMkBLfQ0vE52pBKxAIOKaUse78Uqthy/IVCWIAhS1GBnfF
q2r8NQkh9J/U2TzGqAOD0DVLf+jRcY4rSjuHMGWCKp2SYRBOhUIgEYPcHaE7wISNVNfU8yrzzofN
XCBji08hkhkbMvsD9rFrRKwpqEU7nqMwDXvfQ5CaHjWUm46TlMFw2+EsEfMlS36K3UkG93zqDDc7
N9dUqaPQ5gcP/nHut6gAokmMm/LjyrBPvZB9vpu5ks1/49UOkWmWUIQFV2LHrZQLudbGEK5vPPIk
A6BnIWrDFshoWKbO3KZEC7uOD1AuwSqopUnrRSRPHO1e640xvvAuE57g3S80DEyP+4i/Ud01tUbM
YUXfj5lourMhILFUq1faZdTc8OEb78pzQ5LjnmnMNgazoUJ2KUdn7GyBr9fyLc+BQPQIYe0rrQLZ
fgSb6kBKbs9H08Os2Uk6dj+xg+YJeER7qz6/v7CcFU9Yflsg1ETKreorP8iRuPC8U2lA5yyTgpLD
Q8Wep5tl3pI0k2cySAXt/AyLW/HNIzxslL0qK/e5pF/l94GH8H4xdii6KUDFrDVqc9uK4o2IVNul
FmEWnh7cvMiyrPkVPkH5cn48lo9LwIPdwNNPspZzjqETH5S1/49JQqetH28p15wL+CklTZYByYCU
eW0V4CKYZ8V+3dDZeugmSfTVKnYovvOerg3ZNpul0GoNBmuA2QFJ7SnHi4Rw3bYtp791n4c5+7Vr
3UMqA0msTRIFZa9vDG/DqASuzMV6Wh3awnwcnCN6TjGddUGKf9rO3jQD+O7us1aycpy3F0I/gFgl
YMhaE1VzhRaQQ2DEjc5xJ+SgPf5H6EDmW5dhcbJSGWyQhdIRMMI/FUAkTwVHGHnnm2m8x1KX6DE2
9uYG0Kz4qasGMBhtpCW0mSWTSEnv6tEDsP4uv+PQWmbKFSpnJ6qljwuqE7TgNzBMJy69ZZN84FbE
afxm5zEuOeRR4XLGWNNr+rZ2KRdpP6w6bhqy7QRS6njosSnLOLk8EW4hEI3ubvxwd2j4V8vwD7K4
rxu9p8TsgtsvebdI0TSLOiUAq2T208Ovii1GfgBJ0OhxExo0tXR86zuEcgotoSMVpDalnSC+0TWT
AcsIxU0J9tB0dBvcFHrpXT2403ECM73J5HWamaIrXIHvv7sjxd/WQz1rc9+mJhArxbiV3O/ZU8nr
v5fxJ/iTPJ10WPFJpT6UAQ/HbFsRtWuqKR0zbuu2uTmcy9N2HRsKv7b+yffnFjnp7EFFOx1IMZVc
54B4xpVrx8GKjBLXECcFbyJ1a0av/90v3ascOv9VTGICSHYJNa8f7DqnGoyypaL45Zg62QcnkYa2
1aN7jlbxuVfSIV1V75Jb0MDeat+/OTQXPNH5oIGnfwfUqjWlAfmSEeeB/dU+sFJUdGfRRJ662wZs
wz9OghEbv8tjlpJjq9ysbm9bTYjL6T3DsOxndT3M69efkVHz1xpBsD244EaPuIBLXNi8mEQnlNFb
X7LU4Z5BlsDoh1FmZOF9EZ+GB/+/TY4Qz0pfor3jimqdoQd9oSm2SV0SXOYm6MfrRRqoUx6F0tln
dWmRaatB8wHx8APixpr70CBgZuoEjYH3vbkuTOJCCybmUQDEpegRbC7v65cORuW5QTQXwMOts5WS
cX7g0rNo9hxzU1mS6v3+Mmf0WUV429+XF5Zwj3kC8C1ku7UHvHaww/FMQmCvs9lUDDdWpUEGXTvc
87LuS5rUqiXEx3i+d9TvOFIiPZpnUrxjLQxJERMTmZ3lUQeQS1pmeC9RCMPtErw11mD46lDA1277
aM6RW7DPR/CgmexpzpV5/ZuDsc/g+LDRSwG4uNhx2BjfNl/vuNXs95Zua3qJZfcl7BE30l1F2snc
RGFwzvl5NOctZU6Kc60AHYaH5OZltVNSBTnl+xW52U71X++a/gqE3m3uQ0LRiYFmvJIMCvyMeUhW
j42GFJSSvPgew/81F7T+w3C0TtNI71+BDcqYPGPbFcqQcoT0Fqz93Cwv8pSVusIDk183VuLhtapu
lWRqNwss8wUGNXdFMUM1r4AnGS9DKYHoYG4F1Rh5H5KOK8ti+nhgGNHOjmbtihkkLXIAMYLHQzlX
kwwXR8P6g++6EYnfa2FYGMhmSaDcWSaL7EaKWoZYtdKKkZZ48lzm5ISL3ZcKrKczqZN/ovc2Ia7m
zf1GBfgybSEtqGsD1OtUIymvVk11iiPXaqNOsU9hPBvhXp4Bv5Z5v9EEbZKmHVOKKF9fBu/9PFfN
RThtnfmHQ+fX96V+ehVWMtD6xCEgIAN+aa6vS+gi+7qa2B+dOQgzqGJph9isHC15qJ/UfrG39d5h
CQ+Klk3qFn71QtHEqgQTFyhl4iAKApTKobA3X8W2lPVpwxuqUYwCx0EQmcn15dOyeHRQpBkpPBWc
ITL+ODc83S3CCRHKROHZT+2/4K+qfAw4osE33GdSX31oHwvZuGppvuE1KxxjNiOucbQ0R84aqqqn
NOh6lPSDnSNBWhHIh/XpyhunT+JG2btfRquy8/MPLyY5RSDYuScBazz9SAuoGMXgV8bSDTau5DaS
fnQXO5Hlx4CACykYEDYlhNNcCt6/jM3DOQ6IxlGzWHYngB0YcLXxeJNQbyF8LB2jF0w8wJlNaG8V
8Qm9HwEA0VOFXQpNQUIexNDrCT+C79i3/RFWk21T0Xb8dKXIDSuPsUs4QtjpCYvTStX10j3n2WE7
3BE/QZIcDZR3z+VdYGgTEwHHZpZMM0zG8anMq7mqjUNYpYZFGHklqDzKVBNx1CxSsyRMAVkR8/Dy
/BNHbLBM5K5OXKS+YbClLye76hlOOqGttg/0xtpkGmm+/mkyenIi1u+kWwWW2Qf+Tk8w3zso52QC
+dcXGBeu5bOuJbIqeEz+EOGJkmqs63mMeHdumd7LjoAJohivRM3HvUKm1QyhcpIbGij+UDVabsiK
VBjDOfyC5DQdoMFwO+0fkO7I15SCBmnmBSyYdU4ffcwmOvZkihCstdnlM8tVuqF/g1OdETZDouhJ
Gw2bnywjBsUHZIlXK/BN/ouN8bi4pLRR34EhTcG7gVig4mgs6KfMhB+X6MnyX00eEQOOBUFoHIgL
68qKRxb4qofonRseFhYhr1lc5X4ZcmOJ49KOCh3wfDU9v7sgyJToAs2cEb5JMXi3F6gfAoXr2IEo
8YHIrhJ2oTF8CqkJJ0mgxZ9CP7aLjbnS2o2qu3X3DjVr7xMKlMuhYNcce6Hb3UUzffTmXQZXfcQl
9OzQOZTh5AEYVus/RwKKHRpwoZQaQp6Bvps2dacIM8aJ8dHgywb3Tg3pZLf4mvoNuUbm5+zSX+MR
5oAmN04L6k2qfIpJpbXrCQXVS7+PAWo2sb9WhqzkRwvGB+z0mSbzLOmYG9U9MrEEWtFxvreGviet
U0TLhdAaTcM3PlFh+/OW+b52yH4cYAy/DcOAtE5bMqGpTzAw6HY66wOnYqAusCyZDYBGpGszeyyy
ZRh9AE3TjVK1a4Yb7TuS5iMMiHpFb/0ArPcg/w8WLGZHNMq9rPZtjtu0X9NQ6QljIUHqnSf/ye6c
ryAqNed3iU1oJYOg8AuXWYQbQ8UX8Z7Gy/MUyQPTXOjQWYSiB+ZjOTu0suaAQYcvlk0VMNL9b5P4
lgYg+1I8WYxuTJLRUrCpnwCFyVKWNIFRzZ8S9bWifzKpFGfj2AYBuXHF3qRSqYSEMSSiAtgxrZrL
c+OJSpmF37q3hvyF1yR8uVsd9sXooLXkl+vS+caa8cdSDgZDMgt2xpWK4bX9NqnkTM3vyasWvkfE
BUPemI9arUtvRRSoHdJmBAtIs1Tl6SG9jUFiPf+nhKq0y4IZIi3kqJCgED4V48VH7MJILp1x3BIL
amDr8AfBe25I4TtEDKSC8MTLU3zptAOA5eX/GGANCnJ7ftoQISeod1z5XD0mDXKG8JTVCzxEi7Mr
k33nB9x7kB4/+TnA5pXTYeXDlqdHWhlorTfIMrS4n6gW48AIkgKp88v9Gzw0F4nuSWD32yjZgFKN
vunUI7HAeajOtftDjdnmJ06pmtxXjnVb/PrPQFO72Ei21MZkkofBDtbSD33MMHh4lcxwzkaE7Y8c
MequI4PhgxE2KIrMNaB6/LFL0AVl+xzAKNUhaTcFcM54MtERVeHBQiKldz/9yecNevMNdUMoNJra
OVWA26D99Ymu5AzB3M9AcOrIQc4ctC/nQQEku4WLEZt+/scxamlrbPK8ATXnxyTPCkPRwk2EsFlh
Mz6cD4ekG/hHkTz7bv9v55zSjzpnmDAidkaXKj+IfBtuYBc8Eqtd2faKqymSkShyyXrKzpVKuwbR
Qqgya0BNo42UziflfKsrqUkCOqPw4dri7ZVy2a44ndfwMlg+oEJlRs9S431WH71t/W3S7oxL+S4y
QGPcqojJv9N2JBH0PgkMYH9gozIevjdMYBUTqyBcXmk3gydRnczkDDIC/YUV/Fvruk6nMiEK+ft+
+swKr4EAsMj6aZHCpnO4NxDyizpF9hAPVP11jsls8kgmqb8dx9TjiekWBD6kJNWFkQ/CPSd46wPi
GKl3J/76Pm3L720oOaxiPHi7DKQp7fGFHiDSP2kpHGr0R58yvveG+/T3Q69QsgdWq8jZlBBjfvey
Z3TNjEEI8l/cOiRyQwLdCq7qjmJatgPcD8ZdYUeIsIIENQkhzKd65CpzHFYXYJXzFgMZBI8NexTB
AifBH2+93L2HFs/BbMwG14x7rTgqw5kGYKw5HJKhZ9NcPUOWK/dJlxXwqzCrG7BvKycu+fNyI+8F
Fb12etwTdPukdzMZiqpbO+bj3fd4SwaddVQ541WdN4AKk7nbsziLhI5kxNffod5kqB3ffC0Lrr6P
Z30pL0dB7sIusbLblyav0l8MxXfUlNkPLCGUGpZKEBgYPLc0SBLbIeIML8k9UeoT2hCmtZFnbOSF
MIYiU8s4QifIFTORpK0cYOwx4OnMTf+b4hrVYhNajECYqUAYlX1V4Cu/oG9G4aF710WizptrAEdu
o1MdkPn2HTsga4BlFqjsiTjrhjepQ95EkglUwO6pmeYT3xjzj2xRmCmgTvSWBIIK2A4qIHvp8Xp3
F4T0Wz8PAA8qXsgvvGy9Ex61qH3rJMcOFOMqawZJfdz4aa2booN+jn2XNlhsHVHaAZtef4rVXfgl
QmRQTg9gbWI3IPOL9tZhnfEgJfaHtK/B3aPu+i5JvTG42WDqwJLIOYjC+5cJs2/No8xkyQ6qXoiL
8znbeOIkNsFaoKxHvs3w7jQeoKPQ521X+Cfpt3oluX0Lb5Ti18Vt5kJ0QWijKRKV0Qbo04W7EXuU
Pwhpercwd3aUO8AE5ohlR7AWwS20RwGd8P65s+hb9N29U4FbKD07Ng08vSJ5IATwVUCKWtADr2FL
Q6mLT2JyaaY8UsT4z/YqhOE7e5PKrc72AuXHqfPv+Ssr/wi8k5TqjWg11FXGR416yNGzP26uTqWe
XPKNDBdz4rOBObmIov2JGlIcCOO8KmXAFB2dsiGZnJHbwZMXvMPjtHkbyidbneC1uZIz6UXwRqBO
ePmBUpGvR6tij3QjreX9nHj0ARiGNoRdmpJdXCcXSBiLEWOjyWMFthrpmD9wXiS3UpQFls7h15Rq
HpIonoeYYX8opS3BbRb5UdM7lGy5ALeMSuj9MgVKjR4l9NwCkjS36OFQhR7vd0p41iC/895FQOOe
QOoUHrAa832CG5KqZwGLbkrUyXeFftugrg7bkK/XnkEH+uHuyzCOHnat3G/EQERBkj/K2IsEBgT6
aVWvN5JsMNsMVEMsNoF9FBkDINL/9RB/88fVLdP1e2Y1bBD280Iq54baABmNDDoWUCTw7TsUHBWV
dVIoV+wSGxj0jeOawegAAIblQUlTEu6KRPNkJtz1q51goVWDOxrs9M7fRe8vGrR1DNadD3wg5mPr
OeNbvGwVpnJvA1eC4/XpPRN+iaU206FLdwCX0PZDfF1k1gaJUJ3YcT52dRbBpsj782CDmVVSZeMZ
tM86M2ZvULHWz0P8EIWB9vejCTama2FPNi26IYDhf7LxB3HBAfZX3Iu80dA0ThV6f/YduldXvjuT
9SK22zRvJ1lKO964Og/g3JA/smtPHLuDUuT1GovlV/RtBTTpS2wbUtjtqmMVkSZ9dkF1Rk59xBCx
GHJNLxNlPHXl+p1qBeN8XaUCePgTgsGgO4CrVG3Lg3S4rPX5GPOlTguFRivM88lBimQ53mRZT9F7
e3H9OBpMqs/jCVacivaE9/SkCijFt2kdHhJJQSDde647miSJE0nUB7gAUzQWBMuWDvyS5MVqOZet
gt/v7m8WMAxGGmDD56SrVOgfArUs8Eum/5gM/jUxbkPgdjoaL9XqxLNX+GQGqK+EaGj6/G1hVasK
WuV4/SC/F7NclNWjXufbpitm8+9B6Zd2akiE78LUffrIWPivqZwXbPr9YalY9oNp5CbX23UDE15T
ms9rOGn2K4iDa6EFNquEAL/0ZhFeUqhIoMkTWCTTBJ+5HTDUzkwpPgx82LiC+NXUCCyDXkZnkLAu
giNzxJTxrJjBgycIM0E39Wf217a6vj49yviiIacQeOw0Xg+/jeFj6V/p58y3L/Dykna/We/b9I0D
4xw59mxm85lFiuVopkAJPTMjuFrfbOatHMi2S1wmGwu6FNTi+LcDBz9Lnk91R1S9BLDT1XGxONGw
PIrloZ52h9DSnSLN1WZHa35pgYw7HDzHfNtkCsOPzsqar462lywfYA6ONVJTRh+T4D71SRUSG8pJ
ktHi/uw033o8zmcOlTEMzp6LAI4pwXj9L3/UYcPBqLzY3yfOx726nLdwzL9Nz7Q/XAPGcUYid3T5
R2hhCbvJlqEy/Wv1A9J2YWYDcly/B3gg7PUkGBf2lsmgwqx+65KA6XYgR+Vb2C44P00wR1/a9e0G
c0kffEgLswQykHGgt2YZE4gllTFvJxE98ydoxV0SsmotF7AbcWt83TXddDkrRyscAT1KbzdEgG/T
NdZnOYcefkJW1q8yvIOmj5+8f2Frt/DRUwS+ch0t0vZef7mx8MP6ODSQFckfONBavNiF8Nj5l7hx
i3LCBHNn/+TCGM7c0fRng5GlwqCdE+E1S750kyWn7K1VVN4ZwCyMd/Q6Ov4UwF2LmUq6L1pxFmb5
1Y6N4CkBes6zbjvPZqzA8t/wvZwac7OsHN1SiTJW4HS5BIpXyRACymvCaf+d/YR0wD7aCDXN8P7C
326/2Ql4s74wKfK/2X2aQX01jbB5XWpOuzV7kYeUMc+RXaZm08AAxwsAKTb42MBzf2Gx6TMC9A6p
jdin3NrcDShXO2rVY891tQaCsGuP2lPmRlyWPsRXZsNVA9Yu2iXir5TxdMrHjqNNKox9+2EGNGkq
ummx+Lm/7epQcYwMtLKtLEbDKfW9INWT7SkCM1KUEiBo0FEzbnzUpl/Vw23N/4SfCY8AInhnf3+s
AJFWAIuPB1FE/V5iaWI/mBwz7YsJJ17rTkNEI4rlylPNUc7kxuIuJY3PJQcqXpLzyhfWwlb22huv
I6U16H2Vi5zfN6QKSwCO+vNattQ2J/EiWHFrr+P34zVXIysZ61iqRE+gjPIz8PkH35oTHWDUUBnR
Dk/c1Ztr4Oiwrz96ClpDSgZeUO5xKYnNIP+Ivc1REpQbpyAk1Bc8CpG25nXrX6oisDC4dVW17hqf
e1eluNqBo/Cf1Tu/pjO/UUhvVmGr9mP9eId0py/Qe+pujmQYqGfgOZHWnEPsmFc/WWvJ1CWl4HZJ
2hF+Jc4VDSNl1dRKzB5oCnLMrwe4CLoQNbRXLvVDIBIVOWB3Gq7DNEnVuVa8zyQaobiw08Yh6HWx
9GRi7WzT7HoIV5GhbpK/DH/Drd74vO3P8qP6lDGRw9KFUj54msrNdc03wabZoGdVcQdO6JQjNeB+
fG/LUI0C4zhZnssZK5hc6Snj3fevUzkM+nJioqaMZ35esrG9VCm2xRdUiMibOLJ0BbYFgMB1SgEc
Y17ppY/+xZ3xzJBe6qRy6t2Maxelqt3b7VxiwI0YjaaKo/BmAafRYm+U2m1hI4Uay3gGqocROf/A
6uDNKf0ZQ9Vfe9PU2mFHBoyseSp+HhOaPG4wmLVU59YEKwhmXtQof8ep2IkTTpbZpG36K5BnTGV1
oH6RdaSK32xbLBRXhi83C2en+dRyrmKmLyUlUDNeG31sQ6cgFWCuFxVR93d8SxI3dm6UmfP1DdHo
vkqa9KWkTol+X/HANhv9oAu7+iKP4LzIqpbnuzBOYiVkgZxpYG/ViDBOq6ZEH4jT719lkOaLWdfg
2zQt+dpiAxmUPA5d9qguXg01BOFneBHIM/X6guHj0a5fxvs11AqP6fNb+l5gT+SJ8IEXX3n7J2/1
3zak9TtMLJ/Uw9xUCeXMAKWdlVlXyl8XdNe+BsrW1KIoB2LJ5nQSJHeGt2PAtT1zt/SgHBeEAt2X
s4C0HdjPhS2e2ix9BhWr0aBPU5H3Fbo61OTy30KOK2pLRcKDBSGagdv1FB8R5XI46RHBif3ZSdvx
DdnE9ivyoLtHt8ZCqDnWKSazOvO8V27WXC5DLX/Bpm+OB/4Mr1AZKSCEBhjEI+rCg1i3bVYY1WRD
PR7Gm9RPQ9smUgVAn/ImoSNXtg+OFZj5lmfclS54/gSlBqeSNPT17wvXy2356ARcc5N7yD4S72Xg
f2Xl4xK7Jdete6EA1o4lYgqE7mkOwMfN1RVsvfPznA/1tBQ4PTrdCFlVcmIMgNKx49s/y5aTkkX/
+Z+GfhG+RuYK54wQocTE8klyxE9QmrCwrkXznIBqbmaqNvNjTpoe5Jz7YBQtFaovJIq2KEgU2ARg
w+bwcccR+rk+SCflUMwujyfxTf5TDoDUBx0ByJZKDN7rTrQXu3dD98zjD/bvtLQxDsdeZW3PD4jV
+Al+XmjMNV8uCkByWbWxcP0ye7x27llSPgyX4gJBDZiiAOGC4OQEHTfv5hrm9lbNhnBTIeMA9q+w
Za9GJ2jves5ik9FbHZY12fTprpx1sYjaViWPZa0+y1DhL2RLypEbd0UXxzfD0TBPL0cOxNghjxNh
rKWSVlyTb/NNGO8uUPoOMQ2XnH+kftC61H0Ek17P8SBjkhI5NVVhIv0ROuwru1uQ1SNjoG89NL6e
/KEIb/gRTv6RkMsC2vJamMrXiNN/uUbJNr6rD671I/TFOf+s9megT3iO5DeLPJGvYQ1l67i2pdlY
9tfE3x5yhJ81kbgNrD6f0QaHfXCIj1tIcep1/+dFsgMG56MPQp59nimM0DUwmN2RpRa5DDXJpj5j
WwVJpN95+gmTYQVHJHJD8WXQZgKBngKtRoQqEaGyMrnfaIL6yT8K8gTqF/ckuZGXY34Pvd2Grom1
J99q59Nnq8Ha9UE+8QMGhRlaVx7kzbNoRSK7kfzj21QKIV1BGOPegCqcYpu0p1E55wVns455uFQ+
cgwmGsgkB2nptOlf8OiR1QR/kyqC/dGASr4wh1jLYLjaILzFg7JrBTKZBGS/Hjo3GGvC8edk0dmz
xJ40pAvxn3FZFowoDxnQFtSWtJvS1zu8dKRN+U4D8+YdY8Ynk0ri9duYvcmYVe/phNkTV8eoBDPJ
rBvOS9FgqyQUpm3lhIvnOeVBm4xAFNu38um117SHuuwdVcQKpt/RuvPEis7Gsi1Qdl3Sfpbaw1UV
41zHtpYIzlCHgURqrEfTjcy+pkrM9W17hf0gJmGB6XUDy312WAXvBa85exHp5eWYYzUHMj6NtslG
3CDQ7UjmUNmF7NBK/RnCPNqaC6m+g5kFg0bFmoGQWZD7fDmLZCXTwigwffie6CIQsy6f/oQ1Ma46
HDfBr4lp+Tiw16wa0VeYocj5SrNAa6nABLFU25Li9quV16NLJCP8swWxyL6tQSTvAIfiipdzSEA4
bfkrEG5rI8vE2IfR87/puUlx853l4rTw8f+tEUfz5PuBCeBpMk87Ib9gS0l+ppU8/acuUh6EjHbP
uBvU7ul0iBg78QZ/wEys/BnGp4YmElfZa7hq46Ac9PlS7D4f0Kui6ZJN6QZGv+Vrd5jSM426VUYe
JINUz/8QHtPFBvDIj01hf8W+aOtDbxmz76JbJjsizPoPV4UvmNYUvF3Bg1GcnmpnM0jp2ykZdaq6
A7OdptJyBHo7rB12dXJnRMPUwsXgF0ylDp0hq2b+lLq6yya3BUtCcuXwWbBj+XOikEr+fW/OH/zt
UiPS0VIsXEWeH+fxkCvN+W4+GIWerZ+fcYWryJ9UDMuZlQVvlRV4sOHvM/upHm2zatrbYpNcXGum
G2DHVrKReu9UgSBjycwdUdqucpvd7B9RYHkRhZwjRuf8xS9Jm0liilEU26tX+X+qwmyeNZ/cDqdM
85L0QR8M1mRd37RRNDkwz4thwpbqB88fYdszipWNHfCwdBehG8PcMkoZeWEt5T614nzO1e9+/kzl
DeZnGR2Aa7yvUD9F7cLP+Dpy/R9mpJ0BHKkZe4v5bvzvZMpIwdDvBLwRR8OgcjHQ2+4TAlIF4ThY
cw2+6j270lwKVJ0rO/7MRSjh2OoovUAL/BqJ3ikKuTZsxxsqILk+z84ycmBrRaR650FkdxEmBR3p
tcMLSZQG3uYwtRLw0gLEiDMVjYNadDLeg/hrBqJDpj7MmkpCEXZ77OP+3lF3P6sSqEG4H7M2NEBd
WHuWfEz16FZV2mshQKgbHLR01QgHXTldQLnbvqxJwrlYyBpD20jQ4oM38VgtWCIPkQG+8pzB1jgN
65s4oTrqtWfWpf7n/ktW2pYM7gM6ah74sujjpwC8w5pAXV7I8HaHGem/htwjJjk5xH28ijbYW+MG
OvD9yp6q6duj/GcmnaPGSfdNTrg+Z8rg+3smeXGc71Nv43hFvQS2L4NLcf1j96maS2taRpaLk2mF
SRUPKrdhi4FZ6Jymo9n151jau/z3R294DgGm71V5lrpR5ljGEFtHHLUIp6Dp1Gg6I5WKrwjy1D4n
rUppXgcNWRv93MQbyo26MydAgl8VBEcVh9T+uKuzvev633OpN7KyIFvHmoqJur3TnVLzKn/1PCDH
HCbUQ8xmupGbSUzW385aBhhlgIWdKEs5T7QmPoWJ0xcAZVLQyyUaN8pBsT56xXsi1Yxg3wulFoq0
LeY+DOeRMdwzP4f3L0CZUzVdQ7ZRcynzWK+eEdHAlcWd8FOcTaVTFEXYc6bVqBk+SXELtpmDqwOY
z/4sd8U/g8aXQk8ghV7YtNINLXP2Jy269kpp+M9N11X5oGOfwm3qcqQmPBgBG//Yhio29LvDCWM7
cuhugr95WAEaTH1iFZRFtrEd+OKNqE1TLxHYHAIeNmmQiWR3hVhHNf+xMdZ7bY3ia474vTA/nTvU
bSlce7eOCFNb4apea4SWe23Z4S+Ou9/iN394nCvP8FP8JM/qzQMQKjLS0sJ44b6m0MLL7Oy+QMbi
OvS31udLw+SkZC7DjFdZDSS5MUulANTsvGVsaNC9dH8+7RZgmgJ32zYrb+1daHuuCcd+cVdeKWd6
nA36xT3ePSwrTXWCYrevFd0Bs/XibHdwDIUNMjSw4UdUzHzKE48yZ5UNYx+1lCFu34NgEITwVVir
O33KWaUHoQHTOjGezt/FWCc/Yfys26i4KSXuomPhl4kxKBPgMX1G3b/ghzebykXBH9UJaH2UnI6r
c3oVEO1rithkwCrejeFYJQQ2PeMbphMeWcSjxV82X8ktknTXouBAEHrFMYKUyXs8Zy6ASO9Rfiq5
A/fvFXC8vQC3TBMDJCg9drUf1MuAp+2HPJJ0OeMIxhkU0pLUHxJ/bfQcB8T7bYXj52+LZ0Ns0HGK
6qxht10ql7TcvVx1QUzUlUrYIkZKtrv90DRUVPisTq+ycK8ETQvGNCewviRnFbuarhijdfRlQy/o
teKFxePUOMXQInzmGmgjX1rRHqtPEJOsv54KEnMP1Q6nlg7zHY7qO6HUDP2+LtbbW83jse7PN4a/
b2wR1sB69utsM0XRDfPLF7QryHQMRHMk/dSjK1kfcUDmewTz6dUXmXN9IF++4bGeBnVdsE+4/APj
mzdvz2F4TCTpvvPVLAt/YEeHglQ+zsjava4aBDM1UNZsByAO6Q3AI2WnqUn7RKqznS9erNiwL8wC
UYricWwmeCvG6Ckq016grlcu0741Z3ZQ2MG9Wg0M9B7gyggSt/RRfrZqzx3wccH5VrexwMTGgdjS
MC7w4YYWyViqX5E7YXn7w93RjsjoJc8J8fecpdOjorfPbn6rMVdwJozG6+nqxlbzWwFrqliWZzKK
RqOTlKl9u9HzeGd5Vm39GzPFtXXilKEo9XbmlvfKaZ1vp25VssKuIAur8u9OxDfEJ25RO7SCZTTh
ayCUNkcAQTdZR7NyOTjK0ns8Ov6Ec/M+jUbnttF2XExRa+peaOAmRuFjOZKqu/sRRv7TBGWmM4x9
EgAU8j+/fqj8BTAMcqyWWBfjm1QxCXzze9I2qW+r6rue0MdlhZTMck+ELBoozkoQCwjYVZMW3JE+
0FNPz1pBvHx/7lIMhQctF3Rdc4V//G4mDNicfDON+JIdv8K61rIPQEzHFKKoMXoj5ZsPqzCbT/G1
6TwDZXhB5GTvFore9m8CUxLTlZXE4Q17tM1/ewY5XDcmlferXVUnLCbpU78sP97Fpu4l2ot387Bn
Vv9Rzo7P91gM6KmqDUqXKG/mquHZddygZLBfyHFCg14vhlWQyIlFDKdp0miR4BrZqck50XTZuGwn
NT/hYr+gH9JpHbjJbOH94blnTQYLEGFWLEJUM/nRkw9w7uMkxDOOUNIK3gmv8+RASHsVWnzUQuis
gpGdNrXUYUVB4mPdGukjm/Wjj3Y0zsRLk/qazfHiDBvb5baGdeUUlOIl/S0cFx1Fwg2uSFSGDi/p
LSyvz1A0KMLptaE/DJXrNhjqDocBJm5+TOYdxdc9UnKLjJb4is9+zx/mlJ6aRUJ7ZUHJ8gfF64yk
jgn0blYvhg9BCx/JrQBFNMvSlKtneoaDgkNAjg2tJ3aLHGId7f+/Bd8Hw8ZkxGlazg2EqN/k4bw7
kiTWbpkMpE/jZ2J9ZoMB2jqMNxAosFsPLupUZhgPbzIz+MDfp8XvzGdKqR+va+SEHzRZ6EDU3sw5
lRd1lYVz+vURVYHRndY15vC6OGmLFRIzXSgaJNDGuToss8C0HBGCisL5hyVRY+V6sKbYa8kyDMJh
6TdSwNLj7aZLsvLrbgp21aSGEMZz7+boMigj8Qib6wUWXmEEJRgjuKo4MIv/8u5LXKY6hrqYkui6
qSGW6WLVpfYhMMxD2FBMD3Fz4Asd/vBLKb4+gN23ZCTR9tAjsvgIwbQbrMTmIO4Qkm+fN3NEluJQ
88lE/Og4tRsWRkOD5O9LSj6dz0Si7bGhB1Oxk5rHyvdhZ2Ndwg2mghF0NUf47esyYOSRXV4Wfyqm
mRliViIvcZGFkJ+Mc53aaqcO1+zjpEZhiwamGyU/L1RQOa9IjQlRDifhGkOarvNp0lijpBEIiVT7
hBKJqboNJCtJfRNmpDHefgcfxWeVCdFMBtKGmtlXPUaAPsD6R2YlVN7UKgPzmLa9Wf9MalDNEEbv
nuSLeR9+++hTDKFeppRI8qTfuwhE2dpDuuFPJYN9SL/rWRvNz199GjhqFbQx55FSDzuNlKcAcd0w
Y+N7OYNyKdMn+1x/vcuoV0NYaXkR4s/Kf+gzO9Sa3PJL8m2bOUGTd+CK4Hpt3E3XB/0Jj3QDBDx1
3w7Sp13qO3rmFhDA+wxiWrAQgvs1XWojzUE4uFar/k77FSmHfZJcRoG3HhW0NlZkjxL9Wgt8WV1v
LiZz8IPZi3FA2nnQjgT6jghXDeWYP8nRAaoU/7mhKbmWqVOBwKCvI/2wbgWt5//xEzW9YIjSKnS6
mWLyffckMf094dzGwv/IXAqP2uhp1BNXxyNZ2k0soFHVw45D8rMFbmIOy5/Q883jtT1bkKnDR5HB
fxbWAiiFsPNx5xJgYQCtiBJdzYbW770uwAw+FBergBPascQl/+waH/r7qgw7NzkxHhj4VN04Q1jZ
crxbprtRlKXRTVl5K4ll1Q34HYrAhoxtlFwmiD/tGGvNCA6yUhcKcre1XB21ig3+ox99Kd4CrwAW
z91BhaLy7D6oojaV6C/4hlJOGN6uOzqvyOkS4N4rY2TzAGANpNkLwiMaDmWLd0lXckDI/7Ckfbxl
KVdBI79t+dp7OpmViS4Jx5YDIAzMn9J1RMMoh5/u/tsiWkCffY7hI2su2D7mVXHbiSkbLlVJxNMh
DmuTBqD9nqVLJU1VZ3TFngoFj/0UBmty9wVdQA6sNEcFHUcFqooIj9wgeWl/2hXUm3r918b+RWR+
pu92qcDdxso+k55RLJS9YrIIY82+OKqz8qTWWeGf0Jns23hJZBsOIIY9t59J9WElN6E4v5eUcqhB
OZUprRCwso8PeYteK1qalgKZI8CDrpHCUiWVNSYor+icmNkK26hUF1/7edkwODBxdciI1ahv+JJL
VuuAIePB/+c300Xu+dV5ufbVJfQsFQqclc/Roxua/8Uz2R0YpaGdZdQIA9KDxwWkk/4eUN9IBdcG
MIg7GkHFTREsLm4M6mQYU1NyqwVANQDmXWwKNTC2VWwi9YVbRYTI6NRg18e8txHB8efH/RSxNpwO
3PcV6MnU9Q7BTXk3lnV2nM+Yh1fMUfAFNhYimWAxi5M3YIb00mi2l68XGW4e5PM6iV34K4xvtCYd
pj1zp72m5pm9JIL/5MxcbDlrvimD4yQF7eUUkpYXFjmw863yff1UQB6lxq1r4GjXvfLnBe9YP4BZ
gNvIQHHyLm+ORJle+GdJfJ1x3BTQLZCE491jY8sAoGDuMhnpD0j/CIJ1oSy/QVK6U9ekx5QgLOhf
q98yOEVu0kTqv+25cBZ6RPwmP3XU1p9Pn/OR61uKfWTHPD0YwoKLTvPTiU0xq54d5R7Smd82Il/x
c/0oNvWKdEQWUfeBxFC+acUi2FXhX0YsiN5u8YiLBKAFm8QjB7el+qhCz1Ih/J63mdWl3PKEjPg3
tIgCygbO9r9BvLpS7otKPLN21Pu/nTGEAP6zBzVqvqtFV3ARAix6//c6xlgV82TCn62bFL449NFV
XUHcPgX7+8SPjJSDj4xNYjZlQ79pugSOFRGZXI1vI1bDA5JbPSNg6Tz2xqFzImm1Rd9Xm2BBu8mx
opEKEt+m9C4D27HtVzV0SEuE+TYpILWkQv7ISoEDLJ5fiEnpvrYYGXWfxnE4wLuOo5tXVWPKpS+/
t6jxlLMfb4f3EuziwWxpLpkaMBXwVU5AItAEot6cQO30mGj/QDX9km306Zbq1fkgKBOYIHmGq/Bm
8iJUIifg46VIycNUD1mbh575K2mUrH/2ydXB40nbBIm82ughLIMx6m5b7d27ArA2fcAb2mGvSMnh
Jlhap3hilJG6EwCqA0yodAaXYIC2ENZFNaVao8JoD7xS+JulfpJHICWQnmgSBGoPPFXZT1AKSmJy
r9/dMVLeqCt+jbLb1ZWYq/ZKVES8OmxnU3FkxtuLrbIrSFdrZopSMjim2v/bDL8RG7i0u20CLqGs
p8Sd+ns0Kaxs7hT7wsE+h62/XoEi0AypS5V9XNwM/wR9xZBKJe7As0Qo34jBazX+THl8NTQGAVSl
tuh0lcqPCvgh62YmvuWKG8fvgENh8bUzEyn2AOWT223d3fiBgq017f7vTUqfZ/Jp1QnuwvoDLc/u
v6bWKR1lc20641WOe2KDtEI77IzGvjr4B/kgxum9dhdtnxI8CHORcLu4VZt9yrGArtpDAz1uLKpT
zL/bxFJG0nVBj8vfwo12GEabgCiUQ/TOH2RCESwIF57C+wj6pFZ+vZPwh32CFGNZ60JB7WNMO21w
kgQJC3nUalVniQF0w41sb4vgnDGGfxCfCJMaIk89FRnZdcubBkCGGeLD/nh29ukKeQeMfIV242j1
E1kRPmS40dgAflxFx3OqUHF1augs1yLKrr1TmxjQ0rkb7NIr2vL5om1UtUtOvaLWrNL6kEUPZ9Ux
qyqFbcEe5Yf/WLwB1bhU5GYKJF2Bkr4iUQwsmHPlntdkKNr/4TjS643vtMkyZ/0B8pZNd1ajd5gi
lO13DrGnIvr2crtfj1vHBCmwN100XEV4gbW7PPOhJk9o+3WjtG8opBmtBgmW9G5MYP/BppKDjzPF
zWywhT5HM3iq+nLMLUKpMcZ1UsLq2OT2aoymx6xJQZvMeEeXaJJlogcdk6t5gwgIZCKCSM9eMTt1
Dbaf0UK8d+YotUzfjnEf6Q3pU9p65irqS/leUkqAfUjVgSDO7HtW7QeOuG+WQPpBCH3ahT7durGS
kRw9KYb8kOMcg2qFI8jZju6nZT/s7dnsAHqipcjHINSmw2JZrqYDq5+Or13kPshy33cnkez5/JZF
35rf8z58iUxQlboXCKXbcVxCp4O7Pw+LkinrPPI1DfWYaI4prj6OHomh46oRejzz4Ujdxxij1bfC
a8b8/2ASgEzFBEI7nbltURvqAnfQU+WC6GXdzXbCkLhLEYRPGW01SUA8A0O+TvFwsC8d1+3+jVBW
/49h2o5eco+xUHU/y8YiMFj+LlgvPApO5o5YHg+XcppV2DDneVQ9H87AS7ZCJITIJ2XZx9rbbuD6
ouP3gTvh/9TnTFI+Yzu6lvk6uTpjfMk6kiNqI5Vas+Ix6jrTREM+UMv0Lr1pEA+jYwfPynOK6PPl
gWbuiPj3OI/P9HHU53CNAqYc/ZPLcre0bijM+A+Omf0NFsqvDgmyyQMgvJiNqHx+Vb2sruH91gDi
9IkzC4ItsPbt72q1Kggqe3o2nStIi3g8ctjtXKt5ZjcE9EgsK5xn+Qq91jwyjtKKc8KcjSqGGUCP
Xn8JWITI5JrVYToEVXv8XnMm39MKOios8uarF86p0cV2X66bGxRoFRK0lbsXCf6MMdGjIXmWpezz
5QbWlbvTHKSCzVX+7/pv2VJ3LLJ7Jtx8QSi1UUE3sppDM18ZXdc5E5Zef9MB01YUpBD6IERFDJn+
dcW+wW+c/uPQiPQmS63ZxzRKWcrIArAJ5ukmqzPxpRxzGa+bIVc8G4L9xz6r7G9MMIbVXRMpcH63
rzvCxukHR34cTqAoSR0urGruvC/ewl3ZhribSGwFVqDudT7y1yuAzfZSTSPXzyhGmEWWGXYHEsp5
vn/ZFd+cg6h4P5kTFQXK42HKUtXt88dDougMBR+5Qg+/SaWR+ReStm2bhZz1zithgun6v3stBx6k
isziS3uhJeTV+6yZtIIl4mFGNKglnhDKn9UhLxnYFFaQn5HTa9V37/FsBTBPrKA5xldcAcHn8Wsx
C4AAXZs/QDBBW6c6YI+MaaUcSb/jE0mgs5eJP4UNHe9ytWuiyd60bpWAkYAIXVMnBx40Mz7IqKTy
vn9qH0PfliTBV1U3RyVn+ZQrfC7MojALJcu7Jrm0GWaAM6EhXkb+D8OD/cvnnER6Pb0R8D9HVLNk
lUbTdrcH738pLGO4Pdbom7xyLbbzZog/gIUgMDxizc2Xt/9flpsQeObxnZ37Q4Fd+JUZKb7qnigE
quPisGzZt/Q5RAUEfwlF3xpbU2kIU25bdm+UDdRDzGpwgkNnodz8fMv5M9/o+3B+nmY9l2Omh6XG
jgwIDEykBBsBqtiziCPibCxFvAXDYoPi20kuJKnlqRc1gevWKxJ8RRH8Fz22cPfuIRdEt+FO4m1a
371I+qT96jbSuA1fKx70LfXVqODO7nuFDp5uKzh67qZeoen9u8wsF/sVf7iJdhdaQYFAIeJuh8bY
9VE+Cz2jxZCeDaiPj75qpYYXHNErCBxveOMQRCDMHrPB8bDkXMJ1/aZ30W/BJWp33e+aOsUUoZVw
uRUEqDherW7ztvv5IxrDOIidnIFXJTGrk0FnG0/BFd1NvuIcSCPeWRQ48CySBYyOZ+adIL0Q2WSQ
svsvHfKoCvspImi1czKYWoo/ARFDWnUn6TJtE0/wwQbvVqmSQX0YWSFrEa0Iu31CClTtZi/bttb4
X8B9BeprgFcdQibr9NLHm+0Ktv6iNLMbITREWan9eH5h1zgG/iPp4FMU3dj7uzHtbUrxf8NOdYxh
+vFd9gYyUZsYnt+cyZGT2xd5GRjvy4d7MaxrRDw1+CwFtallbDkwkTwrT/MvNrJyduRHXEVyn8gf
7chIct9khT8fBN7XiYQV4mT9lb7w/86EnP9lmsjnF4lSQ6FNE3bEFvZTLVEA+FDVC8AkLIeogPVW
jAXpYyhzVEsdTgGuy+yHnwleJwT0Inom1OIdDOnSoGD/61+j3P/zro/2bKERcMQVZ5D7bkBy8V5O
4ZExy5MrzomthzUpa7nBWToGSNR8I7JpRZ/901d5M7vb2AHIQsRK1mI/PKgXnHiIWOL3cjONUPuz
zuoaQXUoCsv9LCHYvKXBMWuhz+e0V/BmZdJloz+ruRSa8YSucmXONxq8nm0NJv0Q9MoAh4bez68q
QghhQQOk31M7K+8NGEp3sw5vvwSZSk5zJXDdW8WjIkhfsXpoY7/veKYAGhTAZlAjK3XzDPki04l+
aYVwUvkkGF1rOhO3IhuTf8RaQ1cRL8BG9li1dQFhbczenmFUcU2aq1/quM+B7l89bOCKAee1CIr9
0k1rUKJh71n6M88Wi2MKCcDWSmICLdbojH1SnpoNFlXL0UgDPuaBpJsMwmx6tDDzyFgmPASz+dDi
ND0WFGYOuLOw/7+Ov75ZuJopdUx6JlpJpNzca3CcfMSVUxNTvag03rH4hfM56aKcOdaEkyux05Uo
jTBo0fdq0Y67cqu9aOineH1YJ2isuxWdDi30Vw5lLjlesPVsuKCJtbwimtY3le3M4SOSq081n3Kr
dJmD43MRttPgH/ebf29+eR9/KayMDzsY1TOsnp2DK3ylB+6pS1kwGyDZ1MmkuLaP3EGYNgYJyBOH
9OraBn6E0833Gqa3evuzIiK4Jf0rRuYvh4juXDMtO7wUx9ujNUy3YH770fFz0D379jlhQMRHlilO
2zKHdoLOtBlN85B7L0hZy3cSivE+56t8Vnc1poU6mxCByQjck71/K6FOELFd+HjtXHzPqX9zhf5S
pXEtU2htboXFhZCtc6lFm9FwdchzUHnznVtak9Mkypa9yZjjFuKQ88yBVIfglPCX3GzDY6VqJE4t
FclOh6RYKJllCnuWxcApZL6KAZY2JoxwhF/dL1eubbKO8C+CbHpXvdO9KA18twIB/dpIt12QGiqL
beZnFNU6A7R5XYDnBXEAxxW1Gg82SlXXVvhVlpq2Cu0BNKz45nYlPWA5yShVpos9Sn24n4d6lWk4
Tei1PpSxoNzWS36Acc6MI+Kgi1g43bjRaM43NRm8R2AM5x5Y47LXO1Be3S2YUX0xCuCHcsSnoNPV
cI/HHTjWcOj6cyDMo+PxgUSydwa4NfyXm4YIWzF09CK4UBCZ+LH+jvNQ986eL4W8eA3ffAZ5d1Vc
ymiP+icZe8wdeL4Zigyk/VuwmiKbgSMSmVveH2Hmywk3OROkoaRAMZxbzCPVeKgYGSsO0GjyRpZi
cy2IC7af2DOx7HxhVvgs3jKXfO1BQ2uQpF2dpOadTBGCDNDSo3LtuP00+20Mnb6lXJDFSSLZ0Q6B
Sm3KfcP2pcAPdsJelcoLnaNjilheG9Cjj2MgKKnSgSWeWHs4WKErOecVYc9xLwOTFMtOpK0EdMjQ
ZGO3rgUFKS9FbHivXYumKdGqIaesYZ9KW6le01LGFAPf7cPx4W+Z1M9MlCfykDf9KAfeS1oo9RoA
obsuhjE+o9Z5vw7hNcSNchngBB2h6PGHDdhfosKVAK4qV2L1c0ZomVdhR+uX3YA+Tpq6LsCS3yi2
Kh0bicmiatAQkG5dpbl7H+oYpjL7xVS/9ZHRKXvtQQy/qT2YZUjnkDR6anqKamf9NIjh1+L22lan
cvhKg59fW9BhCwp7EiJD/QreDpRepGOwOrfotv6S7NdT/W/MttORMgkaDBkg7G0NzrGBMKZlfNA/
YbUkjuGnJUhwaHVvo1uAf9/mtqJ8C70DGdKNCXLrGWdX5X8B6vW3YNdslGgfKrCumt2Dp21E6/Yd
+84XWXpBaJG0XsC3GW8OUMfV10TfLr18fFuJDVBhL8t/vKxW4RLahHIZSJmTJqqNaXELGWuDksu8
zwv9rPauyn/1gw4FZSX6uGwHgWl/hEWkRfMGzXKpuvKIVWA+hC18jB3P/f71A0Ko43+V+yB1EIJz
jci0CDWXCpvVnZwXnYX3RZV1q7UAG4ybt3SBANAdNl6L1aq7LOMB5U6ik90Yl7tnG7ErMAJuoA8x
7DgFbVNnuB0KeKm0qEi5JgHaVCJRy403VVBJIR0pLaAq2Cs11KBqap7nFfh+G/CIHbYe7Lx/qumb
pOYX9nCglMz7GUUzdwD2/ls8VIY8akkkledpPvAl1KuQOg2yPHweg4lpuLdfhswy14keQ1IYowJI
VDkJNSUR7XM5AG82mi6YFdxxtpSdoAqV/D+3+KNI2A0EcwAlfvwVGyjZHFTtDYz1FRyhVucwaSAe
SPUe6imJpDqHfLOg3yIHRT4/T/D4p0efmUxehqyBmPBVLpoOKSP82hvovtuqD2a3ZwoIQtZXm8Lh
GETBbjUmcMkBTdv9kz4KWPsTMyDnbn6/Ht9FqOgc/lsr2BGac9NfLAzXg/bl9YaL65S4Opm8/nVY
J0eXaNDLJAEiXn/Y2FA93I4LsCEqJopP0dDxypaqh3Zya9pez0LDjFcLVsapkrE8hoyFGdrTl0Av
ldyLkfRVTxfbBajvqLtxJU3RY69UpY5GzwgGX0rmIvShCnv9rLA25y5sCBFgcdI9tb+ZyVHXnoa7
FIH0LGDLh7AxPgxjyKtS9tTTnrORHsEbwIoXJSVleAFji+Xk9hVpf/PCc2Zl3jLFVZkZyPPQUU2f
D7dvOqKK58wa279JwQRbrZuFDC9hI1hd7XC0irfnW9rvgi9bxkbZ8ty+X7U8BNLI/usTICeS3MG8
kQzSq8VTFfIi87yDYVDQGVzwcSgEpkMyo80f8sJNzyRbdyaq5T5yfFGncxnfPPNaEdTRA4VyZ/p+
Svfo+YxUJrk3i3ciEDkgfABd2tiCkvwbu3GQfNFd49fFBU6JJuATc0g60yV0kuLQr9gWBEiVfad4
nmmtighxdvCKGtx2Ekee7ExflEjJUeuRLqQl1gAvC7+UMDVsZi1woQANZxi+LYJwoJL2nXFa0hhN
9pYw7H7w1tItZLK7vEKlLANnLvwRoFqMfDR9w+7mBS2o8rY3gcBgMXAfZqNhE0RWEE19mNiXNkuj
HH9amd+ktwunZiFahAp3t1KjemfRwcM4f9aI+FOklZQ/Zc84lb8Hc2g6p9JIdlNWj5L+aelWC4k5
1AwQo9Q7GMVe+eKWjvqBjrwbrC3x09J9M5cpYq2S6LPXLW9vH7HDxv9e655KWTXU/yAnuRyIz2Iy
5IpLsWR7qJSNXIIRayPGpDKGO2PHkGCGjPF4Dy3uQDEmVwaglILflQG7qxUji4kQLvKXQRZVeczG
p9mhJrre7okpR3M0gms13AqqyT1Xjuu0Nt40tnIbvYx++Gake9+ezsqdCdJn5SGVdDJFp1/8eiir
XKiD67PCgIXL4m2lbni9OgKQMksNk9cyjlbjneA05/jNzYMyrjkYjMN/O4tCGn7y66PblmHhirQm
CE4ByxQAOs/1KQmcLL7stLF2nymqOf0KVg5rjPp31rhTMKy4+RkvmuMZxspzQrGx0KY0I9ypUKJ2
XSQVUH2oYMa/wE/zrl9bFZZXa82OuIBPDlZ1qqn+VJbvK8wSHHF6plq9rKm8/ly7Ym6WPuw1yF0X
dLmL9bvQDHtJR1PkQHOBsXHCUvg0tHU3y/3hLfNDtSkhph+0hieB215OtctmOwLNcfhM9e8HbhDR
qjnrWVPfo1+KtXDStGY+evvixZwEwufG+0UiIV2wbRJIow9ZiSYlesq48rtNSWkG8Xho6/sMo0Tu
+k3fOG9yxQrNDUvu2U7TQfpBbjk0GUr75mbF7Pd9ibm5joeovp2GfXVdVRrFu41bn2IRNlOgyVn/
zf6AdClY1c+m4ctptag1j9zF4PaHiaZQL299uFQt3/2ZkM6xuocghRNvHlDky2gZJO2hr/UBMGXU
+fVLX1SCYDuJWa6WcxG8m3NkXg7B19CMdODvEIMqXYEegJFsv47rNhAPguIryRh+nQPegib9Skgz
f1KiMTCFy5ujChEQavT54PLI1mjcH0VvHcZ8c+g7nwQWKGAjY5k8Kr19IvNIMQcZ8+WxxgZY9GoW
sxCFkatCMYfE03rumdMuBFKQ0kBmXA+w+xWIwOP+6bhFmSwnaLUQRdHD9efaYjYqtgStKUWb+inU
aedbQNIfjhf/qHYdN2CvLKCdzMo+aVc/WE1CakB6FOiFbD9wsLBxbVxkh032I/mzLT6fsWPRWMna
IDlEqDlo1X6BjntM+8qgllIxH8F+uCAHXnYdr/S8L8vv0TZV1ucxAjnrgkyuepXJ1ve+fr/drJlB
x/J0mJgUNluNCkjQGXz7zLHychwqajCGvOzcYZgBIME4pxAr1ZcN6Wag0gfAur1VhyxfUESEA61J
K/6I2Z1y84TtPNBk66ptkSZxYFOrGXiYNOjF1ncsQpCN178oFnRMBaPUHT6jLADq3hRkKJcnoV/T
F3VS/0CHcXZiAqke+pjel0TJQw8bY+QUXwJf+E25mPdKP9CRAuZZGseX5cgivS0mOPjWEVLD0MVD
FO9LTmID9VUA70s/MaJ9LJl5migS5ktX2yFeo1vSy0kKLiY9A8NFoA2n3dLbg3Je0XKVYIRz7Mbe
/8ekjqjL7rD3MXQ0RmU+VqxpZ8HZjfJOZDCtmHKvrErEXSXB5//y5Xg9jn3lfWZyAmEQlsqVFWUa
pLdQXM20tHUNIYbUDR5vbNFLc3VuQ69e1/1U1EfBiD25+qATpQ37pVZc/kCGhY8G/OFimd/i4HGy
LitGhkLp+ez4+u/LXwepc+K5VOEpJXCLIkGcIxBMiys+LtXjBTl+AYJUwXAedK75zRZoOkOiVvVW
3vZQN4TSNXzVnRSnDWH8g2MJ1s1LN4Ipu2OLMaPRLW0asas3G4jfiObLGcxj9kMSVQ15aNwQb+tP
U2zIIoyECKLLl7ygKRjUdLjiY3ZkTzlgjT2GNBEis97gqs7u2tsVfasJoFvpJ25VmcW0yJIJ7EOL
QvDJHNU5V1plmayfvyzTSsrlMJHI3ysEikvlad+EhhnWluxYGkGPBAqO0TOID5zAymsPqCStnhPX
/nyQ4W630w8GlOIZI8CDEi0Iy6W8CXc25WRnJfgCrg9+Mgx2QXA69tNp/cHmB+9yujDk+f0H9y1Y
PpIgMmCIKcEW9PKju0N3pn+IAdn9Fd4isI427ZIGn2QOO3L5UUEQpAcQm4VuFs2sHu6BYB5RsPgt
5/+ISlUicwXvBQEiiCIA110w3WNVQaRKslzm/SQhszU8kG25drhJMaJ9EgaZP419Uf6NpFIn0ils
t6fFEsWDkdOqIYJvCUiWI4ap1P0gJb7r9tbWm6wMI54hG/l1j6GieMnRj43oIL30VUwusGkJxwtq
2V1NWis1JNxN+u9bFwgA7pCxomHVxCnS/1t+XKSWY/qdbhPChtD4XmvSC9hyjeIQYnRu6ZWpIMzn
QG9uMY0OEj7kRDrkcTroZFe39M1TDIucU0oGiqc82SWMPeufQRpGOvyDk2h990CxpvZ2+KbGT4XQ
sam3VbzbO40Nx2IfAostra1SKGKgAlGdr1RmpnE12o53xx++5RLy3LJJgQKd2RbeGKgImtzp8MzV
W7y+NDgqDSPm/8ZjmHwgUJBAwDwNHsN2SOybU+0mPxRRUk/ODFMURYtHHgsFsV/YWuqsspZUQTg6
9SgLsS08C3Y4apNlwKLM19jQ7TzpVIDEHHTXSfqvVua8A0894kOUMJGGWJKbe4jxxDqUtijGmCOa
fatgEREKliP2UM9ejLPbLbL9/2aqhiwycCP9AVEoP2tfnD/C15GGRVF9sc6NqUsAGj3Cizsih7RI
R8siWHwXNWJYp1TZhFLjhuqYVTH0QdrdFEgyv0/O4YwJUSjsUJapXB/pUNpU+RIU7qR+ThUJ4yu8
aNwyE8LiFlFPIMMPuGv+xrpHAHolI2NNZ9oDFG8DOnvRWLKR3LKGGEs/wIkHpS+UE/0CzNJX9Ve2
P8okiNhfC3v9z85yGpDUNG5w1uYePEISItYe6uw7oZX3HX0eBd5JYEJLFcCpo0P78UiWKnAJLhuM
8eJ8U+WpSGOaIkOjHG8CeyCisCEdTyy1xA7+qTdaGa+Li+i6tYfNHYR/tKmjHGVIhIoqnquKF9/k
t0cvJ/ohwdRcTxnci/Xa6aSwjPw5GuronVQhbj9AsxmsLkj0jTcm/hPKCSMnzVBlhZyxIyFtSDyf
cDG8DR+UvIMz3ED6AfW0s/atmAmRN6eEqVXr0ZcdfsZWqEwC92e1wUpkWQxeP/dR7PwOfP0I3ygv
0kiJw2ugDFqCk3aX3u+p6wXaB1g23e4qhoUMqXh1WvS7LdB3bbq5xzhiuTwPBMSNMEVFhqOkW7el
pXyzhZhVbHnP20NO2ZvWDHLxxBG9lT2fn12yvfTWmSW2N1tEqHQkE3fAuj+VCIvMgwz0LaXkvCr7
W5/i8BkaLD/K1SnEBPdW9NmX5oeHcIGggdwYJG+2mHb/reKw8xPAxZD8FkEVpw8P/ceQkfiovDwC
lt4BT37gengRrsE44NyULjWRBs5DdKAdOTA7mm2WNrJjXgFO4cs6JT6RoWNNvM3jUditkMIYWpOT
A38IhWj1voBqCXJFsuteZrTJsSRmW7qE4p1XYKzHgr2gcaeE2ZtTRpwMMPqwgiwYj/YlpPaPgGcH
v8puLvan5slnKg7MYHsxXoprlv2g0Kqtq+EjXASMDav3sqOrUhOm07FK2FTmFC5BOVwHlHCGQOvO
a2gdaeS+PShPoW5YNw8A4eNdwliz8YNzS/Xkoly2j5bEQ2rbOz702qgs1r1kRgxy9KpmtUB1rouB
qu+V9/sHNEYnJDmZZNZpS4LqwuUOtLoAgnm8SbeQ2avnbCr2w5ZBaW4TBn5yOs3AgM3sWMKbGobQ
hMO0f9Bp3PvpPBVj4kb8TlzNth87w80foI2C6dG08hdQ/YxBhsOC+2clxVJLTEGHkh84DrpSI0VB
6xy3SFYoFWi+i3kZ1nWoHpBsrLV4Hwt4SFeih+s0KhW5qq//uyvnWxp/drGaC4WqyPkPNL2VR/eQ
o+SGmPa6JIDw3a8RXEZ2xIVc2UqMozp5rrfhRISARr054gfn7Rd61l+4xR+F8weXhoshaY0vq/X7
mLRdwx0f5p4fgk2ML1MlLlY0MKkv0sE72bIJAw4BdDsMp3LW8qTx3X1M6u/StnEZJjIfOy6VDA0Q
7FIy3S7H9leJrsPd3CoqHS84D3EtKo0vYWnO0YecuE1di0mA0fC4iZ1woiZs8lEXPQ7vyaswQBCg
tcOJHbr266XEAFa8q2wm26vLBwzHzZQnOZB6LQdrSgSsC6XEbS2T54c+5946B2ha2JqqloaFftvv
mDMAuJr6nc0QKeazrYfzzSU8+eFhMHSsnq3KKX8OkPUv2TFE79RVVmlCt9FQp3pOk9Z9DgWcPp30
FgMoPfrtsWmjP/JPSCK95QO8t5JbfhFWE6z0XKOLzpkBv1jR6n8ZiZfFAkhZTQuhWYLWLlW0AY1K
a/NQ2TS3t43yvQ5pwFe9DWqJU3f8Wsjd9cWHzf8euwV+ZCoenkUe1VuAPOQBsXe43KDFyL6HSE0l
fP4LCCEX8+xXoVFFaAhRcG6eMDqR4krOu7pXkGHzpLq3KNqFLwAxAMqPm8EpWw2Hr55ZzQnmijoO
dDEb7DAtIdLKt+fmTIb+1+nqsyAYpbpSqcaDPs+zPIQMaLyyIMGbPMK867NqvOc3Y3+KUibUJqbZ
NUZgj/0/wsGpIdY5dOenDsEXrR7kbbtwOR99CozerG5RwsLU/oyEMcTqwKu/6URZE0ai1xol22Bt
l/1aHCddiKG5QzqwDx/EybNKjCRZaqJoOVmiY389sC1CYc5RIUqOhPDF7b2pTCFERQZwRXlzdnfo
wabvIerN/hyfBJg7fewhqqx9eo9LDGhIDohxFNW3WB/RrX1s3IF7ThLrfiQyNEUq4Ejw7WyEwwsj
iv716+EZIt6eVdpoKtaGVog/vmFaMzH4RmES4xklwEwKZZzuyn8vEtmoeob/+ZorRKhM/GWkRHir
7ysnPRiQ4hhnANIZq/M83teAEpdN0s3azNPdAbZ605mb1AmyoaXYOHKlbXLgw752i/e+9Zy9SVY8
FbbshEXYyEXL0AeNhx/0aKjQkAUM4c6cf/AVColurChxhWvrttc6Huo51rpsvr1IAxHC9+AN6ry0
Yt/nwXbDJeyMpqmLGPtKBCxH/0W98rC/F9DlrpyjYlXyJ/YGup1imwPuUBZwUIg9+hYFhTHmI2OY
0wrEpZEiMq+QKiUp5oqnPQslmkZg1cNHTYWzdzjK5QBXZqQD3mqXMHXLDYRowRokORFoVCv7JT5a
GPOAAJZO/5Bij+HMy3aUFy1WAtZnIB8RDHn92UoW1Nc5llhabQBEqkvVL9s4FzEihuvx/VQ0pQPC
7ZU6dl6QmCApXBH9rRIbtkI5y7JCNdVmXwi4csji8qS2INCGKwgEd5XgaLPyWtoYjDSthTv350WG
dlAqpX1ZyMmhhSXQPUpcFu4CxprSva1gFLQN03NsIWCsJVCJrqVHSCp4bfVpkBSSfogzmX6anjBi
ZNJXBOxzYn2+QrCIRlzMeBMSOB7wobXkcOcevhCAloHBPPNcnYR68ORuG5zv+hfnhBiWW0F5LVzR
c8quXTSvif6Hv27LmhrWz8dBXbr7wodFypVTwMLg67A2K90GvnyJHjyRFix9aSQwrg1aXjospEjl
tONOQQdfIBsmLZ0gnRez4gXPdosF5DgOEQzJ4/3KbK5kaAu1YTtYO6NvB/EPuzqc6r7JdCQDc4sP
JkASvPH//UODI8UVEs9d2KUM/xmwZlLspxLzf6kvEz4bV2KSHcB0HiRrxVR9FqtBoz2Fs+WgZ/3B
H6+QIIgiakJ93z+IFPdtIlKpyvKays0UBDpSaBtqU/WFZ/IjZMUD4mxpEzPoCgwb9tcZBbEP4qDr
hFtz2MOL7qK637oLckBDLLdIvB22mMFYMhlixKPoktQyON4ETtZEEUQduX6tyqg3HA3YLu/nzGuw
lWwGKd/iu3M3L0b/OjFeAfeFFnYh0VIu3dHRjV6NYN25LCa5WS4A6iairswcejY5l/ENcJgmHrHj
KM6UboZRI6VMCmSW11vYXqEfQpz4jH+zpWZVmPtNQ4VpDopIm5r4UksX1/WIOOn+/Ovbol05f1nk
deF/4ppxrGONVGTkGhyoHT4qBZ5cry+nKUnYtJ25jfpHIm3gNyKcsj8tl+vS+AH6ADjMaYutVhJu
mR8ghqOI408Ux+kS8o060K8OLt8b14PBXJusEW/ReS5aJ+0nhHNLvqHtsnMGsVqNdAM0gw/zw61v
zVp3166qEUbHp/Q4Gn/VKgjCxXXrDhg07WqPIw+hjGcDyk/4xlYkuGhJd96LBBmLWhl2h4A3cj0H
g+7ulS0bN7QVViK4QQgPc9PBPLfeCtdU6sSZcqMgu8o/6VzWBzAtG1Zz/afSwKrb56AormlXMB37
rBaUgsq/GnYXGb5FOJ1nNkn4af698mHp7JWmQa+raAR5IrKPvEfzhTf6P3v9DWw9xsTdXhePTvp2
jyTZB9PBa4fHe+tDIRDIkzaU7ho7HrykaDmJVQuRxyx2H5MXM6TwoUKfXmKVcACY75wFpturTq45
zgfnu2k3YxCm4+iNluRtEDcUo7Bvjlq6Xz/Nsu0PTnGkYFZn16/Fns7mGtxY8oq0ndU7/SBlVDJC
3GJad91hTBbzxE5kW5gR2kI2oZNlNrEBveHEeckxjltC2NtyfOIJeURUhBbj9leSnXNqC87B/07v
7dsgX/5+GravhfpDjZ51tVaXjcaGR5bcchJXni5fyk2pssPs6GVuJl0VYTFOoXJ3Yc/9bG4bLgtO
um9R+6C60Fk87L5hC0W+7iwy8F+sPEp6thEZACjGo3rBugEaegrKtT1JjY1ySAnHvb4AVccTYdAV
NzNX/NoA+1rCWSWl08+hVDmOP6Qkd0fxKeSD9Dob19oHQTWBs56v2iY8E2pV/cJ966CCDLqUxJHu
HY/iXdbJawPZtI4yOk2tmMjGglCLiPbcH30ugqkmnX6EXGqGg9/IcXhJyjamaJEcXh2guI0akNgC
zKq1GyQUqzK/4jWkiVtlmUFOqhqzb2cmjwQdTpDv2AjBWhyVZ8FBIyoacxb4ON2iqvAVTI3dTk5q
RCBLTJQH9ComeRBodo6BzUPpw/HQ+Cz/4UP5bMQo2vb9PjDabntyQgLkNk8WGa8/mWjbZt6f9H+o
6Tko4ygb+hNyTUO6Tf139ztjON3vRw86iK/SUj1i7b+sRfRIf7JGB//XF427ti/vhwWEtozwQ401
SBbZiUEQbHq6y9L+x9Qa/aSZVlG6NowwnGosF3agWsGIv4WlOepMKZ1zJpSjIahgNyOrtzh/qmvU
azvwGorYm6t1V8YjRyfuXk3Eg6Og5poHVLAcH2aij030GDH/I9JWmRG4ZLYK2IPcshtXljqNrPTm
vBfc2x6jKByI5C+JNQYKFQZ6aRwYVlnNvko4VABGfLF7ZDueddNVZmwXDWP1VnD+o0UFR+q/BAjz
HKcGasbawZodkblirbei2XS0z2EpHOdI2xzwHYMU9KCsNI/MwZqNqxWHYX+TaPy+wVgDp5Y6J/Jy
bD5uAOMk+FZkg4pRiEG4IOjOZIh7EzezxZkpcRP1mEi8CLe/KN3TiWXUXuOM8ynjvFnxhDz41sff
fdXJ0QJ2XgOuz8jw8tu32b5/4eskjor+BaczWbT13qWgclpImCwYNlZEa7UFJUMLPQfGcvCmRrRg
TBbj0MZnfK5+d2v8djEwsPoSIvpbvRqTldMOihv+xjMKRKHWuZ+A/Ck8rq05B9zh5yGB9Kj/7E3S
6mexpttzhO+QZYBT2jDtPje2R/w2HwxDNwVJQaReIeeAIvJiTgetjdkmneBD+fLL9Rbtzijz8zh4
q2sAlwWqTfLqJZ/pHbJRYSQWxznx7vDuouNsgVPjBKzTdquKNuIfu7m8bSzQ9CuHP83tkatPsxti
4h7qllPWoHeJ6epeCdpUNzbrob7u5UwA9RCE21g2LgFuG/ma6B1ZMZPMFVk154BpP95mQFG4Jdf6
QdPWDVU4jCJFPB/CJYqjwdfqOEZDdZLSAWrDDR9JDYy1gc6aNIlJuwnfsYv5ZpkUI0Ubdv1MQKiR
IumvBcViRK0lqZBfN7JDaTgQ1GNDO7mU0HB+FaTXk8WVXtIm+aeZBFD2pQkq8n+a9yDzbhqvCwU+
nAt18xMINXc/2lsmjHuxVBwsfZ0ALE2q2CoC+Dz8o1by06ADbAazYMTM4/weojxpSNMjL6C2X1N1
l74kLiyiRfZnYezvdc7MDw+tbaBZEOD6AzvAHsGtY97XS/KYkUL9vsS9Wfz2uqgQvcgO9HGY8dN2
zzjF8//NcNOZ7cBFPk4f7Ig+6W7j7S51uQi3AYnpOMVOX1LiMocN808k1niLlYcYakGIbNlo4hha
SbErK3gdlwxX4JLcP9BU7FnL9mKvZYbxodEr+jMzCm3mU494UwiIOzUWCGRhk1UPNugET16WxAB7
qaAskj6lcdehQL0434w0mIaH6R5UyRRPyKdPJohvWNMEHUQ4/YSiCDS2hxTQeRxatzkPTiLOYRrc
il0wWWSiFeg2bqRQKCPrTDm3apRi3y0WYLOgbRhasGiHpEcT71yD60Ul7n10IHO59ARftgKYcWzU
lEN5kRRaHA8PvAHRC9ooqb9TeWSpyeBMPzjp6Mb0TNTcc7ez6HU0aerIGwrd0SfkHh70iP2QZpN9
F3CwrUqVqp6u+50fwuU0sKthg3+NHPEFv38vrbs6mZTHiSgmWFZ7QNCI+oBqhlOsc68Ska4W/wB/
2ijNu2N0jQ1bPaX7BQqZ0Fl1ddx6UjNdIIM3wO+XqRZ7VrSJG6hMw1PklBXJqqmymikiVE7W+gE8
FfD9NVjqXmF09BUFob3e4E+WkIAWnse1io8ojYGECa4OYFkdZxs1UjROiCzhx/64pUhnZtXtJCh+
Cj8w8JTVex93+qqyfyLlLdgr7KWVQwa9S2IXFyCzVKNA3TwtqIFPxC1bKTci35kLNBJXqNOETG3C
MVeQtNU6+Fps1kQuUR18cExA0HMLNEJ4zVZ8pI/MgsNAX6lciZJAHIe/mM3HW3uUKMI5dF6k5Ayh
vaviBcIG7vg3CP96FZ/LPbzQ8+lweb/xdEQXfEqQ3aw+GOuG1E8oV+OVGGYSiNM5xyt2SiQuiznv
bzyhLnzvvKvIqmHNAYdktK2u49bz3ao5bp9B56fl5Uv4iLaWh5NkkBCF0sbgowaxIsfxW+hvwMoA
tN4fXGlujVAV64tKXl0JBQdcvVjX1NPv2HDnKAca7OqHG0bFxOWIDo1EnU9FiyJmsr3uitULzn5E
rhCZbf5Iq3Aa1oyDYkfGwfBVCOQAt7ezWogG4Km/w+mM74GAR3zbNXkHrxU9nD2pnLxdzcSFmD3h
Hf8/lSWtKsMmOLegW+ObSsiGsSbqyAWiiCTbT2ro75lTe85XyUiUGZ1Ex02vl9HHiqGELBrE5Wdr
LzqolG9Hb+yFebqAnLFY1BMy9KI/pafufh8T2kjo2PEmElUtS7npGKDc/0Nv0ZBBZy7BDimkJ6Ju
Pm5dzPZbUI+BK3seZN0umoEULtHQX0V/iKxCZ0G+mc0LAScVcOWDRCZUsr/Bc0IeAFarqF+57VhA
ao1ypcC5YA4zUGaaY7f2kWkXLFVaplCjzvTJUuTWoiJ7mcIS4709BKmsfxhn1tTUzUxSfGyCzXYf
/R8RFztCEEaGiRh8OyuxMdYxBPD9HjqhLMk+DUK9D4NvkRtvOUXd2wZa5qRkT0EaddIITsSWL9TX
rFQNaFQb43259DOT8rCi6TcNYJdZPrZqDIZ9FNHGwmrKF3ndPCU/z4eZhR4PGTSX4LNMJopyA6hZ
lTYc2Pk2uVyiU8jPBYsDxEyA8oPr/GAONRiWSvUjjLMGdSaCofrUX4jqRCrg423K7Tzg4C8eoyH1
fs64asuODHSrSO+v+O7tEhy4Yk+kFbu1yygMwa/FtxH21MX4T0VojjF7XnUAqzlgqCe77+HEz2uI
F3U9d96EpBFr0xWhu6I8ClgsUZcPvMfIDzZ2gbKW25KNHIs14W+QTZuc5fWrcUcHtF6quKPo45oM
3uWby34PepEGVWONP9+bqpVjTwTwzMTLmdd70N6nqWwN1WZwUit3nCFqWTdURu9dzmF18Reou6nN
ljFIByAYoNiKfJrObEx5Kj0SQLnmjBpP9pQ1wf5k4Z1t62RUE89LMeEnHC31G5lbGSCDd0xXweNW
V9DjDFOHTRpnKcp5Ve+Mb2B64kvDX523NVNoONzh9GOQUbhTYHjieVSTpoxQAfxM2fj3Dk8pxX00
MyhypNHFvG9K6aEUfL2M2qUjAjMTJdewEyb5J3z+w51ZYHP+tfn7TjlRkcuJmz453kmniENf1j4a
5FO/p6aezDN1m/9rHuqUn/GnZUf2TEmg6VWCPVRufvbb/Uh1T3FMKG2qwotb8U9nPZO29zOymkfH
SNh8EjiiE9TsRtHvt8Q0YlHSjnx42x+qD/qHE7T037WFpjkaT5/eqScVEnmRBsQKAl+LLFJ5onrG
0cP9Gxq3QWnwxb7OO5c2lgzqZ1XrnCe89lqfHMNPusvrSM1qzjw04Sqir1ZPGES4L1EWII7q0vz1
XmiVeY3ZAuegYC+AYpMxotxu+dOBs3E97D2s7mbnzvJ7vQhBCV3xKDNSz9siwJKIZTMndfQNGwoe
7yzqLOlcSGkXAL+2Mf4KL2L9+7g7JFdjrCVqBdRMOiHxd9PejGQRZu4YeVOR8jdfgfuX2KIY01/i
9ve1y4eA6S79Y3udH+MARmg+zBLScaJLvQCV3h2qcgGOQuJgzo1gnUrFmjZ+H8LlXrMour9WOOkg
QBgWu9y6BjWS8T5ECv9IMh17NKPkRWl/P3sdh1/JWIP3uiQrOP5PpoVpIF162aAj8dzI/B8Vux3W
oc0bljRVeZZPF6YwMkGvgEVHip1RF5qTQ02daT5KLTOe7TlAk9pyRiO2Ky9LMeF//M2Qd6eQYsrt
PQr83iiIGr42hoHMXlbynjbO413605rMA+d48MvpxHB47jBKUIfCELhwSIDZc912KbultgpXa24B
tS42/mliekFBKMUyhlIJl0TD09MkKTVBNOjJp0q5URUqk4S0wwk/KflmsS+LIoKDEb+Q1WDWHCwM
MQChAvRpvGNotlsm67a0UjOqZl1phwEqsVWLbs05+pqIqQbdRi8EvDDLZYOSqJdPGJa3WIOGtT97
zx7sFhPhV/hYQWD1tc2Ru121DV6Ma53E5MunXSqZ2jKAMRIUMnDWbHQ8DSOfJj1XWXydh7ZX8GT0
aUkrR9vazkwck5b25HK7GKiuJQR1lffmIs1MymAuaP2dFuqPVtV5q/Tzr9ycLYtTQKQO+nzn7IGn
9VuTjFWZqIbCDgKF+08LkQOEB3HEH2xbG+C4HzsETJOs6HWga86WmMdoe14i7/XF4BqdesNUgmbx
h1JObm24rNnOt6pbkOSaMYNN6cca9+RMtG/oC2/MNlHJnAmNqVITdMdlqV8T5ERN9N/mEhkLR7GB
8qfDZ5yB6pwFbUyDip3pQwde/CUqM5Q2TnN2sMdGNT7CnlJoNOQbru+EPfC8S58AcNB0AzngUq77
OPKNorFFtPcR9NBZQRZ6uAd94IEpjrz6BcNOeOBbwVXBO3ca5I9o8QWN4gDnddYwbXORX8fxdbMk
T/PYaEbLGM91j5XQ8MNnOvYf1w7KFHUnv+3GZ/x2JLudBzgY83jbzxZEHvh076Ck2EfvUVFNe2UN
UPP8qkPmAxUrd+Vl5pX5q1BPdwFgcFURZch6Gj980bZ0HIjqKvuwZ+851AAUoN4xTQfkDTKfOTKV
GJHBLbwDaFDynduRQavbEv9bazcww2lSVe6wnbe8G6pYS1q6LoMHElw1pP/SABwk0bCA+kPzJ4/t
5v4Rh5GB99axAC7fXdLg6/OpFrNG5AvKd6DQN5ahcc6Z9TR3NudpoWVAnyWhY8/rdnYx+8+UE/AV
lIHUekhboXXTM15Jer3AcxrlAAlIPYkpcR7mtDppqNDdVPiLpkThtXcbjwf/HaMivQv/aDtRxk0o
f/aIANuqbL7vaulGB85QQt5pODNiXP20iw9nLM0F/kDe7ybMdE9gxj3jnDQl6qS6d/mP1SUzZqem
WCrwJg+6MtgBDf+cJ6T/Q0hkl0KpA7VXq8nyj55boQGQ7gz4SZYACqDHQz5xc1+N6UUNc98/sEr1
lWnqDhLU5aDZ3AtmEP+tZun8AJsJVCzFomv0UChPpu8sJbT5CqskJj+kywM96UOgozP6qED7ddsB
71S23p+QZwmxgIQk6/Ab58I28OjGwDDtAHUS3F+ZfSuqeYX+dM1cy2S5BGawpEjcQquXWk1RtlT+
HjGq1Rf8kWxoVVBvWInrYaNBKMajchkvzCJeNL7+huB+PMI9NNMMjeEmv9F4wvVJYraJoTS9vSnA
IoTPQ7bY6JQ+QMeaN01CSRuT0/rBAd9SQZqtcv/f60M4QstJBEKuIcVNO5qSWM/3WSMwxYd8+P0n
2c0XnheoRdTcn+qYqjEWY81u9JRJGqnUjglFKJBzRdzskALtskmyjdT8OR4WRFbtS05cd3Ky4eZe
G5crcWpFQ538z1C7bFlePv99753EpYF15hbFktcQ9ArSB1Zvq7bjp3tmmZxgRYMNsDLAOl1Uf0RM
kLR26y3Z3G0AwKL+yLrYXHCBAtwCKAmAnszZRG6Z3VxhGICW33AY5rQAlgIgfjjb2AGo7jKGOzIy
2x7irHZ44geBM01/YsRjgiZJgLDHp43Pmpbd4KsCkCE2ankEY44HfSt18BBLxO/Hdm1OEYGZQ5AN
xxdkEeUPGk4hGTl6gSXMChWOPl5rya0E1UJV7F0ziWe3t3Oq7A38l1ZaSeq71iZZ1YkiCSpFOX18
/Eojp0TIPEvio9wiVvg9aqPw3rQrFCI24ovlVXFA3YAfUkbw2E/XE3mTnRpx+1SDrzNtdAH8OQ68
t86t5Ov3W83NOpxjAihPCbVc9Le6/TqtNmDAMPU/u5fu2GuyKwbPdkS3two8nJy0Y3xGpxKDPfi/
4CdeKZBBCw3h0gyGtVhv+gD/tcRynjKw7ZBXD72A0EeosGxcB0pA4d50wZY8JaNryfXXPlWECl6H
DBofHI6hnCnNGA4kJ/sytXw8E0pqlkIfLHaPgzXBNtsw5YYj7KF0NW5m7uHon6NCAOEIn2tAWYrV
C2HwfCthFUdqGKED61SvVhS7WtSr17sA9FndxhFnwYbAV5dw1q45Ssaz8MfY4a++YY8v3wLXJ7B4
hph/T83WnHCZ17cy63FLD13EbrBF0/JDgMAmpJelst8CJF48llfjd2Yx4OjvDvB7tp00vSARWuNS
tSuShELn1UlgayELEv/CWa6HqYACj/WmnKSHgiXC045xMdeV8pfj08oha7UyjF7y/aIQFUEnZzxK
WVf9pcDG7nEfZuFdQm/h053ReaJJztkLUpVS/C4BpSktWd64C5RxY/VKmKq4l6hgKpWOGMR9snU4
u8333GgmM090wos8uAX4m9436LNoeTaFOcWupgxJc/wArA8bqGsVYy1R6YfKgcC2pFLGjreYWDea
UlNHWRlucq0Ym1m1ToQwrC1YANc6FiQroJg470yUZIBJ0pwtUPSHnGFhuGt+fdc5K0pf+jLkflZX
7PXOJAkls/XxqlStUqFiOswVj7YXjsm1qy/evThNeSsyF/elOW7STGQ3f5XMXdzXFV9gSkq9LkRz
hmJkr4DzIGNg/b+WMdv4WnTpv60MsSqx/N4MSHV4jzEwYUyrWCl9hrLVA9kzHeUOxRl+c6tGBweO
HC+P/0jf8lEVJpTEm6IDcBvXueVas4vDedy7vWKz+UjfUq7TUPln+QA2fSCI+cBP5CUfgosFPqr0
oVY1MtoAX/g1vXSBcItf5fUHJW0sbkHw0ovqqd31chAWcZoj9qLC5GqGY2edupcHPhQpZSBzzdf8
+rwMtXuRoQjoQqUDUAPp0KpFA1LdMKw66QmBGdyGJ+doCf9FjbLysNMK6DINVTLfJCA1lAjsOENn
SQOFBFtPJh8gkQpVERY/GdM1T1g3QsmGEzOH4RrZ3r/bgZNBFVa3Caiq4gj/RnQs+dI/kemGPWeo
dlLj5djfkTLOJ+HnQN4llq/nmWp2s9KqtRJvthGYWgKX2at/09aNXbgDMk9V8QUOqOtxWmLPF0pN
TUh6uFhAcRjHH/Z2oBrduzTbcJb9J1cDrmzciFRTxF/zDtojwcDTSeE5RDjE1UqZKSTb8G/a+su8
FNxAPYw6dQfBSHnD0Ogd8rK6DvWP9jVoVK2tujWMxrAnoo/4HjpgFl9W87GmQnJnxDnjkEsyKc5Q
LOyaiEPb5M1aCsXXVcBTMy+xYaTyitamLtZ1t0WwHC7e/gPxKXltlBA3AT8t/NH5PUaTuHhcov7R
CMYzlsLHT1MYPb6Dy7xl9AfdlIfWhOI5GaBzG+dC5ha73dXgLxCBrKjYacHEDEwdMHzoQ5+twdFI
/rNM3McrnqaWkhBul6SwF3qKIgsXnz40XqzTl5IV7OK1pifVOakIfI1nswkdZTyYXenExfRLzYOO
3Wp/ghQq28tw9Iw2BI6fdtxMmQwkQteew6jqgFT6dnelSa4rb1csHFU1cHf0DpHV9nbbjpBSnah6
KSvTdnj+5Lel/ofM6b+jd4Z3wgL/8uYnlsEOkEu8tvcmlAQXqpX3IvdQD3mPNXnZTVtTlPe3ylOf
g5z3fwXsmOO/7OYJZZnuJdhJ1Rg2f9YXxTECFTbhFV3WUzQcA8yf7lpnbrD9E2nBp373NYkuRqvH
Fi3LPFtJ5eMad1O/zCpm2plAwyXRNHofD5CyJQOuUTvgtKxn6CdYoONiL5LGiTSqu1jlluAPUNk9
8Gxai4tGHhdsWKNh1qk4kCHcoAxv+LAza91KaPKIRQbW9v/W9K4QF+unsFbp7gT84NFT8soH8Od9
N3dDPkp+zl5Bi4u+mLDZRaKAO8CcEtKul/z3wCKaXmza7CFfGtK0mnjKV8TQP8RlqXb0MKxIOXZ5
c+1lvkJ065vsBoXYYazHdBJR+z6ZvIITBzwf/wC5MRymk99mG8rx+RazjutndFs0Az1GH6hmyAL6
Zaqj6igwnJhibTFojyF6SdXsOc8REUnjrd6j3TB3MrSRBdr78ev+VWcVUs5mgXaUAfLWGHuNGoZs
OriUgarkqbm3hJVfL0Oho9IyEgmpZsuztYEHX7hgwk4SqKTZgrffMbJIoYL7KHLTHjmTZI4YmBeI
VgcA1orKZlrUCyqq95H7y2NNMrkFrerVpOt5LFluPB6C/oIzlU40wL6GXTiVACG6tkeTJPeZ/QIM
jaxEC+1AdRJey9y5RrJYeoNHXV8uVS9ojMxIr99ye1rXdsQUEljK/T1ptZ2mUcS+XXmN3pnHC2a3
zc5gr7EoEjC3bWxAuX9f5RErHfFPr6hGOmg53B+zoHL6+vXlH0W/+vriw14T0ZUQq2uPIZZXzF37
e8U0dENSSu/YvQlhwAlIofZLK1bSSVFL1JlQYf9x5Qtn40NZyf1SqNF9uHKpBaG2FfMquXnGVfJN
2ZFEk8G9Fy6P8DC7YQzSBnzF8SxX5fceF9aVPUyXTfmf95fYfRwEBTqFOSJBMGoEWA+0u5mwmbCv
BQNovDFvrOF4oqBIDax1Hf8es5+T/W6bnULrkmiXnm8Na9q+pkw5S3RArzyKMwxpuuAYkCspg2kC
ON6d3nkKZOnPqJ9o417w5vty9e+MsKE2UWAHr9ZVre+bgJVpYuPgYLG3NkzxJwbq9eU2ezQOzCaY
vc/IxBANj2WHPTLWinjkgi94ag4EFYb4d9/hFgHTO7LqIgp6U+2XFgjSJLCJ9dyThTi6Y1HhzW2U
bp0UuqJZRx4eMIE6yBIqrTDqX1XI3ZUPtnEFa3TSxn8UJEjosM4SAthVEDVOC7niONzookn07BfT
nyRTPe7+oIyqcYEiEHgGNKm/f/xLl07ydFktDOiiN+aexSf3U2mXa2q36TOFdWzZlKRLlSjrI77v
At4jhH3EF8Fxk/0nCWVfq6rAIMKweEmY3+Lwq1LnuzNMeyCPAiQv2TYloE4zjliSFtUIhZtOe9Ch
vv1qPedlbrg81NHtXar3vG1S5JwdpPcDoMztY6Nzxd1/P/CfhiYtjBnChy4TPQoGEHBvZmZdtFCi
fGltePeBJruFM3N6cS9exI4FX8Yh27I6ZHWOZqFf0Iu/NdvGStGcRHHa+5bn0ebHPUwjvgdtdCwj
ExRN/v5HGWUVd2LuJrVW9hRIzwTEaLFNrbqwYmqdbjrhhX1UoJw9KgV704F3g+1n2SZXqFmj6NMm
ZKoY8evIEmj0PcGlXQbJ5651VgRpb29EazqaAzDj70uu3pSijj+m9OntSh724fTkA9j+Dl/II6xy
JcmERjTkVowkzD1cDb4FW57+gyln8h+k4aOEFSDbgxfMiYdMCE8UN2PsX0Yj14bVJfK/Fgu1IvOw
H0lquH0UEqU+pf4gPGG8Q4E1U1n3oF8UDg0CxFxUTKJeDV954O1WD8tsMwBqykeucV+dtqjgsEgK
FZ4tYPXnG5dnXqWudIG5yxTbOCI0f+EdLl08OIdaViJapJ2bJ7swtKZ+EkIOALhhOIKC4OhsqDQ9
bE2I2wqvbDuuKIG+ZTHgQNYWT0JjFaxspxJe4e4MxIr/ZBVez8hPjkWMJ3KY+SXe/URpMkU/jK6F
8PvxZdWDXUHzangJqP+X/Mwt7Muzjbh31hZyzHr1cH1otvd8G3XI26LiyIJOjAH9p755YFOls97z
ZPiAg8tWtk0ih+N1jmE0KGZXdB2LkZp4ijLHkkfzr2RHy2iRrfTBoNJW8upCw2KPy8tEbbO57RpO
Z1WaSTZplaFpTvCHmC0v//QWLMuyXjVLjJsdofB790Qi5RzyHNQKu2840TyuVjWSW8OYZL7+gHot
ymN5XR+fLR3NWECTEE3Jn+cBVERXh36qBriJ2Vtf+MRIysxrt221Y6EgXnESlfPVzMCnuqzpSkCk
YuzvErPP7nHhj8rZCSW4tpTFhOIjQ/1zKMx39bYbb4FlZVXywnlUzqPjcwPp1YMDeMzv0cbyDeUL
QyIRO29RcR8I/yRRQipguW9/bk4i/YYyW+kriWNXWZ49dMaX4j75Ar+PmQCO+YxW33E1HEiMhnNh
/d0ac+2PoVcHbFu7vpmvquGsnWHW1lfC65ZeyP/UiMx6Riw90AENntrjXwHI2uYdvycz1FKzoCEr
mtfvfLRYMQ2eeiGNZKG4l6SyqEa9YTjy7DSngrvMF17qs19f4Dnx5Hjl2lZ94gNREpgDTEg5BU8h
YtHDt882lI+zoKSgS+LLLNodLvSTrRfp7mcd9H4qP/1Ox4x/ea3UsG8n7/iEvi2jJLY6l7V6fw6U
knQD4CRsAeCBWD/Xf7yVDg1xhXy+U5GdyOdU29TqIH9/ZOZLkRCitNlAwAeDaXTMAmd+MdsOEk92
M5DD/qp/L6epdPbCNrOlQ2frtVZRQrq03cJKOPi3RZQXe33UXPRbzNdlI1thDWmq9MA3UhOVOgMc
9U7g6tqp0PQZpWCUg0wHba5+HBP22adkSYdADjyLhbfMtBHLcXV+UY0ukucBgflCf/zD3LaPm9YD
kN0AP5+cXvzvZ62WQpY8+Seilxq/KLMDpvEChdFiUpvQ0GOWuqTsyOLevavRZQuPzleo0rXYpeWi
vlSqMM22SNtprb9zGnFoaMiDsvzHZnQMs74phIgRSG+Vpby1veo8Urb3khr6qnxP4Z1vJnLegNSs
HlnprKyMKKNs8zfL9jqRl53Z3gpCgd79fAeqz5RCXpm2qVxtlTjbU3hRM0YYUStPzMg7YfHllljz
NCm0hnbM8ee0KOqeUXzKwjgBcl+rXE5PIFJubsFpQLkbix/8pcdkb2lfdGSkq4tYHzzAPXwd2lcB
UlTYOZVfy9oXYeoytG9xUMDIfWkOMovnxMF/k/ESxB2qSsViRBw54TRw+udzLPSDx3+DSMOiO+XS
KE/HygASdMygAB4lTHhEE/7hJwboW1qfWFdMeHIfCKwuxwyPDbDNL4k9Dt/VR6fmOWrrL0AfK3ZU
9ILKhn5qFwNA5GcN2HvXcAZafa72VHu39LNaiiprXP3NA+bkDLa7atCP0YtCvQdLXEgWvVED1LEY
33+yeXjaBPNz/in3RdXK0CuUatUzBCTeTYiFBS6alCFJxTFuKO7f6sVKa394jV+y/NPqyNpAfvvZ
x6KY02A1avSa9XjpArIwORDFR00qm5s9z/JaHQmKxmqunTnErWA2xdG3s7aC/D1A1uQ1AYZYWZE/
Lr+nnTJE/S2oBHbALoHj984diN1/aH9r9kmvzm9JweruDCXsPtU5+Di1Qu+fPOPDQp39ghGS8iVX
MAH4+6JetRubBRBRYReSBSUhPLbDB3apZQU3ByVqzIV7Ztat8dPDdIAg3sTy3/js6tigM+okTtHD
tYyelMOrlvezAOXSdjiQrAI4Ib9wFDMnEEAtHdN782aODoZ4xftH7TbAcfgYGXeaawcyH/y20e/D
0jUykiEbiRVd8bqeCZRiYmtetbxXqvRbgyPt3G0a4/FGbMGLOpGkPTXsiqEUnCkfud/Z/86SSml8
pAS94iQJpxCP6Z04cCUQYACDjKi8nJDqajoGR9qK8PaO87q/Sjro3y48kkyOgEqbpCZYedwUoX1P
+xYNm45KUd95CsyOiZYRSnQWePrDHGuJVRuwSJEysKqoKFfbxBc8XysoObiZGQKlUDuAGM6kEq10
MMuOfco0zY+zO6QvUQx7FK7Yui/8JalOU/1Pg4elMipj5gpoRGmcEHWlJ1OJnYCqcnPs4o6gHF2M
JJiHKKiX/6yOLwXuK/LFzlByxK1A/Xp8Vtet8kA0hBQDixyYQFX9M1jCrOIW+D8Q/ivgcgxyDinT
05RfvKPZ3nXl2EfekHvFZ5SChpcyhd0FqQmUpmIBsUghqoinxMbwg+a2FG5dEiHGCKkyDXNEq9o7
FPekJo3OuB9ZM4f844mgZ/9V1c5h8SZjzv1peoh09Z/qfEa/t/c3RmijHRrM5SEj8oZnfVV6cTBZ
/lk25sTzbpyfGDWmVo1IDvM+NGOaRNLZcdATuItZI54ARU1JWPOlgeTSpM4Qczu2cw0W35f5laW0
UZLpdtvHuqC7k0xUrdmTKkJigGeZGuqpNgQLIGxc+ld8vlXNVIr8pHvsHNRdkIPu3IP3BSNL1/y5
g18B61tce5PBGD3lWTCdfirYAx4JSN35/FcbwvwWeCUHl8NXfrZ7q4Wuh17lffuVM3pxa1qNRvM/
TXRWNaX8B6jyG8OykcRfNfWm1YwUmnqICyuq0cZNNamxtcT1OB3QBnnS6bdMZZb69+xaTxi9waD7
MkLgA4fS7CYQjuW3Xsy2YMNmR+De0pmnqblF/IWRv1sA+s7TBVhCt7geEFSLNcbuncezUmHqT+72
UR7d3F0lIoG5Lp6UzFLy8RS/U5OtpCncRpGF/BBJITRLEBzTLsjdpnmU9qYZ9IO6ItrTMqYOLvHs
qMtn2mlfJhyXB7gHPVjxFGvYXfKvRheciCibR0pyKzIlXU8Ats6X00B/y394wO2T6H6Ca4RKvGpW
lRJxJKBEgF/zUFujGYV6Ir58sn9Yh0BbBT3FznedBpjFju+MN9E4la1tqHU/1YNvUKLhvUBRAzH/
lrdEIecc4u6T1Z/Hb8GwwvZhM4Nbm99oNbiPYcQctboYmBuN6G3MiTwSKtQpAGAPS9sifKtRWfaX
vkenKCbuUe+2gQOXQJUu56UlPTEkANlhcaFm1hYterxfdcArZ3CV3dpVQJX5xWHnr41DNtP0h0QC
cipUKQf0bWAZ3cX+86JgzdAa/kHs+wVNmRW8DuBzeOjR32leiBhgkTN5d4uAy9GN2WOxy0AXH3fr
C5ClJ3l7FaILTJrZf0vWhPt7Ny353Le1HCiNnYTCdgfTNvTPvmwA0/TewZXhjsX0EJe7C3Pmhoc2
dWq/la2eXUGB+pgh5B0AAzeYoVpCUpRiYLkyBuf6Bn5fqAXajYnArquyH1Ro1sj3Dd+oxWhkwrlf
+mdkhQrsGX/VUMguih1oXjIfj9ENhhE88otIyezkBDXB1I6btdZ+AJcQNqTNpTUg/fM/DHgKCAtj
XYJm2zDSCCPiLVCcgr3HfAHHr5CPF9JyrGmP8M9voE6FzqDpKHpdb8CoI1Vps1tb4zrKTnHmcNGk
Yn3knfzIMRMVHEWGc736TrxXxexzCnA7w0AevwIvujZnrkDh/sI6oM//kuBp39GwlS0yGlAvzJxD
cPjPS5o07LATTOUb24bVKIvjXrn4Dyakg1zyoB+oW7YiPOJSVjo9oO2+r5G6+k4L2MfkWZXvPXcN
SWehYYVPJ0UPqtqwNn0PtDqG/9wCymXIXa1me1duwQVzwayUA8kX10TAjvWo/LeYng84LpPX5r0Y
Z8Phc4Tj1Zx4WMPHY+BqVL38GQDXdFoXZJFbRkZkzE7EqWTeNPLHce5Co388YBoZ5VrB6rF+xGnQ
PKUv658zA1Jimv4kIGjm/AUd9AjCydzusUep1RT3bilUmCcLflYaHq53Dv237czl+YEXCuQ/Dk3d
RsRaG6bf++nOJwSDQIKxDyGrRrsIZyjf/yaB7qNcwtC6WaEQWC3GBdDBUWLK5G2hHKsPbt727obz
NwZK1km/umwGv/S88LJv5oLePjPn8lcw+FwwhoJkQ9V96tUUk0CtLnnDUhuh1P8ORqiz952aO8ss
2YkUupQgb9WzaNY5jckJhuIIVNqeUi1mlJqnNx+BU28uncdjvqLjNfnnu3wy85ez5IXfGpcVPwn5
Z4tjiNSZtds3UErrVwTubeo/5QCSJ/LubgdxjXThZqac25r0cpR+ZH1e4jlQJd5u6XsA/zDn2TPF
rzGGQOqEyetjE5ahdRzeBCum9WbClv4vcrABG5soAg/josjCLLW+S3p/6gHQrbsFcWPwAFjTH7Ku
2PjTg7WxKY6H/fk0xBL92RAaWBi89VIAePPfvy62eJT/K9VUijAWvGaBdeptYvv4jtICd+jE+iqQ
uwBJIkNygQcyK0l1QLjdd0XHgHzyarEe8PMye2k+SZyrVugic1OtYWtdmW73ebll9IOt7yhrsr/a
cZ5i5ozJt+lAphE48cC5L2D1x0AWXoYZqHGbigYj4zs1CK04xkDkER76lHbr3F5Jr1mIQ/EFJBuf
uZUcPVuO10CfIhBHXAZv8GwIJc2b2Dq5SOtsfRJ+KzVowQxvyIii5xy+6sLGua+zsiq67TgH5vl0
pZz2AjOOXaVfP8hVI6lyqnc7ohO3a4IzVpBu2j+OnMt5/tr2wqU5tO9LpnUZIp+urSYbPP9srB4E
ifLDHW3Rrwk0QN0z/42dydU9WjDVXHMPOqUwZEVMolNyj6CseKvmhMinNoXC40M6IRULz0ID03ob
GrSiPyskpS5lLekJD+/UdcS0HZLGOPnzA75vgKCUfVw6OfHD7wuHssMbZcuAC720UPl8MaEMKqVM
5tsU2qqLpoVYucH/H8o95f2FTFIrt9xOwUAmb6591zZLnNEcZxVKQtWJyhPJSiwQPAorBWCdD69I
6oF3c0RXsxNJYLR+2CXN9gYzx5LE4L3KSDq8EY4QS+waOlrw165i5wp78bdTezIC+EKWlUn/cxDG
gQD1ZtyivstNKAXd+TJkZx2Rgypk9MMKiJgPa6xyh+Y5acxBe1KwmpcrljrgtwB6wHw9uUa/VC9j
WMbzjdcztfX55vCUFIzunjAuKGeWXNkPxVWNzvRDVHoMYEJy+uZZdCl3FDs6jishEkQf84xjx77V
JAPprEaZvEO71cOh322+kaOdH9g57KxjqP6VR3zDFVDV8QHh3YkIz0A1SjEBw0/QdqTiVo6WJvYL
cPsBK2UOWGOVPNT3HxfHDMGdj5wYC9ZXAMR5x13NNBv3HBu3JXE3ZAG5vx7GogpHlL/+zKwS++ay
TzXpUnZXYd9x+KSgjiawWT3GC/X0aiS6kw9CkvqDXNgHj5kJOtWAmBRkYvwg9qCTD58drLutYANx
KO7DsDxxBPjhpv8MukvromR4S6672eUkXeqdnvcdWWBZs49RUW6VDzoYmrVl32n33xIwB2fkFVT8
gk6/h0MhdPpgOnmybWWTHp1yxpyaXx+DFh7uLDI7KDL+yMnwV5eLuGmEnxvaaNgWXrTwFOG1melI
mZ6At3AeNc0UpTlafeQB3Rdyiym97e2Hjsmg4t5fj9eAGk4UZ8sEKmVkJYHFNf728/ixnuAkp8gx
YLav4hjk3K50cTalL3rx1wO/0sX+QjsliiMFskt/J7q5p1eeELp0yHBDiG5qf0MyhBel6y9aeWPB
2pkeS2SdBipjU5yitNqLqycGAXDZEcy2GK1/3ggDSzR6Q6kUZDOE4vAeAwctRs2o17TgMXSKU3yv
oSiqgCKlBtADOky5OJ4F8+tXvzWuUsmBsExyl0pIxYSiXOul+X3CRLxiJo0VG8MGu5doOaopLHOM
silK4BcTvevk8FzskW/bhoKINGlMQ3wt1lnVzmnHGu80dnbJH7cSC0wLlCF/DWohF9P9RxBYSIVn
TXcnh+AtkuqcgDm22g/0MnXFVIXqydJRaTFgKdkuTfY/wXafumk8xcUDGAgcGOMQfAgAhhgtmbLQ
aT9NwhDSro4vVBK85YG+JmVjKc7nFlFF6Ma0nJWkmtHAggtFj6us/IfvTwKQPWmgKC5wiT2APZ3E
5hTEL2PTrwclRuR/QvUq/ThjxmuMVEzy3BiGGo++3TW+/VKWKqys2c344PzmdjhT+FdVtXQPP2i0
qJMDfMGCnlyfZuuujnNPXkbw2zWF3SWGU0g4aBwYlpBjO95M0cdxM2Icv8eRmJ+Kt51kJRBsAl3e
NGqQ1s67Ryu6suBgKu9zIcVY0kQcZXKwKKyeyLRvQ9KytmYcYCV46Ih8sdoFQHdJPoHwOyzsRgJe
vU053D8RJUC/zwasZ6z9Si/BjEbNDZ66iMtlNXnrdxk7YmYMRhP0r/qFNL7ccujj3mgkm4qsXlf0
ajYOV2ekleOkvVU9otcPHqFjhTZST6aUgw0/aDDOaA1UgTz2xZeIH5G3dN92IWya5jILmoM4kOOZ
rm/VWT5eayKamDHlqtQALkhG72RFREnGGE16q3onWAZXQnuHEc3OCeImnIHqvk2J4GOYZK/iw49v
D0qphL7uSvd0RNSNMsi6tWXYPZUb1s1pzSH0t7Dh5wlnYHpyLhzSuqmZEo5HHXXhpB0Cm+oqfD4f
QtFRf2rLNPQECWFB9L1ME6HPPfyiHQdIqwnm4ZqptiB2MpySkLX5ZA6NSX2gRGmRvph5tT+ejB24
B2xRjg+FmMSF5GdMhhQzdKvQlwMqLfKl/rqrJj2dYdSmTw1vj07ufW51ZZgrT1L1edQ/AXOtkA+T
IgaRYFCwLL7HwHRFMuew6U4bgxIRyT1/GSavJv6HP2kfAz0ZSqwH+0kgvCQt6NHJDwkyCYi653b2
sJYfb6hg4+u1mM2vngGDTcR5ejPFC2AtIW3KF0Rvx1xVz4lnTV7ptbz7O9RppADVzNSsx+Rnce0G
WyLwlj3t2MxaU31XXBSZ9QO1P5NfEIaXC0wwEjKbf7c5+DtnHsf+EGgrmfRZga3tHFfxYxIiSqEW
vf8k6DiLfqPDngh598FR55B2NRTT2bIgWiAROwcEc3RakewjTmRNyMxPy8VSY4Jh/Y+1qv31Iyza
2pcjIDIfrtmx0qh7slkVAJv8QlzEOBAI5WPvO3he819lrr4AwASu5Nd2SHPRfpZw7Gw1hUQqqBge
HSFnFIgBTCcLnEuxC56wfmPk5id8+rKd+0+Q5GccuYwJzqw0ASyMt+Jk7adYViiulhEhmYtQhCgn
+hWuaF5bYlVxUlFHcCOyH9lOYoyBBQsmnvPW+uZA9gTwujPDCZ12r7oH59bjbDBi+SHS9d1XFN6E
qIHpNxoCxAuC6UljnmwLuGrgQhYBJiI1k3AOxz96ybbG8sPskwyAuF/vGYKuc72MDwYfsGVqny2T
vMFONPSsImWjvSQ5eWkdpWXxmZna7oqZtPv0Lzr1FPACZ0s/VCdM1UPrhv1Wo6PAeaxx8IyuHxR5
dreGSW42fUDCBONjUJHeHlRTiJM8vTM4fCyFho3Pm0T50SadvXuiO+hgi/WvBa113MnrXQIJgRX/
1B9z8WoEIE9Dc/EROf9X0m5z1oiqeXzT8yRH+QfGouQvUZX96zxr5Xg/ZX0v0P9szAaY4eHwHxv9
pqAQFkEw7Ua055m9iBgw4rnNc/Qp2XZC6LYQvFKV69og7wwppmc3l5XE+Zkhefg3nP2G6EImZJLJ
PLp8dQVpg4MiFOhIWYp4BvGiFEcLrTzX76YFzWV+LmG60Ekc47jBs4DUyt/mN8w1nLvvsakqsAgy
UkVI2tnrn4NpLkJn/2IqTDq1wi3ZNOHxWT3FxZIy3LnyscDoL1vnyVByTGVitg99AVyfGzHqVZY8
ezj56HlMmBeOH2km3+q1ls4Tz+dJVv+MbibhjhaZx0sxsLutzuzhfxbBIYpXrZfcWpFPlTJalYfv
g0QkPY5keLGzDV94yqp44MzqpN5l/4/6IA/Mz59IEaZ4epd+E7vB6M5lJuMCaHvJ8OcuZvCcKt9+
IEMO3fX/ViBEHYCqhAxlhFslLYPs1rD8GxEOODsSM8TpR4E6Jd3z5SSOM2dz5Nf88zXApdZGWPM/
YacrSVmHoN5mE7ezp4Tpw5MetesrH7kOjROT7bSpUABKc/A/tbLT8l/T534WMMu7r2GvPTs52Veo
kIe1c+bOmBxIzWUZypFKAV1AKiyMK1wwBGYeXVExv3TuLJd+/fhPIhGghRe/NDkaBF0aFaGa4SR+
HVbdahCMmpLo5Cxu1T3+otxsfbOTMgQMWYvErs1FnxN7eAxm8KLszCbMEKG+rMp9gnsI44gRg5YR
eWL/e3YRSzjAufKRzu3SM/pssFJ9MtqPxeqV9CyAQSiNZr6XX6nxx8hzgHbeZQuGsB31yYBLG6yc
jYxeXhvkIzmeFwAuGK7UmbHVWdbz60R+B6bh6Ym2IGI7+nJ+npr9LsG7lDojrFIO1u76tx70d2tI
VO1zRP/tu1MoQV9Mc4Td9jFCVhklVByqWki4FxdwTGV7P/OVIraqLmYaoaXgDKxdk7N3es+jN7T5
Pq7tMRnFPIA8Hz3eon7MJlA8omp8TaXPrO/Czu2bDKNEjlhVf1rlgZ0epd+sfvRntw2l0L+jeY/q
x1+r3rzkxQY7eH/7NXwvwCP+GutbohAEy+skD+7NB62c5+1xQxmqavtGK/xfr3WSDHDQzZRQ/3EK
ehySC1726MUIG9NBe9RCG0E3s/a4tzDCGhPiuOxU4dXmVb67ESEq4/T4m0w4eF7oI0L2WSk7b5xr
OBvMouDhEQbk5rLsXyfTg7fHPpp5Q0Yyoj9YhZw5OVDPuzRjjykM94mE7cOjLes+Qss02aUb0lt0
q5xOV0MBPPNWz91XZllZb+eEg8AcjPvmBHwLGvsuTDmaFpEVJ9RIgJFvFxSHryHyRTYV7fB9Pd17
NEkvsP43Vx3c6+645CPxusZC8lozmwrQmm9kgu1JDa3A1iriEoiDYYcwb0dhUcvNYQMWIr7Ofsv1
/nRhlqR6OK/QXGpf5VfFO3OLMoUWMiod2DGdr8helfBy3mCXbLUKR631HeinwT51g5s1gNpcTdfE
SQ3v5aSYhIiG7048t7oCJOjrwhVQPVmBTtZEAg9alBT0P3zg0p7IFtIEn+pzLxeA6ItQ3tqvj2zL
DYcCtU7HWbrnSiyjg4fx193bIiZigivprKwPVtNqMRlGOMiF61QdKGxnLrOhooRa2v0C4wm/JrvD
tya7wFfLhi7+TcGaUtqpZDEhMzm4oumn4HSYI1bzve7DkOGGc54zk/VgQ20rkAjAngg0rMhAC+9l
3EYpY4ApMqNdXdQawjAJGQhvvPon35c38aa6Zd2BpNa6DrJIihoB8YHqIm5E96ofkAVStEh8PxtC
b/47KgeCyUDN2IEfrbaGliMfxUGLnGkruiWR8yqtKnXEtnv0Gte24mL1KcdjVLAtqqcqA+zSmz2a
9yauDoZqbSASAD/Gg4+urXSAjC2MC7txMMBS5Rb5yBf614e/MCFORvfb9wbj7/A4O2vARa/Q3Nwf
fZIPZApN6gemMaV1lJiQAwSUieaLdsbjCaEGuWeZlNB0hL6hQ4TxmrtHdAR1iEdILy+4A8gtYBSP
Hxrd/HceHQLzbgcDWHVATSIulDWn9xA74i2rBl4P6WUmpsF0yZJLxX4ArAmuJ+FD6PpXEo/eidnL
PMb1FZql52JYXsKySvC7rFHtN3JICa5irK2NowX3+Q07U6ExoJPXuJvvEc8DOORN//4zwaYP5Gsr
GvHP3H2rXNVfAXhLMTou5G5gNFyJdlXNGwaZ97FVmIw4mgJUuGAq04Rp1GSoqQD7NXYbtcuEMYkN
4bTZdiWIr/tFjSxLmHzi9CJWk0/akpmm7DZ0KPeK1nWjYl6JibTmOEbmViR25CSmyAZyT4H7wQPV
LfJg4i8hfDFNDvLViIz64iLjszYLJm9tmZI13jZjL7UpiQqUz4YKJj4vTImsliVTlpGV5AVGx6Mu
03EG1dQTVpkYzORagz3Dt13WjsiNLvDxEFS7uHk0Wlld4lLPDFxJO6Xdl6nt/gi3DsXsjWfFsj4n
j61pLnPaG4UNLx6jdQ/Vo7HR/OOIh1RonUUEtMjHFfQ4qUPl6pJBYTtebDjCMPWaubKmWItmu4te
lMBT7WReX+JjBk4+9UI6u4BNrOQ50S08wkAsAjiFMQjokAhrY1MVjf4r4+ImK6VsPAh18WpnhOkR
pXVptkH1993cDLKidDwm1n76h9UrlLbTtCkOy4sso6fAElqkVLVEEsQcps+0EHXnS/Iutj2TPsou
6Eh4fdASqSEkmBcB/OB8+Ysu37JzuCw97RZihWS4DT1e4h6hlI8R7Vo+A6Cozp3I+aGYlJC4RjRo
1bGXN8r6/D7hVPxnjjyNH6zc0iM0OyiowIhgmhmOXH7clTsgp3DjA9n9xbr8pcXGRsxYn4r4ylJk
DjcNw5fpQ/7aFJgLRMEmJeV+ew1XijgzW2+ggnoEbVF/K9TgOdTgeeo69GMvj6JhpgS0PDy3gC1x
NIa9otLhhI/drLRadPa4r1GfVh+G876wzM8Fm6ar5GrVas8cru0/I6wO0v/IM4PjF1G0gfiCyY9n
mCjzxTUx9CmdsbZlfnOziFvrF+xtU3Lwd+CYf+r40VAwWQyVivZDSTeh0XiND8PQftCryhZ/b1g3
gVTeP0jUUrIfZL8o07IGFZLJSMBZSEzu0/Q3B1qNGNBXPe8/P41yTinOZBwxiY49/iNpWuLpxxNt
AQNXkHrN/3HqvI5G7koX9TxjbtQgowAzwMhsnlrWUHibbBafwh7HbbK5+T7XDFVYdypljairbCpU
nDu3qaTf+ytmCJsz+4p3zfKWXp+NPkbaqTdIgE48iAgUJf8kNLYj9UGChgpawh66wYAQlSUzDzGx
7UKaNvnNEFcm8l3k553f90Yzl04IncvbdTICRNJH/0tBh47svW7AM4kZiOt1aRVim8QsoyvbQ3K8
NdYPdku6zQex9R3za2sznkEyY2IGjZ8477Eq65UCTzMnM8GtRBC61j+y8dD1t7gdzhHrmuwhBeMF
0PAAfP+AbTGrHZCsKWxzmLUiDx933vGD4rjnzbPjGEiLXhnWdLKnCObfn9H0vatUU8FoNEITNZAI
99z2P+6wsax64akGviwMMbWskbGNso2upkYMp42fCAG64s6OGo20hFSceu0FCGCbNCa7z9mecd9A
W5G5YYzHGrkQfP/1UYTMuj9S+OJrbGdfygV/AS48MWfwk1xnmR805+VNyugXtsf+cxZZXEj176tn
JdgfJe16/uVQJpO6PoAbGBDSQOf8Iy9A+b4FVg+jQqbiO9gtRp3oFuNhdjtshQu3AoGp6hBeW7H5
KjsIhJpmO3Qv2xZzEHv9rTQuWHz+jWJLt3baBg4Q1oZcngTzsmLsMX1vX8pcd4oNv9maqMJ/CKU1
iSIHYjw/uNjyeVzv5NLwKby9yksIkUrvnliBLeZx3nx6M2B97twRlLq96+vBiLEK8WOdY6CTp03G
Lv3ZQrlo6gWEbO66FMZKLH85raKapCYIifZnL8fm2R+e/Gl52RMDJl4AHiARF9sWq8x1RxdQlj3s
RhZBmyu1isOraEVSETVfck/jc/Lmi0uexQhEVtvFVmfF6bHxHholcIhPTCekimMry3M5gr/YxOk9
49RaxmLW6ILNQTnIZzXTc6c+iuaWVKx22WdhP2SOutehJ7ry1TTM+bqEAVu/xMqOZJh6LY9/nJmB
ZKpZAuj0j65E8odczVmaFMiAYH2hrtGLW6DMuDoUjd9q6h5rjQwWecAK6Cll+7X37giorgyi3JGu
i5jchW6eWOZpGamwp2BWh7OYghLJkVe+rrIyLze9+eiklB87zQO6N4IiUGirtQ74qnBjA/f08XNB
IziIiWrMJhKWp3JwrGl+vsvwyhaii6UCtekb4DRXI5TjbkijBIdJZ+SinP0ArhEb4zaw3p2j5qnp
6DDDtzrJYhyEoZ4GuNYyBg8bQ6Sr8C/t4orKS2wp81m58mD7oUpVm7SPdanpZKf5jmEcLC9NUUJW
N4PHqaL2AU2O1TKNl8jAAjYUh0elA6f1du/pxDcpCKJFxIsXYwqEWXgRAmpOICwJ5m9Bmp3/GAym
kivPl9aXBKqfFy5SBu+OqJupGnTvaIigCIeFm+yOvDMGMV7WWkgjuTJwbj7dxKIPrAulnlTWU8pi
yUeGQfttEPzINqUnjWQDF3QoyQBfhR5gYTZgZBcyaPVvRdg3a+412l7jRyOzlA/ySOzN5+uwuRtu
bArHjvTkPmtPURWZqm7TP9LQ9tKO96/eXl12y0ZZYUxy7sd5rqfLP5wYszvUAonDXPz6OFZah0ga
OMY9VCet4TMpkBDFK8RT5/uJGU+HpPUPv7JF0TTLz+RHL5vUOwd9vnMBYXaul6A+JO0c71pT+lRo
OU+uZD1u4kG3ZI5SZby3m7vortvWX4FdyBaDmJvmKieaGkr22ZzMdY+MIxLQesfDE0wp8IE96WvQ
zygVlnMOSQiVDzHHJ7UrrmTTzGIEBN6SJe4HJ/F7aaf8ZILBEWHxM2A5Ed8MRjdX5v29kYEvaR+9
Mwk5doHlPeK62KP1nsz1GPYonKBw3rJ3qq3wrIKoC7eJevlPbI5veVc9I4Gj6Oj1o4tKAUvuqpZy
hFbpZQ4Z8NpE1l/7MqMTor6hYFTsJCaXZ5Tiji+HDJMfEhlsGFLframn0vvwQ76lYdYSWFx83pPO
z5AqsE44DH36ZOZbsaiNrG3h69CSv3z5+yqmHQaEE1X0c6zVpBS7qG2jIYMUSN11QD7dfb3z4WQB
pAVC/IYBYRm4gGkPCBW56eIegrtiL4mYfGPkPqnMdf/dTwA4fUiasdQt9G8li8svTnX7eIzwP/F8
X9+sO1e7hWCtns1z6ip7UFn7uhvEl6H84hECtmJPmQOvJQB856J95rYOALm4n6b2G03lEnP/W1yv
FmB7KPNUCvu+Gp4YqGpZ7sqZnSL82UWdwIfcLAIo+ePlAiAqkJLFtyo5lJbnfeGbV/txxwB1AV0S
g0pGJxsVEcOt0Ot6n4h3ko2Ogasq1SLvB+K85bqYg1NAzdEu6/agWMb81mMflSVSomlUN5HZXbLB
qYwksud2BTarX+GsmkRtb0sH7KkFJFzAF7c6PVTuEOyZl5jYHvAmP7Ap5ra0hlm4ZxMHNDLa4UPM
JcbjaW4grib5XVG6asiCw/kibUAEfXianNZwG4cHNJuiWskq5j3ESqTYFf3YI6u4X38RAEXcDi4d
Qm73pVrwgqzS+dxxYjBCdbyWNexAXdqOZ1RSrpSEQP/+2cVYe8YIcjY7/8R0zfdH2nKb4NjogwSE
h1LrN4cXfLLdBp5970nO0EB+isOGxrP4q2C94irrh1bddBgLE28eW3HeCNhoHWfRExWwa/Hde6jO
0xTiEI0Kg6bmZazDnviY57RvNDUtn0wjS2RtxkG24F97vjg+8MhwAroEuF9Hh4d2qoOmt2QenRjw
UF3iYeRVWgs1NNb8ESOdXyI41UBaJ0w9I1heaJ2mZPVukiR/BSha0qPiQQ6qDWOo4Z3Uuai5q6dp
9aRZsNXc+K/JLMJ7NZ+0z/zZxqLJr+udZgvKGEP2Dcb+XAWEmJE/PwFHutDZGZ0HTTtYVHBRKW3Q
oKQG2K/kc3A8MfBvcpsTIkhSaF/qeBY323lmoJ2XPymrXIIgVIZbpxVqF+K2oBsnxWB4S0tQnxfc
Xt2jVqNRRbCs4XT/eE3elGazBQ+LyjOm6qF3ttBoW3NK6lqRrZ2W9UyBre1JQGRCa0psmxhfDLKd
4ClFnunpd/u5h3h8KjnkRv1ZcOE1uscS5p2toKIOXxsd1IYECNCgtRdEjXuRIw65QbLNcL0fCkR0
Z+lDQW9VMTkSdHeJ2909o11c0E1eRYiZVh2TdnlI6E+Ef5mD2BqLUqtcqaM7h3/7UcXMYsvaK/2t
Y++7tpRGT7qqok6GYEx/2l9oiMUKo1kcWsTD31cCKUrdCCNuYpsFRhN2vidpn5gjK5K6pG1QuofZ
rKTZVeXIr0i/EybB17A0ZoFNQ/3lmISV59d7yGIh1I/UgMpQ0H2b0npBZRjLb5dz2bTvbqNL8A84
6vrC5k8gonv/94m8iVRLfV5ZRacbsWS00T8s0Gwc+vtSpVqvEsm+vYaThpYHWH1Npn07fK4UeGo/
1e9pDdvICJWL0ZuDv9CsEtOi24qIs38FEate2fwwwjyF8q+4qGT/YqtzuAu7pk6rgfk300zIil6c
K18r0fIxLoz9QH3KZvnkvUrJ9SVoTqpLHW6E0EZ1QptTzMUmk3KOn+K8AIJBpqAljv86QRSwiU4l
95ZVvi7YvfESbHHUuPrS7HLK1qs9enoanZz+4gNdrMWWbGoDEQGfPGdONJKUoIWa4ZosZJfs7q6Z
IfUBzbPqgnw5fbYWP0g8Dr/sqY8UQuCm7bto0tIVKubrbzQDECVRWafvvq9Iq+IxOoc1Ndws7pwM
SjEUSzbkHpLjWB19aDEuZu84Hfh45zeDZnCa94+SgEJJ3FxtbWp4e9QhJeowtLChClcdl/rV2e7W
x2GrEX7HHRS/QRF/l8wq1YKfZPfelMVmayR8/WiJ/fItPByScWF0HTd3AlX0M5Kd4XJYrNTlDgqy
xslnd//eAoCQ3X/pYVv4Uj7yWOxvKrefBvrDlaTco7mUWsypBuBhB2ClcYvPKbHKHK7kkj3ZpTuV
f2YvjcqFBHAYGDLdC2zibKpAXy0Rdphg2ulAIDRTxmVxIzbbY+P0taogVcaXpOxr0CLbFw6gqsI7
HlA/hjlGILpuX8+iAYv6bfQMP+iXHJ5G5eQa4Olob2+LieTImUWYbe/oW09uuBdTvS5XK7OazfvB
M644X5WHT0oCdf4LPkLqMEFGwHSwfPu/PzmKzgj0nW1uCKKkDRKEDta/Xoq+CQ3U1sKPB0eNNvyo
wJFGJDsLTCDs9Pr3Gn0EXTy1VwCPmqXU4gW90H73ge6Nx4nOpp6W6W8/tj5wNMg9v503bvO5l3F1
xusUmoMY5vtz9WVhOJi9+HQSdo2wXHlwWGiarUmpSp9REGqdvOBVW9KaS9Tc+uFE1r1ZpMRwHPcN
oVsPeb28SO2lwPjbilkbsKinnzRm8DLRiORNH7MyD92NXJ7NdfEmQAyvguajO95Rm+LTJ7RolSCC
Hs4uh72rx2Pkhu7jPps8V6QLrAqFmxPMCRN24rFr/wr77NML/lP1kDU4TFnKjfQQf/5EGuUbP/uh
n4ztH95JKhR0A/o1wYEyAnK7vQruiIOeIjrw4e5feOd9lZGuwGgQFF0BUTWGk8dx8C2a/dhksNy/
111LyyX2PevePcauGPeILLxjFY1UCdWNQOxEE3P7Effia3CT2/g+Vz6aM/7GPaN3Nz/MAP+OApZf
zQDKT109HPb3l4zJt14C3LNOtHb3ilk0UMjWnGf8n5qHCrIocrVlfK19BwA+ECAv7EbmXrCYYEy3
2m7ZOwGUa4bx7Vj4BzvQ/Qaw7Q4c/4c73QFoG6X5FVP64nT23+Gvp5HsHgq8EZvXM6uEercp3AA8
KVZmVKRGSSzFZpuv1LdXIyydpe4cS2tXPf4YQrWYjI6Y7krqPnOAIwMK9yh9SMUJuRL47Wa67dpI
RNoTPvlM7qRVnw2sYpGNwGD9U0pCVZfQcrMW5RdW4GKEVn3oaX4xb4CXAYrSineoaC0jnmaCGYwV
3muMm6T875J4Vj+BMZCUkksQFqUk40V6Be6wiQjANDWsZBmqWiRPQ53YKFNS588ZaFvnuVNRhzFg
Drf3tC45SSMgdO+JjsoxDMyO//A/wNH33BXEO+0R7Z50gldMDdk2BgL97y+fVy/FEl5Y1zbUByIw
/EVRco2SUmqIL8AGfZ1QbFw1ywBDF0fgSNCF0gI3pjmsFTAApWrYyYoDFOvd2jY/IGsHm0ynvZtw
cIyw5MTIqAF9AW14rnY43lZDzvyrcPFOFQ2vYAOb+DSKylmtWJstJHdOhiwK8lqdvmnZE36noL2V
msL9wDDAv8Vr9YsXr1hVTtOyJGl25xSWesFi4m0wt1WETJyVe2t34nugeuOl4cgoyDR1nS8k30AQ
XV6LFCA1SIYWiFNs1uJEHqUYEIg5Jf3qX9+teGbpv51ayma4F/Uc1s2kig0t9RTcFbFbHxCvFhPs
z10CsDpyqb9D/EzXFJhLD8n0kbtJAQ35SuwK5cwu+r9kjQIYJ1ragzijCyuZVWqgDQHaMW0UCT4B
NcvKaia1h7E9cbMgA09NBpiY99Z/tznzHHAJgGrZrcfVyA4YrddGF7vaSMObw/pNfAK/4DYCa0Rq
7MJ2dglLyXR5EYdpnQ/ZcCANsTGxgaci8NnUv9reD+/q8+piUCPYI+4qqcW5m4KzH8Enr6MvOr+e
IKVIteuUDuAzxAF4S8MLXkm8w0AaNRid4zNb5aG74Ox0bolAtHhmtF3g6FGsc+K1EOGxaX+FCLNK
MxyxKADL/yVoEqZ62s0a5nDM4JOn2nh2IZCCHx9ir9hJilqZXUDFCnDu0WX14HDJgpcSXcJ+lMV7
gKkQbOHpWEJ4Wcs731KzHBlvB1QBmBpA7nme9qcM3EZNvCszJ2uiMgxSOFH/w/2gE8KKicXrrhac
E9DPycKaljJaLFWdlsQncZTZsnFiEz37F1OMBtHsmYuoeOzgY4pI2PS7dcUmS/QHwT4EqVNTqt2/
5+ssGHVoT3vsvPPD+913TKz8FgWXe71x09Y82CJh2U83MmGTGoxDngzd96vrT9kqaDe2SLMsDcv6
GrDL1HR2YGVN1KsjJhyzfiE8JuTXR4qy6E1pAWRkeA/aUzqlBe1puJnGmQAxkIcCTsBU7PGzuCap
xsXdsQk6DGoNrOxcRC1biqSyjeD6zn0I8cEi72YcKMuYmVOkB6II7uxr7QnJ13g/WDbBUnXevY8D
ujGwviEznUOZcyJRtko4gOVOxGhFwu2RBQRKRTnBMmgQFF9QMuJKQn5Vp9cxWuBZ/Dou5/rFnRg1
rE1jZnXti8YlPyKp2r86NFHWjFb0jLehq0lbQo+enVixqS1N4pakvvaeK4EAdNTs+/ZwHNbbrhEV
NP2bOnFW+gorhKa/3GiLStueptoAlTijnskcb380JzBusdt+XV0ZasSg2hhuft//ylECSf1cIE0o
3pGLu4pexmyT4UNkKC7jJXu3mWrFy4wE6pRUOVP2x/SwDlOjJo6QHChaa6z4eHD5KSpRUoy6KKpy
EErUVgyXrH52pdZSuA9puxVejTe8HEOGSkVj3p3yf+H4dTPKYpT3LZr7OGc7j36qoIWTARVnWVeq
gpsW6IEOHtJzrNgn0I7NkES1zONsi/DdKQGBaQfIqOfOcdWCrBN7ZywZMTwtORMOGGjWZD4kUCJn
k4KOE2R/uTVTPXfYp9F3EGfqqwd5ngph7fSwL3YGA4KFKu6mtfOXD49zaJgyaOZtxX9VKeYxxBon
x0EjcEO1rNTMcSdNUlzrhr/uT9JGQ3oMPVisn/oSDPJ05pCPjdQ0hxl23u+z3zYPhDgvn6kmffzu
TV4wafxxoRKSjniTJyY/cpheIeRXBD/XmnYkcySZuQjmueBcLbsqZ20oC85Fb0QQfpd1HAvoDYwI
0+akryRrbOej/HzQHSQvuQIXRnV+SiPOAG7WpDgzkspdRTONCzaVcMOiCthnB8xDX9Hdxlq2QoHa
NCOs92+SU9Q1H6epIgcZ79R3GqW4PfZBExS/3CDK5Bgmhe689v88V3ASb5VTRvPc1A8DPyCJGHzh
qAceT0oYEnkuZ/hXUP49OvRdwOy1+TZWFQlju/afkizSphEkaRqfTFbgcP6vAeaFFx4HH+x1Zm5S
i1oe7aVE3Hl6ty+N+dpJNy8W/jruz2lG99ZHD9MIkcTF3tL29z5AZf0UM55fAQs8mtweP76+oELb
scwwU4paokHWdeW0cWagH56h4xds9LCvBdmqbPoKy+FMizjDrrmYsI3vEwds9phqPOkbtCTPfL/C
R3MzEFUY76hZL/XVvlL1LA36ttL3dom7eYRUQp0SM1XPmmloLzo0pND8iwcOaIdX+D+IyCKz3wSB
2yp1ll9tJ35auh8V6AZaVGjLoyDDen5d8+nzZqFEsWPe70HmaYSzv617vedYzNeUd697daHNq794
+o9JziPElsXlfGAyouOqVwQRo+fwZEo7Y+W7wsSxgpm0Sol6A9UxxA4eyRiMLmDrKivEifGOp8li
2Bm0bWbCrt/U1IsaWkiJTomZ2RzLG/QqyokkoerwlBvwFB3Uzkt7scC/2ruQukTAavBvTifxhF+r
CLFLkH4HpSheCxFCTRjov7jiX4w4XAAv1PB3qmP4HZiPE20aJwQkRyvICHqzPK5NPaZWBLkHr10R
uaG8jjChVA/sFR1ZRdFkdVdcK4wowifC8pf7CeBOvU+6KxwyaknI+oAi254YQrVIwybjeCJPU5E1
hy0tx+ukxKsCgw+JAG9U4Lhhls1ZXXNH6zITIuIWefHdTrN6b4Vo0nYHe4U8GQbkjm2ouVtVvWvg
MGd4f5+q0iDDxA3jClBOkceEG9XJO0Dn00mw77Gza2mCKBMOURoimeOJ07s5xuKYRS7D+zR6eo2S
V6naQieEsEreuzjLDS3H2hWE781d/O+U69VhRZC+lFiy8EwLSpolwkIqLvVHJ4PcPT1N1iOJVkKY
wTm32rglMLVPSBacNYzUhMQnKiTmAPQaWu7UvBQPAkurZaZIn3/3Ar63rsM3qTO6jUkyb+DpgPyP
8uCDPo9ZH2Ye3mV1M7Vex0v2wpWlo9+Dne24jduJZ3p4i9a+LJ8efvkpgWddWWUC9wFG0qX2c9bh
QPZ2HYOCdO/CyCJ7iWRkMlfbm1jkJWaNmGJ4Z2wKIozKHmLwV5UFWrCDMkLKy10P1qX6p8fVSCaM
m5gPphQyMdiYdxrnTZv4XtVkRkb1j1K+58RXwdsgmSxL1glueVRJi5ayCn+3/PF9QBIIUQg2Vs6O
h8HmEKWKfefjO4fknM3T+oPH+c07BKLcsEE/DBRegujQc9naz4+0W+YZfZVwiXk9dvbB/82nQn4g
fGVzLUR9j7AkfVUboo/My8YGKzRbRtN7e5lPKLppyXgrVNYGT4QMKVjndg8VZdI26y4F6wX9QMH1
X91EXWOEOZFQktrC6HVc83pj9+93ISSpfXZkuyPmD2Oany2e+eKm4/4TSD8nQgSnIToUcAUKce80
eyQoohO6mk7qxOz7t5wa4iwvSatqu2UPUT1+KxWLmjzFCxAhv7o9Zt+u3afDcU4Fh+c4WrV83scF
UuH4NMrHJJ4KmNNYu8WPHC1Ll+yaWwy/AAcLtfFzUyXOMesache+6922/FbQlrlvMFcqo4xUFHfP
VlcSHXcVE6JgUDIesIrEC8w00d9oEGx+GssysAtlKGkLATZ2qCL53bItkDGN7R6M7Hp7o++Svz9E
aOto1UtIzhm14kqXQ/oN/bdkhRABy843nAuwqomxo1m5EOW955sjCK+RTLT93+v7KLO9vvSk2eqr
m/CpIDzBvp4JcXLv+jkX7qpZ07sISQ/9JLoVuuZOsqabw0PZcu9NvFKLXZc13x6SZugnoojEEUk0
LMA0pWBW5jEszLVGromGKdaTG8nqM9zZ910hzNy7ooW+CM39Albynen18lV0aD3MRc/h9+X3MVqz
zAeSOaI67ZCNyMlgQ3pnhCpCrZfy/DRAP1ZGV3VsJw39ZrGobI7/bDKs/a3ommgjzDEL+8QQ63yI
3lHroUi1ZCLRC2U98zSYeTGUnPLOx4nZHTsxppR974ZuWI5hrFUhmbM8UtFPkmzDTg8yoiym9SP5
1+59hH0BuvHxbv8nxh2BRVxvWKUH2+IafHxI0NQeHUnDgnXtxDjFzZkJrhY9zEkBN1V+3E+6Ne6t
IQYKxqACtvgODkDWj4OBCpOIA6Bn8m2PdMmaHQX4KmtWDDQ4jPLpAQfvrXRthNJGwV0BTHMiTNnT
DXHKRzlGs7HpE9M3GwgJ1G2a4XLqomBJSIP8PDzPp9OZs82HhSLUsfKZZGvcgKwxQ45a6irxt6MD
xMBYY9/d2rCvF7DH71pEDklLbjDnZol7uMi5JOkolsl5BDcM7Nzv2HQc6JNHTo7uq3rRH6AxoYri
u8/RjxfFkaAPtTOL7RI4zgn6S9LfBYIElioe3r4pB7UOGW+2NLD0cO0iIGrK0GVGLjXIUkAovRCK
JUqoSvODvsb5KALYtM10Mf9nLGrnks7Rh/sagn25ThVWe54g9riWyyy53UEilQO10dBNKRKTf6GD
XqFSHLn2dfxYp2G4+BKAwYHtFWWJ9fl8hx55gW6Mpsg7CJsWADxih9nfHcDboasE7OlhhHKkGELS
4zwE8tfiTSirCfLosDAv/zJN4FOx+/MGWY94O5lJF9/Acagqk24kqHFNAA2Xbp7bnsuRuxNo1kDV
jeyi1zZM2qm+S58xpLfbQzamr/yEOmh3HCE3Rfu+3f0HibVYz284F+CkBh/rQba86Tm2tpPa6wuL
aYXiQj0Gu/a8s8Alm6uktzAxogeKNmGlh6v7n8x5AV3wmae4pCEw8LGeZ5K//Dwpt/VnZuHxpKtB
/fnQyZo8vUny8jD9P2e8fiPv67dEzCLEe8zhsjHGO4j1EL3dHMs1i7vsDLdRzhAvA0HJFEly0Uyc
GvP7ZnGKb0/PjffdSHONL5iylsGw3cs6oshS0p26pPqISVObTOl3VFu93lVrrAq0iNyz4PHgvTvy
0tIyQvcxupUUJTI7W9b5nbOJFobze1vMSng/kPSZMbv/Dobz0FM1Ye/Rk1w0X/tC4A1YmLZhQ+fL
hJzNVTLLfev8lq+Fm+d3c6CV/XKR4MutFg+bqqJA4EiJn11iaoq+ZhDyhPmF9d7Z3c1h8Kw6OC16
2QTDza3jMaKhQiOPizQnkyxYUkgUDVeB03ON7JHeby6KvVZbE2dA/YK39vN0GlHCn+dLPfx69qM2
PekJbt7GR5ss4dNJd6pSEva9JHklv+FsBSURDln3BS1oPm0foSGDRsZmc2hbInbobJb/j/HSKzT4
wz+MbtgBdMo2cMnbdnwxRX1VIaU3BlWzMEuWnaixdQQOIjgkuSeOfTQaJNdzwYofbBCMtAlrZAJU
WDx3NhTBe1TVp83c5WA49AeXZN5p8iensELebY8a7+CeQPh38BlzEeY46MXT2PjHWHXdsVcajCBs
T3RyRwzmxLPBCUKL0pBXWQofASRQugUaQkSWhRZff67/hUJsLPnHm02EZCZzC+xquMxAnG9UdrfD
gQJtxMpN2c0ctJ2KwFqRrQ+BEeOXDDKylw7GMRr9OpJ5C6z2PA3jUiHqhYIVCztT8Ww8vvF+36sz
ofLJDUus159CzaIwVAc9AnGQk8mzXOO7/DzFuMoJLk6tIjJn9L0BBCythKoICA3JRhk4FRe7/cB+
FEFlfbfjc9Qmdl45ZmEuikYwDdVh3FSwS9qu8vP1PUzPG7RkOCxDDat44h7IAYDWePpVR+jGAg7W
i2QNqASIsFRYVuBfyGth4ItWwN6s6BBmEqmHYTaRjikV52rfb6RuN8twdDSXEPUfM0JCVQuSstw2
Mx28ACGfcCLdmo+qxwHzkJOMFW+jwyWUk7CYe/rfioBQ2wUCJ12nS3deuQN6nOa5AnLckH1UBN32
xrbpm9MFuo9U2Jw6WNM8oF25ztgBhCiK99A7iGF8XF61auOisdO6pwLbp0ipD2tlnSfCtImGrhT8
dOQfYIJ/r603XUypWlXL1KTrBPk16GM0umfxrJEuwCfjcfwS5aoCp0+Hu2ypIRPyWs1Ehw+UaToV
QrZ6UtzHFcYwwUrZ054aASWKb24Cz7MB50Qnum1EDql7K9/ObvDtdyl8tBzOv2hjMAA8WfM88EFf
QaLhr1RJ73Sa41b3t+Hg8f+Yze/4aYJezhzNuOuRs8d5NRcCmURqX0cA5IK11EkuEp8aHqaLI85V
ylb0TL4AnJ8IzZ6++i3jEKc2E5k1i1K+fkvjlBxaSmIH5o7TSteEO9vNMJul5UBNR44UBCJ/zeR3
7hocDSQ0u/vZz3u6AVeEMxKzhPXIRFpmHQl6NJVnYGShKHRGNm4fT4IYxLUxHgPbXA7XyHNnFrAH
pVEMc9jngksfrkmNVpVyMriVy/xze//TXHcv9QIbLTvHZQ8mxzbntqId1o9BBNt7Z04yfTMUf6Dm
Ym9mnmfMQNU3ch0Nk9J1HwZF9vDS+p3Ekv1FuraIdYXiaPGHw+pqOiNNH4NM+sm/bQqEOkmNSlen
AJXrzTKlVTJP/Xl4BTW1lxwB/x5/6NA5axwCdOGqPN8rYdgiWkGV0yk5HtRad8JrrW1RR4DREh7Q
WLWvSYp5NStBkCnFp8MkHf7Lb2MUQsjXW2W7ABUlKysIwl67KsNmAiqevAiJ5F2UfYjwltrrrscY
6L/jI1308WDmvH0942y6bULHKDi+UiqB5EXbNlGRVKkwd/hI17E8rJGtB6gg4U2BR+UiZE52Tlrw
izqcZnh8ABOlpbKBZX9dR1Rxm39aD3HxqRwZvWwFszHj0b0dlsMnjkqoJ2qvf8WLESKI5Ef58fVU
9c2bZOxrmRCvDgYrfyHMd0FOm38gaGKpiOflHq7hR8Rm471QR2nRDv7FFMTKNKQoCaMY12xpeFip
KHu6Onq7xgW3ypqNUK2UPGDmW19HUNOxF/DiSPtLqF2+F9C72V1hHegFxgGSBSmo2HdeBmwzwoFo
Py2SQRHBGezSaCGsLafOyPST7LKqNRRX8cgEQgt34lh2eC90mdT/slQTnvdEsFgoWA2pwXMijK/G
pa3MUnVInlUa78t8w/aLqibhzjw8LlpNuUTXhqBO+MqBHIIOJFZqG3vJIiHQ2cPWaDdmMWv+qakE
bs4S5tct/Fisi6FXw88bAbMi24XjofMgqFgcmPiMla768Rg8iCFzpV3nEkuL3SShUMcdpng72laz
QL7HtuJF45iqxYyy00JTCecUTsQqHPvetF55B2KTSHHkoiVDm9GMPgcJo/PA2oWwxbKfnhdYwy5v
FiAEpkBPqf1VvNInFwbEJmzm71pWS1+WQrpHAe/gEBlcZXkABoZ+OXxWoC8bsOwBRAIDQc6lRjzC
9wuUwDbU1L3ja31IyGE4gmnHHZ53GrUGmwGabFz2VaIynKpE7vbJlxlf8rE4WtZWEg0Awa8LF38p
zeUcKlsvPHk88nOv02X2rmRqilgPI5Vmxb93plbEY+zzO4XWBQr5da3UFvxZf9MWztJLfJz2HQ0G
lDuw7J3DSDPgkGeIKgaCvUIfP3/4Oip7bKOSHknFoa8y3K6mB/htAW4IYqgOZ7zQvzd8wAN+1cgA
S4r9zVyJ10UYLh2FUpG5Lj5a372DcisjBxb3/oZO2nMHjbxmza2EeIL83TUo9ZB/1bQuIAEVzCWP
BHqrNaWAlIRM3CeDLhOeJgtQSpQ6L0tiPMu12O38SM1+axJz8jrLeELjN7SD0FpRbqRzEK8Kb/CW
TWXCLG+O6CwJldvhDcTp0rNy+nCMFJh7AAyREQZkiRgduVmC55WSxm7C1W9+4tR9c+MyMGnNh9QJ
o47pVlOqMFL2R4xARpxQ5gcbaEdcSU6CMY9Vz2tegYAKshD1bKPywQLWdE2lsTk7tbkW38CvDhbF
1siS6EBiyyc1gdhyv6T5C3YamcAiL/viaw9+yJKKoMQa2K5qPccKOC3GmCgpuEgD1VbxDSM8ly9i
R9pJamYloXOLk+G1+PwLh2/QrXikZjHKvJoJmvfEHtZd6t+RG6FNR0dw1yMOX9KaNUDmmbZ1grg2
30Xkl0siObO/9vmfcjRqx2Md8FJDN17QgyXuCRbCtom23gJzk2b0vwW0d6eRJtGikmu7b+rqtnZW
9yUbd/tsxo+Y41jsSMlEyR74CFv+ZnCPXKc5I1nKrUd04VAIN0rprZeFJj8dJmi77PxAs2QoObjK
rIuM2VIj2/c6kMYvmARv/B04zMTgD90ageDwvnkfaijF82GGFxXXoLxz5IYDg8OP6GEYjahHAvcP
nsp6rPn1juwPu7bIeLLC0BozlyJujG4vFlD5jIauZFTPUsw1hgYTEl/N9ghZGzBnl98dVZkAbBE7
bg3QstUngMK5e8qkKhKlzP3e0MKUfpP73Ju/i+Z6m0Jd8+g2rWdXA+qVBpNuwWbb50wHATrLI4TJ
2LK4m1nKY6yNJtqMvUuIb4Z/nsphFCwAhijdkW++t24wCoHPf1bdTAlST75c0GpKHvFPlP3NsYv4
RMUWwNrbWM7y+ZLZQdr5rjstCuEaWorE5bpmJeaB6CMGTmL1z4HOHQWS0TFc9fSseiGlHQdfTXoJ
tA8GhWp1VUy5XYsdmIEJ0Qmi5PN7OBrKBp55IgsZRBtDKr4pmnvAOTMtWetE9pRjudKZA/DbV7FX
XbcUmKP7wocYhdORW5EeCs8C8psAiVqevdPDgAebt7cMbH2W/2X3jIDNMUb8kcdqMDugZentXW/X
JCYsvlvk700rl/WK5vxBhZnReSz/TcW7GUHRagxdSLb4oISNwVRprfWwSm9GB+5rEH1eM1waxHXe
uzF3EbB6WMMdOcZgkcS5VIhIojEDJYUhLp6Qdfq1qxmBORa2oQVHy0DPFTuho3lKD4gu8Tb/AwX6
Uockz7JdGch6fjRNEKblEnd7mLRQP/Yy4Fx3ZjquqiIoZh+ePmZXD9dhUFVKJ0Orip04/02LLc/X
R53qyA7b3R7ARUmiyrufFma6nMnUlRh4PL1Vq2U0lSkr0mJv12/UftzSFaV0m8U6IvOkt42Y1+hR
0o1vMm2YSOkRmj0uuEiZt32q43pgddJdZ9h/6xeDkIgoj16VtypGXIFI4UysLxUWJGS9Na1E63cr
jVDvoTpqHpUA029DJIrftLIysUctvnlRNVAk6DImA3BMFR9rEAwkgzZFKEAFkwMOpHBGv9rqSrrn
JxPoMfrx/lgHOunu3MwE/40pECI4uKCx2BCDpZfZJ+BLPmyzaeDVxfK0vG6iLCG/J7BQ1/W14ry6
PLgu0bWcce/2+YWpYudkSPa2ixQzjV94jTvXkobEQ0YBmRGmuB4SKzvuHIWYCpF14wTpqNz3jL6S
egq9vqZTYAmtad1eKvLAWj3m8EkAd/lzCMiBFziERztH7spD/PtbdrprvYU8yKySpu4Vd5+J02A+
i6tzLbDSj9VdXPId7lreQPzbgqP68ycxmjDnkJwIrGBk/CKcVU5CjZEb+cfVRNbuLTipRWKE72Z0
jyCoTzkXvSR5S/2nyEp42m4yr4c/s2oSuNTr7fGfbYcioxdhP0zcP18NOlmL+I/ixswZNI9EcXIp
36u72NREMv78dRnH25Dekn6iPVNjuQ2825ojeZOwRlrdkSHmIyUF/1inByXh7Wzp+4faVh1Q+Wch
s+CTT4/OtzxgdTpuyPJDemrWZsy+WM4UjFlD9CIwHlD4QJClFKLSLCSGi3cWRR/Ng0xD9E+O8GBf
NQjS4OAulb8mrKjAV4DcHUwCe/H0H66g10VPZ6wrctF44wfR2+aCss9F+zoNPWHRxTdiI7WRR/Ol
K2f+Ot9N0yfE8OHtZPA5agE6/RZ0zRYYFaf6I9wRtthSjQ0n0EucCkXYPkZ/f1MxiGTk0bsy5W/6
ncKNnirUAmvbaXI4hDAO3hCe1TRzklaRwyj43h4wVIPU0QxaVuwJxi9GcSnnv9d16gHzaExJbIJ7
jwkfCHsj7oncVG/E8CNnj+Vk3fx+rToLYjw+N/OQU5/hop+HB6mQQ45GvgV7fd8Yi0ZrYan80/BP
4c2GWnLePj3ZEq9hErvK7ryNmksLKfbNmfTMX+K9rIgmDSRMX2twxOK8JT7YsMyLqeMtktTAAiNy
Whmx8NAmV76nby5lVEH+em8+rNR3g8q/TyATAXfIbqxZjZObVHC0SR2pRcBw5agpbWhZtISUaQDR
gyu3p8Poxko411bEP2FRjrPYOa+5toRef8N2/3yIINrAX2lReAmH9S25BYIWfY2+pm7LGXu6bxI6
HW/OXLiTdZhH0FVIEXkhOgnE9OtySexy8kIfXsSCy0Y8OGXlp3hMCOAyP0EdenhJ5qnrRe3m2p/l
WoBkxr5dwBYeWPv8sHeMO7SAGgHmqDA2ERFBjPLFe8g46z5SdZQznqsTi5xU44oZ6O3jpEpN8gHh
qNE16z8h9rpeID2FLUr3pGrbhgMYla/BhSu149rQHSowMAjZ94ZCaBmfFGt8GqNdO3qbpvxyUoKJ
fleYCA+He5DXMQlwSqND6GX52xst51iyKsy9MKZBg1uPooYUYRKIEtAs+L+lFx6uhjx254iIsEhp
c28uwqXmxJMhjI9PI1ls1OLOLV+AWTY/GNADepXS0eeuBxmfSeu8PkHvBWGLUySm/TKnEsyO+KT7
wzF7OZwNSdTjvaFuEVKeNmc8NS0FPzfrXMzLaSlz7fI/v0X8+5VrKtBlfYtGGwUQPbOLh1pec9fP
m7/5nrvoMRF3oI0QoRm6cyZqmr+cb02TvBCdI/SxZlZWHY4KN/dmA0h8WUbgC3/TCLy6Xn8EB3zo
hayVh/aEBO0Fkh2Om1TNj8R5Ron63Z77NzqYVMKnXixmdeP1MWSt5XFpiGcG/HBE6M0FE4lT8Wg5
zVh1pDc0lXg8wsVLomZ4uRswsq5Ac9NJsv6q0SmG4CRHgH7/BgPu7TRu9Bhuoo0YTkXqpJ9+OIKY
pF0fRJGsunZdTakDOzGuHOgnG2NdnckLxnDm+8MYQCp/cAYKbYnx8NiE8CXl+j6SeERS7u96etWb
aiUJnoTLCdWqZXY9kUJit7H0iDTvviu+Z4SQe7Asmplw7Wc3MVSMGiTJa6e1szeqDrKDeOeqaYkq
Qkj0DmADTYVLobJM3HgvTjLpSh18bev2a4HYjMpHAaOdheW1yD23lFi0+elXCTwj+xE2GBEUk3nW
4PSkihhU21lrzef9QyXo09BwD+21mMTmEp/A0Uf4PW+n2OnNmco4W7ycDOcozmgfk+jWY5mzuHwQ
gqXxsWHoT0NGuI1Vt4a3qluRfIs3z2WCCytnFTzZKxkkerP8Bvd+ERXzlsVrqaczH4/hXZYm+Ijc
KlAPcRiSBd8TzaiuQ2mWIJHYVpskaLknMVS5KfHcJlBuCFaUadS2mYiSlV6zQcJK4yKnFLxHAJ/H
KqVF6b9ECEGgYHCyl0K9cEEsmGbIbi9CU+41qT/COPMhB2nUGTDQ0S+ISmjibsZAwyYQ/sRBGhFC
z4hy1sdMLs7LJiSmbR6iOmYHcFIqvh76ocqTXtXUMBgw8KNLC7x523BAD5UyvK2Y1MIX5FiHCWzf
z+vdIcIEYI89VK1UvkI8o217lZSSFLfAkZzkqm+oCpvXEEiClFmzbJFaVx8P5kaCxEr+LEqOGDLf
/Jzk/OpcWoCtewp5kqCxl41hqpAWwBi5WKYhiXyTrdBWtY7hIAhs863jHLv8rMdHUGlocn2r07HL
RxwWMp3EcQfENqBVG/U72aWXDKNhqRjb/Jl99LO06Q9hIAoj1GbfMzfO5fwMceGALW/PgmUBGz7Q
MlVx9W7Mmp2NnWXqzxkLQqGRrG8RGIlImgWrSrRWSsQRWbsouGUwtf6JmLUm0bW8NNjxqLKfSSi6
umUYMnc1fVci4u5G9MzMfDe6IW9Ixcr+cpwngvcE8+JcIKyrz67VbsSY3qkdUmJIRGdc0ngEkWPa
BnC6L/pJAbRmBzA+BUx5JWwwSJhKqKRGRb0RHKpNQ48f5c1r4aoTiv8AqWODrVHxdLpSgseB1Hom
4jjFjI3StJ5ICqpNPV2tOdKvHTR96+QeAfa5chzBdNV6CPGZCaDP+VhBEcf/ZzhT0/9wtPaJbH1u
a0ZjH3HQRjlyPF8g6va+nqiMrvMFP9NMLCwAv9cAQVBKsLxU2V4N5QkDsLGGIFQos6iSmiY1pvsk
wAqd3ek8VofJHVuwivORAnhyYJf6VlyJTlPkMtywKCvS1CIdQjQ/kNNALmDSkveDtqxPTIZWWRhP
VLKifI9O1CsOfPzxEmcAaGmZqnpwduu8lTTvYTJFxynWmEsbJzLpXzLqK4QeS12auCxiNBMnUkpn
J8FlCyoQxo3wtj8poWCPQemkSbZQ+ipurfbY8p0cUuZMczp5WIgwRZLqPId6DOynvlMZsIhMgCv5
X09dvEuM5KJWGGwSYjXbDe7WHUET/Z5ERQMp3MsiX78HnyHKh8lVEdlH0IF6IszAhuYBpTXzW9ZN
oubc6GxiJrYAmAMlLHDhyw/XGt7gzRzgoLabj4SO07+TfHf9kdBzNDNhpIvjaK2yOVIBvTmhIS/w
nX+lUkaQGI0FiLMrj+32YcsMCwJ+CHQGHXhEBW2Ll0Zl27GVwH2S7BNwhwh2/qxpXGs8rZeKMYvd
6hCkcaU40kQKfWMjJVm1nez5xQQK2CX2GKWxDRWiKvGYhndwFDmV1lou4YBqJ5PQTV/dHfNkxWGz
8V5RoFcIKuApKEwbOOkIEmwKeztlVI2lFgwFR1C7NZje7LROwkH5BmicF06nqEIUOAOarX8au/JK
+gO6ZbxrzwjaPIK7ivAu7B8HNmm1C91eTQJhJbH/oWcDbk5/JAmsbScgEzv+7uxsEwYZgUO15bTh
s1nSFrILNjC6eTWeXbkk8O7ieeM+Jth/0n3RrlJMr2psPZ62lmSRmTJNREvxRFokJC8dxuw5cMLF
uMFOivJLgE0dC67JpJ47B5LStyRXF+B8aN1wBIwE94Jk5NHMB7Pr0EkQGU48niGVeV13Drv57Zgt
3gdLIg1ucFMVgJ8tusFraz5E0teyw1NtbIOPJuPUbXJrT+OuIJGPydm5o5cgIZeswICPZBu/k79I
rFEVWq7U5hfloWG+3GfJIcPRxveEI03zSPUADZ6oY168mK5wiH42/yT1PXkxhLXDwrZzF1/AWgJl
M/VQVlJrmOb1FPLMXt8uRg1jQh3hJ/MK6PKoI14xljpx0XygrEcTpjtrPXRcSx88MdxBmkQKQKRt
NhZaAIoBGO6DhMrn3SOynyms/e10ZxOSPdgsE9clpK238u/ysndjM4eDr5j7kp+bO3XvFFK0oBub
odBcrvXfJOmuylrTyUq30MWPtJ0GHzCxKMlsygbb2TS9QVnwWO/xzjl1WnmqhF0ukhTb3rdgffQz
1OiKMm7DRvBGHxI3DTxtHVFQiC9vDZHkMVnPsCsjoqM7UnKAWLroWgcywF5qHMgMI4SROeXdjSTn
1M16FqmWqw4Bgz5m6URsw0Fhiukle2vyh28IqR3RwqqEqAybImn6IQeBIEnYGGiUI/tzXcM/WfiC
1SeJp5uKw/1Y7CQfMgRUzhA5DFeitRN5SC18+2MmMFJCEkKTEo4XXCIqoN+Hf0XUm+6Db8o+gUfy
8B+VfT2taJApU+rQbzJHS4akv7JtriMCx4VdTiU/ykE/+HC/SFHdr2br7zqoB9obCWiBhyv/X3ln
c87eF3AQsp35B0Ltiz+PJahQB2zcBDNyWQvnvFztnaV8NPgE+u+FYPnkwpFCywQawn4pYESecdL0
EdNYJ23G4awEpTh9+nDYVcl4ZRHyYeB6DQiNga4prRuuMgERNI7BjtrbXxMqTN+XCkMspHNeUbY9
w5jcmqnIdlWJ3afRtx4bfuBKMh2s1NyA0c9Vc+e8ZBsAfvHzsuN85SY+6TdNM8Rna9X+uvKbpr+6
aI1LBP0kV7manOORGYzBPTp2eaaZe/kqk3GQLB0hIRQt4KNZERuCp0mD52MVK8stkZyw6GuRGfRy
HRzbpZhk4fQGPmcX4h8VOrvWGsiqEaKsDWim1akZm11ADM8lo/IgIPcNKScvwQ5fm6gYayUqNGKo
7DZ5Wvm/9hFVEOtIPBqnlYJmehleym+Hb1dq4vC3TCP2pzZ32dnUb44287/1TymvjZWORpzRm2SN
dcnC0zKZ7QczxK1qYnDAvxNGK3D7uoQ9MlIyBI5rZ9bDTU/nooK7bJsaF8Z9Kz9wEQzNbAU6VFPM
kTDfvR5TqTKxrMV/C/6pLsGqL/OlSb1avFdWrfJ6teoi8j+cu3dos5UPUc8HNhWeXAjCVJ97bnxy
wBk4NiQQc0/IXqMiMsbV9HcnVO3W+MXjzIC3MjW+9rUdOhQpCWcQOgfMGl00fgW5c6kCCeCso41+
xhmW5ZSKvSm+2UV/+BLUh2KHFeb+NoHHsMjybmny0V4NSTHiqj3DHm56f4Z52NOXzlSITSAu3YZV
kfXAbWnY5YxK3EQsFE4ubdz/Tct4L81EnNzh8U0BPZy0NAz9IGG2bZqjLI6nl9MUdBlvFK+qNZhL
hIxWuzEnT/Gl8ijSrb6IZRsp+0wdEY2SlmMXyBVONLWfywNCXUT360UyAKppejeN1ShMCbefgDQO
MlrcUZldnAx35RKC8uptxUBkncTngM+BTTS5mxL/XUh1OFJ3hpQts3st2ZRABA1Wy0S3SqisBPA5
JaxKMvuQdEkXrWKsFOfEJ91uqAnkO6mZxPqr43sskCEiYHEANM3S75UnoYZvQXXeaXE7ixour4jO
rVM9D46YziqPag8ukfN5x6Gvap7b2SdfqHcxDwV25qyMCterVbMBhtLeKX616Ufkz0lNoIeSmohL
0KIOZPlOvaNq02ja9vASx7e2LxYjQXWw+H4HWTRLI8vaZs1voCwP3DUtPSULZqQUuE7OOUYVlgbl
AQ84GgSgBmFwNnsZIpd42U1ZOoKJMIvAg5NlNzi7/bUvRLZ32Lc1OMXJK2N7EkHgh9zl/ir818/y
MOvM1cOTw/XWnri+gO4y7FrBiCSc2nE/Gs//uKcy35aei86uUGgtRN/2TES7IWBZblrfjHlpWp+g
glI7GCup7Gwh6QIT1p0SYSq4ZvOgKgeZUSZUbpmAXcuvgzN2Zncwa5Xm4oZzziRN+WkftjVUrZD8
TpUTl3exdRBemQq8mT94RUK8l5izhfGhj9QCDgkbgbB0bYrQIVZDcoxOP8hG9tTirfnlyBkvYGW0
YuXubZqlqPApN4bsTlnydXIxDK3/x65dn4WvjHckCzv+dZlQ/LatDNzkgeiz7wfycdGjJKtbGQf6
W2fE90IUW7qgWTn/67EdnRF0sW25v0LH4BgHkLjC53J/1XPt3PQkt9AJdWJlP9t5erFYsna7JyIz
1F/ajsedmREf8FmPs4CGaOzOEr+ZEW3Q0mdQ5k79//81EArNrepOMkuCERHth6g6+sfdyp4UewmH
vPFtg51yXJV8FL+uw4nfcVvfqc+JOduMtb2bPDIzQAURkhUogpYbC4fZEUE0vnCGb7dEYNX1ee18
ZfvNQd0g6G+4TNIR1XKL616MySO4dyh9l2CqbqknSYlkgc/OwFaq5nW1QP6D6K6HG3UaWQN5w0HI
RfsbM/ktlFitoX6QcQ/s1u25JmjK7+Gd14m4/Ub/eNZgkA5g5LYAOJRkB12kMBYGjJ9K4kMby6OO
4cpB972z0Oy58EphMgdd+FfZeB7tsX6Q05VNCk+pJFtUieBAh28R4nx3j6YUo54eG7e9AI5bq/mD
xZFwkwc35Qc6KujycN+ZkqAJj9bL9U0HD3XhcYlPwtFcD3/gfeZw2UBZgxCA1lI/z9uyFvwJaMgJ
bEFXq1CyKvKuNxolMowl3IEIvlxJhkTafzqTzdLd5iunbp11KERoeIw1Qk2dUs31W56i5Bubvhlj
G8H+WQiGimqQzZcANRSJlIwu5bfj+jWJ11gHBJ/a7vTVliinKFXsCOw/tXhqllT4BtJKYavdbU9N
CDYSnrycEayxQcTsMZ6SWXXgfMsKp74rdUdci8uZu19oy6vwi+73uB3rVXBBU7GHa5Qi/mrcrycC
8FJ9e8p3sEQH5EuBmWDeWE7cmAl5o+LbDwTvpFHDqlNJzuF94BKfpsvhQE3/zVCd4FioYvZp07EU
5ePPm3Z7/o/r7J5BL75MLthy+MtRKYkr/bEd+i01mBZrMsNBE3C7Ide+8Ino8SxV00aWmFJ5grLn
WrZa8qDXL2LGOHEQyIyzlhP5AEIhdP7HuprmrR0glLfybZFgzZYRBYKagGclrkwG+G6LtXOvmalN
Aq+Za0rytvOzoHWLFGe/1zZtMY+XRNZrRbk1UR5kQo2EII5QRgsvochqJ0yknPNbOxwdaqXSOWfH
nCw1fJIjrXDpaQZel6MZDtfLAzqJ1gCcRPMet2zPS+EZjCE0h9fae0ELFzCp/djqGN4Xi6Nq/lha
XTmb4Nhj3X6VDBi+0BHhKjfirEY3A/QiZdrbWKOtrnTtQBzq7tOsHd/tC4vxOwRi1kuzxtVFg0u+
vKk9cO0NLbwVQTvpqmMqYDYZQXGN7yomkkdkdAbBw2GO6PxC5SI37RQu4/l9iNOwIog1NjJM9lBT
TNYYJ9tC+fk6UCqZF/HGxqkyUFYZJikinA9WCl6VBj/KCGBoGTmDiE2Tmv+np+Vc1wki158fm4S4
7V7dhzgHSKyVEnWKQjUWG4vxqyZpEHoX9OzyBmUBt+H52qALmg0wTFlCmaeQ8pm9H96WFAWmBq/Q
WOmpyTzLCkoXL0zkionOYO7kI5rEiw5aU3C9ZevgMglw4XARIrU4Utove1mxC5ocgbiQovjBrz4k
ws7gAXraJCtF2pzPnp4LaVIGymOYTOoTG2f5kU5mFI3gCs95qlC64jK0iOd7qLci6XZM2bn3zvdJ
kEmojSIfu1H7Pz7kFLJp6jQOdt8O5NJ/QY1YwwKRzqwBi+Up5RLqcthDgWUaHwXGb3LFGcvoUazD
wo4et9IRS9+2KDIZ88qSafXaPY8m2xxxbAqhPALPKnixN0B0Or6Kjqi/gj90vqtENtw8rqwdcHxE
IyOGktcZ5WGV7xhp1/dcF5xHH/Wukio9VYm3Wv8rwAefVGKMcJOFyHuYxlRZZrMDZKe9sQsZeD5C
iUOI5L+h9nMLhEO+sU/mqdFBqVy+1NQJ5MSRTSs2DyX53sSAB/ySssUkk1pPStnVRhHcbRET5JFa
hBL0npxWG8wtwdZXxrjKr6Mv8Xa+37yz72yI7SfSSyHRTTtNwHVFKUQYUuUTUUQVdvdOfBHa8nRg
s8FCLdCyFywZeFL9bBIPdtrBdaBc4BmDOGwDN4J/iKxtQrHaCgYnlsN+t4eHJIuVfxLXPcKip12M
NGEBIKkMm0fuifkBaEfVVsVrT4PZ2f7/QXo70CCqpI2u3aL8YWQSTuGaeV3egR57SKxr+G1K+Ddh
Xttgykiv9ig3tELnCn36tEGIJLIe8nHTY95UBUIRhzgAFgOSeciBl6dL/mEAHlmBUkQgJt0ib76R
0+QJpM7/K8REPCMrxQKmxXlgDT2LQcrcCaE+f64aCrzcbQKZ2dsOs/TEn4PsHdZcnIIOBFS6VWoH
EY4GWOm5jwasf6nhFaW2/OVhowgaBc3D4eJOR49kVzRih9W8ffhNIXzmuolAFTtM/2FPnUQJr9yd
ZGEF0HHaqIt0Hz2piNXa8GK5iRS/ntR4CObxf7vUtLFCpc2etMktlFevISmcpEVhOzUGkjhh4q3v
wCvIhkokuq2rKW7aOaSRCOzKvFxpe3WOgg8EyuvJDdY6iygY73zEf27M8nmZqZUDcwN2p8jYXqzN
jMFr2wA60EVboDwNOINH7T5vB80YVx9eo4RpPGvg75HI1b0B+xEbAWDpjCS8+wYb/Ygr2rOIIhyf
pNzvDoLdn3H0qDzg1PsTqO9PCGbHmTP1rY5kxM+B/ayNmpZ95uS+nEqpMfuN0HdEYOUb8gmi9AIG
kwPtTj4UMmbf423R6HhuFOmf/Zuxp13/xAEFAd3mbjX61jNcXh36YaeofOu9olYpsANRrwvvBPk/
jB9dnIMyM1GbgBQjmd9Nk9w/QQfbTi90SMK6hSk5q1XcNXst3/51EU8QczYMDiW98ZexNl0Yj97H
zQjWTmXXNvKU7UDWyggGhxhU0cXYRgsVTHBXoG9Gm4M3yfsAT913FTFtGaxp5ganVKJ8WLqjnFAQ
r7+PjHfiMufGLsK4/smmTxxIJlAARzlQHXP5ybG1kDnnUKiUnTj0aUIBOVkALrsKJ+SDVRj+0KjH
83HU6RjwKS1M1+tq/oBb08uddB0xV78HU/Sn0ZwdtH0byOzUyrdYhPYiMpBRrIspR7jEXLP+KP+f
RSQZMnjQc/77e4OoSWf6hqqlLyq30T32oVj56WKbFur87cj9mBf0zbHSwYu/jbXbjM4NeJqNiP2G
FUrgWGprxgq1oLEIoFJMOODretsCpD7FR9VV+O60VMG3mJzNhOKpzm7xyAi5fUgotQz/ro+6Xmo8
DJNOIsTbFDbamtZ5FQlFwwHJu572djrXLl0fc3CBivgJ9go5oYKTRpVzDHhAO2Ai3h+UjqaOgG7w
iL2V4ea1KtZV65sJb4pEthZJyhkSsAYWfpoo2PpfNsDHkobnsaVoN5VgJs2Mvvhn2momC98mOh/t
6CAtxr7QNX9B5EdE35XoX1RO/XrgQVIlX84uRB3X0XGYSTZvfdUgXxI6BpgBQDycDhCxyy1uiA1v
ZZjaRAx43E5erD7LyRH9QUMYOc4QJhiG2bkc9lDFGwH3wWPR2ZWxn8lOTp39tsZTTL0rw1Tr0E/H
6TRZqZxzuMSqZXsXgy3o/nLtLG3RGtj0OwHYfjmEN3uWGzm88LFpPNKM9vmNC1nJuxC/w7Rtgtq5
qN3Vlgl+qAFDFOJ47Xj9MpUu9xAcho+0H+vEWSoQbL4sDgCQtmIOzB773NXShLm290DVzW58arYY
mVU5fx5inAr5muTOR0q8e9h8lKJxsFt9zm6mp6VswQiaDQP+rITU/mG5CqSLxc22nPU1lE1nTAwy
bRX0S2KisowOWEgpHLCHFWa4iVsuK85FjF//Q3p3zgfZigcRLITW+yvj6WnLZ95Nt3hYN/RI3f7q
fxeYZGoHZX0wc9f9W+7w1TE3BiP+p9gYjrB2uumXFkLkD2sh+EN3aPst2f2jrA3ySkzPy6motRer
Je1vLSGZs9g4CiRTyd/3T3h4VtnccaNey52KV+RYV7HQ5I58i1ccLhPWjvW6EiAz3l02TJIgCXqn
D/wHCZ/kcZMdduoTdJKrh/JvVncpgFfzuiI9JkJXd2ua1lMDutgblURWOUp2IeYjXp+3PFafumGm
YLe52xEgkuzfulM0sGDIYx+/QkMN3NSbKT/oMox8js0H1AU3y6yPyCPip1wQo/0jZtg65ORL1bA/
ezBnJQJQxodf1nIWT2GUzMNt/jiJ91+MSD3FRXuvrULBQS5FD5taF1GwWzzv28QuctUlzbqAHtVp
237Wn+sVzwQ7UUkAlLdrwc304S6qC3VZ9JKT/hOjGuL7IKsC90kEyz0qch0aEzHrG5V60LFg3hXB
Jz3MtJcenDIiojGn/yQfOCgNA0Vx0A8PCPomkQPT/nIG7R6+Y4ZrQL3AKidE464uu05T+6W1BXn0
GxZVrjJSsVFtlxr9n8GTRAmvQ1eWQNtd9HSBHcTdY7YhpapJ9gUkGB67I/8ZW5NwvIH7PhZbBZYJ
002mqZneI9J07xkSOv5i1q96sHJlVWoaE52iEcr8gjz6Vs9+6yCFKVsaNyVezfnaDGrux5cVP5Ut
hH0LwNr9t9XCWwdsSh09o/H7CKIF45I2nbh3pZNEday73Ie1isTndjJMH4jmcL7XjKwlxBc+wmRB
AEoIJQSoimnPRaU0vmxcFNO3jP3ssF0QB/DXN9wupZzEpR4fWHgH0kwRuGE1ymIRvJWwoyeZqElm
i+SWKLxiEs53Yq+lWZJZQOz0V4PRRI1Pfwy9uZzFgEgpj20WDpxHQm43ERq+Qit0vdpxFSHOJeep
IdEdgmNGrdz4Sbd7pCj3p8Ubv5mEfMGJDaFQPJo0IoAmRyzKzpgTo6yz28jqiu8tRbe8HB3k1pae
z9tPZqWimbrxZilM9/M+On3t6/rl+PQXkPTZHzToev3ebvLHAq4DhMDdA0J+47PaP9vH6KCgaLXt
66J3vAkW7BGyiTWDK3M2U+6nGrEjrWkgbY84P0KoegAxQryf8f3ORImoGZ4PfudHIB5zUA9PzVeh
/xPH6t569tUzHJoVFFbDTUgszBUia5hv1KWaDZ+z2u6CUsssYahPXpf8p4g5ytJvdqwljMp2JOdY
738WlEETTLM+xZLqGqv1EpANnYDGtaCJfAX5xLtE8NJmypn2P4vNxt0n8bwxGGcCvwR2W0GNH8aQ
gbRVlMXMRubeONlfHpex4/kfa1PnjgFD9lLkFtZkXsKoKRw5aOsvnO+LpSNQu87lIldvTOSXKPfD
YX1C2DRIMPyVsNGNOYdNDPci8AhIK6PapM/kLUgZBU4nuHtap7+akXTO2Gk92TRd2DKDnte51KqN
N3iSXlTsy80csrs0Uo97+o5x+KkM/xWrFl4s0Cq8rhvLuzS+yI56lbPiqAeIw3zjUa18mfWLYkOz
6pjICYmnPJTkDkeC4tNY4LtFQpwQ7hJE6AYwtT1XVKhj7AQs+csrln4vp2rI3Is2OBIAyoT6irPY
FwwFFCx1DzdMsbXfkd553cNVAMiOP4f/6EoJ4LsfLlNLiooSs1/ArEZordPIcJ+C2/B6iiMHbqoN
Wlc24HPfcqLCCMeSJZCDwDpCD1TDNzK3UX4ax9Ej+jgTzjBpcYSY2p8+pF5xgY/hRG3OG8Ymb6b+
Yv2MwNRq97xHG+r5IusNaL7AHR+MMK1n+asLxhd78MpLT0C//O6eimPvcMIeIami5t5Zyv5XYAeJ
KsPg9/A8xgTfIiPsGlddeHEu6eiFj8mAVrqyPQylBKjCg9eoFZ6sRRUSogPIJXojQyCo6phhjcSC
iTkiESK3QJjaqWaPn5pLKzqDFR7Un8UFQ64eC2GzwXxAT3Nxnzmk9t8tD15owl+mHFd+kW16E0Ip
s6JJ/+8i3mTQO5Xfq5tm3PnFyIkTGs1DoPN8YJ7oDN5OsnSpyzYtAxwgLUV0WWEwkpG4N1H+wlZp
GE+mn6pftT6leJxS1kooxERHPAwYLe+FYrJDcYlPMEtegzFKNv7/HIs7NJYAbPVpnZq4lz+Gqf8H
3A1qNpxDg5KcVr/8wCNxF7k/o7ZTBg6txGogSIa0gVPqD4KlPAYb7MBc0apCPrJQtO0rcwbF5KCz
qS4U5IdGrJdkzm6O20wWBT2WypLcd+ogJgaEtF475AhZaf8aWVLWFdnjhTzI6XYyPJ7FwvfRb+1F
toEW4R1AdhXrjic6zKsO0SZ4zA7FY5XPJyDwz85/Xupv8rjhBXsgA09TjTAj6VrfdlPWFTT139qI
5JTu83BW7Kg5xXUDluSsMCo/4HKrhlyJTE3dzgiCUYxhcRVixWZBXl3z0m0zE2iIGqYr7seI/7s+
4iYvtOKBaQec1J4Js2H6/Jzl0CdMraDafx3aAWyDOcJUzL4PvouErjt1xpFpZUR5CmDDVjemQWK1
aPAwtYv8cP70HiS/E3VxGEorCPVZ2nLde1sfFYJ3xlhyLoJ6Cu0h8iw9MoJJKiDbDGQigwh/iLlS
bdz+nsyi3j2EVyhd1e9iqWG6iZUiV4+SApHORVYgbnuFVCn/B1Tnruws/umnp9bR45wpoMhi5Emt
FCb2NQhGKFyK/SZSic3DgIxwPLK35l0xVMtZvuzVdMrZJyOr+HAd6Mg6HIX2FvFK8RWyx79xslxy
bjZA9W8PEgx1Ts5PJqRSYRTAPN+R29brEJUHKZb8xl3yLiu2ZJp07l/5xXwPPTeTmcEMxEYCHAF4
RVW8UZj3E0jGYh8R5piAioI1N9kWqr7W75rSrshmaNRIV4HC8ajcbg+6aaLLdukj1to4t5r0siCf
VtiVM0DEVafEPBMl/HRReKFMJrqLBWvIR4L9CYM+9nFK+1qiJcpv8D1lNegZNe7DSwXYhbUiGCWq
DyO1VUnio/3uBvExla9P8VcbDWhMYeWPLNRW13woMytf57zdPZiRzOr7M3A7bmzq/scZLssEoU46
8zUKUmb63C3QUFFcv5yQBRLzP8vv8mHOctvg/Gkf68tN+2O6Ib+1U9+lFS+fBblVRMeAi/V1rce7
j5t6+MDzE/gWKPUq4nD+0eh8H7fsiqgyLeUjcc4C9LqYTjx2vmgtSQZFX2wRpkN6oyg+JWp8xpx7
VWntpa86PKsLHq3f/gd7RwoEtX9WyyeMtxj3bvzXDcGn7sgEPkNOApy7lGDJwKUN9/3csNQ/O1gs
xS2ZfgPSyWZ3E+sREiybUpttjzsG+KFWeyeBBesECdkoofaTbAlqc8RqbMVlZyAAfD/3eNzWakQ6
xlh7dmhNeZCSu5Nywje00he5Fs8XgjStzLHPl2+RBaQ7vChQ6u8hlqUaZPAbfpGAUwGyKuQgEBXM
+Gu8smoIYrd1khnuROOQIAtsys/XdsYJyFIE5KkG4gLoVb35m0UroQ3bAbwxcePqFLe7Of55w7gZ
DLZPdvAGIn0aT/wqO7jvTl0yKWvXto0yKD+c6iXIkea91Ecd++G2O0ytzr0bSWneFwBd/zbghsBb
fB2uns4XoO8ubiGStK144ezmiC1R909ZYAllpLyxFNmbhJlSOc3v2Dr5RrKiqIf9mfZGAJACDeUp
csHAKHyRrtwWZdJq5hb/f3w36Mos4zI+2YFI7Z4U2OjrG0oPwylbkXYx37hsM78/rRoxa4oRWsaO
Qut3fHA8gZUK7z89uk999by1IGxrmN8tH5TwFGMX9oPTYAYIsNCHiszjT8yX5z4wXCaz2INRNw4y
S87vJhPLjn3A5pcYBlPSSZ5FXibSI5jK2S4F7SOKLeaP4a4fLl2DFoMI6lN0+8DXK6RI5rMQxe6N
Rn1as/2UNScYpv8wXo1eSuPQeFUIt7VUokMS/G6Zp3QDZNRNMlXz60ghCwQY1bvKEqw7QJX4/hJC
jpGO60KAPVrIN/+dnvqx0VZW6WpKS+PHG0aHSt3g6UFz2b6BgBu54ITZiWQ7DW7hQjvZM84xdSBd
sL8fgVmD1bLm/1X42MDo96yMjxzhtckFvoNKSItZVhIJg09CnUGhrnUU1VMGp94a9hAfgYitV6zC
zZkMNTav87qqABYR7iCA3LpF50RiOfvvJDHmNS821lmAcQb3eBhLHcuLQSYa2nAVv0hIUV4ASM32
iKoDHaavE2qtT4Dw0qVYgIpvONux3LIB88Dyy+GG4m9Q9bSib/QiqpVAe0tQseCaqVOoK1zZguiA
d7h4iPXLT2wXlbo7FbUa9l6q23RIbG1yTunk3j3cBYzo4K6zI7hVb/IvjyZhIRaylE2RFHKdPTJB
DmfpjwJW4zepjPRZ/wFiqvVFhutu7VYRgvCMp+P1VzhAgJfjJAEchcfMDD+/dNDDEb+f8rV0RW2o
nPBGEojqLGWE8wU6S1U1zua/UZgq19x6GBwyLCT6VpNd1t9hRpPYeuqsoz5kMvydGP/NcygRh7KB
EyaL+N7HNU2q6bvnDN2lLH6g6Q4/eh0DQXyX85Zl8GNzBBfa9sm4YdJMg3OoUoSQazNm1yR+3Kq1
HbzhS8AG6yXiF+Io0gH1MsUrRLpsH3VMLLi/dVXXR0FZcdIC9i5TPUpN/L/Mq7TfupADM1kEKPBm
VgSCPomHGvp3V4cdutPSspb6zjEAbZhmJfHLO98AauM6sTsontF/lrd6s059F9SLyhYIvWzuN+M6
j2mAKGSQqTA2ME5hQPzDBE+ASAyiuTS9JJm9auamjHheiCcObp8Owb121lX5nSWq7i5WgQKKC3MV
TxIVm8KL8/QzK/Qx2BljWq/wmve6a1OaUhzfYCERuUPLoD5ER/KNai3DGxkY8jL4z03lCvu2M8a1
tRWTgZhFj4lOdu2evadG3g4QAWahV8UguFjgd/v7GieF4pGo06AYEAtz2kBS9I0byLdRjGChxblL
785sEji0jjr2PvxQ9grPpWPhLtTPSeI5HNKSPgwJHHi/eM8yHl0Dza1zemsfq1fZY1/Uh1TqvdL5
qwT7DhA+62Xgpg9BAq5ixirDEHVwzC39G+XC4OOGdE7zY+Rryw2NtWj0XWDe2NG2RMiZgMI8TTNx
DU2rrRi1L0azkBNLyzVcopdnoIPsnBar1bYPLh56TzoJvaq7OMOVp5mTzRC1mBkl6UdKJxhCMOgJ
Hf0g0Lt6BTCQbq0CDZVw1RrkY7GcZKjIl2nZBxnW/oUI93BI++Q8FZgc0TX7n8y2dJswrVFATYyi
2n7MUfCMh/Eo6BGLtneQ0sVZ7PpKLpPR5k7rrUWNBThDoLoK7JukFfbhUz/PSxfU0CqK8g48IgNt
8WATGZCOTfQ8JF0PueDPNg498qCetSwkDtseTjwyGlp8FyWT2Yo+h+5x+d9b2SP42pCvPFCd50+h
2dvRewVimboFCB/oJ95APZzv97SljWGxKKI59w/I7KVHKgZW8ajQfJzyC0IuxLTTpI6zLgZk9m1s
qWtybKbPmQGTO4oLIYEWiLz+iQDWubeDtrXgAUs2n01hWC30h4qzJj9KtZ2sD2TNrvFH4OGAUr8B
Nfu6fSSUz3gDZSF8t3Vp9lBOtXACP9i8HddB3AXSlaj4cVSCkOrPh7lPdAM3lWcAZ45AUtwjicdT
0qrHe4Igu4J70IJhoLjvYe8wWztQI69zQdDq4h2HnXP2nhJha/flHzrjZ3ZJGz/n3fIvUVbfWJr8
zLOcaSUfaYY/6C2r67/drglNOubkqq3r0NH/7qBx1xcDNiOpRQwUf/9JYDxVlJtvl+Qbc935FRce
7GAgMMoOXcWiJz4oPeQalps4zY9dwqubcPfpZa/eQ0hoy6ZvsmL8fT6MPDPrArgEhT6AWYyd39YU
R/ue9KEyOGVGj4+3s4PnxtXea8YLa04hQS5BozLm0BBMsCaTkLP39zf1DoWHvHpQIjJaVgMckxD5
JcG4k1vdTHzrq/N3miQ48Q5wKWXOguuMGEuGnEJAYCg48jFGA7sueLl5pcPdj0WTkXK/jyJFvjL2
KmQpQOlu3v25cWf7uUoNzIcB3eLd3NvvK1pPnJ6eA0FRxjLblU9313P/Ttqb8urSBB5wtZ9gztR1
TuBluITQ8AWrNeaD+CgZvNa4bxWZXOQQjRKc3mo/HyYkohmqA+QG0fT5PGbhXQVYIEZW9U+YMtD7
9lTpF45Kp2lJ4A4R5NGPdtYQJPVto5zxGS3uxVyMccWQwTKF+vznS4CGmksYSiKLwKadDXST03cV
UZX6DyUqDU5njLf5pSGulyjNSRdJACvyC8FNlwoY4fLVtXdQ/IMBsekNyHjNSV9tTlPDD8NMMKkB
HvUWwp8R00e1d/xaUDkMxp/tv0uVDHYys6wfJuiF+gLzvS7cwT6AugKBF1+DQQlxpbqgND18ImSU
LpJ8nIrDoXYCDvvZAbXSm5oJRYYdswA+ITf6DjqCX1TH1p+FW/xSjRXADP+BidXnjnNJzcOY8yWl
7aPSwFW36KmJTTRS/1b6Zfa4TNUm9eeXtEeEK63rtIFbZU4vaGmnUAd9BqKroZxtv5fNhvP6f0Fq
eLOykmXQ4ikaiws/TscOpH+7XxyUeVnHLv68czS3rcYaPfV4noNYyg0Cd3UbaK7k3chra3RdMyvU
Osc4In2mT7cyPE502n0l/sWgyH7ruhEZrsiTOCbi7ODp3ejUV7PUFzm/43esQ2l8zk64jhRZSBDp
Hi+/qSCGYoYOrlVOJaRDmhtXInUowfEeFkbp/OdA7VMW6WVCUuhHzp4r/p2FBInjrEUksGy9Lr4O
SZexkfWayGWDkjtT6LqMblDVCnVt1HO04VApTmJ5T2TgQXeOYBkvMze9X3+75CU/ksISX8YwS400
KYJZyfioY1tf6TTphX+Yv+nFxpWkQ+lfVQlrNCMxxJc6SlzgQSqyC9NO6DgZirf42PPR+MDVON/3
ME+PBIMGRkYz8GQc0Bujt7en6g3ik8Bj+d63nbF/+oPIzhyfl5BdLQvxGYTKX8ZtoFma6D5KiBe6
6ju1cFGSN7FbSMOz5Qzsd4pQB7u20H4wHy3ghvG4yD9HbnM9OoptuF9xpJFfygkE0YJTcj2piPkr
ExI7OoScJFHLSzKaYweHfFK7ZJ1gR1o+QBzRK07zr5EZnoT6MczPMuoCf28laOC/Fdp7XJl1DlEJ
cVgozxniWNLKEwour6FbNeDhIiX82AFXDkEACnUPB6ymnWC6pxm36VEOL5A015qqXQdxIBKtc4GB
euZri9In6hRjPYYfnJuII8nUr3ia/9h3l+meI4eTAb040PQvOtR2IqEG5PQiwwUmZ0zFrccMncEh
XlgQsi6FUTSNNG4z7rieakvMqmAXfWNxSYnMJtPP9QsHsNR7+f+IZ8Vf0zeq4Z2j3YekgknyL1f8
jpaiK7OwjDVFl/RIL59gBNxf790qLzrw2i4IZvREdKSza36qTos1qN4doXDBFteYxglUQSTUEoSM
leP4zVdzO1+ka0CIYD5D0Um5l0y4CywMj4KALxhk/bjVsTaOcuEY6nhD2+9obZpH662AQEufkr3D
Awc7XvyVyfruVX5/b6pWxHWGPe+mgwQoaGxsyFCvgna4j6l136sGsX+cf32xuVgAVNmh/gKT5UZa
7jZbn8uyZ3LlUul15Y/b1Dujj4bLTL/OnnM90lp9qxS8Xaejuwb0X+1aT76Pgq4fdPPIFphF2V1J
p8kbFWfB/y0UHVG7IpQ/d+4JLN5bSxRqhLRQFoG9A3nKX1ttX0DoODS7ZYkgj/6VAR5itXBVNRs9
aZWEdTV/CggO9No7vBmqJVn4+owugY/0dLtiRxG9TJWf/4G3yi4i5tK8fvKAkt8pKMyvxCJCSKf9
Ivw+pTB5rteN05PDD5kEUaP9rgPCRlC1g3QuHfcoikAe8zl8ajFcAOHav/1EhXQRQqHypGqtHA6E
gYrl1BDJi7NUjwC/a413KZdI+4sdFZAbHwK2t67LeAbRg6rjQ93RrT4pvC8RPxnlN2Q35ZOPy6+G
cR3utbrFxPFUYyeAnPejRTyl4HA2j1RWBmz1K1FsAkYxydGVXkqE8YLR+7GFhMsm+nVCC4FFEqGX
OOuuiAMYko5sIdsW7S+1yTtMpSigDLAtEB9LRmVpyitPz2Xk03ntDDfrCKl/RtKz1V9LjEN89iPs
stRIpaaa29yOCNb4tgXXZ74kPdz9kqxQIM6gZp1OC/OnC+kQW9Jd7O5HP7D0DjCxwmhIBrA4h0Ey
4F+k73Fl5BKYP6TxECwM8Kz3o1Whzya5j280rBW505sH9QUy5frLm5M192XanDNyhL4koJ5ooILA
1llpb0mE2gqsWOzjunx1EfbDvJe5v4QDYhALWd3M3AP0kioF3cXv2IMqt8nrfeN36lnQHMuf/sKR
AYLowcXMgAX+erC8g660iOXJCUVkJxigMZ3ePqsnY6CoyWc3TY4MpgperwafjKsun19nXD4rT0aH
EGwpdQQJ5v2UylKRrCSqlzHRhEZnVsJgnQfEF42TrlM6wdZOPCxRZ6GTr7mtW2m/z5xoO7B9KRHc
o1goYJZfuPr/vHrx9Q+lI4rvWmtBVGjkcUqUAGsP+iEJjrQ8MOBQ0/D/+fdEKoJJGLsQYjOBNwXm
n8eeLnWv1R6HDf+Vo/GO38ZxUUbiaN0c3oyNR5L8dDGxU+QLlKtEz8uOS8rRXQhPosCvCL0N/YG/
XySz+0JIHFxWAB6eqb0kcrlpQN6F5JN+t6TgRQrM2uFInY4pr0xk5AwGgH1fMiX9v5quZ3rnE02F
j9VlSYJuPiSj4eHwg/sgoaxc5UPkIVtFm/s/+Zz58/aTpjY73ceUDXdWaMsUEyz8EbFW9namwtAL
15eIdBTUZ+HDU3HiPSD+DvJhJdg2cKwr/zAkwixdJmpjYeoMq/7H1tstaYkg7fiHiDalyEQ5qzuB
CkhvHu8FIFjDdJ2A1cXTOkx0m8WoQhauQctuNUEbxYOOO5K5GYYZPMT5F/CSv2/ycmAGJLSJZGjz
jkaO8OOE+K2x6rh+tC3Yf6+/p8hzmz6dRCImLbY7vBfMYbjHzLjhljlOT8WRIA8VLR39pWnDPxJY
P1IqnJVO6BG17gmGup2pZJUhf34LQNKhy+MElUIne5kBqVHQjErV4QrjMxZHfGsY/Fz9+IJB3dYL
u4wLiunEWPlGF1ZkMvMHPGOIUZXTghso7RutJCvKUGSqdRPqVIZkE5x/5AlQds1pfA6rq0mBocAV
e54Ao5kzv38s4GN45hmaElTgEFPbt5IJe0H0rgKHg9+AiSL3e8vNz0J78zUntHmhBrR5HSHw7E/E
9kEDWuX0GCVYMa0ItSClw5hIDcmGMahtExFGuVE54zLrBVdMNTJu6/2Ec/9OWSBHR4++aTv02+6M
LK+ySSkD4Pgji3jOXeBUOC+b2xdvFN5QkU9UMX45n/LiRC06VGG8OUaNgEye+nNDCOdTIZP/jMS6
FjsrtXvCG0smuqt2Xgf+JM6569wNlcQb3xKv9E+xR0dsbV3ourd5QZXnRcPVHKdTBmksXL0ik68u
6fzNmZR7X3gP2ST35nyRMkVxCsicRXqxww8SOVezOZ+YSB3kQLfPRt955ZoCr8VkAafhG3KzIjZh
E5m6nfuAZ0X+8yLo2/llFu1vj5znTgBOqmGIyYTB/8EhFcaBE++/Vr4z3swc150woOvMr5iqS1ps
5i+OWf4J6VNYICA+0S1XUYINJF94/T+be1rW6Lxd4fDfoIoHYh44bo5dmCJ1wcNvWv/sbu4eUj51
HJSpMed5uDKsWmG+JvjggNe6oItI1eYBlHhX5097jhakuV0LCgzpzS8oCCFauixkvteQ3fvdbpuy
zdDjzuDYvR640GtIWdMiRqfWEIIDXHANpyZfHLyu8CWKiXydrD+zOuhGRhTPCrqWa084o7vh53+K
+MEQZnSS4U0H6MyAjmoa22rIoWuBouSFWFnm6WxykgSIVHOfprOe7E56KgFkikAKBm3PHp5P1/6Y
OORo4zoythqxzfMy734moiksJ1lvDmmP7nCCaV1pju9yBws5fnTeVG+xnIo1hFcIFHf1mT26YUyN
7ZqDWc6UZU+KwC3xraiMAYizzvpt2trAde2Bdwptfl+qIYWAare01lVkq85ku6ojxfmeVxESu/SX
YchJ4f7T1OCKUnD5nF9ZBECBglHO88zAXZTYvwWrkL2VMXriFLabEbzchcPHKQRV9eE87o+TAzJO
LENy1FNDeP2SRkTAisd9sMGss/XuL+WhYSgvI/rPCLtagcyj0h2Z7u+URi7MbucuHk1Tco+zX0q+
9w0q0AzNTcjfQbdyvQL16/14swrvsKZ6vrlyArK6vTaaWP+BBbrZbwO3xwEbNiGAkiBvJkiKndlR
ZboKpBiPL1F/TbFusy1+vReDTfEb69mMCNeZZ6kZ4P3N3q7/czdXizivwEARHJBI5vzq7nKVWM8S
sm/xeVsPsfrvOQw6evnhvuzJ4vCaI4bHiz4ZL3dtQObky6WtMI+nyP4KohKJY6D7Q+QrcRx8UNHu
P70vA21v+OvH35aGnO3x4VXK4Dk7ehUOHtoAtIZItt4iIYofb2I8t+/jQ3XKQL2RxdARasFXHgO7
13myL0T7VCSBeuRCeGFKQMxLClSy6PhUSrTIysseXYyRaxapbeEB/FwTBDG03WftGQ8S7l8rplui
FUpfZ8gkSUEtXP+NQpcBQgCLBt9iFbWGuaNdxhshGDiH+KPpM4kY/cdJFL1EDRm33KHFt5v+tn02
nO+xCMIcCEc1nZhmm7irS1cCkGYDlmQ/cf4Tl1c9OfD6/IlEFZ/YaaDOt4lkSQHXUpgdtXvQYPDg
H5i0wUdu/Ueomm+eUwBWVFtGPgQo9scpEWyQRUpG3Q32XcJFiYz45ZY9V+58V6ojB7GfGqeRtKXu
w+IMAGrpJa2qhdvSeQhUDCRi0ApdOCUlXV8IEfZwDXDdtfIDyD8t32VI42ze+egFgQ0r5jaKxNTo
vNScvdPHx4N1cgR3Jz6zUL1LUAiEcczoedeIlSXkb9DRBB039ygShNoPhEJnOG1wr3/0PIegY0Or
XssWSI6tO8HBYc6QuSH8mrMUlCBRVBJ1p9+1wvQRuGCweT5tO2xMGE30/s8lCcjwXrL+CYRO1JAV
EKAiQq6hQ9Q0LWCr5uPLiNsEEf20EA7ine1feG9wq3D5wUlSQ6Bt+0FzkyK03CVCPOE7xezK28Ng
8HCSecIuJ0pvbgsx3uPdSutGW43aZssnglqJHG26WpXAcbbqk6Aiyc/HYR4Gp1mJwXzg0fyEIrds
X/EuU7jNp3qhVF3GkPbR4G8VUTUx5AnoTSmdvmVoIOJntLyNuiMR0Az7Aon4Trvr+Iu+k7rOfcaG
6AI6uaAHZ8IO6fAJIE1cujo7j4vhulrPwYmmsRkCNmbgEljmXkFjLxmcRtIzLBR7v+oLu8dnbF6f
RVLWt2NrtXFHyp5ldCT7/kA638caHFbvzJ/FclePUYz6uPBvTeXo5YPW1HchJ5aTuoFm52akFWFH
T4Xf9t46dfeDoBVZ0DVarA9fGtCmZ8FZjkCKvGD6U8wPg9HKVIPNqDxe37jXTXnN9yk6pNOuVlSA
jpAP4vBu/rOX12vCRf5vaLVj44smg6zpHxZBCEhw4orUo2kUL4xzG09KEs48VuhW65V972iQtf5A
QWmwKhpn7vmzLDzAgN6XSxyO3vW4VOP2XGtsbUAmNCQdvQMzMvBb7dpqjLkXlVI/frCmEAA5+7hO
IuKwmnQWhP3dwQJMCRH728kjOlIzNojQqQ7X64zYqK9NX3jCoI5H/p/r7RpacXdVgrcpchyn8jZK
GPMezGgO42x7UMbLx22jDoNqllx7DgxW68U2HNb79VGQER/Og66HsLh7JyJ2Rex4AcYiQXhzl8id
226G7x+akwSHm28OOWbd9xVjwXHFUVYPes46AdTGIHYiziS86UwN68NAvu13mEGaUrSaqcP3Tk3M
nr1Bb2sVs+lDxy5/MpjkRZVSDDsQqAyH7v3ZvE7B37sr+fGDkNFO1YP9WpHDXfmFsKaXhum8m6Dj
w7xxomhmjZNOFUmjnqiK9asfh1ZakB+TTojoLPN1X/SKP6KM1aFdcYuOfAOyxzB6tJRgDR1uAw7W
Y8uFzOb59cXPMlpBKcQroQUIARKDu+z0efrM19wTFZfM4vE174kyOqHDlQz22SPiYhcqA4ZYngmA
ZzIalIZ0uaV42jabtzoq2dGp265osFffat2Ct4d5bKIri1Dp0nlpDcStgTqIRpUvhrJC1xZ4C3ca
81b7+hKIyYj4uuWQ01/UJFNEyuqBUsJhEAXGhHt2UTgfgKQlin/YdNdUC2o1k16w5XsjDSHZyaDW
FFWdMCoLHhi1uAucZ4TujNxbMORQla5Yl+JRPwSyUL7khwim2cnlRt8ekcn41xVfSP51H7ztLizt
xrcdsIHV6SuHIC4UewYdZXabdXGHiy+ecbqvBlkybp4rRAAc/6+dYVIjw1jFA2IsxGP+CrFkp49n
L5wF6aG2p8+Z30msmxEuZn1HZA58hBvrYAERcsSHDpvKTD+k9wawUvk4xts8oV5zipauXbJi/O0h
fqCTt9raPVCk0sl0jqbQmclP6QefbkDLptQgheS7V6STzq16eQklMuyVGcjzITNFaoTacBXS4TKG
FrQYxFOoSZ36QcYTSXKpvYWs1T+ZPjsOcNiRLdlr4RQonNFCjvjzwCOup56UVc8U3S2iQtSy8qXg
SXv/DJcjACdcukpMC1i0K8q2iGsMV5RubEQuxplyi0SNJ7ZEYlRRW9ynTFeU6yJ2sOZbS6K6WPpV
m0uqeeQrDUeZL7oknYONo4yoKfYyzxoy5PoFKEHQip1oF+OsfnqSd16HGEhVKLptWjFptMzoMmdp
wRDh1kLG0H3m2aDKM5npX071+HDpmhSUhb1WhBcwSsa80Ef9HAioWnfD6/kqgqYocOtJ3H1Vpt6Y
fPS7A0GoQMROf57LkSuLPSZjvCaSj9hnpZ7iBTzpkwh6+sLczjRNwZlEGqLrMBoxIfQGSgkn0vbD
liJ/2h1vB0biRi+BRwVOU89ezEgCLt4GwFenUx9Vl+eRjkFvFGc+rR1fQrpt+EHy2VeoGe9SXeMB
j2QzZX6f6P560CQJQq/jeV66vfzaHXTCtufLypxerd86Jk/XgtsDAAyKgYaEP5usggp+c20YT949
rg0aPvyb+cQM1JHP2JeT13lBqqqdT1Omu9MEy4P1gbCrV0g1Lyf0V9+Q7zf2jBhM/fYEyk4YObzG
dt0iXGisxTiIvIMbAz+GdTWHBp5ZZ30LHhqVzreqVGcM3MAZ4HTXW15in7UKv1KCcbu3iToa0XDu
W41chxUuauhvVIS3i/VHlqLpTb4aET4PELwj1sqv8ElE6JKrs02KEm4crSvoi+7e1hv3sNLZp7C/
TeB8NYCnmZOtysMJC7FmhGWM0Ma73ue8yhQ/cQ7oebejSXOexj9btj9tyGcs2KzJWwTRdRNXM3lq
fni9MSrBvPJqYOzcfm6lrCkvoBAiSGLTSRWLjB6QNKDTMjgG6rqfIeR5RjoitI1hx9uFT/2xJ0t+
2QIM5hOUygxsmWlDinclRU36yqKupRzybHYKaYiYbsIgpNZ5yps7TQVc+LY66nEQ4LjloLSfc+IY
xdGZGA+2splCKpDXbkI7WfYBE9btjN2ZJ7Kk3rxH57vsxzGO6qVHhdNq+CsObNJR+816YKYBzlYD
bojGEHn4ODQxn4uVcC1eYmUanw0HHEzoMVBGLSgtJu+YubCFYmGXbUAVoq4c27MW+E6m+RjxOAnP
LmPqoOBhC/xy0azTeJl6v5f4fo2q2hE1PKdKVpapFt+UR0kyXttwiY6Z5zte3iZ1KzQNlGzFXLLg
royRUfIY1C87iPwUom7T9qtlqBiONeWkfz//eh28TfZb9cLPA3hqQmk9WyCIXIe90RJJjTnoYvo7
n7+uuz38MrN6AzomTgfwCGyGCpvxQAdYUj3/uRXp3wXoY1oNWAHbAiRbVRmqmC8v1IgxmmH3yQ8E
k/nL/Pp5b1K0mvTvr7xxfJY7R5p9ywph+uT6GJ2GM01PBB0ePvyp6RIKvR9KHQ7nDyy118frdc6A
rdSiocvHRX0fCvGIINBI1jqPT64i0xLzHjUulofNAvOrNeZ4TSyLky23Do+5K0jAaZw0Y+2r/onp
vGq99FyHtrTMUzVD6j7gCe2BvnWAB3Sxg5BsP37pxXb52IJmlNdpXgzXEm18akGiiD8RD1Bjuqed
v1n+hDWmqgxHylYFv8UePcCycYTMt4TEiOA201R6lURQmkaI7ZU/G0sYxEBHOqU61uB/M8fSZKz9
2OSB2lrORqsRSa3SxLpwU4wgHOfPbwu7v2jBp/T8Kkz8oWcvf+PhuU42LzH04fSF+IF+a3kCFjrT
/iFdW0Tk+iimioeykW+XmPtCs8ioQwd79TkUs2kN48J4rOUl0vsLGue9i0xc/uYlmsZtG/bJUL/A
KCVEjt65Lpafk/gmUDHML3Y9XuaDSx+g5sl4V4guSLjbsBfRrfwfEtOa7zpqmLyPoB+SwwNEVhG2
h2bzwVLwJSo2qtoNbL4H+yERWgZTaAcr43JvxdJuZKKovr7mE2xSEfmZ3j6F4Ia245WXS17lCHzH
3TIpmpmHql5EbnXt1URh8/gZW4V5rWt2+ikOWkEOy3PBV5CO5iAtdInYVTAOQTvzOHzLncT1gOWV
fqm9cRAyfDSs5k3HDFNeq83UIxGYjQiFupMs+Ognqpx7DEDh+LGNKVJZoMJXwyJfFUNbLZ6Mxo0M
k+KwKVrcGIH8jQqfCSpO1oqCsmcO/J73FdlCGYNt2nh9qgIsvjXqUVBYHPr+8BF0Q4N6Sc9YCuIY
hbAP9pbr8418Il/KL34ofbhxuALqhd/4OK43JUUsGiGd3LouViYsUSjHmFSRGof3U2QREDLe4yrG
4nA2glz79JpSqF01iBaaea01Ww4Iz3IagHWZ71aaYS8xIMMlfVd8nUDmuAxS/gY7u6UwGqBsBxHD
Uq7RrmVOIbahcYcwlI5/kjlsw/GWhqaFzpkA65TES4jREedh2aN/tbUOfRNeYyhpCTxdpL6SvoFO
Zk272XlUinKygrbJp5sb1i9mk48+8tIeeZ+uHSp257TKiKpCbAhG0McAyRBZ2pG9Y8cNw5W09Rzc
LjxIAekvo4aUAHzElnBfFXuNJluPTTXBWoK9MNITpe7jSoF+bMmPG1PEvpE76xDoWJz7Go4AxMJx
8yVt9ZGHTmptl/u3hU8pp92tswHUac96Ks79SkFfki1jso4QU4ecwAqfB2/6ZapdEh2eVpKFCtc4
GpXxugRpjMecmENafrAgOA6Kqt13JoQILv1ONIz7wzMiv7gMV1q3N0zsD9NFumw1CfsYj70jvHFK
VrzMP2Cbv1xOPzoPxW2le8hMja/e93T4mWRUqLOjW/P6lxcs6o0pfzATjM97EBhV2C7Khw33kn9Y
KUEg26GKcP4AHTlO0MP1ib/4UIrSLw8xDeq4ndMbGG/gacyaI1bysdG8ly+I9TOViiZ++ljOqbQY
QXXZW+lqLg51xsel+6EMeRoKfIB15NTig7y67lz4maFXzZDxFa9rY+uoJiCT4fQjzITA6asekTUF
E401y65/UhriNSdl00CZpHDBizBianAlAeAel+QyDTfueL/te2mPc90gpcRbzJakI53/PfvOme2w
tk2zdyiQdUGoYDVqkgrDJf5RtUsYX4+anEfEylonNxL49qhNF3ZTkF5/NL9sF7oAsvGF4PkNY3bu
59XU+mUxRh8RdBnWGhDckFFNGYG76ILEwnUNyeaP+NmrNfq+aPiUzwortqLkELJzvVNgGtZ64ysa
56A0t8qys/1tA8n2kLfrQfud14nwVJmlJK8OB2EMuFoNyc/WTpS1+YiBQCoI7FuQPKhHPZAuBFct
gVzuTn1tdMQclVry/C33GdOStbn10CLzkkLK/FvSgTdjqnmT8scTfc6P+cdsWJJ6iejslcR370Kt
C8SCybimsh2ay+JFQfa187iez8+fXaYU8xKC8nz5yCR2C9Ul21q3LVgRbYab1AoqCXb2zJ0CmuHK
GGwcP3JHvNAZT8hYTlYvQSNHnRhKh8MGsBLIyoILBpLUwQW3TRk7xuywWNJfY8oFy5bMKBopPr+X
R3IXn9uI8z2jxFYkS4NU1ZWam8Y3sgXVQj9RyCTc8dJkdXzO7FON02cWPtg/qxZtmkm62WJvICI3
/QYJGde/s0hJ/wpBOLRFkcPeAfpXFZ7nCgSjPAxDvAbPiZJ7wj/8pWGHsEoS+wdeMFNYcN2kQzF/
dM94Mph5O0ozliRYUmgN6wcFIBO+SoBoKriEVZFzeVJUiaDCS6m9FTVxS9M7fpTQCaWHWN/XfNf2
evLBIDJ95flUIxzK9cf766h+m6o57eUR+Fg9g2AnLudJurgeSPKpJxZZlrSisvKl/q+LbUdRtEG9
+H3F9/vf1l/lptPt6NsyjMqXBqRW9tap9H2PPzFYDlgmj/gIriTqPmqL6/rQRQtw2TP5KmwIAGWJ
6OfYJnHiMXI/Bbo5k1rF02SKxjOizLrUOUNN44Muj+faeMdWEpL8Ft2VzbfPHgtyVnqa4hmamud/
TZziMTb33tw7OPsWi//WSeNxLLIXs9EPbSXvEiHRrgM/CRJbdaT8HUlbC+1UnP5iCbMptkwijCBE
JXyJ0iflXnq7aL6HRlnuBA5k55KrUAhCC+XMRHBsCODIPsjJsHyRpa/5dkiYIdLsXr1e6NutSAv/
POgVXb47y1WHmOr7qNlyVtFTUfld6vbKexfVNg+81WNMpI+XiIFJTuP+B+MEZS5gmwOxgk16IPVD
fPYaMaUXml0q3EIlvk/tRYHkqcMPJbCxpcl1qBYOx+gOq8xLXrcBh1KHArQuy2e38EdI+rhSf33D
zACz3NY/Hg9Uq9RnHbluGPsR+mYt338CbzLoMu69SloZvJZDAYmWmSxm/JgFseDWZIJTPl0RBKHi
BVuWPMfz/jh1xTy1/ZFd7r75c87Yqqugl4qOZc3HxQC/EeS5COkP1qjHvKU8h0o+cHabq61ho8co
ZbfwxEMhu8j/TZoUSZSPl9p3HEa5qkWlcuUBlv0FyicJHmyWcM6MCLnBUDeq5T29eFjJCC0Ov7LG
m2AZm3BEnzF1sjjN6KxV6KplOb7WFSnZtkIe6vk6rxalTzewX9P9vnr25USd38M9aSenQ0lj5W5q
s+OOO8fB2n3QP3Im9d1mbjnxD/FGYQ1sczfbm465x3oUqR30u9SZcuvE7zaTkbIDns3GJ/lMjxMP
TgeJ47+mflEsex25uns7vfLe9FcvlS4dWplhn6oFis2ZGLmYn0Y821Vx0u7rPvG0D/L7vdYd3wYt
Wt3YwJHyeUckdM5GEOlVdOhqJBhwGwsCCjkZ3K1xHZ+v6x006HJl7IuHXdHDK+kHQYCrfVvuID/R
D88K0GfHwm8K7bgQ7MtVP73nlrq/79TnhXKdwuWBrX4ow6zhgNv/4M32hVAjRMLtCFt9Gl6GCBJq
VcX7nU4WAmfKKjNO60ot1QM073SUwDRowkuXNm5YP8zmzOeFxtE54dMyFsescFRuNmxuemz/KFzs
wA9kTavq3wrpo2WGEAFo29WIj3pNB7xIir3a/0gq09WeMp17UgPvmXwmyH4DT58AkbZIg3ugeWiT
9NBwBpFu97Plg3V1+YiATkGIq8TwO02qY1Vy8GWTAKk460LwAOUDw6GJpcapkyHO1LAHGQ49fWpe
mbrTY64+v2ZgzvzfGONs41cNaDdPprTZnOhPbBHh47ZuXEwKu6Rb1zItlz4HoiKDJfABMdh9JNid
dVgnLowiU0T3fzr3g2/uYMJtTG+qrGNY+2Xyuo8ZRMelzlY9ddRfh19doLNytW8ZIsLVm9uNH4bY
BVFnGUVB3+75rovc6fzmltb1k1bi0pIDnKXjrBd5mOYitFgsOg/W5oJuuUPW68FFIkI85rCseWPw
8lNehiQygYy5B+t7K3OakHBqQucN9sfAuWSSYufGugsW40HSzLxRW33I/ZpAaM3x3Kb3IYNgqP1t
gSr+XTZkO4uneR5Z5sgibV3OrcRBAO269R/TO2ETZcxG8dqL0e4DtXzKlDlAD84OjsfDaxpqnaAD
Tycg/Wj6ljDHLg+oCTbLpSF+z8nbzOUDGf6HQgiU9uowCYg9LLtqFPr0GTX3QmQZ0bF0f0DdTmRL
nvz0AQtLtq3Sn2tTYmuqFvzLgPALCBmxP4A3cvuE8zdmwZPxeL7Q2R0/qUSK18VI/RzUSoEJgmz4
SK+LV+394QubkcC1FXJP4VQs48RMzwC3PD2rOD1jQiHDFqe+ewCccdIGjATnNvu2EOEBkTRtnwpd
zy4RZMIKKA9OYQOp5F/SXqIt8qLn4xUY6BmMET0mLrsude/L6Xmvi901+j0BX8iRIAZw8raT74F9
D/GPIdbZXlECV4bm4AklfqsEHgH0tDxuEtJjVmyEGLzuj7LzzfVgwBiR7iey9jtrSIxIxcaGCA65
GczYayHgjwoGfDoLAW4Zq5ja7Br3i0bAhF5SkbqgNwGuajpw8pzNsq3Jdpya+n8O7d/jF1B0yiK+
zXIJms57RmQ7JxkIEac06Z9kpJV2Y/w81n3hs3gF58h8N4aJNZ6yCwhHRoWqs57OXiS+18XCESt9
hd00g7E13A6aW7iXvaQ+u92L13IiaDxqx0ZoghWi2/los0l7hHmjQRd7JWXief1i7AuK0ay+grQh
tATNVRagTbO7XeB7tPkepXUBimQwDK5G3gJFjNSbGuq/Lz1K0lIxy5sVjBGgKjDD52Xk+q5AD7Vs
ZejmObRzIOhCGT/ksdsUWQEFZL8W+W0iA/Ox5c2IUp5LjMZow57g2Na2fGbxkEoV1xJBi6NG6zpJ
8OiLZ0JQRjtvjRHy3XPouANLaliweJLp55+xy0rttdfRk2xpkp9dpC1fLTdWwr4iq7mUaKcTDYTy
lZfhZWbLhW45h+j0D/KhZrwuLBHiFnqG9QmxglNE44PldLg9GZkCdHDplRfGnBK2fhW41Uhqzr3/
uUkHeLjH5zBF/Wti/oOhuzD1Mh9EgHEJjZhHllShtW1kMdBaYLHKqY7CzFl+jcrSAGdiyY6rwY5E
kIWkk+5+CQnH2CHrMQ8JU3Uai7+qJxEDEdfUEHfwe1nPnMMRGG1CTKNf2gDxGg+W694YKuDwUaTN
ViU0Qm1HrgVOh7QMkv7eMnf3JzWJHIo9gECExHkAv0jvZud/98Yd1SOSOLyHkC1bmgvomnpC9A2V
ZJGJV6FKG+QSHxAcpsyE0K0MV1kswRbAitV7wvtxG+X9BizI4lWr/lAPdy67vWHaF+Bi1A2Zh2VO
nC9BJ0BLgmzMeEo/DF95oImD+m2gjGYgQ0zlF0Vm/S1hGzr+o7RZqvzE+ST/z7WyKQQ2PcHHN/+1
lay3wel/w3/DbJOXB7nBvn2yo9VATJQEgHzHfOJ6hUzXimtTFLc5x8883wzUkP51BFHspajk0sca
9mzhTTeotiA6dBA07wGsa65Bh6nWivGNg0nAzTZaLLklIhWIDHLcVFGz0pfuOcPamBYFersXdns4
iuXmiVWAkYypjduTlr+VqCIsX3rDZMchWKKspZ6yomJ7dh+c7HvsF6FZNASDYGUxymMMpWEZcARR
xhNJac869Kd7GhDPnim6bLdRDwo3VJvqeM2XCg99DnA9qhx7oPNgJ/OGdrgVXCNBfyYzlgu4EHZe
2Bvo7Z0aKgsvarkm8EmlLllCEt+cHhRFopWXHL5p9dsKNsYlusEhJb+Aw15nQJjVUdLVKSYs1mKQ
mY1VWXpJ4U+pkX/9tU5MpSrBR91l9NP/EQUznBVEEFMJjwTL9BNasCF+nDwdJlqnVtwabjInwnP/
h6p5NJg76dlqm4WcbMBlSpYt4vUyG+MJ3/FRG5KCGGYIIAFccTBUzIsAeE9uFbvQJq3p2bmeTkwM
T9wqwBD1pX3kWy1L7wQtRZFksDojco3Lyt2bu6tuJ1JBzEVQevDmEJBF5ScgtCmA2LOW3dNiAXoA
k5dUMrlsj2EE2s4C/aKj+zadqOuRpOG09Oz6JKAZ/Dwf3cay8ey6XaWYs+233HdUn1gaLJ0hGJPk
yExoF3PEXsUmRh0b1bypkJGVygdDySZ7dCBgF/oQ+9dFuvUOKNdtOHwxXCI7k1FCWTCqvjiQe1fW
16oSshEXHLBbHABwaakJyMRYguEXI7q4TPFoeKhAWDz43MAbqRWL3al/xjkIhgBPaRFisTPfh+YZ
qV5Dc7zAtU/4RltSv+w0tHyqJQp1Bj4Op4wxTS8F92/nd29iH7bIbsO9Am2YrFuiYjwu2hQg08Ny
YdsDSrBn1UHxlRkTTCSr8sU5U1FMOmuwPMbiOOUkXDhgbNeOmeG+Jj98CHcoYS+7tQeYTgPdtots
tdtHKhb1dGXMoOkYGi6IzLi9kbgWacjSVFwiu5xjyKMmQ8vG5K5CoBGHXzvjG0Jzas1N6Yjpe0PK
bPUXXYlpgQf5Q8sRberliGNW752CDhdrsXfXDUeB7UDbwA9Q6r90mqNXqFslv+72gMxvhBBUuw0b
EoDB1IM2OSKFFXEOQD188PUMvavzBCMD2RufuX2hBIdHLcyeRmT2UYO1c7HQrkSBTfnOvBSO1YZE
UyPfMNQg7p0QC6AQ6MJVzYUzXslS/4ts32TFaP4m09TLR8ji6VjTFy0Kd8PJt5Bi1yufae7pWFa9
H7yWtxWfZIJHfbkJ4awRfcX0/SNznTX6mt6rCoGIHPJXzK3lY5FPRLGI2ckrfr/Zlno1BtmzQBwQ
6CdQkEoA5n/kwJ8xj+ajIxEF7Smj4HYQN900xOAp8CTopn4yGfYCkLKeCRsI06FB+3aYTuuvyWuR
S3ltpOimJRR2BJTEDkkObRzLryd7qCDM5+92/UTMtA/Poiy12Thej2Rx2wCZL0Jh0fvdQgXBgxYD
+hne+a2rMsHT4sIsuby99GkoKBRpZ2czbGPnstV6x82if73tQaFUgAiwmv9DKxC+GM9gfQTAf7tr
Jwwq4+2mO00irTr5gpCRLeri2AzKDtQcEapJcftl7kWupRz+Dsoc4uVyA7sExVfs+p534+YzP2Ft
5A+53n7xw5MgjAXURkqNwAxt5WenGLvq1kJfbVKtMmcEOzZd9nFO68GqQSMV2QLtjWhUDMTmkpvu
2Yc04tnFFOTyaoiiJW4TrCItjDvk14jj0/74Qdm6vsWf92DZ7TgW75gdd4Cz2/OYEwwXHaZxZYPn
E0VV5UXks97mAF4MXkC+CBudVpBx5veEbl3Hhkv9RDZKHg2cMPiqp0ly26FvmcA6iFF95eO3r3ZX
cw9j5+Fm/nlMPTs5rfr03BsSky0FFVllPY9+lYD1Yfy0vkb4on2HEeZe3tgcSOXKxESTb/KCpwbD
cECL5jRNFnyWRUlTI9Wly+tCpEYxnLC9ve5I7u6v+jMMi2pA1qBsVsmayuaCCqxliEnRnmbPY2hf
+sA46LDl7UrvjwA5gT2/p+g21h1g8EF/ayl0rSLIZxNf5aEYi7gorU2uvLgjQd6i6PiTWY2Xbm1e
7eLgsNhHyv6tuh9YonQliRi0qckMVEwIHtfcajzuBNdlYSZAocIEtDzwg1ddA+H6WcwlBu8lWmUg
pwVquiwd9BzEGUQtPVzq1nyHpJBWJGku5g1AdBasnl2qx9Pc0BMy2zfYxQnfS4LUeJgX7yi8xNBS
jxzJrqLdTu7JFVl2jF4vpNg8oMXTiSkQMPg645vr6BHMNPecd/pWEbKmwvnn5vhq6Bc1onBv8FPg
Vpcq5ZeTEH0jqKxp1jfbNK0frpiQYmXoCDg4sLAEvIvC3iU3IPPMcPJ8WN4upeMEVva+NcLa+Otp
jH2V1HjcU4LhzG6B+99QWPU3fGBWbChQYUy86UNQB20r4owRXJzp7KlukUxYAHV3Kmds7riMvu4z
ZM5xtgcqi1t7vWOupcw0TsbGyrzHUZCew/PcBM3PltMz00hlg1u6WHJJUfvIdjXyjQtvz1Tqp2ka
M3T92njxD6BHz/8KnOLUO9SchfwcTbBcfUbQaExN+YJX/6XisAukL2iDBM9HjYwR8oKvIx0CLcNK
3G5p/44FUAHQynrtpKRQPVH205vdMY79w3IqSQXZr9T/2zDyUHy1kKNim4KPusWeqELNs1lrana1
oIbh6afGt2JoLAMAtyUFr9zXIUM4srsfia/HlvAZoKea9rnO6B06nPRsTB7MdNTe76GtOOY+VfS2
IHrw8F07QtHHh0bqN1gN7Daz1/D5BlG0rYmPM0bzXtuoztGzGiGPKSwex/djkyHhWx+3x3qsyOAW
q70sgUwlZnSmjZaJyw04A9CsFEKA2NduOTx/wCGpu+D+x65VVmySayBWGzl0dWQw+LGFsTXZA5nb
xiNP2Kha5OyEeTonZOwPQrT+mOX3XTG4TvsduHhc76jgXT+N+rsaYTaPiRfjW+bqJ4+5iNso0MVe
KPcNOrkJtQIJcUp7gLiyqG0O9xQLxyaY8c6vDGfeu1udHmZgTUDK37mlZlVA8RH0ZTWsjYGR/HZV
vZMEeZ33YU/v7LTKafymDOkVugcz7LK4VvcVxXbx0JyEIPti2x079s78GPDGBg/HcHYCpiwaphUT
0aO0PCzs3kpQBsC5ISLcULsLWBL25bfP/GMPFCknOQq4vrZQEi84YaoLLiA2s3Qu2FW6i18Qh0hm
1S8+F/raDtK48L+2wadPXxfzQlFmee5BRUmSpD2aqOalTnGIub0QHJ5hA+BapAWHh44r2vX/ENJY
FOb9Ga4ohjC/i+yokjz/ShSSpkhnDR2j/fWglCyyNiNbC0delF4vB0W16XTaw6c+vWAeXTgOEznR
+b7LUCQjrr13VsksjwARr58V8DRwuqV+ZMAC134nfvWAE5P3qmVOln+BhhhE2PncUsnJ4I2olg5F
RkLY8avRpyupmSl/37xRC6QP+k3gsqrt2v/EtMuyQK+9E1EBSkzbeNbGivfIOCAH9Jc3BXdqfAc6
WSJJTz/rue+lS2DWq6+lg8s06z3HaCaQXy2xEkMs+y9huWa1kAZ8UkWNXgAYMz6xZNNuE1wStPSp
WlGMusFQd+woY4ZL5WXCxZSmQN/6h4VS0D6tq7GtxH3lY1hIyHxzV00BKdX8ghlu3wmR453wxTQK
M9fWnw2xpHQT1yz9m4ASPaaxVOWKvPZaV8sq/UnGmfAYG+1G74ectXVACroq6glCGy7Ds4oq58MZ
y3iRg53a7jpaKpypOrFkfcG97I1vn/K55A/hvi0v6npGKLuqMWJ2wjQzh6Xm3KQrsXaKIduQm1ZF
pa4dkRYDfoDlHjoeTTX2Bp16+Yy6YLMwD8QBjTKZSvmS7hniCSKpcwFFarLTySvGvLlPwpG0pUIR
IE4fnd3QkfVq+fYRe0vcN/LlaNNLuruia6wcOYg8ojigCDnOGGttZ5/U/S3hvXukumOJ90uCtQn5
6cDOyp2HXKxbBTLGfZakAWE2kx2/c4Si8gGJu6KDEBpBiIQbs1c7Ohcd+3YjJTApVtmQdDxUrkLO
2V9TGyMLOn03F5YyC/qTZ2Ca6UHl3RrMQiN4aqjXxiwFFZhpS25omnOIhCmV0/lQNEgafjAmu3h2
vq9DW4y5lIvR5WGb6PxTFeQS5jyA2jSis+hDWBIsxABTNn9Mx0zzBZfBSum1Ds61vAdQlldmxPPP
xe6RdmBW5G/Wv9juZ6VeFXvG4ttT/0b649RRCklG7qc72AxoEA7s/ADCItVLSPKya+hNS+wSHcRB
I/Y3lgCDnw4OsEYBWCJehOIBhK7s4MTf9O04pp93pWTRv2KjXx7VdkD5wra/N+axMlfBL6ElxNx8
NInO6+hyhZhu0IAA9tXJZrYJqojgW2/8Glmm+bubti10m5l8ArdbVNmlSbdJSPU4GZnxl88buKD7
3MpTVWDZqrZM/TEQ+jXn6aljQKAX3oa92BisJKEakq4qkbr8g+yZAiEurN48BN6XGzzea49Gdho+
nXLwuAv8B0U2aaBM9WToH0l/WUOjvc/XGB3SD+jfoC4zg9KwdIccOEtWyxmH/b2CICjnRSfeFVe5
x+UobEpbkpU/YuV/nKE9KOUQrjvyNH1nOgHnVxwzE/PbRgQ4vmETh09OSP5bHdTPiPxShEf9XrBm
mkpAhNVBf2BWP6wvj/h6a4WYn0ecWE3Jmo8mFD8zHCGfosyhZTVsNlzdZqauxMmi0j2Z4CNrZlQO
wFv5WsiI5bLbE/e42BNgY/wrNAJpE18Q8cPGXQW95SBKnbHbE4bkTPCSaoBjVF0DTqWfsFjkDbJt
W6e0TROEEXv0YPe+j7qtkziV9Yb16Xs6IzXmTXjr512yEjI1WlCtQ5HT1K0TjbR2Y8Sy3lJOz6kn
2kFcn2R4tIO0yUqfk0SCNWrg9bX2BplILBvrrHjeBvdMDi4CCahQl2Oes/GQdZQpZ9z+UeD4JBdD
7bV+Im75RZMruR2wDyEXQDohyJXQPGBFHhYmJs+xGGXcMe+lEor6x2OLd7Uc+pReh8mjKZ+FBev+
j/Pav1yumVelSKT4KeCn83nnDyOXYjFXlRN2DhIu1dH6e9er7PV/mRGczibuLCPU+hqYXreNAqT4
pkqaBzrpTNvKXjpNa8xmAHaTjNGZt6tsWkiT9x4cD9F60+0hM+TBDTgs9cgghrDJ9Atv/RUXFm7Y
EcgxubTdZKOu+W84kO42yaQWOQxDBhsxGHrnihpkH8A0bYAzDIYNOAswg77rJro80atFVtuCf2Y+
NQuSez0SuKgPzQULZvLphOEvDoJA8Qu2ipkfc95jP41AZ/7zlP4QDcfUhE3YnXjR9x6nQZDW6FOB
jgt7uVU898MKgul5Fp1wCf1+FrQVhRz2gDQgBGQ/CpwxQX+T9iIzP7HySp21U9udMya/j0t8O8AT
jHhShZJGHdXuq0FeBv9Y0bi6PEX6rhRteyGHoHQ0vP3AmsvOf2MxeK7O5tu4uEdu/W3P52Y8LE7U
6nFat2BTlVEVNaMc4/jqs2pjC3m7EwIo6ZbGRivHOM+VYEvQGgkaNHiOdje8p9rilFMoxrO4bmXz
MyoCpbh6LaMQsVd56UawY/caJqL/z7WBNCELnEGcOgGnJ1dTl+dhmML1K6jXsflTNVqhgM2R+r8N
ohK9CCgMBOsD3YMri5v40bul71Mt4xqa3ttPDVwGROgcKbHQ2qZwksUp8J+HfCLyTJrraR8lfVlt
BdkAmnZ3MaaYgzBoPHRrA2O7xhPOgimHz9OVG95cTvaHXJyA6RPp+zfCLZstIJlm1Fx5L+bBZNZk
HBL6geYn70p4Oi2QYEUl8zR+YQXWkblqz8DwML+zaJPi9Znjbww946pdT+ZLrWXiDGT+yPLZEemr
0s/zWmXDGoqcDLi35e0yo0me8q4Hdzi2ItZ+PEodtu7MOfUtLUgvaOEPxOon3W9GUxutUJWRNCq0
bFJCAD7NuwMtB2ugJg4uY3zXS8hAUbrdrP4ItW2iU64SBE1cvMiVb2Pk7vIoxhevJOdIcna13RyS
537rT4rlZvm9gSOYZ6f4wW3lkIax7AOb6M8cSsd8kokXO9/w38gmd115CnCsFUadfrqtfAnkJXcQ
c58wf85zPMG4BbfO4ydVJwJxqmAPybDHlD6thRhB+m0xhpP7mV/zRyzP75txg9tYKJmH59ArmBUU
xVOIwFFD/tpn+HD9ifP8qCI4s+0/NbfecSPk4vSjiqq+sSyfrIwQgpxQqFmkTLECKmhOd74WTQJX
fi4itvJGOZMBn1HdZuIQH/AnJSYDMCSx7YuCSMJ2qaIh/mEM0h99BeDaN2DRwA4Ehcp7tvVV2m7W
4y6MNYmE3Mhgn1e/Yukd63thtGZI14MZjdZlaLwGM2UxVz2vL1TOx9eKZ7v1Hy+1gjXAVIx/DKc7
rSCuYNfLDHEKsoKBs0QarI3DbwgI0HFnVP5Bf6ZaPmpcheJPGU526OmrQh2gzyp52pLEpn6E1Zbp
q2fvfGVh6fpapo9RM81EUcD8NE6zswh+FKGRYbrY1ZyUIPU72oUTY6iiwnN6QsGkg2mgmlkCpZ/l
6gDtQvKfD6m6gfClDt2SO9GMzTDC12KLJ89g+XRU4+xAM/M/m9Cm68ygxYpwtFyarkSd1O28qZW/
xlChvnHG5sUHUcE2JH4bRcuxGftUx9Blv7b+UfZrMybFwDRZLH4pxd2/8u8UZabx3w8sglfLLRha
b33VuksZioPXswdPRjhi+jSqGEtzR/EGp/dfvduKyxrvmn24aisek2GjeGNNfIEwR+ITp77JsvSt
u0Iastwq+OI7a3M4K/dYEniFNbU169O/aGwEeQQRkn1f1ubN0XiDW5LuYIMSTUlz4HARZfX84foS
fMXcoGjkiXAmLSZEZO21w9s/LxzUwBXdDZ/l4QGnFlP1o7OlOmiuhLoEVFDu+ZT0jTJcYtG6HYwC
qBUdfEHGzR//aVEUuu1ksL0Hvj6q/6Fd/wcdRot203PeMKK9Byj+fCtSQu91DR3serEIRocq4vJw
fdWQZSj6qEcfDO9MgG8ZscISkBRLc87Gz8xc4GeAZ9gmqS+n4sPIQTtkF+Fn9jsRDPusuvO1ox0e
aDH4zz23C+3xgTiUC3Ikg+Bd02wxXIjoiKaCYjMGWZYo03UEh6V1f5X9jL2xyyBIu17OS/E32A5O
TMLViSEbqExeyvwW6EwbpbbxlEL6gnsHNyrcEV4ccR1EHEE+tfPDrBXEV86jmdRQT+bhK07hP60j
kqeVuSW2tHre6bwoUiW91h2R6f5+xXWAh0Elz+siIfZDkSr2VK42kdjnajqDrw1HWTDrjkOX/xlI
t7KXAnLZHvuapIrt1haDP/KHpYW0DeF4M6uMUKH6YDf3n+l8nkgDlnDj3Z52faSbD273MLwiKkLh
hD6MmY6qzba5Y6HDuHTgp5ZEnVkFMfxy4zuOFEkjmQYwb4UxLjziwj9BJXk6oauh8wNfHWN/t8II
q8cBNZSUrEf9ZkYoU2xFoSh22DzI0XCH9gJ7o3Eq3zpto8Lp50WpV4BiB87gJbOsqd5qnMPPD3l1
TmT1oCw2uPU3NIFUiq9MZLgrMIy3DYX8WIWaxkIBcG+hqrrI96mZS7yVZHzgCUnAXCgTZce+OkRY
PBb3AnTOqblDMY2iZHQLfoRx8JoMGd5qjOFIJ8W8McNVUe5Ek9dQyHqJI354Uh2qb5ShcW5MtJL9
pUQ2b0rM+DJ3tjAHOySC7iNPZVfoudegSOIOrPkuhXBvUqNUOtljlKCC3FCAhSr9iiF7XyOPlrhV
RDczV7IsDGVmReVbVPXJ9qbApPk2diTcscmi/dUEdd4jTvv9HdKGdWIh6kyY2Nizv72UXdyPoZC7
t7mpvcSFpRNwvrMp/xUcaV5UwjL1evIbMsOQjee/KjLMzX2CoYpf7I0DvWoSaIatIXqdMvMA7YIm
xIIafT6bM/pNIgzL72rxMEW6BWevErmIAIdTyHVCtKq++AB7tTXbwk7+WLgUtVOPPmMXz+DUAp3c
PpWoEE0RhvfyhYfrFsW60Rs5oZ0gAM2gmYAhDVQ4lhfznfnmvfbnzvdJT4UcQBpWiMZyUwRRjwpW
/LZl7PdHbl8Lv7hknFnWI7bQ+Cg4NE+6MLvdKIYXPZR+Oom42Zupkfo6R9iyi7XZg/RQyumxxVaY
OzpFhM7VycP5jZ2EdBDTMoFqgqpu5fly8MmINiAbw/cHtp7JAxQjOzKcb4U+4Y0H3CFABL5JhVsu
cs75A5A9JgJ2ngnD074kd3StdEJ5/5oaFIn4LVWhzpvwHJOB7gO0s0y7V4JbJRp0CAVAri6jOjIU
mPbjQPtP8A+h5PwuWtSo1rlsjZpP4UIifJL0aZbejGWupndS9RNk7wR0mEcASB+UeTfwOLJABQ8o
kfUf01psqZ+3IBRMcYfQALnSLMGOKw5HD/PmVThHRXjYTUifvwHI3yLGaHiag1aerH5tcab3dEwC
wKQGa4wyLEWpDi0y0AszUwcu4L5YwFvhSiHHgO/toXC89Pk6OPBX/h26LRh9PVVTHu/nOLPGJeHW
UIAgklqJxlbsG4Cx7Fjvlt5cc/w8Ou2mUGT0Ca+vwJ5A5NJsjbMi2Hru9b/IWYjLMeVgZbQRGD+u
33wYzEsUKeH8lVpR8YFwt5FSKl/URjYRdKobheNtRe4Tdt/wdwtSuJBObb7KH4QAJ6+36NZdT3s7
YXFm+9GexPy4fhhPaaVSoHj+Lv5sIU1+FVVWYshqnbvABU34AzzYmqwb0prbflYsDxAHFn+R5EZg
aQVGTFbOtb9V9rYVOhm9X0k6NizAberc1QipqXpLlhpZyT8quVdJe6fJwRjZkfxMl3/WVE6H5ahJ
JHWxjuuB4msj40ToOKh8J7oKV/+1Md5nq4jhkQm/o+WISANxSBc3JdcGqq19ldWbA+QIVxNqe5HX
czwpKncMeEHQZPfPs+S5HaItZUAwI1UftixwEZhJ71lhVSEbmVM68M+HGiaiTJFez/eJ+a7i9XXB
koQ8lRGrl0uoubctAK3gdvTuCRdD88bSrMuV9VLUMw5FKS3nQbR57M0Fy0N71/hmAoXPFPMQhVXa
wbc2OTSXQuYQB2wXZ6OzrJwzbo2tQkhn2xWyB0ZsJbDDw0+nXn2uiAdfPq2HmR8bduqvrhCEQ+HJ
QdWUT/3hXGV+F77GTL7BcnEeaFR9UQNcXnuHCtqzDKovTky8nSma6r0xh5FYw0aggA87p+1r83EI
QLUPlzSsnVQx0n3no3rcrygJtLWQo4d2+AHO5/1fdQZlMax0i+SB3ffhhno9MTVkZrGjVcoWjMtt
7Q6WVqA7mEHGSAkZs7zXYJlgtd5xhHDjlJdq66r1OW9DNIdZt4OdN7uBzWPobC5o58fZb/axTDbd
oVjiw86azUEiFMvE/b+9/SaW8o9v4SImckqOoeoTstf+9+V2gN8bkXDws/Hn7ZZpVdk/3le1Ktag
k3y/bTTMatt5ASfvOusG6Ii4FoTTI7xZVJgYtcKc4XS/Mi8wDHxz7mEMFW08KOf04zuOp479PogQ
L9xs4E2IPOIu/VTa1FjjFneMIpbQiY9Wp1YCQFnZLIW1oXCNUerXV2w4JTY5rWYjUhFU4T38+alq
uYxdxQ9ZbYAqrQfvU8SRx+m5UNhxGlD/+UgcWPNn7PCzsROBIN1AXPHWiA3iyWSWlU7+2mFH4YL3
IwAzNdyueHwKwT0fLNP0b8/oe9f7K7HUqG5vJtnWAZb5+GHrWezQP+2ls9/sH+oVqzF1PCf2AHjZ
rw6/z44jfhbRngiO+/3o+sFZICCDK7tsd1j/FouFKht8IrbRG8A43pwj38YjDQUGtAsoyG3hfHK5
bTcpseZ8R0Hpk0BR9fODs/LuHffOmACrbOqN9E8z5BaKpgLuq6Pm0eZV3Ws1R8MEWyMNRpSi2Ubq
Xn0G2cxxyFHSG7dkujNliNg327RbCPt3rxbaUoSTDZSN/7zcx+AWEBK72Y0vhQai4stOScj2NwBs
gFkINevbcxtpFFU3bJAtbcCGjcVEmt+6KI3WbotHrZM/mUHXyuJ4BMZsqLxTGTA/F/VlI+PpD20l
j3+ySWpWZDn1IqrJBUkcmkZKruj2UsCaVp9Mjx8VUSaW37FmlA8O9KE9iZlJHbZlVJYn34WGJ6yN
UCv8jdHnKad99DzNRbcp5cX9mgKSDvq3S2KT4jTxTppeTpBEdrzv+CmtyWYXmcCVq+81hAFS6+vH
4k+1x/32sWqv3XbDYFUn2RMLHxc3udBKDWnKXHmOgapfLVXmkgzUCfEvMtaXdAxo1hn4O6e2EABh
ZEBOZEgGXNsIU2xZJhlr1LXMXDYO+JB9PR5ubwAq+BZmfafKvrwGOvStoaMWR7defY8x2IzJxeQS
YvP2AjpyrMbqVIJM/w+tb+J7hEsI+vIiGjscEQBBIdCygjcL8rmsg21ZNdga1f+1ERmWIB6ML4Lv
8b9oSjjsvyt/SuHnbji3KHkt9d5KFbAlVWRRqqZTwG1jVO4NDx4lbHjupY/YV+qlcKA4S/4sES1/
D5rOpXOywPC+F6Hq4RM0o9YIrlnDeFH/td+MQ5MmCGxyjBqT5ivTnbwnVn+lSxWv8ShrEaa+MDVH
vY2gESj7pfYh3pHSdCw51W+xxCRH9pm3T1ZbqfmNRuu9bioMppJZDl1d+mf91dP18Dqjt2aY5ghZ
8xvFGyr3xaqrGMypKGK2g+2lUNOf5xlp5ZI092fdYZb29u+/fO1D8TnhV6teTJon3RdJdFbbUKR0
YyOvwIi6FOOklMnZkXkPpiC5BrTm0HHF2DJWPSvb68Bkc9tX+sMtygh0R6gD1V24GSRRNEkgtAny
I1yMCw9xGi0ps5GMh++vV1cFjFSOdhR0f4IyQYeE0hiSKDBHBIC8pTM9P24xX1lMbNqRfFpurN2C
sfcqjLpf4MkUJxFAbjQSmdpafiZ0nUVvo1xIuZl6I7Hf62ZIgJ4buaad9aNd/lr3lhL7VeSDJpT5
4hliTco/nfBA9nxfevLwOu7s8DjdESoGQkl9/T3jhmDCgkwqaOzBeCSBiInpDM2eVDCXhl1oDact
rWdCqgEo7a6qGv1Dqx2EwnbiCOK2E+sVnRHul3FzUr6BoLlO99AwNlBFybIPpdSlMOEnFs9j/m++
emR3GpaRRibPkZUkkOpHxJta4s3m3a4UxWcbGbYAy+NsSnRJjThGXserxqEdThqz2F+KvFb/Po5Z
2qa6whfd7izvQatjc2Gv8Oj3L7lD9jIU48ePtaJ/IYrx8dfCxo/e4wEuuN3Mop2+aw7oqDOsE2G/
mv80qfELUe5jL1TzwVCLickjD+S7Cp3Dt4Y+pqGC72vZCsAWqOU1PH/cGmd3EEySX+TWyYelp2a4
/gTxU/2kwK2SKy8CvSUNZ7/WqqIVjZENpyu8CA2gu2XAvaR3Gpe6jvQWwpHdQlIUoqH8VdfPtg0W
4F3k5gG+potwAjwRFx2ueOZlZ5gLzcX8CDrHG0kfhNLsu3aOFqygjzxtnJLTY+NgeWxsIxczDuvm
k7/Cge5LhkX2WMO1WgMOaBx2zeF+o24xZCAfxdtX+l8NwXvhy5OKbbUKcK7LnDGoFJTUZvVbroQv
YyxiMlIk8YlpUhB/mHBGcWAvplaNRdJz1U5SrZm+JLLlehn6mlFA3IkI9PG+pAaF+2UJiDhl7PPd
u7exZwdKAZHT6Gps2g1RMiqYkOpqAvg6VLHh0fsv3mtBEbqN7awg0G51WjoM6d+XugTIHz/eUdpK
jSnShKrLGc5ybzcL2xuo2Ibf72t/c9a+NGGDPnGPY5NWDxf8n2vKlle5htmV2McOGqSf+C6z3jWE
6vUvCv6If/iEMJFaEt7TzmdwwWNI/pnRCpdBQmm96Xh5Pz2O+icrPBackOzasC709Cq8nKcSAkrh
cUec4wwWPBuOnidRomDqoRnC0Isb/vJpyB25f92UC6dcPxheBABa3MreSUr/72KOI/1Oc7bY8akk
l0krKN2fZ+Mg/C/+DGVXCaaxcBaQ1WMgTGPGByd+a8vrvPSS9Ca7BWvhuMt0sq2E/rGUSUXxD/MY
mQUf9S/8AXdpsApZ/ADthiMROmBgGjZjCo6//RjOwZXyrV7FvLkadxAcFKPfdHpA5sx1knMp7EQ1
tnr7iUZwAh2uduukOrNxxwZy+M761YPY4G9pLtht8yr9rNdjo26tt1+ES0k400TSZ0C7xvRoPnCd
L8LZX/+iyhDVt5HLY54+/wlPNHaC7HnkC4Yv+mTos4R37vfMLhjMtN/PEtw8BUx9hRCiW4HCARti
wP42BaJmgy2wrSM7e8drpOvYYlSzbBeR+TBa/qpXRCwXEPaJocP2h8q2wB2+jlPxHjbAj8jJZ+Pz
wrthYunItVABe4LtxzhJs46MKyz8/bOC8LCUajBNWq1vC67+zdm1TszC2X541+UyrF0EXl/HNfBL
QfLUw71ogYiHZ8XJozZugzpYXelVx3zYcoFkDHFvBFaXVSdrj1sVgJdsuypZOuvOYBNHi6RvJ9KP
LGh2qfRCRZYe9DkfW6uDqUv2OCcAFguanDcBoW9BjVOniRowHcFjAAEVZ4oK1o8aPOU7miD9MHP7
IvKi+JqGz/RO3J03GC3tYJ9j+tHxpgSDkVvkcwlREUohUzcEUAENL9pIxh78R6qEt0xqIShi2v2U
1VAhGu2nIGABsSxDL8WdAWAioZrR0ewAz1Tjr4eO9VoWokodWV7+ZnJET4ApGYV8AX4ZtkRYsQO8
+Fhuj1WHuKRbR3XX3l67u9lRF4zWsrf07X6/uu/G+2URa3rgkv9S8eLvrJ58yjqxEbSHXeB2ATfg
ZudG5n+PCx/duJTx7yhPJhdNw52dy4NbLqkPAorZKgkKzPq0riAB7FogWo6GX63TvelcNkEkPw25
iDyZxt/MlH6af5+UkxjXqZob6cH0COKVXgjdcKshvgFytccKiGpeLz26nC4Daew2egyXU9joggIt
ggRIkt07B7BmMZwwOD+ziPGv78rm+D9uSXayjdor7OyHCF6W1gpfLVy1ua7Zu5Tiza8XS7rqe460
Sz4ySIb9Kiiz1LoA0B8t3MpBp1Vj07b3a5a12fXjiE83/kQg5GvolRzxyjrp1xapvooPbB806NRQ
h41+gzP91QnRYL5I5JN3Xu27RyJZ9N3ttyRyEpscInqUVkaMTh9341Z/HMF6vSF2wEaqeYEnHxXT
Anj9P+8FM92XfmMMYhcUcNJJT7dPK/zd5FImYnn4orKm7dJ7gaN6p1jehLBHHVxNk00S7IyXUDIM
ru+eJA2Ak5uQUPc+61ErnuxqU+EaDP6s1JWAttcccqBZsD+lLTbuDYj/DwaJOv7vdF2UiOASmrrH
BoNY8voSg63MAwtoPdFniq6e2GoQN0cmV6+mYv4zMV1599IBilABV1UpQYcFII83g+rcvzw/0ebS
qlC6CFMHNBSWtiTWlXJt12rbyXf6u+5posO0ynKXaUBbv0n1ERNL/ZdNReCe8FETEVHzJeSJJJXd
YUF2rtdTutG9bD7rbxXSkXw/wca+VELu4SRfYDVYf/Cx/kqzOjH/4Dw5c0woyCJ3w5bZd4fglenx
7V5gzRVSOilCmVR0ahGJOaIh0tizuBU+kNtfR+gjSR7uX4e5OTtg8KGWh29hPKgRHni4d4VnQl8+
CMfnfM2icBGfciH/XbEvJFlyIHRqsNIUuAAKq98cBMHxhKktJrY/3KjF25QCf1BcgshdzF/SwBz3
zF0jbvZLqqaWdONCAvawXnA/x/bwCu0nvF5flZIjrKa4w2iJ2jLe601+C+PYVzmOdLpa+UuKmVqF
HCBfAQTrlrS5Ree7QoCZqXKig0eVI//5gKm0RmFusCzWIeDiMiUVU3SnRbRTpl/odQYGjN1w/Brl
EEcEbxmdLSo2hmmOv0EJCJsvgA62yAVs0wb273dY12kDTLcnLt+UdNrXjrlwm0P9eZQxz1Cb3PZn
u1ORtBUjQ1UTWnHfOyXB23bvUVzXx5LlOl2bTXAaOX5ltPtbVhkUzxmFEwlqk6bAhPpzGtj67CUU
AqzGA6ot3bseUS8xfXRYJ7yvL+hxp7m4qdudp59Zp8LxTGkjkPQprog6Sh7tZlaIjZkdhPVQniHi
02+CJ1MQxeYOffy795fVjyapHUkLkcCXm+MaVMj6pPSRIVGjEVngENx3YZFuJtF8JUbpQdGLYQ8S
MskqCO80gQpVpf3zMnfq3jsp06PVphRibOakHhLj96IJfepStwZV9jFiets3CJP5eNA6793zfGQj
qpfUgJbPrcHairAXeisXd83tFB1lckNrvWW/f7Ocd6qeaQYXLmRhEvUKirGu1TFZGiSZgroKjcBQ
gmHZwGfagxQIBVOZjFaWDAZyA5yWXLHD5KMwWbwinEISeprqRmEgApYriP8hU9N66y6XJ6MWh06C
NajX3bUhFb/H7TvZPhr55MpU1/CkiYcU1Wj7l78gaJqYe61LRc2CUvlZUowt/Xj/S/Oa0AhLQdXF
4sAbp/CYOKG4rSAv5sVvR7hyso8YHhiWJYS0oLFquwUgt6/E6jUtEdWLOlVyiP9fRyZopv4OCg97
r+jQkhc8zL/KzMaSihcGqtVFH5uR7kN916AbBso3LlOwP2mJV08oDRlqgKbQqr/MyiDuCNAjQAU5
3+WeZDPGV/6A9wesh78z+gtq6rjmSZaRPZZvb2WfU4X75LskzgcFce3rtcGsD6FxDdHCyDPtCIzG
69YDNWrOe/LxfEjLC0tAYF/Yits/RjjEafdwIxOPDxOjIyqnhS/nXOUrtI5aO93x/6qlr3e1Tijb
w0EgZkJWRG/ocQYZ5iv4k1/zOZkCElDkXshZB4yFKYfnactfFpxs2m8x77+S886JP3RFfiQ72Pp1
Ayvy7o5DTiPRVtz16Ki8jGew1a3zrvLr6h7f1VEesx6wo84rdahc29N797I03zpl7sxv/FQLp5ls
33LtiSv8QV7Do5kDfe2nfY46iMUHoJQfVE0uVY2x2PWEFlz74TgGs9FREDkZ24JZTYMOyFhARsXw
HPV5ZXE1CNKZXeFgnOiGRokfteAWiKWeAN+lV52hM9nJ8VQy2XTxa71e+kR0TqhSAU4ebu7k8Crj
AfnIORvPtjlKiqiJ4qECpoPe02YdFhehxterQ29HsOEfsfPZBSBKm+FuwnnQ5e02gqQqgAzTtYWI
p468TBXI5n5nvIo9PQd93pw3GW+DR9A+3sfzPqXqDTa1nNMWy/qARW73JT0keq3qwuX728VQiwJA
JWZar4NdoCUzNtkRB1Hc9/kcSLOOGMoBw3cKrmau5zVJeDAfJGi+ZClsbWwlR41KRQ5MTQlGStUf
QQ1lgSZcby4yKVhB1K+2Q+Zg2/2+67/XMpGUbKfsY53D7al1K7Pwdk57cBI3g+PMOSUKorOEf9S0
aTp/4Ki32BfxFwv4dAd9fT7zmp3EjXhsIPrE+quQzchaI4CFH8orVZs2PWppZ+Uqm1RlHCqnR5Wj
uDGtOJ3mWy7HiBxi66N90J4bNOBfbtMUe9IhUciI5RvCcTpkTUxV5mX0E3qpU/8bc4uzwOSnx5Te
aVNapnl7p+PHfbHX4EFQ8MLmM/Czhsfy8MGPHJJ3jgAlnMS9dNHJ73VtOdOgnMY6q4W/mhSWdEPY
n1el2rlsvIq93Xdm15qcjiR+w2V3UimEjphC1JvueGgbrXUDCI1YGjAUHYVRhgHONtXGRGds3N+X
8lm/VGE3dxHBMEM7yfU/2Adh11ShsORHZUI+b9QAPe/loF6m2WIvy6b01a1jAXFQ+QJpQyJzhQCi
C8uFsD9OlerC9rX+lsx/40msLvZO/qBzduscS/66/JALBjtKgvBEtkQ3HTbinJU0M6rGSLaM37Mm
r4Y/s2YUhUVIM2W2r+3FffptCfGIQj8KgX/VkBiLLvLbsRlX83DeGl9Fbg5XUKEt5V1JHeYGlsgq
hvUzj+lPnJq96e1seRwNBK6+wB1qGCYzAodppj1j05Ypcy/fjySs72lZOR8GuLeb9hPEgnk+RgfC
NirN1/KQulN0nUXZN4LsRiI8p4PDFoBmVdENGmxa8HoaptbGAEAJ///CkSU2UYpACKRb64931eIT
QovovEQXrw+xqFfWHSffXJrZpcOfMMNxfctQ0am1yDnE62oKxJ/bfN4b+5LjzLgm++BCCOqv51Jp
ZlKiZANqgBDGHXj7bRXgb0hozu2E04V31lMHAAKhAc25P1YLyAPME5iKgxDdhuemqLhVuQTgiok/
1Nwl22IsftwxZLW7ONL2DCBdr/fbiAgjqNuKgBxcMdpsZtdwvdfpkGxlStHjZodUMqgCX3PXoXzC
FP5VO8WYl62He83z+QqoQEEZcJGcTxZ4wZ/tzH7vVpZnRHIdlSE6mbbOXi//onwmyCFhHeDMVFsl
mVkXyfaZHI74KCOMjJpoBbYyecWmhrQAqPB1aTH7l6BZaBGHvrjHtu11criq4EengNRMSGMlTJTG
kMCTmLQSVPcgKcn6SExnbtDGNScQ0uK8zstOt+59c4EkMlLurQnF5Gbz9ovIgKIGaEUyGZghMY3D
ay3CXfWw/5w2Es5cuLgLYV2pD0qrdW6mA+6ql814u99FdCDqI9kpfFxtg9hPgouk1n3ssERSj5i2
6EVx6x9e2LTEzylZ3UlJlLtxWmENkgtWeYvdjcPDGafnOqLcrfg4WfEEd9XkAxSYQVw/GTWHFjKi
n6bVdkzV2Cwye9RorF5VnYkgggrtnXO7sVibGDYF1SKrn3Qcra0Rbn39vtMaxEWsu6anRmNLGg1z
ACYXZwEns0gNj3sINWRRfFee7yBbBXBC0aVu8h1EjhWL19hLUikao97DBGVgqG44Qj+UuIS5ZOkw
eInT1FsWhzKKYG2tN+cWgsIEtQ4fh0Q1PMd1hh8jrA5IGbMKJLiwC3oAJmZfk/MaxuEzR1YWINu1
tGXjZOJSVuWb+9XwomgEbyKKRp+6VZ4crNqb+UTxCq25jczvUPCC9u1o5IEB6h9WDpxVLMerZQND
XfHXRaIjfua/FN5pG9ONkYzvMZucSkMxpF+hQYumrKqHL5WEAjQYkHWSy/2gptLV6e4crZT+94uQ
TaroxSTApqob1JheKBhYHTGw5yVAFkvQNAqiSJyIlZKhJqkDBNhbEVY5kagSoTkqdRJHr5WMLm+u
mhN9LN6df14oCl4rw6TaXRUT8HMp/ciZKnohmrUdtKdSCqhg7JEF5EwHybQAPDjxwCmdZAyjPoaA
Fr0jjUIYPYBsP4GyZRU+ULQu5tNXxlEZ78m/4sbNgV0FNntLuB7PgH9u3KLg98buJ8bl5EKlaW8v
aOTzopjKaZF0zIyjiDGrCmOHLnj2rvvCr+PIzxM/GezVXl2TvUbkYEwzvcQy+713sMPyjMRlDjjk
KZPe5Lyb/kqqjlgJ/PPMXdYq7b0UemCL+ZbmRcjOsI1RM8k5ovvJqt2Fz1pp1K2ZubCSvNnXxtR7
wFf3rDkpVCabOyim3ucTurRegMFeTBX+yeMsUGAADvF9VwVEccwfZ/My5uiZarZPB8jyHg8evxb/
I96Jnmxw4qr7+vd/V3ERmYQA+l2TBNupJltsCq9TcYS7DSQ8Yk6Pi9HOETusRrL6NAchCwCuILkz
7GqugF230db3hMiTFHJaY4QR0J5P2pv3y2uebH8YHcVu6TI+Q8RB1oSam+lsSedEGqqYW8WXCoSJ
xeWMDooCI1QVx5Rr9Bma6dDoSY7rKtLmUrhNgN5dV7+ipvaLL43RURxM0xkzHciI45SxfZ8C7MpP
Cx7EVIk2VO/ZQ3bhVAutOwVz2Lje7pbcTrxK+khAmrjd16wY8n+1DOS9JHHbWJuWcl4147Mo6oq/
00Tauk1CSsxUICyWyC1eX1GVvbf94iXXvUe0G0+3aoDiOaGtj6gAeSvWQxgsCAjrl4oCcIKA84BW
BSHgGBs1iNndt/EKdM3YTa71ztpM3H12Ej0pxGB3eovyAwMd5pLmqMlPeiiG2+Ne56qktGEXoqH3
SAfJdSEbLWCfTmnmHp3nYZFSD/zGfKhMHVlM6s9IAju3WAFYqm8qYbmhTHa2QrLo3K1aoP/mKQOq
nvZsmCeSnvNzUzxjglabMsCemsdM7CZIqW4g5v2nXlhnWtbwGAHcy6Vx3hoQhTeLCAdGc560vQhQ
OPba/pTwDEWQsX10OvWPscAbKE6ZpbQ1M7FZewVjYpbmc17AOmzq83JNLdtTUHFfiqICncA6b7gZ
cg39U5D8HQUv4ZwOtG9sEtHKaV7FzJUKwgaEu3N69TtZ76XAH5iX3pN7zxRXkm9Nud7HTC6rcobN
9CFr+vJ1nXCujS7mAKIFPiqwwwCfYYBoDtUJGr9TAA7ZYQT/NAQ4hPA8Fd2fi/YZOi92RxS9a/DK
n221Yqu/F0GedvxaISO6j0FqdFCCEzKr0twpPmkC5zSZx6DofivOaarOW35aOpvo5VsCXjCEf2XJ
bgaCy3FSTzhsf/LDjfAbnvyqZm2qs2ad5p/FVlbLTZRLWhGnSXQzuauqCwt6GeVHAatGCVG0KizC
qQoxQLr/Ktmv5G1XdE+rWNsZSPKnFYBkhizg613VhUC4KB/RX5qSIjsoXmI3H4cxw8oYmoYNEAnY
ttTajmHgfuozLv1jIhqgqlfh5sFbMydHKX23Wz7uXMuB4sS+8AdoueNMIT0+wIBfsl1mYYlSojkl
ARMXYvnWh9uB6pIQIQeiRS3L+LBWppH99wRxbtNUOHkU5TfN1WEIZcglZvWnPk1fEtaeGzLr+b1m
sxf625cWdRdmYoAws7Ywf+ouE7sF+9IRW3016PKBFcD5BrZ5+TCToFhaARYfhvH4gbaOXT1zN512
kz6gsAlO1/4zzqTNBlcfXRz0pzMsonwv05i0Zp5XSP17dY9ckDIdTH2+/ixTSF1yGDfrbCmAUJa2
XbJfuf80bTHhs8Kjlne9ISkz8FUHFSUGs6NWndCvL8sis0GsORg+Ldz+spELKuAuYSqIk0hlTKDo
xstw1t+LW8i223Lh/RRPPFV9qfxYWfxnAu/rZNUHsUFHkLll1oEqoRL7dzhvlwzG2wOo8rSp5hmu
mNjX/3bOsplFMrWhf97WwSStp7Hc8zfR6Md/2rVgZufnny3m6EY92EiFnPr6pm9wIuEI9JNFm+Nh
BWiyWmiYKrVszIcKmwYVoktYMjgkXJXQ5mkyCylWNg3Q8wN+MBhsFZ14078i4895bxJQ6sOO8hN7
iZTwLZPIFJBlNyv7JoEFjv6RExK+R+BXKPQxeipsVVcRT35kk9urrs9Qn17+VLAbaw+JLf14csUD
8qVxiugsL1TeXRaMYfecEL5fsNM309PVyjHA1fXwG/sLQ0DBwzMpy3dVGUvV8TucLLBEkj2icol1
B0yatB+Ltva9dsLB+aLLi1BE8xHO1cssTPZMmI7EvmF+hNpBWQ+46qr6cauUq3rzvk2Ux3wgNI2q
JfSk/kMrFnFRxYUVPf6KCDc39ga6DaJjlnF2ocRyeUxRcikgv5+QpWiNh5cfV8CBkq21qTj0d7qb
+FU6R44sgBVHFvvOHRP5vy8qsUCnPCMXhTLnbN1lk7e2U1V6gS7QyS/Cs8liS17FiY+5EjMzlvpa
u0aD/5pHJb2Nq+S9aDcYmHFQL/HtBBT97Gt8RAq1/rMlVmr8BCPARyHrGNIYnCLJf3GNqHdb8KCH
g4PSt1tg/3CC0NKfFEwyrXgFKQCAPcVViMT8UF487VRshIUMC1yGk42cQ2ziXJkHaIW/SdUmgadN
iJcACNyFLwK88dVbSupX5UkNWHNoru9DRa6Y8RTPR/e/+aCs5tzqzrOAg8L1es3NaLYpIIT8bpR3
Vfxs1t4H5R3IO3W9Z+sQZRvY4hc07XbdoEtiIh2k3zwgre7OeBEuRKvW0jtSz3utOeB8HhP/ha2l
7SV8j+hMkB63g0QuK/4xwStichoz8xNoc/DXGVUYlpgZkxPcLkKxfxCjQtt4lWKxh4eqjp2gIyNR
6NGxURXLbErHfHkSJWmN0FTHvGk1+6N4212H1YUpPhtD1aHf5OJQuk6Bjv0i5ve6XROqKWs0i6+B
C3F+L9iC9FHgQkNfHb5e9may8xTgObha4cr9MakmVtfcV3NWSJgfMW3y7quvsPNBI68VW/kBZHME
ouBe9uW+3l0P4p76jEdHkiVn9XdCAGQP1JnqcwQL4FZWkqJXM61t+7uTddoT3pMXtnUpP4sswlsN
DxGNFX/p3lIA2pJXymE7gEXoAc6X+F3u15RtgvPChX6pQC0lymF8iha/c7N361ywah1N+fHIhjFk
uQ538t/mGbj+t5nzgf5JkDMI3si305bJ0H5teOMhcoPM0NGVqmcmhFrOtk4pdGgV7DgCDbKM3CHM
0jrAifGEu1oQlb99ar29I0g8cgJTZD73CNA19CZGJpA9yhUqTYI4XDfesVs2h1OgriUIlG/hUOiJ
3UOBuWcHxIOBSd1MDI08UCB97G4Mbx2zihCxImKTdemhWR24F88c90n2UpooZLpc39avzwqXhJqF
HNXrgXL9MFtN+KU6HWt3ItDPNwbG+grZVemFqUoRQa81ZHxhlfw3/Sar/LAraH/4CZ1XdUBm+ku6
fgw9rhj+SFuJNt0jqolqTxLA5L+bJYfEzpPEtaWIlT12sIAWYL4mhme1y3UogqGw+TTy9WFbs9eN
2KVEolbdYTSE90K/WoF0DoW2b2fIUNe00kX2u67/GGRwoeh1w8M1ewIuxpA0ZM2NxPgpq3tWF+Sc
40kv3B89Yhm4qmtS3hF8xmNWacyB9COP+F8W3B9o1RPOLrKEOIjHcxMrI9mLZGUjLGCttkLmCfX7
NqInKAioeeLWazb4kmSi6wXkzQxBnm7uDWgt4DmuA+X+6v2PAOZOr5vvBdTfw9RgRE5uBBn+NnpC
xf/e95pxtMK4z0/GGSXxvlHSCrY+RpMBQ58mDgcQXKmWHeF2HKqGGTeAe57MVzOx29RBHBhg2LDo
Tq0ygIyGABLtD5NlhjAdbkoopcG3hDqKScwR9FdN40Zt0ghqWkX3qWhj8IB/on3F2lNMmUtmtOmq
7/v+JogMmFcQ0dsSiy5+dbrgooipAuE2SS8cuuW8ONv+SkQCosLGA4dyMHy/rlSOe/TYdp5F9nZJ
R1TTuDGK3h5r8LzooXFzBp1pBDIZw/XbNXgZYulk0q/1lEnN7K1ddgKhBgSMMNdu/Nt7Fdusti+D
8NwNqzQ/qhMYKJtX66PrY7YN4WqdI7I9jbiULhPko0aceR3AKkTYJbaljzYaMtW+cAu8AWRdLeeJ
ExgxaZrbEQBH24oQbNphtjhad9V9WhQjgcjFU51LUYG29H1l+vQMXbGWj8eoTqjIvdBKOtxwMM2o
VuhiX7rxzZfA+/zI+2664v/l75uIx1Ja/wkvWIljnSPEn+WE7bWa2yahnHRPR4ufOkc3MB0pgcZa
5urJ4EoeISen/XCZlHwPQ9KhqkHZF/KSf/bvFeIrKi/o536NR2FkfJl6iM54CrxnCevsdkpkFu3f
KLAwQUh2I1B+IBDownwimOhN3fBZPLn+/qm2Graz9ysaunxhwDxSSrLS0SgIHA9f1WdcjZh16bb1
LYtJIL5blbbMX+uM5dLNcemyKLb9gNOwilHwiqyK/ltZwuIZECXFlw3Mk1YwB7ZPHBQfWdjOYmxE
jjIIhsc+KGUZ34XxnUBg6t6DSXDk6I/i+JPXqm3V7SuH2JVYgX5nzWXktZPm3Y9UyRMCtRmiAo1g
8hcmyAdnk07VKWOxZo61dLwvSo0mkl46JIMcrQS+yDNyhUn09mK6C4VA3q5veR4HV6e+vVEN09LB
doQA9irvoMJP4xAyjv+qS+BJNYJvfZJw6FQOh8DpjFHPLVBeIHxBBusIKxNrkS8q4x53qi+esYx5
SCXkB7LuofxNzfSHZlNM/UryOv9thQ47HQRtcthuXfpJGXemJ1fayzyzCcmkRZv8ZK6Sj7Lmo2Vc
IXLeyNF1IBvgNIFRWVJHI047HpU9zPrb2Ak+S3+QdArHxMuM9/7HCCGPjXKtNpv4Sv8MwXrxmwzT
NhSg7J1Hr4df1YuplxWoPUbBV91veWAww7o5Af1Tc0LzRZDFaGepoVN2lJqZrVwaLA2w+ILKOfQm
16l5lUtJDjTBhJvSBpvVxQJEIp6tkHX6G2UNNs1d0UzgKFeRmSYTNHrrRP2BPmT1Uk0EHZxSIlsz
Jt+CXCRJ2s/p9zz/kAZ02tOiu71Y/y7Vi0J1zqe9Zc6kKsHqsBhOhr6ygEDNAJgqwN/fdJA5qTUp
577ZzpHPKh+636p++TZY4nGYbwH9jeDqfMCmFJMNpLIGf7wRBxZ8LgVgma+JEtAhQbqsVxU5s9z2
tEUGSgyqkFb+QhwkR8T9BJLyDDb89GCvP3dl9ljIRPipUizNU98B1ua4o1QuaF5AdzB7sLBejgQk
l4sUkQMiuTt1tjz9TAVVH0IgSIgP6oxnK4KWAI6UWezeoI3UKWNbuqUVGWtY2vpxlPvEcVYvGdOK
rjcyNls8+AK6PumQtp/DVacZZOVM47KfwLAMORvTjPkusRX/LpHdPz29MwOtcs05/Gfjc0jDy3DX
qRWvtTkUuFS5gI8Bs4O7veY/rE+DUawPxb+wBe7YiLB0yk+ut/GnBnI2ry0xhSgl0Zy30DothTRd
PDfTLQRyPKM02RNYt3IYYEI7loNOU3oqTASxQFm04BNSEPCnwim/Sddzu5XxiI+4YR4tNG5DTQdl
WeONgmo1yJpJKebB9oBe/MEWzVhyoUoc9nK10bxlyCwlvqf/cTOFh+7mJy711tYseby7jkyU+g0F
gJsQKM6Q3kpqP0FZfr9ROV/8NSeeP4nSl+uelxg/Nt+mRARlBtBiJVDys8Ny+mTia1N018QFi+Bq
rLJEc2plvQ6uN25jrnMUTzYmxcFEUhW8YiG6US9XjpPjtRnxD/sREVC+yuiftBk5HOV3LUbBSf45
zlLhbMy/I8yLU6WEHd3V2UkqKQewKfM6g4UCnR00v20Gw0FV+Pkgjxzl5VP/M4koxWWA6iWPSW3b
x9sPhS2UDyLGiIvE8Bdj/a3QWFtM+hw0cQCzZevPNJNCxcf6vGkCa2+msu49Ud/pZlV12dPJbtPd
SQiAc7CFbvFpUZxrS0tSwPFFuUBYF8CyUqbxIzlkH2aYnTs8HJNTLWKC7kEiHuW1jDpGyCCLDYRE
SAZ3GQIUY0MOfuJadWWyG/ZaZA+FWFXtE6Jylk+VH8YQe8RzMkwY0bgNVDNE9v8JdnefzuSfpR4q
Nk2oX3ND+Xq7z2Gl7b8qY6w+U86Nb733/tha31y8GRzmHyySZdnFcb7cTkop/+alKh4gpGBZbzm4
q+EVqXiK8RTznqegtx7YLisSlR1HoUSwjsAJWtpEnwdGB+gcVa4CvS31Ejc+HUttvDEpLfbunVMZ
Rfzjy7sxbhnUQ61NMb6EWHdI14zCK7VkZfhSsPw6x8oxlkZWcBxH+7SJn07oAHws0TS0UfgoNunL
/O9rPp633G3gx5Nk3Uz6//MZM4ebkcHQWnk4MK5VfgZjHwodDp15totjlirU7eZHNxjJmCHEVKi/
6a4nnIWVOQHXEkVF33zQbLJzzDyRCe3U+IH7KrU91mc6MHDJNPvgd/7iq1CDGvMUdDxaM+y/0jz+
100MujSieB/VQ7Nyolof0ASq5MjNgPBCX8/4QgZU9sWIbUR0xiOblZfCLDLfhEqht8HLGIKhC5uj
7MpLfHUu88eLRM5DC+/ULP7QfFY+l+Ygzg++5+ZuRrSGLOLDkvta9R9egNYvt1UtFzvI4k2cd2ak
AsWkLwnOfqKBK9AbGus2kePRg8qIcIcP6OhCox+JQGwLEEtWt40FGJnGftgpbsINK6FU4F8VRa2C
VZ8A8F8O2eTBJJ6/+bhD3HeOhSNvJzYtFCg/oWGr9Q/bdUjYYkd6z7B2z2xkeERGBcbMAAlgjZO1
SsIgwK4RA+d1Zst3cg9gTI9s20MHQKAFHtVcsnzeUVsU8l0BuyaKsxZg/YS7UfGsCBcL32RGDMmN
mrcwL2Si8i8NgvfPT5U9kVg275xkwM3fp8mtlhuWglHKANyz/mH4M9aedGoeCnvgO6RVsjGd3iWy
+1Sd8i8T+kuolijejj8l4kn73TOopBaBmuHdU0oq0E0j4tzzq07HUbPC3GmuIty+2sr+HoteCJa6
iYYFA9h7KX+x4cVy/NILax8c/VMd3fkDqNWSqWGsU0O9Xsg+FctVHDVL7b4uDPopWH1L4vTSaXUK
SR4CIMlfhehQhbQxqjBZRr5mEiwFZ9eNvL7sMHF7tN2X8Zh8jmqmMOynnxkxt7yrUrolvjra3NIY
JenjO9X3EEJhsxwDaHYf2pcAxiibdopf/vq1lF+jXCdzQ7Uz3FvKkPfHx9a5yGd2OLujiiP1tgF7
byE13o59sZ0YhoJpsgeRhVk+tPyggtOl7YvKSDHxde6sWEwOOeFPbXTMayLJNyhVwldW4NRDCnYf
N3h/sOzXgsLf2cl3jEaBhTGr+1WkBnuPUmU0wK8OMF4mXjwaF37WLjhIKYxVgrdkyUKXEkztECqY
gWC/5TARsNJktKOeLRVt94MY8fzaOfPRwOBnxWBk3uXg53W8HcTFwVkmV5UmVm6fbGyDcKi33XAY
PpaTWPsDMi2ulS8kjwEaeqseQOClg6o9iXCdEkLbjY7byjydI7KHr53mnucWQ5ozTNOT3r3Jjn7N
TCpsjxowIzGF/OMx4kRftSOS+fD1QVhkhe6OfxVD5eWVyf5a++gKwDORJBrV/z3xYxZaTnGEuVVK
UN2osfH93X91rQI7alJ3cfhbLrb7mnXcLPUVtuDWX6d+MhqprnfinHl9QTX7501U3Q9xEgiR/auB
fHHsNVqnKYyFMVhcPo8u8ZQuKNMQ2nwDIQF00gmXUMug1UNH+RSScxyGukq+xYLhw1MSOTOKz1eZ
Vbc4CTrOycfqTXZPAXv5xz5pCu1fGtqjZ2b/PTZmhWmxqgyNRg+MmlfqHwqofw8p7mhx3ptsOtH/
WPHKnQNhQkPDWQqeOvrCSx7NQsD9twQ/5OrS+eaU41WMf0gyOKXoelO/qCALy3y58CDR7MxC3Ust
0mFvq3gtMg+rugRmnZXx7ejciecH9YjzP9g4/vQeqH8G8RhSyPnIVdBApYagLmpBigTnTWGdbP8N
XyUb1Mn7S5PyCJZyAVm7ypNIozfhr7joPEBx5e28q+f9YDg0qVUUF6XuyzbgFK9Ki+RFsie1YIj/
ypvzvYG+x3KeCScm1PcSzKwjGblYCMhmCSQYfJ5UIs0dfdfvov246DqlYuY0alFAiuccEjPtiefb
GfiSwRRNkO7JP1nNaJZVhSscbC0usjRar5X1wqzJ1GKBN7meN9qlIne94E4nQTmuaVDM9z6dVEGE
O7iU/cLEbnJ9wIt949LNues3+13iaQI4w5vSco7XlA/rHwSs6u659NpfRe5lzTEvxjQaBIYsIWpE
HKEncyogjAgmBX6lj27evk+/vt2+xKbyDMzTU5QShgt0TIv9HKjJEddXZ8P56hIIs84E3z5Zi+Ly
/jlctWujrf23cczVdsNvRnRXr+iOsNj/MHuGBZHMFocDt/MTSG+5gTvQAJOM35a4Dulpy6yDbnbT
SxJQAN+zxMEd5+ZOej95H4AmiWZsmdmiLxMR00LvYyOD32ODxWRaf94X6rWeyJtAeE9yDMSENzVM
GLthtKSFrVXWkeUqYLPXTI5YXTbDBvIhqDRpXvb5GezkgJIv8u708xOvZImk5N0KMfAs/G4Bm1y1
NVl2cPthVRI7XViPsFBHqP9TuRvsvx1/Djvyr0u18rxeme/RWHfLbX1FmxFZvnzB5GLD3x/4Laov
u/7TGCd0kf/EeeBDt/ZhLpMeoOaMzWKXqEOv5J0SwCpwEcWsdTJrohz0znCp9H5Ph1SuBaHv7Wh9
tWoW9fxY+PEAT1kBZHVub0ngnuuLSG4t2QoGmgghHHQwKQbNfLSC8PQIbGWmVqCwb88etgHaW0UL
ceOmU+c1Wv6uFoepmVSUAjgc7y1jB8WA9rx8vTJIW6/0XRwSihUlFcCYMy44A3RO4QYZTunGX0wM
24YlcZMZtpXfU5ndADSpz9u0GY7cMLagSRSUva/EzrMmKQ+BLQrxnmHOCwyxz3r0K2mjMBQHJiPT
Wd6aY/zOf9jc7BO6go6PoybruYuTQGrupQ937LX+45Wt8IJ61LZKmk9RUQL2Jup5AkwwaVQpY+Sa
q6SsZvZhc4kGsFyMDOXWP7uUKopWN9FvdvMf2doUMgRxJcxKLJ5ouwoA6xduGBwkC5m1yCA1y8h2
tUkhKGX/6HvGu+0om78nsGXuDbqCop5D0ZorgpvYQTzfrcrhfRlWJAMBnxWU8bF+LfPa7Sb/NoWd
SARGkmxUvwfl5EjCdKbr1OL3tFyeWN5KAjCCaEnMR+NTjKIqA9eGlW4orXu3fugf+WTNhxDfTqKF
uahFi2QYO6KN6r29gJ5sor5DIzIeUCPXOykjO6Xh6nUmMlkV4uIvhE7s2X6XJ8PPg3WmSwkjzU1+
+AqvqClWKzo3sBBq/OculLRrxdBR2vPQI3h4CINPHfeLKMfyqqAOoeTvVCl7fcVEq/LK2/86XlJD
CokX8sKgKipKeXcJyZzlclwmRZlIGG6x0PY7+2jf4AC7O+t3ZOMVAAKV6aOZcbuPf5+NWMTEshFE
8DkKDCfkGfZmTFH2zGdiPbTho9XBVp1jNz4gdXATTsR2JkKzQWajDbr8hvrD92/0xpLSvLwDWsNF
oRv1DkaoH89R/1hAMSNPXTpArv9N3mC2aU+c/78SF2x1S/P6ZkV2Qv89Vbwff+VzNfcXKmgiuaVB
jrIY3GhS3DNN8PoTLIuoumtqzG20vyRxaMjTdw05GeKXebbWtjGf4nAW/XVbApaeCkvzR/5jVZMf
AUVZOh1rCwlK+5xUrgpqGR0QkHprchmBbvQXTIkQkhjW7avL/pedy8B7a0ODD1DTUlvzvLwyPWd2
TFRfStRORCSfq1r9llQGysuaH6pBgvXIfoO761mzUW0C6wYcpRXSDEfguNgwMPGAHAWSWvt4+7rf
awLbWU3G34UV4gjr5fMy6Q/ne9Kh3Omt+f7gL5tmonetDRZ0MoJ88Koli83rPcGNASSQOAdtJLRn
EzxKWKf48G7boXUFTvbT9+VdDUFnhmXLlN3nki8Q6DZcih+GaAx64vzYWNtNLKwjZyo81aw0BHSQ
Spd5CkycY6mEr6f0a9E9w6zLb6cnN4Asc4dcA6KaMavrLpoLMMm0OYl4qaICcubFY6Gz8cKLSFOT
nq0tp9GB9N0vych/vHSQKVjPraIoUpMbCBwEGKlIORLZaMmWWLW5jkv4ICP+mgPewlB8I2Ozt/dj
812oUW3NqjOrVMP+YUvDUCneOVw2KQ6pREQ4rOdm56g/bs37sLTvdruQmYSgMRcDQQam/8Unjege
5MPrZcJYnKJt7hSXEWZWt8M3l7lPRgp2X75iiks/ezMRaT9Tsp+UZYejwMOnsN//6GJs5oL0QaoF
Kqk64m9+5BnKNxsXyrIp5Hux7eCWO04NKV34rmzLv//c8mP2uo5gd7k/scL2aeGBkwdeQ8xAhaOL
TT/GAfzdvMCrbq7LJSnQ6iR6mjWclQqpAwQaP1JpulBGLSQ+uScSSs9PlLJtcOzf71LTGCJit6l2
dXylCtLGXVw11K9/yHP9Bx1DlwNQKa6OWOE3Pedu17WlbnYb4zrs4qOK/grBdgiFCaY2KnkrvmQp
0noL/q7/EDLP6u96xFCHH+3sdE3716q9bRSnHeA0L5BqelR2XZPFaERjUYiwYR2Ww9LXODYVwhja
iJA+hfLGwB6+/4cIyKwHb/Uv7WQqQjgXd7q1jb8y5grmjI7rkA4pFlgpWnTT45qVCiocMK7LGlOm
IpvlhgWjsz2Zh/ya5dl2ZbItVTN3tESPZE/hh8Pzt0l9JkSSfof5t6HhvyOZhwFh3stLb0e/3uEg
CSIUomJsRuGegLxpaAHi1FWn8ZX3SYigjBFHCFIXOyTEJsn8bIB58WDltbPgwM+ISw7/oYeq2TuC
LBYQf28MPRLVefTl/3ciLq1oU1t7c1K2o3b4A6Z9f0FWG238cipJCYA2NmJQKZNx0UnCpWPYhcyk
kwQ1qzz+MK88NkRnBQ5u5sH5spxvYFqTip0V8pYtg+gpCILVgqIuAEcmKyiFlduACGtRmu1wME+z
I843tp9BU+l4gt+3eIgXorH9x8zq8rYxG9vg9YZTNpiyYDtFxJLwaKL05xqfQOXQOBrn1Kk9rIRQ
0J0FxsGZ78rpFxrBRq/rthohhdbBBMZfn78XXSCyQWE8vl7vHTXJKhnxECv5nd01WbTKwP+1MwHF
zY6SHmMfxxOHsoL+WOCwEgMpwRF7doWwM+zELSL76yikf3UaTbIYhR/RNePvnwBZwsv/ePr3o2sN
FJqVcoKYC6lwYFxmWVNkgStRBVSTFPIFYC+1L+qNjOKIcnWRe/s/Q4CYNBCTGOux7iqoX70dDmcE
5Nu6L6IokR9RNn2CN6bOqmjOqpp1ppRxcV2C5gimITEQmI9GPo2Nw0k60YH0ttyLtvKiFLPjz+je
AL0V3uXPVUHj3M5jBOkDL5It1otfftf7309uGUAhD8d30ZToCevDVXdCxAVW5Tv2ufq5ntLfRtJT
xW+ALN/fp0bHn+XtlZ5FdhWE94yOI3rdIrfa/CZfXSocE1gjcbTUnONYlR89e/YrruwUs5ENesg7
/NphwK6gMR6p5ayBLQZeEs3O8TB4HXGZZZYTH7tsJUuZOA7URaH2m/86n1SFJZRYRHWjcRbhGFug
E+Py62PhclXJ34SYXEmkZmAZv6n6mpNXFkU3CKDkUgpFth960S+wObZen+AJYbmcBl9hv1VHsflm
z+E74WEekjAqxfnlUyP4xFgGDpRBkePbmOfr3mR0nZNFQRAt3riNnlAeJtyFqAfvkmziMIEfb/l7
uEAuT3IdgC1LfXwgCDfywLqlEWg7h3iZN9ybKWZAyD2ud29n2bm69ZGz13KEFbe7jKYXFTQ27LXi
loNvhwJCMqGpskXnu7Efi39TbHGxY9f26rPr8ob4DpFOITCmloXLcko3sy6RL0RuxwwgxHH4BquD
rmgK6hML4g/5CX9wkmlzymdPZ321GEarX2OW2aUO4eKytJAP7d/kxKBtIOhTw9Uu73iyTi1fAbP2
CrGBUC7HZmfErezuBistEpZyiWhn0jlaqvsk55r0+zBgOJe7U5nwAxbqzyunzasmUzvEb8lEe6Y5
tPQI1o3kAtWHNuO6wG/ViAeeLgA+my4yt8V358PQhWvxtQBXR4NjkYxEM/QQtI0WsJr0lXUMOLDX
xeAvbllcWnjX56U+llIBI48Q8K3sk0+4Z5MLmtWoy2ip0UiU0zhK4zv9CCUHuwn7Eszw0YnblnjV
E+ozVPsYJ99kyu0U7O9BeQgsSQYEBr5C4a8jlVNWSv1eNYwohN5EsodE+v/2bwHiMqa+w3FHfeku
Q1tm3SZyuA4RQHZakqklr2HXSH6zOOMjONsTKb4SBsUGj9yU0wJqFNXD3MLke5LHJc02ZbEUELx2
TgAfYcUvJ00bNjPT/8lCSTeIXmSlWW0DGjlSdM1Z17+0Ud+jUwsaAK8j6lhSKamq/J/cLKwso4yo
6cLmxC4wCR43UKrRX7CdSf+ExXVjc3rTgWNQPhV7Am07Nqu2U0NiXP7A1H3mwCXBxs5B5b82GEAv
7/mwG3Vf8UwYmMClk1iHqMwoS3wQ0MP6+NLJXzFb9NzLG4KKrlqmwSz0Y7Oumcl+/1oT5vQolD3m
mWGTBClehvu63CT+coFVj/yFtcOgVMf3Vnsmp0nyDyzSyh27MsEscBuRPobjuLRI/VAFe3tIRtdx
mQ7kni8YLj8J/9e95pB659K16Qz/Hc3xEI/6UUCx+gmnR359CnT4RiLv5QgQaT8Y9Z+sCNO8gFxo
XZq5ZfR+Wy1YIqfXQlN2q36iO9MFJYdBXtWL/Y5tzY0+lbIDVTcL1qahTGgRjB6p8jqLos3plkns
KvVodUACYejO9tvEjodTZPznN7ca0PQ+qSOLm20cjCfgKasYxZ2xbi+hJFBeLGwDc8tGBWIt9xBW
z2wti41A7ZPr9DMcdq1Ji1iDAn0e2SQ4sLAJZku4rrHvYQqbr/SwRkJ0ken6SWk91/STIcwwM4OQ
U04on4nJjcDQXtFM1HFFezGHsfB3X8M/brqX8WwyFTPpc4t9xKi2M4JyPuFWSnBC4cfTrF6iADl7
URX3rUfzCsoU3KubPUvDD3gVWB5yd5A0f2a2bgs9rnFELuCdTCU9mFtAJHgFfTwH89lo0TN+2Mr4
vzKOmGE0+wxCsBjljeHKthk0hpUDMwviWa2XSVsjID/5yNW9394lYDgnNQPe8JWhSBrReDo8eXmL
srCCUhJqjOCUP5P4XVvgcmev8S7mPpkE1pPaJoA8BCdgI6M0RdDXDqsEUOXoW3hoWSAcdHjdXczh
22Enq8nJWUh/B7hTRMYle7GFy/hVEaJM9Fz1TqO+F3iSdIDTohQ9Ookq5zlqNisoshe5V27ksVQY
R81eILLcPqaD7GYZL9IPt/1ZR7NARHDOBtCxcP+fQyYfWg8C+CoB39VeRBQ5X1YgnXBrugC/aIeW
pjML6G6eY1UWLm4akMn9IpBDsHobyeU54J+O/KVOAZVgUHNsHYytrycVfoplPwtJYZa2vCnb43VR
/ReUin02SQGhHXPe8+gpCrUuSBlwz4cSFvGxv+5xF9l7ylUdTIIU36K5TXhTBqbyQisdhV0RCYsV
VOiZwBPw6kG4MKeNlrpIAuE+odXLmV4iyEjMwpRkdQHlrR6zqZInmW2p2zTdqbPY1Wx9njuJfJjt
rzA3j51F+wWHg7Ry/QIEey+Waue0D9bwuZPfZygt7D+vQVdF1HncwOb/i+9u+Nu/V+xoHYBJuoNe
rckNkx4OXoCPH26SgpfsTukbU+AuW9IXJ/ehgmwKYFDbS0IzQBn71jzhwnM5KrDUHdLG0YbvFUKG
GI2CA1t3yAQUPKUZE/vc33KmPVShBbh9wT7IiQUnbjVjzh709dWeA0cIgv+7mDVLvREJh5w7GnKP
SnXA/yK2oF34oUnxjB41nlFK2dGAodfp2FXFQS58ezMFLh9qeqm9AsWyXPdcmxPlj/olQ39s4wD6
Mb44P2KCvPUJxdyQzV/Z2Zl9Cj8WzVutLGlkEJGLqfNfflRt1iH2p9Z1AAgXSyqEXWqTBFvU/rPT
wk8UJnCa5M7ybLtSnmqFqKt60NYqVV9jzH/MA2mQQq6GxO+BBPSonpJNtNCX0j9S+9oFpK9Rk8u2
k4Nz9FtQ1LjOdRoG9dqVMRPlxWf7QUf6fMKwMi5OOHIhaaygNC62NlTicIzQAKgcT41UyitKAMTB
DnWm/6t8f7kQk2TwGoYra36XuUiWJlNznATsx+6OtOSdsGI7KnDhZorVnW82gXVtvn8X1o9Gq0nX
qeVLcjFBDTIvrcMmyBJtxNzqxMR/ot++zuk5yEiDHHA1/TAQq9L6aA5THQewmHVcVqgTMabeeTJs
aG1XDz4QYajhD5uX+21GkwfShYGsHHhw9PMnaHcSMyglEUs3EdpYMPl+jbq7+8ok45iHOdCOYwIN
kaD4UdcMcOUU8tbbPDmnCdA4DljR5W5bczXrQpJDg+2e8U37hV5FTW8F1VXh3JGfD3zwxdT43qkR
nj5IH9G4og+eGn71bqQFXYoe1J1JxqdT0KBOU5sq7jCoQr/aYax+3c1cisPiU95rCf8rOZhjNlg7
vTVylNqJiboDmYotbhbElsvErTG0MYuC2M2hsBRV14t99z2Y4gOrKkp4h8xM2rjo6h4oaU3046ME
kTZyoK36ioeEbBhi1rjM6iG5rY6iKwRrXU+HbS9TZo4bRDQgNb+dbX7+cj3vdqoR9OXOcB7yjWjQ
LUg3CanAQZRJzGrHtoWXFKBnxiKZe3R3aXgjEt1wMMPNy/hLQOEdeU/hf97oF0MUi4h9v9sFWczT
m5uhKtUgJnAQj3/ovnM+Sl3iRJyJ3/cqzZsJhkP3n4ASvLMCx3zSS6vNW9UuGD7hIwdmqHV4MQMw
AnHCExnAAnMrlnHL0z0ihc5d9OXaU003JkWUVczJEkvmFwyndnGWnLSE5q6pAdP6t6yxLWH9FfZy
1Uuj1Zu6JnyBKjW/NxJ0KRwmNeep4PwKaf+KS/yRhp1yL0q3nKCq+UhGEna75CbgDbCUl2eBUIwe
gUbGimd51JluXQN+XrWuRmgXdTSfg5+tzk0yjQtebRPa+iKhEALjTJp7dbdzASf87LmLzASeaMhe
qmopChFkD6JJdalpnT4h70bEyZw/5uJ89QFO+lt26L1q+zAcA4QZzAKmhbjC+lACopuSyvEm635V
McK8FUsWwmUJrItvGXJEbIL3+xbw1+efatN+ZEMdQutj6FosW0mu4dWmSkZrnNOcdl/ywINKoNaA
BwdqtDm/UgmAgJoHoQ19YU96KQ8ju/ntz9EQSapzD+1nOgjdhC/XPcEnGsYhEWX/cgj2/W9K8dhk
QESmylCQC5OCaXPxdJ2gSHNILX7bdLn4YUKjQYLPk7aJWwev3Yjxm/n7KQ0H/t7uNaJsznEf1b5J
kq2ahbekBgf8IMLR7Bl+SrdpwTyPV5+sx0iwenoRB6fH5k5InnNBPFfsqPB6MNTiP/v3joiy594W
TGhfLXeXf6Ikrb0xJgpVbeNw6u2QVbh1XdxPoDvdFGOIIRrKnU1aD7JcSLMWlnQxw92JckRU7mEu
awiRx2w9nFk65B6ghlVXiBlT9eQ+Z2I6676dTDt9to6QfUd6/sQCXpBHpCKAuudI+Kbpz6RT0YIY
ZUlwY9akH4fLz07WEyqvJ0D2eJ1h2ZKUj9zqC77FKop6wE8ueriDZurbbeuvMOskUUgIlXaFXnGw
0X+NMnpL6EyBaMsDZvu7++44CUsaPG0mDnBf4RPQYx9SU9cAmJFATGGhMyQcfwhD0VH7bMhcSws6
zsN4hjXYbF/Q4FopTZKOhXZ7BaMsAICYXD9uVs3eyIMjxibPAjwGak41DUColokPx/Y9drJ8NCys
aCzIDhq5TTvSrkxHB8nk/KQZOi/rrT0H+3t2zojOycMoZqc/957DMbdMzkPylE0ove40lvZOZuPE
NgL6+U5+xD7g+kbBDQ/Qp0XVY4Aqc7NrnnXo/Yzegh5t1qAhSVKTgK+cIYA/e9QytguLwhibAULj
KYTzaoQecwSPFJWG1RxA5veIgYrf1NNL5Uu6NYL/3vY9CX1N/V9yUN4BdH2uz2t7jtwBZQaTjpH1
APu9JaSoQQe0o5QHl2POLMmpugio+FGK6AVmyjCHVI8d4qd6aqizRWs31jfZriI5aBWv3I9uEWYD
4vU/C8yhYCMWUf3r/Gpyc6u2i6zrJ1j7MIgopNk/JE/LcVduoQXmumwDolunG2bzUDE+7ihiiEUy
l2uTpr35v5IleThhfiwjVM9tCWnEgBvDnx1VikJlk7KJK05NKW7eOVMxOLHfNBP3EaH86t2L/jyd
BFgiUVZKF6YeeG+4EqCUhBBxuFvKkIgGAQMSH97mQxMIUMvbprRZnUW6Ts8+VLYs0cCJvfIUO3NH
bSW8XmIE0rugb0KB5XlqrGwfmcJMuzyQUG+WOlzj43uv5MMz6VJskMlMs0wh2o/1dwbBm0dTjRbf
57ZScn6enzC6nF9L3qcpsQWtFwlqmGLoa9eQy24Em4ujCxf/Z1jorvDTdKHZAJ81ZF6WIvuYXwVq
B3+CdJ9/gCikngrCnThLG8ruW03r5w8EhWG6B9MQsLNdFo+G5IEwgnuP6smzwBiQEBhngjQKxDe0
Vzb+QYyxD55VpVZG6Pl/HTT46EI6BAa7rQc4BIFCv67gb5W9qfOHBU7pelfNmikuKqw9whfcuA40
KXY/yC0OItODiQQT5Dwdz3/YDz3/8fuL6Zbgh5Pc7ujoyEPPrRTit+9+QlG+mM25MEM7idlN39cU
8EypGDCJClpT1d6UC8A0A0nbpIfAqmt+G7BesyO1zpwWMR+JqUqrSKJtQizZpskrpsvmqEg3RQbV
wB3dXBIKjk65ae2U7x7hQxYQmVtT/5rCMEaZfQ0mUDugK2tG2XwobmLTOXT1dd+rheDkjkUF7Fd1
q6n5wNmEHb8bgnxmRCQuvFgVzdRSuRzdkFSV7O1F4ulKsv1Kfsox820fI0i6gUS+aPfZxvwkEfoh
YecNI04/PED0OJhcUkbdKZi95ytu06XuLgN1TIQqRNcpmehnKn63VfN6TzMzGCXq7K3kLU0kBlnC
M+ZUo7OJ03TnOJHCwtIwWBdmWRodAEMW/8nHjBM8e0myAauyw7lS12STleEXv0s32khPvEQkDUmk
fygpzua/d0IVQlHJ+yWZVO2FcuTGVJsjfp2xhfYzHeM8STRFZ8b8GiiDmk+MQFs6NXhgFNx1IZCC
DJaO/q1D0DBlVoM9i1SqtlFsVWTB01Aqm9o6m5KnZ3MvThwo/2bECAR3MynpKzPkzvFq1StmS8lH
02DguojF7aq3bFyS3SDfNnOKB2VrGuvYkvGZb/r1NzLU4zW1qfMtCRcZaCzHRjNr+siQdTTxyNUq
OhSNiUE7+CPZeW+flGFRKHhrK7kCc+P8VYeinQrPmarWzezWyBO6xTgX+g+U7DHxk7LHVU1rimiJ
ntJ79uXHpQKl6VBvd/kaj9+QLn/CEFysCOgk8MPnaTNBc1m7Z1XUAyohBDhaM+XXJNQjNKoCBElW
xO19/bKNfxDt3iSRQvZ6+UtV8dhr5ztr4gOLW1QGNADtkac9b7kuTPo7dj7J6h8Y5AbvkyephroI
7bFLbqKeoeqJZY/wN/0qOU61ibgSTduyEcjvnRY1qSwsV5ussaJ4vwgu/VU6Bzkf7tFM1ijlogWH
N5onsqFZ9ytYhkgkOUhkp4CzjpJPvn4LWv+si8TrITljPmjzTunwtX2R9G2ISQDQ18hge1xI0vgb
YTBXONFeky+YXg4/QbN7Kz3asJnvUoXpyCoIsACeqs8idHSEHCQSLzHVuAkoSV8c8WdR0VP9nsJi
Z25x0xsgsQMNo5kn+5x82stD+5tukbEXlEZMRQYv2I560J1L65AN+seP2CaMI4/IAauEGVcXDEQr
ecUXeqkDtqaU01WekLD+MVrUUw/5d8+oqKWvpiFegUIiyzlyJ6t5lJi241eBBZMerMapOz3uCcAk
7cKZsnagMYyfNnBPAIgUoM1fdRDeABllNBbtn60C8Aar/DV9VUKv63GHrUNfB8ci7vn0Gi/5Th0m
sT0OvADgVSjwJj1E32Yx9MxVhkyxSbwa1m3btE9rzIQwnuq3EVDrqsTJoUm309Ky4B/I168MB5EF
KBxzfzhxnMhzyDbls+mBWnpPUqWDdj7WpsodFvXFxwYvrrBakLSMOqJ4jAaDcZYmnQEtALYxCpEu
hDHX4BW6b9gvzcdMifZdBGqbpCA7PqlH7jQVXLIhnO2jhJuuWKWfFf+fFDg7p9Lz0gqh7AT47LFT
a7LKTYWfIAfVB1+I9oTdEbt3YyaB80yX4MeL8VIQDSEskqV9PpBjo8vRIfosoNNlFdMDXQ0OjLUG
ySlgEjERelD0XK7KXToSQd3OEJcgyy5SCMSTBAZc+r9GTbQ1JQPNIMF4niD2lqcrBOCRT2nV9c6Q
m7APjoX3CTT46ts67Ce4bsXwX6UCKi0zAYM7e6M6eRdGgH48OGdPAUIYTRoVe06lc8kqOyGtErJ2
RokJ24bxx0wt+35slu6lgQB/A/NvU5jUQSdUIfZB3fqz2Ba5WeFvs04S4x823dIDJ2KaFX2bAUrK
A5BQuPNS3yupPaXmB+6SvNRBukCxZd+KPHgkHbXlmGGIeEA7XLsLcl75yZBYsIDu5SkuIufZCLRj
E85sI6aT/m2mtL8zba/dI1M24aYjXKvJX5NONbjp1T18GImMfJK5OfwYfwqrP06xStIGJ7XRjbf6
iGZ8/ps87ZjByZCMaQHVzY4rWKwULMzYbs6F0ZbWjQzdev1LvrwvxVahZ/I4wzjSq9Kjt2MStptR
7Vx4o5CBeTjv83JS3dx+9wfUlhPypCxJO47bT11GdoegFG2sAIhBILcN/stiRgIHcWaf/fddNR7F
8AWQJmsMgtxVwV53EcXZxTTNPNWLnTX6QLBtfU3Ln76uDC70yglbk1kVzRq1PKkW7+hjWlZ85v6d
BDqD1dBAjc4T7OGLDvkfZ/2G/VBXvNZKhDXZpI0ezO7jMJBNG6iaViAXwSEw9nznMveYmYWHwGAO
eYxq6WPabYW2FXI6ACi2/rNldVv4kGpIUE7uH1MR26PAGg6t+6hmex9IVFJvw7BfJ83po6Lgamak
WqvwX+KGMeTnOJ7Rd25MbJion5Qmq8F2LP6fplwbzysVFK+0J4n6B/VvfLxfsmBnecV3PtDC0ltQ
Q7pq8MD5c+ojeMFZMUK5tfxLnJQMXH4F4ChJhm0WGWNR5AB+UIh4g12IZ4WXRRcnS5nLv8KQARdW
sXKuBDVV9JWLr/072TukBDJYoJ372SUcRjllHiVUqNrzsovoJDV9BVOzhbsX8/3vt/CVYVftAc94
D9/MGuDuwHQ7wth7JwfXtco40BJXlX+oIpB8wYMlKvaflmz+hZBfX1nC1WbWvRVhFbI0rPiixJud
zUBo9/Jly5YOA2DEqBI5tUnDUSCUo+QjrCKb73R6pWgLtiDvRmu8D2ftDbc8vjl3iXAeygNRzfGB
0t98yqWCt5UfM8jNnZ+9u2fwcvGTjHugADkdeJRntzI09oRhzfJxYoIsytoSVdQ9XqzQ/gq3EPR4
sqc9ED0pr8Mwn9FalfNfoe4q3jobd4eOTlAFEco+mpgQGbt8yfEsXvZVxYiAzyC0+kLoyO37mz+O
dACBkQI4MRT8cV71MbuZNULcswdj6bM94dkaF1AQefYGVKw+lt1kelbI8168GojUUyVZjWL4QrUr
aibctwe7hTLBoXUp9wY6jtUOVUXLOumiwIhvtzBp3L9mXtfwlTxla1n+KRLiPsNBt6r9tsTQXyq+
AHC1LRvgA6F1HWco2YDR9Rg9jQbKAt6vSsulU0NbPDAUQvopLaykFusB8EinIgSnf+mx4JaBpBT4
Isem8O0AL/588sKJZFfI6Vhk9ZODN2l+Sw2zWcLmYcO9f82BR2FbEiZXoYYn4tVropzk1MXNMRtR
yno8zOle2XTudU1py/lvTEdWoMUFB1LnzCgw+32Vg7Cttl+OqfUhavsJHfpdQ1BhOHZmB/9a0mmQ
3/cjQMMXFOfb7uKmE1du7Xe0erCfFt98wEYnk+1JZPVhNIdzO3MGDWZihqSno9dNZtYvmMvvKb68
kOeVcQVAyWqE8XW1sFD4RdBk1SWCOCQ5opBCMBQuyIelxbsZmy2YYI0r/U0PYEsTu/iWh12s0N7w
tEVi8u8mCAJEtSYShqg22maLfVJBFKwdkcAIpOjfVotVAW0O+ElU8/q9Abah8As1fzqwCRXaXzLD
62UYrCQxxSLwIpVHI463L7C1cppmDSmNXJ+wgfGohJTdHa2/ag+94hYSS/K8dX2UbnYHKwlKDBTT
2f9UH+W6+9Bd4OwhqPJamdBoBON1Aq7oK+XhObaSJ7T48iFdMjHX1qaaTyhGWFExz3YdwDaX3HV/
BFBb7Hd4+/QqwlSVYx+py949rQFBy0DeDqbv6K8l7v17mUaTHIYq8o5xHuloLu09KyxtVdqzzWpp
FZVL6yunGZMGI0glj9pOWi/TmylMdj75EcBERkyRrBt/lJooZ3P+t695P6xrJC1eVA3NOQuDiqTR
5nsofDMtPULzNJW1w0hIb+JslsAkVjbQQ7v7lPtAyk0zyTVH9Rv1I3NXxdSJnI4n/ES8Sc7bpr2l
e4ajUDIucgbeF1J7kBLEQWUY/m+fTUR1HvpwXE1N2pDQIqUiXR6OhFMysl8pZSpd4hUQ8h9nUs9E
x50z8HXxPEJlYBcXpGFw1VhMRS/88a3eHumtcXAHRL1mTMEx5H4NwNRj0aOUPeKqau1hV/8L3Z/C
uh997cysDP/q1ew59sH3apoig8UVHB2m0jbOwDRn1loFwFlELn2Lk36CGSO/a5ipIuw7+lV1D+HT
mC90uSK/dl0ReKrd6R4DNioIRX2mMf3JLLMkyXYb7mV2ZlMFN2zk8RpyBK+7a0XLJ/+ky9+GfLl3
C3mYAGRcGYErLOKp4koO83dcIr54OJTEfk0n+8GDHHqb2oSW1HDCD+VgTJ2hRVhMPnQGyh9Itk7e
z8qO67YYNMUi8yhzkQEQWWKnLStftWuy5Dnrtyxw1m/X/h5KYNBGWK2B3xlx/cp2IlmERYVP1M7w
czO8dZwwtcHfEzcAzVriJW/e97Hf087ATos+pRaVd/roEQv2dGXUc2XPm1zsvdQNhTLWjPI3WeXR
hoNtNR8aFsHJfHPF/Iael+/0sjrPAeAck9dYVmglmy4ujrobWPX2dKGsiWTQDGdvZzyARHt7+k2L
oQEbAYNnXtf4bOhvsBZ35SIb6pv1Q57qbTgORVjPqrXpmtp4g4SjV+0qg38sVqPal6cdynwKhlNv
gvd7GEkswRA2VoDwiI84TzgsfQKzZnpjIoTwphORQ1nxoqVKSOt5apH1JT3MsTyaJGIjc2FwMeur
JlOWVTv6zQC+jOSpFUqUYNI8PbM8wQ17P23Iz3v1EyoPtozvdwApvjnF5E9O+21AdBD57Qq06ywo
w+3CImThK26X+iUZ+oNmNeuz3b5YVLy1/1csWwh9x7UUNk9rho/iofOoWAyfZztwBKsGqNYEu5dS
35YMaj9Qp/IFplzKHQi4MWmymveyZVimoPM8/UY0O+2KxazkKi9F0pmrLtiIU4CI5doajWWGv1hs
Sc+blpmZ4wx912G2ptOtKe+qpZVAHFiclPRKkpGl8H9LfUu9qLRc3TuskDu96scyVYoC73z1oOji
HflTm+qLPDtfGdTGtBjdiYCh2q/w0wFBvkcR7S4iocpT4bqQOyiRV9zgWeLD05mzZ8d4QPn2q1y4
4bvfTpZKPj0UMGWqRfRL0oivtH/K79QB3PgtBAPxdDe8iLenIeOBTnor9L4xZLa2IREZTBlD1Ba2
Eok2mPv/aegLryhpg9Q1wL4fePU4qjjUatrlKC6MTEmmxTWaHPuHKJC3Qr6WByNa01o2+Yi4XnEK
mX2mL1thxKMwKe7JQHXSz8ZQ6gGIXRcTmazLOUUgoFs2E4Ji1BS0c1E+4YR/KwFy4rUo3YXzaadK
hDieyUp5FIW7J0LK4LXvbi83nIQJSHCR3oDEyhEI0UjggOglIXxf+36104s0u81ABAXtp5HDT9Kc
pVY/LMd88cji9gVQTDsMyacrdG6615ff5eE7/5yqEw1feeTjfhi5QrUuOJczPespUscz300/sZ7a
qxJkSJogR2VHn1UnQY0FqBMaQdG7fyiostRATuWWQaBvgEk42T+27TwIBWzXrBAacWoyBeV9YqX4
kqjLWjrdOMbRA4kvFm1QFw1kQDrpNG36sk/tKXqSUo4BEYQHQwjjlX9q8+DFE1FNqGF2PyGDHn4/
69ms4SLGPUgnaS0A5UtJbi/TVHmpFSoU3niazzD2ItAzjOX4Qd3952CDxHokMfqo4f2ZcIsTnYI+
RGA5p109N4L98sKKrlyp3M3L0K0peE62nBzaJDWcPQUcOAc8MGL2giy37SDeLDCwbKFkQN4JL74W
UsM6+hyK5TbPfG9y+l/7XyvayQgix0rE/WbSEVWknC0KMUwNna91s9gUd7zfj46IriQLnQTxjgYL
coyUKNYMslCJSdORRsLOjOKBWC0Ih2GXmlvGE4k+G+07Pr6jNFYpjYY8WeEObeyPfDPBxIrFxR5C
XofG5fPROHZ01L03rvP9KSzNWZrfMT+90LmzNEvwlxh8OUXc77OpPv6luhZLnOvu/mFEymSf2bt/
QOIxzXwZpRRtJeTgLtbv4XxbHGCLYUvjX0Jig6DWWLBBhFO0upVGNIWUuEZhsvbCejCrWpjt40aT
fRMltUTpimTxUZBxre0LJuVfUaARZ5t2DgdP3IV/BSjtnrGmZoX2V2RjxIu8hpY3C7uSMOqgbPxF
zSpbU3dQQxQcWyBZZSv85WSwRnY7XF7UfMbMLd3MMLIWaMQGjGBqX0lXeWltBFVDsWQOd3aKBtyJ
rgYRfG6vsTrVg7cvBJjEDbB0WcFj/ggyJ5yt5qN5RVYp2AszaSsTpm0sot54XFKoArvEZuk7KKO3
RYg/Px6NY3ScT8LIsHQRzyJxd6e/iX/hL4NXlIT/98jwpMJYoU8hLzTuNjdHkv5LMKAvePk1V+/R
xT6gA473QoKE0M1ax2ECap3rmX9SkVJnQYFPDZ3OuqDVfRVQ8qCqE+bpzVlTIaxlKwVl1fg0k0Wx
QsxKReZd+tU6l4DRraXDDEp/Ik/tJ2Gp5xuH2MexgZPVmp2atFYRCKISd0syFmWXsqAmUHspce09
yqrsoViTjjXvK/fiNHcqapfjZh2lyrE/QKsgLIZn2Q0Inle2mKes4fkz3X/BGie2Q3KAPRdsi3qM
L3O8HmlPSUPfHtF0ADcJvFGPm6y33BP7xl4VNzFOUeeLG9GLdEFICScW5aTGkZWX9CNc1W6shVIR
IRIi/9xRkudfm3XCvus9mF5v3G2cE4mo3aRZhuZdWzyWzPwVaZGAXmXBmLB/Q8RIHBcTxwxdUkO4
2yzoIMjMkoDnoGrJMAFiic5HQYqGm2KkbC1L4ZfYfRxIFRS8QbkRXGY3IdvG7gRgj5KhVWFg/u7Z
fiZaEza1/EgDwBSAzvpqkL0/oMj2OsT0SkuIIfnDQqJ5t3qjuFvLIS7zXBvcAMKaTEexRwOZMfs3
nK9AJMvJr73WRS7cOhC3TBTaYqAxASqIuTspIvzuLQ09SKKhFNL6JhwQjUSSPEkq700uoJc0LrBS
uGpKRNkhwAxdNIE30Y+1NVA2SXgJflLywWCV6rD9WONnJqxwkIbj34KBLeOyPVXpn2toFLKjz/nl
U/Gez1b5JzSr0+1Ztm4sg5G1LMlx4epsGCpyd/qVzSBhEwy2Yhg2FctER0ztem4HihNfGAL5KuFh
yVnS4M+lda9zwQSa86rHBsq8UW9KOSEDumgtHJ9aZPlp5jIl728C5TaqOpVRNcsh1dRMrrhJaWe3
rFh8RPeB+jY72RlfQqqyzH4F7b+wASTe29GHX9Q/q/eJdEbP1KFNF2JuhC5uDxhRR3hyzDgOqhV3
t7gtAnyjKZLvGeRqDqIcmpu/YAn/9zdOhi93k8Ddzd5sXpuFmmMRRp8AmRrdqgNMxKQ6a9M+iO76
kQNAsL8y/b0e0LvlTv4DrSGDrWMELM9AuLCsPcX04iNPuCb6jMota8UJOWzGfY3noKsKiMQFgCLa
3g367M+WPKi/OE5o8jsDKow2bp9UP5iTOy+SzdbXObxGot3LUQxN7EFhyIcp8zH7gqKQ/Nl1FO6o
jYt8EPX/Ec9IT2kEuX+nw6k3s3JvkSPLcV8cd9A3iHL3FH3eG6lcM8sdRn6osr5qbIWX2lJZSfGE
W+1nVGv0fnAPsEx4Dji2XJd2IdpxDBHrO2CP2iRHbbyhTjqqd+afV5QzzBJwJuRezptk6bgXVqEH
UMJB+YMcWPf3BzMHVpywDuhaBH0TwdCWuIXDfNPnxEJ1zNMTA8Tzh0w3v/J6goQn3v7cffF0T+u/
3U7EUuxoel4F8ISrBd75pW2TZtL1thYYlXu3w08a9U9f+MVTLY3Y+Q1fU7G1WlWWkjjMKedzfR/r
1XmvJYEFCRvtZV9BeJ/QaKSrRy4/88nJWvK7iYVUxT5CAXc8oavnbO6ydY7jOOTpRoavMTNWwFiC
mQCkBsctlbTAmO9UH0Cdk/Gqo7S+Ro/PuIsjeSUpGnnm47eHGPtsLekP0QudDzcWgZWtg0K8VeQt
A/v2yBY26p5cPGXPBixmHysrRkQAgu7pFdfN8RUEVfJYsEMbHKzRiD+Yjb9q/S+b4ax6M4qlKzpS
OH8tqR6K2x69a1w/U0WGQriRu6oaEgkYgDr3Hy3XUFGj/nvTFY3AY+9UD6Kkt4h4XKZ4Dl4rvcrf
WnQw4A5w55v7Y2/2T29JBscqpbF+Qz3Ucm8TcrDowH/YRhTdO7sL3Jda+F5aFNGY7R7dWJSZmc8e
js9dOptqB0zoGD/dBPR9ZZ0lJ53za+yjX38oUu5MmECXShaLo62KYBchdV0WPBO/p1zpUsvLLlUa
c0jDTF8v4iiqOZmOiqMtdt3sUrVHgGcL+KYctj1DVbFXJsprD0h5gf82xBMyF8YCDSaN2FKExUOM
HMIzUOUeobpB14+34XgzZrHvwF4NSObcdFYhsGiCnklAFVhX+hE+dkOqdyNWUfS+AueDVxn3syeR
/Uwpahutul1I8eT7ZA2tSdsoGgdPpW6QCAjIi7ypo2wCNRckt6cAfieVcTmNpGm+YkvA94EXKoSW
aUGcYYXQmAUXyUTPDdoDiPusF6YAHXUa0Bh3+xBztEu5rU3UkD4e5MKov0XrCnPjo2baZzAAIA5A
XxInBmnTslRBO9DCP78z6CcXOkbf2COZF2JVrEQfsRtwiH6U983uq5wHq89Rni+JQeZqfQ/tmMx5
kHGqi9Yk3Th3m9odXiNggg7DjPCcNOgl/MSNu9yfUM5zdUJ9XJ1fD9C+o9WcQYT/6I53jfvQPv2B
z+bY2nYAl8ztgqdiQJMc+x88J8ScSL5xotfrgGNkoppAnAI1Xml2rNUstmrQPEbKZHU/9C7Pz1bj
8Ecs+DNqW6uZ4wtJ4XWY47XLnQbo7/0rfBpZPsGTDQRVWGd5pDvZMn/TeK3lua6lz1u1QEZB3wNC
EOSDadGH9BhQ13Lqtt4g47A4Gu0Y/sgiR8UWSpmyTgJxgm1JTp2O4RJtb3lUn+i///ve5oJd6IkT
KXCGR5KrTda0tUnHe7X5wInV7pwS5NCs/MRuQLjUpFJqQ9DbtZPrwIRvZa18Pd4espm3xi6cg3tJ
R2SUiC+7Jc/e3KgSl+wZ9Uk7+WFoeWplOx5eUeDDAOXGvZxhkVaZsZ7ohDs8oOtvcFPgEOFGfVbA
ed8uKle2BJoZILLO4o076YrJKa2c6ZYi1o0eJ5zapCsl5aDkAhgPWETlrG0NCh30hszPiXH2hfdd
WsP6lG59AVXPy1Q7GKJNyXmMGNIjqpkzWseyeEesTZvaTzNzPJ2j+Bst4J2VpFeQxMIt8lWJWKg7
j7wVl/Hk5Ovx6LCegLWZjo8o1g4poTU45AZWAuCSR8IJZBybZ2lUZUWxwonqVBWLEGVVEm8I8lDB
XiztPiOZXuEN1EwS5HOTuJKAK+hNhAHx5lVd2EYjSfpP0OgSD+2G2Lrq7hFtT7HBFeUXNLk5kVI0
kRYGcEhRZmQY87vh85CAAr4mkFbmbDFqKsQu1rVsFSk9yXtqlvmFP/Zmnetgl2+Cyv7nUDFc4EnB
MTET33TqMxwK7QKzV9OLz+mBMETdeQ61+n0pn0845/ALVVhIcFSRGXiTGA5vf0DR9IK9ce7Z5FB/
o6oHrk3ODCtQu7HhoU3aOOPEee9bA6z6F6J1ylu5jFlwp2c6m6FwzNPd67WjDC7XC/6SZ0K8J4lz
oJAGWNuRYDIIYEIZhCEZXtjxLNutI3QJTTItwz4gWjJm8O9znbMYUDrP5q2G9ndxG6xawVN2Mpgt
GXn864v2gr4bKJq2WgvfJcxnlalX1sZsVQm15hzFNWe9d40smZN5nGr1snd7bHGpgoLIPrB4CeMP
Nsagg933qJivFN7RNMz8nZZ+VHv/3xHYubwFwbxT7/rkREJjuKCqRyxP4Xzg/WOoYwjnT6U7ozN6
OJOvGOZ6mkhkQRXxqs+LmG60bjly2xjbNLk+NqsiJqR0JSjTLZKj1wvuW6jgtdLK51Ifj08PAYLv
/Fj+bj6Q4iqMW9cMPdmqhgV1WrVUC3HhFg5Yor02fj8ERLlxesWD6g1wn7HUOZEZPimRwhgHXl3x
iMido1B2oFlImCrFDvllXeLT8Gt1E3R60RSSmpan4eHXqQIG3eqCc2uexmgBPRkFQ/6+Xp8cBgH2
2SLpgOAFh970Ux0cW6x6EYwFja4pcvudYhCYmBEJLPYvEFnp43GliH/hfELHVWHOqgrxufU7AX8a
Bkhxu8HRyK8SU4+hzinykBJhP/iUeWoB5riGR5DmdrQiH7OQBBPgGCCKRogyR84hgniwXkmIqP1V
poMWoQhH4kb4r3+EfBT7gv8UNStFgyUZupsQx4Fo1burjR3yoN5D4VpR642lF5iX13JBXMeIy+Qu
nBXHDpjz6Wx+bkizQK5CdElSDzwf3p33mtQu6OUBoW6qx5FPSNBId+lYJP1JzHHoopaDV5fko116
w74ssa7aJ9TtOf5GJn65hg13RHi1Ng50gofdvVKvKGqD9DcyrRGCfb88leP1aT5EwbYtgcCmB0oQ
zEn3tV5/ZMHwtYCTDgHXOe7tWWKSoV1RaukFHOzvQ4OE29ZVgHk0KDT3z1tUri/olPxkKVyKaLsx
YcyZpzKXz/jtflEoE1MPMHJ39kZF3C+yfeJJEsHoFSGyOfI3ypZUK65PNgI7wU3iUKf97DhnNDwm
TOkpjC+icA/bcmxuEI9iaFya/dtk4Jt54+Dj4t2+wtEY5aeyQs4h45SnYQTEM/u2QfUUR0l7pp+O
waQlvzMo4xv+oRKsiybPs69ljCZeIVQehQNb2+FB1X1fxV1rTX5NujoQYkKYeamVVRpEMvAeNTxX
PzT1OtHvlhTO6Gh5y5oIUZTtnGH+O+ujCEgx0RpX80l1g6X2JnZd5nIEI389sXp66aE8LNgrUNU1
NoG9WEv93P5sKFWlHrFzMb10oRmQ4XQ3t0BWhs/3NWLW7CCeRZYoHms1NHFhqR69ym5shQr7ZI1s
ZGuyroUoU2/x+S2kxnlyPYniRx7rmxG7LLKffyGF3MpbnesBdB82PMkklLz0cdbsVhrBCK11lMKJ
efHhv0E1k41ukOzC0d9e4j7N4GF2Rs3cNivSYkUNlk2GWlq7ZgQ38y/63Wo/htkQiIT9gkNXCf0Y
ZxyrmJQCZ590vXM2awqXRAq543TAtHYPVZRpcjuZBMSgeg4lWGGCbdnsRirCFIGH1rTT4pc65IOX
HNEHwkcrx2vDHzoIVjAUJlSozD79eOkrqCHqHCGPj8R9a8q0TwSK3Q11xfpYN4RB4UO22N2VN0aV
994lo7fEmM0YJ8wJWzQMrVYqrvPTJoVNh12sap86pbkWPTHlEyaCgf396TW4eSgDkfE0dzlgm+YN
uEuHBCV4B41X7ILjtmgIIP78sdIg68r29ccAcOZbDu80Ggj7cWzEu6XWK1tVRqzLWl+gKGmUafCz
bfmaV9nFcIdjkXvnlAbcBQIZt/qqTaIq3R4jjLZvnjsTk/ldBwe2kJvGTYP7qAp+xuCCVOMGc09s
BykT+vnHLjdJXpz9b4LXejBniS0w+I8ZsVf3iuUZqGNGIBkT1WgIQUSezt5Nbnfgu8qjsXZJePQ9
sk3NBdsM2PnwSPTK9k9o9Kyd7eDs+ivkQNTKUq1NMLmWbxXq9dNiOltcASxahF0IPJKoeEfb0cTG
QnaMD5aPyKhrXLblbtDyp2t1nUQtKqa33bEoGQbRWIy4FH8C6okmhHZQytIoYfB11lfXLPu1eqXh
kyOjUYOGikSkTt7W5U/XlrwZxHhzzwlxlGCZyJLLDzzuljz34+kwNIAzrj6B1TfneopG4jqAa7kJ
gGYcvtnhjAQFGHicV1qifMOdpV/hUq/xazWPU3qd/EUTnGsZl8F7YPf3plDhb3HJuo/UPC0bglTe
PDkd7xRHEixbukds8+4oXgZy16yx6f2LYXQTS+scwSfvm+DCYKm0myXR+xDeC6b2s1hz93/pdv9B
1jftNIFvqJOIDds/g5vdnbRy1Apm0i5qwaA5oFdxcXy/0H3lECzr2nO21uJFdeMS5ivvr4QChxAu
45t51cw+fj++3broOODkq5qN5g2Myk4L74uXJ2aPDFD6ISy2cLpk0p5dr+AcfM1yZ8oTIG7TV1l4
DiljVeIqU34LvVlelO7/qVba4iJByEKGJgW2FYuKYVPwcCtqUnpGqUqPAXSMqOoWt+bNesvzwndP
Ig+CHqlVk54nzk9mC+G6sRHKcmajd2iEsMoh3QjJumOMhLQz84uUu4a2UhRReN+9JZ02OTcKArZx
ZQlNgjrm2BUKK2UKAoxO2+oUFgn/PTBRN+sRcO9j8CvTTzAImeonXhDz84MG9NVascRzPbvLvPfX
pQMylhKabe6XvBgQQWqC9DcEGzTe3bfIG7ApSCbxVgbcvwyS0FRrJeG/R4jO9DyBWutmknqJwjQe
aB6pDSUyOoVsh/GvMQhpoa9oWnBHIesXmah2X2JNEu2URxruPLsTL72uebLsho8IyG0tJSijc49/
sgwpIvcGa/tg0N0WpVU/9xDnrEA/krW3DT2HuuglKvLmiz/d+L+OZcR7JTooPfFQhcEFaU0Podhw
IfdXyn0/m6XhBDx7+FVAJBBY0WFAI1N0lBEs56+bj5w7cn2/i1/5T+QVjVTjSTp/AhEi2sl7Vjet
ZtUxF77Xw6mvqoO8S0urUmFK+GtVVNiBm81dMKXFsEkK/oXbLyr6EKZWlc7egeon8qYsBMt992VT
z2gu8BqE9M4o/uAtPBvOKelR+4ePMwRWjNFONLzfTOsLzklNRqIAZu+ky/pwFDxTi9YL95IOLMnS
baglXf0z7s5KOoRP19rdyNgNE4fafSWkXGi2FShYgPsp0X25fJ4XBIuELSNKsfjl7f1DLBllcBOY
chN3YMzidBDB0LP4AXDRYR6KgXu4uhmEHMygTLLiUah0pb3ZlfIP++yIESVnJWjt9B72NyHF06S5
aT/YdlYkmA8e6gEJhdQDAxTNtidxbqI88fbKCdfo/tEgXrN1QWBetrEkKuNdy3TWtNj19dxKwXCG
KQ6TMWJhKjaLYmYDHEZbDZcqBujLJzL2Etv23JrM8SC1VyBLIyB1SHuNu2tdeWML6ZsyjDf7dPak
BWkJqV4tQ5w+frfI7j6LzgxUlHsBWdwEUmyLm+XsAEt/thFvlHQbuWV6oFYSA+gSJu+g1c0/K5FP
q8DmcbDumTO4vby0157ANT+bgCSCravTNMT/sZ2U2SH3nMeyWQYwurWpkGWSzmNa9QD8HMMBc1XI
0Ok53gvPiAm3zrcx/N938IWgWkeTeXnxWGKIrRZxQ5TjZFAmU8yiLVwy97+qH25nz9i+U70G+Rpf
6KVnia0xkhA63obe19WHteuukHEQuZ/yR7UmcxuyrN99g45VZgBoQIJ0LFS+8mL2XvGLL6fDWEdT
1sjNQaHcMC3lJSoL3Lo12kbGS9gqAtbFy0A6ycvRSqMXtWUnhhLFvO0f4+KqTpQDDYL8/gf3OxDU
Cf+qPsyrJS41il9+i9BpP7iaO777r+yVLvzd4vEYQBCsQKSHTYuShL3YMyCiMqZf4BqhJz3Q2Tpb
UcYA2+gd6oYk2TBrJsjNWlFEjbu7D1ApdAQZIZXDh9G/suURT5e5hwC3TXk7NUGgwXxpXA0PnTZT
j6GKJUu4HydjIw/QCM+2b67xy+YsfNqucBTmzwskf5JjN5hg9uMPeo/A5k1kYpHsXxiGlrm+GMyb
nUEJoH62GRvlXKGXxzTRrOy4p3Smp+hlsmbHEAyG6/nK5S6FaGOK0Fn0p6f+e/6HJxTGvua+YSgQ
lU175iE82qW3mGMICQ+lO19ZV0r0jkCqwEAvdCbERBQXYQ7otK6FtxxRnszyZe+qV/J4TcJpRyk2
oMjnFmqywTCTYvJCFWFhmRLLSNd/4BCy/hOP1UvGGT8E2v9yoFnDGdi3428OcKADZB8qCosTyDF3
8Ep8EKO5MUa4XgrL3EsyShjb59JyaHmMhp7ixXD+rmkCGMeqTIBZzC8mOu2ldAwuLdZeI9O+igB4
9t6SQE8EbZn2Yxb4cijVYvyUu2ugCYHf835VOaQR9GYBi3OwO4jCyjjSgN8VUIRgAzYeNMCU7qOz
yR3ZGu+3URsI82CCho9WsrujhG/cLLgnOR2W+U/Ax8L0DKtpK9yBY0AU9KgMQGziU22ybUTXpL9z
hOWM7UqqdUBt2qjK+ZlBOTJerODp1fL9VnfXlsDgYw+QjGOKfmxv/mq4GU5BX9a6iXOK0AoN/zEw
eQ8GQo0In0udV30QtcLn0+jCnfekIn/BwRtbNTqtHuao3m0u5icg3A9x1kAoTlMtFnxOw/2QUSEG
auEmW7bj1PnU2sUdfvE+wNJGdUJzhi9nTSDVzxld2PVz2Wh9BQDdSjwHDdS48NdhRORoFfDFS0Uy
AcDh/bwPuZwg5HYkOU5e95sBse6huhzzNJ55nWO1127b+DcWK7rQvmWBad9dIzoukwxaZaSvrzsQ
q6B44tq1/s3t79Kf+fDLru23oB7FtO/xZmQtDx0vsk6FfnlWUW2svA8Ms0R1j9n0wc3FgQfhXpEK
pocXoqubWaWvPyzl1pkM1vYLOftQndxFBB1N1rYSJ3JWUqb623udD3KoxSRMqIC2inGWorGyi4Ci
aI1e4xkOgJZR2N1mQu88RNVmFVcntXnneqlDfbTBJpAV19EZLeNSqxQdovWHQiECjy1nr84rwPRh
jxOdLTzMNUvD/BxKHe5BT8jCbebzP1992rvMRJZkyDurE1ghoqt33qgQg17Hw/SJ2YszZYfA+OHT
YWJ+SABq9Qe4QEW6bl9O0XW15zGDyimHZvOMt8Sk1c+f3sXLQj2kSnytc9U2wMFHNC93bp+F71bb
k8X7eCnXkEgqWqgMaJ4lpEboAeoyll+nFVl7kNcoIlUZdvrMQUk2af3EuDR2TZCbLEvKZNK98b2J
zzde/z4sG4RsyMaSpAzc1OWtYBE/n2qnaxue923qyjPFMdjwCYRrdmigu80ymA7Lkml69fcDQyz3
c6Cq2ihW50GRu6FmFhSeXfrwAmY9t+kTHEQsA+uxnBxcy0BETHZFzjQxRNtcOq8J9CxJqAU8WxVT
Tmja0MUX0dKs5lAl3+Co9iVho5wzciyeJ+DBIXb10l7Je0d5SGdJfAcoOXZa+I5t4m5kq3M3HutQ
v/i7S3ZGUVtkvYtpyzSpY7wqtttg2spsQiKxQENNQJeE5InoTlpwiNwmd7qGSEgL3H9AfsQcdyeS
4oGlKejV08JtHzmlKakhq/qMxqlVngxy3Qv2/eI3QTytag6gf/nOmF6YGoJa8Ai1WTph9+TwXiAY
IfGqlbTyof7q0DvEV0sWkj2e7Uv0q+K7TRhF9ZeF8dgnXM5W7aRF8fN81HzmtLn3uRWL6b5M/Fob
jaFXkoluXOMFiHDkeVp8IufVD2IYJpeMozGURCOfLeY/5a+e2DAYHP8SGcYhts8IcpmorHilUjhi
6ltp/v792cmH2GQJHTDWHKlz7QIA9C7Zi2qqEkLVX/rhJPT/cq2KRQgfZNkh7qFYHeUzufHbfVyd
8u3qe+W7D61MWqsu8bTRpRLDw1LJaEEUPd/5KfVj0C84j1Ztt1bBk4LK/m2oO0yRU6zhMXOwTSdz
1t0UyQqRIzwkhXpVBmwV+2ZUot1eigOGS9Aw9/RMe0RdvvJiKnx/+JWidPPp+cwX6dgjafiZNiNq
0i7NC5s8lUtMZ6vnSAemsLhP1+gWL6c+soP1vlnjl+DgNuRFRkOW4kU4LqRxlB1GFL7s54e17Kg3
oQ3LML6YJwMZidtod1Auj/SAKlXL5GXLINz2i8LTDCKve1aFz8DZyGMZx2sHkB6h8zDh66p540TN
+5t577sFAOe4v1KjQTzyURpjC8Pko5i9QVrRGyLA8PrH02wRDxeeSfQnYxRMy8oxrE+HcjGOLlW8
qJ/pIWHsQNGfObsGdtsIS0oH0ouJhRs43mEJcCQ2Sa1huhkLNJDGHoTG34GE5mHB1j/5TURkv3nq
Xmn2NZrmStwZ8LR/T9eTFempiaVvp3Pq1vIBes4MthOPf3vLhK/O+bJOZL/SQr+L0L8dRZdWe+In
Lpe0zLmnqc1CCwCOd09boBEXO0/E/XlzUXMdgeEkNofMAxg0ZFt5ANbcxZwk20Mpx+yYEhKSMsXB
88VNrehlIl6kh5ZQscH+N58kDNACgNGa5hPSzuIdVrbtPw/nmnc4X5nlEmqxcef48zBu06UWeDs7
WRAt7nygilA1KC0ADfceCU1WhAxNlep68nMnA+GlKkZQCKZaOpTlGDf2Jun5JhTBFBQcvz3ekXpR
EUgSKsZuwArbNUhZ94KBAzSpoV+8W6iqpFmk/hQej7OMfXViAJxLcqU3e4+Omzhje1cs62ZEjzI1
21la9YIrncfmWSGEc+Pz4w1RHK//sw5Z59dWgL9Dr34xYwdTDw0dRXuqabE/D5bzyH0PA6lti2bF
pigG+GiEd2m8+pVgqgITcXtR76kSxQ9zhttuQdXF6WJ0eah4FjavBFBZF1bEUZBm6OFB+qOtURWU
/YQgjjdAboJ7n3kuStmuCJyPxPnXRqVWFp0hhnBmSOiM4dnBUGbZhZu9VahP7QLJLK93aT3zhGWt
ts4NBy1MKOka2ZWMwsCiMGcqENqiacaO+/gO53sioJ1nrVbms3XQUNXYhWvJH/0KC0QInu5TJ9IM
ZbV2FIgfz4lOSzgP1c/zbzPhMl3a3rGb6LQW8NlqO9TG+2uBRssZzAqY8awC4GJHgcZ9P+OnOVHC
uFEyCIMtEzTBHyx51rv+YfY0UfBuFbkbeGplK/D7MYnMnOTO/uShjbkHzOOmYRxAlVa3/y+puGYL
MUaE2GwrE+Kkcz6S3ngDw78xM2HDCkXSDstY7KHbxwL93FJLpebNPNUQz4fV4MR9+ibwkJ3eSZOT
1RnDz+e4TRmwpXbXj0U20R9TxfczbR6zYsw+IingEObAJPJ5IVNQTEL+4h3lJqGM4Pa5Z4AuoPuN
lUuWSMZ3DtrlLlYB9hVP52xNw7EuU7qODMS19BvMWVEN3El6Pg32U76DDRUksT4wDB9N8/OE3VxV
fmIahdKeSDQaZPb+5mjBAIQo77S/pJPGwHcWg1PXAvydAP7vensk66ONGIIqEDJawj8urarVdGO9
+c6r/clMa6iIVvH3z4h4CABgb5ZJ2/F83I4dwnwB71cQH7m0oPrpwwOb2d3uPCR0IvHxmLFu3avg
9JAUfaxsf7nflpDOQJdy/VxKxzsMj+wvWm7KjCPDapTRlan3UGCRhIfELUKivjLScDNWominc8T1
Gqt8mTt3/0UwnO1hfhk6Wez/Y2RGF9zDIeinQNLRFZJ2PLIQRi5iCzw1NwZxlSgIjTSBGGkdUFm2
sUouVdp2FLJSDcgBX9kWsioJBnXnG/jeQU3qN3j099SAzvMpypBM3vks9UdIADLEwCcKF+nfaVAa
kcPUYsGQZJ6JwQpY2p9TBjqPCPE51RRphwr4ATfIqzmB2PyBtNpMfq+I60kuuTMp2CVWYBQOBrd9
EjhdJlz8RVD0/xQ5HDpoEnb3MDesLXaDrhZgIywiroWqEzU6SM79Za+4dPq4baLzNLJpvqEN2W0G
KmRU1a4TSpFPxEuLKd6kiu1TMpoVmYKBfeCOK9GilvoKiAa/xwGKjLkQx1bnWlM1NyrR9S7vy5JM
UAfrYenWCAaTlPfEdDLwHhCku1CKWiknvCOLCzkej3X7DCKJUWzAM0Fg66QBMjn2jihqltzl2PkV
palHyrjoYiYiUMszHyA5ARqa0gLzfjAPr/I4PVX/C0Y0VfdstdoTfH3pomdOg350J2pcxlzDB6c8
EhYjkf4kBuVQ1emhAL2aRSCLW4/GNvoCgKoNNf1zGS34r3DDf/c1QwnzOJU0eRb+8gFu4LiI5g6S
SEE66QbDN9J04IXSgp5pLIafwwrgBFPxe1TNzTe4Wez0W75MZx5zdfvNFZeJ71K8DKgTwGuO5ydG
Pz4AarP4zchWE7Y4fuE2GE9qQOcY9JiVwbbFgmnmumtws3lKqaFntG39aW/UYmnoog05XuxXuRTN
OA+PZ+mAG9D4aNGQTZqIj1KdS70p5PMKeWMxAkzN+Xv2r52At283oNbJa+WpgywwljFegEkKqB7G
CZkOT4gv8rDLr2xPsl0pS992e7b2fs4qraUNSQeg0+TTUWxTikj57I8W+CScYInqk4XUrIHokB6J
1V4FHwNUVcw9QmGGTaLX5upwONU5Uix735ToYyLsMGOnVVA854JygGhy4zrS6pJu6KCFVkem9sa2
XtlO+VHD4WuMiQhoS3S5X1Cp/9OHh/c27TV9/hh2YtV41lrhaqHwke+QSJL3pfEtAgKqCgp0zYNq
9nPYLI5YXJHlyuKOu8os+33QEcCt5dhp+/rNvCKA+VLkl+8Ysdxp/MtO90TQPwkOy67oNt0u4DFF
Voe2jozrbOP74rPZz9NHiHJdlGFTcetHgBoBLIFlN+hSQSQpK76GAGeTugtCKhZioNLkcqotJKAE
V631L2IuWiC+AZv95lzfLmpr95HDOSiHb9LnR/KQltTgZZQ2TRlDVpKmOys8+7vJZpz48xiNXffh
cSAvpRwnQWdItFPLQrE9bx9p/cUmgBctQce80AuB2cjd/aoynHlAEAguyTRML94ONQBEoG0QQZkX
JoyNeOiHB5Y2u1IzGxdh62fDlAxAkXB/cBWM7pO9VXrBfevkAjI+iQLLE9s/CIG9KPYQrI4Qzkdb
9uX26f5/0UgOfG0uzWRg8vBpLKFoPlglS0V86gd5kdXXce9iPUmzgVPG5LXmB0NZv74/dbF2rq++
MOIxvY8osm16jgsSOx3GCQeD5ORSc9Z8BVCYq9pBJN04zX+TRo/kDHuMBweR9ZiyuRGjJT/gLBUA
WJVWiOfx7x1AGCs5S6ShTD+/3eosWsPRS7+G1i8c/HL/i4YMQz4QB/Nckigd/vTx2jkid+1dMbwt
M8hlFyHK/kExhCWCio7Xn12gDY5l8GffQSz36aKvBjSg83cR13EBDEJCCWu/6hP2i5MgutGK2tNb
2oBVVNkp5L8chuIbniexaRFR2fEYhtSGwSESsWGVTG2bwAODXwAa+h7VILa7YOrw/g1cy1PLt2Yg
ScPSX7kjy+Uz3RYFhfsusRZwnqZ44vW38YE1vi6Bd2Z42Go96A/Fx4mhcuqndnSZqX4J0vqyx0O8
NWK2gE1TKLW6YB25oBEc+iKe6mXOrexXEAy5dseF5Mb6qWWZk/hbzJEjKrgR7qloXzxSFMgsQKSt
UlBWiAfFsNu8GHBzbb9P5W3/0xdKArPWZ3lns+TReGswLAoxH2GVGwlqXqVrLULf6iXHA7KCKU/t
F9DVwGabrfsULbbYPby6JwBjnWntUPYTrA1kNlDZWoYoy/ok9clfbJqh6jjukuLYKe/9fyjaN9q+
Fv+nPIhT1gzQbIza9QwCjG3ohRniYtyx9wG6SCOGidSBLMNVKiur36uH0SopPJmwC4o57K+m/hsE
HPsnEC+2fNz0McxG132ID/doChDrjYY57JiMPPSQdf2mss/iK/230D3isZHjeRiquQTuB3b+0ode
hX3VCHjWL9C0cDDHmzweVMPKMT0KVyNXV3xhxlcRJfbEf8l9zxgUFXQXV2/lEy7YelaUrlW9yp28
PJzR2JSqLzVI4J9yZvQHW9eaLdivjcOozq9fkR9dOzje2e+HClcBXqhEZJ+E4H/bwd8tbSVT8OJT
mFF+WHVAmnNPV9rD/KjSrzG3FvPMt1CZRxqatheIpwBKuLSVcCY1zaleoxqTsoHZY5lpLwBtl7au
Wp1cltVJG/kDdztPqLcsgnRQLI187JBMXwW25lA0h/DClf5q95KF/5sNI9LiEbic/Yjw+kY39/GA
5Ja3HIydoqmhIcK2pIca3o6waV3PsC3v5MHluUp+ydkeccB7TRN5BhRpYUN+B3boBcuTWKeeAD9b
Xw4YRwCYmgIWE+opJDLOqJ7oCLqW3qmSoEMrjx1MjyL/cCtK6CrHwZEmjTv3YePm47P349Xs9tI9
JsJeiPRiZE7XEkQkVOLJVEN1U4fxowtamByIsQq8zKg5aPHVo9FuQMxMLWTADU5n1vpTK/Ws3scp
SJsDOz8Mv4Q186BR9TbNWS36INi0gxGByLrrWXcGGU1VlE3tZtR0DuTCgoK0oTjexS82pJC7xSZP
TrZkq4chV73KFW4BZyL04SWFyaYcBhSZ/Ic/ELNIeH9K8RzX2+0xXbiK9nc5zr8iBypj8jRrkVA0
Gh2fpBR6h5KkKxbZNPetw1s/zxgYhe95fVX+G1EwHuHVd9V+Z8rQigHkRR8I/ctn2OrOpMsDCVPm
++VJniHm1BQjAmi/hXhdS5hzO/8mmchL2o0PHlZ29bbZQp+PKhVwOFw3mtmHw/K5dzwRzukmNKZ9
18lO1yZ0UqYMgxVV4DeklbkU7s6ZvVEcWV5k5QmyeBvfmI9TR6557hra07Ddv4soNs11Q0z0AbsU
aNlYrmRcyTtq2lQat9cMj02C7Ab6KIP260JIRdDKm9s9UiYTBbXRHSvVGU45MF3peKyyCWt5bsyh
KYSfH89hfTDUXelmpGY9GYku3eXbuK+d5YlvqkW9FLGkEvjXz8UrFKu/APE4zCMZyavGOmJhSAZK
FV6Z4lg3XTc508M7zyPBm7d0rCL4Xq3tDBaeYOwfSghQPRA8br/gZQmhGEbHas6hPSBDN9hTUAqQ
IpIRXyv4z7a0dNDY5LfagfvIhIgkXEfURXRlRq1Bu/1roHMn+2lVKcKtqi+58RXp2RLHIlzhD+6q
wClZfK5O0ZgawSCZPKvIcy6GhKt0CsnUbbj9U0zFD4SRwP+BaOSW5LHHOXweP5cgfSOovn8mJQPD
kuBPEpMqx+UZLPWJMURbwTdaxTxGOjG//DCtY3ul2SmZ0l6xaxqya4dY5ii77dK4OiPiqK4zWc5a
V2TtL2/SGkgU/2GE90hhXqAruF8rpMpXXtJKAPrhCVML+VqHnQMuuZvWSgo9PaVub5lklQgPZkaR
SgCMJUxeY2xcsA8bGOqSNga2YiqpTtcl+RR9VzRotvNwrC9nOxqR8RwgZqYqzvYYR5dWnAYtJHdn
MEmQPWu2jb4nwj0lCi9j+m2fYglgaOYG1CCAyop2zWbSK38KttSw3GohoMxVZ+s82SAVqyvccsm3
HAD6rG4xxK6MxvfQrLbRItJrNi/fNPGh6h4T8yo0HvJWsEyqjamIAt1V//m/8KlxyYrxA/N59TT6
kpQL02uKdC+8vDpObUNyFm8tx/b2kUxMqcjrfUwuOfCIRHNF+ONky+LS9M7KTT42BQSH09n3DmzD
XC0ScJIFNU950NnUV1SnaBeaFTUZz5lCmDbp1/BmlJLJcap3ehRg15C88u2QNc+JrGEPh5I6el0I
mLofC27oTwlW9hSafeNKmMAyL1W+jsX5Ku4eCUl9XtDykeJPvkPJ8N5/goCy4i2mYqvrOP+ilS/P
iVgwGJUp63r0Cl2ShrB4ju/M2YrwQxloppP4NBMxT/H5C0pV40ziIEy711H4rmFe6XlFLuMtvuVN
NN0xgNapj2GWWEr5TdM7djL+Bd1q/f6CP8z8W2PbQHCG0Hu8iPGxGi8IvFSTug+yeO0NBzkFpjI6
jO7VS27iQN8BJHZNwFgPzP2nR0Ru2tRJ3kYVrE3XinHkTQ6jh2/8HhIdP9Y0ymZJTQStfyP/dhWB
H+I0uAU27X9hoiur1M35wcCeqb9FNh2ruJXTR4gQrI0rwlKdkzKUIFKw66+hga4TenQGizge0uiB
e0vN16bQc1O6TkxZNiZ9k4kpWDTdnS6cHcpjHW9aEL1QGeCztZzefzmzytGIpYKB/U2uEK4+9Fxw
1cqRd7WnmFD0T8nvoAs9XjNw59CLXxb05zNCyeAnH8cC04rryr0oLMBsewnd54x7BnuYD6RwU0qM
Fg4ixP1X3kWSB0UpomlqqIUUjeMHc94yHGouN0xwwt6qqlQkDPlwhlNuE8RydXNYLEUcbTEIqVqp
2K52Kmb/aw8EIJDNbddFshG4gZ8oPsvvAYb18HYzH9bTZ102aD0qO9wG+qb1cQpNVP+ZkP/dqmWJ
h4RyvSIXrlIH+zmb5ZcuJ1vLxyYA67WAOgK6OxqwQZSVxyq6+MTmZDRND+1Bfvcci1tCxPxXHWZR
igKVGtJCKY6ZI/WyikH8KVkpfwuQpwMJ3+7MUEAHvHKcA/QwkImBCmoRIs+3gYv8LM4iA0KionY4
kt6EOorvj4z4+JfUCqmsY08Ec7yCZTXNhAlHtL62HxCCKA40W07OcadyP+fniJ9g1Tl0nAEEk6ir
dbHK6ogwcUZ+RYk1aQOa86otuX5woUakjuFzMLG2ddt9dfPz1+6v7Q9nrtPmNQm/5ML0Nk8JqSTL
Udbmez3AxyAMxRXeaGRpl40HvA/+eu/JcsCov3br2b3bKJOP16HLDBKKP24k2Ecw2rS9vm2hdpKG
X856ikUYMdf8NTGOag4Msj7sRqm7+EJerthg+QiP3x17v6B4Tq93AoaPpsYYjDVfqaUV4o7Hx4UR
AQ0FSiYUdpL+5r8j9csyIHOWr4R9SR9Xn9LhjnZfgKDs2QW5U+4gO1xWfkYXGptQ3hPjsKI2mhVT
VS2xcZ8OGJz/sNpZ3ieyz3bttfpSrFqYmGsnwsNnRVNxAt6A6fzHeVFnWQOvfdMjhDxOaT6pqCdv
LPTKQgkCIjZRu/CaOoZlW2Z8yqOqsJUteHokWNvYTrMmsVxhdacsqmnkRd06WARDV3nebuzR80+1
wvyOTMMIyDX8deFljwflX8QtzssK40hHCuwtbc8IkVjX4UmDxDKCAqS9svecLj8QMb7NBRb4ORcb
Hq91WSoU6TYBBZUcAWdSqxb7Ykbd20MtA9Tp96fixCmgHhncOh4LkFSrdJ1RYmo8xz83ys/rT67m
b0tHZRdxrDKDK6h1Q22TfqgCyIYJl1leTO7O0pXwWkHBamQrkLSlYf2yv+foKg8vUwWtS6sVZ0fs
Hy1hRN0alGiEt4gJ/kRE5O8fY3anjYjIC3d+EgTilpEspUEJxqMZJRcMMA1KUEX5HPQph6hGoMs+
xqkLUyFxvCSlaA8awmFGzMebHpQGPO5Ts3dbusBlUosQ52YTdrQBYkD26ZinI2KOE3wo9fV0i7xH
yCJWYUPYRhIg8FjzrfKj59OAW8YOc/xYqzB+UitAR475r6apewYLiuyUs7k18xl3F7Mw2jXjgqY0
+bcnn4JNb5i17ojo8lrHxrP2z+PNc+8aapWBJfNn8LFhLsn/FtNpx9jGder6ca6ZiJNMQ+RqLP9/
N0FV70Y3uMU0ZIdGRM+SB9mtqdiMiBzOTH49mtOtulq+mfzIkBM357DlvSi5Umb2vGKmitO9LMGF
hh28xThxnKnS5VTEu5LhDi4rB7id2q84ZDEqEkHc+U23Z3NnnvwuclGEgCE70dfjeRW19MifVYMY
7xAItqnBMaG6etU8zB8RPn3cJKPL0VqaFLCemxYRsmLpobYIlcjoYtBhqD4j7f8dVDZIdLFhch+K
twE2/GMxs35Zd9Wl2rdG+3GQhYUGyzZZGVNs+wWkyyPW7Q8aTuCfdOSjpbuz7vds4hC0O7Oc9hTA
ROhDud5HoNNBnUJdL7mkv27LQbpi9Vhi87JgQKHP8QCPK6bHqEIUxm173sR8r+Ckspy4qceulAtc
47v+HJBhcVJdXAZOi88FulRDsN8UMF938LHXF0X4Pji35EkmU5FDW0H0Nm6JHThgNwAZvgzm+Jn8
DHlx9xtVTgXSNlAJRQd09dia+Fdq2oQR3heLK/6XV7/tiNDrBJ2WI/evBAb0HaakJ9ppAwXLrs/K
XO9e+aaB2FDhWELILg7qDwKnhbzEamBKSJXvYdthfhSXsd6Nrtknf/niPNZxwxJqZ0F/WzLJgaHG
oBt1xZi9kHR9kFqRrcwqgHe04loRykSE2qxL5mpBxKxwr+dWIMJafvHhUIoUBDchVsHo/NmSKmL1
9PyPUhB6DzFD5OEQJ++pBctdUBGrPUayhGsyvdjTcJsHW9fyI4AX5egR2vkTG0XULgLIXqlsPOGf
vj48Ab63rgMZrjVXBINGGxn5d073/go+CXl2x35IwQ8TLzGdEH24spUbk0FE7BOeeQHdyO7enXNH
ccF+6QT4Z51Cnr802rQ1kaWxPdO2o/92waQyNUL4rM57FPaQcOlUuyePY2TYrRP/79ADnxEkDaed
35gChdoOZewT1pbeHFoF5zhvvklDFJ5hUrQCg1wl6+7/+nkdJO85nP2OcTkP5Ir/rCF+CSchmMVb
oxAV9LiDAc4fH/pgrAPa3Xd/IdwtjaWeTgtkIKpCSnHmuNpvrGrecamYIc4eMcrT+MOMptKjLgAM
rv6dJCYw3xPi66mfp1xEuKuvB8HZW1zt0kJHUqbZfT6Z6ays9RY0N9SsDpjwLEk6//vqCoFOdclD
Syu5jlYRN2cVPStReHhinM8PCBmywRfYLEndynHv78SM4rdQoeXN3iU1oyMCzFUJV8NS60x2aNiP
8vi/S2QHLXufibq7Nk/UHDmVVSz2+0eASEOZkeeL/y9jZDIJLve2OD6hpaZ/V0Y7KgFAFqpijgXD
OE6VAF7LXP9qpyq5Dnfxd+oOwAfbPY+n86t2FrNugp9ilIOHsod6O9MzzSSJ5NjG/NVaWgrxOSAZ
4BWWQ4ENMKNSI6lTsXqujZCFC9FlZbpBP8CxEMSHbbICQcrnRI0ziBeWDqr+gNfRL5YVzaRSs9T8
eqEthtNO3CArAuksTRcPCjWbcNfIuxMEfpWD2FrV8nyGkPGX7NjnyPo/EB5Py7nNQPAQ0aKkx2Ym
AvHE1jZDSX3nk9c2Siv9wHjZt9KNzn05NtASF+16C0QfIz7uvjLClUAwq4EHUAJz/q4T7xZekm72
Pq7+s9416ey9++slyFqOTIO+V5RhAMg3t3aPHaViqWNnPSxSNDNnlVnZWCT1q/Yhe+k3aPcEeROn
DAhfBjOCQNW1CBQkJjbAaRw3dOn0i4BkOSqLoiZDxzlmrJjYvT1KI/XhcR7WpnMIUS0NM+V0sdHl
zXXCSOtR56sHCjzHGfLNE/XNJjvvnSEdWMHv2KPye4FYnsy8ozaoP0tr1jQH+A3haWqKy8yRb0SW
K2zU2egvnpzzwDkbK3YO9i+Bns09GcVgQMgZDXF2MnsycuXr7pBqRVMvX0TR2qTLadeNKf24zKvC
Ly2BEJkXritA/k7nlb6Fpe09Jh26RGn4vRqR35Wpa6NKKrnmuYuHtnQCFpEyikPfaOBCYIi7dlTE
cXSUoePWrCJOQbrYwVS27Sgsx/N27Hdu/RQXQxGGbnobul0QLh/20v5AnxiH/dE2wh61JqQhnJkP
gSWgHqhNsZzE0d7epEzCEVlPh5O+YEagJF99AALlab7OgODlGRlDQd7o3W6YulnXszdiIMlm1PZi
W0ZK9zoTNFhyVUc8WNZljN8/rNCxte9MM/Zb4GzVFgH6MJ+Ptvyl9RVJ+PCNo4TW71mF+LpLd10i
Te0hfPLtllPaHrCGUtvHXZ26thmof4za8CN8cZop6PFl9vGDEJB7JbaigZCLSmbTvyCfSrutR8a/
pafteiUIefECR9LHLdGmUmTNJhkcwlGgRRXm2iNozBzPS4S9o6+7b8sYDsVpNlZYHUAIKUJqgK1L
Z0n2EPtn7dqJRysU6RLi0K88CzS8XYKUCxHPZGFxpijsanDAMmOdJTcR76cg+AkTQkIV0869kNyB
1NXq40LRxl36C1QWSKvrm2JgYPo8VltD+/UDCb5lRJqSiiVR/5px7jWbqPpHjzEoosNszpJ03pnS
o3nYPqpfhYdDKHhd2xWM9h3uMn2rk1Y7L/j+uivvfUOmqiAZAoWThGzTsw8i4PAyKF/S3GrY3kMI
Z7CyRuQiF6OQuzsggB0EDf+sdvHQ58F8QcUNK4EuPlkBhU7/KDBou1mkB52282O+wC/agfvZBymU
W+lfqHzN6q/CCKHubXyJH3NaDXtMw89UOu1mtLfMLFTCyTtiv231+m3Y644C2bvXcQ49rt6cDv5I
O+hW5NXLxLXOKHkcbDK8SJXt3MTvyeG82IF5hVGk94FtwHRcI5hm+ywYmvyy7gQkuKJKSEOyH9Qh
UV7+1BZD4MLtIrd8lMzUJr4da0J1/RKu8udlb0Vu+F9SbW0/N8UkTYWutrMfP359eC+6BYpSNWmv
n6xRT6K0Nx5LOje1upY/LNYA8sNU0cYxpGcu6WHJumueyC+Hzrppl+X42sczlFyfM6k6Qlx3ZS1K
VI8QCYpJ7d4N1j9WH8LPwVyYhk7lENghQ2wHhWCFc5417FkU4Mjn7B3m4PK+dhUGuA4fkGvD33lh
KxEI5lOz2cPDF4mBLpNksWO1AAJ+kBCwJkcNJVSuu3UVp5Cd2NezWgSoVHyITJo3uBaaIGXwBtI7
ORreuHyF0CnQZlk87RqQI3z86E4uauHQP6anFyLLCKW9Qu9T5Vt4R40sL2UwyXhCWbSb4uq2YT7B
Q/jC8gg5hWPSDwaepRYJf9sKE+JOIMWK4eMjGDD4OLIv0RKPk05XlhlnexbXepoWra77hOYcUDv6
Jiotrn7Ay40T8njtdrokPKrawUgKzewVYUEcgoRb7n+ROugSI2P22m7NqF5KgkYJWmRF6RAGX6UR
ejYYp7VJ00rlpW6fmFqffSGZBqZhaGHht/MnYxwPqMbZaqR64iI9meEO/FAiKc2mx7WTvQq2z/zL
sVpflfxD+5XjCKVZg1jS7RzxmOl1NbrdC1hfPIlH2MDlyc1hMTsesMGMZHVmUHd6HuIY1wBsUy89
aVXDbik/JioMXBdkdsoBXXJmu6+wEcbhFBi3eCQCPXpHEJLnptlfhq5Lixd+r820JeaUlbPDGRyI
bG8CTgwfnnY8sgiYOVJf63k3plVV6DzoERIhIrUnOG4Cn5QG1GjcJ+/snACBom7XqdA0XFyHXcaM
cVhaezh9yAqKT2yaqDMXt5kyQTLvfpqfsxeryNVeXBHxtSlXfs4Zu+a5n5pqEW7/eL/EdaPOAqto
MxSpnMOg9jYqLNCg/llJz/2GBdSBIFyCS+aFHgHUX+RoQwTB59xQbwdRFyZUp6NhDnQVmRQsNS/3
LYk8jYD+BQ2PynFgIEsvx53a9Y5W03x6xfotSF45viF6Sa9RawLprbU1ZuzGx5VHmo6eULoejvZP
b0XAf5CBi1bHxQqokJSDWk/SFgrf65m4na3KtrILANpYvjoxkzPGAZtZqnZKFCwYiF3hUPl9h/Vr
Kc8J3xIw8afjxacL2/RiKpBCehY/gjC/FInRF6kv/79KwxnkbxX8p2Mxwnk1Rs/SUY1eQgOt54MR
4O0Mv/AqoyNalAPc/xz2ik+hdTPo2dCrH2YQ5ntBxO+H+wz5LfecGCoCUh3iL0e+FjPGcD1H65TI
uBznymEj1HwYmMCGR7H+/6utpS8QjPAuE3yFgFFhj1dmKyMa1pocaorgXNqzw1OAoFbMRvFqawwx
eKxLJ8miAQHSecfHWzvcHDKczb6///7ImwOF+QOzH9Kp3NqPgTGQ02g76Vk+l0tt9x8KQfo4IE5Q
WoNWAIBXj0XLH43JGct8opMKnKzV4QYSaNXOn6w5AdbBN9cNlnQDSCLeLI8SeJGWsVnUPrz3tk0g
PfxoJ5NCqHpSudKFXEDFFpimqyEaOcZTHj1KTks5xilMkRQ2HgSvOQ/6vVh7dR6FcZekFn/OpNEP
oABml5MR+ZGozhQtUPyVKYM4mrOLCB4Z2BdQkmyW39lmBNdju+KkkULH37cEpWIx4T+sbJTYTuUZ
luUcufOTZHG8qEua1CEi1I8ZJAGLhuxtXcIDPng6D0sd9SkHJGsjhlGu4wbdMy8lPLyAyna6+c0j
4qBjHYJ18FID4a8Jo191pb8vf67vDBMT43AUqsxoicLIZplaHB0ggRzqByj6EzlLYmDR+lUA2iud
p4qeL1FQZCHrotV1zmIrj22LMpmrkKvA1f0Zj+kYu4ODAzS0IWO++LKfpyaKUQoluejJxdPJXyjC
lefwOKAWzZ7DmGdjrXCNAlQDoEQuBfZgtqcaL7ULl8pJW1JsIlp3zvWh6IK4OyZYO+/UzOz1a2oT
qluAqNqBZahbAxc7IEjMP6DHT6yOqHzoy6I4B5WG9rmJAoOVo+pXZtRf9TtTkoyGjQrjha3W2beE
EpcPyQl9eWy928pc0BCOIoqYSiWSYkM3EwhJvmoneajnu9lReAN6I4h5vwxbXJXgZfiGtE/W7v+K
yB2JkQ+nrCHnLMXdzgNHX51uW0EC/WuxgT7LzXNFFAo8UWqb1yHpmIuTPdIZm7xt+wC5gYQUwBMZ
dNKjiuqnPkT/rNW0eKhohhzC1hBnoO7TGAmYEqCBSTWQwNSt9Ag4TroSNb2u2ZasOjtX8qSt1Q4X
BXkA/LSHVP3pympZMwyOlTgEcAyJrGrr0S+yGdpfUnI9TFO2rQan+rKodyAGw8Xkakc+pqJlpEWw
MT4kuDmJvj/kBUMZef+OAPTrDNe9btdVGWfRoTLo1mZIKFda6v8iqFY25xDAKFlQmBMGSuduZ3t4
zhpTxEfS0jKxW8AqCaigvhC2HkvgOKSZjvaTJD+1BzBYMavHvLmbVnJd0dyV1OfbpNcE/i+V1F2d
o7x2Zs6+ZVnEikXgTfve05IJBFdbsZqffR3Gg2xPh8OOk7CvqPYNBkv++DD4ZOQqP2jmgyixd7b/
ooTnY4XbOh5HG4cYfi1bx03d1F7oH4NJWSOh9mgZZKeuqPYj6MavQ/QufjdQ1uNFNqtJ8md4Ztgr
hcN4gZE+7mNmO6OW88FLmJc4R2OoyACS93mrfOzf/9GJnAZERn+DoMRR6Xpya2DaJlhb5qiI2YTM
8Ep/oBmEpzxVOnmXjf1NkensST/+6iDPUfMUdALmW8doeYdaKgkhwu7OgQz/E76/YmLX3pZve8xX
mQs1WCk5VndTOyAl8pjlAOtSoaSGcq0q8y/7/8/Db4AHrKw6+d7dgR4crYuwewW7sPbvBfiue+/h
zL3JY5Yr6ydVjkC67k6zUMlj0chZp3QPNTXU8R/FviHR3/S6Bg0ec5ldBt3kDeURrbJ1m/i5vMrw
p57gTZHhH3BMgXQZi6IBfgRSuhYGGQsPOQSNdAff+hRqYoEkAlZl8y0fzoYASs6E2u8VdeuIzClj
lzJYTjYyFmKXCxozA80BPWuQHd41Hrqqv65gmMwCdiP8FxDuHwW7h41jKJ5J9L/GVTJd/UTObfEu
JvT0edVeapMm4umOoPnHjmQIU5JwjHzsDjglX92m5VcoTm0NQCgHuI1XORv/0ZsFS/z8KfwzUpaq
dcSkbU/6r6qKGTqayxCZBLDql9Oh3JGVYYgslOvKirqY9e9QJKWbCRJh3r7RDqBYsiQKu4A8eOOE
zM+S0PzQBcUTaLm1bgQcciZb7pJQlrWHZJFlTUxOfoaOfgnLRMRLsdtBD1ss85PAUwdGyBLTgqbc
LySxkJXl6KUJti8oVDk1RvaUSqR0F++vY+ScZUWCCu9NQ8ZaAuv1b3Ai/xEfi2h+RTfGLvL0P3s2
zZr4J9lYqfylZ6kzLFjsNf7Y4klnuubJPafp+e8YyU0cQkO0euTaQVVO57brArOfXilAdnS+9nRP
ICx17K5a9eLtd/NkoVkDQfCP3j/hqkju1UgDvMP+GtYwKiNvIe7o4ZKt5Lgd+NM8SNSu5kz7eGB5
Q0Rrwlvdt4H7seGXPhsiAVno186Fe05ecuo3U+ziQBVAj/SCAVZACe/E7d4p9Y7rEVtyVM7AS521
zwRH7h+10cwb8IWGY0qKs+fwOK1PFvmOrK3g9DZnR1cjDC7+fASv9txZSiGztRT8DMifhBHeCTuv
osLdVZmD+MdHUeCDwoDhDUOBAVwYlKNrieBRX+ESRigAtM35B/Bt3SppWS24Msnarh5u2Dt1gltJ
djF/bggbRx+PuC1FlTI6OnYPRYTGYRMvoSU1LTAt9KFAsq2HefyM6XrwZ0cB8bKWkaDw/TouPvbJ
HBy1t/kwXWmJLtpztiIeyces+Pw36dv1ieYfDNNtmGNvAJpUOUsXU7DXfYBE0AP/VHerLFYSmUt6
/DnMaTyMwiMUj3mLjfgIcsJHwM09IxSjx+4y9UYiRN3f4JxgoLb4s/Tq4+RTpZuq52I0Pi2WV0+e
WMjhyMS8ZPoCwZknTtwoYsbwMqW+VjNGcJUCkWbZrCUr1etfIbkVsz0nI8c3oLvSzJTxhsEmGDtu
s+5jtrQ4VtreKTEJOQEmOkYW9cJRGA8FJsTIHjQe9r+f4/H8u14NTCUNBF91mPOg+W9cTBtAp69V
5yY0J75bQzTfn8kIviP9TPwAY4CiBoZ+vk5qcv1g90BWNm9OvO/3FyG9dTCybRq7nQbxrgDjwUnx
hNhJgwtq5/O3dU8D9yU58hs20JhoD7At6FFNEZyzNVHOEad9rDDEp24iAsISgDkZVIra5Rgo+Gnh
+vlitMKte5QN9nSjqdro7eZEzqUUzYUyTgXQHbCVC0G14cnYRCa8I+rMg4mxWFXEhtqUCKGxzcFL
2PINyzm6goznvycJgfk0bRJbgguC4tCfnUXUbJHMzv55FcSAR+uokmNSMnkW2bVeyu7u1JRqiJz3
yA2UwXFiskqkZZyBtk0w28MwZNsvm36hIil5LjIp1TyPVH7zudH/CSdI4TIir0JkCz+oSqdz5VM+
019yYw7BBszNObr01ajbAmUbBtfXkEMxOXkTNiPMR+ROuSJJHMANtTFVBEfRGCCuQ0znFqTcblTL
LlaZzMkSTxtGnLl8mGdVb2XjZcoBGeIy+AsbD/m1O4ztjpMXXX8gMTGw327lskOjVq27eylPD5eL
v3e7nRZ9amzWCeqAbSzXODcvjHOroKb+1GcVtriS2Rk8mzxhNCEr8G1+L4ZGBCW/2DIMVTobIFLO
se2/qGyOWI04FREopiR3p8yPLxZi739To5gsfQL6PsPsqv+V4ip2ozadIJ2ZzEnMxOtbLFYVHJpz
8j/mEygWHam5xuG4fMDtOqMUu7/ap5kHFoBkfz81G3yEZ+NpbqgjJVZPxHbX07ZnAxZLgnprdV/i
8n8YSQZVzyuP6ByY42T51pHjAAwyxFavGxAN2hUAp1eM6a6nG4nilNizwz/r/vxijXaYeaoZyR7C
cHmfwgfZ3V87JSlz/B4e5aPA+u4E6or9Lc9Qt4Ga4gyDEtxBHpzn5u6NotBoBAIEaJUlMdGaZMAa
WsnSGG+8XiqcssjnPSr7jDlU+ARE+g7Ode1OeX032lWeeyGyxMirzXV+RreaxfeA+JAsl8D5CnQg
BxaMhJ5HqLYQyyRDHnAQlKMYp7gq+qsbRtkL/qHRCPxcIfXkdGaOF4uMw4GvDnPCPY1eyS8q8iuP
65lPrXmwwxXlwR04EC/pLdJcvvBA/RykckIfoDhVUUHvw8aU7jPoGSV3Q+9L7awOAd3Z5M7vSOwd
e37+WuD97mXls8aqT/UHl2vLPudVoiv0wuUFNV+xHpWGFrBGDiLAesYJg0ZIfB7FjLFeknO3sPWo
LagPF1f86OkVFbklvMynCVDfc94l7guq5Q71Agj7NPY5ea5005pUZlImy7GbL2QArsezju19QyXS
0S2DJMx5WEgLLbO/rX3kO5UgqRLmtU4jKo+6TJBgsK0QPOdR/bEyZk6YG6MP44yUplry74091D5O
3W9CBKmOhTLla4kyW6rtmh2tbp85Gwow7VRPciPL1Tz7JS2EvILa6rD1CyEyYVWOVeeGXfGCAVJ8
1jsNZhQj9N4G9Y+lYgxHvgdJkjZXKM1aXpq7PeyMxuWcn59I0XAEJbTG+TKu0Tq0lDw+eZCUjiM9
sTioPS2lGua/RfoXQX13FvCnsKuqXHXApnjY4mXHHLZSIZ/4W2Q31HfF6nMOPhcrT3TTUifnum/y
moXnUdhdCqXH7I9uuy2zkHJLra4MJdYxCQg0xzXX9+dRuyU4vzX2qemFpDmutgafRGpeiWvKCzY7
H+3vX5Cn75YX6zmGKN7UiHZm8aKlWZdKMnzXF3mNPn8orjq5JLWgTx0eQsbsnpp3ZJYZSQBojZIK
qpMxXrn6JZhcxqeYIP2otG893b5FcrFm0RaGnaGoLuQ9tvtuabu6uL//V6oQwegTwCdgsh1IPWr8
dRhyo23ZyknwFKgRqA/oj6mJE3n6ZzhxTElyY74kegZ1xE/RQU9L7G3m6qWkyImaJSwAPNyFV4ue
rVPYTsi48yq/LfFafcXJtzlxRIjC2b/eV/TQcSkAZ010WgsNO9VZbN9AxDW4f3RjpQ5cvqtbg22+
J7neHfqG3GfCMP3EMbECEvk2I4og8bAfcg1bMgPTBqcXj9DNsvokIW9BTzNVpPFdJAqp7dVQK0wQ
+ZHiTNOoMcOv6H/L6jiQGZkABi7LU9jeqjHehvG8wReWqCknwPdwkC7jOwMa0GUFk58UQZZcXYpE
B2c9eTTi+jHV9VVLKCVsJgKQwWBudzC732uGAiWEn9vlFGXg5khbgTMfCkGI9UXEmk19ZKrk/nuL
T2/sy7qK9ldxYpmepXgQmSVNzkvZIQyGl6QgEcCCv0rlx3+XjUsY5mSt2QRUiaw7T5dCuXJ1N0zS
D3zTcMBFEPOh8ARDUDqsuAywczPK4ZV9ZVjrZ7NpQytXBpyGqqVMT+MMhZus5hYMmSH8cDaeCFak
og7mqREl6e/Noygi7WgE1AEsjCIQMiBmzDiLp3JrCoViC4pIgy6sqmyWKcG5ZzNiGsBObd6DNKus
yb0QEzWipHZiXAwjz4Iv4vtJArjmVXx+ZkNg7JnsI+X8u9Se15u8m0t2MeiWtmLcpwyyoQGF1KUN
2nD0A12hr2H2sVnbUTH5k+Y6o97YCI5/p8237hFe3KQFBMjrQLyq2z8NC+fnECWN0y/s68NgV4s5
hNnxlunLF41BmsyPfRyc81oD+sBEZSGqpO0CUgqv9/wZSSHHFo4Im8lqmNKPODix/dsqGG5HF0AE
VKjuTWq8quHSWl1V2BjYsRHLQZaGy1CrfgWPIjQnVIJnBsqFyLsZLq4piZ9VCQGG0eFtffm0t1Y9
27VAcy6XxNIw2G1ryF56vDO0b5oz+2h6ySVaO0NTHaupmk57sxGea0Jb85Df8Sb6W9sKvG9+aKdV
34qMHmbnJ4sSR4h5b6qVK6ovuTcCZyWrcGiTooBA4CCzUa/RapyW5Tg2mr6uV6cIfkxnlOiGZ8lE
dymeBu44XAwNpEyX3AwxdiHVtzt0xK7HI5dicRZu2C9fH7ufJcaBDY6p6nt7G8N0kz1k1GOsyqHi
hQ8qmLvuCe9CekwpRRO0jGjxszrCeJ03fXOmlE/x2hezxO5PU6dryMHANG/C3sS75KEp8OJvhve5
oLUAzu7T8+i3sAhZlHzpZKQFZw0UH78LZ7ws+6AZ/Jot0Qg0dv7ySYF3PjAYl7th5OQC+2PFkCkt
VqH+ASqQJqokb10zJSEwCFeCvZjCmvy8qfsXNOafXAPWDm5QuSeAydfF/M9s8hsR2CKVp7EkVhRi
T33d0p+TNws1Il8jZXfhQHVcld99YY13T02XusOrB+wLIPCfU07oS0R+w3aliH72G3WiStAu9bFp
Yv/wcrSZn7GhOwQbZF6CmsVtfthYtLh0YLHk4tkYDEqqDt8HOXEagmbdRZLmFiSYqtQtE5pLdb1c
D+p4QvEvuaNiEYR1Qcx9SKt4Tt/aDKPH+bYfnfZ0sTh/3zWumqu4PylymHEKpbvXwRfsRhxp3/KG
bxTZoiofMGDg17u7I8xGpbW7rm4G88B+KHHjslNr/9fHsWdmgbqxTsd9t366Q74F6z2RHoefkXMV
NWAVm3HTbK9oOFWQlsIra0JgQY8kk5n6gmSNOvrtacykeYl5DZfwJ4UrBImeS/E/FQ9PoanZW6QU
U1rtcTH4v5bKkzkXvkmQj+8u4XVQipo7vO2Sx7m+e4quoTJeQVZ+M/8+jg9dVd3W3D4TlGXiDchE
+rxXiTi4g5sz2Io6wGOTZui+ukZPc/Ov2Jd7I8qye/jxrdXkwgTw+bk8hqtUlRJSTLMl9rvZSpnC
gHH+no1A3ggM22LVALQiWvdcayiRJLH4lG646uqRC2/i782sEHeY8LaZVjKt1w3KgTVSlgVxkf7W
ip0oCJ64fOWwt6LAuAHoQNM+y2jw8s5IB2mV5B3rvcCl3hdGeBlJzOy3mXWAdCNQBZfJ67FdSHer
+NSY/wYqgweShLBFD4qqkdh1VtMYRQHegnExj0MEiH7HlB/fZl0oWgsXUvbz03ZgdpsO2pjqaH3B
CuYIqPAiLzbIDqh9WbrBbRVQAbly6lq2LqRAgZcoI1KyROuMIFtJK6FcqGpTE05jh5xUhURCGXEF
RFnVM5brCa8xGbmeWlI3e/bIEYxbsYg4YFs2qoLp02m4nyveKsBBW/OR7IQWNUAF/ws2/e4Sk8z/
rF9hLXey1pCLGG2Me8gAxoZDX2oF+tTECapC0uoJPk0fZMK1qvju6DfQc2lyVHM1n4CUh1olrSTy
Tm41SnTK7JW41QOKsjMoN7fU7quJu+y85ewrrYuRWJc1ICufOqCF2wqHMpag1+ouhY+eGEc1vfT2
qu1h+bbB/5LB0YJwZ/kZ0jcvNf2ROgKz5BioE2BaROypWb7BVGXbG5rT7lAhBmTp7UO3Hg18jmff
oSRDCkympW6h/5ExJVZPb2ptacnXkpDFTM9XaeO+BSamV15jx4ZUNbAxEnQdijN62nEtuhIVTDXk
+jGwNMvaAUybxb4R+lRGojvr/QAOzhujCA2M3ch9DqC6C70+Mrw2skvCv8eVq+XcpySGy1myi40D
MwqIXCaMqcjveRYt/DFV3J8qskjDTsuSlPwjm9yXdPkNsBCRskoE5AE4RPYt+4ou4e2bhDZF3X7v
zR1eYaR/jxOhSse4E0nwkcIi9fpy+5LwmVYJcabvn3w9B3GM8JaszGvULehWxnwV4WmgZ+AQk+RD
h/DHn4uFsKdszE9MsFYbPNwCkAqfPnaIrlaIf0/+XNBSzLUXwQ44tkeiIoTPys6l+KTNjcXUdo0I
VHMSXpq9AJPdXGecM/avRdpZpxShq+FR9AaVu5UVlTQqLLf8jkKp5NxNb8DYB2QySTtzdwmJX2Fu
7P1wPEX0REUOvD6r4Bq7/3mnLFmgX5wrq5Yr4hBPkIhE0kgYw7vuSn6yQZ6/2ML3DgiNJZRqar7o
IA6h1jmjLz8WxEg51Hrt4r5Me9AN8Pu7a7E6DFX8QRGnughbO1YGgKag7b398j7L1Fn2hkefY1FV
mieipD69L4dalOrXBK8UAVXXVrcjmFbwX2oEf2XBCoWClmmBDU6QEUY/wwE7luArUjAotFCZQdJr
NocGDCHp0G/IKr1iI2kM7dA74YtoColXu8o8ekKfVyL65SaM+7yrllhoHddsqoLT0ROpUfsMmdaY
g4WIhS27rpiugCVFH/NyJBYGh6xEHZ+tpJ3VY1m3nvWp1/NTbIuZdS3/VNN2cwdDJWD7wh0tKozb
e5ov6ZdJCf/RcZgdj/jetBKwzs85HewXWbUq4p1jNOtyveL8zNCIk5o9WED0Z9m5aKJ+W2eQQ343
pZ4x43icqdTCgWR6/JKDnK1LKMptZuOX+WcrTO0/quBFU4eRqd2YzwB5n1yDPlfwwCBTZtwEUn2p
G2G7Ugf6y8RjLB/R4pN0PqWXsKH7qWJrjOmPhaN+SuS06d/Jt4EYkR9H9lbyWtE1YSjzP89is0Mf
Ef2gTi9nuDRlhoz2mfLHJSutXts0H/GzKCJ3ZGxI6TxJlLzrGk8un0Yvqvzmb7weYivqL3o7CA7t
G8N6E3b4EBNgUFxtsmp1jV1a2xsjptSj+rlmUIvXUMhGCisbnkAbtt5Jk7NGxfetd3Hggl3lJ5VL
05c0gfMH9DJOQixf/p7+6lMjSi4+d9czXuKu4Fd4RURT3Be77Ivcc5coNeUazZGr7AJCFctUV5V6
+VqmCVf2rLTDxPvBlTA7XaO/2LOii87cIOQYFq+ztqKQSGASXpNxsPjj3/0GgPCIcQkeDQvamO+5
vct629tx+iYVAcIirQm7ZKt1RZR3BfVa4iWbwEzNR2KHcjWfUhbqU9GJ7vnpdaVScBifEJUCxdom
B4MNrCifokGc6pl/Zo2Kuhka8D0ou3EENFsC0o8uq6lwhKGFZGAPwtjGqObNZr9F5tJZUKLSldOa
oEPOw3gF21a/Jw8ikXtZo7bixgN1YMnLHOoafP9Wm55HsztBUlOjaDTXxGBD/LgZL6aGKJot+6Ft
s+j+nlBDraVeGF9tTNzVNxWWh0ekKTYfE8Ku0kjGkXGx5hkVxKyujoWNsjP5/9LtBSt/3gR5sgpE
lhu9crguWu4nf8IVUqQhClRgkUclBLEaEfjsBTRTMP4j1y/jyr62woWdlxFeQH0KhEYHdJHlb9QB
XCMm3num8obVP5GeFg18HVtfkn+Xn4BLgBmNmAsjRdrB7Xm4z73WY37WHUhW8EwqkQfxNCKbnPso
LxoSPuqDOen0HcLsNsslxnJHk9Ix8fWrmxCLNy7+etAKJmsllqte+K953iuIKglUKA3KinTdy6VY
T57f4NpWBWXt/RXfiH2sTpNnOYcYFB7DTIT5CZU0Q2Om3lwXsS27/ZmVk8t0Md+eeXtA5dEdQRq8
zIu2o+9cMW6rDrRUvZhpnAQfGNoN8sdvgyUOismhFeSktDWG6p+VN5Jf3GGQpbKlI9Tp3yimtbQp
jzG0bGNM9AW2p70Tdp+z9Uo7x2iG2ZClEilujP/i+E3NPz49dyJqpdB+epF185kcIz/Zof32HhFo
g6za/aGCGEh66TJrqjnwwfz7Yxksz7Qad+F7xt2bqyPc1rKL+ha6XQhXZh4qpQKjeOGIahGT692b
T//NEMVFVWv55sRjXXbdUF3w7+VtjCy69cigrnPLt8OYhdAds4H+9DopGwMSk2yqbVBJrKJDcIpt
m9QVJBbTI1gqf0fUY9Ginm3esUMzNCQWopQpBoGgm6bWe+SuSFvyslVTiMZLt0Bj6YgYo5zESUA2
wBG2TF2vuC2EABCtu29wZ1iKngEQ25yhfBe5nL9De7LHv3ATKEHEK9jjCxrlgmfH/1bXMsTvtfSK
bWRHyfZv8F48+HBqN46tKUegoh8ylSVxryViF4SDhokRINK53HZ/9unZQfdUxoEXs3s+iEKc5CZj
3ubmS8LTCNGosvVfTGSsA9hhjyfT/YIUZY0cS8nFyAbePKGvw4hf8EMno+ds+TV5x1S8KZjKqNZK
LFBk3L57gNHgatzTeJ9WPuDVL67aH831gxrpZ7JQ4ySoEBEgxgKm1iPMVWPGts5i2sI7mlAsbZ/z
9elW+C7JTV+W93lV2cOkgxS7EmGPS+XUOfmZIw2FpwY0QX0lhjlSO968wM8NE1gu4HbFQ1QXOx5L
k3G+d2LAVLsF/beAp0m2kmzoq24oWR6jA2MU7C+KhLzmhT1m35Bf066nyHbzGk3ESKRDWJW2wiiD
URCPLILPQhs4FRVN+Lg9fz7C69b9eUYYUHI/jSayvYAwqeSqvJY8uTxG6CS2RZ7EqiWhcXlOeXVd
gT8K2/ymMix41JSqscb1EfXcHmSwOxhRsu76/Yq5KgfVH2aChvIGj1e45h/P/95lMj+gNhorpZ9F
mgpjhvcF5vuKRg5EZaZ0iHE+eZOViq2ZoG0gRlFlKZEoW4Z+YVapOJ7ZPCQPyuu+jKRa8bCcXTwo
R5N9O0IKRQQqIxKbVGDH6AFv6YCl64wd4OtC20aVZpEM4Si+VmWLCLhaQXi7FV7KzfVcFh3BWTdq
NSD8VHdV57gjLL6X8wSdl2GFdV+fo4PBenwNRLIgkzXdj42jvjLcVGuqr+xBbcEIBIFAwCV33aLa
pjLgBzVCflyF2Gr6jlD8iLsxWVEKgaUL+lXvxzdz1+VTD0+zhxHScUIqkQbdGFa+W5lDSUBggbrK
P6a1ajS3LmlnurpLOsUGVOee5qpjwW4CgEbZ8D3Tgkoau+xZNEJ+w+ru2PGQaTBIyCOxH5foa4s9
0EQ9I/u/kFl/dIVaY0Kpsi9jsuUu6WBBx/1cOC5q3oxMfCnJdqAbwhiJLqnW1qub+S8EhZTcrLgw
NWnNVURkba4lkwDTfjWXmAx+pop0PlqkCcLN5xLp/SpN/6mSWXoybVoXUY0+ORtpbPWNHssfiH6k
KWqaKebEU9FazEJ2pZRnnmR8PTVlqW4Go9YOxVpcD46Q4ntde0/3Rr9iOlVq5JnAGlOvI9LtAsRP
Q8JRouJ7zND/rvWXRUap3LVjKrNp0jIpjvtHKxDpqIzt7fhOODcR0BUMPxMFqa7XXyWS1IcWbEj+
NIHnpVYNmnT1Hyely3wQvI+R+Pnre2Ktgo23SjKPy/jq6gOUQCjERYAhb6YC+nkUXaj6PFShY2NZ
0IAxcLHpLu1shH3wGrhPdXtDMRfVevWLrQ19rOKb6KWX9IWIwC2eHKRyshtssRmnp3vbzNbJoAYO
VMOJ8Ww/Mmf8+jzfkh7QZXt9fMRJOy5RSiioMRYYaRk/UkQlzsUAKOZxsPJQlsNvwz8Uy6aboAmb
wvD+00grhCBcydIjHT638ehb4C8VEZyBsqc4GuocAvmJLFhNtqV8x38QjRJ/wGShaW1V7+CTuBC/
R50LGdMgE6NzVpPgzFTb2To9z4Y6VvXIVhPIp+XWKbrPkfmpPYDescov/eeUvqC60QAwPl/EroSo
fKUJgZpazEC3SLAFTlU6qqIZSeaMvS+kv/xnDmjmva8HCK9ANgri0Z6IZ6iW5eQqn1lbv7ceyTns
WstEZogEFE5mq14Nss/WOLTQ9Cq/PapM8zRfRky8fIzeTov37yMaUJt660y722tfOCYaYumVB1b6
CZIY9N3St9uz4b+Nf4P1yupsvkKtVSkdiXSEqvvMSNvN76ys88bujL6lS8t+b0i83FOJhY4/J5mF
7211Xi7IZgiwD4y0owaVVvra5KKASSA3TtY7D1GneDZd1+HG+DKkGpjoZVVmqe8ipL69ciS7hF8y
UCX4mNItpBg0WRkrRcqRWsV1ln2W3Dsmnqbgjruoge/To4bq5Ls5ltdLeuHEw5P/jemWTFMD8Teh
x9D0jrMBT05p9+ShzktOHuPlUL0GHkEImKI1e61Fe7+lIL1A68fd1wMbJICU3PiCPobJBHObA6da
/RQI8Oap3qUz4KXOOUbbk3XlCjfQ+XW+Z20+H0+wsZPZke2/baYviybexuIJjxbudm5G9dAdUvsA
1BlSKiDJos98+SWhtHhGW0X+dQFmNMw3MVkDcWCOv6nzy9xP6GIMG0twkDizI92GgwHPAhkBxpu6
Fkax4KI0azai3bxqPHp8ZWqlrEwnpehP6f+zNYYYdxgefpRcr2vQbwfDrUNKe3vuCEAD/n57yImb
pyCXjGDorugI7UVGwUC34XBMSWaTrzPEvQVcKPMjSSLKmpRIbnWUafhD+58HIUqI3u0ekxANg1Cj
4cg4mXR04ayPRZpoD4rLfS+ytoFDwkw+FZ6c8Zv6/2PcAwmO4pV84b7qzFT5h4RfMidm08hLJ/OV
uQ2CvsObsRB7BJdYpAma9IwFgrCUzOtqNufgL5kfGfZ9Y5Tiz37N/zZGkCRu/jGuqcXJ+CLNNJh4
FpS+jr5btxvA90vddMppu5zI52wQBQ0LqkDKd+OCriChnWMTKDqC3kd77pO1zKV6OCYdPvaWfM0O
1k58vPFs/Te4ICNtf2ebF5PxQ1ssdfAUx3hRSmrJjPHpH44Jr8da/gwVRMd+u1VUIYuFDkuo09lX
yL0puqlNcI/tr0IyULHr46gbyKK9qfsBwIlulzvOZKbj1Eihe+SuTwmEI/rrVUbLdxVI/G3ULv+q
7VnVqWed8DVnmq2tWkIchM5i0PVhDL6CGZvRZeqFYroNvmnmUwYA3VtqpoJgRreTWAQwcSGOGspw
zrU98/FKk3CdteXNSbQaA5sQPlRq7p4IVj1YjHJCL93F/hL3DqiwVbhBLRDeRAp5RwsUFSXGbBpb
75NLWSwwIVNaPX20+nxo43TawykK2/CBEj0eu7WfNwbSU7Fm5k8+jSZvsY1PF7B4HNhkyGzM18g+
KjB/o1xVcmtFIHUiHBhPEfR8AZ/P0VwxlK/EG4dhh/VvezjE12yjWE9GSsg8M2ybXaynHHwR3+w8
4i8dcNopr9qdOMRguRA3ewlF/bCx111W7EXbVAiTNxwVe5Rvh+CiFJacI0c44c1tcErlYyV0Jxo1
ibtGZIy3MX2qTAkafLxF75MT0GXlDgMM5pCXPCV+5mZiLpmCnXPKIxvm92FGIWUx4PB/icpRTxiQ
1gkGFfpJklE8Lsy+WqK8YXuFmhE5GDnphi612+xF6nL9keFRekZA8AbaD2++l4lkWNZeG3ZZjhk3
IS1Rsvr88pQf11GaeJG2snW1GAFcCg8CSPy5Ym2v2uru89K66XBEWhPINFEH5QP060RKgS0gS/04
t+XB5sa8tzYjdoCDrApJZi7td/LMDRYnzk0rtb/DmFdioJXXY7qpMflZyM0/IaKytZZNpVbzn2Il
Zc/VFddy7iO26uTMC1hHzmn4WWaUylShyzOwcrmSsNyaJSHSOwgkGIjZzbV024UVKV3TRpGbH8Jp
Zdu5ogQIKCMLRDTVRMrfeEMXB9NwjNY7RgrLQhE3VTj/3HzJ7PrjPlXg0n/0JQ21j7H9z6fkFZ4/
I3mn8K7f9L80jlrjDJz1uuCElnrZn8Girv9bN+A7IFsYLoKQBuuQsWXVtkcjVw/zFP0m91iTdQos
HMnlKFEltmWnT9axIDRdW2UdQNuK7ikP52+eG9daGzmxxzV5cTtMYjWZTFiA5YwClpCI1DiVAz9O
ogM0fvFEksp56mT8AlFxueZMUnihVd9yzEHu5CwebhHV1HY3ESrNv/ero3GdaEUj/j3TpHQ9S6VA
LTEGUY3pPFXyH8Ewgc/cYfl5WZVULSnKC9bxP9MB1xdm9UBCrftpyEmbiNOKhBvLPncFY+GifePA
78HQ50/yXrX8/FTL9r7R/AkvNVl7cgsU+SZJzxs3fUzDQ1Jbx1bHZus57IoNlbLdzsELtoCrDZGJ
Rdrasiwox3yf5t11u2Gxi4niyH5s4ka0akHShdFN4sbtw7MmRvx1KpZqcLashQK3pFhul2Wr7oF4
EPkHPKSr+CMWLKWhd9d+pC8d/Vilo/q7ayDydPOH1u+P975vYu4VyhJWfHjfAyNzB6HqWCNrwEyB
k20pN7YaiZ4vH4GRBOYSXTCU550A0Rl20jBIAYFdK60DtUiHAlH+FUU1zzzGZbnyMX5bK/MsVt2a
0fognKS/2nwXzUBzlkI+iy6IZob5IifFUqS61g2j7T0N7g4EhPozMeWe1PWpU7kA+FNlH2WbLjP5
wh/jQz/5DQ3OliNnJqU+kzaJwLMabAJ6I++xOPpmgGKyExCKuTEU4SoUk/vTDj8ald6ANcxw2wrV
NPW2w6PNatKG+TymcTrGP0Xt+BefDzhqsaHoK0q5Ikr+IWl22Z+jfSUxaoXRry/V2syDkgceCOcK
T3Fy8bQ5xBQkfR6abquOlyXSS9yjz0xtNhq/8kF8MYHBVY8zLUptCTXwHxqLsgpkGQRSOiFcBKHX
cqkSuAfzGVwAzuHzmXs97oL4O3HvkpzII0XXqHksZqLvGaUt3eTm1AMehYjOi+bOGTWda+rChNhg
MgCgM2kLDIZOAggGH2TGDllkFLa397EmRIAVyBpi0M1UmmJ401rRLpak1ZI5jV00mHHEqBxmAVMh
RCwwRze0d7iWx25CxuwSzkA9BzeMcEqCUn5mR3kGeq2rsheufzuobMTUEgXGPvyhaWkkDXB6Kny2
ToYqiUxYQ1V1F23yoFP+W0P7VrR298ds1ARiwWxr8+ABqBCyVHyVDHFaAQtutpzLi6gflPXWChSi
pPJ+2TFKLC1mYt9CWBtriVE9Tk2+ersgVoDZP55auj4PI7sRS+5TnGQzpeT2q5eeoy1ep9XEzcmb
vc9X3QKe4NXZpv0A5fxlKUOJKtkmE5i19lACG38ky6khNFPSge4F1hXfY4XsVnlHI6Fq2BetmWWs
avX5/sbw8+vBNYf5tHEJnBfVnPJgXswUrCgbiom57CJYTQA57a8CiU8zmu74OFKgR+loXulMLp0G
BuhqCIgfX4TElwGvert3h5S8PBN1uxBbriFQErpFsMitOOORlAVJFyiDAvwh9xCKCtD8+49D3mXu
CQfvCztTpjctoi+TC0iPpVfdjTT4ZCitMG5j7i6dRBbWSeiD0KRHtck8uYkrc8gV2qtLd/01pHig
7j6aFE1xQHJ8MCA9+ixeDuqEnlikLVzMMXNv4fDtKJ1Y+U0NOmLOUI6BfIZMNqN6ZNp6D/YmEPK4
FIg/T5P6dzXr8NUYaONSD19V8xORbWnxmob0oiyVqgAlP7pnOehG1j5gVdz1ABaxC3tiBX73WQlI
oGVfxKw0WTSdBonHEVFF8gkpianido8ngOAPRdYYTXvG+aIjL0mYung0zwba8hPug6YlM8Ebb/Pv
pJFCGTnk9xJVIHHY7BZdUsFTeG8ONk3kOyW8hQUNjxJ5hCccPxEOSx4lzypuNRCJ2qstlOVhSvP2
5V2Ei2Y8r5A/A3OUHp1spe/y1jniVtGJXwlIReZWcBYyLvXqfG1s46DBI2hIv1fw9ghFETh2+ljE
7trI2P2E0jXPw9hdAidkiC41QTye8SghTxOxTWJZVBtj81mA3mzp8IB6ARwiIpKHg3mujQ0DL5jq
JsfrjMgHZb9Te2flqP+m/ojZBVNp1lbuQMdkJh+2X/knAHxZfKu2cex7dgRbVTOdzlTdj7V7ZMJG
NOL3mHxIRpc2If/zOsvNigs9dRH+G/W9luwEL2hzHwUmz13FFoPFjx1970kMcSPLt59S4c3mhJrI
qBb27V6NQ1ivq11ZMjkpPErxArdsj81wY2lruci+KT3TfPzw0dI1kyGa94GayVxVC/WfvriP32g5
t+GbS8226O/XqF/FeP6MU7Oy2kSNPgRXznfL57w9GfSVbNsjQ9H/ezzfB0mBP24PiAkzl9Rb0NZt
Olq3JgsT/0ty7YdExJRUsCwOB4rTf5ctBZWy02KaKxitGQQc9jiZv/Pb1tR5kvNc5WrxAr0Smuxk
hIbuYYPvmgVKelnq5HxH1Oy0syVqzweOKyTp8PYjG4a0wxzKmX/4srd09K7wD5PUFIl8nWxFdejf
LTlqBcUIlJAwbh09lcukAdsnUFFX2oMzbMpS7dllIwJnRIaI6UO3TUfmRBavXxoMYjkHshMHJAfj
ag0r2vShOEq3i6Fzwfou3ibO3gC32dYl9djG4HCnUldeVSygTLFOraTE/Lj9akvg+YctDGH2dJzi
ZFKk8XnOl5gKKT9OlQpfsprsrBZq/lPkDohsP1h5ei3iyVtovn1/WJKl2HhttcWlAjeRY2nFjEb2
yU8WQboaPu1DbJhWWhcYMn67O3eOlcAeZc/Arr4dmPJqJI8u0KqBk/U1P0/JPyved/x4AT/i9f3P
LsMPkkNuxdvFc6xvYXi859rGSu9SzaLfmSpzFuBhEQ827tzsS5b5QmB4ghUPXaqJ5PXUhMRQNmFq
VfGPPAVI1B88jTeW4rQsSDQrNNRM5Kvex2FhQzCDDk/F05FwTO++PfK2ms3168URrCuLlcFzjYLO
BC/LbwQo4Zd7C4P59wi6RBItZ+7DrGH/fSoFVAc2TniiP+z+FAKCE0ANMbAQlUTVhKK93xCQtc7g
xMGz08t2H76UISNBC118lO1TelvsWBaJkRXSvVe6/gtM9Q+K+ERrnBGc7upR5ufwhXnURmPlKi1/
SXeJYdfWTBnetCUFGCK2a3PjfdcUD2RCBNL3KbwPkB3MWvBmtHjPXCOExUCkZdhJbQmwvXXitmOw
90iamYCY6eXayvTGaPB4UF7MDo0EjFKSNAWC09Lk3MJFUUnsOQNhf6V/ldCmSo5DspU0ui79VYrx
I5po761Lla74fa6bd6rp28ZUligS4W9VADXxdPbh1CcGjBttSYptM0piYVsxy5TfYJJjeNyLdhnA
5zxZ4pebgPejznLRSiGE26EiXH+e6FByePPPW4v+mi1DARE+kWZ8CXVjVNpZLh5dN/rPvRQeiYAt
ZEpmfgkPmPcPD0MPhYeoVXFisbEUBUdyH8nfGzumIkj5kuMcXewIN48aXYNWGnaP58FjuMI+hxXT
z8Q9jtxaMKIFjS1qJ/WFRu5nCE8dhBXLFxyfO42A2m/jqjq7ODISlnQef1DnO5BV61dUEWfWeDiq
806sT36ALIpuPfeCmw/iRkaXWv1J227pcycv6h8t0z8yKZmQTj/tZQE2lcySnx48YPvkgmURgRH3
Jt8+0/hmWWgUdjvn/C0o98qF5sLX3N97XuA+U4vA/gyCnIreBv+y5aDn/wsBahPoYOBO0N75D6xr
H5ZHWS7WzOzPOFialRjyWTax1uOZoJRLC3MyMcRDU37Qs3Opg68J8faa12tR4FwTa6cjKjG/eW/d
UtCwgrKj6b639VKANfzue0lTDy1E9fyMY+J82MN1jCa9CZWc7LS+5p+DdGRYLuVoXRJgpVJ42AFo
XY95lOsFdAOsGqPJ+/w4860oasvbiKOTCRL1EHVTdkrSdc3o/Sn8Vmp6dfL29JvciV0kwJm9SmS+
eAIBO/lYJz7a1xSXhBdeuoiWOT4RS+rwfV+iZ9s9OJryzBiLXuCODaaiJCqwkgM/spXSQJ1OzcNW
IhGfHfLiZaDvtdRCJrzthz88g/rSxUlO6F6sHlmEFH5RUFx4SFuZx9t5XJA8vPJprJX53PX8AHU2
njUaV0P/MqMMJrF93NMaLTstW3np7t4mCc/G0W744/C5P5EA87H9LSXX5rI4OFz2ur/iJGMiVsan
Xu30/WI7BYlwYgB48IMuLQaxsh6dfEQXTWF6W2h7N6Va/uAunDDGPYy35zBZE5FmrNGlXA+1ImS+
6qIz/MUnlYdVVhyrlUWGFPn2JbI+1Thw3jJGna3/bEasM2pcfFeUIcp25ZTsjxTXSnz2N3T2zGhL
fTdYccD3sPdEBlR1CSiV72UP8YDap4LS/IcnH/0it70VnH9fNheD1j1GHoO02ENCuRFMuEZWtMxd
bSLqraYhUMJ14ERlimoySbZAZz130n8Wgse/ST7mxhSe9yBYojLcm6KdX3PjJ5gj7nX7gdZ+PoV1
1gGHRsd3+6Yj1p52JMbeheUpT+J/yL9LWe81vUUCaD2cKz2H2YhPY0dXUkUpbLHqN85ATNVKpuTv
l+HY4hY5rkp54ZDbxOjof+4bWoWTrdLS7kZe0CajDn/kf5oHE3RHhW5NhdEqUJFmZc6iMIsBS271
/uVnpJOXzJjjH80OXkB8YXbdqJwOmC8VyUCOxnrZU98VAOIwRR+eWZOUNsb1V+aewmlDsLMpzP/R
FTnwJu53augtAn43jlXsEEaU7yKuAgyuwRUjvbcuGmNDw2una3iMO4DUPAhwE2bPecMBj5HVUx9y
kLgruGAlKoxzEVAVk6/ZiQlrue43PL0k1wV1NGOKYXYRC5iDq5TQg37Jw/pUFxuARxNH2OKOjLFe
i0JMpeKJXWhWSeD33mpczsrCzTnQZq2p/Sdr66TSbElSB9vo1l2Ekc/+gpFVD+6jZVaPOPFwatfy
LpNfxmGFRBt3Vh6ZL8PSc0NjBkVs6ov1VtkNTKKtYoVOSEzms1/wBohmcSLpUXunW/nZ1SfNdTVW
F95BOlzv5DUyB5mEKRV4LFvm+AHO0XGh+ioqut0NUcgsFJHeSWYgGSrRL2lwB4CspfDCq2roku4m
qtpcOHUl+acBdd2m3VIYZQfWpHHxKP8PVZ0bxf52ft5bG/AaoDMML21vs8Xby+x9MbSX5X/xr4Wt
aBNKfbZCUQ78iCr0zu9pdtc9JW1VcQYgPoQgeJo7CcuO6+dwAOiRH/iGh689OTpzw4GkyRPob15k
40WCF3YsaHLWFnyYE+Nji4a+wd5sG7lslDGh+aejjgpvRAfPN9dHhfE7YDQOMFrSuGMpbyERkwJ3
FcTUbaZRA5qMUztJpPhjfGLFPf+xio4/nABcdAUL4asVa4+TPCSuHC9cCmPkrEYBEddQ4iY2uET9
4yr8O7HEYo3UgXxHIwTuftS01xkGqkny9+kNpUsuAuZyUVvjMp7p6ITi6csLRcJXwNfTDDXEbfpm
//LhUMiF/2Lun9iTBywz75lTEPOttQ5/ArAczfqCSJY/Qe8tkU/O/1TRRnIv/LciDxcG1xLLldSC
3Z3JmXLizumSTEihpUhZgJe5KgTiSq9PnI5fXvPr/82MY4ZhvTrDJDqinbe6jpjhB+SUMFwPmYTh
OTIRx4xobBq4PrTNJ6DbTO3Pyv0mD1r0qfio3bJac1SNX7xz5Wih+OhD9sZ/G/D3ec2m1/g0L11m
gpu5K+HJeA9LLJlbnx3aBkHNeca+x978UX4BUg0JmhDv+If+lSPkrWce/mbAKajU/6fFPZeGV5Kv
i5Rfu41A3TLrUrEZ0XuD0n+btXRkYsj4lXv0MQcaqjoiU4HOD/gYQIa1p4Mf7NWjYNbCQIHGYsgU
JM1WNVBYDJOLRo6dbj89GxrjMiZKwTbSAJYOuSa+xwCT4SSBFnpp2B2i/x1c+tYyH4QkWi9muAfo
ddMChm+cDRf1bfC+uoXLASeMYL3h000Ejn1HGDIjV6JkXlSdcQnj/OWlpZmlo2jL5gfBbUc916xE
r/rJlaMs+RTdzNwTUNYYYZwquvl47I3xIGy5zw1v/u0P3Po9otgfFyiWj7fzpAsMGVLc9FvxMn8H
HcqpwEUKloa65hHBsqGvAaZIIfin1jxnrqvsl0ch2g3gmG1aujlbBIGosSpcf7kOCTudP41J7jz/
nTTZMgRyGLpnLW+Vkl6431VgQi694Sy7ga5yaog6qEJIDntWYXPh0ICpIDOSFO/yS58RRF6od/bD
rs44f0I1f7bxaIVYolnvV3SuOESpOo2I3jRcgmOY4Wkn4nbBBC/ooK5YR0HdJBcV/SAYaGFWpJDs
fcTcuqgLt1xSeEOYD5u8NOogfo/g04dGdK6nyhc9+ghNzErjRiX+isPaVmyz7fLokGYmtHuIsoSg
ns+8jMAj1iAvbqScf3vt+PE/yWo51hzKQJ5NI+oniVcR6QlsPIDHwlqPibdkNbgjqRdZ7n2YytVD
QXim/UL4QJwuX+NzyILHwpWc+AKcCWIfbH/cggmgFZEH5OGeuhau1EuqqQEdZWm4Bq/UPAsDkKNX
V6GB5EqXu2UHimr6IeIs5JWeeXXodRoTjePd5qOm+32H2pGopQDkv4WoKY53H4sncK7+zkK2jNIv
v5xPsgK58KDc5rUPU8Tmz8bKp2AbqaEysE9mc0DS1KioYdSqwYHRmW6GCM4Gu9DKB7ZgYTq4zx/V
sB4DrzLuGdCF6JCPgnKdYc2mniqgT9pjQmspMtfJXwzAtspq6+ofRQW2oBt+MTYbK45CvFbVBc3k
Y5fLF/eveXewrUwbtfHGp0roEH6/7isX0sUxmTXvrvizPbJkEF4zSgiP3m/2rYt8oMprAxLjsyxl
7ANVgtSmPyAdVdi548yy0iZPJfntQa6fR0/FC7CVSwDAhdS3YSXDUZSI05gDKLCEm5PCOMG2T0wu
B+4OHSnI1Jg1svIstgw2Y/o8b1rswt54vNZYhoV7fRVjNVK3cCIj1EtqwN0Is54uO5CUWSAfoBYs
Lhp4X2G++FH5ijfyMp57LSXCvcwAfIjHEptgiTY+9QseOKJCmyjuZo59YyhpWnF6t08+eRM3DC0y
QuRDAWsqhlJDQmd4XAoifLaHje4k+W+CHzI9iOXMv+SLFA75RbIUKmx52Q1VopMHUrAbgXjz1KIa
gUAFKcHE5bWj3aXHCcCEjihx3zjvI6ozKU4NS/DUDDmw1cPFTudK3OjD95OjTW/gf9x4Q5EL7djE
thPoV9OxrE7kcORropOjdRc/WBHTxu3ovlHvvXT1em0tK30EshHYkQOkIdLUtQLKdj+mWPi30fc6
zI88RMpzV0gkFUWJuv6sZC2iJojAL19D7CW5r/IZgxlhcMlXmUXaWN+/o0tEAPTWjYYKp+UEvg1/
P0nOKl3Q9goLW72ipYc9BcgR5Wz3REZJ+ElCYWlrrxc1qUzaWs2+Cvje7d0x2LS0hlRyz+aM6BEc
mu1feoKxuKSr9zu9ZeSyf1KRAdOWG+LWVx515IEvGmYKYMFVq5oqW6ms8/63243JLnhAElQFFWgp
nV35OroinQDpiGo22XeYxEq6GwHGkNMVGg9vgbqJ+wweHVR8AfhcRhPWeO1f2+rKV2EoirLHk7tm
vdiOOKg+YCCTGOgKAnBUrtEy6DsWzXPFQh1UyPWwO6h5Hh0yI7eFPHFF2C2kSdRvOSFIhI0fV2CY
Iqsoj1Mnge/7If8v2S/yQJwBx+oACkgLRfeHOpvx9nW8AkOxPpOHKpmKjNMQbwd+cjWJcT5gSGJR
uYYtQfDXRTExt6JVy7o/IUpafA5aGDH4xts6nuqceLeBwodGue8sGKRpQowi7nYZqCr4RZyptn/N
rrGH3H9bBKqLdG3rB+ZVOsaEnDXUbAR7M3jl9nGW/iTUj4+QkeTKCCzuotrjspgn1fCKxVFLY76A
qTmyJmkV0fVRFheYzPEYdCXSI9LtUXqfKDdXRc7R4UNlu9KH4e37Pd6rWw7H6IayQ7UmTM8LQ6wZ
yzZf1XrdFrOpgxeHM2c6/jL6wtsyIuJqEr2Qxc7dxbEIqdGAbgoLNvbWRTcW4DIieyVeSgbVB49Z
U5c5SLdnL136pD2mo4fG9IcJx6UFf5HQsu0GsZUnslQCevZ1oL2FQWWSe4OONPUrSB6wCf3Epmkh
YLfz7CKjg/26md6d4HabjGETX8C8JOTSswtOKxwS5Ua7kfK1YGNfnCGgQfPHBs5tSdQH/GhiuJk9
Fd94GLPn6sijejM9/+1YfmzPHN7lPD9cyUMHAzj1wUku9pLnQfNu/ErK1xvf0pm057uXtG8q/oWc
lswYDBqdAZaCFf3nERE1T+26ydgdse41DUfbVtuvdY9LL5FFjAETYOHrdEI6P30KbCywlNO/iZdA
JQMUhRL4M659Fm/3U3ZQ+ZVMEZsgVX1UCCAq0o38UrAi7U6AinY0TnjaRtzON8y56vV1zlrN3lv1
O1AqSYzP6Xld+Opb0aSkpILznb73RBWi9BSUs6dJPJUMI4AeK9aD9w8LuqLjCtNBmMOkP3G2vxZ7
1pDzwHnlMrOMuDMbmeWhNx507bsLM/4C8JpH7KnK1BWUADR2c+nSR9xZOnieYupCSeX03w/Gfa/t
FGazk1DFbicDw1w3Dc3BQ77ijZiFq6pKqm+yxhiGLvIEg0JPbu5CMdg1PyNajZN/GaHghAPLO3xk
yNc0/MpyS0x5KyOjPaDwNbPHSyt/vOtCp4K4cCoLrMI41WEUxdxGmd793S0h9vH/rn44Mn8s7vwl
IF1gZURyKCTKIhplUw8XYoLKmoO8S1eA9bekSOXz46I2zOOT8TX3qPtWuaH56r9WEHbg+JkH97H8
BXc0zCOCji5NfWQa5ev+LFudwzMLp053w/CxjsdhZMCA7EeCMy//smVDBv9GPF0sZAe2dEdM1y4u
ZQR2AUSeC5hzVRxcurGsXS5gJoAvgtnA92SflD5WU1JoX8PasDEptD4XD3cpdomQDunmMUmwQ45l
iukVLgzpvjM9mwgYn3HI43JZIwdk4slPhtNkvaXs1rM+Ih9lwHS36LpVWJ5/SoILh0OpIKYhhvxu
i4kccttzKbU6B9BPmwccBllum+Ta5TfQe/ojgOcRtKBlqsE1UIrkYB+oda5x39t9SV/1YJ4hIPN1
bcrIGyQOpF7O5pf7ybHAMbf3GNLnjIfTCfaT0fZqUT5keTR8SqH1WkZXZZKBRfTSqiMB2hcby1fq
IfULlrxx5jv01JJK6CKwc8F3lM9AdPnDVh4/+YRtUwRGTbWYxKA76nGsP2VU0qWZdrQ1g1ZZFpTK
OskBOtWreJiLIVHMN23H3kfg8JjwB3QgnmPbjmty2VWG+6Xt02RDdjGQ09dMC/0abL7lP2O4sfVg
aEzl4+vPoLt36IYfaOPMcxon8x50R29ETlYpnp3b3K3q7V6ASPvn55B0qIcJP2Gj7YlMD7b7O2aL
y4r0OVTdn2ZqrvOqqLK2vd2opUcxDgaRx/I7ceO6P5ecfQpToV/q61k3dkwrXTWFdUS41bgXlEe7
pUYD2P3k7+BSvqD/LpBqpwYJ5rLwZBXZXZ4yospgCk0go5TyLw4OQWpMHevwKLIWdrJFiKRatDWL
fBrUIF9PjmtXuMFVeEpgYrS7B8DpS975IL9tE/AXYJhT7ZSLxM2kxcb7ymQ3s3YWtFTi8PX/HU03
KJE8fkP2y61iURJIfd0g4M3n15aA9yPR6yargd/a440d3yJpCGsE2cNeQ0XSziL2VTMTMOisbe8w
sFyWhbjMatHY5pkkN6b6BnrTfRNboyPQFd2IftX/oBilp0XeRJwMLLL8bjnn+5HxjpMCtqvWn2+w
CIoZm29EH45mCQdHYeWUP+UuSh1LFQQNb0dNF/iJKQ58J1dCWzmUuuWJh6EXN3vxsD7zz+rYXxXn
jArhSSsAYhvjGsB5mxP7hc4D8Vv+NRfoKWIOXNrYhMCIiqNHD9qu+wjB7U9eYYsjHOsQWn/a2rq+
FSvgrmql5/KxdHTMbTgIrjysRxB8KlYgjlDzubhn8kYYy8Dhgi5m2YQmyxbB0h9mCFwwuNiZFAxF
3e79VpLh0dQxcJH+Vmtwa8cC/zYdBzHyEU1F136tRt5BAWJm7ADbl4l9tD8ODRX+U8BMgxWVuKYG
FIxLJUxBSZAMJeEHPN58311CLk4j2EgWzKmqG7n6KgkD6ncxBd873a70LL6o7nUngQMBKo0xEGad
fWcfv+njmIamQ3m5zODKJ1q8zehhgu8pP5OQmRLKSXIIcLk9Wlx8OZpJaL++6b2UGa0ykshKxVMY
vohxH0twlUYHzy6Guitr6J+CgjsbtxzqkjE9PoK0nxzgMK0plRkI/oJpu8pzj39lcSRGI5dRa06o
OPowDXK/PQJVEronzdo+93r4aGiq8+65ZYNnF93S+icgpUKoOzpz60T+uvDZFd3gru9jGSsX/TzB
brgyRhZF8K1nWCtbTRkjU9/PHSOeZRDVCBBCKmHd4d2BV5DhuXfwuxgBOg8AcHRXwqWUa8f8sEQ5
Gr8nTanE1bljhS3fDne15ebLZse5hAKue1uZ3lKZ6J5dGyJXkE0BNa7scuoPFflUit92mCEX17ww
hYVES8TP6uIzAoV5QYQUQD2UTTf+gnG7BIeYLPWdOXKT0n+otT3lv4xxbhCtsrdW2il/jWAQqInx
QMSCYDgEhqxKy8DsX00xfDaqj24dGyfxUskNmSGXXJhuxPGHsnoFKbSFNBWLzn+zJJ4EBHBbmtGZ
rJXf7QjWLi6Om/nlZhqyVaYfqfj/TtRb5LUFB4g/39urOiNHeLRHFcLwERwpm9NogSOpUxYQgXbH
6AdtqEgdsDMMPh5cSXqFFMSnEp+w3JsB1L5XdiqwKvv2OSSLwFNY5AIqRzKNz+6a1QF3IbcpgpzE
wKFMSa5bPzp0Nmj9CS2jw0ydcxgUQx4tEVnUMnFa0aB5moW5xuJ4mJdBFqJgqM0lPP+HaPjluaF2
gwUShN/QeRAEUQ+V/K3kUsOwkBcoqXl63ZdwplzH8mpvX9kVbUSwYgAg/juZwHJUf1uLNXxu1fK/
sfugL7/zj74Dr6N1K20jful3v3sCsTGRniSwKRuK3qW8H34h9hVMaL3H/tlOtcT+s56FQ6BYfwcd
O2do4GzciBnUerskwkcCEPhYBKT96VM172Tt/h6+gT4so8dNi31v3kG2HFzbGtAwqw7ZERHzePgg
uLndYhDSg3IC2No2Fw0MBN/g4qXPpIL98hXG9JtRuAwwSFLu1i4xSZbxSauvEQO8LJvS9guo8DP4
tfzLH1QKE0Z/niw20MJJ8fUPNqnKOg+cx0o8Y25Y01wUXQyyP9G+bj1XFrTQ7pt9PAO/UntYoah3
Q1gNSwMJw5uE8vLOgMCg/rv4oWiVDv8qUtvlivPoyQIcqMLNJxHsejUzq73Cvc5EkZuNf/9TxnfY
ddQTEKAC2rxPUAV6XiZKIeWYcjwOLBTuy7kybTZTwkAyF8fjMxdC0HA68ZvNUujNneemGx1WEPMu
3/f99Absx35XWBWnSsFNhm+wxyZE7PpeqMO/IDjX8KaJp3g3r7XqHxNtxmTt6rYJ3LRumwS1k+xd
glVeEdBD0fhsPr6FevS6i4lLX6aAtSYYXPXKrfu//2V4VMDy0UKQntnYToZ2pZeFywokqDumxNxd
OACY+yXfmlazF84ubZuhrdI3+nnU7+NWvJSHbGKZT24VLntfrKI6k12/uPR4zK+KOg6EYgGrzwsw
tCCrO7Qp7XyYhMHScH9vs89lI/lVA8JEw/GT9Q4poA+ZNS0aOH5SpzNYEHYCcT9dEZlU8cayEDQh
Bhn9MK0Tt3NbHLvmGskf+GSlvx7vr5UpiCEN2oVr48xzPz+hVHFRoQ4+8QIXeZSlgVrtRA/bindO
piddomLhuGUsZKHw2KQsIaIPOQTt8x956BHxJMWON7ySG/6EG++efDkDQ5vNhmsHd5tiN9LUXUsX
WGrfr4FYdRrIEWyCCZ7oH59G/hWNJHIMR0XTKk1rvGGi1rBumJVfU457bAapKFkyZ8zf0K0dGFxi
g2CDnpfslGxlx7ddsLNk4doSu6ueZ6AslO4tXcU2J2ZAKsYbY/dispLdy5VToIwsrHLpPuCsNmkN
5OsuLlwYrxALIhr7Izwhbq1GhhdKR6vESfRyrpSGYRHIB3NPoajnkVHQLwGsEjzLutfC7TDY2rYO
hCyfZMwkFFAnYpDLfFabveDndLj3JcE8ph3k82m3W+Jc8mmYIsvUzNimNqUVtwcqEF5iGgnxATmI
QOy0hzpslcIk4wITqFPmGphJeORyVuwwc6qx/R4lkqO4MjbMgxBH9qeIqkuMlvBsTeWlfOoN4WWF
02IB8nOaT4qwp90j1scpfmuNmICubEbze3vCm7ADf0AbrISDZtVDHVeZKcHN5V3jG0nz09qlHY7T
9OrjoQPs6ZClucdTqbNUJjeoaHgaPhrfAzCaab1CchyRpvZ9kkHYGEyN+4a5YTxpDyclkpPvNrxQ
fuvFbsSwNdb1apzQgZbH/IZADa4H/YHBrxVeWLXcGu6D8S9s4TdqnoFbhgL80jT4DH3CPBZH8h5+
0tZfxlEa5N/Mr0Z3x6T9gTD7vJ1xFPS1uFwdxZZDYLS702JuWjvvGdN4JN23rGHsKfEV1vhJiNjc
RmML3+0Z6MTTfsUDzK1p7VE8v5uhxDxr+o8IkFhUMj5UhD0AEzhmFzc1AEG+2Dcd+zqzxkZHi2Qb
0Ri7woHT7ee4XPY2rweFCacgkstXh8uW3JBoCcnoeHyAUKcz+QqATcq9aqLWHfscjv5lFGZ5t/pa
2LTrSJGd/ObMowGDFGyOdbyJF++n9pjqyqEii9RFhp8iWekq253jqDyU6lbgMR2HW8UqGjM69V8O
WnXDqzDF8TVFH1xLI12aNDdsI8O7TtkRz/v8Grv9s/GmXheyP/kejleiCY2K1SArtOkYi/nUnrCU
555Xc8gpz0TmS1VXYOrZKwlRt8L2QXZHFNemkp4kQctUuhow/IetoRPITOALXHDBqGl546g3qHMa
PCKYDOFy6ofTXpgpQKJOqI8pAQAWG51/bfxneba1g1XhMSPkF8Ypf2JV5d8Wcg2jkPZNzElJENVO
NBaFTl8EAZAYh8R0f4prAiwJeaVwpDqzvSSI67/4TE+krZ4kgO8HMT5NzJeggpaVR8ZDnTZRC58Y
02AxjXlfhKsBoBH0ApUlOMI8tR+0AfToHY2QCJvNVDcykFYsrbrhr/N1h7YNGwiQpmgoPSodkujH
chUiO73FiSR494CVSn2Cm1ZjA0li4IBIPOHhNtdfTuVx6XEDDO3/6yo3Kpxc3Mb0K3rv2eSguFXd
Y1UTzLKW3VGxkLZjlUu3MYGNbu3AgQ/8Er+Y2qwIGA64wUSfzDTAOs70w+z72mwdVa//D/rr4L6o
f1RXnvmWusRyBQCe3wguEJgE+uNxxkD8jmHMLcEQW+O80etaTKhX1a1QahF923OMbhuP+Etp7y4p
hzpQ13mhoaoNcK/dVGQxpibdGCtsWQW1oj2y3b2YHU9wrNwHTNG4qz4+p09MG7AgYhFNeJDBiXzj
IswXtQkTUJNw+geko6gIKUUKw+HYia5rOsltHeKz1SZSpy/Wfh4B+AcXAUaYncviqpiRgw0LjRqX
zzLHmk23E4IlOcG3sWPXGEvFSliCYwKQT+Z9YLkfJk2cD3E7vx+NhJKoZKO8sbWVkS4RfInQNW+u
Bbo+Zkk6Q0lXmzT1DW5rPQXKln07nKERtsTixTgywVBoe0q6f2RReUTs7ps31Rdg+JdERRW34lea
bojGPRJs19udHddi62LYUxKt0lBaii6SR8lUYlb1hVEbNNMeBPwC4xIO6XupQhKcU0iJXkRxZDhQ
iCqWhBR+egH7IL5EGum8d+/V4/NYIlJsuuhURykXyv8OjrukI862UHIrPvA27iK5QNDLkcvqw/QQ
tfusr0ATMQ0tfMQ9bYMo9qWcxYU9CvTN448Vv/nz1tu5a9LW0UeVtv55zxwm/DCI2w9nkBvWZ74n
bRZ4UW9ZKPxOjy/Gkca+THu9IYOxBipZQBm3qqXZquW0POaSoXFPdqXpW5l56zl2VYar5Gz9/Gtu
+ajockzsGM55he/bjCq60gdEViFBJtIE9jjYkoje36Z6TLEm8hvzImntBCzwIr9b2h0PH7p8iLgR
YSY9/AaeM3zgzl2oCigOzi3EMykhpWeouubEQ6dKbiAyEYtmjxqyYl/vKHeuHEXM2eZfZnOhPIqL
UoKmnUSDE2sW9uJaiac83JmqM00VMWjg1ukLC8AR7WRbS8cIT4pqtTRx3W/n/Q3CNwQShJ2z0kUg
NX7VC8jJT6NMVyrkp0DWt1JrwSSE/cbwOFg8qGWWH+ZkF4mcacIyL4mCbcDzT8oxryLROppCazOC
3GhUX5wH62jx35ZkGNkFEd9hdLOM0JZcpZSlKbgDkqbtRGb3Fevv998WUak9pTkhTOcEgB7quqSj
u0jr/2A74Sh6u+yJdegRw0P55OYSBYHMkQ0e+wG7lc/sjEzDSHgojHxj5I9H7gVxzF+SiS1VRV0n
0iJUtBWwIwbu82iaif2czutPTcy3zPgtiDpVpLdSVpCkgxkwY468EO0a0c9u65h6qSsoteKm1YoE
dQxZ3BWE1vg+sN6D6u6HJiD/y04r3Df+P5z6SBvOSkrbohzPwsXI8QisL5VyXU+BYxvV3KHXnwYE
2ahT/xzySkXjjDJXI60bHT0/n/fbJu/l85fQuUIlFig4QLaRMYDj8a4XoLxWYKPBRaxl0YSItb+G
Es4ctyADBM0VLCbdVxo+sOPSnVTdCOmlS6KBj8uJ5gXXskJGZqR27ips+eQnRXbjKG8Ffn1dTj4c
dThzlRO5rosF349WR4lJ7r3VhURHxuSne6AUwysUJRev8nynIOHSH6RAzGT7dYSJc5Vk0YA5vT4S
EeKaWXKd7EBn2hieAXjPxD9R3eGiAx4huc27Sf2A8Sv5TFz29bxTvPfIwsm0GXfHPjZQNNtlEpJ8
R9XbgN10mvBI+4Vw4HDTG3EA0fQ6x7My+gU9Fdj5qWHZfO4RrP+oBlIzLKE1UPQBBsV8Oee0XVUl
BmdJKE6CK0OQHCzRDHgxLNJ+QKuF0fg1eIQeNp+z/XF1OWUwEZPdYJ2Gv1kFiWfDc5UePHUzaauI
CERWZ11FjRIklhKkTC7Zo9zYx2d1nkGYAjDzBDF6rr9+kCJf1WyBIZgzbBU45JQuRc/0YAEiudKz
JejMDuXNZAQXNodltLewAycyx1qmQ3RKQ+OMjvPrXkL+9n6GTbIb4qdI1Fxs25D+roRPLOFpMI8T
32Jq0jLo5vNDyQ/JV2V0l9ah+v4vfqBXybQln1bZfEVSqCgDBht8dQpsSkL0jkhm/w5aVCdDREZy
es0hbtOqNrNOtE0aWFVPt761d11l1xwCC21Pl6HYrdU5MzHpg6DQC4Jme0Yh9CDgSQQyBm4Wom6v
NMS49ciH1Gy2m0oiZOfDohoH9cGZJ4vdNq1dza/MnbQZLLaJDIwmCeaWiixPuT/oumsrGe/tRkmb
pdBaFlH4zvumNhow6HrVU7b2muzmC5Rfv/tnlh47tXvI2OXHy0b8b6VSewA6RWocV834b6iXXcuM
wcsqoUhsrA1YXrUeGAsnrJ38vRWDWu6wdTtWN6As3gBDMRUeQ5E/cFxClG4hMEHQ525Og1o0k+L4
/yVWa/O/SAEMvuUqY8hbfMIXiUqBIJ4w/Oexx0JugLGJq9mI4zWOVtLhf39ISoxn5qWxayVV+Js9
u9kbGas4CdEFNsyb/BtVza91xirFLn2h8YZod8O7bkHPTNvOCAFxg1cw/vULw8ygUHXh3TUQfDO2
mcWLK+XZic0iQ8NXalN70STRwQFeqCkznWAIYu5ZQj9Pv+SCn/UpSl5o2cJVsP65dd2v6JOSuurf
r7jrOKxKS5Oy1S/8pgMmeHQxlEdmjUW5Kkhg2mck3u5nqlKUMz7DXZc3ztSG+j8tbHKBhskRRSJC
7hgniboTM+0kAkNH6gVKERqeV0dM7Lmp+S0kFX6nuS+4R8WBGrwn8buIg2NldwPOlaBJB9yLkblx
JPtTK+DBEraK7NUIcYcIzh7uCny76IeYugTLD0X/zz37WbRYfm1sixk9FOyeZ/5XmCKZ28RSuZFm
C9VTLW43J2sf1UHHdjGrTsnfRXjkCAb0N8NAqrNbWwGTFTnRPMNjJ/Htyy0I5Ws0A8zuMw6xJdYi
TgMgXj81m4A+M+2FiMc4m2wnzcbuxeuZihCu4kb9a7uP2Ucth3F+rcN/FtioWzirjoSVSlFIX6IH
ajLN8pj35esGHJFaxAwuTTeiCbTCjVfSDdr0Ok7mMQdB6JX9DCOggiAuB/RP/l6YqrhH06GuC1Sh
iWra9i0OOh1/NTmwWYYk8R+TA7BDOa4qwLTLcFBnVZRmX0zjOO+QYsAhrvWLFmWYTM0DjbwwXMtU
ltrl9U5VdiXiZk/FvhMNQ02YhwHhDK8pE5pudCpr8gjt2YmeToJM28pgCtNQ00rQro9dI6M4uTHB
vPviTB1pXQX9bQL4zN3qWRn+x89JNtkmhue1ciO5tuAnr/TKPwehy7jGe6bih6WnnRe+qTe5yn3X
jKF2jDzJzHaOneFJwx/5ajORMxNyD792tyFI8xXurlXjXhUoid4D5x6f2pJfd0QkX6/xq43c8DKm
ddv6TkGVPrD9uvJ8q7oGjBmNUe6lMb6mZzrP2dCUS6d/keQu6QoRCK65B5ZKmOghCrQAcYcwhZWO
HJaYeF+jaoWB8pA1AACINmIL6TqN5QpLIwS7C5FIQQqaqKrizHKO9pi5eXB1nJlLRkOnzyrSSVou
9cqIi56p8DtEUDDZBwfSoMUwuCStRgdQJR6dYVmVxuGAM3E3AQ3e5XcVTBcjxj1SdyfVOvfqHONj
tUYM0pKeBM1Tlq1Trx/IasbpWWSKoYXE1uYBJvVkse2oAaQgCcx9CErieEFgVlR9sTPgf4JMQUbt
sV2Ou6hExpreDR6YuwdyomOnF+YNWYgPM8go+PGOvr2XjQNtMkwjMo5X4W+lehoMJ4GwZtTdOUIP
+cv/2betu6h0+RRdCanSXbeN9ySTTDxwNQuMDlMzgtwMcXNg7vpJ49+55qkaEZBPNEW/gzJ0fWzw
6cyXGMOU+PTZqJXVIFPL77S1HvItCoOPWGYCF4qdM7WfmsQ7OEq/NMHmwKGheeg8xZ2sgtNPlOt6
2cY1qQN3qRvVJvjCCd+Wq8a+9zIiRAsO8o2Um7OTNVbV3BWFXkn2tsqJyMm/9hOcT2A2GzjWbmzw
L87NmU83gpHnFjtolTUTNb2COU4kUMq5ZNqzk2Z4nykEKxeb8/8JGZeEVF8XHAgSndtlJrYxG6TV
Of6oZlZqziXqKt8ZuNtHr8UieUSqPf3YghMUwWT9JZeMIxmcz9BfrmJJH6dmRz0ezaPGBu+KElVy
rD8azjvkuF4zR/AQzDSKPTunD9bn80myoN0CMYxA1GrZUts3Nv9nz1lPP83Hl5tHpf+hBDa5RWHy
pk+v40Wihs5AofhzDQgkk1UfNyPOkIygifTmX1eyd7jzxpMwY6loShUoVpiN7rrHABuioU1WQqXT
1/goYtjT/QjXZcWILJlb2H7vRsj17YPsMzqY+DmwUI7uIAjjqsVZWZx3LmuywGw7ENHE+fMp22dh
hjy/q5YCaEmanT3oflFinjpHUAnNyS9cQG0RkFNVJSNIQaMNIpvJdNED3MgK/Y9v5+MYcAaNFjuy
CS3HHX7CpdeRnLQP4gvl3RiQl/i9YyS+yEN0Zq04I5uSzs7G8GdRtczAUwlyAtcgwl8UOaCU2qOa
cLHdRU0/uLfczq0Nxy+0/s0OpDZ0vGv9hKS23tVHXeHDUPBrUqNcJuP7zLEvmn8T376k7PWwKB/s
Sid/VxyzP4aouk56b4CQsSTawDA9CD02QZxNbiRAZwBIPrGJqNf0YY/XtsFoi44i5g5WN2i9tLQd
Y4uQXTHP276OU/9RH3xUYsE8z8kd++Nf4J2Kk6H82vlhOBKRDYyw/7ukOaQaJYE+0mU38zgmciSe
e0ySE4a0wCa5DW/wYLVpi77ZR334kKF+GzgLT1Awt5kJsYDUh491kOc426NJEdRlJ6rRL2fakRhp
AvL0QB3svtq4wTh1FaIiNfYd94ZjokBOfuGi0eBIfT7qCkPjGt8MErsQTSWWPKY7BDQANHRwLciT
UHIl4DdStpYxYvO1XTZdye75uVXPPjYI3qg5kiexl11xTNK6bw6PGgNi1olOzKZVpJLPRoz1+jQm
+FDaCuLMEP6bRs8sKzr/vM/EJjnEeNIx0WWHrVjBSM/qf7e90UsH9DADxMRTApSNRPpy1alLZFGT
Dk1dbKx9A+iCB0AxZRgREcNDCCgg49TgPINnpKwRiQQcxzvOPLkniNylRGiRfbw5EoUffZ85M8Bx
p5hWiSnn3v1LxcmhV4/pTDL8j+6yMx9t1Unz471uGjvkfilqI0J7DxIN3LBVzpL3bnfg7xIWW3KR
/tRDP+IEAi5ycebQRByopCP7QWI6M/pNBwIjGuhgsSlWriIXY5NgrjM6RUnpa4nvw0qQ7vInoJsz
WLb+OUm22G0+nFheUpZnmWunlxI34rUdL2Qe1c2VZagq51rlQtW4FVRjm32vVlAOCxpvyETP3q0P
Y49MUxXU8ih6nrX7eTz9FrVhb5MwcimvlT1a2AHZEwXr605S81nL+tPhtMeFSFkPnrfWHA3FMDXx
DrCJwVlWWZJsSvmG9P1+WBlhPn24skiwWDhS57j3WulQJGIyVD10etLuYKVYC3D1P9Tg0xHNa248
xKe2M/o0UObV4O1xbp6wB2OP13x6c+8KDlzT/ZJCmHn9YylFlp1Ws9o6KXa2KCOqCHDugaPeQ9e+
N+1d5ZYXdvoSA5H1DDE5ERb/CyFb555ImCOd5evryqMKYy9Ud11yJGiT6XAVTPolOvua6JBQqlKj
00Ryi+MktTZiKqfr1hGEKF7Ch/13s239NrbZSM052sYTPYMI4ItQePvh9m09yZWL4ASUcn071AvH
IpSbfFF5+hr4vbP7GyRszyqhqZivfjNAxtigXH9rqjCsBPqDx56XklJP9o9uf07hbzvFWtpFjkTa
q0fxkQkc5bc7ZOWy4fEF2FfcHJuLxtlXAp6pmPcXFzqooIDSH76tzbN7QyVgQXW97d420dKAKbx2
Vyeyar63KArsm18gy/NjPgvCYd/Azl0PXCVwtGX35yYvo5551SewRA+bGw9Qgi8AjW3+M6RiGPN4
gMDN8wxxIqDk6Uf7/HuJ24JHP4NpQkfMtg/wC9hgmE79MtnQUrqzMHzzw5arC4RkFVeEuqJWNB4U
rSrMP783DaSI8uktkw9JZSaty6xYbXPx0e+pkGaUGk3tZRWflHcYfyu7sRVo8wwXWTZlQ2wioQFR
zBev72PQ7JgddKxMq4GwVTojsQUMVvhNDeB+avvVJ4HpmEeMLOsiSX4tnh6EhI5CVuWhs9tKVOQG
RugQIuZSrdNiCuuXXEPU/A7xkLqd8hlDjekPW4jnay8/dskfG1axHj8afKAN2wEKBEpYNg2MLoBX
AbkDpL0RcmX5EYWUOUd6trSYIrONXYI77M6h0NrlvtP21hq72cTgnNDtDD7lAIfz7LYc1hjM0C7+
Q5QcysIUeNSTOHgHbKmLjg4zqKXe/6uwYBmX4vCarOd2Xz9rT75kI4P3a370V8AgIKLm553B7fWp
/E94eu+svJ0BFa9NELrkmw10mPfGkr4hG2PTKqqKURbTtFBPyuaM0Xxgj5rQts6XZlFxTvArEC9I
WZNRiZX39GDPHrXxlfOYYKamcjgqN7Pg4qEbH39yNnKXpbN3dmHESNDF39Vpq48q6hxM59rbWiC2
wY1zKjoWpF6ipvjQCIHLFENToZYCJEfpYBX663lqaajjvSwo+6p3d2R1Q6ajLZYPPUVPhxJ/VLeO
EkHbwhnlu1HC6uiNmkAUh4+lAZ24oaAnSxBrn1fcj+O932vowv21rMuCrqj7OU3iwX3ZTA41jVHw
3LiK6+mQGPN1ZZdVheJ5hlHUD2uEf+Fnkl9yjuqjO+awU83wEfs29fZ3dWg44Mh35cd4ZgXFZCD/
gmXP+TFrbysbC0t0WYQWWCUKtt/4k42vKjLg9Teok1AzETKUH7ukGp+xZNsJ4ohwO+Wjp6gmoNmy
N07HF9eeucTjA9kJshcNMA8wpRO5OhDbRFdrDOCAhNv6fCkjYl+S1QRTvUNs/pK6xxrUDuqw6eOH
Ji+15UPSmW0IwtzZr3+Og36TQjqOu6qVXEQZ0rhq3McIF0NIT+21PKfey12/uEJqURktKw+avdQj
bhGjZh9rWw7MtN0CKokxIQ0TELaXKrynIz4NwtKu3KP473LNhPyAUkdYN2+Xyv6fBCXP0flt75dJ
6jdblvn/ZGNpcgwudy+SOSXK6B6hA3MKSx2GXczaCyHiHcisHfrBaqHpC9cV8ZASL6xLsOqI5p6p
xO6bUmT05lEpP9uAdNEQN5SJTXO49jLxmPi2USdpmd2Z8OXd9N/ClJpgT2A7Pwnx9+mSRYKEsgDS
DteBcId/gaIp3g8sah0I8GxohJ8vyJt2hrFQYgXTjzpCx1NTeLEoRB3D0B4ppSV8YXrwgdHWz5I0
mx/SY8EbFzioGGDnGxe1qJcbiril4ezCxn1CNcjIhffemTkPLlDnfy5daoK3UYxEEqtGGa9foxYI
LTaBAC4WhwZZBNRMZFR8AkcrfdDhj+qCLQlY8IWt5Yiz5DB9l4q7sX2EYuS2i3a7SXRxxAgTbUx/
aB0GaZMzO1jbUV3C+vEayB3KRmzejYgWINTy0/SD1v+0p96KCnp3c1FNNm1MuZ6CWqg3s/vbC2Ry
m41SAInAa2BukerV0+kQxJt5OIjxvlNMi/5AEAYeUiUemSmDjm1OYAmaBgwZdd5gHKXzGyp99DlR
CX87Q1dbyWFUgmrqEGm4HhmfL/LgoGddqDwzNwtPu0rrTKX9IjmClBCzoOhh/L2SnzALqebtBRPx
41ys6QphV+4abC0zHXXqtzELJdITBmLkQZ9Ik9LSjYjp/4T24w7tK3iLhudHWYf4WZAitC4pF1jv
0sO9xlcbK7B9IxOummZ10DOiLTsLQoGmPxy5yitYps517jG8Mo0MaZuzBStDB90RXBcF2/edwJS2
bIvYFhK09QH526CxIlkprBA3fgd+hmIZnJU4F0Rf9LxNAmDhVuuHAt8RnjttZkvF2AletHIC59vI
2/atpYScCIrj+JpzHDI7XqLCGaVMYjxcaEZjKPcR2RpAqqE6G1oqfoQpkQKk8+G87WbmJtXL7Wzw
5wke/TPrpw1bPKuwr71cxd/oE7nFhwpbzrw/2xk3D9Lb9g6QaFZ00OZmDS8ex9pRA4vmqsXsrKRZ
Vx8AjeDu1pBQiacNAiPRWJvw6L5ekcn1ENOvH2VQp+atMjtVXITIwlqku3mp7xekilmeOnis+8c3
kKmgPMLOUqAuxsD1KomyXlab4cM91TBtEb/JaWzOjf1pbMWbR5DPnkjvb7E/dKiJBnvqOtgPVlUP
Gn5cPWckWeinTJnxwHvvfDb1eTwkIwXnGUhFTXzMREP8GOqg7mseicOvSNtmevz/V9A9fWFjvlZe
ym4CFA8bASZtqPl8zrQ+xCqBreS+okrTWAsQaddHIg5KYxmuWX7todZTERu+bHDxXZlItYYf7HdT
OwgIHRbn1rdXBEqIOHhI+eKcCcXAeIGAhTtfNDWqwiejZJxyQWCMzWP1FQC84krDkZzgXjJJfki0
wS5lZnj9f5IMGl9KEvjJPzMpH/BR2z84eoWU0z2T9yreuBXRlczKk3fizPWOHzSEbYDbhImeji0l
ccTm/LevWphYDXx0m5ewXCXzK8vaPaW4YSffXcI+GGAZUknUSaT+BGUeZeMfnSteD40vnCql3dPy
n3SwNZOBeETAG37nHRXfHAlTUOxBqMboCAIzVLmjvUSVvZYmygxMpmpcKiUtxqeRwjlHtFbJZj2p
eoKkcGa2iArgvmlhjLLX6VuMMcTcFvoU2vw7l3xr9aQYgQfWCvBR+JDV4lIrq+owNm/vDopyp81Y
9PWh1eBHJAKSzDdQUpzArELbcU8JVXChHfKhH/HV1CDkIx+xG5Ica47BIEGILyLxbpzqrIHhfMl+
FMLNfx2Bdt57Iv1C/71GmlDtTRmvztIRmGpa7c3ujRafn8BweESXcKyhcz9dF+FYBbeEgITGMd7A
FjDVmcJTivLQxhRcUBanMjrdkEEtNoyRNGsDflvP/jeePupvYUz0rpMGTBJWUiSJsKcPYvxaYPZ1
IrnYQh8sfOnq6z3jQcnouwdtl+fKighDYuTloP5+iSCEp+2cwT0tV/l2JkOpg12ORTnpKhDAjZH5
03GxfPdZr2sBbUSl2xmTaIM10YHUMpmi7Gr5stn/3CWgob+oz+yHIHmBBKRgtuTrvikd0DmOtmae
18OR+N1P0B46HbKGKONS32BgOjJ7HVkznkiKp+zdDBdPEkb08WXizOz9k1aGY0kPJR31Mt7MQ+PV
gs3w54OpVNiG1vJeqJgtJOrWOIrXAwG5DnRKbTWuKYwYQdMNMv+qOGN162BpXhFpz+dX5U4XZElE
5h4PDDiHqtsfMVRktPlfpurnjng8nhuPB0ycvNyjd27wVlwSCmNjGq/14StvzO45BFKvZ0uo6djk
67Dpamt/njc9SEvFHaw6qeaVh/vM0i9r6z73onNYLFdEezv7455Rx1m6rwmd8gxYEsLGs942szao
VEjKLrfv0JYC+OOYaC8CM4kA+jQIHKlobWkYogyADYgdEIxVFMPHp57/SqzBCb2p5uXKhc+v+xal
d4P1zwJXh0GHCPjt2A+LbtIfSx4G/U0vPcbhwFvJSRAbWhZxd7gSXeCYF/DjTwzIlC7fiBYr/Dtb
SNTjRO1XfWL5rrORXz4tpeKyhKvavhpUUpcP87lqm3i1zcI8AoBNdA+AfG77pcJ+OpYIACy7R5bL
f+ciPZ0kfKoTyU/fgwvPvgnCEsMcwFfzy1QhHQQ2Bq4PmbTjYf/Bph9v1HxFulSwQako3+Ht4WMw
AG3OC8YBdrB5Q//Fmo/19Jg5AcDMM9TwgzmgC/qz2yshszYEs+EU64BLzWk7e4yX6EZ6vHKUKtQU
pdK4hrzX8Sl4Aaeyon1gxhnYd1LxAZGiTpGCNle2tqmhiiNPCN7dy/Kr+XzRY9TOdeDfMK0aK0lw
S3fX1Rasr5NNZFy3iLNOOiSzAP71RvGdDUGLX9cQdVHH5MqX/ZJc//jpgNXIVOgzmesrYPIaZ8Nw
KUeNhY6frSsGBBSPAYMUevUD7Zx59M/ieFv602FBxdqanqsubycoPYw+LIRFB8kU1ibk9wa13HrJ
wBYecgkWat9z/YDkfXGPy7+DCuZw2y0uq5nxYus7qgN3im3Q2vuPrdam36uZoTx0Nxj4EjFCMNWC
Xx/9hqh1y53uAO61DUBdfJeSVDaKyUge75BdOkfHrTTuCcTIR4JivGJCDWPN1flkx+B30mIyPNBB
oWwRoDId5YzgnUjKvvKbid9AXa8rPSkmu2+whTXjkPRri4scemFaXLfLitjQjpBMapmXYiuE5h6Y
zg/xvB7nKuOT7NGgzIBREcv/K8v8L3cWq6Lok2QGwUXngxJ/gm92p0TW9s24YpI8HTCd3J3QOAEq
BZ5HuwzbR4bzM2gEMohGBM3ywR/amnAKZay7TS8AAakjWxTyZb5Dz5wPInMwPxH4F/hckdmtX+Mb
Gp0RRrNaAsCHk3NELTbinUDM1mmYBJdiG6TKrn9+yOMRKO3nJbAwW/Vf4jgn3m/aSwbgK7O3hYC1
kYsMRC3SAc4FHNQPogDTaUgkWQ0XeuuIvgSfjcFPKiuSMdZCJ2sL2MvI6CgfbE6naH5IPGNUYn5e
LPE7gEl77eqGj889brltjttnzg5TJch9+4qm5H7c74sWeezUtFgZkxMmkF4QaZIOD0hxskUQCNMP
+nDg6SZFzu4Etlj1njzAPhzkaQnkkaLV3qUGZKtqENqhB/jxa+atCmuRV1jby/g/7iZ5UCuw5hlH
wMi5EMsFpLzUiu+nRhUljZ94Lx6YfPMYCyUC35oog9jCUl/oQapJ8s85E0bsdmfbayOwqjqnol/z
aanQVty3A+YSDXQDZuzo9Qn+LF/vmr4P/+AilfqXxgAPvhoQ5KVz2Z261YpfKkjl+UQCTj6/9qZh
PfzWmIhewkkv/mTyAR+qYQbo6KPX34Q9XpPYb2dCq+qNuA2YCQCOA4HY3+0g/lqbXBFefXKpvjFG
70Ri6DkaqZxx96ZCsXSHiLAn65Yi+Gy0+BdL2w+I8QT1Qt5G9ViijvBHJXGp68hwPByodMVVgvdS
ePldfUTVNsT5/3bS/N5Dp9PRuoxjW2BCV0tXjlqysrLiILPfPeDoZMGfeFv58nX9xKPRauq8VtaU
Mj/XzyObA/PvJjYDNwWmdLHQZW2pveZ/JVZOqozNfK6GIG8xlNc8hYtkZoHMEisN1VP4tSfhJA4c
JS0vtqISRQkAcNmSLmsLGD1JLM1xQLpnvsJyHlJY+84z3bfWN6Ap9JnTzcI3D7s1Yyxc/p5H/9tu
04/uo7FcF4DcKVwAQdmhAOJzSXKN/XAJ70k4T6vrJdLwfU5t1BecmrwRqHYp/IEgIMkBiTjO10gw
d67TczuD2s6hKnUbZzVuNhQwN1FJT2cbfNdLPkumLCUZvqaGUCgHM+w1xsfft+gKHapKGRzZAUhz
o3FxegiCOnH/2oi5ioOZRS7fKV1ajLika+mqxVnF8Hqfz9j3rd+NBqYd5fC9fmfpTdAl0QWtZlLr
wjnVxwOk8MBGgTWy4SZTKUZqQIa58UN40WQzB5/5hdUCCowD0iJnrfxUtG34bAEZQ5W7QyQs5qG8
2sdlS775ZeuC6vWZX9280MiWSpohm0KIjL5BEM7S0NeIU9PGxpC1xURck8gZp1tQgCmbcGPc6bWx
O+i9OtUvGZxwwa+dcZTet2tYrjg7Mcna1nD69Lsf7cYGvj0BBVvFbgP0FXFZFFRk2HsqRjTgb9sZ
j7WJVcp1FYi717ndrMveCR7217M/lz7ixoRXMDEuY0Y87rSkdy1qpw+kyvVX/8jMNawTjRg52fuI
jvNoZje0GscZhlFvecwFr+k5lwfRrIade9lV+jkbN9qVeJvyYq4N56867c1ke9tQfYeXJeVNFaa+
oIxeIYldsOe51u1Cds8Hkd5s/ve6RuGxQ6GiTrjKnNuxPfEeXW+xPtDPkiZXAc/8ysOqz9gyMVix
Fj3/a+vhRSaxKiXkQKH8TmR36SJSBm1UQrZi5ARvmEtq8NuuW6FiNYooha1jknYJCoGAAd8W+pAK
j4qrHCEIK2yz9rI6jfZIwTVFZw0aN7nxx4co34ZzNmVGB0yOOQtp08qlpGXas3E+zGyCzueP7MZ1
yNvfK0G+Q0g7W2MyFJHBBd9v6gtK+RxJ2sPEQz4Y++m/X7Lv2MidQJE50D1cUh2gXJxDv1sGCVr/
ZX9VaIio+v5MRj2tmHgoeDW5UihQbs06ucbyu4n2i2VKbtoZZtYTQK2S8rNDHwXtvxHalxpMZwFD
eyGiYTSq9KXQ7GpRQtaKfeb9LwreFzIZbSbHoN7lj6rSfjg05MthSWQ65j8B6PMFCSKBsZWpNeuW
PlmjGuBi0E5O8QKRhIamuMalstyF/0iZHpd48oL37cUOiqAuROQ0rzze6rTv9ZbvrzoeBQAMYTSz
c1wdFqlW+/QbXdmFcfqQ1dEsfFQhYEsIRVNkHKGy2+qI/D3eHqEtnJ2zZG1VoWgZKUenFZCVlFfo
on2qJ+ohl9JpA7prOYXn+CekoeywgrPVu914ooTelIJezc+Zwk/o4rtmi4Ufb/4mSJEyc6EhliCp
oGeSzaNzjPR+1lG2W5Br0aRb8CwSCGdBcI5wYoo4Bjrh0n7S08591nt+s/Vn8L4j6zIFhL5RB/mt
KgGIBQ7e0WiHo9ePNbOlcWsDj0wTqSSkYbOEQ9ndWdjuj4yi+RS4ajC5u9C4RZblSpR/kUG0oPJi
2UN2rTgAB2cHweWjkQ6PUsU6oVcuDpz7mIXlQIpPS8VepEgQvcFcA1+bSUou3ttjfT+PvSvLReXB
B43eBngmiJLerLqWJEjWnV2yCNcF2byXvFElcbCMepaYGtBOaxDbqdcXhoONKJHnNoXiBgwRr7qs
pRzWNiFT/gnYFf9ao+tqOFfr40o6H4S6/kKW8y9y0kxW+QuFU3iFzNfuiHySHpJr0iEndF+bCNyZ
RAVyDk7B46W3drLl3EUavSzWaUgv1gO60kFiQnuvptWNQC0HKEM5a+1cpAVQzQDt49MXx/WF+8VW
nbSCPMZ5+ihBuiOZM7ZYjmg8+w4pRnEwhNZSofS3VBcAT9nw5UyG4x11ip9c21hbZ+/HqPSc6Q9q
SFhB65eh572I7gRkPNE9z0NxnXgUvlDykFOLjxJt2YhEbmTHx80kR0h2fzey/VD7pjdWTYMgx+Kr
9wvdXA9YR98Mkhe0xt1lwoY3dfOtrqZnyGow5VhhW2UBX0+lzw3GxIYO8pKGhJKD9goBSrZ4F1Kb
milnkRhZBk/Cgf7HyQhCfpRvberr7pgdd5fOIVI70NBiDIRmWEOr4318UkHal54cKgad18ZSl0gg
o5gKZKug3szVjWnJFN46yGMBIHKb1OHbyw9P7mFOE0FS7F6N05c0VckC84lhzQFCGLbvJVkQB+ge
8DEAHzS/U2MJ/Nm0lqjkYRMPO4A6Tq24NeqnR6DdcVbKheyDlXZFh2yxhqJ2I3camiu+ypFleaKx
GoZiKbHaHWY0C0RSGCT8OYoERfmeNU421uOm21wgqeVI3lRilnDlFHzXoMqOPm9kRChao+dvUY4/
IOqGNAXqguOjiOtbt+hfWtQp+VxpiGmOMS+WGJskEFv8R/KOCzOTCts1vEqFsQQknNDVC1Ou1P2a
XS04QilgTzsLmRQEV0xCd+fZY0fxbcQzeQtuzPfqyaYj0seFgN4AyJqvheYOdxaiX+/coYmbJto9
vp/941SuxANq1rHcad8mxyTLuEv0/tF4yFMC3TToIESEAq3FcP5IPqHkMKmCRQtDd4TbJU85nGW/
s4pFCI5Ggl+xuO8DXI/9A/Bcp/ZagwoykBZN08XiAzSkaDUs1O+CzPWwKizztuWZ9yuwsU1JZjy3
owGnlu/ZVGlmCI/CsWklDj0rPGmkLcQhlWDF6wMZhYf+PyD03GJMYilRDjr3ROg00OVmM+axtB/S
f+2DH1f3jt+jFIF+C8XiPYo/FiIHC0CiQbWxYs1seKJ7PQfmHXOV6FUakMNOCiHlkYzgnqYsNavW
InbyVdMLltSiwm1+WwyifRDj/Tt6vfNFj+jCB84Juz3BhjxC7UnMpvvng6fdepofll5eD+F4y/SS
VJpxfnc7bo4W+vy7mshEqTgKNku0yPWKsFNaWjyVjP8fVLoXG+W2py7GwmjF856Gff/kPreoYgp6
rDsxhI0LAvhAUFzKDh3y/H4/cok+AlfKmRjBqbelX5jL3k1o/ypigK8SJaRV15KeYbNPt2caY6ld
9ty/i0IfyywRZaipsErFBJjnqXIHTRlgYKisqY1nbyZcUfXiRzlfG54UpLW77gaMCHLjf4dQjyqP
BxnG2s02AGfa5GAD17yuEpbyJJMLFSXOHjteUNkRdL86tqRQvE8qK1X31xAPM+0QEKuoYsiooWHs
bOxagKAw5bcAftI4OBT6xqWQ7948ZWV+vkWN74RdAdyc8qAV4n9tBotoTFqLFkrfe0kdqMf3GrvA
NVtMKBpECSNprm4NrZW69HyGqvRs9sz3j3QFPVa4kHd28+ewlmTKI1+ksbpxkvQUhCp1n0k/CizT
8I2rTX5NssIo0kia+44WtdUdaRntZy+kYA3FGqaTy2Y71goHR6PrU4xh/rVcoi5/v4T4DGen52V1
kNsBNiqI2jsXTdlGekR5EyhPGIhnrDFeLpUTiNJMBjXFUk+plX3LvCm/fE7OryCsCcryDAceQ6jV
mM389e2tANe7oKt373QE17AEGEknfdS3Oo78JQPyMR/959jyUn2XMyL7BVDfO9fRcfgl6HD4xuVZ
siYZt5biRkjxJBiVZgW3EU7PD4vtsatZ/YlDvbf8MS979bGhGW+cxk09fusptCf7x2r69i4SgtWp
COBaxQuLdx357DgK0iDw6sDW/NNXYyLlFvhbU6PQupx1M2urci3YfqrlFQwpGqRQxlUNsqTwPWGc
nhUADL3UCh0GUfyCuBOBsg0bTlnSlP+9wqESEp3DHiU/W7h36r9ifRHc8Sxw6Mp/8FiwBGiwdqj3
ZVggtHZLh1uQjKNdTb5c4UjJT9glzd2uYVP1flEstvsgbZJPmIr4jjok+UdGF7y0r/MFDNKsGfSf
sI5Hxu/OA2mM50rPAutYu6a84R3tPFH9HR1I/e2mbQ+LaW1BWsyHpE04JSca1no5sOdiXyuDUquv
xdPZzwlXmtdWYpu6bcFkNp8TdnkXqajfuh2ORDUfjdyGI/jU5P2oIK86eM0dDIGGbYnoi3rw2/Jl
J4XsgD568LGyUQQnus3ZUl9Ted7KgT2qoUzKJr7Q8AfIKQzmg+ZJm7YkbvkWKq/3RO0GWlAK88w7
9nOKS2mfhMk3+Uvg50TAaF3jQtN2wNtm1L/DJhh3Qi6kw6Yk2jQFKhgqdiSbo8JdWRh5TIQ62liK
skkguE1OaXd2OU6RDZbjiAxnceE/uTd17fz/BcgB2/WDrS9JRd2RTE09T/mxV4cGUaUCalW/l4IX
fSpAjSAKVi/PaBnuE9TEL9K50mQPx5mChjytKM+GkodK9WbYQRZvO6q8RCVNi4N64Ez7wcbCKhLf
YUm4ezxxesT5wkViywvEXhvxysaPqisHM7NKA61pROYpRlZVpp+IhpepO/RvX9Y24vWVOmlFO9vH
1h/3xytP6zOdQ54SdldpBAAmlcKt8G7EE8q5c5NhX3oL4BQowIBXPltiLgx1vIWFohKLiTDMVgzk
VrHEHMhUDTQVdYHNmggtjW3WL8+bJcjmIh3nCJNKdAZQJkIfb/m/CYudl6LQ73D1jqna8aG2EOWi
uAZwdaeEYa09h63sggVSTDOUw5uXIBE/i0IXqSzDxqi1SshwWkVleTaKCktyPQIdPkZDL/uwEYgQ
kp/roG01fSwIx+73xcMFxCEvhYXfQbly6VfuopLqqkTaNX+0JZqtvDqULmaIQXd1ZzyzwCq/h9w3
24dgbhXHFpJimVX8SzcyFmX6wJJsM/XH5N7/QpCFUMZWNjSCErAgmxlmFeaucgoHcdJts492JiJO
XwsmvZkP72iH3tQE46o7Z2JSluuwF7gP/wrG61q1a0CTig8Kh/HsiybVbWEj9Q5bqK9jKyTKZ/ne
AKW6VnAEKT4qZqU3FHlbvz0ZcaqtpUXv0GbNq73F7jj1vg0Bpvqecg1xd8KQUk61nCtcN/xXKk4W
PUqf+LNQJMoCsqMzfas2JgV75PHKVo4szUyGEiuhPogBvyXzV8ooIPcRjZ5MaxoRt/10Nv4HRWcm
Bvht9Ss7g/UkNU89O8VAsN9pUp+jinP6xT/l/Y7Efw3rYhuIFrsa1cn+14s1BHlHbmhoXwiDaQTZ
QtKZ5HWtfwkORKyz2x4TFP02ge4ewcgF/XXX9+O8KPJOaE1zEBklDLXpJUQLuO+WVbfYS9c3xOey
bMFC8g/yoZBRa7igf+wKpKtc93/QC/SLUgTL7y/KR5EtPpXZo4rmo+sAbeFIXxFJUUtPF7PsPHya
dIDa48pCkNRCeni9oAVYSY7qYFPUfh7skCZQvDdTMnNUbocgBLIAgSe0fxkyb4giILU/hXSyANnu
MlGTs0q3WEQYO6Cz6D1+7GZG+ctI8HgpNZr0EmtgRVc3VRtldR9OAFux27nRoQvLsVikTqJ37cBq
i2kqTbalBAebCdDDtmzO8FwdcF/1+je9FXzGGWkO/Q/BjEMXU8D3rg5Ivilx+ClX0c/R7aTI9qvr
+I9DBcRkbOTgmZkBptbpL3UwUhxIHW8G7wyfCk9/inu8TQViaTU32KgtKTmZga2AeUfRS/8ruLk6
Xv+EE1BZR7WIdAlqHZhacIDZhJV5tWtrqnXTY6FzYjYV0+n3iMx7LmyKNfu5z3ROBguarZ7hg1ce
J7nntF6v5tzG0I9wAI3QAWaQEX5qUI/zULKTuXHIJDfGWGp0DfYtXRz4yTLbE+ut8acujd9my+cd
lU3Y5C++JyW61sUWXCUfGiuugY+kY+iFHPN4Yn08ErZeD9P3dhTiPMdRmgy9zXP66FAykSDSCg4d
DcW/7sgIKjJdViK3vlj/KMeSZ83ewTk/EdRcTT70VyhlL8FF8mfurL3r4n9pNuDbfUF4R/VCKjSg
V9E25hhQ93r5JR13u4HL4liOyzgGkgJhKGYVVlUL45xih2wJsPZtPnBeu5nCQnJmDPGbMgkgBjug
pT4KtBkTav5zLrTyRI53/wouoUdKFzJCs5D2ghSuieId1MC6JjKmrY6irzDMz9kXV5puJ01foqOI
ksZ7jme3/9VbtGjbEFV70bAsYUgA2z9q0YD+2SYsnh2H2Jq6xb+e/df2XUUKYBcRUzESpkx04ci6
ghgB1VJ32cLu89BJJlbjrayaNwm7vgiv7VCTxVbPBl5P/er7eJJ4OeleL/5wOPQyUzu2+pZYPHuq
khwow0a0y2CPaPCUdMsDTeVbCuYGMkmnR1DkDSroLlKDavatxMJ89vIAynlREbzcfdDThTwZaw4x
jPAI3hrmaDr04Xp7qg4IuMQkbJm+ShhIl8Ih+/FX/iORHfIkuJ618nUUInsVQsBYDkHN9bkviZe+
ggHIxe05QWy6c9CdzeGy3EhChRI7cJCbhu3Yf4FSIIFo4kpOjLbjcOMix9qiQGST7cgb3eciLTNh
7am/gIG1+ulQNQ4u/MBzCVgDdGj+TmXEsJtk8dgl34O5/dkDWqzOhIupL7ufCKi4P/4uESodZre2
b2ezKwN7cuaj8LHTaTQHTduFKnWfLLmY5Ze+wzLKmaFtDdVS7uBRUQ65WVYaew45X9ZG9qDhCPMe
39RYuKOtZxZmiTLO1F2Is8x3DeUTPTutKX59xZba7sqFDX3ssuzD/AXs+1NHRFtL4CW7g/VpT6F0
toAk3Od2vl1LEHVwKDWL3Awjf8Z1VNLYq3p+R0NOFkuOoTycA85UTFaY1eXtNw7lIvYI17/cXM6t
GtPUIpgeJ/VHnhVuxHCOm6Ijk3DkVuGX6SxSe4JjFBK9WxmpKqrkUtKiXBOPdH4vYFec3NtUabSX
EWgWdFvzeBaCeifs2BNGc9xKVaaHLIaVDNLuFxx/WsoUFD7cE50WHjTMlDrfHuYn14bqjCf/Vo7W
LkTzR7jQEgtlvAZ8zySD7u01yECZbU0Na2liPwC+toeS8BYEVsHmXgR8UUqdssBcUPj1X2DxxwoY
ehkldN5pb66iadmNHISzyCKPHhZKRLRUeqTbX2pp7np0Lw8W3In3Ox+2PB6TJE+9Esmrq8Bw6moA
0aywvg8XZnsGTGTdmxe9p7X6xAS6Xrol8v5rm4vqcMPrPIdmvLnWq0pXKZ/i6Jj0DLqr7rxUkywL
4t5yk90AIlie2Ul4LCUupCLoWbcEV8pTv0fiZWaDFhe4RU+vzKhIv6kn1/IVa3CnnGU16eTTBzHZ
4HF9GOwatIKwiFepqJKXsDiGBza72YP2Q5WyOSKBelCVW3ic6lcMleLkXMYnn2rjpCpcWEjMIBwZ
i1dVqT4x+/l3otF0f1yWfTtRH+br+/OLZJnRYfsCz43vJKlXuDS7AC5Z3u8SwkleypTGpbUxzhK1
K+gX/xcYf9kvpTXGysH1BBEd0T8lVZNZGHkmeoIY9+htPuBilZTJVOdeS99AHeOD0DNI4epDJkaG
QVUn7QpmisA1a31sjLKZ8OJUOk6Z+qbef37jgl0Z7rUBTAnK4WYbKjmLP1FEHtv24GLbED4FULg0
OBMt+yAloNgb4u6+Z4WprnpASscZyiOV9NJsB2+3yrXTfzXl3X7DlwZ6OpXZwUw4jO7zYXxeKyTU
CM+v2efUgbLw1lbQKPejdpqEFbYfa3KvVaLPuEQU90GIWn/yOMFMss7J//XePta1f587WHnfdXQu
ycKRIIv8DrBIMjBvNduVNVA1HDva+k/OtHdZJ/3xhPEFifHhPPwM5U2yllTpQTgE/ySid5ICVcv2
vVujHECgaNVWmTGqKMXTJ9IaHKgxEGf4FwTPEBoL9HLzcH7Q0Gde81tcVHTjI4gHc89plYeBP57/
nCDhpLrWuPuh9EWWpABclRj88M3mKfzLxb+nnsLKVqlOjZEA5qLgl+Nrj300b1N8kKcvivgnvGYO
aTDwXHAJxMJ4J0NSTVYvtEXPdQVCGByrk08wsA5CFryWGiMTKv1Un3VGxfFRGaXGuP5EWj5+u0RV
eBhJZE8rk+zyAac3AeMrhWSENaTFtDZbk54qlpomfwuGoehsV4HhER2rsMlFzxt6FYeyHEk9nOFm
EfTy5qb3fId6CVoJ/VaZtCy+qLZ7vVmWPhDqcJrm2+6v1HJ7O6Cz9v2ALh3C1iWjDkadsAiEZjsp
QOkgDTMyI/odI/TprFpzFKSydoORoUdin3qKwSGaJfe3kzCpdrDeXVqfH1+vwiBauO0EOsSsLi03
hPpxVOuXHmYoRSB66micuMPlaDFZdAYK23+jU1a9JZzLp95Pd+BFjtsArFzmo8oCYhUuDJ1w7pJ9
FtSP/pY9a5Tf2h03xx/umMpdLPlY+7iMtWSu02lGFvDdOAoTb9PHnelnq/BDhs3RmYHfCO6kqfxc
GSRD9Dz0E2ScYShIWiwyOBSFNpSl5xXnEaVPUkT/qEGMfZzlv4RdeK8yhN7LxGr0zvGHcX1P3JXo
Hu40nswmflpq/ukU0+CjU0fMEgV7YDnSPj+pnf1PWjBddHXy1zxkGJpHh9XIgaFRGnEynFO4AJX9
DYt/Rt/EAtXn+7SxXqbhV1OBJyGUZ38AKjAyqupyyDgvMY6fx9B/Xi2yG5Egy7fynOC9JfDJSzjT
sksO0lqFFjGVmxBJFuO2F/nMdnHh4wYwLn5ZMV4SgyvCvcExnuAT31/q/hHuH7chn+uOYJ3cT70y
LkvAd9xe8UCD10Ym9j3fbo5OogGQCsBcKu7NjtiyRfbHKs3loe4uWaQH4FT3aoCVmuMisFR3zIUX
b8ytMknmt9nsMc+yShwu/+3KIEJqKfOOJcqvv9ZcHOxKqKfBPjxtLGQruRoAuuZRijc7w7BveBwH
ER8s/Ve6bQQ0D19hnwlyKwNP2CqAq8yqOjLrGap3n20Az1PmBwPpG8hkaWzmp70ZIFy3nYejCUVs
0D+99VM333I3r3Jjutj82z9ceRBHAywbLClZZtzn85JTIAS3RXWpJB8rt5ts3vueP/KQeQQu6oO0
gNK8e78kGZ7amjfBUpsyCV7UeoJHAUr+4sDvF76mUiV7/G5fKBz22bosdiz/4CU30SxXODIIPG4X
3Z3Qu5fanmyK3jT0MATlHfjfYYBQwp8yd2R997jAKy9Un2WuBxT0yIGdXkgobn2NsMV/Xcio1gQj
Rm8KvP6B6EHsUPC3wrWDP/QZ/ex6tJfSBJ8jf1k51g62YG8m7Evj8t2TZKi2qlbUOpm5Xdns4iql
s/bvHEwfrdiwTSA7rqHTuNnvXkE+xjajqbBTYTf85QpLIAhKIQfyf7oz6kPz+i4Si6oVaRKJO9/0
iB0ME3wJ0Bz+ZjmDfJkiA7G/DarkbAqM0/GCjHzlZY+LZkDl+j/q40AUTNA+J1PpcLLXU7XhTzA0
w73wFOn2SMr8lvPzr1HA3KXw0B7NV8ulik0T0q+8o7+8FsSTjks/ZYEXoDMljedl0Gr/yhcV3/Kr
eysneCIQllzJNaZo7gVb8sfQoJi7oiiNRh2NpGSd0P+TxKBpuKSgTe5XtrVO0I3pHPN2sVvX+C6b
SE+a2iEi4IoWk5t0B9Zd8XbtdIL3YFbwz5Uzk+62g1XFqaiNOpVCqb94q6kJZMLUHD6J9Jc4dI+x
moSWHBMyK6wl62DLUilDPIR4m6/h5LjSyxCXbjduNh451BddIb/KoXE2L3rZ7lCKejMBv/+C4kLn
mmrczFLyfcJOKmkYN2xBGW2FZqQCDW6OZULQ4yZydWFZ0hFu6pgZyqC381gk+ZbvEm9NfSp2oYx2
UYs4klnzU4e9mq3eoff/mIayxDGCCo9erYeuLJOOeEp6j84sDz3NDl4RO0oprejQYciq1dII2Chs
fgA2p+H686keJF1GefjlklQQdYOw9uqpFs5N1O1YMISG/lOLkhloYpXc8/yV8zhNe9viYgrhUyfU
rj5B+YJA3TR8WIsdI05uNvodH/9AFe8sCEU/LmYiABkgUG97mKMQLrE69IHLtjoZYNHAmKf5OVVe
4ccQIg2pBfiru3H/7jMKXzmFywtfxHgi616FEz8A5jSOBF/QbjoIKDnRjUEEjIo9rwHX7o/33D+B
711ayKBt3AWne80mzbyW4osL3uJ2F5a9KrzpDooFClbOUalnAyVQi/Cabnbms+cVaUJuQom0xAb6
MKPEOi2+dikJf4eiqOvXYR1cWfwwCvYnijoxJuVw9g/nAO6IF9ZobacvweG8FlQL/dFCWakK3dtA
wHuTGOKuPTlj64NKrCDpCOg6km28AOVzvrbl7srFbhgSi3SaLF2JLhZo/zi2+QJpBc51JXHLST3k
Uv8QJRzb+fAiMOSKtJ/SNwoyzBP2thmNyWcphnbJdlEBZu6qC3HF/hzxQuRnSiTe38ln63j4G4c2
REdQGl5MqcXB7IfFN4oochvveSGUZbp2Cky5CBEjf3b1w7wMeNKlOTOE6Imub81oNbPB6Ee5K94y
Wp/7c7HAZIOX1bJqwr4FZlX6Uk+P8gnIvdgECi4SCC+EKi7Tg+Oq7C4Gjs/dAfferH6PwNGaM54X
7HsPsA+OcO+WgvW+XhQvo+TJ84KmlhwnAUOcnu5F2q0NPWrYiUi1XEsmCYxvh+hejqDRRXuKqNDI
zP7D50s8/y55NTIsAA4vyujOLNGNN95pkOvM+eaDd399PtejNwT64G+2ljh2Ae8oeGPdIa3mYx7r
Y5KbunclkQa9WT4n3jOUWUk8j9+gc2/2HbImA9TX2Qj9kiXvsNnRAqdHn2ccKnn3V+0bai178r9j
s1QLQ6KMOC/ttGnJeNbh1dtHRs+l4l+gghUI3eAJuj2L34a/jBvtYjcrHTcUBF/vFoiy56qaAuTR
/Ss0vjHMN58RxGBerWD3HkEAHJSDT/htTJsXzs92xCzs9DbbXQAubKaQ/YXPe6/UNXfRSBaxwVCJ
afQmsoJV/fdXgsT6erJYzrgvdXAWg4MQXe5FmYkk3PX3i9k0Bp2pwni0OHk49zBJ9g/MYKkJ+9Hk
D9g+I4m13JHGbcAy0D0yw00ReX820nsdN9utm9IrV3xd8ZudNAEyUTyfOqxCTkfoRSp/lHMuNeHT
+Pygx3mK91VpFwW9sJD+VAtNi2k2/XI1dtocRgzxBfJ9uVHrBLzmp1qo6EK1K+VOEqFgOp3B5+OH
9i0qO1SLte/Sw3EknkEJYhM370RNCzVjT5h4jva4H53mWOf9Pc8wQ0DKMNEvk3694/qT8wOC7qKy
Y+Zeo8nKOBRZaknH2G9z2rhpVerb5oINvlLmZk4Dm2Bi4B32OTIN7XWxNWW0qN5m2jGyaq/PuOjE
LGywrPKZCafsbaXyUbmCL2SJOUN35hCM0wmw9IYCLBoJpRvnqOFFIbdTazqK7dv/4eNcZuswXv4N
OLlJyqj5cOIK0eRiixS+DHUWq1kqZKXaZsUM9GD12qYB08410UspEcmzxoT+hWFZ6Dg4KdeLVbnH
qVF1VfSCMCuR3NJcAcmxdq2wTyDReRQVqgT+SBVgjx/xbpfLmANW8QD2vmmsMZ/lJCH5N+dN12VV
7NoK4WqON/srzHZOB3aGuFGnPiIGHPzOnMCAA18p53K+4qhrY3jtoWjNMXKB7K9bze2J81i33yHh
OV2050N0oKmTKzSS73p1czl9XnjkNUe+LALODxsndhGz+rnoQr56r9cDYeCvZhG5DpvfxbBLQkl3
4gupWuBRDKIcdVvndeJR6XLFP6+5UAbReTZ/YJlvrtGvcTXNIjqBr3fLBrdtskS4uQopZmKJ0Y8n
fVaOFY03yYDXaHkvr29F552eGi1+gq/LVlHjcbSCKigXqFwNsIEWxGzRY1pCYG2S+J0PVjzEj0n/
VrhIkkiYz47VNbPDhMctV+9EvqZ8cesrbJ8bap9dSqO7O3/EFg+fiibFGTlnBa1P6CON+UiLK3tk
Cjut+9BBJQFATDueXyv5IDXCKlfmDhbLQdjZYe8N6NLMcirRUG3IVRpcaOGzCTQNZ4kN3AQQMYb5
a2iT8vYI+Fck72MdwLN8WrvlmXW6heL4VzY9vI5v25O9MMfbFwVGMW6gVf4El4rMBAbKTAHuHyvH
DBMdCS0A0a+6zB8wXYzjbyTiY6GHnLI9LQwf74ArQqNUeTzoD4yaX3y36aDrKnEsx4ma9hktsLht
iRxGvO2Bi55DuQ5TDGFoBu49iliUliIs0/HwvKXIhn5cvPP4d1Q/K19knqyu3hFvj5WJDXpBk68k
ASXYNIuloFCdp7n0K7+64kj+wwKe5EM/OlEfPXtXXUWRYJG4A/OUHH5a6HIephdw23ez7Y8fXsiY
RzEvrLI3+0Cvs8H71DhKmrZMk3AAzvfUURXsoIuhCiqoFU1YvNxXQd5M7qCubnJi/eCTcvaPVLrp
attKEF2fMDVt57XAsn/rC6OK1PxzHsKvj1L4jZ2FvF8Wj6wm08LTQVeokii7d0vzjotjWgEl2fZQ
U2ltSfbzI/d80XWpwgSar6Hv2zoLvwqDeE8iqc2JO75dhDMkug8wQlJw9gGb/DLPe0M4W9GJ0rOC
HmZnToad93svZQL+VUloXWSGCQsehraf3RAXe8Mtp0xnTaFrl1EKhqsi7nYqsM5qiE38aBYp9WI/
bRWZimO5Wap1Wq72Vevt9YH8gsxS0Vgg5irxj4Q0LWQjByFqRTxFUBH6kJNEx+70cyHGNJ1N+gGL
1kl4z84H9n/WtthuDezhmP6fobapALQ53C4UlWy3j0LMuplMnDKgJlato1Am1kwhLN+xQDxLqXyW
nmSs5cWWEtBoYj63nA0kRnUhUuNG/zkuzZ2owE1v5ELFbfd2zoXPLosxo1tKH9ZWaHWxBApHr+Dj
FidrubRVTwTM7jyKh9TBhrzgsqiFKrqRZM0PwK+5R22m91/3w9F7DudTSgUofyork6dNc0BJDLVH
FYRj1ujypF7+r4YEy66FpNNw4klPyQ3lMijmT2d5PEjDRhAg3c8gEZqBnsKSKjfRhboqVc2LKu0C
5/hxxC5Gm9/3ZiurqqFJeMiYaExTN4CCim/xVXPzHPDm4paXz3vMV1f79hhiTbMCJ3pP1NUf+YI3
vyovLbhgHHynYuXL0NyUKicJNRoTQtpCN3/TRVLVkj9TBEbHVsAxkT/fc1WlbFlm4KDrsfq+FVF4
AeSosazt6YwqLF2AWyX3iMCDvh9mu59hetH+FiWeEjrEuZuQ45VAYAB9BIyhpsCV+7y9QsEkv0i0
LAPsLZluN67E3+3+mjUNMEPYqCnLGO2N7VwU9BIWEMCu1KDcZRYdGyMEvePAvurjeuFMq7LFs4ro
CLb0HKoWpgm81b//K0JayGRqkb1DquBfGO6BPAKeew6jd9VLFeorBtVqLu3pXgvqyr6rW5vUb8H4
Dg09B2sECwAV7jz46TpGXtXCBriYLCSP+ykBHtp8oLp9Yl7BGm7oV2in5llham3FRklvz9EcZLRL
lR+Uk7PhUrR9Jsmnj0dIIN3aXgLtzzbP2Td/QEc/71is5T4KN+Aby97gnBSFQ+1yLC6YSzAvw54N
zIh8RMqEUvw1Zimhza18ZpMG/dzIBj9sYQMnhoLIjFLrvGPxP+365a+SAdPxkRq58L/rvDIIhzPd
jjjsHBVZrmBctXX++p/JwvBJqJxQBcsd0rFN6a05NT940lwU90fdKToeLbfh0hqNNTWBSsegv4G1
8kg/dMJWxKWG2nI5p2pA81i0Mw5B37L/74TlT038W3NcHAUVBdSbFisxKHP3O67P7rS0ykvCS7C0
ERP5ax/ksLWIV+/oYKL+RkjlufijOZx3OIKjwoQsU3F0athEiCtWR5j/2hZU6sb8N9EMKOV7OaCZ
gr0v9RZz75Gx1SJ3pkdIWGGWzwgI9zLwOBf0WSlY0S2HDzw9ML0YnjbW/P1L6IwO+psY3avL5msn
Gmt9qtkPY5LU6Yx01S7sR16rMHAJKVCyt4aKc//Rem3eM9hGJynTBB5sji0Nz6C5HzKqZ5EVTq22
HMQZaPcC5VdgiHFkFfxm39F41fr+HEOWyLmdAILM2gvyGeM3FnGaoz8EnqAGtENfRd/enBNFoLy6
BS+KZUZ09djZwj9LeNMnymDutMilTNZqH3hZ9g6JiRsTlkSVoqb1epR1c4k474+8+oG0Pn5VHzOx
7MZFDSU+qax+SNI/MJKUBsfn4DQ2ZmOyrXXIugVMBRrnzc87rKxLWtGbwrVxpBo3JLwk7N/gssap
DZ7cmopLxF/cz9cLbezE2Wf85xeEqDWRQg5ZhMDOuJjPiDkmOwqKyLHSlUQQkQ8USNUA4fPWgsIA
dteDAc/CcYYdp4Qa1RPq5q58et7Xj/ddCVwttfucJgZuNXkBrW0RKm9KF6YV7uM8VTmZeGUSmK79
q6CB1NLGHrpFyRvXyza+BNoRQ7rqBxCcP4nrnofYVoQ1da3JAkx8Q7pgyUqGexQn4xNhGO68P+Ok
dkWaO5G7nk6wcpKiliqbDtGYhR7lqK32nhCNCCyJn3reIst7jtrgkg5+8+r71XdUwhZZmcfubnvc
98LrpCgxNYf9KgcR0ynEsXOQ+lYQUyftwvmnbCbHzP7h5qFDOjecfvVYixuayVjX0ksKu5+LtI8R
a1xrTaRsogkTUvW/w+uBjhkOFGOQUVAbQNBYnGUNPQltNCDpGR8vNTfUjD4+PjfcxkmhxSERkgd/
/gkC1BJ+GClFkoOhn9DzxK+33XVktBV6X0cpQYvOccLliizh0YV+UL3SrTJtVCHG6fqwepp/CslI
uHfQYLCUHh6MGTYIopogW4dWjrtmV5j5swbRHwzNDjFRrtSfthnjPRY+EpRlM2lZZkwgeApL+Z92
yquNkjycOi7kAiCI8qktAfT9QeXVuGyZzjqQ9sxHZz3VC86tk0qDcoqJx+ebWU2GaKxW0SvDiI1t
9OMKuIUQQ3CHkdAnjKwBWESwxfK/L6HSkVrFXEAxD5IZ4itHJfSVP0xuwK+KqswNYivId8ZwJ5OV
VHI1fEoQ3hducezB1MXR/zfyW34BzKuNzZ6yZgDXTHOrRQDkolQbG9eNrewThlQ6jlXNv8B+uXnF
A3WIwOEvuD90ayDTCBpTET4MBLQWlaJa05g4PLKn8zL5Om19lyLeQNSHhKtKUQGaOf6SmPPZUkkH
qc5Eivprhi6zdFlSLHrTxpkAuwgwkl6UReK+jU785TnRaRoLJFI2wWVpPPZTf5nVaKpxwu+LHHpp
vpKSw4HlpQ2DWkY3eEg+CNdsPMSQ+p5VTrj29D8SX4K1MGBQAK/QxYMNdd/CQ506sN3RrC5ZDRHa
2HohqjRDM3zSY5RGA86i0WgY9Tzo7bRMuQ8PGJULWdi77sLG3D4ZJE3XYYM573y9+slZx225Osjp
bPXPNJu1Fvq43PX4TS+0YXojkhHsM/jJgjDpKSJu6POV6fpSt+LEnItihw7tPrMqoR7Jbwa4Az9C
GIwuVY4qXyVv389/Di7PQSouQYgAOX7tIO9tvUW8rIT9DM8P+tZzGKEh7/riZK47vzo1WEO3jMGh
ixgeCudsRQpRoqM9RUC+8LMpG0AJM1Iuut4XQrm0v8DCSBiWKACYyoYhZQGGE35/bnkXnTCbdgyl
jCC5cd4tf4M32P4ViFbYM+hgBiPAhmKyDCOpyFUT/BhCfWbSExyl923w07ZAhWOccHARcxV0wx+I
DPpOSvcJe/a4l+Bb24bgWe1tEBwq7WeZu6dIwxGGpIAFl2BVAXP6AP4iyR8Lxa8OoQVcMZ7rjoRk
dc4LC5ssFVQAcAAaL2FoKbjMTYVuZiFI9lXqyZ5QnFRpC3B7Us2IEA/EWJzIa6eaiyO904+y0a4G
pAnrS+girXD7kP1gcBdyky+HRhPQpXJAv0SjezAKn8Ptdq2muvMOM7aNusqGx1CvCQGbv5x7Id5N
pv9PEoRmVuMY2xuYCbfoGqey1rDCg9iDTlhEw1YBh6/dHBD8gSwLZLd1LyE3WGW5x6dM6wUjmMiX
4AyN58BtRDo7xpox/zk08hEnK8/BSIx37j+BbMM1FOWwKl2SY9LB5DWjkKA6NLL9oUILQIs4xp3W
81+gUX824wcXWlHOVKz7gg2NkP1uqr5R5vWmDdtPtK2YMWfpeaw1BtzEZ3YvQ3XRzyBDBmFVAPAG
nnT3Ky7pD4Q/nxeSnUQsEYPoVxbVZhz+/T6CVPlPbTMX95/BfAsXf7meh1q5ndRxGBmOZXwTHLyX
lg+1VDhbuLQFcpVd5nhH1bGofK22yVPe/omVAxA7nucpzuqIe+NZf8YxuNo9pwKcixpLe04r8zn6
sxWcGcVISSCodyXnxekZiBFbp8SBmeQWPRt06aagU7krwD/wEXe9H+ZpkB3GQM2voVW/KtVwlKhz
YT7lTcNe+VVvVbAhFhw10f4GFE2gPXwsu5xRsYQ+8cEDQvt3Q0tzgftqKlGRxo7aamOnez6m0BLi
RUOCawAItZjzZa01nstiXiXD2OPfVqJiNruGotCc0NYw3Te2N1u82sLOJIeFngmsS7EvI5dSxqRE
xlJkYwtdkSQb9IHeFcsqqHk7dsr+i/Xwz6Vx1p0sJ1X2649X9+xvHT/kM5LUNr0T/ubnRsvFsVU2
UXPy7QJRIeVjx0daUmEULX3mCGxKoijFjuzuMe1+0YSH8i8u5JYmdP0xFjYgyOt6G3h2HAHuDg3n
kPBHNPKGHe7UGyx6f16L4LGc+DWeVXfwQ+T8zXJDkr5fmpZLsShzOTAQPTGwxrX1F47+mV1htLcN
nHPi6DbBqQTRwh1RucOTaekPncAyX1njz4aWeyVjQPTpQFScspshILI1Q4yVzbh3MVRxk9QcRF8P
YafUO2gH6+lTNZBMt3+OeArLn3ThZcKDrZH3cljNqeWA/Y+o41aYS03T/fRFM8cPM7ykTCCmc8D0
nIt9ZqD62nyGz6P5mcomkkCae0vdidIOdFo/e3MJT1o0a1dxm2Bt1t+NHP+kKblMAjea19AoNV/k
5DT4BYPB4v2VyPHs3IKiJukHswzDqJ01x10I67h8v6V//jHw3eRmCzvUuq01zk9K8yKS1jlLNAzO
Z9pA7uNK2WqIbS/dGA/t153WrIBDSARdq1yu47vZnAXVnjIlf6H2mFUI5iQO8SGa4+Tzty5u2qzC
XhuvkSH2JxjTS3eHQj8rdh/sqVlqLk5HWNxxrpAdBB+nKBMt0n4/KHDzCqtKX3YcvhApqFDSCEF8
cqBEZeKlYPw77o391OQCupuITo32aDXXcd7rvES2IKWz7nNY3Vuz+DkW7lDIHRuau5jdWxTXKVdD
i/V7Sl5dJNHtWP0Ku5k+5E2l7UcMhg2r5SB1nAXbaB1OQHtYnDd7MWJuCWaEvhxLgUNdZE3wLE47
QXcRkX48O06Lkx9/p42INzydLlw+J8D7kt9jIzDUW2M7PTUofwTuhI5PANpGZKOmU7oKqQD2FfOb
kair3oG9QZ/ydi4G6CS9FSpvUBlnGL04fl7zdxCka+TRxrcI5Pp9Km+UZO8E+sDy/nw6lx7qK8kr
jTN0QRoDyJWjbc6B8hOgScZO5hFRohW1wIfsxuJZbx3CmYLEYYCIjTjj9VqfodwZNsmM838LG82X
OBBpbRN+f4gfgVWokg19IBie6mObTHjuSeQ3iETvizcOn5Im7mIU2sbh9BldYIvgVgYhR6i3GmCX
Fs1xjPR6TSI3s8VonBWRsOuDCZ2MSFWH4GdBHZa9d6xRxTq0u22nczsHyfTpEs8bxXnV72MBPLOH
fRF7RxKO3LZK+eym0wDfQ7JUNwLVY78b/l6G2XYIgx3Uiosy6weriDR8Q1EqDHiyTLenakf1Resj
PE7AvkKvr40M7oMzANTZS9IiWljPeCWSO1N4/FjjgzZdwfQ/ngIEborq3LaviGrMRONfXqROZ0Fe
fz8EnTZcBK3Ca4Stw3qgerl7TbbqnBsIn9932d5bm7+XLSZ1iYLByvXTt7p8tnyXi+pXhxrsUPAr
Ssz/RThFpWXQU2d3eZl+At9yc4uTwBDVE8nWGSuIqwBSw53PTFTb/Qc+MOXUC7lEBhpUmPZRXPPN
m7ZVEFH++3beQUXOlNpHjFcVH76lvM5xZkFRU1aHXxgtV/vDc+I0jNUhv1sxzo+79gyUSs2jJ6eE
TNnbBupUx8CVyz4k2+xxepIOLTqXlSDXd7mTeivB2rytEoUcgjuTCee1Y2G1bfDZBM9jpg9OYXHX
nXTMREAeyCF6RvtZWsA/Lqr/eJLSNLKIE5vdDE+Fxt0Y9HNbRM5nQme4xxd+QtLDPrh8ThUcj6Gv
LfhbJxpsfZgoMc6s/7DDA+O5K6tf3Logo3rHcsMMGXOrvuVoCFPFlUDQXvQTuH5xRuJyOQvTNAtN
Ui7zm7goLKnK3Cw9UbnEmxBJIL3Osmw9QohxOoPxZRh/2HYLU4OSPYzk+FwbL72JMnMFN/nZPd6I
XAj28afpVrK6CB2DVYMUn1/6Gk1P36szEXY+SQIGShm/PStmk9cR4eRTcBsRq/a/t1KyhQa2n10p
djVgIM/D1vo7dAts34TzsvRvliLa0hMTk9qIHSw1l4t39wrW9bdwMXpiWV4aXvnr4ARjHqh+ymjY
iseg5mo2yvOo21qDQEDO10rT7YTwXA/ls0iZWfK0U7TUZYAsdt25YqIyvDuVLCddJwE29zdbf3QJ
OH0wVNAIeqdJaIAGz9iBo2JOqDNmbvs/Yuytgnm0R+2WxyMfE77zlAHtTGmR9cwciSBneQMTjlWZ
FJdnFz5h3fPedDhrrsZA5oQGj8saPHzPp6LTXc/F4FzbKd3Ie+kd0zD4wAqDC4a/GuEJE4q4syXi
D2rqJHWgZ9DE3CkyuniVcHpqtflt/NmiXzWvGvbWpE6hqt3JQNOZJwBgWOOuJMaCmU2sajjCi3k7
yOXIf5f5YGedRgBrUeaYpVR/BLr35OaFwZgNgnGu4G2ijokCU5xfHLojKpPXCF/kljDvPkFNYCkM
Cm4eLd5T3NC0cMOL01doYcqcIVDqG+RjEG0zHyJFuv7midMIKQOz6j3Ytv4AkypMPodgpX1Y1wvv
BPGO7hS6voI67EZUPi5F/tanVIhZ9LN0mvNXtgyhaAym+faXRkYxry9KNxH4RRMwSf7tB8aw8dC+
ok9EBTy0OMq75zXSHayANDbd3CeuAqZPDdxM3PmwA7vtlFlEw3pfXMKKJIfgIi2/Lfgm8mhmo8Fh
avhAXp3LPFIW/SUa4Sl/ZLxnUD0/BaZR3GbcCmZ9vh2ELkeovb5xxHw5kGotyp/CTa0NukJMifmR
KpibsiafjzIDJ6VnybCnh4TMP37kktlLkD8kY9Sb2xIjUPJJHnMr0dkfGcmcoqN2uJ2+ICWYj3Je
yIGnP8s9DMxWhyusHxEayusxuf12Egu6i1lJs7ruVD7d/QVzXQJMt85Y0lTTxFXpa7g4ZctFojPG
TtqSvJz+Zw/ye52SyLWslZgJ4dSHuGq4Xl89F+LEghK5lHU2O7GfVLJ4rRtVcBHqNKKKMdl0m2Pn
ao0fWSFJSOa30bfl1PiyhQ6CmIlP2jHAKuniSZqSOiLw4rvLfhBFnyV6Fdgf7uG+wXhnWNgZ/mS0
uOL4+7bJWQ1EsmGGnV9TwltatuDb4IlQBzm29HrJ9Ge0PSW/WmiTWELk0QxGhSg9ukTHLt4ALK5b
glgwZ392FKX9FV4iijRX4UZ6en8Eu+B1XZTNeyyGQvq67tzwulkZdBGkzSf8CXIt+AfINjPgh8zD
LZuynM1ZSiHC3TOVbGbYLU5EDe4Wiy/PNU9aleGEVYr3X1ahjbHWqDNrd/0qY8xyMmPvMa2JTs1N
hF0Gq8SgPiNx72c6Mj4cD+1Ccg+3JYr2BTmJZvcX8WTvoXT/XsxNEshV8nDiQ/GpaRqR3ZhOsSL/
4EzPwzWi9kGPnj7Ji6/MqKejhM4WAzMiL4FqvvqZPfFKqPvTA9MOi4s1g5G6CxuIRzTjfVV0KWDK
hcQJtRI4TI2MaEATJ38kVyjnfexd50cR+qPGVs/D/EO/dc9mDf3GE1fp5jkd4HPj1DoTlWT4kR58
khP/fcwLcJquNAea0iiSmkFpkIdw/OyXdDjDRrFxziLeGELijQFnoONwivBOMc0tCSHEEDYJA4kq
Vi5d4xDnW0F8g/7/W3mwSFAZvoAgvZ3h87Cai1QUEOakPV8jhMbhFbkIQRq6ZBNNYUg9b3yV8j8o
93+g1JWSmnggvovXKaid/1+XDb43PEJK8VGtcugJHnDqqsFLNMpQKBG2rqOpY+xHssCSHW+IIAG1
/SYTohxiGbITm9Wke+SuWSNW3vD5MvY39OOTKKYSV+hjgR/XijnwEG2wQsBS2SDX4tj+ibiCBGQ+
WKvtayWN+of3eFlC6Gu7CZxYMcj3mI/xOREjdsNj0CjOkO63LnwkUkawvz/c3/dYp76qkPehUAlx
Ky5CJ54NYZjzd3ZUaDL4w2bWrLFo86z76SmGbcAkinoWebrxVt2u7B2TYc9vZSSTTI7dW0tyUiMo
/Jia0tPhu1GzNHYhEppSx1D8yP5iCATwf4xBiMPtOrmYyWVbORkbDSE4hR7wrQaKkn4yZ/wnEuah
RaT/OUJvb3jdGDNqCSYfxIRDykcMyUO4/t35PFA880+S61vJQ+/v+cfCbVpJ2o4De4lZgs8qo7vz
4s0NiPeb/f2ASOIPj1e868xTRLhVPQNW2heGPs1I87dTYw2kChmC8g1STSdS2r0j8eTo1u/PGXov
cAnEP5qokh7/DmTued00VDTwBPTa8rxacRPEyaMjTtxuBTv1XRgpTm60lQH4LZjvepq4L0FoFRl/
XLfKpZB40pmQ+ZGksccNq1JjzYr9Sze8rNVi7/0bxM2+O4RH/uwQyyVlPyqxpymRwDo4XOKzlFvP
fqYzt1HxDWh3NXbLjRSs+i+IYARHyBdfcoLfckNEXPUd7c7IpfRslXAMiG8iF0N+CK0iA0fz9pA7
jLddMBlZxtYDr76/YvrExCBBD1rudgGSYZDMkYpL7Gtac1xPrheNNept5un9USMmne0CqskbRynU
tZIlC39JI2AkDfBCd/7AExiyEMkepBT/BC+2Z4GafQWMgOdqxPvS6vYo3+re7FOHBkJM5mzHukYW
/UnUaEg9TUa+rkLCDCTWa/1qEgAdLzUuQxEKvqvOrEYopDysZ3k0mm7mJICX/qFbQ8sdmzkxCxFw
BUGxAid2jRJbb99DWvOXtEhY8UJd8nAK2iKowkd+AoXCRxnhr8pkd2saS1kURJg/z/TxdXHGVvL/
0Jdtm05JbC+ge3BHD0oyOfonb6kzOhXOwwLpSS8GTOKvp52vAXOcy7CUItbv8ERjj3fkpVuzZSOn
tckxF8PrYERT1xZlSS/5b708bIgRlNdqmO8/VTG8bEUHITIg7ICMaChbvRdD89cWbcwnTBD6zSgR
2oyEmDkovLBTnvQO41XC69UVLg5Qe+rMw0yK02YrFMHyiNURlcuZ9M1daMunWZif70oAAJAQ6vNU
dSQIocJZ0x1EpigKP2zeyvM0YNdWrdVtzb8OgcH9vAiwnSO/sNURPMYmTIlO2eFwd3+B1am3tfAT
fFMSbjDgn/nCT923mjxXH1Kzd7GWXsxRRB4T2XI21SmCAOpJuBBpLbRcC/nx9f/XzpximeUZRu+N
Xk3TIaHa3c+Bp45uLMkM02U/Xm8Az9rUCoQutiAkkUlxJXFY24ZtdQVSIha2lF46YWKBxUfIn+y4
1pVpc4gEmBMIP13uCnL+LSvdXccyC2VXM8rY1GoKnHZ+8EUxu6Q49NY0Q5dGkfyxgVm8WRfny+sp
mtkWPXGA4NhaBV2A+bFoVqlWFd6e0MB/nMjFVTE95gpjy0avsevCgxnO+en/CmbxeJvDErnzm7Eq
J5wvzdzfrZUT8o4KvPxEa0Ad0IRn8KuKh6jcPEZE8v2XNIolysMO6EewnPv5FVa8Pu9dutZJi8N3
+TY81Wopy6t22rXZ8a0gWImiF/HLWcsqRCSUMVsMwd24s4VhSDscOIDqvkV1st30fnECyn3MYll9
RABBfNEIpc2Oka5FvBcexafznbOFo+eCR6e5sntHEQRcdv9BDZijZutLVdX1idnbKXYTtuk6B6kp
D7teRealxnc7QEw7ggRzFlK6bTmZkFTuh5SImy2O+yChP8mgsDcsLSTLJcJg79Pz8oeG74+d271l
DgnCBH3jw5RdKDIusod8Z9dXOX4YyahJRsFEJ6/RRvtv83lG201UVoMhKNxYIiFsZeSYI2NZt3jx
4HZMc9zdpiLG6Ld5WanWGOReRQDVb+oHmWpGd7TyhdoiCLXJZ0caIQN42PLxCtulPgGu/TbHVmfs
6MpF3VtHLRdjB5sR9CziDh5wiElcb1UlDxi8bIJGT8Trp68srU3SeLUkaoXangAGOiflOki1OTni
pU00+jDwxdWvquziiVOSusji0WxQSi8n4Dwr42p9SgsAUdOE1syNPbYQEAn3MdJX8w2lYM4i7kIB
LhOzZwe7ibzM/QYl3vnppNQAg7vZX/FinpFyAEoS7kVRXoKtWyTqbqJa3i8UJhwq5biXloGeq49K
nn9Il/q/pLwVoshEw2y2Qrd2LsrBziUbUfFnKNmHTjTNJ78ue1KGrKvQqsmsJHr6xwhnCm+hr+MV
NOvo8xH6f6RbOKshq4UclAkla+HQo8Wvh15WraP92o0k7vEuM/XjcLrCJrU6jWIKnuuNTKbwruyC
+nSOkpF30UnT4vI1dp8Cbxp4FX9gNYSA3Bp/fPA5WPMkHzMtfERrqOz3Q1f/sI9Z5LEO+5XV5+xD
bwDmeFg33CJDwTN1WKph5lOfViaBR/Kz2EPd6cqME1c/0tFRHSp+CR0JnX1yBcHVwK3HNwYWhiWl
U+60A/Q29Ps/1ybTZhr/v8Eu/2vqHs0YYdpI0LygI4L4SueQzyNAju33SAumYQYR6YqDnbOx8kZF
UOASQUFYKhTqevmQj7klDtolnGHvlUi6A/JAmtFZ5ipRgb88wgqfQYa/yBC9dJxevqM/K/XIKU8U
Q+ovPTZnMx7mtX26mL25HD0IIBJT/uEGvHepnz67lmv7ZTNKD4DbREG6TvLPEi0yiLDo8xki62zZ
H1JI5Hi5Iz3ThHdOyN/uxg2sVzJrit+wQm1Q7i5O/Zoj8y9i9WC5NDNdjDh1kY9dkVghuYyOwgTi
4yKDa8JqS4F4Lq4oNR5aj74P2YGGXMnN6rBs/Dlp7VSlI0wBccXJKuJRUudRIoa5EHX6h67CTCUe
2AxY8PigZxnuumO5d8a1UPLJMGZ+xVmD8pY01mUc2ypE0tdFEabH7Nl0HO8xzuDkJFr+VlETipcv
w8jW5Ys1EtpcfDjU9nArbCU/hHd4hh+CBX1BZDGoarK3wDxZeh0nfsep8dgyXJKyFlsHVAvcFXgp
kjV9jNnGfHO39N52606AOY2aJS+Uj15rZF+14s4O0ii1bhMxzP7QwdfEq0g8twiv9upj6SS8taWx
k2tRdnoFAj6MqD+xyVR0SyJUmWBPcE7Fm4INThzEqW8xjBNfm7GO7b4qRCJ/UJiqmRXQcA/Mzwak
PaYrnVIiVu0AQyyO1amgKy5qRVl1fKnsAZqS30Bbqbq6odTkueSFryebHdq1jNFSBgY1wDGI7Fy6
jODE6Rtxnesg/27UkYtIX+2ofqT4KrS7t66tivWeYTX14f/iofVu5EuxVp/J2VYZXLzsDJCtm/fr
sY5FreTL4zid1bZbHq2+1rzJGXHNbQPabowic7m9/3cUerelxHcIp0nGYFndHaMqGWnsnDIFvBXe
/s0jEccKSirZKrNIQt9LdIFBKueyKZGWGYOaIRFqmCuI626ut4ceS+5z6T5Zw4OBTotXWw9i1+HG
FhqFASPQk0blXMiqvNj05j3cfI+rZS9XAlmLSDpDLENJ+/4CKzp6ve+wf/E/ADSwA9478HU4x68s
w7izYOt/X+9fQW/+t2vXRWHg/Keq0IaLjJHQXpGwec0R1UhgrMA7gxTETL+mg0epgillRGdyU3cn
pnethAHlMwfqc1PVmlECcFFE8YDAl35j+x7mPynRo8VhnXTuBH+KtAjFuJ73qmMEjtkRGgLQgO8z
KZdGfLmrTPmfyMB65t4hUQwOQbRDwfc+fkJKfmbvHq33hvrNTpxnLTX1meXsOgSPv5ApeCQYLcpe
9bfi4gpR+x0xCR3zh7IEq5PBGTgjpLBjp/miNOAZPHiFWQcfB+bjvI1uSy7aoWMwhd7Do4g4n2Sh
/kpiv+DvxQui0buuqV9cMnhXOPCzqPV65zqwtX3EYYI8sCSx74xK3T0bs7y7rJ0MlOZtRL3OLlH8
z+RZSW8Oy+0JdXClHGlJq/BbM1pFJT8IvuuYjozMz2ZeC1hFEiRICwBha6NbQCDTYcdalkYsLb9g
aiKpoZ8cjTz14wn9yKALvvOHJDvE5D8fNsdqc1Vp2hr3BMqhODrsqmPY2xVXt8EBq6posJz53Zsu
Gp1gG0XUIk3s31AxplMn+2gdgqp1M+0Q19uoks1vTbSrCaJN5Wne1R0VdBjiKzEnj5psODA7W0ju
W4aw63dzLVPKeeIZfn2rYSuMNudZ14sAoY7lILrOrf4at7uxoUOx79gGFyrL52fu3mNAYvybe85h
SkIH2Pp16cjlXsnSuUaL1G514jtRj71ZYaH/acynale1L/RHZWs84NOhFEfcAJ+7vLX48dHXl4d/
ra2uvImMtHdZ5zFR7OIoLyNCxGCgYbzoYFpvknHaLfATmbUz6CZlJFto815y2eJiDdUz30qJ29rs
uDJ+ywfhzpIeE0vC6zUvt3OPDcYerAydFHc4FR64I4My2BASV7NzUoKaGJGKfM7724qGACRxVLK+
Iqhe6GjFwo0acxAo4N2tXqO9ZT8qM0kLFbvh9sG5mJgGJXzpkoVc2+vUldDVj4kI/BZ0pltr9KnW
vFejmmD1RN8XVQwfiu7FUpfR0VJqoxZiUbgLSJLkXzw9qE20DW7aZOsGbQB8aKD64AgMobbRNSfx
I2Gy51Km0vPHvPv11VxybJ9HVyJxQ1yZHLnn2k7jSWP1nA10pGE1LMACj85xSAasEpSZ3U74F1kv
4ArR/lXjEwf17NESIfk407Tx+9Zb4CA2EufObqzrXINIgGqiwdakG780tw1GwlUcrJCCuiKKLehY
ohhQOrwir/bYObyBcQxGfPzdQYau3mH8CKiRVWJJzQ5BLF9kar8+UondHmjXRpH9c6c4dpnUON7H
9sw/YcSUBWB5dCeTO3/5nnkWrehyGEG+LockItFRaw9lHsb6xfGt5TB3YoRzbKXUs+YMlmdaFBm7
VBekBb2rEA3ebPUFuenuwwHZBbIfElbij5wM2UBi0S+EIrg3UmMo/VQT+NVxTyE0SHrJDTXwoCCA
mPpydPxtjoOeki1N3/8e67PvDt8LNJrObNconQWwMHRKdmJ5p8Am268wO0CJMHPUixpnbhesHFxk
Y2AT2S4pD5keLb9BSui7Z9UvyNC4T+Us2TX8pBiO0pf9qXleF+Wx5wPWLNwtkc7GHYi/hjA9xDJj
tZBVCBkB8RB7nadjbx+BohYGxTUT/HVniUKNjSo9EJ+lL6WY0igYamCeuCEufbCyv0ZU+OAAbA7B
EyL1+/bmlYLwqcj9GOfFDeyxwTtCm9ie4uEM4nrXxPMj2B/iJgIpuA5Gp/D7D4iPcOHpIcztwcsS
CDjNh6ZcLbbHKsoJtVSgQqSPlouYs5H5rNKiDXQ9wVxHklvr1d7/heY9hDfYodWpl55wRrm0E3ib
3of6eiQoFTV6rvy2IVEls1RFW8V6HKLtdztEWF5XZbTxEHG86307sOdT1IU+fZ5bjmqV2DfSPAqT
kswyjoURNdrJogL/mPLaBnik8os29agCR5TvpeId+J+xeLMMjTFQNtGxpYRJH3UzeKPJmhOsDnU1
nCbfkAF5ObQR66jDSG/gzQb/3XW8cd5aW/Wh9pd1ZxSxLRdiS0JDggiVjKYEc67ALueuqn0UGOFU
sQG69eA/dCn9QrBZrSGtkFQ/ow/O/7PSWe0bA5txtqaB2KQbqjQN2w4FWApjKXplLX6vx9QNbxwo
s1LulPGhIXh95av7QoOojpjsjRR1E9Hnxbryho/M080tS7IwV2bI9LO2uqVOhTscg+P4R5+nOC6n
FYELI6LV+76pOGGH08QRQcfUz7zFg1FcYKQOuDLe1x7dpJaA/+fGBz6zhKuaz9M0uvcxBc2TgKFo
7gRtEJ4qAMn9yoZhG/NZ43ZR8QMCoVGlHKs8q9c7c+EOMxEUS7CGdqja+qniPV6RlOSB3R/dqpoi
dTpgFcTbJkBCRORkE1YAZ2kDDwvF7S0fiAxT8Q0ZYuplKepXvVSUagebVvYGeIpSHrfz7WqD6i2b
g9X1CTUnKlL4b5oVxQ+pK2NUsD8AiQTYrt6wWca6C/peG4Nd8jEWltrEtKdSvFzH1D+VKi1we8mf
hIQLPPKErxaRnsj7dtubFFiLc98ypQWolPkqAA9aslXu6yVT+D+HR7AfKG/FbZMzxKAbI4mufZAT
8TeyigCWYv/cjlpU2VtW+gczAeUQiUKv5ZEQ+0VLidZWqvfBsCXoQmYNbuGIkx8nF6/QHtZ7e4Ie
6kT10UclfsuEnwE0WwGiLbOx+9Gh2icazZRpsQMAnJUb+qx/Uosmc/j8/Lfkgtxt3Aern6g63OxE
Zo6aQQOdGJyT2thwtxIfVEHp+z8qDEY3XVfX24gVqSnCSh+V3VW21+WTV5D4x7oC+gwEdADGFmP0
2Urq3WEuyPaA5UzuDLsrGyDrdYVYFUikL4Oa1HkSH6Ikb9OuXtzbj6c1x6k8OpehyHL8G98bkO4N
7VxfjyxZYVLXohcflUN09GzQEErKs4EPKUYUdCZrTHvNO9FJqfdckiPQYkq5MrgDtOrnhIAWnCHe
765ib/76UrAMqaAwmkTHi26y76gjvg7FNnMrmKEGMroe1Zs/NqZJzBOUYw05kGqK4qz+ZW7FzdTu
lMavCZh8lrkb4r1lqiwe3o/c/u3Kx+Pc7NenhalPEuSmGfbleaJGvkC/p6NiQiXtamiLKAVJL4tf
CPD/xF+uT/+/XAQsaFxwA9bbqyOHgLjSaQXRzPO5z1lj6dj/nxZvcgPcOvErft9OcEc3vD3VsRVv
galz6XYq4/qL8j1OJXN53pCtyOAx3dY0f+6ceBD66zJGHHZ5IaGi1WmT6drQ7nYdREg4BYqMc/5s
6WFpTeHkuWAxVMV+L6ghjoZp8N4Z3IL28neHT5EiNJ/AaKOq6OY287aSualPNQow0nhlVeqHivJ/
mwaYw9B3ZKNWxpvxWfBZUp/waZoofZfXjONaMSZh11yqgDRJ3wIXhm0NTuOrTh73ttAkwAh0T/SM
3+7esR0jD2p6c10rUGvKiTyf6YkWb5EJUyg4vRex9jHc65tNUBJWtMebkeQNFqLgUHTzq9NAVFlS
Rip3Uacyz4W3+NiyqBJjXUQdefB7SHKCeCZULQpzLmw3qtJRGognI5hPDKVRmByhTuD0aA6tP9Y+
rLNmpuEQH/QhhXnOFhKCXlGMZmNx+hz0JiQ0CvVBL+5Ek8tiAdfN2XSOcyhI2VS+Ftwj3wHbDPjd
xbjyuZqd0fAY+WALe/r1O9LXTtIs/07iNd6vmrM3BunDdner0pIQp1mYmDQnbWLHjGIt79HGAsyr
6W5I2020E4j+B5VS+cW/pH8nDRSolGMsRMPC0nC45aeKZvoOC+ltzD7yv7lNOkcGHvQ2I7oSNKfq
BMAJ89TiE+pgaD/+Kplck02qH0ZTpemv5hmkQbLs64AreyEby3ISvcD4HvzR7/9Y14QsgBG7tDD9
jIPNhVkHAhOLGyJ5DJ0MY2k7Vxdq36GST7TJncDJxo57Avuz2ErOl70sTjnQ8d2Ca/42/mtr6jX/
OEHfiWKvHsoBT8II31xKEUQQTmI5ojQvZeyctsubzGs0j3z//XzvDTSoOIgqV991waC8//VjVmK0
OxzQUGe22YaHVs+TFGh19CusMNfIivmICqRQpRDmM0+hJaeUCk4RVVc/fhlL62G2M4hNvznfNyn7
05dNXvY+d+D2s+MgaJ90IpmyeGrsvwiOYMa8H4T2Y55QRScpHGbu93WeElFsFDiy7MwFQa8l4+BC
3QyyVK7YqJlAElSg1zs6BL6/sWsnR4PKS1cXZtAu5g3OSi2M7TQ9gq53+1NiOUJ+TXuW1fA0zMfI
b54eXZ7ahPxEwQ+Br/7/cYR7ObXIThKFYrND8CTH2gR6if4AgQzsW1TbF11LHYPvHI3wePd4byCz
Yc3ynVoF6+4RmIQZKhmSw/4xNXJbd8LLMXD38i1n6fQTpUy0dxR8j56bk5AxM6lp9FXlIHtqeInt
1xIdgwX4gOZlggeWXSmKCCjfIfNqoeZUeDuven9MKM3xXrlUtoyVajoYlp7KU/LmdSLZq5lYMSGV
WR74Y7fiP6CtZz6ON4ZtFxazAegOV3t5QMw9paVMcdAvIbtbiP/wx3JOS78BRI7AbNlS9/WQkLKv
U3WUWLMsoAKBT206gQ+zACpBszLTiQeJMKNlUvnglqePbSCR9fX8M7Gum7sNzGni+XUV0Ir5/eBk
Sh8rBv9tHGtqbquN4HE8xEqcSD1TL3+2zPVf3rChvCzo3k7mRCedriBtQBIM34KLKppfb5wQ+kqu
KLAaaSwE7QzfxFVu9xQPpRsIhyRUAlk8IpfLqyKfZP23NhbEquVN2fONxM/++UjKOqC1hCm/wTop
odjvgBCp1RVmxx549aI1S01VMZr9XcZVx0wCRbfZVP+ndA3sloMW0alQJnOBhYuC1LRXlTGVrOc5
S/71qSsukWeE4riRfXbjZegkshQ2cZgqLYxqSV4gf9yPlciPc+zXfSZ34YXnXmyL3VTpS9aRcdiD
a1A4F+NEkfMPA8aIDXf+XwvqMhtEVBabXciRmja7S4gaBc1FrF9CF7cqAxUpKXChyVqNDXu5ZbJe
GdEGsTQHMJyRYKmSxToNl0pEbp0swcjRdChqaxnPccuNDcl0nh5Y4/Sx8f7FythuPr1XjJ+3UDy2
jXa3yM7XebmPgBdEY3ikv85QS9aJDHhpmdpPsOY/PfQgfrpBatFgUeDZduD2bTzfcnGsTarclwXE
qxQTVi2xKjfc5bv3RkAWLp2s7JdrPI/TLKXf2HefF/tuCftENTLohzQ543uqDPN3hEAhog9loRq3
NfsK3JH74v2L2K9g+wlkSAMb8WAh1su/IalOhY0DPKu13pDwR2YDsvMzOBKJd/M3CfPcph297RWH
bNEa66NGpy8RXe8jerCBF/Hu8neaBx4yiaLnG/nxG/vueploW2/tyTemb4v1WZUPlUF1HrQjrIFa
T2H9Ue4LtHWqWZ4k3ZcaZlYD3mSBr3pAVfTH5O0EBRWZePiuuYTjm/+x3PxvT8AfBL1ntfaFdC/8
EVyFLJSy+hqvToEW3ntCqNI3MYmXAf/dlng5G7SY4eTXIS2GecCQ6jsiyBbOU5nvF4jw83ddrffP
vzFpVN4g789p+3aAChEtF5NSRnjWgMZgRTEcurpeIA+hPI+lGi+5BzYx/FQYIoh2RKaL58iahUL9
caAzOvGMrdDXD5zqofDxWlus0E+X61jzcvR2GX+sSRs7LFTiL0m12pzQn0+kicXC04uqP7dUR74i
zHgsjF/MYNf0htDzeZOqYYkyxSJkVKJwyOCBZMbDnfSsHt5ka44JTmdO1sjuTCvaGiTwAWNbA1+h
nVsr4nxL26udwNFEbI7qUfVKwbNz00NDnfbLnZtQSLEn6uVt/qF97A5ycji724rpoPmthaxdWoyy
rK4W/bJglIvK0G9tuylgjU6h2JQ0iNpLxyLJimkZu788nn+uXlUiKUatjVzC1PFZWvsc3O4Xv3zu
D4ywKt9yElZOTF2sZ7ImqpDLXIk+/Djj00OJ4YaTD716EG7R9xLIUP9UYEHayu5KfoYXXEineEXU
au1Fri8lf1svt2ByoTKjspA0D/nVbHXBLiezW/oBwyUiA5RHPJp00nQ16mgnj7sbDy0c45x2ae2R
FZInt7bSuuIS2Y80lk1ZcRZp+iQ+KJamRZC0ZxgN47Qg5nwk6ZFXFxCvt/dxGAIgqab3mEzv1aQh
3ZX7Wp81fXJW4oACV41Z9nqkUtr9GckbuzRCo+v1VI2DUZmyzulYsrosllgzsNELxd/8JoiCkQK5
XoRk6HDQzUeiA6M2cDeWIMJcQN09rSOJNf0eJ7LYctIrABLOYbm/eutWfvxmA/TVFn2oJQS5r1ZH
7I9tdRoGgwlNfN0NdoL+ANeOK5N7KggL0fpUl8EzRhcAJOC+Iin8tdksp6oT0XZSu/LQrlh9iac1
kbFjNqvDuTKAX1b+jpkOqZ1+08VmprBo+fnrrc0mcv9GvUI+bfvVAInxc7kxddnkeokmMuL5ugpD
8LIgeS5RzGLkvri284rfKyuIH+Yibc1dja1F79nrrrXgYl2IxZXXZLbwUuN8Z4gt4PlUapcFVmcI
s+dssFzHFNczQM7KweLltr7P35Vt0GxU0KDnM6uNv6i5E/FRsOuYKxxtlwn4vfZc1A3+LLOnLU8C
zfVFkzpKgl7dTCjo6czo7k2NOETyqmBGpFBiYeosWcm4pBYzZQOQc3aBYkjm1+rKungeF+EX6GF0
bEfw0JdqtHGTKkyany4+I28eho5MtlVehdjrMA6/zOSRthOjkNlayKywHilfPaU5VXJYaKVLnyI4
tPaDtofHGM7FdmCUgTCtocFI9oEPqHENuvNbxif/cEru2bVVOERdnXrxbRXIW7AqFQWRBRzGuHyW
ZXDCI8Hhpl9/9i4wB9zlQ2IhOHpxUfASrKgqu+0yXyNSdW4NpVip0KeXytB4Cq7a4uHIUURBSG4H
NAR901SZX9fXsusEDELldZeUNQMBRGPFWm/VA+zRrk1scmzB3q8G4UpFFKomrUR2xeThYmbQ44Ek
YvVfOFrYbctwoOizYMobFXfsgegwPh3s2EhIb7n/EslWPqnWVXT5Cw7aZUBCE9iBT4gMD0eJj8c3
CpytBTBP8IvhCBw6l/0eOFBUDBjyPSoAKFMMPd4wdRe7ygXOT4cAMPi9m4P+qW+dtZZQ6zL4F+pB
ilBfzeXfOSOIV/6dSwsMGjUuitxRqUifmlcSOJAZK2/aAn+vXwCW3ps9/0gkURJ7Sz71mDFLG2rD
YZ9DW2w9x5MP/EDT3RX0CpbCR74lVVbuFCV+pvLl6/KUWarfIlsPdQWK7meRnjUclUJ4+m8Ww4ke
sh54S/U7y0pv34CCtlivgKpC3WSjSpKTlUWVmiQfubrA969pBNSfknxwHEwCjkMrXoe9GwJ0qVFn
nhDOhHwdOE2G17sz2XG7kbwNIJxuNbHi1Yq63nVqJCVA/SyW4syADyTLipBI+mAceArpxPTrLQAL
UG+u2yS8CTNAd68GO/GPexYK+wyyY1mo/UQqp8586DrBs3i3P2Mbo4UGskKBQJ6kmAiUcnOjIpSB
AxLLMzSxS55G4yjPnAc5Z8b3K2RDY6mdUFneQJa/6NpplRLNRWSvoAPhczs7BJNegHF8o6BBBPSF
PeL3b7NPj98weMl000CrN+dJB//MRpdtUfYjQ0YdLLgnS3yAzudrBZBM4hkKT56JeXfar7eXpx4v
4kqTSdZFt0ns7X/fDMHRU0bXWSLdSwd+heaXpNGvnjXCbdYAZm9UXhBiHZmu3Vj9wEhNZqumUvdQ
nOzS6cq22YOlteH8rSIzeLuzYdCcqwknWEE+NyKxrS6eah6Er+3ZWbaKh1T1kay2yRD5n/g6PD+/
kzdxa2upRbi0jRYxGZV2y7adY9xrgT2qLzhBPyzaBdgl1rLf8ycpi6SR7as7gy5BahtiCumJaOJg
g7Xg+W9kdwDGBHBWWxGBNvRjFrxOVVDd/8CtUU3eXVn6ySTrys6zvdBuXopHcuVk24YBzJHA+QKq
gkmACtYrpwVBwOfBFTvwGOpUp6eZz+75YMm7d84CoYLkf+e09ay6yU6VgsIVm/s0BOpfVOdhOg3f
q3Sl4tIKi2rOWsBj/a+xaVNMU/eDVzf59I2kqGsiaKl1nBH0ImLjAJZlUEBCoQgC+NSQ5nr4FNHF
2bV9EZJdVVYSBlmIH0VL0uRPKLVSAALOm2mQ1Hte9TX7Qpwk4DZyiwlYNTx1f02p8rpakdACC8EF
dOJjW2eyuQsi/J0SMEcjTFXUzp6GT0DRhlfQxjQX/fqQ0ZyFCq/yeepJsJybn6UBbbeusHYstw0X
Fskn/tfYaAyDtK06fJkYXslBYauleYJ9o6i+T2kBn81xhqZhIzrrnKPOoA0m5jQp7hUhsPmT+vTf
OXmUWMTF5Udq90wCqb9NNLT9iSzV+BYQZ1+4SWpG1Kplh26polbrQc6gWdklxmA4Hhmepd63/gU3
Trv0wGbKPtkL8noqMVaI2i4D7WK5/0SezkuQYf6nLEUoZp2srsWsUz8gcKZbX/GuYYdPlNEtPcTF
n2XQa/qoyu++xrO8J6S5ubEaydpOo8DYL2D9C8uhbTKvjikZwPiYCVM05gP9ICvFOwUeOOzZdqFp
hCmEEN80yBRKeKqdkr+LbjvvZiOwEmeLe81QkZMqSJJ1Z8+Wc7NB0EBFKMK5+y0SkCL0gwxCRAIk
BfWGBj3sR0Vo5ezbVcX2FLn4/Z61S272cjzhPqXdv6q4ohwr+jkQd2k4JbzTfGaiw49QrOQRcDM/
vMQnZeHGR4EstM7TA/pjS+6ln1c2fUFEjHibjGLNtecUX/u/xd1yCGHnW643rbiZ1US/5WYV28nT
mNNLsv56kuOnP1HdIXD9xWdIHYCGLlI5vZziaH+gQN8zkJI9arlmtWaWyna+RDvecDRyvT98fHMK
euQsN0O/a36TA7xiTDdnern1XAF9rtpoQEQe+cQBp/19PmLBILrcsRG27C90DrcpKWHh90Wmi4rA
mhmkr1B2QHqMhcP1MwnOKpuLtD8CrFsfC61PE7IF0tCiCnYgdFE4IY741hzZ1TNGqO+pZE8s1j0l
NDpbn1GvYcllwwPTS438PliXKns0r8HR0yfH6mE1e7YTjxFaatNXsqWrSAoRuJl7jjWWMBKS7aiw
O9M++gTiO9yXFK0vf1PAq4FTudxTi3c+9XvZ4ejv28rc9mwTpjR3d1Oc4Vjcydq/aREJFnYkW7qk
UyjEMAE9rGHmhF43nHp6iO73ixN6N+HtuRgqHek8x2AYzAiLMIq1r6IfuWATs7M28X6z+X/JlAG/
OuLr426bfxJOQ8FSks15zXeZzktnd2aZUEUQqv0e5V6cnwOkiGo5xvhGjWVp7XpZWVDI7Q2ETyPM
RCI8Tec/mUblV6J33LVL9d5HDwTcvZoZXJdO17Xp+qwsOKttxAKgEyOGJOnNtwxGkXfZ3Q0MxUZx
eFvuF8TgQ4sC/nU/3Uigy7cCMXmrTYHX2+a8Mp4Ro/SzjWDIOO9YUM3s6A1oo4qpCzXQ3XFS9Myu
OVF1HaGssatr1eejiMPsnfTIbHERMwQ7jhkiorfkeDGdrFgbnlf7az6sm/WTl36lp2qR4Z1XJ47j
jvAKexgW/o76WzrfiCas8Npn87uSAb4OClPNsMEi7luzisQ6rJY4bgqJ3xv+Ik1QEGZahr9pXd+S
GVLG7aF/wYDPwLTKQQ5ulD+0NhAJ86EJvQviB++8LfgjcwNuBb3Z4fmMBschFi8JCvBnNpFliRUK
N+wkd7Oievbfl8p2+ABd55HzrAb2utrflTTBs/+Ah14q8rfhaEY8gD3KZMUtBtRNwHkEoHmtpvAU
owv99MykY2SDV7meh27VLdbeWkLTYWT1zGPGSvlVfnzFH6YTHYaBCTglPyhLZ79wu/bBLthCxdTm
EHdJUI4gDwfJ+TUvA3igw652pAQdU+B67CAY6x6ShmVBatZ5tbPof5+wQSgcjxg6vQoioOCwtj+q
hFMzeg5oF1yRkkSB0ix59JE9YmRU3DADOXpuxOB0x9T4iiCo+bVik3x3B15eE2OjlRaQuJyX9HeD
lzLeuOwIOkD9QdjC1WdXGXXW147E+mowwc+JuRZsongb2bJfTXTw1qai45YPXxvdGDFeDC0/Az7Y
pe59xOxZ2HLIEf/BDLe9LwQVro2HN7cV+ZPrhv0OyhHDcbEXHOV7ODOnSNHg8bC67YC3q9Wt1ygB
ul5s49QKuNYCrW18+LzTXnlBvijV1KtXlFNl2ZXiz3cQwnjOnbl4KshM5JzmTjGlNrJePkpT5kWo
LT0qHYCgn8hS1T6ptC68o488hKHQgnPCc1qcGevHFUkeYz7ttiIMRUB6I0v63ZmV1vBj51ZCVQ5H
L18dNhOFfx8V97lkzBtUpJ3M/opLQ3Rg/lMayn+fktPOYLbjPjrKQz8I66yKC0vBVkCvWhvUsYJO
J4fNSRA0HquN8s8iY6ikRhE4hmz09jLIwYNgUl86n6QERE0IeuafPzcaQaNjbUhREYB6NYql8WFB
oZZMGa1pL/eE+RElinm80Nvfgfi1R1EPvADEdC2sBIEbMI2cruwys+fhpJHye7eJacRzQi8ODmbk
LPPtgY6ixYvAq1r8Lmk6uiXC6/N9vL5SvX+QSn75Untv0e0DF0t8B6AhjVyiO6Pm9J/U74xcKiYX
+fAW/XnA8UTyOCKqRRUtgOR5OpQOcWoMTUf3yH861l587ZD8fRy6TMuKmdP5aE20dd1XeWdJ3Ska
gcKyZZvSzz5lnDDrbo0GrLZ1kbicQyM9SVinTD3r2QNUVEmJ7gQsTJFJ7z46oZyvk/02tO9C7D9j
Oc/Zy01m8cHgrxyZNu/OOP7+FWzv0GC3tGB0nmzrlaFuwA9tCD8bs8pGhwnxjdCEn08Kb7TJVW53
z3Zyl90C4+TuHmXLSeZjRAsO/kN5cZbPL0MckV1lT9D1uABJ1x1/xPSxZ/2oYE+XrVQF48dRz6R6
9Juyh+a605FtmAh4SOGB8238K3kD4JUGzy1Zl5+4tHNEZmMNhIh2BDH3/GSkZzLueNOSQyV/yQSE
GkzQnHh9a8qxo/a4dg8k3QYkIKSVM9491KeP8QeCCTcNmZ/mhEixpVeMJsdxwzrKr4R2qFm3uw87
lSBRCD4vz4AHeIy5bTsTrXVl3uoyBqJ82DRFnMXwNqUWoXTHzjRhDjUSdctlipITORlxRQAOXvRR
ja97XoLH4u5FHFizC2RodHBEqczS2XmHj+tg4/l8dsBwiX9nLffEGiweV2LefXSUs5fEiPrr+oX9
cREHXUxB99d6rjwwm7Pu3/h7DNS0Q5+FCFPB0N8C/xDfjmZZUPd8JbO0+QzKKjn54U4sqkkgmdG4
rr8bFF4JV5bTrpcIQeWPy7gqykJfYs+g94K5Ag9XAAsdxnpjjhSiWWXv2Ihw+J26NS4FXVLnrXGQ
4xDZpP6s16nb8WqnCCKl0TOHv9NYooaMTQMWqtGcBY6LHatEfA+FC0LB6OoRUCjIueM15PdBc/jF
eQVU9rFxV1r8jZgnRdf0zu4IFd6HZ+NM8sWQLhO219XkduSZ/bJR5l0U4Jwq7UpY+26MFeDERLhH
S0eQWCsv7r+b9oQqKSxX818rmGROPyfXVrC3QvfL7l2MVN8OZtwnR1hFLKGeLMAJbCTuyelRyyat
iDvUtE+sxhTUOVO1F1K9EIkjkXgRRnVdP1+/7bIawbAtlLTJTsDwZJfJeC+McdsFaTmhW26Rtir8
GGec9Sx5Zug6x1jjTMdMYdK6jNBXeekqsoIFFdMB+YK6sdLlqI6RR7BTJBT5PjQjcBhhgb51VwBX
MQAp7cpJh4B0wiT50Sm/wJTjtlpW9ZXnV9l6U355lycr9mXuI32+x5/P+5ElwoZM63iZlPwQnO2j
SVEprOswBRkohYgoYPBB9uP3XbTUM4pg85v4sVRrSBVP8D1DwvW+U1YfKtXPeKlq2NCj/OWbvrKR
Es4z+BCc6iH2te5SAFTka82uHWTvRaidBgJ1Y1F0JR0VbV51VULs+b6T1EG9v27Mnw21vgmPW10q
MIN9FPiX578LIW0skFWfbCUOQKltWsmEOKF8zFXDeOgcCPUapTj3BMMbEtQZ0ftPQKm6uFjD7JTt
5dh7eruZCxULzf29Br8+HRbjNI5Z6t6HhHyJzaE3b8OHL+Ddz33+1F5QH0ai3JFQIdzBT89mYRc7
OHaBUbsvB3lJy8lVzXrZujLjfYxdeMOoNpOmx8PQ+jGcrAO3A0MPAuAtfiTdRCST05NDEcLgIFGU
rNv4YrnRH1+WtPHJFROLA1M/Pkr7j5j1ZUMFQt93pUvYSpNfRy82LUNWabpXmcFUq4FMcTAiEgmn
qL+rAyGa4ItFifvyJEFlzTXzYSItSApvDhxzdUlYppu9NwwA/bwxln1AEC06Dl+ac7FJU3qWh1yw
R+HSHAOEiaSmjB2tJ8SlhqqnHwVMBOuhqGSfiNwAwIDlC598mkW8AjwvuQfY9Dpb5jTwAY6/EwXj
kXqEzGBpyCFbM/WCyxWUHa+rkFDLlBG7Rev6H1g/9PUOCcpYU96UuizxdVIaCpSN6DRxm1xZVjNs
U76mxmHLS2wrgRal3yJVtIPyQMxfcAvOT7CWwlLkXA7lG4pTHBNH1uAjK4vYmf4aOA/fiOnkLnO5
Z51NlTIdYpJTklxUn+XgMcbZp5JpkDu9kfl1huiXRKOgY4HTMYv78y55e0+4xvSoBNwJugUJODXL
HN+b5BRTHFKJPdjyghUTUzsW3gBxbVo7xI3Sx0IurodOav9fMmQ382vS3wfL1jp17hp3LpdGt7Tz
iHAV6QWRxCn5FOSOd4FNVKwYRr+HlQK5HgrlalEhN/lEBnU4+7WHKlqoVxJwHti/2NHIwFU7Xlce
xpZ/Chm93bzCsKUM9AvIUFjPuMMCxuNkT8Yg++ZeWKN/T6LXsQVCn4k37BKa8PaKEAfcQLlPlq9W
UNm7sdXDUh+MNPYT8ZNCWgdH+ROF6NgrvGAtzu1+S6yhswccNTuF9Dd8uFMkpzXbANd4nqVjLBom
PsqXYf+AtfFPpDwQT1ipi4PoGb60mWrCpVGYUGxraTZZ9Vk1nYERciXwCSIOKqAkCIF3AXX5scRe
NGTL5UdFo3mvXivxLQNNQt2p4vvOge+9gUsvPRWY/3hBCsSD8eZoOxAAJk/L5Bp220RLT+Di+ew0
14jWsCK6zpP0wzKihj71WlVA5rvtaJJPH/3baHF80l15USgr5PzsDCAtbGuiwTShd8du7KRcYnoC
0OVF2p6JlU7CEqijefvXzPuJn7J8WAvLgDpCwmGFbuZlraURWUXKBCeXRQAjg3KnTA0hF9OcVgL6
FmYME9+rPWyHJiSoW44HjfTcRdL672DFEs9ZNAmOJb3zFqp7TcV9jKMi1tvl6+LDus4BkmaJGVjh
bOGHSoJQwm4o5h+sO/CZNTiI8qgNX0rI+heFN8oL2sD77LP+x5tGjEvL7aH2i7EI0JPLqESOIEQe
NUkwSXfeBpZsq/+GjzoCbK/czDAGpbQxF089GbK9JScmUNkwBcczd+PeGqAlvog9kHDYNW0aQYtF
gh0DBvI0TgHE2qTbPMoiYaGbsxH7EZ4FESlPTnHCfj+I3Uk76wtoKgROgfv7hQkJRtEuCsJpRUzi
xmF7ldbiSuMQ7oCSZqSMourYHHxuShQPBDWO0GP+aRg1bpCSwSSDEZbxDxElQKP35Ir1m5C7oFgq
9ZHrV65SUs8RnWrUwtYXOTo+OdzwtnIUcJwL7wJVIICfAkCStxHFYy8u2DhM+xODwRFWV+sBFOZI
vf7ZRI99yEfMYN2sb6wqlibgs7Pboku99lyWI4xUWhueHW8kc3jXe+4SQFTwkvKhaXIkKe/xZryw
lMhVxrx/reMWA2jaKuJAy8cZKgekgscgjxMTpzUhGbtiYVNSkLzIkRLbAKZJCv1/JyG665gc7rAX
Nfan81vo7lcfk4Hoj3vDpvjI6MGc4NsqWxqFJlrcanhuQuWqXcaSRn7RV3NlrVvDHlWhOroVTakq
QfAsCjreXbpe8xTZIzxvYMDXbN/xgpKhMs8t//Ez1D7jp5L/lDQgF5eJFryJtLQmJqL9OeOrsFLD
0jluEITp6aYJENAnlsK8gT44dPRpvTob9rzOFvQ5lzlxzosVqYsmKA7bpjm3oNPvAD8f4MZuklMk
/4BL01oR1y5Y55Ag1tufqvFmlX/wurSynmmNRPwNRR7cuVg8UyEf19VZ6E7cTLP0mZUjy+ppJFOR
eAWSAuYuHA3jt3657ZJ3WeoLqo5kykg5OlYp7IZ8ehORcTVtUx8CyEr9JHY/s7hNqi2HLFTOQ+oZ
vcxsTM3gm3JQ+HVYz07bQQjHsOuEQuU/+F0p3zf9NvM9RtV8QGat64h2gCrgbzobLucCYUZxfLkA
PDYFUT1OSYb321xRf7QWasxI8cuC1FXWc5JIaxT3KAffEiUm5CzWkM+YgcTKjIHib5C/bkRajjxM
TxSpd+21FxA91QAPZBFbw7nRjuFc+pbnj7mZVtf+oM0bzlpjVB8ZBRYQBeOGfwXQiUXuMvSrC+q6
FbWxSyGPhGdV3+8IdrexXG4q5hlIDOeoEMwNuL7c/83eopuUpZpBhx+/SuL5z2zmTyA/t9EKY3re
xlLc8nRKp8C7YvnZTbbngF3SaiWHdbNTUlQzgE8oHXikdr/ay0CqO9yV6T+O0aEPhQTzKjEVMQi2
fK7C8amhLmnG2sM8GK6wueJy+9tQqyhplvyZV8uPx5PDVqynKLkL2PXurnmge8d886fhhupGMX70
EJXhbVkjD11pscZMBXwFIpwxYFHNrgiXqoarnJATxGKd46T6vzswzkLSqzd7NfVDh301ODRYNd8/
EckgC6xxXy7O2AJKr6LSyaqQkysb2bdMGeNTwpvTnljyRkPiTHLtKrb7gQ/r3+J7gzP27LK2UarM
ol0VANrrBJKLBay6BSQIsACqbUAQdNMZ3dH4tf+tqNlASEMJsXT7nL5H9ySiUmfZuamyDCkRHCUj
0qtNhmc0xX7L5ODKF5RAIJeCZGe7i4QYCbkUW9AXaY+mOKq1J97tndlvfF5+/WXij4WGVoIU5fQ8
JPsXl3f7R15OnlOyqYRi6FjpyXxPyPu/fVAU5CoOs7tdxCglY/nGz1xwvd4cnradnF85vKN5/okI
qGHznFMSmeNkWyQqcrIu64VnG43QiazpX/2bhxQRdptM2MkfREpjoNivcXfq8WfdXtIpZzdWdohi
KVy0FnCZAlcHrli1Xa9wvaE+GbpLQIVNcSlmKch/ewvmpLw4xnpzbOOYY7+Hqo4wil/KN2TOqYTQ
618/UyuyFAM+9aCCxQ6kkHzHpo0zViTNZhQn/Ed1qaJzl3EWpwMeIrS9GGXohz7AFGOGjx6q0eQw
6KwCfKusyeTLOqpFDBKouTdUg2NqPIoGmJGmka6RPAH30jUnxQ9UL26cC+vmQNXBkj4S8oOMqxby
QDzKss42VAZTeXpZCkD/jR5LRWwDzQknW9cotB6WmvcAQI1pobHEOOqo2VEFuvqky3cfW7C1a5SO
+yemwl+tYFKPhxndhJ/Q2iB3LTCghK8+PjhZ0lIbiuTQGgaFKFOvVmKZ6id8D9ituRGdCz+Y3/Wg
TcjdrAPx79BP9FlecsWdZrDphikM10r1YIm42jXcpe1HWz7lqkXm8JpQaS09+2qlE/MHdh9PvbFx
KgtXkl9HTeJ1TgpY/ha1x2+ebfIFXhwG28i6xQkoXDUY5RDEp+QtWgprlozCQCPmOil/E4xjVVzb
OzMSjMOSXCt7JI1XAPJ/Mf9ZKklDMmgPB8WVCRRIfBfwtR8avbiROh/i3nz3MVFBhDCc7lbYEV4h
2KQqrTR9TVA4VUJLl8Z6wwEez6b1iJAFtTtmBhctt9YcFt2W1gRrystU3I7XOKkGrPT/Nm2sn6xT
k3R35OZIzrwqCDRCr42BS6ca356ebu5/Su33ZQyfuX6sPAkpFPpuATGngzdYDErQkYVM9eoTg8HF
6M01usIhuUMr94zlngBFLcx7hy6a0uMusTNuwlnxHPMKd0d8l0rpPA2hs+QDa2EJzI7NFgleOHMa
j5swHUAT6VSWb7S67HJ5mNhMGeWqWKgsKlNR3VgDNerVaqRB2Z+dTHzhoD4wM1za2eJ7w0bSa7Q3
pIb5aIqaRGEioRDqKqMbnd1VNZogSxzAhxc5SbOt3apEmnF54vjbKSMHwQNrGW9GgSDMNJ+gdYre
ORVVIB0/+WxPkvavrOMJN+yR+TjdM8QSL5bmsBN2QIQAeb7UwuBazw8PbyJtAKDDcNYIJyxtsAQc
3bsqlZBv2f/1MaQp625h7KrYDWA5sO8WNJfbxHjWchH1yECqSpdySBQTQtjFNHzPhxIUG4o2Ic5D
h5AhfhUl2oK7QHp4bkqvhQ0Cq9yb419PLGU7zza1pm+Yb+KUVR3r30u5kKyGzcWXW5Pg4Mqe+b1L
vbLQ2lFUnQ6nHRI4zjd1KDFfiw1VcCsmhcpfQAY/xNxtJlfoPuRx2OAbhPtJi06E3kaK8su1dpKn
LIRz/xrwzgj/9QhZgPQta2Y5d7xV0ETwN4qhJ//+vrwlv1telyEFW6jS2Ju/xKMJ8iFHOLQfLUX0
pCrOMZdQRznFgjVT5jgyVzP2vfY+GO7+uAEhzmmDQPC7er6VdVcTMjQfuoPI+4W2jcDZ1hOl/29h
8YI3r7AjO5n9mJrq63bgQqJ/n55wwfX5W5fimkONj43pv3r0EFb6iNkYSGejUKO6bOBhcBerLWRu
/RXorDsY4/4JtlJNJRaikucwkjk/0Lh12/mV+ZxyAqp4zrJ9HFkdwEROrQrFFjB3J1uGv/QfQxY6
bI1TMBrWsfGqlGNbBDfLTjlSUGey08uP7V3xCo+cjP6uzhKYvTSNZV/95Fan2MH3/SpXEHgAEcXc
xSw7i4rjURqujtxlvSK9mCjCuODRHBQUDVV38rirPNEwAQx3crLFc1CXN7LK1CL6BdZL4gDjC0IS
aNzwTb7ujPPSVMBPVJn32z9NtKA9BfXOTKtBgdRoQ5yHk3dpQI81G72T/noo215y0ESlEptWitb5
NfMEi/3NIF49aGdGwSJ4PSP4ECPID25kx4NmzTCvOVXryJUYSa8NIboRBZInlXbq5Rh8xQYDuSQg
UHLde8YRQOLPNHUnIYSo1quMWJ93O47tP0BqvYOcx+2e6nHXxppKNZoKwJSKT9ip14r270THmFR1
Og9zevKG5K2iRn1szCNdcYQKvAU5Jkzwtx2qDlwHz4gyQClKR33y9ExQ2VtgUB+6WKlqKnfx8Pah
pTXRn3hAQ/HJqPILmGSZ454xfO9Wk/zGDlzMIDT5VXvwgEY5mFIN2hxH8XI3OYaWPwmDumkEPO00
a4MGaIGimSr8POIXyRB7broENT2Xh8PWaJyA7kg4xB76If1OIbR2P8kI9fFi0Bg+DquzTgi4ZXh0
2Uvop9DB7l4frubb4EJTJWY/QGjdweu5kj53bCI8I29XG9/NLKgR4b5CGNJOIeL1Taa3dl7xs6m+
35hXRg0xmX6YH7A426HEjRjkDk5Ls2yfo2BotgtXzlWn9EXIND+c8SvgKKhjgA7XEkHFuRIKXIRi
0HF4EjWbZnweb32SBgMwBpIwvia6bsrm7Ic5by+z5DxkBz5xMOLl4uqlxa3a67fyWO5x5ckktsl3
8SCbfxwfQHu366uiA/jQEsL2MYo5JiFP1VmgU+kqumt0ScrrxyE35IHL4Yc4g2qumzNQqIUxGyA2
A0H9GvQkRkQH2fXKdhSsqAOtbQQoX71ttyBXYt1Z+pFbQ2uyWSEYqTdZNcuD0a6tMcCLyqC+GvFV
YnGfsGcnH/NX82hv6h/gEysGgT2dMClc5qwB9Q60vSKu/sKSDvfwizY+dn+hC167KI5o2zu/OUt3
MVvxJUTZr4KZGcwLe5O6HKY6RhtIervFG65faJSH0v/JhxSz7ATq1l6ORsCpb0A/y0H9gUDJ5ng9
ii5YTyQoEQtWu02xScZHuZ3xrYwqJTbUXXXFw0pmHiH4fFwgf4mpp1ZvTk/+vKjYuS4GhOKpN6gC
InXYgQxmCgY6X2cdzNXOr9d4+4l3++odHIATM9kbabQWUGNeT6Bh7hRhaQxn/e7WFVxxRxpxKv5h
4aqFyYCbcLCU1S0aX/xSskHYdCOOMQwF2doJhFSXQnBBA3rCpLGEjolIGXzO/F+VEtOhEErPKd5W
Oxt1hQTP5Ktxsl3rwT8NtlBzDciH9+XP8vI9UftAhtDCV1r557mwK0KAxiv2E87R1ilYJKqboNlp
qBwz+3jGaUg8oFJXTAivgaQ5ZWE49fuJdXZuRCfepXyN+ehOD7JTTLmcRZhOg+aIRKjLYGBqq51K
t3ci38aphT4rej+riHQbMfav9SS2Sm6/vq3I9gKR6pQrEtmhcIUKLKqo/HrseDztlyQBzbbNzddh
ED25Ea+JM7vxTeaEG6w4IEwCbJRqlS2/j8lwGscmpLTK8KaLetYU3UBh21fCEV6I5N90FcOWWIk0
1n5wl7LVuZ4jEQb4w02T62OGTJiAN7ymFIAW8BBea7y0MTmKBhiinbG5VNZTjnNe12muNG3OE/fb
8mRZWAnDfHcqzphuvnvGMyJGPCuU8bhgR4yfnsQr2OV0/l9MPzjcMcY9ZihSpEDEiVzfvJMHLKyh
3TU33BM7pK9+MNRGJh+o5w5aeNl2KUstu1sMNGOzQDVeIRGgIzAZmjmOF9d/MjfQdC+h1CrxUDBu
ZnLeLcnnqVixy1LywPoOsvjYiVCfuisUfW//ZIKZDvTobQ6WlsSf9pzYZuinXesRpbZ6AxaybJr4
ajUBnHX3+dls7UtbC+SteqMXGPhWA0yayQFw4O5Kzl+j9RanNuuqxsaOMaVnBZ6x+9VwLbxC/33I
ydkwiDfiwOBCtEYsKdVNrsyVdFdcmx5KOIu912DbWr1W9vBB0QN6+YOkCOHtBPDv5db6Vk/Prwav
tj2suRaixOyOplS13ZKX+WylNZlpkyahontM6DaFMfNMWABsyW227re4TeM8M6t2+NCWckyiqzHA
cCL2Vdjos1OE08HDiDyNok/d57AtuJLipBmA31ECH71Q0ZLbMwewFUdwwj49P5jKR3D93Jhfxys6
0nuzcnDZAnJY+0M0NbqprFssWfGpLENEHpuFeCvX78MLwzamjppfurm0qtKIdbdrPaI293rOrkBn
jIM3LLCrj/d+1BDESGws4vk4PlunC9jZ5fNhLNEPTs1cfX9QpyjhFEIA/a+X3gwKOJnJSd5Rqtcq
HKXNSwzTd4U6Wr2o9zBK82tb8PCICly0ptbrSjsNUy/iDLxsSBVsJp3ix71wrUryq+3bE7CZOt/L
WKNwA+MHO3hApjiRkehwk23s4SHk/pOo+Ifve2DHzxZT7JCMlIj1JjiV/uR7Xsfoy8MS4m1/mNHr
q6D5DIBjDVKDuQHWB/jOOz2Jyqscuj7wqOUc68KgD8Jl6XU7X0DR8w7Ug1HhvqrKqqW1neumYhTQ
u7wBMqJehqmj/99PhclJMafGrLdZ6SdOeGww5nlpsO6LOeBBiTxgs6d6gxMR8P1q0xEYqRV6Li0O
ycANQ0buoIOAvUmUFN8cmGgDGj9R4qj+iQt5u+/gmDz+q3BVHd9+QPf3g8rkDtoiRuh1ZJ/Rwx5H
Z2dqDsrA3hbTnt2QKCF+H54RDxPvI4G0G4xQ4+L5WrxFjgLacT3RpXEFrtoLFQsi+j2l6JYKtHwq
VtzQohEl4dMza6SEJ/8znBDHur7EdfBuANpx2LDL+a3TLA2urp/X6rkWxCeE6i+rV6MFbt15QrMv
um3b7AqLKbxyb9L/Jtxyx/8HfQ/u96v125Yp1BCbot6GzAfpLtmFiNQ8xoqyHd0l9t1uj94rLfj3
N31zVjEqThWxZWeyx8yXc/hGFv019Z8AGGwfrVFP8mXuMu68U8FyykjFpAOLanN538C3TVN8nJ5J
/QqEYms120MlAJgukbqtFysYPWB8IWDvF+0R09GBo2sqNaHqzVwUhMf7dKgqNl20IEsMNyAfBMaB
q7K6+2r5TbIzHa7xmV/JGEOTrGxqakd/uuq/u4Fy0CSh3gGmJd7+xHs+/59if8WjNi1g16M/id1+
rGwLrl/29HIvnUDQ5edMZ4dc9HlvwatbKuu6CbFbKtoJL+R0zgZIaQ3Z9Hi5f4ilDudyYIdQaZ8P
pjCiiI5553v7zLFaiTztIAqnsKhvuXvvAFO6VzjFLUcXLhhA3aMAGF4PV2yYfUUYp99TqhKUvasz
KnfbCsmFG8d4R+ODed8chK/FSepVoz8e1Dr12nrkcN2YMfI+QFHzpGoFZZjEK5MJuqmP0R2x1GOH
PJ3vJpVs1ApkBfo0hEIjmMxt/HFZTms2kEji+Nb37I42ip21fHq98YIOpxeQc91dFB+P+BeEpdIw
vmbUI0/W367kojnsUFdxyqDrQ6QjGUQe0d6Q5mr5xlj/pBMJG4lqyUVcsYsnhakztr/erzOQH0e+
/tumIJNOoh6MVjBWWEJKtMU3Su1msfyoPX11WT9LmnulqpXEinB0arySobD9oQqunHsK+ao7RXtX
XmwCwBxbDeKMh6kAozeyuB4WBCdyi+3wDluyK/7CdoiTLMsY/iCBNzWNYUllPDo5I2D2JFjttkcK
xKbzozT1fadJ71ai3a6QF+yPFU4WMzg8BScdwKPzHB9eOpmSZUAK5J+Fd/xgixyCSx/EhilIAhTJ
o/jvyfkeLNSK2xE5rSp8lEiHKp/NzUDaCQ9tGYQvJwW/QmlC9rjkaoGOGZfVI2S3pfEy2KBnUTIu
s99pHusre3OFsX9TER7a8GdF72M4sHZHlmifJZj3hnYdVSai6r4f7b40yVG+XR9tMHzRoYWxcwmJ
aN+lytWvUCRwc601q2DnIjus1b3Wdq9kTVpJN33K2ARmZrkWfpGZ+/JRytV5m3yDdBHwe+dkp+qa
NBsmquaQGTCKWYgMkhrqowxvwUosgtyo+Mm4PP8pgZ6EzL0oPZI/3jd8UYGollzAmkY8RHXaBkVd
VZo6ATo9G2NLNZy/zSb0NKK6VLNxicZyNjVatIvDomeeTmMfkPWSWIQ5Jw7SjO016Fxh/lsPJElI
iBaf3iCewaDlxXVpFyt/CY9Syak4yAxpzu/5DDx/fjeOqfRxbFP692tMrBeZcQCSG43NsYW38RXI
gleixpkv1EbEuFrSeUW7vRkzouR+YF08mV8pXhwmqQpOJB8Bv3RA32PdWn6sekeiyqWXiOthX4N3
xTkvGxrh6MS3AtxpcZlaHT0yQkP/kSI+bVnz0s4Umj4jMq13WpxRjDCWUOkpNgJoFrmxdirsIT5O
lacSunaSAI5/Q7XAeuFdFeAXhP3VSj0SvJR2FRx8sFtpGqImwvJhC5GoC6jnR57oJ0g4AJ/d6JtR
43hUd7o0n+Rz0vdH1+hIna13aRDc6fEVCrvaYL042YXqbOxPOxbpQ8fBkP36yCEFSc0PObH5KOlM
YYtzoyMnQnKSU+xSytYX2YPH/x27bsjxQmEZa5Hwi9n2PMPTFDnhrFYW90J+vYkFyleg/XOJ3AUz
uBRtjIrpUr4ebJwrMVu1mOgB81Py80H23K4HEijfr+rIMQzbCQ28HFGF7Aw9xTiCsCgm/jypeSa/
e5OecgQQIJqhfb4MVuXOw6EcXtHl1dOJFbQKneYQZwvoUr9ZT1++21gufTv6SGmGO6uqzLpI3Iis
Wam9AqkD7Nt/mex/gszcd964c1514ZxRQy7k3rFOIZWa/n4AgW5uzd6N1YSS3JKuEaycyWEv4lJq
foi7kFBcjMTW4dwmCowTzMBh+MekoZzqBvYUJu51buTKEprTgmZaxHSXMwvTBjtfi4yuXYazLoGr
OTmSZ7avqSHNZExNVUCftUCH9BnVnfEIhDYH2qkJVYf+dm6sh/DTYZNemhVtMhZ6BK5uyAlp/Mb/
tm5Uv4QxifHb5EjIPiez5VbT4ls1NHEw/eKkv+5TpB3WVz8ppshrTRVPf3wJtSMkmFx2J378fspW
WL9B2ZduvLCBcQCQaGCSFYaqpWu1Y2Jj3be2dsu3KsoPzmJvOrYjT3gsDEsjjVkIntbGuN4OO7T1
8SlR8/21fmYnMHo69fGmyOJrB4ULxyfcfe8KFUrvrTMdW5j68/McnTsovakP/D1mqO3ZBxMkJ4Fd
Dg3OirKAqhWXBZpEIK/Xb+pdztF7N9LVpiATXVihmaGbpSKQCbZrVuygS5YCmASXlwIQUqZIUawX
GvaD8xyji84MzXNMie5RxUpOnynNtZ9a/pFmpo3MSIziwekjnCIi9tukoVKrmzXyqTjdCUyUGK2C
dsomBBh6OxF9n+XOfhTXusRvDOhYqTL/jV4losy+YXsEscqFyPk4F1Vv3UftdSATL4oEwOkm3ABc
mOsEBqMVl3/IgGGFlyoIxgHjg73bm5czbf6nTji5lKN168TIvrN3PTWpUQTei8pL1BvinxumE4p8
V+TWUCbT4i37NC4MfB4avmy+9LzRln7S+OHImZ+spnfw5cPgyxwMwAqtJpt8FNPftty96KvcmRjV
COJb1Rnx32QIV4KsTSRXAfjNu3yRGeTtzHiO27EUlmCrxcK0yu413Z/eYVVrMjYjBoVu3SzHL/Tr
7T+niNph9AgkXEN5xSamRRbVTRYUshA6byoc25v/RCJDAKmE1UiWqT8sHjsXKLx3zgzCXS0FKZ9v
c3mwLyK1cV+U0GWeYPEgT83ZsbLkgGqK3pFMwQq+TWjAFs3x1FVp0EL6zwkCgOLvv9BR5Ezmuj7t
GAuyKr2eSW3IiGXdmkLfyfROFY07FhlwCrVy5v7w5kg89OCC5B6g77gvQBDMTStNdOaE6HHgl0N6
Ma2CHT1Y4X9lUfpA3cGMyZboWKOfLysrDygWtIf+KdOLHjVo6zXUBaXslJX88p2I5pmL1KMywgcr
MiLuzEHYFI68/zcrK7IQv7fpUuGaQXya3APksn77X43Bp7aq09fLHPYxfsI5pqUv0et8yL1aB/6v
+GwHkQGXHPWrPoaObGrULy2TKU85szH2xC2gJBItmifoGQg81AykH/b5dBejpl/w6zisb35UZTS9
RdMjwVOl8fGX5kcTj+HtAYXEq9AMUq5H2xHhi78saacimQzj+2vHujXXlSt0q7f8JHv0d4MGRqCn
SV8ogbs/pSzncfHCuFa3dYH0QmW6t6m4sk4D7ljGNh+rw/7AkCKiRSMlxqshUg4q8uWKD9FxJdD8
uEKSYXRzX7tl201+wFLkLIB5vbTfR0ThRPTCNTLRWc3R1rjM1r8wdFazAFDS9IqOfmGZxNFkoPYk
J7vQn82nj7aulZpfpzu6Q7twt1JMBVgqB9p8GTO66sTJS0Afnf+2IT4uE4cdfthDbyRksQBI+Q/v
PEax7DC6LT2UNs8pO8Owq/mE3OCZUcQbxgHKq+3rg5Oxsflkk0IChhJ1Qe3hnt8ArPJ3mXodq0BZ
jTIMBQyKcyJPLXHC6LvrzqPhbZivLFItAs0jXJYqf7Vk/nuk+ybfLODXhioRMG2wXpg1zCzlfqNh
jWsQDoEgV+Hn/ClWRzGO8JTANqdwdnrYs1nTIbFKy7/ZtPqCklpRDYxEQoGn/PB0f8dCnMKit99b
5t7b6zD1rAa1FFfIgn8CHtqJWbF+8jD2dU3nd0uVxU3kFlKs2rEqm+9dvxEadeJZEo9/NH3pmL3B
X7RA+Ir7edL9eEQluWEPxE520G2oJQI2Ksu9QljNbV6aKxJ6N9kIncjxkL39ATbU/f65H9BRntwv
5prPLXpsnAjKq6OG2eBRkp7I6sF0xkTFKzPs7Co3YIlRuCy1i3s96daLV1bDsFqRN/p5gO3a4yUs
h0T7R2LlW0MlOdeANVlDzfDqdz+9/fXfrVaudc5svNYb2i/R21/Em5a/FtcHaW4JmVGXO29nB0NT
2JFDJUxwMl4K4plKauPZoCBVpRL88Xuf5dIVoWW5Z8p5aBZFgXgtkWXtBiW5AyYHkub2XhxDsHZm
FQwudkxwtYYz1c04UT+xM7AN+KCgEADyfKaCYBE9/XgM8MSyKI3JT/LhGhbY6G5GFALCYcXTC3yj
ALhLH/nTOobh8fbt2KqHUVaam4EcHl05F5ZwunE6di5iBudnknBtP21uIZx3QmwYKvyZLxrtlbG0
Jc6+yIYfCG1QCqOixIK+4GOvlk+hFMVZZ/Fo1qIJcNSygJNVRxJAY9GSqLOyx8T5kWZAoy/Gf6V2
uFZQUwglLCOH8I9v/TrtY//SUdoa9ysCMEUpnhHgjTwstFvhQJg8AV/GwhthBIic1/+uZ1zdgHLd
Uz9nScg+6AEiOmvBvnEDXZUi+Z04QQrjV82Njlr+fUElpaILyz+2mIceb/oI1EFpjL7UJt6J4S0u
Nhm61Fc9hWusa+K9NrXrzPyPsa5Dm1ICVvMoZGQMdxA7TmPdtSRsz+8LbRtNApn1d+iWY8UBt4sK
jQKo+Qc4vzZlBlpwj17Bg1HN0+BYgCSUaBkKsaV7jrP2LoFMw9HTJ0HZ8rnGXx4nmkDeBQIKJeiB
soFT8BXejF5pWVWpkgZGAJwbNWs5IqLxh9LmpGeYJ6qeIijKWGuUpQZiYjxe8qFGNqOXUxX+9bm3
4YUZ9KNXaENdsEBqOkOJMbI5IXOcFYaeKXLcdDy5sOgxXB/nRtBQGfct7RD7+kSKu/NyxFmyKzK3
kLgZXlHZAfeTbRbUFjaIejOEMNt257fD/JglEJvIHdpsAtfu/pZfNdevyd26IK5/Eb6LQnP1tMM9
vXVzsM0FDnU53KqDBRQqTSmoywL3a3RexTAGpiyqqDZWtO53eU2ZL15N6J5X4Tuz53TXpgX/TFTh
gER7c2aWwlEOr7XcbZw7NJOVinY8hrIThoS/IdZtBbUh1jkZ3xi3knRMCmrP1zyX/Cqj1N04mVeB
ngGGNlMqhzD8I99vHIKaUWZbQ9zdrA4yVKndQeRSjTrjnTErK8vp5PoXR7GZXHXIQhnY2CqPEgzV
Ewfe8nHP+T+jvOqxVUdUUpQ+ljYQK28lzcrn2nkGJBC8Wz7I+2wydt/WC2ZPLoZGz+fKew0cxTPo
6f6tEsONzVOty4xo+xgIsyBREYuiS/cnQr8qjKDsOzrLwc0oD4Uzfd4ND6YQmaA9av12cZlh1R3t
rcRavnZuEfifikVLwhrMgijeG0/B+82LN4dgi9Wyblja2zKq7UybG3feiC75IroS6/xZrOKg+2Nj
orKpA7XcmxFk6CsSxm76Pmlarn6JDGxg/cB4PtCDy5Hk3UM5nNuGm5CoTWWCFuUHwNBDVJXJXus5
82buacAyNvopxwLSIDIVHbP2O+3gmr4YnkRxEy5lr/OqIfoN3IotHVNfGPtz8APpJFsOsgPh7Xrx
dvhJBl9t9Y/gFWPMxdqOt1MozjZegpMoHcYjeySZ7TmBJMizs2DUAX2LDI6CwO3kTDa9rtOlwx5u
SNW9I5E8rr2SAmRtdihez9eeDwg7MUbEVHfC+rAR9tGMYzvvhfbyOvWqRf6i74W9CHF8uGJkNAPS
dULfhzv5gM/WfCMxYwerwNi/I94CP+19qYm8mdlBUeK8td8/Y4eXtmhEwpe8kqJ4dSOYEejKqD94
DiL+vqLggI3AXmxC9lfn0328NLTzRE/na0z3WNvoyihh0JgPvLgUNea7PWl+yHJvxtP0Vm0zIATg
tpu8eY+LeD/nMAhRc8LYZX/w97t1eX2R8mZVVchnbsLDaXT55Q7Tv6Pf53QSGZWvIvgLzMNApGpH
d87PiGc1Wt4arMtcV6HH3fjDl5Z7RStX4Hh0ghhU/TPQd2NktZi5PqAh3u2JjaULaqkkcScmWF4d
nnCm3hJgpqrWGKg2+8iySVADU0iV3LpnmypGSxWHaeMylnuvKi3OJDbWG9YOCVak4+FNrHm5MZSR
QoZeO1wvcvsGna2dFlo7kX+b5lRRLmCj633u2EnpSCyh+fUGIJbWa7qSCudQtBDey+x0MLtAiCbi
erQBCnIzbF6R1pAxpVFllOzSHEkucEhmuaZvJJFhOKGcfR+dwMTksqXYDs2cUjyq+35oZMB5QYcr
/GaY8SZY7t3l5720p0ZiRI5UNJACMxpxXlFfz8Lo5T45+sVIWivYcQMBfaxKv6Efha/rf4T1asn3
OqADePcNbUuagi6iDnL4RNfdB4sNGyrsKh4DzllzmC1Vz8bs8JmxLLgeAej1dpjGUTmH1jrGgpXq
uBOOFV3PWcoxgQ3grgcyz8nncI6x5CchqoOXG8THm7qt8iXQpov8KwEXVh53RTRDuGhOTJM3IXVP
yiL6FGNH+fipd+5r934+bse9CDn0HNJKOiK7TxyWisJgRTxIPf8hQ/Pbbpez9iOcxxPt+58HQakt
rF8Xl+FGMcPoXSWUvi0if28UQjGrqODWaL4qQP3UeNARlDFpGjqg8nqUM5mEGdISzhgLceaVQW+U
PqyJl1B8hxdurclsih1XSr15L8JO0DDVfufxlX+Z+NTSQlhTG+vOHnTRbRhk4BL+D3/3YnnKlVD6
SFSUKVwQQCbAQc0awAQjNpK0efa3s5AJjTMpVgbVC00WN1L2SchU2TqXBnMUK1iu+iRcXbbcRZFL
suEXRppHmkMT6UVLjLHLcWgxGFFfK1vT0QN0Aw3vvZpU/84PulIhVW+62km6ywdFVfOjbPzAWlV7
gK/nATIuYC+8k0/eoRQ2jK/3jvOGgSIztWMrBLETo/wC206Wc2tCkCp8VinW3eXWhxJv/up+OjIs
TglrkN6YGudCAecbiq1pTJL/N+PC7FrqHLWpWwuNqQNRjOB9odwmEiERDkLYtL7zyBTD/rczeI6u
7KA7ue70VSUzLcE7e7JpVvi7LY3/G1KwnwfNFSsn+rXwHgRye1BLteO/L1zAFfAFZaKCWRdoPcfI
vpgY9h9mEBXLbvojUO7shSYe2NqOqDkIX4tpQNff0BCRPSXFmWd/+I/DEl8axWN5OhvxwzE32+Mr
th8d0nDAnI81W02TY7Ug7aMa/AJDW0f2M3EtYBS6sQX2WzhBhnUAg6in+on6yTrqYMsQIjFMhPg3
hpouQ7JbeNSGJDYXbE1y7nWVJaSiqZ86vXD1IiHCYoFKcVbGaN7PvGnK91KkhaoepiuxuGizlzrV
L+P44j2bsTBqk5ut7E62VL54hQMVA1nbUdpG1RbSYJZ8qyUu3Tx/rL8Qk7peJChqEXxONNXVADn+
QYf9sEHHSZ+b8BoPCrwD7ogeVfzotEsRngtxcDjR0ryI7acEgszluUDeN9n/HReX+8uhnx4Ry7or
yOtmudFukUbnwnfPCv0PHjaJfSDIWfj/TI0N+P42ctEB12tQ3g7irKDjCDqt6jrpyb/Fz0/2YNK8
OC6Mapv+cVklgG50V3Pt1G2wgWrjDEyo45FFE8yUaBCr27ZUCN8gtXjW/Zfe8+slr2KHnwi4nj1d
IATVJV3hkuqCkCCAePUzt5RtWwmVaN0HUwD/W6RTh4lXSETwzLOI12O6Qu3DHhvs57yJsSL78h8k
BMiN3q/YIW+WSMynaWBt7BIc/cdxwmIAYjiYryZnjL7ZRUZtfIxLrBxqDtNC/t1moDOyforRzq/C
p9j1denzO6JwyshCxrQKioHlIMjSwrsipfKlzNVF31MzvRSaK5ME25E1UJYisy2hqpJ7q9JSeh1D
ptSTf8kDUJA6bgLbj6lYypyCB1QJ0c5vAAkYl8IzWOIG4HTJjCKal99YHuUPOmn9WA996haFtLmm
YNObgLyCg3uuADbVgvHNrBWSGl/oCIOvA5KExNBSi5uGWdTVb7KPP57RhMrUY3Ucvg0Kfvnugz7V
LnxhzOlm7ZSjK3ReK1Wlly1aU7p5Aqm7RM3RDvr7szW5bqx9FZ1ZqpBUDxAuP7elFVWSTAQvUt9z
DREmqcpikQnFFV/DtMO3T+0figYYzAXWxAniObmKiTfMFzkdf2bt5qw6eHaPY3VpJZ2dcI70a88w
Pvld8cYNYBavbpVr/5l9vONGiLEzSjf8SOZFbPWmnEotSLWF3WH11Tgy0af3QdoPDtYhigJlTfNd
IEax2Q+FzsnFpHnKBCYKxsSzMvPb3TxFaZzhNEMMTRJRCJPLgn8lozFi2lqAzv89RFIOSz3ssI84
6GfRd6ievuN4KnsjMZF0ITsa9CnyZpw0hipfSA6YFdAq9Z80gQ9DI7oWTv2yUikZy3rxkZPMGs+o
H4hONNVCWYmUCN4EDxX3Wyso48PHl4e/uN45SkqweYgy2KIz9FRYdXskWiKwsjn+ua1SpPAc1PZc
ocgwgT9Cn1uIgpcb0pWJyL4/DzXYyN7uxER4HkcGSQMYTPGZBv23evHUTXrxn17RQFFeLj672LL5
WwW4FvR2IiKtvVD1I5aSyr/039nwkNQGfZd9cxqPS+XcVjaIOXzRJiVLH8ogDSQ89NTR7qiE4z+6
RRMV0mDKXTOT6DaFbCKw7vzhw+1DtsDrAc74YWTTKmtYZd6SGe4KalPL4w9X+u2/UJS8NflY+N4T
nO8xowd5tDjCuLzv7b9znvH5kYlXn0tSnMlt3N25yxKhSVsujQgG3WfJU+BOAsoroRNwKPKOp7Nq
ACr0Zk87amk7RBolr1uPPfgMVgo4wpi0zNs8amYrp8YRvKeM4m1xYFqlAMZq8y/oiRm09PO2V3GQ
T1++PIbnjPsokaUiy4u/zDXCGHrW72jF/VZpvCyJpHDBBbkyXmcyNew5PID8eduwCv1Nf65L208n
PENt6Huotb2uSIMsynP1LEBIGvJUnanwnxz43WYkduA9bJH9V1Gx6/eDgl6E4eDa5c9+RGCWqsDV
ISVr7lK4glenNQUhnLdQxzRUHlRjkqAnohAkT3OoYfxqjtfhPqAz9vz0Ri5VdIhLPEU52YLyK783
sTR5vzSzR4zcWDqy5NlrUru6HuSVpExOYgx47hXR+i3yUhtT9tTKNLRjEV7zxtNY88kVUcnhSFwp
pDD9VKOf7eJS5RNwK1sbe//+WTrrIO75UjO1cHpfCMSvUo1HjfTR0azhajum6jXp+8hjoISeE5pw
MwDNtsi40fJWdlUroxWy6cZpvHI163bgz1Upl+uG6jq0Xugcg3I8pd4PFu11g+tIieT0VnW4ogo9
edvcpVUNM/oD7x7RkUnVsF4pECJD4KpJjE7b6A/ZWODaMdR+nPSYEnDQD8CUXd8oHK9q2cGiWD3m
241eDsEuzyF8uuB9am+Qp/ZKwP9PGG9WsGfEPbQTaRP/pZY1DmXE14eDrzW2i/kNNcnjAzqw3mnS
OBn6+S/E0ouXlr5jCAVaz//N4mDo+QwCFskXleg+aKuDB9529OHK6IS5YP5NlxBTG04jkbavUK2e
vr6KKO/xwAbmWRDCpP7eM51ToAh9UEVPx3Xvt6msVKaQDPt5pF/UOoJQz8v0ZD92K6Fbgx7e+o+O
hsAroVCvAZ2vRGzA0DJDDYjd7nSieMI620u8akW/JPyGqgbsxiRf/pTF9AcesGtcx+hmAH8lHj9G
LUQX0TRLD7mlkLP6p9YKoDIG9zcB5kyz2+VvY8Qfc8rbogLePOZEsq1T7rRBHU85PB/dWslmqh0Z
rVqr6gdO4fCZVoGAsq50F3Opcc4p1Mdy/gy5dCithijoFxjgi6ZVu2CUjwmCoennEeqmJlTNOChR
XuRH7xi6KHdG4P7pnO3zKmzNjzyyI57AdE7NHoJEOmu8EXIlwsYkwGkUgx1lhjoApdiZpefU8xko
VB60F4z9z0ytkefVXPSXW8uhX6Jao5VvdnWHlK/MutDHLXpTnxsw3U/wyjFvG9jykj8p5lO6H5H6
wAJIQYyqDpZkZWWRg/Ed+T8tNaT4ul2um/K0MLE35q881UhEEIfSuS162Cejr30wpYEOcpxSAJTf
QoO/FSAwmKmtwcMGqf/DyAB9pB3YyhimJgVN8AYlxUExj/vOiNo/8SVqQcg164pmuy6zBQSTK2Z2
uIEcLMkIr6alERO/04NHSeFnZ7A8MPpMVEJUr6SG4Jm5t2K8RtlF4A5ryIwRmEecPE4aDrP/3VpO
q01wdsYZY3ddy9xdrzGObTI0ZUMxW8q41KqHBi2lT0oiZMkrlrk4xtiAwbiQj5bs32Si0EtjBH+C
ru+nVl+qgNnPodtFPMMrl9E8AL/QVPTkP9ktHFGQ3vQnGTpI/bAelEoqqjUYwQtDN74WT5HgUOUN
KvjEAz+NeI6DxmjZR5wzMkU7QRYT8EpFsaQKO0Iy81ki69rv4djK5zCMd9tBri4vnh2BJ5K0aN+C
Fgj/CcMHWt/pGSJdzNwWOLM47rdzs9o4B1RBaP67J1HgAvqdoN8I2sPT6nbnfiWgm5mFshVumca1
vTAYQ8EqM8jaM5+kvZSglhupZw8tIyJxkMf1nAi3dIg53XWW+TymLayl19LDGzvCZ2bfuVTBsHYZ
Igf0+XejBOyGmcI4GUMp74/hRz99dnS/RI448iW1QDj34v6RGX51iDAAn3VWk/LpPDPgJNB5Scrv
/NPeqKNEKAzC4eag/Q/KUCxwgRImJ2DB9bXEEE8xs5V5mHLQpZmlp4ckden8BYQxyzZEz3D6hbxB
tx0v1hY+LgrVVxu1Y9kt0rQVAIPjIV/lH6/agaq+dYg73x/iEsulJnKltAc8lPMfdKKQhw9gUG5f
C7G8ElJyAQCj9GKSrdo+EukBoiPuufMjhM6D1IGKUUjS39TpWrDhScuxk9mjfGWKDaqhSY2W0o/3
35jLW3XqRRQvLXvdXebIAv7N+M43fUvmGMOK+DnOmamkWU6RKtqSXe/mMRfNab8jPwW4IMFPHRjP
MYRPkqXAOSmFIiqeXCYGL4DdYh7Ys/WsXG1xmXME60l6JxtpsZtZnxbJm9fRhXoNSLz1+yQIjnS4
ze9CEKei7rILtCK0bACtnv+IkzicuwsmGxnK89ENWpe9JfIJBxv0mhO0TT1k/4P1ZZs2TJzUhdOv
MMgEPaYszJ6yg2VvXcHZ5qjqMsdz+7LcmyW++0phSFu4RuYTwjUf7AgRC/y0pC2PaRu391oRPoZm
z65J1kGxZc8m2UojZbCwFkBh4BPpwKmHwWJLvvmyLkeu7LuqEx23/s0KPnxQeyQMx1aI10FtTrPN
fWxcDS2JyPQGKPc9+yLfYAcIVrxAVrQwydm0dKM9c0KNMTb5Q09qCz6poHtdwywtv803+9UlihQc
rMak87AdtC5uRUoUUTCm0kJkxc8E4BbNsHDTxQuJG7c4HJuNEMcsHBCW07bTv7o6EoagTIK98Wka
gbS2H4okkEg5cMHa/DhtZ8q0YHkFsJvhkXRs353RUW6eYt1sb0ia0M+RXvPF9LI/XQFU6owZXAuq
wPcaQTN2uWVtkUTnd3FetQ6+lEq+HY982JNe0wo9r54TirIA6JxHxMF4i5qJaXmwKpyM92wTEhHK
FQ0CdVKYRm1xUy92x9EafCowmUJTj/Z2ZGEJF4qen8UQ6cm7iG/EajPLk9rti2F1zeEMegAq23yJ
dtMdLVojn9OgWyxiOC5fzycFD/XzVuP5+U/iUm7pIAR/OBVIDfTUkMDb5L0rfvEYhViJTe/U/obT
l8blDqDzUSnLot6j/zAADXHa4MUlQtsl2ZNcMqvpQOVqtN+3FKUnlB+bcFcT0SXeHBW7zaAJScqq
tI6NDc9xYhIi4cyzQ4+ndpvqN3KYN2IngidSUGkUkp6/hF4w9BtOUlNXKU1di5KEunohRuJC6iXw
BH9d02UpyFjJoSoZzf1Kq1hxs/nVqIa+AEnaZPddXxr6shZaibUX8wvgClNxE9y8qnp0h4bDCfs0
zcItTtEYr9M0qobnlo0QBHHpVNg7/gm4gWXu9YNMi3p7n58tu+CVMOUUivWloUSASvZUOB6HBsqJ
CRUe1UnUL1CNUsQdLj6lj5zZCteCtFwkEx0epww0GPCw2UNoAT7QJTFjc+eB+SqrQ+D5ixFs7tfs
Tf5tWnQsnXih8pRgCrCvgx7w0RyUWNARwtwP7lFZfihlIYqNWqUivNyij6+0YHg6QJm9UutH5KMi
nRoCT5PN/QxAoOCKyUXVCv8hTj53rdsREn2ijnQ23MClHApEJXmlryW4oJXqp8U+8N2gqNWpKMpn
8nLx4OoDs2Ns6InGUcA4ocAXMlgJNoCuDqaxG8PFrwQ2j5dZAlDWVQW2NrYpXRNbPQ/mp5NLFNcg
cOany+G6ixd+0rF6zu1VbmNoEdHB9cKYyftpQTZ5ld4dHIY7aPTfErANp/FfVitrgiINR9r80344
tGFTlSilNaa02eLyGtMfUVghSoz2LJ4cDEMacq+rugGo7czU35Iw8I0fnZcg+3dyVyVw4IvlB1PM
uqlg9XqD73cnufSoy0f0p6IcXPtLD1Yeit6PJLidU7IrmrUBjBvVNAQURsBwomfkri7AXVOaq/+W
40JxcwOCbZiQa+fWlBCQ0OhTfYnVcNeMEV+FAr9JolM4nXpH8vQIZhPbsLigjowFTElYnXjJTUso
uDAB95+qWUfEF3mHihMHXVfurt71EaW7OgVAezqvFaXctshhYVKUGhbGh67wilDlD5QpZBWDRNhq
NNptxfKWLDgNRZQgCGeypNYoOVJpZACoseYqN4WGVeOhIWOtXUbXQuwBpthOdWmH5cNzzKmI2fx1
7E+5gsqbMsbXsiUDqTp86IgHXZAvk8BF8fwoxwE77FFGTWYS/j8bmQm+LZg59ylEF0SJmKYmz8H8
1zSWs9uh8sf57zXgkm7/Nv2mIGQ07nri4J1N3vGEQfK0opxxEjNHWj1lwomPl0Q3SIaYgvYTJTHm
skVOiQ6U/FYRNGMsalKLolItMLEsR4UC7II9q9fjCKlFNjClj5JDDcZjM9an3Y1Jxr0AolLFzKBY
3Y3HIGG4Zi7QoRo8/Q19Ew9Prhjle0UKX0lKVdvBUBbin+IqXXG/JMSgCnYSOsqGsjHUskfXCAQh
bUCn2F0sK3wSkL3x+Eok9aJkoXElyJGWxWCn0JON2q6D7/EmWDK2q3rp0pCB99XavjUwBIy2vevn
KwTfrqT5trN4SDZBgRtWG/JzPpJe8IYqFa2Vslc6h4Ycdjoo9aKdUkKOHJDVftW+6sf3bETB0jrt
rfqdfOtfG4mNB0XmwHv/MVqqXiazwSgOKBqzaI3nKF88cXuC+eH4hxfMA+oiF9rNH6KxKW1A+qe0
7VtAYfWDhZ+lsBoZuMxwgu3l5gqoKkf87kPksG0512B4N6jSZdUwXRU7X9wUGBemyuuPZ8c//O57
WBDCmj7PDImgvScMKJ1xhyiHVnSeWJofQ2Nc/AjO/PA81Uc75Cl+Sn+Fc++JETn2kSpX1Pf3LunY
POvQHsfRAJj0gcy1T9r8FFaWRz8jtLM2A0gOYDlVviHTTR6saUhz+Zkuy9D93SDOCZrQUv5XAIW2
5COXqzImVDPA4auR1uyih1NIl0dYKKWMo++3ar3os5dCXWJ2nsDYLIETuJvzziQPoqcrpU8ueoX2
7Gsm8Cu1jf9mFz17RP62laKGfYRDW82TCoj5FU0wlMcf4+YVr0YG6yH9MDgLIrnEvWNbUCXQYeyS
bjjNVxqJN8HJRcsh5ga2SNCr/FfllkvYm94cNXtoKp+oz1QbT84sWqsYYSQTTC2o+ia9SEUQNjJv
e4kMu6NrcsgLyAB5zZ0kQmRIpNH8MRrJBiUG9gVtU/TLXwGZe7vhmC8W4wmkAG5jliYAJthIJTcm
/3WNiuoBAtZFojlJij2/bniIx5VtlfUDuQWJCpfCdhQkqK4njdOZ6hiYrSewkUq0BipSjpOjZnim
0sWX4+0UhUHzkp3jsLMU2lMJCRDHBXG8D5riSOkuuOqz/NvriL2TqBnmBKZLkLTvmhXOFYTXwWjL
D2gqq6KF8sgebTB5tNfH/zuwRhaNjgzx7Xo7kPvejOWg3x/tNnyXohX6FcereAcfPRQdmso4mZdV
f6v4MJI7oqLPawCApgWh+Us4vvdJ8z7OvC3ersOgDpKQjLCpSbZ1Bjp0wCZ5tUAKZlj9q+7MwMIz
AFt2f/ZuVC43pfNWT2dwVYLatkqRah5gUseKDpnfI2wa+u0ZTDwOv7o2Tiirt38Y+5/AiWWFNzK+
dbNvXuTMkQuO8JBiSgsjVXKExC6rUfMNevKApf8Ro00J7YDuEgTKBxnYiS6sEsWVYOvXJ4mUgd6r
GPsJ1WILgip9mEvQZ7fxO+7RrYu8ex9qDheiaEUAgv2WStWZ235BqQnlsVr9LYjCOe7TFyLGjl5S
MPJZYfSkXOMuNtfsycbLCk8Gp/lCEMd6rboyzdMtal+TJZBmsFyVA+Ub4RxbU4gyv0LqjbyEsThO
ADF+XxtQutQji+ZcoyuPT9Md6skCaIxXKdYQ7uOUpXaxnfQDjhKEUs48fManMw7ESERp3mATD9rm
rkRsAHidzPZSF8Z4jKCUoLHnWUAV5X1vhku3IDqdGy19WsofaoOoj3YM0SBBBDGA4ZozC371px1h
rtU56/e8X9PL41lb+mhB35e3A0JykmC2pW6m9lc6Ivdw+sVKgKUVsRu7zwnO6DnwzP4nbwMKj+Wz
5dytHK7DwcUJI7ZefU3XUVM0MXg2frnjPd1X0upON9LGsU2rFAH80HyXprvW35MJjrw/qtNW9WL1
1EBTlXKFeOwaok8S7hMAcuauMfQvKzqMmvR0a30e0Z/BJR52iaLjGyTOqJjtRJiQ/y6Pw+iDJuNV
uus2KI6bAmwkucVEYCU2jQOnWmrQenfcrre0Ql2o4ZrJKjMV6a+5DTzN3DM2KTn8wfnR5EDSeKli
jRvX10DR67c5TwREh6gM7HNfPiEqRdBi99GgoMbrCKhg3mxD62qBjn1FYs+mokDS/y+2dIy3fkck
Ht1KBIgTQt/QjUTKF57MKwoSNyZ1JxjwGoOCk/MfK5gMmtAFa5/F9B3DU/X6vX7fk+WyELmFKlIt
OapuO2dz2BP73kAnJxThpGS+N/56qqb9UEYt7jLqR8GhQ6lLZQ1RAVVF+/4O/wOdeDphcVFWhnM9
bKUpnZqrOc9OKrS8VFC+cs6DbFEt4qEA80l0xwvp2SQsRrRQZ3Nn0MGAWsf6BF0Rng3qHOcT5FAL
HJmRKRSIGhUKbTCF3lvQdxkT1xs3qFzDdblEF4wXu2b/h9bbuGVX0kTDA/Ny49IXkCiEuSk8u2VB
e3craeIk4/akmHkPpv8qnRMcLU0k31lmdkawMsTAXdlDWy9A2UdSXh8tEUMVTAwYczWtRYoF+Nxc
fa/9c9cOs/e5AFYXE8pEY5qbYxbPToGk2dl/b7GEDMzCYRufuX0wJde0+AU7lAWo86rqjj3aoIu+
t+ax7AItt0B/INV0zazN6Y84hCyqKMjAPHL8Z0kH7g1NeR49NLOtqWD2uKqa+VYv/JBvb8AhMid6
+F6n5TMiO9RT9dbVq7knkjnmxUX26PRxXLo5m4OUlz6OY96xQdzfr0toxEyeDoKQ78YZ6j3n0Ebv
b0oJshMhHrdMB0VQm3HZQzNgst1v/vaDq3JE8KVfZEyundFbEv/4AGcna+FYDlUiXjdW0OljbxqQ
JAA/aHR7yAJakcwu3KY06mucmxiZriSS36varrYSvgU6cP/8b/j1q6SIAxOr7mG0O9rW50K5qT7x
FTLw7VPVnPwnnrRIjozfW5A4JLfpsL5gYtsHmCewhkVP27FXA+CA0gACugDqwLdXWW+w9wUYUaWV
dP+z6sHpXqZWbitn6VBURWiuvIg1jjwvHnrshc2Wc0zj3p31nf9xCPI6MhXdpNRMes4TqYeHsHKE
TfajvFf/3P5cRtsTu+DpTCwmxYN1mdL5bNEgFBDjyng1atH1vhNxi9xjWfN0zFRMtjA9iNd9UrLL
Hgz4laERxJHyLTL5Cvw6VElUqXEZHlK3KiSyVKEoBbPzub+i5tIGn1SF6EDnZpOaBhnJXkbMCjLq
WfmKIso8nYw/PhSFz98TonlfnXUGV55kwDTemL5MGjaOmEnkw/O0FUSkTSOzvldXjttxDPNa7Cu/
DsGg1ZAdscNNvYMsd/4HVykHAnOpYqXjDFkH9DEGy+PjwdxoOOSfvVqz6srDHSYxxra22oSULq5T
TqJBal28cxDHTKM7pREmehNOCVhsh0Eh25nPT47JMSIS9Yz6whD5qOega/wXMSDjwvs0JLp/v9qw
qdBg84A/FClHDG9utVx3Z5TduS0azTQ8FrcliiDN2nK+w1lGXsD1kxKXK+kIaqXj9iVE4BxnBnYh
gMmXS6/YY8Xg9ztgBaM5shXMsejZyRAPIwabvXGuv4/UCJBseCxIPcn12BjHdoGSWj8fpPUEM4Fs
8GkUsUIJUQjWmCrTzazBeUVUqQKHYnLQYvCsoLZBRtfTBpMnuPaCZ7rfkCAJeoLSXDvGZ8EN3L3C
wd4LSppIY2hkqnlNZXSunpWn3awlIzsz3WKb3viLsVqdrYNFyYpMd0OjwPK8aKvhWCik2bIzkUiK
ITiytLZaURKA0OcODeu2/DDKO2g/PTNnOdi7a4ZyVFDI79ESgk3sYRDYnG86IhjeCu/zRyXXp83k
XG5rCgOdyo55mSAYfgz16GYqs/W0adOiRwGztcHKIFDphYUkBgQUwbZXYvE+2fRi9UeW5m87tcQR
W2dGC0MeoVsBUMrcpi9fuq00LjlM4NJ89hWZcufLNudGiMKRsP+tgag1PqgQ+uKRb5WWvyqQBFci
Tfc+yDFPDmNsGVrYAXW31PFdxre4LdJ1ufLceLJDOaXrKmJIgbiSN4r3cPNz8u4rrQJAKeH8t/i8
/nIAvDxzpoxTvJTBOsHa1k2TZ8nQG744ytkIE7ocDHwlj3AvrEGsyOAY20nK4NjzroXt8/UwpTw7
tWyo8T7Wfw4m5jqjTpssjnIO6fO4xzrlSW4wMc4C46Xf9CtcYmLsLm7jXk890wh7xLXPltM8ykFY
bfMBYiuyxE713lXNNgRb8+v1h8R8l5tmvAfIjdxyoz4rRbtAlKkbZRYNKA3r3Qt8MnSuNTSK90xH
6G+qG+yElqHUuzBAgw5S+hZRCHxcU5IHXhymbuGBZKBgYBFhPQ3jQWo4Wg+vzSTACFPNwPYYR58U
j6C0xiFQP8YXZ87VV3rTuZh52iOGHIXpnpT5vN46sUe/0QJpp4HVO9WF6hBfqikk6GDybbm7sLnw
6iCZD2L3rLWhsooDRNIcxTmBGMTYt0qz4rBOJFGJx093RQcNWmKSUYKqCTC5H0pCRC2NmNcWwjCW
7H1AxNMnJXnM47Buv4cueN52nSI+lig8EBqS4TllaKzcPVMyu4ePpmH3T4OwjopW+ZZlZZhwIzKy
ueSV9qBbS6/36Q40u8rdTQJEUnpHe1W1SM/NrpQPm9gfHtlLTMOmxfYpwCzI4O0IIjBX6QXFQ7BB
mfv6dZgB6Lm9y5dIHGBnUHJ9YORdG0+mMIsBaqMsqNmCcB63OSoNmFB3KQ4Up9tlltwieP/5RpVm
AdbB7Oo3VhDugGf71ouU3JGertbujQGeBGAxbp1aBxS5B0hwyzzyxk86CmJnQq+dw2iTNGjJMtcW
1I7bsjk66SG3VEYPkFyHCTc1WJiTvTlT/N15PT+fJ3E9XYcZKl3XCjj+8Q6db5nxBD9OIxkDZdDa
BhvXuH3iyU6lULtUinRo3KXkmR4gZ89bAKknFVp6oXYhTOBJH3nzM0OqIU2WJhRvddrWE55Oy50L
cqHBMTnWMezo1kPFBvZQyoSxAvb0wSMvEE/c89Ul8Ry4OuYeiePRr5a8W/SFGp/K07Cwsj12mzzt
Aegs2WoBMRV6eNyxl4TSohBnDiVIa4s5Epva8Y8RapGUaFGCZLhIvRhChbwbpRWr72kHnjJFN+Hv
6008dezcxPrjPubtEA0MdLutfNYE8QYsUsEHCSQBT08LhMYgpYQRT97YAHF3B0jOVPIWe2fGOlsu
9XS3UdU2zNlH8bdNUVOzn9u4THcQGnKl5KehmGCN7RubOkASs+Smtuu6l1XkEZFsmn+zgaUizDuB
p9KCQiWkA5Ewm1svPJASA9IMjBGCdx0xXrioEjqO238oD9xio4G/qs1Ed3CvW4KhBNK0QWn5yZ5J
7CBKw+z0z7cWF6SxkykbM99sJcysm1q9bo/yIyF8QwAeBImRjO6SyyhRzhuR89mMc1inAhLj29ML
QFIS77q83Gs6ww+xHkdGQXdgkf5KF+MB8EdLH2t4qc6/c3TqygJZeTuBa+kmas+pEz0Y9qhDnwMC
2X7ADLKavo2i7030FFWkLFAatvj/bclOyJmRLxME1T6Kk2hEY7nietlTzkSPrzJGDGmBofIZOmbd
cu11PS6Lc8KdyZz4Yf5x+GnR8MuaZ9E2yMRv9KJLFXK1cX5GmrIuUSfD4KKiQkQQsglUc6aF0ilU
e+uLSE80gLk+pf5/dAXtpzdRFJuADE/UgxFTgLDPg22ogymeRQhj1/BV/+KOPzBiIcr9DJryvfaK
EujYpx2FIgEIsDD2jJeEIlSKPeHCZX8vu7LZfMERoIe/9j/StgJmsxDHQlwedByL1hOA6B0wI4hf
Guk3hnMmFiBGBjXDkQ8YZIfLleoQ/cusIPagpIBcOrIZzSZeVOqRIlvNydNoGbISO6/HibM1KPNb
CLjTs/mRWSX4+LOJmfxZ2BL6z6mp/9BCO1/D1R8/bN2oFK9QD9VgZ1kpgmGJiiNFO/UijRQQuDqu
OACQNs9CiMsaP8yrwd6JQTQMEeA1oApsMcmyCGcUdzOhs5dmPuSzeLBF7Xd89HkanHvOZzqa718E
rK0Ddbv9c2BBlXNe0YHPzeMLR3Vq5DP5uTNOcRJGx28UxYarvOAXxdQaE9hEfeNUXs+bTadZGdEb
hF8oFPBPTLNOgVm6JACvfYHGBAAdF1Sl0d4ht3LIaPXWOoyzKbdAyR0kF26Fgnd64qQA3uD+8mZC
F+JGBY7dgciPunvdRNTcyt32XjCDqAkUNdHBoEWAapStPPsbB+FvGqJCC8cHPajYNZcNaVsiotIN
3ip6PwHvdhDFj5pEjlGMV5JkWpVwls6hWxRsNRnA8MyLHuRQtm1bJn5vlS6JX/hVURRd786Zc6O4
gRPoxzQDzNHCXLhJLn46s9g4AVSYzJAGWrDUWmZMWglebAcBetrIh6o3rxeYROigaaaRxkLPvTIz
/QQutITTHmPZtypBEbKQaZ5nc4nTzVdt1vftk5qzleWALPq8B9pR9eMcnJgoQhRCxxHAVEDRgEeM
iMFngCMsTjyytJutU679frC9Xiap21pTgBzJ00zOkoILelbqU5GMabMKwC5FdPlr1P67GCHOsg5E
VhAiajY8nMZwhBHl6Q5AgP6EuyRzWd3kH/2ot3eE187R4VSjd3b4bT3LIdzMJr0bEVTsRjuzHQFH
Auqm69HSkh78WCCAQaKPVdYXnCO4Inabn60QlMqHc/JTuTQGl6SYeMrENYgcor2p+nfejSpHgYN3
HS42DK91AW/68+zEiWZ+lysEoONWeSyZJSRTEnTXXqF6IoIC4jhfkHp/qTGZXURjmlhKLOW7oMiG
RrnYjtGbO4I0oTcalSPqtRDAJILwH8PWGI1O6zdR1t50kEZAi4q0DQ7bP6p6IPsMx+zzWOffM1lg
0TP0PksfnIdVOo2/KKdGrQZLQeF3VSFy3LEpKSSWhgO+RaDOn5beFiabGRh7AK279LluqTv4UoPv
qYjD852uQA/O12NKKwcNmkdW39bsWpZpf/ULtws5LyvU34u3qTy/0zg0yGv9FfIw4+Xv/EOOS2CC
m9b86AGUZkjRATPQg1h177TB2uVQjGazA/qx1kZBJJUuB+oBu7OIfd5vkk3I/Z0IZf8vnHXj16QI
kNiDhCzt+dq6uuWzQUtX9G6AI5u8C4TKQS9jAY8rCuV/oQPyN4J5GCzhqPmBzv2Ti6ncrPGXxZPy
NSpqx1JkT4I49gjQ6ejR4snNlmRq4psGbXAItR1z5vRX7DVkTSJr1B3ELJyw15CTUwHNFQe+RJg3
u6utB1zQkosxXr9dbxlgLIIeU69nr3NsyuBfyAVUz/vDhyxuUlXHq0m9aGP/ixQRM4k39IJ8OizE
oYF5E2bToeb2ICTgR8TBP4S0Pa/RM6hzi2qXRVB2A2t0vRpGCqIcz+a8eNK89M0fB6B0jvtbaA8w
EizGY5JJYUwEQqpvzTE8ZwaRCGl0H4IDmgZxjUzttWrYnhE15MaUiwin0mmWcFgpoWEItJ3Yarfz
0fJc0d5y3qRayVYOeNip/xdzQ3NGnhq711Ch2YXef6OjQUZ25uAHhVKfm8Fpw0SPIvaX9YkgEaEc
hhgSguOrt7IfKf2B9h1NyN5Dw2FJht8KleVuZ/PfCpCrN5cUGM5wIb1zIprmxHMlWl3HcZDeYgig
8jLlcA3WwCNVyCJdbg94fbM7AQYoBlxKhiSu2q3FiwzHOVa5vOCaRlfpWlwCfs4FMRnaMrFbI8XT
y9jRQ3/NvCxob1QYt0cy4VAWyTzoRkTQO/+P/GgLxq0T26JEAHayABCreVJgspquNhxSqTJg0T57
kJhDa3U15otNCbME3iRoQLE8cRitslIP/nX7Az/QJzavvIdYk/49UwXZkfGotH8KOvoANc5m6235
HJrwE6JolDbrJpsIP7qIhcBKHbImLczL8JNLqMKg73ANYt4U4CI5QG5sPtLRG/+MLiP7ScosShy3
KTXzMFoes2lbGrPGjXOJHqALttJWcQWEYbbjwbAX34zy9bHry2qRf+EJzmGwIxog3qmMXRNKulDs
Eu8f3i9hyLqRbVfa5mofhEwAfNfclG7mdTgK5Wm2xTkxFAku4CcuyQDTGfDa9uP0QPcKa+XVjXb3
7FWW/GQ20lPTK+8TLKzek0Yneh53CsOJtYx6/fZp+xhkdqxIlqRhS+rK0iwnmGPiJkaY4Ydpu01Z
crZrGK2NKZ7iz/gohTVJuFCer0j6zPLc1dKUZrJkh5502VQgw6g4Aq5GFw72B393S4JvhZU0z+QV
fVLuOufjYf6V5CMdqrsxdl+PiFOmp5vLLiNwz+I+uz5rjnP2oAttJwVOm+UNKlCjaS8ZCmNVuKxF
XoA0PJAudE3uLp418WH7hXaoaAlQInTyer3vRF477OW6oOICm9eTlXKHVk82YFnofmvYcH69gajg
tNw8ZGcJFXnEDBvXzAq4kjuP/obJ2jMc3aKeuugYhboeTucyzf1YN3i8hhlq8jayu3iQQOI83BZ9
OgoYyxLFBSGmpUb5lA7aLVauZL3vtL5b33DwbkzGcw650xOYDUCB5wcWnOxvFWmpYRTKOSk9qRMa
UBXvmPbe7gwgnMz3nV/EKfG/QOB12ViGefaic1pxOgSbWPMVceQUfTfQN5a3sdQafQczUhokUCp8
nPNW+v37l/mquH3kXiqiNkukDP9sBdgwJa6Z7aGWt+tKO3UVQtc7Hj6KJEw52Y2Pmr/q51z7eIo8
61Tk51nSJZra6tD6QxzMPdY3T5FbzSLZKh3UMroFT5JqZ6d8MTSwoNpeqiYMmI7uoWyWvLH8Xwq2
O+Be1o8RkxRX2eGvtfNOkYmQ53Bs9Au+C6FkWNR+Au2nh1c/rrGHAPsCK+ToS1aOB3urIKtq7nwD
2kyCIriYAwJnxCosnp0k0zWmhZQkUYY9F6UtuI3LZYEyFoj7glgH9kuZ/SeRM952ivvTI8bgOzAL
Dq818P6QKq/vcEGYwTfy1f6sfg32UKRS39E0AeJvYfaHHdBDszd6NEavzAra6ObtY9XJFDbzND7S
smFFczkMhlwdELoh326s9Fp0RuGGU/3+I2G913lKgMzN5AQigO4tnF+40oPEawVxOpqE+EaOHgs7
4KUKVGY/JS1eebgJ7DimmmxgiLwWZqqkDcT16bWBi+UV1M0VyHoE/vSoF4vCJ3B34ZTts3gSLOTf
jW8Ir3w7aC82pt3rn6xY0IA5D0/qy2Cs2tGR8hefcaCluRNS7m6H5HoNo8RBfxUIQ+8P7fc3L9br
ji10J/v/qySc1kOt8pdIkXXLYztzzeoPGaanxFOMuXZ3mEPrrLYXV3o5mg9VsAszF8/gMNJc+OHD
tGuFxTg6QFiBg8Az1zlaYaAm9N/NLDwALANJ962xQAwI1Hlf4qaCFP9VoYjgK1mvddm7Leuv9Gxi
0oKpIlF96PJs0vnQa8CwxixNPmrsc3dI80kqSpWSqQPHY00cJILzXWb1J6AEwQbNZJ9NzW9OZslj
j1N8VB69uj6DkeInsiguJS6DwzitzVQi0neI55xW8LAOyUnusoamDpTtCMa3ravVuQdGxRx1/C3n
4NUcBTQKDkva7KK7ptoODdm80pXd+8HmTgqHG6O8JgKSa9ULOf2ojSbjobhZ/O54nHfoGqMXuw/f
RZDmxPZT1pgLhAXI7n1b3dcpvrlUWJZ8OnImPLwcGg7xT6JuWGtETBVqGxhffkcQwtg7YId7CzS4
CkpnoQKzQ3ch2qWBCHuA4L9syQZ2G7R2JYbfYqgmiut1c8m275+gni1FZXtmnn4H5c5fERfKPKEQ
Cvg/szESA8MoY3gzkRKlDa1RntH3fNNNmi1k1pzURTt4lc78nl7N7BxuJSoWSBO7cfLMEEEVXUPT
QB/AxEAt697e8hQXxlxRUWm68hC6lyjolreS/Cv8LulV3NfnL2jtvqERINGR9rKRgaMq3AsxZsFJ
ZQz7AtJDTFE+PGJnz29yD0we/43mJzIq5tT2STzRpbp/Psls2TzKZ/vUXrO3aJHdn+oeyyiMO6iC
AzuGI4byrRoYvjsfAMwedqftnp3lM6CEnMD4QWG6g3hvN5hUoyE4TshxDFNlvZ/pn2lDAqB3uVBW
2TB4o8+M/M1J6nX0cBmuwEGganZS23yA9pbm38frQAaDmKK38nQLbg8DN9KTx0EARpdVYYKVBm3E
3oCKthTkLKBufDJF+FOTgTzRpaaVdSFB9eCfFuasFDsYX8PNXrLdZkRrKHQfWJxPJ9h8Jt+GWp5A
VYRstyNIgsYeWA2FSISGsTdHYiyzb+/mL+n1fOXuaxkZcBd6eQmeLqeo729K+j5Z5nNuHkD65uV1
ZEQmNvd5Ce/nX/7R1UovjIHqSrQ975rqo2gu2hdhz75VixuebyIaQiv8b+PNUtL87yeRaIPQeV8B
v8Ymkw4i7p6QErOWqxpdW42BckhIJwI5tu+CR5wO7TGhNTqyYi+hJayjG6qCtjffFdXrF8ptzNr2
qSJ6OcJiTCDp5d4oFEePoXN8NsGECsoNYhCNMcbSgBeRl4/hNaGVBJx+qRMENeQMA2w6DPDPlG/v
/xjETBU8fD8Z82UOWpM72aI1YLe+7d9QYBOaBYF0eqCWAwlo2mBa2Y5+1l1VzGoFp90eN7pR9+Iq
N2qHtfEO6lhOSmCHNflEufhHO0Q/v2HShzjUp+G8af47+nRlW+pevNHLP1sQE0NSEFwLwx3awIgj
5bCwR8ni09uFLqrsq8emQ5hh/00qGeCmBNsB9smcAmWER3yWwHE/RMBKnP7aMNSZ5gKYnkdhfWBf
L4kc9+GFxpUxO41128QEsnrh0zZQ/kpwgwIJV2CovlSCUTYKxn+wuj31UnkMsVn9el5Ly5T/pxVP
dxc1Al1B/PdnDryM1/0DoBMVjf/D44aJTt5kTUe46889f7HUL3/OIgIcSy3yvDgQOAIXb7TTfRoZ
o2lxbyAXkolzupE1RQUxFARQsIIl58udge4CgFwHgZUoJIOtBTpnGwZ28QOw8+u6m6p81GCrySji
iaiDb5/NNKtHxm+BWBSRQgNXd7Ok/iTB83ZF3AYAQsE2+TD2fBDRcKKApiwoOsN4MxBkYTDDMpYY
Lk0Rk8rQ5nr2bKOpzwR3I2R0FMBJHPKXf/kyrCfmb9QpmXzDbFS+JeqTjnsQo1Sh0JrDcCyorDit
8p/F8sLcx6tKcMiGjeAnVKlRc9A/HNHu5jWROGQu9LRS4Z/QJPm4C+eH0Y6vzlzOv0l5H52DiTP8
H2LQ17o8LXT+0zqv4nKZu0SMVC6aqk48nU1TUnztdwDhzHqlZUe/3U4gMB6KT9VhF+BCqc4jxxFM
RSyOJJjQAISRgQNJiSapY8B3eViiGpwosvan/qH+kEqtfv30jXWuGdrOtig1xGo0LM5zm11Q3vSL
T+qDFoqbf/KIe0/eSzYfOgTCors9/C25XB+M2U2Lg030qxdJBBoCXnveXL+l/1z61jzMac9KrC1q
Ch1X/xbdqVuohJ0Wb8QU2tySjaoP1pxdZcDLY2gzDFt9FWonYqc/UBH78GP16IAZXLilckMgpBam
+qWzspVtuG/1gAALlysIl1dVEAJEcc4RuHizCZctSrGew464IMqFrkM4bwxfpQG5ZlQm1FKlJRCo
sS7pbd7lXg+ZcAW9ABETRJJ26Ku+8wLD8mV8f9GTdIM7iSR4mRiTtBg8Y4nvH4PaMmQE64FMUokK
4TB5ZfbxKRkGgaVSH0IV+eWg4FdVVs5wtUgotUhLGfjZ+uiz72L4qRTYuiwOYx7fi4PFnXhhbe2B
UZlN6EjZAcdBWYHJQAsFqm+TOz1uvdZalJJBccoE+F3SkalMaRVeKfqqMe0L2XMQLYOkRCz2ePCu
EsoyNOcUYKJDMeI5T/WafkkNtFy4J35eV0BZrYoxeshDfPwlN8I3BZjK4BwdpJuN8QopVF9vNXq7
YkP3wZd8uLtQrnqV54IuUK07b/8jNa8V122G3AZ8QbfV2p7UFhYwpHsW20jOACVbLw/xElHe/lOn
ZKFxEz8uJiXHlg21YXg51eSBB+sMAY7XiTisbRuktJx9oXRDmQVQqlxGAIFrM+i9+IVw0E/mf65b
Q2zO4jB11fyN5TSy9V0odNTUGlvQNMCqU7AVN15CNgYhx7FCqIkG6B77BQ8XFvue/ITFAQjDf0rh
/VxeDoeZfRUaLUsnCcjvLs0MmXwgM1pxgkR8V37gi0spGeL7osN2EgJqtDdbDZPOdKWXjkSOUoSA
b1VxbiV16V8/ZMaPgkwgW+EeJxO7JHGX/5pCGkbBbnctrp8kmTuG/Y835uEm+6bDoaAT6Wz+quau
6PIOvL3IvcVflIobClfyC2GD5br5G9ZjtuzmfCU4dlTI8/qpvZypn8SYTjIhF9UnqPLjeNum8d7j
XXiurt6DGJF3rxPjsNYRmZklZzT8ZuFc63d9qf2pZOa08aznJVvrujCSN6E2f4EjrqIMGH21Expk
o8E9fwKyhphTKMefNgcwT20fnX8TOYn2hsfMgbg9c3fKtvi5vl1SLcuQ1r6fDY962Qp4jIB7mpFd
U73NbR/VC8/72gsMm5vkHGYFsGVUjUPHjJ4F3I1XI4S9AC5gUGX8QeYFzvzEkr/M6fsSqqdb/vVZ
0XaE00TRTyDwUznPHbpPQNZ3FLgKKVzmfF4arDEiVeQpBZfB3nqI2/6+Ey+0RU8z2+aD9HTpdH4M
aTY7yBtcaZs21iO8fhqNkR7rBViTU0WxHRtaOmwGxzEYYjV8gWAnOm0jYZKc7O//dRZyIWA2gLxj
MTL4B1NtPffdlKFkGRy7iJE2t57YtYDjjpT0+Jdli4iR5zWgf+l9xt77qiJlupklLH4yA5Q27e+o
djJqIWTRNUmSAS1XeIxiih+bJXyUPYAyH9z0YABZM1C/Xmu9r6x2RaSj4C8LzME//LIWcztNWOJD
TCm+lEN/FHFxvyCg7JwwRMKnXDPn37mzOi8rQrcXOn92gkuznM6maKSRnFQ36/IL0/Nlezfs0PsG
2NaoMmCDiA4PClFKPEI/kNnD+H/mWFtnYja6hKHGk+Hu2sfrt2zmCbUVrTRuCSYgZ+8ZF3PWZXIN
8vKySMaYb64Z0jL85lb9gyvdHbJ0qQ4sKgUxc+smwhhA6RgmEJ5drtrNg3yyzg2nz6t2DeajXBvJ
VGtoyN+bjcMuQnFL1bult1kfAKLwtrwuPQNrWNW3f4S7H7UGyDFmxz7Ac/dbOyq8iPURSm0vV8sD
UTqGUDQ21blvuMz/ExGa90FvcN0n6eq5RWDMIg5kOoiodzBYrEpMUXPbE+wlOC3O5GGdxMBr7Yn2
sr3mKTT4R71d3pvPk21Hq1H448NeJ0FLSiXo8NiuGnpWGGz4NlYtZ9zmc210pK9qXngJigKezSIM
g42cdzOOuv55IicPp7d0zxlPiFLOlhdX1kjwJeWPfeX1ZgJDt4QDFlMl82zjNjRngOe831k5cGyv
KO6xF4yBjqD9CcG6QizUP5kqRY5MI/JsdH0/kb70TyHThTJZ2pzpBWrncDBBoA96Lt4c2tPjY01q
76eJbbg1Rk6wpkPk26ehiJv0CNDiEvToVtzDyHe1wAcU0smbT5qiy85vXurXbdHXKjn/ZXj9XzDs
luNi3CynljJbjWSZUVM77HWrzdUevxhjXgko0ApIDY+MsZPWDU8NnTJpMiDtJO2NaexgFhF5HAhU
CKUYVei5Wv/IMwRrMGYxXchIJXxE/sVbFRwyAnShSnXULtTgZOCTkyMoe3MeO9hglug1Dd2ZOnGk
ur2Qj2GTkxMZTMZGyn2Bdq88P8N3mOLrPEg2sJNzSv5Ii8W0E0KtDIipTkIB+j3HMCCija1X02Vz
6g3zCdPgh3/N8pQHOVNqaDZ7t4+lVh7alj1uBsXEeV+wtSX3xXpcLqLZqGPt2qeu3Y3R/OQy8wsf
/EP8kLov2jdY82rdna5RhWBaPk/QGB65CKEzhkvsh6jvh50lXdD6NL7p3wBTjXd70aWm0qTBB/TR
PhSC8VhdhwOAVqRSh3NpWTBlLANWEBaDx1D2fMWXBvLFGkmbg2dTEg2g2scF+MYKwuzkJBlVhRjW
qEuvwSHdtjKJOQ4iFynSPpV3nYQybTd/2U3pw3gGqDJvnU/p7eWSrTyUQw1V28l2TjXBOV3sppDB
hf8Un78At/R42PXHPk3V6P074KmAtGMpID5KxWBhRha41M+t3y1s83+XQFRDJwlc63DRWaZeDZ2N
UpWgfOlPWFzjI8cxhpg2fa3ccdky2L2wYFCpuk1VFtngSQnIytflLTuPBvTnThIQlwdXD8FJy91B
3jsDkj712Ubavqbrtg0Pmu1uvoo7jjcirfWM6LynK5RJclj/U+Q6LUA9PSgjESSf4PFo6ZroyRJE
ynRg20A4+WdVxPzkUSJR44M71m50muyHpug+YyirwMfsJnXS1hRG5OOiaEw9QTyBE6qWRDaJzYMr
wxPEsVPCx3DeHQ9GuBZfo9NvCcoGtz7d5Vhm/1KF4q+7RxT3OONI/bRiJBN3BZJXGF0/7uDdALaL
1M+Mf6600E2+N3hXxzLa/6xLbZWhWP7cgJP0C98bx+OfQE4DWeRVSLoreZK3jZZvKKk+KOG8+Dxj
Zdbgo1E3YAYZlIJ//H0B/f/1fwEIC4szyPo6ZeQSL81kGim5vaIoo3ZS6nCvwAl0rwTvESz4I56a
D+ij7BOBng6MDS5DMaRNV0w63D7RdHqBGWIkadC/aw2FBdCEctE3AjcSP16iULm5t7FVE8rh+DXT
/LaFEOQA2ddtucWTnLeOAYtYv6LNkB+xQ7yp8X/c1ZYxGVMkMpZyZB3GOncJQwq1SJ3detoNTk/6
/pnAlLnEg+eZnXNU06QBsETsXzWWDo7zqW2Ayc3F8Ukb4e3sMalom3vHJNB5bDHxPYv/Pakn5ytM
l+6ZsZyxRn/jzXbbizRZC0Ii3m2HAjtdHx4UBOKR6tPwIk7HOgndwWaCTjs2oRrRNf7bQgQhEunr
F7SuQg1XytUnz/rIjlB4zytrmDEYJPvA3T6ApZY6OJw1p22B6FiMfcTQtxQo1QK+kt3fAc61/ZfR
7AHZCdYgGJyhgUISsbk20+EZORubS2VszqwqrUtXXe9X/2oDFw122vS6pCkvKy4hCwm3B80EiI1K
PGdsNP76OraUP0A8rBy2uMLBJv4Omx/Rr6jQAjS7az8xXZYgTqqTLm50+PUWj5X63yBCGsTjfru+
AILuMEWHFh7LwOt+7qJkMHOpc5J+fmpzQaz9nzVZo57J0SrmtTKYSXyjTOOLyz7uWzzh8cAxJtGA
g8H3NgkocbknfsQFA/R+G9oGVr78gbixwPg3fOw1wi0bLCqKJ774zIEgQFr6SjCgTekwrwLbE27B
iylJX1a2IeKOujJmWNY/leyocnLfU8RY0PQYRcuiaeBeG1bf6IOPwNookRpDGKwawdZ6/JbtAacO
1JcWD6YQhuT6szoAbSPVqbNelbYqHAGQ0r5pW8yoHw3Eus9ORcgkd49QD2/oEXeoGn1me5afAIXm
qTy0aHa2ztT8Xrq+XJdoMYLvk7H3eVBFWmRS3knm84cj8AofoyADXl+P9pb8WM1ThR7wc1n13IGF
1sZ60NFrd/HFjfxWILvvimey3uC+qMV1S1wFQANpbvn1KtFLIeM9ozemDcGZDBrrcQHF88k/5ZHK
zf9nFfwJBYy48g1K1lb5pfGxw+393nbDLNcTYmOURQRKZNj6wXLayIrU/LV0ZGBfl+urumoZlkWB
fN8ZA0ajIQH7VJmf01oew7koOjAtYo/PL16NvNn/hSRYVFekm4O22HKESlvgX81keaOeLPoSSPvM
PD7I+IzJ5OV4g17mcxk46cVB8qzk14az2+1V4Z+16BqHC+7h9Dk9k2uNyhtwITeUog2nwRH6B2eA
kUL/zu03+80cMlzxPSATbvKsB2dq8YdcFTF84CrWKl4nfCeCsv64ixBso6h7f/Jtj/tnzKSFenpG
pC1RwyEmObZiPOOt/MCdQxOz3LelSCAeXbIWUJ6e2Tvet5KHIGSx+oQHFOhsdpO6JmOUcL6TLyfV
9DOS4FT/CHEWk+0wAPLBqlyO1UmUA9QhrbML0yT/EqNYRetNaJ8OegIam+MJXEs+2WKD8YXqmFRF
xpfAsIWUDbCeJ/ZeWFoyf3ZXYFTFZ/b7YXJMIlW9eKxT0kh1OaKrLp49UcBtCTloE5VGsXa4Mddb
Z/o2lsqmLCVsMsijWo000oPlOmREK39M+lapbrFN2y5c1C6p2oG54Mc52IFAOmXwVymykRFMedBV
spYlzXOooRbLxtjIpj86nojW2U1qEsGsfoDWF4l0N3onouUM7qZzFxqr4WxtzXzIm5UEaVeU83z7
aP30rzDmRuPf8A+fK9O6lj/+hnk2Lbf6mUdiE3zE9FDwFLDpFDfxtJDms0stTrsa/Xlz0ek9qxiM
sUXT8+ApG1SKQiZ/6eIOE0yliiS60bTn8hk9z0gQNvGAkC2sEMga+vVXhlvF5dUeUSNdvjL+hXV5
9qo7b4wEACb2Ht58s83pFh/J7G/BYdvaUEfd/s6rsxQSeJnr887qPnqP1A6C3K8l1jW1yhdGJSTn
wfcxLN0FdH3ZWvoPvaqkYJjrue/tcQUDJrJURBlsCofeC7dGax6VcLerribqMuOX9SbY2wt5B0yy
7dbFRdKXSk55KgliUnQAFPZ6iwzy9VptJSbp3wTtVi6cLwJqMgRToPlYaZx+P4UbaMWm41h7YRdV
wrZIPC7h4JZP4x6dYI2IRkUGy4QD8Bu2A0xtrSnJNAm/faqo6QTy0JTeKJvbE0/078NgES+Y5p4R
p9eFUUhVg3xfzcTXVl+IQefT2tGpOs5MTcEcvaOO7TMUHXoVSD58FSAyMiJS7ux/1A1Q6n7EhNvg
N6+Xhd1GjpuHtk6jVOswvlpXYUYNiifpVQp32/rkHcg56SOf0WNnb2lk2mzHOmvC0LI5uQAbhzo3
wkZuBRyIH7K1cUUwJmACvOXVRHAjCLtd6xUdaRXmL+OVFtgDrzguQR/VqQiSEeCQ6f1tNNeEGaTT
ZfhUtqxA88ftWgAbUj2fsFIOuetDE8BWwAiGZXfE7t3Iao48+Ux0ipv+1TJ0Jo0ZmMQgQDHm5Okv
GXrzA/8cNHQo7fYPZCZfuXV5Z1KYjqjVMLezuownYNYCt/fqE8xuYiTVVi4SmQJkKSdsxPFUH4xj
ol0aNtOkY6ylUhBorV5kurOM+zzBT+mKyf3W41o0rfO+Tku5oHlf7NaO1YG0kR8lJqePNEvUU6q1
tJro6/cdau71BHPHUVDO0g8q1nNx7zGI/ak0908goWuy7IK/bo4fPuiCwMd4aVedVy8GkAG8eRfj
fORSlLTjBRRVIVVdkXhcs/Ui8t0R1yd/5STwI1aIlN9GtwRIThnoH7UHbv5ZtezF6YpmtyZfd9/W
jRk0HOpKFWz7qBpSRbI1rMEO1KNuDtGk0iStgATRAfzC/ZNeI2PLVD/G8eC1Pxd9e3P5BkQLi3My
cwAa0hlaRKW3CKAkiIdvAmIhdbTGuAlRehZnjzj/FxjCFuBDEi5YmaQAmlWzZaaf3l0+T80aW1om
OOXG75+efFYAfOX4nMva8TmF5AOKFdzjq7eYe5o/zeDBrg03UM9pb9Z59n+vWsCae025iCFW+qIv
atfElu4DLNfyEalIqsbSVhm748u75NEhYgDu2MPJt09MCJlljXUwQ7dOMlDo7G9K0o1PvRqc6rLh
3x/YlyF0VsxqPuuqjGjqRUHg/oWjDQjAEpUdm5a7z6xFnXWG3rOZbfFm+W9bR3dYORW3u02kmF0z
f70y57+3VKXgQ32/3UOPjJ3CbzptgQbbTa+WukGontMf/bNf6gPX6GFxtirZaIzC18h418tdDWRb
R6ey1cS9zwP9OK+srhTW3BD51cCkQ8TIhTo/729TkA/ic34HD0L833/eX4DnAmD5a0FCoEC+Crzn
77e1nX1XjgfseXzfsxsoVpsAI0OSwnuhbHTvs/JJSBmFzWJHbe3LX2A006pwqIXBasErAJ8P9Jd2
AGgiBy9YtGFW5q2jEy6tv0iKicosssbItMUqLTVYgxJX6xbeT5leVnhjEBCV/QXcJhcv1vwYhwvg
UNqnD9Y5qSD48PkspAq8Vo1i0/+YxT01TT7HfR1WiwUJVoxjAe+r7/kwh+KQiYl7M8qx2s6x/Y+j
kgDgdobEL4940xB9CdFHsZMdrx4dSRhalMzV3QS+UlE3w0/ORMnZrbcfpthHPE4fJKnAArqDHQZ2
bZ8mjG4F7YFcGyzuuwl0/VLKRDnSkmI4oVv5FvW/mmQC52rnVM1sja8vqm2QzJbOA2gcaOXfVSqp
pCUPeonKsUXt14Eiiui3ofsfxk4+jusj4wPKAZL/R0b+RkEXV6OER8giUQGR4BdF/xrqKdoMCUR8
QvHWfLKDYVqXHyOWuFXuJbP4o6YeCZ5bx34p+1HtJKne+m/nU9VxmGMaGfxMAGxpDkIZzO+bvP9G
aRBd8Ll/a0E9vN2sqE7M061fr5eO46J/HWM88WqNiJQCDqN+/qMA2RyaII0SJC+gcEVtVIPd2WBZ
Mkww7gE63snKLONX1fNLEzRggiC+5Z6KvwuUtKgcTcAntNcMyTM2NSFAdZ5tMCsFGgnxQSw7yTI6
VD0PGWQZtYsTMt7eyrM7pvIRy29TCnn8rR445mZ491zftw8C+NNsmGfrAwP2zxjiakl/1oGZB4wE
CPRO5Au8i5OVi3hztf0jQ3MYjRpYEUFQEq3gABKwbRHwWG+pGQUmoyg+dMYtOIxIu6lXgYK85VAu
x9HwQ++5zL7XJ05etddcmIea7N2873G2Zo5KIhUEcFf2QKpdkTyPUlcxZVEXfMVuKxgRm9klR9XD
Yrx0csa3l3EzZmkh/NV4arAlu43gAWp5BM3CfygNaLn8e5IReSU//zAh7ti9O2HdybN6q29PgTnb
/KulX/2EW+FCRpXQ4xSBQJtv3lZw1//6lnk5BE9sNQfazp5qWDl0Yx0F1iut8WrbQNbjFwcxQ/fG
CExuRYkJYJvLilQED0cw5VCRiSgGi4558TZOSOjx3R7JKid1QqbbFvDry8fnQqGfJeVHy/dnyl0o
jTkvKgfRewVJHL1XerSpxbXMSROP2y/+X7CXXsU6as4Ide7Ku/DdedHr8O9sOqub1J6b+uVhl5lP
JBQi51IGH8FiFUL3WR/jPWDDCtOZKQaOE479/hrKmQ6OlYBcsdWDshZ2qm3Af8i/mIWd68Qgz07m
zvf5rArkVaIldq+JpDG4mWeKlSxAgbSon/qByhbyn2K67uZvsj3xpcjyrs8hKGKGrlhrXBOtgfdy
/8W/pt4jvU8CGEFV+UzY1xsUE6MilEQh185g6jPx/LErUtjkEkP7XhKTYO1euUWXvggLkoOVWj7a
X2uTvXw5grMNQMRHjaV226RJXuOQvfFtRo4k5Y23HBVcAb8nDMQxuh2xdsFBU0OxGrK0JxXnHQyc
ln1h+Wuhs9NHr2rgkPLBQ2mqy8GTmDjDuw/Hwmzg3PdGS6xyOAIU1HQZymETfi/OLM8jmX1i3/6J
AoeA+D/s884b+AGwsVmHew4Ikrrj2zjeDK9IdWISOHcA0E+yvcX6W6dbqIGzrsjOKsOQoMPAZC69
nwUFEVvhlB8iLhWRi5OizfYiVwcdTlDVzmep/TecYNbvToMpwobhu2aYN44TZ+jFhdG0roZJ96/z
tZ/w4/tx4dCi8K4YY9bRZiXhxhALZrilqLSzrHqU0ZE96SYxOpmkc2tyZW8GneJynzW1ORREcguz
lBj3VLC2VtW60jobM5jwCi436p9k2BRRUDDiQKvff9SUDc8S+GMZQF27Y8GVOJiXVe8WDFNTCTSq
M2DeFp47l66OxVssfR2GGli9RjrS9afjlqoJ+XzgwmoJPup4sbF0Mq5A/PrKbwSqR5rITUeRf90r
5ijTdOctDampJqIqSF1xePmqnaQ1WAiWhqFnQvmH5kq7roKfXUZZW4FNATOdA8/1OCGZPJF5+gQy
7hXTxAVxCvdtvu30AVRdrAtDkFOzU54MQQMmTqqmGRXl+0UY0hSNsTZuJ7m/dkQUb6wOue56poTP
4RduszsG9JWa5sEZz25JEgkN1oM5kMMKx160dliS6WyVl3eMeKmCwk6kNdJ2+X4+PKlIhVxdD2vW
3c0KaXSFc/KJ0phv4qpIxHQVoAhA8m22VXyaLukPRnCLffUKal/Z1T83Z+u8j83R2izY3LUWaMBM
tGolxUlqHmD2DOo42+Ukej6th2WRAvR14hMgVe4gOLoQc0G3HFg001+Y0vtv2vuzhS7Au4HQuF6g
xLElEEFPStSInfNl3WN9mB0uLrNSK6T7Yd+74QjCU8VhLm2AazlEi1oqUY/NW9l6t35dKaaFZbYH
viirN76cyKNdQ2yhdra6Zeay07KYcGWjcbnLmO7261RPtTbzFGsJw+1gnQNVvtoeBbZbl1bUQbFn
n3vH0uNjvBhCPO46j9J/NDYBepLcbxIARkbv+FpA007gTAkKMwx228InODtZl4peCAt39dGd8Pkg
pPMK9eMCe6HDrhBrUE3gQuZSHMyYk10GrwXH0lQrF6atNcpUej5FxGrhJ9uLkGyvSodCIBDzLbXv
l+jgcFNHz05EzkshcVH5mWTfGoNXcopQ9j/sUKlw2lXfDU/FGVWOfzoGlfwj7Zcd/VWWjtV8SFO+
vbkAZj17Yx6M3HWdY8tHqTNwA3Z3DrGtWjtwrgwT3nRbTn5ABzhygNnWGeUPURX7qvEteaop/7QF
2aTg8ucpD+J5uM3NoR21ZBVVwbO9w0E3i9jtcFL1imdjwt/0nV98lgoM5c1FCHiz6juSI1qbkcoe
CLxofmXApTTzn5MiDJNR3rXdBLdBWqGfs5ZVMMLQZPnvEtGP7H83XBJ+1zCgfJmoxoIvdPhRe+td
2EBS4EzgUGnDa+luh03+568jUr1S3ED9r0NaJwtT0b8PV46BovirAXCmwNqBj6Odpur/MrhykxFx
TL6jgon2zqan6udZ5ViCXnrysppPfPTqn21qUuSDXvChHIanz10VGx/fhgp447I1XUqU/SmzaIz0
vq/z9QFXi23gnmgocABWYaFJl4k1htkGgMNl6GM9SLyMdsbvv9luQLFYuzXwA1OFp8aELKQF9lDg
uECMhBBgDp2I+vun5KeaMSzhW9ZwCXQLzcEx1lFY8gGI1QruCMNLQiKQpuiZ87jFL7pmd8vAzHV4
CBcuvZ+MXfYMbko83iDW8nWbiBULZR2a1WqO49S1llxyTDYSVTa9DF6Y9uLZAgAYi1fzo0JbG2Ft
qX39N/252oJ7pBzhlwkfp3y0N1Z5bD+4UhWoS2MKGvTODr7utvPDe1TZ1t13YN7+C8HTL8pCSMId
04K2/YLAX6WA3U8BrpDiHHnp1atfrI8OqiGEpmJh/9cJNKs9GqW8U9P8qgmzeEkj7zQui2XTcnCx
p6+AzSvRbCAln8mNbDu3/8oGiNkChUMFB6fpQJIkdxhGUOqzZMECKpsNPJIlx2OzQIzsMI6yMegT
Qc6GH4QwB0KPfqPPJWj2ndnKVUgZGzxoSrFuvaVoBUoQEWtw9uMa6bAwcT9c4ZG6fdSuafxH3eNo
nF/4jfHR+aDeb27+gklcZ+mkM2vDx09gCxs7N7adJTteKUQyDQFH++Bkk4Qy0aEzhU+KE+8kNP2u
k61M1X8+FxYI/V3zwZcBKgMGuabJTuqRfslSrkid7DOlAhJmE9FEGfzJpucaaxNZG9R4VyQTwCR2
F7KKEo5hfbJ7PxmMjfy9wCdtox3xlFVdYJGbfuYgw78LPArAEv2aLUJqVKfZCODDE20Ccm88RPNV
V7suiymI5MXSpJPzTYRozli2m6epcfPXysNIif0xRlWekTQixXwXhKKgMxLHXKwQy1IWsWtY25JL
Ya7wsaaQG9ppMsUuqUM0CzGOX5l8ieJHn3kOWl9+BuVaQesZ0tA9gDxZRCzaWJ9xCeUyZTQPfV4Z
gwgnif4ghd7Mgfbnic9ceSbaiMwLeUoiS61cBoi08T+k26VGBsEX9KVGgZxYl0weHkHB/MLIOYtB
7iXWI0Xq6WNNPhoed/lgkFzMM2xhJuYq2fVG0WIPn9EHi7xpkNsEl2nBR8IHZN1dQaDkM51qxj+x
p8iDuWJNvu/bFnXKGuHLeFXdNg4g5JToxcZTQHhD6vlR9VcgADg2m4evrMrlZVSDYbwlO8kRawMy
5bEwhWnFPeFKA6eL+GBejVqXj4LBC+VynVpqmmN4dSHf+sxYBUNRHKHMPwldvk6i/CuCxcosBP6b
RQ8c/uzLDy2bEfAI6yjBKwIjEtMIHONk1sdCN/fpnzrowFPc5ygZfzYQwif/K6HjYGiLpVDZGw/l
/hGeeE0M659wPvL34NHr4BVaATImHEbsMJCLrbXmSSj0KmTZJsiJyTX52mhQ+dOko8l5FxdXzevq
CvLy4sqBqtp8YaRaeSyQYfjjQOypnW1WEgLdpWRSr5IMNTSf1mM1AfYXmjGdK/6RXxQeDUVguXZr
Kwq0Tp1mAXpbtEBbCG2AN7G742tA1WP5dWwdHZrvcJ7+eoSkGTUrCpoO+1BRLeukEI6HubLFHcRh
yCTaSQg8Js/MsmfjWjEvBouDwxQ8yxOU+xhRmll8WKsG2GBOXtEWqzVw7gMDwJB3XPrNLdhdyfTS
jCmudM2bxB9Rk9Tr9/jQcSiCwLJkAcJCjXYQxlB88B1WYcFu8Dpj5By6F6Xf4/91i9gGNYCLl9Ue
eOCIBPR1hy593u0qRJ5iat7El7p4XVbZtuTsreDHAHO6V8cAHS7unFxO55LKGZbPtFJAfpf8TLGx
FIqAAgbU+MF4jJHGVvNvyMtgl9mZPL6i5czu6aAB3dZmzaH1HAOPGa7yXMb90+7UeOy2ir2igV8E
7cc64IZktr8sTCkbyeNl3vVJD8IHoCeYhhfLljS4iOfdutZliwfzT1eG8Smmj5V94xVIEOg2/6Dr
YwarSeJPJjcbnlaENCaUQWRJJzix+cRLp2nacy6+SBp41K9P5ukxJWqV9CiTt2AqlVYEL1iZABCg
kNTtQhoF7j/4+8JYyGy3traLB4IoaxBvDQWbRUXrhx6gGqLVJOJ11AqURT18RF365tAKbdcqLhRH
gq7DVBhEEc2LvL8zx/pMJedr4NBOHaKEwky11bpFDim3EVTaLgGjJYdq7fBd2GUBVXq3KAPDCfF8
KS9W/AnXmLIBJuFaVz0ILqMFaxQHJnWBLB4Oim6wzC430h/vu2gfWQsmR/efvhAstzeXHuPgTThs
QWOlKI2RC9WMJf0in3SCIXS4Z9jUKtKjV3XvfgD2Ui6cikzh3oDdi/kZqhJ3cjtm6CASIa2BI4hz
li207TFQNNIKjMEIIcZCjQbPPEFl/BUjflFaorjmfC0JMf+bSHOTFIbi0IMzupQ4+dKM+LuQiZ4E
s8CcvU6P7dhxpVVGRJ6YNGR7r6jG8lpF1qtBHbsCZte2gEyMfmJKjuN+SgR22j3+txaEnkul+LOJ
hB8/gug4XYmpJVxmzvJCODkoeLecJo22hV3uQ16FvrE3NZ32Z54O2kzQ9jwIS8RCjFIv9gFxcSr2
l4Ohpt1+SnCZSW+migHaEunmbbvfUsXwa0+SwaiCLFsPWCqhZkz3KQB1TIEeRoHuQVqDlBfyfzJW
RISvjYvPX0drkITVZ4/T5hsX+NSudJpDckTt6qDCa01zU1TdKjL9ZW3TsrxPpNkhD4Qusu5pf7cv
+PuuyL4Cnv0X++ChpMbm+a6tMJXM+KapyvbgPSj1xLOychf0SDGFhzT8Vi3JxUuniEAveofRIOb3
kq1G+jzB9CfnkygPkr/KI8mj/YBxZ/h74+XWFOkB4WCfAjQLE7V9EC3h4uAw5z5OdcMnTJfgQtXl
aKYIdlvZP64rTsEO3l7iY+bFIcSxiTK64y6eXn/Fiz9iGwtsArALLXN0A5/XbZRqW/lPOKqG5u0A
dXRsLHgdPodou1LqW/g1F6jbORgdGWXcxmqN4ZufNf2homNTh2JLBiq0cfKp7B02sMvbkhEz3jPF
Av4D6wjrtPxzVaBZhA5TLI4iPtROjtWa3T6sl7apSVIVYaRQY9ab0W5DB5SMV1fW3t0CMxVH62X/
vVAFGQSWVW25gNZU3y+F1A6XOh7eDNRdvZrbeEftdms1hFWjhvM1CPum9iNZ1TYvZXT4RHgRs+uQ
2QxPHtjwj3qEzxEW16luNIZg4zyRWSHPCPkiR9XVnmHf/sLzsyZQXtfNcxJBErMf7FvTBfxbakgk
VlSxsPl1kRrYMNM2btLeF5a2lRtuRioWh4wmNdurd3hLWEocVDuAFRxfEHYbq3u84vubDYg9KYhz
9IjxrRMq3/qM/VdrVJRd8oF3c2Dl0sOwYGkjfgph9Yw86fvrzAYTwTnHIDPzcsdW7spvnTWrbpUN
9ZCm5ilVb1KtQoXl8N3ZGcaTvPVn2xnf9AY1EdmnmjoqynJ9B76NyrgEJ6XoZppEq1/ig1Le9npE
XsNzAe42ogKB4vMnNVUXXVg6D9NlkqtJsEDDlbCy5Hcf1bXvYFXmtOX8DWTYCfWewNQofewIv6wG
3ctAldWyPLkb47CeQg7njbFItHsZk5ESkD2ZJ1zl+8s/d2o+LR1ia04hlaonIRApwTpsusUoEwBz
9nqvr57C68PhgAVwvuWi9RKWhYyJtJ6VmyeEuazynrlLQhEPYPEVBNMgYahj6PKQ0Dx0UM4focKI
308hW3oE0MQPi0BGzAhzSj8v1oX3V4f78f4KHmdcb8WDJ2wGDqAA11XbsVtMLI63E044+bacT15/
kUZQriZoIBRX+44Bi0bXxSjbfodnMoqUPBfj9M3Mg1xQrOTc7QOQdh2oNUE5Wt+g2vBUYTOh/LL3
KnAhOxgysfBuAFgP2+X7mgG4g2hRk+N5RRwCESD/X+jUIn7csggSkt4PgiiU+T/5PuLj3r8qAapu
lLng5Y0vwTuF58/E/YQYwxNmHqXJ+SKKPMlIM+SmMcVTj2dtUNSvTa5L+7buNZMQaxWgNQSjGaXS
+t3ErjWJyiuQkSvphIj5Vtk9rtEMH8u2MfC1eBagcBftjS4CJdP8laNmHn9SUzOHU6zBrEYHcO1q
Wh2SrnaSO4ZyTevYwR6mNNNBeMB6Xf3nW282EhhpTPlBwvDv//9pR1xNeL1tWQ5M7uQ071Yy4i90
815IELC5iI8Hivbk9YtQYp0/n3WJblp6rQUH/CXAw7EETdtf+QnYffGndYx8oupcdn4p6iC8yxaU
Sf0bglKDyY2UjJOBBMCzRv36FEWshMasNhPUWYPL0wq9EWGGVzYiDB7LTP6+6JkXo5DYc0x+IDb9
qUtyO0a3wa1h0LV0oRgjZEYi8XL8y1G7cu2L1FXOz0IiZCWSu+8cJASWXSRbX94CYxykmCT7z2Lb
+3IbRPuST7jzvmImdRR3DCmbD0NxYqTe2+GVeU/IpOm9+bTKvlOtwZT0GMZqDu1lE8oC+MnHMLnG
cb64EyUx1edm6Llf4pdLFxLfeNP4uFlDtYDyUlNpDB/ayFilAmNy1zezmnpzuGhPY3GFgQPXFd8X
DCj2Ux1fHdamNniOPhRSvkH3v7ZD+lifDsfj0aApXAj9mnKd+Zn9e85a50LI3sf+5XnzQc/B1Ok7
AizYhyUmvyWJrHgjwln/ceGdO0+TB4kUc74oJF3bL10IgzUfb/B2dDuELQ8AkRzbe1jzo+JR1eNt
eE6wI0oYt0jWThOFV+P9/btJl3jNDg70kaPvb/5VcLRBoS0K3hJixQTFNI5IJ3EvRTjbb+tuwW09
j+n2pyAAopaW0mbILdSTdKpNlvooEGVmbHO5UGNudw/sCUM+pK3urMNbLDkQ/TaX5zCofqpU+UBc
opZBgDIDsBFETthtcEDOnRXL5Tcm6TbPPmuQhp5ugA6NxjiZs0XqgSiJ4enwpwNXz1PyTl74/gV4
r5O++sL6/jWZFqpaEPNLSFwm/J93vhoeumWRCqzBstVIKEHy8GZD0u54XwK8syOk10q6jeTHFV6H
Hd7YCw44512TNSJ3FN/yYIEwG9sJyZ5MsNbm0po2pS0zhFMgwX2emJyGkkEWMkrVc2TLV/vgm+js
G8cTQKR2ziKN4fFjB7hA/qXSb+CoSZ8dTSvpvwOWVZCMrX+s4bYCSm0OuMvAkfKPLoGGoEucxUTY
yXdz1TO2wAQAzWWJj9mLmL7W8jluf+s9PXUfOc1vlhau/o5dgiPHhiXNkEcKddp/dlzhBTF3iBbt
NVgSFQ2z+bGJAmiteaatrmkgmbCzAGir1b0mlR+th1X4SnuZIWxZIqNSOOCUJapq3hfdgTKxESqc
a3zPR7bY+IPdqChtT0knSfmsJHcxf13ouKgRmfP0FWsldqu6bnzDfTKGaoDqI6NaAhw+CLc8GXwe
/oHOtHID9uGMaw2kvB07idAXBmPb+6bmsZLG9f5Yc+2lDO7SSP8TUwXrDt8Qr8Fqb1mPY/D8twmd
qVaP6ZOGJkrPptxJQL8FOu4epn+fNtV9NjCgjUkKYNz8ncr/fRoWk7m8FO6q1DTtl4RKbYt0Bcgm
U+7kt29CZlqDdch8OFDDFi3S05p1NV4mauaRYi08jvQJSO1Z8Z5qke6LM+Br2irtvAq2TTS/sXJ1
FbdpssUTfQkL1LugSDKWHrne2FXormDcHOq0IMiOot605GKZjjMg4S5D4/jIg3bMzHPAl5oUWslO
0vvHbLa9XgDTDgoiNWGa1AB5BQ+vk1F7oFEJAclTRaait6Mj+7187ujE07ItHos01irqY1y2CE4c
1IYH17MJ0iySw2GJMo8gig2FZz7bdPMfb50/crLEASHD+pNGQITxNjrPpeme39p1602QHH5EBipd
xl/r9ozEq9jsXY6BJLuG4O8mqV0e+/aQ8QGlUUox+zUI59JleMQqvLVm1nUfbwN7MShzYf3Bzegr
VFcqDZv+LXRQnoCKlajvZfLgMr0gE0sONjha90fRaIwalnHiwdYk/FbiV65yiZs2XLE1CZ65iATH
Z2d+uJhCKsAIhwgIWz4g6PPxgy+z41W5GRT2QulWTzYMTdp6WYhrj8VOOyCnge5fF5CI1cyX/W8D
pHHTyOCNDQyc7oxSHqNpOIOC4l8Wgu1PjHj0hiKRgRhNF0JrFDIpaeSfMP5YoemROxCPfASCfFLP
X4FqqysuKSqBmnu2kprEcfCGpKIENi/uGaPWj5J+hovj+bBssIOXABP9jyae4iMHdzq0v+ffPQyb
doeLuPISkHvrQeJ2g2j7sVtHXmFem/umH5xzcKy2vNR63q7mCACzAy8OLkJQtFximzsorCiN+pGp
bKc6MFwCtXjotzd6UUE6yYyLD/OBniCXaF5RaFvKilInyTH3yFT62SARqFR++zJEOPbQmH0Fz9Mc
AKRvrdUU1GwJkw+jwymeudKQIIZUrYTQ4tbYcoDbmZ1N3zrVutSNgywBovoiVBANAnu4zyby1J4G
fABCWyHEwPGxktI0dLPJECGBuVd0RP7GuWHBjwkHIQPUV4QXUolhZXFMmc/ETKA+PqhKbSzSQP+b
rHDiZc0nrrhKMwuT4j25DOfWjVgEZXwnE/AzmfkCfw3yqnR/kzVvfApqvA65mVUi7My6BRgUHtg6
eZNtlebuVITDacHSScCasQGI9Go/ZRoxmebqWcw1ZbRnWXbY9vDNU1Vi86GYIh40D/x41imoQm+V
S2EMbWr3CKQV1rl7LlSdBdDruI9nFYrMXzlpAdINnM8BQ4CWNAx/O0ljBCVWHyj6WbN6jEQa7buX
ZKI9w4DxqjR9Tt3JzgUquv2Z4xopG/3jHrziw2hURldzQE7TwTY6/tXv4iTYsrZ5CfCZ4gTH8g3p
4yZ5ViNUgagcW1AwMa5wHeIhDxs49DSMzP/llEU/pd37hBwH7MYjdlhzX0swf6zeu2fkDsjMj0q1
w+cWZIdqXDGa4rhUJjjJxi8TPPJZzd/DpD/VOvTmAG4i3Nq9gQVIhDPLPKryt9pXv7l+W7PloO+1
5SBkLDZzMdcghHrHOBB+F2K8c/5C32DEgxZR8OdGuhjyIWv50AN65fuVuR6CitXt0qF6HzBIVic5
+NfNgSyZde+ulI0sYUICJ30Pt5qvUPJwpUsreJaUJfW2q2F8TG4lI8C30mhAeBtVIh9KLAIbII3w
7h1b/rOr6opEnG/bbCgX2wrTIvaHtWQJcPku4ezvYN2YrqMC5GKBG28v65hfphNn84MmtB21ppqm
oB8Sk3j0YBxAO7cq0d/kEhHdRTJIZ2NKd6z/REAfpeVkG3SMoe5y/TsV97yhYEWqI/akMXLcLpql
i77aET9VTSKmdQztVdqkyRDBPMXdWe5yvet1rz48I1r9Z3XMvKXIteZ0HQN0LYdW5Aof4ZEsI24W
W6jLPDjiK4DmL46sETzRw2PYpYtLfGXDuXxlMjGvwAg+KYWxahEkTDmyl98lW6yD+kLkyTp8vX6p
a/Fso4Zc3QsAq/5nxCP/vNpPEpPEARGVjiw5CMxS7eSlGTegWnpSm9vyV33b+0qK62PW6NsCnFQY
LqjXfi2bV3yNAd3E/0tFEWxf6Y0PH0LSAwWsDzqjEbTknGjukfSxccUCgLYS82JtRYY244X3iUB4
Ed5Yubocw50IuD3VrJCSRCNbA394GTW6r2UAuUrkJFfyaTnWWkyBTGu0ovzxhdkhvxGkxpTJ1CaF
3QPZ9frw4A4YWnkQu2oxQjsoTGhtyy/PU2s9Xd+aovoZZewK6uSSZ1io4PWW3rUzK9Ov4vzAoVKA
+9N7seVOaWew6BjvPnl0QvBGVq15BmHxHf4KGUybku8hiH0tgZsufAf10NHI2fIw7m2qF/35cVDW
T+UgMVoN8RnVk67Mt6sjZTMbi4JdNAY/qf5E3nHaXmNhvzLgOJZd9QWdftq3Lar2NfaPxtEMtDDB
yA/NaQNsQjTulXmTs6COAomhizfUKAG5Fr5wIH9t2xxz6jq7ho1ve4Oe3MaK/ElB/DRoU/+f9MdD
X753qjDyC8cstvnyf9jBf1MmAS46TAyNPAL9RJxnqC9dCAlUMenvgBM9ekjuKSh315pxxUnMboab
fjC640gjE115gPhO93Yf3BcvQsJERyVcrpCxg8y3nqHfLvkonw8fqFHFkev6eFQe3gDB/3x0lzQ/
T9wEaHixDjTFie2JiYrvRTUZapy3ji/3x9X9UulAPdsDCj3lL8BiPDYrX1YLvUig2Lgz7sOQRNwk
ZXJv1Ep4gAsuhwGSwRpGul18iY1SlkwSNzVCTuSIy90MKMfY8kjBV09wRKtB7aUNH7IRXB88I6mY
wteTRacGsc5FkwypSWzuF5Gh8AE7xJJHiIzsid1I5LLpXMEoblx6KOseHx3R40bhtjami1MAzLjO
0DJ59+gibQQtykSNyyfHdfNUCOfOr/friYK+MbKwhM3DNuHvUzkiyoT/ITMC1mZxpOAl/uRyDIeE
u38Ceizrk7UDErxGSA+1XWOV4ZY1IDs/qACv8T40x1LKdqwRygMzD0JzYh1OCLgqDldHJ41GOWp1
/LL7Ik5R7LG9vhakmUuiNnjnMaWVPoaJDUzTXB9r068bje5lBHqS5enl2nfksT/YEl6Kpw+weFxX
UYJEfTCLrRT51tnAD5Guz1qKVXxsUg8oNsxcFp2SJ8U0qn74bLyXmP2XF/z7SZQSA3lOzT+JV9sn
uErzisMpeEvM7hPfjrKa80DFTPtNbU8qXpMyl5pBg9NCr12Ot/y+B7jyZHT4Mb3qBzf+h/8Aaqao
xcOSYnsc097/ePBaUe7M891lWhC4CyItVXOq4gP/ncEsVaZYhejf8buCYN9RTrl+3DrtQuxN4AUk
ZdmLjJhibnZZytWg28aBmli+ro2JEwyYYWb6qkmDYU8VR95heY0mSK7CWeTXbVwdLuk5B93klgSD
aUEb28I7G7xjmU4dHw4tfEiwaMl8iSvDkm/HR7RZnGir6fSGn+q3iG6AuwIGwDRlHFrsDMmsaXzp
wTI6U77kuGXYUPmTeL4hRBBMOSHZI0g1xtIoBBZ6HIo2K4ovSJFaj1RWIO1Ic0vQ6iGomjGYTowt
lw86nX20+dgnUR4pI9U7djrd978jlX4mLbUg15ZyPOa0nOQBjkusaUpgXzoyIHBZzKSY8POtndTG
pThHzTENmtYJwxt75C2qohCVlWQ38zoXshDuXK8dDkQuOswHcR/08Q2tXBpMWES72wJs5UEsiYB+
g3TwRb1n9yHkifbz9Ak9KypZ9pYwmc1wshWgl6Jd84NH0KtGZxc6viQmSy2sktRhtijyFg7GibgJ
S/OMT5AC7BxrIry6xSLpH6G+vDJtYI/9LANCvTjuwmHM426M7WOl5GitbiaMWgoqxzhTlNvs67i8
DqZ+zyv25LT6q7p51JLFWy6oMbQgQfMmvTnaCC1Yy3tCgMjJYRlsYwi4iOzyO3O3GfuzEChpzN5g
FMgJ32axbgWaHrSlrsrxiExn4El8xEEjhoNLnd0HdRVz8PyRvvdQiKDxMsJtFTqHT1rnsxVJhh6K
h2uBZ6gimxv1d6p3kahjJ8q57AKwU3hEfB2jCGlB3yHHorH10EyVJDlka4b4dO0XCqMyfN0OX2ZH
DMSD8vpi/TgjJk4zThdvVMrCdqecWAeqwzKzLHYtVK8qzqpLEFnwH38CwcGZvcsbLmrXLqf4ZshI
gBoa+GeM1fLhZrmjXVdmnkeQDawuB9PumdQTtSWcSsRyIphxdg41hp6XKIaMYGS7YQbBbfp0jSNu
OShGqWfHXBIWBu4AM+KxHrlT29zOeP0EXGikDxofaOwP/ZFR1fB8/J+8W9WcJDmxVfV9KhKeUWGk
BNMRbZR6GYCMHDteOCsZH5KothIoGqpoAwr//9CvLcrAnt0u3qZpUiTT3y8crETR4Rqz9x0WgBuw
7lPFWL9+FWCzQZX/SN6RHKJ8GsOHB2Uk2YFKeeiba6+lcvJZRwaMdLc5dT5vwPjMVyLua+cGIWHL
u1jnkHV3UNr+arYd7QlP5UFUYEn26gJv9sl3lkn4dPK2eQLXn6hLRM4Ic/yIDw6sqRchlsM4/Jul
pWd89llZeixM54w8ah2ZoTSP7yofeHh3lDpOA9GQpk9BrjNp/J5X8Qa8gKLbhz/uHK9EjN1ybHSu
Fh8lngIgj6DuELPd7IbYY8rEej0tmE7sKnz0hapOQSskAFheLJhvYNcksxPiu9jvT1/k2Refc6bq
q8S5Mbjxc0xgxERXPHx9gk+IeQcGAW9LyexwqiGTwZq/3BwTPKeopS0dOMQPwcoVyB0rKrBq6s3p
SQNt10fup8XsBITl7PlBEM0A+Ob8EnqKuJ5X53dPaQjJnllBnlhuwkZjourkAoVn60v9pMELlIn0
Ph2q+f/IIkqkhzWBef9HEnOonxbJogKscNgGoXgq6Azm3uaq/sSfZJA3Y1AA89tedlFrXRwV2pCQ
vPHrH3/c3kFbjJi/FbFGozRBIWdzLGiWajnexiEK8Gv4grocfbOgBdB98ckegIAOHQ17Sn7cW5so
KpGnT0lTdITPC7n9AP92o847SrWCw5qGV2LVFesj1+Tkt4HtbTaXtCufsuKzzEIeoB2B0taDwYTd
D00QIOnZQvi+YKhrZtoWeYaAexjkbSsXipdJosxLqphvGwgHGvWIPkhnKuOZb5Pz/dvUkfCVuHI7
7Fsnjp08TgSGu9kFFrNDQHhMSbvSXLsbPVfEOyQnZLeEjh4qSkJV+/k2QPCJ5P9GugqviJUkRx/H
kM/v4ebhctOY4ydtICHqE/0PBuquOgDR+srx4zi37uzwATZEJYDWrXHXfu6sgkRiFOzIkXfrIKmF
RUAKiRQST3TSIf8CQRwwABPcFdjIthlw+VvVKdZIPQ+8kIgmhuZN4epPTovusWquMM7dv+yKTwf2
v9PvoHKeOB+qtvbPY3yHG8K0n9hNjRyDZQlf151Viy/d6O/a099gpThc7TU8rQVZc/5pDIk7KF1U
o2ziBYbfkldoqSPWkXUrZ3OzkXrVSP0OQ2nOlP4fMVjFxGLqTFLgPe9Ux/W5grTc8E6jmC/K323Q
Y7lsaTEl/pEGnbb80LYXrO46wBNToDSJcW1xjIx3kp1tEW//QsQLKT3g9a+5gnjN/uXjYkTdXYG9
vApQWH2tS7aL7Jfagp5Nw2JgP1mtkcygSQXV1ABFzWoOcgt9R0Z+03HT64irgQgWP4Q+M8DaNj6M
ugLx5kNw6EAbPUjVsfFvdINagp3quNehrbL4mU+GR/SQbXLTaZ9TM5tTQ98WAjpehq/2ANiAxDDU
UPCI4akHmfQ7xxdbs3czAfQEB/wK+LrHSd8r/+e4c8ya2kwgevo/OoSoes6x9TTu0HxS+zYqq5S+
EYmMKVvl3pypBciAa3DJX4lKKOg0JRnZyYH4yQKqB6kE1+dxZXWZMzXXczZK1g/YDc3YzykkhOa3
PRpmD6vSdq4Z6bAhUd4A1ieODL6q4E3ZTMHlb+pYS0JZ2/50rFLSV0SjIvwdsroXsul541oat7Je
enZOTJHEbPBB6B3C10lyl+aoQxlpqfEYs54a5oKEYHF+bNjRsSGnZ+qfSUoT2bwx5gGWer9k6DGf
mWrGq2CFZQ9+yAL9rq+MBPxbZEDr4XoOzhJaOC/TlJTumCCeK4/kD9vB0cNcZ/LGbSyNwTcWPFaB
KX1uGNg/HLZABbPp4i2RpeHFhPA2WAbXLDP1yoJUidZnQ7lj266dnb/SFK7ZKK0AO40p4Un3s4zT
jNNghDcmQ6ekOQTZnaGc6NTZFMkJnQp8i1i+9GcNQCN9l/XtJ6oEmsE6N00Yaz34rBLPeKAgJsDA
ld/H312w9YRjyc/L2eXmWvwOdxj6chSXLujT3yCR29Fm7mkSjZVGxc/MiqAFNCXeE7u7x1GbadmC
8+84ixKecPNp1BlN0kFJ0ivxv+atzbJi9f5m0dD1U0AUVYI+vwfHXtPwquPfGwGl2rKvt4Xe3Hhm
rO4KGkVwEdu2Ev+/EsIeR/1Z0IOtkXIouEAt12NWNVUuAmnasimdDlzQQe5PHucAV8108JDQuVB4
t/igj5Do8ai1n93GpqVesAMGg7z0l49cSGhIWOK6RT9CnwM5f9tiBsOnXoKBCtn8YBkiJNIYC27P
0dK/vnimY6iuhlsGqZsKqlWHAZpE4IUaRHaQi5bDTfp3vLe0rb8Jm+PyBPP+Tx9yV2KmsjvqgMF5
Ypa0a2bKXZqaBHjyK9LGsA/e4hSKQ/0zj9YLclyJfEIaIznrjz3P5FtOXhrq8kgQGuH8V4QXTuru
G0G2+IJutw7vUp6Du0g+qj2oX67yV40pKZfJqH1CFevWTWt5LY5LGqYLn0zvv6+Hc2W9/XVIxC1C
DXq9bOaYByc8A/hECrPAxhSioaI2h+i3WqlDE8Oa72SOKxU9Ad+JE+k8QdTtGJJLME/M4pHnq4/m
EBZPQKohhCpEi1W7fbJlXK9t4kVTg873leJSNaamEw6UKSK0d8sOhBqfIG46373kJwK/O6wrHt6b
Yv/sqWo6l88xj9WRp1rTOGyP/YLSM39Sdw7fOkZvmmRYa/AmT4yFEFtxZDXTXNEfA149CaS4yRLp
XQ1eGIDDDzhnq0RtHR9ykvzH1G8e3XzKZ8km66N4KX9J+USs4lUjsk7BzXgQSe3d73k09n7r1tzs
GE+BMQm3trVOPwLaWuLbgiJQj2Wzf/Iz+rAH28HNCPjKGX6akD32cgnZ94n/waP4t8Dp8yCos6Og
Nv1l+eg9IM89A347Pxrfr+sg2n4YRwauDwMcnYQenF0gyntAq+3cvUHAoVYNhVqRWtGOikPl1RwP
+Gq/oqo0o6ZXM26PYeIZrObOXSRNmYLslqNewpUyv/U2i/emWoIyTdx5SzqrrWka2MPmfwTeLDKs
aeBrA5gU0aOdB6mcvqCDMN/jJThOZUy500Ahz4d+BQUAYusfVG6GPhmtmlejs6KlM8LtfVCTLYwB
PaK6MX6ICclozhtcQqZ+dUehtYtkhEdXPJMDAJIGsVR3rpYjt+zwNBZGG5cBmT6qx2Vo+4Twzqr+
ilO3X8zNPfFpy4CWLQMZfyJxT5nqamiTCcNP3xzDQFRbRqblbKNjDBx/QvoY0nWI819JB+DxZlEj
S1NE9wDANfpgKRQx0aXlQt6raIRf9ILzf0Qbqxh4uyO1Au6Z3SZ0SUZJtNiXemdldKxMv9jPFQLz
3azdQ/vM1/kojxRoC4r6vGmZGL6HIVnMnkgAchlJFacTOUETx63MxvG7NGqeOsB240cPk15zAfvQ
K7ah2YVTGaugaFLz12qCZOP2gN+/pZuq5934i0vsTD74uj7CplLoOsjQAyvfi0PFdyZtpCEorvnP
KjHdmLBQQFELUHVAcveClShrGzenv9AYGIdUfOMb2SWhlSybiKzr2TLMzM9e2U1Lqpj+jt3Dle06
66CQYdBTNzwJqVSpSk2I6NaB7vWtKNuARweQVtoehjaBFw6x6gBJ2Cx2ZHZLiFH0vfrMka7wnTsi
keITmL/wZa4mfQZhdTcCxNvi0BhKzeh4lcDKgtEsv76wtVF6EagLukywKzaxY8crIIqTmK26fgdX
24OsCbGeMBUtQ84qq22Gg0D7dOlyg9C9cv32lmoyxSFQ+jQL6sNMUKPvmVLvjcRhaUsX2pibWyku
748bJJ7WGpZNaVtcMEDM8xoatfPFok7bw/f9dMRKJsJtoCbnf/BCuAWeyBu8uz0kCbG3mifK7PLu
0S3k8ZCjSMU5hI7lCCHI24oaneuUAEHjtrsXqI4LhM4GLwHhBSb9x66+Kd9AdhNkI7rtIK22EO5U
VEu0XT8zheEabvdes4eK2ATO2pWa93nzyPvXc192rHCB4tZ54ctKLnLrY617e+fhVXFaLGa27NfI
qfiaWA5qnSU/N/YDJv6b40EqQndYe4tgTg7rtL3UBlgjpocv7AEd57sLgGTmMU77CcUpgK4Ky/1l
ZpC0OEgSVSz0SiBEu3m5fDFDTfcHm1qqw2gkIkRACW3pOOc8v7S+Hb29X+qee/PhOGSWfac+Rj+Z
/+/1Rxufa5oLJC6y4EGWdcDjKsdpYTpaCbHMXjkkxeKMdViIuVAJ+c6vN0Z8p7L775bcug+m7zT3
Ee6Ib7apvmWEe/gBXriAav/lMns+fPCM/XrXuxxFjt5tybLhNCW6mjcPsGaPvQa9OJ8qRy0s4IGx
dVr9QoNNu6TxhX9gWPVnyEqT3LTEFMf+nK0uoznbWaWFui8WZDEocboijcyJV54meMYsFHXse/TU
CfmI48i0KOfui9xcmXsPsZn42Koaw3PAgOIz3eyVX+PBg07ZtQjZxxU8ttdqwvUp/5aV58VZtuyy
kI9f1DcJE5OSmWLSXR50SIfPYNBtFRRDUV4GWjJ+pmyS5maDWE2ekY9s9xYxPvJBG6gcsKV0N2IR
OmYHXnfgj/8S5IwrwSzlKx9Hdlf5ur2kChhfBS3fef2JBYo9ZZ6tyLxeC+ip+pzvrETkc9qVrJmi
qTXtgdouvbZutgF2oev2uGsBf6SPQuiPM16VI6oLROwq9mEDPgGTX3JtBHMvVnrwJV4oTfPS69OU
OYOsvNlOkvqrrdUUSMEdgU0YGFw8AHZV82cT6uESjveisKBbNMqnrIoJeBewupvSZy4yMAjmKW08
/Ntmo9dm6C2KaU0RaBddym8Yfoi0D4AXttrQQQqqUbX1ZdMvTWTuyAPNorfaIJpdO16Mg+xM75GL
U8MN3ZK28yRn9nmFdt5yEuWkQkH8RhDESquydxQkFYie5CCWUF4/eOX6McPJtaVjjRDVGhzSfdAV
3FAaZ5RTnh3XinaY+UZPb3JEXMuIkzMKaePytOEuayZWbr48/GxFB5Vso8tlg8wlZE6pshMxHNQQ
hUDgUgj4Wxl3xvlKVvytRohbtuYFieQv0+VkO32hQJKWqMzmXlbyo/9ThP5c4FOptAMKZcNEapq+
YcRQXKK4gBgFjp3kAKzw5DDacOr90L+xhZaHZVQdd10Et0Z20Kvhrxddsiyg26G2djNtwCONyfmc
2wbUI3ySygETtagH0fNikuGq7gCSZPfF26LwOIsI9QgvS/JJI9UoJAOQl6y/Gpn3uRZH/aa3UxIs
IrG0aquVsfZveiWGYGT1cHHrjpuQEvFT61X7CUajbtWhBbCpakzwypD4mBjUMFZG/tAv+IM/SmLc
rQ/OlujYPROWD0g4RsyEbxU/KOa1ecZ4qaRk4mVVZKCnNy5E7Z1TKGfeoQLbxjCa5JUrnEmoLN76
p5ryuggi+0eZRDkTU3uXKUZlnYSfR0UAhR2mGrbSvArAQP4mWF0xyd7plV1mQnV3CTN/q4pSVJ7J
FJk59UrlF00w6u0If45ftU/CwiFFXhJgJvqvUIOGSoUpzhhzB3QqEWSid085UURg7AvXyQiuYpq+
3ZAzFbqMIptbzIQuOB1+3SYSrK12Ua0McDpnfXhhQepXfz4JT7W7HrQ7a5ZkCuuMVniTZN5wHCub
CXQt2is8bJU25spF53kS4M0KgLqSkT7ULILti2yOf32AvHxsWmy0LgVcWVI217cyyJZpKdNBM3Qk
lEkHXjOEkyVmvdL2cXD9zzEPLtEjpzkECtrb/ED7GVO9R5P/HuMnf4MFmImnZbQeb3yJskMIYO/P
FZiF7raaOjWc/ll9FIbPDRzWleAhCqYOH82mYDzjqEEC+cQ4sYG2wfWoN2hft/349Biarq6fy+tj
uBHfJ2VGBMpgsZ3RWSIS/FfCnGUGdmgGZo9CQJxUFL5+34nHgLiaVA5Bk7PR2yMDvG/RHGXe5v3E
YoZJVgwZkLFBsKJifG6NHuiw+lBkpht/SskM5WdRwPBpdy7K6Q6qTrUd6aOyCssr2lyWqUsdjQb8
oZzra/x1IoaUsEcjmh2EbY//j/4o1DveGvPxum7yvVrh2BujUdhC/+R2c6eZSWhQzq1t09CVvDge
toEQEWo/e45vvGOkLLFV+6jkO7Sy9K+JPtwPqJZeTMbpSYFk3S058jCDqN55YTAFRSm+ZqVGlXQi
ZMTSFQ21DK4zm5hGRmok14BVncH1K7pQPTV5p293UgJ/cVZ+T+ixUFKH27/O/+pW2m4QSUG88cmN
hvc/v0Qh80HFVd0LTKr4+uLW8dO2FqzwVE3mfVaDAMQVuoun6cRtW+1TtjobAkV6IuxKSObgWlxp
ko21lWQxMNZstJX+yD7jCpQITX80VZZ+pfvhJzJGCrR+LtoIO39Y9nwHoaDnWKY/pBFoiYMCleia
Dqmnexe8yRyqgDw2940tzJ/VRj8w8e3F/Sp/Io5yCNa7CBMCtvzzfKYoGnDmNkQmxp58D+LqUhBx
aTNpIqicC7+VCX/MjO5EuyKzPlmXWiEVpm5CilJrFHliaEQrOtz8ije3TDpoyBC0jFq7PHoTJ82w
eWLUJ6q5fcmZzQ8ZxSgauv6Xm67qCwJM2S1z/b06zBMNab1yjOu60eHjwuSELJ6rLzbMf6CdxxXK
AAya8CcQwff9F4aawO/iKWhoRiHrBdunKHFp/5t8mWTTEQrbf7PwYLLJbeoDtqLXk8FC/NPDn3hL
0wfcrU9ewDg3OWmJ/e9cFlnFmLioANFovBRK+4C46tsylaMVKcDNhj7fOMqj97PHWfIrfFSFFMmD
gzhiVjHjwd5jJ6ib1pgW46vRvfghFy39CnuIA2chbOj7zZDhSaVs29bhQ698jd/wHiq5Z8SPEV4X
WVlxjjDOXmFS4vxYGTdIiwJVEaziD55476Abkmk1+zBhoWbJ4eP15yFFssGPC3jOp9KIkHwuNa4e
jUbBLgJNpnbuBDw5lDipniSMOSQee8Y2FOnyM7v5gtvFZUVtOQX08eiC2kE8NseU1vzgr+q/SN5i
zjrEFEHHLLMjTU8epyXyrMcEyLBWAcYciQOHCzxZISr4JkX4hk5V7gM9bL4J5VJDlviGIY4Ruxdz
1k7Hpv/nAzxayU4xUbrFB765xCzz7hyr/PND+AWl37tP/EWw0fXTZD5i+VmKMkE4IZTDgW7NV7ih
ZKFtqXBLJtghM2uNT/Y4aUrEHzxteBdxtxEWmRxWwftdjPa9QA5vEPpB4yqF2oitee5Bwume3yD2
DgKWIOXDH9/jMjMK6Cc2Rg0SGksmj3IpqGQButPzaM9a6kCPnBINqF/i2msj3hHL0Y8ja4c9abD0
SkDVuEH8rZAsOz4f6Q0zWkJnOG6kYRsl7IlkH5NT61FtVT5GCTmmp+f0f7/m1OMTImP76mTIRB8U
GtAXwAnpFr79ApdEYHQdd4F0UX7su3MbbXg7h+EaQ1gfU5U44v//305rq/pc9jKY8QZ8G9+ITT9t
wEikQWaUkaMCov5bmMqEs8OCJ8PIvz6pO+ZE3SwVqCZbwNsg/6efibJ2dKHQyLqVc/X4aoPCTLwx
eniUgUWqZO4hMENqmnHoI5XAs5o92o+PiEGfJAFTHlVwpNqr3DhS/qlO/49j40QpYXRPhHOhZxgS
2HAbPvnY/HdGZMWSUrBDQkSRORamjmpOlx3usUCOmRB8+3UxNWuuqd7zbJ1z2iQs3u4hl14hoW+9
fqqRA+6hHkgYtIbk3c+ISL+jgt6/4Dsod4hXLwzrDFXOWLAcUpckDjWTqVaID2GALq6vjtXMZwKq
ORSh/FLQqE4KcR4D5WU+PkY0Uo1BK8IhCJ21lCfyxwwFJy9Pn8KcpiFq4k9CqMWdFfzvpFCqbjPM
e+Zll1ArzW8AMWz1fekxkdytIBa9/MOBr0WKBL13XJWTXiibHDkCgvxrd6Safy6VIATL8VDvQc9k
B3F8VZazlkqH+CWKq8gN7IvYIFEEMp1G7tOjArfeYxKp9saxh9qPrpOvp2KeF8uv2sl2s8dvZXuD
Prjias5GsEGDETAXCtQ8SKQRlYQMUgGuFrRyZ18iTtOeQtrXl1V9hdE/6BL86Hzr+VTsd/COvrpw
wpuy0cE6dJJTi8kgAhdCKTxsHZS7R8jelmTt2n5NaqCSzs6FOs15qKMH8E0oCv+dZf9kOThP683o
PDmC22vtl557dR2XHfH6/ICvZyusd+bRI+YrBInym2RamX7rytAvT9e1S8ZknbnOQsBdlbF7YakN
gPLp3sP6+/ZJNBw2X7vdfewm3Fdzf4En24ny5HRKXtp1sNEzNElFJW9VRnHVncxo150l6ofXxFW1
wXzmKY+/ICwlcBPEKEaGRDc5YlBC0p9SUUtQkCJ+bQzrT3tLs2qdHd8G65tFvmvQqLFOBWg+BaNx
g0xCAkGWojFd69pq0MhCckXdhBiMpu2KvwDJ7yOESTpDH8I0FyCiKUIt/1ODTdwKCap7Kr0x2lWV
g0+0y8t40JVmog57n4tef4YA03veGVoUivVz1sJJR1Ll9EC1e2qm6JeYY2MW8o4rBv8DWByCBzTB
75S2wUj5TlhbXEN1zCpGv1iAWXvAJBRIyWkU2lai7wDf4XCQLD2uifI+XymGV4S7ZKo+W8rxc4Br
YLauzDmNmQwt+4ifGsj83Ed8I7mvueDpRa/V7X8fM0ZqmULEKDbKKH86q18UWNLqz6Ss4XHJ2TiJ
ah7qlEK3QWLTMlnSxPuu3OTX5PhPK+awub/mhLxeZlhdesyXjLWi85d8XiyDELNXD164JO8jLX0+
TvrlsnYcevsA/kqFOlEkUdFWtgIaw+1+3jZeJDS/rF0j1Hbmrkm81RGwne6Z/Ucd1geW64Ket8zh
Kez7SZxxiL1wQmbB/TeEExHxNuTzHbEXIWann6bzs0/kozJbcWnp7zh4U7LNRtAD++ANNsu67uUB
X9KzWpvziZWWvw7dDhFlO6nkwHITahAN/r2qe7UkAHSmYdd0dc2coQwaJ3lnDVWiAIf5gHJMBSTA
FoCPn61ecsz93ZSnywU3SJXuXd+CIPX95V/+4PlCZAVl05gyxMGUydnOow1QTgvAWwJArmlbIMfY
AIfWXcLzj799g73T4NKL0EzTCc0VeWJ3Zune5y/qvU/+AXaDdWKOB6U49P7FNc1HcVOBfvKA5tX5
r2iUN9QFXABBLyIRFqT8LREKTp9IUZRaZI6h3cTy7a+m9KmpvkH9jG20tLOkS+2AupKSNG7IqaV4
y2peLyLMdb1cuRop90nWMKCZsymb3xt7uEOV3XOJhcbp3ShsOIYqqLwmIkn11wtN54sbLv4g9wJk
2+UuHORBh0IJoodB3Nj+uRzVZBxQV6rxtoZ1GnjILXXV0qfmwV+Y8WN0UWxDqHSSnRNvRRKv8ps5
OivwgM0+VUbzWYkVNrrT+irveFAlAOwsq4Z+6tKm2LEmsFf2Em1EOlcnmevc2jO4+0FfFW8mrljf
0C44QXslubgNpeOMvZyJ7bz2NcPm9Pgf/eAZP1IhftBafj1AUuMEQ9V1LnH7z2cLArG3OwB5QR1p
kz+NAwFo6Ftl8oLK2XBL4jMSQtwZfwCVe1Ym2+5OXeXfsCm5YfKx1c9yeXL/COQwoKv72hDjQA71
41SHfRoNG5Ck0MPT8+GNwUwIcaDAVn6kI96MbKJzcXQvgKoLty5TEJASftQiOLx3CYS7ezdMUfHy
5ffhCHFwlwq6WQKS+gXgY4S28nQWTzFHR+fbwjAoQGFc5P5PmQNPxkxQHxZBHDyhENovcYXlfPjY
bW2AlUGQ01r9BnRPcys+aQ1vx4n1zQpRxDSHnCh+u7gQ089ct92VRszxbPtcPbp4lyC1V4Mc2z1v
clR3P8idaxeK9WlVrut2nMMkMAjlZnm3z0ts8PiCyhD0J53GN7zG/1lSqHUVK22nfxDir4Pkf9iX
kGUhYbjB3//MxB7ihqcnTkN6fTcIi9ldFVe7kO732HRoktl4aHtOo1TQ3roebYdd0Sf/yBWI1myX
xWqI1K1eYvQhX7UxC6PKX29RKojB22RWv7dvP4YO7J74+wA7mHJ4KScM1eEE3oKz9GjlHOt+sf/8
LPPStRqaBJmd0koexyLNAM8Zush0xhREMDhow3dJJMUg7a/3pQzUb1hlYrhFjd8q0JsTMtf10YYL
2mHunqU/YZoBR4IOrwUfeYhjhELhXokAcjrWCpCSVWpdzCC+8LpVE+Z3GAet0Lltlg5wMwd9umX9
FLCwWWmzo6uz1j34JBOP6Mv1HhT8Btgq01rBcEWKAviQHCww1Qy1U/QK2BjEZwA6oHjkCtXp488J
xCUqty+poyNjtXSxxY7sW917Al+/NdmzXI6+5NFTiKcT67FNDAUEf3OYivlqKLkJ7RNeUUHqc/d/
onimcpddgRL/0BG0K9pmqCZ9peVTtZ/1zqGXuzuIZhC2pWHSeM32cTUu0yv6udlTMUIvmmh+abZg
QtjqcxImXjARyB5PzlJ8tk6pZAraReSfzukYi0eR8SKgZTJ8SPAB2bQR0PHltyBL6dsk3Ar7JlzI
AMVjnQf2+JCqFMjEQv7f24oWlqzyil33CLTz3eoRhF6c58MrdzQXTd3YBA9DIW+CFBn2ZYWdS8Na
7z8OXVplJi1lsBGQ7+4aZRUawgd2TrpniuM7KT1i+w2mnSddEKBKyXZO7NBKwDwhKp8UeuzvFhel
32QiTxYtqmyx8fcns0Klgh83U9Vvu6ueFgIwd9WK+GU8wee6sa2JYkzQ3a5wkLIqubOLena/+sSo
Kt3e6QhQPJ97eY6TYJFSnpfLSbpSE+d9EtJWwv7Gt8VW/E+95a15Z7w7vulGJjKrSj7vUWh//7wA
scPCqptO+Lu5F14xQLplaSjMQBjsWRkmRPU6VohgeFblC8gcwnJiA4wh4GJyYTrN1cJKOdBfe1gY
vTP9JUXogFwqbLWbO3WWJc0IzlEQzOtxVZYCEGIZPt+gXW/dP+npQdUV81Ryo2khw7xWuy9ydUM3
3oSiVjDYMWmf1RWmUfHlSf0VrzXZO4rcUcKPisHLzrvD8bGbZ174mJABIyRI761MVcuUntv3eTi5
jU2IzYnqP3vwagjtQzIN/4IitPue2Yb1teUmcushr2CRQz+GJJgS4/WqZDF5/1e2bUWT2S7Aysfi
vxNQPIaJjPyjLsGbjycKttmMTDUTbWLepDA54D2O4FGckUNGo+K7YezSNzICy/n3tULOVRjz52Me
MuVCN+7E7tCilCbDdtbKnrJTPG61GtCVUROmmjJuGaCXvTep7XMoSdc8JnZVmfPyXxGFn7xzs6XB
OLS4GXgVUkrkUPJharTHaU+s1iNWfHPfFxCE4QvNKyVupgvZ/AUYabQOm5pGqfywA+83lyQxYFdp
sptz5KbQq2IQiotD6oQDL3ogElfmxjRm+IA3HTOFz5B4k0TVAdUklleVxbnvOP4SNtYy3nL9cMmN
BXwCfV93Yo7Y77CRme6182zcAPp5aP1oRXK6/Om/FFCsFYvQz+SD5JVf5hdkRVUX/qJdWTrFKuiB
KeeLPoA9Z1djAA7rZjSoOZX3RGSXOfvwZnK4WJ//wLSRRG653r+a4S/bXItz+qRYY4AeBfVoJ7xZ
PDVgDaqnSW/y2Q/6+jQ3MhK77r7Dioe7iSVWocd1YcXduSNfs2FMRrckfIiaoxP5ikhIXfsY56jj
cEuqkgGHMWpnDcJaJe2EsIXSnjbpEsu93CMpcUwXluDc2i3XnEHYI+0aStce/aUj/T9S7fS7U/pJ
9OI2f7poyP1BU02PsDg194qxCpL9r64lJOmYW1d+WzraedeUeS0i/ZLTTZQE8Ml/b9EyID2w1Y5b
29v08t1UPessZ851+6T2h/oKw1j0M5rjqa3m41llnA3g6ScVIYgriFjygSQ+xuuBC+DyVA65yque
qPIUR3gxCvtZE7N7KoTixEm87gsO314qWC5lZzOF5uBqb61dzTbyhx+/3p+BawgKW5trOoPbOL5A
hvtpBkoaYtSEFQTPGr5e4QF0unRbDpfxMJggsgeIPe8dhRu+weII8x6PhGy/tm8NR4TAIn4/NrzJ
1VIhJAdDaNywijvIVgDR4ZpvNqaGgG5RzIv2kT9n4n9eZGRbYBRNn52UDUze7QEa4bToYkXAXlLv
rn0kTATPVfhf9v+xFBbc9uP9wgd1FtZSmkCwZF17HcCs9v0rsS+Ks7Yp3YrAuFxIsA0sTvM93kUE
qMJ+CVRl2B4luopzPCXXOnYh6gMX4vzs69Ej6j+4zlOhvzxYNfzZxpD+wijkWoD3tDaPnJHvNn1y
MWzgdrXLzdDKUkxq8mlxBUCKbY+ZVULo/LykXuwxDRh0QiugllBwngskQSlVyDHi/Df4s9w+12dg
km6kAxIQYY18dq/CDYX+jLbavVmokxwtKY36bTjkM4lxpOiWoux67K6texh11ni4E3An03GylC2K
DW0N3m6syRJSu8iGBNOpVhXjnfi01p7jFsKMT/wDy+pgg4aT4PGNF9GKFIGDrPc2hRw+Lxh7McIb
C2/7VFJxmZrzv92iuGgfHCz+wmNlHnCpooi47/kNGAC3mxrLiWF60bzG/e6hwgQDkJKhIJzkFW89
bawj9IEXiNCVGNIFbMkfiG5/QD5JAFZPVW+p3h/3MTM0vJ6S6Qc1V+Qk3FgFa+zcnr9STQPjrHdM
AZwjxLK709QFRqCnz/2fOqoJfzmW3vTZNCMT6i69zaeWs6sUzQ86AlkCm8ju9IY8HxjB+GaBsSXe
INvPTX4nhoXcVD6m260ERTah+NcA3W16KBfh3DfaMtaBfXP1U1a39IroH3O4dpLGAnAwNMzopjyF
lJWvUF4bcCrRaG1FH6IUOlbpM4i0pIV/XGld9EYySOxgrhYau4FMlwTYxI1VJgGf8reLCqtPvrLL
7y6DkS7gMNQGbxkrmUKkPvqHnZPVI7Ep8nSIbRJvSvwYyYiTI4nUf6xMD/PVi63ekHwtVadFyEvr
+RvM3npv7QkPi30LXzaQXaXQzS4QWXf01o0fFgbSP7JnXPF4P8sRix5rTSC2Dt1tGq6jJKamKck+
Nooxu6rILCAJoVX+xAmLkkp9stFBzAZZTVnPl+0lV1clj+zQHoLo+KI7u7epidpqe/Wkaa1QYY2h
NBnl/uFmR9eJaIueBO+xroxL40jIuc6E3/xITYue5CF9i66u7GgpCBafPWNNfryiaLIkCyJ3a9br
DwVUADxbuYRP0ExkYKYKq5OrgvDHUVoEXJM3t4KPE0ZavA6COKBz7irfZqgN25bHG7Lh19IrBHbU
1+5KbJbXM/iBzGRqkSYUhIJsM2UZPaxwmix3fz/4f22HL2Nqz1ub0Mk5LeccuyE/HqSh4zU3YQUg
2kANg6pZYpunV4rDb3hiGb6Cg7HQ4tFcvUIJ/vZmk6i1+UguotbHaK3Q1Kmi8XL0xDBot/2Nti5i
tgr2VqarGH/X1/BezPYFDk2D8nq07c5RXq8RX5gl+l4M5ReVqzP/OXdmDeLBymJZutrJjFSc4YZt
MPR0pg/2vaMB91bXxBuPOAzrbk8xA4LQc2+X8uJq6jpJ66/7CvTC1iNG0TB7zsdaM2PUJPHbknDt
JD2FrC1CQlGbkDzXQdwzEpwDFSP3ZXmY48o9iRtjKLMFEexutQfKrxclKGx4EKzyHUeHOrAWdgGM
5KTiiNxnjmzHfic9WV/JZ6LdmLTjVQ1YPOgCCaP36rtDBHkP02UZDF/zYoGFYf1kN59gTyYCVc3W
SgqFeZzqZy2ebnBVZfT+fW5oiB3vdoeuxqwBqXHiAtJEmVOqqdPHMhwioi80KVQZjLWQbMFzFBVG
l1q7esRuTRxemRhLC3ffhoer3VptzTIVLT8ZwTpmKWOHsVn+YcaYdAIuryd1PxRIxWVkxI3FZKVO
u2M88AA3JpXP0wkXjNpxfBTiaTupT4GlfBom/bcIDeFXTapy/6VzVJcJY57V/HSm6AoVcUoU+bMV
kUgRnMrEKC9rN6vhjOLcqbvixhy777NNXv3y/2FY58AKbIsoynTo25zkDabsihsE3Xt1ZJ2uyEjm
Yz6IeHyPnX6IRTfBVYZc5ail8MM54AwqwDsogsQ6aV/LHRxPurp3fgbFmONEK30pr8Rhle2ZITk8
CTCm1qzQLLncmPcuKmQyyOBA3vtAiHbj5cPi0dSGXwuvJZg65q+CdSb8xvVQfo8iVejfJkSrSBgF
Hr8XSIMsRswpzpFu/Lqpb8SU2hsVrOMKD8gkSFR5Aq8QxwM8SpNB2aFfULF63fhYBZFrXk+rzln2
PJpZ8uOeSzRjTgl3A2551nbbQg42bzyNAnlZGP1x0EYFKWSieOd4AsSJcF0FVYCTjBa3CzDvxEVk
wEcd3SPXQMDiqzokqqq6UC9WRnWTlG81TKlggbt5yvaHKxjphBPC8EENWBMEihVcoFTTGNWszl3H
HedLArMOvJ8OA9yBv3RkaOjXzjsislO5ak8RCuJjuBHW9rftVa2QGuVvQsxYmMNU8p9wNxLh89/W
jz/fWds+zSSdv5bq6QvW+IGcf9OBmUjiJZduwo+t43DeNYnu/D4zS3lpd0RCpHra9pYKpIPI4IB/
dJAal6VX9sMldrBMpodTmGKjt/2PkfhZRL3SagboPeV5FNGF4lWCelACgwcFxfnork2YmtRcnshG
3+/YE3XHhu26nMsmJptgzy4QRrqLqcV/1bt4CaiS0uWT55mv3YufScLYO+sBTeGgFB8e9vgobqCe
87noePmlka19iLuVSgHb9r/NKuBLVjjJc7mI+3WBzLwu8WjC/Q1eCUGAxdyGLRrWkaciRhHRM+kY
u/jC353WigcUrFMqLqoR1Vo0q8RvyB1BQZOsFd7V35gOWKzmNnIsveyjBrA8XB5tzKorcDwEu8Kk
kprvnwW9ejimv5yRkbxcc9yRclwu8W441K+kgeCW26+9hZNCpXgRhfznjqXE2XnFUvIUzrtNxUEz
yhH3PAbdbGkEEDrwBpkbSN531qmMVX1njIr6uWCRd3Jju+ICCNA/z7PkubRaEkBvyWFVUI5Rd9Zc
ehazJmnRisMeDVm7pNWN/CifuMY9kbb2Hx/0Tzpbt3R5c9Rfd96Pt0pBXZAVY4JyQakUMwWBdDzL
C6bBgdUHx7iQyj9mDVggQCqB/9QFQc5XpP2CRqtQw1JUpMht2PuQHWUQu3q0wS74rGm/Udcv7w1M
W+j5yChf2Q+qkpjSKVRxxvtJNp92B6un3tkuLF4dvVkOIVbTa+eDEKsLAP5jGiY0NGb5T4JwTFAU
ob62xFe34hcKLVE1TcZRQg7UqJfNjwYJmqeO+zfTY7IH2WcaKTQg36qv6zgW0dzED2wZHMqqHI+1
5Wgn+EZESyhJPHI6VaRfqE2ExFewmWNLDrMsR+F537kXydSofi0DU6z4rg7bBWCKiQaeynUGZhl4
rS19WcDJksn4z6+wBzO3lGGfvtcEEgMPzlyfb8MPp5OQ//oDJksuToYmY2sJQEvMtW0tV35Vcoqq
PPliABrqyZkh7EU6ZDs7ejedjEMwVZvPyQ+zmuf+ZwmOHsuOIC3TRV+cczLxjmPeZUEyoKaFgXkf
0ymrcV1H7p6N5g3B8x/98TCzZWztQqsabqARGZI14BPxEJ15DGj8641QoaQ/rZGmlQI798oBe10S
TM+6ddZ5E9gSbLOzGxb+OEK/E8/YEsCFarVwCGZHHe2W9IgLLF+VYo3kDPgliVCYph+n3VkLLZJI
d3zfR+RT1ghIMEcmPIOLnv5WMmb+opD75eu7dNwP3OuVPRvrxCe2+gix+UK1TdBMCRg8d2Ss6V37
sMfFcYLWFd7zAmAcCu6E7UVC3ajOJehqw18V+7V7Cl86+y6arlMztNwpcPo6y+irYCwo2jcHbEnG
QLZtqVAEyjdfHIih0AcI43LBYXL0u00hG+sM6TAioPqGtrTRUYMmUJZ9TbrLjvEfjhSNciW7/kM+
LDoforuTQg4estPW9ziRG7HfyaQgx2CyIwRN+rltfKUramAawcJX4mpj2pygegdBG5ICSaYzdPIj
qVNTn5x3vy8D691SgGCt1w+60gJfk7oZzLYQEnYqWg5jpFbVAt+e0eXqOzIKIeGuXS6aBcIyFmav
Y1kaXQl6xTb/dIGwQC22oc0gRO0wuZQFv0DIDyh2fnqCHG7CsB76dsF0Ewu1J/a5P6qBRUjJ3OoK
WOtnkE3GswRSWulrRmD4W9lPLFZvJqce7UJZj9a+xthAbIEfGASzX0EnhiVPckf1O5006YiXaCoC
e0ub1xYXxgjvgrHtfaCyuySYzUJkhQiuG0/T4iIXSZ1L/Apk/2vOoiQxqAl0wlJxxW3TUsRSD4qC
wqXSPdJ9kLSFOtcYFwm0OxW2/Ch/hYzFvVzJaN9C7cC3mr5FlM1lyYkRgWUqwGMFJ61keZRTlnqB
Ce4eanvCYYei7OsqjqaKaspJcgIUio/443MWZfP5YY+sfgZP/lIS23NDeeTA/avVjkQVK39AVtHS
PFE+/FyJOzpmUb5heI2PqPGhYyWHevkBaPo5A+v/8+fdu9JI6uy0dmT6wRhG+ODT+22Rqr5LSn4J
5XM4B33ZlGKZzVX4pLGMJA4HtDra4d3IVkACeCQ9nguASKaoLrVXWSyzRYsFJId59/hdYLrPvEyA
sr5QzUeFlirdM+oKRZgg5xazUYkynjX+4lD2mOxxYQS2Vu3SkWC4oSm40WCnilYIWaVfJuQhmv8H
5DxKvvLVDMTSTp2q/5vHFaX+SCn8iNdS2C4zH8xuE6qzOPdo2g54unX9rltROZj5bxLdVz2hYOX3
pLjQeRsl52Wh1msyQqzsSfeIDYyWLuP9GZxh5jBvN/CkaR9F1ECx7lEfIKEkl6dk76g7+aEZVWWk
kmntmQ149JBA7HtW4Kj/Mh3aycJy3dIn7F5dAyAqVOFCeDs5RSiN2ia0SoH0DwwnXIkWxGKGhp4/
YrskEklhdjXTm2Nz8CkWOkunvrlXz/7Zgh8sr/P/IKesMrSRjUT4wYCxiTteV3fgSvIb5TfGmPq5
LsWkr5Y6MQ4aSax4rMxdrGLprVkV2My7Y+de5o6IxWEL3cwGqEmiIInEJYfx97+w1NhqR5MWyrH9
JKerfH4PpipLWhLi9tCt2MKxiLCQRv+tYjet9Z8EUBrBY6jxcjbGj1r660cF8Xa7S1XRitJ5zPws
vrIBnWGtRu1vEWBMr3wPGb3M778j9jL5Iu2Ufq6e18MRyfG3D5iNkrJZPlyq45h+MYYlGBZtNIEq
8a70+OBlqq/Kgyxx16Rn2FYOrJk0rsT/2Wx1NYMkaS2GOH8H/CCZCq6c2bRp8sHwofIb7wkRfY/r
S6FlP3NENHQ/2NMk+q2zKZMzcjvo1ZVMtognO3IyXCxckxvHRAPkXwWWYLzXTZ+eyCIHsnCs5AQb
P9HGtaHVZQw3nGZNoAMLXqPBkXCXoFkLOcv3DUqvQSYsgPwqQ7xv5abGlP/rjhZ2VJvzdJiap9NZ
KRP5ltsoTIjLE1LViPxIbT6C0Aj/yK67VxQln21Kxl0IRJEzs7MbZDiE9HJwJVgVfSz7YLg1KfJb
vremZ3NrXLrzIwoh5H/BD3mZPPsZAnpExvqvV02hZnedLuXKxH8vnCMXM7T6gRsTYLRxVj+vSlB7
KYNmbUWkMjSy+9OMm2x2znKoCb+OqmjaHuiyUTnGuPgPwfeOwSJkvpukj/D0dwyvDliCBVDGNmo0
vfYlD34R4xkvSUiuq9lpO9opjiJ2Zn08aqLKhCEr+O/mPLhMoTA381iTEWD8e29faAGQoEiX2z59
X8O/CqUZ/09NBxdIrZBHMe8a9JMu7VvHpHQsskZA7RH2/m6DhZBDaydLGHvN2MzdZ1wiLAZgPGCt
KPIAZC0Hi28CZAzBQluR4yQMHtkKbBZh4/26uF841FogGjLKuk1+Raiu0MLgnrOdYj3IrmiCKSbR
oACj+XpS8SdtufNJrum2mcPQ9roShh6sgEaU9ncvFnFXR7SvkHhInKqy5lhSXo6KHuvU+Zv51FJy
W4FAjwgkx83S9IoyFUPQ+rx2gf2Str3K1oa/eNIbnrra362SYX05sqXT4a6hzifpAlsVxyOV3NvD
PDnqIu/s/lRaQiicOls5zJ656TFIbFjNa8JmFtGnuDzhvt8Am3J+4D4XxHl0++4k1kvPRL6IP1td
X0H7qYMWq5vW2O3swmr8JL8nMan7EXXiMz03wwqi498J96OO9IXUa8CqQfwRP98Nnufvri12FAaw
xT/HWPSHuxrUb253lI+c6zy0yN/QP4rkKtMl6oWREqGzHdb4KBudLJJGkp3NySlxI3ILUVWa5oOn
jSEvMS6Pqh7p9LZRDQQbeQPrKC0OQAYuDO3WKQK/Olt6P4iwnf74xDGlb0Dx5E/f1AOI9gxi2xHd
4Ab/O1yNiCuzJO4ghrYhW4E8rkwEJ6l5ALajV1vxPyQigGgfN2y6P5cNOhcdbGnDnp/bBZ99y7yi
fC8ztV8gQg6iv1udZtAKIsSkKxdMKhbAZjcT8kiiHI3VWcCFWehUOWfpMHyCsVQF7zI84SXB/FgU
UxCVEWPr4o4iz8c+8Dts6WwpF0h4BP9w1pRErQotzbShXSMXd7ruu6GH1yJbsUd5vR91UFivjLhi
H21wcO4f3Zn+hXqOh7loj8XKhOnh4NR2hXv55KkdVORMQWvFMy1HZbCPH150Jr1aM/rZley4vEWb
Wl3BR0hjolAZow55E58SaAqXFC+sCou8BEDl8RSo3af/Hvt2adGtVZwVozHLG8hPu13fk/4oaO7A
qdhtpvAMp/6I5qbJbAePplkMTp6bkwqmLbcPbvqyheUruptDLBFNZD3DLCEiNisNJ/gWuhk2Md3V
bCv93OS/WrewgKy1DCP1TQd51G8OWNKnkhejx7bfANc3xb0HBVqPUF4l9M7DLgzKpbxgJp0NaKCN
lOBS5Byk9yWgl/XqlVDx7dOZi0fw9mwueiyuSZIN3y4H5MfOBvnXPlhQl89s/3a31vjs9C6rixG0
Xr4IF7c1q21MKqya5w7pa4e3NktfPQ+AC58c6JEM6g1S0CdOdomtpBiHevVxKZorfeNLn1mzhBbZ
ERtvR4APLF25sFQHjChUiU8xx4mjpeM0UaelV5ZHKL45IDQKTaZU4Uu3r1EFYQwWrs/ZYVyiZHBI
wDDNEpPW/xCwDET0klRwl/AYZkVWmZfR/236s7omtV+jcFBmR29mqXEviX48M/7b2yM0Znfr9fSk
dwXQIR7dQeHGcJTKP4NOLa8iGGFL/Ie5h09qbICzSGstQaBW01Yi7XOAqxJleqMq4HBWQENPKuU+
L3euKbsEW1jUCJKA6emq43XGalsrlUu9rLS14F5Jfx5jGcEuc8uJgN/33zVLsXBzSo+1tLDEiBhS
FID8gZnnLdXjgKLYndqXhardBA6gDKtfyjqMxuBQXOCJw8VUwgu7sB+kj1D3BNqUTdhR2zLxmJMv
XHRT9UJ9HJqR3RRwhGONPTcBuQN4ApWOhYidXmDJmJzG/l8qQnNAlTf2UhXBZThsaUqY/ccx6GRH
FiJ9Iv+xjH1jOV2TCPByjLSzFJWBuh7XnSU8X0Cd8ByzvKM4eZWVik/9e9gbzAl4z36VuRJQmHNU
AbR1nAjXQBHrs/rxArZQuRmCd4T3xiTkWkKMfJ/G0BsyD5Wjho4n/V71tJiTbGA3qNUTWV7WZ3e/
Nn7Ccqw5/F/VEIvKtYdSPNpyqH/51kedVuPkYgiTDVcyLcjOecn9IIT1rK2Qlr33nYcREp0zedTE
9mzGUf9Rnbt6iwoYpRnNqehEyQ7VkvMngPLz5Vu4l3t/XIyaIfZa9jOypSwrmp5ETF5Y/kVQeIxR
1Ph8WX3EOpVewLssAHItIKARy28ZALpwStmM9hNVXF/jbpdk4cLBOllmXbHL85VauNL9llfTafkT
OXc7k6fylIhfNgWQ7fgG/m/bngs69t21V1umf2SGxdBkKrBLZk2ZUBoZM6MHudH7mkMSQ1naNZwh
/oNF5d46+SWPG0lKAXKoY0q+i88NHAAQNhVz/He2Px6awB3wZfku1GkKckUxzeP7ipS8FpW70DOa
/ABmd0UTPstH1kErLP+K1GDrxPPiAJUzNx9iLO9hfBEXV86xcUecrW+5LVwt3WSrQyD0V2jbma2i
/WN/LLCmT2VNFtzVywYfUJERhYMZTRhMgK+4FyNmlCKqjs010OYHAIq3GeI/NJ2BKSqmoMmgGCAn
jY7IDtacyeXSLtww/m3tlfhllshMjfZmo5w4niVCCB6adEhnvzUYMRWcSl3tGjzBqqTDVrGqJqMZ
qT92dsieawRZoeaeeIcjamKemodX5psdZu9C41WvTGzMkJvKp8f9ZD3LGHnhvzuqLrAQtrlJ2zkt
syF2DZ/ahmiZBW4W5i9L3CLxJhvmM2zcgensQ8PSroZbGlCvf7h0fqrt5IY920HILU6UXSmJKX8Q
xgUhoiDUj3qVzqLqa2qudc/tyWFwPTdPjP6s+ICMo+VWZt3l1QB+bX94lRI/1F8Ot9q7BPZroFjN
jO/tNG3dHj6l7BFjt32YQQfHoT8WJglALEYW2afcyj5xUNJX94UChJp9pHj9PwiB8s4gBkdSijYs
NjBkNpI52JlN3oAxg01uCbPXpxIWheFDeIRpAV1U6CrAQNegw3xLvNKA0taOApVznnZyBmNuXKax
/1dwF4/PYc+adF8oFbZkq6fBn5H8qVtqdprzJcmcNFZ9m3p3iML7aP8qNAO4OkDxnMX5njzG1ffV
xx3MUqFOoWcRYq6UZKDlStfhHk3mrVUWktP94S0VUfDjQ/ENNgZSiw8msnuJ4ZPfu6V1QGqJaLwg
ngKh1GCpBnQbHEeOzcsIqOs5WuBrR5ZL7eyicUDxLbXpfIIVeCWdbPxGm6ZQK0ZxIN8aNKWl411l
ei+WQ0I6k0bHpDs5S8T0FfH4tzI52GO454G3lVpK/EHECsiR+EajEApFy94cCpMZ3uVh7saUPzCC
dqXw1oi45vMx2X+3A6Xc8bxc+Zc7gW7/DevjTJ1EWQhRJqgH2CYmX9x1YpVMdK9R4FRhgECc2CX1
R2NGyqZFy49wUjKcwg205sjTdYaEk8C94Nt0cJIguQ/zsuour7DueIEy1nwgK0nxqX40WPVKuZd0
axDApbDtEmIqLxUcZnEc/yGvEx+7PiYB7zp9LgYhWm27fs6QK7aN70FOkeQ1mjNPbF4lBNE13A9g
I0bnXEen2uv8XJtCWFz5zI10VF8oBDXFccA7uWodPzGH7WzOwoMblccmA4vv+ujd9obT1Yip71fv
VeJvu8+betG4A2r52tccDy3q+eGAzl0XlHG811CsSZnUvW/V9HeVhz7FUd45cFfv/NiSai1G03TR
Gu77Tf7JaFlTAa8XBs+xJbOHWWbgUqQoPxq1V8z7V2jEJPiLzYhFbxsFy/3ioTANpwdrq/0WA7Hf
Kg+p774MTpQBcHBQ5phNuYee4Jlo2+p0rw92wCt3jCSEVoAfwm/mp7VMtFbBNbHcGzU9pgWDVjzo
4Yci7DHqyrW040WbZDynj5KBZuWQcWYb7zmCtUBB06GMUY+88kMCYJ5/OmSO4vO2Ncm9NqF722om
WSz20mpdpeOpl1dXQad3T7tt0j2BJ0mqtFV7rkNW8kJwSFqXVfE1B2KkBmFpDrhjhaZyvqLv5DjT
s6W6vcprx13H543bXCI2ICv7q4+XR0Gdtd4+Wk27S1hBTmUGXUDNkxIm9AyGiL9lKR9alj5o0ObV
WoEqVejIhp4SlTgyNN1WYFFch+1Z9FUT692sphj7ygVeK9ZbjVmaHbja7x09iMTzvr4kTWybueN2
eFhi7Nxt6/3R25j/cSNprTQ1dfyel/w8YfggUJLEI/0rUUcO+yyPYC2EKH28cWBmNG/bm6KhElnU
vBQ5Ll+GWs9/O9gmBSfDtSDSDg9eIKT+bOluK8CGJrD9xsHorP4ehIv6pii/UyrhxxR+FA/8QR6x
H0LwYe6U3U5X/u4XgOpbtcZM/RLv9eS+YzCoIlyRMalZOW3SGcsl8xxpb/ZAuVDcrowK7cm7qkfz
L877ARdHPc7oBcXC2DAC33Lvhd94hcpPW6zTPzDjUCQ/uNjl5eu/39inKZ2K9TRErCkK9B+yXPPH
hxKeUz+WkNwAkfM/yRN4va63IX+/Hp5np3zAvAas6sG/AUt6Jent61UgjxGeRj3/yawtya04fsx0
q53pkZBAJ1CO3APtNEM/uC4VWL24u6F573fnauJ7i3Tr/NQ5ija3vcU6+f86UfpH+iRu6FlF75+P
RhL2ZCxCOWrNUIefPfqg6mUCi1QZMNEsYF+gMxCWozksnQsZ8z9f1x7BKrtkG9DYzE7s8Q08YzBo
+mgdVZOH0SNO1+aKNzOqwJxyXFVtjT23tNbQU4DE8J7UgpKrrNQdUtyxyNw9/1VHgnYu2tPPoGkA
XHh2UXRGWbjSC3TK4bTg54K6IAbv1y8Fo23xqrGoOpeJbdKhhSi8bqyzGwMEEYyLSjjOu8koXn/a
7VcSsS4PMc8A6UnmK1hwEAt1Zl7ATEXLstOrS+cVUyr6vMLA6gh1YK/zL6tsUJpFtua5cvp8EXA+
1Zt4+8XitB1PKQW1R1PvKeXhk5I8Mj3RAQY1RMcvFjbL2vG1jzcKEViG2LH2pBAKhUDhp0AdS/Qp
QhFhxI53kQIwODvh0YQfXRoq8WRdbV2RNdntfbp5LWD3XMf0t1Hbx/tUVPvIy/g40PgyWOaWIDw8
hyxzbmczKwnmEqpRYwk/0hERPXZbH9AWcaIkpV0qGRgHMqfYeKB0DJRcG14BgIV7cIeRZBIvoVDf
yqc7/HBFjo+rNkYxoNBjCGWY+Ob2k6Qr7qbj/Rnpwakm29Y8NhCTbBTtWrehqHbeFVkwGfof3s7q
lhdAQYzkPMB05Kh9BgD698HU9sQ2CTWoNf46vLF8Oes8YwdnlqXqtO8HieLJNlUayg6t1eID3ATA
TjMWxsIyKfPYAP7WoqnmSkLurmAMOPtuG67/qtwfQ8wBlDnaMBQs6xq1qZ0cjk1UiSsmWm2f5SBI
ThTep5bl1Gw6gHUIAEZQnv421UwwQ6Ec7Bt058eLWJ9kNXAiPA2zZv+HIt/0Wo7Mog2ZzLK8lGAJ
Ze7LuRwrxYUo5nvPc0OUEOV3NxOFt2iOqgI+jiL3H/Fz2BFbdev3SUV51b8cg7MTCfIZjpXQJJrm
0Y1H9GNjW5G2Xj8jJ5hfUtAfTpOxq8dox2DTzDWdHbwRFeY7c9pMWRofl2SopcCSAL7RQetoFh9T
miRTmtUykhg1x5T10hTOqD6f2mHAHFEw2mNqNe5O6wFpXYrnp51ioMCEIT//Gf7jA6Ut+8OgKe81
0wYzCuXmxWtI9crAKUv+ZnNmaMLu5k6hPQ5rvQ321BTJrxYlRRpXEMkzplyyoW7lMzdWMNJG+Vi3
8JSMmBXawWXyQT1XKeUTBEwnUhIvsN+fHTbUWeClPkDyfshsIgFUcjQjCJOVrXAW7HddFM6m8IlI
xs4JWl6fiJKF9Ci246GxwxpcwlSh29HdR9sazfB7CB3KF8kvYf8aADy9yxfmU2DLp9U9pXSLlBvQ
Qzju+iw2i4bohLbsrlrMgogo7upqpSaGUEaaPAYKevwO1oNbjFy6bvEmZJ+jlJL7AetOqjyioWpC
UFrXXe5ApTnWNPJbuP0/HWD+PI88bwRprWJdc8BjSfalInQkLNiHZEjUmS3twHHu02lFZ3q4BRON
bd2l5+gbWplz5LdTLru5PMqa10UO8V976zZY3qoRk+SvtCELzcqmCpz2Q58/KuG5LCnLXCBDn+wx
KxcogzpmvGoBGs5v0x75zir/NYLr9He4nJFPdhcE6kk8G6I/Jxy99QI7mIyq91YXwSLi8fEeb8f5
jaCGF6+6v1PAT/AdXCMX2IzPkP/lhi66446NeNvfNPY+0jdfzOugDQWSjEM6b64PkqECKLRTC6xC
zAw4f3phJR5VDy/VUefZZkED8zYmf6+J3RouUffscj4nvY59fu7Xgg4jc9jniFzZtcezgmDDktJJ
RuPmKd5H+PzFMbAck3UKMgyTUaIkUoeuQhEW3TC6UISxrintblDGdL+rOjA6UiADoTXt5WKgHQLM
+zOA3UO+Q9kmfeN48HFDbP2lxloLafQP34FwAnPlWcJf1kNDXwRBkaBVF2+0mjG1K/Tmffgu/Y9E
3jkPNOTTpCO1bMFGwuDwzEvfE3zOYi2/a4WLAoMeFXQu+9FfqCxmEUzjOPluex8Ckaa2ifp0PJHd
2SF7inkQv6z5iNIu3AswGq7BfGf0iQLF4JlQgxYHutV9gAfMjigK+5Xc9eVlBiXk0jTe94tZ8lBX
WMu0jMDScgzgvNtDZGSdsndTaHwi3LBIFwQarI2vzTHhYAA3JCStz7wPftffROhtnq+NzDcvE7Px
LFqBDKgi5FPn4ruxR6ywghA6WiLITVYy6cAGM05s437BLGRuZ4uu/ibg1uPz/tSaKTbxj5ob8tRw
CiTt7c7ghfkwmjhrmGdPUFD4sHkfxAgGaZ00GslXkq2sfSp/G8oxQUWUTDUuFtMVKX9zuWLCdaz7
Qfr+a3ZhAkwxQppF7JGZ+rsjvxo5xzpT8HA740BIiPMMCfZILYUqEsb8GKjaKT8jUa9jso/QsYle
sgRuu6/e2CevNDvN6gtRoWDwRWgpVEDyEh+j21c80/ZEPmkCmhwZrC1hRQ/uWBtrKsQ92pm/pPcu
87hyA2dhaw+S8GgxFP8Hh/LVlJYxTbY68/f240lOHMc/RAZIXh3rxC/ReFBKgxl+BMurWjDAgx1v
OjaDdx/PUQblEMUOCBUESv0MuvQOzo4GClRJFiKZkxwO8T1GluGi7RZH22KLzKfvvxc3kZpknTJT
scTVcX23ISl5Rwv+OdpGmPjLRyhhQRLF/gh8uTFcHIGT022et+KC6Uiw+9lrCHTwuW47O7cFX74U
VnmGLk8kA9trREJq9TTylc2Sgos+nzKHrpgMuAefLNg+JiHZ14NzXFEFH03lWJYt+v48KVPC6V7G
gFdsRV8uMCxasvy94V4NSu0xmvJmr33lb+iMyUzvZj9YulaIJlINvXzGnxs5PsJX/9H0uU3Ndpam
kr6b5WpupfoO/fwxCG+e5STr97AfqlEhuf8DtDxNdvQcpfdrX1jp+5XpwEzGj3tHHMBj79FyY+DL
rJfq19wKaM/j+12ypzW85xt3z+b34Kd/t58uhiQ+9CqvL3clHGhFpaMDDsrtdWJw8Y/+JWAQhKd4
WlkLRt4ERiI8sPGcA3SEl5pkDHQAkMBZndmOaE2HHKtllc482Zw66URo8lQaMjED69yA5GRU8zGD
LjHo+rXQU3qxZTe9oY0VvcCHd5048PNaHScF5a8ByU0hsoSsEIter6LXl7zXtqaTRQoRwuQK7kYx
1qpndTmHcgpakMYQXImqbxhT5zVhvtbJte0Fg+yQ/SqtFwP/Jz946OmG0CbbQbjPCtFSE1CWJdoT
+AMpwfpqKvoftOhoiLx5EK2ZGRihd8obEsjLbyInzCLRebC0DKFXPFGzl+c03Z6g5OUyTp6w2VS4
5Fo9FKbQKGJpnxdKbAySaPvkzUmXQpwbbmUAqkje6GlPA04AbGqPDf/JFQxPhkxMIrFb9GdFklWw
IjBLZWft0I5Ov9zelYtgMMwK0rMd9ccrZHy5oE4C6DIpU0gfsuom2X8NQC6J82lN06zl4E/Ee9O/
W02AroHHfGdSmPqvaVjrVnSzwR6UMEk+newvmS46A0Q28AOMdvLBn/UbDgAwAmKllygfhtb7JYSX
ASwNrL7mdqnG8ca7caelO/SiG3NX2XSlxrtxXuM94OzlqSCmQCcNP7fJHb2hvjXpJfhfiNZLrj+H
QOXT/3vek6iV2jLy0IujFYF9iSMLxQXcu6Ug1KaSo3MkG7elgMlmC6qADybYTzi7rP/92nv+SSR7
MbbmYJVzq0YnP3Bvuilgi1VFggBod6mXHqciNp3VgLH8pxRdfjdVtG+up7N5LgTMiIUJXVD5IJjf
FVErHrBDpSmo80GSKPGcrtQZQcwyn+ROo3zSiDWzPDQ1Jt1SshARTneH1V6U/N0+qN0r1A8WrDV2
p0Ah4A1cuOdY1mxtVFdsXF1xU02pBKZ1XHdqp/gavEa6XltI2hE2iMO1Vg/wdDkhbIF53RB7lQeK
Rhg0Bi1RzXcBk/C5TYZ8rcL6o2+Gkh7NVtL9y+BO5vT5jZVgoQgxpcnfDCYf6AeQrifvUi4TieZ6
xAJp1tEzqSuvgvL8G2n7vB/OIA/GpttJu8Nl/MsZkeKy8SswFxtF8lpwlyMx3C686BHDPnoaKDCk
GiiIH/BIDj5sfe8czK6eLkHhli7tmRKhMJueR4pPJ7a4MfdkQ6U8mWvXKJFKoIMkdAafeN2++0kA
FxJSoUtQY55p8I3ztug1c9nbp+9bF9l5J+eTMhGkjVk8eeUgnQOMrkywJLmDdBhG6h+/ux0rKoYd
PU/FxdYrD/08m7GAF+lFSVJx1BU3E2pBqwXRfsAGT64F6jZIXjtmObUYo3a59nYxN5BOqLWnJTDC
mn3WlQpz0+alS2t8zjC7H7wUruOaLyGc/B/l2xyVNrY+5resNKOlJE+lhjKOtv298hoeNkjGj4+h
o0/m3CHrE5JZGbD3g28LsTsa3b6egw6cQehhVnBXv23sgJ7ZrWbcepMTujSrNQQGxalSg4cnxa2l
HFYRy318SOv6fS+cxfzXUI1LADjHCesVl9xK/nzonkuuVGBVcnWwh78E3cZDkYSU3+urSEbB+rth
oxOzzXrIi4wxRZAok1R43yuc52K6IRibVCE9Y5Hf2FpI8S6BNc++hjM3e9+A6ou8g6LOudITvTvJ
ZdYtFS+ihkOGQAlCXeL3Na7HD9oJ4X/SnyPFtLvpU5VyFPVsAexoVr2Xmh6B6R2os2OwjM4EkueW
5bV2xxd9nFHz5peb3qMwt74yfRlCHa2hL7P7XPuURIP81M876idAL1XT6PCdfKdoiyM+kCkuct/S
QlUv3uvFN4JmcV6TxcsvcDcdJW5SdYEflDwm8WViaOw4SkQD9cIIE+Mfktg24pI67vwzsFnotGXD
zxxYju7sJqBMqPJVG6tqRWwQ2DOFzIkZH1m3+yvQcNgzkLpQtk0kX0GoXhyF1aZKt1yo7qNZmLuk
TlUPcjkgmCXKsNN0/gcs3YULqLmvDyODmBizPzF90hjBFOjB+CQ/49ueLaCpp+pV/1gtYI/pk4q+
ExOuv2JKdH6HtamdJsGN+JCAwziUccB3jsUfAkiz95rzYXeCIURpy15cLhZyuQqi1Yh09W9fufVT
UGAGXAWxT+c8sam8FcRxR0dX5kee3Y0SSAHMO70EnQbU4baXC+rTSr0/neoBc7AaA2AwfBfB7+YY
2JYfqF4qEurzI7+yY8cTi7y0fQ1SPg77/bmlzgh6x2+PZyaDduMAKna17TjMShOGsmOtOolymm33
bcD7Pm366f1voMlM3kudgCxuBA3sxGDR2+vYSgA9N0F0pvLYSekD5WIJ0cPWN2QeGDl/9Y7oMZmu
XNhfkzFsb8HLg0l2HPlNnZugo+bnilbGLTEUIBYnVaCRo4Dd9CWu36pyM6DP68duxBZaAXHnP8hO
Z/99AoT3Jdtod6SLjHyLb4bR67bt4JhQNLnFqu/guzLdcNymcGbhMM4QdFq5sU1EsCcvfHvMNkvc
kKjENws8vTEaS0b5C/dEzTgeOWeMKQXuFgm9JQCD0DSPhX9VaCxWxcnqDS2xuFtv7Jk5i0RvfF/n
2nA/1anQHUMQXQdVkq0nkDXFlt/TrL+Qb5aLBTZNzjuA5RmEaSevVIk0jXLvzEMToG3BHjgP/0zm
YrnFiI61wnSryeBVHzDXCYLiUV7BDihJfbMZ/BSvjWlb+e6oKv4hF0Be2gfR1V+CTHXxroaQ+OOa
0DRXApW0qBJz5fYVv69RpZDjnsyV/6XC3YzX7GaoT5CEo6t09dM++EX9m4IsG6/k7pAAtsYCf0eJ
HgKTybAx4rgCwbbgmiirWbJPM7gfFbKIdcoNDcAmt2DN+3XtiAAKgQ4nysQb/tQOQxnkG6x/ZFur
eCgtXkzksT/XxoOuGAPJRj48NKDLacqbmbP5S/8rEWp6GzAfA+PlXrltTH9IGoXCnmrueHdGRdgt
4BOvHmBQDzcTTSqUzsFgUN/GFoeAGNWD4lJGVdQDfc9gewz8REfqDt8nt5+Z7z8y7Il5QNsBTEt0
iXzSFNyfuv8zukVtAaZfcXEkcuAWCbHMlKWPWipdTB77pGwNMuAluZNSswXsj3CGsIh76jw9bcGn
z1iN6zAfEYFt53bRbWDlRbcf3WoncsUpIdmVsQO4L1QE3kFBGfUlX97lTrhY8EXJcbRhdZbVM7jH
kcUC0YF7iEubgS+dYqZYD/1QA4nM+pCzGT/JxGvz2AqbRpYa51k/oo1LXhRsVxSzEAJNk2joFlf3
+byHv+5KW79UR4g+cMSWCNu6VluHy+xLgMI0P6iNzcDzoZ72auCbqvBJwGBblukUS0tNVhWMyM/0
ahdAs5j8cHILH2aQ0ByaM+wvsQMg7iWyT4MsxYtQ8Zyyo2xYdKt7GuvMDvh+ZQps/D4WZYUXmC6v
p20lN5vhdOZyhKrMx2QxREJqOSlTJQe5tRxZbW/jZDE83TjLVrXvkZ/KDkn2+vbRZELcHp2gwhIE
1De/JcZ4VDOCmkTydIbUpONXheEkVszANbGv5zCSFRCdPe5POAiwJl6hxNE4gIN7Wq4dmNyhENHh
zcSzivc1uqI83xhQB1Hi41bXAyszNMFCFDiAqpkqFr0WMX6rtlDa+inwitBs2XadG6WZODkOUlO+
pNjQXU0ShMOz8i8AtvlKScJjmdcgT1SeR8w2ju0c+b2wTFAlDCzxqsPFZ2ZVXKIF2Gc9IUI2avNq
WLythMCdVYb3/WJnMeMgipDCiLRBus/kEORSCkZEIzqAc3hQ/2C9rcfOIhGdbDlrOqQNqSv908nx
fxC0NLEAotWEMgAxuQ77Z8T9yM42uxgNGJ6lvGddlvL1VozpmukpK557fpZMyVvLP/cm7wuZZhxH
RfIMOV6nJAnCkIMRG3mBzhWiJplSPBUuAYxxsPo486oedS/ba0PoieckoB+uO+HxHw+EvSdUkIsF
RI955pqa57fthR3w3qCS8Bpyn55aE9UCON1MJOje1YvdL33UJrq6EZC7aWHQxyupJyeDEGfSEMuW
uy4C07B2a1p2sxNW2RU5e/5gvKsuIsa+366vGZu1Zmscqfoi0ES5ysJmwgixFuBbVTP0HOmxJGd9
d+W1Ep0bvdQIWELvPfPz5r6jsEsTWxfjoezbO1xvxAc8PpmdwsakqeMGhz9YAQa9XOVJ+4bfAgNB
nTBA7OwhD67GqOKFSZNecO5o2gIkAd3d2bZ7RsUt52xuqL2w6/iBcoAMtSPHxk2JleMYS2/8VBLL
2Hw38eRKhjNsjcRQ4RsSuBxamNTCX0UtXVVkmQzpUzuqfCGdipPJricE3zd2FWH4Hwanu9UcCgpR
C2efgmcW4ug969yW1yJ4g2I0orckwRsPZpZ/VHZRd4jtkDl3BRL0d6DzsQmXKGiQ9zUrLD4C+y2Q
1fgAGw+VS1Z0QsVstGD/w1nstIPFqJ0bGB0mjnrMhXYz2yJMNjyvy2xQJDn4rf0dHZZR3Yi+6U2X
mABjK0DE342hxwY5tfQdyXZFMdV0JLvcUw3TmY2+xknwYHm8eflVY6vXRt/L+aCuFx+GjN7VHfw9
gZJF/3l6PR5/VJE3tIcUCc/lzr9zQjGLOQ/MTMv1gnuNiUS0xZwzlvcr/gs//nmhEzGljUz+RvpV
FZs/1JEx/fF4UCwrZ7PDUgqYxVHM1U1QvOATdbK6HHYc1+uqDCskuMxqWD6SBi56dTqZH0jZ7V3/
U71Zpoiva+RYNOZyD/0clUmtGc8Eh0zGgSNazfhtn4RpsllpRW+o18PrxOlcRhQ3xSYjmP8CXfif
zjwU9ILwHqu9lBuLAc1mwzaC+Qq/2mhrPZmONjWdMLQxthTxuvN3vVpKzIB9goaTDBwqVk0+1KNU
CrqWGIas8fIdhsjYWD6KWHIutu7EJIIg9H76AvlL1yDJHoaRaLvm5AzBL5hUzegLH57EXmzRY0BC
B785We1bmymKFRPw/X40i4VXhE1CdW6Xqnick9AMx9IO4oc86D7xXd9Ahaxrvp6R0VaZKzYxG0tK
DV2oVBkw7P3L+Cyzen/EfAcFKGVtIHJmxzLYZwLzUiomIEyd5Vl28Y6RiszASD2C4yz6uJ7tDbMA
CJj1peM7zFmo6oXGtsUlBm928F1nv4px8iVeesBEEEQmSd0deTkfJKSACDP5STloxbvsqO205MpE
ZX4ufMbdIN4ricFVmSMMTrc99TUpNB/6XZ5L2xqjo9BE/sLSiwCnn9YOTQXejd8P3IU77W20h6gD
Idunn1WKYw3sCQ+dze7HimsoJMZzIOT6EXf4j/yW4afnprw0GhxtYgfP7ekdw+yMM07xcgPsVwZU
LIz7/zTY/IRmLNhkA3glLEQXg2m2oEuPOz69UF69l7Ly0fLu4O0BhPC3TsSCGVqdEurDRTRMWiM3
0TlrQWF9B3adqPHfMfxsbIrmMYbc/J5luqsuwMsjgmYEbBdrw8wwXzqwDPru8bv7JxDBSZSHx9E+
bbWQ8MY3vg1bwzp1oM//jStbO+csCw8AmNaU2o66A9T981D+x8je+u/BmosJuU9UnyGfv0h63KJL
4DHwQxlKtewBOvxqzXlbbiF0ObgXAKrj/D4jpQYqTRJXO/0ebNW+vSkPOI7wDRuRA5rS4UiskWiu
C+ae1DJtbSuIC3qVfNEsvHfWjvhw/KZZUorlHfDsJcQgQvXcivUaW1wk6JCuxcX780zEQAnIQmuu
aHWTO6ABfePAh63h70B/WIXNvNwMlHvKpGnZkQo9hkZ2Ess7ZqBqzN3/K/Z0gnQNgdhotSaMjHC7
VakSzE3w1njYH/a1ahlTl+qeHITP9su0YiRjeu05538ZUrz+yvtPLnbS/OTs0R1WfJoSZEblgf+L
zCnvQ4lP7rl8w4sKPP78W3VJmnx52HAbnWGruAo7rqIBXdW0OM6COuipc/fgGOy+bdjhdbTs+4H6
5sJhCML66Iwdgr5ei38HBQTp9mVwh2Iw2jPjYoj9AHf/KtQv5MTb3CvNcFFEw9/5zKehLYAKNCsL
KQo56yEkmPwulIbwEiJv+smQuOmkphEqPagNB+TvaS2Tx4N5w2ClR1F7WLn5H6syXq3fow/Md09b
NqsSTD783s+mJTkYymuoJbx5FbAU+8yZzIpdk1IOi4HSjwTx7vw3gQ/WM8KV4fj/6hHj2NHhMKG8
LT/Wn9E+56Zgq8bBn8UK0wpS/4skXDxHOJh3Slvmmksd7O0RJPr4rrhylFtvOXLYcbaCqRphpX4A
4ep/4vz4pzwjAb0hh+w0WaXupLXuu1NtK2JEbg10ABeMdfW9+K4BasCIP6D916igPC/0HnMtWnzP
1vo7sPnP7uEzhX8RqXd6Ksd0Ux4uULNvobW97YUQcNSQ1aewpZbwE7zVmbUTUVyKWVTh1BLjaP0g
I1rdyyEW/UhEaucASH5EvQbbItDthTTcDM23ci/6GmSSyhzPFD4uFEHiwdi+qqLzEMGYWnuzs68Q
pZpE8PmNr5jQXRJLnt/3hSywMl4ORwnf5idM3Lw7YGX8IB743g0HJc4G9z++bu1nRfIX9yd2FaRc
P8Vt2xnQmqE2ItiTucBinjo6L9mwA33PstP38oZgLtlKjqO78LwufnoYTI8aZShid1Mvgh8Iapeg
7QkLy5qUYzHbi70FXOyabIhOPCl6dlJ3nZDniXqKsRJPrP9AQueYiNXAvckeYR3fdDjNmhskAcPA
Hta1e0NvjsYOc4J+C5pnHaU3gUIFlgZcCKi/XFwJES7R5T5X/j6b4DMReABAiWW4nH7DA7R1W6bX
GA4J2JpnTCpXgETKamHkg7Sw/BQQ2Pbk8xUJrTXlFunU+RqVbfjJGgahsrlsthThxbaci0euXFGF
UHv1roPw9QrOoaGUXIMOnLXbAnCa9H9d5a8uWvbXIijLV4ZdrEwXzlpt8v71cGFLf1+cB2hejB8o
0iZq47oN5YfGTGNfBfx8J/kJc2otFBEmCpAUn3Zbd3FydLy3E+OcgDPJXdKp/4vXiVKo6GMQnXTH
I4wGRHgVRbmAOL96Z4lz+mgXW525+co5CO4D72v620HC4QRuSz/vxVU00izVB4/eO/j4nMVgguG1
QlpnpVedxIQk8UxwPQWZvzwub+NPN8pJ4eDuVLm2HDZ4AOjS3ZgZ0h8tc27GWzoYKjSHFJ4LvodX
BxTzqP93o4qD5NRm3rqwuVSStkfIco2MsrAXYhlqprdzmc4OV6dpLgvP4gt71QGQKeunbHxlWwlS
seCI7T76dP/kOZhvDb+Xfo8xP9S/gXXpW+zhSbbVCFSl43hLTXwuwMW66w1UQoq7j9SA+lZShnud
rLj4Q8a2OPj6ylOhtf+FfscgVbwu1xUqSTW8KTVVQ05ArISvhnfxrwy9yd/EvRB6wPTiVwJfdEjF
VrqPb5HR9wwHXOaer+mdAqm8TO7kXGyTtHSuZgkP86v6fKsqbQ/hlWC8nhfYVCbsnRl/rOSeIQqQ
UiLGt1hcbwk1HqTpaHzXFL5OohDwivElEXXFXF/IN4t9kLK4+pZAoEeo7CXwA0MV6XD4jiod4iEo
xgEq7o04dnmwkCrHx7Z1sqUe9UQepu0gXYiowfT3FvONlZqNpxqS6m0KJmx+TPR9mKtG4Q+eiKB5
NaeRaogzuy61arhpKY+Nd7HGe1wATRk/p6s7zVxlFpXcNJjHZyg/TndrM4dnNwsfmtiggECvp7xZ
wNIqWFkLD3SQO5RvMFJuHGGmt2vdyv/j3VzUlCZkSquRZhJ2/3wDpl/pGOEHVCafoKd8ao3wXhCJ
pRJmSab6lpY1ArOHSTNTMZPo1e5EZPrRXimfg8zFdQHW/yWQE4TyNxXU73X/Q8xpx4r6cUU78igy
dm0VXwfcmmdRW5IYi2Pcps5l8CFtzsXs1MlwkjlDAT6/Hpv5Ha/hB9m5+VAof5haVm2Xet08eDam
0k1DqwbMZ6B5iq+wfNZYgjf9zAu3F3rr7XFhZz6nkp1l1U2w3o/SaOZSjrVCGj1VRFCDzbnikAGU
o7Cm2E5xcZcgRqGnrupPVunkKvQPnJe5ESMBgvV2wQbb89RhrpelXCJKixE4DDE2JtD/Vfg6NvyY
FkjKYyK2oWUutfn6eoCD8bKxRGGbuktI6TCKFOFDJg8/Fj7q1tXgobFIlIe17Awf+ZpspvQNkBOH
kUdpueM1GA44YrXnVPGhAzW+CS//US4VMKZnOT1JyhH1e+QkGKFIZacyWGL++UUPGQAKBr+hKq4H
z7WXwEQvREWCWHjzVyMU3Jk7KFPoWwOBbo2N+rYiNkJj8i25WAL0MCOosKVofe5aAHQg12v7xELL
FLTiWdXH9ug+YaZITUDXfVDpCTIUqurcKJxYtsLj8lvd/hKQzNSXe/CmQ/muqWCVCiaABUdVlPqC
VSRJBx0tir8R4sWSIiksbdxKb1FB+EcHxUzHzxWogilB+JlzDE0a8UgHQ/qtB0fQdKta8EN4hzDN
bCyyU3RDutQcmxgMI43yMVDDJyTHdy80QZB/ZW+rfD4RJ0ROS9c8hXiaDdsDkI4zyuV4AdfR/Ert
Fpk5H9TdqZFRzI0E1+V8WCfpgxAR5AF1AYiR6LilsXgrXRcdbrwpm54vePvc0jDs5xiz1DRH0q4y
/TA0n9UxaEI3EubTZJkF/2lvaH5OjBirC0wbenjqeK0vb2zde3sYywnuRMWjZWl8APnbxokcaLem
EsmjNUT0hn5pm4oNmYiSgzE+A5yXAPpWBjpy4o7RR42dNITeVNEw2PPeEfOp3dw3XYFVgBfGfUHw
YHXXojN4SQOiHRxzzSh2dxwOzvoa+CzckMaVSpCzianEwMmk3WrsRTeyG5bNDFfT/LX2hidVicH/
q2bkk/EUUoSDfwd6y80jUvtgYSD9aybeP4BKKA/SVtaJQFH0tfU2lMxXSkv5btG67ae+RssIlFEH
eqPBTw/WdAra+nSK1ST87brfnUnX9c8YBRFvlFzGGNXRzsrDkEpkIIbV79AxY9gvaB2aMo57P5Ks
x0Z6PkUDys4fFRW16PkpvCH62AQcrrun0AzBFq7goTlCJcJOw0h/vqOkz6oIMMX8jWkRH7JISpt0
yRCl31kkBL0/WTT6Rnhra0Vooq91uyVA+Jigc7rBU+acPnPAzOX5TmodE4vW+wPy53cOipWtxhSP
pYbyiaAnRmVq3nEeSf3+DKo5CysTogSkiJbk2yjYx6+lVTCyLleNiCxYXkHmvezatfPf86DtkXO1
mYa/JuNEuh9+O2kPLuiHKpldQzrwGKT03pb8ZwYHWLapPIF1uZN/JBdUVc+o9IuJx3jiAlXUlL/k
BlgRJPYIGySL0xbP+yTWN01+AxWXqUV8fsXUljmEvHGhWgK14NtG3zooJtaz9BGxq0tuW26Ak6xM
EGzS43NXdgPE/bX0ewwZ9AbnYJ4prhL4/CNHg2aF52ZU0h++mlKjkpPWh/jY6FSllXesfDLeqGXB
T9ykogqgLQis9xxeT1i38c9T1cokc6OLnobuavDKwbFHCKyE/HBQk/2kPH0ej8/w+fwBHKpP1qiX
exJdhkcQDwbwC281LUO+sdu+/M584Npi4rZmjIsYmeaprL2LeS0hiDEMPBql0RB5l3L2UspcJcjd
czPhrUqaj3SrA5cevUMSLu+6ZZZOiVmb1Jyd6gg/AfkB425aZIkSjaTWk8IHQHRKwwO7KLcV6BqH
m4ZRxUpqORKnGyTC+9OIkBDrSSKtZ3XF9JzkW4nrkG82cFmnqmqFL0d7ccnB0tBtVxU/eKpRaag/
fTkpV2pC6/xTe8Q9IP4qShF/72HrftDhLnU2yvy5SLaVFRZL85vDu9HMK049aCt0Ygpzq5Gpx3gT
ElD00IgY5PlMn5eDWx058JGl6PPTgK0Y+l5JXqhwdRAgdJ1NVHhd6vvgLc9z2lxfiVkPDDlXhX2B
I6I7VV4f0v4DHMm3F9H4vRT/+Vs8REh2cl7fBB4iUPM1uRDRaU5GgofRbhOjLZOWD1l1euYgQVmx
JNyPpG28QUUbRoc5TGkxRe7H2C2vFoDKiICFkttiiZhleAFMN61IQTyKYitNXGHGH8rgFECnw/OV
6tjDP2NrfOw92tLqTdkOyujiUA1J20sJPKfSWywjQy7UY4fxPPH+L+8MwMdzZw4wgvk3WXpNVkOV
78166wstaG7huVaSSE+yDAhYSPGwNFF1KTAqe9qC6qQ/iCTixgE8LnXJGIGWmBvw6Hgz3TzBE26t
C200I1f+M8n1mV1k1E+3ZAZLuKvHBq5HqnGHIuvT6VpYhaBZebeojmOI3VGehjeb1psLx/jQd7cP
o7lmSLkdqkPVzs9lodwQg09drWGgSbCsSeN87Ieo4KCewEJcxsP1rp0uiHppGyvHwgfuWFELsyZs
g9YhLE2dTfAbiQFO77oVNySbxc7zR3gLqiFO7INt/t0wOp3WrkSyDHar9PxC2pE6LP5VkbmF1E0P
leiY3CBBxJ+Ua46E/6+tLz8uIHk8tRhP3dngoQqKDoY8b3iPwcYZA5tbLiIAi//irvf8XAy13aTf
eTxh3oucRRL3KN6YYlNeLKek+dRiuLGmDNV9jRlZEj4Xu2pqKJbbT/Nf6tj+CJGi3KvflSYCCfKA
gDkjKy5vbi2+kbrXc62P0b5Or0yREYk5Ie7ewyp+5OytTnFHJYf8YH8tiQnAopCEojkZxhEAoBoE
17dm7XSPBwlRAWot1J7nPGXkGSL31/7n543N1R6/wNFdDvwirKAMGhjs/T7w7202doRFeo5SIDSA
BBQ0itU2h2bqub+1f54i0tHSqeieQb3RFb9UD9Cz3UuoW3fVcJAjSxVzZS7SPCBVZP1+0PgjqblQ
NowWfe3Xk8km8k4NIaWZjytFXWwpcTC17wwP3qErXhCrKGMp9gBztNRN/XtsyS+BnzwCKZdZ+0WR
UDnDMz7nxcnhft53lMNf6nwMFwp579KmIdgMWANfzxWlQ8Mk1xPmrZDnx9ps2qFnj8733gBbZV63
4N7tn3tpiJu/L7oHpBxcyOmuzMhTcphe3FnoHJRqjEPKN5B6fbqZYRORqdOi15WYoXsuupoxOBOs
AsvVf0GdySAZqHOZIp6s2WR4ScDIcE3if2PvSBfeAx7b+Te4MpWqAJxRcqTPioRQkWC7e6lZqQt/
CfbMNWkbGgpTo9X3NZ7H8Q4q69TivZPf+ZXV8+RubsOm4XB7R9kEdiGK2JoH4mNug3SvpQvWk6pG
tpvb8+ifsA/GHkEgSS1NiNqCJ6VWnMNcKbR0JsOjc3p4x+PA+gK5IIiSuPCnxTAOGKQ5sNCc/7Aw
+G4p36THaWKNeDNlcun2daLKEC9FZk6wziFIiljAGP3eyyzQdi1bAvvbQX56JqbOU0RkVOwIzcT9
uVxQyVCsGQ8QMiKHkIhdgsrcfnJfPOLErp6eGGb953uJHUqszzcuCOpgcJ1e4n5qkaWpSBNVK7Gn
kAJ0vFhjY0q4cLxRa/GY2hlu+3ut8R5Yl89WXZX4vV5BohKjFbHVgBsBhonk5HNQ2jHSsVVnTrh6
Dm3DcaifVzsJELVUzqM4KLXR5gQX6t9wa7AK87EjSpakH3+BztIgHhRZ5ucP0WNDQUMUwOcO/Zjp
p5jBEVloJWzgK7cTnFaprvqctYNDs0IH9CQ1KAevAvKZe0HyyMfYc/lknCjYqqefXVgRu6ADHodZ
3vVcdXlRQSRPI4CnpKShDke7wQBgxtkxkIiDR+IcTSg/r8mLnhoGNy/SX7wycpIHpEVdUeecxcAK
Ezi/e7jWxYCx8vt9T+aCaVxPbFuTS2jGYcgp34wgWG2UYZjbjxz+Bjk0Df4WexNhjnhaQLG0J/Zs
EQXtHCnUHtzqxLVNq6e7BdAICSnAHofqERYqfCW9KZENsCphoHxpFLE2lm5XG3CHBFhBpP88UdIc
QU2+NE13+l6dT9RWLcFn3eA7TnbPjufFJdizp3zsPiMkvNFZnolQ2vuojKsgRWIFLcyx2RXgsA1+
OjbRQ8TMsNtNeTknp77GDotHBm4aLOkQrOn2vlcimvU9wqmbC34HqM/bHJJnRafQiuakGbSYD8wZ
M3SzfQih5qKdwpqtfKihPmo9EfWP1nC7W/NeGiPlCjUzuiGEfLAb6SbCVyt4BEcminb3w9kWh4yl
pmWIcyPYlABEHWFfJYo5eIL7+bzZfiCjpLJApqwU29bbEDYzRPL0K0wDnojYzb9z4VY5nWb7naMu
GCdZcOxjaoFOMcCXkkENJ9Lvy/4eHbRKKEIFNC0WFj6hv125bru+bnZoD8Eoy2VgWyfIfs/ghS7z
7J0xTJkX0VaMBNQ0H8RnNfnE+VYa6qxGQU0jAWi55BzB99O1KX8gXPBh4hQvJ0O45MIh1f7OQLsF
SiFBBipwHV34X8/RVr6zjh2gPFAkTZnm/5uKLmYS8JcTRTjxxExvioXFTCBzmpxkCq4lqpGdkr4s
wRyFVNuwypCBmZ3xno+TytB8/LkdzvxeWeHmDEHNxIuRb1GekKDidaq6vog3YHOqguhwzumM/ao9
EjIs5F1Edz+fs2GXDnk7t7r/Ve2iUNUqLH+ZqXZuGXJbk+Oi70xr/e7P8nFdOu3BfpsfOUoZFXBU
7AZdYAORhKGm73o5uj1ySpluBmBxtTYZJWTNOVFgiIE8GTxx3PrX5s0wtqHnUNnGKxSkSB3X8dRN
bbYajHCbGbdyTCbe+pgZSB/03vLEJvPrRWqljHKr6ZERWZfmogN4PWElfWi5NzuKvaT429nGEgvj
RxCbesEF8h5VEb5GPXHPF1Hu18oaj0z2kCDGG6cDlnYzDNnQY2MVKbNWYkTbXuFFpAsXtqCIWGlE
x6lTSgeiULw6K6yi0jpP8SiLlovORO74yVGyUcy0R+evOW2iHPOhwyO7gSeuzJnvXwMNumcD+Dsq
doWq1JPO0yCNw8495wy9Wgp0rZgn7BDvjdj6Mj6NEndKwvGPMOffKG/VA2zDGtJNbajSSrc+0bRQ
G1DiJxyqp42UPfwGlp0hokeRpyMmTCCo5JM8kiT8H13sRnEYF+hwV7kClruxOwHpEnFog71JqMNP
+cTYPfnzxKNh+oBOM9RUJcmB9DwWeeL3htasEqo4UU4fpAyinuv5+ruWZsHVcekk+v9XZiJZZhcS
ohScZ9KklkdKe6+IIAO/buc+GUBO2sj1kmXzxxdmi1dk3CcDJ7DEdlKzZMob6Mfz2Vh+hyGj+v2p
HlWGtogpc2gvEA531c7tEFA/UiXurC5xkElagDYO/7SPn+IBMLUwFymg+Xq/Lzr6tCwEF/De4mMk
7qSa/RT8OEMK/BdvWfPZyu4temq+nM94F9XuZ+mGKOjBWyCJe5pYhe8yOgbJL6ufBPPeubTS2lEn
FfI9jAvbk4xrwFkWKkknZOZ2IPae1orLWUrrP6boHbt1PSs72CazEcELvT/dwdmgeWBr9YwPKOXk
Ruz04BMzcnuw7NAJx+qnsjekupDsT6Hnw4HS6pqpHUCfDU/JYeUzYdmkqJh4FYiotkIJgdfFuQif
aUErfBY082QPPK+SsDWV+nbWN4vDNmpbbrw8Uv0CmtkmFSUDcJFamrlXiuWbTYq49XLkDayzo3Cq
NdDWCgWRE0G2pd+P5IN4ZLE80UxgECee8LAEehRNdBx2CAbkE5AT0sK/5iTH7e3Ql3g44zdlmw3n
IUMDNc47oX6rNA/943PqlgkoynrkyfRVowlfM+nQnhUkHqPfqxORauPFb9DBkyXO9MBAGZk5qr0Q
EpkCoeEEVZOhbCm8PHBS6GAUnvT6Oi8mm2Ld6DbDt8vC/cmIDhvwYFTLUUvEt5nK56d4w/wQKQaI
crscVaPx8PxV2O5BhZwU+tcJTBYtpmTVMbrrMyIajBL4WV1hxcKoEtYU1lOb1dyCUgGkcxzkqk6g
kiU4J1iC/wOINjrlHQz6+pUUsBjALP11/miJVAPOia0fmy0ct9iZqajypFMpTlReEnSLBNGU2Hww
GZfQZz2MOmfNLoitFDAZgSejjhy8nbqK01B3IjriQUFo10iFh3W/6/azijrL4N/onPqf91F5u9DI
b/W2E6HO8+gjeVghHpHOM/rXCu4pj03LhPfxyDEMRGg6c8KNQQCjkkfixj7IUwt5vI0AqPty5IKC
OfGCvUpfEcDIvh9tSYjUXaswYJJDzzyUF0HTds6bUgi7XTvT4y6Tx0dJ9Xc2EEs/YYX51/vivXHi
SN05B07JQH6XCWj6knKzPNaVfvK4sruIXnNoPYqlxm1YUgXbZLGoVaITvaHVQHsz2bwqVJgZa8NJ
W0xETuC2SDVEU9XEss1tG8/2WcwjjeL8V2jERONrYNSNoQ28bafie4wLmnrTEEiLo+eX6h7e4YzR
+V7qiSu9PrXhSRNUCv0v6sfpBoaw/Wsju7tSjNlZwRwZHzcGIvqwEZPkI0U9L0O9WxSOGWc7TSE8
uNH4HJDRs7+fxTmfsIr1MszDQflfC95SpnW4dSrF5XiQilItUyUrDenDVj8pflBuFqmXPNldAtP4
HoCzdV4sxhCCNU4I1farCKESC260qE3iKmxYiQ4fgKTx+GbpY0I1k1AQxxUSXYcFfU6EY9zsjIph
xRtpysJMKbwLaEnrr7v9FNQ6QPiIShhfy7fQsXM8uCI/BVj+tiWH+e3Clc5oajsDIuBohBCIir0Q
W6sJ4kv/t10svlQjPjEJOO5WDGSVKD09m/q6fGAQ6AGSe7oFUqBQkm+KgXNUBIAls/VOgH006xdh
CRblsY4uWAxedQbL/MkuhzHo2g9Ka7jLVWZrt3LEVGzwHFUPuF6sKXHdGQGbNLTFxud4ppzpTogM
xA65MYqEESag+x8Eg3gVtahwXcDnvFrwlGfUoJt8Hkh1p0bbJS8uoVIZqvfrc/Fng3Xk8hXC2WCa
U3zhZxwqucCWJVeuZ2d0vw4Gh1h3kOzmp8l4Y850UuGTWF0VDP5WZ79iBY+N85PSFL3H3Se68aZt
c74oaaiBxAccA+dg2A41IWb6E+FZ51mWBMoAePk3htm6k3+KhvnbiWnMpU4T6kU6Gmu6pZgAYZkc
pEaXuTTlqZlhYZh2IPcU/CaP3KY3Der9sQl6iD2GNTnZVIcGGGr1xyH8V5qqpoCcJSfzHYJF00Do
wkVdta4hk0q4xIGQWm056z6XjJWnypCa8y6DEPhFb55aBfqka52yCqnOwK2eUmD+Ft1lzjSDHefN
Q9YLV5+5EYpVXeKPC/CAcvPsLp5p/3hTLpBqpRBRWF/wAx7z58qRdbAIFtgPiOP4CVlUw1hfeNrb
mHfVa3KhOsABwwWAN/Zog+Z5bspGjKhLhfSL/dX9hrNXGAOzQTUvnmUitBjCCSYggkqMfnhB9nEI
IPjV4Z7xPXdA7WVWvKDlBAkMy8Ic+ZdU9HLuo16Hc1Dr5kmqER1D2kMa0nU28RnwAF0pFoTF+zDc
uTHuUdlOhj1T2o00oVKQZmXdlQBkwW9y89fVAKJ+MvFVYqw5O4JQ5HA+jLAKgoy6UERrB3iL+2F0
6EZFERurqdB/Lr8VOqDZ1DfuU2A8oTBxMuT890jdGVR2nFXyIjWZXuU/Pqp/lb4vVOkmn5kIYjGA
Ja8h/PJjV3qH91IV6Q18x/9NVm/9/vPG72j1otjT9TzJr2NrtsTalan9EuX4ents4lXWzSvBsMkc
fgGV21fZGXMvJyTixHNXwO5CP5stZ44iC/pVRCeGItSu2HhdoKubc0MLOZievHudhMORYaCEYfv1
fJ19Pwb+JzkaxCIcYnl1fS+hqQkWJnmZINXTGsZvq237kByApBR4t4I51iUMCGWxpLrKMLyxBZhV
yes+f+AQ2t+wjndCA1tVlzJIAItYu4X74SYf53YhUHKmFMysSZRKsv2r6gupddqYY7L/0ZcJ42T5
WgTluNIrE3n8i1PnYonaYxmIu4Znwq30MydIp7HkHHbURIgvhpNPOqxLwXki/zMICU/EyNtd14FR
tLrEKKp7VkL1z6h7vHqCNMZ2bmYoMIjmYgTur5cYHCbSRhvn5Ad8pi8qQ62BxE+MgZqTTLZ/pqMX
7G/Y23fUXOkoIiGZkYIUMnaqrbxF7mta2zyqEoHFbCzmcVXYsu1YkKU+p0FZHQKBQdVBM8Waaqjg
txcoK9Bvm68cVHA5+Yp0Er2X/urDmWgTIgIgKdQuTOit+ySEo1/BpYNtUt//togB9EVK6PGLpeMw
0XYl3fJ8Mz8tQgSzUWMi4lI9Wxkdus+3nWj2Egg55OWr7Ru5hxTPvMnHalBPWX14vazhN78Y6FNg
N0MDrJbm4mQbl6hALaU17Z718/hIJfT3YF8bw9LUX32+ikFgKXOVDJVOZi9cGA9OgmQP1SUTdrPP
4B/9vQ4Qxe8fSb+hRYURUIywV67rU3NhELSAuAhUK/95OvZGRp6eeusu1hT7ZEr3Kizxa9d63vgw
SxvdoBMZdaiSUHq3USC+dbBXEsw/Z4F6k9zj5lmOue2aGdboAB5tU5/N2fLQKzzmS2Hkiux2dl70
h/yFECi7rzgGxHVB4s+6LA9RxBYn8r5rYsCQELLwOyuIrWC2j2grBVWoBYLZLlbkhMR3TOlijaM2
TmpgWuI1pD0poGJWkrW3rZZK75GqHAh72KC71+64ZiMLDYqzEzpyLdCCtnD8GWnpqKekRq838WbN
23JaRqCRfcsnNyIQeIi5MFuDIMS7kozeiFCIooai14TbdCIZDk9Mh+0BeLqd1929/UYQAxKT6SXx
5PvSqm96D1Zp7qfsKxFy9uwDhjIDYvvQR3e2Sf1j/iTlPGmMJcIrQR8Zv1uAqqctjo2Szxov2wa7
5WP6JEXydTKMcZVqECBbAvDCY/lqnKms2G3RV16WHBrSykzaIs2SzMgvcU6TRV0V3Dp0fDEyhzS8
ID8QrNx/3Mx39hUe+4kZP6dL1pdPK9SlWzi1n/sH5aLlxq7YNBzxR//oRfrFKPEsHPw9Avy1qERA
fSS9RurGA/uaHZUXDBXYsRDHl7GSV1GVrJybF18eD+VgEb2QhZ6M7DB/4b9PXF+y9ZHwGu4Jz9Ph
Gsp2bC9TW43kL2vrXwzrjdnVH+eieOuZmPM0gB1kgQ+tV2jd+uwWliLG8XzCsS+VKeDZW6yd7qCq
EK6i8ox4yx9u+ZwBxlnWKUJn8u/oy5Dkwse3GKF1wR6Kk1RzJs+zexUbFF+TWIOP67xOhwcWimtU
P2I6/GwbeXZqK38t5yohnyeE8QlaLsisNAVOIvdP0Ls0K/d7bWFV33a026+NUCwW9IQocRQuLc05
apJne3IOC2A2MkLWRV9AIxpJL+wA1zp4ypHXfoxFeZzdIsfEHaI8loN6IRH20TNTEWqrdQGgA3YV
GwQ+pBWVbAZUhqsvStxgUxIIttPDv591FQ83cIluT2GyboFwMSLE5SE6KoNIhI+FELwy6CMZdPHc
5FEeB8XQSTWS7fFo9FmGvfvR1q9A4no0sDsc9cdO2E14rn91KA2JXATS5hg3QgR+0LW3ASjvh9CF
dlYNumNsX1OwBvKqoNogEwlTfTLmNFd86fNrri04ENiu99JKghkfS1BFshoDrhkHhGbmuQgYpw0j
A2udMdjebqjWWGCVnt6/AwAtUF1xf/J/VuDLiMpDxzklRFy/M+7L7S8zaG6Bj3Js1LqhFvZypYe6
py42F2H14+oEEo/q7E0cvoFEDH2uoPQQ6NZKhVkBwAmc7/Vk0abi8I/S+uxiCC74qaY6sKbnWWf7
WizbHr/uq7qg1Tla2gr6mVkFdxsFh4WDl3A5IXD/Iv9lJMIvSP8BRic3PyXbR/oygxxpwO0geuV3
eCTIvZg9L5v2VNZFWVdsZkJEXKfJYr6Eq1P/wjDvZzericRIxZnU5izzCtXjWYVfSDnrWJ9tSEhq
UIY3H27Xans7ZSofgLJwi5zrll9FQRU6J1bdfrslH3uznmzozzLkBX/z+AllvH+KcqxP3xOZ/hLb
lyqmuzttxES+VDdp89gim2caGWbeYhBnAFtJUkYXmNiRuKB8VFfHN3+ZUxpA+jH4JWiUfcSK1UbV
r66brNAQy7YnXV7QxEC0yM/V8todwqoVL/fI+wzzUW3M4ZKHyNxF7ZlRcOQzNqDlCGeKLrnwyi8Q
iILVDnLK3veJRz6n2dLorYTpdASfD/wgsV5z34C6wZsAI5xWCOkxRqx2i6/Em0GAmcSv3GbRqWpN
6LLjRZujUioCCapnoSj2ig0p+obkQgCH1HWjtjyEKk1HLHA9UFMpcogNw7pBMwx1+hH67zWC0I17
UBcGiVCUn1VmF8ueaWnzjMwTgQYJ/7H4qOucBd54DdlM9IkhMOJcJcFrttS5EzpC0vEdTB6xtfkR
4n3xkJm8EOw3OQskrssYDBAjzx7Gne7jTdQ56WMvb72isS7Ds2FZjFjcVtMVAfvQPMPY7BsqyCsK
Izsr+ET0gR/w5km5xPfh6U2UmMIXcGO6mz7Bb4EEuoGonxhaUb+LLN0P47M7NJ2r3xBtYTURYeu5
1CM9TJRrYeKYMT38EV0jDKm990U69arBFxh0LBSfOaQyQFkohKQx10cdXzEpdTcwT7iLYiQENUb0
Qlclsq0WAGXcyuuQSkQOWl7vnRTMRTfHGB2yZHXspEnFz3g1cozgPHD7RVlyQYt0qXxwylDkzvP4
tZER5wTsnXHwH4dtJCOEubpcO0FE+mK7CWn8qPfT0xMfyoDwfu+99KMvufvZRUXQuA1XoQevtad3
Ii9673N7orTqlPFj5hYS8fQRHh4pPis6qK2HlCbVKB8dHCk7KUcMUpObFCnO3JWpqSk1sR6XnIc8
gSBo/Y+T2E7ktl86qGXBV5P/P23IzmFOTmTZHcWA9jzDUZfLiLf9KXmywa3Wg8qy5azThrVAfL1A
t3FIIBAtqHCGf80hyncxlKOj/dM10MDk3y+g5SAan6WG/2zd+SqkxJ1ijYI2eB44Hw99V3DrQm9b
mLZ7ZIV0ZxlChdsGQVU0SY6hEvO9/XG1QSh/kE8pSepJGJ+1+MagWRe+A2hXSSo1EQ8si/rxfSQN
4XnqwgH65bKRhXEYC8AppZiYHLgbamiuUkNfzNKVfy8VR09npSFeqZSn1XI6d+smD7gnvRT1dgsi
WJ10vMz9nqVU7TavQJX20KoBidQADGPetg1UCLdXkJaaNjWjLuZOQHLf5ga6Y1dK2HGYaFpXSX5L
h4+cQ8USUUJxJWL6zBdJUIY9TigkCyRBkwZEhw+3APy6yWYQ/DXsjhxv62hjaJozNiugW5a/UP7a
2vVBFYAfr0aiDk0MIlURjTwChdE/ijvEXAHGbFoHzUC8k6zUc7FVTn+k88+5e2Uyz4sAQHxT0TYw
dqSTVq41YwnHGDCmWaRYm+mAArKpsM0i7W6c/vG9fMN09NJ7GY38tD9y+aeLhgJhyUebI5F4n5LH
+rPo0LkLnkAfanuE5UH7zsoLt1qZhr8GIVR+kVnUq5sVfPLGIU7+yKPj0I9IFUVYZeaiD28g35i2
dsZCcC8T8f0Z6Oc/78LT3Z6VSX3NlZ0ZKj7M/dM4943G+ShoTa2uG1AV8Tv01AS7oqSOsVpabml/
Ophp57ifa6QuMs9Kb92BbLB2cMQHtIlNuZq6he7PC1Fcd05HhSfY+ZuvDUug1z6W4IbU5He84ZY5
GPu9hOOjuggokpGuWdMWlyeykRoYQgb3Ti+C5TBJ8jPFqc3T61yyZZGA1etTvueO/pCX2MJXSDGU
9aOoa6g6LbIHtDGKdKZEF5SkCzxlrlz0TSvqiujHSMExe+UonavsIpHyD2mkZIHpFA/vlLF55o8H
4QNn3EYu5mujdCUs66Aik7RJk8wSwwGZsSwpSwr/aRff8sIP7chGvE0CQkwQX+dP13gJWpTIM0Lm
mXqOvjfiKeD2/7gJXoAozKnp+Lm64RPZE5/55C7Y7c0YXK1MrrijwdjA3Cyn7sPy4OXieCNmTfTN
0ZX4E6p95gxoIOsbkSSGtPz+mGVWNgl1JhuggRCIk6MoiHJkm0SNQlodQivdWiU1u8f7IVMDhSLL
iMks5Ks7krevX0QjEKEeqJVh1aS7cGP9gRHsTpgpC0IsXi71XAm9fd79y8+xswDh+P0cnRxqWGQk
D8955P6B1X/xILMrTdWqZ3cmYAjS1JaLAurVfXXg5kp2Adl72/XhwqFut8A4se3Xy4+cUQzZSfwW
iaq9naLr8bKymM2UIE3U5Cbxf++EuJvoVrGvHSCCs+GaIxEQpJyeJwQtR4FmgVn+p1fjNw6OKBAt
ox/4uWKSQUnpTROCZPgYN+XSTgcZRXSuNLfZbJ28DqGG7Yow/4h9LtPA3uAqqa/BlDpf/BrM2IDi
6CpuBvCwx5GfuWZ6ECo6f+WrqfP9LQfxnq3wStKiRfXPJgkEIDXAyGcahjlcEZSC6tuXaNR5KVDq
BglJ2+yX8+9mwgvV+Vjx5PtN3SKZKw1cSMXn9hnJiFNPaXqxKRLZL4uHImQsCK4DExmYv+zuBVo2
pY5HhtzjYJ957rTxj41bK0Yb9jtRCdrrYMwVdIa0UOZW+Xd6Dwn4+PlurzV4y/sjzZaQ7zr9+uvn
5OsMpb2ay78+UKHEr9v6K5ai+g5k3Z5t9Rf6lJLViDfCDV4xbEKX5KmjJtIS59QBVpVVwWcA7D21
aY/ccJ67p4ijK4Bb3SlkV18PBlhIpabmjXx+TEK6xelnQDMpwz5sRZh0w/+WvF+24lWD+mFHQM8e
OFvbOM2q/fH4dQis30/VyrXqpEjXzhh4N3z3p/eTdAhpGXSOz2qStdQ8wbWwDAbcjM7XwmNBl03B
0wZpeKwViKAiqMiY3rSNqB6V3Nr/172tXABQqrzNI+WsALRIzL8Dal+tV6AGaRL2sln4qNQNjnaN
biPX03qaa46Al+lpFGwnVwBIDK8eIEKovItddU80/KguLnCudSlhBtjTBwSbDc/CAGR1o0q5aGXS
le25KFE0CppDjai/qr0/azSdk0OFmjqaEpVbm08JXe9ZTiFTzZcyDWgLRUrBF2hHzBUmfSIQuYS/
BlTTn/2AaVW4a7ev1r3Phfiapps1CIlaV3FYhS+jB5CWn6g5SBuV6ZWFLK5L2trKdRIURqDH+fay
1x3exrnc6hty074EPGgGNjfvElVC3N01Qjxxg5Kh+A3pFTOXTsfDFB1Jtk5m0x32Ba42J+7nhaja
SsjCNFTXn7ai3CfA0MEUMTtEFjXD1ZryoTxF2fkPc6BEQ9dk/b7lkJjsyoPpptgagpPtxeY/gIn4
frvcTbKsLglAcVoh085nb52hNhrdkqgz1iKZw171QJYANnx6p1z5iEjthq2xffNiprwZXKgMwBee
EtQOqb2W1agehiCeGAZ5BCAuu5nh6FxQYtYRReUllRq4qR5Ozp6pvgUc2rQT9OueocEn7USC0iyU
CfWVl4yV3dt7fsFFqd5yFkQb8ld/mPGesbBZmZFenjI5T3z++vw53Si06KjJKlXBmy1waxL4b+1z
mmBy06i4OGeJZVy6N1LSfo6mMJF4HBVZ0zohdEUOkLDnspVwqnl3nKkPfbdm5brH+Zb3y/2bGFrK
WFZ3UyEcTgBgSJMZZmW+0UXyhgOnHBoW7gGCijFLArJQUFM4Ey1u3xWrpMpTT1PDsZN1qbMkN9ed
yivHzjVLLtsSlDotAcN9ZlxF7iFfzDLlV/jgnHaslj3bQm339C9/e0xEzE/mDtMm23MxB5prkY1j
TCIB5H5P8+2WmAaBGz4duH7mC7k+OePsBO0Jpj5o/C3MTELTXBZM7nQg1glZnzeqFFKKzBkm7AFY
M1vzbGljTpjbiMbNqKNgDyHOuo31cGoSl8i94ooMvuPc3iwtRPXGBko2UAFbz0k1SvQorSoob/Ml
zLhJAsipEjI/qNU6R5pmsw+e13ZgRYFqVrd0tPIk7o/y9etAHUkXY0M15GC+qvQBBBNCYYqQQKyW
pxkLt5MgHBLlw/pfJ2C0IljGuLy77/gh3HKHL63ZOYnJx5qCjcdGgmcb7+ihbp1tJAV1gV01q2Ek
oNAlaqO2h/hYRUaOeLitMIAdd4yYTiAwP9gfZ9mCxyzVCj0TysnXovnA6wn1X2fqtLRJxdH7kYlY
Qhknzjfrnlz2qxqI9qY9tVsZaeN8T6VVQwAIUGDlV8FZCRn3tPYNc8KHGb2a7wA3M/Qd06Yt2bJ+
G967H7KjbaXJUSCYm0B1wj1BF5AO7oAgNV+LJSDqcMwHEs+hy49GAHxLUTr6mEMNPD/YL1lZQj1m
8Q1e7OQ+J8pAID6hVLM0Bfc3PIEnJzOBv/LgGMb6VnGAbLVt98/2Kos7uy4qQlDFZZrdO4qVqyCN
XydRiO/c4rVz7NctTdpAHiNJunDXbLlboTCICJn6/2/6Ov8ryL73dIyEyDKNK4nOZJzxNMd+77ny
GRTMUpdcAHdRNHXKcOGDHRmecq8O8i6IpDJvyNL1elES4MzVrEZPhKm0aVOj3y1ka+KEzzTxNZOf
at5IyGnebw2oGAy233niJQNYkrYS9KpE/xCqO6XTmoTW2/iQnFgoYnWovNLqvGToQM85d/mDgVM/
iPEPCNCk7d7bYagrUWW6wi6xU40/ExMiZGpYkRWi5kkyJXbEv3tyJ+SWZ9jfpD2Z4fSeHtYu4H0/
CrGQqkjqKTTOQQ1Dx8kcvjuLnBg/Ra2HkPQ1urcE6k/bSwmuLFzuHFxulKhPGKS6Xlf+W+BXrv+u
+pkSmu+OtjzfbysvXUSVhtsuzJ+iMRw1RjyR+hV4gpdHVTnTGNtTjXm63QXPmjtPF8tLrqCjcwXS
dJTzUJrPXrKt2UpoZk2GFCDN8sNxRUc3X/jOfJzSIZuzbY78Wcjy+upm5cY/AjhNmGq+7zC8NuqT
5udNt0C8a0ouwZsxXuIUBq/5Ma+DLohzMs8i2OosvFQeRxzWFbXk7rWKLqgYahndWbXt6bd3i9Rk
L8aK7OvQLj6mZIF84XDe1U1wGzBEngadc1i93EfVl2FlfizIpE+RXZbnuTxONF4qq65y/BYwoqaD
hbQTIWWyy5F341/KEQfU74qOxzBLeLJN0z81BQs59VupSLiQiDD3lM5tApO8wr2zwv9NaVqv+2kn
617SWROI7d9kK0SMS1DHkPwMOEC9T6l94STk6XRvaQRQ3+HgkrCgcD9FZ/bWj069AynA+heddPz6
F0wGto4ZlIlUNZrGzoLhX3vM0/QfZz0cXcN0RtSCAr61kqg9s314MK36osHgrEpF3s0VfQrHfQT/
Dh+Hpo78zwWy3YzLEjggc+OaXhY9iLFAQTw2ZGfJHQrL3/pwf8rhIK7MG7qV4KtPtPlri5Act5IF
ZIvdgpgAalSB4eOOS9hn0MNZOO4eaIWd1hgpTiuFJCjwEASBZ5o0NVyQ4MiGQcpfCtOGbv4eLWQJ
V3coIXXzUuG7WR/TRunLNMSn/e/nDa9ZbuBIa/ese7oDOySQz9Ep7P8draTX61UQ2SsEEeNxsx7G
NifBR2Sn6GhDUJ7ua1nEurCSjqUyPrkQGGE2FyGXpNreM1tWxtniVVYmO5zwILBethgV0wdJpcxT
U/JIZ4+vK2WEJkNbBuF6e+yPPjFz5jIiHdxOMmxAnqHo7vA3L+ySZcEZVIsGBh222nEhWfxWmFkQ
a58SsXQB7VBaCZvi9FXdOpKZ9nHKHH2bmRC+s/Z6YVaqdeOIMZErvezQO9KIeHQ1ZAwGZx+klKwr
tzrqDocpnyksgeHpNf04Gy5h47E0YSkZSRZlIIDu45oV9VxXcWgM49nq1cC7frheQ0VJYqQfRwFo
H8irCuFQmNK3AZy6nk/mzavGjrIFotpeh3m4aeROb3SvExqzk0iBlVbmSWA32MOqG8QwQr2EbmGr
QYjQW89SfyqCdduzv1W4Tzo5DsWAsI6sVSs031Q/JBfytnnAP26Mu9Iotm72C3u8L8h+TzCZ6EMF
lSDp9SuOdlIxIW8U2zuXuq3tw4nKgs6BfRqeBKQA2bXjS2TJuVmtOofVcvlaKUpuzQovX6vAKkIV
TqyLNV36OnSl1Q5aDutSIJhTtVGpJAKy6nYSZi63o3J7/wAdkTCPFV5gRmwtfLJ3qFuIqvK4MFjl
UdURIHdbfrESX+ffZ6xPgWaT1ed044z+WVyqnC4TbYrPBSGGoP2CCKJTQ78/tu66HGm8qZefMwOT
jnDFoJLvbfsZnXWi1yXZ3p5aXZ9WrUtIKtY4T5dhtaYvG4PRDtJx50MN2AUep9aymUUQ/kQM8WER
GIhZX6Xt1DL3AGyQZhoPPI4zTKWm8Ur9Z/tNjcxXSxyCdxpd52XLoLNKejyJizVFjxrz604jr5KJ
R9Wb+5oFIqf6gRkrI9kXpPMG6PELHzovWG+xltBMrJ8eB3Nz1D3WDoH5x4/BllyfeLI2K9THVx5I
3vtsth/tkawEcJHwV+FLMLZRjGW8WU12Cl474Pyx431UvgjbAx8+5BpCPkKlmflpl85yjJbkbFOn
ha31NYE7R8AxShN19Gzj3NFf6z2JbhkJOh7EYZW0Khvs95w95Pblk0e/oTMgh3pc2cKT7ceSwzXk
iEgRKBGtPu7iHrPxapOxwmlnIMTXKx0yHL8FF1Uz7Q6D96mWyx8DSBqeoOWZSmAJB4kfyktdotfN
bQMMKVEtU7hQmxKZ8l3trXCnX199Dnv+/wCV6RP7ETFUm7nJldoQuRGr8aDcuLFbUsJGkWk81sIX
pJsBV+vlFSWPZVQIdGR2JwybgmfQrFVWHn9rYvLNcTRG4GeVbZSpk8O3PryATzIeJPF03qbVE1g4
CfutI3YLX6hXALupjpjdkXPMFmT+S/r9lIbkCKNgkfyE/lQfpOR/ko2Eak5pIDkLK6BOwwXtATQW
B/b6a9hlwiVYHKLAOZPDGdBF35LE2qhYPkGA7FtIr0KIRYd8zwbk+jD1Ag33VRdansGRoLCF5ikP
oWN+gh+GvFe0gFjFIN2pyedNTtFJADoli/me8pgkbHSRnH7hPTpcPXtQC6jr2qGovd+rIHX/+DHN
nmOuW7Srs86R3g8TTaSq+7rKT+M6BP401mTVblqmpiP+D1ePBrNqKKasw1H6mhQGB+JplCUH3dmd
M97+/0naBIIctp9Bz7xPJbC90HevWGG7M/tHzQTR7arfuxpzpY4iwTbJzMMIFfn6Ns46qAXXQgpX
YF2jLEXm0sRxwgROW3DUbWyvKP2vboT140ofc4XL0aXLzlKmprego10iTlH7eMzo4ZwiSjjVBs+O
HFK2YoWEDsbG5hx/9wiyBZZGw0rAFkXz0DofoqEC4R67KQ2NaQWIW4oLZqTJlzRm6p4FuynPJctJ
QGCi8MCskmm0rm7jPtyih5lqvhjiOgi1jDK3pr/r2YEaFdmjhYiiuGpBIzpID7305ROVCKVjOUSg
6k/BPzyv5kSt115STzncf0dJ8nvDuOePqNSNUaISj4E4AQ9UCyra/iNTlJI9nyiAQi5mWQQGa/6M
V0PATkHduZWskpWliyNeg/DsAROAJ+SrEY/6lveYS3UNAlO5yJzHs264G3EuBt/pwGAm6dCpZ5ly
Y7+aM2LH3xmDlSthjlbuJDH62ISZtCJnlXuHCaj/LQkk8diEdvVeUtw30Oz6NOpLSCWU9+iTRdwe
H2PDsqdXzzBTGmYtzMc7LtnWz23yTZlO4l3BqoZfM+9kDhiWaIS7RTXFj6gGK3BSBlcF4PcDEoCR
3nvpiYiB9N6HCGSBVISNFmoDiFjW+xlaG0Ur5/0WuX3UxNbUtLfSBYOcb6RO8v2lo/zsRVTBhl49
8dnemTNTfSVlQ7bBh5TBK/2j++y7EoRG62YxX0ecNNrS3PrFe01tKuoJybSTLDzeJifRBgaBQf5N
RkoTX24WlcoV6sKCYSf9XR/Fm0k6tMT6xWdPAySxPYZazdj/oWUl9GGpn+6itpkSGlNoBTqIbe/z
gYa14wQ6GPqFpXHSCW1+YeV1NiZDVCuDcZu1nnhszl4E9nQMZYw3S03pJU7rA0iyi15Ffynr/3SY
lV3hWTm79OHoOCiHU+KnbYO2fHJl787DombzKYK52ven/k9A4t10eZSXAd0tDij3hX7Oh8RPYxsN
zk9uNRiQFrYydj/0U/CGAEOcObIvLVz1l080KaDkOe3kHw3rFP4FEF4SNmgz4T71f7DtJk7fAMzJ
54jdeB6ZR151eRRcag5ho+o5zqPHW/QT5qP+UEpoWLZ3Zle0dFJlZIAvAzfherMfsfsWfiArJ1/Q
6+rjWNGOw3DO5ytpR6bYd+stKXwtLpzN304gln84bWU6Hkapn40iDN9xjDBspszWewKONTM9q6Nn
/42LdUXepGVH+zYUmzSSjm/MJ3MkVktMeIen9C8HV04s91YaHv6GxqMk5EX8MNvi0LJimkf2Jpg1
XTaOATPld+EVaNxBCIQc9RrVontfHW6+olx2MyUdTvCFJR2R2srKNOSrZldhpKAUysltCFzMv8HH
d9voq+PGuJBW/idMLSQUQNxFc6OCpegiO7FUCTjE9OVc83CWKh0o1KcnUaoVIFbgdrPNMbvI/HRk
Pr1dA1v5wB5OMarrdAYXANEJWZmkfYBjDqwCghf8FED3BXkMY03Eiu/aQGFKvO6rIPVvjQg2DQz5
3gXWvri/9erSO2+hj2y3AV9vX4aWQd4knB6Nip756QFYucK/ijcOqqsZGS/BifAFsRgrPAAuov4+
xmdY4EJ3MyFb/JtZrB/BqkiYqmN+8ophxP2VJ2mpyo3/oYuZjNWuxYzs1Q37jUeJlsG3EufP1yff
avszeTm6mks3MWuon1hvufIkFGePyHGqTnAGJXfQYRc8+ToTywJyoiuPb096StVb0QmsokfLgRCo
JcjSHMFAG0VpJoIsN4BYnqDlK/YEVOa8axZAUzwUftnGrdHhDMBi0DcJiBMgr1N77T3A6uiXgEgZ
UqlnZDQNriHcQ0DXY8sx9qbDP/5PZvaHJEhQsTBG820my3BBCMqpbmm5uN3DlnS2cDuJ+CnarjKu
qUyqKcPDmliCfI1Fsg36wO5bV+4CV5ZRDre9peTIKsSRwDPRa0bNLPaAwsVCg4+uaqnlDkP92Dgm
NudSYL9XRwl5W2+g05NBDHCf9RthmqUYOlZrCYQc+WLrxvx/dpT5U6DAK1Wi/ztbngCrPiSxw0bD
qUGXdXon4f1qCLxQ3yJGZhlDtbkF/+Xy6Us85gqxVmQ9MVD6y3uFxlLeiF2aSHBBEvOYL8Smw9tg
MaVPraG6Otkuh0y09MQ9Gq1nE0ltBi3simF0zISwL8Zk11aWFsluCezkRJhLYHEBIqvnA15v2k8M
P4UeLSdESTRvz5ySmW2aK+R/h5h+mJhMX/jaY1In50l0W5yCdxi682Qi3A4a7+GrHsM7GXV/26Gu
1RMtZJob4jNm0JvnRkt7W/RGg/DN0GogbEPBvDdqhUYKxod05U+Hn8F01BKoB9FGy4w85LAhkcG+
HGs3nNqXSdMTr1PECoCDd7P49vAv3+HR1vynY4aEl5f80/qSwRzeVLWMTKQ6puVLPU4r3ncR9nrL
uyk7T8agiBJKvGHk9n+Y2SQZFcl0AZE2AmnUno0k5wJz5PxLK2L3fuKW4tHzD6GfbUUK/QDJtlF4
/IOGVYoEn4vq/NG9VZ19K33vDqq7W9ojXp5h17wAfuvPEe0F5VGDxIUYqjC/VxMGLgnFOupSaUTM
N0DNpxo4o+s2wY2XCOpOZFRHidQZ4au2JJOLK0RyAUrc19niIdLjyAZWVPvHqTRuACYoI0jxBk42
HrR9eJ6zmqnRxjMOgaYjtukHM7C1b/7hGnGjvgQSL2dIFXeP8Li+JRH9r5JTk6OpNKmXY621dH+2
IJoy+SzMP9EVPZ1DN+S+yQsM4U9+Y9VUSlp6dVnDClxTgXKA70Fu2bF4CexcG2abNw6jVsTjAXpY
Wxey38K6+oDh7xF3olKZ8z3hUMK8oCA7ssjeGv0mdBfOnzNp6hVFpkL9IY+x8WHkKijOrxwsTqhk
vxBdVtDmzAGiu9MHB2jwsDZbhpFK66JeI92F31aKAZbKxiQYpfkZmnNsY0A9eqCey4BhwkNNCvEN
kRzatdU9DxaAeTOP1NQUWvcszYqb/y44k8xBHniy+3CqbQZGdzPRA2K3m9r6Eao3rKROPslo8VMB
dWs8XTv1rM5qHWJyWFAu3B/DgFvSQB71phxa8TC3/iwtotw04//m8i1qVDIdvf85C6lgCV9UmDwD
OhzM/ZvAHILABroQeRxy1BSOJ2wce/UsvPMPHmXgIYyo26dDFKWCduNQLNx3y/pIrA1s+W2G7Qj2
ZqZLwEM9Eg+4u+01MNkrD03T63Z129DyqxitWNtboYMoWIi3WcXPNozDvJFaS1IWeIF2sxjDCeQk
HR2ix0lbk6Z38jsAc6SdcMjAJPf2WRYGNKHJZf50G0oZr95aBWcy/7s8amliyhRzMr4g7Yo/fvnL
mduE1njQ9vReuRTpnRu9Ewg8BZchZVlrUrJu2Hz8BhcwhhWaQ/1692TfBmJTnJVcuKoKgSckokw1
6AU4dXVI56Xkkj9lRGQeorcfBLc68/+OTsFUMEITTKhyV6x3Fq6/GuWLY3JnrtGVZ/AgcT4LemRF
bcq6zZJ+mIhVxS0hCopk2ZJw5fohoESt1dqD+2Ll1cj9bwOdogcgSFZvYPqpginoVlRd+8qfs0Zo
b9YjGsbg1fJw2ookTzF+s3w400ons1Rfq1F2oHO4eOSrbTseY/zhykdWsp5NjQXNnYQ+B6rZlVt5
6SQe4u3oEZ+felgoyJJ7XqiU6mK/p5z/hcmxgTq0jzzea90tcUzUt5Q3rUMGafpJgY/CUjhisUnP
GWmdQU7FGy0fhg1/2+MN3wzimGfaozacldtBvczV+uJ4ZAez9IY8UcD7ZqxPNtijp6Ae2uZRiz4f
x2xriELiAZtCmNmg2c6Sq6rg9NqpSu2XO5zQuJ0EXRdF0fns8yWztonfbjQUKNx+dOoslkRfNSDw
DbxJ84jYSmoz9mezGKzykKkYzZGt//9vsnoYfh546Jbu0V/d4YUGDUg5ZMpzvT1+pwBhU0lytiMh
hNYFYP8+LYmC0e3oJtu7H4JVH1lBjiec5nLYlgDAiuU0UhmADYfy30dfGSZ/aDDw7lbyzRrYjX0C
n16W4Mz0ionXitoTLvhwX/DBHQN3XriML8YXF+8gCYZOPrBvOF7d1cNz5e8jhqYVldAEvhB1HQWM
pSaxzSrzx8VyznHyFfeUpZM4hJ1dpjh3UwDACSMx7KNK8m7QUDf5qcMYhCdeMhrlJrzz2AO8Ydaj
cVL+fdvRZ/w59LUSDjT5WYBNZaqc5U+04fvnHUxJPJ+M171d8/Jd/VBGuCZmkt2bpkTQchfI8GeR
gdXemA3HFzxsf2YmXdHA2JmyBJL7rdbHMFDsWbTgSfQA//IcNL5zhG9jJMqtCeojuoLg+y2Qc5E8
KpOfr/RitSsE75FyNIq3e9Rhh23EcewtF5E7K/7tOmrRC0I16mze+Rb2SfSg5esLMuzqtLQJUAdR
0orIuAWRq4Vg26cK4plX6tHj4S034dD4Si1mkOcposmGey9ueLbaVWOtrqOh6DcQWNLaLZJ16X5W
JLFR5TMQyiJSG4BJa+Kz8q2BrVHtwc/7U8PtQCUOWMUQ36o3HyLEYL1KSJCjg348uhwshAi8a1zT
A0kMAa3S/vZ2raeJ0QxCNxV6iMdZIVizVeTfO98Mlw4gEsha9KBoyP/t95rvNJs8sIgm8+BF/mBU
us4MKzM4lwXtQntEjdLKyHqN91YUDywPoHAZJcUb8xNPY1dfgdVqcyda5vBAvVFxXS59Rts5b1Nq
eUdt7+BxnT1LYfdq8nEdwwjrexIQxZZnn4GNuTScUMZMTgL3rfA1AShFjxK3O/no79SKnaSioBns
8vLD614YeVbDzCI3+TcaLV8k3BYtrzmOxhEz5UfKkWFCZwLCjLGyZrveadVyQYzQXtGUp/4H2FTm
2F/e0ezbQx6VVcdwW1Y/k7vK4ceWJzyGa3Zi8SptbPcf7Nmm04hk9lPky+Qh9tWFwGFEi5QBpHFh
PXRXdP3CDw+Qm7hj9X6lPcsO5WNPWMr9BUPPO4L4p8JGAqRx3sPgP51sg5ES4qZymTztxGGtj7x+
Z89PPZVJXWkk+d+JYFRQFfx9eBBhMxbCr3LrSq7riw8rscRk/bkgs3bOn8dR8hfzbGhYwWA/LavU
h1fg6J/XQ/wBEgcgM3p11oHa9sKEC+gi1OfOQ0kOTMb698wvFifj+VjHvoTo1upe3oJYjDfRHQtA
11RB0F1/pj9LWaoWVWD3iXFZ070QUsaaSBlQuJfJn+kUPMrSBRkmk2HqFwEUVs2m6ZoLtuslD+Zt
HSHpvx5Bk5oNWg2PeQIkQziCNyzoSQK8+PurfDD3OYbiL9LO5B46lctcTTF5PJwoVrxg07Wnh5K6
KXuL62OHGZicOgSZA9j1dfSTvDuX1522X9OOQimddrPWCrry/I8XByDSzWM3Eyf69icpsi2Arjf4
oLo+qoH6gMnblw7SOEcHQwKxjc0EijIpM5VCpqRQYPyw5ziLh1n201PICNgffEQRFgSFBGhQuEVc
hn+WIMPV0L25YDvmLHDEuZmsjF6pCvVAiCniXph/YsaQkCkqzpjKqEzsQ3jArni9rWuODfV4To8k
Dgh9cWw+K60jBMYN1vKX1BdMTYKGFnqVruFqew2bC8kYD6H6kIv60XdrUS0jB5GREVS1QLOws4Sx
zeafC/oW7QdpnOKu+G+j8K+JTYuM0+Qln/ua5FlHCbTnvYFl+NZTehaivmKirSE9cIU32+N/010F
/NGbFwQ6qMsAh4yGQGzHcI4rnG/2X/6zFlzeMNBt3d036HVq5LPJROpgtCsvA4DKZTJHCu/b/Fn0
Y3GZ52hh4QIL1BugzsMsk3i04lqIb1UDOems3pLWS6p9gQSUbiRIM+xMgyZYwB23rThRH0xqRMZs
45mvYT0LJK6DollhsRwBY5lpXLfVSYEtJxIJ5YuzMXI0OJ5pkc0qOwiBwcfrofDg0AbCWXRx5sXU
PkVrrSPetFsbrg+wsAxrGWEh8t4mR8xpnqej0lBt2JUBp0zuLReXNZrjX1KiUvYyGx3gUD1crKVd
PXEYrwOyazNxeQS5OaYLs5523LIUtJ9xSh+tvVjEumXgkP14WsoXivLnA2NWLduaYNpiJ4HH7QfD
2PUJqjJ+dvvQx+dJrDDqLJjwLcJCqbPLyMCJDm5A3zpxY18VWXv2tI1SeM3pJzeogRMVraRzxLSO
AYh/f0KsmmVJkO9t1bVIICznmSpNCuhyb5cDnoO27uc8Yca+7lfatvqDKP5WoTDwBDdESJyTtqh0
jPZv6i5+b4Erkgi8wXyVMxsbevn4dk8p/IQ9rDGw/CqOgPky/9AvixnoEX/da5W5q3voUj9f3l3U
CRdWkEuBvwk/bx9X0ugR9mDDANIyNMlkNO/lGzoBzLuXG71abTsO1Wm0lQfL/e2Y3Z+mBzGTN1/Q
j8ZO4rGpz6PUXpYryxalW2lxxxWpLAMJKAvw+OYXqCb8s0HXHtb5R6iYvYhgq+a5OBbq6PuNGOl7
eE65ybmHQ++NklGOx7iPI79s9LGodvXRADdueyF3+pQRPCqfZvqKmi6ZWxgPhKfAijTC4V0Fu5UK
joShazMbL81RL2Q9UkRiao3rx10IKMYJmlaTruQ8wT7D9QCp/q349O+eYA1j2imHIaTvUSQf2B2H
EQCQV8j6LQ7Pu2fQs/yl1ljPkCZyzi2ACAESRGDqWK0Pc7onUkYTfZg7cIOU/dcpX/rhFYcRz0Kz
nVbskAS6GSQqlYyyH4Yb4ovTbIIf6qoS43Ptm+PlKoRHrkMjPyQcFRT0qEFAGoDiL1sWrgiG5xQ+
8ItU9WNXa4bJtWblzr6d1Y+x0o+NEXkW0WrhvuJfu7689OB4h92doa1cANzGHwMrpNTT58e3Qimj
I7/lISV02pMAxxOn0VMjDPmTPerT0tXykV4r6SbXkfrwZBjNef+o4Bv/MsIAEyIakAOxXbvHaqBs
wUQbiwPywtBUXX/zxdnzFbKeTWRsjvdm/zuXG1vHB5EUeFPT5XxWLto7/e5000inZ6DJYlgadNTC
pia2E3GsZi3DMUFM9T8hYcrDcmy8bAWNI9BcLlro2SLV7hzgWkngWa8NaVJCPjpYL+S6P7r7u7Wj
ug2Fs1Z5oZJPAR1VdxWgb7wAZkkHAIg3OSkqpgLsqz18fqSu96JPSF95NWtgIZGazA1YiLkV/p4Q
zI/fZ5Kyv4537KbGNns8aA3dbdPQR27UcqRi+0COugZt1P2+0zJvmG8AucR244MQHzpB9t3eF9qQ
RcdWOHZoRZ6HnURP1uWNlYNjHYwaTx/lGdOPJQbyF7nYLGoepRvV5EtDOfSmZd7FCWfwHbDlzZTd
RocvgIUfmGy20FtnRJc2WspsbnQOKXuHetDO15qMNqlWVCy6f9Og6SBDo4Tr0gi774IXWNoUy2Zi
SM6qnTepNNl8FLUovdCJW/LKG4jlleQ4UB/p4NUeDL4NR+glcGgi51zB43/lAAS53It5AI8au5yI
9QDvxUo+/M2x1eAoM+vmyFPallBkHSVDjkhNd6uVU/RTO6qkNx5+OYBfymGpEJjBXP/SJ5C+4j95
yM7o+Ky7C0KdxUmRYsGhMkzQsLrZZluv8pLzX/I4HLxSaj+KQIWRgnpArztXqqHvN1ILmDLQ2CMr
UYCloFPMbxWoi1hogthwYktxAODZ2G+inwYOBwDRO2A96kMY9f2Pl4vMFyp9Wnzc5031rs/YHirX
dyaEf7tnX/9syVQj+bmTSqc5eZOrV/R9tTZnnQyvAFGDjMvQsnvEZ8BsnhhXPwnmzBfapUEN8zmE
u6zH7wRhAfJSxeoWc5mpwOJzIbD13+8uSVqR5rtLdwqITSKGymDSd2UPBa1w02J3+RfF2uzLdPQt
gcofaYjZHFny2UhXNW0iFhhfsvi4rE82aghFhWquqAtl45zcZYO7bICM4D9nggDSOay6UwW31Wzu
w/C6St/WOCBB7BKAegUUjKl1oviCCSY7xBR5t8F3MYkFrsGNPjaCkH8IAK8zYXDqh/MJWOXy+8xL
gilcXHuIY31xTTvMQeRFMZBy9exXOFDitlLiaFPXSFHzh1YqOoG/14KLxdRbTOpoA8iWb++dZQKx
QjrecTUmcCzN/YoMxdbzemNFET20+AYr/AvnFX6cQNvVCRiaxnIAu2dNfl5cNfHybcFjFDOjADM0
6K6ZZt2+PEnxUFkNAPgF8ZIvgNdqAFHVL5ytcsBUZ2ly3FSgwxXltsT9WTXFus88jLXPCLgbpDT8
RNCHvJqxuEI5NfsL5TIHl1um3P4KFYYXMJ+6FIQZWaTikMz7/r0R+sAmnL0BF89wzN4oY3wRygLR
wpJ3jV5uiDGsTahmHdDvW0wROKHAhDcMT/llXpA6i0Z7zm0KilauCU+XWiWUQbVsgYsRi1+PpPMA
h1IkYYMC49PCHq4u/XwSAjtZPArCM/K+Yu2jQonwpmpwKIyIDVosoKiEasUDIz0qc3taor18SYzJ
qNm81NeW2ogvqs9M+ZNvAT89bIpFSdk/Z5hRRJJvbRepdglFI2vf3tlqIjYO91XSv0WTeFHRY5m6
aqabHhwepT0DhJnEhmxxgV01i3zT4RJ913sUbqodcM9/rWUGtV+M1r9OTKMPjihK8MAndM3R4X1x
QHspV/GYO2pOhXkLBh5pM7SkvW3mIcL+JMQUI5FfscnP1n2chDzS4iEuWzPq4knK+rs3uTRMHsR3
jl8pfCp0KXW+8iUGPsKqfwKmJVjhLD94IOBoxXiQ19RhRSyFSt0au3htXKojU2tj/LKbnNuhHy0g
37SPASB/rZeWRKSVEbmngzHOFIxMr3D7VoL3+yGVkOpvaR3sJBBLfU1EPUHXgPVVH4NTtgcYchby
5lAYVOncSYW10s9dr+I8PwbjOioDR97X4FzU5ZavG4el0fKwbPpXWxzs4hKhwyniTp0ls4wNV4p0
YxBqO4BdAfi0UMGQzK1N94uBm/kFlvbgHVT+Zz+i5Hchr5uJlu1MheSLLSGinnOfFUWQuNf0sfVr
2HXpyHr1E9WP45ndCIY7pYeH23YaSGNg1erz48ZuCeKFwe3VA9b+C68pE8AQX41krkEHYJm6kggu
wsJhU9AOUFZzF8zMvPvpN5RK75VZ5tLWOB6EueLpKumks1sK8uUE8kmchTKS278pzkxPessh9Cg+
c3YeY6f5SVaSXEvHnGpCvXhBt7eYHWc7xvpwZZSMZubecTNPBpjuHkFc1pVE/9ctewbdaXSMaJIs
FsLZ/Gb+UCYnk5WYtgyUy6x9JJ8/OTIWa3AgOSFiYuT/J86qqehrueKDvwCsmu/ZiilMsnS2Jpvr
ZvZ4VECxhfeStkDnGAu4k6zHlXsCYKiElb0/+0kteva+k2qXVjCfbSVi51U85IpFJZa3fG4zHi9n
UH4oQWEkbE2s3NE3PefuA+bCgFvo4jZbMjLD9SJzY3jIoQKZzv+3MQkI5hjRj/ygmAH8TwZ4xvxt
WGl6OVy5kiDyqVKm9HZwLRCeOr4tbclsqZ9eJXtINO1rvPvY5zvLh+7JppfbsisreTFHv9o5vaXy
y+xf3oPgbzfZO0iaD0CCyPGmlqG+0Z28tqHoHGgWmHd1igvkmGVPER6cVYrV9Wb2GvYBCDd7zmRj
j3sqDi5cwfJCaOKGJtDz3LYB3oYsidjt5it2uRbzJYoedrvO7OsqRIJsNi//uVC6J8uwPJSK696w
puyn1SqWlEVpiVXWbQw1i8Qy/Z2GPArSIu0Dea9v8QNVj6I1c47CEfDjRLHn+fpbEO5a40VR7nsJ
V37rXTG47GbWFnG+80Ny0m3YzDm9le4lHw7fGEV1vIC68fs0dCz8VDJc1s7F9q8lMO9w+4I06ztd
RGkno+BJwEXUutXybsQGF3/j++ZciayHqkn6JyhDAbCSDnxhsHiVM3gFF8Hvod82Uqt/1BGV4p7/
ehVWYluIl77hxrR+DpoCOZ6XjinxthMZkzgFAQXn0E/2d7gVFCZw4jhhh1LeQSMXX418Pt9A4BSL
r4CzLttxU49FoovOUw6lHoE1p3pi10ZdQrztMqphP4ehs4xbWg4Bs0UCF8DZNy/lsLSnxNQIxSxz
L8FQwS5ZecyzL6KicpO2vKu1bcWrs+ENwLNimVXsjVCjKZEP7CEB7ycFZ3fzCvuy5HmxgUzDye1C
GGRJtfGBo1ES3hCd/mNoYyQLkt+ZfxuxmVY9d+nSv3KT1lYGcZzry4SaYyKZbBDeF96WPWQ9bRFL
hR0vlkKM61Jgc/mfWlfCg9peX6a5s4F1fQVkIIVPSuKms5G6DX8VHjkHKBFLrVhsWely1eOiY6hB
70zVBKsAr/PYhXyaPZ2WYAbMrc0HVoAsQUXUetCn1Xkd24r1RWuzdupjMzOAGivQ+P0qMcrauIFE
pY3JtDZdKtjVgk3CMQBUY2yFwsozX2dRbaTt2Ka4Z2YjD/x5TbKW841cHIEwOUfel7WIzPdwchGN
mVA9bDE7i10bJzLAWY9myFyrbETMFULkbbScrNQlLn22YBfl/8Fa6a5C60jsCOANX2o0prJM8r8K
azRpoOa7wye0IpvzZd+ntYJRmgHGdVbNs5voDlrR/mBasaZ1HexW+YbEcUXz31Jcgh2bDUsYbPUS
TlIBJx7lUvIfqXOWACiQZpt5xG4v/nyEkKo8Dv0ySX3XmpdcyduEppYueiesmRQWm6dSRjRustqX
wn0ujutwf1BBjfZ5vAQWqWz/MwT8RQduLXJKbqyJUJkqTdCMtcdQkL6g9V2FIS+QbRfDdw4o3zHN
s2rjQLooOSTOEbNQj1Vy8XHOWwx/wlHTJd76Hbi3S6IG34YLfKfEy0zKzwkpPag8jYQcp/M9zUcU
3Fs58Y0kcCXnXdEd7vXxrXSKW9jhFy/nUIUAO7w99us1Bkt1Rnr7L+TE7bJbAWPXgh38SUD/oOtd
g5Y5GQ0dPlqVG4FC/OkxRQMUsERHElsjL7SEN/Af1DrhoYEqkM+XqXaTKmtQ+dNsZIeT0/30oNZH
wO2P2HoBx+NxhU+at1Ye2C3eGfBiFZW2bq/U6LavwmZUa0AnwBqvEx4rUPCNt90lm/N0ut/kNkg+
cB9fBzHL3zS5ihGl9TyJBUT4GlliNl1kPqxV4NBNmkzR1DFgoGABxQbSriQj2TESenPKkt2jVc/V
yIEab7LdENnWaQ3bowWWo2doTSU/hhBUXS6jXLO/a8DQjBUbdrndOmvJg5AZjwffgfO34lf+81TU
VFKZ4T8O3l3vhFWZKtnsleqzU1j0NDZgNU4GzPKOmbCT5Ap10nrUgrAeFW6U4lLkpMxmzqQqfrr7
dOc0KnoczCxSYA/f6xVmcdaDQr9RLC3HCc0NkqWwkQAfuopBoiPJpIWihoviv8XF3ptHjjctGGUe
9Nvl6fBz6pW56z8qr9FyA7TLlCCXUqxjRuodWV6cd4psEcoIey0ECU9prKLBPzq16VvfTriH81Eo
dg5goBSr2ySsbzMrMF7/+ZKKCdde0BghmQm8LCcaSqDViPVtaVenBcYdXcTY+trZB3Jf7B6oIg1B
FroNUpweFQtW3nGBrgQPjThy5kTfd5ARfwo8X4ojG1NHjqof4cYmflT0CMQRkW80tUn/cFtsXrCk
tcRr0XBvKq/VhOuY3TUgx7HMC2lZRa8S6ljXCz+jD+tgAyjI+OpL9MOCTmHoVmasWTrZkHDa9TKH
0MFkxdYl+U7lEYCEP3L/kcRDejdresPYQrFsJLABp7eHfQi930FqsrQXatZgnlL4HJ2bu2xoSxjS
9o3ciwo3nwcF1FzJRS1uGvVFBuOaDxwEgQ5lnjqm5H3BSdsykbfiZOx46MuJM/tObMXDm3NRhsN4
0igst5IpIHpbnoOR00Zw8ZpgVmiPt2tHSQib8cnHecyJ/oRPkH2GrvRZg7dh9CYbhso9V3nzVtSV
n+Iu0VKU+JiF959TBHSs+ZcWYbZptZjKsCWIgP8iPfM9JQDpifaaOuabXpX1XFzTKXEV8nQ0vt7C
GXxUXagQ3o3FOmA7sZ525LfLD5+symVJ5f8/mLvn9MNffCgGRF160oWQbX6GKDUTfrBj6ZsfS6DL
iGUx8B169W8KZoe97sFf/R+MbeMmkY308W4CGo34oKpwt68fvxxmC2pzRpdxN1cXamGAhZDYiiuM
59mRLI99hIQbgQuFqhzDOBFR1P0wSsWfKe20nFrdmAAEZvHZHAvfxq0BDbzMHZD79S8j0VgN6ON0
2MFuaw8FbKpTB8mzRv7ZrSfsm301V5ANxvYKesFTk/ziY529Ed4wCZKgtbfIJ5zfCvVdSkYQUp7f
G2Vt/TSFcEo4cE3JzhUSFJclOY+BZ9ecAjHZjXNQ9hVf1a3Wun3EzFvD7je7AMbhPUxjRMzn37Ma
ZZYrS+CC7Ij7+Puy9RKKoiauLCEkk8ko+qnhf+1ghi1/Ws3UkI6wdkGgsJWcXv5OpDj+XwK56ENb
IKis8HgOfyVwY8fyxsK2F2b9AE0pTIhoCDi5J6uG09WHbgG29qi8SkZvn6VkE3e7vfRVPPv0Msed
wAee+HsNUUkX/2SOO+yRHV1RjQD4KpdAc8EZ2nTcCOCdUH8vI5kFeUVxbb4ovCQ/fCpJaPu5Wm1x
E9VL8RD8daAPFHcCmokiysQq4oN6b7T/1DJPXM1Xy9D7ExFoR/yYKjU6o+mQ8xHjbd+9NPDzhRo0
vqRsdVhkazyTAz9VOlWR1fVs5kQTpXXhNPLljQQ4FKG8QyqLrxF4JVBIr51bW09PLjgSGWejMpBb
KqCwKnqpsSRRb1yNByaP7hHLeW5xT/8nEjtFCHMUcMQK/C3Sn0XJwCNCpPQdcMCOprHeCKaRt/k0
kYoE9v+BScX3FBDMgDoqcTsth/TKro4gka8BeuSBp9/QoSti3JMaj2BT88X2BAf3SM5dTPOGUJqF
U9KVOHQY7kUI8D1bNv0ndWuSgRoMYg7Tbx3O9RL+Kx1qyLMuISAhAZ3m9l0aZqVqWn3wL/Wncg3o
E3GgnSdRbut5qeIgLRZu9piVsLCtreaI++sIIOFw/QajDY5K7w5TnvQwC56bzcYUiWeP8w5xuJXJ
iNaDQgKPzEKks7QErirWcIXAnrd8ceLE9rUciTsl/r+bKb3+/ozo+C37PJWLmiLNCP4nHtaJVPRW
0gCedZMjCnJSTxrTndyxxSKb4gBZBS83opUrlK4/hM8Y46fun3TlSCW6CRbQQBJujQzZenhXjUQM
A+JmW30tu8MvUGRzzfbC+IfQNy0KwnHz8cF8CmbW1fAWcoM1BBAAB3QhRHKaQzNdqwzrAcFR4Gjq
Y/akeAODeMJV1Bd8DSvTdiJUy0WBI4HhYfDe7fdCAiaYZn6FdzCjK0B7+onrs4BNpdltR7hQtSYp
OP33899DXUdeDwzIOftRbKGbZ0ffW0ZqBEgBG4mcKGD+x/ncsVzeCaXbid3yqymtsMnHOonxetHN
6pMK1RjMByorYMrAXnsmQugwE5fp940DeyRR1+YpF2OYK/RcHCJIHB/oioP9rd79671ChpDPMq/J
MZNzSMOnvAis3atnBKSEfA/zg5z3v8hmMkvVeeBE/Gj4MS53tkotH3w9TZz3d0OqxzuXkJmCpQT2
QsbhtcHXlFV9+MEN/8tU1qYEjvchLBVAvaKMZ7gjlff+Cy76zb3yFrVwVC4j+/WqloGXme90kRys
0I+ck1Z2B46v99FhXS1iTkRrGFWMfL5737jZVegZsgAGJeEU2c9GDMv0WLm/kWhFwoHM2Dme8ZgY
UwMC2Lp0dgzstw7BlkLusyTlxRjAr3k+C3NCoN1z/MmwbAbV38kmkF8Ylt6TuuY533mw1+jUnsEy
c/5cNcppK738cq1cUoNJ8l0tNvtbxc8U0opDo2QQ82/cJfSkbxWkOXR452x2+2f2jyIw62xBFT0q
yaUO24kzE3F8y9mMB4FlhaTqcaq5j5D5hmMUnstK4JoTv/uPIHHk3CQaAc5rV9JipRrsMxvB4IZ+
HU9x85FUKWGtg3oPup2Det0RmVLy4vn35CnAhr4Zes11Ly4yOC7Hw3R4VDWANPPFSKIDXeMhBwnD
feCmZn1iCsXcpAKn0qwe856J53gQBbmvHBrvLQH4GbzwAiNIy5ZFAEsGlZwe3oEvgc5wwp1szC6u
GJlIBgEeOeVFGr96wic7qqvPnznWM7zsb2Z8FSi8O9gAee6XE3RB5pQU6Uko64MvsD6xHKgjefwH
JBwiqx4CVEYgoYhm+O+kWK+XseTXrClFzatwffafEPeYFZL6M8gq6zcTraUnu2Q2j98mvEiDavk2
hcs+tfStQdzxFonD9Hdw4w2tmyV2pSP3uvykVxwAVMhZ4grbgvKefdI2S1RjdsxwhKs61dYPsvCt
qal/qsSzo1Xuj/6oACH7+Ps6n4czmAmSV6upV2AVh2TL5utBZbmNbA4FGDaYpYK5XIo5YeL9A/em
ADqYLqSYGNgCd+uthvtPuO1zv0y+IX1QLSYs1DXEAOm786+e4RDGahxKAqydL5a41pkLUEDU5ORq
Y7tO9eryQOXo5yeJEzUYBuj1QE12B81pV3ZBDi2Zgnej82a4eKbRowpDrT4GBq6WZmMVo1lIsT+0
0Bo7DP1VKS2U9BO4m0MjUtLD2R8ko6YVXqtg6XK5UjSQ8CXVANkxQqPVDho+YG/dMDPIJyi1J/VC
r28wLGRme8HkuH9HP1u559uMccDTJjqvJOpot/d702OVf83iW1JLQtiLJAFvAgfP21RcoXOyr79i
8cNTjcaLl+yZirdNl0n0n+p0iLUGQ6T3wEJ7/aag2edMA58ddyFSxGH1D9fbCkL7wGY/aW+F/zl5
nGsUXy3ENa0ENxvXiJ/SvuYP3LbGzSGQth2ClPcBRVYjroXRDqyzaJr86hZhfCjPkziaRD2HWqjM
RY574BSBVbZGb39wlTRO1I/jJuWbo//5TWvIM4FyGQzmggVSGwSn7oTMJ7n0Ul6+DRvmu+VlAo7u
Q8ayFVD5EDaz5GIQAEpqVN/6UhvZ1I1nNQfQnJSPEv9y728lnR8bDT9EV02nSgxuYJGNEqHR50v0
Kx6NC6XU9PAe9ysYD/4XdiTkHJZVZvaFeMi6gQLreHe5xpDvqcDFDAHRq1HjjYnBJjJiUi3Uk44E
EePRQeT0utqhq2Z02D4vT5/HyOohRUaCOFQQYZnhliUSTZJcXyxAJqv8KdzzIsKfcsJSF6AAYgIV
EAIFHrjA73KRUKuhFlY70soGaOW+tSgKDVIffzZ/4+NZieQ+CnFPI+5c54AEV6SxB87ZqS0L3OUq
KhfuOx4v9yBWyfSrNYj940MNhNY5tqIGM4tp0NnsJd3yC4bBvjjdM75kowZHZnxr1Kj2ybMmcqLc
e/91dUn0ogG+SgoXTgZwqjF0i74tdVbQDJ8QrsjUPKAb9Q0Nlojor7tGfqfhazVxomhzJlhsyUS0
7XFjPSwuGZuT90QtPZIaimF8ZTtPBCRfci1/SFXe79xhjAUGvze3i53Nz+x3FlzYWsYrtv+oyzNg
QRU7fw35MelOnSF3QkShSEhC+67wmPL0uMGLXCmJLxXZijLw3V6f7T0oljEf86c4HzOoAsIaOAD3
s/6EwWYHz62VF2YmVc/O0KFicisZD279Jk/rkkJaXivUwIqtvoLD0rguFGgfnQ+VKTWS1ClQ2pWH
vu2cd2Y+RhvADpl5mZ9c5ZFln+AB5hhUR5MKaEnuOh7+s0c03new71djIrUK7UIUrjhdNHkpMObY
qfLAQKuQp6uTKnB4jx9mKEXNiXsGNS7rVx03jQ9aZiGpStMulh230ODgYwhcjmvxysll4mBS4r7S
gh2Po+3eOT0nAtQT9X3jF+GX+2t7TIpCYanr7/JMpsac65n9RrWv6Scew14m7LUeL0YpsWWRRAX4
NDcqBUIulJhXCVHaiIcGkTa0i3+EoHaFgWIxUyue1rQMG30/hUcgttK4sKZQRK3TR1AmvcsxcRSY
tY1HjooPbIBoQ25oGR4V6Uo5ErQuzeqGJYWvhmnSl2bbCEFLtb1KQbbR4eaMIfVB27YaRT3NYov6
FfJ28GF8/iNndIo/hcmF6E7DZI32KpesD2qOXdUUAyJoXeAkoMoItnPCmjK/toE+AirfnkyjgY9m
oROHQjMmQk4PROAWk01+k+YHNyF9K+dLYngmx3Fzo8vDFcHFI98sQPPqH/P/kD5GVBlV5dn6qL+i
sW8vrc6vxNDJts0XcYblodFWviXUJKQjO790FCKGXSSgWgWkwbEXyrI7ChAzAwiqPuVcHN3rDEOM
7r2gI1VSNoeLRzlLh/yAqe0YR6Elj58H7TbVh9l8o+qTCONd2CYYOaCg8mCX9f2FqxTZsBZ9VhXF
gepSDELdyfbOVZAEPZVRUAoICAPgSMOWneU/HJT0FS2NbHnJFcDN/TelHolLGHJPdrJWBKmlGouM
g0+e5NjTkHEUhidovm+imKz/cqbuRaA150Mobb0TEk2apHL+hVJuBLqO3sqh5tYFv+LBd3d/TlBz
ZrCUXX4rkmaM6fjwAUq+i0PRI+P92nNQciw9iguQhTyXaklsgF4Vtjmg1vj+RS1M97RWoissMucN
Wrr+YJbYFbbCvPHhnIv7DxKMgA1dXnR9EUXIjrs9zMX/WqCzJRThTO666Y2Gys2G270KV9VFcfnJ
nRYDeIF2b4PDAjIRd9tRIdx+wQ+JOqUP3a8YkXaDe+5oSmS5NWP8MSiMuHUkAp/4jgNubAp1Kos6
YRISCj5I8NbZkLPoCaeBbnNO0m+nTwMQM/IECP6qcGQsCO2LmpiLh2hsJLNzrLTduMi/lRYJxPnS
DCZ1IVztSK7UmnV6xZDl2lk0s9kk6ljuLqM4w5aU5URlaBkifoCbLYRBPY21OyG2jV44KHYBQy+J
EKRDG/9icJmmQ7h53UDGe+hV5UHTrZ6XH4W6LxDqTX5kAXkF1utgGGnFyY0oQRmHV1v7qYiYKQ9p
5SiA2HeQ2BpkP7C5quNwpV+ayPJnyVJIOZ/zrkC0S/6eELxmM5dJOzGwY/YkQz1yHJVdwoQbH3Aj
YNoDeIkXXe9+skhgiKcLEMImUb0CsVZG1UGh6OZO2nbnQEi3c1JsOFXbwFDf8Kz7XVKNnsGD0jFS
l/WeQ9CP0c60FTs6qxHYSKlUwbNa1JgZd/jI3+P/d9FV+TS1jnrvmnzVzXn23i7lg5eNYek3CVdt
8gG4YHCdzOzhV/GJGDsohbbMFY9I1tERvY03fgRs9E6L/mU2ePHHp/1iXla2Urdyo7lcf5muclGg
CY92TV8g2X9koRczbAAEW3OG6QqK333rpM+L03lGZeN4mI4Y7PlfgWQ3x2S0eg1S7SvmEusqtixN
bbb8q5WRPfacRMtp9Krpc4qKVN8dRy5DgTAQfxOek75EXM0EgN29j/gF+9coeOeIAxQ/JW6PhcqI
fgRBCdPkl/iZH7Bj0gKKM45tTWYthJO1kGRSpkqOYqnAJwWm0iQkW4uveHKB7gD3EyMuL5hlagwf
SNHIkbSX7okriaUN3yS+njdB4Q6H7EcqDPiO1pJEXM3lg5gJF9ApUddAEeursv6fNj3bAVKLGG9t
yovX6eYBPdTJQO43/JCVCu2FH83jEtC4He3teglCYSqa2Is9GdUvvBEuOM1t5O0AFJAtDKmgi1Py
s1nVFCxIvV5wPAz75xWRR0lNzY9eEGEl1C50fW1sIQZAwMNffTVrzV1DrUWY8JPVzwhYyqoVXntF
jHCSHJnNeyfzawciJ1TQK8McvkxSAkiY6F3ZXR7QIpSeIrZrKud34Rm1YxLsYOfmWFUcV0c6bCYs
AL6zWM4wWcEmBZzOSeUgsg19Ki0tyO81Iw4+H9zvye3CuvSqXeL1oibucaYA08l6dql7a3pSreiD
e2wqDB8zSAhqEK2RSz4bMaOWx5oEiV4XsXPmjGn2vBhTo9GBZx+WCnhM/R2FLAAsMRa+4TCjVdbg
zkDsexN8IPQxIHZjViPdnHhkmiaxallaSa4EuIQLw+aODkqRmDZK9BDylNtxHWyROeF1xpDW8a2f
CENPbQhwpx3Q6D6aIOnu8cUUNjv4KQrxmjxEzoSXlShRJPj2tipiJ+wY1FyUxy9WjZJ+ehplpXyk
gCIdctFac53ZdNQRA2lAeqfDYRRclE2W+8fVDdaJE+lu3xdueG/+HIUgVxzmIDha8++4tcsY5DXV
TN+HGThZs68xHFCn3Z3hZqZbB2WDt2pE6RECrglGlhNM8zy5YdpcaHC26SUw6cJ3HZlgVdcsJ48y
Ik59OOc5vPZQj9jnlQMBVrDNJOKq5yDsaReMaDqT+azEXCUBi6uc/jZLTH0z+W8CmCM/DQ78dvNp
uFkjMI9Pg2gcBVQ0Fg2z5ljiPESoMwCM0/wZifgeCWONMJkXKy3Zt4ikgnhKHTj+M5Z/20zeKcgJ
YK5S8g7bbKRd92G5vzlBB42/r/Y1gnQEmKsGpui/uXL051dSjWetIXvIAiKR4REEKLzz43lXtzDD
wrn3NqWgazEFsMoe1oTKm9P9CKo88dkGit1RSZFikBWPlbvzwTO0OSmAqdcR9ZPhmxjxdxgrxp4f
2RIeGla+287L3y6OOInV6IrsKN7G3wmshP9NJZ6KTAeq30JcSJxmt1opjF+ZJFjG0T8uPxx1rp2H
hNwlcGJQRvP6WIfFZ+THiLd3nAuvHN5w2a0pS7d6E9GuyGbmzl94tteW5mgM0D0xoaJX8Qho5b6p
boO8m4YmQSjLXIKEy42q6m9n3hmc6EyjjyE2Pm65VLQscGSNpHW6KnpRoFKKbeU0gVKvL85lKscz
XBzku89KKqpQd/OnJrCAjq1m8e9LaldtiHlfiE2m55gXCGeziBYxsIfQ/RPc0qhHkCTzgg61zaoY
Lw8FO/B2Ncryno04bG0AjA0a0/g98WVlR+VavQZDZSlQCXA2Z93kjdzI+CNomUUJfL6yXkGXP0Mp
kqjeLubwLD8PiofLw0Q0Wr2nK5Z4TN9dsndBGzjpIiSiN/5C1xW+ne3RkUi5KLLHMsnbbwbS26fH
U+sYrL4t8oZl6tQv9Z0Y59VAibNBgaMABdQq8D+nzD8KQsK00X+mAl9DtVXMxf4by6aa4RSm1frO
487PDE9C2taIjO9NuGfAQbqS58zMpNTmEfRnpvSfU1FperP7DQ1EdVFMbeg4UE2v14OUUeQet3Zs
O/UejPpzQCErVxCFv237ltA1Dl6DG1PboB9VGgF6oufrc0af8VpGf+6pHWm9Fk5PenA6eew7Yun2
2SOSFRXO8tfcHvQj8etWqRpIZxi228ZWDyszC390qkZ/W46Uc32prKtsAiHeHQRYnQEGDDeuy5Ik
kK2gHFZeHYD4Brpi7kLnpzpOLImtW7RLqs5iuYCoLkPQ7p+M+VPEPV/RczVk3ZQ4MqBMi9M78kUG
eZowxX9b8s8I04EEqMlfoL0pBSDSDulI7BF6tRZv/uusWoBUqnaclN3Dzit1O9gM0RQC2yAPDwln
pcZf0vfpNy3ibdWI9qfgW2YiLTj6H6f+aReVWokcoAQkIvqzSmjDoUISKjEDnvPvtJR3zq4B6P0w
aYrDp5NehnZPCrHWUEGCyRdChNq9bwT/YJQmAALsohQYVmkCTxlKTvkmRM0L0xEYfVA3AFmTUaM1
sSZ5Pg1EpCLrJruWJjBzDZ0N4VZKxUtAbPU9fkXeXOCRmAVX7c2YDK7OAnE8PsdXsvSNbljMw/cv
xDIm7RCJWwMP2oaYajfiuYqmeMgHlDnHnQDxo8S9cYgvpMbsuDUYC0JqVOy4XN6d6J19jMs08a5d
LClm4oJa0mltaqSjmqOujFJAl+ggMCGUTYVNVAntcQk042b5bBGsMlQyIox42UqyE3t6jWOdPEQI
yofiOtXjy98ENC5WCsieQbc5psaTPZbJC/LGF6F5+5LWaeFi5EqSwNwNa6RrN6YtW8CGGFD1c6dh
NycP7nUIpsKkI+kKE1Nhxk/tPwpv6ILWAtbIzF5yFwzIYvQZPwJV5rRUCAdmR845E4UcxFjBHKMj
ZORh28P4vDB7FrX19d/+1ZqpQxb8uqjSPBfCabzx/YASSfdg5cR5nbQBBGA5ewk1efGkAR0d/ubb
EscTuG7ArQAgfDH2QN9UxLQWXkrUwLEaNQ1XznHHHQ9syJGjUKA5cCCh/Jo8jTj/zYFx2ULIaVs4
LR7nVAze2mxRws/Q/WM1WzE3T5o6MTiXIzsD9IWM6D8kHaHPZ81n4qjH6v6oRSvjIWZ/VjmExjQW
9JS2+jWhDICmp/JqKerN35a5Dzd+7h1Z1vWjXjKHjn63Usx/uW49IHmkfZQ393MCoYIrIoEWzJDc
uZYdLTrpQRDREh+tFaIe4J1yEwemJKt8XWF2tX4uLQcUBrHR2XsgvABxW7QbMiMoyLp417UrK36m
p4RQhRjg4ViAGmJTJAuzskQEwldBIDn0B/SedKfHUc5PDySkYOZEY6Tqa01fnvgYGwDmLKGYYbvX
3n9D1UG/vVkh+91mr/LoM9Gla/OP8FjFVPQR3GXisDd3Z7/MgeDS+F3yO5AtnYYGt+1BlM55cs8i
SHm1osh78PooQ8dzLEy9mufD/73HfQwiotz9Soh1vlYNwiRs5T0bbnNuusmND++3oC5i5iQsUnaj
OxnrZGDy/CbZYBYVJeL2RlmBuAkA+76EwYCA1TIYgy3vbxZ0YDLmCyzBMciEsj80ybwAcTO/YuAN
ftisrbyOcN7qSUcTf4yS+mOb3vfI7792tsFMfW5nbvhluhk5ETQzXQPS/18gwwCRVnzeVbt2DFq4
4GakuhZdETYloNTv0P6/ytrrN0IdxEjy1vcoModMAm/ZxxPoCpxghIga+olmUHwi/KgZBSjcN821
uPl/bQ06MssAb8dvTGBxLQLLXOzFF3iApe6aodP41sVAva/z2QAc/pYraejDBaop/IBPEaszkXb7
Z+l0ej0APVsAoYAwPUFvyUVC19ChkReqwlied/D64su9mDr+InEk9ivKxeMi4h4g6OaP610ZO0jx
zBmeNKAbGsRHwqTtz0MxGuhDBTI8mWC3Sie7ERRbnOq8dXR51gh2biPzMO7z6ozeY4Fn7G5RfcDZ
tkOfdpXiwdGMEKek+H7UU1h9IC/mKxoVf7rH6hj+vvLKj+1jSoF1qG9H162qB6kukm5eUKn5Qkdt
oAuV5HVk0jN+bUYcBAp/9uSaC0f0UFWcAmTF6tkuCjWrhzE/8OTKg//Sc4YJDXO8wosKKMuQMyeL
dGgQ3gw4FSDI+5FtbFajNLGJfIEX3qJWk4wqrgfWuWaEPhM4iPlrp7onJKZGho4XmTdV72rd+k2n
QBcLt0OhmY/6/9KhNwRD2uHG0lyzlMScmdP9/+PxoNSz9mxiEKJEhJvc4NKyykC0kdiCTZ3JHpJn
T4YkoYt49lXmMVumPwwfiyZQr1J+8XsaZNJDD3rIb5bd73m3zBi/wiEH9ySFb+1wp00awyuaQTkq
FsJDriNF1gDNWD0ZNQnxFXK8VekUlwo2o81EcpC75DRfswctvGw/jP0QqWhXkmModS1HlpQWuUnx
1KZeVnRTbvjV9WuHRJp5ACJHoNIYWR+L9AKDN+qoc4qhA75jaWUBDZnVAw9wFH2xAgkj+EJYzHIy
1x4LePdlAC1l5h0RGvlMON4Q2oRS5lv7AEWgY2qkCZYdGRDBRQMv9N8JpLB0dscaUDSEjheCRlRh
/806qr9HcBF/bbskBuZOzin/f7QeULp06kcR7b4o56Irf+ySBNZrEQ3k76bXUiBuNuF8UEsrnnjr
Gk/JOrsAtvsDO0AGe6iERqbT1r6Hi2uhhpbNYY3Hf/S9WaKPY43iIIy2Fbg2MqgZNedJvD56L53/
/QsjkKmzeaBEPHTHrYDHg4mMzLFm6gv5UpDgsvuAGC4zxUFjAIwGwIGrnOnA5cbxCXZTdTm4R/+Z
5E4y/GyZg5G3TDW/4bfPCD83z6OgGICODaiVDosKBNkcHJACnhxvCUeM2FsobrHlL806EmGiCz6k
JhjZlfw5rXYIuSmrYoT/7+eIsQ3GSUCwhNiYJQuD9BQfRcWSz552zRF42+uGOJFpPNPnjXFs1Ncv
iVWDbg759TP/GRvz7VD+73fplnXbgqlR2m7Rqh/t9SK63uJlk5cWoisrJeosN6sX6Lja/EGUq/Qj
Kpk36u/qdeldlI0raTSplGzAjxEeLUoVKmktMnS0lATemmRA51G/0kYO4v7n0pQpBXn81YfeMkFU
E0JPzIVa6EtxUIYpEtOweHePIrzhO1z/gVt88Nxh1uwM3agM3NckBneyZYg6/t1kHBWNmBb1k77P
EaiUkxjn0LSt+bW+HSSV9+SWs2o6Z6C4uMZ58XgydLhBq6vC6qmZlWWooXNOp8jrfQsi/5wFd60O
0ovaf3Wp6ipn8BZsl/UWPS2FQJM35oTLSaPcDG+uX1JlnZBOEvzRwL+3OYE6lLHv1u6ghYJ6UCj+
Eu6pBWGZIEn3W868dFgSRvHAUkocyYV8QvKoGY58HuduHjN7zUnJcfhFpbs5vsGat4WOinVfChoC
gjqgWOHNVCYrTrvwVZr/O3Nv1SB/b2CHkpJ11kz6we/8pmC6JAkJ/wpJQCWdkkT4wTN+N5pTUX5u
CFKVqxQe2h/VJyB7/ZlBkn6KWnj4cHqh1JAA4bQPmc+ZxEQQBz7rRYqd/PqUh0pWWlo2bn8QupH3
LHM1tPEDn6Q+zetorYwQ8fjzR6MeMU+yH6EaABu6bI12Y0BP8OkQ0sqjty7M+MBFY31uVuCk+lKS
2Hj35b/YuUKTSAtAWXwE7H+HdZVzs8M84TG4vWave//OoMbglyfk0OyatikMrNq5STo6DLwe5Rrt
0k8Xut7RMwRtWCLTE08iQaNEl8T0qY+cXL/0+qyVDZx2xs2tQVkQyYStztFvoWlVR5FgtmJ7Smaw
z3o0EvQIuaY1cdPNImdj2tdQAmtT+Z+IFEoPQoqVnyECcyOT5GWEVoXc9wvBqWEQDtV/3re6s++p
HUNU+ejNaE2nqUSQyPtNuHlK4hFC3+7K/r7L63Q5+UA2FeAmKRT+RpN5v8tPEdDeUPnw6O39dWqV
/lxy7sOciNwxw3D/lZYYk2DeH81iTj7TLNu9+uBRG9ixcYFmCQtrVzpuXmoS8VifpW37r/hQgB4C
NIfsfIQZnpL2bsoUQyN1UMMbGbBJ84PLGWaW+rZD8yJQlem8pqtHBt58sZXgt5i5D6+2hCbj9WE7
v+aCxQZnWkDbQUizz9o5UVBuZkYMVHPpSstB8C5T05rBtdqfkhkT2asn4sFTIPT/xsLNYbg//6vD
RnPkf39/dHrv8KtggENKFaIQoikHp9wP8jjAq7Q/yrLJ0Ve2ZjI1yR0WTrcFqVlxoaKYWz4fFdzI
FAiooiBB7HEtjIKkvVEXey9Dulqx9mENsUv9Q4x0ahUfTl0z/5NkRjwGQhPoBgBkvmHg7YP6inRK
iL7McHtBmorNgudHFsqpdtGqn2a1TyvcbleCrFq8A6tUshB0ltux4GVBQZBjkTvedKm5sgkeNTJg
GmxLsiLHfbxXyQDUvAeElaRV6iBnIpZujPBZGhuSau9b1ATJSmuX0vOZ6x9p7RoGypoGV784bBUW
7etKvUlRyAMyL+VBizC6ikPJqxpnR3WsnD2ia4Wz0clAXUe+TAwb8hJrEBRsKnEeHbaXUuhpd7nf
Kh9kQRYzQWMLbxvQ32s743FNajbpW8E11Wj5N9qYl1H4sExuMuJwhDnWOREl6qRpTgCQJKaCtVcz
2dgmTiil/nc8citRgAHTTd1FIzMoLENU5z70WKc+yjBvhogpKK0bx3R57vkYSFm/LvdJf0vS2N+I
AVWTngkuGIJGWnOV4QUV54uydUykQH5yt0MsQeqY9e9JzknYf7bQGy3W49HYApybdjgCmYpr8/BL
IpQPkWz4BSvl6LZS/Y7vIxqelOjQwI/YvNUDhFASMSdC2lXh27f2zDIk/NjOdQqlm+SHVJbg6KML
GxNWpSB/P5RdwZStfYX3pRr/JpPEcp8I+RH0uabNwo2o29WHOMEK01uKUi/MPlpNlJIy3+unrSQR
ibQNzjcsqTnr1/tTNSHEkqNEursFpj1YuSiuYYCMj80+cU11heSH5OKEw+w4mgxg3G7SeeJtZiVc
VDTGRqMxU3bU8UWr1m85mSPOqgEwXbaka88oLjGFbRdLVKoUdRF/fjt4/Kq5f0dLGMbvi99tIXKp
ZwBCD8d5hW5y0YjbtPJP5Rb0AUSFWqDBfCngDA2ywzKBUwfG/8Cc6F7VcIDMTdjcg8EHHxcF2nss
pQIWfRVaiSRtcnetm9D+hLSn4lA+awABkdQ3Q92Uesg0nGmDAPY5oPYPYAYE8O8bzHF5vwT0yJdv
liRyXaiLzSsSU9EDnH9NWWrAIEZIz3J/3GurvUecN+F4rpUXAm3vJNU7FBQCB+44U3vAoQqw0+pn
Wfd4JqeKeyipNS3qGezkWzOYZMOQ07BgoCYKV3v6aPG0a6w7SD5kb10Z8sFy5pFkfpeuKYMKpaM2
BeAgloaWdZ1CK7aEtrGSBrIB0tBwPvMamVPFrMMXRoK0shG+P0NhTVRtG0pleQgDCxnUba+VFgt0
4fnP722BP7maOftwmbRhcyo5oPpIFdUOedBqlLPadsR/UuHJ4i2C9XtFZcJoz6BS34z4+CRvxMks
ilm1ay6lONMu+z6yL37ciJsjVAuTc+lq13vJrxBBLT9Ccnw1q2BO8VzKYmGZ4UaWJjO92K1/VFPN
vY67UOk1XLLHwOBqR9iNuKnbp0r22HjFeHuBeTeea/rmofW68BvYpq+eT3z7Baz4QPEbhKOPpazt
5xXHMUF53byZ8Qet2UY6DQOIR0PL6mhuDFmPcLpSzKDqB7t3201aIo1hHxPwB2DC8hlaKvD+KcFB
9upc37bSnI2PHsEmeyY7SsGFaVIVV7G6hAKmwnc2i+abqTX1uA5eLoLi/vkXdVgquC7y/llraJHk
kCUJ1JCQAs+IZg/D+e3cS4GnieiofF/vnVq29rCQ2TWdh/Epv22QEMD6TcP3B79EFOCpF7Xq3qsA
CRcViulkDSAJNhA3qVPzFFH/XbW+DSTWRzldNYAhKLsErBoFmharT3H9OaI8Jv927MdWRrgJyVFF
y8xqAQgr2d18XfHKNxRpp1Y3+IAke8HW9w0bnapFQpBguk2Hj7pXV4ABlutpu1EhtpP8o0mDnIeD
bYzeOknMozOmgX7vpl5EOJTKF2DTcun0vx9TPOeLaRLMEno6Wx4pCgGBxYj1joyvRJ5jVz2AiGbf
e/AW0n940ijjruEhveALOPZlAHGTujgXaknksnr476sjTw4E6dXMpQXo2KAUX5Fnv4IYPqreG5uY
brOybcYd87g4KUW1Zrl48XkJWUuXhnbYfdAJuFyNtLim8HtEu57S5m1OnGTsQa+Sxfbi+26q9mGT
eHLfw90XVl7eAU1NeaCiad0oqgjfTHBNYLYu2nOHaiQRB17xDMagsWAW+znYXHl6+2H+lS3E8NcD
EtK1xxg8E7bcuIxSR2CwkueIZqJ99K7jlKihVzxNOHh0JQzNLO6CYCUzPvZXosMuoOuxaMroo/Xu
7CgLiUxWc1iD47bfMWDo5Zk2Os/SJMlViLymKlrQu+LyRivaQM+fi6Exq8HD1y+BKgUCBBAE9tnC
e+ZNAp1BJ7lwrIfGT9Epa3qzHkb2ZQM3ljS7H+SXal+CFyYV8QiN2tPk0hNTf5LMWOvxxikHtChO
67nzCDB1yzwKFIz1PKLjgkFoIowl8Kx6BOkOeNfdwR+IKelPnNOxdHlo4ElxGFhbOBpsCqhXXK2K
3/UC8Gc+m8EXpvASgSFjMEnWaYAXQC0sDXl8z36tUyexMmbMcdkg7kJyk3UAbbYZ+lcJdfhVRLP7
IU99qG6J3KKBI92CbSI+CtwzTfEE+qE4NmIqVRKW95d1VqP1tMQby8Kkd1b+KSYRc2ATxLC1ywYk
wVKQa1K+9iRORXksekGbjTyQPJQc1nlrI3wDUR2hR4B/LxKPXvKqCQXe+LZt18/Bm5f0GvbfQaOG
ebWqKv2vjTFVPq9GIW/sZGQiaDUI4jxohCHgqZIRZbiiP8yla9JwRdB6UC457mPqn1HGbZOyZ+EX
hTLYSu7IV+0VE9pFsupyNuURwDQ88k1i/ytQFJAubxwqc0pW0FCslY7NJE6jjDcDCs/S/w7gjr4K
H8yKp/jNyNyyaMEgrtBWcYMMzsQ3hna8C5i8Q3dqjfhKXpPK0zPkR5uPXiHeJedAIaepHi5qH4rn
B8Tbvyc/1+9gcyDG+bHOZ73Z9Omt4TX7IdhvqiCIfQMjn/JFgOD0rrSQ+vdq6PvJnxtgWIBASDL9
j8J1eOnWl09C7LchPZdYYWRnVQRSG+70j4Xb4w+/TIb48ry3utg0D1srnuozriIOftcdkVyMFK0S
huVNj4II6J72is8ZIGGlbXgnP48oOuC1cWknfjgl3MxZpZ/OMKpJsyvB1RXlv7YXS5oqW7ZwVpw8
mE0gvK7Lq0Qjt6aldjuCXAVfhrbqmNnhR5O2QeOfRhSfQez6pt6ipEK1DoxTYMVXJaBdMxSqNGmn
ieALFvEF8ADQkwg7ZjZAsRZpwVsEE76Me9S2cHRpYgrMCF8iAMrtMTLv/Mj0a+UH5ZZb1bllnI8p
F3IxxjaLgRkp7omUJYr/Ds++8VgGlXUms0gZVi6oxcZ4T1u6o5w0D9hau9w6yP8VtP5fLe2Sqdc0
E5vHPEyAWW+trvUow2LYT11XhodMZTgkdwZKRNGaVil8acJ6gVmMUpUh2KNeD9HjXXcH4Nd5BUmh
da6j6wGLE7Djo8bECHJusi6Ep0+/owzpZ8CTNqGH1m3S3krj0+jz3QGRdtQaOAwiFJpSznDs3YIE
tvNgB0pxqLJMy3rdv9b3dirGFnwFzrw9ZxGb0WsjyOnDuZNkWTlUPJc6iIuAz3F24hDjr9j/kx/6
5aoJoZHYdb0lXemHwmj9lB8Vjr4Os39oTIM9uuWvxKL+dbd7hIV2H+G7U9G5Ck8acxNPLE8V6oEK
VmFlEbYAHuWsqk4iJKmiqFTsJScRHtRyinZ7zTQKU75ZH2hJxQ4dhgyvaut2JBZPQ1J4FCwqAV3W
HQCEb6XDSJKHGJnD0pi0DJGNsAhbDMzPHyZHONuRL8fWPYZfmxS6g8Hm82b0osrq2V6GXafYnihX
RBOQ/W0eXxpNV7mx+PxYUNey8r8lMUnYRsWOD5+XVaZXpFGn+8rhWZWLuFy0qUxALw57/cVWCxw/
i/0A7MMWOcvWB1g5hHrikE7OgM4CzmGPoATo8pY9/KNQQly5AkyN9bKll1rZ/0q0prgxdsja/mWy
o/rMZVpUhaEdv3HTp4/VMFxjLRE7LCDjXPko8EL7KZNFQj28BqIoWkL56DnkGYEn7NiiiAjB2ESt
rpjVxXqp6tWn7szWpY8ze8ym23D8reR+6UbLMQdTYleNweJBYK02WIheQcw03gCBzlt0tkRSNMyw
WWuYjA2fxJMgUMGLkIDan0WVYdA6Z8pNFB/e2Ep0HuMsMNzouZB+diuuNLTyyDBR3fUuW9dl9Xeb
+6QiRBoyv4K+yTIaeXyHmSBho7lo6MLmqHb9VCI3vwndugwj4BW/YnVYDHdt4L9A80X10NTGe8Vv
o767uN7zhZS8YVRQ+3I80eTdNlPiWDjpCYSN0AdFLWUT99nd4KGyUQ+wZh2S/ZJD9+k0vLJzSaIP
ni/qBvGOPkt5eJXcNgGgzfunCvpGZmytM64ebdn+0POOC4EGdofPPB/ZVNQJUuuHKe/YQ/hGObfb
lECrQBUpG+h3jJoxr7grjsVssbONyaTefpgirJRAyP0AgcrEj9XvXIDp68dRN9dqH2hJCVF7iR2N
3lQRspyxXAv6fk6vwQ0HYKnpRmEamHLYDJwb253Mm0ph//Eujc4qsE4yL82TVPyrigp0F6AYnYOu
v+U4EZ8gSB2QsSUc6ytJbueuP4vyEGVVVJG9zPYtFr/i2hqqblHLWII3Pn1hWJBa5/jxGUSS683C
H9aS0e+WwF0c/KGNbKxOt+T/vnnumdbik3X8bvjyfrDzFZbt20Y+4QGySn347/6m1PyzGEiZUnv6
EVTy8WYET7yvJ+qsERpEBvyDYGM9Z7cCtc7yRJfsQQMnO4yP5njfdaqIbTNSVUJCO288njzWv1Jh
C2GfooBJWd5SI4cxG7njAcqsZ/BwJHcdUzXvx9gjp2pqE6FDot+uKL/LMBtZmh060bKKk9s3j8US
0tLBidQHIVphcOEY4noeQpkQW3l7nNLalFE7Y/nF0pyuxywPwsS4QtU+CwbnNcpb0izc1iU0QeYZ
vjzz/idVGKHVbnGyrFyDzBht2QEmcX0zyeaNrvExww+AVAlOYbJVCXNBY6JwxnUdU76hYCxcGfT8
O5sJWkKzxms2btiCylpcaVlEN0hkBOFdfLmeVS6Uyjg7t43hZgNEG1BH9p7y8q27PJGgqu4gTIsF
eOh3N1CIb/tbBpjcElV0N89/CjcUwfH2Ltf6yTCME6FReNDxADW6rN1Sd1q0IHYcTrD77ZcDKMKl
7GndQppP5UY8ebEuJcaYuyDiVlonBBLzh/DKLwcyHqK9haMFlPPzZh/1sSRMciyiDD885Lbniuxi
EbakhBUs+Bvh+wZyEcsaCy3CK+LCGkd5bNA1RQBH4jGdnxuDWASkeDeeWU6HKLbd0HxvQ09MjYh0
5bnYhfEBeSadspfT0Pc+aYMa6h2jMgfjyjfGpQIGJM8o8MmKQKboRRi4NtPwen/ykEKMVoxk1Ydj
GTgCCAm4PO+1Rsixmxe8MVEYGnL/ZdfoqpGPUtx8X6QxBQgPDPXHfOnLlpUmrq7lOuR4MvoJAz31
EkmLIHSBHOqhGsW3gOZ40r0NAqfoaCNGJuZRNQiT1hmGlw2qrHXUkFRDrlFO7mhepJzO1svsvRS+
ajgHeT/SZ8nn//rsSH1/TxzqMbMCuTWWoeiiPqJ6KxjT7T+eahMo3f9CQ0LWADRwouDAS/M3W54r
IWmRhBfsVdR9N1fGw+l8MBfjOh99NoxyR8eUbOXF1hozZbaokMHVgj4KKgmofpJ4jRhjWOzrSek6
zIOoOcBbewY5feCrcMf381uGRYWms64cxPTSOPT8xrcTTvy0U8HaDQ7c1Ii2EIuEdGUd9C/RzOd+
xZJXRJOLxyS9V3vJZun5rx+TVcpjRjCRicgPpQeoQe0mYv5sbS1LCM9ed5wiWREXqM76C3L3iNko
ird/5Cp0nADGvB4YNbkRmpU2RweweaFVJrfC/v38pMbolEDWZFaRWIq1M7HqO1WH9iPAPFJYjkvF
+2lJHY/nOlvwWc8qPlMQd2POUCcz4rygq7N/d84l+hUqCX3kEiTHjhefpeEJlncwszFIBpP/prH1
BwNFTGnXGVDWNMisg12f+xyrKNAH2p5H0j9EwdFNBFJDpkA9mjKZJm2befsEaV9ciiEAc7Wqg/d1
jROfQ+/J6MwlFrnPd/TncHq9Ct78CRd809VgRtLjMpr9rkKngR2tN5oyaRUT4N7VjBUv55smbWNL
SlugyuZ16+lkovYEM2xLKDoV31GAQdlciRt8yG+vQynxBRcRDhVP5/MwSGXOer81v5ghwMefZiyO
qpLwwzpjiC12kqwBQaa4C432o5SC9ZZ5vrb88l9BCcmTXRJPVes2sNe14ARbry9fE2iVpJbPtI7d
wnZ5MU13d+43vdiEAv+bRoo/JfN7KNqlQyOMrUS5BR0VKsp3O4SHfPVsP3WWQjvndn3XTdH9swBn
QMr+uhLz4i4aLc5i4Gn26Aw360Cvndw0V1r20n7f5SNLmOi6qXrlVMMKP3yFhw/CW2IKZexM16ko
S95AhrSUxVxHLpeHXHHApZf8YfZ8FrliBQlgkx3LHTNu2UtHMndlTwZCwuZrYTu9ZTjFUgNx/hVO
ZQygSgDH7NwNfp599WJCReVSE3YhwhnNG49ze+cVcEhRBkJewdW4B5mp7S6vCnxXdzE5KxG8BQOU
aCw9WznUugXlPCh1UuMvhpauj9AFa3qplLOMprhQQe4X2cCaoci/qrVGLT20/ka03LANEPfgRRRA
1XD6OLHCTrVkeX4ZDKhdws/lMy+lj7Y9ZlgumRDFLsSt7CrK2qZsoPm86jCPTBg3o8q06mKdOrMC
/nLkTsAisox9LiqtK+Xv2s9oxjWOV4WTTnBFDJXnkpiDSu4emgWMrN+n8AwSOtkc2OTo1bxNypza
I3UBG69lj7Lc1GEZQzeCR3EeSpY6L7+YCiSoK5vP6lOmlA5VLstcTBHjLKVC67d1IhTkxtEjH8qV
p4ML6WL7tMJMUjEpS/q22CqipEH/xOPhwjeXzdBbnw/NsN+Bxi0+NtePLgaFrZxsknemXIUKF/Pd
K9XUvGbSnllg8na8ZyatVvY1CYgBssiGnVJPNIqEmEQve2q4+VVTpNMFzehZ0XZ6TnU+UK8q9plO
uVTdP8MlgtO2bPfsHCHfg5nMxyX05sp0BEeYfSDmm2Nkf0cPXQH/dlIxFIJrPbHysNQp51wefhzB
LjAJlQwm33GwpyCx2gtYUF2Y9PpiZPW7U2ryvG6Dm8hTdG4RmzL+GR+lGRRQPJ1Z8jUyoBj584JW
rVfsXgejocttfVyINJJJq3BDSX76+gk5RiEwAWQ2eFCShIgvXowT90Xon3HsgcCiJYSaRYDC1bRi
hwXyDC0Gt091tPFlBVXBPQxCyVKylR2O1pPM3RST6T6hwsoz/ua1CvmuuXwfoDaRe+QfsAD5hkdm
Y6bWxJBYg5c7KemCEpic/Gvy+gIlUPLOvkvNADr82hj+cRdRE5ZzGTbBZUiOW9H2dHL6j9XVTjnV
JXAri+0VUIWRoezQ0ACK6yweFQQelB8fgND897e5ZTRbf366UGm4An/g/cI2WNqNEMxqBOmgiAvq
RC5rJZ1Y4ZIDcl16SikEoqR7T1EJScQmERZOdx5g6VjAA5lgWt68629eYL11Bld5mUQipucBFKFK
eZypd+sQxlO7SZ8DaWMfbJjwDbC8PYfb7AB+yy7LkFpHLgUegyXSYFRAEtrasPwEAmoESaLwkpbn
DUePAzrS7EHe2a00cTKUgecUciL28IijeIFZ1y0Ti329yvG5QN+w6L0xwrgt8SWjDopzvPb2xT7a
AhGIULNWYQGPD7ndzEUdGxhvxoTpqY02fpHTscIS05MeP+EGAGD+EoHcXSr5geozUHSA7BEpKZNk
C8aTCebJjW2OvKnQ+lpSTmqLPW9Z9vtzdAvN9u4F7eiB73U7dJKusSCE3gtTkC0/MlZAWE4TTTGZ
DVdN5iHusZDgYmllq5RlrAqddOsmkigYNmwNa+Z40adHByx6ieZEKu7+Md37YujpwRgkJTA7+vTk
t4BE1Y/Kn+4lYsn38de57DRjV1aXfDN+BTYehiCNEjWCUOEwZEX3ZB3O25r7/OopANrD8c40Rh+x
RH9Gv3X0o/aGjMJZso4QxwYxSDW8UoJDCeZrwNpcv1BILNnjwlinDmXRMQxZJUiOTSmui7Sm5bfT
Yp6bZdhzG8zEQlX5pRafeknk+EnxTS/S8QP4PBE3Ib+4B7v9vm+n/P2SozunMv/NrD5ZPgY3AuK1
HJ1QvwYLwDs4Hws6XnDk5GJwdGs8slqPRQILfPE4HGylvM5wSgAvZjmCYp5j97K8fiQmgg+img7l
T33zh1mF7ygkKAaKkrspa9bPLCoOX7EkCp+zFC/oACTEehNWc6IWqTMge3qpRUuV28zppf8KF/bA
i7Eg/MaxOIAXdmr9htYVCgpYMT1Z3rxTbs+Wj4qCC1oF5UYUTScrxnKpoTqf0c+MC7XwSaLuS7NK
kYaOkI4uQF2bXp4hQgsjKv9tbhZuHVZWfg1eneUd5QpIoDfQIWk1QzezNfSRROYF7p9DP9/kwcGd
FuhFzIVbuHmEuhoeFU8H+5QougMZia6Ht+PoREsZhOR3nWgX/tYSAbIPC6XZQnMPa7uc3TY8ZWwK
ucDzk4FVbNY8IvGcwjFPEoDSo2XrpDICCBMu6EmzKWFsWPim74ps5P8SnsCX40Vv67ZRGtjNJ7x+
THc/fy7Yw9bS37nuTJd2U6J51yKMbYiTaVE9sLCbrSjJRKQ2jDVOSp1aiGMueYk7VHHtsjOI/V7N
FFS41OF+Nkucysu01L6h99upZxEemNZDwnUxAHj8/XCDuioBjB5ZTROKMkg5OFP+4nBgq94h+so7
dt8NNvOq+ZxCti/cqjmj9Acxt8Y0WczHW2JPBCZ8F+sSxhWgFTsGJvBqeqRWeXAa24AyROxyg8UH
m5n1oKuROMZQoZx7Sec1XoX50n/gMgyfC5hqPALTxoRJDUiWKb2bd9lfM124GB10u6wEo1FYYmKF
1+MKpCeoiGQs0s9P8VQQkto2JwxCsX1yUFHNOVzycTpenN8AYvzxQXl6cs/OodX9UdTuLvnM08hl
yXsOqmSSTAmn8AJivVnqnuXh5lJQg6EyE2uKXSYTiieYMT6ZM1Qyxe/IooQoFoSRvN1Oy8RKoQNp
Zesqd6UM3YojB6+b0PlZWTjnJOdlGbzr1kFksL+teID2wPiehgn4NqSw1LMzSZ2FkD+omqoSQm0I
6TmV7ke0JsxC+1CJN/nG6rAU2Cl4NdIGsb+PxGpPtoWbEjrnX8edGFwu6oKNhuESoF3cES0lYnDz
bV+NDW9r1N/tQq5g/WGy0/WxNHYzOG5gUXUDmgeDeXeoBl1d2hcVjOGD/+ClNlJXv9T6IVHLwoCA
cg0qGKuHtu0SkV9NaNwUdtYPlcRi2Lt6HKfoOmr0x5FSQf/NBCRMeZBnc1ES1xBDI38MhK93rRdS
QvCj367kpfFw1ZI+H5zM0xmNJSL3r5ktCCEYU2hqPJcOMUuFhWihPTULAmITPxlOg1Rx1uwquypR
p6IvmktHA4lmejXbo4G5vJu6huTURtuUVcfY4VZCIFTdwBFk7y/PXzeu75fPkkQsPMBqj8XfNiiS
dYbpl0C8g61wxqvs9THXXGNXMXNEvwXB/6y0TOO7cVSz8zDe4DgvCOCbSMrXMX5O3pr+N6jTTS8Z
VINJ3QLATToxwDbRkaXXVuSSdT1L1hQbN+a5ApmllBzgWu5dAdKCmsQCZdUtsQYevTQx4gFgrtLL
4H5uhWoDwq4foytMeAek53ov0zhfoLSBagoHgUJwmxzj/tAJTq16jF00TnHRK9x32NsVhpcRKUXS
nptena1DxE7+AYRRmFNMpuQHKtJc5ewB9mXb+O6e5JvLuyd+8/BLmCUfvjLQs21O5u39UFE8KpZt
6cdot6441tjy9doXEgWM+gScRhyBjhzSnEe6fO0zyxHn1b9KxX+GJsK7aUeWj2AQgTsO8o99/XVs
tskq2hZeyEb2c3hoPxzR/bG9Hyq5aT2J+bVX8958iZ0N1Bv+Z6I2aKtafPQvp/X4VK4RTMX+KMw+
rpKu1yUGYVj0ptywIyTMrHrpbibogyLWVY5OxDtMtR/TT4O/0hnA5FCFK0p0Adovh47+JhrP29YL
jPVU2K3wiA8OQyIXDUkLqwZ6D6VZySJ9FtdhQ/eW74857vQRxijeTI84o0TgOuZhtsmv4sd/UE5z
/OrS4kuDiL5nd+tdZti0KL6QI3FmP5fIEvpk5ksvYdUao3fEu5Vg7u7/YPR8C4ehnyNey+K0gczb
Wiy+N52i6r8HC+/3KqzbmRxYo6Yu5czYXjcGl54VS3bXQkHg6xOaDZ1bQdeYUgOX+5kR9pLAgztH
WkOjcpmCmJGG7p1XD80GWAnoNBYUCUy1zlehgSNCoGKxd4HiAyVxqpvaN6yRTMSUFPAmvoM9OfA4
RxEMu40VhAGaFfHcM+yd5/HScD/SmbcQfouplXXyGhypwgEC3WaFg/8v1tWT/Ni9Wj9jmxt1u01E
z17uUTPcJOBwSj0YcuqIAu01B22MDy/ExRRRN8ta06nwqSDdZj2dvVSSynwfu3/LiJdbwx+ewPEp
UKCnRjkbUwkTpNjZonN80fzP2Qbl4KEg1thg0AlJFJII6cA3BkrOc6Ofd5JQD33pi4WFnMi0nRaG
Tr54aqXH2R95kBvQCU4rA77cLALes0EwKhYgLcOAuSAuvzkjiszkiXhpakruMjs40Q4gTgF8VVBS
H2iyKLU/2+S5iJCiYb9A67MJ/Zvx5aqXG5SGjeDF6nS0k3IwqPynV2yErHw/rxxwQY3jU1yVwYvc
n+JAFsKokbqzhubvmtneFI3fTSKENKi/OQVYBHUKw8UJV+3gx4nVEXsISi64VSaWeh7JVSE7OPlU
XcOImoN6Wmx3giDID/VCRuo1a34PnM36GnVogKNv5F4L5k6NScPCc0odfoiB/qkoea5/AUf86iav
ldjQAjiz0afX/4YEal/ayxycAEpJtTAxSs4w4HZxSjvRgDAkpLA/Lkn3RDgSb3PD98afEoDd/DUM
aP7du648/5iaESfrA/d3NDjt3fhvdI+2/HMThJTi3GSaTbVMns1NP73d66x7e9horQU1vhN3CI5+
WInuVnomWclRkxji/sJoIlAKidjUUHMAZTxMOm0iDlEJgJoSHx5ejIheuk35UlRTzkxzTn2tj/b0
9ihtNbCYIT5Z2U5jVa28Ie05+BKe6cvkLyWkDEFXSbo4RfHbBthx0CVW0Y8l8qij1CphB6rJKztV
GW040C9/eFNfhbEBGatQEO/4V9vdo6NlXppV6zHxcCvO7Us5puRXBZUJVSzChsImBAkojXzou17n
ncdtG2e4rL1FrZlzm5vk8PxWhXBp5EfbxypccB1QZUwE9Hjy1v4ADilnHWcpkaNkPkfX54sHeTkz
DliF6zDCk+VGgj1DKIMsWNuYWT6RHryWv7PGyOjlucRzx+Rtyszqmu0VplbEn2pQC+DSobEmA4iH
tqNJtGZnIYHNAik50A6wsk+/mbWtLgrQf/dSe2SNcQfiwYZUzU6AuOpN11GpRPqtw/PdTxVKJpxb
TZcuhNKURETpdqw3viqbVz8tG7bGmYsmKSXuTfPQ2VGO4Ka0nSCt5lgsagSEH5f25ZFLcr/W7wjT
JlDUc3eCpDfJFSmXQHGJKa33qzEEJyIemFsWSeGz4XwJKBWzRr5ojYMxNaZrUbOlB03Y4o0cvXs2
/9ihiEER8rBdLooBPBwjZuCkHSBRcQqnh+4bxc6rrFvuxjAPJ5y2whQMuvIRMSP0b3TJpLxOSxms
ZrkPL/j42MR6vvgYxcI1/qkYH3l6Wa6m9uxNe3B1eG3R4x+s7VIPWdePsqco5+jjVI24VlTBHupa
q2Y03Vw/5mRAllTK4t4JkwPey/2oXAnidaT6PEOeysvdDJJoMrOkp1itrki7VcyQ9bEdOTXCkWbC
CEKZ5uShpObB6vFulMmXdErcQd+7aOPA0Iqo5VdLxeM1NAUHvhibGC/obyozShp9U0vJOiM/lvxA
Q7K3md/yNvqki7dAlOXwAgx4G//i8XrMGi4R3cHA0jbX4z9iL1yhJWBV7ZSK6poi6t+Q0OjnCuji
MVVgTbDem9yOnJ4/zil16DDZRzTfQulB2QRPmInOclU3AGXVW2YV6PNYk9AvXQetjmbZhRVJjyal
p6/ls+ewgmEpOEo7xNqYnVj4yWta7fePwl/bWkQzhXx7WNLP20G9wBaivC7h5mgP812K5rW8j1a6
tijr3g6r0jsEmcl5zY1Uv7Se7pWqjQc/9OvuNu4rcCqyymvyup17H5f6wUA+xHRCrZsh7lNGxQ38
5TS6wQ8YkBO+wilnARL/9o882M9VwhxwiyJ6+SQ5Cqtg2XdhasfaNl3eKxpiH6JFgHE9fs7g8AG0
5/zxipayBKwrMfYLw8eq2AE33rE3IiKBmxGMDqA9mhtarkLiNNaBrKHWj/waGWsjJ4HR2E3JFz8F
aeawEXpHgEmUQDwxOwhpwpaHu7vOjDBBTzAUGeNuLRgP6+wFRB5Ih75UYYC6QXdHGntOPc42mWaU
QWOooqCOT6L0CCROEeQ8fyRmCwWHGG56AvhS0WUqwY4nYX3IphnwGrRolEOu7/nHPqgsn67EZ4Zi
KyCEpDNN1SYkVm4+nv8fcnb1hOC0VJMR5xWjOHDYt+PSx+/eBtOHxRddRyLh0rbVmmPOdp+RUqUb
uQbpJkPpwEEdHF7xmrKPK4c9rtCAUYbfKcoOGMD0eE31dxfBJ7Vn2eHGJo2pzMLakyVxaPxeUsFP
fM5iMhCJfXDboy0Do0WBRWGN2aFjLfSf6lEI5o+1C/T95mYQd+tkAREJH+SNIxfPdS/4nnR/2sm5
uQxQw3sjo2Qd6dBrJ/qrv6U8Ap+tf5yQYokY006zE5mkwnUiT/8qqja+bsuAhVXzjxhKqYViELGl
scURyLIN1w8HSL+s0+dNuutx7ATE2WLvpmmzqFs8WL2WNEzjjJhjH7+ob2QCqIvA4ANCrwbDHH7d
VL2qxW71CcDUm9CADNxu+UrcNMZ3yo9ZFuL29lMjh1suPI1RayCBdFibmVC+yOMGgQb86ehO75WF
bGWr2Z5zSKJxNSwO70V4IsPfQI+4/02cKolVMpKWGDAAu9QhxgAnujYXVf+y0UTvYn0qzyd5RgG5
pYYTmgQZz6HSDDoyt3oWw/T/ofsUoxQFyAx/QXBAXN8bCvLoptib9AmS25px0BuKAFsaEO1iCMdM
/s5YTl7yhE343+3d9Jqewb5cABvwZgRAUFM17Vh+9U9EJi35N8EIMB3YfHNzqSmYeqQGxEhJawMX
14s/i8ljU+Qo5fhjmj/ltoNfB1cEWsdzFoFr5O++wRqmDuG3pVazLYTvuMGPk7wl1i4m/68eSeSz
MhmqM8kFWJ0Oe6emnfeFygpitLNKqVnI0jVfF4rL5CFznxYoE4KQIsMiN3X0t65ridcAhsUp25jK
k6dGfDqj4uBm3WTmY81ZdvDMklxruUolAqVT//9zdDU56+xWIlIAR6zUAaT6a0GBrqFVwf9eGOOi
WamivkcMbohb2D7fXbqExfKcq1F5+T50B0Dii0S5BMkuJ9iDUYHW1dwUruhF6ZCiZe9XQ7zyxwwD
D6Htv2oG4H1gsY9s0CeV+LKPpa9JGZN7foce6mbQxgn3l8b/B789dNTKHPZ90CxoeXtNECD3nz1w
pxJ5ASigYMnTXP5ZpymJfuIA7mVn//a+VhUBcdHxOPKftoq0dlIwHAjiEgMqaSKY2G+elgahC180
D1rNsY5IPr8mjWPLDlz7TzhsQRvmDk/irNlbleqgvXad+X12hCNS9ubv6zLccfuMtRcpazNywCNG
foSzp3jCLXCFHvDgtL8On3vhDb7BH7Hk284wYq4IezVeOI/S5x2B5WJUpRU0QvNilPvbceNkrYed
OlddfjKOJwAuVyK2oqwLpwpPTYA/8HnIWGD5xH3p9BwylJX5K/4gPcdlz2swtkFXILkkd1979OWf
GZIqRtC8qJ32c03I26TA3n0DNml/v+WsDLP2rr10Xc9OGLgTs1W9wj0OuVW5sjK6vlk8Te/lWE9y
Lvrq5QrngPS0iD7Nv39wBwYHU7ebvptc5uMRz7wBt8muRFv7tgnB8qRlccwAX97rpy5mjLw/TYtx
pLQREnoGc23oghEI5JVSGTttuJYo4xSe0ANayOg47yjRYuDWCaG0poenucyzv3bL9COhUFj/c8ov
8Jb5YYcAjFsCcQOJDBsFijgrDimkLNymzRaIRxNASgIE9vHVLgn019DKUKxuwGWq9Pq3bgvw5xUl
Tiw0rU+uemzjuIZahShCa9ElZ6zNWi+oYq6SWR5zJcfn8eoRbJE3rkiDzoU3s3oLNKGbOQfk3dvs
unkVCl2OjH396jktfzo+Oa4ZAb9LNUAYLSg2xsAJWX2u0JSdRzZWcoKPTTkFdgKaVCO+RgkviQVu
cPAg/rv8iRNmOB6RGCXXEDmmgcvlLXup9yIttdeevei33gSUyWUbuRbQBYN2aBaOwAIC/lwnQfTV
x1P79qzYgHhvtUVjiydepGPdu56xyCO2KEqpBapTP+PaV0+anyYNtmSTAUU2AU1uGPQcWDuUS/F3
iO9Db0yzupPzcJpro+4N5pQpUPIR/0d3iNSlmHpI8FZbDO+ZIoHtB1sxBqBOpgfPS2YyWHp2uA9d
NrXmyQKKY3eIyIcxWU3zt0ylbiWJzILUXbHoaIOY8BZZWcGFfqh844oPfYkK3RFM6tZydDqXZBvL
blRIt1XB5+H1Dnzg0ngS/xoebdjPwcu0WepTdkkrawG4KAnK3b8nw6JOYNKPHbPEzqdA/P8LElrg
rKO3ML4a34gjTbpRbIjf5tO/0O6akKKk339fM8JFfpawGAtImg/tTCtzmUoTUmUZQRdupzUycgLz
exkBFuEoAfsxqGh4eDRNGbsKeyqrUNeV8tEvZOH4BcwGPytXg9ChjDmvCfXXT8dTAzCpcYIWR26M
YWus/js6268nN2TfppmyT0NOUBL4WS+5aOA7s1XnjEv2e9An9XVH+OL9/PWaBBDIQomRXHuHkCmf
7Xy0LcbkarJz7qxLqtuKSqJQqU9KweaWsPVk5nKRaWZKfEHxQTq/ylbdPSGOSeqvSmFja6e4m9H6
2TgV/o+CG5/hvf1YgFqbE+cDsZZ2umN+A+zl2NMXBYTjQMWFyYJ2RMDa/HAYDJqVyPuTwbAq+hYG
ySmqO7EpUEPrHYOWmmNEwmFdpeloBcOiKb2dGhVxqxo3cfAXfMlIAkAU7V1WG/uCmBizJTgm6JIQ
cmVx3g/QjuWvxA8ILu1AIXJMxy3DEKZK5XLZUvHUoMAO6oDJvyMedIvBr/tTTGla5fCMgG/Vg4TA
HHvKB88VVPWX/58BAwwCi0R3+Ffb7CeAWYAIiKeEDgqCtVwN7qqrfLVBDNGoShYf3ozzLBo0WSEY
C+xD2HGfKUGSfw+uFY15pu6aGsIVOVmWnoZ3xmxnNs/eLaMYrnvjc7ev2GfRmcwhFaQTV0lFRCLv
JelTrENRYSVs9dgNhXj3nl33rgPwHKq9iuJtSoV1uluFTJNsQVgIq9S4KuCTaF+uMLIzGdPD2VEd
V744o7EIwfTm5mlXhy3O0XM6i7ymt5GaFtyfSqZRLZYvHdqvRKlUsas3H2g6jCeXgeYqNsPQtUha
obevj+xKqlPAjfo7pNsfGsGyl/iqzEnv3BnPDA13irc3UsyUJeTkvUtu/+q6oAO9DaM68BkN8dOh
AtAsZKeWJAXJlkZgs2OShXI0HeKWuQ0EvfObb8KEMHIUzOkcTHhVaMh0b9V9NS4DbW1X1QfZINqI
/pr/i0P8KHHwaSlOFq+xPvROEvi+R4wE+xIZkI6AeBGlV/s0hTcLm6RrXsTSL5kH8stpjZ9IQ9sn
re7FzvQd8YKM+ApluVxF0SOnE4cVPu4jZ4XkGYJFUbbJyeoWlz1slhlriKyvA6MWisoNS32N/oIg
zsnZM8dvKkZ+eWkwssHOAtjxSL7jqRcqdtfZ0TX/DnoQmvLH7PKOyofub5J2CA3pko5enYdVYw3S
5pa1YwLwG0ofZf+eHdcULehJIEL282JnAgFqB+iB7kxXR6izNs00ysZF5C1YdUJC69noJDu/zFlu
ANlAlTTtfW21bnBhFd7Ge2EnpN9kRI+LMLLGyV6gqKYszSDOyuHNng7nLws+ZyDjWIShH3gxCbWt
AJj95bmfmNjsoXwIJkHAqAr62YNK6RCvFWjQmzZwcbCd0g6DQAuql2hE4rk7S7AU1jYO2/9WRgMg
TxdXpZYb7Aip6WMT6JKgGYFzvcK19fPjpI7S9d/A+tdXATK0d9UYwXRqI8Ue2PETCUiC4syWynjf
qoqB59v7o2pJlNs1M+iG8ijaSESfODh8dEspSdTT4dXswVv3vs8peo91jpC32I+ESp4cV3GBf4NI
5adToTpNIfRVmMrkkEfrjwLhydEJhXBzhB4rty22ioGugepsrDhMUkmQKrbzExk6RUbjhlNt6F5A
juTfc+8QGPViy+zrewCEaj2u4HBuy8TcZG+785q9uXZEqLWOvgMSeTsXp6xnqfuZWdAfd7IvvXME
T2/h1UoPWpCOCZZ3XCDHZjbli+2pCu570HbOP4w4gUBUfNRmbk94uj0hkkssfjd45pU6tHNVIsHw
nymJWWBTphm39Lv6r2HOFGyWxDh9we3bz6Ja0nC/cIahQjujNTW0pQEgRI3aXgKaGgr8CVs/4byF
mABOiEjNSq2uEBZq/12X3BLKvzmHK/sxAeTfv92yNIyYz+VBQRTAyKwLduESD+Y/0267wHuBpUrx
wOd8wqP9A7DSRWfHKIHBTVdJmqd4jPVreXsEaG1e6cnHjarfB9LNTInA9qCCKvQYZOnVaOZpeMtH
E4irYjYyXd6w9FnYSAntYFSxRCLIQck9IX+VYVfqdl7/U2He1myGUKFsFdVnU/vAuXA0H1rdC8JH
NKm7JvqMWNPA6b60GjB64KfIOXXzrv950B+gvrvGMy1hlDAK3jysH1/z20PuPSqApStvjKJu43z2
W36/EtzqqGZwS04LjarQ5s1QKKmUvsk89xH/LLsOa6KthRBkyDgqjoVAH54G0JAQyeDlJiKQmqb7
pIneb0OCOs2/HLRIiBN7gY/+y6VSpN0tt426LTKyqla4xro6QUbVxiMPq0JAbK/zgKonm+Voc7a/
IEk7kNH2VKbpckXY3U6jIznEQLCu4sNCf4U4ua5aW9/0g56+QE086I8caFfyycCG1eswtHHlgwul
qxFq5JfiqKTuDXMa3rUU/3mD3YvQ56Pgw0i8GWvQTymxnnPW0bdhVCuD7fYI9vPpBeVe8gz9Y0fx
jmaGVrBc6uqgUGZD+tAZaHzyMcIazXSOp4y4ZFUAWgBRnf2Q0+YYKrFJHZu8JVwuj1EQC5Lrsu01
JBbPEW38wV+fcIw9Z6yTnnH3m83rJh8RCWMI3uK4Qa1BwyHiQp2v1wwoOmXzYZeUMsRiNuMdMwOF
a79DQsjUfA8dAb9yPjvCcuj0FcnoosnV1iMAyX9Y/4Ajuoa35I5E/4UGJfyeuvbAV0FILUqcTEgf
dlwE0jOmcupN+VInxIkM3QUyeSpICMBvtHLbKdfyLKcqXc1/PGU/wwN22C22Q+sVcC99PlMgDeRJ
3bZhSXPSYjSPpoFatE2cTAhYpJL8o8Z/NSrMd2d4i0BENOVd7AmvJcXXw/TAPqAibobGbrh6SRdf
T8HS/1IRQKe6OPyEkdoiJiXxugwHU5qNvnMQM0kWuyEtehFaNh6ILx+VRt5wT5pPHX7pXVWr5XAf
L5c1OdJcZ0cfSK1s410pFsD9+8uTgx+VecxDHETI7jJg8KtagWgtg1SzvPNwVZaISSQ2SFzuhwm/
hVesDHTZBo9BuhIpNzvIkfTvWAnZ0P48MkMk5oDC2jr8SDG7wV+fP+53f9rYNw2nIPf5ClfeI8XN
ZAq+fI7S5CnEAmHzxt8mLUjPy5jQLgoeFYrRaahTWvtRBolbX7+Dc/1ueJ7K68bUCvjZg30m7XZl
XJoYkmDw+5MM7HzkW2uwq2XQRBnwqbLKlRWIAzfq4I3UpfmNswKm8WulwADfolxH4Mz/WMXhJwDk
XyzZmM7f+1fvyivyLX9p34uLdgvCHxh8e0mdOFInJAabQRa57E2y5B+7bGZLOV/xdUzzx6ppcI2J
FYzjbafMkooAV16KG+r+HLY+JSmJ9D7gs/hqNsEvEqdCG82MkI4Q4jghPbMReOOD7OoZ067v39WY
r9BbU77rqmdaULRsxzTRghP/ZqzPsJkkW4mNYgwwUloTxRyqtzaSwIm0eUGHmwpepp4bIRBaht9+
Byq3s5GPu2xk1y3JqMPHj3+pBLJdQsHmUEnjmUAmfNVmZMTChV3OtMGVPGcwzK1jig9d7lU3utL4
PWFQE0i1bB3jDnd9lFu/TeRV8h6tfjSLt5LS0evudlj7s1FR/FDuaHG1AANbGa6rDj5mQqta5gEm
zF9sAle/pW9Jlyb6XV+2R96Ron3Jv3B3D0WvIsdAeypmbTGNr/81cuuSvp60nLeLPu+iHfrgkiv4
a3fRqtWZIQ1mE10zhVTZW4XK+T7QLf8dMfo5ZyX/yOuSRccinO5rz7HNs2IwQXPozVhRpX5ZO/Ay
PRNHNKRMcaN9Mk5jHVkGzdONAgb1WdqrWZ3GoiE4V9cRf1PjHbFFOTst31NwGTi0XL+frYGrV1JR
UbHOqTuOFTPUFQW8gP9v4kvtVkmGEvKcpQDVRYGIi/lSl99tkys+RU+saPaVdOJ3nd/9NErqDbBL
tIgfZtxYJxvNtpuCVpGLYmLasEdlpUZK62n+SgKM5Q67Wsc7w4eVr7SAkskPd5JKH2sMBpmTRi0j
ozNEh5Ee+KZHhUzDZsrhpUbve+bv5jtPslLb69wGdsGUe6hRM1jA0cvp2IS8pz9GaBjbeiWp5ER1
se14YKZLR0f9mx4Id1hbz+AB6DDncwqTh7kxw19TzAdhbyV9pbvp06ETJfu6cjqaiqZ1Sx+fDTT+
ndGFU+bZZcliPsxg4ueCHLnM+BfbBgbPZSeqmcO8W1LyyWtILxJ2qF0fDnhpsDmjtNCoHh92qfdY
QfbQq1BZXPFSAl2GZ++8SIwGuANv4/Eor7kF6z9KeW/3IqJ+/LtSDN1JnNVNw3RPFdx6dZAyen9W
mRJ7luS7kW+ngL2tpLH9T0FI0eD10Ny+hs04UoCZiBMhGz/1gokHhqpf4KTDeGFV+W6MulLXX+64
+0Ow3H+s6C7v1MVKszYBQj2Bviu/w83PW3gIR2WO9RY0M/b28ZmGXmKemRD4QyKcKJOjtfYC1/qa
NPXjiHfAFQx0k+RmInaEVOzjYS3puGQ8d0UT4CZUrbro+hdReAJ4xjKDJC0Ae0iwK9hsfYmZk1jE
XjF19mThxpeLh3VV/9Fx6bhVo1PkEyhVTHfice2gSuz3PD6w2xddjwZzPMH3jEta2UaDIrKbkvcX
q1qmdAkxOB+4Bm8Jrd7pv1JT8VkU90vr8M62v14O8nCu63gak6y6hHAjnR7JFpQ/LSQsOrPlLMas
gOKdpIX7RqaIFJCgt22YDJHmkb2JcO6EQsKCT8aPQ7e4uF3a9JGWKsO7FfuRPEynHINFOpIDTCLP
kpnbSwEO+5UNRqmFL7pxk81Pqie5nCyMLkSZkkRXSAquXXq+FF4Ad9lcoIz55qm1KkZ5zSP21n2e
PAndAbl81R89fk7TlV8TnW1AXe+Ja3WWlcY3U8LllnOJ3h8B19ZY5skZK6Ip7c0CPGEY8THmLOdX
JTVBINUN6rQ/0LmzdW9G1wjmzEWspvg5OiAhfWDBPxJ6Ioo4jjCYeLYCc+8wyj+kak7bmJI5u5jI
Lj7MW+Q5gnYsi8RBqVvXuneYvcOOwKavGsOXMBryzcR02T3ec3dr+0Wm/FjItDuVsGzoKahy3Wlu
ICZsRKmA58wBBtOVY79zvsjYGf9SDA0Jrmu4WM+5f93YwfpATQqGOFej1MNp6XyPVwDegDWDajSX
vGGMtm4HZGqMeYAKe9COn0KGn9RPLoMc6I8ZQTCblJ1YQIM4yEXca19uJKYaCvNPEafe0I/5RDqS
OLFejDhn92zfM3+wQm/Vl+wg6/2b0vRKDkbj80FNRR619hQ7qiyv59sgOOyH6ij72NWl+jj2qyx9
1faZ7AVgBLJMsN0DPgf7r8bM/vewuyDwhobTuYisrOUrPoJ3CQQQJIWS4wPjlJARH41/0jQEtxcu
Q/8DUEVnFaf6kyZoaIUVqdLuk+qu1oGTOv2+MdpxAp+dr9fkLOJSDlWs72f4eEYrp12Yy2Pi8R0h
LzoFaY09BLvw2FJ8H7RI2AHifoVdCyKTtimlxUIlehXy3x+5N0B3GTCj/6CfIulF0iCOCS5KBsQS
6Tx65Tn0PkqcYPXot9Vg0qIrklY6T0drxHIP0gHOMe0o5kyem4W9eH+8Yejup2Ql7jwkhpbza7KT
ewx/Hnbyt0falIKNeHqocJsKtk6tdOGe7bX2X0BfpizTfI8l2SpsfMF7suvanyO+NOJKzUp3NQI9
qqbRlDxoP9lcFo2+wlE+8u8TM8KCTRJOkCSugq1FNyadPxtKn6DofW6mRLV2e2l/hiQB0kJtxEFd
rIJUZ5Fy2MlpTHyqE4AuiNr4af7p3ZSzW6MCvreT5S8t4d0BS9qNn+jfFfA7Lfazk8y6taVLqwbp
e4F7o2peHpUHhR9zho/zG9yRtKRevkXsgomoKrhtb0uE5D2E6ykhir17ZtpDkqcAEBfSl053WEHv
WkXkS/iqxH/Mt+LOxG5W5yvwBptP9oz/NIsivClBg7q0EJhDPfVSzV+H1CLs/HqPuN1lLte4pSWR
PxRFi0SWnC5xBDxMZUo/yd18H9zGGhH/pKo9q0CTuesV7M80qUqHXY4zRZZjDJW7mCmdyhOLLiww
wguqWib5T3wX0aMa6/ZiAL//c1DuGsqa1dlBLiCxw77zFagyGOVL6a66CF9wDlvl45xfYsFrb1f3
qt02zKmIaCOXsv45c9a5gMvGooCh+c3Vl/sfW3ORLjtlLVjN3bjRa4iFZPBrsG599+WP4lB4aj8r
dzT8QZ+9ulfz8KM1S42hFzitkARBAIRNpgIcP7FKgVfzg5pDKr8axZfASJQ99ddpBElj83NHNKvV
/ixn8jvAegY8/nQxRhM7um9ujq33zAC1hkws4stQYr6AimQItNxPyXSJlNZ/Zr2fvd+uMfTt7NHQ
UROHfrZgODUItE5LfUly8BT5mgYN1g3wMMilOk571wEfbtfKTbK2SPtrKPvYuDnZYKyXCuCKsI/V
ZoHvUV7e+AVEEZ+iC4vLSm118AvCPAjuBNxVQJaJ+ttgjgGEXRxG1SjlFOoJCUTClgSYb+CioBYG
NSbfMivBOud+npWc7LFFSM3PWUKNyDrPDZbsjLRD/eGwOm32SJlljBz/kdvBYdlA8xwrmhMkEyNd
OKx4QBAReJwhgR9udU3wOQpl/QLvBpqZ+8dVPm0sfROJZYKsGibAQxjgT1SEjAEuzdjCep1dQO1l
kduBXkhnfcpKV7lilDYl2UXnt+oTqHTwdOmJsf7nGOIya2wkVilk/jalQ7P0k9UbiKsB2B3TCQYH
ch49kzfPCttFDAmqxnfQeqOgfDACSabTB+jluIS9PwLcZoWLIH5lj7aviOTxR+QBiKbfkImiQEI/
HbOoT9jfmnpyGovzeqgHGKnFCFH1e5aiF5aS64ErnVrOYv9ixAe9NSObj65Q2IfDPNC7+XuoCl71
jvFqhLA7iAO5x9a3q7GKCJPCZjEIyg/C1yTaMYrZ7jJmoc2bl/VlFft+jXCO9X/l/haoOagtwic4
V2Stq7Sko/vfze2tc351UddhFFJTDjNgz9YdMwMBEkGQqnGJREZUK7oCGXqiWQuQsNSo+lD3WeHY
PDFmgxUuB7hVU4J3wWF6Sb/ctI9VGzH7SyASNhaNcbpsw54sEpoOESIx1SMoIAiTr7MROAwnz6Un
S2rrLI9uhZ0crRPTCtvtrc8AupOvLKrniofgMJGv5q8dIqMBcH3HOWJiLW1Ky3ZpKx0I6LqvcS9V
SU7a4seggmGwJlw9gFHEWLisXe2TqJ276zOg0v3x1MoxTw1wxieqMQfORWBl04TnPO2RNUr4l2Mz
qxxmB3muRJBuKKWT/ed+gO+fBmRypYSFgueUEgcxj2uP5FkyGTuso0OyOGkHHnq2eK4OoE+5JQia
0M11u+E0hB4ZgD/UPSo/F6VbPslqW0IcqfFkfCH2sC1oFf6shLs3of6eqH5qQlsoCsWEaFZXlREP
U4aPQi3fnY0MD1l8RCKv7S/GHspCD9eYAhuRLZa9sWrqhsYvWbu9ptZrZgr21o1jhw+eR6g/7jOA
SBtTcczrokApmdP0t8CRyTI91eNXCz6mKLWFNPsBgTbqL2zM08frk5VodvENS6Gr48FpBkvupLJz
XN2Stj15jjr8MUUGigMTZ6jXxDeSXJJ5HGAJr6dPB8Ur/VUSOgEIti5C+538DxANNRq3ZVusCZ0E
A4yUn3T0o/RFK2cgS8KIGQBKY6iccuW/IgcYOr2i5/P3qoOwXpkkEnp89p7fWEn4yQPvdNPuAuFb
eQs5Vv7c8AFxUxDAznCu5l0BEy6vFAWiKSyjHyTtq6bjI6rsUegpXuxfrNVrX/6MtZ02PUm/UlOX
Qb148LGkr1Mv2h8VVQvvsNkrJZOUUl03FRppQjJ2/3DLbT8Vka8L0zIrtZON/DT9xXwq5mKBBetE
QFjSoHREy/bsIQhrGSQJmyGzeoVwMPiN55bo+oCJPON3FAej7Ryd9vEbKO+BNfNA+E09ha74NgeE
BRSd8DwfJnNnghF8FXTMXSyPEdGw6lSGdEPraUMeRSFxisRImYHsDWt+l1TqmJQ1O/FkUslsQsKa
4kXMlx80N3ZypDQhe7I50kcDhGLDFAZh3TRerwoCQ9izRZFEwCrSkJzNH4eQ8D8c3x2HiI2SDkIy
XyOiJYHG72nCoMlG//iQb21jACpN/1JOioS4Mnwu40sb0hGSHZUnXZpStIPvsUXO7/f2OWyzK6wc
hRIX8Awk6IKrsKKgodmzvT75O9ZEE+EtfTKSyQwY0Su7lBIGtWFi28Me1RPY2/NeQfigpxIF6Ser
W6JsJsS4tzI6jtTsV/bkcKalgKv6ZKYVi6j26JqRchRU1ixtFsDcdn+D8EN0LtmtobSO+ksEaGqw
7cOfQhDjYdCC+jTsQ1HjdTXxQSVK0Q5RTTiXufA4bBVYHnx1HnCl4ZGOFUhSJwpp/F4AEqTTV0Ul
71h4DJQUcTjy8DUgU4KCeRaaLL77DZKYkyybCz0xNfA9FQKHF4j5wVjpCCmrS9eBWOaC//cmUOKK
DJ/fo5BbQMUeXctOAQq2ukx1M+L3tJ77lww0Dki5MIIiFLLGG4wE9TRn7xW1kSgKGQDfAM6at85z
G9ab8XnFUactk5NhPPF5g8T1P6nlTi/uhq5r4T0JexBRiYVUE/Y51qzBbnA3y6vk+pXFJmgDOuBx
mPi6YJx3+5gxdpnrAdb9aQCjJJNwA98f6PLT8HhyFdvwggVBSnUDbffFQtg1KLBh1HPZZa1nyFOd
Bc5LfI6NGDMQj2NOWyrzyWX3LwNt0ROvojfL9cZVgWvjnfGo5RqCQaLw+Pv72y8tVSCwka4EhE6f
PIQiLbDqix2iUd6usvx+9RoUApLuXKRCzS7cDduUqbyq8KMpiLm5mMcgidP5H2WnQNSk4JoJXdeN
EHdJokP4rG8D+8niYBKnIS6E16E49qop4CQlFOB6pnJWVMhBdV2C554yX8DRUDV3e3THCo+nEDjb
OnZ3aoRXaziKSGGF+NTfAH4qdzhGa7E6FoOW/FhhLW50EHBLoyx3MbB8xOaQdJ7BAtVzhqQN6a6Z
ujmvsqu3Kr4r0irhgT2BjhfysQsLriF7G5EUg0pydaw5Is9iP+3lFFbeUzx5peftfSTUA9dPlczv
eVPLRIQOyerzf9/UWHX1kvWOLc/rNoE+uQUBBugUvgBaxbIfwIR2uc6tpDxwfRRH2QOrbOoFevMi
p9Up4ruSH8vElAMYw+16cg4QQSVCbyA4N/OSumDncbOoaBMQL9WzWThe1aN0vq/ugDgn/F4G6Vh9
lHeq/tIl2saJeoPyBUyp7/TG2qqYAp8nAT5UKgajlu3RelZGxwwwMr/dQzNyV1tJQb1hhyl2jMWu
0waSdYp1SgPj0qGB0SSvYfqEjI+Cl8nlOS7dg1CSP/mr0l6lJwLIvXt89WbcU4WKkJiUzWbOdBkq
Pmbxl2nrd0bNGUx4ZJOjHk7TY4l5ctgcQ7roxDKGlzhUFJ1LTijOAUicO96Z8BGdXTOsE37nvtRQ
744Uk8e3ejsjLth1prJ6XAtTOTD6Kd8zXsoM+vMiwYiNE9MYgMOeuKZhFuZUoay/FvEg8pz1HQyr
J2ykxM7K+4k8LlTrhzz5OR75En41Ey6iNFLv/1kWIHCpYEQla2PiMcU0/anqwsaH5u28AbrMBVLD
2xbkD5Obsf3QoPSN28j4faOhESSAacmFHHXNiP5uG8ykuo03/ItKbAxIZPpqCKRdaUVqabgepcYN
VZ2ccTPglUrMAjGGirE7kBRdh597ET7jpJThr8CzvKiXXPsiLXm+qCPhOrXmqMgqN4U3kLN6MRb9
nztpMXY214l3xfrD+5xYwQ0G22g8c4EEmeZ8G1StvcVEMFLM5zOB2WhwdrZGeBPe/otDJA10jDEH
He7utJzTg1zt2lBPjlZo/Mel5CLcB4E0wwRqDrPAu5xIfhEKj0b8Xw5mhQH0TYNzMw23j2glhDFs
UR4OwtMbV/1MBNX4tu6nAEd1dTBFw/tW4VlCiEHgjxLFFozuybEtSlOVcdpQ1J2kI1m4svgpbCD9
oIXP19tYGoT0Klzk2pn02od+/wJJquJpqrf3JxWZWAvn89kNflx5Q5iYpUb6YvBHeT3mBQysY46K
Izw/A7JmrngHeghxgf28PwGGf6ESAOtSmAWvt+2JWbic7NX+QGH6l5/Ro1DX7vZCruN9iWDuzzO6
Mlk9bX5srv8ExPJEGyXQkXGI47qg6iI8SLQ3CyeS8je+WhTbPAFlKpOSOmmYIEM5/Rm0KZY7Gdva
VGu47xOvHy+3RY2cpAKthgvcz9izy5f0UjCZNP3VVMLHTNrvKKCX7FTCChNwZLKOl50j2XT2KCTq
ZFPiByHdDeCkcV8cDNZqHkqKEtESUAsAh00HklmhcQqbni1NzOzJ7O2s7Y2G6i4qNP6fJviUPDZh
4c/rH7LDWzAGsk+XoYS+Mm556o4IzTjSou3c800UvAmYV2m6/WX+FyudSpOnZBxwjgiqarPg8Qcd
wBTWXwwx/TpadmOWNJnCnzT/GXWu3Of0vGzMRGNcCElr/xLZ6Uj1181fGn3deGQ1+YpUeNF8JKej
fkGmWiJHzRpKi/kJ39T3AQHG/kOxEU1OYzvvweKyBCg9bhRs2r3pbaF6utAwocthNx9lCqxr427B
w1qK/Ir2qYDnZJF3xtJFAIwlsVBFxxYKVB8AfLS7m9qznecTlUjG63s3dA0v/efqRe6p6fvGO0qq
2vZp5AQ2MXlykHzW3/DsP6GpCdVdM9ZtOOT5CJUpkYQ9PhX8chlQ+lliL3DtKZr2oXzCftnyvUk2
/dS2v0zcBU0KJ+GfEHmi2+Azn5jxCe/FE2jwOPQrYk1WbWTdpMf4mE/X1GbnaSTQlj3mwCmjgoWM
mMSjSNHagIFOBLb37INaKsI+kUS/FcAw7qFCt7iAk5szXWpgdvoSbN9RE3EhliD9+7bYlY2n1+q2
VtXYn5NdkPF0RmAM0dPrXN8+o5QYvpE7mLsUP6d+sLEmEHlvFndRewteQZLTxnj0lUsIheDMrQCR
1qrXqlFaFqI0ThlIwl/dKoLMZcqHhPIq5OU4TsSZdV7+lyVs8lM9bwRASSkMT4feZKaIx9ksrqX7
5ys3M0CE7HwlBZn714xVneMxClapVBJo/g4Xm7fVz26xZGGhafRi+IFLpjygbTiDAK8tUqosJXFT
iFb9r9kQC6R+6vRYDWJ6KQmEGj9ngqj/PNT/wOdp9kUU/b95imIstYDD9OMCtL707SgiFU6D/ed3
CMFM3XR9L8I9NEJZ8Pcddn82dv10DEH5k6iI/mYfn9Y45cdFnKSXDiw6bEJO1UXL6Z6rlj6mvJW2
I3kVYKy3Jw45jNrZT3q99YkGQWF+whfkr4c3kE5DpGLq7luRLphQS0nA3luo1tJjX432YW1ibeh6
Y6RsyBR2xi3X1AXJNwVu/+dHfsGwDkpw+I676Yat/SQNBIigXhuPakRQvtvQDmTF8Yh1spP8adhj
RAIhzjLGzLmjM290Hv6wkQ0XieHqoWa8J+hDTsrK8ppdSm2lFRF3unX/Tg0Fm54t7hecEiaRB+xw
U2uDEwJ0Z0t4rQQ/6eeeN2cSA8ntNXf9ag3AoiDXWqUNsdcleHhG2CCIrz8sWo+MUxQPr3BDthzE
q3QHE9msNfdF0DilOk3w5tMqzW3XcP5N9w0dT+ma/S/Ntl0gXwTmA0y6j2UOvsBJy+73iKj+W5U6
UPak8G4JveoT8wQh16T6YW7dhnCwks3U8akeVvde8Wz1IWWCcoaEw35fXYpTBh2S2w29O95uEu67
T8mwcY8gwBligykOeR0x0yMlMKtdCIJ6TWU7uCu1zakyzaEGNr7pIXPRKmL84vJbYZ76tsJTVbrv
uV0107254Y+1UM/Lf9VSkepVgDLo+BOZFyCyBBgGPxRISocQH/VXqwfTH9luBimrbxrQnQdQvz1T
ClQfs4DK8OVAqoC4a2ObLM/SkYZ67eFtbwZD3fHWPWFOazrAPX3cDcCBAp50Wndw8oUhSZ9GgFh8
lVF+eJnnhmufgZg0cq0IBX029q9a/7P3cNubHeeJ8LxUYKWZzyG3O/MvlZ2o73m3lWv7MHGvei8c
V+LSEX6V/mFumBKYFe399CK5O06gtWoS6RWrWBA9C8sbw0FqNdj/qgs3OeN8FhIt5rjkrKqhARHw
59rD7f3O/bvN55JzjbB8+LDdUtKD/LwG07UB0i1ec7ZLntpJlJmygtw12ZIz2PFK8q+Ke/HlMZXQ
v0sy1lKwKPQlt+sltcdPBXHk9suJmJmXRStqeBRH2ZPp7Kwldnk1I0f0swYyVAFi6KLLG237sAhw
A6Eyyorjg6N7rTZ87FecP2ybPBdLp3oPXPA+VgBvGZnd8NX3hdmyKMprqipV2Ed51b+P7uOvfkqn
MKqKTtM558fmV+phUbmqVKvOYFzz0D5H22XzB08R5NUH/9ZOZFCSR8TrvNPAk70LnwH/rmNVnn8A
7WjqC3fH02CozP42s+6qmqzhPyM/AIUrrF/N2nf0gOe1z+ZLac8LM6eZAWPqPrcMJOxuV1YF8ico
YZikCYPNxhm8Pc7obBOawrnGOPXoIhXJIPLgajl+zYOJ6L3wBBcISbjdhaIvUfQgSFxdXA2WJJCM
jr758Eyk60aJ7S400TDT3crL8+OJy2sxoBr7gzWZsbXHkHIsn4TlRWVo0t1ZIwuENim4SyrHXSXW
bdM6jrO/kQ6mv0ysiRd90NVgBkIib37BJHMYc00QEqXwzXJv4UOoDOulFOt5TNm4NUR1U0Baqy0h
hGaFnP/jMu1PUmqYrAwI/77s0F5/bo/SQzDrzeW1Kwbul4Z55eJ4m55yZ/9ZrlVuZKPmNW4GSseM
P78QkArwWDg7FG8UFBBM4F2LawbYbL3aORv2HkqynUZEz9BsmR0iBX/QEJZVCNRcaCiO3ZL6ujL6
uzcNUDsZQNNY8q9+AgmQZEh60lZpIOVe7ImTZ6wH3q5edIexj+iPj+oU0TPBytQeNIdmkr601jf0
2jDi5YfFGrJqw1zmJZIWm7uhpntuXEjYXqqd6g1cXWn5Av1B7IAVRzhIEHxzLu7m33nsUAm3/7IM
BlpvyihdVYewnK8g+UphZWkjbONgMmvD0PUC60eu4HuD6v0UPvBglRALFnJy7YXMMAnRrKe4gSZr
xDKPWWP8VFH/7Jm3OFbVC7dsU6+/3CLPPeQN/fjeMDZCs1ndX7e6aLdFCS9PRIpmGKFVRfldvcAv
SEfHuzPMEdVnLiIwG9krXJY4d57aA2mToQykWjvSJXsWuPvclPegHo9S/TIW4ktrE1skivsHnFkN
1nRrEwSQVBmMJzmJP5Qhju8eGK47TcNQY8fUxHC/qiWBmzzHR7IiMScg+zCxTgNgxi9+YUnaeXIS
Ma/pFj5OV49Hnd6a0iIpwjSA/k4AVTjMPOQr/Tgb5gbf2x48IobaZIrs+tKVF4M8U7Tda9ZsCdan
WADESxNTlC4mdNaLHDjYMD3Z4kKa8YDc/5cMjTBsxO7Vr40pOIygOUs1jAS6d8Ld8a1vDFfUowTf
gIgiWG1jW8mhvPXeJdDtrkNG91qnunLvnsQj9SSTFCJi0KlqDi0tUYqPlKXhey1/rzoRDGmMUqKc
l+zm+mMr82l7FhaHfKJl6SFbns+B8hA2Yb1T7ADsa87RXOZ1qEKmjQ1YDS+ldNObI7HrW588EpM+
jMDYZ05OvNAP1NQUl5RLVTfremDne1abdIvpmtVVtS/w1PYzQwTy3ppAYJCAOONsZZX9zFeeIFF9
GDPDsbybhokWvnKASsKMT2wDQGcOhlVrvnMNC76WgSbZ2EnH/GP0ndZMrK9gUaoCTZUJ5gGplhFh
GPYDB9x9wJ/pSAKyMVkUPOp3xBrH+6lAWjwnvU3OoVLjr3We6/kDS0KqLz1JBmw7I1y031Woqiw9
2hO0kGRHxjpAn1RrHiQp4IU2J6S9UE5PlQZMCjYMcjeyzU2PsM9OR0qatT4PBalNseYJKxK1apKD
D35ULu8Ag5n6Iyk/7LJH2pBMkdEt6rHq56bA+JgEVSEVLwNBJEAA9+dDYQEmTw/tuAQ184nF+wYV
Mc/a9jBdK0Sxgee+1NtlqjEoHEeUB6aaRywgsh+ZOVql1pLw4+Oe2jw0CKCjuAr/1lAf0+OkekjM
hdu7iuhq7Gi7rilJm/BOsYn8GFt1iZgfM+rSHkPdr/YFXWZESmqBbfGMKk7KwpeDlXf7Gkq2k/gO
t51QVMssQNj+NAWK2w3u6rD9UDLxsPVtPz8qet//QestmPugaUiHTeikQifKH6WZD87syxZAPcyu
rVu/nCd0Yn7boeBnkDlm6mehM6JMHuBBJuN5d6IRqV7OsXEpcqD8VSkZp0MDKZeDFLBspGX1WZmu
EMPA+V15tYmtP0LH2gSs9B9tFZhtEtTAP2YHDQgT8jfGdhErzqR3po/TWJNsiAfBN20wE8G6g3GB
JyLJtYjlsDdzamKplovydtjwVZtadGWMWiUs/lG2CDzpITCJN9g0rC+W2HLCh6jKAyEuxzSK2aay
KerCTbWk2LyRdDQrHiASRcA0CQgKdNw7rd7JZLdVx+uwX0BbxEd/k9XO6We5xQd26tnvkWzBg328
yTq3Nlww9NHGRhev7fICyXwLyUk67QdfWkpeXRgtdheRCU+Zxg7DoSCd92UYanTuLEYPmOmcaVmo
C5dHxgTATY7YJG3cSflNqXo+fjuki+LHpb7BK93hnNFoR/wq+wla8c8b69jLCDN206NpjI4vV6g2
x+JkjWel0URS1kzGNJS/Jk6KOdSnxrD6krAl8MiEO83k0ZGWtrwizXd6OAIfERMrEIM8VqFuRooi
5WJjIvtRNxc2Sb8DgW9WedOZiPdkWMl08LnWmpLKhASX2XDSHGARINiCUOU34FYCnNpaNg+Y1G0+
d48jsppNei+VJzhBIMEJbX+YwWJr2adKdN17zgujWhtNVHuKFBWfP9f/HlH2Akz7Ia28TPDFFEIf
CY7AdkNBV6a8Ige1DdkSMcOv0rF+WWIbtZ80pz4Pj4N1nPzuDNmwzE/X2RrCE1WwyZ5o7GQSeqN2
vw5MSMnG8Gg3VZ9HZse6VKm7XAzRjyIefj8Pucs7dC/u3ixO+q2O5tmQECTRlTKf2tKJLKsppC8m
l0M0QeuGlWUem8SLgKDnD1cRfmAP8IEnRxdX9Xgz5VDyyoR6UHH/lfAICcpj4FqQFY2UmtytJ6IL
QRvskRNMN9xPP4E/Rj5zpCI/70t1gmRzMH6vR4tYjQC602wwdB01e3Bohd0FM07YxdPPALyGxbq7
fr8iExnWXQXCP5snRSjKMci3bcVZq3fS8MD9YVryY2tgmQTLbBQY471L695rvZNKlGXHT6o+QPag
ZmJ3qDWR0YvDKvicyS72X1nGjBYn8E2orJtcByR+HhXAFGC/65npf7mTRV25PHWsWHY9Lz8J7eA/
9xvtN9QWN3yQYAAvxQjyn61mNRfFNeYfirKQ3PwPbbHLw+/5iRQP6XveVSHNvXeN4dhdDV+mH6Vo
ojXd5N8n0BEJCD08vH1PX4yLFJoJxYLIoxiAOOBJnXt8YCqUNOtzq0niStHIIA9yxJSpt8EuJNOj
ct1i6SpJfWi3rUv8KN2VGNMpZkcLZ2wKPz1jvENXbPWU2HIZcQsg3tQYEQlowOYWa9azt5Q/0yqh
eToi+mypM4d+h1A5cNwdKswn9UIHX9i9y8LsOngklkpbmmI+xKtrMwQWs9X6/4DyRPaFe2VAIEpm
x7Qojxd2nTcWqbd4cjOkensp1Lt65zfH76VcgaeR82q0n7J9K91C2yp0EsH5mY+iYsap7wfMvdiY
oQKIc16bULp2Jr1mBa187U/EgfPg+0xSXIaqnab37BZFzFuJhxY4fZa3JAaXmALVrOc2Wrbydylu
fXdxLwXq4Wv0RXrj7gFeKHqV2ZFNZKCdytvm0foxbxx6k2spCoH6i3FCcncB5tBTxw3dqRJC0zOl
mnVuaLGx6P8OV1uDuZK+Dy8fbmDC6yM++bWjBO5/lZYLbHacbMndT9X23lonE6zZsmfG2++Z2VmT
SBWDLGCQlLwB7vB2Zs9D9TlzU6mCCbuK7JDajX80JBmQGRV5j6V1rOI3SdqRKASg8L0BOGaakM5H
e8TB9FChqKTE/C6LIqCMoE/qomnHAETOxSOaxuyPhgiPhBp5LLckvwbcJtUXaEUWdnnYd5yOStV4
hHbd3I/TfGiJdv8dnpP2juEWrD5Y9lJC+5JM5aaYAiEIehgNPX259gia1uAR2teuWhR4It7l6sFo
s3a9pVGsg4aYCqqKSXeqh0RsneGwL+Y4R5mHj4Y7zx3wRKuNSd9qLkzijlUWxqEvI+R4YxvYZWGv
H6x/KNg9vmnznFYeddZ2npjT5VcS0yZ8WiJYdj6qsOVynkV7zhPYxjqamaXuF4AdZs9BzsJvq2G5
D39WxtApwNBm0SfIOFJ7WUj273reLtqk/jXEDbY8EljO62sCef43l1sjvdgQdYzGmsVZpVwwnwmd
JPP309ompWRE5X43pfuak8+T6f/qA50SB0CZx7T4J6PCMWEAbxWSUphSnOxwnZo0vdk5EJyX8S71
vCQz9DbiJOBiorJtdaq4mq1fFHsiikU5JGZiqUOW0Wv14IU7EF4IjTfB8TA4vOFPzBZXm3rrOuKY
5BrH674SIwFjgoY94andQGzdFWV6/AEQa0rq3aaSuu26HN9aWNT9UBhbyMaXOmFwbW/xb+2NKzKI
WoxPRvJCa+MHWXeRybj8eyHh5gSs7DygYjqbSQfAQi14J3jGePEqivjPBTzYsYPvAdYLCt+2Y46Q
AKiPwMMYaBRghVCNT9NkZaw+jXU9BsJfEwapZoWpWsDW0Kr6IUAhrliw4YnNOxi+OIgKdG/8K5lL
TUOJrsvFjnylUbnH28DMUpeDf7vriJoojAfuJqsuHXKe9cIar3VtFxca78s/tYFUuL/xG3gOcvLk
fXmf9TP7fLwf/uKYAAmZ65gwnpEC+LuYBdQHORl6kJPqyGtpIncvgw3zKbgkLTx73lRi9ysoztPk
BUHVByLf5kTNOZkliPg4cWokwD2mhXrqyVar7p5FdCtpA6PKXF7jAIqOJPWmu1QWNA36p9DwYwJL
sbCRykTFdnDFwqiziuzR5xLJrkKnyaBnPkAZz+j7MbT2FH2VyKAxcYFTCuT1Ifv/aVO/fK917FVF
/DQ9u+tPWTHusxX/Tu/+vxstHpjeogy0l+8qzr1HCPThe8Xm1mMmAIxAQdG/x9TB+H6js7GLYoXo
fjJyVhjeZBlsRoT7tM7o1E6YvCkPc0t11rUkJ8WVLlzTCAXumAZkTwvTKW5AHuL5tD8XVNQRec7d
E7ch+pxajO1kxG/cHtsQ2NllVQ+dJv/tijp1iWTaABiSP+Fme+pEAJoudhl/ag/BpAe6gxQmaseB
eXMZK8lpW5zsw0sbsVGOjm8zk/UT+jHhc63F6/mPaODWnZDy5KM545+WTu8tb18zbXYqh7KAs9yQ
jmn7wlS5yS9B4tew385srVi06WeW7eGSJ0wY9X/21rx85XGPruEsev90ID0DPfRE4gWs45jXgvGP
q+Y3PfRKII9Rf2i8bbZshsWDCRXvhWBtDYnRvG/JWSDrpx1mYtsEbW1X+AlmcpI0wl3c9+bIMQys
roOFprodeVdPDJh+xUbDDMsAUwGiO9dygLCj3Tcgak66OdoiRlHVfV04L/YqPqcbgFY4BBFvNDGZ
j5CAgpkP2yA89McsXwjCo3PSqfE1RrczDEUWOp5CyzZSfdi6RB77UYTzui22CalhZbLnz+RXdHaY
X+joTB8iv23Q1xYaOfm2vxNoLiqD1M7PVfhPHGzyrRxdzCeLd0kKOYFJ16Qn3EWFJVnDcQAPIut4
peWgdRgJ45AVoQOz9X0bdP6Xk/Bzj7BzNMYZ7kV2w1liRWeeuF/dUHim7PoDH79wfeI5yc6nUARw
gCD/aXRcS66Fd8TdzQb1md9z+GYO5HeJSsdx+F+wTY6tHh78cME0SXKQiFghSVlEyQgDe7sI4/mm
xbwW3wqKGpqwJr6EvtZafoCfPG4DGLPgFfkyBLysz3Q2Usg1W4DlnmqiyCXV2n9+wX7ybcmfB9Cl
Wftp/Zz06NnboPDUs2wtqnJ9P00UUmDCTK6m924QWn//27Q08xGCG7+e+0Eg1E1zgJHBJfBijph5
Sh5lvQUFPpW1YfiAQ9q6rIzAskzZnUCHVfkZEZPvJGZKKvG8u8M5nDGgI3Lr7RhFKnf4B6r7DWH+
rbiTCC2mSWUc/oD4cZahGBlv+ITY9qaPuO+bQM3U4AcXEPqGNRy40aAkIkZZwXWEAmDGUcsSWc1t
rwzc6n2yr8ljo9fS9+/53yygp3svuX67UEdx2nG9GQZxuRO44wxlJ8oWqIv+MXReuW2WMkadtgUI
HFCH5wy+EC5CuJMeK9pjqk0EKdyLmq0x/O6+uHulyeAYGxXzCkDIgFVhucEUff83Wfo3/FhuH5nL
Enrsz2U0NPzND4ThFt1WFipCAFmnOSAVqV3C60VwBkO6B3k2Ve3TCAr0jCwBc5nXxDmpsKzmPhMx
615dnuegpeuEHfPkdOkuYDt4i/D8acJEjPI7/AaOINguZGndECtc0Secryg+UYaNgLTXNFLtisMW
BIqXmpn+vkAfl1Iz456n5FhDYuUoGWw9zO9vRPTXdKNxQCjtto518/CsZUaUpwi1PGEaqfpph2VK
Wz3EHEhdm4VEg9Mzt6dloYyDAbFthEHwaXCq35BF3HO++p6kGa1ZIlrCBXN1PEJgA+rCxMcl2MJD
L5r/0g1euLR2cEQJFqtZhuoUlT3hyT7ZEtvxJOhF92+Bg1O+VIHyDdi2Tr0/PhGyyea373S9jIyh
WzVVzXSpDpJrk9PkZytSfeNvWhV3mXw7zx+jw/HXvzGuibewagXeUPIKVlHk7aq2s3n3MPcehL/w
rOa61uMCLgcrwQtGFuklpLSLq29isYDQbkb3wEVtKQOJPMzwYOlq/zhLq9IQnsh7EREr2IaqtbNx
84GScKQ/Yi4CN71ncAgO1POyJdLM3gjbfzK8MGknroCnysFBGKNSDYIEWKpryMGe0lmzMQdD+qli
7eZZQvt0bv7PgVl1S5vCj6kIXt+HfM9cWZhfN9kW0n3IHXXa5QgL3suXRRb4MqzfjnSSA/O1wUPL
HS1iPY6QbOK/J2u57GIlxiS45J2yrxtUZfVMb7TCne3JExBittI7UBnuWpXGROLDyhjHeZoFuBeI
UGkGPkYM9jfU1rhw23ZFNycMp8ckpWyz993mFCVNgA0ke3L2jezigfaz4lOflVvToJuJHteJ0S1H
Mv3ELis4cn9D+slNULgc5T4PSAXwUMtjyEKk4Q1XcJ5eptT7yddoUOJlgrjkwEsk2Qmjt6oY5t+U
16C0wu30O5sHoLVhSeTIVTpkTLAZknfc9f2FWpCiGx+hPJlkeGvkv310s4qj25ybiGSpm/oJ8JGz
lQg95fmoY8c97ChLIQbxoixS9X3egAzk7ERkdvkjUeVFG9OxeJq1dNkiLuLic1i/INRMWb2ZzOfj
Lp9jigP8yNpm9+D5XpEDTYTPuE34/Lo0qgls1bnk53NYixjLnN/RZEX/JkgQ8tlZi4vjTypU+m6a
+tgObDUXbTd4P7VpmM99625I5pcnB+QDtsIDWgoIRt7YIRSdzBZRhnAHRUclAmT85sV+DpTjA8fe
Vi9rffhhA+1SG+ZG79TaQyH2gdNKkog5jDPfqULYkJmR2uxVoC1V4nzuekhDzBkaUxjBhv0y4R4Q
9NQk2eND2J5ADvamO716v1TMfPQGI6yQKQV/1DeF1OGWW1p2ZfgYM+VvZT147pYIfHiXN4naUumu
TfsdTsoU+FgzcnZujjLdT039UmGnhs2g6g3AIYx0tV1Zg2pZyy3bvgImzYfLwXfusR6DY2Pw/7zc
u+AWILyHy0ykMq+MYD3YebWn3jB6GVFTyFF9qkB6Kx0E6uO1sSB//Nt/K6v6vS0HhfNykhCnBOH8
Z5SnB8blR5Xmv/QHXW1ScuPKoTj1kVjw++1714p2BewKAjFJS5SIoK1+95nemh854seMx753g+Vz
dFVH+j5zhDAap+QO5vIthXNn3Jq3qOn2nn6T/TgZfoZkmCohbJP1qHQ0i1O4BJk19aWKqhg+qHyC
RmHDo2u5ulmd3G+Th0slWH8sgOJ7RMxb1bMZQOd9SHZFFwGST86j12eBLpjkoy2ii9rCp6QlRoUs
byzH5juBmX9zIQMRI+cf3Wdm0CiDonBN5vrLGJ9xohhcVoFcJMXpFwmyOYX0nnRFaVsZ4WHrc3my
SOJ6TzL9A9iknxZQATnPBItInyonhoRK2W5euTgmNw2rkvNYGQVZSHU4zZTAUkTY+RR/A9ASX6b/
N/93SUqjEWssCiy6iMGssW6k9UFC9lnbP/pqu8ivJqrM+oukmYqQ39u0ayz9q3pLW/WPYus0lNde
LBD8de5QVOX9JPboINlr43xsOB5zbcwyqq6NPG6PoWR1tcN7ga8rkQ//4zg5P6bsM64gN4Zchr5Z
v9hmsY/3DjvPHmGNjxF0o5gmgKoMVrNcYq4gRYClyGqVjOrQpOd2Psr/CIblCM2AW3hLN7NpXxMe
kACbG+jbaa4pJD/op+uszJO2Be7vOo0tKqN2NK6M8KsJEyB/nDCvGwO3gM7c1SEgx7hSNpeCSIBm
RR+5voAPZcZCruFyNUwjvQ1LtzQwxGtLMCGpHkSzJbaH9eteYfyokPCUCmvRMusyBjlazg+gyMo5
GDQCYpohf9eyhEvlUrtCqc4h3GSY+k+pwi7qdj9/rkinougL+TOLrMlpdmmDHkheLeHcN7nnb3mx
rq5eHqq1CE7PSUobxBG+RwuVQCq7cSuxncjgwg+3J0snobQlCp0mrzhrYsXtzABeQ024WN4HBpmd
Oe8p9sGcWQteW1Cem60Dcy1/DRSug5zBBxQMPFAvYCj6yWmTNi9pSoEWIOjSvXdx9kwSfvxO9Hm3
yFbifjzXVANAwp2I8Oj3EYvLl2fD5ksyVLrKbPurCO0OufktntfweW2HwFeKLT1z57PKJhi3J1Od
zb3sVhngcZ4pM/ZQOcSUyULXIrIAefUQFqDIPoHnzZvFzOIWV1Kmk1i3UFyOXc50KR28Gtha6k1c
xS608iVzS5/COoCVfez0L7gkfB6E4PYhoNQc8EKvWZm+GDckvXvRyF1T/1WBF6thhtEdis8zisGv
J8KJnPBOAWwFrEEx7qPKXtg41qu6oCdBS/n3+sVMT8WssSAND9oV0fCwTs9cVlLIkwOK8gNau5H3
8J9q5oILHKyLZSgDw56HYzre4rJOhMspyoMqKeWyDti1rECUjOsX/bkETOtH9Bh17IX8YiIhjrb+
615Cg/sgHOeB6GFkX6L02K6KX+D819n+k4LJg1GS+W1QQFU/FdEULMaA738hKC/vL0Lt77yX0bKx
2YNc0RJ+EtEeEGMH7YngOPYj6Zr+r7ZwCoUBr00UGt9p9O2pqaNIN+hmejIiwpGl/RId9mZBdZpe
ZYYOatx2O2nmcnZ8a7lNtHV1ELK20e3RCXNpACkzQLF8RFUgrIy41S2rDO0nScqweMF7SYJRP2ml
y2LuIf4RA+XOIBT2hndDEBUNHtebKwSe1ktm4gR3Sz+N3onndxGSXWF1D7gnFu0Gso87ENmyH9+i
v9d+rKqh/tifgyE0pRpUXF8+B/2ZYYoMh3sVdi8OZtfs71wfanPLroESIJTqFFsEFknroENyhqn/
krYip3DvZ0xesJRdlNu4Xqjs9hSmB9YVDhBbFNyzgp4R9HDGDDoNOqBReP6vuvTXePKVEm1F/MXL
m5sbjrYlJqzy8GC485hmruGS2R67HD9chprmTNS8LOb5WqHRd7MDHq4n4Fiar53jQ2/67RB1IKkA
TMtFOKcwxBMN3AVWFL32+pfX1JNWTfOhx4VNvVGz6tKAtPIZOGEVByVIJraDsK5+sPo+9HJ8Oxh7
nBH2NnYlSK0GFKYPCADG78/xskwxouJFv8MSM61hrQ6B5h17JOrLFh3p81op84QLRgEXlBVk9ir6
yFrfkAvwIYFgCiic1KFC0KfB5MmiGmjhtqjWVezaQkp74KF76HCZWwMlC/SVKj8PetcM83YcN7xa
zbX6U3+S5HEhiFayhuMR+0TAYfkX3iFa0SyFUOxDZC+iRqdqpor514Uc4mZEXqIu/4HDp01Dn2MV
Uk/TGE3vEtyW9/fBNgsHSnqmB1ifCWSvp3gEFiQAmAIBskz3mCOegDHZIFNrECLWRQ33Qey3SkJh
i+qZLNxT2qONGVUigxmpUSJHmQ97+Fu3BYH9X+mMmnaObOnrZnxG8f4WnKKhXrGCWNn/58RI+1oQ
2RjM+dZjIE++QMeKI4GSvIWjIyU5cdU6T9kWuDxnExbf4xL83a9xXQLtMlmqHzCKbaSPkqKPCL4B
/HYZVA/5u/7s4gmClGiAd7n/4P+cGGbK2lrTcciJO1dG6O6Wz2B8wjrjmGqUhFMePWKDkoINsee0
qrHfpw6SZFsdr+w0RHP61+6OywYzG7GLjp0SrMMH/2VhlM4fNpiLOkcbecksSU4RZWXhvRvwf/Sm
IgmwZ2HxIMgdPrC1Alse6lOMW0Vqu0VvXtykFxjUxRM1xvOvEzLvPiYdHBLO0FBtMhxAWZHL5lRv
Deu6ePZ46FhuMyaGLOMkVgg1guRcdQo7nEIbDTIBKdbA+XwyBHNaY302K31itt28DhFhfqNDEu+H
/IoM81oVY077QCe5fx1FPO2uClctuJ0O9NM9sHGZaEJJfHEBT8S36XLZ4AT7yU1nuK5xKrXjOkHk
22VSEovCPlM945AqnHsYC9ZN0FpcfcLC6utc7tnUBF6JgYy3SCHiq0vBo/0psqTWUyLodmOU6WQp
eZrrzC7ZblksWpvs731xE5rhtuQtRM6tVUdj6mZdjL7p/JwH3FinGzw72dLL5Evccg2YNDh3Crbw
Y3ioXyDixXwqYYEt+oahlKbijx/shM1uuXDg/uCiPu2QZmvuxljQ3NPrvUWoCyS+vs7Nb0K8SVco
8vasTdZmh63ACoANIKciFH92QUhebp31ScUVTLzRLyUboYl/wi0FMejDo8Gfuv7URmYiEac1kLxB
M3Xk3SnOuGyFN3nKkc+lyJTvGnBJ3FbH5qkOxE2PSz8BY2PIzAAza03rWyCNZEsCJffntwpxwA7i
W4tP0tzHrJDLGSxlAOJe6qflwcopZiwIwE9felmeX+rGl2mFL1kaGLcCWoQjQaWUvvsWdtvSu+bL
gSDEfCWVBt+TxIYTr4CohdIQ263SsjcbOeSiAJczVke45+NGWiag+9XXvP7YgynU9121nvoZ04mh
WrL1GscAnPTVRKTrBWZ193yXwew2jeVO3/jyoYOOmBjDdvrQt8xb1N6f+t2D2XK7AcfoQUFo7zDM
qAfnY0JjStB4GnWLzHxN4jRzYgzKx8FIFITugSHX8K5198WXpibNXSwhF9kEe7TK3EiGyXgEc1Zt
LRni7D1ybO/3z+mjjzroyXsXM2U+DDmvF/6SCeCDn3UhZiS3Qj/vaHXBdMT4lLa/SOM8fcVbrTgH
DWkoKY1bBDj40neuUM/mQ5PWHoz8VqJv3DJqWmM61HGqGnHLCrKbf/txqP5ctVzZxFkeMmNv3noF
EYszwJ3EwkADQWYqyBlKFfrYeA0vysm8OQNzhzWeOUcKx0ZNM75mwQXYDUCCHDdbRhW6JKt7ogGU
z1R8457wkWKyM4Ql+dRnOnyar2N15Mhf7GpnI3y1DX10BQmHju0MGQMhb5cz+bweEVUu7J+CS/kh
kmLFSfKcKCnyT1l7rLxKZbOxYrVjOTCUt5sMQomZFdhFEsp3ptJQv0G3UIyN4mP27WCQnMb5W0eJ
aGbzfRE3lTk2sIvuITwYT7sascedVGPqOdVLSTrpiS0+RENunnr/Q7He0rzFWJWmlsUkGW/EXx9D
wlOW9MHmkpVC55jneOsDS4Flcen+b3peJFTpS3FK6GcKF6YLyshAyO6+tIrIglI1oSNlogySOVb5
I0iS8QmqtiZQiNQ715QoRxJRnEfh2MLhqs2cCqMhPVzvqDT4r19GnfrsUjwNmTnupfvJNcuBJdsE
e+0ojQMEibJ3lWxP418i1URqjE81ebIe9xJJvZa1QNPUEkNYP64AmZuN/YX/0zf1NfGL8ocrxFB7
zM/rhtuAxtqw4P1m1ZOMdJq1GELbLy4Unf/SzFVjIQj4b/pKIN7CUDGcYpCCP5EieDOiCe3+eznF
1qLhc4dK/5h1s0Uybopho6jW5zEgMnsDeycZZQZn+WOd9a0Z6x5MvAgFrZ1bpthdPHs2WqZf9f+r
ZUTrwXgjFKQNntU//0CrLIFESFpZ2QFj7YdRzxFdgaBEOh5PMavaK3EZfZr54e7Hrs5NYr1FWAWz
0NuHg2J8JNH8pFEwbW3fZ0lEDRkv8boj5lUR+K2BihOgvG83arltEk26OPjXXrfyDdSnjM8662SJ
4/lfUBPFsxdVrYuugHX0xiCBIblzOGUdN6MMya1ntz6cNKGyIGWTery6z15yBDLEHupgkXj1Ct/r
zYGu52U7jH3V5DYx+ouOmYxKH3XlLaas62pg2OF4XHltltTdwyk/DHijNkGndKbNdRzinDir6TNq
GHeqd7YI02QhEAdlNv9LlCakkaV4fqzBag3lh+kcyMrEii3Y24ee3rCI/+m27dVARp7Ni14DR/OK
x6Nfmed0BpuCh0Q5M+xfga7Uxknj/X7zkhq4jE2HucsG+JDqqgpSIYiHvewZ1DlRZKFZSenK9zUv
dK0wHOyQLpy5dLWMWQP5PxrtHZegOdgasBMPEfBYkBGXEELIVhvL9P6BUbMRhdwsr4FJrZRFbPDB
+1alPLfJCSG3ThIAAOGymEr4rn4vWk3N9Wo1r+PJ40dxf1BCyPR3pNch2wuc46y72GjaptcczSe7
aI5qthY4ApZ0hMAxydcJ+whwIA7Bl2lOB6u2RwUFjXugLGUkxb8JL1x0nWzkIbKHW6/9wRuH0baT
7bnHXlheDUHqVnmmRPXca7HVvuqqRcB6G2b8kXAzTU2s03T2Fxszcq2HVXbR+xcJgc1ZsRPSrFRe
FAgBgdwqMHXHJyzyrKdJ3G3oxy6CWDkNeeTl4+97VfH80GE+now/faluEHJdo429TdR4v+da4suF
gOiAKohgz3pNCrPCcApF8G6VidQOk+8lq4HXg8mqCAKGZVt/03Q4Z61GeJr/1PXYZLoqd6JFzNVS
YwO5bJeMAVsXjx4TNsz30EvRGEFWXp/2EV1rMCHV/aqL3Lg7xClUcFQ6KHNVKas4jlW1sNfLbqYT
FSDqq9CC+4ZLkOLev69xPchj3NzC5DgBnfDBqaEwYapd3eM3WJUF92rstXOZrTCN0CT0eJab8e5W
xeGsOFxeFeZpeuCfhnYA0JxTEIeDhmp2woY4IIowUFWdtLtJTV+qXOz9GOC2YWFOZZZaCqXBKMW0
7yBlxyszL/CRaxXaNpPSA+VpiGHcL4v8qDHRZ2ZkvaNz6U7qv4Ew9p/jbnHuyZRRKIO21DZsTGci
MSF/ARBSnWnMNl9Ov1Ct3tmvQjnwxTQjvuJaC/KjRMsdfeTvKUTn9oFxUvfyS/xQZ95FsK2bKG9p
bxwhxVyGivlmSfKEuE+lUaol+8ihz7OznmK0hLYIvCqBjg56WBfSAQBALFE0/mDFR2HqxLM0uiVU
QWRwxF+Rbg7ehta3SkgkgOehfMizz/HJR8B0F82NNpD/osOS8cSkfH5ZlRpIhhgrFXzO72HfiYDW
5KABq9BjyJdAscmRX4qAPxhCFqip+zxbSZCupgbVMTG/j+8qsN2jcTfcnxalhuf2tHugThHfpffc
IvRjn2AGJNBBs8HPIBRBSsh3fhx1aA+b61Bpw/loeGx+aYl+dYSCZjsUwV6/kEXkiMPWVPX/aZP8
pRutpY4E27qRQ2tWmY4wXOm6MBLoLo0OF/uABGDiM5emoNAcIBahRWFF+FNfPGVPh/KvA5vd9auS
bVd2jUFvIsl1PI0kMc0nFJ6nmFV4KnPsW/pIVuc7W7WoBpdM2CW40N/7ajiJDoBddv97WNyuih87
HqrZ2bhdcAWZuft9BIn6W9s+X7QPmDrokSfID8hWUbvmk72HBYHodRgd5SwhstRhbECEZ3DHmtFo
70RwPcb7WD+SDrCtuJbTodK4gnBFkkRASv7H/ihoYe9Ykcg/JfWMtlZ1foS80yRDMurkfmnxmItl
0JYL0zPfsnG/iofA0jXAoUaOX/+LGyQGS+pV3+Do8cEa67/h2ZfjFIZ83UaNflT1GBlhGOhqLpno
4nTFVoQnF8Iq/7gy9VhOwfkscSuWdLRE3DISyvrmf0jvY6jLsaUHgkUpFILXeDstHK804INfo573
frySC+a66mPaKj2A6F2KFjKqtnZ0z5Sbk2KZa48Zxy9g6GY1vimFECF5DxD7Ii6T42Wcdz4vL0NQ
wlKxbcWjtBB8VHE8VvD7L14nlMrwtKvflaa8P0W3Oc8N/ft7sH80UkGUzR/DSSjpLXR8hphJFg5P
QS/fRrZKsZjmvH02JHh0q7Vf6o2OK7/aqymy4Zj2K6TY0oI6t89/+1jsjgkxLOZHu2HOuWw3sew/
1xNTAMxl3iuJq4yufxTYpaQqHmxEgEkRyCf560TdbuDwONnWNm/Mwwa2xY542pkI+90nPh8hZ28x
5Bi/Ok6vwV21KMjXIeNYnLaQxfxktTPAi/DZpOk+WeBu24BD3/l4OE70t5XNIhdWnhYso8fk49Rd
5u2r2QBzQj2WXNYvVAWPfOWdNoOymHrfNLg7ni/HNJncXU+IYhcRddKaCyxXYMRQKEGS+gW/zvpc
HihFe2COvBZuzqvBNP+DO8wEHs0k79ZwA8F4ioR+SVgYo5WEXYMn8Td5sZTuE9GVHPkBPa6ms+Gy
65Av9epO06cAtKzWe7eZH2FKFKV2wUNasOsYA1wHo41hLxdu5kL5SLP1XFgf7n7dg+fy9v4EtW1U
+Ko8GaSiQ1vDNa/5FhhrWITP+CZCaSwt/0hT7Redt6DkKYWlzN4sk0WzypZSXy7xPB8VaoJuJmxg
lgeGZakQpdXHDL2YwyAKdcA6fLQSoQyLlRt90FT7QxE1zf2t0LtNbC6+rpmdLiJqtDbW7LgU46+7
dfEWkZQDDMezi1VH/TtpKWWxXkDWRXNIUKanrRIwvVWgta5RfoofLXE0Zc93EHLQv02gY5wEKL+Q
Gbua4i3KVghUpxUMsquc9+ud8kmSXQ7srguuR/kfU9NyR/vWVJd+wFYoRMThoSYtN4gK6JHk4iLm
0L502rkduu5Vtazo6wLFuFyLb1T6QiMuH6r7Uz4Alt5f3wrEt1UBuyaJ6KKjyyljd29vcBeK5Z5+
f3T73ucFYTIFX64/Kwq5lyh522aELTk22eMkFXA4aQhetzkMA6lP1AuNPwHapTVla5EfX2KcmPqd
4FnSGzf01+4BVHb0u70r4mbOncOspvk+yGgSQKtEW+ma7BhFnv7v828rhgJCzWfRTWo30I0DMQBu
tU57HJS5pRe8qwQolvYOw7FRRRJp4zEqUxpmWH1XBdkIeIVzJOweoIri7bjLBc2NZoSxtGdDVfvj
a4LtKAxsRPiKGmINx6yIGI6VivmBHQdlZq9kGN8LthTul+dwPoPMWJb9dQj+YULbvn9LfM4jLB99
DQIK/dU//7Fgmnj/7WSdtvoGsrOiXroBF6eOvfPEyciKci7mAzfaODOs0vK9wMU+uu5RU2WReg67
mxIe3IvMdUESE0h4EfimQ/ZoY7dnsM/xHtAG0PfQ5WKgccr64e/qCbNENZebGBIy1/xkK4mVImHv
3wn/dat63HA1JNEGjoDwiru58GuJ4fMdllvuholyFKjcz92MxHkFStifcHCFlvdKzHcBLvt5qVib
PV/ed1haiUusu3NaZgJPsi7uY5oZQ5z9kNvUtSehtR+Fe7kLl/vTbhCPBxq7JM++oij49SpLOIsM
4aCMhWtYZwMl/JNWxUZXa9SpKheT5wVAqh1FwY1W89k9rNujfwjYG8svMJtcZFroDKnuVwJnBy4T
qUiGSuRC9MLfW0xM+tyjau5gXmpAZWabXIWIvSLJ+4vIN1PBCfi6sxEaSd58RJKNLVTb3Ti92Byv
+4wK3QXlER6D4+Dv+MFASnnLMj5e82WZhMZFN6axw0kc4jvextjx9trDLXYEU/C4jkvWsPRAvj8k
2QHKOfYxuxozudY+4Fn3tSc1RyJqTYDwsmmDT33TDuTJNo6MPFxyzn3O6bZnLR6OVeUMCxoE+/fb
jhnUkmo7/q4Aoi7v52NHCm8P7hQdf1UbR8MFH4czRusbcNSwcs6Z6tjdOfgLywDdAjfxm3yn0eqL
df3nw5YsPRdzvZ+8aPTQdkYQ1wqK+g0xZQ2wBJLwsPSzRasiiiMolN+rQYtAavlPmyBedgHNtg6k
Rqx43/GsEtSzCIYSM7qqcQjaj00piqHY44DA7VXIGDWjRMGf4gGTpilPymorJF2LuoUDSUYVAcD9
kqZ/+4zqyfiQpiKivYouQ8iDliy9TIXa59fYAVekZYmVD40ZZU+vUAQ/MH71j36U2ft7CnaIomC1
U0dLNsjCK709GrOIc6vCKYc0iMDXFUcYR6hUguU2oC2x1bJZEJxzHEuQM1x8vpwL5Uea6W9x5CDO
OKzRwoHxqoM3XaZSupNBu4g6s5uyKWVgeFeUJG/D0tGC7u7su7ABfrb1/ExmHhpMtGTcpbaAB2+V
NFgT0/PcXLqokY8hSeSDE3F6831F79S643ffGcLR4JlIN7rb/5vuRmtGjZlMAaI0TEGItTeJBStV
HLgzaacn1aRtQ9r/MBErvmqzsoZC6cxJEKxkt6xY80Vo7KY2hRdye3hqh3w2o8s50uW94X0a44oL
DtJWGjQs7FGYEN1pZbznMYSjDpbg+JXp/CP4NSxoAdId/KNKMrpIPEAHS/xcSjnUFVZc0zchUAXe
xOZ+JV3DZhdz9TpPID7r5mODGd2pEnLkvAMvswGDrez47VkzDxOBJSR64slr9Bq/fZVpW9Emge9u
7dc/ZqzTG0blVUiGhL2Tlumq3rkwFly1IroDJ4mdcMyV66pjsTPnOaWAFWOjThk/2QWbSErUP/el
aJ+S0rNChG2zvV0/+hexfCaiH0GzP7AT4FVvNtgnqce5jiyVUtwZwXYxCKnC4M5OC4tfba3urplm
qIQLSdG726S/Ijmmk82Nr0u5tBZ/RBfRGrCICz5w9bY3z3YXzLn7mQxREu8FSCykOB1KKO5EpLo7
5iZGgmuXi6T9HK5oGDBOCl/v/MOA4FPFu1Iqhri43EvZbPpaFWqrEukfIo+AoAtHlH48oVUqS2Mf
ykHjLlEnzzM8v0ag0XIxhOUHY4bQngkhyjD/EeW8r7CIS77cz9qbcVBLtZvTJJS6Cc0w4wjoN7KG
IW4nwMeT/6/PyHer/W9PpSEEXEck4ygZ31Cygt2BxiLBUDvod5BQ2OtDZ02j1Xdb3eW5H1Qf3czW
PFwjx9sVK7Ku4whzcTHs0cm4dQxCzPvGdpOmjFeYQR/sLYx4SJWB5sZcwqGtjS5SnwUaN8xbDS4a
X0W03X0kc4qJejfCBfhc5P8+m5CXhEEGCE7nnXrLuWoSgHnOicH1cdm7u1p9OScIg2HDQeouDo2y
RKXIHk8WBnBfeCHOxX2M5H5AwJZAa/7kA7UpQiIMcghw5i8dIHRBYY0GAcVgs57W0451LZBYQmUC
H0RO7bdqCaw9yBc7Sh8Rgl2Tl/yowXKvpybvVE/gCHz337i3XOPugPsRtmkyHb+6DsG4J1Wbw3jM
k75GOR28hqoq5Hd34zlT1re3FvT/xeNaSAq1jh4X1Z6SOtkfRqIHf+LbYpK6kC0dEMAPW2Pt+h5p
8+b4mlqjJ25+nAoMHF8LXzlmeAVVIsG7uFmsMT7YbunA6LWVkMBVbFw5lOjIWExGij48SGn7wk9/
VDJ9sEIG2otKfOyRcsj3/90fvd/5UD5d8miai3xi07bWUqTRaMJFEtg1lPY82FVXa/TKsmE+s4I2
hBAvMe1CokW1n4F8MEfbr4VgToRTPYVECVppaUlYLqUtXt4V7iG8ZOsvTxxZWGOTirSMOAHrHRQf
8vl4dGJEk83zCelbD0KJt83LmVTu/RoMg52Zb1j33+vQiO5NzwnXRpIwQHr/PKZ5AiF+x+lzkINr
HSriuplGrf33Mq9MBN0/aNHSjiUsgGmA98SdRDNisgl8of+P1j6wjAe/H2ueVov0lfWnsG8tsyb3
lnCzoC2xCQTFcJC67OpIAGfLAkppF/Kwc8OdaNFchRKggYstmBvi327tn7gV29j1mJEyuCLDn5ib
D9v3hA/HRGetF90GZeIFy7QhFP7NrY83BrnJ7Ks1p+TaYQkel0fAY+Sm1Yv8WMKM2TUARd1dNJsj
jkQKzyo/Fin7e/lw28lHXvtXnQYeINmh91SlWsVnRH2t9I7R4mAOMmgjiIkLKqhsCAnl0FMKOYGl
/aA5JtUfbMnoshVpwD4ag+7igsNL8PjOcTkZ5okWdTCngusNMekjes8REtrx8RB6Bkw+hV8RFA4Z
pfnZduwMxPicuA4aycVWD/zgQ8anBbP/NueGwP2eN+Baz4s0P0UYfJL4tDumip6WFzsVJVEzouVd
Tz/xWrpdXAOjR5psrHqyYN5n586+ymzmrtXitoi8H8I2MFNd9Fos5oO+F+NT2fqSYw9nBHplFxNO
nvWoKv1qwRQDSDbbUGNJPK6hUnQNL1qdXeQfIKJVN1pcV+xOwiHm1n5mDIgc2CePoBgFB2eJlGNY
DjLnraarkLARcrHdFfb+nTCSQqFTWHx3vnMvEFQ9tJlUzDaTJmoIiN3//eAZwtJIfQq9gUQAFjkl
gyWnHOZl6widDQF0lWKcUqzHeKxDpea5rpZRWMflrrUHOk9y4P7op102zVlb/Q3qkmzeHnEGz+Ry
j42FZyiWJmYjkH6bLlz8OZsxdI7dracvtL3x5hMizgj/LK5VQtctCYVdlJYO3Ob18FDyvFHp4rR1
WTqXcYzYSR+U7pgc9P1al3/p34wGUayee4D1/xDqMkfhiiSFqsfWZ6QF9nCPWULQoOdIoAPofOsZ
xqZi/HhTrmEFw5GWl4g8g/aSEbmZHOkO8D4exM4fcNyhufaXcXKGJaPlImlPBZurNfHNLdqPxYvv
QPuMg3dxtHliQVs9zUXyvpK5CfQRVPLamXP56incnrB69QS9ZPDW+yn4j0PCMhILk/heVNNhl0zD
PWdVfbSHlXsRUrEVp6+npqsvnHNwvO62FMfJKK85IiTd8rHFBWmAahlhAp9iDygDz8WqxRqKtWCO
ansWdtP8vzvvxBG1WUlogzz8IW9BvXLy1hYA734CaXuuLws95wwLa7f0oBaqphiL0WgLTfwivW4o
Bf6r1p3K1fInDiW2INhfodwjahN+jZ/8z6mGqVlCMiACuR7uFR0vC3WUNVe6fPKZqZDxvuYRqXYY
UInuiYe40iubuFO9BaDFDT/XsDT7blsxC8kC84TrivWFJjqYuckla+v4UMJZVRLF78I4ARwZhCTH
zAmYUkyyWZayaLWwioZHvRBxuSRsJVe5twNGEQcEAdTU9pWmvyj3wsL8g8s3/4h6fvf5T3n62u3k
1VR4jdVPQwmFVfXssCf0XDIj0BJAEp+Kxwe5VnvxHM529aCahwko8nUd9nzcjtPNhKYrmGXfB1O1
ze714VAZ9IiNKKlNdGqtg207gUHxYBn31nl76U3TdNJNsXpisPHil5tYqtqjbUvKuNdlqoAU59de
p2RZ0dZE7KUcdf2jpDc7A/C2p82TulvHIsHYiLijvyzInPHh0mI5jsy/MvTmhmCp1N2v97aR8y2C
tA/2D0HDDQXEK2Nkq9f2cSLvZgj63fdoEvte9X4Vf/+HG23orf0OmDO1u4oQL/v6STItRIK7RNSe
gLQsbqLEsv3X6KKpHNqZcN302erx9r/1Wta/bZVBf2yh4UOULeX8mhF3cGumv7haku0H7XCmNMr/
EYjaxJGQGXpmR3Wsq12FkHefZyDRJ6RjBxnwxtLJDjD1YuD8cpTMOA69dZLyY6eO9MWQj4umh5HJ
oIIcztLHOIKzX7KyUvQxY79jwqLeimJnbRz5xF12zz0elHI15al343tYp/xRtfnztldp270Pa6Tj
viHNE/v2FnAqGUHmMnykM4WomSQKqsI2RR/ZZWG6UTIrTstRptP1/9+3elZM5qjCTcr2hNj6yxrE
rEay4QfOzhDtU4enUKhd7E3nlGISTQyxYzBD/2sL3ghneAi7mDOHhIo5uL0azfrHYHp3yFVT1oE9
/ITdhBxkAPppqWbjfGBF8IGesZeY2hCqSkqwYnKZpmkOhBEBMqm3LYTdU8i957YEmjpHYWsAPCGn
TJs7T2Jvzo7PUAYU/KKfjIe8BoLfB1C0NtVcdkNZNswFIcOVZ9tsH/suwMIynatzhOMMM9RofPlb
jFCBeaPOVPAB4oK5u91cqbW9bPaUqVXxlBYeFMMZywBpd0v3Om8JuZb4QfaLXgNrOQqz7+pxEJjP
iiNU4sS9sKDXpV7BNoQICjYEYcbA+BC81a2ROO9mjlZ/Wdg4MSk16OpR5/FeXSL6TTHBI+u9BhB1
zpFh/8RCrhjG5QjBuvnbxmwgm/Co3d1/hhqnSUnG+lVSjIpQMMcM5AfX/96uBP8IpZiFeIGdxpNZ
VQIb9UpROTF3WJ/XFQSZkPCdRPejzgSEVMLE9BF0GfWyPNFCp23EwjWGDS2Ajh6VwkF822ckfjPe
MC0VoO8Xq5oQ0yXTRqKrIDMN3myqKZMwoCZ0S7gBuOtEs3KEc4aX61XjQPeFC4bEfJY1FRUIMGRh
4EZgiP3+vZfU8bPe31PLNpldYpDruKbgzKxl3svMkJK2161tKRCFDYJiahHzxGDnMo4zXkX4uosL
rgQaB2rZlRm8JR3XxShUyuE8pSaVQ5EKd+SCbTcks4OXMWxlROuAHtuczNZbGYD7QCQJIm3kdhvQ
+nbsFfl70DrkVtkeZZPaB/xJTO+/tdIy3yUHg0zSOD5u70WlQKNfZJKR7K4QqFBJ0MybqGQHBNh0
EhDkG7iWcH++6D9miFqtK2Iw+78WPerZimXSQ4TRPk0ZONHwmvlIR2imHhgb2lH1zed8Xs/zDrYu
p1C10J1owWejTwlYfZEaa0++5mgqCXeoHjc+dNzhP3ADZ6t9zHyhHU6SELDbolq03DPDNe/Jxj3Z
E2GcHNiTfIVbO6Nh/dPepegzTLabR358W8PvnZh2cteBxhNK1Awg1GiM00OhsnPZPnC6/manGYQo
/+kfKhdoE+BwdTM+/mFE/htpXYMzb+5zt0Xk6rxKcmOD9uaBSvrHaMALc4U2Q53G9N7rqt+cN7de
d85X48RThBl2kkxYGMp/6epJaMy2QwrF5R+VrF6j3CTvHghSZ96+Gji07Uadg8h+Ao60jjwkypz1
DAa+HcaiwE9UMl0eTPz67SFZ/EMOjqvNiw0gWpUpZfVlKXmtxG5ZqH/vnLkfSfdE74UKuKbtgrFo
UuLwt9ePkIxx7+RVRXyPaSEv6VL65q4x7rcyk1omg3s3kooqz6GiceTdFetwKWLqbDuzgoyGUPLs
+fWnB/UkxSVOAgNgqpZiMZiSEyiCgdgsTInSyFuUmTLk5JLC2PxeMWbHKRufvDILfbgK+s8Pnq3n
QdCSwFz8JfLCqBgUHOcvkO04bj5f/1AedFk3jcQZIjlziHvVuStWnPizpQ0qmGKPFskCgnNsQvOj
YvAI5YVSwJlmHwrhTRoIgY7dbbtWb/vmjHlWI3mE+qgYiVS6kd1WzD8ZnqX38aPNPw7Tch7+th3t
CHukjloseYxKSZqWEPGoInZ/LJLCBGw5KbNca3dWzb5+6qYoxJ0ocZzC1E2gK0S8QWbNf15PxuaT
vo0Uz0JHjubbUug4RjEwBKAu4OPTGklf3Quja/uGJtXpIaRyWnqpD/749w4D53Zya7YZBxtd1113
+PLFn+MlYA0c6nmIR84RJCeswRgewaY6vgG3xGmYeyEwB7JdJdou437qn9QizJXUwEjemDXlS57V
xKjjY0edyoUXIHF/mQwMyOi/ZjF8G6C43/FfePZk+ID+dBbIjuLiM+wYcvJVXT3rTU85x/dn5mbz
zyYdKoBW4ibH9+mggdbOnKIhwneilINpUbHb6d+SK7M8Jx4H8iJnEQixNkFPlcb4ocs0vby5eUOE
E4O+SgdLI7in+VigvgN8Uxwpawa/xyAhwqiZjejFfxzsRRGY/t3nJQ6To0jPzUCWbbUBgYDexyZf
iedWiMT4CTdpogi8nfcAjafhMOCxH5kNuR6fMaR+8S43uj3yfpKdZbVvkQXJocEP2ZFTgB1UqMkf
8eu6wWEq7zTXv+FVdHj+FLe7GnBb61ivaISXMFKnwFceowqiRv76WNKE9fEauvAtHRnjyvRcWY0L
eoojpVO0diWNtOAXOxBuxNBS0SdfTKF9/fTx9mJPXlk0YxDGjPCETHOz5yoaOxqyara0GXVnVUJ+
MFNShofRtFTmn+Ji46qGvfhZwWBb621gTIfNCPiWnLSnTFM8DMWo1FHzlHcah/0R5PElFoHo42/O
wITOwbm+h/Az8pDB+hNZKGYgSLhF7QEpneu6e15hb6Yxtrw53ooawS2gygff98iOCcRYa83L6r1u
PamDTFjPU0DkgPj6FPxolhYOaBlVcQNqHe4UnMTlO1PI0U2VRsieFJ2jmHX3KwO5yW/YSQNuGM68
vV0Sn6yVwkuBgOi9QgT7Hw0E43pxpR7oBZr8vB1Wl64CSyxWzfK5LDsELR2nDSChVpTd2EWjFpod
eN9f4QIgYe8uu7kWmvEJ/c+zcd5pK2URkFk8EMYqIAFFWXr8Ua8SRbP0nAB30e3rss8gLcs4192A
YSL5dxGK0q9OArM5TvHZZRaFgupsr527AzyC4onwCQdZZQY3AmTY5y225Q43DoqdXBZoi0rfBN2T
5m9oPIWkbQ2rSweduUJEWXAl/trsHJJoi3zzqTzUK0iZlaXy34fCsVJIqSLCcCUiArZciM7YS1b0
LTy6knppVEXENgpNH0PAcIBcTQNQrESqisGpIWgbFLpPzHBFVYKvsWAz9+b6eQXUzFYHSmqkkL+s
Iq8FhExIkAs8MFT/oBjcd64xBAO0mzgsvaWok2ZRH4HdJ3YU+mlIW+TGBsTeWDlcRQQO28YnXl9C
jOWTosgho3H0yhMRSXTLaPNrXrtYMVPKat4pHH+lPrYVajEEXuxYV1dUbql0wRKxhq1inZsob6Ex
0jDpsBLDqOalQzPjt3StSmvDKPaWDGGZsImkYHUqBto7dwRwwU2HwzJWRduOj4cloD574gRVw+Bg
dIH/a/PwoDXPJlELJeYY31rul8U4UfHB55Cl/msrq0D+31mvKN9Fv2/t30NiCE69L5pkmlLLIeUq
KKG4GnFYXBg5NQRmnSPK7Gog4FAHCVYZtQyTvT/ZZLPcrPFZ9jTt9e5MgYF0hcElL+ipwTLiLfMc
Le6UYbPLReqWbwsAgwxap1vGFMxQUXNkxNFx+UNmjCE+esUFKTXF/2GdZRc23EDFJPrTUJ+D0tw5
FdxDe9YouEEpmtIFVaHdJc8P+nE9XECU5mrKs6o5ML4zkC8am1ZEl9QWYLvyY9PgcwFZ2Q8/G55R
dbGZCSTmG7ABfcOJIS0YtN++qZNXmxDJwWPzWPqf7+5HVUu7Kjhc+DOdYQPm0+IaeQct5mJVIoqL
DtcaX8l+DD5o/TWx3Vg2BG9NZkuw4AvT+y6li1uwdHKdFaM6BPY7i8qeaHGtuE670ERO6PdNIgb2
ph12yuSi7VDTJlnMr+ADFHmxiK3qLPQ7QW7K/wUMQIuGgVl73rZ3sA0YjcDn7GGK5LIiXlGcPsHV
O3gfDl7WFtiAUl05PIr7kJPOQ9l6Fzis8WC2nNRuBI0IgRD68LOhWQy1suNR/nOtEhSG1g/BOWhS
/Yyc+UV4Bq/8JjhUiM7jJ4FW7yTDccUu5o9Qg2Ckok+31217hmf65VvW8Ej2y7h0GSTGwQbf+JAX
SQ/lAhXJ7tKlJlR0MDB9qcOUbgmjFIyHtThWHB/POHfxrrfJzuWAJ0Dq0LanfZQBSUVX0N58ze0r
swXfyO2hZ94w1kj/AU5ZPjKddaee5wwh2+mK3rtSX+HXwoMyGCrt3owi2g/ySzpQO0dk81NRPIFs
dxBgmmxK2Pk6SbVWaSheqcZYSmEiHi/eWIKObheFI4v57HUMGuQcqyepNqLaVYmR1yuKJ0aKr88v
fXkW2VDWdEkeHw3KWMv2Lf2OTC5aMKM7LhHSFFNCjWPXqpdibVjV7pc5DFnkMeom16CRo+16R5Fg
//c7GA5LZsmkCcmsKgu2fKU4qCEACRIhf/ujlB5V3KlYZJlBwIftUCPC0n3hvHpVKdBQ5bHE8zAi
KNwdfFrbNZI7hFQ8xlFEwCsIKu+LFDPvCBS11wAPc0XdyormX3ryEZ4ueBmxax39xbYeKLOtEefC
4vS5prjXKmFfiaaMQFz9PyyvUJqvK4JZ3LHDnYWS97SbNbJcYvxp1TRMHnqPMWHixjqov2O+h6nw
qVj3QzZdUYyEpcFPIwMoPz/FJj8Fyb1eWGkR9MsURHqSWri9YM+FvbvO/G/D+A+VLgEw93r2h4/3
asDVVz5kRDCuHlHJJJfbqIiPZtW5+Iql53Qb/nPpIjHuCqsmMCaDWhm2ShxC2DB83Dx10PMprkBR
1rtWGMKRBhAqgrbRtw6942nAfe0SfRgIkZyomqGC4DPiEhXCh8WJMyMz668pUyOnsOxANm4w1EN+
KQi5Is90gpMhe1Tphl+GpeJw6HyHINbphyUceYOWvugCRj4o69OHS22wX+Ii085HD6DYQ+Ak6XzQ
vD7Mm/eEHRnylj/0OH5/K8hQvZ4Vnfx751UlQz61aJulOE4l8mjkwwJCG9IJWbD8ZSxWFStp8i3z
W41VovML2PnHtJvtfQk4n3xV4E7HpnjqSbh81mUjqEvrYoBtdcmaprNa+qM/hAef8XrVhrOw9OvC
qxtDQmKDj8EikuMqmKkIlUgIvsn4GsMy+/hwvJ2Fb51YZIV+C6jHw0+S/nRAbCXIJeMHWXlk3SBa
6gm5iG1MHf/1HGmrkW0w9eUaqUb8QkkS6B7M0WhoUHaFKPgqb5B46sQtbGTNJeCG+46yf1UJoWs9
xTNwbIeRxwlAKMZLgWkfZga5qf3AaGHl1rkxNj61LrNS1Veu+CksJsRLkTfygoZLrpbC/aJCKM+0
hTmE76F/SFj1i+aZI5Fki9qzriqNVurXSKZUdBXZ3f0B0oMk64FXeqMwOA3HPpp4wVlRdO+Bv3vF
AuQhi04IB5QNnlHkE1nauNOZlfB5G4Ou3ttPkTJYR1eYeq2jKXFfixlrQXQsodNuMDyUgMxuX8co
RlhvCyrgnyIBy9KQ6WXEnJ9F/d1jA/KtQ/1xSBHPyUriQkMfXzKYOZ4GAAM9g3U9jopcOKtfuWSN
VUrZinoZmR9KKOAXGWDKX8VgXwijfRv/EaLWMNG6HKF9tteXxMm5tOYi8oTOfMQOlW542s0qB3it
bGP42gw15kPwisyvOsRF+vj5WXrCpIOBPf/9REFjA4gl1yEgOJW+t1vgV/XF2FzExIkuZM2xm5bp
MfqRXhBHMMxhCazfiWyun8ErPnm0FGOxf2x0PeHxmBWj8CJtpfHmIC4bQjLL7elIjYZf6IIzMo1i
9lb83UQ9W49YIa9ajbpvBj9B49undidSM/KbBEAmS5HnrS7mztYM0/HEbmg5sUjB3kBVcTKsHtCG
ehK7xdv6vgLM4RYIighdDVVE5t9X/lpRDl0Je6wcuYHeB4mNJjfqHda02nwiqSx+aS2QNP4Im8aP
Yy1VAt5g22Cc5qQhaKvXo14Q/VckzICPsD7akNAOYFTCLwnHiYGsVD9ApaH5YtxE1sxYowxvBHQG
rvaIwnn44iUuQmnlDKXdXaQxfSM5ezTdQWiWWvf6V7oKZo2nL+lL8xRE25NQly7bHIkaBFwQn0SO
RP7KOO0/vBsYwYX/L33H+YcWLNCjAXew22zFTW2+JEIa5FlLCA86gia8PrBx/BrPe2sitWgE1grQ
+/wwsTQQoMPV1/zODsDArwClTWBfFfWkjmLRQXOg41CwjB+Kn33DPmNFhynf00gmIprh+DxRin4O
8Xdwz8FxC7UjCLyGyt5DoIH0QuZfn6cYSmq8K57Si0JRULpCoA8nkd6Rr4f0wxciQVt+dPpkmga5
KUdbuIL+nqIQKvhyDfpAztfGpi4bbGAPGQNBbjYFZWywf6Qh4z/FqmL2pQX44PD/dhx/E0mSwSlc
2eqOdG8LYok1oEMGPslsyuHyjUUaugz9YncEWvluT6qjB+9GVLKnDUnBXa2GFg+qEu/8dip7Kbbs
Cp5O7vQFWm3VhBcoc1G6XJOJcUD8AunkVsHbMpdUEMwKWfSIeI+qMO7f1Er9JU7wiX0lv3KZVfux
tIej8/jG2z+XpjOXuSx+gNwvckCB4gZ/ocSaWCiEEI5Mn091UfY+Kfhi7I4hqt0INsg/1NWOTt6n
vnLDH4P4r4csIP2IITF1K/RjdptaMP2qm76Bw3pSKD6IMmpxWivHBMoFvQiTEcbc6hyuoGhRa/GP
mscwDO8XcUiBwOcg6jns66AAnH8Mjgi5blztBDIAGPYXT3boCMeWcHk39b6if29gVWIsQC7sIRwL
Lr1urd15xGOil0rpxUwkYXCTBTDnR0iKM8CdmpACTHByVhIQZ5bq5I4ra0l7J0a0EOFmIhHs7sTI
jIp5IRZcQtbuuBHdnoUhpjW7nIvzdVKs4ZMoPf/HXw7r5fTxaLpXo/KWtDRiazTih046dJtHrLyk
YG/gGHe9MlF6aRwuoSOSXyz2gAjKNAzxAnyw5pPji2d835Fa12saiiL2U+JKP6aF/OEfM8emvcGV
R2JYx2PECI7UcD2Rjo4t85HtmkZ/YxyZhsd+mMZOif2nep5DtBrVyXpNHGO+pQQi9KvcHkBX4tT+
AmsLcr+r1cK6YfypemeaBf9VbkXlDZ3Y0xZqi2O6z3YgSrgrvgb0KzRS8FSZ2VjigW0r8T0sE6n/
BBeXwaRjYsICwB6q18Td2rY99IJ+eP0asy500ab5MnXHv0TJ25eTUe6NTaXepX/GLh7TeoEpuML3
rBoad1yKFmbATPb9ADm/OitW6ufP2S2y9ZBq2ud/5NzwFfNGUAgJQcnjFql/kHLbL8z7DgCZ1ueN
Tvl5D1Ioy3SSqQK06STPhV06weqtCaV56A+v/MNIcIe9qWpIuX3+PFw/0N4HXz7e8Q2WJSbXL5FB
a6lOxffXkjzMuO+sfXm4jT0YjkoRMecIt8WJ2HeTBSVlLowLAXHIE+wx/irfXiBbiZOXDHZ4Y9jK
Pqqr6WjA7I6Ah6zK9MEi3QPYzKDLl0CWALNdAymcrldjDfZqGmKFwUDgqXNRut4sV/LKHXTq4ddS
1eHouNm6mM8WSRth1D2LW6S6gCy/DIJMnYJ9Ea2PQkXx2p5ixIT2DWWxN9dswVivrd8ukYuFLCCA
mcUmL2P+Fh292t2qd3iSeH81ow3jqOP3l6ZDITGbvM2b41XNXn7eXn1rLqaGJpmDwVMJ75XOYYC6
omqjSN93NVSWI/D+gvaE5PSoItAzGTHpeAG/GTmBPAJIdER6uoxpTFVpg3TLFtSVn2XlUMcsMAM4
NzCbv7b0NmrK/H7fBEHRxMS2FWD9u8/4IyTaAOg97SWOTG9IoOXqMyZBxCmz9RkSHfzodfuhovB0
aEpi/7YLQuU5nn67De3BaJqj10lRUh9JLqAx6zbAnPOLZjyfiDyQhMbFl0RFysFTVQ3mZlwJFuga
XBnlA2633lLeUpOXTXIBeAMbE0dtvJgYTZy4rv36sKgVjaMkVIHZh2nRaNwrlrD2d6ixpr5Zw0Mn
FIF1GhCvzvQiM6IuZw8Lv0cWchSXujghLtP57nLDEOFAXkUAWf11zPNQPOXQTeuRX/Z46B9AgGpk
bDaSCQL//Tiqdhqe0AH5O78QhyHpNfd3HlTDtkuBWFWw7JjKFjF1RIPsS5Iu+ADHTICTdhdLzyhn
WR0KOUTILILJsgsrsstkyQ/AsTAjjJ936BV9uDPTN0oqLF8c06tROLSe1gEJ8lRl0TsCSdWmSwit
l0BTE7mThX1uO1t8gn2PRE27JmaFWSEiwYL7pc6yNRtcU+1iDceuxSuB7jdVZDJXYm8A20pREmMs
jIsZdIVLhPpM5MhD3kzAploBY7JnNX+j5V8B3pPlgnfVXDI0K754oMaxTLZDZGP2zlOOuWJc5yUk
39umQoQY+efguqvYEw5sYlCKiC0FHM2GKrFI1IMxVcU3kW12ZQsgY3Mfdlo+T76fWMzgxNTiRAaG
umHc0UdlP0wSjGjW5d+AvSOO1Upc/6Y6psErlt4c8bhwpXeYH6byljKSGndkNOpBnMp1PrNIiylP
GgsmCoeyXS4xfy2AJ1mQKZjX96QAmMN4C5IjES1/5WpskNoGiAern4vMKzd0vtyxx5SoZkwEYbJE
JgnqK70x0w6n7F6octC0Re2es8k2OJry+s+GV52x+br/fccsVRlfOXA5tIZ4ahyLWcbKp+Zxytde
P7n7PbkLWfm8/BJO4dIOeo0QR8VSPJIhwbA3Vcu/c1nCxxUhR3TGOW2YIDgkUp/L0kJUFlDQWX6F
kgD5KeYSBI7dwhmeaM1psJxPUYWA0qXsvgl8CxRrY2BEqLku8tLdmfSmxH0moYXelDP0hz/KKB3/
ABJvSaybIx3kq5fxsIypL3jFDuSmqydmljdWJgHCqqjsAiibo8DWFohAlLLvwohULLVuGZefKnW5
vXjeYyLI/3q2DtzncDf4WHkvPDSC826QGEZhDvSrRzgs9hehxu6RVmyPniodeZJ3jkWM+FpZumjs
pOqXW+tFOWjwBUYW3dcWQVR/OCckStUP4KmUKuaW6nEi4QY5A0lZIOWN4rUSuoM91vTA08xbxHFP
rBAEh819RqxHp23/cHvHnECTPakTMa3wXEIzWPqFTpsf3TliHyAhTXzn1RkCT8z3EQNawv5aOnBV
yUODE6oDE9fqAslBCE3lU6qnjrtRNEzk7jlQmHLm4oIJ4F6vvIcHKuQiSUFqHdqF0K/6tfLEr31c
POcYY4DBxg/qiAn2cYxMHPbaEtfOcxGz1NPpp5bLHMwF/uR50IoUP9t4rsbT3U12choGcrTDtQwv
JY4CTemf92Uu71RmF+D8iLqeu52gTMWKjvLG1218b4Pxs+jsemW3nio1I3bZ01qjC3otM8UT29pN
fgxeovbhXuPdfLNEwG3eiU79dOZidaw8/yKI+IueHIyTCuj7UYQBuPM113teD1rpan7iot+izy5t
nTP/uGPIFvBwNpjlK1SGyU3ER+TuCcGlZXDk/w/7OdQyZlHzbpHg2vvlKRHCnqNgDX+4szM294dn
WaF31HSsm6O10O6Exc3XgPJ1l1EvPh4HrrWiQjivUEyEACMyMHIu70xGdTbkpPh9U7J1fwxQy1zA
wv4wQ1UaCcRokUSBMBIULP3zFsqKNgEjK0bjB+b27mLY2aE6+lgiAEV7qZ6TrA3Um98AzD1d77SL
hDh8XfT3YgU2i/09OH2NYPWoi7zhyc0zctD1zmJWp6rJffg34Wzm7w9CMbqgqYswVI/0P/bECXmK
dOwfZDsgNuLkbnRTZ4BhpQwuuBTkYqaIryqc9/YfbU5h+ASt7gbOenlzWptZGvYRvInXRaDItQD0
dBa0vehHcPAfjNc2Om9yn6ipBQd6Izs0OjKqzVYz49jvritzuGpNA5QF/t9Hm/pGLp02SS1LIVVg
QsmsCVTsGvnKkM6FILExsnsMN621CuZA8TevWvK8KkHbmz6SIGP39tvtE4SHAhAVpC+VYK2L4k34
T1fX4mubEfrjbVZT45h6kXFhVI/OzYNHQvQKI12xy2k5SJgvCj8/bxSmG48+oLcaciFGfrdIqvf2
3jBhyptgrhWSbKvIdu8Skth/D9fOK/P4qzDyxTrSBe/6fq/YFLQcA0bmcLPh8zGK3EnfGgL7D0sN
BVrj0aGLCsmTidK+qdhkGAjsSwnBIyjBbfBpIJ7MOcl1KpJIj0f7u9gBklOriPdaovqTeOmsHQWw
6Fd79Ord/BqKYdPSR/b8wbnx0uPt68c+bHS93H3xHsSmIJjyRV5kEM8jWgrOwJZMNJEW/sOP7fin
JLhDVhWLdBxRgioxx1o8317sZVOX2ieEKALGzIW3gk/CeT7v14wHRqzQOYmYDO7RkYJ4v+DXAETY
cTKscKM5o+EKaf78l+n5YuRw/aOWsHQjYCQfb1ZspqQ8iEdUVZuxhQALnuGC9JmVXUsOZ8jB+idK
6EVOPjAw07S4e3yjgrvggOyrOy6IQd+2VkM6AfVg+mzoxKcJxlzCPecxkrpKBqsEnVJVUe3TIs4e
A1DRiF0qi1wMr66eTj/X+FhzvlyQCmaY1DOOvx+8DsG1KvuE0clNvN6KYDDLzVxNeCCdl9lea3nI
vEhpDQePxZrlRSDugYF5h2ndchxoer9kkcEz7mDb6R4XnkZmjC7drzueJhCpy2YRMcRSHe1wIu6W
d/o2vzuZl1czsnRz/0ZeQYSDXPs6sdMItzEMp9fJ4by4XjGm/prKo31s3ZQNvU7c3WdQQ3Hdxu5y
lJcvLzS2ATWKcqpMMGNeXp/GMt2wTqSsbKBo2Lii7KjK66Mz8j5IIDcoHv3S+hVgN8KoVYBNQaGB
NNZy7svDhB9UBCTGcLw57xcPN047/cPN4du0IZHquBrYD4BLEUnxsaekdg+36daRpBLrGRa7/GAH
eaAjcz8+HloLz0SnkyR0WnKLWbM4V/21uFoZilM3uF2ohPpRoLtafwiBTzPBi9xfwKBDs4qdXjnD
ZDkNtSnfL4ZEQ5EX3yIK6aKaQ3XhhpiCpGiN9bUKClTjX94TBj46EfnU2PUB+eGlulYmhk3wtQ4h
T9RxnJJ3TUI6B6N6kfdCZTBGWFOEBZKKuKXNgYIiJnBF9qAg8dWPzr40r1ottK/fiyGwMFUtP8nR
z4N9Kh7u/iIqSdXEte7T0WqW4fRLX9moTQad+HPTMuTjaQn6fbSAdDh7O+B3no90taZ+rucybxB2
I8bworaNUmruXM+6fGzMb9Q5506AcxOl5CbA0BiSftbAb4XzID9f7NXQBc6Lk5r/A+g8sAqGn2/p
n1RSvyzpUSbGeRwagfxiVaQKJQAtDz7DzwUsP1yu3IsYnbDn9RKaI5jCWaSPvoVzI53KCu5HbYyQ
2oTUKI1HGGQxLHpetIq2n+74AGU756GEQZf5yKeLb4kzjcboJpHs7y9SaGdoLJAZdUkcX9O2QkQP
FPmV/ZCfsVZlOHFZ00O9+dG2CtwZYKlzz1lPLnVCuwZY4a0ly5L6owOp53UpFGBTJpBJ7HtbvB7u
+pVOTSHRQ8BVeXNNYSnksoDIdRVYlWVWyxZDl6Mk/zeOES3EsD2jFd3SDZbuZmIbpgf39NqVS5tD
fQQVtNZFIPztIPMyrL8DxTTcVIMA5vp0ZDYqhl9K3XzAYkxtWQr/DH0u3XQV1BYBBoxapAsFq0VZ
MZ9mn7p1Bj0lrHxTzY+hccrugREQev1zcprrsowoHhoS/JqH4TqB0ZJwzz8lHkCqSKIMbCZSDrSc
+oqjVlPCP/9+r43PoO343P5xlTJlFQ8BUVCvLpMj1C18/fFrM7+GAYksockf6qOve8ZLxVPAnn23
Dqabojty8lOvyqz28nTMYhRIjrw+r5U9d/oavMwLsYfAG1TaQ8S5rIWL4V7wYLXFThZiDKEY/7ev
kPutu66tCeTqqGx/6XAgV/Ox7Z0ZL4iyI1VzMN/kdYpxGWCjKFyPRGu2XdnLJ90T1ICuCdMRYHDf
is5rKtg8fle+cjTyCFgpPauTPnUffl2X9+NvBFJXlzTogtftlF20xx26NDzamL6FQnmNqHFXYEtV
jJx/mNQVQsB5C93XcFPvfnDGeoYY2+V64MdAJj8SNEyEzjUe8MIVN6KckpNrA7oiPFfxsO/1La34
mifV4qZ+RaNAbMoBhCcDbmbRPDLW9mZM2tFJQrkyRg2RDWZrs8HmwW3TxkU5WdCufvlcWmsPEiVy
5CvT6gcUpbB57e6GZcMeD7R0waJmPt417mDMMBVcoTSUeXoHTNz73KwGqv4mfYLLa7Pe3sjS4aYg
NRBhpdb0b2TY+SrybzGmigMeMBPSVwbgBWFxFyuz22F1UqEGL0Ab/NXeVaVvsx7c8LIb8UwSrXji
QCYkeN+0lX6Dm/QKw/TclS/MdTJqQZ5ffpd2Est4N6bT92/q+f/cVBWVqQTgC3RxlSpPeyeyIiSX
DkxzFHlpTia7SK5CU4kA3dMoCsy24hSeo6b1Fnm/A3z1318GZJrHP18lUas7DLfBQf5kVHof1DNo
UYEvyeMZxWxCksyd4C2bpSBm91Fzuzvr/lXkYAlPAZGiF93Lbx/9AUPsp2QbFhjGBJtyh5odArCy
U2uMzPo/3AM1qKS2xVWCno7aWH8lk8Z91WKYy0/R8y9WmyMoG6nSTmdSrOpNEluf/iydeN9SWAS8
/VgD1IHdstpHat8HUFyza9HHTHMxDu8991/NAUVW8W1OwH0MQnmwcYwWgsSf8H8W1xm1iTfsDpMv
oHIoPfwk64nO8OHlLYOu1/0Rae0u+Bpv02/sIcMdXCTmnXl74aFIyTMfEAFdoCmSx4eUXjAxXR0Z
nKzGyzEChrZt7yvyPqxsX0ilOK7tTNSe/0s5t1dstSbo6ED/Aemau3HA9aNoWtM5rF1mGZhUgr7D
0MAD1e8ESd5BaZo4q6466HVd+8sFaxYVuyexOxeqMh26sKKPbkcSrMfsKucC/xsQsoz1Ge7vuSOL
Ge/cIAjwK+T3f4a/dxQNB6W/JA7jyhSKqLF4ZdrB8lWxPvmI540FPccSSpsFh8/20kFJEG4FDxFw
mqpHOKGoffgjulQg44O6ao3R4w036GRpQ9dh+lKtZ/MuxjVzUCSAnqHG3qGZJ4SO6vfUcNSNI78m
Ym7CxriMlPL6VpNfLa5YqDbLbzJKkxKFbBQlHZrG7KhhkjCsaUgwuqpjUdEn0Cko7q2azUx8tWxb
5XlKdykCdNk/5bF54nqsR9OLGeSXAEW1jQQQeq8DQ2QbT46V+JCdHvV8FibRyAbcQs8ooD2EDn50
aRJqZbFOyyLuKFIgiUhgoasRJz/i4gb8NAMtS+7TLjSh1YZIoUew9qsKTEyGClZVqQekwdZOSKvI
gEKdkLTQfcMzd94w+1KAUK2ZxJOCiLtydMXMDIbwkxw8AyXXgUrBjimId60OCFV4Wi7FxiMKxzH8
ZP4xYIrPUCry2VoFl3A6++tgeRnL/k/W7HnZvNQqrLyWgyqvnGr86iX493K4Bv2mSfYlumxDKUwV
GoM85uBi9h54YRZmwD24IvZ9a/rrhZu0+jj7O7R4YxUrnnInT7HBDrDnixswhlFh6RT/RsXnsRZo
TdtKgdJta1T1biObg92u3n+Cx61PtXTQUM4soUXr0/VkE/WCYssI+xH0fyPaxM7KPPEBO2r8FDNU
1bpu7oxv4pjXAcON0JIMDSGee/9W0TnimxuGK8Sz+IucP5ibtJ1gBd7urXN3r2rVy6jhHmxAL7Ef
KqJwS6dFaRVdWkvWbnTvKtY7F6L5vc1j7+CFz3jb3A8vzQPrwkHqVA5Maq5Rs+Qu+2CmMNE0xhvN
V1zPv/90vtGpri31bRJYnBbWRuQtoMuMgZmWpmDX6xAgTPEPk50AXjAKInvJvIBO7pRySaIYUnMB
+v/ryEkTTMXtn4gCmL8c+It5CN2586cHwmnkTkRtC4JRttWoANfWtODTMKMlrdnwrLSnYjAnzcBh
jAnjn+zeAly76gbB8wHU3f6F4wYJ+h0spJvkB3LcQytctoWKD6YkCSovfu4DBqYOK9Fx8PeW3wrY
rOqPYqO3qJUZmRvKY/NTOcxX/pQdSmIz6AiXS0e7+p/U8WHAw04HNlTVUWAUlSMmAF9aH7fUy/og
qeG2rg+WlYI/8KW6kG1fLujAdIjRCo65Rsf3lzA7Zmg27YtTR7xg7nTNVVg3cClxZaNLoZYOvt1q
09YsAQP218Gu7MbF7O276u5XeqlIvqOavpibt/QEAPS3jTNwCoF3z5I+g+vgegayijbAAVLpzcfz
YwuGRsismI20UvSbFwiViNlvFEeIgz+JKhK4o6SA6/bDYeyq5HCUMfXD4U1u78e0iXHX0W6iKoog
gUc7dgu9yho1kEMQnlOCCC7qxgnSEsXUf6BvAiwLMR3B+09vyOj2XxlkzKKU/icXRwnxdrjsG56E
5YykUICYFqxxXwC8UfFtTJAhT2aqVBkZ0oPD/KbGD2TlYQDLHhb7b+fPavR8XbnEW/OyVpvus2gu
KJqFEVi+6RSOgexg/+gxMjgGQ8hC+a9C5mXXF1Z+/N5Hge4mo+r0zvq12jOpGXgk1/+JRFawlOyh
V4d7gJ24lS41c04tTtPWpWkN8YdAqJPzK03HXo0T+vhuhO/OZvfRZJFZivSrMB+g6QlZs+3DUmOd
xevsPCtROflZ/r+yH8MuGFVzRSSXIN4PmBRh2wLhxJYaZnrkjik5VzSdf441wOQuoT990Njyc5ge
VWd+mQzeAvVQ881jh+qfWXh6cPv9x40iwEOjBZv1nDgsVHApbjlSCzOxz05rHoVTYxvkLhfFh5hD
AlSiZUmPq1yimooQHChP6OgHHykvRwNtwwi4v1H8kdQIzfxo+S21B5A5ha7BtBJ9VOnUvQqNh92Y
S/dk5nYxI7x7r6GSgGph99B4NrDcRxzatqUp4ftA6np/2p3rgyU6eWoXW8cK8/WcKoaNxtgqFaeX
7CxrBagmycxBt3rR13QqbyykOYogUbiosngbNfIDy7Mk7tMfqXoz5BAPAe8yTUt496dbT8U/ZZvU
ArC6Oy7Wi5E0UDqDB8ymXyZssn9uqB7e1jwnikA7NxOYutjA2/S5LuAJiMzS4yCMVhhRYJ3FTbdd
jTJgLVaYhOhe8A2qOtD08WRbLbmH6NzFB295hr4nJQTd9HYuvjqiTpLhVKSNLLo9qOxpVDUcok9r
TGsC0aZm2RmOi/W+aTsMtbnXLzvwUTBQOBnlZmSDRVB/wdeLiiQsRN7/moptnB75jKOxzEu9nts3
adGZY6gaSek2hWZptl4xYkIIDf5sh4lDjaOdxUY3px5QIPqUpkiO8sjuL719b7ENlQsXlD4OgR9R
HgFsWL7mn5gw3f1kh8ipSPw645YRqSHp7iQuaOU20+j0KzSGVM0IIbKV8P4fjIKZV1YVXCRs/zR/
rTLEpFamyz2QXAnVLEF+nQKAkYoFq55zYWWE9iCnMhvE8mxO3qw1mr/HRQERTqqC2E9zOEghfv99
A3t7paddn9B9oRCkCi1h8J1v9ZFLIUc3QvFeyiBD2sTeJw2e2AxN+bjRnhK4M2XfcwRW/x/C+2dX
Vm1ngZgRwd0eSoS6azIt7iu5ofoxV3+CBdnRsBTPVFgkzhRuobpcUdI+wlbWKoKrGgJPXLTsiGcl
R/ZfL48GLLwi1t4YLtVAexl0gHMWNlFilYIMnL/CYvp/Pr7g1BBcZmGkt6f+t9gyM15LyxNlapEP
bIC32O87ADZt5YmRtF613zgOagjFHNVIot2Y8WKtDZj+rWzmCIONBtJmYQyUd1e86bfkfjcP4g9y
I5ayA/zUa6Ky6666c26ASLPgeyPaEgse9GXhR2kFbRX6VlMay/EFsgZ4vUB+wx7GHgPfuDt/gRb7
MLYRojBYJYYKY32l++F+SpL3InwnX/ULT9FgnOlA6WxlqygIu7Y9vcidZsbujQ+msV/utfnHTRSe
eZkGvS0kHNaa4jrMQKoA4dZt/NQD7bEk79CEM3smTH1miGpeTD1gapsPmor390HadClUa0I0DxLd
NJ2b/1BSFDHSA+PvWYZgCjMKW8IFNv+vxDRTQ+qqLD5L2X0TQX9beTH3+QlnUXJlkxHXY1MJkDoJ
qysuEhVozgU72bSeJzK9xlrfTSVXJEaH+oncCqucfsS+/qv7tD1oBFYuXlhU1QzDC4rP9B+WF55f
N/uRBKdcl2xRuS/tA8UZgvif7Z6kRxEfxhlJ5Zpp82J0dY4T97FSAZIJ4CUh1w27cO4UrjNEbXPa
gUq76DMzPkd4FaleZ8oimzKxtXWr4vuJWEE/gp8Icdeh8Pte+JWM6bDViyXI4ZejpVD+JaYrZFcS
qYktivtCxpBFi8BXLiSTggdL/Qet5fvdiEOb9+i0dHa0RZGncXye+OuTmytrs710wZLqbs6pdC2x
gJiQtVEVJY247SQVT2zZnjMm1DVSqwQObWA2BduzX1lOVvvFvMOald1mZKb5lYb0E4ufIW1012Lh
sntp0XTOHSrFlPpsWMO6vnuCw1cQHhPZrc6KHLeuCHlnAWGOLPG50cz9b9fos7ZX2qb4dPXrFO1o
iWEK3WhBc8YKQIU62g6P2/hSOXeMipcSXKbn5UZfWs79QIa4xqxIfo3PJCODj7D0G6IEA9Wj4ncy
fLLkitkbaKuofZCp3jBnhkWh0zgSutfn/QDVLyMO/GPfvsypQdyBoj8hQsrnycyaZtELCRcsDGVs
8Y6MUzYjxDaTDfJ/fi4UKPHMToVU92Qz3Qrxe5F8S5YBJlCrciAfb1HQLZCQAOA8N8XpxH6bLesR
+xGj7OqPEgfY86iLbL1xKSss+aADzR1rMFHKdzvgMlRpt1y0PlPHWXX262yYjHd6JkuLSG5bfxTf
IAx4NbhRJChu5P1ghfM8C9ywPX/4fNlvCGmGMKF4EAC2osEPsAW+jVy/iDSY38LrrDyEge+l/xQ3
dQlGreRiMf24/Gb65C0oHD1LweYGujWDloFsJMoA2Lwjy1Y5Vq0ptsyUFoF//2nXJYZKW1IN5Xa2
a62xDRKCXyksFVmq3rlMiiT2uu0dEm7mSR7A6osFDkr622QDPy4GVWZloktxshjHy/0AtHkgpXqK
fU3sgSO7HYbe+WK0UOtYw3llJZFNaDX2AsJMSUd+I8ru5UTBoAvZARv3CPE09jwUhc0VCrj4VsqS
yPE0mLj4nIp4HzhL9OIunc4e9UcoZw1HM5ITcg/0oWt0mgAjAsRCnOAldnWH+aOvyHZkkUPM9SOu
sgGRR5YQk3svxYSZDSvukw5Qb6zavHABD3mZOkucdTMgdyuIPyL2YJ2tSFpH+ImotgqGPZVLoSVC
ysRRE17FXRbdrNothEEdscZXda4w2Cb9ypV6xu8byNluyRl6zzrOhBkmjYBHjtKjq7yiqmnzIoTZ
XDkycPR0jOM+f3PO+Lec7XRnAWrmEhp8lhBG6qbzVPp5rNV5sIxC8rHZLccT53TOOAaIzUnWhRfZ
twYHwvAlT7w3WNR8CoGed7YVYBxx0BXCZt8NEcP9xL15tuxehDVukpQAKrRXNqeCS5YwD7hBlr41
QD/fDfhW9Stwg4LU0Me4ZNNURrdhuNXSLitzTDZNwOuP8+3KbEuYqd0e6OARhMuxEtZBPe9HjbUl
yzVd6fVf43Zpd5/a0N4ptlgS/oqfFM+oNGZPgaOOvw5BYi0VJ4W6t2ZfE2X2NpJX073RVSTEWEuM
N3UM5Nd6Wqs3Tz1T8vm1lUs25W/orOHq4TBcX6eVMVsBy5Odtpf4zswJgreJ58VMlamsxe29woEa
FxtX8+CG8BaFt/taDOW/nGw9gm2LNXl7GextxJD15oXjv28+Zl4aIU14t2nC0zRxtPyVqNujqn7S
YfnfEu0UQ+BKCjBz+nPT9QTDFmZpVnQ8kINE6aMO9WAUh5FS56+zyhqlvZKMDQ8oH7WtA2KfQVMB
HvugM17BIvSApyRdkKMQQ0N0T1ddEuZSkZ8nFVVXDSfolV8jESrEs/oti5FYKF3XB84NTBQl1mvv
qEpqeIciMRT5meZnmVoYQ2/S6U+3WJ/LwIgQiuE69bMXjtw06VT3MZrME6Wxs7SQbA/KjKB3Ybb+
3tEgn4PrErN+77r8WiQwgSz/cbTa6IbaZaAD0jEoU0BWvGe7o7B3CAeV3dXZ+egmqZvpJrx2Qsd/
8Qh4jOl5dahFc5G4YEjdEuUje/H7Zcn5MA1K0RC9KAb4o+P9JOof/HlYKm30iuxKra73dWu1zg73
IOszff7+ZFIYmWOO2a/WDBVyy/S7CYE2Fptj459picHCZ+/xs7Vyo6n8p5jLVa4NHKeS4/REDRMG
DMndJlEcvILAghVC1jdg683h7b0r/qCZ5QrfuPHy3uPZeAu91yQH0dwcJ82/gCZaj1A81fieJZjS
F9CW1ZOHQNlgtPG4rH/cTjPbHlwfFJBAewQKzRf8Z2GdisZR6Z/RlUa+R2Vs0DvZ2/fRFbe3WFgb
a/1prFAwk/sIbze5bVddEVX0usjkhtfvBX1az7TP5uF+I9Zqu1hb1q70NAh6J8g0BNB9tolSGUXS
o+LxHr+2aBUSBSIgL6oCYvvjgromZ41qjHyjuFTGemNGTkFcysxtQUuGmIAPFLvjuBePIfTwPfzG
yNQpLoB38IDtpUTzdtuc9+Nc2cWuKOCvJW+9Ed71HcKci3aeehf4bmhqUidfa1F7Ys6GLhTtUQlA
njcf0Zy9qrPP3cv48x+3+umHZ4ujYG4Ol1zch9nwMFU0QwA3wFGojaBoGLuwbflPs/+Aphohyu+m
TNbyegEhDsT6fKVi5Wfo5X4Xdfh0mkmV5r4QT71no1GRFMB/sJQBM2DwGlTfEXp0ECTAlG0TKSYj
9koO1ZP7cLRP+07Vabul2x4JgV4bT1dr5UZzt/8Fxzbql4eRO8A31nDMJBDhcYBwxB3HiqRDsom4
nXAnEaZzn5i6K/ELNbR2qPsY1PQJ8eifubxprbG9UPqtlsvHYjmmCh+u9mpp2ywxeGVbmxBFYZL6
ckh+WFwxbytgZaTrOvrXrVdXvGMV8pZCeAuITmhkiLP65zZWudM9ZA1TVEIokwq72UjsQc4rAGmI
zi1Su6THUBI0Hgr89umNIO6UjG2FujGgRctsQr8J+JIJa1w1fyWB+RL9aAOhbGibR+k+ix5TE9Su
S6gMKj7tQNgI/rxEZ2C+U4kw4ibbxUkfKz7EzQhqAO7jONP5TP7UnmpDS9fUqc6lmaHjte+8LTJM
udMxURG+6i9u8N4zXYPsw5Zdp6yVkTWVPcXFZAP8p3UcxcwJcTyXfEogE6iWaLq5cb9voVsifFQs
Q+lErK2gsSsu+nieUGV0BPVwajM4fyZLzMBNdTmL9PLiYUTDLmlpZ9xZMDy8wODu8XtnpEhp7L/K
VhSYzWHjUUdYt2mz7xCEyllrnKhVANQaNm74STEpEYDQgylOiwg5YiLSwyqRWSMCkMNo7EtTfK9l
p69nlIYmU+yiNtxsNxAW++xb3RrIi+nduqHJ2tKBLqKxWJltPz5XP2aYLZf/34xkzNv4WQV7i+qP
kXc+JljnoSpjLqdwwGsxlnEW2GfJROQ7az92DwpJny5i7GxpUllMDorRmR6dT1J1bARIflXrRUm3
9a3gexlc5Lj4hqoqMQz11ZQ6KOpmztjzFx+cnMapLF0Fi/i6Fx8lfkY51oXOBcHnhsJwv0NjBlo1
dLDOCzuJhyqCrq/X4D2gu8YU1Y06MdVlXuYnSBgVkdTm0Sbcb98m4WbbAmiVUTOZNpn2vpqeLQOC
ugjz8+EKeWao8codJu3Sp5SkuQalcvEvNbud81kr/xQPLWWDMvTnIgpsWfev40soXKZiZyH/Zqes
4eL12ijbk+7iwyHlypI45rGRoNbKQKzc3+iRKAE6r1W9miYaP35tksO9DwaMOUBVB3rAXsB01Ww1
oWfnInwrOu/xmlQimfh4G8+xDJomu9+0VX2Bmm25BAssyz0QMGdwmJ5noXqOpM9uXFF/uMVc6tzb
lNo2Au/0izREsIGwiDIvwtnpDoXOMqgsL+wFyxg8AdG4FOdvkjCeCRKM/E4ssGohSRigheOnJYp8
XzWEDU6hdGlhMw/DxgdKUHGhOHe7N2vOB3XblmdGTUOLaKP0zDjEOcPxGyuGbR1zRl2O6EyfGmzE
xsSOtytfStXfUSvblTj2QAaCyeykBd72QQDj9JAXMeXHWIPPYqBp1zgkgg5racEpI78DUPsEXyqy
mNmTHK774pfUimPTy9iZ0ukBION1Jph9f6yy9bU1mJ2Rdwgwfya4ik1kmkkSz6S8CtTRHySn8Wek
LrIz5Ny54kPDSFz8K9YU+4w/yKWGuLaZ1hqc9Fnt02FhacMxLsTlrk3+0G9DR1YFVf/RDFlVfV5G
E8woA8GVyHezUh1Iqrwk6Ev4CitwRdEleH6hJs0IWsk2EqWH3Gq+sKANJ3Gf/v8Asn59HoquJ6sy
PzD214oskTFgt4hXLHN7a//4pwLsSnRUEdYMG0L26Wb1yn9QIBM7QcuS+rGS6sGCy5qGpzuCWJOf
HKiy/zZbE2ElPEsh0feLR24hmRbhAIidp1uz5fpWC575lqwUXze+LA5E+WVItiFHOfoNUysspwcl
FKBzeFnmMvMZw9N3yqIZVYDWhLn+mjyUenyI0lXZzmi6C7jei1cVgta1lz2we3vb+KjyJ7PDGl5Z
JnkUPzUAdcCqazxtUltUw7Vd9R2iMZeJB9VPHE917QWcAMgwUlNLILo/j5JkQOkVW1xovjqCeO/L
4o2pMDKnjaj5C1pmezHRiXDafhXUoVPDd9628uX0+9Zyc9tlvpX2xU3gtzPe0E5uLG7K5gzez6SU
HMad1MIEisfizbuaMpinzHhvGMcPNChp6uim5gqPixF46OrORYFeBWS5HQRDHVma4I9EI49wEqZ7
rqvx2jZuo5rBJELN/8IPfryQlpf5XQr3Md/zTzS+YlWX7B+2SrAw9/8ANxxjkwEkkrlpIX9LsrcG
7ZIL6YjvtQQNycSSQEOwsHqGUvaWwCgscihVpwuWAFcyOoTZFYhMyqKyNIhlygPhY56CeUjqGuEg
+HZYOL0AxLc5Fvcl2zdimwvcWzzDEtcemd3st+zH3w5kaBzEWxq16tdu8Bo0rL3IWd+gGzsTs2pS
d1aVeXi7GX0YmYcDHAO8shq+o1orIXqF1CljBrNNsJ5t0db9C7o9VhQq+GkdyAgX09jxUBGY+14J
RNidjipdSfydewTgYuKSt05/zYfL719aWCvW5/RCPgZ+W4OTJUMWMO9ePGYzT/QEJ2kylPT4zGpg
NEdXVDJDyJtEdcmtfKdwSnuFPQzgrrnFT3/I25jF5Xca8gyj2sOgjNRKC11XSNYAXs13SWmZLxJT
Rm5MvYOAkdpexEPxayEqD6C1LVAIqL6xfMq0059zQO6cyUN6Am7AL9IHHjwSMmD/8Xg3jErKnpLw
4R/O8fkxd2qPt03J3Z6dzg1Hd6hy7dL/DrhWN87C7b6nfeiIa75OlkaHJyOI34oX89ApF829FTJ7
1sQzIr+VDBCzUIVgsICOWrIuhQck42k2kcvZO+K22CNwdswOm2aKTxPYpCibLkR18qD6yK9VdaK7
u7OxY0fxsLSeC2omN+yTCZ5lAH7kUN7plC79PoNBJdMri1i7rryToId7iJUasjSz+AJErou9clRb
eLDar8puLroqBPkZDLdgqWsI0DuaXUgRSGL9sjUHOUxKuY3aAVBFf5ksI6i93dvZA9MaSw7rSn6Z
NAhG+8C3giijktNkgMlUDgB5yVljiagAOom5iKaTQU+trHaSLl8CH6rF++DYyAiVzRj7zf1ol1yr
/jh3YNjttZXi/M8wVhrN49G/S/tiW6D4r4DQjFO/GiqsfU7TTCGwAWlmv6sy4CuqyCjGCkRFLaDc
ctMpp2zxoupbFTyb0c/Co2z1yCPUwJrQkiL3ne+HcD/2AZXN0rl4kGGp5X4WVPYh56o+xQm9Td8I
+TskBkYE/MLWdUmmcGfuEWaz1G9nanbjOobZENTKF3IifY4o1VLzNYyjYYL6BsOuJxE4d6e2wjju
fnVct89I+umYTSNIGWt1q3SC5kEOLYw7K3KvgkW2YZ9KJaBOvN/ys2/PMAFUjg06il3Ewy8hU9y5
KvsvaConeJ+MkOwE/EnrExOWc68T3LVwfZdpJKlDRD6u891j1dZfrk/TnYlmmgD4s/gjyLM6VZBh
4qR4AY3KLhwqw53jV4mis4ZJdKWotSHnn4jpQ+12YuU1ruHXMNB7eZ/D7+Su+jXUdpJXkLTbtOlO
GrRB083vtpIm7lfXmIP8tMoiRusGtYrXIS7g60tS4icPGPWBIamcDq2m7nHtdpElV8VuaVcGBAb8
+AJAtYZPwz0fRzmOit/kAuDLb0Vi8k1/qpTwVAiERDC6V4llGqq+n0ts26tnQ8XzC2SA5r+3XW2p
yhxX977eYOOOHerPrFVuowAkb0mvLB3oARk8vPOz+AJBz0kfX3VOeb3VFduOLN76/4jNYGVbxxdS
qrLJzCwjWxPzEaFNl/YgSsc+mVk/NfVIKsBHS4Toctn0IFT3fBmZ4CcmFRyOcM1ZZXi1fr30d89T
oyfhe7rW1uIZzCyuzS4i3fazpr/vPK5nUHqfxBXjWoQbT5dXKVQqDlBLLm5L//u1oM771XdHwxir
xa+6yYMhvmw67apuEj9psgwyA69BZQVrxe99rKPZTqKcUZCZ/va1//VF7eJsq/LbWs7Cp3LTJymD
MdJ8BrLX/Jt5jYc722CxwN1/I8qjewXe8M13DBLarxY2uJRXhV45bXPhk6PbP9Xrwf+dEkyOT7Ev
HlvxI+L/qMTDqUlRlrDNelHz9e9p4lrwum4YAnxlW3XzdQXTTmqjDnOITW6vEPRs9wXTPOczTlP8
29Yz0DlRC3kKHZxxuXl5a5ewFKSCuCaGUy+wlFp8qGkAXpAjBg9rQWEzS/UTd+eBcSGRBOWJ3Ecb
Mb6BLlqOX4d55Ewujg2uNYi8a/gKFb733F782HVYLGz12rbMZhfk3uDjqwHyygOlomsV1U5CRT1p
M1ej1mSsU3YnzVSiiC/gTBzldYUITdoHSSSlTFEnXuvE6cQpP/FBvxFkpa5AbZ1I6JJwa3e9sa0r
NXx92OtpNwk9IFayR7RqtVkcVbA8ArTAmQkn/AV0YG69+Lu3AOT/Lxj7hFMUDpjZuLMdCRhPIenM
akaV2OYTJ/M5MLapZ0K7m5HcAkX/rmGtk1YtoN3GPIz7FB7Y+FGIpR3J0+xQTqQZowa+F4nnkNnG
Eu7MVkUZhnPe7Lf6wFeIkuNGg3N/m8Zq2Jj746ARJ+VT59GYC/7jKxlXnWLOUezKj9gpQgrjOBXW
KgfGYyTNqNFA+6GPGDDGow6YqYsU6SrUBLbxI6clOu09ymVV8LiJtZCNBxajvFfpPw1HuHieUFK5
/12n4ngbbNMbUuxnM7Yj2Yeb2Yok6XnXbfMP8uAWeVLAVkF+TAN6lIIoNktsO+ZuFqXCPdduIF/U
aTrst3RgyitGg8CDhDxRb9BkdgmPM204EAaDihshmsqLU3agBSgoZdlQszqQbVO717rTdNtOktrM
uSTI/uwT8dET1Yh19wqnMWuBd5B01ZA0TZ2MvRSbDOqsyMlJrq2oByrz1SkiaKABQ9qgyLnJALWO
qYx5lqyp2ydG06ZuVJBZhGejPSL2m/sNqEaCeCbZ2UTAyQA7BUqki0rO3bhlo0tw9QqaAT5LYH2f
nfnNtbFAlSRU9UL9heaGON5PWpVA3/4s9Vps4Gn1aci0A9orF2lYZCQmd1sy/ObDPtqz5QXR+KrM
Q4bquvFpszv1SYX2SdunKuD470C+0l8L27aHADz11ymwOPkSlMSwT6TA74spItUYd3rs/JwoBzOL
upzB/UPM0VSnM8k5C7e0AkH8a3L1qJy4WfuGrnhOijWwfAY6rEu8KuiiDoPMtIMvf5+LOUKgTGEI
ldn/1qJk+jhbpMAx4TEzb65fovBhe9ppr1lY8D0eLxWdN+9CTBrxQbxUrHXO5LygbKK7vvUX5fnj
HQIybYHVZnkuZbN2xdFo04hHFokS3xDDUWAW1Q9UsbbOW1XkOJCM5wGC/RlSQi25id5cENtdkIiK
uLiYI0asejJZFfaZ+ZFF0tzJh+Yme23ND5gt20EawixBvYkZ2d8ApcbqFeUuK8mVfR0bINNDc35p
z0ggFrE7E5VrxNOmYBO8iBEyAUuRqVTqLi+8NmQ2EZQiLF+bdjjfqiSeCMV3kuK5nz1g4iNzLna5
omUi8QX4EBj3AxN0cDDX0ixLE2AM4uK5c+4nc776/PhnUlj34RJ1UdWHs3BEHJGOD1bQxh9nKaPB
QDUMeEDhD8V7CXFTSncs4jFTiSuD1nd9WfwMUTNVwJ4cRnmzOiIEd8s8WkhABDdMzNaNHa8EJi5F
PYjEmsKB1Vo29IpTB9D6DS+ff6TeRCEMBY5BUOC0nHjJgJG/c4fxH95k0t3/M56I23F5pKK2bfAH
40MA1DcmZ9sidTCGbNwUDftFSk/NsLqPKkIELUHbmgFy98id5HqhkHWOnpzONiEM+E+J0OAYZj+h
3MDGgTCEShaw+Wg9LTxLkWAkTY9VxgC2g2abRaQ3IPawVHyvF8dkhLgp2ZdERegPo9NsflFIRzyO
JrWXBL8hSka/S8Ql6Gy+DB4nWxHbfCszKmUtzu6sA8detK69q3tDGj9eJakB593IG3+c3Uihqju8
fbZmgrfFbDlTUVJThG4gnSdRpwWdp+f7xluU5y3OE9bIPShv77veet5fGWOPgOJY9+c+RVqsBeLz
T9GrpcJZHbocqefysWT1BDt7TylSmf4E3Cwoff+WAkkwaHcwxK8OfXKQy0VTHJIQIyncRJx1/Pqo
ZwKYkyGLidh6iuStl7GD5MHwX95eulel/dPtMYMbR90ceLv+yELSud3EJIYZYy147qem9Nyaivrx
14MTZGuOkSYXEeNfO4bNPGNrbbi+KBwFPMjqkan8Pmez1QfbhIK+OiUZYeDGlteZTRj7j3Cn/y7W
MfjbUOXClwwWDG1MvSDD7ee5vmxfUVdRYw+Vip0ngpEIxEEhyu6U9HJ/NSkJ++6tAikv0IqxHIrx
/tnCgJUl6sahGb+ckzq/1UQTZKacI9HG9a3mPkwTmQIJNlBk1UQMtbKY13L0b8wueTeaKqJxNG0Z
LST1pYvaI9flWYbevhleDugyCB93vRr2X5JmU6tV1msDN/6lLP7Y4H2QgvtcolXnQBZeASRYrK6A
yRSV6mJqm99Z1i/3xh5pIVz+EtEsSQjYiHAl0NKk8VcKKGSPSI8b7wmLitbpYY6r1582caK+MgHP
kMJ01SwJsfiFPO/KFdA1towyqTgsRo3qjNX7pwMcLuogiyCOaxJiWzsS42oj4Vb11o4L19wi2i+0
vxhUVXaLIAb4+Qp27dPHBiXE0hbTN3fi6TcJLlBflwnXAZICD8GU9GVBsRD4Ju8+fRvMMwhJOEXz
+rFAHdlFp4eE0tWvlEX1zCrnbk4+q5ByEl7DiWHI0S2TQGWx08TSnXMHJlYISzCPlDMn2mMDavYs
Am0NBRK4okBxpQ12SLgjJLeQEXf8pnROUsDBuo+tZUXZveSh4P1vf3EJ6Y9wXwdZyMuNPnG8oNYd
FVrvvojrGOTB/S5+WZFVFoFppARdbFlvbN7jYwc3G1NwvqMGEXFB6YOPTPg80XbPVYvw1auXp3EI
0VAW3dSSPG4XGq1RcZ5K/v1gQowq19PGaUXDbjz8PlrzQQfkX3r2R1PSLjmYwPLup3nk1+IHHH3j
/8oX2YFaQc6CAehNFoYrkdAPHG1iTDykXRBPIzzYnM0iwx+ztyRJEHFBaYMiokeDd08pGeL6w0zt
hSWW46z60va3rtDDyltnwpBmVOUwEvXuOgwm8/S+iy8srcO197Pe4hEjrsl+akYwhqD3O/b33csY
2dkfESoUBq0YRctMoViKryAu1UV71mlg5Zh3uWS62ek6sRajSiGnrydFN0rm1xukZlfkpX/MYQTR
KGCjbmwKWQCfmpVqoJXxGKMAgbovUi+Hc7EkABbSu9RofLFVSF8Dm8Rq390dqYZXumxvCv9HHF0q
S2+SYEro2HT9JqCjwtovnMHegjuRz5KNtAuZjambgJ54Vn/xnattTXkk3TgvC7OY55/VUQYE/sjK
P+H1xYyofKP7htPTkxEkIh5Mcg9Dn1yswAVMdmOJwe8oB2Sy/qFuUkuwsDNv25yE8KRegMJ4SA2r
4xDcFnk/Nt9ttsg6MYmfBy0tft/G+3Zd7r5f0LZuM+S+AhUGylBYgAGE9nv7LFlCOFjfOMe8Esde
dV5vrL5ClB36818IQ2/o0yG9hEOo3Hchyu7iaQTo9jdQOKs4kfciLywqHxlfeJtxIKB3iu9LAFX5
IIG+LwFdnVwTnrkH+w/8i5EwTSgOEW7y5uFH4VSMNbZPQcULjkT9YxOvWKV3WVJV87kXYN3pOqdI
atxny4XJByJVPW2TxQGEE75IgxutC47+Au9syP80o/TFFqGh2Dlmhp6LtFRm7n2ZVUQuVXWgMjrc
inGul6Hbmaor7yqUA4T3ug/fmLilER4D3SfNUn1ZvAWsQoCBtmWdsYZOH/CzG7XGONxsKK2hYyIn
ASg2z8KEfPgzo5RSN/ApnqLjl3BdKTID4Xjs338AVlKK656xuZ2dGZOGCrinb6DR2Vz7cgjmOaR6
ouANN8vVMUOf8Fe2mY5MXY5UihBYktsP8a3s9nHB7B+sq42rUPHED2n9MPihgGhwkvwk28U4tayA
sz6Jb7wtSzXjTNpmEZ+HGGdizmy/YAZ0CNoTZ5LWsCn3PC7G5q03vabyfxZaojsI4DcDsoArwSeo
jHDkHbfB7tT49FIiP/IXRYU05x43KpcYq3yjxLBi1HY0/ysbnYsPAFn/K1ip/+AlbFMX00BfWiYz
vwvSAIoghvHt3TPESa53MKF/GS5QYoP9nO2KWKIrR+IhIvG6MWJLvPGL/C+ANib/m6SOQ0dr17g/
q6MGgf6Bjcg/jQwcSO2D4Kl6yk+JBgg4cgRDavBnoCCfiQjWdYOZOgIk/QqcJLxjAW+nR74+uFrP
bs8/0fqeWr8VRkynfxb+4jSqHdTM3fl7D0PijsTTva3nAS3fTiftdgbJZ8p9yIgHlWOKSsWEzFpJ
MDGnr4Xcox77/AJSmdG6b2xBX+x6s7SYAQR/U2vsTVv8Alcvjmtoey6S/aeyeIQbEpxiJPO0ormG
IP9z22GxMrytv8zOAlysneR+Eg1xgZHjrIZYWnGmdOtPefabsOUA2LY7sV4Ek6azhhvAM4TUko1H
v9IQEEO5MdDWmLwIPPCw10d15DIPS/0yuw75H69ASHzUXGsd+3k2yv2EZ+cPNYYQdMjbME0WR/PF
5npx/xBcknqdqH0UjZV7cJ53A/zwYpuTMdJYFtrA2kZmM80wU0MIE3nidVjaxmh8mOnslH+SiXs0
r8hdrZ2b0j7mAvTIptO6bkZO+YTgtJXcSPvvuLB7zOliAU9O6xO0Dm2oOJ2iNjp/GBC5v0ilGeqR
MAb7/mDzVS9dZ0iUMCsrdJFa8dk+JXE7r/wrxlU2lukF5shyA46EBXfrrPapcRB1Awgu7lEnUymZ
kMnpVWvJ5Q354LBBUUcAZofi+nbiLYCJSpAinNA5tHh23kdjJfnqnGUGIZKvzbIwmnqxTHwp9Y1m
+qiAMPT5xmZ2c1zcFFFq7pzELsM7W3zzJHg+RNUtrIiKrzxbL/z195qTsKvQl4SShcYhvipeddaC
P9eV0Do0ty6/c7BnSmBTDVtBNCygnVDuOwHL+5AJhljPqR6YmF4pfFjbw44m8oa8U10WTYRz7cud
0vBCdLqSIwigZ8BHXpzXJ4O7McvooXsKZfTkDcgJ7aIiDY6cYtyJjjdBwie1mAtaI34TKK8/bfTk
dxTQOQdnkPdxsD8X64RVbkUrwvzd8nt3IMjnZMjGlJeVPcjvEpu/z0C0S0Mxe088ountUfzbWMpx
0lEjPuYMDHPd8CobUwi/bY27hpiOnA7XlA9zbrIGQfF3milabls+hRe0jcQe3BYhRaCH+aMD7RzQ
153sd0FqiXnDlIhk4FpfqSDHPrdyG/A7Ba/9RFL0evCoY8mG87/5KFfL8u0GUUAfGny7vKcGzgBf
Gem+UJ9MSTKy8Hu9HBK/exoxI8Ynnrrmlbma8Ogj/Ty7x+cy21TPmgzyLkERqTjUVIDxuD+BPK6q
CX0qbGWiZer0ldY1gTYyBp7V2cEVqOVpbYQTCYIMq3Y4FGN2+YoS9mfwBh4Gdk0Ph+8WgvOz8rSh
6c+r5hlMHZNDds1Ux37sz7v0sU6yxDuCJgT4/n2dZckcNrJMNrpAXMJx33/D/v3sVW+bnmUbQlse
esu/ZSJsoo6GmutiOHI1DOqcOmikCoWjgbkqniGdF6JWxjaQ/QxTT5bbUtYK98rmnlO0JUQWOrN/
8Sj6rnzc5i4jF41b/zTUuJKzDB5CivW0SoRVa25DRIPxHSnOArSvBoX8xiZrLqx55+kTLeq5ALJW
s3Wr1DAmEqTE5Q+gCkfrisIoUwSNDVCTtMpO3WEpFcHrTTyNoMehA0rgQL5HtpItVK3TA+8R1CbI
mCQCKcr4GwAYpGLMy5qyT483mUs4CtX0Aa8yy1Oo++f+crYC2T4riArabSPq5qkHQ3MoN5zeUlNP
Un8QPs1KBsCBLdNPw2i9sUua1gKKyxezz4ZKLjLVv/LaDIG5G61+9NSNUDneAdZ2dL05wXwywz0G
/mVW3pUo/h7VN2k2yUNxayhxPvZcwXtE5tZOsHMpRXHL91yahxKwSzqlgWZ+zkE/Q92oqVW/U+Jl
5yN7E0x2d2Lrd3h5/73SmMJwh9GR9tC/cegr7c6iIi6auCzV604WkBNkEW01zr28ZsrX514skmVr
uk1N8AxhfqfiJrVryaPw1kQLfgyDeBCIkKqG424Vk6NxWp1MYqfYSlGhiSjsoGFlSqI5Nr4Yl2fV
uGrhl/FRnZuLPHKkbEbIq29J7HH84CSJyove6WSuYxZKi5fTJ0izs4kyuCVdb+UCmPxnw+tt7MzO
Nf6XZOAYOmjCRN5jqj2mLiPvrLhYzWnnFqG86BMEuiMoEkdc7Cw6PWqtL+iqeqJEo9z8glx0s35G
D62v2fZ6KIhDG+ImVkdjETHTIIcCdr8t5rdQv8RZ30TM7sMJNSuRA5ekdo4DCfiqri1+TgpiJuSX
HwewuXAWz19+utUFwAI5Zmn+8Bjucg1o/dGDFXkh5FlBvL3pPW2kbnRTG+h4z7uoJJ2HxW7z7ySW
6VJEkffD9FeELxZNZ+Buk5prqHyihKbLRA/uxsA2AxFGJAN1MIIXWCHru2zKVm8nmSED3gL+T11V
1E5bgXpsDWF2yVAH12wd6+AQQsCVilgVRf0F77qMnT9/IU976AulHk5m6uUiWQbBcf1qLiVycV8g
wJ9RD7DYDE7CrxDAWYrU1TBFR0VbRnkazbEejsh3Em9unoJ47ILgxb3zqCaIwMKOS3XJir66jCwR
y4z+VYpIc1moZokumtWzbPluZC6EuUn3Gk1/cE0fR0tzAaJoY0j7WxLmvn4YDCtTRRUa25CMKvx1
87q4y/RkrqKTpS5NV0/xqnUpIuAzxtr9n1fnHwqt8Aqr2xqzWAD52A8Iqe+I13skLKP8dECDgCtB
Nqa6xAeAtYHeSzBRwRjPRg7sFkZXMhrmWiSvXsx2Akcwu43yTZNv65Z14G2rYWGTBlM3RlR9H1XI
R0ZB0IG0j27CpU35pwtwkJ+0yPe6hngRYE4/QVSkZGsLKp0bO/NuJug6RFFjEkghqgvdY4hGT3t9
TXhkR18U906SCMSsqraAUXy4cwopkN4hSdYDmk0yjvSS5kcCgKM1HwBvP3IGTs6zLmilRnwuxXWz
qAgWbpz+IJNbY40m00EgkatPytzC+C6xBysBZ8m0HY5ykO0cQuPzD7Cdw/ZIdshkKDX3YQ/9YlVk
f/s+B2CbozrxzY3/MfEOAfP10FlTdNBGMaV47h0JLuRxuopbtd7nrURhAORB4US66HA2iM9wPHEV
Us+rY8yuFlfqpqWuWI6263MooMpde/vJTuRvM+u+gdIZ3/MqEGiSIVExspHYya+HP8NVbGn/GBqD
j+Jbz9qDmEDtyqxz2DF9IeMR57RNvyTLBxFZkUPVDUx9cSMOaZ+1Hs73jY6CRj0pvYXsUevIMrvB
r9YZ0mZ81ynRgXcDMBQHMSmtn5iipvlNZ/Y3k1Cfjwh/0ObdaD9UM6gMRlNAuY6ivF8tBPZZKDAW
KlEDxEmpNaLzNjcgzvhtS+/wU49B5TM/pT0kYyG77GUrXr5c/Dz8Kc6xmVRFatu9X5D86ssujIop
IEt/5FHIj3WKXkaIHibrlUio9sF7L0BdgJ9TIKeuvsRZKjw969tETtpm8AzbrY4fRTJ4osXOAX7y
IXNQqa7/3ZWW3mqUdUjVKLzAtPMvVFtz8boHfICp2BaR5Kf2zN/nDI47m3rIOqctlJKcE7iewrNX
CAjGgaO07aB7yxk/1qMZHak5Hs2GU99bhxgNFX8u8Ne0CWgu697QGV72vG/msN4DqUrWmQxiu2xS
oI2rP84xUzXg99TpJgf0Z5JMx7XYAMgqz/gzvee6PQv7C2JeT/HyD4AnY7wTGbtsiMIn74EF9PQs
e+iz48UZBVGaTI8jDcLgrS98XIssN3B5rk/XBEaj/L1mWLLEYfsSnTtYcbMpOGSQx+yDUx2tunx5
C3TuxXkuyXnKjU8dWB8DVP6aoloWsfkr6vUC/kEl+MPBZY5h9KCSkKfvBYTiZFVlF0zdFMRycgNu
rwHC9m5A+Ax0230dKMAIFSr+EZwZUPVXwMaKIjUTBFmYwETkUepQDWDoLvFMjHRu4jfCevchf4QI
L+hDcuWK0L5WqNL5HacXJMx0tJSwDmSgFh93/ocLc3QzngtJv8qyJ8B7yZkTxO1DwA3dhU8fGWTB
Ozg3O2kEOPWHBcM8I2Z5APtxeXnFNw64Jy3SmJrfitUNHXkN+pMXEl1pJ2MuQ0HUh2QVNws9qjeG
gOvSFp+ysIia2vILTtQ4S+pAY1oxD8jSeb5AiRrcHRYwx2Z7r1uoKUp0NyTkvsH8WdpLeNl7nWt5
c4uL7qal7yDlGWMlyK2Nm2enByLiE58W3nvozfUvEj2z1/VGet6IW1rhY67jy3vOafOYZZA9EgKj
Ritw/VQjBLXEPv3Q0IUwSDQ6/m+ckYAMn3gxyRussUKlRdQiLzQxxPTwghjnuVCu0K/Ulc9m0xlN
+FxZ+XB47SymUHcziABLJKPbKddhAu0VV9yk7oncGOiDLdpLXJjmN5P/exj/Dx1leVp9YUnEoSey
uRLs2abggPqJGtCs6/6YoXOIslCndMSCeGgfc3r/2+4mxH8x/lTa0tG7GrPFvGq8pK96lCo7AhGX
sy3SNtIL0wPQpk1iKZ1JnywzPIbbFd+CtsmMO+d4W68dEz7gUcpMc5yeEtjjofRytUc+xfUQK3m1
Ky5JI98Pz1MbZM4axULlVuYwwOi8V9RHA+GlHahEKNPPjrsZUntpO5K6ulcfMy+RRInZXNVk6QRl
wGIl1lOvXNiNqkKw3PQkm4QWmWqdAXWQxJvHeGfejIhjaSn2kjy5o/RhShp7nX2Vo9qdy6Jy9WtD
0o395/SyyW+gBdd8pApMF5lNystQ8oyHzBxkD7JT9quQd5Qwn6sElA4y6jKWSuFbxTSUC5nktn+7
MJc0/Yrp7Tg3xB+LB/HVIiJA833BdNXgZNjpDn9vO35x8RDWCYT0+GqdjSbTG+2/OJFzUjbIgk75
JtIY8DEkQSbdZounkBp1OWUCULbzoudAHVZOxEj15Hqw/qwA6Gsbn34l10pvjjjuc5K8hYi3eoTO
tblGYEOtBVW71btQzOjPLykAKpMM6XP56X7ilHA50xBqPmeEedRUQ4oa0MBHPCnthmCMBGiCorsC
WWvfA59ruJV5IWYVjdpi24smFasS3VGrFkl3/spvnH+3zIsxrAqa326RqDj5U3TBenptkbkaS2g0
y5me/3oZqyN7YhK6xjGAEdslbNszKthLUlTdcp8c8IbRdPcbGvcOeF/xlqYRO0MXH8bsrYUpTixf
zha7qNgCB8hKiVuY26ACv3FhfMRoLVEaJkq5NnTfGCrLtj3PpQleY7V7Daymu1coufEjYrQYtDbF
2ZDduIRgENWgMU1OqukDTlGtOsaefYI0/gcTkMqN6RpX34PMSfnMpS9Sg0DvVrdbPaDfleyXQqCW
7RHma+ViraanZNM4kGBXgBJu1SLxT/cZOKt2KhfZ7yM3xP+SZlOyg6+WaXeBm5+9QSYFRqjcBawK
AZoArUfgBPxpKL2BqgamwLOnO/YTE17D/FHehSncMJTApd+J0GrMOKZ/7Lu3PX5po7XBSQOmgHZx
0bCusHCw8ptO0E5D7hvF29HhHbVriXfDrMrnGi5kHr2w5n7bNwOovdWDzdIU+luQYbF7zVgIjdYB
BR8ccBJMPuA3SM/9xV60HvbfYsGx+JNoUZZvPzddeGKV5+mnGhEaf8bo5YWqjSytitLLX9AVCCg2
CiZeazNgI9QceCkH43/mPvdwK+udFTQZu9Umeq8S35CgQgKUxRXnDE01zJYqKQhP3Q807DD4i7dx
4OdChDZApYNg9eheqfifwwK+T9sJNmty9P4LuoFT9q6HEZl2nYblCDEopUDrg7uaHvHzqv8IxSrN
ED/fd/Cs7EKabkNN6qMrTfL0F71fVdrRAr+7k698GZKj6ZirmQaQ1Evr5NR5K3wjbGNKYoDlrZJ/
xDCNoKA+sDqXUIytLV0dQpCJsZ6tocaKU5Za0fSY7h836EvEyCdop2q/VyhZmEyNFwaT20hV8xON
nZxPafTOABykI30C64s4g3QjFewozsGDUGdn6CKQt4KbH9gLD7iaOjRQjDXsjmWgjN12rqcz4gor
CKqwX6nUZHAkt1dIk185tGySdEISNLMBHfIP+fg+SaoD5zPTNgeYhGF2UhYBGxzW/JWOsjM2wfSJ
fQ1l1a+AcmlewvuKWFP9jE/LVPd9HY39qo8R+wN67elRuW9onaCnH+R8DKp3hMpIhhXgvoexAVy2
Qsv60DWeaec4rhoFzhLkOyjpb0ZizNJQ5Qs5XaBEjRnJEmq8rSHbJAzStgkSamFNa28bcJkYxviY
S98W8Ei1RJgo0RnM9LsfVxrFwKMj7DwqFjD1ZIm4ib3bh9Q9Mfw5yesSGHZDE8Ry3TlmjNYg0Y+z
aTzz/8szq8HHoZJNI9Gj9HjGLmBuFuFRFyOp75cfbIYaHMvHy8k/I81EtyiuL5hGOEl8HtPefmFn
CMiChbaGLXTFfew56hayyJYbLFbjWn0mav5+wiDPLq2dcv2IbSpIjuXaR1NSretEeny7ef5Xj7ye
qoHl5nH5AdXwxdHQmg38359sx3W9VhpZKehl383b0qQQx2XigoHK/9H3oW6H5MNsyfoiv5KdJFwT
O5ral62QcBCXrtv8Cs04hkcFHeX6+doXmOuaTKsLlEA+zta2Ix9SDpQT79pZDmANEC7frTDeUME2
hBokPwEanlKijUnOnwq8fp/8DVbjFxfx0pL/mq1fzLVCNrSWWbaow9RJ9pkamI9aXeO+BIIuEPwW
leahkidI/aIDKwu5i+hn1CPLkJFCFsiqeIoERNJvTK8Qpo+2bMinr/qOxcfK8nuDKwmSRe9Vj+UC
QY97f556s+16vOHPHujqR1cDNWBuOemFPizCO/Mt292odNm9LQv4kpL8Dc/YDhmoknb0H/kaKKlO
5O7aur8CbvJYmUIw4YZjjYGoEpIOzCkl5AYZF3L+xrSc2P4iMBm4PAXdLiYXqo32RC+2vT53ak8a
KEVE3ewfO1cFKK2E5QBHcRrwwDUWEtaV1+RFzdZeS/SjNrN2PClgO/pc/zAtKKByLRWpmWdzEizl
8iMDMTJ3x+4yqTwhGv+tXdJQ83qKpgXjtq7jU95HwCBSJKiYs03kljYEWdVl3aX0ctVP88JqhB/k
4A+Mn0PXkQhxNr4bCM/sf2cyB7drn7T0x9gzTpXHIjBnVF0jQa7arjz7t3LsQdHGO07C0s7Kd8Zr
JZqTR3rPzjxpbrS5q6xdqxaaFbBUh8Ydcvfw+20WPONK/Lc61GAAQIYduwMyARKn2iufn2ELJcYT
EKOSR8OeF61vEgcGseMJ9NWxazBXZQtUUjpTZwrZPjpf5s2q8eDuOlD6Ty07e55Zq5MGwmy7CI5F
vCwBVYSfaVUHjzl/Sui0HLoeuUCNJvl73XsOomkoe3WirgfHdq7VS0MkllSTVGZrMipsLqpYM/To
V+dYo3oqjbjbZpX2hcLR00OgUtuxZVhXus6u7rhn3yr+CUQmvDWaeRlpUjzrqKgzrLmPeWTAlMIH
khU8lfRc4iAVDrg5JEL4L6fzxejThOhWg8W86szuvUvPIFaTiLLamOGs+AbzLqO+/t1rDSE9mntn
uyh5cTRmuTDl7treRAyUw/UuwEIr61C5KqKFFbZGG0XY3cGMsWNc0L5a0Y/8vhXaerAdALFSNFEE
vBDihwq+QyqIEuPaIHcipYzgCpNenmuXqs6SIC2Ld2kmQw+KUUn4k62h58JnkR22O910J8HUTScH
O6IzBuM+9TofB3b9TmXjl5Qv2gOtAmKXwRmf41CCvHjHds+3CtD3b48diLlE/ygpM43+ZCwaSBdB
ujFWZuKacvKBa+h5755nAPQRR5QssDjRmK/6XspE4NN4ChnpKCYWGlrmr6mFaZzwoOeeGe0d4wlE
rW97VrMeAFTFlfZ+6X9p82d/rwlAZVvobCWV1t03B161Rz0xEYAAhUcPRGdXVKcbiMGOqC54NvVz
tLfyKwJUi2bwSjOKEeoZBtzxh/THsmGLnD1nRkOqPcnHcndnNiRosUbTUaFnfROCMCFoIfBaqlXn
xNZT6p1y2zk0l9NwTxIH5d7Y0gyr1I3TSe259nZxJxEWaMhfJu+qq9U09/sWToj87QNnMw9QfqNM
7x5WFETe1dFzSIdxB+DI8FITpucciGhFu4uctlsOkzgxleGL05EE0VVGsb/JSYFMxZJIj7E/0EbI
T07p/gj3NchA4Ngn2NC1JVgFTCS1cn3fbKXv2J+a9l5QdeTg2L++Sf582VppCvrVkQPx5LvAH8mV
rAP/vfh1aZxNS2E7G1qznkADnPE6OZRSUmCIxYxwyIkcVKkKkHRIJ4A/ITUz+RJjiWZHWDxow/+s
RvJRzYgbmOy7IWD/CsKfFZnsLoaglQBhT72jaO9jvH4KlMp+/tr3bdfpXw2ckU9CeSOAzPFl03VL
IYXCEHmUv2vpfLoFTJGJWTc/JqYO4jVH/3OgZiRnu1YhRQA5kdX7YB4HlAjLJ+WknTybza/AN/4r
YlkIMJvjtFjwQct71rX6O93iz29bReeAr4ZDfLXN3F4ZDFFg5ukR/0MCq8g1gudIf+m5ZhvbUZrJ
sLTQ4sOAUPHuYBpqi4vNY3MBWVdCAbRlBdhZuKgr3OlKng1GWiYkwG25rpfV+yHuuU20FZ+YsDnw
AKhdXKZCcPyL08AfToS2FsegzyWwd4+C/7i0G72BX2HZJulzRgbvgjH6wKIoegREmHrnv9mdfn54
3qf9pcnGWyJ3swk/T3MG7IADRhS0sN5+O/uMn+ROUCTxusQ9QkLigonsvFSkslXPfBrzCPDCQ6eH
Y7zWQ1XT/aoYbm8wk+0JpblOeLdxBbfr+ckvEmk5jhvBZJCLTd2UebVQLvrI01FyIx8bbfkLdaSJ
9MYBj82EoBSQOnJKaypSTx4fs1JgZ9oLOq/sgbVvTBRBXuEkHoDdewRgAKTSZk+fQBTXbqGRnu6B
HKcXdFFbeebVj84JYoHM3EdejHtfglxqABhB+EMlJrv8G32OWQdDTYUf670satImfyATUKYh74+J
YJpwc2vBHgqI/kbTMHAM6p+ShswJ7/FNWl801PSNLO2bT5KtT+ZSQmrkHFICc42iMF7MueW411Yl
NoAD/I+DtcHWkB2X3lM0HaN+V3pn7tYHhULr5+BoMmCL+5HNv3SDNblFt6u7sPhGJ9JDDyqhNgg0
EH4aN93KjHyXbDHZFNwVJ0PrDDmp2//mGR8vAz7M9929Vjab3WHN2S2GqbJ5myjfn0zlVAYGSY5D
Df7Hjeko4WdP3ikQgtLtiq1/sudnMnksckiDFYzXgiE3CjSgHolvMQS4jfYiVtHwt+OhNJIc3wzt
7+rrDlxNGUnb8opMUGABFb/v/Mw1/9PfNBp+zJ3bFJLuwIAPzXuT67jDEb0PyOT5d48JqBjMZW2f
640aOcAjpJ+nwTEN7xvn+uDWSx30y6QZMngq1ciDHxkmImiBZZoTVYhCUBlhTsngNnTuJHUlvTgf
/nFHct/43z4h1Wx71AokFAmEzqoge+RMUWGHDbEb5B5CkrUnHg4R3nVI2/GsPNXpLmnZm1wRK4AV
916xzHB9ghCqjRhtSNHwkjGRus0c3l4msSamTY3pcuvxNOK7oOmFnwi4M0lfkp+42hl0s6XUep5h
4BlRtTe4MmjAm2MRG7520W94k82T7NUHdQsp3mFs4zoJyX3qpdtS51/RdEm1zynm+yO8tl0lFhN0
s8xhs3WjCu0+SZWuzQZOXZXx9Ytf+YAK0OyBwJDnc1CjemAWfZZR/91tWUqYijxupb3npiiE0fpU
b1I5sZud1fmBsD90Xb1QgnzDwrxyM3Is42eFsoLEumnmQMc9MucMAV9gCXaIl0g8fio76sb2p2Tl
tNGY6sYESaAJJ5hKZ0VUGaPnecIaGnbKJfYaEjV+0eneYCCJDwu3NUqqy3dGsv0vB2yhBfvIgdXz
0SQJkxqdmWEfKvhDtw5Hnv9Vi/2Bh1rerJrD7hpFwJ+ze+Lou12Sgn3wtDLHl69xS4K2uwrl1FRM
xXjD7mGZkTsqNvYKv3k+ZKsv3j3z/Hj4xaOTlIgezIODALnFuPDFFliVgoWLl2XoFbJvlrZRtWcw
1Opcg/OoRXHAR8glgPxQ3xkmhtQo6dABeZvuRpcu7wjQe+Nzx3N+4VGK+OsXXA9wfRjAbTaXhOW5
503lxxUr1dzVf4QZ/LTRVpjHLVPlmaeMLO1aD58azffY/gO9CCjFFo3o6XafqElHmbqfs3n3wn9j
2TZPbAZ2ESAW71qWGGWmDkHcOLZzfv+IrBJMHZZlPqm8Q4AtM+zjWzyJrw/iQ4Avmks49N5yUlIy
rLew4CtNTEnpAwIGlXjqyptOlQFgkcElZz+aPBO3I7toGOUnwDWscp8f0rn3RUzcdXOINRs/Qhio
K16QY2nQbJmGdGdY4+Bxef38Nj3s8kmi7JlSbC5YtvUYIdof0sbwEyZJTKV7XNNfEQU9NVI1aLrN
G3e5mvJOCpnv3BOHwR9DixOL0DCs7llfgLvivECAmQ1ZCl+Fk1IjK05oQTRQqxloiFxKS/sWMUUG
/Q28FrIevVfAnr6fR/0ltdR2xLScvBQZZp8eXcOO/41SnwESPzdbgM6VeUw5y0VAGNFbXceLjDTp
19LjzpxLyQZ1SPHuid4O8fPaZkDX/tmCvmBDiaQU94Gy6fLTAUsRt1ju8uADGloJcaH18dm1ySeM
G2VxASGCBynh+X5o/KUPD5yqwNUilrnOVE9wac6Gn1T+ceizO4GqXJnedX+zr4JgPlaSXLhkN1SB
46l6CCixq9upmkDvn/84xMEjsghS/r5v75nLgBzyb/iVsYC3A1QXIISFR+HekHzh1WLup6Mp7J/e
wltiPiAhbwnL0ATMEgltysGKMWsRhZzYVzhPCdxqIpYp11/zoNU/aeUFyYGqoL5Ps5PtJWVtMXoD
YmHIEujHtCdd08/hwvKcVs17bzdjRCygx1sQla5zXgGiw21n6RruSDuXbcXV3Xgi4RUt0OrWrOC7
KEklq264SZic02eBNLpzik4DNAKY+tJKPwaoc/Yz2c2yLgGpx3Ei1tyQV7CZ834+Jfy6w6xCwaB3
dBUNbOqYOGH7Ox3vTyACKAdHDPvxED7nCLbpzNP/7uLjHTM3gSlH6TIj3FVq258qKeUUKHPN2RUY
qUZC77LUFDNwgoaD7xAqHblGF5dwvpt7wyeI1TPmeNDBD0dhPqkIIcYKmjBEmtELWTenwZRQwmrK
Mo+oS6oz+ZK89Yw9EtFiEatjLmEu2PmGKCbLCcOfmq5fcDNLQqEVBWtBgdhE2YM5gU8UYcVWtyGi
HKFocqWv+U/p/YHx+MgA2yvc3Hz+ONVJ3w4M2BnVjBU8k0LVTWCUhiQHKio4tvyg7mKOG1sumQjL
LPlZgbFUEpypIiscfotqkVAoXQ3Do3mt2W53Sfstp0AAZK92dQC2i4uvRr/KqcyZz4SOnwXgjrxx
FCo5pFhAqjoQ8s5pHfethfMjTPGplkjQfdf5sdMjLTepaZKvGnDv8dZQfIP3zwUuw3b0+4d5Ys9d
KpW2KdzoN/INVALUaolHH0WyrKBWZVHnsuCaQjQ2z6M6/htMIzukDWtHgA9DeDiTDIP17wFLhYZb
/mGuEjxpExrDNShmE1AhjDDlrM+NzbrU+xvENNkrNjunOtkKHAATkpP5B+0n+s7Pnmj1tYd0BbKa
hCS8bMKtvEvdQKy3Ia9Nshnp02XJ15VI8u4PJFJ2JDoM5pvyPXrtr7NtTiHvEDLYSODGBo/cPIpF
DuyRVsJIQNe9YpPgR772eV9JtvjjMW/NVTfChIDc6we+E07xwx/L+5KzLXJzr4BxzrJJzcQir9YU
Ra+0cwYhhr+BpUzeTGembBGKwleET4iw9SJ86BBzfx81j6bIm5zdsjhw+U5JXRek4SmPj4k24/me
KDzCs7EDxw1KN3xOiSmyS0Kn99eiA4lZo/m678xCHk9SQLO/XHQSPrIklBbwkQpYg9YeYXwSE5hB
FH8ILEQycX9/2NYtyd2es23yEprQXPKK1DXoX/vVKv01Fo8tJQ+hk8imziqrI22TKcvaF4EgPp3j
/K5wLvWLb9cBFpGrzh0TwbOsz61zvOoxeQ3b0TqI+2su4l6nFFq293TgZvcX/wm7xvHHdbVt1g+R
F7NJCt139etYnuoB+avUucVgtkVYIzfpgcWtsuwVbZOdlvv46JHEbgGMP+3G9sjbcV6gv0/nrY/v
kb8Nt8fa8UbCyNtQ5JlWj3M62a/0/1ooJiUTTyRkp2ZenE7DuTzuu+mIzQjcq6SbyH1CAYgrXBQD
cKBrJu4dk6F8fSJ3dBySJ90M3s5U2VVt+I6zohEtvrt2PG21K2Qcjp695zD/gmk74w/mV/4oEQlS
zgYJcFbYtXzApf6roxT0q8bTg9NjmQrGAktfuHuiWdMLFIdQ0GJSjgrjNMFDn70ot8vC3WCb/NBd
LTISBX89vur79CtUb6L6UNk3WpKxh8DJxjzCG6edPawQt8sGzEgfNgMznZTyBObGFU2Xe3BW+cO0
5VWdEpdfL4XIar3T2qUn8N+hSs+dr/A2l/TLV5lAp/w/4dMoZ9nlFeJSqXWSd8o1kCZebq4rjjBL
0TcIcWEV8RL7d9MSMsjT0qIMRuJOOeUwXhXJudek8/9cH+T+JG1fd0nMIuA4XyhZEIEKFUWcn00D
RSbcUdtCKZ31He4ySqP2WX4Z7wQyIUiWEkGX8UlAgXoTUU+vnZCMxwsJlrRG9oQKhH/mIjVZZPub
7y5yDb0aj6XBzsxwu/lu4RnqxITGF8HVWXYovqU+8vp73Bvqo9UB2m2XS0jCd/8kRdyryhLbxZVM
piD3Azg3aE/FXYsP5yidUdXDw1kUqn0xCOJEdFfLf0omTo62QzntPz0tqhC+bqSQXq6K1MoWCnnq
t3Fs6FOUP0I1jx3DWwNRL1rq5P4d0qM7gHaVwwrzl0RV74DTSUovRkfG4aIYKDHytV8Pr9d5N5Dj
U9spT1bIfxyxVozhXlmKR/4jrrhYOIDasIJ7G5MZ260qGCKDolQkXXGyof+KLvsCtleSHzwhZsNm
suwHVzuX0foSNWZ0SXA06S/U9WW3a9tzpk1GOrWi5kWYEiXAbtMlbHOp5S5A4mOmpOyD1dY4wc22
G9igEFpCDaufXGQzwOcv2b81NG2w4rNCSkUdqshPkTcol1Xuk4+hgroeScNBvD+eWYmFOsN3TgKs
AyjrG3kIF0BaQsaRbX7AQiGCL+ScK2fPE3qssVwEMUf0bTklECXpC9WCBl639fa1I6nPxdZ1lmdV
LcMgg1USlKTbPHl4hjBm+siYSHLD8tBK+xrkOTcd7EyzaL0Uj2hQIcQ1znMG/JyttoHK+hvoW/0Z
y48PHEDsAxQ/+as6WijOS7o/8nB59QNonaZsCVaI9+mDYZ0baVoDnVKazV1EUKzETUed1aGPQ8iX
sHuPOVI2d51bK1KY9rx8V3dIbKLFSpxM+g7sNsFYdHmfgpsaeGoozzTqDl25GBfKxeqPcm47GcSE
1SyX3DePyjpBqvnR53s4eJNAghphFYJCpmLC9zqYHVTAV1NlNU8scpnNtPG63wA8FjFK9P45t1oS
x+wjdeFZ/W1P0H+jL8udlIQ8O5LdOn/c/mqG5am/jZFn4Au0k5zRwA6H0vWni3ugDSX59NkodEb+
BwzsDEWyd3Btjs3znnubV21mMzezpHU2STVV7Zmwn/JDaQyr+fpu1TgVN8/m93zpgVHwzZBNHQBK
mVXvFqRFb9w6mvT16oBs45iQ66yrlHZTJaexTWVNcpU3MWWW7Rcj6ygueyGBC2ryFDefIqjikf26
Pj0oyhRFzjRzbNtdOGTwNjlXD0CiNohY7fnQWxcfqq5KO1XfKKA/AOd3pG3o0XgzxJv0zWbhDcz4
0Rm/sbL47Yfw1oETGT5HtwPFi1MEx1xjB4SKF1NQnlbzzXwo4FXSUOk15FwQGjuG4OXl3uJl2tIt
6CurNCsL3HR45XVxZtsr/KiwVuDztN/PM90PoyZXIOWgo2oJeCzXN/o9hX6bUcKD0z7EbLunJ0Qu
xlJG5kI7K5drHB5grcFrpxJzGCapDA+fZQymDQ5FyefSQjmY+v4bn+Zb6fJIYN6E9Zs7AF09If6z
chK3QKlc1Y/P5Akqm53Hm+FmbggoIxN1ACY3xBFN0G5Dkv6WP2M367g63WXU4XVtGXMUBlyuEaZQ
CDcEpKmE+wiFoNwuJ3xbLQ+G740+/eJFv0B34YxPnEpUTieD6QDrC23Qdv4Tp2kSP394Y9JxbK9i
tUUN0CuErN2z17r39YnW+v35QXVYGXQN/cAwNd21DLt/JxneYy2Yyh12E3tt1Gee4LIThoi52BZu
+xqFgp9+jP45C1EdZJ4QbVUISwNyQCM9FpVnlk+eZLkyIN1oaqVqOULGTOybAWDSe0amAmV9JInx
gqDdgSuWJeZkGpV7NkC2uTF8VkE43Ku/C4NBZWKlEtpn0BrQDhuDgPWbeo6Tmy/QNdA6LVujNrcy
eRIR7B446P1A/Vn2T51YlwEZEIgewLoK/oYVuyLu4jFrDDoEtq58wyvgdk18UoPk06S1MRPIwAHc
u8qWbkbP7MH5CA/U4ZlI4/iKONgyUi64oizkAGIhYE+jzr+qRUlQfck+2Z4cY8NHc0l0IxHGVMv2
+hCbyD/rKB6j9D+9H1kpTqqL8WcS3EITEULDs9PCB4mKZQMwvNY4ArDyvXQ31hvP1meT9PWhcKjk
++jS4tnlNILNXbcXNI9ESbyiMuS1guVwXIg40Dq1oqAZoMGIcGMzbQzPOXZJC9wYV7VSUtFdFPV1
vqNnmHEva9RyhPVso2nR7WqkPAEN4MjE05hXH3OZ5qE2q46crW+dWG0JUPW/9r27qHlzMsTRstLi
u+pgfAbt5+/mY1KCuTchdiBahjMB9Xtj8/TztSk3x6IxWMQtTpVwOQ4E3LpAx+eXlMBcjZMyn4In
XkEnEAqa3xORPDylc9PLYZPocKcPnU5xIhyQrBssYYqXZ1lybmk5JfVdYTbfjzS+GwAXtaLRPTxC
z2mQNvvsg9rQvaEESDszfNPPYEa01iMCdQuk5gx4iD3+cs5De/Cjou/RHtuQ7RZWvKu+97M5XJW/
mbNfSljLIpt+sg/2XZ9bFzbXp02OZrmEweq0DKz0DKKdOLVq777vSmbJP6qL5+K6E2PdcxIZF3Yg
+ksAo7rWA3Gwy+bSyZTZ0YV0oPy8e4olA9dWtdUGf8OzqAZHUirpW5DTn3sKgjCu7Mayp/m4lD0s
hYYL/fcHxY5FugfJCgoOJC39PWiw+R0hXQDH/mzT3sOaJA4V1x+m6i07IO4GtFUz5npgZWYAZV0i
kMQ9uxHNQM0TcxKG1++gLpvOpMGRULPh9oZK7k7Mabw2WRLwshqa/EeRFbgBXx5DzL/nvRVt5sAQ
ENMAuMo6s84b7lSqJahSwS1wGw3cTv2+3Y5oF3edITO2XmyJs2w+ws7SWseZubpSO+u6IQesRTkQ
sscgpk7UKldNMYtL1ufLWa9XlBPWeH6uKuLSaIlfVuth0u6DCwpNHujVy8DyBnUwAL/M6yJ2sjKO
CIaQvXMBLW33mrvlEtYAlEWRyGjg8MA4/snc4ZkAdvnCCpAZpKk/3VZiN6DhPxrY5EjJCYeTaDFw
6XfzomqtQuRELhnrWlPpVfm+X7NVWnsh/eaUo1p0QNWGTzH/+he7IxLEX5hqN/F/Nj7Zk/SarsG8
nW6ZaVHmTQDg5O3OWT2V185UYyIZiHwibBP3SfeMnThyeBaKHRjFtaAaacTXN5rJPPHFOxDg6p41
LrYO7ikdmDhMUkvpeMGjxDblow+p1IJZSlCgm3cDeL2htTwTNmY0LatnwjzeUOP05pBCYhl3+l3x
JTTUxRsHHZLwamq6JtcDFfE++2xaJlgT/Hy7M0Eda0ywr0M0LduP09VukAkbHPhcwOvn81XWZEst
6PYskSHLnjOId1T5rXFRgjqiI3+rGnDvbGY1Twm7XWdtJ00dgmaQlPb0tlvXJyegzFgcdYsr0DnX
7Ts8dq3df2xIFAAcllNfG/WpyViuB7fYPoL3kVBHBKM//Pr6wyooVRPBTVLCVRK9f8uyZFN89Kba
dMsGC8L7oNfIqM99dt/Vn2loLIZ37R/SGwvn9Xhue9xJjmlRH3ihB3Ze3buayYw9SQpKEUgQqic4
tIWSn1mdHXHbjLzC76dXYKMQckPSvGduCl7PUD3+qZ6wLR+mHEfnnWPUcHEIFvt0GidEtCUruLQo
Om/x/Vnp/f5NtTNKiVv/Pc/UzKcPBBDng4yJ7E/+quisC/ADEgyMpxqpbFLNoKv+GMWX74VA9/bs
BfUXeo0WJhC47X3WPi+f+/n16DpzhuD9RUvlxDuFJMWG2Pn1uAEYp/Pz2sAMfEWsMEyoE3cvTWZy
chKUMNkdHDdlpjgYEudn1NeVArXtDJFMdBL4meFmkGjDzws1R5cJMQURPxy/8ib0pUmPsg/+3G80
4+0oNvDsuWUrYfO0dlMRITmfeNwt7pbc5Sd8PfNOGydmR8dkaO8uaPww3+bigmV2klAmVILCZMy9
C7aA2IE490WC+5ilr2xWgkm5ZhZjZgcuHeONkWyL5KZ1zjC8bonZPRITtS8gjIg8sR22AyXANQKs
D3+IvEfUKZwFlf1vQLPcRtu9xE5ep+DO53VtxBhX0gbdNENWlgxn1u5mhaja1qsGwbdp9k1XfP95
qoXDoxi7sN6tBbZ1Aa1ctM2R0ZqyVZs+EXGETF8hIxUkNMNJzoNAmbVxbrRKePu/q/DUP3Ev35n4
s14bvJYPg6AWChiwPEIWOtYDYKaeQR02w0t9hL0p+jPlwTreVUwcU1FVbJPeL0bAMLOEwmMG2C2+
ilnKYjARqW5O9b7ee41WlqfPGyHGZ4Qr7QqBCxGRsYVx9baWsfewpTd2v/AnTCLdNUtVagmduvH/
JzbzGW1Hz8ZaZGnHdZSAr/XnH2ID90VyQQmY6Z8/1Bd8XBmG7Ad/qZ/MdX5d5xHfSWtPAIIi7lTk
SfgnJC7S+6NLL09rVNts8Vs3NAi+ubkXYeSfNEY82JnVi3GM5IFsSXL14lKBHjMwMi724vXjzCOD
4k30n+iE5QDzT3QEXlCTeUHxdcaXhlSgezKBtfOYdE8c2i2m7HwCYKlLDZvomLbsk1Hh7xKvWfOn
6XWgUSsqQ8Bbmrc3K7FUw+BC7vqqwoGHG7B4ljJASdb3booYZy3ZjW6tTpmZNFVxGJGs+qr07aiC
Ljwl50tEjWabC4RVQVZOUWOeNu+Z0JEdwcDCpw0myusnraUpPe7pXLrsMSagqb0httXHTTQtMucp
9dsHxsOv9tyBehGFlyDO29dnGOPOipMVeo19aSeqHUD8BzOUGa+91bovHtLxdeKdtAz7Hsq9tOYv
z2e27TJpzvFjcw2Vl2mVeaUKgYM+v0Cdd/XFb4OvBQMGc0QfeVYPQtUwy96FAhQ9b4w41KBfvKkR
W57OxplPKTrHmiynGnysADL7dTh+AowkSKQwEo0Nh0kyQrZeVut1BQcuMLJSUQQOUOgSsJFa/wX8
gPjo88fHH63jxmiyjc9/5+lmnWv9LMnlezkPscZSlNx50I3pwP5IipQddwujjkNFpH4KusSh5DjD
UO5lg6+hN3czPjQVGGbfmuwtn+NbdjqUeIRDfgPJerZ90r9ZK2Ixli58RRQuVgu8PLFrN5/O/eKx
C2sS2nHT81gTbvYfEkuqKupMxy1vH1hDJe2yGwwznrVElwOX64zWrjg5IOlrZlDZ3OumcGkHGlQk
6mYZYyqt7f+iQUMqP38BOVIuarOx26WjpSZLtpvD6ka3pgxYkPDweE22EnbF/V1U0aPc+vBG5CfI
xl/oLo6Yk12XjyIY3XQKHpA945/1fqzlnuAJV/kIweh/5+12ahD/6cPzoXGgrjkGB5M+LuJ9uQN8
uJNSUmAajT9KRewz1BfYnypP9Lf9AQh5EHurSw7XHkvr0VQ3Pg5zCOgCd07hKtXxP0p3SnugPTC2
4OiQG8D3VAm29HV/gkzHEOKayUwWXo3v3R5nWOw3bjLEfO+01uvBS/63IDd5x/c6znhDD19S05Rk
6XhuSJjUNXtYXGngx0QuGqNwgEyAK8ElxkcU/bCZlS/vnor5ghXhVELcIVTs0tzeL2yefZiLDG8m
HJoXaXk6ssF3A4QLm0YmRMYUN1EXTetb7xoa0IfwTLPmKG9gFA1RZTgjWfxglhxW87FMb9pyGJzK
XDLHoPu2BJqNufanmtdNpm9FK4DpXfRNodfGWMSjM4KqgIeYrAugQz2kJyD6F3++9yrVQkDBq7tb
gwV4AbRlpukQ8OqrMp756X+KuNCyJHYjf8q/VTIKbsXi58OpadQiY02ITIC9PLk7slr5MIEbDaP5
Yw0w2WNQUmauAQeNMrDUMqzGnHkBhpSoCPSd9yKEbwlHw6QausRLsBLf8Sd0wAzwUI27fM/SISQu
UuhCZKDLFQ9m18USvYECA57Mygg1CRxDxK6lfwj435hChuUIVovDEAMvLnz1ZQkhnQWIJkaAkfle
G+Kx67s6aanfGSIU93WWMNjOJ33FIOLWW2jSATsRUkpmmnETU6mQlMhdVkdyJFftGrHp7K6RdBGd
PE92VulIkOoezNaAVaDzpqPOTg3qxQu0Y2kh6fa4X8Eu0079lo9olY3mOFpHZHzREoxSxlVGRXOJ
KwDAkID3t/J4hVh5xs837REMYU+Ogqk7P4SrZ7tCfY9JitWL05dfD8ExDtC8w3Jl2IZOwIKf2duR
0lJX+u6HdRQt8X1RLQtv+RwhsWDqMTMn8oA6O+m3aPhdemPLCt3forPCfAsDtYKIR+53ZMi6JDqy
whqd7eT44LK5n6ioHPwERMDbQGzSNg6Z3VBfHK5iSf0aOQDpEmEnXqxU1K8zR8lrXkmXPfBlHEeC
j8ZpSLyc94SODTOkUP1qINHFabTmsC+18AXzVBvx255AQLn5YqN9/wkTHxEEWqWXkSILJslNFpsU
mmnEFbm+jN+9rN9PAYmf2YFsuHbOX511l4QHDIZme/X0eXBcCsELM7j8a7g47tvXkEHRN2Chsd7S
grmsy/SDXHOUXwTPsWq8s67iBNgZz81SELpimqCis49CbOKCWTFj9HamvIOYJjz6411wzqIGcmSs
ooznrRPAzBZhPqNXh0KYl5a9GqxFtbCBC9+Q8MGK3Gy7YxP1Sre9PZFuUQ2clIs/2Xtpa/ws+CwP
S6Y8vIh8gLIjAxF2PRaao0iN1wmJC+ENg0DjuC0lVZPzDXTiL6573uStHi2sdp1vyPGdyYinsx4j
AJLabsOj6ge+b1/0JjJOHAYj3S70+2IwgXp1UgfJgqxEUWx4Gx7148BdhBbQNjlTh0m/KUUNU9ru
l8BaQQohHvAZLziQEXwN8iZOjiCEjQlZqiAub2pcOD/SWxkti4SRRzNtZXTJwLwD4vNvP1ezc8uT
FO4eEPeKGxtTsBtKGamg73wrCtpF22qd8MivI4u2Dz/RGqT+7C8vPTRGxvzBMnaEdX8j31duKC41
RFNHQBq8cfvKijm8xKdBeS9HI8xyfW44CfwwjvI6SK+xanbvpb0p1O86Av3s4sEmnm6/U325w7aY
IOf8GVm/xjx4VliFW31DaPZPtDUZ411uarfHCe9FkYbrgruxk3/PsB/VOJ15riohQaZcdn1ahp5+
MB6L2HcG0BNwA6Eyp3yF4YCcHlL2FleqQvu6r14ipoV0Zr5RhPkDluvqbOP+zxb4oONAklrgCTiE
Kql+aMbtbclUAmMmhnN/NsQb5uNGPMq/KStADK5bDYRUr08cCyBN+00onyBIxvXdWCeJYpBj1+up
AyTPwSO5H1IX8fx2IKwYksIvPuqsmpDjnxZGbvTrsCaXEatrZpxs6SvpQF+lpsFfxlxnYIFCu4x7
jVuAAAS19yGQE8VznFZi7QMGcXLY2M0wyqumRsPpWyy9V2qgD3vK4ZwwT/a/wts1BNCCzLSMN/dt
JS9JiVckppjdtcVJnEEoX2qVh2z5G61WD/plZLQdHTx6eFtdgTxMvI+xpOq37jJKTBqL6IcXdOOm
VPz5QFkl3oMXGwNhSEcAt5ceUn1JPAmDdr7U08i3C+IQSrgGBqZ8PPHrvzJ7vAswt9jLxG9AkVR7
ADkVJkMg/s24NR8IwJXSk1HzYZ2RNvUCKOlzl29UojYZFmO9az/+uSAU2zEFGEqOvwDJl2dWfrQr
Lq12B5h0yIhQs1nr1LoiEvhG+PmDRCspeIQyuo2FtfyZfkPQt6N1qF422ZJj8kKUTnOc9YSi19ja
7pmGtLSKBuWVAgA7hQBANAqM/eTwBYhMKw9/eqb41fxEBXVllC1bzfulKD0E9QmT541PDQIoDYs7
oZhU+euGxbuv8h27A5DyvgIuVaJ5+Y4rbd7HXAvQh7//pCgPrN7kX42HOMLUDeGWeKaugK35dpQI
MlApj5NBJFWtx4d4X67C6mhB0u0iM/Av5rclWvau7u8NRyF6keuemYtNnn1ueTILwIqq628i8Tv8
m6n7oSvLC7C9FcrVw0J7+zfdEt9Ojudg6O30pvdtNE+EeuKMZa+yv5/T0iBTvuyEjka41a8sP6l3
/Nhfk28mhjaKQOtGah0daCWZvgIB0CmIBW6gUN0AXBwjs9bYbe7ZawenSrVnBIwHzY6ruq/gB10s
j21ULKqv+tZvRHxecMRoXBltJOSY88MmV+AWklxUVgnVruJ8Ug+DpqRQcT+xEUX3W9Oyy1EJzZjh
YxfSzj8x+iw19VOWtSzBmezl7YzJ0vqj1ef30iy8p3eOEyE+STKPlJ2E+428WtMnH9IoS+Fbc83n
p4Yru5Pf+VsXoLOjPnsopB8wJhbvsAgiNLcEockP10VGWli/y1WetO14NdO4/eRqKFMUJAon+cM+
kkZyJIpm6+xM9NXVJHvOASYCPXQIDRqMReYyU3YYtGCB6iKz+9Fwd4d37tGoTGtpZCJ5VUDhX07V
C1Dv6ZALIhrA3h/dlzXaZHm6Zl/nxmUrLpr9CYxxP4vZ52GOdr0MO/hVD4mK007PzCM5ljsdLkZF
zuNd0NDPk3EQD9GMB2neb5UtwSEgGTY3KozU/7CvMHwDPWgvmfXiZN+vR8gRjZujgR+iS74dxFMQ
2FueisI/miM8uFnOHquap4HJzQpQtojXBrx9cNZBweGC4TwfOkvLENaoBbS47xm2H8FQWAbQ8fTs
AJ+B0cxOLDJueAEmTT7CMTmx9ilK3OiACNGlsU8wzkLJMAqy6azFK3Di0HmSnQC56HDq5LdSWAGs
eb77ctb+6k2DONbtSH6/Bk1ErNaQoeDVWBOHaB+3ix9RBF2In0A5c5bQ3rzqiS/ch8A1jp6QaHUn
HpAkG9MQ+pGhzLP2LCGIMYb2z6eEFJVDW/qtxu+tmmgH7IDuQP0EJwDvWGdY61i6LTOl4HyFLkKQ
kDQ++OAWbIB2Czwf/PHy9Vu/qSTkR/a1n5XSJNW6bmY26oWUjbE2qAtjVBM8XAZ11Hg+TL+kLDD1
QK1qqzx7K1mA3A5yr5xrYsSdWbYa5CHBNyRoDji6VpIZoXS5kEtmx3tTWmk70BTc0A5DM+Ew8Rn/
Fh7HCJBpKy/KY45kyKelo9DxzVJLDS9WpEF5rFOwhgkqDq5yJyqkyRthQJLcSGcvyg11JFiej5hh
5E2gI+ImzzkxPzofLoCm6lk5UEdQDGNm9GRZB/d1omeQSZxph6bGJmHHdrGiCU8WqGltWjFu9SXp
0rntKFR+tlUVDJqTsYQQyO3iuS6CYyFXc5oEcEcfQngVj1NFplKUjTeIDK3ixf6kaCQ56AeaGEyD
roWAblNc4lY+uD91zJfoKOCdjiuKZ7WV9IptO7l174hbrjhKzMvQz/llYzgLq1eqqSzzVd5k89ZM
BJtNwkQWFlwq0ocQzfX6sUSllhoeGZs8WUBqq85NZ6tWg6bDzdQPfmiztXUo3hZ8iTxEoA/JeHgq
GAB5ZaZ2lDJxKKrFGZ3grUA0IJ/zziKOiMq5eTfxeQNXSlaSdXa0xPhQHtWXhQQxy4TmgtL0IqnE
AbLGDpZay9xwQ7kbwYLlyld/mf/2jxetwZcfsgtCFLHbaGv5EsWCdY2kukIX37C+wvLIxdV6Dk36
F28mMUUFSSZdj6hXbptEwt2TK0oTu9ri/0sC0uw/Ou51dcve4mIRcpC6qYZ/oIJwN9ZOLcUioCiY
kOiQjVqzxEv3abjABkFQwbjs2e74JyQWuQmhXJa8LUZ3Fb92QPn4yaL9bYvXDP/sxJWRagVGrb4x
eMtNzMWYGe29NZrK2BgVTTorG9NtWnW+hckrbMlSv9LFl7kxRANl/nqbrHAdMvyoLs4mhwJXf0Vp
s6eDStWjI7uV33SR9S/h4vvDgFlMNmsJH5jqvhEHtQflZfJdTf0CLRVZMLdTK+qM7FX6Ef7zKqzY
QHMloykVBAYIpdFXm2KdPwStSG3+wP3atrwhawbxXoSC4olrXjq3PromU8eFkLQXE9kbE2HptXTQ
cbrSm7p3SY938mVuvd/sN/o8hLgoHxuYWCBVPQm8TYa9rdygssGjMKTvRtuCTDQDioo6VlALVeZx
6wFzPzKi2zNk1ppNR7M9C6myVUUHR7JV63BEjRFxhO5cQfXOHcoxo0WgRwpwZl7iRDLnuO4RHRqi
B67iO6t6yG4lMeX/iwW2nRpD6nbavaZXirOr/pWHT5Mx3nVIvU+7BOzV+JFQhTM9UESF8/lKI+wF
uMlojXzWBmMT3UxRHlsYSBrXsGCek69SHmEElwnW0xwPe8Cw3FaUWek5JTpYuMOfrYmqYsRdPSG/
yuP5wUURsMo1wRygFfPkm9UNU9Ts3LXOIymfCeUMMJPNxMOAtxlNCTNLx9/i+/4aSbNkgAojtvtW
2i5gwnicz4KRt5Bop59PciD8MtZ6fZZOwfaHFjVQeJi9FK54u1WtbfNtdqx5ntWuOcf4ORwacb/T
ZPBIInHLgczmYt4oCdpkVFBpzLElUyENwcm5aryaLaqkiObEkC6/7yxkS/Hnwp/lG27MySD1fdyO
GhI/qBTVgampOnePe/rDnm0tV2m9JNfXZw9mI25kfE6Z+hdOd6nIoNDh6vDyRcEfaVB4tMs/WQ2p
GebkMu7xhv+kPutsLkgAT4yQEQrNJ5YSy9VR+ibQcb56G1LFlo2VcY3vKvpcwJtUHNHInJKSBmgg
gs1qGHsa3/N2G+IBw6iefKr3JkVL2ksZxT0IldyYc+5ev21sYtRjWtUtIefQYwmny+U8auXw+yf8
9o6ujQlqZYeiBEFrmJThW9dAU69iTlm75dvB6dpyUJH5VN+K6z+DEsXT11GLotw5wCe4M3iNiWKZ
R/IS+pE+uunW112MDrx5go8wdC9X9LdWcK+HGJ772BQkSBxrKgTIULGCHWa3s8m5ogC92zrJytY7
zjO1vu1bXftLWYxk33YGsNDGPLELosFJz7oV24c9vnmKARqnaAMU0CXqCduJ58fMWEe9EFFIioKr
NZXqjmRNHADEr0UulfSmnQxojZI1vlwszBx2St7it2pcKcvveq+zQCLE20jFkObU1cArc9bY0pR5
ro0q7G5zaiWucY0/Y1QGnLHUPeVUDLRTh70PHGi9/FNesuHch59GbzWxBnt/uJCg0MJjIats4dcX
NOGZz7QF1yUfepOq9ON7p7USf4qBq8YZqxBKLWRVO0WrESn2EDo/phcKv2Q/SCMU+jh77c/pHSD3
hMIfOSMdRMnHyWZAubN5Fv9iBji32HAjCzXd3EjLe9IxC0HHxGpJuGRKkaeZf24gpvzh/ViVzbO5
LX3IaK+0QSrf08XJIPFMydLu57XbOjKMuPjLPdn13oDudI0ztXciSBstMe0BT17A6tkH5Xbo+a//
A1s6Bkvg1jI+l1yaTINBDVbEq/v35OtdSz1Ax0TIzyMfe8VqLuQs5Vbc3G6SlMW+7iK7X+vgqdvH
aW6BMzNdKd93TXVa3hqYZlKOr8kUqM+CUQ7PK6y8hOdInzuBbsciwJKnOm/cKCzvkZcCOp13t5To
YmX4Inrz9h5iobqMl29HhJ4VUSOcRdnNmMI9UwoDIq58bsV4e8Md9JS2FofELYz43s2WJBqMmrf4
eoNqZUJ3lxUKxQtzVtjJc70Fxf2ayBzwX2vUDteKStX5u2bgNagsE1VDUI9rnLRLRmdtUWIzOvLH
3XwvlQRyV2TNvsJarsypOgBvFNCnrUXUTj1n/mQvoWNiGOGCO2/DujmAwkxieZK7ZxisFpa7l4yy
RqTkXyc577CUakDfyu+xZ/O5XV6S9ZE4B/niKey5FQuxDCElkFePUg+m7W+5DH880x38pvXU8eDo
2FcEERyub2+PknFRSZ6G794ydcCvQ9FmNSb10GPg5Q9l6AXk22ACOT10MVf3RvPMgFwjp/PjPP+t
uEx5REMmjwkiIfrRyvgl7bKhSL5JvOMs0/6PvZ5utW1/bDZJ2l6XcFPQcXBk5WwpxcJhGBsRjLBP
YxI/NpPKcm0parivJYGDdkG/Q4FnRTa7iUOWOstMGKkOafCc1vmuxI3aZQZ+wLgHdOgTbtmQ+NTl
9fJbk0KdCKVzN43cLSCtHnEm/taFs6/ZAIUhP4+/O52BcCI321OybauDbrsUoIWdlUWEVUn6SDw6
h8eJtpNY1ue3eZlp3sAji918mHsAaj+IVKzlQG30jIf1XBHvCCaw3U19R0XZ2pRYs/VOVJA0v+kI
CgIVDfdfJzuiZ+8+Afc+SFGe/+KNrOnJPG8uaECSh17VITtWXAdx60t29jetLmIDY0tGGcyyAxsC
5p7zKvnsxH1DkXjmm9ba86KACAzbNWFm0VgCGz5GAD9VcMNgfBq0IWIQFQgkEMxVmWUuXmJl9dGC
OlggPw/1yJQTk0UDpD9xEbbkxcg4LbwinVCxQEAGPs28yp1vhgaphGrYjknSr6XU9nTG3RnpEgvd
6j6qAbFpRjgQLmaD2K45+D7sbTS189hKalrtNkn7hw/ac7kKvNelsOoEiXoV4skQwpxIz/PcmGf6
wzDlLka1RawBRIKVwFOatT83G57QZJJ6o+EFcGSp5NP2+spjj/3Fu0ifJjkwZnSG2834qzgUWfU4
7PDxvl/b3I4ujt/d/1QDmYZ8J+sqMdmmAfUMiMl0z2M7lwNRhTtv5dEazdJiana7cn88HqAE1K2S
XpcuhWm8k2sJO+HCarTcAIeJJufo2rNLHQAbESepQFb656MOxYaF49akYF0aPVADpqnJ8qbBWFqm
/cPzf7K2BKzKyQai08othIlvK10C+wtxO3Znv5jsl9cugtjjcG1ZP31r/mYOLJuqBGUh4NReGEwp
xSEF8yTLEM/u81QDgbab3umD27mBR2MlkC5K6sJlPvts3CNyGjCqUK637M50tRZC9ZVfSZod1mME
4+mr9yLGLAnowYKkMetqmRyw6bsmcEYBqcPd5P0kl3OLSadby+PiXnbZaT8fdQeUqSlODA3QavF3
mrCO6DQDP8H/q3aUCRNqQdt3ipLBye76mBTzL0rJvIbPcbbFpMdDYZ5MdFl5eJnTp9wZUUAQTGuo
pyzx/camCEpLgVo8gVfnMCTXHubG+ZM0AXFXuKGgMgRVl6KAqm7rVDRX/tD2NbzzO1tacMstXy9P
dwXCEkZcc+WKKJFXlYKPMMKD0o4OGAMfy3VoDdjY9D68OZa84nmAQZmUxGqihiPSMcBiIep4mlRb
uocMMmcvbjrkRyNqkbiymaPIpoSKFAWes9I2SD35SA8m0/luvr/sWY4jNUA1zst+XfXbyMm/l0kP
2FqVh1zW5BNav8q75f+Tq8ehFrTvCNuDdJKpzn9yCL96IEMtU3RsTn81R2v3v2kOuX1ikqo59XeD
GUnBmCwX0ALEt9xJKxrqEw3Gma4soEP77wJDL/AWfgQzDhhz6lHxMJvaivpq2ZU684FhcL7XAahC
P7LsPc9UlXuDkG9r3Y60l7dLZqp9q6UfTIQyY2lKu1pwybN2LbQXFi86k/pUaVMSiNmMoxlQglD0
PeTm/NHCFTU6PSJvnUNHoRWWKHulaweMEHL1KC7Tvx/YptiAiSXHHBNoTB6ty3JaY67stk+5N8Mj
/nJ7QjDqz3DEZv1FIJuY30ZDLb1zzSiPA2M7nXqAgkZqXRBDh6+1TyQwtiQ3vrU8F3+v2mGObhPu
cgFfwuJsGI42d/tFI5/BGUgB2/6TrJ0YNWVx1QP/DV6bQGuYLvc/WHBwnSi0u9UCq22Fuz9hnRFL
3Q9aSVI/ZhCbmrhzhCQQ/iFN4x8a1sn/ZOknsmTsxd3OmjtHIv7nBEfUFo9tqqfNgEXw+FLn/07s
68/ZZK2pUcnz0+arEYQbGZ+KtkB0yHBT1DRgH+/tIkip+oVJfMNP0NYVqWRBWnh+HHR6z6kUlhmT
a8EaxvyoDyu+BqgwLUgVcAVVlNzIqxCtp/A2tDY1Bo1K10jHigERVPeXVsyHZynIPb9JTz+isHno
rR0U/tyxAMZ9BZ9JyIY0JC8VzlP9tAQ6w4h0YjArQ/UGBt1pyPtU6TsHW2G+xcehFXa9YQNO48si
3M5vQPhHy377Hv2vKYqh5wxqikVqRFWvnuJuDsml5rv2cOdWJLqb+dEZeZjGuWmiAugbY5CzdDMB
VwselVSgWHb/2JdNWLuyQXyE2ArcHBPNYY6mqNgqK2eCc9P9UJz7tOmzE/9KylBG2I6fDGPGAPOn
wsdo9V8sRhto6Dgpf47vCk9utZSof5v1nYDbhK3pjpiO6OjjE7BHIw6F1+YbDedWJ+HM2Lf0S6Mr
l4lNSDsFVmaAm5iUgEmQNaFbBj5+ygAwZ+xvULKTyMuzsRHBnx+IYoj+TNp9lgWarUM23QPPXPrm
zlEfZv+j5wLsePMz1K7dPpB90ePiE6OTifQVlXVy6yKwHjdehkN3RiJsl8KOeV6Yz9NwuHk1QMl4
a+0PP3dvbUfKWzmot54tOkxiY5uER5KDppI0XvyixXJw5apuBGi2K729kGKjhwTgk2o+pSfHeD3Y
UrMS4/VGkLk1tUF1guj3HjxP/5zrOr7iWl8hoFRHrfUgBuTxUsMrlXIx6HXAOutVGC7Nf4Rwp0tQ
OpYDN260YVoL9rxTmtFtLbK2TpyV5S7htht3D6Tr75KBXg6UUGXSdI3/wQs2YTe6qa0PKHb0h5Hr
kYYMJ0IyTtRcZ8S8G3XJwFdHeA1hOEf9FTmD/OSP0BSrEfTgYDaatogO9jnbaYsCIgwn1deXtvfU
UghzA3yl/r0KUalnB7vbcU9IQfNZZuTlJQL3mwa1N10C1Ga/PQr8Aj1P9cs8urAEQMDcElPXcUaL
+/jKW0MZwwV2nI37O0kSzIJkm6MydjNcPQYidzd8QX0LRFmguf0I9UxBNAKLoXvZmv538wu/0JGA
2x/b2suXvQi5qA9HREoJpgfLi/9jl9j3u3cDo7qAZehCt8pYm7+HzMjrCFV0y9KDICS77JOnge3f
NUXB4lM4YZMPGRmRokn+BijBHYiFBn2fDd3LcNJ42SWcc5HrpW5DT4kwWt7tkRpRtJaVQ4vt4iMy
rCZd97CzOtR8mOZG0Fi3yTGT7uLwJwHxbN4LYBkp34sSepWz/xsYwoV6MX1tl/Oj7Wk7wnIt8vgx
0D4IVLg2FH6stmf1G7dlcm0nET9nFzjUM0l8DXRhjsVaG/8mXZi97Ys7VCl5A7SBsneZSij7uuM5
Z9iygFCLZAJGiht9KlSNN1+LVGqgQ+xe3CeQnMqpHKWWtS8oDwAsbJvSg4DGLN5EDeLb2b0pbm3p
VFkxI1+DyPIti7nXWsZYC8Lp9N5thY8stfb2T6ArfMVXgxb2SWW+tCUd/mTV6mYbJbnrlw7fIlYT
/Px9WQXsKKGdHhn/HCj3SVQ/D1PoHEFikcsZg2zkgiyNePMLsfUEd0OghFhPr2DKWZ4ZCl8myJJP
M6wxDDGSFsUiN67PExaHcA8ne1YgTKrFBEXeQ9DJ36FMZ7TjNbGiooQK/tnie0NxuVCL1VYQChn9
RomVIZrHud9mIVHItLIhBqi2nD/FJFlA99A5EYZji3Z3aGDzxT3WVzwsCMzUdOQg5y/yyTyGVf/u
GyxUdVNjnldHcH5mRnVR6xrnAl07sT8jVauuLTtWThSKPpMuOVjL+GAOSEqZ2hyimCOLuhKD8G89
9Gbi7wP/kEBnvvn/mnbblMeM6CIcg3xlcIj1+sijwWsK7Byet6g36732lJahfURnGDvKiP1JBBGl
0YDDEYlstMXmjw47aACAGbavCh9f5mdTeW0hMcj60EtpJsSxF43ClY4BfnVJQb6O6KB9W61v7tVj
VQCz8xyn52kWhtSWx4hTa9Sb7vhzrUBs8PPpxQlzHKFeoN3zTap1sOMs0ZqilU38DssyPETM9yku
01MOPO133dsFusn7h+aYpbqQa3k2Jm6HoEfh/ypqxA/oFauuwYq4F12EZHLC/dMCc+E+m+mI6ffq
ePgdBLqye/XnwSFiOA1BYKpOcOOEJJXWgk0mf+dXuTBr6/rmOQZQMV9siJDTUbEZs103FgkZaPSw
gv6qt/GCo0cdZZBcW8d+ihzCg7WSsXrmsscbslcazFltlD1XCQ5QbQ/PeF051JaqXUsbByOTNAbX
nOqbYrwOt2ZaKboCmLpDYlyk0bM7sKi2OKYZeHpzNV03QyTl7Q6ec2bQ1qd1bw1Xter7qfkPnCzN
j8kFhXWG+sDE74dDUsEhUgINUSZQwNAcc+t0/GRE+x08Xo9zspy+C5V6n0S8U6F1rxm4pYvzecFz
W1AM9MdNNLH3fm03mZP1RId3mgIRugv9aWeByduWVyZ6yv9fbXfsHG/fd0K8xNsIH841xVmPqZjK
48hSY8X2Ru54q1uIEz5jw4GQVJ7d+nt9e8OcN3UgzwGcYI7cEQvlUt/Nv1AKPPZNMsC3MFfDQLoY
7hJUNOHyk+aZ3VOZhzs0ukS7zBHwUcad6jnaZW3NuBbwk0nJqYA3hfMEKDrfGwnz/kb6Ewf2siBM
jK+qShJmyaPNBE/Fvi46TLYpkoS2T5blHGZIwTMa25ZsgUgL81P1AX9humgjMBm6Aqlhz+8CGrcS
qaMg3kD9SnQC5+p6BKb0MzjS4BVoMdExiiYWQBtMmiScr3JKNahnb7G93a8GKy8cRO1T8lgBaTKP
HAnTGzWQBglTcBP2Z/eQCDuBG/FlR9vaozmESzBh2eaQehuMXzuW6RM3IRgH53Vs9ynKUTTWMEty
1N/xcylXoefTRvha2q8d7TqnRYEEvXzxCylUbwwf9cmYkuGrluav462unfNyXFhIZaosWfWXQigk
DpO1wkFjpD9Jrzh7BMRpnABxQg1yGZ/bTAy7ksr0+iMtWaKDv9K1Qq7NbwbQYN/065RuazE6SxQD
RvY8bTKtTKdXyUw+QjBSI7KJAqnc0zDqasJ2itzJg90Ixk6YwNTfepV+LR0PQD38Q5Iqut3lGL6g
afR+Oskebd3xOcukuJ6GgwElkIE/3udPaUDlN74mwHXchsWefI4heEeouTJoKaGgqQh42hPRU/KH
anzHpMneTSPsH6NK2fmt0shZcZD3KAi7g25IaqYaUDOuPysIaQEWUXqJjuJmsKqKkAMhd8Uetd5h
+jdSGWqHMs0w2RNtxJOPHt7V1iksgk0S2iTobXHZFBxyyiuWypvlpVQPfD7tXmXZde+Oa/CTaHWz
HLVcn5LiqFnnEVFFrdUh+G0vzB1nyxSOVoWeHPx/AV12ASyZucKzWeoz+HSjCTxawgQSn6pgW1PY
izcpkQWGNFa/7GO9Wl4xtpsGlsA5/1qvwE27PzlFWmoaBNNw8M02RPsLeKu2dXTRN44+mF0HLn7R
tSmqotLDhPujKQIdQ3J6rsX9zN8nUcGeTVlS4sDi9pc+CdzgfVs1TkYZURBJLeJAFx+sjkS4AWtN
AGTvGYK1w8m/+lt/8fFgvvB+AeNuLmajyd4VtjDwdU0whd3sQJl99FlgiLJB5bLok3QTBaXR7ESd
YAsFzXnTOaT3mCDtecSzisrEgxHrRCLM6P+Pq4yJkoV5Han7ks7Lr3B+Flr/JbOh97TP27JPINw1
P66I1+C948v5HBEoXkp8+p0jT6nb1MjSO8SJaHAELLKGjAKStrDnJNKzqdOo8cqC3o/fy8h8WNYy
bPvI9aSi16W+uFPZkU7G+0YQhMSyQYThuMuTxtBmoE5CfqiGtrLSEO+S/rBt/vEQ9DdVNv3PISxb
xwkqxplBWbm0h+KyGO1S6XQaBLzDeXw5fp2zTPm4RRmWB1EvWzMPB1EsCzI/4DyZw0ekns6lW0h7
/h8kgkfgsuC1+tJ/PzdJ2e5LteBra64daLi81NyJcbfybpiFfJAFJwne56mqlw0K27FItrmfuwKe
LKsh3TNWpaPMVDAjDvUTfcN8zS1f/9VwpkioT3hH01EHwIORY/Xb/jLFPFwWtn1iHxBrqfbBkc2r
2q9L/ED6Qex2uqmeo8jXtagcSU8pW2Q64utYCRMN5h6bCVb3V1rYTU1+VExdTvM/jlatidBTTTX6
w1bTnooJPm4e1nNNtIsfBVu/x4I+K1cxo72D4KCWwslZtKG++CkTKMu1GPXtB6fO54jc92ff+TLn
w5GVAniNzMyjy7BmAlYyRhNwCrpu7onPT7zCpS4eiPwxP/yotwDNIs297PclwuNddvmTtuWG4HKi
z1rHn+C+oyri811+2VbeZRlJ4PHxd/d9YHhSlcbFdcXObzsW89/FpwW/6+XbgDwzRyVSUDLj5RiM
m2N0Xthaej45z+tuHBEm+xS0zIqnpGFCaD+A86MyanSfHA+J7GUjYPl2jBekBmvER2wVMPIA69lh
nFs5irXCokl8fZT0WSg/a4AJCuWAy+qAcb44j0FcBaegOublxF3VZdgxTvcPaMvsJPydAIUrlESp
3I8YOxSK6Xn3VtbVQX7NXx6m7aFWahvDd5aV2Vo6pZ9xDM+36Sy4DjEwYrghouErGcQ2oXAd12Qx
vtv+1LuJZAU5qxtlGZK1WdI/hbaxxRWx3euYgqxl2jnQFlyd4V7djVf2L/E2bLSPmA3qMxXuaSR7
6nRMXneVxs6YNv2fODGsDKc4keXC4Q9pGB1Xng/nR29CpQJBt/xhXKvrzg5vE0uCuhH+xhYYfdMo
kkAznIj18Vb7QI0toVOA8PmGaXF6YMM9pSQv7xqE58nwbMHzo+m9sFjrY5RVO0rnsrqQ0y14LlAs
23qujI4T89sr8KhSM9PyGFyvawsUHcyUWnMynp0c4Lu3HLk+PSPoKJNMxfJc1DabZzR7o/8Re+do
drMjNpVqFFrtmlaSMEQbFC3dKkj2GSyUEKjhUvGvoDpaoLqybeQdEJzPP1F672v4vMwvs7E7gG5z
/TCm6iPIRmApa8XX3V5h7tRJZCSGNvq8GA6Rz74jCfuj1dFr4joa6NI52BqJg0/38n8lTwHIImAb
Ng3nmEIS9QkzMG0jGHlrgexW11tG57j1VUAWpZo3X2FyL1rZy4GPTA2fKtxd74t71/gdqn7PwAy0
HEv9D+sdo/klRjBpI+XeB5ttgRgfWktzfGEGlbX+PVeHxjSw74dJxmdZRJjXx4rWa3WLQlw51H5U
DuLjg9OQUgogI6Q/hMeYPG5BnSKEfWZAXzNrQmXKabssqqaHj5HP0cfz7dUe9Ca59Fgfsyj7pR0V
AXrPZuh2b8YaMEFSRsC3QSaVZCMI3UpHbYmC3TLg0hbYbJbFANmtBvrLnbOi0lJGaRToy2ILeqJd
Yq+Qru0tdkESgCPO7huVZlJ/GTEs2yuLvMBKXAg68qRTXJ46WNRzuFAuY7XyCdLQIoLGZcElnb6W
c5hByjxRmLERB1lVCqYYR+DIaFmcYiTMuArgMTYkd9+ageIiLqZsSoneiNPJWzfXZe9uVBAfk1Kv
Z8nbDk7UPyX2scsMdEjjsZFJ0kNBSmg0U2ceiernfhjOAMwe72Ukj12g2PHkloFWmNOOhEX+7dE7
HKe4eEz3lKI1mmO8CIDQjtau6aThv3yYh0Fcy89yzP8Wg3IfRmjmex8PQVylF6PYBGOi0CvsG/FD
NHNgEo38DEtiDDWPNELbbnVGzPFqiCJ7M71qdiLt10IAnCb5jjwhbnHCelzmGezs7axn56I6aCn4
1NszVGTnF3Wl1lGfADfdOK0pqH2MCSar7I8BETZIdHYtkKxYGEGkGcqtRT3RynfuYEPQ+oAn8+eN
8tRPE09VpvTraTSpdnaEIP5GIjTGYk1z+Q4D1HuOdsNq43Gq09NnJi7NQfjmdYPjqVk3vSQXhlZI
fc1pJMCNuUKEDvEbGqxIQi05/1X4bPBm30q56m59jmWZpKCDHpWf1Hg8zjMUPUpR11JSjgxe3CBW
m3FLa9fLtqJdkF3UdKNF1qeFXp91u6cOZg/0nV2qtaBnR4lCp3tx4M9WlUgUETrhR1B8yVPCYXJb
Los5rH5TIRkjgo4ARKFPK+q8iqAIo6dggKPm9JwDJWMfR/RXKSKrdaoP7icaoqodEdcUl2YL9ylX
Tn3ECtginXKZFU8UuqZspyBAb1/xwd0nMT2lQwk+JqLw0BTzjUPsNHOJl3VBifDuHYVIS8d0MZm1
0IUEjhmJsvNXsMGgWRbW0wJUnU+P6pQQd+lJQRz8Oh50NyiLESQVNAQIMRAoC0H139qeeaAJNILa
9qgnczIfCpkanmqtugCCoOnJzqkjXYWdrDoL0bwbO6nIZUBXLx7xVcl5XHFZDmJ1ku3yLZgDMC4O
nxgcgQ8yLwNSbMv8BF9uKgYhriVgnjGJBPHu/GQz+aGHXgowCCPOnfX1rSC8Z/x1GLLy1OmyansH
mKpuLaBbItvQPJvfvmwXdXi5VDwgae+ApS0CnTFDokNJNp5+e+WjALZRAw7RF+g+GAKcVjrg4u9i
SZYtsQka7rUyuuAb6UA1zj1HtzgqnmfetxvespxtlO+Cp2tLVZkkv9XFjUEKpki9VX5BHp2W4tXi
RJGE75e/kqPA0swi+K7teR2LsA/NFSV27CUDKpHn+dWhBFjebIQM9o/Shy0lvopqhh7ky8ZTaQrz
PbXoQuHh/K2GnAr2aLbX+w17mgc8atVls7k7A7AcTCSuO8dtPgoCIRSuEh2zYDsfOkTM8h98nmFO
3Zwb85DESkRUm1uIKU/9ROEXViJP5Re9d1BjMglVfRNLvrgCCGfLNHe6XIVRVpsRfKaQ9dSJUT0P
mTs/MHZbSou0jvSYmbWOzZ5G74VzchQa5uW3eTupBmfDMoh4aEI6J+V980LCwWJs0ok7Ph2Fyk/g
glDvpLMk1TCekdWlrl5EI8ygh1VcpoDyWB37sVPGA6L9yhwi7DCyLMgV/T3yTyl1LYWdUczImxkR
+j/pxOhUmEts/2vBIfuHpi52o4VKl+kuSAtofPA0LOrW9eBDiXYSyJeJ9mtKnZTLP+hU4IJ5kvxm
OXI6kjPd5+d4IqCQx9x1NsxplxLikDB0EjW9sN6I99d61+UKgVezRS/XO6X1ARXR2brnoXKYpP27
u6rro19C0SPk3LKlXPfuMGthUtrye92N8RdmjGupClRwsevN+NYovdBYz5sAmo6qGLwuVuln+62i
TAeTk6I7VRRQrVXOdZFQeh1REm/1TmjDlH+C66OZL+4JMqaTvWP3FR27YmFkP9H8fDAWHSSW1hzg
Q1kx/D7oIr6EeExRsU0bEu1/0UsbwZkjPeGF/Bu4qM2kV60xHZ+dVwQ/J0SSK1ySU1gOkxE3Pfck
lzUrFZUXTLdg/YEs42Lq2JWB3keexaBWLQdXhtxLOcJAUudZ9hYyGe1IIju6tHgzpwXEBgDww5Dt
K9P/hU6LYZ4npUYDktbho55Tm/t+PRaM96tv50qMultT6iCeOIHbfVFSFVo4ZTX6ziOtnEAUEf4J
Yhf0JW9YpvLWZJ7qJN75aGhTKSa8sAGpbqwW/axxNw+aQFBT0qHau74g3r8waPcR/yHU8mLmUZ/I
iVqbzNjYbM9b2XLsHLoMcc5pEp7V/EYDCkoimnS9LjCQm+pE7QKC9PSbupSaUuUUfiPTWH4qfm0S
P/AovAaITapcbYMTKKuHpIIT9z9pll0FPsqW3bBuE1bVjw8PNfxOx56wfO3K3CWOEwLd3OLQ43dU
U0Gx9SqS1QMDhfZM3Ys+E1vYX2LiHcsJoEFp0FFuBp183KzfodnL4nQybqjPb91srWK90KvacEhq
ca1gkQRtDF8yua37HUB+rmtLt1oHly6eICtXjIPCEF7/2x6Z7bErrJkkybcwFjo2X257D2lv7Kjl
UYTS3mKxkQ/4CmuTUebMpbH/Pra/jJn5DCGwkwbkDL1M670KIKn+yk6H7c6unljLuheBLYWnIQce
CPzNotJTea8ZjLvDkwNsgvUQwfCQcjAkmUzIpENsLT1349C4m+fRrPqlF+cx+zNlbZ/32mbv6RaW
Ipib1LOR5oWtrVA4FQ8mSr62cC4+5ZOtjLP/UGdE2pr0N7iH7+8T1KBugkFMJDPudb1q0sFd+upV
I1dkFiUNCYdHrCEVDKrncKyN7uKUzb3mD7qWXMn2QEXpvkokFnGsOItJD3JMwOgTkBaDnPUX4omr
ebuxL/HRV+gIJsquVAzHWP61IK80OtnerrBT/ZrLP3CvEhruMUlZIfPYw8EQEHY6A8MDwV6DdSE5
67WbHU0kvBnATr6qlNJ6G0//qGfA6giIeTMRT0ILBz7NL0pusR7IP0/DedpfRbBV1bmOuMJvsD8w
lOP+u5/SnNXIdrsGV6EJd5NiC8wOSuODqCAoQgu9lyVQG+C7yNtCGA0s0G9Ema0OaaDaE4exTUUk
FrK66RTt5z0rvgLqJJ2KMJ9o9IZms3a8RCqA4Ug7lmG7egJwF12L4XjADn7soL6J34lqleGxai6u
jaqZ2P2NvklVd27K5NHPjlRyBneZvK7AW7rUHtN80452mVbF9gwf+VwVzVH/4u/5zitL+L/O1waj
4M+PuZ0SSpGJpbGijSloyLwNDyEQT/TLJwGFqqSxn18aF2EHJeG3ofj96y8VJcIL/38QRdRurrct
ZjDN6OMyjWchyPx3sUsGEezZlL+3rnks1x7t2tCDjPqZfHMsqggtQuWjS3tYDEocPPdQ8z5cOa29
KKmDlBScIZJk6xVvFk11ZqkKxi2YqkToS/Q3licWTJ9zD+Gx1qhobwWDji3Y4L3jXt0n28V776sz
bsGwyGTA6nT/qvq6ktJpkmZvPFTRPR/LMrVVDvkEFpuOjLiNfH7CuNEyF8RgBHIWDKqG0Mu4fDPi
ZiQ8EOOIVfxm0Y0VwTWrz54uWwutqa4AePo9Wcc2PpTnVBzGcM0MFgSFdhw7k85vdsJeu20kBi/g
R9SqEW458C709B8wL4m/mofN3gSoJO9slGDgfRKruiaUOIHfPo+1Mh1n3iiMe1WQH+vEuq97yyqd
pmOPKEm+He8EFyqmIZ0hZK46Ngg7q0KpkYvwqrC04d2TXsCC4nM4WM8ymrysbnL7O+57TM2P3mX1
at6ZjuDgl0hQjAoQGDsOkDZKEPCUxogmgVuPXvdmPiKJS680jz4a2VRjaNjjV9ObyruaKwOqG9Yc
v+UwaMATc/3+P5xXtrkuK2TWzL1lQg36Cxov1PzQ0dFjgL+/6ulxVG2+psTtUKx4RgXnSRoKMctq
+IQEB9PuRhuDa91gnh0QYyQHlvX3eoeNzn8qxWn1GAT++docSrxK1mKN3ESOsuJNpmQXFWxRtgnA
OACJwvlKTLvIzOm3R1GPt0kMzTWrSm0d7wi2nuTtqrKD6KLJ99bzQjl6x4WSqvGQ4Gvbw4JQdmne
mbuRoV9eoPU2LZWtsGzmirqoba1a65BtM4hx7tyF0SWkroi8QStCpJHxGT65joCkx4d2ELvGBkod
/PE69DgTn5Selu/Z09F+elb3766OMtnHMs2bBTZHVsaur0f8y4sVuH3Yk5jkUBx9z+hmkru830qs
+VCscQ6q2LyJg7mYFcM385Qii7BRi9b9XMCyhZX9hc0citTmpaRPKm/q35we32pxZZ9hPNaRA0WL
e1AysXw3eLn5Z3Vk/rqGJCC3cyOJM7yENsiQKyrr4cjqlFiczvMePOIq9kCnLakB2UXYGqUXYEvh
NRC4wqBp3TyJbLArQgFcjLHOa9bDJN1S1Dc9oaKhBycZrlZT3gM3EbQ8CuQ4LD5fRyNVTc9bIO8W
UmgmWzEy1JMwu4dAd1oPjwhm6ZLeYHR7wXjpO5JODQDpGf8VT4HmwUDgzpBgM/b+wcW0mboLRp1j
CHSpveCt775RSc/CQhGvbs/pwOHtZ+zTN1EOEbnzE6qRZIUQmW8vGlh6xx2n83wPGudjo8MrUOd+
H3xy6ovBM/JtLy4w17WYEXoDkz29Tn5Co/9Jn0qpjUw9hlIMKvd1fCNIowExRw9VKp60EQ6zxwOu
r8W4vv/HmaejqWuK71tfo1lV30/UWKQ0PmbrUiOR3mWOs1pIG5Un17W5oMZeuql5sImZbv5bdbiM
bKQmuClf5mfiTAoj1tbBK1MpfL0EhnvGXzPs7aJqiFx80rD8iRoET4SwoT7Un3Fxkp3A84D9fV+T
5UQDlEA30ulnSvK/kNcPSdbjob2adLxIVyHP5pTxZ9wFxq9F1mLyYxDtB2mJh2mT2hfOXpij0C1m
CIf2e3XJOnfEe9hZ+cIHum0hw0/cOfpioKwabWk6Ug+bMAUUeO+cB9Klr/fgLwWUjGW7UI6AMqm1
obYyJZXelMx95w2JQ5QfZNP4irYHGvYdfCaQIiUQtYwB+gx9ZM3PI5BLMKab2hP7l8Xn1yr8z4pr
x/p1Dbffk86P2Od6HAT6HWjO6bsDzA84mivOVpvR8xSL/vUBowmUBWiTqxhm9FihW0e2UVAhpm2w
zwWiiiowyjAFbdQjUVGzYqHnQktDtKLk5ZwAXIoCVUif77HBpssUPTIurg9ont2y5BnACGu3u1Qe
JSAokVjg8/kwgQfJvaijkWhms0zSWJ2q8jEUOhFJIYpM+4dlO/YNx57rZ5e3oldkCtOwEUX4GswJ
e6iYyIguBjBBVyxzIOnAUigOygvFCD1e1YGQPAATSH1dsK0/iY9MqU2FtT73uRxsHQhrN8UYAxOo
ZMm1Mj0OEagZGorbY5JLzoLHF3sOEqnJ8yECZg/CkPUpjszfEjDZHCG8rUxicTNoJ3rrpNzIynaH
kRuKOQYs2gzT/seoCtvf0f+nP2d2J4UYjTC66EglH7tpzZ1t25BGbFPdgBF1mDEyADBZhBPHHEUl
XMdlos67ARoRczK6vPk8mq/DugIFi9eBbS9pYtPYNIjON83LhsT/gy0M+chHiLX3ySxuRlNIan5f
4lUktrPwJvBEi/Hjd8q/jx05rqol2SKAi7K2RF/ppAC72ed7Zm+STFEc77RWAnRQOn0XqZe4j/Qc
rc6Eq1E4nhgFmotCoEK6g6tszq8pTKfgRFNTuDEFbJbqBJagSLS/OYC4X06Z3I6a6X/k/Bm/1Nnq
2KiKLLpqgpUCGf2R4iqrlljghbG7++3OzuBGlp/z7WLNPMsHQ1hRdW7VNzsh3FB1FCxi8Budkjr1
dC0KdD8j2aBK502ZZyZ/efT4HHE8Yt/BGdIDj5ZIsiQpNGrI6ssU+mbaSx66fE9q3dJ6ymsguMxE
4Ia4zaZ4xTfO3Df4DfZAWmjlL2rWjq1BuO8fitGFIiJeVwwfv01nvqxiyLCem64uWJfWK1PhMDDE
C09bzE4dnD7vsx0jacR3q3Q0E7o3huTr9ILmw3+yq0QxASibQCwH1X711Qd4+s1r91ijC+420nS7
9u1wROdxSOqVE/4MjRPj0exTssA/uUlnETSOQwX2wah+TVgQ16wF8qWMpKkFIMt77athV5Lgw8A3
Zdw40KehBaEtkM9n/DXwU8D1oHqt9uRKJeTIaVB0oHxcjbUVZYUl/h+tCzLwCQzL6CCVaoIHKw1T
5uun+NR90cIPxNk9WEG7+tWbix9LSn/7ZfR64OHdrxiYSoPAeQeWpsVeF91yn9melT5ekmSs3gwf
FiyVSKDoWOjpEAfUnhpXWrcPBltUs4DcypLyR/UMqSBOaPCpaLo2QlOQUREQt8xnrhR/TpksMuJU
8lCY2r1Prw3hrlBplVZ8/UfrU7ouZ3Ids6yGAUDkfAGsXESyW0ORG2xvHczv+P2rG9TEWpWxozOP
W+ngUrO/RSyurhfqce7Ua7ISd915RlZ3lBq4MvPBwBdHErALud+IOaEVz3p65WK2WbdEc7F7lVTs
4Z4g6uaFPk/sV0XLXT0YHiCuuA20cgF/K3NGLkTov5y+FmSwwBnG/Hi2BDlOaziAZ1w+rnyttIh8
A/2Zq44KAco5ysVrTay81h5CiS30ioor+HRuqD4k6udU4pDQrcbxJRUZgK5vYGw/McIyLV2ok6Ge
CT6kqlsVs2DvhvJxiKizNPHbfdZrAS3rr0T1kGV2JqQCdtBRRXiVrzydgsQF2omevWNPBF0wr138
UGGy1F8NEzllrVgAWKRFpKBGtEweogcGwHDZq9OGqcPaD2F709D8mw/NZeHiQyI5wcT5EgoBtSUx
QgcNWnVOFg/3hKfc5kH4vG+p/3/9Y4oKedpTXnD2ZiUHSA5zhe6vqGIYtmsrnR58J8/lYH7YAwxT
0B5NdKJtS8MhjApZUnKNO4iaWwYSxR2UvrWv7mnjdWj4RkZaQaQC5KbR5cs6pBTa7s/jqL0bUX6d
W91uGzzkecd6H0sXVBxb6J/V4ztO/bNGzZO3A2otsQC/zNnuKGM1qZkXDp7I90tnLYzXJpkZYYEA
5S3tOO1LJnJKqlC5d7k+6g3/yxTdrVcy5eyYn5oTHkhbjI0emXAZeEOxVlieH/1Ji21RwyFi/65k
6UdCloch7wNup69A/loWJreUW9PDvH+zbDUQ/pL/f4kd9WotBcOF2SnESX92mfV/W0qMRnZbNPYk
8NyPgmO9Q1wggaNdb9OFg6wwxm7pSMxOUKoBdNR6ysL/R4qOhoUeWTtmaecOGJatxl10y8IFpqh9
lnwniOTMfyhvQ+DJWCTDeyPvVfonuNN9GRWeUoHlnpVE5gm8raHhLxbIPRi0FCZ8FvXld8dGp72g
We7drWOT2yGlQ3ER7pssKDel+9GaDtmwjgjT83umRuf3Cm83FGKC/gQFg1gI3wpqOFJnmh7jj8Qj
35YLJhbRh8w9cIKzkV+opWsOZ+JR4yJGlCH9wWY92k6ilSZurZlVPiyfR893l4IwQfvIPU5lhi3P
IZjPTSAY50+blSuxgDY8Dg22tw71E7O+UDkt+gdMk7r2CJyLuK9bVE9pg+Otcgych/G3VpnbojFW
0oQxq5v61WZNzYmF8YHjp/FaquDmwwl8W/wqeX9yz8KxYbADPk/fd8B8fbs4Tyak+nCJkbVuyZJ7
fEqQxEDuq9KBtUsn2rV/qysp3gdVcgtBvm7Ur/5p/wre1nAr1mAS0h+niiJmCTrmJwHgbBEqMgQd
uh0z98oLOOPs5CYqSwq7G4xIV3UwQiZiYk54yLMGAYQdBBVrYk0U+YEZw7nbeQwlnT55RHpdhDeM
+i4oYoH51yftxDK4+LGZ3rqzNwdmRE4DieM/qptpK6uGjQyfGL/OMOcdZcGy4W7afLthblRN6aIQ
LQWhK/SK9+bveNDtGNrWHeuqPZnzB0bc+f+KaTutyhy05NufH2fIX9VjxkL1kcqLLbyWR0wVzmsg
lnACIRPejpKemPraZIOdjZ2YvaIdp5dnaI3937nVZ5Q/vURhWWhCXouPHXNbX7qS6prowZNLOv46
jVF5Gv7aLNEOrUTC7juxV7DOsn09HqN2qKHTMM7P8eEJoKw+JhPB2lRSTleK5wc+MSzeRiu7y3Qq
fUdNxdBa9NJd7DPT1MWMCovb6XU/y8oBClIPkpw3gz610N1DbzEXTvq99Hupk5pObqBQFTFBlVTo
n2mdtvfoNTwbfg4pYg7gobh5F781XJ3BjtPqjuI7PoIt05XhLNbY2NEVIy9VOtzGRtBB2+Fhscfn
80F4mRjPytBCeYOxVcnWn9+olkWJXP+su33eXe6r0wsCvhmyAL6X/DqRW3DiMfifqH5sXsaBZ+17
y7P8lIVdJ6SA9kRZO1yOSiQ3eGTFTzSzO0J3H0C4CSjKOO41UXAANiOxFaAk1P09KpudxQJairpm
Xk2Zx378b5kt4OK8zPt+yGinJ0l/jSCBYw36v8BoVqjpTCzx/k3CXz6YYv9FXwtuXcjRsZE1ASrD
t2Wk6ieSZ6ARRh88b5zuefEmaTzVq8y5ZiEVyV8/MnbugzeWyWgN3aEJpp3MrfYGnqPKSQd9dBF7
cVb3It35D0a6OvTOig1X44rHpHot2jxO2yQ+09xqpzHEIvQxfoFTYbzP8MPzM1xqft/kB9mwgBS1
mKFnlBKxcclRenHOjEsezTJvzt/SFg5/BpCQjs2n0u7qPzWbnOr5l25JGzFJxNQwkZJRgESjwn3m
dHr/pyHXQD3fUJFyCB0SjyWaw5SjAHm/JiEIzMMRbYvlmxktmLFSSL6P/Pbri9r7kX6WR4PUUmV2
VsyxWb38Uh4uqFlAN68emSjzu8/rFzrk2ZcK5nnAasQA2T0ZEsHSH9F59epW9dgUPHGeIiWTTvub
xhz/Eefl6rZnUxd34//tyHzxkEK+mP5lyfIOEw/1W0o+r2FlyVrA9bXaK00/XtM4uZlBRChANX9G
eEYmdpy5AAsX0fKrGVv+32ExPW0cQTX24Nq4pG1eGuPivH7VzFZbC1c+vLsIn6w2VfX30PI6QI07
4w3TZfhbRhoAjMcvq/Ephix9hj730lXRSo/NhCtH3B3+syBgyEPgoF//SeHTG7DblzlltE5lHGwO
xy4Zc3rV7JGtHTdqMx1fcAN3oD6Q7CpiDQRdRZL0kgJazYUXjkmSL9yvm0uY+HSetwlS4g6BnRO4
yVWIDjOIoLca8DroLkhz7ll4EH0CVFkzI46+y/hJ5+1e4Vnr38io+gLWe0Gatu/ykkCJusBJPtu2
a/fpEURXpvFqlH+5GlKfd2TiiC1yVOzwNnV8Lk1NtFgR9YV/TVscosrlmwxdSV1pHW4liJH6LjGQ
sn6w/APHchizhInIewO6n8So5B961AOEyL6OZDbsUHhtaDAUM92cIUFEFbvdveK5vGyt0mAV3heb
PR58fJd/xz0S40GDYdZD4+SEO/3Y/AdZmLleQzeEiHEOvbENFfwtsBBtZSaTMPAiUd/q0RhOyhqn
8vrfQxPRs2Cdv1vmKBgUpDjo2/97wpv6/kdAxOQnhIHurVO/gdBGeeKiGhFF20mp35ZKhsg/1jNr
Lkaz1PjxQH6fZqIKfCWoG25AEYvRawezJGHAq544EVQChb5rfcKvFd7qF5mUs2F6iGDG7e9rrc4I
dA98Dbn9mm6QTfwwVF3aNCyq7iPwG52GtL7sk3eFb3GnLcTV0OCml+m47PwqsqDUJ9DXI0C+yCc6
1HFxWEcEAXHJY14wKLMzrpMyXuBu3BGJUw0Zzcdfax4sxLBZB3xaOSTuiTcszto8HSGJqbwC2v1n
TGkn091qTroiGX+VnNyjQDEbTTlUbhwLGyA/O29RHjBRB3sA3tepZuDGO7SreLIpt8t/MOpnSOZT
H01/AY+1WFpfT4Jjz2N8u559Q8jcmTGbuotaksz37jUATY5B5dhLyYIUHWZS4av4mKGV/90LzGHd
GV7K4bP3JhR67JDqEgyvaEXGglqQCHVxUZsJMhh0vmYPJTTDPg3tqdw8wojq2g14OJ//6AWeVKvq
+0mfW0VPapdZXMmnNJCLuH5TzJtIAj9SmgwrUduqkX6HSnR9yWZfh2se+l24pm7pAXWO506zB+XH
9P6sJEUAEPItYSrGp202qR2CdATk1sy4M83C/IpQgdIzH5CkyRh3Q/lsr8uAQNJruFqDZEj5dsSQ
wTQ19hmdAodokmrueRH6BGOaCbMqW5oZtGOYG/eOgYk/lFYEVaxk3jRpIKEQYi7D7xNulCSq3cCH
J1iqGF2bir+oJzOD9EHG2OrSfiAiHCniEJXslF40PZV8GdOgzkuiFX2dTg6PUzIKnYHgGE+hyUfw
5M8yJAdEUKSJUkl/9PNp46IZ8erKGl8ce0nSrOfnsrsRXmu3GO1TQvga4L083eb2b1rRxPA1oa8T
EQWosJGXx0FhfYtLv/SaF219iUYLEJjWd+0xtGhNYugGPQ/VtP03pdpO55F4KgV3broI6kFEFDNk
1rwKSfYjhfSGDjIzw+V468GSgP+MvoLvExXyPEjTls2Pl7x24b+S59YFzsHthYwPAgUbwFJwjwQE
mwv0g/P3fcUU6nVTPaemx7WmJLX8PsEHLTHgUlktLTORh5KoiWANp48NbB4rUgwZ8gisCuuwuCWi
v8+p+UlmAdMmsNvKqQJm5hrrKv4GwmEv7p2zz7bTAeqMgc9N5AmzFQd/xoW/QjfcgOr/64xW4AS6
TZEpLaMTVHPFgC4Eyu1jS4CNqvthDRr70K8mVK+D1Yt+QnkeJmnb5xqm4umi+xIAzz1NeE2ivw1F
3zR1EAo6rUB9/qelM1q+ZCtoIc9Z8xQoOQc9Q3b/DSAPXi0w6q+ehIwZJZJ8qHnrgfcdq7Jl8Vgy
A7/Ki4f7co9NXv7N5uPL2wAsVcbFcgbENQB0qiOMp6D9OovnaaQvDvIbVfC3Ffo/gx/IEWL6p6Qn
dllf9YMz1JitQsrqMycEWUBijWvSTLd2pAGsl/K1EiVpQN4cxYgmOXy+pLNHauFwuJd1PPn/AsLD
nnReyUhgZOeneobU/+tsOgAQiWzBhm/lh0BhlHiLX3nYsdsXkcXCFmnUnZXLOqmjxzf+Yo8RfbgO
s4c/jlv2awuUPuT8kGCAAz9k8ySRGYNefUarmNt7Pf/Pm6Vz94IW0JM4I940SLWw///6XWqya90p
TSEYWPWRWV+H2QPOTVRzjS9H/bBKgyHZ5B5YiSfYgiEP6aCyaAonkZh6CR+9+ZNK8WARiLs2Exht
nPL2+dkIX0aOs1JeD4GJ5xyNEkSN8rRl7yGCJeOV76CJkFQ6UrERUftrVaEZYwRXwWUy05zZRCwz
xDyrSe4A6s3hKvdD3klXMCbAvFc5wDHDn7O41lJNr1CygsrXkqVKJ6Diei4II+jaiPeNk77ZxQ3w
eMd2bFhCVelsHGt1MQwBfONv3fxD9Iro0y8xlOlRxUe0ySi5qjQONJm7N8/SgTOL/4sCiH20poY1
lQR6+mzKRaW3vDNHi/ljz7577DIjfpwS03QnIkkU7zcgkGHILyZy4AG7F/2A80K2kCG/uhOAiBo2
TLmF+K9yzI52dPzpNwjf5O8VKHpgJfyX304OOYSWzNaOwcfxZ1a6V/nWYKaEuWMpuz0sU4EycgHa
W57XPHlR8ovyKKPMC9TPyOhXk+mly9FhDb273q72fS2rC1YkQuh4A6CcLBwrLFBCQKIfIN8mtHia
3UM52yCmcxjP58TYvTT0ZUaXnZ/8yWwzLsodY1ZbkfIUGrl3Qi4vwCXfIQavFyq16PYFJuINgK2i
HqzvNiGE7NJcmgKy3eMe7wlaLsi9cEON8fEVVFsy8u2X5/60c/FpJtOtEqWcfU/Fd+uyqrYWuEXR
mnSeazWEKQqWir8Ul3PYt0IqP46uPL287ImNKtsLBVhTJ7In2JRObAHFjfCFPycgw13OdjpFUfhr
lLEr2m2F2cXcFWa9Lo991E25rWFM48qWCHMNT++m41cPHi7nS+UcbWhApwKpIjgffApncnMGtKw6
SstZVZTAnap9zmjmyPFCfZJ83Hr8W40GeWSSJfS8TIyqlPb363mEctqGBTibM/GiSWr+SKnsN8Cr
XGzvONtnTWG2opOx+j2DZ8marTDHSQe/eufYlt7XCfksBqi9NmiXRGxedGV5hLr600GL3EV+hbWv
fvOQe3Rlz5rxhMBQReNm5sYutP7jhdz10mLOT4uL7pEiiGyUKEwizl7NW6Rt6+KqGfl8QjuPlJtg
nANux/Te0pOVfocTQR8WumY4lalA5PtSY80L/qELXQMZNZ2S91DD9zmdx9U0LKuvIrEaBRPNTMTm
SlnBqjdyU20kwF1Fsxp4tSpVrRGJPmHSck5k1rndHBfVjE4/0rrTBFa1wfL6gk1AATykTXfv0H9C
unPY+r6WQZCVCjcB7MhmKJUZIoGt4Si8UP9/QTiieNlNB1SUfAVrzSNjfHIBYESyKoKutyrzDq4T
qP+lnrNxR/QEjfQ+8VbjAzrLJylVqCzIr+orhfnxhUA+xUiQZ2HJZIG+196GvHXGGIt2o5dTYm95
Bualxp1aSJrtvNknFiG3UHtPDKZ07k7V0I3sBGwGGneRjNNKZ5JF/lhr4daO2zmn0phHBXZVXNGF
ML19OyKwgVE5h9wQYds4MqikzKBC/Fi16aCpPailb43a+tC7xbK68D2wV+mYAIDbecOyb8YLe8M1
wCjc9k7LpwsmHCdfcelWcVim4sLq7N6G6ycH5KunWxXaWhEStobSwhEN+Retvk6V+4QT8hnZi66y
UmzG/Fb+ZsUna3KUO6uLVTQNJPAntYg4aUArTANB/uwF4fSAF/LS16I+TollZ/zW6EEeE1/6bk3Y
D/6C8P9cmM1spXBSuW+F4gPUXiwxE9hPKqRXZ3qXwn86nctcNVyO2pKtoc17zesW5UYoEMVaulhB
noyVX+4ISMZXxVZXLFOdaO1ra1hAoK2ZDszXINipuVntpNMmBMVICn93LaKX6Ry7biUqJW2FpSpH
NJnS2iED57RdpwT7vwQvNhEwUD1sefNLlXzysWv3AwO0JCdV3RLYbe/cfQeaTUFdR/6/NrXpcOJO
dOxDh37QIm4gTDwgbrxqmOsf15vSxL/H5EVcLeWNBvVDHji/q9iU1jaeRZZ/PoWn7rlhvvHW1G57
K18L28HBxlq9lkvlTp1oeiztEx0bVBNnuSbqhlZ6I2X+VoEgXJloUybY3tkqYHAiGkio8HCTUVRl
ZfRTkQQiLhgzxi34eHWLxI/MpMMYkxkPw4mxq3W3xAsHeibpdvyCorPVcohF9mf7Xu+t0GAKQwLf
0azNeOO4nrsC4Iy1xn7ER3VxVdWIUUavF/eX+eslF+x7yjuyclhsTl2C350F/8j85CRozGG9KGKf
4ZcFSMmZKpYfmKn9ZdtxwuKMqL4xsqVqziE+xkk43ABPMAExdPYA3idHBpjbRgTtXqoqU1a7+jyp
tHWa+ah8mYKp9hl30hxQwpHwZMiQ1tMdZdbSBDu5OEA5UO4xPjFoF7hbV9jwTMyw7UCTXKYAwop9
EwnPiUZLOCFe16oxoQ/0sNRDEYlf50aMrqfMnLDqnfMLM6f/e7sntjtnsdOSnL6J+611uUN3EGTM
Lvlzz4zwrOLiJvWsbZhNRljjmKLPv/rNCjjz+lJkoiBhLkOeLrzWGyuoreEvuFJWo9xeST+CWVT9
TPy9BeYPsWuMUaLblQ6Z/FZRh264Z8kMcNYay4iq0gfLZNNV+MXTJ+3xGMEHxM1pTaKUOhtWeCBL
GafEH1ynLICYaQOFAKSyCESOBDb9vNwN4uU4khB0qfcW/3GMQXKAhFmqI+0jFMljyvxOrqLaOnTZ
IT7gnjknkz/0Q2b06eC+a9ksd2236gZUTjTTHDQgTXint9moO50YyJwZEswnBKYclR64Kedna9X6
K5V/3WgVM67fcizfeEpxP3jy7ng42MdboFFeUx1Aeu6ZOfx41MPtvg4D7071XDi9MSDNVSEaVVOK
xfN1yTVHJrtEJPW7l4PyPuO3+aaXgzLLaT0h9XX2Vp8+Y7Lxtcpb3eRAuuqtegpxOhX+Uh7ajYF3
hf2PUZcfXM8Zq35z0ZBR2cdAMXgQ1PfhF/KVoFbLIov8vlqZ4krrOowa1vuIcjSZU5U/6OWuljTe
tKFWKkTUQu5+uN8ToyBZjCc2XqX9QtLAfMDIhiV1uh0L75oEPVx48KaZHiFLs4bMmNl8RiYQMxHM
beqsWx1JlFbpmqOxynk4ii2/edMOUtqdLLctnw01vczzyX82QHvWrFc6GJ+GI6JjutQmp8FZhwta
AZSSR4vB0xIRmVeRc+GuTtIlXUBk550/XH/lmKQNmKp/QNz1otv8VOM0qCwyWQQf3hX0hDd1qzFB
uk+vogo1lXF/NhIZogPBQZhjTtMu07SBowtDQcti4Ho2WSZLELaVquQxTHE1xKl5h3RM9tKCEgnG
tmRigAeFFjGjB93Cbi8cF6DC/s+euldiG2WeprxDcgsYB9yIZKWXf3OaITarmgJ/TZXuGzY9Zhet
PTmmuRUMMZZP0F50VNvcKH/Ld6fX7dXIGBxeP5jNfSqjbSmFo0bw3vpFi6nHTq73RcIU35lVvRMB
t/+tHlXGzjOn+a1Ki3bTXTRyDkwmGSDC2p+acXUofX1+UmtKPTmoEWvqUddMcFJ7dlReOxzuzaTV
W97rwYUoAjo8VaPfzmXey9ULTnzuVdsqj49TkadoeHntLTqejwlO43D0NzNinTCzCcp4NmyGIDPS
SXDWCka6auo573dfA6VguqmHQxDJWOh+bOnvSbTCKyowx5WEgm9uJA/pIaT4GYeCjItUU6H409vd
YBeGjfNV8VCoKi5zZ5UiRmeG9IEQvPEi7LZAyIAlG/OxszKe+deSiqadm9yeqghJs+Fz3E68qpkC
B2Sx9pQxNFlyj2T1Q2gleGRGfDKLP4j6rvAeTAC37yrSk5fINUHrWtV3stvU1gKV7n1CSG49J+2g
YmCkW2UptrDeFbgg01E2NIBZTTjZStdnjuGU+zcpL5QLvfOT0+KW6r05t5/dTJvW0zqlfgiyqrkR
XHqFDf8xKalu9el1MsdThkuYNJAcR4QaUrNsQBUynseM5TfK9Uuke1Q4NbeZ6IlQ0akGw81ipBLP
vYOBLcJTIKZj6YoUybCdUFAxGNR2IrowIXjwqjeFPwS6IUOv2WJh+j5TNVrj7s/LrIGYaxTWlUZQ
CFyiHTx6i7bKW5KHAS3fXaL1qSXu3Dp4xUezqm6DGA3/4iK268Wfx4ztMyc64j3wtEydjnpoAQNz
B+Dh5WMFPncsy+Q9T4UxAcrIclYsgjMU3srBWmKFwdqwP/sBaVo+P3QPVJ7fJhg1buWGN8wQB8EO
d7wTKG6NX/hN0iFy+YiHX0j0PBM2UIv8mLh+1b5msvcYvfE8dIaImqTW9+RgTSeVHHvnkX0X7l9V
KJU7XvFP7dNi0T2QQ7IWHdqFnUTEqBjSRY2nGgTO6yY9GCiyVn/dhKO/YMX+oJa7bro9iD4LOhCV
c7HO/dZ+RlhIVHqzgdNrxK1evTOTOOi0MQnDqrAQTn4ZsuUkVKVS4cxTUeqXs4b4uRmCm55jbVjm
m78gNDOduDdc1Buu6jJpK5dB33rnV6jUwnyKB3F9bJGyknzerKSI3xrcva9Q3ZBep0RzKEpdHIsX
Dwg/4JPi6cOuGQgdZ74JJ8NvKhjkXe02389kqbPqeY1WYxW6lZS382htHrGfRg9j+qqVSsJf0AXi
6hwC8j5E5Cls3Avc73BME1YEWqtjLeetrfApHALYvCE8g1KteX3yMGit0Vn23xg1CPaC8OvRBnW2
cV58XDs8l5LjxrtAp0wyNWW/ci+YS/iij1G3P24eNvZI9edUC5JWhvBf+tfE3rGD75ClhGb7WybY
ckWepzT0tpgARgjXggepyOqq3SsRw3FYulqiyfQl6vGExesCmSe/uGC3AKw82OndR284/EmHn7zB
jSApF6BKuzSd6liTWWjcsYmdDZpvFY9iguxnum9irnjY9Uh5Zf1AztWZeehG54iTap1JYtD9fCGK
D1sofFu+L8D2K7V+InBRw637jHpOgak/irviHGf5QaqzCF8F1b+bn6XrABpZH9iApgn0UNWMhZzm
rCDTOW6Qa+nNtJxH0kgp8fg1l58hdGHk1qD1yvN1Teuw3RM39wNmpS0Mh96mzhUnNITk2hKPQkd5
QIAyeMuy08RKPwNe0ETP0+hO7BkcJA3C2FRS9cpmLO3dx2HVeLvQrT/LFgC7YwkfjBbKahyf6ytI
vfVg//wPAsypH8bpnbV/iF+kfhvQm1VLUqkqb63bO/8+3ttlG7+ohlzw0mEUriTTHnHcP/15Fimf
WLfguROMtXxs1fkFjyvJq9Ra2d9cNd9LjOc6/iztM3c+xqc273wYfrBkPcY+m8bzYzdnRSxuxaB7
qqXkzQP8eAQPEjPLK9e7xFPfRBOCx+8189t6qTSvUG+F4Nj1HVi7pjmqRyEtc1gW/2DjoJuxpRhi
+63jWK47RA5Rdup8Qzmo2dTFsWyVZhnxL4oRGVrpKNy0CIpZcpl6YhZgYLwa+pyc9Pb4NPeGXjWy
qt3dKitFxUBg1PPAz2/uQqEkLtXvJXMXRZTFZedY1eYhKpq1tOV3QggdvBUJs+wLv+/C15raWn9C
D8jJs8n2VidhdkNZWOVyMfvfAKSS+qW7iQii/yHXSPpz5oBMNluceo+eze47mla5qIk2gaAonotV
IycBdC+TiQxbHUrcR/ikYAzjQvdQjhOG7mubx/LBNrQKlzKseEyXSIQBi/8aWSb7gR0hZTsnjt5+
SJGk3nVNArQ+L/D+Hg8W7tNuMTcGRWREibV8D6q42UryjgSntr+dDYoFnvzVjnanQLFWZfYMbhQk
dCr5J/deXZWPVwOmG7eoif3v03tbZ5ZMRCHEjgXYa7PmWP0TA3cxey1F83SDq9no/DHDcqwsLV1d
EI6knpaUStOb4JEiTEJHVPqVdW3gatIB2G1YiBL0dMblbZLNnU3VQoGTG15oWnxjxWsA2GLyHdCn
gyoqFDGZn9Zr9a/h2TntdVz5rkSGRzJo6xKhjoj4kraDOJbQAcP5BADEbxgM1NQ9DimSz/T/ddcP
T8SacH1AbQdODiAD5OGZ/y1hjyfFMVZ6P+MS72zpQIpjfRjTHlYBQlkrAJ1oS3dlqR+DxdTJdnzJ
lT8OSEBxjvveFo2Xync4ejRviuFJwSplKIOGcTjfwYeUiK9SK6up8UYjqGRj0TLPoYwjewLUT0r4
oqRmr1TZ4xMNQsHDeO8VMBrmF0pTr2XzDWlm1VfA2Zo7fS97T6sOqHUCEXqDh5ocoXXOn+eTsHUW
tnx4p8jYJpdlPcYVO7qMefk0muGA3ikDsLX2LgLieU/n4scD9+DS77hSwOiW+T0GE64pZ36dE9/t
65SeD57/QcMAxuQuJ8hOnB+ICzICOp5U6aC+4R9ZERKpQlwwmb+hbxhFE1vuzSkZ8/vCzE4qi6jR
upFwK17vY2fyEdGsU1KtU64brA273eiLzJOcXk4umAxXQxB5eTf4s7YKu4eI6kknEhSXrpQs3KIs
QhKRmwQtJrB8d8f9C0oY0KXH+By/aGH8tNo1k0RFY4CLFnf3I58Y+qNpuI14/WORlR9B5J43bWFs
TO9tyMAyv5TrLU1dmkm223a7fB5AolGHuTiSSshTKwvSND47XAVzAHaaQg0JncGnLyHce5Ypdp30
vcU2/iO6wE6GSygshlD5B7i4qpgnqFrynvn/NK7GlyR5u/iytJdrc1Np2s0Nz3XEBLIKoUspUU79
sZuPzTrz/FR01DQ5k+iztRmXDpKXMUuuNHTfTMYQtx0zUvmMwlsN2+2Ucze+JyuFAML50AdGqgsC
t1rwbYuH8d0E6W8jNd/8R7duLQMJbqPvoYGi1YjZDkd1Kk7xTip+/t0mfH+5TJIMnUEPdNeGT6uC
ihpOALLKmhnik0TY8tpxmIyGBUE4rYVMO8SEKg+xLBA7WVYeq+p3JJ60hvYjQqQ6hdB9lmjAEgKN
tHL4Msis5AtiV2F564c3JijsZS5n7qqXvH/bCUOLZ2oibSrF28lcVknyjjrBXplh5draeMMuhIwT
sSS2izI7ZJf/Gi0sESCuY1E4C0DP0qLuFziqUNYWYD1ehQBFXgUCGo6OlvY+w2uJPiB0ybm7QUKP
HTtURgdkb2eQYBEIcEynbduW2I8MUId8UAOuuTsGdia/DEb2tIh2e2LFK2Og+ShI/2MRMl1SvIQI
CDHYi6dFtKzc4eKZRJ1nWRYQ+Tkc2RYA7oM4oo1lcDjq7CNhpPY3TjHhGDpkKHtWclv41vNckaEs
9x6aTQ0kpQ5GmxuCrW4el7AaMD6mw9VqJM7ZhgTN78973n3WE440cX3oo0igGrtb00pj5jreu8Ds
Uljw3avRlGvfNhG8HEMNrmoN8PUUUQ+9y0SxgMKX8olE09Lh5C6/kMhdAEMITdF9hKR+saayINcl
2S4KodcQoZdi19GE7OS6sZxP1q2ThAIK2P3bxwS0fUEYOrt5WnyEAJhPpTNo6t7WU8kODkt0MHpo
YZnvfBPziuO7S/E5gelwKgweB3ZNKpNCo/q/FoGUaRGTrgdgNEg6TuvYn1zgAdDYZjJrt6Nvr03R
BkyNnOtip/3u3trrmK0Y1cxomBFPZKX/YyWpJu8OW5w00EQq0IFWSq/vc4gE6FI1MGX/cC5CSS+N
s6cF0CLGR2R2iK80a/T9nuCWAe+RFczOXQkxve1F2XK0XPvPEfHTCGmuNZZTS1VCJB98CoD/Kb68
j8sEorDbCBzuTlgDdw8RqkCtc/LwzxIHdL+tjLt67k9CQaXz3RDu0Ts1yuKe8QTRcn93TI43pKHm
mmZpnynGAlCyZ3D2lef5B48a4w4bAiQA3k7nnS/Qm1dqQttzUypEe1YBzlzIHlynNF1ERQfByMUw
1fiL/a11UkKQ1ueIu3AHXCYLt2jpgC6oQhaxbvF3t3apAAsK2OLIWrObyN6n37nBmmgPz0b+s6jb
pECkOE3fCgcIX8TbqhIxnNj5lxP4D/jOh3FHYEQjTOm0azmxo7ZogLTqHL05kORlYkemzPxirs2M
GH5McvAt1+74vR7BuYeLH+WQtUyZ+gDq1/OiAPfFSoJmnVJ9sd4wfQltuSQ6c56fp1SJJlOa4hgq
po6TrecLqGzGCZKe6rng4IA4zIhfhdOWEp6K1JW6gZrTgKg/ZIjJr1wVCnSGd4lESdtyQ1CX2XwY
rWL6mnhafJKfyHMYFqI0AUaBQiVDxT2hyel7bzt2CDFfrilfUJq8Pte3KkMN6AmMoRqeG3J2Klm/
tvEPkB6gMpU+7KcBqaYbkKGB8JEI7jrFtarcIHcNOWW1GXht7ZzqI8Mouw7Xx4DqRl2xk3isrAM2
AtA1F1GSdzKNlFWqrSGoUAxTb4e6bYtfgKMcg91hERwOYbBFMNYNj1BkeFS0YGpNVj9nFdrznMaL
M5ixjiasXLl7WtTQXIWpvY8mvZqa2oe6rM5it2KeOY0+b6vXZQt5sVbsoJh8+zPIS5Gm6lPxu0XU
0zhXaS6EKBMQ6nW7tBvpGw3GZ7gOgjKBqBvQlNyIKBJ9MSJ+uUDHR21j6C3AaQidKziEUW4KV14I
fYIiT517vipwAnDCOLXT1s4sJdW5xwC6mCFHQ0Q9HzqSePaM/VdUiHHRZuIgeYvdqINtGPmT4boL
gLg5kLYC4dvklFQdW8BzgG0N61SzdpgbXKfRPWk5Kw5JGJx+G1Mrb5A7CePiH6ZblfcwkyMMKZil
lpnS3n7XPS3AQrgWJzpfavHSM7Xzq0yUX+InSwWz2y9e//nTIaBSJNQBZDVPPBEfyc0xecOy13LT
nxxwJdPVSeeSEeZS4nGZyWSAMjry2w26Itr3gQSobX36FMhBAvIkhmMDHSqCgS4api6IFfSvLMk+
WYFkq7OQWKmIx24zRN2ayDml0LuTxEbscOenAHfOshtltrqY5FKcQYFiN+0ppWmCuW+OXuu32OBa
1g/iJutYV+SysPcWULIt+vP4BLzxcuOtGft8uQNWqqOfWzEt9r5aju9qBglZTB1OSBpk14Nws+X7
b3THUUM5tcKV+OsIGWYVhXMGyrXjzeGrBjBlxPt7TmzUagVge81SX7q6tO//1+5f97IsSy3V63Z8
mNFZJAYzpTZdfiP5ZaNNFQXpfdTCW5Ku6jPTNvfzkLHqVSldrQCDH4Q7bAoSMn6vK+65U4DHvB2y
3NRUgwjjhJ0LdVlSxttLY1lQy3ikW0YWzctdqQTcCEVre4n4vac+FZ4CGlYLtKYeJfcsTEEs4Szy
rITR8pWSk1HeFE1wjeC53COxbSQJ9MAYofrwaXA4ZXrF0Z/Ag9s2Q1vJ2iUVQs6qUEzfeqBmbjAv
X7yc5Lib0vuYHFFvwww1DuWIYraJtAwz1rdF1Mfh/WZ5gJYaNEqsLlDG52bB2Pec47SUpVhQhs8H
yjOXO3ofv80bn4nr5nvkztAZNda6Ot7BMmsaJfvuC7+WtN+QYa0ngDmbBuearPcyE0HaoZf5/vGw
6n7EpLM01+K5cuCIS6QPwX3Y+Q2/ep+dU/SIWx8SlvazTAkfVE1tNBLCt0s65JOWQozxtVIWRTdO
1Co63b4ggPaj9owW5SwteEDptig0tDigclsu4JqRLh8YlQ1O6doio+5hA1a0K5lUA8MsXjG2C0TU
q5kS18d7wp7aL6DxTDvegg/3qIF4P1ESyCuvfJsYLeHnZr4MaQUXdaXklRYJHr19/wu4sGtExFar
gXMFTCTCp7YI+4DH84mMM0aPPWOsWzg6hjfVu04agbRSXK9S6u4jsc9AB5Xcieqsc3uZitkH5+Gz
EaOs8I8+qe3EsaKYKJdBlRgXSYF4YW8s3MpWAOhRuErFDdBQY2nnGX/G6mzYzIIHvu0A2Y3Orx+q
wqNEKJX//tFrfYGCf/0M3Twn9TuvTITgBOK/cGA7dxRXVxBETC2YPrIPcMqkigNJR8A7tZysePrP
8Z+SKy3udstWziqBp/nuCK1ig/McUoP6803BEzrQGG7SKRaIKa+l/vHAgSLpgN2pC+cObsFMtGO8
ugHQOvuG7QAiQxzEC8AdquNByblPmB+V+tLifAl4IsWhe/PWu0egk+nx1KWLItox+qdQKI68Ty8Q
t91FqdAvM3BacfKTwehBCzfxAMp8OQQZvQTGZJQRT6m4ztV8mRVkqDFKGgNefJMOaE3pMnofnRuO
RAaVCPZBHRbshWHMGVEAmVh1YRxL7mzSod6GfWvCKBHbYDnKJ3FjT5TBuGHM+nVrZoA5OekK1kWJ
XbAhRYg0auGe7h99p19AIasIOnsKC+szJlnmTa4pHJ1FEJ5yaRt+6ZuOipL1E7fRuL1ga5+ukMZN
MJfoTBCl7Jg+FYzN8E5hz6JhwRTf85S4aqmeGcFeUYDScF7F3N1aV+FbPAXHT0lOLGpWLAsEPgRG
oqpTkDqqu6ijULQtrcvD6yPEvsm+wna2wpKHZUDMMlvCXDKV3ISfUUI4+LzsK4hYuCRD8VhGzHxp
3dTqnycRi27p0oC/ApGctbw3xMc7hS0o3D1kBhiFYIgZ6wKM++o25QjZ6+Ng80SiiFHUpCZB5n1A
U72YDwz5YnP1k/6nvJ/VSTd7KAGEdE7WNBSnNVBNAT4b1ox6y3q72ZzXhOaBI5aX2HonaSsOY+vW
wsBQyg7phxKnFSEOkwiN6Lwk7ySVdzY0v+3NXMFrchoAzYmYOIistkoH2zcwKr1+05MLnDMMPgkk
vaMRb994jXDj8aANGAIfMnTR6/JSG3LXgMDCTDRuQ9wM5L1nZER+3yenrgCGbLYCQSJ7ltxdrSxH
cp2jlgGzid/uYBcFQz09cdO/6PwCN1qw7N0vvUvdOO+cMYkhfJ2PftdkmbgtPVRs96i3FzZUgAcB
64Q6p6ZJpBM4eW1QfN97xtILlyTSSWe59t46hj5Ns2SX8F4uz6BIfNtR16IyUOza1N0QxaMuGFgT
UqbbjlwouahAKl2zWMLRi5vk2CUFCqHUt7h/vejAzcbKhiPLnrjPVOpiNeLFVZRZ4miP/VBJ8s+e
GmpvSVWmo+Ryuwg7v+sgccKzwOiRcMOXLhNk+Fsu+b68080faCSFvPTiicHhfMNyTmvIgOsxwRJH
/JcN6GU01RvF+V20XZNkAmbqLdmUSFfL0RdD3NfAXleIOrXadV3/4RDv31/cOyTku/lTQu5Jl4YA
7euzMEjrdX9WE+kr3SPSpjvQlVHmZz/A75NjWPXCbsEVG0uB3IFvme55KlAHebm5jHE3xr7eIuM9
IbAYDKV0S/gdVqyzoBqGYuAqcMj0oTqqvdY1Ozx4TK/bvR6X/M/2OucbV9aNnsw6ROaRYZLwtcp0
d5Gl32saF1GX4nRwaF0OrYOsLhECt14ie08N24CU0O7XXYgCc79PJMiIsJg71Z6Xz+WDkIJW2JuH
ErMNCX5tLiYNNGvxdMkzVcxlMTavSWMEoS5MKULfhwKKnqY4pUWA7q10iR9kfpVaABrSGPO263CJ
Xfv/0d6ZfLxqZrZRJRqXF8reEvdE7EGX/HLP+Zt5/ZxxOfCC7A6+8vSq+t7Z4K5b+7tVVtCq3f7P
+Wo21tlDqAKUBPtRiJrF5U5G/PeKdfpRYLZgGOsB6bCqHpmh0GUuP9l/SYTE7SyroeKaKDvA7EsX
+u5N2i1Wuu88jMSOKrZV4zcvwqgN35ERi3mOqtB3OxPqM3bzPKVPhiun/Na+zIOI5iiyQkE9Qom2
tuEayMNOvfhFtJmklOxtzteR+03dc67gUiRoz8EIiYpZlKZ4v18dEDZSW3uFEvCDWqTl5rbQ+Jnb
OgwwpzS6AIT+zN8vhVpQEN4Ab+8nSaIbzlVaG8VrudyrznFW4I0N3jZpTcobNRCChx/iQUj5KGmR
kSZBseBpjuDwLp4KgIc0JFGGChEzK9zqpmlEIZU/bmXj+F8V2A95sGU9U1Pc/G9P9UtTyc33yEso
zgkFhIYQfMZim3Y7chPiLoo8nQi4TE2r0hW3B0nnxLoqRnYgranZw6YowRwjsowOpTzrJYNQ7DUe
rejfZpn6NdX586uFFYggZkflv/asA2MiebcVzA2yfLZR0IWbYNURedxdncMq3PXGmt9ccsRZt8QX
VMe8dE+RVxLq0QHx7+wvBFGibK7xT4q+v9NGC2Qh/kqwHoPA0mWBzxoyKVwGAzCtE1nR3mTRS8Ka
tyoQ3aSqoeFFPR45Wv4WikM7xC1CWW4RcJ1Kerspy0MibPmoOq9NC2nJRBhWfrcdl2N+tBEauxXB
SAXKspqb1fp+w40OMxPQT0GubBPidGhCEwYLEiCjlGxzSnH+9VLHkMOWnK/lT+KBA13GDq+CmOA7
b/Tl5pjQvFsPRrujlYqzJP11dMXLSxyGqjxpwPvWe3Xf5bH410VVU0Oj6sSM/Vilu79Yh5d6+ojn
EV1uPU/Ifo6RzzdRHiDQCJ3Pz8S8rcA+rP96iZuMjAQPt5JU998HlDyAu26hp/gorN5j4VrUGS5E
wCwnpFI/MefnV2vth7nTkDDS/vbOKAMaEQzafgmdLblgxGYkpl3S4CHeJeX2pbSjfi+JRzoKBOzI
S3ih1RiKAZMM39NzaTF/98dFzSKDtQ9IUpxogcssjPTlHPlDgwF1NeZlIDwQz3yd5Rirbln4EHF2
eyHFA+1imXFi7zxXsoL2eGcvf08bykRaadLamYiwhRigK2LXkQwukeJBygkjFsQE/5sJ80XIkPIe
JPGXU9/l9ajbYjo6ZozYmJwKPobosK6AUG4MEANm9TsvwJpR4Of4R2VKtCe0dXho8oJ7KGxQF+kA
6QvQhjbc8WO+GBPy+kCUn0sZ+HOraLQBnqjU9bOPPeVevhHdV43xRjV6UuVVY6f5mvV2feygOVKR
bjXIl5mAozY6JljIrNQlGIYS4rcCXdnslD7J5uwuBpFHoTkPzYMKXHkGF6qk1hZlSn6BvoREVdoD
MjjSrmYYviKZHnJOHFhqdKYjnStPXAi5SVsIEv859MXo0uJF/qu4LFikHXxKcWQF8+mflwGCwu/i
KBCv5WSWz+mqbZBNJDfqs3eOSmdyOmwp/O87FGNUHOMOVHVxNsIJse3ZsVhrksXNcd36hmDC7C6I
0/QRz7XjSxtrCSzES3cteirNtn0DrWnS2J0DyGdFCUlO+KW5PfHdoMSh8Q8dqqUVIjojDomi/UjA
tvCU+CSi9x0WYwzVuX/jyLe8grSPEx8/Y3k5uuk8HvTDyDJdcihTj7ntwW/mriC4C/eCOUZpyK8d
CT4xS6nvETLe0/wRTpo6u/c+C6JKJXAGhXEH+PVGiPMMSgrrSsumVNQ00Z0OW0ez4101TEWVyF2X
DCFdLgV30ZYxKlqKHj0SomLgGEN6JfWlrxzZyFj+j3ElFDIPVWo36N/mRq/kEJXIAKKB4Pyb2Y9r
l6nJRM8Zj/sQB2C2hgqgTzyxybDJOqhc6gHpIS3xj+0zK3JuJuQaO0NPY235Ssiz4RGRUu1w3SwQ
CtyTbCYbsILbMpVPsJPhsLDtjYaZi3fJCuBTrEmzTHPldw3tM+viNzXaOiz835mBEugHfGt3/+31
YLzCKsxWPbVaMSQmOETZD3zFafDofCYaZaSpsjHkUsBcT3uXOYDmcXg/NEYIcpAnL//YUjar7NLn
JQtXQ7vP8SqRoOdxRRSB0GvkIGx+Ri7QYlDj8Vjv2ecZFNTeqnDi9yTgqXo3KhLTlrisZSae14lC
ObnN/8j0zbFBJdZoaNzXZFPIjmLkNs+B/YZ5dzDYkO+NeWtWjqZYq5jITIwiqhPv/RR8JOJG4Ypl
6ovbW84lK1FgVp+78r9SBtr96pfQqctLQrqdsWxcYcp6YU1gFvOnruCyy/V4jEpPEP6XQXippzeO
R9F48FOKwbe2+ycKez6jP7UVljzGGlQgSDKLiDE4yyKzU/Ic4+Pf1qZtwOYAr5huBtj1LK0drZEy
HrnTg90yiWnnUc1gE8ED6Cas6jYs84gTZLolXv4hEoTcg0sFLw9DRQ/JYRTgi1kZG6LZriOIPv/0
obbWfF/uzOYHOiVGo349ymIxr5ywdeiePO/hwhBvwS8ERYQDGe2/3bKZpcg6Rc9vJ5KPpxIS/OvF
orEAt/zoaXf2D+19HgkVPnQHYo3SqZfjb6A4kjh4k5ILusjb2gJiEnQ2gu/oiU74slwFksyT9Ew5
KbKGnrFp4uqNxhcdwOPIhzo70bJpJcUU/gKdtEc7ihY2QjMFqqrnDMg922HIN0FjE9HVHdQ0aLsg
fsoJ8jJB633zfQCDEuPpaz31fAhoLNAoCVQm4kndfB163i3qNv3VfRR5jB2rD2ssx7NEcpFnP6OI
/cI/yxeORnQzxikdOpx8yMUgsViblJC3J4nbISHXDsE2U+rM8XSv9Z4bwNOC+CvwSvf/FBUacXEY
zgB3QkIqFkJddZ2IHyHFseNxknsxBw/JZgmaGRi2lvNlyYblaFgJ2tjleLMMxcdjojSSOE41E5VS
U7aLG2CnBKaLgsqx7O7M5h1Dhvalr77R8faGsTf3TaffmpYVwadxV1XFaq/C1+dfNNJWXPkNxBw7
KBLlvMeT/E84ZV71+NiIKL7DiimFJtOmUok2CeAwwbtg/efnAdBtsBe2re642xeIFtCoui94VUdr
E/QxWNVvYl9NXt7zIqVUJ9PGJVHKsCIp7Ax9cXgYxfESNscbbG8MjRapaMJKlDMoulkoFIRjQIRd
25BDXVZuAWrdxSEVAAODu8KoSyWW+PcmGilIIu0G/AHnvKwsYQh00zYvJC7nHoSztrLxNgIJCvUb
Wzx1TEfmggUaUL1t5P7jlby6hjbGkNEwUwNeTz3ANnCRvyWYrygYlJNnYbxATTdYxhsbCBw5CMUq
gCPeWTo2KpngUr96GELZoxPICPOA7r/pfPMhYvyRjjK+3QmOS1Chuxnm9b005NYGjLqV/IPPPcJk
lTGsgxPaMcdnqHiRXu2W/2x9kx0kXQ3jTZfuZPQUlXQlMd2SbXl/4NaGp94P0N6tvRQd8zIfjDFK
bywjeAQqZwX9qRU9icDW/Mmfgxghz82KWXbFLnh5NKdCO5rlAmivqYqZZfxnLNXlLp8ejmlP8aiv
8gQ9mh2+c8W2JGqc/1CM+LsN7szTZpHiEA+XlZtOIL43kdETFWKBSYCNPEhVu4nv1cV9Xgtun+SA
vzEyedekefhWTWADw9cPDZBy+BKyGtGjyga9lg6qA2JRN6k0cNKuOaKDgyjSST2lyz2q3Fgx6i4X
fDUn4vnzlie2D3svehCFr+0cyaTrW4J6WQOnOJN5A76tamB/D6hnqG9ECLjEwUIYdePW5MCkVUf+
Pprmx1ENT38Fg2poXs1I/ATLqZEPq/QLXqIHStHxCW8QRSAapNHK+rPHidzM/uB6eeaLccMj24n9
jBNX/eYrmgC5qNwv2r07JCax2S+WlRB8LCFPKQOctPcl+/S7NKzIqQkmfOoEyhx7CLF32c+9El1/
pbskICTJrGAhCKWQkaKsPBgvMOcgBU+IHmro4R4Gfi2aVQOmTvQGPex0+UJMAQR2ytZ2BP7iC28N
jG3Ran+qBZQbIjLuMFcP8Hqha4+m15NsAhHiRMu5nelE93aQx7MrTriFysXpy17CZoasoy9ouxVQ
ALUV16YJJm/8BpP9O09fADnmphaVAkPOzROLK34Qd86VoM55W7EQyCfhDBDir91d02xQCYcrHOqI
bgmwWxqT+ezb6vQaF0l/22wsNLNWFNRAiq6tqFU+wSis33La5uGVwCrmX940d7cH2FQl7NbOWtkw
TKKTkRt1+iFSP1CqG/FgVBYeXlhDmcOA7x0EkWbq0RLFpoJEIWInMkwgOReQx3tgEiuwm3FJu3ex
h8T84XlBWoLy5+MWcSNpYhiskEep4MXbhtPYpydSiD8BzZo2d1xtGZt7AHbzlm/9D5BaDJ3mWAas
7AcTmoHegOIXIhkf+exGC8XA7QJsI3oJzFq8M8QE4Epdy1dprjRGzRRU+wMN+N+aOJj13LbjHH3S
kAq/6CIrcLTfoMnVWTXBnn9050MJjqnl8HiCirYGqFgxD+lAGSncqDSPGv5gDg6qo9UOkcrrK5ro
a66ZID/sRdVYRGLM9/Zpk3+AaMieKIh7Yb5Voqc58sT6HnMeezBTzTJt9pNUp4+8Bj9gJ7mzJOob
8ZuaLxpInSkc2Zg3/TWbTMOc6nRm47EW6rcKoVsCOSR9SL8sR3CH57I8cP4nEiRt9BqKmowVZpf+
yIjLPO4L/7GyR2iHZI73F+s5mWDwE9J+HFkxLn8V3TbiwV0vY03uJILtc5zJUjMvK3YdXOIIWVGy
symTztTu6waTo8LRDgNcv95SIUsLJPJzN6UHWdUw1sGZPxfa+lFASHhMlFUIY+xQQq02QGGWnb6N
by2gefp5LnruFlZmw4GuzoX4fwt6OOlN3ZNuPIdaADvP4V8nzNAdCVgf9d3RkiNEu2l+hgcMeuj4
D4jV8UR+glAM6YqIrjLl/EETQ9guRjf+hByp/r5Fvpl8xFcLC/El50+bzjufhpY35LVWv3K0X6Ku
sryyNmNIn5OgKw5aCmf969x/1lqKIYxaQqLDOiaaCvY9Zxd1y2OYwwjC4DVpQa69o9uwfzVrDxMM
cdrPS1RnEOjaTyrpSzmYf8KAjV3Xg8Lyj3P+MNilAoLfwuYr5aTgE1TJMW5Y4ATgCihhySzChVuj
5x0obSmt1UeL11G4r8z3hN6S6m4kwK38BTf/LpPqWnMq/wTPYQ5dp4XtsMgFoSZoI59o/YFutOZv
hshe9KhwxfMPm24bW3HEn4sigD4Ew9naLlcwC4bzaE8zMbc5VXPDjrgc+alxW7JwAL7jC0mFMx5A
6ogKEO8SFWIiu8Uc16Pmoeknl2kdKbWFLZDg+Q1cA3GmZ2pKwAp0ELSzJuyW9KX4fEixlDKcWlpV
JVmfg5paVSyVGx1uMrLt2u9rgFy7Owev8GBj1GkKiUr0Tz4VohxoX1mpcInQ7yxzu+p0Jwf76A4C
Cc1ZhGWGgR/xa4xcFvRrrvrpvNDZ1q60pQN0w6ipMsU0C2uJXiH/Gu19PA9WZPTEy/WSOWj3078j
4WKZ+00hgWLEOkWKHsFwH+XBxbiwq9e19LV5ZvCgHuNiAUeKkRFZQB/qYhotT058V8w6I9/aHEEb
633JCh7MFtPufLk4dEvHJmXwhi5sCb7VcSLgfkaZzJxoSi+EN5ELWZS3ppMXw9ZtHWP2XDqguPa9
1F/FLb+gBTfnTf1sCbejangTNHj7HvxVyuV4tAYiuHkZxJi6kZH4gww14evaCSb73gBc8Shjp+nE
ulI/zyOJYHqEzYRW0F5Cn0ib+cE+/ag2qhbz/9oY8FgoDnHhitgsgrQTim0wVcoI283dWcrKFbkH
dk3OOlMLsR9/eFyEZqpvez0/O2mm4HrMzOwVfb2Z84VRprda66JfzMqQTHfzEyUDVbYyK28FRcmW
7PzUyimwo5N9TGBFoDBUMtgYLo/QokcGVjRHGjZjtF665DKkr7ofzo8QYupFTLJLFNcu9OO8cq0W
Opnwbz4CCJqAXN8SGrxl2EmqDCaDu4kBS23SPlJDe0FriHUf7Cma7WkFS7+jtfhch+ismad+gpom
sLExkW+zF3AqEQS7udo2SXB8uzOV/1HuzbfEDvWIINc3rMxpRNZTgBAdorVJ/3Pymeit1A5Tvv6+
PyixXL2ulA3EasTuN2YnNqIOrPhuuIb1ZwN4Z1fgny/x7F0GGsjcq5tEp9mTcB1Fg5thsbfOkPr9
OWb44hgelok7pln812N4VgohifWmISnBpUcGZE3peOSVAUrUQog/YwCxszqWBAQTkpHvSJRxfhwv
tuoDV1mRjgpujE/Uz8SgLQJdF0LjhVdB5mZKZod1Qr+0iEN+CXxu5g/i3Xmtf4877TX/Knss5gpq
yYX6LfxcBnwkC+89glAPzkCR47bWRd8StOTTHyFvKWmouH8r5biPgtD86pOtY/5jtmMyheZZg9zJ
5LTQd5bAWXjxm7KA6kj9r8Ja3M0805uWC1vKal3xnuSFLdNc3D4QhHYLPbacMyvV82xF2KbaQNf8
2RhZRiOw1QL/JxEwO3swh+BQMHAKppN5R9vsNEOCAeTAfTgREb7k5b5ypqy9tuckz67/AU/QY1qy
wPsWPMRaiiO7W1rnBEpAG5fcFKsk1i3EetOjvASFgwUgKBZNw9P9sgDfslq24Txd9FQs4jCPP9UG
xAgOhVRBBUjzPw78slZH2gcBYxnOOGLJ9+TEGOUpLlGYyDlPVR21alpXYlFsSFwukM1LoqWFar9j
RWc3YQSN8aFP5VJAlKB1AK6L34bpikFXUnu3xiFS4Cm123wNKcP62ontSxs3shF9juYkJB+VIxBq
+yljEOxnL1giGFnOWSd7aB6ozVN5lv4bcJNLjDkTc+mGrh6FmKjTrLM1pPvl51cWO4F1TzSztRTW
1pNWN+8OUSY+HDsYTtV8xREgyRqZdRRU3gQQ5tw9H5DjyJphCGl6bgk1VlISZLg1KGVJiJvJHJoF
NeYNh1zXyrBNY9239TLmPu1vH55TJUftVgf7wI5hOio14GLx2IbgFlymUY/iqqxaL7750xdqIew2
e26xPY+k8uGSErtOxalcfkk6rEX9G4kKjvTn6mdLix0LP+jD1f3eicAkb+dzfoL47A6gfliA5NQ8
yeHU7Rc62gl+p5L1p2sF/oXQBXhfvRshawk1D7qi/4CB9fiXdznhnOTIVTThahneuH3gmRd0KPLB
2wUqwyurAaX8STRuT9qqsV3ILJKjWjjH2xo15cauffbAgf51jWXVQJAFb4Aw4i2ieCYIGclsfKx2
SUQtbQ1tJWjl7dDtX7DPZCvVGbNbOHDTlb1gOXnrJjHLdEPuC9YLQUuATnrXInlJDCgbK82XTx1N
c+bVYPfA9uwBWPg5z6y4Gg9LT3I2G6ES607v3HdaJM6AdgwePfkWaZZ36rN53q7R7FYgFoQVBM7u
S92JTXPmN9SSinQMxgVpHN/jrMtTqVkW3EDX/j9kDkVcmJOAWsY9HLYQDK3oWVIXOyaw/Ga1KplN
AaRGqqwrBBJgdSKliHmTiAx/xq+N9owJqBrAmWAqoeoAfw5nUfpRe67CNbjneaqcj1lemPY7+n5h
CIK9+OpbHU3olrsl5xvxgbStAvXtB6055jMj9WACHb28xUsRkG6ffh/r0e511MEUrJHYnk2RuOCK
2rrMiC6hkj8aE5f7vs0M1ngB0M3j2p84Nu/J5+44rY3kVq6CkhzAfxRhjx+4jTJd1Xyvl+w+skAq
2CDhFSOS+192PqswL6BgS6/GzfEYsPbScbPm3N/TMrd9zzAs+ruC/k1ApunOIvAMQvqTozSsKa4V
hQTgKJyZmiNNFNDPZbrrBzM8Xuu4dLe0KFmJlBGBPAhQWXnGT3cQmUyAnDFzTOTRSB3siOpOPgXD
m+4Urd6oIT2CL/dRDsMQDP84spAkbUxjMsIoqKNLnegip4ZrzNROW8RoqDqaQAVWx/bQ6/BB3Hjx
Yt7rHy1k4xk6bS6enflw/7L1/EqlFOxiGrimlluS5qz+eeB4RMcqdV13S26/41tFuKunJllBCY3o
jI6oBF7u2FtrAYNUoTkpqAnhxKaTq0kUogwcchAjUQD3do2uCFveg0wcV1eGrehnfVNCP2y3Vgsb
FtlXpizF6e43XNWZVgKUB+cZyDamEBk2KKgMmetrAim2PYelp/x326ZuGzr8tWEPfdVx6+Xt4Ts7
4TZj31o92mDKUex++NViUR/3F9GuQXB1rDOropMMQGvlsHdudM02FYqCudHoB5oue2prHiE35lQ8
ZZ6JdGY1e4LTlnbrycSaNSA8Q/RL5uKdRpNNbhuzGi3liSpvYGa3kAHaraoyzhC3ANoh5blNEZXT
In21YIqSBukal4US9/pqDP01TAZxeAKFsK1rCPMvUnA916SYHrp5rhE+pKhCZBa+FY3UnlElGcVU
zV/mpPP5zf56Y+SMjvo0fYVLY1u+ZOO3mnanvwBBJtM0m62ajwFh72WDTOCncX7+u78h67fRmoK1
ij6EQyVnRyk/Peg5K6sZI+ENA9RNlgPa0c6tO3BzFIrr4Wp17kVR6rTw70M44mn0wf0zdc/JO0Ee
h+tUXnutrcB9nOtwvmxd44fw2/oQzZjzGbXyk4WbxmBvebB16Ix/6zKcPqlxWtEI8w0BaEBfwxQ5
1NqDxMgrpfjcInPzNXg6/m/i3aWyut8h3Li/lAmIMUDznn3Rbnx5cqQ6qmfB9t55HkXWNz/R2MV1
o4/pjdDdum+5frSK70PDkZ9OtnOOUllxLl7NSNF4I5Q28IdnmcDmWz6AGttcjh8MFq5NSwjVsN/O
LBh5+gE77Ur/sDBn4bmj4SUWPgHG1CksWzXSuZeoB2g9HbsE85dWXil55Qfi1LOCHRyVKbVse+1E
71522DId0763voi5y2MmAs4xvRyIIv/PAFT9FPR0eF9n74FB2nUFRCFiO1nqkxiJYpiMmyszj95N
DlGB4cTj4yiPubJ+XC5O115+PjKNty+KDkXxwWuz4EepQC/4Xa4NFpu3xE+opGGCFjZroDSsEOXR
t8sZR6N/GM1fU/5YIhmTThJDTqkvC2J1Ydhm1icdOIn+BP8DzeXnRiBNWsdf+G4T2Vn4ZhD3fc1A
C+NCgk6uQYcJMsHJp7S8sQcLsmhnokUpOWeh0oQ8ssbxnNFStGxZu2KRB0omIqJaqdmp/6y4xyn1
pua8bYUnv/cQ71Usnq8+QMwOjevrNsXB3iV+XjrG+fVJW23Ohdn3a7hjzUIXDyKgt5CkLvlrif42
gw9WdldwD0muCJAwMtlVml2uCKrtR2nMEY8MM2074U/IyReVntnKIlluFZqkcsi4hHF9H68LHUQb
cM2qroyVQt+MFzRuiDIEX/uD/h15/7TsoYBR/+Au7W4uKzTCMKv0jjzrb1hGp8dMjXYivA3NGdJ9
MK7gGOm0FdX3hVJ1NhOPVjgMiEf5j5BQcIwl13VHe0Bdugo1MSDXeMUwVbiAb7A+VF1hhfAC45Fv
GIQcxzBYDF7cBy79ub0A47cud+ygr3x1uRbzLXZhV+IsE4OHE6PgKOFuegqbOE8zb5+18m1XvrRN
ehhi/FjGXrMk5NmflQ6ooxiyJk2vqGIgRwxg3/dCPdsDBKsATa+RHgL+ibS8jbUYfDwz7psJghha
x6EHR1lERcfpHSwFdTH1YkMgE2YjjrOJq3K764THCpUnle623f+ei7yqE2n3UVZuA57FLt2xwH6x
dQW51zNKw9hNVbt9hY9Ci+4aX75Q2xd4C/ZT6x7hymnL1GKL5oC2tn6YEqcku4HwoDYZ2UJq9O87
Wq0EvsDLeD/W5Hik2/sw9me2KxJpW6lYnsbstJuGI9IF/0VaWsa3TwDvPYc6XMq4wQvWSljuBbnT
lVQOaoxm9M27sCCB+Kclq+3cVHJ0hKmxhwnYsFf+CZ39F1nzrwszp9dTgUkMZVgtQfou7p37V/2H
u2+xYugAfftcVPSFOLgPEmjngh0fmEofKgYkEv037BUXqhbOSD3daV2C+/lu9TBub0bylee1kF0d
qu9gD4vJfhQSf0fkZZJh57edWJ99AIWV7slI/iixYIqBGZr798I3a4dEy5mqWs+k06OTiwvyL1E3
hk641kgma5Qockl9OASBGBHWpjTWICh5tC8RDzJpumbgyGcghQJ6zNXlM7R2vKUlix28M4wuSJHU
cUzX1N9wQBoJ9Hnt6ZvNfnTgu8DWdoQ3Cz3MzuQG7KmoeFlC/VZfUKTPQW8zpvNa8eNd7o9urjKv
LuYzpT3+uBqtFdFB53hjT5zLHt7dcLkrMoF0iNbQnmHe+l4Uk1UVhJs63pGPvyodE/pEMYqySUkT
FKk2dq4/nAmN8popET5I2LoWbvn7HCLKwbf87aUA1FTlcTiXWb75bG8HwbKp2mRcbWWP5OkkxgnG
8LVii4gOU/FhkC2QaBGJXiO8m2QHY99VLpX41rtv/FsQy5uVExJ50y5YHfIjxUDbH7cMJwW/y0nU
p4SLr/5Wr79Z1UkS6hmFhTo+VS47vOmMDwegYHZ/gy4hSnMTHE1K7MiIhGy6yLAhIQL5KJ2+mG+W
qIcw7fGF03VuZAO+43lItTTbBykKWkWNHDmzyYwtU5JPZh5/nJtzACtliOUvHarkGMfZyUFb0JlC
mujzVbqXQSTSj53P6RtzYcbXVRyONhHE418JV5SWRieEw28z32Cy9ttl2AMtiVXRAs5ebXAQq8hO
cAzpbnU2ArfnKJZQXfVHNVw75tHLNst/uxz9cAGYzub0HokVkbv+bpuvcC6oD2cI8afx4ga1yYGU
5LBxtoeI21N/fRlzybL/dTT68qTwmiEqZU26z9nLXLrgOXxERMcAXW2sLgEr4MjzkF4Ip+ZV/Eb+
JOww0TpjVpwfRgxiVh27gqZd+Tr0JeLuLeKelZfeVlQdPz/WTTPU6PZAJHlG5NHsaDnNovdKxzYw
pWS3Md9x9rbKHvz7rAe4Gy1VcjR9eLiWf25PAPEONeC7/3v0zEjlj6WtIKyG2UXwcj9PVibaNn5b
leW85gNUdqDBRHJJSD7gUMap/f3Yr94Uvq5xnkp7OF65W5u4oGd3Ulbz/yP5KNeJ/IbXm0R25lN9
TviH2WD70tujdm6d+ph1eS/wayZb3R2FsOfPrHEc+oSq1EfcSUrZlsqZ+4BMeH98CTfnJx1D3b6G
SpeTI0Z7j0OxCetgjxHEBg46UQiddHKndADnQp3jS4YJeWUV3J6bOY7UYR+cGAD/bIh9j8btbHsT
DOMvp4NphJonIjvCMgjBfZ4WkoZm81LjK5xKg1Wwgr7bxuhNd6A4srFLRNbQnIfBtyU2LQsplmki
fHYj4ZgB9p38ISfiihMjr2FczWs6HIQ7eLVgzOnUEOk5WPi4DNemPxaMYZSbT5LKD+KcQVjvfRTw
UXL/jctRP871ij/Rt5NWuevZjP0v0HzJxUwZVP5CdRCb/eGxpNAYmY5KLX3HtX7EGtwk+0x+4owL
oVd/CvXhqi27KZl/2PAoPubLWja7Be1tlnGkqYL5V3Jg5F9kZDxAXxKnIF+ibdBfBdnIBVQpExu3
bIZOHJO6tJBDbFKCaLNZo7SmzzVG8XWzCPDTQedB5ngUU+F20Guvcj2TRTyu7ukmMbsUsVwf0CpU
unAT2WC7ReBcm2D/Ay1yU515c/gBaUDkDT7mwYth01OLOJl3ARMLrVhiTwn31jdCAPRpZPyYkE0c
ATR/t+TQlPCQVIBuUT67XeB2bmJTQrnmJ1072R0yqn1YTxzrNiqRPU+m/5SI1Zd1pcER4Q7atu7W
Rri4KPuBfM2OVtMEumIp9CZEC5TP3V/0oZ0AlA1DSKGQmFCEfRYzqsyJI1Sd+B83VC5wZtFl55za
jTVFl/IP803CojVPxdzqPDxZbf25+h+Ehyke59FsAvlFbAF0CpoGd7to0SAnGBmYA6rLPMEsu5rr
edXn/KRecCQMpu7l/EE+wN/WaQ5WrQ3rz3D6VFWdqRAHWvTFJw6mARBZa/lhLhy8YgTBuyfXPZZm
wA4UxUGsH8tvSAx29cX0ZG05IqDU4Zf5TwJUwyWDl5U8qi/3eL7sl8Y+UAvQ1smIv19BaU/mu+pc
0sJb3Lte9AcXnOiyE2QLGafztS06dlENU0EqZYtouTQtr6C0YEyQO2BRGew/xPilCDna7gD9MfNi
Py2rG2KgPGCY3PgPUUKilSvL9/DDQwDHWk1+aMRtVrJvM5RaGu7J4byE/ZjXFeMfvwVSTFatK+1U
mWRTHKqn9uxw6HD148U763ACZXbEWaRSpib6E50sgEgVuwwuyohtxh9DbWlouYAqr9JZ/bBXktyB
Rp2pZQxqtt/mTwmXayVmyBxEQ+NwpSZ1255Xayegvzih+5z2zBxMZlVhA0QpG/4fiuXDQcPufVvI
2hwGYpk1Q1CvyJ8ZtN40omzKv0S9EbN634t92Z1+O0mtU62iTDa+atgqjN5Wul6/088TDHCf454K
dvDLtXhyrAIufQOp/BYctkbHsvjzv+Rf3xY3dpyELJzejOw1CsVOyRKHE3J2zREQihf+5Yt27nNP
pe6WEEcP77rgMRDyiF/9KgFFVWPXDkRPVuVIPXG0jjEADmwMNV32OAHhfcH4/wBSonyPA8ckQBAM
Y76nSkzhkAsuJVkxea5YXI/HZfm4v/sPUyRQbha9uc6LWgWRCKkDqdnDEAMJLyOm0CMLad36nkWw
PxSIgt8OvyFAas8X9E+Q+S7DofBdYlrbNRp2Ay2KZ8/Gyh7ODb0JcG6qtknoH6xh+QIx9nqkKEtr
8AITHkmWRDGhsiDa7bVeBut/4j6U00pZw2Bej4xItS1gTzXoLz8NRNJAZ3NrMsOfGtQ0Y5R6piRS
4aZVrtFYHpuhBUk+n+aOIoOAm9ewmfS5KDKiCEdioHOeeEf8KPuxrwNqevswDJ+EQ89Zd6kROb6A
Vru+kH8UPllxKKOoz71YHMDZIZ4aEJgO1GrOwunRUdNLHebIlXpYEhFH78JeRVvq28Xd587A4WS7
mOnOWILmBRQFc0zyj5pdRFMJoLU9lUzZnFhNlxCyIIhwiQyWpTJ+aU4OhsWRii+LqPPA4L+siCFC
qc/ZM31/uzh2mMUVNVO1v0yV89wqFJ1C/trxrFG0QvNJD1u8MXSmw+lxwd/uDvotH9Q0C/ppLTn+
ysNlFlQ3O9CvWDIKcFDzUHyIPaKkbqafkfmFXaXFokjVQCeRGXZhSfrgxp6koo6LxiWNwYjfwXrz
3PWGElNoTYzElrsUkI24FFTF4JTTi3BGXNxCRxiWoh5W3NPKmUNo/yiF91e/Fo1iP1z1ZvUCSlNg
+Y787GQv3f92AxoBWujAGoWbNVvy2oNghgDst0/xhxIGvWbtuqx3YGA8B6riNEKHKMO2kzQEMvck
MW2aID463Hzlp661RwaixUDP1i1B+nqeY3n3EgCqYVFLq7KewVzTSQDtmV8auIJIEamLwU0/Eyi5
K+gROyQGZz/ieuDLa8HtrY/Lpl7Q6xho0bRyswP0aoXdT+8vvVRVKbxsjImtORUdrNpCmVregfwu
1zmQJ8m+uT2bTlZqLrDuSKLQugUOW5xy+wlav6tv7GVmU0esUiPC5kdvLJMOX9Wb2dw5sdZs7BeJ
x3GKozmj0jGmDUxS6e4gRiluNAER+EtDE5Q9ij3zrszWDC5yNLxORSodPqLhRA8uj57YmqesVO8e
SmAbIoe0C6oAUNRifAB+DUEtlm7hW6N/Eo5H4GBFjhAry9KuisJHgU07zzXl/fHLk8ZsdTG9meXB
0oL5Tt0rDoDjTw055olRWbssGM+T5rhy/VcC5dK302dKZlj3NrlSLsqf0/WDMW2cUZ96bPgrZWrP
HgRnvRNwt18aDkA4xXeuTEe+k5N5HrgHfixEXtHUCr4vgZOBXmS91TkcfBgc8xXwyJCm6HsE50Ey
kqGJNqm2gJrk4YiKWQRW1IsQmrMNDsEnmos4/o/7BrGJfZnVz0O8V00JCXqVzb4hWxR6PsKW32zT
Ty3KhcCgiAqOwzsDlGA4ZlMnfS0v9Zkkg1FTfuAgCHXzO8C5+iJGX2sddzdnQKapNhHXq7IdZKT5
NmNknms1rp+iL7392M5MrkFiiw4wqqRUvGq8VJO9RpknKTg3FPvU3QnPY+diAceECJmXQ4DkMi3S
g7yM6g8Q1f0FM4WNXXwoVetjV20N4T+RTrr6KstZAt0SBp9Jb0ZcSI8f0ETdSoNoqCNvHRhs7kVW
cADfmP0xh5nhfpM7p4y+vKgMcaOVtXWZBPsjRL0bLdRePdCP98gZWeGh5f5wVbG85mJ8z+xgEY/M
u4VBL7kWvKfxL9KEor1BpjGF2oOwvqcMHzWGdiK9/S5StbDW9nzKuiJCM7eubJJfrIIjPn5EDoAa
kmsvnuOj9Sdc93o2n+gwfpy0B0kOS+3QR/pPG20qX0HQZe3roheDcZeQ7sHRUPoDnHRvWHoqTH8s
w+VnaMYlmYvAZ9lwgNDu/NYwJapSLSh50zUSurXafasG/e9unUf6QVnS7hT8Dm7+wfYkDClJKh70
DqmQTHWG60WYYxHxbsCKfwDFVJdhEGCoZDHnTwjfKC5VibnKJ8vxyif1yLjHglvIlpytsmPdWnZ8
tOWTRHitMHHceeYD9kn5CZTz26l34Hq1gP+PEYPiGTTxcfPyD7zELe1wpBqQSEELEhgC+VYCAEaD
WW5MNnieqacfEeg0oH+TAVhkLfUhnf/hS558OQhkce3czFw6P0gSEekFqkTyWq1cQxugwPCWPX3O
NbIxXpqPyOEi5i2CveF/DeCWTGh+NMXfXAOSJN1zn0KnYyzvWJrJNtdaFSpEA4VgXgTJ9DNHBCI/
hJhM6W66/yX8R4GkR8dCNfgSzNlmTPWCb1UiqhbGV2F0LGwkAK59mZmQJWzLXfL5nq9X52jFkh4y
3prhMW1K1lMLmxS4EMjSLPY5QEbltW9pLz5yF3RvzXuE1Tr+l7nILi6jU3CxYV1qOjsvvIr0wdCp
0Vq/KsbiWtCFVfGP+9iUiTSbc/jzeTghlA5wJ9fgtd7lMFI0aJavLT4AJWCn+q0deBaAmXtfkEJY
S3X3sgO/1nUQ5tuO5gmQ4Qwr8qJJC2EOtbG9kMyjvroPoSkDWER9+zVcbBdE7ktLcdIsH0b076oD
2R25Td9AkBvUbjalZjXmTkdyHqH+aDmFgrcMNLuj3lysQb9WxxhL3qfQdIw8GSaRcl5EMq7KhWli
7F3zrhQhwOgGBlGQdpxq5Q9CSitvm3DdtSg0I00TebAqoOt5LV7Q+oM0bv2PP4107gb1IBrVaVWn
KDEFmebPUs+kMrghuRqT0IFAdE7vmrbYAwJtkzimtKvycp/AuAenBVgXPKzYuwnRYBXlrxdDEdwK
oWNTP9oMS3HAk1ufp0yNaqZRI2RzD3CuASekDGZsYhS97CWhkzo36kdCO0jCiY1hAQ1DoWfO9Amk
2Ml/x0Rp0o4abFMEmFlAxKR5ibbOxivBxlcQh/0UPEmK5RFdGhvpUsAlFlUrNkLc8qg28rt2Sonr
JaxUUwc/lIiPim5FH7AiPB0AJmHgLzJCyKPQqJu4YCN2MGKC9K4zYdPadaiXwfmCIzmF5rxM5zSi
nwLsE7//PoCKV0PyHFMUzAjNTwsyq74AsEse/iWxahemV1oEE1kM6PacjNpFaLa0NuCNGwSRoook
j43HRmFgqGwSYtdDX1gpCtvLgEQOjvuSPM9ipkqXSDudmt6sP498A3YI3J3CfLpJriks+4ly4QZR
1LBax1y3YQodjRjp5xnTImoyXfv17DOHg1bX1eatXOqnLF6pakK/cAmMYT2K+egZZ/aOKCBoiw6T
8x2RLopxocsXuV5Si0+r8XreeAhwbq6EM4XP7WTMcgJ5k/4XOqMDse+n4UeaOQiJe3mvvpMtmldj
OyNLSN2B1dE6V6FIEmseBuVPZiz7HI9Ez+LIcSA/GNWV8mwa5LMp+R++eghovOxBl4cGSPp/DBUe
/wvlxD8phi5S5B7+Zm+HT0KOyNuMSeH4GT3jIJl8j9hmp9gyZWoVkZPHK5MdbMsZmNdOzeOHaxrc
OcuDknw6TBzyMNE9SpKlEH5XR7fglLPDVZ8A4HK0gl3Mw0QDClJcgb5FTYSqY3JU6jFhHCfvteGy
8zgH4TJs29a1LkMeOSXWu7f9wPXRGUkQnhOJkbejuQ4JnqyEXw8so/kvDKAQLB1oerVJXNz9XJuQ
meKnnzz6V2v5rIYZrZ719MozuActt8Y68XV0LZsSEvNM9NiaXpqhAmkkCEnZALuf/S7vtM/dqZFD
R1wZUpKH/8x0R/daRzpJ7rMjYARw6fXIprSWp9yisNOvwtCNrN1ExiBi4ei/5CBryKqV2RDKG+5f
uCavivdzyRcZyltwN35yT5e5h+ozqPMn/sbbKKoi1jpjvPt6fBxLQeTMJaYSS49oWqoQFXCQjnPs
a7f2dt0bSCQedyJNz4fTs4JL9qTl2r4DLZysVqht8WTorv2FwtoufzvxEIHGwoxNSO6sk+CSMPKD
NoAcwzT2/Etz05AJ/MqQ2ziBZk1xb7Z5yK+jXKI9SlgXxPwmFYsinQ9oa47nKlwwYA6b9itszddi
Re2Q9I24Q5V0Uw7fUYVnDRNosQAEh0u3CYvLKZZ8jI98fwLfZ9QBC2s3MEBWmd3bymyi4LeoI3rg
5GmZ4s6BhQM1Z2JFKrFV+Y3GnosUHUnTE094TO/GDsK/h9wKtiGdLBvS4Qefp25oSE2Sz0n9sMyN
a+LrIUtNWGChN3dy5IaSbXjHIj09gWyUgrjgM2Ig2RceWKi2JnWstv49CTclmSBdcMYiQyclOKpr
ocKQdTl9UGrQmmAZ+FFD0AuUpLGwBjcdFM0QQ5mrVgkEPF9Xd3qSeMur/b7lCSFka/mKl/bTEyVw
179WhiCm88nr3vW3Gvf580j8X+DG0jUtHPEuZ0Nw4kjs1oTKrRHqBQ86cqZgj2OrQsQPK7ZxF9p5
BKU/+/8bftFPe3DhEEvh28s6MEgHQLyLdneJtJYtyeX5KEKP35etHG64Ngi1dNRV1rFHRWZqyQ9O
P9klYUL7TEj4xLDs1Wul06GPhkCkuV2xYdjKnJuVJUMRfHHWqrzmNb07YmsZL43Gri5HBKwVQNxD
prYTGSSn33TAM3uKKyum2yWVkCtw+hGqjrFmr8r4/B10AL4hgdn4jaFD+Me8vSQ/pUaaXCVc+Q/1
BOMrzyZVdhiAu4fjnomqkzCmFUM3+QdpSI0qPJh/ZPhcKlhmoW5D1Ps/YLRuvCLl+waiUIiaz5bF
UmKgcAiFHBDiQfzB0IsR+ILvdOuawSzfc5jDklYUlg+PqF0WeHW1fqw1Xb9TRG5QwgtU/Azoc5CR
CVc35GO0sis9vOpt/2/2kvdz7wfJjZjwx8IOqSiE7GjCtu/WRss2dabwCGIdpTuGq7z8qfFK7Ggn
kqkSbiT/q5SykG3zT4pa7HU7on91QT2XkBhYcGdN6gRWlDMWz8zJ+0GNnOwt9VZzPHj8uK7gsCtj
eaCYGwQMwEFGCX+vtR42+Ug5yi+TN9POKo7qr3hBoNw4TaylKHtTjqV6C/N1mZVN0ruf3XCHhFKp
yiz3VLOy2yXvpngZ9e3cnWyXgE+djBbAf8BbqQoT3CPStrOjbjtoF9X4dSiZJw2eKRkk7degFSu8
iqG/XwIBjn6gD/HPcRGAo+Bvwncw0zd9J2XLFqqyi0Xync22RcTifvQXNw8Tji6y9iFBKF9T9ewJ
qMYYQkICcNUmWsMhOtS+yjevzI29A5x1RfzG+4YzfEkyHCAfraGeW70FucBNwDMiaNd4tzJ3Fj1C
TEMNrYTQH540FkVN8T8FknRjGc4u/l3fLYuCvPIjlt8jsZSZbSPQIjl+ADfmUBItfoNtrG8SVr4n
KZd6zp05m4be3bn6Uko8owIo1WAPuUZh6Y13/R6HXxpYywq5COLESugGYOmm5pt+pLGALSQk3xgi
k06RrP7dvNraTMZWA3uvuAU58m2r5MACsSPbJ39IuKuG896IiLwQNn7HErBXB0C1oIUxqv6ooLin
kiaZHmRqsZ40/6dIPaV3sq+LkoLhLXpyAW+ZXDZRHU9F8xuTU1F8IvILwwy9SihbkxKfi1GFRpGu
5QwPVwZhYq1s+SmBl743ux44kDJ5CXaJZJ/JS4XGMj836mkM6IivFIjI9WMhoW4ae4/hyOV2zgag
pDt4gVAZVCOByNWi5MnsgYbTgWeINwEV65j0DaonIHInUET7IituTaovHkcedkVDYXYKenfzT367
cuA9RBmPfDe4zOy90rOLyvyv9hNDdK2mP4NEz1GK9nbz2H7QgAJVXrJ1U45dgR3yFEvGJwf69McP
1TIxGOVP18fW/LbF2iYPfa63fYa4thXc9MNUKZt0waNBLT9/0pwnKWENy1takHmbe96wZYWjePA/
HRx8zQa233SDw3cUgG7tu4kQH44vlsoRDMq6zYYhTjpp6LUCanHbsZBxLK6m9khJ0+V2lSlLMtwm
6No/PYysE1krUzXfAbF/PsZrqBaOCvXX6PjMqaSZVddyutZ0lyb69QVEQdEMldcZQIyE9vZUWEEV
EOy4mGvAa0tB8aQrIHXzMjwlaEIYPpkp2/Z4e5SZLJkUO4pdlk+IZSZk1MSUPMMlHbZNZKehy0GU
iW6rtPHZ1szh2LfE0l30UASVeXKYXPQv0d2QBif49sPOz2hfoqFBtr5kUM5Fs3ycoqwyN94bXX80
sXI/7ntZZmM0ySWshKer47OunS707kJoLGzeainG9cxAtw3RDQDd6bOBeR9bqbPsSxnQlge8mJCc
Ex0BXtZRo4vDPnKd9TeGODT3oQCgebKxMv6GGBKZSS4f++evdzrqDskNl2EYyXIDOIt/nuYtNEz7
EJMDOLhFc7o3wxdWoLOAxvJtgwi3+WGCIt7hE4S34iKDWE2BXmoH4bYVZZq9zuuzCGvVVrDpyljO
2TRNEntXiXHPw/B7tIND9vHHZhVdLmSuTeON8U4/wKY891VUP2wCE+T0fv0c82tHK2SFRvw/wG6f
aH7qQrqcbVk/8HBU4A7DnK0uSog8JJi4v5xnYDTbfxYEIpZDPNsCjR4RU+lY70VKPECMUwstbeSk
V4engo34V/dAix/aFi92OcB6Y60RMffEL/aq53YjRPw477qp2Uhqcd401hhqbhuD1wVeGAS2E8Ve
zffFjU/WFxjjQK13mXXapXDljOllSun/KYXs6xK7bHb0ZYtg8ab+1PiUL9PtCy681lLZEjzgZ0Ee
CivmKZq+RcFaDf8lvcvDcUblSJEW0LHn7mkFRMxTRBijJMzkB6kgm7dyXmQdGqG8IYm+sViI6AL4
bpPVj5apCbPi1eGBGen9xMV1Zd7meADGNsJbP2k1M8tJn238hnsCIkWhPEjAUFj7xWIM2nacd6Yw
i4Txw8koK6UcwtTinRBf8Y81r6K0sI7CbYafd5x3TMuYGbc+2Dqji9L+rx/c84mFPd6L7+L3OMwi
fUMSIXQGl/BAwn3YLDHQDwnrTuhxuWD7lMZqbxhkTYVp+G0iAzCu0OdCzVVyzF92TenDAAtlMHkY
d4oxUaizoqZpvcamsw2tF8o5OhX2zqAm56XpYhkj7xfkT6Dn6x25am3Egs0n5kx6Wagmy7sJH7oT
/ru1JjXArQpyET5oLBEnV3byQUGB7xkvqSLCV4ZygQuhzzSbJfd4iU+wvbROXlQEeQOy/KjnLBri
IoxN00zkIDiMXhehUpXKpLA1Y+1M1G8ZPJD+UWKUbQz8Nj5jIthpba69kZGckYDmneUI0OCQgMvM
extcuEGu+G80P/hwsNNjPcA7+iFVm+IJV6Mc7KX9k3c0LchN1I+9r8N+owgLdNel46p9SKgDvAVU
b9twBU4Ze7QyOFNIThiWg0tU9uNFu8A4QrIF+k1vr6OBIckhITLs6jGmMybDmsiiOXz8c156Pqb+
sn06kcRXuoLHD5vbYH513CUCuV3IDDzjPYeEw1VLXmcNjV9Cb2MOF1WIuey5vVxtdNAlxsLmbIXd
B53xLMLc6qRItGILlhEfqR1IqRuKjaBZf2F5Z8V0ceykLHti9+Q+MsEBXcYv6te3nNxBjIZ7GzSc
CDfUn6ej0a05reAtt3BG+hG6fzr9Zgk4y9/d00GsT2i35Z54oCabyDO9gFnINkeYgUrs5qpZysaL
254dxGHBQmEAMGFcw14SnawB2PHG2sMIsFW+Cmrt915lxfb07zoj8OnkWq3R8ixSs98HIca9of+N
tnGtiJ+GOU/uacCkQLSH1VMIrym+NVb9cCYon0NJgLJJSzakq8XTWDwszcFLl4nPuK8baTdwz8qd
picthCL7Ce4Y39XNLcH28cZHXvvs9vyVAQsxGBi3M6NfUxT27UpsT6C0veAQuEh3VEOHKhBor5Ih
9TZUG7hxShjDNrrOeHlSOCH6L5jc9sBjVtGU631eLmTDgfIks+SjqQJRdmAf57mpip/S6qHXxgTr
mDhyvO2ZqYCpV2jgRgHhknPTXQmHcCUpQfZfXMgrx4qtidN/eELGmqDhRv5l+vNnhju2aubg2+KE
fsZlrwZ33oPRJRB7sgAIChiYIBBIBy44g1TABj84pdZQwusM20lHPq0NqTbzvV0TxW1Ou4bBH+d7
wuRuly63jSukd88Mz1lZcBoWklaG9JTYNl+iFY96A9dzQbcJvgOmFdEbSXpF6mnVytWkQNUYucXW
Om9zyVB5Pm7SRy+5+GOR7cmh/NKSyzqDuXPVuabeKp09WlvsnEP04qk7AQ1Cn+deH5tTY6hp43Iy
CGiJ12F3uxl98nBigXRHE+SMXQVQzZSLuwhC9p+dlG7V/ygaJjr3B0brDqlLqw1crhvwlXKFP2N8
TRlDA2CD3N0WSMDF2zTqcKlwI9sotSyf217lPll+4cKtaJi5IZNP2cKD7QliInWTg6VbYXvTIp0N
5SVR0gPTwGnmM/LavfYtKgF1brBTuoKhnqMoHuHtWlca6cyjj4kz4dinMgOFv1PY57OGSvmJgdKf
lFy1275Kpp7e0UPf8jC5hP5/x4QN9kfZPklP2xDSgtEFh+q7ae8Cb4GkynFAz+YkIxkXUnzewXwO
JNeZ4v8dzs1FPhq2qOpCGQz8+tf1hqIam6IYo4bWS+kj4+vMBJiuoMqSKdUJosvv+WvP6k8eVG6R
DX6zGmOF/G9J1AB87Q5/dAezXmkhaCqvCS/qWgx3a8qbqE40JMqvg5dS+e+dHNgScUPbVbVlHkYA
Kgx6KViCHxnQerqkaNr7moCkSvH2tUVxG2qseDRTXJioJgDJh0+x/j6R97buUX4RngXQtr+4nQhU
KRp5KJPab7QK7AI7NLXFTXjhc6a++cIJzVu3lZM5avzuhNjFymIwYFKKiaQ1hmgXYqhO3CEWH/3L
v/lAKY5ZbDz1rkh4rlfy1WZVLB76XAvQPDcMYCC8rr0PXYxoPIlzGN83HfW5nwx1qk/KiwHNwnoQ
hGYH1WmZzwGA//jOwMp39eg3CNVdtJsld6xetTVhmZ7uf4cFNX7J0Im2pPvxGWP9Xgodc5iT1Civ
353RYGY8bclCgz1mjkjSTwixqqtO8zrx2OnqtTZ6vX0GvY1+Grc9MHUfpqTqxT1mhAm15gSy6Ocz
fPeipaNiUwBkqBh1kb+afOzX7DKuXYm+HfBJRs9GoQN7VypS6Q1B1sXXq2C41XAY/Couk3oNNqQN
x2ww9KXk6GHKWEI+jPCf2FIgvOZTncCcWs9xtPSB4/IX8lZKtJovxOsujhzh6RzQqdt2DEw0jI/x
U+DzoCxLd+Exmf2fQMmLs5FgADcKTyI1EsqOiaesCVUiBRZEJBfGl510mO85r4xdlACaOR/6pOSg
oriAsUFwYZfA0o/HgUzT/ulAH1Ty1yFpiqTniwsC8PTObnjm1fUTbSoqymTlXy3oPvhyndNWOgA0
RkYC3KF7XT6cgLOqx8OGqHgstFLW/xjTsMBdtlkT6A96bKXmg/myMi3t1ceWN6Ovgn71MyM88Jq3
Vs9si89xbGrRe8HZa1KQTUSyt/aBoDxVe/29VEO4xEc7MKhNS3j9Yo2ccerxzl++X1WFMzF/u0W4
6TiAgxDCRUWFXEvPPjMK0whV+PDrcL4J6L47lUqx1HHP9mbOxkZtp4pzCVGwP0rYB+ZkVMWvLLHJ
YKlZKoYfLBARDOYpdSQEo4U0hdHCUezUpsITZLpEKeKn4ods3SRHCLipWC89a3cDRFg74C/QUkiI
TS6wCYJeMtDsOyZk2nvYlwkUAp73DUBD0up6vqBw9mn+9Lhyw4GVD+8d6mPy7XKRgrphwDGNfEjC
JKbgNrU1mmfRbtYCkmycBRfqIVW+yVGYwgKBqV+yIdLiw4EOPooJ/i6/faSs00MYyNMDo3MUner5
Vn4dI94kquNYmhtMZZ335F/bHVHC8Nzz06r3WJUiWdMx3GKfHmpen54t1ppL+1iogqRdOA6yFZNw
MH2DA/IckQKGVv+UxCli4fetdsM7rIUrNcZlL0hrVitIeSXQ9vo7uDfT1ZVWRDSpyf4kMaZ8yKK9
bQKHq9t/eKXwIweJ3OSsubZSlcIHvOZhJwN5SF6g1WbHZaYA0SG5ov7FHK30Cvb9GpC5h5hNZ/X5
Ogy6P7HXSyfVMTsEjGk1CduvXdEiZ1Z9FQ38eI3Il0zL+StYgWQUiCxljuo7tUmyfCXl3iHZPNYI
ls43RWs3aRRETGUgX58WId3XOVTtJQNB+LrJk6H8f0Hq4v104pcPAsb45F1ZpgHYv0dbe5TIVBsD
PfS+593BR4ic1vFC/EP/PpyhrJmILF1If6wZEEB6WkFWMQgOME+wtLDGw5/RLQpBINWTctnZyE+Q
zuVtKNP2fKSNkIsBtMfw1vdAO8VrgSgBwTiqnUicQ+4ZYUsn1rUFmsiPB4IdiPlzNIlu0LFRZ9lG
6PQhEoNGzI61rS9Q+DN8hg5G3Oz1ud/7LSLYMh3nkCgaBYAg9b6XGWKpOlHBIUo7Gjf9r3xCgAxQ
3lgP4WmVufhJbsPafMFdlg2vrJBT+p8jfzlucqxz/30nCei90oT7zpSNZ2Nmb+lLZtHnS9U1AFIY
By5HkKMR8iBNyahPgpbJEHMQWxR3fVW5iO5497yLOCi1D/yTl+kx1as/e5rwpdzyR1znRbSPNzJH
QV4liaM3hJUSGCCrjej23bmngI2uEdVpYDphYzVAC2xNNPfsICFwlChHuFjh5jmM6wSes+saI5tW
F1y7OF4HvOKOx4LouFaFpe8kgWXgwWJpTGujDNFe0xS3BVCoX4VBttEaT5Jw6dxIQXewOYlBCqh/
nFffXpDaGXMK54em9Lu5quTFJ1WHqDjbpf+Kf/psXlYYrB8hkKaR0v+CC+PEmWmuebKa44YHqCv5
MCywnM7whIRaX83UmcHA7N/aKCqzehmKcVYLj4X+36bfgA3WLq2/zcGABPGi/uEBhifol9Ogw7b5
fB19X/oHZPSLTLn5LkdZL1dR+wW+Jl9uHPJVmQ+DGPTXrW7dQDX3tQ3UK7Jd1HzeY1CCDRGqOchN
M8YTTZ+a60uA35s/8vLj+0ob9BMSr6ppdqMrcJcp9juB4a9Y5ulIDiiLMbmKRaIRALMAnKQyox6Q
6fH/s0f3QjWqhfjcMibKmg8v3XsBeiTkT8YHli8e1q2H9Ri5on7L+KJQhWysTySh0M3WhHfDrS+z
Hfse8NBzwWwXI5V9RItQ1eYoPMFkySTNyK0zmMbBEZGPeb6iE5hEP2Fcfwj0mILKP3wnnFtSl1yq
z2ZwsW6RComEGaESaXB+2gAI/fyXeLCAc8HckEwpu/gdcQ+Z5zwBww3B+fKYX4UyrUnwF4zGSFP5
TiSXwX8ViGXdskGz7DLYNHGzS8rMOm3doYQgE7zlmzqmU5S/XBsmo5RrvoP2lb+/rGQX5S03w2/V
bfX3JRS7Jwha6Gw8uDeU2NSW3lHfa1yi135L/lX/HFWBmN1IRDOI29uM/pTXefNubE0WxT+PgLfy
cx3vVOSQgCcUQ/sz8u+VBkJHUvCU0O20exTfoj/06IbWy5zipdjkBkVBnwDBSdU2vbbU25geWKCQ
upyDlxyuIYlO2f38BUkLCRvTRHCMVDazlYMVbm974T6/2mw05hxW5KXvkm2K688OQOhY9ZWdX5pL
52mQA36vvtp3xzPUVPIcX9S+MQ5BSwVqzFQ8XiFTgYKdLc3Nuej1U6TgYsu5/TLozL4en5XqHK+N
w8IA0jsORgTO7ZFN6/srn7Morx9wB5UJv9UCnhvt+rscf+fXpwxSeo4DiogaBwV+QJ+XiF4jdyeC
HvytVL2JjnpuECFOvSjowfdvCexEVkXNRZSwh8cWvKkKJrdaVfYJdSVP75StnzIkPU0sMSoY8trw
Dj8cqZB4Bk/ZO9zKCGPxCDhI5c83+Fh7STUm4CPzgmWISCsX9+V8mmmYeYc0QULBVdaPjFKyWY5x
h2HmoX2Og0RetxpOMFlT7f5BZMzBQFOR8628/pZ4LYR0HJFYtReJ27Bz5n4SVw2ihFpS4OuT3k19
lABM6yNvEiMQ1JP3ETGhCoDntSkGqg7uRcX+809VrU/xL9zTD/bVy4NGZllu6euedS1aGZfR81x1
AVxbvemvf5rmOQEqNUqqkbx5YoY0Ln7yfQpjupkEjoJn8BTuRegXuyAn3vqouxo+f4eFU4E9Y4AL
/ongB5bwzG/F6mI15eH2khCGP4GA70/m2ANssIgxjrf6bW1IfyOKU525EUuyOKT+j7I6BaZt5/zb
HrAb7IPESKg1GTYUMEx+HiDbZXz9lkoyA4gHWxdzIpJT5GSmrHvTgC5hflcz621QjVt07B6J/f3f
TPJmaakcA2AbynFOIm1A4Ip3RD0VQFGt0VOUlPd90yAT96Q9sdK9nAUxg07zqctoAkRqroOBT57Q
5CdtF8QPq9uaLhhko3eNIWiC5hR/t2mJNvgkJHuh7g0+ah7V32NTXZyIbW34uZCzuA7GFGdXuWXw
CGxNAtDdw/fpuSTHIdxtv99M+UbuHGqxU8WJiQ2FJuBNPluviaph9VzWoZxiU1mD7K6PKcr4nnEr
+677CjHT+EbSqjdKYmgSqAxLsySj4vzh6ZB15EVEbOzyqK1ivY4FRfawqIk1pD5hKwlVOqCHyKgS
9DT8kVXJ2dikteh/dg+1XmZVs7VR0R2fFfjNp2iDF1eEMiRStjyjN6iRSVG9Tud7FUKpPhwjoKnK
tgE1gu+wefuejphfF07X+SzM9Jnu24zoiUOWC1d6e8ANAcwXbBP1vX4Ixh0as3WjvWzGOp5xkKCj
R88eyLaclb2HzJrigfAaoMrAfdzsqgBYrPOZt22NUzBJ68AGZoExiFYbQ6E91Q+F+HD/CfBktey8
dw304ZFqQgvY92PIK3r5kKGzdJRxSzIE30O69XWjMh0664pcnyN2wU40FJLADv2muazoWJoSY6RX
QlHPKxCINjqvSPGDo21ZylLUhnFyXmCWANLbUvgD4FStgovD3O2tdlD6K3fSu3boCh7kzo6bWlUN
FRN2d7CsfGtHvZG0xrp4G4U9rBR5MnEX0/4w0VJuN9SHHidLXsYybl4ztA9dIOzfeQ0Gl+u4jQh6
PO6VQ5T+M+LtN+JIOxDdGttWtVgnvITePSCv7fFWJq7OZh+3YT5sIcWpQXPVj/1xK9+OBJkiuHrm
O84vsFu9k6vTqOGrsgITv+bfP3wVX9DbOMGcy6CYWkhfmHq/Gy6Ulm1zgjD/eL24LiVz6SWYyquH
Bb5D9XtAw6jD2/XLQ59Ll2/l4LJ4fj0mObiI5VQYtXlkDdywQ8x+wjgFztm3Srz5MblOGXUXKgJA
lMme/m6YIUmqnwHG202FnqSkNW+33LUNEXuUNzilRHO+DSuQlhbj+BbAZMb9iEezb+daX03eIssK
jdsICBd+M/dl4MPzZ13q1zpbBHFsWB9sleTLXdCYPB4zPN+yeBYD+Nue/zPC12iRkxtgyCiHR1q0
HZkHmChuBGxlniHkItgTlkuDAHSA65gsQzI87kQmVa1i2nLDPYT8azKcqbDJzta6ojwoIuKOUQWl
SXAjUE6J0jc5VgmjANgznBO0ZxejQYZK7ArR/68AkrbfFJqkXvtP/6AuN9QBYLG2bO8Ij6PLnk5E
cDLwBQBf8cmteZ8qsu8scN8C4A7cS97TQPZBU+ESsSmjEnsyiWzJqp1rYsJwVNlVR5k3zujFPSVE
TiCzU6vT9oXCGepqh40RScLw16hkT6eQdwPOSL1ycRj9UNiVlxQ+vTu7jl7jeMKg/lwQvDmMjZtt
FEuImzM1YEY8vkQpAzZ5TeeYhABNJE1+wR+0uAYqQrqumHTInrRhCvfkg3ESzWZaq2zudg3MrUFJ
jzd74kNi1/CYvpT7yQwuuQG2VGbwPxyGClBsKL0Sl0xnJUHW3v9ML4j7wlQYXlYlQI51vSMlzdcM
iUbobJH/c6DgLEwg/7BllObbe4SJZuq1OeC3g8OOTeZaA3XUyLpMwQFT6eeQM2EAmWgL3WO0dNud
VTU9sdy0abSODCbciL/DZoDrdRozuVdovZgiyaFCOgUqxRUhAvpeQZFRS9B0NkL+nlitH2004Uyf
XZ/CpZ7cNbri40rbRmCZTdykXNQwepUT/gs+8ZD1bEn41ViZ5GzFeBr11x/xU20VRz7youCmAtGY
d5eBRCtgk0+/GvNRGX6qNAJqE3ol5HVKX0MMU4ApH58hmeGRcEK1ztf+QBDZS9agHVUTXpabnAsY
dxWcI7XExDT/XZhzuX4O8etopmcXl8nhHeW9SSQGeXXuJfqwwETn/D6mEuYyW4AUuYU6UvEnV8pB
ZmZjDbAaAu5OhkDE2JMbwWUR7ldT/UrgdiyhdxFW231N0okHQJaNIiYQX+RF3wvVv0HpWK31cREo
U8Ju/Gyf5LR+PInpXupR3Ko4lvIDdk3dmbHlXZ0NxGXnJxGlVjRoLqVUX7RGL+BsrbZ0B3+yACMU
GFU3aWHQLFfIaaRCm5s48hhkJ3rpbqIDLr0bvrD2ubvqATV6iWm5x9pcE8MuYntxUmLu5iKHbsSl
72m3V4tdmToZaybaPT2gS9Rc0PsTHEsIFy0Kr4cUkxpf3SuiDhNlj+KK/UE2uo2SQip6KABprPxW
ddJM3Dk1z8JLz1EuoGi28dfPCcnuMDEJ9JgFvqwQp1IJ/vB7UjQRjNgQxODA/UNc9hQdBuy0iACU
+gv0xd7ztgmZS0OECzDwWqcmOPosKnoVnGLlYPn8EkjB/0uc0Wlfdb1ZL8tLs9z/R1fXhoHwiFS7
hx7yR3zRAAcdj9WQeuoGVYbdcsRaQb5bg8pWiBK1y8okhnLndeKpMpyggESE4sXiW4CckGgEu+LC
QgUnyyU2QiLYlWUCoLLU78tREgkdbN/FttZwTP/9A2qbRkOVNQ/xjc2vNVpvYihJqxfk42fJJkSC
w+4uwkXKFl0o6weY2TX3w34BrveBp3pzsXvVVThti2aAUw9SteElCSQvlPNRafLaTzNRIn66rgDv
MhRv6leLEAUjM3Ym8H9D08TnyShi1F4mK/Qaq6q5YpNtJ3+/Cjla6NsICDwRxWgL2eZDOBsB8T0b
gnNnKvNfkSTb2lNgSIF6s/s5HNE2WLv1QEMt+eQyR3o2zhvt/aQoMvKMOnlvBoNNgzejeUu3LQXk
td1MCsfW3Eb9/6qbuQYB6NuLY+5LYaQUXAXOEmLNxkO6TogBmUzKAS6+CeYZWubXbhBza6c/N65N
g3j3QQlpEcirkbr/NLqKL+607Hi9P4yuazm0uA3ZercSZmDk1t+x/vTTJdQTaDE4HC2tadgvpeKN
AdvkbXN/i25ofY9dDkihbnkRevsFn3zEdF0KRVy4l8k1lE2MmHi4UTly8AgLU9+gxIyhJh+9FFD2
dAGjO2bP0VJ/oJ2kF7GFzAPWkKVRDVcw/iHnXh/0Cgo9MXu7wer6TQu+QJ2h1d1esjgIBEHLVuk1
7pG93eZoDmuQMGReU/jNuufav15zSrgyHZ2gbmTEkxEXkvb8qxiw1KBc6QYUN4h63GGgRswOC8qq
fULPBHE9YWXzYEC1LoDsohbQIOetilHHvHY+lmQMMxK41zapVCmw+H1ztKRqkrnO+U+VQ4k4EcHT
nGYP1/jXhd+9nlZO24Zz+cNYBcmEx1k3TKRrMa4Sea7muoR8DRAjUuL3Flzc8T7XrsXlNJL1HltN
zJgHyL2FzvLtA+D2thXpVDtpxocvtdB9maS/UX8LJ6So8ri2kxx7MECobwj3OHKYfSu0VXXl8Lkd
iGmPMrr45IqpeS2ErNNQz7y8GvSMTUJtelWqhowfZwtzcHLyMhgil9prdOIuyWZcIS1dAx+64DDo
P+1OagtQOdXzYPnZa1UHh+33yqGRuSBCAXCI2n+gOxj0IcvBjVPtYTwhACxunKa8zDe5iLzAl57I
w7+dzGSS/olIbdt1s9tQOQrkO+1W8FguKOXCWsc8j62fqrM5TlQkn8E8V0EGprDYPFJnlgEAZ9Bi
8tKKxD2m271PIt2enGF4FhWDg4mYGU+Fm38VITjCYS1CASXjWEvUBpjua72tjQg3BOgB3i8iOJGV
appRFIBb6fRV7Y2UcT9emPO1IVXPqqndQdbWHCv4XlhlaAHwwR3rEh/fA/8Yl1iUMRSgCoHAk+c2
jBN7K3fmrDthItij9D+ascqsksK0nVBvsWjO/+HRYGjlzYvjEu7q32thInZNrAn8STHlqU0p5viY
SpzUOJBYBE8YcDPd6MtAMw2cdByCHQ4q7nV6wH9wFxlJYpC643P5HPHWYoJpI1+TQNZMrBBj3nRw
6mDddUS9F7Bw+l8NpMKAw80qvFquXlM12f/ylK/BefGKSIeHvJA6gCZd8SbcrJ4q/KDr9kyDfHoX
NMCSBDQtenS8+mYU88uLwjydllUmPRnCdD9SfPkErei6UDIxnyslP+RAAqDN37IKp5pZhpkfozaC
/MsGrbjebAJ2G+HpiNrenVJMf+a7plvVguZR1Lv+adCHr/axsEaAEyEMOFmggJLwclL711oaK0fO
ipedI0+dXLyB5W4pGZW+9tkgvo49fJzt0iupQBbt3D29XYUe5FIZTdGXmk91hJmvlAkKngxvup+W
AXqv4BilNmkxECfOK/7rP4smn7Upth6HIlML7mfRWEBStgOdpgbyTKl0Q5lbGbGLA/SJ1cF8ZaRK
6BUqfdc129pGGaxAUtoLravo0TZ+HlPV2WFYvzUX6J4oNY/7GHKAHE/hJxPdYluW8eXMPe7uaah0
TcJUYS//nPNbcUE3IT+ZXHv4cFcQ2JohZRCsBVSvID0fOlYlRSqBYrVA/EeOeOhsMdFBeqYqZZek
rZqOAViVlsPkZCzyzRaem4FUGogOknKAdtascwwOU009U7szcnZaEGDLYVbkOVzUbRfIW76X76yV
3+UDQf4pzdmxjxf9dvXqPo8qr9dQUDcCCDXEyBcy0VN7DkS6jG39p0ibCCoLEitTxaZaCbu+lALp
xrSNpsrLFQ22ERqhLwZu/4fEYT7wLFN6PqdobnmslwpJ2vTnSqiQ+8HlzQ/mxkCz3izSLaRPzH/R
EGI1YmMIuHahQojnQWVtFHGcGZ5GH6L5XqbQzLNVZkGBY46prMJQQWsKsB9QBIAivm6/kMUYbqFX
+vsp3HFm+IHkvQ8URXdoCbPKU5L4y0mOoDf8IpNyd7GOzw4YZheZ3RVYiG5pL4j6zCQINcSlfJll
1tmHth3kfZrZ5ZdS0cZlwsvK7/3R4Re2j4Dic1t/oA32dBPqI3yUPcz3dhvp2loAVKBpeOXb3RFd
lBgl0J0mzmQ4eb60VgISs6SP0WqvQJ8htoHQf98x77Yzt8uioAzXUYs3xl1DRlPVy/ZoWksavbfm
rbkn2xEquxWY9PFfQnx+otrDi37DBGEsFhfolpkK/rGNepDUKQNY5s1eSpiXmBI1YMGLEgJ6rCsb
khBcX1K8nFPWGwoaompLRRPqGQpw2oO6WXwIlhCmkArM9pcphqFoCkdImnDmQB0Ff3YikX+i5u5d
Wy71pv9R/3KrvuzrRIBgJ7hoTObW2+mN53kIk4cfoLBT3TG3V7NmXpQyNs07zkqkIOZWFN/xe5gN
T2zmAQu9slHddohjDnyRaaJm+TvmN3HDU+qDh8Z/4p6K0WY4eISsXUakSGfPmzvbKjfGV+vN3lG9
NstwRhG1ttONtJ1GswcZI/dzS5j8djnNYqTgIke31usr2x1gslV4LGAAaWQI/aGFEhMLsiGBmYgz
x+4VFGGFh46PQf+h91u5UqOQ+Jnql4yGb6oa5x4wnY7Ml1PHgIruUUDCtcS/Z9yWjVtpnK10BJj2
08MpJbfWGurPgY23yl6CU9idXr2tWYeU8SR8k0cyg8jb7ML20e+S8RK/PyP+XivDvZXQDTOotxKC
y2fpx1yETI3cO35Cpo8YGNPW30MTnkatsvir6dJW5saNjNaFJEsodFprrkaM/3QBAkRZfpOve+PO
BJqA09f4SFspmwt8gjlBxTP83kjZN4MFhnIYVGjDkiiG7UpMFzLWy5Gctr1tn1jvVw4c9SL9tvUb
o8hi/DNrTrHQiOKn9KJAu+xxnF5I1w/OH6KDq5CI6MzYz4hl/VXhuaj6TuMuUxRCba7tVqm7tMSg
51COTIdxEDY6fdXDzQvYwwYjvQlGcr0Zu7NPSYfgMIgA9LeBeE3KqgEAArYYwJy+jQvxDgc8phsD
QTtpnY4RfqrH20gFK0e/g+x9zGilxDduabuL8UV4iYu8dftj1h83V4Mvs+bO51lQsYE7do6VnLBL
hnUtmrpQu/Glw26OOBpJ3+GOJlcJSE/ZgpyQ5IhbiR32iozM7L7r3tX7mFxcvbm7TuveBcN7c71U
uSKkANnVc6K5aEMBvx+jDhJPculGPwso1OJvsyq89uI98hvH9h4ld1lBlevtIEnedptc/BdsBPCU
EbnAXek0W6QQtB1Tkbuf/02blCsZ4ikD4e4hNnW7MI9vhYeLygD3q4rTnFr790y474kVucKJNTy4
E8D32Ufau8M04hyupAe93F1yCgiA3MlKGVbO117wpM22qKj5JnQtQ9Hdh7OMe6cHB/AqbfQcebBW
JWvQn9rL1K/c/KTsRFZyRsIk7RqmtjmFRUFS9mpsKq8It4ZizXSdltW4pNhFoFBhCFozY0E7REUE
QKkD3I8FS6ceU9xQ8yRdWDLfBk3jPnzu+SnKCHf2MYca8ZI0cS2ez0cvJZ5n+Qrrh/QICzmXk5vS
NHk5mWWFCzyuqxPxI0oJmTe5o4RmS46qaKl7qGzavKZqFQebwLGVupK6lBJ1hy2NGHdhBY7YLPEG
Uv8gZEbN9+MqthbYj+IiMzszk152wmH/2utYwZ5a04lqnz+Q2Urr3M7QC5yOByCYqpzihhVOPMIM
0Gd9PVeXjeX1BzfVHaCn6tyGibfSJWCwJUQ5xH0YpXoJgBpHTOyl6okOZtbYW2j+03SkMCswEo5S
ubEtLT+nro0BhSytcI9Jf9oVN1iTaJqVDmFMarXzmRD2nCQ5R0KuCCHwuWYhomSjRvSDVxj2TFGG
DGmPbb0Mm2dCvOh3vpoDjtgCNCKw6fssb9+ujquP4P/YnHns5to//C4KE+/clvupaIC2wE1jiW/F
4F2TRXAh/CCaEtDlu8EGWY5T4cyomoMrGRSZnKj5usNEMdHXZ+/2WYqA8K1DLznBYHiC3unr8yVh
9p67J0NiZ5NPyAQa/TPqiDJQ3+f9Wd5UQNB+iW3o2KyuWgov1EoZDJVbrvqqyUdCLwZ3SmGzrQ5j
MuRKZSVcN9EboRLoGqLSU5b5CbYTmasB5VX0dIyTytQYe5m8YAkUtBJvs5yYG+W5Kjq0lvrSn1UT
KEuPADP23wFvUJCuRpUKwgeXxdJWvD+WrFszVjmezCZnc8GabsyqDFh9/bRrTYIl9QjkY7VpmajL
OvuKrjO/tSWLKcxFP/H+p0AnN3X83PjGkgsrxJl++V9aO+JbkmBedL4yvMBvHGY2mztkIP2y/TzL
VKGdpSsWPhFeF05akXWNhsDhhmpevwBvtcQAxDMWetvDxdhxjuPOYWspI/5I1Q8jf5ELlXrmIV97
hYJ00Eukh7slr+yiXMckRnTO4QQ+XB/ROzU0KddzJ8nA2XpXR/jHYAlpP8pMlUrc32aEGxWkIW04
Nz73P+ghF6uXSJqIz96rOqWivCH5dUi7NT92JHw6RD3RkcxCVuuQIfbQz8K16J1aZ9BjnqoZ7t7U
U8M182fwQLQA6U3u0uwOaym+4REFv0F+PPr7r23VP3X31AtQcIZseSKtVDdAQBijXxHGmv8q4hN4
Z01QKDK2U/k33i11YtgYmU0/G8pOtNUPpGIFYYrpOET5D/YltSoEkxqki3SrJJUUyd7GQ+ZlpZsg
nukUaujXR/JyyA4mf3ygPaWIJKFAOxqvsbxRUof8RLGdoNGFB9MWiaBvPfqmvvS0lADu1ptrWcGh
KdIKZ1KYJOXUOlZ9QMteo9DnKdTLKGsvKSzEIQs9D8aCE1ro38mlqJODO122n5k6dBtMqeiuAB+5
GYKa4+iWeEeTLFCC68yxnzbrAzsmrNklU9uqHk1wBJaImAysKmI2ZNufT/FO6d57AhZg5Y2h+pou
qud8VqaBCNFsY+t9AFMMo7s13Mv4B2OwbUG9A8tGGGO1C8S6Y79+21gKj4U+PSv9mczUn5Z7D7TL
Fi1CVQXCH1L6qVqCvdQFaUZNZEr0ge5UGlJkaEK2mtqPeX6/4pNkXNuoY+aV5tsC678FQ301iJGD
nw2ZhHiJs5pWalc7LSKSdqZ7EAMR+c8GlF8UdLFsTUxVUwRjWWPjWLdXArbJLompIGdjQ5VmArWa
y+5s6S2G8o9oFfS+teEdO/detFNt2JnPEzJfVDBoe1xHH6oc5/I9PIjWw7KJUBt5x4TlzXih+u7K
ReLrcwhLZxIbZsx/KY4TS0DxL9LtmCJCdUe0/DfJIZHAYWtk1TftlVDtbBc/+4UONoTeHfQYvbex
ma+qq1GDt0mg/aQzXX2LmModlCRZNJ21Ydoc0MxxPFrY0iCOTnpQZi8OxgHgiSehR+a3J1p2zD3K
wNMLjb+hWlFEjUX1FSa7O4hhVjus7o9TyJ1Z27X6upP378Eh9/aM1d8YsiIOarydHAyCHS5P55HY
xacOhCM2HywbFmrpf88rsKy/tVLkRQYA8fPaJ8RovMX+Z2LWe9UN77GsAD9Oh67KrCobxXHTZ37N
aOEdejfRvF5EYLFwMIENK1Pu1/cEwM4UWJqtA3OCr9tEQ5XgYQwx06PPedaQhCA2OqCFn40wglZe
MHq9HN7aCHA1yqkkBVUDMmTXzGWZ+j6+YfR0du/l+OhdZDLbW39b0gQME5UMg9G8NWfXKVQEke7d
+JUvFebj3Sb6GcjK4qyXgkOwtsLk+u2QKHMjPNTa7eA80NBGqvvFXA3ikDI6TN0OS/1NIFoxSEjR
vBKp+1pOoG+yBBM6j2yShWZstmTvmTLSSQUoSdkIqJRe18QICn1I1KnWBJ/6RiaRIs1+iJpao/4t
yexEUjQFlLm6vLhWy4ao/67ylDR34nlyA7cn77MFU7D2OsYoLg4phbwiIw/teTbNquFJFyvv9H2b
QIuNVvnf9S/A81h6hu1HWtgRLjI9mivhtJoJfq39egOH0mwlY7jlSmHzYu3cK+NkgB+KePxKu8gM
oq7Hf2E+je3Y08UnKfNSqfR4TCAj8CLSw9o9qR+c26RG44UhmbhHvlz/bpB2FzbUz0DsBoMDaHV0
9aANVsVlWGao/GLO9YDr8WxLWi3soYZ9UKRQc30O8KZd4pkvwZF7PgMQkk0MW45j1zM+WVxgB7Ct
3hwl4G3NoHC+R2h5JMt/SYuLpmVjiuAUBYgASDGwRVVVxnfRCu8c6kyzzGmy7lq39InkmMXjfb9o
k+s0CjSOx1uDVbiipeuShfBUPEaJY8IyQiJ1IsuP3rRn3WK8TyBiLlCquClPentqv2l8MSoqhA04
or5byxE1RzfmVSQIhr7qLjO/TSYU/LGUf9vFiMqy7E6+n6y8MBV+6EF0GTUNyvDYBcRIJIPEXa08
qEIpHr7HK5zh31OHIx09hvJ/4g+qXs+anjpKWi/Fmw/4FmFFdLB2/AfyZ2cIVoSUqqWomUDWYnfU
CIcmgjTDhNCMpPiWj98NXlErpBVJh+rjO4RtxvpppxuaU0ruckE4s9cm+uLegNF+q3815znIIzQG
t61ro+ZAQJtIfndrtL9lAOpY8JM8nbSqNB+rs1qvi0qwal72ztVzFs07IGaRTJ8Lrd04Gq3JyFo1
PL2w7UL8G+2CgtUy3ma0hjhO+UmGAOxbCHNrk2LvS+AvuuMDqeRVrFFNaaB7EqE1lcYlFqKbcr/a
QwzXOEUQNj0KsTH1Yvt4qu6rbjKMRZ5gXwmmcM3bxZORrmfW+v8mF5MrjTDaA83FO1K4+Xk9fxtK
xQWoojPRZFa2ZyCrwdT0GpYCYux+5xYEUP0mq68/cnzqMd4CTE4x+nNGxXuCzA8C8fcISN1Z2FRi
5F3F2FgZzX16lQvbz1GkWOYABgexvqF3DuSiUXcVp7ytHF+D6BzcWpvMFwmx0RJL/7q6BYvzOicn
ROz8eXhzSWTKPYW9iwxHjgjhDqYHMjFxosptjQS3In7BR5PltrAMz8rf3iE5Tx33cwJcRCYtrVWF
XrNzFd+hvpJo7y0gq9quMJkKpIL0Ev0xvjkYco12sxVcVJOO7pwNdLt5ODahi78KArsFu7OSSTO+
tFVpSQuISzzYPig4R0bmDMKq+sJjMpFKEI3Qdy+Hf9zwkUyXclxmskzPHibAxhRRHFmvVTnUE6kB
qAcFUOvl7HbMmY9a6/wuNs5EshlOr86lTtugQo11u2eU0jiCXgQ6BcYzkfdGQAUNospDgj/bc8w4
C8RyAqpHMHdIXqUijD1tl4/gGyzmtkJbBIeYN7sIsfmHPerzD2GLFKn2ky/2lHGURV+JW5R7QhOq
dSvuHhihdUaoi+XN5mL6KxqbXCttVXpVvaC7AGq5VSL/Frxqcc7afCiOIwWkV9rikRBxFNcznhhM
ZtbUbwjW+QbI6ocDMsufpUJlfe3XJcO4O0xZDhYvKH8wKLCLECxreJwlvyClL9YjBRQNAkSDjmQH
A5GFcq356vRcuBJVi9vysQf1wMh1Cmh63cVxLZ84IcrhoSVwtkuxJtzptlxYZGPIajUaPXjz+8ub
MVzKOTiFy0dAAhJWBVyORs5650dQQb3wwva6qQlURwVQHauTs7efyuRKMHVExXueGO22MSkLu0JV
mknn6KGBJmHZH73KzY8YCO5nRCgjhMhzCMCajnI84PVFTvnKUmthGU3eJejOrQarB/HdHdIw3Ibl
SxQxJI3iqklOo5Mq6nQmgkTjumAvi1t5aOuLY+vGxxAXqPr6MZjDRr8Cqntb49XmQjGHZfLOlGNE
X2aLUFC+iZ745NtTfounc9aikk6O5GgBhChZwntfs56QvpOGagc7E5HGTM9jHI3ccIBCbk5Nz3tV
epZ1MIssSkttw957NhftwdMIJQlinrk0OISW+/E6H/Lqu5ds0UU6bFH5XSvq4659TZRmogk/ejdN
2v8K2sSW0rrWZ+kF7EPMOuAmO6PovdLz35m0EiUb8y/u8XVDoXsqLTzb699Z6EQpHZ+/3pECqndq
LqsIzQJJ/SAheHgTPHlsHOomYa8YH8XLPx5GlNzo0fSMJjyA7orGSXq5GyDlnIpm+oIyi+XBcRSX
UKj+qFVXUIMZ186Zm1Tk2C5uTB2MWB/34yoleHnFjIyMNjQX8kvCWb4kPsiu1GlPx/L6SvWJaPS7
ZeBFZFYeZ39dbtkXC1RH5XVF/DS12sicwXvTKch+IVvFqWpZ/mml+sUMcrNhV7dyPizEzr93ckPJ
Vctu0+LVZgWMAfYe22mHGi8nsssNricw1Z/4uzmo69k2keU7qRw0gyVNsHrzluebIvW6DSE3f5S5
ZTd1aammKtiu4Gl9EEK6OUAdxuWia2hjk+bLwd9dPPF4UAB9sXNrj25Y/e5fkGsSeHRxJVOIUaK1
00ZoSkE+K+gLfOEZAvWsQhtXgQu35meXG6T3+Fh4SIrBcEoIWXL8F7NapqNmeMYVsGlMmYIjd2HO
FIVxE0H6kVnZeHj6ivhDqeF7ng7xFuNVooTuVKYoIGCeGq7SUyhC3P4WK8TuAWtP3YEcEzg2tgfc
R6/z9ufySX4vuGyOWCqDBQmsuOxTprnF2ksyJzBhTWXVIpz+LqnlYSKiAqjwuzIAsYstVYMK3IWk
ULyGBtib+OuaediB3pfrjATgCFu3WBW/+z2lM7MCDv0ZWWe7iiBKN5YC7mFBBy72ka6tIKBia6g5
wMotklX74FG8f/Rgu9q13zu9lu9vsplUTBkr29nFdN8urQDtiOV7s5U9RTPba1OndoLOfwAPK1EB
GQGlwVKfVfiPoyXF47uNZlHC14jUKKyR/fgHrRgA31kyhA9j0id4FvHQKMtvG2ltvpYbtM1ZUOSq
EFVV4CoVSngxUgLe7RJMf57+MmIxoipyG4X+SARXwWiScYBfsgrLnoOaAT3b28nB74nm5uhdxwEP
tjiusRfjOARY7oClw6DxcxSBGNW1hk4OEq1x930wFnT9FVMOT7TJA7Vr+i4mv4iekMxZY8vI8doz
PkasVvla99NW2UbdAC8MqNd/BQVf5DcAH7v+AZtABfkGAclyvwpcnBKpf2LNrKJEK5LpPpJEX2GB
ATmRDMrGXzd+HBnQE1ZkpO45mhYZuaItuQHg0t5T5Y3875Ofk56lZgZUozXarPWoC2k6RYPeRKwX
IFShID+xLjA/7TFxiNmpd+phGh3+BWehHZngGsozA3vY6XwjxwH2nAU1i8qR/EV6APLiwmbHr3U1
FoQ0wDvzqL9LZkLwB5OrdkAnNmHgsNYmNk+Q7tf6URHmOjUCCR54E04EZaEowIqHgTnjYBwmZx7N
zeBUvDOq7ykGTD0Gag1GARHgxAShrgWVh+fqW7T93QRqJej8SLVzFkhNlLrrXWbe6sgTBn4KIz2T
ZqplACjyAZ6WP+5xT+vhJhg06DuvnuwvnJQFl9G1NotN/NX76ija2B/+ANEQTW9stz4HYHsDmCCj
2jl1p/DD10HWW/tBy/F9pKVOM4QnEnDnyLKeHrrwWOrZmV9rPRcNekHJw6fetIRawMmDp32MXLKa
oOUsfAYvE4P4GL1gsrwknyUszjXr0j/F8Op6Yz0fHo/rOHUnUHpdImVIn2Bo9r6pE8kZQ2QQV7tA
Kt84cxXgTZq3pwEeYRmUM06Zqx6MCyTE4awWcZ3dNpPd/Vy+t7AMbtbzSa9b08DqapV6jNuTtAF+
ieppqcsVS9Bo/PZVQh97YW6sZukdQWZ5njqrlT9WDU1QfzC4QsULWnMRw3SEAF0IYBap6Siof2eJ
SS85Z0zsd8hHnNM7LULXWZXEPJjSPZZMifkQXHdOLhCFAt6GN31rCily8wnDv6RbGJYg6UQZUAdP
y9//R+TcnVW8r/PCQ+pld5s9r6WSItBWL36tiM482OdiH/UuKiijgJ6liIvkA9H0+1QQoicSwrJc
DF+Kzq0Ii89VdkdKdM09j57TQPqjFrsVhpn8hFCjKgxp/cd+z1IpcnjWfPS0/FfiVVl4vv5ekQud
bYZ77MoNOCJy8U5YquWc4n14SJG1IvQo8PlHyPO8l6snlgdk6cLFLayBo9YwewgyZ+2opBvQKHLz
+vW+u9gtWNnVopGavDNDH22AUzgQj+PYaPPf9JpDKqpNbVcyzcNv0b61OUAuBn0k6aEFVSqKDnuL
1hYgO3WweraeHkMSzRxAt2Gc8itF2IlVmvjuhPGXwGELgjdP+4TtYuBqavQQgN1zk8cwkd4vzK9d
JPxJjOImAL4lbWYIFLzzoWe6y/ve2NHKmgY7/rVFAQiW4ubEOpidlOR2zskr3erTcgR5l7lmmf0l
sRfqjL1+zi39Ulaoxpv6vX+Wr7nGiBr01R5/o7atszCO09rAHa9auglLqfduQzNmGPuJDlvXvW/r
2hyUcj/PSYiMJRvu1qLQBi9cj40B57CVDqe4fBsS4he9dcRCpcCEr4g9FZwGApG2DtnF3K1rUg4P
qRBTYWPgJuAedJjH/mxxrai0Tb3b9ru+PIg2iuOgVwj/Zc8PHBf0v1VaB2WqQa/VOo5ggr/ICr+E
ObblhKRjHQxxUuwxaDTVWoOCVwFQkKaJWrz63W1SogHm0AwT6a4iCeRZ+KhIpke2EvBsTFpP034R
KKosxfgI7NnUiKkAx/G8vDJJFNLlZcQPrOEgfwdtxCZgV7egY1S+tGs4bLJXRROuxlEDyYQ/XgvH
mdFOcamZgfQEpHyDnDCuzS7NRg3OLi1dtSmRzFrV+j2r/jR8TrDdwmEX7QVZnuwsDsRUOv609pLv
JIt/fHp7jEC5epdYJxaKh5dbIfL/EkvC0BTLBUtDcFXwaH0a3g+MpGLYdNJaUqn/E1gs45wvTNN+
RJ637ymsw5TrE45zaYNGHrqtNCq1tOznOXaCQ7ZqTMDJhh4V3yg1tQzBZHCyIgnr6u7Qhk+6mDGn
YmQeK+4LE+nx5HKF/Xszaj0pCC4uPEoSlzXSFOc+NyQaC+cVMyrfSfSB72wFcmc4X70AydeWJMeK
l9ekcnVWKSy2ijgQN73Mk26MQDRivxL89r1IJUDNqqhLQoQqlb4gku5fuTXqp66xopRhD5R/NUYg
P3qd32xk94dJKX06cfbhdg7hGLr+NFvSTHFOgTfz+gdFxz8f9xSwC0Da6i5wGm9e5kirJpPwmNEq
R77pdFSPg2eQvQsEF/XqMuZrqUO/WVCLmiD9s7QScz9jaFWQo3GaJCfyAioG5XntkAAUrFVd/CbJ
n/fdNitWTn6FMmQDXEmorexEb1YqqzdeRqRSg/eUv6xmy5o5AxWdn5F9uwhl0kqzdOl1jge/ZAwz
rnuqDNKwlMF3i5Uho00bdzWOJfknahBpu5FxPznyRaVY8pGFJxqfJSaG3woo3xtE1JsKkxGWZC8O
CBbgbjF2y+BRKs3Mgt8f4iGCxkfukHTlf9JFi5KFgSZbX0+1gHEED4CQ1ibluf6DyVJ+W1N8D9v6
LTfsvXTVlkLn7X8KaWZlaYpqM/LK0qTD2LMsYVf9z89o8Hdh0g5o4RysojnaLivMlCq0mYWFmZoG
Th8G8tJq5YiRQX05H7Mr0EjqzhmHzRWKT3RjNcpVRj746iE6NDrlCHxc+B88mrMwME/IXAEmFDJx
rvIlEJ0kM6CkjfriSSTvn+9c4nhnoEL8rscss+IKOqSUd1VVqIGePOEkP/9l9LFbIQ9AIos1thBx
zMj/UcyOYc6ItImhsTF0/smYXUyVaQgduKP+7VChp0dhYJrf7Uo49eRUsVzx/6apB281pG+sYX/I
sLcR3M6y3qSOWC/YXeXtv2MqAlaZeyfuOvuKvF2f4dAjFpAnnRaHoULFlm2KK15UIX72cKUhaDKZ
R5fmhOY5v4xkGiY6nuRiUvsjB0sWSXa+AfGuTXz7MxY0+cC8OjauX34LN5CoVIbF3r+uIklwmj+b
H4LKc7/EpmbSSMVybNpS5xciXsWAEypCSNe0+/8726kRsWo+FtNRz8ZnNZnMUj5xFmBPHtMRUUxr
hnKoMfxVVr2+0m0KMgiZnEUfJsRnVGkofV1qXoyyT6nUFQXtwKIRaK8UA4PQhu7b4RxIhsehpbN+
KUpObAcSjnft5cqM4FoD3ASND7L7z9LsTSeyNo5GdH08ivtVkUp3A5O9WyNc1xr5qOMd+QDkaotD
D1SJZ0PV0n7UpowDY8HtcY9e8OtWxpIppsEL8b7KDJXKCMFv5fFvhR55nSOy4XxrJeVvDSfPgQ8u
lBCrZ8LnBUoY5DYGyLpYqXPt3SaFj0bvCfcqiQ6TzVWzue5fuaiF7hlgW1oTXmFnlDsqe01rE70G
KceyvZxFYb5TGSuIcQSPTRRBteV1UZ+2F2VphYDuUxS0BYm8qvrV67MV+7fM4jl317Vi1gxvk3hs
8uhqLNDz46VIxGi7lJ+kliX5nYYbeiJHDPZCOrXxmq5bByHqjlzKqCeIFxigZJg92+o69CNWc5Eb
8KeMewuCQs5TL1T1QZvb1ni39FXumnD2pvP0wpdGvwUR6SwUyIVAHA88kRKRAZJX4oHQB4ydSPac
/YGxZ0pZUHZTDf0re7D7x0LK3aysF2ikG9kwO0RMYmAnpbpeg4YT+PSl8iSLiIqadaUoh27zYBjJ
RiIUN4PeVUgXwMdtG6Mw6suK/fVQqZqJ6y22AShjRRiQFd2hXUsm0OThxjBzqFBJhMH/TJA6dfqC
+h0l2dtsAdkb7ovVGKxEhXwCg88jjLmFUvwbbNknyO+nIXzi86rxmJTOdqI+s6ZbJ77GgkZIVYmu
5x8IPMviOSb39z1GmQEbCGRhR45/ZSNOHKBcRYg8m6p+rNiLSX1ckg2Fh8cXwAl2e6J7LHy6muVZ
unxQVg1k8Qj+3YeB4rZum+3M+L3KFzXzxSuTLpAdmhbZK3uTOi26hbVhehARMrwT1l5JMHaF+kdm
pXLIqiJmZ+6l2RR5H1igOafi7zqtgRyYdQ1nLHZSoLaPS839/0n6Den8TKjjaUWARy64XLnCuSpd
LOibnXuOuDws/HTr1rlkdvF/967H9UPVuUz7Jfvy4FyhxLhZGcotUa9DugClc1dExHkSM4wMYU4o
QuGGbBNpUtaPbP2+eABFRIljAomyXLA6GzJFA7v7ezRPC0cwCtKH1Np774TUt097Uc4Vw0BzHNhn
x9I/SqIW8KRg99jVMNjdc0gEZRIuoOcw1D+SRzcuo7z070nVg4MBZ3Fww0UE7qHn4RIswOT0pSp8
hU8Vm06XQLpL3WtD/a0elwwClR5oNyXoOUDICtPEU1kmM0QVu2Hj/SUh4jlRzjOFlbB5HM+LLkm6
Hy9MfeOSj3pCGloZQ9TrvE6LnE7r+jZUox94DjjIwI/R1xKY3ay9IIDr0BKeE9kzonHm173rBepu
KSoYm1p01VOH8Xwb0+IkXZUvwb2JD9hS/YKSmWkivYeISOS8UYgkn3UuMENFnAuoQhxNoyMST2Hh
VsHQJXomtVPaax9VdquDCi1NtlBLb18IJOcC3479S3yeL2ro7eC6mNO71eaAADexhUaaRgkefshj
hG/wkWDeCrUx9enAGj5iRUE+M6G/G2nstAVoWzCrfKUHm0hmoxmgFSuJ2GlMkmRKkkZDJHMTTxSd
aASLQFz02CpB4ofeCdsUZQKRz1JJD3TUZ9ytgkBh/PAUcPbipu9fyN/SrkVu0h9SPoxvM9tu4euG
83NUPeLne9/M08SAHEZRYPjG81liRd/wkTX+AR+fOV95wE08WHKssl62MnvbzNb5hePHiMkpIy/E
jGZJImrlIS8zxiwcPP+Uj60rf3q3OGvuv4gQ1LR/XRQjvFwz3fpKAXAgoGwJu2NUfJ5Eb93dgRFA
8talfLdwQKplYvUuSPwVBldfxJiAdDrqqc64JmmNY/8e8XGB+Fgg2OyDctKh3TMDfuttYHPS86tG
wacIK15Ao3V8cpIPb6a76UQGVK+88czHZ1UzLySR+pcIHeJWSJm31412Lu4dtoDGGQ7KLQ9Lo1iZ
7VEmAB5+e1yBJlCbD4Zahf62rQoBXK+UNFRM+X178RU4GIDD5GYR7iHWRhQcQ2Nsw6ZWpB3XcXKo
tL2B+XYP9ZNE4EgZe3j2D9KrDI45N44QTgqTvroDWZKxaDX9RK2ECJC97UZ7nY9WqeOW3gevenKS
yTr5lahF4IejXkJlOMuGM6cCnt0H9JtObgRix8AwpoGZmzRIYEosxGJCnj17kthrZjleo4JyW0wj
MVFiRRpHbENjEOWNjebCgCw0mxoNgiWGz2SzEQS031a6mc4+nmNHWmXyxXBsrYv0OnO0LpegmMWz
kUlhjm+q+sxPG3Wr+o53DRziJh7VBu4KBeMn2oTLwGxYvF3V7bHfxxe44sYYIyosVZJtzvWnKy+Y
bK4FsXXRM8XebQ7PyODZLxomT7jX84iMoKD3Nm28z8655pV05jYVj8Wd+6LpuKh90iTxm522t2WS
l02rN/YvRWTVE8E+LH2bs+pU05jH562cVj30X7DFC7V2mstFfNc6tEuy8tgpPaJ/fRmSYSMvUwEA
qsfzJEtSF7BWKyGMSIWFkJgRw66wnP7DWfCJIJD2SxVsC/w/o3nwZ8cxx9idUuXLrKYJNF7RpVex
pVn1e7KH8odXj/4CiRk2PLXiB+q11UoT3VBBk2Pq35+CSIcuN8+MFvTOVZvUshrXvddXPy+IPlM+
mrnPiySMtNGxKIvx1mnyQgeZ0IqUElnWKeLLbyQ+OBQKeZQV/s+8tcW1kuOwbIOWLpSSE8W2Q2Ba
XevLoRSHYnrQ/WWaTp23ykKjBA6m0GfAmCL5g6av8Vs3/EGxOayrxueq+St0w7LdFBR4TQjsp/57
XE+8HYjsM6BbbFHxQL4WRSLJCEc4oehE7Rzg5WzJ2/k00caKKa3nnAgiGhUXYaix/1p7pXkF71zs
hj4vmrfEKoR5fhPltxYBT9BkUdrXIyB3i++dk4ZZf1LRdlyI3joKLHIJgsmm2tv9TxQ3neAtP9cB
zg+JHRiJAohZ8vP/lKCQrOpQe1vo2BWVHf2vHb4dR/ZK6RvNgUy8ASC34lCH9W0/u8hyC18JurHe
nSAYSQBmpxko2Dcl/E2W+clsNhA/woMEwLkHeEjvKvF4y74vlpEesEOJejBFofoM1URazJqKv2eW
YoXRQNOwqioRwFrM1Er7WrePCmnoRXnsVIT3WcXYLaUXS9gjZk0AWHn/1q1NyRrRnx44JytA6ZA5
z8Cg4ZudrwgPK/R4764p3/YQW0Y/FE7YE85ue007p2GOGZWqHpUM4NgRJroAVAmrB15PtFfbHAX8
YHtbmWCPCH+oY1J+f6nQ+ltRMvzFHnu2lBqer2OHpFZDUvBOBYHmpRjnJYSaCHTa+HNc/9StJLsS
ZufYQI1nIWEdiEm9evsm3b72YCGID5XMshuEfgRLfwTWOPELbIoAkwrZJIQsgVLSwifE2nOu2iIR
n2Kvp76iGUC874QNEr2lrTeF/IBEr3zg+D4UnmGKI1xY23i0azWAoSgJfmOUf+Wc5EXCO/Kxi6LD
mWk/fLA6gytsVlPw3Xa2SlQbsfNOOH6ivwOY9BfR7p/TF5Enux8CFridP6J0OMv86TSGSe5JRpna
zqvIlupFraZ5gblPs1TdpzEdTdlTAwRnXwy7lTa+Q9hztrJqsqVcOhd4uH0SGRXh4aVvWHwxFpxv
z+oKJSD+AC4vq2vhPl+MKoFhBvbgRO6HVLTATC9CUox/bp67vijmOWaL8r5aN7XyPn+vvVfZNSi4
wnzPdOsKsXF3iVpebhZiesnAfWZH6yRCjc5ew+UlSlLsyAdvs62v8tK9ycXvr5jaICZcAHwLF3L4
9smDK5mxMEBu7kRTB0aFc+es2egbD773kX3Kv/gvdqRx3FP2rlo+W71Igf1Xe1r0hPiF92Fn8opM
d59dJ56Gh4tT5qSlwXc1DsvJLU+wBEEkmnYLwWZZfEwnOP35OlTxx30grc8uubWwP6dxE4RQr1cZ
S64zyty0U6/I0t11Xo9Za1bAqPufr83295x0p5q2diV8WRs5iY/GDDSvJQrEysie9h3qFUKmZicG
p+eN2euv4/3aOQGj6fAVCEM/Sie+PvFXWaqAVGo95/qaBDA9tfIEOLw2/pdV0QAXVdghrFUnhXlB
bb66b6uy6jvR2P8PX2k5E6T6tBJH/eZBlT5+Tpw5RFgA6ihva2zdZ8a42H3FkvbZd/7eDvLtEC0Z
F97npbtR3THOG/EV4cebLgpIzdhPpJL+rpYvt9kQhZ374A+n4KE/JueUwHphP0812uEWBgQIbMum
pH4MSwk1y0kD0JZRfAi8hRHgbkBQnzmu+kNzJDEvhY3OFYqofcrTbJu/YIh7dHYudeuloH+hnZ66
j9LSOFkysZivJPZCzZA1W9aFDfv8uVSyRPVYxJK8zUm1NgKBN/2JwqvlJ3Zmn3fEECFzZOcJ86o3
WR8gpfIWbwq4fsVnJg6o9Gkk9iNjyAQqNTjcYgtK0Mec6VP2pWvt0RaxogkG0EdEeWEwPUL9VbIB
srTbjci0fvEXpp/UAq29hdkTnJ8NBi4Ss/xkA3ScjRUurO0qeFWSXrUivmK1t4AoIrKGqrCZMHx+
lIvzQuSnOQAlMLLRI2lIQK29PGwHar6ssCusaHyV4aJ+rENBDdXb/bbi+2VR+DpmGql0AzxxmT14
J3PqrObLhkaO1bBgDaGv2XaY9HMp4YIy3XHDIhPl+W+p3mRl8vZIGVOG+VqLjdeFAbaH635SQ+Uz
7iAPIHasIDdqzZCfokRlbiCnZQ0IRqKwU23DK3Pux7liFyfW4q2domRn8AlWI83ZFGA7Galap7hK
byNabbTYuvHeMz4r/GQXV5AbvVypvTy9UeYbIy50bfaPaJRAXq02nqMoWS6OE1ocIlKYYiGYOAto
v1KrDyhcwKLF4VroGOO/qQBlB9vOm9mFlMuHILxObHGybmwjDrbpD1gPvzvZKmfJlJOSzNISVS8w
otqUPC7LHuRnNKdO67JY7E41hGnxl0iW2ig8DJoQg4g1hi3bP54IKT4IOs7UeaqpONGCuYupID+q
VEHOv3dsTHs/H+kLRjCvi1G+0xa0Twgzli2uvrKtkU/cPdbJHtnP7oAu6b9LNmkvsE3lS6eG+1DF
WIvN48gSA2AVvkmK0+rptYPOSWrJcLkK830UTtV/KUdGDCnocZWZ/kYvC6B77BS1XH+vrrdY+yhi
CcD1otg8VDYhGXrB18stbA7fHpK7GLoZ6I1PQkS1Pi/FKO0i0kNGapIBlRagY9jKMllXKGFWkyZs
eTDzCyadw/MzlYeBCcqyUuug/Y+hc4D5rOrsf+lCT9Zcd2vKvDkC7Q5zbQYjY1IM8dq4ONGgGEvp
4vxSsGyb1EGBKYql2+Nkxkuf74c/V5zq4ka9ItrQ+Jk4H5iNrNpVyTo9RZ1y+36X3/G56Iu4RbLQ
u75YBYTPc4TyXkZB+w0yd0OseO+1BP4PK0XTO+c4ctHMd+W3s9/U3GQQQ7EDpQaQuGQqhRik+A/w
1E0yvvbUGThNoArDL9UUie5fHf5GuUpkzn+HR/lbnSnSn/bTnH8jUP9U5n0wPKw47LhABJU4fSwU
wtlN6VpPTDTyIXTMPptKtUFOrLy80pK6GZFb+l+k5QW5qMxwUMUWic8kTDGNUR0AykjkH1M2IW0S
nR1zQ5q2594Q2ebL9PGq8Xf4CVCJaXfXOFnn93UYQeMONBSL4UGMLypcFcYzkjisBVSfhbw30I9L
t8bQFPeopmmHvzY/wtAvlatk9ZFaiL4BKNRQgxxAIaqw6XNJnA6+hekakiD/Lq+BC2KRG4yHBGLn
GSMESc3vCVUeD0MWL2R4iT3YNfnaj7LI+vnEUOF3BOA5HjfuBdgWlVuu0l9q76RRM1EwI5nCLToW
hJEGxBoURFez+oCl3ci1xxAUC3JlerfhP0uhANNs7ml8JeGX0QsDM7kpkPAWXhF6tTXyEbB/mbPM
ISZ6qH8CvIBNMgHrNCuibOe/ZnnjAM8UaWXwm2kpVfrxCz6Alw2ZYXjuFat1Z9GAMS1SxYXt46HI
CP1nDDdCvMRj4AnL9JB6cj1KR+cIIvfN25M0UbrHc/VUlAhG2bEchtHG4y+Da7xfWER4MZNYMarI
0xIEPPX1T6Nv+NFwTYC/OKYkSVCk1oNvCsZLwTD7ZoSrOsxkZy1pv+qYasW0qjGOd9+9r2R33fCe
1+NhlJ+3R/snpNLOIqf+DcnxjaK0mTE7GFcXd5Tfx2ds8f23KQCniKCGOBKOVtRDSn30AKEoTOKR
HSgxiaql8NvdEBH0Y0B/nbbMZIJeZ+stjoAgwMsMP8Vs7zav2gDLNTJ17W5G0Zh/Wq3llvW8VnVm
XQASe39kWnU5o/ZLpfY81FqaCcsFvNStLyhgCuXnLKlFVL8wahjY2AZzlCsBZXIi61uJbE1E6M19
jypv2k0w8yy7DEVUulA34tpfzkZiibIC6GdxL9p5K9SrSEzQCLhTBLYSw0n1wel17QYsC184Ow4c
bao4z/BRQgjPSi/WLGnX73WRuf3M2k1yRbtSLrfENKulIeQKLPloy0e4mVz6eGI3PstPHAI8Awva
Ysh/04rkv0xGp6A9nV6pVDP8W9ozDYeqVto4EbuH3k+Pguf/kApsv/0ICstuvqKO1sZPO6JD2kFQ
aym/ZBNX/eBvh0/j4cd1NY4+ACCAU7d7haEYCL+8U3ByLcAQwXZKqoqmaalP9pjWeKSjvdu1tQEk
7aueQpohOpK+lCagkXdvL4Cl5DNzkGEZMzt4c61lQ2HWVqtwJwPSGb/cqvn47SCpQGWLINQ+WsKk
ASHgkfFlxPrydfhPC0EXT9HjLkPL0qhtiFyB6JbCNrLFbCeiu3q50rBfUez/x1aWs9Gaq26EFskj
59p3Txo5m5gvF6hYalrRetQ6KiO0FM8T8XBe14Car9akn60bBXdn083Nzlmqstrnq/t9fbLrHPmR
/DyGnRfeRRRLAovZlSi8/JZC4L1R3DaYVu5MxH9l07hWrWqR7LHtHtHdFRnqu/oW7mY8DDaxfX1n
CpaFz5S59vFdSFE6jvl2zdEBbAvfeLzbAIek6eVslSLTEIFjOdIh6ZDMEpC/j4muLHJ+3w3+Qgz+
wPhAr1xcQHfB0P3sZ5cITANRvpmuhuPKikUK5cM6SesKMCYI3OjLcHI2fyaAgDbeu6dTJ7T8bKEj
9veoY2bMyJVuWvV5ZgDCQdQAYYfXZvY1kZsDD+4h6AftoZbghiA8MrWQidNwp3/hrXI/e7ci2spU
J5D4GrhVlEucUfqmz9lyop1QZ1g3FeKW82NWsBgyNdX1qWqII+QrYxSrRQvajIw7R3JnIadRB8xZ
T4yx3yg9aBad7p3gcYF6pdINAy7q4go1y9urBv2vQd8CP16kLLR+eJlCPJrTfePwW7ZvUinBN0KR
qLyg8GsXyNvj9oa5d+R2lmor2w6voZ4gxUlMtLjq1zDzeWcgz/5/4FuWvljhuZ79y3ON34MRhMP+
A4dgCfY25o/1RBUaWjR1Owc7X5TFzWx72mRHjoqZq7tS+9jgGBjWrFD6jlBAdNUsQ0nDhjcrsmBz
V+ulw2elJIfKZw1HVmHlhXoNYdhcWCSm47bhFBUpsH/ymgjp1X+nHeYROKuPbn0TQhFiw1BDL0vt
4fsjNL2bopfG9L9dVtnDh8KlvK3wZ2pYJ/gWwmwuUtqus38SXYDYGDLFZTX2zmBzV2mweJ4hM0zn
bsl0qDgo/7eFB5W92crj0ZvbC2d/rcAqj7DMuIPic3khLXH3lSag0iK3eIqgIcC5Ks5dmJFx8Suw
kv2014dk17dAB6sd+hhh3mMuyANFD0lbnWqxddAZB7kFxXaa0dz3Zy7xxlL9nQzUtSM6wwDnPNSe
hz2jy1fetQEQVQ7oEhXlykHNQBVDgZXE5oleBwv2v8szbtDkn9GWrPMV11nyeBzR1+rsrZbkdJh7
aVhEqFFSPeo2EiLo34GUThhFVfr+M/lABCRAzt0X5slsE7WAkuZaxCq5KBBlJph1TD5Abj/FlpSX
Gx1T6WcLfwoQXWu2kvOFvLJ8tINAJ+oUtm8QU0c4sO3XCZKIwNlDg7y30FGVCG0TeIF1hFDy9Q02
UpxQcwpgqIGabpvuwr5AutnEOO6Cqz5k3ADlVH8HOwIY2qEq0RZursfs+Z8p/6Jw5Lokl38vsSX/
uzsT7o3BJvbg+q0YXt+Ch1KTGipooMS0lMbNht1bqua5YPRRrGeIxI3c/nwEtNotGAOQSyAq53i2
uT3Z3rJq1U6HMGpfCGI3fbnaeaAhzcLnaqSJ22zShKKDMQWuI/0DfGRCBY7X6NFjRpS9wr/ZmBCa
e3sYbQvGcD/wEFQ/ZkiYCFM2vxhlUv/FtWvVNEP9q1diZo594dLcISh5zQhHcgl7jgKVpp0KEDpB
bsJRrRREooOwLDWYQCB4+P5MiMmRNjcT9xYZroKa/0ssgYKFo4MNRHa3JoBthoOk85LwO+813bHo
Rpci39WcZ7dwWvcwyFt0iDSqi6p7KSIkB+8l3QM6ZeIRuHI/zvcCjUaTfozi9CBwrYRfeay9MMKw
fip6m++IcLRTSmwB953ofANslF92ZMnUsbnx8eAIHtMEeUwR/RxVQGl2z7j10o0O/opdEciVoxe6
YIoph6rkiX0Bf6hjoQaQAeG4YSQ2hw7ehC4ugC53csXGgYtPNWs7287g8OLFOirbYLVIWOqqOAXC
DioIE3zeYVRXoKkeGlm5BdHIQOBO82hwEjKiiN1dhplbCkSmCxyFK3OllsquoyDN6Z+QZouJYWDt
84OvXByznHQ0uK8OsdDoefcumbPdQT4zTPU/QzlMtk2LXVxWbOkk5fUr/d5EeP19j0T2CAkZPR64
0uPacoP/2EXy/Ezm/+NpNep+w1rSMMEb8lzmBWN2lTfRtsZBxiOhpmQj/gjUVgj6tL0DnChl26ki
+kOKtNLaLcDCUPCVuuNlfK/RMugGZW0lO2xGnBBbSpS+w6ZDtZjQD6Z7vSLo+iUT3i7V2WmXu2Uq
GXxySq71R6nw5BwqvE3bIzyMTLQ8NB7JQ2/nZTJhjev3edz0CgJpQo/T0feFy2zIZacY0bTFViPA
YBDggcpuv8lm+Ok7NwdsA0pOLjaSS6ulu31f4vU93gc6yd7a7ugDinN71Wr5j9YQxyAzSQ/mrvLE
beTWWFWGfEztV6miOwBUjixOmhNFtgHRTkj39aZvrlgGsQxnYaoW9sOwQ/Gp0JmfBK6ANGEMDaRn
tIGnMCUj1wjlmnM2960vivzmUF8xLJ6VCJbYA/Q18gnsCYX/6vO/h+BAwjV/hKaXKAjWbVxHV3fg
gVHaGqNyxg4zMlD5rZ6ZuhIYzIwF4wl6Gw8XRyO1PEZGvtw6YeNODkHoQAHaknCRnI6C5wuJp0+4
9h90KOp7r5TShqzPMO6yGEmphk/9xbFRVj7Js/qS1fQfAuUcSVmwiIjjSBPgI7+wZVn+cEwzMdL2
97SlO/T/EOkkvm2brzS4GzC3s/ldViEkvs+mbfjqZ7/TR9IXwMWeCIQQ3/YkP1wn7ksP6xC/nf5F
uizMlaPzTxmvnVagdHYcWJgDfIigamu3JTcdg150CdxqUETDmwbv4ZfZWMUxql6kAkb73fbr9IDn
Sy2kLQg/pAVqAaOwY8rPJCmLZig8hKX+i7Cp6DOgN13tj+Xb0owWyKtK04uZNzfTkoGVaE6U8ICn
gJ+nq6znopmFzcuCIuYps/mFHTfjEsxO7eU9NGjILWpLVYWVZkctoduXB5BLkgFR8gOD3NUZKVDG
MftZh5c7IovjY2n4glYXMFvzv/h6IlOoUpP0pAe8FUZgtoo1EUxGUTKLIOUMgC0egf3Y49dNIVeO
06QC4+LD4+YOgu6h5oVfrE9WlUdr0NNhZv71URX19t8NbJwzPpJAX7pyyDsZswX0RSoS69Be2t+q
C11CTYpGW9C9lTrcyd81UYgY3e3FSlK9BwmTs+yQrrXO1Q7WS5fU02tPo3/mXKeC8xL2PCoqah5y
WhrL49bdx0TpL1aaWaC4uE/nvw5weiiPxBOP36PY42sI6HdtNxJ7HKeSMiG3XPmD82g74q6NLfng
tlKHYztB9S6+jbqykh2bNLoYuwNpN6kHQ6Bw6qAq1U3cuBTHHPzHnyAk8D/+8drG31yyrSF0ZXBm
g0UtzokKk3427N+PDnhATTEonaP42D45331awdkEMdFpo8ndfAKBxKysUL7sFJtgOAmxLvDoVv29
59kL1LIKwm16JEkBLVmI+rW+xZPxxq9bbPOVtFDM6+jtQW93JXcoQz5aseAl8vZl1/CWXfPOAaHB
r8Xwki/1FGCISntD2eOhwYsLQgAPTEFKgPeovC+3Q/y+i0e/oBtM+1JN/RuQRTZF+6upnrd/mAl9
ndOOU1JeOP97vBpVCs8gDCQvE3c9SeD0PRZpcifUI4mqdkE7jk5T/HDeIIpqdcJkwFf62+k09XgV
f4ohi8ueqrHZ3CvAkcq9LSWQrUow13d7ZFWbx5QS9CuwtVfpmrFEmk/DMZXMD56tXMuMuzkep05m
MDEKM6Foc/hz2Y2Es/CNj8FFIU+KCH6XQStnR9Pb7zL5P+V2J/m15U99bk30NJkv7U0lmUbAp4Rr
N0b8DK5a0LgIgD/tMqv98ouPI+ELb00wycQvOGs6cTY8cJoyGqS3aPSOLblnHFQ325VwtPu82Yap
pxphUxeOCJoPkzKk6pPEHyqsdQxXtL5MC+9IVRI7tNfyKL1jLjyizM8wrN8CxSlFqNvcwZ1RBuf6
/DP2lVf46e6NasLrBqJZQyu5aB1r+42qC4A4OkV4jlff4gRXehB68WFCnX+SM+msVL+PfWlLEAHx
bKK9oEOvvorhWR8goyb/GaRFE+uUJJlf9WEn9By2AYtv+wDe+crLiffDlwh0TvoqeTR7L8GYFIHt
YIEuRnQutgG1vmu4sazuUAonW9Oz1zgavywEWjNq2mbIC3Yk9jF8xsvPy1NImEPrQgMGEvYCM63a
SmSDIcLJuHBZZef4rlfYRdBNajIZ5vDG+gIQ5rZoxlx9b7t68sGReYoTZXPo71mnsqo6DCR4l3+h
ijFtp4qSoPVNge0eyBvZcJee6pSgh4iGAuri5+321TdZ/Olj9U8KbbKf+TE6BAUBLw3L27jarZjV
bfVc04IYeFwRHHtOxpa1KDbjkqsw7ZRIsHHHmViOZaHao13pgBBBAKmSIJ2+4sYI3Q9afXDpe36F
M8hgJCMUDfkRhvMBgZUKHgQieSO4Ri5euCdIy5qvCtCf5Ir8xt47i3gbDx3GRKMbYj9cr6Vc4FWN
2AhuW14Caw8hihvKmgQFR9quZvFGK6a4wbsRkiV7LsLwfHyckz0gBbm6guvbkVYYBr7k5wPS9H7y
Px3iMhxDgWsueHeoH2bJhQrxgGpmT2zVaqaj0x1BgDnANLKXPVD5bFkYBuHJ10olDqwnLZ0lC25v
cmiitS/jNGbNi71gWZ2lxpgKs/rR9PLVO0RJ6mm2QiKCl2mlIHH2MXCuc7EorN+m/G/eq9vwSXl6
Gt8mVxz1IIBWog52NJRMYhHJyHzA5kC7ICH2h+Ppr4oatJS1wXih8RnJK1ofUOvMa0JeWujYTLQ/
OGo7pSw3hd2nX0tM2T/sRHEsIZY6Io8NabX2VtkyZMeA9lmrJ3grtV8to/5KjpYc5RMNtN70jU0Y
apWswpwyOKfdRHiO6Ddx7ks8RHIzmNgXUL+tbGbScw1wC+k7zpy3g1pF4tUNvM62/D41xtFagggx
wH3iX+/Fg1ZSQYlUyLBkiIN7/5Jvmkdh8TvuGH0WHcqg5PriKHy8X2hVGSiexkOynSex+n6npwbD
Im42fijscxRazmLbBtktcEHrbryFFOXggdKt2NInsDSIvf1lWzxauFfSDKJi6uDLlVDbNYb0QO8O
ul0ZvCObwjHsIwu2evEEAAtCIldohA5Pk1dFvfY3GGPs4PiX+NKB1ZhNiWQTdOgmZPCIpPZ7XE9u
dt1eiY1/boo7Rk2kuwSKUDLRz3cDL3x3INC34w9kUGuACmfICHaS2YwRbsU8DmSbah7OLIUOkU/j
TCmxS/eyz+BCa01cFP+bc5Ph2KR3XpdiJPStInQNLdnlDaBf/n1mMhB8c9YfgnbND5hfuV/42xNj
GWRJB9xaQWqrllCn2jHe85+tc8w3l9jzMkK4DdGA39mANUcvd6SXaPGXmVMbL7Rhv+P+M4ISAYZM
At74HXNA7Ip81xwZDBdRL699ML8g2ZCaySJ0ojzIZg+eIiVTu5elULsBFaudU/og9sPH7BIi4YBu
ysgRTK9tDNGUuqFhe3vdz7dOWw5BYsdYg+oVmX76EMwce9kHqrmxAhHCSoNbH8YzbhInbTTdhiSA
Gqw3EC5Goc0Ny96esVvz/rzF2NrtVk52s14C2BVvucP1dUlkLx4aDFs3/KNpYqUH+Mpm+g/Et/pl
8ceU8McVfC3lZkvKnhP7mA0EsdnrfzK5GlW2ntvbFaexv4hl4gWUCEiQev4wNUwh9eOLhLiEUkUc
tSI3vf1ZyuwtYapierR7XMBbx9Llvc3VUxHu3E5fE1Ms7UdVCeGOKH13j7Enf1nmQfS+oPBmTiB/
AAxeYGZX+/aGeC7NpbR4FzO1krQ3Z6W3/ZZyOFfPhpPZ/ovt+bvkoKje8szEvNYhsfjzpqjuDWJl
wEfYz6YaBkohDzbUyRaCp8u70z2puMpygwheXCnMMX/riiRflTDoZooNREDLCCgfKhcXgrztebUN
skz6yXMkJHUjt+NJ9ot9aqYs5FltSMX2pEr0C5AKMGNvynQ0lCEJ0oYOF0sBU6iQPHOyhCR3rsgm
ceeRli/Ttde6H7ArhAkh5cEv2sX6Zo6kSwQjDaZPXA6zW1OSvm77EEYOLN2sIwW2GJw1Ib+adyG5
qAmfWk9uz7dBx9GNjgor3WZoA7HRjI0tT2qW9zevTRhS009hfatR9t66biKA9NlhC08gWcqts0ix
dzq0AaYjI91jlhPP4wjJleOdDP2B9tchaoXJnL7pNsjtECvXkaMpzmPNvmbuAS38prEfCL67vvF2
Y7d9qu/ywkGk/u6cMpsXh4WXPJwfT87dfsDO1AHspQ6TWG2dWzDvAyieadpWje3N9axVJQSycZDK
RHV2Pt5+1ktl+qWB15bZN8vyhXTJlUGW3rRDWMPkjtvVx537AAjiteUwrVVFAvvTsGlQ/7HAxls7
jx5hlbLaHqkqnsx92fVJ+AMGpQ/CZFyrCGJmLO2INGCoNM7LFVf3V6nmZkg/8X3EaudYor4FUSaW
h5gIIIv0oYRyt1ehwjvIby6m1o1Y/k2ugdwST5VHOiq0WIiN3bVAiEzvoPv5I/g39f3Pz3hAKFeD
oXcYTmBF2NPv96PqNCxMssrtsRQ/wcWinvdr4FycsRnRJnj7INRzvxcTh7kgMro3fu6e0EBiOU61
XbLZcbk1yZIxfPSFvhlSooaw8gklW6Jnn/XKsKLwTzHLtv0j0RNF+Z65jU2X9AQuQXv97YDx2WLO
AEiZM3oBMI/uaNVlDqI1wiBokWoGj52tbqzMqXgA5EEQX43w5FMKTZSs79hEbHc8AmGqTaiFrD2E
8IencXNOm0Dbcw40pP2fjrPazNVl/Mzt08oXozhbKkCskA5xidSyEOFcpS5nTYKJNyriwbe1jdf0
ayGPun5Hm5luWvLCNiPIjDybkqTED6cyZ1kmN9P8cxR/klpzl4G7yk75TAEKOzrOWbX3kH1EwqqF
D2DmR6lnLJZxRzzQ+uom+9DP9uOt5H5I0p0VX3RVVkWEs/Rhdmi5Tl92nleG0YZUh7ZMSX5iPdTX
hLL92lnL9FyE7Ecq4wj+Zwfi+S7fqxWrVg2khMTV7yyRXwThQtlBXg4CdBlGs3UqkDVjDdAW3ZPB
C/Tgzx2DX3ksLDZkw4kTvsLdOOikXmg48eoFJkbefRVoh1xeIbCtCmsFWBvEOr4g7n7kurzy5D5q
fN4blW1Ioh/3J48yIMKBExKzNL+5iyvpE93aeSYpAGB7WdvLB60HS3xXlG3uTJ09Q0idseiN4a5o
um8WCAFoygO0N4QnYqnkzHtO73dVLLTN49fN2aXtnPtLfHX4Ir9g3dO0RSAIvAp7GHCsGPmls/hZ
3q8vC09jlNiRDHIV2PSTXOz34J3WM0GXrF0YhqPSspAtCHu6fGnytqxoziHrSB0/PCUSM8tVPRrJ
Lv8vJnnCPtY0vF52W3T4YIGnMXRGNO5VzGLx0ChnTFAeINy+qNh4TlgjkPa6aOyyrjvIaLbfyvlI
8GgxZbDy51w9OGcjljE1wl8E7UBYuOstCUu+qYvA3tqHIiBUQNySMF8q31OcT7ra1y1YFJ3LnSMb
y+ZXRsmrGS2GQjclBs78e1wXEF2a9UEnn9kvZclDDAR86hGnEbv0p/ejL5mcVIX2z25QQuagebwS
Lf0gEYPN4by5mpTcGKm3Dkx9LGogrGuh4GBEjnEo7cKNBmXWnvClYrhkmcxiE6yNMJwQsL2pIGx3
Aw5RzQv0pEGT3nuaVrhg8iVhFmxV6WS1BGAPhEDUEA2vd/ybMW9f4Iq4uOmY7l0SX/ZPH5P4J1/K
iHKwL57bQA15NqzWz+d7Nug87pu8JHlGxgevJx7aV0FlgCXHjEAagV8qD2c52amkfWX7/Vz/cswC
u7hERGX0IqCZjdHJdh5EexRgXmkpnPh2d5phq19gMGs3G2PI5TG6AcuvtLaa9mV9gXlnE6V1IUD8
m9l5jjIUTPlBGaBm6aATNo+UDr7ya9vf5fuGzS99Qpns0GXtzGP1ryDJlbZe2xx49fC+c1R73VKj
8t9rRlmOWIWbJP0aC23sDAgavRfy9QSA/ujYaRLWBzOnubqBdqslivGeU8+Ps0uYpqswlkfZAtBs
NY1She9BKVi8L9NgPz2BAM0W62kDEtvnM1dImpIkG5NYaYfeXq4ZRemAdjZQ/8qA8WVIr6pkSPWZ
hq+Kg62fNriHrW3cPIQC5NHAXCqXjZ0tCpuMKKmt/8FclsZQ/hs3oYAN4Sde4u2LQ0srivhQweB5
G9ck7+sv6N2ZTxUwh9y8dpDr8AxHNHMBxVxa3XzUbA8a3FzpErNAub0ziP9uT3bfWEESU5lrN4rd
iUiDUWvKc3Zk0MgDcHtKLS2MFttBoLaHCYaXo0hcT2LOhnLnV7jk19XmLOI6AG2YU57geVzIJYaM
AEjwFYJ0jRK7q11UrRXhcqcjTMGxSHqUwFPO8GY0ax5bnkrIl5FsCHTNgjLywVDyEwBknmju9PDd
ZJy43jH0VY2p9psSK10lIPxhvxh2rpFkJC9HiMru+i6VJE7qpWTv+/yGsGou+IhL6ulm2/f3LHz5
7Iv9gOQYLjEM7O1HsMfAjuqLjxxKXpTB0rikv2FW0RsWhXDjw0zjtKN6/ms+tVK6RcGA1BHCxRM3
jyjXQjIVVvQedjqhzkpgJpllo/B5GJ/c6/nTAd6qGfjA4viyICG5AA+OdVe29dOg3WfF9xLDgMlA
bp5ay6l33F2wxHeWLwBwP3cwuy1mJa+8S5YW6ltgyKK9/sYyxy5km9N1SGmLxtAX835VkRgwu9RP
bL1kqOR9gB+9zOPJ4QheNlQjcRIO9sFrIgu4EHcWGwe9jHYFkA3++IC2uO/HWoe1Pa7X+AB+Weur
YsScovOprauPl+fZ5gWW38jC4RkGcUv3opY8IFjMZYntVgeVgIXJEEyadOKv52lOWzMf+GOte1zg
dqfNgNEqSStaC1H4kgg6S63MObC1fnpaeywHYVQf3jM8bsVTPhPbyinlVr+lbLAmHoGd4hc4FbFm
XXQzUXO0V5eVVMV5lIWH4X1/CxnsqXtt2B9J6HZhLSUex1HXsidiUf5NCg51WfsR6LPduU12n3QV
BXiEpXleYGhOnytoyIg94gyiBt5zAlBSDUN57HXS5ReT1y6L0z7VzCizjKjP2T14MuRl+4FOoNV1
AE0l1Yw9b+7BcNLfZaK4c1Ke9QlSvqOxXqf+uQphE4GOaGTXucxy7rrGW7vaQ7FeJAlYJh5t2J1x
PiIR2O99kVAN/AeXuk1kuGanfKXCPNMR0fh9WlNsKtPishrHMAMyuE1z5r+hOWJWVC+K9/WdqD6X
nvrcLRa+E5QFeGP/QCkp+cWW3kuR+1RLFXW+VOaHnpm+A7DpeqvTxF3pUf8qFsAAGlcqgN+AJQDI
Lv/AKlqZths96rnMvElCak8wDWT8+qAF/qKupRqvBMX5/MEdLlsjfsRc9FkHta635vPiHOzMn9Em
ZZ7d37WjfpHEMWe/InyyjlFTSqyNr3SmmGZIRUyefkkNr7oksIbocyUBws8IT0c+n2nxeJj2hkrR
O2Zz6w34pmTfG/f/Sg7ezghd3XjElncjZIZaIfJCdY6Sib7Feac7pDmCbqnd3dAuTQCXyhVJbIX9
GAKoXN6N/6OMKAcXq0IvwpUjEulLR2WuQTchmh3BBDiENJkdDD7OfZTORy+9dqN6SqktOyIlkElx
L1r6KoF0/k2C/mEW+dRfic3m4Ywjj/V9p1q6GRbWVxnIYyP5+PUeqUzvmBcwtxxd/chdJseJPxl3
XlGx4BUbSuP4pvC5b01aOsoTVSSxg7mM6zrJfTyWW3UmGy2pfQBGRbEyquTlHTwEy48mavmC+9if
1Qp7tJVM7P4WD3cka9bmhVgJlNk0egPcXXRGqIL6g+5v0y3YJZBGSVMs9Qa58T7xvJmD3KkhX953
FVNULgCRvNrLMy2vEQ/e3/50iULbtB9fWCrmcXCrjf6KUTpO85oKE3ukVTi5DTb66xVcuIjwhQ0S
LV0ccl3CN8dtStYzjdmXrPYFl6XugEllYT1/UVNqZr90S5fD4Viwm9zPfxdHIXwu5JrZq3W8itF3
HSb4sTs22SQb2BTzgH0M3zlRFisvpoLspZS3lEmLXOgJFhRmTxr9CBTIyE+uHOQQU1PYK8I7OOBs
3AuZ7zSzyVDLm6JjSxEBchCOMnPonpBjCEWhwWGvw3COm0QelHaS9A2eZhcasYTiaYJ1Y2AxBp8l
tUGyTv3bc8zIZVA37F2qc6Ix3C8FWygYPNXbcZgj6TOudzR4EgIp7iMhL80ajwRgCQYiIcTBJkLl
AmdCg2Fr0a91B7dlyGUpNCdqW4yk25r/5xe3iPIQi9L/O04nwWYGUw4aNlFPD67gUwRcC+9R54Kj
EeXdjNXv+u7kibCu9bqsoZs8mp1UwgByziUnMRXs9cZo1TDG1seHg63tUCLFPu07eBn+QGbBx5sp
nZi9UxVzxiYCNpfJB+q+2ISglWTDLQF3yVRd5W5/XK1yn8BUng26mX2mdAMHzb5PlWIlwKHbq8PE
M0l+5fDRHP8I8ycLiPe78VpRp8GEmCYQc5ncPcE+TOVAeeeM7f26F0bF/DUNftTxJBglYZntdObJ
s1ByKtjSFKgO+Vju4zyrY09niJe07hna+5cjZ/bugAkeF4G6upBehxnkHew9WHrV+L0MA7HPKry0
pHwIaWt2/ZfooKYJV/oLkyL3/k6fM75AsSTyI1bzk3el9DcBkuGSxqo5CZRh36sVUX3nUjUxxocS
s1xMlf6jjFkSD6K1fKDRPB4HW3QyxDvcIttvtbFJKcO09m3G24tAXzHSok38UVdyPII8ZUP/HALr
1QuMfLhAJGgUR4aTzaPKaQqOnaJdLZh93IcW+5Wqb7OJiIUxmO3ffMMigfWix37c5NQ6PbFI64OY
E5hqjorpFVJkNLSTaURCRWOgK2V17MHC8vlYgAzl6F8/F338B73NImPwZX3AJZM0k5Ld8jPzCj0J
b9CIwXUG6RZeXFZxdzmd7Fjpop7+iNAxFa+m09kMmqOHTkawBLudvQL3h0OA2w1javYIp1IYqTXC
V7Twr6qaQTHTjaTP+8QqU6EA1BMRbc1ExgQVvXPm0BDnhcyknVTMcUP5kQF0EJQzODTRyirPbfR0
YW2dKsC6QRoqE1vTzE6fuIQsm4+64B28qWvw5KAlmGprykG+nmqvgM9JgEva/eezoxYn6rJex9jN
k1D0itrc3CmbSbb2Z9GJM9CzIn3RqrO7GKaTv7/1kHY1rTNu96nXcnoEh8t3u5IZ/fGy604wziKy
Fhq+uoJr1pHUeF0CbJSor+X/AcIbvi+pIEZAxFqolfLFceEFFaaf0f2es01wqQJ0X7csScKUw4cJ
nbdpUYbe8GQZ97Jq434TlkKFAO+u3FfQ8a6m/HmiJy7CMIeWwQUFly2wYLGz5c7O7LtcjLe260k8
FppgSo+S1/8wcof408l458SW2vhqg/2edzme/kcNoDO4VfYfwlAsevulR5qCOmlVntjw6cvXYZl9
kblS4ppFl5NGYvIZvzW7spNASnG3s4O40erHC/MrSpEF1g+pZAc60MnrUlIvp7Sz83ZInjJ5kjh1
0mNtu22cKGVGDdLHecfGNcnqg0bgVYb/QyFGdZ6MAhrh6oyY1+Cce6NdtoK5CbnDUK982DFYBCMM
9kOfknhFOxRLsqt7/y76VgT9PoU2RLurXYUcPrsetNVCGs1+f8hwPXCE9te4dyDEpFbK9SlBEATh
i9VCN+eA9E5pOnD3estmN3kbAbxeHBsdV9/VA7cWW7qiGR5FcL0G/x8xj5lS36KFd9GlzIb18ze+
j+ZXFhRFO28JqMEJO79bryaVu7HunEXGZWttKDRE5g2nDsPf2GsVpXxrq5EAu8LNxTilQWhKICsQ
OJ12hxaPm7oOv9/QAJ+CXzg3o7PjibfHFfGJTUlMWCu0+rGZTh4xiw8tCV+4/R/vTs7TQNg6sxkC
4z13ec+swKdXqgoXVeqO6pgvBIRrSYuZZqhpb5/XrUS/GWC7oy4EQjUp7IZ4SiMGq+XQd1aYXonP
+nu6r9Olc666B9Xibel27Fc4bBVrfNDv0xnRqhBCFGN0RSze+E3NqPiA3h/CIhaulefTfaLuAwkW
U6oiA9XDRE9auf4I7OIf4npYhidNTzm94AlFKGPak+H/hXFQ9QYT9NwSRNpUtkD2kiRBU7hZSJlL
iJEqVHQqI4nRXDArH6YyurV/DfEWu/sTQGPBEjPnSP33F8y0xHZZDGDf0jRuQn+caz8sKOsOkmsK
sFA9mRjA+wwFCvQUd+JwAy8S52rLstec6USHS4CZsTPqy68xHNmBIivi3dEGDa67nGc5Hu7sRC5f
GjgxX1HOu/VQ/5XBq1l0+OXo8Ce3R1mNPJCN3aCmEJgOs4adnvWDpobZSh0ZUnAgBq/nktpRpmHl
Wwpe9zBc1MNaCneaWJZ+jy7yNNUjaiuWLdDe8rwPZy6Y8oXgJBZFv7MBwIz356FH8XccNDGC3IMg
P3iXBt9MHMUzjy98cUucSB+13qY4J9+9EFVk4ewrGs9VctFyA77CwNp7HbSEjpzzXszkbBIrqZYk
mPh3VQp9eMXpDa0DFKbshD22/rWUPqej9q9NMHTNnns9uz14bcL6ga8KURgndYwIToxc0Mem629U
6JctkrNcyKqHGO8YyW7tiGAXi04UqnubuZD62mou+suct18/ZTfzV53u231KOy0YOmbuS7MnIKrx
e8VoIhzbjF1WWTci4fcv6XgwU0BRRprpS6Oc5wSaP4BtF3bpHWgsvugmYuaB8JDltaw663erU3wu
L9Ok/SLTm1mZ/PJvVXjwQ8pkRJXMrIaFH5wyFXJPcagNhoaeXTianJ67/xXfzBdENW5S7e4dhLRV
80exlA0DiRGzn+D6nVIkMY7XGi5KUdD5bBeoHYKlZXtPui1z1I2wfFHW7OcIzOj+m6pNGOPuwap4
3qvsoZOrMqvrmJkoFH0pECcs4ZYhMybLVHc8erk0Wtt2dAklX+wCB+T8HxqENfRJfoBZKFRvOPMs
iG+qqf5/UsZQq5Eyb71q4Gcx+Knq+PBi+8R8DQ64QZaaLTPgfq9PQOB/PB/Anqe9ZOfLRpVUwKIA
7hP6OHNU9m4H6C3DbyT+4vZHO0ZIEpdTtE5VSVe0Na2vyhUpUSQF12kt+HY/gahWKjl9BHPvn+7Q
jTV11/H529qd7jXkUt4WfpvAnkZe16eV+/2PMbnIdHQr5vT12F0ym22yYygma3sL5lV1aV7B5Jxm
XSeqdscakv3jDlh5Et9IDEUdGPK2N+RSWQxxZDlyRAv2xAscGR6Cfmr9ub7fq8svN6Vhr6Y/f2E2
RNnJHb0x1qz6Ea8BTzqbzLGIyBSvm9nXRDafFRfEdm7jrMe/UHyYMZ8FVIXTyKRBSfzVhfqDBdf/
eZshzIlFuttuXsK6c6BJ/EzsAGmsJvHWWiJMd1MYFFLYHHybU91O1WNT4m+WwikW8meIHZLU5Q9/
JTcLFHOqMzjT/npMfis0k7ueymj7rlmzbgOWSHPuH1msEJD3qNoEnkHHJuEesUSvA6eE54Rjskyb
1hvfS1dDZ8Jw3W/En1lujdlxE9e7/2cUePE8Wk7Q9A4usKb8oayipkbyxD6EK8N2Q0wfkvO2K3B2
4SqlSGyNGsA82alGUekDruVTBgYSfW/EjdMNhHZJJwswW225JPzoSAvpZbSaCYS5cZ/BdS9hsvU6
XE4A6rwCTV1XrBOn0dWmJL/59q5Xq6mVt9CSEVBN1kR4yRR192OAhJG/ULuXFDBbuT4OO/w6SkS9
SEZ4wzIEBAsZu527sjVP+37apeKDqHkRzolYnmkQhq+92FSCa5l272iD9YUYlfnMGSBfCmQOsEO1
7PWf6yDbsQ0WZZOgjtPZb5w8MTnXc+7HPbAjq/PT3BVlYvBSrGR9qH8PoCU87cIz6NTltvS7cJO0
Qm1tBgQ7ttni5JEI2HIfncIsufTcUDN57Chd7PRXOMoIAdWhZrwP6a7/sJof2hhwzgikgcS/Q0xj
J5yJMj68dSfjEcsjaRD5LjuXW/fQs/P3KJURlGE9bp27GXwYHiUmcq4lupyF+6dk6hxn2u2PrTqF
K5jaXANEiL9cGffVkw6YSoJqqz4FSYdBg2Hv3zfBnC3ZHudi99Pp6UH9StksiPzxrNpUhiM0unJH
NOQ9Tru6Zdiqzl/uLayzgRdbcbjwGTKtBy+o2hytu2xCalsn21v1jUTaUdwsfAV52F5Vgz9HWcbz
fT5b5x/fLjHaqC5Y66m65gFkA86zi1xETaQ6q4Eqo/g6EzxeHOTRSRG/waFCFwTVFpFhs/Fn1B39
7I2K5t3laSIC9DLDlFsU89plaGESrqP8UGFzd+AuksnBVw3eRx+NZWJTXFfIt+FOOqI17UJ+IoSP
aqzAQwUYTEjf8WEc/7wGAdUosOgUMI6rMlqps4xgQPDkpEgQP3RD6qpBAmPyKtiat/otsqxA/QbP
lYDZGLs2a9Vx0j+V6fyYKQ0BFfuO0HSc8ZlhSfC7S57OfTwCE4UqC05mGtHTILkX3E3UcCnyYA80
UQJoh7gHZimiaR+eewzbS3baALv8sQp42Ub6z01emR1QFPzh84QlX8TWt8ypnnQpfHFVW3m6OQ5y
k+OkYDT08G57MorRx9aeKV6ivl5zq+b2Fb/k7LibbmZNQJjJJZQ6kAji3aAofrBw+TTFtmHEqRwg
17IgZnP/uxeUAxMueNX8q81Sum6fj6mdg4drHzOczDZYwnFjevk2sfH+dlj4JWveQ7ZA7PlKMolt
SkK0dd/2f8RNOAOjk4iCCfbLAxvxlNgtau0RdBOE1RYyxkrMc588aqGHWshXLvg9cOyPeUsirDFp
e4ScRITIRXBPFlDApi0egVjUuf3vdc41d2LM6fYuzV0WQLa9ck05uBuu77cerInZWzuFF2x30zIN
G3s9FuhGan/6EBDs/TMj/aSNOSEmkvnhR1Li7YmVzmJf7A6wT3andB8IZpTRwwAFCM5ETbSYzxmx
xX5RuJeUClZMj3YxdkWStBKeldpTmMl80YYQydauHnPhHn7m2RdunZF1owR1tuonqx2GLedZwxzx
+BuYEMdskuKsHAWV3ntXvlgI0xcdpU1qUHKq6b9eGTgdGB9f9cU1qkWt5+fenOCfFDRik+BHoRSX
fkyKbecQOP6iSFmgROr6Mz7pKPvyBkcq13fPxm9HnEFUtEJzYwXS39bWFQ1yw6MqhQnAHjHY1gfY
JBGrRyvcm27O+EpXRhxs8SqPo8AmtHcTl0BuW7Sp96wFi7CnPyTLqwli7kP0I0iIOZFomMp+6Egx
WxOaNPPy3i6CXGlWjPgIuFLQtrzFKk1MJyP7vkymFhK04I9Q2dypz3MzAMkZLmAYG9i7wC5lUNhq
A9fb4CNI6mpNIFs6Tghkl0AmXjE0WFyCzjWSZNgdeGumbmmHav3VIjR9MuPYuph43cOFiTmJ4NFX
px1PvQyCTl+2UETY5GNQWkeTK8IBklVUM/zFjZYch+tVjJYlETTdjV97nURMwxu3ZiFkuWWqkuve
2eHSlhJM34WmTyz/J/YQNQzhvchACNCCHj44CrsQmLahR7lEnd/hxvMBAoaj/eG8+CFd+OeWLTQL
U1EXKJ3e0bjFZGwWSWuU3ZHXL+DsQSIXPDBk8Rpi6HthLja8Q9oSfEx4QS0hRKR241qeZtLAA0PD
cpav3A9nBlloPmDSYRFeUC8Sp6wI7ozP87PoypUgnyIAt2gJNJYZMsXiLAnfesnPRnnYRKO4NSZI
/XH35GriY7R56UpE6GQjfvXUpSFv25Iqnab3wKjNBw+ZqRzDLX8j6EfHofXOSezSQuYlmoIYMbHX
UGxOXyzgcZMjng3DWvGBOt3tiV+TRsdBP7WOO0Epp9EgCSk/ql9hyakEfqhO2cvlNr28ZWdvZwd5
UhamklGkX3ilzBrIZsAGctJLqmPVA9SEodFqGmNlP4JRyZJZSAY8WUAu7PKlm76j+guKUz/wpBWu
UqHwPz4YR3qvXoxZyWzj/tL07/52gyLshcNn2YtK4lFxnvpJqEl+K+AhJABTjSYGiZj+XgJgFcyH
ukneFyFS7WJmSYn7DCJeZv/3b4bX2d3uml+czxcIijDxzis5Xu22JdX2ycJuleVtvYBF0IQdSrpF
lPdUiv9mCguXlKjNYyPBUOoBzQbRVhdYyskhAha3p3OxmKrB9tVPOG+SQQqJdzkHiYV94pKvUMCb
EmqjPD0CA6pezABclRFu4Qax7yLWMa1SR/MZ3sczE4A0dY8SUBjcEg3sKhQzreE1fr4wJ6vhHsie
7FfOPtNO8O5yoi0khP+s+Q4t/olv00nAHRA+Z+ytcjRktmpEHxO3S0vfXlPWypy09vHZWVjlbtII
hIRsDB3fWfrq7X0UrR1OG2UHrNwy2yGFAQgUkH8yGft/UGMdS1b1kydhZw0yLhu67+886n42UfOo
bi5+bKTBjzMGSZZTTiMC/GR/ltERaMk7r4siTrgkE1rKF04aRaGPbXrZ09S3TrkwXo8aHd946fqk
62/0yOIdiSpegLsSdgct/UMofgBbzlZmFZlJBfyY9THcl5789FAayZlyUPz+vBptZDN0AC+z9jsj
rYvQKqjW/zC7mHITTj4flvAeyM3m9q2Q9LvyxEd61nFs9fMkbtd7K8Baj5yVyImiPKotLES4XWFH
UR/NXG5n6Er9MB8gn3njpyOY8tNey5jYZ6Jh0rzPAY20g9bncjOHvaKlx/yL1XXdrzZtwVkyzflC
RQaqqy3zBgovkbtJNQ/0S6s4Bwz35KEPnH+NrXM2bvmcL3hcOmGQuThTnT8UagpSgsKjoO/CemiU
6u7yoiuUAjb5dmd/LtqOHCa0aXUUx8YjbY7fZihLOSieq7z68LgBkVr/wVsU59D7lx+BHn8YrOBX
iV1GyvL7Bfkqzu/L/uJwhM3QcfPpbO+gzMMiU1BEsEc4kKtKsuM4XRxyVYSfhljVngVFoUqM/AkP
6sFjqHktNJdT1G07MKQxYcbTrZYskD+7FBlE7TaOJ3QEGxFLsfrPvf59+6VEkScJLFJ10P9YDMl6
hpdE0dvnDf7le+lYyWZMv1esJs4RxUMdj1ZNkPRzzKaxcj/IhkSFAqmBzInnMjIpbmKLjfKxB6M+
L16rs6wKlFQ+LWYwauwaKompfkczhyXX00gPA1kU5FaWMKPVCVINQrQK6/Q46S4ntleVYdn6vQLd
xbuBKVa8LS6hiyxPQRnXtKWTZ+TeyoErQexJrWrYWkOUVnoU+exuvcbKByIr5ZY8FjC0WnEXhRDn
2IFg0hzehQIdPYQAvHs+mf6nIsBkvH7/njkKFUMnWc/eNrJoUCKPvetEOEFPKfhuJkd7PY0Z/3VH
aWZkJegfLUxpIhB/MWjSVh1WaQKzjfrnqmwzODYsHs7p/8v7VuJj/f64BNqpwhl9FnUPLHCCdxsj
99SEI21dvcI84pH3yOqvcZSlFEjKj9DdTxuWDNKIi4cf2/ZA0mGag2qnSVHpMDZjnUaT+fSIfgbq
7xa7oKqQoFbv9czeLYxEYvzwQvptyn/ojjm8JeZ77aaHWbYw/aWvPlxxL1V3fp2ozAq2I4plfhQy
QfO68d4w3IpAQEAj7FfIkGyrbORE8ThDOIoe4VIP8j2A/+KT/Gr0TEGuwY4FC7Zfe5SGFZCSgl/n
GPBfwkM2QE5kCyPG5auaeRvg4bKMBOjwOfEcIAOc0NNvMoMwyWpWNmtDS5KPB9WRhBIBa47RLQS0
gZrkBO0xwOrEfgvIt5mKOKUNbd92zfHL+3ZRKJJ4vo8k2fmGSgGSmwlihuJ1Y1VHBsvq5zWpeiwr
DxfmStwQX+r+CEKy+a3YyBUzjc45qFnTQiXMVAO9o7AQ3a7ifQZ+dEpFL3iCZoSGgfTu8EauHftd
XaZL9WwKB+TRhz8JSXHKcs+alYyPN+tSKcNizDrZBxVJRxO4pLRCphMpu4AZIoG/BGzENZ7xs5Js
lPDirwKdRmzbN4R0MIm2Oft+snS8Y6iQWei2BFRFj3RyAG4+1FQqPCluQ5ql5M+wu4960JPRSwIE
xSrUEDZ4KE28h3oeRll9sR0temFcr8hm5UElU15lvgZ/lzovpAs4LzBmAv8PrTJNeZdntl57eXsl
jX9/R7893K7mhCQIhmdNG2QxUKHWjYF6X+bMpFsMeFRiKHXvqe860MkED3SpY3aybwncMvO/u6e/
+nFMZdnA8rTyhpV0uTsu/0MtNlqkFLizJN/Kiu3J6qy25yPp58CzU3dHfmmSKrwpa9ggDlZeQoN4
BBR2zQlR6mLCkYXSElla7ffDDFBqKIM1qLjwFUBU50o3Ts9Db4wMUt7IwSgDAVl1PxVC0HLA9N+J
E6JW2LT+mclm1bqukCFYKRk+2bNlO91KdtOvubxjEEy5fxKSmJx0cxKcJJmux8CIRu0zryDc0b7a
atiJvZW3QZBAG1FgLrqr3V0dnIQqBUP6W2VXSaCIuSJuBReIB+73iRlrwVhJPjbVZqDnQ2q1lHgz
4RAuramGU3ueZhEEqxil4yL78/M4zuG64zhfdj3wrjUaKgzDG7aq71Jnlx/h8WPz0Z9dmJEpaHDf
HXAgiblfFUOPK16uIldGE+/Hk9A61mV/vX/JzDX+nx7J3VSmQ44e1pmwku6BcdCLpY4/c/x46BHW
g3rCwSfp+AlO0cYGluNYY1OaRlMLMYu/Cimefp3NzojTrJZKM3sioyv/jdU+9cr5C/ZMdOWeW7mr
ZjARo29Uwi6V9MlyU68k4qwqi3ji8hUZ182JchImi/EHSdQAAK4/tVm2feL0ImUndxYKuzpHG1W5
YwPzUcRZ5bXzS5ulNn5mwKUKm8Mb907bPYzBqEFtivPP37dCS1Da6sKBLxAnDIOeDzZND9psaglg
oaEVPCj/lG5wrvHvK7KgfxDCMKhgwxwa8hxJ82J17J6llfY2+VX5jFanPrKi540yxKBW3N8gjHJv
JTAIA5vwpZr7iMvKs9ivcwNvghMRa/XVVXDd1gvUJpjKGaEByWiG+nzREj7W8Vq6V3Zt7ne8/hAy
fRYh3dQVhvCfHXyxCh87MZ3JRAkQ7EBSdXsRsl/gXECXZakADQ0DW500rrbVX+ynTn9v0fnCIDjg
3QmF9oehsb0Okdi3hHK75Tu/lgXPLUqQ22c6unUm+TOJdvvrjVe/ZkOq6GbmmAldypqhltB3GPP2
CiiK53XQfMvBlDe99hJjCucF6zLrCX9nd0I6h0IqoOUuUhM1DLeb6VC6vS99EBm8H+5GWv+DTrWI
XFhtJiODlqxllhM851yRjSRlFXhKDQC3FZA32b9e/Tj0L66kR+rKlltd0TGJdr2eWwdGZzSWJ7wZ
lR4hoKBy4OqhBBP/1WH6GkwDKRamt7XIuWqoGZIACBNhE/uI7ApSMmdSyA5NiBS/hNQD4IYr0We0
6PpxAQkNMCfv6Uq0WHIlHtbrmvDmelip97WZXWFchzA5fLT6OMojBK3h6zRoLVjsy/bYUmpKqM23
F4mZYqlnJybKu8an5C5tyC9/77artpKqMvIrYHBN2UW4mmccvjkZjuxHW4xsxzsHYCu0RcJjHube
CSyIHf5irp3oxCURIllH5Q2+U77BU6TNF+6ghN/JZ27jVd9ZndbtLRa3qDk1aZx3sI8otUhV2yMR
pCt5Irx6kotbix8zQH8g40lKYkrsN3AA5OxNfnV0Sp1oY4GigjUUwFINAvyDdvb1qKOHoPEwny9v
AnNp61KAESIyjuDZ/Zze7QlAq8+b2gl91MBw6nOdHh6L7duVjfFTPtOhGSeMX7oQJlEoXywooaPJ
28enZ/CXKGva2z/L/sx3ERJISyepOlcPCN2KMgmhe+QjTxEQeA//RR8+u1nIXEXv2sT1qshShBEG
txmzeUzutxHoKm/Q4NWEplPkrh2yxDzpOZ0xSBafB2n5i3Nqk/1jerzULb/W7MHSFZcEvjNQJ83K
eQmdSJtvFDN23fllKzJh5vOoDzFaTjYcCDCgiEX4+PEt5FIrVfjLU9vZfjqJSJLo76+FnJfSrF5M
guKPG9wqWAPQnQWNgryGVfR6fOn1A8kX35+vlESFqKF0KPEOGwxFPwlLzI6fmCPUb4gicmqbZiY+
ltGIsXKHRekEVMMIBTP8nLCGkngMphclkr5CQeY3Pcswl1zozzJdwO+vIHC40yJKvi32kD5PL8+x
NbXD3Tv6TGpmKu+T1EXOMMQ6ZrEJ5sVePHyUCqvO2+cHaXRXMdf55O62ZW7mbI42n+CMssUW7+9V
QEKkRsiZRPB9+WP7DYQvbebQwGoasd9EiJrKenXZPNWofnF7Qrb/7yiloem/f0z+hSfIZjRy5YX3
OHP9xrmm+rl8JX6R485fO+9ntbrgy6wL4XTds7qvQWNt1mjvcbPueA9LNhhS+6tustjoFmg50Wy9
xIgFf87uXS2Pa4A9aL3VPuhPJIyGFejsTRNWX58bBpwG3oAb2XEGohRXy+w4Lt6YVf84O6/wQsS/
2DW83iaFlw1fSQqqGw1tDJaplBadsaJ5E1f3j7jDdvBQk8ZTduPTybJey4Hn310q5JH7WfdEeG3O
ZTa7Rs/BY0FmVHP4wHo8PPVRWj1im600iVDP483eNjXFiRyKMjI2q1Gc0Cbns0FljK5CiyFSJyU9
mduyP1MJz826/i4Pd1S35A7tREst4Hkp4hpzjUp2p5f5pRlNyt7GmXSZQwElR+KqtGxZ+b4gSWxP
BAwQTfy6HgvUsO/0tC5r4Z87wki+dhE9m5fX/BxTUWShA+9j6X7tTgEuViSYCCxjX2hANjUVwKm3
TgVRVXqC0zUFrSbQd4WOYr63RV1BXLQV4GqoXHETx7XWfOY56tles40bL9WuPq2Cp11GvrUHUo2u
lLQy7VyuapUZjpxXDmF47pWvJIEfzBvZw1sOX/7nFzvPSNpNyIn3v+bzBuOe0F+T32NSNYOBNEQW
lyEGypWXF0Cq5yEXdnTX0Ny8ZNFpd/6piPf6QxOOGpT8W5dY2ho14rf9oACKtbo/ZGLEBCTwKmRq
iOxBVJYDozluZZSxOKyc0lVIdUBUOWoRzkuKL5W/d+02uIyEMlANOjQax4dWO5+yqB+spJalZGKy
JGXLG5ffRPelXUTeuq6FAFQS2Mf8n/L1BVmh4SFj8unKQf3Mw3scALrKVjlkMrNs9oVmlyOHroqq
V5RLV4Cx2Okf9WUPJfXdUcDN+Xt3wInyFGfSV06ioXj/8thnzgwu75W4A/SQ5ANGb7SobX4+9nN5
wR/7I90uaqZ5MFw2RDgOOh788p0n/cRaYV0iBDb0OSzRohcOzzB528wZriEZYqByhjTsG7v6V1Mk
wZPpb9tC8QBb+oDq21DVn6RSNV6WJM03vZwMeyIAUtVzKoYwRu2SwiISQi7GXIHse0AV8txG7o+j
hI62QTEJSFSrqfiBwIOvJ2BX8+0m0xfPvMDPAl6FFf4zi4txtjGnB+WcCgtMeTcucUFD29IolIKr
UuPz8w0Sth86Lj5Ffgkmd7c7n4O5kPZydWWQM3WGoINJ5ZdlYpBqZjB3KTWhKdWCxZWIh+kZD3Xe
833C+MC11R2MO99IBF7yR45je/tcF0qsezk6stQTrpfjN9NVdDIVDCRS/P00RG2etSg7klL8nsaY
2k51rgrSJhdVK/KAiRXc4jldKcbDo4AQ79V9NI0QbZSG3Y6pTwR9Tq5iQgt6944dUpYgbeB7Ar5n
iu8YVHk+aFJrw1eSiSeo2SSAyCpdzdRT4mc8ZQB/7JmERxEjPG+gOs8uGCNFuTnKcuYB96ojcCU4
oxa1mwL5fUjjpzdv3ntrBnaARo6fFB/URq595hCidhgs+dVERbJX8LJBhMpOr0ctDG/Iq02ro3EE
Fb6YufesQasNwCk8OGNfI2MUJowhPCHxodiiTvnyclmOtdYaNSbkyKJLcmLuOEFIDY++rDhsC0tc
LxtrAFIoFum8GyiMvNV1iCHd4/MYnCFoha+NVvj367NamqwVlfLFHNnW94NJO3YX4cf8DZHfDlDZ
P2o4E9jg/IPqdjFWfjMuIhKTsXkoF0aopslFfYWrw3j6pwglwNxt0uQxRhdNJ6URm9t2/eHjtGMT
mGn8XnYgRYx79IhUa3bN2U5ObsNmF4ygCnXqun0atUZSamrj0Ex0ae/EOn7AzbARkhquh9MTPID7
10dlhUW6DNwuFvevSBuQsta8Tf8r5Lb6rLPdlisoEePX67BYKNEDBA5oJGz6ieM65EEI9aenMMCi
mZ0zME7IqDfx1pCPHNUkMnUbDU4bySUzxvF38j5NkrVJR4WwRoOwe7cgyAwT69Z9sHcJCRMntlJM
Fn4y1H5a4b1i4FUEd1GfhI6dIzqzJ25hSoRn3FKiqkkYaWeiV6yHXtSiSi6gdLGsH1Q5tArxw6uf
orlA3LcomI56r3x1sSjpGU6DiMBPmh1Bm4hNGZKODrF6QLd6/uBQrTBWunVkjBm300AJNtRnsyOl
hCjDnrKtSe8bGxE/sLTwXo52ImRW8XFS7leHLh31q2JZjzus56N6iJvtXReA55oiRjHTg6HVkfPq
kX4Ba6QuBRDNL0qTovWXhWBxWZLJ8NAbwPnvUGlli6tzDFS75aKxNeBr2znoxVybDhq+3nKP091q
6ot3rTH4wIPdGACb10wf9/Jk9pcTSoJzSgwXof6Ao5/9Lz8nAQheGVrRs4QBgd5D/+Q5q7/JKHFc
Fel32k+BfrDWEedvcQD9lMOL7NImx5kVMn+RE42ns2Ci9N08WTBZDEx1nZBU3Ai5t3YwyaRvcAil
xvhKwjReuFLWKYp4ydqKjfbxoucUIEl0GqbBraw/oBJ1VfwBgDWogZvIeyzDk1agJDLYuIfw7Mr5
yRamSg9Df6sLZXt1RgaFukziVq7HjyucsUymwGgsOstUKxqZB9B+9L7a2QqlvEDyKZK5EOg7VzAt
IanyO9YqUfozpP07J6+DMqhG78ZlFPt/k+lkZpwNe5LZot7s25mZrw7yuEg2mpM68nfjIwcaFWV+
WSqFgmfl5XUvtKxJR8bah+fWlI0krU7+p/D3jtruZ/8teXdyEzXeKaLS45kw4KGkEo8N8RoccbOD
HdlW3EvcPU/kypnIrm6b/HR9M+Ee0kRpK4dmu9lOX6/iSS0Ihjnc15ZvD66pZsdN5QOBgMHqRLXo
4GNdrzjdIHdxuNkGMoA9g7fwe7zc5BFILb23t91Z0Q5EEGf6LNI4AsUEJeilctv2NA0Lj1Q/OVkw
IVRmBDh9V/I2Re/MzbDo044AEzxnbc6a70iOWPl3zKf6DJgt6IO7sqPsyD4JtN6u3pUX5Yzz0COl
9Yf6FBBtNspTuyGYMv1TL842FShFI4fOhu27sVFJpZYmuYyU9fDN/jhmNBC+XJTdxIJ+IKckOAqa
dj3IbN+GxdgrjjkdNxO7pjpB1C2onJQqkqDe/zeVcZku30+vSOsYWvKKqCfMYwX8Hfks2RGApRkK
bqAxy/sSyL9zFVw2Ji3QJn6CJVE5Dbb3LRnhmq1e8PNQm4zSiumbvQfuPgoQiIuyABmXMil4VBbZ
e0sS1pg+2jsdCxk8b7qRKrWvKplKqiT3Pa5qve8MThqmZudAu8OM5rwnuQEXMekh6GiY1S9NrT4o
3j4XHZOwTc76ejKqrRUPRIhcantwjxE2BFl8AK12F+pNqYHemN7wHzTXqQySwvsw+6qzWq1RApcy
fHWuL3xZnQ97mZkIYJmXA765YmfsJi67CBKec32hapeWIVYV9fYi9et/Yq53hxiXUI4CxjvQD4z8
iFk0dE69WOQrQBisSFJE79VbREDUwsj9sYjg4S+YoLmfIEhqnfRARjX0tfhgvZVbC2QgBPgxCdVy
4EH7vu7PqixgLS2CFUSqguuNihop7lTgVlzBWRHQ/KBG1l24GJUY406zWe6tARhiblVK9zfGxIZ4
VF8Zkgv148QrzAB9qY6bVu0orfsj/sET51ZQUGqCaW+KhzpoLiepfxmyim7fE1r5BvL31K0d96bD
R6sVpKWE6UP+8GtSKailQFJKUPJDh1Mbh49hOfCUcZFUkH0sBHut5nNLumo11xa13V0j0nkhtLXT
TespbYHWOHjkR3iReCRVFTylFl9WwANGkDUecQxrHDRR2plLjvcvgkBtYjkQdIyFwVXGvIliRRoq
FU2iSYJoisqVxPuX2NWiiFIrV5o5PN5KZthlt9oj7ZEunydcjIbAN9e/FIXjcCyLvLoYDlUv65uZ
Fv31mfr4wTulTwAqwtAMd4zK8sQEA8tbYAAlEq4zMceonhD3eGeA761Z8/He9ywNWsn1Kmg7XyyQ
GPodjgQi6lYGlFAVRTy1rLsLdEEJFSO7XvWNWT11iup8DzkYPMmVXRYHs6dpm2+0EVueWes7hZNS
+z4T6kEEz+DgZyZqq8WX2z5Wd1AhuJTQspJbXk2GN1UE6h5kgtNz1hPAgvYA1cOSQbzCqL2ECnUl
AxgHs4Vt1zp4HIB76Em1p4KWkQ0kL38VykD1PzdgUQGmE5Z33kxJ/2I6SayIXadNtV3ATSbzgPDx
jlY9QtMzvadf4RGPiYqV5MuH8+soj8CjQW3IbFmYZRYV+Z7/0ZuGgY+SwN3kPvOioAV+bEQwKlVH
oBDMuRaEz3sYYII54nKWZguN/uXtx7LHYoTbs0Z6lNHTQKFFf8wEYTcr8TaCj5CmIBmK5D3Pc2s9
2mI3Vhbn/WQYDAHJf1Y3S700Tr57eGLm9BGtlFJfLLdV6pe3hChovTmdnZSskQGVpPx2nVfowsXM
zrpGoTWn+kkRjUGRTqCUFJRyWjakPKaCCW7UW9vTaTO7iZRH7+t64RnylAN5nihIbhI8O/57eZt4
X6xyJwjkZQsjCqyA4X4ZH93VvEZahbv9KLh8z6oGx+pq8ewYhSt/Tt7LZo7M7pSu9AWr9Z/KpMz/
62F9r9yzeq1FllU/wqztlBqWZXynI/csfckbZt7OhiW+X6jUmADWq6lM+Vv6nSV7rstPLKcLx5/+
R172g/H9F7RPA1QOSCmg/6HsaPvO0hqMaq9YA52/ysxcjfb3qYMaydY6VktGU5MXnNrEFLTKk23V
CxYcDH8BiV0RCu8JDlKzp2XzICx1cRM5atdMHKSYkgSd4N5m5ZRMNCSp/9XMfXeG/0uSjXcvxNAn
8ou6w3tW8C0nfp6Zpo20/A1K7tYCxP4MhLU3jZzUniOxe2S/qrKksWhbzotuAiW1SWfDBnDnt5s1
jAuu2vb3T9BVE5mGEJEh3787aE2U7GrSxhJrPzLm/quZRVI587eoacOzOF040E4UNiwULl3yxfxR
BSh8ot8UyRa33xEt/tZR1oLON/GLcHqeLTQPNcTWdlzr3YsPBuOVtVdrkfPp9eb020yG8STXiwUf
LNNrudrXhdEx99kyg1Wi8T2zeHT5nzbRhaS0avq7tgqLo9n6g+mAMVy2tGLldIhkdOHGQrSn7/mL
e1yu51wQ8KNxJpKVK9wi+Fczk+ouj6dcBZWmB08J4Q/8Cc0safGw1iZBkQ7kSaMFbkNYmzKgoygl
fh0DQN3QpU7SW/cw5GYfbPhV1sUwjH1ESlRrZhlTcQp1uJRQeVbaUqNQsomAsrnLEMevR5wx/wVw
xhmWvLIRhIurDIdzq+IKLQtrOpsenOb6ZXpsOajbFgH4XqBsT83trEzFGL04Ym7v43TQ3KWGCTW7
t3x/VjUuTrzE+YROaKO8YONpLhAL9xe7DEiXFl+iAFbt6xr+wO3ZZXA+5mvv6+JgK7wyM5l1R7KJ
PRGfretBH1evB9pCdUX34U5JU1XNaeINFL/GmXRq8TvoTnMA5T5ZN/cScVK3+EZJ4NQ1cJZcuoJh
C+kiji0dPDbQ5DKHCRZCfB1V5+awGf8MUql7PfoSl6V1EAzQUdLfNvP/RVUOBhAQB5cfcR4jE7s5
V84WLdo9v9xTxjfBUZcHRufnBdBu+ye03XWWQnftbhbJmWnazLK+hxkVbDnr8yPdKLLKXyRw2GvW
c2M0cAaJXjfkHty1TkjNn8ZM33eAPJ42WERd6MbpxEYlh2XHBnFd5H81wAt0ElTr/V3x7PcWfCSg
w8/eueM3NDyINqDss4mtQR3E2tjhomJxweKNeN2wVqaQT1lnVFM665HHi1v5xTYOiXWqXU1HOp4i
w78w+BQiI7UbgOrp7anJVQkK6BYURHnfqUK0JFw6JwbCUFz4R37YDobmDWDlH5Iv3Aiz9ThQse2H
wMQoBFD955Dob9WS8JbwMN4MJ2u9xI3W19sKoRCoxGdQ4lwUav21/QACRWEIRuDsTqiUbAq1kj+P
MClOKmbGC3t3vs2rKMRqRc5o9/EI2w5zuO80dOlmLiza5mt4NCFTIybitRYvO55mb2Jjc52Adahs
mwX3dBp3X4MA1twBdUusDWpGfapwuYCkdOFTx4yNSvKN8Y9PDyX+Sq6I/6TFZp6ewkXBZWlTLgrz
fu3zPJgC+spqFyyvHBSmGkiZ2y+MyOV6mTgS9UPZiA+h03ljb2WoXY1OGdrTGt8E1dqccd+JYMIs
n63vVPNVBRf4lDWdxm/w9JLzbpvq8p4Hu6xctywJC4iUmkdaSxHD5CIfW1mcrw8sT+dGatU5Ezp3
5a8ET5sGebus3OQQ0EUvlMz6I/kdBu4DUGWdTmhBCTBPgXgBr3dtBooXv2/tl0JSV4dZxCNpD6Us
IaZMaY63E6lXhAiCxsta6TSlFNjf5ge4w98uGWZaLjiHq+pz0K/JdzcyT6XETIjzLkMYMlYKzk1Y
AaWjA6r5xWTupb9omcW/pp3vF/Rm6VWxz10jLBwPiRQ3ppNhLiSWqIusUVUNi4XtvO4FndF5BZdB
O30KEldliFcopjJiiVKsSIoExo44P/UiDjtW2LimRuvrRhjEWBL0QEv810hGBSYUZ7ZLfqdyz+zJ
YTKu0EEvdX3dRSCTHLYBBQUEEo6PSpFVjqmp+WNMC1eJzHg8h3tnT8Yf3RrmgMwBQ+o8m35gOLsS
IKuL5crx4yEYuAXRY9lCWlm3/L042kcucc8BZdUKoEo9R5K9n+PrS5BkMB9CECo1URNxZGmOWUEg
zmgyRrl2sGTPDg7mmGJ86uyeUyYISzq6eLOl8QhT8vDF5Mv4atddyRjRt1vm4pt2SfQYtiE7s2AA
T2AFIQCH5Unit3t0nl2fr1HG/oVcFcqkiFaO7EaGTAmCILgpbfp3lfADaPekuyhnXFPfSKzsIAxa
0c9Uo+kAIkesbGO35ZklSHI4dq7kw5v4BEBuD+XMVWKZ0z90Q0sluxBRFj8pHLxyo7XYzJZf8kyU
1IzaaSSv8ZOrZG+XTQOFisutESjCL1mvAfLRrPw4Qn1EKE5Erq6WfKeF0NlmQgh3mlRIbRqDCzL0
28rk6v6nBNqxy4oi77P4T++kXGpi7ceqGi3MEAgNzuL9hgeN48Q6l1f45GGtzMvmmr/YtxQZA34S
fhr3PeYa66dOS10XpccriocF962aTgCL1fl8vH92epFxRhABX6r4q/9PnmP+cVfd4HDtF7WMvTe9
RigcJBVq5Cy8O4Y54Jd01dJt04gYRVIS0DKpffE+UIVLV2znY9uiE9uhn9/+GKGDu0V+slBwEuSO
o17MTzDqt1HwAWru6AIwb4YrKw+DeGnIqktigWiDFRiipY+ATlfbNpLCuNPk/ytzPBhON59+eeQ6
4QV8XU9g/slDEFRvh1C0u8mF9kuIkS5rZWjWM2kBIZkLPvZ+1lIxDAR1fzjH3NThTCQhezfthhRF
4zSbdMmPAMOO4rB7xr8uHRVUy2GpPl+EbWMA+U7P4wVjQAangzHJeYp5qix0cVW8cQfjRcrVrx4I
9iQJMWQcbheSYyQN6KqnXicNBUvPb92WmZTXA+cj2x8WkT2qVsFtt6Hr8QftJIcQ7m/DqD/n7Y9z
GApYsViDQUzLt8DjmtS22mpx9O3L9Rm8VKyWNanej/Tj9/XRnSMZPvBVr69J8JWyPu5fW5ksDIaV
98lCp5NP0C5GGCjoWX/k+8DTYQaJxy2bXRMC1TTv7lgMhLLZW/lwzqSK+5xRQYGaoDDA/Y04oqLH
hhr1noWIuRcN36wFdb99nv5Enyufv+J8POLZuWpctPPhjKXAqGBvI5xLFtNFVHqIPTMpoVeqlvg1
Q/h6GIoKIVU4tsuvvWaVx2Xu++WU8iaHv8vfPGDjheRGKM76Zn5P6oLDnErM5HSeN0xP+pasMkiA
HqDwA/khZDatC5BInmHxPEhWtmnZtRmsdbN9LerVkZuZDjznnGe67K47Knxs3vOac3MCO5UyNl7m
Gr8Iy84XNNX8fnL+MzeiChTc7FP1j7YYmN2V3ZDj3uVNXc5JktNskW2979lDITJjWGHbzF93Zlkh
cSmsZstc+SCa44WvS8QyosVbfdIz8MyyLnQxqFqpL61fb4d1KtVC4j/hApSrR94E/Sjjb60anVz/
l36xaJM4cY6MpDFxk7buYuTP1NAu01vlOM09OQO7W2wteEIOgen8JcgPSm/6TvCQTYgWl7widxks
2wzlKS1mlpqfVsw9h3IrVtcWPcN5C3L9jRYkfwzdFiA2rBLE6DhjPrbFTVbGo1VIZwhVOJycMiOs
Xu8YU0Aej/aNLGBT4CzSc4mnHClGYErDX3Iim84xhuO2Hrz8SL39spJ2aXDFdgdbT00ng9MK8Tt5
V6qpMC8cYyDOnZY3N+S839/YyQgx8h5tXXmlPw4KBSlpF+ycFtdk8wqdCxLnMltVrWoUcdkAIFvS
GSdPiTxOK7Zd5gi9T3Aa+dUwIqLyWfSp7tknjkm+0dSbWibWqDq9a5GUSA1y1OUjN6373uuy5jAX
Wt3Eia49MGfUuBwJfEFFvkn0Lc4CFyIug/QAoin+SLpyr8BYFhZPML3QJH1NTwrhuSk+QlykA9NB
fIjt2+ih5UNw9bXZEA0tuciQMz4Ww2sKiFQhQDqotyVPuO4mV3I+2Xil0PvT+dyOhRW3PybsrGFy
/Se21yQHO2Vwe7jLyQdOhzbsqgGeAPqKqNJ+tgbYwQPn9DDonaO3TuDGvjvNRD/E2XIA5JKiMrEd
My9b9zHzVjEQiMzVhL9foNaVVrVn9wEi+J7/kJ55RrQXnfdYin3SiGqGp3lEggwK5LUX6tBZEBaH
7e5MEsT/FS9vKGfBhsguhMbHOEr2weMuBv1s9qRydiGhpWEBua7OVPQ42RxblKMAd7zjsjNjj6x4
ozVuhFuS6M+SZYTJ8JyPBDZtBk07nJjWV8kz4HSSKjiFGFl9BAuHvp3s1pW8xHRDJaDN/x2UPQqx
GZ6Fj1vn/erenJB+sYjyn95+ku40m8o0wW5Gm0LU1dTyyxJBQwUaTy5ne+779Xg02cRM85CVoxNS
0QGA6QQn+XQVjjVCk1YP1fcddo9BNiMfp3b/bW0VyJILxJjGdWdnAw1apW+X81zIxu8vgl7d5lqy
5NvWp1VTa8ytajo5xyNE56gf+i/5rqCbP8B7rRyvsSRt7scezSfwF3rs0XEpTr9gKTeaDKFYGuZg
4i+htdvQ5hoy60qphmC0tYKPUrfDVq+nKmoOudjK5bxamuqX1VEZXgZIoEw58cwk5Zlifke9OerA
ObMYjZJFrQcs3vXfnCUdRWJKXqxPJeuIbXKFdQwXsQe3j3r4xLMo+scf+tqp8D1X21arQMGMZ1li
oIyP8Gddm9OCEkovLr/Is5McraoFtfdn6IRKmShTu8kwnFLVuzNNNMeuntG2C13jFVqOex/DHmg5
slpkEcCB6VV35ZjdURc+TROJhVSbWXNgGEvO+v/T9M0MIizUjTmJp6rOpGrzMjXwMuLLDLOs7b+D
epQCAoNvoo2eMZkrW2z9PltpzDyk02/J/OywAqTcFCdzaHuKqeE5EBTZxKmFDIvPila4Bck1pV6U
G2qin7fnaxKO1V7ox6DLWR7JkuZGL7uNVLGQVwFcIl+UnFEVx/RX3TlytSxf51udTC/SqS8jzSB6
6na1iCxHkhcVoZK3ExLMBXlTzMIpMdephLd+UBu2n9DJr4yy6YZJtV1sow7O4l0/1J1HUz1S8pHo
hJ8/Jcqi1ikI+FLz+foe60NT6Ednoc9gvCYpQ+3xxC/l8+yv4iSEyquNmRjSB+sbjtViw5B1MkSA
8xWXXsrFM+vrmjsGbJ5acKUmviFCNqBHW87EGtjy2cHVgKpUHj7m8SW81Cln66l+6S63qmBebwIJ
1SKN04j27GztQ6kGMuQu4O1YhXInhxXsgC9YcASMOb1XKEN75RC8Irrdoq8naDYBnhnK0jC//aGr
CO7jpK3Asm1p7ALxopMSjT8oQ73Red1leZyO4iMBICd39HAZeNa1VlMcZilK3ZvadqFz8jPEfgmU
TsfhbOV5g3fRDtA0zdOqDqUwULyl/z0ALn0ZHSwYDLaftY6n6+Vq8zrbmPma92zAsL4CcZEgKxNn
VY8G7mEaY72g+ahl16uw0YKekBRD09aLAXy72RWMvqsdOHXFTXbJcswAxr+8OC5kkMQBAPycRSPL
FDgTtZdv38u37I69NLL9tpf/csOWvQaLr+I5xINXo+Ro97rC+fUv8rgy+fu6jTMnhdesxU2VYxts
3hmq95pkg95F9KQu6bxvi/THs/g8bXV4owzRvNILrqRjvmfKDiRj2NyVUhrFgZhntI+haovJMavb
fd9pNhWCEoScobm7TPWEzlgp2/DostTHQ3fzNNa8w3UrSSMxJx7bireJxHrWU6WvjDt8ddePU54B
iIFqHKt7Ku2dzgvKW1VLoUAbAqoG8JuuYbUCX55j6PUb3LjyNAeoIEOZuT5Jek97/TTWiciSCdu+
XaYY+fuhb67IBs/OTK0wRl8Ltg6PJeuEhUXAQYvlPrmAqssjDEWd7mugI7usvg/42b8QsALWQ4G0
nJJhYB7QOxstRCC7pRjRjmL4Fh3KcEtKXcOYXoS4fJ8f7M+Xo0V71dfoY0b7pLqq6nEnBFbXaRxi
t0sJmNPSdHZKXVjsAEugOQ73fCm+H5qBKaCHkhBfEcf8szxoJVVLicibQnPdZPtMv7K1/RoWpmZ6
XRwlhaKIkIf2IuBpvSr7xppRXK3qr+ayj6lav0KJZFntoyBGDyRYckZZCr2LwX01RrboaJDedHt0
2SfUoJJrrUOnFc0xQBc59Qr0MvM/rSmRHbE9yJHeWNZReHvIsUIdfdq/xe75bUQHBwaG5uDFE0zO
D+ePSm9nqS6ZPVES1YMewYhacCCT1ALfqDgAFDJ3IdOANe8Jy3YmkU3he9+rOG3fhUtqY9ihg3pr
UwtwSPvnB785pse6TQ8SuKqI2IAaFXe04zuUUNOjZnqX4CRMhIsE55UW4btfO1/U9gX6iUyH/oZx
E8nT8HQH4VRWjyq8FYld4IGJjptTF+orLR5CbV2YHXOSo+Cg/AkKgwY6L3h5FNxhZJfzZ6WYjKyM
ZF8DrFZ9pvzkjdEsjaGJdk8csebWgRpI7GxIPe/3TrVK83UBSUBArxcSK0s0KR1oqncDI0HdQFs3
Uj+DNd5UduPjMMEg320qVrqCBs2Ik1k9ZopiIMtkh47cpdt9KM7xBXeCigoCMlvM+nLcsarMQu68
QL4rlyS5XGLZeIxP1PPFx9JRPnn66BKYR1Gkemq0LeKdOqOc08cu63p+gW3fp/PvpB8Y5EdOxrWb
arrgUaVxpElhXxBPYEiJfzOfKe89SQOwxO4eQOntByI0HbJ00rTCKuj5QY2JgjTdjP8qg9q30tll
VhOb1V4h36bX3uyi9g9vXGuPW0YVwyrSK+3adlpSrfW68m514RiaGKhYCPns5AFMp8Z60e4TMZJf
gD7Vp2ynSf8oh0b8jYAsF8Z/gCPUn/2aOVq4gyExhu4vM82oJiFn2tYfOAxmoqtEvwLNnBwD5OYM
mho4/0LWGBW2jQZS6EA+mShIz4nPpHHZ+rN0Y1FHVRzvIuuNIdbG2rDvAw7FgEZxUFIP4XI3XhIx
PumWe5oP/n90K4dVtMyb57Xznp+xYNoiIZyJKtKDmTCAGvhXNdOuUkRbVk2+fGvdt7LZrNwW3zD3
gj7FI1m0ylzNIH7RDGW8flQ/i6Bp8NekhaIa3MLLWEWcH0sCshHZOS8i9ZquufiIHc03I7ZCiR4Y
qvvAou39VuaRdNXfz3hkQSI/edGr0Upzr6bd4DNSfoi1uXbJH5ZsIyeVkDuwIZad03vbKQn0O8EV
rmxUeww2vVQRcz86Ul7j3X2bc3bLD/pPiCaZKlkueS19FaA6UBuQgTDU5ePayCwTh+IK4RHfE7xh
jFf2npsymeWfyR2sgRLe4nNdrtEUonwKxb7f7YAVNM81cD+vIh6lwIVGSr1WPYJg8ieCGhLayVqT
SrhD8fp/dkt1/1aayD9smax/qV9r1LnqazjftQhwvV5eHqZac2fydrGD2ckZcXV0wlVYAgBZNn80
MkU/Iz2LOE3TUSS57EnwkuooBHbdYLins/R9jrZzVj4IQtY9ZdJxzDSP2ZT+5s3cSl8LEi09x0AA
/JBxFSllb0rtgeG6ADnB9knqztQbvz/eYNVR5DhQbQTJzsHVfI5UwD6ITupk86WXnDguPp69oHEg
vkIzZvY5FfpCHtzKbH5/Gjlka+IqNLVwtmI7wQQLArqD95ybzIExru142WcIVbR7BW/AYuagXWvC
9BnUnB8/NRacjiSPrdL1NGwxgar0jBqtuxm5qTGFEolUF9S8MUXxmeR8VKbHwRcgap5pZ6Zz6MKS
wybjzPvVceH7nL/wobFcbMIPWajInysTjs23A4cg6qt2rk2DHe8adkZNSHbcow7WP3SDMA+exJ/W
GKB2C6f9o7oWU0jrcUUbqJO4I8LlXl94092ejzVOBtif1AmjAcQHP5M3hpbbJFXZaBLnaKWaY0dI
j9e5yUabJA8yZbdL32RAwyzmb1oK89foXTzQBYHci+V83cIiOY09heVIGHiY4pUrC+o8GHEJKA3V
7A2nwbIKftlGPcqIOtOO2TOfQiK/QlYIBOiXseoUYTjIopEVGv11rFA6yQuzYsnCSQdxaCULf7y2
yrp5M+wK6NJKmKj6RlvHOHa5/05Hg1KK/hT48FNQl9dtY4WNo8rVEXInzAgTeJodiZdRSXc8tcye
Jh3xyFQPDF+PLHpJ46HOhBUtrqliBQTsalZP6djOvdWNiUMgVgdeIau/k5hPx14u/803cBAKO3gy
/NXNOoq/Bh0HLUXAhPyteAYv4Wb8fD0PoqSH3LoLS4OQfnPkXnfalfxzScdVCuWsSrNvqNfs4RJl
xzBYlzMe3uKRwymXqXh1DVAL+Ahc3b4Z2fhQO7gQVtAAbU/gXNAUH0w3bRl7eOKoh3Jba7Gr7YzS
+2+b6O6Oj/WXdC3AaTbN4EPKus2Fbv1hOrlYs1Q8ZnYMCT6iXfNQueG8DX/UxIkummWV/9djyYcn
aJ0MKAAJFvG8IusvPez+fGLy/ACBuKSrXJsNAq7I7E2hZ6ya0V6Ew0HuynYXVQ/Iubf17ECVcpDh
thkoWcsya8qMyU+mK1PlUa9P9zHzH8JqqNcMYhLSeXrgOgkGq4XLYUOBvglG0M/AlxKyl9kPA3lm
WWn0xsRXP0v9/6XU3KnYvJq+/hc66Vi0eCoQkTHT5OO9CS4OYkb4W1NHvLL1Nss1ZSK08CDFg1uI
2G1CbuIFFeNfDNDUlrmNVb5fLlJhYjC3ouU/ZI8MWxD553FQuPAj1tk/ACBeoKoFflH4UbVNCXP9
VKZ74W/a1znpjZm+wZ8Kt9JHyh8rVgBOavCF/GMB95C1dr0XOyr86QDXrm0SMewHk1R6l24nR888
71zsi5Qu9uwo1l8IaSfNdDPgpXrVbovXslJVhiviyJtkZexIIX5nJz2ZlIRA9HGlTPj2MQGTiHwH
t490VK5D2LmKJP6Qvhy5c5lcWLn6y2VGAUUvM/Sv+ekPC8a9ScAhgqjznzqKQIpIc/0YVfFsB85b
L3NQyWzHxJiwnw5gOR/ifoxOcIYRRQVMjpdAjxg4BjSZF+5Rf67oWpnpHdyCDCXFh2e6rUGINvkj
dTV6Fi1p0ql1vuiZ7AHoAWb/xGDIEKeduMfwuDH+jkj8cROVxcHPh8nhqOEhyqkF9IyvFskaIvjd
gfxIDtOzzocdVX6kiFRFVV2h77sInYx/N2h0Es8THo4XMK97I+tQTqUtwxJ2Eore0ey25nBZzih8
yBrXc8g/ZM5zqh2qR2xekdFteeWUqFbwFvyWiGy53+3YjLgqdVBThFIRVeFeyorigvu4CtP8mOK6
BrxaqdkiRJDo/uHAhISGF4U7O5rkIR74c6UknqyZvriIZ3oGceBFsyeYrmqvv7pwLaZm+/WBXfeG
4VXwUPHWAgGg3RvkVr4ub1FWrcz9Q/27l06OfycU7/HJKSxqLG2vvraWAE12y5t4vqb8Pmz0NXA3
Yop0IKX9ZL63Us6vcPZ2CxalIItH1LJOe/+FDNp/Kk2JE88DRgq8ws6dU8RljO7ctvDC8HDJCl+4
NyFBgKurrkIBMaUeSnuvFPP/TTwH8Kk9mbNb4DHwH0vuNZRcI5MPy4MQpx8KVPmAeHTdu2gGeGWz
Ou06N48yFDB1wVcw16PAbaP8uKSXjfG0TD7ahpFiaz1PsZnRGiRP3D+2u+mvRudNGwXxnPrM0XbP
gmsB/Vp1F3fLMVaO0ijLy4GoaXldrhMiIm7ypQwxT4IUEmJyoPG3G2tifA0383P+ZvZnY2iQtPLW
3XO+IeqhsbiLGedqD6h5D9yez2gcVRqgYCEPPVrtdky6jlCdmTO/8ljpRAAn8bx9DVnZr70C9F1c
1Yqn5p0qX30nm2eAxP2O7g0O5kRFQMyjvNddpXwSVYoj+xE2qxI0QO+A347pF+7ZJIQ0m0CqClQG
CrTYJKGAXljERPTTxcHtbw5MnNPhC18JG1faFqA5/hH8/l7bpt4CwmY/qwZ8lVOxZMjLBNQSv8lx
0R1y1MxUAYPj5RQ1Mqa0KsQVvC+4J0Z/wsVnd5ruZX7swhODEkwyU0UOmiN23ec7OZEOQ295TGW1
ZlT10bMZ2u+LHpnA1xuqkmvvIo0DuIwnqXwBXzBKCizNqthj3H5Z0thBYQeZt2cRW2gC+g4+NK0X
vtR/SbnrCaLmsUroNbn9WQvvVLnVppU9MwimDvROE2DyeNScybfwcb+D5qhU2wt+96/uHRj8ZHEw
AgjfH2khrF48d3qCNxnYiuNOyoUxvWDSpXG0CG2NSJat07+FSeX3qBa8c+ueQzNrVg932p2lDhoR
AlgGJH9qEEroMu2fUsqaAeIkR4k/MqJPucz6sy0ARUtrQNny8oqiUpQBTMcRuwmiMc4Q9dagOgz4
p6R7Q1Tl+RkWaD4vVbRmYVIIiEb37I3Bj3topKd0zbEcZOk0YS+vB4+62OY0a5BCdF5haRX4DsDU
KkteCQMkrZu33OPWFpoKNSlm+K4DjhY0gzTlTrwNPqDaO5Upa9LhLSUkM8Dg/0tEJTd2E10dvFOe
LgiPtXuMmLPs6EA0euZZTchIt6ap7INUjAsxXM8AkRwiOYjdPq92IPcMBpMTDVv/NvWwIv8LACtS
dxBmN9RKX0S+U0zbn+9xCNfQ6sgrlYSeF+KwBUffTdW1SZ0QjW2iTihVdpQwxNHwbzmljKeBxBgP
gRjPXUlLIBwLkXeInIcHL1JE8bPxtjYyzu7Ni+irM7hq/pVfyMwI4fq7kb4ObJ+g+pTHWndMVSd+
u1eBolhWN9LH9AD5ETWsBH5hdaAil6LYW8XbYgGx4+L72SfFnnbW+JYzy14UIoRnmOtz3CTV+waq
BD+3NU2czmvwuqh9P1ADI1tvhBro5pYyjzfEZB3hnE2JZVHYu1/pkR6IG2PEAPAaVFARrXZRhFmY
0Us5SBRp9iibL5zGVZsrpiXXj9RIPiDmrAxl5GjzKXdbczp5RTK25iifypy8f8ygCTTWlUGTKMEp
zYNI0PyKTvrVvvLuUrDdEOhFccpq5x3ycUcVK2l4lE/yBYj9RVPba5IyHSEXnsSZ5Mxr6jOWIhH4
+V5KhvI6qpwHBPTROSYLPkX6l2cMkZbzBfQiUM1AuVgDHRloVK8pyvDmc5ZZhm5bw0KFdEhZBpx/
oaGVW4QVH47tAZxiFFVxeWNepvnAU8hJowL69kW+ulxflC0mj34x9w/7DZis4I6AqoXbvKjrdmlG
6Z3a7zm9Iw7Fs8upyKmwzjq3z/UZweKjhlzbBNUy20N5N57k9VZcsx1SNtspzsU+ykVI1mCMHNRN
I9dLzzZa+UG7LnPyOZ4XuwalVohjNN898G5icQ3fp/rcBtsNWQc8BC2DdHXuIBBV84iKD+fvVyPi
gwawB3lH5PZlAKFCoA2X0GlRLZUtSr6DuN7ffqHvo5DU8V9RRe/iT6Pc/HcQDbphvLdBzUisi9fo
/V5O6fkyBGdyQbPbFC/yvtviEQk5ULqhXYPELtoS05AnUfGvrg02uz6afYWya7+EU1QujMhp+BrR
2G4AzQNA2ORpE7x4hmfV7fcs+4T8MhGQUNfmYEqQtdD6Q8LU92qd0ohwCZDY+au9AQWkNyXAMXx2
eAMdpEhThe0ISfWYZ6ycuQWBryq/96M0wezYDqy+cVMnylHjtyH0oYeYvh7G2pLI4eUsAp9hS+ME
RAo7RKsTsbbZuyLxRvbCKhtHzBpdlRkD5n7O4OY/X0aL/ZD2TVfLrcY48ZsJdLnKnoHmBXLR690u
MvwAr+WRCo2YPaMbP5oNDB3NMaqzHn/QJxwZjY4wSv+axs2MGP/WrKZENJtRLf6/WoxcUWJs+8DT
DKfGWjpI7Opf9O2PlWDsVwkRwXVrdwoGa+7vU6t98RcuICJAPZ72YERzgrOX2B0hfeh44p1mETBR
aDzy7TtH/ObAQKVOP5Pzqf/PVsZ7J87BSnFrFObveuHOayrp0km2ali8+PVM77cElKUAUWnLCTQP
p3LalY72e6esSgSDguYQuLAfIKAPT5jml+UjiG5v3um5mSwWb1xA3bk7KI5LDnPdGS67Va+Qsufd
yuRcLKHqO/5jllXlgA77AflEw4mqFpxbOyBzsjhjNaHv0PMHi1IetgVy+ggLCU5CfCVeR2BzP0AF
mrPLYt0pwJyuAxXaSMjp2s1NLUzWC7g4eIT9XdaramwxltM0NIS3txYBlWYct6+rg9hlSo+u/OiG
7Ovq2gOz2izmIs61JRQ6CB6Pxhxj9umkM7IyxBlZ+3YFIukiqpsK/aOeN8y6h1qK1ZeqBIo6HyLF
VVLE6wWpVSWJ8GY/gL2OwT8t203aIV7gC+dIoKFCcbp+SpMhR1iu7cPh9bVgQKaxZciNWN8+VaLX
XkFO6wP6uOz0dEogFL+aXYJe4714RtKmn72oJr2aQyf/YuBttzVkR+6x1/JsuHDk9tpxF61Wv85n
i9YdLvYoAM9c/HItssef1YBLRMV4ANyVlO3XXbAQGoB5lNvSYzoU9rIgjPV5labWo5l5BNNemOme
Yk+a7wawojpHDaznAqSO5NOiRVaKdQjcjPa8YjBteqd77VPeWc+0eWWMBAblpMF07L06qnQhLBaU
+MDBVs2CJGfWjnPNv/0SkSzTL+YKMT5ednLXS6pwrn85pYUM4xcyJftt5zYn7C6p/9HINe1RfuDY
gAeQT8fN5tcuZm24g0N7RsQmhKn5Zv/p6F6DOQrPO9fZg5+1eXf+cp5IgP+PeVybBfSXEySBgMTD
D1R6uByNQUFh68Tr9JAynsnnty1EaxUerxfU2ol6u4WY36ghFokTUaMeCkTXfPq6zcTs+5Ka9x5k
M19vHQgaYKk0ujT6jLQOh22eYhZmxaX7D6ZSsYoYtmrBvc0v7/XvMNf4pe65I7g+584iCII3ojnj
cOlMeIoAZV0ZJS1LQ0uO5u/cilblfIyMGcGKOADzGl2Wjf65YrWRINqKb1ZAnnObS+RJfUallOUW
/pbGkMgX0ym3gQ7Ol6tH+OIK1A4dCcD277A9cvDzcP7aF27wt9s7GabcDLs+xRvQLlACqzv/udnZ
7jJDCu4a+EaMXXyBTNonTG6DYVY4oKGdxF5Zp5aD7emdVDq50TW0lBjJv/bjzxxbDdZH6mHSZxPv
UbWhrypQLFqggqN7RPvsrrw6yaFuslaDs1Sl6mSgdfu3sE5+vucNt0XNg6XR5axdoWr2YAf4mQYB
PmUkXf0mv2xj0D2v44PnME/GcwjAxX/dd/h0A7yRlMKjohgzZVb8V1Q9kxRPPE2ilx2JrXI/TpHT
p+ZQEun0Yom1dos6olpPpjkiklmOjNPvqlzAIh/nadttN/623HdOxft6DZz27njQgMRgeQMLaIe+
RoksQdfj/CoJ6HBCHY+GgmbGO+OxtYyyXVDEKz6FrIWqYmlMiVQMjALg9cSsLkhkdybywpzmak7f
AbN/M/KRbbBy+SyvnFbshLg2ycVDQ9NJIZiSrlT0Bxu+QKd1Y3WtWGoNy9KPUE8UR8jbBwOmSeM0
IDjU5qL411Jfw7nhy147Y6PU6+H/NhfbZLTFHJho3A89qUb2yo/bVUwRD/gn2phzghgSU/Qk11HN
0FvIXm9OLGxCN11KrMtwFUDeg4Ae3ArjxOq8+cSV+Egbs6WafuD3U3WS+tRfK9iueeHnsTYsKSUe
FQyRIGdoGfreTghUbefQpw29B8hc8Fx045CWv3SHMve794I0N69fm+bcNECCn8sb1N0YmJqvQ44o
O3INSs8G+4jMXckiih2tZDUGnyMwnpzreihxhJswqdtYSDszlIGmE0yL7QAw0mSmtwnx2KaZMzQH
S3xxSmpPfU6ms8CWhIS1vVkb6Ota/xZZHV7CLkWaBgwp2dlIldISVjsCQucHI4DhukjsiDsm766J
IB1q5oh2AmonJ/LANB//vPji6v66BPdJdj+rmVxptk5OeazLI5rvDyJD06sjfaYagHiydoqvfpg3
TeDVGMVDE5RLHDUcKg+W0S1paAQFrU/34atH92GEh8urueZFvENl61vkQhnSFqGoFj84dbwXsSq8
rCfH+DsJNZtjkEGi8pBXY1srunrPy2+jEXyqIdC1iHLzgpwYmY5xIahLcv6BDBovb1idvJrbZsZL
5GnjHhFe2tlC0hJqu3NDMRvwu7nwQqIw/dFDlNYSVBurUqgSHWn0iggdLUjcuhW0nFV3I+iXCsEm
yz9iq/KfKokJm3FPrhvLQ9zpcZ1ffyB5u5sT5J3fgJXCzFZWddj8YDRufLnW5CFBbUzPkxBDCq7i
k1MMwRHEF3K05ACa/D5tqAwtoBPUOr5yajowoyvppP38I2XsnLiILZNMRjro97gJOgP5JoYNKkHj
ikQ1aGd1njbN3sw7pH/Mxb+yQLG6T9ZprXKv8eoJf1sQRNc3pfoJxPjYZJd81Y4hVR02eHB9HK41
tr6uqBAZ1v8pFI8xCRnYgcKzwyxEyoS/Hk+8dUYRcWDxpJVkVVRk99++SbW3Liy+nTSRPNzQ/23v
6JTAtBoX4mUXBJHoewbIZx+c0PhO6MSxcOna+EkIWrIHh61oUGEJ9XJvrzzhNVNIKgB/IaHFUPrq
H9JUCvx4ZeU2eNwhOj3aRt6oNmBhIA++fScSRu/7aQc7awzt7Y2hrXkQnKePWEMZND9hbJVjPw8/
jff8AJ18xC30vO1jBpkug3V/jhqS93nocEwhlt74bJSvpoPBUBgqNloySU6uZRJYgiNo3DF9N/Uo
vGBjIP9uvWjDwbq9I64z3IZXMj4OvaVJumPu6HzZZRWY80OJ7t2xfitwWtja+UZ3+RHCVh3i/UNu
ycSUJiGsQ3SuPaFs7+uKua7B+RHjO/AIBfvfrf8Sp4fe7V8x6AjCZEO5Ju7jxCY+6hfr+6pYCBV6
SAVqbCQ28tVyI95TUJIclku6JCI/PLLuliEcM08LP63YvTOFk+KbOrcP62k8OZWpANhh+KBSg3LC
LtxtfvskrvTC6fCIuiO5eHcfc9EoMHEhau+anUV9McOQVPou4qHp6+lUZhKbNmecHDsk/pgC4vhh
tF+vy3GhQ3q8uSQ0LxY9zQ7hJQ3dR9BiMgKt7+LZg+BH3I5MXAwvkXaAtUgTbXVQttKvwd2VQEEB
tGjnWwL1/ktJhJkyDfbm3rV42DY+/wPKfvIrfE2aeLh5UnK9nf7Ezq+qioDFYzQAka7FOZt6Kshc
H8ngu2SwvXLkne9VWrmnjpTtpwu1A3XOc5GvRgziLtzPLiIIxkx3nLMMGD2xKWZS9almBDE0r9Wq
sL5hSPECa9Bj6Q4c75Dq0PIwMcL3vyRdoQxf6LPOuqMsLeRzQ6B37lZ1LGQOhNkZacKIKh2rcCpW
w6MHcJlF0tMypgu7akbnqiJeOCWNYcS23Fw+8alBY6qOoDitBYNvBoNeP6WByxmptSJum6RTmXkI
PUQWJ8yYW3ZGceO1YHHenzmAudoZggSw77hLnAImy69UqfLHKE2d2H15b1Nf2jZ8QVu40Os1B3tL
eH1Bx6gUkS5KomM+MuxL6FyVk2JcI0AyFLzKiIfcRGi/6lMddvSukoJdUcPRo9+MoWd4O9cBlQhK
qth+fNsjFACxZYTeJto00KvycKeE5jj4WqMnLPFkWT2ymOOSuLUaO0+vLl+wz2c9qhlZRg+z2Prq
p5O7U6AvKhMLHj4upFCqwAOjGdQYnQaqTs2POyMt7eH8IKUNqv0jwVin9wnSh38CLgMoA1057NId
sUVIiCwsx/PIN/LiujYAee5D06kT8Sy7tCMAVdUQrN0A9tAMIxTIH5XiW9jN4TKEtwdQbT1wlDWA
mJPzbturBFLk04dG93+kIK5mlbrdP1UMo1ibRPocy44S4CNyKZG6VsHg9nuLoKc0GZD4UfVSwGNU
b/lnORBQ/d0LsSKz2ghQfxIAT74Mm0XJ/yrfsENwHydJsfI4Q6cmH0NU5T8OBuujYaAkngL/bvME
jTebi3jwg5SYQS3EB4ndvu8X2qEFKZmWZrFdFxNV10mUHfWyfsrdM3skobqNTZdtp2CLFloLANWE
57EoUEOaeQh4smEc7J/+9r4KpSwMPP4+jOhKFhuu6d/CCoAprfXRzAXpgt9cp1WVED6vtX51w2u+
4K/qNLFZ79D1GygUx9Xa4T1ijjCnBl8q391koYsOywZVXxocLUaqmj6ELYWnT8IFJzvGS50B2H1T
OYFCbCiNh9hxuNYJVthuSyEGN3aEcC0Qa4qKosktHmrLVKgJtMWJUm37d3sHFxnRLhsny5hlYQM1
5nT5BZk3/R1+BlaUCLp3FE5jNsObwlCCsSUhY/UmAaJGQ/pYEFlSYCcbTOjvYIRMlbiGqyU/jw1W
DK+GkJBUyNiRlX9hL+mpQMJJxR7XkActmb8VXHIkRlwQMNrdwlqVKS+/GomVOXYtfM0eidOkU+rm
bz6QvxWn/RYLCJweF4YBWmG0xY/YMy0/JfJj88wk2K19gOYSw9OECR4EoivEza194+oiTK/K91AH
sSgHL24rPYLLVKgUFLzngpRRZ0vXra2uDeAzxW8EfWvZUGIKi9JvocBwG7PIVDyAErOI+APTdSRQ
6mnt29dVDTQILfAxcCY3QjP5k2o9Lv9kQ6kEKY16uBIFsqTFBh+VXQSOqh+fLY/hZGg5f74ZdbZj
OGMng9bKf4V7qk4iZHJx2NRUuook5MIIP9JmOTpnCc19MllbcoZ/6bX0qeJmug+Wchwv54uM/YmK
7JIetzzJCNZyxHZc6u6xy2w4xQN4C+p+62VHnA3PG90xfW4EY3a1Hzyzit/iDSVhwyMleNyPFkWw
oCFc7xGCeLXust3xxqt2hyRTnH9CiJ/HM+gfvHO6wLxfZI2K0YPMbiTdzJA55FxgnbkD8rSiCNhI
9TxXgTJnGmCBHLEYUfYoC6TuqIv5CorpIBOq+Iy/I008Mn1dZ5EPp2wmNVU/Lcar7bmvRLaQzFQ4
4LuDVB/Y0LjnqtlMdkrRB8Vzvsrgl7i+jobO9/+sO4D48L8V/42Ie9Mhxr4XxShpTG9i+Ppp14Jf
bk3UiAHWJiOhyDbuV8hhAKNm6G542VOymJ5DiVgTvFJtoCGe8koNl29dvFAmZjQow3G9/UtAVPbN
JtT0fpFkOIWUaTj03gi/TT4KjodYoT3raMYztC5TtGdosEC9eDMQEpMblPgFOAq3HaECwdp+TXaw
PRUhWTVXdsoo7TFig4ZXkOzNDL4nWEiVg+fQoAvm9ZPjQiAQK3lv6hObzKtamX8EHgVbwu17S3MJ
Jkjd2JWcavD5G0DcOEsPPJte6ugomrA93N8knuq4mtEWnvSmJEZaj+Jw3YXJH+jwPReTj5hwRjMJ
7+/W0BeCUGb7bvkOLhwPH7iPEEfVBzxoR9jqTO+ffAlAWPZEUVZcFsRoydEVqfBWynStzbpHC3Qw
zxmKYHnzJgzEi0YEuTSU7Rysoi/iaia6/A/ntjr14ZsEWC+8TV9jeu8IcPB8gLUBbeKoyBjUMZSj
opP2nyvXT0rdgxp3lPECxRro6DuG9LF+FF+h2cPZo+KIa7U0EEw0CkIk0FnTsGGpyQb+8DJVPz1f
chs4vn4lU4xPKqETNnzrBBtHhMxvX2KbaZ0Sq3jMpRr9ElGi20s7YxwRnA1VgPMcwv3BAZg4vZgg
x5WAMJn0e9pxMmp5BAgzqqtJ56/9FLXssKpYCsCuFuqePn9C6fKpauUmgDJ1lSq1OHASfSHsDlEU
4Kes6ROn45e26GTWH8CmpoiPbZN2ge0Cp0gOorDnLOY/6jDvvbonK6NwNP9vPeIgIg5Qxo+0nUFO
n1Ttu/5ko7bNQQfBqeb0P5VoChZiIaeoXfggFHq1Usz1rs1QrwKDoRhEkh8Pnn824Zlu/wzgAKG2
F0IFilUGyLa580wb905JfhMfosYjmAM5fsKaim1ztMyFV45OMRijrXGN5w0DcGKB9hJ8f2gp+oX3
3pY4TE2kROJSpiV3FnD4eyQ2OZf3+/goXd+yeprpUS6dLKow+xjARxKPF3hzzEdvKo9mCKyOzyiB
zIfnQSlHRyvdL5iz6hY4EgWWJLdvbZOqL/wOJy4RgFN5sBTTf24LCjFpWZOmnxfBG8552GbVym8c
Tdk9Ye81cGe3DWHGNRtQ15iZBCspxxyut6QI5k44g9jC4y6Vb8XsV9nVaHZ3o7iDNle7Rj+d9rKy
1TM40V4v/ZPE3ASkDEoe/yx3HyTQzaSwccEMMo0jZNk2290aTS4QBrVCJ9KgI1rqrMlzeVhdl6r3
esiSQuvfqXrSjBlIjdOhIhXj1IeSQwHNmi9z0lc9XUao+onVCGHtIDJFrUIVIfqoI27yfqh3BeBZ
luvdZui0EpXrqBpNf3CobCG0aiJ1ocBokmRyJoMV8Io3tD1UwztUa2qsJofUNlUzwItL0yk740uA
Pz9EYMU+QPaOBHLwmyMRPvN3h42RUe7MaxV1NpFWRLNiI5t6g3jQadPSTKwlZo5CAFU7KhhhF4ys
S+nKCTVk/TZ58LKNCfCn7HoDAKPoXvY1ds9H51tWN85HttHnShVlIy0n0yH2+GAhKJPkWrg8Kyw5
fMMgl2/gANDLKFBpFfrEVKcpLIaH61OlnUW+k0Yp+HD0ogdeRfv5BOcUlkYzcl7UQXKQigDcyc+Z
6FIU8SPWU/tfg4q2U5tzuJ38ZP9KMJ6zCCDNJvEYWBVCP5vhVEiaEEj1SPJ1QweFH9Jpd7vlPJnh
pCbUWnwLT5nYAS24pSy18WKfSu8qNHzKyX3kfEYAsHsgUzDHhj+0cCsBQGHh0ot+ld/pPXKHI88e
g5s65EdZOYLcExvjeaJXbk2RsdLg/OvucNoxTE/hlwH2GU0GmOGunr5JlBaZAPBK98wkwXb2nC2n
2s7yWyqV11WgA/W1Dlt5AHRCTSbCv9inz3ZMzt8qeTqhgu+U2hVVcEi07+bUis+9qT5IxOP1CmjG
e4ypSyMJ4puIIVKdbNyPrLnPt4RENA3AEKEMLALs8UzM1XW0PE7vUDAw7EomjMTMiMBAqh5o3QWY
4TCUF/z3bFfZJ9m6CtEMUTcENa7PaN8/NvPFrJ/IIfc2Y1cf6ltiOr7riOEJZsgHOxNRbhl3BjQT
9Bx5mN5y3T1YA42dX6cw4oGdlqBGO2sI6ZRP4Gsvm+Pu7KkDDtBFCKTsUxjnpmgyHvlE/PamVCHl
HbowVNJpeFJ4thZty20An8ju3yzJQyr4B6TRCMzIrN0lkDUdgheTkoxEvk9JANvXGayrVSJIseNE
SQR9brC/72lqevRVvEVsHhWBzqdvyLcmwzvdBQbPxXgFs1TNcjM0TlCT/L5/KkBmUGaqX+EgA0NF
dKpvIcNGq3dC4DmVt4GJAdfDnA6gudeKDp0/XE9gX46ZMXGStk3xVyQJHZ1vh54tL8DNDzDGtc/F
p+giVXeQBRqlX2TTl5Vg/f90hr1UUdDAI3mlDN5KVBh689jyzwvAvMnM7rReROnWpwUMNPUuVOUv
mXU6/PO4RijgQwed6IkEW8yIQh7KGPbZc6DzLODxqHRCAPn+cfGpkrRJIbgE0VAj0M/RM/TQ0+I5
TCClLj8N7ZYWDkRe8MYNRV80Sz4YXArvbfPF4XgfFlNNxsougLrR6RrCU2joAMetp4vcCy7vAxUW
mBCMUE1Ue61Ssj9Ukus4xV81GRftngyJFUWQY2iQofxG7dZztjz48BMNqhRiaOnJJCJhhWVRJ96/
FUZSUzHrSeeK8xtSyhRJSirGh3MeOOszjoQCmdAKHeEKRv88kKkhDiaWUU3wiz/rB8QRbokYah8W
RnrvfJOeoOOQhf78eJgXwHUQzkRGxOZJOBhNXOc63TjNgE3Nb0OSL09EUZumqsm0st9ksHoKs7eX
kIfzamvJ/kEVLuyc8KcjRTvrl/Mke9ylklwTr3sMIUI7ETj5KUeJc6u7yYHi+ZverZYpvsdl9SbO
vUCvJIl8umI/U+iXrkUQAIdL59OGIKpHGXxjmHOHnXigFSV1EosCyVGrfRI7RGUK3HsLH2oynagK
Pd2xTs2BHmmmtzyOhzdXasDrtdbRniau5d12ZYOpRflJmIVQj5A4p2IFpw8kj0lxIDEGFNNknxPQ
F3iLl1Vnyf7jPdekj6i41n5uWj1xWWvUGR96s9Fm+Dy+QsnB6sFIhN6jJf38qid31cYiT0Yubq+n
+YRnSvXRlbVy8ktF5BokYsrY4BfHg/qT36M586mUXyXivk5mOmgRcRAB7s4G6yKFuutVNEoJIyRF
BV4IuBzabJMzirGA3m2s6Mjs9FbT8UM22o0vo3jCI5IvFVv/5OoyCTVW5Es311jqYonbsOYb7Ogr
Ejxt9GEH19n+SjMIHaJzgCKvimo1j4Gl85KHVnzzVeiurTPudr3BCVYcObSm8FzMNkNFJGyEX9NW
GdgVUrojO12nAuCGgUPlfKMhBSDi39W/FffvwLDF63mVpZRaLAzg70MKKNvpO2cLoTKb7EillHIT
L+OkZmHOpR1t4kL5RQCtU2zcyi0MxSRdSk5/MFq408WqaUqAauLYy/Vw/HeOo4wTLb0czFzpH2Tb
k4mmp5LWOosKoXvJGu2pE86ytTdt0V2ngEHv1g97bTdaGtKcw2j/UIyLRidnhNgUEZlR1BSE25D3
p+LtWaZpcr57kQ2naX/oMeTrZxAguw68b18H54gsMQ+IMIVBwOxv9M5qefZdzWhmD3RjI510RPZH
6mXhlq9YNQ/XUWLrKHUY5nwrqY7188TxN43rDn7vnetCXP79NzKgI+Ef/DPCMPVvN1tH7udIMPrd
lcKY3I9lIF1kHPj/l8U3Z5cbdzGUm4g6di32XYBUfH3ir3GxuNFJ+HhbIKm+Cshzc1+AQO13WM8K
GtVyoI/3TynBOQDmke5c4Cw6gS4HogNVJVNif8TN3u75kbbzfN4s1fPdt4ZMZf7Zz2yw5X4HfN+Z
RVEJHmVm7B5nOi0cSTjFWLrubnGBUGtL1Gqc5gtIwguVAwrrX6nhpJryyBb91tnffQnQkFcx0kLy
bF5ZlusZELI54aqNBcF8dRLrk5mHGWC6FdPVt9goTp+7PHLHG0GnAlVt77I9lf0tbR8gnGOo0Tno
uF6LNa/7LtfPQiR6MAG2EEbByqYyP/C8/PL4rdIYg69pkH1ecXEOYx7nyOZzQhrzceBnpeeE7NuK
fUi63jFzIZTp0Mh9nio4WWulWsIFnNN5z7mH4T4XX8HmxqHdVnkchtBbuXK+Kr3ZA6v0d/rFOptW
he+O42u4NYUPwlIJbixQ1rSh3twRyKkavO6UaDL9ug1cvm62Nd2+toUfTfBsK3bx8VieqbjU9BqX
fRxpl1gtyZN6U+KXTqItKeShBM6KFJ1lkiDaQefix62WffumM3kl3xvpjLZIf8jWN8C2NpNLpEEr
NGFSXr021FlNjS7fEIGbi+JHV69iQxjtkirJkHxIUIniikosMyPeIH2wNjFKfc4pdWUYjWgmDIDV
gGOFRaMbTncVrODIBmD8JnsAhjUgHaaBM/gPcpgkazWyQo3kwMKchKdRiCfPqTe06F3mABNFz8iR
459786BbVJvzhWWS77JeHkoVz2p94XgVCWjhhKI8HQTYkuidlUJCNytBJ/4P+GMegh87eqZgtjkZ
/39eluFAQaXrm4CoPnPAta92lMHKF/IUgdQjTDi3dSa2IhO2paFlY98rriknLc5f2CVfbUP4twvT
BH6ZVbIXB6xhyChwWrvvrFIHL4R1cIQjjPVWwiTfAAdAfLRfKqOp5ZEvSjVlVXBuQaD/9JhXPRMM
CWemhwR9wEgCAwIx4MJhBC0Vyyh5ALZhqwHPI0LSB4xlY+6vzx9aT+nxxnLA0AOgAxed/Abm6vMZ
bp8P4lDXQcygLuHKONzWH3NLR3TZ+V7cRu3G5NieH5SSnpZCrTs/Wa3RDESRAmScfFS6/7N6tU14
9I0BzfcYv5L6AtrvR8eFuE+I8K48XRYPPOerSbiKJowydr6CYS75/Y2Ybmysogwqn+fwJGkWZSLM
E1lNvyiS1FpOoh7MkDVW3DELwUd2g0XUASvGFhRYQq/g3fYKodyx8XnNsuaUiDTFV4wsevE0EXuC
t+JjSI2IeuwG4RdoaC2tcpfipuBalEAl0JTpntInkIAXjvm7uWwl38UBaFepX9V5eSv3A9EMChs2
QWaJbkHU6owgYt1U1P0BTSHuXphbxPIzNQTyc+//TKgZG72uqtlnIOgns1pR0W3T6OCcrp1gZ0xf
LYa/lnwTN/VRKLLXDf6rrdSVmvnrJaMPVPEqqDwSU0+Wa1p/+fVqEz4iS97mX57ezPNzUoRSa+9o
xbw3TXVHx27zcL6a1MUdMGeXngwj03M3cM/QRKpnVvtExY0xxkBzBfDws3YbOKFfQ3EYEx76N4/6
Sr5mxmYN7OMicjLfsQ+imVU1qp9LdjGwbu05pkZr2r4xjpHThz6rkOASneTFUc2fn9HYbKlXvVJZ
u0tjJObBRbl8po1gb6NdcZ3Oru45oHro8O8YX3CgxQ/KgpZ+JABoC3iKizWJLpQkNVK8GdSoD//P
03HyzhYqyGcidZJtMfCBISFjjsqbovOkAiQ+qfAoov/h3F6LKtL7m6qfZgrYLyCtLWoONlSA6n9J
aUIAVonqtSE+EIR6MTP3DH0ReLni5WeDG39svanleM3wm4ESQx2G2jVyY47CTFctguKWiJBK0R3t
Q9o5tRsJUATHduotNnAXculYCAX0dOyCErFC6edWONDXxBCchmsUYsvsGWjXzoFVHwfvX86O/RFQ
NAFca3bP28TnNncQG2yEK9isQHJHn3k93oTOV3lrWHWZdReCEKkvpCsnAzQG9W9AkVTqunnpXXQz
bypk+Ubb8447e7HjfSxLhIRZ1uAUF/xIIyqWjvWlmXNbW8D9YpdSvxvfPnChpV9YX1lrWJnTOz4x
bSdqueoES/kGuNzgzhm7BX5Hwe3nEoV9kyoc+kn41i0ooAq6uE1ZCOdxq+UQgmy4QYgddntY7ZIn
+cm7PI6e3pFjN9jJ/+n3VCILjYUN/HQXcVD8hmBjoVbT+/SQs/jIih2yM2Nt9zbFTZg7c6+/nmnE
gEmkN6xJOm0jKezSUzkyplSSKkd82qsYb7h8Lbd/sx/2DJo4e0rcQClfKyZC86BlADiw6qnvEJie
LBdFB6H7eg56vYOa1bkIHbaPB3GwigaUqzehgDjv59YkWdzu2WVlNkBUy0tFuPDFMXAnNS8KqNtY
u7lZD3j3VAZsLkqUfmvCLTDl2M3XaSDYndHhqB8hITXNEH7sL1EGwh3dIcYGt0KmtVVp5eOT8j2G
WTgvsj3WM4yrm9nFKlX0i9TfHByMu/yR1/5P2A1JLzhgVCvJnpPYiHu6pKw5rMAsL+9zBt01HsAL
9QVxFNJ3uQVvkEXKiodFxPfdG8oHOuKivrQjiQq7CDhnLOlOhXmQCnYTB2u0OA/ZHyGUJFx3vnjT
6eo9NopeCNJhkZcaBbqQ9x6NPhy2+PWm5J1TeT3nX44F3tvC+P3ptnjkm5058PP2uGx1VGVYQIaK
cUXGeloJoxjlNX0FXdXoSNpnllKUv4HQm9FknrFETOqeaf/T2nSWz9bVYatfzNip4UgNNBQrYUCZ
NHpYck3wVisgXJ9vlzk3Z5nEcDE+xb3MQnqM7d2l63u/DzMl7EwYzJ0pyGYmyyMoJsqS26kQzm3e
2Y1lgsyeLnEr+IXsRMZ04zg7kF8u6RofJbj4nDxSyLqLuR1HADUuwipgkxM3bFBtGa2jc2uNWyAl
drU0qRa3GujosCyePoGdhdyU5Qlhx4GfbheoQOstS/bHVLH08Pgtgn6L3bYEobAmKGWeQxTY1kE4
F7fQxIaDc0mDl0GGfJ1lcaNAFheSBcEjcTeixXTgJ0briGKI7wli4qWZXJjPHWu+b8FbuyfV7Rnj
191+Qp2/7W8AkWARzE+ekQHdOFTGehsoPEVtUZ9IebzCk++ZroEsshtqAqqH4bGMzeN3iCSOccCi
1MmeGUiiiev1Wl69+QwLUrlsgVHH8rOZRAyYTtA1H5p0n9nhsZFz/u2zeNDGzhuc8MpQe6dKJMEd
05HlOvFs1h5Ah5ZM4FrTCWFGuqknb34ciGA/pIHNALaFAFm/khInqgi6GEmVC/0URroXnNPW2rIA
7MospxEaV3EZyq+2637E58lfWExPn/aIkLpp1AUiOQ04mSJGOsSjGCS34o4i9pe++cfZcdydQwuX
fx4PvGQhgL6HL+BPJjTWVIxGiS35wmGBDkXg5MQq0YFYOPCPqPOgIA5cLe+nGX09Ujerl1VMomcl
yP+vhkJv+dALMQ+7T9P0fp8Qc0o4IBHDpHK9T15/f/EoLA1/z07fXLOuXmwYlRMu3bA3f+RrSpX8
Q9zGHOEBsHYdAvYLNRbsSktoXlE9pbJoEp5DZDEa75u6XbOO3YYiUcqrLR4T7mZ6y1BVNKwpG2sh
v6lVk6kScoYjAWllo6SwzKxK1Sqg7sSh5yki+VcX13f+54SKlWkar0z+yV2ASEuw+f7VB2Nr5kVK
9ZU4w8pe5Zb+4Xw4GZpwQpSQ4jv4AmP1i92xn0rfDVuMiPKMSa5taFEAwqreuNiyB2L1/NvQpaiL
9lOOvSTSnbYldnI9gk8LgHnPgEZAPEbP9m4qI/Rq+wWDBawaou1mwEqvFcDjaLedgoww6ukOj0wu
O/stIMX1poKoCy2r4S+MGWj6Ftgz+itDerIxRImjTfJi4bY9DacJSCAn+YG9SWbX8tduly6T2b+d
p2orSN6/RXS/sL9RT3ZPhiCBaFHmHqa3sKQWrcCFwSXTV3jVTPzhRCi/B11A58WlFRp+H5zDBj0T
LIKw4IBtwpzIlMDPhF3JHWCsISNIk+i4wp8k5AoFpVgtwSwGi3OqKsv9jIHRv6bJCUY0CI/RDCjd
SrVFD9t3EK3TtDH4O3JpjUp15J+YKbMifyn6E0fNcJSpq8rF2kUhCpF8ipUP1wnXw1NOPggKfRTb
3EdnC6jrBaxRn1PyMg09wz3fXWx9LLXKdinWjw6BZ7FLVz5fkdhG3/kpO5fHBa2Ozyeqv0qOyO9i
Ne6TLa7XM8K2SOG7dOueN4hwUmxz6ntP9gWqOeYChoHG2QMMlB68/Vo5yT7tTsnPdTb6bDoaObYz
o4+EyDIdcbKvLMZZk+i9IvZrU+Q4MUcqO3oIwZrzdncA13IwSU5lBdmfNaIuZtBjYhtB0bdRAZl/
q0+keQiK5MN7nNy/hHBXRXd/OjZ35VnOG8s6vLBlAkOGGSDKUIRQr9OBkPp8xrBJmd3PsQVMii65
Mga8lyL81g/kmVCaKEpl0zGU9D9NWzZiV0JFI5s69FbQUnO4CSmxiUFslcXJn30/nxH9T4HgoT20
Fj0Tg4F7dDy59nRr4qBSI096qEzIJt8ytp3bKUOf8hhc9HbfV5cHR2IUXeFWB1nMAR2Ud+6PX8c5
BNPEGTAvQejtf7jZSlwM+yvyiuo/fOTIPa9oTjqAvjv13EIo5OfNLOuR7Z9AzQNuNqGHZfc8fG2N
fZsBxc03/VcrXYxsx7sOcvYY24sktDN0MnraW0ExkClMPSDr0UNZHlFKsOXshj2vu67nbJXxYXwR
GgmT0EghRd/9v6MW4LVAB/OA7PBNRgWjEQkTJaneNDgxkEnm7VQJQaYPic2bO40M7fSoOGklAjAJ
bIXMxZfgAsdmi8WTFrSd8jHyKyWxNiPJIefrJfUSom1Y63dQmChSKKTO4EFBUdykrUl/eIimM2H3
ki/E3qa5EZEvS6bdQA9Vu8yGMInHkX6zWApQaKOKSFKkr4e8rDSlnUPtENIgrubsTccNoFMQ9sRD
TZDSUlZ+0F1vSyAvtVJ/aW88ZEpvxeZYdy8lV7dePvOsO29DN6/NIUKyYlyQPiCNDrvt7hOACBZi
g9j0KFF+FJz1j+zQ5ST/S+RGuGr7XQl61pderzTjWRLGAoqgl/xgX6tjN5KU/2XdBVZxher10C60
LyFYc32kObfHM1SbGI29d7tIH3DXK0zWFywAQCCVgRZ4cJKbb38egV2bo7dyQ7UZJgCboKTZyJw9
HR2S8lqkbodVQsKvXU3mJlhLEcA+PC+etHsTFLOo5ivq5Dyq8xZgOXXGr2qUJHV2qgDL952z7kHW
SBDYE/P12VGcEGcj3/Ymf4Jhu7FksBIkl9H1DJK8odc3TZMT0F4lNMFNjiP7xj0FvuvU55fouYQm
nKOUmbwE1eeU63hauDpZozq91Z+7ZXeTtD0VsPqOdlcLIolQekehZ4Wn1tboLVfVNCveqNKT2UaG
a8bmqBmtF5QYnesa0Y9shKGV5gXGBSIkyFrpbjZlFYvEfTDBAhqnSWNgb8q0X6uPGgkc9lDCAnFE
5HNMhIdDJa2706+h1npBVLGYqJCCGZ9gyNRgkZGvT2pKKdZ38JllHqSx0enaCPr3pQLbRatTx8aI
hdiDtpCvJYT08ryFjwHdeKUcoTYuWAtEGdqiA9oh7LvNfQW08cLFduJpS4d4Z38FxoSdCWQzTjzh
LaTlrAMgK3QkdpFxpAZU/y9MRhGVoDtr9PtZtONZFDT/6ygRuw38FdoNfnwhwfmhjX0904iONzMG
ilcEXEDsT0WlUhaoJA9VqTX9XVDfdsm0kr6bwt1bwEjNSFPdPkE9FYXBr6xcHsF/y8Vr/DGfCGUY
YgQC9trqpm2ly4AecktTCslG4IlC5MRbL8IcOvIwr70YYE8jjpUw56Go8P95tlqc//iGW29zA/yu
6bbPQ5W3++BslYfPHtodTt5Ok12FAE+m0JCXj3J7KaquBQccjHx5JH7OI9NvEwB7qWpXkOi2uIpx
nokhIKbKgkuHc5mHSVjNmLZgV/KRNqQoFTepTude2f/onGV0qoKIa5oXah5/293O/Kni8DyOLl+s
fU8QeapuLszVXfB8j4R1BONjVvA+zCvug+utUmqN2KbbZ1MFZwke1p02X4choDmoHp/dVFJsF4eG
zr+nd4ZuKgME+wmtXsterHYKVPIq/VYPHbd7LXuE7tV36hjSo45yplkRuwuWjrzmLtuxLYjlkNzz
Ccg0xOVxWO6Ju6JqwXmJ1Z554NwVqWoI30j6vTGofSmqnS0I0152WLLnm7SNwc0QJqlc9D7V5ufG
Xz8ysrfmixZCBJZqure0NmV8mQfzco2LM7Cb2YD5kBf2A+3ULXuhpKZXQYiKUsYK6cNRniDiejsi
q4eM7tRmSSMM2bGODDQZxAsUv3ejZQwfJEkdRHteCQfocGUvk/6FFscempPSSEfoI4OUIfXaqVC1
DRI8c8iLSpUZgWw5nwTeTU1VlOcJ25137TiU1VilfXjWTfA4vGdHi9npdDmqhqK/50PWbRl2mEGt
4v68bXliTZW/oD0aAzVvdURqmHb4pGXdqn06/ANuKvyNlYZN5O2b8IFjdIJTKN1GiQhinmY1uKpc
f2JpHAFY5RYtx1NLD2JlEpkizTf8uig0KzWFXV5ZfIMYF/HgbSlmvfokD7PkiTy5QedMlwcInY5b
xWik/zWRXXYWxXyiSkxt0x72fp5MEV10zS92tcM5xSyp7crv4+WccLZKTMa1eI+IJejMGUHeidOo
x0DuDyusYP+dmGc7ItedVUUNRf4WoLYyQZmvOT5EMRX4R/8DtjB6M3iHhf1TGCmDrBZCVmsWkzrp
0MJo9KA6XbJF6VCnCl49QIGCzdsTbX3Dkoep09uC478gX/jA5Vuf4saopn5N21MxZ7mHhdH7SyEi
gFrCxtXY2aazzMw16QYe9or4DhYWbeCOeofh8Az+FBFwA88o9vAamVppsv1BmADBapGkmETpdOPS
Qf9j05yo90/5mLSba1q9NEOBrsfM/7Xsb3Ver6H7pK+aXVj2CSl/OnGcFbxYN7l82n7Z/4xLp95N
t22yPX/4ogkzCrrgb2wJo1pkwkJ7I0xyW4bGb7QxKCjJ/rT+58tGw47yrfKRWqiYzoenXBKV2yxw
x5TQeRWzStv1Mi1dcyeVAzoBZVQrB7zt/ZLELeRp/KlWiWGq2+uxWdsbXAENV+WZu/Oo9q5xTbaP
P7tbrbM1IK6N1/6K6T4JO/tiXMCmDXypoMymoEY8u9qmdn5CVE00Lkou/ghmPC8a2uSiYYBAzMBg
eUJnyW6roOAbfnUeta1aF0NdON0N56Tm9KpiCG/t9Qty9HH08zqXZjP5nFrlm3WFdfCBkJnBZo4w
1TdQUSblUoKIxboHs12OYRjfe2Fc5p7mz1Ag3Fa3/uYcIZYdSHGzTWpom/QgAV/zHe9QjEapBwba
EBw4tmJ6J3hh+7t+0kiL5StCScN4HnyCIiSwSNnL3JZmJonI866a0hRt12oZGnk5ejTCPPHcdRcv
x5em6nj0MhXXI5CS2SEs5ur0POKdJ9/xJwztYRRufUzIncj9Es90g7IYNfp4mCMghL9/XL/VKXuW
XM5KmmXtlPIgQcRGHgzvoofWWx/yhYTvVzowBRh/dhA5v+iNGobn1ZqPwy+Oxtfy0Egj+cqRxvGY
jIXm887bvBosQ2unDdSxuppx+2PrNVjYfw4u5YEJxVsT1Nr7YYvTR5vHScYMslCJPahDv18Xfkyd
imOfz4yHiVnYQc1YV4VT9rvk9tk51yUK6hnqPTYeRe+ra+qabZADR5RNC/iDWuoB3t25979PHzBH
V9abp7Y5181JPb+j5tMlK1zp/WhOp+PvpgfNwPQLeYMz3IVD3y+8luHsO4Lia4iaTVihCIPsPJZS
WwpMd2aX/4QBXAIpys+blMnGKO17FajzOsr7SBWwkxieVEmo4MMZTJFxvp2f0Tj1pzmMs4DDFbiA
qN5caErVepZxJ1RlyuPAIplJYqcD0GwMxpwP820tBB88g7rb6X/MIgdPknhg294GXCUwIDzcptBk
SgA9m9oUgESJbfwPWtJ15xqYCAg50i3Cxx0ZTsonYeUgkKqvRAYIhDUktOVYnXjvySL4W1ZRC2b+
xDym4YI24ia89x6YiY0G55Od1EDPrp2/Hyp/ak1+qnOBYjVWPuYE7kC5j82HB9mcaLtv62eQOkyP
zps3pwQERLUfHI9I55CQArr10Y5wO4yhQPwD60i6BEVTvjEpKAHF+9MJ0Wb9YUWkCasCSX0VoFZG
/F6HVUGjmmIQTC1o0qR3z5TKdkILcZInK3lSJRdxGkA0mdnGZ8DCczbE4jJ8A578kjfDIwjrYNFa
ogycq1huGaunmCg3KgqPrUB9sz8gomHW1MRKnHen07zEl4EX2kSr06SY7jZs+2eJNug7QTPIfcwi
8vuk5wMo8Qi6JiW+hJ8xxyrJLEWsX7gJU0qR4Y+/nUTb1nZ9snAWuF9Yv0HswMAkXxPK4GmVLB1U
9i8bzBywXfxzh1Ene2vjQea6IfZ42hTcQ5Yg+MJqwRSAu1tkp1M6wG8jTCWON4XxES5DQkT5uIi+
rai369lX4NGyK5AsC1kgUMDyqwywAWdebXCla+PqZVBuspnldccvM77Nu0CYR7QmLSGDae7pkbnV
00s316s8gNC6ZxBRhnyX1eveFRZZ9qwn6wLkaCR8+S6ODMZkr8my5KyQh1HO3AM9bGNPvtCeDdk1
aSExtTcKsNwRY0OOlAM9xpPywSMtS0WW/B2tJGvM4i/f3pwp+752khXWbrbZYE1GbgDcpU9KWWkl
OguX/GWVFOLhhdjW3kvolGXsXxQRluDxyXKJm53tSHY2zVGr34gnbvK4Zx4XUbR51FHlQ60XGr2D
4tK1Wjr3tzsqAo8nByKB/gL3G3uV/ukApl5HnYyqi2Kk1SyH63LLDVQ6G/nLW2xrh9mFJYhDZwL+
RD3X/d55locslue2JfumDZHDLk7pnUdOahgH93s/K8IPkNx1Il15wqWx7RLpylPD9PvqevQFy6ml
K8W/B6ca6+BvexY3ry44d2/CLshw2y4Yy6ru/MlzTdHeZF7dYWJIdJ5a8JaWVE64SkVfrnkat/fx
vtmvDjO6mdmvO1O0DWht2MMWRw2mQrNQ48nfBlAg0I8gV39ZAstohPabgPnOfWitz5mCUdsY65g1
Zex1dGZ8L+0LE6eIWxNkodJFWeIm+sjrVGGshBkutfEeBAcYdtueheMNXT704HZtq8qwTIrocOEo
pC0AAc4VKh/dZcb8SyykM2Q1HTyRZZrWpnaelKTud13MwaDLXl09FKG66cxaKu5SXiXfYb2IxGU9
gubgeBtSDHo+TPcmt/z8uB7p2sWGoKMNwCAF+M7DG0lDgCFl39syYYLCz5W8DkHv9MJ2icx576Uk
ZdGyJI0phTmg+cQ783dgdMkUYNmYIabDMSJhgVYWQtOXn6ZvzFGlYyVpwbXt9/paQ7PqAIdWNykZ
gHHUVmyP3IiBDAFStZuXqsO8ZfvQXELM31FQG3p8nR/3e7f6INrXJwKD69k/YSn0mrCOOrovln1k
eYq2vRLJrzOspwZ5ynNPqaD7UYr90hjzu1Qkj7hg90dOlBCyne+S/VYRB1XQoAmmZwrw8clV5Nv/
3b9KY0vP28qEiFoZ09VSghj8oYK1v2biqkb1yZyoCZ8PpfHFWzUjbmak7FgvAK3H1U1PoUtrvSod
npKr+4TkyuWj55eB+5VLD0667zgsYnB/gZnKhe0rQ7ZdroSI+KVHOAINeO9EAl4Teh2UoiSZFPNM
GvbsHFK6btJWalsRgTOkKm/9XAfkYK4SHaxElh3lWsg4/Ak77owKWrSRm5EflSBIsA2zu3LWltgE
w+PX3OnKR3i+CVEG+nj9qpI1z2cN8nfWTRgFcGHcqx2CzioCSDHHFsLe1x4MQpoSiDmKNEEKmso/
glMrRYntL1Q/Iubo4thTpJz8w/UPSTI9WTycu+uM49osmmaXlb0LlTcwfRUBwq7k9mOjpd90DNnd
8gu+Gxy5fC+hToiITaaFgBfgOjWBCOsE5ZHDbumSY0OOsJ+1E2Lb/JSEG34Z+WP1ks1SZmuJ6GIZ
CpXin6FhKAWbbLrA+3IHPGGsB3ozwrNxwpJ3Nb5C4rkLmryJzsJrsNbtWdWVD35lbX9v4NEwZHLS
HjWYtDe4sMel8xcM4oSzpSBbe5Hao/umgogzSu43LCJyE85Ajnf74tfEDzS6z9nfdecu2/gvcZr9
SPZaZyIYqJUSPj6GGfkU1d3CqAONAlBRAuJXdhs5MECCSAPcFq44K8qMGCdb7jHDjKo193h70yxm
1k+P/C3UwqUT/pBJEM8BeBgWwwr08PGtV7t7qEy8PYeKqw+bsLTABnRBD0Ykx8YmE5s5ROOoVeMD
6zEEniS7eix5SjAjifTx7k8Ygob/iLyE+SjVDGtFOpM7Ks7YFO4aHg/7nJxS5Qty5sJU6UaPgaJb
WYZxizc6KSrZxUjeJSxvvoW7O3FRVXwqtcyoh8nl58gDoRDdLBMwl6cpKeNXXn3Srb/fDfXKQEcR
bvFrv07kOC37uOQBnO31VE7PkYDoTv3IknvMg9ClTjrrXyKMbufB9aS8AEqO/IT+2lwiw4ceVKo0
u0sz+hkUxiHvtzzYVS1rgRQsBEv2ZSuCPXdMGnHWTvdjI6gC5OW+s4ncieSCCJr+yEXaC1Az/iml
cgi5woTe+f99MYBUHFWIHFrJM8DzYsvhhRkXqLe88TD9mEvGUEVkii9CFsbeRaNaCvwvV/S/5ezu
UG/iFrJoqcD9tr/yqXbtA51tEiTcqB5Q92bm/ZQRxkE/2J5rqhqzQq+3Yt/npSzGFUfdhZLmRlv1
kRywX9PUkugJwdpoQu8a8Bue26jhD33GWLtYaOtGxW0dwbhEptrZe62BEJ+syNamPJgFnU8vf5c3
MRBnjPDacaCKAf38aBMnZEKnjKZ6nr8pCfmz9BfijC4MaHwZoBMAZkd/Wj1KDyJXbt2lMx67J80M
zw0euMeoPJ4Tqg0GsXPd3lHDrMfRtRWQoRzRv1/qnfU2EdyTgjgV8mMkhR/Uw+FXT3JOXm27NY5B
F4y6ukzH9EMjyHF09OQvmsR/vjchDsB4/m2G6ZLM/mG5OXSXwyVUo/fDQNRcWURm4Db56PVQxChS
fBd1/M88x3GYRyg5w8DmxOGNLXOPHANErPUuH8emidpNUQ6K0qZfQKZnek+pexJ9B99/7Yf1w2sR
locpNxIam3YixW9NBVAcR0xhhQFRaR5I1uaeRnzlnuUVJTDbqZoCsEkZC8cSGCWopVqYwkZrRqMA
/+9INWW5j2GekZAyO4V23p8dW98qCqPkO7nCgIiaVPyQrhhm3X5y+cIC4wMUq8zk1OFvUF74Rale
YgInc0WElbl3DP9Az/JLbFAJjl4nev+Vf91mgvr/ZXCSp/mxmZdRwGQ4GUspV4EFz9bqVbkkaXaD
CaM6/N6HqWSZl3NI/kVYSi7jBebz/LYv45w5P7123X1z5RTdaLPmJU1++KuuDYhcoLTxDRWHDsar
dlzQtym30IoV3XQTxLMCEmxpLMY+ewOsDYbUdUNLJG7Ctubdpcs9mkmYLbePfhrsUImeeWsnBSSP
JExvL6O17gotEVWozLBAa3mtmTdQXHOnu0Q1fjbP5f1/SXjyDmgyQNdHEWARwCH2ITxvWK+r6Px3
WV/dn4000yaum/3qDK+jsnKU93OP9w9LW8KO99keuq5FriDAV3LdR48cDKK6uwE3XDNTyYe+v3NM
FkgGTYHVIBxh9TLMJZqzgdySJnQDVT24ha6QERk8MqsubWE6Xts54B2YdH46q4ABTydox3qyY5lh
0I0wrOZj6c9FK/Nb1JwFlbQnEpxQ//RkJC47so7XBsol4Znm3M1SlqDR297cCm0g7dISD34KFLvp
nxb3BAU8ibqMCFULJmSPbZpHrKiJ6WeDdMR2ljYVkpG7wl3AzJDNG2Pn8IsQ/USOr1P/fJ6ixnhT
A4UpDo9hxzr9GmwNk7IZf2D64kHfpmhJQ7ur2oWMvfom49igFNXst6uf9M3MWeId2Y68jLm04ngc
HAEBbt7A3NGX9ShC2PUCjm3llQdS7o67Aeyr6kchJftIsHOidOi2zSkw8/1NVfl0jhOSmuqp277h
KmQPxSpsif0AuAi/NZXL7rhR+JwxB5qc3nKt1XTbdKDh7wQclaSoxCcsE8bis3EeAwiuMT4PxXjA
mPEJnGwBghciTsFyTN6W99xPkn02BXw9CkgcGbdO3llsLhOlX8qaiysP/ULemFhrJhiRLvRJC5+w
iO51EXZ+soIjO+xjNDfmfB9b9E+MuGZ3wDvwSDTt5pvfGIwYKlkTTTO93+0M0nGbo4iU+VQLYcoW
MrLpDr03siCn3orT/OdtdRrGwDk10l8th1KhpKFSlYE0wPEvJqBk5atkVj7R1r9Nh8RwJdJfYKWl
jMUYX+BnFt0JTI0zQqMDx39s/zIyMAOe7LwEe1aK9E1tLOnfvaLFqWVyAfQhQCWWVmHa5YGuYvbj
5JlhJOTeOk1JFikehKiRYGXwZ1RVJLj/VzKZRuQOXgccqck6dk98fYweSVYi0WtQKmGTOzZPwkjx
AniXmh2OgegMgAxuYzaPr4FerUsp8+o+numwghWO4RZJiO04qL6Et1TkzMBOiIRGlRT8TVd0dEjK
wUWL4DJVGBAc8tzapFDXobFm5GDvDViLYjeRJHFlvD22T7a+BqRcbz8+wG42AEs8HSwinv1SVxPl
FIS6ZpiF5WACO2g6MhKb3zSln3D/NgKvIxwVpokegCUXijkLuaywwUWEVAlY3z+u8k8XLePKLFA4
7KKsdfceMF6cIgb3Bl7owCRvlji7GAHKWI1mHUBTUmsl1w99GQ+9LxeLy03N8x3WWUZEzQgYFPIZ
z5yUVfFIsvf2avX216rgUtCcyFEc+rp0Kq+hCoj9MiVmZOflnCy1jzWgg9U85j0zO/Ed3OTBk2Gi
93xaj4GUAjnA24ZeTRxlY8j9NVEhqSqV0M9uQMcGgm9fKyiKFmTxfpJY3tMPowq8L34TXb7zrlUO
bD9No7LK7rGqe9hkZRRXYbh+Qfwn598Ugbq4h7EMpQy+mNmiAPvgFX/LFuzhl4RCYRhelIyGFZfF
3U0uvOPXLBZMLFTEE0UhImNf/59pLvuzu0pMOGd7vQhG3LDyrzf8V9ri9UNRMAgO/rslLm1u5uJG
LtvxAB09AhvSxy9/+UqRa5of2e6xvqVkRKTiRkkp7PASpEIBdgZbwfZDLzptq1d07WJcX3kyTdBI
vjlK5eUFbTqcPGCFiD7agAcx/hGMoOol6h8ZvmxFgiaFvb/MguFHJMoIn78MEVlqOpRduAcY34zR
fp/MgeLwboh6xlJSxIUsUqiVBDCZT17yZEi0rQlNrrinT9hXcrHm/4yrh7KPeO67IqrkoKC8ms+k
6VSzmItU6X9Hgtnfxtfjy3d+Vj4CKMgHyZqBVwg1D7RmjdAC8G0pfBtNUzNy0w1nN6W3+wFOkgHY
EexFnGXKO7OoSq3frXfNzjYmOQ+X71FOyqW+V7xXbT2RZz05W4BpOsDw2fLMim8d2IkaJf78JK3Z
CfgKouO281JojbyyScMtVrTCUSDNXIVbDE2mndumZcFta9f1RwwukDQyTq2UfuFJnEASir9A+R9w
d6xH46NwAubjrJyhlNFjeCSuXGPeiqX4oXtZmHI+1yF49cMLLFtjlwFlCGzOqwouZ5XnIYMdVyG/
ksIshSkUwJ1EwxeHMCJ9lusuHXxmf0vJ16yGYQsVUKJ2awqNHM1tcTRhf+mpandUfO70/2RAKxK7
Y16zr89wwgVlfrI2WF8eGC3NoukiKWTavdUk5zzAv1ikaVQKjNEQSVayQkA9eLX/kPLqFqTgTtkP
o6QEabKC0A4q40d8JRLKzGgoUaPV/iNozaIV2uiYnlCfHo7OL/8v1uqtHUN6oG53lhGnoLP82pVX
ZIwEl9DGYeMnHbaSaBsOdyW+HcKsj4KZW17REOBuv+8C/VS/tESiN9EWWDQYrwr/p7GotnaUMXOK
XGL2i4WO62fCesz4JoKlqPzqq7D2iuxvIrS3W1YA+9bNPZ/UwxLEz4aHQ/WTNlN43grtS7llRQUz
htjaw0QVGs57PbMc0J4BAORKZnYSIcGUjBguuhaDrdV9HLrqXRNqUczd8Eyrque/NYPxdue0KhJE
HnmPJFR6PtmdvUC6QJrQPWv9aIL1R/AX1m6krIjDxflLwrvDiZ93aQgkiWopO0KQnQH72ZULzW2e
iuXpIIfViiXPlgMTIy9vkiFS36EmlVrWdaLLrj8U7rLhRhAvpGcgl3lGgKwVcQ891igvwQSwMnNu
S5rLkcXtYv7rbSOlAMl+V5ibxWTiQWs8+oj5RbhSXRVvWvMKsjOrxWSRi+bTe0H9Lx9XptjLGSIX
KEeVB6Urv1DmVi/exh30CIvS77LlffvTBTEV4PJ9NC3yBy+PYJP4aZISRRYPrlLg5eLYFkh9RCf6
o90GMzbAEZzB8Wt9xsRfOaPdnTJYRPVinYOoWdcx8xhmkQKX6aOwai3AxeMijimG3IUFWNRDXBtE
wVwm3IKKdzTysraiIbkL8QHHIhSxPvaKNQPWFMti9JHaAdwek6+YIIjoEkVc54tONHOy0bL5uyD4
h2/dJVqfw+n+L8r1mWnZLZjV62/hwxzN4t6xZH+5Zi72t/vqYTFSSwXEGKPKKGLsCdHtjzXXU/Xz
T2NpssNilkaB4sjbIWd3eXO3SEdUCtbW6AWOXWxAb5XV6XY69gcXvXVPIa/WtrFWu4dlSRZumLXN
d8/ETPkajxcHBw1XMjtQB0vh5ysRwM7zidSpzHRjqbT4zHM5X9UVq/29YXe0XAgzkl5zLXf4tZDZ
vPEPmmwoRkVI7S8MRzN7llSOqy0i8UwxnlPA0pejaYfQFJSsBBaLAEUqI7S0qKS99LG+bJ5/iKK/
aoWfMO4l4Ew37VDa3wZ+mQCS7x1FKkiiGwdWgBj9PIFMwk5MMn+Tt4BYXDurcAYAxV20540Po6XN
LghYMEaz/bYOO5NYVYM9nxx6h2W8nh53IqQQcLOpmerkJ4tuze7iqthESoeasgNfSJHUAiB4KYks
N3t4ijJQKpiI+4m7k1sRKfXjIpNgZKLq3suBjH9rsDUXGWOsZhM3EeRaNwyy7cahPa41XoKacnU+
xlFvsSejEjHxF8C4dQ+WAo2modiuslx/XUwvBaEoXUZponB5zVQYmPWdTFRTobMTAEZB/JeoL0qX
D97StcIrNX/QtJhfX0QEqjEPrkwXNQ6GLaDBzZeztCGJgiNetrR8Kog97D5S4lyT7NpHSgRcH2et
guoCNZZ9/9L4FRB/gObeOldDPtfp2/wW67FbwptqyEsRAfQ22md/z63jTnIs5wrsDO2rQ3g/Giqz
OI31ENoUH9vaJeZA+WlhnajD0Pfb2GRJrrPWezZgToUKNQzYCix/oW2VoDXnGgkV4NwRp+fBCWUr
W9etTLDc4o6FD4ZAHxyLLt2Il74FZz5JJH/4NEg4iei7Rqsx2SeGrgT8pSlPa1XTiTuJzWUJULBw
Tnd/P+YRpli5lTYKrGamftFCOcp5XfqadwpIdoUX6xpl/+I/vaUu3yhYz+4naJEnMsWdhPfUfLNc
BXlVvAF/d0gmi+zawST1DAVzA3OrHYoF66gGF35JBvZf9T9TCBxbgd1ZjyRyFryORfUz6/pst/Th
Bf4USHXvCUAf0JyJ0D5UBwMWdHfI5z25HfNclN4KCldV0XMKSEWA95eK7+7rKVX5aNio1xXZTe6N
3/ifE6/Dew1OIdcJb4PCltzH3ZGRj/If42gfjhTGZ82rgVDQeHD3meDCRRHL4TE/yCHqUV1TOX4Q
eKaVvajRrzxcPCqulBRB658c3v1CMrKO2Z9/0x3y84eboY0BV1w2WwsZcFijufhB9nANV7hXhKZr
G/9PpITtf7AoSBRNuziKzQVo3IiWVcJyzSJMRCXaB4ZtHu3zFYSFkUzNSsJ+04g2sLIei/4rtAWK
3CKUQGHoiZd5QH/MEvp5C26gJnXjA0ePrhv1CDWqMZYkniiDJW/wZP3IAo26wdpnwj4QTuJVVEH3
Bs4yH2zvTuZkQ/L3g42uZdW+zijvEUjnMtSGJm28qQKunu4CkhBRz2SZuJWa5fl5YBT4xn5C2WTx
ATxXSocWMf38B3r2KbT1A2L2VEL2PLq/4UlH6DcJ8kVGxgEefcCGxqc0zu6ih4rNgKe9KzmP1KLs
PBB6ntajmd/YUX7kraA/j4sqAxEfkkxYENkztgZ+J683oGQ3MFlj4e6cMFKWn6LTGes04XBmoNF8
uqnV51VUO5YqNvqx/ZjRQW21dir6blJZNNN1y6sPM7/yzqbwYzKaMOilyqHY1XhGW42KTu+/OqfQ
LlyL2Mb9QI4X3HPBUJif2PpO/nXokl9zwQ1lPxEsycssdAKVkbUX8S4YfIkDAlzwS5YVS5QcQPGL
bNvJp9dJwRlnSHVuVjnW9/2meyBMvPooFYVkE6XLkSpOXJVD2WVVmvNcZL+AbBZLbW4juw2PRxZu
BArs9MPwX6v8qCPygoexebSrK0SV7qOjSqBai99p9r55BhDj1scSO+2MzLW+dQb8UK/ZrnbOvp97
jeap/fOUuRoe26cXfvXQNzMnPpw/+47Pxy8GHmZtMsFnrBb6/NYjgyR5x96xTvkMzO2NiNCH1AEg
MOzy42h5QBnnhSvIyl9FsIVj0IU49+5BUQPBICnG98B5AAfGztPjm8g8yxB6ZuyIkHwOPkp8YCIu
7siqZAv3W0cyku4LuapuKgbqEfH2+VfDsRCnfD5Rciw1IQR/eYFN/1ps5I6qPeNCubwf3rn/RRl6
5Oje3KT1HUx/X1DM929ChFdg8DaSND97dlITZwseBGw1RbzkRb3YN0SacFGxqc4DPX0luWI8A2ck
KDF4nqf6GavY8aMk0Be3+DgakEuPdBwjJECrDqrSyLnKaBRrhwca+fNdDXcgJ7LRXXlyazRBQUfo
jnkkgibkL/91w2uepTdFSPzHdZ1Ia4aqVm3gsmmUW2hNS1Ql2nQDncNcGONaoGsEK2ETxiHJBbXc
dq8S7hPmcSUqEweJY/1BnNA0tdXl6fX521/6M/Zmt0m/9TSHLIQtiSRJ3cQezCUw1UE40G+ouwlK
AhvHjhfdpk6kX6uZxfX/9h0hXuNEhYncHmR6uWQxv4K4ERwdiZK+yACdRPDu3PRKGg/nWFNHwwpP
YS07KQ2B3q/RbQiG6gFI8GVwoykG3mmRFUhX1CNbvwnPBLYMdQTrsRkwynuiEZMiHlRqvXNuGP2B
BDSNG9WZLL2ElfJlbWXbNwKFa0E06yMlo9qE1zqopvB8RLnU9bkDW3z/F39zc6DXqaWjWfGlPEGj
xBKaJhV+qXUgyOJOHyarhU0mIvZ0xQG2o9OFXC8M5CAIfnwIrhylTyTt45ltx8PRn4u7+mjeNJDc
QeKjrGt2v2cxTW128F4bvQjB/jbYYSUq/2ZmXkXbrXdFnv6yuptl2fFDJOb6672oWbrc9bXFcKy1
0uUApK0hqxvEM/ZU8rs19oib4GulQTSee7rV19ORZEuW3H+dE4RkXUmOYU8zvNE9P3XIxRPOBULv
Uu3CiYetdiCzDc37yTVc/jvzGu6p65CVCK52BVAO2GiT8/D1536nZIB4pIGBQzD1JXd+sTRYLZeQ
KQY32pt+7wB8KqPHbAGndOfinrRlwzJ4n7AvgPpc/Z8OLDEQEiRyx2DO4fwkIUaRZ+V/UDNnBpYf
nFOEzKvfmmZ2vHzF3Y6+mDEDfq5RJeUpq3XNEpdBDYh36LO0dLi0VoIRYRQKst5VIcsJUFDLpnTS
EydBVHbLzwkTXFKPbnpE6SiuyTVHit+UzcRwLo9VsqovHrfhSrQSbgMO464Y6zcis6DvsaTqGGzP
yMYGorFDPCurpUpJzwQ/jKI7fBaS34ZHk04oXlMXuzRYQetr6ertswp7G3JxP8KRFG/xU1ewROXm
Fx1zjBC1NaN7IMjAyxNG1ZF+3h9sBJvqyZNL2NjZegNoHbaiyTM62LhP9PGCTmhha2ZkeA6JyRuV
3W9xIjltXfjRgOmjDuDWBnQETVGFGHJwZy1VvcUK19ZMix2Sqk8tMSS9s3XNWLvrvSLOrV1uIB/o
b0wgnLBPMraTxZVHPbTAAQnrja8je+0LSQsFD8LlRhGpEduI0t2gMLCT5MzDfyHVdL9Qb0YxYS0p
PRBaY1LGy4ga5Ok84PlamS1jYe8Ilg2jI5wOpHo8k5//Q+z6tST1ujd+AftvQxVM4MMIAQuxOYjG
IEGBnkDew55xpp/yKH2r7lxCG/neYkyEiwsmlMmuVLiau1Y2nMMOoxqFBQ2gqRJ6tX+3EWvSw2GD
92rdtlos0dDLoDXUPEb1Xz8mtNrpTh/e5B1A4cVvFKic1/sf4dCvRYYFA1X86go0NNwYq3/q9sfD
2Tw4Y4Il68fbaK49pBRkkGQm/oPpMj+fUTCGPF5uBroOKcl6f/lNM3Odyu3fE8Wsv2oEkOddE/48
XFY0Ii70c5XMLaZsQkFaPtCnbnH+6eHwwEXLW9avuX22vL+4rf+afiGvO7B2NnA4qdlIKh3Micy5
BzpHu/+K1K4Jonz5ezkDTj4KIEZ1iHN4fCWIMP6HmuxSx6lx4PMd4Ju8STYkvfIls1wluqDuC8Wh
kv5k0UK0xYEEQbUB8oKoiqGjlB92nSzmuEReIIYP2bPro3N29atKGA1VMSTR0dogqqTdlQ2gSs+e
JnbXkVbe72wz0aDKWtbO5CrtQvvN+9ztJm7qxLeHw8pw7hp3KuWiF/16BUvuTA9sW+kJJZazJoyY
SvhwnyXOGlrdrZlVw3/tk8Ne+VbxgBxoDHzLQhF+t3w3/kmRuTxhzki7O4fWK+g+NaqOPG+GXLll
CgVM5DkUxc1FSzj9e4EBK4Fujifiat6X5XzpJrRBTCU0ncwyaGh0KToMSMRevvPuvqma1cMduAU+
KafbPDeqhAXwU8+R1N3UOq14pyhqZkpccF2KiKX9B7pxoKg6V58Iu1baeUuR5NVgIaySjn7e06Ba
SIz6+9FREFF7eOVXO9vhzhki2Ii+Qf1AeFgj01eRbnunpiTGOE+iA5+eotWXCXESYZrQeq+JYGgO
dvOQJg1MhY8Z57E305LbvxUnQlrPQjx131izn+4gRfIJV23sSefQjCbdRF6OpdF1WPU7SWxjH5l1
PkRSmdPtS9z493ZuM2r6rGSu9WRyc5CXh3lVneJ/+O55xamDYIcYMSJuV04ebpnh2LP8t3o1MdW5
3U9PdgEVgfmhQX1J2bpMXGRE+EnUp2LjXmDirJXzmZATmvt8pTpViS2+QIhPO/6AJFL3olUs1WEf
Qa6FWRGbB+v+PxsbXvwgJTYzhY3WAPPlBKcmI7YHeAES2T4OoGnLJKnv0jQTG1/3nQrh5akNYreZ
1uCae1dopGhEkIjWNa+m+SBMQzU5RrvEEfep1rMp6COqUe/p45Ni0+Eb7G3HMaXkOqgU8LGMPdpy
iQPkBy30dRR98EccRoGJ4hYUiU71rJbREoFgGJ4mVzMn8oRT2Z2EI/PciNpzP5gDF/Y6ctQwcUSZ
m1gk81ZKkU85Ag14NROe7/32b/GyDezJudBgc7fAi3C+f0hkOBweuUAJ3DFfw80UWIDEgDKSz9f4
gK1NhQxtRpbidvN/enyQR4HcfCYbz859AOqhZOCP8OtraXTMW2VCIQwYDZLIVg0dR05587KS3gkG
JUYqPkHg6nbAZEGtE9uLn8EaJQuJfTgOmL4MbnjquqzCfuRLCkaC5Wvfby+zzFYVB/O60Ju2PCyq
4982CpiQrY1BDZiRzF3ljcefkIUIcnQe2Mbznusdut390/+X/VyxQKrff259r0ke4bzNqqFdYycd
Ct2S9d8oPsyCLFkS4N8Z5ukx1qbodfvZ7lIo7EKEx9qLrDEiXODD8A6UdrIF5WSCHu8TzSun/ZWY
wUE6SzNVX29aEd19dXO1+jEzVwQKo0ivcD6aAxTjdnLSJWmmxZxKUFHT1+TG7HC2QFrJtFaxwzko
KYFYw41RfmEieHsMpTc0FhwcKEJKSuNTLG8G0uParbLFZTCaxPvcjXoOnCkupOKYMtGUZn490Tfu
ZoY2ljY1og7tfnBMpxMq3i+HVw4KcruLXiP4s75oF2O36XidOhvsa0ilnJzfK75b5/8CDEl1mZdY
KI4kfOPrEpoYG1nMFbI7jME9lLKu8a2GbHZIo+VQGALek/dOP1ZdcraqX3FOTMxTz3pX12p8lpeA
LyunpnQCshPP2QU25Mr1rdtAE9g4OGYaL5yFey9kcjU3BSFIWeFLz6oq3nrOENGzl8HHT8kaGQ+B
UdMZ1GYl77witp1HW56WqHMO+krAuc0TiK0ymdCNRZupKFOGVtKmggowhq6wl7wVgA2N5/IR+twP
2JaYqkTd+HHwJ8+5iCmmmj1KBdH5cMmad59pAA5tSn6yQcj+8NWtorS1otVVrx5np4tIYpLo6F+z
0l7UGraEyiiZMuwW6xvmEUzHPlvLnGRxk10cggR8vw5v4j99XA6ZH36Y7wPrcErWMBAehLzP54UK
0a+Fjz9HshzhMeQ6Z0ulHyk5RRqVn902nlCnp5YO/d4VcDO8NH42p+g24C+/uxEpG01AKnM8O75T
M5eIG+yiyiolKEHsx2d+6rUMcHVeGWwKzUDZ0oMBX5I8MZ+ncDf9uLFhivZ4yozdOqZ9ZWUDh41A
bs6aNRgOcvbr8K8CLlLuy0vms2j+cE2R7dY5JUNXl7WhukXqRAlA3wanWTEZI6tRqOVI8+BVfW1E
4+LlClpjjLaZHsygS7icCSEnsfsC9TUtBkYEQGCMaACu9zWHdkCN9Liv3m1PoBIYgjS/Oe9o4ppd
JkbEU8ynVT0qFc5UwP8XthYYdwhz7HvSjHgkG55zZf7vDglsW1sk53muX9L58zfVILJDs1sUA3B0
qMPZvoRfRbDV2ko7reqV0Sh79YbvdQRBMqM5XyUWBcHTytQKofaCGBPVihddTzizHDQc3bjZSMuu
jvOgOuOAN6si6SKoHBud6NQCuUPyB06ASbSCUfUR2gD9sreiO6mxsh04/ji7Qzeb9Nq+GuF21lBG
d0EK3Ed54p7kAQF0LR7rEqcOc+6yvWUeUaygCL/zhq2TIjwof9e9SOPW0t2Utu3yD4k6oBA7xAKm
mv0PvN10e3/tMIkQ8gEHa+CVjrxFfXxEyZ9enH4TP24qtcRczohuqy2s4MQaYypGwWYbB1YduyMy
5kcsdCX8w8DzPOf9yeh0+6TEr2/rXxNH5U7M0MryPneRnI54MVo/NFh6oicwWIUZkz9tPM+ACfwA
jUQbmob4YJuUltg2QoyLvyhjBeNgacp7+0uHIH26OuHJwrTHneCNPPvmjgJjZPkbTLeOcBmhDRNE
3MrG6/AqGh7wUNu1m7alnmBACn5vbcFj6yrZtB2CFfmkUbZCRUFBiv9dV/SYdvRu3krMRx4JWhIr
LF3Gtacx8JItkgA8hZ/omREsO9X+8W+BgEZQsm6IcCnLaW2ifd9Y2nlepPRiCg/ZntEB08gtWcBl
7Bpz9TYMrr9XvUPL2oixUh2ghqDaKVMkIL3VBDRbeKeY5GHWqkYQmo6LH98yLgk3QJ+jACg1j/h5
ZFbYn4ShH+b+1KDa9JkLlotNLc8ns2Ry5x62fYA58VvBP6YQLH5TYZUGvwXpQ+e1Vw/pQSQQ/qbC
9Y1Ksc3WuycTEE5GUFQ9TzsD/D9oUQQAgfH5zq8gIFWWUM3aH5JmUS6jjg3PFh1EHjdQMiFs2vuF
P9YwahWRW08qGrY/qh2YGU64kJR2d5LpBONVL5lMO1S23k7bPlHxP8W5aZ6aPEdw2asnTnPy9Mov
VojU69dbyZkAQc9eBxE0dx3/t94Re+baeIDY5xemzS5XaQ6CuYio988MHf1GzdZcZpapMRW3Ybc1
anTqVkkE1NTye0oHjYd3wGxDkXyRgAgjTp4pRq4BgZZ58F7Y9UdFquKUaRwKVIBQqLXjaffZ/Owl
6/3ZoLduMKr8zj6IMXwfCBeUAE+absT9YhPDyjqLn84g4ylA5c4yIobh58GgLDGJodROMiaZopYx
KgtkObC6rODu2+8E0ktdMVUeqU2pBsomRrGvxJ4qJGJaIDVMRNJOZjugc19+6SRYnP8YN52LKfPS
b1aRYmBh8cIgW1ViQGRLk4ryzPN64z9gqFBvOilSFqJaOmj/2EqSK1uFVFWoop6i7LRf7k3jcrUM
Z2uzkZBrpEwujHHYQLWG6VNQgZ4CByn17HkZI+RW82YQnfWIz5tQnCXVgK/4y3RM09Ni/a168+2I
qLS7C/O0yoXcCW811K97Uel1qArSg+RUeYHrS4RMWY/OvMOBgMxwNIp7PZqw/9mF39hYTp8QTUGj
sMMGihLWkhfy9W3RYEjNsHTU3bXh0n+Mh/R6zFnXFo5o51J121goFdPEtV7UQrTVyX/PKoTmZnbB
tOzqJ5CujnRcswjjrtaeyUtw1KSS29a/8SIflJgaj+55zdyucbi+fzNXyJnnlOa3Q3J/NCwEXUF+
dNjlL1wG2UvNqnmHqY8pLmqx/RsDD2TZmDoyAZdfl9iKEY6GuT6GpjJY/+KQN3BlSyLBCCk/3x3M
e6Coj0aCUav8wXXJntLc+1RljysbyI0/yUlwJGdtTkOBjb6sYmmYaUR/mP0pUhq0OHzwXmsNiVI4
iYxXdKcYAa2T0UFlf+7zhLyj60EaF+QjWH6ljQJrZ38/LQROAkmTVIDWWlyyP8XA5OEOPbn+bF8I
aAcBdPHkD9ojz8YGY1WSbJqJaxhrdVhM1G25gVCs0SdyXYmNrZh5jtfdcFWc3M8Y/1smm+7koeAv
BKBS+ub6EaKrQ1/KwFHKMDBwPHL/yxgMVDNIkiDkIs53qvl9zbdy3G5kiFkuKk4zQvHCXG/9MaAz
uqZ0KgNk/pybxB56D9bv5EEk+IqR8KApHBd+a8rbmuqurpq6d1NGP3/YchZSTobCT+LbhvnFpq8A
BwLyEB40MGmLFw4CO8JP7DKP8k5vTM9C6zx2JF3RO4IG8l11nOXAuO5gr1VhvkeEyNBnHNfObeAY
f9zcQ17JgByCe1bxFXVkG79VbkPpsEkd51Tgn4oiN9OThSGEQHcpv+RXML/Mm2xhWhrbrTKqoPYT
nh411O3m4z7xirAVsWfS7CLYIH+LiSv7uC5EbzoXdwZtqlJoBjz8cu8A1LK4F5DFzPIb4e9Ag5CG
5SIHq68RTTq4orQC6z3esfe7YrIi6hag/FmO/epK7GvJwjQC/U0zEkOXEphafuNtLXvBEQ8Wk9I0
OoKz6vk0LBLdKeiZ2lBlnNNgajVuo9fdmqLWqsBI9Lw/JRfE8eAS8jGnxHq8XAAbUaRxVObn/UAT
LsR8XX7B9fjMl+YPtsBnpImmNBcylKVXG6XwsDC/eN2fbWb4bCLmCB/5GAFx91ZuHAJX27WABxYR
GSXIvGR2I6lf2CKIPf+KdykHe3cf2zBRVf2QbOws3tNlcsLBI9oABIj/+eoOCW7hlKtryu+O+dLw
9zTChbpJ0/4ZA+82XDbjTlhQEfveU5bkWY9LSiDGDIsLmPJgPuv1dvg5VcZMUP8eeBI5JE8rt/J1
pnai9ZrtDaETXRuCj/lQdJgimnQviMwyetflidXfGBQgrTDY/wztsp3fdc3U15GaomLPFboMSCks
NtPMcituUjZ6YrcISkrUc1LDOEGnKPGC7H+DcJpgjmAhzJSqISBZOEwjLxkiERJEZOLyvV2z28an
cWQR4mERK5aU9+78xI1GR3mA2rPpEH9ItoK9it4IFRuR/Um+nSGxKRG/6ewvOuR0a6Yx2GY3fOwS
VQJQWE2Q4lNNqqMx8G6XaCu2nhaMVwz0g/i/AD7wWdp/Ux/qysvzEP2JTtSZTOeMqUC/eNTDlYhg
8n7ExKgOctiTO8B6ycCUjNUNAH/YPYSXrKgWazxYokBXyiTd+8GTX7qRCrT6ZmVWj33N3kTB/8ES
cvjTgBFqzRZxq16zOEzuWCH/hLs2j7pqNlRbN9VRfNiagKwaeabqK3Mllp+QAPvj0IMEUfv7qZV7
/MQuC9+VFGbKWGmW4Q+9M04iyngTyjlfkwdj3rr7XaiQRIPqH92MjJqWFMTgtB2j08sAgb6nG/DU
v1scV3nRCfBtxIXt15TDGk4b5ws/8zkwGIocjHPOfWb5IYUWqmOPK0uW42Evof2XK2wbuXAC0OxS
fr+6wPVKcK0yUmiFm6AdRfa/5C9lb4FwUJ0uPInkiN7EyS8/S6mkkWe8dXp4UUfc2eomh4FsKhKp
Di57QNiaMTjTB9vob66keeJfhW1R8YypeGreTAYzkfBPFL0GZ+52a0uiddfDG0z5YrgGUTluAA6o
AV8OcX2ggpcYaPrvp7nRfcfDGIWVjlQVHB1Izvdn+G67HIM5C3XK4RogjOjKa0ittAjVZQL9NgvD
ARRizHNGzR4Xex00es8FVLOdfS5KEmxfbQr9OH+p7Vq7bF2Es878dz08xvlS7aG/x1fbkwGzwRIu
YW1azx/IyY+VHmL49xkd44AHHNHsUaX2+pEIa4HLW5qjjFDc0M8Ng4xGv6VEe/eK4utgBZsdqy+K
UydAVomaGVYqrEZrPcyLqE30RK2a5G228z78n2FGcB5AXfcHZJKzhoC9EmOlQxik+WfVkT0BBr8T
ADAScAoNJ6CJ5MHp28fcFmQkNhmYrWyF0E7UArO5XWVlAXzy5XuIGy6eSdxhn97Vf+gpxXJH17py
FWpAv4tVMF+NQHzX1C5Gs6uB3v0qBZPGNXrAfKYOrUFHNxsz73gF6d42hdWzIDbHO/M3shkRb9aU
YLyKbcShhAK/iMn/zvkF/N8fKaPqb3dYL0meamyUz3QfI7jVyLjifpCfwPuSsILmgO7Kvq/Dj+wd
+yh4QBg/5441fRVItr7ZVGNv08iDQZbyXVpaH1nZZeX8B/+Da5ObvGSDOTdS64SHdHwwd6t0i3Wv
/2H6cSwaMJEh9i5GMtXtLDKfwfnuElQo0zPadLGUQFmBAFNNIzriZzAhUXOzusfx9hox+AVDrr6D
2QxrdUQvKrXc4cyde3SlODWwqz/N8vM2nFv87fynPny7ciSHGmwQv1Ywvcxs5og7PPjVW3cZcFoy
Ji3spoPiV2kAlxQfEWCGDXTOiRuvVxjp7O6agl+FcjJedy6GfisAzYPZ3ot3csthjF1Qy4Tocbzg
Syt54lIT0iGlCSzqxVyUX7wxeqGgu4dAP8Zfi42xQLO3dnncJnODKMWkW0EYuEp88O9E39LgUVCw
iAF+R+01idUv+tkTG6DpIttP4FIZkZo3aSwTaKXJz5gMyYEZKYoC9sxuRb1pZVDG1bgMFH1yrJcH
k9BxkU7DF4y8y4SEJBJ8GGpjT6UPoETOJN/07IU95vqX28+eVN6vLifbezEJj+zu02XSh1Aw++gj
EsbRzQSWK5J4oTDbo2U7EFIY4EggPItVYBvIxJlazc+MpKhKeN0Rt7cXmQAD+B/HAeglANeVnKLP
XoE4Z3ANXsdckVUKpJinXEbQeD/NGvdq1urOJkMCHJs3cgFL5DD/3RtSuLyauPwix04dFHPVUE5i
zRtTYzRMqSPB6rgwKKkPz7HWlid0w2RNKYeDOBj5gho1wBxwy8KjZ36Ak92lFBUmayWJXbQUGqIM
oMy35U7Ng72Vn9woQ7Vc1BGuW64C4/zQaHMjynvibM79pXxISAcaRueZaKGpkqa+QF/Ryna5acMa
bEaaoXKeuuYiazo/MPsamQBG5WaSLO8a+E75GACS6tmaKJFX4YUzezWxWE8k1h+Dgo15AWpgdaz9
nZwMIh3n3cTeG8MkUXZk7ZiZgnDM4gylt/V4mGk033XUEmXXB8MKapRObMZc5dDNYfNPM5cygyGw
VAEJpj0S3pDvIBir6NodZ9T1dKkqHMhsK34r1UQgazFEcdhBN0EHbcDTz8zp9ONXlJE5XBFxZnOr
oRfLzBhBcUb+um/MVWN3auZAvTSfplRm7MoUQyUwUn7u+TZ7Ia2X52E8VvsqOoiaxfhu9JScw9ij
lheqTlYBH0FwuiSL0MgN+cM5IoCZj850seBy8Kf6UEF6w0xsnXLWWmYYXbnX1fEZvP1zOlkED4No
QqdSa8BJQqtQm0mSnKDyXwrMsyYKfkz6KBhguL5elRvATqI+q1BrDLSm1i5ICKfUGr3ZC6UCsrLB
jhBN+ZCeevZAd+wTnGcyg2TRy83NGo1c77UuS6ut2NLVXD1qE5phw1y+BiJu8UdQqCLv+xsaXKwg
86imohctuMKQzBtO2/8P/uIU0FLMYjsSd5HzPmr0yFV0JdsDwdvQ/V0l/3bt0yu+ZtyS6nU4NQIK
SWfzx5ApgNIxcUj8JQJ9m6TdJKUtlalop9AAnFzUc82kuDiemOZ1YOYLQ2Qe8A4f3of89AN6PCmV
N+zvogOuhJmd+RZp5U671XvjuBOH9LVdKIXjQ64pNZEvtuxX/ID7X0dKeutrIvhDhkT5Tv+YUQv1
3W0JGn2MhQN4dmZNlUt/Mynj2QbfqbMP7r/QZl0OLlzvqtFuytwzBmM+vaVInKJyqz8w9p3WiTrA
425v3HSqgwR7/y8TYveYTYkqj5QmBZcOE05rDYRUNysIdeWYWlJ83SvGDFOvGnSF0W4GSqX+Y0Kv
WRE1ZsQ1rKnVIP/y3V2fI1PJ9trZ+toEmwMCuKGVUXVCU2t+ui+4qttG92GSM01j9lZFQklw4RIe
DIEminrs3+YQX06CNdw9yGbIm4iP3hSbHYPX28B/zL0UfZNDr2/VCPC/iGeAzKdxsgvemSZShlxJ
bBlUNyIm9rP9cHvrphHzfYyFreRaAsI2D1bNM2TaLRR/eXQxWL5khi9lcXNkiQ3pXHbiKRcKqkLF
Ih5aoytUpLFrL+TG890u1PkU7EUcU7qABhxO5XYJrUIYcGcQ0Bu004lo+ZWBjUSm/23tvUqoghL9
ZDyxlu3giUYiYlw5sdX9L5ps+inRDEBJwv5pMEU5vA0/3PR1gTe+WtO5ZDXum99heH8On9bxQzXK
p/gPGYhKO/vVT9oHh7Oc0g4k7yixFyqBUtE1rtwkPyUHCmc9A2QX3XInu9Uf3Qt2U74kotqzJOMC
huxguNniRHMncgfVf1vxGCKx7bOoUgEATlEsPNdm95efAXaGBp+qRpjZ3v8rGi6amMePja88P8kR
u07mv6ch1HUR/jRQBJFkTlLvn8JMU/Fw9Co9XibUkzhqQM0yn3uympD/aSQSZYkemE1jw6CC8Uru
K+7I04ioyel094iPSX4IinomIR190XTGOu5/azYSSoZgbvsupsp3SE4iF4/Hj96eoYUtslcu56NM
Li6RihPh1v/4PlVoWAJBSrtTYEfLYv2I48BnBWPAu59K5R25ZhMPtYg/75vqC4QyLMwLS2TAApi+
LeLDqyBuVXYmRwxqR3rir9gO3Zm/y7BSsmB9N9q86RXRqoJddnlYI154xYLMPKflSLho9KZLOUbK
UWj57DTBDx90vDjd5XRAmL8HdayQ4shWgDW8m9T9xWYSr2JzG7TYTMGJo1amU7lmgOSCmCOF+emo
7a+C8dRlkgYnIXv5zPDG4SLPjKehMg05xWsDRH7stUkZvuGuOVPeGH+ZD9R+37sjKj9stNlVUTgt
i1wBWBBumcMAb5LbZslG1FBJhTFlaoATKdRpQ1wD/xfU3sLUl2KCy1Y9NALzfbVECsBQ5yrHflTc
N88tGf+PzF5oWRRAvg7GV7/8/gxniQJCtGnvfgvwzgX+A7iw79f+qnG7k5w06BISeFN2AdR8wyLb
ejuyPbo/zm8NO5cFquAbjQf93fKOd6TKEkdqR0aIwtcQm5crQ8YUZE3hKQe7b8sLra2gWXrbtCTS
7iUdP+VrxNZqXIXNR9JDvsUugwPiUHcgGnQDivLuY9fuwqO97PXRjOtgePufRxaGbUxRiYkwwUiD
0Bbv/neKiJI1YsaZl5GoIwXpr99ZGB9lBKx3bhmM9dvT8nwqkaqaV/okjbO3/1FtMmHdb61LNvgx
wy4vXeyuFVTMQXp7C1Kr6k3TxcKZFBy6zK4dj2dG4gI2fnErCfkno46q3oXjnFLYO+hfKmI0yTPr
/eTqtIa9m8yt3WYfOzAJ6pKuHzrUdD+TLKvUgFcIQCryJGtkF0uPuKEkJwFT3jrDi1jDJsXPAMl4
2tF7D5ZuUu4LbscVacMbfkfHw9DF0T+qjXMoaKVbBur7I9SEpiOgK6ZycOV3ow5nxat7dkA3Tw8c
FAu1YIG0n9O8QWKiFsmSqqbbYSbmyqJXGecC7LL+1AGQR2lKXbMVe93hKtyusyYF84JM3I6mF5CR
HhJkjMirFwBHR/yq3CZfX298Ah/5yMwM1cUIGbsieF3FCFaP/Pncvn9N1FexKw/meA7pH3vdeEqJ
u01OL++LVUl1xRF5AAnC2HCzKySvyFiMQMfPnUFIsGGx+s08ZJ2p7WGtbaOthxXEClu46HXSQmcs
yyLUM6A8IyyK6tuCw/YGSy6Ezz37FydoXGoFH6EKry/odtWzW0G/7cKkG75MZglUYMjiwiyAJ4ZA
YxuVzBCgRZReADUJPE5Qlp2OwYPWOEmS2RcXJmk/NjpTBmVZNSN+KNruYeAKCHuLblhGngQNcHjm
fc8asb2myJKjBWpDJhw9sYVXpI6rlvcCNivLE9NVZqG9nrYv7Vlr6IGS4zy7JcMK3O674EUWEbLb
25ptF/0gTmOpnRHAILicWC4O0178NMeSML9Grr+TKpedvy/O6ZeHdusMm1ZPueBLiTkPjb/sOya5
VQa2ixUAyKnlEf7/CG5aImRorY4Nxtrz2hU9b4JCqAx0JlSwKGFUiZgJ2aIeo/m68dBqjUygbwO0
YUTUYE+Em3CqJmyNZM6mhVT04FVaJWhQZPjCr2ERym7t2XbbM6a9NGbDJlrWrL5/5BaOzAGQkfLt
fS5gEX1F1XK3t0jJK9ULrBeK0yqeObYYL0Rov5HK3FVp+uodI/FurjlIQJcDM8YFY0G61QlPlBSC
HfSzk7sxBudIKitZKoCxcClz+kOoqiUhjfuUpmQZ/Zdht288ZZtFykdQwCekpwNNRIlqriD5QN/t
halvLZp/2hCVqK0mjP/DmOhIjlLU3zg85VdDGd3e5Ar+wXR2UdtfjbBcpIekoHfsTn0pLRT3oUls
frj0aeQ9SsHGMMASQdXN67u34zZ1FmRr3pN9WYnMp6YTXAK5l35vItLuZuxpLuOGCr4BkRQ5EpAD
HOOSvzwnUoyvMVGuFRQA4D5RZJyIp9LSX6oy9CL/kaGTo+m1zOLx+nlm0cK8fO4hJQq5uUEHsNcf
fayn1/pM6+/BCkiFFlFjkw6zjp0g+NMjwa0kNOQAYjkRPGwSqyteMpJQUmnNS7hUn0OA/o+P4C4+
blhVQ4jH8xUxTckZaSsyd0/ltd9JAUXu6ZHkR8j3RcKofFZ+yHxdN0i8eBwNOxIRbofboTe7EDli
6KisSblKHKrQ4rx1SApHKKER1Hp3StItgq3NFl9hmHPyOT1yqT63SfHGeQSbSUKuLqUL9Kz+6yoi
w6dnrR1m6+x2Iab2UBg+jYYdNJ/gSbQmhf9PSEPKrzsMoy62gMsqUtahZe56ZxDFcOz9w0N4+a2x
J7TE3WKcW1O725u7S3nb2uI2p/R6nVeIeM2DsvXSjetDbvLXat71n/95WTxXV+i7AukIMYW6AAay
VKmDfLa1B5xMFJg+lNC11AkGreasiBz198gKZFi//qQafjVlwxujB6ytWpJrwjO1naaBzJ3ecFsH
+iF0gRwpCyG9EtV7MxYeRVOeACZ/qqpO/14Un6WWpDdoft83DcPSOxKDCEcFHrXAHAoocBHGnfJx
A/iR15tAIRntgjJRMMhFSNsZF0OCezw+laKiMitBW9NTvnMpOa5LV39NiBWrvs1R3xFPA5gKgzHP
XVOccsREteku7gqbxTBKwaDzHtBQBkiEgsRWaeAr7yaQxYmjmQyeav3jgSGqBe8IULMkWp3F+oy7
CS52InUpRQIcMCQf4pUYKdCAQ8zqHSprO9M1WS3hKOYG019X1j1v6Iq9dv1HYIGsxHGsYOaeXko/
P4/+IsrL++yoeUC1HWk6OEs64PaPx/A499Ka6OKAN2dacNEkpBdCfLhAPKExoBixCiWiT5CLNsyT
wgL5u0LXytzJG96Sl0Y/aURRtjzkxIthUMGOyfYCxHjm+WZvXUJbAogpz3T8NXCNCMAhB/NyklxR
2TDmSM4uGuj+aUWO5uNbiElg8WxT3KY5G76oFsiYO81AmM1ybcmzdDGvDVjuZw9CwBVNMFsNEOOQ
5b0gF3XZ2xi9HAR5AJRF5jz/ufxn6eiLrW9Unfl2LoX0GAZxVsgb+kOPr3XexxpEYbLehnhMntPz
kjWqnbuk1DuC2IQ5yulBs7TTSe3QXlUh4iRYHVpz56tLhoW7CIDEJDoF3f6xR3n587abx9T1Vqgj
PHv3z47pWxhMcNjNfqsu84dPoF2atCc2up4uGD7E8g0+DGWJPtY+o+F0v5j/kXLSW2Z6OmK+AsBa
u4mkS6dtDkSVVZlYQaEX6rXDHe9eprUBS3eJwHryGEtz/Dwc1QsIMQ0M7tFlX0oP/JxuZbXo2OXw
9Gf/0soeMBzvdUe6iPyBn6DAOoyJkNvm6Z2yxayfWrDMm1jvnQsKV3lSzQC1SWFdikeSMh45gPZs
VNT8PnGwViRQkAhtau7kARm5AAFrlsNzM4Vhg+ScT135e2yAzOloOV71lWo4cBk6zHr/xLQmfBZG
v9JmdyZcDPqQcigyQVyBKLVGuWupv5JBiUGxOKFXRg1I/xgj2t9uH8m815LCq9VLtG0y96RKuMRv
b1xkfssukv9kQTpxKcD2m4uksS0ODZsXqKDuTHPVBYnA0grAX2jPWvM2LRiqQ46S43QBS0pH7ezD
oKsQpEMx9//UnMqXWjpZmLZkBTcsdqCelXeDaxtUmNFIPu5qFT7An5QM/Qo95GAHdg4Tv+FmtGxf
Cy/Nwlqjs+sdI38qoJQ6GeZucDgzJMQgkTqiUekzuW3uUkWKD16XcuL38reL4BVUbm2FfJX6eS+w
2xRYsH28Dlu6liZGwW0G4ZlWO8WUgOaIXdiELPhs9j+BxgSgdAixghO2RTqdly51ce9018WGT9uy
oSNyW7+7i5o1nqSWmhnj4rb8zaGHxAFEGk9Ni9L7NykhWeZpO5f87pKtCGHoXZk/+T8amGcNIiY5
a8LPh/XwdooQD6ScipGD6S5hG3ygnzOyzugawPmmtY1AGPw/BCzZX2iawvKQ5irMA7pxRU5TUh+a
d7B7AoRehkTvNwS9gtgOTU0fDPHL95HR6aXsPf3GEvZXDu115a7XsrUJT4QMMR9kpXzH0qVYNrcD
mdXD5shxPNUZYJyg3KFt3xVUrknytdZ0TsJaQVABrI1w8SK/ml5sQeh9AZD4e+XE8RTRa0lLcWQa
fubX3/RF9y2dWtFUfEUr4KW9jZXvuTRrjXz3+m1PnBBo5GUakXnH4dARmRjMjsEtGfX/CVPherxM
HhmxKg5ghbR3HSqptc0D/ahaipyYSpNjnQoyKg6BUofZO/MQDLi6pn3gEDMX2I3V3rNsDDhlQCn/
4eidRmOgBWVJ5WlcWKoWZRz/QtDJmIbt4+DjuphlpdGjK9yldAYoIBaU/Rb233BQ0DIxqLPtjbak
xzFJX2yQILbyVgIbfPJjbmyHmTCQ1w0zXyufD94J7koyiz9b0kOBoYfU04nJ+I2LTW/ScsLnVRmE
qGTMe7zt3baOLfEXzxMJQT8mrnqEU+Qyqw0dY2lwFD6yfMHiMUc0g2NrrrEPxrHVf8UNlxKUgC2l
VpAJrd9gGpCl2uJ8fAr921Z8RLX1/2064IcQ8nCsbzq3PtnkuAl7fXwY8+wmDAR97ruMaFUVtSBP
iwJZfvmPL3wQtzypkjYQUThP+gsYhcSLuIrXctqTa3rNXez5yA+Yh18g0t9UaXmfPCQwAr3uHeIC
atsx3sngjmuHpcWG9HNSUybUZxdGXHZCWnITGGqxYWndL9zSG3faTATMXM8S4yH1vx5hW9+eAV6y
l+9yUFq0T5ajWBU8ptWSAOEZvFTkdDGz36Kr74q6LjfI2sQjXHviAKMgAOvdt3RJpKsBGZBxzDS+
tyX4E8jr/RMncqEggR8NV62GRJnGhPx463uJv2ppoys3X6dNcVckKzfWsna8fsKeMQ64proqKkuI
iqx+gnTFYVQ3equbJUShGkUVWafLiZoLbmqVmVTz+p6lIfQBg1eQyQdyLMNQl5HLk37BafeH3ja2
lZSyitYiwiIv1q6nODQ838voCnJkcxIhmR0y7CVFXpeFd2Idioil6Oq/7UMuv9Bgpg0tuv+ifxp5
EtMQdQ2i6kIMh3ATEBV7MHHq7j/nlcYhbO04M00fhGunbKL4SJt3dByyvmKiJFTs7zStT5HARijK
BgCy9MHH9R4B7wsMHFr14cINWp2Wgbk7hQxikaQ9SpVf4DC6HJay94w6UlOfoVWallaQcBX1VdGb
WJ0s5Jz5fqLLjBUE2j1rmDkLqjxVIVsbOjA8pec8n4MGK2wyxEFVihDO3vvZoI70yWLM8fipo/S/
JAjvSwInPEvWM3hCyfljpBCTLGJZZh8BCLky8sm0bxC9AH4NX88wOFcQC7b+848WeCQ4BGByyoIC
EF2XT3YmDkROAfICGZNJe615DoL8L+Ax5KmPVGBtZeiQdh8FN0IAm3b+YOXrgzaiKT3cSBGj1HOM
UFlt83SY7exQckawHqnftoULt8yuE53g/tY9u5ZDqjTc1QNMz3VBHrdQQFljI3wGXW/LhJ2/J4jy
AEyoom6H3a4igBY/3FDKzC2Yua16771bOaTiUVnDrwS80OtnwwUqlY9QVsMMEOo2Oq351VPFDcBj
x2p25A66WKFjqZHbNLwA5hNo7VPCi2NfzvVovBINmUk2S7Sxu/zODMzTypm+nIac4kOcc7He3WLK
R1Gkpr3XWULo6zp8mN7tOXQji+h1dl9umP84oc4mWGSrlmPWNf6xy9gj25hLeNasGcs7hGBp2Vih
GfoDJr6L+XwSwsKmTN+x40nYBP83T8sMnTtwlwN6+CkfcysZj3zQN0Hs6huugAASk5U0eAh87RYO
xhrZjtKcwzjldzoXXfwoG+G2WX2CHoCRcv90jPYXUmXVqu1ILycEhVlswuZq3P3Yv8O06jGDx14R
rQkJ/REGs9bF9kEtfVHfffzsL2d8sdlD1KylPq1J/vS8fCqrg+rChca4kcHA816/9uvIm0lPwQ8N
iDfwjO0dSPG4/eJDmVicTlMS5Y7CNXyg3lV7+ybk86GfTM+5a+5NRDUoohdo4YAIH+6Tt55docKV
K8Qm+1WIhkaUmNFmCGoilAzQ1zI9Tps1eJXtWdM+g1cbuMKhfBS3HQYXDi/lD8HAX7hcQrQ18Ejx
BlyRPjFnNrd8Mi/Py+FQNdSzxCAnQOqHDkozD14RlztLkgGqmIepyWS+/k5AvyTGZnb5IQlhrv7V
LEbT9Y4JLqYTHyfM1f+GZ0prfwZdJbO/ZlDgmSg9pUMHlncC/zG+IaZyLHJrkKf7I+P24811q0um
uh7dY46GDs6t4I1O2Hg/bfrxe1pmGeyzfA6dYcOuGkGqYt82rnmlGOjvWgreHTQWseUN6kebjoff
AtV6WynTkDWLKq8FCM+76Wo042mWEWOxEeuIMM5hUmgrRJ/7JecdGLyXheZgzZYx+dVG3GyiV+dS
ERu0c+RsYodpFXIAfYXYAOQW54BwcbmtAGshPrren+yV8w+6WrTLNBYGrE7sTMKssLgxdtfBNxak
KUmakfcbsY2wFc/tWV2HaGBZnIADLwJfbG/m7nFIhwjj5FpuFYg4oZipmnKhndGAipb8hDrqCLlA
dm8lcKTgeKlub+aqY2i0TKi2ylLdy1e0yetKiGh2Ph04fKlPqSac2ZMPy0d770rDxstzgSozoxOc
L9nriQ7jDah/AwanU5nM7vh2SI2QzrHLfd0EVrCI8H5yvXMcNwkWUoKfft+AHqYSEP9sZJ5yWzuz
CUtFETKY12AkHwAx+9nLVXNpZl0tQgZojSBabrfcF1t7eDAgi/5UdX5SQ4CTvkMsFz2++U9YUHGH
HZrqPa6/NHsJvTcEoQ6nKyFoNzTYcXAagLYo5HWzzsVXas6wm9v/GdFHLelVqPFFUu6ZKs+SJzmc
jcFdKDTAv2MS0phrfo4w1YYaW/ENY7fH2nz5jBKFGnW9PDFWgiB1fuqfNnkfLTqQGpe58uGLgdXr
IRlLosDB7IH2cf3iS/4rkiW1JreI+sOgHmmSBlwKihSspBTArO9sKjK84awj9PrEbZWOgA4Yv2nw
7qO7Z66NunIDXK6Xk/pz9Fey+ViF+2x1UKq0SZIkxozX7HzvJMvw0dZ4nCHP9klwEFrDTo3tBEyx
9FHBduPRlHZtX0dBTa6+/7Z6e9MS+rjbohg2et/hV5Lrl34NnXDjsTJR0antOWXQkND5YLUEWD2Z
D0Sw6BCaRqB2IEBzxoC8wrb12AupceBILJQqrrhGXnnpseEjQ0gYH6juLdrbzobVjDmbIw5ja1SK
Jvmm7IlslSQeuYNsivagMCTXOAFNySlrBJOqm5t3CCRDasBZpJGcUeRC0TvH4FZEWgDjbjHf5xT5
tNoLWfjReXhe2enOqPtD6qmU4a8IwU+qWwuMr+6c7/ALYdgTaoXVLC9Qy0N/aiEIvV3ZJk4Qy0kp
zm4kPzK3pyqjg/Xi5yeWKvEptAd9jm8YcAYU6K4/xHuKdn0JNgUF0K3mizbhyfislv+FR0c9S3aJ
qKnlpy1ePq2NvxA0u0o3W59ppB5VqrSRrC1lYQGsSmGLsdWs50Bxw0wcPu3t6lffOggRKvQG5cc1
xNyC2cxCPnkE1mImI7UJnT//cWJeQ5YVaQ+ltnRvW4FVDxSECK0E2yuPquVkw1kgw0rsrbCAYjh/
519DF3Ss+fhfBM0UOpj5FyJgpYjPh2UTW3p+uPZbeaetL1Dm0bBW4Jik4J437FKAX3AwRvU3usnZ
odY2xwDGzICEaBNac8tBlIwcrpOKOupiUa6kqEPv2QgsdaofJwPQ9Co8PL8/XvrhBgRTlKJzfYlN
3+Gs+bNjrSJFoDHQVcAjHZNmMwF1MSo8t3eAc1N6CRim7rdmNuNqIVKKYfptX9cCEH5dmZbrcSoW
14xr3PivTENNzhpjBeYrzuOCR9dkfHshmAlmwLMfs9KR7r/t3/na63i3M2eWYn6B96mPn1lRiI2f
Q5d4h0G8caxYbcNaS7wcreT5dVB7Skbknpkxag28bO3lAwl8vjwhBJvR+s+tpjsSEnHAwMASArWo
Af8pA861c3iL2jG8BzPk/sNJ/cPpE+dnJQ9HuZkw0ROHwp0AHxjHB0G5TBWtvWBPAsphz4MWDhdN
uIYvpsiIm0gs7UlQW5RVlOrCTxC3CIPP6KAt2apnDMNZrhet1NE/c1SyiVhrD3hYVi38sHL7eRsP
8dpzNoZxK2j/ZsvxTyfhOQqv87HksikEtYnXhJLfUVgJVoJPYNP12tLWWDTXaeSxIZ0pkk6HhACf
lc587ep/HGqwhOPrX5JW1rvpgbz/S2jH2ggUcOXxYv9rplMTry7kM07vN60bBnAl4ykO+K9F013l
DV45hutXuswn2NZmrigT0ijLHpxfY2YfytqOJBHfuPhUq1VVafTlir7XvV6C2lsiJ5N1fz8uE5Z3
5TMyvcV8/UVyhqj0oi/bRMqdWEPbYm9BHpOUCbkOM4UtOz86j+jfpp+0+aWjw+BGjHJ4Z025BoR2
3yD1D5oTLGgJLMQminiLzRVgfPwcynzM/aScLItpLue9zr7fIcuum3LL5NXt7cKP6KmIK9YGZBzC
f21Gs49HFaW8vaOjcXN+mvENDqRrApI8s8KKA/cQUuYzRSGRAEcfu46Ot/AX7V7KIkCchrO90Zp4
76pL0+yGJl3fMWUR/Edfj1XaC9tVtgsACe/LPK2yRVjQ/DnOXW30bM/BrWk8XtJKU7BY51yOjHVQ
aDNFO38DViHRr6b3xAj0fYsowCFTCQNB5NAJwXHJ6yOFPrfMqYTexd8sco0kvfobANLwbqM0k7wg
NcI1241ypa2/mxd30cOFRJTat191w+M7YUqvTNYnIJ8PGJBo2vwoyPEptCtPRbvjQHvOtPXBB7+9
3mMlM4uUfiP+iXJ6DS7nKfA+c0vY/iCtPhUq31MHqeAvywQdFiptWI5qu0bVk3f+Kg2XCTG0hhLZ
apWfnLufm5E9aq7nbDP6VSj2Yx88/yy+N4J0aVKF5dnsYOThv6viNLTGemND2nt5GN6Xr2koQtb7
2GHxBUDgpLajOCMdHnxxILgUbb7riibwAobxwxHqThLZlPbrq06cCTEM2pZu1UQznnGv+38mGZ23
57ctjGuk99st13joyjiHZnJzVZ+Lxh8eHEDN1D2tOMs4CQF1BT9gwtHEjt/r4WjUS/ByLwzXHuB3
lxaNMoTLqFpTv3ggf7a1/EgLRBrXswa4ilCUCa86vhLOxXd2F6vhNg4ormg6bnpHQ1mXGViGIZxj
Pvfu6JTuZFKURM0WzJZhrmICtJCrbN4leiaqteumHTvRhkNAXoZHgnjKbt6uibMIeCICULbGXwFj
geg0pex8zluL9vbrFQcySAK7ZWgpKD9XxTTJ9hGHuxvGNtrvOcO88Ynqp62UOTpoji5o+00QGlqS
ZtnrNJRBNhjxdG+kOQlt+irmPiC9mfReMKuX7mXP9g6rQiDhlI+nEwy4N0t6uWTbTPOOUh+57SIy
QMktTp5jJNDR2YWQyhFvpl8j4T6dPRTa8GlthJq8hNrW/G1KZnPBFqwLMC8ATsuN47Zq/gIhTWhY
YwOTIT00tqUISxaQL4+86qzBnEy9kduZCTvtKIPO5mSvZI5PoP1r2KRC+e2f9mI1PwnEPwDwBq72
mbaud6A5bwoqlOUziBn2p4Af0E3/5kB8dM1evVGZPjeMJnkeMG3mqMa0wBb2gEjJqGqv3wNXOT5u
ZMemPLOYcbY+FFvBYL8Ae2N9n6D1s8gpjqK02yClzTWc3U6L2L6ONNZkH01Q2GWRveyCRMfgm3pg
iC+Zt5VBPSmQ93XxxzOvmI9NnYlR06hFLgm16fgl1qrBpAKeUivMFiJfvBbBYuB8vGTUlBtMPEmT
/R5WqxoVHHJ3yKyOblNzOPT53/6zQmw3xYuVkmdn58DiBndZXnI+r9sg+Bvoyy6yw/hKPWIG/K+b
57lcS1tDRGrSHTt4TAj6aeBV/HVbNMsZihMJ5oWf2DXUYNQ3Ogi9hRY68/c0sLXcgMsU30Q/6lYn
agIVv7ZyXrnYDhXSE5jL2eN93n5XLaSPJ9L3EnwkmuL/7n2tIUVIDx1ervzve8n4X0Co8iiorOS3
lIEU9o+SEnCdvanokQjH5//0n3W/ihkCKc1md4humDo5EDrl5+OCc3WK0wjWG0RkWyA501aNoqY7
XzPMWkcZSSIcrPpZQ5N4+zFBti8Sc4xct5bI4lGKNG70g2OrOLKnbQwl0R9ubkr7vcw1ZgaUns8S
tvPxdB8kTkJCqDCb4iWQvbqn9N7wDKm9sKtLgMiqwqP2pEbMUgQlVEyQLyQierYI7wy7jw5NuPaa
ArgSJ23krt7VDjiyi0h8WVRCBcxSmZs7qnokqBpfYmHGOE3GPCuck58j3jT+UdH1ziXu6ZVr+XdQ
pgZGVrOneAoQzVAh6/l7pgQgSaXGQAShQUdMchAvFmQKXfgB1/bEeRjV4oaF2xmGtnMKk+TEd1LJ
WHQHUvaVlUQY45jluO1tDHh2qkGylfz3MB/96yWrhhnN4ObKR8zFRi/fs4i1LOxZbAkimbjOuTdz
dPl51nn5eRgTbZtDQeHhyy7ybBaPNqtl3TkV3R8SuZXhoTRt7EECaFUuwzcv13Fgp4Ll52tuPOzl
HcOCjiqmbTRU0dOb8HLTH6ZKOKHq4UtMxsabVL+tQMVaFGgsIfTrLoO/g7zMxkhy8W/+jQKNbw/0
RcLVNnXQCZhwpQZPRGVyMDF0XWDUdJWs/1PBMujPJBi0Elg9Tdb9MrIf7+ExMbZW06EcfCE6tE65
muNdWlTwl2YT6NIi5cMximpE8bvGixhRCVf1FraoOaIfdG9rKlOb57RgFb1EyrAGDJtSNuBjqQzF
eX2gAV6gdBbc0qVnQdNR7byR5UrqcG8Z94ug0LaAqvVExIOcqafo4pHjGR03jkcNyJiQeKVO/BBd
oW34LjlO/q7X5d8ukOHZvsAk2GxcVpgUWPKDgHvcB6sMvDdSLPWaZlrPMvZiqdau9HkvZf8J+8mb
4cB44LmxI3OGQrc8fFbijHnPjwSuBOihyV8eQ7oVw0YGTkOR8oW2v+18nGAW+FWmFQwYsHa0PMFz
QHh+X25PrcgeU+h8qKr2p9Io1iTtxRM+Lj4pOWYD2x5Gd5YBaXA/80NA7tP2QibUw3sh2fq/69VK
7zplNCsHSBgsHDvKqL8R90JSG5yIyBWbhdvy0KCqZyLVq26YKOHq43SDcoa2NsXhjldEcpOrXTHE
i4jc5WCopqY/8JJVbaiiOD9t3dkM14VdAMF/xenqTDJGvOu+7f7cXcC79/oZaI2liu6Utc6T9czD
TtGVNuRer3QadN4gnWzsXAzNSV/RgShpjitW13Ks8OP4UowhisJRzmt+wbNXy/6TKZMpodSfcxIV
w+WOixNMwWwXBDE+4FanMirUIy3aM8emhzNcDS9x0bRJY1pPwGt7P0EkF2d0psmlCFCcX2YvH2PV
2hU90LayfX4aGdBfqNKrPgGujUhoSElSfNBL39vlFWf2Bw0kP6QobHOypibcPRx5yIX7Uc+oYRPf
8lq3u7Zi85aYjgrlsHNVU8tlQvfqCYNco3c7UYzQWTjcSH2pzHL5xNaztO7lMpLYZ7Sl+2zuiUen
gQt1l4izRzY9EP+qsgBuW0EayrRC78zUsdvy1LSsnKGDcW8VpM22+/lWe9RalETyMpWoOMTtyLDE
fMIMX8yQUdt9t+tM14jMjcu8PyVFuv4lJu1kEZJUN/U8jVpus01SBc0H4P/IQ7JQ/svG7WPl3KWo
zs6NkkXwVJem1RDqQP9WZfc7iIY+euOa10jIwidMatWOtcaIS0TRhRpvrsfxDMVSEASHGZpf2C0C
PrE2z4VF+e7/gH/6xYjghSh+diC9GhcRdpIGdh2ZYD2nSB7NHfyDnqwKORQlOB1wc5tlngiXC3fi
op+4NIk1l4Ljy2FbxGMwFXmpBDEgayGkdjoJv/GwyQM3dawvzgr6T/syRKVVdHcTUa5gpCKdkDd8
Z9GWID7ggNEsI8aXhlbMUNgoaqiA4ftCd5TeKl5xk0nEyV671+rAe9/9chG8kOUST+CJDQItgVqL
uNuNJ4/ywdXvmp/Pv3GQTF6b94MUHFDhx/+b9sDTp2qkU8HzwASTE6BioetkwkhMQedE2rNDCDDz
eH/GS2L2IeoX3pBHSoBduRq7uVkVBgAxsZrDQF3c8HCEyeA/gI5Nz9lpWpEiyAWdgOugnlBnKTl2
pktR0pWRrAsPuPch7NVwH70clx8NAcc8Ht1A/AwmuOumv6QDYHRQlANLPRpIJj+EeFjutLDyB+cG
yTX3EETGKg0aaVNjkzTBb8NhTUAmjDdE7I9JrcYinhkbJwE581DpQGA6rQoXFSN4OoRQWK8cd0+e
vJg8rF6P5fVd4wPMFFlNoYDzjA7qyDP0B0/vLSehWwn++6rGgKYTValcYsu13V/+JCMs+6AZLh+K
oxASFuPlyTWtuSfVpSVNm+PpOs0gnYSQSLbtnMj4dalSVTxz9sIHzrg3EwecMu/tvY7Q9MyMGGAu
Rr595njGAUPTbDTytiJi0oGYZ5eAFef/fEVjFshzVLxYuDHlAbe6yFicj2PvNkZsFnCQJ8Nsefg/
WrP5NMbOCAZT4PmT/04cn5mz76ZHP8qcTSMzgEh41c4BCril7aQNSMC/UCZQC9O4j4sjQPXPqgxS
ACEQNoMH4f3PQc5SiZiVW6ccX+R4z0Vq9hBJEzisa6kvEzYkW/Wqlbf61uPARFB9HSHkzg++bkLQ
xkfpEX4/prUjDn7v6P5swLbJo0ykO+226CKPQ4WlyYec9WIA93W76Q9Sal3E/ROc1zLe8SWp09OA
7D8rUQ2ffQ+I0UVHTCuM5xQeatlNDbo12C95xxjPIM/bvoIgtrWGWTvQjUsCUEG+i9SMtUQN7vcO
WS1SGtwJhNiSFV7peymB0I2j1R3TQjkUld9aPQOjItUl7iQqaReXRipI4cufGoHyHZbIbPn3j9jK
S4I59lS3QBS7L7MX4DUx2XGcfjsK4ptcEeUPphQ6tb0VDqM2EKydCSpyGKNa4PW5zy0jv+eCkWdG
9Iy6ASLqyP6eDFpcyS2nI/plLHSCOFJzIc2Qqz0+xdEQvUK2SAhtsVC9gdDJmwDtENI+dZ4Qhugy
wsu2Elx1qaQbOWum3if6hb843Rv5S6Me3MTzbVrbXhvoC1i2CA6icY4mMlUG6pM6F6aNQN5cGapl
qdGF9fA4Pm2McUnL7SFGt7qNQ3ANIZdkGeFgUsJR2s6mXVVPb+xBrH5EDIKLi3lWjYmgYmXfki8O
HIgOzXKlCyZb3o5yHD2deJAgTxXQ1H9qxESA935GC0qnDbb4I8xmVxuekliBwI1Dgv36hTWYQvrN
DK7TNjABOB+HBOH6czWEfBY4U9zzmimjOXqUYUYBkAxb4uWffR38pm4kgoGNqo3SUNYzQVvD5iuH
Ef913ZUARraiCo4wG33DvaF/vAfpkHCIOhxCk8qDtr761lo3qPvyqx9mTYwerqF6oj5knyPh09AT
j1/xI5np8/lAgyzblFDnL9KORI42l3+25T+uZUMuxv9+XYsgaucxNNyt7l5z9zSDFZqGNh7LK5WK
ddV8BWjrCtouZeg+s0kAljmwlgrKh1GGnAz7zty7t2tC7hCpGLTCnoiYLv3eI8NKdD/y04BYdhe/
9QaIl8uNQqEJx34bFWE2cqh4aMes3sGghklqhg+4hYPheEwWkXxvAa+nhtqzFLXGVqFV6NRyyt8D
BjlTe6pd/bSTG6DPsrjuY4jfhEs/0W7hXGWu0JLA7n7ZWTQoxQfw83PlJ0UyzcQU2tHr+eHa7j8h
f/dqp7mAW1R5tZtfM5t6ATmzZF4dSdLjsaX/4uFr0TsZ+Zj68hZV4/C+w6IfFSjDfW2YCrmm5hC4
Ha6jES4cJ/JEu4WQ8udXEWZ9pfg7e7/ZkQA8iSgcPRYTEFwa528/qfPYRakeOhe5uWHX9yNiNdba
vrRRm9oXM62zYiy9LUYRfa6qmcDQAloy9AWTU851QPO/kDSPjX/BdmvnbPau8ueT2NVkAbqVXdWS
NTHwVWuUKIrSwcIbadE6+/2836xqRyGoHVSqOVy9j1yVuAHGamqoiCTWZ5flwjaxcabLbXBTgK87
M5u716Sd8awsfL5I2egzXpYt8pAXRiYr4udGFKkIxNHTHXA//cF7ql16YHjXgxvyoAe2ldABDlET
YjuzNs8itUhflrZKfBpGK3Rh0l8RsW70vHNRpmdnj2lBI83oCcfcPMACi8hA9Khf3xjMkfG8onjA
JdhW9I5ph7HPqvYCuyjNEINmDi+tZXdR+oXsWh/qb74NOHf65zjgKE+ZA+ICsWDlghlOMa5mzr8t
SgDClgvVu5/UCcOAwz5xNw2LE5pnOatqFNrJKlnptL1W5JcUeteLeoa/EWSyOvRUr+tE1QPJmDu8
OFSwdgA3b3AvhgJjodGJmI8sIZelV2BXfrFiQ7PpZbgqS/zx1FhJ6C/tkpDPABEbHmO4WnERiGOW
cJRXZdjn8ejzRX4OhNRWHzMs6Rnjv/cUbyf39eBNxX9DaIufzH5eyauA2+r9txhlcw2J3a5/Lq5z
oL4JAGcY46gey8ajNVSXIUVmxtPErzBt9l8cmF22q1SDUcdCbIOhVmknbdpjy+myQQ8cjKwaHN7y
p2JRxrg8tXzxXoES4Lwoduc7Z7xtYzjIa3lw3wghgibRHyFejFoXw5Vo/r/V3lfT0XCktr8IC0II
Ary6lDFA6xDAcKHcpao3lFxMwegFabnAyu4WYNIJxd1E/J1H4koGu3byZ5q+DSI6crL+WYwSz9aJ
Yx6h6xZ3qIYeB6rRl6rN9Dkffw/qMH02UkB61EQNuGk97L4sMV1b2lp2cmejZYPhP0mk4n+aVEfO
+fMjnG4Gad4C2bP82OO+VDb4Kp2JD4BbRedAwG2rzQjTF1rWlkDHzgSrlm1d9+G125aCrqg1BuqR
2xQCYTodKSzB5Q19xr/ud+uQNJ1jx+LHbpSxk7XgNeDWPAIsUXT4wzvLOQ3CUce0hko3qvbq8jxV
1lp4ZRfUdSIhDgDKa+AJsSAsgdlvGZaOpK2iSlACPmJzKLiQ1Wgd3a2gAsS+pos2CnZfzY7zmFYF
m9cZK/TkjWODeG2rncA60BTh30GdPSEiaSq5ORDUz0gtKCNqcHB1S1QDgCWfaWRqFdMcfUPhuIIc
J+P9RW2vrj2U8Woh1bCP3FJ/NLTGWMYn8/57UeDskTguNIv3J2mkVJzL9T25YFPOy2tK0pfBLz+0
eSoN9+UYpxTkxM7AouCLd3eigpt9WZ7YfZ/j+HxhrX85f2rVgV3HLgNjdUn3y5xIoxfWoNgmCtxE
1Gvg592+0niESFJ9/bl8mNMzlBFoU9UmuDw9mWjaugpm8OJXH3Mxkcg3nRvmG2ff7GR9amZeDAIS
B1PirLFYol14yzTxg/4895hDKDb087tOOnXVuGjum7qKzjpYJB/VUxRwPPGOKETaDEJH2XZBS2+S
+MFRbwwsJfxAcuW3stpOJDqw1Aaaf1hllXDfwrcQYb5PtwozlJIBhCRPaFP1Qt10viOQj3Pw35fA
XCRjrXklCC6g1VstZfzRmBTZApvr2HYIfjYCI2qGn/nMwDfEN77TrWGwV7NMaFR0KcY4cGEw3X+L
2NtBZAKSTIqOgzhHcZYvaUdFg57CXKzA/SNdVx4N/GrOCBrYBhABkLvkRk6M8VJVtaPZKSGXKAEF
4B0qKq+mVpVjqUfhv9V6WSb3OlIT3f79ZAkTISI41dP36zW7L4gNzQfpE+XKwJ92pElcrvrdxsnV
mzBNwbPQIoaBEHnGN0X5eqEJYhIavYDwhu3OVhQipMmPr64+G6Jj2etMECAkW5Yto42p1MyoPIFU
Q6KvyLp8OCdl3wg7cDrLDMQWhwi52JO/9UmpLeFOCUgcrERjNPOgQiU9nKY0aufTc1VFPWYN+vyt
DiSnPZYjluLZ5xy2ZWVUOFzIM4wsOA25ksZb9UVQlT7w4og+B1D78AAN0LbbFBX1/0r4zjU+DDRc
UUVBWTmQUcEY0X8MSiYgfVenXMD+jTpdbFTF50XTZzoOI5j7Uo8A1HVTTFJuz8U7/gYdgN8zhKMJ
9chqJv7x/DtIuLlGdM67uv74bL3rhaPc73gvVznEwQKuyznMwsv3DQQb3QCLrIP86qn/6QTH+b6/
whopWOk7h2m7a00IrKs9tPxPMgrYfs/oi4l5D9zOPakfz0M0R0W/NJ9G5ua8yvsO50hXUf7EKMsK
3KRHtIb9kyzdFOhTUaqGZiYQiy+6IfXfFYURw4HYek+qi0/KfzRhQsAAtZaIoIh18j4Dvfy/YGww
2XkMguxPEgfpcx+dt37YPIcKLS1CVr+5oez89Jg0eDY+a6ZNLDmST213+e3iJ7G4YRqeC3wzg4is
HLqE8b/POT7uHVVC0sAsviOZdPPVCDyeka17+NFU00mcnvfoC71V2fnh7s4za0RBBwUSe2drNdoz
sXCUY6vnax9Gz8YMGPHZA+ZrLdhrBBNJVOCelqT/NhZmap7UDuzSCFtLuaCRYwVKRQqos0KkUlZ5
BBMWHmfJo9nJPa9QZKKpYEkiLAYmhDNi3zCakmPti1fXD5T+gcnBRBd6rBqB8gK0eDgEYAxOsPPC
nbX8qLBL5Q+zgLaKIhcC+Kk7tFQsPkhNRh0jZE7GMCsQmNFsoUpCl6bLL63y7w161ssRcXyl4Mw5
TFqG6kQeR5vGaj4pFdx+6E6nY5EvApsH/dm6ajJfT/KurVG4z2IkQvIOacj86VtA/TPJ3HiLm7VV
R0rEQTTOkr93GzUcn+UH5+GNSU45DhgXLYHMic61n61DfFXYnLs5+fH280rW+PKRU+qfqPx8gJGb
f+SnocxoCrkPn6SUnaqtwMSQlJc6BLyeW4epXXLyd7TlhSBNOR+EiktTiyuKIT8az+G9MqsiPqu1
M/9NVTC63jHVeUo6Ww+HZ7ecf0ivowF55GYf7JQL2XoqnWqxnIwqw1uJnOn9589yweS8VP19Vb11
LE/L3ELXN9IRkTJLrDDUtifWfldCCBaalJqjD0cBXkHPs3a667Osliu5CulxvTIUx7jCM6W9BGJv
hDkLMhZbgMmaBbjrizJyIMOIPanDWeFAL+BP4gEQtv0JzXpOtpnSWy79KBY366HEck19Jqj6I1co
LSJGD01qLI6hM+Po7D4KxnDuLfHHiA8p8QGJqvkL/3jOD6h+cV3E56nVDnBehPw2uqYgZsY4usw/
a/6T3XYMOTauvP76vAavdKfuPDQkbvIoGLc06UmlrqzAMNdwBZoLmnlyYsxeuVLLG6EV/rAV7rIz
mDgDYdSKGQj/bf6tDK58Wj6zEWtG6ub0TKkNIVx4fFoSV8btGoGlS8MfPOYodF8CcTjp0fa2om+4
WsGVFZlGy5tx2cT9J/Dyzadw14WSwwTykk9S35HzLGwrjH70QJOa2z+N74Oe99iJTpLhkn7SChs4
Tr9Gj2WsPbvAHQ4SmZsTUg0k7pnDOIxotwf4goWFLqS4zG9OIw33jUPWv3GQcW5HCOnK22YQ4Edr
rR7YLwz/jRPFl7/BMDnCx5GHxWFuwvh3xO5BkTYc5YuXzmauQpcXVw6fifpruEk6KFFjmf8CH3n/
V5wXatc7j/TSRsSWz+QMyJlnVGkwr64KUvooDL/fZgZKYyuJ7NVdLIOIZQctRR2VOEdj4m16aAs5
5MnI9AznkUtRravhgLOJsK18dx5tSGglB5XargWVzc3DjcnvQMkc0DoTf7Ymzc8iIrx/RPmq4JO0
Vp4CROn0Yk2HcspkAY/gm6gdcEw1ZSg+EiOZt8BXZZ1hciZfOP8eY8GpnfIzGDQSWzcYkv1/hJkO
m+spdSHs1MM0XWYIGrnYFcRTVjOSHmwkcwxZoHGVOSUkgXmQIYFN7ftKZCTNq8j3+/0wwBlAoDve
IzahckY9ZoHP90HgfYhZZvNhqaX9pjlDHZg51XlEzjpfuXhq0TLWyuQDTiyn7Wwj/rN0UAmRHoaN
xDZ/KI5GtRO++/neDWdIbflmVJrKBE8e7ddAoFjgrqOmDNIYF0qETKqT2ZfKlMSaujzmZ2xoBCsZ
6hOGetB96v5YGH2aDK1RrKGD3gEUaZp6UUObRUCTuygiO6GEgK241AQzWxRojjo5aV6ecbhA3LD2
kKldaxA3CluoBJT4hLaQThKKRPPQhaMUkBQVd4sVCvBJrJJKFDJpL/4LBRf+iO2wU5pPYqffnAkw
NpmtKHwgjIll/Q83bQ1e8My+JAWpil7OIPKqU1Xu7ewh6aLGTGWqUSGvRLT0/jua2B2UQ/nkuLno
Hc/LwkVkibAl7Cz+dapf56JBeWL1RYLTv9PHJ67przU6FdsWCS574YbLNMvqLm4Au5nz4tnS5Djy
pQwvkeA2nahboGHtgTlgF9ziQVpkSMVBheRjkaYpkW9baCzc4H4D0b1xkK6vpEySqZsmcAV/NItY
MmWmjV8KTqGG6rbVJAbh8pHhbmTmgngzi24VVa58NgVm4GnpQ2CGDewFgsdMgJ45bfOzHKQnjTSx
k5lcA0lmgjPr80oNQOE63kZAmYWUR1tW6jN4PJNcMWU1r/8zg94zEi4q20gKfa1eLv2e0L3YXDnK
h59l4jLD7QYt2Z8qkJnnU4UryNnDDPc8rubNm8LQUM3VKm1mebGH3eHuKOjlvXsl4FxisNTrwA3H
yqyqxbr7EKxzoZ2dXr2kDSsv7kLBowziaoW5uTCcsqPzXugUs/lzLeFPiyaKZVD29l0wNeOfSp85
qhMhgPXeFDpmUHhTe+XEeFdWeVqMv4GE4VfLOrVTGhlHjhAcaUE5nBGYilBd55p2PpuR3e//GMo+
7UTMDH689jSHwvX857lR5zzf/FY9ML645UmFjRziNPhQnkG14xEIfCUYyyFUx+h43lmJJYaIMZl5
lVwBeUszaRAF7oy0s/HQC0+fuombkwnBuYQtg0c14fVr7gqdcVjV+yD84oxOAcE2TggcJN22bR9J
M3VvSb+SdDoVPdsGtwQ2coW6R/rIjWEneHLUW8eXeqTI9is5Q2kLreA6laELQf6epZsDmK+xGITK
srAIHublkRf9a2YrTBPA7Frulkw0SO8Xka2jVNPoB9Ve52hGVIdYRt1G3VWzKQ58YfPlYP6CavWV
ui8lMTK+jiIPmgTCIT8NACb/tuF2ii32q3lDIqNVt6Q5OOaqxdUJgAsjJznfKbTJPc9EWDcLxpjM
a8hWr4uyVccZ5kmI5clTnmypoQEiJIz7H2kDmCLKpCd06TVPDXbcfsQESq9afqf0VfHzKYBzl4if
ngvuLkOpGSsaS5mCYcLi6FvPN0O5ONboecJijO7wM2DJdBl7JKPcuW1TZt59UurtcVtt6ZGYjP2q
Lq6cNgy9Qc4xgo0ocYw7FN+f+SMGXf4dfsXNO/by9Jk4sQOIOcl+QDX0r6cjK9h8GHM+p7kBGhN0
KV3ViV83nHqNneLW/fW/+cPPJ0tVOIrqzZAR/WINoP+5GbSIp7l6G7P9RT9alSAupcQ1J7kQlI6O
LqQTIN3S9aM+atoooFzzOQkzO6c0K4urpVtQzcZwpEHg3uO8EjWHGjXJamnxMEtMKTTkFP7HhGtc
SFV/ntiw159NCYFJEGadOJf/l1Xi15AJ5l/0a631ZYNI55WgJCmVVYiAVP2vzmLPtvdiRHEL+Y7k
NUA4jByDOieG1ts8zUeIBdhSIITbsewRvN/R5FXYnQ7KlXiJUisEwAo0aTy8BlUKtUuR5zcs8mZ8
yIUWoReNHRk33tLVKrU7rKjCFs8DDwiqSANc8ac4dwNTofp7WNVub83WA/V/g5G9rEGNDWTSonq1
5myePp8PLlkn0DN6s/5hQiKqaiaOc9LG5+vRyQ8EG6zC+Vq0K9Z3TZi8ALtJrhymFS0q7O3v5mx7
2xyfjT9mBHokbmh6l8aVElaUr43YWKYMVJbrIjacHLLh9dieQvpdpaFWu6Q2PHbysofMSTJKjF9P
M2i8EsVgJgZD1rIYk4tfyRPLHYxpZIG+5wE7xbsou0+bPIDVyLpsFjo/HgWZdQ7bTj4Qw+LNLNKP
rtZXwSPXxJE8IzGr/YVpIOfu370q1K5C/UQPEz5dp3XvLx0v+caY+6rFJyksUyJsL5k2iIteQPgN
ClGsqlZTt7mdZhn++9JyoyMUsSPTb58Ekg4CGR2AKRqEDyAOiOevWmV4Fw4MBVI7hMiDlKs76omF
8Lga4pUhXqFEYXtUW4PQr5K8xUaCkTVTqaCGj3FAcpK87VMl1O+z2GrGivLXtWxTYSljDYb2CxsL
BRIfu3Ffd7r+8JnuAr6Rk86f/Qc40VhmaotUvXTwR688aoTsenzspBJGbNy70duakTEAncdd4Z2T
K3aNyjWpB9cDph0b8lf9acyrKktGtqfB8xNWk/ZWoorHsn6TjsN+dwZVhbarQ2Sd5be7747OYc4v
WCK6OCy+Z3D0Si05ZDTpJIlOjVgEQ9uCH64DpaujiYFgJzIb4msM4uNtG/kHUk808vV+N7gVR/li
8QGxrnPjKOzYUX15xNa73+tQJkE18jIE1aJsg96rQEj3EBN4dIaNfLzGR6cw6Ml/v92+Zf0Q2/ct
vjuYjPg4cMTFMgtxvr2R1Pk0w1ZSct7o/HZNdIB0P/P+kgJ2OCt5lGhR00NcyO0cn8cutKT2ivNS
uEoLywMJcZrNFf51nw5dV+r+m+rEeksbXi6W1Jk/OrijHTK7NbPhLE6AuaWrd2t+MBnhuq4YGcb4
1+fjZA0MHN++vzFjAv7YOAhVv1kwksUdQjRIupx0c0V6qs2d0ggjUnKwBjCR2sRnwBtFsH6l/Zjm
Z66RT2dI3qo0tZTDcC7SCJMe9zSLv0OaXPJJ58w9L3Tf5r3RHMv5fE7r7LYVKGybTAGyvQbUu2Zw
YZSrAwmgy9gLvNvTSnNhCp6NP6DdKlB371pPeIVkLiRXEyOl960kqRqTuOo4p8H7kgIR8BiqwFH9
WI6Aqh2cenp+L/s2YXf2lJeVnUAzpw17/fKq+qpPIYBN2LTF5LiXJf9pSYyKq3Cth29w15T9hVn6
iJJ3oVLOsFFuNAg4w3PNce5NebdKjWgdUa6QSrZ2NFqZe+wpnrYUFZRTscHEjL88/hMxVSjBNF8x
FM56CsKGaxydpTjhT+I0YAfwz2nAEooGAFW0SXOL1rjsrt/gIo0TBsuaiVW1j+mOt2sE2w02LPRL
HEviq1f1q0JlgbD2KAzN2LQeXss2CrBJkFPhzyzKNKqq/9PzpCQd40SFUsOyWNgwdOkWyCBdZ9JS
aQxEDA2B6URASFSp+6WLsMZuPWo71/inL22AJzCQnLwlPRHkpG39Adw/oLitzpAhj8ZCkeHn4tO5
aHmNQZwRGadnWcmCA0Gw8wSlufg5dqufuZygq5V6yyRiqo87r9vzU9dZa+WoPk2mzwxIPm0s091c
yVsePMD583y8J/shDRMeyB/myf/641CYUYv1ugXuxrxiS/h27DABMLHe04ZOqYZMeXXizl4l+dvc
4EC0oL4o4BJQ7fZ9SSnfwGc7/ehIgUdiwOotzNKJJEZK3Yhf60m/8tgDNHxngn/ZT15mmGKh2z+o
1upe6QPA/Y+v1W1cOCkL0nrNFdtMtWNI8vXfgkGGVrMaSk+pDODOSa22XmM8y9o/QuP4xytX9mYK
PI0u6Sn/tBDb0PdaOws2tzSazCLiauBMnTfqqsQZr0+ZRXwxENhTtu4fo1fBPrPWMLT6U3PMBm9i
ktC7z2KGN8A6rFKSXMFGV3NvYBlXqZPSarDGdQ9zP3bU96GXam2iRCsWqKYQsaOWDUvKuxWP6Pdc
Zk+vDxIhGxxotK0CF5O8tyS1j1BniWLW6RAl/3DkVHfk644c3EcAqS4u6zFxPlr7Tbz8gBxL2LQm
ugjVNUzT0/+LlIFRL3AeyBeNrU3wyV7DE/b0k1Iw83prEKXhkleWuMvfDCDb57ZWOtCOpB/UN9KV
D7iPNOtwEfT1M1HzjJNyjfp7A2f9a+wUDoT/tYKznSNrzkW9nUpz+nN2XGRcCtlEdOJ2SE+CxfkP
SCa0T4qmM0MMd1LYktpiN2I0ITfkMdH8PVIfS5eNmeiyISTEjbWirzmUG2PDHw/vlk2PMcGFbMMQ
/sIaqVzEy4IOipmOj6t//X0FvsNJn2q6K/LTiVP5BeRrM7813sARM9juIIeHnHPiglCt4IyDuGvz
FN4NURJGM6TEtLeO7ElkUqN4YPTTyBH35ptJKdqGJEexubML/WfoW3msfWKz68w1XA0xVk5jXV9A
ZsPySuXsNiDy0czoEKBGVNPyZCHOeZ/jAtS6mnOUO2lB1TiCTvvZrJ5dOKnPwxSAguCnX2GCAZ8t
EixmpEKJ8CPxTzuaDlPFGpLJBiF+boW3/KYpps5zw1LFZGdd/cYdFesae0Hq1HOMzZwjQ+ajDssj
9DodeinlsrOsbSvhCD6QQnURM2gO3J6HKUewF6k3pXQwWGPhDsPpYJXH3FCwGYrqIlLA1N0I1DdR
cTrqprlz2+K1H3JfCffoGAB5cTy9lcNxyaZ18Yb5xG0UTk1lU95wv24CX/NGRTrrFbuVRSFTA+Mb
mIiOuGT+WuibPU0xtUFWmKMyts5LOGkf8sCD/xaaD2cJste4OQ5joPR/EcpyEPCZt9Xcs1K1Ao6P
oLGo4kBNGDdE9ZL+rBZIoM1h/GsO6pNIXAyIyTtFpDxgMlwde4JS9pjCnmM6CfuxFv5ccEAA5ES9
SmhNTDpJ8v1up31BAmClJ/akhXEqZUPMd0rKskaBkRA7I87h0XD+zrlVvWkCfO80te7wNNb/Tcuq
EVsDaz3m5bWBuP45E7T4i8XaKWyEwKfXVVlQhYDWa8sbodnsqc1Lluhg9mdoTVM7BuuRJYEYB0TV
O4p23s8xu4NbYClL2butZ5n+2Vw2KymNo9dRLJ4dCPCw7genHYyXopVb1dI8XSwhbfaMP+TPTbsl
f/jiSkGVU7iQNbPIma8lHer3So6S3pOvsnljxllzGatSZkDeAoHqAnwfM4qnv1Ug2Ai6W61iD6Rg
ssh0N7pRWEp4WWNTruPi5Wt7e4XDlQ/qwHoXpRexMC+KA68mQ49FYyqofsCou4mu66Qf1/8QLit4
awAFGcfL09UcDsBP0t/RarZPw2kswGYfX2GzaY62ww05Xk6MYog2RBbjm395j/F9kEMK+yycErt2
zi21rq1vGz3VKyQbPc2trgfrjAtCgHgzceZIunVGM/6xQW6uRi4EzZdD1FAtqM7NGc96SYFCrzKR
rl7tOu5+VDwEdcmaZmUCaIOzkWlAlN8CND1FaeM7t4Gpoz7S6iJXcUJsrZETCzgUKujUl9oA/dC9
DNnjrG06sOk1fwUZULkiF/YWExm5+bTLrTX2P42iqsTIhodmducrtMwBlG8mB7K7SOvaXa5wGrS/
tSU8/LO2CAse3lqOjVfE6aPR7BK5mstDQnaW59fT9GwTlZfsO6ZSb/bSAtKiBZlyWI/B1p2Dgd+6
49PZrQjiYEQCuQBw+/8hcNcIdA9H1nVubvrpSZqMOASMs78djSStrFCiX8nUSdY04MKsxMjSuyWa
Hy+wSv6LIP1MJD5NfdVniawKayeSFdPnTjk8JjkcjoGgv8Rw0usBgWFhDrDF3ReiKchi+voQUq6m
zRSVTtrFKPwsTrmkjRgiVZ6/rRCCC+mR1/s3PVXPJrZ3AhzjT0jwMv+Hx6oemvViABuyXZlMtBQr
RtPjitD8dStTdFzTgii4ld+vEGLDKkPjfxkOr4DxcyZnbQtKTxh9iWbZuxC/tHv9uQ9R7i/73ZRI
+7OnnJC+lT4aTT5xZG7ajrGw2JtNwruXMkN0P6C81sDf47/3abH09fWiIeeVgPoK5OvHh2GFqcFl
wYdlrlcvZCbm7lP28nDQK9d+XgGiprCQCcXrYODgWqJ8Qu8jVzX/VVthbyKXoJS4XXMrPnCUnj6Z
GLbr3AQ2NoVgOPzKDbPcMnnQt5jJeXdg6qBl7Y+hymhqW+qVJZnU8+wx8/jgv0uk6/J8pcNRV12h
l1Vjt+haAKdx1BEkfW3RauaOjelXPYro7itTMkURO4rzClkSwaTgEAlQgprN+gEBJem7SsP/WLFd
wEW3a+Snm4ZaZS+cND62x2VNHXHcwkTYMV83ZFop4egp9RagfxzpY8bcwZJRPXuh6kSO6wKl7ZoJ
udavoRz5s63e7BMc5eE4VTrLMWR+hRwHKYbz5k/N4V3pBuHhJtJJ4dzHILgN30hNNgzRescFdHVi
rtgiFFoxR11wmHBYxKF2xok1B7szgshmFM48FNXgFN3hl1SsUrwFBnw9gdY7K4wx4vwkWoVkGj2M
z8E5S3nV+NP5yzNPrxlPBC8jzYCVQeL+AMrVz+S5o0SAhVmpV/ogOXD7Fp1H22O0eHXIHimhgl0k
o+z2mqRD0XiqqLFSuIWEinE2jam1FGWwV9+hewIom/O0UsAmcshFvFRwScAfjn0+BPbSnXiojNse
xJisY5b0wcboQ5MGujr/2iBEIjhnVyDDMsFVhnQqqnPJGEHRDPr2qszIqFAMy7SQTlS1dS+dhPvD
MchgvsAvjVDpNY1TdDtWlhi/xGCHS6LEEvlXAFnRwFKVXh14MIeOGX4020tafi5+KihVT8KNTpov
gMHcTWLneYpZGMOzgXYznJyHXjGjzUcDhVg66FN7iSIWhteZX+RL6NLmqHkRR08XT1cNac+lUSos
1P2j+hf8i7E9f2oxAiFZrVCBSto1Mt+kR/inNOSwjQg5oe4Xw5ha+G92Y/ERNwTy2Vx6lrrR0chh
m8tI4pA+Slr3344q8wQxWmlZr5VbHmeaJuy3rDjKnLGS/wRqea8tqVTEtpFZBvy/J5Hg9C/me89x
qYtXlmLYl5cpVhRmNEyIrJJF87Kd+M05WOETPl8WXaOT/TOpNnHgak+PhdK5oisAARpgYO6BAp+u
Q7+/x5p3HN0TZoNNBxFgXe1UzsOMRT05u5AwqWr203sSqosPPhvTIUuNbHmOk0VEQvqXdoMsHzRI
zvZZjWvOKvB20Fyk/40SNJW8O09khH0Olaed9yayy5eqb0g6sME2C1C6Q+uEnX/nbGBZD8car1qG
CX/DxzSeLkJSNMMNzrZsgBk9laIp7O0siCBC+f9wIs+Lorouuzoz6NfzpNX79LTYGIkj6C+yQEga
I/ArIll/ofDHDkDL5vEhSOvJtUVObCOIA9BidsaIWp37ZGwwkJ8vJBJogorNT4oSoXH+dQZRnEhB
Rn4FSw0UxGvxt4xeDAPOkCyYvHUgd8YMJJQKzg/XZ8zO9O9IPgD2KaxbPJuKdvQJf3BWh+B/I9Yc
rZZk11ALK9fyliPmdxGVS76XNdp6LW22mu9POSH9VUtaxALuBLf0cZzOtWYt2vOV3crCF4xmzTgc
1A+0CJ3TinDCQbciSR/2DLW91offiqU1V1ALG1r+BmQb+G6S3Rr6ld/LegEZCEIUZzoLTmVC7l2V
64gL4YsFXAfQpAVLOp4ymClDtVxppI7AOruWYC92noU+LJ3FXRf3d0pFrjQ4dhMWI+9nktWFAIBH
OeJnxeNjbzSy3tu5VjqBxkyH67AJUHWZJD6TREXXpxu3TXW55ZC86qcBp4mkEpGctYfykDOt4hR1
MqkkwpdOEeTIYK5TCKterfih3Y4Z7VJhcO+np3XEqAxOn32KucXQ/FiQoE6enXwq69skahtmlC1S
tQ38s+mzstvyKht1OfCDQzsMVBivlXwKGKPqADUqb4Wx2dNSekE088pl3icjtsq3yn7vAP+8MUPS
JUX789nuqgtp8+fmAmSRLxY9/f2D7IAB4wWk7jUV9NYzQawxOxEyc/gPaOCd5XiA0NPC3Hrzr9d8
whFuRS+0GV3geYjqyqwSL4MpSZhuH/8bu25/YQhj3lWhat0gQwtAw/9UZqRfp5qJRgSu27ug2GyC
79GUua3PdXvw5gDcmbudddqK3dkPYCkOyj4FMOKHtpLn+0VTVOUVx6CyaLkG42fsVllwmh3OxRUM
JN0pqQ2IudTz185Fq8HmPzeqAfo7IIb1geblaTvwVFnkqokV5uUAKi2f/dlf08pWqgZ/0yxZ3qFM
2KK/riEhKKNtlOaGXVW7bnPP4wlVvY+KeviY8KjtlY8o55qhJ0Gb93LpQMgTM+6jQTyxMFvj7NDh
oMxifToNi8yajo0X9iOTeS2w+nd0eZgyRDSGPlL3eSJkGfWrgREWO39nuD+2r142/QAW7EiKtkQC
yhCOwbXQF+i89nWOp2deYp1B9fterj/RRY//zQYiA7N6B5yjo9u/foiFZc2sG5L5xN0JrvFkC3XV
7jljYwzJf2WAaj5Cxz3q+tcja8zLqIHDUIeaaJtcrvpsKCi0ttOqTY8VjE47W6nfi2for077A63O
EcxkgixxzAuCOo67nMkkvDD+H71dXrX6WmZ/XoMYvUTlCKyeqHwEFEVzegJwfXY+bWvzCyRv50SS
1ai/YsJn+sl005jO/2I11d+7lbRNx36Us/A8+lEglP2W9IW5EdT8XjxZRiCV6IaGOy5wKPmzBaJE
N81Mn39spIZGfbzgG43CSyP9k6m+yFvtE7OGqMP6z+14P4SJgtJzyq+Op5gENh+N0SaxbbSKApkV
j1w/rwbWEpduftZtvsa34Si4Agx5auWujpWibkdJF6Wj16sNZX58c/cvUsev5ZyWp27XrXchqGaM
0wy23Ul4BzGj327ShNxxMXlOD9hGWQD60jUIvqtKpl5xmCoUvqHQkKF1y/B6Q55snQMypSq99rAY
kCScY16hsDDcfabRH7ixB20VlmxLneCcQ6WLKMvjT8r6qeQ4c+tEfCSh/21cls2H4h0x/eDy+ADK
Yd0b7Td2oSWM44wAxhaLdVTsr6CWzuyjHqjwry0opHljtjvUcjXSAgj8f+EoFcpSbiZRVERc/Jqb
NY6E0guD8b78ot439h8KmWXGXDXu1O0jValhvC57716or0aXMZO/u2mw3MfNq7eUwvBEM9h86DpN
Txo/rQ0KWOyn7DkI20qVT6v0IroocgTV9M47/uSOswMNTYUhVco69yYG7eF7LL5u2vrzJMmdoDNr
Jopnn9cxNv+p0X6gHudk/71ErF+pElel8hhk2SNR/cpXuTVVZSehedYNkRBn5umrGsJxHG9Zx2gQ
k7DEKrRcc3Ui0teCluz9s4k+5OT6dissdkEOI0X6hj51XUhGfWmn5C6eR94g6oK0jNa9grss+8cZ
tShXrudsfKMKfO2PQAoShB5XSN7Iacm395V0aYHL43lIF+x1LyMzqNOmWqDRLWDa0Ep4dInmfGeL
Ghbfquy34SdnyR4KTAu9eLw2UtXe2OIVqovqfpAbIhFGQEauUVjyx4VVD2gKP7ix1mMXy+394G1j
JQ9Ao+oN4WpmGONdjJlDT8nHb5oMQMv4HJTD6VJX2d5VGJ4Nsmtu9ppRnIkvIIDdBsF+/79EwqOm
dD3hOhW1GyKKRE5rNS490IAIVJXYWkjgieLr/QoKvSk0KhW2TRnEHhWpxy3pItMMISXdjp330Vly
Wfhcle5+4HfRlX4Y5C/znweJ6pb4+7YyuTMQW5koQ+gYiFsw98Jd0XFnGh9Z6kNN4Zoz252oVkBp
tG8TG8iCgERkj3jIZZBVJUnJJemAq+SfbR/d3lCfKMbDWtR26O1QTSE73P2yMW9ZD7ZB5wW9uHRY
4UVYoAXf4WwUfJcAZiuWFuu2SwdNr33cW0gmqUNfX89XJKfMXsCg9l5FCkke5Rhe8MDzVDjBw10J
XObfk8MeTnO6NrYtP9PxNJ8FaPSsEM5pCaJPGaz4r1kk8P2Iaxb4yYURBntuldfDGJ1bIiyObstT
5cphbbAN0MDa8HHos8dGlc7DrdMTrvDPBhjzAZ04anZi/Zn50G+qPDDFKxvbkCagETO6hQProp69
kMEn9MKY8EPUM3oefbzd4ePXqLdadMmKwYjD3/coUDjEF2BBKatKaBQV8XDxIZED7bNExdWGp9Sf
cUe3wjxE5e1kUOunUww1vYA+vH+Zz0fP3rELf12PKMEIFmQxbdTKECYh1eDdXeb4lHK+LegQce3T
6AkhYU0JOF4iuAWns45rhIfsQx+16wcn5uSRFpyBrv1n4yyLE0Og/880T2WLB9Fcoc2hAp+ZZ+GL
A94Wh17z/XhzL3O2teqmIpWO/PLMk5tm+Wn9RLMWfuwpEIInRiNIl+aavoevaEOxtFAiDpjBq3nJ
i2vEj2apoAnVu0d0i5ULDwTAOROhhYsVjGL/4sMQDZ+KPCqtUfZqgPK5y087HsOkq2yG4l0eBwhh
50sywllNbqMvg6mRzuPBIVgJKgJwpKLFuG2AWh/occrTjIvFzYWK8w8YBMaruRRvgE3DsfmNqmgG
T9MUUeGw727RChA2sizCnhHuvxDeIF8WkpJwYL0VVhwJVCv+nxmh3PqiEpTYmYMjTjWPjFORs/zS
VgXpDBm9RKHZ9bCjpHuwDM2u/CUCZbVouXKUHimdCGUrryqyABYeJgTlugAS0GSk1Ckzmk3z3NvI
/ap7lSOwBxZxQrQR3q/HOH48wUoUNVeYjO0IFz8w4l0+jVkdcXsn92qlIP3UQlUtlX2t9DXx6hdJ
we9gzl+Ij0ytUxiHLN2rCK3EpQwgvXj9tRcgHjTDYFTIGP/UZJChTmQEZF48S6pvcM3jgyInuzG8
/sDW3ewDePS2146Vqc90h1BJJlIyJYSSRKFix100uQ4Wf8aMBXM5rc4VQ0fjH4Uf0E+GdxdxMUFQ
DZ8PP2yoAnWF6gPYval3vMIZAwo6v21qY2nzjHSgA0lcrdF+oj0bKm/bdPGXn21gu9Qaeuk/1Dyq
mBqLJS8j0f/SYJ7N836HYWYO0wda3LhG9BrvsU2qa1OLCvY0TJMxdrt7g1PNICMbF3uwmxSqVJMA
37HjZfVVPXRcxc4mFT14RLPXQRG1b9+du76mP8o/qxTXCwVqaYrT4zokidCWzhBQ39mr99YFos0N
NUlaoxmPpJL0zxQtute2drkiWLOA4H5DMSEnadERR+4b161QEGFRCq+AC4jrjXCR3+nOYXGfMB6x
108XdmRq5POe3GUlAJU5zT+/PvvL71dU26vfeYas8iJAubr4qRheyUwrsxacISMYgk5nefU4kQr6
ZjobklERcaHRPGi4cbTqrNsb9HV1nK5QnANpiBOrUQd6br2bysI3soEfc2PEoSWCLS0CWSwE8TGC
Jw3VJvHVOkhiJvxCG5IAzmOce4fpco+fZ3f8O35BC/nG9EFIYEdKIPAAMGWR6ZZ6T4qHXtDE7p/p
11Ar8WCJnfON9ppMhJqn94u8Fz+tkF1FYZPIySbYwxqsLQpWLzyxJzSreAqyjCvANDgG4pXHbk69
wZ3rMHLqqJEeHnnN/Tges7htpXvZpQqhYsfWKVHt06Dem8PSwXgMGzTDfTY9X32XvIQZmsyzLY5e
hTBVMRMRd44TjeVTJL6P1H6hMdtcgYKvcJZq5beio7EO/iDqaXuX/y1sCWdxdy/+DGfTC3pQV8Yz
U5huHj9EE3JIR8a+kmVDMF0mWYYYR59gGOH89gY0R+1GzbaBbkkSXqmONe5o8s15h32jfcjGGUub
FpHnknrt+qgK2jC28t45ccLYHjW4oRjv60EiO/g/kXOAv6ZaIncuKTKQBSYY6cOAwP1CI29V4WZD
4e+m7K/3+cJkUIELQ/hhGyyf8H2Pnynpa6d+F2qKzpr1g0cwLBMkIyruJT+fnE4eM4+21OhiXXb0
Rx69UOd+hS/TahlKhTVYc4c+rkAIGuoT/E5gJAeKSTJkQUdCfDCCRJkadnzj8QkwrmATYCk4gGGI
17dQjXyIVB7Qlfvwpx+p4VbmOLRTuOcuGDhHgn987Etc0eRkzw48H5fxbuZPXEavaKc44mEdG9DM
fZQuQU20Iu7N8zEsgEmhmeS70MM5D5p779C0wwUhUy11ZuBpPtcpEJiY9Q4OJmEVnw1shDY7nP6s
1Qx0PhkaQ3uhKfrNQh7q2ByMTn77dUOZRIGLNM38jPWIB4B3sOF1deYQQPVWwg+3wHRuL1Kp3ihM
pUzMYPzaMgexF2lqbVL3ikDlvDSNlJuHlUhQ6QDnZAVYkInw8Px9icgLh2RHKIy2vMkyQVAFJnmx
3EoLT8Pu6h80WG0xYpqT0Isi6A7I0oI6bAT6Cg2fxIn2mISEMsHzYUWW8A3ytm9TpWB2R4/FiOX6
/bhf15l0aV4FaIPH1C3XyQtLSq5Ffs8lWIRA8Xp+t8hRNy8sQOPpPo5/87dw4J4Pljoxl2MvADky
Tl83KPpUVv+vOL66to1Y6FEJj2V5+e2A2HUHLdgEjr1DS9Lp9F+rZz+53LGlsBm2fIyLVaPBl+99
z1yWUiFlYPSghA4SWNRNlQQWiemphRMWnWL3JXE9Cyj1rVoOR1HEsMlfvvgQlOgnTcLt+nx+IYxg
j1YszzRhhzLH8DprQg8ffH3WzdCL5mtl2ubPeg51Pt4lkryJjrn1qXrkfqQu5UHMztqbZqZpEhQm
USSOOeJGStp9xiZB9mRrOjlFTboM9vgko1A9VT2tphTHuGvgkNMimdsBqy7ZYXTfJspzN11BQ4bP
6Qo+lHlB7z8rt7MhY2znk72da0tntV5ltvhuunIot+tp+GOTp23Iw1CzM575iElYgK0PUS0PY2RJ
E4C6L8EsqXaLytAXwm011NAXiQQ2ISC7mglM4Lkdj27CHdDNdtHJtWypHYlc3cCISPPjZ9QWFvkI
y+IiXyb2ctvJMDRH4p1WIHCxzJpkX6CCcKFTyMqh0GZ1PEi53VqE9HKspPj+FJuTnVUdkHm/RU9S
9knCtyLulJxzUi+BugFjT+doD9UoBipgs4jur8hPftOv9jDYfKo2vq7UJWAU5c4PcPiHjUmtkMeU
GbFyfefHDrnZzl/ES/p3ti0mzL87UZM5iTsQNtj5xE6LrJIosLfbaT3bWIsYoetEa1Jih6Gonqb3
1it6CksSaIwPXwvpV4L9f/ZGUOs63hoNrUDxzZEb22Qtbp+bVRPG6ovSoDs9onRHpH1TZMuI4LQS
8aGOehc6MguQ/imDa8Bv97ihFcFpMV4Xrr+eAPbpuxZDGSdGkbylR8bEluNr+sd96D4BVOrcL/eg
2BLX2xE8eBJdnIiYY6TP6RsMtVfEXFgFh3Nbl5Ma+HnWgbiAIwNXcM3zU5CUmDOAvCXvVJMr5oCY
MfZ4Yuki5YUhwsr/QjZV9/fiaBNYVb2KpfXJl6vr6XsfMzV9NTMca6MpvgCK5WlY6HLeqUajArlO
fQ0hnKrWAJ7UP1UjrAHsxkvZAQwexU306bhqwlMFtlnzAL7R/s2Avs7GPoqk92FQ4gjDMTAepB53
lMAst0MvsVVorXG3e38mafCrNgxGhn5SLV8A+n9gxclHa5emDbrzvgRDW6+ojAmGy0LhRoR1M0OF
2hrLSCtf6Ory2Rr1HwiSIo1WlayJ65OgYrvm1mYiJ21jplGxy1Mm1C5mXOdp1jPMXj7SE4thsXZE
hHyH2LBDgLCkB405IZu+0BrKN38V40gqyxxO3sEvmm5HUuTtHCsF0549Lh7BsWOeF1drxJ0hL8vv
/10Qvrexo6kcrccmSV+oSCR0aeh15FMKIcNDEupVeFgPqll5nSAyH+Sgs54ixCkpqfg9pe09clQb
YTMQ7BfnmQ0o5x7ncDdJSFt0LzelClINFkD8mAgsCFjb2mqLTYuBIcdh0sXgoDID1XaWbqqbeG50
pv6PI9izD5Ha+YYzCrnPaWHrKK+vQeOshP5OvlmN0+8tP4SFdmGLsZe/ezfIUQbBwrDdlTaLuXX7
zJhx68phdHLtOa7ns9QDTbfRu9uaTlK0nOvfN6aauvoOE0msQ/7Hr0FlNq6QL6mOD1DPY07pcDdW
/Cu0h23y6cWPyk7M/dsvw3WZD6F0vPPpX/6FPgTbe7PWHEdvpeNYBKcqpsx1iP4rG0IWseMNR1gG
c6kPg4ynOurHt5JfHkR9BzIneaixO9mZqL08SfzLKSRznZiAtdIPK6+vXOX4nTFV0w0aoNL5i1YP
/SmkdqEQ1muadGsS/wSTEiKqcnxmVojqKTvag3ce/Vn0sI2wqAKwLcEMrpO3mgtBBK9oK7Ivmgbe
BDXBznI1VW8GZJ9mbOz426gPkTLwniQLn71wvxD3j/t9Hc0WDphQ/UndcCakmq4fFezRJUPk1DYD
Cy6LIn0R3F9ywBx2GaESnk+qtm/2rm6HtaNQ4Rq8toOc451W+vdPqtFewp/Ats9dWqezeeGCfDQm
yhCLg7CYT/4hjWootHqJ2mJzAoKOiqXkGdwVbRV6eheiivf8EKKrsQjV3iPgQl3Ew4hoqOg8LPud
XJs/xr3DnmVJxTI7jFVfA01vtlLYka9fcYt2jAVKTUXjn4OmorAbxxJxunx5t5+e2wAdDJVEThO3
A0K7aUWdkRvwIWvjG32cs5PaltiDERzqYYOg2HfEik7BXtXNxmT1B1deVaRUDsmr+Jc/yPIAFXRl
2RfUvl6aQo4Wwe9v/mcAtDnxIG9w0xAYEMzgTJPabWJLqLoQWdt5h0JrJ7eWi/GLH8KHF7vydiev
w0e3MW0d4YLj5BbloTITYl3KBS/xx256cqPGnuQZx2VnxYB2AjVdHC5J50+erXjKskKQOy3wYC/T
4dIq3QLw0MfLoMJijUlo2oDz/DmF1yU0lyfCzuGwQ0wiPF8N7W5rWr9MEWCuhmvTOQZkP0OwpPLy
7zQAS4GVxr7AYAVE+YG6LeZK91x/Kfa5xEArjM1TAgGLqU6uyeN1ThJ4FMNOfPTCwZBq5xOSy+YL
se8j0Dti7wnsZgWM/sxyHLXBupOIdsotwIFWTfKRrBXij2Qwf/w9X2WCOco8hkXoegWomM2TNG+C
eJ6TdT8T4gA3PkOYvmJ294IhgF0geWsZxrvHZoQjy4N/7ksXlL9UmkT9RdxgsTtFBIpLW53pL8wX
u/FwZONl2IXAcQZ+mym9N9tj2I1KB3JLKejbQ5wDChoRcJKXeXieS/KQ1/Iss4XbKZZLn3S5JNVr
a23zA/ApoMsEK0LsyhWuijy48E/0ZeINJjd0LZUDR62ADTm/zxg0vXIoV4dB/F9o2O5AtiIh2fEr
tKdZ1f9Z527l6LIFp2N9P0VR97qkoqWxWi3Zl9FixXaohP3JW6ztXdsbLI2mAdro9W5cdaPS+rvh
7VVf2hFVBRJw94ZLYTo9XT2k3LjtzzNZzo9HD2mMZbGxdpuS8Wkos6lWw0MtjAFkuSEiSXyAxQMP
6rqHe5Na/9FeFyU/JF2/ENAwSHxyW9kqY1DxXsjREIn422MbIXWMBnOj/sPtB3a7larZjisJxxmR
ILFQUE0pcMr0TtCFmxXM9cRegoBqOTMdzrdnPKtnL1qw5THL7QVINePgEOZhCWRz4mYQFP5W7Mnq
b0XImH+yRP1j2EnCdSB1+QR9G2LVBLgcjBuB659xPXzVI3fNx3FLpLqrFXJ73h0nkOiTq+8Vsli4
Kqh/oVJZiolOVB79A6wf5yIdbsgzd04hvfQmL5NFtaTE2Z4wlYFuwHVUs5H1Sq+MzPITmaMkpali
2NjuKDQV/DJwbddneUInoQ9+muqkpdjZeJ/8tlnGKhp5ZttIqfxiu3EQ4uDcTsGvdrUx6bs/NT1l
YTlb52ftOw5xMIGqs7zg/yKi99X22KOtikySnUPR4lfrgqTEnz3iGixfx7hEd3R5tc1vGRVBBWOS
ignewrmhn8JWRAmrWQn/Yvo5SeRAJ0f2WGv2a2Qzv/gLjOuVqGoVXdcHv2a7aFVWcmhN6lLAU4vS
m1TCLKOyvJ5SYAOkfKVrvkGK1zgWQpQUj8jjwc1Qc9TRzItEt2JG0o5/zi6OI7t9aEWE9MvogrZp
xPCJCzfIcxqMygb2ncJsg0UYPGVDAS3YJs1dVcoq/wKm8xOHyB4vgJq6P/EXDgygf5esOjNTBxCL
6hzRoXpA0NBW0Jf7YNc84FGC9SCuKRj3+oEvLCPODshqtHgsVwq7w2otOPoh6gfY1UaMYHDYd3R/
sZKJ4QOMOBaD6b9mn6bBpbKmSVcP67JQweQ7w7JU67yuSgyRqxs5a0CNxQ2x0J/eVkTyeNy3xJfm
UsebInrw4ebDWsgvQOJ3fyeKFBkc/i13cRLDKYgtmunR9ZJeZVtNHG0occ+44eYVvjjEqvcojiwk
4/OWV2e2vscD3AGmNPgK20N+gt7JlyLY5bz9F/vzo2FeW9B/vLCSifhOMYX/FYGg0kicDOkaHxjT
pSyqhIB9zMvWGJwT4U0aatxm2Esqz7rQoie/Fe9a6Ys6wxo33HD1iJcYdlwMPMPWn5cVw4ZZKk8h
5G484eIarKr1mhOrDbKDRGd1lRUNxNmXw38p64R84moEpwONAymh6mBSuxE2/jRvKr1SdCLJp28+
LIngMvNSLZQIxDfV0xXxeQeDv8yci3T0quEB588vEBBOux6uXCT9aGv1VKWMlrRN+/Coy55cIgjN
K5SsBZ/tAy0GEBht08U6AoGN3DwKclUu9msn9AN9w0CXtzi5B71+PwZGrFP2M504peNZUgf2ZG2s
GcAPGLwcv1Hh0gXVpZVTtZQjj0lXU0Bzk2AsYaYRg2ymj+z0+awZXb87PAyOfxkVfwLPvkbrYe9X
zxau8G2thv2rEPx9jPfMYe+TxnYfkDoasQuMQHD0dOlPY5CG9ujJHSJIUgF34AFEPtKc4mROxch4
A+83EwqU+7LKa5mNGHJFrLJFxQUx4F7uCEwh8D3zQM0x+rG+/tj6kHLThd3gBmneAaBeyJu7B7Ze
CD5JyoQKcu+nV/UBnRkjAlajOq+KkrNHp6XM7x7J0UUYlOC1eMteA6JPTkw+hRlzXLzaGw+OQ5Jm
5Rq2r88BgSOdfsPCb0kZat1Jdt+o2XnT9+q5WjsOsHW7qJiiQob3LpsfXzMoxGp2ZV7n07o16PZc
fint2OkHxXp6vBod30BorHuiviBOHGQqZKM+1wfKQdxWfIle0EO/vIT7g5dj5illR+c2boFQFdr7
5Ew1dfTxWMrO0KKvEbWSMg8eVRIlN6KwIrCto94IS93eZZGwRCi9spAMz42TEuwH344SQZAwzPy1
qIBSAIOr8+6TnMchRS8VTAggUJOz7tJbKzJkFz5cGMu7A9gzbPWXGS2leudNgkJmjYK/wQ62Gz3z
jUWCjidSvKzRI1uAe2jDkNBgE5GL5Bwqot5efUlgDZtNeNXZyfdeQkTaYStCq/rDIkN+7/eqm3fG
HHl2ubHj8zFh5n4ACGZhXP99RhdPmX2MJsqZZsegwap5XMr5xzfWyA6CkeaPYGrCG04bQpLFkrkw
qfF4tFXRPWxuaF/FWrK01N9NZktvPGPj46ZfXM0rPT/eylRi6KU2lzSncbacNudHiRhkZQi/yx+3
wQGbOYsBOgIiGJcEsVGR0Kv3lzTOwKj/kJYJARnjmg0nyCCmF5FYrV24nF/25qQ4SnzpVoTGl5cI
Y1KBuM1GKYdd3lkHXIS6DIdaiu+ckWXTpzYfmllFbRo+cf8BWSNMmJ8/qW6xYAgvWgILwXmdusST
Xj8QFAqQjP6OeQiuI7/qNcD0OD3Vu66cwD7UZDG+p1agi66HV+5iarWCJTex4mSxQfXCZHTiy7Ei
YotEuTe9O1kOadFSpxLC6mqIfvvvrsLbxioDOctOh4lDIY95dp2kBpbXbmANPPbng6ndTJfIEs4E
vnjbk5DzKcjV9vVixXVLHEAzIzfprA9JLyzDuAuqxhgt1hSPTZurlwc4Yo2+hzKu2icXTWP/AUk/
C+uWyjbdCsSNTGmo0OHrYno/SR5O7AjW7HrS9a5QkhcFM7e+vIeyLfXwtMN5MZ92YhRAL4bR69Pg
iukehZrCM1G79aUdRN4vYPJkRP63RVY2UEcHgTdhrqzDOHKGY3Omr4bIGT5kdIFqB9pm97IuSyPy
zZLfWCuDDMxC9ShoGyOyaZCYnjfm1zLqvqjehUkGnirCh9p1LmZ8kpFJPfL/rzeAOMEbHsCFqqub
nCeoxK2JHFbCiysEpJGdzD5UMnhWBJiSox3Wjv9U2Z+nuJ8jW+VIeeV4r89n/padCM2U6h5zGKou
CxQKpkk6Gb46Bx0NWBt9BRVZxCMDcgtJoaxjAzEFKl7kDRpNidFvuZq79bh+z5hr5vo/9mhaWd23
PMFCqnUwVhSrBOMbqrnF3uzyyjGKvLBvL/pntvlGTe6I3AafkJwMeDwvV7V/ivqPdvBCVvAcNDU6
85DKrt1pG/FAPUNb/W9mYOY9UmSuv+2aciNiakhA6wwIDWzaHNwCgwF0zbUBlERh0krNmROuN9P8
te/4OBSoNVfNjTGc+27I2JuE55SpezQcAU7KTgMw/+V2hbokVjMXeIOmFaNcB4byIyD2aUePrUku
rc1cxmU8y0d1a81L/bKmUOuMDxoSSO1RI7sIaYTCB2vU9k7r115Md93jdmqLGyODkTP00dMb6YgR
kblHNRDlLqFPRImn4B4rkHRWt+ku0bOEg4Bvr4DANeNxYDhq63j00f/gDbPWSyuiLKZbTG/nNz35
gcJM1W4lT/bqJ688ah1QIj/+zobQHDfETYpF4YyWRlmZpqhmKsfOG3fxk2MURO1JXDLBV8yXBO5k
8vFsMr8OgrbEV1DAAorb+7JHrw9O2laopRMuCCRDU3iz1SNvxtInPcai6VsibTlTYHSCyUGhvgg+
7180ydcNSga/MZbryChgVnaWuhQyslaCqoQWS+OOgcp8TmQ34imMxY1xpeWS3AYjmGVO6R9neyIF
3xpnzA0Fp2XFaIt0XpTf3KqGrrqs4Z6uHu8y1xxiHrkttD43BHz40S4arvDSIaXMC+Blh9RaCm7R
fkcYVnXqwfq+9KiMVWpns1pTwHCe0VDetf91ms6CeyemdX6JGxQaJmsJYBECRikW3fmOtPBviBT0
RgHEISdMTorDXl6XnBFBPTcbF/j2pXtUWwzzS+3iD+7mdwfiXTnmWCaCHouuBNO+ECe211R3L5Xe
efWNLtm3y9NI+pASvJK/T0P3ygvyjynic5dJobyyDKzkq3BkAV03oCp6otVQS216atIBojWnEKDi
eG0nwXlgxfr0D4L1P0bmQSis9Wswj1D8Eqa+dnNIJcQ34CcPcZnAjYww4JQgK1N0ZbMu3Dhf2sV2
dMrdpNsXUBOq5RVTYMCzo/yOwMvxe9ycdlmgVyYYZl9zsZWaUBxPgsi60/2LfVCXBw0mJj3vKAqh
CwNaObS7BCNSyxGD27X1LJPzzEd7UtQmCdwyQ3dvmVDHroUakAweqYUCGd+TrGY9G+e9byxRk7/Y
B54w+i1gMRD3LdbAkEbiUFAq8ORj3v5hirM+xkbG041t0fVQCxIqWigBvKF9aIA+8q03ODSm8h5I
rCwvWFv9LD40qcSrcTpCT6QKBjdLE6BFSUn9vsvskhK1Nsb6UEoeY9TxRRbQHda29my5tTo8Y0Et
HPghuXVPyRlzDSGvqM77NTyDF77AcL6JphC35VwfMEcI7P6Bz+KYqw6YHwHt5Ahf3MJh+gINOmlP
dqYRxhGoBxr/FIx2DUYa1gc+3iYIwrkvlY962Otz/jcZqUxZ1BFY0Kr+7Uz12bvDiCsm0oMsHl+V
tjctTggoDrliqL0T+kz451bPbatKX17y4zMHVJRVIAC3ozAmEK2QGtSNZQFbIdun57yAWA4B+gaq
NiNvyn9ZBE/xdI4tLmjCXKRt5ziF/a56vK182ltyDeZuh1eNlq08V7/GCSIUfa2oJB7iVf2Baai6
rEHjawQ//uBcnCjyk5QP814yEpB2T/1pPS/Ss11H+v8RtJBqKBgy+JZ+AnvkgJUVql7v+mOHGiqJ
98GHo7/z4GzwotZYIhAj8YSF6O1TGRGMo5Jr5JB6tr04tjTtkhtUP+QvfFl1iqz8JUQeGRIAtiWK
+bpW24Z2WOhkP6EtqAwLxi/Glf9S0Is60DLzS5XV1md1uKerUCtJFjxFDzw8grRgfhs25qFvkwQF
KaVuwHyaL8L3B9wwDSGyw4lTtajYFWpovEWzFihoq+mlozu0vBO8DDef2BW66gr9wHmw0ENR3yQY
q4otSV3ssSrBDnIGVmSYk5mx4muS5jkImD1BPBghVNtawiJhXq+F3+HgbtL+AnaFm8b69T22P0y8
b1Epw5uLppI8y+rdjUU6W2FAaQTmVsp7HixKZwJBK59EHxGGNGwK5crV/2+dMWyg/cfc2KISQXkr
f8oHCRe/rmMQDB81k+5ItCn6q47teTGfBG4nlTveaVqE9XWrTIIih/VEK5MQLiCsKQzUZxIAtfMF
CZu2sxhN88sDzeE85OUDEtSFha4v2UfS+PCIp5YMYZXaZELLynt95HsOJJhKflIZEUhStvqvhdcM
Ruoby+HgpG/kNtPcB8vTJk1RsKFZKj0PtrIh/6UBGUg4nnH1+adqPKfwe9qv1q90Ha9zumxLnHcm
j9cVwqMscZwkCVVjuzibNfaRTykPPn/2GaT4lLi0K9PxbH57mwtjNLp+Ogc1/TAzJIr/bmMyqfM8
zKYuyk9N8DzoW2gBpTYkJ3KX3oDFbiynRd5aZ4i4VA9ElQ54yNT11SG+BKQAG8t/Fnm48Xa12Cuk
85C29m8j85Gg0y5G7Im8WqiyLdXJlmUHmSGSApxMAAJK17yRsB4NVx7xULZOlPcZSqRhdeJIv1YR
M7qGK+9OuahI0DCDu7i3pai4od/VDXA8U8CJsL6t/l0xxBNdZe9eAQKb8r+mzln0STu2ukXvDgIF
UVrqx69fcG7cxQUhv+56HN+80m8VSlQnL9NuT3SUzhK555fzwW0VCvCf7BDkzoBZFHsC4xLFG9tX
Ty75EUktPI8fbpGeK1GaZOUOjQjdvzxK+HKqasAaUXi6R7a8uFVlUrbeteKHfhGwT2nRJwLS0iFg
p7LTWYlxr2lX9DyB7HCfepR5J9phUhrpUZvyKnNTCEgJErUyN2NQ7HNQMV9N1uKFe7uaqTsnxyLK
/lNKhSoL06dUEFz6YsY0WWbcdKr9v2m/DAlRZB6yDE6f64C5K+tQrFvYWb+LbKN26/IkUYmbc/ti
hM81CAqX/d3PTn3mDqXh45IUGMIY2LnBIok+vgAMYjU886UjajsyJPBq1J8GuPX9iQ/q/U94SnUA
ZTkZqWNbmN8A2UtnSDpC831YuzR1CWGL+b8Rbgf8TFLrUG2KHBQBSnUB0sjXtkBzB63ajk6wivW6
vgx6Iz10P1ySyoVwGAvyCHmCXL59U2foG4FoxPiwIzoHw4MeKslkgbIx27Jv2LdhcnJwEvvAsRrV
nPlb+6mCe7FrC6sOR6HoC8rHjwF4AVmw6bUa/O6T+U+5GE5z5IiHPrwBVI3x/al/FVS54XvbED3O
aFTlPJJMB5SllNE6EJVAOwwYXL3UkjsW+jo5tJjU2fdV7ZMcPSZd/uf3MGTUb1M4We8flw5X9tlG
/h60TdRvGucjHfzx9JubuY5J8P0AsSHCdOgUBBpsdPmAtXj9DigEENs4JkQU/QRT4yGKtSWxzhBR
veuIRpHKdMOY1oba0TUFkphBknAIi3bCEP5x/Hj9kVyeWg2q9hIEKKMHuDIGMOOXBBNHcwDoIaW+
VWcNA08mBETKrEePEMmhriPvrm9AZ+vBrC/rg6gQZr3IeFHRdoUHJo3DVGEIUOj/uUZMFzJ/oxSO
SsmSLH5KxLuDogObWMKsRl3lDovSnYQ2nArdGhEt4oZCJHzZCkkw+V6+yE38YbjXEcAMP/+ZJZnW
rFlCD1SCUe9YiUX+XOC4MB9lsxAXOQ2ks5n7GHx5sC4qJxwy9fqDhxZMzQTexcKebl0pijwKex1u
pOSre5/1Tg+5Cij/MBfxW//gD1Wu5lT5SjXcEoGx+ulRfXvrt8OLmSbEoUpYMVVw0e9XiOoQKQrR
odk5KDbx06Qa924Cm1fAUWf1XfsXIDqyRLD/cMxdRwvN/N7mDa+zTtpktXENaKxtyAi6xwipAwzX
dOt/50w/frYGyzeXgJRXWTpOdygFyia1EGRYbHB9+OgK9E6wflRZ7PyAC6FyAR1W6rcD5f6H8p1g
lOlDXMZZBFE7kuGaHD0YPxSwjiqir4ZDKlQNKnd1cov0dg1Z6uX1FLA/UCPqiZZbgHfknWuR6tFQ
OPdA2nMroInRCNwtd3hpafr2yOxTGI6StiUWHxUfkQpwqfr1TUX2bD5VwNFi8/D6OtXqT7rV8kFr
fIFskWgharebLP4QiTt7+QsjOH1e+VKp08j/YCDxaTcIrCWsxf25HumVrTJGMrwS77X80DyfyXyV
Use2PyEohQQA7N2FoVAe+o/OdzZbSESZeV5OgUzbVYnLYQIgoV2vDSCrScfRI3Wl6hIIfZtgRQX3
Sj//feSBYMgcw5kqKKlIDPOFNec3wUdqlF+zDLxO1v/9MbZTN7fDx/7P92/4mmwNoFL6AHohtKP5
yKHDrRZOjI3PSXRqzBWHfZ9g8RQEsDDKrrj+bGDwMXatSybn0Z+aGGvQcet+yH/85y8ie0kccJVB
wiDiZ3PVOH3U9e10y3VWJtaCIvXcANV+/XGapeb3jERz1bXdal0O50VvufXdcsZvYxUlEOmHFDbD
JpHP0GfMoqdU0E/a0NFpGkTiNgOwlOiQyzox6QitGwPGchcCRYSHxCFBZQ8H09MmPbAqt9sdaBqt
vVFR0V6NANhy0X7ri+CF5djcvZg1SRKJ6OgL4i8Fp9ZOFOmOuS5upjDSNf4YnwG5de5bJjU5aYO8
SoI4BpmjSRMfLWyXAKGm23Cz7MyeikChjmiP/I3tTFPuG9gS0G5ddG97reShko0gsywcpVnJUVsj
rMwfkVDhInXHNMf/bsSxUuDDtC+C198xYNZ/oGjPWg9s8n/rDHomubJ6W6McXT20mqhbe1BDWF3f
Oc0dnZAL6dEYh8vlzWA0lhDROBWXHqo7esCnwCQZq+TJm3s0mdYxpPQOEXdGuQmngWkmw6OLadpQ
+TRweShJc4Avj9gdvYdzU1U7koT/KyTdmsK3Dhop08Arztlgi9e71Sy8bi+0Ugx4tniHgPpbhUHt
/pQ9LWWigr5+yaX42E1WOF+TsN7VuAOK+73ANqk/WOA9+rbu18GOxV5a2pL8xnJnqlwvRVNYv6V2
R97BYixsqEkvenSN6nroY7nlStnGqH+8r6Rg0qQU8dJ2+Qynhzcfu5Zcy1+o7E8GO80BfBrvOOMM
OODIqr4j+ihmIzoNLhDBXysKS97/BYdTbDHfMNpFX5ZuBwcILbsZpxHdgPtZTzo82lr40teng6Oi
h3XGGcR3J0T4jXEpLFy7eiIIcqAIc5iOHOYQICiSjMZI0kimLXDvVAv0oo34AlFsZNsGjulxlMdY
ewc8r9ZGrZusE7aWXXlf0XxOnrvp+PICshP1rqv+CgxaPApriV53VGIuEOG8ClF0Kjp3vH83BJjE
1CskwIHk557fYIVbTHbEBEs0QiGnEkchuQkJykQ7s1QcaXjH8lt4+VUk3cB1v4OIXvzeEUNW8o1/
dGFmf8bOC/FJ2+63ul4zmaRj0lMBIbh461ZJB6dXbkZmGp7ip5Rjtb7fcHa4PVnekFt24MdL0EZX
gr+B9o3Dp5ehtuQIvNiU0NgLMZwUx6ywbU6sbfpmr05bXIWo4MfhmJ+T9GhSJ4CIgN1cATzRNT64
oYlMTt7o+FyJ0PkW735IKZZjygYfsNJW3FSwlbMej8/zIh8uctq9vLb40yIYn7YTZfPOBj7jkAlD
z2wiWrsu3pDqW6gdALBcApocKeAWur1mkni/xvcZc0d1+Or41h0HeVatpC7vVjPNmE1UH2Rrxq05
oMTZTNxVzMka7dOrKOsASRAX6lL00ARrkuxrhZuWz5D8meAhCL22Xk77YCOrtp454iMY8gO/cYlU
XNYvlPxLfTQBlbh+W+8FuOQ8RVI7Dnq0vAArULnZNUvzybwYdszWFTFv7rPWo9d6YaWMunbWfO95
bKGCC42GDrQjTK2VZycrlTBmbx01l+tQ66oHbvZcUb3osL3TPxg8kxxixVFxTHexgkSq0CM73eNy
T0/xVMAc5DWCLjo+WzazMh79RCGOwsKaClI3Ai8rdvXZWxKYzzuBjIElf1apD/sPbJvP7eHD5F/6
FM25ndEp0rmuIUe7DsUK9ZQrtl7C5JKvQokvGnaDoXew5cj1NDJ+XSXT/kABr0bYcbNXyPJ7Bgjz
FGb9EqHFWq7iGi7eIVLCZeFUkvLUIRj+6i/enbGrT87NHKOIAsO2jv+0b6GIYBBH1Ij82clZU7aW
bJSTMbjYSyswP/2CexwqYByQOpMbRSKCwvkZXjM1HO5nLqby8e2GmQ1A1fDzpjLve0N8UY6V83yd
+cMJ811HyN5TDhmB6sVIK8vK5YeBElyJWAhrCaDOOKrX9Vg/ekz4OBjSKbsC9BOQKg3vxd1zOO6D
LvkINFhOVnsLpZvLsmmeUn27eA5HooOHmhMJVWnf3xwm29ZNJt3mKjf9sr8PKMUDORrHbxgttP3l
HuvCDynUAy3fb4AoQGrSsTXBVwdDe7C17RcXrD+F8Xf2gOpTh5/EPvV1ABIq6BTXzKRbVcQepm7I
C5Ko2uAPiasbSCeE0frGorsH8kjhAilgDNTbgF7leqcLTT5ZKTuRqwB7l+HAPz5u3+WbC6zN++dj
Jrf/Baa/6YIdpAHiLQcyRv2QawsBzPI+zUu+m3YeivMMQGSuJ0CoQ+cUCV/j/LS0zRHOqJzqYlyy
yyOtJhgfNLU4f6udzamP8TYXuu++Sdm688ldYgmMkSCUVYnq2LU7B1/9NKeIzKGY9pOCTQ6ueUCu
SLCjU98cFsqL6taiJQPgYw4lZxooy+S4edjO24H2Ly81o8t1R92eRq4yiT9uK6OgHBWAHRInlqiZ
sBweOiZtUJqsouMpyZE+k0WeY/yq9lk1s3JM3XZKTYj0k0tXVNZv2ogP8W36UorDsTVE/Yz2wqrj
Cys7v+2nwRUUX4jsURR+mM6XUXD65uLm5XzWe6UHYfuNDa+nj1G+UZpZOHMEDemBigkuL/s6cWc5
zowS80l6RwT9crq2T3SbAm8kAq/f7myCp6RoG9wchOJyLe06l5YtKOY1TqLQ2yLvLqy8nwBirD4Q
aAFzse3mqcst2FKEgm/toaXDy8HeENn0s2UPAOhItDmab6QKmb/C6coR+i0kJPcte8MJAtOiau8k
R29YmH1fKVvmYiC6LPZMdhEV1JUhmFGKaGK7MCfPl4mpJL2XSCgdJLgpNRLxwkAn9S566ixl2HdT
s0gcDYZImNvT3d/OrysUXRm3nEKaTrx7blscqnKWdRypl6/u59+uKMOTpum149+/65zJufPtArId
DfpORoPBvM9/2Rgeoo7Kb0zZP/VvhpMcIVmn68v4YRkPc6pNDIYM0HKoTimB4+bT88CJP/nyXG2d
t4Wo76/mY+FmL/h4VVkEpROvjK4furS6BW1dd1T2XbLb23+c/5bnWdhG3/z+ug43muSnQ4FhCc5F
5+AXF28eCdSf8wOZ9iER6lqI2z1gCwRJWuxzAnY9BLU6r5le/RdhuSQGlq6YUSAf7TFpwxCwQ/w5
fWk9z2R7mHaGn3K6ZkKBbSejTwAMRNvR5RwKewG6gGye3aVJ98XY2xc4WX3tTKVvnOziOj/xL4Zi
OjXWEOnbiT+8vxiCtVNDUlwvVynqsBmBiYay0wxYlPWyLG33iwY/1PYdl0ILgZ5wKxvWJFM/2Pr+
nDnMdiyAE5x3/C6B8JPt3cOwhxfQeCoWm7C3N8Yfgbi29Md8S92kz72nacV/loEBaiP04narsnjf
msOZybYow/8Vn1IX33qo+KRPLbEIIWHCETIQo/QNlFeSpUSiUTrgAbI6JzGa0rtbUC0yv24i4MqM
4aQCByYlB4PWmSeb18RT/jeJE9eebZwDucsTvQgVKPTQF9LYOMcbumCDr7CiESaUcPd1kSZMNNpQ
giCM3oykWVFY4CaGsfzU/OjEn8iEspBm7FXaR2yRUr2mirwaD7isRuHPFsCwA59rDkydbo+G7jAW
Mu/1UGvE1Out6AoySrF7jEAfKD6h96zbZzzwazsTaAV2g0CJ1sJF5hzMEpgizXAv5Yzi2oDyL2GS
4TozDbGh1fXvLK2xhAyZFf5jYh1+E8PGzsrAWkAOZ9T6/YLc8xt9POsORxBkj6/gUgDYld/RhMCw
Qp76a3bfWuUTk+fWROXsTdg+oKKTQugc6kjz8Ft5+Uo278VbLGeft+htYdJTSZyQuSuDK7cILHTJ
yV+iMENtq1LEcxe6UDfSZsGcXD9durW/srJIHY0ug0LK9vc04RjkvbYylgHuPv/wMm2SmOSKHgXt
ywK4FrUorTJcKsMrNspW5KoZ/LEIw8RUqgDgSlOERfdSlgxtYl5YXfLKvno5noaKrlkZuF7uXqc8
06IepallOg/WBYN0tRhB//0ytkffCg0MYYfHyH70/VDJl+ykhJb4Mic+TYhh+cdZqBZq9/n7g7ZN
0hhOK2wCdSd5tDI0PG4PNxCaoa3Lmo+vRoBiAs6O9sGPcAXUSgshocZAyNlgtcFQQrBnTV8Cp/Su
CkR1+AQRPOpex0JsT7GnqMbCowBjSxRDboyON8R/yNDZeKU3pXATYbD79ncM8hJ8x0AQ+DsmsfXn
Dq/hRcZglY2cH8/DEN1pUHczRTia/2uw1p1UFz009iq6qt59I2KKp9Cmo/I/A1H99AUwsutZh1rh
QNrrGN1TXqdqoaEw/2yNEe+Yt5TSx4GK3xNtVFq9X9dk2G1aSVFvbu+xOGbIutSMwFZhJRc/zyTf
GAUUBRfky7IsayYvVDPjf/CRdcOUXVBg8rPQaKlJNL9Vth4J0oAeZ2gs+ATMruI6RNy6bLjPM5uU
6dVbfLRT/sUFPvNpuaLF56DTLwwBu/tz2BFfbqd8DHXbHcPzaGxAKPOz4U9iidR+1NF2O+a44+0n
ygSxaDCX/N5P/X3aSMoS4pK9Qy6VmSBNjhKT2daTDn6ytfEYiLae+yAMHOn6sWH4ntY3/JV2SEdX
BGXS8VcC5Q29viujTdqtc94DbgITrz3feYRFuTzTQ8t2+8oODP9vpM0Ce9QEPjmMo2ZBxbAhiyZZ
Gdqkqa97E5CsJ7FEIwyw6LHxt2KA7emgGa1SsjhVYtbgAwNhXCDxbm0rkw3FumEphsejkSKpIAQP
W66+MCYbXsn1ZUOwqaq7A12KjC3slNCly5yILlvwHA17sRsgswuPq1daSROE8lrIt3r1D19Jov1J
Wa/p+DIbFCpXxkG+IToePQ0XkTyVDDl0MfMNTb+OTrDpn5ywSicl4NqiollS+3fxEgPd1fOmAApf
9Yf86lZ1nA0zN2tIQz13mcTe/8xFpLgcd6oqfy0PfsA6wlUfrpLfd09FGuvfW72L81mBMlYBopGD
2Rn4WZIDQyQEVTI9UnmcOEdTXN+00NCE2puZ57pToV7Ss6kfokCjRI9XMkz+VHPh7wttdsSmmGLX
agJLjJ5mRxSRR7VGLCKjUIqVNXzKejor8c6TN7vjrRAhnR/V0o2EPfXHJX3/kLmGGeWexJ3hB/WS
wgB1VMBQ4dRnrQp+pSzoaOOKPhXVt6hDUBbH7eInamLUUy4XS0D8AwPLfBxjdxO5pzBb+443SYq2
oZYXWC8Qk0AZdhXKu4kb69gkM8efnZ1TQADtmaV5RAWXiTeHGtjlhBtDzUUz17aurGb/2HP5CPYD
wtafy2NOifCBhKZIa2imStEta1FpGx7wgstUxf7NRn2tuF/DhmOvqOveAoCu4xYGqpghnwDc3TVI
N15aaVqi8HQMMNkLv+AOC5T/7hjY6UJVwOUL72YkWD3F/TB/74KSU3/MFXlMqVUs45u0WbsCR/tE
kbZDLgDhBBOyyZfQjbCZUaBw6u4Cbo6TWog3T7W3+2/mynzVudEzj+Mnxv8pIT2wdkYRlUrO4x3b
YX0FmDdNCdno3ZQnRCg33rVy5nAhKdB/N0+T0X5WWghMZ7cC9UmqdseYyoDgskMFFEwODB1evqLm
PcxNQx0aYxRo/zxGNtfT228g3HW0Hvb0Y270ib+tVItxwAfZcrbUUJvkZNClQQCD+JyjjTndYRKm
es0Mn4YrVjuzmJ73AxHtcRl5moH5KUQ1A3BZmjY02JeGMq+f4AQN3IqG7x6cZPAu6IGKOHjWWjCL
LXwQRa+E1CezgBzUF/Kd3QZB+nLoLoFr91HHsTphs3r3DEQd+oVjzgE6gBVc/I+mBdl3Q6xGMaYk
7P4Y61YVU0MRx8HQBtSf4PhNmd7yN28goyHJzJUkSKH+DkukiGs/7fnBl870f6Baohz72oR/qMV0
rCi0gFkkD8SMbKvO78E3H2kEodq8gxKddf3xJWPGzXgrQxBnFX3Rgy6bg+VbPeAonoDxSnUYX2pe
WR9fRIiPikkxPEJsEI9FKj40qwLiLUhDghwVObkZNDMMm6wZG4g+LAWQzckUIRl9j14SMPvIjezN
hpDKTf7AxOJZPGSt/VXot5V5geenLYtPHYhOYyz1vYJ6ns9mcnIT4o5OzCxS/dSuv2sJ7X4jjKz8
AkMKJXRbYwOvmxBfXP/MSAozE+ChSi9txwBBJCq949ukCSSYcpQxkIkbXeFDZk18dloDFxssRY2n
FZonIyfJuuz5yN8t4WhvwmghSbNaEXQ/lfvLLjE2TYF9pFxLXVWf0GZFNtCclbF2arUeCUwP9lgF
IwEbkEPR+3x6kkZk7A49J3upDZN2Lim7BhXOeqiROgRQBSsIXbCSicZWSQKSmPo5eAw4CylcfTtH
e1yMAMhtKqNwlz3WjoX/L4Itz3ne3/BStyLpyQpzn9leUpPJcXO7AiBf3g0wXJ7TqpCVmUJez94/
S6FD5pOW41oMQbsLAWfQ0T7DwlAAg2jO0fnfVExSh9sZndv8+GKAXAdcVWy+iuHxsLQs/bKO1Lz0
a34H8cmwYiL7zLT8rEmP8F1UAL6O9YnkzE7TwBisqcmdbSVRBNNJ7kqO2m+jXYY/eJdSuZjpzWLT
qg1vnUtL2isrOSpH1/w6mgCbTiz7+kQnu6l8OoymQMW2ZOt/pWnQ4GyN/2Bvhc6UC9YqvQw7UkO2
0d7f1PhtP3QZ3qzqYlZQeRXObvIzHEIJvtxjuSFXmx3Adl/u0uMtFWh0Ay2jPFLjVLvn/grzMSou
8HW7+Q5dMdooS9LE2bByqY184Ukgntakl8VBLcaZ+PRcVN0ixgwnSMAWxpE3I+bta+Pmv7og/sq7
T6d1qcJysem6av4nG7DjOHtJtGc89BLEZ13b2VUX4OWcWALxt5CrIH/H7S1VItKhG6oCcbzf0oDU
Gz29PLVMvfN0HdFAoHSLRGa3glHVMnhjRD4p0nMzAWcnyAB7h88eDGJlNtzdzdD39/J4xSEHafgH
yQ9zKdYd0JVlcF60xn77KXjaSmaJpisYM/UfuQB/8wQBjJEScjMK8RgRm7h8TEQOnGSliTBWa3kL
9LsQfWDc8XJXeMDKOmNFYcYlOcrLMClEaVdpSjOTZNm9cLlm8mlabrw4bFdumvkG8XqfZ53N3+3M
hE9KLmGLrDCil1UAkUJ5n9sa0K1WO/Y1f1Ue180J24WNDtkDH7x3R2GD/HpMDvELIMFP5Czdz3Lo
MM2NPY7shCK2HuVek/PaVo+BOwv8YEhhVfML/1pj4SpeI3V2cJFM2+3zXYQSst8nKgFoq/L7cq/R
67nIe8Pgdt40WMyB0biUqki8ZHbdIS0mLi6g9QiEC+Q6l+A6Gn9rX7gn0LRmKH1eNvFoSh0XNWGd
8Uu6raWE3nQH/kFP1+ZhD486tx6FBuP82knn5D6a/o6xr01FLJTShx+SQj4igmrnM00XV+taAaHQ
RvhGPsegu4LWvR9ErHBDwleU7DRMlnV5FmkpKnae6UhT2PdfZ0EcsyMSJMijS5u6dqjKZyZ0t+9u
IEbn9OjZwM2VMeXZ/a3DHkrjDJw6/xLCqFQJuXbhjXjWUxddOgAJSqxNJKlIvknX3oAFlQvoRoWJ
ug/zXMNQhubzmLp6FJOWa0Leos4bvc9PxeU22UkO0ySdcHpniL7kC4F7Bc21Zlpw7gUg7qWQ/63r
EICT0ox4NQ+lN0XaIM/i6pqhbbHw1yAGXHsEG+RybCOu6AEIuHsKsIh4h9xN3jH+qViFvMEC7CHZ
0g/PFEaw+ea79LmYYTsAMXFuHofsm1HmyLBOGiVNgLCUnEgkBytsdrcvmV5vmBML/cY6NxC8yp3i
hyiBk0RmIJ7OcSDd+8+6tDX+YkKVeBTNtjcHBAYAduXN1IGsdj/7LlFZYY6Pb4iSmgK5326goxfR
7NRryCaYuMTy+v2CMdE+daXHn876H1r2K8CXhSroFGF8UPmvv9gE3um6CMyP9vPpP5qdM2PSfFZj
uv0LuLHMirzdTaLtieV+c3dN0r92dymfSYKuQMO4XL0oNehy0GB4M4Vt8Lameraa/XfflMYBX0js
qMBNo1+xC2nRScpQ6Y14DW6Fh9xAeT12nE1PIjcJpUvDdee+J4VO9l122Z/o4+iR3jlvBAJTHgIG
tzRZctyuLGJeBLoRpJHdHYYovOXk80BM3mSqclCsO+/CECg6/GXTCh6S5SL9hk39tQUc6DYxQZMF
X+tvvlhTaImAZ3uzoF8AfBI2AibenW9AYqUGp4g2///rj1oq071GphkFQ7jt3bJk/i+vWqgCjmh7
bTqhLABqv5qh9Oab4LBEtGFNECl3Z4CBkRqQ0/0YkRfBymuy2I4T1/Z7590nHodrTN0SNz/zW0XU
9mm/xZEBUS5mFpztLMr6nVBkFUmYhQc0jXS1uHcKlvo8mebOXPFlSJWAoA6Lpi54wp6AtwYKiROO
80rnT5cx51ruMbKLCZzKnbzEuFMlLAOfgkE9M3P7MJcjt3zx1JEsXwZj5JmH+Y0vwDlJSkukbFL+
JMDYQ7BHjoMWZf8pI8Eht2eov0nd/ULxZIpTE1nZtqqYGGDSiuQWNvKj11rhH8Vm+CgvdwS1JI1B
RgA38emAezDplvagqmLKoMeGwKnM6lkmgisbrITLvgBhY7rPNHsML+R9l+gMOlYMnzh76HeeOpj2
jVJoR/KcYOZa0sivY05r8xleWDYN02Md+Ik2MMwhTB9ILvQTXGN4tfX9g2k83UbDl0gvXOhaLIgb
/L89/yZ7DXvuVtIGptJbrS+/Jl3isd5nvmstEPnXWW1woHpB5MzY9GaHVs/ePl9hKM3XKbuYRwIk
WDCUsdyNwxB0YbxIFLhertljB1hDV8PUYqGNbJMHwMozODhNrtrKJOv5ddMy5eiOqhhlaLBDK6kI
C5iXobVLxiG3TywxGeWsOttRML02WZw3AnO35oSYnF59F6gM9OsBgTlQ59zBqiM8OxZswlr6ZW35
VARU03yZFZ6aUxK2b0VTngEC6sq2+SfGs1Rfoqh8FSyEPBwCANkh2LqAbMuZNU8yGBKn/Ve9mCrl
LZS2yo1xmJf5L8xDuJ7w/2qoHAeXqt63EDsG96T1GoPXkboSjPZX9GrfgCeHwB1dV5Ks+K1VvfAK
OgHOOeWjXyAuyeiI6RN6H7CwBSvOLBzI/LhwGz36o4aOvdzNMzDOE5B4j2fWA8WoBydea3fIIqhl
WcxwVonKKwhcalTl6sG+PbOXeOmidiFtZuZ7YVRzRK0G4VxtXr/xrq0W0LOPf0NJykccPCEzenvw
TKwpRhZYXOpNqfJpLEyDhdK/mVHmihHlQ1dG88SqMli3Eod2PySA7I9EI/5oF4P5vxMU3nlpex4C
AK9AoRe+JZ19XgJNWKFXkbx8AN5jJjP8ZoNJBv9Kqh3VWqrZ62g3/j43IjKjp3XFmeWdt3eQiPJK
7ROFv8ft6XY88EkkIDYiMe1C0IqoLTtFCwMZquMq1lRbwd3QO1bfIBcpTQpN0qYQ5LoaGEpS1Yyu
60vgDo/wFweHenGc/kZqtZ3HUJHC+fGKPMEntaMb2tgcnUVRvCxvhb+9twNM2BBGnvAKl/JeRD7m
y/CIykyhs1SNUoNiGoVDcvXY+ODtgheXS+4biXBXTPyFc1QGGwREs6XlN3+vhaJF5tSeSqEu9Dfp
4ctmnPOHSt3JQRNqTwE73V+OXcBTofrsAi2fCXswQtP+lsCVhWTSrvTwgz/jXUfh1cqXESxcl/mX
YIW+zYlfgcchMhCDX2U+IHSkGetXVLwACvbrjHCqy5Q1oHHfcM0eFzwoHj2ijNRhAls6h3FUITkn
OK4DHar8LHrPU7j4/qLpNMv8EH8eQl3FlKmoNXz8c5+6VEquQMKhY59VqG4wFJS4Siuf4JsDVzvY
yYxpDE31s7512ZEtX6MFPryy03dedpKfht4K9/rBWYjFwOYecz1CRCMnZW9r3Gyo1wps9lGvCOdm
AnUy49NgkHEYNIK8AplRbrUt6I4V/fVZI8HK3sfBOZxtaTrOrvxqHskwb4Vbb5xseMON7k41Q1o+
CGSBd95xcAebu3w+LfCJhH/y0LjNAOwAVc1xuoSuOdNw8LCLH7Pxg18zUZk+qCyVMZcu53B/fN79
1jxBJdhiDMPIyYO1+Ue7I3vK8148awHVR0Jin8UcRfdfWZ3ANyvRBgy/QsUTBxs+JA4K42DE4HKo
P8oXXOsSOAuTJ7eRvz67+lH3XMqTvom051PmrrJEJT+uAN+T/onTi2yrUrrunkH+ZkxkQWNXJpay
ccrI0eZ1azQVQU6MFb+Dd+/PaF7n0P163GKtbTIFyPmqZ4yfZe4mSdhxTJt4YoCE1z0hyjozPI3X
DSxuH1P0md25qF8ClmM7D94GgOjlVIY8dCqD1ORz8NaLJQ0hGa0vWc/NDWug3taiJgoVSTs4G2VH
fiCiEHeYTJiXDClzZjy4ErwpV1ce+FRDUAP6EwvEL6liI6k/TvgB1FDBtUkcMtpSuEsNOzBF5RKz
gjTD9nnEJ3uiOwGF+X5+GYliATJ4aWxRignaPDzluARwhHTxlizJMcJ8uXQNjlg2SOBqhEnhvjuG
XhP+S/j+Yk1b4IuDVOgJhOYjlJF1uXKyXYjh8mY4vunO+Z7fmk83XTQl0zgMKElovG1E4dMYYPKw
N3HUkdJTScI9jFGzwyMYwxm4LWhyLyVGUXaqHlSMaXrcIZyQPxa98Vd6PaWnqtZTLPfTXr2UVmaM
l1qhnHjpURIKrAc1h22FupFxcFo3a7AqXCf2pHEYZXVTL26uTeQn+J0Z4oJfKwWZ6AlNYCAxRAPo
UouBFaxOn+vQsKVKspf95LadFfS7TGw68WaxaTiy5LnY3GwW0LvrJm3YWUXDSSXpwA8KnrhdMuGY
6PSpHGysB5WgD88Xo4hdfBUzeSwtdrscrHBEIN5LFcRuAKkJUcfYuS41+xaHyUWxGDoPJGX/vSHA
zfNyUyX45qI/d3muJY3jx9J1JYQnDkwr+AiMuGFiyrwnki/mEd8RP6f4C+KMgzuriUZxtqdaxc7X
ZFAtu0IQzyab3t8mpz0UzoWQiebv3xWgb9UUF2HxvXCrAbYxQjDll8eAxW/FGo4oYo+iELv1Z1NK
Mypgp6i4oKnhOAkK1m6HOr4bPzKW0/XXU9R5eNCG4CdG6YEcx2h3JFUIHyiXLGeKlEn73+CP2rk3
OU/ZLRDN+pI/d/h5Ntyt20ATuJmy6DjEb+lpFqJD6xwLNMYu1YC+OqiNodgCnbO4Vv3VWrcLh7gD
PXcc+ldBQkY0tA2moy1WbVoDOk9zuzYtTsx+3MFO7ks7mzFEJXomhfTkPMfF4AYXKlbzMwbiVJSv
6imhemgni+hQ1uSJp1VVTld6KmZYq5b6/vJhn+PcSr9iyKd1zQOk06KRolT7Wd+3l4fxz9dTk+VS
FITtQETLwlYOkfXXjMJctR39Af/KqIGWDvHKmbgTed/4exYe+sZSWTAj4ZZQlu6scSgWwPCXuXdA
+4Louf0TPBcP4JMTvuTGHYO/2StS36nCs5odvMkhfdsMvHeP9Bfosy3/T1Qxbr/ov5OE2ga+RYvW
FRczCwZL7Ih3xo8vsYBZIFB/xImUU1CQX39isp9lcR1r5bmyr94OfRggxFl/253yHq78F3lMEuy2
MR2M794ybUMotQKq7bCZb5aWlnS4RrWGLsL2EC0nscNcKaB1hai8rrXjGshWN/fg9EZZ+H8R+Szj
M5DV9VTGBv5+2F/fCLinzswkVrwT/D3U4EzqlyjL19cKUaG/R11NgD9L17eoAEkrmkUUeSA2hGqD
GYgPRc9RByonKxp7S42qRFT/Q+SecO4ckPfuY+AaQjM/bUXtNLeRekV/r7efRWeXnNE97lL0oyk4
XTwWrZfpzJYK0Ktia0Z5uNKQQMU/wtlDCC7k55B5o1ouRHtPTxwmUFhJZzoGrsQTjcsOHx2gEtfv
V6gf/fXoGlxRMGLneXanP1c0DIQzXcWBFWKqLrq9MNCpus4QM6DRIcRFLNJLzOUEcWsb3PE+9o2o
PC+2YRLlLiSrtFGLAAdktvXMNIl9Du8RJ/68zPqvm0QrrCucgji7xVfLmFZfStlnoWfxEGwgjEhN
L5Sey4N3jrSYjL80p4tI3nEy3jFvlMR4Odzqiw+xFk/SZFiJsnRZGL/OMgJGjgIP7RVB1Jy2Soi0
NzavOtqaWJIJsSzWEbN4rlZgFLelvWkTafe4vmnE6ja3/tm+wW2ZsSp1I6rUH4wWQnS16qSlpcT5
BLJ6JuAN0D8iwtHEqtWl1PmD3vrSafC/7MHeUIjLOwOX+sFzZ+hXjCPkocMSfEpbZymFq0Uzmf+N
Hol0JMTtvgX3KwcuALBild8regj70PQwqXhVvAK2AiDiEzLs1yGXfaK98pLE5gb1jJeSVJEHVX9A
wgeET6riJzk5Dj6aSPGc9Md2m1tsfOpA6p/ZM+AVn7A/JRiQtXMx+OEEBDTO4N6NJ6dJvwb1alvT
2XRlEkPObmn6W8Kcz6RurdvsHlZlih8angsKzZ1oRyUfwc2VYOhBX7V2EE5nT02WEyt7FmUEXwCI
+pzw1jB/m79h/REw0BZADUTMYGrZ9qYUgJyfY38qqIrsku5rr17Mo6BLlMusmZ1AinQQ3dTunSJw
347TeRWTHwz0Oldo7Mrc5+/vONDFrf4yydf07PBbTT/PXHbs9VWvNeVlmdqSghTrfiF6aAROicLn
ZgcImmCKnChftiG63PicycEo+AYxYVoDwOnBEPuiUgNxrQ7Wu80slxjcTV1+A6rGwJJE4pGONPjb
6mw3PMfoJ3HZgtM+x/rItBvW1XM51j3qx8LnBUYtLCNhHP0x4N2HQoB2xh8fD4NFabsML1Si4GV+
+tGm+PO5Hqvvxi42DEVFbMgC1HvyjatEUsH/u1yhMITmLbQZegM7luQ91nxgPEXJO1FJFlOA5Qf4
/GkmBAK/QVITL7VT00XTbUp+VRkRbZmcm5DAVWkg9oamteUrJlHAXbQoba2VcWj2AhMk78pkJeK8
REDXQpMwPler8e6FFeC+kHVepd9snAy8WgIEmgKIc1gSdMyxrhMizb8yebq4mI74GxIBQH9UenTY
DUc2T6UPELrwn7E+Hnu6z96x+j4iHNRmAQ+4YXunqVDBhXDueXQ8qDoEAD8U3BLBfyk939m2q/tO
oT6ueq4dwztszhFGCJUhariiQHp/CyHz3A/g8adzmB09A8mAG9tJ4Iq91gCHzcXWUxbaSV9BSPEY
qvVkeFAOwnqlcKS+Z/a+WcSopkvolJEYCQe+9qIRX994t5zij9wvEhTCmAuQDdp3In4GI8/TsTM0
PBp/iBNtPKgTHIQgPTQ/25hFIaEQP28sjUcV/PNYssqfYS0KBvR8LmRdLFuCYbnpzPGUSrUvpcWV
PqfAIhGOXXvlIiXQX7o7U+JuGTpjeyEeYBfyZRnBlJKjPwfFe8CCBSWcuDZHSEWS7MHtLlR/27CB
slsK6r+1PyGQHmWUW6/SWSdpoC6NP106Y5Ecqf+CYlERxj8UE9J7xqaOEIUodW+wDmJN+7WYEEmT
ewgi+Ra5pu6nuwFSxHiN8XCh25K5AAnqnTvcIyMy8eBd3+ZKrXQWVgKZWx93ntJ8qT4e9lON6/Qq
wqUmppoWxYlLBJzKzuBIT4LLmuNY1WKJDawr0M5f1a1NjRbNTa5hK4AtPkqBGIP6I5m9xKPWsGwB
croeklqYe//+t/bciqPg9pDSPCTEKcmP19jMSY0lHBTMEmcZ5pA4qbSjeRm6/yzLcBoRTymdKq4R
mcIsniRM9y4eTkMl8JvQLE7P0c8Ne76JhZbbogmD7l3/6Ch7ERoKV5pWLh88V0W5s5cqk6N4ipV2
2nIh4N4AL/fLkWAi8tGzAkLhfv+tE/6uxNjhPPMMHj8he4NPitpTkyjQZmGbJZw3WVGuXdssqzZ3
xLrb0oJLX/bSxLIkSomrnXTARb8rpr+tkJiqh7Zy9Z6vyeJ4F8EdTXbLYbDynDOrT29nAU6uIR5M
qauR+ZjiqvpkMnr5xFE9H0T9LKNLmLK/W9xkfzpB1NT0wv6pdTm74efYT2adv/vg8ehXeFk9Xjis
P3oYFjxuOlsuC/KgwIn/aIiaXqgnU4w1hZ/bc5SqkCgTTZ7jXgdSfPWAV+42vneO5DX3Xw8WMWjL
9alyhK++KqcQJLlJ0kpaZUySemkANtrhl3R4UqTPdMfxiT1OCE4c+87/D2/9w6e17rn9cmSeF7kh
nQ3pIUNfHEzYQrpPFRvUo7f27NwJBLu2Hg5oVPza5vc17ginjyRzG6C/uj2LZcxQ1KAxO4qDHAaS
Tb35h55USKEFy62PdodIbELo2L36HjDqwIHkMQElbwVgMfjEd4ShUtLS9LJ3M16+OBECi7lNqoV4
stHhJAsxm1+/3vEtAy5Xo1WS3MgZvf6AJEHcIUKNgWHoez9tFbVcerFrcQdhUINpfwGh2fdpwPMM
HWEIWjIXLhzuu2HuQNrxiBB64VoYsUT/vppQWY18jvlgRk6iNt8ilcDzkEvc9TGwZT3IEw4Sp6W1
xjopOE9k39ywfJtuBGqZeNcGB2k6EKSCb10YsmISJEMw+0MkIKinp6r5YORItMg97CKA6XuIm1PY
CiXnujk7DoVY5au6i1q24tJ42KJA1evWK9oVzsQlfP7TBgoI+hVMNS4pCu+1zRbX9pxiVdd/HTx0
uUZBAxH6cZqgqeTc0kQx+4K18CgxHwD30oSO1zOjfIUpvgCrI5nLUGJFfPBd1lE1URzExYO1cRn+
w2xSvBxmJ7c51zM5gWzjUiwUyavFV9are/C4mrAOH2SBmRoEMKAFWh7b8BnyIxcZjH+jkZywzr70
r1nzsq1wLQ4iVmq5KSVzBmnY+v/qn2L5q7GbcamjKq1KTFd5I0GQGnIdofoyug3/z+1vX+fu3l8W
ehxUOYgTzhUsXSVhxue7rsHyPcAHlEDrUUzwDCBQsYjBdZtmqYBmks4C2LkhU172EHXC1Ylix7vg
Wt21HW183DxViPHzds15i8DEY4snvkuT2180LqcG/nvcqqxO3jY2R857tUAeFYLaV0Yz9a038Ccf
yI1Ia6Hgp2Rn1X20+6ctCUtAu1G2Oxlo8r3qY/NmvlFq7tBih1WWlznnHzYvEpjyStb/KycP/MrZ
84rCb3JicWldrOlwF6GszHgncdojjo1snuB/nyhA6+qSciKtA9LqTxpzU5dfB+tMgj+1l10wGUkb
ooNvOCdlyjaifND3bokFCrLlgrxX/r5XKU2tlvpiDAjvzD9CfmE+ZMx1p2Sj8qHE8W/51GGk1S+N
lkzjy6zTOnWXDdD/EYD4nJOn/GVLzAhpJ1vTXQBlqW6HSeuNMEq42fQu+KgzANNhUZspLNCQzOjE
S4/hNr+iBSReG1n5yiuphH2h2aV8fsZmIYy/t2ENSI4HnJ+P+713mTfiNwNSKgjob27d/1pL1FcQ
uBI9OdA5+5zx8Dmno25cq0d62PHqUipeoX3LnFB3c4nPwnV/PKcgWNwl1xfFF2APDI0H7I51mi+u
U7vpps3zCSHMHCeQjy7KbxvLW9bb3IE20TYdJIdHPWC5EN6tTnlQYy960LjainuZrtm33maVMd/R
NVdc9abDzc3iodiwka88g6B3XyJ/1Ax/JHgPz3+6WBv6yzbl/ItfX5ME3QCRu5i9t7VVLLeX4t8H
8mp+stumiET4EE+WahiO55UFtnMaQNdiqmZJ9fWJQUSjFjwS7scH+zfCmRxJWjnlDgCEQOnK6SQY
rMhLT9Zxa7DkUq0JsrWN7bb0uKxNoaI0II6kdi7D029oK/zGP8onILEbUuGITRjQVMVmj+5lPHDN
qhs+x4Myc6C24cDK1Fts6272XVWzhLngzUahZULsejrWlgBk4oOGxblHFqM+TLfMR6rbWl8xJKDn
f5UDeJ0h47hhui/DNDFb55xxBhuQJJoWEfgWrl48EJnA7DxDCFhNbdDt+/4MmiYsKVv4p7tXobNp
tVFv4cviGAykt7pHHX/sDcNfwn9tN8XmIS5IVpPX3pE3MlRK5Z3gOQ8ZYU7fn6WuPwuMgeyZFuHa
8eGy+qjP7h5N1+L3V+FGT5kelm74vpwIn71Z8FOSpx8G/L931B4ArryKyraf/fu5F1GEYzZdoYq/
b3WIxeera9Ebor3Sd027XIfs3EcJaxXP3JNBeMH9W6NKD/nL0im1dvspw8MmXy81cIVuYD59e0na
1Mb71WFPzi6XdBpLOsat4vTVkt+BwDvLLyrAXctXuRF2lYI5kmjoP0eGy97KxrHVk8sZ+jf/krpE
mH2Mp1aAtcbyKsb9rkjU16SNmgx869eWpHe5mheM59My3uBKC/m/U1mLS5/fIRyovwgUyQ87LDBY
yFry8xl1l/9pUOxulmhhNLCxAqSMKQziKPgDLJfaCuT/ItDqu326Aeu7QxiTdfZ30gK1rxb978x/
/gaOJqZt2EW0oDsMYYPrDKc2y0uRlge5nOc+i7jQKyjPq38vDcVwh/sxbZsIkrIzPlIOr76PiuTH
LDosql3GD1Ahv7xOvT1Fw/KwdAayBon5rjStabqW9EpQiNPofmlfUZHVGmZxze1Hk5+VEQpbRry8
HWqApKEz8KBVw9f2Y3eVhTurUSheESQyBNuc6dcLAyA+WqnNvfjZgosePgA0GNG4ivMvLWyUBeHV
dMd9LebHVHTDM40UObMFa6QPOVVjf1i6/CULrcLZfPSrGBvb9UrhgdzIRwXxWaO2zlYfqPi9aQAJ
EJjorVtkyeKMvEoxov6RDz1Uz25f116BaQr5UETv6FA1KyEMr4j/BqS94bDa3R7VHnAz5VbM/CXE
lKOoYKW8At5GNDfdWjh883gYFmfXZafOxVYnnEcCU5g7S4KewBS9MiW2hKyLKdbOAtSBi0E5sU+a
m470xJBzUQ2p4Ni72auBWAn4gUmQ05aNrccEfYZwuipZ8JM6q/h267S7caiW9C1KvWPeERzkinAO
dXTX9hefxmZCpZX/p1aRe3XCw5GoqMRSpnyRsKdp1hIqP55t/zcZl8X5zagLyriA88WT7dU5Ca0h
oY4xoUOi1my/LdKDElv979vPrGXvdtB7ASKVf++C8x0Mflh8gnRTSCiNB11bIjO1x8U6Eo50OgX4
6Hj2moHGogYb54dN3nVGl9MDmM6t9HUmetih1gUTQnQl+DBaCDXSbgkJODsKVqexIcXADbYFYUZ7
1bSOtFxuXZtD7A4kgADtZHa/A8d7b+qVgjN8cILnhq2mAuNz0w/jNJZIQIpPUVfofIq3FLYp4Mdc
raciOH146ep3tXSKiTRN4TiRUyTRGuJq7+Dw8Jvhy7XBRedVdCCPGr+sR8Qsv2k1SGk1SaMMAgFc
MshgDr7/mcSw8szTg2CZdQ9VS4mFoBVCQ/oqtgQMV/xyjXkvKbdGHgZPoA8V9ubM5g9Ytj/4T1CK
DPf0RKOPFUJu0YCR5VIpYrv6ugKdSFT77KfMX1ssgm0cAsMIG8aLcpSYW6rDUBCojuWSMVd2SPzB
RondJn8Sf3BX4F/UZ3sCeRSj4RedNbhN2iJDcSBTy236CH8GN9YexDFe0Kyhd+R+ArJ6LLQL1pFZ
MYsc3SX6pNCKRt/Ao2O8IPkY1fHnEU4iCf743VZQozgMpcrDPh3RSYHLeoEd9ImY9XT8tUWgRsGs
k3vdm7tMN7OIMtEjPTIWNgn935U2lwqLYTqdmVw/mWKD6YUaNATOQgSz9Oh/M+DXLAK+HLif2PJv
8jh7fiysNIZ3cBHUVIqeF8myKgKez0Whjfo9GVE320AXFcIxGFjAgn7zupBwsUizwEQ2Dc8plixv
CA5BlpioEXBqejtJtoXdhrf5dfgutNCf+nJkBRkkpvMIy4NqFk8clthlmjszwVSLmvi9nU4IJVkk
ntam3mYwdu5jR53GdVbvJkCc4XMMfSEqPWdnIUG7pqpAL7XJGRzy+TwA00JCr2gGEXtH92s70TqF
+EiSpCjo7W3sr9fxNJxG6NDAMHuGhu2GThHAZZVyUS/VchGQAc22+0mxpYGItyEa5tYYHji/zWN6
s43yFoR9yCn0NYgoGGdoRFXsxV8nOmFj4fgJmsDWI8Qdchn4WfaMAKd0YDAmAEUvyGgkQKM6WFTK
8EOGbaSJy03YpR5IU60JhyJznCx1A0fJqE+lSCNgSpMF2y5s4VQXlg2E3SL0k2TR7oxJLNtyyIBs
c7HmM8fvGmHr0BiHFE8lY8zQ22H5gvBADB0VPJocp0ZtUYAJU1c8ZEvppYhFhDee/99Otx+fkz6k
x+zACSExMcdVmC9O8ob0rE5mlbsuwlbe4ZzQQHEjqhMqIa6r4LZsHuJifLDnmAJYJS1F1+gcugJq
RMdNsmxBBQIMeQWKNB+1MsCVakg0gzM8zNWIPifI+4cOeYm3AgHRsoKRio7Jh+ngu3XwH/h4gVSy
ATtw7hbg+1UtuoAgDMqyid4TbXzFTNt8v2LTSnBgHrcTJ5JbFpaUdVdg7WLFt6vOBsWRWDCEBIPb
/9Nz0AjBfOM3z/Rkf/qX7vt+6qrJdnyG1Ui0Xz09KqvBaDrAtkQDmMETupgQXeXQnWOJ+M86RIyp
WG2h3fPqbJ4gGAR136DZFLq1lxl5iaS5YIhtMYmpUTYreA7VLXkyap8jkDq3gRZQuw86VzHmuQrw
J5eTIIkwCrXO20OkpV9RST2NjXIMcjfGyZ/KN3Ienb+kGXmBIFI3AYlcJcOWBogC+TaiLavSR+Tl
RzP/+Mr0lJ1Ez/MpZCQJj0/lGBml/QWfY3kpK9I67QSbpnM9QeFw/ZyZGznuATy2jzjK4JTGWoKV
cNVCpiAKYqIyNXNJzEWXywiBtm2dN70MdAYliyDUQtMSNmct/3xNuksEcIrZ9+Oq8yOUSsIp0hZg
5xVwqit6hfKv0OGGoF6u+bgNxKBJyNSHJomyRYs4wRvyx4phTtn/M0DkM+/NPQgLuid1tDmV7/lF
aIbgpctBabjucxfq/8EvVrs2C48HizbmtVyFOJO2TzlM4vJe8cIQVi1vDAp606nq8u9A6WiQzXHC
rCqaGShz7D4jDPghJAmYU9xderci6LW4SLnuSWFruoEfGCdEYat8AFylLcVPaiaxqwC+vwUvpcL0
AJPtjuX5PWUnQ6hAiwziYsyATC9Xr8XfYEMMYwekBgHliABuJd11QSxPIeMiXPSC3yKDouWxZK4Q
xfI0/yjy036na/OiPATsl/x/R+Lb0PAmwI+AxYDeJg63U4LGJc8Ak9fISWfPKT7PUv4y78i6F/7O
Tn+ghrUsTwa08OA99TD/3u33hjxNA5Ti1hQ5EEY425tS4iMuAf5zLJ+TZeJAqvbrDvAW9i0LG8f0
mRAk+KV7vnfCJUv402GOtpLbALPe/5dgVCvawqGe8vkfP9JpEcm8RfgvHLiFvnl3KiONGKOtezBJ
USPEMvZHm44rKPG+BU0qluzUt6djlwDua1KwpJlAf8x15ajo0LQ9oktVRJ+sy8xI3XzzTdq/avDd
s9BOE312v+y3G/F6ir3NtkjfKsgDTfep8xAeBmZ6KvvQesn080XRhI9G11Enxvz7Kb06DThMrFAU
1xzaUAwOlQcs/Z1wio/eED+e2sDPfWtRmPQInc204aQdQHGvS3ak96CDIDTUjB6llmiN1m5GVgDr
bQyexcVwcEatfDzwjQnoUl0M6ozkZOYX9PEdQgkCR245t0oLYNUbrU56rlUF+PpJsHmyDZfKMq3m
AW6GJOj1bqf+UaM1i0pWWa6s8pGiOClLX1/SphULgtGfsvs644JUymCjLQnxT/xLgpRZyrfKCYST
SOOp/kCE2DyW3llN5sfN7xZknFKX/eBQc2VYovveWfQGT1HxxwyTgyKfB9GnaPPKgLulnCvq8joG
BDZR0R2JCZ03LGNL2LOROo9i6w+8ty9RiQR3soGE5KGq/010taBuDMXj5o0p8e/FiaI+mbgzSFIL
GRwd+1BQVcaCmtIEpU0MdGpZTS106JGUaq6nXVOS9wRSdnq7+pQ/zPqyE/r8k/VZTknIRJm06L9u
08Q/eV7MMedAv7ZotAe+xeFutBX05vBL2Z28T0qmLsnVnDW47C5uvI/6cL8MjWvzxf6DNdb/zjlG
lTK8lySuRHj7uiI3nN5c5e0N+RPw2iVXk4/T82nLzsyb+iLWsw0/KZTsKMkSTjzl6u6CCB2CmPOf
CjbOSL/AXbjqJ9tT4R5vBxfq6p5s4sHnb4xDvZBK31Dzdso1Tc56ufe7DLF33ncwr0MHkXepiLdd
d2eEuMLHlMpOCGhM0tuX3IF/cuEaYJV3Vy/KddasDXHt7JXjk+VLCOscR3H2a0Y58xfydzDteZP+
gtVzzdnnCU9Rq1o3QVtk9uVH4yaIGBCxujg82Df9r62vwArVeHE2jCEfuPNK/D6rTDIdduarZyMe
zmnyBJw+K8zKD954jBRdcklUQZs7ewOhc3drfZtvmdYVQmuFOIYTLmr2rw4lE7iWZGznEfQl2HeU
f6WjtvIEU/c+9i9pGc49cJIqlXSKXKoQjay8CqMMpwtRljhxL65iPlWSZCAzXYJrzVGz3iXnDXJR
DAVp7N1BeK9EGyIFc/idkRGjQq4yQ9sn8aCK6P9HdoBp2ncWn4ryB5mMoZdZAIRIYriNXuoOgvl5
sEpTaDJ8yvRf/aszBHVCFhr6IsVIbmZLV92ptJcvPgUVLggSnf6xWbJy+p07+xEbSMh0pZn4OH91
uUYATNyczvfl5jQyMbsCBJiHuDE9t/7N3KQjZnYxF3RrtY3QncaYe4OKSfx+4Ja2TwuKAv97+q7Z
sw635YNZiX+qTtKswu5kfADfjQgRSqbRt4Cgf3GMrBIwet8ofc03rxjcaYRxBAF37EupbGrNpxs/
CJogcFc0p8mdm7IgFyo9hmhX1FBm18SyRgErDaWHj7+fLK/etvamcNhKt5XxP+OD7gWAbjcn+Hzg
GZE8njvxNka05n6VhyBsDgGRqK+vLRHBxLO/8UIX2ZBS5j9f4yMlFYbAghu2rkfOhqGZniM6lPcC
f4Ob2BTy7NBJVOHvwsrui50UXJK4aibwX89T5tKic2yJXONUbItMsoqSdYvnBs1/477Dut1xNQ1v
GdeA4GY4ZVJsS9XKzp4Ci7UzZJk0GWgMt6Cd2mpmTEZWzvfRSIhvxS4BuBxgDDa7Bm7JDTKjWmxl
1CCmP75Lz0DQSTSEwf7akhnG0WxqLKbjvuSBqVt4Rt6vV74h5HfV1XBrlODOk60vIXKe31ezRn1h
/w0cu7j3FBsPN8BVYbqQubcP5NlmsZKVeB/4qaX0/ob3bZggiRxXnwiWA8wxDeygPjGSyskXODG9
yZV0oTLh3ghRBkFDrT304kbAXsMXvfXoTqc67rUu9f+1eFXRRVg48R56c4edGM8gEl24lUIvKyZ0
glFE1qYUFwHUxIvX8YE6AYE5YSN6EpT3Vc28K8Y7CzAWTumO7f/5Cwak3UlGz+jn+Vr7NhrdrJDi
N+EGtIbpyE9zMYifW0TB0XfE0psfaD7LB36BCrBtUe0qVJ5T5/KCyWu1i/kPJvKylJCipDNOEjpo
Ck23tWbB5gCtO/Ma8wgXglSzsBL04ccWiH/JvAifKLxhZbKFakR3FFQ5PT7JZp0FK/3TZMgsIPzT
L7C5cjU3uEZLxdUihmHY007olgFUG9Caw99q/Z2n53ynArlkAvYlp6nHC0dh1KB8zoKw4DHbNd3Z
Hc5SDzX6VnQRyJFQeMn7kkOKQIkmXoSp/L2rFdC71xWvrcB69H3Am5560qaDVE7XfVP7OC4Zdswd
3ZzFJk3zd4JDYzkTV+j07tqq2UdRCmzwnH2RHdrQ3LSuLMpukQymNUT9rUROLDihWRA6rbgGvb3B
c56rVzNqCJ1NYIM7U0b+NznqT5JbKp5uWqi6nCX9w7g1ru00rPQk0dCPZoly2ybVBLhufjmJsEcp
wvjS73Z2Hzf7CGbqVjn6g7S3QCEsJvXNttHetxeW+0oI3FJhomnrqOLWM/1wRV9rQNTZBd2kuyEK
KqsC21/trO2qhSbXCHbc1KrKfrfHIxNUVlWCWXFpzB5K7NJ5ddIHgw5HjWEZwRlm/2G8wG/qCvFk
XHyK3TEdRa/gPA6s3klVNewvTA2FMNPEHmB08C2h+b/R/FXTeoKcFhOnpEfWvCd2rktCnW3YOTBk
AtFHhiqc+iBn7Yjn/qUOxrp4GoVYnsBzDK5SFPynVavqOtokfpq1kblmKJ1t6yi3v4CYyyfbsbTt
ZGdaxfI++p4l3KCu6FB0i/fKdmVm88hDJ8m3Xk/CLpQbigNfQg6Akd9VVWIS7+1s/Db0TgTvKjfO
Y+9PUPIG8Jj6Coktfk3Bzwo3GYiz0PKeeOZQu29gcCAugwxQ/2xDHc+vSF/c27ynS7xZTG5H3QLB
16qS6ve9qDaecLpYzPCaUQEN9ulO1Z1ozkapvt2nSnScDiGujgiFIHfDzVFWQdwjw63b5qVfoTqq
qzhWjZInuFTfdQDq2+PGMvQgfiZH5nH5my8OG654r2fuXXeGpWU2wvI+HLbW1a1isTMDHPnaVkib
J+ywfcBxo7wtTjuWH6lVWOPHgLuFhmthVooKr7Af/ErCIL2uiT5SlsAvaAACtzu5PJhyBPbQzN31
u3EUNXvXpoWsBStqj8OGzEz367xPJ0lfmC73par6dX5DXBG7VYhgzp+RaoD1o5cHxfF/xhsCYg1/
uqkWSs+VNyuqxNToStq52XPnwhYS+poa376Sfx2qdR98/QOi3sHpiUFuOTVLUL0dblA4JpZTEJDg
PgeuPLL6keJei+vcMy4EMW+fVaXolOVT9tOpQCeGvnydhskLTBtYOE+SmChIJHx40/pVMjXZYNz3
ehNr8mZN6WE3PbSUEoNph8v0tqDTA/zCgnj3s1vA8k9B9G03t13PFqilHfIeKqWN+FRRWJ5XJwNJ
jK+aaVQ6e37/njvMB1nQEM6v2OW7pAId0z0twuh6lzxGyr2lcn0Ma8CZ/RjcPZ2xXUeYgOq97knj
W/QSB33nYYzj331uK1qtZAkAfbBuGCtIN8jqmu+9jjBP/qDttcI8Z6POWJNYYQVpq62nemsAPxEn
hn4Dr4ANwjb/D4TmoVa09GmUP1Ta4ISXDjAjntHg5dGO3zoPRM7AGt8Qm/TPQhIefn3EAaYSZrgS
GMQpbkKTEheXQD950HRIWN9xtU4pSThDCPRLtZPcVIYQLSv9kkdbVpV0dKOtwtw966jkZWm9eh1s
REkqSvNiTh3rRDGTHIfPuLyyU7bM6MRNRhwbxSbUpUQWlF9zaCES6ceoJphQB4GdEXd9iiZYwjJA
m1/qjOm4uImMA08SbqCSJW/17QoslT+QnM8iTDogG3d61TaTtJM63dA1TlIIn8CLqq/8QXFok+uj
A/rnu5C80CMlk+QcvcsgbtntXylsg0uAyMCsk27VU9x6nG+ltGcL+9M2V/RBzDAp6TG2abd9nJqG
idySC6lhXLrK7h4sLzgv+oMCTR3dCKwZsnccSEuRB6VMNHdRe5KQsqikkJMx0R/gSwZsoVdOWPVw
ZuqssuTAjdZbTevxxq8dIPBmh2M+sV0i3DMuVwxTK+pQvnGER/BHdGb+p5HQPy0xnwasCzxEmtOW
8G8LBaTHwn2C8YRS4orEClWsa3H89dIUbC/YaOrymXfbJBqvQvn+ym2+lEetBaBNwfeKmt7NkdHu
nG9ywnjqCRx6iFPIYKVyUKG5rHHrZcpp5vyn06DcsIWV9PLuT+vgJoygPeDBU9JceenR5eFZ7ZjN
jA70clvxE4sGBATXMtSXeUKv25gDCVSriMskR3LIuKvnR2Xd0JTzLmO0dC0SnuDX1lyrRLynQ3qa
+8J4U7oruhsV/kZPv6p9a3DhxFLXlkoURDn2r0LCFkEXuQO234Tn3o9hm8VR731efOAStsURUWaQ
zHjX+w0xj2ZAbX6HHvq1xSvDuTxG6Ou2SdyIsz8g4AP+0DRI/lcsiAmyIi8AsiHse6b5AxEo7+EO
tDG7TsxzjEy4vKotHGooBjFw2ViRHuzWZFyC2LIwTtsLavE9oeoH8e8pNzIgxdLZHb0peZ0sKBsG
sGW690FxMwl+/bbCKr3dRC5hBxE/YK4EezW8WcRPmeCaUZDynhnlmO6CU6iTCbL1yHCVK17Cx7VN
VxI7wjvmrNdaY14K+NyvMss1U3n9lXtfGefZdIepbkgRctNC8hYvW88iFyocnw03rXrXczRwUnlS
P9jxDZ71P/QY6N9II0J1jxGbA1BpMXQNFYjQZ+U47lOwGxgK518viDYjhul1GWKrvj/fmlMnrMXL
nVnRXNXbX0VxFVigD5Ah2ME3mj2PQ7ltk/t5+AsooBHV5kaR7rDO5nOy4Rq+dx5S/c8okuYpgMON
XKTjAS0N4+pD9HKuebwAArebWDotF/xYR//7HCt8pWMPwy5UdCW1ZKMSSDhxIJRe+pxf368XQl3K
iUJhRyuTVxRHBH3A7ddPWp1NFIWuC+YWYpcuV0jnt0k0ViwmLSTs2V12o2WPKb1jm5CYYZvzc1ew
7MUoMD5lGLOseBSqBRCahb56AyDT+KBDS4ZrLcCN8MV83WUsObZv0E/dlS/JKWarh51njbh73rFT
Oz4y3byhZQiT1qFZPJ2dWQSjraEHX8yl4IMpT32sCPaOEOX/ky6WRtSNJQkFo3xqbSYmJI3LJVDi
fxkBA/F+TaG0xXD/rDSHqs71w0XIvt5LU8B6WYSWL1sgIWX0vCVEOjc5DYB/Xro/b5Y7DRxvK0S/
Y1Vm9IVcqsgviaJZJqIcuPpPcvZMJ1k4rcpsD+mnJQg9XVAmzM4zgwPAiaSlrkf48ye/qqqpUdIJ
Z+ZW3dDC8ceCiNpvAyBHRR5yci/3ktpV18CskISLqWPNYfQik3yOVy50eLdZ9zsposOrlpsaqJzO
Hqk0TdKwUEwZPBbnhrEVgeaydwiqLpfBe1+iJ6PQ2XOUQzYz2oai0V3CYWmYL9dPEqphCnhb5RWy
iBNq/RZT6yv0j4XRVoEgHfCZvEczSUmhxrvfsiPBqoSDuFxK7Tfqw/I2zszdkRqgN7+t9rd98yz/
sgFFI9rGTFFij3YJJza87BUIEOxuiE2VMfDfPNLcQ3vSx1IZoi90Pjkdxh3c8ZAALD1bq3Q9RkwB
Zajr+hWlMcOLj40Cu1U5kAvCS/j3mgjnGKtx2ipHrcpBA67ZB9J76Qnkqv6ksW+Vdab5tmxG8/sA
RwQXNHzhfC+5XkV6a0hK1bqv/g24B366PkJs/AbBhGKTgMyyDtc7QrxW1EvQjL0NpAtd0TuQ8T24
3ePosk8u10HutIEHGOROLEerV2BvAdnJCTuUs3kfL/mtK8ky9MFtUquvg7ka4Xt3tt/DP8ZIdFeK
yarULYpFeZaRpKXnANA6r5MfEzGhSph3s3zcDDpWhFensgK4dnDc0sWrymOD9/uZ/mY06XgZPbpA
m2dJ8BPH8AaZLmTdQJOHwHpW6uNKi7TrMSft6tYbJtx5jb1xihU38XvbW0R7cG8LyOrcw+HWPgX+
RDFWJxaCK1gCRFhBPSyZTA8VBPGUfHuDalOAcXfH1O+0FwRW9XqwNC8EVcJi/H1JNBdaDctkIZiL
lQq5lQLzb9PKuWOwenzxH2s7YpNrJSVVBr4Q/5hBLrrIqtz0tYnf0asoWed20pFw/Qew9Sc8n0hX
zc2CvXQMSzcxHO7fOzNeMoA+bfQ9POTljmq+JA1SZGMN3JKKMl5953Ci55tuAEylM1154APREBRU
mEHrbCiY7wl6IinCZqhj4C61/yOk+KVw8petMNdhYChLnQ7G5RDy8mISSKyz3vTNstOqCjnJg87l
Ma4Wsbinn3IICL1cKwtqKImX5Y7mJhBm7gf4PdiNrYzwzs0bqYg9W53RPVVE8v+Ynt5+4Dnv8LTv
phv3/3ld51P3ADCCin32wLZjsKdtKwPp9Xl0RNvaI2uksUDd6xnQcpab8RX2c8LpE0DxXY+j3VUU
ioiK8VB6zV+CojZktnqfU8eOWyKAalQWo6heCRoQtZuzvm2FuW/CkE2vM8ZHFGNmqyaELJuPMAUW
BH3u1MKcObxhdpa0GnkqON5X7iVVlanaGuHUjO6bewThamkE6Rak7kVdDwY0SchksTLe4Rt6uFsY
ihHaCBr0QcteQyRLQsDxLsk1nBUZqch4S+ggm8MNUhfbw5rOwLz44Jtni3YbDmW8dHECSR3m4z1h
k+TR1SMLNUIM6B9r9aTbdvC7uVBEzPBVksscv/nlb7FZcdsb7S4b0ISJlskPQExd8t0Ebkp0+Oni
zHvu/qQg3FILB2SAmgP5mXpXxWz77Lg2PEerBqCRWQm/zIRBiMQdwxakloXsaa/ZTtFuc3ZorZR9
ntsFs+DiulSjglCmlFsXByklmDvK7hSkzAvL+gCgUPUlILmQYPzDbbwRMHqpU5B9ANWpWDQ3h/x5
AsydQUU1sDZ6KN1ekg14uXm3utPZbvAEKfcIF5OhnujLHU8NcFMPOL1AasDvhpjD6Upsrmn/idjK
rXAhWE+V71TZGMlXqBJA+jtgfCdup3EV040eGXBL8PgWBbsUCMRJ5h5WC0l3voduzw6ZUPzlxgok
qJAJe1IuVjb2kfd0ahtVciE9Tmv624VyJ4zM8L/QhSVBLDlhXivy7edis+72J3Jm992TCwQLWR1T
5IU1G6KIz+q7qCwobTalrkJ1RuSNkgnVGHUj20TGKgxm8+fivmnNscfWnoO16YVdzLRksYIgaLYS
fwe1UvPPErnNwWETL5FK/760bOpFMMvLaBuRX/5CzagufXU/ikE7Q90qZI7pQRuOVur8myFFHMNw
BjWU1o1N3UyMNNV9dMiGJCGxWMXjQ/EuUK7zgDa7jD4f/Vni0B946Jq1In0NWAqYfOH+3A+Loajv
Uv5+dqptZLsMYatEenwiAzNVzPDwgQ+rCV7RVc47po/fDWBQfVOdpGbgf8Ph2MITxUCR8nZPEqlV
+kuYemxCxXPtseikvQQDdQudbuSd/cyHWE5hIJhR7KEoEngXnqjOfypdG420uPd7Evz6hsRghxlx
OY3VRk/hkAfPltMipJU4w5E7X7TtllI8SbyVD7bwziYMXuhxg+DediMMTd/NLPIv/IdUPZLjkhcU
nqoD+THC6znDV/ICuJliDGWYZsh3QUdRYEpTgzS1HraE2MUaeWW2+zANqGvZN3RaaTC7fOI1mqoK
P5+1ifrnOUHRmJLzNXxBiqUE24E76nF7H7nhQn931tOOCULKBPojk95+UBNMFnS1qQ3pSwyPxnzi
h9Ek5TjeAdTf+nWW+MAHPpGaPPpQNskKr8R5tWzHzmft5Zmi2+fz8cSHJhMr+5tzY6ouWwHUnAPS
byfNeHkWX1ps0A1WFDWQrC/0uw4EZ39FwOUU1ce/b+uvXu18ZgQmezJGo6SK1rl2hhwrVzblRRzm
jKpIeOw3DU6LZnCSrjOp1oor/mt8frlpOwgg+34QyI2kFywY1S8EirAxmHABNjDr3CmsYXYT/Ram
OYZ1wwG34CXz9bInGFYB2yl9yR6PWznFtdO798gGFSnAuR1ML46KuzMmqojAl3/LTL0jfCd4BaFB
hU6IK+s0YC0RC9DdPZ7ir/hMLXw2Dkvv7Q42xOPwAlsMYC4tIDkREoRd7I+hbxOiXILau4yCKtQi
gdEOIaHTIdBxCI0W6ux9QJKoZ6PEMhohsGYju+zz0RCgC45gEy2zw4fNYZg5snBjkTpC+xtHdcm4
+4HoUtyAyinbc5x4UvCboz62RfD45QxUGR01yeOZy/H3gGMa/f1cR2o002uB1hTH4FCCgW8JDxLp
TDoD0vGQNzb93g9K0DxI85SyOkKdeQh5lgv5q7ZeoJlP6EDZnNRnSmGuTLkHWox1tumm7Fiw9qPZ
SCrxCagfgOv5Gf3i8aUzy5zJhHJAg5XtlNnWyZD/nExYzaQ56HB7hPoNbXipCI8yBXyL1jGFnQHj
vuZPE5g1x/5iQg0cUWNaMVduOC7Qldlfh4C64Xpoczoh1MQ7mHvKbIQM0DdUv0t5YbxUfDirKvjq
C+HAfx7GcFF4A6iU9ltm6yHZmK+RX+jru0DRSteJjXhOh9v1sHwXaO0sAiEzOErEyhvhd4FR3kDg
lQcMvoefcR7Det5vepztAFQ4TJmldn6riEFw9M8P2ioh0gmRHdp7QjTHpdbpy0VZKsMepb+HCycq
stjrFY2lNTTCRdtIxkX4qxnnnpMRIOi7siAhjFW8fUQH2jNKj0jt8J3lGrBtMWWBASxqpUvhk+3d
NPXphzGphFK6EjfefC6YiaoerURpFcWpMafzZFJ043coMv0O1xGQojITzUlcrf/OCDKyoUyo7BaO
vhxy950LybGaNvIGWfxyL6cK09e4L7HnigThuCnd8QjHlB/ppWKQBszpYwEm3wNhpLJ1Kei3G1r6
0WeMnRW55N/b6xoYaCE+/BQfJq5paxp7t1aGYuMBH+nEcAwLvbAoRk824ZgPZN7YVruRs33bZ8o8
CCNmzMlW2CrtLKWSNocrbSYLIvPYq9TklPgzIu+iouIs2CR6VKBl70cKWB9MsihyBjdAflLjyHZK
KNJhFSqcNQCQEjzDMNIXF4WgNtRhHcsjPdTKOu39UsvwWSaoj3M+p1yv6U0GgwRHGoRZdkGfw5eX
FenOgX39LAydpEbn9IMnjPmQEQPQnLznS0lvc/Pt3ceh08aWiGW41Y5n+V0mtsMB2gYulceR3HqH
CvBbp5ZRlH8Ez6aqji7trrLrNgd4WTcESrMU4255eRL3vgX/BR/8YZgIiI8MQEfy652bKS3o1zV1
Y+aPeLF4dapgP/vrjKiT/qNrBl61Lik2+R8KtkfDlPnJ9ZE2dHJKA+OOVxsaxc4w5+Zj5Dk466RB
yVaZ2eHlv1NwcQZWXolHUuRKHtDziuts/uaH4giQj2hSjugV6O3eYttwsDeVKX05BsBufesN0kP3
tIZbkbDCtKcA7+pMK0RODEAJQeOImSZhnNdMFv5INg1bVXl4ZLcNDCXz0mNPiQW6gyFi+3t3U1sS
HkO/zqPhehj2B5XEsabSnX64xVsEMnPmGR/apKAUpMoQaUKaej+IL5l/DfYwh6d344J3EM98Fdwv
Bn6gndIMU2YJEz7+uryZXwg59v0CI6EpbVoBlY/pP9F+q4j/oUct2yZGk9VtZP5haSH8mEEsBSAD
hKlkYUU3rgY1ZYFkIOCqMJ3XvvmqLiFMqt4+e+vQsQsrStYqNIiofG0gkJpCHMvrbcQRIUYi8RH3
OU81UYrolHUUy7uF29uRN3B3wSRf9gA85jR5HMkAApKeTs213tKwwm9G77/D68YdCjpnwt6f9Qo1
HqV7PLxyk/bgO2h1Db3oqXhDF50IaYekuF5qczA8MM8QG6lNY9rMWmmeIOXQUzNH0txmaAsGqyeJ
oS6jQIRjEipurdKudl3loSU2d9G9tKoyiZXBUKBhn7tqejSPtrxsKZpQUtVmx55SpZGyZNvUGmdL
6Z7is7wI/nEGePqw/qi1WzA7VvwfAUelzhZUxrI9Y78gMjpCtpIKzp9YqyfongwP/R5g/0HmO/OL
M5xqqiqbyWNZPSrBMK0HyPiVmjkwceVDTZvnnvmlKv999UrgkYhTcLVG/aypaKQ7XMJB7sYWpngv
d7kNhjxFREVczNDAGND0h27K2edivxisLDsq+r+BOcEBYHeSis0xDiYpNpg9SS+v4T+jet4lFHb4
RsdkZ5P5qZd97et6gNNizfry4+SF3O6E4eLvxazs5+xl8exm4VCjT34dSPGuC1g/oKbcnAeaq4RG
mgsmjUBca6sn5TIQBXnsAb84Bnn5heamO9enfpygi8II6vYh+2SE04YB41Cn89R+5LRWV0iQC0Jc
tXF5qWEhctyuzzBojnTCsjMRMdSraX7H5Gzkct/heXHrAJkBfcgXytUb32JWKVtJ9AMormHPUf1X
4LlRo+XjJc/HhRv8ZEzPo4r/GCaJzgpWxikQUYNk4X1d2lzKOtG/594K1td7AFfhACh9Ps9I9ANP
EMu+RkPaNIPZTNjizGGYtI4bDwrZuNy2uXGf+BkgiMTjcEzd6f3p8Si/okEPZM5s8aBRd4LE6S7a
3jMKejgvEbspU0mX88KX1uTQOpzAxGEDAs1XxS8F7EU0HiyM2zCB12VpRUWPn2eK71uXqwGBSf9U
66oN033oSsZT848VRGo66XOkcb+taYxIr3aw1JF4VgVVID3UMKRqrTABF7EGxEbx2eG0bZFUVqjg
Qvygwg/mO41FelTebCngr9tDmaXZ2XvIln9sSgIFHj4Za7Zj5IQc1Vg9qMBP9KEY1bjMSdzytszb
LB0T0eqGrV4XPgnQPMNEhCbKHNRO6aZuqZhC1HG8/JBa4839x8lS+EaVBONTmKQnFrrOBF0ml8RF
k2G3wiOrhRNRVUysjU2ImRVQ0+71lFpft1YNdH1S0mRJTAT0fUTGIjhBFYRsMUafSzmdpzxiKl4g
EcgW3ex0vbzozurgq3nmRU3wMKbz07iVzGH/N9GqAaNI2nSJTvVvPaFGkAkjb4/mG+VYk5bpD8dw
xZbCpWsfO0Nk7M+dNhqhKpOmkvW2WMiqcxsmPnqDYK69vOT/bwbU+CYDkirBUlOwmCdoEML3JwmB
t54D88zBB4TVOlgPiP5xvsnretCCv/LjSAvobkKZq7jqnpHlVMBDuYD5N9ec6BrSd9AR6EkvrAUS
SJvJadWizX2K8m6pQVToLrPKy2j222si50F3GUZ1Y+FUf/rW32/nDbPOLxVSdC7Tx86TWTARuaaL
LEO7WNPb3GvTlPY2CQ77bS3uS0ax+wN3a4qYTWMahdqJkrgWgTYyx2V49VVEK/czg3FtyKPoCMVJ
wkR0NJaCmTcG7iwbDKuugM03gQaF2EJAulgHnfkP9oyIRamLAR4T2DQqE6hl8WmumsTZqVAwiaOo
/snhUojw+5Kviec7o5KTVSr2c6WFC4PZQfk8QQ0WPgdTLiDhSz0M0lwh6+n4N4lu0iB2FuyvDkP/
/yCs1gHOMyE75eUoUrx8KAWL6J9oiI2UgaxFRVeJYR5bSVQk1vX/o4Kn1AXaMh6Psx9ig/9YFLEJ
R5R2QRY80gzbIxSbdP22Vceuqto0j9LOBe2Nm9+x3yUfsls0iXccwp77tTHcXcLWX362vOLQ3vRs
hMYPUPN15L8ICtAc718fGNzo6erdvzgXhZwh2gm7m14AIGkagIXhnyy1uGoswmceb8OAFWitVKZi
ZzJ+a1Bv/bUZSx8wYmJQNdHPmEHYmCxioCRtlD8aQF2TvUMlEkgJOVIR7/AZJpMRrsZBh2IjQw9n
SO1oPdhpJ12pXz7m8RmSzhUTJBlt9zcRJXdeoBy3VSI9V6bjN4Fm+7USEUUnOwYg6wfUY5Ayspqa
5HNZzL1/EUn+ZHrBiDBpSCUjNDH4NWHXXAiOD+cFjo9nndEoQlXX0CSTj/D4uRnHQn1L9XssWL3N
1w+nwGGnUv4r6yHLMDdSsv1rgh6NoWraAjTmAWZpiYgfmy2UG+OnIN27Kl+FBlSH41WHGj5vJX8d
ubHIUonU3G8gjAPbxs1aQpr+lHkLhFvP6CQYUVwsjlFBGvs4bvHyNdlwwbDKDvsAnyT5iJDegTWF
hkXl28jGyZNBJD8OLPPYV9owiOmYqpZXAU2aT/bPHKaR/G3emu+imSESyOoIrr4Z60kQVwqiVsNi
Y4UVe6v9GNNb9gOHSwTnMu3apCkEbffSRtAJyl6M5MWMzKsHNUKPNjPT6GlWCJUKllOoLCESSkky
b7mZvjzWpymM3NX3M3oOruDyjWG01FrEieNLeqPJWAesaux8T9i6RR80T9YhZ+31HNrDQabWsY6P
O4jpLoEW52Rr+3TD8hT/xjBHJr/8pcwyCWT1+zmSgdp4JNC0xuwbGz4ev90aqWtmtDOlffKbq5hJ
IIjPuFF3KsK+QeRqXoECWR/qj1oqusFIZ2srSYpJmVlxeFJCk11eBKF6w1r4QBlYPsMstZKeY5a5
SFiMjkqSFvXy5n3fytZXaGp9b/7lQHoAmdRrG1HFyLpx6oxWig4oezFj6eBENcO/NTFDENKI8PCC
NfkMoQ8YWRBCrTWN6V2194l3rVwVQzsUPNCOkFSeyVu/OrKyfwrCfj9riJozHKLs5xgpsnhy16Fg
pd7m+6mFkBB6hGbrk6/sWvtG46WETgsOSdkU9Vb9YdH2UVkd5lldWdonI+trbKFen/xR9kCEYDZC
LD/tjSxJOUTiG00Cv/2LOyrhLmR0UTTM2yWnFdxNPG/bNvcQJj+lgU7x+F3oGsAij1G0sD4qcHUc
9cx6u7tumKkJCOOvZUYOtlWvg7A+nK8DcdAUh5SI19Tl3m972PmRPXeliESkWiHh6D8OXc9CHDdW
33Cc+VC45HuoIDY+1NSYm7CMZcBgGyHza6Om2WY3UkZUZuk7CV641qAOTZL/gRzGomMaYxScIPsf
jPa69GVHXcUit3Kg+0HmAkeElAKXqIXGq4xjcvrggLDrwkDr5zz8gUpVTERK15vgeQ782kF3woF4
xMNyH1MH4hRNviVyjZ5UkOmA7Qb/HKOoP9bYxMf3t6PgRL6ULLoP9kM/P/AHHeonA9rzNr8rEW9W
Nh+zjaDzus2CvlMssUw4P+q30vBNHWHta7fHMhQvTPp10cnFCH3R2LNQ72sK+bwjzYbUvbvcMPy3
XAaC7+8kgkemkLX0T/aaFDOsfVjuq1mBW2Lr9RRbOP91f+VPH7rZ9vf4yXS4ju0LB4Lfl0qBZz0V
kdT1BLRzsv/BJMqLZZT78dK27cgMg/j7eEA+MgWyOafOqQHxlg4YUcSlmnfZrrjC7CxP3T68S/+1
op8TSoUtE+XmOLJkeNhS3A2tdYig6+pw8Z6RE3CCkfkR11Dji0aakviNNnZ+oF+axu82vblo+WGD
h9cxZ4uEamiTOWhfPk9D23mVX1YUDmaXQqE6foiR9DvAku+sCCwCQ4IWB0izMtKFkHQQsDmdo2dv
/4M/P3nnV8qttCP1EK41xkjaQSqiZPvJbtGfnolh53Rh0TrqRDS889NtHjT6cGt+OlEr+RlA3j3U
Ejfsa3t1Y8NV0rfF9fuohca9zxcmVdYjkNCodvRoB9xzOdCTvfP4knE+jMC6YlrNO2Lub8zmZ1yQ
4ulFmzWhDZ8a6sKF83OZsFH8H3/rhaIOotm9CbnyCm1elwOI36PlK3/Ms7QU4Lp7EI5izsv/LZHP
M9q2q/81O2PyUKeedxFE2jDZvGTA+jzRdfaPCNcPk7FpO/DVjbB3KyxB6z843rPTcPhWltddgur9
cBmi46LpWnzehLOyZkEZoj3CFY2SzyaNo5z3dDuK5vgRfpGy3zDQl6+mqsmI1U59m4RUngb/UsEX
TKz2rgwrw7pP5Z1SuXB6qQ8abgHvF/E2mpJpcwrBmeCmIGmOZT44e3Ix36rULYLMgTmMQDGZ9jGn
t5RVs2jPkqPyh0nlC/4NThZ7mtQlt25r80vZqPNQaQeJQrOlTetjXHKzkeLm1d1abh2bZrtxAAZz
oOT67VKOLkljwIZ0BpUxcxSgR7uuxlYAqSraQInVWyv+z6ZtuW1GBFCSCsVnzii/dGB8El9AsOe8
MawOlpVQfsj9UhGsFPOdWw0csaoRo94xzSG/A2c17/Zlxjdb4HMJvDtLvvw8seHZg3bPKGFvQOWc
IZZeUvMQKJqedApUJJetO4KPgBYgn5yjIoTuIJB5g4bVGq1k1epKl3ZTD1qnnGHVuqwPH58MLwqn
l1VV2IjucVJ7JtpQiwc25Xiky17RnnZmTta6TN1p+cuLl3CrX9Dhi5NLnfwLq2ZZzrUdEJvM56lw
3vG0oqUEl4vdPbqPaYvJeMtamhR6qjbWLvehghsj1T0xLxkCVPAcu2u98DeXbgVEdeBX67xe4SIt
Ob5JUlIT/GR788gYLXLrkJMBOBDdEyoBUwADNh+o3DQbt8SuL4Pcmiv7k5ksyCGQO1HNHR7JTiaM
AYRCNjUueg3lfFd2OaxGK8cU4ZHmRksTLJHagXvWhjamToPesu/8pHAYT8AKFFSMX2tyn9IS3aUf
vFrmR5onQ10mf+ZNbLE72XGYOfNb150O5NCHatW+MKG6bK+2AncrvMFiCm1RiqYFiE9xgjPSpUxZ
+/xhZYWah0f3ADmIwnCUmQTqHEUGR79m97y9ScghFoSv1MxOgXaBIT6FCxi9uBB7QYV+uZteJl4G
QZ1Xz2DR3G7HYD8wwIIXnwfQDKCaEXCqbB6hUKdBJFTYu3b6rhwbPCZ16mnPAPKNJxNpPuQahTBQ
OEppuq/eQA1XhzPJlU0RJH5cEnTfEqduYhNjPOXOppSzz7fEjwjd6Bvatjt8T62hZvglHngBsMkI
w/TXIZX1RtJFGxiU7NQuMGcLe3ADU1Bf7xCiIcZeTR/3AhcmbV1jJ3BFdJhy526zHlk+/j5KVbeT
muMuQxeDDwriLi/2+ApSNJ8naikOt0QWYEwAh1pn4iSnVSwEUfeYRsHowzfazdHGSVbyvgoA/MIt
TV63F/a9lxX5ZAITdelX0bGrO6/hz13lGcCd6OVeO8+iOXgB+aUCOLdMBfsgDjdB7oPgBm3WSKio
eelotKrOGkk335lI8mCJkHDqAi8RrqV54YrwrQw1tJMTuAnqlXsAu9kaM/GnBDUrXM7LFFjjDXRN
2MX+0ZMi+jw4T6VJdZPiArzufzsF5eqa7eAjMhpmewoHN98y7ZUq+2ymLyZseEdoUQs+5u7uTbQp
Vbh4zzHcYoHseYa0nI6xIFbXtPen6+q1O8b6swCz+uQroGgjhGWyYXgEXVPiFHNGwvn3rcP9ntu8
bRQ3n8A5qz+GWacHdvXMv0IE29JmQ9slQit/o4+KjDAC7VgvT5MAhmZ4LJq2SAu7iFHSFqorMclm
FUmKwrgPfPKpW6VylzqPSjl8UPNQhXytPyqzOhfhJ79g7bUQGEx3YcMViOk77/bd8Q6JCc95wvFM
u64lqI1SoeTc544PefMsuFR5v7ci/e32SIeT+m717oX5uLQqF5o1b/IOoCNjx4hChU5gE9GUY7lc
iCVCF9PAsHvGExuiLLhDi14HKOyKqZIrWo27x5W/uuNoZ53W1KGkj/JPEgZmHgsqmEU9L2smxGKX
ok+WuFuk+0JFYD1UPw6N+qPIUwNH976vk7e+v3lF2ebXb22qOwVs+t7Tydi8DLwpd7xIbzcVTKBd
X7vRQCKzZd6kmKgLMEPmhjK08vCEIBdbI1KLbpU1C5LQGgZxCs7LPm2RAi70n75L8VVmfc5IUf6q
0HM9WqF/a+NHEV+6fKu7i76ASjI/dHZd4rKhj1VpOA3aSagy/NJROI11wRo/rbUqF6ELwBYYHaFw
ClXm2ZauLhR2Y9VOziZCzjCWc87abKHsPDbO+2a2W/6v3+2RVvcPXaKC1VQBRnzcUwIjrBQTzjPj
8m98y3iMocJaOsfpVlpgN1a0EhU4i0pIXLrqld41ZwyeVko2Tfa+uyTYrUXEL8NfNCDGIlKc0Qc2
RukiDwt6eO9i7/J5tQOZnxDeaQjXHdubyo4ZvkL8y6CAzAJ5YVcP8EbzdEePgf00GrfB8SIgiG+B
de8Ldxj3wgVLn+5OXmAY2sxyd108PK2c4kVmgPqocWQpA9yFEz3rgfUWpUuROwtoOm5oaQAD8ZVD
LppA6jL3mULxH6iLwLup1PC1IErTH/a+upeQbQSqw1ZapxepE9bDULiJeGJK7AvJD5QIid4tXzj+
yiYuA2wYWxw2HkAM/PgKNQaP+RXMCwIkumTTmFHiR3aWyvTeBhd2W7Qld6IPPgHdrhvoc1LZyr5H
EmqXIbmrPyjWWApRbI+AGU/C9m7lsLDoDgl6YZsX9JeCd0kfV6JuPzmb8wv/sPY/Jlg0g/DLfQTH
rm99mTQ0CiMcc38uI3U5t7TxyBnZF/YkkHpunWXjtMIDmA6ijPmAhu/28A64oUlhpa4ExJ7iZOow
3ubR348cQpDxvnZf8KygCz7mclAleHvogsL9FNsepBWaMh6CQvbXkXIh5jocRPlc0FBZJAvHVXOr
hMahbgQqLGSsTt2xwpVbPm3rIJFWajfHH/gd2RuMwrwYZYFimP1AP+5pjCXrxpg8GwE7P3C3ScjC
VsVZldQrX4yp4BHadRD/UrNv5QW3N3n07KKEVDLNOas42jy9CNkvCa/KboxEo/4t2ymGsR8QbacY
Ulr72zM5HXJ7MpMl7RTua9ng9H8yT9ZqSkrvS5cptJmrsYp129NF8jSKPPVDdqkTtfCdWuAM0ao1
ntgdG4l1bNxw+yjpEsPrPgL+bSijYwpTAk3Du2w65qTCkPYDTN8esuEkag0PAIdqw+sjQ+rzAkvS
lZMZqmT81JQCgOOFVkNWCpBDgOOGuZfceYKDORYjPFvhZ2onIYnKNyDPl2MND04H1n/DUhYJPkiR
dDjyqKSh21sLCFMcz3yUU3HA5lTdDSVM4KRlMBH/38an/+Ss7B9+AzXPZ1VTBB6L8GTugp2wyDVW
kkl4Pgel5ZzMOws99Ypw3Dr7XMDnlhHA1sK6azeEkbzPXUA4j96+dsmh/In7vYWXS6Vomism3BRN
gHOPKFhMuzhHczCQ+FOu3+tS/C6W3Gw6L/kil6cwo2OZjvqL/W7itvsK9lvgjEIoTLUUu8ulth43
pTLQqkJCHeL6YjHZeKprm+oTDkrozjXeHNqeBk++XxhqTOnz6XloTAXy7WjbMGGtgATf4nkj1LlG
LuF8UhmyzujdXeDty1iVQmWkZ6jpuyF2va24J2GyDdMqcccCzf05DOsYWiMHV38NZtGuOgwz3KsY
elZSgWixU6BO33JqIMhIGRB0VSBcX72D4XRV2XAGsPS9vkpw2RkWAjpPvuBwnXf/Qs3T2nDjhAFe
JLpIWtZE9TYY+ZyHb3I/7mQeSPD4Ao1xIy98FHpmECd9T5lizndsPmebu4P9bmpz+fFFI/T00na8
knAPEcoDbQf0GQ2FPlCIul6Clx44KPvigvX3QStylWY26FfzkeQkj9DVvF5VIsAPH1w0s3c5anhM
oJ9aDf7jUX+L5jyhBbMAZVIQfgUdI9xoh0vPi51rKLhtlDEmd/SoIBsmYpImdmCc93JGoCw1DTga
HgKfaV1zk3tp+lJtF6WjxvO2pG7MsPwHJFE4w6fgMcLkNtaHJkiZRyC5GMqS/o5ofjsiiygHqynQ
/dGAmKFp6HlCQ7BX42s7GE+xns8Tcqxs8/sMYtj6Ku5dQtxH8C+CLaCD+ODslnkxsUk2I62xpsx+
RJKdOuXB83Q4UH9UBmCFHnENHzes39ve4X4bsY8Mma+TmNt0ShB0zFQb0BIxDeorVjmO6go6GC8D
HjgbnMWp2qHYWOb3A2ykskBJrVps4pw2lQn8YBds8ZP/FI2nKBrmKwFxH8LQfqinMsdfrNYg96VR
NxHfcNtkTo37SgDgmRF8gVS9oyaXAObIbWvuHca6DIj9TIjQA0FOKCifwx7jZQMK4weTj88L1Deb
dJrpKyda54nhEpYdAgGXJl5c+07GZFZ4n+dr88dIKtnJsNV5brPav3pg2nZ8VxAM9G6cpoE70sQA
GrA0m1Uq3A8yJ4LbDHf2+X6xEXQp8cwngfZETfH/Lm5g7nqNmpflrjpZEF/N56BuT1Dxx96qm0j7
rKNrResAwGOr+H4CfN5zYRK3bAU7Y34whXX2UptFMQ/7BYNJ/jXeiwcFO48updb311YOmJe1Ngjq
nMf890XbF/8PE8VtoEknDGBQcmh0BGCiJ+tlwHbzgK1J/GxHUWJm1+imqEmXiaZ0G2GaQJmCVkNa
JuyCZ+IRBPEGcVDSF2/R+aR9Y/FTVy3LLKTFXl5mGVKcc9Qvb5t90ElMYtUrVG9paSFmc/h9mE1i
ftz7eSloOwuTcrGn1r4dcI2FYYpu2kiC5X8G0CNhuXwac6X/AEaAutWt/jgJbKhfooUp4gJPUTG1
7FlTc6dxVYGNKCFOupe8kYcMvx19PSw5z4WcxesAUSRwMSNvUrcxk+1PpwbgqaBYCCX88EdqmOz2
mVSG0HlrjJtf447AhT4hdYL6UNUW5nSEW1R3deknbeIuCL2Rsl35Ha5VWPc9YumQ/AcY1poyfBTq
yqb7zGI1TnvEaZFoGJEM3LCF3J1QTjZiuMerpSNbf4IKYFBxj2YJwP6fr2ckn39U3qlNf5vIOBq5
5N6B6EDa9yQfdLbxi8E6m4c2HORvSXI8hm8wOWIYHcp7qz0+5cM3OKyrJnuFUVqGiwpE2l6uO52W
VSqyLV+NnV2uJhW/i848Ne4t8gSjujVTejnHQrJoJZILYJ/4o4J8J9V02zsXWSBXIEjf3rx0vvdB
bwZPKceJc+ZayIs8OvoYnqNVKCrUgfpELhyL4Np1sdb9ax5hgVUdbHeeJw05sbmYqqheHFI+6YVn
JJ+buixStCR9x+gulsclGHD6wYMfuz1mRchpnBurEhLj+9EbvAeYsrs07Op9wqoHVtY46HhDZ++J
UXgbDBNKPiBnBZomHetGXVRZfvLtR7hO7ErVT3nMx2CGDgYKD9LL7vqfrungHiLYanQgX2PnZYMD
ipoSr5dZSi3Q4VYEgsTrurSdaqavfd42sqJoq9Zwi8ZbovCX4VR4YP2aDHi3fUANdTXI0Jz2ysch
AUk+1lBEl4nZtkvl/5jxQDHznv0cdhcbHv5qvRDF0UQ+2WgABqYkypuKr9yP/93F4gAHhwq0o0zi
LsETL6aEjeFSuczlaxBXdaq7ExM548AyUwmQDXSCh32/8veQkthvjlMWWcluQdgu3hQBEbmIvZ91
o+CP7ArSSQGaGskwleP60ItHgvWytSV5kILDgt8HtfT0DjFcFup+cQ0uEmfCJMFCJcr8NjE30wpB
3pre0XmI/ITPO68OjHEPwtLB9YyaWr0QEmnDRhzPClir/HG0c6jlMnfqm4Nb1tTIKBoUMISN2d22
oyyj2js5WOWTaTq5DEAB+DRiT2dg2CbPdOMyVC16eoiS3RcCITF/AQhNBNkgBthc3hF7Nt3F65G3
H878EN/hW9Vj1w871QWPR1vLvVlh5R9Qpucyt/l6p8xTQ1/R8pHeRuJtXpATtfLcb2fO8BVmEiWf
icEg3HnrwU8WUKMLG7CG9zw1Q55AowZopR0j5VtQu8J/hCLmAbs3jmTvgKURsdt32YmjygBYEr3Z
iMdNciyWLZneJmf0WZsrnlsULS2d7GbrMSIj8yyNBeDHzijhKhxtVXdPYeoyWehLsc23kzXpmuZP
+zCbhRzF0lw6xPn8LNWqwZVk371C+LqgL7C/0e2qU79YcmydjGZsFFYzg+GE8ZMqnEVpF1XGfkge
jLWF1K36r+noDiGsq9kEeg60CEzvBYiuJjdBBpEx6jC8bCpdmQ5RYP/feN8OkxAYewsFn7hgf5HQ
d47iwngJgeyvmYwyEU+scIqSEq+GKMciB3Z7O4/+5DDpNspILW66wxRiHPubukyWLeCn1IcRKt2Z
9PNC1RhP8Up/eouMjdIHtRjQdQ6pd3V+cYZ6dfYXTmlJr42mBKaGGMFxHhmca8txJDsc6uq7QrGn
r5sVuw++cvzBcNhYAklC/AvDUTyCYeOt2aFEw3s/SdbWFWM4Q7Lza1GYOZ5oXhsBLR2C241RtyJ6
ax4fC62LcMpS+BlN3Lzx6bhGJXDYnMN+4ZvnGufqA/rwNOGmrdJGSmgNEQ0Uvy6tiUq1TmfOkzjx
rFrkeIG9l5vkD14fsVVWSN03HghkEDglBL32s05x8MUlZhuWOUbGol+mKFYYbYXm0e+s3GnKwmng
V/l1L0CU34gV3HpfjR2oqfZ7EYMGjmdtyxKWON9zxQequj2L+0PLvWAgXHp0R0A92pTZ5vSDDIGS
9+gj0mgoBRydekm+cmr7MB3Qa0XO4oiUrduW/+VERyaqK3SlNeq6d95BKrASdFvlvmcWKFWb4OSa
L6cqL6yQUnsHb/I/L/rKePGe8vD4Sc8fYT5mm/d0eSHQjv48F1MesgNmHW2RYlLzrHda45Xfa85c
HG26+BCFOwl9JkGzuCTIMZJU7TPMxhTn84ifk+xROqjkjISQCBLI8tBuWMSVCDP5d6VIyeJN7Nvq
msqeA/E2oCkiXge4EkI2NITOduVzeA28h8NJ5+ZgQw+8ZgES+9uQ55NiiziH/CHfUj5GqwWZdNdA
CeGa7dRph8qvCt6CvDo7VHDMFMlhfav++XEwZh5xhfjulwTtW6MLs8m0PW1SgEbVwzklg7bNOCoH
HQpckBMopYgsn+g15MMEABQ4hXYcYf4qXdxUScoGEpWnW5m+hHzMATskJeuDvOfx9/pNpwyM8KY6
uMrmpwkOQU4Sw3xvD4QE+VK66Qm2ppdOpoSfc/qbI5BuVHKPygYC+NxsZb23RHWfoVpaScno2gWd
K9BywP6ER5uY1F6OFgF44emTJPqCSJiPSiB9Y2pD1cecBr5Y8yoKZrZzegllr+/41nYaS/PwGMTg
XomeP8XeMawr9zqj/ozXAeqMm7x5zzJHDyO9i66is2x1AGwOFFsfIK31Rkonmo/tI7IEgn5edUjN
4E8ombDUCgJuEDBKfC9/Pw3RlDMSWNl6qfBXRQ574i7iJYn3/2YQSJwYwHqEvpapYvFnRrxVEqNH
p+Mlz351eTXAKW2sgmi3Cd0i2XeFgFAP4mL7k2NnO/ocy+e4xAHYOCOofcJBoFZuBbjX34YVlic6
bqpvCbikrP/xl8Ykxq1a7PNHP1/Lb9WqvfGdYNIRSO6nDMJA3Mce4BaifIK5yu9WAdzU8gf2i3l5
rSyLBX5gfZA7jkZ8S4oC/Zzdsuzs9F4mRhTCGFRI5WRzzJMdv0LSsyy5RdbK6NLJCclCNYw8GQMD
ThS7LNnmOqre4FEELxMqrodm9vK/v4WXf3nmL7fVSj5CvKQ8jhWj4yeCcXB6kTDQozvepdUNUOO0
dF6kpg8FcoPBjG4Dn1vLPNlWyUctxlBPO3urUFPd5gUybcrHcn933PW3m7SD3AeuBOqEEpEG1616
ftB6GH8ALsKzLeHZ8sdLE92zm6G1/N7IY9/Tl8CmTYzajTULTr2CmaiXIMpUiBphn1VoqRIkoLp3
w5hBYDrsB9Z0j7MTG5sTI/GB7u5LQ9pVif+ZseoUJFJ/AAsx7pmIf3pVgVtRcmq6PaS6rBh/HPlf
CB/no/v1dwxOeBTFv0yzIX35L8kpON6hhSlgT9MHXqbiIndaYP03G1pUTNy3K0gx/bj4ite/4gMT
tP0l6IGFE8BjWgfMJ562ySybEj6DDUJAlIDbDPIxR8gpVVrmaHa1tPio1Slnc25dBFfLWiTQpyTO
uxg7aSZcqnm2fMyXsnAXgxfYMV0eeG8sztG8/shedK50XnKIGCy3lS86H7bIKU7OSj7kDishyq2T
8XF7Kan2bGSNVvZQuEIsjJ9G538IR5/N8vpuLwwV/PPYBGNoJIMkDtRfggdQw3lqCBzeyGtiTrL+
t0fq81TPGsGFBE8zcRrzY93ORU2JshgbRP0+A/Y7Fslxe7xQ3bQNjV6VbWLOfjCE7Z1BqZ81QL2y
POy/j11JnVbDBulauTsYTkoEuM/gUnE05dlzwIX8/rxykRxtW2dFwRwBZOXv8gIFgNdObWtCqdLp
Q9e1Flddr7I0aAP8/bbCjOTSiMvMI8GHD8+g/h7x32SE6YCKgSKf2fVGAdtG9POJAereFJuS2gJx
w4t6fErjguUSSeSJTy2EWzEASX4L+kgLWrgHk2qhMdcX75uYTX3xgnUTGPU5mmjWpfqjQAw3o+5N
FsQ2UK8a3A/Rdx48sl+Kx/cq8alTGl8CJmZn8JClZMvVSUF1wFgAmh+yMDxtFN/sNQ2Dzvq/9K8W
fJSFNlSQKOE+o5FtiZJWSHLANZ4yyu0pkfIXm88x0SwEYlAb049Ea9b39F4nDApON2GKueck92NS
TmsS8pbtM1sXq/Kh5O8lMfk9BPijgjjHixDgoYp6LB0EuRE/4aKfQ5VWir2ZoxR58K2vMC4wpj1O
WEy+ScMyCzfBJ0N74z3JoAJeEGmXF0vbKyDtr26j8/ZDxq+a0SfSxPsdVzYlPYjJ3xylCtaIp3/D
pMaC1r92C5+ZBtNNo6YqUGQLK0ybe7yxbubXzHT90jbe64Unyq5rKqmdOewpjzYs8UKiwkRb6IS0
E2THqE6Z9LtXQMMC1Bt+gyHr88tCkJn6lGjWejWt+zR+PkTJB4/e2HBxN0MT9/iBCHaXaVBcRIZU
wNnXSnDalLWXEdTPWZ1JX9ycq1HZphlJ1b8flGJEERAEiRVVCOYBFwXDh/BNAxU5X9oHxEqk0T9w
JsYcP1/FEX6WQkT0Y1VTzoc/Kz76CL3u2nJxx8vOdjPScxg/zsYfHNnB1jq7QPForHDMdc/01IDZ
6IYVSrFzHDxE7DNaAs48syehiq/C9pXbOAOokNWRMNXjZybTYPEzqOD+fpY1Um7O3mz1saboD1YQ
ELBpwBHJWzkKQvObNr9vZBvTVV47iuoQDx0JI9AYI1Fz7F7umi+jmbhma6qlYB4jsxt/vQ4l0Rok
lShl58MC4WduFL9MlX8gc1sJDeXgZ2bd9l2DNJB448kplgXD+iJOCoRqsVb41T41TqIQPQTSIcGc
FSNA/AZ6Rw7GwrCessJJgLwDzPlIWuZkMv/wkLiy5uGXFWqsS52NhAsbmacTUXGEaLG3bk8Ampjv
VcG2lqwD0kvN3kyhIAEOBUezznJYK91jphKxOrTrSEbDVXjVmVwSK7msI0fuQvDKIHWs6dXjngow
rRRav6uA9c+j3a/1T5egAi97fP0yGNRjjtndiVW8jfQnsSAjIvFEFbZmDBpkr05C4i1zggLqUTHq
BG2A4YJhNIm741JcAHnSicHmf/qlt0EIivlAxjHKZ4k8s1oAFcsuNwRkoHkBJmzyidg5lBkOTK4Q
z7h/+CGL7xBR3Db5aQ0V8Zmm0XCYYL9WrVCVaeAnbZfaLe4U2PdA2uEBEZN4nACt8lHKAPXtATbz
VPlQ16dbyc1WjYN21KV+nXy1KRVRZR+xVHNNWiERMpFSgsRM7gFmyGI2CJlj233Eq39lNrNWD3kn
oA/Jr8xop2LWa2C/gxj4uZM+gtj9d3wiR/nsBRxQkBjL5C9q4xtbwyv5atk790+670/UGnHIe+ug
bjl6uzGHSHJc5ozVT+TJjEGPfC0y6swFs+dmJdWqQRuSAY69vF4KniJH6UHLPOfMhVg9ZPRqMbPm
xJDo9pVnF8KzPIlJHn//ZzwnMM+LxtvDJJYHS3WShDVpGe3GBwYKYXjwZt/OhKCmCbWf+5T4VspM
zS+GRrpXr4VtVy9To5MUWmyPG9Xwa3hnTgy884QBIAEa/wfg4zJ4YgmwstIESMcJ9ZPOeXE2ZgVw
HY4EIM+aaZtaQJ36UsnkNcqLQAWp0+SXI/xFGOuVSHdWTf5dOT/3vitp1jMtHLtX/Dz1hRVxFlON
QzRnU5OKQW3SyxknBszD9nIAFTc9G1synDIrwKiE1yc5/eMYNb9JjsbE8l3yeQ8AVwkS6xVGC6ki
m04A5ib/YEuFS1BMR6+ikqUY4yjOS7a1jC8AKBkBoD+vyKx/ClVBI2F9w/qhSK9qcnzkH9/H2PSY
UT2ohrOSj/qRriUPbaGxBFolBfejpv3Yj037SxPph2EYeqZ9DCvZ/Fnef6gFXDVIl5t6MFOh8+qU
HyzVKm76pWI0BX/JXM0YKwYh+rc8hl8mQ/G49xgRjeaqu/3Fs0AKWasegt2DCOY9uj/drc9NJyvC
jGkhagyaOIB3TvZwvHFlqIcjfzBtiWXgSIIKQT0q33C9cuwS92RCkdQ3f1QK48ydNwYB7wDEvZnO
gyZ+ohcD3gGbDBqZPqU4XWxNghgP5wrZdlUji0Ztt8O4QS6Zm8xnZRy7syvpC+NooArGuzrIJghl
9UkJWCKRFjvCB7bsk6m/o+93QawcOHtYiJV3xDQWVHkN2f4Y7s3mJUSSY1VsH/+jV5/pYosbihkY
1rTcrTsqM9ToHVjZ8CWM3o/f5O74+lLzaF1+0A0C/Ju7jfB3dZzJXrIMS2HQ7oUvtQUipnppJzWI
aB9v+NbF7AEPjPuJRPEbqTrwB0k1iFhsBtM/nyS2qTgH+sbzWHNP2jbJ7YeLBILNHzYe5wLB/8CV
En/OufyuAkgbCaS9a8gOcx5GTtFPJciKYAJiDJbdn9psiNrVzHh6bnCnhzblUpI9oMB7QK1qgWps
RCa/iNdZrbPbKNFmbxOai3gFQLzCu8DOq7FYP5NxWwIEZ6mvWgR+A5HlgnPDQEMZ3bs0NK6MjCVS
4wMeQrpfujJWCJO5cjwhWxAUpr8rS/S2MHd4KvMQn5ktjwrWiXYyNfP3PgZZORCU4yTMy9++iFnY
B73FBanxCdRDHJPo9YOThDhtUPi+K3jJg4Ly+tCfg4O/rr7kj7DdiBCl04PquAOrmXgCyve7MpEt
gwjV7Wax3E4HllXhcbs/Zkeke//twkiVTzCAR+JhF0USHatjAapz2cK8BgvL8SaF2b9K6ze2rFob
mJKmd5S1njbCVLka6RCxw395AilJk6GcGmR6xWs+QLSChw1KBZIdBj4ee4K7qG73VFdbP/1Ulq1/
B4w3v3XtKvhIHNV2/TxkMylvDVx0u9jpQCLn5WHu8068jhGzq3OjnysgPFqjjbMlyl2zmqWv8ZPt
62iKnNOW4FVjYLGqX63zNCI++kqJy1eJWCgshUqo8Bn3hO2g2hTnXiJHyLJLYfepx16LZ7mC0Wtn
DfmhQUDqd56uLGSrDkjdpzSAHxiq+/PENSydZxgTYp5p0QQg7PRiPjVCqCx9bI+QDPA0V7yM2AJG
qYAnRdLWSYMColgct726242KHeraZRhPTWpHJNj/uRzLWtOEnDq+M7TLHna+foa4X1ZvoRurrwiV
+CnuRhXorzvdi/zuH/1WXZPu2mYIzgJPLBaloWOhiw2hGzKAYGrH5RzFm2C6TkwFzDq6cha6aFii
pyP68Fwk9H4KcQzs86CdB07mGNIqCbFwax6vs9hTpPGWc4pjoD5cRceFF5yED9tu66YATa/cQBmg
SGfa3o48+d9dS4Z6pHR49OpRGs7tYzkDxuuinVlW5rTAWmdjGtvXxDdkI2IEPu0YE5J+XWRGM7j8
3/dYVeuzD5MDFfBn1J8dPr6Xp0YHYG0p29A/mFqcfNopFeCl1DI7RrnFruS5shCFHUUlUaa85UZP
vLjvgQQxJkHgwunqbbOnn2B0d1jRzZ1vn7T6kMia2JvyhsasrYKWIs5tKJ2pus4jlrOF+HILxe5v
HW8Wvx0RRwKynTiCFEzSLkOTed2st7Kgj4G0nBJ+j6u9AbcUNQE5fR+eQ+i0fziYxHbUfaxutpyt
lpL9C4a/nRAoyOLt6G8/l3om6eWC0YTQyKrMwIweGYpISV/pt3oTAoRoTb1gluSnPD/D2Rb3cmQY
Ym17/LcQeo6YYPwbDmX8e6ercvceS5r5lfYIKyNL8S4+bLwRRHj8Ysye2tyUFzxYcsSgHIT7027Z
FNAXcJDuQ7B3SBcGcuaBcoY9Jm8SH0+L4Nf5FPH9uIJ4Z/RQRDA64hu7hu3tArHOLjlVnWImeoO+
6lgXCdBerBIKO0373lSKgNikV37hDh05W2tyrvrmiHKxiw0A4TZRCUnDTutO2DMmMdUiCxu3iClM
QLNnaNZvUfEBQwqJ+4DsFPjJ+GbJhfcz3MyyN57Ac5ItF81OIcINU9H4tRb+XUCm6yiKsth7jMTW
OZMu+75iMyx6Oy5of+t0QgpNrKy+b7pNsMU4BXcaWTZFWv2ExxcyLmO1xGa0PI/L3Q/P0kas1ZvL
moxEmrsKzRt+QzXxb7uVZmcYX5QAve87foi2hHzv1WMOLOTHwlCJTYxvlp5YmHvFrTUoFuGf8rpt
Ac6pR+tArbAEtOccBy+BlSevY3dfSnxetKu/M77uGuStiF7I7Rfy5riGbaJxBcqmW64agCTBOpxf
CcPMdN3c6+e9OVLgUD8t4O2rvGnvGgXccao3E1XXh1gTTlMUBqnBeVpOgOpE7Lie9TMOBTZ1rbyn
8Ha/ccyxJW5w310Mx13fykUZYOEqe80Y6n2DmwKHNyfg8urxLkayHX7xqNOBLlZw0H9J3/k7rbwl
TKFxDWVzgCBqRxcHT5Z1vv6VJTDpIr3RwY1Uw5ZAnol8J1bvUaIYhT6WX1xDzbhed7bDX74FM1Z3
qNHvjoyg0DDdMwlxFW9jTDR8JAq3tGpcNzNzyn/h9zMHtJJJqeLOVrjkf9wSY5dwXM2woPiRoEh4
1iNe+vrWG/26xEhtNxT9NFen0SwGvJ9r6pBqdBWBRCFkYGz5KFsIe4mJHZZD3HHtMv7icSfEHPYL
fMwmW8LwVYHnJarPploaKVBlRIASgapKDOuE7RnZZ7SvSOmlBgDnL5yFjhBUB88cZ578P0p+eTyW
XLUDZFUx2gU/03GW7huiW0MpbAo3Nw4OlD01MdrLq19IEIuR8vQVuv+LN+P8oLEB7hD5bgeqAeXm
uAPGzWHA6rkOVelVmrmDG+PZk3zYQzMKe62EZm3RkRoLyUUFRkcUnoFzskibhFvRUHKsmplzSLrW
48PO6Z3nUtmypTXCk2Ln6zewGQxmaMSXIOkKMW2n4kCJRteazoVQIOKj+euxXH662Qc8dFaS4Yc1
nhReK+pDEgUqBfAEi+tkaJDT4XyF2WHwOEw/lXrGM3QXK2kWE5giaRiyljWmbeKHrQCQCr/2p0kj
eqiQs8iw8sISi0EMAO8kJRVaBm86oru5xadk2V4ZwSu8FS7YoqcVxEPmIhZdafAk94HBlzTO4c7E
JMraD+6GvHGp6d1DCRPxGDFwA+5396lsHzbfmv+OxmD1A5lqY8UDQAHw0qamk4Pu5cR8fNREL5cw
GbAWgZg+6D8iiQKRznjc32kEFjL587ShhF9PjB5ZcoIaliDatP32FAQazREnepLXHyjj4/Q+BLe0
K3ZzoEscXCDr9W7bw6kzbjSsNlHtu4QSMPC2qkB01NlNQr1zIUqY3WTzqeWFHEn4aSlCaQBSzyFW
BIHrl1+XKCWhtBGqivQUvqXuchD/NPcYidHUyg+8cclQ3TyjMlhH6E5Kwzya4p5c9cvvAPPxSP32
bcz36zaJatLa9/A5Hxtl0E1CpphW4fssug/9FPqrdbTGteCyRBkWJ53CFhLyET8c6upvN5uvl4ZC
3b5kcRlCJTKyfLLFw5P39A/VHlPkiz6LWjgiPdFMAE9W360ccrmtNkDAyjKdaY6kryfBHSgWUDFx
j0wQmZqxvuWehZBHSToNByfY2BNMjV/ymPN1nloqyjVsTReVAxaI8V4FC567gp50Op3igwxiJ8HO
6O9QPo7RLqXRoICdNZd/lWMzc9fvQ1lZHnE6MvveC9O2uWifCBJkqUpFpKicmx9EoJL5DDiutwmN
ydW7tgOa/dpcPiFe20lWHXeY2KSLkMZxKIDvI00MJP5m8EUlqYh06AaTn2+CZk1wZW3tWExJhw3k
LzVkbc6oeNNTOpfaih7jl50+ewb5BXXj5CPeCPIm1JWxTXYml3rmJ2gXzXwD+WOUXVFqQsXn+YR6
Bx+JNSd4IjaMkjbMqM5PcaqWPO8V8gTBAju8JJY1UZnz488zfkVosPIi3Q3vh7Xvd4dFccAakgpU
jrgTzB0KcjiqeK/MU9OKnxKMaIxgsHkdF5P4EcbuelX0eSQGhMn7kF7acA2vNVdBcxE/poWPU3LN
d/Idrb4sPaU/xZnU3o7ToUkCCn5VzkQaktFpV7h9q2XI6VQ6vY9VmfQ/Xz4APgE4DK0gtIAl7B6g
MqqW1yL0FC+z/HBku3mjxi3mpdFmU9ByLO3/IGpjwJVdxD6G7mGTx6drmnvSLOEbS4Pcfco/7vlM
wOxZUoY7i9EMwT00ckbfk2IoYIDRUBFmevHqa3RIyxNVzUmT0F1Na6CeplAP0iprjit5rqbeHegg
0OCznW485Lc94m4VudC3bZ4EF54KjPrR6w1mtZIUPBlc3P1NYPjlGoajPz665MaJ8BFqGlCbHRir
WqeXQwVpae2zjPPtcn1YmIklnEWSfsU3CAWNq6Nhrf6Qx6eT4z3ifnq4A73v2jYmiTcqz9W4cTS+
6jC05XCZ7PfLbdMM3q5K8TavvqgERsT36NyPH2N3ANbi7F29qpdnbfGd/ZMYGDdzpaxslFp0dSPU
161dSTTWo2Q8RNjoI3y+aaBbj62eg6lV8zOFUZCKjpqSgKuBfUicZpcE8Jw2guIuzTHpPsX6Y+VW
oeqI0XH4vafsJ7lDVorrgMLQm4WmfTgl87wdQ7+jRkGnLUGp7hrKrRWpRXx5jkJOAUYdyGuARdC3
2n3H7c8NDVR50k3Uj0Hg9qwmH4evNeKf0fbanfnb7d0Nzhfbgzx4beWmecTzvm3nR5FsdLAFsRyd
UG+FVcXYadUOfcXx6yB3OKoVx+pYcRS7z03ZzP7aZ8k+dhI7mLLr47T0KkPxjAKUeJM3M9JXMtiZ
2FQj83FjvUby+6Rad+xb5OW2KBe5C+6w8WEegUIjyjdtngmlOk8V35xF2IBgRw2cDsORohhswNTj
zslSjsG0rLCKc7YmteAzIwurbEZfn1RNwmb0m73cZvrSctY+rEaBWAswVmDkdz2yUyO5/L6UI+Yf
EsZ8AXd4I8zEUyKqLluEIbslbM6QD6QBhKuE9EljcJ6NAHB5Nurueu5i1TxI/Cv1oXCwAzzu22yd
e3JMIXs0/0KCD8eDnwuGijbVKJ1BzoKNYnvkjivDVvO+8BqBG0sJN7+hDuA+VTLyN8WDpEMAYu+Y
gux+bvDSUhiriAPGzfj4fzHZrS6nR0WZR5b/6Fkop0VID7exBmz+ghBwgBBll9njjHacb1HCvRCf
gFpopEBGMoqTJiK3yL4DgTjUbK0b/bG0I9WvNcMWc7pYCmc3NvDFiWt42BioYe6AVFwc56qoIadV
h6D3574gclCnbA2LwHL7bEQEGYCCiHegi+yHsPIsVy4Uj0uxAhHKmKnNk/qAe30ztUXwsf+loO5m
gAT+mRotgNsLK7ojXyGWtZi4tTKMIFGMPi5I8ytnQ4S24Ir2fj3petOyrZjEisyftQW8wLt1GINT
nwCdaPWpodYBLufEQLClVpLjT62Ph3lli1/4Tu4/yeq+vg2HBZYv9Xbz4Xx8nlO6UN9HP1IXqUE2
qaG3ezD1px+7ztaVcl/n52iCXEhC1zGzdtIxhccfWZwyPHBHcuTxSDpbdY7Ih73CpFy8PaYTrwuN
ksQeCx6WkRlkE8QJ9xiFwttii2KHUP3/9fHCkzqUdGN6bDHIlBD0p8Zw9Twmn5oDCr2sbTf4/aCE
80QEUBp4oY1N8xB0aeyz8oMiunCwYxHRIddmYEiulyXNlZZ9sJXXXZLMmixn7tQ9DS4e5Azz6DWZ
nPErcgJL7drDy1nH6/LC05wwrZVa9fmB4Qa/uXmDfbIzzKcmjU/0vjrHNfPWVpn3JpisELZq3yFq
BMNEzONPxNect+OS9UH6FINM/ZPDBGV0LafMrttHIWfPdsXl4gH53FbtN0qu5r6rUl33c8frm1/h
kLaX7JYkmHrM5KsODx7EDFHNKpZzKXWLf/0N3WZ/dsR73Ou3LFDlnQye7gB4qK8apeQ36/Ex5TVy
G6nk94OBkspD3+nQalVN9wa9tY5jfa5Daqn8Y94orF10nj+Fvd8R2tixOmyY4zXsUmcyZjbsEp2h
l5p3clH859fBvQpj8apEk9e7A4ybCMFS6qBK0ePZmApuo0wwHlBifYdMX7aTE844D+VYwiQkNTeh
ofxycFLi31dkWV5uzzq0V3Jrou9RcXuM3q0XlzwCwvuUu+SJ4Ksc90C8R5/J9ODiabe9iPNK+Vht
P5Cv0JT9vuyBv3pZi38h3GOAWNBUDsiC3WOXdK9LUgp8VF9mTTK7ZCFu3G3rn42WYsQKC/BAR2OB
9k0MXOwpzMLtiGtO0TxM+61mNh11fWj9AgW3XrO2MH6SVFQTsfzwLwpFdqmg8WCZtnj2C+bc3YfV
7t1UQnCK6siNoM5bYPnoHOtoQJHdEM0G044cS997E5cmVODbn9goeUrp2hfnGuYjmLXu3gPwSljF
03UH3UlG0G8LrOR6NMsA+Zv8ZtKGA61pX3SWQ29t55QtiZSzEodMqz5TJc+WTMOIHXJGLl5mis0M
50cZ06dyTy/BPNcI02biZj/uRQS1z0ZfrJNDeFv16lxFcRRE7cieqM2ML3zW2TsbGoyWBvXTVMkk
YdhQ1IC81INoqdf+4oKAWdEeTooeWUaMCDXDNJagLNesN7P/RIYT+d3x1Yp7hGv0CslacckWg/DA
gUs/iGiu49tC91taqyHTt2BgLdXyQP53bPnbb0i6J6VDeiaOPsVGYQYzt/3uln0RP7kQKDtMJL6x
lp8wz7P3VsC9AVNrPYETMQhiAUaL3BuRemfOcGwk5/zTKrRIVO9tnLxqTDepfmyvJ5RVRooCTWDx
0JPjcjw2iJN2DXSAThImt2dypfB/Iu6/+fqkTMsfv2riLLEWC4+UFE+8smnQkJ9ayQRmR9QhCF31
58d0uO6cXpjgj1X4z+njXkie521k3uhn9UV6UUgSoolSAE/YRam8L9XQ49Y6hArVL1hRTjSIbBXr
tJq+w9bxyMqlpxTmKVAd9xOYYHl5JEPW4mkTkKh7mxbrkpGyK7KNUCDgPxM1clLSXnIimD2KmVSA
LZowkB4ZoSquvuK0utYm3UsQ1f0aDnaglrPp2QbxL+fU/an7DZMJUshXoez1h4oiBPxJ11Fx/tyb
ATDqx4QE1JwG0QX2h5yMOOOpqptLjCGsuJ814CMRSWI/pABv80MPze2KDZ+PjPiVHv7lXxwHH5I1
gfLlcJVPuO7ul4FKZVbjXOWKF4+Lhcta5WmKdY/OY9EAeAxWy/L4SkhWd0Ew5hvmX35vgrRcwPYW
4cWjnYcID696COqgU+jEZC4koR4xNtND8E3HYthvatljk7kttzfVHxCg6Ky8YqOEEs58tcsZ9sBs
CnxzainI5FITZMfL7nKLnXiFEEu5tlfs2DU+MaU9UjaVYJ3rO/8qmdoubt7DK9KvPvzOvAaVO6cf
qsnub9pkltqaKcHoz0lREETND+yB7ip0SCqefBHXSDMLphE0rWpttB8bTLnHy/SaUrFrn9KYd+yb
Uh5G7BeSUx7XoOJcnRNVMI+z9Wn18U2jk8fg0uBX1I+n11eZEmYcSBP7a6F82oIPHGuBZXH2SzsB
Yslbda01aFtQiXhxP9FxTN3TvCTyrFhoJGycbumz/1C0lC+JmjGjEuFkrU7RdliBCYMM2fLGGJNh
yxMURDTjWalbQa0crF0nVOddpOSV3ja679pXkz7uxm+yHGK79nV+NvlnirnezSkCMt6BSvuAr/wY
GrzWHVugJTh/axiulfbPUxjQBdlsMXzyHl3ko9BbnemFLuj8FHfR4n5+sbA4SWqwZvU1Ti90wTux
pUobnzgoO06YHE34lLUc/vuFdXSP9npjbAwKOjcy4agtcxMS/oQVsWMmPx20WhHrahP0GPGhIq5U
mynszytCfUMOYK+zqEzWoWWhW3vEeRDB0yGb1otUJoyrow4orjLsxsQNTKjh1X0cpF42+i3SRIOU
ww8RnVrGFbJJ4i13kguU1u3JvByQfiXLAo+U/wZrjLlwVHZ+FWgsrua1alwj/uJqn2RNOs62u+LY
+T+KAL6z8dTOCfKlMQl/e21jTiJSEad4XSQPfLds/tFdMJ+boSpJs4QrCBVHs6xJfYnPiSHrdMmt
ElP9MGWT0hbpz9HeZS0vUQJfyt/KdImCurFaaGgfJKwL3GMSa+pW6ias29bi7AuBsi//g9p+A/uE
0SCIp6QpmWcQp7q5ECIoE+a46Isij7ltofftIMtDmhRK36GX2GstH7TE2QBhnq9cOlnEthi8n4gq
H+JPohQjStLXUIZdBKL0/vnQn42hzRG4tHWFek6xVtqjGUYw6N7SzVrSNGKYnQsDq2Fl36r8tnsj
UEtbcQjq7iVZOyTVPO8SAXg4yLz7QsZ8vGuU5ABLBdRzA67hGnI9hrnzlGEcekdyYz37Nq1v6XIm
BchTbaOoRv1rw3pVQmz5qBPHOccL9Mb3DBSUHz9sJlNiBC+eQ+nmi58BgE55TbYzWwDd6y6rWsDp
gKbV6hvaOn3flHKzGz5QfrFzZOC1q5JjLW2RvXCVNS9WuBhXHRIioVQTkE0ZAL0EUi/8MrDke8Ke
MfwF1lLYNV/Rz1KXOIQyWBEO/UplxEk5Z4+gF4y1EnIQm6OlADDsWc8fH36ofKguOVrye2qxVCqy
y6WHSwHgQgbcX7TfavfUPfC6HBw0xvyzeTVGsQQi0hrfRPwRkH+F0HplXWyo9n6gLNmUqj/E2D04
jKoOavyi6Q89FhBnuhb0rITRpQaLm+MO9ipcb5FbF7iyb3YS70D5zR2EC4W60PDvxSt4WeFq58vf
GKRTlEmpymILxlyM7y6RPGbiEMuIO9+M/rn9S3CoZdeqWXblP/jmm/2dm846euHV3vo9nOrOSjl/
Xo6Ls2AhgzR71wPjwmviRJe+IQGlk2q4CoUosn6QWSMG0GcQDpOig+dmlNw4uP5ajw2P1hqhT/PF
nmcloxvFM1SvvpsqVW4I1V3B9W4GUzHvkv7ACoXOxG2sJjCFEtJiTmCk9VQD2kVeH48KfLiddvUF
UBWHnLmJWJySlpPgLrpNPEBMWHESYn8mPlcuNWFP8A3QButI09YOwd69C/+3khNY0FOfJwDRjaoL
eyvF1DXdbah+SIHnqPA3wGjsfl6AbSgeLDsWKpaVIIqnMstCUIE2uFqa/NG+/GNDJRaCfqyOK59l
TZKppPI7p5ZNbZkpK5fPbh3Ec2i/ececuy2UyQZvsaMeidxFRpzR+FdiGdGCVYaJmVDi8Lcd5H3P
OnVgGjK/8StaD1VlnoXrGHnn1kZefPlQnArxnYNUX2FTqS++fiBPtXrpNlZgJ8/aGbiZZZRyAHkO
OfuFpLI/r1Uio5hQV0fKsGnJpQ/J0J4TkQTzKGT6TkboElSCnH5ICLg/oLpR5aZobanmHL5pqb+H
8CqgnLlyfFRq/2WNALf592yaOUsDbkTbSmTudEQinVfdOZRsR2PDJIsUsbvvrjz/9ARGsVNz81I2
6rsTJ3BydlLv4hGthoR01W67apq//5apGS85fh9DNqiXn15R8qRef6DZ39TCPMJBVMQwAhRnWNtV
7xEyLx7wtt8MbYLgac9FCJjV52ZF9I5LmL6EVIFyxYyojNY1G1vXRSX29Zk4d/H+aIcDOIHgBRGj
VUHZOjAOMbouPy41fGY+zXJjK0B2MkIVe5Cwz3CmC7xnSzoQKyWDFYaKXnEgwmFuLB1VfSwysm6y
TirRShBOn5XCHM+XnEq02yDpcxzBtpqPV7HP97q0yTfES3Z24jmFmfkxzICT7OE/fPyL2wK1Ny/M
DLAkbSISTjmL82CaVLSJsso7IgU7rB78h3OYvhq/thKu/bXHKe02PgSRCD4bnQIw9255UyNvJzF/
2e2DLBvmNPlH4tiIZTh+Rroq9Uuf4mnaVNKuJbS3p53JFQrjPFiL7lUyKwQJqqLw4IIGgE1k8IZY
g6OaB6+Ru5/fniUiMuJtoB3O877TaTOB7aAuwEpenO7I/nQYdtPXWlpwjtQlYJurDnKqvJHH1qyy
20X/3EcFnd7++NDyspiiQAJKXaVzDcw5b3N6uk8OkVW4R8MIW6w7gyDqiiVjMiviWG730Vk6GoUS
3R1zvVANg0epgiG7KegLu0cXRxF5jgSEZCOfol6hyKiQ38AZc/3kO+i6FI4mmISrDV5wUOSkrxkD
65f25Uncrxac73wNc2WYJokkkmQIFIczZaBEJdLoVUglX7FBLSrIM2w2FMiwAEdTtZ0iXabNYI/X
45d0KXXLFFkOc+0mXkxvdBPElV9BJi74E78lFkpFAuhuiz+wRxHUo0+etk0CyEHeKtqmpwpn4ViX
sdzLPulNb+knIUFfvljlSASOuj/BddGP7dWHkhx4K3TG18o/m7Bu/dCLy+HOB/q/D0qDvYAtzEAd
Ej/k3AnaeqoZhuI52LsT+gHijqeQI3ezCp5TaD/UxOrueDfCJjmd8syKAKKiPTcF0wnNuf4LwNEC
TKfbEJgkdmniAY6m9VyvL0RamaRBeQJG7QFOWBdcZaVzpedlc4IcrwVfUISkJXL9BAB36Y/Angor
AoJ8nIIbcRQAegHrVtaovfOYs53CXMFW2l2sRjWDlYb6zOMWOWa5bDs04pzWv1ASRiPtEsW+Bbl6
HEOrPUk0bJhbk6CRudYzqeB/m4QADmWufTj+Qkpy39cCJEwlyQfV8azaK34rFGIxAbNDiLYOk/M9
WQDN28Syh6vPRUn3NzDPP8kFLL03eC4GSIkkzfP02G3uDhb40udn1ufNYm1rT8ywJrZe1eAlyWE+
ouGR/EL0syFLFVOIvjQHuaA2MdoJHZmUNn2+YuhAiOUzA2Qkx1S9J1jtFgS1NUM/ZuzZWC0pe/Nn
AOxXeC22h+xhTXUqLWLksu+eYmX/T1Oh6kU4sXQReGNqMJYjyTAI3KQM0tV/YRyt8x0/8HiuKrzP
5A2KHNUGq60uIVn8h3lYLuyeU0WU4Kw9R0q3HkFYHpl7pkHEXBhQEnnYigdGj8z3aSefivcYK87+
hifQUXinxpzYLCHk01Ds+ooYp758s2pyE01Lf0O82zFZVn3LYVAU1IEO+fFCbX54RM10qKmP/L+H
u1hWlHg8ldnTl+hnMx2lD1uM677QK+Y4yJd23vqu7auflnBkdZLRohYU7STxcNuFqV3ETsFLOogj
gdzDpLrQksMtVAAbu0lJeOfTV7Ci8mlgWIsidleoJbnHoLPopnCriwQWw1vA+XqBrZgX/7ukoSVy
1yl+KGJ8iGQHxxdaYMPi0qR1kr9/w1/2yD+3sAvRFuD8HpHdg3MCS9/laqkFnLtQrygyWVxcTdo9
W2MUGjV+W2SU4UgDeYXYlMS1Ueh3dkxI6UHM31rTWJzD/OcuGCfIx67u3uweF4s6eSTl7AK68Sd8
XfLzm+cdJBLxKfHdiXctadCTIL3gBRCq++LsSYBBOtLl5pVhjDJw1LRXD/jxlXpgar71j3A03mdB
HvTukVF7va4HfSZHOwY1qU9mRto+EiQ0mtJg5NamWaycapNEnPDlJgLhHjV4QhlqW1I4D2HQzBqu
RddufOrnxYxdBeUQLtjVfWs0heMVsW6z2MhyV+y3AHJZlPyewhJ4QcK1sFofS6UitVQfQLK62RvF
SsfokmrbBvT35Ao4IgMMy9sa334nUb0ki6HkRuMaGG55BH8g7XQDcr0df88E+1LOfPn72Qj6kg3A
zHIqKdP5BbKgVZnDNNgTRwF4Xf3K01If/4OgEd0sUJ6vPYD2QE4GrzewTfWPy7Da3nW0V7pqUMV5
LnUsioekYAqxtP9A0jGIffelxLRD4ny/Kd7l0Ve0EMADOfsCa1QXxvBSv82qsrJFHGizCNjlk/yM
FsnId2Ya+Dt33NnMHt8QLr0KjWDRt2nZKbfxUQgp3A59+ZX1Wg08fo1TCafpD8tykKMi9xqP2wbK
K+w7LSt9p/8Pkyn2ItLSRfuJ8PxxPa4KGIjMmr6qLYhUFWb4QzgQ/2Xnq06qacHVsdlkuUF6/tnU
y1tCLgkLD+g522KbEyep93Z6aZ8SbETfcCn0Rq9StO1iLK1Du4xcomFcqnJ14je28wJeCgx/4hgY
m4lef6SI/wleF4nQUHcqAAXQNlMOdyiU2PNR2RSPF6Yo2sNPK/ULCyk0y1LvTV6XVMzHqu87PBY8
Zi9VQRBGQMw/yMz94lVz+FoJHEPnCAYleiDJHF2PAeUMP3AwyUMPl3e0OyyqzFDmLK8sYh+RPu7B
hcD7qffnBb6WDnBhyJXSuMGutJlrTt4vROK5tVFCWYsTKr5hpfqsnecfVp7Zxo1VQfDPX100Kopk
fbXoMz8YaxJ6cyznqbTcVdrxgA32OmCghqvLTRK+5Qi1VGua7qgQpQtfROvW6TBwuP33EiTpyLzL
OhQMolorn/BLGgzkZubHOaGboQZDIB9eDY33wWfw/1wPd5r+Fb05YAxepX0t1D/5XaifOBV+rM00
yiM2n0y0mpuT47PZG0ttoJ5VAWvq+v2Y/2uDpSIU54uOq79McK516kDxFTmMQUtHa/othc+H8Dgr
sphZyn2+DJggV1aUDbx+hj4TZRb/JuxrqjIeun+f9lNsQqU7HY8IBs1wKd4glLURhcjESA6XELhL
B4LTPp1CY8x0p9L/3SgM9gbbYbesX30kiHcHcdUTxdbpci44kf8yMhfgMVruVSSvhb7UD2fvT52n
Pb/dlCu+cKMt+kiV7tzvhRxbDcRiqvJEUcFQzxjbLaM0xLCN+PR+a2fcM5v7i53v1eTRNINSYnfG
iCQRdErsy3+6HEfu6kVwYXFo5JWcSXa+E41aR0VQtKIOoXASJ6KePlypGpC/ZSraembehumHYokZ
qpoeCffjYh8ryDTIuDcllMHREr4f/evoEtxpJ9hlY0mE0DtS3/i1jz7ELA+Huv114XB0jb1cO0jf
F+cvIJmeNUHZl4F+MiMJ7AUCRN178m7WU2L990eHZp5immLfkJfJ9cpJZuzfLPBbMsrA8oFMPyro
0T97HVs25NWGyfj9wHB5XISBy+7ewB5oDDUS5dyfNT8524V86BMmR8yvlAjTitCh7RFANx1zFLvN
CxIcMeDmepZwyq4ZkLGoTcGXBPJ8+i6PBfPH8GTWLOuG7nAQsFHIn9YY1xrQlubBc400j/pTacw8
vEu0lXRTwgOCL9jcF0lQcFt4P/DSoOgKWlOS9QCGmgfns7kFz1XhpU5FzMY2syaV9SMfaIfzdQLL
1rlVJ/DDp+urseM5/EpQJytsGq2M94OxO6qEKusf5xcIy624Xcg+A+w0/5Ks41EQfdSOgZveJaZr
kSc7723stBXKnvZEXKlN0ZDmKivS0o503G63pTTSUjBxqXdHLrQAT0NRj78+/K8Q6rLI+Nep8A/Y
wxAL9hmWx97gUn7iNggwNWLn3Gm4kFd9sn38wHrUjx/6tFfnAn64TWCeKFw5E83jTb+NvWrTBBau
oml7P/eU0i0UDT9GGRL+nS2aGigmu6BOpbUo/Cf9h0N0AlQopBDa6K/OeYIWoYos87WjcNEjeRM4
a57vvgRbrkupvoDgxE+virPE9xfG24Hj0fIG6O9Z8JWFYvwn6H9U4XG+vK390rMnHLZS8zMNGQ7u
Qr0+Uvmc2T9wXjr17sx9WwSF+IWfaQcdZDz6t5VQFh/W0aR50ma1luqvQwVhKVGZTka+wKXxBqrb
UlQNcFho+a+0/QgZ55wwDmS7HUyzJjqDH2+keTBLCyrzKViIuCyfjepvClbX6aZsrmkoAp5a86N/
xkMyjMkC7qqa4MhPLnnT8vls3/WSiMbYfRmRNkC+CpOi4XAKyY5ZodU4ivL/cUuTVgerc6iE0FFp
rD6jbaXvTCgNLXEvRdtmti2q5rTS13+ClKzT2WqWQS5kR17NTCykWlCRdddCoHj+K7TVFWS1c5FI
vzUizK5v7OJUPpm9fuvFOL8MUTMa/WCsOZTp5PYenSexjHEEAxvE2ASKLvRERkf5I0MDrilzb/LR
w64tp0gEhQGfz61Kk5eQNzhkioa5Zs1bVuFTS9LbdeacZDqYQNOvqoN+8EkgO+lAqPkuBsAeUBLm
nrMOjig6oDWPEjlAZgqrFEv43tuWvjK4fOLKGjFMqi0HeTCrI6Uqtw5fH9fPhwVo6a+gi61w0ukD
9aCrrJdpRxMl5ZnmqW/XbnJI4b6FKJiSXR9kJecAfaBtyPGWd4PrNSKp6fpbp5jxcgQxOEy0apkc
YNy7ZDCHZxX5CP7HByEnjBeLQUsVOMGh3pOEQEP1jECLWKXBczSx0zr3NqAB0NM/EygwaLouLR4N
Zzj4beB671ONZ/xWQQsKwTMjleYhrxVwu5P0eAJqWw5ES4L6a/NDifYCf4Qc5QihlMhnQOlHz1Ah
/xz1HKZpej7oaWGuD50/8LbUJwdXpB13jx7SWE8QG1/ZM9mRWmlndIjaRl1ofPxR3IShRFj/aJtR
jhjlQ58YEwm/ateYblr2YWUB3TBFusFfVmlVPmnMfENexUWisb0/jIbeg+FP8VI/Vc88V9Xozmho
8KZVgNXP8e6GfiGeJJGnul4QzfGpIDKXoSm2JrME2mbdOo7L75G1oYO3f6Q/BAx5ZjnG6YFWTGKA
yeES/W6bO9H5IFLngM+RUzApqmVRyWsSJvbxuia1tblfF3M9m4KqoNjSWba3YPIQT7UNmJcqsyLM
UO8E9WPDhCJa86sME/Gu+2MdifSNZL5x0MMc8iMRTtqvXbnOtm50NHLgqrhsDrwMMZyZF9xB/FVG
b/rrl4veZXFwMe5ZIMowHi/+RgMvsUrCScIeWm7s1MRlsDujaPThJcst+ne3C7eR4wLGOgqJ62av
7ApcTemkxhYSrpAKIAmi5boL4B1c2YiCYIWR7iz8U4spPb/KZu1RXgc1kVnp8Xg1Ax2vVXwPtebC
chphbjO61mRXYPpcXUbc1y7dt80FR2jHzwly5/RI3KY3kWI7WVtAkh53NDO5nX1pmkNpksIhDN8Y
2378oWwMd9YdkWdkMf7bjOim79h+3sfSI00m3WBtBfJnsWO3/M1FqxZpDAePCC92pPAfLjJ+Dp5B
ORI8fj/EBQmhyymtZlzcTE/ExxBNx6uGW39irzpyxh1Qf+qzrIANT0EhXrPSUBdkuNJpqJkA6HY/
lxOyGcvlf8GruSNKcCjek2qYYaCrLezawJQK9Pxxs8nLuG0JsC/9vwmYme771n5I/oU/oLlTc3o4
ZIW1R+PmonweZV1cgiahwC8rXzmAzWo21FmA7SLpdAuqgOHo88F6NeWPTEWDHpbo42tO4JhqFgKB
4ulzhoNShgCrEtvgpXTzaYp8/A8W2CVWRUfqfDUVQwiQ+JJrozOt1oO+CudwoZM+AytUk0oEeKFz
47nc0X4j7btONjE9/oPkl5v6aAJ1B+mWUbbuPOHGMB7wMvAUrq4ZfWy78Q2xPVPIkjuJxiHECeSU
etYt1TOn/93PX7zi2R5jaI9TCAl0M+LNszm98Yc/dcvsBO32KGKhxyipePsjikxHRqKAEnqphf5m
RGI4JfQZ1gVPrXUPGEiOUSg42VAz3QwS+x5TopkOMaXPbd+BhTJx70/Dx/vm3zovrEiH+yq4W7zM
MAhVCQzqZr/YMKxgAmFQoUJ2tvJQCYSLCY8hw3vc/CPSjYqaqgvqody0lDu7Zj8T9qow4ls9kHTs
zmWU79qjdyEMxq7s+4TX2jKHRoJDKgHRSLqSeBGIl6kvZHjiLskbVk+/YiAVWCT0Il5k6fAvk3Yb
Ii0zBn8LRpz41hqsyoFR/ebeJQBjpZxa4uFYxcZ52gSMA8h4/z/tNVJLAqRYVfFUUfJqYZt5xe1H
jy6MU7GWntnMC3v43uM1OWSc4sTDlTE9zLps/6Gak2oT/sYnb3gZwPF+qDPbj6L2EWWeWSC1di3P
KGpQZeIaQ+fjhuLqeJ5VgJyR3swHZbbZzJSKvRNsyDMmzBJpE1UiDOyE4pYlysh0lmMWKDTg4ntq
3f93Ipy0hNKBh35bb8qSzscHERu2uGX/SzrvJ5m4LOzzGsv3ZVUS39LFkKVFuL2R2fqnXVm6bKh2
ZVM6mGOEKQK+VpUYUtTLNdaZmMB2Y0Qu5TOkR8VX18Ae/PI+N6CW4+pIPVZJviA1WwFm5/KDB/U8
JMcw3F/pR8Gut/UH1lF5il3I+2xyQ4mIWiCbtCHyfdt5sKs9n19alYso+P/qnQd91Kz75Th6L/iD
IYV/SjYd0H2C75FlnsqnGWhJEAmG20LUah0n5Bd6hfuZZ0cACt/z78sWsqfL4PZvvwLzzRhOn2tk
FJboaj1N0Q7LT/WWYBUBZwuc7CKju57Lu0Nfa0wJRldS11OSgzcbRzwLBUNy5d0Y2aYzE/4hpM9L
vheHmVcF47A4Bw7qHrhbYKzeEy9Y9afqk23YP4wqQlgW732FUyz/8AknxJ4kf6PzajdLnYl6ZxJa
mf+osAORHxqPhOcnj9CbHkl3IgkLcNtGSX0qeuiKBjwDDYZl8ByCEuHcXeilpwEZlMCE6no4aH/Z
RGjdT4xTLXREE7gzjPpp1UYyA+Ic2Gl02Aa5QstfrhgfmuqSN7XutM0hJebiMInPLQZMlUWh6pAW
gO7m/tuTli64wFM5Wpz30bwVzg8G4ZVgE14CmGUmCA1IIWZbXkJ5UrvX5dZ9CLnDGdQBoEO1YW0+
PTUc59UY7WRvmNAoHnNkipqL1wjxj5vWm1Plk4hlDihsncEuRnF1wbCStumY+36Sur5ZdL9jOaBb
E1INEVUF5Q9qxbbSDS+uXYFDbZIPtVBlwcvcjR1CoRe6I3ygmNTQq5B2E3XznM/owNDjlrY2nJiJ
JGn701N2wjeXgMJ7Wd5tkgAgi11oXypl+Gy5qUitts4j5Yxtl72zah0+g4VFTk0GCdSFZqawgwzY
nGbr4n4crnxYEfnDCm8wWC4XxQ3XqXpCsnL9ujEiUAG0pqTGoNIKAqSx4jt+u6ny5lpRmZzPJ0SB
He0sZjBcnwecNecrcV6e/0V+gSsk4uVk/BaI7iEKLQPRNuYsvaaofcPa7XklVtx1swpysCoiL5oJ
3ZE5bnTKhcgxOl+m4HCC9C9bPoV9Q/3UFDzRBE7GA7Fmk6ufySTP68iqWx8HNMRHnGch1Jyuwge8
VrccqqIqmBUsyF9PtUJFBkrg6tJaI94iPM7NR5jaHC1kk9aChqNSQPIEyFsJzAW97XwWGUETqc3b
4BeOWHME0P/99B6dmELUzUU0/E1dE+2X4wh/IWpqmTmnPl0bSvkGGutw1cMCqb4PZN/kEZkNNdkm
m+fjwGe34kZK6G7JCgJlhJNB0NI5VfgHEHWf1lj/eGYf0f2mn4oxfnyQeG+ExUDttCR1ppC5R1tw
tDhq+c30OoCXcakL5GsC/sAwDChy1PpjKxK17iqpbsEmKTbW9kWVZ4twYQnPJ15tTnyzoAgPsIDy
HuJqQ4mGWNa8APeC1TZ6e3YhZF4ciRhHSx8+NioRxxTd2/5Grk0+FUFrVlS8ulRNwg818RIIEtzU
7IofKzbhwQez+/I0hFjoKhcMC5bpdaMEdc5qYRDLprwpRJ7Kl7xQgWiAN4D1SaztcWglb14z7zmW
NeEYc7DHkY/0XKM1FtIL+N76TMlEOGkWqFA606mLb6on7lqz21eDh9SjeqAB3K6qC8csNgymiHMz
O2rufGweVqIoUJXpIrxdFGkK8pFWbuWv/xDFzN5BQw4toFSXeJFc6VpvTNO3F/00mVacXK+7eszN
cJwY4Tcg+MCo0Hai7x81cEZHDFYsZup+Pz2KYARsZclJdz3i/oc7qK9oNHc+EM4qBd4JIbLEnNr3
miixmgEa6TuQl03GLjFbV3qYN2KBKiNpscI5BIzqAAimB3tPoZOsY/W2k4dGh2gO4yrhHjKaAXN9
sq6YERjqOMHGKuY4bf9KPx1hW/aT37Zpic7f9mgq6qFVdh/Nbfc/r8wLpBvmIWIJn8+RvPSv7fi9
6K9iFiIUQF/ealvOazC0VCz6dWrItlymE2FYfi8bdRBSpXQxQaafs03RqWGFKV9ekSSQ5flgHHZq
P4vQ6dAMS14MNxKz/HHSAK5YT5Uc+3dHK636mOwfHv+jpsPT4C0F7ovOQMqqHqNUuvAU4J7yX02M
2qwOpk494QLCRA8i62cPQmzKGABRB07jMW3A4+Q67xmYD0XIL921AWjbPF5EapQFH7Y9qOH3lIc6
dab34jKR+TwkHnN6/sRczbW+eGqat1x0VaxM/a8WqtkJ1lcb7zE2yHYk9A4lKcUWTdnNXblUSnkq
GPoZZYPrluYo7do2TTt2wccEycYqJK1zAx1aBuDLHwvXu5I6TUwlARiV/MBOUe9b9gHe5sw5BxeG
3kxoNhKaCTgCmrHIgKh6eTbGtRtsytKluEvYxNxxL0TNoB02hsQcXR/9BCnpLXIckIQhhplZoXZv
XNUJH4HY4nRzjieludep6EuITTgr7QpIeoRiQFEltEPr7h3hhbkx9ze3P9e6bK9ZjS/74XRSs1eE
oFTw7/1qG5YeF2vd2jYSj8qp94wbHUbvITmB4aijTrq7gVxre8m1lPdpIra6Reagen0xOD0K8Sdh
t5kJL/JlsO6JcafMg6e98rRNmmdvJbSSzyaLp5pTMHrDqJ8nfBZ6iH2aMyMitwQ3eB+zEWZtu1dj
EXXiVjw8Vy1ZIC+zfhdg6BN7RcUtjVbLGSwFmpO7InPML0l+ChRbUCll9Jje9pZZs7be4tNS+BNY
1KXr/VFCo9kgV8eVT4+37r0IQHec8+rVmHlbYJeGgAmVM1uWydgFKG22InOrbVTl1aB9q1IJSCFI
76RvnkLLyEVs6A2V3op1LxJffJOE54rxsVMJAVcgcfcawId70kJcZvNjKTdgKDocGt9pVGMgxjFp
y16JlK8AEfpUNToWBDCiS8u3Z2moczKSG4lBEPUH8dBqf78hhUFIjHe7aT41qlic/0pEiuW7NtgP
I3tKYoY8D7Gf4BptB+1lYR4IQQ4hJ5BcK2XpraA3up1hek0S0/DOvKDglIEJczREY6gXzXsvf8pb
Ur2/BL+4bXVU8ZMz/9opuIFJ3f7lJ4+u7W3nM6Ab0yq/uxrkfpGFWGLuZXbjmGzQTO6EMxWPCi1L
d/7vOs5Mo0qk2uTGG6+Yj3inEr/4cokjZnO2+iN186idj5+CMVl+X4oaeZE04xjfTOzZERyDoLXF
LnWc3+FfA25mUUJL7oOi56EN4sSStS0ddGY6s+9mgtJZPv98x7afdVgaUCfi3o8hhkYUsw+9N8uw
QwCYypPE4xPQ8w336J6u5R8i/p2h+QZoq8v0hZdkRA4uaCktkeGN82INT5KQcFSbfyQNNli7RJi/
HhDbROa3FY8gzXUe+WTPG0nT3f4x+b+PSuBce5GFysMkDXAxTPpvwPHrxOaMdipuY3AlQS0u2xCM
XCFl9YTlJRIG+kTx/ym1fLAqyFa1NVdcKBgTfflKaUg6NecTDOxhOVZRqz46Fbl0OUlPEpNXiojN
OFnZikofXYWDv+GI+NptJRYXjElMLJGzXtJoqKu/6ZueM7sw2Lfq+ldre3Rr65YgTUftbe5Iy+1r
/13eZuNbSyKn8EkfWC5008LlU68WTlpQ7vDUTdIndIwZ1BJeI+/niQR7+F4vMmb7mmC6P6Du52OA
lcqg5900jhEJVImlSnuqnkAQd+emKeqaA9WwxvWPHpCjAXN1Gk0syjGtQmLR8vso3GCdS1RFIop3
c6U6UYgzvUhwRns7mfhFgQul8KiOXaQ09Cv9e9b0TKkTPlEDB8z9Nc9jB1zQDMR15bS1+di/ue7M
bY+5TL47iXTodtUm6bkMvpPakXl62Vw5QAXX/iEYt3mJ/iAcacTbn94OO+0Qps+HyTdJJ49QWLm9
ZG+8e2H1mMfeslfqHl3I40zgtNH2sjn4gWAzeUC5JUNi4uE8+aU0Phvz20OuMrJBBs7gm40Bc8hI
JjsCZSONip+xnmWYUnWKDZ8trvgpOWXFgSCnNlGlIBc8mCPvYrux0CAj81K55Gxx03RJbInRk9cc
UsvBkt1TMF5e8roAywIY7ESmA7SBOhdXae+eRbN9vuTgBPi+Ixd6jiibCld5Ad4O/e1ukiwiXzdK
f9OprEFgdrBixDttCM1/M1cAW7nu50JYgvod2250xyF4t27IFmEdAnH4ZMhnOhmrraBsFk35x4Oe
/lAfYhSayWtR786D2DF3VnLlzvl9SQe4CCdyvfrVX76yDY11mUwUD9DumnaMH9Ypf7DV5emQvZ2B
y26hM3ZcdiWOlyvPT2lltQNKT1rKABI3mqeax6jVpPyMHwYA+IQ5T9Fw3LeQuqZNQ70Fo2Z9YebC
f+8Y45BQVm+poxRawOi9AoPhAZilRxf7PS0qHkvn2kqIxWflNkev7NY0wZGtlIoCr9xLugR6HAK3
OqrEzusCW0nTLoMy5MomwLNKCnlbW26ESqVbb4X86fiw4jKTkzjh+XfalDT7Dwb9Z1bXUlzXdCLn
fJJCPIevj/p3hnBPSnbX+tCmsbcdQrNaNXCBHHqpq4MdwuoZDXG0jRLoLrhoVKGGGptFWlAq0YJD
wUyjZJ6Csmshdq2MDrpA2RLKIUjui9Fz7b00OzkEvejMbLjNDo+FDMZwvnbFtzxca86SG+YsoUfR
G8ArJrLOXlpjHI5dqhqexANo+J/h1z0AAmOyiBkx9Rql0GfFStK8lO6WyA0QKCE4iANofJVJbhMp
CJKT9aZ0cMkRl4UwYW9g4JPrpALCSOAKgbEqV8iRyRubU5vHQ6ORBxoTxU4c8eb7qhu2nbBZF9tI
PRwiWmjXSPxXQNEy2LjuupggKv6ckf53Yfvo4sJSiohHPQsUYgqznVVUa6aWss/+N7b3NWl36ux4
VCjBlQ47QTmu7XeGqDNF1oZUBedHNI+2oHstY6Cy48aHZIIdYhs4KrGgmXWRKdCQAAADXFK+EebA
Mf+kVo6BXRBTwQUJttW4mJrZY3dbeJxI/eoEfGbYFJLDezpvwzZRo3+1l67oSiTDs9crzNxXW4nr
V8Rzw6UWIt0ypu/PWi/N1azr7I8zJaXViFiV6l4riKBvcoizZwMaxJPeL15mMTjjMRCqO7hp8rjW
0pb1TU/RFFQrmlnITP8kKIYC66PqdFBO0ThAqflBZrMY6eewZYlvEc5mRz3F1L+H1wQL9oao32Qx
AFGsBz+LneH96gZ7BkxPCUpv/+BS09BrQX3pYVWsQgBQhhp91NX9IIjUNXlnYvLx4AC2AjHI2IOQ
/IcRVsQY+Neq3zPOylARgKcykJeERZEQ/lrwLnfYghg2M/cSDmQmB+q7azMfH3M2M9TO+AvKO360
NXilEIH8UGPK+7TXpQflsBY/MTJzfId+q0/wu8Y4gS7D5t0O0M3voXa09wDHBezH99RHHVAY17Fc
k5Ws/NpFGf1ECs1veup7t+0v7XPZzbt1ygO5wblE+ybYUZHXKHlc8cRwvd5WNM1mNPiV4R5L64U+
t6uijRhKhmYBcyjba4hi3VTHPJ1xtd+ul/RcibgntTvIfIj+fCJUMvUd3xDr/clrHkXDVXH1n/20
2zxUNZMgnhFXVOvp7/InSkS/fkUt8Olz9NFmksOBFObYYxBsIplBftf+WOwE60Kxamn1yQ4hFHRQ
oMrJ4BdgXumRwYnPFdOoHMw7P/K6rLu3X9gLFVnn6uITZnIUsFG16oqxCuHh6QHdMEe7Y9oVzp0A
F+bXrlnb/FOWgJ3MZyguJQQ8/AKyV5vNiaPb8t/F22+rtXeopm8M6H9BuUKzwVRy1fGptUyuI50n
JZBqY2+3jqykZPo+Zq0rBglHYggHPNQ3GgHRqXPVvDsqwiWvPhvtgQkC55R6JCr0J04kFeKw0kr2
dDGUxFHw6nZgwip1KfzFfJp94Yb25zG5lICOm3/X3LkPtpImsv4Ut7vjI4PrlGX74EVqvzrS41qe
OMt7xQUi4CxFPYw1q+R/EznN/2PCs9OyioGcsAv8gD/ybgC+h6UeWNjBv0OEWPUEcbbN3d99bzNK
wGgOG7reTueZ0IPAEERfnHRomu0L+6US+Y4487Yjm5VlKe2pHGXbMb6pAoSpDmKXKJo9aaMKciy4
1CBaRV61dXRQyxipbj+UvpGxMm4BmCiQpmkoUFduAU7D9XWSJVf4vEDOSqPYJldyrl6Y5Y9x4i1a
Xv27VBgoFoh3wXg08oFxpxlz4P+l8S9JmgA5n0F67mQPkJfX8MAjXetGEO55AogD7iQB33tLnwxY
5TBXDgwyT6ENTuHR52Xn9J0z6MvxaaO2T9zCauHBJNbJUtQV6Nrmsz3hYHlt6i+s5G2QbOyrL0oI
fiFDOHtgt3CmVUlEJCvFB0nBBZ7O/L3Gx9PFyiMPoG0PUqXIbNl6ZUUjjRNwoTl9cqTg+jvFxt9B
LF5q9VVFKPz7NiaJOprI5+ZzemxdSCePAOIKFg8Y9oylENAXdMh58URMfrJ1i203ocH0mK/bwfh1
oHNbW/fGfXAp2QPHJmi2/PRxtgW5r0jnpgNHT/kFAXjwBfudeYWjvyJaT1i0pbZp/cQ4XVjSOl3o
61CjR0NVjc1GmtLxJVmRTLuXmYmzVgQCnfR+6WXk1J+dbGLu+8sUa67TAxeZM6lzD6DsdzPuHw8/
XBh6/JnYy+eAqgTdYAayIfRO7dJI76lSGdnET8hUhoMltKhJ9P0IFFYTn1MErAtWg4UYOdQIUgmV
hbLJmp15XyyYLWRHopcVHf/gN5eK1mxEO9oPGIZo0WTS4/soKbPixtjUFTfwozSMPzHUx2xHDj7A
2QFYn9ibm2+LjowHA+lkDta0iqWjU8dCs4X2lEEVKiYhqie1efxS9BDh4DtCPZPJaNlo079udkxC
9o9Hz1KQJnDy93JJwm/aZQWLsqlcc/KvS8dgckZ7GREVJxNXS3Gygjal2g80YR1Ty5MquFYd6Oa9
hwfjEJ9sPJiwjqvgbFO8crgsX8nh3bJyrj/KZOdvM/FQCf5kS953ogGadb45U8Q69sOW5cA6qsEq
vJm0dytqQTc3Fr09Q4RbruhP+ZCa6Xct6QlKuz/cflUcO0BqCEY0i4ZTbykXgFoXhDBhGDmP9P+F
irkHETAuwnuk3tI/eOBW2fXTrWvzE6dsfV8KYNrjpmj1FoxHu+bEdZIoA57Vm9+wkfb09+akRI8i
sRkAmUM2V5Jrk806M5uMNDXfFlfaYY0t+Ae7l2VuSBAjl5TOsOXAwUF4jEW50qkeiiJpjbsA89KG
HZiz8r7x+Uqe+zQGxXL+yoqqkvtkIWLs+AP9IHwUcZ5MDjlME+OVXZ8flq7fNaSEOecBJCQX7L4+
08wk2QTJVbaYPWGl5cUTUBGVSUGD3P3d5FyhcB/VwpqUppOVHVnPGzs7cKqt2RtjozERfdnUiXZd
rjTBaMh6R+fxTZ+WuRx/PT9a2/dQkkFmXahGsngEmYU6DMK1ZDqsE87b/BWYXgLyS2xInBZmr+xa
QZd4FpdrAmYTAT9ofw5gdMWQXruSd8UIL+W6PI7croKHC8FUbYkYfTrjq2qj9UDipyrJgU8u/lwh
N+d1GXhix935CEgnNgqG62oLrsJvC6eBaAO2FYzJGj6SHvuNNH00U4p8NG57ErTOOaXRru3FqfzF
QhMj0juvupYWbyi+CpTfGzht/aTFEGDKku61IIK6TTmx4tdff7O1asP/6/ofVG4QNDcCJhb6Ll5U
OxwolFHcBHC48OoRA7yoUToCaSwJepw8mHcc5FQhyTOa1K29aPxs/aE19/Ho4LJbxfzKvEUjHTjD
NOAVc1qlCYOiAZ0eO8AHgbI2U8QzQPVIz7+/WzSW2wmMu5uilkJwIkyHdFNiSW4W8oYJNFMuW1Fw
CabSNcF0Fdomtx0Q81npvGo8bgFs86S79LG6f4lZ6M0nHQBNSRA4tYlj2XkHHr1N01dOW5IdHkok
KPJ5+t0Rt35wIJE677z52k4e62LTg6Pum/uhjRm+VIU3viBq1BLuduznNKP/w0OG/NaK0mPwezMm
Clgyji++0AEngOh33PHWlDXX/rFqPrvrDmFFyUeK6svbmes0jPBXZF5uZEKscpOxk07I7gjBkTIH
tLNH1dEpDw4QZmL7gS3ysbynPDalTgdYjBPrQr0pxsNfWm4+9gTbwW13H9KdNSrkFqeJ1s/uEte2
1TYb5S+N5wp1Ju3fdWlgHp55sz5Z+aetVV+dQGwgw/zBJxz0u/bCW9OPlok/wKqoz4QrE4Z6VzkF
N6XM8tT6dO5uGuNroXC/+C+9FNROweGEExQ+IfRhv4LrXw/+yYMKejAFUR6B4AOSb1LvdyyGIKNy
gNjokNTFTBZkKFW9/BoePyN2Hm+L3iBDsjul1UAzuAYZOGZYtrhAsgxlHMNi+TzpKUpcl6a/iBYR
XkaFUasOz/Ewp0BXQy8FR+a9DvHZj/v/Jqj0U6Nf3krGB8f2UPIsQ69zKBHj8XDM0xneVnCiPvYe
nkzY7wGQy0K10jpQVzrjkpZTtiwqzPdPXMwr4KDG2C+TaMzrLVDHCaxeaCaCThzTMLNu8cTFW1NG
cwFamDFschMfkiqlhl9jWAViCPtgFqy4ZF3c3+fhdW2dC7h6/6RUK/Y0S+z18dR1EBX3vIUt0EQw
QdOMjQY5h9eFPWjlzevxKXocHMN2QVaFXXEFiJ5BfawzrGmZpY898kf0m47vSDFnlZRV2dD8tLRF
/DZzXsINPa5Gy5YHMjQqQ23Em71s6OW/clV85nI3j/GIG7m/5UXdhbxYqWwyqrFSZQtaocxqKlFE
cMlGrRYSLlSmdF7rlS1PeYX0GAhnQ/XNn2cyt5flZyB1dP7d/gscjkPXqBuWA7eRrsmoPdiRvPBm
5l0c/5t+bD5crYGxHt7WhTvx4XFSwZEDRDotUU4H8meu1yP/noARced+BRy8Ngh/ZwJvwT9LhscI
kKCldzqEfnNMth/Jw+OJPht1bgJTcM2+eFkF/IeM2H4U/q6t+WH+JVpRFrQ4xrhiPkYc0jxDzm6E
XbaG7JBDbx2mnhsklGgYza81bIoh05OOACL9D+uznunburWMTdvvac0q3Ax62gy3S/iQS9GLcZM3
Sk7hoOGWuqbt7KflxQ3T2nn6EIIxFZy7/j7KeiakwMqoeUNoLN2YuTJuaA5SR7g5CHEaNYag8ifX
gok+lT8ZvgI0Lbw/rMrC6O/UmzjByl8WOgHu05vLDO4C5MGtob435vaUsDFUNAMnThrM6GC+U3go
EYk9RKbx1FNbR0ETF4m2oPsXIFM1EvoXYGwKETlEttbnivAiN98x+AG4fWjhvds/8OWydUAieTCO
j+Cr6NLHt+TxlTWFxq52586umgfQmgUZFuL7Pekd6rBJPt2JmeOEPTdRaxfpoC0D+4lFlpbUpvgE
3XeeA5CUK0FCO5ruPqQDGRX7z9TcjWCefBS93fCgOrne+EhpyYjvuBFZkxgnJeypltm6JzxzL/Oi
buPsur4BR6dE1XkpQyCwlcCBKULEjpGijr+8+IG5pxePeL5choqPAkT9jMdZWuMwD1OtLLga1UPT
fqY3/YQwvMDwZjEn8okTUZYnLEEM/bmZ27eYZzl1pLfDsEoe/U+SQlCxTdnfz3m4Jhc8uqirTeXm
dI127oTzt0N/p4Og8DVVRKXgvOQz7yhqA2mnET/B8rI+mCeOWpDOJlzgm94EOZVl4fExseRDZarN
3rHXKNtWaZFbsg/bonD2Ys5tYggzR1d0In0dFUNqVugN2QwwXQk4uMyix7fUewjulZbtGeW7fR+V
IRrjmJuKO+tkx00cVlZrJxelYzqySVjTVfgQQHXdD9vgiT72E9AfcTpaJykzfihVIYcMIOO9uAPm
sRoMb2o3nJCps2dGcprs5rV8LjOga0OXoWgwUFkmROyJnDWPKhTPkU1z7Dg7WB2ROG3ihxnLIImi
OYsl/quS6V37GkEU4VCSMd571XbgYwPaW1aWX5OjWn18OH1xeVOELUGgY//IG7R50xZTPa+bMtW6
wm11xAh2GX9ce8hyftH8Sz1lBg7kTndPzc1eXWGIYOfKaVjcO6IH1hR0en7SCHqPzGESUnEBE85g
PpJQmgYFvJUmG49aW/RuTg2p/EyNO27e5BlHZ4TKG6p0VdNFtC6chpRDuBs+7rOFNs7NYrfrFd8Z
8VJeikd4CxNn3kmRirhSAXAc++rJED1F1nZkv7EmhhTodQKfhwurYOUB1I+SI4MpTIkUWRzgLpRU
N6vJeG5JA+PPitTqda3sHe8nyP+O/jv1jfaxubJ45uJXTsEPeIqSFKKsvdtSv09FQGHz0iCRui4K
EiackutbUhJTWUkRJHSNBLr3mVCJglx1w3uAk2kBK6BQ0+oadt5g60f1D98FrA3na3uf4eyAzv6Q
JVopoD2DPRPKqBhPN/a0t8QlLMtqzF9EkhmTpboOWf98NjhjmdASUe17q7w2W0huQZpm5V04qyVX
mgkdlSZXCVC8XI+SYSl6fybgv7XCu+xNtVDArrGRG6LLMUKboEiU/ND/yerDEv3xc17AR+maYJHt
Yp8IJJBXjGAfEc8SpJU8AnPbaIpYl5sD9w1nVfoB4QXc9Qv0HgLcP8akFSCHW6CR9eRYurpWkexp
hQSljOk0GvLNwcdNrK+XSKC7klZ7Uc/qYMHi8XyuCfBhwgUFrE5kEVgGn/HxGrhqI+SuRDPHhRAA
G8xzY2OEv/sOLzBdoMI5N4+RvLxEZlcLP4gk68yQMABsazdiwMSzBelTUkXlkAv6DtqNYAqjYqCr
eSXnt0JSn69vfv8cDRIEXFt9rvam2S3nC5NWQz2m2lxFSE8suUdptDDss4pGBAqpbPKeZeIXbANl
o8FxFUrj5/u7NcUUroDTd7LVC4WNLgeDDCAA6tNhEkbpfpr9/Ehi/iy9Lo1FbKry38wLDFqCD/XO
Uj7jB3cx0aMdnal2V6YV2ZAe6oOo66Z2pv5qe1nBHa5kq61efuYTzYS40Yy7LJYuIOEMiLWdkfZx
REJGXOKpjmbbsPyWu0j3bSfyY0dj8h7cTxOPgngCxDRr6oMxAtC82wGF0q6Q7lHMIw054gE7Od/h
+r+ogI/pSzXSGwSn8gP4N1fKRs+UvyYxjomkBs3Rccd3uknFCwu5lH9tfGi0B8QAEiP3bw6jDbik
ZzBMJCT7cxgQKEBozOqVtgNF16lXi7W/vm9mGX2EHkRcRaqyH/w0mO6AVBwT5lOURMDx5CEIxto7
LvwLgoztI+Xrsn2qGpO1a0OQ410wPYHlmZwm0rZDOrkmGXv471QOo8u1UCWMjHLhEpqqYfOllIWe
uCbWZtKW25NtzGqx0ttFlDoV3//fA5myf9zVw7OxJex6QB2hBQuo9YEjwcvxdOM3Aj60hT9M022U
QutacxMNx6HElaSw7FOXSEl3ZkbKFqGeDO/LH70cpaHb/5Rc75yA9/Yq2MS4JbPWgjIDoMAwbYWR
oPB56ewjZDWdD+hU+rSS2aEEYkS4VbKu9+aS7wGuL6Pi+ENVfPVz1fNmdeJk2+qYnsZ55HwmNNOq
Exc/SLM0Rh9T+wXZF78kUKNo1iBmCxwGuPpaJzYYjSdhabpAQkXbFgv5e5bQfKszlb/qdf+mJbX8
+PGZjawhwgbB5/G0zr8x5ux6G3JFVcdT44OzPBULgE2a39Wxhs4+fDuOoMvVSMVxJ6fjgGajGR0V
sJtgdXwGg7ru9dVNOYTg+lD0mJ1WZcbOqqeF316MFjdSINo5ka7yjSJpAcdc1QiLLc56gj1VSpdR
geGSMGpLSGn0Pua50NVNPW+R8Ql2AaARF94OurRcFpws3EQvhLQe7rv6JX4nkJOGhrCZlFqxS5v+
dI7TBPhP5TQDGr++DikROlvyrJr40ReluKvo7kpR97K2S7NKx2BbAsON8dmghV3FHkn9z/4H67I+
qeUMRLtlDIUoGvTVV98WSz+5wvROzgH97KD2x/f+lAaGuWZmv3KEwvUPWoBfFAp5uxlsIm7o3una
2KLo1fEi5yDoKGW7aI6Xy6gTSGcm1ClpxhOvJYxgAgmJOIFB5mF7BH04tQ2+DRpBjw6rsJ4xl4rc
1/vgu4bN7QrObK1k0Q6SJX+Uu+q9Y4uFS/WwdqWJhcl2O0eFt39WkV2x01FQmb7tU9K3FrxCR5a7
N/isQso66SKsXjqQFseT4rlTpaDtcsBZJ1vTKx1Xyp2J02WaXhVh0Vb1AhY2Qg26oXu609SgOGX+
vLzBVGE5/h4m+gemYmBFGESKXqRdvkLqxXlvcCAmqBwIlp3m8gysswmNxmI3mV1DqU3YUI2UNttw
QNzcbIOW0eqo0SP7loW556xT9/lW9YbjF4Tc1XiXToaIUDkHELi7t/X/unlF7Y549TdpxRKQNU9y
v1URby9sXWMhlnDx1c7JbXpuz0bqL68qdA3pSqb+8kT1L0U0ZeUzPgoo51p7tPH67cciqKBtAgR4
LG/AfKz9GBb6IcQTAh+hOUKaVjkMPUxmjZMODw3Ru0l87N9HE6z16FGNaG6TZMIof3Q6BfZWf/Ip
UOlBuuYj0q+HSbkf6EabGtGS7ps/BrvVfcQmZdAVY5b+WM+I7Z7IJKF/0g5yRwgIKBuPJhjgStm/
QvOugjFr7X9U1se5zB2WI5+i4Mh99LCxQxlqvsEL2lO5xi85XKbe1AJYZMIV7WkqHuEzeopZGfIx
9I8U21HF7eTv87wwYwlxCbfc/ppPXT4eANwnzggZKQhLUUsYp+XIgyAYUkjmSrwYG20LoOs8stXl
KefkDbSf6jMQUzOKWb3zQkd/lSP18UOp4xM6K6FSsuXBYJh+7TXWodBLqRNOo/6Xlf9b0ALw4R4F
y65tHO4k1c5B6x6ppB62B63/UjEeDf7GxSOduDZW6qyOu25d+8b54GSHjwGOMUB2l9ZQqcj+4Gxc
3n8jdw3Df0t8zH/lFWMNinDIJshJ4GneuNQCmQ6+PNzCTsE0xG2KDhQAW9eQ83pYkVrj0pu3b64W
KPqggRjp9jCr6tY7p/cYHXCilX9jTtJbTtx8QmjRSdNyF8lPO3WRJFi0EN0HyVtv/Dngxomx0EuH
QMWOIPD5GZKxTYriW9FTOwjv1nzDoz6RXxjJx0e9eeHeKHs7kuOdaj0ienVEoVi1FKOZh9q+egVd
V/ZWrXp5olZXmjsKnDub5XvSWXFeXoV41n1R74X0og3DVgqWGrncNVtNI0JHR29YSPZFSjco8WQP
fZwysEdslKWqNS+oQHkSKvCFdy+jBuwuAywo4wOCW/l1x7QsZ3+w/opHw3ncu3S3DAEZFxna6TIg
kIsagb6uuFBOUHd2sqiC1tZ3q1Ay3WtQOtgYtZ33Gfpz1w0FFXNsLxgWVnUf8ff+6W7rtjEpbikO
SGxLQud8QmoKAsD0bpgiaD04yqS76dkf7NwvcyCEq/HPYZAKsoYHWkXyVF6ogr8ncEG5nMi7nLdF
Ejq5Gw0RJhYTFQD32FwJ19M2BpbIKAJmOWac8qHk0n+8CI5VWR3mRoH3H7dD9VDF0GpDT3PhgQeM
V0e7FZzAitVT6/Zq+gczDSNmkH/PLmmz5V2UpbQpeipyv2omKXhYzPMuhs0567cURbeGayjx5aRp
nO/G/8fQjroFXWAHaKmLsPUXIbOjTgU2YP+KudhblmfqDrzHorjKmUsQCraEv4icJzfpY52yJkkc
y7AmPBfCUfDx6j570ipH4MpRUNmggkf/CMXBtr9MliaIUvlPKECpikkH4AXP+wj3fGHCop1M7VHG
VH4b8KdhtyEj0VudL8NLd2TjrjYKMnMebYMid+VpKDjeSkmQ6EKMOaKczBFe/lexHEgoB+8q7aR3
jOJq/AZuwdCLN/AW8vGWFXKkOrNIZ7kNTkofkMmvTLvI/Ao1svsanA/cL6fePzxJZrh9TIqpbzmX
OIXW1LYnQVWzIFxc+GHey9jZ3+FxGFf27J05vZ4IWos3tS9F9j0U0mB+9SFfBnIWy5WrCexsSBE4
9hNHLx+pT/yjxRxG8/JejdLHYQbiICIXcXAyetmCxzbbpMWXgoIjS1yJSNmCUIX5HWdof/LFkfBz
vYTBU2o2TwUv0MKfg2gkLR0fMHrsNRpvE2l31erDjhpDwccrIB1cBRc1NdQXdpjSdK49cWMqryB+
bPVKIR1sItOHSjxuYjH2V9wx5FYSK2e6SvprdmmlUI/URDP1VT+/1CnktmZAsbLqFHS/uwPsW2k/
ZOC7KzhmIMgt6be1J11EDTXTvS+5ZgJHJc+WNvePbaM/kr9L2t/JxvXn8oUJcmEEpdDs0sL1jy+B
/dVZZdpD+gabTUli08UkBkQFmM0f/HfVmPDq6wB3/QszK0leqoxLyU4Kvhb7m4QQuwE21LStoG/V
DHKEkNGX69JX1/MPxzC4Sqb+DwY/rXQbh2Z8hqbyBSNO4KXdAMyFWgtaPi+XSPimwaX8R+44yGXv
SmA09qPeTx7U7FmRyUMLdP56slPbdE+avqHVLk7rbh0W6SUtBdEen1PAf6g/sxi+xYGiJjT1/cIC
SXJG08ow/2EI8pVbPxPFemb8fGUR59sA/nfFnt/ceq3NyRdj8qM0fqsouwYlBv+wvJl2Ure3FUfk
/DEDkMC9hqw8Z30EmdXMG/hJy3CKhWOs34WT5Q9YxqncqjFkhNTYOt8cWVuvUYBxHV5g9IZ++slh
lr26bq2aQN5u4roIEEMpGPxCe4gxqfS3LnjIPKPwNisq9QhlPTpxpLJRlyarTNJYRmgr8abq1hs2
w46+GSJCmi+OoaHJEsIZbygsW+WeEduQvXygqY/OventtaeKwU4RcEnviUDV4aFPN4ktaTi5BfQ3
ar+jtxe68uMFoOnBa6k9g1QrDljhXwohlYOZXdVvu/2I7kNUZ3IaSkGPYvepYaCKKFxEJs/pBb90
kfBrEJgoXaanBsHRR1+hZxH60Nogf8ZOg1CQfso62xpX3WjqqpaYVXUb0mpRssQrEnY9SupZUnN2
sHdgSPI7D/Jivuc7PpsNw3v7O8/jUxw9sjST6wNvf2FG/hTOL1djRjxGKpH9IjFzqtKfCLWxkTzw
Rd5jfRDtjj3wJt8GzmLeLQWHsQ3dAV3vKLh3D4PP5vBZGdQDz6gcJN4dqHC2sI4g/mnSga6/tH5o
c9MZXwmxoSxEeULmepa9RxxzpTLgCH9Ui/12niRtc7dIQ2ybabhnG3/RZLeOl3vo2rPir5/W7AM/
SrSen5ulMC0zPsLEf4lh/Zc7wvSvlyTHalthSTo8GpsNXBzbH+0Q6Lm9wt+2LmhHuNgbhvl9yUJp
90jJQmOuYZNrZYDoKTwr7t0eF8go4jEO2tqk36bnceVMIltdz6FRrabLfxcPytJblf7Pize0QQyB
L8EQLtJ8fuT7ZbFUGyp9wmChIVqi129CH8aOFAKhafh69ftaRl4LRGxhU+2VidI4+yIs6PbL3yTh
QTaQ5DumWrMab96YaWMHX9YqMC6kxVxyziYZcsYJ3PwXy9sZBPyO3hhuUbjBltBOyA7kMy8LRHWw
xTgQJiEyu+ShMB6yVRvEDoqfshdsxtVFK4ys3XSwZAPDUBALd6iTUUd7pfpWyHcIgoVIaPTehN+W
RowWGwFj8CUcm1mwI8JsTuQvHgvDEpOzezfrUhHB9qayDY5L94SN1Dp1sSLAfQ9Yyw4VcVmE710H
8kOb0gJ6fZBlSPE7FgKrR7M+Q9nWym4CANh656xTgAVxnGwdrEX+8Irw2zatla/bB4ZO1oP0XKVQ
g3Y5d/wF+G14a2m0huYYErMhncmSuimyOh+8QMGhN2uqIDmdMG8PPU1I/vM1LeK7eNQEqADDQ+WN
hfhaGjpqRHiy/7c9VZI7Cr+BAOHQw1+ZXYVmd4duFjsZmhOTuYOQKqvr6SdH+penQXwHzWDHkTV5
wv1XeVbG+GFiCvErqRMHOh+8AdkFTyShkEOxytZVvk+c6BOoJqgnps9De1ek3luV0xpUFXLbAaY9
F2Ed7nRCxEuQBQYZhbK2LJuHv0dhiVSdII2NCWrAph7IaF4UOanoj/D2yihal8QYCJidL+0ccVrF
CHqzrIjtq3bFMreUytECJUpBWIBKKvEgLx7SA3Mt7WrTSm0YfjfTOdGEAm31LrpwkC+Nrg/0TMsh
hVcragJuqtJJyBjsrE3qpEElb+XypKUfUudu1JI0rE4ngdztPY9iAAvf95znRXsuEn4VHEDwNdwA
K6xocc2y3JdxYtU5iM/NUnW7c4SXejaHo+3iwUq/9uIqK/+7Umkwmf69yDTvBS5ifHqTXVxtM9HO
3ViauOKsF3SrMPM3L6rkmL4zrkhHecg2teyVZOv2LmDzBUlfRsYs/Ljp07w2TLewITR8xonE6CwE
HLkmLxCXBBXVMgIpPkORBzpD0WN9e41Y9xK1YfgS3Qcaoino/PoIbhHPuYd7w84Y9j/pcBmeCjWV
dQiONZHoes8oDVzulqZ7c6ODGYjBpcKc8NhfS7sp6YkufzyA3SpSb6RAQb8mcT2YzGmOYxxuCdQm
7WqfPaXPUc00bZVL1/Gkc8fqerQwgjq48sXdDiQj78DHYVqxgVOFvqh7tTJWfxTHuyekwbusYUAN
ygv5mr3w1iivwD7KogGymuwpEr2ORiHCAzLNPE34v29oBpQs0fp8IBKND65ngH8S/VNcF4Q0Y5Pj
LiXuh820OV0jn/L6sn4KfpyB/I70UvugL93ui6UBeIgxvVFaK5aGBXuMy4+eUd31+LiL+PnsJ/zc
o+6qI4D7hSRZ2pOzLKZRHHp93ilk7YuqANKVdOcnuCBl+ISx2herVfhBlbrzIG4/XY9x4p/vHFkE
vMtEA6uv0004ixYiHk8bs55OGrl3KwphMqHoqrOeYYIBi6Ycm1vijdT6h1ktsoxM4rGwGCD7d7Gg
8IKGePYwONo3gNXyRB8RLrIQGMcmm/mJo0mCswDnMP5cRmhhhhysd+52g9IO1EV9vvRfp/Dvmks5
CljdD27Nhns/wzVb2oJylr7E7nLbemblIyMW4mF9qRkL8efn4nocloxDLUiFURufBvvj9pDJWu3X
o4AeNUa1cL6h0QPuiuLiMpRHcUq/AAVe8lF8AsAcZrAjOIj9YkCERrhLbVSjYvyM5uxSUz+2CBb3
jexDi++FPF49pxVyVwKh3rp0g9AZOvcmbdCV344S6KElBfpZcSc6Q3qM2DGHFq+axxlkIVASpd0Y
RqZ/lXKKXRpdXh/coW5czlB5UssXv/XDfGegJHwWWHR8OzRdOprkDO4yMNveh+WUXiPQa1ahU+8X
UxEmZzMlcpCCyR4hiJsHSV9PQx5k/ysrGNmEMnaHVxIVKb+HfzG0itr9C0fksrep/frL1cypjnWF
XNNYWW+/VymGTRj/sjGikucx4jBI6qB8B1FpSH8f9t5sWCtx61N0h6zh3JwTpXVpRzsA+kc3otqq
1rIx/plk4hSZs/gdFDwBCyNCw9mc8WscwiXdbF0v5ii0LvvK74fzWjzVKxRR/1Ba73nmfed0To+c
M1XvKESmv6TpK5RjG+5ag7A5UmeHVVF2MVWkIAgwaeM7/74ctz7R5AYukKtjGZLvetBf0l2SQfra
nVY1KDVoUXj6t+GgIK3vZHAcnYImpMnncf4XHTW0EThXY8Jy4s6eBJKNQYU43fwO1J5y9W2TYona
WOLkQZGzKUPgIxkzPUNclLe0hMx2R6CZbObBlB1cBxlUqclgBIysP7UBFadZMbQdJ+Ewt9SJddj0
eOra7AZS7Ck05da/TDLI7f3GmtUPQEH+HDi+pg8OWCezEbTpuJcLUjnyqn2RTNM2ZNYWSQPIwUXu
LBLU3ocrEdm711YwLQxXFpucu8D4Ul5As/pduZOWO2ExG4G9MFhUf2fAL3mXucQMxN9xXFg0AfzT
SF8mbJuP2TstsodJ8MznqK6vrcOs7dKRg/IS/Ofqkjvh75qeZz9qYebPCnrXsWTZKF4HnbxxWngA
pwCRgv3WWDhU6nQxKTy3VTOKRbJElg3PWUknSJoSJ/gB9d82ZEPMCNbOKkU0NYYf18fmU7at+qb+
z1U5zO+6nn7Ge+xUIwnrNzSpT+k8L6/rbsgdjm0sqMRkQs+Uwl3YmUUlacBE6JNF/uT75lNbCBxm
s4JPMlqB/vEy5A+gQwMG8nKJ4EvF0FxhfxVgTqsuQ9TG2NC8dTJneD0CLtwsJxjunSkRkrCUdBPz
kGddAGmmBlHGGDEiI6/k9G4mY9HiSSe35L8VxvGiENjPTvG29aZPhKUtaeLYuPWNNNQAgI/BN4Mb
Djv+ihOTr23zQUWLKNuhTe77GSXmeGORCCwheFFkGl2/5CboIN7yGMQSiv5CDlzOz4dshzL137XJ
Rnmk3pbSOhDlQAIxIJq6zggdlHME3y0cBNKC2oyXs8VOcEpuCyw+5k/mkrWVmrZBMMIK8qDkpzsV
3tbfR9ZTDJ05S8j8LsfJCty3zkk5rGVKmAsWd0jt9PaDy/9atacLhG/2iQbZk114OcwYSS0DScM1
sK2dMrn8OifMNl89TfFNzn+yGzaQqPBWrlitGk5mwIl7w8oPKBpPkn3ViHLkiUKJiHgDqQMYxhoy
Cl8LnZajdEhJr3uJU+PZnYR43ajKqWivkkuBZ823jCv+pByViqRdQ9STjRtz5dI/27oAWjLQ9Mtu
jJ0DhrFdwbI2xkQcQcdeiqoakIlTbP/u2XeKdHCR7mqiBlY2VSvTycWxcoeksWy8DvalBA+Pe3h0
aXIfkEt8pqgYIVFgU/51REiqnD+AxkNAOrVue745IV7UWaHpJVx7XS1cS/NuOepUJGg7J9HFzye9
Xi4Ryl1QaqApfp/s4yI5DNnDCx307g8bqnGWDrsaiPwEPT+AjPKO4mr5/bOJD2lKwI7y69DnYzt9
W5cxHy9gDbDhPZ0G7zlSl5apV2PWiPBrFj82Ye1x2VsxUyovPEGDULFo5FAoy3NPdQ8xA1QbaQLX
IlFCUfdG7fi0EOT6E9I7SyFjEJqMSB9IrSIX6WykSHw6JnJy8fkvuo1ReP/VgdMNPL5Y1MxK9Mlg
Ri1W/+TjNvUr3L4bx5fE4n0lNsopkGuyI4U5jGiQPYU6s0AYZVYMU0JrlnD+FmC/IJZOg8y0AVms
JCLa3u3LE9L19tQidHEfBuJUYdokgv8ogS3ZtJjGkNN2Vlk+KzVOlXBPZ4kvLvS4tdaytV7mUot4
ZQi4Y35na0ZoXhQMxxu8MEO2UUkHuuoDuTztEkgaIUohWnYejXT4Nx81IyFPp60qMEndw+YKrHnf
aQkteaF4o6YJYBTVIuQSofSvQgJy1xrVRTuSjjq7m+nxULejNjDZ1ier4wqqYtSH+JRfZ05c9y9B
byC5uiUNjHMw8vAfXeuvrNg9YXYRUXGXAgSvsX1UPu1SqIIcCvKxFhEQLQdlZidubMJ4NNEQdTWL
o1OEf9kEnxYYuoZ/kX5P/N4Hx3fULhnTFqJYJfusWnW2Lp06ECI5AkWTvB1rcEC6LVyhR6i+BIdS
C/YJUo4Dk5izd8+M5ytNAUZhUszmIWLO8A0vcTxFeH4ytXzSpcxOTuiv+DiASfyWTiX+avhXqatq
ZfZ33Vq8z5RupUXKfH0PN4XmIHt0GvIYwgF0vEVxKzTlT7rl5OA0nExOny0UlLWw35RoPOP7XRbR
Tf3mNiLQBGwHgiyALjIcbkJ4h/HHVwGWOE55Gty8GZVT7018nKdKeHx1SpzZp33LIeXpTw0tt9Uh
pthPbl5OgIWcNJFY9JtTbkBuPuZb6YG7Ojdiiq7PT1llDPqS+C8lqBb+0v5HCDv7owTC4B7Mh/Ce
YPt3ll+8SggJBOSv3oIPWotcheXlzKUDMbz2ylBdtqUH1KFdMxtQvhI96FMJ3nibyZcT3zi2dTrV
ucbyl1FZMlIJTSVQ1M5tGS05MRob5ig6qABl9KabSMY7/Y5jB3DjGR+ERpp2Xx0wx7TdGQfolB97
rUQvqH+pMowWPFDG3RcwxX8/U+BNHam32gGeoKj8Q9W7AuGjzMPIh0tnS0q+HMb8AXgsYd7QmVcK
RrJnquR1UVcLdDJaLGZt+lrphqDW/LPc6bnIAekYhQtkS0orfphJco3c+FqvF52h3fnZAm8lURtV
omvdhlkhEn7U+OdTDco2ZgnKtZTAYFrajwZ/hPagw1kbMoF+Y4KT+HNpClK/i3EQvtKZGlQYKMJc
URTpKReFTW3YtBSe3a4gh+FsIG8Og94hzAzkwgOt3hAFFhY6T2MpyaPClkC30o0++wuGEpPxnB8n
sfMktjdG5HlBKK6BiEP0RceQzsZNEvxGH/uNgILfL5pdaW9BJSJA2Iv6xhx0dAlyiqHt46pwx+Z0
imtDlawMLpB2e4vvZXyEoN58/MsNQtPjgo9eVn3uaXQYkY6lsSRd0Kpt/mxBL/sqRmtgTrBwE1o8
FfCDVWaspEAN0Wye4/IxrTfMoZS5r+tBnN5OAcvU6Xtu/GY+euYRWxc8wHTzlnl96X51wcS+AsCf
2zKLJBhgzjYhno6AFbEZwEOq/RJtDFowg+9xGMOTdjF+8JWycPVOAzLi8Jjd4/TqyKzO2ChMXD5z
tdKpBq0KvI1EpM0mdswq9dN+wOsj2GHRYghsKrkCHKxWAYz+hehjAXC2qDFIqUSWHT79ZDOp4/gB
hFaGh9CJrnpD9ArbM3qnuZd8ZnHzvK5+UPPSKOuF2MnzelHn9BtLvoqB7/KVdttBzn7F/SqocIU8
Hxs1wXI+jRWDfUhjQnzfcwMVAidu2KkCZq+MG4zZsvImr5/Ocn0ipZBv4rR2nU72FP6qgnLXacx1
z6JsUal0hk16eqhBuaM/DCR4ay5Iga1r/eVH7E2PlX6Jce1PuTKU/4f3UlXlqoA0F3vPOPAWI9cE
pgcGpHRNUUfXKBkMFX2kJSheTkQGFYoRrOIxADZggHjr7NXddZfK8LTbIGfrEi9hixPXGAU3LZ3x
UF2gejbZ13FjaLpMe4zrD+AXQpQ5xt/DkmufPr0sGRd/GHiFJmKiDGAIc5Xh1m6XN5iIGxZYGjMI
8X9/3R0KVezo5aMRu6A8yUrpLWMojAlDSKOKaNBnxXSK7ZrqyYNgOO+ttwYLtiUIXTx+WRkZJx5l
0REsppjbpvD0NF3ekf2S+QO5HmH9Lustv9yGGdgyS7El11txcUmtOD0c3lgtH8KV23UsaZ4jkQMq
u2D0RYNQwIOfnnBehlcHZVmALkgN5RI5NoYDG+XprEIV5i2gqJFaRBds0pv2oqvOmdg/+tEBzXJh
e4CxBedNrqsGykR8ZMnhADSTZzq8QxPqR0NF/vbsqyskCCR1g2HlrlaIjH5Xx7o2PatSjgDsmw8l
z358oT0rC0Yb9mR+HlFFxr/xRsXHoOWXqZjqUjkMDqC8djGnGgVeAECUbXTUNkv8+H53JKVL+ARp
KqqylgwZAaU3JiocVZkOr2apIoIo9c/4F+mHEEzI1Wayw5fiXs19wNp6Y3kBN2fIRDdt8nNlW3Lv
hyVIn987/SRD46X4CHV6hXqNU4iCYWRDp3OECE2fWW+U/ivu0Elne66Xe/Q53OX3xCTdokOqR2sg
l5ntJJEC2I/X0bCZwL0sgMG9UKxZPeNEhQhpzsYBS+6IJveuibn860cMxvNLKDdgJW9QqZLsGNvc
R34HJtzPk2110DG03OHH+QyhrJqlMrBKr6+HcM7zfTLKthb5ex0EHr6Q1Xo7WcoIjNc0VxM3hTHo
cUDrogkUs6fbcgje+yU8acJLCV5pqGED22ccWEgz+AkypJGjp6xhaZHH+d5R13JwLYcXfNbTobTm
G+wwKXOxLvwGR+JvKU+CExP9AtKRP28RIJ8ZvqM8B1V21WR7z8JUvsAHeGosw2eYhOWkL+A69vsf
bZ+zaNbD6rV2B2LwcQdDxRFsdOkg2BsgWCNUMcVzezrhJFkSdrJd1ksftCthH9tYmsJMT9XjOJDE
ZR1Lm3dbBRYWljfCETWehXAsvTXfnop4d2EOW+OqDtQJrNzcsUpZTK6mebb715a7/bvbZGpX/+fR
v7f0xBirB0qThIRzdGj/dLjabAo/KfnVCgMggYUJ4GdF3uZVHCdrfBTG+5Bv5XJUzlDhozF6BGpn
m9rviO8ZVy2ZRtvA7xOF0zlCoxamGzayWAr5wgYt8iLnjH6PUjhKmTl+Tg71xOAP1RJfZ8L8HoKJ
80kLvX6RguI5lY4U4jJNav6Yojrs682MkjPzCmouXPf962WGzV9z+UsAItxACdO239aWZ8RJruAu
FEN00YxDSk9ajUuAmDHIW4hD9K8BqMP4mV2ioqGf6ItPlmh/ALLbsXKiU3X8+janGsIqnwxi3FpV
lACFJ8nR9OZDTwH3E+9QJGYfNCG83A98XbjDVRCuFmDgQoJtM1ySL9O6Vra7vjcSDty1jEU3JaG9
sb93aaDatNIOESIC1NzZz+9I2uBuGe++j3+zwwplo0vU7SsFOqiH5CuhJmn7NdlRttcLKmQMKflU
+jE+n0+Ae/ZFpTUaWaKPS4S8jNBR56JRW6JJBFq2FQNcMMamthLhvGU4YOzSCLAmtfmfOItulgG0
P3arZT+d+tCVIdHM9myUPZXnUf+8pC5dFvxe3BkEe3rvXrI+WaHDBBOxAe3MuLiQ4Cz0Io0ZWKKC
eCjsrQcsRWndqV9IEk3Wk52qHVTQy3oCBTEMJ9HbOtQQGzNGwn6/y2qjpKyBn18QnOLiaa04wAiE
YVDyK1+CzXhrmIMOESCID0nmFsQvoWsFsBpjIVD9VLGeb7eMdqQ4xIlVASJrlV2p0l2yqPl3wvlx
uEzlmskZufUn/rCgCuOXDSUoLKVpVHxx/jmbWYVj/dpxgMSbuylmZZOzzXtwl+/fRNvvNKOrRNx/
ghC1nJVHDyyFrXfGqRntSfxxYOqC/3X0yOKk+9LGIzywZbEADHUH0MfjdT1qukUMx5+u/e49vAkh
w4k8a0x4L9RYIOeiGNYtIXGNB9e/BAa+cA8ZHe1pxKuf30MxDctVHdDCi67KPY10TT4AebGS1+Mg
qb575VbLEvI8wUiOAG6dl7SmoahhDz6SCnSRXcw3JO0NjxcynwJJDlG0Lv+6f8i3h1Oec3i5Rowu
Vlo4BJj74+2kYXr4+zuy8dUvxEo+9XFrgK59w03vlwyCyEz6ro2QZI/zoDGW/aJ5xAHxwis4H+5W
QpjSSAUWxH1V5UClwNp6zN9NJFJorRIZbnclPWvjBtWyuF14O3c37IINDXe1xBboenyB4ivb7MGa
ZnB8K88SRP0RE8SHdOc7syQzWW5qCkc3PD4O2A9Ju7u3Tgtgsecg0JuVZFoMVl7qmLIb47fp1zLl
JL4s52Xs3FGyztclUlEhseTklT3B0w19F7Hd97gwxbeMgi0AaI8GzORxtla8yoi6cmSfMf12BOI3
wMVe9s22b3PYpSNQbiXtEQXdHST+xZDCDSzvl+n2lYkVkysa0Q/oXgSRpxIjMDirxr6gYMF8KR41
QQw9emqIyxsRCPlL895fAZZm1JM70fhzVPLgTrG1knfEMBc+hv9SiEBvvzFEH0aiaFcAp2CaaaIN
tLdEmEQ1zJEwInOEjXqm46xQi5KZLknhkiIKvzdBQsHY5u6x7ivSWL8Ct5ImPUFlbHxDFpM/5wHc
dpCC9l5TJspQBLB3Tm6z8IVZrkik7urZHd4z4x+o2/phRynbDKwku/U8fev93A4BwWpiSEcjxBO9
tTogNZZcltYwlv/XThU3jzVx+rISEfesGmriJSfLB8RWBRYpbHMeafPhuIEMlvCtTkTb//HKP9HZ
6z+2rkAhuQYJueKROXNhFATHICz7Lxp/UKYafYxoUp4jSv+jBLtw5Me6JAq3NyL8ILPVAXws4Ypk
9HHA+4NDAy9Avqqw/izCxTyCtJTV41i1XX8RgFiS4ev/k9dqst1mjyFm0Y4tom+Kuj4a1IXQjbYV
vrumG+x14ofJhmLyxLUMn5f2meBozEmyD5REfJZ9Syf9j9TRlJc6x0Gn+B5UoBLsqdN57RjMtFBU
9hurH9jS71/rDhQmjVZQAxiPJs6Jkowz6lP5bAxoGGyakcvOm9shZ9o4fwh+fF9KEV6mR8eNJ9nh
5DCRa/g0btcHA4+lH8ZYTyUT3rMOWew2poAOlM5gl2bsaH2S/PU6rwPWiaxbT/dM3X94Uwf5T8xW
NSXtKTkqK+6NuHMhz8xUG9cEVXxQeMK7QqTB0bKwIYF6UgImt956PhKYRxMiKRC9z06GJsDwlhvK
8jnZMHLckw5CxfUuuOxDcZFkREtg8V5mtSeoa20yZ2PxRw8lfKutO1d/PvVzptV6lLlRAtseJ/+L
5EnpgpBg96QiAdO7Z5nD09HS6MMxiBIuNvf0ECJFWC7PWgz+a59i90kw8TQJe9M4bRJ/u0iAzQD6
ckiUsXO+jRqxX15pl3N8uUYQjQ/5UwUiN3KUWbeLslyLEdVAXzp89JTAU+rSqA8FeyA2wsLzZ1ZW
34j5ikFqpHrx+5WI9z6/bcMrJISIGBpfNy3o4qYzC4BhQHICuXW7wbk3z9KIoU1WS1TTtB522Zdf
Nm4dabcCbdDATO2u2EL6rNQm1zmA8FQDOIgNS5qgRitmjp8WCyNvHRv4Px3I2V3cAN6TGjRy1ZcV
4prQUqmwbPIRLrcn2xHUsBvXNwRotv2uf5/cPAk1JZk4MpknCBgTrgwh/Km5k91nuHCXTLDeOFjY
/fCG93l6396OTaQgtHNToPb2SLWT5i/wViLeK/JfHR2UpBWqdFirSX2v8x+40HL+JjMS7Dte5v9W
2NeTWpz8UKcsFg6VBMc0llvGQx+QigHzBuzNYm8wX5AW4asg9ISys94WqNZkY0vF9r5XYrknTaYN
I8UwyCOolxbQ6iLzoKc1hXBdawYYrutIxO78DhcfYoMAmAjV2tbFwRBil/61lfe7A8Xk8oQaDDPF
xAswa/va7lO5JM9nrdR6Ewn8n1Cq/JkwC5JUtau7Rd6zBpyascuAX9av1j/4mnXTqgoV9O0OVe0n
tsHyjM3vghp4TJXKn4urUzXUfx6jWVUVooCuYCl5+6zrgMPHiLLV8oQOCzSLHCqF8PIZpbMCkQym
9Nro6hSRszIPT1qlSDeHxjvp0XsMavzLOy6LJUyNFZm6hxDTUild3S4LoW5jpmaJwaGBZTF8TB+7
l95M59VMxWuCIVeuc9zv9Ekhs1npZn7asrsPolvSklPDAIvMye1cSAWBaIgTfhthvQFM73aKz6Q+
uSaDs4uRE+514rFgxzkTcC/SxmK/tznQVBKR5t7zZMQ6u79wTeQGq6Ar9Acw7ysNia7qZfiG1/G1
E9rfilJy1aRGnVO+H4+HjEXNlWirkw89ToJjcv1x35Ib/8pBGsv0uOFAjNvQrSrwUNkB+gEzTsgY
Km1OBXWkISaBQBpqQdNvX0ZcWHHv4ue91fML0WI/8snu1MukyOjWR1upDjtEW+3oaBrAmPppUDi1
KfASVVPH0uyQuWA/Ctpuvsl98xdOgQ3CDimAcamuSInrW12JSj90Lp/4BsBU3NQN7QMzixHenVGc
FoQLKDFvAv70F6Xc7LhSA8W5TFYb3jZjmQYdNIt49Fp/K1d0DbSUIUdBzIDmAYU7n61hQ9eGcElr
CtUEGRTKUQhg9xo6S3HUWdEclXVugjaZz5/yfJ/e6JIeugFqpovI3CIJ216B+ZmVrhucQsnjylxP
DdKVEMcYhm8KPSL+psViDzpKSchpgBDvncti4JzmPYpb3tH8TS45Hi5W2s97BLVi3bH+Yv8eJruk
pNDppv07Nz6hus/uMCC7lIv/r2FS5rOyRWCsuZPnJk/NLwwi65CS9J0DD71yOrl0EaKTRJHPq+ns
HGQxNTAq+5j5GYIN2VAshLWOeICsQq5gSfSWL4VwmJEmRTTWF3jducI0MHnhm07tOLqAOWUiey7k
0yBhXEIIvQ+mLxyxWRYzbwYEgoLOKcux+S6xT0rb6YApXAlHjCT4IIXbNLAOqw2+YXhjzawQlHen
bTbp5Z1rYu4Mwvj9/lJzqyHeVlTrBdOeMUB+1C/6Kewp+Ke+yWBccWU80LyPjHwO4mQLTOkIRYy8
sRGkFIoQ1iU6WOEuKjin4gbDBPKOhUqhW4mxalCDtbFrLfFrV7GrG6UbO8MlgxnMB7freRvcsK/g
QpIuMkGRlNBaY27+M5p2C5r7WR3R6yidSk/KDCIHx0VImqGgk3yYdrJ/un8y2xNW4Uea+ZvUjQS+
bzF8DSMOKtWDLnfW1inl8xNENpeY4lg0NssK2O6zQa5rBJ2Dw1L9cQSMASfDNRut+gx+k6Fstcoz
QoC9KK8ieqCx5x2AUfJUbi0PYRufLTqcsNrlpALQuW9ihJedUaYqLQVinrrHc0BsCwgCPpqnXEu6
z1ifG5BzkfVwegIJajWHLTkciLJ51eGkjuiC9QV2IZhiCSmMq6vZ3/iTXoH8AGUkROvgK73QUqfS
luxe/LalcX0lQYcam9Oa6ph+EBK+sa51rvywrnmj7ISeGnCQiwKYmgPAgt0ZzG7YSXGJp3syvbel
0ql73OV1vKPeG1dfbXiUjSkaQo7WxB1QjzlucT3eQOTowbZ4Xg4342TAzAi7hiUq4DXmB5o7qDq2
Wlf2BeJ0pZAmMBqG6ElpTVXDouL01omyNZ8gO2KgHJ0CjGHjj6305V6kIGq/DRVU6Pw8TdWsFQNa
RJqFWUDfS8RNFKzix9wnwdMGHf8oN9NL/iTBbBS0j+oxV457WRhvrAE4oJStpwNAQeSq7koJHgg/
t9ise6R4KfBpcjAqSGJ/tzxxq5WP7R5KrxKzUYGh9kNzMibALM39ZubzHp7MFtJohzzgT8Q0xt5+
9U/Uy9RKwHD1ZyW6x09xzkgE8Zcu+bps2XM6fGZEqnPiO+dcntWEvp741dGfFuz/o2wuQW7tLnOG
KuMKe14wIzGF0FnrgAfQ7QduL2pkAQ7Zosf7LSZ7TIAo3sAtIu3th88sDqJrcZ5RGimSqOChi1ua
uornVLWpJR1lJo1iGffrbwGyoQ2rJ/RuXptQEFkdS27xs8yDjeLvj2fRE0WMQsBR/rBoYSEk4hBs
HAFtU/dRB8ZI5nrXJVKTrlvrjEuy9nSWKhBhspKqAbul+A0xaNxaKH3NhleUU+vLAO0Shn8Qmkpp
1qm7t6QNGSlx/Gh8smIXOANH5j7Blh4QAnkkz5hQw2WH0rGu1XBzPRA1OPStYtyLcT6euBTnCj9M
nMFp33aU3DZ+bVYJ3kadqcZhIJBmAkgCyOesF24eofk9V2xEM2Rds4iLI7TMicMrFN1bpWzP3EH3
DSIlaQG4qtYQk9JRuo4AN7x1zov0OIoW8JD9BwKogTE69ozbf25tkZAglhFiiSN0NbFLcN3Yp7VU
69z6oBRozalFm2rSYboUjp+pLk946pTvHm/p1N6qqYesc3yM2mKI90WdTZZmirTw/uI8+OjnbjYB
2GxlsEQGQvfImIUT/F/PTx92n5WTPa7vcVlzJmPlA7KIFeBLHibZXL0Yg4csGqfJAuDDgC3Mkq2y
KhBMgpzzw9S/vcSvyf4k/19+gRV1vThRe/bAXGeTcHTm/1jhYygOVVo0GDM/jrWssF2wSBAgEh7F
at6C0yJnGQHmuyYpcKMgMEkdKZ0Ln+PfU/DbYWuH3i90dcteK0/RzNBIlGVLWS+ZogrtjplHtRRr
3RfQRWNv5PhkaarY9SDEr8U2q6HFJ2uhg/EZmHxnAMEmMwb61REeRODNYrfH4oIQa82lJNwtskbJ
8q+2MWOdBThSBtQ05FlBhUxLAdVsCM7Y0HGbeO0Pw6oXqGz486T0KVOnYKkT0vk0RTst6QBGOIzy
1RRN0pixBHfcdZlHkH7q2nUkF5k+VmCM1Meqb6F4BhkmpPK0LvTvs4Y2pwhOKtg8cyFDuPqa7HFh
DYnrHWV/qiXYhgp9M0s6DoFdJy0Tsb8yrijTyf07i6pV1as5oeX+Yni1qx16cju7kdIeCp6ALFve
5WPSp69jlpl3L1yi6fKdXURkrhMHdc5rdYDYFN84wgnC8GSDAXEiQ3jEej5xRNBOlTJWyF9qRAr8
UHuYnHtqjEq9znks7pmCPMNUjGm1IHuDhusNTZ8nk1r4VRFR0f2Afl7G5nIcrlBwdLn08TJ816my
YblIej2qN2TpFnaTp4501ltrQsxNrjVcSO835b2QNKuhWBFDP/omALe9iKBF+/OOuuUsB9wTN7x6
wS4OtdphiMwK5x2rD3KJ2Oh3Gw95oIgPRCdsEyYn3s/9SnqMX7rRYGMV3VrApA0RL8aFgnaspXDR
74jEJCOOS85eQ1VECu3IK5J64xyE3TOzCnpcqNu7HVo7vGgMaJFVJBoQLMURODNy7PfszPItBbR/
CqsGJ9sivSiFjAcypqW3vlvFC3iAbaX8sfs7EoGxK6ObF/6tbKaPi405tDNK0oWJFJMofsfkR5Jj
wNK9ttUI+wMCjFefRnDg5YH4Kvd+LN7bDdw9ruBoomOJUWu/DnHnMJnqLqgr6KVaLWPYOE1JWU5U
38T29Typq/oPrr8SR0hwL8cH/W/pzMtpn8Rm8wuoP3kRlrImCSdCrt487418ipq6GwYW05p9u1n5
Wdo9V/c25eqYKWnl1An2TBR85KtPsUmsVzXL9JyndYwngGv2SVnLHonMCHRFd9IwVB4jdjHjksHL
XH+ekpXPMnRrzyOsCI839wF8NKT8KM5RIta4Iaq5u7sa6ChrlV/5jz4TY1lLZjaWeLp/6WNpUbk3
jKcqr0TVcKF0UvbMp/Ldh84XE4gTpqyodMudJk81EIbL3mMyZJQm9hP6dJLmjQ900IoVxDWdpK3x
9TibuYjfFRsbFZLvQu1UeHNPc5gYkA2vg8LzikqVkRQYnp7lsEpBhuFE+MrywYqKxrY7JtASonjR
agdc69p4HctKqIKjS51Qu6QjVrd1DGSvwPc1hOOuG5ja8aTM8wIkZ1+AmKLGRKQxecHEIZz0EqnL
DtSGIPRtiOf4KMU1JLww7RqSIwgkU1WIJ/I3BSI8lRq1rIFOtBZh5q0uSk12uS1NqKxyeUcaC2Z/
1gkGgzLJaoeTmHa1xXG+VEnBwbxuIzjMchFw5749jVtIy8YiONU1wpSAx5BfwAddNO3bcA6wDW6y
Z5UkrGkWzXLP83A/+v2xeJCnDrPvwHxcENInoxbUxW2fJIA4z/gSBhMUxVg/1quxVO4uq6BzOYrx
6w1LwaAC2TwYmUUe0XT96acGHcD1L3YFrz9STkSqVC9CiX4mkw6Q/fG9m4gQriTl/ypF5rA+YRLn
gSF/RAzMeslgOpOVsl9TP8F3rT94dBP1HLsMYG43sHY1rWhENuSC4iMH5hFiImSyqL2uGnZXRdMR
vtwY67YhyJNYAvh8La+mL5/diFRnXXyRPBprIPEmDr2PjjY/wy1LP/Ht42tVpKpy067GqSS1YOPH
nUw62Lw13yexdqp1EjQNJgXv2hpEAoOwE3LlbMSapiCrsGI8jdRS7ZrGXdy9YRLxRwWWGjQjj8Mi
Sxh4Ava6AkWJ4CH7hNrDIa1zTmCCBvn+evFjl66UOQIA+hc7eqrcOzbsSPVzoxehbT0uDqN7V5s8
Dq7N1FcSGakC/T8Mh2QkJF2fXd3ESk2N8XiTR1EFS78bHSKbDzNIsFKNbFFqrdsx3gwjh/3jljKV
QeGrRvIi23hnXBpsfzG+FIImBvnldl7vSvTI0ICiFIuQJuWq8CMa07HsbaW1uV09ugETqZytzL6i
n3FlKzZkuLnksgDxghAg8kLGa6bWnk9gGwxoeXEPhJ6fFs68tE6Arpkzg5IRt/MDX6aeiSNUHBFo
MXOi2+Gbz2FdZmEeyip7Q9p4ldpls/9d/4FaXmv4O9Sjw9NB6EcQt6YT/9+WYW/ej4YCtkpyuWT5
LPxdSycnTBgr+N/LeGPoxqMRDY3tMGZDkqc22F3EcmTjpdMAKr4CvuGjz90thpSAjpinyi5041Ke
vOo42QKHoqbnwaCOHjbTnjGlBWDxExLMJEqn0hhEjrxIkhbn5nlM9f1uSEaez/OGlHn15s33uGoL
I+JFwpDuSLOY7nETZgVKMgAcE8QG9fxuaDT5I21wLSwVBVH76RHUX56+aNiKkDaOEL9bsDEx3diL
NmsUtB2dPfQ1TWqbGJQqy1MEzXcTue9cyAsxhPDLtzxxvIrfm3jPMK5YBgwHbFGGQ4tliO70Vn1j
NWoH6nKYzi/gzv4fQyW0os+9wH24nbRPR6mjThdpurwXkPLUCH8a7YZfDa6rmh0V1IDtLa0j+2Yg
Mc6Mt5mLjYkeUKMVSqjSNAKC3+UWfLr6RUwMQ+/EN22seq++fD44CmYPGFG5pNCF1Et4rDq1f08y
pY8H8L7I3Pd/+HvbM4h7c90vC2tsrHstKjnjeInHjWi0sv/E/5itekt/A3kcKqES3OLU2KNhJXaU
mrVD39Dd5opPXS1Zq3t6wivoacEpMOX9sr0khPJkrSewrFMGdm/2EpgXy8jWkrCo5cT42bd9aPZo
tvjg4KoSrC+KqLqPn1SsZISG0AIKFkanMpYlcIvSiS1J+K6FypP+tfjbf/l1DK42iBVFbDJoy6Wx
GRUVViqeUGr+x3C9z8yjF6g3lfMPXCywwvKsP24OpxgRHQ0ze7KfHBPkG4sSFEv1nqkBz+86EBh6
/DvXMBbXg9tjLgl5S+SuIE/u1LxLeff3Bzh4L9HW6c0vMBXKe19ENVmg6X7XVwhsOFWCyldbzg1z
Pews70AELWyS/OKo+I8tO96OW/55kPnoij8KdBj5sln4Gnny5EGbjpwPFfof941lt40Z8eNgYluY
4KTaEEne2OfGsXFh4R709eSWtSeUV2UYUZSxIZlVym5HVaFRxN4Rn3yXgVuz0FqyY3tTU7kXuGsc
5n3Zmhf4Or8SF8ZMsRoc3+YcQGpDzPkwYkyVAlVED8JG1ug+P8BFVoh96tNI1UNfD2fl5IYgQ7/E
gdfal0xjqgqU4dHW4ZnOi9mOACXYBxlIV1cAEWeFZ0F6PMN6wGm2FosShc8wyGob2ztJ3jNPs9tx
DkRC9vkl2cogOwwRo+sLjbf7CzyXnPMcsJOnmqsr51rerN+whxKX1qVtMutmhgnFWpot6U507DXa
WQp15dfXpVe/E0gQUayBgHH6C2tu6gRnbyqGP5QYBMUA7XYpWT5g8NTW8qpodDjvmYwdM7T4IugK
rswoF9IVzrTEJYT1UDERWQwIS9aGThNCnnTA2i4U5ayU2VyOVSN59v9BDNU22EqyL3utVodo3xUX
t2jgOijgtWEdmFIYWEt1iAAJyjmF53pzuGQAEIDZfiv0qH5X+r2ec6ZiQlmax+nxnWRq8BtSDl5n
loZ9vmJncfdsdr06HNrmwD1cXn5zW/CQy84fYGeN5le44CDQeDL5mU7OsjmZSGhAXE0DG4p6re7a
ei5wDScXN2Lmnx9myaTT3ODK1r//TP/pwdQy173uxtKhPchnxpinfpndm7UXyH+NdnReTf+HpnRg
JBC1opaV73G+mlOljrus6c1WPhtZzgPGqveWPo6CKx8JcQF4C4AscaFx5i6lZwNTPER3RhgKyTyi
Ifeeqka+AbVU7G1zs4+Yp3wMWSSac5aSgekHurxZxbe6uYD0G4LN6s73bjITW569zYFdJzz4Mfq2
CfEq0b2O88ldXt0z4bTW8IzaI2PRohYc4Hraj4xptr0djLzHuY/5rcMq6H4XgtyCgkqwbsR1f4Na
J5NCtTAJvv1CSHqmIPOLts/ILCa8Jziu/bqFGxjzb87Gv4d/8b6LvcdVVUgWUKDC8DuksrBWomi4
NaFhYCijBu38kXFnPtunbuC7sAA/iRcr/O2822jZF6uIwhKvtavHv+EZYCCdORh+i41wP9btN4Lb
j5/IMuvT+g/aGbcJpsLlDrqkiPRPquL7TNjuE+GvZnMTaTU5SIlN6nL90eTWjRiqAkA9QMZFL+hS
iJ+W5xl6StSrAR82yHxRuncIEjbrLTbkubqiYTLBx+8P4t93oJ71f7TkoW8PoGLOrlzseEIS5hwE
H5t6rbJeNMl0KAn4gDNfqHdxJ/bf/1eG59xH9THKDQDFPNTCl4XY38n8ecn0Cn6XU1FGptmvHCVn
126ocMSRkEPf1WV+XcqpsRhKZ3Y7YY2VtW8WrW97jH77Nv46qevoZ9fkwoPxacZDpWQmc40q59m8
jUddE6In+m3wdm2yl1GZHHkBXxzST74uWVCMHb7jGgEWQsFHadSCE1P2rpLMAKMocQnXOpT5XmxX
EcazWeiClpZe1AONVI3iJWXcEv/2SKqFfBsf+RrIKo61PAQo6RttJ46h/tFnLrA0TLLRo45Fyx7/
OZeo4TZL33LXW76YLXJkPgf4/Cm2fEbhzo3O/aHyJwpR2FIQ0hE2O9NHXI9PRsho3CI0vIwtSOpo
eL6QLSjQ4W31bRk0N1bFMNCBM4AOE8egsqA1ePlgeV5LHFYMvb52j9dyLAzNNTVe+mEWjXsocybA
P6Dhkkx/rQQJdOtFKb08oAoAQp5JSWkhnpCuckB6pQ+JWaE36IUM9YSt5AT8IMawfHybSiaOUFkr
kbxHbaaskKYxFOEtgkJIS51vLSLFrIqo+PxrH9Mp5IBReju22/VZ1bJO7C/oaXB7WmK7xUkH4gez
B0Rm39Znf2ZVPfnhXaC24f5Mgz5hwTIQf0jw9fFtlSFyJtKIGKZbObP3oevGUiJvX260ZwbuUa8g
7gu9VC/YSotWcd+t7fPPuc4OCGlBXiRfurD6lCkvYhHGcUy2MmaQqS/3Qt7uLm0d0T2J2hwSw5Gd
57XFsKz7OChhhBOAAi8BHJ77sbJ29ygawZUEVgra/Zfg2kWCPZtHocy/Xr8QkLHsTfUCV27wzPbK
e8OvQGU+iYQlyRvOhMBR8FPAeSd7KLktY2Zck8uR2oVbGgYlB1ZkQODwY0VQ9yoVtG1FClm0X+kA
sqf/Wd6dKd5S+KdqtPqG3jflUCpCnZ21HmF66HOTte/sjsx/BN1ZZ0pyKlN8UcYBjxpt4TnVV1Py
yNr+7toVE1NZNQcHUyHdSrVsqpkyOZDHO89NvtEaOER051NeKYCmqoiKi3VPMcPijYJxF0EU95Dc
P9D1f+Mq50FktuU+Zk4XmedC64aobZroR0EGqQWJ5H/n6vOqcYgCRcHUi8IqUOkVVik+MIr+1mMn
+j5kevhjFwcE0lP/PRHwBxuR3lORX+tc24YinuKQGVGaxlViQASUwzijs1F0aLuV6odw5KyV7P0d
R9VzZrZ+OQebYhMJ+TPcckEasq9fHpPSLKFvZSmqvNoPB1ZbDiyYWUjQxwD+QR7dflBx4tbsjl4z
zMWqITkVYLqxL8bCMj/sqckOVrI9zzPYqXSdWdiSExgQjpPuEEvOEnwHFjbG5U6NHkvwCzodn6KW
PZXqXRQ4+yFHJcS1UbzDvDL8tLmbU/443SzqdrLdfKyidGr84GDpUqHTI9yd7Yeww2lzzJ5x0AWB
NrMLw1OTpiolHhte+xiLUA6BULkb573HacGy6dlIukiOChlu3+A0HtSD58rs9icM9osWWJgqO5fu
b/AV6XIfxIAigNbJDc+anKEDnu4PQpKqh0MTF6lhQSI4ANb4VN4wFOlgL2wXrHf/hv2O+occQFdZ
MhK8QsaFBodEkvLg8HQB+hRQy9DvSMnAe06QaBPPpCfCK2r9MURdgGRAobclWYIuGO+mHPxjYZsc
DP2kQLqvcldp86SMH62qaMrM2rrSfSZGTnb3e+oqNe/Y8u9b4XlMXLUBcZsxequNUv4fyqNnkMhi
eNLmpsINC7pLKcLKfkG24oUvkkrUIire4CX404B6bMIqJ0nWt0nTwPSzMDIiDQe4rPyZt2MgLqZj
vQGgV3MgAi2K8N236bUSm+JyN1rxQok4GdH5H5/TzKiAJdxJwxe5jYxrPGkRynshoqQ7e+nJ7Hii
OQlG+dSU+J7lcmjspib3ScnP8I3ZIILm/kyT9gFudf94VhNvzLwwX8ZWsc4GWchDq33bZKC8IxSx
UjZcTI04Tfj87a3X33+zl2UQOE2r3tAp6Kdiu+CEuBIHSImxrm2mp2nDBDC8GO4C0Qbh3+0hEbzo
vj266l/IWiH6+TRy0pUJCbDWsbmwBJrIYXBKnk58VT+DxsVlILASZ9Qgq2tiufzWoxKNmepDBEF+
MFBqhnJ7xllHIShObOXu77cejP9evL2S87FYDb5BtwixeKiNwmKpAD9RtFaeALmih79LNwA1FfHW
8L+xBISOG0/56J9Fo8CzBQjhYQ8RPjbDO6nujGFkosMA0odN0aQWxVxqomTSUxo2FZack9GQGwji
+F3z/gdxBFMIzbK35kqTJC+8MBQ5xBB1d0v1lVg1xSaxOGDxjdIf2+KV9IPEk9nTm8i0On5L+I7a
LGU4NvX3nttwHfO5qd+1V/tfaVbqBEqGeP8kcO6/LJu1CsFE3PHj860G9iFJQ8S88IoFr51qqOyk
3+WKqXLW2zc6X2BSLa0Y9Y2BdTDeWV0MW3QSJv/zQKL/FwdWXiAL5WsyrX8eSPC1ibWUlL8lha/A
guBAM9Oxv9si2TqQ+y/J4MaxRRqp71PBrPdBU921gPtdyvtl884gW6EI/zcAtqN1fXixa8Kb/AfK
Fxg7cf3MIQ39ZuTNzf5oyyDcXQ6bIvAb90f8a8MF8qDL9xxA4OxXrNqq3yyt1z+A23Vo5AkwL+ZP
Kr6vXV1PbVuiw2fbe/Y4PmwDNQdN5+ylyQrcfZSHLMAN/6BgPv2CjIBUPn5lNR37uxVs0QsC1KDf
hmkw5cI4j3ioqvBBLi1/wue+T4P9RUqifzApEj86xaoonkWhEE5WNqwZCRcHTp0TGqFsO/9VFwG9
Qj0O3D/yhyF42pN6+dFpAEYLJ9RyouCDqdDzQE6pbm4qzMLQVt69GyAOXUlsnUDzSXbx/rbcGGD6
tt70XHB1AHJU5B3FN5YdvMP361dwZzGEeOyujFzedlpfNOFZ41m2AFwrRA990xdq+0PCOkQckplh
ZbpfIvdEn7wgB+W/qL/cZsLp0+pTu2nUHQwmszactokb4vHfJuMTkA2u1emlGiuy5e3go6Tr8Br3
8huaLUyFv+lWq0FpizySInS+g+q5ATh0RFKTp2hVlJ03X3r66nnwUmWCQ4rZ3BHNArlT4RNobPqz
wic3aUyBAeh1vZRvJVU9IWSU1ummYdUT0ePnDbzAvzVqloJ6so308Sh3KofsTpCELwiML/K8N/nL
VRxAQMNK117WdV25n0llpPWbmyavBF3xZSMgOmbyO3ZDFrxv1Tq8zE8BLVL8r95Zn6i+2ZvD5n8H
trMMEwt2I2l8YMd1eXdyE3J6X0XRlUV1vbI92bVK2F38moC+g1WRAUWPrqfvtBW00iYZtX24Hacm
UZLLySUsLgGknDZgYyQ+Iq8zmaPIsf13HuH8eP0AImpMwxoEYxQKiU51JLRYWNeDRG+Y2GT5ZR8c
7uNzQbuugNmHSGDzkx2zJtYdhC8GWR9RW6wRrX+1jb84cOXlgKg4oGgaT+GEjyaLGKCf4Ae2XJAZ
jDr28/ggduLKLPB8s/UFKgTpKYOjGlg5T31zJXD2Npv0PfN1PJ/z9/56Wc05hpWIZX+s4WD7nqrO
p3VCEoxalmmU0COvnm7akHSKSST3Y9en20+kuELigV9c/KjP8pc3IJXtN2CJZfw6u6RhIg2IZZ36
sOSeRih9sPhIJHSVzhFqLfS6ScK5Z9EifyAxwI4NNZ9Ap0FnacE0437TKxIzc5ufqac0drLIdD/T
wtNpXh01OZDkAvEkRRHdLL6gvhSOGwTK36dNnbQh1mTgxhfA6bTIkncOLzN5xI2rQhur37OFz4CR
LL03QzGnnhU8vYyTyUNkblaLgBIREF6Hlso79NZxVbY+6Hgzuc5m43npSRcimkcw431CtOUEV9dR
l5Fh8ceP1erYR7YWMA6JLbc+PVYnGmUqpUHJ3wBDc3eP8UgaiHmFtvhqKD5yDyPZLQmjfNDVjrME
BF3t/2rmFpIE1VPSs9SWL3gC4LFAQF3TiONH2MeV1M9uMAyP3uKKSKNG0Q+l2ruHmPNGBRU48gJq
xFSZ1FtMVATImMUWCY8rhY9oFbasJRPvTkJdmpIS4B70EfpH8DpRcA+kN01EFKydHdCYVL9ckbXH
517xrRL41SxoB+siNrxmzfwGUXYrQiWK8tfu+rtIl/LLLDUFGd1XjDrs2ZnWt1oKBXupuhUC5nWX
Z0FrHPgKbbVU/MWFqUAjob63h11H8ufjPuNh8OI9tYgudjMhap2x8Pxy5XGJ1NO5XE0p2cAN9oHH
lZllJRzaQEtc1+kbOUYGxrsW7apPClxKya3EO3tiZ5dk2OUmnC57cRXlhttpJrX34TW1MZFl5YF9
TysHuVKqSDb/0326zkvQ9gtII7yZWVaDm40bbyIUNpH/hqiKSD8GZFqEMb1mw2cJjA6fYQTwjPV9
ujRG9eSxE78HrbPPxrrnimDS5tLTxg5tIUS4YH/vOq5tkvRoeDBMPoN1Nf/AlRf1CySXYulSlJJT
07SML45oY06LyJZ5Y1obOT4Mo0sFkVDgCk5NlYxhBMGFLXagVy95rikcHOSQObqIG4LaMBLmIH9K
kO5X/efa4S55/jSI8pcCdQSr54jpKvwROACaJ+QDF7xYflvuncepVbNyp0g+NE7EHg8kqZcD9rXy
Sc4lk7Wg+Es/nJaF6oSAEcdKPjj9HMk36K8FSxNg0b3sjS/99MBBnqlAvZU9Ar3A5exlWjwcXqHE
ULhonIGmP5R6qM4O5lFvcrjIGe+nnlxPij7Zb8bqpyaUfkSNrfFIV766azlrQw2WR7vdw90ytAIJ
uRkfHZ7xjTpOahQ3VzkK4aAPyDdLwIhpZDpgercneFumOXZG0TpTRj+SIKrpKlvkhr8RVD+2Dr5m
YXRVbJwxRCQSN9eeKSVb+hNO1PWQjwq6Bg4UsC677zgfWm33VKQu9AeqDZz32EVDvrC4CXLNeq/U
yGNlI5SxmirPUiRSGlsIRJ1JR1XYYboOfrrqyq03UizsJ9K6XpusAgY658kaLvVpbXP0SU++e3fw
RPaWbgPfCJUdgwDCL0641s7PD7dSZhObm3ydwqHYg5XqGDT2zt6Ko5HgcsIMoulPQO/DykNWgjaq
6CZGJodOPS3fPdRSW9I0JIjtLAfsp/X34myYwqMgh53Dvfj2yv+Tsqe6XqTSjj/UqnYJuNIaPNh0
SIMa9fmY81GlriFITcj8xXoGg3wCjPes/GBGiaILQaTcrrj3+/T59zXI4siPoQ4rtExCDPq5QQkX
bq45MDdHkPjqUWIWLKiUjlFHkP3hDdcn0Ca4dX/rrju8EwJM7nP5YE6Xpti1PYj6ef3b86dZqYJO
y4Pf9N1CW3LA84OREQclEoHBLzktmh9pmTJOC9IY7Sh3vzawn3LgGNpLL7wouSvUdJdVFOqk4EH8
sJgnZGv9rHtZ217AmuxUF9mHzejeJDrKhb1hRzrQqk83/uhtg6rNv5AVVukkaCHyekNwJqmDDXCS
98NhrBnrnsvOf8zSZejp3xmAB8nKyIgo2YSxlty2voH7dPeQuf4P5gpnZZhNQ+oEJe84zz0sBdaw
Cn8xGn5VIXbfpR7QfMpHS9z2YPXaLqTQAruGglzyLHPyZLJA+khIadPp4J6yQX2cUa7w+Q67DMOR
qEcbhiKBhyvaEeR/E9O3deQ3OUJlO66/vd/lFH2tS/mPeSZXEV+0rSU7m4djft2VMcK19ZdzI+zV
7ZtV98ZttSKizGn8VIYkKhI2dja7J6gh2TC1wuiBzM112nbtSjO61VUWDfaz3GBvwbSJlgJjJSPF
ccjYRX04ahpew6L83DQN6UnSdfINgO239pfWugb434gZgeKQz+KtWsS6dDhMCnpubNQwsz3IONh/
RjEzP+fJf7cWEwIMRBcHkymRgIp8bs3rrQVCr0o0fZJucuFIHMSI2OzisJjUwO7tuyZ+CjyH5d9t
f5TNod5dnsJhhpoF2cDjk1nwWpncGH1Br5E2MlQxOTycGhIMDlc0EW3XZ5tFuSBSuGuOuq1B12Se
RuuVfN/b5XZIP0ZKWIkgizQR0NsDrl1f/S7ThrkmeImIQIJIdYhHsfMyTYNO6+MhbxU6cszQM8lj
K0sGE0e0wY6K/dTqugRvTgNhID2Q71uedLIxquuNXD4WCY3wWpis0l0MpKR4e00DYM3A5okEdBG3
iAi/jF0QiuCPxrvWOHKLlJjf1aSTlpnXVGatfxKFpII3jc9hDCFqqlQCsbYNUJxNEgtYm6l11qRC
LM/Ai8EuC34hgYFUC0TuO9QFAmGrZAXJTBY7T/h8GIQpUy0hD7877fV74O8XTMUqLV5EiGexqTdq
JMpXjIiGpHlttNL+7KqUl4pNJhbbCZO+xqc/r5aPWIZfMsSNCHu1gAu5y7tRJ4PwRs3HYke1LId1
s/MmC/Q0lkRz+Rluwj4G23xBF/mDXjOKLIHRg2am/Kwi30OsgHPeVq5Al7cZ+nLoo1X0B2H6I5IH
E0QsJuUsDgKtI3abORvfCT6AF0AOrkA42CYsPbxQqQvIYT20liJV3dAnd3UieBOwCsAmw6vNxtSQ
j/sM5YZm6gBQFmwq2/GtBtiRMCIV+/vGw9eRKE4m+d3ymReO2HE1LH3Ql67hEpo7n/zNnqKhaiB5
OFlhA1jdMNnAottahNJpWEKpE/mIjPRyjuecb2dCOjKdKorQi+Nj8MnFONblPYFYY9Y6Z7Uh+7vU
r1LsL+NdOfZCypBIe69KFx4I/1ftqCVyYCGC3RR8BU81IWoztfQTufE8tRTPhyghKfy2CTdEbfWT
gCSLKdxSA80GehtZULxri1Bsd4AZ+1PIEa9/X5wkC0jZW8qqCkpddKtU+Ckcx8+EYejgjnC7tONx
4XyqTjEGGWTzVyy6uYm8vXkj5xyx93Xw0swjhxp6caEv/NnY3JaC01iWSEUe3y05S/3UqR3g6Ato
vDA/zdWpje5hYx4PSyl5qb2WkPP6UzWVvtwCEgCQixQfdGQUlvemJQYHvka2W5m565mRUjirrsFY
M8BTa2d+u3LYPPWvHbf0Pik1LN4JG9pE2cbbjIDZY1BlpruFIwFiHCtw8nd9cfrK0rHbU2AXYZBR
Z+oFTy7z5v1BAI+QqBeIGCj3xigJdKGjQh9nai44pP3Zp/pjo88DtypXS62+uhY2Xe+LvWks3jo5
Sn1nKGqpfEG5qD5IS+2HHmpyDzEomCXkadVtiZxBCehBpUD7Sj47U4f8hhGx2EZFKYvJD3uWp34e
sh54vdrpKizz7S6v8pu3RiNcUusu2qMUnYEXY67Rx+vPQVK21NpnhnYC1UXKWRuLx+fy0c9uR8sW
6faKI7t6jQeorr0jJSuOLl7mzmTtCT0Nzdzun0VeYyvaZkvie2XfZ2g1exK2JeQaZtB9rJ/HqEVA
wBR1y/bC0WSldN/7VXbXGKgzDM/t2DjOl0pcbI8bEHTVhY2tifl6WFsRR6yL5VFlX/ScjudmNQy8
byTo42/BAmd66ZxDGudHaNwhx59ieNEHWweKNSMiYbE7FMPtuEWcpyCr5/80av9Q90wS9skKaBBA
z8tupZqvnXqFv/X/nvVmRmBWtNiGFj4srsifA/W7DN2KyADAyPAzWxG8Kyf7jdhS9CmJlMVd3Je2
x23cpEdl6pCNagZwLYpUQu3Qf+Qv7xzAv9zAukVhKxMM/cSnbOjiXbPn2bnQ4to/amTguIrSuz+B
DkWxiPmaf+Wz4/b/mYcFwJOqKDsKN8cTPxoyzAlVq0F90QOSNNKGtZGH68wFz4F/P3K4yYBiP6Rz
gjYeE8nANeXD7KcWD/kC5ejLU/3dv2rm4g0TCi2hxz0t86Ipie/1nB44NpYJ3mPSffS4N4qZ0NDi
g/Ftbihyr8xfE60w2OFIVkFyO+++bXdLDNC5F/LdakiFPB+0UNNdtq+7W3PPsyZR5oREX8qJXPM9
lATBG2f9TIWoyquWk41BTvLV2O3BzNLSTUvzpUiwy4fvaap6BhgwsntcBgzpWGo7xfDdkqNiSIHq
IIdZu7Vzsv2BOP0LT/8p0apo0dut9xDuD1ugHBhVc4ETU4jYN3RerzZNhvPYxdlew7vwYP7sQ97p
FX4BjA5gjIlw/3/CZzTA+X78XMwQw4eyRee6h2DpS9RvQDFjFFC+WcrfSztu6kPSmpv+ly1Nsmjb
kFoVYTCnxTf/ThDZGxF1C0nJC3KixfThwHtM6VJ9lRJ1IDaiWoHJuYRAwQ4+hAuHtA4/gET46la9
VJrhwKI6XNdAf97xLwswVcAQ4OuELV2z6Q3V80UPNIaRzH8ucwwCAdd1S6IwbzWRhKrx2fuHSiyT
waI8JicMuFoiKkwqSTZKxDgs9LP4p8VTyECIT6iLjd68S0N4Epx5yrpM1NPcbCtF7rlwscbEjY9C
bna3vH2eq/hmJTue2YeRX2tbjqw9CW7HINF6eOTWAEaq8JhXbB7AUlzbX3hx/VCcIaLVm/KuZCtE
eowWTYhIIgVF9/HsxQFKlK/IvkXz/fPqsfsLrKeUA3ibsu3usyL9TsJcywDk6+PO4gamYX2mF0kS
6fa5M5XebbC3EnJeJXZx4JHFmx6PuMTiWBqUSp3S36prdHix226KxKn0tOnfWgmnxZgKxroihHub
pUjuTKvexKOpFsEffzUqvb8XlOQgNp9y4ptijQGpAeWUQ1jKcOKNeGaNiIAiFEFf5s+j5GoQMGvV
3rGHVzxVbMwyg/3B6wqM3jzCR4uywhI+popdoz3IvKRBnqGb/2MLZdr8eqBaT2qLbasgpBm3S8yc
IlXWJkaTBKcFYdoO3B5FZnwieyHOdAf2lP07ViipO+ZgjMDvZ7tXCsI/aVbvTfv6WdR7U5susdby
Y3AGR+Cxf/ECTksA3rtaLuHmuZY8ktz/ISoESJlXFzQZHNSTupVa3VrP917sS2lNgdLavVRflgvy
B7jVUzAdkQO0m2N21RJnEKuIik4zClulG/gqr2smdtiqW4aZ/6ooFdFtn3daaUl4g9B6Dor0NUK+
DJ+BUIS/3R+96pCD3XPtLTEUEmf84aIRNH9tAbnCzZJ3d4cZsvlGOtp8zte3W7SiHoPk2PiUQdPX
vJRf1hwMLsMtXJnmjTJkKol5yMLpSYttwFxGRjm6RocyepyX2C0OXF7tU4qZ9zBFONpp6WcjFTgD
INBmHOaRlIQdFjZH+Fom2Uiqu26K1rAYPA88H0hTQzQJq2P9gT4ZQ0cIIRUh5jJRrMRf4T+P2ssB
pkWhrnyqu9u/LIfuHStoUL8PeOw/r3JBRi94UPd0Tm3Q24jqEFtYiZMZR/EUy+MQvoVuEIgv3ri9
p7Bq9SnwYithGMmVnfKCRiyiEdjR0VyU2tTYzM5j1N0j5VZZZfSFFF8uRMm2lJnCiCl/3ERe1bv2
yyKTu6q/jIv/e4+ObTfKtw8g2Q/Z2v6lMsROWIVPoGk4Qixrh1P/RLp7/AuBd8znTd+CmA3M7HW9
TbjceDuI8a7L1aphHTl9vwnyzZrKTV6U6PZYbOKejwQGd/TRSpmGhcS7BGqTn08+anOlYtl55eIJ
ImdtCoB19u5doilYJFvP2X1rm2BqPogIDPtVQJP5rpBZUtGwXYjD9/9GinOYhEumixdM/lANFgyu
2Hu96bgYiVlWGiANYHk5PvgUgXqDDOVcJNcrLlilBkgtaXVsgtNsLW+HhazmGuZ2epK7BziWuWz0
HIdNMnJ+/+5UfSw86DmO6Wig5bD1U4lVdQj3JbcTVtdK6r7oZ/GgQJcDYO/j/parC6Xy0F9QzqQ6
AFlOYp0X9oYkw0BKft9Ny75W25656Yd0Gr/5d5jGubcYoGtF6EnDQqrkQWWC51vzPWpwGiF1PIRw
R6fF5DdJxjaQ5LINY3h40QjEjxLG631yvk+SUs0Rl/eZQIF1CKPreScj6m7temv41I7HByz7HzRa
H1bLQylFZEMFLgRVOrqc9BpmRj1h3+ToadRJHMFIlitflfZfnx5EvX4YXEBuWF+wFuO7Li22hLv/
/1+pbGp2qumU6LFw0Xl0+jmStRYcesLhbV1sYiZ0sNx2xkgBPsXcZ9bWBMr3RkFs5Z2xLZ9D8210
NneaXGr4zqf3xiybD3fPa8WZG8A8R578PQLuqp3FwrWVIwuzx59Y7zRbpiEiA7nnPw3jCxjK5XAo
ENCiQ9ScS/97Cvv+B8E1MnV1CU7KgzebyPehw2dKoVcvxsV57PCxUeRWcrirc7EqSlgLud+kM3Dv
L4fUh8879DLiywVYTHq31WeIcn1pc2ruPrFHccIytMZYdNBCeYkmkjYL6JrW36sXTCXhce2oQVCa
Q0ef9ljgAV3C/DcImYdsv8izUpgntwwQrHybbCP6RmvXnwgmDGL4ulx7CPjx4MKDuDBiX2aUSwuJ
SRwTxLtNcJak5U0sb8ZEOKngQ1XOmSq1CJKfGrg9chIpccWxoj0bm3LMTo5i7aWJo7LvZ5eoQ6hu
qH7eZUsgBsz5vTib/ElFvP3T8nRw/3Px91tpMGm0u5YRRIMuBAzQdTtsstNK3T15JD/LD8l0YoWu
jiEYwZ9BO9QRfFYHshg5yDw3ePN/DOpoW4YOB4n5YaQz3iHaRdXI5x8GBa1cEEqOmdCVk4iMEQQG
WoTc1R7VYh6mh2lOwUXVH2usEKk4WJeUQm0rn2jrZ9LEkFZfF0nmjuVmPNXR1sL72dY2AGXSnLSI
ewb6VMlEB5TX/ToShvof15xW47/MSoMKaWGrrM6DgS0wC1GWkXXTykFYb1CKvf8OoP7g4J62DY1L
BexODCSziypQxcL4tnOiGNb4zRILS0c1jUHpYKgpdtecyc7BapKxyfkm1/o3LnUkoPG1zWs/0jIg
dEooVVB+pyMiK0rlnObLDrrO4VlBCZ/Y6QOFGdct5L5DHprXlhtXJU95bUOGoGFI61DMzvFzNw2u
HaAPj/SuDUFLVqau9bGf46zQI+pkZFBCtm3BntRR74Y25J9EcZgNEJaNCIt+myM6Z4SDquMMsjpf
EYzE9fgYrc9DdzWfLJXmQaoYdZExG3o/lPE651X9yWosU7NpR2O4wXRisqdUkpq7jEjwdN7AvXAr
dClipJrm0mDFmewXyFeCzTgH8ErN6uRnyMJKKSWVAeQdnhlRR48KDPcREX9USe/El9AigJPdHoAC
6zd6JCz36tw2/C4xs91I0YUuK/pAizzPcwib2GA3sag+VVlEDnzQPp/D8xLQO45FzQ7FkFZQ1J5h
xj29E3fW6iyb96X4XXMAhnwx49Nq+rzaRbNBK4JomzKFcT4VaX3ur4KczxAU3nI4gO3HX+Q68659
6vL6KOe9fY87Kl0d1vTDqmuzr6oXkNRRAM2DqHtzyGZm+nh3xpQZZ5OejS/gat9i7y+lbN/qCLap
8JCLc7ZuX8Oo5uDt+z/3cPQ8Xsueo4iJyTe5d5mpqbhfzZZNEcAJiDixdpkhg+ytdl7EmTzt47eW
ZBdPLqLH2clMsPgVU/WbCFIh0mq9avNb3CooPMaKceVl4HUqba6Ra74tIJ+4mtcdTjj1xv/HBJfp
Oyb9HdUT1Y63cghCLAntdmukXE3R6GNrwBZJnudXzUm0+NzsJeoEOBozBNaUpEf9GBaECw9rW2Lz
eR63zCNfzfJz4+b6CRODlJaFSzyk1xJxJ0C//DKk4VNWa5oiqp16r5R8ssy2iSdK57lF4mUNBu81
v64SVIUCWTa9SsvJ7424SN9TXPPOAKusX6MZUq+mbACJ/1GLzaxt8NwFjKMMIJwalVA+ueV5bWyP
qL4d07cmqLDfVTLdbI6yDBep3Laub6bl7GIEmuBqaPg+nhNeTHQQJu4aXM/DDjFlGsii2/mXf6X3
IgBX6HQVbbGwF1kRWEvoqwHdr4PRK6v9NUGL3UkSAoqiDB6Pa+ozKhMwvBbx8o9DSh55W6AbWLvA
lEM+ZSASsec6sF63qgdTxY0B96K2xi94OoerBG5XNRbpvGC+K4cmlZKo+nhTFqh+RJZjTOhx9V0m
US88iL2q4hlEVfiD7ifwIeeqyMqG9B20n37JYmx5T3RjDILa8+cs/IkplA1HqTx5sTth/hzcm/0S
T3KERZLRiE/25EDSoGTYz6EAS74TgMIFXhvM+wUhFHcJid/rz5QwGylvBP4MCyOfJ87FE3eXPnen
0TKeax592AY8rDsziYbQq9qjc9WzxCVYJAp/aMZlSdvhxUeBMlGq36gY0oRO8Wtjr0UYk1gXROHV
ApobP+sUBsyDqCwgk2PdsF1He/VGudO5kecUFL3+Hb7WTBrK9265UZryzuYeketsMTate9GsgMWu
0pIk0xI7248gbnviPb+96xaGg/Hqrcf6KvkodTaPtanJp/YeTM80Uzu5bsX5XW1/YJTOrTAuNNN8
IWQ0CKsvUgjARxfgVWyy4aoZe0WGnvF/Izin+8xapYm+rThxBaRPOV2wiU5EmyYCz1BLBLkaqR/y
jgMHd+n48bkyWo3T8zTXGZEv7kB6HebBBYa4bY0BoIEYGuEWMpvt0R82HCaudRcllTYucHZeLs29
xJffzkKF1XUuFuRl8/9FGU6zUBzBmB6ikOPSdvY+rCUEbz0TneDjucZvP3F8bwPNKcv+LQx6s5U1
o/U9jrV6Y6yLKP2wSZuipxOx4xftq8EdenJRDra9UfDfcvnJvYYFvBetIeCJnrCPQ+KDiGMqJlqA
x9quH/jH3wshdKtgw0SIEccv29/vizr+kBug1QBd7QEWuKc9Z4k0Kjw/nZVj8FxRJB6V3F55hAay
23LqpQq/CHL6X3pa2TC3YeDjAq5C5SUFx9kaa+yzbblw8pjWtf/thRo7+2LrIx1nyohDoj5wAhjh
vseCyymB0dAE9+jAOdiczErafOJjpYMY09AvF//Z/nHKiT/+8I4heE1QDD3X7ObJ8YDrxmNx78JM
FoXb70LyM4HRKW5QnO7pm+p1OgOTBLrL5aQb3k26jjYfpMw5SSsCbdIu+CUylQdMv9xVfNgHYVRF
a8GxsL2JdIdNTgld4As4ynG6pQNdqfh37hoYBGeJCwQ2M2peFqTc/lZY1nOvnZmWs9oqPfRwfylO
68lYXI6zsMldVyOXn/P8cEz2gh6q/9/K0/xRy2V/bfWIR6bE2IHyRHvp/dpZTV1PcRudhNdUsVc+
dS7wk2yZP/5PiNA1hoDrWJ4TY8h97HBGkHVHGyPP2e6zH1zo0W6igOkNqfqLnl071PSmbL1L5oq4
xYbEPuOGmmaH5CxD6YXxZ6FA/C3J8taOHpvaFUa+yK+fHBwwCJEOHEDx+JWiJ8lEZZUxMW3Zf7hU
UItDvGqDOTl2pWIascPL55d6T+oNmZl7R0uEwX4oM/tF2lt6EoDtYRy5K7mC8klndicxbiOTScd2
6vcc7ixfnERR32ddefpjFrCHUyOGpqF8L68fYgUpOrhpNkrk21Pg4ERcDl3BlE5kPNakZipWq48B
CFRAymH8SB0BuwR+9GiV9lsuH1gZePXw9pSG5e4bgq+SGdURoVT8Zv3lVKHEi2u2tlvsyRTuU1u+
lW7w7HoLeHoKWLarO2bf1hBbU4yhRxd/Brn8KbDxDncpp0+ztnL1vzhmCPbk8r5gnAXG1X1+pqPX
DjMdm6pbZ2OWCg+6YQrTrP8HMRlOt1vcN+1dNS/PD8mM3SRy7Z5tpKk927D0fuvgjB971m+TZJiy
q0+Dk4/8b3oWyOMbsQECPIdwcFwVhml6M19jJI55Hz81+PL6b22HPiRhTKOTKGkL29FO9u3w3Q93
GDNzY0MYF0xnRhHE0XQQoQxbVXHw+QwwpfpQAdAHOAjN8di9bFRka/h5HJ2/jvQzFIBbwdgwpUqw
AF7Fe27GOqyzvKt6812lnhDIVSmUDDfz0n7sxxjIiuNKb/Y5aNAYJbjgdS93VA+/6kWrH9G7ZZ38
YRT1+sUkfUPePAfvq+69iFRhFKPrQuty102V2GQFUJ+sv/6GgxdEEaca6CnF9L20XXhiauz3eGIL
6MBWR8PNd/XYGCwJRXCAiR+8EMhTrstd2bCK3uzG0gGh0mLos6teDMK+opp4nUbQzZ6d53EUqic0
Vx5fuJfT4Or+HDSNo9ZgCIq89e2GkJmCTuJCz8KKx+DMZCXDqbQPsjP8Q8X0+Za8LCqFJqfs/KKG
qU+qnrKTRJMCuagThlItwWxIT/rL4V3VB+1sRnkyT5YFIhdlHzWT0SrrnOWjWMIZpK0e1zgUwlMc
RHcrSFTiqOddVhQ+4h+ZfQcpy304eS2iQO+qXhr8U3667M7PUGuZJuzPQFxuvFPFrkxBCjEmJtYb
wGJ/7RNjR6JVrfiYW4gVRs1dwihiZHKQ2lRWAw7Pag4QeOCpgfR3D0hcNDFNwAANKq+Pmu1+ys1y
F9cMbspK89JdPo6kWC6gixHAI6UgbBC/PVZUvLg0wZ/ymPYOTzzWy1Gj7NNfILKd2yRUBTaqAS97
uthHbswczXZis3c4fXo15XVpfY2/vamH5P3JUXTQattbVEGzAkmMtiZYIE4TCKuOYvw4I4cxAbRw
iW/b5zSGOKzWVCByY0WmAB3CM+SLkEaEM+RIPLw/tqyFsYsARyTHX8kuWu/fWkDVCMka7VaOus/R
YEY/vFcUEgDAaMMOU1dHwsjngpT2EmP4yQx8fiizRFL3yg0t/5217gstlwsFK4CF14Lc2v7mMWDF
Go8WwyhHCWiP+2cjxSoWDXDDvL4kHo46M5nY1qsSi5JXDa/s9YP+8++Xo0rhjXWBpuqfk80xRhpb
cK/UO+Ksky5YOxZtkJl+Qp34jXyakoAYe1c4ugMntV5Ci/ypzo3eIQV3yeiCI8PwFIUDS6AwRZUD
EJMDCzsjh4L37H3L/mVa2cPCUwPmU7nf8mBpbzcHZQCQcGZVmqxRgXEkHmdvLIAiw9vVqnmLJgev
d0hPcIFlrJw7xbGnYX8BSb1BPfN/FJyWBjY5uJZ0CxF1XK+2klFS6ElkO/Ynq8wYHN5b0a+O9mgx
Tcm6jY7SNywPI8aV7jFMMQSNg34+83nYOoc6OgZeZ283UsRIkOG5gHJ3Cz+a1iCX7OphcC/OnNIT
H4DEfokQ/Uy3upe7R6avUdJmUKz/PB0frGlzT7FS0f4p2Vd6AX240EUF/BnlVsSGBEYujuXqsZ27
FfYFa8c7aIY2DPAJXlXwNBDepm8AwAHv/FAP6kKZund3FiO7vJzcG+HZXJkAn+nPy8s6my5lrro6
oT25pkYg7WDUPFnGMWEK/SsDNb33srzdASiS4wb8dA/NHriW/uuHYTM70VTnq0lFeJSqqysC/+XJ
PepvfHfzcsD8c+Yz+Vlbb4rZNVFj6yynl+cqQ8+rCU+yHAt2FTEIL3P5ZZgSHH3BeaaZ1Iw40Gtf
9ON55y2DDPBNXUPHRIjQX2gA0020CoV/0P76DVHlzBSW9GOHwlMy3kofk12TryQ4ipL3ADLCAKMJ
RGCEhg0IIe6VKCgiZJGDe+9LcrkhK71ambjUiKz8Oo2u7zSnUikZcPtGjlmptZ1U94u9u5oeoIS8
mYFeOT8VuZo7FziVw8bbCRlgbiBUXMPIzmeRrPt+UebtDK4ZhOm3Hxu3d1WxiS3ZI5d//5yk0Dsw
YIofzfDeqwc/4tLRF0jmmNaMPgKRMH3Dzxqrki5Mn1Uv67KVx06pGpp+giHMnMajN3HRq7IBs4w0
U0UGk9EKhrV/ms4pzDN2xqwjdMC26JHjiRML6Wi9ucPiePD2580MpptVjV/Fa+qzo6BjXxH54ke4
TelfMIQzfsbX4at6T5L/7xst4SAb/D9LKGUXnmDPjducJZfzc9vWJHduAESn3yy0u0RyJGlUPhWK
KxxUF0fJihX2wUq7atoDBHkq02ZEXmzGhVeTMHgyXQwy2faRNYZOFFJhpdWmoaCe2Bne3xoXbp/i
VKCE+4OA8WaCZ1vZJxzKsesIddfcJN+mo+vngLxT28rqKA0/0wi4O9oFwMthAAdnvDpDoQTMKn2U
mzcVeXZOvkX/OxCEE5BoXnM0UIzIhdxgmvXLhwv+6nYw9UUPJCRk2JPxRKNMf1ZhVIV+jK8D8vsF
p0cYTM3Ys7SLHkOTowKq1SUMjG9hIqhpvc2uUG88bnfHnitpiDpKLX1LPTsvt5mnNQyKsvsqp7xX
fQJHnRL9Hh5TLLMfMNYKozaf13x/wyxOK6C4PNc3j14khAbE0MsEaeOd6Akin/0WzKQva/fayg09
xwctj3zX9U0JE2OPcknQzBgAOziV18UmuQGf28eBi3UlFNC1iRRxY5AZymYgJPdtUpjCRGWVxLSq
zm+8rrAQtVpN2iRFSjiicUmwesNKul5mgKN85zQT4ybuSxY/YV65yUDUKrt9rQ0oSM83YNKAwz4g
k8fEj+ajLtAFG1tUSmvf9pLka3T7JDX5s43WucuxH54CwMwoFeVcCvUSF2jrgy4/2ijPLDj02zy9
7G7v/x7dmA/vfHEqFV5wY5NSy0mqiOP6w2Tjp3Em2RRZmTwjnS1NRAtjCc+erUC85kl+Y6bcyOkS
rUpvqxLCbdTD939hvjMaEbUStq/QipFuLYNy6ueLzoA3GJaZDuxhWqkXfhG03GWA+DTneG2ejZ9c
aJd/BpXQ1AXIpKZPCdD3/0PASBWhL/9iWjzsrLlKLUXOHwwYGp9jVwQdpnUxt/OZZOROagOJkSvI
gC0AB7vDy0oJbOAyLU9q5szDwpwUxE+juwvsfhPcUYD/2+DE3M0JT+lBdPz5Hr/GLcI6YvGKbWRH
cqC+1BufBITt1xf53l9Gat9EAHOE6SC8fs73PQIh1CztLB6sWePI8SQueHT/eQc3GK1r0hIkapDd
fsnpdx380kSlqvPIUFQ88K4uJa5cq5mF5ko1GmcL37GqvWbRIR4Mgc2LRVcefm+Covy1fNLhHNyE
6BfwP7XpSgLB8G00vj7yEdJMOsS8eamHWleZ+VEKsa2vwujivWECVfWXscgTEv1YR0i+fUyygZbD
wak8TPJ77qh+He6m9SIeopmiVfzhsq94Il+5XLRJ+FyzT5cpXVh9qlJsKP/5R4VTOyjKYArnjYqL
w54E0gzITxnKteG9xajTA3ybx0rzfYz3Zs2a6yIlbgXyHHWbAaIAFI9rd4oGEGkj8gydouFxxWnp
8zPpZymmzBs9srywjtPm9nvSUIUwuh+KSOUh892xlKBuiDD9sWvq6xghNmkUNjfYqB3LwjKaowpb
2CC+Ojl/UPUBg1bGE7wAoARlgWzxAy8lH7Vuzz8DI2OiQbRcbhUEuIHK5ZsRVvN+jtqR09dIczpC
I2G5PCOBGzs8tkkKN7KLZyk9njGQYEai05mGeeVALc5RCitWHK439O1xsMQkrEb/Yc0l1y0BzME4
W8ojtqyUHb6dkJIMxyXhLBpa2yb+9uleLj7r4I/5fVS+vb8AtVsJn2ATSxH39BpCdmF7TpL9AyeC
wck6ITyud04xPD9wOW58nGh/QYG6nhpKG4jgun90fRJBl7Ew/MlVWSsu27Es64RmuAPUPRChjzY5
B6qB6Yuw+yqieuu2fefUOn1nmXUmtrQDNk+2L7vlDVnRyfyKhXibTWTpUEINHq+/LTXK1CRn5AAI
t+gK/fVkF35i9ePEwuO0i3E/oeuSeoJZA0n1HCX3CwjaAk4RNVw9thAaLdJClpe6YazeFKcfmfJW
5y2ooeYuvk+e8/Qtp166pdFRRhh08k4a+HZBBxt9+dMEL1Cpy/rKi/2TPyK0E+t/N8uwIKuQOBfg
ceVdLUGuE/xr3NNTSxhtOyoI5uNWGm6LUW+1prSvhc9Z+PDKUDTqCUlFzPh/f5ZoytMiN+iFJEeB
BX+trBlKz18cTqdyCDy1fnfRczl8ByS16LhZuML7ScrNuMxwNTpD0jRQERlyiSNAas14qi9VoB7h
WL0PPuhPaO8tpkmEu2UELGX962+6gl5GgUJNOoMpM61VFQGsU2cLQhbY3VHKmeWztRHK6dQVFO+J
8Efqmo4YYcLmoVc+CpfatH13n1CRlRN38YwOCtVynHJtLHMkFYehQqp8xCN85j0PhHOfC0nyNocB
3eO5Yd7x4aXiazWtnITIHWLAloQvmfIbCee3lVBBqp47RVt890J4btrSeCaMuxwAOlaFa2FUN2lv
eeMP6KBMamJAkoHmp7k8yO54jw5xVM8G08YuflGjTk3pfY5XaOJlUYDicZu1zJGbZAJi4DNAUvie
38JRGHuA4Qw/DKsv7zyCqdqZ8kG/7g+uot5F1Yl2e1ZqPJCLO7Ye5p+huIo/HtTgKG337LsuUi1K
Q1EfPccNrU8A8+857g7y/1Z3B2fvvgFwsb47UYggXBSs3/7x117G55V+BFtJJjAxdPwXU2pySaaY
FmLtvUZykEqno9p9O9Ti4UstJ5hPuww2/I1DPjnsnqDWRo+yqmSdO5u8rN9BCDMiE1hSkRxrUVxZ
Zjg/DaVafHrRZ7NoD01FltRqdDwzf2zfr1LfpxdLMNQQUf3xIau5I8j2ogLXJE+ieqjj1q2LLUbh
j3lG8BdmOjuej7K2WAlsaP991kgDLszaaCR7lEvqXhhHhChUy6Cdc0zT34GnuuTOtSUqdx/8Cki5
VC/AksC8mkIil1jGjOxEW4ojp7F100zPsFRczczHcTdt/0ZrmR5GjpjasYHn5taDMHzR5t+rpaa7
VIUpR53UqkRJ5WeuNj+PtmfCPlz7xGMMelbSN/ehQDM4Tgx7wvTbm2RxLJw7KtBsVrVJYbrABTDd
n5rf7eFEmIAi68iCbZJLZkNXWL20RVDjN2ZoQ9LI/mE6U8bSPSMHOhnklJYpxdGjqnrMy4sFAeoR
aT2ZGjmaTTvXclFGP9u/I2XDs2zbanDagaHyUx8ISh+FuE5bI/CQFzhl46dnvFDG13YOoJNUntNw
pQXVCifrGsKJv8KEmsZRqHntk10yqAOAks4bDqLNURMDxjjopQ/JskUWAQmi5ZhtBZvfSrayXYKn
T5Kd/is3V0yimKCU1YOpGQfG4PG7cq2slK8VLcvaLu40Kn0eFA0QR4DA/tDj1UCtEw1G4+HS0I1J
xQMTvKJQR2V6VpHKC59zCQHCO1uVGZ0hYKDJYsEiVPPfetnOGCmKKlFhxr1jYxL5d0BIMB4FY56U
vUBp+Wur/Zhwrv7XKUmnOvQHjnYiGvhcQANZ61zlFsjCg5eewJWbnGFDmkCemWKtPadQz2nqVFWh
RWiYPbaYg46KxG8+fpchPfbJLdEEu5Eo6iEQQF0xKm0cFSzBTCFZg4UzGSVKMZXndLD2xeR4/lLL
v7vAXd8tgcJrRn5nNGguCcPEZ2UkteZBB8cB+MkyKDF+9ReZS7mlGyPngpVcpWZef5XH3KCYRG3U
MQDbXRNUCcF+93ORPo8hL5IawuIqFRuX2DsWGawRQvlZUeGzZtAktOvDS1+Ell9YiZohF117HiHc
cTFVJAR14Mmu19Yy1VmPp9b6RLz84YnsH3hZ+bCXchDTitNsdMPL6y+LmnJ67vq4GYxkR0Lw2g2H
Evekr3F26YkrCNJzKxucDkAMstjTqMfXdd6kNboZ2y1crWAxWZLDJ1B0KRi6hcNq/ZALd7g1J+OW
WXPCb30y+DtcTD7Dm5Ir4bf4A0TcIN+u/SDFvN/xHXocpT8l1klBBFtDXG5vdYwB1RpzEQNkJLLw
IxaV73YyOz4wRs9td4c6nkU2cDv7EY9WuoDdI40ToI8lLu9UxBH7l2UzUR6FglA4s+KNR8GBxalB
ptBAH1eF3EBLywXEBn+DvvrpjL/zQa2JAswT6zjRgJ76eCtnQhsz4wcgEvBlk6DGfMoDRCWPExmU
9fOwQe7tBvw5fxFWLiI3y2Y4qJvXNjmmFDjjPbLDH7FkR6qGpE05o/C5wsJyYypCstW6KmntTCQ7
V4PMRO7UrZFysUUgSnfwn3t/L1Y2K9KaRVgcICAhYRTM3qWblaUrwI1S1Waq4gSiN0NbtjNk+l18
Q5IPE9KMJSMpfBCF3ksM7PtAiXwvgMoCgusc3AxNeFGDTVzamEcQgwsRFRlCzq43hAcJysHmKPkZ
MvckmnbTUZghzsSbgO5KWfI3ZuXKHOD6L4dQ4uImnnkEY1GZ8HVuB+92nGCCzrxULPaHGafkEpaX
fn8uvto5KviClSTQD4VFwFl3pfNHYiMYpvpezdRO9lFE8Oaec3eDL65yeefAtugLih1bibNpykcq
/UmFeSqgHAD8EL64RT3e3EnOL4fHTVAhgyU7hhto2CdUoca8B8ZM11H7cOnGKhWMG9cVqtjWBLDg
CSFW1dCNvrY78OGcypI8/BaB4HdYrykb9fJwvh/STyMLubHDaTyTFJjrEAKnPbvxpgv5asUxWtPi
RH8ntfeOjnmkK7Roil5Ie8qRqIIJjoKJ1KFa+MUWZS7bkaBpLsw7jwPlKAxVPUhUzfLAjSA9zsd8
S2m5Dw1+R813O+WAaDzqub6zO+ot76jVOLSBHZGx5qrEwJwFbwf0Dk6a+T26KEJ1FPV9nSuBbbZV
W1FixFkv+WQWvhjIQFnIDSj8Ur/sX48+G4PQlbbl8oYa1hhsWTIfIpxFATSiYv5iyI1x7btMQhQc
7H8c/eXwVOowIp8bAFDCx873P4nIkXpa5N7bhA46915RrwjMTqWcMreVFPU6iYIVO4y9z87wWlik
/VA3FbrWv3NRhVHPPe9j4CC0ylBJNd3/+7DmoX5bmX2ch1gwY0cCZipGbagAAIDXHpsE8SstHAdn
k30q/x7kImE42HdA1dbmfQ+mHaoUvDte4jkKD3ekoNWVAsjGXCFsV00rREq8y7nEH+jCfI5owna1
rymupeMOGV/ttXnaczzTUj0dX49xHYAFYQ4GlPDZBfM2H0n6n3sFOwXHQNtOPsjaxkt/PGWZg9v5
AAYSMAx31q6/asZ1BDoSsfjRf0u4UGhpVYl7VrjUrBvYSTQQoMyY07Pz3z+9tTpiJ6VnAEnUuTvj
bso2Q9y2L3Q9qNCCjxvtOMdHB1OdM90c62xaWYnvn+v0C+NjqKP7EBLhaSsnJPmRz/6cDJHUcrGf
AN+Y1td7SGwnePjHRkCCsuBWSk3KDkk+WVs3GKuzSVl4FMTdmQ2kUSiBEqH0P7kOIMdzP04b9e66
xKxBXgpkPlclNc1w/MRYisMhqs4ErKHFY+Wx7LmvncaFgOjlJvaNF8BkSavZcWLvHD3GvzpYnzth
PMoemn7iviWHPeklu110Qi1AcE7o1Y1rVEB5gIAOl1sGG/6yt0LRqttFGAGnx/HHC2lvMIsHh0S/
aDrOu7aUiSiDfNg9EvRJZHB6bdLD6sTXq0YL6OXu5BHc2QnDu5rwjZwl/4xIB4aMEaVDfZK4g+1R
4D2rzFdHH5k+Ytaos0AL+RqzZ6Q0BUoVrPnLnFfpMzar9eqwfqTvlo0v4zRUDcMR9yqbZh6b/Z3E
8cGZYOe/eqYdCkyOj7rMzUph9QIRxebNgL+sfOSkOLTpyM75dL9v4QKAU4HQNzT31eXHR/u+2lsq
a4jrJrCVWs5BcpypI5zejoDhFdLYc8T2ik4qzUGxcPNL6Po1xuxZlK2SnN+q3C4BqsssVKiFfN1G
hNdHXJj0cUg+WMc1m6yVQV6nLWos5pUjVEtn+BTPD7Zf0R5wlbd3dp9UlWI7yRD2ocCO6WINB51C
aTl9FynULo+3FKpgqB7X7zibdm7RPzr9tLxgSiJcoXhrdrahOsIGUCLIt3ML1eI8CVTvevt9qK0w
r37Qw4gCcz97VXgU5ysAgkVV7FntEL3e7L+g4uFnJ7ff7UAEVpseel1ADKDNgkk/E1WDXB+a5H0N
jgnOgPCbPytRQ7ERCQOZMCV0ROU209IJ1rw9vyaJXMd5MxSZmqKSTkGI25QD95XKX9JVIvTemU5K
ZbaLqJUOI9XjYEzNx2PsFevnOv9jB/LTNUSYigk/NkoYe2QdDmgDtCKjBB8krqCVC5Ef3VnXfgDm
98XIjd+CaNYVkyla5G/nakR0Fr2RU7uZTWooqk09RBQ/S9qFFt4QrDKwk6YuIbIFObWufH+gxUkp
naWY8gMO28bQEXAZNSZ+mFW7LEGYvad4IbJhOE+Mr2V6A66MQS7Kypg03J3NaJm3MHh8Pqle6HSx
Ra+gIEdLupU9lT84Nzm6GY4aH+OorbaRVKi1i7LZtYy4s0/2TmIyDjK7MA3C/D6dk3fqPpyldq51
lLhqyQ17heCDdzkdV1VkTzTs0XCUmBHPdWpgrWzRXBpy1R0StQFBFnlk48IXRrk1eXhgNy0bYu7T
2QMT86KZ9r0YXggDjrlGHY/tSb1Ygafq0pU5Golo/4dGIPvYfeBXNHJbVNFFRxTntcrCus1VJGwY
++IMc5hvIQiE6BtiaiNKI7qJQbR2L0Am5bAxPAxkcTYCoIRa45jKu27KMT1+em8nsqpm3Q5W4k/C
r53ZYsmiS6RixsBkL/HjSgVRRttRQrLESjmS6Iy+0JJZKk6Z73V1+/awh28HfbvE1Z8VL/WsKujb
CFjaE4GWHBKOyItFasLaJs+TJwFhYqEd6EfYECSM1UcqsDjka9B7LUVx1g6E46U3ugPXAxw4M/yR
h84rGfu8AudTil3mbsg+zHiC6e+3bEefScgXgkXGBk0IUQpvxPxwQpnBNNskOhUcu8VmttzDl32Z
1Es46mAefzJoSDVFtb517A1paGBTiqFQOqam9KCjtmeT/JY7q8k+S+lmad8ktQ59ksgMemHLJMrM
sTCfbaxeK7I6jA6xvWQS082U24gvs338vCrjr9swy/0C68rhoxxw7EJjuQl2S+V8xoMFD+Fkh4Hl
g1KHshy/zpe0WimqF91EZTYWBJsxwWNt4qjQGfbdqW0zWBNALmc479m65Ap7dm8ZpdSvYIrMawb5
7DE0V77t9frdeloroEKpbF2xcRQ7uCaycnexzJLr90MKjuzgPZwy0uFvjL32YSY04PAgfmVmxPUx
4MVUrK/VK+YGL84e6+igUXPltGjFtYL1WKdI3G930x6v2q9BusFJKS899ZMtw659YGS36NA3Yrms
lEF69pahfmZFWiHgU7NiegAYCXFctYUaqCPtHT8skWO74Z1Crto3SE+gU3od9iilbFP4aPOb7glV
n/if9GmyGWRP/mi0rdyslZTAm18+gwnw3qfFbzieWNUx3PpAOmdxepd/xRdZLgwliJS+bmCQhMZA
GEXhl7PUvsOqmwHQIB2wEMux9LPVhs8SGHy5OkLcjLyYVlSJz+8uCbGtFU4ZRXuGrMZpPG50S0Q5
YrpCGdWhP69H/B2SfTCug4+StRaDw60sLmC/VhrZAg72WmpgcPe0gIlU2aJTjC+LMXufK0fLGOGs
k6F+M9HK+669Af24KeoOSJpeNfz491jEkM0SBj/0Z58mU4ezkjz+jtbgfBz0VpGWDrOwDnCTIjiK
1jojO+FkjpmbX2HayPGTdTzcm/Ip6lpZaU54liXATCDn16/MAyoM7+devKV6866p7RjXNFcMbjuf
OxwaeVkXeo+88oZnHGfZ11EqarYkDgctrAW2pJpjC1QZmYxefZ1WRqkDs5ol/WsK8Fd1PKouyUqQ
3Xs8Xi5pTARj73w2Srff+Ao8+WfzIJ7YDYgItKSsR4neIOnR8CYdGODRoEuIh0aorKNjF+VtdkDk
xH92w5sndv0RfrpIhTal8BBzQv8wpqDfbaWWCG6L+1gqO3+u/o5SEVqLPNgAGrHYa7VxuDVaEHde
igwBOUcEzK1XJ9jjTyf5xd9L0YD8NZku94ypNqPdk4xUM/vSewbn+PVfPhFlt+oKHtER7tG3SMJU
4GPgKpIhsxqyCi/iWFM9pIOw0/sEijJMiV1zGee1Df8+KBpLT661S8PQoN0N4R/msDqXdASzftfh
KnkE6JYybL+ji3wHKGLZ/W3SMOcS1u/xA0dhNRnVsNQmS9H0Lcx8UeV4d07dhYmDuEDfJbKnW2Fs
2hWVIidq+ZfGm/fuVc8ekwf3P1pSBrr/TivwH8d4lFC/4LT+/otOjUFAh24kqf6MLLkJ6q7XEzuW
j/NXlYAM5adu7YTJ/tEJ6nXOj6spuYTLvjmn/te0ojsK9G11TCTnsNNOzvBF0yx9ev4tL4t8aKPR
G2xArDYrehiF1G9jN5kbElW6Kfv+JmoEwfMIFMK0+VvuEk8GCg9ugPxwNlkswq7VeuPHIUYLR/Av
3tG4JocyzIbki5lcFga+ZXI4+qIwVxK7miaU85s24W139dIyP+STrK0ozRQn4F9+Z7H7uA/Gm1oX
GltYledUaB9CFS9eKbTEuU3/N+J4KsX3/vChQivnhyTwNchbGFg8JU4CZDQSdIHxXTRZ9ozZyRi8
pTvJwR5jiz9O6NnWE6HuSoQEEnjGZeN7ndJnOY96F1TByrJ1zgWx5npyYySDVAOKbe9ne6MhH+pJ
3MI+hwY0roor+/gCNOTRjaKH9GsYWpcwSRInSI1DIaSKWfH7WpxOPehqtOcJj5xZEoCcRiul2A+x
Ttcz423XyjDiK8+AjXhCu4zVzEbyiAuEWDOkdXuwmsvcdc1w+Tni1oVROT5c966hvwe3o6RlXLQX
d51Ih93gXpz+w6Wu0O8W2OCoYn63gJd1JAwBNPQHj4UMWw2mAZs0w8RQh9jPOBznUeo6+Fy60SHJ
B7wwKOU0ZGRb3SYdHGhASbAYJbz1KhdUz65TvGmRxtH4dJAnNDS0sW5zyWNkDHme+sIzG10vjJI6
i4mNDfSkQh2jYM9LTEB//Km2Y827Tvjh13G8fNigVyAaUH/lwkcpOAyXrDAh9cUrF6BA6qheevqt
iT5Mw7BizQbj8IlqG4nzT4pXODNsKq82RKXI7kKxhaQz+V4sD8RelObblpEfrwGU7qoeLhIn6Ns9
/7VkfcwZjkl+mZ56t6qjpzg5ZyQDcVp8Dn5UvqUJgoawlA30NyRX15CVwiRFAxaxkNi2wl3ZJUQi
f5T6Er83ngljyufuirSuDsfxbM5m2znJczz3sJavkR8W1udXpv8qhrKcZP1t5FpCJOPq6LSXsQ1f
/2JyB4yACbAQSFkPaPIbQNGNDEE13p0o6NbEKqHwqEnzKc85NXYZ77jmWeX1vRD15lBYXJHNOK7c
rjWeaM6REtJ1Lqu1aHonPypjKt0gbTDvrl/QHqE6Pvk7A3r9wU3Rp6Coe76yqIniRbjwap4r+mcQ
zR2rs3SxGjxYzGvQ2YS1YfkbY9PgR5IfafBEpubHt+5Dz/SudCxM3laECXGCr5Q8ALtn2FPcKE2l
I7ecbasitj3pOvoDYFUsan/eDo1y1W/sq0A3PU6/X/nW5zQhSGbd9/W2AlJop+KoJoZc0n+uOPeA
JO+UEg0MFvMxP7Y06mWe2VM63q4wuZuF32skyzkE/0iP+oJSNaSuvTfE8/0QWwirocy9amDgKzVZ
P8Mnwkw4Lq2L8zw8wivLrL/8lyLj7i67XeGCGguNK9ykMkqaQvjQwoG4Oc1o7MvuzSuVu8QZpLHQ
kVldBBziilRjFkNOYQl42wNjsNj6IUk+oPPh4isXSsuB7ZKcjx6kW3IVH+nZ7fzup/V2VkoB1Fpu
GXENVGW2N2clkvY6vxma0sWXrbEW2b9q/w49+jKraBfmjVJnCAXF+gmavUSs6TXDbpSi8/3sfq89
hE9BtEUisaYP4+meWbLjLNECL/zfNNBpE1zXz+spE/LODEeScDPbZ3qP2M1QH/l7C6aRm/bpYD2l
vT7/8n5c39w261gPgc9KiDWmd+Xu17rmG9KVNe3+fHxvnQiEYn8nLyze2gYJv53NIWwDxHmRzPRz
DOE1YzhvQjl8tQZ1w2oxJwe5f0CAD78yxMX24bcEz/j0GVoiaOTcYsCqSTHQgt9lN3XzH7kddyuX
a1RHCNttXVtev4F9rzAePH1EMEqh9fMn3o6SZNGtIv+paZercB4/7eWDVcWdr8mvSlpt8J13/uEc
UIXhffpNsNjY+PAnuJkLujfYbHMoa35fPV7TAnyVH4L277zf73ENyVrbFVh189NH7oHRoGxamFDb
ZChU0WSXZdi+w/RZGdBxyT8RJcSm8uPTG0wO6HqBJszbiRyl0dwVdJeSjlZouw0Tb6gez13jImR+
sFCp7kDqlFxac58i5JsKOJCsmUjfHP406IK8QdNgjJS4lN1MAyUDf9wAxwkAXfe/IZi7JJ01d2EW
qfJvDa2hlU+XjwFzzzFIKwoibHcYCdOKU3aqMORlNrmoS6Dv3r6x/APo6Y4Jmxc6YHBpG+SmjvXy
1qfvejcQ1J69tJ4WgIzCMFsEj5uEqYzK1gc//Dd+RdU0Fwt3xNvS23j8XYmqmALR0poZ3ByQKXRz
Njg7xGAU+7MaNBH68HZdtIs6i8n3SMtw3RdhRuCs90TURj9SWgiQ7kO7RPP1JAUmdbRxAc7+SWiR
Yr6vtHKjLcGWxpUmW+sh1/rJvGlTokwnTOBZgNHHMVr9K0UnkqP4GIfUG9a6TJq9OBmxUc5G6jTM
wZwfmrgGB9Dti3/D6dAwTxMtyUr3mjkUmzZ0O3qnk5fFd/2F6Xu8Uee9ESSHjRlZqVGHuOT/a5RC
lgTE7JdSE3lP+7xY4wUTo1gaLUntuk+Qe3ATQvZz8t/ynnsm25L+4KLqz2SlycCXA16HKP4+6WZz
AJoBDwZHuhDi34IPkm62s9SexmvRvAs75SAyxLS2AUbTebbkoiCtxxcQJ8WB6FfIpSy2Kh6ZolYC
usTbUCGtRPYNM1qXJGOeV9nm4oKWr4wzBkfh4BIMPnARrSKfw1fww/7DjlKy9iiOkHZWOl8ecnYj
Sz72V2Crv/k/cbD1WWC7SbxZ+uOVmOH+yLWyQAAq4W0peR2xQ3Aqo1weXXb0Xf2yqD7VxlRrOIu2
zpFhrJ5reBJrWJDkjMtR+EfQxwlCcy6mrRQXnOiOFD3XHJK/zkpWaPi2cfjr5q2L025+N+qVgU2k
L3eKKmMaActOGQ8JXO6/FfTzS+02N38ix96mOpMLILmTQFN2bkTn3GWTGx3TC3iGV35loOG7UzS9
G7flUO6gsiiqB1IN4JecVo+uwjiGIHlXs682VAGJu8zsHauTzA8toS8rhMKCJlVaM2Q21khuk0NI
NWE6DgtjKXDaZjx7J784n3b73mcWRCfQTbRqigpYEE+XSlx3xJZlW2xBlXUx7DzZTqf5zV0ivNos
TploEX058oKBsj1fXQ3mP3d4gyayDdhEkdEc+0SCn4eV9/EAJSXJBBjREB0lHt/f8lWQbkVEZ+Ag
ySTx2dGM7r9qTtP3e8Ve140sKagbJ/aeYLUVsUvq6OruHrZmb2oUSWM0RCllyTTH7AhuLpYqttBd
wRcLVEBTMK/yd08WJgnVjdf7JTU5d0csJh9Ane80FoNTk+E7IPmPx6YU0ArIC1hYg+bDj2r+qsiy
NXY7T3NHskLiK2Nf8ahFAtPjXu23Nrd9FY1RHAvoPLSXTVH4DKrruK7GvppcI9yq1WK3nYoTmqkn
DHsQWEm879bt0Hj7Ify3gIZDPdV0NpQeYA18+rxxBBo+cRe8D7WaBtJ9VMWU7YKbJouzTSJvamkL
+Qz0lpDklqMKDDf5RlJObFTg9gw1Ko7gaj64qSrjK5QT/BpBxdk7fPSNXjcfJSgdn0HN2nXFa0O1
NrDAqylkxNvSdgJMCLc7LewNzujjXRMrh/xQpaKTx0oFTkodlN+IiGXH6YDJQZQkJPSi5WrdJWjz
FGShiKOoKlWPAVMAi9kHmj79XUOyuR/reDL9BNT+eOMLpsMoC8TWzS6peK1JaouMPGkxZ9ukZTBQ
VY/k0OxfTZa0fAQjuOHvtxb1r/2MfOPrRLfGiOd3D76bdir9r5MyWmLcGED+zClTpGu4ueHZcRfk
M5y5z/+Fpi47r7MK6u7lFbIhhMcLWfKLI0LY8qvlJCRRNRFrH06SLWEhdAA28iS8s4oy/cHMVtAz
PVMNxFce1Z6hjPZqwxxZmhxxYQ10XknSANRH3M74jF/ZzX3/E2M8bq/8WOZ+uMMWBbJGzwOVWqk8
20r46O6AgIvsKWKeYaYxLgN/pvYa4Zh0G2GqCxy9kgjz2ZOeJEXn6SSYUdhln+TBfnwFx1q4Ott2
4E5p4+1NcewUQ+URw9z+xIU+e2cEF7l31u98uieow2MajFpi5QIa/0G/EbdyBGeA23c+7PdFGdwx
V9DRwrAqZxEw1vUCB0Qlb7ncIcX6rzyZ/N3CnXzVIkjFN+NT1IAaNDKWTr4+m97XisBeSwfsyGMj
+X3iu26ZBfXZmDo76Pk5yX5szq1ZI3iAtEp+vc5nZ4qygfq9yWb1YDs4klKz6ubBq0hYKqvpY/Es
PvlykMG7Jk4nNjVoaZgWRSFY5S95oivaYIZ8ouh0RmxVTR3DBpRueyj/nac/IU5OGYrmHbsZZD1f
pFlzuftXth2MXNRWzsYcA5fgxpG6IymPonULj13a505+fRNE7xHgnGHcTpqHYimqqLAiz2doqlt+
uDUbvDuyVk+GfpKZOVGdpfJSUPy0pVr0uyTZPazOChzQfUCiqWVrgzZTsL/GOwtQuMs0r58ZCt/t
qYqRst53BeGEc1F2tNT6hXG/g+nzM2BxQ2e6aXPqb1dOr9LCyDujCDdzfvPUOXwZoqQJkBABoT5w
2dFOZyZpvq/F/P7oyeetV7RTFIxkqQjAnOcC/XxrGHJ+/jBQH35+ivkhOYPdnVNlsry5VguaCvCq
dLIPsI4/b6JXNTD01/qhbPCZmdNq0vZrtkA6pmPtHN7UL6jHqzklFfEPy649F2dZLikxLW/ZrjiB
NKt/2PySpC7aZ9gqdLtMPnjiAHAK+prSSt/fxLI4A/fVOQoT21aK4iMsITZtOzB6i1jw1xsoXo0C
v/7LUS7h7ay3/ZqHsKsGaKs/4xU2urAXLM2c5jm+3TjCSsXIwCbj3OrhsNHKru/r61uYpj69alVf
1fkGDhEJtEjVrwaw/CAoqWqT074a/uJ0T/JkoKIXCJSkmObSFzQN84BGJzFUetP3Ur++4hH64uX8
Mcjj3KpDyaYCn9v9GWEO6Th60J5M3M6XS58Zxd3piiMcmciJuxmHY8Z3nPhn77LOFb6Xf6FrPOto
cs/or7Zq5iN3TKaywj/OY+PcGlcI7YCLh45hwAXfUm352WxCb+mxZCYpMAIrONLNNKnWEaR2r7f7
g/kSz55MJOin98GgmslDq38rRkYzQkNd+nGNKNjQ4mbu2itHR1aJLw8Kyyh7tQ6DNsYgryIbFXzZ
xZST9qeL/d6q/tT0RuTPI7ASKBdZIMH7PeYKmB7xRZEEedAeY+B2m1dUJEEDYRmWWmOqXuohxkAn
ThMdYAdbhyeJ79924SWTiL56GJoFeZzhtNEvoPZEYcpaAuWZX15Kbqx+wQLJ/++zepjxSr/+juRk
GlBas9rhCHZQCerh7t5L6H2RezW7Hoz8k0FUGwxYUqr6HgFTmxuTlV7Zs3U3qJ4QGS+IZWSbtkRv
hymD74wbLz1ridyhma9XpNaUQkz0qDezWkcbkWC0ygZFa6vfqO1W9eHxgwQzdE5XnG1f9vRh8oGf
StCyIAHmp+g0jl4B7Dp/GnP70BaKLXoQ3ysprDX9C6jPLAhYeVoFVIqc3B4UAy3YRhiHk/8n6djY
fS8FWCUKuqNtyadxWl2rGjSd/GGeax+jiJIJ74H4vFcX+SM5AcpMFiy1qBzf8cCIPLYCZpF70TWD
CDXKQydemUz+MZJjQOgiW9mZWl8ARjWtNd2/IpHCmVRZtPka/umgLBLh7gLO4rQEpkTe354tZZkH
hKjEmMq+uAxVCMGki5F02CzzFSgGtOA3rvkxGrZ+fKzXfXgEPFqKgRR/xqI00lG1g9eOZyXy9hSD
91if/HpDMzCULbL/Jvgah/O0eP3a0OcLgtWoLC2qQj6D8zPgjLq8/tj1xcJZFeHsPNdX0ZoZJ1d+
pESIrjS0ZCyBTr6MlujgpwBuw2kMCtrILX86Mtwpy86poT84fXNH+uH+sF2Ed4+0SAGYRjMdT1Pa
HH/jR3tKVKb/BZTh9ORKiTdL54VU6CfDSPLX3bLQTP7Up9jAr/4Yhc60kFFVi2na0zlD80gQTTCy
WfOBfN6E9o8C/129+vGeDifxgVLqLhdmlUr9CWHYkWd8D+u2azO9T32paOlZRDQJ4h6b3HF7IgDT
HrCzrKacdE2E84bzUCQyfK+wTzs524gMmQM6QOrqlZLfWnw4vPU/rvimq3hUIDWNXos8aN6iNqC1
xbhCEyJzvccnGGH7gg1OjZQ/dslB/53avKXUyQnybT+hUf/1D3mGCsR2Y/riDZMpR8M55X6rg3wN
/ojNLK0UkcUdaAH0RZsmqLgjaPSJ6Pg/ZxCsO0PYVlzd3Q8NLrFghmKoVNM6/1Gc7LGVVhHrHAmh
9aJ+AncU12J0OubOVLjVwk/u3E2gCaB9naG6rmATMFkmFtFSt7qKpoiYr2EBsvS5kwCP3hW77/OV
HvtKG7G52NrZxyidEe3NTzbi3LdvzwJ5N4PHoBbm/p5NI9JASoVhsC4I8JKSTomLDQ3a9C1NPWf9
6ghn+5WG9vGWY3N7Pe3qARP7t+qXiRgEC2keqhc+bD3R3OjH5eyJAt3oHw0sJMQpCTXCpFYJeylU
DknYUXZd/hJjFEJ24kACnnNJE6WL1D9eTfNwQ8WR2Z39VKScmnjvcQteO+ykiC1OqDnpTeDTegQh
Bf3Z7m5wEDTKOvHMM1e3xIdqR1IX/2o5z4QtBv2rRZG+O6rdrD5hXgJfN/lLER2+lQBhWFv9IkK0
+NYdxJT2UcIAmdUT5VhZUw/KUX4qZ5qliEekPG0sQLJb+pF0YUPFDfoGHaHmW74uVMBgb5IlYmk2
mXaODbJUFdfnq7jz/NYQ1zSQC/YnWemVaOOIPWIBIumo9Is6eL3B80ElQEm1Cku1ULrCZxOJ7/+i
djIOE9JW9ZAGQz3fMCVQ4sMEp24wDPbbTt5sC/tEu44ndUrWw3IIijsjTGLcN1Lx2cohKVpb2dQf
0rfNuYbuigvUb5qGOXE52C+Ph9yIckoyU4gPvZJHiB1v9SZ7pBmobzlB9GAV7+YGn+r8PbIcrnl7
zSm8abyJJwrRBmhCCuCQ27dfyZEQlcJzpYhzHKk0+nbjrDIRjdL0uWIZmCkuiDfe5Qm+RfuOhIG+
75GewEf0F9re7hb499kpx2eM1jvDEOgaSLzx40kLKhoK0M3m3IE5NVR28an2pGiiE8eVVqBDKqyX
NFVCG8NxQq70TrwEcUJY3kG+2iJ9tIl2XMMp2RZ5ya6neXmRHD9pm66/aVIgyqjoLRZ2A4kUIXYn
UEHTYQ/WPtHiO+HeUSypnjvGYR1MDAK5cbSsLnriuzUdQTxC5HsMsZ9GlcBLKp8G3SLxpXFjuVk/
00Z44VFnQ1RMlpEz8t0sXQg6FdPaUs4m7c8pdqZkCl3x/ndb2nzYYYxGWmoETLPwx0q/jpA/ZrE6
8GZpCHloG2FgeURLuDtWdxTjxQHovOXL5uBBMj9WH0PAq60wEneso/mT35GihnGXdOXBQMIMhhHD
IoyD0SViXaIN4YjHlTdvSWjQGYYe7ScrsebnS/vETsoOu0ec0A2KilcEQJ5HOZuiwaxpNYDewfcS
HQuY+PysPh/jtNTmknWtq3tTjl0AGETPs6lCWe8Ar1eSIN7uTWQfBPC/iKw7wyjG85gU3AlxKgd6
CKSk/zwLEKN4aJ51YYItZwWhpg2EobG4gSuLJn7txVQojuAs0RRNY5Y71qfzTHsgHcbXqsPKsASM
5rCrMonFy67ke0QsKcmHGlZ+uZO0fBQRHtRV1pfsL8FFunkcpPbnmK9Ir+bStLk8wNTwCHSPKQH1
JIIl2ElVDnVHTYdCiJpOCPB46tmLSGq7tkoFw6umLZ3rhyLnaL6QNr34XLJhDMm5Qbh2fjjaEnXe
ksizJWS8uCmUqj7SadxNJXZK7Qe3avgnu8C9StxLQT88paRH6bGpro6HGY7lVunUgb/iO092ztEU
ZpqSKpQLhrVicfHNHjrRPa1d+suifmrCDFVCFw4h8RYAdrHwDK19HVCJWlcQnfKIiQgtkDtym1qn
wRW+eBhLHcHKgx4J3Xvn+rDakjcpWgAN76BcKGsaQ0ymgnxvJqDMy6F+9BgxTrXdgTTZWW2z9fic
b3WGcMH3TPF1lazOUmgKYGSnOQS8vRRSn6EA6JNc1xcP4EQRAKFGASctVmPCEFA8uLa0dEFI+lfr
+Li8LQhrFuj2J7cIKkskrmejHdtITW5YcP2OofzXcB3XiFCQxuS81ClajaQXp8XNVbR7XWGlOE+f
NsY8CMZej8271h31XlnZJWj/fRX4i3Wg3/OSmKo5BRYEyeLPod2R9YOujidGZCf/oPBYjcxybZ6j
8Scc0mDVec3IwkrjVbMEub8xcNkkcvdXeGdQ5aqEXkWYsiSLfPM5nnNIhwIPW6PAHrDgaiZZ1s9m
+o/ICT1SFlV8eypa/u+3FBCkS0l77qTxEW5mGO75o8f3HCYyUVZNhDR/Kkg1c/Wi95sSiqmueyiD
ZPC8mOp0bOMM2nH33K8vfM7xWf2edJzdP0Wo176+5v0QOHuAhbLnG2ylh9RwYWxG3C7rQIF2AMJ/
n3R3Sv4O9zbYc8nT8LCqYDOACKsjZ9dVRbk+TaqUlzMmusuQ2QVzChL1044/xdQwi01Rcvz3cZaD
DBrLpwtoe+aewSnNA2TnnlAge/DxDyq9wa88hhVIzThNETl34/mcSM+Fu/Raibu+E9PcrHfr+/oF
seo8Nq1009j8gKx/c2rhVVsxypGONy89NbwATx3ubpUxxdmwcBhlItTLLVxaBbky53lQq8cNRx7J
jyAk/tsJ77yuJAzP6bTql8tr9Pbai4sM/2stuFvmNreAIYqe1qakqBvskuncs6uAYUdyseo0QR5H
ZT4V8y1+oxS7XNPRDFanXfkc/Qkf3uJqdYOuG97XE+XK5dc5IGj2msuARZU8jiNN4c5CBL5lSINQ
SOKBbP+/KMAngpaAZ9RyqWxRV36JSxOqx11Nn1k4TZuIQN/BgZCnR723KXWSQj0rArAlrPlisAv0
GKSD4/2D9Q8dqbQgqAMiGMy9DBFtw9O0WJaCw6Z362cD00WEed9rlgxv6nmRFcKfvwIeG1aTmEvV
v1bTFrwB5yAQ1RbsZiJNw8AtcGe/z3C9G7OEIfUrFmsqD0Oz3vimFW+pAof8r1MS814bsdWa5ASr
Kms1p0UjIkziWF7zMVX3ZSlBxzwu99F+V2ukny8PnqdcFZcOcbUlWBELila6oRRbBiKegGGuNrOd
/JT7ICeMnPEDq3DXyo+7iyPfJILaqiFaba3XvfjI7Zsht99nbJxp/bNBfY1kjUX21/N5xLus8TkX
9lhwL1wCZFk9CAE4fqkiUFEtE98fAFeBBzqv86uX2EYUdZH4B1dhfP1aoL00Q+3M9yrLgB6sJYgL
2JG7qrEVxR5mlmCh6Oq0BZKolgeACwJzy6p3mkTEd5u2IIEkBeXT3mIRqSCcin4jueKRjdai7u36
kk+1NzUVuuBfV56IGwG2+mWtW6gapocrX6uiZc66DVWcICga9t6jbhgf358U8GMH3122nJ22VQsf
dtykSFZW91gQIdTL6g4WJwQwuV/0xroqL/KQ9MsyTfl32lOH3zCeDVnXvPOtCk8K9hHsUx0WyUOl
mZL6ngBKO3yxNDbjPz3ICm6+A46YGO7PddfpPi16tdiTbDhaQeSXwctk04r8MDBn10egOuNXiZjv
nUIIX73j8iksUvbHgQqMee+a7BNeRiKu7dLVf0SECDm46kP4n/GTyUhCGwvk5AfwiYHKVMed+Klq
gAGXbq0SW2vIiquCc075cEoWVjK7lidK3MSd/3NheQOsoDielAGLLQP7XtX2aCGjREvJbm/6zmBI
oXBEt98zAHRm2Meh7usoZB8WEsm0odd2muyasToC1ucqipZIepaS4skcpQ+oou4M19bbd7tP2ngj
WBLvsG+qUgRoPhJj+kE6/+p3258hi/SY52cl2bVFQVvvLMic57h69f9EDhgdJD2hQwkDAW0bd9TO
FUXTC+bfE/54wAk9R0983+H+3DMe/DH1au+m3MuaPUNEgwcIdxrfqY6ezCfjRm4Bnc0wStyg9rhI
6wtyljL2mofjLe8bobgMDmrTMr2mxDNfyvUCdF7cwDE3Ki1eYlYmMupxL6su6VMJq5ZF9RGztrs5
f4nm5PZlL4wciJR4D2XeFlQCxZvuwiCiUaG42AwXEp5MIpCHHE2SgG1fLmX8eNkF6kP4g/fqENiP
cFS4BQUyqe6QdJetEHLZuIvaI9kjZgOGKLnE4nkjrwtlP7NHD/SISz+5S2rxo3/xWlpddES2n4ZN
NkKW97DZxYO7OLc/pPiQeCxMrFHAFchueLUFSPMg52qXnoK+W5/qAD+C6zCpsN8WLFcFYnGt1j+q
AO0/HRiTjPeuxEl7Xvs1gzA5PMU90iPzwKYRMKGQst6RZl0Xaa861XQthangJPRWqwvthcjmqSzV
nWnrsRVrvENn2HZSnWNHGnkpTdWKbRLZHbi8NDaQK+SxWkXJ6h/86W6dCsVQjOhlJ6ICw6oCEuB+
t/sXjRT+o5LZo4H7xQcESoN+umFtFKxsDin3GSMu2fW+KtI1SjoCMdln4AjOgwd2f4GPZ56IDLhC
hi3tbits2oruRbBd/9JEscbYbIU3qDpUyEKBs+pZbcSZagkR8DU9OweKfbFxy53SA/0y7Vy49QAx
tyzy7p3b1dldpP07h1rds1YdS4z1MLDtQ4SauHWWRZOzQZ19DIpXW0bxsTiD2rxnE2dUWkvFyrLW
LuUJLq/Q80hLJ3TXdHkioE0VD3MjPhRcS2GKqHniwmVx1M8DaCTf36LiN532wjSqZ3iPmCN9nROL
rK6Qaj5T1Jofh4ownQaMdKxMOVgpWp1hajJxC6OEWAiNa6sPfOVIysEDJAoWQwaWrzufGCUM/7Gw
y4D75zq8W8ezSIWO0oMQmNgSv4PNqPPRglvff9I5uQpMXEz2qvZbGFZih0LnrplPypQz9MTqVWKQ
8VIwqfMPljcv2aTpH30iqsk0YrXkaq8QdHoD+WtOUQVu0ezlOvxSAUvN3zCxzq4V/K6XJsuq9a5F
QZZHtAWmHWcOLobjC0dSVj916npXW+4jJwz2CfC5z/4OBx2wPzOFx4HdOwYu6+yFreX4xhuiEJmo
QorXAmj3hcgUDxT+55oBrpg6y0YTAyFtKhOJKWTwfG19as5YHIbx737TXajtuOan2jup9k1iRbIt
UiuqzJWWjbfkywJLFFbVWcsaNhZAz7qisw8209JQefCGL9NWYgLgEIBzrrU3McK4UmFNutYSHAPw
DWZy8MdZf95tNtIza/Y79JONiaB0NcUxEBNQYy1jZMd4wQHv+h7Zg7LMt3nLifV4fO11lfXBO6WJ
K5KTs8HLwZPHNNKBOhjBpohzSFopt1/UIQVfPEj5AA973R/4/cW1lD7R1GBPba0oohGY1mN9YJzE
2j1Z2u17MSPwkJH+5BGRmkZdrtevzK+W2JoyvR8t63bo2udBbgcBlnhpR0Md8SvAqMsvio/DjBKa
d1cGBj/b3q9GWbPDF+FYdPzyxWZPd6nnX95//fDSnH4OgFDflZ5jFT57jxJ0qPvmjXg/kRkRv1Wc
/JAQo6hDGmy3LmXeMK9QhhffdGbb3+BqeIblG0HEzytsx0jdxd9VwYz5gcJlL75zCasJPu21DvH7
NWnlwzPtXbj2AZtBp7uZNBg3UzQfRZeZtxqYuh5C1PpWfsk2xEldI7cegYCv4FjnVA+cd65rHQFs
Xm63JFzSbR/lRitjzYWrsij/C954nnBM0D7+9Ja1vEdxGcxvby85EkgbP9kOTcfN/y5daEoWZR7a
GZTKaeamMc0bM4f7OpFXQ+IOMJoQqwxCiz8xyXkyyILmnqbRUF6UyJMq+Bj3cgup23hq1jUxIqOo
6m9lbl6Xd+Xqq3+FY48ddHfxbkAiT/jiWZRe/P8qelKigzJmPr48BQiIyK52SKFYFMJncE+81EVm
n5q0gpBkPRwZx71dpdDMqJFZHLoNoGi3kq/7gYnreKWN1w5ujv9DDnKoAr8tJ2nYgv4tMmihkC31
f5qFbp55j/h/YQdpDSQIgM0znt1gUp+EMgKXkiUcuJ0YbZUwabx7ht6HAnA3rBz5IQ4LCWyMdSCt
QgmykrYnUb9kl886Jv7pewfbNWgUEvUnWN62jtA/BC5opEhJc2lQjwtHYDwvp1L+DtCKYxLM4Mzc
yKUmpEQVSWnhN8NegjZ1Dkf63RePuykRRvqffwsBQW7QkjaT3Msw3xsSILKDuipM64riEKD3JSnb
ToswlCH260Q8VZvpE7PlZzmQFH/n6RFgvXgEL5KvYkrVPbkfdqS1tXJmTbHjz5XbGls4WDogv6CM
O8s0zabiaL/c33fNsN1v00zzETBlF+MWPxVkYR/jMEvJUVQtbZ+bImUZsItWOxEMdza9tNOY6EMu
rr9GXkIjOeqItZ+bfAlhKTkTmorhZFTuqE0ebC67llmqhLjK+8Shpx1lbWu2WVVBc45Jmfqs+CMb
k44cuqDK0sNeMjVzHiDmKQuWhQvc7wI0lpCZA4LXBhU5qrHQItI5MqFa0w0xfc0+QTpCiTO2bwQ+
SCGDyK8iTfjA6lKgqv46HhtRjpQB3mTa73UzZkxkOCd38U9kb5b/He4c0EMFJEalyebRuqJuIqFd
rgXAKhehk+ZROezNzxgCiYf7TrVmZMmDB5NzqC6kkUd6gxWSORORZYT53U9HvWjj92/+QwBQ0GGi
5VEif7+PslJCKtyskWiQR8LYZu8S5hu6/ULrhEqoG4ihEb38T+Hwpn6A1nisYjVQCGSVFunSj7a4
37R0Mx7M3M+ajEbdnVpFMBFU3IH0q0hqVj9jQcCJ+D/PNDHlrFnYKjnwP8ZlIShsPbm1KWTmJKp+
38LRGGL/VC3pUkIuC2KglzLQx5cIylUYsXkrbtwUMuqLlhHuF8x/O1xRVNmVyToSYyWrKTzS/Nag
HpSjARmy+yTikpMg1zEa5RNwPQI0z6pJG3k0Nu2PKMxdKVyz3tL4hAmhJ5G9bXRGU6YhrwL0tzi+
dfyxlMU/eHBOakp9Y34jiJrjwJ5Ac/GAQCVUXh4n2uAhEUv0VfmNxwz2X+qS8xDnEmXOLL+b5gxa
t26Y1HBWjZxySCiwGvSlVoyFMZmt9RA69i/jfI1QVRbdFhnIFrqm0lVaqkRsouuSCMcVanpau2MN
sgWEKYijQ3t6uO+9nUmp+0B7xM4BWj5nri1SQoL+XboO1erzr6Pwk6vIkhKEMOKqd+fKwq6OJTo4
zOpsfN6QIYUsuaxeqzsHR29twxBIhIA0fu0jXbhWNwtgcnMlMGMRPtF1nPMYvaZvSU1O1GGUISAA
RxBrnUY1NR8HwWRY5V2cE46f3u+QNcy94CBEiMdXbz+fpMDDPWAwBSPsG6tGzOaqS+zB3/q4ZVpK
Z3Pya1/h47ObohwNOctG8YWp3d2aBtxKr/Pm+DSPZ+l6qnKn5LW9OlKH4a3Xkn/HQSxsCpzmGuJA
vg6ZwncnbgylkwZj3xpdhA8+TF8vxEE1o5eqgIrLEANwk6STk/xLCnIUZBiS08CMwDr4QNvOtK2W
Qsf/Pa+lobWtxaQ7HmZlvoiW/1YYi0T3clfd5kajAVttuGiOImjlIM2Mx7kmcsFjIUABplQu4Foq
tWZGxxVN/kMNsHLvx7FRXHHQdq4t211UixhY4xMQv7SmbasbAsZeqvZVXAJXKqO+2aXZ6m6ScC7X
+gE4YGXVOwgniMwwB2YIVVo3500JwBey8LxfU1eVRdAvscMwLISXNinBkbrDyceeDPgVUdgSKVe7
gmE5uY9ZzU/aZ7x2yI7YoTDZw5Dl5BX6goLlGA7A826L3hLQKarpnHD9Gjn9QMEznDsLjcq3X/uw
QkEiIg4ezghJPABbhp6LtHopc6O6uADwoO5BY6pup7vh+fclYW/pAVP5y6Q96/RPTI/Mc1GbEIHD
G/qGvi1VBJtAIkJSiCzBBxugSqjlB1AymI7QaGKen7xwL3MlIaMwLCdOCTtVb/Y918+lqWB8viIf
ofW4Eio91FlinLOl6ETpjpT2G9gTISohGD/iJQELmeTCeiPaSF3GG+y46QIjMWPllI+tplsw8GPj
0xy65qsATlyC4jtzxGKwHJXAUbDA2VYbOQnSgZ2rrQSzEDPBsscLOg3omPFAoJ7jkl0H4d2hoLpy
mgG4+HRf1v4RK+j9Pt6A7ttvUnqxrgFXsbopsnGZ6f7/2MJxFxV9mvnmv1XyQfk9ejg43uteQaWc
6RHs58WaS4FZnkmXsHauIyWFHm3m0kr2J4E+9hFcqV2MPM10Ap02NSXoXcvtSlTimi0z6cnBk2gU
Ry4c3Jb7BWoxNTVDNw7AsXZgB3uqgkMrZVf42pxTY4odSdf1BQnOb4w6k7G7ZBIs3M2YkfePARKM
O7aPEsR24q7xJ00MlcE54JRYIdz9yYzDwqyuqDRRSLAgL0YwAgxxdBJJed2jeDo3Z2pwkPV44VSY
/Uik2MfDWP/w56JcDr6kBDI5Wtv72v87SW5NNmqyoX5CLzkyCmE4j/L6UhZbChzv+Qm0B4dV5Jdx
I5mqFaOdlwXnYPT/zRWWxhvATrZquShrSwfTGvivFKxOi4VDWR9fZE/32CMjOlwh43cpQ31PbNeK
Kw4YeebMzeC+y8ZjQG090tCqRTlGYJ8dZ7hGoyCiIqmZ3Dy5ctSVdfuyzDXALTXAPLBIb99wV0nc
dCk0s9or1wTBoyjvqMUz7rgdqraG8+ofPisu4vwOn9snsZWQmr8EXq/9aADf5scPQgjwZ6yrYaBE
WaVgWdAL/8FNRPJ+JshtBkCajiTkbXLlOABWy2BkTDddUyMhlrUK7HKqxt+amsvsk4WWVtxATtDW
nRMOyx31c6dEmNxBJc5PpFbJ+ZSdLhk+MZUkuNm5diitCANSf5pYsxOv2ng+cgt4GLvXzus30gcc
1EAEwW0g8bLdiTx3mZLSosJOAK5RgeBY3Q43pgBwvXaUt08+d7dJtVzXok7upBXM+WkRFlYZbnEb
CEE6ahNVIwsjS5nRk0VDiKp/OLDXuysUTjN4V3iCEIal87QcFMVmIeeJem7FmjOu8P2ExbnIxxZs
xq6ZSHUM0v0UXj8HvGUIfLKpLrocWbT0fIMuIA3uXjV62LXyXY6c0ulFFoZBpFs3MLcNg4sZMpyE
Z+XbSuONhe6qpoCFuZvImnbQ/blcJ/WhRDfX6FW/LyRl/vqGKIlHoFQHTB2wNeZLpOuz/9mVmXtS
cqsBPuMelQN5rSzl0hd035FrGZWgdv99gddb+Fosj9PJPhOALXyiOZUmhakCfD2+38Hh+3fwPS7+
xaLgd9MgZsL8AQqWKiAHfvzzKQQo06dkNMUZV6XAvgFPb00Hxrji+T2JZePkmkHNnT1cNY6oTKRX
RvtY06mZ8d6A+ksf000TcWRAx1mifgJi6yVfJ+v4mm7Ph1s+XB310VCfLYR0cSpM/lwAbQRBYt9u
HyKCzcu966HQAc2rU4easzyuCQjOohp9j4cirM4sP2/bMBChg14quGNkAus9CDgxQdqWse2JTMk2
ybKwcBAXOal3eVMr4HKky5MjcKyfCMBNn/LC6TPd9NFJU8fTnFfK3FYnE6oCsuIDSMtt9ZV31i0a
bjfGekS8SEOyTVlnAAZQfidKpCN9SuF/TkF8VJLMCCX4nwSLnjqS7WIG9U2V8qhAQfgFDo1Dn/9F
6uMucgcpCC/RXvBZJXUr3KFG2ZP6lRsThee4BYmL1KHYwHpOn3bD8rQaaoo77BKqEUK49ZR97z6y
/59QOQMnCfV5MdyPoTDrVWRh9Wem5GM+GDyanwREX3K1DDg7m9NqzZEY9/Ry2SJOa2U2V6ih0hX2
ya/RtMqfhBHU6y92YzcnwX73e3g9hXmF/2blVGTDe4ff6Wco1MXDtyEYNuPXoLPSl2oSev3uqGyL
zDXed+F4SgyfpO1T8xmQi4QEe5c2jPRlzscl8BjzC9bijVnmP90hV3GlA1WOWhfXJlkR1A9dFW7Z
rhUpNLmBQNwd/POQr2A7UyqVxBWipVWLcFItu2lOYelGukI4OdP8RU3VfdCijdl/kYfRqDhq0r3b
1CkwogRg2BSfjV98NSOerD+mWjMyjbbcBCD79EG6D1jtGAdbT4m/8HghDmybtT756okHr6R+qHvp
twQU3NF2HhO+ufZjTFb2y/qGoOxGxIWiGVfDNCENih/jsvbdzxa9fyekqPlFobrk3APPz+XsmGLq
zpxiu0LEO6fLUqLQSgjxK/QZUHwbY/ZMEK/oklJZyO+Seu6JOEGYMymRCwWv3dAxWYjqw8cOK+22
GLMJEsV8tB3NyabZdsUR42royQMesX7UiByYKkNr1s3+8FxxlmL/n1mFr+QO/XHYLZ26c9g0hCLm
19S5FcFkvFHM8qHVbsEfKJZ6gSJa0gj1A/Nq2P0WiM/YrJ1KEA30eSfiaBufNWhqimamhSqYFNAd
hwS5TlhA+dx2Vk2BG6kHX3v7cf7OSFMCrLGUDXNZGOueq8alGRf16DZONOYPUQrzFNryPZdSoGis
Y2sdkuaRfclxgieoVIXlrvQsBC5XOXAzYFjQjRd92SHmpU7eoytK9sd4+SuTCCo8xAgCoFsWkU+S
sbbAvdOuHtkg2VG/VRcx6rJKksWrWtljyhS8WpKCy7gLcFilXS+Yp6igh7WuAWh9rk1NSemnSn/E
1Ljec7hjxJZzCQsw9VWloqHJtcaE+5TgdrqIsk+uwqGsLnR7xrDw4O0aONizzs3+8GdQWKo+1+zr
CZwpc9v+QveMueedh6WfPczV8+A8u11YDYL28wZJIsyK6LUibcFxuarv7dVMfUu/TzAwhNhCXW9g
z8eUSza3QFxgYwAcLN61phFfQqMAeWJQrOTDNzwaRW1PKAyfUrLTaD075ef4AyYEjnPVle2F7jK7
qokiTjPe6uHm8B1Vcbg8GZ1J9ihSnrwxLUuEtZVHoEod/N4cl3+I8whqUNSvuk48+LQEjbSTFupt
bwUt0pF8EVzbEW/87IS4RZmKJ3xFi51PJ06nD+r+CKLXg7uxOEuvBViBeoPtY19GZhyHIMlbJGpp
XQudRT5TYTBaf5AC5VEN5JVcklZhJJQ7RN4F0Phvm4kE2GlrGKtEKZQ+vxR+kn+AlocD99L71Sx8
wdy0xLFqsYocrcDNGVHeYAVVU9fKyokIIW+nDP5vYHD0yFPFKNr8osytoyxSMuYfLsqT5+7aYOe7
m6opWQb5B8P+rK8O+cFE4lsb3X1sOmAh3zXRUdadIOQrPYDAAKI+lot0dec2y3TUH2uuV9AQrYBi
Apd2STlxSeKiZL6dtv7FmpWKFZoeLXkx7LlS38CBAAv+bWGcYEwQJypSxM+1D2z71EgPqNohNIi3
qeViDNR3d/VmFjCCcvErDidq6BEmaYCF8ja6m6yXWdPuEmGTtq3PaOZSyHTWbSmdV/9uuVeJyRVs
DeopiaxKBt2csx/9n8/PSDvjxYHsnO6AHBsmU2Hpwy+BzS80OljISF/+HdirUITBfFYN1jXf7rIm
6Ma8iOtInT+45MVRnSqDZtfl3mOxfg6j0tTaNMP1P6EZZUS1PeN2likYmiriXbAKQ3Kmt+c2V/Ld
WnQTgOsrR3HNcj8efI/3ccLBkeQQYdnBy3XPk2EkV8MBYo2pQB6ahgFdhLqSSryaHfJ/Fz24oKRr
xv4jZbaQWAtIv2cgfa76BITJa45NGUChz2B6VqsgENcRCERAQ1PN8zq/YZhNEnA8F7pzRk7efWWC
ruTJmLTUtqOMR2nhm2sHIWtqeBiWHJHdQLg+eU8WuG9EQ3P5gf33+YkpON9h5SYr6xV1VVAMu9RT
fIYi8TKGyTfHYmlcg8qCOdn563BLjVuYz6Yh2/Iw0sFR3cOJGOLl0extCYHpxBLOcLjGYlpuv4vy
uF/gCrRhUXPSA17mqIoOTmNG61HtxU4XO8Enuf8Q/JgiO6w8EZPAKfnlWtD1XDdOAVKeRYbXtx9h
VbyyNmVBxwIl7OxthY5ElVHSYvEg9XxQmLq4L8dwe9uUgxY7jFwn6kyyC3txPOR4Wd/TeU3dYI9b
ntdLf4ysOdmV4RdDE2nXpSsldSRBBq2j6MYwUMgH/QRfOsNEcV1rnAlqzoIz6G7ZTbP3XcbJuesK
rGWqHhNoaQk2AkoUChdPbaSn6ew8VkaAJTdS6qdmNyDnb1fQtnG1IR46aLleUajeIbbATwnLU6d2
q6qN23O2jonQEVr+RC93NvCJk9Cf2VH/SeZZnvYbIXfkydvUhAVSYMbn3K0Xmy8fGfANpJecyrw4
9R3IDynJPspHWotZ5CIaXYoI8tRqEnKtP/jaCOl0PCxV1KJu/v/ODoDoyjIgrEZB2KOhjf/0GSvf
f9qhnXaehfIJpV7DmtxWBB0c2dPnqdARLrHph2W5eOQYT+/qo4feDstHKuw8F8G8B8FNHNC6UbvS
E7jsEAeWQ5LtwKMlmxuM/oMACVe8PyfCt7ees8DmaEyx9e7Aqop1qNcaBfIXBpDW9PW/VBOyKxOo
IPDB4ugLxMv0KkkL7jB4OsuPbu8pbefwzIy2TORMKJIXG6STTWqQXDBktLkYV85Tw6qjbbaEFo0E
v8VPHbkC4VU3n1zY0DHEO7o6rUnzCCvCY0v9k7vRPHzLwsta9KLcD/woAFRuIp0Fu3oBZOnfLGvf
GvWoFj48jFupc+LOGpb84hj6IwtJcSfrOTou5wfWC9SkzZsi9JYN/2nAiqSGNU3jDygOWIg2Q93X
1i81ckRtfpQG3ybPXK0jXROKOJ+I6A0E+zIFYOpKztMLB4jAJkG+0TlrUvUG46nprzIeY7tX7w4C
cePfvOWZjNjit+hJiMjNMiRwUwBJxy+TgBWfYtuuNoXrSGNBrPWcF1+0VENS3/okbZZIYLIssMVv
WFAXGR/iCWMiQs51bxTZq/O2s3BZHmO8fqj/HI8pMRfEO7y94MHnbdkZYH49VsWmS8/A6S30bA9p
5iZVAtSykqi46kgNiUTM+SZR6R28/f4j/VfU5qmLUTePJqT2cKKgQka2Mbb5Ncy6V8iNo+EGXcAL
4ARua/42R5De3vbD9OPbnrAeHPPAiElBQfrz/V3zcsovVJ+caRkqy13u5Pyib7rYq7bkImoeLJY7
UNsWhC+dBN5mXRUXnDnzlyCHwKSQ7jYPWKB2MvMN7ugMgBZk1bUXaLp+WsF7P2UOtcDAEcszRTLX
sZkfFPq9bC0UDBrE+sxA57IMBRZkUtLddkSe3iDkM+6JvB8Ju/2E2j70aQYErrtse8Nqr5wSGBhE
hszHDLfeNC2DE7NHS1kEQSK6t/4irDKo5KpZVm8agkoHeRCIWZPdOIEbjmQn5HcYIy/RKnvazsgI
8ofgV6sqkcZCczWrjm0SkhIMyV/B9B+HWLAUr2EE/1eOn8japskInKzg3AC/Y4LAr63RrDSzDeeC
up12Y85zQ6xkupZe3JR5nZ1VfnxeyMlbEmTScT6iVAHtM3CnNnu1wwaNMS9KMiiA19jgKMt3m0LW
whOJ/OjD4/wSw3btGtJtbeqR/Q41XB8EgCLGuhctcVz5By+RCfZb70N0NUu+5+XMWgp3PL607FpE
QkzRsWRCCsvn/IZ4CPtO1TLWvMz9Ru3pm9NjW/t/TD8RZcqiz33q3/sIww4hU7oq58+KOfk/PD+S
NSTPWKhbKtrOXqwOvjR2eMxSAdoDteoGYeuo5+KoXn6rxd3AXj1HjUFLvyjS42XpZYlbEhCsygIB
Xij757rmr4F6PNs8TnxeSpu/43pWtsFXCiu7y+WPwlAj5uGMXLwSiuJ3qSBC8598+4emGKxoPIrI
MvaHzS5GdLO/5gS7Y7QSxfYdWnW1Vlq4RD/lknLZYv5RoE9sN7pp5pSfd4ppVNNPPP4dvCYEp1zm
I8/3UEzuIqFp+b8MfpIV23tej1e8BDDr9Tf3Bge3X8dleNh9ENcFi1RkbPIBxES1Lp66gXp+omfa
ZNubK25gpsZZXUmWG30jZ0Rh70hEeMB9O9XGI6JAoJ8S6R7gT4kiL5i3NCHbGRnmJPmb3URdEl+M
1TGiZGt47a9833ypL3mR5dQ0/n7A/KLw/ZLc/zVxjYrgKZ7/K+e+33PE1HSzKMpMQgYPB2aPgx7x
2ZUpM13V+O10NRL7qd4rj53w+atkvN7TyA2Cl2Y8/9TbLNAq6uZ/aI9JUv3zA32hZMyBM7LeXRdq
BAfgYIWbFoEuzQU3GNmG2qHH+yxS+dqyuT0TYB0uln98MgU8FDT24XhMN3XwHffd+pKN1Elh8Eml
IOm7U9RyToGNzrPKVBPecJ7PLWsTBFkU3CZ40lAeJVri6X2PKqAVbA8n8Kd4wzZPwGCeHCqiE5pi
nHdNxVtjmtuxkef7PklAQZxU+qZgHmIuzFxWtMqokw7kK7c7IyaYcTV2+kcuEubgklwBlJg0aTjy
ZML+XQq3vzibklqhIHi7LYRSSKelatemK+B4Egt6MW2RpArCpk1w1smVw4MFAbKcCMW5t6Phl2rW
VkMeocGgitiruO/+f3Zo7wlIFPun4WsOy3r/COKEb2FH3rL7WVfOf2cOOsuy4F5X1yNf27cA1WY0
t6d+RKW6n/YOFL/FmoCdTDCbIER8xzNfCN+ZFCQzgBZz5GwW37GdRMEUZzj2fymQgSXDHb31hQCb
JGzhGjFsjGCEDhOj35R65t6KAv6TtAcCM+QNGqIWZIgkzyyxtuF1Uapkd0iV4CrcA0Zcigt9bNqj
C9391rKVUiq0uWdtRA5XYSzD+lWEwWrU84i1JKR1BB9p4GLePhkwOkh6BrCk/LYD849Z4PbA3qXM
BDM6MU7vJN6Vxb1nve0ORDtmbUXWvJanHabUKK5TqSZf9uvXof3eSoEHGSosrX25n5lAfa/DgfJp
M07AcMboVA0agy5Auojz16jKdkyHUXOGFiDoGNfPhA6He2i4+GX1MpS1srBp/cJzo/TiLAJtb3dQ
k06WnkX6jVGsKePhJs+HUAHr//ZcrvD1zDWBLVHlmGjWRSyfq+begpbBJ6Shl6tZ+kPKcfgsdTXg
Vv35nrYrFHYN4qA39fWVsjgH/3fJtru32o4RGBDeIVYYLfVSiXesbJ0PLcC2SBiZMASjdMrHhaqw
xOKNyWfgukqb8DgKHrDzxYNCVCK6T0fsCGVsnTVFTDUZfJD7XYPBeUbHvH9tPuQchrTmfA8IDVHY
ToPN9p4DcJn5ONcRlyL1ZMdkMj+MoSDod4s0ydm1lLFMd/4Bh5PegOJeuX4AsLA7rkxYEO/oTdtB
REhtcNTxH/BpgIOWxQxzCIEtx4XEJcvukNBCePT2+Ad88uaM0s9b71+gu20XmZlE/xxBq17cVmJn
O4OOGUnqVmQbdeGnbT+oaxexUtpua4zIhwQlzZze5D3+zA0M6bVmArPkYkwf6ge1OZMn9Sa+qQ/y
lZLmwEYSPMUCXgVThd7pJC0BUoXJHn9BBtBSJcA9FfBEnUxH1P0kBAC4KYNX8uuIxHoTVd++nsm3
b+Q/n5APia2SXtN+M3Aj3+SM3c4FkAvn26bc97SDS3UnowLa7b7ZBAd45uFlbbuKO3m4sHIBmJ/E
QA7tLmruVVuJE2Dhk9f7gBhqKHFL2UQQ5Ci2YXtgnXvs9EVkH8WJ5X3JEfO3fgp0d9ryjJXapgvG
KkNbb+3sYM6xXUiCTXHu5ULFVztloJocmB6jHtQ4pAuNxdZvmCE8s7Ce2ssEJ+wLIx9f+cjTTOyT
Qtb+4qO3+DDm5X0J33GMQAm8RBWXYq0F9GY9L+t6JzcpPFot/x53SlVCX7+32nXnEygL7h+fEBh/
pYzXB57cqc9zXZuZx5erm4iqnhYsqFvRrET9cw/gj5dZDK47yu3T6+ukQ0PDZpRYN/gGcWMozW12
pwYiUrVRIyZAEwwFvZTSoGYhT4XeeTTTvu2DoqDK3Za8SF2zYRXBChzYLkrvtPnKnf3xksLh23Ld
EWsCge0ww80rpdx/u606EBZNUv+0YePgsmuQNRehcMAZCrTpgFjhpz/srmNj8sKVy/Sqd3CThYXh
sYTGE/Ae/7+8KqyGQwLmNYPx8ap1jmB6dDs7LnEcy2gxwy0lPuJ35dKQUOBHNFdipRS21oG/AekV
326Wbei1lxgaSv+lfWGs3A3GuhZIzYirHR3oi/R0kwQu1/1TkQJQaxFbMgiUGDrAIuE1y9R/Q3Ab
F5wJETWdeRqKRnUqmdtL9rj/vtRT49k3EvfjBDPt0KVcnG0+JHv+WquV+BbgP39GenJyh7Pt77vS
LsyTi8NtxDPdluvSnTQxh+M3osf0iOHoIhaooOELfG4j8UykS+6uabOAatNCFrPg8MRJHvVfjvJF
eW0qwmOZdd3NNL5ZFBiaWXP5oSZoPix74GPcRCMKurzesZZFVSG8Ds8gwHh/CInCf4y1uBAyO9zM
S3GABbV7Gz3ZdGKBgOHw7xcJrVd+HHBU8glg6I+Y2Slk3RgUvUs/hw86AWs1T/fQ6y3Hmav5xdRK
Xuk3Ls/QneNvQv8zGdzIBgxtJbpjlUWG2A10URYQLttTSBa1v8mM0GSX1Tz9Xpc7vQdfSlzEptuL
JJV5N0j6IfZZhN7GlvKjYQsycKy0dcV63EV42Enun/sTecPMEiNGeVdLTPZ+YmSFI+tAEe1qugr7
vscAaKjEgzXzglabMFQiv44dFAkiEhkVRRp23gp4o5dpXvqqFPYCfuEkqz17SJML9lWnjLEmmv8o
wBHqUotkTR57Ld9hW8gJUzBIZb3J5uRtfYq+Dv1xLekuxvjd7UonHRX9Z8TcmCeoaN0DWy5/XxIG
9+Vw3exF1K1kSjgJIOW4StOfmTqmn9zkk7Js7OYrFqrRUsw6j3yQRP2Ih+kXJLKw62oTwpoMw8yI
qYUkHpvD8hJ9kMxlTZgcVLF7CIRUebbOs2D1xBcuzmziDKOan3OEeubOZ3tRBcjwVFOqkmR7b04+
YT2BTjglRrqu7GQQ5s8tJRN9ZQafmwiaHzFw2B458KBUOLe2D88efjLxl4acm8NxQLbvHACK8aG4
xIY0QTj9nwKRFEExJ1wQMY/1oqceSkDwV5Mqa8lx0GVIXNomJcxFJLE2pHCf7IXXEoZkV75NjXth
gI0YI09VMQmsgJlMFNPXgomiOeohuLZR7/h5PB06OTBY3M2ituVD6rSDJgHymZ/svffVQtQjGKm9
6YLyuE0O3sEvVTPoKoOJlG3i7o3dRILJiMGTtGKOmrPjIxWxXD0zSeuqoIp6WINjlcnUNNUHO0WJ
8xNve4CHtpRIJpUYbLMh7u1dReiWXytFcEY/EE3DqFDoqhILhVTGartIJqu7H3maNyCSJMchW0rE
bNYVkT6z86kuUd8dZfxPtAELexVS+kswfgLVlKFEZXpiImdh2XGcgJytSDYfjHBD5RNONEYuLuJm
yY4Si+sjZEP55nklJSTKKNS20GvWQjW69TiWQkZn6NqxbIEYVS6f+JsbgBV7/SHuVmbR3wEh2+Cc
+pIEQTNWPXljkTXkartFq56kDG7T276qMN8cJ4Hu3K8iiFfy3h+QnkHvnOMVyVshDlBCvXScAOy6
xPLGkFjjqb24eXDMTOSIJ/SyUgNuFuaRMlA7Rm0AA42Ubt4qu1Ag0iPJ2b1AM8HsZEwucxNxYAlQ
w1R9Ss1t8dmbwdni9GENfPJImLEZlbLNekWWkpLTi7BsZFkoBmlGGQTX+xc8qK8QMWdV3IK+AtCZ
WjrN/fBdyJasvoCnF0ip4oGHG49TPRV65gRuDSdqnI57dhTe0xPB4esfvlcPwvoAvlHckVIIqhid
Ft7a2jGT2WVZdzp4k1YwW2ccb5DdeyWS+QIMlV5iSAKhMspcKIuSJcDTKbC2vzOqIzp5RqlOiEyL
hkictArlqiipEGGxJ5bs8ZRIO1KafH2uqD8AgtJABmifPtANTYWyYxullIObXF1eThOysEql65aP
0UH569vSFpM0uCSShlPxuMOSB6IcPwtYcqPNg+MwxDJryMxK1G5sT/lnU+86VbmT1Z/EC143djZk
DBGP9zR7YlZ9n2zBmCJa/7ktlJIUNJIIiY++yKhI8mNflS1ZnPfrd8CfZ2O/BJ1aoa305Px3l4jX
VhqrmaPLx3s4BbKt6+ia6Xhk4JXvNcSEdsXY0Y5+peBlreb0Ujjdf4WNBVLwb+uOTE7WZh4TiaPK
qguYVJvjtGGo0BjzUu0xqd7RSArFVIH5mqQDgUUPN0lL2c8V7e+0UV9I+/gsMEWgD5uCVXj2CjAf
V3sD6kn6qPhky/b7sz7B2V7Rl+UXeznsQWHzIgyEiClDu3HkMQ07vfC0yVNuzY4j54ebkI1QPE/T
56cxjfaX7UrzBS9f073IbXn1g7cP3SfNPGyi2DrgSJ838x2OiUGXGBROgwndhuWwRrJYQKs70INq
4ZIBZi/fozelgJcZw/dvaAtXNB/S1HVes8BIJIxfv3kzLDutgRmQbgGDqlzZrt8pU5WgxKgpAXjv
7d1EEnhNsSsSoeaL+bfuQFgYeIRGnZYUgvCtb9G+eF0CigeqhYL2PhaTFS5dKse4JMW2+t6DVKxW
QLRtEyJ/5g0RKVkyLx/eLZTyOz6JYbWLbR+S7k4ndJ9MIgBbEbhxmWZxoouOl/+s3DB1EUa424pQ
08sGCWB0ZWoErceKYJFy8VNu2Ibg2RC2GquWmzSaAZ0A6uovJhngsyD4w95Zs44jsDvPel4vFsvR
rPGJ8o/IRvmuiHFcs3h6CMv+eNnMPKwChh31R/tDB/KQFRo/hhA64d4VgYAeKnoN6hqKNK0to2Kj
Cn5rANfr6igHwOGrne2WSA3NDMQlng1tieRsfoqlns26oW3TiOtZMPFASfC36i+R1lET6YLZcDhd
LMmG4te7ORQbM1YAILLoU1BIdHsGJXxUkXxgB/kfgA7kXu+eW72/nuFXMILzc0Fz/ZIjo4GhHfuu
0unhiOox1qKihKXPR3eK24kTmC+Ev5nGihZPGbvKMuNLNCtJ8y2zDOAB/ConKHO6sQ1ov+3Rq2M1
Mhln/4SfZfkD3j3ZYB6c4mwW2HwCpx6kKCQyv874/JDWFZmbXYQdbK876+eyjH1p6bc+ybZ5TP+Z
zt9eKvutPXjeavi6zc7pXuZRuJa5327n/HGsHCTVE1xRAv5GwCBIz4Jo5NJdScBCwB7Dx60RPvCR
7sZCEWZsLLrJEq/sajYVLxiaoq2J5sEQjcnCqQ+JiIrPdC7OukwU/bdqqmLfgfo7CiSSuHg4oLOT
V/3NQGlf5WhU+e/Ujz1SnNuSczOTLSNpxyptmhlL2Uqr9RiOxrqY6d+dedlUMiVDSpJV4WBUVX9d
EdZVCjVOO75dVHb5ViijdvocTwPLAbqhNS7+pzq36sUqkAnPMGrBM8sh4FtXB4P5su9qZLBjGzDM
CDztZHPJwERt3WR4BIcBv6LRUkBFh/lUBH0CS+oJjqVQyMcoxWHhEcnxGL9oOcCiqjeFpdSB7aPN
0kcrjcz0D935HMe+4iPkzWJoMQxGX8yFj/p6SDDPskngzcqbxRxVlhtncE7h+TuBEV+YbnRq95PZ
bsGpPW4d4mqwlsPLjsv8Ie97ZhrOWm6nVm25LaxS7ddnxzx3VWw3MsLUx5Y5iyY5uMewTwGZfxNG
4Rsh1zuXTioS5VSEXZ0CZjPzWqFEzllRgt1POAPe77OYI7ENhOsDMq2ZocQBcaHUVEXTd/b3PRhq
RMvhOHFIuCnw2Z70ZSoOkDf9B06FgxhrvdUaCUUNp8XP+K+a02lFzAdelozX+C7xD8gKVbJVV21r
xdn16VO7p8rFcYNqVlOdG3g1FZMNSROjEaVVReI7LSjOg4w/2g5JDfnTDs9bhxshba6d+91fCyOr
Ji7SWcM2IpBFvRisceTPGgdXFLT7HKpstBnI4nenEAOOqOcPNBtFf8+gA9BI2nDQYfNEl3Cb6Wdp
nkTasxdu17G91KSw6ZgyDNXnSq9B2Bb3dOmRjMKnjKjSI2MQ0P3gQLNNC0rPAb1HIAaD4rrZ3Z02
OAp8VFM0VTuTpoZwEOe7Y6gBAO/dvXpXLbOUXOcoegpaOUYRM5vwkMAvR4H+unTIPA7WmQtk9ygy
d7rWC9eFsEHbRTv/o0jncEmUWp1J2rXVRynGS34B6ORYv0K6BRFznH1Zivoo+cNXUJu72Ixmwz3A
muHbLrHQw4iOjjp9lpGs4QCFY1QZEE1RJBKc4hZKeSrMSoCugCp26Bp8I3cxcDStlNyn+RASUVoD
DkCxZ41eYylhxOZ6it/rKfl6oyJ3uZ1ENTVPICwONi5nOpHanDr85UCfjY0iGJG4C450HkxkNVR2
XmitiUPYMdzSAuWmBTjDei305sfsHYEdPLl2cRVRm83NF68UizJ311muflsiJM0dImemDm9V2ovp
nopvu+Av0p527zH1QuNmsCyn6n+wkJzT/GrVmqJ34ImcPhKUQ90unPZXYQ2wSTFzMMWPyHvWpMKz
EK1ny5y8x24AhxK+Z5Ua8KHWwkeO94bE4B+bPwiOOW1A4e4kSXZiL6/o5b51Obw3BDwg3XYggMP+
ielLBXhWQHfBmjHyEm9NFcsaqlLRYR1qnbC1OPK9c5XLxWsiBjb39BSu3JY6unm0rKnsB589nsM1
6qSfZ4fsBR11GIkJSQSfU6VjlglNh4b1sSm6LlzAbHayUucLMegtpl03TTx3WEO0gZzjDjRmOW4K
8LCGnq/PIZ31YJLzPaVK7Z6DGBzkxRav0KFjFhKzNJFQ+r0UCrG4jGh3r2Z9/jPLC32fWJ+/roq9
GaMz4GYtyLxw03/+LVdGRstiUpwvN5h6qfx4JkqI5CIWdfZde3c6ly3FAwCFdauYSTVYi8jTRmv/
sh50/TQjTGZh5+HYj9jeXJ8P7otM1/kN+gcNZazgLiD27zXzJb5UHwHfTEwrd9JeDArVxvBcvx9S
Ter/nWFqJq+OfF2AjT0ABbsy1WEockTxS8jAMsFMDFXbzoesUzUOQOj4COmljCJXFjgZbbBPIcUa
D8oqwBqvOpOwqA8tG6F6h7bX9AoGOH76DP4WxuXoqLRq+QzZXENDkbkee69PJyiiG+TJf561n/qV
pa2Pt+5WTfw4PpsqYVIG+VU0bjFlO57UyMo0qphVqzrSUmudYD0ZBqOnQKC/n8Y1ihb4oldUtCty
sUSDfCMl14+5dhvwH3hlK07/pXY6H55rkanPQJqjKJozxDw2fCO5YpjJWBPHDcxWT60kiUuJKSM/
Q13WM9nI/sVEmxaY4iMRI1FiFAVTebRIzth4J7/qCw81wmjXMaNqP26p3iP+GpJBSpUrLDh+8Yt0
f+hhHITmjfqpSkz+RmIFnLZv42J5xyg4CnvCPE2iLhGmjOHwQE+CwtTqey6zpK7YAd5SO8Cfebbr
7GGHdjGZuauWu5okWgyT2geSYEa3JyPDFwspVX7EIVZpagh64erVluxyyEzU25SdHzMScfvs8iE/
MEPx4yjvYk2AIpsMYTEuTuRO8fRl9XGHLIcNUKXp6v19bsCDG5C/osjMJuXChO69mMiw2drRfJyh
nJ5wXTBTwOwUSxpWk4qOPENxjplGPEuKr2104LGv7gX4dqLa4RmG5ud55EU6fnik2Sta7eZ1iKis
6JOXlg0HpT/5EcWJcDU8rUwCaJYlyaF1mEqF/igUPQK1sac5SxxuZayfqtzNm2ZK1Y6RWExbqXUL
If7zjuRwOxHqkgcgOGM4WlfbJy6pREN+oNZtnA7xlvRCxTPxH3GwCYXu2J6l8lRmaX3zyOLUrX0N
8CNuQj/2s1R/AyN3Eo0uIRtzypZ5NObH5GZyqyOliLOpDlJ6/gKUCwN6ZDUK4fZUw8O4uG50pQ3M
dINKvoOyHI4EL95PMEOcQcqcRDGaoNiGrtiOqyO4uaAlqQPVdMhIJh7D7tf6kMFU1lms8Lu1p/Vs
28tsgSKOCnMOR7dKWXd0hvrGKEljQ6wV/E6Y5zlxZ9pw6szB61ghjFf4tmysg3BoTQXo7EbLYesn
+COPcTb4RK93PN6HizxoPBMLoRuuWWgWMH0jTg3C6mYEtDIj+Oo/E2Hcqc83E9IfT2M1EhZ1B59G
tCTLbFn1IKizJhj/+FBBIvvDNKQCIv4V5WcOCilQ/uMUxKjVOngsCEg5qhpdkvdvjL8cNkRAYmPa
43vWSlhxyOKvGXFbRg9EkDyUqfM4+WBUJJrYte2KCkPiq9EwfTddH9yJ3MkMTdaCb7REz4dnzXVa
ChPEVGI+0PpBZa5/kXV1R1HSjQ6iE0MlbMOJHEHggL5DoJQ2fD+MH2dVfymOR4Vkba7zQNZ8Jla/
23dhv4nwGWGcSkPK83r8DKES9EtDv9H0jj5M1vkVqt/1Ae7WyMn3nc4T9UFqP528d6QvF2ojGQuq
/43MqXJwIUDfeMZBIyRQ1sPrqLVSES+MiWIW07Awm/l446G5kokMRT4NUAK5Cs73Gz7bUwAadIO+
I+GLu96T9+IuaCOpZJYtSKsVem6tVHi67Nn3tsaEigW7OCCTMaWg2EmN1+TzFEyTROJ8CzDqrVrZ
KnF+0E+a6BCt0uzhrZP/kcnw5NWylY4rlvLdFKGhQYJTBWCSPV0gyRA5uxPx+oWrl0nQKjEBu7MF
vowjbaopP3xezNJ9OOASMCl/u+KeddvR1crN6AktcZldZeY39sd5Dzo8dMoyqfia4RU0lBPh448B
W1441+on+IHkcl3BmAz2Ddzxnh+0dCmbRSmpLxtZMqHdbg1RuSgLY59/94YYE6e9/p6ynueSUJKL
KRy8zYlbWNee3TfiGf9ytTZqxaLIu1GLTHYopaDpRWcg6t8JpWuyGYvKvaCsR/q7/6oLxfneOKoX
RGOitqvYaVi+P9q0mAJKzJjg6WzW5wMWz/DzoUlGZFEUPQzbu91k0WS6ePpdGqfd8xTQXafvcJF1
55Sd1dO6iuJ6T/PJFIHaAwg0LSOMYHOPz2Mr5RpZkbbS6Zj0nxw3Gb7mW2ivtNTl9C+sKVmuhPyA
yauE5ruKmiDleki7sSUZTvL42lPA9lIsxoJMQX4bRt+NtYxVOaS9hVOMUXRW/VWJoBa2rZOEfAZR
ggmjQPxtifzxNr+QLuCIdkDbtgktel7/gi5WFamSMQ5ZZw4CEi6rJC8KT8xOQFK9lVYCsA0nbO8C
Bvq0OdmzazXNdEH/cjo3WTj4E+KzTjNZEfdqHq8ZyvJWuS+KUHu2CTthfdXnIuNW3iREPbhNFEL0
aZ14zCjyfGanIdXUSxYcmb8AFHsMM53nCWHmsB2ThxfvVdGTj8j5/LPI0lzP0OJRrV2IfHgLCxlG
OlTBWBJmjjLVHXZG+h5eKwIhgz5rXY7K/ZX4PRscV//oUA9l9ivG/DsiQkxMZgjF0O0mElynz/Fn
nlgfBwfHGoL3DOUQYJIulKJn6K1ZjhhmB4rm/DroNQZStyq+RWwA+XfHfvXEY/PAzsitTAJ7FP3M
Vfjdw+AbmBxbFZvN8yxpZIrYhPmUgo3fPNWvU8O8wG3bUL51/XGgZgxgAZZwODGuYMJE3vrTDhST
ON2/dO6hYN7Ih+BUMTN94QXRHutMZLxyC81po8UQdXwQpOA+CN57aK/PTy9N9LpxQ+ticqK/KVSi
0QZ6fgrYJVPL4FoC9Fm5K9aYlC8FIX2fR0fN/y8BwzTDyKVH4ZQWo1ea1RLvdJY584i9uSUQrQPO
XbHXl1IJYeSKyJtwKgIvjmn+X9BjP557D+JCe83g0UOezvo3uNKUz+LwJ0FJ7+lWAcHIABUS6V8R
E2tkSihJaiURXcfn2G0L9preKUL3tILmXf6G0BXKV/5at8d3UC31O5KtTnUyzdzs1edZmuAjuy/2
G++xryArgDzFHRYlazqwWrQ05/RHTsHRMlwF/uQdAeCYONccm3HcTPj8SUOpcVyd2mVcikf1mxTw
kALfvmzvRn+X1fx4SM0X4hsi7DW9kbM7Aex0gzUIHrQ3wd9B1D8cONw6jXNVH3BU9Xna/EZeOZAP
Nw/xb9kQsE95T1Xbn3zBRtMrn9Tw4kBeFkyTsIsg8KAlbgdkqtjCqOGb+x/gBEy4aP9V/kTRI6wD
TtZuzpiUrP+yjSTlEH28L/Ht6Kt9X5kQigNAZv8iVykKrwzjCshTZQI7pN/P1StjHIDZ8ZSpuLii
w3MrjXXtm4RR9jmxJRX4KuSk53OjzyuC1qEpk1bNNnuH6YlZLGdCecV+2I8uND3aWZ1ejG7/suMk
WPKE+n0FIjxkps2d2ezUnGIL1u2Xsw96CXVpePjhQaq97q2N4mH2nt084leE751kbVWZaqfLuqW5
b9SGrge5AAXvfBdixuLRJf2y3FHjQvP6nhkenTUY1x407VI9W7/WVhVM1hFzGE5nm+GXFCKAe+/Y
7wTnF9EY8QgvKk2Pv97Tn9mrG6LiVTg7GqhUu71DhTFNoDabmyqE4K6E1aTjc3qw5baFmMCmk4A+
iyKw8gZhfqa9ZJsKuRu58eICuOMEH1MyTZRVtBfIcpOUfbJiQKFNGUFMloMwpr21Fj5zg4vNH6a9
mkwnDDRjsxYbW8J54yzaKFP3MHqkdWfOFihyLG1l38oEVsS190lJHQ0+fTUgZJvMaDLUaRzCCMSV
81qGKd42b3R/GAjJoBQr4SuF4oLVOyEMEq/dnwUnjU+jMK8xq362DmvmQA/YieNjdn9IJh1x2tvV
NVJD+BzvV6g9O84iLxSbpJ2bky2aQjerX/jTem0b2iW71kwAAE4mLrInNtR4UWCPfH9YrZwvFpyh
sBVAZJHzw3ux428JU6s50jIrXJ9g1ZlKHXBgwli2dqJv68FlMgrvtd+HO3dYX1r0iGoGtFC2coXN
XWDIU+p0hueb4LARE90GkYqu9LrSH5IKborZ0FNx10D/Z5oosLNhhDHc/zmMVUHM7wof65KrVoof
TLBP1yk7IESudJR7gFIex06ITBBOJtjCsP4CyULv9LjWq3u+1W/7d8ZR0YzOR3LBUkglJd3X8UJv
AqgO+vTtD9KlFODDQag2PRK1DjCeCw4Sj87PGK+VOSkSF6bIjg+LtQ8Za2z3KfLD6XCguM7UHIZZ
yz/TVJbRbtTRJfjKEtTxDjYj7klyflltx+2Pq9PK558ISWWZc8ODyShBzUa8jHtOEHSOQskbvS0u
A4EdRAgmEj8tGBru8H5wwpzGPQjnMM+GTHU3RO+rGyc9UW+EKuwrbHA0ChiuJ/eBP8+U0mOCTvFo
omQRQlRyjlVfMAYUGPqh1NO9p+ed7Jvqh5mgNRQEJl+3Q85fEvJ/o9IiicgUSctP9THvBTrxvtEa
I0pknj+qMLYmryIvcMyFzTMu/HGKykYvioUFWw3Cb+G+jUsfjYR1syjTtKpzrvt6vC6V//CnCr0B
tiWDblVWL4qxHepbA5SFijffVFJxWYzTw8Cm6hknk8jaSWG+IIXf75DwfIvqGZOn7K7HsqPhocFn
5FCp8UHRyuutddPGrfSRq8JVYK0rar2VXIEkaEq6vCH8ON9Hpzwh/1u2yHwV/05ZR3FS1pjhSE91
jZ8yzaUGyHpjHxsF3suZh2mzPudAYUUeeJPowzqHmuiyZu0806Gps3I0/DdvJPqrolwO8RePNId/
JULZeLyHxtLvtuAlNVCvFzFsusn2dAnAmTYX4EYzorfZ9EnviZ9B+bDiW39pR627kNgwcKzAetvg
QO0XE6hQA9FsBQfdowKSEDweW/i6L43J1dZ/EPaS2t+wNmpK6kP6/3Et5hleaKTKU7Lmi/Dg/cjb
65uBeiQ+RYKG/2Il422wtx4t2QoCkwfD3bSapx0bSsHdot1rd35oKTrKE0R8hwCgEwLKqCLL7dPJ
R0ipA+11RVt3uLcIhl5RNTGlsiSP9T9Sc23Fb6bIyUp0Cz/h4HBz/x/IIofePTQU/uboIeL3iZr2
1xiN/JXGVN5Tpp9mFgoKcAx5UCfO86kPav3ZDoE9ZTnVIIeCdQ3sIzr9PNXUtJH5nZ3JU2Ovy/QU
nMoEBgVK5DNoGZUzd2Zul1pbopaVm4IyPPJ255NpjGHECfUu8bgSSVjVlqRIikuFIFPHYr1m/Lyy
vB13hJqT+dtVs41rK090mp4z/nppL6t2zIq/cB3DRQsBiT4ea31EAN0ICKMpsPFIN/HVaaHtTfuA
gkaI74XWjCo03ij3iASvqvETWOOQc2A1UZLc6O8RuLlO+IOaVq97wtulu+0vQ5tDz4+fwh8ND3mv
nEJVRNLMn0KUfmftBT8ZvRsxDKKLBSpilGaIi+3mNhYwlN8u9zqhQscUkQv1tvR3Kn00datplOfR
HMFSAPkMNAtTV6D/Aom2MnLfZySEtpgou0m1Nn087vIFR9Cs6+OWnNbEsu43qpqacLLkPPvbEpeq
bpkvYsrcp4kOSA3kPIXkV61i8MHiiFhdjF1TxRQwMyuCsWVWh8u5qPQW3fv3v0oSFd5TAGmfHGhv
k1QUZPor2SSWaYixw6jnBWq5EopFo6V321ARPdmWJM4ntAKl9+jSM0AklYD0RdZpdMhoysXjrXvE
sR0tZjbxcOhvcqcspON/ytINmYpEKHI5c76ycuuziCTWsEOq/PRSeEblONJvEu8SY5Ccwyy9l7r1
vi+Ow18tm/CfcJrFihvMM/92EX+HXXbt6SnHz4ycD36OldNOWFzpmWuTvmgBQHgwwGhvEwKqhgjW
6tPkB2MIGCySUNs0Uytz2mehlgcYGev/xhdurU5HnTYluegvWp4gQydEay9l7Gl3CfFww74UMUxd
816k16SpmKvj51NS7uGUkqCB0xXJyr/ndfGcmTXBymArKLWnlswIcs/F3WM4LKJ/ncANfNuccVTV
W5MSiCZvJEUJJxcylOf4HtUVXAaE3esHltnYeJ/3fX7aRQXOR4khrrln0M1bdA9VshSelCvZEj7H
LfKpBtW/7iwXyO3T/7bd5uU1MHR6mjH2S+JkK7NiPMmGYcIEPrWRehz5asyptqumlgJJHyTMN16U
ZLcfp03If14B5vI31hB2HksXfhRkP1EDTGt9IRbhuzcssBovxlg35lWzMOktvBAbcC3eKGMKMpBp
nn7d1EZDj7emv78TYEhST4YEkwVQH7C6mDomLot7WOBmUO3wBzWhYhWPq4k5RbPI+iPEfwePwtTg
7xld7MXO5taLmz9ESA6nL0NjXqhMiZy+0nI5lx2CXZgi/guvac/ZGCLfGHGwKd6vrqa/M4zLZvxp
VZA5MVRfDGXx1k+Eymgys5/BFhL3ERxXKGDmYGbH52Pi8gEWr5fWyWIrPG++2l0oigONHvZa5Ydw
T8yWBd0p9vyfE5uh57lAj8jO0Rb8RURfinnfpql61ppD57vbrQtuSmk4SMQALdxx2V8Q8COmRmwG
/zLXzYxY9I/LTO1xX1tlrEqdu8SntunOb155wE3NJZA6eDfthQSNaQ/li4ZyoFmAamYMMaVIFD5A
j4NZBkIGsE0ILw34QIvbpOT2NBQKIt/k0gVR5BFQPK0mJP9QJb5sJ15srlX9Ft8qHxrBlBg7t++b
JUtRQcr0hbhpJUfcbxZq3mGjeSZ8aRwNTizwmKSePoVv3gTgdFaDLcCh1H4hoT6+IcZE7HztxkeH
uZBGylwBIYC8ybZc90vrcvg1/jVWnmqfHwcIm/OSMN9xtfx4Dy9N8dx9+SZhXQAAO82lGHVXywRR
bFmPEIrJWAkpkBXsWAjdqdqh1yz8x9ujFCjlZYoPsrSXMcTAql+mbBPzifV5zlFXWmYnqpFSv8m6
sksDDDNt2BNR80rfgsDYouvPdv4PJzz6LjydS6zJLePbKxMv1iVp/B7+JIPhipYWPjwm0XPwC7i8
+eeBshJawl0ep0D2IC9HxxZMKUgKsuFsNSNKctnTKWqRc7i4HggnepIGBPbT84FZpylgbnS1nnsc
DEOYlPZnBOGyM8MnwWPxEZu7JqZRWvIJAum0SS17YBH4ZRoecge/pWs/R4pyvUzpSsxh2FRqGYwE
Uhcrg4Am56x+Q8j6d1k6IJj96AaQg8X8WiPq3MXRMBri9GMW3KY1iZG5pquwHS4z0bX2twgpPGvc
VfmOT/gmIeQmYbpVXPwasAUlVGNCBq0j2V11w1hQ568+RjjZo78qxhFnFjsdaAiC8Ubw31Hq/O0T
pvHWdUx81zgzgyslUp2dy1WVNveLleTOuvHA++oWdkHkFCEM0bm22GhJQ+alaU4YbYdsFfI9CxlC
qirGkV1r49FFz4Z0fyuMhl8wuNMFCu2K8W7ifWpdQh8IFQ5lTMv1HGScNeC+lRWNRGjVIlX/Q6X5
2f1ti5v1ivg5lh2niMKCB0EbYdBDl+tPE3p2822H/4/oYTIZo3gDgbAnrzIuKkc/PdllCB7Lji8T
phaWoGSJtSHXo100NMiYb3DuG5IidevACk9MSdae43+AgM2SAT4d22y2ax6Sbkz3dECZfR6WFkaA
sTRCJ84GZ2FmJdq6FXxn3rgWX9dP0bYsqCwT7smIdX+dlSYM7hJmhdRmkJ4wr3gvpvKhNd14oxgJ
EiURG2NY9+272hxkuwp6d24bh97ytzZzB9GyVAK3yubLr4u2i88OtTNZBwF8MMq+iwCuwA7bIxnR
9CT1zwAFHc6Cz0KcNou0fUCJEe8XOPKt8D0Xi0pICOStV5sxd+cd+w1Xr3L1O3jFHu2XXlEWglcQ
tXeY2rYJaO2+JpQabPdhpRJoRvbx4hA41a/4Vt/Dzesfgw1RCNqXpvIrECBaU5uEq8I8M7rP7aKC
0kHOxWtpCiDpjGvsw6euUDpD+VwohlsUXeioWPFgd2lPTIZxDpXwOqjJheVYl1PoftchuChLiZMq
eTf98M8aFBaFE0hhLmxxXe6IPMLLTizVKQflWcYh9fxOvG4Jd4PjAJL1cu6L6Yz0i1GKJBPVjOGe
O645V3WZs0ChL3Yd0FAHY+XqRaS0r+aK4CMbjLjUzc+QqRY9z+6XnyWU7mevFzscXzIubuGZKaRf
SBU4AOuCfKwn70B0cAzVGrqsVcbIVhXpklohO/yCask/dbYK4z7SOXMrBoB+t25gJTskTjUa+ZD7
dSokn8z0jqwoUUmNv9ouOh6H7aMVaKXiy2ix/z8eVbsHA77fWRZql1bd0HRY8Toa7FdtumdB5Omh
Dn4j3rz/luB56VyiTPNWSvG9F2mXmlUoQ6rSgK0ERowI/YN3ZSExSdy2XOmF9NvgJrRZc7gMpIqR
iSMnSbFsz2Nmp7F4TK0lhRhPI82I1XbMDMfqQyVwZuhhgEH/1JCOyCEpjEgWIxT1eef25QdSyo6r
yEkoba/F75y8ArZMX/SLIAkI9/ABbNR06ggTBd796lj8JLrv5XUMDzCT4eR5+CBHefbdOTyxx1Gy
hVuJlLmFydnsilN5biZpXKNwkkGpv7YWIMBPh2mmVmmUJR/FnbYmnb8mcMaWYzCAQHiGet0vxIad
9a9HV4ezo7h8BzrT2JSJ/9eK719NwFC41rJCr3GEfmx1hhMPaWu75+JqVbcelo8jV8jrvIPuYgbt
kfu0siTsMqfDswNxBvc4OwyrevGwkPsTz62cMMbr62iO/coe458VcylKSkUIqDykzK1t6gBYRrgZ
CquaXlBaHokLUPQ/HSKEAxbIzYaEgkv3ey9C5WJf999QuFoeH+MD6YYhjAs58PD+6pq/1MWhKNk3
At1y1j/folhXMKw2GLMoMNFMJLQYmrB17bCUBc8faHz5nc2yd5tRXPCGbT371loJUf4xxmKNs3xZ
xyO/fdCzjLFE0gBrSO9TiSA1qjxAgbBfjzrBJFPrstu8woW8mKdBdbTy+A91UuUshJqZtFnM1Cfb
mqC0YHQdh3iiKlwSwCJfe90PcE8z2jScdmcP9zG+7Dvl9jNdjZn6izYFlr/LGOJ9uZsHrhE0ha7o
s69tRLl3ac+SR0ypit0YDXZ0KODMRDxp/ccTm8n/oWM7Q5thXYyGkwG25odjB1fW3uTcIB67rtmx
AxE1lb8FZy4P0iJAGurcYOEWyxV3R5BcTz7QrjLL5RViGPkdx75EnafC15AVk//VPG+ApLfTxR5A
DdDQTL5s8PhbkzpcaH7nfFPBllIi1HMIhlsTtq8gBELML2KR9RfJ73cMtgwdVDOFDsDrokEHkWQC
QeqLq+J0A53y8I51aAAYlISU/BU7KLl5jhEhAcii35o3D5omRbxQ2WkQ3mnQHDIytpNtlZBXQXl2
LVMzttf8om6oyLeKBiURwsMq1rUOONQ8Cg+oRhvi6w9x2BE2/m4FiMol6Jb2t2Ss8JRwGJ9ir0Mm
hV+Q1ocWz9n8cVQ1PLvb8lai9M52ghTEDEScSmdDYNTxO2Gdo5FN2uoIxdBX2XXFS2oj/LPHHa2G
LnSKIR9IDmceCGYhm976xUE8JjMXww2zUmEJywlWKIeR73dDutfYvcCxOmWrta69uSdy4UemgJZE
QaqCSXvOgcNKnyLwrs9eEYQ7RSzmoJwgt3/2XI70qVxhh6WybHZiDMTmdYvCuznsUq5WebOD+5I6
J3aoENrN+4RBAiQuVyHVd2XVBHSrO4smWyFSQ7nqVMnkbQHBJDmuLouGPqMBayLr617w5lYHgzPZ
KV6qct9wlXajtG6zIg2Puk4/DQgSJZR9DjUJLXvToG/gE62RtRDgd1zTrXLnPp9x4inr/lGP2wLI
w9dTNRrFhdStXWrWHUKYFnzjF7WgC+1g9PDxus4E42eRFY9ovWVog/6gMWrAknvOde+IcSA358di
5rDDKp4EPGgRhnc3LYFoXYQQWgCf2/vA0mLbIsSs3Bhpe9U7PlFJhef07Ks2nHLLb4nfN9EbSpCT
X0v7wwCTeHs04HIzMHiqwcuTsfYl74kze5eAmE2LmAV7cLcGMb/amP6e6luOon3PSZF5cNoQhClT
P/UPN8jojgMEVn9hQl9oRW6AOqjkGib2PDyJ1hJHsITE18/GsfCYtdf+uH4KeinbfV4CsAoOdWEU
d4pJpErzvzgyNzDiQGFivGiaQ8CqrFxyZJ1wqvSOgazGd5CHQPQlcDSoD9x3J0BCCybm+8PDwTFr
8kOf7Z9Y0sIEojlT/B/VxF+8/ecL+Uf4BJw2iRp6OzvgRjtAYZ4P1L83tRF3LPzptsomyc24TsZN
eTcxfdKmGvMSuo3Ozam/0dHdAVfEa3nCEBoCqtJzxCtVDgHCVw7gurQJ54Ll0Gm4HXJuFozXcGwg
f9P6B+yNWZtZgMjKxCL2m+j3ceKjjjuIrHDRuWYyLrhmcsyw+BaJ010MI+eSqM96CMtMKLJRS+dO
9J6G5OKwwIyHWdXFxL9ieyThBbODODcUs83mWx/CtIrqSKIlqOeI4B0bSAZeWPcm0jx2VrOuIDnd
rfsnyu0nLCsMpbaZ3y03E7LsRmRz8px3mHDj7FJ6c3n9VxFs5n6Ffh2QLAg4xt5SoNUnoblvg0yV
BLcBMkM7FP+5n0E3i6jrZxXMK2dTr9L0njGOqWxUlQ1vHOjvPFG/q8sHFlrOTj8RDGmiyzJom61V
o+vS3YOVNOt1dzdsj2KaMaIe+JdlXfMRYryxPTvHmW/Nan4myCYQa+aBz4MhN+sED9lUjVyyr/F+
nuDO254zqN3h57HIe8IaCRWNA8VFk7lOig+mUYMvmax40Uo8OZ8Xe/UEBsEhFad8tPzb6c16+gpx
x0GOVGcNTqX4mhwbmYuTNLF1jySb77tFjXaAuD7rhrMXMB1i1woI6WZXhICZSlYst3VA1cCjwsrP
TABjZayki7zEL/25agOh3PbVD1TwyLnsA3RHjEflan8AOOW2lxS0OGS84gmiv6BQ9yFZrzhmoYZR
RdVF0VH7uRxW7JJTWSG7/G3HZiA/1V/iAn47PBHKQUVnA1gNpa/5ZQ5WCL1f5L0bN8FZDC8FdmCY
V/undbaz81xtixqQUsd5vSrQhPQ/DgiCLw2+6h8w11PNxD2/cpeYsIpnrN4rR3hcUBfY3y853HX1
B67OXFoZ+ODtVoCYikT1WouL4ecJ3ovdvWFQdgAXRIcMQCMv0mRf3RX7ndfqnLyTDViWPd7AlK7M
zNkJQpTK+8/+H/j2dUT+4pye6kq09wG4oks8zJwqHI/XxwbdF80N+Br0iswe6OHoGYy72pemqgK6
cehqbipMcAINGYi7n1UlKnQCn4y1XySDrBgpy3WYElN/1u8/3TVoYFo9kFNc6JLhS+CojYP9RxtL
xpWVsrLea4KuwjcZ1f690B+TJvryQeYKznhx07C7FSojeIn3NFTsIY+VuOeFNT4FQ6ro9kjHTtk2
KEdggrioqangdrIKkiyQG6OF87P7xGZzugCIrSq1wjkRjIheNLtIAxDvc/ravWUIdGquR0CqNTDb
XrHPzolpVnDfaMzrE4ym4/lnKTG2tv5gc0VsaFLFaTR81eXIpSOrvhXTdkbCL/IKr/jFW4bOtHTJ
6UNUNNLIA2iVkebFlgVI8wnglzHwqpXLh/WRx6BK4aG3B3LIn8CGjF7rzLGDckNaPUtFhULUEny3
MYFGfR2z/m5sQ81LQpwT2hCWFljt1LsTKQjeTRmP4NIj0to+BrDO+0B093Q2qH1XyDj2/LcuDEpm
tF8gxrk6AZtgIO3r4flfAd+aVJ/4Ba16aAjAt/KgP1b96/bwAM9GFN3v+VDONW4CViZoFlJOJrQW
gbm187AZu0cOjLvoZMKqyml07xj8tdVhNlfM4zVso7gF5BSSemlOnHjQHPLjnaKGysgPHfXaP19L
yXgjSHdlrPlLmuBUbNi3b/7d24QjO291CzEKVUZ+tMXvP4OYWR5DwInRa0b09p/tDgUIWFKqH2Jh
ek7kONAyLrwiD4hl1hvQulCF5iRFKTNp3fKLoA8edchhV4Dgplk4h9t5YTPTIJGjtmU8+gjlegPI
gcDKbQ1+2UX+31fGvS1AQiOutY8TnYggUnHCfm1RT5iPJGMFUW5i+CX0M1bJrMB1elADWMAFuDPC
/n/COhuT68hYZKuk7Nel7Zj68/Q5ItYHXJH+UyYLZGV2gTanAphzN1p+r2f44R2z7J8QObjJ2rpl
xWMMWzKXlKPX0isLFiERBntASFXY0ALtcKqS54l6qK9+/2mcfLAXfYo8t6YmlWUFAjnluL2TmmAT
oDPalM7UdamSSYlI8NGyxQYAn0oioGcQIdH0765QD68SFQ7A8jlJgABMxtF4PuV/XgS+vhDUOUjz
19So+fe5i/YETN9EEhLUutnzkJbh6C6TsuPW1ejKW07/lRjHO2fTHkrLG12zT9oGJvC8mZmz3Tqc
4MjpAl5i+D264HZ/EALQVdhSBFT/d6cp4/mGUmp7eECBTgQA4ZrwI7t/KgbLxY9mCYKB8Qi9Zwk5
4CXEL2XNI3m6Ddc2bHVFJKGVmaEEbQ3UIrtb0uEZBIH/G4uhxFiTt3oDfi8AeNXtMEsYV3bk/vGY
LXW8kS9JU/o6T2Eux2xuQgFz2d2ZU3S4WkkmQoHUJbTjyH3twnGDeqLXHbNrLRT/nkSu93R0aPUO
PDlV9D7S07atBlW5vlJyYy0N078J2tnFqh4Pw3BI60gzw1QkazruBnlQSPVJrV+WBFXGVEN+oKfa
qs+tPZQF9/FRPFZcvbMgM3fSbNjaKfgkzXfeEy7Kp/GBdr7oDSlSbaPOj3NFFZf7R1iZYnheRWNG
7cQTG6mC+Z5/db1lDz+/GR0YdDQnLd65SeHMtSaCmgnIm56lMQJWe3vRwBvKdhXHG9pAYKFScR5v
HhLG4tJn80tHUtZs+KeWAKkNGJy2x0VDkLdAuMdaGH4SKufzekFY9lj+ciwDFvFap/Jc2zMe2puY
WRmPyKYUsXAtA+MnCFfLv7BgcYrlrsXasegr9KZiMe22fKB1m7WPwB5T/Rtjkq1ABS30NdkW/GZB
Ao4mzAFhK6l5X9gXYsc2ERyiXCI+dNy1Dp5KJ7Mf+9AIrs1nP+bfqsNfzzEJcI9oklnAP5PWVRxj
NknfTbC5EoWg4rV0Zz5piit7mS/3s/JgKnga6BNHkeW3yWCaoIcxuVKHO0cS9ZWnBM46yHMHN+Mt
Wrzv/+KikrGF4m3Bcfsm/FRH30qFST4bLxikjFwDWXMbXt1jmQvQtEUBHzQo4618wI9hwwXOXms0
cj3VmqgIHN8+EiUfzYGGXeoSUnSo1gscFLrTNMr1H9ZRtInU90ASu2poQlU1fm7vja34eJhS1t1V
J8pe5+2DsCbbAN5KrsmMofnbzguy/63NOmQVM3PlBm1Oi1wzQWyUzPp8ouKbnnl7v33HA33Lfveb
l3L8Z4LiXe99kNjwhfqD/HT6PW1C0L+7pSATg23fjEAUvByDcRwAU17s50pogLngiJQmT2N5VY6j
vjwcEUU/mkJvZPzB52HtMEJKp1br/7GAMKYbQgPJRjUGunI+xjtGe2S4Sl6gp8QCyByYoXxqmjF4
vJdAjFlgU0REIrRq4ICVELJbonwj9Hz9yzqOHEYUBF/Jt9xdAr+lvk5gLaRSillSKU5mIyaDbQzI
vEWGOwyoROTuHsnJLu5nKhThDhoVuK+6bomN/A1Xj4+ZBonS3PFD3qf6mAsZ3KIs3T6nmlA0Yxvv
9noVkD0Hz7xLXIfpMETW48usMEQNhCFBWw/OezRlFDS88XDBSuQl6aHaEy2WlGeZt/eueBl0Z2AT
NikQLlkDjaGNN8MzRBDpusQ3DS2N/MRz3rryJpsvJAaspvi5wY93Y+4zXMSIxINI1bsHG8JKimai
ZQsxmQmQGIDWKV2cbr9k2hZrZUIW64QSWJCHm8xoSl/nKt2HOjYMt8X2E+ISpYN2JtoZuqrD/RGP
bn0iDeszb0rjHmKdKlqWN54P04YvXZgu8awKcoRa/k8lu0unAT1lhx+AIqphrL3rnBsVfw9pXms1
r+YQvtvF+Xon419SR2bkXpYsyg7DXMeezz8yaoUx1SMMv4RhV2Dc8el6+iWLF7JM+ryWA7KWux6t
OWIRHgmpHeO+St8pRqGBpBCMZZUB/JKpjsGz7JgJQMJU2U8zCWanfX3nZcy9Mxwvbz3myvp6nyo5
HqsbbIjJTfNSRYgpp7iVnazl8fEs+eNNpujFnlm+w4oT0yXeNrRVffbAWuDO1qUgyFtV18/CyegS
jM8t9NBHeEKgfWJrobehaHA1hnLhbSSQp7qabWfxd9rze/iqf/JY//Gkanq7+ppifaA/p6rfGq5d
XMZ5wPbpMdRnwqO+xK127uGW17SjQzWNuAntk+5mvDqpvloO94TTLfmZLvqbYziF9X5Gto6BPJ0L
pL/0wTmAmwSkBcNjoabRaFKje4TT9ZLCipSlbuKnDaidPBCARdSZvdaI1uC1d04nUbWgeUpBET3/
242Lz3mT78NKD112V7cLeBdLY5QK/QwqtODntojBMYlzFc1lMg1BtylezjZEd6AS0E2kUYeWdHEs
kwBuipZA/sfhUdzs1u3lvsN5I4yk6GIRhB/PBRA3i7P74OgUZ0rT4Jj1qYfx6YVfC8hKBmF1zfI9
UtxKtVn2PiKmRRfVaGrR8gtUVR3dFfMUATDUAoPRmh7oovqSqHLseLSVYn6p8El97KNknVl7jBRW
WHdyE4u5Vs9eA3u3dgCpEzKtndRXnRm04TKLvOigfUT2xrpzIKYayUsLH1NL2H8/G5fZJr6dMjQ0
WdzJsPzY8oYXCqbzPy4zR8lpH12ZcC/uX3gKeWDmTH0JQk5OxqfZFRFt++P14aDUicYH7Riy/QTW
idXkHjaL6L3LpQsbtelfeWtD65S5hsTOz0vUU/BFFLfJJJMaK5ki7OvhKuFWf41ihyss/qi8BUJb
NsMrPms4DTu9AwxRUrmUWAICCq8wKbhqT1py/0uvBe6pkGGIr4CtyYhgDbX125p9z2OEAia+7unf
VM2p4V3bX/hTrIzVCdUijKKshsAKel/D5sfrAMKr0duWVfFuL0XgL/ZI+jReLaWUUBaZAUlhfAuE
apVrucPkeRF/3P4/+wUWo+DRpa/TT6GNHLT762voIEVM7rno9LA/sNiKRAH0gWxisfIFtK/kK/ll
ecwdzrf2MCYbhkG3J98JrhbCBtbPXWlTqzixLukHwhPt4ZnmOEDjSd4xYAvC4UhOw2S5CImq9EnP
g+hKsdbfQlDfAg5Sh/rrxEPKM8lyJveJ7bOp4PxYkt53vLjpEJ3biqeFDz9Ldi2cwOxoXk4YDVwI
H8nowZQ+4BqsZaBQ75VZH14i42jEzlPJrGArAfnGo9BgsphN37YJE+Dp2rA0gvadKGo1n8zMHl81
YS0PPD7IuVpo6ZqfRZsqUM9NF8b0XR9E0c99Yq5l9WWk5+sGBu6iGx3iyF/Q7coAeQLfZZvo5QVR
BO93IYVMyB0RTS7+y6ynQcX4m2SR2JJqPd0xflmS0eiJckvnOTwmvq9uI/IotbdXBNuHZj50Bgsl
MtxHNUQ3ULYsAzvy3AMOsDV+y6+1dhO+XihkLcvRoW/mWTDZHcr4cHhDv1bU+F7H4miV6soo3TSv
sWQAkZ7azqyaftF9UznPRQmr8RQbm1UEsjYT34Hl3V+kcYRttPIiZm36GjjmLAGS44Kmm8hDtk10
vgh1xT46CKEnz4dumi8GJa3m1CcbWhQSaTwfiGDp2EkAefWJsEZl/MDxxa+J3kb0oKIOd3JHmOJv
GtlAbR0bBSwb7drvbd5wbc7mA7nY7nW0IMhJrBMR053xgqn1EpCD6suBjHFsnlTOYzsvtKyLBfeR
t5R98/rvAosMyiQ7ajAvbPNnTsx5EdaQ9bpiedCj1JYjy5Iny+o2zt37usv1LrLZmjTtt01TUwnt
zx0AgeZo48v/FC0/6nnX6U/h149LPJxZiL/3puKQ0S1SicWTl6A6HQUVab80o6Adl/tLgJsSCmFM
TSBud79PFdQ//Yip+6bEq1sjN/jvzrDqEU1vm5knBeF0sRnbQ87BlPYG8CE+za2zkNRJHJtN2eHh
ySDu+K+MsauiausjrIggjgSQnhlhl+A20MnmGClUfNYbdK5sU2se0AliJ+9CdObNTXQa5CV+I2n5
caFZOfBunK12JZorkmL4vSH3Y6718+QeeFL9F1cQrOTRCwc51qfkFfLedPywqPL5NaKGKpH/JYO5
oTfdBvlwxg1f+hNyIU0yHbPV90IhbgpT6kfcuRSOArlXC8cpe/fnSqMI3nDEfF0H+GawJ5sv04U/
Nz1qU6akrlITm3YU9ijNiVXiyn7YKW/BSrpE2WBCvM8XkrnzZlOe+3sQjkzuRRF2hW8K5DAQ8Mq6
4K08fNTc9r8+DvpBF5QgPffuNy9s9VbEO75XMBigL1+zt6oUm4KiGhK3uVSYTAvr227bYLLijHgC
LSkflxh6OvMiFezrrURMv5qWmA6qiF5lDslRaPVc4pDfYdDMMxxIhFdKwGcWAeIPtfdrB4ZXsS7g
gNoaYQDDEimV08HSQQEE8Cq++JK30UoMbxr6Iwe0PdNhZvLfp1m8wP5MWS9bP/FYWwjPcFzYNMF0
PA3V4zO1sWST+7hvRFzYnL9Oul5IFy/68+GyCrzMzPRae81mqadR+VgbNfkEh5luJTn32LXCAmZ2
Wkgr9ZD5evegTAqbWX2dCDIr20GA9h3V2jTmMJudsUACMkXyCvj8EUBaPi9RrVsb32r7pO+4akIS
dwa9ecAgb0nhRw2UOMMb+0bRbfLtsW5R5y39qmxmeC/Dj31ojgEt4jyyjOgFvG6MVTmkAa85rmwB
IY0x2NubOpypwWlQwLuv67GXYIM4bT8JWozikBxDzuenhkyFPEVHP5v6Pgu6dwdNm6OJJTAbRHb/
QdwZ7iO1r6UmOZEafvSATSWfaVflFk/uRajex031c/ydMLId+sCXS0u2vdKLVnUbLBDocaFd/ZTG
5JkQ2dO2v2EgpRXeeCNYP5jlPtqHl2KX/e7Z/CQySDwG1nRIDeRJELww7KMVYPMRbkFBlb5/HP69
1bn1LnZXVdP58qHTJUGa2m5SUXbes7u6UFfVrRFNotZrpbxD2MAaUBZs0DOMFcMnpb+H9T2IR201
dlJrrzErQf34tpb6YxZcYKleGSLsoRtO2oiNMe0h9KFFOR+ELvy6wY1qhgBwNA5z3x8w0WNIYfAZ
3nLyJ1DqWkqhBgp3QebSRImNTlU4IFqJS9qJXNNY1NdOZk/sfcEwjkUUKHki0ZPH0LEaUGCg1uJr
wLM8ei9ilXCUP4oVKB0FDq+AMM7XYrzXeQnVGYsIrBCkF3phL8TOLTglFVtOm1lt0NPnb7533OQK
kmsu6XV9g8rcxLYEpYCYF9E76drpbLlYbaEa6VVQKCPEtprL+Y/QadfqPwrBZW5UeX8y1uJ5icY7
I9kELejnKJGk1hd2rO9iHH7tp08CXnhUpJgMjc8tyvVN733Zn6ZSHs0XUXjXBy9gA44hUQcJRF5z
tmOAXURK/vTjxsQOPVuxCQg2ExoF+UrZH8JZgFs3RCXUMmDyfET+vAaMekxnAHIGtbj8VT257dd+
o+a1a2ptYmEmpV/SPZmy01mMlTNWdQ2kAsHgrBeSzCpdTvAeej9y9fLSlQjTIDtkfe0lT3+F9tC2
DZviJ3r5QQVzAZiosHvWsR8jlrJKV753kyZdO3s+5OQP73LapZj9kKeEwoms/361j6fSfA55W9ce
q5IBz5maysmYIFhaIp0tlkD0YW8swI9hG5bnLLbjEQ+c3FZZhH7jZi7dDjAtaDwQ3H4/vU3jlVAn
JKpI54o2R2nzAAkM+AfaXfTY59VOK22h9C5W/ruGnbrcUVtp7RhYLak2vrOZMhETj797SvUtboEI
884kNsVfmMG9vszgpzVL2tHJ168JABmza8nxL7WB7ZPqVLQV0SZfVH9wxfvCO6h8M/PYZ0N4QbC1
4ImWhzw37FWnAoDg2APLXKnzgZdVa5bg4ZGeUbaCGfXbFEkBD5lGyTPVsr+Em6eAe8lOXV3Bwj4x
q56cLjGwW/2P4bh3+aWen9sBtYF2SxUBVGZVUDlrOQsplR9fpdzOGrs9a+kf7xK9TrT941P1r6EE
dJU9RFVU4w6s3avwaznw98ySRUW5tcwWnbth4aEcQ946GS7CFI+Rw0f77WHrabN62MjvGHrK2SUk
EENdMNU/KtL9z5dKU/FKfsMK6AWxnidvg0vvcgx2P8GuDbricE7Od3s+ag5LElKH6mmD+6/HxgvP
ejDYXqaCGc89i82JnOLQrAb3d9RRfuJiFP4rWwDKaaz/OosJPZEpdcGaprcRBFLun1ABMxU+WyM4
kbvP3x7cqyqp/syj00GFxAk/ZNl/E8a6GzeWzt46Tz7ppU9ySDyIq3xgyTca+U8pq+ZlUjj+HZAo
9Z/ljo+xHqGQui2KrTw41j0XyZRCL6VJ0QaDEJAnDnFqZ9FwtPIbmEtaTvFHpVfoCkEaupTNrzI7
xKgT9P34y6R/75KpToehGiayiTq4p1pxAgK76LG+oQ5+zCBpmPQZYo5mNJfPjrE8xSOlDuw1Z6RB
7StGanmRj8IJpMLHCTqv0YbEj8OT8MbTZydr57cuiKYArASGAtBSpvEViGI9Vj72DLXbRSm3hCj7
QatN+TNOmYWr1tWR7yXr6ugAU9tcaR2y44AWlmHukoYw94O36/hReyzYZKyKr6A6bYKy0oLxi3EI
OkWSsuFZpzugchU+3NLoykajgtMwcztdCv1hNTmUCHrUunsDa1qb0o+yr8zCNlTb0TilZR44cYWw
vNkZvhWh/yONoA5dWL3nPd60DBjpJUeZBZCfMHLXLR86B6xGgsRpmwP1V6sn3qXvwbD+0NtU+AR2
+FYJAcsURu9xD7giB8exYQSkqIwzjbCYpJfvy7jkL2bygU64d5XxIJI6lpS+3UimbY/IpvzxhgoA
4XcBmbwv4mLHx6/SQVZOo/BiE3w6mCyW3vYPuespRCGBXL15j5pGIcJFdOIqgplhd4uBCww7h6/h
tMocxhnfN9Fir3X2ZPJ+HpSeQAx7l7Su98OrE97SSW2LQbCL5xyM2wsNIxVTCGZzb1naiuJtDCNy
9p1iXK0TXp+XVBj7/I2FFM5SgE/tyMhJ6ewJFAmFN556Ke0uT19+BiwvtAKUwh88jRscH3sm/9ZX
vYvo1Ka/Wy79ghgzJyEv2LDNDy9dSQ8yp9tMhMV8bCAU8mhlX3okibbLuiee5AXBNuCdhfgQBvP6
V3umOJnEZF54x4uG5dC542HIkCBdRkgGGC81s2P6UCuyhfE1q4KUI7Eo8e9S2AMNOuEJriJ6tdEs
Ggu2fJikOf5MDH1VVZANr9NI7mbRc88zL/5kX1xeueAGkrf+apLXcbWLtY2oeP8ocF3wpZwsvvTc
bRRqoX+aB0TLWXtjHtUj0LvNw1U9A0taNECYrb5fX7AsPevk+zve9yX0XwIL9JzdUdGQ4iOSm0CI
Aly7Axof6GLiqT//eca1UvJ/M4KG0WgB4dsUAz3QovT9Osn799rWKpw1UFg2gHTL+VwNXspbBdrS
J58dyGbYF4oiuMf+8MeA0XT1F0KQXZvc8fAfaDkYDdJuPcrbvA9uqoRGus2LHCyfLi2VFDY6f5L9
PGPh7QFTkEIWyH2Dqq4aio1/5Jx8zMKaPPQIq2Yg0BmceJ1PHLesCPUwZSCGoIicpC8ldKhCBekv
vNeYhEVGRtEL8hVkO5oTddoAbPhFOyCqWdzlRzceOEQIFGuCpuDBRsdAcqCC3/1+l4AH342B5aKE
8/g5vWP+f8nhWrvdLO7uTUI5XBUm1JLxWfKdytsJ3zN3V21agi70tWwlZU7CxbhhGMDVaB21AZpb
3VmHKQoBGCeR1RItWoiLFgDyxEI/2t5omX5qVGaTh4sp1Glyef1zhYhxvzfaOLgCZS2GqoEbxjVX
yBhLLXGnrny2/Wvj/vVP6mugPFaJ64JY8TjjrjPaDXC7cZZ2J0YA4Wv7/eCLYvx7+ALE2ybQKD6Q
+FI61ajMH6QdheWCw09k8skll3As0QTYVwBzF96EIJQ4YJ6p4MrJZJFJrIcqFKyoShH3xr/PDA+L
d40NBMKuXl/AqTP0kxeSFaUwjAY7vv1Go23vJnIvQcdFIZVpcM7+CS2SDWF0zqdfx4L3Ow2m1VDc
K6VXhLwO2wNryf4Fkv0ifF3x7HSpqCUw7FUAspVVOIqpiCK26vN+Pm02k2Ktg+4dDbGv3IeulXYx
WqgVcrYRp/z/LPKoCBVLkkQhupOcio+HiJ5HqcF+EEhg8w1WOK+E5Z8WLOHVAzb6CoeflNCzZx8L
gq94RizLzceBaY9LmnM8roAmbdzw2l53qAiWGWKUwVAceDIOELml4Sil44fO29erqBNufTeZenBG
60g6OR027n5rwIpKl4awryy/maS78w6wZuZRJ8TXFept1NepFuigtB/AUtlZXn+3Mcscyso3slyC
K09Y0jtLLzqVuHt/0WmlOLVIy4Z74XiQwATxor7jGFR3OcnrpfLZMPR8LzZxavS1PmP/eYNvOvbO
0xmteqEVZKhyi3DHmF/ZMGLfE6zzdCfhRksvky7m5uPNFVoWjgfCtFIiXOkE5/zQZ4J9Bkv7VpEP
EsKEb18FCv3+ola64Nv1SFqC1KN0BTSGQx6XAGCrs6XPzhIys5MzMQB/qyUTHwvsLijcVeo4V0/T
Dnow3PMvCuQMHWYrAuM2xU1Xm8QAVHPLDDrQkERySreIJ4XxnI961gqwXsZivZ/V+tDBmHYiokjQ
JTh9/8FDhLMynX7JaJYSfVxyuTouZ2DhbRsy6xMOHYGz8kvlRo5AqwhyZ3P/EbLyQ8+e3qbkUesb
9nbBk2BMESqjl/eGXviGM8ckzzJY7iZC+L3BB5MyVzmmWU3UNWL8iIa9sk3fLD0jzNuybIb5reov
dhtUv6FyrDnQgQHS5hYmkxELfsrCo1U9NaXItf5GNyt1niS6oLsbgIlh9DwxwEHARLajU7d2/F2K
FFk2EAmccNykOA3pkvF2nK+fChVg2EoKB33tJQAhPPropRUmuVc8Vmm2DYKt3UkTS9hlsa2R16u6
xA7t9AzPyk6dA8S9i1RRer0fLXLPcDlLypX3ml55u9VdPkGsS60JmeCCKgrEJde/UoG80aEAosYj
HH3LVNiqTJ+uW/Sl19NkcZIjn3cLKGfTLjQU8L+qMRSZHn1ecpaoLjXNBtUxV6dYVGcy/VeuYECe
01TM5e/kBspb+XCSZILWp/IaNqoh+PNuiLGKGB0hlL5n0U58qv5WNN19Gu2tbz7bmT7YJsGYEKVB
Cif+nCgK2XhAfCciy06xuKXyEZUQrBrZc0O33lsLEgFsKRxdvghIrK0fKYw0hdJuBrhGb3VJDIXr
ydpgx3nwzMufUPoVuQG48tgf9Xz5wsm2DJlvYChPnxJ+/5G1Bvm+/GUgRnnKggDa9aZS6SqXGRFK
1tlcyP9lXhPSLKDq1Tx1bfEJo7vMfFTPuOJz8+pBu+6Ozvna84hYFMpBnU4N6dWiRmBAPLTeiG+P
G1thxpts6Q+/xDpFIEflTbB3Ty6aCIGpTDmXheeUt72znPThycs2bZWhOodGxMROZXnXpO6Qk5rV
qpoXzn7BjL4YyKGlIadTdWYaWiLxmgLuWMIsDrGrdHBMy+F6L/ejAX13+1TMM9djJS/Ys6u37ffa
2REE9VWDplopHjoquMRzb29ISGyc7k6AouWOeq7MhCu/Re1DZwPEIPGaBHFaEgPvxliVelQvXEME
7kQGZR2TJ0Nzx9lUY1bTcE763aA9t5rirCzcvm3d5Fwufzmeuddlv3TVPpvI7gQS9KKlJvNqb6Tf
f7ah1b4oaMcpq8jcjnOc7v4mWbcjkA4Ye+QD2ZlG5gyxyCAqZ75VEoPZDw2MxBPbL/j2+8MJHOOX
ic4+d9mcePzhwSe/35E0E/T4iIYQ74Q8LlV5/Vq4otXK1Wq2cyqpHS+k2+cbE97zaLton60BO1fw
nFdoGhDhgroAqYKEU2L6uGCspI8AKkLcioMyLB3xAOLqzg3tsKjq/5XtgpSX4xhVWzwAUUeHwwUk
Rao0s8egKrjLPdikHhIfto3MMLt60GLoMyoDedC90dE1GdlpIZpXbOg+mZjHE3Us0/fYrAPA08pX
P1YGk3IK9BZ8Endam1MuY4A/ARiMf+BBTr7Ik30kW3alnRvIT1kyrZuwoaVultt4M/q/67S9vGls
BBMKKkTVX9C6BZ2sIDjL5teh8p/TIY0pY3Co6VE6011xV4jpvw8sFGc2rlPIMFOhHOs+GJDomPxX
3zGL/hiPV8Z8/uwENV5flah1deLgSfuKrR1/5KTTl/CUkUFpVt47DGqgEE7hiVIURBbVZJK9+Sr9
O8zlU+6YRvySfcDAHtqk5Wplt2POIqnFXjfcTI7zr0CX/GWfZwTeiN7wKBjTNfqXWakG88I3TnCq
VnfridQVLc3bQrH2mRLLuSUW0MUnhCyZZFA4y5FIhPUhFHB5hqMZwuTkMrqcR/NVEQKF86RXGsFv
dzD+dJnzF/9n66TPL14rZ7/9mUGQ7a71Gz7bJtXvMkB9XOEWJAjm3N563mBk4iY/xaxjgPPIDMsZ
U+VzRvAO3H8ZhgadDFL6Ca10HYr6dwVpXypXfgkg4pgQVutedpQI6IWEBXChHIhtDQP0L3V3eXfn
CHdsPxKphcPHa23YR1WDqU09o+Xkdq3yzGzK8vD3FEpX06b5uf+2qb7oOSpwK8XdOUs4tbm0PxSO
1GhguhColMfatRV8Z2XSwPH1jBY0j+fR3pceAlcTryajlBiuNdvy3uyzSefPuUfPVeId/cgbdw2h
LbxAqEjNeODwla5YZr7OljcHPNH86dQdqIP3xzvVnowyM6VueiYAe2Z+AVjdhvybPdJhOyY7QJSR
jm/NpGVhN9GnQtA1EjU3N7VyjX8vT8nCP3M8nKmmysrOhkdZ1xKeFNwQOpxFNiu52PmwHvKBfaos
HcXXumSpUCXrwxgXZBw7FndbF9CIAOEoPg5kVJ/iVSYJ98/duUMPf61KvTAjhOxylTCvcWUwMnFS
4Yrjje2ci3gRdibc0srZHs5Nssvsmb26XHF/aROKanjA81FhvuCsEnVdmHlmg0gag/Nhe/MYYmKC
7mSnvwtkHA+YnYNNHdy2qqfV3ux1aHg+Ax4HCcoQJtJZ+d7S0eiVOIiLZRbipC9yRovh3DDBH2JO
zby7uwVYZhNeqZbBOX4AdSHxp7kF8fwz37s3RJrlzNsHviDOihbRE86ISA7+vbcu/mGmU5U6Qcp7
4iNuf1pKYZdawyThFY2hycB5PwjJxJIc+L49xABRTKW1TLnlbvdFRVmtTUWUbed9ZIKB6P8vWuvs
/7HvIjD2pr0ciB6tBbIcM4xqgffnKYVf1f0r1FUEUKYeBRPQVw/4qivOJnnX7KnVdgPpvIfxqrWM
FqbOSV+V4QSeRHvxPrEsuMgszv/gpjUlKyv8pWPBL85wjhF23kVL1aVoQqwS4Jls8bQPi76SlXAN
e4qXp0fefgtjYLk1zFTxjZQVCsNyct/CgUKCRvWvmhsIGN874N2MWuetDEnOjavWoamj1kBrAbzg
PiRHxF95Se8Ly0GDyYyRVXoz5IilPE7SfosxJYRykugkjkdMEcj+1hu/Wyu/zxHE4HpqbcMTky1k
mZyBR1t4dVPr5DV/3U/4t5TtjIqjK2kUUo+1ou5znHGwtk95dcFhTX0CJEpm6kNCCGABbJl1n2ud
Kgou/ZfEJ4uvOwGe+EJeJKNGt2dqK6O8np1ACW5nLMMe9xhMixRAQa0k/8syRQP8er5iayzAMaAX
YHJMhmfjdiTZgq/gVmlXvJKZG0r26q3Du7aRJ68b5aADwZcsn+n66GPprjFnOUpunAzvviJwYHLA
N7o1amri1CRkmfFHxW90Z8p3NXpOgF+Nv2UOWh9Xdl5eZPZ1giNVVL49tskwtybEtzKLt5yQNhsk
tmKrP1Q/CAi6VPnnJvDVbaiy2My4xf2qDvgFlWIEef+CJWvymyo78XVVuFp0rXO20tGcHmtTmKhw
tD3VSlaV71nlymHQEEDXB0LLW3dw/E9A2t3Ks8n4zEa2s5Gdwg/jKHx/MJFf6BSyUClVxo2FANih
ZHOKwvEzbHmnJyCNzNaG981n4HOgHGyklgZ3J1SL4daGcLJ9wkRVWiQGE8P5f+dOGm108AqbPcBN
DdtIOY3IMYIz8ZWqtmOGK3gqX9m66URVzFbfemoG/UjK6hCkUmTAEtdT8gOa2/SBbbg9EsWh0/P3
SEzP/qfIyrjEbJJeuWrBhTtYJZ7BOGPOq7iWbxmrsPFySmnvAroX3Jl2W5CAJshpUYv3AWGP4BhL
DtvgfTtTqGUW05rpzlw/dXjWMPw+Q8R1qf4fHqYGTluO6MwT0rNo7geqtquPaFBo3rALggYWapVI
M0QglxfJ3haLRloKc2Bz69qy/PJ/UugFTM6K7h/LDdyuqCL/v+DKcWsH2Xzhs9+5de8fbIUGVWKe
F1XfcVzRNtEZF4AvCOgrqvW3l1+vHUj4ORzl4V9j+QGbVWur3SxoklYl1tikMtp439AuxG9hBbpY
kJqS8pd5J2AD/2UApJzti4GrxflFL2p0Z52jMwR5sCV6RMFeSXTxcxA5gPnFMoYbhba80FVR7hbT
DGpCcZ6Jh9HBo37rBwrKEozAAPWDuf3Lb0UEU+GjNUxUVw+9u5jnABknY/W27ZTs1Qiy8wH5mPXc
kr+OEhbJ5A41l29IXr0xlh6bV1G42w52RNcubrGnKrKWYh20f/QVC43LOLhUuevZXY64ZSk6Dag8
V0ALT0n1Xiviu2PWzHI06QKRPTz+42vQ284jb4UT33ztxD+CMSR4RN4aIXzv9tNTvt5cIWDWTeVk
bw7XMuChff2EM4gvoZxo5tevArijfdEyrIhQeFqIHNATHSCc24WI3Kr7dT1T284d6sbaW0Ae9nGE
VYQ43US2EZAZLFQQEC3dUZWdbEsqgq0FzzMlN2gAjVOHVlJ5r/z3iNVZ1zUB/glHNw+3DNRHhw9Q
XWi4f39oDyA5Oiw3kXc5uBwGmdeM78qdptQ7UOuhCjLy4rDH3Ch1PBZ4izEaVLCzdluDoNwYae2D
6hAgWmYy0xYeFOFMaOu6PLExDJ1Zd4OcEt2cTeOvbRcllpGBnFht8pE5pU697TV0Ta51CWuFScQ1
ydp1ZA9tVRbKI4btZgszQUUzSQDiNQEaCGWAqSIs4XJbda+lCU4GGRWjvAk7UfRkloWPiQ4MqD/4
JkfnkOHovg502NzufCy3CrxtR8nOr9Hpumv4ndQ/tajAxVtY2xEtt6AMY+xARV5WgBGDa7zxKbFf
zZXZFYLkHOEn/Ka0pP7XDoIllk2LcJsUy2aNepDbLWPgCqMsNJW1TophJ4IeoioglDcnhjN5TvyK
stzUHFaeJxb9AAf20/SVeKDgL4fP2jWPwqn5itWjWWKXuXWxW35kYzVgZe905dYrmGaiNJ+ltZEk
+nExt68Lcbap7HGnjMOufPjMiH79YDp1sJYM/r89RAxOjOpx6++5Ar7LJbIa+HhHs6f698XZ+owG
BoxE/8eT5ZipKoE6i+oiU3mRSrDsQuz531dZAAJaHnptFS2Z3LRwDnPmw/dwzfKofAEcZ/9jI+D8
Q2CPlaojqK5whMEi3AIaz0baASbIAuzoibS1gtXYufDe4tS9mJYEvNFN4uwDKP51+BBkTgoUgwmI
OP3xFBAmKtmBNz96kGJO+7M25Cvo/mnK3MoLQTyBEoq1pJKU9loV4bGjMFDI6UR9BP26Har7NMmw
yNlmLRaB5ptkMRSiDCG5qT4T0IbKUG7zPV4jmrpPyIB3ax+CG8y95gFNPZ9FVuQ2ok3ApsTCIMvl
5DcKic044kCflAzzEC1hS1Y4PLij1bgVIHZIwXtfOsU3jXdYDi5Sk+bH8FEic1REyBY+ktxFw0eF
eZlc7hMPpZSvyf09u1y51a3iKjomqqjdCcO84zY6YHdDZ02shN+QYJxPYVwVZyIkOhiBScaqcsQv
fU9/cE3ewZRXKrqZLpYXSAVsDVhPEfPt9Gtq8D3M1AI4hCVh3o+GGcITEYFXlHjs9/CrggzbLy0l
bj+rPA05bSWrnX4IeiU13qG1qNX+AW9vdUHKr6piO5qqTaH0c1z9FzAOq9Zx93UOAKXbH8WpjC/l
3Dob5fu2jCzvnh8U27pStMufnw/C1TtulJBxr8fzdPXwoHkN8CsveSvB9xRxOjDRlNidCSvx6lUI
Vup+tGwZGiqel1eC84N5OqUdj4ZBaZ1YEpcjJaWyMRxZ8BcJ2Y0sBZgl9R6lOPQdvY6Ae+M0Gn1k
6bdHKttlNf5dHbYluxbqJq7YU1y2WvQ1f6CJK4+ImbnzaY5GiRvFvTOKMxnJOpHh8+0dL+QaG4Md
n5lcVC7uXuoRsHrp4rtpHIqcoq/+pjsqCvGODtSu0KcIcBGXvgKR7fx8CR0YfjF99Clu9arDKS33
l9gcqtV9msSQQ4FCMdSIKrsn/Uws/MwMnVXwov3rYvrxzrFUNRmlU3es/eMZ9ix/t2gEe8aMZVQr
nLl3jS2iT+NIo1ritRr6Aenl15Vtp32V+AeeJo3+/9nrdfrde2eiBtH4J0Q/BzkWs8xETBlFqxI0
/mrGr9efG/xyTmTIEcGgszwU7ZkqMyt6Jpw4Km64OHybDOp/tLCOJ3QdTMMByeTavc6TAmxlvrLM
uwAHRaLcBvs8N//drkezGvU17bbVFCTvq4MlhxZV/xnOBOtUH9Sm3aZYYPPUQB0doFqUDdiLxoQT
4KJNn5EyIVN4h9vUR5mC/W9sPgwv76GB1c6gGOd3UgMP3LhLLNjOJhmSMfIymwY8GXEHKO6I9dGE
PX34YscTMhPJVR5+yr0tF4kYI4SzGSEToLfhyAUGjn8y+FqIZRon0w05/GW9YliXAbd1GqnMgwb2
vm9BO9zVYoM97wewrfqWnkOtSdI8tYwgChbiatibArpTyfooSF20U6hv13rin90S4iD568IV/XMu
A6Y/dWpKuhHEARbQWm9xunqFBa0OjfoR62tuzn3bpJa5kXR7c8n6WVocoB/GiVev20ccjs4Pj4kF
atUN48TPVRN7H4WBcwkoRHy/lxmP+dgKOXwg3apT1Z++OKB7udnFvmy0kE1b+s6jmxePvkdQ+9ly
HTC6H7ZCx1Bwv0WUDo6OV01R1BMcc6ixiz7jL9yv0KKaVaBn5d6Rz4FFbVDUZqse+TFbNOG+82C9
qYUqPt0ldNeVv7JJKAfoOiOB9cg0WQqVM5pNCVaBnPy0tlM4KFApfyts63ov3rihVTq3Q2yjQoDx
SlNl/2sk3pbzj51pCJ5RqEjRQ8R/mL8l1E2TCfnkAU3TVY/0IYrKIi/nO7QS00stWQkP0D6K4rw8
JEEk2S71+baD5QdDe6Mkv9XQXw2MXweDjjcLA3jhHgjhfSECDn+PxqiXDlC3hw36JjnJAc0SPmz2
qomzslmE/2Pg3gWeIkRGCWiMT00Txc/VfjuPOxhjvUuBwCfDfHS3d4LvEnFnxdsBEVlBQb4pHMRi
19u9SgrHZtiN5Kpqf+l32RVO6H9ImIX22Va4nt9Xd5AIY0/+AndCEmZqULxvGh7evL/7vA+Lp2Cd
ed6l2OEcP/dznnuHkp2ulrZDpi7/MYHncnMgdSD6Uuts+/tlWVw3qwx2Sa7nj6Fs1AA2l/Mo18KU
/MgEsSNYyRZAJ+3+w3Sns9BlBaxKUiWniNCYgjab/MtSBTH5l5Z/Yt4fO8mHoQMNn9Tldpj3Clvr
U66EFA9aaB1jlbAUtjWYJyEIRIwbTlQQw/oLMJ4Nkx25G7Wh4o1jc7noStjo0XjUZgrdnfUYN2G9
hIRZAGd4xHIaDoT+2+LJKa315w6ZQAfboI8qI8Ik8OveVQiwnoE0XTdPlBaPoGQnzHT7YDr2FKrr
PZe9MiXGAwvd79f68zVzu6fDYCtfCAV4hC88NQcrtLIpJP5hNP/6OgsTJzMntdzBER1PIwLuaNku
A9qndnr1d6IgwMgDRtyCi/8Jp2MMgYNk69y2F5O2eF2KTyckk9Dd8KiwebYQOrrTR33YfnKvD86x
Wll0rt5vwcxV1q1z7M1Z6WDPMw6xI+Fi/j6e0tg6Oe8zguCwE117xjLUsuPtlbsQEIKyUZRy8Z7o
bu0W+LLXlChuinhGGx9eaKcevohZe/cyg5q1stPkzs+vMMvpIufXfidsB/yQOwZP8gE5FhkUbyU+
JvcG49/BdVuERevp/6P5AWqU0lyYxJYEXRg148YR9QQbVSDfnElXrb6OYJufIj9h0hx7Gzs+m8rW
3INrU7vGj4YTwvgVeDzbdIzyk7IdRC6YgYV0imb4QCSBlJ22ulk7CSA2qZ8fz7QmVaQIIS/fYjZV
8b0ezsESFV98kqRBFfVQ92vQInICpiq3E9QSEpbT+BdH93HaG4JOADPL7UP0Migzr6SsB+2IHrfv
uqQQpDoK6U92YQAni+pngO1do8AI2SMnsN2lKd3Tqh3Tnij4LjRPR5QR1R41xlR1mPsouzb5pdfn
UkmAEr84370UpaR1KFEOaCpKv8ihJq3psNfHH4Rmtpdi638/Nw4dczG4if/4zA9v7LtDVD//4T4G
CEOxxGzApb5DgjZTxVZkHBHt9BTd1SOEMsjqdx41Q47bB7UZhoJmGxiruW1V3/BSktz/oUYfjUXx
Vny4E9r0zKoswaLaQ8GwmgY8UgRhberot6g3rBxl1ELXW1njxnc8ju71xXnWRu2TjuWwDYYPF+9H
QeAfZVHVmPMlgySWyO/n7CDCKJ0bevPaTXrZ/ZG7i+EOSse2QDEkeY/LhiwlH4QtB3VMk/IYsGc1
ChKHazC0J8t9QSDEmjsQGmL5BASNsJVqgb94EUytl2rX8iV+BkjlbEOKJDnLCfPKJzm7FV6LLTry
t73+UhAeO55Km/TK2x+7snudG/2/LmmnUHUaZbhV5g0sgt/9rbGzAFaf6zDQ62pos3frNBRpTb14
xkUiXRshYBfbRoBLPadqCtbGHzJp93D5ASmDImW7K1OTKg8UBxiJ7t2OuJz8Agmx0u2o6KBcp2I6
P3eFZ1bKaqUFSZayE3MOampJBZzbsMzuhsJk9UonFtNQAKQs4IMiMyfcSFlWZ7nNa8JRMa7J5QRG
HliAH+4vgBGtFsDDU0UXR3MZ2nEB+UL+xuPvxwxxNolAl69MoCPx4oziHQnBgiitm002Cg16C8vK
jX/xx1MEVywFiN+ydMjxyZVRca73A3FpeFNt3DWSGmiUCKsThvh6nWIMK5Jh1NnVIZ4DjxgE2Xyc
9sZKRgeVfmYb/x5Gbd6jKtP8rfLS5np/P1ZJ37wO3HZR16kXXj6AVA23CX9kIX0prR4gYKuf+ZFD
3LCsD0dX4SQ49Oy2wXIzJbnQlCpCRSY1qiroT7gcmWSlES+oSVhJ8qUoDDa//PzM3V/kcthz/gZu
2paDeqkj0FtG7+r/FO2Vbythg2saz2LOQJFL9XLl8HrzRhjzgM2c05UchWPOZJ41He7eQoNxFSgy
HdLjJee7CdWxwNXGGOILOTXwB1uSHZI0D/4mVTRPfS0YkW77NB+ScNsVKVlY+KasHHROASFXropR
GtAKMhk0nNT9/AEraJ9yqcYA26iBJDlrraOFVCYThGdOWf4HyIWhY7NAhdslODlymBd5SVg/4rEb
R1RIPRFv3HYMplDinAK4hcBWSCiwMaPs9s9qrkejXaypd47DDwur1Qvk+R1+DaL4ZxAfaeTOZMBE
2m2yEOBrc2D6eQJ3tQ5Z+/AXcnCevyq0r7d89Uhs9gF7dwddrDgQ+ma7VMbOpPNNWMTb0hQ4QCnb
miU8Y554Ma6fV0mrv2ClhkI4T7LjmMZ4LJlimsvUxmw0A4zlteVGBOtc34UVeiMRKdgfubsEnPLc
36vV++67L/w3BDoUXYx6XYwFlRsj5KXZjMjT+LH1dh1T81VtJRUWre+YsA7UCv5oyt3IB1rwlI2U
DSHd5xYKn30NvPp9/s9L6kvLbHUIfIlAdDMtb3W//suNnA1DMTsKOBUqTfC58kv30dfCmCgAEgf9
fqQeDlx9KWMdv7o0pdNj4yWNLUCCPKunL4if+ljfrCENYCQsGEGvm3zqTQ8x3bG1Ftu/XwdmX4dd
HZ4jONwGI4FqCU5dHdmRflCyDH8NXjy5aQSheHcuqtH9Wnbhr2P6FMnhNGD7KZ2v0x4GOA3iu9IX
hYOzg3vGfKd/2OKb7ajsTMU7O7LEWnjcASH43qKeWrap+NydKe5//5jBjn2M1xz41x0P6cfgSq3f
PYitpBESg+Qdlsa0SMGyFukRHtD+7l0e163xw60vcpoSheOsBgPS4kn4RBKbc+wEk3gpmphIkc9h
DOVGw3/g5teQekPdwV9XxzX1pG68ItNRfxym6wqg+7mby8f1fevaacMTbvkwvuBvZ4kFRzdO7VqG
+4/qALZvA04zkaFx+VT+Nj/6VNePXn73iHjeMOOSr1aUwMzWlZ4QwhbxxGoMWG9n7t6XoOHf4gsV
LLq3ACfo2D8fP3AmIv0Yu4BxpGo6lYphctQ1wDs/71MizJYv9JkXILeC5T8BUfhAVbGsRgVCwwHO
3v3ZxI5TkmA10LPNfTwcyL+c7QSrvCsUTj1KAH+LGAgORCuuNoTsDrutKEOi09jm2+jm9fjtKBCN
JWMHK1BDEBbkT84n+bYvPryLKwBFQm+LJTqlz22zL2r/8HOHF8KsiZyYeAvmH2MTyNOXr3gB2Cjl
4QL2rQUQe+PdebmEQT4h0Fg2Y+eeKxAp6lfvdOd5oaBZ4DHQWR4BWPSg75RqizTaKQszBhkD4f1g
YmzIBBfdocipeGPVNEiBYlG7maC4/Rg1xtvgZEJ2Tst4pGmkYYeHc5XsepKf5R6kfexXQVp8L2uY
sF3gVOU5p281WBr+mrERD+DQYtz6mlklDtUKJA64/hV3MCYG6LeaE76HVERYf5g48MqXUAsSaPJD
ZtmKSjst1yRiskHKRTu6OUihbktW1m4WSG40raz+RqUe817ldanVNqg9JLbXkFEr6h8LOZeAo2/g
nQw6m0Iohds0oue7icc1wRGEKti9FZ0mU/u4TTmwB1wuEp+bS1nS1OFI+DuW42TE7YzM/1FthRNR
Oe6CNcMHwJq0yQLejzfh72XOgGA+h9oURR6fBQDJdmkhwsGSM17goCy/dUkSJ5h/UPuWyU4Xryrj
l7EBfHtiGPB1EEwHMVDlb34/0vgC/nd49TnwspKmGqU4NoaqcWnghvaHN21qF+dn21vmMH/r+FWm
Nwu+lUjs4MCRtvmwWiGpcwD6v4PtOvb8nBA94strtDiE0Rh7HcJLj9TP5cPHuGOOaTbMwOQcJKCd
LO5M8/X0Lzir+0/G63Rv07NEjM0M5IH29YVvOYhZnLyFRkqIh2zr7ZPiWADis6VwDxcpFkS/0qZ8
aNJ6dnDkTozsb8OGU9y98fNGvR1n8uVYLse7V77Zth71t1XCDz9w4l6FCswyL3y9Gqs3gEVjYJGJ
o07Rx5p1WFrjkWwl4jKm/canui4+SZQ6nTbX1xBvvUh6FR0WbwqkLDhECiUhPItkNHGZqMv2TjFx
Gl9UzjfD/PWD9H0N/U+ukNeIWhxtg09YehnY/w5PL8PZ0omnDr3Vm/+QF08E73Ls9+wspIuP0kjF
cSNjqciXcTwsP+BTLP7+ybfYOW7VHDiNBZ2AJ4skV6xi8COSQfwNBUpDcZ8TNrhMt75rOejFzDBU
xWUqkFgrV8dGQZT3p7pcNgT7b/A0BRxbgmm6AZUJq8iu3J8SaucJMrbGAm81QivZXwW5XV9Vw3gh
jxBUUDnahD1z1gMtaTB9WVS09Dgd/qM8U5uEG84FubtwkUzoT+grJR5g/L9bMYebAG/Q2R6CW+W0
5af0QlcHn7qT54UyLS+iTqs5crtD9UhjQod/U9BBYWwC66TV1MaWwwBEiztXxDmUfwpXrHXpdm+c
LPx/O0DE7XPOXmW9PP4474bwaniyn8einn1ycOei2Aa6FrazSwe3YnbHW7bw18fCSvBEFFzuhMHM
BBk9Ej0I6j3AlFLIvjimMuWKRa234B4VKzm6SiUt2SN/lIyKtp55Yx7ADzQZJUUeIqac61GzuP46
sxW8vNE4ZvM9PKZFdz4tKYB5/bX0DQKWN8CIMBz0nNS6iPnGlXHyIHy934Z8A2pftFNth3Jvx5zI
r7dxAdyxEIKvPZFU1NLM8shFWJffPL8mvzHrvP2n5WPCVgq68mbHJ6mWzM0EQyU8j06kPwjtzoIo
dNAShiWfo5mPLlVyEEdODgflGitpOgmmqRKLX7P8Liy9QXqcNlWY51v+OKluSWOgcHNWPcRbhzLw
r1iG3CNl+SoQ3F6SiCyW4k0kcxiaPxwGvV2RHN4A6zTkL/UB6h+ggDiA2I9rT+AZN22mphA5YX57
LgscUG8gq9lcAk0VrYrjLvv1zq9L0MIYSHFCsklPn7uUTSsP0vJnExoyWq+bFet4lQBf1+y129m2
ShDU06A3vw4Qs6AtCzUVuJ5mq9KeYvpEBBsibmO7Gq3crpuihkn4vYg5+mqRoyatOgWtCZSdAawS
gn9Gf6Iro/g/5F2wuaaHafXXvBlkLGsUgjIHzVXH+Eh5r8XwpRB4QszKhWYWwIO/TL5II4UzGzxl
kGz3IcunaJIqJEkFx6gGoRXU24F/SxIZacRmhAUQzd6bnSfBihzw3BpmyGD19oMPOE3OB9Q7v2m8
7i68JRy5yBsnjD4q2NL+Bo60Ui7QX5kQMgv9xY00desrSpQ3IK6C5ryKO+uVELdb8yZ75a286Adw
MUe8vHhIcxHm23fUhf8AgWUSXTodTQ/g+GqCdJAmireyfcNQENBvpRfr6vdyki5tEN3FiptcDaGp
KbGq3gkmWm31nd8NYH8GFUe/Z8MpP5cCE4XzwUYcYyxKaTVkY2EVTozmT/Nx8rRMr6uyoy1MTxnR
hjj/gpY1o2jH4lxWxxv4UR0r2aaYqUB86rRDS4qYPhXjsf6fVuyZDOuEQd2H7+HAGaq24AmnqsNC
nRvplPF6Q3/rmnVvO9YcoaUr8ENudzbVR+Y348+wrG+frv9+Igw4dIhJaVwtV65v7j+0IU6K9D7d
Z+huIr2URv/Nb45tmNzFJ89ZFmaqfKztxuFTtOa96Cq9mBM4cm4E4e4KZE+ZvCc+nlOe+QxmDS+Z
TIqnzjFX4YGNSWKc5AMLuVqWdxcZBUzdxU23ZxVX+EWuFV89Ap93IxdmIoxTjFyiEqGnZ/aIgEmq
onV7WjAZBgJetaHQ/nPHBCEqdj8fAUvwF4o+oFVJnci1WhH3Kta/xaE3oHdoEtMojJwSHX+VukRe
7SiOS1iTYh3shP8pGsjtleP6thfacNQFvYyxR8utqc4BLb8qCX1H86rZTqRnKzfSlf6Aos5zuamd
EyGw3M9pTrsc0eBe2BAlU5IoxFpauqkCbzSqT2doqfkTrTJUrkLasoTgegGHZiwgyvE/mU5yTr9H
eNdyn5/Gp49KuO5xaHOrKxri/0eVaFCbj59rNJ6YV63X/C5DWiTrTT1U0h43XzncxUxD/EduFJ9I
X3DLwcvYOkEKGmpnKHhMwzWxNJp5zu8C0z9W+KnRHt3ThDGflopi6H3F6QpoAIWTzeffER0bFOJy
8mg88gaJIvjXTtvbE3D9Q67xKTLCUyfSdEe6Cm9agmbb8OAIs4NpsuQMLr2lzP4HkwOpv2x0NHKQ
T02XTFFpmUEyPrbF+EgnUnxaWDtD4AI8M6JxIN2F7ScSO9HFNGl3MEIgehBMWfVkUV1wJAFNbf2c
REyHxkoSkcLJSkYdtnUSkk7sqdRUWwy+NTeMQyC8/Y5QLDaZosQtmydGwmYinO2EUwVLwnSvRE5e
Co7FXMI+WIC6XokLj/k3nbTwwB4+mvTpmEfG1ChmuNGVVAXOtWl4W89QxR7BNwqmImeOqJkSy38+
Poe6tuvOFxtt/LfTZCqPse4a3SVdmnVG6mIY1C0aii0ty28vlYqxe4V8Xlc9cSmvRv/MoHCl3d/r
5KNOhF61sS6MHd668QW0IRZO7Bc6cTljPJcQiMmS4XBixtR9NLeUI3FEXcW7l+fQ6yk7AGKZrJHU
cCDigq1VHbFuW4V7bFzZWYzr4dG6OEektannmMIVtzJZFjx17k4DIGIIklTB2L4b3Qs/iUSuCJes
jWa/oaGRWxX99sRB/9T4GOGb5TLUziqTsKaBDBKIfJxsNNuzb7QkTE5UyHZeg3IDhXR2OBmCRT/O
MzScBY25ORwPDjy5h6y+EN5SFMUHJ13L+L6iuyP41GC/beD2OLFMhcDg3IsVY0rFFxNyVcrgD4Ya
ZOxIhe57kncNpFLrc7UH1ZqkOzZWhnb0/VfMRJGSUGzOnEtwisRgufFKLpf7+LpSHgSY5ut5jCcz
fLWZCF+2I85by74ga4oEAQRImWOGKxU19UK9CNnKgaHjda7aX57CWgW3X5ytRXYsJTyTfV53rx1X
SxGh+P6uW8/lU4dNHdU6+Vq3LiJ6QkHsd+gk/jEjbyWIlDhuDNAV90uTWBNRFqHG5xHFaihMhNu3
vCWROCp4ZQSIi3nO5FoSVLUpEaJM+WTLZ8UtAJ7dOH6my4q9XRL9lGA6wDMLysWFRECfYrxSX/eD
6f6CmqKceLSKb22nBz9tMk0FhOh70qbUXtCi0++nEGNjKIqWq2+wogZ1shf8l2eFG39YiUddGwjh
oyqTCAk2Iav1KIrec+C23t13lNbKK+CK+crryOmZOH55MRthKTxN0iQbzLp2F8ESxEXt18c58+Zn
3iT1Lo5ypuIcUmoeSCZ9vzGSUdvJtRkR6I3MriT9wfxNnfOIlpn6a/dxZ+LeyjXNhy95BNj51tcJ
cQlvX4z+AeWAEnd6jrOC62l+02T51rPbTmJaicUHEsgBjnDK1oF3dgdZxBgaiMxJY4u3II+JmD37
lfzfO+HzIiEHTfXjhHJ6lbHxdpIarIrVLa0TnVGQreBZy3MWodedvlnhjrN9NOKeRiW8V0/0ym7p
/jyFme72rijYi3Eo6WFUyGtgvinebonZrqlzsQPT/oIK2kqm1L5NoTtB50E6oRZ3MLevqZYF8yvj
MuyZhZII5fTBPYnLpVcEbiZV5E4sMcMf8iBIegIStBdJcY9e9MMr9dXhOJUhw0phE9X+xEyj5aVk
PwBzLjUaGX0dZAkcwts3XV/lBqPLe9iUWjeVc1+sSu3p0N+FeQioqnG4Gghrr3j+AWahX4s8aJdX
hp1YPOd4woN/ENxOzr7r5iqufbFSCfopb5kFVSC0ZXDODL9niILbDbcpEMyLNoXZNCNjZLQkk6nA
EvUmm83h7+tRfgT1DtioqcAiRqMEfaBIlOEaksLWz8bEJ04+ymJLJC2KMKZkUu8tALvdTXUflGb+
EwLhcFzjeGEwVo+MeB0Z5BoIlsStCvytzKxvvcabVvphAdC+hHKYHXgsSCASni12mDKqaZow3SmD
5364aq8xNXU1KjRTCm+cw8cYUXLEUXOxXNf7GakirX3ST35xyLkeWN6PDiOp1ToBVnO5gDoOi/+x
jGRRu8ltw2giGVo0OrjnBhFrYiRIohl/JTLpI2lkuVJ/sY8AjtR6cgw3yKqlxf7MYX/Lv4aNC9BA
iZEnvt3l3IE6TKsqQuOSyJRWMkAxW73+LtcSvJCR2LVjivnRvoeYhHx4Vu1pvOKFfwHrbwUGzPxR
ZweygUEsw1LIRCbwZ57K/OM0OLYlwXamrUTkRC8+dvbt4w4H8vJxPq2zflOjSIR66gjjVn237ZKq
A1UtPzLWPA7G48n+OiytSWsWJm77Zx6vGbWADcMF3+69pESJgjSbtKAu3o/fxdgtiXjpyXMU/v1d
RCOQsOMRNvIKA3nlh4spcIpBbXFg8A3KHoJ7BAqc4wrKwESHDiMy6edxPdsHECL81IIO4UGidQW2
+YGy178Mi+osnBpZqVGYjk3AjXlXA0Xj1MeKsH21oCGWAeJW0kyIg6VrOuOfjU2tTWPCiUKelvk8
MP5iARfjaZPSBUhcin8yx7E50JOcfAAkgpzp8LvkQohVYBXC+Dd7+O7+AdgZSb+QGwIIzD/p3Jzy
bzBjoaM9V+QhaJ02cZmwjJ7uHsDo+jhqYhj8+1VTJd+j5VIFD4hre4TKpfrVb0MgtRkRodpRtTbB
PzRqu7ZWibC9ITX5WIiXon/43Am/8PuBgZZsaMfyapgiDLiXz/a362Uzwy9vM/P/shWpPBxTPJ/d
/Qo1imVkHJp3T/KIrpKedoUAU/K51bCuQ1BQZAzo5jNfAp8K+csYjaui3ynL3aBnS5lgOvWcIcH+
UWUEG1qR82AtH2T0popLJixAJHYqauO2WOzOKuX9LgtZsUOPEasBDHV6OIi/UAvpnJwWsWwxDEVc
YizmIXo1ZTT0etNitfa2JNBZBXfDJJVQsLn1zmDlF6vAQJt8zdgxKeBd9VYzWvT4UQQ24cFDN/iZ
x4kh6eAMxZz1WI40JJPLmdh8LJ8XS5H3kU53BxJhANXbyLFwmS0fdY1bE0jNKHHB6kn7Hi4V39ei
52KJfZlLIa4dodxmEflYz6AxvWnzW0mpKJt6Y5zuVLyIjtDlNGWNdd2v3eoyj2MqkNh6KAFZ3rwE
rF4Ox1fF3gMEn69QzO4eHj7mlslkfCovtt9XUJ0Xg4OHhu61rjmLAgYP8qfRMDpRSfZuclmvg5CH
1v9DF47e7f634wcW4XXzVGrI50TTejbaZSbdN7YJU+0SUT2SBqrQ29dujGhzBBQhaFdQt/U3dfkc
jUTn2q1lUJ6p0sGv8g5X6hMDxZ7RgYeGVq1nBBS7voGQWoY5RYSP6JjgywVv57JbGFkMKBieAx0v
T8ACvXwOzkwtlVyGIrmlZ/cfnhxHbKfP2Ap7FZ7aQ/LLSJPOvt/UBPuPi/vAG2yiHO8a6QzbhcUr
HrfPrj8Won5ckTyUWJqnr+EZ1z8OV/grVnhT4Qb86eSATHLqjP671xaDdnKWe32txtGAtuGLUtZ9
6ClvlQGVW7mOPUC528DgziD+0szpcGgSyRc4WDtRx4FO1xfoge8Xz04S2DcVIKOMjVLTx/3+Hob4
ioY29LZYhgLvIekaw9xxLsG5HO8JTIuGhuNQPzchL3GOWChkiLJCbxF8UVD0AJ7dryFOAqxkBBXW
sZuesxmZ1J1zc8LgLuI4qp76X895prxCV/WfMA1xSmaet2tYDkxTGR8Y0hiQmtsAT9lOeP5N8AOQ
a+R0QdQ+UhVInoUt4cR9+FNhY0GefC7FszuC07nn4Bt7AGwBfMK2sbwzy/m5m1kjDSZiTSUwvFFg
nsBuxkcc3V5ZdjpmQ1nj1m8yRbds3G4U1EJaTJUwMw1Km135LKX55LD4UvpV+lXKbOC7glQ+9nnN
ZfAb6iBvPxjr5eJgsCJjMdg9QYQYbA3AUpmzskWql+kWH+2FTiPxlcwEg29wUxUIxy09P/zY2xnB
aSuRxUs8ZxH5TrdFCIQVZ6TKktC/jG0iI0J6bC+i4wUpMiC6tSajFoGDw7cO0ve5AM0WODdLdStb
ET8BuA/QUaFlAHuGkq9ImVQNcrcUc95dtsq5OXUdn5S/mDCklL8Mk48SMF2RRPFUwDXMCvZIAo7J
2TUU6vH+5ERcPm8L9NUPmeM1jDXTqdXFEmSBSrDYZD9jcQjmR2U8KbXWop4StV41GRjUDi2CLeug
+IdVKLCxN4aBn1nxFtlYekH8lORGjvaPnCvTspPqke1btKeWoYO7jbR/51x8KLu5Vpa2quMVA6/N
3O8z0TxN1CODCR9B5jcZne44fd1WWINTqba9x8wGk0FSl7Rjeya1OYHnfbB32zMHZnjWHEZhH3vK
Un4tfxA4IBlZ3FvNrNIn0yKdZO/HJ8MB7djBNFyeZq8DYIWIWiJgagsvUSs1FoXQr0Sr0etzjl8c
H6DmwPwCUg5pf3mCbkgTgQLzAnm39liQ0XYwXsyOUZvnbCSts2Ws9GWbSwyW8ObEa2ciSR/0lxOq
mvHXxhfYWd3tYc9f8ItVcx3DhJktteV/ZM1cV77aOV4l5V9/qDXYu1+BIOHLulsjKiyUekmgVQR3
tHBOYwB2MEjPUL0fVTAdTvXyldIG6bZ+LwDA0pzIHegkN3DCceXa5eOGi8Pl840/POqMc3M5IvC/
DDEGQ+4CUDtx3rYgxqLzb6rlaSR0N1FtM7YVCW5X79fPs6j43pD4QYcw8z5g8IwcADciLdyuInD1
PW9db0gNQA6QfE+AgdXatatesfKMBlisLZlcObZ6Om5ANbZZilaOuSoZLbyZXGDt1ngJbpJK0Nny
xEYPk9gkaHkDo3lmzlg/ZUI9hS3xBm/tHFy/axg+6QqT0QP9d7B2PntdcsLJD3gmBVL6szulQ1Lv
vRQksY8tuNbObDSvL8n/Vsn91xd/FYA2GPdNX2oelmEmHVUCJA//3EaIjih42zgigzpx+0hfoV+7
5xK/aJIWwJtfMLcTjgmk3lo6vrAuFIqkCPfKKT7LzQh1qQJK1xbXbJGqGj/Qj4T/++rkvAwz7gbk
Dgj2S2kYKfW30s+11UNz+AZdxhKgEibsQ7t3DQ288SGpT8h+Hky94zzks7aV/30dmpZ/pm24AfB4
AkgZGJfyJv4IR4NTe6JyPbiRj4/MQRcxHO5fpGOlST1CUHTy6rDutwQWQcEcX1X7NBZj70khAJHg
QdxQNyrgL2jXc3H+peoQY0lLX4RTI71xNsdoNN+0SMKi/QmVBUwV17HNX6AlSYgSa4aJ95m6c9/6
n0WbqT0bv6IGx6Idn/8exC0Pc09AD6wgufuOrN53qYu2Nhq2YSuX4MyQN2tEwe8MqOtv0+bG0U7e
PXnyimH2zCyfO0o9sfFOB3388cMPGb65MMxo9XdMP8MiWTdO4EN5t33CGbixz4p+YLj7W/Cv5b+9
3Bp+/8fHSGiJa96gyH3OBvAON+FCbi9mr9VUS4BPV7HfivqEmAyiPzdEMKzXZjjSXk54daZyMBaA
v0nwgDxkOUB/zq5BYYYzraxcqLWmYfaxrw04Dull8vB6B+eRE/fSxdsOYAZPSRcGeA8WIhG3KRJV
TD8R3pzAloknsSNs50jnPjVnM7wjN0UH1F8VsFybqbJRwQJJ8il/lhaUe1giHCh+QPdIvhh8TEmB
DGS++fYS7qXpiZk8GU58r4Ohj3E6XD/mIFUV0M6U3Z5TvF0D6ibAMBY5VVnZ9GeqMxkWxIA/F7wa
HqTayrsZ1YH/ovZNkuC4RrBbhV7U83ZbOUMyWE6t2Ew/vo2v910ZfUD7SukBLUEuS2Kkb/01ymwU
Ek1pOhhYh70Js4n6WC7akl987VsoHvoVl7VeSM+y4sT5T3xTa1zWo8+aEjsMmYL9udiUOs/9+P+V
7fdoIz5Jnt2do1HRavlIKoymk1HOYw2W32zvDJlNuNrRvum58qPfpxLGl+JRPaiuo2UdAixQtm+m
pyYJowJS+h25QivHcwFM/+Cc6V/vCDzPX80V18a4u2nLbL59En90Dp+e8jGhq9Xb/ZkL1X3/albZ
G2EVFMZ1aX+hW+9ULthxB8LzdqD28HgvMpim8UqXMICRSkDZCSzdYOHImaEIlBVKejKr/Id+sV/K
RDklxvtJeRcG9Gn0LXFE748PDYLtTC1lF0MLgqn24d2BZlv5xqwpHA7usfxSOSlo7FYiJWKHCCMo
YFVQxLP9b5iRRqcNeWxcEdmKoXdJhefyiU1d+ActWyxILB1rSz4xiGOZ78kYmfiIDPYn5ABL3s15
toqeEdKmcQJuc2NH5ht7SKSBQl7EtppMmjIOH6Ps698qyo7rLY3Hfoa3k7RhlqBXOny+CuMSiVbr
Y0qgu+nAHLx8FI6XqVo0UCNZVGcqivkPLGLjhWBjndlJEz2IsQwnKhmmMkD3bfs7MT3KMVwo11nH
dKJUNfMFdIW6qfg5Z5l8rsIiJMwUy5T76cqk2E/ff7L0Au5li/Qturg0ZAQgZ6g9c7qLgs+gU06R
srEjDKlcH6wN8+n8m26WNIRYqscRpWmmwe0wzHyYnxwAO21SmkyHQ42vCDnc9V4lVQorkzRdImB+
dPz1OurSKDhnyV2CpIc/zmhglugnKrf78EhvXsjtwwqIe+GjHK1RoWTvslNutp6YrAK0mbIH5Hyf
Mm6ZH4SqyWjatPwUvW2kIElk77LUWdiwXerx1fZhliiFIEhcr8wqtaSDWRV/yltROV+1LYnQJbX/
k5nB2u2IP1Ju5Xsfgyq7/e/rrOUe+pd627TDbnF0OnIZKI5lvtrvOPHFuuC20GMCUDcH0kNbww/S
DQJj2PwIHQpd4qy4OAVxIeTf2ibUeKrIvkvYVKkH3FERlCNWL1ELW5S/91w/Y8HAqC0PlyUNO5+2
+OZ4vdkkjDGoW1c+pHWBWphnnsRTDg2zf6sh3wGxyTxJu9A6ESri/rVUryxUtJHLueU2kNWxVx+H
zdkEVJMC7vUPywcjM3yqofmww2kCUPqGEjo+fpXk7GmzRHuBMTNxiANjwepSW+HMnM5RjqgmdWIE
6efvpXk2KtdMpqhk2TS7eDZykJCr2B210PB2Vu9eKXYhyChYPMevAk/wHwxGWvE917XpJZ1w7xVb
ADtSJWQsnQ5KY4qeQyie9thVvbHNVOnn56Wv3LOTFa6w52nL2WW+ARhZbL/yVxPfw+gTDUWeOpnc
ALPBBcjErJPlT1JfFiVP6Nqu7w5lqYx4FBnpej2T6Uapr78aN6+I/hlyIr++56lPf2gHT9MpnD1f
W/SpRSMpo5dEkirmPG+yJAkjZVKHMt4XatoSLJpbxW5cQ6djcBgSo4xb2HR7E3I7Mz0hb2NAwMuh
F5IAja3I83E+W0Dogf3nPCHIVCunbfnKK5TI2YoSHlZ0q3gxt5kTbMvc5Q0QbQ3QoKLjkuHsmfQ7
dalpwvcs7xiBgkiHVUQNjyFJF/GeEypOu4SlZZUzR/EyLPT80AlqdAqPjlpBGGTJ1HMHk5JM/5vH
skkYCkVGvYDwOGAIAZhRuEz/kzWBekWVZukos7221WTjCm+7I9wy5eODGbp56XFAenN7WNNq9AP5
f/1u+0fSowl7I+akY4fK2FUVkAxXpq+/I6sf3M6pDttydE4yPGZPpPGNGjPaKb0VFcSNsT7QOHxN
LKp3Y9fbHWpskCFgEf8x0LOlz8qMeeNzWP+SZmOqevcLI/u9P6XYy1xbT1SOjejnP0T3zFoN0cGA
EqizknVU+c/QkqK9JCMDHQ8Bp4Low5bBzNrCeYNjC8JtDmYML3aSKMkvaicyBZrQoKJAJchFGv34
H8UfSJ27nx561JnMENLuCgdBB3rQ+BjDoWTPT3ZBJZHWNS0HWpavp2b9CQj/Uo4DOHK0/vZQgrsA
1ZGGJ+58xfIvOUPIOOsb2CwlyPwEGPOOLxnvtOVo0yjy2oqxXQoXcklkWjNZoS1XVmRCw+U9xodX
5uZKgj9TngiFyWd2uSwjkJbfJAur+qF7Zw5/QiooYBBva7F5gsN/DHM7XL7fM8GlW0iPnoCoSOtH
M2uqpvC3Re5FNjSRl6i0Y/ZikogcsL8cgDMeFyCUft3Eo85QU2jP7YCfGjMEViYHqvs328vom/HZ
ZPHD1mOpYMpF4/zgVge5CBiW8BAgYbLE/d+nl4MlPU2PXUTvYxUVcqVdukEmeSol3VoEgRmxlB4v
Q+9gcllKQJ96XLjs5ypI4PQMVaW8ooyA5IYIePJdEiYYTCWJ8KTQcYMA+hxlPkEluGqyJmyLz+++
wVB2AT9TOYJm9+qBDpZW9Mxiaj5iLiI1r79PvAZaDznUIIMyKZYirQDbP1szQcjgU8spxPZevek8
MePX1LYZZ+r+/P0/96emis1n9E6q7eCVjIUBH1jbciAuo2HYmmTYaH/BK/htjK3n5xRTtEYHCkvc
lY1PeIL+TYF2JoeM+Tdm1h22gX0dCOLRua7R6d7rjN/AsAlrBhmn6gsWLBqVGmKAlSbX5L98S3VX
WWC7gc5jZ7pQUFlBwWNwbKGqdj81/FfohnxEdNYmAEAD4+xOaIGjdBLmz0vABOznkbCAUS6hdas4
42q50NU0e2xov/LXBmCEOiG8bv8DaKIsBT53Z7chOVXDKkVMxCZQydL3dmkZlbIUntuGQntSeIru
Yn3FZcDmUdfuvG9MvL8Fp7vCC/fT4iGglJhgbgclH5b9Jgd/fUhs1SKboRMKL2UnrruBZLHR8QFE
MG4OkLRiUBiJUk7A1qUhTtY3G/ttip6ynt5odnp78RkCvtQ071ij2Qo2aEY1HLYycgi1ICfN/k19
+JJVD8UQC7mENv2pIEl5EvBhR/9gnMI/EXql1DbieZ/kHTa52aHn7kw12R6C3vXjnQ6o+Wvifa2d
AGwx16LvFLY67N++f8jDZTs+lZybIkDdQcptkkfg0g1H7HUi9/Pr6quqnCdduauzR9HwExpjqLu5
XADmBWvsv8deHn+6t0ahRvihbBxBdXuwWhxLoepP6FhNazenJNz6n9C2XhEwQtISVLTN798s4Ue5
BVXTTzZggmlmhQCSerlBEFjiIPVCL/W8/fIAfmrdMGeaTYC2H5SpADzz3aii0XafnO/b+BpO9fLi
oNw05q/6RYmZPrLn8byHNJhG3y5IX5UiwYBr17I7e4m+Wkmubn6uoKBrx5Vg+l83HUfnjsjeQlos
nf2xKtcFE4+2UA/8WQ9Ng+tOIIMae3WSmPOYmlqObchq6Ox/0syMPYqnwey9IVejZ0fcGqu6CYT0
pQU1zZxWbSwmDB9ORoBo+2oxSbYOEkuBZ89Uj7nTuLspJMEh+aVog0ZIJW9imTq1L+1Csd90vBjp
r6NEoN81V/Fh3n54ztzUttmrGn5mxomELdsHgj2P4cpoOx4LChlyqZg4qAUEA31vhmxqNDOYfbB5
T1yk6TMgklz2CTEkkc3PzS0QnJoTwrtbJuGz+EZaSkqHle4/MT9VD5WMeQYYq8uZ3T21AC7uejWY
h3dAbMrIAbb0tMkcQRi8jPjFB1BlHg7coRnJA+xcCtus5JXxkhczrwQi+8lz0vSOgokVIgECj+Cl
63AX+EyOWD055RHIb8qQiWk/F400uJVGe78OFASmeTh+pTwUrSxYXr51MNgFfv2K/en0uoh/Lbdv
YQTY9E9ZHgD4TUz9l3HWFOTRS09I5exSRU7BgMZDMPe06gv5ZW61gz5XP/yTZZl6b9V0LYkQMHQv
wNd8wvrj9Q294N1WpnIqC7zHF+iBh9jH3YzXjUdxZ/etAbOsPKtNENrufyAIdlG3tafHDuoHBr+X
m++eBw2MJLFsY6R544vUniNfZBbq1CF0w111rMcYp/+MyuiPskENhHpO+TI0MBOZOoykm+x+jQ1v
KfL5RlY3Jzqv126BnuP9qnpn7akDEfVIuODHGQO16oh86hTIXu+4hHEpawh07QQZwFSW6txFhYrA
WjQuecQyDCcx6JTO31cUClrlMn4HXydJvcY26qe7P8gttVzUAX4YIXQtioRCntmFSY9W2RUKrQUU
PvjNMbrwdhTb9/XsNyXuiveHrflbo13nRa66DmkZpxoh+Ta38rfoNpM4MoXreI3EJ2gOhUrHtKZU
5i8/tQYhjCUe80Zu+jxZWdwrwbwAotX+pSipumlCEnx5psbw2HyrrjBhSfGe5iesa0vFxJnrdQ7q
Cv7ZqVdHRDzswa2m914vM+LR3J8zxREOK3fD4I8Pccc5abND4KWXRJqJlQYXRhhIG+ERDsqPEcR+
++fqTW2259jrW2OYn3RddX2vLBuS1NFf4Wi2jB4P+pm+2Ck6+nmFV8OjJd1LHQamVWUJzXHpkeva
86soCOrnI0OEFD6psj81HBFH3w70nacSVCaBveRMar4z9LOl3alXF4sN7mXDx9pb4PL9NyngonCZ
xUF/8cqw7ospoF53nBuBCFQ+jc1g2w33arRUxqeiHQucgsFa9zDewsY+ns4o/n63eMaoxcEfH/++
+Sn3Aj1bGOOw7Y7TQz2R1Fe+CqmrpqtWqu5YkqMzqSzcZY++BgZgi46sd6JxyqRvRM2QCTe6iW8r
1vp2ONUtPS6VzjEj9f8UvitfaTYKz/Y86QTfuiR8EGO7K/Ugjr/a8vBpGYo+crPurc15GRFZRCts
Zla/7uS6BENTuUwQVQTc9zm+ZDxIqv1P2xMOQFawl0Z/Qf0KGgOi29ft2hETT+Wlkh3vWUbax87o
S1yg5WOvCMoKzQcaTuXwyGhdZJ7MU1Z09JFsPl1le9hum15gKMLGwDtbDG3oPPcnAZWKDdhHpoHg
UNhd4S0X6bpDOTfb2VPpt5gslOFrbw/crouXuBcB0IRRmxnKT5RW8LGscAUFcXbxc2BDoCBktmCL
zTcWVySKSlH9K22Nl0dV29SyEkbsj3GDvDm/5SrwhMeebywuEC6PIarIsMklyth8UJkr/VD41ez5
oHSrj59h5h/iKmJEyKvS5hrZLLBJNPWDF3uizcMHe/RNOo4tBEjxr9XEfvKEtEmnX/9WZGaXwQZl
j+cWeqsyeuJZWYkpJxxPYsckx5+QtN7cHbbtMPDvJwLgnvPjutUZxO70r89vTx5A3tFR7aegHS9m
RR+KJyMih/M2mD9PcUfAodFssMwoQtfSwmglkdftGlLSju0oLlW9a83rjKzRDLG/L+1iyv9WHF4V
2NdV81cjfo5AHjN6xUxHV8QzW6O+6/nDFWt1ixMCZ+Rak/ZAs1cmkD+CJcvk0JTXWTlm1xWl8UrT
u28VB2gB3bCP1c7Y1aUo3ZRGQx42aZMEs6riOnvwfDlltWdTTt7Xs3ruAkpHuChAdxgxWvQzz0ZT
FiyJvau2tgzjV1IRNosmKyv7i9kzQ805T4P7RrNdQ588b0C8yDYawCbpq0AffyfnRmn7uzLqPfQX
UxIpJVo1R2QJXZzJVsTdY3SlznNQcc8x5J5dx9GldWuffW0uWwOIbktkzu0RP4vXozlrKM3dW120
dNMA6xmu9lW/IiJskP4szkH0BKHh7E/7Q6WZLAeoSz90h3uUXIYY0e9b9pOppu+SAK5/9jMKR8TF
ly8cdBbyW74wHsC0gAftWG1rnnV9yyQb7X05HI8fzVXn9ETlFcE8NPnawqhql2tL3voOm1FIJVGW
iSdsicoMDs8zdw7e6taOBp0IbDYIhMW8qrxjlqPt0bU41Iy52d4xtHPhdS8teMtAtx4pdzRwtYRg
FAdq7FRq9Bg0q3qppBg9FlkeVn+xBbLzl+7JtBUaBC/BbbYMs7vzTjCi3RwbXQPTYnrlnz2n5moE
2bKsmgA5iDWgh2QyD71M9Fi/pyc6Kypbj5dMAm155xoBsqShy8Oqv3Yowv0cM81WBe/BNmDN1Lqn
H4c4rXF8s3Q818ZYdudkBhUEN5/J4v7xLz2zwZwzTpLQadzsTcBfH+hF1LvzQaKZ9krgh9lrWlOs
vlFb2/e+vEXuJG77BJXu1c4WB+5p6tF3QT3hlsheL5ivJonvH0k7lbnNuNdn0LZjinM585ZoNDUh
GGgRjcFNQOlb4+zf6Xrx/ypIi6TwZfCOhspEMSgmWV1T2hM7mPvGUOL5kS16fEGc4FBFxnyEntSJ
sWFV8w0x4dhQHPy4o2hurIJweRjUaavUtie65oJ9AR5+KrEeXUaH6usKQ4EDt6G4UgzupL5zQ8V1
HnBW8h8fVJ4CtXt6l0lB+2/90tHqcP0kCSvI/UAl/qTAEdv4V6AZgeeUKX+ZQ0yYiTloFUNgwRPF
vsQHEDQw7WsLmTm3JPU7yCR7wAuEuSXJfmdmr71zuxOux4ZU8TTMiQQApirdA2dAPjOjKkPCVdN5
07WX7rkUgTIGwwj0JXQjd1Y4a9K/IKLluMaH9y40MsV0CItkbDQRN4fUPpNCcDKcET8Q2Qbr9yvJ
u6fsqxGTkJNKwpEMPKE/hC8f1IsI72/4L9aLHZyvreD99mZ4Ba3lwouHbX3D0futSYzRUJbEq2Za
tvR7TNyQ1D9FU/mYTOZU2rysC4F8lR7EX6oYZ2AX9Qlh6SEz0SH37E0TrlJx/BOrAh5hdARYwTnn
4zwWRO6jN60wYmJ/7dqHXk1+1bCC8G/IlWlkCIl6HqKR0I7MpI8WZOrIm/xjwQ/KYxT193TlsEKi
tdm+jDyjS+tlqy48uXygryZCcDKsIkDGLNfR5npvV+spPSXkMeGPpbRf54dyRb66WM6PH1gwu5sd
ua1rAZz9hM/r1tVKPA6c+o92AP/oOag3ASSjLwVtoCgRzyicuwBEDJHiRGauqzPEQGM9sBRodqrB
nngaLoVrI9eY7xMOF4+dlEldyGcTfkzc22Of/hzbAICAS5xiyuhvuOAUmnEqzcXfPduStb0+yPnn
CUCGXLxCibdbVfdoZhiNHkSH3o/KMK89Z877JUgB7Y/LPbuDz7yJG0RCp+pLhzPS2HImao/v5cwT
Ep6d8x4Lb/UDL2Xis9lrzFAHYqB7ah2fMR7pN0Yi/QZDgOfl6QP6KKgbSudiwZlOKehKq9eEF6Ew
tb6YKGAYxkP87DnxSLrvShV/lgrIggMS2g1CVcBmNcNMmN5crPeBVPOLvAUG/Qnyyn5tdydP9/+k
ybGm1ucZqQtuNys7pcggl44iB8yVcXYYnawH07cmfe+gn1LQp1MrkcqJelQ5ZPZ37e3BuSKcCwie
n0jYmCHa2UKD13bvulCZtsefwt5wexrpuA5WRCjSOYW03vWbH45/yqe0FvaOGOTRTNcNNGRj6y17
QaXD+CA24QDRtiz9udcKA08ruES/pAb80Ypwka/z8qjtbOVFEQbprIF8QlYMvNMQGLTyEVY95j5R
EdZkrLVw2iuqbmkj0+4evBBOGcVn0W3uS9JcYiUa/hz1b3euL0jKdMDzTLdgq+1nfU9SBtDRKrZp
l118NRcEpXqL7j1T5fAaRKg+BFAq0b3mLTYC3Tjxoa7TbCjijddOX9/JZXqM2g0NHQXm97GKQY8x
dhWBOjKYGg2MXwDum5he/U1q9TqluKx9q7QCqvKskdnjyG9G6du10wfJXKYuioJ2Utym1CnO+MSf
S5onhxFLLrPw0OujVfD4Fifa7E8Jpe4LMUzdlSdU+nbt/4OU+vi/jG2nUkmxSdgb5C3ZfDGycmpK
qy+eS9IJmy94nzFRLN7AmuyTfmlMLp0HXlMmplvL/YPGEre5+OGWp5PvrYqk/DJ81hSFkJIm9stc
gx4x28i3/c8yiccwEnU4TpcIs6N295z9x61EtAT+H7iCqvxvN0KLFp0NLSaCu7vJP2+6zYH8UO5U
1Hbecaxy9xYpwGXz74BEV1DGBNUzj4jD8i2TE2FkmaDFa0DMzkmsD+CrVbQYcwhW1VqIWZDSyQub
1MkReXW83PP0iuseL9FNXuoYtZ3yCI3QFoveO2Ds6CBGZlVOU0ueN54YvyTKKZ263BH+nz42ILh+
uvsoyQxKSNBZiXmmACGtl8WV2LypPfPw1fKbyPwIYDeO88GNdsbjCibed/wdmPlViOOOhIi9M6an
tYwH5vyZaGEmMYMok3q01CCHTpcOSfLE8RlWefyZQZwy1k+KceX+Dcs520IjCa391G9svQPuN/0Z
whwtts7Uy/EdW/uEZKN6+fSCAB4m2vLC9pLx0spbP8+88yHzaiBZ2FGLm2o7/EU2a+5k3cE711uM
ccf/KKbf/AX92l7zDiG+lJhTtzqfYiYNMSFLlar1eHueFYfKHmQo4MCwcYlHRoj0fsNLILCOrJ9u
2OqgBrBlcQi6NhFXd6YWKtgMdYgJKpW4jr8kskvAT2+jg+5nLtXgAUk8U6E1jBrqPqpXdqaWt5fE
8LRkYzId/7BpkTHszltcqMqqjVBNrYDlP4HA3SnpC/fYSXTH9bh7ufSJ45jfPcOR+/whivOL3tqZ
s5tHLld2Rm1MRclC8jpdMqArbsnueSe+R5V1C/C/EeI+ZlSytm1FcEZo052JCic94pF6UhW+4cH/
+ERlpXfRm9m9vSaCXLMS6iBGxv3lWkB4zF0yZKn1xiYl0LH1MdCO9HoZaEmDcR9/Jm786Y1wwlQk
xYBDnL1fRPwBEpLvrcRJBMuC1XPJd35JqPZkcxTJkubyqLr3rRfjSrtwIVUbXJhmNCBmvpx+zAOh
yfX0F9ofYkGv3u/2MGyYViKxBmjrk1YRhN11CEvOGD0sCkgeuXLbTX5dljfdS/l5NFsChCXIn9sH
IyHNwxDpD7qIsaLeX4BXb9LM7737g9S1xTJHUia0KYdl6AUy9C66Azc0t+yGM4z7bVQ7ImDtWu4W
J2Uh+zmH4WR4JlQgWl9qrLDAhZueoOTadbgsPuVdPqzzxRkUIn6+utxLt1GyprGDEVfiuBVWTGZo
wNZh68Jrr1JwXojbiHRavQJTliSg4a+uheCwt9KkP0vW0lK1KXLLYhlBz370LyEt5TqT6ovv22lU
vtPEGyms1ZdhMdhaYmDrcD13b/3kccanMByH9oN8j3aa7V1a2WyTkjHA4ys0iIb46mDA96rOGxZ4
1V1Yk8p1SlVl2fIyjCJd340lb6atOpZHMFA9YN5PB7IDrtnR4PqyoCtbYm4jiZM9VibfcfNgpdEx
sf6fDt2k56eP2Ez+QGMUX0kWeGc6AHDoBheqDX1BF5QfzlquwyQ7yL8phJEHSR7ZrnH6jWzZxz+1
RELpKTJAYRRtUu7yN40MRY0kWuWgjHiBxPoO7QvmdpQYXYc1DMyCoDRcf2jDCforitwCWlbuPjH4
dWV5HnM7roS6/Vq1f7zvJaGnN2X+aibaSEMtga84cx/8IeL/DulQ+MNx0g2ESUiffLoPQCxL1R5e
e7i8d0As8kq9/hXmw9nfhFkEtDwNtR9mS1U5Qtj9jtWkhlz3aVsU+j5QoFzldsYO3jcOVGSmgZVG
vyivr6wAfV4UZtnfKxmDbMq9xoxvLOFjcTafSphxGQ3jK/nQBmLiXz8j+JyTXbBM1e9Yuhw5vCCN
aAV90wc+BIjuo4XDFYP490w6hXsjzqamBRj3KUekT7eyTxMX1U1GTiAJI3FW1r3AcB2sYSW9Vtci
TOV/2LIOQu1z+b7c105ORaJYzswddHl0mKbd7pbGtiEBKGLLwNbbBnmKZLsLMHeDZQ7DzKKIX7En
fo86tSnIq4lKDGbGFDiEyH3EE0wMgj3nfkz+AaSyZu4XeOcLJ4p+mypIcjPW5tS5Hrsk8fLXCksp
QLTlze6uzhfQWPwGNPOXcXpLKTs3D8r1CaCBW3p/uC7VeFK1mOB0kmhZIOw0PwsErUOlPrSEmyzi
kEaLjPv6xCEMhUG85/4Ez0UXIGnrGpkI4xY1UPKfxfd7FbbmDAS5Dk8fx96dWJU/R2c0GPjAmiv6
oMjp3Ha3c2Ne2dg+/cOKDC6Rd2wr51yvSp4mmyrlfZWnWG6i/F+sO27aB82MW9LLIBKQw8RhBGVB
AWpmoE5UjRZgPOF8wsXPlvYEUBuowkJRAjSqCNsn7f+Eqla3AiOp1tIeGIC9SLsblnt8qA0tXnsG
VBw0lX+Pz4oQ16YnCvsXu1qGngP28OMkLrnyvTqGhk2YqQGZcv6eCnmVdVJgqblnpDanjHbRarEk
qAloFyfpxwtEFu1AZgMqV8pOYcuJJl3Ch4nBMsM6GWqBpzGAFL1LmczjLN6aJYXAk/jgQb7oO5Eg
fLh3rKKEqKKH5mgtNLhQU15ybeCeBw4vFLBmptGGd+wihpQfgOzHQF7R1+6p45Yczpu6qg7ZwbTU
tN1q7zLW69iGy7iq+s82PM0e0H27P0IZud7K4F2N7BG119BIeD9X2RSfkchQdzJCht54CzXwqbWo
gZjwk+84jIu2I367SiS6+Y6Zcd21M9sXEfpStHaDbIBm5n8bQ5uLszpAJdVT/wJVGz4Wm8MEot46
MW9IQQCJw8IHJOUTOcz5j0wS9TNqQy+HROoLDPYrmjr9QpuaRJDdNAXjNoJqpDtyAOxqR63fzXIk
7oT7uzIxNSD+y8dThP0Gn5grkneyzy5L5ZRyT2YJ/pXSjGspbTXclkU/WFpLIe7bvtUGeuYaLH6N
KTe4RbM3bLhNGFEHwFEKBoswiTYA0M4k7FX3M6jZuYa/8m0JHAqSFMmusOQShcnjm4JY814ZQq3F
453RR7tJpoIJjyiEGh9QmqnGo2rcy17N3e7HZ6X7OJL2GD2mSZdO8IU3VExYmwHjj9RrHBr8vHi7
DhFiMkq6NxXagZoVPcGpfSOWX4HVeikdU5A8iOB4q/QGZdS2chNUSSRGxWnEMkJ2SwdWRGCsPOy7
qAyUoFequIloQvrhU4buxlXJf7BYaKDr7sz2BOqwKfP2arSDBy+H/rV5d5DsqJDDVF9SUpGS1LyM
gLdfIsxvYvPcWWvZWthSMu5TtBcZMorm/6v4scDhStl2yayMZBXV0RqcgOP/ieqVxW7/84w3i9JC
D9DDz+7PG0ecFPEqouGgfL/OFnw9lEQOJlfZHshKfUPkd4kGc9lF6n2Qgt3sDCMhFWHfj/Ixjt4N
SklrnjPPD+Ow2sUo8F6+L5tdyzEBayWcym+3j9GRbh26L6c/LccRaVMphFB83IBXStoyxOAKDKyu
1LykPgrqvkmbp6BGcZGg3Gy1PD99Bz7HqX3H+nr8tTeMELiE68CGcpZcnxHrz4eQHCDPPI/fET7C
9aDsyWmimq3kSKZJE9UrCSlfNUDG7vF0ANsFJhI2qWTbv/PSUDgNlwb+onAAT2fKq8XA9kNtqwun
KyMN7jfkqkZEMVVlMi3Hg69YpZ7WAN5ymspES0Bu/VpjdN4XEPrxcTZlXMYG+4LF5PL9cZY+dkcM
KvW+gPPc1wBRRRoIfxkeP6ZWkIKwnl4Yo62EyWt8RQ7YVJ6in3X/ds86hgO17MUQ5sPN4otUaoi4
vgew5CmM0mwXy35Npd5FhVFicY3mjbSXRFZdSoYZ3JBVecVjJ6rLS7T3Nsg4kGb0X9dgqRIwpeXK
vdDU74Eidj/khA/iWGWDVXE3QEKHZwO4JSJ9sDC0u8jV5HH2KGx+UjDjqTtSkZbhJTg5L2pavk9T
GykmYpw20pp0RnWr1LeocnHoeoEiFns7+pjQJMe9NYQHSJe9xEcnA18foaJgUK7LLrgm9HcnfzFt
EGCjWITJ+OWoED/qlqGy4lODIDZGswjke2Lwq/ZKbQ8lytfHrDjwsDuo27XyhXD048jDpK9nWXHu
Dv+VSvx8pVScftjh0qJ77EcLXmJRcHztD9N1VtHYnLB3wuunXLS67PZaOWpeBbnDKF2/4CB7S1LZ
MrDxPCB8UHZAslqz/QHdTbdgk+XYvd8jUIddmQucm/D1SeGdKEVgMxFDnqmkg6jmkA/ZuSSYL+v5
wRzLRMDo29uLyyp/pBodZPCoQ5sAoagRhhPOEWmf2wbxBuYz0+IITYbEftaw4jDKICnhjMMNrfKX
jEt3f2CjeOD9ZzNbNZHbLZ48j6amKFvrNFhkC4MVegeirgmXTP0WXE1pSrd3RFGQFyLM2m2eFq6F
erqosx301Pa7Fi8SPpBKSzLohOi6IOZhXpCB6ZJ5picbCMSSFlcywFZn+3u1AndhMqS5eLVu8sEE
zttZ5LK99yoX8DQ76w1k00krt9Zl5SvXC4uhqfmXEWoJ3Xwe1KAntZakq0+AB5Fsq4cpxmTytRT4
SKikkuh16nao9cCQgh3QAqvSl/MO4Y8sjaA2ZZlQajfKJCToFpavqbcPyYMNJmPNddUC4UduGsrJ
gHxDsGDjeNTvAnA4dbJvxgi+8fXKoUatwXrgC6YUdibaDvtb75bRHbvagi7WmvtyVs+4eJJ7Ju9F
V2v/b9aFdIX63Qv1X/3euLRA3BFZnM1pHjE77m1lhcYDRFzZfl1uUg3jKhKFno4LWTi18uOAmhnw
A9nebGuff2qEbwyJroxpBrcFVtaNtjhkNsw+87UVWmDQGW6yhbA73cUbPL0for+li3rwOCZzXBSs
pIeowx2Ndg3MaKdobUs19+ps0DsliW8+tE2OSSvqDgbX/kBFpuUmMz5V22QD6nOm7GdkySieoixo
ipIPenNF2BZ3GLEUxIT9/tYomgXLO6EBneDQU97Y7YQInAB4W8AyYSd5Qup+NN/pogp87P0RR9bv
LShVejezj01hA9YBJgFpygfNi20ibh3rIxsXpQCV+UsipA2ICHE8dXsPzxiSeGJiwlCSPgAtq64F
piS4hSo3HF6Dfqs+YrTdT7MYOt2tvWdhbQeHAaxZhGfBaY9HnzYT+zAZgYyEi5tP9KwHBaoqRGJT
PfwWa9wKoXN5FA1PEeNNWQepU+i1FQ7maDYNAF+Vd67+T7XR4hkz/jEb4LytUUqUQiPn1OHiO+0U
VzPurlfdcrQ1tZdFE8R/lAQnRkDtp3ImbEL1qY5kKSdWqLemVobLeX/YmuN5WaEhISe6522vTBlj
8/ktf4SwbNwzN7Y+UCybJ0flpe5P0+Vna7ygCdaJvRAduhmN7uNAcEMVTBVHTD+etZPBjeZMXFlF
BTkLJhOxiM6CG+VkWMxIZJgwi0RADf4pFsqknurYMbSw4nVu+34TikBhezk++4HtL9AFS+jGc+8b
4tEz0ILsKYedhiBUU90Vo26HRKY0pQ7ZLMH3Z7gJXix7YU7ehpgRXEFwZMrbFbkY7ksl0ynDtl5D
xu+qxYGzTfi/Mr/PFxjQ0Rcj0L4Z7zp0oTFFnjXfJKZP3X/Yz4NM/nWnJLZlgboauR8/dUt4nSU7
5eXco84pB3Wk5B/HjA1Q4ZIEQwWd91hpnLeQ0u16Ma+aOJd8EMBWMUKmEPyQC+tR+GwquLhQAmY6
nLC3akoIzsR/iBthRUhY3tNjM+2m+RJTzuEZxt6ixnLOXcPwDiAovUrszHm84VxJ3ciI2V1IkSGc
YhCRlbcwIv6hP6bbDt+LgI0ZPyceB3t9OfWcNp8x6keefpU8Gt7d5S5jihBRrJm2VUgp5LdFn/7e
QC6z/3M3U/8yxLpps5UNgIWIDEM+WrPlyb7I+yuJ0PAOyQmxBOeZKeuiAbNCbqIpR8IIJcOrISLX
x3yzW9SyRkaVp5mMHj/RoOb4/qioaUwqwXJ62Tu7OsS3+LSweIu3G/Q6BHuBbVhIUO+9z7wcIPUC
GBxUX4l6ZVJm73hLnkv4/vv7taeX2wDp/SVhWGBrXRP9Uyi+ZD+oCXUC8uwAxd0Cl924RQZADI/W
hqwBvfS9edah4IdN0quQGATcTdgE2bDgCfU1X/JWL9/SMNH+AyJ2RUpFki21khje7zA0i/qUjhb3
WRxLgsJ+I6iQ4KwecrZY6FTUZr7Uvj6mYFMbiJeFzIK/+5POuRx8ZhYkteqkitGl+8hLWCbIjn51
A0pvb1iu3DUW+S6Coxo2jCie0QoqmEbdZcI1r75LX+lf+Kr63mif3Zsqd9EaUF9ivMZ30ftEbDDb
F1Kv3gyJVce5EWWngAP5JogIEUp4VUO0M6KdEucABDBDeEfqWTtnEiuuCGpnw/aX9MPOLrwoYc2b
5oiFqYBuDUw5+n/aoYigmoqakyJ9ZxTRc5WBrRrqUUVN3MmHMggdDrUX+Q6YhoMBKZ4aFtgD/XLl
Wrf/YLc7CqNgUyB0F6eyH+37YnnilvyXBRgwgz1NLKUsKaOh3AJth8f0dWI8wf2gYNiuJ4y+2czk
6gfamboCdOPsA3HyeJeZLD7bZMc4cEcAV1sIkxxfnhcf1m7YIGfg1+xFkotuDl9CmDDe8kLP7aW1
kbRb5OLB9wfJudi24PuqaR4Cjxl270h/b3QC2S0pCZw6trVqf4o9iPLv3tF20l4w0fsD0lbFYbwf
ifqy9bk2IYtwQj8L1U+oXHhRxJ+ifdeFz2jpRBLfONV/kbym4T8VtO2RUMZgnQdZ1vuTKCyhRiQ9
iOsGAm5mM8aXD3BuIwaTOI+BnDYGklxastlUejymJbFMmdYjdsZ/2qZSwnuOwqKnrUFidoYrXxDT
AfS87NbF7pS0eNx899eMHwf7CTyjlLt22yYK6JUtJ8BLxbaccBenCy6abw47g7uJr68Kj4UDOfVU
6iSJIMC4QJjgoJJQs6zM2731MrQ6oNgxu144zYq5hD5aE1vkT7yPi7MDkkjk0SvU3ttM5f8SxYUz
R4jHaLvJpWPYZ5mWBsVsIJs/jAy1jRGOawstFXN3UvpwztI8Yy+5NFnM3J3dV3iFGOH4RkcRL03U
snrjLkepERnMa0ysOGRGkSG7HgFH2erDHKvPZ6utSdGPUrkRq9s2Qo57jrt7bvSRKdsmNRlJYx9W
P+6LYlO0jmK5GZaDghl8H6gt4yXs0qEYtwUDJrOPvfc8kYBjZ8IOozP8tZONYJMjqyVQTVlH3RqH
4LWvTbJF5TpfUtFP0iBdKc38P4lYsvF3JKFFfxrT9Y+wi/QKoxiggCgQOUeJyr4DWRVjtyXIYGXm
Yldqirr6q+aL8ipnh27t652PIHfyqyAgnNo6VpGgwp9irunhGJUlD9GLPL19sQ96G4IDdfVpr87r
o8pP6goJfza2mQQi+etEhNxdsqtlEhPJ7K4Y5myAPrCYns5G/kcD32I2jz09PFsNpFZrnAjXbxuE
K+OiB7gStlssGr/MnjlpdTTR6gOgla68AoFJjpJG2FH4YrLxT6Ag90vn7xBB639dXvofvFfovA9k
pNRnlnjHcDGOWtZrXkskqKR5haDr7ZWAn0q+dTVUelDADDQfUpHNFcuAzYkWlOZZdaJ18VX/z/+R
/plEyssfcy8UlxxPKtdxKkR7jfB3g5CAVDGO4qoEzfB04zGD3iTmxXQWOgzlKiEkIfHm2US/W+az
hoEjhNVEIr2FksLKC7kKbTYxRf3sdF2z0EbV9x890zvBEflzHSauq9RSyBUjJBMEL6wCO5oFYZAQ
b7ePxVNYr4HY2q71MrLKA+OL9F0iQ1vIBtSCRZaMWAxqCpBT0W7Xo46fcC5TjIULSgPkcUlOzOCt
gU8ANrGyUAnlCcLXV6ESlAQLrB43jcajnEqShXTiPLBFeza5gf7dDo4V1Id2kJU84ZtB+jh7WvSm
eWC4g68iVmyp1J0PfcwhjQZezzzUc8Zbmghtzt4PfU7v2Ezp/zJwiXtEPtgGgv18kSG5IQflOhih
UHIojFs/mMckdl6fP3tzbr/jHjy8LIe7UTwvSAeuU9U8sCbzzsb35oO/ALgs7sSybPbGm7A793mw
aVvnd3Pa3lTuXT77e0VQew+Aipt9fZiZg5HnagWFLG0ir3QCHw9TkAvrdCtL39AB6Nv36PXE3XKK
zJeXAMfqC8RbcUTeut8wHUVlVtZ6OElGdr6ngGI/H0z99tglQ95KlAAuNoTO3+V71gq8T+fTspQ2
BeLxJdTXuYtlAA1dSJM9SzFwudVyBr7egGWdGax82FSs9sfkfz2QVwV6viMaY/lpgOpWsDyEwg1X
19Eycm9uo/mmRs9nW7xSYMMT4FczlenZxE3yof5OdE6catK29irTFL8cY5+rI+DxCG9ac/UxmTye
0bPJNj9JUeur0feLzym7m3FhahxixmIubbvJynIjUBny/jfa4PtbdRibfbPf1DKtcxwgMBtizFhh
TzBCVJujz6h238yanxh5VBVVAhtCuVDgVsiNOVl6A8VvI8b92C1YknVtUfu1K/KaoNG9YHHjA4b6
poBv3ru3WzAT02v0yIZGuE3cAW9Zon6CpsmHW7bitMt/CDWguQWxHwKmVZckCoElnBvJVNh6Zv5x
FPzzll5Rb+QMtEQXt3eSkpur96TEo4pLtY20sgIRoS3BH2QfwQVeQtKYbIURCUoAB/1vGcGNXWcj
BDiwkulBlqEk9YIcIhYe5Ro+DMYs2bQMADsxtiw4JfmJ0y2zvLefEul8nufUHs5mp5YpRgnKHba2
wzUKaMpzuBrAnAZBTnzI5hKD+dA0JfwAinCJ4XXaNGSVk9GebcuCW/E5xbg6KU3Cl0LhXH3etno5
7Fl+ZQBD0zTeo6dYctq23JzFeBW05evF2N5wewWsG9NhByxqOJVRAQwcXuGnsCirH8vlm2l4paav
bHSSgE4m1OBiypSSxQvM9hGoKM3ByvD6RCbbgQXWs92vTKHTDPa1Mh8Wwom36ugHuZFjFZ+W7r58
4OSUqiw/FNYPEcTCikfLg5meeICUPTV1l8kCPUoN6IAiajMnU144VGCS/9kBQSUqBLzmxaZmn88f
+pyfb1EpIz1owD1NmwTzr4mN1hDyyMnYoO7ina0lK6qqQmQebDzOyn5xRYSLE9Y5HjGFBAT35kGh
K1IoWDFstYbPAt48feMefK8/NTYoPj0Eu9NFHQhlytNxNpY0a9y++iZ8YmgWbBjvHX4dOGz/5+Fc
Wu1YMpNsT3gDSkOTBnVtDdHsYXdqxi0kO/AfN/9XllCkh7VcR8iQripzbfNMBUN3rElgaPxmpZ+K
ea76tJzO0YiDuA2+UEC18i12uZrWE7V4ldXwyWG1+wRUaSuTv9dKA4Q2lUNXni+b747XUR/WPqki
IILimQiDpAKHHAAIUeS4oA8Yh90AST/Deu+18Z7o/Lea1KVPmaVg7DtLRy1ODF90wLkOCpwLYAHS
MgaNih4JmzhybKdftbivZ+U9pUOQavl8ADiRnvP+g2d6OPgp5omvjZ/jdDbjBeMmNCR83FYoWls2
U49p55yCK55ClBXMmM9ImvSxQFVoA8TJ5MGnTixlGWvujFQLPxTg0tWCwXtm2IvrXw8/Qpd23sHj
z9wfRqi9vO5ZiLZXsnTkOhhZbL4lLiybY9vj6p0BDW4FiHLPoFfENlmf/20gDbSwHkfcZuXdpDdU
vfET5QMAecEgs4tbqVizhnvmJGir8kuERGYfwnk/kduQBn9QxwteLfL8qlUCqo8LjSurm60mCX25
GDr3VB23G0vhuYR0AHQaqEe0Fi8LQgRSqIZRmG2+B+DrjDvzxlZ08NZ73WvsLC0y0fwg9w9kVnqe
g/WZBE7Azq/2j3m32cp83MENV3/9KbShsLogn1DdNpRJSrB5HiFmcEXyOy7DlGMpb5jTTaFZsm/h
7Mi6aapIq+PCPipBEEDGWJg27/DBH4cmRBnhYZk3Hko4QoI75M8kItteIrsqOYrhGYqWVilsHB/f
BSBrqqOZLkznCmHlnZ4QBe6r1KixuAjX3PeH8zBt7xvC6uDDWm7uDPeA88/JaJf2mqmz5SIvkG/d
Ry9m1gEYnx5JrK6RAwusHuA59qQDr+jXQWHM+alrGrUl+uFPb7Kak9372MJMPKv0/t5pR/SkYFiz
q9lD2Cb6kP+XLCThxfgErP8FHlx2c8qD36QLK5sEUOUAHOmOYK7bNIs+mLHnZmPqkikZ0ieeBEhs
lWJV0bOtzGYmpgyw1K9qRR/8TqRoFhC8wf3zx+H44vf4m2BbRgZrolb/9GnPDaeRzjtwCKZMbcG3
ZWz1D2Elc5pzbDxQ1F6iXr2GYjPL6JJk02/yzZ14FMSNpQScQBwcWcOYBeLVag12SVJJUAnOFE4n
T1Sr2glaZKJlO9f6K+dKJVr4EwLp39S7gbKGmMmJPhBT42tQkLbzNR5Zj0sQdtpZ5qyAyd2z0Cnt
Vpna35Hs8CSj6mOPu0X7HMIWMeJaZubi18x8qODCKmWvy6/2kQ00LzkTtrqk+pjqe8TTPcENyFHA
KKNTAaPUTSXDjGscIcXex/bodUsOoXsx/ZujQYWStlMi9jaK357HBAOQ/L2jPcUggl7iEEHm8P/o
mfZwsuIwDj2pmYHgejIGhFWz/vEOz4OoY/9la3sURiNJFAm2SGwqPXwwELBN05AW6IMW5HvpLqq8
9ITdEdb5wS7XhEhKCq5cupnTC733PSxZwdkGsjHDNauWv1QqOqM8S6u/8TGtmzbu9AYQ0cMJxnHB
XsBFsABMCo5eRug04mGPdKjP8HLI7suTziDwpij98IsWXY4Sp18npc1/2t6MUB6DLd1vDfQNZsph
Q3KsHzOSEXGGbP12nbyqPc3hF8U7TwnjlRjQwwhwOHTve2eRDyvFdXdHz49z8fK0CQNJ7NmWIV2R
7CScpYSa7mHej0Fm3kaGuiDSR99d1GUugu1QrYX8Fvikl2wZcuyJPlMBTBo8ezcPimL7Mu6iB8Kv
zkGazG8riVfypftmy2vKRXyhZNIbuygXt+2fCBG4aSz2Tp033ol5NT7BaoSMPQYIkdVKb0wFAZci
Fxfng3gZT78fpHcxsEc/LHxGpayMTqH2adKq0nQYM8ZYyCiTr/ubvkfZEXfhHmZIWrXKQIdmv4Cg
cZftO/I9XeS9/J2miKlJ491bPwZU5oXP6Es3zRq1SXkp2nB2agHB/9jwLff014kTDZVkZhDMS/N/
jzhV0uoCe50sWuF9fuPXq4OhwSeUJl06yf8KO23u0YvaBMW8fWf3ao78XblaygXHVu03H4zPoyZN
2xPG2X8mp597Sj1claQBTgkWaeqdpr4MCD/6T+vB5wH9mOUGKcNqTcr4Ys1a8l/9nkRYAnKF2RAF
K6FfXSK4XCiYDcPZcdNfsZlRUplW9lDO0NVwL7PQSQs/6wReowliJx4TVPjxBQBO6GUkA3IB5AbX
BckpujS+2b6/36QBGaOYorrIeCLStDsFopaDM2eqnfD9PEHYFKeM+ulFSXkuca4W+tm+AFkD3JxI
pUKiNtB26/+7wuLiaBuSFqbWkwTckGF2m/ZDOguFhNVK3kfP1w4pjBagucanTGbUT2v6IpGgXLPE
84+bsgPGqGRqnjVYZAUwsDB1wEL+rsFDjCfjM2u3H6HDnlxeBncuP8AznZPnT6I+9237zGUKtHdN
0yuDEpQ5F4OrNqvDM93zW/jUvNXY0e4upAwTCppmB6TmVW38QUw8nP6KJjY1xnmCuXfhjxxXS2JC
l747gkWqupbAgG6kHkoCoME7DdLtEIYDBkCwFPX7RxvfYPwChc+TEE6s9aWocSFeU6qI6RNEWMQd
9QsF2COfQm8kNgCTTtBygOzMdRToXcmKrX0h2bdBxZNRSHF+GuZJfca8QcQK7rtPUHZGS/FfTwsl
tUmnFhLRBDQqxGI8lpehnO1jVwCNR7nFfYG9vE0FUdvd+HRQvYybpnkGx0jhmOobcxYwDhn8Zx4i
mGs928TFCTMQJdShwBxFn/0LRfnljKpoimN87rYStXOsCfFbalz6GQhKMx4IbfjaMml2SQqHocWr
QtDozvnOuyLDa+lRhQkCNEe9E9X9w38Zuu23j6Tpk8FXE3ZL0ALTtHgsVER+wQrcN+R40rQ7yXUo
IQd1zyjqDvDSqgBegt9WEtBCphnX0m0sfCAor1bIAfQVz2VYDn+ejMvja49K0YK2Yn+n5PS4yUzD
dUEAUk451U6kTp+/bQDQ9tOIuZc2bHujoIKI/ujs6mvVSijCqMYzBuy3AVSFA+u4niplSVhH27iJ
3wux9YFjiO1LgTnT1Ln1WmZaJYydNEGb9iKFlSj/UW/5nCCFqnRp28zHXtcpmgM5h8hL/wKrno9H
5Ve+tGLxY1iDrMTLKzAuwjfkngesoE1TqMCRH7QYW9yLouAhm/ebSW5d9tJ91sFxQH21o+3NbATy
Py66PCcm2knQp62d6+U6KQmzlovT7HK0kW1M1BBbyrYs6yQqOqCfyWXezAnBZyyiZDGuKJRoU0Ev
TeHzvy85s9f4v678TUdQMtzP/876/kQqJ4GhfhWqL57DOzoxwLWbpf/Qf5c9J+MvM9p95u75+0n+
qLdXX5xa+ZD1R6lzFJaZ9OhC0nwL7xRMh7L0Sq9RcvFdIypvfaNdky1CnwZ8H8XOaWI3mBxVusXf
k0s/DiMzsinKQbTKEzwPrfA6hdalUMiDVQI8m5/novRrhfHp7ehZLFmSdSYFe0t+AaUgQ9ogQdaI
fJ97XlCoYH4OU6JcjchmuafI+IZJBBdWx1bb5B/BfS6oZXuagUEkyu3+c7bwzqnKxsrmtk04XgP6
1V/PrlkzrWYB/oqCdP6kiWjAyID5QEithjfWDAIFdQ5YXeIcGWHDTQnoD1I4xhg9kMWzo9SFLhZ5
ewK+Ahk5exMm0TQecoErdG4EkRZuJ+tXWOVFSeWdJxwqAAia8EpyZwwDie+8GXg0TtcA06gf5fQ2
Kg9mDvv/fp3lfXK+Jl/l3giHN1AJSf73K/SHf8YW0YrMOvnbdwZMADWaPW0mPLi36Y7xGCTMAdAW
2+LaoJVIyEjRbs8cVC+dYBrmtzCJqBAoJeesH9mWO7mPHtlDXWVtBIUEBtW6EuVt6gknTLkrHVkp
hUNr/WJ8pR8qcCmP9xBWdCuqXLAWu5PwbwC3ulTeYTW8C+BGtada2S5T1mQIbXr/9XjNyG2Qd9ry
1oNFFlfyGX+wsUUULLSo0jGVQXV7oLViAYoMP1RtwB9f0xMggLZzyi1S2S2McbjY9faWgXCCgriL
ThuZXmAHaFPc/BAwoewAxQwLXhadyTAUzCm3ju+X3MlpDp05ZKQn3vq2ma3uGe0sTG4KcOuYtsgD
wEMQ1JI/x/fa0bDrYJ+y/J0DCJp3WOMaP+NXSHgDN5VxMvqJAi8zIUuBirPPhFPQYMPduzPSrOBv
MCilWUcfFsfGjKHYlACnTl0ifnP6K/rpgqmmgikgvvZkXsYzTUe9aLzWpHNvd6T/ucibEDba3IdS
GF1aN0DkWAeeCq4nfPbIJRSANYDRwt9rJJJqfP3ngrYkenzXVKeBfamTiIpDUGcHHvlTo5wg2yEv
fZVZKzCBP8eQJlfEi7e1sTKiPadAW+jFKa1F2SUFgIz+AiVcHnyZmSsAL6Js4yZS3gxkPbxaonFt
UB0N2eSIgDfBevXsq+rMQKEsEzjg0B2nz0uI7wdtJoUu9r5JtC3XHjh1bNeiPrI3mditU9LHYuo7
qpqZMVWLcIgqOymb5xYM7VRCv1faY4QKf7Mibyu6wnJXlOMxFE6OuhTkesay46tfaDEGr16PSovg
aKJrLPfXPG6usPUQX9cGb3DRE9+FMJbLTj07b1IKrd+QiM6EOw06Hpxq73p8pY/WgfV7ZSpgHter
mVvuReDp6oLZG+kYD4cPLy+gICPhCDn0hNHQt+59Uka3GZ+iSJuEN4/K+wQQQmiPTWiSuYN6EfMM
DE8Oth3iGYIMl7qXZxmRUBdBjRjqCLeISp++xiiA/UPbjEkXtSfa1fU+FegA6IJgxM/FMt5Ej0L3
zzTVomHCkKYBkDNma18M12tV1tJNbZcLpC81DXbdau7GVwUveSLM2+QBiQc79DcGUMFPthlZ55ZP
g2dkvVJ9VqWJmquoAKWSsfFyJZ61I1AEePNStqfTbrh/8/gOId9guFFOQBc+cZzncxdyxGp+Gf9k
L3c+qWxC/nS10+mz+vFzOZcXHtuws/5Ien69Wgd4odfx/pAlUD942fFiRyRIg18MU/kj0D8Tz4H/
ZBP1w9yUmSifDSEZFdqai5mOhl0D6PUJLd8wXSOqdEHRhwHi7tLONdFAKrsPS58f8Uz2JJ/m7tpJ
dhtGNe253ksk3o1tEWjng5I/gc2mVlGuXXi/tYMhkRZXJl5fEGcGEPYFddDAN80g13vBIkpvFHXD
7ZQ+AhPya4t9GXcI0nc2XboXUc3H2o4VwxIQTcy+NtC6cdU226sQC8yCloxVOLvD5NdU/dsG4AT6
x2/1WH2k2cR7v9quXxVxMBe39jzcHGPlQDRwC0zbRWWFqd2VVoqZDk+E/3cstYZUv7c71vBSSDJ3
jirmrLQfCQoa2klLH9e8Q8pVDQbR2/fiKB8/W/OuKeBjyGZRLh3726vrF7KWvSKA19IlKsH6z85q
HT6xpYqBSoTi9TqIWAAEkoYXNfuio0I4IqH1V0pZ+qZExB3Yoqwb0quolWp+sjjBNq6rs3JoKUJv
R5MTxPlykB2a3kCyg1BDXoq7HnFkKUMTnmexM8+mJfViC40KamKUzYLC4lQNcWzBbAs/AFaFgH8H
UawTdJsV7wxgv8hjYtafOxUCXBa2YF9yXgQpfVcfZESXzwpi/l5xQuCjbwFhBw6l6dc9DzneFqGR
UC/3QkI8socGoU1jC5JDlSU2MXsOKMY4tT06RErKdUj8C6Pi1SJvluMT3fkxCcQ5X+IEVWuHfusv
6iFkrkQCTFVpclJJzRSP+O4KGKdT6Dh9Ty/GUT4B5TIztUZiXPVY/3tmwFl+mehVTLQcFZhmIitj
2CGgBwG9uTyv0S9PYsT+yxv49oDgvKjnEZSCNolHUbMYVXoyUDN/Qjbl6JTj3g/VzNtlKzk6bNJg
/DepmbJBPzfQsTWq28YRM9HMyCd/LQ0frkgkNp3/QB6ORiaNXAXbYoY9e6IPPnhodIerwYlFLC1s
UAZCNPKL8XfnIJ4uifDFfqHWCIt7zCie+9MzaM4Suj8Oa+T4xlfS6t8bxFOiWQfN4eMx+rdmAY51
cta2ArpoQCE5sG530ntCJ1ROYIoK0Aj5MmFiqqPU6WTmw1L9gW0zm1GUFnQ4MzBwFJcpBHvoleyL
M56cfqcM8j+MAM6WFtRjVwfsqerJPQ5tG1quHwPU1MBkoGmQAILR3xnwd5TJZf2nXm00Uuub7B6x
KD2PvVW60zqKYGlQUMkqq7SCPvZu1NEpZDOHcvTgmLUNbQwu7qQcaGh1a3QAifLLkosFr5OrFt66
Y58gqULX3/td53ulQzk3gLx8SpRdNzFOVhujsPs7VI4fnF8MclEUiE993WjbCdiezMkEYiL9c+ef
SRtMPE7JO9jZLDHdr/tLnPMlraw5J/jKy8dBgBGLfXmm5mbtxC5yOLYipSvSQybk1UbqJ2bTFSji
f/ehYYse8mL6L034hLelM3GXbwofCO8bGBRTkogt/dXSj/fTglYK/d5C+mdBqAifyVlUr7EWI10u
IVpkGHa1QroqM/bBTfd75DKdTKdm5hbW3QcD1NelN2oGxFDtk6lLf0SJMBKRvVXN94mGvYNptkGY
FILwyuPHBe/wixvmeOmVDWo13NYdvwjJhLp4+tZIqYLIC5vFQv4pKVYEKhyWMHhCyD2zTzjr9iHA
KI2erQYslPa9RH23bMOfQxP2AYyVJqSIyHuRWMwWKvEL6rD2BZWJmDg6qHke7q9Dgt4sUrHsCCU4
L8iMgsRlS912ocz5F5/UbNCbGnB8YI9Jlj6TweF1aAeNiHwxKwgslWiZDIklmVDK5L55GXVfma8u
lex2xQ3Pw4WVz7bTRUym+yKVtfiIWi6Qgrv15mp+w7LTnHSIcMg07e5pFc0kP+kWSD2gT4N07mOL
0BZubYrE1lP7D0pcjpuerCzsSvqAyrEVZw2NWjGTKRW6YCmGAzUjreFXCme4f6xHigGc7xrMo63+
dGQgdtjx6aZTT75A2SvUQDht//VIFK7nGJ23az2kJoLmz7Xp34jurTjG/EnFFYfFvcHE7h7ReW17
eDH9PgbXhf7kP7a29o4yfav3FcWsh59O71H45kQSWsZYa6GY1ygJS2snvX9ZM3wLs9v+5vvwkyTo
D56alpwYc1lPeEDQhQhWgxSlImwo2vbK0l+UbTV9kNIp3VMi9tgMWATLJzW0BLRvl2mOsRPVa/OE
t9SfJQsP5QQhCMS+1gcxj9mFnbD7xobJKtF4YcPyJa7W0d+ummY0iNZ1vcrdeaaTg+rMH1U7IVuS
Uabo+c1wrvQVaXfbKgkAxnpGk9mttjRfCr0vJRYfxU0b3zkAdydctQKFVebhZv1Fr1LGsb/D/Iln
/P1YUqqJS0tYIkdTw5KqWOKUELDSFPC4hlg1RzakoL/Y9PZ4uGCSOQ/Uj5WMdP+U69pLgI101yCA
zdYOWgW4T9oUMWICDXShXcXuD6HxML3NlG8G0K143NBJrNzHghrqbPdy3cE/oCJQb6F0F0LV+MkF
RfCAkaQH0Oc0jXe1KYtAj8Axcbum09Cn3IlGIy/PT1boOqYAPMtykF50QdFiUi4YwS5DsSclmss7
qwa4lNNKWvzStkvRhjc/9DOyR43qhfmuZFNKNmM6L7zr0c2Xw09OOjbv2zdmy1/s7b7Q0MM5DB+w
20WxNVIrWPvuRWwFwNNRCCPh3xZhAxUVJOAWMDP9v2FIOrm8R7GyZkqph/aezuq1L6D3f3k4ka5L
Em7WfXtuE0VHDLAa7/JbBkj6DVPInP+t8/5T26ZD9T+mBTxRyLiuEsmw2+GJYgQZMSVQu7zk3sTG
zcY1KNydxN65fcKYCumN+ced4XatTBx71rcxr0m1koqfC+q1gAqGD5BdF/eFwMHoNl73WjbfbSGN
YXyDCp6R2WV5uiGOj2lDtFdUNYB3mQxC3WtMqM9WfQrdmZ/OuV63OqVYne5y2Ls7ljjSxtOgKcGq
zyCXFtzqrfv8vxEjwJr9w5/snIc4PLwhU0o4y+uOCCJFE6D/epoDHjOLZ88eZraqADLoF4Vv6hSD
VYa49Lg6+AcZrQzQyhKs/iYv+wDxZAFTjs6vw1nwTbmLCL1z45lJCAiSGheMS8BB8U1Ql8cMSHru
IcZbzf8klzyfxv4peMRSBNRHXUlnjYMvHRBc20HwXZPStvWkfEHNiUUi1wmoZTFB3ajnYXMF7y7c
k8ZQj9Kind5hIZHtnwSSmuQvvVMlNTlJNR468SsQvfqzlH8qx2GU4JP0DgxAg+Nt+5rTxuMIk9dq
kBeaGlna1PzPNvhw9RM2VXV5Bvq0jDcG0v9Fl4f9r04Vt8cAJBPTB3cNvUJGyts6Hbg2bstRUTjw
OnBLtCccRe5S2EaYQIfVA2I8xLvM6R5mGSmqSl5cCwlaPxLF4rXc17eJnPJWPLCYVPQMUNRiadLg
sGFtJ6fPbvtdHFbU3UUZ6RooBVUUx+8bwfTJh9UWpQ47jh7izzD5RSdLT7Irm4W50pXeCEzgGxSv
Jnn3LWEH9Xq+/GbtZveMeD38Ce3EFqjWjx865QmdU7FbWbn246HdprD6eDoEpKN8G+66bHjEOvup
r+aB+rnP8Lefwhen2DUCcIRACUeTZ4FItSBeaesN7L8NbSxf3Qnnd7HlCdY1TIGzXf3me7+8aCj4
wl38L59fMZM9jxSMvIRnUx6AtSZyvoCEgZJQf0IdoTHwxDuKTnSaco6tpsts2HyYdKiqcA4258WJ
yQ3xr0oHaqWAhToNGm9ybPam99hm9zaFIVhFw+AlaOMGsaaIXX+oxpd5WwxZZ2lkYVgwjFUDvvjJ
Ikz7r36TTjOb+YK0MKLtUUQGg9WxHYJFrJhU1ZH4mm44HTRzdhbXu6ZOSfNLm9/0nLY+EPGFM59b
C0giHWMjr67SyKZ2M9fCD9EqVNXMrxDc0RkvaBphotgIU/6uz85+/NOgFuOSJJFyiEx71EeM3iW9
fchPo8V62tbqNZuymvpH7Zsc5M+pJtY5ag9KPXfnXd0gknLwTCzgws9RjFIL64lXoVJ9EIvplXG5
r6hDtPAcf9u29vCMNfh2Jv8PqTBOPcctTehuThu/PFdeyVofzJra3aGZGMpU854dswnGVX19jePu
wIRRdJoppCGn63qFjoDalcReM+Y7T5IkyWfn+UCXNcpRZczZ4pFkyNA1+RibNam8TX6PE+/MNMk0
W/3Cc/Dpey7R37xAALYq8XGCg0vVK8WVQanGwvBhKJoWnRZ3ld8HDieC0d8xsflRbfpyCuv8iZlA
ZQnvUr1tno82wTXwcqmByRvVgmkjbu6EVTPb6Ms5xEcLlNwTE4ZdFoYUTAcU2gw9UJj5+ZeDfcej
99Rup3iSYZJkDvPbZkfRFZgedMf+qxQLiYHTS0KAd/RON701vUtpM6zxARCVOihyb+UtDY/Efhz4
PU+t2WWY9ota2iSWQz4WyX6ZgK16gkI/4hI4GHKKYNHMx/L9DObEoksmBT4FJzOSSzHvf7I51QlT
QiDCHnWoXVrgDSsWxk363SE27/Zs/qITby/kykLkZr4JP1XbuiSu1UM7TxIZo8rK57dhHyC2Ywzb
Gv9Lln0UjzEZZfwW5fCuqyzdv3XbD9zJuPSPGpTksfFLlxwS/TnJKQmkfeaPPayMrqTg2hJUdGB1
/SeN27ysEj28vkdIQ225KW+cJYsdg/MUTpTRAT+cascITwefndtjam7raMrx8NmSPkqZ51Baz/8Q
OMtMbv1PxwiIF7sK+R7oCR0ltqRqEaEBwzuXkPIdzuCMHQik2YWa7SsdhOSrxctUbpLXn5qFiYOO
VIDf6p1VI/Xv0o4l87vxmJBR4HzHHhSYiSna9YZTmUNWRPGLUtlSRehLxL/g6BPVmscQwSkg43qp
FIxUlqj7KwjNe5KAvpSQwn17nsoqGb1p2dj1kLQeU4cvtmyJ+LFaAgqklIoec7i2BRNsqhw1pvgK
rCaRpnaJUhmNKem6u8q+KgNK4AfxLYdiiaJs6n+7Gsay1Mx/GVYJ3jEhH5qs+lu4HHeaH+4OJszv
zl73ZGPVLXrS0I7mObWV+BTquQmiVm7Fyxw4vD9Hkty2Ixi33XSsnccfNtXsxWDUQqAVGNK5dxMZ
hbQ5Bzv0kNJ9YTkn+tY0/ariIe6Kv2t/0+YdIdndsSU539eIg8VywE4WzXsCw00Y5g53IfwLxTwD
oAxpoqAqBlt1qNEfpfd+2Wjc6BVuss0GPoYnW4cy5TrNmN1FX5ZW4Ftda9lEsQLUCa+gqANyJnrN
xyp1VhEcHAIlz6D0K7MzK8jUnoJg7QC7U+YwAQsEiU+tAIyNGTx3KHv2lprd1aIGNl1mHmPucWJz
woVuuqIoqBcuqUUve5EEAQOTfItkAKQ4RPs+GW9Mgdn9p+KC2QbA2r/TGlfyunL5yUZ3R5G8VGw9
Vdvu7Kk5ykO5QRYNGxwuKSkrlF6qBKDIZOAG3eXtTHnmQXyRDftOziNT7BFlGUXdSEBRidzvUZNJ
wFjJwoOsaqN4Cxy+4rpB8+6vauqh+peBjaZ8yWsTXSnGZIFLZ5SVhV3KQGMD++w6AqSv2x5r8Z1l
DyBikJ4RSfmP/S0W3cXPZswnv1YQzij7u4FBJb3KBiDfOTdEviB/KFYl4ieG1xWFB7Tv0RcC7sHn
rDVXaqB4fiqI4CUNBB5wk/5tZ021lBJKB0unEx7tapVcyGbLVZohOI0Yt/BWUTG/QnIuq46V2SHC
RfQkBC5rr23vEdcuuTOGBws9QN+/6J8jEZytVWSlQgtXz108dadzqHTLHdQ4MaX7ImOLWG9uys0o
7iUZTLhcv3MackO3PvFm+sLPoyaOEm7N1OIwocLE+rAtasPW9OJ7DCNnGgxxX58mXEfqizVdSLnl
XKt3BZUblejvoGzN3efhkzd01WNLQ48/HKX9TcJ+fuOArVq7zctL4h/O/mwk4bfUNaeGZrUgcDu9
EOcDMHouBW1opWgbXvZnbRRc8uXZGpR4X/MvUjOkWzNtWUa9tJAhlSQBUKLWgT09Sp2RljkAuqOI
Pk8UMPOH3KAqal1CyfGUOxOlXIrfMsUYg5sMkMDqNARoqIFkMNX6kkspx7D/kZkujuVnELYuZSK1
346/3fmnrNkVhNXHvuJ8DoLlih2xj7Sh8Uh6sFRxZrlhdEhvVMhjxN7TvUOTshkZ7ypUXIVv6r5F
jF8zZ/dVWUq/E9SHsQpumTBH+YfhaOEmEFx4QCurKc7n4yBlqF6KPeLfVbGB0ZZl2AkOOjahZfTf
qBzdkXoFIgIQMpq9/eWH54ZN1DJL+OBZg30g3fi95Kg88A+6f46uB4PD+QlsEUNuG2bLC6U6aJbR
y80ddHCqSwNj2vQumhddbgv+VQ1b6d2OuOWMHOuvP0F9uOVioxa6+7o/6osR7yqD2OxBdXpwwkB2
aLly9afC88Z8eD4ucs8JaiAb2Bj3GpTqhBbKguEEhWDzTS06iWEJziOHtEegWefa/z8/s4kA7oZx
x7CunV5FTvOcG1mfabhIR3foVvwk5/zlxJIYsbzfPc99bJ76Solbri0RSzOYMhwb0lq/zisnY4nY
YrFk9Ms0suyLwWfRjp8wHsKFYirqlQSBE+37y1GaPouswRVrtXnVXO9NGVVqieSOcR5W46GlOAix
fxMlUmFzOhysyogZ7Fhs0C8emaGhwGAnVQTkcKIaB9mNaZDq16K2FNpzLJ+WMYjQmfAyF9iY4By/
N3BJ8ZQLmYXdas8ESCfB67DMLKRzqV6sjqGhmFVH5KiNR8SnJbZkxi8McueX20WOFB9dWp9O2rrG
Oslzop5YBdbDy266/3DjU8v41rsjC9c2DlL7Bvt6hLnZkn5yJdPVsCwRGON82pUNTCNm4/nk77/Q
rFkJ7HoQ0iwEoEeF+abBqmrIbEBu5+RfmqxqpMaAcInK2HWELUSfJFWnde15/UkdyswH9nEwjuW6
ZzBnS04PuS31EjT8FTEUz7Makhi56Li4wPkz2GLeh+Bh3UL9IlolAEOqypowg3/XOx+WzkaWav1k
D3vrB8jcfgcBEGDj4GT07crJakrc6FR3dOnEEC9yEhQ/yZ24vNi8KULFBYin3AIqy9TdIicpCnKG
WyO6agxaA15+HiHvxlnEKcNJtld6qJeBOKj/9JPKIQf2RyhfyE1nkHfGp2MttrXRI3AZyOOqxiJ7
dE9FyPEhGZw4dZYNdAOaBvoYcE6DaZHHS1U3/h04nG3iq4G7PxPMWICfybVq/HLVJ4W8K+dV9WEx
eABD+iO87aJGq9uE8mh979SzgXqrA17hgEr4lYBlecNHL45bMJxUX2VkuPEAggv6yuEjH3byCemr
Ef17JRHd8KJAN30gzh/3rMyStuck95tJuOOZ8QMONysEx+BOVn7LIMREbulghdIfjub53BOGGjf4
TOG85peniN1D4L71cdQ2JoUSkr4gwYJwaO+vlL9ZR8i3EqHeQCuesVovmyx7iQ/hTL/nMNKFM4TK
L7mhwOdp0RaseybIuYoJ0/Rd43gl9ZGRrKtECeqlYcsVhjSrqXjDNkyarOrWdVBRC7Zy8ebVVuTV
zqXmGjmwiefU44g6tZ3sZx6yaClhcWfrc/QIZxHw/KT5wLn6raHerN1SZ7yVclg1ONFd2qtXVGaZ
bGTPWKusDaabuS/rh/zw8yszzDyTvCDYxPBtej2eiT30Li0/qtLDQ367le56JNkTbvJVsLIvEcf/
qxXyJnQKteoghU6M00QIDhMonKNZHh3fGQ2yhVjyJ1CwJH2MhHc1woQ0GZ3hqs902mBxqhOssP91
wOmEMq3k19K7TzVxzFyWDSf8SPqnEzVXwc+2LqiGFGW18A1Uab9atgmMjFs7wxEHPzxaVXnoFS8D
75IQAeLo/a1kS78dkinnjh661fDS0QeE6Bblrg9/y/3PRVGMMJkhzXJMhddGw2WIWA6qZxQh5Ty0
Wk8osUnWwAnAxoQaJ/aTuv4dxUZQjTadRaPUH+2z4/8gaFxBqWWSla/cz0/fb1+GL5LrxazWuRMz
9JCs8lxWlgmssttC3T6O1IyNMm7var8gWPHbIpLlRnSlWXzizaaCMlhHARavjANb3FTUw3MJLB+r
0g79ynf658hBOMsKoHhaHBVehhzmiwa0tbcfzAmWrbEDQ5U8DPsFjpO46EGA0lbt2pJNne3oYEgb
j3VHnSJ22LHiwj1waJDwYFRyzZbmZ6cGRxPhr8VOFRI9gPTKR3FldELjamjX9MWMY13zq5HXCpf3
gdd3biXUvyxkQZjxb3B157vPGUrYHQCc47uVDC7CUU02d42YEGjTJ7iTdz8DlO8bkWDE2ftEKRy6
dVPpiuZvmoDScTgcoxsogyzLTRSaosL/F05h/7MbDuCm3/vl1sxP+c/3L4AIdcnAyP7bwlRspvzr
GhFnBnDbxSmcgV959sRZAkkyt0L0N6N2FTXvVa/9QMkjiC8nP/fXe0iqv97iTDw1ljmRjZwkzT+D
r/E6Qc4rFnJ2O1lVE5MXAxX+V//dMABSUHTJBzvF93UEw6+EkacVh2NskowmucOdLzgd9gDJKAEf
y9hmkVJTGpCvKvX/OOaEMXtRKm0T5qpSTEsud5K9w9bp66RZXbJo+FZJaUVvJgoTgpOII8jgiB7z
YWaZqgLHQ4nNdPIn4BmF7Efn17vC0r7r/ms+/NdxW76e9p8ZXPNVyBVCShehj+6vl9LNYUs99OMP
5i+mk5anb9LgcSgfw6EO46PWhypcn6yehMre7uQBsgUt8W1nhbdVdvsSHKnbIEiF+Agmx4q8pva4
T4NK9Mnqw904xe1WSN2ildK62cRxrUI231PVSgQ5WqglBi718jWkktAAB8rzPRd3s//fDjz138Ol
fNKB+/hReOZAEd5gGWp/ODDGZ7QEiJIWhTl5REh53tBBbkK1uHy+tq6uTS/g5lFqAbOoCY0b2HIw
Q07NjyjG10GalyTgUUv/HeXLl8whpZHCK6sOyrq+UVxa7ogoM5AkfKUV+uMuyxD1k+JE6VZroDrt
0ajSYt27VSsM+JYL3ehg9vE3qRH6ZhHZGG6cOgz76J/2RE0d8MCMF2ISkWeCbTTuQ8M1zLt0986r
e8u1H3HWItYmLDDDfLLrsYoq7r84Pklw1gQxCjcMwBccs0K1AFvQINLrOEgCzkjRBaTmRnB8fy+6
xkORsmLWw82ZFsbQm0siUOxghU07qg8DO3A0b8f3O0F4jkHFvbP3+el24XeroLrY0FjVMco7LVbq
F5LRoHQ5F7UqRc0a1O94rgUygJR45P8eUterfCt5iY4EISVSDFKGfAIwHTmTHPd+FGV6v7BLxRI7
fYfVlO0f9BDCcVJfCSJxrXCJiV1JdOo6fQcj58TD2c6iVAQaZG7tSBLJqgjqVw7mNxDaXYYGB33H
aSef43wOcbMIvNNs7b8//koOH5tF8JVUZI02V1GjSmfIjalzBy+V257XjOMy1l2Wa06F+qpHYwLX
h9aEywci+w7X9x0UYHfoTXiH/JvgT84C7viomEXLEImWEe+F5LCEgbmMPPtURjWR0pY7NkwtQjst
nLKS0nR8Nb7GsyoQi81Inkc/U/q7ji/ID/BX9PFq5J8NSwa2ZdWoPndTM4hXvdLh2yukOfLj2Edy
p24PDHSgop+tPM7G6HGtoYbbpVuwgAa6hdEYOfhCaR8+Pgwf0TxbuNlPfnunnmwMKDaAhBUyHa/2
PSbTPyYgQCp6esZiUYvUKm8mCroYMZoQRdyHu60v38kjEdZWHZbxaBYKmgfvjgZ1iC5tO5HveKOV
PRCyGAWrT/bg/p01RXmZUk/F/8VqyoIgwWudaP4z4B80bzJyKxPlHSdfl6zx09aPqzOPSjQxnJTH
JqmiTgo3jI5Darz6bDehv0KxaD8gINaZbeAO6Zn+ALBw8p3NxoObQPfYZ6CfnwqWPaxCfXkuLg2c
h381qiajlYkffpi9BkrV4j+7cDwB55viUY60X5CAO/2hmYOdrD+GEUD6rjQovm/kk+8tlb0p0clc
sUm+FEPO8D0SuUfbsE4bBvIyj1Fhp3K0rEh9paFeDf1M/AO/We7+qa/WtJgOLEy13TyBJu3Jt8Ik
mgULcgPRgoDmBM7HRVHDMrqcy33QLfHPIpBn5F/+dcpiu3FDPv3N4csqNU7RCcHU4g9Tjby63TEN
eYNYvw6c7UVMGf4BVLm4Szb6cRCZBdVyEg6lNlWKcdtJvMzPFkGR1ZCEwd/bObJPZ54KIiIPxapr
4qafBRUh8eghpvVj0l33us3Z3R5ECkIveclo9S++MkmPv89NUOz3V8zd13HLUu+9rkmB+CC5mrNV
gAgsNiFnL/35jUxLsF07eu0GbazTvyV67dS2tcA/GgIqz9ZP2vGY30vzOJ1HSAA0wbnFjogk61E6
/oqK7Eb2lxM8CRysUxRMsP5MfamrKFZqgA1KeofGZBM/05s8sBNqfg1OytCfY95Hr/t5+nwoJiJm
lflLBQcGd8Cclu0J7l0mZ0TRLglAm3qmzGn/dbO52D0puCkSuFjG3RpKcGseB8My/uCVpGc2NsU8
wXu8LF7Xykzv4AdyRMZwvLBHc7t9Z5JwGaA+tZ1vh/m1iF/4S2xxURIyds4p4/ULPhoJYB2jiq1X
xkOeWIRV8DklpwqVX0larlNfkZcGj+vXKF2evSjh+KLq8rY7wvMgxC4Q45VLyhXque5w7jXNgpS2
0iehtynL1DyM0ZJU5+rCYXVRpfK2F6xccd439lkCiR3CNol3B65f2cfHq/ie2t7nRifZRdfvRNmE
ZtbPu+BKfRBQLqyUNgyhNe6ITvTVcTmwUrf6jKqt2h9c97Oens+F4CnGFNlj2n1LRMrHRGWx7Acf
wtGIxpCWt/seD4kvPV8uMP8Vb77MjMuinbH0uI3GJJb9Zq25q3LJw6cbUmzh/OYZuzueuJTAhS3A
BOZPLejBXJfu+ilUAVUfchjBpOOdSG8PsWRd6MVMxEeA7Z+XQPF2CfbPJITxqNimMnzeKLAYMyfs
pQjEZka/UQ823nGFzJCwLJ/9+ej/a4CmMH/2TWM9egTPrILr0Lu7dQ0mxztxE8Z02z/q8ehAH8Un
13uZ5CFY1uYGOIl9UG9sgoPLhkeoX/wY7VWRr64gAuoiqeVDoNNVTJ22sp7Hb45Ru4eRdd76iB7T
eY2QrldNU9wFCxHobx01r4Su2Gx4J9iZohl0Kd40Cqac2NkU4AoDErD3X8gBsMbNix4LxWd+4ucO
/4zMeEM3dw7BdDJXrcH2DqyddR9WjYX1ipn00SjQJooCBf9bITElTtfad6efBLPwJjujt7qJgZmE
7+Y7VKkemv85qkh66O8SaM+LDmmwe2K6UcOFMNe7oAxE4obgH7mlYYhXQVIWGJMVO38XmFIQ0gRT
ijSihpQZ04Y8C/tNSvJYNsrwO0nAEFVaNYA273qD8bh5a0q8GlGBPYUB97Zde/HLWvqS05dekx3H
XxTQSGZw2uWHqci2z1GuvPxUS9VxBO3cEwxQ3HsvyKaJMXhol0XJvHpAdWGcylPe8b6zj9lOCASc
HjxpzQsDR/k3yGj0J2gC30qXvVPwX6dv0gesoH1bCeQhPpF9X2/6uJIAghQFJcHRVz7Kwu5Kw6IZ
4hRkluMs2CnEeCaPLyMb5Ffc4sgq6yh7iV32yaf9OIjWaeCfhAMJDQUc+oHnWj3WcTVE+quXvBPN
aP+mFrVqUcvugGW8xnJ3BkdCmsMAg+njn1GYiCUmqq5Zi1Ham5UOZ1vOHTVz/aFUEBjWPgxKo0OM
oQecZcG0raM1OkyXS6jXypVFA9xT7GoksdELTxFHqOQ3jreyGwi2HQGUxE7QeinXfwf+vS3xMsVN
vrVGAppMXf0Dj1RL1GK3Eh+mTgz0s7TDvGqPZ1ZdEx18+7l1FqnolBYLwm0l2rl++UJn2fC69BBu
7tHn5UF2C87mIk2KZ71YF7m+Rc85PN6hTnKnRz22uFFB/RgCgCwtUWw1AwHGwMFZ6lfkudLhOt0w
NxbGHj3I6jFQRi88E5FivO4cBoxnU/zn8e3qZNePgHXlHEP9E+qO0szkDossCWnUNIsPdGF8Rezr
BAUsOyAWiM7jeVboC00wJ9WQrUKtZvbAYySWVokaNmcUrfxQJEWOzDEYZQsLOhHrwMdCCpIzZ3EM
vbAL4etQYFjSmAxAAKP/EtTYSLoemv6H4IChrjNecnI9MfHXmWpu2gHMYdo3ni3GZkQMjzQcut3H
ZeolVaAV3qYW34dkVDQ3dlkiuy+iN1EctBHFJngE8XgSvlfwtp7Wf0eZMrBp6mK2dC4X3T9KkxTr
36hx8QpBOlbni02m3Z5eqxtI9vqYUOK5EnP4563oIUxKiMcB/NWv8nPaPv7qX120QkVv7xYJnmo+
5GXnhs4ePkjajOnwAwPNTk90vDBgxUp47GwfLTKBkrz1noL5AaJAqjzWuBZKrCBOOEIGrkXrmZN0
W/H+Z5OEACZC65qGFIMPgTD+mv2Q1Djn1ZLSG+dq3oRtLL7yNzUc2erUDh+YrF+oOvcqIMzMTQjW
6kzgOb3FNMKQlfIsdlYZZ+Lz5/J28qLgYm59Vf0BouJ5wk8yT9lZMYBxOElTEG+2m8oiX8cUC+xF
q/v9ng5jsuTr+67Ig34v9v2WQer28qcFCxgNqF3UyBi7dafIfOGTD8CXkeRLdpczb3d4I1euCHtz
ztnWZLph/Wvc3tSt97ZapcLCD7VfOOHoLzks0lDy5uLDcQPmqUTESN3ZzeK91UA3pfonZ4M+5T0q
Vsr8Y/KOdlC9K22sTeWVYfVPUPghLvp/lGhVoSNCZstsSA64MQKWZvn+p8Ldckx0nRJh+Jq3R3gF
OM1xmyyKbqe66i+lHWGWl5rkjmYfRV96XqxIO12JZgPieNSlwlbKaQPweCAJduvuidUEd+f2eVk1
cT/Z6x+Ocshz5w4fp9/iBy0LN+as6oAlMpoBIBT4QLcUK6W8huXAfBW+vUPEWvBEQddjqJkWPze4
BJYKf0yNf/cPzE8HgqB6obe3cAEuStjw61LN++JN90haHFB31IPMMYpyDttebDzd7mYpuNIeYv6L
FO1riEfhcCkDg1YYnQ/vuS3RA2jgLp93ALQE2WBrixzyMPaQaFthH3Euoaspvd2oADGIC/wUBpI1
SQwzPo1YCaR9r58AdlMESdCRGRCV1bwqJEDpTuPeH6Rm8w+Ai4G15gjeppd3EqZUiRdszcItQBHZ
o6NjiSj3Vv129WVVWZif3HLjg1PGQs2ABu2C3UEPh0g/oAV4zTs4p/5xdzn/8u7KkTp5iqNM0PYT
KrSGPyZYo/soUXs3ae72i2cw0yp1KTdhABpbk1Rcp2qjtzekG4kRmM1J8H/qJ0+s4KIpMB/N//1X
BTspmwv8fDUFdVlBvtHXF58Lsf9hKlej6ubvWxlS7Mt9ljRwAYVhLL62ZFvshu8NBuWMo+trbNWk
XtoEVTmL/WOEtSLfNbzcLGgNQ+b5RocusYD7BYvTW9j0OeLOvq2ZZ9wSRgfIT4uwjaPCNwtwzoIn
Q7IopBcW+vsq+xSlVpN28qpZPSh0+8+w9fAvDVZZDPLs/TwVNZZhK5z6+tQRx9XikEqcXQV7mcEk
vLAJBaSfjjCkN1eEvyOgaPGRHUE74lXyozOKzKE2wAYEbbVf6vQNKekNkRtbjJIc6nVhccWh+tEi
V4bzNZupCElLoNrY+I5JUPuOhb+fccIESuhB2l+5/Fr3+E98d/HzshT2xqftuSa1Sf92Lul5n0Rw
rqJZUR/ZWFGwvejxeAiNDhnRgTqUclC+PGogn++tbBcZtTlLYF/Gxk5zJUMVOIHoD/M+kRPOaw8d
NxGU34Oaf7SbZy4RoUZYqU98LkDXSXyLWxGj+LAhDU9ocEwFezWP97XObaOicxOLrb0qLwRugh18
ueaXslO2nFmnialaK+R+qw5wyUx90iLtNQfMroiaCj2CslqFcNcSx5K8d8q+GZoGeulbXq2XKhF0
xpIHTosvI9WVRqwqNrILVet+VMFiAWrjc50kEGmEgJYMYBiPC1hQJ+EW27Rcmaf4qOW7wl5slwE8
jEFRw78J9Uk2FR2Kcq5iBFtEow/kcU+NJUJ2LTRIvSFC1rdK2Qbn3gKZ4aYXgXWp4dIH31TFp9bN
nCT4sFPV5kzBtzG5+RSLGp3giI9JDz8C/frjRQY2N+iJ4LaieZKHdZ14v44okM4lS4QZAL7PHVIq
8zxdeSSu1pEvFH3ZAV0nE6Z3E1E1W86xG0WbMboRUDjIACloMx6eAS7S+haewV/g+gOwSuzqD0SB
wtyRSBa32/vdB+5WHTftXFspMueveydOsc54iUhaBfpCJOHyDaPLXIQzymwbqaMHbwQSCWuRDObe
rRQdV4KIp6Qh4DoLDI5OqwFnFXKWdP/Hc572p0eXdWXK07go1IV8S1rRD2fY2vE50rtYj3rYnJy9
alqq1uklVA8mfUi7hun7aJlqUUWZk9KOe2MH6s/UsmnHWQHEPkdZd3udDEEEmGvFkti6aLGgfICN
LYK0Z1ufhc5H8u0oIviho6HoWEPvC4IKL0I++qXP60rXBLFUYTMu/W3XySwwbaUOEhD4fRb/Z9z8
vvJmAQuaK3emGj+u40Shb31hIKOpIRNip+hdV3OXLUvjQwZXvsGLJSNSwO8+f6lJIGUqsmR9bUL5
ZHo4wFvRYyIO8xi9pX3+BeWy6QEFwRVH5L6GCKUAcHFPEwWGUyMFYKsqTloa0YEa+Y+307Bm84G5
qGK47EtWwAgWIYl3DBOVf7qLLQYZAtrHgffVAv4u5rHyuFGCbpQ0oGf5jsfbb/3y0fP0srcySAVB
ggg+4BGZOJQ01vmDbXoofl6nvw3MKA22vrZDDGTMnK/Nf6At4hSTpYQOMn2+V4auwk5FrTCDvNzq
qhbUJiFa++iNzN+102j8GRUoayUcOK/f0DVtkdxwX2nQ/a1QhAQEXA1jsCFYjoQ31ODPyT2Hi2Z+
4nyJHuMmrgeIbMVPzON5JxeXNyYEaFv9pp3gR/Xgeg7tLexTiZEKC1Ri5RaddBsG2UovJFtiM10M
IFACUS5JXztL394ns9A85O86RzDTwPNJpPgbShNE7brFf2/NufuaLD+VAfG2b/NyDAvTPMS/I6dg
XnW7ii0VO2ApHcvPi+5BiXlc4GVIrMDKvMk5NRg0guaAQxJEN4gly/N4Zr5ADggTVOe2yExlr0gc
2AX2nXylOUtFXDCZ59jRLD0Ed8Hop3+pNuhI9ttjVIj10TpQUozZ7/dongjxQQCEItiJDSA5XP1X
pUvfYUu1mmoCCwwjK+NKPfDdp+mPWRcNJY17umXe/OHzrJOVzAUZodYj1J4t7lh+vH7a1Flm/tPm
qAPWkkSx/qX6gNEPI+ZxW/EHsmvskdm5pr0jGb+BOspccN6An9lh8cRtpcu3k7RRgDwDsAm/Zj2v
Uc2p0xYsX3hE7EVM+P5Qh3x2xBau9y/yDG+Za/Py1DLLOJyl7PeOFlmjGW+9cGdtSpsXW2qc0XcT
WpzfKGnaUjgrZd/EPOPHgMti1AkHlDUINqFan1OkoV7sVweft/g32t2NrhRNPlT3+IZvYW9lOm/m
cXBMj9duKGaSKd6NZHABnMlkRjG+LaQlgjAKbd1PKPNERuGnd/R0m098p6f4fMzESJji7nijTmxz
IRu8WKGArGpwKMfmk2SGJB6r+iwGUUHjYWltRCY4shlHeEDwSpjwenVqbtXn7XDL0yEw6JzqJF0K
5ZrULaMx1wm7CcFubNtccKKHxCJtUTlV/gJL1BPydf9yhcXSZ+J5fcK13Q2vvIG/X4iqJuzY2ZDs
TsYhVlFLWRya8v68C1J6H11OJSukjr2M2JUyNeGrPnFfFksocemw8Ur3EpZx0DiE1nZYqTsH+wch
jLn0q6oTZNBqdchCLrUnmiAIhZ4yU48qlZoiNfGfxYCoPKd4R8/e5tsNSA9XkFAUeMdq5gMU23re
tXXM1t+ndk0xMnnTSoW+Uw2MiwkTEYVBGJQZAJ+F+2LM16Aqz4JU6o4gzjgdTtWjXNqVbjboX7D0
rCk/4+35aVxF9oXG364Hfu8WrEFjo8iOCeAsJpQI+oXAa33fBOWjJvFR1pYlwlpyJ5iA5hTK7GKb
HFqJh25K8UuJLygD37ctX6dcY/5OPJV0NkbPmPbHCju5NZG5DcJ2LKcQwY5sZY9PDcomHLftB/za
PBY1DtehP7KCeF8xwCjMPtsGIXzB4NdlhiRVSg0yMevgtnI/AVFD7PBSGCg7BC2D77g5e3SG/bGR
3bngxkMdXkLgQSz1lXoXSrT3gqiksUMxI4yU4lN0voypG4ZMt8fPx27HGfKhMzvifyBIdaAIkrh8
p/HR0Ovag51NE5SmI/v8ad7JpujAu7lTaVXFwMmSkcHhXccKo3Ud3QLGLJq+MfAcqjvbe+NQJZvY
3w9fkqwSY7ki9QLdImNOEEad6eDXkiiWrVEz5m/BWtiKoAFCCgXkdHI6Mnj3O0jBCGRvtO2iZXrv
PVrhrn78bOPGHC9u8umK9VzjQWT4VuDXwaKw4yqkFolGUwC2Q8VbQyW6Xeg8K7S+ilZ8JQTO1y5k
OYF5Xa9/veitjMfnf7SlfFa1kfpCdZ3xg2KyGDHKnYP16T8xQOqTY6QqiSzh6b1vwaGz622t5xnR
tAvqwr09j6XatM3s7WCRoS5auw+YjymzdhOgCZkwaqe8OQo5WyuqldvgUXy0k9XjMX3QgG9+dgNY
sLjaos8qku1Xkq1nB/rQ8cobLq6VvyCWAtpiypZuOhJUrcr07PK8nk4yNneZTOd7igOC+Q9UOc+N
jXl7urIUPlxMdYuSsKlszeWVpNcYRhygQ8e3ENsxSneNbhQ4DB98nYkBt571K6e+x7MHojjiphEj
HiMQGEBye4VOa4PcIOvp9727y1NPb4MwGz93QW6EFptOwzW3uGUKW7VDivHtgf3zcQo7gQNVXTO6
bR/QuU04iGPDtP2YPfddWkc94soWHW/bFZugzxr0Dly50zH7bJvXFmEX1b73MPUK3b+YhhapElkm
ehoOWLmxxpdyPcemfryEelHj5GEgVoWUksk68JJkuydrg3hrSzN711kjHFi6o7PKwdMpwHjaN2H3
HXsWlZTheH57HIteQglPD/BxFN1uzZF6qPOpDjUDigPOoChcrPKmZnOKr1TH1XG5cjJ1LNsewfSC
NN5M6PJL4ncOOYP0LawXTfyLp0qe+NWHJSHMy5pjzF/teO9Rya4hWHRBZGvrJyK2aT/AFFYjLyZU
PknAS3xxpxgi9Ihqa2CbxQ5uLxAwpgZfUDdB4fQuFYQYjmOJ9fOegjMUAR/dV93YW6vvYgo6mp5h
ocyUWqGtEQOISpiIM54Aw4Tv/+m7smibg88LXshPaIJ4dU5aY0BuCGslZcT2UfHKSkFK70Xoo7ji
Sl8VcVFIIz+xMVyNLJVm82AV/DJd7G910VNzPae+6W6CoF6SZ8Pnoq/8kWA7Gh0B9CrZF7hSDFGp
ttLhBlTCNVFpMUGwZNeke8wHrdSBVSg61W9jhck34NRj+2vdhW5oxrkcXdCSFVZMoHxBGk1fbSaD
2TRqQcxidoo+zw/qeGEo1KomCDCVj0Q0wqPWb2r52R202cgaud9G5Rp5lTk9OoMIUNAxPkHKYs8j
vTk64QZVkyNhtVR7hyaZ4wYk0iuZu2Fv0GN4oDln+MO2YalQKgrRe0A1TNPAF47+9cXQIurcVBBs
kS6Zg79jExSoyxJiRiHbHqQP4VJ63uOBs/OXbk7A8rAQIRTpdQzIIPJtJQ3Jv/b2gOu2WkicdMoI
dyHYpcTxe/4XE+toafgx2s/NBQA2GidNEh821uBxVtheNTLOCP5sMIh9d2+c/JQ3NTvYdS8FWnCk
8ZSU2wTn7hbPNbl3u3/gukAONhzfXrY8QvnC3p2W4CHBesoOqkarTnW4Y7VaoknolVMvYDeVpz3a
nrKOMWcDIZm+mJNEtTbxxwAoUmMslNrT/Yp5k1vhnQBN1KZSCgbAOI66xwq+tibUlMTS/MgeU5qg
lg+tqu5AiOhJgVZWxCvjz3NXX+EglxRNNl5rTRD5rtR/lqso2RXUEMdOls5JHJpVv5csYmawPmIN
mI2F6iArH+Kqf14EZ0zcyHY7fGNFVHweN2JYCmPQaSsypV/arx3lK/rYNPaKYXaFjo5lQnH9vV1p
+GWEzvhWA2vU6GkQgsQjZknZCgGXeqzxiDop4gSR/CVZtfT8SAMtFs38NOzUzJy/OIafzkh43gm6
ot3i7lZHKEgKUHwHwEjZeNVEdbwBp08/NC8VZS/fSPzjFLXCYvMxRXr+n1xs/0VlxbzcZtqvD215
upxZ6lfgohBmnHC5tj90C5WCZ0s3yI+ZA2+j43pxP/TlUpOjlaLlEcR3963OsE4p7Nr5k6xUzmAD
hv+Nb/b1epnQ8Vou00TuzJEDOKeHW4nZcmeRkRd3l0HHcmfIKUVMDAKC8gaTN1hmudfYYJzye4e3
QDkHIAPs37KKKByoBGnjvjf/M8fuBPjIIftYZfs83xb0RTc5TytZU0d6HsUkfaSQAKMrHjMEwECd
Y/YkVFm4QctUAYuthRHrZdXpo58wwC0bitylpXyyCIYZGYW7bJVN1Ms1D2sD573ipYdTR9tNSSEh
FoxYuV+4nzK7pDSsV4oJSDqTQOm05bf2ns4cxWe+7FqPRwRWeqZdhLRLJejqAX0I+n9Zl/9Z9tXo
EvNyum49+1XcBrlfGL6ylscPP2FlS3FDPvkilz7GnI4uwtc4gaRJBzjE3fR0rcqi9KlLkZF57ELP
231/shUcD+t5gBYndp7nvHqtTG23ljRgGSOYffQevtb+0oQjv0OSuZkCT9qTsnckxS6UjiA7QExh
x98t1hBK5iTKjdTs3cLyzpfemsl0O0e4NXNTPYsAI6Ish6WsQbkFVi7XQokdKmECm5Qhy8lPa9fn
VffOYFjY/bCghPZv56X00SUuZx+XY6pR2YfDn2hXMjmSNS4tIQYuuwn26CJRhF9E9rU+KXjJFUJ8
qCE6HJwIHNkiCt5jY8S+pIQaA+zHa2nZGlnlCS2XSgvXtptC2CDIPoWqjPN4QQlsU+FIOq1GT+qP
8z8CWJC2/pDLd0t8LRyK0EKKQGVPVAZmqzVMF/vUH7rCxhrgrG8alg4nY/7zM5ab4jHj2dFvBcSA
f55cdJi37yGY4EWLCI6ZvexJi93QnAafFRId8h2uEZhPY2hKvy+uxffbkXOIJmLGaRPBVN7R/FZM
4yiqCi8AocbsOA7n2eymBZiofRRRejVU8pY2HhTaXKxF5FtOIm4ulnuT8RYevq/rqQqlVgfs0QDQ
Ll8oiSWGyKlXr+1IBMRTKlOV2nPNCdcOpp8W4bav5IeKcbDulw7WqJbJHoHgfdNFf5zc/WLcBN2P
TFfW0gNJv9kAfgSs3Nd2QK1FCWNcl3UHscV9eOXnsx4DKVwiLj4XKc3soJTfOyQHro3AhINN6ip1
13BLAOlv8pEN+x8DSJU4NcKGoKD9/rW5wD/QJevvEXHRrkahlGsX8fjjtCifxNLyYG+P+Q/NG8pu
QeUvs9juf4soXt0NWUvAdx9l8MlPDTk2HXk7vsGH4bdLOEUkToPeW87YdANYMrfIqHOzufXrq/68
nPPxu25EDoc8XScxFfQbQ13tnrECZLy1F1zZ9rD2a/ll0wr2zxKd6SCn0mhgxDP9adDt3l1KPXfi
SHp2Ik8OMwT86+G8zVVIUeXy2cMoy8raVIjIa30QngR/xzJuY+bbnQSI8CA6NCLhZp6L7ZrDfyvh
bpDkAeqAH3eMgE05wiuUa3mQdkwbaQcEbkkiRYUGD0lEdWhhc/0rQ7F74FZRRCQKRGBHlLko37jL
v46yi7Wo4jXOp+vJCZ+XgQOV2jp9rN3fSIgS7o1Ca506PCrJFFbZ3IsU+IjPwQzj8ETQL1WsxTDN
mat4MOAwbFD087A3MDKAyBfKeWkpn5t0q+JiwbbMBkjFY0YqMx/T9+NvhwkgUk9vgiPbJRZI1nop
s0LYBgATs34T2Fo0k04UajEc34bdzP+UZJnYw0EglEfuX/mPnWngMTyjH9VFXkKY1yIY3NAfuYPc
sqxk6Rszd7wmnl1EzxJTFtE0gvAXRJSmi27UUIpO4T2ccQw5XogKc4Z+w/CJl9g0Q+XBFOQgSIJh
vCQUPK/NXZFAaXahpkFB0ZxvzmNP2wzA//Y0uT/U10hjpB1EKVjKsuu60K9ic1i00uOKi7g6r58F
TBF8PmYPXYGuzOEURE/F3g9abkxr0QW5QxGZAPm8zaiPz4SqbnTHnokoIl3PpWbxScQG8lzBjfCY
3yLJ0eXl3L1YCmiONAgIXPFseZ9Fy2vfscJaSd0tPYhF0MmH/pajvg7pIrt81wL5wodAuiOiTgd+
SDL0hFUAt1pSKm6nhA9gpOulB6iN5xbkAvsZdpVwcR4w22k7HDhiuTIJLHhmHxz0EXKk9O4CIK8o
n5JnyZleDvOJli0qEzCS++kw9gBPJkeac0IuGXJEJpIUciVnWLFIWsZOwHh25yTxs7GfkjNPPV2p
rixFnvGBjE2UVYXeKuZXQ3q+JgoQfrlEtxg+YnUzsVZJzakmOBXzAIK/bE3obxUSF7rtkPs98N5G
FlXpa0vglEGdt4UP52ItZgzjJPs2A2xvYBBXPHZqG9szcR9dO2zDttWcpuJPR/Oy0mfMM050lzc7
tsS9H3exAClCT7q91NHlnLAdyaKnedSqXx9+YtticcLzeSU+LfWtdBpaRuqddBssFwhxD1Hfe1Hi
a31DRajE0jjzQ8Q3gPVublyYkonHGuUZiORIt2sx5ESVIKi2fXNCBQxhSPM01ct9SMhTKYm2+aKy
ET4Q+0BkXHYOOzV/tlVMHRwlnGywloLFHPumOQFs0PlaVtVmkqShK2nt8l2xgzyMbK0Uc464Dx4k
VpsLqkYBDwglD2CSGB42e1InYKRjPtDrTe22WF7Z60D8EUDIcsa5K5MmK49XtSqHUFPuSiBUM+R3
gTe5kkjbfonrpTIcL1LE8qcqosveeIs9L49Shmhx5wYkpw2BUMLqcbUf7wWPYfXcPoyqs+yvpuD2
+gEr9RJeddjKc7hFD/8NSQz+HT8gNAThMdSQ6kPcbUCZmV4fCS5pZuRtwRwpjKdHJVp98+MocT8X
sSCqM0Khyk31WcIvXbfN3GjGbmLOlIdkTP4/rme9BhAstQVB/11stIeMU4U37Vzg9qtMC4mK+19o
/4pkjzMTBRaPWSpIAyjxP8NHMboCP2NwQewBQEflErnav9W2WvELfvaqguf6sMdzNdcivmpmh4J6
6uNvfKO+9o8IXOKAyvkHtCjCSKDe8YcUKoAmxt4VHWMV3o3x6JCEQP9jPa8+bvT5uqrjq0PC0HX4
6Sj+Xwdk94WRBMxOfu6uidHbmbNDupZ7zzC3WZQctyRyRTAN9zUDkAlp+jowhbUksHQW26mcC9eL
h3UsXxNmgVNoBRJjWvKIM7/QXQoB7c5clLOQNGHR70sA3oBtsRaVoBR61xwfzhVIPGMCvGFOPBlc
NBeBJFXhMeyrI85f8+RnaplpXZU5yV5QiQgqWwRIsYrNZDTQGfkoJi7oDU0W8Y6lkh5NYTbfTLav
67APaCFbQ+6ZxPlnizTchIijBFpx/8UmqkzwMNGhNrms1gvk2EQAnmIREwbsc+3davLYOW6u8gNX
XOKnyRSyJBc2Zf9Jo4oHv2xxN8BsCFHXspN3rD2tol67o+vk8K7PEXc8VULfE6UbztmDbQMtqGKe
yflx+sq+d4L0Z5HtNh2c5znvctKQky79UmYJ7fDg0/p1JtZx0jMqaXLvO/bz6KOdaphxFqsuM2MQ
mGy4UMpKiKHi3yflQzJKn3FSKUYsblvlsHikIpM70VEjTcj86QX8yXebmiVPZg76ja0rFaAbvKtq
k1LyzPyE8T6ufk8eLofZ6qd06tFMSFcCR50ToYL5Dc+gI9Jh9+JxqtkO5jcLsxZ23Zr1Am6OwpPH
iFI+60EdGdj3XLf2O2ExNahQ/OACdld0E+mHwMZkkIzfKK4oxJa8hSZwH0sjRKcSV5zYVzRSdz45
fZH/Cbr1GSvWellJ6C0LjjJLURZq2/yKT22JfUFcoD0e6o4CmLVFRi2AhxAAcdbQNhzzyxFnvj8a
e9UgRk3sH4sxEjwqlgtV6HAwsiuSF3z82DdS1uvAE0HC4tXVKp0rzp7B3D6Z2ChTOuTBcsdykExM
ZwR+U+qj7GFGmKmFNd6mfE274408Q70ZpS6eW2tfJzJIo4xvRHclqKkrMl6NlpvPd97zOdgtibcg
zpAAAjUYzD47YTqBs2or4tCbNwu0DlYTzlpVA4nKgQLSkSUR3IZ0hjvf6bzagHFotlkjI1GNZc/O
FdFD3Fgg0p2pfMIarAwZlOCefq8VvqrzMfuL4RdzeKdUunPWU/X7oUeXWvXM1YyBGjTrkRDexj1A
cV8pK7cm6ldJhRi2aNp2LuD82R4zau/6Wj2G7t9kc7760q5VPNXZBkyfQB0ctTc7JXVs2erIElXb
tGrf7WnWctTz+yO5hr5MtrV0MassycCzUjWQKW/i1xyOx4GTFrHCg7FMJ/PxRa5Yz4rDUgWeRCqC
r6h2MOSN1MMfGFhiNpwxG61fvxZRPKDelCWro+O9vuLACSrXTkC5YrXERlu1Oq2DG6lLs/Cjh0VW
j7EP3sOYZR+L9ucgzBN4ssfC9pmAIzWGwpORbSaaWTQYjCf0JaCR6hkxN7VyueBpdnEa8o/LwjJL
7kcW/UxO2FJ7kZs1StKXLcnyOAPms7gaxp16t4QJ9SAEYO5YQExugjJwD8wFAMUQi4TFzMv6P4zI
yqUM/25txwFkIh+hVBK9SPl/DEjQ2Hy6wNa4twtbGFZtkaqcOrccLg8mrDFbhylRvNwpzSKM/GAZ
rfac+AdOd5SiJEEDSxfmJPR4R9pVETtHY6HE9LaJBGvBuA8VPOCp1SEebHJrTKp9kvqR+TMhMvbx
AC8vaFRLPAWX1D7ULJixEsUoETS72+/i2BdnOg8n1LCqUDtVL1Rr8OR2LvcRIRDx/qkmXs8iRW4x
idWCs33yD4dwneQUJVRUWhb2JXyYsd6R5GqtG4qcFJfOijcAD0mBDhPPRle1jX+fbuWABnJKU0wY
li6cSKB75UK6vn5N8Ug95kTtmAIdFWMCKjiotN+UbHxS+ouOveAHEiIaSzLyMCE7W5EMXJYkXmEs
9qUmP73NuHRw5KocifLlTVzQf+Tz0RYjxGaIKN8ndz68D7ig5Dv358N6wEvF4RENYlhCgaGxaUBV
GLGHEGYM3r7sa+i5Nlo8pdJ3GnEnWGN1zjUK4KR68UWXj/n3IWfcowzveVW+J1Q7O/Z2PPh7y216
t49rr785LFsgHg82ux8XbKHgS0LZk7esEENzgpto81GT6/r6bTvF60GQlJn640WtTWUBhSdsu/rU
/icgkMWom0Oidpt5+vN7Z1sJMLvtmGEANNTVUnuWfj6gJhJ0DTKzjy9ZkJ77HRNiehsbeKKDfBh8
UW5l4pB8JfZN/QCGXB6+Gv+E46lQrefQU2lIqQz/6S5MjufDhls0qsec6h+zI11VZX3m49d305h3
O2y6nF1M8sL/YJ3oVPnwGS5jY4xsFie5PQaIbGujXAcNzP8F5KpLS5Ufgf/qTO2YUtPvTU77CxPN
Ai+OK5PDYh7jTX8+7DJBo4tYLC/ARIh0UNXDJlYMu+I+Pk0OVIblhpwF5NI2MfTZ4MpFpeFVhSzl
oWLIXHQFvGffHkMfR0reXH3ywrT9XsEfth53kPfy/QodjzElk3eEM535oRXd1uzh3jYmXmYjRzPK
RQQKsghM4/ayhtBrmV5iW1vkDy42hXnshppThSjKAqercgdqaAxfT31dPVqM3nuXPDPTLrnHNSdd
PQOr+S9KM012dP3FbctaxcnPwlo2CImggiFQcHjZrkCAlj8cQSAwzGEeffBJwQ/BYjhe3m6Ij4L4
Tlq6qvvQKu62p6anPfXCvcO2BTKSChLMIugzZ2c504UPdc8tLnvR+WLje3WHB8BuK1KCrMCdimxu
YrBLVbOHVO74HqO6AYpU6NBAeX5Zxcc7boeK4LOZfZmcP7bjzEtZyut7fDHNvfC9IvXXrMHMX0qV
hWx93RPTIvwtd7YGW8MArAZtWomrB4HJ5iqL8EmIen7cu/TOCG+Vbvp1pdO+2PGmgRzxgUE0Lw3r
Q6/A8AQ4z2U0Okutf01D4fiXdbSOFuiGCuRpRQ/9BEpIHUfdvpQG6njcjrE8twsDOO1EPjDweARN
/0B74buzeznMb4rsQhGwkCcPjwmtdMtzv17iXnmTpT13S0Lk7PI2XemOSzJLbCIhGLNtlwvDryCM
c/7g8Rjy41QwXE4oaM+R9xqT9d3nB02qpNjn7qP40PgELUCgGj8u7Ggn/Wn6yTxZhKlnKYrkrQnF
nuWKF6cU9BlXOyRjWZ4LIUXrCfmxKpLmIIBGPoe53vDgfu4HJ+2MyZMEt0Nhr9eRLlbkjm+8IRy8
TUWyRmeICgGB66sIrYdEO4vZtuAkxOtd5hRmXSQzKudafQNxoNM6BMbHvTXCqfA40JlzisRfabeI
4rP8kPIb2tqzYRAcMRh+X2/5h4luyV7isSzMCuXRnrGznPzgCP9/jeTOitXHxt4536vYhHV02Ryp
I4rhVctdo3rm6nFYhYcTJ0FqsTx6XyTVeg9c1TU0F7xSAPXCBBbExTFeaYEf98bKiWKOD2ZI58e2
9YEfRlf8qGYHnfuDUS8ipRFRQOu/Md33ZdoKqikIsikCrQ/H6aregfHyn70rXfa6mtvEyMk/iJiZ
GHIrAIwJ2X1iNvXRi20XeJ4X0ilL+/hMecHHGYh0KUL9oTYepcDkKQzjOndsCpeGksjozSur+x+k
SLUfpRFIuTkidiYsb2pJ7zR3DjQ9EU17ojIczrJoe9wX7GroopgjL7uRYPXeEnSaV73gjEaYHcQP
M7o0tUBRDwpCDx6/7jlPgcAT1A0gu/8kJbHavTVVO3lBn+0Npn6gqHhAq8ehQHxufi3TE7yVcBEQ
Ee3AhKyDu1cC1sTTRtUDoYOYfctxRtzfwV2pbUEL+72eWLaja1eaFFfNSmou/ZLSy6lTKoKYbGZk
kD8wXNkizy5+MvHSnABcZ79EemhZGbaEvBatcwsQSpsKm06JVycKHm2YNDdZ57UcS+pKMI6En949
6A+b4kbJGyuDqCjTgIol9fyyb3sLV6YKUeBqS1aM/8M1CSlK58siRehs3L3fiSt7Ii+eDeTlF4eN
hG9FIsh4y9B0gohHMZ3LxV3mPIS3JxFhHYkrmmjd3Fk7oHYpohkg6PNQofnusEjySCUXql7W5xsm
0TLrV7gC66kAAnyuxrOBwNzDJbqnxFCqllXUWoc5ofMxQFOzTtOObcjK4VAC/5Oiol2rY96GUmSH
bu7z/yRx4GKJjrF79Yg9HOFgBeM0DKKHtBoSZ42esDA8AULrZbKQ4TaL9R2u7FHiD/o+5IZ/qMUi
XWHruRB0Z7Ni+b6orXwbdQQD+8Ezt6W68i2acpii8/OaRPMFNYelZFtUV240b2bpoDPM4cj6QvpL
Fc/8bdFA9Vjccd1Rdo16+QEnf8E/0W2n/wFGdKs/1B+sURGmmSFAnA5dRl1f6XRRBMyTxGlwz89y
eSe6Zsx8SQpzLCr4IiCfD9yw8TqvwJj6xsTc9+K3fBLoZLtvFIuPmKjx/93cT9FJSVWDzk7CAfqt
7niJ9jUDaDt2vlkEXjbqXjHHdzHYjGVHIX+7KXe3dhOh46dlh0ATa+g1zZ6J6/SUNty35XEoh24Q
VGKhkTzajotSo6jBy3kQKqKyELLk+7ZzvZAiooKP2YsBSOCVEEhxPoJqzSfNhcYDTIPAPbGqoip1
w7tutJBtprMz58Wyl47b5RxsU04CDNjXjSjXMzzjaYDAVnuqsASyy6PTHumLXmqXZUmSejIhG1sG
VAo1vwRUSiDL/5w/jpT5T5DpYZ6OrdUzn/lLdh4+PZqIvBEhbGp2JaUknIMm9ytvW7leDYZdV6RG
1ELTaDcU4JbNH6quwSy4JwTCj0a3BRbio3FcLXDfOAS7Pmcg4YaFYKLSn57vS0CcUZTtreLL0WSN
GYiWwoel9s6ul/+g5DW4HFxo8pMeuhDrAmi4xizopkq2/EW5MQ61rEHJS6AduvJ7oKSEXdwVFXa6
I48li7dXaP0kDHLSgT0tw+TgmGTNrlhexUjUd22UT+jUQwLkm5uzoBm+uLm1BnNSDqMbn6KCS/U5
sgSgCOQ8eIIFoV8Pu0ugza4gqw5XmE3qaNJqlGHBtAg/IwHLkWLJq+n48RRIhx6i3+Wto4ew/iNv
jxbKAv0wratbbY6VwalOyN0tOx33ijAXeff9ohIeSYC0z+ZtUwCfM17kmiXkhnf0m05kjpH45gPF
xQwuwE5PxJQZowAF4+Ll56KWQCOj1VN8/i8CtRnZLnS2SZgWZl185y7md7WSEllgAM5QNuSXAAqL
iY3BXOSYlA3igClxMA6zm6CKrftKdg8WbboyEBM63/8EqLH0HpC7NxSaw4IlTjm6a9ca6q0JmUv6
38kppDIb0lmEaEUEB9a1G+dMKTHJgfbyrrNDB4gthyfuHg3UpDFtRA1dZ98NRjfVJdTN7f5/FK2L
Z1p1PqAeF4MQQekgvDRfav/64G1325cwaHBRO9hjYe+yRYQZ2c/pREh+h/SEMXu3vhlV2aDaeON4
MP/ndMH9yV+sOvK1d8C+cPISo3EhBd6gLAyx85ZoKy1AZqKnMRqsGTMHRqx2pgms1boT4DIO6T7q
0XvdwEkfZt6aMHuC2B5smH6Xyw4ZQkbPIra/TAyE6KachF7mt1YjdSypZWi3hxnzwizbbAeQwgv4
7dV/60ltVKH+LaLM8TSC5edLihx5JV2m9g3YYdn6CkiGTidl6nGB1sEqHri2pfH+NSdo7yg2wpdL
IYUdiv/Kr6TFl/u94pyL6C9gcQBjWM5lx8MoFhjjPMIeWhBrR1u1Qj9/fI6/30KwuGY2lPWVCZS2
9JxSorkktgwgoGJTAG6SNlIZ+ppVJ2YkraZHi7TO3COz3XpDiypqrTVjJO6V5YVn58oQqwciT9uX
D44ywz1MH74thcBRkMhV/J+TDR8YBTLrPt2gPJw0IBfsHhtjIPPFNiHhIOqxEvlPS3ZVaa2nCLbg
8oEfaEK1eaPirgBPl8Mb4BYmJ0efodEW00yFaCUrK162ZiHhssUccQBfjB7ahmpt4RU2IVMqDUtj
3dkSE1IWniN+Y0TlbLShPjP682OfMo3cUHMCkd4Ozbzbo92+0WWsdDx+doSihH5gzWSM8zlPMqCu
6geY1RoRUNR8xCsyku2piaUJ2lmmSNmcW7JZQT2LUX+DqGLqz6uPt2WPyNESaxp9KVK8EEhe6elO
mDXON/tSAJf9QLBSeNJGtNrhgdxbCWqcNWtZ3gX26LpweNcsPicjWfV/cikD460djvhQStwBU1in
tTJKKhMGU/7MeN2S29cLFMyndOJJyLltNyi+NKKKjQRk1lpfrR4lUmMpal2W3kYicBjbwrcfGCH3
nVBnnYrIV1pbGgR9VenDLsI/Bo2yt0rfXnSsPViRcNEaN0WeUVb8BYsQ5cBhBGYACuTRkgCk6QFa
P+zh6H1y5JvD0PCao16Cq8hUhojfXEvOe/ErVei1uIobKHUoTIHIrDqNuW57uUfbIleopVDhik5o
rMEjhAOYuGwPCoIkaUlm6bkmh/zGA/if8y/8db75VBS8AViZ33oUCIDp+SNAbsgAanXW9+mq8hw/
UtCaUSOsn6dvZRULFueE7QMxzh3sCUQhUuiaKpCRjRm8HiSkhXC0dyawaDaF8HU9xNWoZNBRsg0k
cIaL9pL0gh1bIaLuJnXWfjRrqhQ4ptCkO+k1oVXdVFbo0u+c07abqRkYycY+p/GB8ntyRjSkd+J8
IoWyKEAm+6AfK3kVamve8r9+sYjvxMth9yo1+byZF5suB+24zyhgELPw5eSJoosoZPzLKyH5bNUf
hg/ptZv2ubWu/Zw7vVrVPo9CBR8MqaDtQ7yKd8VeU6KhhqTtb0SL58dAPfAQVnum2ed+/pj2ZoS+
FafejVNgd9ZdwCxD1gvI/lA5sYpeXL3RdDiwIeXAO9OpjYmc23u1xFixyl25bupdHjvtPUgc9keK
roCz9QLZmErYE9b7ETCp+s4+eg0bUEX6Uaqhe4sAOXK2JpkZNN/7gAm5t531sP9YH2MV6+zrfbCt
vSBDKbeYpZTJbhN25HmL9bBh38ilclAOyLym59e1EEKalJYnap8AHQ4SGYLPuN0llRn9sFzlubLn
xWRkm29wG7N8oFNdvhVQMgzOw5rqeJCxE53yfZCfHRutkkp2vb54+Gd0pnNGnyHAU9qt/KymuK3A
o9V5ESV54QybhKBsqjbd2DYKEZU1uB6RglBV3uQJDzyrZvxGDi8SIOHGsmfpbVJIgfjUc5gps9Ym
gAfwHDLfk6/TyiJoVgI4tFWS6lpGV0ieS9eQ8VU/hDYh3m+V1vAxQKhGdHBpu05TPCsjiUJuw/LM
EcGFp55Z6v2/UbBL6ffZ6171iVgxNzdeQ/z9E9/8o+/0q648RDijl+a6bCnuNy+jSNmv1Y6Z5ZyN
e2C55X7pGcfire8spzb+cUK9W5p0JOBGqPIOW3Goqb8oZt3XavflpexSI1O2/Ekic+wx18Y9mu+H
6rTVXsDmrO6LfxoLR/T4IKi7Py7YDQnrTHI9jATyFVLfJmbddmgbf9AILCyO2HycRShEQMRMEXHW
jPE7ccvGa3VSMetzmGvD4gLJ2OqixQD3rm5GDjhbEYCeMXfFTWYUG7eVhXDDXlvPukO3zCSWxeJI
BNyHH7neV5k1MR8vtWMr2deUp3PIC/+4F9QgaQPoZEwK2Iq1L7XiSaQ+d/CbJLi1u4LSZaQIOsFn
ejPiwx1AurIqJSyENKsWVVlS3SC3bbJbCQQ9S7cnmE8932NwhLqNxAmn9gSV/5H61EBHqbVfZ8Mp
jGm/pMxQTMqBFK4l8x/Fw8soQwYTGRMdI/cP0YxVLl9ygRdnl2RidQDeYwtrjb+GRKh22Vsa2L6v
z58lUWUqpG/wWKVt3uq8P8uk+LbukEljvZhnDrhkuINn311FmRsvEIGjxqpuN0rqsOq5EBChEo6O
KuuP81mWpLjcye9ipsiUqLh3s+yuOQWXFx88eHNrMl0jYlRHEtLrVl6TP0icF3p8cezI018pN+6E
AU7+S/Ny+8AXzFdeXRH5JKwSkJ2mdXkCRWh5geX5LhuwLoKBvsxSg/4IHt7xr1OrvxxfRKFEzQDO
aBJq64giqf5U6uuemvigYuurggsrsuxzZrbdgSfoczAts8xjv40p3jjg4GR+Cwlff+qkKdIsrpm9
C8Z7BuoLNy7bgnjEZH3lc804VuZ14Krrh94EYlnmwO7A7MOM8xSBHGZS0Tzu60Hp49sESdZuFlFf
oFpcTd8GfYK+mC8mOiGp+uqSFm43ywo/NF8/Q+zBmtI0qytTwSWykWDCSdUyoFy6w2es2pUUVxHY
Vn0OGl/yi9c83WgX/RnyeuFhZmVlvJZGW1ep3Z48D3XwJ0N3ryZOIcJCaQE7xoE1v5HK1wF4BZ+0
ez1mYr93Nf88CufYMuJ7vxovOgc6+2aljhD0XkqnsBcyTkrZ/pDH1j4kFmzFuddtt840fy+ICUFx
elfHucnslZZsa2Bmhnm5KVXOc3XZP6PToJNYZY377Z+vN1WPeqNXtOq48si0pMA3k9m3uKt0O491
kZKm1ZWmHMtplj3f8OXEXioiyAxy4KZ2rSARMzCfQjnrZ/dnblVLgEPSHc7mknJ1biSD0rOA98T5
AiKoUTtZaNIGVmmR7rHbRBXvKnAPdjDP2bYrnUE048ScSdNj9oE1q8Fm/BRlD5lcuGIJ3gmwmQ3c
NKlugaB16gTQFOB9vrQ8QvuYZq5eViAobE76TzgjK62FnG+SDPad8Fzd+S3D/kqzEo17gS+V12SG
zi1+aOJukUaHm0SbTpwTH1wt/6Val2vbhlyvuA8gFx1v2mhf9/a9eTdoqYlhfq7LzgcKJ7KiRJVr
I5AdE9HAqtdLYF0kWKPqMUthu6Frb6I/TeNY/YsCv9D3S4mcuYIn8P85rDgKg90wrjustE4aC0LM
Jcb94D1bvytIsSwdwClTzp0WNCXQRdfgQ2VRXbXqe5dZpEaoQ3P5ujry+SXjVTxUIT5EUb7x7syK
NZMVSvwKq+HzcyaaJ74AXrpzAdBAIvA4HX5QNyH71Umgb4a0XzdcU0AeWtoDF6rxetDyixFYNfdL
8J8tq5sPP0vrTwNj3BBu0aHakGcMPL7O/7O0BHgm6B3Tw7SPvD+Yj4BEBt2GdiEmikP+VASkorlJ
wrx+4180RVP9+QY0kzY2AhGEzr9vUOfH4CZsv6JiPJSEQfkbFYds+T4Fbira0x9jHRTU7Ijb4QiQ
V7/5Q7VdIiZztwALLvKEDcFrncsW93wxhNaa9iYjkrw8DVD5LIIf5tTn5DtDdkbrj63mBskyVa2d
R21aXJFmQn9lS1MDfV8qyDtNhIYboEoLg36HYTNFxenQpzoe6vRHN5th+s6TemQ+eAbZiL2DT+Bb
MYyRm52PujPulqjfpKS2C99JRCZaoEZh6lKh/6Mvrs5akeNnxt43NacRHbTA9k9kWScBO1vYzKey
Ve/XNzrFaklX6ZetMIAF+iI5iBYLzeKvu57O28nFF3bd4zdRt9r7D19VNa+jpcW3aQtJzCZbMJO/
TaQmIij4aJd0S1zJeqMet4TWhZsJ8O74LEIf0kIp++k3wIhj4fQk5grDxcIzdTtxsv/VDIE5a9xX
Z8Wd+8/X/VIY3r6gfOMYQZEBoABt7fkGzPms7UwXtljOUyC5xHXi5AvP4l6hE9urhYTFVeaCkzOU
h8C31tXltwWtqhIDF559+mF7yq4Fb5JHUXNHj4gQpiVk2aREtrW672R5itA3gahkZNPwL4/E+yst
Q3CHe9Czj96psPD/TcR6tUF6uk7ZyX9O0yb2F8UgzmeqQzScYhQSAoOxTgyvqnc4lY0R00j4UKHA
kivc/+/PLHY8jTll+SZHxi5t5ZhwbwLoCgrkH4+6Zx4U+2w0V5gKNUxYiSGm27RIVI4WK4mqW34N
oyuPmNZHKvp9xBO81gk+LumiZ3kZHEBIkQlS7eD00IObLqXqhFKk61dmertQWElPvs0Ts5Vx/MLY
BtOKGMPmsqlFeP54MJHA24TrEzx77272ynbi2H0apXzIYhyzx5iXxSgU/6XMd/HrppK6JUXMG0FZ
7+H97LyEsKh3mKtkTcijYIX6Be1hMIfV2FKHaHrJo7GoUa3xfcD/NXj4Af3KiKOgJuD6zYASm7LP
IFKGYPxK6L9/mbg6ijsrGm/e/cSA2O4w5uv2qh+rVpXWexvcRr8exfDit+KeEKIwNKrrtnZ8Dbr5
qNGEa6pcnmEOQr+3gPYXmw0ptCJtSHWP+QWCwhLpQ5qxwhh4/Sur1ONisHg4Vkg2tH4eVzW2AvUW
aYtHFbOGj5QY/FunfWzAsI4eG/Ey2tn6r0DfRSUveSU4EvB84VNoFcszq59h4r0hIZOyQ3tev2fb
ae/4eWqgIjWXbme6G0jDIBwFyUArOgOj82JGms/5BcmLHZ5sYs5ga9Wq52ThbEXGAKPOl+fzvPgy
NcavxFErqf4BZ13WNbdoCeXOZQZrxmDzsZP1px/53ZJXeSiUfK6y1ID4XoBlQ+HUqwKy58197A2D
fvz1vEYTqjkPdpTCKW4hCopKooG3+JHtRZa/J4Qe2nXtw1+yK/Jwh7HNs+76SmQ5s3CIhescfX3B
05W556v81vWv2qZY9LAddioDbgJaD+dczXyKxJ0kslq5FYWRDjlt4TSQ3gqIXvFqPfddHIUslmid
hR9X7k0oUTHG/JANqLuflQ1V+b+9ykEBDtHBxfwbn9iRly4NbCwzMTiG9xbY1lhnR0X3B5UJvNHn
J8lzx8LVs01TUF529+z+YVYlnVarW824hF+AReCRaUDANJGSHoFUtlxWDkYE+aHAxPIpfchw+Gdz
xhh1ULUju8CIREnHZ57W1ooInFujAgxNrMCT4tnL33cQtcQtUa8xHFDPLoH2uuNHhotE6VxKykpH
k7XUp5jNfTe2Qi55Jfpp9XMgcl+nNRk09wHb3kbap9hWNjRbSbtmvoU+xlq3Y5RU0qTNI4evt12T
zYA6V3/+nhNqkPTbDroIn5keUKVOtouLHKBSFUp/9MByznFvEwWBc/FMXyroP7MDn+RLopOvsC0D
vscdyMjt1/nHbr9ql/dRAgl7psRqE8yNsGsXitL1Tmb7jl1dLhyY19hk/qJNAaWo2UvC+zfVjQ3P
J3OzjCHgEygKdEMOlMXBpF/UE5KoL4+KA+b0WW1kyYUSCNaJWVXopcibt9TH100mZt/lcZ815Rv9
bxPBc56PX2kI3NQtnDTx7UKpOQmP9qneoB1JbZ8l2EnfYBJ/+Z5AgvM0yvQ5+z27XbjNv3Ix80Zz
heTM4SAHs28pH0Mjew6ivZatIXBpyZKqaFTDmAu3sgeNl7lu/NNp8i1Dm23dsEt/Fmg8F7+rbGpH
/mVDtYX4EvgjfhH/ovgS6lNO+5qEZqTQnF5m05yJJWEQqU5oQ3YwVnSU5YA0yK4CQXYvywSIYuSs
O2hMDTr7sh5sXxqiHp/txVcHUHCSFdmTl6RHxEaiYQVN95Bx0SKnrE6XqxjLN4dBZtdObks2xt2G
YXVdh5bbpAr62NuZx2qQvLGdpgM6E/XBaxFk9l0rZtUICrbZ0guplPsjKgQO8vuwIATL0qFgXt/n
NQ0uLSoECSbymn6Bs3hf7QhtgLzaM/rEsm5MLMcNgu741hII8xu1s853M/g4s/u9UG+Dx91xDBvb
hHMfeY9sd1hhPi7nyQGuAVLiMuvdsnoreGlYEFSAabXKeFesUenmi9GK1/9z2by2TCoTU0rMed+C
T6nWAFOnzMyL6wS/Jh6hMfY1BXJ2w4RsBQzEWgmBZ8x32B5Fyz441Clu1wDRg+IQTQLmQVGqICMr
+9hjO2O02yJdK8tjHTyEiG4mXnp+IQ1fS6jiEBUmzMDNGdXm1xEx1VsVsG/dVvXOR2BF4lKn25Nz
t87IukMekrMgPpRGZT8n5eboVSU4RZ821pq2sDXaBzbrCH/zALGcmRKqYZ3e3YEdbArq3axILCAR
2ew4J3lbji9HrO2+iQeERdpwbm7/1tPmYTjbCctMx4UB+6T1xa4wprUODMMatefmCY7mtKLJytrH
G3tG2j+cOql4MZLprWzpsO4BFEsw0gwNyhatDsmI69hu14/5FShuh6gAVZtA3NFuogNnDN0cdxAd
5zEWNMUXEeCRFPBfZiAVi5LQEr7BGfPMT9bvIwAYN9u82zGxStF8g2TLUHqXD0SDxuV60U0ub41l
rHlEqjK8gKvKawfsua/q4U/gSnLj82IKRI0sOFo/stnss8EiOnjKmxHlnQzJlRBULECVQIIRkdUc
Dy0FObmWlNAnf0cfJOR7c3lR4Puz7ZZMfY0yJXwFAXiZMYWNsrtVPu6u6pMlg6d1xj1llT9CevKI
EQCpN5l2+Mn/83EmRF609azxUThZk7qWhLUGzezlQduT9Pql9hWLFoY7Kf1owviUUAkFJxZgLf3k
v0zUlB3we2a3/z6B+k3IYEqc7VY00/iYOpW2ThCCHEBy1gE6YXyQsFSzTHWjACA9umAd0f0TUoHo
6CP0SZkXI6bhVi9aMJT6RsGYZxIv9c/WM2M6yYoEVvfCl/kYQEBj+ZdU8dqp8osPg649oWXFLcIB
o5gXNJBrk/0OrjsrQugqTE5MHm7pX07EKBvkJDioFzDUM3Dbw80URF2Ya/97vY+2Guw8NVha9xdb
vmmxxaJuZZkiTI/h1abptBDbVtwnb0rBU47UhVNyxVo9K+EbRoxCrUpQAc7HPqgLbnkN4OkhLFKl
sEAHd9ZPND42shylFNSWAhUMduxhwoXS1diFasTv7vsgCNi4tBrs5yyM081FZWO7s2QzceOYQxn0
ZFSon1/1nzdo18O/OuUvnYy7tjOD25h6E2QL9A6eSdbV41/w+f7ChzUgfeXVLaCf/4ry+Gyvwzds
MIcsTy5r0irc1DBg5QrW9RKr5AOhBDojYo7Yd8++7SdCLIAbq+LrWHvSbj49vQWNDqogn+QCoBKD
O6tf7d6Xj+ZN5pr6lOjC3D56tU44syaL/+7/sSEz0sj2jv4VxbOEZ9SXJvolUxzpXtk60nTSBs7H
vH9tTjDOzufke7gRcwg4RJVMmXL0+h2NkarmnfH9wFHezyljldvWTwrxz/BuiPfSs4hWHFcp9Zvg
O7s1Vq5nKodAjqVcUn8GssucfLNW6S4gNJqV0KhnzJaXudwe5lSLzD9T9A9LfpHyFjqoYN6XXoqD
MyYEZAnVWO/tjOI5wJ+flG8fYqRiNwic/7xlIZ11M6OHMndrV7EbTUVvBVvbvZnTkIytaIQcsaau
kvURxYfXPSl/XpT0VCriFWJOXK+SwZ/IO584EM5xySGMhyrYGMUKMRT2T5u5bItG8QjOiHAtWLd4
1OxzQrw0KYKVlmq8Fh1+kYQqCcHmcsPbGkVo3BQnr9O+Q66olYGSzzKpacrenMUV0YL71bZobyGm
ArglXbADwkJokRCGPncEVZyEzRk/U5AhOeEwnXW1BtazgkIsh2J/aJhvf1pj2eXeGRrn73NHF4w6
9vDItISfzIHWAnxorFtmvLi2X7lyLn01GQgWn68kEWCo77gCv+gzRiIub3emFJiL6MdjFyp89w5O
QQwY2sbITsOezr1cQqfB3lW3yZEFztWh+CkBXX1uijOL4dpO1ZUL+SXZ0mhnANOShMsgv8nq3jHi
5VtVxrHB7trc68d26psnXn6Uvn86MQF/gDWJ1AH50TeLoBmcvuFQS8AUZPOjNbfsDlsmgzXx+/DI
oqoUlhuhmQmUQBDYOsb766EFI4rH5e3v4pLDnWF24CUHq+3hcJ2CyfPmfBEo8WkHqy5XATOUbn6Z
0FbRdtYchaBdEbQB56xf7lg6msWb/gquw//SiaiamQ215BRpRGu/35TruxKP9lK1sGkZ1djs1gFy
W214K8Ittsbh2OoQQu8Z9snJCfVpyX7B/+ZXHhvi9aWR8+K5kG8dIQeGOqLNDhNfqTX/zf0vC5x6
jx+cs5R/vPmTEsen4uGa8Kjt7ycu1YGUqulTpX0ErgLHEcN15Ub8E2GxhTYEunkizoF+AnGEiFnv
lmSmGMZSdAUCXg28YOpH/ldB/x1/Sp8tOGV+DJw3u1GWCWdeoeubp3d6jQ+ap3Dv2qZZF5YuRyU0
HobDMy5prfWuZrePENb5bBOOUP0aoJ3EqVUrR8aLA9wev2Pr4Xgaxwk/q2fjTKGfHHq3Oxql34fn
TSGqnLZMTFFG3TqG0XES1AAhKn8fBv+oFkWyaW5nCWgTeh0v8RfGfuQVzK9h0Ynb9+Y4Xs6uyM/G
skslhwHX8mkHhv3LzHcfz5A3N66GfXpA48cmWmQH4dqjCeKeh4/rwOZtxT5eQDkSS1Rvhk+cu/b1
uWeKfMMRyqWnjW0+LpW0fpvX0fxYv1AxrAhPSEOT0DBRSxQEY+HnlzpwO6hTcwVPKAqDMwBEYEgd
w2bsHO5utndSWGeruLman5TB2koSfzoyEOo+/QPEMbp+LRpbkRvAi3+mRsPZT2mUI/KOaD6o6PXG
C2MwK5FrlxKgySbthvGOnMvxIj5GwQYOXUQ5xG7M3jTlgFxYQjpnvY6lZPIZT5Qx5dQZ9tgpS2pW
lXMKw25qwOX3QOk26mM6p27RsaOxYK5BLTKOUgZUpbeGvxpcN+J2smhQ/4RE76qZsPToJLkN/olh
OmiEV7qkhO+7uZN2i+kmwTFW2pkO2N71IczYoajxN05xhELcaEv0O73wM8v2hJvaU8PihftD6KAD
0P+rAz7UgdbYZScp4n0F5OAIDaNKTgQJhk50AxXysvlaQ2svxjndog3GMmXIrYgYD4ZVE+a7bxvT
JTVa17hLQE6FAOufaouoa+ERmBiK6XKoe58/ThZj8M4s4/2WgFLiquEY9wIBqfx44KpczV4aFmA3
AodwDyd/32IbelgzgR0IUG4ATg6Ac1pgw2FSB8n9c+HIxEGXJBmL1mTKaLhRSqizs83HU565kGNP
DLTp3j0YksLA4C0+957ml42JDS3Up4riC7Lv1qDaEe/SDXeyol4ZZEsRlToXMrcDmCEYzNWmVO7W
7erqptSv9bIpGkmUuTaZY/QNEDbfGpaIURsMi2JHpZg9jF2lsFn5iC40Jt5zgXMUAbMYEXdv6k9e
7u1X7ZE2yB2Yp7HpXCUFZ9Jy2MnI7FBm1p+So3CPjsb05/HKEkZ8Yg6vE9388d9BFX09ug4CG0Pq
0UDvTD0XwDy9UrFIN8SW1jDWEeVXIxhurSjAtVVH9pndiTp8cxzcr47RK/C8lcizrQkh3S1P5ydM
t9A2/biT1j5WpXIaiFgE52Gcnk1ZlvGgdDenfQXEkvC2jR2f5/J/5DgIqoxPvLcu9iVRxXlBlRZT
6TT1ADfUKptYx/pfb7lmhk4Cv4LUriEFLNF485INEb0pq97WZjQslg9AqTtBIFfHa1IkQ2Wwdiha
ySFhYCI3WngRpNWEfXkPOVUImxGOZeNFzdWsTqr5UQlxZSqSoh1d6THPvsc0rOsYy+vguq9bfDIy
f0DFYxJ5e9PlfK8vDSWagq/MRtkTginydX23cUBOaWQgdCKDzqbrB9EBP/hGKb+x+Gev7SqcjDGl
7iL/fn1NpnlwUZDa7wOQOx4cLo2yv4fc2hQJzOEECnaFxO/gxu0anFxLTKUbHkR31gf7yJpKmBKh
IpCG+8i/8phJtiuCrM0AMdI9BmI4pBlAp0So9BRwZ1LWedAWPeExekqt7o06VAy/g5SoZ9LOX7H5
zp2cKONXWZNHjHzfpIdnIhjnuLZ9RphAgUTwsuUDy89HbY328RtdG1cd0QafG4odj0aRAbq2q/vX
C3kX4Da1ohcHrr8Wdv2LcKEO8hLKMeSbL4fZH+Jy89nHei5/LkUa3OMg/Z78ZuTJD4JK4UOA+Phd
jOV3wDAUFTIJKiQ6TwFhFCQb95XQ6s+4svp5310pC7rlz7ZB9ceohHudlaOh8JAn8c/Iiy1ADtGF
zkmWo6FYM+GVBeAZHYz0hlYbtiAdoSWeIqyhKLzczZYSOvCjCzIJYADMv6OdVDIK6S0L4mclZmVX
W51jB4bzR9LYwY3EAf2cMepiJ+1hTC1WDgxPc4Nn69nn22K+GaN73M0gxtTQQV2+PSOn4bn6PQtC
fk8ez2v/gXCy20RTkr+WnAHBh9eRxP98V+kGDQr4FRTu9tcpvDc4jQfyscc9E9gpPL49D+d4BxFr
8kflxdxjDTDeNgZtMCH46CDQ3MWDVeAtWmieOHTjtt873uDFgYmDLYU9k4dlUefNx1gdrxMf5IlY
UL/EJn1XZuUtq5acpRL/4F6PLt80V6OHYpdLAMKmKaTfsFXMfmGwBU2zNmwHZ+xUpJ0Kdny8BBAd
GJ9y2RA7pazORFq2uJxXJO4npz5M6gtUb+cX7LwIS37qDM42InbK0GN1+tIOvWyBO9TbRddqdUQ2
xaHh2JbDJVkrNFFwPN4Vf6gW860gkiPirikTgIjQ23CrbEVM/4C9pdWP5VFor0xt2Cq9XxuE5aeg
tP43lub5mbmhNgqZBuC5HquCE/eLSRlFyFpuNF9Am6OIKAgvAw4HU4vpV4UKGgKANgSNwSrDQPpV
I2u9JgN1XJ3R97y6huecK7yXBCROOdeGo1EYhTnuQ8MB6b9nLB4v6faLgl7yCLxcexBtW7xk3y2S
dxRVYFlLCFHuWHlCnjCBm9qiWho9zP+61t+2q0jPuphLOGBBqAPysMZf42siAkyeTSwKUL7xJIhC
roiCzegZKnFfgFE+z9i3XpoD/0VlNknzaR2egE97kbFU+TvQsxMB6ZrADZ6FJoqRZh1BUgVu3YLk
sz0gNJKzPW03ybIHvxGIoYSbVd04/wA8Nxr4CEBkfer3MX1cPSaFymbEQbyfVe7pgDv5mzvhfpdx
wi5B2+APbMdwYUMHe3SZZx8ZC+Rt13dw1/7c/Sp9h6/WzOtCGV/eD/FMTEFPQVZefBH6EblVXs5B
MhC+OHhZOguW/8vtAHr37Ur0hzbtiJFA0BQZ2zGb9JIjucR0BjzarxXqTbZ3I23VBdtLsifUrQ3e
rKvukmvalb1ZV0M95tEAl+9cVPnbgsIoqgZlAzJM5JX0mrsoP5TdCcZ7hEpZE88Ckbsk0x23KDzn
uL6on469eqvXFMC0V3gvKuWz8qmxBUdaS0tWHCuBS9I5CVJkKiLz/uRtw0gVfYSVnUTiSRgVRBie
twbpwg1Z+tdC+/AwuTknXLKIdRkkXuPNMKJNCzMIDlkzQLxfcmItM+gO7QCxJ88Pwn6glFuigDaN
xaYa9c+iHW/+jQJYKd/Lzbh3lGmkTFU5jHbVMeBXoh6L7Ed0eMpUC0ZNw7mgDOQXgEne2GB8lv5h
NR7s95+LnT6OnWjZ/OeB0Ud2kgJanyCyru88I1+aRwYs3IWWsF84k+lkXZ+1hahJx7SzsQQiSYxE
qRFQb5jo8OG97ohJ5ytKIVzWRtZ9ke4R7s+FXfQOY2O385Skd2IRJ2PRhNnZWpvmgX2aSSW6so3A
xXQXMxSZstJNtuiJnNPq4Pj/2B/LYlEsG33EkyI+PHF6vOmFjdHC/2s4+Wi+fOK/l7aZc2X3mMHu
fB9k0G2xyWKvl4SPsv32hIripzULFLBzxcBWB/E82ZmaUBC20h1HzWsiphpI7oXlO1I92yRMXzAH
SjHiXCA69SX6NqVcEAXryjNE9m05j1c8pnsC9gActigQP2tjy/Ch8MnhuOYxMmKQQOqN9WSGU3gd
uOQhp2JVa1ZgllaZ9V/RRAFts3SExO/PKU4J1RNyEmnyp+/kdJQ0mryVdZu341+YthAxJx+UPJBa
XG+IWiKUU40TaHT+ER9kID+DF50zaoVpADoDlZHKpzWuZYU3NjEHaCttxMOieLMhSUS8WTWhWvSB
eIgvKxz111pGZLBT8hWpoVnzrOPGgtgcZuEbwuz1OsLbeEzDIkp7QrBFMjR2/1SYaX+ripAbrl1g
8LRED3n7537ZXl+ggVub0ULovut3VgfzJXjxkVa6K7kDOplp1qkOM/0BgGHrzkN3YkGHdv/+R1yi
7NBgxbm7+OWg0hApql/rsrK+jNlA9RGqbxbV6gKpnYqM3s5VaS8boZKEbmbpWJvmpLBQFUJlgmiP
lIlKu6FVnGph3tZR8VwY6O/6UxLaYF06wJPSSFmkZObtHgQwzso1w3VY19RV/BYRmlDxJu1MEqGI
EJvZ7WClEBc6OVOElyzSmBiXja5iM5QZLv7WLQpMiwuSXv2zpCpE/wphShexQDYnViGUQwhvifwT
Ym1dHg7dPtFmzwk57GDocp4xxUjySMHXv08YEWoQTB4k64uHWUjGwAdO+YdI7bA+hb8WCqKec1iM
bXEK88Vg0xgBBjJkLPjoFFd25ophMeOI+jgrPT50Jym5Q7D4Cyy+wsEDUQ5FkktQxYFEJArYcsP1
8maM2uMeYRmV08aY+djXA+0PSyt51hDUjWosbIo7+bQJNVQPcaV3YhrOP/vyUSPKMX5h5zHiexWo
fQNVSRYKN5DoEzSldIZJvSthsrodzIf+jxFhY2qp06IdswUQ7oNdlFkAh3+KPRULaTwoVFoAzdDa
ohHnwuTZZqWLHay9ZlEYuU90OsIx2IdI+jPiN8e8Xg0YMXV6JhP8z8ND2Xey2Of+eLxc5ymPwU5O
4d0Cw7pubHTnc80M/BxinTVr7ssOlow1nF63qf2DpYroGI7vvTJc/3IixImu7BU9cOK7kLZ15xyn
ZqtqRLFdcvL69Np8ynIF+OLCKX9T179RTyIdHXdTLM+bafOUawEyxRnMh+lX9bSJM9qI6iw1JtWI
esWsitJAEU+AbfLplyn7XuYuoQfbknQkxhhQg6wam8P50exivmRMEv8MFhHg2SBgH9i0evC/zlfQ
NYSEPzzVqlTo4SZIh6W8hYCpa//r9ZVLFT/R7yk5E2/yYFPNInL2wwA3qu3vNTPSA1pK/6mxeI6X
iYHY4QoZvXHwG1Ve7+D+23CWcHs3DrPACfz99Di1/a+gB1f/bsIWw0cpG3ZdIIw9QV2m6ngVlIHT
QI9vf7NnCZMS7EZ22WnK+8NoyByUCKOv2MclOzZ/EzmrW+HL20LDXsSTa5WHqUs19Zju/8QUZSlL
ztNI55LxztTGn1h1WUjHZelWUuLR+X+6DgZRrirziE7/swLyP9tESly498EgiXzgaAT3NAYPoo1R
JKmRVQJCH3SZQ2spvwjwcPxC5kb4aX9AprGzxM2VR60uhFZJe/haByn3sejdSGfS4mimto8ZormN
Q7ONn99XT3IHBVqXBHSnf/pfLozh1K2xzXf+QXOT83PUJOEBZ6gpDAynfignE1R/TKxgPH+Ud3yt
NSOBpb1Y5W8e6O+esCnDXKnwtMfgXySdu64mGIOnW6X+RT3ilMjB4T36Bgg0bWQh+H77yuRduyzC
yPpivPCbAGpzFV8Q7X2vJ9uefPL7f0NoIen5qAf0H4lIuQ79MONUtWv7fqLRINE0KEFObIi3cvEi
XBCl8ry7ievOYvhE9DyxOGrclfBVMepVYfQOSDKyfsLYqf1BiAaA8EGh/ClJ3w19nPrbYI4tgH19
z/+mfCDUkUMaDSkVflo3CMIWWzpLF6kGfj+dL/tTHFO7Rq/AjfOCz2DsyRvPMz/WJewVEiHYUESK
4Or45i28ZwCZtCZj7Co77OQUcGM9NjjXaeHNIPe8ZO51uwGy4XPotVrkTR9EUQRSJ7xahxjcPqQf
Ao2GfZKj2hHw9YKLmwBuFuNle9y+C8lyIkh65DtA5/+BSnXRsKzJWQeoYR0SmTDpLj9qoN1IiauC
N/g0flZVjHIiQJHOD1qpfl1G3C4DTJmObYqnBV3rFm9jUAmXHB4ljlpzkGf8ztDZrcO8cZp5O/Kj
BPSXocQtqG4QhCuZG4J3BDRI4y37sg4+13COxbR5direJeLGe0bMTa5TKJS9js+3qJaPbtw/pKjA
9+ZZBmXuV+xggv1t7p8dDm5nfs44tXZnZ7XxFFxHjMWqPXp5SI/u/YUat/v0tUbgHNu06cqPUG0s
Xym+UZtcBKlapVpWcO+myfib8WLz3tc1kcxAvuBcAyJC/mlPssx69LfQ4H7JmHwVt++NaX5+JY9Z
jVAm/GRdsLqQ+wzo0sAt8bQ9sc48cxvNPJBiGvDSglW3m+tQXgfOUOb+8ARzUrH3X3Pgbh3OiZCK
GUtPcD6k3i1IV6E2o8wVkaRQPgMnuqhBXf4G3BVXaH/hp6bgUnkbPJta5/9JKcAXkZXUiS6Q+O4Q
ijCv0H2WGTy47TAtspjD3CpJWWaSlJtaZITfAKn+j15A7i1LexVrMr+4G37ceUrVulAB4M4nbaBH
+fx1Bf79g3lzA8RqGCEDuacw9TzryVgfOlL/II7TFdN4gH+794Lu7O3pjpn2IN4+TehB18DqbnfY
xwZbX6GKG4QROzP7g6/TqCTfro4HFEHsvdKkOwxfC34GGfgnaqj/JAt/DMu8Ez00VNW2xUurN4yM
+14u9CzBflGt4obQzZzRgszAfBWkrpZa1fn3uamcqpMbSR6QXPlo/V3pLPW1hbVCmwiaTAYXAYpp
ABeWc2Intk1oQ80nKQljqtUxOyja8dvBf5N4NPY3gIqaDWY1NpGhgUd+7MF7AbRMQzCN5umCxFGt
KV+jvtPeC7NN5YpOo2apXGZMbvcEnMhWAofSaqNZvurL/xYmkmkLgpTofErl79NrMbpM5WuzITS6
e1gPRF+jsODWHKeDs64gxjVP+skoWFYZYE98EAWp2KIuWWwtkKHWGewJFhNCfFFg+61iFXIBnXVH
+d42sC6CJ16zlTfx2NV5cX+jMtqKzRJezTQXmu8uxafal1Azi/4AVp2BARdX652+1ORUue/NfXmn
3x+9pLZkv2iIU0U+W9JEA5HjBH9iBqNRv+oZN0Js2/396JhAc6054SFb0pQfN7uVdxfI82phDwRb
zg8X9WF8wExTwxp/eAYVpPJhF/XSkC536Kvy10dVUjLhMdtAEna2wehXswluFTtPBYsanr32AO6k
0JLMJmqSd5oVeeDOsi8xBbFLfOjRvjpM2Ulcec/UMAjVWdsCMJ8pBk9csGF0FfOcSzz2+bvVajfz
ZqFDa5XqQu+ot90Kc2nLaSIb5XO0GYHtll/2UfWDsMFXdaNNkcxQoIMsg/bLn5wCBAESzL0VP4b2
K1JpLIS6MMNas0E7z5da3PxvnViHef2H8g1DYzhLJkf8vH0KMaT6S9FfigyyfQ2Eccb2+d0FBIAz
tVh40fYg43lMzjRIsUrWScKu5ysEefFl1r2WDmrP/PnkpVSzkXWSQKsrE819EB5bpAaj0/TZWM3T
fOxI8OUTKIdFcomMAnZr8iZt2Nb8IppUwxn2vlq/hz/apg+2Aotoy9Zn/wJYso5J6ymUCJpI9W8P
nLHBWiiK2LgzagP1NR84LjNs+90Az8g6/DWtOLWLOErJjgiXlAUetDDNJdHuYOeEalGJR1J1a6FC
E8QLAgOq4yiYiezRfFWtjv1NS3yzvhD/l9dI6kmZmbtHniNy3mhnBpA1P4+tcLbXpnwDEqSwwgAy
+7FIz7rl8v5QZNNWEJ/Ws0/k4YakRztCRIu7GeN3TdzsZkN88CUvUxFjuJ83ayESkQrLpFAi83Yx
etDFtaY0bkYf3JY/g1FsX3Mk4xO69vXJhrEBPVuxK6xPXh8kRMcHMhJ/6uNfzfFodnhhgHMrejfH
LUjBSi3O0vsfJYLNq7FsRVXQRgCrvAcSh0t5SozZLgIlGrJDdehJVI9ws8ayDq5pHI1Vlc03DqCI
8/eyYS6F9UzXFhl5uaaQZNSdGIcySdRGaLXXIb+wDUxoq2o29C+DaulL8dhqxvGSkAN2mUlwsvx8
bfHcDKyOnvgTY1YAD/ZvlS7BAEJ5huWDFNahdMcBAkJEDNvAH5xl1FR3/givC8aTC02yT6sbeBQ+
9n6NngKxGRgltbOKP919XknFiAr8t/Zlp5MoU/uc4cpbV8lvXLCVpBLCi0kYjl5vwEmKntJPHT/c
fpeJ9JxvdOq4bhbWSI4gT0W6bX3bAs0U/QkxKzSt8GBCCLbQWKqwMctuBsR8knd0f0kn/wLFf+Jg
/VRamr+XrmJlsGRaMVg3NZSB+9iXdeoSv/8rVPZPELLouW3emXoEkzNE3biLruDrN887SkP8wixA
SOtEFvql7tBFuOCs8WLv4oj11RmVfgUJdL+qJt3BtTzv+B4hwdbOnQXJGkFHjbwDVWOhlUzXBA2F
BwY7x8ws2RbFaKBvdgR11Dp+c8AqjXxfU/WilQyCz3cEZ/O5grPz3Y1ZADyvzmipbneNLXNuLlBC
v2ZY2WCRvTYQ5nXMpipazfyXNCNvjoPC6rBSiBIG8HAVe3EdRoF3Wci80OBkqUVUJyN1A6urVyUy
TtrSwyYijJ8XWHTdPGNV9Y3H2DtCODSSbjAHrrtiXDQLTNBj1nAKnpR9mBie6NbJCHahOkakklnc
t/AoB41fzh9Oqm5BhGVoamsE1kdic0yXMuOh9rSk7jMjxfV9pjcQQYFxwJypaIkrGgEnBDr1QwEc
+qUXF+HKPQz/B3yKW2PJTABjI7QJk2pPY/nyNGJXJjXc2eMjrGKMXKYlQpdh5L/RVh69jtSYjd9h
VtoFtwMt3TyE7/DlEDHdXVSdOCHoG2mk23qZyyPO/amhmi6FFsHJMs/G0LTosaCGOW9r2Vqeur37
H5mnUwz04t1HkIIEpiGUYO4SI4zboflBkwoaoikVy4GJm/rkmRrdZzHuZ06siImYKQu4vFMmHayq
+uFUZ6rAiKs8P1hVlbyBTlA/Gwx0ZYolYxOCpeCpDQ5fUVPPoRp4832tQDZUT0LOnciyRIRE41/N
p/RQ0yyOxZnpAUriZ2as9ygxfMXAmbvlIeK2XnC0LnXt4kA0eBN3whvq3aJ9WOzTMmjn55dG+dfo
yU0tj2cEvP5i/CO/ARgFvUweYrwF5UqlYsWghUmPRJZbqnBo9/c/xpOa3D/EP8yl5UEgVgP85tig
NyYGFaMYWpQSYReTJlj4tLXwAsj1q1vVJjtMYPb+YPMwenuQccLx4rU49tjTx6BBXq+TXvjHetaM
1a+QCfMBAPoh+L4Up+YQF7uPVIw3MKHHgVRkcMVWsU1hh0j5NTFZnNLCl4LHsbgxKBYOgOxjUzsZ
Njq/7vp0/0X8tGQpAM8g8KsUrnN9YaJTq412ChWrXWXC0Kf/gjlQlJ1EnmRvjs1upooduG9WMyA/
RwvJ2g6q0JtSJp1DiFzWcdN+kJssiV1gfgSE9pvK4tUZsLyRXW5woKf/uvf+TaHYh3NyYGQsJnHT
+Ppan1OALEVlg6IOw/1U9L+CBBMo8P0DO8COHIBcA0sZvcTc1HTH0SvIQjJ6NfvINzANqWZMuVZu
TzTdpQu1a3JMxct6x6zajlrLHjBKT9fhVJWVBYncJ04ksaE+ffIj3W2IIXM+QOsY99syffMu9CvC
L/E100GAMYGoFQuE+k9CVcsZdCrlQnW1a6dMbACeKVmbfoqyDdZVGci/yUw1HQZhEUqJsslCSc9Z
S6vYc8sGh0nWYI0e877Z6zIfUaqG0zcOvbHJEOydOBjLa66JIy+7aprv146MLs32RSIX2XSm1aN+
NkfCawF5B35pKFuP0d1qt81rKFmgyteLDvZX0HjkqmGVSwedJL8l1c2igCoY9I4bwt2/repFiuQs
+wVBVbEhChybAdEJYrE6PKg0/0e71HrOc+ibPwPgtAIZJeRk8VWd1sABrjcCELGH/wZfHS7DboL9
ZVLtftZT189z8crtUjn+P4Tfh+RlP7ftmiKfy35aybyUp+6KEcpzRnNCNonfwoVwTmXSw6U+HD/J
g0Feab/SeTkCDZaTzjBbnSSQTvLYgavYEY9cKjxsgXsJIxXpp9p4ncgwanQRSQBRBO6OhNSAVL4t
ZDiPiAGu/2BWYlIBTV9MoSnR485dYXqRQZ8AQsJEhN/GvgpPOLiG8+U5fNtHqEt2EDtPDuLIvV4R
c9xM54nJcx7MivGO3e1bOKRZERMb9KnTYwNDx1izSmXrL9XuPOvHPEXY2sNEKpsXDmw7amzE1rPi
pPlVYnTI804WBVopXfHZzDwfp/S2kfQgtp0cJ8m1xpTxef4d274BLJUnz4XMMurggilBzsyE5x7g
/zxehuZtYlh4VIzKM/rj/EeHFt6NwfOE5h8nOjajMXs1XObQ97OHnxPLG/TYM+gHAFohDh37EVS8
eFNHAZOrzeYZdeS7LZW7BysGJgqBHIQAzDidlutDmx0rslmsQnx7GSKzLuYPNv7fVT43apoA782o
K0SuxsRmC9jgaRetuPZoedf88eF2G6sTvMHwra4fU0SiCdbDPbi8jBnSo5g2Ko1nnk5FxiTjyh0a
l+zmFh2mXx9ZDfl4FJ2bqGpiMNSTJs57uRWrbICFVak6iJn2IgKlRiYBk31TlWXd3fjtvIKcz/Hc
T3U8ZFehWCwuQv3w2heOzWqeYvO+u77PtxR13I+1eWNiQNt4SEula93Y29N0CSqXHA9aVg3/QuXd
DVayEEeWiHH+b/enTnd7J9QUk4foj9UQ8uwCteEc963WUm3X7bHkfwsDyazyzJZ3HEZgexwP7Ms+
BPVx6s4YkKAC4sjedbt/yKH1aWE82tvlsHgkVf46khXK3AkY5aEDWOzEtnqlHP/MZxfS2n1KP8rp
vTLBUbGG2qg+HqmYxJ6vwSfnEbCOSu6LoCCc6um+5mwaUEkw89Ylj8jKw3dY9zzhqT1Ewwmqo3+w
e5WQyDAyvYtOcLRKbi4AAALky/Gf8jxA50YRj4Rv62pJ4lKWF7qZzI5qlxiinLbWA4C16bKJsBp3
4ciL5HjjW0z5YgIBslEVBDFRHyQNZ2Vxh1mdeO/RuP1UGMZhNdGS7qIq1ug8Qf3vYqojw9qdcziY
YogdErypL3kb5MXZcBwgFQ6U/Jb0uE92p/OsmNbVnT6IapQv9/Ud7iLYhUJNFDjShIbGEW9RoY/t
eN/NjBVsWjzrlgeLUbQu1pl537BfYBwSbWaNeutswibCqN7scYeUKWjdKgNXlDtadE/uflshlxoa
G8eYggDuwfDFjgPAZ1+QUIsLszv36sssz3h8evuyaOaKdNjfOoOzDXXcNBLM5FazZDTUKAVwZG0t
7kwKHvLNzLAnMbV7V5aUqXpJzk8X8DlZSKulmewy0QF5wxhLpwYdWG8ge93D6VwNNBe0qDb1tl2l
VOnc0GotWrM/yQIru73Yvf9BNKaVp15/u7x7GD8EtiEMyP/3tTI6vp5IBMGP/MaFnwi/oUsZsEuQ
hC2so37JCdUCmEAmqI//v1Rjev7JdZI7KeySkh50CfvYrWk5uPaw16oVOJ4k0jfAW7p3Ox0B2qMA
2kWCyfPtzKIV9mAm2PrknHY+Sku2mGB6SzHsOoo8i12DLfCRMiI0O0fmYfRUHKSAqv8O681x4B4e
jq/9IXboOuM30+Q/DJ/nMKhZJZVw5azg0RwCcKHtm9E4tkZOtPbDL2Dcnp+vnQSIiWk6EaaacdIE
6JHraGDu+SpYc/mq0ew5kY88nUvq0vlciAq9AF9Soytq2K+SGAm2puyXo3nBRZIHc+TVB3f70eZH
2yqQuC1L4Q8+P9TBRwUp+igibEMYnI45yZfUX40+u3STb0Doc5AEYo5HIKi3eIotFsvh+s8NsLU4
xkjqHPFx40JRU9LxromS2AVFcqnjRXpM9TWH5Z26wlCyhn4I4bum5PSplTf7uG4bvNvvEXF9Q8I4
NldBOOAZg0Cg5l1YWET7Zb7WORcRz2WNnU8YNUJMaI6Yn69o6LDBln4bFIdi50mfl7lIp5T7nLzf
XGbftNoUcrkkfDNAY0CcMK9i8z5PL4LSb91XA1luhZJHlBCGI3+kU/To/E96lq7JZ1Q34Blmgu5w
fwR4pnaRJdv5vjdi42cNthG5FHx4MTOzYyfPdRY/Izrr8l9vlBlWuLrdOwjhaeo3LtiHAjMnFs2N
AplPqpXX9yrTtX3fUicfgRP5ra8QtePS2iUUtxyE5lIt1JCvS1KoXAMzedL9rhJXXimnMipK0zvz
R8qi9OcaoMWCs6qAHcWWYATnNysmyljfYSoX1kH3jaxaNok9VDuP3mkzhW2m+SMMEScOAuASF9wI
f9N448eV6Sipn0DgCRTts6LwaQdw8DkAa9GTcQtv4titcrnXIwuR/o4gUZ5RtorbNg9wR8cJhB3s
+2AyPJ/YJGqdExEsciSufLD/4xP91rXURXTNrSSTqvZkl/62jBUUAWIpqvSsT5rNJeQyxLEWjooM
P30yComyC3i4DD9i9VtRSgeAcXXjjhCUsHqGqMgtVCVjKzu6p2JWegdrrogkTJHFx1C1q44bybkq
rYzabFCPFlFtvDYWIhTU08yA+CPwyPZblc2SGFM4k9JndO6C3pkVYYb2yxeISNhpFjv/zu0D7Or/
3NU1M0dwPzA0Rt7G4oI+B0HUFP1e+Wsb6mR4AImx3duNtlkEc0/vyYiC4qn5LdPGkvyXkGXtLnY6
feaZ1yQwB/nv1Jn126q8A0m0roYvmqVLyDMjdQzGsWoN1+rGoFQ1EAfIhTtTtbGpQ8VZzZmtV8EG
xsbWCoKB289aibkqEXc7CbuucrL5V0RoCpYvT1ER2fiYPaMw7MANPaeyKDquksXxkTehW4rpLxHZ
621d8fu/hGNXOrXzcP1DnYT32hPJp2YRvENNCmvFxt9wOakHWndPwkFvlVzUQNG4iOwBSaGqZk9e
P462SJsXLGeNdu7u4skdMLy7CEcB8I6a+1IP6xV3Led6ET5Rjrz6mrFxQ0W6WifHufqmyz6ZEkA9
hSnxAp5ivAFPsIfxtLDMB19wt/OxRSp6hs8DJU47ncm53mkLl/L9AVyouBDl/TYtl78CSjCf8xy2
mAfFVf9o1TeoJLtBU4up6++35wiJXSVOypAy19XqgdY5pgBQxupPUNy/x6r2T/gws/kO9QVKgdoW
nmC4B/SR65Bo59jD2tf9Wqu2SFO2rCTGmxHCSYCZ481ecYeldWCzzAmzxrsFnGrHcgTFA/HIHvMB
QWvJRXdzXrt9zacktyxJo/r1k9o7YQx+YDgTHx+aUoupzHkSyasUwHwMM0gapcuWMe2KzpxYUgQY
Fpluee0xCAy1O/HNRaLHWtYZkZzrmH+mHL/m9UDBvuvKekAfKRCKb3n1p5WX4KqTN17x0IXwjE6s
v3R5vYWAUw0NB2R3+3datqhqaorIm0CLCbAwny9X4hrExgyYU1DToG14z0+Cf32suV7dXsSEZ12I
VaP3bRYn2yxOBTJNr12wsggtZCxLvUSM+CTgSGEzk1gPM721NzQKyZREUVDzNUSGdR2Id/89R3sP
vyGCxTEcUpg5/+n+jymvLDCR++xyMrjXpQq/X2Y1XmaJn5+auW4mgsFWEErEm6WJic6rOfxbZMyM
qyHVxunh9cByUxhs1knJ+ttqQGNUwn3HTnhq0cxv2Aj7dd9GSju5Xw9qdHitGYrlKzGGHNnm5T1F
HqwQnMjaPZd3z/HCvEAh57kF30TrGAV5C68bA/nfrwZbavE9ji9exsOlB2B3u38zfXNWDetrnHUL
XGqjjTkInm0lK0shFg49x5HnN39xPB+isZSOkhVHGr7bltWQxWJkAaIbUoB9GyzASXH1gX1DWyST
2lLsmL/jKtxqj6NLR0vfZHtVjFaexEZHIUMzUY1g9F3UT1ofULMp/RLoxVdoTqxiia5SRyObWSnq
1bgQYpu91Y+84zVq7VN9Tzd4ca5T4owCOvAAlbXfbQXAUXc1UNIfQJ/0EfBsBXSKWPLKnw9t2xzw
YnjmmcsbKAedFDkg2XrM2b+k30rggB0aTNysCApdyxphAa7gyIIwDKTks3+BMkCytCuqbmXWDTlp
Djy+r1kJwHbAiAkgtSA7PN5WFkx/8UM3opEJ61h8noUyUy9otN2Q2j+JOYwD1kkjPvoo45VRTnD/
lVP1zW2zwLPGKHvs8Fvb0z/s1CSf9A7OE6YFsAanQV5LYklfMahykSmxqCeYJv2WhKilSqvm92lh
D82gOtr/Hk0Pq44ioHZr3DCOTwWVddH197o6S1BvmrGjpCo3YIWhT13HjYq7XizWASbD4nTii2K9
GeZ0Vv6Vw5Za0cG+l2IRKdB/p2FNKFvjQ29fDr66UYFhHS9AiVhFqMOnn8UAzdIFAtcPS8KsvlmK
RDN8rJvhAHzM2XQF3QwFcCzjLXmkAugxvxg4oG6Bu97//V4mkpJJp/KWTwDSR94fIRIXvWekpIk3
OCSjE7ppYCRZZkCi/zs8xVmLGr6SHvk0JD7YTsDG9Z8WJDtVD5rPAY5IOJFFLk5bA/Ui3Nl6Qqor
5aSsg/+a3TabUjPZcp01eJmBU5KDtttfNwtpQuihJu1mrP9lx0iv7yilRzYH01Tv9MygnvI6d0SH
uNFXOoYX259HKv9nsS6w3/CUrG0bET1rmjxFaNvDrOAbLdvHbHxvrRt5t+i00cCXG46uAdHMhCzT
nKzNnc1tLG19EqUscaUIOPEIFEjfKcsJfVGI2h7nYBbgD5qDpRhzPiaYg/oDdfMFsHgaaujVmASz
ghjr4/XQAb1fhfJKwwhChyM+scQTpq94H4pyFaIs9vKGTGoHYCSuxD0dmDsuKQ1iDtOpjqf4C/fl
rTCC6sueAeAZ1ZlJ1TVcf5dCcC7rXYcfsXguTEdX0DiiC8Ny6zqOl8cm3YPaj0nlB4CG75dousZG
27/lc3em8JyH2V63msF9sFiYF1/JnlS/fsSdn+DjEKwbQVFGjpJ3BqA2AGeEGflhTCGg1DpbfveL
Meq85DIxZBKLtoNrX85Mo2EqRO/M4Opsole5q8sonm0NRKxqxQNRHFz8ODt+gws552C7qu+0zAvy
sNlewBRLhnI+ZM074Ru30NtrEzUBWCfxSnUwp1xCYWT17obIyRoSAjOds8TYpI3o2NjpIscF9mIH
BIj+KYvXKqMeuw3iRJ/OcQgVD0xajb70lt6tfL4weFxctrAiz7gY7qIjpu5+SdwEzcBkBpLY4Z3M
qIsxYDbg1IpCv3J+vP+XQTZrTkDC958R3hXm4yjDufYfkQ9PiPEFL8cuvNdbdOsDiNoPPmD2d6QF
ymyictJZNRt/8fRtBb4tNCovR+nKgqQ3Y+pCNYma31hy9VpQd3VFByGeJQwnFhxQMFdcATK/hhUi
ai5j5uLPKzeQ0DkKTXqR9rMOJn2HAAhBdDMxjPKPOeNZHXzVxGMVJ4eiTEPE/wRpYJRU7TVrIr2/
wDA7gjFFBzCJRXtA7e14PmkptXTlnmqBUoOYWdGR2vUovjY7FnfefLx5pZSYkJqlCuh6Ke7+3FpI
pdJ7jmWsNhvuAjMqv/GqKwWMBAxdxCIMlyV1JRKYJ6OYmONDC2H/BrgNW4uvKB8vCp07xT3w811r
zw2ntLdHmy6yKY8Y9XmbF1Z79t3u0xR6zXjNIb0Sls65Q8aAX1klvhZ0qt8cWydh1uvBn3nFx4cJ
iMVCq7y6vWkYobmYBDjN2B+ZI/HXW0Gu9JtKHjtCNlQrAtqYdSdDEg/IDkH76TVNWkaw+DeBeEfk
eT0U/RFy/2Nd/r10HiR8lR20CH6u7M3FeKNFWM81hF+MK4l0byVANYodKrjwujhx3TRBBFeaRDMn
bpmIKDCM79vfCW7aMpStY481b68G+UzI4LiaeGp2WA2GtJ3iCRGrfXkeQj2uRIwgi/WXhGiqBjS3
RLfBNFtTG6DUh8wsUhbQWir2Co0FAu7KddwQ1EAlsfcRI0+AZtlrEnBeo0KntPaZMG7PTBkppLlj
lFp9tm8uxR0+E4QMxNSmfUQfLJdTSxVsGyI+M+SlW3b6nEOy9+TJ0Tf3wKevz9+3hSbyQ6bCFj7w
st6mgOneOhSh6AL3p852OmQkPexhHthL87eaFEcCxGKJOMZej515wuQYFuEmXyWapPfkHVajyvUY
bmyCX+CG8D9p1RDPK+IVRQzcGFoCg2keuOMBRjxCRZqSyaoK26CRliersSwL8SgAQBZKXTGVBk4E
AkwVXlZjHLP5LC3gbuipDQA7ZyFvtBaRd06dmhgkPjddvExxQ5LgCDP47/qwNUKocvIYQ7dja3Fd
O11ymmLj3GwS7c8zW+eKssRD40ZrFS/F+HO8ENYZuJKMcVHqusBaQ8U2DEMmRFEX+57ATnOiR2il
qffiN7VvEqeTAZG5ypfIpkdK2MAZzlHkTlCksf0q6jl4cncBWX/hVqclu7mR0gqWRo/4NoPpD7F0
iNMlqWJlG799joNcunJra7a26gEwhJA/2mBEBCa3RZG99BLo71ie0yu10rFAve1AL93dKDV2bDgO
BqGvOi8tpLwbJvr+0Nw0zWmkWkms6G96a0ndjGQishMt0NrBTXRiW6RH9MlNJJKSfU09A+QK29bb
gAYDaA7iQgZ3Q5xsUh8VZDXeb+vMTTJB39eMjUmAHS58lzRp9yc4uJ0t8ZVAKzAUfcQc/OSeJI7N
Cw/KBaTwwBM6D/hRU0VXySQ2qkxMK6SEcjbNjc/drsoQLGR1WqAUeWBsP5nLf1cikn0q1NhkkEIk
r0aAiM8Yuvouw/H5KJSBLMn4o4VRiiwtcQ+ml69hC5wzIvijKmL15Wac2Ng0bKI9BGTRysk1cnTE
FqPH8GuM0jsatVWGa3xQIwIZJmH1/oaTkPQ/tqRhjH5HbRfR89yQXtTk4i/RwkpWS/6W7eMzuiBC
gmlbqc7m021Ifmb1uza9pepsD2YAYsnFlVmkB8dPg6oS2Dx8oz3JyI6r9gCtjXWEFPqXNETIvOo7
1xoZ3L+TPgbo8v2QhE4FFSubhkbqsRlZ+KpJTdXH1kPmQm/twE4LqzxzbWDnLh/EDD+H1OKmIruZ
C/r4VS9gaZWlT1ufbXtXlb6HhqExJzfpsxbwbJW5J1YpzVkCL7YCoNR7UCfUYl7t0ZQvFhwPmBSy
2PUnwt82zVQX/b0GlrcK6/DYzuBYwVkD/sE82+SooTEfDkPrhxEYax/ELb1nzOzIW8BN8sLo+HpX
CT4Y8FGaDrWdYPIdT17Ay4HP1pa4SSQCUqHNnEQduVZ0FEalOfZwkuzM2CvOAEf2daFLPkYvJuRB
U0fggg5IPIEuGKnVcPyXIlyTcwIQXJDQacnl/1DodPlt8rbdeSo8etQFwzdAKe+ZDE1HYsAnBNlL
9LJAAQCYIZfySDLLEoufZsvbFIf6hqP/6Qu81imIHwatcaMwfKIeWRv3gtP3AOlJDofjL5uzzaFo
K1u41+19BstLW0xbkBI9fXoUe3bsHw1CzR/KXochjTjYwNHGqEAhZQ5xoa3WE9qsabeN0GzndcwU
4M5NhQJBOFWiXpF1D1fvPW5I8ObIxVWDEFRBflbnxgsSQBTzhu0SRbhXTTJtCebJqpMlEpX0tdtz
VEvJ6zFXxtlhX7/lTa4bHdFatiGME3fC3W6yh7defIzS+0LXl0SRSn7LKsV8rELLl0dwhGoRfcPp
4b8t0WS6FtfWKAiM/toSooE85wezIOwBRiucjaTjg9tGZyewSopo7s1s10HmtrAqn5HWlfuQ52rV
vbU33TlqnCgKQHu2JprVYYiR4O9PVXX49gAe3GO4usnWqM3Msrczg+/amNVuIte7TeXZDOHr8IOy
PCKIOyk5gOYEG0vtzY6thx6xTU18rtZRy8oT+eiw62mVSzZpygPpPs+hSqtyrimnRIWpn3mC0KR7
Z+wD/Bz6x1i+GovCTwDUFVCYFWPcTTDTvPRN2lqzf333XpZcuMIxdrf8yxETjxAW7A4/OnmCFpGR
jHIvVBjM+fq0Qp8kSPWuheVD+wrZA9U+g3h1UIyJcErofYgL48AqTRNncFqlp5BbcEuYTimTqr9s
U8J70cTzij6DJadlrZW0PrEAo8YZtFov354nbD+Cxbt6mUhWR1+WUi0HmA/ibHFXdGgkf0PNnr3U
yxVsNnSdWly3lk/gSE5BxWxMLw0BP5YbQMv8vdBTtlA5pfqQrJQlwYu4R8gQFR+NKtAqbhdZFWvF
31kPZ+0mv/3qW8BHiv3Bwco98hHpIwwOOo52TkdGQcoWwqDE5Gsarti/7sdwl0Yq/Xrc2sX+ldU+
ZWPgGdREhFZa5Qc8I1o5cDiCcU4jK9lhhrBrU0sPN096vfdP0cr/ustTYQrHAf7mz/4pqWYzZ81P
C1OuuYhibTWRVCWPkPegfbPJgUSbs4SJa0OBVLnE2zHPNfFnqgXrinKXrPPN3gNViniqy3GrqGuN
5OvHOZC1AifDuL7T0pgbkH125HTfw5Diurhm9Y8CoYABsACsDeL6PB8mzgrWrg9MgG4UPovQH6No
f4vcwpE24oICazYF7vr7f/DBGmuz4+7HN9C/DaJ6En+LbuaPIevbM8+hEIGySuIt2/9abgPNM+bB
qKrz5weOHkUVm5MiIAsP+umGnHpxNediVx2A8DMn4buU93x1o80UW+tfhMgSJcZOkp1AWjHcASJs
WewX+ulfIMR2Hbuq/ByNyaVv9IF8+1/icK/yEmbOTstluEuIUN4iRQptlzxYAY6xoHHKWgNQGN8o
NLHXBOKd27rP+yYbXXgbKfbsXk+ny0Moo15Wp1BhUE9LLJEPu/9gJjvB+xInX8o2D0Tfc8wP3x4y
MAJfoDnl/oMmPymjmLpMznXxwLiiv39YA5I+eZV9OAtvsiK1g12qReGRZZNzJv0JdRiOt8fSWniC
KPSvDpjiJpz0EBkPf8m3SnCjzVDnW5c+LlBG3gIyotG2CnNvMzYIVa3ifysl7yuVm45+OJ3NLdQ6
OM8MhKkwpl6YMtYEOXCIwBnJCR60b395vKakmwbiixTatLpjGyefRySfZBmN/TlKbn0egJ4hecFl
Dsd4ZPoO8AO6ugnnTOr2BqysjOad7dwgocC7rQvTxqikhxVpIWBZQcB0rBD8S8/VmG0Mr73d5nPR
1+3oMDvFu+CvcV4LFDd82g59UG68TSRqXxsL+S1AgqQhRrXH0IoYJEcDOgFDh5PtOQuk72Ed5SZf
hg3M2gVJYp2DVy6sKyPE4TcH8YBsrFNVJcGS6nRA8MJxhQNlA5oanT8nbV8YRL+IYrdKDdNfNx4O
48UwOjdNAzSwxdXotLwFSvnzbwbmkkdPWZnaqwBo0fUMVtF9glupr4b14/bo/e80EL0tMLd14K0u
6++YxGqOrvrGVPdjVLf2H+0h7bhvuUBuEvAxHO2kQivQr01RuFRGRm5ufvGPMmIdmFSRRl07uTa3
uwk/ERa4GzuZMcjpLFE55q2Jl6jIVUlVu1c6xtDz0ETOrFqcWEGCSTdHNoOBlxOnlFe2PDZdWvqu
bVfGjZNrTrPrVQwOlse1Url+M7G92PGVu7HhFnkQ/hvot9FADQGAk51R2J7b+qaltivh7rRf5KTJ
yJ04ljRyVZYnlAzui82h+iF0xDCO4JvJ0tDNz0G1n0PYiX1N8HtLMGno0zifrwV+hGxISV+jSvYi
FmdDqRsTLqp75nky8uVfWnav/ll31GhPNkJMG0fAHPZji92ZYueHzp/eJTfA1iMbv2/wHu9AeRJz
sRu9r9c1bzSdnmm+PJ8Gn4fe/zeCCvDyjl34ZwYbP/bVsLx/ux6bc68oACBKl1/AeVCx+N84xt2B
Db9ZOHbm2hT67MxZ0zN+c4pDYufkMGY9u+4XlcMsXhEAS4mY0p6DW/KcAZrlEKwEYonYs+HLrC5F
QLqgk++upoUYJXALmSaEDZg9LmSdGRVAH6J9/+ix8Lwo+dDgkSjiTbiVTotCcoUchNgInbuQjj+D
OjflLf16SK8EcLEH1ghlTjHndHyIxKbDMmpQeJKQjg4tPmIXU1seS+B/4cpvtW8/hMrNwRa6AlKA
yWt31K09TvzsIdBspDwTSpnu27eCwbPA9tMfgGjWqa8jsbmnyprkmpVCyIjasLCW4Zwya8p1+xIj
OjVT4l1a8R3VCPxdXaHq9H8V+qtT1Mapm/kOD5Bu8BFgSqNRJWwkg4M884ABVRSzIdM0w9Jbnyl1
xWHVyGIP9D+5rQZ5dhA6UOezd727xzfkn6d1cpIVZqtSyBof9c7+ef3vgW2V/jh2fjpnnwJfnFrg
pooYtInCGk3UNeRi1PGgHUMCct4gVces5BlQmCGSG6qij2sHGfgti8op3NZsJnXEspS0awth1H/n
6XlefWmS43QGfNppcm6LcCNzNOs1rtVlkQoCxO71V8bO1Wk4ilqg5dCiCboM1TRd/ihDY4WnPHW9
pxrtUwt5Y9vlfmFfn44VS17BZ2FOjz71XvrbLpwTvjXrMHdGEmK4IioPl5lypeQY9gNdNN1Ko7zQ
CdNvDftG4R3Y48echGK8DA5sjtwhe4mdyHni62yw429x0eSMnB0sJ3M1jqLnB3p7UlAqcBHDm0W5
29h/B4Tr+oe/tuA3jHKiqWs67S5DW1NxSTPOM+MaizTY3mcF9OeAnQLWT0vUF0vYbjJ4kTjHv03y
9CcmI34eWuyj3x30PHJ2OXyV7vCan0oaLrn6aIBPIurkMtODW83apwjKbW/23M4XbDkyxSvpeZn7
fblpR+8tIg38EujZucBrY8Z5RA4UehbMOyNvc6uAlb5wKFDKxbET/p+9KsrsgBjCftFhO3hsqekW
66lHL+4JUnCpYzWlOMvgEKGDxaT9y9ehgiKQS/XNo5xccBCq8iVc/VYBV2vweAfyMkRyXqzpirUZ
ebD3GYqzgEqGY+6KfxLG0CgrH0pS2KN1m9XbRAhril/XU6waPjjUkqSPGORLOeGdM97sqfwuXwWC
qn0odAc0ApuoqGuoKjmQ3V8OxKUp3uP4Fu409jtAwHg62VR7ZcMJ9rduKv9wGdvF+oxMgZWgFE7p
lggGobUW4BebkW3GKk0UrhqHiwh4g+uSwX9Bn7Z1UqCnqhGSDoloIHwOYdYfSvoe6jCAAuh7mmhK
puB3Xr2oFyP/dTNyTHGjTTv6pKrFO3A7T/eLkJv3Jz3pHZxYWwOXDK389VTSlzf3nfF3+kj0ZAIG
Pbyk9LdBvPupciu3pSL3z/f7sj4gJub/Esf2Z5NHwnkSZlt4Wcccj71AllYPHvvEzTj00bN7qY0a
Nq+Iypp0rtPhIIfspsNcx09Z9NsZr73dRrpHn9hsNOMozbI2UD8A2m5s2yfaG9NhN+aR7JivJo1v
aJBogoKAILxjDuJsynsQQXOhUuin9Sp4EneBPbx2sIYRNcZAAZ3qyf/k4i4obxbayj65DCzI4TZ2
Z1LEWpbjJC5wdPHWpG+Po8npF0vhI6ndD7b3C38y3kYf2KSpyqV29yJ+BKu4Qx7IZ9VpWEny/hHN
z0iqj5gdJ0l7JYlGGzHPStXxUqLL0S7aIHkGuETNiwjKDyv8hNj72wTe48RF9UFvbO0OwNs2NR1u
l0cwHdXCa2WnP98MeO8vq0FuWg4Vaa4+aCROAd+TSBilwW9aZfrlLktBoOeiJb6stsxRrusECIkW
MecA4i+SWlEgIGM8Xc9ITqwYydE62peePhZX9W+Nmlc1RdJ5QGCfNyRWkizUFDbRs2XDUzovGmiG
JUHojF3Tp11hUzto3F5CEzlMaVL47en+CcoPyzx/W5cKzhXr0q5La2OOQnZPUB1/Bbt7dQia0/Nn
RqxK/f0o2dHq+cxw0TN5X6H6q0IArKWEHTQ2aZlJKwsSfmkL08ktFpUQEMAecwWeQVsGzetafEiV
4ByX41O14hI9//+EVbIJf1ajoXqAJhur/CrF0wlT9HMvUeRi+vKR0cdyE0celsMDvH8iZjRfG0LU
yu9f29fUxWueoA29ysos3S1pxY19ZFnffPXTUIRBMYUyp7RZ5z117KavmIocx00qYQcahwsVisKU
+d2U6tC2qTgQIt/l3BZ3ElUla2tSDyRutughgnOCT4FUlrCS4JTW5wZkJb2e0x6MxGXUDcLvlRgt
zd8LVXeJVSSQGJIvvTiAbubAIk1HlhGaEqP8HXk0z7WSWCb1CwCw1VwKj97EWdSeB9KzJWbRRprz
6t0uf9+8ZWQ4ODju51NBzGHLcoKgQitQkjM7uLpb6sQcgAs77EWxVpMXablhfdmjkzm1BOqSwTmC
MZgZMfCkd3Fw8u31uoCuyDvbNqYlBcYP+0NVATwBbCwSxMGzKCIj21Qmo5vJUtjSu5QchNVx9/0w
lGuqWukfEJZFdSgn4NmLsB6VpxmQbLDSfOGUAVyvQZfwRrQ7L2qfLDAfSpS0p+/ZA2EI5PFei/h2
2oWR3sBK0eXCcrJQFQIQLnmnlN9rKGh5Tn327VRj9BERBw/KwMfNEH+OdnznZAFVYr/5Y9NkrYd2
2k3rg6bzLd2nyWKc1HyLdcTRzp+BRyMuy308WlUt5KyTKuAAcHKmhdkH2KZ1rD2rfQIr3XMA2cMk
s/XjzCCkpFCVXSaRCPZngsVKK0Y9dTzXSrOW/m65tCkkBQQl4GIhBBWCF4dv9teaNCm/uZ8gO8hh
9uI9BO32hSo4zTb6akbzu2dTTE+3nrFaLz3FKYkqKtpm8DT1FlSuvICubIUHOVycKIjDPtn0esli
WwyyXniBElUPG0pAQh5ets4BJXc57N+/0bW8L+a23Pr8EAquAxzHmz/AEMzr7YkKvkXwiGlY+xni
1q34V7fvif1+Z/kQOjGOVW0OjhVNqglrnSR5wGdgC+KUpolHa/pztunTeaNBtC/BovgN1Q/qrjNl
uNgh8qrxLo6iZGupKKKR7FJ8aPH4Xd/9OvFZUEvdcnnKubx7Zs4sPHHxr5etmv1/7ZrmOJhtkTu+
tjRBWWXCH3FBI9wYNBNnZGhgdmft5tQ98+QZ9OF5HE8OlWzEM/ENTxGy/9Hgu5oNlpG8qneUY3yx
ZPDVToJJJsMYb4hPAiO18V671lorgBCGh+7tdZWT9g2OTkDCNcyujrZ5QlB0//dvDdI2cJJ1J+ol
srwpl5choZqX3hznwXCXOzZee0SIPBWS2tf2yS4R0A8PwhKa6uK37gJ35XjckNe3zhwTMtP1le9/
h/OiOy7kfp5m2felKIXf7UtnTAIzibDasEvH2uIp6bUj/ktQYcgALbx7b6g3420AscSBPoyVeeB4
CVcWnImXWfsPhfAGzxHrI8wesbBxhpmo9KXNMMNjTB25JIK6nEBIeZxhhR4velwJkYtcB5SFnGZI
kBD37ILWPn0ol6cSHFNBI0GhqB1PBM2uPe5lohcU1zSWUEOqW35R9zwPrYCFi3uJ/MUM9XRy/DVy
tZUvrYH1szGHycWwKS9CmdGtQvQ7CrdsUIHtf7FJRvmSkdk4MPbGn+t2o8REZP4Mrdk7aF1Zwetf
Inhw81Y4Xv/J7Y086p9hW3hw+M8Qla0g112uCRaFQb4hRoF5RFStl/pvRmQ14ZiHrChFr0v2yyYy
2u9oe4Ao0P6ORHmB71on+5FjAZSed7lPy/9Y9Cc2t3yCt1v0Pks2rIvImgTSkpRsgRYQ/x9x87N0
W5Uz6wtzqrQAfG5eC5NU619QkyVNUslVYcIccNsS9QoXW6i0e0nkSvmRbBP2EqXdpkd9udndHWCM
WpFlzN+FxGHt89hpTntvO/tvFbLww0MJdjMk5OtTi1K0J0Zu5eMYFwWQs2q7/m7OPtKZKZjYGy5J
Z/vjwjh44+GwHI3Osmh3huIkee8NVnQzy+BMm+2DcCEQh/a/wXmFMTwrYhFSKaUQMH1e+sLlDu3p
MrRrma/o02ZjHlfM0QjLywVQ7s1IJMH0ec7x2hPPDdVVevsVfyFroG2m3yUcEFcJdoUV2GsfYGMa
nxZwxn6Qo2V1QukCDqcQjuEFnPT6xsh1mik4GTpNp1DHj3sbIDWu3ebQIyxSpT5md7C93MkrkrS+
6EMRo4hLCp9TbkWw0SO73SjppTOx3y17lelTkOozhc3uxEB+esa1NgsQK0g+rZb0cogp7nZPsfhA
5LfXeSyXBmXmZcaaZLuCJZTAnbK+A1mzwnIdOybt7mCRka+qtCJL+/W/v7FU/KMfOTUulA7bWOC6
6BlHUcyL1+faFNfU76+lxyktDRd5aGOlq29rG6hmNbzyfyZgbal/VQ9P92ZoxVE6L69CaNvtBD42
es+0591EyTdlVbER2t0GgPx7swvfvinRZ1KbukiqdpLmDGxQhm2ORiMGv459cSqkfNviE5xP8jhc
pB/sDY76HWoqj3ILaiJpfXppDvaaOBJ6CvG2xDpaaVi4zBYFTf5bVtBhAeB/mUcdK+CTxDq25CGg
iF9z9coW4Z2QSgIgtdyihlRllYjeQCN9gtT5X2yEwA6BVq6P2+Ceu6w01T9+qbLm3FVhoWQWN0BA
lKhcWMP2HkVUvL5dcPHeQEFqZZ3nNfTJQvbmEMlXRMa433NNggulfqiidhHAXzhq2EZPBM9YHjfW
FmBt6/sOch4gN3zD4rXXKSDR8B3acelYXw5Mi55OD0BUlH1h7UvtZvZ4rMOPLK1QaTM/RLcinGQc
MFt+YBVeoih3QV2OpHOMOjU9GWGi8kDgJS98eD69YkU30Welf4N1in+1sKeaD8RiWTxpgF3XbWNb
q7oXonFovl0z1r53Von/BO/96qiS5QopInKJIQvvcC/YT/Fm1nQ3+jGlSMn8RkPCIOTviOm97gqr
/qADqXr4+x9Z2YxCo86O4MDoE2EX6X3EWkVVJkYliSaXec53uH3x23ywkakmqBHbLFNZfo5AoFQR
YZQlFs5fYD2JubaJ8pmYoJbzUetiYFMxDUbcidFDqssOV9idbpbb0fMTOwkGHPmkDg8iJ5hCTWO0
Oow4Z0WGvhYBYsEQIlFFILkrKXqV37wStnYSTNLfXr7wLPf/kWen6BvaElFTly60R2DBDW7r3R89
Nvt/UdtZy1mW3RZgXMBY4LcRrPcQd9bRiqYmXOme0WxCncgn7CGgaU52Maz/IeBQdjNLM6LLPb3u
PkuQjiZMtS1IBsQZbWCAThIepuntdOOLdShjGODzQ+ITshjlRDowwM3q5iwYsHf0q/gzbw1t42nh
p3RRvrhPg/iamEK77HNL8OMOXDMDPo4zK110LB58rBQFF6mVqGceaJyrHkfS6X+y0mwxH7nRlaH/
EvNXFN78IQUWMHOupuhQ8WrjTWzi1IPhhklTvNE9FFY7GSfeReeD6CFgFcPL1VVp643/XTotwNMk
PYvNSml+A84veO7AWu2O16h1hFeVlgs2bm1zzwVCqJ6nVZak2iiOmnNhhbeVzV5th+uKiEgNLKrk
cVZyICnm5ww77UpoH6MxeqS753GjOPGN5cENDHJ8e9+ShlG/6M9pYR9iWbkkccyCy3RkUruYQ7i8
EVTB0n4D7u79uqgYis0P3/yIszZV4B5ZgTUIoD2rfUnL+f3SaDNyFGuSyEgZwe4ZpdOBuEXTcIMh
DAWlJO94+Q4APTKAlEQhm1qb+tjlyaoGG0nwz9LGmTr//+MtFD08gcHWaHmi0y3E61c9jA830pd+
QzW5WjOZuf+NFVWm0OmstJNFRa5tE6Q46LRV/JQ3Z/4wzb+j5RfkZBMIC8PGOQ4DtSdOXCMIjmrm
zBTx0oEObAPJlgrN03Z3/XvgfB8tEEpzfB84fIOnw4nTkUC6uXiItFoYBiNK7banqtnf8ehKdgoY
3JwV3NOSNd0TjrZN5l9+h2NUhHsubbWuDm4Z7azLJNCjG6QirScu86j/33daXEtJJ3D1WkuMqpVJ
K3gEcRAcQDr81MHdDsGuqswTpRSKSinYLJ/FpQFe9zE3sO7iLNWZxoJmd4pnxQpj/YpPdcINa1Wt
FfEgfPGSJLVyj+4gAp0xS8vHzxZPnnWxvY+UQVgM+SrimH6fo4M3NpGclPFnhwNqImRPiD7kAK86
MP21R5CRzioQBrz1fi1WfAbHwsKY9dmWcCXlKgzFRxDtFzSD36RVagnQ9Hzmn2Q3Q+WSNj2Eb1sa
LRdyFJtXgaSPWEuw8xz4EJfZtBhwZYvrCAmt3oS8APRWOauqql4cdOpZFh8o+jGL6OLW7lm/5sUr
vrE3tAzhln420EsDUhVNDRQg/Mwevbd2PQa3iCkyiqLV069EXXcrojbue7p/JaU14LTzRcDk79sm
LzkteQjRR+kk1E+ed5crjDmy4fAJ6o2pH8TyArVbf4OXxk623CnEdfsGuY3mxnYZNrScUoDqDmig
fVb6uWVoSps2aza64nP2AymJpBa4SpNT/tIaFy0RAVboWSOI6Y7CRrK/AFkLTioY3BBTfZ+JHoIS
Onejr47rjeO2HqzTFwk4ESCSPpjzchRCbnHccpqNqMBCXvWE9+EvTa2fkBqF/7fHt35CmQG9BRAL
YkjStceAaF/XYMAx/NKzZ2g2g0tP1xfdIwAb5QngTHngjocQ4ksBPeYtLTrvcUxJ0M36fGMvW0+R
W/dAAQOZGF5c/htWerGdzXkF1CBGrchYRjZ6ZOjEKyANVmdz7H4/3dU46A8yiN1X4bCQZdCE8dXo
xvARv3OVnhM8wqgsKmC0kmfqAJ9H71YwU0p9Y9Kph24CJbYo0uJzi+hcNb5BW6wmyNGJo7t6Bi6+
PJguLTVJ0pPEUkM1lH3MN2e5TyJAMiXJevNEhIeAXkQBcKKtTfMEF7IcAQAd0u9pbGNYY1zDxe3s
BIcT9uDEXw0H/h8RyBHXGtzT+v/zjQbpajd/4jyQVh9YwqoZhoHs1WJ00Ozh1wX61cj9xFtRjZvQ
0Mzd1r6BM/GVTbd6r2qU2Y28O7TaZ3s8uab0j/gtcnUCFpFsW+LZP9x90Zr4MXLB128gcRXkPLfB
D9DSpxl947aG1kME8u/I3UwJmzoB6G6Y/iX71iE4Apf6T7gSxgx/nCZ84n72Zji3I9yuwU+jH9R+
MHT+YtXMwfwVk3Ozk/EAsrE1oj5mw1gVvPWHpOd0GEJ98M1N3zCYZj3cbFxHGPhHlE74n8+FSn4v
XZ4gNv4pbMZPtI61JLp6CUk0S97niXg7rcu9x/tTrK1Rv4bF8hLMeytz9zNn5QPH0MdgnTjz1mrU
8g0SGKlvvQPzVsSHuBEocRSEXOppAwuVpr4lx7YjOTZVbneW7SsJJzAIraOqokLgUPxDffPGoMPX
RYNRv2Vgn4+khAspvXqOm7lgt6EK4Emv1X6RzmnAHq+7qOxSRdbmgcmY7AFKcFTZaaMViffJoK5S
0E1IR6jWszvM3dG1L+alo/gwnqgQLvkX5G0CBv9ImqFnYaq4JLbws2g33GeQ0C9Dbw7XvsriCLy9
MHYtV7bQ0zUqChAcNSK1QQ2FZR/eZM8tSBkyd9OqSPWrpnWIiUuuKHce350ly/zYPj24ofgfJM34
Z1N0MK+jGUOw6wWUznW/eZrRTRar20pj72WTHiSZgigYpUDjm243qPfqR6vZBckIZIXwYcqhE2++
+ILz0fj4CbYalEnM+OBE95tu76ZQJWT0K2RYXFwa8se+k375I6QoeICFC+JqhI3a/o70YFJaOESK
pWB21+sOIZksnCS1MXdmnq14zqvHIZLeliZIvnbuEMR1+MSx29q3RwyVe/ZJMId3YPWvv/8DVvrx
1wY3s7qRe91OBl+IUi8rkTNyO2mc1ZDQpcYmY1h5RtuwspiAPy2M575o/nrZ4MRwrr/srm7yXgLo
qAh/Nf0v49JkRG7zWtnIprp0RNsHs7rmFiqfPLaE6Ahot97qmjmvwLy8Qtmbv/OxNle7QGLz0qHp
rUHjXu5fciqXUd2MFCMEkVjGKvIbC/gio2cw0pzI6sqitZlLUC9m8p1jBNPmiZLBY6MtFGzMSsll
FJpQ8+1+aA3P6ldFulkOUueyrHE1DKtoqzPnVTF427raNtijLYIRWLbFRW5sQMeSUH6O2lyC0jWj
HFSYvsW9uALYZXbnk/mqvd4OuPCfHriC9Z7FUcUyBEGHwgVTQ1QFmBoHLJZjlMt/nhJna08D6ZW3
Gte03VvTFi1j+ltlrsvsbjuzSWjA9IpySMZCiH/og+3ueVLUzJGRXxgwhFCfLwepIvjUc9A65/00
AEj+qb/oipTBZKYAOG4KTxS5WiAPpqGT0/C9n8UPFjiWpHvZ8X0vThJYtd7IN7hHuugyz9oM5Whv
LW87pSFj/3bucDpFN0pPv0wbp87znBe1BCdT5lEaxhNYEr99l6QP/slnY9U0jlPQ5iW0Y9kdRMCx
eGB2oGpKhu8gG7ABjbiWiROWLtyFYqJLunu2pjzlwRHagOMoklf424CI0M4asgzbQguo+DRybaYh
VqETL0qq+SC4kPe1xpfD6DUa1OjntXuDFjyIlOMzyx+bJgVPS09OkH9dIVNEJact1EpzY7fy61/u
WqyXfl+meeMtRMUfTxUbTiUG5a7rZq3xlPb6EhVygP0btiYTj8MNH4AGkiLFBuOeKc9cii8bkDbF
KJnN0I1fFvQJZ96jaOHlMjbBvYCDEOaLDgf96bQU1ZOYABgHd/nS7ON2XHv9rovf5jBCzICQ11a9
a0gDCrV9NL8hGtdbxp9tb+/C9xVoTZaYpe7cXxkX8kMxEHrPWvAssCzmBIiY5SEBMYCd03brttWm
oa8r+3u7uvDhjPXBfFiMuEQQUXWsFjo9S4nW+e0+ZvojFd2DJUr28Sbm7kEbAYhgBmpKhuu5rNh5
B/muZhG63B0MuJz+NXwqKiObhXNZkR2a1AsmiPRkwbrve0rSDPM42PUKOrXdPMwjjG8Sy2DpT5QO
U9ynLAzBpMX+PDLsYaFMQbguKvfmMVWDPVrN1Ru0GANhxhmnC84sm1EsQsfZOAc+z/trgHMvMy3X
yg5BAUjQjY0OyDIz4WKzUixHAwSIy2zX7ebF17KSFLk+Vp25Kgh3EYoFlqjtktHCF/6ESg/DYzUd
NnCaS5LR+NA0bLiGHon/qm1rzV8S+e0QqeuzlK9O7Uxe4ZKeUy0k0VAkl43Ad0eZV3hktZS2seM1
dXlGAhdlNI9PeUWvUAJZd6DGmNlemIUCgnsxOv93lkh548HZoVMoDiu00HXPPD4gtWRDUeBg1atw
KkA7Ysl01eqaUA99Vg+5FSNbVXG351M1BnQqkz54lBPVLOlKlg7Ngo/+psvlWWlVModzUGcmtqi/
GCJvfgFFGZCZyBxI7nxGsf7eItHcM8/eTqrGfq2H7RQ2/kFDebqHFs3ahWzSG4IsoF6zU8sLBIDv
UzKFoscjOoVo0sGAk7CN/1MkZgBLZJ794X8TmScf0VKcpFIxBsKH4WS94/rREEYaORQxXS4KjiH7
7sElMYy45RkNTm+GIV27+fX7uW00u85l/VVrSd4QIG7q/jSKO9nWO+J1n46Wr7B5+Y2akIhc6BgG
7lWi+Tt6bCs+dcNgw/xHha3rw8mEN1dWVzYDIVIgBP8ya004s6xm26h4rVBHc5W2vYCYNrPjpZd7
XB7LccT0hHFXQZVqO2laphdzgVjwy3k3zWTcgsAO1wl/m911IYsOyr89xnAtSPnnudsWwANHFhnP
qtOBDAqDch4QYs/AjzBmV2m0ovgCAZwP6MkKzfIwWU6xBWzqU5U6f58lKOFx4YkIg5APxXUi0ml1
9nK5OMggf6gcrawyQZHNKxExeq01Aoi6B2oEdP3iXpcRavWEtSIWQAwDMOv6yzQ8Tk7tXpsw6mm9
LQ5TWUck8VOiv6EXd0jIUSAl4XksnLgNCkAIH4zfCfsNxn+nLAMmrMaS9tbsWGs05DXMUf8GePrv
wQR4vJiweJ0E0KJDEGDCDOyBHmGs1c76h2d1gXqJjxY0aoX12mxp0pbb4KcCOjuUtz8knPcnFWkb
+jf0Z54NqQVKczNS7w4vK8mR15hAaqv/IPNQKYn+iQMB62HtNoNbNiQ/vNOWhfQkBqSwdgPmrLZI
5NUkaNi0z/nC8Lj+oV2n8gDr99MrRGGeb0Kj4YQcN2FPNLb5WUFiOtYIciIDuaq1s9uCC04drLyg
Kv+StkMbfqPHTaEpMm3kqxwLrTJMkrUX/iqVyQHinQ1YK56aCEt2mLWU16h18EKUu6hM/sZKayxc
/RicszXXiicUB1+RBobfrJyyCObaAZahSXAQlHbhuuCEq40J3u8ngRh4v6XPBgRjXFd4GIeoJVaB
ULW0wz8vhrrclIO9i0NPKLfU99dp90ktNSP43UGakiuNkG/KApB7R4stt0TwbdqtvY+1ATR99ZDA
8VeFkoesTr/M9xkQmNb3pT+DpgIbb7kU3Wgg1n38sm91KyFGezN8isJcvR0xZYd5v2YJknlUOlY/
Su9Y3jkC8bCMcDuKnf5f+nKKXGhy8eKwF0XOy+cIJT/+CCtljfK6ebMNrpYHJ9aAx05Ycy2UlUVe
O8mXYzHSVRJOWlATvu6EKIJaLJ5cFhwt1MlwZeofo+XlYb7Cdj4a8dpLtZOCYoKnBJNNjBu/+YRW
w1RZPc6x/W4pfrHQpqdbx0StJqxyfdkZ90doScbXnFfBj4OWmUkMbmBlSaD9bB8C0AHnmH6ejh4v
7Hzn0/8nbOYwfiELxNQrTSR8w2+K+e55uZZB81NnPxt2TGZ7giaVrhHwUTHJS6/K24t4LZJ0tVqW
jMBmIybjTPHkJbwEzBUcdtzcOGAh4pHLClIzhrofGau+vyPLnDmTrEuBZ+gbddFTrVNLUskjswMo
xif7rL0bu6RtPhQfkc2lYYZo4rIEK21vAx6Q85Atj1//nTwdiz/z5Z4jqnzwtBvAM+bVTlsSJgdU
tOZKOnW4QZzktErlAMSUgqVvNAOLmQk/Nj8AJwLeEvYCFARelVqM81eguvyhm3u5ztV7Ytf4uOf3
9fS9IMbdDYTatVkmFOneJ3l8ozPgq6MEs+GyedYimfbrjNrDdkCv7PQxTkNQrPfFPqif2HZ/qXJw
gFqqMvDgpaprh5uViPQmzDqksSe2arQHDKijgyi3ftUBwAHi+AL/tpW1Oz1VilvbB1PJzMaOChpS
wdhNUXh724uxNlFzEK33MfX+uvg6XbzKhi7zvpKe4FjRTdDi6c9SRErAvvB36TpIAqbcZzzobVyI
KsMxPRhPjhKI5sZCM0CU/+cGnl5xIClXYPSY5wqRfONwLuFgTeU4fl4tEM8hTxdZ3QEgu7al/qQm
Jis/4poymvPClhjFS6Bik9RCe1nFh0fLCSH884MFe4rfqnJExlfwCj75WiCA263wvagsOEyTwI6n
7+EDzWly9vmR8vKZarFRBfRAr2Rh0bHVX7oRrxy7pfo6cTV285COtGEUGXxdugQrdscg3SqShCDP
X6y3ba3o9PgAMAC7Ytbc1b1DjWj85RkdZdv2MUjNR2oeoDdilX2yRqfi0TDIip4YTI/NWmEJWwIN
X6A3xP8Ux86OApom0T7kCJUhIt5HPkFAI1BiPS/rL5fLdYNFjv7wzckOg9wLGZGPtM7Uuck4miVa
d4mP9ywHtvVfJ24wxYCEPd22vJiLStC10G5P2XsyZU7L/E6ovach4iO5CKvhX6IqdaDkpncSgoIa
DqY34Z0yoDe3qS2OeQDlTbUd5uIdanD/7UaSq8ChSax4cNuW8BR12MaBdvt3QwlQJkeLCLw2XOWj
wB/leBHBy6qB9KT1uh5CDX4QGaoqD3UjvbTFvE8VAh9nNKHLauO8D60ERzHVUYxpviDcIGce+WY9
S/HKxTTYM8Y9JbRTJw0Syu5xtXzoSFZhFBxza9iiYtN4Wq/27341YDwWPDmuDMwe3+R8CMtEtRaK
CdNhZ1wA9YpA6aalyP2PtVqJsVFwO3PbY1jBgUo5vpvmztsarhPjF10Ot4nJ70wQfYy1TSHX1BfP
T2StCdWC5nOGPEEKF0X0sZ/0K1H27MsSxf+6wFg5pLckGolr3SEiASLIpytM8/a4T957NoF+m+KQ
47EahskHRE5Cr5Y4mSkeCNZ4UDQQ9n4CysuDhcgcsnXRmTcQoz6fTrJNGDd/tOtotY08C2jTArzb
rO0krCqSPaQAE1aepVZN4dEhwd9eRecQBg7kwBS8o3byrXxYH7zn6d/CDSmmZEO6MJ+Qmg+C8Gs3
/41yih/OgRljGOJVP5JBnmzL5hl6UTA33dGXmD7mSJEg5Fopt58RDK3VGy2Gv4fErOGmr1TJCSJq
kSZJW2+wLJUxkDVGSZ+DJSFrkBSDCSyD+sJxkcXWhWLWJHiUuX0AoYi1CNkkv+kr0C1Fb/tZ4z4i
+dbSZv+pJ6ZHT3pymipBCaMWBmUHEyrovCOBldFHo1da7miclkWNeR2G1wNX0m8eWozH3DAwySs6
/4FXuApxx7fTppXvft9niTwWGzrB/yLJMnTFmGDvorF/4hWRD3KTkBkTdplv0mWEE/drPRDAwRpA
mHcYLl+qZCSTK1W7v8KCa7WwBsTIcVQrpKgEXPgIqD1j0rF+l/GdDBOR4+SeFDomM9bdgC/seN43
GJiTe4QL/TCXybCADE0oEAXgyUR0ecAQPq8L7gzss5v8C4KvDcscZyI/JGxSSvtZgcmfsVbYeE/O
W6AcT48WrQAxpmESgqEPhVpvxlL6/eEKTFYtqCvPZoZnTw4bXRznxw4mvrLI8RauOWZ0WmlVpiXc
dnMexp7mU3wuNhT5Ak7IrhOAOJlphUJig2bFqPzm4bG7ElRjuKhNv9vYu0IaSVs86xCYhT5+T1O3
GYOZtHVY29R2JGBT0LrXHz5BmUEYsIC1g1f2D0YoJ0srBhY+QukJVDVNCCn9VvW0SUs5a3liheoY
vn/bVAKktq0sAYQ1Y5+YSJd+7ZkAtxnO9qlyffDD+9lhIUG3IgbOcHOIYPPpcNUDTQnGnkqkls7n
vBWhLeyz0MXHcTaLW+McuMOOkStvrSn3DBp8DoYOEMByCySdr7xoVAh4Pr8TYgEOLXrAlIxU1QOr
4ze9hP4q+0Q9WsPsn58OdXg2FBac/xJFY+A1UTR4hPx8BGbZsNviiyGfCxstFdqycRd3vw/hfWpU
Qn+DRWrXMv26jkm/10qDRYk1BG/IJAdHX9oDZejqkg906kQEtuxuka38OqiasLGLirdpbG0gZzKN
AP4YrlAIF5IcWmu9yoTqwb6KBNaNC8MPkA29ubG2WlqF2VynLRS6+8PjcfhUCTP4utSihgtXyWiA
GuVWX1n/TvdhTbLKqlTYcHLPK7V51Og7ObWHTFkaowM8iXiXmxKq36Nwj/+Nq6pt8sdQ77sGpmCB
bXeqiXLIAKMF7Fz0/Xi6dP3J5yLVk4CW56uqkX5GUzVpxRy8FkQ2DAHRSzrohP4m9TfDDvC7ijUP
KoefuC7xguPPMFOfpnSpQNp3UF0qx+UGbTXZHNogyHpKI/slzbXvnY6hmLbW6e7F+mvPyYuID5PX
FJ4d6BDPMcpaDFULh3UWzTw0L6uCzbxiPHZ7cfIisGHQ5yPJ9GgBMNPnmI2ZuU9pea3Ulkiddmnb
5sdquA8Ezzv7xn42o4KFbKBpGcgNzbz+Tn0b69wCbMbVXmVE04UGlOtEKPuJ4mxNbJTrohokfW2E
pJ3UIgVpBh1ZyNlnVm6UCMTWU++g1YHEf+e08bL+UiDSTw6OWOJMDIipRRr4D6LnNkskXPQ+iSQn
k1u08eO+zaGvd+APq4lcKowqBC8nQqNt+bHQ6qQnaq5BWQF/zjknHPNzhCCEESjwHPayLU4ebr51
mAvMiPxSYw/idzaH4tSsTjzxLs+v+C2sJWC/3Zx7v5EE6/kmApFRNPnmnqbAARq3SEJB/7fmy6aO
YQJZ7JmAT++Bpx2sZPXknsqrs/1sbnClzEW+qq4j0Fa7p9AlbkwpN5zF+GVC3zBs+4PGH5Z84qxC
ThhytcA7IP7kqBJdvS9A1py+LV4jCjCM3CEYk5ru47C7ny5Yc1kG9OIjF17XuDWqU2eYaRMo4/Xe
5e0He1LUKWxGYqB+gGTTtd5W5QDbZ236EHjBV0lmpoJ9HaAbCBzIMxA6c2cvbzSvRYjHQi5NmJV2
fwvrF/B1XTkqoFrezadIi82pSsIRF7L/DKrWpdrLDl/OudwvEDXuwsqr65ttwDuq7i0ILUkiC7m3
unIb6/MC6y7owWXtExkDZq0qWVqaVcv8nkX4A6QwipfRxLOetkDhgxiSKjqsiCemWYXosgddQFMA
9h8XMhljNpzRFrX9ds5J1Mn5DkavCjwhdbVNZHanxQNmAwdvAoRmT9JB3XO+mnAowz1VQFYflHwm
xprS6kvWsDjfSvjriWGYLdVlvLQCeLb1ipFbPgEvoQUini4GdvMc1eCf1EVgF2Yv/UPg9IMON39E
F3zduf674YMnCmhl/eMwLVl8eeg3eZxJShrTpOK3BnKT9N6/YhhkWLyYGHJ3hIQ+gsxL4faTHY7i
mSyIm+VkUUNhrI/gdQ0TCzWcUrbKvbGd6GZ+VBLycPzb2g9LSRmGnApymF5oRr/ULYs5icHadbmX
bvoYI4fgz4VfYWn41DfAiMCryTTyU/CTh9tBOqzzGRGQ2+g4fh4bkVaKEmNf0png21AqviUSc8vj
BnVilVAJGfbmlFLXeHF3VzX5sKhJmQibPXnRoOelCuRYCSSdMEHFbPIg7XTZiEeOWc4jBImRiYri
YktQzgK/Ui6s7U8CTVetytQPfCaFmDj59RhEcnUxbecKYqa7GFr+qGtDlAYDICHO06SoQYJs8wY4
AORoMWqm3ueF07AGzQeQuXMCG/f4Jj9I7QZboO7/oQFqBGeD/y4VT00eam73WLa6pIhsFiWGkTUD
DuQSebtbCbYeoByk0VMsGAHHpcVzX3TriHiic6KrKoX19ubxHJCGGhYuKPuf6ksBo9baP2yuhWPK
ZiCmkXXHHPYvsjLAP7xl+cl2X4LnwkBzdf0wfkZ80q42Vb+MoERufV1to7PG4yZ6Cg+x4x3WfJ3D
f7E7vpERbHRU4g0kY4M99WOhkpCTYhpebPXmbuydJ9N5xW2rru1EIR9NjkZY6TjP9PtnkSqitJHk
UIEyZ54eBkk0wscO3FcOAotprmemPglhuJ0rhtscsW4s7OMLCIZQ5jO1eeD/lO9d3mR7UXTrFi8T
98BfOPpBax2djpJpWeSQqUGjqxO/h0pzRhWNn7W+B8Iy6DPIkehd3QaS2d/DQihU2Qv/bOMU/vrL
j3M4617GJ5eH7jzV/ifJYUYF7O6y6t1Y8XsHKsJQ56UuKWMQFPhwYO5HgkvK8wrDHEwfvC8di92H
jNFVu4diPyp04LhmeNPPzLxQnRFZWptQ+speSvPuVWIpkxNnpQJbepIqO4GpZep4VBkv07zuNUQo
lAocvzKtY+tEBlRIhkNcKkGtgE8PQh22qLK2wKXSCG4mrkw5W8qGSb32Agasmv8rYFvHQFLueDkP
gKDsn8o5eoqUhRSXK4/gOpA81GGk7HNDsBg/S7BbA/CppsKCd+OqsH7kKb87nrTdYrYGgmvuNOfT
6CgzZ5YZImbPoe6Y2/LcBD7Xa8WzmvwH7uty/eO1DLx7sff5gDYAMJyrwFAWZ3WAbgfiyHwafvxQ
skciatUz6+0SOHLblUtHqI63QV4g9QWOGHxqZ9AHctHuaA/hBx0ynr8/vihtJVM2F++I02fr7Izf
XzX2jD5lQs9zpJas2xnzZ3L3vBFeEZ190VTLaYoH2G5MAPV7QlNJKAjxJeVne6ywjUcF/fzTPD20
kOfdxJOPQKfseVHqBwASvBTb3UlJJy2nGAMhKitrEj1ZTqMEBqWBWzmL7OFL0Eyh1VFqKRPk4wMV
lKgr9m36sAbtbBOc2/heJE+tb6aUBZTSx2zwRgm6wJxtHwYwQ6z92t9mU0c/xQqT36wGVEw6qRjL
6mSTvGeO0kedRN0PB7XPhyaMHZsgEbpqigtxBDhB6FoiJENxtqGUl2U24EzFzCQSXBDqES6pzKeS
lvVqm5ZdWRLB8lccE8exXvhNEpAKb523Ntdqxattpl8+whyP3j/8xTLpe/StdCikPpg7N5mVh04D
G+Dpl84d6jQ28TQ1Vp8kbyjAwF3snD7jVcDECf9I4TxWFLAZBL7LSDMGbbTeeq28MBC2rHmrB8ZH
Des1cO9CZ7gsxClvqlyIpPDomBiHFRuFQhpPCcwFgIWUOc5hos6UTER/oQjuZYxTwGtKwmz/CfSC
+M12OEnyVVe8Ak/z9MMSowYD7GHRiGJDwrGTLb1A7+z3QhLxxFWFtIgZUjRIuY0bDyR7Z7w28RH2
BEk5n/BzE+R7QnB8fR2xSjpDhon7LWfgEVU8w4A31AWRFeHfQSjd1LNudzeSBavtLRrb96Gp2uqg
SI2hOw27ajwfTrAwQWTdw4TzBeoww4/g8n41bLjUz+iaty9o2NkFqN8dZ8857JvEHWeEYMbuLfVn
nxAzyvVlx9aJduEuplbtedPEu+hueWs1ad0tzYbh+K6vpiMpEqhcpxXHRtesVwuD4go2BwjJwu4H
5+p4nN/jO/KxH8fOBlazipe+DvCkPG7M4fGDWkJsExV0bmf1E7cnZ0dkGpsYUqcD2gkXle42pGGH
QxpAUIcQQ1qgyWSuymboNwNQelF8pHCTjPk7lW7uUK6REjs6HtXnXXHxmkf+3UJ+NELm9AKY2KLT
1+mRJ+Je5/Y4aJsH+MrWclhfB3Dw8UwKot9jx/o1i+AQwiw6IKFJZsSQ1JbskoxrAd8SOqmq9cN0
3wlyWwFgZekzlx0h9HfPwfBOjz/ihXPPfJ1uNN2HDCPRaP1dbYWXvdxHqtZY+9lEx8jv+SM/Hx4/
97PGLNpBjkm+NiPl5ivvB/C1/kZoTQocf5Sy/F/7gPWH5aBA22/085lePupVoyyPWnQXHX92yDrO
KCeiEBv2GBUV2wJhRCNYT//uU9xUgikaNXmzSO9HK38dTWJ3EP9FLEWEU5MOuUSiBMiJq9KY8m6i
/GJkRzVWgAYeH+oyaoslbWgfs5KFoqs4tkq6t7NnZh5kuiIvGFVH19gfcLqB6aMT+yscjbZKf5ID
bzL5F/Ttje0ClaGA6r6zJu4siUmlk1WFZpcyVRMjLGPKiOsrB7dtWGtXkE2mIRNx8BezvLKA075y
n1LCkP2Ob924DlfCFyuzLDfZv/c4DZcQg0Pj/xrFSA69CRb0UGTRm1yyIAcPauOMgFPzYqZKgS/E
mgQraCFwhw3xgzOHdbaEyPkrEFG3wQIxgOQel/p6t79Rc1AOGmpcjSNC1TOw3nnY3aMaqRkqCwpQ
HpGrGOrVYYQ2xvK5E4fDgWKDcZDKpv+bppfeERtLoT4W6y/mg+ItbrXb9UkejJXiL3L31BQB4Ay8
khTKkiUwODSO0o62wl15sYOgSntPchK7SWMkjAJc44Ytl071twIRnWeI32xxoSkG6t5RqH0FBcbs
i+hIALek42tzXhhwWgZBqGW21DjzH9QO7XdrruAcQ1IBFaoG9vFn4oRmoSCQczZjW2JsdUqlJuoU
rO/dIxaSboiM/NwDULwUrCRyzJCUIhjC1d+4Js78VqBa0hN4WuQjgdA7hQBDwF15W6k9WsjcTM7H
G6dtXvPmKN0dMh5K4PXrl9LPjQYNc4YMW7302gwp1vDjiloAtFE84lvtuqkr9UTzl97V0Q/cc027
coxIPMFxSGzCVQkhaGfpIct+Nn4V7Hb25LB5IvyYfryPEGktf9ic3cCty0PnBnOrQFf4eQ7CUIok
IA+cEhvTrJRKta+0CD7HlKKmKk0xaLS1knmkdZJBWnPc45OVnoyUtIJhownf9ZemZD3UE4k8Zyj2
9DPrK9Qh5xp0Zcl0gCeCHEC66nPiOTQlvLWsoVqHfSgwFdkZmiHtDRfuKZE6XXZKd4LIT4rClPQt
GGVMQndGztbEFNrhUXVM/R/JEy1m7JTwhhE2PBMsIJ+OgqgvbqQ+iEHYcoNQDXgn6aKPMBuj5ytu
Htc/GNhFI3dHCpA8aSXyzAmtE3QfxYK6FeTp/jFS+lS1LMHbA5WxZ1A+I4ZMuRsonyDPO6UgtF8F
ITE+wpK+BAftcOnDx3A0e14rKRTTiWWyo9l1S/1NCftWJjAkt3rg+CBhTQwuHBX3X+3BavPUr9e9
NpIuNah1U0Au9fWEXb+3ZUdOA2RQ7/v1r3sX9XdBNJXJX0KVo9Zb0rey45D4Yx5h/Zqtd2N+yzy2
KvDIkvqkG/r8JXrsfkb8Vx5gQzGcrSps8WprvUgD9MnLvdQj6c+/6xwvg8bHkHJKsatCG4CvGjew
VMz46rO+aAgNPGfQHbGqCsKTqzNG3LvKBEfcYFzG8h5Wgjlepq+rOCIBoPOkt/ZxKrmF+l+wHVpR
KeWI4vGD64tzeVY+fFywTDsXIdQ9j+z1wJgMUqc2JqK+KBpDbxTPdznMmHOdWfkMk2NuwtV2x7zI
wG3h+5sUgEjihex22iAih9qFDcwr0r0vgO/nj1WYUw8cEl7HYejy6z8nZFARlSvp0cZ2nNM7TJzC
N/kgFNQQ6QXKNfzm9MaKqkh31Xv8vaUJC2Dtx+q6k+QdJbv5QFcQkWDFgOvEMBeXb9A2DE32Vade
/A4e35tYQR2xcEiO/XYLV+I48YxlGbpYx+WCF41Xgs4mRRhTRAlRPglADbcu0yIeqd2Df2/myFNC
4ZwjM1w39BeY38taAPK4feMJxtOEmlzjcjeS5x4P11X9akKuO8c8qfBHvdcgy/7XdYW6efcWVgFl
yMQhPWtjJqK7EOX0xKLckE9vQdj7xriFcB1X1JaRRHktYYuOHK+o05R2SYX1n9GBB2ct06l9Bw6X
MxfoKEqFVfY3xWHZrcot+u26Q/YmF/LmSDnelfQgW4Q9UM9CVPtalOT92vd11YLgnjuA2ntz++YM
Tiy0YnDlIOLdxtrfXN9Xv634Hi7UENBtiQctR3hxsDCSFGH7adxvcb2FK3BkKFhTTTRBS6Dwq8lL
9207mIXcjJjE5BaMX/Dcpn1WfAw9jYgAIPy8rzbbjd8QNKarok8PY5pkfIX2fQ4rLVc76hPT1lWq
k4SwbkYrzqROUsmKa2MofVoaWOzpscZZ1iuSF9OEZKRQShBQpiyzf4dTcrnmvwpuOTpgu52ykw3g
IJvJnQl9V9qvS1Wtf05EGtAS0bh/AOYqLR8wRz7xfL3Ak9yUdY5Ctr31T2BYM/9i3AQXc2TyReLv
1WytJDpt4FKAXAGJuUZWyvv7OxGKmR1jyx/PRyjU58tAjBxH/Jx+C1445IKTobzkOFuEx0F3GHUL
cjJWz1/HmyGouWaqBEBmIHF3LzDAKWxoGn8DcrbxjiBXMuzY4bWCyCN5SVdKjgifv0dqhJVzKwYm
WcG1dS2SIj3c6nb+8RfxkaN9w7kypZVE2I0BkTFT39NJjL2e9lpVPb4d0mNNNTdSx2AOU3/PLjwJ
J5ktMp/+a7u4aPI1ZdVzDjmceczBYG6F7x9yGdrGs5uLXjz3m88hojfpNv62Yfjslp2ZcPAo1lys
GtcxnT5sRVHKNs/D5bx4JKfoXvJ7Lh11c0NWYPACpPxxi5RSvtH9JAHj/vYLAZUIVd00KLUbY/tu
k3J79008hr8KHh3UpHJxrfqmKNwBiook+f5/uABTwrv4r6sOSmGSgMNdD6eN2cPHwKGxpbacpXh5
ez1Sj7zEAPs4Z/k69kXBMEkPa3Qxdu2QlPZOMTIF/2Wcqc1uJvgMWRJDtGcs1b8J7PmDLyeD88jf
kIDQRSgy8JDxo5gpsURQoUUQ4SMv0sfcJvOFThPZFKRgb9lP4s4YS7M935YRA4MyRPIuA8ZKuKHV
E5QX1bDxfZH5H3GsWICMTYCgGGeHQAOtA7WRDEByz7vk7H41hSlMmZF4gqXuc/4ZTZ8oBfRlOyJC
CvV3tLtS46/0kqUdBWGkPZ3RrW/mG9vwNW8f6BuoYa3Il92q0NKRnvQP6b5aVFti3DAbB5g9IG1E
63bTHXGQE+4eDENT4i6Dp9saYpODgBnXo5svZvYuQ2TeJ/OvxeKBiXHi2938yN+7vv4Y7/o3Z1zM
F67kNufNqS6n18rLlCAIM0DRscS994Kov8ZlNwN/ZrpHnDzmeXG01Q6V28Mg3elJRlMRn8GOuOA5
DyiUcbh06sLt46E1uzjBsY+uY7FzA59ja1aHoIAir+wl2pnA6StUHbZDhTytQo4uZVKh1tFZ34q9
UaDFezIhw1se1I13oopa7nCoBH659WykOGKJQO1DRomgUnaGGS1HbJlWWnR1GbAMP6lCiSV18/da
fYZ95+QYuNeOJ7z04ioCA+iCBGG23ngJTD6mZJ3s2v6HVbF84UVC1ONMt7xCOSetITqSrz5S6fHh
rELCCFWwlXOjhv13VFVyL+FkVoVoH+lTupQ861zuGHr1se+tZnxCeslRchqdhZWkI09K2Mm/tx03
CoN1ImCWbCJ2ygmykM+fF4WoJqS836wnyb35nL+JB0SbqBa+gmeswOuD7qtyh4QRBOnvXYS1ZWKa
Ak9Hv8qPFdOw+JCfTTFkU5aAhSS1j74XqbykfIrLYtZ7o69z53DbNbqjjqhLFe37cpo/IMcbeXKZ
YhmLOEpkrKcf9eRyfRC6Wm8d82VsX+PwwaG/REolrt7Ao6ff35eLDMI5X4DvegEx5aPX3cj7i2zZ
ERN6bPncZ3F2QL1FnLE0NiBGjn4shBht+tjjQmVf+JRs8u/Zx7yyb1cTcJUBJYy812F3yz2TK5a1
U3F1DOK7K+xyp5ap27WejRkcorsb0vADmQ/pnYENw231BROD3CLlT2/j7d8HP2uXz/LUNBwSQA82
yapC/0LFdnTbv7sKB1OQb7I8kT9mfyqYijn9u+L2MoTGsIzrlkbPNZPuHUIW/Jh2WlieyZJsDGDq
csE2ciw4AKctRgEDctPMF28IgswRF9J5t+IkvJWUkZTF/+tFUF6bRtHGCjqP2MLsKiVWcKsKsawN
jou2fsueowzufnTR3S5EuKLBoKtORMNvHUhGdvdtXB+RULYn9U4+czwdoza24TRSnB/XbypSJTY4
oPyNxbfVjYMk1aIe96Iv7yCCH0YGU4NEiB315p/owFSM1ml2TTc3cOaEv6y3rylr8KabhH1+DsTq
IU2AzofN9DhlhbMn0qsQhXlgPz1i03DSE7dwEXmxchXbzytN3dZscHnU3Eu6+1K1UwKI+W2StHyS
NFJs+D4IAkaiPAtJmhuW/mKiCMh4PxQzQwoXuKsSpSokuwEy2ayHrWAoEsvJ6/na2kDSIwqiqxqI
FZ6mzy0BxdHPdv7f5KD7T5WULsIdaLO6Lsvxfb+V0ioo50qVyy300z+6SxNpQINhNzU3u47gZOci
ET63q2nxFALwur66KYEGmq1Zl6z+tPZ4cXR9xEnM08faF+Lsjy4L959kldEVj3z9AwayqmAsbTbA
U0BFma9V2KVcfHWrTyiDebMq3ED2fcbvBi82Xbr9G9Jmf8PEQbuT94buKlVD4qIlbfcNn3Mnkf0n
X5ZcQEYmX6qhTDc0CBFx+brFokwKHmjz7FF+XGJeUWjlk8bEYlaL0F4zRub/+FTvyHCJb/Nbf5UT
uXcFWauCdeGHxpKJemHhJc4HwutqQAF8AX2GzMydoapV4+5Rg3okQ/gNzEpQPDzZ/bMJISfEMr9g
REjxJJTsnGcNUrN7yW2cHAfec5h16S0qpW7jzJfppQIaaG4QsIInOPth2I3AwFrUdjSEH2mrQ+X7
z7L4jCslhcYFbX9lGJLC0DzuNyKtxyuXJElSTzUcIz3uYDTwIbT1B3ebK8vWPK91T/+aR0am2WDw
yEmPS5/EPXeNseYlcG6bVaHeZtlsjttv7DCik0tNSzrFat404G7uVLgEKrubTBxgdzqa2QFN9Ezu
9GDWG9VAKxAamCYZ/M8pCsh5rLItsYNQA7LOjeoaeGmIilFO8yRYH7Lauum3BWuypDnU5ALjYggU
F67I4rVBfo3L9Kvry1BruTJFCoG2Iwn4FgmzuOZFUv+/4yyCM+/0yG9u9wiWN7fpBKKEvsiKIO15
VEKPvZxlL0EWzum25yg5sgGXwQwTDNRHAvKIVpyoufT0K5fNgO9s3U3jahO2PkgDbuPQcxoyE2uE
KyV5tOb9hvD1R1YJ17trV2sQ+hCFHKTSXf8RHcduoxeySwurM56Upfpq56vio1EcnzYL7ftlzC2h
F1d26L04Yuvy9RXhGwiIudpuWWBRzvMTmB5wsstI9Zzt49W/hoU3rI3EqQBZRuXJbYHyqMp0ilyx
0heDIElkyPtbzYQV8AVWbstoYj/z+8AtchTK7Ox39JT4amWBtB5txf2Wj3AQrQjgT2D7O3DhHEB2
QwzKxcMaAIBxD2L0k4m4Qj1SeEAbfoh0rLDRCERGmtMnXiqN7tS4GWDoNqgLk19ePsJDGfevkoDy
+ZI3vUyifnZv9xeI4CR+MnIJKHc7mzAbPPrHXxTEImzCNKyQ7JC2/9VLknw3zJacPFIzWBjghaWu
Q6rtAMiqFUJUiVplgLbPC1nHbSjBd3MJChdHhHRy21qJ04vThv7BQGy63aT1GZVI7/UEmO6UFX48
9NqU7rwE5QEIabCYUo2Q/bShdQR2m6VQCAmcz+EpJig5svFwCEbEXW9QponYdangjsXD4axOryRB
EtXfPe1xtX5Gfj5KgOUAT2At8cR5HxBC8LAEmibvdfJka9O9cGe2kZvrJVxecKder/OhXzJULEI2
DxcSXFs+Zdi70Rjd6VpzDhBLe9BssaWXZ6uiZ7l5RtwtYkf+eQI6LkJVqz+LyWCH+T6r7Cr3Wzxl
1ecBVDnOrjE8yekr0m7glPuca41aCJ28j34jk8YQlJ93nQHQufJ1QSlZWWUvA9q4Oy7wcQk3ZEh5
HY7dM6Mc0Jjso4SZwBAI9slIsjzwPvjc9TJbE9NS2ko3jGb14mv9XP8OAHKEW+WcsNGLsz/qBTv0
yE2LPs9mHYGJOEtt5Piy0jvyQJnqUzWDpDlisPG08+1w4Xf3UPJlyPR9reodggw8MCyI+eG67VIj
HFBjwfmKlc2YnEe4ThCTcE6rAgQOZv7Ss6RbFTL5/rrNWBX7y4cwJ4DfoqFtWAHUaanU0IZKrCFu
a/Bd/tUcRtuNPAnjrQwcMgQ6C5h5tG9ks9tQHSrdo5qx2OumbJMewPcwjWEiD5itRW0iD1oObbpc
XIAK4/2IgQDHiScss6sxrLua3V/DcZMPfw37kX3oQFfSIg3xW7g/QBxASi2WDkwvDiGXAQGDCDnw
OlABYfZjZrOXsFugSC5x4fia61/Bws/h9kaCdutrzPmI0Cwx4T306xg8LOZ9YgXYNfk4qsGwoysI
BQ0oMb/xsoWS2Cfu3L/lzYdUTDgg7nIGiEi9L8CQHU/4wiz/Wlk2Os7Q83F2B77L0yVfx64Q0rfl
xmCD5v6KcbwNNoNKtVT9RRWb27ayrxOZ5wet5kCeYYjI2mVNrpkKgLMVPR3yUhIdLGxr5fM37er+
x9DBLs70kncmD0juqMsE6IKbxLGSdWt9li55MjQVqbgD73BUTccxy4aBwq7rIGNrC35RFt3Q5h9+
EsmG8C95iezYdwBeZyUEmKN7pV12SJdc1Lq/JvCv8RMJLUaXMsgIaGYMNHHHDz9bM2COejf5V2Iq
xWRfXKMyiERAy61U9OxGCOQ9yCBzskkexY3qCVhqmwer546wUkLdB1Jv3vb5UR4K27hkPu7fNEiN
bxit2W03/ClTKZ5pYQx2fSG2+AxtSYgk8kqIqRFyolhoyb7jJebgn2Be7z4TxYD/EC22x9qHMtZe
X69UJV94giX+Oq6XuUMvawteOfVF00K0aFkv1o27YZCSe/veGEtP0qhVDK9d2CZYzxK4PWt0EnG7
8zXCg3AdW4v1J4zzMMUlKkbTqrN/0qNn4nKTznWQt6+V0XNgnT1Ab1nAWluXQpDG5jeJtR9UjKPc
hwr3XQ57hZGTGIRLUKSAUoSBuq1XUCRb1rmk4ccpDa4U0WOB9S48Dv3Is3NHT+GaQpLCA2Wr5wZ3
kawz8E+4IUqS8uxIVnfYK49t8IlEZVboZ6ijfM4ZfrsDMuzLCwtacNqnvxq2kokfgKWtl0gadhwR
ts1NsTS3YtufvqfdcoYniZuyQYG4E8OVbqmd84vb+IWsGRcffv0PapbuSPIVhsYOfdhVB/c3rAtA
+7EXffbpkvjEpkTCGeJGtK5PdTqKXeGHjXlSws8tWQneZHD3DMMIuRk0e8Rz2qVxFkjYODDHJDCa
hZCgogIn+GL1UVahhdudjzMyoOPFXc3EFaQZsRXvXI1yg4UGYuPPN7I4GbB7tSQJ8wkd8meT7UDN
hR3gTdxOpT8rOzv38f/dfrFGUH0MjrBTYp7Ie10e2+yS5Ixt3qevGNvFiG8BP4cjlknxG4chIgBQ
ZI8lbTjzonFsNy/cJpaDTP4B2ul21jI0Bzle7THCvyvTql1lw2Hm+4EZeTSIcyk56RRNh3NICAG+
sG/kmlJWkDme10d+E8HnYRW4KnTdgb8hZYclOYJuEMZrW/eMVvIxVwp7efncn4xqWRi0a90LdP5Q
rxxDBuDeSN8C5UPTdDQIWiP151UQYe2GsDMwJjwm2MsrL6DpTjA2nqUl8v/zJ5EbsbdLgmdgA7Bz
lnJ4nHt/gQwdh5ILTVOrBYLW0fP5QA1RvfBib6HIRJSnRJJMUkMcwV0sw8HpaE3ZRjFq6wFUtcuD
iZgK+5oFosuDMBnoA+zLJiRQGAZwNmyQaweyKDMREMix1NTPQoOZ3fijlfYHzrZw7VpG4am3xxNT
YiblVRis1DmXTmmhefQpUeJ/InUVcpOOzcovakJ9dakd93jZfiRRPKirZa7sZBXiO/q4e8ispzyX
SAKq/aTh76OBxl+y+jA9EC5mL3dJaPfcZOwGpXUZya175FzyGDfx43XylNdevGuDAPaRWdLWrHjL
vWdpjJ1uuCTSYHsLFw+to9/ZIliVr/tYeKW+LmR6OxMM3VvkLaZ574i+zSjKgisfJmp9qlWYq6r+
ApzRDFDV6bj2nq8iVRwvWbxIMSXGQ5zP7brl0F1TFbeokbWjVW44AjE1Evr9C3/l5BZJ17/gPSkC
Bb2FbNwZvrj9uMnrlnRtdvUPk3HiFdCPSjPNu9X8J9Jwr8eMRTxuWtwebav4AAfEtmK9vkOJAYIQ
P5H/l7/QSI5FS9vcfBksd2/ZtQC/+nDYlrIC2um2ZPMyvzOnjlTU5wrXXrwdJ/DU8WXgAhmNbUof
FZJVNuZeIYJ1xkBV6bHD6xXVoXf1sfQy+BRYu2pMxju7eRtdB+LhYhof0cbkHp1dyF7YkZTYkwFe
fao60+1+Q4+YRnn6A5RfbYMJO7hwr1BPtqCsquV98dhkJUR1gH/ZG20Pg41MnSbqNytiHII/mKI6
GTMTxtFuDGjlzTFHtQ9HGnI0VYKyL8Lpcb/Bui4ifQBaoR+07+643TWUl8/fs3BO0JNyCm0Syv5v
0LIjrkRWU85iec1xvOvk3RDnk0aF6fdOKx/V9oerM4/2h2pPT2/lcpdSAPqxPVIcdXTxFKKIIVCv
jWTRJziEPPJ0pxjg64Sjo3wOcX/S3E2t0q9Iz6b+CkN0KOTf9j+fqCbHu11CP0CWSGNlw+Viv7K3
rxx1X72PkE5ybfz/bJCd0/RlRjogYDaCxCXia3WhTR+hbw2FcokmTly5Wt80QbRiZkSnslf1dTAW
BsvUPqSmPljx4pd7d+GmkdrYZLUMNX0q2COaQE82goHtr6YW070dSM4/XFmgO3mPtcN06dz9IhdJ
HojT6HjGAclyDPTCvQkBUhhhKqo1I+G9f7bcqFre2CAB2TypC/swCWWNJP69CPdda8JuXx2PQBkz
9La4f0ENpo1u7hbf3p7Vq/bFXJ/mHMvLK+yheJBLvfDRF5Uxarka+MUS4I3QVucOCQd6M3TxDbL0
nm3slVtfg0IT077iY1R4Q8U44+F+8wdfgmqvp0K50nxZJkEn4hKR4PrtBKLHnIhyq2+cMKhYx/WD
Ct0BNrIGP9W5D9My6vlepiZkupFHOLT0QowV4DxrbujKImuHpFwi+eL+wPtZPeky5oFZ8NPWE9VL
5UdtQ2PJk4Wy+biw9H9OZZ/+THyBxyRXBKmVwu/imtjS/0Th3ME9f/RsR6LSHXWsoMpq1tlHOBgY
rFuZHEI2ckPDu8PPmAGJNEilyo6d+2firnVAueXMxyz8OyY8XLfDdisgvPlRYdS8SvIOGP7l5RMv
lZutn0s+vhmrY9qBI3HiI631ghKh46PmA0sr2WfTaRfaCSjyBcJzqurBMcjtSopJJhXXf08uV4F2
p78omY6O7ExfMIwmjlXk5nZ8tIpIy1soY8zeE0lTc8QDsVsDSn8FWqlfl7X3BzNZGNMKMj5sj3b8
TZe6FcFVgLmMxjXhJXt2TZVRG/iT8J8W86Kvg8XQJQCahHbRaKpfDlGZdfazI8x5x7HpvEYRHLT6
pQHnb2HTlUBgsMV+OPz42s1WG4kt5CzE5ChK0l+Miz+9LTzw/pvGPhxp1lmb3o2sb58bYbKWGiHz
nsnEoIOtZ8+nexl70Oq15/Ak7nV6GeMsm029kJPstJlNpN2f5BvzHrP+5rNs+e54xIRTLpyxpvmy
1hkFX+uw9Wtqo3RK4TpfX60gls55U/t5d0DAN15t2mHUSa3dz1gAJIioj8IrcfBqo5DOXpuQK0sU
/t7+qPqCH1AgQoTG31S9bIVQVPFIDCrdnzYZh1bm1Owrk3ckYHgsA9i/aSn5x0Ik1fZqylJQUztJ
t2f3YBdRwf1ZJP3IUdVnOoiIy2JFUWwdCzq9jSbCsD0QLqWcMCA0buvIA6/aB/omFKjMk1a5UjEu
kFz2QJzvFEnfyMQ02RlkDAV4S58ttm3ygtU3qGRoJNFpDVS59xyjSsHPimyDHLmWkINwa4i1hDsE
gGFXupKonGg9iKAxttdegC9Vxo5YH7ox8ePITzs8EwCjaBAinMVHZi0WOLua0x7273mCB2OBG2yo
6hS/mBylWyjO8frPyM92Fl5Qq1olWqNJX+oRF/LvOuWN3U8koUvKN15s9d+Wlo43WDYPpdkKA3CB
C2VNRvbe1zheWPAIoSS+y073AZj6H92k+3bEHEl9Wd7/VI5cHVWf8EuBiwc4FsJuR2uvFKN8mOSg
bFWRKhHhvDYshJJKReVR2e8yZ07imZxfbLWIgB/ZlJ2bU7Z+24p2QarjQfYFOU+K4xe/WK9DShXX
115Mzfwof9j0v780WPI1FIS5x7uQsWZX9Nm9rVY+Gmts2mIQne4GG4JgVl2I9KEsCXRuTJ09FmEw
ifD0sbkmCLMiWOPFz3GaxeiWkRQ9vcC02j5BT0Moi1DQkK90r1hKXvHnCmGO8jxkqyeo5d/Fe0iP
ohR8DNT2HXT2muYcAgkwIMTWaY01zsjtmQDLcsteWkKN5/PCX1RNSOlhkCaMN02azwDIznVMTcU7
8CCKuUXZxKPTqICMFqAEZ14Xwbs1Pwgljqzi7fAmZ1E4sBHMOX7e6PLIMw8IlByKJ8acKzB+V25B
BTS3ccSPYymvCuTrvGWlz6KFdP0z02w77x1WPFJnA4tUrW4UNZIJlCIbvcMqr2uYc2V57tNDkx59
A2NCg+kGZ7BC0CuMOukDcbMWmu5lEz5qTBe51q6QL5wOcGVMp5g+VdTV308KkLvNiVlF6tVqlsrZ
B+YynUD8s8RcDab1PoGxQv9/uO2uTwWZDj+8+6e5zPgNWLxMrHB0Sc08/hdnyyXaZ08gtJ+Q1P4F
bf/QYWdIMO/nAzXbh1y073VQw5lQ08Lk2nDun8YemibFldWxEavngBP1+NaORiIoBate8nO7yzfZ
R+OyQniL5VJp1tzZlLt/JO1NMHEuS3fQi7o+/x22qjPyrS4X58n6qF+wHDbxfq+SpAhuafKJFtjL
wM2+3zylwnAE00zWMqE0ZLMelYpm0VhWFR2tae/c+rn3nZOFaGUD8r42HkQ9HOPvmDvPNL+3cS1u
ppMEnjfuYQ1cs6/j3JyvYB2mbqc1LtX2dRMki3xAvuGu/vmtPa8cMV2ivDNHrDTMWXXl8QMsleoQ
2U/2jSP3BMXuQC4eDyTPwCWlaEKDG98/ZlV3s32LU1EfuRh00AMNtKGhhlvamM1yYVyjoKeDJCUG
/QxXMZSDk0aj8nBAq8cXkl/DE0EmuRS657MDXRFnwmPqZJXywJTiBDB0BASJV80RhYHunROd9Nty
HmAfpV1iHtqNhn+MQU1xYB47alTo/Wb1036RZL2AzNiWc09lR3gkVXtCLfQb3ZWWLGIZlKl7jz3i
dotQW16viK/UiKHG3bko9eR3Rm2Thi/3nGfhuwNzUjJWpE7pj8+zqjHcJ6TrYoWXHMlDhUTWx7Hb
wBcIw8rR+4aTZd7LpHOyfz4gcIPewB/YfQ7xFSM8Jq9L0KtKeaFQ6wtjKJ4Oq97WbogDCGl1lG5C
ammAmCwae2a8TKtn1WKxA08eel6C1fV2VMcyGyuvIVZJucJ0N9SLMluYKW6J0MOF9/qtY7eryMLa
7HMgyo9FqD8NfaFi57sD7CZR0JgZXOe1BSn6GUGB84ydeSjKMjp9NPDRFavP3JF/ouaxNPnDZknH
CD1OM7/KTZd9QC7VZRH/44f33/NxfMons7Z9Xgf+99mq33idjDvYWiUlkz+C5Tfv40hnjRnqw2Jo
NGVq5FGcCy/94h/cMFVnMoUJ9Fq1kAqwlbnBBlZ2Axz+c9VpyMpLi+Ekokq3crcUSS75dnQzNCBI
YAiqZZOG4nyMO+ijJcG68saPn96p3jN0SD0JV2OFXkVa+koB/xz63EVv4J0eBg4Jn/G0a3d4wtz7
Pmy8Lb1n+F4IcjI4tFjeHlsjTqtiAYGEnnOVCYtaYSjbUm/KP2T+gbbxahUeap1INs1LdrkAEPIM
XO5iVq+FbYIzZcXd98Uzwqyeti3RJz6vvQoE5/l9zNrkSx+COqJK0dZxFa0xExII0AvfoerhE5on
L7IrnfKjO1grLpGdTyyGK6usdGtxc0kK1LOSlpjTH3WKfA09MRXFw2eFDUx/2YeIupEj5skGc6t/
Pg0FMvEp3EG0r9lq93cWBwcLHmEES194YQvpaF8yTahTTtW32lno2QD4CvGZK/djXV5Ajg5NtRxq
eNmjY/OceBiUALZbdJeOC3gE7h2syN6cM+Voif7EQM5N5D3hgxVhxi5GHa8zutlDkKZStBlDBY8X
uRiZfrojZe3rDhpAc7wm0YHZGgfIjHN+GEvEmR6SlxHjXD1fJE9LDhOracMUaRvdRfP3xh11LXMJ
gP5hSyNq+yLQBMFjjqmqDCRsTA83CQxFjXr1GMGxjtqjRZ0lJsoJZWDnXx6Musp6r4/zpVFogcfx
N0JJ9sfwj8ivn6IA+WOAV8A8d/nj+a63z5a2vfK+2KJA12d+AXuKsgyWumOqxyWGQJFvsfmd++fo
TT4kUVCdCDxqLoW8gRN3+vPKNh6cnB6qBt65iISItk5CkTVMjs70iZZcFu7D5aGN1yM9TnqJpStE
wEHh2QueD8Ss6c8ZnOE2+ha6vG6gffU0xyu6vhxkNU7gidlCpD87OdWhoj4i3OENlWZ5Ucg1b6WW
gaXum0iwYHZSER22yC5/Pm3VZRB0dTu+AxDW6w3hGHM//NgEgLuFmRrbsSdt31m+PzKKYYBX8Qha
MGSJmOo5X61l8baj7oJk+nofbcRI7NMv1D6swLBM6sTb6Tx5BDXciAL833zdAF7P5lUP2sxYgcCl
jSp8WQhfI7QwiWFh0C7HN2EokgcDBpiT7Muxrh4KVbJZnm84IMOv7au9HXeyEaA88fMO9pzua1sw
On37k7A2IBDnuIWMFmLfBah6hGp7P4Jxol81SQR4T6GCIWq8mVc52gHdG0WExTLq3KDXDnwakKuA
4yiUait85e10fhvnv5J9e/OZ3EAm4SjkQX8Md9KjzFyWVRyZZMcPlHLJ6E7pXBiJVXqF497YbgLO
EyEItu0sfeAa05DJc9EBlZT9F6+RpRxAN3MbZaO3g+rhNFIaf/ro7cNFrrtdd89JlcxmpmE8KSJe
nv/PcOziixS2/fjsj+H8RRwLrAzPpCLiCSvxYnkXbHM7Y6qnkzoL3G8mTCGBHpbzVYYlILYOB2dB
KKdIuqj71vKjSQ/Zcpav9wUIyulYJKSKDTfwzn72qtO4EF9KuzEejB+LuvUs9wiji8GJP7z9fBrp
kE/ghhP7r5kp3vczDnjzhsyJ4ZifzCPGjWGFZphQHrv0ndaqIAjaPkAf2AtlPSIxZX+fOi+5nEeF
BUGASHXktiE1Jz1kA6pd9xth9LsTZGOumbHoqZh3xD3/4Fdx/hzma+jvnowHGCjcL8jYUW5XChay
IHAugfOAL7qs5e36XljSAn8bYGfH2WvL2U020gclZIRRtyqQeev/VhosYmyVG03YwZ/l2XUJKq8e
EN1VBXwna5rhi6NTSX5++pzxLtCWJgS4tu0AHxacIbA1PS0q9hS09yNYUG2IdKnLMxWmVpAZ9RIm
xuODkJMCrUqYbt1Fn8BoAeGEOPBJfvwuyHSi8Oo5n37rSv/vD50mHfpTsOuFz0T2Lu+d5YQLc5GA
T9sK3HkQcovkKRbROr8mKhyUqf1QMdSz3ZXPMKUvvGG8Fsb+mGeKzzBTPKILH7PDgLdGGKlNzVHO
s3Roh6RznD1dl+ZBQQV2GHCxVEByFwR1TfJ0SKM2rnNcg1Gi28KthFOoB4EPSuzvbYn9B5k7s2RU
1yf/JYLVhehEIIQ5ZROip3yVi0efBSZ9naq1fLj1HgbKa9sbtbVBBOJiahA9QCtd+Yc/9KdUt4E9
IjtsVuyDdjy94lrNe1m6Xf0rQfhuRMJ4nKEtuWRIXu6NZcRLuoekQtUEc9ekQZeTmjGuK2alPsQ/
VJohEkfo3Z6lVNKxkIyswTdUcHx1tNOOd2Qkt2SPlrzlXJw98ss4EmZUoxbkOT7KpfLqVsB/3E/R
nVoDZFvDsRiLPXFog1zhal5ze7E/ljh7SwWcp5Ur0cdqRa+ZbKboTeh5vmTT5ffSa5A/fEfuSizu
JcuSK5lBAvv4ZItPn3nN+0XZnQsDeiHO5Mv50EoXnZAGVSCUkCczY3OHXPPyD3F4XxfGgwCiIjcC
Ktcx694Fm9mx9rMXxw0+NVrJ7Pm3qVbN71/V4OjuJKTFhLB2rTzYzItESRmAaO/Cs6P4XNx7QiS9
CzKfajr20Hf/fkb4xcFThtz6+b9wgN26AV01VYqm7iWDJkjvMZDgcnSZqh92IC1M70161NRk83xm
BczUVgciM//efoUeJHU4X+IlVr3C0IfojXFQl32pkT8/39q20F1hkfGZmaBChcLiCxmm2fwmB/NF
SVd7hTriN+0IhfHMqrEGJafUPG9OeLtkI0sHgFNAaEV/C8fWmaP9f9KvXLzbYzBgp7RPgbBXYLwe
WoQmVtIfeOBmek3CEMyV9/MRZXOazR6DuMkhVk1iAORKW5YvVYrcZ2puzmbiyBftSvjOhr+zCy1I
IhtQ0QobkW5VOz912xPt4iILw/SP3xo/vVyGf6TwpPV0rVPlEu/pQ/1eAYI3POqTiuLckRcCG1F+
32BFyMzBuOZopnCLPe9uxwXTl3RmYTecR34gvvt//IeYT1L6/sKpu7/ALnTbCZoHGNmu1eljHnQz
F7CkYr1KADWkZFMYc0lauScdifRJBesRfoXanCPN3zlRCrw8g5FjGLtPxbUx8CFgYBhkQ6jLbzxi
5YbYBqKlumHZTMx2ouVEEnDx2jablZjCLiR644vE7FSbhhEeeOgydZPwtVOZ72a6IcDR95IidjF/
1He+9LzsGcvMcw7VBLRB5jMQwFt/MvJsFGStg6uOkRYiPC/pHge0RfplabNiVD7j+8VogZwcAZvn
Z9ZTqw4vc5UdEjuZynMPkc1qcGdBwxbXWdCucI6L+osdH7rhtH2ixHDgel2RI9F6j683IkqIPol/
ztn6FCh3aWhrB2F4zM/gR7RuvyfuOd2+FxB0H3BE9y52xKzQ3uYFTOM5OSGH5afffsW6h2WiTNl+
WMvpUhgUmWr9nv6DXIPeQyqJGSGgG1FURBA7VRm+ftI7u0AQMu6tSqERMRbU2U7+2erkP5SVsMi6
M5obZB3xuFB3Zpr9+WJ3ZJp+3AXjpSb2kr+SihmF6xdsFA+LK4o6smggDzurh4trqjVuRgVG89Br
GOvPaUlDCgyC2XvYDm89EGIVqLMdnhErwLlrr63XExGBTD1ah8usnSp5nrSM3In0xKF+0zek+4rF
VN1jNwxhwz7hmlJw4q1mlv8k8NzxhvmprUAr8NXOAAfp4wPMcMJTyEYWiOtG+D00bGbNjIFvCTbb
IxDAx3Vo7PxPMB8XL+aBDYb7WxWxTNsCYT4EAVmRGgNUk/Rh0Jsvg21inZGkBGazk5jNWUfos7r8
GtAvXsT6rcsHq2KMEBm2SZpWL+4MGe/F2nQrBguGXVhqbICEJoQ/MAQXGsKf8UVY9X/IvnYX81nF
BiWiOR1kiVO78cQR8bz1053O+Cak5EROQj7Z1g0CIVdmCBovz+ku1xKFMrm3XetbxgkFsTDwatHa
BJXPy1mgsEe6ry0b2S5cD/viHx8+8NvYhnCeIb8zaLbsb/n3Wi/+Pg29KXfwUXCkw31QPZShATgB
U7j+Xs9GOe6zF1H6vOJA93c0vm54VH+NDxeWCxsPnTqJNOdkhAa8DFXeuN0+bQj2q89p696MHzdX
edQUrUJTDrj6/32HvCHp883fo8v/W57WXLprl7FXcYou8dwuNI2BanvcgwnkodAkcUgDYReZB9AY
dvwmn16lsPoGfJkR64q8Dt49qQvSluW12HFHBt+XB/chs8Fyzptnxr+iv0CEkEZvPdZZ7z4QzO6/
HsJQlHlcSR5Ftz5mGRZ5raMdMHlFTuxgTN0Xi/vk9t64t3ZkcYsFq2SNCXdTWRBEh+2XAK7BzIe9
wShwtC88K4YPonLr5Wtmp+nXfLzqsQSlhPcuraeoxyO6SC2vGafImqkli5o7veOavkF0tF7Zrnwu
VpQrKFlXEEmhsL+qkrbqwZPKLVxu9/IV610FVFOmR5WXeOGw1gfwzLArjHl3rW+tOu9SKy0MkS+9
BYauGaV7ldgzVuQoo6nCZeFIWlvBi3I2qy2eySfvH4fZvl9xadJhx9vbX8P+7UUep5Xv9EQrItgN
KVUPLPexrMZpc3VBq8Qfb7xVTo+0/HhbWtwZXZ86qSTP0KM+QfTSQHHx1g5yYt1YgFqJc4/9grWO
U4auwrBeJyHU2b+ulMyotc+sdzhRbixTuGQOA/zvE6IP/lZ+0epgr0MADBCP1xJ3PCck4Q/2LR+/
ASibH+iZ4zDJsSSqeHOfXDfpeyL3XDizhqcbkgx3I9GLBPDTgd8dTYOZSU4bRyxY/ET8In1wl01M
HvsfkTZYb79e7kpXiI5N8r97nKB7yUFjryxIOcfmZS+Tw+m37pOiqIDpD1KFVN7QlT2d6BOE1J+D
MWLbNQjEU3kPZYD2lWZWp+T+pLD9KXuwFXmXsTVUkvSDLvur74PatDtfk7lUUxi7sh3oUriQzkrt
nRyj6ccVl2Tw3w3zDLiewvYvnVzT6Ua4zFVblSz3jmapN8G0Hb9mqToaZ4Pvttby1gL/NpUTCmvO
wimI5UiLqEQg+txzEFjHW2LwS3F+Nqvr7aBn5tuUuTE7HBAZjVT9stlTGR2+YzWvjeJgPwOTDHkb
OPQGmBA6riQc20lgMl2E9v2TEyRimgaMjdHHya4z8W+zfAmN2WLeA11pCyTbUvOlcaBEwyyC9/z7
OAvkovMSaQrHejUGovaQus/UmWLRucZ+OG9+Rf0XDfmQ/X5wf9fj0Vw9ADvhcg8XkPMDpYCNJ5cd
qsXbvk/snjCBh073bXN4uGW6V8LnUFdKEguPCRQVytSiBU4TbirmOl98dbjGXxwhw9pW1dt5I+zA
zKNY++hfonOZaZNX8Ra9xzs4VgcIfoq14EAnqsdtRPKiULR4Bn1KR620TaAQphgK9rYaIP4AEm++
A4lduCpN5L+VdV0PlSn3v1iE5HA3lqXoFFHWvaZd529swjHxcL3k1efebHtyyu4R35MkK2jz2ED/
qTwC0yRdqwD7w9OHbX5XIlp6odgx6snp7wYK5i+rhg2sOdY9kzksUuOUU+i3E1Cfo1q4ccPpkz4y
QfEdjv6Z/oIwSagcK5NLK1BAZVqbDEYPJ2lScUetaFaC5nOHG6csQKMxmgH0EApVYnlcwD3QiEtl
SCGkCTHy3ofbPFgN2WjgNnA/c8WS/+RqT+RdYHU2uZXAmRYM2nuJIq3WC8Zd8+/kXMjz52i86WvN
hdLlfLo4zkWhF1+Px9WQtgSkCoQsiPRTvWQ/zGoF1F5VXYbajhLS6iW/yaqhudeZknq226z1lS7t
6p8Tp6omi5Ho5WW6PVVKFhAC1f2XX9ch0nkQbqlMa8KV0MCQfw+aNkokQX7majQLWXH6qsyTNJHH
SyljnpevRh6ynHneOlnqE2PkBMPwEcfvzaCSoivBuKFdCqjmoMWhPsAYnVV9xAudDwse8D7TjRkW
eFEx/hOdkh0N2E0BKno8va3UY/3/gSrYlELpx+/YzO3kfLD3MnqMp/YWENMqc/+1YRtcPKgNhFUI
LodzEI9S/8MxqstlsjqBvfKGI0py4L4RtACGRxTHZWTJc5LlLKurrJ6U7pmjmrXBmBENHcw5uS30
/6aXA4/OK7nM/NAD9E3JNF+R6i92SYSBSIVNAg5c1HiqwYM220AG7or4mYI638KNmPLg3LfjWVP2
NZ9CWVsL6djcuUFl7jR2dsOezEWjIXgOSDel8Sb9rKMJBM8V9nG5HfsU4YfkQecSFkR8POk9SHDq
7EAM6xGr/G+EXi7/eWrsXjeUsnS9imK7c4ew5DdmZ9rHPmBGZhj8N3hikiNh92FSr5nSM4ornojQ
r3U37M5MMeulHjAPHx2ybL1BFawGvc7RYOh6k3z4JaokiI9YEaC9hyEWTdTzXGZc2DJzJXH9iKoD
EvKs40T3OE7OuVJDJ67lk04bbY2Umn30s41nb0yFIanTeFgIOnyarpcelxOPvrqy7RMqjXZsHOpf
5YuyMrO8FZhPJPMmgZG+Ii/GXul61bc43kkK9RplP9iIbZ0hmyPCFwli8iPUQ79+6lF+td+TNvIs
ldSY62LMUXymDQkGFEJRdiuIqyuu/Uqb77Zm5CvY2/aC5E9OvAedt5tGa0b07PlT87jpkPBfCdQH
3Rpn69y1aXRjhQNn/JRzyjoPHXnAKtVE0HLoPHFp/f8pTPUatjIPENoxzoYtaGvWzueoF3wNU/9H
dlFzPBiufChh29+/p4iIgxbwLMLTL9yech0rsFzu9+T6eeChK89LUoY/3nQeYx8zEEfNKne3K1NJ
5r+TZicckgnz/HJ0Re7k4pL8u/f7DIE3RLZo0StxxNu4yZmokvU1XM59kRxP0nyQPf7/TEHwENna
7VC4v/rDXPHSeogeh/WYmrryQVe7tARdLBOugtSqQIOcmPY3qxVinZB5c0iWQ8yV/V0/4dPbyYrm
+dfWkIjHG7WjxGSU12mRbq2Wmf+BevYqUlvbUFWjNMoMjVleWoOz7KFV20NDA46esgnwN2GMArpN
3w437Gv+JPxig5PhvYSCjnB4NGoP1PeFg/K0jJ/4oPX0gwT8GrFQGtXBFPLWL770Xx+YyZNDbRaH
+0WsGJFcLRPugoHYWYOnIkyjwmHdnQdBEhPT0dFoiQztIMQhFkOZipqaZmbEi00PQtv0wDYOr+8s
iWrtPhA/l3gEjZuQ61Qz6+dh9p8asHfSvsDaHnU1+1JyGN3khkGpChZzIq47NTgtc41c4DAgioL8
YjeVqyLX4PQjW1sZn16MtAcghr9cq3O4CZA9Xv1L2QDBMavD2rgNwRQA7XO4yzM9prX8Yrj13Rhm
nqTmqROQYU1h8uYUgFP8tJ7duuY5m5o/qbi0nwctZwKV3ApFEncuNat+JiswpNCrAQCCRERDqwUj
y9SYRHzwJRaW4F84EsA1QLdaEcOAsHfZV0JaKTtAHYz2kGjVhamVciBYLe2gkwIael9+qxml9vGF
N1bAa90/6zzDIqVnuu7FVYdkSXk22ntPzT6/7UE5ghj9se5/6+P6p06sYHXALfKp9iBANG2058ZA
ZRMxEyKsOzpmfBcB0J/RiKa62aORo3QsBtdz9Cx2vqsav71NXslg6+RKBSECTdcJJEdLxqDD+/1c
d2sDLrX5u7HiHZun+hFz+QNPKohQH3dUWrXAYWmQ+JppgZbTgoQkykg06d1t+Sv9LftPfONncY37
vkOEUNbYmE2tF0OIGFqdL34U+Vec+puA554InkOnwQsqVzvaRxgeDT1y7SWSW/dl16p8n+KGJn7F
GhOV8XqByi1NvZ+hQE8XYQPYAWzmb8pOo/fJhTyXr3CmHzulbbUkCcazQtL/1/WdQkEv8zrmnpLo
4vXAs3yQZ0XNKXB+VWQnZ3VRhEuKdpmBKPCI2Sus4muzTmt3QwC9lyV+lcHAdBGfRwCtimPf0fjf
PjJzuOcTWNVErjGkY46SMj2Br3cBp143FDecLLbHvnau1WtOUxJr15HDBA+Vz3YkKRqgX3VzXIpk
nR/1wH+qyZieEl57GpupddGmSugdVoywSxMixW5mrJBR0k/JeoNzkePrXDu0BNjvgCG8Ps3/tTGq
OG2mqgfOEchoB2jK+6hNaXU3JNSNqPyFIs3ENW0zsgafcUpH2N4uOnYlfGSylEZ0fnJmSSVm4Bpo
VgcEVefQR+dzwfHF+PPvn7UdSTlJB3SJDNZHBL9JP9CQp0W+0Ga1QnFG7kb5Pc4qsfxHdU0I0e76
vrFmLYB2B6qHFk5kauV9p0hyjPdgkYGchmEICKw5QmeB4YiPt71hNRjoU4hSuA+wcEV0pdpEpM71
vbW+xVJQrGbATt5Y8i52FrQVDcqfQp+Yii+Ob5VzcSYZ5qT8BASjouh0/D+NfmhR6udJ+FXeEtO+
RM+szKEam817I0cTFPqYwjuIfRrSpDHs+SJ+VUyDe3MOrJo+/V9hHMJQxqDIW+SREzRLtMGcLL1z
Bf/uQyl+HWxRVWttIRZ1ysrnIwSy2wDrmiQ0khVNrJ5oZujD3POk7oPiaGNF8IJ92uII7YWpMdu7
woqgNG1LJZp/Hb51H5zQFFH6tVFEDy8PLWuOstU/LpNwhmtpamspHtq++rHUw/jikezt+pWEGhNK
lfURRNXgJ0vZDvocaB4Dh8rFuIrFbxGZD2OF4Fd6sDTu9VhLN1rntvZpFl4n/y22lMvaAvocybDz
XrCbDdnObT59H0W4btS7xHoWi/7qKbC6NBAcO7xnNLPtbaSxF5DPLHmFsKb/BpM3q/IdI/cBQtDX
4j4y9/KY35z81BfFe6uc20Q1HvhfHgeqrzOnDmbvtH7fULUrvtcbzJJ5YpJGMdCIWjBw7p+shL4k
PxOiLUsuDAMckrzmSOxBMjLAVSMwhsmXyh34dq4tPxEukl5oYUdsk0KjOtg+RTkiaXamgTDdxivR
1ISjuC9evYRufWeb/2ZRDvUl7R4F7GNjqb12Q6K9KOw9huwrd9k8lRYzHL7vTjb4dYJs9yrCyJr9
zgSFUIJtj00RM2ahWRgSZG55F3UhhcyvE+55Jl73/DffaNL1Wyki8cHBib4PKGnZKd3Ef63gBeSm
p9SLCxoTzNkSvOUNmrg5Lt2uUC4j/SBQ+YD+SLCRH+XVYvz1XH3YYVrmMXyCUzH5Z1gA1LdL+VZs
Gnqhl2/yL+bVAA/aA/NrseEsZiXIi0WY98LhzvxDuDlBMtm+pU2C6YI4xxenDOMm59t5eZPPe3bS
vkvg1E5bqBfxrLDfHea897HCG1YJw0AWCp23FoQAvC1S3KmoFf/9BOfS7vNfkoUulUNv9hzvEvq8
u/oZTa1E+SXfBIiXx2PZ30uYed1Hvm8t1aHUT9h2KWkoqcZJxGLhXceGvInBnQeRGR2Iq6dFtQI4
641youa4NSb7apfKsmzmVUwpkv4uabTsI9zEIVvey5iejFflyx/7ageD/nk0up3GMYnuXg6bUSMA
BpFYm7LmtsulEDPRVx/GrUhiOceeN76b7DdlrxIlnZf6WFu6ADLGSVvn/wBwn5xB3iXeXfN+Hot3
TpEKkMqzOYEMFjflwS5Edgw4QhdMsOSEJsQRhPJ++5QzxfAEjrZrdGzJeSAK5zhbAtahrDvCdWUu
YzbtzWartaydb4XvEeyeJ/pvvQq7qTrl3n9Q35E0mAyfVUBzekUAA3MEn5Tjj84taMpV9qK4KyZj
gusKNIHCrYvrVd0nWb3jKAt2B1QIhBuWUQdYUH/Lq577At5EZWTCyq4OJM4BeYqT2eqbg26LM+d5
2M4EBCUVugBgt2mdPMNV2NRLcgXcTNmk0i6+MokkIWxVyRuFKz1JuM/p4ZLx9wdn2jkVS189JQD6
T/JeMSCTv2xlsk7ZC3rizTX87vIIin8T5XoPh6mpo1RwGCgLWIZc44ug1vX6QDsNyTSiQY+bnGK1
krXMIGUPyIMVqO6LvpP+RM7j8VC/+sWtW6tPr50IvLrJs2c49X0IJNmKWIIfC639hKUqwUzI+zkg
ILwc6wjv2UpdukURw+QQZnUp+B8W/HMHRDlrd3ec3o/kEMu8x8zYThXRVef2V4iELKKFSOnYx9yS
554cdrIYZ1adtV1i0FF3Vf9ApoHCYZv4OT73l2KNdYwY7s78m1JehvxGCpgQbLNshkK9MkNnw0es
mOVhdb06NS2ZdjKTO+XFol9P8vMQbFywFtTqOHt+RkWYWlQ9WD+x+jdNSTBsyEX1RhZzFqElDEa8
lB8PrrNEvfS8t6ffgXKo3MDY9dUaOwPlzbj1LKu4IkS+5DDw0bRTe+rhFUoxjUhQIz5edrSK9ABD
uAVlaNbNl2Pev/JvJaPBRiQNnzcDwAUlJITRgmUApnfyegkUiKdY6klIBMNFus9L2MXzDmqt8ZkA
LuS8PSAvLIduBk4lJfoCaP+z5ORCXnONzeVNyeG50WGAGaaxUKjCYO5nORpFGDTUzIuNcCEvJpt6
eVPoEcZQWaDy5Ihklabt0nI2XOrpvSzU4VxQARm6Ci+gryM9C7AP4EOgiXW5mYq67fo3LGuwRO8d
9u9mIlIeGQ2iYA32eKTgnmyvuKSJt8sHA6iEAYXC5KyTHtrikQVL/mpHjCM7CP3EgxoJfNmgoIik
G5PvZgTAtzWoIApbxotRKaY6vTwrMGtSgRO5YWEcK7FB/JQXs5oBN/6A2RNw59ayZ62qsPvqq/ho
f0/mU2kaY3KzRnHuq/1ICt2T9rEqryZUUEbOp6qWivDEBraVTktsNt3wRUnRR48+KhUvOKB97d9v
RKUnVCKYC6U/wcVAjLIUZKe3XuP50qQsLNncRI9rb1+iiS0yCp7AoT3stb05OJpvlKhIn80M+I58
8RT5FyQr6kxQu4i/qrXd/4pQ8xnMiT/OmyKlPKqrzxKrLuSkIP9QhHRx1Msxe8LbD9MyJrzel2fO
eerajXuCs5FFOG9VdhIFHPGO2jj/U2NkRufoSW5DDwu7cneSG04XiZ7EUsgMlYYHZy3IrHyzsnSJ
CzBBde9Rf2dO9vdL8G1ZolV6UJzxy8q2juYC55sJJMbdzUNUtyLmooejO+ysaGirYL9a9wrBw20W
UxLI5+RYZXF776eWF6wd0Von5eE//BhODpJ4J3sKhBTrD/vWTIKGiFS5fY6lIRZrKgwjziSEqyIY
t88N7W8Xu3v+RHhgUgquAJoqV5KjCslDSVpWrvsmqEnfZ8i0/SuAmrOtX5hXbg6fgd13w3otjH1r
A1adbTky/1JikSrfVwBB8xhXauZal2/oRBxWHDUl9F1lAyC35Vd29RKGW1pwotRZA9/7OCBLeeXZ
o53MfAAV9tmf/P9B5tppswI1S2WQjtHbGF+u8Sdei+q4sM7Mdwnqu6yZ9zqPhCQnsjmKdDeY2xOv
4Yk/ewnfr1E+rUsfubm5FIJOBjEGpvQfjQmPn1d/6ccmDbG0OVQmQ1tilpQ/0MhXkBHmLvGFiVCh
kVkWU3onINvhf1PmB0n0EjKQ47iKWmwJNfvxlh+BwZ3CljkNKKqxrpaG6f7b+3EG3UCk+bkfUyIV
tZIcyZGswukyNxBD6krzMLiNdWuUpVGMFkrJ1e0vNkmMxmmu9Y5ul3J3Mx3nKhgx6+b1UYBYwG0v
Z1nqO/FR6YzDig170l/U3QSsoni1I5TpuZ5vVVYktDWnvyei/oJFH5vXd9mp+oPatJFMAofkeCWT
ZUvmt6BlnM/t+12+keyaQ4Koui/HSt/EwriHhRHAO52zFDxEhpk+4XhT+IyABSKHF0CCaUh5ipL0
3ndcHxAlajbCdfikUEoo/EeN77cIHTyo6sY+m31HDNgkI2CtLgUrSSRADU4a+5PLyB/CMA+G9Hw+
lQay8vetqW7KYkY8i+nB75cCdPoBK/VvtLZE4NFwiZdh5TuMDwVfKXBy4IEnxKItbYKMUexGoHRl
wx/keQgreo+gSxq7Ev6Lycyo3xNinG+YpFsq6jsp3CgHjauIkHvzjzGIEIMSVEpEpDlEVwvQbKSp
LjvFp/fusRJa0pq7Q5RZwU+GkHFApD1p7DnA9pPgt1b+IMb4joSpI03AcaxigQHIbGsIN+iDlrmq
XXV8VX+zAbFEr1sJwnDBla/7fifOj5YDWLRKD38ZXESPRMXosALTmajQBJhxTPO86YFRDf23SO6q
eqVF5yP9nNjq38BhMO3F3oCY8lf35J7jrLSOdMUmhqWvyu9rynOC4+Tjyi0QStFwGBhqRJetrpeh
kst1asqzO5DT/9dw0RlkrqvOv+lNh5x0XdFDmmKKpYColC5oLUuQ96I94RwpxDRGlqLOkeDTfm9Z
VyD5J5fHCjGvJbH+lWGkmZ7GJv2CCniQP91/HuIhPRqMK0ei8zm+U36JQL+HKeVVMc2VIaykkPRE
s+6nMGhxA4BtXLVQjy08YtT482ahNccJ0feYvdLih9ieV747+iIjjXktupFNG+7OPbqYIlS3JSTF
xNxhTzfnnQCLYXssn0RxDgyNX8xCGiFIzU47dxX53+s+izCVTBUcspgEsZp56jT78qmDIXfK/vQ3
yButUh5yclbVvH4njCrSr1uEwp9ig+00LrwDtDGrt3CdSXhTiJNHudpvLm9OmhRIeEPGwUrpiGgI
je90Qrrv3H6GkKioZS352iJfn2zWzn1dds0WiW93zExhtxnDD5Sb9jH6ilDCa7kL8KTCRJa9vXOd
bgw8DfwGt8xy2ENlVJ0ET1pHfWDwrhw7gZdmtkkhnD+TMjOE7wo7ckV4liva6C+P4aHb8QKsudmu
T3CPox4HgGnZII1a1GgkwVIw08vOJiH0oLY8dnqXanyWRKHKNbucKXZ95epHP4szoNPHwki62fcV
0i1oC6oTa3U2UZbaP6tLe+cNsB8HbIQKdw3RvWLUrtdGjDJBuJFv54Hrh5ngF71nLlYlaLz5mvQV
Np2TWuZHxAppTVyElsv2cX7IS3oFe89ehO3wJegn5sAAh0t7yhCZtS1vOTy/UCHfSGP+aRqU68iS
C9k58CUt4qGEjsubCiOVWaAMRiqHEoXW3of7uEwEn9debMD1fCpZBMKu2V4uppCcbpHOVoEYo2g3
8pWgm/kyakdoIP8bMdPgUSCyPXdfB8ot1FfXQ/wZGps2mLBI//qYu43pP/Bi0teutKDMAhKA/JSb
bVQZYzZpwBeMCiqkmFIEXk8hoMzN7nO4DYa3fiYd/cuVYS/6QIsX2Ibm5U34Thfl8ThRpITrLM5o
5Ch+U5W/t9HVHnKcQHzYh2UG4vDE62lZAa25XqjIeG74tVHKJsvGiRZQ580Wc0Jnus9U4yKs8+k6
UK69isyO7fFV2AjbdfxAuhqYH7KP+AD1bZnRiwKMME5tyF5QAcYvM3I7WTFflPm/KDHRrkIseVYh
BKP8HU27tgEESydErn2lJE3cqGojEczJXDx23AE23RSeaLlNhj1amEbHT4n96sVNkDqje3blrGHC
fJF/+Yxv8iJM/nOPgWgZ60cdj1aO2LAVUJbaXQVz0t3EbspzX2JnrUMRfEdYDXqad5IAhEeNrUz8
KbPM88XB98i6CTlCQze9cwH8OfibOP36PgjxVfxiXSeBgia3xPFcbbBFhjRj+eedBH2XwpuS4W9d
idlp7MyuIqunSyndtpAZfw+VSR3D1Fe/xZDWckkJuxaw8UYTClXrmnQRm1S07XCKivBBS61y7DCf
X0sTUZqD69ilwFpMLM8XlPlZSyxzkB4HpQv1LEnPmrHMmP64oucY7Grn4rn5aC3QtWeXPbhXYCLN
DK6OH+JVLSTk5KtrdWUpdrTFOVbkmgHMh7KwL6XxQfXiEbSIHYSPkjIQKworNXbvk26+yVrOlEYY
GxancS/BcM3ce57QYeTT2j08bI7SkTeAEmCS1S2OOOQ/zgRxGZt81RldHsKKciQLwPGvqSjU6/OL
aNv0zB93slIpi3GAeOwPXea0Mv2OETzDsPNEiJN21YVDEswnrRj7p+zW0NsniBv3hxIHQMpIF0K6
o09zoN/LqRk3fXTRXGMHa4EFgMye1+PAmsLJFoag5nqJ/b2B2eG5MnloaAGHazLENn+5zPWx39P4
UOWWPVQpX61U3bnVw5vDraK+ht+vWlzKLWeqEFB01WKYi+EUjLovnvPhrhUnDasXlvmgDoiwwT9U
aqTtx/WMH3j4TBTyrlK0EupzPVHAyr2gIoq4ur8qXXEq9Rfmn+3bfQJKV+v/C/a4izi++R6JXlR3
5Sv+2c4PwtQA2dRYu8Rx1FWUobcX99kCLwYcb663i1nnQATMjx9MvKWqunWK2E/DtcBCdYrz6jfp
hqXaZxd+FggGHjqUQS8WaV608omeTZ8oiiQwOzvWKPpg9SqAMsmS6vpFqcq5HiD+GhBfTT7zcSjb
6wYU8zPU8+UXh/e4+8MrIkP9Q9JEuzB18+ktUJkHiuC1iJHOwdX18AIBPpvDOupzKN1ymKwHczKa
8iS2rgLgkiQESpFx+Ulhoo17ItUGdCJlSuse1Tk7ppJOv2Pe3Tf1YflDxXYY2FlfdQgADXb8+Gdp
SyPCzMvddDJ4OKFYesyigf0j2i+1xZriyB8jeLsybrve0Lmuq2pUqttwMtRRVSf5cm4SZjawd+jW
KqcjER0wbuAHcoIen+uVNYfVSpe5plLFrA+0a/9dAOnaLpVXa6CAb5LsWLWe56kwH8A8Oc/9Axxb
90Ctkk0GORS/GKDiW17Um5FUJlS6LGXQKAf6ub1gdWgZoTtEcesNz+e0rMWasftFB35wHxM85OJ6
BYO2ijVdMO4cOq/kk3XTbFqK0xU845Kbi5Hp4nRKW/ZSeRlkAtfQJgxAuIS0t9DjWTiR4cCWHHM0
4/yTJipSynn8lMjxD+1BHiYfF8PX2cgOSwXQ+kNsl5LXvelFuY2Tf7e1YxAGpKaxYSRHckZTx3Un
J6hBKVyuR4e5rxGCidIO+f8rtKXL/UePZgTFAryCtOitkcP84QayKeTBOsp9XSjGmZlcBTfK0ZUG
U1OeYZPQlrKnQ6bCWeBuitZYmSATUPTNM+HZiHVEK+4XziotKHtE9bqjaxnQCw2DGw0e5DcQytRM
COGfuUhuCG2lFv0WlJ0/PsP5hNi6I7ozhSrMBtq8h1gRAZlkV8QhY0u6QSWuiF7OKQpP384X1bt6
RcaT8ctKdxDa6SCFuFJqqh3TCHAyzX5iRGSaAoH4QOWY/P22xY2HL44SDMfNa6Rz5pnNT8Ckht+R
9WzRJSK0H9go5TSv+hD1CmNlTnNkC3ydS+7wP/1xq4eOoH+bm1EvrdlvwZAR87kFJO1OjABfUGaE
lYimEVDQJZl/NpuOhHl/NAPn6gFJt4P3K2reqNRebSJyVsK+lDSYuaB7MMykf8CxzySOZeFy1mqI
eWE5Mc5Fw6LQBoaU1nP8867ud/AS2xYQckAU0KKMeCVOFLbt5uAfeeGX8O6Q6Uq451OkPEpsK9+H
lubQcQrg428zvYfgTVAJE+NORdvG1jLIjSF7s4YTYfFoMbUqfStjT1CI9+RtimmSkRG/88zAwY33
q//eR57bGj79ZkDAo+61AMamEayzx0lRnyIQStXdywlg8tYUr3CfSjG/XUzPVeEJPEXOp5V+dOGE
Qwj6CexrOshVl+Vl/1D6TudEaquEUQ+uSc2cQGTgT7mBXnxf4k+/7tXdtgxMaEKAzgcCHUN3VyJc
fiKKcEg02EXm9IsPLT4r70NERjDQEMsvv7vif1uj/uDviVzO50W6ssFH/6bqhplXrFiGAzhAGi+e
tULQKbPg0esTfkHCMZfyWey0KSvg+SSjLFaCJcwydt2O9RjLLoGh7nBo+JuMoY0YsmhWYHBb9aSj
iGML+D6ne0++oVhNs88zXdwcgTGpbWhrXIK3C1TNKqce7L6yxYR0t1YZ+cZiDY1dhZCMYdhL9p1x
uyfiGQAK7ZJk2sTH2iSMjsQglz3jcdkf6Ww4+m+XExJu417XYh2mDYInnJcEs7UfnKW/fybsiDLT
OUGXNOKAPJYJe8LPZH2WUYKwoBO8+AH9zrrZSvhH8G4qK9QZMPorGKbQRFzw6N+dSIJ7sTqylyGk
WP45yaMOWNHoZTA12zbLHOXXFRw9zatloGC6LFUFBeAy31iOCTOEqRm384RXhWJnr/UTF2ahW+ZO
ADdzZiRrsYaUHZL01F+pLyCQowVReDBhIBry55L6kgJJ+KNfREwMVy6nwJ0f1mP7g43scthpzQaN
GJWzZI8zwpxYJuRCVjiyfk4kyIY0AjarUGdOhfWPNk7f4dG/HjKl7uapLKs7845aMzGMUzNDrpvG
lx3vmqRkQhRUseOZybYgae+Jatmtjxh7xL8Pk10X88CxQbiNFlrr+boDvXKGX5IoppckBhdG5r7M
syRm6r9HKMFNcIgiW3UwWT/og+VSHFiLhDeK4gH2UWXM2ioV0Ysnh0EcAj44OQedcnLqdMZe9pxU
gZjOlVApOs3VzDOsjzoZwwzs8lLhaAGgfaLk73jE4dkSR/g8M2/yUyTlurOKYP1UCJVie0/eb9NH
j9a4o/PytP/8AtXumIuk0XKeOdaANcQ4ghuQBb6MGe6fEePa8KcEM/CHG1TfSSPrRmlfFSjkam+F
qlnW+8v5vfSWe9Rvf4dmQkU9BBWJRrjmXCfeFA0kNFkBtJYlEvd0RP9gV4//io+rRUl3J3eNg2U7
3NMVyv2fiGOMuMJh5gewMP8017cNj/Jf9dVrDSCFMb6bgtgbMa24XUwz2cBomwc2XH19ot32+NVz
lR3d7tlVXTWFgQcQV8V+hkyuK+8V+6o/BQjaIb0L22nHMSRblD0MvypBNF2h/Uboy6fYz11Gt8VC
O31CkhDzc00bzjxeZnLeClbBalbWezKKReXkhTRhAfqFVxgd19W95vgXejaOh4+f1sJJempSBpbx
dtLp5pcguOb6KKYXJR3fIfQVxYtUc8cMkY0v/e2j9/2X1e1jyVonRYkjcGQCUy/0cjR74CZhGA/s
n8uTliQWdWqmBsb9TCG0GrGASms5iYUFl2nnvMfDIukUD9JY2zHdoufjuB8ksoTR98axcoKnOI7C
900/JjGfiVS7ywuHqW+Zi8jANEbvZEg0J1tzCWuv1xiR/5+UYJSruam9P1N+1Y5erDn9bUCoywre
bURIRwNz7cMgNvQauVr6lAyR4JdL+XcyfwBqmRY7/eOBOstr1yuKcMxOex0/6V7njYix82HcGLuZ
R8ZTG+bpl2hrLUXwuVsrl8lUohbj08mgC+Qo/YxZxTt2nND7FIecl8kBDzGWdni+yhoK2U7YcR8c
qKxoQIApeXn9GxapaOgN2rs/4ZHmy12f8GFtTNfiMv3hiWBLhzAIBe5LJPsySNDfjFebVxPB2x1M
fvVbmRRm436s8qXrl1ukuqoLkgW8AgSUq4kZKOBIeC+XV4oj7C+GN86aU7LUW4k6VNSUm8ODCPsB
+XNMN7GNSWEgKqXtGNfJ+2v28LbtmItbN1S2i4w6HPO6V5VjT/VlS5TYUN8cYxnhwt9kqx8dzeP8
eK4DmBumT/YGbNav9FFORVJ68gvjtxYT4NSmkQAFfX2v6WmGwXZTgrB3XuMFecuUs4CycDpYKWbl
28t70+9bmSpTldyv73qaPd2E5GEO4Y5fyh/AQs5JXDv6ilqXhT4vBuoUWlYRetSzJWIJJo5slETE
9hpdColxAe1y0wRliZPIMV/rLPkWXCExWNcy8M+0mJZ52y2WA82pO69qbsieVuw+1NRYS60VmbPX
b6G3zLt+CClzYc6RS5uyQ+H48iWTwHwuWgxmzx5stG4yDlycXHwQ0FSLU8+7/G+wXQlUxGdDxy2K
uK5b+2DKRtG9wZ9ZuiuB/YzLL4TTQ4myNBaZabakvRiIOUheyaWSLvrt45q9X1ZAN+OajnPGNaF5
XcbNhA5jca2kfB6wSVOBh7AKrbveBN/5WL01UwfnU2aOQ49tmnj1+N7oYUr8x1mtX5A2EL7SV1Bz
PbEcIGcCWY+HQuVy9UnOoBGXW4lxQqm/tUsPQ6MUePQoK6UITPglIqt1s80Uk6+6w4WpNFcA3NBq
rctz0Tu4TqnBN++G4FB0w90XGL0emFF72MDER/gnKss26M0LB+L9+BnV+Kb2ApKAkGbVYXnZOMHs
DsZFDSxPSyI8d1ZP8dUcXnWbzQfVdepo+w6GI8SXx+r3mTdut0Vs5jvG2Urox7ZGHW3ojttjh6kG
HLxStA0I//KsB4+0eMKzKNGRWQjyf3KZDZPpAqLbIRYZwmM8xM7o8be4K4HqF1PS812bnyQQBxmI
XFXQImHjivVT9331Kkoin1WDUsHieI4HCU4PSf5bsAdrlvbPwzK8SX2X9hvIrCYIALSDxPSzDJIS
f2N0BF3Cjy5tkbhX+f6PLZNKSNTbHRIRYfz0xtoJYh2e6NeEGvW6NXh1syn8i5196DiqoAuCQHK1
8G/PUwW6ACNZIEkxKMW48kpvwQQH6+DH4uaEKBYQcCa+YAOvyzS2q9XTYF89NeEwcwpd6z2d9HwJ
9FnWEirDxN3Ur/41IGKDLOrwSNTTyBXZkyq/xiUfQLcHhDBAlunV/DFaAAEv0LqVlXP2CBa9otx9
Q45IqYtTc7/iShGEEJzV9CZ9UghkEFA8v1wEpoJrjvAsEoQLMjpv+KqhT6SsfP6Z/l+TEZNYYy7s
RL9LZEo2ijZL/b2lx2VGG3XvF76IAt5TX1N4BxDu7JxG6Ed1A8hk/GU2SqsdHu1v+RvO7mLRbrRb
RHgSsf76gB8DycYyFTJgPJWaHfGopB2DQlzULA6WO2tkaA6Ig0Tyf0/8Dmb0svdss2GObEFLTBrQ
U3ncL60WdyHmn4sDOnBAKhJZg/QDsssi06NKNdnzfw9j78H9mmIZqYmBkA9eWcSARBMxO5SHot/x
5v6aEmkTt6qKzd6a3sYfm0BDIrcKhHGx7qKvyWFsxp+EDg3gdNmSrimmYo5LAhR1m+MQhfpV5vYi
4Ma8D3DscydiL//cXOEWtOv8zGhuJ9tWMyaXh5GA8h/mEc1zdi5Po7KrAxjpzr6SfGf+D0QzDVQs
PH5YgWoepbjB8MMH/JRKHH055yySgV96H0H47T/ExZF6S18Mhfuj9W6pBXAU0OpiWPHBI7Yiyxhv
g1w8K1f/7BhAOtqjYdsziVM57/cm3UxbaTtjsix8SdKw54YCfNZwYGnVaVVPWIm23QTrKOAzVPcm
n4+9NEj7AiVU6LGkgAc7AGlhoajMTdBttSlCiQleN1RcrT+cDJmfwKQP8wRs8jkFr7tLeT0HtGX+
9MepguqEPvcPlnZHeGpH/KLE7zVDeGljt/N8a2/C6JJxQc3ui49Ue+rf0bly0vOICcQgsKf1/hOw
ySclEgiLnqt6oP7hAfFx8ZFiCfV3MAq+teoZMeq6s4H4rnsNDe5nP8OWdu+U7tlco8ISIyvMjaZz
Ax2TApSSRbUNXf0ITeEoKQW8PzDYwEUi+HbPpUnzef8VpbZdgrlpz5mVin8WXSUIQqI+Gbe01tny
C7g9DgCaQ7LC3C4K/Gu9DH+nNN0VHe2CcdMYwe0t3JoFNdxdKHjghiTxVokGKIqnNMesqnn4fB3M
iwYEmV6LMzEpgLD3GaDm88o70xTxe5XyEjx5ewrG1XhX23sbAqyXO+ENNwVDaoh+y//sHd+HugIz
IORCtHWYeIBY69XryS85GnvURrwLDzIBrKljfJ3L8/P7eJdAnQ2vfDtGhc3Hn4KDuC763j5lIZmG
VRfsPREGDrAk4N9MOYf3M4/ECi0O61X655zz+dY+kjB4CSe3V2QQrree6/vm/TURFry402VeP8SC
gZtBb9cns7I3jCH8jVyyQBp3dmaLYYut2fMls9FB1g9v5BMnhVysiAoJxIkKI5pK1XT7GhMquorx
QVJlZVo3lESyXcefAlAjjmWVFHd9JfX4hakAwBTjqZFSdJwOC2iQg3pqMCxCZ3D0zkPTnwhLjxOn
oPKorH9ZLy8HudV5YCMmbIGF7zndmAjCSdrpjhm27GrizhCab3w2Mz3xTaMsvv4pqLzMJonGlEt9
Kr3NFO2w2njffLWZur7ysrqarR8ekyVEjek80QG/ExU0t1oapqiQmLPS5bE+K7zT1CC6h8NTDJfz
7FMyIV4CSmCFrANzJo6ktoEFkaNzYdPTJ4hqR35DIuYSfkRdSzCq7OezqC4PDSBnIrwagj0fyNgj
H2+8oA6+JYvO7XPLXpqjBoUPGTuEa88rGw9pSllxf0Hv4qlvaeJl0wbbxxJ6znSU/S+xunDolYO/
9kWDVWEDGMIAoFHs7p8EqoUW+/3bl3FzZplDvY/xgPvGCHYFCaKOk0bYrExHAevgbu8kduLDdZhW
mkPUrvpSzHGcsJY2x73dHczVc87B4/JhA53ZjsG6mJe/rh8p1oSiwGhZqVdsm5Y0H423axfB2MrL
dQ69ph7qxJdumB2QoSHLa3hEAjKQ4TSgRbCArke/jgZ+K9CqaQcYGXp5F45shDlYhl7IzcmbGovg
n25UGSAcPoGqjER3IfzUtaJ1acVAZ2PMr1vfjChKMtknTr7FhNmIUVBtIWZ6OVZJ+PeKVeTsykwu
C7JrDQVX1yGIid3PKRXxUkcFY5RXW38Uysj9li8IYJaTLZBm70JAoVv9rEQccvS1g/sayP06jwkN
Zre02nnwmNo2A+OYSmF5J8AVxWdvS4svjTtjjSyX+++XzgtR+ILQ59e5b09r+JHmCUqVoGgfuIb0
JHA4qtjTLgAwkEG4ExiY9jpR+YS/FflwNi8V2j7N2m0gDDA5BkLx+EK+rbvF7XkBA+Olvwao87Gq
EoXfInlKiqyadF0jwm791EYz6DyN9Vu9ru8c2O0KA9Mxcjrz9OpLVAU5zN9aSzIl2gg7YMaWmIjI
g7k02YPNZZPEEKpwHoJ1kxnHCzslVZmjycN1mj1LvBPGfwSkQzOF+dmfEa70vCYqbQ+MITUP2NHB
IItHXGtzmHKzKoVKlEtlw0yKeV3AhrgQe61NUQiKV7uDaW6C9K5nSmrPElTNfv/GLlp4ogIDaUv/
VMR9ZSW0e4lajl84hWeJsIzdTxBbWEQqsqgJsiiBXk/m6enwqE1IG16rd2PxEr5HStpGxCMnT4sH
zaj4SuykXcg+N89FrtlpmrY4iiibJVgtiRpXz9ZdmmdkDfUcSt2SG6xiQo/4pBC9IhNbeeRZoor3
2GQkJODCaXe+2Z7lGnb+iNsSaSdsloeOK7tbAlCGwZohGje0FAOwq4KRAxcGTM10vJ+3dIVrSJwY
XhXk9H8E1GuG+Q0aFht2lPkVvOGcu1EyL/CSYNwA7MA/uS/SYUmaGO3ARzRukPUyHty3Y8ciYu+W
37P2HqEqQ24r+ZQckpJClo81WojZ5/PB10UBe0WTiJDKuEZN+nQxFxmJtmTzyRxdLs3gLfH4uKzf
G8A2LxetIp2c4MuNApFVWZ9rkI6vOCnRmMubL5ciqWDAkwowRDBzRDs4DBpaq8yqyMxhJ0lqIjTG
LsgP51cge79h+C0M/yv4/5KIFzAtr2Y9xDY6Z4baJQrUMW2fEt77y0CfdZNAg/chLl/dAyejKfbp
RsTnuhoNg5RM/uwDpf0Du4fL5aJwh4usQsG93zwlOHAJdk3oyveK2wuTg3p3A5sVRk6LkF0VI3A7
ilWASlx4MZ50Z69SncCJU01pFmnFdgOht9SzFhgWMrqzjgGgyMPJPO4ML1/Wkn2XxHUV2cvQuaZ2
Y1ZFeZ2m+JnxNY/vBt7gax9hiRX7xfXET96AVL8KX/+8ZkKbUz14oH1CXrPIUzO44yxEJOvM0DU4
SfxV5khXNEYF5jhBQ+pzyDMjzLLRtoLz6ILN2UGve2ZKwc+ufRykkncPo9GRYUqFwPqgIm8WJrSa
wQcDRb6DoxO//GyrapjKCVtr7OvHwLeA/8sHhrnei8VSR/nI1kM4zEmO+5+pp9Smx948JhgVipX3
seHiSIRgh0PpPUhO2Qo5TEVEjTrT+WaULWA7AM0Zqscba+/5nidNSPNXW9CAVAb/L3e2RKNnyZol
YGMUAiCxVyH7LYrpXauTlDE/6mBqnZKX6kkx5VWU+CfbSfT5nL1WIeewNnen/PvxX0rrnC3K+I3k
51J7Oc2KuXiTmg1cp4uEgxQXJZ1m5ufUFTqUp4I3T0uOXPMOQp1KfJ3G8/oV6js8PVWzUvASnrqk
Au7m47YdFiFEVP64ZUUlEehjZ2x3HWxhclVUSxa3M9sMbz7bKP851EI0Hxw3zs4Sus7c296uzQxY
smkYJb86SPlGuB+ARM2dD+ugQrEWg+kTOtnNBXI7BNVYr3Zi/0LjHGNbtJFfl4B4aTBFatrd+Ace
OlF9hwyh4wmUKXu2o9aTvBVH1G/69dY8wjH/LxqYHDJZVJisxgxgny+YqBYsffUIje/v/ryaZD1I
KBF6sE/VF4sUHcFIvSplJ6Khv/CJrBbTKpvYACjthnELZ6iWOO65/F4kwUAB/ODRAN75boAPNzY0
D2x+6+G68vtp9F1gMcWw0uJPz0bWOA6SikLUMCerJChdsCR81N8lRur64N5uCK/lnvhN/MZA6ya2
3dkXZmi4ivaaNA0t4E8YGXndzSKehJROJKmhPB5HBtBMlFN6A/LL6b7ZzUnt4khuz9HooID3oxjc
3+xW+Xiji+P2yLpsKMNlTUcXF9RhGGSniTNEP+t5A8wkl8bfjyXZkRHhHFDzxpOMfkf2pCKojsUp
L6bw92bmzEy5SWv+uVjwaBZ0Y2qs8DiUdY46AxdZ8hUHl6MA3ZMERdz1CKphLIxJVSaUrbvpzKu7
wMjmt1hdXMjJYqBv7EWR4BXS8Ds3u79KM0huMtBOchbwUb1C9q5lxA2XTcMkS5IjrvajvEKAWFU/
N+I8Hjr9l5P7wtOAwJhG7uNORZzInSdfo5EkS7sSBsZ1TSMP3A1/I8PhgGdMmNS3CbgoKvGE3U9Y
OrF2eg3IzPwKixAas8QDIY30o491uvRSQ30t9EiUCxRceQpFLPq2ioZKxe6aXvhznp4l4GfCE8J6
RsyEtzhM8ZJ9VfZLw4lTN9Th2Hn6tEk6c98YjQpwY0GgTR6JJtwblEoAppF3FhN+EwrPj66urd4B
e8pT4GBZ5LSp4u5C0FtQyy4/vNkpfZIsKGmiw1JtUrePIEHbHxkGh67IzGkAcQusKVuzZiv+UZLJ
C+rywHDlkgzxEZu74OZg+l1+/i2hasF8TQykZTqf+6Xvwc+soGJRsOATvEDobw0KxfqSOLvN4GO1
k+3c2n4rSOO95dHJkX2dc8jN0+RSdju474e6UjHctc093jswp0bCT9StzA86C47YtQOsG0HDcjkk
bTewP7s4rG0Oel1TJfhw0pFpB2BHuGMbtQMCSdNsoQU48cIwrian8EEBmr93tYCjpU8DNbtWR7DR
+oXRmCdDmnZuOTzH620VXTBuVxxc04q9DFtgR4YLSUq/quf7CAiHzXeyfOrqSJvJpsrrdSfbUVnW
zuDw6OFbaRxMs++hRJoYqq1jcDzQN349F9xqjM7tWKX3cegxNOGEsuzCcxXWuhJ59KnpiF7XkQMC
cQJIhfjwy4kw5DxnGCOR3dFPUkt12mIYqLoxnRpMBwDdnytL1Lr/1cYjBNFTqbJD/g7yf44MiUQ4
nAGgRBMqYQ5QBbtOVXZ3ZuG5vrMzzP39RA8tNggSoQcYTBDZyzsjSjwHyJeDPVToDVBeQg3gtqT8
PDc7zDBMYFp2Hr+UbvSK6zynAbuiXtRbY3/08UFCaYK/PBmTitEeGlNo8GQgW/91kzi1gpOKXiDP
cIZByrJUhtvIj3vUv4EHdLteMUKmedf5Ozlb5m/xgsdFEkXIs3fVYJjccL6gWExm7Ak8MvJRYTed
lJD+Nde3IzT3w9rv4S1Jo67Js19oQRzoFRn+HtB8QC7qLZaQdrnBSVExIulU1hB8hVYJ1pFdASS5
kj+lIMedrvOFj/iNXoAshH+yKPJjiKXdmfuwMV9MF7IPko6gjFDQhp+UnLZscnSgFT4yabpZ9D/V
6VS758bLq1JAsK8sAflNraLQgOZtSG4vq3kZJpk9R7fqhzPaoRtMDLdGOxndpx/fsZsr7bF9xDHg
tuC/BzfwJCIfSq5ZgfGfP/s4dNUWIQWVMmgnGbhXtwwvMuvJtDPyjnpccZRDjX7hUxvlHmqMW0Ly
9YJvMhYAUVs89HzAi+NQFiaeYgeWdnynybUmzabGf4S+qSdty35qEAoFwKrQ0loceuUV7abSSeGA
Zeejx1RISfzbwDTKba/V4NAsoABzxz2LbCYI9lJcma1oMqEbtF8fQY53VlTMVj+kNTH3f89iCI6C
iF7HBeZY+V3m/JpIVoCQsUo03sOXyS4lVa7C4hl+vfRIJrw2bNoOfaFp082s7DEPlOP2G3Kn44MT
GNLBpExtfMplb1A5v/+4CXacdTGSmHmAEmN65Bi5b95CVYArwYUSggRh9WELG2BJn9RsyyeGVZ3s
7habwxq2bJHGro5TRMZtv2oVzUaWgvGQs7uU1+pg/Sqkgv7RDKhPqTuD1RXh0BREbBfQqOFtT3c4
BwUeWpbHCrWRyP/lAykQxz7kwUdERCWgm14hgWpMjq8PhcP9fNimDcVWABhkM3ysFoxZgy88cFmX
a5ElVm/H27ElGzhVL0KriVg/g/zrKro22eWW28Wz/xgG0qcFDXMvsNhFU9fAWuhx0HwxKlfAvdvn
4COcS9ISJfr0fqNMboxBXTy3//78eA729K1Dn90v6ou21qmFOXMKX/Y1hz6Ggt5dM5bZ/EM64pOl
5CCBI/2hgUGZ6B19ZlCMH1jnGGEaAXA9v9YHfXQ/tabMUYIkdHiShtqNvXvvDBleifeeSPMs7Anv
ClW7CmAFSVs7lSQx2dfXy3jL3DTHbgJ2TBUCt4f3O+gCV3dmzoQIpKreBTTn8sGj1rXrBkBo2aKT
1Vx7K5ZZxQmCbIirqkKfEoystfbtnkCcirD/tliEnyilgiYOItNjWCrlcO7Vb5GTDNOr3X1ZRQeC
XzL3NDRQYqLmKUpWhDctfHpYIToys9gLwou1oloUK2BvzlOkXrRTWzrXecbiXn/E7FqFKXUfxc8M
CsQ380RyVDjw34sZCWom7Jdnr3GljGzSc5iuG1VTgzbg0z/IoKdkOyLxVmM/nkt4mEydQkVsVyW2
PDiOvPLLTN+Wyxh1F8gFKogyaBbnTLZYVgKicYUJ0/XAidr1jVO/MnPSPwB19+CVqAdFkkEZDTNg
x3cGQ56KRyZRp2+Ef0rEfPDZ0LvsFmNgUzLpNIrNiTSbHcDIDhj/IzC4x3UMEu8AEfGOwz78s08Y
Iqcm5NVOVUUJArEpye8UJ0UJhE+FVGWpSd0JjBdmWy+rPcCWVP5Nvjf3/KTfU/rQwK50xzw8ZRW9
eFC98pp4Y3glVd/AUe+ztHBtyLKt0IJwKNG6Tmc5UVZ/5nAYWj9PDiFTcBj3KzpPFwO/vyM6y+EX
rBw2VwsE2mizIMiVTZfdQbgykzCB9DYfdiUMI3XvGCjafBJhuzWHWkHHfbNQwA0pENnlv4u+cdG0
Cgn+srmmWb2alqZea3XZpu188zhHy/TvuzmC11+zPok5Tze3HvK/cVi2HIVC1PlDtHTi8el7oSrr
wbJxfjkpBeZPq94KIpwbfBk8g4N/HCb1yWgMVnxX1JbClQjYpILspTTtI9Th4jAQ3JPC/9hBnfUF
YMqg7xoDMgh58o4Yi4xoi8GXJTcl/BdJv4oYuxUtdQ3k96RvUEoa3WoMIwfv0mFZEKxcVPwStcpV
IkWa7ABs8GfzMNifm0hfQqVGxvWPvy2GvWtNT+GLX/LEX0Eekg3gnbRatI5Rz30hUZX4Un2+WDPJ
Uyty+dOmeQrWddgtOZRiZaeVR7+DJ05824V4sfHpr2yTjlYV1LBpRWDsXbNr72ZXaLIHTnLVipkZ
YaBYSA81jtPea5MDjV0GO2s0Uyb3B8mKfa76UT2OLPEmmcgHoUfWQlcx+jCyznK4pmlE3YxAtviF
8DJQUViy/qeSxcRCqcKdV9VldSqU9CVhJoDA65xzKM2nWnINLYKgVSX0RSeMzo9sKzLJXn78R8fC
T1cEt8Idze5hblB1q+05K27fWIbS5l1XA7GMBxoRVtnXrf7JcTVpidA2ZRI7G0n/d1PNtbmuQR+l
WmKSpRUFVXVWgKIDpc5j5RoHwfGaBzZ3HPwPCLbETmxGWHdIqbmZ4QNENEjvJp6ckUPL7oBlr1vR
BOeq4T2Xj6ZzKVo9xf2FR4XD/DCXKBBJBG4m+m9HPb3Y8G9dS5iyD/tpYPVSug4A1AaWqf/++DKV
847rIxSOpTngozMQm9wX/Oh26bs0Cj20gt4CG5PH/of4cQtDHzvJzv+A5WcmTapulGc+5q4gfGFW
Z6yrjzQpFlSvVBiKvhEGJb+Gkv9RCvH3RFpK55owFszKKeAolC1ppYt53g23APuMy8cM6aFJnLeu
i1onva9Dw/SSEOZQWD0eh5Z43fRaVkKge0FCCrUNL7L+x9KVFnaJcKz9E3763shqvsW7orQnweHG
BqFJtddTNi3ENDHEGKqxfJ4fIExdV1yFLgQ7d+XqB/MxSPk+nqSx4lzjV3mYRIIfXT5QRmMCbBE4
v694ZeL+fQEa7cdZELp32YVRxXb596bL/sjZ5HGAbchEK2p7oZybf3qxLoFHM9rVjA+XmoHlRV3b
tFax2Xtz3Cn92t2vQh50s44FjBRwFIBb77t0f+laTaqeHUok5xuUyGNPyrLTXU8keZyvBRNzYiRS
y2mJmmQ1ukjpGK0fdq3RE/frunEfVaVlq+sMqP86Y3QCW66rSJknrK1Hi1MaMy94pOHCFD0eYIRA
zE6Tr8EAhKWbI/JWkWd1aasASxo7CEguCqW6KqHOL+UlDwX6G5IEWf0eEJvk8SjZJ8ziiEbGo4aO
/u5N2j7WGWeN6nUh5zmRV6VTMKZZSa546jUAkiddAQicqw1oa2z+AP3oXqURU1VYV9Qpd0R2mv5t
QJ3IzSJ3ahF0SIMOf8Gd71nNDAlJXzWZgugLONI4i0sb4D7gciicNDnDJ00g+9ldP9WFQDQidWoH
OYd9D/MMu1TwQnR8aRxD1y+Kq6v93R6HJGzo/FKlN1d2LPLORIja1vVpNl5k0HndLI3ULklUwAna
F11cXslvIlGgH1xtwGF9Ikf6M6w90kz8UkhZDkxZ71aKn+QPOWyVMqxWcRMk8I/OI0m1fR4R9JpA
Bk+q9WqFdnj2e96p4txGlyJWUt7nwYzuD4j3n/Z6OiURcGB3PSxpbDonSlnvWWq1nlLB7rKay/7N
N8y1lFreoPlM6jb4tYES17nKzLcxZC6Bap6s6cqiln6plntSgPMNo0RHNT9YLk0khOXOO67F8kxe
yDWK9K5yWnMVvpVTP2y+RjHKpENHqBl67FFe0QIT0xAT0p+vw+JIIvLxcWBQZLX2l+aikMFrnbZ8
q2yJRjIBpo2T9FKcnFUs4BGHaolmPhAI6gZZPApzS1pS6w7vhGRYjIQNEzffCn+AUuRmMGzHsgeY
/s8Bd5NVIIvW8wPY/bcYoOqDR7GgEWdSG1XAOdP5D2n/I3o/nYAu3MsJkV12n5XKWI++xDj5SaQh
CyHZQe+7RXRWhmoXip9XzyogRsD2yXE/WzSSWHMw2xKrbxplXe0W8lLyaM3F++wu/D4zet7EBGXr
xyAnBKWN3ND+81MerSmzQpYDgT3rMz1ooev0w52qBvP5+tY+9uRLo9xULyq89bZbD5CxbNv7mNdb
30vJaX1FChzNzWPy+pYaFVLns10jGLh80IXO2qoQ8jCq001f86Q6Qex/F5HwzdDCe0EWOiP44PrI
8RFfS43JFp0VuWCAjh4NYqG+SVjThuI8/f2ChxdWA8ZbSAGXFOcvGvv/ChFrEiIcP1pZgU43v/Ny
gT4l6O6a6JmGdhrKZcTwXQbo/Z3fTPxUJcqzZ+SBb39AML7cmJJjZsh/5ZzDvdxs5P7SOt3EAv6p
2FgVVr1W5/KFLqKCP4/BVUORlB92Tl8pWprcRgPGM5TozmRuVw87GykZzkuaYGm085UiPcpeWYPP
mvUIGkg8AHGIJSE0pkbBFjlGoLJABVeepKMp4bx9CfPHv5XYshY7eRw2Y85JFpzSH+67PuDj/SIr
eAAfWHSpRPfU+c+ihFAz7utNTBr5YbrHe0hhuNB+xzC8CKF4uD/Oy5VgyAg9E6Q1nABvwwNO9gXS
ueACxUsJqd2GEn716G4i5se8cphwts0saRRxHyp5OCEZ0m5xpTLK6cYtMcj0v9JDZmPxbz2reDgT
JgNAqyeQxd+x6X3tzpm9vLsACZeYecHbx4Vq/4ii1tcgpIYXTM3BsiAUuxYj17BgLbbXt9OK4cbU
YYXkApTmB16xfEp3ObF1xmssIAtGOcQ2N1kvO6ScTmi4lLnTnriS01vujgMhXpI8885qfxJ81/Q2
s/s9q58VCU50G3ZPH8MxHiPrtXZdn5xr2T3wZPCsqLkyYqDG5LLZT2UKCnnH19Rw0SNiclhhopP1
ZxtawJ81qavuzqLgZUIkDjtXr6JZFEXnoc8bTtypeh0xrUqvAQejfeT2+1i/OZ6kWEthUgIeRCjA
+303wRuZ7VnRMgZ8z2KhUNZ6Sqpozg0drttTBw9dDULMGun1MkzP0rakeSikcBsCGLupslAsTI/o
Y4moXwOGL7nwsapHr02sL1uynKQnQ8DBqCdF5QC0g2OhFQGFNiMteDAne40gftHkvT8zR91lCdi+
vmc7d29UOicQ4In5rWxzlMkfhvP9IvXR5dhXx1Qz2YrGrOvWASpnS+mnSdEwsjRkJHV0boRwkcMd
PtSzN2j3ECFYdFLHwG2oJKJj71H8JPNSsOhyvj4kDts+WbzrricIdWFsyKSn+1fcFxJ9w3dc3+Y5
CmOPZZEawdXDIl/hxeQtK4IVWdAXWB4a1G00rdk97UY8Ak955DzKB9oYaGa6ZGvhR1RNsxEOjO4/
U5pmApbFgB9UZpshH7bx+P/RPn1sxlaCEQEFuny6ECj0iEX1NmRPmEdSBXgdKYkXjQEoF+KSzfM6
9fqxlqbW9nUBDVeDe/a9fBLDrd5vJoG1NF9VfTUiH39jasdfy/yyjoFfr2GnncXPUEki5qkotWdK
wRgZYGVhtfxAF3VVsieRuyFo0qdGeI/3Ly4OKiccfkUoOsltGNNP3YPTLDlNcwz92OPdd9L1nIJ4
2EmAq3FZjXsTrR3mzkNK4Cr2sOYbXDFpfNrbhRK5ruqHSzo6KM+AwyGA2nLKEnWjkJs0zNNC1N1f
VN4195lPsSIZUt8sNHLk5rIRL3X6RkbXzqDRcMb1h2SZYrEmD99ysYFiY66FHy2upqkTt4iKVrSH
APurseEySWi1lnCUagmqsYig7ldefzvt34EYQ8dBcrXiB+M9n/ktkMSsAJABqdkH+JFkADJDDnjT
nDa1bX3sCAjnm20N1r4AZ7dMkRn2gxAC71GWaexe26qfOkEc00fnJZVqREVRHqrRsCt62NjqqazP
QhjSZkSaok4n1oyQRWXnxdCCMywnkNlBhHFoQSKBxB28CmrRArZ1JLUc4MhRS28zbX2C2AxrtbyR
Z4HiU5AmYCXEbAZ4V0q5AxojzMYxm4ICAwuk4ONucjpYZorFSsoH126tdsMoS6a3SR2KSCSD0rqt
QbyTaqGkhjuojIz/v9+3CzcdUX8AHuOixt+APSE3pQRv1UgZ/asGavbNlUyVas5/8vbt6Gh4grhZ
3MtE+Q2e6YjzDkF/0EBNYWohBtoXS2AZKTL2NxixZqmJ46n7a90Cam6c3onG3mqDoS9HnYmP0R/S
GSH8vW8jsLcK8kc4MKtIiVaiMvq07xvBkpTvHWWrZ/w3IdWR1Lj1P6vxX2Q8Nq3o0CcXQlYRfdG1
nkGyirg4hgecbTAzCSFTiHGNRc/35VUhTiNMZsPrkU/gS7FHbRWUNSLHoGQ7MSjgTXTxjFXx7lbo
EljjdzKAw3BB7z2lrgb/g3gVPGYZdEq+3xxuweZHVdDvNjmR5P9K+gvPX7/qQ91N05QWZcpT/lEV
5WcVhfLTb9iliVQj0q3XLuNbi/OBrxna//XLQ0GSZx6Kh3010wwYb5jARKoUASv80ezDg73MWYb+
xoaBuitujobaI6RIlqoGxzKNWpfBGG1+B/fVyv0N7U9vGakkYw5JTV9Yr/JrL/gpGvtPTCfysJpA
kNlTmbvdx5vE4DA6+N7FIMlIOR1NZAYosZy1WX9Ea12AYeh0EPA1I/s+euAIb4iCCJdtGzt20FB7
YRUtzN2Vo1y9ba6UzyYuZrAohHOAFfkuMdMoRDDnfA0dCCMzS9qYSRJpcO1quHpDRNodXNQmJ5PZ
O3AV5cCBBdDYhV4+3ujEMRW0K+VaEcyy26ysJQ7LuScmXE/pSa72wpXHbq7oAeUcEJsGLest3yNP
aUw+kfh9hHOj8fGHPMa572BTvcHTVzDQwwEkHzm0o12Qb5XvGNzYWndXkFw75FY/eiSR0HHx3KJF
guIMXC0+JLSl/+/J0Mm32CjnTmZi9b6DqXOTQTuUcMW4TAVStzNMz2n3FNtMDFBv8gSHhfQ7B7r2
G6LD1xApuo3WDWBLBbDWBdAnfu4zpwMDZEDWBC1frxKA+9JgbcAZJF5B1AOSzkw8ktYxp6GQuv5I
u0Y449iIf0k9wal6CVLRgTnG23Nz9sCkPwgZWSNtS5bTXbXVIwfZkf+C4B+BK2EEdf6zYj6C4QA1
aqkCZE+WiyD2jf7WF459ggWmZH3N1hrDgqsvFucHieUeai9EJSYVzosHEi9Y++DljHe46T0/dite
PcShssOEbNX5PwBKwMYGU4+UDeFDxCUa0PCra2f7UWkv7OprRmOToTfvC3CHszHvhfc8pQZVWf2Q
334dISlrAUcdoAFbOornARVeZEOZPBwoNDpXybBVnDI2ZEOd13jG6Ab2Q3Jk6TrNL05vD9ImEdI4
KMuH7XeZmOM/y/n7/LJjMNYl+kUgEDnDZOGo2f8b6Gs/bC8BxlaaJQRQuJp9t4dg+LsrSuvbWkep
qR3PbJrCHjpg6dqSCMYo3M7h66daHcieADcIWVUMvvLk/ne8h3A+DzvbUxlRg5OhOLvPxb6HQNjx
Qm17qb9Zt3UysOdeK5vi2cXPHZGp3qIxMUxZN7gw2Zhv18DsUKLElwL7vEPnfaKsjbbFJSWr9hKp
s+BQzehH6OKWkKBN7KYbdEMNPKsKvpcwmV75OZSuci0LzSmckgXjlXKo6uZT75T7MjirWQASYDnP
IxHY3RPU/rEBuVCQ90aC7fz6Z/SLaWTqhHA46xVcmFvQJ+feLSwfS5Li66Wz/sZhYRUjWIw7MDj6
/DNEuuXWlevyRekfDNaImDvl2W9zj7Z8NoLExbhVc98YdCdb3wBUvdXaiSzuyVimTbYVPiKIIz8R
/8gOYwdKl7QB3NG3sD/6MzgWWC8BEj6A7SD801sFj6GX5zGxph5l11oDAOW98DcxWjld+mkqkF98
WlLx0Z7vw8A19x8SAgF7ZhDdMVBMKKgspbjoAdtdsni/VHcPyYyHMqBOLleAGCqQo6dB5WKxVAOt
bFAVv2Laq9NOYPPzhoy/s/cO/LWI2mrY0xUvVRxjTMPU6xLqvnJKKKfcE4v3p0QkcQqJzDSGWe2v
JLfQ8ktKARtnAaWhuprfY55LDR21rt4W2riueTjQGgZtnWDovALKeMA4jDTnzYQZ9SjfBlu//1Mg
TG/ziehqjSfL8tdZBsIutWF6XvzXX9+trgd94MRymmC17Lfvwt3HGcIinB21IMUgjBeBF1SMDSxq
b+X8YHG0fE7SKqJEh9Hu2V6PmuzB8VaDAw7ZJCp1Ph3nMtKUUn8N/0p2oFvN89IOypWxY9Lc6pKs
WJp3xsS3Gbh8RA5KMZapV3aXk/yfqgPxJsFLEkJ2Q1o0ykUttbFUvbJ2O369Us6xt2dC5O3yqBNh
rc7clHZb/ep0jsosvcN+wSgDtnJsdXkvupZecemxbGJMhyyH47N1rYl2N4PEOqg3t0i6l3uS8NjT
P60UrwNQ6K7Ryw0AjD/z7Y9DtGU0eiqGjdawauNbiqG/PY6Yfuks2tsm0Uqw+UneqYGv2L9NOYX8
c4ccL+mkaANHq3HxoUgOCnNK6JTlHi1lCqDtt+B1bvg+wOBKcI0U6PmWv0sCfbP2iJ5K34E38B1Q
gQ5YYZH3wLl0J4PMjbuxiT3WB2IXtaiWzXuX35n4SSdgWA2++bv+Mwivuwcjk9cRLu5Qs+Pctcg+
BMEmdUAv/jkbdSlcEMu9vUmp4DUfJh3kUIOdVjCiSbN9rI2tcN1VESuNGWfojlMyv1xTlbEKTPQh
tOi+Gr470DYMH2un5bJvSNFT7c4oJz29F8Mxm1cofm0hfEaIYUDeLeT/HuGnnw6DPn0lNClq3MR9
VT0zArTA+ehxtQkQSwnpILfuoLsNixtAJowrL7Dx+X+JdvIqM4IqYDTmb+lSYyPlppdKyV5ZMpJG
fzXE1Wksdk4tG8nacQpoerehwHNRRemZXBru+Vi5DlMMzN/96R2V8fcQXM399mT3iec8s+i0Yd3e
M8jBGZ1O05a/uZGTZ2ElK409gaYWBCM52WafI1nJ7IA0mu2rKL6gHF9ElIWmhw/imzo/Oz5n438E
VWZGtG/B4kx+1zGqDO3XyyUhrmgf5vtDvDyaF3PiUBtmxYAvLPR6khtrogXPBKro/8uTWqwVpPKH
boFvlJxyr+Tc1Scx/FKorSR3dxhqx7aOt+WNlO7hlu118XNbh/OoftOGrwfiQ6TVGkbva4GtldnM
XpW7V90StMFqtncQoK7hu3cK34u6XCuRIz9DkXOTBsCFu7egzvAxvNITCeHKJIXCew3HkaV5FHay
6JwOGfQvVsVL4WaaI7Mw4zV7A/oIh//29QmdFifs+4VeUnpdtuAaIih1Ag6CsiYp7aK6WxQWlQ/q
iiKs2h0Td0y/XnKrTa/1OHT8lGEXPtQZyIm8LJr4jXoQ50tJgs73LEZmYRvDwZOYaQPuz7Wtl5ri
F+5KYa9UDchxYXR0ulNakff3aOIXtGExqzXbkx0CvleuCTXkEB0guh2SfxWEJxZRTLaLS0jaHzwe
0/c+kf67B0uR2FmqC8UD3Ukba0vLmUG9jKZzT0JlwdSn5+KdXcZDUmJDbaDPRHgzfHb3tgGaq941
e81DH2snoK3LwEZZZyW29HHbmD357//I9MvpnrawenKlxTFNKntRFdpBW9NeikLmp/ety4Sg+mfR
fJJSxsQb+p2k3EAelO9BUoEaQ4wDTBr2uoABaCkf7Q8COgq165RV/SIFYPRkRLwxJMpKN3/1af7u
5CDtR8XtU1nr9b+nh4Hp9fPgR9ty8MAqzI12w8P/VZPSg7/deEP2JQ2JgJ1rgw0D5lVVGT2B8/uk
1owD/TbcPpMt6Dj2Cbeb7MFpnTp+DyLZ7xrz0z15McXsIcIJn9rsjEuCeFveqH6uSVRdTBRzGtrr
AIsmR8skAZjDp81WFJaVPSsca1GErK8+t7LF2nHvKivRgjPHYgvk9rsGZNjqUkVZju58E7TgT24F
A9oaf81lQDdzlS1zOC0MH+6Sth0OiBKH6otr+18rKq5oSGKeGQyBy0HbFWmlJYu2amGGRqCWoh8t
7pHIAy3/ZWS+TJKJrDQU9c1CGWYJyg0tbFXRaZ7hxFPy6LFGTkrwQeHZTQnACUzhUs8Y9WH27O57
MfHqjMn+3Ma2WrE5yWzFhs8Sjq1YPxY+D/hygOPBi7wGrCnZ5hHadX0GfH8w6G/bnj0zLRucKRx4
yc79E/9ZjAbvp+8SOrxsZcO+Ve9dQX4vbMI12qBWvJNNinOs8Pe9JcuxHF2NbBg8I7kOBwGInW17
Y+5Ve2nnq/E8EsKDEMP2VJoOQu0QBrJcWugHgBb6BVuV6LX5fUSlxRcNglJH45oUWvI57ZOrYtO2
szUihGCPfeBFgBNQAc7etsD3mRghn2Z20atg+GZ4iy0lMeOCQV70eWoDC4JVvD23KLFGe+LKEc3p
d7h/EQO0f9dc5dn+vms6DH1y2tRAgv/r5fcJhZFjmFM6/KGcGVj2K93lGGnxH+eB2y6iDKXOSYuv
xWzOkWal+C29uDLyFo35unjMhm3pUZCsBeFpnCUtwUyMwfCSifjeyQL29v/UKvdDfvNyIvE8P3AL
tiiZLEmQj1nO9p66C51382RkOB/wpItwcDY5IfVuIouUzOGQxY/MDhJTocEM1kmJOQA64iLvluAD
GNHQVqvY7hcQAzzTDA2EP3U+v3UYw7KBd85r+nWj0il2HX3Q+8mrcceSuIUnDaSO//uX3PLxldJL
m2yUd3ASrlilf6nQM0krVFJNtjajDK6XEd3jXNu3cGKEPBW+wgDUEkRWQ+AK7p30UHsfc2DeEV7d
slSITvugE9Qp8m/ARxNie5L9vNroJDKnsn0ppyY3oxY64LWFs9TrlAXiPsEKc8YAzZ1FbCoCOaKi
z4MHrgQxoZsFhqwQuQL0l8xWDLGUxPKjuDDU17UOTyZuPrncTRMZwazD+05NrwoWMtrPUdrxwlI8
zT+6m5LiBKJPJ4OUIN0cEzsay40Cet4IA1/0IkLhZeKChqM7OkULzoBhwJI8VApheK99QfgHFlyn
cgw9C0/zFesYfMt41QcY7Y/jP5zY0R7BrattgeSJ3pp73ICyQFDViBh9goIromQh5sHAiexlttDH
ADPZ2MHL6a8dNF5+Fl8BF3JydJJFHVZ6uuRinXdPgUdGftDazu8EuxaLokOND/UST1sFAnt6Ldv/
Kap6j72BlAWigzUmq/Sr8m0QvTPiAulGLUienRewNg0J115hE1dt447Rvd+VKJXc8xebHdACIIfc
/2gWbbVXO5s9gSfc3bdLNtG5ZgSJSif3Vcftc+O2vl46piBSkE6003H7mW8IHcN8gj1qJ8pmElt2
S0pPl7OTA7BeS3lhNENg82xXXW0KS+1NHNr9m564J8iTBxVZETlmw5SILNAGgdPJ4s4GTaJqh5EH
+B1dLU1WkQWUlYv4V4PsS/Rw1W1ly4/iv+jwDSRoS1AchF8m7OyKjvOupYbjMQPlrhdkQAkl9et3
b8RLd9LsMZ+unNwWyYtgbg/6THhndfLl1qipK8vWiqH3U874zIcqSkvJiVjtTInJi1b5xzyYSm8+
QJjPv3c1S6v8y9yVIwzpajiMwkG1CQUi8OsWW/dbhqI5WWctZWwDGDWjuzNVKKsy68UJWmHnOVDz
qJ2EbShXlap6hyDMvySORgppaERL089kEeKrWkOEGP2do396gGFrMOR/a/iwpb0Nx6AiOa/tGUMt
pSB1o5a5oBXrLI0+w+REsHdjhpTarkdPcu81Zm5thPVkTZLbUbU/ebHTNQeWpV+0Msh6CZvIbMAX
g1DVLcYWHQcj96aiIFkoSKwP7WjqFsrva4LYnFxdg4jIiqPl/u4sI35Hs2psR2Bv/KaF6oDmq27K
pyAC7AjOo6GdMMlGEAIcUXaO5CMBFnxVCcCBxVwfrKVrCUH5lp2kncSFYjkB7fb97HHOQSZXJ7+L
AMUfMgDsflrYJ39EFj3U/+xxf07fceE/EfXaSaRRo4tWTv+rs6SznzCx1zg71oB5fZNKMCHgOovo
kTSfip7UqIqd3wfz9pEpJB85CfBmwsn7Hw0023QfIafz5vyNR4ORGQakDlVJv6yNie7uHVHEZ3HL
URCtIbt/EM/BTZKkcF9yidOQNRf8ykTFdosyQrWPqu15jLeozRAtvAHk0k7j10Qm7iemBkrZnho7
KbMmHWEHRE7Tlccg7TxFNAfReAV2yXdg21cTd7pdhrZgr/wCpIGx9o3yJovyDjpV2AEAFLb3a2Ts
a0VMcvR6N/+UCYw+CYLnI3r7dFy4nAz5pxbkl0YJoQfPUs45P6Nw0J7CwpakYI9PvvvZPpqujRhZ
jgX4VDOo3cT4CEMj6ZQGT7DgMIKns9KzLiENiMQoNUibTFdoE8E+tHIrBMCFcDVF/XnqgwozHmMP
XooIs4DivSKDKGmpwMOiwoE4s8Q52ajctjyPj+EMEnqZanoEmptqoy+vSZ3XI5CmKjNlhj0B0nqz
Kfig83JCFwgpeDJKAL1APk6jry+Wj16RAwHc34Yl2sTE8wCPlpgwQtBe1IzS3rWcqDg2/diIEDkt
twU582zVSuMQQKGbDWP0/MpYmdb5/QyX/aS8WMqPyXpKw5uvJSWCTyvl499lwJrWGzvx8VLKupHR
pRdWHRQkE1V3eNkHtS+3LxYQO3ftYzdLQsuuv6cjyOzSB+w/RlmrtdU1wyGtlKkQaKi27JmXuYFQ
5GZfkzhxcPWMc7qPPveKRKhcHtKhqx2dC1k5GdokSoZmEQU6KOe8Lt57rwUM9F/p7g8MrwX2mwrH
A2tmHHLDl9QtoWvx4b8CKR5dCWULU2TtXL/BDRvm+f0R9JY69NUaeoQwuHZw3pvQTEEz2McX30Lg
2j1N0/ViY29LICraZDH9cnHPEMGuepymDpo4Jr0bhc4e+oMXB3W0PUCVFt+Q7gN9rmf4ps7+am/C
+Y/nmHOu+skm6gKtOhaTUuzYkRGCbwTr+ir+3h8FeDMRJxoOwcZ/B3+q2OQeGNP4HtVghR9Leyq4
01H/256P8wjO7BIi34Mjb55MLqUZAboOzLU+40VIikGCwGwsMLA+JYrRExCxtu8JdIDVkEKOOlK9
0bUmNpFEH8Xw9f+gUYIaq3vT3AeLtf8620aV7KcnnVJ8Lh6THI/zJrJ2MfD02PtwMu7RGaoUSVSK
MiaIm+oQVtVWW/NSQkydYyA9fkVTKCI5CTyGZqDpfHU5vMfMkuK8FXxf2o60/pKtUlhz4Zibzwfu
WCnmXvh+ErtAVKGRml6YDKiKN1sPKL0kgFuaTueztvJiekBW/cIJtT8a87RJhamnenq4AwzHsQp7
zyO1xCUWiwtoE0vsGtM1lTbs6mltQYX2mP7IIF8LAJvzM2s4gyhu5h5xj7rUK63Y1G3Oxyfwc0Cs
08st9lBqqkHMUgebp9D5euqxyQCV+ShAf6DfUIRt0p94jFEVfki46NFfW87R/Zp3Ubq383dayflX
u5Qi9/gja3mm+UNpNaG21pYWHOdW8AKvmZk9GrI3PG6pwTD0tTJVPn7hVvbMh9NOml9FxSSEyf1l
7C/c0XOeI0oo+mBnMsZvu3W9Xyvr30lZe0Z1XNeVgOrErpPyp+ji8aM69XG9U8TKvscqGLnA/nyW
pUtrp9H82xtszh2RtIJgGidBGcHOepI5iCCIKrLbnecCOrVO4SKZplTGCyMIG22dxc/mCYt3uVQT
xaz7ZRMBPjf74p8cFcRzdZLXcI8TH8BRkT/8Sm8hZdMcvkAcSZWK8ZBHojDe3FYWQXWkN3/Q8WHt
HMwRvz46D8tdPeJiJKbIEiykmiQaK+6/8ToHUt65Wik8E3O6OMuVBYT5GSh7be/lj6s9iShJuXSF
bYrgYOfWXoRqHFQWKthOfLDIoH65gJNqdZuy3ZCGwNgFYxg8KbMBElMiYLvaz/91NiULndANQBqy
UhwsT4ieMGhEnUpLDoi1tFGPbwhDtUCMajFhtgv52uaBn7rCpGuXmgjVg+NyrZQnV6nTxj/cfIJq
rJnkFpIq1p6jmclHiy9YxU0DQuK7zWPXirmYGy1T3wAUL9h5dXUyHklkvqqKFkt2Av7W6GndAjMr
k7uPSYHSCbuurXxfSsAbBCjxPLpwUBxf1tPmkwKPduIAkaM+nuDPVgDJb8XAgWxjdgD/OIOOV03L
TtHn/mVU8IiOyc3KRbg9KYXLXEMwopsJoxDfOkwvzkCwIi/IEsyxq7lH6TDJR/PiGJiOA3uNHJ8r
AhfzcFTpeTgx1c6SJ7K72CdoOmiPhhyxTVqVrBW5M8r/W+52lXBzniM/neDYnEb1dqVA2qqD9qwE
F6wM0kwJOEbuHpy71baQZ2b9CVulS9rqc38lLMXSRj555cp65Y5vI4itbIJgWoo0qGHca+BcSbiX
DjsbF4xcMeIZpsP8iBV4a4CY1hHnYTnRxqGSFpXjHV17FToo1qMLUzJoOVh7mB5tckGn6wIF1Eja
4u2qDVAYTvcYEJa7tRK3sM1qZt389YEtDMltene8mdUJr+z9BAItVtRljGaKARHTf2yqjhXChwRo
ZWnmTyZ3lEmCR4HNjhA8glHs88Whj/n3Itlvt4qpZxLgYWJhMYVSWMrqoRwZy7IUnp0YLWzs+bBY
twqESZr8x2Uu/U9TdQKbglUGbP1cEg0aGMUnARspsZCAR0yLSHL+dkH7V3nHXot81Z9seyedyXR0
aJwLEKavrwAgmowp5gxFD+4gstvHdWsOD3o61TX7uaJXIh2SQxCoHrxXAKoPXL37ROM9L0Gbx6LU
TDomCVA5qfkIhVlpTC0Z7Y1GOol/26wfQ8TgGLW0a8auLn4uWtzmuzEOwf7Ohq+IqEoqxX++T8Jf
1QQFcQ395jJOSvIn/fNpJjV69zyCgY0p4gUZDysrX/qbiAwB3VzZE/37ZFLyy6xEglIQbADPIxJv
CSdrWBhZikSsDn4133UQoFlX8T73chfTgR68rexqPjXPeyg/JhmGjPZW9xZ2ZN236EHQklHVgbw+
q2bY4dXUOZzD4vzt6VH5I4xl1YWxTPM9x3LqTQTkQMYW6PZFnp/KCaFqQImFuilSHnIr7lA+sLu8
yhsptpO+ohjZQtUEao5n+gBpP2XFEyCOeDwB74Dl6G4BvRNcAHuJNuJzTCjrsGYrhU0sV6gHJzwl
0L6BFx5q1MD8xQCYpRy5WGct+GQEo6NRdeNpC2apqVBuqp/uOshYI8Vlj3rFJM9ftC7GvMPbImy1
WHp5qTP9dygaaHPVi+EU7QgYh3JQAq6HZJMZn8aAN4Se3U07oBbltexmGKDVHeqtVGbAvW1ZR8Xn
5UOqbkMFvdzJKqfUBobf9OCWLl5ED1wgbPNaSgFTiOkOOnfwwP1R9afDlzMAJ7LJa1uW1FOBx80G
jWsLiXwIKoqvpoWa4lW6Q0ImSSKUjDJKHpB4rVhtFDJ9E/LhNyNAxkJvZuQnGV8zbDCKWpWfe/ty
dnKNK9ys+kT0mwAF9Vr5gaM8Zja/GPmun3aJ278n0snUaDn99mR/ziu/ytsB1PLHrMU3+7GbZqe9
HHeVzlTG3aXcCUEAtAoTWUr83Q1KV3k2nZT8SArldc2E0g5zmEG7CZ7p32f5uH7NUOxcTJce33t9
5TPn2NhPJkEnoyff4LS7c5jnN16G6pqqIdqUdqHQi9XnbKiiS74LN5o2PVwCCoC3xzW/WFNYqcVq
cpJlP02UJk/72vF1609yBAWQj12RiEQdWJ9zNGZoK3JUC9kAL+O7yoGgWNOxkgWc8Z/WXY4dvfRj
jGkbn/Ews8oig/q9AJqp9wew73lyKL4zk+NiIMMDpsZ/S+fo+snxhG/vDDdrZ/r8pLX37iXGHKpG
0+tS2+T26oShaC+uM1Qaf6myP3+GKb1wrpvxK7MLJH2B2xtNzCd1/3cqTpGBLt1LK1xkClBjBX2Z
I5wjanl++QXkV4SVqhQ5hpG4cmywbmXpSAFc//ymlPfvFWYBrOipT4wCNJ3i3xkl25gJ7H9AX3kM
eMUm1ZP8EAELq9cAGnFKhIKcThIDtKTNLvveNnM5gDESl/+CPgH8yFP5b9y/I5fseZ38FR9+QAgP
1BKjFsIdYklDKtxqHiQQGj0SEvOXs6h542fYMV3oluMSsNR/paii228RFi7Xlv5jz79n8A8EPVOu
N0Wjs2cj4xBwtPZo3mA1LY2RXQvZzoLcGiXwqgM3k/gd/y/EMahttbn26L9l3/qy8CHkjB9UJsmp
eaQLEmhcmgQpb6toD5faRA/+W2NR+PWq7TmpJGw3mgsUHqN3NYHqzn2hvbKgITgGnjkgJrA7cHtQ
DXYjnsnW4TMb1ZDyIYySeGxtpkPVe9py8E2MIrve/qwhSmKBYoWDLXsrF1DYSWRs9u99qsR7PTJK
N42VFJMHEuxU33wfEtPpXUPTnoHGx1Ftdcs5rTIpME2rwBTyCPcq+mL81cMiCLZOpV0AIqROf3yc
4ANFKU3LXwJ3JjJUuFmE5M7HlXlwhlzG3KjI9ysUEHDEq4xz3ZDDVlTagj6yIelr3Zmqplkk67h+
AwWqrw3AqPOsnHfJovZ6fcCgw2KE2iu5Me+WVkBBQ1hMDALBAkR/zXApo+r9cjoRukNmJKekGpCv
L/g7PdZHVFsOhsoHEhEfZeUGiuObkdCsnrRKFoTFiuCD7B/S5Qj0Oki+mR6JLJ7cmmoR4IGnJE1P
DOmFC80KRUlGQoU7MY+3RE0qzHI7D/yYJTmb010RAVfBg4T5X+cEKUrVsOn55jRqegIi85ublNEr
GnscRVjJdyapQs31AY5rDVDUGiCX6P9UPHyqkvFJh4kWDnofnzexmjj62Y2m1zq1opzxyWHLRTiz
+bZO/1LUs/LFVeOnHaKGStnlPu5PzLyfFLSJbTd1JjJAH4wF65VCrSRTgK3hpugfavHZOCIZwHPI
0dpWqwzJjFDqUSJHgXETtnBUnVjxRLuTD4AU1cHm9oZHXKiFF+jQXLMNYt8xxdK3TJVALzssn3kv
5kXJvTGmMPNWVZF4dJj+XTjlS61GAtrBxXjP9XydcNTzAbJqgVMFaqGPw9+YpSZ7SWxPK4kvm4uO
94/dP6kNUrbKy1dN9ntPWAyixumSCbt9YcTXocdn10KoRAh5jk4aoYn/ZJ49D4BhlIUh0aSYd31N
/UpOHtbS+QTXYGbtdBluLQFC+Tkhb8TqcdGihPZbQEFnl77+5Da0LmYwc3mjBqw01xZYM+IYtO+I
OTRSwPyK7VvDzSp14xgYb5am1MJxn/BHANb3CgEf1rD13N5grsUa+bQkXOlKrE3SYDnb9vZgijpY
akhwmUwNgkZd2HO5L1YVP06VMVeITO0AakgM6JCdQtbnubT4ohAt+cDUea/nQI83L1s0BuyOGt2c
Cj4FM/VDz9Zey/Oigk2aEnhvxM45l9yz8KGo42EhzfrChZ+CErhV7m11XNWCiKndkAwUJ5P2e8ZU
DkIQ8vZ99V5MbS38JShj6Weo6WnQbruOypWDISkWI8VarspmY52ASnnonYr3vIoRXCsimTL9wLBr
HU5TXfsfR88y8UOZjJMGx6TfPNNB8c5ggv3LSEnfnwbKycZPTxY6bB3r/qHTwPQ+5srrcpxl5piJ
QUcMWkbekawmHLGiqqzWe3ypwb/ER8YGomb15ZRZXzG/YDIiC1x23D66GKX9Mx//0NF2ZWmi75jL
KQZxcEr9jRPHYqtMhj9G/E3+yHn70mxxF/ZHvT4oAtIOB/1JZ7d9a/m/PT/kn5vQ6yP75Zt36bNu
KZEBhV+u32miWDuactg++NGq8J4+Jq1j6xEZVRUOXpK0Tc3SEg4rKbBpBnkv4dq6pnvosMV2Wu8F
CWfVagrfSB2vLsykmO2cNCKaY5jIBnG9mmDfje83w/90Vf1FChj8t4RcQHGRn91ZgDt7jsmDVYHq
Nx4j9TG6Y3V/U3GMW4X3DVCI3UhiBJjkYjQq3Db9bAzkaUKJOD0Y1LI8HZt0PMxp8QZBlVPo60V9
Wk+4ptReYl+gtYI86KT51kKV8bTQoPhPYLcUfnGAU8MbGjf2TOK6B3QhfYSeDbQRCevrAS0Bofn9
TA3Y/04bicrYTk9n7PcoITPwfr7R9Y378tXLimUUT8GdCIzCqojH5f+AaEYsOH5/8SigVXKrRdjV
Q7eDovMwLCYRR+YEb1AYQrvHBNu30Nl7UoSL0O0d17gu7YvvrZSW/jCr2xCfEkWFU/2MwDM4seUL
TQQ0FHrJCWvMpLDqrzazp7ZsZVE0lyJiE3yfNOH/1FJYf1gJN9daG/kke1u01kwHQdA6NsmWjHn6
j/Ek4Fd+ETDDLkcLm64od+B2NidlQSlXqJLoASQJ3xz9ti1k9zRnYgIGfp7qWgV1b4rmbADwO7lX
m/v83SuA/cbfYqTkG9jBR5iJA3kvyLH6OL9veHHU2S7kP3rKUd+sJowje++5BXXOCwEi/3GtCbiX
yUMJo758jWoSDpEqnZiu2kRGk1YmE/eUVj0rrpJedxIdfPuTj7qecns89yXJVIOMUIN5T7MUuNFk
EPyC/kW6PztmCLHij1FTD9dG7LB9R/+AYUmXHTIjmMzLcqEDueEdZYHC/NPR2CXtUC/f89qeBDXW
tendYnTdRz6IzGkAKYxer+RedTdcOBVMfkSb16rt//6b53ZHyi5WB1vQ6WUOMzCEbTD2T9dIOQvh
Rsh2FOK7mCpEIPphAJVPx0sADUJuoi6/FSXuZ1v46DPRXpDC1sVmVxxYPZKmWPqNuicqJWAUVtBB
3EHB7W4Jj+wYFPVyhS7OUl07oAZ+a9rE6w6pOdLr//AVRAbHWVQaxD787HX+ECM7JSOOw5GrvBuH
MJVZ8annB+4jebhJYYCEknDPQ5UgF0snGaFPQCll0QATJL+icvb4ELJi0MHePm2Y0p5xJWm5l51W
JbqucoIXCr1SBODYGCLBKS5k5/rXAjONIbS1cj6YVY5/79k5JWT2AKeS5W870vNqU2qi10rL/iuU
AJk+2jQ2Y+NezpmU3WYi6ZzICZbzMxIoXmXUrDfGwuK70gs3DAdyuoxZuqe7Tfxlz0ohqBiMRyD9
9cGuoKZmuBL0Z+8PFg7gtFJ5qsFZkzLH7hNY1Rl+aephzVhMSmvcaWcFzwWZ9MKd2DWVBeejBBJI
Bha29nFfsJIp/Jz7PeodOOb3enshsJhsSj+IElUJuCeKFCc1CpNNE5SnjhEjTCHdTnGgkPi5tZhw
A+w8Tr/vem6r+9SwiJr2N63Zx908osA5nSHTPTLGFArQAZ2D1o6Ey99t1xJLZDBdRcSO7umLQCY6
VS7AlQZ8GnLBFNH8Iz/GK8n9JNsTYJgn5BmtjYHmmYVM+RuAURdFsrb5oPU+zelHy2UQVCQG5qyy
gD0b1KiI4EcblNYTHT/GyoXPCvBf3aw0pNn9/9zpm23pr1FqDGNMsCNjNJxmyzGrrvXDoOEzu3dt
YOK5RDJp1WfzRQMWj7TkIzEI6uQh4ybO+9oSPCJBm2e72U5o0+JK0/0B42CwdkcPrvrLXO9jUou1
IhZfQk+T0EJOynvN/iHE9rwLy9HXj6acdTd1ROLjkPMktfuJSbHGkB/6N0/Q0rsrXbgHmcccyMnj
GAP72DQEqO+yGqso3enqdRBy53HcoQuHXjdtEMcbZx4hXInnIGfKwdqTip/vbxWtgCfDqLq48Ee1
YMS0IexmEPr4VPctW40YhzyQFKXE7PtrpjA3RanEipbThI/glAWzt9Wsi0n1r+iuFrs85BfBTFcC
KBEoaqg3Fq9WK8V4SEdfO4Bo6GEIMczhcJQYI1e1mXMvN0t0nBGOpo6kEF8aHhretUJ2jxg7qAMH
aViPJoR7SVhncnnavaLp6T5rQ7blwoAZfSHDABdYPE2nQYq22Gtdphr031A7M7FSK3s+jF5RhqOM
2VB251M+glCKtUgglR96NiFPlv4D09ZrCannYPLgPoUCjpgAV0nhhL5+dKcqZ3IgPG3L33t3T34C
AWsWV7dYtW70rednYHPUILAdwmsnXhlcMLnEI3L5cpmhm8g4AGToh73wzWoOIt67bre3OpXnCx7J
jOXGlItTWBDMHuExsX/vcusDiWdJe76hcPENOpQH7pI4vqWVv+mt/BoShBhiHeo0pl7zEzQIE2sX
sofKtU1EgxyzMb9XZf3VonK8nvmCcdW44gB/7USonxpkVMjnoeFNSVR/z33S9q4gM6cfnZFPJsiN
oSgqjZ3i6H1WFMbiFic0P0eO+KbZG47gX7PbGGirtqmByN5E7D9onMLIqOO2h/uGz2ttaaqm+0WI
grbZpnJyBzIQcnHjs/LTQsPNwJeexQkxM+bTNb4JEKYi9hx3RD5ZaoQNDeyXKBGDyIdORJQRwY+X
xv+XV2Oa1j8CfzaSffT36b5sssHAac6cTTVDgk0sFhHxXaEV3juVWmjf1IKj+Bxqz70pwAtLYR2i
/ob+h+vAwoh1FabK65Q2IUXxETQMTzwxoTf4I9EROpE8hrsvUgOTJtVzH724UHzkl2hTMlwe9deS
Sn/YTAAS4Bwg24yVVX3PvShGzYOeaiRZrcEa1F58L8lp0mJQ9hst4ac63S7mDxe+w8Thdd9LI7xI
oDGIhEtF+Vr41qrpJOCwR1hwCauv/hd1GYWfQ6tI1IAseu02LwnKizNjXnJZrPrQojnU1atPqTs3
34gwIDHJlKVEUpj1RTTXP9KIwQzCneSDzbGSAnNtbnnyxaVoU75xBwSUDm8kCkqSMRHv+uJDNF1P
/vg5MKKcIfUaq7vsDQH+4KNw6R7IFY5KCVmPmBoD7S3aA79vjlS3ZzWhsV0TI/LtQaJR+WxQ1biI
NX/EOJyynnoQc7f5bNjlASSbUGc8E1kEsuymlBflS37WyL7uRVrEG6uqS/DrZSb71O5W3ot/bu/A
zVhdAnsJvZMQ0cfAJvIzMwNFPoLmesmihlRP3BtqFNrUeGsw4RZjAMASQKE8GtPdQANFyA8btT1d
W1jiAfa18jhBYZR4g/Y/x8gs2bC4Y94Zmliw7ENnGNvzVG/YKfp6mK8XZ/Cvd0lPp0kWKo5zLLrr
bLIf7XvptEFDgqa4VWxOtub+JgBTdBHZ3LDA5xdHxW21S3VnGCNRgaGivZw57ceaDNedlPwhpgxd
YdK1ZE7rj+ibaUq8uNY2KVoqd9c+2mYHi7mYPc/O1Xns1ieNihQk4sFL0YG3oOzdfKVfeWKHfwRM
KEZe7Y6bI8eXGBzh1YugYG4IFwOloY1lADg3M42uMb+dY/97hA6APHfEKHnQZ0ZwXixp8/It4ajy
y+HWSQ9ySCyso+cLMn6LlhA/y95MQiuZ0z0gVO+lgKRLznTZUlGqhRI2xg0OZcHnGd3RJ5dca60u
auhxk110bxvCIu3xG0KlXO7npSeTfwFnq0o/XeR6dTMXN32JA2RSRN97VQBZWkVGLiKIODuvW/vL
aZpgRsXIbzXhWPySimaFf6El/+n+20cEFEABwO1FVQe/0quUXdgsk6Zo3ffqG/7Ymt74WMvESOJt
8743hYN8mGVnaotmE84hXHdhIR0NYjq+aqI0ICpf8ruSejX3xN0uds1eMq7hGgNrrbbNld+HkUMU
sDtmdapQzvTHf+dX2p6X1esWrfrMfftqqa4w1ZYcYd15q4lQhODXdhfDgx+V4LEz3FPm8p5ibnbA
+snq+pSIDKFDVvvhnfNR4hcSu2P2coOCQFndYcaIp4nxIDxlj0uLni/DgUa6UIPObmwFYgbLoupD
rrOWNna7vku9I7ZZZCR2Hg1GzG5cEPQguIyqqSRVWMAXM3HMqkZQH6vvtGnzgQAk0lU4E+fmwUt+
sCrzMr7eyesho97gyMo+18crlrJ4HJi3xHbiNTniyLNGQm3ciMozyd6jRxjdA1lSQP854in5ZHNy
+pGIjZbx9hGWlbiln0eEeqJJ87NnK+jvHxDXIOuMBlQy8Plufn92VD1k0w8ZnPjYFXJf4n+ulw1G
kfB/0BDHDzSNk/bwnQoTswiUhitL80sFPCfCq97eIeNK0uAfUVW0PxiIzaaZ7Whn0ZHe8GX///DH
K1n7uU0wnNs27BpxAI4YOFUbnsyQxrvkGJp5KLBvpqaHUcnwYLqJPkNNu3A2gN5Go710Jui6QmmH
EtD5JcDWHKFk18VAwTdsBU64V4+nOQN+atGtXXTIsHRtGPPhsw6JzrohUAdzR4xWn46JHbS06g9X
toRIfaNRMEZ5gu+2ms2fI45K9d9e+q6lFftXSAc8miGRyBGAqefzGxVDU65lZ15RgqiTeWW+kN3W
JFYmV0QZ9ePsmdk5htc/pHw5SDnS6Dd7CoOI6z1yi9WAXTKkIG9KGefw1ITP8abms0Ag7PeusM2j
sJ3prF8tNh6OBFoEVjI6C/s5NCf8dcEkgxUIp+2+T7Ein89agLuD6s4+1vZuoxJu6tx2YFjQWoTH
qRm6m/DeYYfG5DGXr1E5Dl86P8nncqBY6N3eXfp8WU+gVwZdDIz0QRUCBUDzC8vucc7//ibYrioP
+VV+PMA2l/GoqqlgVJGCqtCtGoYCsG8C8WRLim86CawBWVuNouPvO5kA7mTRNZXZdmzEfKecISMt
eYJ4ScJAZ3MpoIOgbLUoSotUg/coiL8xDo3D8vFIoEARHE+/1PBWz6Zko+P1fZeHndQrum8TiyUz
QDSGhG/UnVbrhrLootx3xXG/5UfOxxkCh0AMv0mWkZ0xgNNuKDSeOPHgdSodMoi9EqjBR5dkfJt0
pbFlP9+jbA1OqhwNN6k94l9g8MkKEWltRSxl/ChkOBX8tDTkXkSXQeaj9TD3uI6MsPeHLyqhNjga
DxQKDv6twiPz9Fw4SjLFNs9d75gp/IMh+yRPR7DWKJ6vmPjXFzpUq/4NbcG4Ac8J6fogFkm/ZLcm
EGQjt/txTHocdfPI8IHnwRfmIFevDyLZtFpRDY0XjPPNrUUiJJPTn0cdt0mU1AtU7gyguoJ/veo2
8ZuO/jUaIS6LWjpq/NlCrz5KuEmp9WPpcoWryQ9UhJ5Z/fBeO/GlzqfX+w6Jb/WasBLx4pU18bq5
e7qHB+XDfU+QHWVt5zoALEnNiQf0PzX/N6lADoa6DgA+Cip41AqeQjeAd5G9EahI6gtu2tG4+p6d
o/aEhkihsE86qvoc2UxL3HmWGzdDCmS6+fLluubX4EohxTas+BzWtYAHaSxEoUvFLg7AflA+aF7J
kQ8Py1tPPTo76eZ8l+NpD5Z1ZFy/sAMUypVP43Yi77n6bFkmPQ4SKRb5ht/ixGPsNLt+CbEgH7SW
TNgvempJsX6Aa7MftcPUJZQiwThVrPgEzDfBOM8+syP9akuGloVaqYSpKvYE2Td1ZPlvZkkGFHJu
4guzERTCVK6p0wRCeyRvUYztzX5OZQ64X5yTy8tSFn8gsb2VnHDxZXy9QNIrFCmUgjuQ0RDMtPL4
qHbUa8uTw4QkbU7/YiXBi8NUka14ZAwu/ODMBYYycCMDHfJGOHBAF98dAsS4+/eOPXyZtdBb4JXn
YQkY4uukCKQBN7MqUucTxyerA1ijze/LGGu6BEdcSAu4d1GvjvkZlDv1uuB4xvaO3qAP18H6d9WR
OGK4vyx43fw2LHCmC9DFv/h0szIdDnG1flqweMnK/xcmrlcZ9wRzMN/ZTWwF5LEbNoo+5s+Od2gZ
CLKyi/OKFE8iCEoXaLYU4bAzloLWeYjYq3wRshmQQYWZNuGB29b8xMm4S5kZ/zkeoKlIwaGOrcej
aPIXAX8ydGAEyEAeji2YLtn7VBv4FTnjNMnnLfac22+uhWrOT0OLMWKg7dENc//cSK2MXCiRpbV7
ucJ5nx36GpUOXy3OCgbOPmbhCm+4o5nKZIZCBsd1Yj7TtPo+76I12JhP8RhwnxiYcxlF3y+6W1yF
wTWXJal9F0u0Mii1Qk3TRJQiy18ze4+B3oQKhFTbL1DDWzv9OHXOKivK6L1LUFsD3J5TbTKUoZ0o
/bfv9WlxWnn+HgOGehtljBTlgsC9KbaP6hrgGCeQCM69D2bGSbI8rrFnOU5DbKcHqGtdfLutiPyu
uUgPn+QoksiC+oKJnYE2XPKGpYN4iKTa0B84hgT7mdydgOL9F8K5kf4yzRRN+vc+FqRz0aASdBUE
m5zgBAScDgzQWnUqFF1j71ZiMUu3xRgg+2r/GFLgGWa6WceXqMkFFHNslv9fYSBru7xDpbIdM1le
qUqB1OTjYhmu03oVeHNirKQeTAoLIXzz9Gr/c5CHlJtIOcCGN9jfkMZedJzi5tNX0SXYvBvDR4ER
y9MjdlkK5+K7UA6sVRwFlaVxCd9BFd00kCGS7gZKkG/N+OKs6MfUhCf/hYXsExffEQu5QKTUzMJv
0ddBtCdK13oJrp9US5BXmRfznwDZ4c7CqFVe0czxbMyACAHYEjSXbDYS2J3TujIdgvUxQURa2ZZi
qvkNz+eNPJJVzJ8G5THol0bKcbgnCcfu6nY4eGPx3/k/5YTrTWMH5Z5jcRnJeYedvaMgKbsi2onE
I4vjwDckg/LLTnBADDqkseFoeFdHLudz6YrZMyEBpovqejkZhm5f+fGfYAcGSuhnGKAod5nGWFjs
LMo4Q2ZPD53cnB9RCpWC+sxa8MwQf9oFhc8NXVeDpr4mIhPtvxsIIoQMkC1hwIqCY+O987gQvWSN
bUzL9G9SkG9A88nlUDWEAAeavucNQZgJWHf/UckFxdMhCiXY/hrM+75KR3TQ2nLdSzCUgLobksgA
gLMRdZXNTreimjbpjHJRqafBd0iFa3N/wG+sFCMhYPoJ11C0BF5MDIeBSuqc2+OYoM1BITLTzMID
6UB1Ckmc6e0m11qEuPo2BhAPkjZ7nBiu4gp4PcxKOiV0LdDAYQ6N7iCi2mb0E98eTsq/o9UccoXh
cChRIo2HOk3e4oCSW1OJDInelZ6ZMR7rfJt/l4vc6M38Ue516dePugz+YjtJq8lnNpYgyippBL3B
pJbg8wqNzlDWDpxAPCGQqM5Gu22UdS/uVed+UtYOIDTI+sSm+4JFQ/9OV3CADMiSiRMeCnfkXIxf
5xUAk4ydPJixYtMB8S6LdIdo9tuTNmq4nmMud0ojw8dUkRog5L+LFSsVJE/fHy2wHSi/N/NvCXDD
tXQYNEGXthMt1yahH/rRh/pKRaKs/VKa8gPm88GJGluny/c3pSs68+Gd5bX95VITq1cgFG5H9W7J
Tze68SUtqIje6v4rS47SY8TbJbsrIJu43NyISGTmfmFCIeLxQPRIvHSlgCN8+GJ5jnmxH4s4RCMX
2aZ5YbIpyTp8JG3+ICY6fsPUh8gU987TZGmIlFS2Od3t7tMGowHbhuTq6DUWoYmhJsGNgvIB6/1H
/70vBKcBSCTT5wqpdU1kFDFUdHuacNhmfA6DD//3viwGRUgrBs04jCkKU1D79/e6REzIWvJl+9Xv
PmvWpb2EUppO+dBGRLRJl8QiQ7mRaqrE5YZjMdub0M5NQnHJVpC5MHi+Sjh9PzIiER/ucMuODTFV
Lx0Mnlc+NB/yfsQK6EySihIGVA7OFk9SRIJRH9HUDG55rnCLNjASCjg/OmFPLFqlSKAlAbgehqvQ
UUMglDmstS3Wluh5ORN80aOZ/Rq9scv3idOclSzs1MGSnrORdb9mTFU3vJg8rfX7FQwNAvkm8BuC
j5HnVQ8k6jFdW/Y8wDYyXxaLCTkTw8UyuIo/o2SLX6kA86avrhu3NVSHN297PG+PFfXxguFLWMII
TlfD3jAPFWlZEV7CFwSPvg4ao9o2aKsWt7ZtBBHhx8qqDZIWKQelxcBS2HdXhlb7wBmvtYaa6mnh
exhaphJza2Pe6I2WOMmSRovLxui9PPWVqf6cfsIEmTMaunJ4YacWRhKj7/xjvtyZEp9fPtt5FDOU
g0uFLrg8G1GxmJSyJZv6fy0/Csn2O6Bhp553MFyz6Htu6K+nnIx0Hbgbk+zP3XLyhcR/eQEM6EqJ
i0DBvlCl0Wa4y7USviu4B+bT63gx39brrti0rrrUq+Ub1XM39WtiBnJc67EPrMH4TVTGWk9UisOC
4shbAONWx3e/RT7+PTUfBPtDdE0oyDlUcHai/EWmF3bTmVd+ZzdDs4LIhkez8p448pWm/IikKTQK
+T5dl/iTzFdR8pWGcmWdw88rf5OKiBF8xI3idRzK3E9SzDbT66x9mTxuAz22EFWcJIlrPfBkRzMe
9xUgdHcpsLCDKsXh7xzGMOw2EWscvyDcc9ZbQsiJ7KvMjCOXDSjCFggiyZspzZERplZNWYemrWXM
mrr27sLDSoq78Fvi3jLIsn+WfYaAonv9USIvwC9hZZPnI5wuO0hSqxRXLNVTnHBD/PwFLjHuVJEm
oIQYs1cX8UkgtXrJyuvgOaa/VqT8YTev0an3UIWdbnFZ5rj73tk7pOuR5x8YZvtnbvDGydy4Hl34
Rz6qDj/X5bYEHkXkgm6Lvk9IJ3w98OTcuKHpnnZd8aKxTX8+IWQcHcE2uTrgyxN+Jbak2+fOvhnN
+vOE4/h8yzY6tQCwCBrsxufVk3GSbZSSYMx0MpW9hZj7qYimCudlSNyXpszLyH718DOvJ7TbLHmz
BN2gsdRVbYF5MOv11HabRjvxDZ+sUyKGEEuzHhrjFzy6GyfXnH2l9u0BgVGcmwWjEwOu+SedPHcm
Gw/ZmxCFQUIrZzsLljR/Qp4Tbu+xaNuD/Nkppz2mC+1fGYU12PmBmMsG2mQSx2EUJ+MKUHsG0xPs
VIxpQ+uHIMHlFo3x+6FaZILrzv8WSGCo/4U+phnEjDFXx43d6ItpY6U89Jl2laB5uDlhRryIOtcR
Ie4lSg7XTDYT83yu6hUhCJopwMdS2OVGO4gMD6tJ3/yJSASyI6IVXhMUHYRX3RHMJF6MAYFLvo3I
lgWWzlE1FCn3KEqMdKCHxeiQ/Y92s6GBJFUiu/DEnKxDTHebAEdouA6T7P1MwBx9i6NLPXhqNEmD
V1FnjQ0qFe/KF/sZ7h9bEmyStyG8ey1vE05sMwMZQqPXWhde4iiy5h/7F9VKwZdZSEX7V4IobgUJ
86gsb1OSNHrPVLCnj4xKNLp69B2KSkjyjS1NJUJdR5bBQsz20TP1LS58qsi9/qMSS+9lxmFgPkDI
p0vkgb3o0pjreV1C8VTN82ifhInDO/rmm4mGsTNsuBafvs03Z1Py7RqSybP6V871A7TPFftGdW4A
geBhlp8gZBlZKST40oYhunURPU6iDOgUrEYmrQ4baB01RFb84HpRoEwNiQlWIYHIMX3I3Ge7B44g
Pjrzy2BCLHZoY9otQVbfuUW2KGJQ+LzaoVlryTBmzIjT2+3jZt5sfNxifPZ8p7YvmRl0+Nrv4YqN
5V8m+mYwUWMWxBmOSv74YvNcMAAidc9MrkGfm/FdXMbvesojPTCgsPG3xAKIcJECkllvkLI3SJce
QL2rqXaJhsO3RqhyoUp2ZFiClm5smjheYncoPjbsUyQnlW+H4THKaPzZchFr2BI7cyxkQsViURPB
Bx3CfZ8Z1lHRZuiMp8WP8Ijs/Nv9OcqdzpEbEb6iv6U+9gz7SXqt5F03C+kR3xQ41wDa9AAm+Y/p
w+DfrumVfVTMHpe2gu7c/X6KA910NOoqqYU91xrIbYs8qMgC760MxVtfk+4YY+RMBxpXRhqIeO5p
3MJDhUuB5kPPXXStMIpFeId5NDtvjJQN9qc98wbkdc01nlAN3mm8hsJsKTWGL8TPB7VGyIOzJuxP
AyqmJiEXrfcNfwzborPLwKw1kzdvfGX71UQ8dFqZHMLeAiQTi7uXVjBQ4oKB2nsd/RDZ5xwq2Ch6
bhvuqKjgRONFaAkY1T0/ITfVWsc9LeGc/kj7tJ8TLGd9O5HGZj7RNjhzfrDJ7vxY0jTVpmovjP3F
eSxJEaVtOR7DdDtgan+uJzUJn2dwH1rYN6T/K9qXvFp2F6G6bTJjIAhGFzL/Im0q7q/qk5fcb7XS
vZCGyt41mSabxOBMw33HSyG1Bs8L9G/RRtgnm9ZVATg0DqHb4bfNvmxaXYcxUcxudcOPIPBGKCOD
ULGCYw8eVaSj10fe3YHqmDhLTLG9IdpaDlGb6siEeVYx10xDnFh13Kokwzmiz3MjkCLvQ4agyLH4
gw4TRwfT/j72QVE+jawhhrmR9GV6m96vhDODz7D6v0S4sJLQBQXyQ7ntmPSLtlfL0edTMKXks3jN
xfS19CpA8hfO5T8xpasCaY763Hir0S4ci5mzOTRT6Im9I0jDrUWLwIbCij9ExFo72DBQfXJVwEh4
w+5qiugiBKgnCWoZE5T7RBNSu3LXKV/XztAUwWDOdBoEEMDhrmnQwv9stMoM+Du0lDspxZrxqNZR
2USX+aLizZWWcR20JY5wfTUv5HpvAtHH5AGYn4BNKoK3Ry8W0wVH71YQ269VSyFbF6HsE2smsMvb
mNmDUc0CFQ9gBoLx2FTtz+iZK6VCy/9UFvKErHDcrmBttoZv+plHDiv62cvVm4gLpO6880HOhfUE
G4EEckl48IrtasVnV0XKQna4TfueFAs1FcR3bf7hIrT3dLm+CEsxy+1PtQsps4FwCtor4O7r13r2
EGp77HgZTevpPk2HZzQYiyoT/TSqFnvyJm2txJMeVKz5unQQGWgfGnZMwJAJxDCv6vpq15RCeHfC
eT9nOpkC2TjH3rnKtP92jjYODcK7cVBUInpqQ446YOlJZpbh7tuyGXNvZcI7AWVoFaWOMptAFCqs
gH5zDKLE5xTVtGAP645f0S6HVcczAt97alS5hsRamu2zUzHPSeDktk4Ix7TRF1AEpXrHDYjlep6I
DSy4C503fm0sgumwYXSsEikngV8AaLiCoGFFnWjvBqHD65fkZbDQVZC/bPvDD/FTu52g4DBJwdTf
soZGlBhNAYGs0WrLYp1ARzdcdU5/8n6KeQ/3IGid2Y6qfA84wkcXZyg2XU564mNsmyW+Gl6ERaqM
g3qKKWT4Sppe+ol621zNiLVkDXyPoaHaLK1Z5D8UGdyjD7OUgVilJh71fY0r6IFenOMgjgFKoQKz
BL6PtoX2szhUv9jZHFWS/j/2bA8Fk9hvXOxc9p1wGU77hLl3NG+5gCLOmEpH1ThPZEUMJRyOmsed
GhLKJ3/thPNhtN4L+cORtf9Pq9iGQoMa4DXB/AWwvBk/nvWGVCF8xSb7Ib2GfRAPW1A/7+5EFzcS
O8SYxnn7t1bbRGrB6zbiixcu7Awm+o0nrWPaT+OVePtaHIeroCyyid4SuNnVdCosHuk8Yp3KXJad
vxfmEqlFaA4YXLACa3O7eY9Dj7xPzyy7bU/u3JWJyDtlF3t+CjGd5hhQEqb2WfPvMMtJQXhWm67b
n528Qkhk/B/xyAv0p5gdzNdHLzqP52WtY684WEQx+AYf7udcFb0hnkqaPvjcwB+6IOIbIwWeckjY
TARDweR+heOHl17uYlEymB29oKB+QBdIkzBn5rpDy6G58YHnI0ZZzEz5ujfbIGn9SjAlccF1w1VE
Y4ZQTWAKFG6dXQTIBp+hc6JbiuF9qnbZpHjTswuqZxOoTQM3JZ/QoYE9UCkvwFyUJvBNVu8jU7QF
g6AvCTNj9R22Jl9WV6FrLShBG4P7REbvIKUJ6DSzYgeVNopwgtEdOwKbZOi2ePGUM95/iM/QWxLO
dKO7duWRExESlzfHDnxGuzGAYSTLQg+C0xNgkYFkgvM/ZNLXz2iheDs3RV9lmW/Ta8gNrMLrgHUf
BRu8h0q4tR7JQjliJ5xR3n+y1RTIFZ9chcxSMzfD5ZYtQfjxk6pizTzR7U3zvEvhyzpLPOxmV6El
8dcFDu1rrayGJb6Ff3DhGLkffKD/ivo6yvTwJ7g5gH/HUiMEXVB+jQgEKCg1U9F1y4fILQOxaDsQ
47v3KZE3g/PXKAXkn7bKH0VGCFC8D74zVs1uxd9RDP+n/7D8HcBpHSRGA+NK73b+ISVf0cc9l3iU
zkiPZ3sEuid7flj/AUIaum1AHEUrdXl8C81ZMhUFeIJb27RLeEOY9r6HVaIlAmn9Mx5ipBR6y4Fe
JwSKu7CnNwwwS9107dy212DlZ6NnODsaCyBi7RPcUOOlL2X86cEkxV93hBl9zeZYgvxdl6Kqi/Ei
00H5aLzq3SvtW5N/XiUUMEXbxuAcBuXRNl578nF9d3A4rJ79xBBVjyZKgzeZR4h1x7qLyhp4Wb52
EH4dwYgGRUi871RXfbbPU+YIlMNTN3/jCrbmMuZ2jqbs4V8beFnXmXT6jmMK72TA5GWQ52UhrvZG
LZVdI8xCC4FOGYOxI1t/H3BZcXC3+w5XiDAWXTqr08UAX8CY5WtINJTbHuIpg5FdMk4v87YDsXzZ
WsUCAdVmBW5D2zPN9m7Dr+tOva36XkYd3V15mQ+GcMtKEeJGwphZ7ryMBWgTaDA8DKj0yK9C7Oa9
7VjCcAh4OKBoL1qZEmxmqX4/ax3gJaS9qhl449yLX4bCUWl5ZN3o5A/K0xnxq5mzYSPU2B+n4jBz
qLmdU1H5FprkFtUSO8amM/Ah0KPoAENJaI/tFuUIUTTiehQAYB6PeKOlJxtFte32i+kvl++2kljf
a3E9NPCk/KUXEchK7C60AiiN9w2HtUd2MtYWiX+D4V/NJDBssXsoM/e8tLVYtZkR1vzaLjwEFM7O
vs1sPlOPzdOO7TEv7/Es0TDjoQKTMAaxkb5XPp3hRUndROegtyne4GyEgpRZNibSNKo8cwfQVuUU
0KWUx3l4ZI06Z3zyuxTJPJEGCJbDToYbr2eATOqW47oHaj+bIOUY6yOcf3bMSc388h7DoB3u2sOE
pQ0j8yVdGlhrMbSs/8PlZ4Eh3pqwtV9w4cVn7Rc3MVtgvToFxpPljpv5LK3/I7yrQY+7G6oAHBJa
vdTu9t7qw+9OOxnleWWx1pKf4oF6yzXUOqw37m51jJyeQjPvE9bdsXQxl/+tSUnOi1WJIZEg3vsq
TpIRwgZ8OUKDbe+l6V/r2D5NWrCr5TylFgzi4mYY/LnGglkzj+cg87FyK2q3rmhJjMaJ1K7k0Hmz
IJ5bHjNMw+kO/1usrMX7SlYv8NozeseP8hDIZsOo1WSF/ORPJhEuStZC2ufAiaJt+Zc+jBas4qwU
v7bsg2WIK0zVGCGR9gzY+QFPnEGJEwZ2v+3mY+7bHMLpglOHbnm+hTIQ38Q80HEOTjKKL1YPmoY7
oPAUHorEHgxwVd9NpfpEpAJ8YpC9/6gsGWstCJtDAoYnAqK53YhoaLEtTZwFWJPtzLlwZ9fMxUeE
WDr/xvyq20aWMY1sSJ5qBaoak0+i2vjwQCSqVfW1Y/s6RLUZikxn/e4dCnWMVFvXuRU+yYy/hOv1
2gN4N7EbDBOVYdBJnD7VTjsDbc5lNkwx+puA60Q/mJaHxZ9gKfMVf4VN/L+VqWMIbLpcv/bdFMH7
DzMK0ZJ91GJxwxR+VzOjCtrmjSWP983Bo3SLlO62nJARwCWzd+SRXguvBBmwtNyDa+stVlEUvFKs
ZcO0j8p4FxYZaZm6QxYMmt1aZ8Kce/8hc6p/KNLQAAy/mVekUiyaveRH1pAgrwChv/Bj7NT+H11u
lPAzLpprqcbECOutYRlc1em3yeX7NUa05QQgrnihq5LbzuWn8dm6uQ0k+cyVT7uF9jgv8Y5jIFAm
R/NenLwRiImM1bMWZqs2K6nUa3sZxF3SBVjtwGj8i7NeSS+xn2phyqs2vaAGFluUKHY7k3wgBXiB
eK+LqHYAUF7WiVzXRnO7wsnk9Wc9L+V6ZatBdXGwIaRYId+X0XNd4AirLk5t6ya2aGosi29VoweF
SAckU6ovJykJtwsyHNP+OIBGchPlvYOWrnirYtQ5+i35HtfBkZpgn1I1sr+cfu6oAwU7o77t+sPA
GZGJPyrAlOazGR3yW5NWZ+L6rBmGILW00DLZaFMct7mtpMieuOzuMbP0uHgyXD+HyRm8VBeoRFXG
aIJy+nD/s8iNojKB6ERZwq3JFhGDcY4Sg7fqceBm7n03AmxiTp38Yfv81IfzfJWKbJH1sWz+9YNr
T0oZZhf4y+nYSpRsrVH/wkEK0B6WKqXBspUgF5TQ7PfvTART2iwdbFKe9AgtSqMVoom2p88zuvy/
L4wxFM+PwV/hVbhfuJXa1e3mi4ljD3G3qiyAwX2x7YSeY89EdqOmufkbw4GRNSzOyFkhNaMbtgkA
JkPreu+h80iDwhrsdQxcGDM+7Ee0ak7nK/akZHtyPu58tdwbrv6YoVo/xZ6AV3u6O0NyFRi54/UK
tu7yEdAjw2+Yd2ISGus9yklhSFRKk5pDp5Sqgvoc19LUh7nIJNmoPQbRUHMAmQgoXcQDMU3CrnV/
tcWOAs78yA3uK8xU/V9dqDhUeO2DkrnQSqmCE4J8kXAEXd9pvRyozSLLWMqwzGBBEFqX6OhykjH2
yRaxowr98aaaJvoBBURMPCDDaOw70o8seLJHXhkiFe2c5BOCel6yewYKti42M3FqUpyHdpf8Y2H6
1mdJyhEdx/vetC/RBPNzy2VpihVDNhhNLP7fN28BCCrHKL0TM6JQAx6Ol9J5XZWIu8Y6wylRhEUZ
hr4HTtwQ3xgyOmhdIVqhiJ7M2Zrr/eueLZoepMvuZgCWgafG3doitOAY0YJ2BvzIEGYDKP42/hUZ
4OUsAFLw7DF4h8GDbunYvC7HMokMRUpwCCPxdDjdrgjXvb1spVpO4IA3WZu2OYdzITPDRL3cESsv
GiZjDYFgY/ZoanKlztMonM3Mentt6Sz75OSFvKaU/t7xvv69kkRn4pqYLa/+CJSfNcJaxxgk2n9D
e7tllGFJ7MU6STuxPHNiezKOE5kn6oZuZUJYI6dU1mj7LfppJPiK8VKBe/pZy2hsAEbDt/zGjUXx
iQo7qeWe2JJGWmAueAbSFwWoKn5HFekYn9VGoTGjhhX6F8TW20hfjk+amFXb/QnUam5GyhhGKPkS
U7J0Oh2/Q8pGe7xC0GwFgwNrRzoa89eaZGeoenyDkuDD4jryd9eeuV16ByPk041xLLCwZNgWFg3u
wvZbjLeZ6trxeiyzri45Wbwt5Uetirvbw1AmU8Ga3c1krIuhJICj4ZAwJziVZmVOZsAPNbEQuWBC
1Z+87Mj8I31ZMYmRAMLDWPi0EcFbl9chAsmMxmLeh4uZ+DHRNLolk5/r61AmQ5nxnx2bVBhKYvSx
ko5NWlz62dvVAudowHg/axKA/EaJ7xqO0TxRCcTB0lahBYQvUDy4VOu+GyFqOe/KTFHxQuB7RuHC
BwG1A4Mk0M3d78OEobaYHMJhQRatGARc99C9l1iwiOKOLMnsnW3aNHqJ0TVYizqFo9JBf++s+owh
nqqCOln8mVTEeQTG8TFY5srviBI3mymWqCXnwaZ7M4GWY2RWSyjBoHCSwC4HWglNSf/cpqZ/PluO
/dil/uaIGyo3ldwMTQ2FOtrQ9Rn9M8iyVL5heOJA2Jh+WYOE/DaaBFnYK6fVwshKsq6VCPBR1Zpi
B2MEM/Rl5JgSJIQSDvJ/VwXTHnm6fGU+WMlg7yD8mcKJf8GJj3YaPRh8O2T6TBHuk6/tm/eFH6fh
0y7bPTNrqc7JPRvqTRhgoz8U3Sr6U+aKPCU6rxkGDquIiNYgswmC8bsDeX2Y+R+8qefYFZAgMh/P
t63rUhmcFdPyl4I2aHsGMj3ZGoIYqTnOv3ygr9HNHHWqfCVblcFe7qyt6Jzeu1M4U4WZWXWEnBPu
NlNXK8yEeUG7XpN7BpYp1aX2DE4mObiGcR4uM2dpxd2xd67Tt3QAXVVyijHX5ulKOfOBKag30Ij+
lVYrUTXPzKvNrlKwnUCaUIAEfbjFAKrMDFiFQGw2H5ieaLm6jp8ZN0mIfwcaWavGagd6MDIjMXP2
nslp04/KUaqQ73Cjg05xJE8TsEMp93BzZUnwXYTSqiBIIeYGF+yp4rQxpjfPzG0J86UxaPVXvqhe
dC5ErP+ntMiZb88WqR71ZSHV+pA7jRU6j/T/l1t2GcfKLL0Sak58mYJJyX5skDhyj4Vy0FS1KBna
qoTGAeWeHx2RDmAtLA68lRhB0koZH9Kik5H+XYDirYiqe9P4hVGZX4bAgxnfZCh8xWROipunigje
7vas9l+P2ljYZG3Pk6m3MwoOuAyhRTv8x1SojLqoUewaE60RTg9E4O9KEkRag27bTm01D/YISXk+
LDiq2OimWPyxJcIaRH/XTdLr8lnEdOlCm67nJl8VsXmmyEyPcRC7/JBIJH2/p9jnNNCDzQEFDHaN
ACNG679g/5QBj8xc8H2o7LdHqRz99bmm6AG4nyT2T+qD76E/tcupX5wbn98OO8kvel715KQJz6Cx
mcDIbY1RhqhPgMh2hv1J3NNYwNDr71m3OyDeac4T2KCFUmouDGYgP0/mEWmBSEsiIcuFyCiWOvdv
4PwwcZeOcMk3pTFKzG+P8NuVFlbeWJKo794vzUiM3QxBM5LlOB/l883RvcNgw/fsUi7wf6+S/4Dk
DZqP+GQ/1lifIYMjnWJd1Q8n6t0v4sKtYWM3QwcPdZfc04qxnVjUYunGQREztvBo0LKwvvXuVk+4
bmBs7gdbIlIXFaIv4jYq4c7jIy4wUbGQosXA3B04TE/iCshVJ2t+DUC6ViNMb6GGYP+5HmWr0pIw
j5qaBzBurIDRa2eyTMGdbSn+m7dqg21myoGnWAs7/usBxxtv2wJrfJNCP5CwCha/Eu3RACNc5pyt
L/Rd/4DLU1YIbTcif03HbcGR2cSwlKr9q6F8j8dscxuNq4lENS5LTkRfyCt8LSX10UdaMlyZWI/c
U1r48v+nallWGtoxZ2df90lK6SrGnosbQdxeRalvwRW/PLkbJGW44OLtwy5mS7QsUt66brCwOCtt
58mwCl83ao4q7zJyDoM/ZujMLLg2P2yPan2A87GAhkgojOZ+yPXIscJmjhPNRTn5MomWoY+Z8/kK
gASMDlCEFyZNPU6BQWKKih+256/2/UvHqL5t9ZETbl3ZvaZE7e2QwSXj2MX/aUM5litYbgP81nDk
Eq2QUZc+1v38907/cwim+RNg7nxPZGrSOJ629Jxok80ys2mYPv8xV5xIcwFMqDnbQo/YBQ17zRfC
0lERL5vd7/bDWrFveuBgnsKWDIVrgA6dF0kFzmQZSzLINb7oYVUKoNlk9gmX8qTtcd18p0RjpHwe
pONN4rIg5WIuTvxzfuLQruY47AeQWB0AVx/XrqXWF19ygqc8Pd6FQXxrQWJ5RQlkwnfJ7FdWEgop
XJQ5ucQ7fr9Uslk8niPPUzqT158gM/SM1qEULFLQ5NhAkoNLMmlQNDbctQFKg8K5oQ4dMjghj3iH
R7zV0SBOoGxKIvvRqCtqu1eITNzRaFbcuvdnKkPgFJ/qw4d0OwZcgYHdCdGL1vj+/9qUA3FnvtvF
rGjrIDblHLMEH6joU8GyP61GiogPIKhVWt+8akaQQdgbkmvTwNujLZmE3BeASUdarIc9fpt4RXcl
LJu+m9yKGO8Yo231unVzbENK8lj9KMoHFmRK+YZOPgvWi3mQIt41NJyoeEvjDynpsmvHf6H04B98
LBMK7C9qOwv0uS7TKgEhzRY+Mujno1c+K3EuowOYuH9UEbxGeVpO6Oj5IbvPwj5TowOUNrI/kTLV
T1Kibk2X9y0bLa2HO3TYXZ7U4TCR28B05Duhz/DSUR5dcFVXPpKIyIoE8yCsvYgKslSPdTgLZ3Ac
wRPdPnVDICE57b0lHjzQrY3AHl1sMdFpxL6hgHYNqrNelZmuNs5Qe66PBd1L2W5nmFVTQ7WZ76dr
Y9qFBS06U7cQHelLMY9N0MLm6eju8v0C/EpvKwTdKmFtD4teE5JYHdC9X7nsejUBiZrAWg5a68ET
iOv1bHm9h4q9SjgGn8TCG4G16rQTGsbBbqCj96Caur2zhubmP9UXZFbuLt6JHRHJ+KNsAHjKSO+t
rOIvX58V8oo6rAaPRI66/aXoCV5z5zAFwxtHUESVDmd9aQCRMFkekrWRw0JXCv6NqxKURAoyRDoV
VpZuRJto/i429YPd+qq74J9Wfm2SD73RGPTx2QNJaMJxceQ1oPONnQQx6CvXhFEAv10jtnFIDYLU
1rbChL2XRIGw/1eiMhLUtzidedjXwDdj8sj/QkOvrl2WSesYYYTBUiJnBihw8bTyqR+4IhawPQMt
jUWBlTr8GF7AcpDXMCZl5Ncty/7vF2+LbutX50TW5FX8kIZ2GU7sQUFZ75YOPeDB1t7EmS7S2Jpm
r6SN+MgMWKR0a7blplRgdeL9pv2Yeu4N+sYB3vNc/Yf7K9/g39D8Qq9G/fMHuTkKmbD8cu1oP57L
dabX4KVvZYvJx3n4oCvq8Nb3IvL++fZQXJcn0djJMRgTa+DKqSnsWku1/ZwHCOyKbPjisGMduxnn
0WUv/Xu0p9sPgSb7Iqc3klgLjDFXF4UKY5I5PYbegzB+bTuyz0jzM9Mu+IA6YZBJFqg5FlKWDe73
/RcGvI27VoEJzDbgl1PpW68HMufggHzWQmRFmnaeGyzceQu3ZXd0igwQfAC3e8uzWYa6jtCH2JtA
z9QyrlXnl2WakuY79biclHyQPgmnGQF0tjGoF1LJ5jhOY8vVzX5ZOkafPqBa1Qn/5+hTrNoipw8c
gfI4UxESZWRVDsB68kHhLJ7mk0pkotFUzLSSlqdoinS1+bG/7ZF0NqplhbqPveiDW94bfok/o8BJ
2Y22wN2hZIuE6REOh2khM9PznNqtMBtiidHYM8CcgijxHFDVg7Vle4sRruDtRCceV0pcbkWHjW5d
dF0Ds4zoVskbZ7FzsN2HqUU13oJXpdXgVm0jy2r+GHbTMPDfCtgJIWS1TTr+0N5ctmQNqXQBAUbY
6Cuco2DnzXE+RuCLqixBlHDDnPthvBpTosAy2+CD3CCmBHiF0Q+3ODEJfHxjJc8sXpaemZzKNA5V
2gYELtwzup2gO3JMaA7Q0l1+Ro/dVWEOCF6mV/SMHq4EezMDlTR4lF/A4acxAokd3vBdRc5ZBirS
+mEg27DhFbRudExjt37KUWY3j/9OqZD3OgQ6YEIyIISxWLFJ5EnzpSUowKsQv3y2dvRM+7XCoKsB
tyeh8+WWwPujJEUpPKVZzvFMeF9UOEjnyz7YQyAax/5tHe3LgLzNYn9ifIHeNe6cMRnVwxxDgP8l
Ev2CgmkjCUwaQ6zxC8sWtmtWEGRFJufuooAMc3WFFn65ltnjDC/7dekKSPxkNJ8El4ZAefhY+rSH
Dgqfgw5gavMOmH8VgRGEW1FeFE6WnaW/+coj2Qmyfxd07g7C4lJSEaiTADmA/nvvaNQgcG/LeUwQ
hKVzMwjXqKxCI5t0rgpRYpT+hc7ig1xXGqcnckZpldzm9guiEiVjy5aFt1lmZBl5BxtNvO/uINzn
NPls0hiDADt8LsH6zAqN4GwpbMXv9IGyR3IdjE4RLhpHDRd8I9mYvI9CEH+TFAIPfhoE1WLn1EWa
F9Ba3TQvFHGWkw5lhFocCw+jtYzklqpNiASb1rLWQeW2Vql8ixU4+4Y0RSSTJmdpmIIKje5DrozS
/o2cLUWUmYXl0+r7Se/rT8uVPtnPvBLdqbJ5QBsIZktV5zz99qiKl4LGFWK7tUat+NTzKXogek5R
eTskXWRqdGqx2eXLtfkw7QKRJqJCqIHqpeF3/NacQdE+hIRH5juu5jNh7oq0Jbcw8OCRogRV4ZS/
gp/ZpNatFubRoUS5g4Z6vkHBHhlQo5CdGgF5xQa7M8t66gTfLp+EFLQQkh/E+7McjMCF8bpW1ur+
D7jt/HTkW6IBjvA6ueb9gXY3q9JjJFKfTLV44Mz0APanrkrDcx0B85KOC68gT2rQhn1oaGZv96e8
PzlWvBauwr1Pjs6ZXYKwc46UQqyGfhHHiiVYCcyrWFRV8B/MV4WT0Kn0JshWiR/Uxy1tLfY9Qucs
jo35BWFPGAVmqKY1tMM8PQoMJOgR6geC893UdLWpTlxdXDKsj4qAVFjmFZoSOH92S9gJysKXtP3j
SDjHVKapKUmRqhnNrJ/wnPwXnPjs/wLgWey2Ku8r0zYrHp6sYaenGF97JMQQICecURibP6zmkY3e
SE3fW8/PM4EF6OMgsTTQLOU7brQcidCTSk5QaNCGLdCpC539pXMaM03rOldm5pfdCJVdemvuKEUb
KiGrBJRetGYl71j3k2CgWHX6gfA3V0t2DYnQVGA1OCLSQv8wx2UnLvf6ECFuRMsfH+X/R7a0HD0r
WO4i8iiYcgNJrQlvUqtUlxllU0vraWMk9xrVWHYjjwXORm11a/PmY56krXjtQwhlGv+m0QO2fwH6
gqT96LSB6B1NKn6aRJWim/9GBcHD+05pn7j9vtJnvDlYbpAzapP/M9XhJf9cQiX7wEB7EIWVR7BH
bFneumr3TLd3h2XiIXR0+/5sPCF6F1z/7yQmxv1mugLW2KWVCwu6N65CHdEK3i5m5VdTrWjHbIeq
ZC7/o6q6uiLy61uzIX9uvRB6LAfkBhyIsTivQ7qLKKXCRCT+yOwfX4RmCASDuBCKlQ8+Mrd8zb0z
A5YMK9IBKW9auPjtQFIinzbbQXsNEvLfsflcfC04aKNfE5FM3EZD55PdyDCa1+XTQal1B+wefZmQ
HykBx7GJbfwJzn8pelikgj0hMm2pQlrYZTk8bzkaj/QnR74DcC807N7a5aQaTLI5FsDi5L1xerNK
sH9Ahh2GSsfog3f9wD4lxJ+RAW8xCuhboCXrHyyd7hLaBMeMXrDTCkU/I4y5b4RqtPa4HAzBK3ir
ofeys2veCKJzRyOhadS6fyWJcupH9tdPS1uLBJkQbOuQBNrbD50qsvrQu55DXg7m11sqeNBYCkUW
bvxeOpSelVSWn4xid8pjaZgCL9StkkZgSbAf/vzcpoVXEkNlLn7POQUwcsi2lk/U66F4CrnmBYiR
b2P1hfE0rNM86kGK7I6/w84loOun8TKLjVMdh6HhSTsmB1nNDNXkIgwAsYS/czZgivwX7EhGa6I8
V40apaBgeLMf6MyvkjFPybSfjglOuZ/Ofg1woKOLE+3nJ64OX4IWJlqgyCMaBsW0Unsz/2+Ejepx
M5hXqrMnwjT5AxR0OIllVQDZiha7pt5o2xA2WgD8gyIB5RD7bl/UJYsd80/77PPHTDkxVJJlmYIR
6s6q9GBSYVaget0QOORP61Pl3+dJQOJ6xOzOQQuTqlNaXmOr1baWXv7pCSMhZpJj4daK7pho+68o
OXiBUHT9nY4apSNXeec9mtChUqlS3QVv9Guk823n3lEuAIbYryA+KMc6ccjNkWscqGAebg3zM2Jk
u19wtmb3Wfh7iFTCuGo+YrpKaSY6bmSceiEK7nxGdFAGcRj+2dgOCNSy9PKfeGsSlHEa1zExvim6
B/i1WzbQf6Ryc+niZJMUrEeR8OV0hVbCvHOMX7i4OmQnt35kndWfyYWLkPDQFez31TXOoPJeQu1n
JIqB0V00Clt4HnQzyMhrfzX7/IfbKK7OsLaj5AmfVHebA5rXTPkuH1oAyDo85d+dNOicfvhzXMbh
vCJnGDKhdaZ3Bt4WON605nFX8CCzFN2yxRgruv0tfmIXYDsZ7Nvrp5rXPvxPBgTO7pZFMzh5g8c1
nA7M8Qy7yvMhaCDRmAPfD0Z0QnpwYMSHBzpdvCegXza+9zxX6d8tZYVj7uhGrVJCrroLuZqRs4QP
iLeWY0wNxOFcfZGqS4/47pffSOab84j07hkgRLU8H3HzjdMcxRF0c2Uq7kQYUOgiwcVRZ8XsTiUG
6gbno06bSpJCr0jayVIX9QhlGPIAkJWLwRPnSXAQAB3XWBY8Mf1SNAvJTuPtU5MHVPxxRn1iENdl
rNr+88kzBYBWaPbBH4kI31puN21/8j61Vub8TselytHF8HQSftOx1lQZhMm5UmV4cQYBRpc9pnr/
FWH6TCwBlWFMrMB5VXOOt5U4g4RuxT4llz5wrJxi15wcX4UcW0+A0GJ0n59dhgvxT2I927nQqOCX
6QCTKvXKpLquSEv8a47cyep3ul3ZRJAcSEejWVTAA42/rlU28O0HTQnWoS4xeXoyW0tFId+oQQRP
Bxr9v6KGdHesII41ythUmfHhQvR7kdDm1I60kOfECN43BfPrjs430QyXUXEEGo+8XHOmnkr8iHPB
HpliWZPa3Dc4+q4Vzyu8LnUEOykHkbw//enHLf6uzPtETJINClkQX71SrS6tlrUMJaX5OATXLgky
4ZXqVJg0sZ5AbugxLyRol0VQ3qqwNS/frPC36Ycv/skK1RrA9hB8BmnTQ6x9UG5jie4EMsh+N4GK
tCXATv5QTMJ7ELlOcXgLzKQUS1sLEQBqNXEi+g1bxo47vBHl4JxGy9mrOQzCbmMd3TN8jjOYqP7+
dMSaoF62JIb2ANb0I+rk6eB3KnBLYvZddDGtMBBs4kcQwebXoRd7MjFx/S2kU05cex+rbUvBEOTH
/nvmysO1NRC93ajNs5aaUgM1e4VncIXwrrRpSVMM7sfBDrHuhikO6cT6LwVsQ0Nz8hbsKNRbRZmi
InBIvHn3vGh1yXTABWGvaaSFLZAKvnyN3dwSBtEwpJIOq07B2pvdIBl59hbUbHA+MEC97q833UTJ
X04oIKw6dqKB+QpLHMHg/8ofKggO4XNHodroM3ZSoBSG+csW1WH3am3DYoASox+a6WRgV2GfBWjB
vybXy04extqKGOeZslT7sZhiyaJ2hKeFBI4skucOAgQlQrD7NspS74O0Ned+Yi364hnf6PqDgbP1
zrDerraAzYnKejNZh1Xkhuk9m+yVujCvBFbZcXCRtcxTf+XFEKRmsBoCfp+sNDIVp1yCoAB9m/VE
81S/3kmriGiSR6UFEDa+moKydHPULpSDzaoK7M8nxe4pxOmn+n/uABIYFO6UFGA+oxoB3sA8akOD
ncX1dBO0RH2oVb2mIG5rmcJdZhNQ3HVj/YmxHucl0F1+WDGW+9a0nf7nA88gnSgCNovISu4CQl+N
P37V76zWPXAy4kw02+4N0Xz+L14ljgetlKf/yO2ZjQfnVH+4XjLHrRXq3SLEwzcMYu07m3E1Z/js
XkOBKm2TvKckl2mT3CJ6M2k+gUpbIcuuigizHBJznBdiSISWhLqKZQ8L9wK1QWgnn9ZxrnfCr0ot
Fd+GRs2HEBCyuooOxqcg8XfOw0ckhnvjhjUB7CgKjxdmBP+t2IyBrss4IcQ8xL2SRJbKQxv+GDj3
VBPXLk8mJfDlUINY+RGDxV/jEeRNj1QbtjWPvAkYsolilmEV/CcecXgcC+TXQd8MP+JJt9NnKvEa
djS2su7m2oP/yXC87fWitsc2kUR1Euw1yqe4up+KngqwD0H9cj97gasko5iJ4hJp8URH/M5oGzQ/
qs60fAnfCK8qZaQi+qUWek1e6MxjjK0SXSvXdNZCJKKfinA2akoaalHlScet38GZEXOWemnrIT3x
GlbVgPyQjPUmPxjKw4awd8vTAX8MqMh+/z44c6gx9WbToKoiJA+WcQrQLo5apDw7SMbwmVgjtKZu
zkZcY9VsDc8Tglup9XnRMDVhQ8/6dOqfsMJI47Ggh6qRbT6g4Y/Xth1R6SdtMpRO7DrwsMpplgc/
tl7ubkNzTU1K55r9lgvhQqcEDdEGfmMFg1GtraVxAvH+yoG585mpvDwcTKjpSdOj8faVJfoFmGPI
7kqpqbRvJU7FWCdFHRoLcQLsiuLpODYguKnEERKITWxV8Dflk/kCM89/1ugJzn3d7XoAJxQNsCIl
FwwJaWBt5VSObEq/naO72cItmjsYdXjda3lRMrWeUxWFe5ZnzLpNkhER0PrBRGjvSWX77VZLHH0T
Uyx3bY7XSxImOuEzH1irQWf/YmQtf3CoptECMuMIovh7R/w70uNc+ff6POPpQYKcPnfucwgdc4ib
1fFqtndkpQJC1YNjEuBQ7mqQrayxVxKSEGk3QsVAsaPM2taKGfnkXBVLGxzsPpRr/1HNl/lA/Pmm
8JcCcPj7GizIve2I9dD/5KSQACHpYt3A4sejz3N65ssnpX5DXxPyF3EofdP063GyOIZNUUeO5REa
/eZgeeE8R8nnSh+l+LLGbWwMmqn6frYDvMiKY626VamrsdZuxoZgbHbkGhZMooIITn3Hr+xrl8Qt
499AkfnOaaqM0/rsKD/DavVJWRis2Nq0pMoUenHXynUBS7/lYZdmMYxudz5iY9Oh+l+4zHIrvyN/
3hzYSTT0U8n4P6IpFnioshfsp8ArGSfnwOPl+IrHqewCR863jXOeqwv0rm/RGEeeKbagtA5z6dh/
PtiheDNE3na+O0fnO4BQhHE8vp4rJiDW5XVSHou6c4luVGrbjrPR5036pqMefsM5rs/2mCRT13xB
5nInTNsiBeNHor/RSOsPw7CM2mV6EryicxpacZC9Atxrubo2Z8GFj+c74KBFxWyyduianvJ9YWm6
0DgjBnwNIayoCX9eIGwJ/PGu+nDnuzDDZ9dxFF+rpfeYDloZzNCZEO69DdrvrfJ9hT+ttZHx+yhV
aXRx1vNenOpZt/JDinWbmD+nkhUIwFNI7vrkUlQW4DXC6/5t/a7cMh7xu/HJ4/RZlg79thKnA9yG
3AEEnTco4kVRu5TdmHRjEXO95aFDf/ABX6G30RGCeSN2/XD3YpecZiHuHYrIUSCU2jojc4KQUn4b
ye1CwuQ550S3qLwoGJYyBsmp2ZGB6/T5z/X56Mo6GX+AWvigAzpHWgWCN8ABy0YLSmaZnHJRnPtt
uszNVW1WmpMf1gEEmK+MXNFXiPjfOAGc6J6V5FiyfKXjYSSuW6sQaur/OeZm4cREMxQtJKFq3cjs
xN/DLOsKfqcxhud7VHUEI8NTyIvomwFn9g356Ci+5Jsezbp6VGzG0wJ5XeS6Ii+BWBcHMt7Or58V
SJXfrRMnxtVURNCOwvcT/oyKg3Fi94DwMcuQCUhuwFIuq37b5VuoNw9UBRWJ6tBnF7xetDT0kp9K
/uL96DF/6bdzJZWstgQx2ifwjbvA4ag4ZkN71CcoVVue6QDeQF6CrocoKfdmu9Z4h/3nxSPNvosL
L501DLMoF2cG1sVYooI3u20VV3EVkf2jFwoOsxBLVkhHalhX1rri+9TTxvCdPtqbPSixjV7TiikK
kbFeRHYkWVuZlOsBVIysMafVTF90aMbHWUAIq5c2J8lUHxvCTbFBOwUZlSkLCaZzKZIJuSwg4ANt
Obyj0SQd3QOsMkLCPatcwBDVNjooZDY3ukwoUpjyewEYnddTusp85n0Cc8d64EkaxykZ11GTdYYL
CIE7EnNqxclMzmv6H4oLeDSNsd1/aJx4nnomqmJ44gS3/4AKHTdMLxNdSUoeRZE5wCsHg02S5AyX
uEUW9SAMznP6qcpSoQ/gluQF+dTVVC6HAQzpVS9Ij1SrdbmXrPbcaifKs7fPkPsHkO9Yld2QcgPr
JN7rpiQ7AUL/2Tt/7d4eVgCM5u0OJhhVas20S5rglbARM1q1oEeJZ90f46Kkl+WFnllhF8p4w7tW
LQlMISDPsfRjJrYX3O0tj5AtL/ul/IC4tT7RdMx697yt5bsQg0l5bLrkK7mbevXNP0NDzeAgkt2s
dPRFAAayHJVVgBGtmOVKggFuddjYBBTexN8rJHnqjOviTocdB4cvoBaopkoVxiol8s0vfoquelsX
FERYe43OKC3XJckhjJvmm0XSSvcqoWjzVhXemK3gQWYby1tT+iuXBEZOfU78EpEhzoRFrSDrF+dl
bZad7BbOugrPQe9sKD8Ng9kmvr/3oqKkjOMZph24WzqfGyOPV9K6DP0/tSk7mE9b+IKRPwtXTzYc
Mk2+/zgy1enrI63qtIaoJSOxACE3c5lyqaSP9Y5MYu//9s7kacStJ0Ix/kgQrhSEtN9TVu21uhO8
9SPJxqrTDZNAZ8Gn3c6rnSmVhG0fq1hyVoTGRu6z0o0ETC6znwVgxMiekyNi4Eieb+yS/lbEa3Ae
1qJue3+FlHiiShwUkAdl2Uw3qJXiXXmzI5vIiAjodiQ+aIIH+SkO9y/n+e0L0xHSKkWJjFSRaexz
Skj4cpxgkSn6EVlMO4VscQlva9KJe7zfg5KgVCNXHGois/uivKx2DUzOTxxJ7H3Z1pgvnKEDVqM1
PMKTtdhdJIaAshlXTD9j++fj1MUR4spaeFMzDBFTJfBKPB+1MxJLvF6E2AB4umKdx6eikacqc4yH
jfRgslhoRyTSy1WIVDILKOgbubTVnhm/B6lCgCc162v1tl+BivKfl6iBXhqQv/vNJdmR++ozqoHf
kmxo6EYJAZWqwmSja3l+CWEHKIBelRiNJlEHxbHbCfOMJh6Lmhtie/Ya5EpiUXw2ttGscWyfaFcj
lJg6YW6aNLzK+UXvCAJOhHUBVZxBte0PLQ0mKUxB6+Pu2DOAWyZffwS/AHqsnGws0/kfPOy6Luuj
iXQXAsWsh2UyL9OynfqRBzIKLQySEwMk0+8MXEqcwHm1TuDuo9QuKO7v3jrEpM+2yngb3a7QrJA2
Lu703OCrC3MlxO+fc0JQ6axZBPLHZFjyZ5gfbJVfoYlubpSX8hH8xcN08A+wEoIjD96vSSin2hqO
10GhSuRLTnlTHd5JgP0C83dLxQhKfR64tokJA7SyrOg2W3l2Vg2Mu4Um7X6+/qR5oJ6cHCzZAmzC
ryYLw3ZlduTwLE3NE31Jir8cnMsH91oznCpVu14PKjxX/87iT+JXNnBL/RQnuoaxC87l+jNNlqX3
GH6nBKlIyq/Clf9I6mKt5nnkL9xgujd1Veb8330HL3TSbVRVr0Gfl3CQjsGEQS+cjCaHUjG5yI13
EnAtSQ9R0h+/KURdAVZ5twmQ69kVzVoFvFDH7ZjMUAn4RIDTeroUi7dtkRmTPFzV/Hvx+1Iwk5/3
WiFCLcYVrN1DebOqnFOgGC3LIrcgx4ssFygI+Q8RYYX30EX4CqBMZTLgU05lkuwCkBRyZSQpJaRo
R7UCfzBEVAc+PZiAy/0VscVYuujIHqIEQMNQlep7DDLApvN2xNKYcb216JIE8cocQC02jCMe35ds
cEJClYYSpQu/Fm6cyHOJDAmDFfEKjjP3XG6stwgLKltEBxoVuxUxqr85G0JyIJxDTOPkc7RaDLuV
S6Jl0bQwr92CT2pj3AHqfiHncdb+UQCf3RjjRpreCo4zGpabUiBzRyrH/Y3yztWLPCgC5ICsuRAn
quogRnsmJmpkjStGoapDaHV77VnxY2mhI8qw079Gpuyv7Uq4MWz1lh8qPLvy7Gwv/ShXGoPJob+b
tgbFjs6bzBv4JRr4kv2sLU3OrhndwJ3qHOXdmSv6LFIyXFmBtchGJ0kplAB2uMjMYhqnxZ+5eIwq
ZqIvave7mGVwOAFZQsu4QyzK2Qxbox6dtE0ZiILW8Yw0yrkpkz/y1j0Uch2jjN3IQ8bNZWhysZf6
jRNqv7hAE+2JhPwF/LbPP8VMtsrFqwlnerSJu9N+YQIHZTMzM5tstcfEvVsvhnS4r0haQZCtCxk8
CbwUk+r5rIauCkvdZexU8TENXt2ItUfffRifDDfPge8rBfeqK5VBVWVNJxM8vAodnuGU+yZfsJoS
teNS78/Thz/xwiY6a2bI5ThuViuD4vrIkVIPPK6MNQfNR82C80pUsQVX/1zdmz8uj6UsNpB38y2v
e+ygs76CWz+VO6MH0nyxBjf6E0FneVTlul7YfqEKmNVpvG3Vr/a09H8ZJaeBt9cpsueOITYbFCy+
YSFgyLEgSN138+CXd9pD+vQ56YceoPQCV49qTwZWIsMSOugoKxHCY+omHcs5tsqI2+50j08QsPeE
TWTC/WxSLvrJSeCnlDXj+EDgz3+0527SPe6yqVJxnbIXyQkwFqXyMbWppwH1rA1DexQo4f5G0Rw/
jIqorbDM7g/4vg0cnAfAuihAS3AstnDJQNbq/CyBgk6LuMsaryjL9DhOGfSD4AtwtAt0m505iEtO
JBnLlH9LsD09m74t7zjQyirBzLR+HJxQOyazhc0/L2emeIybpzTIFoHARY5EA6xc0tX+pJxPXgGF
4v1R4geNK9Vs7W3TUa/v3ACb8RhFlQz7O7lD89fGg3lAIuS1eIkvZzF2xXFakQvV1SP02B4lOPmB
2cqK3vwj1QJ864JqQDhs88tcB0H/hZYD9bNRFov9ogFtMdVSFG+lAGnvaqKu9bgq4N3BRB3CKOxf
8rJsijgbAREAik/SBZmkKGpbv7ZSBmWB2w14S+lTKFtW7AIFHZUSKqp85dqhUMkDI8OmS8ngr3UZ
BOLctsVy6r9TXfrqnY0ZGUiwIVxeKu63ZM90e7GXezNgESUab/B/4gr8aAQSfjFjk51nSmZS7KZm
y5WDiaBHdOX/d7GrtgViTxHZU2mHuoKvYADn3fTdvW5r8AQdoqgCZsFychDpzT5SQB3c7lK5GKSl
UB6EFQ55K0wmrwZocqP67RUQ5y74qJoJWMp4Vz8Xv/7g7bW59UhdYyL9DiVzCfgWV81WUxwsAgph
Wq6sBJeQuZBiEf0UIrBds14J2czx9oR3ruO7adMPUP4uUDAvfU42R4wdlzqXpzTZS7CAO1TjdfHL
vBtSB+HxzgfGIzg0DNRSNJSW1CJshbNUStKpH/Apwh/2X0dyiaFHL+l5wDjZr/CDo2iXdK3QI2od
UTcP4LtZA0vcAMPW5/sWKTEYjsxAaQT8ghpUxPrwRaTaeMl3N1lymbNuOByGlUuO/xV2PVL/LZA+
iB0Ynb1aOe8ZTh/Ze2mvDmV87rCWpMXX+MuKdsidO8kxWfvQbnn1PX318zHvbmUnuLfSVViMLRtI
C557iLBOSQrFQjRxTr7R0u9fZ/T6h5p4UMDIDnS1YKk65O9hX5yAHw0ESFtr6ahlUhteVg0hZa1m
504XKP6ALGiNPICMqD3pPlu0QbkejEVmpAXl7EA1tj09xJwDzXEo4i4VjDnxiA65q/ERYG/mQVRb
ayBre5+/+1c0+PuRX/c9fwvQjY275NhlLnPJPLGROd4fOLKcxMQ1nrurap1Md34eZRWmyDGR+E8o
CQsUAcYso3xz0wcYnSK84A4CaQ1Wd6Ew4xZksiQ0XPiZ3fQy0EbcA5XTjZkcYTc+sXkQvUoxE9Zs
HMhvOybkvXtGj5w2FoTDryOIqA3vndnXEir6TngrnSQK+HAfUmUP2iSH8+wccWXxaaa03NpjlN6E
Xr/HKvH24kaWLZs4xos36dh0/VFaHGDeaxqN5XJFaZN/1WbvHfLSjGWoHw9DB6yINqa5JwsT9y9c
R41yrmPAF1EjEa3WewFChNSuxEZmy6E5IPAgpmVm2S6Sp5I0s1rxjCia9Cx1i1eXx78+BoKPUXHM
kBio3x6w3rTHnUTv8WFfjt7kp77mjCqUrkobfxZiLo/oSLBNVNn+U1udPzFIpmhkSu+ShUOfxt1y
vzUWK9nVgFLE1JiQe2m5eqbVIJndPITVcJqlUQy5/n+SKhIa3fZiLgenUGoAV/ZbvqKHGksPrO8Z
u3KoUmAmtI5z+gbUp0eTV+Da6ucPeACisctmbblvNl3ahTkBxBloJpBDHB1/oFE1DCTJumLLy8Tj
bdtfqmLtaA1026urLM/AwT3dSRHwvdQeqccUTZ3pNfsat8lr9dDwIk0PSVr05bCXFXD58TQ8Gtyp
Z1EUmAvQdAolTwU5lTH+XvZRI/BJxcF0hXf7RkgaKk/0KK40j1wmEjxgN6q0W6fS5AT/Qmd8Zrx1
RK9vL1eE5iMoDkmzYDC2wTQuqNUl8Y03hG0zCr/vWIIxm3wBo4sg+6n8oN7cgJyKayVq1kIIubrO
62pyZ8XMCKe7VdKQS2dyR4MGtNhumcMczrqIDjX9gSLwVTxJjOO1TDX2B/61P2KXqQ5L3zoMc52/
ZQi8lA6wS0b1DW3NCANf/QqUbFzMJYDtmMEoC9NvVtKp0et0FGJklCsfm2MeAsY/0v3Y6ICQqdvQ
XiX73SS63aC0RMq6BGrf2/VD5lpln/tnxUgdlmD6PXQrikr1h4rXImn6+E9AwJsgl2yLltPr3aAE
Ky679VXAkpT9dd/hRIxrxDrgTLJ6CdDD3wJJgHdKC2wmy0Ig/AUto+t/ywhEsd9rPi7dOqN/id24
G9Zc5chN1HIXZrc0x5ZUBXjQzplDUgOojWI15ZnCAkdzaaQmxe/CuHlkdY4lbo+nYwxmGDi/VNoA
bRmTP1pBPHsbrXopm9FoGfOz9EZY81fyJO8uNXyghmYfsdigzd7omvS/eTMYHorj8ZiUIMov7md6
PUi6uodpXanDN64S09LKE2ezwaf6UQqnLscWW8EzxiBtEzEkyIUD9X83McDHz57j7Qnn/pXctZfI
oQfNaKzW4aYRnjdR/7cWsXJkD/IR20/wd5tN3C+sk60nzcpNHeCD3G7GBsLhCBOb4+/MT6g1ZVAC
0L7Odq9Ek2sQlXLKH68mSIWjDeCPsX+dgWuLxeciMYoLaiie7QzyGXfgQr6SORPUlUAYnLmTjpUX
hchNkaJSqsn2l7uAJaX9a6AEuhqDcYnyabtzojCjRbC/02yUmZ4u2xTomBIEUKQNDDJz8l8F5xTV
yb/IwliyxPYdxCLxUzTBfMv8su5b09Bbx30BlMd68aTU8ojqEE5wv1th+qGWfxEZApsbaYq0qSJQ
7qan+8YFXoIeed0IV88sbnlMXNvvVanXi2qIcrhwd1U/dF64k7zl8RRFznRZKU4fqo9R0ORWTClT
gQQGdWf/WosFPNbHdhxTpSek2GdlIsWdA3HqXSEUYVkIZPJm8IX0/Y6MTDXtMKY/MmKCUPCBuw6y
pc3kYYKNAs3OPadgZqpdJeZ77ZHKdPf+rPIbI88rIuTfOBUVPpck4xAPNDGXDiS8OMknyLNClCPH
RgqfI5/LVpDxnz0R9cq29HfaVmnIGQBsHWlabnPxhFkj+Ipf3pHnn/EHN2Yuc+132p8PyuczKY2L
WdTGcO/+PMMXhQO6gQNd5wrf0i8Xp8WMxFL+l9xkke5p3/DNc4sUtHy6HRYg7tzambE6xCXCQEZI
e8NSjZvrk5Uh4D4HMPYHp0Q3GxpHn8cTDb9IoUI8gn2PdKfvvfWNuRjr0hMP4NT+kEOrnWBhmH9C
9yBOrhq6Gbmdz2mzC1f0vqYS3qdqmfyb3xdM3INtBgnEF80DvhbeYjiEp8Bemq4dqfG5/+ux+xZP
0FggftN8Kb6qquXEiyivI9uqXekJmhWIWf7G3F7qhxhhkd+FD63YyiEAzYeYmwEa4Thla81GvJY8
0pyCNf4JVHuL2qNpfXS4GKThGf+PtOe8/NMuETScWsE4K2U83x3teA87OsqU/LKzehsjd5mXLezo
Xw5ksn8sxeXSnSLuVap3FYzXorQ72gvh1m6bNOQWmGJEMPag65aciPcgFFXtR7eTYqllo3hFmFfm
7A6GvxEEspiY2EL9QKUa2ozLRKv0HWk+1tBCr1rj5M1mIRzgYLtM/3mZ8hGTsPNuhmwYIMqTK/hl
OIhCUtG09+e2J7IL3toL0+AJ0pmuYUVnia7qde5YiKfZ2LTUBJuyoLOU5K9JZzgB2HyjamsmsMPg
7jEtIyM1nKOUtAnhpNUIp1zwATFZPnd2f1YVUy6ocFOmdZ7ZpGTEL2mPVrz4C5+9DPMD306nX8RT
UsgBHE/76xLJV28WZaAlovlEOXWpAu2Mq5TCd2ujkeFapEg0Nq6d5VRL8oVPUoJoae7obaffJxNY
VhFW4+0XPLZrgK5gwH+2NE72iCEwS+8VFBb6Wl0or7+2xfrbte15Opwjo8WwwPLXlbIE18k4DH1g
+qkNuPxHZKJxlNtWLcty5vIiBkBRRtqvX+oTl4c496jig5bwYbNyW9z6zG5tovb1ot9YdposB4TI
NWXwLwmsgO8FDgEnb01YRWrmFa6YjSQf4dG06eSJ46IDdEch/YwQOPa8jihNWbZXHaGIQvTmVSM7
fpV+mkc2u0qQDDKifXzBUrqYCs4AtoaieNRY6zu7N04OJvpg8Ty1xja+X/dh0XtmIqSeWotRel6M
P2wQRDRLXQ5EYmcy7VR6DSD9B3EntkRZc3PXpOh4Y4ZNa6UTMHUrAefc3XYi9mQ7MZcogsEQMmn1
dMbPvHoUF3GKErU8vNP+FN3QDbcJ5sU9nTLnoGAGRvUJ6LLGp8OXZpGdm2j9KleKZiRNFkEggBbW
8A1tMseq0VGtinG9JFwgI04FMYx6dDwxGaOpGY1i8+4k4umQHojR35+vaYQA9UrE/8Dfj75SL59N
Tp+LFJ14Lr64aKyJus7b1iTTmmIUA1WzNs2vWj0NYOQaPu1P5A4YBFA7BID4h2ZxHh9+yKa1ZXN8
3VwfcZlJwMINCexvF+mWx7lX6HTETdtZ/cNb63BG2yzKv2GYsdeSqmdSGDNu50+mGeIXELE7prSL
q5rs7jw4e9/QPG9nzGH98v2QNdTjyrEHKWQKf5NrWepQv3VlOsmKziv35om89JXksc7H1T69q9+o
xUqBXhkJnxXY/Ca8D9JjWQP3TJdfRMtZ0UzcdSW+NwWh6iwoCR0+0Gs9lQpaKyKH3XqmND9cPaar
GapK700smInVxIyOlMlQaeDve0nE/uemjtyIMxs8blRwL99pUfsTzpFxUmnVTn/l3RF6oH8W/jGu
qrbiSSgtq/bKzFgwAMD65rN5FGqM6dzE++su4ZsInbWdcN6iQjEoKedJaFPUH5+2phAw/cZnN8lW
nLlbPD3hv5up2+l3EZISvBOrHHkWuJyYuXuLfeMsg9Qe5+nlsFFuy2Kq3xDPdQJAUbqeaDf2RKGz
MkQzYSomRvg9jwIwYA8iA7SWpCZW6WYvazmh7257C/CcGkpv6XgSUGsvvpg+m2I924icdaeJ8LYP
yIYlqrn51Zf8qLJIbjRf9AqVHkV2RUijeW7AfDoyu5ufo9S/IV9A/CblDvSHU4fBHU7LJ/aU6bZ5
7wyNfq1xSjrPkmMOWV432IM4CN3g3DTCX3TrTtuZAoA4y/1FT4ap1HLPFn9rf8ljcgm5OnLuTOpn
UYs3W1SBdPX9ND0tKS8MmLmcj62bhm2Cp/kWO+pWsa/Oa8r/IC8v6cGg/SSSriRFqzje4pgxsaTa
Ms9ncYqR7MDgLRsrxcf++78RTNH+LV4lxmyTsALdpcqhU/JIcSuKQl+5IL6lwEBAdHvf4M5j+jmz
ruYJI8DOT+A1pBtmPf3NNkg/tadvYGGbSu9qAmFuxY/mn4cRIVSh3UJS0ou/sm7E+MalLd84IsQU
KQAm5Ebqjqaxx+jb5Upjqw4lVo7xTmdJ74e478048uHwCWG8zszJJCgR2B8En7JkNuKYaSV2yhn5
3iX5qSrMAkwZJ49WS7lwcRBiQLR0VW0UBDotNSzTCIzAYoZUAI5kE9X2wDiLuIFGW5G+ksebuVgF
O3kXLH05aAEyBg/IBfzn/tjltS6rVRQXyAM4p63jeB90YPSYqSbSYgnYsBr6o93B265HvlE2VyGS
IN6JpWbNPaecF2OJPR2I6WGfMX5c2gEN1VGhXT6FntGeX2E/Cf97LBw+n3UmGACVP888N2V9W2m7
0iWXs0wVhdA9w9r1EAAjpH/gOUdV5eesXYL0tCQR4PHfEiUNobaURyKYwZgf20O8SWRHQu24PeDT
lbTnJUdjTqbeR+2ojpmNRAHofjZ8wkoyDebBHil/S60lSDS0ifuq6GIketa4VNNzjq6jI6A8Z+Yp
G59ouDdltJfyf+/oM6XHnZrEoe2W6VoPFvOrA7NbBzB2zl+0cqiGkJ6O0iMFSQvQb7NLwtyoWlEG
Qe1VZVSDnlY55SJB6/kAQdVjtewhVjo5PKk1CxqopO55Gpb9HML8qI9qn1lNOoz7EQLYI1GSXCcR
q2tyY0zDjmdlfkQqWkCIB7kSh85NBkJOMP8SOj2hvay1IpJU2t50ka88ucmDonwD72yWLuCRx5r8
jaRj1fDaS7nvZ89nx0b398m1NPRNVVzSPnAlrQWyvk4lvJ2yBNHfnsnJ7keMp80NarlYe/j9bqGd
lyAp9TkY1Q8TZFJyiAs8ms/dacKfkf1g+0b85wbUFthIEOK9HyuIcsq7SmSycheJE8Ywu9D03Kx5
DJhuwj5+198OFV5FxKgY+WfwF8qXbyp+/DMEE4xGWaANTTz3Hi+YNBlLKjsS0JwEliLQNhRAp3+W
oIJdkJ8ePNf/+24Rylhietr3qQzQFAPrvTpwewUchCB+kZLa3O2zAmS4KSiIQCVzSZKqVMp9wPCw
WkUFpMo5LJmzyf5VXI1g80+Y58HZTDgWJ3imTYbFmHP3gVMab+o1ZJNxNLHT2hpVtH4S41/7XUKi
35PTGXDWQ6Nf+ihm49JvZXhl4/zunm1cP+6YLtmGFa4MtNKJmZ7z2zjW/wwYkEa3K41aFzGKH+8R
bzkgrkZsBJdgyag4ZK+MXoqbC6u1d9xa7H+iydc4e044BatFYSpi7fNEyphpvF5PfbHnS1VLmonA
KYfWVXNusCvQYl70el3D8S+csOUZZwiqweWSLNvBi8U69EomWo41lFE9wZUljJFwzgSTD8GQAEEM
9gD1NQnUOlPwpR3wx3/3eGUaSATfczbr9bRDrSWtLNJND8HiKqhlsgv6LlBQmi3jJ3pWH2JJ1c1t
b5cSLXEvA+gcrVm4rRutmCrApKdHLS1NfSmdTbhmlrw+zdUmzZ44sAaHUvr07tWvFtfPtXva+qC5
+l1ndiYkm2oc3Wxo33oGNrl6Kksn8sY1/b4VePuvUfUnT3DGzhQpMZT205aKHPpu9du3RNknGfPR
IJhENY74QfeuzC28tVqxUCYMviU4aUOMtfIcQWIxJEb7qHtOYWCnSoO/imdhZtkmSb5J4BSSvuof
ORcKXUn9S5erg/0/nRtyEc7nqx3VP/6ney0ionBwS5AIP0RT4dXVwXXqXCkkGHLUX99vaJ4Da3JB
o3Q92xNhac4gRj8mQEECEpqaOsLg7uyr+vh6Uuj9z0pjIoVuR8H2Q646+vaNZe9fzgTwToxgbVYm
ewV8dldk9lAE6pnvsY3Ck+R1x2xH9Ix0mx2313c4953Om97Lg/D9q2zzVfoL6xCui4e/iu64J7ar
4515vOCn67jnMiH3FvakBJiB3MFnVeJIR7lOo6GEZAyQdOOavmKPv+eQGmDaMIA7bRE1F+T15vu3
zHACtH2WGB9OzLaQ7xUaww6Iwq4Cpu4RtTJap+uE/asWpuKixJWwtdhAwHcN6BkdGfidDcPeZ08B
vtZTf7EkVT5BY3i/47cdp+QI7iKo6aK3B7yuSiOIShqfx2hCOR1xv84HByoCpzSsvGKgOKLAivFz
98VPpoTJpfQu/1OWsGNysSqynOZC4kQmaxmMXLF5fFjmCRYvJQDiX/2Z21ARt3Yv5KTzZClcrE0H
39bknFWb97DqmPCo6ngzu1RMxA/7JF5/uPV4oABSSgpbN56zEum4kXJ+D1CRIhIhpUIyb9dHjAfD
KRrWGUWF2E0+KugLv0uRfIO1NlZLbnbpdrAuAf9C5tPL0vwQDYPuV/kyIiPNDU9kehwXHV2aoVUe
ORVyyAepEYNvV2oIkG443/WUvGYDQK0arLV69kzlLnZM0qFtUoQZTELYxb3fenqYpZNDUe6pPBHF
u1sw2eaZqm186UfVg7aUDxCBKPaZv6h90XhCWYLxk4KsLSXRINilBHboPlM66/vA0FgsqLlKwSST
IKgviDAfHCtTYKnung1/EjTbiSPKTgMTyunZtc23tLtGNLRvrxKEyf9PSitVLyWtkum2RR5ds9cm
Uv4U/aKiGg57dCB92QULAMndUa1whnMuHSRbbt1tSjeeNr6Z16lhhV6CS4d4HPhiNO19jmjNFdEx
AqMiH29rDQV9Ut2jcT0BjcNVVeISuh426RIOkE9Y/7iLKG+6hEExJnFLdUVX3I2AfizGIFRzTxSc
2vFmZtghXPc+YQYyaraOOhFQclg+hRgRZ4WjYQDiRs1hw6JOSfWRMO+71+s4b7oGzANrIUl6+5on
rXKvX1rf9wcnLaUySLdnPFl2BaIqIrjhFDdbY/1c8Prkn3QtgpUz46nS08cU0VZynb7npDpSpwI9
D0K31qf08ZK7XP8GxoIFPQJlVoFMdtwYR1jq0iZ2THzxvRbI5G1Uy+2Du/nN1s1F1Z/CPQjd4Qr0
MNlsWseQ8sAcW27pTRUhVadfEd+xQujhDhzO5Pqv5gpIbw7W4osmRcNoKr1NyYZo3f6mERr4CyT9
ojCxQyE9N1XsmW0lzphpiCvdAje5+eRwoLQiMUyboiPndh7u5viNk4EKv5ERYPND9l3fJa834yAK
MrHdkeUqVbZ8/ZYHliya62H4wDvwH2or2q9bWfRVsl0EOcjvuv8un9JlME5ILrLy//jbFq88ecnA
kOPpHv8xcPH2dGcndf/gmS+EgLfKyLWwR8exd32CiVMeXaGubWGKRsVo8SB0fRJdgQBXyPZgs3z1
WLIqcSVyp6swX5u5WDrQbCuDe/VNYTZhn09DqoJ4lAasjXgF35pnd+kpXlBw23dLkwRh/tCwDnM2
znmHTK48jNKxTWK+8e3C1AJD2TQwcqJ7XmJ9OnkfR0TPwcAsFopJkWymnRVC6EyvW9cr6Oq/veT0
5jDQ+XX+kp0PMRSLoYTVtLWHZdc6sO1Mhvoy2TI8Om7rOKW6+3ikEHiFZHV+MS6kQf7Ct24O2SZJ
gpq+5x9wg8Ix/iXQHYfeduVAGzCAWGMFahhcVDiSnanKczRDvG0DBk30Z2YuAA5K/USlQy5MI9KD
HeaiO5AC/CIo33O2ZA6XJ8ZcNvRq68GIzy19r3e9KFKHN4GJsF87GoMX9/6yY2WtarP/4PnRFZOl
pQGnooIAMxU3vltKRntdmixMuCMEL/ShZd4lUD43jXXgoU2QmEC65mMoqPzjwcoRRbwTT2u1y7fB
xkzhYd3E93t/uAa+NK/fG6xfC+9fbQTX+VZvDm+Rb4m2IQDKEbTwjhmCN5aTPmKKXF8VIpcGvv/F
L/N27faHPCdPsA3XHFjPcmi73NpgXbFJORjniPWzsIUYDyoc9EPpiCoP11wAa29p0Tu5u4sHpmlY
T1HeStEKnHUGSTHF9q74LDerKtl7xJay5jVnH2vC4gdDaE95dfcPlR0dFbm1TxKWItGxYNuEZOYA
zHxguHlIK+Wgr/qixlwZNG6KhyrXY0phI+rupf9/Ozj+T0kwSW7K32waJl0G9S/C8exNm3c436g5
irCU16c6DUiMwJ+dVBCPVc2euoylhwHqVmf/wRX2qmMTMynjUHEb3SHY1jOt58+RNmDKCHIeSZ4O
w5Xc4fXtWmi+xyibtX5ku3ZFGYWW1+S5Sr8Y1bKq1Dq1UDt87UZj1RGQxQgIFoUVvEF/D6OfkwZn
SnJdH5COOv45J5NZxFvOY9mVryKQaH+UgyaTAGqOORQiHVnf4/g0kWlCzZAvjRuf9nuXcsyVugbZ
EOfXPn6xsa7TM3EuTAsWU0zZhXaWjnsK9L10XEkj6vLDJfYC0mzZrR5q+JvHDIz5vrHW2cEnRZLt
BZF4iriALcnupYQD6UaOobM3uDgk2+Vr6Vr/LdMggeJa4GxuD7LEgyau6bnwP/KVuR75WkIls9aT
dD5l+xVakT+pxc0k1BSXRmhz/9D6iJTjvZKrA/8h76SNhPR+f1A7h9qEqgYWJE2CajAm44viDmsp
0+5KlFO+9BZrBppeQTcocpvKQAVsgAHO5Zzv4CPlUOQDvm3dI07xCTAz90GYQlQUe+bnxqgK6oY4
uCzvE3+HUBRLdCHB+7p6a60oddgDHNF3BXffmv60ouXMqv7gu2kAyQ+QGRAO3MmDa3NhkFM967gy
rvKFNtp4YNW0ikeJYl4ybBBQYly9s8oUuGRECNNZMRDUnoLKwjQyodkqL+xwXvCaVDGYCkDF7OKf
ovS6glUf+A0yzHFKuCOJQoqXQEfNx4xhfSP/SDlRybdjH1kCyLMQ6FdXDhP0W1ZGpmQGC6BH4yPy
8bQNEL9AsMZl/dhocSmxXvxQrc44ndLj8tH/v1H57foFeRsfo9mAXXs4ULj8ePK7//senGTL4kih
CjnI4y/p3vMfHp8p9c0g7QNO5tuLR5oc+KjrCAdcezc8BIc6VFafEKr3YZns0aS1LArciKNSBBnh
JIv/2Md8shT6A72VxQ6VZxxWpK766Ea1dcQ4xsGfPhyuugvu9QjjXapy5WB3fA/zQUY+Y/64GVS6
4Wk5wDg9ahJW6kl9Ha7LA16el9UJXlbe4RSFe/7A2HOnJ/KhGONUcGc/osC3ds8g3Qq5nWGPoJU3
QUSxKjWfVuaM7dl/RqYJl3XRdf+piIHE4aIHtJqwSDWl1w0zGxJQ6q7obit2XdLQrvCHNCg52phO
ehyiU9OyzTTfmIlaUGLQrQ1foTbAA1VuJQuAP26NRhYLmCMhLoHQnROuNQu6k6K47jXtnbd3a2rJ
u79pS4UkeUfhigSybmCgj+5/qcLPT9Jvn6HUfRYu8dY19pcoY+Afd3/aHj+uAWYp5Xk1ARu5mbJb
f2oxav+K8NHWxBA5fq3drbO1qS+JkBpOkiEakV05HCgAUaN+uUe/5D3nlmAZeAeezN9ZgA6UH1mI
i4EF5hpicWVISAo9ksD+qUQzZBViAMB9VHqaoHALAjD6QsBWHRhZfnfJVBDYaAvZco+gXEl52OUb
Vd+J58iaRggBAoUUtiK8lCgLWiE3HHARJaInoR3LOlg65hu5KfVgZBJzsuoEf+vBsWKrspyFGmR9
1cWk7E/Dn1ZV6FKIzVPwO3Fw2O/lW7XGZMl4aWWrJBOqE1TuT6rwMDtn5WBWr62/3yiP25BzdOLW
QQL+ppqlfqZ3Xpq+7/1SKAq1L8ouhwaIoP9+iEb+r5A8y0DAGbFWJ1EaYWiyK9lGgO6HjGouOR/+
ryq93sg4XC8yy7+SP39EaCA1XO8+tyanO5rPuFwUGCtfVTYJBscHNXYkKVKNl96OED00lhHsq1IJ
km4fAifXXKdv4PqS8U4sUWWKx8LOFvv+VfsaT0+9LVlKmmreXC5PEOUUy/6MwpDCOaD47LoBIDd7
B4ocSR71nu0BVEdRMjoGgEvIJzEBbfbclWr5eCPwgPK+3i4qHQMF24K8WVeCFXg0+082BaTNMWti
LE9S93oVC5XVTcaxzFBozNaIdjJeivtJmTk0O4TYZsmbXHMEPgv1nQlUcvd+nNyxifu8nE1d4Wj8
446kmT/UtlqgqCRZEzr919M8iBS9XLpFH1IbiEjaCUCHWdyfvqko9W34hh7XjqJePWeVR4fXSEKc
NwGvjLknb6rEupJZcm4bQyiIJ2XPJf3W0FHzMfuBuyjJl8z2mg2ifyS53lpwlAfROU3jiF68BOP2
JTk50FYIrR+mU1txfKzVjWrkEOcZQm8yHfXP99SUmbx8gU7WRtENcdgvdQyf4tcPOF2rr8dKqybS
qHcegTV/Bi+44fHy3hlXYGY24prOHnELG5S0kH9uKmO5VM++8l+VHXis7agL+ZUwpeC+i/pbj4PN
xO8pcKQp6mZDmsc6rbJuvacubVyy7J9v6v0AB+QGF1e7DcucvhRxMHquPCrFbjm1tPTnbooEelyV
FVe0OU2XCC14p8AlDlD0LFSq/knP1DgCg2g7vW7jS1iNCn3T/L+ytXN2gFwk0FjuaUA+y5Ob+hDX
RECUrKsjD0zvCeLFJHgksdKlMhwfPPJsyhp8sAoeySPJevbYsDEVImgm+XZaOwTRYK8dPcFy/TSU
88qkf1+JF2dEsNTgqvIpCtD0pwVQD9CPYDEpFNtgb98XGXQlfPbUMGiQrnPAe5pEApxiE/4zanfq
7pWDhLl5eXvwI1A6BHs7JlK2QhS4lsav9WBbFUlECckYWPrdH0fYiz1xTeYXNqUK/SEGZ00MX8S6
0RXDH+UfelyHpRmmk0Z7U/IiWcXG8e73nx0zgikzg9YrmKItMq+zSAnH+JR7c3yO81o1y+Xp3hyF
HCdGPdduKRznlhvs9IwSABPfBGoDOMxrMc2dWyr7WPjMpV+AhOclZjy/ho+btwDY/SMA4r8mc4mA
7hACGopNqHqT4gNp9LE7Rvc9ISh5rMginC2jBjMcx8/u7fMIrXPBirFIsMkNcWwASyiNrAkAxbfW
Q3/YhfHkTd7ZF949Dvq+QypYzSJ84bVbRSXLbFGGShW/7fQB/ylZlHXvi5QIXu0vc8kVX03/bnEZ
GMfJ5jZPQ0ctC+BwIj7oUSus5ceuZv+r7aYq7uB0lUAWvI003LLYWt6U5WUQ/Smg0yDZ+zRk/SWy
10G2J/oTpVTOv3x1IkgH5rm7kMfRCr/dC2JJFjNBcJVQVAi8kQ+NIt+yHMjQ13klxbfTjcA6sk+p
0Fb2bCGeSkeyCj5AO2pyEGKTN936TWV0QWZbWovu+sTOqbHTKZrh86YN7ti6SPGQEynm61Lc4czL
UGXb24Ddwye7d+toAJlMwU5goIapi1ytv0VJrX+W64MT8gEep5AwfxQNTnm3pbr7X/5SM3d6xYoz
9r6PxC2BUJzrJf5gT2y/hM0q2ony9HSXH4m+navjQJFrTMEkYcHO53GqL1qAcx+gqDkYWMb14TNL
JVFRaKYnz5zNImh8ci0MiB6vq33cFr1+yR/pdRP5l8AOEtCzmAislzqJjp6xEBCFcntF40ePXY4B
X2uvUauJbw8REgJ/QZob1tYl0OERyxZ+qm2CUJXCYXXLlneyYZk7/x3xYTS7X3840hlAuTmOFJxg
T6srCZB0MXI2WJkHfCGSUsbvTabmJXc3EqZ6eIRF/Tk/Z9WM77D6mzl/sRnm/PhweWuwbxD2DB9V
OykSLnQ8D+553wIvM8g+2Bcvrg/yOV0jutx/m/FveJSCFHiNAUnhlHn56o36croxidlyePX6jHt6
bUh5iLXf2Kf5pAbq2YUnVo9EeX4zh0+nrslBSvoc1tshyRVUkdZrleCjVkirMrNziIzqM435rEBb
6+6z1mCN8Vm6WL4z199VcZkgW9sh1I8KHa0O5hZwxitUpmFz2wC37kKTijnsDxMz6yXhXEP5ksrb
kLL6489kTke8/aeDtrbD9LwO/p8duGJTY/8Wo+dXiqeize0RD9vox2Q6rTL9D349bND6iUmMIi6+
0hnJDQH3Kfv1qOSWtNqQ3BAMTzpa2ebFC+jodyeX4kDDvQFr5aXHoE/MpBh1nySiE+WRLDhgovQl
im/K5fTqyKIgod6DBA+BhgaYNcfT2XPIn0GyWbh2+YVKzw6ofTeB/LQLL/vEYdI/Xhpo4UDfifqX
0h+5MS3kXvByx/eQu8KbQrViCOmkLzkVciVfQByM42yB+AeaPwrzqwtvNHKuou7I+G8gOag3pXIC
araV5OwO/LaA7dGOlT5GFiEQ4VEKWJxOcMXhq7ZwhbTXG0/W+yEQiycXKidgbtf7//ve71Xx1bMz
CGrV2mwK5ekKlkzcoyrY9Gslw/Xl+g6+D1xLMSCV1yXWbhXLd4KcrAPJVNFuJCrhufr2U4NOp3YE
y0ClIxXGJtLnznlVT00JMPYN+tum7lQEV3xvMX9NNsYUNRSVOcEJCXSBgBve/jX6A+kcgZkXNzbq
87J8rbsPnG8NwMdTumQtb45tWoKR8hlRNfSWjAtyunlTKW46iKrI4KTKP9WkhD2qvwWGMGFGyuGn
FP32u6ud7kE7lcvKNR22eTtaVDsk6BPbOb6q59SRRvL8SlMf9Sb4p+TM4s2Ha45o+Xt0nvnOe0CY
aSv9ABLPYtNeLodZH8lgx8eYTEqB4sh5zfXJLNG4xKcfxbkMNrC9tsj7EZb48ebq/e1EoC8/NMFJ
mUA5SYre+P0zMIH6J2uovzPgFUv0SUGi7kibQlmn2neRO0Xr8b7w6aff8QH0xCUu8sb/QFJRwI46
swFcNszv1AySlv5l70ZXpk0SVSlaQg/9YRcwNAlYp2eXz6vsFvUbhxMWetKsGP9TZpemvc2K/d81
YL/c8AARY5FwvUP7I4T9SoEkgznMIKgkiJHOFrn3rWfJOLdST2gPxrZZC3sizTYpQYqrTlpYSONL
oD1iWhaZWLdNPkRJkUtmCyEoxqM3lJrs1VcGjNkEHgSIEtMchItwpe83ARAHyH3JN34dRALdvl8p
4TikgdCtFgATs3ACHDhMU0bFxQmEVrTcvUsI79G+D9kNaHaQ/04volwKJEL+OeW+2Wlysll33qfx
wCFBrNAXtddhD3K45dRkvZks2XpluBKZNpLC2j11TjhPiu1Yu0paGjhme5hCWuyCdePptuyhwZH9
pu2T8MxvVFUIb+mA66d9AuoHEBR28twJI9PMg5w3zmqRvpgEt/mKJj9HUxXNO8fcvZvEDntvDc1H
1zyVQvFQNIsZOm4ziFSq3gva3R7JfDwsS5WOLbknHHFfyawbHYJZCTY+cOXrS5RrxQQE5NoH3PxM
vSlyzGNGpDXxGS4mAYNIYCpCcNJtjkBByvCTXv5iF1c+6SlZYEes112g8txVixpF4+/4DeOn3WGY
/6Oevx1zjUuyC1pY+Jd1ESsPNTUSUgJPVV4bNzWoHJneDtUAqXSekFUDzX9RGkQ094pU15EQ7iok
BduCZtn2NzWEqSj71zt4xODsgMMqkYH5OP/5zFUC3StJMGTr/EUpkMudWUDQ/FqlRutcGAnzXQAY
jFY4V1if2yolxr4Q8dE7dFaVEmVoLhMvEu0V6k+rZOmq9+8mVH2U/uUlHy27hqrDLvn/a9Zf1X3Q
yr9mgsO0Wg7ZtEDhfETA4K63iblEKX6uHFQrBjRli3ycY+tQG6fsNzYnWD1tWUBtgbpmNffxOQoD
A4kSbLSq/d0Rhy5aEOayTeKrPA1TK4+Rs82GX+Uks/WuLR4cwBZ/KTRNcQCtAcoAJRY1wfw+4hXK
1mntdkOZWuCyrWf0WxQ/yOCQjwYmUSNtBOrBrcIyYW+1pUdhM2EyKS5ufY/sES59Z7jae/VJlWSS
yEpEBapLUGI4mBq6sgX+bISHn/8NTysc4MWLnxcscF0aWO7jdn3YNvWF5dbBbJ8ou+G4Fz9pm0Bk
bv1YwAlAm4NyihWnbgPTt2cOboqYn6/KzASMj9+a0jWjmIkOAY7j6rEiXDXMMSMKFtiPs0qvuDnc
IeMMC5t+/cMod6vdsZ/KwqqZ8N57XJtOx9peWAH7MCkzuPu2MYykHQ1l9w/+AACz6VmF8diHehLg
gZztq4DKNci88q68jfpBvvpeYsCF82PpSt5QrCQFnKfESl1aiooRsQdnmRlUz3d/uDmJdYJPYhXw
oZVQzEp4PVvHcSeACy10wIpmyeVFWcPB+ZzF9GNhYUEAtGTIpF7vdrZN2MMqpON/ryFzR8W66ehk
nbVRDQ+rWPkCh74pOWrzxaF/OV6of8550r7Mn0Xx97+fQtI5xJG0+qR8rdRopc8g2D2ywMxxeGrS
08zNKHI+1APuJLdt2LFCBUGpAYRcvKcFKJJoaaUuU/ckKfU77G8gXRhF44D+MIbFetPvDLgvuqMj
NXoHYBbrh2qQO45MVxJoOjSNMewNL1o/TlHr+utIl3TUNODZuVfWEWjJ6n9YyNpMf3k3g0qPVD8i
ePKzqh2pjZXU7vFhpsv8wW9PHneMNYsA+PXsla83Z6HUYkIaYiznJBQGCrPcSbE54ioPZMDhmHlj
tGX9UrLpLFER+FDEEK3H7mWvpC0uQ20iZ5ooeFEolLu4azcge2Q5AmPd3uMvjWvYqnrWBZJzE6aW
iXaTVO6IIZv0VuDn4Q735l+oz+Y7F5gjmkwYXBkBZ67+u/c6vIab48GXMl2bhyLxZC2B6gJAUBCp
iYUws9DHTaVQqAGAs++FKg4IwNV1njY2QCkV5Ae5Edv6hqDFn70a1u8cZevCtZe9yON+riWm7Fp5
QpgmOLrDTGxRRQgxfnz03dlKc/Xj73HNbUqvZLXSEUh4lZbetrxXFjCmc1whH3URlcP6iq3q4wGI
YaW6KydIcjWMNI8Be00oyVehsTUVQmp+TN1yWK+Y6ebuapZOnYDqFwNSe1XUJN8P1kKVvEIU3dtb
sjmR2ePsxwcmVs0NLjF2eYvRTzWpT2Nlin/JGcEQEeexNWHmlVTjE5AuJWVTq9LvuL5gt779Znke
iOlOR+d38tvvM3U9Knby8UqAEDaA+yZxPNYtrStvyTXZYQVdB82csE27vAy1l3VbBRN9+nauCD7+
EzwdgsKJ0U+6xr9Nf1YAtIx0GQDcJsavr6NVuhu/u+2mpAoSzAXLBjspQ8CxlpDq7ec2bRZ3AtTc
R0qkjCRmxVLw3cx9S/t+Znd0p/9TfoI/gL1oUmmorOw/n2eypoyAZyUaf5Wn4TR1AMMIsyBuPdjv
IbM+eGDk100sYvi3GMW5P9VgRH1S9d/Szcaa4qomXIEXapUfp3c8Bm2p7sSCIxIfKWWL9A0n6a+f
iALgL9Y9/h/FwIlRkG4Hysm69JAtUN7hQYcU+eV82o/wPqOTLYCCTEULyHx6aU4OVWY8t4l/v2Ee
HtDCfxuGhXOVFM6HeWs6ORph2FgR0QXPInwXRn4dtdoAoV/maAXpKbTlTqb1YtKq3ykyh+g3uL+z
4gDlBQa0xaaeBirEOAJvQXSQTYM9q1+DWPCfuoAyFL/OtdNzTGJh/aTHZDy8hVOCcfni+9JTwJrB
J/A3Pxl6MfUUIwWxkze57il9q6wlvC7T9RQH80gqq2utK+y2wX0KXJajTvCP0NRVHYO7cpd1/njN
x9L6t4zSs3QcIwGvt4OV/yWz8yZ2x4iWRbgrJJOOAaKMAH/OQRCrzfTjf+V555nei0RKh24Z3FKZ
dNhKBsQ9uH9fkWTLdMjoNZDAdGbEzvNZd4+fKI+M62MGKj4ZplHJLOcpdzN9nXT5lWCEKAQM2c7v
iluAgK3Lt7XRHdxgmAVLBIYYr/z4hEj59YmOazr8OXsZT/BI8D6C177d/LI0fDFjgNChXgluWMrT
yf5K1Dpw9Ie5u8qxdeJK21lls+hyuHqsbjSzPl/4yAIIGyjE+FQMTwVZDks/wfiqsq5AOhRt42yC
ErriogVrXJ5CQzSBh4LcnSLmfjlyzjotAEP2gEv1VpifOoNBOAkpl6Qlb53goDOQEd2tI/gznSEM
N3t09Lsc4m2uj1vqUKCSoYwy9y890lgpF+pvEqjr88Xf1tRgRKyzA+DC9cStxJCZFm4xChgrmzLN
2qg7UMD7eeXeBnLDc/wuFi8QISiswayG6lhPHlKfwbSDfSzwyMOtgDai3ff2OniJsPfmDAcAEgYC
K91rT2cedwr/5zheqM/0D2xwElcmb4hza7i8F/MiQy2Hh0AaWsP7EIzXgAnNmIrOYySQ1aXDPd9i
FG1jJfhAvgRl6QXllbSQLlWpyqz8kKbgIWoh9NewKrYPWwQIEb58o1AklGLYS5oXGFFtobxIxC/i
rVwS6O2REF+W0Bk5BxC0TzDTa/VjV+LEoV65EpFrCRTxRr1V9sVl8Hp7puDtcV6pEhuFFKdMh8dg
HjE/tVID3nCZLaNieC531+MsHXXm1b66OXLxiGYI7ImLvE5PilcrxagCrCbc9jLcSNfpZVG+hkIv
Ty2eS42TPuAQcjaIgq8nI7HSFjTGQvwHqf1mpLKdtmaiAMATrXiDwxk3+PyAxUbm3S4q9ogBmCJ1
3UBasseAU3gLhPKf4x3gekd8OtURxq5wJBazVkMG3OFPAcVR66g5qAIDeUSps+VD1Y1mmy87BA67
C2rCf291cX8RtOaYKvainIq6T/2tx6SaOA2o2Q2XJdQ2/Aqa4J3edKk/bQ2uZ3wGA/BauXkKiVKg
w4rVqMaLDFjl/fYfsYkKrTkpYGWmOMFyD4toA00i/N1y/fdSHvHdYM1i7dZcjv6TeCN54GHihQ8+
Quyr0sjobXshCKVW4eCBygycvkiUCunlWKPevDeus1UArMKjhZTmvcfolKCxhEtuLZdPdRJfP2in
9e6PwxNTOnwIJcgY0eU88eTrhb+q1Dz5e+csYwf1vtzCFJj0aNsHyrZvVfmwzjLhjMmbUCTkbzFf
4X18CZQGcLsnN5kIRFojKz2eW0i0IlAhi2akZDDU3bdw857vWccEQBMh5btNT1aXS2sI1AW1TVi9
FulEekCi4H96J3JSmCpNhyeMJdu4jfG25xHXBahlaUj244g+sBZD3DtFfqhY3896GdUPGRS0sveP
/umzOPUIyuTM8x4/8zdqWhapS938UR7Tnrk3ABCK4k7zvsg3x+bW533I+V48n9ac2W9GJwC3icta
UWZKV00N2tFzwsn0idiyNO0TiKy61E/HSn3Eu+Jyl4QRXw+4H0mdu9z6p6DLHKKt2lueNevlZXVt
n4RHHbpa8RvOnRxXt3PhyloPCBEiZhs8tYLh7NixqrTti280EB+QJLwUQ2VCFFNScAz0cOEa73Cu
mzc21oIEhI5mF+txTuajAARr0kdHCcBsOGRtDHLTALMWpS+ROWVMfaAOPyteh8LotQxZkSEE71aY
hRRAYMnNEPHt1luNbrNpS3eTGL6/SVJyuZGJxaVRPZRl8Hc9FlqrvR/mfcJS8D9WVurq/clCr2tM
K5jlhGZYKm7eYSn8fi7AeRPhQmaqSBd+F5FOf0MSW8AUZO7mffHTtJquBDs7fLvCB34o+jR4iggh
FW1jOunAQx91weMpEngIhF1BKXd6n1PBtgNRP3JrS1Miy7HUP0UQh/du4iJnlWMOhEv0OC3kUY8E
rsZQkn70zPltw/NkOKPP/nros60Gcj/hD7VoOdMcHSK8fzrf6Ak/KPZ4pEedfIbfD1gSvkYi7MdT
gIa0ZiCGZMVHdEo9wQe4MUc7fLy8ftoXGb/muf0BpBDxuU7wq2lYhnqKW5F1evKrhIz8U9SN4xmo
Co9RZwfCUl+hVGrZbJ22FSc9KQ4mPvGsMQXS3S2CW7gErYuPd1aCPKW0yKmfBfUhPnljNtbD0VbN
m7ttLMok1WzXr2aaEByG4joqPzMnFFsmjZQKPaS6WWEoZO8E5SbQSvM7t5p0eIjNy8lUz79U/DPq
4MSNVuy/CwvZV2jEFO1nakXA3Z862VzLBCfoeRFxmLrOveGB054+rjqD566gvBjEMmvLUNkYNECU
9sOZdS0WQRiCd8MUJkv/VBASUBhtw02rsZqyoTZBI9MLhadMpi1UBtTXq7TOv6tq/LSq9MHw2wPm
PwOrynP7iQAnXYGw02ce8v2NDu942KC+VkaoLRGvnioDeV8rVTf3cJrOuxMcGir3UiNymES+0YWg
0wUD074p8BYRZVWDUVxpIIscY82B2cs+wW4TFNlQNHi3aCIBUEU0S35RdaGqNd4nSSo6r17U0uEA
wv7FP4wSJye1wtxucJEtNz2fE8CFFJLjqjpWUyMvGvtd/tvHUllnAh15Ej4wp5PzJejak+vN5+jJ
ggAITR3xz/lrw5cJbS4HSg424DP1yGNqWBuR3U6sOXiwpks4x3Z6mYKWe+pqlnYOY58n7lB9rXCM
gbTRA/Nwxeqqc/wxfTZgKP1ZlER0FlzBGTXppnHNa6ACHZutn2GmM+ZKnq208bM8EB2MjpiRXPD6
etCz/eXAafj6Vw0ptd4xQyATFXryeJo2kJIEbecAl/5a+Bzgete2db99Bx0DbarcTAk2NgbJ9Y4y
ndS1535Yw1Rqc+fKxKhqLYygl6jprbNkW8CSWXL3bcHPr9Ne9oHZ2X0hajfwLnm1XalIQ00WSWAY
Wja2mUggG3Qhzk8t6nOmajAbROwtPlaZU4AkKXIv+RmPJ2cdRolOfIXHeKN32vrt/gd4SlOxq3Rj
nds+Gosg5NUfff4uA4x2mdH/Jl79syWnf01pLIBFRt/Bc3pIjWxAe5Ydq2aXQiYZ9+5L1jsW45Wo
GNKQa723q5/bsbQnMLyrw2MmTz2LdJXz5l4D8vP7e9+Y+E/2M5xFsGBZXaKbqnFmSrTwk4BNPO8P
C8cP93rrNG1RWkrGD9k7DfcenOMGeQikkcRPmkRZ1tQa+aNueazm3bJAJS4lgaaoCQbuxVWh/ZvB
QnSVrm7ajLJwb8anXWvwrY6YO4Y/TGmExT8cpYsiM5L5Iw+gKCkwCeYxN9m3Ddt25WU3F9q+fa7X
AleWT6YlW8jYK3PAVdBldqFYC1aQji5ppHCHzPn46n9whhP5jQ8vjPoNXG2oUEKR0KCtYqEC/T7Q
7V8Ym+hgkUV0ZNhh0Kiwyro2ouezprzUpXnxrjwoucheArZriEWRSMnZVKkvg2+fQ3uGVEKWWiUh
UM/livFkeG+jxs4fX66yk5+qcGoDPzALkykr7l/0rKws4Pp8yYd4ol0nbDrqmvL2M3CevXiyYVF3
u2a7ueoZfb35na0myUh4ZaK8GQcW2+HAtMVBGGfq8GuNJ9NYWhXS1kd+vHzhhiBzEG24GbbcK/ja
2OmNopA2bDWFUCzOo87O1w2y/OoyidIcVTHcP3TP43H9ZWoXJEtxseutTmzNpxA5VuJF0cjmewrs
zbwuSanH77xLzjuyaWSuTYXJfmTJeFlcdHMY7ZB+XIkYOf20aYPyJTx/OXJ5ikZlxMq5BY7kHQa9
eD/nghdV8rsS33otr8ditf9WbBRq/pmTgc8qTC9n9FL8qlFLLRUKJ/n6WPmAjIyyy8c292oVAV+O
OvYOYTCe6dtFnzjG0vklmzYYfIxtRDZSo0fNvlkre4xJjRpKSzUOPcb9Rs3ORxIsx5R/fonyugT0
huMhlqbLbzu4saZWmeGGBApk790FQqkUWgNOsfYOJQEE+y4L2Qxy0wbt0mRumkPdQCnqhbDBv7E6
VSozvnzk4DKNkyLdKfu0/A2E0u8oR/h4bG7SAqMVcM2IUXcFWUDzrF2d4wJpKsDBioV/dzP+JAc/
1AYPRq08lBzQHDkDvGQBZaJc/owuwSduRu8PzKtuBwLdp9y0OWuvAwxYZOml9VlTt6/RL6MzjVkE
ZuPBA88Ed7kzUxa7W1ifolSdTcBDRyGZjH+QygXaax33XpbfIuAFyT2dPj65Dl8xO511w1qQWgrt
QHJVYkZUo9ZmCFzgNT4iSxHtNIJ+jcaL0DnqrN5Uk6KHPn33BIz3/pT6L6mloI3054YW1U+XA6dE
RuVfkcido5sdE3YMQoc4cGLseKuTFAO13KNvJXsWR/F6Rtcwz0LI436r/0YEsx1cLav0Jog2dz6l
F0U5klV2UzWCdyGpDXqDsbYVjg2WaU9hAa6anC1yY0w5+GR+oS04Nvm+5SIvBxhGLll3q6VmgNFg
nXevVTS0x40d4Ew6CLt6jeK7vtGGHvaiu7mrvdATKQbBStqtFTJGdx4R5hMg3SxuCLBV8o6rn3li
RnslcbLHdWR48uyfl7Ljoul/257Hiswg9XqpQ2YPY4ZkooHxwAQV0WRQ0hwNa8Eezg+CndUbWB7b
FcdL+zHSmjT02izo34o94MXGXGVdqDnzk1oXXeP34W3kIho8opVRhgvpjfqyQlHJ4VqqmR9F0bMU
WuIo2+DMbKIngtgNnkjd+vbcgCOTSVWzyszTHF9Wf0qBUsm6yqv16Tg4IKet72lqVVHPThLXwUcd
3/TWlBQVH4mysEvYw2yW6Dnpl13BUOsM2+NM0rtJNugLKK8UbC88DVB4M+WUTmOG1z5sgapu/x3W
uQoVi2oWp1JBv20JWqpNWb1agv/Brnm5tnWr1WwzLDa5RchmKMdmBwt0DGamNaanpMXxFmSLg/RC
DFAhQjEOsVjyAJ3//08e0TWlio+f9w+0jYz+MX3uLDkRizF5AG1L3GX9s4P4HXsOWaPUZbUKaL6N
nlhIs2aIYxyU5/P9yF2cRQtdyaL1CNC0tcsmj+m5Kw6okP/6PF6lui9P9tdBrzX/mC7OUPOWDyt8
kfoESdaOxkfHrTWTomSc2AEeZhsaYd5D83oxtPUSTo8vLnei0874XO0P93uah8N4atNSKBAHVNZy
jtdvySck02f+py3RkJLTiD5NFxke3jE0uJ+WwoXOQn1jzg7lKb+75PvGvrhunfuU4N9pLa7L3Z8q
9uEm2rXM1y8CRwSmvI+oZYl7pffdd1H45s4Ux2QMRcRSs2y/8bQ8Mia1xgSx1pzfTw9ia/Y2hwVs
pjcr3ycgZAbpi15IoudjU+JPbalAbcAtnXS9b+DoQLfu+DZdCm79u7AavdUTQl7xYRBGN4j0Ljqp
ksdymc11PLI4U8VBW7T0T10UtjGVfL3CI/bXy1hejCAKQzJyUB6xH99+eaVJZPzBnxxvNjRsyeV8
Gr+ZEq8r8a0CrCQ4MLiK8t58Kbt1beYscrGhzj0AzIK1VKymyqX6vY80U5Q6SixtLq2k7FPK5be3
VD7JADEpgqUMWxpSZ0BFZ1jszwK3JOrO+pTUqjBRxa33722P+p3XqwtVETIWP7Lml+gMKeGkSHEn
1VP6B/s/c6wtFxNx0SCsq57UpBg4PJkqQA7aEdwqA9XfIwTLfWsLwDrhRSLwIYiKe719CI0NkYDt
rgXRloM3CxphW7bY2zs3sb9hpag1oLwOFKQ6AbGzrRE7igW0Z9qkbN+Y2VxwKP+eO3jEFCuNFBaZ
mbLDCWCnm59DzTXqaYPccKbgK3iGTq2OjFna7+FgAWtoBI/nC7VwJ3YVm+9h/Yyo+BpeLTGQV1Md
JhJKY1q7E9S0hsdvxNYksw/DKxy4mlsI2Pht2LPmxFxLTOeKRxK5/hXL6XoHRjo9t3PSazz9DIa8
+srTIfKxH0dxMBQqvIM5kShqSyeFF9NLJTnSv/582aVG8oHeN9n3AwYnOeybS8fIkOjM4b22KD+z
Z0oIRsNlE1zMtcqY2xhYmzaRFN8caxz3VvZwYTqZoXlNLAI4gZKMQfOnArCiRcj3rVSrqISygcHU
wQXIgyJn2O0kYM6V2O04CdvTnXXBVmIMqrJa4cktqJriznjbOE/r3dMurOP080I2gZAqOvawCf2I
stpBvfTfmV/3deDKDu0QuNgDMNJTg4NQvOB/fT1Bz1q5nxE6b5Vwx72iErcBN5SA+pJgRLmWhu4N
GCqBozUkB/3/XB9ozTDDwzjbO5OI+/Xiwomu2+vCP5IPzPmJghvzKah8WH/EB9n3kjtcG/FgioRR
uM429DrALbZr7K+33ksQRPYic+8nCBJFaWnqmx7y7IgkWtlOQt7zPwrBKBSKQNLTbox5L1PwXPxA
ssEUfwddnr62SV0L6y+lp+ZW3QVdlGE9tl4++J8rQGI/mpJtDTMvd7P+tb1UMqHhi7GGiqPa3HST
/bp0tmdi+h2s9o5blOswahoea8+TfsOERi+nTBfGSdRRNfHoFafA1y6LNmWEox8iMNTtjWK2ALGd
Ust7JT0UdM6tU3+707AuRMVDkCttbb8CVQRLBPM5YY7PNJ46S2sQb4JJa1N50QJXcBG5lZx961Cn
eJI1bOubNrj2jNmeoo3eAqUDxwQ9oH1IbN6gj9WNLvtuwYGMF82xbS8nMmpmUZgUMKsqPS+4W2mB
Quq1O0AL/8G94z/b68qL74GFHPCAz3nJgCHr1U37K/iRqoGJZik77qPukrcjcJmoVrEb706P+nvV
0tNISDQ+YCdzZwkybl3Ff4ADxXcdSmeXRWhdTigoq8pLZjvA2seTbMobxsWP6NTNwp3KkBijzYvh
6sPn86BrPJBkE/FPpaja6f1RhnCTDqsb98X6oIiXH3E7u5i9/EB5yU/VcrSiMLZBvqxSM+XPROmc
IxUgi25KOMlUtE8nv6s/J2q1WE2PQXSNOvTNVOSUJfFQoQhV3guS5adt/spzllPmOIKqtkt0eh6E
pJS5zHLmMKx6Xwiihc29hHhV2Qq2WHUy9Xud4Oxyq3yPZ7b+YKKLl1lCZ/cqfq9A5Gbcftf/M6Tz
n8RSbUlnH41GKBiEvjzgIfIDYC1ClnD9cqzWuI7M2J6yQrWLbnoibt/RpA3jPBOnlyEwPtnfpbbU
oMa/M++WaLw8LWMNjTN5tb5c6qTKFG//f3Lo+dKZocJP3dXZAE1H7VXpeNJmMtw6kxnjmFNcNHsL
URW81k0drsAqu3XIyrWa+JysmLhd8sqEZEeUFc07z1cKmzWqewwgHOGplA7dFefhiG23JK3K3ZCD
BVsPBimxfZqcyAUXFRTL0T2/pFo1U2kTw90PnAGolv4O8GAWPp24ya78f5aG5kVhAHjEVWqTzBsc
FrBJ7D2MGbPt14fWV+SpJAWN97FOaZfIfJJFB7x0mydu3SmuOaaaj8+z+W9eYE+Wy3LfkGnLZIvg
kWQ50T1rkoItFA321szf5TsC2LQaIgNZntMrXlVJtCZGJOSLnZEZ43F1NOZW1+9vO0wHujTWid3x
FXDgEN32y78uw+iQn7Ns262iDt9NwuYzV3HTKxAiyHFlkuZncQdqKU4j1E3p79u9xBMG6yzY+ZW+
jq4DqslAfQUl2G3CFMD4kQwaoYVamJwRS3+wB2pN6qQGKdMuzH2La5hXMIElsr++8c0h6t9D23Kv
tDDZ/d2I0ShZ73Ue6ZusWNp5aCdnoNov7pszbDay2Wfv6XW0+O6OxrzBlxHIeL5ex9I4kB3ka3KM
ImX3LSxDzVbFehO1SmYgmA5m34GiGdHBww7POULiXzru/AnpumZKw07soOO3JtEajX/0WuNHunWe
JLNVBsZ3jhPWT6JK4LO7peeHmuTg/gCiy6noIvXz0EJPGulAi5y9bzlGXwRPOIxpBBfEjEh7DDsf
8eZA+FBdvIRUJELbxFDm+bMWmA2T6WVgIlE07Dqzt7QDSxGwTiNarGmZPQFimmJefP341be9wSRy
lclPmm3+fEt194cjYh5gkmU98eT4KFWfDqjNZjlvAYiTGmou0WfkQ2anFw0KdK2EPGkLRzNJPNq/
OCovAbgGnQh3FasmtX5aV63Hr09bGMju6x42Kax7TsLcoar8Xp1YoLq/Caou46yAw8FsL59Szl5m
n8sgAWPQoAXSstRd7/+qPgsQDV4p966JjjQhMwhNPgYCPK5W4fdREbT3eu5vKDFbzuqcesYc6YNn
h14KiZ6jrWg9weH2MDz2Ntem3Kaw+mn6TQ9NGwn5V8V94HF5qe9mi2/YdmhAsvYf6ru72uv34uYr
3VUEJtuLgaHF6W8Ovk86cmbhq1qPVw2fN8EnyoFZQlFIWshoRC9yIZYrqFVUagG61dgOegsEy4JI
53KPOW5AMX2F2496U1sTW+P/Ay/f1xIBhlgIuGagyRATgHADpGntqV4C1vXzIGfaqzmvQIbehsLE
3YWXMd8JYNKmNnKSOX39+zgZPlu068kV6RFmZENOiPdopP3vR4/NF1dMATi0uoWRP6+jaAooB/RZ
oa/1185MMpbv2yYVHY3mdzqJt/ls+FLcUje87pplNkvJ/ksGP69zQmsU5gznvRNE4yskeAspjBbm
2WlU0yPfUPgIsv0H4Ul+Wtoi6ngkWj6g7CxcJQ56RsrU8HAwgZuUp0jJ3Q+d1T1xM51ztHZjNibJ
sFM2Ucu09fikmBccMxWM9y3DJrwIUXAGUlqDqMApo4EA048QFeSoMGFSgpQjKYY8cwi0zLRC+wBN
nYpqrXpoQd4R1SxQ/h7/Q44mqb5OKLqAG7K1USM6XocJoGl6QtjNKd/Jt97yUl9gARKkUe8QhqxU
eGG/ElXYBPB5jg4Ov8UZ/eO12xWQW/nBIY6TlY/13f6Pr4zYSO2HVEgAk+r5Uove1T88JBc08kqe
nqPrPWuNFC9X5PuO06wRE73NFhG+0Zrmeqe5QyfTFsbwZYghse7JGnsyFuaM8oKd3J9L+NgES5/p
u70VS03CMFHWjNOXTqk93TEyxVB0jkKGoxrHNWMjF0Ox+AIr3G3CsN5D8dVkzupUvOagPciaEkgn
Kaop7vGwUsJoZlaEXZFr8uyOxs+BxfletiwzL9PVBfdysuRs9JPE/tsXdzT9XtuUAeyAGffcgIVo
2vKqgnQ+jw13nWwv89o5oplSp+DUyg1wVd181o5lvWN0JniaQulHz9VeZ/nL/S0Xfr7XjX/p8y5l
86mDFwkUK2qTkUu4+I9QkNlAXKtclJSwfR3U9CPCSuIIajqYExtmZQJDUmDu1rJoMYdelHSHu1jJ
RM5CkdhdmRaYJdvbs+KSobTG/W1sTHuCAtVvnrA7c4FIw5Mvz9K5YiBrAbcy7P+KW+uadq8Ei6us
GI1mBhRB7JtzfzrAH/12FRz8U7QxGRh7nKSC4vhfwK8pCFGfdohiT1mOfzE4qjt1mg39v7PFARdZ
zdk55dJLeLKs5nENRTkRmZL4GuYUIEKSWLUzJxt7Dn+9kkl1V2OiWzSIuK5ltiTcoCDrW4EnVBVD
KjlRF14T/uQ75qEevpnHFJGua1ucDvJ9csCssoF9h2eEd4ImmiAyScbEDGs5v0YJj09gcJeno/Yr
lxMCoGcsg7Vt6yIsgPSJGpmyPa73lV3kWO7w4g2IYhcFSWGCKm3tsa6Jhq86L07HodtJh9rMhu3K
zdkprL/am3e8NScvomkHmO0ovljSEXH94r8eD5uxa0FeVOGjHNrX8Q0LzLOjtgyigb5lXfSzZ0kF
zmPinOvMHTdJ4TsUXbp0iL8FXHOF5uKrNtAF9M1GMKOCxs21dFM+rQM864Ad036jeqoWrcHLXEWi
2zKjJp/xxgeOmRH4ys+2bXYKAOeSf9c3th35TdmeuAyZJV7AYuyebGJD5twDYT0OMXgG1FpD/i8S
Zxqnqb4L5fFzs2uGqaybEpjior7D2NjmoNIQGwvYv2XACfu/8XnoFFMnK0MTQngANiTaiXiS7jHh
xwK2x/CYd2De8qqBknWd/q9SVO/i5+j/Rpl8KBOnhtLjESeOLSjaoXLhWXaatwzemwzUgNadwf3W
F7nvyeUWBUKC1P86nJE1QBcwOq+nN9uQvgsjOVrpzHyg+VOAwhqItYvxJ2lgq5vawG+8lBDAr29u
NyFf4Z2PqjDp8lCYqIhKrvM0hpjBh0MxojfthKYEJpEtQ2YxWXQ3uSD1ZNb0Y73YS4q7+rQHB/38
o9k9Jfegkty/YDWNOmSEGX9KeuAb0hdrAj+LGcyRodmIOSEWrMZ+8EqsVRltvKir/j6WnH0ZDQ0g
jzcevF2iE49ii2q55MB0IBTc485aWMSoL3EoQsl4pPdYRWwRTUL2yEvF8V3uGsFmr8ouA2vTMBLi
l7nrNdajchRvX4HHGp8sFG2xj/ucQgaUmQ8KIbQwYtHyPvcnC3WUWF9AHrhowAxIZs+9MVhp/hmb
ynHjguWWr6L8dgylsFpt/jhQeUHT5aA0DsaEnikskLrMQcDbPiepyzIzD9ScQi1VZ7bOB41ScZrg
HKyxkPP9ii2h+jQSUAFTf9CzeyV5gDqG1ojSPNHiPcg9X+OLQaccYeiE2UD0uFSlk+JNk8EVSOx5
mKEYv9XajZbOP7bntG3kjbitWkPKaLZshQiSpV02ka3zebksPaatsBIFQVZgkCa829/oyxMa7fph
nQQ6H6BZWC4pQTRBWIPRLmSrk+CMe7jgqmLQReTMPJwkUbZ0hIR1XatyludYIemMaQtWka99cruW
qe71crbDSeyJSQeVZVOj9K3ODm0hCSqF39bEhCl7yV3EwJIsXVDsE1nPgEJgMdH2kZjiqRw5g4DG
fcJs4m2wNOBIikPVSfUkc0mnuqQkX0wjN097Eb2Z5Z16BJ5doA7XnzkkYSvvTse29INbpto7CEGM
RJVcxtL2u0Xxb4Z0dc9ONU3KWlPmltwATpVlldsX51ay2Ym/4QhveVm7JzE/W47yk2wlZaNv7l1L
p+MF4xmeT8aFl+RLayjpUsILMBx+fNsrh0mprCdiTdOzbtpAFqevstmQeDf46NTcCSVCA8luxEJt
ihDguAs32IN+u8YTxZ+Av6rMBqVsinp/aQOkbfQYdScMkbu6Gw5dDUVRwMSg+0l0UPO3UnPNneb2
giFgWKGxh0jIzqp8iiq9D28J/Hg1OqX5puAqxqWcG1RDz6SFv7lLIgmmr+S5aQTisPi1eD65nBaX
1B3EtC9KOzIsfVX3xaqhlXlO49hR6uqpydUASYw/Wr5RC1E4mx4mU6m2yH/aBk1a2DpXLrs0T7nS
Ln8qc8JHWuHas2nNOpLs6kVi35bnem3tK16G0oyrWVk48rV0SrRgSltAohMWb/Yl8u62vy5S6zSQ
u1HrvHdb4LD/erVnJIvDlgkmtg3o16bBdRmL7kUbKg70lj3XeKqyIpCPUCxeYUnXe0rGB00W7MD1
nJIZyaz+tBRYqCkeOVk6NrjJn+J0agmCwzSJ3LBJiGioGvF7pj3qqeZyEDOl14jFr7Kp+AGMKcg/
OfIwpMAW+Cljopra4XCQzGZHqPO09x9ei8riH5ABeX5mNzkTWEQB6zynXPT36IV0i9ck3RchIh1D
wnEOH6MmNVQlxU8/fAEaLFSZCLA8w9skOUNWBSNFd0RPAUzzqg2JrTahdDEumV0wppi+y9uETwvB
M1bH10arKl1eANV1DZhRVYRhWE2D75Si0HjIZTOd/I2dDClwP3nOZ/2WiposxdsDiLgqGjNI3XQS
m+ZuLQ/N80M+6iZQck42h53D7d+RuxLVws6axVa8t4z5GXwi4M8HPnnZC88EBqBc9eLIaYEwNPGy
tu9MLqlVWCQSLXvFy/lfRFVHM2XUIYX8nArtQOI6i36Ah/qbuI+EGyVp/B3AdoPqemc+ZUylJTeP
PDI6/yG8iGb6qemDIzwYwYMHP2Nn6YaT3dtf7ocOQRW7ZPk4e5irwvyIvxUTkEBHSnvKfKSh9TTu
TIXvZ1dOABxF2nbEb04qUlbykeOQ24FCLijOItlzTSB0Rz8Lc+CvJpEjXrELnUUQqGn0xe0JdtnS
Hva45iGJHh7JVd0l1AkYi3gDVc8oqEDwJV+ipZmS1sPbersYMbGHDpX0Rv8Lg2cvtWhgVT6Dpnjk
EI9iW4VbjmdzQJx2Rvy1DKwFFdL5O/xKw9OxrBkVlxD66nPOJau/m+AW/346aRuUoG6xW27CLiLG
Jv/Qg0y6O5wgEIJh6NBGyTxkkFm/XtHRfakEs4/dcPoO4J0gMNBwgUTC98DqPfCXtlwJ/4Dha8dx
bx8NZJygyx0PD4PRjnGg9a7PAtW1bGNIRmxKEormFO09F1LmjlTd4DdTSmkc0iuWomepATBd3ljs
S4PZV0y18IwTgf6YpDZSm5hbbCzMd7kSA4jAZDL5dCTFw1Wp6wKa6laXeF4Tmerx7No5UowwigU3
i9aeB8QyqSTB/onQoYRB8ZMoNqFk2YurF/upHPb2onrK1D+bynNjl7B/roqMJ0k9r3FU/2yqn9a9
LiMdp1RGoZ1XBMYEN8grVJz1uJNhzFIO650RcQcjuFwecGSxMPF9Pl0u/4BZ0m9/6UYqO+PA/ZJo
KMNoazSLIyZDRO3V6NJx6cJYj+WvWdTXBxJdRG2E34a/k/pW+ELlf1eKx6+805JLGkKUTxW+WeQK
3phGBnEL301v3Oo8k8I9BuTxI63G4syQO4i16+sf1HA/ftu58OLUVUgYCkzYwYkhKzSc2mff4z3o
ekJiSFZ4571he5vqCgbdu9xuTxRkDY6kwP8Gll9DjiSP9JxM3+xlMp/3DHJNHUnmLeYyy/cbi1a7
QOMuWJnkuQh8HozqHDTALyChjlAESF6guQcTbAoSXUyY1VZpDZ+ZEkCXBATD5I69BRHSO9dDYB0y
3QbKukQ07vy73gmABysC3MndPm1Z2QIidP5a0DxRBvLCPMQAPFohWp+NSV+JKe9+OgicIMUgo/2F
Yg5KdyFT7wSjiQEFB8d7Cb9FOWcmxBsDNB7KY+fxaURgvjhd0oNMy1vkEsYzVeefGwHswZ2ArWIp
ipJTAbte0St5TckOm7ETLcHPjLUhdiOMooO3AoO5/60aoZJfxrxztJwf7bsjk8JWAbpqSz7iZtQU
SVZNO6L1bWSbpqjNzo0uIXtIiAC6MYh4snTSksWgHieKkZIDg46RytG/n2A090sJW5iQ//x/13MD
LQDkj8NZC9x0u4zdROz5Oos4yLjXA7KKMmGk9YMumO01fKBTBoo+hXX1XEOAT3hcRgWTc8yA8Kgk
d34f/WWLPCA4Qc+Z6L5C4s7O+wWWuivCuqYdi1Vg53UZDdBa3wGqmtS8jiM1A6Y326aGU+3fo4R/
y33GmxY8Sm33GVK7fflMOQsOfl4qS3iYk7QKHyNrFjxeTdvgzZzHpirYbzQ/ag3WDhuxOwO2eIW+
AbJEU8JHvyy+fmXe+ASzw2bxEZU8VtiiQRRU7Z7vOxSkT75P8et/+JFyJoVYDNEAWFDkEWmnXZLG
2UsMaZ8sYTzjZZU6FSRtYctPXn1FH+0jFpWmiPkkPzaIvmWcWohpeydzbV83bQcDamFkMJEVHCLM
haMCg9PM98YpjqgqFi7hCmeAenZ8/I46uyoqdbUcsz4sCoEuQnKf1qWE99HpcyVpXyvegKSo2zXO
gn64QjLMSgXpqS9aDvIVnRwiESgpYDWlTkYZIQivb1v/shQ21G1TYJfqa/FQ3dmcWc6gNr2XZFD0
Oh4QYF3ZPK/FXs0ESDD5rFIFispQvQYKRbL/qFAvhFSQz0Rl1nHtTRzKfK1QpT0q3DofSqmQZ0aE
CrtF1z+JmnfgHWw7j0aUuNT99FXcMqL5xTMFcOFinh0q8pjoAQMspxlshvpu0ABVHZZLomucmJsm
HGb5wwpy1UX0RQwar7v3w9KxAqb1k6FjdLgA7SCjouQD5mtnsLuG+7QgvPbJTKjX1hkiGnk2OIxo
mi/WdR4kRxWCx4RiT96IlUJ85J3lT7knjEi6tnuPYiRDuNXgUFwrQ3ZiGW9SGP/UX+mQkqRJwnTm
JcI23wuzwr3yZKcsD+fGWqMDfrrgU1YKZ5O52NgiaZvO3Kfz2e87JLwDaSfcfmHx+3YEMiHQxgpJ
DNQhw2S+4uOdV5r2NKPV1oKV00ck7imbxgZtSFepb9q+DvjbetczWkaYoheVJGzjaevGCEd2QUBd
mCPeL7YEEuO9G7S8aEQZwHCjykVvw4cf97TpWdKhhfr+F3SXbJKoRiGwLLpzQJ6ChNFkm3eQrKkA
dWK1i7W4ZMN4ajKfTvHs97NNzNCxtG+xHDsZYfEYy/ob2DxnWuo9BvzYIvUmnFFeK4Zu2Faa+2zT
dzwP0BMdLA06+EZGhXg4QewN9VOjj3g54g6ImZcjqSaSokvNqfctLd5Q4twwcOsHN9LaBzqPjM0Z
u/ho0kDTcmgeGDQmjc7B4eiSpIQET8LNHuf67NM5KqKQS0CkHA6dFH1xujVE77DqqZeNXLaL4KXX
sf+gxk8PUfbKcomVIZSYr03rh6ivv8nWPNUNX5aEtE+81Ih25lfV62UkfNfEROI3/JkmKkmHTTbP
aZtA8zuB3pGGImZyHR++I4IHRrHJ07yzrSGARxEScQXRuX4RGicOrcT0HfAOo7aSCpGjY7FkACog
P25vK8Xqb3r6z37Fkwk9jo65U4udOHvKj8FpRAXAKFBYrSdt7zRf/NZ4aZvPyNCiuweCf14XuT8y
lWYEA3tcNoA2KdLEE92hwaA3h1SVwZi46C9IpJgM6REkZXy2NKPLI6s/IYLyEMVRbhRbF3wiSmuQ
DRt5Kudw+dldE+qrWy7wKzWsUPn5MYGuXy9qYeAnltNWE5CVxeStjAcOAKNL3UOXkdObB76WNjqe
h9T8bEB/x1nNIaL3W+4FWmPjTQZNoN827aPSOIm0cvJhfNRx+j87SUHea6p3P40MDoVH4wPMwJ2S
FPnRiiPa2w7yB0LGUpoyezsDRklzSmc/Cz06bHsWllVPtZVRhd5Kcp/jxT9pV+KEuyO+681mpQr7
5fFHBdAyzRsfl0vqATqKe6tciwcA15/csAgK6WrN4yRe5B2H8UI4wlUj7zLttKwwTB5siGbcudTN
buwmWvN9OHZLfOKYONguYf3XG94XPGIamTniyN8fNJD1yU7P1GMP+U5Xk6Z+dDX/rPwo9k0hzP6o
tee/WK192JLAcMb+napwTKXaiHUf9tlV6oJK8sdWwKJpD6QTyDqejqQue8Yq2O+5lhLj+BTMmdQd
19BQ+inM3VGPn9QhnNie0hOTlSAGNKO4ybXxNJtD62WEO9RL/MCHFzNGc9V9UlAvhbY+WbEFLz5J
Z5eXiq1GOUghTQuuXKvRhIp2j3gx1TUsP83YGjFQtUVNeO2ntIdTpcIAfDxXhn8yEsyqE4Yhj0EV
h5aqh/RSmooaRZvCL49vklWGqkwli7/hss+VaGPJIS1qcifaFEOaduoDfcIcJDxonCX+QosS3lly
4FIgR3tP/i36UtS8Vbvjn5xv4lY4AO5Q/C4fB73Y/l6ykiz8FX4UQk0Auz42NMwfzmgxWYK+YHXR
s3lfdBj4NFw3r28vEvCx/e+WzHyXS8Hx7nnfSlIv3aSJh7OLdoqNQfUkiqd7AOCQAYSHg4CqEjJZ
fFJOGM8/LhbU/wIM4HaV9vjbAx2+zHeZFctoEOFoxbAwvWjAveIXfT1vdeFGfwXwP6W75mAtW0yV
C5sth8fvAJU6b+S5u74SFkuPYUFj/kxVNnF7lYgWu8rnnjGB9516y5nZI1QmZMMFvyg34n6foUC5
wOD4JPJq0bg2+78N6VqIPGK+kswR4Tt7jzs+/KNVBne7B3Q4Ep5X94NIMrHVu5HnWh4L2G3F7Xrv
VjfwX9mIk+clG7w/+UTEm5HXr5U3a21ve1juYyw7wpPubJg/aHU6LptPoRkNVKKIo23AogvV3v4v
nI4fPggS7fVcH3OKRJz+c3Eo22d1bpu9eQTE0mYXAmOWiL++cJYNenxDOBDElO5IX18r6LuNaDC0
Fo5AJhW+FiQCK/rVfCupNobN5Po6spKZhwr/V43eSNeG67i4z634MbX5wwAhPaUDgFb8Yohhq0p3
y6VYWboJTl5Ne6QBJwd+iv+GB0Wz2Xb9dy4RrDWZQjvEr/hzPDKJvXbCaWT5OmNdZJB9HyTjnM5J
e4Ya4g08YGZFmN1IPBEMuiinq84LHYaH0PZbzRNPY1V1gaKUsS0Ya3uCJBqAwNrwkMUVbOGK8Gaa
1BGl/UG3lO+C0eAbgXLrIHvTAjf8YDoCXatku/0A6yhfCzmCy/la50HyaN3v6zpfgSxEFg/AznbG
ROSH0iAPwf0AsW58AxIxWdsbww408iG2W675KapOMZnE0dBibDrnFUoCH2XIeUMkuEUwGnQIsPf+
oLAWGxSPhQLsworBI0LITvboYqviPpgR0MywFFqSXga3KjjpEPMgjrfsJxqTkWln2XRTOkogsfhK
AWYIRvps3763pTzuaUv3iACFBFhuzw4dUNUOkvYYc2c2KEql1c3KDvOLntZI/ZqvjdN+RF+tnpII
7y1qeeZxCRNaQOMOXEjA7Hp01phCWLYb9a5Jb6Z8S84DCHQV8lUiiIvsK2gLKHy3BlU9x4g8gla4
02rfo2jgFHcEIBnAIddAvB+ndvVNtE0mNBmILtb6dg52gp+R08oG9yi15rk/AO9cqESc7067kNR+
gdq2n/RQxpkWs+gtFHuHk3y7CA7bIOg/44PfLovLoxvkv80HAgIsOl27pJ2VJHKH0J7xQyDUmozH
j4cPIye9Eoq9B/UUvT26Ta09OYs1DUhpys27cZL4k853GyE7mVoef2kCQJtiWqtw7tlcjplm//LH
3mXwDQBfM5TbdWjv67z+iQAxcA2M/LEEBJNAw2c58yaiopa6skgCZrrWWEMst3TdfDF1lH/hZHR1
5GoZ0gQNtPQ/3BrsIrHW2iIIfqPklqlu2qbINB/VAF8Lx/VtqByu5jTTh44t7rB9o7C34L3EvI5m
hVbEwKntPYZbyVM2kVLrWGSkpCa6Nmaualc1agnamy3kr5fCTLqRxvlp/34JmKr9PziLCqi0Ggx6
ED92+M3mxW7aKtt6ag4KXSPifedcdfLtrwc5bXjtycWSbgJKn7SYu7Hs7uva3w+PWMqwWjmPu7xr
CYnvDO+HUqS0Ccqz4mqoiIq84I3gga4dt1CRzk8A4j9xtfUR6Ch4WYIiNTibo4DsCxdNmGGpmvXb
49NVWzR8kgh7CH4pDzXpFcg9VholOzT2nrno6zu+dZLFZvro5RXovXeEC+l0jqeJKPSCuAr5oNYi
24DfzRj3D+GF/uUSalm4fvj32e50Uc+YwE6xwDgJtIc+YwBLCrNn75tNjFgnOtf0MIxtvGD85kdw
347dsJ2hyb0BFBvJgpqpEgxwKbYzDGXvsD3DFaUJi0eIyGWjw222az9bOChNPhnHCMP3CHyjONVa
9x23n+aUHQ7/n/TStSv5UO3r141UmGpb5GiBaORX6HSd/AT/tdO5aRT8TuwCqAL7V+pUiGZhPgL9
Br53Hda/5Fd9RcXGarDXW2l4fOTR/Fw6p/LQmzWEkdwB5jAGKqHlboStxQYpb1ZYWz0FgI04a7Nb
+Z/uZHkR9M6j+BF5QPuy3boHc5Bj8BIJ3D4CNmGVoL0cD37tj8bUSuPUC76poNHTpysPQUWYI5bs
fEJQ8j1IphcHI7D5UgPhfwqAmOb6eSGs9XUkLMiTg603A+f+ZbEfjMalSlN6a8JLX/o2r8CPGhIc
xCsoEPPLv/pXknsm6Y9HUFytZ8LEFaKsOrBNvMKwOduFiXpZXbZBQ+4jmzWvs1fdQYI2EB8YWb6W
0IgG08I0d7EfXb+MFVSlim8szz0fdEPeXfeELc8qF0XsCSjeTIriRZaJTKC+P7jwy0WbtwBKFNqE
UcYgvxtkF2Qb8bi+dJvrxV0ZxBep4kBdm1tmd2vABCfUe8mximGHFcZ2nYrYBLGCkYgRvCD9DhIL
tpTblzgLdRx3U9AN6+BrA0G7oxYhGyk5TN1aPY6MehBgY0naAFdXDKdjeMC661fWDzTP8nTzq3dV
+dTvGDnPY+bfEBOF0meZssBVoLlbl2RB2NDzTYGNTqcJLklFKiZ0uT+D+xczT5OKj4Zqcxo/vZh8
fe9B4H85pJfibdoKLAv6suA+BPZICjtK/73sLJdEtzjVQLZQoVS4NEqAsygeuNN07mdyXnltQp7J
VkwUubSxdQViYDqkEInO4cw+3HiYZgLmj+LAvLzawSOd9IlyPdMn5/gBPyUcjO8E8TcUnncX9d8K
cxcIBDLkWqRLoERO/RNxlUPDQ1/HemUV5fCVmlmhM/GMYKHraDnHsZ9XGN7fNS6lRhlP4awJ/TFN
mZrq96K1D6KIoR7WeUHQ28NBiy4P73DQH8AJyW6G5+Zxl867j6iicAbc2a2rUDj3LSN4YyAK72WQ
ny/UHjI9WNBR3pOpbbgBkQkB6jI4SUiMn6CVQAmStVbF1Rt5JpK7O0w7mhhB6zpdSfng2PCvw6Xu
iZa/epB9zVyL2in4vuvpUXQnT8gYHKlo4QjDtiBnOqF98R8jD1gDsokUkBTN0RlyXnqmodu0PT9q
Ts1qDmwnJizQGWvxU2NXfDmMNeqs4u8p/osKddrswkPJDn3seUsG2haig5IW2/n3E8uE+Qe/rRt4
5X0KQOKoeGKVqDaO338xlXsgatdCRdRFvSkI3wfesPwBzpw6MfVgLIvrsAZ18TwR//DN5CRJm9/Q
E98r9e7v+4BlsMtb5SMy9Ym3qZR1HeXGbYO2FisnF8OEGEz8McpeG4jefF6s5EOXTimtiSHJWn97
gfPqEBJHNDSWhBGnv5P6UZ30lHqbkhn7mOWtM0/gV+H1nciHqHG6GYW5rQYL4jK/sf54Kmu4cJJW
HPQ8WpihPwa7sbhGLKjvZOFb911y0i9q6RbHyIy8ajHtIhVg8Oth2JeWzSd5QZn14AosD87mCCmd
fmbTxa7Hek27bB3sYPWp+JqGEbXwUDrDXfLS2Hhw6NMymLj4ZSfc3o6BNaxWyEp4k1Oy4i3S9II7
IS7gpmWpaj/Nfg0fUOyTs02i0qHDLtwGkOqV3AjAUmA5MZybfskc4R7wdghw0nzo8OwndwfpuVyQ
/P0BU31xgrqzs6qdmYCHsJ2qF7LP4A+dju3iwDgadTeWUOcoucY3KWlYhLTw75HlFoMWGkBiVQJa
JbOmPmoEzkiwsvInOSYdPm5BZtwiItAxRzLC4K8kym6laXcmfxeDfNzJJDOTntG6grqgHptFQPsX
dNOdrHj9J9ghyNli46FBSohjSOjuIOoYEedtdgmEr/iO8c0QJQTeRgAazkwzDnAwvAYCFKls7nU3
RO+a/RWvzn4mjtwYoQkGy0BA4Ma1UR6+0/l2nCTxEizHAu7mVD7d81nMJoiozPZ9DmxodvpMj0Dh
DyWQddp3pCM1TPDhiecXDtqSimsIoH/h5RhKNryeF3CxkvnZWLRlKc93nUpZIdLK0i9g34p0kIaM
ffqFJD0bJ+Da3pA93W1fK4s9k9Xhsw888BHQR0boHvU7mW+4mz4aGpgd/APeCeenaN0sEsEcFYEb
K3r1sY+PHH2/IWiDebF88YXnGGGtR28843ey2nGGOR73jpDBDu4O2y+sg5wALLs4N+bFf24i1FKE
dkiY9auc7oCRLAykG7nx0ezLB3mQoEfpSDtY1N655sOkyGPzI4IUuOZs73jn3RP/LXMPaXBQoAk5
JPcD02N8AX/9ARK3hyF+fsxb9KPwwhbOaHfRFPaSPjnpr9gpyF54pFuswwXmE6od371K0tJVGcEC
FGay+neNYKHImMs3beuoAcWNnz9jHB7z1rSPC3m63vvfhmXxT8KTkf7Uqrzgayz7NMWcAA6FU/Mh
KFoRafDnaSEsIQseKK4q8O54K6McASiHBzbz8f2MmwnqfAy1gXgdNk6d1uIQKEMP5qIKCwCyWoUL
hJHB2ErsYQH+vNV33MFWr/JFu4StZImv5eiSzidJ/j8FsWJCgio5wRFUWSemITYsI1l0P+NemMB8
gUmZhVRYVhh/YqZSN5Gd7RKdesxL0fJ+eQgp7nHH7oj7UwS4jTKYRtq0z8iDp71y1CfsfPRXd9Ka
R+RwJirb9yaLtqNti7+uWBP4guR8eo8Rc3NlECC905EVv4L5Zc8jDHSjno2LvMNoJQDoq2VJwko6
OpjQEZ6DZJeeYXKvLzO/rvpyznnB8TKYV5k0j2jmLPTGJPBQFLQPd4cAGUw4cde0KsJY6JN3rDtE
6i1IgvhJZLutE9RgZW+F10NMTQlPjNoBmoC81No5YCE5AwL2KcxFVkX2Sc1Xz5LgktURnFFyDLOE
W4y+dyQaUlqZtYsSuULwWXr8y2wV6JYqSjoo78VHANWbzngqqTpRE6UL5WAjNqzVbDxfQVOBTr7Q
LTRyU/KQ+rnJWs2FrSEamiOwtVi3RgO6s6lBH1Ujo0yO/4SpbLIooaK7Zo+8dD0Fr09BSShs3IXl
GEZnmZyneq4qkNcrJejXEsdVhHxNydAod+XzGf/fi+KFFkQG6vrG+PLNz6reQKL62yuexBjGcgFl
3aZYjZ6LGdAXONm4LnY+cob80tlBq2BSEr0YB/dOY3u6HFaXlPOfglyWLLBjlrwqpLhjLr8hHpi9
AAT6M5zMmG31uqME18bfyLMvUKf4e4fdh4fwUdh6BhXzzErU69QpYUf7/rPqxF3rXVsyVg5ociwv
S3AwCxVXQCNT+8K948EGTOlW45BYIisp2UUSh36vV9AB+er8H3nOBhxvCZOOIhGrPv1jR5kkEziH
oikefyeBc0qv8PJhtqxg/iAxP7ce+pP4llou9rEEp7AJByOBG3aLL+W2ZxYMnT/uOlpuy+DGbAfe
B/KbtczlSz96pj//uExZ5d8V7WjSbyyganxc97dm/79w+g+v8C4QTYT7N4+xV5qWFGe5B7G/Tc0m
3rqxI3RUzrraGyesfSxcQ0oyrmOA9WI+bRpcNb/H1E7jYqu7QbejZ8XVCpA333tuabCaiXZ9klSw
NbYv44/QA7zh/erbUui056JEm/AyiD07cn3jw9R+1VG2Z9A7XC4oEc8/ba2aWjbiKZSeDSER3kHH
RxdCGVufA6I1DAPJvBVnpors1/QjeNMy0XRPdi6N0JFLiL7SXx0XbkXsjLfBFcDKLQnb+45alLbF
KYVV+pqdOKgP8JOn9CyGY3LzuvNlFTXdNv3/1up4W4RXfdBbO9FKsS/++wDPM4bOu5Vj8V7CnSfh
241FPU+9CHxJf0k3aqQsR1QDkvXRZBKuCTK2ZG5bSeZmuKVdA4mWC2IPGqb+YD41Hk5TlsbgAY+f
WRz09eKrpd1jJCVYa4Km6fNF0LOm8aHWqzgXeP6YxS3UUUq1OC1GzlhCj1ro3oWd+Gq3f3G7Iz+d
VuWwUXkOatAcSf8I1kUIGOSyu5XD79tRfwJ7DIJbY4xRpEL3s59J+2JVxK0Zo95o7pj/myVv8AvE
XB4mCec4WbEQcc5muFM/2mMOM1PVK/h0npojKTU4c3CpsQFoTYDib9yOmHmNWbo66DD1/OByAQs8
Psz8NV/X/Py00pWhE2YGbO7xRa0aBrhNjPRMVRaanCT4JfPmhrtADkp6IRT5z5S/xwgixBz5LlUk
lYSqzKnXFuHRS+elYAil9YIE6ruGjAu9N5Qv2Paz4Eahjt/pucLKM+U2n8N7Q3SwlvnfTJpvnnCT
ptVSI7vhZHHD3cP1pg0d21JiDtdt/sCH1XU38y4cKEXcK5Jmop5dvlvoGJG1Ty2L/rguT9zJKl/G
Q8Zmm9gUTKlFUXYQJxXTEmr1eTTfehKuXLHpGx0fI5RO/HgBFtMl5R1BUZ9eFRyaF2uTwNzUV1R7
qC3AcogsVhfxl6AiZGwliSiHzfAWbtHTU4EoATXK8yxoy14SrDLfyGnohr/1Fjdqebbl5zq0rMNb
16xt2wwu9QbNscxUe1/MIpG4T5Os2fG9cvKrApASXbwDqs7bPOXPnlWIXsbSUErOVHGt+PbKe27u
D7h+iIT1UA0oqt1tr8lKPhn/dnQKiSwVx5+Rz6YpIP8tGjXFrUzx+TaAoO1gfrb6acNVZJ7sEnWg
6dhC2EK7rAQaNsdbvHTgqU713QYjCRy15wlSGwcqfjfCG8r8kclrOKTUlJAhEgRKEV4ODRZwtt29
+mSGj/utNnSuMtPyOsN2wfqb3+5DHXMqtzi0m2FX36DZQjIazBxRO8Y7DrmSdEyvpp8VKOeylVUi
+yAxy47VIOEupIvSx4f35NSC10dd+kqrUdgcksYd3UumldHAmMHXTnGZ89k2kiHumbLKZSeT+NIw
p07tldZxaNmElj1MWN/i547GrIrMhOzyvI1ZB1aM+/80KO7/WxlH5ljTPtryODogQdn2letSZZmJ
l8dcVyeGstPK/Qdro5Yjo8bc3zv9bXym6gY3bX7PgaWqKCCPDX06NJg91VRxuJGydYIVCXz7EDBD
Eo4QuNV+viC2l4oWq8z8qDoLKasIXfsjZqi3iEthFts2vjmxzojZy1qLFGhbU5exvpDLcAuVwV+7
Luwrd8okiI3U6ByVyij+EMys8z3nnniCjaxtYyuVwUpqNszybUpvMNpgSBaWoF3E0lQ2OCCS/fpK
SPmrL+suS2nXoXpjJm4I9KPQhaOoFeW0Ox107COOhUJwKnul0NyDukANzV2OkiVLAuD+yTL2/usB
yKRq8EvdNqsxbfFKjUoehVQZCLt+Cnw+YdRMbzIDCVtcKwAGR7bJrpCpXOnPiB6rJ/paPwzO2qKx
T4r1dhA4oaMx50DakOuKNMgu+/R+ETPNq+H2qpd8kKVj299kpZz6c3HiFAGezkt1pYs2SX2ut7MM
K3aboljVBCSCDfq0TRbfY/E/96e32/t/3nUc6fprPrTNqgZ6z81mkaVDzikMW06zhbfn4Cp2E8m1
gYWm6GKUXCoIPNLUHrlxUDWYfh75gM3fdNh3+LXNGstpkvBNBJCdJtl2UEgOQJkwRILXxbncUey8
EIV+5tq8ZqtU7cg9PDKlBuJp2kTw4+LknOpTLyN3ItggRYHbYGeqql8i2CI31L6LM/xLh35bOknb
E1ZqD7+v9LkrrRToWQeEk+7pUElxLLTZkFAy0ulijcSFxXwxHw1uh5QiALucCcXSQ+fEZa4UQ6pl
/HPbR37bvsrbsSt9GxLxT0+cZTXqvabbydXTx53XRFMChzKahAn44pII4XwKzhv2xP3ZnykTF0H1
KCglck7C02q/0XeQ12vucgeX79bW8AeXOBtvKe2ljLzDWJh4uCxeTq4k52xWlEObtg4ehE2b3qe4
b9VhRhXR97SZ6p5BeoKAcXiQP9bFdImcgte9aSnC4m3P7B5RTVSyAJ0+0WuJNbz+eZt+sMkfVOHv
DXUaPZrQF9FOHOjqzbApRJTRmUs0iO2UntfHa7eVTwTznzKAdEpXa/qpt81+Eko1SCXJBAObzkpz
TslfFL4I9+7z2uv2R9yeqMIAHFog07zo5hlF2QAncr2iLctk5ck9Fh6QU908mDvxGoA+sXaAYXt3
m2s1Z/U+86FikqmDuCGaEtRw/7f1tjShpQIWODLYf+liloX/OexLcaqTXQdpxgnJNsUGKtrpF3tL
VYli82DxnhE48+dM9P3LiE95Ar//u+rFgo9EBUiVs/g4dL64dn+Pw+/Ih9R4kE/qrX8SHHbIdzfU
GHhA2a7zrL45mEuNxsSeq/U9mwURkLVhWa6k7OkL0ggQdN23NKuqU/bsWq0I4/H/miRdjcJOLcGt
9NZQd3rgnaA1qE42ZWSk/a7UvsKwzUCThhL2aHLcF7jbkztAkV8yqDMRMoQa0HffnLGOMnMurRuD
3rVeJ7YbT7um1SiOft70eusOeOj+fRT+F3NAjJMY3FuS/2Mh/d6BnoNDpY8IoAhnogwR6Lfp2h3T
viJSBAfynGP20qk6DluiOtxqocu0LwVTt5dUHEadsKn3TmUHUW8ntq9gOy6TeIrQCx9B4fsFaWHT
+cLvaOBlhroVBEa943Vxyfh0CrQgKifpa0sShi9PLyN9CE3kpg5Zq6iiUQrmPAbOxeuIBHENwnIi
7pRuAVMynHJ2h3+Eo4WZTHP+uou7egLYWwBy1ysEed7/wyHQqZLdLj8lsQ1rtUIY7bl6MklUdQpF
9KDwfqxVmPc2TFevzqKxv5Eh6MYGDchS9GQddXTTLlCMOJnjDLpUWz4KBUZd64kJGjqC35SWW8UM
ZPDpCsldOP9qsWNVpc/v1oeJE2SVjRDO326S2qHOyt9S3+FJK2gU3bNEWr6Z0bnA9fDVlayosvCn
/e7BR96/SeAr631CjtF23+IM3Ccnj/rdKpm/b2oHDPV6wUkd+KbS2DfaSuIGdVaAAtj2PRwPmzxO
/c++CpxfIjOGkP5py4TYEiG5ivGwF6PXzmAv2mWXmqg/IhQtH9jRtLWvBKpZ/gvRb6UTGhG0yEzY
vZUFDqUMnVtwYI5mvUiWu96rddYmwmj5siryhEiM8Ct7MePxaFFe1WrWD6XAgATMJuRN2xja0URV
WZxVWyUtrmQexAqTo8LePLZTii6c62BSMlj/o2B3HpB0WL+iX+UIbuaFEKVMz6ncf6TZEtWplziF
A+3W3DuBuoAF8lTWG053TzL5PLs4ZyCtoposrZ9qWH9M0/OOEVTPkdrGwIbPVPDl4XvDlTMkIbbI
LIRScX6FoEdrbX4M33unu0qtK4336CHStIyNQfNwi50OQ4doR05pHNilcmaCpgAWIMIlVKOTGpuq
7OkMWGQbEypzXfIKIxC/cWqzle/LcLkwcd5Fej0SjOCpkTIYkHj5GvKyFRV2Y4Eb3vMfOaYRQ5xB
e/kSIVe85XdRwrYpuc6e2CCwzwSNq4+Qag/LiRon0WTUOmNABb9lZk0sw1s0SF2D1N93AqyIqdGz
mEEZNDFMTnVAtyv+UNpVrxCrGWlpbRlBkvb2c4dUMEJpbcsP9WTJ4zwRSIuhkvaCsXsaHKBA8LP5
AK85Z5HG92o4mFA9J8N//Cu5lWQyUb1+1nYWX2nedydbK3SrduFqkOr/AH6SEYPFJT61WKyWNtdv
6vBLw7HxZhL2sBaymO2US0hRIeIuSMT+jB/WufKrD9krtph/ik/KPqdn+lRrSnqGm83YJcoYY8Oo
oxqSFh2J934j9DUknlrq5sVxZVsCGryMMzrTPwO8kgCn1Tvw2TvlmuLKjCwWkFxzdIUu2mPdKVVF
bSMDI9a8KiQ58hpgmLOZcptxK3IEaX0WrGW7kGLu9bHzzL0BVhsNC5rOQKzZOwywP6td83rZ1KeD
qa9WIUPuXflo9WkIpS8Zsn3rGPuuO+z7froZxWo4szleaUy9MD39V8l8zac7x8ha6ezxppmKnw9f
WP7EQC8vOCxnITWaqJV/1uzuajzNfYoVx0Ih+t1BOYKWqQUBpjXUTzzZ6LsuSWj7HPQXe/RTi4Jj
zlb0VcZrL8Iz84CQVVxpR9278rCZHunQzoNVXa3c5CBHL/SImHNXWpizckemAmI7RJZtblBUe7Q+
M4abtfR0iMk0NEdhnN1/xHDNPOn1R/BkZXEapTdyxgKY7XGaBKeK0zQtEGjAMLKgsk9vnjDP7X2g
CYEx7NHpbFoPYbMRCixHiXiKCVdYnL7JxUlweqIMCrOGiz5S9IrooAnlE2undlXSVZK6vptPOAEz
M2iLxOAqIMNopBASt0/Un5p4hK1ggfUFgxp/EA9JvpjCPEJUv+SroUTnrnmx6SxCL7NUQAP9BzGl
Xc71jbkCWuOmLcl+dxkfwUga1QikxpEX7TZx3xhFBXi7Gvp5ZW1f1CurEsqF0gArp2XrPGk8Mgln
vpoBW+/w53E05N7w5yT/7b3AYn7d3DrAGOTg+O7HZUbcGIu7lRl1RGYHCGaCDYrfW5p1Kl18ynpf
SEVw91QMMsMXI32EMXK3Kvw6cy9bGt9jarFC7rH7ikgg71OeXpj9uQFtVRcrOWSdT7n2HnkzudPa
Xrf/jZb0Q6pg9YJ0bXrs2IGS32/iZ+SxThJdW6XY1QB/qRqMPcpkSOcsTYgudThCTbFeOychhUgU
pr/5Io91Z47MNr/r+8FGF3goReG71RiVQpgvMC+nIUZFHe2/3XbiFSAPFPj3NbD0SkSa57oYTT5m
eNjI2jJoe7Vq02NmgU0q5UosYPwwtoLfWoo7/GLiMEbRkbSmblYhvTiUlMjG3mBAVTu233zPEnUJ
QNwiIhFgeKoRCMW/qLBAScEAfZRz3mjbLGOOJtL32F0hcTgq2qQXBf2BDLUsJFjVieTvMVniiQXF
v3uyVrbVemxJ4p8raYlyf9/RGmm/wsL9Acn8hnbW+/ItIRldU5tmB9JUQ3m0kCo1gULKoS7vEbJQ
1zlSJtK38VUT4ljlNySIx+66GjRAHWYtXNFtsv12Ifq/hxywIlOFdhTUllM1JTsf8JAM4R12c/Zi
1Fd80g4PxywuQo5pxF1sNODUbaZbH5IFdr2yivufH7ehyO5Sv/HQdRw8VED9lBzuobnCcsEU3nie
iqLfgqat1ww2hhEH3F3FeAn10sWne9KgQT2T9oKX5qEEYXv7ExAL0tymsCW1OD/3OCeIUxUA/uGL
YqBNeFqOEIzIVugEEb8Cj8WwV8xTSpF1nFzEWXVzrNGDgiTF16BTZIYopKtvDZfjD1uVuG7s8gcN
ihtI9u3BSp9YVvK7UIAreCEmh1+7aEDLhrjy3vDNx4BFDK0loPh9SudbK3UF/9Xx58/G6ZIGWu8I
pGQjY+iMsPi2S1EwtnXFK18kOYcSl3pPHYPH8PA7KhzA4P4NHFwcv2JVsy1bWvSyB390OGOy0Hz/
4sQkJ/eR2N+DB3b1oesuYS0wN5Z6KZO8roAQ38AVdeLZ9fSyEDAtjXD5HRtr8YOR63QeE8npgb3A
ttaPoLtfHgf4g9t1DYazTjRHXG8XZlrjF2jR5eBB/l5qBYMNiYOkB6dgkbmwEoxeS29wpv3pi54a
kTXz+qV9cNWItCmReZUU7LVyjRIXzq/nYM5Qrdig9WWw/YRy6iC6KqAhqebQjsw5QzO92aIf4whR
OQC4IR+KfFqJDtVBgMJa51kvT7yKkA2hnVNSHyjnQEkb7MnH0nfoO5unjzmKpQZ/7E8wv/jD75b+
WQf4YrFwItO+uueqMtJfm/HSYXshJCs45Dg0I5YEMHTglp3yycZ/6xMZ9/vhBAYLs6FOr1wszVEw
Ea9OsuUwIxExtlmW/Uyg2VkeQkm5V8AKCONQjX4S+invvVbitU+jnKB4I93Efn4w70FUYyAnxrLI
tuayZy6fhZW8zqLfvK+6GmnY+Q+EEQHPKhG4+fyHGiZIy7jEGVdblUoG4kgnHcLda7Bik7pGRxYk
bpjmVmKMwI89ySlfXKlTBfmJT8dSnVk6fHNLet1910FGe+N8FUONtbz2iAb6dz/gC01DqbTMPXEM
kAK9GckHHuEw7rVz81GFCwHbno6hlWfNerP9pDCoWfCbWDgQ3JhCvMWLyrdsi0z2OrId28+jUZ7G
PdAvHy5k3jYQHcueAS15Kyy9HhQ3TSa73WBAZ4t7K/AqB4sqxVgma5k2wah1knKOk23WPAspGzJv
qmEYUKC9tBtOZcNmvVBR2whvm+cuStuiMsZoYoG1syGwhO6vqXCiJ6NTZ2mps1lWIv6IaNXTzIe/
ddwZ3esS2Jhfj24ZxQUhkfJNwkQbtZdaLuAj8VxCXfe0+GZJCO6DDQ4uisxyGbt1e1bVH/VV8/Db
SiDgS+8UeJaOtCv/RUpwguZr6jyLRAij7K9ZP2OM8BkGH9yg3CoCLsQtcanySkKLUOxtgzVmfajb
ov1u99df5I3osnM1Hz74/wAzs9C8/nZr0DCmyYn+4ieYKRt0pq29IIV3/oREV7+qX4ye0kS0zEWv
REUjhM0FniQFRyLy6Wtj0yrUxIVM/P/7Z+jCmIYK3WbIPjAqojoAP1eeEAD+4hSqqWfSaPnv0DDB
NT3HcZR6e1xuCuzKUYjkwlq+DHhs5gj4wrQN7kwDNusqII4cebyqy71oluoEkBw2AbCeScXHEd5j
3vvbSbZMwJA6xLAtU5meB7K2IndrlSuFWt5/KGLO9nbbxP1dDBR5lkCk/PNmfaMlpKs8/qDrTCHZ
wrcdPieXTj7B4OYnkKIVHx0s62dscQMVJQWncGZ1LazYgXZeVRWCPHqoH+dAZpxhbiu7VTaefwej
I2i1DwTuS5OPTPd9NCFW5VGA/slhdlfpEkuMO1jd/yKzzfeRXrSHy25uvr1bhBXCVRJ6zS5q6Cgy
BmFIFmSz9sXg6JT/HcAwUYvvQpMjmljZCN45yLwVT+AdqIxfNn+MJH4B3FVUDn7/+dx2OowJg+RF
rigyzqNXarjkdzBt5pQRrvwkfA3m9ZG/xQ8tVIe/dBCGVtwjbvAmvajm9XPsAJSrR2xvn73aJS3e
MM9k73k7SzxQLCQSMAEdNI92gqr7r3pbDtaXJmvofq3uKbrhQYgHG93zWXNqFRvx4v1d2Ij0eyYZ
n5WEQBQnnjGG7xXOk1Wke0IcEZkRAMOp4VE8dinJbcNq1NHspRYhW9bOgn5+H2Xf4zzOHfpv2xCG
6nj7e4di+O2BcFGTyryrBtE1D6Fy0ChrX/2IwbTctSNhM61gPcnMw50US+OLXPZ5vVzECB7H0hDC
rz68tw8L9JVg02CQCJlRaOJVoc4mC6e9MswWvnVqNw8G8Df5Ok2SQFVZ0nxJUgEzblIDIh47Zmk3
W97YdZ3gd4y3FrnTilIcgxhnLWkrb7z9csthBDxugcrUQua/+I6lcV4pq6LxyzWOCGP3TDu3y1uB
GPSQ5ad43Ay6pP/bVBcfQZ2xp6ZH7l01hvaMHkD5VFC21A9IB6KI/d41sHygANjyqLca8W8dg/PX
nurGOPWtW4Sp5PGpNqzPWiBQmjyBkOVbmKFNKbSkDC+Fs3ihkfyUZjEfyPMKfCF0n5rZzRrpXitT
qyET0abtBjlT3Dego7MjvHxzX2tiCIg1itKnnZPzVcPd7lH0N8asCYI9GKrA/z96WhEmmUDeH3AQ
Kkn+AJYmStlgq1Ns3wp4dabNRSpb1ivo5Yd+oNDNFI2MObK5XcikUjR/iEmeMU8Bmiy5K8ajx3Qa
mix/VZcdIcCA21njHw42NUVYtKrWo0w6HBE9RRebwujp+7ONQ5cHlAHxkeWf4zEd/Xhbe/kLZuL4
2xNe+kOCZWxE9nCVZse5j+sI4KxQIuGNvQpShAZ8hY1Ya8OvCJTM8SdV8vZkW271DJ/7Ck3pjQYo
fjI9g+juk5lf0FQbRCiNZNrqsMJ+kIbuo7yJjQjNfj6RphbJEfM5R4DtnQ0P9raFXosDoiS+uCv8
CDI3dVK3RW6f+I1cjcGVYQ8Ew0zfSn/OsU3ht8VpMzDy3ZYq7KqxWjKhw9RJ5rxQf3LflWg37NKu
T8DW7OZzv4pPFIUQ8Kugbrglh9bJodVe0XlaZLEPYTbCEmFLbk/hHlLC/hGRwfc8JlEWCiSbDrdq
96szkELKkZafQq5qUP8OA4IPVEOmM59sZbC4yTwal26TelVOZ8NFPLfF3Yjls30yjdufgeeg9BFN
Z0mQzU9II7jLMacG615G51ZCYCEWYLVCGak15gvM++NXq3xc/b5MTGKp/fGKJ3nG7K7OyDL82oAK
TKtj4hmvYUA9EYLfoMI0qyAN4QiOX/jmWWY4OgkZ07abFi0zTkJTKsTM0AzDQOLe953BBiw7aEYz
Xj8wyHNqQPxOyXAY/ErveltBDTBv4wI09uLcEqJDpzENfZucsU8Gs7jaADMz4G7JTlCyY7wbnbQS
EpfjDWE2jbw1XF8NrmzniX/IvyCNi2wMVbVJBKJvrabhwZg8JjX8PwHHVC6Q4XXFYh5SuAfNVysn
kaesuXFLcPXN+ROb65fKDy8bjo/Q1M5e4afKEwsN+tNQh487qk1oOaxbzeDHhgrTTlfMQ1uoB3SW
n6B1cFYqYsZKHg6uFaXt0JBiCssD9gCkbJqoGOHr2YsdxgSrv5KpnXvvMMtQXf73XuTmgeHlzguU
rywUvVlOCLzrYSx0pN/O+Raf+SeWCo+Kns+DTnHDRXS2lVh8hEW8t/0nFCJBRBJVG62sZtJXet3t
D2TKurKCzAmjW4ohnp79mBhc3np9FxYuuEqaNynlCL/swPDlbkN+aLdW+VbGNY2QVklL80gfTDY/
163aLSjG7wh3pt/kOK0dQuOU32Zj/yi5pDHb4attrWKb12LKdn1X4VB79WmER3nP0gpicY/zDKSe
w95uettaq93x45ZLQyaVccJKbpJGW8oZfjinCh+i0UN9YfUXzEPoeb8URad2pW7mQ8RyePETMANN
ZQDK/KJgR7ClbIgHCB5nyoq37CHmt0u9J5fytDes6Mtwmo4ddOjCdi2/aHUmNsI39Z0iOFEHglwY
LNN0Bxz/9HHwFZn7s1IzPd928AfBPVKq2fdy6XZPcqdV8keeXBKiDcLTvGDGgoJ6Kc+1J7q09j2D
uVHArz2blKruc76e30UonABDqByglzOgF+ZYwwfP/QyS7MWjtlhoQG2qjpB+KsY6uQaufHq0xG8l
A3dLZ0SlypNUN/50VbRgK+Y2In92DQYGCcMbLSubG3k47poan7dZlSzocIMx8C2ZTMQiyZIjelEd
h/gIH4SywwLTwSw8Wv+bpfHONTgp9iyu4O4ce0d8hc12kqwBcbQiuAyrdg6OWV7NZLsmU436GC8H
fXcpKta4Kw/3kKs6QyTaGQmI8QpkXl9f0L+3Yph3B7Q7DqZbvASyL2el9d7R9QkFCE1Z7jH1AoIA
11a+6l1rjz+7KQJSpyCQURVUHZFQK8OSRaCofK5oQ1vimDlMlnNUKIqmCdACNW68uUoN6YOLJPud
wNMFFa+bxE4h+F457Y7Q31m8mN8+2R+2o9be9cAW5GJsW5qi527U1JrUTM1dZaVDDadFu4T+EGVI
sm4PW3J0IpiQ1+v1f+Zlr7nplT9+iAAE5pzy1jW4fp/bww1TC60eet+fPUlmmCwgTpVLcy2Fkiwy
c+f5r07rCvEeZ+JS26LZX9ueaMqob6SbV4o46SgckVTpWIlzQLvIXUi+l+CY7eJT+64pNOTyWt8i
vgTPmQa8Wsrd8D8G14aLsFKh3GdZ74ZvohBZ8VHn6ms/+ghcDDjviheOBxY9/TL6sf/Mq3YFlVE1
BqbkJSAIvEjOVuaWoGMq0/AIMyjsWZQOawTSUrFmafFyjTqBcneHW1NI+rVOOcD6igqrxwVawNDk
vAIlEA8HXJU5URMi/vQXwLtNA/2XQNmFwB2O3NR2DdJomG+8Nm2Yd0lmBj860Adif6pnBlpuo4rx
JLzYwVcyxJLLET/H/Ch495aSdMWEbP0SAjE3NdUwDxrYZMDKkU5ErUtaKw1/MJvMLzYj4NcOq7Mb
cpO7oCgbXaUC3dkKbP3GWhcpsUunj7Pu7U/Px949tywBaJzaqEUjbV+vkjIxvbEILSxnIuNccl8/
xZsHn6z/pUSO5WdUO0yyNUIc/A4YMkVESqEYRSOcgO26TJm6m4eEiwKqTcYj0nlfN/PXWGGso/E9
KDaNclPPDiW/CKZzYtUPJv8oER8lXsngBDMIc5k7Y+EmoInwX8w2mzjaTUYls8HYhiaLHWcf4ynO
ZaLBo4Ub7R6/bE/DJWGbsGvmFzZUXk3t/a8It+uQTeOLOpOHkOq0OuR+3BjgZ0qDDQgabdprXA0W
PT5TqTj1WPirB56VD3hPy4PtCVf69EDJaxXVudJeiwDmntyI9jeZyPyP6DHJy/TvPCR0M8Yg4hLY
Orv93suBNPg2yD9yTpIL8E/Wzj8hzMO+b/611wsy44Rew87FGyN8sCiuKQ/V0QRyt2CtYuT/qkUT
hZXQYNS46Sa99D0u2tzZ4TYltMdhie7UZBMuU8wyMjNNKoIW61/1v8yWj3K/fLZ5pecXYW3uUq/g
QJwqOqRjqsL39WN20A9nFA8knVgOmIJ99EeorNpM3GrFrrZ+hM7GS3hGNKnKv1TINdnLnTZXXBRI
lfeFderXq44sAYgjRzZ1PVADFBj7Zb5g6RLg3q/+2j15mPTKmy46O4SxhywlsPYz3t1nB4vCuZOd
SzE9CODDvor7PDK3+tLN0g7sTJvUtmv3eS/cQKVXP/C5fedXKPfArAbR4+REdp6EBx6GpAYmOY3n
d4sJvirEXLfpEudo7LmrmRQ2JBFgfoARFTQrMchpOpkG+YbfKKx5bBn2kfLF9Uv3vSJj0KZtOLi3
KnT5xpba6zEcMSddKwS+gyk9NIXUNqr/ObPoqqggsWzM8cS28C6xLpSP/yoixZ2p1hotdvIetLOZ
9tiw44LKmt3sr+NRLsREtnyXJniLbUD7UdEiQLu5SvH0oyu7WogpdT+LxM1HOaFlz27+clJGmbj+
e/QGODF9Iwx4ZSvQ7GgJGt1YFi5thmUnNOj5D1zwV9EoEFgGTzk5Ze3cNjat73Zvj+HeJWSbAH1V
5P7HUsaqO6xhHvgr4tv+IFa/RIzujdCBzn+3uYdpbgtzuYqq//zM5NnVktY6rHKOG1D7GisVmtu2
8LAVuN4AphEn69vNQyUVbvGPcGOre532T2qvmdv0EcUWO7bsowIQ8UHxhcBU6lWXnVDnG6EqdSEP
mot/U5jGGsiOntWwN/uePgbyF1aLP5Pt8QUk72P6QziD2TQe8GMWUJfdwPe/7qqSoVaMOGYBJrKK
TKw3zXnakulM+xC9Q5KhKM15B5/XG3uoUFuYCmhSNZ/1LjI+0dZFEhV4dBvphnIO55BGRBfGX6ps
W+645ulzvmjYiss/awtR5yx1QSI3N6IECTXdwxjy8Hg/b4nwiqYPkFO45Q8LuwoTPnKyC8uYVNOi
xtwLjYWkH18hh9sGgbSBxbWpUMRnM4hWBwOcDdsnUYzFbYGzvz0/wGL80ierXJYbHRtkco0ghYSA
WyfICaNvnTUfEpbLfU3NkF2RbYm6KOjuyqKr6R27HXs0bmLUVLJ4EUbje/ncCPK2UQaQvYPb6wMP
WNchr6uituxpW4W9Syrl73+Hcy7JFH3XDcXIJ25vabYgrf4vaJqG+KsSOtZvWJu1o08Vnf399bwx
XQAm/nEJ0YdBzJO0MLo0VL4BSM2q6EfKeGbaUl/GMM2I29SherVDGq/wCimHdAdji4Arm0/DNTxm
vm/gncQf7TwWvm2w7hPPzw/jQPVIdaC/+9OdmhEKz1Ff8lO9RrEG2Vzjpd/OHryIPuuRDaGgLtU5
YfZE8cS635qcPDU0+pZRjJG4XylyIKx3Skca0lFmPnPdbeFWWZT/+or3K8raMLGEA29j/3kRBDyT
P0krfBTvimbs1nGIpKpFlTlKJfgjGv2b0a/ct3inn59EKKKk3odu/nzQh8F/ypsp1iMptgtCKVE/
FTkcqOW9YcuqSysySKxgADjCK6wK94Ke1UoPU7zgVmbuusTVvl6CkSMhqqkiUoaMnKgT+9cBD1JQ
ffpObpSzZztUF0jvsLsGHxcNJ2i6HTJVZGNuZ9MNr1O2+NM5HX+/j+qUwCsuJaR057MSvDypQ7RY
Ngcgmy0qPeAVpVWJl1QwnHG9MmZS7eTHCY8LkL4nQjhYDbC/RTNzIx+x8G4mRbO/trO/HBIBnmZv
e2W5YiRdMMqJJMfC0rublzDuGB10Z9tIk0WmPkhcWY8ZWirJDX/dXVJeSzBtUtObURf3eItgD8Ad
GnVUScISNcKiv2hRdVQtAF/aqqHfvyUW2Eg73oq8O4A934dSBUEP+L687J3dzcghg4sjufj4rnya
5ifUCxkPL2CY4nrqjRV/tgsnhw2ZS/rqytTMpO5dOrWRJjd9GicHX5t3rVh+NL3YRo9Q2LbQ8hPU
+F3wb2eDF+iFCn/VDTGWDtOFthXEkbhw9w9XDRHh8dsydZG2hnMCkwYtRarEHvCUBxOKCCs34Ytf
X6XShdcXzORv9scWl0EH29wI6xQ3Hl//Qoekx2LqoW7M2R8ZjRwOMdyat20ncghb6kvOehQTpKzZ
+83u/hWWib/vqzE1fWQG0y/rguNsJ8VYSmCabcmWpRU/kZNpCFuAFrgLxgK69BBx4XtS0nQAusAq
um15CZmObaKecLvQS76hAdlZetdDid8pi+tUkeCxLTJF65Oe7No21Pigy5zIAjwOgc5BPh9jWRc6
Wagd/jDyc3ue/+FDiI0xsEWjP9jH5oc44XzzinXREZKnfavuN7fkcsZSKS1J0ZDHjl5umpLfrj2X
fqeJkl/ypZ2WSeHxOrklDGcFrCtn1qZeTwOrvqJSQWLIyR2qbwT9+8M70Uo3kE8P4UgEA55sqIvz
A3OJPjymin/HgxbEsaeyFOTdx1cJl+CwktVY1uvxhevILYhrMtiFa5klfxJjm+ldEVa3xaypaKQT
308c6wmuVdisHIwUGqey948Am5Oal9Npb3LpO86/n+aAqF4Mxm9Dc+YkXkHlTuj4lrY55GOuuR24
XN9JLuZQTJ+ATAfM3VLfrVnkFpsF2Gg8BJsPgVtzY7xTn/h2qYVCCIdQ06mvW+YqEi7PzOEQ5mqu
V2V5sB+3v0hanI0PGLWZMiuauB6MmH1ttfFxFwVv1T+m66XPtwXT+iTFuJ2xUP9pekhptpDpnUoh
qIy9WxHN3znk0ZB51/Yznfox9mHyxfrTz6CDPpIEtvY7mQHTaALyjv4FvVix1rtfUN7b8x2xsQfR
CBrjU8JwLHHWgGX3hgp1XdhZZUEHU3L6K87VpZn3A2lz5twQ6KJjWur3IOENvYxph6qtJyKx2bcK
OuzeT4WudMtXJnwtfkjcOeJmtrB0vdZMyGsZUjcuha2fYS74juB/P5nA/+PNTkR7l0q4t92ELwkc
v6WLYXI8fuXOeeoAKooxmnnlCNeSkk3UhR4EIi7Yu1TWHiqJsnzghLtdpI3FZTHPVpgOyKft+v/u
EjOKqeNncqQQwNKRNKTJPcI+J9nRwxlL9TeXYMEPPj1NFGDMSESuwP4VnrRSTF49pB/qmRRpKV5z
R7bIWbfQOBX12q/aCLvk/XvBWw8mk050pJtYgdQ9dbRDV6NwHIYDUL8vXaBqD2XzXH5qmN005XuT
uy73K366Ha1w2OQxc66/vroWkJRutAmMrkcELQhoX6GZlGZujM/lDCGiBjrwCibv7RR7whrcaLYA
QJdKNLGH70ujTAELHJKCyp63iTEqMWNqJxmgUjCqoixPuQ8PAn1OkkR6iwxf8cHW9yh+bUC/jtvS
2+7cqujZdakVIRM6SEDPkMuAUW91ujQsR9sBN/XvR+KL0gVWwW4EdSSG5hF19oNpElMmrl6D2Fp9
HmoUPslLoybnBpM77KGo8rAWMFIbKqaNf7lGzs4cKu9PrhY32qhbQc9OMpH4/AJhYbO76nMwbm2j
fO+o5SGxrcCyTnUhYkoGWvBFnRLZwDK/i7D1YeOErdJ6ARsEFAjcZR5R/Z8SJhiIUELEGQzRykRt
mXZL6p5Y9EeXDzttpQszTGZ9bhIFulpvO75Qaw2cFkUGDQTYjw5e2/9ftQ+yENTV21sxSNzA9UHS
Lo7hCvb5G5hcvYTuuXvWROHU336H/41wOkmDmC1IKjeR34UqEWoLZsA48uDIXl4rqX24y+Cf6mTf
eKTrsLKKbiUGcfnrrzM/StKi58txQvQfsPiXGf9WaMqjZkF1pk0W5Um7TGT7l5lE9yXNOSsWmKEi
GF7tlE1IW6oOZCNUy0wrOY/gQTqZrUfRX4CO9fLaN0RCWvvHELcw66gzcDr4y0PxpE073E4RTttv
Bape3DEl3F/Ot3SUn/4dlbmJ+QqKolY+kfU4fcMMJ8SV1N6hROUJvCAZszvy952gO+6vOak0Vy5M
WOtEQLwfSSSVJIejnksmJ1HXqnyjTOJu7izkJW62U8FrnHqdqf9rVgEoDxm1fSERw3Ba0DQ0Khn7
Kq4ig2fKtGr1Se39mwQbfgyL675f1oN+Cp8Nlnt/LEbGLYcpkaWAWnGiDBUWFsOVdZJYuU6QkyvA
mtwFACl2dWchHRKArw/K+uE2egsSS+j0MIOQXm8z3Fy7oJnonz49xnomDTVeAy68OlZ/BRPKO0ZM
5UG0NBrf+OzRsI/DpFcLacgJZoB1k25CWZbfrUSkXHoiturWsbPIC4zy5gMdhUdTNbjiYkHhlG1W
WG5fshb/gjtM02APGxILuID4pTvTp2Y5Pvx+LzSgN0AVVtveeSsowvBGXr7chg74C0tS4mhGsuK8
lnOGZPUosZKKkZOECEq5ObakMjOYF1yWK7X9+qpkPto4LRl9dyU+iIDEWHsMVXV1BTpLfeHSbD0B
HbMx35+Rfs7PB7zhpcmCQ7JuZOzEc38bgxfjkcYCamTfY53QD/omZCtmkJvQZNnUuboKIX2dmA6W
wJ4xuOHsvxxdwUwQ2GI0JSU5QWLo4u1tExVoDiqOX7TIW7Px/grf56lRX7Vf1LiQ7xy8Akgd2w1r
rFAq/TNXeMlEMKxmRdMpkh3SzD6HSIDewE3MD3InP4eonFIfI01/NRAqTYJs5hnyhAaUTsLq4wr2
eP3x0pYjgILc4HAgs0mOTvYrOwSGfIldEs7fT9l/l4PE8X+WvKL2P6q3N5vARV1pU21kxlsdvzHL
ZiET9rEBqqL/qg62Zi6KJpT5bAB+BOG9UFnIFmkB17ljgGhus4fS9TTkeKXcDJWipHETgvUFLHyq
ruagRnEnRyZ+Sb5ON99noTd8Gfhrk+zG86FZpSlx03wL8n05vwXM2A5HVio448ABNABLf79gXjPy
W4OsD07dfyt5FmY040pWBg5+7PTLLPqKmxtZ2J5R/LsEoKnjx5T5PzOUOJ3UaBrlPW3+daWNp+4t
3833AwAMATHFyPh2eN9DGVfuhLqqoaVqNUz30lGvdCbhZ/r2q/KlWNOI40kvx/kDFp1jSR66sWmU
ZvKC3ZDRAm7HvAsnyckTJq5W7VFD28YqQnfvNeQQzV1AuX45AVzvRwWFAgLbPE9MC6L/RGIbX8Xs
AwqbF4Tr9fQFVSB+JzW8RTONXHwyawZhvEeHXnbpyaIBml0+yNK5kSibySiJWfr0XZmprXq0biaO
K11bCL+udy+Tl2NgIVrhLMngQCrF7I6bIrcUzw1WHiY9IGckeYPT5w0yjs9f9GYujQZGBeyuxZtl
T9mqUI6JK8hggewezVTgalON0iSDeV90Jyvcb11mgwmzWJW1zXh7tXi42QK7wnx92U9go6J8YxfT
CT5F6MLmLFOqsNtkGiUDKTbKtYz/ObLdTMi6xAFEYK3kwFYtfXLvtC4y9WgHjBXlsqbSjtTOcylr
ZuuBGNXcQl5meKEJVKxtAg/9QyLSQpzHtIm6tuGRCpUMuBsSMMC0CL+LjwwjsBsiJ15Crrms8N+z
1+ai3SZkSckLZLoMdMO9c9+Vz7UmUh/+iTnyfg27wdPM+FMLsyd3Ya8ZTi/4D3mGPr6WmYaXAYST
qB/qhOATcXtcquUc71djl2GcbN9FHXGbc8HYapeXdNpNBsuS/B0WvOvOW9uwg/8C6X42JbZhkbrr
Y+3oUnihWzkyaRoh+d1ppTCAa70An7yTn+q8YMeqiHk37a6AgnS6bUMXD/VGzdlnS6uhCp1lKeJi
cf5c9rp4z4RDBk4Cbro0Z2phmAeVfXQMVuAW7mN3lNMKal8KekhSMJOhmeAn7u3Q5li2oalJwO3W
rPaVA2StRV9wbLnkIic9rXz862zkkoel8Bj53g1lg/fj3VmgCSztDftPQJqUnok4i9/hZS0XOwc7
jbuKKK2TQpe88RzQtV1GxD1Odlyd2yjxei/C9AtyTIXp1bP4LvIaOLrInssO1CHD4OfNC8QgPqq4
Vc+t2sRCI8D5jrhGgQKCI43kNKJ0a+EQmxyjov2gbAthnfaZa5WiKNkUEqnqjAEegUn9T+DuTsvq
u/Fgzo9TInr/nhvKZbLWvBzfvbFM0x1clY7nJYTCvR1JckPjARIEeniRbnihuFv+VAvNfddLCqdV
+O4Wuic4ewKOmprsOgVxz9ng/lQW12QeOYuDRN+/WOi0bhMEuIPkribEfdfSpXjaQuOq7lcAq1gY
ADc/xLxx/aGJjuGe6eayGLN39pDN/AoClOjs6rnkIzLZO787NLAlOyps+FZSuAYjr1S181Dnnsxy
MhFJxy4i/pD5eX3Y79imHlBT3YulaI6SwVoUAxyZYVq7M6ByhZOMq+QzxxsfStFUZQEMdf8VOUGe
o6GVomb81QLhM4cJPMBxfdGpeeyOyFuVySBAFu4Kn1o6dbKHIYLZche61D057OhAkrZFoPqDqYQp
LHzH9UQ7KOZjoZlo+RYbsXA5XR/U37y6CRi/LuJj+poLbxBKfRR3W2mYrtMO0I8BZh6yfDyr1ot7
/t4tWsmxNbiij5i3ahDtLbQaq0jkRSPJrfH/CC+jvJXuCWF2N1LcdWaEhtAf687CX5J13L09Nekk
xgmMAG2d+6cmwQCNDSnAXb29Fj9rdWQFeFNVIBbvOE07s4fPoJy963b5PXUdrkhFAy7JTz3piG8V
7F0cUJr7HtRfSczxJDtOmuk5rfeawgLim18ut4RocQ3XwSLc6sR4MRoftcOIKybtPddUvlPtod/M
KAYh2ta1kjtMjE12bspmzR0QVp+chh4/bOJGaF1ZIrVzN5f/+vCSds+DSxI9Z6kPsOEueWjexkYp
Dh3Dgf34osxYfpX5YG7mcZlRx/ubD2VlU/giyP+nbob29iZ2OlA7OSqxiFXvCc0GH/aY9uGths4Y
29OIwIY9eYa4TkKrRAM8FypbS7XGvZAboSK78T9fQYWaEz6DXhKoyysVCYbIKmSeZOf4jYFQMKEy
bBd6BoTeIZEJJ5qm1mXDaZJAdIovCTSx/5NYPb4xhslrObnXLmhcaZuMatPPaZUslL/5AUM9pB2y
aMmqiDbC578w+Z1zvCe0B2bDVvY9ETg6aFdXWFG0fIIqEpIJC6TCJMApTxxMgdDiVoInO0X50O/1
vAQizO8kPL/2H/zBq0MBMHyfEEjp9jYqTgCHmFYWknGyppiF8DP44DCGk1zZOpEFP58i3+F36Xic
364THmYWnF5ys/Fd7WJF9Z+65297pVd64leOrWX0MUGc3pwaSvhluK8Fr8d5KHR7Kua85iTspGHd
EUaJD3p5FK2sHEWWdNlltV1w76SMc7bEtNAA0pTQqqwom7Css29sizw7hRd0nPs9CPOZidSpsc3A
hMVuwIeRrV477Wk5hPCltyomDCVm8QvJslSabQRoB1JExA7CGr198HPBWwwLWaEUBQa+RFR1mQap
hMk59VCTq6J3+uFfDcF1PoU2XkE79nNcqCDsJmHl67gamkY/FFNECe1ux1fC9nENQpl2536fjYFa
K6jbXpHLgbXRb5Kly0xH51sWmId6F8sJslr2trWjxCq46IL86e6qnHVqgmxOPKpwu6kVvqey+2y0
FYQDF5kW+pAp4SOyOHIAWxKp3pUICm8lwwEBbhJX50jpDuLk8Jj5Db+ZnV7n7uZmvY3MX5c4H8+p
PnWMH2QBCWMExMeN1JmuDastuY0f2rZNXlj57eFVIiqLkaWe2JW+MMiOpPBYL8dcYxkHry+y7xVL
cC7+m63I4WdXN8wNiextd88HnwJO0zhBznKJ0OqZyeqT6h5cEHQ+/Dtx4BoAIimLrtGg7ccWY7qA
+dLZiyG/NxZrZOwOfvTCJdviOueXm+DMv6hR3nrS3uhWb5c8Q8WNHqctA2QuSc24eRC5E2xztdPe
8Ve0bg8QUtQwDXx9tMLdM6fiLfAk1vDWl2g+xhgfTB1uY+jJgkoikFylg8X+5z4mZE5NfoSGeP0y
WBos0pfpi1j6dzHCnrQQ3Snddnxim5NjAsqAqVRaOykgRilDfw7H3aKkl/Vhny+p4ZZDnb3L2z8g
REB7YRGPP06lto3/iGbo5gOHApuhQKncO6CpA8rUYoj0uVNLRf7O6DzteLrdui3EyFec+n3auYEQ
3nBqOnArbv+6fr8+yj3h5dff5CLaIrW3R7MVHUVCLL7x+EkrEugP82AaqYCjF+cXM2TolWzjiS/S
9cyy/35djtuhcpNvp/6+scrU4Qez/ivSLJZ1bn5IL5g127TpV+9uaHxrslWZQbhBKs1bcg72ILWL
GHlZlpU5USLGY7TEVOJ1ns3ryew0usHjbI8MVHB+rZwAM8F8MrTDmOCbVbGlmZnkxXnALTnyjvvR
KH6Oepn2iZKL4jKA5TqjHdAlEC1LZjGH4HXT+OjkUgf66tZOnfEXiOWQ+fV2kC4LpPOJmj90R3L5
vowgyqr2uVvHBLn5WEq3Vie06cKxQnUwWtDe0q5QH6plqfaYw2+FL6dE2e2bdjrlVWO0OFOBnjuT
g6xPFaDGK/NE2fD8TRl9eqqf2tF1fORMmdGupgWA1mwlC2sqeMbCAR7psK6VnUj4HtPFF1FvYFLo
V2bsQN46iJNLiyDq5R4gqw6IBnnHdFqIqQGSk4WVE1XzR52GMVN6wc+nqw+h7s9PYmu0usWCvMIT
ndG08w+FoKsOZ6iLB0nslSj3VHZQBXT8622GMdIDyGR7DP6U39BoL/DWFQz+9yV7EnPKXF4+VBKt
L4/I++7Z5/tfk5/rrudj9WgI/W/SSqxc1ervk6PLyyNK/j1Y9ZA7bbXV5P4t2VOdy0IP/P37K6rK
k/2+ERzXVfYtRp1ysEvJxjh4/9tP/w09JpvmIs4MkfHopElvmv0RvJGGXlDnQr2Ofj0DHvf+59LO
P1TUIK8wurrJRHYIEsOloNcXHH1JY95t5TB/0zxOziMEHTKBSpJAPJPjaOwaG5O0VDfuFTTASyk/
uJmQPPYtj85sj2D9h1ybi3W9t0540ZWl8LMSaiEeTE0UZ1WumuO9qNY0SKAV0IM/yKoHZgZ/RubG
eaB+SLQot+dfZp3iBKm7lQaGDsQ0l1I3D/ePLSBybOacRMjGG/T8n7liaK80NTU75VEIA0ybOJ8s
QcGOexqhI23y5uVygbc37CK3/fb4+efw/4B9yP2ihCNK8VmgW+qhS9YfS7bM9Fxo9yQGGmJ0wmbi
fjmzJSv1M2L42UAeMIhrV8GhIVV3xqDNG7InDS7xbvHFXzu+D39KZnsTSYKYSu7aWiCzpffa9e9Q
2susoT2yDrGFlreYhqjahdzd+UINpV5j5EsDfq4oJD5tE7Ho0eCHeV6VBth10mVzT+i7p2owBTp2
Nt6AGJ7ODMak2u1+czudL6yfWi6g62m6PZn9h0gv93QuRmN/gtu/x4sKk/N4WXsbNc6NU3VXKd6Y
9DRdvFR55FliipqvzcPxe3/+ZyFR2UrlRCZlVCvuUE4CmJWlpL6x3hQzx7D1FjsunBXUqs37Xpx0
tDVZO1gLyobmr8jBQCdYEdguzDKG9vlGPrjA23Aya59j8qd8Juw9FJus2jNEvn+34u1y+kYgDlCf
dDOhm7wPczAdQaeGYKf5wmhkzXc42tIx9PzzrN9UwJVmvREjDUBqk7HrOi9it5/hfHB3/U7qnFgs
uRceJ2nPhJFlPI3B1YTPGtE+bFNTsstjsb1mpyoffVBqkYIDUt2Ihx5/3rEnRxyfujtLtKh/XIYA
0i+NjomqewtSR+2V3jKwEBCoSLgCd5ugdgwI40aJe1C+IHjiv4B4KdwqDnh76zkuS5IZG6o57LnM
Ps8hi/GJMc76MAfdFf+O5PSGzy69dqllY3wSF4mspKVBudm+1sc1StKwVOiVlpR/adkP5JELhh8z
JQKhlzPWRhzCT+HJ/tGMBAED7XXwe/1WHu6vt9bkMwcFxi3pEb8dgaJe4dwirv+UklpizYsXhy2K
7O+WgGoMNs/Z0zoFxXwZsTY5EJeVRjpjrYIdhjU+Yhs7iBAVGZ9NGdKklHyfaNcxcH/xqIVhYvzq
jnbxoZ9poRzMk/g1tbnB0GXgueyxvkVqTXevuTg/5FpYw0qv7uWD8G49s0SzmYnWijBujCtHAI3E
/laXyNeoBDYJ/sRcAurDXOd4KkYTq1utFw6wJLeSeBVsSSPQtmHiZ0wVhF3MTSDAsoUM6hVy17Ja
QVjlTMjHt1undYLIs+L8zruaqgT8RLYfwxTni7PdOzr6gm48hnj/ooG6xEBHqd89MV4I3rff6EmE
tOSIxKRkMXPLO/LBF4CVYyMo16+h7B5s+nHanYg6McpkMZvQ7aF4fMp58zC4kcARIShsuenHjyc7
w9br8N669/MyV+0hA1HRmnt2wW9N9AKEv6WCMl1refmRAtjBRK5Mf8YknhNr0iZPJ5ujnLomPYuT
tP6iJw65MEzEufniO/+RvAiyOo8Ht6I7sdvTiEo2eyxR3sdybyFnPApA3vr4Wei7qA7Et9mSIP5j
8thIe/t28gTJLiZuR0VacbLjZCyZMVTWN33BXRzKOnCH88OuoyzsWAPrl9hHAonZeevW10rjPrYe
+2DfY12SXJLNwhHHX5YWTUPCidPiyMXNM5AybsQdt3b/rOAaWddWiuVqrzPHN3pqO+hMaQ+mHUCe
E0NIroLrUJgewmNHNMpy11AG91FTaEe2DRDl16JRgl1Fiy84Q3VL3mP9UcGGzq1LqXWMRTqd4iWv
cPp3wwzmKReOpvaw9BvVL7MTkR7jqXAm7KcLSeWPkVG0BQqyrjufHKGcugUzb4Z0AnVT/on/Bshg
dPI0tnhQisxM4lQP8Yx5Fv5T6H0eWDZ5gZDUdpyJZPnKgh0n2O6dPVNGYLgoNq0KKwmzmfB4zW55
GfDBH8VFaXJg9Ru7V/EOgkQRovqz/A8K5bsxDXkmGuyDtWYKtWES176e3bi1ImxXVwJUgvvG4+r7
xShYXRc8+3iYVawu6QbxAiQFP3DCTdRrnLgZ6D6EW13KtWwQBfvyGFLqTEFOaZrjNV/yrb0zrW70
PZGurZjBVGgRZcMtPvhZJAkhukpZ+BsKvYgHmJ1SIq9pK+zWJKCne+TMmCrtagatP/eVv2D6IrqX
Rn1EkLcS/TdnhZM1+8KQstbFOAOEgvNq0lbA2BTpvjEBaz7uBpRWgjssYR2qTGThtG2pU1Smib+d
BFcRB1usUD7L6sTE2RRpz1cRrqeqpQ/5e96QoNTBFLU0kRSfRBrAQRcU/bwiCDr6ggYsX1KD4PZX
NcRJrGZBpHjmiwcJOGW5p2hcznvyD27g2AxTshlEHLF6hEVwoKy6p40FYHTZqCHA8AWKU3AcZm6l
HlxfcEPC+CHzKPxHaCHR2Gi9LvNNIP860z6XX8XJCARUSL9wUOz7fxUF3qldgBid7sg0ucjsgW3v
r7rmi9/rV5RfhDVER9sXYYVSJMHqBgmX9Npb2MLAU0X5tpOXQ4tsD5rhBHMLoNL7Mp6/yfzVHQ1z
N0LGwXHQEAIJ4yzk9r2tyWDCwRcBqGc2wcow9wsMg4Q73Bk4fb7qYgtBsqfjjFuWS+xLGcTHj27R
Sge9G0vmhwnKxuzGcOEPHazKA5s+aaBG41H0Zl9HX0vbU14KqSO5oAdz/jnpQHahTSdwQjeeYhe/
T6VeHCtCOLPkuyKnOdOQQx38OZNHtkEiltIVJHnx5p4JnVTm5NcRfgUFdQKLb1Ozj4k4uNkn/F1r
MJAncJRi9csXvQg0kiIFgvIym++AVEBwaFtNSPYLi+t9Ry2sbhb4ylJ2zGiwuRoQu32CWB+HTqim
3kvoirBjm8wwRXH2LNreFE4EfvS9VLd3a37hibWle1y/kRR/rccyKdC+gkjkhG4H5lKb1WHWXhqE
91gixF1CYYTIrWRfvrpOYHXOswzJA73qsINVI7S3tNDNoJCpXJPuhAPiYGsYXx+ooFKIJOziNis6
JFeGz6lqo7euEtZbNrYf67UhlMKG9FmqH1kWNiqNNTIUsNij2NQJxDoYduT86oNR3UB7CjbJis1s
/ra8U3Vt4MJwSBy1UWgHEjB0g1CtlDirzBfpjHy6ylI9Q+hsHj8FPY7hoGIQYATMQQ47F67T8VQ5
d4Bzsb5r/GDHlWykqCmK6LFHMsyB+5LJAVeuF6Ql6oQWnVGOHpZTs6gcL9QcilhT8C+cVC4r8kze
lR3a0igJMzdTfGdyqRbpg7T80o2c6cktJUUAiEsMyi0w2N2wExDtKPA2W8Ziqp1XP3UufywOHtuV
dNdzYC+5AfJYeMI8u5CzkP50d9yNuAGMsD2ym798atnCs4tUZc3hKpEoDz56m2eLT4d/tsrZyd7E
4Bijxmy9VLHQicUqyz0ifBqyuS5yy6aJ95k9jkqzFhn0ecZ8UJJUhW4DHZlyux/hfTHzFr9A9ppm
6pclulbJSXoWnS2QvFnWZ27+UfiXTpPsj3dDZQ2AwKJ7ccyb06chjXCtw//vVr7sX1pCszuJ6b9O
49084z2oFVuzKHKuEmEmO30hMfh/nKpAwvz2tpfjX4GKLhCSlIg7+AnSuN7Lc+Of+O8dExD8hi0H
FMG47q7WVbVq8AlMnkc43Q5XZPXIgPp+/qMgRHfZziHG28+LCxCqZX9jIla2a/aXG2Pkkkbnyk8r
S2wx5ooNkkRC6p9/hCCRvIn/VKraQZamSTUdL0Ba9Wnx8W5LsVPpceIRo4mLPdiQPy1S53t8pmwd
iq/f0HstpGC+EQ/66CN8lTT6NfqyXsD5xg/7khrF32mo3x7tgTin6MRSDqdH931dxFQd24EFFSat
rdN7XyrECYsnpPT4wk07avD2mdZ0C/CI/QZX9wWRMnLUsITbZON5OGnYi3jbUl2m0bD1/X6XtVtX
WWCOpS/P/C3+At59VnS6Xgn7oOPUW3mtfwM/qrj8PqAyASTUFZaL4xYxr3/qWIakwYkmCLKkkXqn
llb/Wt+xg6MwKqBGaDbWi2TwzFrCYHCacTuaBrJ8JF+uOa6G7E+chtsYYWCkT/nbK5vKQYlbmlfq
SC8Z8rRSSszWcYdCyuh0UUifY1eSdZHe+ex8VOUv2Mnl+mj3NoM/fELBCsw0c/avnMrTKd3Gf75H
rhU7e5BE/nM9KeEmt0Q64anQkH12Ffc6vGK/o8k+YJ4ATciBTHXZsjgVocbRea6J7Lsu35bfMAH/
E7Zjd7+TM3x36+asbHZzO94pKnoe7kBSdeBtZ+7snbsFYuVaL/+VUpQT5Zan3/9eGGKuq4/nLAng
8YlUF+rkG4l6FkOTB/jTu3IkQsmkZSIz9mCuIGV6M7yrJYuZhyLauXzeM9X3j7WMp4OGINFctzpC
7949ZKs7i+F8cxGy/tyGEx/SoYVUTT8RvOsxqIzD0AjQhxPU6BHdICStW9kXzzM9B2bpwEQj3IK+
MwDf09nA/cRkDOeUlCngOkJ4ymezsucvtl2NRxX+0a4ofBPfdbajbkQ8wR6zj548mRDSKOrRdUgr
m3lyIlY9QYJ/z8da8v8TMbhWAG0kbHgkrEviNAobnQ5lghnDry5sTWEv/SaTKkzG1YuZSVePInMq
rcFza6tSXzRxeZq3cNOm7lK5IckwC1YF512UTPAAoiwsDaNq+DSBxeO405AJkPbfAZptsD6rDjK8
reokels74Anraa0ui4KFESU8+F34ZWXnU895IRMsU+6mskMcXG8f5PNQerbjCbirrUQkc9hsnhWk
vxcam7NpHH0qRqjHlBm4WyHjqCipHM/0ZgVLyYsQYTahbt/3VgIQBlgTG2knzqsW4TJ0eHv+eElr
fjSCY4BRKAJLwAffLoADC8iGYpdnrQb6ebvtFO+5p27FMHukXmg2PtMw59HBiwAbwOsBACxFulAF
vfGlgY58igpBZ0BbMey0Nk/6eZ9O/LQRUnVoj+Nl/oQ10/dogFu6N34rogby6eFuVqDI3ljpuuRv
a0GNXRdUjzCC1Rrtd7EvJdhuLuYL6lH1/tm7mpX2RVdqP41/p4zU51z6q/nReUll7LBjMoKgZ+/i
0n0k7vYw4fuZDAANHOJq4muwhXVNVHXZgzT2MdmkjlmMgiBmMsB4cZ4/54F4/5Fu/uvtBNrs4El9
oDofOEWjFAdmh0tHAsSDZb9M/0gHYF3zU2WtYYZms5nxpYknmzk3zR+TU+q7BMziuicqsebjHT1+
hxg36ZgxsRQ5hn8jVoUiLhYbJ1x+Nhevcqb8UgBn7o6A9GArTSiBFNzdSFaQiapaN4jrK7w67Ut1
1Hkac3LWlQiVKyNBd3WbxafjrMTecUnADQ61Er8p+dVT/RIs6yqHUXf7lFN8ylH437v8X5TdsUZw
/mfndO4lYCI1G6UR293SyH+phqktXTcZt8Qn2TBvGl95Pq0gwskVFPAGtcVKofD8EJGOBvDsRo5p
cp8HOIOs1qEjV3FxIowrZgYtI3SvKrfdTok5B2XaAe7OAga2msNRD4nDV6XVzztf3XSfnxTQggP5
41OrAxwgCfUkO6Xe1dzrI1zgnaejxfWvf86jMvZRXL5yvDV62BRF+SxoLxLJ9p6t0agixjptNX68
5vpqJdOud2I0Zs8NYUAWcEjz28dGvG/OrXI5ZUriv+IqU1VmofWOwTc+qhSEJymmvQv7ckjONuox
JHXdaKaxeaNd2KW269eGzkgNMc0zVUoqcAYO823SJmzGWVRFss5/t+NA3R+tDVuQnGY19rAnD4jN
GkA50UZtPzLZSIKzrKz8JDjehhaRkryvxBf9MRXut+wjJ7gaYd7Yt1Ie3UbT8jcLMGfi5GAfQ5eG
oLmDW8+Iclje/L/AcZ/XCxpbi98nHK4wTXgbBfK1xZSh5L9HVsdTG2BKEAJqk4wTYXvkzXVh/i6S
2ok05RGLnclOQ0jbM561Uoy3sAsW20Lwkzb1w6csJTf858SIp6wlaagt2JlA76ZnEYUgfhcu88so
ECV9JEVwnM8OS8S7FyYwQ1ssRvKBaCIGNJKNbUnudrL26FUKcvFv+fOzpqbBqY/pZfCANDYy1iJ/
QCwQ22S+plWN3nN4RJqNa7Z1ZixP+nPKKhvHb7kYt2n6lHftoPhtFeobAgpAmzQRVps7tBxS+2b/
LH8Pl2O7QQzfN27TU4soI3G4EYN/B9Ge88EzI8aQKfFrx8GqGs2vkxBWLsn+m9YHlJCF5cidqXgS
jcAQK7N0eeJKXRTfDO+oZnc3hynQNeQbEo14wiSiRKfUiIO6Zvhx/g8tseLn1Jp2L4pYOKywJvql
9Ln221ttrDhkV7Z8dRW/Yz++Yz5h5ZmTVw74gwwtwEG+jGuTprFwczTEKVhQwS0A25xAkTCfgY+G
0zBRoCz2LxBEv0p2x5lPCkUtvUFHT8fFLGn+00AdP6o0ok8JSh2DkrfUukswIGA2kzxwsEahb59l
e+S6pP3nM1jqTDfADSvlEb8va+jESzS4qjDlNF9DY7QW9YhaYd8Nkmb9adstEDG8qK/7REJ5p6ef
K6Axvxc7bbhg8ppk2BRivzpRvwD63Je5eUBQ4qMUwQhkQTAxwDMuMmRZ+ZwLcsJfK0gO2k/TdSyn
9/vso8Z+w86Q4N5dUi6PTCRSe0s52a1nl+Nc/5iLEkUn3gQIYVArO5IAUsF0N9jDTuAGx5HWTzyF
cVzvEeE/+QLj7sZaQHw5xcShaPlRNNruqihgaAQilmoYyo54bD2PwYFsMUOSzTl74EQKmYeWXukH
dJ1efovnHHTAda/MaHiNfs1sgDV3l852OWINzFnO65wHC3Iy2WgxzmhNjnlsAjiIFcdFX317vDPr
c5HwczgAuqOnWhGL8nzuKofvZ7OaQNOikM3zzTVjOtFmyLwjkBVmHti55LqWuXUH/G3CE86+uxtR
yyJMRud3774Z4jyren5XvsyhJHD51RwsQlrbChyvfStJin8/mfc+MP32KFxbjstncaIwugXrb/AL
1xzZfXl2DgdFjI217YIIp4sBe9gv0pvppo+3THNTxc3C4m31ss+Mxd0g5RU8WfvRPNmifQ7kYHli
+C19sTozYW1t006Ve4esHx9GJ2tI6lVzGAcYGdRCAmng4Wi0SSMJuk0N7GAEFDIkuZz4S5gE4oER
NqDZdjgNuLVIBohAPm+torrvWmi9uaQwExazD2xdfQ63N1/YE2okzvjvt00FxhiWWGn00/MvRTGa
uSO4d5pGPw4/TeTWU3AhonVwElHXRqcokSq/kE6g0umrv/cGAHaCeJlyMZf4dM3GikJ5QNIp0qZu
MKMwFbW5etQoFLT4YtJTc/QSIJxt1SgSTgBNBGEB2EKfdtDJOK9HAejg34tuRqrha6Um6scm/DLo
qfDj3cRdlkZmTU9UrldAgdj1wHzJg2sA9C/Dp0IxdkvBBUtiVqsPzeH8JDIaplaga0k/sHFsviox
hsQQBSFwU/VJa/2oyTZ54i1bRJ/U086ie84DlVjSYvlte4AU+0g621G04/VGdTGXsKuVdVfP5esE
xJzvoiYfQAuttGylZP2rlTi3eSb7/xjyp00IbE4JcLtJYvskA6JacI8sOsyo3GCMdfgAIaOMgDx/
OgbUfAp5JPQal5mgg88G00rVCzIMFULAm6mRyOfHZyb9c3n2GKVT6Jfj+OPZf6/rqTi/YSqPGnyp
k6CxcsFw4rMkaa3baZHsJK+S5wZjrRwDE9ktOG4rH77kBMLge9hkqbs0Sh8Tc85rIFoYIYLGFG7G
OKPnu7RuSU87Qik4stbgAcya5Tppc0D0pu68/+xZZDXkccIgCI7KUU/XGaNpBL5LPRq/9YAy7vp7
vgqAnBTGyrfp92vQC3EaFUYTKYr624Tep20idYV9drmXlfgxBn9qRx2Aqjx15OAxgQPZMmHMo6Ca
u9vVeOfnrxUR3j0jBWW/N7Iji1volvFulmeJr11YR+7vCtInRBIIjB0VKyp5l21NIpaOEiaWhZ5J
fu2+1aO1Y1GNfbMXd8+5sZxc+cMjzpSfuv1U3QzxpEWYrHYEFhwNdRC3SVcyQ9ZdLNn6EURBqfxq
JF/LmpHsi9DeQxX0mqpVdyA4RM/kKWeIUo6GDS8TosC1FbLMnv3OEsYistrFY+ZIbjNAMLEv9BVJ
aaqNY4sC5KyPL2NEN2fC0CbY/XcxNXrci+hSsfTLOW+Ik0je1ZUBZVmpzH8UJgw5M6p4AOO0xKXX
/Up7ZKZbvuxPjP/9CVz31q0/wLVN1wCR0UX5QqEc63WLYlc3d9JhLeVlu1w+AMb8T+nMNXdHCt6H
/wIF25g10Vr8O2bPjCK9TOtYbTC4wFgDw0/ep9uJT0Zj+WkQyT4HfIFlhrlP+GSg8imki3sTHh5/
DJB4ehmW5/9RtwsrMLHDxseakPrrmX6wlgBBWkzBSZRQ9fB1Ar7mgsEkXi7w90v3jq6XXfcEb41J
WdZm1wOWKvWlLMdNvJgca1PtHoAeOBSZM5EiV7IUQFDEf0Py9z1G6O/8A1i4T3zzxJs2aWPR+rRR
zQpGr9f6ehmFKbF0cDq5YkeEhFQotMeIFbVWjxdkDVpx9AUNCcVbJ+ar1sTof8JvmPgYXsJryBQo
GxWr44vqTu46ik5nqgXU5Bs5gFki9xKuqt5H591QEOg+jvevvB+zrs97tzVZEeg6StASCI2CmeGz
Uf72wlM/gyM3lAL03FcqSSgxGqTxgEIq899XU1KkyhzNMTfkEU02FvH4fBNVmMXSi31Ixzunbrmy
M4zcZoHJDLMN4cpuyHi6KlqW1My6C8WTgZyqaBa4GTiFTrBdsiEtYGDqqhv6ecDX8CCp5z6Eto+X
sS8eJiFMskns+l+XDeJHgM0A+vCOYveBmZIQPhx+nir+UayuqIhMRVmqEmkqFiWF4i5ibmG4UCY7
k89qut/haFRDim1WLHwAmIBeVQ6ZH5DvniCbzGyUbOL4qbuG5jmpqVRS6ejU8+rJzmvFen+45SUC
y6Ih3CYBIYZX41RP2p1eDS2nt7WFaEsFry0NT5FnpGopV6hI6D5+8KYW586D3LFv5Hu0dKXjvUGw
FlNjROpE4+mVoY1kSbUZHJi8sk3rFVhzMsTJuyNU7kGUNXaKE5aGbAPVL0Y5YmW9hBFn7UItVIr/
BvY6TlrPod1kj1mrPPg1Ez/7Zo/v5LtsQgD7Yrss12XRUg/jhvkfZg5L7Guva82KFvU42bmUNctn
/dITgiuBR8jZA4OThp73AzhHpcj4kdc4dHutzMMWfgGox4QTANwWGPGuY0wRoFEPIMTs4nnuUd1n
z3DrOcZmySpCa9sub6Gqp7EDkPQRRQF8XdiR+m5r2KaTJ1hMkpcJcwDXilZiWrBKq/yBjyJXY9MO
jlhImtvdjVvZbAM42r3jh2s03kZEnUIhFqh28UgEhpjhLUamKfa+L0cTRpBzS8zQBMxlqoe70gGH
r8LjfwFWkre+1CU9GRTBgV1kmzJoLD0OHmYci2J+dfqt3HUAHEjR4fnDtM2R2THYfjdZqTrM2yRr
BbtISHqyCoVH6UjlEQZYvSkEEJYyL63ggv75pph7TqHwzpTpqMNA+Kn8AYuFI9xXPiP3Y/yjIaAO
bJKby4dc0dgiySdSXbNRvXs8iCkXWsYK+s306Dw6ktR5uaK9wIU9NRsO6iKGUHqqPE7FBCShAJ0J
w2VBWGijeB+cIJqO3/ZpSgW3H4FY1TR6kQvV0p/JOZjWEksn9c+DgdgcrNVQaLf0ArS1PdKmgDbt
57Em7uVm7R6OtNmSpEUHGtGPQLGbNJcOFoSpgxEQ+A03T01NfgB0nquTDDEgAzsdbS/Tld+YzaQ3
MY6XaM6CjAvqq/mx5pSUUyDsqpQFxvMBxPhWQK6DDZx89nrSUREHJuEPnay8l89h75uqaQcVyK5W
oJGqN9YutjTHxXg4H5Roelzv+zDYNOZ3ombD7RkxX3dIL+j63ThOYlVgtnlqVelIjjuJuQrR4TJ/
Yx6Qoc71tuxpNosRVyYV4qzbPiCA6JgkbUhNIs8U6P+gZPp+2HIBHO/PKDy46NlVLAEYpTH4pwNq
JkzG4aL1rzyLQu+2ie7ZgXRHXBSQTOBbf85Wc9FrLjJ2V1LX0Ef4eSXTgSTqbTm6Qv2EHdZa7iMj
zK7RLANSCAc4dSkndmhB340ZmqSnyNznt163Ia+XxEt/XNgNCYHmcJSzEMuS8wfwvVJqVHwZIMYm
zoBFp64Qw9qPhLS5x7Ma68dmT57VrIQb6shVRwAgXuPUt81J1tqofiFpaEiNuhSiNSaFkRVLT0HR
Dr5U2sTRzgA4CZlWaULBNjILmpGCuVuTvlNcMiKPPqPdAmsl1FB1Q+gAzeOqJtFLGUo2FxDXoMLP
ehe9z/VGmO7TA924nmHju1nLTBRQ+Lc0g4vglTlma+pb8G/NnwkmsQFyGi60dmQ+LznvD4SIVszn
tz0NAHAY/3p4HAi449WY1zURIHS70VpofG/GMaamxNSArwnoiSmoulbhzstlk77WrORzGCJyopmR
7kajhTaRpLLVdIoxkZoOPBcYbu/CYAb8802UVWzSPS5hCJI3Sn2K9HtHYtpwA2UGiicWUCUqJgbI
afwGcDgfRMW/B149VDxSj0hCbeZNROhtMs2J3JbGDiF25UnpkJSs98GldxD/g3KRf3woM6AjhJeb
YnzJ79nky1DDSRYPhuI9/gmfmgE3WgBkjx8XPZCDlRP74yvvngrvq5d4fIa3kQRhZA+2IbsLPXGg
rzP1iZXiUGqlHmOLOJ8ElAGazvq2aj270upn4miEjq/UvcpYpeGjV56T5G0V7HxALiPBqYDQPQFh
pa89mSGyxMGjLtI6qYRt875HU7sWtBBPauYAwIHm80rNn93UCO5lpDfiFYNsFHCS+CSE0HFOENcU
iqj9hRZ5nNdh8nnvjxmm6Z+X9XCAxB5q5jVAy3dM4SjegzjZ17JJ+4q8XwQkZwaEEJjjUkPEcocr
XOvK8isSGuC32QJKeP9QAV5Rcz5t2DuS4bCauYkulhernGpbin2qLysM8CyJ7/MAeW5IZvcn3si8
atXgH0tgFxYO7UqbBQ4U0ohEURC9nQ1xXuIzHe+AilnwhYa2SZdDgKAa4KuZvnKLGdY29ZCEjOHs
OSlMvusuxn7GgayrpeaHa0FCU/FGZTSphSWwwIPTnWDuG2HNAjw/BND7S1tsOdyw3qJA4Hng+4Vy
F9ZQfrH/Pa8zWPk0HzXNugLaIpH33AcDHDnDDPext1w4QzGhRgI6V0flYdQE6g+W8RqhzkY3sy/O
ipoAVQqutv6vO2D/dAd8A287p99aKuMy8Xcgc95E1YJRYGMGP/ap6RG3zoVtXaZw1b7UIYG/M7KK
LnzwkhgMP0y6JUagy2JAaj76OMP4CeyDiJtqnCMRMp2ndjGKLyww3p73YmUohxAVwEtDq/hWq3l/
XmwzeiuLi3ZMlrNwG7vuQbPV+RJKAUbLIsTIL/d48DnUL3fZqWfSFI1qE38l491gqdRVk+cbREZn
G7hgwWYpqu2jx38mbXGeA7Uqci4RbvtX+jCpcBVzGWfD8r3jJ5+pr5jV+XQADDTOIiJy09ASjs4J
u7Z+g2DjSgLmOM7VG+9iZWnjhO3OOetPLHU5QLNGH4QUtGKF2yp4wuyo+syMasKr11mcDVCsrnuA
V2hHoQS3OQybO/rKwncqDor637Cygef2gv5nR3zUgSWn1AA2UIQeffGOJXLXjJOanwI8m7REAWye
dSsIqvKFCOOe4TY/GtDuST/z19ey1Vz0sCWx8bMX981uHmCBQxD+acVHANwth5sh9maPYVG1su6h
z4GayX06dwS5YSF0ONpUoweBMEh8Yjgu2KKRRLcbfu1MW6e4fvyH3I3WCv4y79vxvlF4MMPMWL6v
tCnrzuoEY+5nHnPyk275hFmM3EajscY/KL2htVnz4n7n08TbeilBOvySxF4K/R2WJ8a8FtqVF5Ik
UQ9HhrBZUndKgVNKf6Re52Un5QiXdKISFcvzN03TTZDZqjknnqfpxwABTdFGL6QIbzUDylMdHiXK
cU7GrWzSE3G2/87M0IpDHGGWsMaDwcY+FKN/DdA3Ia9sNRyg3PJF50uAN+J1SmTuIeqWfxC2wolv
UuTiiL9Hal9gUYfGz2+F2fnhsq7teqpi5UC96ddK2NOX6A8gd0QHTxgw3yd7qKHR4qbwjstUDMBW
PW3dwv+d5obqmFfxaCEl++JYsT7RinArZbt3nsUyf/PF/ZeEd8kvjCk6IXsym4FCfZ9jt6rkIvKt
5G7rwq7NwHZxQJ+0POu9m5omzVOBBvxMF0jxKGXtzjuk0Z14evrdsE8KIaYdJYIoHJavZTuFMVO3
FZGD12ZgKU/0fapYMVa2aM/YbW+cY9OpuYRUiWlO4rJ3A/ncVweVDDw29vDdmMxBHHnhFVpBELiP
PrrdmPFqQhGDuBvo5D/nSYaiWuIy2bhZIvuxHxBN2O0QMwAD9PooGvOtjjOb7SnftgZ9oJN934NO
URcuf/KL+62klu5EpP8+8uRHT2fjskLB4lCPwMO2zio+8xFcmvYEpm6r9kexNDd0I8M1m0F09Cbq
t9OqhzhkBEd5qyyxpyALBPl7ZG7mDK5hRdRZMS9UTbOobpLrYiZ612pUf2DoU6s0TOkPkFSrbq8W
EUh2xVy5xZOhOqvkEthZ2fZhuMDZNM+yk/is7ihHdOltb1lHWBobpvJA9FDA+RdnymocvpmWg125
GiqMc9x/dGX1I2PnS7+jJjqx5AOJYunLPRLuGjp9NNRXp5LeBYyVDjPViL7eEv8Lc8PPoXd2kbdn
z6ciBnu+4NPI+YoV8ztSBuXTvJRGJALQFeKFqT9siSrZ2lJX8B907u00uwbr+xvDAo08Az7sxaiF
fBdhVNAJn2nerpPxcGIDZf7Yj1Y2V7EaipbzO6D0/NQsh8OsWCSAWt75MIDQpp/kPSdJ6DQRF6QK
5z0U1wGqMyuS7CV8ej0FIb+6JeWGKoe43dDuN6er2CWtUNtgirWS7Oid9V8HeUpfVyjFACYc6qva
FknS1dm493uoLt6/dUtdSfTb/OlxOr4O6ek/Ctd13i+W9WWnGge2RB1S4BehAKXHRC4sXMZqugNv
xxg5jhY/F9iWQiY9psAf0nIOs6//XIBtLwmnM4IFdGH2h7nFdjfM5rGYoGgQayDe0Kc4Ley59lWy
6IngcPpBGpq20BtW4WfReCPr3itOiw6sgS3uyZH8jVFLEQ3pGNk1PgVaCVzOqsUt564GCoJTQBcv
CFS2BdUwBLcLZiA6D4mGfriftnc05/5Nc0cLRPkHCeu75+VS00CqHLIiPBcOfISRughbdGqK84Jb
l5idP6HfbUPC7FtR5x3gHNmXfZumv12RT8JOJM3zcd42WgZy7aTJxOZ/EDVadaDQcKlSrRR97UFr
2Ei+c7aaNDasbVgZBgKO+4HN8sRYTRw2lHBL7Uqj0Fc6NbkT9MevvCNqkZbt1zqcK+jWwRRxnBiq
QLFj27xRAHi7Vlt5c7gaP0+6ny2yExfmTddg+l2TPtdBjhBS56TC+KIyw8SgbxSoMCLS8JjLZ1+o
Zp+GCPZMDkVTdIG95GQRbtgKddTsJbhqu/6FQxiOQYWNC1QIPTiP51DhJCuKnmxbhjDNTKB+Kd+h
La2kndK6A93KuppzQ0Hf9ZVFvIBLYcILra4iIZFl4aVKc7vXQoPZX6CnQkG/e75+6Kk/FNmMg6yf
2yvSJOCzxTvWOjL0lRAwSuAG8z/31fZYFsv3efzEcq76Y95KiuEiPV5/oaOvtFqj0LTLis8Dp+ml
h3LLqIc6XgSszeAQzCwYM3TtOmBI27MvlJ+CdJXHU2CWdSVzxqunw8OX8Cy4jIqOf27KsBuWjztA
tEZ3SkwAiIJa4DtWOZxa4RYaJzFVSiKMbNlKhBG9CThlE+JgR+7v+nJ09pxhSzrfKZipioLgjQPu
DjUmpsnGp4LUyMQUik3PadgdClb5kLhGTaNJ0321luJSUDVjcxkSnQJmcAbBNFj1ihaHZPtR9mfx
BCS4tFM9Boa8syV7XFbDsPPm/e7aA5Jp4GcCnhg8Hyu4qCCU92Q8s4Pqpe4gxohN+LsZ4DH3RbFk
9ISdk0MuHq9HEiRHdh+bpvD5NHM2obGFIfu1NkmnhEQW2qYt3jOwVane1I5pzdD55GvEBYC9r6w2
Q9tcKTSM3MlU1G3K4NHoDLj+yUL4hX3GZMqRbOxIGpcY3srp8i7iNKSiwix7C4gg0b25T9UN3ywr
kg6bGXCqAAs0m0xbPBdZFUZIZFQTugBs2OVEp6wIjTCrJalSMfQVpJgA+PdU8wp4sEny3aH8zKPj
A0HsLy06zbDc7K7xwk6G1NjZmgymrQSMeyGKMbXa2QG6Ux5w2dmaPI/2P2oikw+WDts1eQPTEkak
vcHsR1Y7bEiyQBt23hbJuzwpJcVsPjran/LwMuRTH8+Ygsv+8Z0qdz1+xvkQ9g/oguHm1Xg66vPh
ZhZ64XukvUEVlZHLyrikyZoySXgqthw14Q3iRtT0uHze7NBNbxK4T6EFcVg20HvTKlTJCScRT/q7
5hXEslAkqxLiv7XGvvDWU1++V/OekMOUS8G4uJGflrVPU0obHr4kcPrOqxQVLNUH9NReNHp/LIVW
xJp5R8zblnEaFrmkAT1Vfxv4KI9eyEOOIAnOMSoCQy94jku4GB8Jss0a2rWTeqcXvN+PzIS4WHqY
R+n002ezrm9eC72WKkJ8KI8Khb3fHlLs8h2dMJTQQ6lkmeLoViC/9gsp7WMPZ9vjQSowRBjWUh6b
gll/aNoNiNQ6D/BMCN6BmNVevJb7WrVUredYWDbHiwAbxU+ln2YzZWpBTlDCux04BZqj53Nds8IQ
U2B4fIYuPHDBydW70Styxl+6TbA3xEenzEI3e5Zo74jKJKF2B4s/zdoiFuqb7breBwadM7sH9ugU
pu8BU5GIpfGkn2GofaWSy15/x+5oOvO44zxS5K0Z+VgwwRqoYFgF/KAz5EqjA0RaYQFfm4hEGIb1
iYodcXIA2lsQKLGkIyAl3DcwS04W7YpsZeatebMm2tsMmj3mIqPsoa59P50ZIBFI3lItOPT+QAQ/
oyXtrx0p0VbPVy5BHOyD5b7J8H8IxPkouz5BLlkGcjgtCrLZWnrcuJr4hpBJxn3EFoJw0hvuJA44
hykAOGsi7fIr46sA1sZ8A/V2T/gvg/Kli4bzosbVwu3x8klRTDDJBH4QBewORtn/jcxCWIvuxbOQ
reGm7QCwzqSfM4Y1Qvhi/gO7SUsxYTGP6Sfjp4sW9CjWcfL4ZOD6+ZCN5Z0lOgWt4MHb3I8lI1fo
cMQAZaykrfkNaVtAv/P4j4lRqSmZ30/bEn/M6Q8bbkpgafGmJvKNQxKVcwgQ7qtz6uSQEqpS8VJR
eiIvvQvQdb6N00PyiJQUBIsBLK/nZ8KA7fPjYhjLTGB3lzJ2Tl09aJG9JK+MpmKoW/5CgWUNYGsU
evSOFFjscZCXoXwFQ4xzaHVexFLjvot9WkjinXmWZhy05PgOXM8D+Wo0Del1bNhqqDB9AsGjPVi/
5X4Bcqemjbah6dxDNViTIAMgLI8sTJCOEz0E39YQzu0iK4sq1veuVr2We9SIAoYnWzQyVqZrP996
/l1uD5jAwZc0aFFN3JC74XANtyg9Zl+8qQgMliiSOKKICs1beG1IM2mhVC6pBdv5OUfcGBW84DOT
dIyAmhY3JwIwpt9wTm3o1HazhuvXs2AmS9QDS4DnUPesEVUWcW8r62y19ZpZNRNtp8fjPMAOLXwW
4L56tW1y5T6eyL4Y9lRXuGZgKbkVNqemi8itYUZzwtRMnvX2mphRC/Temz3glMaGC4pULWTcgRVU
zV6s5vHceAGQ33eo0XTPPIiP2NVIjP2lzLad63jYkePzsrlUqRXU09o4me4DwFpfRb9EVO4Q4Vk/
2Pe9075IgJz4ytljQQRuH7jg2w0pvlaDu/YDbeNDXwZx8V5GYkqzVKdStwjp3hBtboGe38Wge4lT
EmdI78mU5fF5yeBq7bUROmjRL7TWpBglG7yjBFGGf/zm2kLM2YGwoAEpMOVV65wpPHAvlt0QHWCO
gmf5tcnfioP3CR2V4/mPnw0eaClGlsqPh+jMg00n4Obj3f+ZB5iIQ+7GAuBNibvYL3MWYs73IarN
pcJCajqE070oUxe4kd8AfpKTjZ0KCECVYHTpUrebdUguIzRl1clLeCWhtPZBmWr0KFe78gYO0ci/
wgWq2NoCOMSeGVFPwmqZ5B7pQWA7LG46k4aEwJCcrRWKysVWY1uMTvLAEHqSLmMbJgiCKz6vofQT
8II3tlK2njh1nNxn9LO6JJzhCmzfS389us2rgEBUwy/jaVgmtiHrspvzZe5LBvvoyJGRuLRGTHRs
EIy/turOCypldQNxY979BApHPtcjGBnJx1+XuTLfAfSYyLuVH7z/UgwvYD+NAmkl2Fsrdo+2CHDi
N3uTIbqXflK4WSqDjxSsM2i7wVd6lGjQtZPiTmeiUzthy7c2xVNKoHUjC24Rf7kMU4qzxHyVAgas
bc86FajLnpsblcUqA0C3s/6LyuuRNoDhZJG2JBk96hGKD/Y0vRcjgPvG1pLSiiYU+0TCCA/sgPE+
eXtSeFlvARiounKmt74xvWrqizzICLjHMgZuiR6LJR6RepX/djb6/KWfQ3xZDHbSv6pxl2b0zGRT
RcfNkiw/rPBd32QZ6+wvoy9Iu8euBOlxp+mHsLOCLoaJdtRtvYKF0PCcTJs898d5oye/X5+tB5H5
0sPuENa133tY0/Nakd73BkF38buFY99CDPq1hfzfSwi7sb9iuSRRV66A7KLUESptuiMBMH7G1fZK
KS/GSTuREt+Ngo4mRJKB7Aci5PJUHvNjA0/E2v8tehZGzoXUXSR8ayQAGXJIC9qayy+CcSQsTsis
PBuh72ojdRqu/c4ZCo6A3nkCK126/OA9TbHb2apyhj/s/T8Kc0PYrVbP61MYYxiMrtPZS94dJAUz
yETeAtQyeCex3fS5qxsaFRVeiEiv7ZUsWlTaKZWBq3m8UkKsjD4uNwfKIvnMVuI3/nnLRdD7EVBg
bTm1ihE0smO2Vljq1eBjr9i9IovEMCFzEJGSWX0LyI6h31pFHUFJGZ/ToUScBGcAe8MQ0yCe3xEF
Is7eiI8W5RYhuAL8H59/VIS0rWuRHoIx+QK9i15zgHYijZqg7UT/HJrypyiuhWJ5mb7jvrQ4cmdH
rfCIgTk7vV7FGJSFAwR7uVq2dlzkFdHiK4c8dz3puE4jn6DBxJcK86meFPa9CTcOQyeeGs4kQbFI
oOHYa9YEVWHHGv5U9u9mPP2iEwP28SILJcAOHQqpABOU6x2EkAXaS7xgDv+dLGE2NPZGYt8Nu2fg
fsJ4xJCGX9B0Dfe+Fe9Zw1UP1e8zU45oiicsC+AePpLDTr11EV4j1nHlOxk2XivAHfP+pnJhwdIk
pscf/HKvrmFvNpqkdWtl7pBFBtaBd9/ZNXP79EDF/5IPVGHpMCR1SzJVgFU43mwIh5MgnePwKZyr
xq3qkyiXESfVRSMQHco3kPswysPR50u+W0vE5es13K75mjfy+KoWROjkCGcOKrUtXYDFU+m1Ysna
UDEEPiOnPKJriAOJRArobXjG514KMEydZLMwel1+13jzGV/3h+euRa68mcZ0WY8nQS4zkuS3ObDm
w9+qzS/00vaIXNaTDEIahM+hXhh0eyaDYAMmsfb7gWgPHQdRIJtpxkwRZQd8ZR7voSqquwAPrUyA
ZhclSoC9vbzHXPh4nUSWvutg5dACvdmUzQqhyD1QPYSRkppg3N/WEm4h2q1wVLMyNcfVkDPMI8/O
2yZOsefKTDYvQL7aPVuCTF+6K1THbze/UfJoOj1lAsRjlxj6CjSaCQ3yVsrDzBRXccxvW5XaY/kB
GwIdtde4Nl9gQy43RywokDk+mJeOItDncnGB4SEoXBVd5LqzNG7rJBi6TUM/WP1KBgUiA/VFd1TB
6l8bzii3BQLVyTtGlZ/Rs8GqIu+z5wlo2aapWGt8Z7n47YnObNYM2sgl8T4vex7zhn0lM2fVMI0A
BmgzxTY3p0FyCcq+wcEQwGFN9anOvxK1pknDsfJdz6ZigG0LAxS2Vlea+NpV77U7mvZ7clCjnc+V
fnJUiW6E0kW/CUzLPPCS/opwkFSzqaudOy2wBM7ukgQtsQnuvSpYxaz93ARpHk8jNZDBVqxDKFl5
uvFmfTMk8blpPXYWqbFlU3H6a8TwWWNP4jkpktByACe/lOAMYzGETsCLYPRNIjRRCuiUO6dXEeFR
Nzx6kTYGV8iXDU49/sFXmlrH6QRFZ420eLQ3kDIUmzd945acioDskO+Nlw2s5haDhG0ZvsYiXMzr
vVTBLP1ym9za9H41CluNBzBjeMi5awlose9x1t6zWx/MdATtryQTTQZjH+SZtWraVvqv534vc+kp
kUoaRS4Ngc43PnB6Fhn0s4tqpbBe8UYD2YXmPcbp0hNES2bHKcyqM+hTTE9I76LsZ8ryP+SN9tnh
c+CLQNp7L/KeLMB11NLWVDq1csCWjcOh4srTztR3VghwZW5F/JRlh3Md5qeFrnusAU3/FzTuYYqI
0fTCM/qeH2+tu0vQvR/Avxs5po/7b/WgEdBJDk03/Zutx8QuxojiE8S6DNGwaatj65F00qPPBLcS
yPDQ6+GYnaEsYFftsPlHgnpQ0KOEM/OQZCBYAhmBvhXGvXfCo5G408EMTdVZGCIYz4Q+kXewRoED
ih3Rx2yHlTpGZDNY4Z5Zr2hxfTjdQgYG5LntQnIK2nLIR+1RXnhM/vp2AC73DxtyfPiI/zUAMP3W
G3okiWaB+1hj1JjBpCrQdvGOJRolZdAGBA9adWCHUV28uzyL/Q5b63XreD6TnM8XtcivpXA50pS8
gvTpcekfDiunXh/NSo4tDf3k5q6lhFVsowVfuA/WQSPBYyJKG6NZiD/PzYI/ItiPYo/NVY3n1rqk
yTviE035i+ogxt1bi6ugoRuz1SCV2/ZO6MqzRxnMMFiRoh06FoUAFk/Zhh4xekCtlIUnW7FORM+i
+f+2um/JJnuS6LbffHj2eOLsen3XZ4whNoOE53Ai8vN0eOBH95VDlEK0ChmsKjpeQYgbabJ2Ib6X
b7/dfa+BBvIGUDUQBaPsqvySLKcPKQlvDZjfZPJnmSunUDQwfAD61dLLwJMtRURpc6MnEnbjEqH4
nx2i8IsIEdWSPrmpv0X0U+vUOgq1ogn/eY51Fao8rNTLjJxIjiKEEhnufn/Wb4s1OAPSumDlvjjk
rfndT7OezgWxdo9R4OJZf7ElEVXGMWyQRUIqj43AQP3PKJCxvaoFXkouEN4FxHIrdZ8KX4wKtbxw
qc9lmlfguFyvdDQhiOpefG1ogV0GraZBNvD6ssDrQvAZ0J9gN60OucJ4y5cTtu5sjDidjcMoQuiz
QRdCJYYTSG3OulQBQkmWEvkJ+6QpHoIn+IYiDVkHbil7e0uLHy8oNPBiyMVj7mg5Ptzk58aghmKG
sQPbGeSyZp9l8clS5KbKlGYSg0uTaUlkJ2m6+gO/ztSnVSHw6BQFUpz09OH8AUHU5FbtnZR9LZN9
4Yo7ymrYnKt8ImS8Yq90Q8v1jYWRW9hrM1S6EHWbtALevbInn1b5OCeP7lwzVePkJBFNJFyu2lVl
3YBoBttH3hyoV7nn0F1k/yDLaqSzAdFWgLi9lMiomF1c2vXrcomItaelAMFUTZJJ/Z7b1+DR3TjZ
ELAAZhEP82FYaALz33qmSMBIcbhUwAsANX4Xxw0ltfiinrFl2/14o2vylULz8DsgibtlT3BgQjgQ
b++Z1zHDO4ZqdMUfxcObJTL0zNXfoQ/kf84o+M9Zkvsz/8K1kY5i8qzlRMHjo+Gr/lQMNeQX6ru/
mDWR36I0R4ARB3DvwOEZJqG5H1PmdDmP5a+NZgudVVq13Q/HH3Rrxrd4ijlgqNixEqUaIi3v1fer
87Mqv3pauX9kfZdKJRisNWLca46p59+jIuOcqvATEOnsGUxSX77zNB6D2mX7jNYtBum/f4U/mwVE
p489yfBEpxeyHPjxqKYkMlqHJ78QJfVCFjSegqb7hMcNYmpArIqIJKt1T9yUVZN+3NeGawS2TQBq
/SgQTFx3UVJidTX9DuaLDTQecz0v/hNgqmIgb6a7ht38ssfe/J33MRycDT5UnMUsYKqf8m0zXSEz
Y7UnVrLZ6tmdqzkNtenPj2VUPJYCwiWiVSedlOWTE/f2dHvX/ePm0uNVBnEvlNdrxQ8fN+Yx3omk
kmuHlR6UUrKFM2Gmhq4iJB24QkQUhOSLDhhBJP1/co0LrQyUkrNTQ91JYKMdnYDOVgZj8A1OQEmq
hMuUzkyST8YMeJGOC/pCqHQu2nh6phoIvszGduuQ6vpcbl1J89+mcffAlRo3WcNGzvKD0Z2R0auv
7/vpoxecMi7ljCwrt93bGBdT1YZnLAnmE+MsZgU332dD9W+BC1Ss+ozTtKDy5eVHbc5I+fFnQHbg
MW1fFxQ8DfBN1e/qVR+CJXNv3FfQAjyRT+IbqOZqxCG8iL4M9JZ4FZvFidZKiP9GV3RuTgS7stwL
oDTKhgTfVPR/3tf4pCW2S9VRL0kAkusM2LStKhGQwrcRxPMf54hcaoEqBqk0vaIv2No2kaslxFWM
+whM4OKXvAJsBO1b+t4cStno0cCBzTTWLB02o+MP8behAW2NAU6u3H0rOsK6KA9F2KtNb3izK9fw
OV6CSa8DOtsK6bQFGDPdWBHngfG6Wjts5Sy0FJM2Q92kO1UWuE8A/8y1mnbbqIAooTiTDWc4Ju3h
7Z6pPCVk/VvzLbhLkgGVfkCRPq8hPE1C6TJGe9qpR9qzbgBFiqhNmYBRug5o5+8RKC08UcFhXxc8
zKyQBuR/OnMHHhOYmifJCuTv1LWadnMyhPpN0PGHexj/KZXB9q2Cgcx9JQyLtk6NyeceWr2xxQa2
R5MaPHKu/T2s0Xn8Mx5t4oEgP50hN9EuRvF2tk7AifBn2FvfUXq4aAa3tOzMINb8caqacCB2InOa
P8jMo6vsjCPnVL6wYs1EWL/NDgTc54u/TBTFvXFbcfzxSuEvCI7ONlHU4CBXMQzsILveKIWoHTCt
g8wXz9965cADsqdxpVHgG0K82tU3zZ2pJ8S9rB3Rmooahonn5S0sHFnmLLX1ef/Pk0BWd78/MTh/
hzmennFq/uWnWM2CwnhugmDl256d1Z1WuLI/P4k4A3ynH3swu1ylsJDLWnowRRVXI2boufvYxoiO
T5aKAWzza3eEr6lgH0YgYRa/i24oM1aoVXcK0Hqc3bMhNbKc4hlKfS/nrykU5wdVNp9JO5gKM5Tq
hPqrOhVnc1meHm0OIbYQkFQvPVohBxVmJFbuqXmRO0cuK3A+iH/AKWdLknq2KH0eH9SxDWj+FxT7
HZJxeNZu94gAXWZ5p9kb81RE4pbSJAZXz6hVl7IJ5acTbklCgKUzxsLCtyINPvBVntLrgKgtB9aL
3c7ciDh7GdtcCFdlq9DQbWlrNHESD6WU7hLkaMFjU3SLZkqWFR91JCIDdcZr9YRP4yr8nrvAiq1S
oayWXBgewC+T8NktK2Q0eE65LwVcM5VwM+24gYWwY+xi7UACHO6cUSZl5Qsy2jRrAKytkxTEFVCM
6u8VZfXH9Gf72kVqwfZKoFgCZWbs4vyCKOIsb/ERM97V9Fq2iZ6tW/h/GvmtvN3edv9XXPjGGEO1
B8UpvzPevsL386egv3XMjVqctxK7o8wY9v+OBuFdBAJtGMkFMWOYVp9MC99MlXeWD70UoR3e0asN
WIf4mR1ZplDppYrtURC4eancstiUKZuj2keDQbsQtoGMjgAC8EDB9NQs6CJ4IysPFcb9zthQdo7l
HvzcPn1mzxDzpEb0YTomoZSM1cDHOJy1K4l6+Y4tTtNpWnzp2v/Y4hP9O1WeE3choM5RGBUGD+mo
f18sBWoTUgshe9qGZl0GJi8ap3AFj4B5KKuq/4n4hYMrIMm52NxaC/+SmqeXP/givHVWTf3qh2+7
1xUpTr4TgWPqPUXTlYqwFWlEwYTo0g8ftSvQsoiDe+zdzJze3k8JqUdBVVfVDE52TFvyfdyFRYnw
xaLvDaEdh8vJ5thgJ89NXFf3qxvJ6VzOXvvBeFXhEXdBGOk4le4bWxVpVUF1/axZ0l3tbCPrM8PO
UjL6ixXJO8xLDWEBhbTQ2d8bFhHzG//5fo0Ctv2ScYhf+Z4GqE8myPdGaL6RFfmkdzlGq1Ew+kNR
yPDddS3ShJQuNRYRVy/sUpGwvlSijqUYIBrK0NI+KIlRjLVwdxd7a1YiwhFBCYo+5jJzG7Gogwiy
o7AWvlnRB7swhR87Bqn3hbcXHmEQNA9+hWtWPsPpHTqzIb5x/kicwt5XTi24Y9Js7eScP75TVbKn
+K3APaX3o+5k+Bu1lhWTbiAJH4CU1c4mgFfcpPoHdIGcS+x90o0+4DwB48D97bfKiWjy0BVwiOLn
H0uw7P73lQ5WJ+u8lkOkqH36qF+WsdAkGJ/mjFEWUb1egQXXn3AyA4C1keQF9OdiBc81DTCTqEzE
syI1Fbf6ei3Od5joyftAgTYax5CmklQUQyDOMiPj03v337Awi9Diegcf2CcuvaBukqh36GQFCWh6
OSCV1vDMWF+SszaqDcRFUiY+K/Yp+TKJM2Ss7e4Fioy92oO8AUrqWmrljMpmwoQp4nQaclGa/7KJ
AMjQ1CIscgZAuebxmHB3pA9UBGTZxZcp+gaUM2qx4E9ieH6RrbI9giU7+3gpK7Je5js67j/YZQ16
CFPyqdSqiKVrgJwZyQ5fSHeKJlrSCYw88jhOFlh6yFe1o8gKwnI/YUpdW9Xd2XPBn1goHX25DVOD
wZsw/eLmicWhf9yxJ2lX0yYrQmDTOvD/aw125lQBun8tMGyaoqCa/0n1zQD48UUtjEL5+YPLu5xj
XfZYRttr5H8IrA+7R07KANNXMJ20I4cOL8ReHcTK9RQbPaiTNJ7PkzC2Wclv89OqtP8rwu9K3p9k
Oab6Hd4oVljqB/GRF6ZJDg752uYSsOtmXjY4t9vf2OISYwJX1L0PFL1yDWLl1NplasgwXx7Swagh
YZWwr1ZNqLc34K3UGSHPFkndXlVb1wQqTqjRUYch6pfLlRAa6zbNSY3Px8j1pKvLhKKTrQOpI+lz
+J0RPSJ6uSpLpKErBA3nVKhrFBUMi3P3hycJI34Q9JIKxg6KTvSe7Zr3wrNSGamGDLslGxm53yV/
5m3t6kulkP9yy6mvyZ5eyr+fnZ8RzMSTcq/MH4v5ZAry0rftAEwuunSmnRGwVRLJUdv6V3GUXY1T
YS0tf1MQw1yG08iHyZ+8idWZvw0NZZigkrRdhxnRpG9z2dc98jDWJJAdngqBV1UjXlCVRSYWpTHp
/SAPG5k5CdRs5nTCa7JH3v7CLaXnYuNpBT2Ka0u7YFEHybn0mj1xmybYIMncYiYubSM8Mu7eybGg
nCS+RRCUE28v/rbCQKTNFwcyxyEUsW79x354zp8FxTTPuCTyIceddWs7v+fyRGq3rBjzHLfyO1ta
SkdDv0YMfjA210puVwPOTR4FOqi61HLK8hy8tBT6xlDIWwSMcdMQOIuTFDjOxTIcNHnf9REkbvCn
LHMxhPMS25bBzcQq/FLsHkSpdlEZaJeColN80j9Kh9DaPuda41amdnASl5mezN+d3xEvQQdgsSnQ
3C0hx6J0tLlIOb3SU8ZDaErFwuG6xe9/2b3dVaoPox07JKBVn3sDklD3nBJqPpfBCWFfI8maaKu+
a7j/Lfmm0pL149NBB7fR3rQEnT12eWSptPe/G/rz1NMWUxUHnAZo3gsiTQogIYspkmINeFOEt2e+
eqJShAHnsuyUVqswQ3zMS0+9wI+jkAa1BnraZtz4WYlwEQIjpymmO7DEivy8NUK0e8KT7Vhxntn3
PtuZr5ptTYQWYqxUiXjV1FAGE33yxd8OIgtZ4zcXuIlWlp99/w41z1VH9LcHnjI9sd/w6qlj2GEM
m4pDy50QD3IJf74npcpTRwRdUkL3qfci5RWJuTUA7G7uH6eNiFY3GM/IVpYJzUPDUEoa5OIPHeNH
bTGuaeaGkwTNiHUvJoa2HGOpliWglnsQa0TKIv9Zct7uyT60yQomg+fBpYHtcJb7ybD9hOvM6ql+
6YLGdZVom3evSMiH5k4BjGLeLXq7UEY7XKcRgRrvTV0SIFBvG90qgvlsulfT8Xg2q3/1tEukTGIE
H8QLBFoCZMj6vRcBVrj5kw6bMymE/zMtik3TOk143rVlYUMFVhhkMwuMqoVZKwO+MbZqLdP20+bv
/NDSaFKjCCIzkH/2neo6n7Hc+qwLD99hsO+55gHm8yX/XW+Q2mYCTVPp71s2ETVFNxW6VCoLghwQ
kzYDwek6DGS0DWUcFh2h1iMtxzwrzqSUiSG0jbE+fiJglXR6ehaVjd4O6+0QPFN3n+dxDrw8pdAK
326p/DgH/a8oEWciAJN9o4aBYsNZEzllGbWtD2m233MCYGQIYdTeAFnt2Txsumga1FIEjFW92far
/ilSfNMrJ2CGeUDY2dRAWzAPMgFgK/u+SA/WCMkXN/47Zc91+aO4U9BKMntzlvQaSENU+pjNEmTF
VfoRY4du2TFkUTnSc0a60dzV7wlprdRB/935QnzFxkXWtj6XPsuTVrAVamBFZkxui7lnnHKcqycn
0zB1FI+YmqKeVI8VW4zAMCBDVO+o61nmhUY2DRdunuU70gAVSnZfh5hjQC3IB7i2R4809QY/3sVh
HNLWZQUjxybppQWpdpGdFgktE3xDKmSR5CXloC+9LnIkpU53klqXbdRYihH+v/pySQJrSrDBP+1H
6Z/obo9WsKEPZfkwOiMBviKth4YuS8itr6LbCnqqrNpqCNkK3lNlUNXUzEBRwdD2e+59Bow8BHBz
RVkQG5hyIPeCcaRr31rK5bvQyPOSOz/Fr1dZP8yn3zPvO3/LDkS/Dv7/HBbuOYDF2duJtz4dL4c9
srJbHHNvL3+9qLVqcWBTr82/sj2ITvZ15UUBH6etsihgEVN9RJRjGJeBRe1Uf++bSIjas8LaFdbT
C7PuT+x55N2YEhE1SOwH75Ul1CJtLDbqalsQyY9ifPVtOe2hQi+UCd9f0xQF7Mj4s1x3JepCBXkU
qilLOch0vi1GVYBSpDaq9/u19kV+rG98t7EjlJSgHoAHHeVwGv41CtHpFMbJTbGCcQ4z50TXC55Y
4ICNNeA+ZmrEe0eMok6ci3Iu7kxHITwL189EZBH6LDrwsXb96WPM+PLmCMew0zpZdZfjns2Wcrgf
zHh6h0aHuLQ1qdpNEsUTuBPuh0V4/BU5LMH5SdfyA3Rnj409xQ+eUniVPdWpnURRKapnMwyphkaa
V0B8WyQFgi/JANiLZtM6F8bGfODSm+XfuKdAZmlQZ7vR7jLtTIT+hhu4pTp1osOtmT2tjm1jEvFt
hWok8JS0Uod0PawEZhRsP7IIHyQhyHx2cQ8ixf8W8VdSTOCSpOWKKy8nOLCiVfGKqFdDJGsiRtU2
La5dUnHrHyOFTTsSjjyDsQ6OuvGSTO0BZ0UZRUM7V2TwOxXKJik0JPpSCSXlUYS5MkSxH8kdAedn
IxkXhxf/KbL4azzSkpOWb+HQWf7P9LjqGAW4falo2zSKOKbyVoWISkMq3fKK6fTjWqEoH48W9ZW2
0rgAs9nC/o7015wJyiDHMdxLh5fYMg4JAGtbIDxIyqX0fUup3QumCUivSLV5oFFLmae8dT+XRRxi
9czz6auKGCBfSqJh91UApkqduLif4wyfuQtu13B91n11A+HScGKbDaIR+DYh4/IB0ifSGRaDPIxq
QpacdJACN5TUZcgzKiL7pxxGFWol/tTpNlf71L9AdjBtj63dEA+VOXZFNwUmD8+vQ0PWHAgkW/ZQ
h/dqd+Nf1zgXBKM9Ac6TZIVXETQcKmoGLLE9M2op0XtM0pYBEFct8X5lgOunPDxXP+3ySIjBl7mR
bITCbyKu5yER4mn9oQ7LiICcTLHESZUVwLOVbEOP/QH2h8Z/7LewXCV9WbgasBTG7MFYcFo5Fntb
DLFxAr52wJdhIn3LF5L4O5y2KbuFA5nGM0Ivbj319Dng2lLCs4xplBvN1AbdxurZ4UeXtwBgldLs
/4/1Bh3F6bo+ZHPN2Y1AEB7QpFMeSFYhE+A540tr2AyXTUsjSrA9Pp63vgQsgkcLuQxcJMXF+k57
JjoCFFS7ghMHjQUFgcGo8ztW45EgVZpuV5IiTYY4+kMUUtPOh9QTkZHuOwOScD5d1qUt5V136Q3O
j/2buaaQwk8kj7aKhOP57wrfotM1GU23Sd9ZrFWGwzZFLsOGchU+e4B//JsKFxu5RqEqzITKtup9
Ld8vq7fD47Wb4zKdlHjQSOoc+kzuYjF4E8CxIPdHrlh1V2F32q5/NqsUNxAlYVwY/AXfGQo6I1Ty
4M7ItYryCpSBo8KPA2zwsKUjN1Nf7VzskusaMeMX488I6zvUoEOTJv+jSwKohDnwpESdHLDzVdlc
HzbVQy2AKQ8X6NmEJjrf4U9Jb99F2HxglfCm/JdDdkDdX37EK2/P9tza5/PI2xUJs36Ao3O1a/jC
XK5jKfphp6McWtdVVgJ4yzrRLlXb/aLrt00796JoGPJRtbv4A3Ta461u3QyxAPa7tKvmftRowkL8
10y607mkcaX5QhI9iR6XLqdM3gPnqgVPYlNiTp6vj3IgwVrywUHnzrePtKrc/0YxvpvoUeNl2F5L
8eycmyMkBnheV/F3oSyYJ0UrCcXJ5vCipmN34J/Ha85hMgQ1e2yfA7N9FZSNY6ggnJnMYGz0Ll7r
3q7xj6nN/hrxEUX8qCcM8XEpq0KcfS7HEmhzYZJy70SX7LcKPVW6kSlp/64UnDM7KCPT1juaPzFX
rGYTwmbK7XS2ZURmgyguwb3AQp23HvO4hlADbVJnv00dkRRQKXqjqzOlIHSwh9x9w+ov5oGEa7Rh
Sur4rDkItXkVEIzAdROWjUsooP26L4zbJTF07vTaxRaOnxAHZih9AXBelDFw+NM2g9f6oWK8fAWk
FEly2/59VFHF70TYJ/LUnPd3z9gpxpaqJaaxki+YValSdqvncFuM3UsVY4ysgt9/8xtNIOrPaxsQ
w0NBG7f73vdqvJQENGVhk7h/Ygtm5nfpDVFa/BTPPSckx1OhpYFH1B0uIIynZJ9SxbY/XsnNawRX
06HYu6fHon0VBkdx/1sdn6eddR2tq4byvkbV60I+v4NUbIe4AhsoQICpiMY9AeQJcqEdtPP+rrYe
r01wb8B/GVXNjBsucPkCkFJtihmCCD9rZ90hxJe7N2d/gkKLm74u1oZy0vzHzvR/CbpwJKjo0zAQ
2AUgPOMc390DWfbzalRHIuWCUikD4f0+yCQ4FveWP9LMShn0d+Znnyx+pgjeapLMk607DOzdboPq
mYIEovhRVV2hgPDBuuUasWxWYuz35v249ubcq8cR2A8+Ulvj5P0d0x68RKCvSpMAQtbLX+S0zDj4
XIQ3LElW64IExJ6hcdicU1R3+l+It3uUaa2koZjXyf8bPh8OulUvxZN28yWcYeT9qgJWw9huBOWa
FF0SW6cVHk4igua18q8b5DorrbJbeNE1wkfz9/hyA741/HgXyLTZ/JlHCY8xLEgLdsCGsxm8y/ZJ
0IPCBVI+0JeEWjK94CcJOM0wwJaZprF/1QvquUakQ0yQYq3oIr3NY0TwxDdrsMHe1L5TxOGhuyhq
n3o1nSdRxGC24AJU6hs4D/p8UeICzbiaaoXIXz272AHMztK0Mef6WiepRpo6od75U0BjDebq3nxI
WexGcnL2MtKQG/r7Xer0wgLvA57515pEFGL+YaqXxMDtOVGE5UivaK+GYin4Xzeq6F9hVLbMmHGj
8e5QQ9NLx1rPWu1NrHbePVOvE1d5xDtGwHuxx2la3S0KMMtwrMmrMVCUtiQ5OvmXnZbhmqraie9/
CeXs4G2BRrPw5GLqqdp+LBC4WZ7QMGkm+B4B+Zs3T1+SlS05g2jUEuG56zoJFCwWS5zghfPQ86Gm
/QPbODhACVbAldyV7521TAvxivT/s3AGBfyzLqZQKmtagFeoMJxbzc6oDW3jrF/I9v8ASq5gigZU
zHMAl1/KbOmJ+DBVsj75lduTjoGKrWCRAdcrSiGPzkNKm5XLoE3C4QWhV6QJ9Qjf4sJosiDF6D/L
BTSXlicxSMZ/ZPaWGH9szhde/f/0zoIafuZSlym3DJ1g50ru/sL5JIX7T7uaMHiMkd0Woh19pG6i
Bb0nE9RKMU5QVaG92RlV9m8w2fpyAKCjxjLSz3lI/dpM2d0ksxOfUyTvuCps0jm3ebtOGfeLaBWk
bndn9XqkKKpR1Um2Slokss7a9Naz28kosg0ISQNn6qzmy9HzV5FkhU9C4nUyiAYNxvJdViJkU71y
CN2rqDGcac7KQN39XvwAw1J8nuaMAQBZDF5SNKa9cPrQv4tKIIYVdqZJ1Rsuk+yR6AtxBHxWdAgt
ZXUXkB9i8YVEd0lq3cf43lVM/1agwWTOmgvk2LN7d6UGwCn0AZ/OK9H7Wco8cqj/jtzMCaAAGbqE
dFf6ulFMuI/JJtWIZ+s/RBV0huHijpCtrROveMRSWZcfvbHNyo4f23p8Re7hL8Kfo1SeGZ+Mh6by
gq/4MElB9jc/bHJa5LxZZptzTtYSWdgTBRrjTEPCQv8GTIBZ9xWvJwCG0FvnLCKkhsBLvSUeWH0W
GSGu5EZm1rj8qOp+cc0N3dxsICStFN3O12CtHiFc6CqWchv6Tr+xbZ3zovz+kqoGrmuXmukdqS2A
S1PyBWdvjTppkPKERrTTP7DtPKeOi1cWU6ZOxxBJ1Hm9wsVJsMHMKD2CADAacG7YRTFvR6o3YFZ5
CnlTa4sDUj8H1IEv/SgNkbptjJfDkUca6BXJcivHHlQ7LYxUvX5oPqe7kanRPp5UWQq0xrxedek3
WAIJw7aG/zhGrEyCoVWDFThKT8Pg5G15ZsOCn2y1JcV1IRqj9MgSoT6CoPuMK0JmcKtdFZ7iHmO0
4tZAE8VaZLiTsYjg/6yrUYujWz1ByWUE1UKdL/QcOv8JWUx4XXtAP62ylgPiLBUjQfZXWnacEVtp
s5M0d/pUz7cN4hos47wXtezmzA8dnvdxDcw3SjsOXL+xA2on1cYfZQ+OGlPp+tfxWbDJ7hu6ocOu
wCtaMBni/X/SQvZIcJ64IL9ohxdpeTGGFC2IoAQA57Dmf6f5aHbjw1eNXgDpzPU6sjHD7usAEV/3
XavQFPu0Zuo5834nNW3yEt2inOwTtOI9SLn76jjqEM0G2gZMFV+mYQp9KoCsFHMPfXYghcK9Mgbr
HquYFqIoiS0cC2tKZKyzraWc8gxYn+96cKPVeQWwVf33r+TNOGGkVi9cZCOxnvpe9YWQ74JDkCfu
+Wea18J8iqAq6zOwDg3Neo7xSo1WRK+M97FUvvQLtP8Uzq0qlle+JmQH3RowK92BAGmx7kdYDP6X
xwvbV3JpwfN27cS916vsLbq7Wxd9oGCIHmUDDDUTAo67HrghfwdcUQVHJFSnzTQcoH+DpGA1OhAS
hbZk1kjVHjzjFlVT/KFmI+NJm68y8DqiNmAnxgh0o8mF20hOD4Gv4RLtz+Jnj5BtWGWMnrA2dFVn
2Hxl2XVe9Amuu/oX/MYayWoZ9sLXv964M6Dm2kQTc46X9xbV/23OCKKHrH+XTUlpG7nz5X0ZgM2h
oRHUS4zVzIQruerdDk1puoEa6RBY0/9gGt5nbT4uGa9GkoYAbLStLqCQ/mD7zh4wVMvk5KtfN45s
MFctVkyFEJ0DxZWkSeUPIjJeHGNAhxjNXRryOmB2oXzFRTemr0NYvmIEc3w4mwz1VqvrKxM8/alI
l63E5XLB6m0ALYHyfVzhK6Pptre9GBMNc8Sd9zcr5jo+F6fYLImW8YnPcJNt5y6MPHstBDmytV5B
He5CwmPbzcFXHzpB73HFze1FQB9h7osHicIIRRivOZUTzrEzXx66bCVPQuUr62oeCidatLX4tvvg
AJMQJz/xZfyY/thmsprp76mt8aHfxr5u4sbOjHTCjqhe8nTEMJaiMvdzjUOZQaMHJbtbUjvqUSN0
bdXi7fZe19ekMnI8kUdvCQYcsR7UqNFx9QpZs0oZeeDrHjeAiPCD/AwI0PvrpvGau+hFZnOCJT1y
SNrGwTix2C4+kGXR3eFzRTqMp+2Mh4AUyIo9OzjNzXALZvwyeRbYt5d13RvkrDWykOeycCovNRLJ
BWWTQwp8G9rVDmtosdpNKevTNf0yDFbjF9WFinGHSxX/xw4TTwcqz8tsZ1iFbRK22j9XkInQNFUS
jfktsegO0q+pvRL5VM2UFXlsur4FADmHpUdDi8cw7Pim37L/QrbmtEXopN9X0wk5cy8wsC6tRFdE
IT5+rxyzrLzPKbKawigwBHcbCHDOuBw/QgMK+p/N80ODHRYOb24y7QEkTipv4bEsZLCqqP+BYwCL
LRbjPC7UNgct0oz4fwHatCSTnulh+p4sOE97PmlO73gEg46RT7uSVSrT3MiI/0GhRdmoAKp3gU1p
kbsMOemQQOLy1hjVmunrES8G0XmF1FInc/g6urzXQyRQ3souV96M3jHdPR4++wUNMYV0mgpDORFw
fqtVeZhmSgxXDD2sKuxpdGjixIN7UyTk8jfgtSqQJ+fNqZZbPDmK2+2K6/052rgshZxEiZJL6jmw
Q1Pzij4gwrEqBL7L5EgB7M5NbMAGrrdVWXxdloqdOc3dQweqUPulw+z9VYNdz4xHAwuDIUQ7oRbb
8yMWE/qVQHCcFMqq5hhNpF0aOYOJjabKe/UEt+NFihkO2/QIFBP4SHPgKmPH9nOLWeIWBGYpc+ok
YSzSDh1ueSi4bGQgfZNbXBrZ/7o54zsCi81i5j/9mbTC90QaKuXOy2MjVCbPIILQq/PK1JmOiD8l
sz+AaztnHLgvpMLhCe4NWsf+4EbK79Zq1hW0TkqhMQV0eA/lvTVJFt6MXcjIZ12LgdBpkqC/eTw7
Dg/ow+fdaizGAwL6b014VZIK8S1o6VpE5I8qOwEiXKlqJVAWlif/Dzmp84SsXcrZNvjm1Z/qyvcu
Jk8L7MOS4nRv6z76JIXPJF0UKTkACA2lXnmZdWcVm9HwAaW7b2GtmNVx5Iz5fWpKKHQvjKZfvVHx
sJEh4e3fccjkyMKERkuFrVV3mT0TbWl8YxVEThyDxPUYs7EwGlx3Z+KMyivp1bATxyylNUuWcLwf
7gFO8II89Zf3ocUIDR3VKLyVpm1S2J50J6gTdL3RJtG8P02druISHTufl1VUwUwCOZhmaf6yi8w2
eXGfhFfDEDJz82TjVqBBFRooXWAp+L3d/1C2Z12hMEtRXS4bgtcmf5gTicfgni3KelYzmSnRdFBt
c2NAick6bMOLla7dDR0L/8usOs/CrcZhSPRCIgcKE1D3FaYzSeoRrCyUv30tE6UxoRvEzCo5PiwB
Exi1SqfxpH3UoXycJEuCeT9PgnhuGp+683nLapbV4pI0TCwrI8gix0REZzfUXMCDlinBOwNJu0j3
HzfeU6agjXGWwJn9XLjUYzGgVQjsoTA80L6VSRevO9vpzJJThCeHhUMuctaBk3Zqgh5dvucyajhB
fZgXBsDfLX3jXcsmAFuujzp/mJJVv4xdvSHal0nKkQyqjDy2bZ2Xr803bcwt22YvpQjUw+kI9gIQ
/gwYCJHddN/2EYPOczB7Y7FcyCj8oVFdFaWaP7rQOdugblMEM67/i2RGQe+NouJH6yeTiw2i2k8d
Sl1jzYUtxjwoJaBRQkjIblXLCIhywuxdAFpq8Xo/6zGE4D5WJnUn7IIWVELIlTtVU8ktm+I2YMD/
vq7a1oLOjTOaA4zCRRon2H/NvJrOJ1AISdR6kjKOcreCKSzGB+w0ETfMuA+3y5actRt3CB783D2Q
dGdjmGUQckIb4ELhLlKbWCYDaQHJsKXk+BHMY9LtAvw2Z0Xpq/t3AVZVvLbxBNN/l5x4p3nuk7W0
lKyrFzpS0FnwpSlwld9zJZccPiSO5902Evwfkcbio+dbnzP88WJn7lB19jN34YZUPOQfQD4yxzQ/
yebg0l0OSmBhqpHpfU4AFqcYfSKWiXEDMaPZx9EOjQ8rh/aaYMLMteHeqonwCDGCFIdqBtR6EDVb
3fgI78q/5XILNrpjquOwYoJeuwibp/hFEMU5EGgO9LNhKTWwu+ZltfL12CtZaW3cgSfjpvaR4+Ze
K8URiWIOeQM08YukB4xpEXgLnXVWvo6Et3lLw91X2yGuByU0nnyK1Mh2VgF6Af40Our24PWZ/7pl
M20qdBaZavkfGNWNW3TQ+svWjk7avs4DFFEKxXlD4Z4rxjZMc3Ytc5szKRyEPKgKF8JZRYpGPB/7
1/DmQWt8ofUK2ba488EzAfzwasY9jC7vLCgWv+IVC/45XS54pS52W7tqVKoNGGoe4/aBl8GhEAfK
pGIUptnTy2eGX4B7hC8v/m+SThc8v/uPBH9a7QyUUF+T3ZdNPtadNsr0gFGxFyM/diaeQf74iVOz
ueMJ3175lfkF3o9G/3nd4+G1/FCLdfF0FYB5W6AJYhX0BRXV5thZVg8VoqHa1u/ymXWlfNX5Dfm1
k/AIl3qgl/b4gV6tlquqMMMNQmTk1o6RvXosI8Y0qBLiEeu0N5JeAesh8dH/PJXBQ03CeBxa4jfz
N3xchMpCxSR+/Yt4qCNvR3Qz//W6dv3444BSVSlN4Da5aK+qu9pOT+FSNKGNBtRtJty7QSZkH8oi
uVMiZhB6EAoNj+iBdTipMsR439SZXBm5XM/F1uX7F5W75AZvpqxngythcu7Fi5V/gCY/Ay3ZElwB
Ds/e1Tmur2C5p1t/ag+u4VCf620s3fk678EFgL4Y9BnfS511pnLLrd8dGL1hX0JtFuoUlBE849mP
HoFiI/xdSpzMLOViWfayEVu0JL4T6z8GUfMaxaY8h1ayXmpsSuOyzNU0LlwUDWHbC1yRGkWoKrPn
xh8sjRZJvn9/yAAsYrdi98tuy2o1ecCj+JDQKVvG1WMU8xOE3ii0L9npr0FOmA04OxzGtdLNtpml
jRRGd/V/Nt33TFzNlU61bA8UMLm2GbPRik8H9jSLuWyajroKakTyOIBi/D1927xPFSqTA/S0lqSU
EPZlZjPgY5LIluMbfHXYhcVKA6Y7REY+MH1hwXcthc6NQcEaKbHmONymGohCZEjPnWIhM5cO7y59
rAvcmCJVP0o3kp6WWqNMRfXamK0LF9MgjJC7yV9EeA6Iy6Vw9e2ZBpmzvMq06SmuWYLcj1T1KgKF
KyT1GdFKleTv/ncHGOqpj6AUS9fPAuo7KyB0J/Feji++RvH8av765EdU8uuWbweVtlWO0mmOYlFZ
EEBtbcyqQSkwtfiwfP5SRo76hT5tPODevuZHzo3jF7ZRPcB+O2IrwfyLtZlW+8MJL9b0Xayt927E
ILrPGEfkp2Dk0B47XHpn2qk/MF5qrjoj3bqbyQ5pbLpjPycRFIVq9ut2aZWbBlOczA5Y1Wi4o33j
N2v97V9TZaNb4xQhgRcBwM4zzyVkIDQSE6doTOPkq8LKVHQcZRMZCNo5Qadplu3b6T8ZbfzcPfM0
NyVNDII6oKyi4Ys984S18GFR4JI88T3ER0+v+8smK1S6OfVVfJMjNcvJlpA9Ho5lgH5G2drGAKC2
E6ahx2BFpGkObiidKS89p7Hs7EZ7KYplK+SziUP/XfDeN/PevSIAc3Jb03xB0UnPqrvpExgjOaun
mPuD35reNLoXPck1+JS7cwf5AsE3V+oNnKA1vFQC7lVsWkKFzNXbHC4ds0f9xrVTGhur6e1vtKlr
cu7sPZU81IH60C5grOy9mgWCbB3NTIW2ZkC27FBwh1k2p221F8H3n6B8xuFc5ZV5DbTWl7CQOzCy
xtBRuXv4nABvoc4EKckCtjIBYRSwWC9yGm3DqI54EcJr9whTrXBjazVajHgUYUdVaRiavrOraJOI
banMz/c4LRBmF15BBmzeQbbSwu/WugTAx/WPraxODn1Mn0YLpt0x+/Nc4Ji/Es3n90yv8rTUJV0S
Pju/R5ITj4hqrK+hEsrcp8bnojE9gVIFit8+p2wi3SPHWAyHOki192gFou2/dxG8Rg4/0c6zStNU
9HNwQYJXnUvka+Tgz4jV0pL9SfPJoTnBCk71BFPgFxd92Ju0N5H46fD1xNh8A4/IRYWENbflXW7L
tIjfX9u8HigRNEuVkf6C+vx6izqESJPwAUq3zTQb97cRmYtcp3qWVenYEF1ahAx6RrYRs2vrqFzL
rEr1D4zIH2uK2lVtwAgYNCy+QplHgXRNmDxrvIRhp/l7ck3OLpklJ/HGg9ckYmR485nkXl2fnAKN
NyVK5J5V7/do7GHJQ1jSURekG+fWlu1dLbNDHMCXoyswdXY1EPGkUjlmxXKKb1DqUywQl/OTn18t
h7IHWJbpWnQJFfq6wlZpc4dUY2M4RXkDGO4n3NL63OvOME9hklO6kO0p9q5mC/YDY7DjD0uPtS6O
Vv+3LSy+sGe9e0aINLLOIjNt0uDri4oWzRahLG8PI28uqDQujsPpCzfipPJqZqQ7hYZRdu7mXoox
v3IeYfQ6HoDWwEWYpBtKxKDDoh6PV220DXBBjXY8lRwbyy2RJlNFAvjAJV/RwxLZDMYntREFYt60
rQojr9A6C7iPJ83ohh41Wf+8YsFWfORth0peqUEsHkR/Fkfs9NI8mxCOYHBWi6JDHPs5IPCHOATl
Y9b3ZzG7p+Iy4lQ6eq3hjWTiXLVzli6AgDV6KenmP3mjSNnwEVgc3pmWMwOC53pgewIRUGDc2ImO
Z9j5ettzW7cfVQwmwwDaDH1Ua5T/b7fz/VvxLNaKjJdu2Nbenlshkm6DerOU/VSzSTNeF//hT4mv
gaOKVhY3L+NiDoAIs0RQ12xAdjsZhtUKPTkfzGN8FBc0AnpT4M/jCCUjYBbOsoXSh3/T9lIZsqX/
7lQyywoDU1QfY0bMhuQfZuy/a/YOMUjST66qrFmCq+LwF14e+pnu9aJvBIym4EgqRABWlmqfciHB
kBlfdFBhxcPXKTMEN9m3RuigtnrEc19GXfg9TT9TlM1xaQl18D7gDwkZtyH+bdoH0c+4fZeb6az5
VNtXtLI8to5bHIR9UVAbV+7MdOk6ZAFurCJRQiBWBVB6b9yuY87CX++i3bETTe/86YdH0FaoXJ+z
aJXGlnKi/GMF7bsi07RumA0BW03a5r8WaXIdf5ls/9HzIot47EDzwdUr9+oCHjwfFgN+yRSbjuX9
vc41N6Ygwu1m+tMFEUgAZwM8ijk08xO+GMoM/MIi40jjlErzF6SPhvRTTAh0Ym0/Kbng768pnLT4
k0T0KhzY6RYZBHjQLwk9Ya/DngVJ3pHcwkTVRUTlZOD8/TLhBpecPcV2H5nIEsbtRnYICXe93oX1
AUoC175jjvtWbNnG4mJNfBfi6hWCCgbaPml5VUpxrWnwsRtsq8PLxGwTWSzk0QGcVy/mY6vrItCR
x3PPcrqSAwCsGYvraU85UzXRWVo18oBuIGrD9P/VJU0jHsqEW7Mrbn+TM3/elugMWVQ6RlSMJbkH
DuFdIJBBv1ik1ggWR1f16UR8Ci3KJaXrHS6f3BIZMhbtrP26iEPEvOmnSK+CkqG+7pIMDmE3GzVc
47p9m4fmdFkbIMGB2MpqgMcEWltnAI4VtiUNwTG7BE/IEWeU/FEkGEtANu+eESa46oPc1+s6biBZ
MlMCx+poOYnHhSlPo3b8WpKUM2Og2YkY/BB6U4OOJQ/gV9I3eDbIHS24Aq4aDOWAhkqz77yXtyat
tHacPM8i+1nwFgXpe/nen7XkSEXTikrqzsCHOziTTEr0gsuquFbWIg926wsz/ljaGQqkPhjlUILm
rBINmlYQ/ppupiXfAAKfF3fe/f8l6NIHPXVhKrOHos8mo+WOkerf9AWF4HtEkiJojz8+Mh7UUo+7
VnnFIifaQHFKPXdC3jQPcIvtXP9ZxPwwSdmliw56+e8/FnRHwisfRbviwyUd1baMgGSpThUBfEFK
Wc86WYeF5rEw90nqgj536KPNzxTCaIh7DuPVsZuIFG0NNjJgwsBv43jM+QXyYjPsPXaB02MnDjLP
UM6IlCLCzttG0D+In/5OCBMbQL5cS8aTTXU7/wN1+Qgxfuooa52zKydwzKb2SjkbdSAKX6qyl1mo
FDzB2qvvhDVrE32yqabCJuKbLJczAdyURLSBqnV/hrKm5BHw8ySqt/gLImmhmBvLvSL8CRHDUTLa
GA1J+Kd/7IJ4Ku5cbvJIkFpTwz+c6t4vhwKZFUxrLLopX6gfX+lX0uhnhPdDys9RFPF5ZRe58erv
9gvx+Npv4FDxaEPFhaTovAjMUBcmPi2tUfo6Kpcab7lvlg3YnW+Pr9HbrlOnPG3HLd7Z/NaiWGQ4
duetJcAscNC5XQ719Y1qqeGDppyG2RPMOnu5clEtyezhADfFshZz+E/zMDzb1b5nm0mC3nt6aUqw
YzUEWvtCbKtqXjQR8NNw0bW0JTfG47QpvZnT7pho+rkE6LtlJN6IOwBtQufzB4TOnzYro52EmDki
HfbxR4ijoVCD51CAsRuiJKXLQINH5I12nei2q3tv5tNfmwAiAvHMuF2U/81YpPLCQQmLLZEZMgS2
M6LDZxLei8GCK9NyJW/xysuJsIU/noHMQbcsflrEwurv7cZ+RQ8ZJLu4pohiBlployWtbFNZXDOc
SRunl0xeiLh7th2JeGS3LVukdNRUJoGCpyOzsw2WLB/n5aV4ppyvg/t9mntL/Jp1bQoVxdFYkHwc
BZ38T9bdPs4wGrld8+LrhJY2QE51O3vTW63gjkTlE7fOxNODNDzepFB13+psZ1zb+G7noLeeQ/5g
LG45UvSxEfgqA0OYW+QQGr5SPJ496ZQkBAokPHEQrl3YMOR2orYVsYhrG7vosKvKn0Gqy7NRsljK
DCuaKcvFbu3QBTTrAXUK5l5U/poGIPI4J18dmoK+Ayp6fbNg6M2OgCLsmDJ7lOR9NdcJbRot7Xfl
x9Jarj+kG+d7L1+BA4XBVhE+WAWL98ogMGlSLJdo3JHcaZDLI83LDXe/Z4lxQHPMn+ZrarMtq3Ok
4gHLBneIO3+OHjssgoVn02rHLBi7qQwtjbXtQyc3HCUC/p5nmSGvTthn2NMawcJD4QMP0yO9TYQp
k6iRFMmQHI8BLmIyNXqQCkGU89GgGoBYEiuhHrBiK5qSnKobPfeisuRm4zDKGyLWYzJIhlHTSrcn
6Fyj4FW+wvRK/mKAg+GlbWGQAtVNslAXzFh2ClaEqj0E+2e2DsA9gawucJ33ILputhT5mvvcOFGn
61DT3//ibJT5e+2FpXko7WVskvC/nzSFdrjQtwK6EoMm/nZLGYlGJrarm+MltFGfRoHMy16hdpwc
xaEfEpIqc3ehsFD1p/mSArduvI5Uu+MUeOHOPIQMezFrDEChs9B+1zKQUb0R5wy+W/q4m8UrkSSE
fQjaoFRB5BhiJffGTxmRdD5upgZWn7/sgZt7X417C1OJrpxD9uHZZeDtcTsbKXSDe6lcWAyXb4Dh
ZMEd0vbxHSmZGA6OCPIilk09BzjDvwhZdEEen/K6tZPM1dvYb3Rf8+sEDWd4S9FhXdU0z2WmlGlO
l0kyoFPUw5NNw7EybLQulRt7NHwgLFPFeBYT8JWxTVZc39KJ+SV5wXpIybOtXowYUENqcyMCyE03
EDbjRfZufd9Dp4n3rk6GTIq5UmWTaHm0ViAeEFl28bkL9gJEXpvWyc3BHX+Y+cYyx7ROCjqBYxQG
dnfAbHPfW+eOi1m29ffecsZjind5FaYeC8AteSR1k9QFDW2hBHBDU57MlE1czrY1eXSOfZFT+lWW
+A5AWtBgrNls96HuS/M6zhWoQGhNytBIkYEXKgb7SOl2Q2KoT2+4xlkXWy4w+P32dflqaduahjF+
566jWcrMwHNTf+d6Une/Fb8bliu6ZL/LdLP9Xf8AfpBrt2qAM4w45godqjHAUl54njuEXLqJJqVk
K9Zg/UZYHEAzQ4NRA6jTiXyRAV/In0fU128tugCZ1N0b2n6XlUBXl9nrqAiZALsjtOVhEmeXLDPA
s4DSRFIbjiXmCRCaVIzDp03O3zWELdp5t5++3UhdKBTYEvBOgiDpYq8e/Jd1Vc8UbpXA+mrzNXy2
ClydL0J7m9aYn+x6daUk9KOsLY9+QL+Pn0ef2ORZJUDz4AgdcKpB73XNGByEUW+YpqZJtMkuQGuu
7bBrFjcYQsyPIupIhQi/lh5DCDRmMGeiBy/A3lkT9vhJ4iydoUrTR93Vr8B+QncN2Jc5lNKxkmOy
E+K2m2LOAvDbRegtpqZRx+OfBuxu/cD8iEPflhmriUbGg+Q7fa9RHcdH4DUeI6R17HrG/60wC346
oZgrUhW6VT7Fqr2UPWIcPM+UINcg+RJuclOCs6eEwEkxr2ioUqPwsZczIaWdHL5A+KT+rbvfQVYX
OYNMBxbUvX2n3fRTgToT8phl4Z2r605iKlbKeLVLLZuIg7LTeV1EEC8Ssgl3k3zeYbgM7XAu2c2F
QlRc3CpyJ/pQaNT24F07COZFbvS3dTZ4Jl/7by1UXTqbzX2JX6K5IhF1lFzUmTi2ElkR9+C8ZBUP
K/7/JQB8beTl452H38lyCl4U4Al7imzfs7GI2xOeECYH7JHu3GyqAt8rQfR5ttor2xq1hVELgFz6
2DAZjjQedBm+izsaDNNO2PpAClSSuojUK6Cx2DW9T+68rNh6RlwZqtgt9++KPA2QBs27M5l/VhEV
wxKW2Bgmv0txf+WPvyZ3rhYk2u/NZYl0G2jqDRZ5LxyAdKS7Up9flo46t2cmhLM8DB/s/EevN28W
J7t0AYdfrwOJOUJIIRfif4m+bjxH+r7cGH0s5/ea+qpMb3Z+rQhP4bD49JXXSZxCfALleitJuy/b
7ZsENidfP5Td/7caWwJ8Cw4B5o9l3mzsFCBSBkSvV+L9eqrcN3R71EERczlU5upSk03pY7hqv1Tb
3jIk7Gavm/ndRaEPb2+r7fqfCp+ScyEcO6ePraieBiSF8JBbxmzuddny4IgaKtSFHVmshAohA2XC
UtRMQp4aHHEIlFV3mAi9eiDzC4ahj8dty9YxogjHZbYfS9tX+E5GcFctH7bfqnhTNzBq756rWeL/
wwlwIcBQS5NuZv0DHAKr2cMaZiyeK+3/EAA7QCp3NlTRaj41RroD3uz6e6IVnhE8v69G6f5qhDsj
QqTqAYdotrSc6foOF8YqdXRYMUQCX/rJdJtsDo4U4uaAxbY+Fo+pLT3fN7k/OVqDn89fIpLDujwg
MFRWXVCY9LBpq9bcYI1WgWwS7Pcu9RptD1uAbw2d9UjjGy04x1L20iXYmzI0Su86IVRqgsDfLaH1
SmRwuXxrJy1I+VOwXCii1r2Zr4GFjIkqpy7jFyItY3ZYlyifafAlpZSnII9fvIMszgrdbotnbq6c
GnF2GU1a0+bCqLJ6F1jvsv1aF0tq2yYleK8Qu1vTtmi31FijEYrL0Q6MehtNntZydMiSdo0QceY5
LnOBoYaEzzovhqFtASXqq+EDoo3orWm6yq5QISsYUcf789KLdRipPNPm4b9eeclp3+W93Gjs3XU1
ZdEbjSwhEiCkmgavNajZSut/jeOsfAKvPRl8O10qDx7uhJ1dO40ZHEvq5jGavc0t2i91xLjAQkOx
pS7ouHvRnEZw9HMuxOqUmB6ZS2VTYVJ5weHuX9jLtlJEDPTBTwGhTLyuySPqNB0+DQCfJANkFn3d
ouqLmo0C/M1kd0KidgT9A1VcbygeBcmJhF9uV0f1W4b2AbwRvVpAoS/hX6QcnKx0fNew6fjsNkE0
a/ZfCzYuxVLxwiJrUGvWpUNVWt0VniHONLjwMuL3mCtRvp4QALeEJOj5n9zuVDxDXuKC6KPnKYhE
Cm2eUTgrYSHBSV6aIL9lfbccheFa3XbXTYUGDjsmJIBJy/W3Mqde5q2Dz7tU/0Gq7OxqekVVmJuH
OfGtTEJpNWEdvluIMfsysywhqPEa0DjOYtIQRc2txFNcYqTgRC6zQ86V5vj1+09rdFrv8p4pjQ23
IdGYJ34rhCVgg2Llx/OrLpAS4wSDDSTn60F45t0sjQgLVRaxLTNhsLtQ12RS7SmIzi3GMEfcKxQr
UYheybZP30yBhz0jrNrLMHh3S2c21JCds3bSdJlzqIf09PrgfM1N8fC+oQhOHhME8b22nM+ao59S
pN6ksoQrRBKulF5GHdWXAp+zbsuYGuzIGePEqDawwNTyKKB/Fu58pQG50A7CsHBqNTo+B4BnRm8w
LNOAI1VkUzyaTvTAbR3YaaM5XnJbs5MEjGew+eEqvWdZIrazC4Rx87YwTfRsav95esyF+4yOOZtN
yfbjDRpsuC8F/Vh1K+z8PzT5he6pGD6MJiKssmgfIXRhbeAT1ooCnMM31c1tkjzDgCa478FUmNfy
blz4BNwiikkNWglbKhjpv27JP+/xcAJ/l9sN0G8mNceHBPFywr5hFQZOwv0uc9omOor3W21fW4Wd
+KiD4wO/Iqb7QukGDzhXfuIJ2DJ3YbLazyZp9FgCF2nYuM/ePJkl/gGg8Ko99NjB/oJLGbUsNJ3L
hOXsXksfvIJBL/ghoUQB7rR/LgacOIRmadvIb4TPVKMDy240yJB0DTKU4DiDOR1gRn9ZFNpeJOYH
3edSWgUxGn4J3g6qRd9vGAwNyIaMfropPHJoyFET5YOhWMPx9LAVOLTEQKfVKq6Xfd6C0HEvq4/y
HWGj47mB3cEH521bu9zUIhbDQF/VE1VqYwmKDcyKLvMDPvocPba7OTwwAdyoeBDMBgfEdz2d1VNp
DZiLWijVoQrRa0lqSDWiXVh2eGlD5WR4ZoYr85ptOIcH4+jEzRURHXlUQim2MPOe0LrdGgebLTce
3FgmXIfjvPYwlWsOmvXDQztOa5wxEpBsTePqr6opx+P/Q/Qvn67iDE4ULI9REPI5Em3wexJH9vFt
FnHH4G8op0od5L6NChUhOGWp5hygSu6wW/Dw1C12skudCzYk43nCafTPKHYDYbfMR5fZGjwtHVC+
si1rPUcy6BxESRdepuWAIGd43PfraxeldXTisHnnoTD0+wYO3h66nIne3XxQHzpXUJISpkmfVNqp
l4b4onIud9vU7Wc8ygLLAuO8uY2wfqLgNE9p9KxDDaGbLY6pJpPwKmahz2SSMwwvtnvJ6ADj4dZ8
LdZ0Eiwlmwl250zEmeHYoxoppUpWzxkhENjL8XLxPwu5zn2TprqVLun4zDxm+LoBnjOwvSa6epco
Cj9E/M5TpJiXrUjWWCFO4zngsL2C/8iDYOnl01dwytwXp95xxWDU4UG6aAxP96ABlK3tb17Geagt
ii7ilgYPHNjiRmKdMJmwbFtTUawAjnMsyf2jFHYGUDkeaeX8fgJALj/jl5RnnyLBZCcR2i634Gv9
QTcbid3j2Zci7KAhc7CrCt+UcoeXClCGDHEaNoXKV4vto0YVaHYDbuxwdJFu6mvYrBWrf1yGZWvp
P6C+G4ph8jvSyxRM2wjtO5OhSrj0ejIHxcm6jWKFR1peI0SIOuBbIP2LdcsdnnJzsRb3rNKahjhc
VNPgaPfNwgSh328jiJsQ0w6vO5BW+lNI4RWq+QphiwZDhhUg3B8E4RnvCs/prRgpts3lzfR3Dthl
g1x7tCz7Ou6aX+AYLLykLgEGOeh5v5Fuwlw0AmR0Xb3X4YtFEPcdojdBw/lLAx6uZdEErDqhUfqD
Zdwk0ogagx0r3gp0a/G+xYtUjZBk49NlggVQBgX14k2UClRkKlNZ6KkPPmjtgbASsq3TKgppESB2
bapeTvXeJlQRC2dZyk/AHUB7S5vbsimeHQjHgkdwdJp4VIwcZSiJu8YKrfxCtuQwrqFEFneHj4wg
Uoc4s1vBsCXA7/q0uoAK/H6D2Ie1sEoqivxVUm9tuwL8AUJuusNl1hKsXj62hGCMT9sIQ0ZTftoa
pHwIld43d0Bs8VZSVPNtB4NuWYhoq5+XJued6KZcrjthHhzwtcx/ofO4bcTY8V8K/WlLb4wDGuHx
62wHFQ09HS4u5RBMn8i6p5NWCBCD/7FRN/1YoJKg5oIfe3ig5myxuR/m4mFsVq+TkO/wyXZD1yqI
JBR71A8LCjnKyroTl86ynZiajfskiFPp4hECq5FuLen5ehg/Mj9j/YWtMa36wFDdW9BTJFkoYhq/
d/3WePvY6oh1Cy9OKN07lM7s+hGXh+yiKQpzY5zf+smykR/8nPArZWkf+TD7CMsCfwGnwvkM+ooZ
c0WZsQAi04L5ynuWhfvwDRiiHrkn4r804vmxiUoB7ansEHXyJydo+FTLsegG/2AKfX1TJP7nssNZ
6zWPrLowiAWRliO1BqTDt043+PhQi16WUViDQPgQXbxRRlRvtjHEBgPaDvVxVR3XsB58P0v4XOBn
0ZGpZkGtWGIoGQwxh2AHOmshsH+cyx377Wo4YHCifHFqIz/nGtFsMfCMdXhuMSgudscQKz86YEXN
aouXizOcUww49L6c7SLkJSFsON5uoydDmitGEzLkbKqOlLIGbi9u8peCUP3oELB3IF1RCjFx8+Ml
oCj2SlO4WrqWzavtSmfyTfdFAtv5zJKAToJhCDR0iSu+y/WqlkI5HqaIUcuYQniQp85nH5TIqolt
MQs/zyOOhfsFa9EBw7HgL3DEQPdoy4hnvbnxDmogCHKN6ANia0sSX6QexYRSQ3IGH55Kr+fDdrcS
IQ==
`protect end_protected

