

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
px5VQscCY6Ikn37Zpcp1ILfeMqUABKdTg1DYgjtssW8p17+5AGxXn8HlpYhowPTnVABTcqZBYssq
AdObyoeM3Q==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ULCNP80NmeSESm+VisdoToUB4V3BI2wtpkjqCJWHR3avMOuOH9hW1Kzqfa87rPTMl4dCkihqP6P9
9ZmBjExh5gD+h0lDqiHiN5EytFhUn0BcqqpubbuthpQCWA8Oxrjs1bPfbx5dSTIg3Nvqp8n9XBsg
3zIBm4RI9QAchjygG20=


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
dpxwD/lMzAim75xo3jZkKsZtfZe6qNlkwrVWbOSfN734kpIMJDy2GDoKNkLpwDMDo+Zecq1+AwiE
tmbFfvaR5mEtpQfPg2uzfev2LBtc078lTLd8ncDvbmeBwRJoKQAWH0neS45DPlcOejtPpZEQIa9b
uP2mmz1SR9Z61xN8tyE=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rr6iRR9plfwfrxqfZPPK/a1GI2z53pneLmml9ARqu0imrXUHUtUEyFMo6AEqx4/kfi5+Z4Rxjm9c
IA/bKhDetMTUI+nIsWBSQgLcipv1W8mpcPT4ZcfmDqpU8haFQInt6nyU7K+izI/Vt3RcCBYoeiN/
bGIiqkyCSRrthP1yjTIbhI97e/tLoBbkK+iBNmPMRfkzpg+bewkn2OODAIbCn5IL+VA8pIS5uJe+
VUOFnrkxw1o1YyzTM9AjRmjDybemA63FaJRJNbFAfUyvCpMIascoIkE9gGHwPUqjE4uzo0rztZBe
UeXfzIZSyusOnktFXuJ3dMX7oTItjAu6c0RYqA==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ASzWOmKbEsU6RfaEV2ecw2nGdGqv5D07B1n3NC3ShFAQd/w4c5bSkSAeC7JKsUtSWRAwy5EUu4du
geIW8EZPtSd2pVcockFIFPjVTCstwnzAkzk6zBWiPzXCyPsh2TMr2rueS2uGUpQYo57ZlPl54CYM
qVCiNMkhSdW8vFhZ2WxrOT5I5BLTXGcccwAaSQswGuUM9KxaMur/gE4rT0xFdG7icki8Ey0lIB12
eOpXev60WDh6GD2m+hFkzi/rEM/pjGNRDkKwpgNd0ZU75yNxA+J3RBK3SGzHww+WkIZOR8/nBv3r
/uAr0WQsqKl8nzEC22SgL7YL41Qy5cvgLOOiBg==


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Mz3sBTo4agfAvSjl6hbjqGw65Ht5H3/pguuwMPjZNFVD/QYmZuv8tv7Duq8gqQ3IZfohQkzGZAPq
o9lRfdhbfXLxHxkfD4WKD8WK0ZQlBndVhi+/4BEcM77/9KNwgxrYgViFc6eAxsyj8nKgiRcHNA4+
8wjkIZnQtQp61nQ+U2mSJfyu5xp6/dtysq+9iaBIpHAndbuu+CK4cNrDVq3x1z7JQmS2Q6uTy0PY
iaW04x7+SrEuLUC2/JX2Or5radCI/q7JOETxwHtFhCDZJa3sAQJyCFLx4GnqplVFDMc66mZcYGng
6RJ1oWrP2cziho4GCU6GDdrh1xMQcq/5zWDopQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5120)
`protect data_block
FLA54R9Zjr1EVrk0ON9qqgiddB722rjk3iVXnxvEGqZsJh05stHMKhmTSvOU6nuqmr+OqHW/FL8R
IkajomnOJvFMQ2+6nB2mw4uSR3yctdjvlUMewaH3/6slMNoQi2jmDSjEYUaHFe+UV+lrIwGSJkI7
WtX3F+bOEIobo0myJx4xw2gVn1CRtb/woOcHqq+XTpzaJTtTxQk5J8VkP18AvPWzqXhql1SYbWgU
kyiSgdVI9wydwo3toofwiLbReNmDhgkUSvMwzUDWAVLSFrS6K/kJFp4yA7ojHlXQIZR7jeMrFqQE
ykyH5yEaDHt6BcVZt3Nd8dUevm7shko26JKmZGQSQK1vXKcdRnnM7si4Ww+CLDjCwTgYU7npS5Zi
s9e0/L98alRV0c3hwrpnup8lbxF/sowh+Y+ztyPdNGzOPM64fvJrk0V8wKAJu+RCyGmuwtt9mQUU
3br+X0XBMdy+mK5tsD2PibwZ6mwUT8o1bYbVGb5z2qjW00w9EaOtLVk9QvOfT9jPVFqgIU5kAx4N
JpFXmxNCdIo8rQhj75lQpjGgfWcyrUXQg1FjnVd8qmU+Mw+n9SbZANtP0lAvo9vtw3ij8+SzZr7p
R6SiBeZeJfglmdH1+weyL3qQiwxCk5bFO34qLAwbkWFUycb/J3XwnMy1rTtl4yjmipd8h7nrRz2P
YMXgiepyFSNORq/VCAW48g/sYqdHwiSVIa9KBajj0iBuylMTL2i9ZriQ7pHFsNKlorZmXOoJ6OBo
qKNyT2bC032XsXa9qcvRYQb1yFbpQ9rtZaDMSEirCfNA82GCUS3Fqxt3csYZE3Kh+kgVOgvh4qjq
zw6Ga1KuQ8Qo6uH4VXYXHYnljGQ6AslqwUPOI0vAjMA1SFirNk9U8DnIsJHwA2gVqfSdhth1ub63
mwNzEf8zYC6p9AlOAnhYxPS8Sv9hhupvb3oZOpOOEri2oI2MvGa+hVTVJkIjqCwzmbAyIOn2/9Lb
5UGNDHKevEN495V2ZHPEhX0M+rz86lYS53HHLrVBuWlNbJ26ADr71d3kOeDc4iRrvU/JqlC89HU+
tk7LnQKve2WbajnXxTeUos/abssLWckb8eplsIqoh3Nui8k4fKCBtMz2+Es6gqBFSJzIcOZ0hg3H
r4ok68TdWADlrMdEiHAmIvMgbl8gyqKZSwc7CPHqKDksV8rYj0jLGvZqPO2o4ZX4PZ0e+ZEuUy3U
7xQQXQtk3zpAFBhCc9JVjf/sdwCB5KsygK/pIf3puDAdOq3spSMSvotWNQCINeuf4PFkX4nZBUCI
fduL+zcjAsTJHC+JTANy/IH7Uen082wcAd4cV2YnzPPRFNoGOF/2v0rmV/ZLKCiLjXeWY8n8Cr0k
1N/OjEsBfaNplAkfct3MVLpXKNyAS/D2MQL1ZYxblyqI2ThgCWkQkvCS8tXFoo/rPSGBJLviC1rW
iib+svgxbEd+/HfjlAtSow+MMWtzMs2LBAp/z+YzMHznoJbBPDPRh3ODLKHK70+/TZxaap67J/Ut
rN1WjAF7Qg77BNlvtQ+/yiQsnw6nU5Uk3Z7EAP/lWVvdZc9tPjpiZdncSAMVh5gccd+fsDR7cGCl
fyZDcFDWERly6qThUYrKQxs5zwigKyqzAv7Ru0npSdVBuoimOTAmM4Vx0vkui8ABSJHx+Lb8+S0T
nL3vgM1BKnqlgxlYzXFXvQvciCPGdMqRU2WxAlEuMDbshBtdYlnsZTONi7ILpB8XBlpuJ0jcxOU7
z9SAflNsyepeXkk1RwsryPh6dpEMk2zhS4qvZwoV0un3JznppdpZ/QOIVPLOL81xwh2V/FJT5HE2
6rc66+UMajB7Cgn4d+leK33MxxikdaU796HupXxQTH+8OwIqrqxkXOk48vXmUFDtl3p41Yr8i12e
poSQobWMW7P5BY+T78HeJqJdMR6nWQvRC30MGJ4KkGyWsxXqpncfPi9LhD3ttDUXHBISQdvrTvZH
SHQSqportrGHsMJ8v/ip4tjv2laDP/mc+zphIf5qNy5XRxOPkBHomkgQCNhfRolJfVluzEckE4Pj
I+N2e/uNURZ1Il2sP/DpijbGiDnehqnz7aBjk0J81FYsD9Img1jk8Org0cknE1pJgSZWHiBF+O2C
4k+2IpHaQ0kjh9YwvPttOMXkBOHYLVCxVY36qVYWBcB51homdDzXufuMDRD+IagQPQn3FDnzVJB9
RFPUg5/aBuR9J90lP3AQUxOUsGeurXtmVU7cnFUO50phVsspbm15Y/nwSYsnMmub8qj6siQLUL7U
VKJjR8tMReoHYDH6P4WfsvLzIuDnVmEoiZgwjJ6dOzulz4pBGSWCQQi4TzR0VzhR2unEXbVPg8xK
I8JafqQW4dFQ6ERWdOL/lpesJ9YaP+MKrxdpuakWC89FdQ/hQNcm2nV4EhD5TlHzhMNsIrlGUqry
Bh5UDxJIxxhyRSYvf8KpizC97qTs3ExTb5BQQyAude4t7+NrQPi+AZMgMu2Qces1gZY8HnKA//6A
+WzBtgqCC+TAHgZWZM+wg6nMqKp52rLnHIPk1Lwqqi4BhKUYpNlWd7Im7/MQZJ4lUCsMX4cC8vfo
Zs6ELHnq8xUKU2dxeMuuXAPp9x26rFz2icGh0/TP+2WdG9aZsClGr35WS8WWQESRQcQsoNy4PqSl
wd+2DtkHRWC1wHu5V6UDoofJg0enL5G2++1MQdr+zy9Z2zHy8KaXu7aQoPJuB1fkda2rVybLaWu0
wzs3msZ65+YmwLubGCyNX+bu3N/EnC2aeSQW6ubs2zDZqL5c2HRbH7vEPjEzFgAxCnuvtv5j4S2I
l0glo82zA1TNK1JTjCOkOxycQzwVrPRSnAH2i7bY6+7ORtEgN+Da6SKA7PySNaMCVHCobrmP74kS
/twGRwxklaRaFXryrGM12QES3iVdsDshwN5X7ReF/aOAb87ERjjihwOxDgxUzn2SyHcfbhX5yR+w
iJyo+GWyQ24AU3/Izf6uBZsNhgNZ8un6RtNVi4oWpzTs7Co5aOQYUmwnnM74ScR5uIkrd/YVLBvg
KWMkJT7dOBsdJ/Pk5AGq+Ve8IFzh0dNmXA0DrLfzttjKEDpJBjBHD8f6F7IyJOlpAntnjF+u1a/a
t+VB9a62UzNczlIFhvsIU0uq/Ixk9awV6t0u+gRUuF5jix2GBRg9snzLwYh9WqAgx2rZY6AicO4f
BAZjIKRSbRjPTFpUTuV7Wr993AciE+zg4fnRa6l3Bz0ok5lolqhMnpXK6zkSpDpe1/7PNrm7eRGm
Phd4Lie92n7AfdZX/wOvbpu2QErPBpRTIT6KRCb1/6eiNC19eiZJXvbXib7NHhqhI1IisvveG97k
72B4FHrO3eSNv6loAuLeJdYXFqMxwIOp64MIW5+oE23Ji4gG7p7jw4n/6rqUq9xjjCPZj0GO0zH0
nB4NIukG69XepwN7jnZPEKB2vLcSXntaaODng0nZ0Ezq0PuewrqnFx3FcZ888vPoVBxXpM1NJuvn
x1gAyZkdPCopWRXhuAKkjMWYq0Jhre7g786mQ+EEgQ+UMn9PX+BR3ZK1Ryzdv8GrX0vZpYw6uz2s
rNDfrlF2suN5p5hhwDd1fj4H2FvaKex8NAEpSjbLV6C9qjhDcSj5F9Jgsix6xf16GQ1mOvtbZ+zv
FbeyfcXDYltqSIbZsvTYTzCELC7GfLBNJUYnrosppKaV6sfrrLNcqSJRoNe8xiR795UiMFG9S5EO
DHwhZ5KZ5Nxbgp5ddv3JmE7cmGqc/SsiXhev2GwetKJhHqRoCK0I3Jul6M+cJEuGzDi2gZlWn7Q4
fKXdu+QkK+LTcUrSAZroQKRNY/gABJYc1JZtsQtAm7tTXhqpJQZHO2J4CV6yPRZECscENJ/UZFn7
pIcrS9p+QuYccUqV7mDmWJ82d2S9LRM2z7l4Zb7TlyjedJBGSRuVkNQOZCftLXpyVVI6qPLWWZE/
szS9O6dHQwUUPvS9Ee89osUxnY9nfsfiOVEmDSnc1CxjQwzBX6hOi9inNcxemfiQ7N84axcVPrMU
KemqSaegFgeDgh61yRsBy8D4HYvFwkP1AL5ijrtNLK5onjEoBWpdAgMpIZnAL3ebxa3+38/7+XGb
XpjXriQEr0u54JZ/J4X/+9bDnK1uImp9mlSr2YaXOd1CVBn3GEojrQAf8/iV6DuR5F3zdNyyUheb
JkmgXbFW5IsDb6lfUt0lFY6YqbZQT6YrtdwURfoECQf1inBUs+HloVofle+DyTs2zXVKkug6Yb4m
c5TNHzvWc9+CHN1/XsxBzaSgad3lzGs8xeumOzORvKQondxmYe8rawNUcNHV4nTmYEV4kSSKt63w
vQaIwlVKsUq9cn28ElYlt3S+fkku/JqSzQMRPrF6q5ingTxqzd4zl3wbEyv5vZmYxD1KrkbJivRY
gmoqqAbczUX/eN1kaNtqeLKGdUdLKojTgcLJMpNI6qD9ExkD3XK+N/jIWUX0NXRGPcsuj0avhm+w
a8at9q5tEb0UwMm1ehppWBdRRhUpB0YR2VWYZiV8iabn03zHTBlNQ1gCL82Cn2YnFc9vp884hKQu
cm47fJ5iYBDknZyBfgEcPOSHGXc5eWMMVXHAe2rc9zhRJFCxn0ECRgVZA/8PKzlGVcAGDF4ulrPW
tPsoxx01cABYw3Z3uhbzHdwmZWABTtitgIp96+xtEwoNbLmxeaXmyqteZy8auEZQ6trNoc9emm1/
icD7xKb4R14dTIufRMnRF3CliMk/5IchegKkkmZeYfgDGJls+5/GiACJnFWQjf9cZkrTJO0B2hcr
SlIw9HYJRl3Z5NR2bOYqjbojRABimowCb+ZPreBTOe+JEStEt1gDKJ/IYCH9eDt9x6GyzplLowPJ
J5z0iq1bUrCZAi23vh+reqwZPAHkffTKBDt8lOWe4fLoCeOO4SP6V3pMFX50xZ5Asxv/PSe6Hdz8
FEjOXdRrI0LCOYo4eBrxPxP+RdVRf7GgpAMuu4eK4/kVFv33oG1mpL6nno9Kdcp2KP+Gpk7miHUy
cmhVvzMnAkRaed/4Q/xFOg/0ABwygadDarTDRxj7K4qIpdziCbUTyPNdPti3dcQlt3UECA6kLVVN
4C4d/yeVC2oWegdx19LK6NoM/zYrLISdw/m9SIkryq0uz02AKszpTj5nn2PBxh1r74g4r4k4RUHk
/PjvIMz1VvpCa59YUli9o4/Ce079YlG5U+rViT5GI2OVOcL0HVMHXKrl0sMCy+rvIBrWpcIFL1yO
5wNh0X0aK8jXIqtU3y+LwdeUIzN9ANk+Ico9fCMQtIKBfUYNTwoJL4tkmG9XSD15G3RDkk0MgN4b
YqE4R76uVLcANYCcfSnsql0wj75w28GSSDRfitYIhuGO6PfBEprTIY8MUXYu+9CxLMt+2VzIvHic
WLmQAt7L1KGaxdtVGd2kzqWJv0poN+l8wainoiamxd5M5msEMoN7p6TxnHToCwJmzLqaMpz1i8dg
vyu2kMJ0ul/skA4SlvUjBalyavQumiPY906KzTwnUi8hEEnjeN+94IWLxB59QJ3mjRWl5V+26yBm
fu4F2Tf1/rQs95M6WyfFrpyUm9H8vpHW5diYSfKXBL+of4vy9foirJ6t39R0xPKbS4L/TXkdu6Ez
3ojhScLtpCnoA2D3wBBCxzXKvTTGFl/efr4QaGqB57Y+qkwIEDEMo+yEVubdG9bFxO/Y/p2n7oc+
EIFUb0wEPEk2s+NeXU/hTvRmLGNWCjhDks1oZ3jLTkkIUgivVXFzCJeyO19WYKlRoq2jon8sWw6e
Tyz8+MwgxY/z5Li4lbp1ghFpdYZfKt20MsIgaZhgnvBbn5j12ka+lI5W2n4k8vyT9J86bZh0pkkm
fhhKO2X+SLTIHE5Nc4pUGEznU+vPNBM+mz3egQlk0fYyMpriRNLsyx9/uKzbcbwzXKG2yahThS5q
VY4sUbM5p/l9AqGC/zFUDZGB3J7ywXbq4LNSu2PG7jd/50WuC+O+PHp93gonCq0rBsbS3Hgpn4rK
hPtBGUEC9yGJBkkhnnqsbXLdUo+h/hKJe6XP9D68uXAYGA9U4GlnlR2Ro0UMtOex2g4EUYEoiY8g
5SjGfdOo5OyoKffom9QkOe3SJeZCmWu7D8d0U4vN4kyDS40x/LSrRPq9C67i0RZnBaErLfJN5aVe
jdlQBqfikI61Rs5t/s1iJOC080jUHN/vt7XhEjmX6hXav21/A5ncY3zYOkp+CfhAk7ZyyRM9aG/S
P37FqciKnaPnkaDkj5JjufZWV7xBpaezueda0V9Vhf9GEx12M1WUZPNMVWnS7iAjXg4/vnrq1rIC
aDqoXFB6U4hm2h77mdkQG2ps5O+9Tylq3TaGAYQSLnXe+zIIA9DtChoODYL0Zt9dzR6iNSabbl/K
zNj2dAAnA5zaT96Dsoojll0F8ce+bpTi2ArlGBRXxqbBkpaCMOOmKRLxCgLdGxWuJdCxV1KcHb1x
tj6nzslGhfRzYJgpTj3IrHG1+vWFWNcU1uXlJUhLu90mKTHOL9DydKE5BzK98OwAi4b0qU5ohCml
WMw+JvweDivVs0JDj8ZNNIo7GDt9M0NY5a4wqD6AFNJIZyFNU8y4tDmNsoiLmMCTv8M611vy4fEo
8QoYlhsZj7FzS5UZpELpiLme9xsCvL8VuikEwlqQYJ4C6aLfzuLUNNPexEC0rAkITxT5/L+LDOAG
6Ms6zOXKbvTzCQc6rZmj3jcnhWsBDUK/KfMtPLrE9pJjv2vxjhneSFLbtVBeqrc2ehhh1JdrJtvQ
Vy8wPC1OkMnFoLdo6GB4cNxii/W5GX3jyoRpAQeDhWqfQfho6U6xpGVp+utT1qk=
`protect end_protected

