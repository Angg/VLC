`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
lSrzbkVRez7TSrqtMj3fFBoVDIfcRk6Ys0Ryw08YT0xybeh4Imxhh4Xo5waHds9EoAp/p211hEtH
U6pvrX+agg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
icUbHhj5bYGT0RXX0Hkl3qTy8gXjmaBdYmbJdfGSlDqT36aBG1MHxVot4QdFfhzT4y4EGe95lWcG
bY7yIo2Z80wxkaYltPsUfmPKSryRYnC2RQpCalRwEyIV5kwyjLyH2PMI318/DGe2zOgfAhyaJa7F
upzBPe1dc9VfrYuArL0=

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
PxuYgPP9isSAWV6BDGFF7E4+ZyEAPJFkhVqMkmalejPpQU0gnnWwnBm+iezC17JL/Xa/VJE7sfaC
AKrBOUostq0vvu1xdTV/TiVQSkSuCL/ILd0KvrM7zY7byDcLHbE/HiK9qAiuHZ9X9afXOA3LUXa+
NeIijoXYNpcPKApFE7k=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
MiGbO+1/w2LzUP9w4vcJyQmRyNSWoFP9CtT7NIPM6EmL2LPHcWpvAOqX6yz7ntfA7Pj/Wid64Hgu
shoIM7ZLSfclvZdj2d/qq8ODrS3OvMB2omZlH7/9Hf8BNQx5cdlMGt2EQPapbaczdAOSVlqfQP11
66CJpcIpu9PYPqIPi7gr0sPciFBMJNEeJMdBTGrQns4LBfJmDRE5WdPDo1iDs7+I/XoFMkZhvL/0
Y91WipnQHvefAAlRLwBWNzObJ2omUnJDqA4fEy8FyO94l2UP+gXZJY6q7Ahrfb11AzhWCQy1/6kO
U8WeGtgOmdPeP2ApeGCjofaQkPasVPK93MY9gA==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
J0hRzoctT5uNrkbAOYhG/C1YYiqLYlvZtqfLxqcUZK7708gdRGZirVbjbqEBeXYlyHsw5AvqFtqw
52FoZUAEGkFlwIgKWxiJl46IuvZVYEef2NF6y5tgMHwEjkFVh359FztlWhDp38jj/NzWHKBOuK7b
WD+057fNTohIPJ/bd3naYCO9ZKinhXefS8bjBLsa/MNn2ksi+KfipLV2LY3t2pcBC1wui2dHqGvO
RvXXOCVCULpb1KAf8M0xySyzObSjDR2pgz7PdVOuusTxXaD7SgOSTCuvcYLUI/CgGUFhDdSfpo/T
KUE844cAUxLN5mN+SZcv8YXfgpboB0XGbtZjjg==

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qRYjS1MWZ9AEGoXk7XbPnWevWA7a0pAx3waQwdjQYrYZZwvwBmZMyfVb85xxDCsnqBfY/X+z1MGN
R6wP+/VkRwqWybLkCI2H+eY/JIxV8wnXukunleMgiWrZralQzn5HM8wFmhN51HFEHt8MehA+1v8V
GkbvyB+NWGe5V/g+PjZbUP7Rip9Ktc37bLfQ+BBs+LxyODu4QecoyoLN210+e2fQTtiawB4NhORz
sjQ8EkpqOIGx6NCgriSXgG0/5bBCy/0+EaWSre9yzV96ovJXPqneFAFAykHGk0lwBtE2N2jTlUmq
4YOLU9hzvqdkuVeyE1y7f4GZCgyIM0Ch4LciMA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64000)
`protect data_block
/PbXr1dFiE9t0bPa/ahRG5b5GwV9F0+wW4TFPebdMfYj7fVqBoHagJ/mhEfvdaUpKJMsF9kmVMZV
s1S1w3dHyYPHOjFW9PeYMaDfkMVHGDUaHp8m68sdo/jSKroI8gqnEldZmmNhFIVc3WGSuWlz1Aw/
5VM8GvgnCfC5BguEsfWx0ugOdlMqsIotscw5bXgMI7fy6Ve6Epjl+wQjEPBx8bYp1b/5BuRe9aM6
H+FhMzFtcWklDKAF0H2ypWCG0Ioc1RkfqAwIrymuCspg3ocUOR/Jqua+CqVl8q/vgoRHPSlLe52J
XRyrJh/bTsMAJFsJtfnkCvGRVxEx0cCyaNipCaiAY4g4/Z83OEqn5yZN2pz+E+89zaxTsCLdLgY9
t7r1BWeEvBgexca0eHXfhNTWIbGFfVj6t7O/G+3K3lTD7ygDTzRUzLatAqUJVXN8Pdr94+I0RFs4
8FS4m88o1m0OWydqdmd1qIXDhNmBcQeujP8BeB6LVKn3WYuixp15jy8+opoVi6g6MixRBUWAoHMK
/ZIxygqgtJWtN7Kjroh420b/k9qsM/QiPq0WrHRk0t/Vh16f37zou4xQ9Hvwg/to5oZRkin27BF3
PzisAAPVY8OzkALN86mBnF9eW3Z71ESdifdHYlS9kHzq0PqKJ0I8IE43hlMmkJOavvOdxNQUYRMe
XZ74IPaj7NpM1wRwjhiUcV+Ago0lG7zCp5A39s+KDk6zfHfT5f2nE0HP3pCkDn9xUtxOECDmIR+K
hEIpAmSxfe+fhLymOijlD9hVce3EOk1Wdf0bDyIsWI0Svn7GcvPz+mZrFlPeIWShcoPn9FPieysr
mQgxJCuLlgfEr3gsb3u7zZ8MpxVW9jTRbuSm1mGmzFK3KvmEr8+1DuuhhGcNBPq30R+bju8cNIr0
pWyMhkg4TlwuoMkqrWMZYJ2JEl5Gm8vrzc5wQSo3FLqlHw8h36XhPFcz8qRonD0vEr3EPCIYwro9
2jaIH1exUS3hRcfwJ4PuAcPTz5uJqkfSqzwZwXafYjzvra5N9USRzMO3VaiHkwPmULSE+5F+NnH6
xq+mA/Lr73Tk/mdSL43Ds7DwknFPBE9yhp2HIVCnsRQa5h3fwcFmLiTc5Ese4U4TwI0IssKaIPEV
vjaeiMkx5D5OaPpaaC1/tx9RhKZVWCcZkKs6YVVvcWE7/7BoNtkugzASbMeeljjuqXydGAjVgQkq
BT7OWQYcNPRsFXxCoC/2MG6AQnhqzVTAqK80cG1Jm18+w0jtzZvJD6R5laxZ5DAeVvxFqhy63+0w
SKePhcDBRDS6x7hm3KU+hh/gfF/PSo7Q4/K9Evf7xn3wV4B7trSQ0B4gPnKWnJlVE6yoj9M0dl3U
TecImVw/yUrvSpvxxs0tq3+fcns+4yYChQoJRvaOZ0/P+31F0P6bb9GxcdIvqJn3PbhHf/5vwTcS
86/2UpLQEgIcAIMwqUT6Psasgolb8n33OgsOAOz9MoSTvs6DnztsLDvkWJqIllLGkNmRciHKAvWb
RRs1ibVjgyIB4X2q9J2RvzBzsB3GVaiQbKydF+0DRqRyPzX18YENqrb8sgoDrvHrJBiPGusOExH+
KtM+NBSdMtFQ2rI14zt2UQ/M/h57RANU0N+gfdT2ZC4sZP9Lee6VOvI5UP+l4gvQ3pkYG0o1uBzO
Y0jYKNelbTQZDWHY0B5bizRRsnrOLWqbelyEJaK5lctnCStzUVU3IBX6mk3JUPzSEJYsvrObMh1G
sBirBVd8Lst5yBheiePfHW5Kp1tllHxtuve4Bi8/xtUg7u4D5LzYNKwi2/vkTGHehJLeR2Jes3pL
KHjjWJnICNnHS6CuHcEd39zXXWn4wjnTAW5BeaAF1FnhB8ITUCRC94u8LTzvmgv2El37Bm5RfU9q
RTzOE80EWTyeL/BEBrJoSEPKJsZnFzHbsEG56SOPXsOhVO3HdZZOSqryCA44sIVyqoqmyVZmohIq
GHrEqOP6tYY/TRnw/vzu1LhHNWqP2fLBrRudoxFvBFbMvoeyDGDfNjNv4g4k7cTaobp0RKEKOn0h
AI1G1bfxv0a1SUHbj9mpSkiJp0Ph/ngWdb+BoBYUvHBkod4KGCjlVR5jJsjNokJHDiv++fChmN2U
2zBuk1URP7v+pwLaypc1UgOiVHoWbQU2sujCJ2bS/rRv/kPdhTO5V2MWvxhswF7Oa0QBzIRpSwip
gqzuDce1urI9jqMBuvMrwxQTU2CWvkzG0kbHSw3q7CviFlZ+oFYmkun5vOqE790WliUI5pk5ZA2c
s/S5GAzzGY1lGwDDMgooh9wJccOaHcEtThakd+Sly2mJgjLMe9frjpL3lXea6FnBBkOXiIonYACn
ty6L4R/SJ0bL3pAkz8w9j17TrUTx/IDGeEk0HFH23Z+2e1cKGdQZ0EFVRgI0HGqyOtmwajbIahod
rG9CzJVtYJ9w6VO4LhyR6EXiWleKy50OCaG734XJrjjTZ+WyEKIdzIksL+FWs2YFwDP4Ib9ktQNW
Q6sYAUcp8NGjBpjgQMysRY+Vl6lUQX35ILcqIsFQsOlfAjpyri5/XLuXa5V1/sPxn6VOmjAFlZbk
F4coI3VVaxaFG8dWg5jmnj0Ta6oCnIyxV0o+M1S6w4pJ87lxIXCF+r0/YJ1bI4eHIPtXq5s2ZB5J
K8ydUiIOuwj9qIj2s3MSZ5t3btuMBjb5yIBF3CAd9hcQ2+FwlrT7j0fS2avfVIfdLR/M2W2jmh62
FnGaajbuOzR5u92Muyk+olDATEV/DKwe14/ykFzqUnyBg1ZxkzfdZ7tu+68JPDjIF5ushc9U2UgC
ckFkWzCZXWstsZl8vmi4Dq44RQDoBG3KobmkaqiREIIFJ6IF/d5VGfNVYkvOV7OYlcSUCfHZAN1F
QyzwwU1xUEKkoIvTqZOuQZ+O8Nqx1JyHEL6uLqxerDiWMgmqP7Diyc15n3E2qkhaH69oVIhsmZ8q
cBkjyLRlsbaP0ukfCmmU4kCFjjgNNbW7Hxg2an6T8oA95sM1bDwhGPLSCkZCDMiRg64CE5FzJFDg
gAXl4xajIJHg+xiQTvMicMCW7YNCVO/m54ORUlUd/5gTZr4z4DaOP1TRYsmuV2F6NYVRsNvaSJnx
2I/Foh5OlvibckHZL0bpltwWTZdkhVfj5oXXU0sIEoLpsqhsms+z0MlqW0n9qbrhdwVdrJ2uMCft
G6T2QNILJa1o0DjDw4NKaBpvzGbJxWXordxNxIqRRDlpNTn/wV5S+5yyUBnzR4tk+qb20YNsLXG7
Fn1QnSxAp6IqcfC+LUHtPwx4jQ+N3l2rR9c1PXtdJ1fGneEbwrBYubdweN3AN2NjEVACKzQy6T9g
r+XyL+w0OhCgvP2cwa2zue0Mqa2MD9d2Wb3jLgZ+vP+DODEqq3KDd9XPdpNyPuDaiFKO35HuRAL4
OpebQZhqInuJWXZtlkcgvYafui/ztB2qlZ6vlrtym8bBtgLK0CeYWBXMmyoK8nivvkjBNgEETMAR
E9/E9lKiwSwguFHDoIqde22CuqMIUv61g2zqZ+DFmoRkAUcZGQhkPU5djcYFYCCvDa16g3RBv0DK
LRlEzYGCUsZJwy0oRgs8TB/4lQD619sfkM6V4y7hBWX3ntDlLiw2Y+TmF52KEBDF0tfYHphA63vf
xtws5RaZ6siLMWBjsvwH1E0kGa8s3jKYLYMqYhLme4nLDdcErqOot/YFql/5aK332U6CeO2dQzOl
s+etpJ1u6NH+YAp6JhcvC/ed9+JIYdEZPqxl6YLSTRzp6rJywrhyq6h4Nlp6SaO3BJYtKg8SQc4H
7mkBQM+A4+1pdCw+pjg21A9N5/TdHXW5+svo9/p+Pps3RYDxNTWV8eRcJ14zNddMRdFTP6sH0Pu3
qjyalCnKnoYICXWw6ZvutR22o9W+mZ3KCsPPZCz+flFxU3YMuKQCWzEDxqohUoI8uoKIutzaL71j
JYq45Kfk6OyZUIDVbLh0u7wTYX9QAarRDCnSZVQZKjhFa/3ix1GAYRQX6ydmpxVogVK0GPq8LNL9
ADP81S4e4tWT9HHX2CTk9dwct2V47ITfhVikOO58rjVCcTkhOr6IKE05GLjauhxGyIS7poxLe/LN
1jMDFmlv1WlYMX+EvXszIRy9yKWLVDS+4cMUethAlxSxtiVrhhTD/Z/DoFx1isigU2/brZ3zjl5s
1jMl237Ltj4UjHBamd9pEuh9Ezq+dGdBWhltFYKGrk/VVPBxjU5bacGvWa8X3LjsKe6BpD7tBfnu
mLmQMuX+OUaarGq/vtHGWEhjnzpELg86YRnNpqBSpO7UIkW/Ao5n3cFxlnRFiQkDZbkGPXJJvpeT
xV2XAGRakirNG/UNDsiTtRfY/u1+UPVn5ctqT/3SZJm1uRaXZ0FpwjgC5f0THD/uZqOvu7lyUvcf
JG8+XUM0Dd5ZNc1YKY6OY6t2YdJ/4hcspok9j2y2v3BCXKMDgYkyKdYY0eXvHfluoxzJwHDqhnkd
UTH5tBO+EhLRgQ1jGcjT+yczG/tORVeC98xrJyIEhs/l6fWXPlxU4PMJ8l9IZkhn1mlhi1hmKOu0
zadXzKeqyeYKOnIlfbh+Ollkba37pWwPYX9Qhbd4/J+G+eY2STzo9MDCGqft6ffFyRt8Rbk9Rzr2
JthHnE378N4wFXmfwi5XbLkgU3dIzghilRFIkKD7hbqVSvBVcRCKsPSlhUVEK/IdHDu5BXgO37mn
zksjobu69+EzIi2dY1aJRLhXyp4EusQTGqr6WZ6GdJeAbZtExZbidKVxA0ITQ7WsL6oghgcjpzxf
ut/5s4lh2bOrEo4fp8pnNjwqIrLmPLjrAEJteEDhyJmTyL1xWLOrfFD/QLI6+680s7amYr2RpJN/
VorsPaw74JqVWocztyn7seJ+Ern357iAcUUpl5FL+jcML2YSznPaqm8pN+VQg2D5XzswYGLhDa63
tgeKE9iq51gzOpxXXQPeHfidGXsIFeDWHsucpIbWTd/EfH/0kWqhz5jj24+p25uywzl2HVuX7+Kd
zjNwag35WfuhfxS1+n4D3Dnak7ZL6L3ugeK3KT8jKPkPmAlNnNAy6jJx4ppDFETrvY1W51mcDFxo
Zwhg0+319JkGIZ9iW7W0EOyvbjZ65ce7p/SPmDUp397vsKQrdW+53OQoj8y0H3MPLdJ9KziaLxom
D1I4Tro0YVXarMfQpTNCgpTHwtZB6ga5rJmNIYSsiPLygkCEVo0HQKECsrQItwL1q6tEGpFIXrWU
IbgJ0JCYj50Zh4nhec+Ae5EFoNbT9eRENdPqaUd2W9xETAOcADOc+wBosZWCQIzvWLEcdgfT+bPR
GY/cThLjhXD5s8wruuzuNqLtYBAwKvWYlcHQfgOnSqwKHtLClI/KiN8SMKkKbJOdp43l1wFAelCj
u8J9H3n1upyQARxItvTejsuMt8b0AzJUASTlC8ELDEk0yOITwAG0F95X7UP+u1IYKEL0OEnY6mFd
5VAsh1BqPtOkvA5VxEpFm0QR2Yj+QoAUqn7gbt/osZMC/bM2j46rfkJZiojhTYehiP05fcFgfpwj
DYbnJh5rmefOHrqCS80KLHrRZIBQ5jjU0t3k5iuBJhy/X5EK9aLEfRVKbLXsvT5czNzQDc6X3D13
pJsDOlWegrAZQUnWhoZTRXVZtZD1S/LoaFShGuSnj/H1cMEoVTsID5y/dfgQF1ccjPkiLlOpDddf
Dhuv9E5FfFlJoT6ENi70g9e+9lNQUsW6ufiR039LGgmCr7Tq8lNI5nH/aYkRs5OX6Bdj2xfeAoC1
08DUceDB1zFJFK/7cVlA80rCq4FEhDrV+AGe7m8e0Rbt3Q3fivhAgsO+v+/sgfoeKqlSdX6lNbuV
4DApvZYqrOkeveDAr603pPzqq6gvkestjOoN9CPkRIQYm2y8CQtOIx//ScNcjs0xJZUDlqEvN6kH
9VV2YgFYEeP9En44ZI+MCRglpt7wAhCu6t96/5wLciZNyiZsEMQFwMQ7nQc32v+3p7hRHjYVvIbM
8D4F3Y+08Y1RelgN4+/j+d2G/3IzCu28U7nf+n4r0RBGdH84nh/YHlgerwO7pgQoHeYPN/v0MR2E
D2/xbIXzBrVHdSD0JeD0yI09f7v6sqsDPuE71E5OesWixW/c4y5SLFs2/k7j5ZsPUhYJj6xwdT2d
EyZngzsAu27SdK706SXRGQsVK/CTxVLiTkdVpqr10Mw3ghSWsh8If6PUW4aXeDrwtykCjQRoakCv
aZeWKE4k6ecvQhSGgkKbKMNbp9xfKDCuK6W8DyR+KukwTQQSvGFp52LvYAZKsYvTehJ3mC0mBVdI
aqVyyFYzBQ87DY8CIJG0ev09BoLztQiYjENR9rXRWuI+wPyZeXOAc/T+NoYTiowKCQLQGcpC7TMs
6x09PNHax9xK+Mb8dRW+CdTHbTMCjHpZgpqeF8alVEbhaXB6DuPmhc4QXYZQCphz+m5+1Xl3506B
M3Cdr6oIaXYbDEsaue81TLGdbSWh0mTFef/ViC9HRCAKHZRQBwaMIJN/5nBibWr2u5axXIJc4yGe
Fud/J+3ng67a8bK1sxQeizV6XzoNMiBCLFHCNeC6lVzRi9FtunyV94L2rbkenhMqIluJPXTx9ufj
h5l80kUHF//GUcRJOVGtbfCSzWNCt1E57vzzJ7FESzI2xqGCzti4UONLOg9mzdqXm+WqkJIKTPoo
JFO9JH7W/MoukhEh5VxRMj6bK4R3A6N/ipV9SzuZxOxMOp9l0J5q7as7bwGL46Q4JBg94VtoHPnY
U6ITnJIglt7OJJWbY2IuM+W26P5PM9D9wQ4YWPKpYLTLMvhbJbLlTIQwj4LcQKuPjcU/cfolVCud
pkQE2bvuIg59FwkiXea+tSqP/0HrWtgILHgAbUAih9T7emMx7Yro0xpkpKLfpBVMVHkcBz7loEyO
CyQLAedqoqKoJGpK5z4LHQiQ1fMw0TXiZYtcTqHjo5B0+7FfavbvjfoPc74PGzoFbqBWJMA0qTm/
8EJnCwbPzqknoBT9xlz458OnNr92zokblNIULLcCOptoYCma9vD8+iwBf3nsatJX2DR4aWnX3VVx
v8dfZXvvtoKDcwbdVEUks6UwFk4pEsrNImX6+dtnUKe3tUBpQHoJY5dL4Yi7q/YToe5Q8tBcXdqT
cYAFt3NjzaDnDXi8BOsmmxtpH+J5w561nwww2fEKzmzlLYjOo/U0d6XvySBo+P5OzKV3s0Nc07Cy
FJjsi8/sb88WleFw35lK1B5nsDYlrl+pYuoEP1uH414QfAFI+UlLs9jHNjdnUZZ0pxjDmwDUStVr
XRe3hkyu1Pb7Z2lQeeEGBYZaEP7ocBTpD7W0gGuqHkuvd9NPBCIr19vpUDpUK8b0XON4vvdiSbFf
wGWPFCuZbWB8P7mhhg/bN6QnqoGQdsvv/P6n8XKfi7p3LDTG5Q+ge55mr0c9fRCwJssSqPbrYqJ5
BCIs/dqXVzLEbSm7gn5pa6Dsbjpe4Df7goKMWBGBccc5Mj5bR33KmI1o+FJ05WF9WCQF/vORSFPm
z3Q5vg2NzIt530J3kqCB6rDB7tITzmcFnpcpHY4TzzacqTX+KT+dpg5fIEmI/vgplLacofDlUKYK
izc14wyKMp+ntceQqlrPU3ZpOx5Z9KbjpAuXAPggCaULGrOAgkm2QpLbdC7KWMtMlCOlkF1Zoe9N
Sbuv9DYeQ+9D2s9CX+8zg8GxP9rE6Ev9KOl3tOKQ6786heGo3ANc3UEnniDDt+TGPIpGWFIkn5gQ
KXi9rEl9LHuK3bPf8oPX3+wKSB2gz341lZ8O/YD7mwwMAgX510dRo+LZub3RX6GCkPqT8BmTkHNU
Xc5ko7pqEw2OsiX+hfTMz8NIzed+e/TJstR75tUACQOClKZZhDNGx6osmnwtkCo2HzOXgC+8u+uV
g7Pux3gM7x/WdCy0DFHHX85D9omU2jOKv/n4uqK+MDh3eGw4glcJxPcoIpjLjBRESkRNnGw1Zmb7
fCsgumGCE5DpDtfmjp97OWnMpV4us+AEGo9wnLXKuXYKc+3rP/jZEFDK7HzLzyfTM2Di91suHD59
yiTRweqZCjpH1QpR2odNkYO0V5IRmqI/k+2qIez4kERJajyBH9xcJM6VbADjqAyCvuAMKPLfGAmq
E+IgGG4qDmoTCcVabyfqTBcDult4TooB6O976TrqGHK0sdoIvuZjV9l4aCXRJ98KIszkFODJbhFB
yWUzW5b8qY4ZaulcjJ8FM6TZHipBuG7GtMwj3dEPHkVnU9aw4Yc+PHvcvEebLts4Pyj7DtOfRB0m
1vqod1OW1LVRf57emVp3GN/e+uy+M+UejI8Ux/v3ttXacCtcEGRCV21NAwHSurWs6fPsAk+lPjSR
sPwsr1bgzGbVSk05k1KqRwHYA4ISN2RAy172zVcaum+l84WYXWwEGxC1SzgjBIizaBQpOnUQcr2n
wIQOiH4v4hi/lS+VLbreXSBWKMO51O3r0l5NB/omqMEH5lLok/cAx2w2a+ICLGTDls2iyAYblsQE
dE7UGqGodbMV3mKHrSzsSZuoU50QLOKyDEJ5nAyo9Q86ApBWIN7EPV+7S8pH9d9KFZkAvUlMMSj/
1HnFKkWaDZOt/ixT1rWG2xkkOWJ93bFyEdF6Rs3ohmcVSVs+GSCJd7sw/ZlPYJhg83+HMWabDNb2
BFMGRu9p1Uj/OWG4WT59froM77ZPe36WppOur3O1FQtbJJKevOmhzhlE0nab9oy1wRoHc943ltFT
gBx9nY4BsC63iFJdJJ3sDBrhlH25dATzjqTW/anZ8lubWsD36ZkjtIkBXgEn4jFZxK6/MoTpxJGl
s5Yawzim2azdk8wASJv2sobb+xWED0xeATQtf01G+b/5I5CQTIEi0FivCev29f0ti65n0irWUI3I
yQNirAV8Jg2EIHXeWlyEXU0pXtD+yVc6OAtAnbSrg02U+oMEpjamDbVVsPqRZFvna8Ei53WA71vc
xEUSwC+Yd4htQ0+tgbZUxp0moISjgrgj2n9f11Ed8l7dvrZpfP78DYX5LOMGtQKHvwm6lEsNCZAm
JbAlCKdWyGq5I98dMsKE5YsQJSNBkX3i+Ov/H84taaLNwOOVFb7PUGhU6y0BlhXUyV88xYhlfbbQ
4wuR3SvUGIe5yDpAnc1JigVjg9NTtUtPkcovRBr/iseTqNKyUx1QEVLQj/1pSnEF+rhgqfzVRjV7
xbJhHqoFYNGvgoGHXkwmKM5QBNdwXmCma/fpzFA40Oh3pbusz+/Og+DOjkzIcoZfJiCzA5HcKJ+t
LhbigOkpIa5U84oYJtzigVlNCi9IPuCqKK1+ffq7vjDbgcJUfCwmGe68vd1zejleT5nD3UWwMbkd
yaxKMiPRxabqef3JJcWoUWPrw2p9xZ61Ylk7+lkrbpT4SLuR01WS4ob5NQJS7/Hjyl/Wrw/68OOf
mOVVQVg0Q5yOY19THTDkrhC3HSMxIReSm3Ho7BgQp2U9N1bRVSKaslikINTRfg0Y3otQQgAdZWao
8ewon3x8tE87KVqRGF35bTjE/99cytC6qoL4o7adbIfV1sJUPSIIY5eIGJvcoUj+sfP4gDokTZwt
fawWhiTiFlIgS8ADrzNd0XbMhcGqh1mPYuLQIIa4uYcoHjrteieSVGh8E0lVdu1hDCb5fx45bEep
bBrUjgQUgNDaYVq+bMKYxCqIYa15qoNf+W9+NkFeZSqcAzYGTLKlYHHJKhpl4XOWnBtg88+x0kow
qDfql1vGyT+Rs/KgOTqyHVJkd3NIn6l0Jajo8mpKHj2TAxaLSI4vLw1tX+s8SL+LDilkzyNMCiGU
g9njiAA9gbwxkaEv+frQPcj2HBR9Ah9C7HYGmtUyNVkXtgDdZawH1+efJTYmf2l3M3rk3m3NsQQ6
Qz8bu53svyIEF4ojtrB5dvHF9jik1i8msIXAEeYcqCHX2LVnxjtfp3uVfJLGetX/BFZiLkwc0Jhn
R8ArxF67q4V52lJlk/kprLzGHIVnNHOrosQpUhoqkRkUzqjA8UcPkErP3VxzucfBj+qp8r+8II9e
NL8XGWDkNVnbG+eP+7nVZifMYK4Wodtmy8LsduR4Br5mcRpb5EDn6W//ad7FF3dMT9DXgXzviddc
tPGV/L+P/sE5sfxltdomfvGlqdKiTLSVXdo4o3wny5/v5c6KeP242AVjlhXutQvf9nRYEeR2tFMv
/Eji0XjYqY0shDTMGtLmrN505xMU63tMTNdEjauo9vv1+7nT4DTMbCA0x0/iVx868VPQhfuxGf8F
HAv6L/gj/a4CjUtyVrcMCvEu5Tw5TtmKkhy5J4aeje2xwYeoAM4jEsA8gVlT7B4kEBYu4apqCWJF
L6BYxUg1WuDskQhvTrsT79hXmuOpTlSFx1E0tWeHDHUdyDU3VFMCDL++qCasHk2eaejvj9Z/MyYG
UxHnfdd/nUjXNP5nKrFi8VdvREB7EYHgx17DhMjFDrj+q6jA/6S1fA/oNHJZcFCEqxLcsfad9maU
Tgjr3tBQQIHvyjNCQ1c+zpAlPQavne974bqpe/GGUiW7XAokf4sLZGIKRormj3KAcludL7Aqn8w0
JF+c+Hix3g8ixjMdpDnfm1m13dmS4gZqGaZfmDRzM59Hwh+ZGKP9MmEqywRr1DxoJsAkOo3JbAtZ
KoPamnGWUKvT7AuTsYOeFHWxa1zlK5r+jv058y6Mk0zOCjEPg0jIVuT/bQffREZXX4LiCL+LUD7P
v9mQbJqJO+oOVnbaK1GhbE8vi4jd3sTlXXqlkp1jUkBgsEnX/Xun9drcFUu4zgHuwww9VvqzuEI+
pqE5GJHsXlSlHlKlFVK2bbQajPvga/mmtq20w5o6o430yr8KwDJ83y+t66BQnu+uFifmP/59yMNM
RTJ1fPLhxgh1Ebiykps3RRsAnQczITE8ZwzNoI/E3iO3A/ApABI67vk8J/d8SLTBH6c9m8geo0t+
0GIDcp7fkHSsc7rt5OeiOQfTQtI+1fS5/S3qSOpS1S7v/zvIh/Oiu5AsrT4JYg9DO0tVdUKlWuch
gQALxLMr3lHmbSt33hux4jGmkhS0fAg9Fn+HG1ZaE1IxZrBg5bJTk9k3OS2M/Wu+WvL8e1KmTlFG
H/nU6ZOE4jsKG1MeLK31sBFrgp+EzcUDnvqixn1M19ywZpzeiuRzfF1vCFdvKogTUIUeTExGp+O/
6zwE7rUqm+iEtIVUwXeGm4EQtV1qyPDI2eyVQrmKjiKOi3obOvmtWapeoHKthvEjTyWerKM8PKxw
SJVvUYSqGBodR8i7ocidasAHYMMDMJcnT/WlNWnmhSno+VPBp47zrsVXARIi3Mlhbw9FRP6+F7sB
tY0LojnMJ/X1Ajid/zkVxR9sZpmezJzSdyA1kvZbTIsVWXsgVdENeh1uI2fv8lx8dwDYINrlh292
HYCIoWV+NutwPifKaipAETLccYiWqKXOZWZhwwFfQLuxjjgMAKE0/svUkdbJx1SU5lj1L6jIF8/N
WfTl+xfcp2g0DO8VnKRDz2re4iWx8id9uYn1LccHTy5zpHzYcpXreQxYZV+8ZRosjgOrkFC4UtFP
z4M1CUFleJo9ODiEEqDyfAcJOe9SE9tqmJIJwAdHxNaCQPH9z4Aiv40GvkIz7iBLzTPYeqPVEbzA
eqeJckmb0ES7zn5brr9Yh43l/R7iqrkv4NYEuMbzwbp6OAlCRDoreUWwUs8H08cgDImclw+JnG6y
g2KklqSyoo5lAfceq8Th0Iwug9r7jGaMvPhm84NJPCfSQgbKlXMIpkCAx//R+nk+m1PeeRSp6GK/
/7tGBdM3/OQslQgClFhLWN/kac0MYMfz4Vd0NoIajlyfTGH+poM8uzTuWf4s0NYH9JKbdzOBzbej
4UvgtN5qeNsM/gvurN6eGq5pAg3DQd/+kixparDdyWUVsEa4hZK/lUGezMNE+CwA/L1S7wFgb9wv
HFbbsLLESHbSOdvC7Vu4QlRVPv1O+LlyI5DbnV0ZSwOvYBtq8hDzDd1pE0fF6wjaTyOblQHI+dyv
imRPCxpZIvhgvJk9lUugrL2vMgF51ZWqYVwfGqsru3FhBComndc3YER5rNhDwk4s/nf74wmiYRM7
k1y/uOq1kb+0AlMRRM8cpFf49eQaEDWZWoFw6WO8+QTis1P9dfKg0cJvOEnFvGZ8FakVC1Xobw/v
GvsK6n4ShqGUtBLl9mA7UueQWry1wCBRHZZKR3+hX2axwHcaUxKlHuR9jh1yv9wNyh1BkG+L+eky
tJFgSjaqxrJnJlfRsvORManXXALzBQmCBuFDzSbKxRpx/E4h5X64SP6OfyAXSWTO/3lu6G0ufsFz
Mk75oWhTNLW2ZiHV0wj59VbnE4xPtnrJLfHwCSZB0OX6cDN/w918l9U5ziZpwB0gibau92LvA7k3
RdmvIV4pAllgIsB/pnKOu7uMeRSVLINBBhwSN1Dl1E98u9BGCmk50U2K7cAE1hoHqqWRvPk/+Eyo
GAcYlCOHr98GrsuCAuzG7u4ob166JZl/3KuMGEBTMUpHreVoBwALe0i7yxLf09OTlWa5i21uFIFB
YyyPylxuZnmrwvCc0TgKClN+vrDSfEVMVGkZyQMXRcd0FdYCJrK4oVQUY7Xw7AHPo8K3XWqt9sXJ
626bgCmyaq9655LrxHJrk2pO9sk7hBjJxHrfZwl4ca/Lfpm10sk9OGff4jGHWkN/aECMACExPK8Y
nPGkVokiCSTiYonl+s3hYmp7ra+e+7hk5egZVcNUyThu1M8QD4LWCMdSx1vx737TmVjpD6pGtgio
diz5zXvX2HFaqrUNmE6/I/8ODyWO4DLiR9fl95Pm1NmZdP2V0H5ZZVAI21ohTYZFMFu8GSeAkAoT
qKzde3nPjQOivuJx6ekeXkQ0mPt5eU9ig45WLJWsSbY/6VRI6rW1I5SMVRHRI/ngr1zSf/gYKVTR
90LIeZnffQOfphPu3aueAGjmjEzW8ERGHuMxwiNhfpjaPJkr5oXHOoz6kONZQqWJaVtnKpA4CK5F
PQdfqnFbfBuPlUxqWlLCXm5joAtkLW/M5SSbN9m9Er0tbhm712ljwuBj3SZJxnRMPM0T6+rx8vyd
A/Nk8OHspXax5GaQ28+uWweE+zrcc5t7dFc6C7ZTfR8glZe+pCjgEA3TW76O0Jr4X28T4dq/oS3A
DbLhLwcyF0VpZlqMDWEe2zLaVfdePjzxp9BYsbeg88KiAWAKAaDPoSKApnLPnj4gCSAmb/9ULYLK
ga3F7LPfcABQ99d9ifRDArZfr9VyFbHDAc3+bQvhoo7bSP5vs35JLFKsekmCcQxW437/qguKBFfs
r5BE5U2IW/3K1vticd7kW5BFfoh3fsh0w/VM94+fI4lWppACtJ6Q7u8MzKc7BLnsu4kJVWtu1yZL
y0s97WhhSIDNUIkvmC0Slt2efe+Km9/9otWIl1DC/Inauk7lQl87qDuP0Xylowiij1Hwg+LNBmzP
upYbL6aPOkvvOQV/srHovmXeLUFQenQx+5j41W6kmWuwXnGSrFgWil+rHgNa3aGdgCSGNnO6KhfN
hqjx37cvDhrGRmdPe1l3MB3dM+SyWfGTsH3X6ME9p23kxmD1AQNCzmEmxJfGe3qLjOiu7+YR/7mq
xfQ7F6fywV2WjeFpZvYqIEQjVaWNEJZQpwmz7w3n6uNwMphITlsyk6IdUVsQRWU8T1M0pPPCe6t6
FCXeuyd1mShORABho2qr18S+UtaZj/c1YAIzL9/9/Ma9ESSNPGJ14q5vwMaDQ/ZhLyHqlkGI7f48
c/4CdWHVTynKdOq53K/3BoFgi/KtP7joN9K1DAw8cqzdDb5Hl+HSIfFEbGbb0lOWDJXDHmkLHCAw
sbRRLlGwxTZIdW6GQTQXI/q0Agvj4c45UlZdbaiOp3BVG7E73TAftKLC7YAB55N9a21/UA68l3Rx
SMJqOxLzyb/sQpY2+TAb+yF8jm53M61q+zhgAJhDit+J2YCXXra/zlRyGQxUNDZ0Dhbi7iS7Dq4t
CyxSNtb39HsZXP5R0Eyli2Iwf8gZWz6zrm503GMiPqNjxgzYjU40/4PhgNzJ40qyGyX7Kv3evgFm
LN83PQWsGhuHuvXKB6fyyBDp5OoaoGOe1N3EDW1oI1pghY3AQaFO8C1CMqNkgJXQOLlf5NNWD0Fr
u+CrQLnLeEVZ4MPoCcjV6XWjNjWtFOZra4E4LwECqGq6fHYoFhYGm31MWbiTWO0FqQtfC333NosH
ME3o/cdNpu+sZ74K6dGrka+Ys8eZppRjfiOOPiavVrmDXaQCRGajg8ugKmtolZ5aL4hbG/AWVjM0
8OiShYC8LuCbnI1FsRmHXpCu7+8HCJshc7LzWet3GTGuPuuR/Lv+0/N12o7SaX2RZ1rg6/FfQhWT
i2cew5bdpFMa/o88FZVFGsRdrvyjMgvup7JyAiZyJLiGI7TTjaDnaMjvZrdsvrGftvs830oENiQY
tC9FkGKskjiRmv6V8QlMlHQviIO27cziBd7+eqOCVXwoMKpbOmS0wKMqRW+jFjJUcRwwhLVvukcT
MSu6iEAW27Z5HtLg7aLa7RwjkdODcdsIasKCd/PbVBmhQCJD6k4vvv86KMOx2OH8bLh6ympBKJ8T
XWpGz4HjzGm8qONNN2NrsJYW4pXhkyVk4tZwyYnIj4uwnx1CEhmCdBHIdp2xpSEA6UzLiJXCFtYq
92gKqxgVtsbNaYuwvv/QtlULj2tTvWOmZ+8PG5lxOQAIdixoh6PAiE59qT/U8DmmlPfH/d5WeGKA
b6nA0lKFKLSpmdW1A07YYz2tl04RKbgjJhRF/QsxKqLmH5xQZGHptS2nooVLZfQZZ5rV2NsBXlCq
r28NuQirsmVB6ajp4onerZO9grD+aCeAsJGN0Pv7BG3/ChZUL0z2NG4qDJ1X+SR3HDXZhfSd6jg6
542xLXyeY6O+MhtqldDh2OG62eKsN9RS/adxIPsFz7kgylAy+Fg40laDg6ZW+NUo//nu7GfjVo1s
GkP3NtCvpquEtdfF7VxW7So+s54BKxmLYtdmRfOleedV8h+4gNzb6QWV6b+eRzS7itSNxNxvEG3S
m+tWiqTMpz7BBoneQ9f3D/VuwStrdGbc0pjLiZnYvYIemczg98OkXPkdQljOVNAoHBmxxGQ6dJOQ
oiP+vhOiD6c44MOq2mqTQGC2k2fI+zF92bpI5R23ztxc5rJ3QnTl/L3+f3/iBuJEe3fQ3rzxSb8f
Z2d8Pf4wag9+W/fxDcbqddb7AUIF7YoKbujtCIxr7el7zrEiumeyd7I9Nx6043N0DaefXLgPtsFK
kECm3eA1OOLjzGL5T3+Qi/6hSbg7yaRe799FbdSAPSRSTKtR8hwEYXjrz68v38Sn/d9t/DUtkK+p
5b6YcYjEfPEpHRl8CFeMkg0MKEoN7SZSt9k0ODEZ+t9NUHd6RoJh/cy8AUvgsYZPfPUfBkkaXQ2w
5vhhcNXqblGnwdXVudbqOd0Rr1/OKJHQHKlD/EF0Y+hRmXOwRnxI8nc7wWNx+H2oB4pX8qxYM5bW
Jwvhpy/Pz6A8ahk9eQFgNKJ8QQd4Heiufz7A8lsfloMw+mmLdm2BHjAZHOpear+Oked89DnXkh8J
9ebJkdmhMXO95ie15lbva8S8EhiPVh5t+A8A6rEPkdcCtlqg5btOHu3HhQ13GrUlXFxeD5K2mGMo
OAhe0uBk2FZDz0B6YecG2nWwVfe0f4O24y+qGLNgPrD/Cbqmg2j23PE+7aO7agb01ULSr6FaIaOi
lLm00B2lH0aVNKL48Ty+WKFCA4zzyVXtScBTXV5RejwtMinxw386i9BWNNGCyJw3ygU9R0l1qywH
7GWZLJ/E5WJqSN306oG10wgPMEkMm3dxnLsQ56oc6EjipcU5MKtrjnxg0BlOWjE0dMcENvVjWRsC
u76qbJBjVQNP+7mpv+3dTWoijF1L/LPhBRrTNoDp8bE961uwiPDmQsLjrUaMTCeQmphVRGYDZhVL
WVAkwiYnKzMfREVJN1OhzcF6G47GjSS9sQ2rozyMol3samE6jkm4JaKRxhDtHLpXnoZbUSeMhB41
OUGkq4751sxeRaY0mSyReo+dqcUjaTPcXYcDR4NPLuPDAhDff3GqKmU2ik5oFIeaiNRUcyaI7ocO
Ny68RU/TxI8QlUCTudYIVTww8WPMebQ45kQETcaEDlEFlxeW6gf7iig/OtW4UBoP+6rJt8+VAzKX
+MM1ElRNApQOxu0YYuctRgsy9WolwPdDO+zyKm554KUJB5WOo+ZZtJzGE8lzKBKYHpgJJQStS4kk
9YIU3xAPBfAQD3u6NUZz0JPu7sSquPqW5aKLsxu88tM0FBTZ9R3tkXKUCMc0RwvJxs1HW/prIWvS
HU2Lbq9IhR9Vl14R0tNQGX4lZGvjbqH5eSWJC75rLn8dq44mvSnN34x6p6QBNQuBKRUP7Cg9swu3
iB9nFVqT5pRhQAzLkhkqSOcUSDE3KEQvlO8yYc9Ig4prAzAK1pCjr79s4qIf9a5n+kUbkVPevdoB
1Dqm6K1Bcn7WYwCDylfbIEzZDoGqECUbt48prRkyjlC/Xu7T6O31YBREJjnakDcKKjIUHNjEkScx
9Sq37Ak5OkALwRKfS2A6ZyLpBd8rflgtZeiE3NiM0MO224ZVswESFfarRvN0EaWtNjPPYD8HDmPR
hzXKyQInpJ0NaKE/mnrVdGqve7ePBM9iLM9BzO6BFltC0XX9ffbT41e5d5alkFaG9R18Ju7zu3dK
zVE2xMi6Wu0id6923RGFUS0mEPzjZLvnnjXvBsa7AyIY3dbvG1oBAISOZ5MYvaBhtwXm2+IbaSIK
QmPS7MhZeYv4jwCZWPewlUrumFsCbaDmdxXlQuQJUyKXbDDpLanRAQvjaJna+3bKWYtPwXpIG7eI
h0VCDqiM4SrhUSFP+YwrkyrkqTHm/wlCu9shKzMVoddLc0lJcaejqnhY56UV5v3/q36FkNxE7u43
BHgRc9VtF/6HWRMUhw5m0MboYJirMMB+MWFeyvZzUxAZiRTw9ulufap85xJc1dqOs3rYGpdX02uM
hvNju80STk+K8Ms2FHJv7FTAKZgh6l4yY1D44SIRBk6I3iPv4XJpLfZNN3UTuY+W7sk9JyE0z6oH
zB38SzHK2YrS5mO3bVuycUBkzcqlWuGJ78j/TW3zlVf56LjmD5sC+WfPbTdIvCvgyo4gxf0YGzG8
uhr9RhzSiVF41gIs4O8bcEz3MFB+geqY3LGoQQ/CTgRTK/C1K0RuF9jYhtkVR8AN1iB/T8T8lQZX
WMIf6lK98O7gOdcfmfNFSdgdOkAI9anJHmGyfkEXiNpAkjj/nPx4X6QBM4+PYGTU6PQGclZ6OpGY
QyPKYaxWq9yiHRcNN62i39gtxf51TDsiqkYEQ3SlYwy7pAPEOJ0cBWT/RU0abqyVtbNyyQvHYDVi
HghCmOBC15cEV5+oG4s4ciJaYZ6RaR7z02iND3ADGIsCa4YztP08Xv4brs0Na9Bhn+1q28AyOses
xN+NZWCRxahEyaDhy+WFXe5l2xodrc2artg35UIXcTLUBSftbcbYVxRv+Ft4xGlAUn+XTFSrm6g9
lqR3Q/sSoXvCRpZWo7b+DOShEDz4xSP1CBhwfYEg8CwIBL8FMm2U4c20n+BgTOW5h3e1Yq6KR+5s
mzzLTfD4KyFFgpXt/Qrf//XhqsE3svvBBpemz18zGu4rv4qiiygDJO9zDxZx8qphadFGU4YPipbO
3TY6TD5cBC5RaexHnGiYNT+cDNfyRMwoJS/Xa7+YS58qHQ2VyKbE48AN957UIfNehv/hPRnVu9qH
CnOu/PAWatA7dgCRypL4XwR04fhEoNoNIuR6GbWPRlPKMr6OWr8pPkwHwJabcQAf1x3TCbFzwBI+
ojGL7ENI4T+CX8PcSVX7A1fYbi2Nvy7pzWOoBrBMMr9ysJTVUL6B7yskb0ghIFEup8xqF41/VeB8
Bz3NBiFPZqJoA9oW6j4lXu6XvLSsmPf01APaHyuICEIlYl/iYOjnXgi/xRtbmZgg3tfkxQelMl9n
caYuYQ7x7DobTAHhgAC2sWE0RNBiNVIrjHFYZp9/sKFoB6nxTWsMUyKmz2/acSDZBTpz7iLLhdbR
siTwrCI3Gd9rgSYXH0ljeHbuQrOx83Ov9XyKWdppDMaq0h4GeXYLXBwByM/tdD+9QoWNJlQUdhYk
VEqYP7uqHCn2sDln2PUWqSeocQoXYVW/QmDF6KIaSfjOfJxA5E45gNuc4tougSIHjcxHWRHtFlNU
x3yP2LAaLfOnBKXk5jzQ8zzLphHhkP8LyF65RGblpgxBFvBQH2FYYy8udamoHEhQy1sVfiJYvyzt
0hZhNO3K799KvcXV2b2aiwmJYnVC2pNNKv/NoMEFkYSDweSQe8LJri6WI0kME/SAcVbpLdg2FYjV
/FCkD7OmWa/3DEcrRWIpXlM3TcOwRPjko7N5VhmmNMN4/sVcQPKuw96dHUefrArsXH0G5AVPqyyk
8IE+Gzank6JPV7sjLCW57SV9DjWkojDDgcnMi5t/Hx+fPCqLBvgBotw3ExhY6DNSmq45EWGsJyiT
NmYRaFf2vVkXmm1/77E0Ek7V8g9JL9DaUkJ1hf8M9YP3NZxK25+PyFY3TiYM67KRJEVnJ1IIcNpR
t4nQbyQADieNlWmWKIx5OxRXHOziZtT2vJ56sIzi/gzkSM8y3a7oJWQ/yQXlwMObhFhnRHJSafFP
kpe3dl1wf1DW11gtdOmKk5H0FcfRkKcS9yDCLc/p+vwNSfSO7s0bv5jnxtf2TYo0inQ5YoR0l4vK
BcXcTCX4plrUKxhhf6kAqXJdKLwDtZw4Ysf+m4CyL2GkCrSzm0eTctyvEonqAXcI0ARq6PJajHyX
xJte+V/ekGRl+QcHeEyP4JAmRs1keQ86Uf7IvPuronQSgLosqJQfVLolBbsAs0VoBSGfS2qk75vx
PS+CTR4FDZI3IR4Hj1w8xsPunFG5Cd+jGqmv43AazEuK0nCgJ03S1o/fHh1aqvU0x4OZ4ZFf0wjh
NELFoAT4/uGfTHVvN7k1qDUjB5WxnjmO6L5iQCBaoDhmsyvKc/px4DTlPWD1Z81qiO3yvRY+zOFJ
qvkO2RhNSXH0aQjjNYh6TeTq0i23sBHQfRSrNpBS2rcOka5iVqiOGDsVyfYlYHAduULdLxyIDBi5
alVv8IPoOLNlAOP53gu3s3N1312UU0zTTdh69eH2553gQ9Mjk1dDD9EvQfnwz8FRCqqyDUAXBJVc
qauhe+jrEOb5WqJEYErlUv075geIJHUnedIJtcSq1iPhLmJNmT4wbFjGXJlvW9RHOItcmrvNis5M
zJDyIUUe1p6M86oMvLe6u14Mh6VC0Kb9x21re7iuXnKQUXIDr6ww3c4GgHzWYnjM34FEJnUPl+lS
uigxZ1s0sdg25IzQ5TS2ib+tNC8tDYMSxaDqCK8HeXKV5WNTHo5ip3aZRPHHZDzACP0jb8Y9pHKN
yZ7/1m3n8iKB5A4LIBEBpIcnxumlGZ3KjaELQARQJJb9TDmRIui1v4spy2Gjqxvbw2wUwk9+/+ye
gxpI173u1xkcW3z/ka5O5aEpSQjw8H8kcD2BprwwhLJ174iTMwUc92EexC/ktg9EJey20g71mA0i
kB3DNwy4iuamwAfBJAoo3L1PIyCf8qRi4+Ameyy47hgC7haopWku5L28em6+jfQtvwIT32zk8XnJ
10WGNDu/cTzg6DirXC2DJtsuQGT0GcC+X1fDynd7aH0np1S0REnbG6iX3V8WiLrCvzlowpz3Bwzs
nhUlxhtixDrkCyInviqVrWxNz+Y1ikc4bE5+QfMQ205eqQMbTYQ8kIyD15pJClC6Yac92IjxB2t2
fhNuOeLg3A5ypz4EEv0xgsOhZibMMmt68Vv8q3I4oMSHI1wHclA4mjHxsfCBGsq1FWCYqueKvnvi
AHh1anshFhJjQLqAPyy9Qe7f84yfmtgQusDWb1A3rOpnz7sDk2OtCrzlKDEm35N4yLnsrkJ1QoLL
lqRZ+5O2za0Rk2gn0YO9bXdRQ7GKEm26SBqY0rZgshWv0M7x2o+HYSIhe30D0xbLjDhfj+VRHkbQ
v2l9ON3QIxds3nxlcV3/n62gmJIRcm6xb90KZxkz32w/zMzrURE7fkD5viQcCvWSIykJo+BjqEgk
wzg9LTC7oNdsuEo49AUmkAtppoTdudNw1BYNCdZn2Sq5OSBn6alRP8c/tnkILJ50Rz7nfGKJ9V2H
o28KdvmxHsvHwyx315eSuChaICwNwGvlg5ftGJETbTdFPVQCd9hsyXkysaDlBcNFkhCpbNya/HKC
9/hhJnoezhVljimDLSA/XYKgCnQiuXoboeSUxLlIzKtoCcoDDqHvD15UVysGYBTjM5ficA4pSs68
FUiMn8tBpgAaV7p8Er0BFbcAGzq6dx2jComAUlEsA/QExKu4mRYjZx1BmbV5vylXeLssR7m7SDZZ
I03ZdVZuU6iY0GtcjKqlmusogucOP0GaAC6XkqkwkVKsoQExrrm+SmPoTQZhfPxQLcZl2TnHYsNc
7RanYFuYPCDJDe9E87P46qkLTSEXBoOYqcdzpYEj/Stj6IEZTEU2V20DxfSDQ+xx37mScVisRLjI
71vpEGks+oiWZeUwUN+zmPMgin/HITTvF8x0IBCGTAYdnBNo2H93Tm+Rf2cxKl8VI2QXwtU/Ookq
WOK75Y6Xb7/AWjhbB0xmgNnEES7HW6K043DVriW1JiNPI7CGEgKDRqQxbtLLtcH6cLllF7pZxhHt
ZyMZr9ay6ZG0W+MY38q/4fSYeNo++7Jraoua7InwBf/QvxPPPWKZThJW7pVp12V6+H4le0RZL3Si
ZWZsuDndzCV2/JHRtBhzpaD6wqv1sl0cC+Y2RNORBD/tRejWzCw7Ym+cQlExbiWWL7reufOLtRad
k/MEwVUfwpR80zdrMfIKFnXOyZqc+loyvUGXHyswio2j4bnFxJyyDJRqyHuFQ4lRnRDC68a4gbcX
6APwMgZH/9/XpQfaIzx1TGao3U5kdJjwqnsDkNq9uJ93e+BApp1jC96Ym+YREnAQ8q+xflKv7jhU
Cdni1R8FoKLDk9YBu0ndhX0R8Pq1XpXNBViBjtg22RCLLTaIGXDajORl1gHcMAHgjPPse6k3nS7O
dklzpXqSH+X5syfiEo5D7Ma3LdB+sUKpSefZzScbN4yi8OeYvzV9XebWiQQwsPcOHxjEC60yB3y7
6B6cBKevrf/s3o77eyoeE47kJl9G8+BNN+dADk1VRjBwh6wrH81vztW7KgWd3/GfClps2hvaZsPG
nTlrzAUc9l7b8JhGvInBgxxiisDlxCpaeyN9lqSKD+x3YW6sROAB1JIrebt60N60jlONd0elc/3e
fVL/cpKAqD414YzfSkA1T8LuEAMLU30ghsPo5zxKA8mKW/qF4EoTOo5oCVODLATDvgG7yg6atdPU
E1I+fwhjWAFzgoH1K/jcNdbPphMi/puXCp+/eGvZ+HCocbd8gJHw4TTVyuSl49PuCb0dSkZAWrI3
3PZeqvVoPLIgt0ZNgMINtaTDm7KLKuqUfUySWxuyDQXYDrEaOzQDBX/SnL5NF1WcPqNRrtcKvAag
avWj4VMYfGuxfhIk1a7hWnas80c7QeebwHmYZsC/g+PVU94FG3hu6PNu4w7eYd/pEXDNpp9L453K
bBGABCT+IhkBtJOy5DYV7qwWr4p7/lgSPSyyh3fv2OajdCfEq4NU80cjfDg2GMI+oj2UDthKfGFc
okOLek3tbnCamXIPco5VtsyErDLbaAcj/SqDTUbMWNarK5tcSaDQKXS30SRRk7M30yNET9A7y1lo
dR24cA3/RtEIeB8wNTohrRqQj17dWKgm8j+x9jVVsjr9++9T4w2BWLFkkesJiDBLsvFBzAombrt3
NnLpzsyIdXT8X6Bw6IwVCvqj9TOt41uGmAir1Vd7tmdj+CeLOVK0Q+ja35Ke9hplGr6KVl2TYnK8
tQ3yzSsWnhZyh608ECNoatRwGLZB8aJML6yUjuMN/2nHSeWqnaCzqMJAbgfK6PX46vONjuz1c5so
aqdgrY05BFCQ8sNZ6P+S5man24jRDpgEnxHS7F3Bltb3+X0UZu4GwSR8EQY6OqxCvwRNUGl683xQ
Vdo8mdjthh1LYJNdvWQf9SZil5UJjzGjH4FO1Iit0tu9REe6izrN1wr8kYxmLb58pUHOo5hXaRWR
1k7zTbMN18vjLqNcz8Z0p6r7w27flDa1FwNXTXkwY1vFizOTKGls267dFHlNW8gkLDrNuG3a128/
2DaN6moIUdlwdXCFFy6hnk59jNbbAGu5So9wMstvR3zPzeiSykC4TQDb33+2bB4PCO2fZwGlnj1N
TuFDt7j6EdnCt9aYSKNF4N8w4kNNz0pzWwt98rQXpDkAH3o6rBKqPy8qKhlk7y+j2YXtqIShW2V+
6uA9uuy25P9cCx+H8Y0ZsCrcFhlbS4zXPhXd5tSl2K17e7AkvxQZAnbSAVHdY5Zfh/+rQQUKGkUu
rHaElx6kRu2lzraSKUrT8QZB9AGv0LoyPZ9ObM+fkIoavo1+jvd0nURfk7xwbcKEu0HHERFOW5bW
0hdHHcFFZeQ5unMFtY7ia2zQ0C5PKvVsxpHbGUdjKargAw/C7PIO+pyLR4R8Vu7VZfmPKliEasHu
k0CdCJg62W1KAIEBbRKmbCRVTAxBtg+0UgfIN4C4qGX7cg7QHBWRYkIO5ULn3qHpRkGO5i949kJT
xausXaMgVxgHvgAXhStntiGBUkbUQ7UckNIdOACaPFJorDz0a8Tjp211xx9OSgckO/DP5EnJpSzC
Gn3HffnxfQJXbadAm+wHc6fRKWQcEKAi7wOYEaeYQ2iqWShFsH0eUgxv4Ni9+NVcdXsPxrVt2Fbq
v2TvEYhtx2AcJ3kfCCpwXPTj+x0qklDCUVgmdQ9VM1or245M9G8QLzNEq3wX0peyG568Vlb6Qvv6
6t/iaoGn4ANSKJSIsK85wFFqqmdH4f6cbaVGQVd9D3/M1q4vvRo+TQEwJiCIsl/l4ifX8a2UPQ6k
l1FTQ2y79nnp4pzwxzW+QxJJLcgCBw1MyT8JLFSiWDt4h/LK9+35+kie9wuKEmwnX8ARkV6liiAQ
AKvZC1G0A40UCDXoVS+yqqooN+eX8WptUmlaq9N+zXuuCgNyrqbzL13S+WDaIltmvxqWUtS/tTzG
NANCFNJkX2KhVCAyd1j+qUxStdchuIXt8om9gXzsJWe2yb1lEYOzeBxej6EP9f49hqxDLDYV7QUi
Ej1vyPBQ1AWWYyyBaaAnucWvvN7r57axQDxRPKa1EgoFGavX1C6EuK7IXGbX9ws6hWBUvU7zLjfL
+QqMuI1WDWxX3JiVs2N4Rk/ZHtTFv4d9LwTEJD4OUozR6H5XrJk2V38teTxYW1P2i5pgbxMpkO5s
Wpp5tANdb4qqYr20NMwTiQK9VDkmgY0JN9OA5sd0J1tXrQz8M6p/XoTtcneAEBEzlSulZ/WtdrQw
8eMafQGif6vcBqfiM+FoH0ONrOT6OLDtIpTse7clD9wptDrnbKDy11mG0HtdkjmjxEK/93prpbKB
62KJI4xffiDgsGwBwf5VZPC70TRQv1mB4T110ga30xDzFDp/ezO9kFutfWwd+aalhYU21zXbOLwe
Muiez55kVETRYWf2MjwTOEUBDbFZXczrUkRK8TrbDla0CdHFsVK3RSy1ifSrnZXJdg5Brk7x/7Hq
K+Ik7MOc8AWfi63A/Kax2hd6h+CWxTepq1ioHbqwYjaNx0/1lAmfPGJssAUrgwl5RLT39SgOOpOO
sKj/BPtaQXbRPoL922xtw5+t8KObD3FHnSTZqGqvkL7HDm8PkUcRM0HCfa6JNBSkQd/ERT+28PrU
lxHsJdMESwT2/MZ/uLXuZVmOrWRco9aHXPV9zK9c10pUKkdZwcoD17+limW9Baszor6ACyUOlEAx
1zNce2OS3aJtCit4o47wUltQlqPjhE3M/9S2f4w2Yg/uJXtUL1KhKsNe+0LlGsWx6zbFct20RPC6
btx73ax6PARdsZ5mftc5VpsyMLIzSaoZPqNHGcF3CmDexz1CjVlvyuwEjOX3RwUMMpJDutL2OWM6
r2mt2br7VMIcHNqGCSd/yms59GSUmRAoLZVXASAagi4fItiIpCtl0U6wBfJA4w//+6f8IZ/QP2If
K9A5fg7lY4QN6qdKdwRCK3btLGkA7AcW3N0mcxZh0Yj8qTyxQ+kC7gdVkeUMWluKHpfuv6mtpyVw
f8HP9pmgwNTRWl1dqP1nLYjABmHeXHsxAv69ODDpghQpIXmf9k+VWJ0dDLv3NTdnMAMULc9Fb7Qw
t+1K9FGeViyif6P5BGLiN1bdMf3+m+uIOTle2exUr6+0krG58eYUGzjlO3kuRJ+rwrgTFp74QxmV
SR4BMgrISp74y1/r2C7/LceNGfwajWClAAf4kcI5WoAIHFJ7Qox32M569ggzk9eqpirSNWHFb6g5
1XVxGj8OdISWy10DYLfHai6WDKxRKIEJYk3KGV7OFZ0cFWLzzLatrzSh2Pe1VhiJbg9ISmUH/7Lu
u+h7u8eYfOVWH7tdKUhinw4jZk0+3CJGAO/aK5O+e7bfmZ2tQzmJhMpV//IO3ufpxObyVpVPWPfF
H3j4/1D6n2z5KgTWIYXxkvcv2EJPzx5Tn1HHL4N/CWb8nQ35SIehmHgzEX5nBhuNOectMVshZuUq
UeCIuMempnJPQws/xFrcd5u3GDdgmdy18vJli4VqHFkFL3A2HdddkgUqk9iRotzFBOsc06/msHHA
Q9SQnX8zsYr68ri59MiTHWKGaHK27jvJrLiyGrA0vyyuYaelUfMCevU89S98Cc+0DDy9lHkA0vHn
cOWIoPEL9ZrI85wFhWZJvNi/EjwnJVyk/0MC4heabU+q53I3VT6AGdL5QAapW/ozOQGE+BqwhNfp
3dDWU2pmPYT1Ua/7ws3Kh41nCBH696mXmC+fhkUMJ16p4QT6OCS2bUrkSsdJVdMkPl2aD9G2pkfE
lLau5bSDuhDLuEXAlmLoq92/GvRhtkFdTsbf1GebOqm/bfbD5DzGD3E5APSPKYpUsIQu2/o+14Ng
aYpmeEHyW4w3iatgOEDRVN0pIpWO6BLkStrtBupUDmx3ZjotgILgLfxglBahPyOGctT91Q9Ay8Ym
ckWYjNB5yleEzLd25cyAo/n/l8IT/oBSLuWA8wGPa8s+IIPE5jTMZFlTayqvfwMQrRQwcHNjijDC
zcbwt8RfaOEnNH+ZleJb/Z0f5SVQOQFv9f3AzKYwt3TrpRcfZB7o0GsU42dWEPhJo7fmRxpsTUVL
JFXLCs0ZVT3GHFHDBVQXF5UQperJLjHcHM5ERqzk8xjsfiju75IEIAlmd/tPqvZXmrsGJL2Iz3Kh
DC5U8eTpeW+9bMwnXLUYcWuVvtNAZ0vra8Xo/afh7LoekHuH9rK3MzCT2XorAEpLUSr6rgX8vvek
SqUxj4qplpp/93pFQEg6l2aDDEqVYZSAOA4opwiUcGEyKqgewTYrhOip1LTAryqc22+D8+I2lr+m
z40Uv1NXvG/sTTueVGaWtq4GyOWE65v2a6thkqNXX+txx+SDNmlu3CgfgLe8R0JKj0vJTEpBnDtC
73xv5VpZxdoWiVc9jDbQBgTeREBn43GRTeY40juvaptj5BPuE1TPooPJLiuVDDAOP4KXoHWkraxi
qn8RKZGi2U8vJ3K/MjKAfWjAT5i6LaXKyaDT4s9eyCcLN2N5fj4CaxUBWys5QRbki6xrj/jr3u5R
y852KBMzEKG7u5XVVMO1KEZnaUXU2mDMd7nvlZ0rK84jTltVTYxA94vouHmN+VLZN2LG/C2p/z8c
MtwWEBi6/EXjUzd0E0zMRvP8eVHok7sjSRm75jRy+gg1HnUrqOqGgGpJUHoz70NZo0AiNxlHjqUC
FhjNV0TmDC2MxTeri+7dMtcdFvKZvMQ1q9Y8hA1BbPTJQcZ9Mo3zWGDiSdLFQAYrbyYHvLGyZWaw
m3Dt2/v0QRwRHgQIWOF7WIRchxenchCXEe0X94mdR8DP9e7PRyh8lixiGyKWbfIhJkDfa6KPGOGN
4LvPD4nHlCRnGGk+K4DgYGUqJLuwhrqApJ5sPRAMxJnStfoRaXn+C5MEpuyZ57jCYY4avO3cXk1+
TBy+S7/lvL+x1o4KuMmUwbXDRrAmhZqr7qa3FQ+X9PnzuiQyquR3aCOnOLAa/6enMJp8iDXfVi1m
eKMbosVXZ2kUc3FsZ6ps6NO+31pJXj8Ayj+F9eKKTEk+CPXFB0M7Mex9d0gUHLrJ1VoH2qF6kZz6
23EI/deOrkq+/aQN6GkLOzHFjVE1Wwlo5w9htuKnWIe+FTdgZtmYMEtlf3tl1NdlBC85NldXSK5w
tf0lw9zrMzcG4wial0u5+GRKTzyXNMhRqBL32G4W1ur0d1aR6NEfLIheBVR/6ZdPLUYLtbijX2Pg
EcTCdou58zHWOmTrD6v977zX+Wc7o5jExcU9wSkW2u2V5pP4cKopAzUj20tnlqXrnc1YoUWANKK0
6v91gIwINzozbCC/NI1tgh143tk5PX3AO95EHTaLe2cHHl1hNwnLJXneQ/oh8Iulo6lQCQApK7RV
6Etg+DNJFX0D19f0q2/MeWE2kNMHVA5JphCtcyslvCmN/YMXGaH0D7XXzTzo+DiiSVH9xT5Ls9pe
MPRozwGhTqs0/rTYYa5YAXj9OqU2fh2rjLmRgIUTxo88EqP+GXslW3bLHxC7VE3i91s2CRK/pYMF
NIBIyGGd1KCJWTtAedrOhbMHdHfilgh15fsEJXmNwuNrUYZ44ufdTKpfoCxceq15TUnXvwqHXPLg
9E7jFKwTS0yzK6xDyM6+/MObwkFx8FyPtNXqbD3jBsVEg5WTwcP6rYupeCo7+Bkj38E3OlZLy010
Hp/9B3GMBFxSf7gtrSlLJkD931WPcrLIneCEbG3QfbCusSLVWTKrh+NTp7U4pL0OscMK44r3XFl4
QOeZ8TwubEMJLmFy00l6pp0pQlEvAw5f03gk8h8DQN14EiWppx0mJPihNR2JlNFlCZDLGS5hhjvs
jv5s43aoLTRJLhAf0OBmVdsoHALYJNLuzZW93vkqiIDhwbHXa83Izi4hApJ7x7J0L+jg13jqbBW9
Bznv/AaQtUBxIQGRsZrlSRIlTn9R4cdKG62GBuAJW4hi0tUkxel49oqdcb+5mtFqzTzVCQtm3b8p
WGvaRbw3xvnbzj3T0Jm2c7SKodyF4bE8btQ2sSYcWyrrvzCeQEAadG2IkTL/mvIi9ohkFjNbSPhl
ZkZm/mGMKt4V5wiyTDDbgK4E0vo0TXBluK2L19iN5W0QhQ0zOGchWQyt3jhDa5Fu9wUKhGfceQuo
4tsZGk+wNaBOx9wpkfBKv0DV/cGVpfmrmqG/uyKeGl3CDNOzi+zgy/Yqp1qp6sfIFApnFo6hdOfs
NVYVW7mkGYoy5EzQ3B9PX7OAO9xMk0/8gGkJO2E4d70wVAKdWJHB0BJoL4uKPnkCQzyCwNkyHTin
EkmyjOHq5Im/H5q3CBMRGNQ/Fmi4uVu3SbaIyvInlyrSV01G+Ga08q1Qy7YKX7Cof1DkUQMgclvx
D5qv3mSKdr2hxXGQWPAoUoyLHg0c1sfrrK3z9SyRzVeqKQx2ef5OqH3fULa1s2Ia0MzUcBd8A+n7
fMnSwKVQZ9f5r9h9QoUFgwkzN2cujTi5DQkJXmMM+OLHD5WOwggZtC7FPD3DAGh8iNhzWpLxQ9Sn
En9yLvy8hMsVFY+2pkPgPSiTdMeNXZaZCb56gtozjlMPqazhlwyaQsLgnpp2hr20uBRTj8VKet6r
IbP9DpfH8FJk9LVkZiM9ZIN87C1Jny6R55Bggf7jMGkShznmRUS+TADUagU04JkUAlIz5g+zQvpc
OA+EIQD86KRlLkg9YXK0B4T26IhltR9urL+iuJj8kI68YgPyF92INIpsd411cpgAwP55dmOEgZz+
O1Ld5V/QynZS7PC/lGLt8X1X8KfJt9pMi9hZL5cJ6zwRl8s5N91Vk5FzvdAJmqKOzikwxQb/v59a
9gDb62yH3z3vuIytG8qL/T+KEIHjpkeFCWerGML8oI88M+z9Ktc15s46p42TvgDgCuuYseGF8HCu
jqBk8rtq7tIvKrWHglXzKFtYFRsOOTDWqSx9GpF5YCCrlWyoCHobH3lrB+WDKs/LM2u9SdaY0wpu
mQgmw/9VkIXFrRi5amTRQmtl/JBUdlQwrP+uHut/+vaeP9DJ/dYxk7FWohW9edtM3QqWDSvMaa3W
QEHFgoW5a1SQNYSRRbarw1BymOlDjR46hklDy3pEtkkeFdt/s0NY/bTp/nMCe4Jac0tCkgKc5GgH
j54GV4uIjOGdM6wFHooL5tYhDctNHaLd9nfW8EE3D4I8OADXFoEtVhyAdNa8fO9W6DaviANtOXt2
2KTSdnUCLX7xKdyLCA5bv0Takp+jj/MKsPpltPcKpBd5SQ/8KHulo3lZR6UEz6BSibPBU+bXp8Ri
RCJDXO8n+veXuiJ0aaCIsrsCQVyZVbZTJO5MdZRnuWgknQC+OkDPvWYbpug3L7sRjuGyBtaFIcyz
4OCITIWJAkp47PdRxbZWZtFz5+w9d1bdRvgD1r0QCAY8ykYL0TqEbNUkdT4lmWrdhgqY0N5HlFdD
HAu9hdvEL8v/YL068o0+BhVFU3mUBvUAaGWc2628WE5Ce+I+rZAGf8wK59DzL/el23LJK0E4e1k9
T4k8EEhQIkw8AgtEkRExvDB/71Vnf9wFBUufZDBZ9yhrkpk1rUXyX0p5qhN4w9rmfO/k0fL5Mg3D
MBiKaI05mwBkmd6nuLxjmwEaTWxidTSr/lcRIOM/wvud5xtVuGYJRN/Qtz+Hq74bPMphvAtaALnp
VE9F40rj5h4IuBW8Aiq5dgs3shkLuZmdM4pxONc/isqdHwUXXDioL8I2VMzjusqYq5y3795tw2qJ
Otf0hrW7DQL0EeVQBS2SCiZg9spxbVewfVQVUWV9/qL2wMMpXTr/KbJ45H04PNlc9597mYB75Wom
9/6Y5DqEjD6SLfTz7NlIQz4ZUzughQYNpKzmIeQgpHq4s6KSBOd5qsxDp0tNWNBEx7sRfmlgfyZp
Uf0MR/xUehYTlQh9mGrvdS90kjiP62VZKKUs6qAlXzs/+F8X0tMUt0Pr3NmHpauHMYHZeQEW0grH
1VCRKGXHrunB/K0sxWhGJpQvx+FGZhiOi3z8lI/fDZLqNa1fBb6ZJrX7VNkRPhH8KTesleGMZDUl
C57IEfmg+AImV8UfMk4y+noOsYRD8BJZoOCVWjSnMkdqzQdfEHU/RodxoG2F2m1dD32qqmRYME7T
2KObtwgvpLBgbJ2A9ENngnJOkin6wZklJbhDefXUwjJwi92QA5paBACEgT6IrMCe6PKvcN6zPMAk
iYE3Ql+lPGrWslgm9HVtZgXx4yxh+RIz/goxl2TetZdZ0CNr1Nw1lMspyFCLPc8cl+4ib9+YL2aE
5OP3EvUEsuwoJvnkppkg9+NVONRh8Z+AH0V2I/7EGz9mRN54eMXsstBAf5cTwzzMZ/9ogPGk1ilR
riAaoajVjQDMsKnIqNkCbNqAYNzByvnWsUDpp1KMVGe4XW/CjSmtj0XWeWvogDE00190HkaPlVhj
tquCewpYXGi3kMqQ5rIoQHv6tUW3MUIIXN6vuT43gFeBv79bnXUdlwniX/lBCSyNjscjrCD2NuaG
dxf3a9qdbCx0nros9aOVzS5xspELnC9lq/DVyFN1yLs1/jFpSVbCv8gKe9ILFD+yEJoihlHTEGR4
1jbsIq/PyNxzw1LaU+K8Fi/lIx51YDY285imBtD0+e7ncTibwSFY8dHcoZRuai5ATm0pdXAzpKf+
2+i40fJT/Of9K8WgXlKAnP3NBl4SMH4k01lxMSPUNY3NWfGqygP8LjE0UxAoSX1ahmhdlwXF78kj
j0XiqT3//9I8RcRz5V8RIswNlpYwMTY7Cp/QDgFE9sWH3oY35ulg9XgEr54WPUuQULH7Sajj2ZtE
AKlPVcvtOVHb8kGOB3UR1KBUWY3lczsIfAbtAh3tGuBQrU+EQNeuewDyCk1ZogDaPvNsl6gWDyKQ
m0rhdZWMbwV4A9mxkFCzoa94UKHVGxNj2dsk+WturIhlu14CBsEujM3DvP6EgxcdOkDFi6UtEeOT
NAYn/bZrEClIrxhDcFHxUpdkZ/gb+YpmIG0zib3d++TXJyVlPeCb/IdIeI3VUasY6LM1yQzd/snA
iiPRkX2w4dCyhFB+JOls/1hC97+7lqDhaKQEmwBVxuPoyAuSFeUZ+z+9CDevICtM547w/GnfWekK
koPwyrNZ16W1mojqQdg5PAPRxKDswYnZoGHQez1aOP4Tbz2bD7Uc6wEYUQwJGq9BLdB84SQXzdWk
ZBwQkphjridygCgFYj1wTXlqA2Nuf+6EO06Bh9pq1gNrkGyqI+jZIohTPk+4fH6PZzbHQktKMnL9
Y/WVGmbzNzk2jpksySE4xq8xt4CdcomszbsXCVOCe2mw0JJKfASFO9xyopVCdIH5m057D/bkB9NR
5Bhgv/x5xHbfrABKqCgVR4/XWjeTd7hyb8RJVOzSSw6/Hb4ZYSA1r/EoGBz+sbxL57btNdJgZ+Kq
Ij9OMiaN23RfMOjY62l4FSEGYgTWG4fR57qzQSMHBVvIRJGekMeUfWn4zECbrqcERO6XkU2fsI5n
sR4FnKz3J2j2eeKldilvXsdfZZXWIhj8MlrDlT6A3nNA8tnLUFzJToNRGAGFZBY/r1q4t0nQGIv+
RMbJ1vA9Is6VqrEhJN24w3eESyYe5c6FsrlJ+o+oe6Cl5foOsvE+5c6Adcp+UaiN8jbIGRxqo4iK
jWBSqMPzdx3LAWxgqPQZNgGXJnISsXeWrfhgj9WkEj5m/by7FhB/V495GCkEj2lOpfmu6kWsUj2h
RbB12vJT/E3f07fzUeK8krW7KFQKLFfhBiYE3e2MYWAhj2fUg3Lv1Oe0KrtvxFmgj+w4WAl9zlNE
RC0jIEvg706aknR/9+9cC160Zi6K7EF7Mmk8bkBi2BDa0R39XPagGNJxSMqdTDRQeONp1rTTfPVx
RpCRYLQJ+iLpFmi1OW9R4LhAJldvWyi2r1zQeH/btboaGA7iMWr5HyZGs39/d7D6AgK0N7U9bYJ0
lH1BfP1/MesbnJqktaw1CMQKl44HM/edmHN5cqlH7xwKUzoiQB5a3juCvSbEt9mTz+tZ/h7vV8fw
XQe8GGxyfcPFcT7lJRJdh+hG/mGOaJ6JdVLlWQ95wYHcBKQSmZvRUpXo8wFFsNIDT9KHyBo/pxS3
o//8uHDKWL2vQAVJvvBn6sz3Vohbd94UoQHR9570DlQSj14vzQlSL5igujR79oLYaxINdKjjBumJ
Qo4jbsfnUN06TB2o7v75YmRuc9u/hdBEO3NNQHL2NF4Nvhm6+Iss6lGtVbsXQcM7LscYJqqo/vUw
XI1yUpgf/eqNc0ljlSJ6OB03wF22oN+ZYOvPbH9HCdJh/g6TTC8bw9H6Vtqxvf1JAxrbuad4wW76
BiJrdo4h+9tU1KYU78GXphv2XTG85uRaqDTsqL0mBondPgt6tC+quyusrX+0tDAp+xhPzf9WrijI
l/4HNfcNKtyGNNrtNp7AmPoaeuRUS0Vf6KQ8jHHF1Ut4u4Lf4OmeDcwJenjyT3pIpbEgwangL3Aq
rxQc5QmtWSkawS8r1rLzSfBpY8yjCLkk3H3qfiPngVEuVl4ClPFOX7gzNzCfsuoLrByCdO0aFgmL
MhJq+wKArfQ1/opmqQqzsIsUXCRdSK4g3YXx7HauCUBlgBJTDqeY0dRLiI/xRXMc4gBkr6919Om4
DhbjY2hPiaCLE+AV13RncEAubhYWTs4veJsXMlu9JTCIYQ3RUczJ3d8X5vaZ0fhFfSRPoIL6gCc9
skiPzO8GocFcqfxYDZUpKE1J9xBkdMP93GSY/LPWEprJPVyYfdEHAviZ01vhMoHocHxsIjA60slo
seSaL6LZniLx/Mj1Dwm2jw5QIWYgcV04GThyfp6I8rN07c6j3ai2tLZ0gkk9s4pwXvAgYqvG3gih
R8JfAjeFLcILyuOoi7+Ev5lJZO9rhiiJExB16aCIscSw5LEv3ZmmMULTtl61SFRcp71xtmbhnGlh
3sVf5FUrelvuHMHZIbsYNBIbnTnLYHLrm11KqDg4cgcGkELfGN1MWzq45nDoWa7P1liCerfykGw5
8W3ovY0GuUBBrrssdUAdDL95bZaH1Qti1vhlhAvX7mUJdtRS0yU3Vg45pTHPEJ8Nmi38180sA1i4
Z5+lzOZmLH/7fx2UpqINLA9E1eaQs6IJEjRij3jYUzrHllkIQPTh3oNxN++2lIqUTLzahKsqCIpP
ggBw+zyFYiAYuMBriZzs5QcTu6tpqDq3lNX7CNVb8m3fvJh3rHE9r1HeOM9yXnNJ8Lei4hXhjDji
v6iaemdodNNgw9voHNPqljo9M5eBgshkOHo2OuOcubfEBzswnWwQHMB/uBiCBpGVPqYXvTwN4Hx0
oyEPbP7BnxixwdIx/Jcjt/PNe8zWV/mgPMUbqfoE5r4i5IuC2lY1G+/wLVOpYQyzzXfF0svLUfom
Gcmec6UG/4ocaA6uvSiSEELQjGzmPmPqp4QqqV3ksODiTEtr+v7vd4PWL0cawWhxN1g6m27hQC3l
68MtWLN96TASjCHl1Iq2zfMpsCqxsSLhlzuJRi41A7E/mwdY/KkAxZwDH0qvox744XJPMuR72Cpj
jlaF0eSln1hnTpj2PGrHOrx/uBhFaEPs6BRiWjP6oiJOpkQ2Ap3g+IEqphPCjwn+mnKFdT50Hpgq
2//cFS3Rx7IhPP3dDeMm6b8KJ2KN/rHL3RkkoBJkclX4CC8vu8w8dCN+u0GeIs3Y/t90YhKJI2eX
wsQV55z3+Yo3Zx21ECuaNCxCmLaGq6hnbE+wiUaZvfS/oFyEFN1ehFEg7nZkW/IW4J2fqaSErGwG
z9R6hnhL+t/eLRZ/IADll0JO2r/ah1KTuwQPz8S5ldanPUFEbUVJYoibvNys95A4XHwJWJEPVHdb
od1GsD/IO8t9OoFGWnH+uP6PUUluB26m7H4oKBEDrcSYeW3LUTLkYJ8A9JAxRMG5CMVawG2PmZyr
olcWyygavyw+E84EBNHTSuqyJzk50EpuVfGnIA4392y+udv3c/xE149/JeFNa45vUEeTfnJ7KHDV
q7pMvcD7bDvRxWDIM99hSrX/DD/E390HYy3Z4jqxgwNa/+XgyRAzyc47lZuXYoDzzKrh5nIkwSUp
JA2mEqW2mNH7Heer/W55tTkgoNZYPSgL/4fkaNR3qEaNgS8/pbC7RJnG30ti2BPi7KQBAEEBHLf8
v/8fq4+G26sJ/nBWOqWLTEcgoDQFMnyok+5jVOMVW8rPgQCqhST/euCYtw875jNiYJcs0VH+qXKD
cZquMbsKNw5gff/MJUdwCGHEVB7z2QI5L71KaGDMhQDNjPTk+WUUA+a3nBNKETh8Hqub1C6J+AAj
NT2eY1xNxBjrozuwGkPwJAExLZgDSrbwd90RoaVq7p4QRzrtnoGNNJCMFSAX4B2Ys8HvrcDAPApf
ilvZ+ndXkeYMQIqmx3S2zHELNGAx2L7zINqJGYv2kSMDFf2GeoCshGSF30+731fJ5+SqcapPD0Zk
xop8bwrsZoJLHNRH+8RSktzZ21TyLYEPFTu0FbxT+H5G7TBF07FrqQ2QW6hHC+lvOcl1KoDERlnT
SnM8FIN/kzPpj2jJ0m8VuQvzVTZw9wg03NgAgcfFGb5FV4dNb6mLjbfJiv5EdplkbwZy8oda0mXc
ZGYgRveNf8Gur4sirez+iDbVV0zeUDiPX24FHZEAjQACkUhNabtEbivXL4cESrXelPpP0SkaOVWM
tQZvAAggplkP+SZeqydbG0Tv75AfVZ2icrAvMwJCeBV9jxKNfIw9clHnp6RyvZDZhMnRbd/4KLcm
B0YhkdXU4kgaGSFDKtRFoJA38o7WUhAREDhnJMFt3Fs57Lj/3fYSc2ClGLJnyyJqSgYu4mGBAenR
vdWFh1pB4jeFvlYXaJbbqjW3ZFuKcGQBP0BkPuLz1S33cu31P6LE0sevahurs+Bx19iWexi7YuyP
E0ooVps/QQXjBmzckRNwr70HleUAGqyFJkwY9skJ2Y9lroW1iURNFGalRE8n8IJ+QbwDS9zasXL2
unABtdNqdabf+rOtdjNo9nc0yiD3GvoPd2bGsKlnu+FO+q8lFAir+TvRk0fFNtOmwDKhWNpsIk5c
f5lIvaSkP3H3ocTnFGltP2VLTP9y8ByZxx2eThJElAI5TjwAVqQ9yF6tPG9SpkiU7c4jxDLMNq+P
sY5Ov5sWyem0KHO1/0Ab/8FaSXIRd8/vEFVv+mlNrG9fuiopkj0Gr+WUwlmvkzpTllzkoixdehk1
NEvQdadA6jVT+CzazD6jGYcm0Y1VhhsIdjdflMS34Tl/1CoEPK+TJokoj95L9e2c0hCZOKSC1Gjn
b/5DVjXdyPBidJL8lFM0+q+1zgOJaNwsaBATgTpLa9ml+WlGAxhyQYpU0oQSsrccJxwBIoVl2bZ4
KM/hcnYMElwlDRPCi8s6q3RE2sAvcLB8zb7pEFafIlAqotMfvm9ONL1irV/fwiK97n4EFUQfzD2f
WBldM5qwqWRqXE/ZsEIR1OJy87TXr0VV/XgJML635mcs1tRlChTIVUCb3xBqnQUTRQKJtEIcn3hh
tHVjEA4VtYmlecL0B+Mcq4ZHQHGCK3CDGSRpzNgwawdbHZuqrM2cIMskn2xFFlPUtJtucok6iH3X
dG4H3SQLQ7sSk9AySpwWLyBF2qSk/EKkR9qa+fZmZlL733YGgbPzg3M3TnnkYhK9By36CUKjEj4r
H2nCYmMvMfXRA0nv5yXOdQi1RteNVrlwAAlBhcDo9ZTL49q4lRb7mgGwg419mXl/QeyrVPE6YfCJ
X6njRs70FJMux7/i2bn2A3M8pfe88o0FY9ROEuIWn5TUpokwlF/ZDWKpwIbV6t/SnwKF20eK3UQB
SSz9zo6EHU0iVZRbz0eGghpTnvfLxrevRIvUARLnLMhm5DRdyZEl2yHlbqjn/KBNZZbhiMTSm1w3
0bk92UriyzYFaP1bm+ulk9LqlJY94d/vQsEnie3+2dvDjFQKKnpqpp9JFQzN+v/AAIHVO8CDGI3l
g8m+bcqPZX8U1v515GrG+HP/G7mI8Di45UvVOYLfvVqI6AsBJxuW0AYD3WCBWCXugAH2ntjPiiVx
+8GNqyp1OcpXx7jY4sKzmQ5GmFK7Vv5gTVRJR3S4+Vwg3aUF9IJKs8miSy1F/KMiyKZ/T3LtUe0H
S1fgpwRV/yseEnqPi+/X9ArJ9u2a/Vo8+Wj7o51QNY0bJMrkm72ObZyYZJvUjHr+Nx2Vuk0euTu1
j6b0J9G/2NzlxqLQbWo+ra44kEv9sigDbwMBa8UQeuSYMiIIyt9Yy138a/4zrr47K2MLt3MMM2/Q
ACkbwdiK1MkxKf1Q+pMVhOb+6cXAdPjS/0ODW2D1vZljdecOE4vQcp3HmKg6Pz8BJfVif5mtQCWp
RSHcEbMXUaJX2lELQ06VcWWCGRBCn7yPEvGM0LPRb4CyLTEcTCZa9t4h3O/t3YQTZH72P3KEYnL8
QV6yjOn22t4ohlHsiIM8bEMtPaslpRxAIl2KxyvVAxglUWf9F6svZw/GkgcHKZ0UMAgYqrTkvVs3
zYokrxEzGeOdLYrwDx7yZ8xpxyKwucgomqj23ov+bI7lVYmu9JmDcCvSJK9/Cf9WNeNaqCSdAryU
3IKGdhIoFxy200K1MZfamVK170Zyvw+vVbm6VqiAV7+bjUxrkcrvyRSM7R9iS6CPFmjDdD06TzVy
+8YUjdkntQ8Z83kx1OiIaZsnn4NINmPPatHnQAZoFXAQt5VpOv4a+tQlfngCOqgTSH+2olD5FLXe
0hEwaiz2yymfcM5fNAJT/QRDngP2YHaALS42CotBlM9kR0B1ntrcPaelHgLQvDlebHTtbu3e0y8N
PV49ZuwW+obzfyX+RTqdTPuCbaisk07+uQH3zo5ysd0VqqzCbgNyOd5zNsOgxDGHvnUuoSubYi5r
mFGVDRQNGlM+Q9OSD21TqutOLSgSQEQRLlLYjO9Z4q0u1ujStLflLyh/5Tf472JJC4p6a0jYVbd1
f5X8zUck4vfGmB4ug1LEB2bwn2MkWsoqE7UT3c87F78Bn6MS4j58usdK4SlgzzZklw0HxpmRO0ql
Jtw8AtJ66V3ERHVW+cpOYJPtj7v1MdjY4niEYbPmAohJiu3tnXQfTXglU5osxp+5b5Ymo4sovrQb
3t8T6uAz1fFRa5t9COFovFbIq72a0m0SSwH2vhJUszf8khNLzyjur2+S85WnOkdW6Ac5mTuwqiUX
NFz9rNqEpKMrAo4EhkP7ZxOsMPuRDmtgQtKLUolF0nfOGtr45QE5h1RhYAHy7cVnOy6jnrq+ujNM
5pg6GFxweYZ4G4IqwfCOjmCFtsJ0AM+yw6Y+mqg0rI7f3kTkSVrlM0mgiX2KAZRzH/UHUUvQwhMy
dh6fu5OMhxLx6T6+pb/z9DVukdWbMO6fd0DtuieDlX+zaitK1C0BjkXRPiFKVNX/8//RxdNRrAp7
ul25W7z0xPBfmAPrEVX9MUjB71Fdi9EN4rZ9QRXk3TcmOEXai95yW7taK7gDJCKIrAPnZwTlwLCn
/P3twfH/i3xny/qaC54MKwwsrWKK5jFg43QI3HCtJ6KaqluV2CsscL3e4jr7T7rv+H8H9stwRMBj
ZMyI6C1gLFKKnpbYKLmjJEU1siYo1IZOdai/qCAuLCJ3RKTdlk7sN98v83Egw/hZfpJ/XPGZ+UW7
e5iZuWIW1sfBtyb02Yp+wFRscTKrePYnymm1sVL6eTc+2zMslZpkU7pqIrzf4Ogl2ISRSbJsSSzg
P1ZsbBxA2LO6JqEpxnGQIt6I0c1J9gQR3hpMKqMtjK8FbY/ijpQ1qZsTCPwb3XxIILLCvS1iwOa2
dPJUNAkUuHgSaxJerOqKkXTHzVb3ZAj8CuhJSN6s68Zy+7Zkr6G4Mw6f1ldN8roLzVJS4uXFnrdD
5lKrcAEoWBkjWnD7ykw90Jhyxd5yU6PsK3XiErnFErnPWmxopuur4HZ1vHtiO+aoaTqk3DLYF+NA
BQA5n4HZdEwIBDA3ICK6ZD+N/0aVMPiEdcLKts0R3tPJF7mPoQEKDkhd7VeZvkt4+uhirc2W1Njh
w6+2zkBtprJAVKUwv80u2O/ciwEkTmzZp4d6Mq23yh6bo9cA6TNsIGjMqQr2aR4+PcQO/EiivMjd
ImzbCaxZM1NiS+yyRwOylWPIEZRPyVdbiupXVNwzukooDYKmRUB/eu5xIeavJ+L5OyvYrXluTMfm
FPWnl83ed//SIQyJ91rcnfdUhytmQy34/1Hv6/XQwVgOmTmc/HUlz9yeml9pkVnjDKEwKe8WZUhn
8CQTYh0KaBQf+Uvi8yzAR8gZfw9sr0MgSb3Jq3cjQyvMRPcfxZ7kSHQYcYDHR4A1D1l7ANNKIva+
uRLtwbFgAftRUXoKZcT9kGoeCAUnRqK3YAl5MiSHuodOKSvfYSUzlvogwcYSSRLSd05AMvIeJMLL
ztjhzHkv4V0KMOcF9OSPTvQ1EwF8bx40uCo04DsytoSs5v7dKGYqWmAVPrLMiED4HGmP3u2g6LZ2
NIkaPagOr++yrjfgXIEptKYO2NhB6VrnN/GdWcCZdyVmYLinFDz+LVqlCCCpbEkDz4zREu7K0GA1
fXbV2160zycQ7BeMw3zsreAHNhEROsXqzmvdoZhLZO8pQniN4hYWwBlsCHrNmoL8LTy9bHXZiXLY
tIyNia6zqW87Q9kitHnBF1sNBF5p1iwVTUrRARZIHniEsvTQLhj8rLW0PNTkkYOgLzqprp6YjJVF
5GwaLf/i0APHAgMTmc6x3S8Q+lcNvo0+46emnm7JtXkzEznQYO7anPD/6TG4HRhdYD9fFO5rrKDH
ydv+aiZs22fyzA1Waa5FbSpGGftQsGhjMi35v4c5J6zNmGWvluf/vdJZ427rye4fWN4Py5WoRSD+
d/j4JVGCM1rrVGbgQ7GNoWX4lurd9RMAb5P1v7YZbOJflT+z7QsdYgIQPOdxdE0MyB0nr/P4iULD
TrfybwElpuAmC7FD+1/jrWjSxr2GOcJkABu/tC6S6a03yI7qQVxmQ2z9xk/Af3SJmaqKzm1s1Kg3
Dr/w3KC4J9lJZWa3uPXgKuAuJDtakrgVVWOzV2m59zUoIip5sDl4fengdlbTYYPSdjm/q2r9reBZ
7zAuwaoy1+5378FusVTwo+LhC6CmW7GPI9YGC5IRdiWnFDuGGi7O2a20bnvSXf3grQbj9jZzdLo9
HcPN8iWf1fW715qNEBRSJC9W7fFLwaX/doqmNH+dFMY/ZUMSASmHtbwCHd+SfsEgXd4UuSkfQPRu
wqozHrSawXX+6TCVFWPvFy5BW09pgeC+7gHrzYoELJbhtRQF11WWRax/dtPQGLK5tnNa90EPiZGV
rpR9kuPW21W+hT/ULKnK6kaGW8t2IfUWG8liTMrF4IWMZPJvKMhY4o/1sBbrRIH8zT6TW9n3G4bL
qBtmACxpycEPhgiM39cFzh/uNJ+X9wTiw/laa/+O3X3HcRhi9JLxngcSx0NSLbnZfFzf9sgUUktD
RMD9iT0YNu7zduo/YzvQNb2eE5uUwWQ1e7DP7yoLam10xEoPjIhMZLScS+KuQKeK7rIsTzToL4s8
RGxHuI0MKOHm9rLzLLAfW51R18bCMCfDx0DWBjVUshHpJZjyQmp9m3FYz8J361LRzF6MD6RqdHPy
PcBFr6NRJqo2HFCiA13KxVzCUSx6PFfSe2jq6dkavZRFbBFx1i7jFhG4cs09D7YPS0EYQ9w1t7vU
cbynq2ssD4f80ca31/dHfFYkTkOZDmuB1l0vhbCBL8ZQvD2vs+Yl4gSv0pawGsO6mLtPLqGaB7T4
g9azPcIXK6UZvvxRKOb+ZQz4f1D9D7l1US18x3gzoSlq2oThulzRnp3toRON7aK+MIYRJgkfCBV5
E9aEpOwNYNomQyVu7i/QqML9qwafv0O7g90WE1ly+KNi5nO0c/annVK1ssLcdibWUiKnEok9OtB7
jpRSNmmt6JM2MGJYcrRKxfIK5qeCOkJV4ftCfg/gBkTvaM/xwAMpQaQjDXPtKdhMl27bGfP2XHzX
RObD1LU3YrGf2v0Aje88Gk+fhiqhJClU/CqDm7YlL6QsGtjqz4CrHMuq5Zvl9J7SLHtJw1PIASbf
uQreOkKj3wAbUMdBznMH2hpEY8pXX88H+MdhYygu0mP9SLHzlR7W0zE43S5YaZ+FpCUcobymoZVV
tYP0aJwUcnk7fLNcN2kGjUD1YbhoKuUFc+Lv/KKYWpILuOi5WGhC92/GgVOw9ZFHyb6V+looP2qF
kALzBh4jCnfzRPrnjEKW4rb4dVEjBUFXrQ/bOq3YWKZ/mApGJwqVvhUmIxRVCUcW9psV5CIDCb10
CyaESnyWK43QN1IpmRuWIUrqnj/U0FZ3JRVV6Uyq0/zwUbX1w2JnrUp2t6epbvo8p2VMhpT/47j0
y3CbsSIgW9PpJbakXJZ7Uknsb4Fo8VIN1JoV9p4hVEhyPaMi45C3lE/I/1h1oPbm/XDAIjECxSW5
xbUkreAne0b1XWvFiE9NshNYJveiNJVQQN+JfTAmjen/obCVEhyXRoXLCS6wTDLl99fAKyDzxlHN
mG+U5saTk7f9hXsnXvwi4YIN968sjl1K+gBxI3yVn4odoPDf8DLwOO88jzZvK7tNwDmQ1am/I8p5
5T8l3RuXHKC+DGYp14g/ItSw2BbFEodwUp9Y4Kdam9MsvRVkdHPeWrv2OJt7rO/bM/u2Q3Qm8dCV
E10IPWgWkQZEr6XLp+Tj+Q5cKh8RWJGSZZc8TJGZLMjFxUlp/D6ss+5ZM2U7QZWR3x/xdgmTZ/l0
+b3GvwCKH9CsvYlN4901C6Aj9r2WZrRCDkRztwAYrdaC/xoDnLK6Dxsl7l5Fw4m+QgUKLdUPHwXK
RdIVnf5bYZX7MpnnvyqkH/eL2SEjnxNfBhenO+JNTSf022FpVoF3IjE4UksymGgqRlXY+KvOarpq
eVR5ur4PB6tNv5+9BLPyj7Wcc9Tv7CYKjnepGCz/f93TdKDUtU2O+eHxgeviiI6jaIZC0owUCGsH
S4X870AdlKIsj9zsZnJoqVEeRGkFsdapJeSqbt5zdBYFfAeZmwV+z0lOKISfhXeafZzWr8cwBroX
ceRva1/C8i33/C9/Xc/lM67/JOqhOrf0xmb2B6nWneYBWFth0BgQ3+LvolehBcFWebSY4mvz/MfC
VhnU3fCt+gVNCd/XC0ccVMJciXmt0FN8zUHRMaxRX1MquJXAfXEZtZG7pD9SVb4pu0b8iLS21JC8
y1mkRdNvcYyj5YFmQHcIYUVnJI1X+uorDPL6YkWp7w/QQxCQxoB3lF1OUuCFj1aaUZ/RJRpqKRFN
RTYC2atewlfUmpRzl9Z6XQzb1Il/nfQNr4lMb78O0kNoU37nqhc1SKrzDTEqObwv0FTAI9Q4NM2X
6ktMczX6AZaAn4kn3XNVWjsdqZ31jSKcKZKvpTyZrNNjRlKlcq/0WiD+SSY9P86/eSYVPiGbr5VE
axZroLrCQzEWKQHSD/Inyviu0n5+l5pfNGdeW5nA6XQLUtSjxGygNLENyOfgJ+suKfqSAEgc4QQP
06b47pPtstEvPr8zCyULbtkWB8U1FC4NRVSwlpJVLPSn4T4oqsWplg8be7EseN2JQmY8faEHMwng
bvtnGKFf2PjAa+aRIyrX9iX5rL+jD+BD6eGZ7SekyLAkSlanL8zXMc02A1Aq5z/v/sachudT57RI
DbRxcfy1bCX30ZSTbGjLcZ6rsLZS5pv7Mz+VzC08cnZJxhGe04EcJiuPfp6K8ja9fvJi73rudKm4
2ouoY5NE38oOjO5vOIOKWJWfn+P1+9JHbu9Tn23Kll3kPfNZwdCml6eeVvGc2+EnZTo+Vy0m9v23
Tqy4i6F7gzAoooHSPGx6kFtWctBvNnkBucq1N3Yvrnk0Vbl+pL3YFuuWL3RKXTaNIdUxkuq0tXBi
ZWRrc5IupQAwCkRS80fASyDICt88ovvZjT/zMeiZUDhlTXuNK4TjG/QFEqgwhPMw9OBrULBGmbPX
O8xQZbqkdOY5SleGECK+8mIUuzn7oyRYAKYeCI1CJZYCtjLHnXI6O+8ivU2DhTWgozsS9y+RALjJ
vf0HFD6vaur4/y9An+UjmFWxUGOHz2InkxKGn+lb7pYcXC3R5U5a99eHSJFrj7VS0ebUf+66O3ok
K42J5cSGWtpWaocow7DhNyI0j+1UATCQLngsyE9b22uGXSTtc35Aw795XERG5ZJjNClKC/oVnGzQ
Qzeqy9FSywxO8V92kpm9feLM7ubyJe5MXejkQe3dnZGWjGb0NG38dldhoGJPOzXkM7a/kOX3M0nK
OzddsNAJxeLYXrEVdq7bYqEst9nSE0UmLkUhyouyz4sSoqS32mxygdY5g15sK7HI01ojYMvmY9eb
1OpZ8+7V+jVDpMe0xfjXyRZI8SKE/P270xzmQ6OHLYT8kLp3XU9QzMT4+lcRuy6faobeg5NZBy/B
iT+VNt0lu2zVbEQr3EaYAnVhaazHHDSP60TI3jZhJhisEPN7cUAy0UumKIfGzTB87aIJRokFzJnz
e+W3do/ztPbH/aoSxNh6IRYJo4IFw+AxgzZ5p1Fe+OT/cXAVpRaLn0lNONe72CWAfIxishXzHYRp
T5rbVJL37mEMf/SJnFx1sFc0ZcafePfLZ14mMue/pDa9ptSbxyVJA/bccn3c918Ilep/iBBsMwIe
8k8Q2qHYhulBDFlbEoqgrGcU6cNJeBwCfvylXmYd9gkBgPI8KBXFNq23BnH5N1/acifbpIi9qZLY
J+jHoBDOvEAeeRDDQPzq0snURb6Sv303LJEoVHdldbLSTu8KQ8vDzmRNKP3+f9/sIkw4UlXLRyEy
cgXYmAniifj5sBBRMxUhg+ZNW3juV1kmZaDnaCt33ufmS6gpwqvdo4IhREIxejFLY1rcEFp/1vSW
5XY96y4mcEHI42djA2rN8LhN42dzhzTDZElNO0NisUz9cEmi5/Q/uVHc15lWPgCHfmGhE1T6U0Tc
auBMcj+rKkScojtIIeVV08jKyS+CApjvAbBlwl97/D7OSsXNnAk45VAF13zQ0onXzOg+Uhu7uuzB
b1oclFijsxk+Jgdo20Onx8wdVbdeSHDqc6O5s+86b/bRdrsPe2cboaRgkZqRj+u/XWM9ao3EdmKe
rqpuhWsXp/YUkNa2JTw2lQ7MQHli31VDct36pDlZGw1PEelJIOSo9q2IrwLQbW7wG40av25yLJUI
lpppNqukMxfhDqvrpNg500KW4li01BasDR0y3IP+Vxu2YTY8twc0th9e8V4C/M+khnajIZ/xfkeT
XlCo9HsknM+F+zi8qxfBr2j9GFBxBf07e5895+fWU21wxGLwV25jtjFyvE80t+qJyLDLdASuo9bu
GkrWglzPrEqpECimUWzOC7pRntUjFM78tIVKq/Fp8qnYkcJBQEL9NZFLqAVK9l5VqrssqK/Y5c6K
cnn7tSdbyixtPp4NxeNivz+mYSlBtx8V6NpUTDFadd/XFa9Mrn3M1my82hIzJZBWeW5gwmAbgKTW
rWcQJIyB8hq0cpnuR40gF6UNFA61V+E9aMhOUTf5w3CV/0W4rS1vtoM9YFuSoyBRxSXvZEdIPEWc
3r9HqLzTOAfeugSIUtLWi2Mj7vH5V0zcCVI757ECbJB2jNo7G7+zc6U/HnQhx6sZG3Zd2MFJk+Wq
qjN32DKgnoSDNJrsi15oHWzfh0JgimnZZEbXRXmiAF38DXVcKJD9wKIRfQbslmLjj233CLfL6IQe
+JLEQ42Fucl+B51+uLHfr6J/n4luMwmejwxGkAFJeII3LDGG1OcfAiqdqo224b5UTWq1MLp2yPi/
uQVYVx2m9+W8HqNjgFo5EOC42JWuRFPh4wtFdrQq818jknowJBc+2fb31fRVKCnw86FBFW2Fi0b6
ppsXvYL/1NXD9SJTf3ImCzFUTZs5txKVs1y9aSSaionhXXv6Pk2pPBge+bDTZxKXaQqELPj9ybhX
zPdZro4EZDOPUzgLSUiRCy2cymyZ7JapBAswBsS11iAQiCAQR90XRX+8gi1ZxG0ugI0g2JBTxuY0
fjCCTARwAQjFfRHriMrgqkhwqKjZjO5na0dW5N8PHv5mHebVHmhuneXJtNVt3ku8DzId8KNhElPa
gbojuhR/K4ctvZu8MdttEErMXRqFL7s+1mXBjB1CjPnA0b47/aYgzTLl7y+HWxde8CtjIZ7j+P4r
14kP36NthW0YKmFHXLettiwDta4j3aljheZNcP8lnLnKVnhMNECKPaQRd3+mGAQ98i+bs/RSpxw7
4OFiZ+Bw7OoNvzWwBMcux62fkzCPSF+RZmX3+U3ZnAWj4BZiiQBApNzo3xiyDejCUOONQiROTMLt
oJZ0aIyfm/IP1OqFGyHN32Uzi5yeZw/xqC4kguLmOEUOB0hPt86lPDrAEgCyaKBGsNWLCUjPSvY3
W4l2HlFQ9JQ5JOvMLpUeVn6+bEx7usL82b/I7TEtPUalv//hF4zddZRAz7t4JrktWtQ5BogaY9sI
gPC4d/7Yl/ea5WR4xEEmZzUQWwkqpnvGEcv2DBt2W+9UY56+JzH88zEvhGGEX7EjkY3+BchrEoDD
w1xKPA/HW0MonAkkpK9TilhqzfdellpQA+le4q10qGAv+hMYpVsC+R72KjJnJ0iKMnn1wFUUenIs
bmWe00xVDWX9XIK5FO/rvOshYeZp5hZs/zHm+TFedSgnrv5i0V+DxkvSlAqUGRDBjBgLJP5c4vBR
+FRutCZz7a4DJSi6xk8A0Wl5hv1RQnPw1zmHxi0yC8HYnDgtsPjMieo/sv0CFNV40kSxhm6iUaBM
58Y68yAq+l6eb2gQMHEXzN51d0DQ23xarjdHtb/oGWHLjFxGXzTDiuPTFOiwlXyNkpA4uELrar0q
4BaOz7BC8QS+jDBROWvWavFjO02whacqgsNjYY/2/XpRGHLufOR/vX99sqZfM1f1tstl9rg5Q0dH
AX6HCKpExCdPAXPqOmS6fPzsbkFb5l/TC3NjHz58W5vDEJ7o+4e5v8jdfEX54Ub7FEeOOOXKmpVD
EaIkLqnRknDJcXm61lcsxE1fvPzK+ItyIl82wM8Id/AB9XfUsgGELZ+zRZUwZ7oh9ieC8vJxUU5l
wQSVNUS73RX0W4+11gFnjGoUVOrQCgdfuLZpYr1x8SFhKFTe0+ZAQ54CZtnO+reATzXbPDSE96IO
4HDOhdde0hX2z5heSsvYjUOgs6mrq0awL6x+KilEVIZ7XqOwJF+Ws4gk0JuSufUPWEKLEJ0OznPJ
lldm92zBMicZxbzRZi1rbsEHGtm5AKN+i6o3ybmTH0VYzsrkYO5V5wrbAndtVyXr9Idie1/jU74b
szyg3Xm4GMDkftYxAv/Ue5bv3qaQgFq0mzHXGHDtG3xdxtumJsmVET92jD8C64FHzwUtpcUICP4g
5ZJ6emzWyt6vW8JydmzkqslTGlhGgChc2UVLad7iocf8sKrjt/NQZNuIzBz6b8tQpamXWUYi+Ew7
jElBQafKWvMx8cqiMGrYt88IfMCsgrISgriF5Gl8qeQqmjFVgi190U+YfPbiPb+LqE4+Y+5MoPSD
WBpDB2d+IsaSq6aYzWgTt9YfggrAmJQUdJh0Tf8KT/PwAXHnJHjTNRzMksTOY9QsQMo6SvXpMr0k
//iRtQmLmU7tZiyVuyuluMnHQnRqs+9lVWYKDUsz/OK25Gt4paD0LZG7fvTroa8vsQH6Bt4Vz30k
8HVVfjS6XiwT/smQgks2gajiqnP7QAJXmzhRvjtlX3Ca8gBX4q7N2fwmMHE6H0q3MNpUAoklGPHQ
djaiPkpz7Cf+OCPQiVmVD2rP4+UQ5lILw4uiwRsvJMZZYSqepit2w+cenRnJy1HO4OOcczIXGDll
bJ0VZxu9r6W6prg8LrTLW45BOuoL1mIwEs3avPHKFz5JI/ZXtC5jfebMs7Ca4hygTMvs2NwtazeV
18dh3jUbieUKXcJqRc6x7HBn1ln2VOgVbuJW9rA5vDoVf5VZo3qtCg2Oh7yyLcIyXCQcYSIdX/6V
A5BZLabqc+PbM9uro62oQ7McsIFpA5HptOs6V6gnhJmcW+xyWTihQpNd6rV+k3JdhugoaBeMKYU/
e3Ab2eIJKEt8zJ7yHu3ynrCxnvUEdSxovzzn16IL8telvhOo3hmckQl/nR0OUu9IvTQzpIrabJcJ
OFfe1bGHE/l12s+DdEse6GQLyAPAsGb9PsTsDlf6q0mA9gKK23i+cjez8zmboVgVTH0OZFGuVgC/
WeOfxORLkJHsT4iYndkmDrUIbZk/c4bS5rm8VOtfmFKTjRc7F15RyVBY0UWQ9LPnRi3u3JWH1N1f
L8sbaTA016ua3Pfr22Pdz0wD2/4jEVu1FUSvbHq/vKMXg5WKUcaEerXWxPIZiGhJPERXkLLLJFxm
XPPsRL9DI4KHfrbixfif42ZS8uSkShaiAYYuQb7H1+btYRGsLwRAwVzVan5SJVo212M495PqyQ6V
3AlD5VpNl6JGQyioimxeVZTSBDKWjnSS9f1tiEY9O5APxdPPMmK00qGV1jUivD4F927g0PqDv9wt
xbIJnN3XHl0Hhfof2IIKN3Df3TbZEGph/Qx5fVNgHfFQtoEQOkxUQDu8gUaG3sBPObfo4OR/c/Mi
StaJLmHntLoUWlUK492E89w6s0mpPEobMEuKyD9Yg/woX0TKRumP6yJJvJz9pYElZoV8oEbvfKpw
xzHnupLzYWDGjHCVitFU8HYabi+3c0VxqvXW4DPGzq5PsXlSDZH2Vg85H5ctdX6WY6VvqpUI6raS
aGOaRZtydN9JyAUTvFTMjxyRwHebWa0q0BKwHEWfp68C3lrJjn/rzBkB4LtsI9qXWZUwTuyYZReg
uomOjCRd8L28nKfW0psinV2SuSfwsxAeH8Fmt1Hp+zfvoLTH5SvbV6mc9b9LcVW9GNNQk5I0R3qn
1RDuWrh+HpfqmkvG4Q7hS4nIVdq79PAyBEXHgBb8N8gY+y7FhUN9ibR2ImbWoLWTNy83fdQF+rSl
p6juqLu2ONUWDQLkayRcpwqi7ySZBcd7i6pmGVDo1H1M+g/WmLst75CgT/O3lhs00hG+d3ASWk9y
yN5Snr9TVgkX6YGDiSY8Qisf6+eRaf8aR7exXaxZAqL619lNIFT2vWFFJHicRIpEEU/CwPw4Teq7
cx/p+H6hMXsEbAr2O1KLIBTkbo8m2dEQyOfqB2WTVCzE4zZUSCJl96tv728B3hUx2VFcgvmil5PX
UkFyzZ19E3oOqwG1ZDHD8zWZ8Cxvb1eFo1gMvFNiCx4w/Q1YTRXCw4OvEJO6e5HP8AGxL32uPksD
U0+ipu2/9qLA5oHi4X/mgRap4OfWjbAkFAi3kQ1lkehAJQTbgCei5mvXwaCuvEVxWRQX89lzrrTj
qOOVRgc9hfcwfRinoXtg9ojaw6H8HXn+CXMkCC1N8VPnqKwVRTP5wzBlR/GYt6RqCAiisFDlOfcb
wGOfQmunU7nkKlkXS+mHxNxoVWMHx72aq+34Lih03ES57eN0zChxH9Ql5JGQVP7t+Tu4RHUtJRbJ
TNbxZjkIEHGIHvkEr9briHcF25rdPo1AffN2DF4BtYY3DZML/gbb7POCJ6elgRv0fVDTZWW2QWmO
0Lf/JAQzrt+4jRKfqKFNQkluByHZa4zW/RAdQeNsB1L83dtuaxfYYZ/HD7/xuSfOYXNaVo9xIQBi
rbaR5/1oUpFw153ZPA7KHQXMtp6lWZaYaxxHhg/XRybKw7PiR1jMccbZZSle3MlCJA/T5RYwUrFQ
tRFJoPaBOCFlm23ot22sd7BlgK2kq3BVtDvQVLYN1tmh5KSKOimq+RcIUB0Fg6s9NntCkagd1ovk
zjm10CKXEKouO7Epmfdm3S8QFH7fJtWNnPl/rhhary2YLSBR0p036Q4n2+mnoXFJnZWl2xWi2Fi3
M8qYz/fota9PybUEIlLSFzScsXuCFq9a96tD43ZGXQdCmyXSyeqvLZflEIDa0ujSLUt92Y7afZfi
pFF5jLhaB/UCWqn/YBSShsuHFM0Si7LooQfCzD6BRPQmjOP6gioRny1e4L3NP6LQO8A8OYUJ9rV1
RPkdrGl4uHkuvBWnd7lMJnHEg4a/+HLimKZpYsV0tUbpMEsUJGDyCS3HmM8qvyGr/EBiakbkvPhV
wb8ArpH3sssT7lAoRVsilGm3KfhUg6Zrta9IJRuxTMMo8BPRLCc0KkFJxsFKIl/fvvHOcP0u1aEK
H1biKIW4xitVGTHXzSl7ypOFtg1B4nZDK4pfpEMPjP+PJVIUgyU7SJdKxPQusbG6gZ7NJLXv/xQS
JX3/Db98AowpV/TB6Wu5QeVPjIJmPA06+PEuKKEsE1id+JD/55bJblSrAX3tYrKEkMDERIDlGK0Q
S/1w3IfrzQQBooM0shmRc5Y2Y7CoWJe3EO7aWMCnCJ2lsmReVLgGOCFqnHiB1vbxGsc+/CfFYLeR
klyFuZ/MriYfukOxfZNSUY8Wz8VvMvO63xv7u6q72UijugyIg8WNuN6XmRUkUTvBLjnDYDuINOPw
2gt7FGaGLXCku6rlMzho+gY9DnWRMvnWtQCk9gTclmVIJZ4KsMBhttsFhUd3QKRSUQCfamEfTfr5
NV+0iWHETH7vKv8/xmJOV1nfIAce63v4VmYCDjJZnHvbabXlVR+bjTTyjuLEgcWWlHuvsHTV2vyP
JDOW/nFnh5JdQliOps2nk+t7f6k8ZYJdSESqm7DMBVzgvLaC9oTXWiBixOv4EY3cJHkumaQRwgbK
FYRSRW8tLqgv+gej8xXHDczXyDNdC9Gbw2KbQjiMzKahe5LAbxi2PNGz0siIB+33gp3HnPOmjCHL
fQ9uvWm2Qm6U+dFWXG6RhngwnqNLpQFdrgtRbLvEt2SysfEcNCCxsqOwTW9IJlGgUUHy/l1hwjqb
lyBfe+ExSqsYAEbxoau4PVS33Sd+5fl+zzoOxGyp8A/nnzDUnFrUGfbKGimX0QxJKezs6OwmSV1F
4vqikIfjjyAQYOwsoWxnaGjypAhHDray7dXE5eeT1QahR5flBj3WDhcVYLGvkwbVDSy81N3KdF8b
6KR5b2z5/TP6dxmZt9KDrqS8tvGho3ubXDwwB7QyOR0LesTwlclqTx/IzZyZ/3rZvAesEulBOlUW
3rhO3isIpKB2sv89jgyI/5AYS9COaM5yRo9fgg9Lp1R7TIy4MCXhtMBnwfJOSM0PI38FAB3lNuRa
E8FfAk1S52TTPJFyk5bGJBMOaKAYZnH+AmVFTek/GwL2NQyF6+c99BAfMaWZP1ARtjQk2eG3t6YM
SplJtPP3beM3szGhmRnEtzSO1SxUv2YH95Uj2MZHaBgfdNHFur3XcIxEi/BQRZmKn2mAfZ/4KXsj
cZ8E4g2rW96+MqeslHdT3gIOeWnugyMWDAG5SPhFnQnN2px22Ze44UwYwpNeiqm3EiYxqKSNOlMa
AGwFjh38nefXU2Ym5QvMobW/x3i5xP24eqfue4HL2Bh+I4e0ILm3ff5x7xM6Tg8AZNPjR71GWjaj
+AG+6bNOIN1CHwgsj4cXl9xEVD6DdyAj7Xw8t5pqzW2cM50JgQsiv0BB7SLTzMJjbkr3Ff1mfsev
4WF/+ot6/MBk+tMITo2ClJ8DFZc851SiJSq9aWYz6mSotNJTCQLCAcZ+haLijyDfdp+adtJa4WKE
S1fOF+03di0kG6LvFHEXSXx+4APLoVK9MyKuDP7y8L8jWFfz42YvSTtjm1HWIcaWer5OSKAGTwnY
iu34/pzutDPM/TqZqQMbbG8cgQSSIZ6ypvDvZouEpdgbZ6DAmp/alaIGYh4LgBV+butjQrgYoiJ6
OGK37ceywzQUQNDbpicUljHR6XSMKUZanab1KAWbNHkSYVRsT8pZzLaXo2unILObFZxksLhMpjsC
WXKpUybh/vzvhaVjk61S3DlWds2BZs9UE39LsF7CKNXKVYdRfMMgNuiQrz6Ed3QO1rhPzPjPEY/9
4ZwvvK6WKOmOKhQ4N3HMtwwbdoGWe+sAdVI12g6GzkeUQICGwgl4DpGQUIpcQ73Kpd+DXiWTFOn7
SJ8vh5xf38KU11qPeC8jGes21wEchzTDKWpOPbL1p16XhXN6GNHyV7NyB13mR3hlWY0s9smW6Brs
acw7GvSd3IoMpQqcWrq/gCn51rdPjNfAAn5AcWcWKKJa0ipGQp2Grzkp9w1+YAg/KfaCJFE/udUn
4rOWM09+URumkcQornarShRn8lZOHWsMsppSYk/jcOuQe2lf3Q6zJncWSa+8vPlFZDti7KOiDubX
JtW0aP6SwklSO3SIcLW2snLY+VcKe7d4qyJSQOjqGNo3rFESVTpcsKGH1DCvGF8yWuRsvN+kPnQJ
NOoGKVi0O1Z3y/aGQueyWtGMMcEgA+rMM25ysJ+eYP6LwD8Gz64XFYAARPI5J6puANa6i3JOb35U
vf3GvFUff9oGUjiqMuXLvbvPxGGLWgd783eBUO7BgfXyHjYe6nSqZ+M6AGXgCbR83z8ahgCxVbU3
sra/UbU1skldJVYPcC8+wYARGdev5v9tMVMONdQxA94mHKNFNK5hE/hR7FkOfYr9Stsz1344yYZb
DWTfvabFLxEa+bUDZFymjUh9ZWn32YHfdUAKTScMq2W+TJc0z0cvcb4UqCIJxKiXWVYpVyHmHOe7
Qw6DlNc313yhvSqzpDihat12e0uWjesCUxTK7dO+4yejlp239nbXHtU6fOJu/pJqpxWSDKTeSSXQ
yGwJ68C7xT+MY4RHvtU5yRe7wCoZhW/z83n8NVRYjAFBaR/flOEccLZp971maH43H+BniS3ljxqb
x/rIB03/ardhJhS1IizOS6IMfYrEDDR5fOFkVPJj2HR7TSixDIgYbeTVaGIZBJur7kItHF3EaF6H
41zcoWDP6ZO3udjmmamEBUHfksnz17e7sxTNhMMA4m0lACdsfZSrU/XYJQ7oweI+AnHAH73hYWgB
w3otGL6KU1K4Ko+AQKaPJLwZ1JVVMNq83S9vwkS0LzXSxA2gn2/wg9v2+aLtIz5w2PHJ/77HFuF7
9xjTNN9Z94bjOpBLOxDlAH0Ahl6IbZD47Qe/8MsyQXuI0PJUTSLOqO262KyqKWKb3eiJx9dja39U
QRtMQf38OrvFMxq7vPJydYD1VyrItr2K/Nu2OVPs1AzmKafPhV76Ylx73HJ4XvEd4u4no5pw735M
68b2t1ZYFKq136zALAahZJbdnUbhs1bAz+yV4uSQHoL0nlxpEXR1D1AqRqrI3DyuJFwGznJ4PIEV
fmUDYUPT9rRTf3zZfU3/l4eNIjdN7G32u0R9br/LZWp/bxxY/ULaf8DDV6/BlEFzd6Mh7ijCIhSP
Eh1COhTJv/oV+DCTIXmot6/ThfGB2MlrDnln8xgvKKvhQMT+ZjIWLJXDdst2Q+s/2489lIMGtHpr
kTLDYhxPeP3qgkiiN9arMezWZvQ4x2UvIGXtu/TbMxDjNEB+Gh8NOfhYOZcnGpxE1NU5vvhaTmQ2
fsZon6OAYsG0GNQxdfI31h/IGIBvztDkpk+nkD/OJV0EFNAYFw9Vu4zq5vMJo8SWEtXY68GBtIHk
YMCBPhMxZTElDkRowdx/jblaOjN7sC7DmZ9AKGuCszb7C0hPb9i1WfC/YA0agEbBg/3ip7eDjR7j
k4lILaCrWyuZVmkqdX6+sKP/D8WeELSevs3u4BvP7/xZ2Vr+1lbXtyyYwr3elQgskO5oGt4W2ZAY
bY/JFMyD0jjiwGaGCShfXKMjLL0oHDVvRCk30bo4DFkTVO+p8DGpIRUqjxauBHxnAYvUvVDYFjEG
a2fABV2EIeSvVMG/73KZIBSYjR5lQ7MmQ4DKdTIXuOdgO3vesucS8X28YmlmW9BGUJoIWlbdxnQe
4MZE6vKiSYu3Oh/gMa7jdwKqOWMIWNRRGRdIwiPcOWo5wEOpopfRcJwpsO5bX9O6nwPdsUJ0lda2
qoAZTIZziJ9vArcfdYcVxO6uiv/7k+cLXY0IFfGyc3OVjCV4csB4lS9EROnNX4sxG96dRceUiSwT
y6PoArb0t0UHdgejyijtfEg5fPovVO2anOiH5Cdmis/6Rf0t1OQ0YKPgPhpw4MKIl1yxDGCJ+9fh
W/5+dZ5dft2iDWm/OJYXgpH20uDGsTHGhDsm6sYfjPknpH/EANZQkRBzMrM+cd0mDrz5ofz7eY1B
3Mm+AsWvBjOpaq4dPQLjm6MO3amgjvXp3qxhYsy+gPfGddD5I6ETUvS3OtABiTe3bDAZy2di6WK6
dhK6ZT6Ve50vJwFKBbxpP2jp7lnl17ZwmjPDs2Qq/oD1DLX+jWsT41rGRc1bRtQOvbHNC+1ZtPoq
ZnR1Veakya8jaxMoL0p/tsnI6/Xd03nfAa7eOYevG8FHgle9UFCsEtHi7lYuqftFETZegaLbtpMn
KyL6kc1eMVWXNSGtUboVtkiNT8/mPPjZiYqEL5UNEYNCL0GCqOlPtfMUdbYU++f+pryMcsZUECLX
ADGOvOuaQqEZKXk8VaUPEXjo38lFzXAjBCgAZsam51UigLH2qVXUq7PqOfW8XpjnwSpQWbxGMvP2
VwN3QSDe+CLAKkS6zK3UeMQ6+QRwAW65utTseozS8qwss5fKHnjTjyIS9SZpiQKIZq3tEhy9BTVu
GgdRLWce14OsueT4Cfu/YpUT8V8SCtQG9k9KW+uph1XhejwygiiH4iUjH2nAs9ONHx+0H2lxjJRa
L9eHZjfTrQxWJYiecST0VRetSDTNXXSd0oV8/DuC4to9apeHp1YkeKHKRD6Om8AmWpSgZe4WnDPz
esfuDn+2SWaNMAXa9hKBx9+39SqDDWC5xfSfrj2MHOu4/QblOrEcEy9kykSqsw31CZINnAKOtgu8
+PGqmQoSZ4uZ/O87Cxjug9HJX1QFh4SaT3QmaiusC8wud44W7PddR5oQe+NfTfPGMkfm+w/e6ltn
N1cvN+Nz3G7iyH26iZ5Y0Ar7L8RaBUG49nZmbWJkVhfGfaYW8yixm50UupXe8gXt9RBu908KEaHq
z5Qfj1D4QTUZTTee4TpyYQJQp6HaWsbEuIZwYl6+YH4QYAEFYs1y+TMmsekLf7RrGdl2NA1DCJRd
qLK01bEeK7CPVwWEv/pGEVo5X7eWMj9VNPx2AmKlkeE4b2FgAIewJfB6kzBOfszqEJLfn+hCYFlD
cWqfsweenQYv9EgBG+yd1+dr8k04M3tCk9pFcgnCIrGbTS5EXM8Zyoqwi5AdkDZVLN6N7KfKsRVx
BRQBhii3V12Zn6LNejKvhMGXvSXlysN8XlcaxHjgV61xLFOEloPFXcLWM+m3k5oXrqRFk+CxkkVO
g+HZ0hvdcZ8kdwt1xiBV9TJ+HEEleiimorpsxDCM3UPg3EUhC6T/IlV4uKzVdwkmH/iKW8FDBJmk
AwSRsmBwNGKUbA3J8QTlRjFaBkz1JHlQ1CO+UmcwLAARWFxQl9W7Vhr1NvupHU1XYAd9g2piyEFE
Vhpj7OWH3W/ibKACw4mOKa0sXNXYhrmoTFKqA6Sliui5EvqpzpEZUpRbu7w+52BsXpJIB83d4a9g
qgQx7XcjoyHEFDuRSM48ATfKM+hLRofca3XNVt/lOcoCH3fEYNT05K4Qh27vsMx6fhMS6YiiRRyj
3AO7yxGPARGdmJIWbCfmnOYmp5cfqtjWFKV6ZBtbhu6VrI9vNdFqO91HyF4NGXRVLfJ0FcECi8hR
g78znXt3LI6dvOAbLmY7KSBPQK21Izc9Mo/SaDWre21wuA7jspyMDpFZjJwXixip+cS1vVoJtbMk
umpl/0wCP8/JKAmFBtQoZMUE9MO/6GEORMT8V9aaZHgkD4Kp4mla9dA8F8sVwuOd5Sx790YP7yLq
Y9C4ya+dGkwxNpsF74ztNhkHr4plMX/sxUitFU2+KJ1MBWcZP+qcgBJ1C7uVEKLQpoYZf1sOE5oC
cI7Xd7ue4IXz+NmwyR24a0Hzuh8ImRnC7jE4q1DxkyUwPh3JSRnWK02BPChcJBkekWqhudF/WmCi
RA4Aiagqgcf7l/leWpfoALJBv7B7P2FFlxKdG6j891NL99g0ADdEYOHZIUb+3TNl197t6oYg0VYP
0AYORRmlGwx8AV96JbCW2fiMO8u9fWECi0LfJFdTLnLy8kluk09tF3SJoY9oHpPfq/nc9usgCCdf
aopEnDyK/x8upwTIoKuI8lN54Il/0Y/RbztFIKxTFbngo9vuYImaDqG0mUH2HRoRSGoO03zyw+Hk
Jrko1rEd1Z64xNqGMJ3+7H9H2sIf9tIuoBkMBa1nD09gIz07kO3t96C74P0EwaHjWnuyanrhfLi8
cI9XDUvRCi0arq3Bld+y6luHJqmihlDTLJkhUDM93bWlrb8vcyiUdPWlQGA4HAuWzn1l3oROJ6JB
r4iq6c5OBE0g5w7FTBg5rz4vIIIknxrCwiopLKOpvXGpJSZoc40vlPCfY5ypQiNjiffr9aMECa4k
cjkU4EVXVdpjxahXq76IyLnog1zOYOfWCSjLcFvu0golfbwAE0r7yFaVRJH+d+8XPEZFwc8VCCue
4PmMmIyuZbxKx3qizIIMMIae4POH0yXJj8/ce6i5OCfHFPLNWnVHkwgyFH8l3sbnZ6rA1suTidG4
yfDJ8OCV1uL6P9dbxGcFIXnHTyZgZj/s2T3GDWl/YAMJxqdY2grUMtOVc8Tp63w7FMTBWRNy4R2e
SumgbLy677947zkxDFmq0fYv834fQl4tP9yDT5e+C/oxPzdKkklNdh8A2Zd8JAKqeIxuhEK1oj5Q
TGgUmGe5LLDMi2efmgiT45IlIxzIlzSqcJMbskWfvR9WzqOASC/n4qxFH4q4IWicxywVNETd0p1L
HxmwlsbNw+lqAuhXlWFymixOP+lwciGUEFyOsSWBiP5Hdv4FN4RPFIB+IeUR24QPhZksILQK5U1+
V995svmlonhX8p5oGpLEugC9EAghDBbKyq1pyloDWl4To9HAVt2GxZLZsEZo01fzLWvwg2pC1oGc
PmIErL8akbW3DP1WoSdiXD+Qh7SNXL8tj60xtc5xaGG7D4cXKo989ZGXGrdAEs+0RbKD//O799oo
zFQDmOGnnD8fXRjULva04G+JlvohmGhaeXm0WaI+YuKBFXSwjnX63W8rbWCuclLB5QH8RbvMQiZq
jaulEUpfsYvdPYrFfxSBLzb6WlOeQ9Cm+LhGm/dty/ZXOUTZpPzlLdqQlm4CZJT0wB243guWtAq+
uEPD4E6ii6q2jm54saKGzx2+JUlQEFJ3S9T1/IVTs7IsGo/zsd7ANcE5PNYo0/F0UFVp16CRMm/6
jeVYV4FK70nlB7aEghrLKGnv5ZK6MHWSKQNQAeqmCELWVa1v9v8CCYpFkddIUikLsw1aOatBYnw0
seDjjI4RM7PfLKl+o33tILditb9Zc6snYbREj43pCOBP+QdOAA220LvmTufyGKZLXtoyB+SV0cLE
rpkLwnCcqNwVK6PVDfw1f3l+W1nMfw1aO2b1cnJZBH5s/eD6c8kj3NpfX4SIlx6wesHSp6UhT/E9
4TiLe9mrmyHz7eiiGgnnkQ3gGVLDFediR4btvx+nHdnRSKm5uXbqEYazSvw0GNcHKBrxedhZ28iM
qsn4L7dqHi5Y1i91fDAS5cNdA78Zag+B7oMz2PRDnrZoyMGOuv1jCz8T1n4nYgx0fEU3l8UKzbL9
DmbqiB0Xk/W2t8qK5s1xgIvQR22ZeQpRZ1DaivWv6ecfEo6d7WaPitGjK5aqkXF0PWO8e4vi4zKP
lh+USBpv9AAolJ7G8bavU4OrtGeAau9spZOsXG/P1vnpXekHGZ+A3v1ClKO5Y4Ryn4BSIfPMsbnQ
ZMYnzTZkjT1/qqmPBZYyOMVowkk0zd5GyEfrpjWLTlO9Fw4l2SXktuCpVUJ8U3olfCoFDzgRZ7RU
9aOzWHv7zOL/qTUNnC7aOaRm184/fnp8k3A49KGJBpRreQn1vZdTIF/Ygo80G76Z3CmrXQ6+oqoq
eV5E1mUozbFijPDE90pfIVSFRiun22Tyo7I24ICf0JGeorSMnYse2KxMbYyQAwXUclSyNi5bf3CU
zT3fs63f8+CRl/F7L4hJUgJBaaeAvwvzBLuLwaAXNTQ0Is2T5XW54XkWmECuGt4yrQdU0ThAOWuo
6om8iwDJKpyXiY3xtRuCBYub2Tq6Iu3STRO8Z5uz1ZMNemexGMllihhmOjGrHMyMM7Qs2t8KLKbn
OppJu72k8ytI6xEYIFep44nogPVFRN8Q9o2WxEfT4hf3PnTMmSdUYVVFlvrHJzPIfZ34uTCHIarz
HUDNGVE1g13zrvz8gsCCGau1WdZCwhWtpF9qmyxzRiFk4TcB7WD5Jr4/jYSJxL4j12vkGxD3BAgl
MxZmfGY3Awh1H3lfXwCaRRIazgmlpmWBGZ9y8h42XREHytjSSjTqb7wGlB2TZf1h7utOl3hiQnwg
BtTfGkynpKw+6IOtR87jUgABtx1hPZBl9U+N23BvBguo4sDAS27OJAMY7d29VRBVlHgzeOM99vNW
95INFy3ZZkOvUkACef2K2SdrdzqQwzkmPaMyANNFiqDMtH0FMVTWUYntfqNGJLSYJ9i8C7kz+gD3
TqaNZ+T5OS3VSzeiMuq+dT1URtNhDmYurGyiYPlL+JOm/+7VFjRgx7AE2lIKspGhY4L+SXntAKcc
MdgurUW2+3Q4sr6UoffdGSfQr5LWwhwV826C1+1UPGfSerA8mZEWdwnh8Dv7mekCJhCFym0aknIW
0k+eSzROHhOCKICQ1FzmYgladKr6V5WB1lPvLR2z9euySywgC5lDGyi1bj9LeX4muvAc7RK2E7cS
63rvRWFVn9DvKJRwnI60BU+4TQAvmScmS7iEewb5P6baHYaGGh8WC6Za9PCOlIWNAMZJPcYO1KbN
G5b9C6Ke2jsAry+bRMSYrWmwlMyvK2bM+2NT8otXqgmaI3u0FrTjKXX6JLXP3XdIGcXsAAM/GMdT
t06uuWBf0cv4Lzu8pZcDxzH+4UkGQ1+EgTypC86ekwVqz0XSNgDGZbte47Hm7YoRo75DsuBC2/hD
4APcFkG8gEIt+3wuMyTBbvWHS0FeCzcgXIbNRfvLh8yQiduNMyluy5V3Lts1yWOYMEsiSDQuoLgo
8g49V4TPBLuKduAK6d60P0GtXPL2zlPRhTawlpH+XR/95LEHRpYGaJ7ezWVbJmac+00mJ5OR4egI
9cTATMGEmRRUIdQkPHt/hE8YQrz1lZ2lzvNcdmX0/WiPNhuVLzEvJKtPnDqIeJdCGlDdi5V/ghur
hbww0/IAdl5EG5RSqTKl3jdSz4EHN4zaKT0R8NI8OaAeWtO9K1XjTBA5P8GLGjoKUAr/GI4qd202
DbL/DtrPycejDdcdLuh+b4WugR8cgpIkz5EXgPID87OTHhKlpXYKPos7igw+qDufz3SIQaX/1iYk
UY+iePdxX99zHz/Ea1ehmFZN1In255KxD3fWsbZkQ/4Opdx8bmNzg44tpWckga6JPua+KA+C5QnE
tgDgmjj0CF+iBTgH9dZAQkQqRGvRhpTmpqe8Qdeoatc29Zrm+HI2WmfqJt6j4b2e/vnyFUs1yME/
h3gIXvRsEaCf5nTlv31/RZeQfDOWSWkpkPolkshCoW99KCwfk5YbJVMBQpWJDISQxcCs38x9dF9w
wiJ5J0ZcF+gBLYF/Z9J9MdN79JVBhwA+pwg9hWnQPzPhVAhfjhKhGgbXWL/XZsvEyzk8nysVa2Yk
E5+aXKetMLi/MUdALK7a4oJgtW3abC/HyiKBBieg39dMuHA4xcUOJjQ+NPGSqVyre6YDc1r2bUsQ
XoATAI7Z+zkvSdP9j+SqjHWhffapLapnbxOkz3dxF26Z7ILEiLFkRD8gt/ZMEJdg7rpc3TbYNbPN
pH4STJQVgWvlV3xeBESiCSbI0pJB6LLXwdztFeRMI2aO46kPNiy89gcflbkEDdpb1ztsZIm9x1Qs
6VH5B3BkxJNzVOZQXG2ilLtT708EFKr3458Qgmg6clFEOWeQyLh4bHrt64Wc2GU6go8aT5+6d59I
NvLt+kehh/mEP5T1VTEZQiuDaowvd6cx2EVhKlw/rc1j7igd+OBnshECK7m0OkUU3otTiswZl5Gz
rJTTknf1wTu96l/BSHBIyvNh2KMVf1N1nXyUb3ICjDydx+E8iRk5vD7KOxsYS2kFvUVGfak1Fd/N
xvkVJIof6uvSeQb4kLg1uOLs/+OTviJrjmzDLCRLYwexXEjHCMSKWjrLvJcvxuxDJyJ2PlgnBm6z
I9z6kdBi4NPEpJD8kIt4NVxbKdJKbhyyqTd5skH/ZnUln93WXOEMG0UsJOfeHF4eOamBPEeEDrQb
TMzQg8yAK18prcv14zk5hGzy7jusLevAJXhkaaN0WhdYDI40gfzz6Xj70MFFR6VZvVKDQEP7Y8A7
MClkiQRQkfqTkmH0gOcbEkWsEx8f5DxrdfyDbGGFu4wG6FLQtO76KSk5vTAQD9g/4COzjbk5RzyS
fwe3Yq1sq9obTqmTBuZcdxisjju8Z7R5tdzhIJNzdUPO2RL59LCwo6k+4xX6SMK5vF9mrbyWXIj3
KzEtTc46DFWigFINr0zSuJmW+dYXdm9a0+lly5fZxAoi1e8kBDLFU+TKZmfI4XAbPkscNpSsIz3r
iToKaevKp9ebinJX5D0/r5ETPncYlB6SreTKmu0D0maHfPYxpDyFMyvdZTPuCB6eBcVf+pir1xxE
W4MNiRIe7Zetp8t1/JGAG+1O55tmdFpSYQGlNQ7U2QUxS6PRdgPQfPs9lIqi2JW72lMtdenM2gWp
OHtfzhyfQc+mAdoCp6n2qLlAFGaTFjyqawjSObMuT3U9MNpqiDXy/PJM6WYvmfMSIiiondgU9AYE
dnfc6Qkg/wZ2rvFqymF5coesQ5pwTc8gJHGdUjU9GzVFKDsq56frIXtDJgbJRHvKadC+K5/HzgGS
aGj9b/eEZxJpHbQIG9/qHHmqMM4hLz9NirPYGYmKL3ZIoXXEk6ebcXljtg7+QhRBLWtclpA5TiMj
mWuZiQm01h+WhBZH+4ox3i9y8QMbepsNfUBiIUMoeKWCB70ZgeM39OqxwYS2+p84+sC6xBP+aLWp
VFK9WFMwDsFnzrsipDoFxqeq2KtZcWmnt3oH1+d21oBVm+SxRqS6KwGtbbTnLZB2hkrAGvZsmdCM
1t0XHxDukUWuvlYIf+us2GOVfU1quDEFtms4GvtyuN9WqSbcjHkboDBbazlpzu89KECnIExsAzU6
W5mVYMyTSDj2DrPXNkUOhyUYGkHQMVbGEP/xwiNY4N7NCNy4P1toTGwgsfFXJYt4dYNritCArctV
fajy35s7I8YyRA8OD29kR5aHtpmh2FCM611MgFw8S7OMEXBIXLgcA9FGCksRUakoTI5PTlKrV2gP
Ree57I1Pf5vEomXOz3CvJCyC4oMj3p/qNh9GEjw9cpFRqhxw4A6VYhXk/SvbSDPNIURbg0szOX8Z
qTKGK4nCfMxMcgPGJ/KijcpyaoVLsW77VmJ/ojPAoe0TED6cnelmey29MvNTZ71DDo8UagWTF3F1
Jr6EJRUmRG87hHoU6WqDBu5Hi/td0IepkTxoo8iaGR8OOYHS4EhgUS4owLFD8ge+ruDiLLl8BzaR
PrwKBIuXX0kbcJUJB40Qcjak+Y0vd4Eam+LbAHYQXb3o3yBoIQUawHgDGOTpiTh4oqY7t5SnRHr+
Qwu1JC7d+V0BqoQfDz9cAMHG1lWDxBPh2S9I30YHJUq3l6+1duqcTdtk/DWFlmsVvEoPLu9L4pAq
5Okg/Y6xZ9/WpBDRutFV5cctkNSI2Dt/z/+dRPacQKz3SIHj22tSn+7d4TZ1cBMlrVaI6C13fJsX
on2JBmngqM/QAe9iMhCGew30RIf09+3O6m53fQGob24yulh/iw8Dq51Nk6GEt1oK+GgpYGox53qu
m9v9Cc1fvuVVJt9Vch0Mh/sjRebp83KJjJwfyPcwzHxv1zLxBySAMlxk3r+Dr/4E1pzlqZs08u/p
JSGEmnYDkQqIv+Syal7iMsuDIzPpMh005hiprXZznFnSXItCCyFgQtfB17OMb27UUVWoCdfKJP6Y
LaZ/leDngGtPEgmvpP/9A8omQecvOFtCB5pbWXuQeEB3cuoHgajPzpyMuOUO5RKxe5z+PK6Hb3HT
WGFfprr3DBWD0M5lz3iM6G8PgvLRvID/8oc5w1lkZX9lNcGVyKrYlSVy+GDKv6HEGBGhhDIa9go0
+eiVjQ4y+oJ+e1CX8B3D8YNIIjpKhZVEhE8Xj2oVxPEnJn4Uq9nAqvmEwf1bnbyMobNUQl8zdMpN
RYuUVlmLAArQ3GvQTCJlV0YuiczP0Pg1uJ9AbVpz4C/vkIcjMrIY5PRlJdvU1POSLvDXIKj366fo
D9Bgz/9Ubn6oA7Ynvho/Vy5g+dTAVCf90NNEIvi1zd0K3P6tqueOEaTko46odbyxHZZ/S9tNYHSb
jRpfDyDHOvuUQG821yGmNJRSOxeENabGLazK702VwQEoJcwVjRZWA5UeyZXf//plmZ4yxFaey85m
y0J68+Fu8m9qLo2TG6xrowtFmZ1L3g6ARiwj4h/+ukEa976vggztx8X5vp9S8BPO/TFsoVmZ3CsZ
6W8wlM1in+Hrhmk50L4GCgSrBGUL+FvazgxaIGrQV5GA2edexoL9s32KTRhkv4V/KZxzzfmuCOr4
6RYvUfvNqycdnPc0XBdUMq+IbuMw32EQtvCMwnJHVUuUNIQirzaTvfpI7/yhY6AgVZLascvizTdq
MdqDhaXRxxfzgQi9yvLXNkQ7WA1P6x6lNpx0PQdlzduvC/0UIoZMj8kDLeNIxVTZ3ovKpJTRUP/d
3PJOn3E7RuSEW6emf5ApCvyL5yHGotgZOTgMmcsd8sNql3z/CmUn0PHuqOx7OYTpR4sXWpet+eJc
MD+8L7RXl/yPRtGUslSa8mSYTT6qDC7jtAIKxWuTwjVqJE/WnMmrn8n1ucRoDto0X1HGsxklM54P
DfYjvTdhLNsqVGu6P4w0oR2+ygIyhFCbZ9XrOc67nMAUmlT9Pyyyo5DbHf037tTZOrNq+E7lnBaN
F7a8dLpj/UYYdf3ZXn175qRa20InK3Uo9ZzUhoORKUyb6cjr88mE3pvm3bHZd6y69g9B6W52kjwc
2CcL4j1tgKsihJUrEGKzN8wM0qST2O7/TQirzttLd5tyRjOK7Lu/fKgxYKpZBXTcKE9EqXfVPpGb
hfe9ZuavOPU6HiSC8Q4O1xnHB5G4hz88rJSbKa9RolNyaO9AuUNYJMArvgRAWHZVnju7IlaTG2MZ
1LrMBO6yuHY+fWAmPPYXhXAt8FsI0/EiAS87MCbd7GC53v+AlPkk6YkNvZ8Fp+cEimjgivNVtG1C
tUkGXWpGWZX5Pi8z3V56eWIOEvCpK61RnQoOAy4Q4bMa517duBeR08jzlmsGzPljjfQVJ+495nOh
UoY1iAdkuq3i/1PdUtxDFi3hktqNgAv5UY0LvZeG80tMe5ZIIKwvNePG/qUqO0Wq0IglTSxbZDwU
IYBwFok0Bm57Zn76U2nnMzhuLdPf416jTbksLdsAebQPnGqDnzJsbgAMUWKU/rWzWOg5xoVFcSxy
iANcydF+rMKJF5zXxiOPoGG+fycXSpAafNc6+pMLTStp/i7oOgwBG1hfqVsaZMmMMIqRzeFXftNz
IUsJUR/zZHUsmfXP/H6fJd74VCIKVTLxIxWxWkX6x8uA/kkeVJdcMAFSncfToMle5y6+sCRQQeyT
6Ys2YGcCuyY6Sazg745myjvVXXVxPm0kV9eUNvYv947A1lgNbQiLX6y7ob6EGzxBaLkgZQIVV7XO
XVKi2PZmev3bATBPI9uY7Qh4olx8lY6JAiAU8W6+Mgi4e43Xzyhd+NZxQchWF4Z9IhBkTqAAsxEm
cH1M2e0IeB8XCaKoZdJbuLQ+HHQXQRFYFziIYqjQODP9NAjsZsnqhCeuchPIgEshybBg+jCkPhcw
TvxQmXpT7l5PZrpGrLHExAlacO+FRxGIayCAwqFU3P6R1j+nSvSGHvVDHGL4QRebSo0ZPo3HdZHi
V0aU7te7anfpNiHZZJ9cfZcyAoRa86xlXBvTviI3mVtt3QmfXO3X1QGxGeJ2m9itv1Y4a3pEFVX5
xEitwuSYHkomJ+wuRDCbcZPD9D+np1PmzpblbkG/+ymjVPy1zAiw4uBSlKDJVXucxdhHaZDQio8Y
g5FWTuE1uLkxCjkuSta7d/+pdsnfq7TC4KeZa0yLSYHvpg/rbZxoqgvzTLCgX4KMBO/mnjZXc6V3
lhVT0vm80DptpELukyLO2gcF8hUmeriegL3xWJZWt1rEamrwkZNRVFEAKuGxFOdqdJ7NE7tAW/qf
SQaSyww5xBFK9EceTqVvDxHS5aOEVxy6R5xBwdew4PBAIxS19nc4xSHi4gUp5WX11JQarT2rP4lh
pOLGoibeLCEKXsX+3eFi9Rs1STCVGD3B98u3JEywL4CeOPMVep9/OE7pVA6szOlYdn2cZOlaWIk8
P4oC5gqhbyhVnbjYgDBRaB1LkxskeQhop+xHq88T7/ZKpr0F7zFgBq5TFuMf01qEwK/sdOGBXhSL
NYNCRmhVycKO44J1y4cLtEnA7bBQ3q0UrTdhb9d3nhAC065u5eBdWOxS4xaAHxaBrWl+JnQruuG3
Ofu/96SGwFBl0Z7tIV/Ko+b3wVeTV9wiCiBPMOxTuNnSvaulLf0JIsSH++0Vp2j8fjK+IRePfuCY
9NFHc48K55CghaLsYPM2IrLAU1gre1YScnFhPbHdkKgVuxlqDmQy6CAgHiZfvM8ANvSOPictdA6r
83EGv7XpOHfpswiT+NhIQy5KOWEt2p6BeRfuj0H+yxJK8eOnqQD3EPZWJs9dRV449daHC3I7IzUO
PUG/VzGUVL3KGs3AuvHckER0Srl3TVZxGMF9ofqD+ezNvkqi9tD9iah5xYjTay9UEAAlb8Swttp0
sgLS2ApYBP2oSpwllp1kD3bx70QXQgaTIoUofkQQOXfgjxcED2kqDnm3go1oC3S+0d/s2Mwiiybg
z1RWhb4ny3061rWMVBK1mmCz1+X2YBEsxH6CQ3ANIjp3vO3QgBUUf5SswAHA7HD6ZRJ7EtVg53kR
5YhkhbfxQvPhkfhHHzFwNTIFvjNladSH4cf1mf0nA7gLxZ7aONXIYq47qXjsRIFySi5sDtmMn3x6
Hl6py1ItoJ49+jg+3fNASZnpWnu2r5hlBP0B4LagJRgoX6Z6Ed+7VGutVypqF9G8NaSO4FT7oRaM
jeaZkuZQ4uHROB3SQPZaWlMR+z5xgYR97RLafY8W72I5nqu10v8JqWuotmsJ1TlMwhl/ufErRHA6
e4Dysr7QwYW5R+W2HDFyfdFtg60MorxXCDgRSR9Le5xyMJM4xya2aMkzykfUM1JAMWpn+b547o9J
8c6ZJJBWTOOOqzCDc+/WJr5m1BDo/+f0VX7/QeKla9JZxQtci3ExoZrrd4ta4VNzG7T3QbNNUJ2d
tMKhB8SGReJs4CfJ5+hlqvYIDblnwyC6EFy6XRXqAQ6r79y2rgD4EbcwlK+im40D+TOjk9vjjrps
hAnNHPsEr3ATT/RSYmbN9sKGNk//kiN1uA8f1jU+ToTq4XuIzAjUBRNHnJiRX/EyJCmMiive1x2G
i0dmQGjy4HYLm388RVonsKfJaYQEIeKVscHUqpmWpbjOe2A+euAh59nT+3ipz9ikoHxF4OffrJDD
FPtlOtVK9HKnUhMLm/f33AKwdxzKhMMRgrv1fmpYSpHl+XIsNyjfd9RRVzlI1Itv7G9DOkL8EzWH
es2cLwayrpdSP12xxJ9thtICP/oirLLQnNQ/bI2UOycOlP4lEWOhCs36iwr23i9oJ6/uCvX74g4l
j5jxiUpXrr4v1BAC85tpNayMCuJT78/a8+fm88lN/PxbTXNa26lKac8jxm3ZA6h52jZGiSdnQXAQ
gatQ8Prt3yFpSTQIfw83GypI7/gnj/zEIAHq1MyytR3mNFum4t5PDc2VQ25P5AAVxcSN2EOcjzqO
n9OHGaYBpd5DTMqnYbB70PgGd/5Lyj2ubH0WgAdJagwQfBNX9fQNWJ8feQcEZIETCtgVUfraxAt+
OawuyLGXyEXW8dZdbuClAlkM3/Nevf+wO/5/2uXy/3jZPJc8yN10/pFapSqUYAcziJumKuDwn1MB
+4HQHbrfR1IByhaKJK0QF3OaUUENgtuAJr4pFCAcIHVL4N+fI0Au3cl2ajVN7TD7oKA4G0qIv4zA
mGZAC4f2jp0j+O9iWFuMEouIAgpmf27CxPG0+osnaGdprOVyMpEFKCwCZTtN8d15tQ1jgIyyXfKg
nvN9noA/eEux423Pcd66IpogflMmLf6m3CEoc2I2uprEX0pZPbByPbOXrMY0/Yhz6HfPgL0qgUlV
S5hUa5QKTQBEFUezHTpW46/KbJhGiHRIkrvvp6ZTabO+VA0yBPTLOF0sL6aTAa/Rmm1vGsp1Q5sX
JhZrtfhEcLrYuYHbWExuFU1r9hzcKt5E4CzkgRQbyY3Cos5HoILuYkeV7j9XJHu8LvBtTBzimPm9
bCr5lmXnEx/yjC9YAXvhl7mvorY6Y/dH32GGDQXSfXxQO3ONkbFF09FIUn+YYvmTrTBN8ogyxFAV
s488xCR3FPkvaNOI7bBpaNywoUtbPBLx52NRiKiELW5rH1vPrEIjSR8MRfmUv1QZX1sMdrC8L75a
QiPoUlg+tnNKBp6ZbwaegPYzB3mMvoNSMNigAq1n4u48gHkJXMk3hwuzvRoLZAilztAMoKUkx8Y0
O0AXGijNWVA+61WXA2I5PXt8vKNz7i8/JMhQDa4b6vk889QCpqgrSVFmoQ9iJhK0eH/hnkE3rTwX
+QDSDEuWOEnARr8EA/GSBdJKDs7VmtscVWECtpPIyZqlgpoHmpYiwDAHxWPIJhZtfOWCS21Mn0AI
jamSPkWAQqrjZuexm5iClfG6ZlEBxFxyQNRf7b2D31hkUi7Qnd7BaP2Cy+y9Ik0EW7DZuCTnkD4K
HnokoXSWb4J90wc/H11sXvXqqCavUt7P3q4i91HBsDBPJH6xSSwUUvdHe6hVa2Sjp1B8pK2jb5Cn
pAydGkeBfLVX4avJfvqXXVJFdPAxGlr/PU4yfE51TVMKToXECcFMKFCJxLiP4RK3nB5EOUqPSiR7
5naXF4pHLfz1dX9sFR/FeXcyGoO0tMnkUTrzOoTEY6cT86hEDDNv8lsjtMr/i+ZSXp2f/3PQI3EK
WRWmM/ebc9i9rlNL6MDcNjBw30piYAUfpHVi1Q5szP7+AI/U/YO7ZnxNqhjEZTEUKe4Pzotcts5S
iIfDShSPEBMEkc6GPWJB+VhlyZg5ruWM819LgWVwHumTVwLrS41ZnU6DCQIVbtqpgJMTqh/RN0zT
MO19H644qD3nJN9W/iaJfG4ta7vXlGvOFTZ6jRGaxJ0ocQx/XbnjhTmss3PuF2xZUvKCyJSgr7sG
62rnDUi8ZADOYszdirAC2KXik2yGQTf/lI5n3KlzomVm82P81QHbkaguppMdOYJTnrQcaknk+8YG
7KxcpxHQcqHGEeZFgWin1GhLdUvrWdh+jnbtSagaWWtARM5ytBC0pekXxav9g7+bFaHTJgAXYl1W
+V6cTl+Iwxf5pPjlTIPToonHBuKouzAX6lDbeGauBk9wY/Cg/Vvh3//fFw4/5/mF7AKHsAexj0g7
Tz/9qcp1pmteeNQI+3KbJcqNfT+FGsfkxQPLPHe8iO0Ju/CcSmvX+ubaC+7M0abH4GVNl0u52+4W
UpzXJAF2Hl1gvkO6Ai1oy7++vm4n8/NrQBsaDhMlAfU66+Tr4+9rSuB+Z37uqcPX+9XqvhmG5+8b
PZG1uvsoaAUhAB97VyyAQnHzE6AqIy29bazRhMzly5UmsjJDbCLmy5yl0AuyVlB5ozAg1/89BLNV
yQnadjB6AtCY9cVHl6BrwdqQTWbTHNMxYjx9Z5s6dIx+qb9sZQ+7NW43t6zjjy0/ECdMYaDvo9Ff
ow1HFOOi1L8AzZTJjkS5dSoiPbjpCA5V6r+G+wT8BVHeOJmeI5GQeHoW7PamCbWfx4g9lacQtM/f
IGEoY4SkY3txV60Cb5kF60slTRODCTdsNlcBl6Fgl0xK4RoBvDBx1/OpMQJrOogQxUx+lQ3WD/a+
FE3781e8Wq+h7F0XK3ipNhVMV1i5s6gM1vJyIPo83j9SsXhI0Tu8YNZ7y8YW6Dz4eW2C/er5m4LW
zz0GMNkNSsACsdigToYtTWdqq8yo3ryCwb4wo+v7+eT7tS1ppd9k1qXBUQs4V8FnEgARu/BM5VVo
iTrVydB2t/NCk9A9+oIn5L8MmQVuBx0aiQlAeIzJz5SbIH6rYq5uosZ+G0VWI1foxelfvMAIH/wH
6744VFK2IQkLF+fu5CkRjyqhlMsu/WujH8t15GqLBTymQXu8UHA5VZjXH16E6DWocAB7l+m/Z0ws
/M7FuKXaDxVKw4oslq3EOJvcRQg3a/OqKFFETIyx9K8V59GVuNGV28JOnefZ5wgerKvC5oM7qaRt
/pWnTShN55+JylhqUbFAeeqQ4ZXc594F1vpM/frpanooP6ovZj+Jei4Mc7gXTICfM9TMIKfQBVqy
eq8g7cijXrajvgryUKOltNJDymJjhkZHLn67qwoo1e6P0XyWiOwCyN8C59C05wZ1+xu6q7GJPTr4
Aatd/RbDyFLwWAyuxSsZLtRezVcEYUp/ToEfDIVHGNBrnfIuFzg0hz2FFzXyw7pJ59pftZLaeTcQ
Dzvowg2F1GDe1pzmt00KfajTF6r+IwJFF5z8XlPcX18lwyNwSml75RmTIAIHxGxklwwWvynZ68gu
R0IBrMzz9dtV+t96QlVBkG6Y7h/kB+HYYfAhcZBF4cvB65mBDZekP3lNUsq2Qm87DL4ioJ+CiGZh
2GoA+99mSDwVRp91lIRYDTcnbaNNyoEjnFhMHnuM1Ax9zSBYzgD+Q2pItvzI65LdjR7/eYtY5eMy
fkmtIxljfXF/4Tiak8UTkk7GS3lFpvBidhk8jV0VbJG9RTi1HwouSq68AWLgqZxIQei55UeHDWAO
VhbgZkGt2Z5Z0zT7Rp3Eh/mv6C+Fl+qqQiamIIkpx4qZ2axkuuDsAqnj+FL1Y8p7oS/0c1t8q+ZE
BlvFrju0nwt3isWyta5AGDaZP4EcMBBYFeWT1fQy1haOLfvuBPkxJvsj2XK0dFRzVXmrNWgifssg
U+yhzLOjJxFhcT1onfkMXyTyZt+ARlrai/07IIbDiuq3wWobHiqwTcjtvNDkwOtWKDBxLPTDAa1u
j8vy33m7FFaypOmF/yOTJnvpshClapLplmZ6Yb9dfU3SzA+X8kM+TdG2fPVNCbPpL6L2jvzuF9Re
weHO/574CDU2iQHfJ6CE2UXdq0PC02C/uoz/O3keQK0eVQxGm92a1rNnoaJGmjXZr/zOCI6InFHT
k4OOHhfJn6CzEyEGv4uLkeznKYfcGmiIhKS3dazAC7whwTSDAD/7yqFXaMF2E/5TAAYbJIsjYOC5
bIwx4I7iArKtFCNBcxdsL4IlsDWwKS2IYtHpZctAQWAmX2lQsPdor/YsFTS4P+T+/8UpApXhBW45
V+cl/0KO0sfhphA7mA1RO7QgMNDjEIysf2zGCYKoQYMNw+qPsP/BsB0u6gMH1IsMRWDxwKk4vEiR
UFnE7KHB+Xj2PiayIbiYE89druikiDp/oRxC4+ee2DjndIZ8gmRVK15m8k//5cFmeR5QJgSuCCZ5
K70vm9x5EbvxgPrIOqQeLVuSYlqsfD2Ip1e4kEhpGEcZJzOOiGL/GCGVU/5xs6q+UH0KnggnvU8+
ej7wbWAMQOSo/IRMLXiQhTKfQJXYVQp+ZCkbYx79ORY4X/LUxSRiC5mE7BM6/CYW2tklUb/bjwq2
V7jHgA5KC+e3hzSG3Hw/mngN8ULxUoll9a3gh3YqpMfTJFEzvxI5ld8jNHsaf0dGuaQMAp9X2meV
vyRszhDFfrNzvuxuHmkbkTO7nqgFGUszGgiO7iv4wVU8dQ7Bx22GmqH5yl/bX8OTGZvd0Ueof7Ob
x+K1zqFUv+c130j8PIMFR13jU75LIgcjMfIKfnFBealmLfu2jSKxiAT/C8t1D9RZwvoOamDW2r/f
3YzkSkPBKx38noLyLEXTvWrgi3lCfMCuTGk2EWSRK4Asvt8Tk6QnT5wN4ZXZVrqKiyfpsAkl1+Uy
5+sUWSvNsJBCb2Ju3QVNXwj9tkJypLnor8c9TnPuBEmQ+WrWEO4Z0WbnYb3j6bdlMUKQ1Akw3uX6
VUExFkhgLgWsqTS7tOdFa8ZDNww2RGEmHfq/cjm6K/abJmMAuEl3/swwpRu+6thUUXpZY9oUWDFG
T6UTHDz+IyIEvKqbImq9Fp1jDUw71I11cgXwK6SFz4zqoipsmwD7YwzkBUGHsB5gvVymrCIpRnPv
gCiNA3Qxqdw7zkGC8XbrTbBXtf1ZkHwHOrnmTC2Au06flNtTYltLMRb2cWuRLwETkX85ztzaKA+4
Qh1wc8xd9Rn9U4qhMrABQrsvT19Ptw2h0Tq2vztgi/HSA9ZvRmltKwS53MWTA6Cp6GYuftr49pV4
k+3MJtnIQWNTj9wZnLHp+dIrgpwV9FQPYenhUqAnryKq4XCPPC2K9JOTX8nxn/kKgJBPUbS30Pu1
Atxci/0sP8OdsPor/T/iigW1txkpoBetGQDgDYo7o5YA6R7QHnlPc2lvxP39XftyTeO0X21ZiNJn
n1qYCXtXyKaUoA00ULImF9rUTbelX7BiKP1K3+iPRz4NWlFgrFTCXrK2W6twEad96Y4V/syhnh43
zWWe+ZzObmxECbEQehIpeDboGzaQBAEOtGwTHAc1SOwLkgW0whhxTjAaDJvagziEZiWaWTs/WNnH
L26F6xSWWqrvpPO65KxHD4UA1vl6pPKkTAZfJtoQ0VMB37o9extuhBIyEaSDx93HZlmWdpKHE9T9
pRbuNMUSEyR2INFShAyxlOoiwXuXJPfHvEmEFuqCmgMO5KyzxKnOeQR+i3EDVSG5Mgx+uxWdo9hT
pw6H1ZXYjmiqJM3jKwzRGFexnKtf1RS1pX+ILkHxhTopMsm+RIrkNvrt/8xMXEEHAMeNeP4lTTwu
QKBvdI4IXmHQBVUoEC4Po0X0xvTFIKAfjJLfgIz5YxIYD++9f4s6jb6Ldp+dn2Xbjl2uzXD2V4mU
IuLKxCEmv5tKmpgV6lPDB663XViGUZ8paMhofqmE10ibc1mbwqxMQNRYBni8bd7y33Z4a+gS9N/4
ylGqCQxbJIKt6bQNX+cJEJfCXWWVAUrn19/21pTs6Jfqmvzn2h5JEcHxuj2u0Ulom8oq336OkVpP
1COStzo7/iip9/rD3i3M58aumYTOP/7+VI3uOzcWP64qMJ3mvyTaMBu2dgwU1Zbo5devhajJDsXq
CqtiC4dfeFX1MF+OXi+WNstJ2sC9xNTtiRYqbxUKKYE/AaHsm2lrSRbKU2WwUxbo7Mk/wWQaMzUo
r/lvFQ24f0wfC5rJyHHqlV5Kceqxp6FK3N7G2lw34cRD+0pxA0MXC8bO50koVgxYmQigHsxmBBDS
PPs9zH1YqHDT/jTzWCQJQ19uKEmxkc4ZmYRYWITp5Vjv6+VDNfFIF05qmCjad/UY7vGoRHOr6Z9V
C04WSeCjDaQoAEXJF5uSUIqg5EvlZn8I/nWrKHIpdW4e01LuAID3s023sVDjVFZKu04uydJscxWA
PgsUNp1ZdA8B4PkNIF9Fx2LRS1/vh1zZF5QDTpAyAyj0KQlP4uIjK5Y7G2zy+EnruUMa/rnjqi70
UxYkqUOJkSXRmGB4DV53mcCeOsPBR5QtpOiqNHHh2OCX/Yv0aiCb2Jy9ebbvXa2J83d46hN+6m2J
S1TpT3UuUSppq0vEK2Fct4jHH6krnTCfrvqzLf4OcfLqpC+YEAwvF/An3LG0Mqeg2CpX1JKeTo6k
aAn1WehQfG5lwbsbqy3gBxDr+7iPvod9Qm+fEbEtH+bldc88MPpeIhh2h51ZhgNq0TEDIgR7bXOh
ShHGDy3B6KuEl5RwIln3+dtvAYUYMVu3BESH4uX4CczU2IDMi7MVq5HwATlunTP3IajGj9tu9EQQ
pO8PegRojMJgWk9MqYDwZD/gmRN1I7w69rVehTe8ijDHjES59jZSCn6TUMv3qq36y5uIKtLr1Jf3
ZS+CjmgDQKkQGYjHlgr88P7PAaHJ67I8RSywlZEHwyx8sC8YmaC0CcCWzk6hBSkDFTlRvdH1Aqnp
Gc4EbxzzY2A6koGRt7hYpVaHqDdljPepPYJ4BXgPwUZnCC7J8iH32NceEOzn9KtMEPZKuSi7w/aV
Y5JZTz/BAL9ZmrR4SYs3XROYUdscKYKmqdBJ7OG3Nyu//PyRw3l8YcrrNMczffz0xWq7XztJnHrO
UzI3WL9R5lAD5py2gL5ommfPfe6tEEH/PQxCSSoBq4Uto5OG9gwhBdEXp2CkOTGE7VKd4lAHxi4o
ZibeVAJdYKtbe3Rkd1ZP50g1NIPWoUytcoD5CvTe5lpDPshfGaYXN8L28ehDOJIktxwMzHPA0s9y
ABJndmZ+y/nImX9a1IWh4mjCyDswQj6tqXxgBNsVt0UN/5NTrWn898THj8kv9irFqM4nwZHuEJMp
0hPlLxx8eLnD0yMPMzU6BymZ5qfLO0rdO6Pxf2McWJjlbXYtg2b7cPJR8UsGkSY3RcY1bEnqPgSX
B590nw03E36M/LzM171g2t9pPTyyMkki90jArc4LUKY8dokrJ/DSUoyWXPVCTSe10KwqDfrahD09
dUhmERGCJvWeif22TRimO37xnAvtr6KDuB0uumA/I0nVAJrYZ+cLphO5WdaJ0qxj2wHSLZ7aY2RV
MCauYpl/i6H6X8KlDuCd2nbY2SOrthYMImpLonuN9L8mNmdpmDwoCWPMu6zZ4RBy7mj2hfClqNxa
e6qQkhKQwJ01caovwCECRutneekOxr7+HTXa5Ow/bwG+JjhB12Bz8UsGt+P/PdYfaUUUEbkG7Bio
ZgeHA+ZQUsqkPq5/7RQK2njo5MzIdeff/h5GXC+YzRA63it4MjH+CjU3bpPyHKJTUkK1QUHc1jQR
Beklu52oJbZh36dnGCYUm/GOqZmDnIcBh1fLE/oHqecW6Jielo6s4TBTyph3SVuatcN0MiASoJHz
I/CaA7ylhSDJj4870QI4vx1HcFFdfsi5xnmGUCYQhvRaJdYyUDtb6ZbhSqbgHJkJGIAJgA7/ujzz
XAG6nHC37StBlpiqP4OfMZf17uVFrYKML+65UAip986hUAkvn4y0dB4XUABxFQN5HpCZY8zyWLKM
cP55NuVzc//9UGsik567AaiBd3v9CJObDHfFdHqsHygH2DTnuWF/MYTenj1EM7XsjHUZpKokfAJY
7qzbOEX8Cy1CJOW2ip0LZmjrnapuC+mGcvLHSvIfihPOhK9/d4tR2sJAYRlYtiNfDZFo0WPBWiS8
4bh2iOXhBEXCN2uCsLyZOJ2/Lv5ta6o3fs4KoJ8bwfvbO5W/DY88hk+VQ8zTg9bdQh1CDqoxyWrW
zWkIlN3D0Mm6kKVggaVtSE6OvIGgwun5Xywj5fCA2WXHvPJN0Ndh6xnEMGC8WgMPm+f+JR2NdrAm
DFUBUgGa6EQdJGMXjmhT86x3CdXl/MeRhoEOgBvCTVFeL2o2AhyLKqMxXgKjfJsQeorI6Y7nPe1h
GuqkuXXoF7nZwpwPBaYaS1pHqeeBclfK8JZczJ1GWe+rY0AVXchj+hbTktCZrZJJVnQNEi5UStd+
z4JrCibUQKzhDoiFSzp1gI/xokjW79wr0gusDsclPWpPVwpm2XfLDFhHGhofvutXvSamzgMFIJwI
s3Pg1Z8wtbN25afhlZHb1A0vPgElzZdxGuMB9iA+y/G3GvuqrKPPTO8Kgw8M/JBWqtOJmG5GJSD7
5VIuLaU4uQqkDpYXeeesCGt43C1kvd15g1KGkTzzx66+0NfHw4dKKORWpSKKjysfjYHU2mtruLvQ
gn52755Q2Cg4GIuCOYItqLR2n6fsJURnlzLwEfhboqqFwoJTp2+CWld0pIubU4G2YWVB4aXpkLgd
NOt59Hy2mAUk8FoCxicp0zt08yYAvzw98M7OAdIMHTQzsLThatigvlUk4Lfc4cZnjz3E4YMAI2+T
oqmGYrUoAicMaMV17qzl3fHi6qi5RIsHPWs8NOJernzJyHvdTmIlYhbvZ4SUPS46VktqatSKImDx
l1mG6CxaIYt63ShT60YVffVI2BqqloBCb70ScmVYuStVJ1z0FdtpQEzC/X0xeFrmFl/ZMJSSP9yD
kxlgWtgUGMQvVsGzp2ioRthRhMft6BJ851xunylgjkhfxYJGXljezm1PxuEKWp6jYBdQ1qMxiZ/2
0rSie0Wbisb0OoW7smMv6a0pc1SG7yptlYd1kRikihCp9IUfDkBW5qLxnqBvXF2aI5ZZm+NgyRPo
ROP7NrbR0cLEcqjSckNK+xBC7Vs1uwt3WtN4v/hO7LYmqNxppqccDCNd/CtJQhu+2ZYOlGFicv5V
3SDFO4daj4H5joSOfLENAhgG320xuMFINNsi7o7tUbV+t4c3cLxuiexjfZNgv3yqNk2dGrsRSmq4
c05LoP3fpKxS0HUsRYewopJqA3L72XS88feHCh1vpC38MX70IOpV+Gt1Gs8RIFR+zxQPYw8Hb9Xi
eDF2eiIzfBDFly2y1KT6a2IDAsHDcBeEPAmDKmKQsO9HSZgP2mj0etYB1tyzC+duGVE5h+rGOPF5
Gez1cJjluZcEYbTovDvNzndj+2RXP4r7grrbHVX3LV4H9WbdHCsTEbjOBKvyVncBjsl8MRWGpYdN
Ud565VArW0xgvinBHgSF6RUcTCq4Av9Y6t6aYysbSN+uuakjVnO9nLNZ/mp/H5wT4nB4zkIekKaP
q8qINiW47f6MQ2cQ1tlV+ItqJxY5mvTJpE11yia/htSvIXHRup7PDCVKBCfFHClbKmHJRqW5oyuK
r+/09wC8vjr4aZ3GsixsicfLKjagMbw6qXsJnmIYC0C6MKHXKOct6otxsqFj7PO7Ja3zstW2YsZ2
TQzRjsv8AVTbAn24BzuFFjLR4iV1hDUWZXuzlaLo1bA94t0hcX7rya09u6rYBpSO82hDw0hBI4UR
LWeHQWWexgtchzUBpy8ZD6hKAPqVyUR4qFTJtFPHZkjmn6I7H5Snk0/lIV22MYwRR1WnYcMlRBK6
MQcgGqOUVhGBUa3CFqJ8On/zqbgjKomudg0M1DfuGMb6gEQvBVX1Y8fB7RKYAmUiMNlRa+y/KxBc
XEmrK4S8C9KdUN6bsAIeamxJ5mgqmobDzJ/UYl39TyOXsSnk6WFHIdpNlBnm89D2SvBFcVeKv5wq
FdKwEX6SQKvbBy/1yM3EJpuxifSK5MRwxR2O7BVcORJhJasnjlP4dQKbaJmZ49UJpUH4XzpEy+J0
R3CkkGCnM/ydPjfD9GILQflxuhjrtxZd9HhOTk/ughjPrVCf1g045wIJU7p81UNMvWzcvzjDVUux
xcLlYx+z8sVVsW6kJx5DOxzlebhZpNAp5BV9pnKvbftt1qJz5nUNYjqDhowQwxmfuceS08+HbJVF
LHQXby0D+ym+qWtW4fWyJohaqyVl1zU6bGjKAhwtewarFkhO+AHPrjDtxkyxUPeHXR7ZNMLdRh5f
da9DA5CT8M5ZzZaBG1B4+NwctmZ0XnC71NFu2IbDqdYGhq9GwncHapmzvYME0W+oehHv4EnK26W0
aLu/88pRGTBLBPyTO34NnAXWt8uQNLtlBobnvhdGmEvDo6FJ4+FIOcYntv8JyybTMK3vvYcgcWHP
P57LdEFzrcSLL0QmcgRM7zY5O+5E/d7oi7LSDvAHNwO2wxASkozLjfSf8UlYd1ztmEVR/kQzgk0n
59P9bOP47Y2JMXrr3mAQUnHCah4k17RbBE2qFJ5JanHYsAuTCmH5UMttSc4K7sqM97sCQcI/R5tK
2KUMTanl0f/dI+L2dVNjWNQBherRdp8sU+oGx8pfOEBNifiMWN2psaZYfvt+xAQhNbPtjuENjKB5
mO0jfIpEU6VVBWq7QGe312SoQd2Q9bhn08R/zBOGZ0Z69NYZIHiDzY07U5FCUY5rF7EncfJ4hhRl
pHsGwQH4KxXU+1G3ha4nUIKt9X77K+5sCdinA88z+EQMYpNzaRi7ZUblTnk573BnNFEbCU7cmAjG
RLemmuRMyhv9aJGgRnZ4C4WBX9AHp6pE1DC9xudlTeJ6c6l4Ls+KTDBfjLNoQKp+P85qNxy9Y0AU
VpJhchlGmUxLlgbT95ZN4jBG392VJW0Qs8sbsWxyF0D/dryHgFi7zj9jXm1G7Kbz8pthoxxmffJI
e9RgllwEfv86rfZsJ8Gqj2VwoU9QXJeHdHSqWU57GWgkyy2GyF9njWFNA229lS9WaZhWgIdyQSI9
22JL+Qmxf07j7YHTu/QFn9c1CR3xa2OuSD3LgH5UUmcxQUXh/veYYLG95WGUmI0GLK4zZX+AqwKL
PL8Rw+uj1QkwCk1e2m1AAQ6YNmO38mkMrjCr2s75rjcQX/5PSPnGI36TGmprcQ9a3+0D2JkJ7fPR
AweRwToXSBiCBEuolRGIm4fgkOZedUi8F3r56/qOrZrqaJk502RsZrJs51APpt6uvwhcxVa8XjCd
ym7fKZ6Nc9NzjiPKwWKkfrY+vM/7XfHMIwD3jbWUvdVVfR8I90nfIOwVKhZ6XVZSWlTbWtvAS/eu
EDMkWIZAF7ga7XCfN30nQLQTIGikFCUM5BwGZ5/ogT/NEz9Mwc95TJI74jggyoTFqtOs2Y2xCIaN
vio/hX/0qlLRVAzsilkkie46AXmHJuAV83+nPrBFtnd0AvBLbQAr9DAcM6LwUjyyswcTccwO5UUS
pdFx9arPiNLi14uQsbJ358PFplgUHS50VcqvtyCd9mOS0LpwfxDZ4Ttr+tacNnEVR4APUQYICVUv
LLjom4eleGLozR2n383xQtpNkzsD58I59QjQCmTduSC0rP3dpV8wVdLPArCJCDCv1hTff97NpsDj
UWb651llcRzBHz+uESDgl/bVgM1+01AEZgrA2CrzZjzM7FEQbIjc88acc67yhduMtuWy9SqNZcNd
jkeXw1K3C1ZBXb1PNsRAIBljv7EFw+Gay/sinUsPQYGtEn1gk8VwhT3h6tepb9hSz2fUsF2cyywH
CpMxHMmye3SPLxCRFaPEKG8PYMk0u4EU1qaxCb1d9D83fjmcJxZDrWRu2R3Gg8NEjx6STGQ7VSGI
lb3KZMQvr23cREUgHoAzPopgS/BvTLdzm+HuB/7+DNWUbW/QqSOvFXgs/NboW+HADvkNT547eBmi
fTpD7hXpMWrqWvN1cYx1exJ1M1f6o8sXdki4RPqY443JWDpQFugHLBy59femVLkqw85cqFl+lKoL
fcjxfl9WawDx+4Eu4+7CeR8jzgVnjciSphs4yHdg9t3BuwPoLZN4uPpeK6a35iHnauBgw+OtjtxF
GN+i1WFzfYeZZkC8AnwXi1e10km9t0wcdZXe7I2l/K8RZRiLWoFvfo5sq4rjj36wH2tPFOVAFHgy
C/PSxNNupoiYQKsG5/MGIksArDr3uNzoA25c993ebocvMMSjaPUKV2Xi4xlrQbAtplE8Vo/8BkK7
COTYC0cW3Lc8NhcXt8Yi3zzs7GBgyUjaNgcd0XCR4sJSDQQTNi9NXGu1xrdbuVbT4GcXI67vY/fh
DywZbhHTSZC6egE6hZNgyTzoZm8cb8QWwWxZL0RKJ2gRUujMZKBQJLpQ967uMdjZTAb5poqTQnwA
qTi/s9nwd7qrDj/blfXa7Ig72FeDmMRmI9A4EKyOUAchhpsDmXRowabQAPWWCIX5ohU+9+DRhTml
8URAXDRZda1ulbSUOn3rspcyYj13aM/O7JeF8is/hvxZOYmfzGjBRCimFwPazTFYsfkyz3F/VEgR
+BjXpO9/paObTQx86iFRTg8OCNXrky98RYj/8Ydid/D+edj8crzb/6H26UmRHWpkvGnRNacH19Og
MeMdwrsb64GLgxrleFr/XSmnGih746rwv9JooMZS/16whTl/D10cmmH56lAqpqfp+KZ0OkwyP8qn
5gNCb+zjPF+XqsnRVoCoVPbFWOSXQYDEPrBj/Cp6nDu0a9sWCb2EVnWC4LkR3lNPOjo1nxkFKMG0
QxRqZrz/TwhzzdrWj43e6bxviV+8ztLCmfcYfS52svU0TBRJdJL/BrxiF4gdUdyq/PNjiWVTH77w
wvCqv/47FN4JWXYfgHowFdtgb5ZkU2Aixq2StWUTiQ63dxrVlZQEAhELBsqJnYu7cp+SDEeoa+dB
UnXL+q0R3xazb80cdGZ4U3ghxEw7ya6q1STf4Vbgo6ktGRQIyYpW68ikRBuvvjnp8MrZfKmynLJW
9uKBgPcVMhM0Tm7HN/uI8IG7tjauEhwCwNQY3ViopUsdLYBUE2HkiJyXE7vA7tNfIkZimvUhFrIS
zabKhWsEAyPq5HQlfZ2M/skN+3Kfie5sEFfINNHOxyGLzCGWOCiywNp9hsarV2sd/p6wTwq0EiB2
ELtra5J3LsFgDbIqig9G1C6PuAe7TK0d29f9QXPCkzx5hMkWqz27jJ6gsBX5tgiZXDV/6MDo94Sn
KWvHAADFw56a9bKAjrYoE+C2v/TB87kuQ5E8favfE9nkhwyjoPYmimPhGC5AJjXJPT1w8ywfifYg
4FwTim7Dygo5JCEb86K1l4TWQ8gfLI7OhBuguHBVC79KkkFXFyjwWoftsZdSvtA/VmoYECqUM/iK
sdic9+IT01JLohKKwjUYg25+BX4rFxhfp2PjDF+9/MmYRPjsxKSuGY89E/88GiytnZeJlMMj6ZWT
3NSeHfqH3F45iI6GhPLer3GrNY52EPDmGeA+35tazsSrA9HWXlekY+jcbs5QTKaxKHDTKa6CSIsx
C3ndAEzOdO1hHJBtjLjeQx3Tp8No7W1c9u7f+v3Z7y7ZoTSvodQDQS1I+d5pOjTcPW2jJnhx4EeM
dpkoTV/nlq2gMAjkAL8Gu9cEq8aJbYtNQP8bT86ERzf/MBRShkXxPM5iyi4oHDYB6dpSPl6bqo8m
zmUEzfAQJ0V+3THx8fGGpewqHO7CsZkqWYCXl+ysPegQkbrZa/NywuEeOWw1zsSdB2rcYrmq6R2t
yYc72BGRC/phnxRGTrW5MgqfoFwMAz0J6ge+wC8XO4ZE+/fDSG+roWPSdGN04zgTrYsDtx08dia0
CdVHI8rIeBA7/sZuH8KtlfcpNQVdMU9Oc8e8laucFhuG4ZHW0aW62HHdyu7Jps69vfittTgQX5dw
EqBie3TEqpmXPdrdNUdiJNNBZ2cKRfDARYaJyaqHdimDx7N7982ixVaEqUF5chU1kzg3hljL1sX/
zZ95kW4naE9mLSbe2PniNr0vawb6lMFzjblnLZinVeyyCq1ba6VkBeuJ65Q0B6flkjJLJaaKa53F
gU3LXHoyxdRZt15FXNV1lug/j85duLOMqIGjnPjaTlTntw+UxNSHEQaTvl9ARhDqeXnxh0Y1KcPq
uNABCre7YOSsQbefuhyKjNgEDa/1flmjKZkU0E9YldMM1vZEuqCoy5HtZBvoXdkr8ALUUtsPCWKJ
BokKxcBrLwIGaACv4jGwhfIPua6YBAZPhWazIqeOwjXut44bEzNwneLINcSN6LY6kTzEpMkaxcUh
PIqZwXxCe0klrwMsrj/ohC+KhBdzjB4nari0J4kQzz+0YZz0ZbTdgmo6DsDSVhVjLXUNOwL8HBMV
nabVi/CgeQCcCHK6edC5obulk+AywSh73KXc1oKYMUlJLdjeToKreQ3zbv03zqaaOHxo+nwJZtIC
sL+femjg5UKQtameqw74J+ZnXReVfBDPPz+aUDTuLsgsEFdNtHdcAT5GdLRR8U2Jz8m7DCAUrNj8
3o9cjhOdvjy+D6E2Abjhs6asld37rkC8TN/6hR2wVppEzjx6OXhYPctFBy1bpHxWbLBrjNS0sRts
fMTg+QJG/beq0GRGhaf69WVKr1OHew5qIT2N5yckw6kR5sUqKEs9LZaeGenK8T8CtjPwyCI+bwIt
P6dxe4Nw+J+LQSGC5tPtyj94CwAh459QF6tg5mX5HmtFPUPK+CGNOWSM78bRLCQ9hoFZwJL/DoiR
G8vmJbw08scNUNzadPcRaoX9lJSXWeXsULKdCkyBkBpqyfYF+JhWlJYAfr+2V7Iq9/HL4ztquELz
9DjbZjz0LEyC08vVaTkl6lzZeWone3mFsw/ghVk8q5QTdwW0XXfkDIapsAf9CR07xh6kfqPSbcyp
J5U1i6q85P8N7q/Jkv8gYE5ZaMKdUUTliF8kNnI6I9AbYW3J8dozlXnJBA8c6L1Mquo6AS3TJr/1
HPNnZWE0s62OzHwP/Z0i0pkc83B88jQCBtYO7qxEroDB+WqcDsz/+zLc7SnkL5fgV5sU7yo47jHc
3+ObCBne6m4inio11QIF4DD/ml/+guPFB+1R/v+8WuTLhls4jXP3J3eSClyrUC/88Otg4a2gTPYM
Wd/n48fSzexUDYVHIYbUeyZCaWhtrjqz/NeQAxPkehznaCu4oS93fLAjlEhdMQALoxcamhitjcLu
WbPeeTMlbCPW2IqvREjywWPD9kT5jtSt9D8XQ7NV/zDFTkaXR6Kyy/gD5vlc4E6q/qFe1+rT9LmF
JNEj/7BkBLj7GKRTRroVauNleaHPXyVK20+Xa/dBsGgLKW5AwHVVJ8ncZcwbT1LzboYruH8uWEFJ
JI33B9wS0zHouakNXU9TPeuyHL5VzzXwfiwrdi4+ogp7ddojtxFdvwiGWB1/VlW9YgSP3XT1BxTw
utJE95ZA7qgZXhbbuHSWucQNZt9J3Bb1vRHSxyY9cS7MXoxEr9CawDcVVML6JJLZeYA8Kr4ZFK0E
ybG7ezPM4bY7kiJpm2b7fky3hrKc3U+jyNB1BSaGHMZPRCmGKaVw+O6F7Y+MPktuyIkIhiXCNk4j
7DEGuT7+awkzCXjndvYkDZu7jsbui1rsSbOI5PCMIe0fRRmMtqKjkJXV0fKcBjGEl7eyVJ8Oi8+j
0ve7U78/nj/YRKfNUygQSuk+F83yQglLdslxIxXJUsIm3grmB9r7vpeuLgbWaYNQyb8QU0m8jOx0
TbqS3Rp9QPXrbD0+3gT5CIJ7B/26dq/CvJ1GyIBceSJgMGHxXNXWVivYZHShLKcqtY+0hih3ZulZ
cj4eNTlu7c8PbyITnJxzEzHpfu+Q0u7KK/oAPP/rCgZY094Psa4FegQCCs6iOBaRUxRiRQ7auLMl
ErPeIlq34qE5wysi7T1/tVOqbJEGlRqKLiSfgd7hY60p39mzlYNoNjDuBn9AbKg+PgYr7jygnUGl
edbUDrPqOQ0i97nJ8GSfkVy2AT0XgkUqllwi/+V0+SY49N13s93WJ/LTt2nAN4AxvR2pqW7PF6Ke
EO4NZEvdRYRfSA9/BzfFuNdtBn2q0T3YlWuDSCYThbihdBE4onpFR7IGU9F9EUqF09p8rtc17yD4
xMgMWT+B1+osdZGgnhtioAfcXokx1lqIOt4YD8WyeugWxh6aov87LJLPj1Eo5h6/egqq28q+9V0b
2plAOOT7NMvc2WCo/7oq3yEK+l2sxWHIKF0XYHAa/0n5BxZ3kRJIZFwTveEU/r45VAIS3oEvFI9c
hmNuYw81hykNsuhrPtAAe2nUe7PJZA7o141Ad8ClCbLMAsb/lsh7i2SPijZWVyXwW10BaxP0zs27
rTPUUZObi+73HjtCHI1GLixLCF+9JHr4XRkt7fl+EgV3CRM/EQXe7xemq0S85lA/rpK7Xhc6tuHw
XaGQL8QW0ZQ1RbEryCo8qXSQVEmquz9wvj0sSsg5agwO2piuy3H/t2z09/6gDi3NG/qCWTGWrvO8
uJMETss4nMQgfxO2CplT1UwY9aWGFRkr+rLlFxLXphmFw7nLksQty1c5oP9DlFlmKEBmfRSuAKv1
mrzYfmSBA6EPIUSRQEbj2Ta0EIVcEmhv1ZuYzhAdKChyUqbhzv5JNhgOBLumkY8x/WXjS7fQ78iC
aZWllf7KUW6Gp/4RkUJUTgdSCtmTm4Tq3NisZuI1F2JcPk/rdj81rv59W/Zic2FH/G1R8NAlFT3A
gM0nQz4+FjEpIB3oBzypg4lTUdVk0eIMrrylPNbFPI7yErBJuUo1OpCc7ZLTpyCr/8NHHUVONnQQ
evyJd8N3oPu2lT0eh7XN+jOIisFwzXTub9teCANUZyOe6PXaAU7uQBDnlR4mSyUegQkhU3111y2G
NrIYrWeAA+61013BSztdVgLA6+9jJE+zsSNjiNRettQ1bi3EwUaPrcOM0FRoZ71twKeuoIKDCKLh
A4JhPemoPhXNXSqn4AH6lKc5HITLjw3LUeVAymPSWSUpWd3xiYtQRuJ08gL1Kp6tw3k2gmonQ4Jq
kVDr85Vs6SaCWL3NmPKRuTzYpvIVYnyVKIqr8iCGhJw31Nfhorb2VmvqhBp1zwe8qhiVEueAEcLR
7zHPQntBWGHXaMqrUt5zibVbqFhoXqAPNpFTCu7go7WJwYf+h9KObAn2cfqVWWv8N4EY1/Sb/5kK
n9qNjMtvUqhBieMY9VS8owhwJ9p/M8U/WydCqM3joS2I3D1netHJrf2rikzPab7tUkaRXujrjgOH
zKyUf+iLitbxYAdx4AHg5uID0UjaXt5NtOuzss7oEZoKRQIYPBrpDKYelMW9vmGk3xfrCX89jd8r
QV/tHKIjjQpJgmiHif9okVUySwg15ZbbvqZ1x8+HgUBIUPAK3U+4K4Mg/iPC+ZC41/t+xcuftOOs
q3RSxbxUVVJdNW05rqlOuBbF0aJsl4hPY+2fH8pN8lEBGbh/EDukSXlZFoX/HOIk5bwhwThtpFNo
pMvOlDUjXczjdXOgJ0qAQSW8RnHC+eOy6F/lFzUvqAPmnAkHthFCe6T6Dsnhp+yDtFrOZ4VD1Yu4
xIxtoNm/zyYCkgaw+YvQqlsZ8t1Y5n6XxMyCvkpIH67RpowgAsFEvMVg/Wc+T19MKcd9fmv/xHXL
eYFXqHVPKYsKMsF7HvqgDifEsItnxW+QSmQDf2a4j4QJ1Ex+faJ+ku1vETlaVLL9sB/fWizGbNw8
5A2JZXKS0p3VZQ+TqYNVttECwAZPzUz2nUojdN/sA9aUql0nSkI4y2iwpRnwV8GcxfzuwSRHMaXx
o9qbkEedgx7OylRg3s2m0oPd9SlSgH/m1IbbjNV/G/MAHpBpMf19CGmY6wmCjbw9SNSclnHJ5OlY
WJqjqXjaOJ4wfDxvw33DtT2hdwA00z0Cinywr3bmb9MM2pwApQk+deueMxEAVbERcXyuxuMSQ8xf
wNG0xAgWJJAGaGqhu4pdVm5skuXlVK0IJ38mHsv18INxa7+NvSpkG7nD0x92aSCaZqQ2J3U8ZJ6Q
4Iq7YHQzj8E+tELLsi1/SdgNwteLAxQPZM6pnaKcRyBBD7dI8z6bEfrzGXJC2nLLYi4bIQ4/T3UZ
Ma5HSHTi/hJBAMf/lAgujoXCGv+WhprMfKQbQJ0bOBKuHi98TKzRCsI3XlfTgsHzzbDwIO2MofNG
iVXzq775KMPG2E9ofTtkwbpSMHLrBO4GowKJZOIU/LkTW6QDGgdjev0QeXuv2Tt5JBzCQDrgkCaR
bx6O/V3InRBx5MDAq6VhMrPyd/Q3cxFFzTZn1vyghyuitEn7QHj7vrb/zOilPwaGcamUWdosKqSl
FuTEK4WgW6hdYr7BlizJmPf1cPII0GxyX7QLxpXNIB0G7qoQ6ZGbQaVOZGJWVmCtdYeki1Ra8gBa
7AowWSzIS9H5NzdMAxFqgpuYod7zAcfMTrk7WVDnnDN006d8B4tn41Kx7SlGkFeyrDy75KtTwEk4
avrpRHvED1yEKJsjv8YPDlrlXxJInNSv68QHTVl3IdDjYYyk6WSMpDfSfueehkgppMQCtJgBBFRe
kZB5DncS6Yb3kS4e92Jz2TeSrbbuQp0pWOIu0+tF1C5wQOF0FP9MhyqdrmfOU3VbQ5x6Tq5LUKWa
ii9lRG9oD7LA5Yqji+hEoDHEbhqSf42ONcBRbRv9YsN6YWY2TRuwXXrk8iO2+h6JGF8kFtqk3//m
wnZYU+PmW5ziuxF1Ihov+KmWiTnXOFBVZsBSDvP/o6T3l3JlXfa876z1oDmdQqN4Axkzs910Q9aQ
5XjbZnyuUohBT4DLGh7dmdhzb1StusiZ8FRC65sljFeXAb1RWzt7J0/gOZpmHxEyMrlTgQ+U8iSJ
RhebgOMLegL3MMCIU3gPSLZjuNfbFWgqjKn87rdjanHDEkD0fTM0fqeB3hKrY+E9/BZzFS/IQo5v
YLtkycFlrs1ThgAyVZauOLJE5nE8u2BOr7IPp/B961gPCtdYe39na4waQ7ZCwEEOXmKz6VAEZH1O
dqB6J7ELf5C7GgTgKJUn1tTAKHaZ8Hj3NCxzRU3dvWD7UWwd5nvJyKZt7Xl74zaZgtHbmkt9w3Eu
eQgrGCBtbPkLDt2nAvg5ZWz/iKhoILiMjw5mWQ75uO5l/Er7lAt/12YyrNISSZkD9zJKZisawK6t
B2iqx2jbq/0TIfAe8zFEtrx3AGt0YOzs65brnHEj5f2yHVasn/uZaIz0DDJl6/xr/vV/xVDCbqY6
6KnuX935PsfLAMadtK4GETZFYEkxjJOjLG0WKFV+XSf7+2wz+y4IU2N4jZ/vyVa3Aa6ODqxSnJat
oJP9C1GYnmD99UL9WkmCuds8SqX3DHfBnVwD1MvsBVYIDe5HtdVPFV2MXHSKYe/0r2EGJ/JVX3HX
Rfs5atZsbfl4Qnx80YTibYf4ZqRy9tGrfSJnzBCIjWTZNGBM35fVGoA+ZD5j0igLMbRwXXdTRBZZ
TkOsI+s9IAlAivG+6WKxgjTXRwotr2lOpyQlRlASJapwnhI1ECoHvhqi8mef12jwPZugSjAJnPyv
ySPOQn677S9NlPrwvscAlQQ+YQZ5TAvPYVrzd3h/oGr27VAr07Fb/2aQ8+UBGxzY4ejCeT/GFa1i
HisiCHY7vdcL6ZMV0Lo/PEJu3hCyX7iZrAqNAc+Yq22Tqwg//3/xqatLv4n/HFTts9A5dTv0b9Eh
9yt2ShtWs+69bBGuwdCgzbVcsg2Ezzn0mtuLIyg1j5IfxHByb2w6/UJUuDpb3yzxx/PylV8thNBN
YZYFATR23lr3xtlanz3Y8iJXwoHeeMzdBqq5nnmnupPqRcGkjciuVZ/yuREKx1H6XekviN/Z6hTu
NkUaHvkhncUPzFJ1SmKLtBqsh4JCexpxqvJAC4UZtXhhHA8FvfdsAloj2y+ZH5KPzIP4DmBRraJM
H4j5VFplT2hmLP4JrZEASBxzFaOJky55ZOM8occOllhYge2s4zuCXSwmZtxIGLWY++7BHzg485uH
yTiwIWqS5Nr2s+4to3z5H66MCMs6iMQPiwuae07LMD6Rj0gvWIYQQzcTdP3t+2ZqYDv3tny0DAUo
LQhvCmwrx8ZTkmAlh4KXvA309lmn+nvtIDCOp5Y6YtfMRAondgQvzQg7O5jAvI2RHCNg2wejYSkJ
7H7Gl9DN8rF+E5yLkTcTqRX0PgUP74M3Vgbp9LDN6FVm2xFMRzjYhRXCU8/5dKJ44nQRXA/7odwc
jUFYzKK1iBQ53xcuCYKLhrp9NUYVluwSoDRB4QnZtOL86H8BiuXHGHTmAOeQ4+/8QPqnKeELWNI7
c83ByCrMWbunpd0uvT1rvy9YNAYskEvEe8aHzo1GlFSMgeiKS0pS+nMbLdSxHY/zWPMT+GzipauG
FEypDglurYsP1zdmF+nkX/NnUuP/15qUl2rIrNTfw+hSoLfxC7P3mT3yFQE4owWInxrCOdaLpAo1
o1uVaOSVUhNELplwjF03XK9jI6XNc4jQAS8fN4FP4Ffx32bqHxGEtxPfRD0D9S5z2jftrvpNpzSZ
NAm5Tvp2HXC5PEf7jYBbRVHB/XLS9A2cxZhdvsr2llntddHYMMG+3N7xw4ulGB8cY8+lYPfPsL14
M7SaC359HLKoqJrQTprk+5r7+WLZTtjxwp6o1APn2B/AShz9rcj2FhAjCNRQ9nQ6wgfocmxU3V4E
rqiUZuSwt9m2T7KXXqIB9yb2LAz8ExmSbrCiRZwENRg0FEAQnpyMlFaYVbSL1LaC9tKYArWpf+9o
dsjPdHaXrgTfZATh0Z/kvWmfNPozXBZQr7cC8zTl666rWKs2+iWvoIIrLAQlWBfV7BBWSYdYmbxT
b8KsISVPuTfYTjKXqyDz8gC5QsGeCNjg5wwI7QBXjacCn7VO7yE0HdWmyGMO7WFVb27+s1Wn9kMW
T9gO+N0eJDD1hf7eHd/Z9JjunSn0C8v/SQbFWTjeQUpDgcGUM2e/el4v0sgo0FCThNrp9N8RuU6s
0G/SIIgyzm9Onk46wGPDe0sc2EP6MzKoT38VqgjQYyn6Er5chXPuWY+m7m8pcio/kC/ldjz1mue1
eBO3qEPjXiHj0+SxEihKTjp43gHKWZtYQD+RAt8YYXceaOctYAfBzGXIILlYyoP2UtpPTqLg7xLT
clM36cfZsrmustqt6oyNd5acaEGhpaTXNhkeMsR9KnNwCVbSNdCepkh35X6YU1av9JQnCVetS5h4
3i9xYiYIsNHIKKVOvMB0zbgWnm48ORl6xL4qH/uVvokw7J4SRCd7gv/bL6APjp/F8TLaUX4Q40eM
jIgpq8hfKmzKFWRMIFmMbOYUmofK0Zp+6JxE/U+QT3ZTL0uJ0i/GFZusgcVXLsYOKfcH85dtyckS
GkLMSzlGYDGIgaX5Aey+lRp0QsF8Wm4HlZjJTfyT5IW4kl2EK3KuwY8rXTpExyyASZRE3K+FtsFJ
gcO2mLG01h9us9oVXhT5fReNDkEqzP16m8LfVetwvuJgnYebWGUkmjQWCtIY3e0Coo9kbEmpmP8Z
1iIbUO2dNOuCydVBjcOb6rDRKmGzxuDD/2d3qcM4EmFogb2VMwLcyGY4FTRXSNeXCse1DXIV6cx9
zGI2OuEUJ16D3JRo6gqR3YvyG2SdyBA+DubEiFNSbzRxbjnMLP7J3R9W6J4BphsB2xZdq1/fBB/F
8U7dMFuuaedEZ8X9o/oaXNyerikQjs56332TwOSVmPS81dLxxaaEBFBj1xIwtckRdW1/C9PdZieV
ayIlK+F3ndlugeAIFkT0RpF/bScD5d44SwodSKTCtNeTNbkBwZRj7El+TcXMOXwlQqfCLsX6iJkj
8qJxfLIQKDdIyHN44uFP/xOvEhVQvYzeLeyl3wGmI0N7scUs7B95Dw/z0dkYDagrebn0EsY7dx1H
/A2Ij4KdAHCLj7OqEaGFrekR0ZMBEAw7dF5JJFlJ6BAbYsxyYSf98yldBpKeO0L+IdJcj60QpLjG
91hRrXrNB9/JIzQgtYKJIUu447hvgRs83jydyl2dVSAZb0VQA2V4k+pY6fDzhNpbMjFBSMSXY9B5
Tnp0gXsxY71vJk5+zNGkdhkQg04yqhnHgVvGuq+FcWIQefNz8j13ZqzEAqvHo7pVqVHdU9ktlFYA
bEj0bzH82Kym9wIM8sv+1vhf0JPg70pQd7H/ZnoSFZkofqJcPPEzBJCYKLWrTvYKJRjNT04fBdqF
W6wsmRsUCT9ruWq4bz3hIFL4xPxsX5cQj/yRjhI/fnbeQ8XPyw05qdQnBMB7bt2YxJmCmgP/qdS1
T6+IysSGjzrWxCfG1WpwS2zBmAKB2Amz2gIza7HD8R+4GSchJ1aveyWl/GDr1lASCLjD142jT3mb
Pv8RfrF8WQ+ZafYQ6iGvF3NfVTCIrbmRrbGrppOYAH7805N/2RN82SMSXCM0vpSS2fFTegQB5/qF
X7DUXjMI1+2U6OdKM/pdOdss81x3QOXG2L5suhgRyr0QujImKu0di5sGUHOr/pgXW6daUI69KhRz
P1SsyPxEwJ1kdfs13fI2Y3xVW/h19q7xgjzALzHOtldVmYTsmtVR7Uu293HmzAKGiDM4gwi3O769
gn7vfLF+f2+hYvwdoXrhZQanXo+ZpO0VwwFUltK1K/DjMhiAaqBLEAmHtPtgm7qydFHZMtx2Fn/k
DG543WtNG2Znhp3fPwbm13sZ1Yy5tmcjfPET7n1IWnH+2U54qiOXhGHO1rjgow==
`protect end_protected
