`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
YMyUwJK6qq7ngNyEOxRtOJumC45yjgp8AOth/G4oXUxDvG7YKd3JDSxbLX6CM9XqcObDWVwwh3J/
EqblB61+VA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jTrfdS72GP2+inVXWkxbFW/d+djuSWiimmeZqu7jMtBg5U0EWu8RIaOUjhY+DTVWLTCgziQAwwBQ
LAMaoeRrV3GVLKCkhyDkgTB+WjpfbJ3t7yTQaLh+tOHDgiqTxdmkplllFIVGcR7hxWZsQ1elpprK
FtzNRV0PoAN7RM6hSeE=

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
XDvdj6WGCKA9L6/Wd6ToL0K8qy9cheS75syoBR3+X1i9fN8v9yYtErWq7C96pFs9d4VprULAtqIW
tuVNmJIPztQlnUDO4QO2qGsEcM2TDe3SWp+vO2vrYT+YxK+tzuuSoeJ/fB3m4eGKzyD8RC8o4LGl
DavPyJcSFbuY6KHyiLI=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
VS/RxRP6GlQlom2noBD0WUWlGAtlBd/2KIQqfDEB3Nw86nw0XOFSZmK6d9CQjP/Kv4JrF51dMevo
0f9eqQlJ14OOwN/3gN99iAoXqSPzAtFcvH1yC6pFVO3Vh3EN7DSFkZG1eGqT3qHHk+0dnPEYhdnj
cjQMAD5pnSjX83m11zLdN8QSRoLlNkkZWu4Y4wBaZXHmIo0W1yud5f8oqS8OxTXGWwGuJeZubuEv
gYRS80PkKI48UQ+VSeQwJ0et8/RQgKUuliSlGDu1xY8oDGNDCZzahSu3f8YP0F+sdBtb8Q3GAEA3
JF/qGWC2065O/mk7XbzcZCeXa9y0G1bRqrlXDA==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
DUs/Zdaaygt1f2BUjXWq5roA9cmX4VcJboRptEEUyKLnjbQ4WmaG5RqvQPluTbauDbf8FIBr5dC0
W2NBW1cH6VvJBxMcZN4XKKniSMqIknq/zvpFLGjP8N5BPGYWXdk8qakisl0b40m7gsU3mwaQTrKd
lLVKj5q4wrpFLvlkxkF0MNAkoH3Qjy7INVd3iLIGc3v/0gj01OlpW6RuHU4Zcz7QMNxvVtpVImMQ
oo6TkF4LsBijPq+W2HydwWC2HSyxte8qomweBlPtrraHE5hlbPf5HtL0HVrRmxdtoKKL/3BWMDAe
UZ14PkBWuX7n5fkpeqXtXO/zL39KSMlegPJZMw==

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
MIO+wxMOH46jXI6g/A8QtqxCNmtyx1Ih7OkdwnQW2HCatcxQN5To/Jt9KCMTgryku7ACKg08NovS
r5cL9aPAoJUE/fqhjIp0osLChUdCZuOsNCSdFmDwKnOUBXTSXoeQ/kpsDtti9y7DlDaAvclgHNdW
pE5ekqV69xYq1DzaLeYoLeIjr1ZQLJ67Ffzqd6JkgzNvTwpTfoMBpkIJAD0pD1xLvQ4nIXOXjWjW
aEFKB78E0EFEWEZWSnQgjQjGd1ouwoJLrJTFHM0gHrN4R19ojSLve2FnawVwqy011UDqERBPMZSq
i3BLXBn9isxh/aTeaglQif2+63ZJuapIXQyzlg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 302736)
`protect data_block
GIeVGPtEz4e2OLj7nID3O/JKMwRoS3y2kJ/F70fRgLpXGvTQ0U+hmyK/P3v2hI7DBigIdkvlPX67
I/3ez+TJL/rO/YcJA/qmg9uc5vyS21gKglOkBJbs+KGy1TVrls4u7sDDEcC0dnqq7yJRPoTp3ZVP
jjIpR7N8qs0OZOYcg4UHeyiy2M1uAYurFsBZU6b5VP9sETD08ftm0DoQ/DSQPBfWC16/qoCzTLhz
ObJIJQ28wZ1kxgb5t0K6Wu2viEbiG1YnJkM0Bws2picI3NlFLmod98hFyZS/ydlIePMW94GQ2uQE
WBZ9LL/b8avMaQrNn8UTJ9r1XyJUJXW9iWMGrR4V/zrkNBwdzH+I3+O9Qoy2tSa1T3NY+Hpn6ok1
ajVSaQEBitz5pJ6K32grtzzCMSKt30+lnNfWa71SXoiQ8Duqm3hF5A7vDqLrfJ4JIx+cNiJuR8VK
VDx8F/4CrnhlFlv0Q7dSMmUQao1PcFvS80iCyoZoRu1zYZMvHFIZxEGeQ3LhV9S+WnR2Z5irQ/O0
iNk4Th1OLitlmjRplF5y9n4S17zb8LbPc2j3IWIBa0z26Kts7c+dr/f/KIKY/Co+Up4REDU8QXZf
IT4MujQimf+G5JAf8X+OfcOjxFLPNVjJWqt6Gk/P3J/jJETDgb+nadBl0Pt868jvZxsJVHWHCwgf
Vrzpr5y81+3FmO18jKlCikT8nRFFA5bxLjyAIOcLxFn38Pt3nIHzljzXqEvO7Mzz1AzNw6QNq9MC
rV6HjFzu8L/YWxekW+mGlbfGiTUEH80fdzWKOABpJHhO6AKv9wEWOB+zfWwbk9cFc0wPZioXU2z2
ECFO0SnwPTCEMqboIeXoH9dZvZkwNZ+DLhQznuUgBwFtLGUqcBpnOAWITWOzc+VdR93GUXoOXqNy
NOZX7zezAF47xji1T+ZlnRRmo+40JMsb3gOMyoOT0FQ5efO1YVzaMa8XNXfa+zxokHKh7bvr2GYO
b5yVuizByGjjnIWqwm5rm/zO3KElJXC55GlYG4q375FCeBH+LCF8bdiOD6hOtCwe7dDoAO2GMOSk
hZsDqQtFSSTIbLLfWLo4IzUHzrLtWu0orSAjBFQj0c+7fsBFgnYkDWSkQo4rKTJcfYsWZuJxvRlM
KAS7BXCvyuiUQPzmCoS/SmmnGBWBU8YZ8TP/WyCGlofH9Fhcn9syhpiNe51OCdyHUlromYwLmyef
/1bYfp707DsM0mzzQuAQyP98yChHy6jk0lY/ak6VK1MRJjXX+e0r50tqqdLIm3XaM1/SZvmV8nxZ
ExIaWBWt4rGFW5jZhvk480ypNzjEpkXYbgPvbITgD8gvha2dS3gf8uQ8s5HKa2NyU7NDdgCFqic2
Be5S5HIfElIBi6DIuRylSbBJt1Oae6W67/SWMM/uPudEzfE3ZyP8vNMfLvnBeAvLAsJMvR/y8vMl
dGTNOm61q18jaMIgUcpigv0+W7bOQuM1LbNqmCulgdwhWi+ZFNs4hZQx1Do9joVlJtbpcQHE+WMC
JB+dihOEdtobFDcps4uC7NKSCxjCzKj+hXAFRuTCyxU85qtAgVCKjRRtiGC9thH8Zx9BFPX1SYe8
DpHPBEDhgE6dtiSCkh1kaahS9fbMaEmuoiVJ3FqRqP14oaN97LfZ5UJKUczOr8jEByB+yiy3TMVT
bn8C5Jbjq90d0Gz+bwHiBvqczYYZZkUX9QCd8/R4msSPLXMHGf+DbeqYlapSrri3H39Gli1ypV7u
CH/5ik9EVisvBPl5RzHo9AxwEKuJDYTaN+21ldHJPw5OaA12LXgr4kM3yVY/N+mSBQjs7fgiSbnH
D0y3ALGSKgKAUcc8s5sFWWpLfdE+i2lVFmC47VKUswrdwn+3ABG3B1uOqFvl7Tp1ArgCv343oR7j
Wk1qLPtij1g3bbeNxrtrXjCIHfe2xSSW4P8duYhjMDFFpYpmndI5GVOSFfq4gsOhv1d3zehlBwmQ
bMF1I2N7VMSYV4396Bc5UXp6G+fJJShXdzFyUeYNEsYt3GNz5hrz3giB+Nmd0dfS/MfSD0zGEHXK
l0kohzgiX7F4u64c5Vg55EkD4mlcw/sHZZhTT5D1DALh69TZLqrwZt0ujY3/3kAFY5p5c85jnGaP
0/xOizyloWgJ9PbmA1SOIQf60TEsUZkzv7q7W6ocbsqg4UI9przJ2zH/cUeC6a5KSpk3JWXskejO
ZkmauRjpm0rvyf+FewcaUDTLj4TEQkelSENK6ECl7DBqQc2bTfRcNUyp3MKcbI8+5s85mT8kXiK7
DQVp0bJOKj5F5ouSY01+5MAS5AWU4S9doKFv7PXh5sCztjHk+qWRzHAMZ36WtQIR+kID5HvQAHMS
XHB6K6R1retku8JQjmVtuKjB2jMinrU8fSQAvPEeMMfqoNS6SbfUBkmVWLP5Zq1L7mZtbhWW7yCi
5i/QKvsoBIWwP/C04nHfUEtnx5GfOj5z8+gfe4l5VZssXugHRFil/+SrBAKIxXHOsOSIJPxnKEMd
5snxlyiQcrXB2S9O4zYwITFpdZ6P1nayceaoLZdY2xa+MRA2/H29spZXFkaUK0rE0Lp7iQDFDbVm
q8aGT09tp0TUvwcuX09l028tgPDnKP4jSEftdTuBslWipVOWWnzzm96P8UCsXwcTr0TxX0PW9q4Q
XEAc9orzXL72Z6+/l6El6d2DF9tMjHSWhil3InRc3IAOYW4d884lRAcBAcifmHKwFN7FKDZp6vZj
pQlfISe7I8eaT9Om079L0vu+J3IMdSFjVktsQswPVuku5zJxqWLSGXsCQqWjN3pUDt6yc6oB9Mu6
5X8vxSP0wvU9Zrl9ASYHwYxsTjIbgkxbqQg0CkdaATI6/6rSiKBG4DKLmIhZ7CEl9fc+ti8WrpbP
3bpfj81spJS/RpgpT8/prpK65KAhDkh+kpFhnoYeBC9WN49yBOY4XLTvr7In5+lTsg/MaoR8HC3n
0lpOJZmi5l99tiAqqATI3OgwCW9IAoqXhkXnZT3dIixpx+NfuXH2daMEzsgXP4EkyEvu2AJGBxFc
7uwXTwanOLFgzZwbMpz4K3RyYFVBpbF2dF7pPzJie3f02+1oOJ1A3F1iNmQcV2+XZ9cTLVVtwTmz
wqwlP6rpr4Yrf28VEamHikU58SQdZiiJvu76ynxgaPVRymQCnjVxiPCnxo5ZygDLjseY/qBgSCgR
ZDqIBjFekvUmVbXIHhDQZ3lc6lDRQLJj5SLjJA3tCYSB1yJ3/pfmJTSsBHdek73MAysYHdHmiFCi
S+euG3qOhltZvjUvBA42j4zoldpVNF9Z+A0/pFOgip7cLCRLcgwa0S7RU0zQdY8ZllOvUKfVzNRn
h8ZCY/FXVd38GSj03v8frPrS/Xw2jT2UetD2318MLUGDBx5VrwhX/n1rwj/xNQTw00c2GfOXAAhV
yNPloZtSIvYmNtVNRg/UlgzTIby4V5svOEiwYsOERQn2AqzGbNLrW6RLd6BDUzRmjusVxzKHc/Sp
iRt7GPesUXh+RBF2+S6gGTPrG0RSbfPfnErhf25REZ3RvwllBZ5wnlWCw3bd2rJpSPnd3jATnxyt
/5vr1QRK1S5JIeF7L3BGnJu4/4k7Vs4u3dvyzt7CgVBe7n8+0ZLN/AFgzYES8L+YccH2y6kvi5V/
znNrzK61kchJzw3RVfGD2Ai1XVkW99n/ieSxaQ12j3I9bMT0F8e5+liptLb7NJVckq/kvHwpYGZm
8ulVEY9XW2rIAWVnI45Z1Bnyu89p8HftT+cMs3+oJ7jTzj4dFsmX080qqUnH4GeTGR2j5mAd4yh8
IMzsuyB42H7H4qi2gkLxG481dPhiRsit/09lbWewOIPEYgqgHqyYgO8ew1TCmIwh867p2msfeRKY
JF075NHtpmLDTDb12f1TjRbWAPiEG9xnSLKru3tgiMV7IJfqHSZ44ysll3LosL4qWE6b6ABzvbvg
uYTTSu6CDypVENhBJavfqnHMnJyU/onjuYo/oyPppWtl4mFipMcI27QJWlkz/0VqQZFQ61lWCbSw
BxQCaSftzMoO1NVCwhd9207tZGvV/OXD7ypzSAQVysRfin1YIy2fqJxbPpRAVswZA9/qhLvtweUZ
IU0xJSgYkbKgOwrLL+Vb/qeX5OiqRuDy3LhI5UVeIeg2/U5aaB/uAJzlJTWOn1teI1BF7rpEKHqG
0u+qNhxc51oOzTR5HKcnY4IjyxL9QUKqRlfaC6BKjOOXY1OhQZ3khPyKAQlGc315ECtzMtDbkqid
6eVkkTWRCyqj1GzNcEKPFjbeW/TmoSYkA5Kbqg4psY8jxOaOg8EpcQ1nT/xdhvvM/CXpZPCuypG3
bVI4DziNYg9SsDKSkJFat0PNr66cAmbHre/Gn9mW9ESAIa5jbzb/gDy5u08T/hUBJzlgf/dKoEIg
FKFV9AU2dm0+ttnFnCHYS23e67dfopBtzWcshiXSsAzCknB/sIe9W5TKCF4+2mBzAwhfOwVH/rlu
BDqAdm1oRpkbPRLzpUl+0edt5UTfU/ax4eZ6QEhVEsJn9hFNOhCzlGcGuCPUh9cEqF6AV8Zpt6uv
6wyj6WGKa4VQ1ji75RJT3IluJRi8+otJgYNymATiYADXsKVaIJPudmPKiXbe4NoCGgsM0te4odrd
1THPtKmzzBwf6GPbqBoq0JKL5FvwewKPJ+hJKcyRTkc1mtXzATLnJWMFp2E+uxC/yD+rKlOUZ/TT
aflHklR2qT6OTGMeUYDRFQ4FfMlYw+Urc1CMELb/q+j9v/0op/6IHXJ6hNwTOwHZZLQYvN1rsJkK
QggpPQjJNjVCI33vU+ahcKrT6J/nK3bK45Amzv2xMkuvgmY/2pw9KKvc5/Fj3TxAqOcGBTPr/FOb
s5AkKZrxL00PQ1NBawovaUg2oX/y1CSWdbjpjjsyeTx1H20Fwe9HPPtOnf/461fmoikWemj42wzp
o/x9aBYPpXQWW2AQDlCv6Nl5AOPj9jJGueTjr25hS8p6+YCJK8xe+OPw9Okukvz64qqfgzQ4XKVa
1G11jYVCu/H8vOTDvVb/IicFQWo4G7Gqe92cr/rENazOhoG9vgfM3FFi+GbszPq2vcRk8F0Lwpjj
MEF8Hr3Jdtpt3NCvflj6EPSHR/2+z0bs8YpqTtEYzZuqleTvj5YAkKNgaIA0F4UEyzQDr+ZhGDN8
yxomWE4AjMrAn4zPE/gCZUviSEwD7iwfbH7NuZEowTxfutqKMnHcx9kpKS6XQOJDs/H0ToWhVrYv
MprUBzeEMcwCO4pcW+WtqMixmGul3AN/B4lB+f4JAaKSxNCn2mmtCBsFwyC9lieaZNb7u1wuYxNQ
PBjpwQ+IyB0o8ys4tHEs0yH3DA0rKN3W85Qb+vZj38M6/R7CnuA1uTBXVMNyZndL2s0w/iHGcBaY
zyvTNZoo0QjG06xjF0rCCVX+yyClRG8x6mznuHdo/QrdLcGxA5fkRc/rUvtEm8hbYp5bz1Oic0Zn
ovnegOtIjF7rCeFjzcHP6ZjOqIBU/Vsbxte/mGZS3o2AKgdfKCn4QpWxmaJDVqdSxaJW4sH/+d9j
Ha+Nb1OEG5FKD7eB5BFJCUgZc/wSJD8swzKY056efj17Q1j9dDvoPAqVTWmP+1iG8fZ+ltWuH9ID
8At7HU+PyC/1CqTg0xnmkg536GcLFzpdrYU6ox4igHkklH6mq1lPKNmMfOTukkAPiXmLyddLh4jv
94zuZmBNPs9pYKvrGzc+O5KbgTLp6ELc1lzMl4+A8c+BAApUAjvPM7Mt87U6jO+6XkhRXBCfs8Ps
u5PKIsiXUKl5Xes7Px0TOFIszIOcKFcHb0vu0t4aTNRmykoVZUlBf1ENlqD33wFlW+zbADObXJu0
HnGNL6Ns6O6q9LYo+91w/+TzHIweTEfdESHLZtXQww8qFvyc+gmX56wSGRF7YzYrhqRQLqAdh/bg
kpj7JHLuGibuK8yx9iR9RDqJbfZNm+DEK/6LvU0QkFNcSKBKw5OoulrvzOv8BR1evOHOIZ/GHUjo
8B93mCRHdb13RAyLFgx0GHjH6k80wTo9q1xlABmpK0RZ3Re+R1m3LfQZ8W7kHnrtkCDNjhjy9+oU
0UfEeG0zXkKW2E02H8FW0oR63k6fgBlRE2GLPhyQFvEWmfd5P9w1ejxBCDexhgYvemEai82n2ejd
qfgDY0txH+JghMQlEirLCdziNoIRzfuYiisE202DX4j+coMrIgAskrsh83h9RodNdb20EFniSHIh
+nLG7NSlKle+3a2NJQWT97aNMlgT1vEfb4IOwd3FsatI+yEswO3U0GrSJpCGLN69sNoWRcqKcb+m
vZJHhVXlyy5gqmW7c0EOLRfLU82fruhFcMzP+1bQZhnRxCqTDmlkQzKg9J3/wXUf2AEt6zIPGHvH
5dpR1eY1sAMpV101J6J8dodwnf1qv4rdyOZmg9FrZoeCVx0K//gX3q0mZESyItpiD37SQ4/dkwD+
XGui1sG/05fqex2pnF4Aw/ygOCHnBgwN1Z/ft+DQ1UZ+jvy13S7UqE7ADfp6aEvcN/JAlhlHOUko
aLhXN+Bes0pndi3a0az5TUr8HGCg7bUTsLTbyWEZnj3PcKRfWBEJMHLRGYR9yIebvDPeppP4UHFf
SAEH8Vwyt6KdcKBhwJTPJymm6R6Su7WmDujnOO2EwCBu4PZPv6/uYslbXY5fh9OdpMVKm6YrcMcW
BK3Gs11FOQPfhqFi8jLE/ebUrzcT5pe0MB3E3rDveXR4td1X+omEOlIsYRswhRRdeIN/oFNYWVWS
tddM9S2zCJ00zugRvEvf67X0dYj6ZVDhWqOPB4o/YFQpjhTd7/u1nYe2bD8+fWAyzDhVicrM+j7+
MSn+sq9j/gTrfPhytQ7/GhibdRjSGTe7V9kV2c5Mww+EQHLlmkZpGSXAY76YSO5Xektvphs/ePKU
MRLXNrUiU0J9Oc15+PXMKlhGARh7R8WBFp8pDVEra/2jgOMF03NLHGyd969CfLFo3rBm5dNgxt8x
N+xZ1UaB8djCZ9cUuyU9/MYLBcXHd8iJ4g/ItWYOQUtxcRyutK0TZW0ZWYSul1VA/rUZPiAhaIaw
gfLgPABQwDpqwPv1KRpiLS1cJiy+/ObA3Tz79XBQYvLfgZ6LX7Ly6BXXIEbCtWYj//ywQThM+hs2
fGFj6A1xD1dP7/+QblibmGOvQcCGHOllCDbQkMXWmFWeSQ/KRfaxFR86dGwaPl1TapCcg4FneCqw
zwAmYtHFDYdCEL2d5bP5PI0oAiCF3NvuyWS6hrmFIUscJ4O5Lnn5832mcOEY4/R9JSS2kIoQ/wVO
ABcze+SYSose9BnmWH4VX+AdVKvyh3y9B6lPUVwmU/QNL2cF5v0CwiYEPzBKXsLZ4gcx2aD6LiEQ
I9Hfl1nlGwy/rDQ6CFs5FOom8jHtcCn6Ltj+pAELP/REaeyw8ugRCvcu8TDhy7U7j+OaQ8a3AVZE
3/KS9ozcMsDsvO8dXLcxMeaKnZkAfbd9td7wL7nY5X2EeqDDa7KJkJZaFPjCMwAJAq6OK2g1MHhl
9WF5LXTw0dtkLo/IxmYOwcwQxJcGiMdg19UE6n3gpg8+Hu3KPzRnLERoJnT0NWl4SigGlvmY/1bI
3RSNa6y+3St3Ii/4FHrjYd+jwuJKBCuah6DJFr0NNltwzsdgpXLlwXvLgITW8Skd2O7S3kMQi/jh
ESWVvbcMN/NZk1hJKZb3reJVvJyq55lRuUODwof9Cf3D16K9tV95tQgnICFzlLoZLxlyCWSaHKjg
nsZxe8RUquSf4bm0974O4//KNnv6ryvCBNwWVwBSiSlTbxBkkYY0qjbmJg3XFNR+f/su/0F9VF5m
aFDwCEKK+it0jM5fEuv22k54G4x7XJGqZ5UpQ9D2+afDCURFpNfexh+0jqgV1nj8M/e2SiwlqESM
iFsbwXHnk8S9v/HNS4bn+V8a6EI3MDa3q35MDTGb5zUNLQRR+m4kAxKdBwwJlazk/aBjucI3UO5W
HzFcyUe0qXCYTEt8Dgp+ZN6snuX3jRcb0GvXGpbUWpyHc42Nj9NwXHF1HN7xCmB1I9FO++anNRw8
AxBb778KRk1oQ8pRUaQ1dFkhOaLJyIq/7ltWsjRsqg90EMtJEt0Fnp8md60G0gmmCzupeYWDfQ0a
GNlOAy2gVhTk1yNjT+I57a6R4jdWxz+Rf1mVYD5UnfBvgNfuPP5D1GY2/IDoaP6xZ5beNVvJPONm
nKEa28H7RocklR7Mif2GXGgUU796CXShHENRRf4fJSWoCnVSYcd7pMt85KFBznNG3elRQ3lJBh8+
PKcJJm+VUEhh2R8+FnT8mmI4CrtGVqPn+o8LS/SWyxz/xA8aXBG0jJgL90ciTPhLQl3EYeARfThP
HDCfwtvkOfnAOj9XD1iKltYAGkupN8vzCLbDenMFg5llrsprC7g/bZaWKDE802NMfvjUDg0OqxKi
zznpekkDYpcXzEY57a3l5wrRxFjVMKOZrdADJNhsPMQ1QBsaHBDRjQF1o3vW64qiHgJL01TLRCwe
lRQMLOBYjKDNWDFnaDo/rBVxPfwZJlR3LdJ8ny2BxpOH6krYEZREfbK+pYLO56UoHK62Yf4BImEh
qoQmL+4xOb2DF2xhwpnQfF60wFRLSVx0WT2ozYclsAEjOko6PKen/jDr/yI3yAbmixAkwxZABELH
7m261WdDYbyekSvlPWHJDI6Vplhta8Iizz5jbqf8uBPK355APQAltQj9o0+qfAvHNWe0he8KaGlG
G35dCruVu/j2B7s9th2ElkHz3m5lTOrAMnIf3q7cqANjgzg8qLRllRfO3mXFWg9NmaU/JnVjPdqH
orLDi6P8Hw185NyLHoQSsfd4LM837smqSLolB5bYVswAUbtE2uKwnx+dzQDLClIhEmdmbNmLDJgL
eZipkvY/9kaNUwx+1EZlvWi1aloOxZZN0nBz6cY6cx0k7lgcNK1B9rJ+bGq/3vDtdzHYa+7ARzbX
8WUcAigp535N4fsvSTXHAyUEt2aUW41nKWEAEKKPJ0xR+Na4rRgFXn2SzV2q+GYalyVy/LWZlvt8
yCTtHZS9PG/x3fu+4mczRjvHD5yDVlMXLNzea/8xeVAoN4Vg0A+AQLAPsA8zrLBRmBvmCB2G7y7a
6m9+CaospdQz7UDmwQnBxuQoavcnleF+7gGhR6OLm0OuAxeM9S0mmIMSFLQUem0Y/2rafaINgPbF
rfdU6L23OsQhzATorAgyt0pdzFPOleKBOa76LvgPEfe7FFxY8c4MyxejOBkyfRic2mQc99EGWAzj
86+fkwZXHLq1zgz3M7Sto3pNal9AiSq1a1BZEza0IG/Em3SrL+itXgNd2YS3VyXsXJXq4elMy6eC
vzXIGdypKzEj4aM+WDxKxIqbdJ+NUMyfYytzVBYtaoL8KvsBfjjQSxsSqvB89zaXXBvfKIkw6Co4
MehLxRADsJ+mpekeppugsE05sCxTkFyalPyrYis49u7kU+xCtb4NwHu5Ro0yH6UIDHtfd0amWKt+
4sUBob4t73tF0MMl134oiL0pi0uGMRVc0XXL+9ez6JBoGwGa2uwlH+nHpMwSA6aKJzYZ0YYboiBn
FYb5srRIYFvImdsbPpg6Qw9SaiaTt0NLp96A/FZS2Crc5Oyfe+nwOq+eqCfJlRa2a07PDsV9Mxuw
TDKvpApEw6+GS3mMXpJr5ETmekLolFZc+A/HqkLIrGFW8NVuypBSdTcNinm9Qj2I2WBrjqsE+Pbp
3y6AJt1nTD6BvbQ/G9Us935TRU9/GHfmZmRBPqyZSH8BdWf6qGPA7kgFnUhsUyTopeeNqaT3V5Nj
BCHqnrMc3axhprcVzBDsLDqxedidPyl6nBC4cRhkM4urTwNVaKzIiUE4RK+rEcbPCqwG6sgPqwa3
DWTKJ7MEPNn0pWiOwVAC8oehwbRkId7hBHU8AUgbc29NeeN7qGRYPfy6yamLMT/FFMHpEmYYHART
Oej0/TcJFwahE4evqjjumLdO04l3IC9qEToZjMOMka6nffwlEcgUAU0Wz6lvza5tHPvkNYbATp3W
QRKS1kcJQoG7Mkt57ccNR1gsHqSmdkL1Ky+D5Dvl1cjd4sKRnpyVAx1zjyXUyYkucl+GaV7V6Ylz
fQNE/9sV4wD8mnJhpWJdK9hefxr9Y2FTYO8bNdNRa8PLKQzBSC2CwarJbvTH7m+fCWil0KbyDI82
QhAJEEq2MKgW0iwDGat2+rqI3soIlRoPsVgJbHZ5zM/GiA9Xo85J2qjHc5sQzzMa3rnTINOKlEwr
qLUOljW8lVKAh2FmfCutGgjaQhZ9qlaAuCU6iwLHAvoHzui8uYjpQqffPGQGz//CxQfSoK4azb9d
wIG3crFu+xSro8tc3dn2LpLr6N6lDjQuXDQ+heQiTJEWZQ0+0bMi8ArB6oREqfRzJp6bigYkCbHR
1kIMQw2A3OKP7vJwccQmUV48467EbsjusNkc2BtGCWA7tgVrMtWTebGSUiqJFYMpxfCdRTF+3BVH
17IRsZZtPXqZ45S8GslnzwpSUD4u0bweEazv86SLbtvCs43oLC1aG/8SCXx+dSwlLiAJToHz9XvZ
THBxpuVUmffdjShmFM7hJg3vQKj/zB4HZ7dgIQs/+Zf5QHkiJwqeDMqG7PTWbEryRAez/PdWz2MD
32IY7NFL9m989hCe52WP8W80umZ4z+bNSJjALyd+sYHpg+RSPg+mVM38O2bQb5uBbk0+geFf+Rjs
oFwErkMosD5Fb5gkuKsPV2LduTpZd/0TaNbJkpaLuKrOZ6ZZnpkd4bjvdWnWljAT6OAi3el5PTxu
OcjkZJsh9Mtmc4GTI7bDAtlO/lkM9KLxUhup40TeJ+SdQHG6tb/FnipjTgxd7y+K0euWtcRKGesl
Zr4HxUWhwVd4iaNrKTaGaaKqpmRfxjrpijh3WQTaOIaBzqh8+fqBX9WJ6P5RHNxy2Ja9wIiK4G7j
n57rF+KVrOlDdcUpIjBqzg4j0SkRZLt12m97kPadJd+u2O/O1naPMwjTCv9/iUsjeyUy5/zZVAM3
T3PlSjPTqNBYO+ciBDAsde0O31xjotBtJqfmuFDv1vfoDNa4JaulEhOOtswtHEeDxrS2BaRJ/QnN
h2CIXB3sY78Thz6Iql5zv1j8A4DHKM1hjjhGetJQMPdyPW3LwS9EB4Cu1VKsIHSZhghgpR66uKRg
hWY9JXvxdkXTsW396vN4MRee+fqDA5yuX5NiWGZlw4L9vQW1iUVULXkoUAuQW224hAw91/KOhOPy
DwvOAWfCTDp9rllvvmXpOz8d1KEoJ1rk05/rchik/FdjysMKH0lU4PwRq3t9ReoMbkF20w36IxlG
32n4ytRqNkRROdhhvLnvqdiKTBCo5b2MWd6JE8YZ72ni/pAuRFmzGmlj5J9SPgQQWj8oKBslUIHs
96BHfT9SXa5yhYcVDj2FublcQyw8ciZRCbl2C1XFUnZoaE1b2y7rjHOOLCE+MJXxc8bFHu9dsdyg
WuKh/Rt+190KPfxtqljYZbga9NwFZajwav2p7haSD0O8in0sujZengNuIkFuVuo24l3/ZnpGwjWX
0/mnwJmI1SJRIvMKHX9M6rdT83cOh42uXJpdBFbC7nQaE8euoF4V0pQd83Lx7JoP28nR/OULe2T3
Ff859524/MzcU1FU4h1PEj9lC6I/A+hCCur8CDhtDJaDoXAzX2P1UcP+WFLDVjmvreIdbYJVgD3t
AUIfFS4Kb4gO3TL2jPhpK6W65XLzyBaMg6MrqaE9xgsuPJxOvSuQnKeG8TRtxS4P7QQiSh8mERma
LEmI2TSEO+/zQk6Kynhzye7dgPmf+U7K9YHVqfTFLB9ih8OpL194Ok6Ur4eR7+JXgaZApqggGzYu
qIUkhw984miTeYTnjwT9S4p4QeM7nzQZ6TbtXCB0jHE/IOgDr61QZzRUUOBCFFMAYadQ8WDfE8OY
NVEaLgRpHMdMA87QBclwSFtOLGYBdfSg4joasDoP5OzLcv5UD4IvzmkpkQogxbGMoq2LHMTdZp2q
P56FjFoJHyNvNHaAGURx/0lP8CyLHnDRaJqLLUOigd8ShadA6eM7BLb3ypBVOrzzVu3JAl4M9xVp
TvU06TIUSdrndret5tIx8Yro20uNlGGRIVuyDPNNvCzSmu+8BuwH5Ng+CVhcexAXZ1G8YYr0yua1
BH0N+0Dv/qkFlw1klWDFkkaRqs7z+0hZbDjT7rntH+y81L6WjVd66fjikSBeKfAPDzFnAirbeaWI
2SshCjAHs87D4RG7agcbJ8W4ZPHsERS16h/rd64j9Y22pOD6FHDF5mK1Dvau8MeZRNysSQXHh0bS
BFqgsbk+C9JZ3gdW0et4Q/1YR499SwoFkGHded5eCvnGr3am0i9zS4+COPuWCNJ8gv/mgvejBunZ
kXHJ6cuiN9K48JGToFfBJ6PzkrC/GbefTgvcjz5R3KA6+eG/O//+coiZ8hbyRRAerW3sHywwGSK1
PUUf9X5kWJ99lFjOStEGad6iqRLyIYX7m6q8W1mG2/yLbUfDRBvRJ1Vi4s2RXXLu+7ZbBUSlYAg7
6VSjzG8b0SE9u3b9pvOfLUiEpyUnuRMBpkL28LgfeW9taFvraJDHLPTEg6/yM3qAhnhTfhpEO/i5
eu7bJJ6480swbLs/wW+TlMbu1UOvGdOObk5VkNmqJa9VCWq55Vq2mfiiuks//MW9pUkinmTHOLZk
vHFgGNzEebx61plZMBOhDFo+Drz60hqd8hNERRjA7qwv0JfOXAkUdOYtYxjYlO+2Sqn664pvWMbP
I8VUAnMvbV2WOvfRESpIdUGNN1Be4qi6z7gom0RtHwU28XboULNAZ/e7wkiMN6BWNJMgYdaRRBWq
hTi2qBA8X0Iie3MTtWZAeVhVpWqCCkJ2z2iCd5XfgdKzJ2BjLdJpQBQZTY1tVWx/ZT5CJ3eQL4M9
/WT+gW/kvfHk4W3vyiffO/ybzn5MHXJ2EzuSH7R1DLvzOxv6k3TL5HV4v0nKEBWOPB3Irk5ds24Y
aoKiXjIdt7t8QB51C8nC8w3PzNL4hhpssHcGtIVvoXaBcc2mBAcLEf+fhksVRK9QB6JrFCTgEraT
p4DV+7bTq1xNARAR2I/mbWTD4a9csfxiwqrYidpFxU29XClYsjKIwa16zqgk/6aZTg2huOIxGrJ9
fNOollfVUUeo26Vc9AHe0ZZ4NJW02IlRiMh3ou+ZmiFcHDp1d+yl0CFoy2CMyxM2BBeGYwFCwb1p
EVnzw6Cz6cLVnH0jz83YIEXttzdUaTs6UgqNc4WAiPAGSCTzkRH80PzB+17AuSsk2T/I0GMkchD/
0bUjW4FhBl4E5h12iBLQV7cs9aBHupKumOKIaLcusM/Rx6Jl2RYcN78E+8AxGPSxFi8EogOavIc6
y/HgowLOo/b6Gt81SG9rldTmKc+cSozSTOd2w0Rs+QSOROIa4CsoYAWZ3+Bc/6I4gBv+SBuCxaO7
I0Dpz6cNKHrbvk8npBgpQJIxb3dedTu7J0jCb7gss/XiZv3fWAJTLv5zsfDxUUb2d/feQWGYfVTb
qtyFU5fONvHqoBV7fWzXUPjrgvSLJLOQHT6CLaiiV36QJ/V0EUS4FiIv+VFfeLVKstA7pkF7gX+d
9YVT/s0XtPa2mvn9ovPnqit3ROg3RcHdXkbf+3r+QX0Bn4tOINtos0eGz5bdbhioa7D7WCranGI1
qZdj0nRAAiBI0d2ntEeeTwuyHmZ5GjuHzUZ4kWgBgfmd79F2yWq7rovEhjPAme4R6AoiGh7+jZqk
Cogp4PMIK/8vBeZZu7ulyAiFPiX1sX7l4nTRNv7UNI1NU+AOCKl9liSJJWOehSaFpYI+PyfrxY0b
APqBXXmSlzCDGj+Kvl3pjdyPXFQXyYF84Pal4X2xFvaZU9qpNuw+MlPTxHidp6Lp995RkwseRfCu
AknHSD8/e+By5aPDVlilT3VVVBpWdaVmiTt6Yt3KyAluyHJkRtKZRwLFYKRg+XbxxSyG+ZbIzY7C
sp/dUbvrHTq6m0N7VANWlaREgjzRCOryMFsczLTc6RtfOdiEItVfEGSj3aWspZ14m2V4kLcsE/O7
YBjF8O+evhsiUqfmBu46MMZizs6VAfnu0sg0BDL8rUUp+zxTYIHGixS18HvbMyptU1D0Q2WSX5JX
yaC/ed37p2z4s9YiU/cV9Lzavk6VzsHfMHAxiwGCiLmGgx6J8bQpCgr+6xmOKRS010Vr2KtUR+NM
FzfheOwrvqHa3QPVbyBxMb97hx61FOx9/jsurC2N4MadQHBI96bnNqUkhPAQ0tgAN2HnUyNyVJMY
fKz34kJuv3RlPJrKbmsZzd3R7/eAsJwan4kxZEFC99iQS3R7XSaVRoLVuSkobsRQgmnhLGs1otia
ajFhKELQemAitoNn7c1YWHF7ksVxeXtLeciNRvmSWVmA9Z11dkgMHbjTs5Tg0B6goSJUvMZxrIdQ
tc9sMwFzGZi6rW2M4EU+OjuHu9nfRG9QOleTYXa1MHD+J/tCtQsr/O9zsnTJUdg3uWWSnyTslzaV
TZYi3484UW8tri8ssSwvJz8DAXaxg6sh1wibLZsPpBhbmuiPaVQpbJCSfTmT/blIj4WDwJPJyBkU
dNcm2ZtngT8S1eAqDiqCsOb/11mh18mEUmkSRQWli9243uCd2ayQhXfeK0X+pLeUA4zbWYTh+qBG
1egAB3zjfAxeJM1qU22KQewFXHVQDEOS5spL5IYWkln4Fx012rinTd9Wmt5azRnuOW75m6nlWHXj
zI5qhfbXuonpxl0oObkpKGRebeUPTosoWsyRrTXWkyd5pzSZgH6f6JwhOu2tv63olxsXc7aB41v4
Gw5piyYG7MOO3AsqEK6Y7WY42BsOD+CWCQ7suAm2gOTfI41MnY/0NyRgescuZ+Sc8dFD+GPmIMJr
xYVZU2Oz9gCAgt2YzcytFSRjy74FYBq1IDCE+Jgld0dZ1HG7NfQC9Pu+2cZtRtCtiqokddeAUbpR
l6MpX9T9R8QASz2QSEjmJ5zzhn2wgo/rxYPiDIQzl8NyM4wBfLdK1SBuSooSNjjRXVLxdGE316HH
nmM9wm+DQhQYthtRc+m8zv7iq3q17NXQfclZdtp/DRah+xLR0wr5tlypE67LEg3rCsadwxEUycBz
ZkLp5cWcxppjR44Ii8WlYMstnVDSkGSHpD4+MeF+lgTxsoqGjyADyEuD0W2v9LphZ9OR866kGQkj
HY9NS+WQWmnDO1b0UCggTsq9mAI1OnrMCxw+6YclOx2/FuX1gLPeWfFhK3ercGulNolpDfprHm0O
KRbHx0L5mBt5sVwzXiqxlKA+V9KxYLj0XTNeD0gNEje99pqQGbRyMkf/0JmW5YVMEq6PPKsVJ6E0
o2dM8wCYDPoPNJ6YGgiSmtnaifGRNxGMiFU9Mdag8aDFlF4JvbqXehf07js6hKr4wCCgdafiNq8f
JsY41tt6k5YeCTZJcz7uLWQUeJLgtm6BovIeCDwGMIP6CdeJ1Om1x6LjbYXjndXF1u2Hx6s0aGak
SloWbphbt1dlQXOUXL1YLJsWNl5rVWSb1sAfuEEjF8D6XAbcGvlYCOqFzhGrgdCodwDX6jvSk6/I
rAK6XQ+Q3Eu2ofCWRQ4c+tl8WQhstXSGh6hmbOUzopYT3PC+Rl6/xs3NiVxTQd/P5ZhcuQxFjKIp
n+lQM4NKgxUP9CxlHXKgZZ463yO+0uWtV7uWyYBVegxxh1EHO/eYjmmSFXi2t9YOUGFFbGV2cVJw
osMHazXRTSU8fUKLRLlQsgAvsF43+UQjxUp+gZB1lFO/Ij+EC6/BfOjOriI8Oo82tkQDciTucW4H
upwXyjmdj8ObhxKb9OdXBxbM2PfxmwlhBFqAoxOQgcXRGckqMtpAIIqU2K219C+opHXXOGOOeraV
qmtTf8PxWMxgSk+jgU4JGHRGiLAJD+8qPrh5VS75BXdyEEA7eVf+lIxalPTbiLZUPvtQa1mTuBDQ
mQqo5+8e1KqU8AQqcVGDclvYFRIdnDg0QdwKZT0GWdEIPBJBbgS5lQJOhJwW+uRPFgyGPQzCaFKg
8s1pJ3Tt+mocBlsAxVN18Ogj/y5eYyr4uhft6Q2ZAw468hFBiVtBow88LiudwTjTRcf+wJixk6RF
6xYYaMbMxriej7hEYZu8BPi/XM6Y8+yHCSzUoLYS8saqfsiqMiqiIXQFkWntsDMK3HXCvYpkYvNe
BF9/01EyDjAuRkCkbIgCABAPYrltDzkmkiCJzybIDdcKGDBhyrYdfN65LfXOO17nWaS0PtUbhWeB
AMVzS3DUAOkYrZfyjn8bPNgWJNcTpMjVMO2IF8rAaqJCDbKTRCGeU9WWefiwBR1Pci90HvhtJkpU
Q/zyEIZJQk8cCE3OYrBt8Yt3ygIL+ZBa34FAWCEprsb5zzFSQ5hVSp4mLhpjpCyPgDtoZA373h2b
w3r0QaPlbWP22d1klE/DgbYXUJPn3HYUDCqyQlMyKPvka0NBdRwJZReq/11+YnM0bH1CtRmlpoZq
hQPBr/nxq6xPQAoMZijC/JNdaReLJhMJqjjzH//n7+1B288D/R5kmbjzYrej/Bdh3x/dHV2r6FcS
eFlMz9+qS/kG/JrSYKQ2s4my5fQAQbwJcM13uV5Ag+xeocbgazOwirQmiylaGi3yt5xjnt1ox7Ze
KgSZ4xPTuh/6WBkskqfE0pRziz9Zf7VTJyCdd2xr5HdzrdoFrDryxqn8sYbfDPfmucEi3pmFc3vq
LaPrzu79j2HJDVOuW66YvgetJ9vuPjF0C3uDH/ehYFqrfAdK3DYq+kvS7yarTokvaliFY2tjYoT9
mcYCl7gwkL3EpZcQaMoeJFsqsNLfHqlws0mGFFr9AnLkJVLoYAftnfCeEWgXpY5A5CCW/2DXboCb
9qk1mSGfkBpc2RjjEmxOTleUN1AQD1M659J3lXGONmx9shqioCRgHZLbux2KsmIN83285YMxB9tM
PvbaqiAb6Kt9PTBfDKKoUOHXNcpw2+lpw1T9pddAUD/mrHFoaRXerVcnb8pvxkEsgWtOkiDGjbAv
+F19HaWQza/7vDAExy0NFPyDF0ceXNrwvo51+gi1XN1lhleXHy50wA9KhX+RWBJHskgCJisz+jn8
VxHt2ZiqofTO3cpMvtfkBhAaqnFN0rCp5x1Lhuelx5oDBBzjOoh5Ld56MqHAop+zUlPeejFK2hL6
QpxIy6FuVjpVzDSdmgy+q51RDJMDilXRaRX/DGnqDkj7S+YJkq18ydGVscFN8JF/fZKYA8a1lMtg
OO3PXSJUmNBZsU89Ex8Szl71kTyAhHld2t4ag3KNKmlY2CNBEtkbhsfezg4t3rgDuW3OVuGiKDGu
ICcRvrl3SgKgErkpw3LuTkrdS1M5DcXxPgr3InY+PIHdwX9LG9PWZzmJ9eJototqYd+C16eAGqbh
SQjHSJdn4qLZHK2I5mz4oNm85hJ2ek1GKuekYqwNBN27foVp/ZHbs/mSKpYmXQgFiRkrKsRnT+vF
k46Mjnqb5tX+nDEzXBo4/rf5NKPs7SRDui7TyKJOCLTDfGypfFM+i8HmNUQk/+ALpoUVlu+rXasl
dHk1mMySKQ+yegWSH3TvLNUF/tbA3W+IJtrGObYqXPBAbIAa7pHtKfZeOH0P7Cr/DT43FTD9+j6E
mr9nID1VCxslMVvZFjX/9yC0Xt0iY63zdYDjwJLeXKvZxBllZWqFao31t20jeKI8QVQnYuekrvil
coc7SyamvifCPk7j8fpYag1k2fZocd26za8eDGvGitbT141gzfD107t0TFwCFtmmOO6eWVGzazQI
NIUuC4bIwSuaiXFHpROIP88+DIKYq+EpoxL19gruIQi6f6alBxztQB/qnEr6CHSuVzKzdPWMRJ4g
KynfhVpNZh/F/WkxVPLW8RjHWYTepitmET8837TzOvSf6IxrUaLCoOGSSf8C359BYUrKOmZlR1mP
5XXWdNuroJQXVizrdkLHNWwYtln9HQIJJ4FYgsHNn2O2p8VetCg+naThpeutOj/5jbXho3m2FB1G
7OV162n+0zMVG9Xu1zgjvE04Akpw0nN7Z1y+e7hW5X19qacjQJ5bxxpRM2BSAUZxZYlffKkd9RH0
EqAeE1bsKeyaBW3ITapDMEN7y+tybwt0QmIYA686pdhBIiUrBBNEZFR3R7up+zhC2VP0FEDTDc3u
MuZlpDH8UR2OkUrYomBD7tSojf5J9bUVM1yGM6ENbuYkUKSeBVP3JcgGgtIjRh1XgPTx7kV5xGci
gniWRiy/ZB7cim8hwYeOhvyLQlbz9cZAsM38Td8IKS4Zdpj/NvCV4RoqgKh42D23wXhKUq7I9/AN
1crAqVpWznTA0aSmNuH65UhrI/UY+6D2ItF//N94hhpqHYeImrTdLT3/Htd7O189UfmU96IQlbMi
Bp2VkoRb/qSKqBlAlv2mJ0SvboFrsvbNo7TGLKPZamAgyW/0KyvLbCRe2ZvrNgwfS5UsUn8FAeFA
JpWVSJqsl5ptdGhSKWk+s8kGiSuKAOnqsrFhKnjlv0lya8MZiPB8nD2mkYef3PCdcnwNLRf0gXvo
D3oZKx9pHxlJGXXKp/HAJF2Jhls3Su+l+uhixWDREm9DaDGWZzA0I9CpPAUaIdKO8Xw+t2rDItck
hbh+MTIrmwJP3S1LjXIRbOHkDb7ThCB2kfxxegRhsqs9haWNpBN6eZnyvhCvz2nR+P3mHwLGR5UE
GI9wg/xrLvoKQX7KGbfuBi1/RJ95Ibqdu1yLYU2j98czeecUtjXnZ4zfpZvFJd9BbY70P1nuHXMZ
qjg22Ax2IPdD4N+riwjl5btS8fsHmliJnn3b/wMfqHpqCHH9hX5yybuiIWRkNP4k9zprp0867q21
UyQhX7spe2JoiryjRJBm+UdLTX2xEbNSZA1F+/ESYJdOnNILgg/E9nknJxa9Rq9yaV6MxeFVdmp9
tggyQyTllsGRAFDMTCyJGIyP7Yb/TsYcVVyuUA3KTYuOYWWTH/8ZUILxSJk6OrE3miCFLJFc1fQ2
i6cp1YbE5Rb58eGvjGieyj3cEEQIhQ7blW7tV3NNT/ftJZwC+n40ArdqObGJ8lgnopNdBcwoiUHX
S046OQBfXyIyvQrd69mcDbRfmVVuK+GCOxytMAnmx58lWRcWe1eKrNC9hw8ilkdOdJd/ZlkfbGLT
fWF6FQnJdDXJhP3OCC3eHZLzKdnkx4E6NaT+6cob3+jI2PrtHsAx9CafZAqvdmC5dMAZbwu5ORKK
7CyII5WWt1vQOKzHkPKL6pruK/ZqhrDe1HOPBd01gC/fScXKyXPIAofLWyinAY+ZKNkA41J3Zb1t
wljMfhWJ1e3DwpBuC9ZQl9k1Rhl843YhQQljyGZYpARrQAuS1wXsSld4wRNyJf48AYCG9lk5ryzb
BQ1qAWq2UmuugH2LhCijbHffbV1l8GA98XvcOqpURMxwDtJo+bHjLesSq/Fg7wTSSkrSE72aC/ox
2s2PXERZp/7nsCR/3MiE1pmuAkAgCC0AyjDy+bZBseTMLuwglp83ljrrbLKJLmsDPXrCFm3m6jbA
hDpjpHroM4V5q6KbiVr3es+Jg5mftDw3I2jqKRIvvqziXronPvtht+MC4tujb1SrTMHnVakieizb
wqlCMxosJyBCAvOYjeDqGRcsU5vLmTWtymy9E5/19oYfe8qQ7UV683xn2pIXa1/g3TR3PL2IBBbz
5XcWUK6C/+kQml25BlUO9o9dFsSniRTQZ04K+I/r6hAb7mr5+4F4nmraQvyksKPZRB7Xs7Hz0pt7
5ua+h3puLZoH8elw/kEarw+TKOhQJYawZzGfsB93lFPcoTnMArlQV1cj/z6cPgRsmBaHepeGL1Nt
EQJaXn6xQST5hTJbQLBhEjM+7AWZXwAo64y0wmTmwKKjf8CE5h+ZA992u+MT7mXMOcaPFFKyRPMF
y7tXKXOWGPcXLU27SLWVPXKnTGXXS9+Lxf7h62uINhHj5PSxtAcbTtN9MW+KiiqWABFBhm+0gPp9
I0trvzYuWLAxzp7qDPTDcpF7Xwn39lwbEtgvu37NmCjSyjuFfl8+V6uPyU5RH1WftEoy67opd/tz
2A92EN7XJuhhSG+5vIA8M71f37bt7dJG5XT0tNx16aQF9NvdhB8QQ3vzDkSQ5oP/DcKr/2r8htD4
l+6P10xuXOb3maHv8l1EEOdmxWud8/E01UhVEXQdCB4e4A5rXuUrAySJYeflvtiRpS5QmArC96lU
Od+munXXk1XPmkxckiw9CE+A6FdSrdRCBPXoJu0FBpdgz9CxrqvTAZI9aGO+AP96gUC0X1xMQiAS
DGBhElNN2DkGjJ9MYI3fJNkjutuq5P7QMJiBtoWPA/cuucyfYJyj8/tYdhpTekzWIL76aBmS0W0j
tVRz9ODYzrJl22H1P5z/5mt+e2cb9DrKcp2GODGP8UHi67vCNfDD81cPgX28p9d5CZE3VGfBKEBY
uLEmDB2Swzdd/2Se3L7cjMz+IwTYJgB5/LJg0eFWpfWNebxZka3nG0J7wql0x7bYol7n74oAPj35
CFT2XCY12DT5+UZTvemSn827OGrDGLxr8Nh6TPMEDKK4FvC5vzMIwOQo0xZr10Sg7QDuL7qcU2KY
0wENyUHZMsw8NyARaEOANw1MsJKxOzpX0P8oKNPL08p5hRvYzIeS7CyIhHoZsFGW7CIbRLJws86a
qhu7YDTzzXG+ChyuzEpQdu5RwQU8iFCPr97OIENo4DhCvL8q0iFtIGtvQKKqduKCuuk2reN+Je9S
gSRmSUA9HX9Jhn9pop3RXfANMLJvkAZQGpovKggVD/SmgQwz4LvJAZ1ZhWTa0J7j/9IAiXea23z4
KJIoXU+WF39VCQ88l86YmKVe4+wk5MUgGRUPiIs6flTVKlieE6FH7svBVNU/bX943qdKxBCeFTlE
WOPtEDGrdQ5NGAPFNSx+itKPTKMiTvOONRuXIBsU+97sGeBIuI9ISGUe1aDZJAwkhptWJH5cenQt
P7+RJnd7s73YvgiypVp09lw6alvhpSBiCu+iURVDX7sCrq/n8ASm2/O9m04MlU9n0nhXEmQH2Xmf
9oEWGH2FAvBb594CX74frZBacaKpV61Ff3MWRZB14mVinJFY1GN52OTbhiDUhIAafB/ZRVG/Szzb
qvENR/sjEWCrZFoeRiYPp4kXeYwTV1LvMnrG4kC8f9kPxMV+E045dunRQNmLeW12h3IfO2qDvjPl
D84Gfvllest5k62hYnaLJ6PU23y62QAhpVe1PD+NH/FCIhzWCDbAqD2rXUF/B2LmCbacx1iJ2RCT
DLp5/Q107KtaaseutKzOmZdjig0XsTaJcmJWYsCX2QrkdVCrdFsL8+mfLPJkuqzh5aGUmEpL/kj2
oUO8cfp+4VH6tgcUBJ/jsBr51AWLWGOeiESrVMFgL4Qik/4hpWphk7+9P6JhDgO4Ht9qtUfQ1S6p
yj1M9ueCTSl/9tS4vCOc4JmoHdLcdRX7sWyAJIaM+ZMz7y7w2Qo+yKXrgfyt1nhlHKSDlV5FcOgO
YB1QpDIHbMqfA1L4SGb9ZsAEstubK1jPj3jsLvZma0tXA/wSIW1Xz7hKoxAr15zMn8PAVBehsrIF
Tvc0UURGlUJ2yJUJFTejol0yj8Ketav4+8gh3l7n2KrKSc/H3943VQ4qkTqLNq/nxurFbM4G6R9z
0+uPJNr+1It+VoSsmxY1iFzH6gyXy6skmYZT9muh2nUR+snSkloFECgq39iCiiA+cFS/gOv470zU
OIN20MwBp/CX12BJjVrmLfYvEJjJpkXMxoGxG0hS+mbXwEMhwX7MuBR57rWobi0n1uJsHEaNids9
k+LXJAcnY5WRliXY3iZpaFjj5wF6D0NtJNiiHz+MfEdorCZSvKIBdf360qQWO/9AM6flHyvwUMrI
Kx4Mmsh73kdXdm9g0ELA1miqDN+r5pwNzLUceg7tp0b1b2yK0KTeZ51oF2Ihl8crmJbHOsH/JUrz
P43A+zOwTc7TcIvL9tR7SYPKTV9sjfn/vJB6eEwVY8QR5LMPEJpTeWC7zyoQ0jzv0Wxxer5o4B1O
ih2/DAXkCqdEchIv9ctZT/62wbJ9HiU2CKBlo2JC3xLYWKJm09BV0fez7MQGXmTNaHSSCM2hiSpG
0XH2fFfnR6MZFQlUImWJVxVDu6bmdbjguilw6UsTJ92aYB0rw5rt1Bx0hOrmL2CNUCxYo2Sz/LSg
H9yZr89vwrPy2wKFMk6ttb4/D2DxOadSH9BkP6C7IXOUEU4lkOtxh0ZKvJ7upYEn/WiTu8PDhG+i
tRJCW2ac2hEQxde+A5cY84fwY/SFNZ1XnNbmiKWFgDhZCa4ZbboTBcnm2yzj/19BOIzXkq4gpnAO
JTL8OxbvLSjRNijMRIxzfO6cIu4nZxmdAXFNzlHPxQaDxgJ87yEI0CJ7uy50mhKRj6Ywx2GWIrmJ
YVVxF5Zu+ApLjely3BP5nDrIYvklPk7vYOcE5kcD46nXQu+dO6vP5tjlPQiCOwyxh3P4XodUUJUO
+sk3UNIxSpNfO5y3uP1zIP4ELO2fdnom/vW4vmDPeYAICDEqRcu1iOi1xovWRctgjVqPDWodNND5
HwBUE+0BwGnWurrHRM787PuCH5waa/pBu3advJ736Kj5v0TgikQHZEb0LfnLF1CIukvMUdHVmuV3
jyAf70cz9Snqp0JmgIH/rYHb//HvoX3bUd1AFEpP9iUNWvZuz/KF6E/djTH6uPu/rhbwtXgvt0W6
MyPPCAncs9ugBn7UTLENpiENPgOtv69DJ+IN04O6rwg0Aeb105EKzGP8R8Hcb09hOBzV6fcfTNNv
j7r+w7uncsZ2l8y5VNrLq3+vXyBmcKmND26RX5i6oxVwYv72CFtxoUa3DgqEqoFAKvVyoxgCfd9F
4Xn3z/TNOf7mOxp9/MBx6XVyJy0Njsw091tMb5ijtACy0JV/ToRQQGOe+DbzfNgsYgiqDCTuB80D
sQH/qC9gsj4cLs0OBxdHEgWajZCak3MpGfsf0bftIOVfuinDDjK62IDlm4Y+jBowcs48TsnPPpxZ
3UHSkIaUmhr9oDcn6+Z43DZ4tt0cxhdaVKU9JXDpvfOQ4waU9LL4Y2+I3vwpiQWymvCiCQx/NO5K
/iiSWb3kHx7+Zh0p/O0AcBrRwTMcTLQXQF2o9hhQboVgi0zvrGUH9dXFLCeEOVSuAhK7Ve6a4IYH
GLcPISykwnup/gO9jXeaFYMqYpoO5OOb3bROt8wa+w9RRvKfiVBWe7ylk9ma7XOmmREXabOdYNCH
bYMOIqP/DREqmDMIRf1XBKPPRziMKqRdEk5Dif8sytSWQzLpjc0WUexQEEGASASf0hGjUloReug+
5yWwO+QqRR96ostpAiMQzp2K20lEkCk5/58IBOJ6gCtYnieez8j371x8NlBcOQZiOatUWIkOwQzZ
YdjTCtkfahZEZZmLU9NJhM5bh/W2D7iHPsNrouuJYHNVNcCt7lJNhF0yo2+bmAyd+VfwBXo/453S
elcl0tCd+jZ3XTklyh1fx6Jd+IBMHc35FgjZZxyubt7vnaL//eRMFanP23c5p0cW1NM+7fmT+ZTK
uAV/inEOONXTp6Smi+0WDyFG0QnHKwoxIHGzjrJeGcd1XrW0eOzp3IdI3Kw5Dak63EJb39sVjRz8
VnNbdZ8FxUJyh4nE6RvvLBIet+pXGdRz8a7+lIiCBhR7a3XjMkdU+CsgFmERJtgRBBpN6LsJkeNV
32XFKeYvTTMLNgiyZUNKOUMRvYEn7KzPaMydk1qmG3MAQIxvBa7olW1AidZu7mi0QQnjp+GRmkZj
zjFTzmtisncKHTToHsiAN8logMaZaElLcAbeCwI4H0bNCfivGRfmaQQNEtjEDs3otfcOvEnGqPDl
X7h/UuCkHioGgGXeEp1kwuxyVtNzZKVeFizBO1zSIaP00CdwbVOhwYQTMrN1DIXYxgHovmiaIPwN
JVOQMPLfH9RMyxT5LxDTgSecSzpalHGtOL+Ku/Nyl+G/+ifS2y0aoAcQ/+4deVpFKfvPOpI8Afsb
pDuKV5RIVk78WIktLxD7Xd32DV6pgUy2ya3U3inHqMK5qMTW3dPUnL63dZCv+saMNkdu0hINBCZf
NNk3Qjazw95nM8bNGBAEB7O9Po3wXDbpWGAZpn3H+NCRN3+LFfXAs9E1Z6qqrvHxvfU0FLPufU+B
zXYE/NECom120WY3BE/AyRf0NJN2jSWn74nNzDiFPvOu3+xM1nEkq9ZZkQ9Yq2Q91DmMR6/qQeAc
flZ54zacNUqEvzYMW7V84O/gMaeLB+nGPMYUCRiyo+Y5kxAGBrNbO6gl8yRgkpCzbsaDX3TvSOEO
auDbzWVYsMZW8Rp84sVtPqoPmO/6iI5ohUbmN48KtnjUPMDJEri5a5K78KPVQVgEQJcBaAXPYvk9
EHFP3CjFRGFuyiXiqLtGtThYuhQtekJAJXfErRQBPyt/qdv++d5+8cXYfaVVDfLecYQcvkmuFmAU
xcoMuizEWGaY1K2M44t6bUqcyx9PsP+7X4pw4B8mZhKdDREhTjO8JyU2bjfCwmkF+8kdkKiP1exP
bWg3Th15g9cwDdySsMGMN7xJits/RJg4NIg5iO5KpEdNC/l96WnQXHTUPMwv0DZQJbH/VMYYW3q3
qlZAl/IgLUZffGUva1kzHJuoJTu9gLTYFf5OvI8Qsz/BIEDrxbHT0HqfLzIINnmh0uNjuRgntBuM
drApW63H2vMpzEMXxuzD55xgjUZYmjM8+RzU0cV/KAiCf117ZjrOek+RN5AVl6AGDtfq4r+9BysB
7UIWjTkVdE40X/PeN84JCSyQkqmvPGBU4KyYVpVgz1MdZ1cSG8pnxV6txQGAG8JJ7vOioCU6oKwZ
4ygWtOL/R6fuIn33dXbkY5H4PtqxpGgKHBkwnkhbjom2ZaSHVbsNEZmT/WpxgGn2LIkj3lPHyXAc
SL4RIqIq3i+PtMo3xKxOzlKoj0KXjfqyRw9xV13UP7FbMrAGjfHn53F8dT7p01NggqmWygOuLIYo
mYR+FZxXGL0hBNzccBAPEwa3YcJAxdX9jK4sTqMJu+xuT0KRunNpLs+5LCxmrUpGC4xZbr/ICGyt
5UEXqZU9xGdChb6n+l2tbgvbrY9xeAimJ8Gr15HK6yWTJlVc2aPI3U+0XbY1u8LOZp7bLjtnqQ42
f6+2hax0xkboTn/R3z4tGqGRzglMyMqbd7jCa5E5FSqPIpgHYRX+xx0Yny9+km3hsuV4o3M67tLZ
INP+bkzFxrFqGPicQttWmprFc8dZhdq14CP5bRzYWbpEvpmI6bvE87KC3zGDM9zTJsrZnvxuEQ+h
HyzHSMe5mwaZ1Lg5sdU/rGb4qRFlMuR0lZE/K44qS6sr/hMq3dF3Gaqpt+cq3ecqBDo+RiVcTa+d
OH/L2JyLZObvTMzs+g8dsyxr5GLBmXTwagxt+PTNxTjVZf6P5hj7L8u3m34b9SXwpDuZatFj3M2a
NWuaRcAXao6Udx39+L57EKZIrPEuu9dV08ESb2v2FO+3C+liICBdPqH9EbLJWUwd1N7TaY0s0z0g
PqDhKtBJXw3EbbWaxkT/97kfkY0CrxF/K82qAVb8Wy8Wn3DjHkgXJMPblCk5aUsJb75UkjrVVZvT
Hqn8tkhLO4TR1JZmwJgcCcTUh6FwBNUv2bupn0agLRBIY8yffbYzDw2KcnkZyVhXp4/cmCe9Sh9C
UZJNndQ/OLhxJ2fTzbIVbNHZH22MPc8jo6v4TzGlpvZhJkXJnPFo6cVKqmOPwwbrv882uHPP5reD
h1M36S1gpd4t+ADOzW/o92yXzMeMUcgTvnEzeMnLavU3P38CMBMAEpjjTQb7sizyVSLH+P0h2+/J
eAplP4k59Kfs07A7/UJhlaZKKDSTaBFGlisWKqkO5p4YJ3Bb9rfGgHk6HGQ4n0Gzh+f/KVrp9HgM
Lwxx/c0GfeQY66vKIozqdktKsT6PiVLMuFhl57Zcv7vMgvgCC/2k6iwyvB9KE2LI/1fF74+RXvr9
UjM1B58fHhbbFfvX85Ds52ZCjGCEbsBXbvb3Z6ETb28CW809dazadINI/3X2zXgqadsYvPu7SAM0
+LB1bUwP9IU1mB6sYy+RM/HSIm4JGOGUEeTCbfAzMGMzZ4D4hoviIGygO2+J3BJFKExc6oIqPY6k
KgcGb1JKWLcPz1m45V6mFxuhoIoPMZprOfdPTbGxycKuosd4vbD63h0usveqDWXxZbxYiD0KUnl5
R14JpzDfY7Ffp5+i8ztyPl37xhItjNmVCCAEoLCFCJPdebWNEqUVhYvZrtrQnibmXNbu7XtKgisM
T3qw7r8s8QefyYfZGUVfOqw55lnO5hbyQWShotb0uL/VHrDIiLd5FvdHwLrNnCVCAexm6pYR8d4U
OMMB4bt2qiUBwFurXOS4oN/yGzBzfsbxSQ4LSUl2kzVJdGCSiC6ir3VF/QUQBQIm4cXGh0IBBBVE
Uo+UliFttAcgxz9zwrkTfCpI7PGw9UXjfOCUYiPGUNUFUH+R0RzV1xsXao9DRVVYN2LEdZXjz4kf
zFs8bnNu5wH1d0kV19CmnDe5YPiu4BCHooiCn8gccraooSuDg5Ec+OMrXN9ykPfUu6n6VgE5GYPf
F2OKjmzQWIB0x9CM8/swPqW/9McOMad0NKKGiqyH3JwQ4aIaskeCd4+AaGiaek2zL6NzltXNBURu
m+LaMy091bx+6hgi2QxDIBJq0kiSlMJrMx7ufbUgj0GOFRMFufbO90QHBtvy9LIBUMK8Nv2bfyq3
sdxKv8hFEJPMPv6DtUWgNiQrxRJ5QyG0X1aQObIgHfcEbF68KDBApATDAxGoTkKqHevyLEh3yg63
r7c1PHEG+agVgQpSMnbRSpbHsp4Q+wDCz+L4qKdaKPlrI7xrRxn8cHyvc9u9949OHPfiX6G05o/3
xD6IH7fNwayWzZSpTmukc5HX7gdou/BMsRjnpphJtBsm9Rc2UiN0nmHfvLy61+Ns5k6LejVydtNs
o+4fECSIhratzVUHJBExQUkyiJHqC4AiKaHB/W/QM7vWBeMxB7tS+5AB0wXez5tHRKCqsLDMZoiR
oeWgw5VonjRBujKbsm7zrWcBBIsCJpu10JQxI3huCWjMfQEUlM4NkmFLbdntbR9LYQB8GWddazQd
kVCUdI3V1qSO2ALylegc0i7u/rYoHr1P/MURpYFpRs5wvD17DNl6G5r0M9qjNtm5l9F7YK83dU8K
DnG51u2G2aMyrrxvXWjihuno2Ip3nMkqN/YLBaIhOyDbL5tudIUnHCOl1XzuG/Hael/U9m6YW6ro
L63znwW9ulBMfNDu2H6VgZOQXmHhfCs2gHPV6QeDRhd2a6fNEjkAEd3IN3uzjKWwDWqwCnZomdvv
Q8IlE6EFpSHxA5Vec92d86lgv9oqDaVSop+2ylUNPIB+UPfNV9yclpa9r+OQ8CsiePy3B7v4ggSx
ifUtjsdMudsq5WbhTnYNgkLXr1bjY9/22Pi9hJq64nFCgZNuk6QNtbjtN5PmwCXkg7jV6jlcGSzi
+tkg3t/hAPSrDbra9lBSZhfc94u3iJwPJTt7HYwzi37q/psMj0J0XFxLLgb0K43btCTV/2F3LI7+
DrBG/KwalAAkknNTgf2zlGHxQ6qnKBWPL/3Drng+RVYlPHJVS618g8LGlFs19ZthI1k0lxQx7Q1F
IdDyX90MXZJh30TGFoRBa8ydM+SMHd+EnHvWZnHTjXAN4ZIwPZYFg+rJDIMjYmwu4Vr0Du5mPinl
XceqzQ9IJzJo7PllSu+ozckn3p8llkJrN45i3OhMD1PWm3qUkX9LFnm4H2ZtdF5DqQr6iYdamxkw
exsbaNOvPMsihziOQaKC02Z9H1ETt02S9/1dcgQ/mHtWwasOgJJCYImoUik9Tggmm4hqbqY9C0SS
UmVxUytUbYswXyfytOhXvz35dmSwMXO88L1dkgnyU1rDJ/647IlV/OzClxNEbw4SZXNavygFLxgg
heJpxD0CmDitgUg75NL8+6K8vXDLoW3S2Ym+YbP7zDEsqOUd4+Rb5bw9hF8kpRZmsuyLO+y/dkm8
VhkAnLKBpftoMQsfg6ZEZeXfDyNXPG/IBcpm0bX7C4HSqmO6hgplJ6Xi1FGqJSLGMwISMHN30jsb
yMHX5iFtkcrLyG6fa2GNsjPM/PYPDcJqxfPIxysweXW2hXPNMEPE4fQWl5SAJUt66fD7AQqThvq2
TRIGpGbsP65NqH5lW/thRXFmvUp78c0fvUnv7mc/H+BWT3dloiA/8l/cIIlpn6rhhj0wigi446FA
gAS8QJrW4nl0pViktHGDKP78tPZ7/hUQD+1Oqi+AAx+4x9Ic9Mp8Su9Hz+PtZO/1AKN0PeEcxM2A
3FOFNNFiBE/oYb4iEjW0VUUnrlhHHoHRLZ8pTNHaXDWnkV+fDXLEKLDacpwc5PIw0+bBvIgoR7d1
kRsbQ6RLhu1FsZpZGGfe3NFVUoJmz9SPSpW17GK41dEdTZY8kVqG6RMzngZufPfDtQAz0Yc/eVnU
4rluYyUEO3PYX0H9x+c2/hv/7xYvPJoErMiNX2BM+SO2UXlwuWGsGEPA4zHEod87AaTS7ispxwUL
rzo9jUYtC9AS6RuRSdQlyuNMU9IbFo1/9ZV9MBJfqb0PQkTc4ZvcEL7MA2YiVhJFUs9kH/SAdAa/
XRBdjdRvECEBpN7x8YLPsi7v/8sU/+IsqPu/qQo24p3yN/TqMKNr0NmVSxssDhaHeEHTF+fc+YSG
EvqGbRZZlZp2CS+rFojDN4SYoaJ8qBLdefQ0A5Soae8vPXp1JEBNlIkW6c8ed7KTZjQfZaBSnSQ7
CZx32QMn5LS6ZTnUU70GiAzeopzzSHiaho13rRmkybPMLyaEjfZ2+GUN+56rSKRYqgrK9BmJBPMu
+HZJvqU6ZT1MSpC8ZANYja4H1zJarhxHGXDgeB3TGCTI1Lj4MJq14y2jbDYtpWzS925OcQFdE6st
aovuw1gGoPIn+EV5+TACfFDZBuct+Gac4bo9AGbqFPwjs2D2Q/PVAXRjgN7wTSeMszKTTKc4K8Nk
FKk9ICiGp3epqN6ac3km2jzDWNDdgFWictF2z6kQGjqnTKCzsAD0SZz8DndbiRhRxQSMUdM20vMu
SyaRG0u8pDdTpiO2r2XPIcrA242GyNC0BFe5ZuQRHolC6xw3x98THXj/ChW29Z1EcUSqkYNgdHpN
bIlvC8Nx6ix17ezO9K6YqeY3pPrVUS+mxm5a++8adxeVjHsK2aPG2jVyrRJk3s+pdFnpN2gDi5E7
NUPoNiPqFCNwwCG/CgcAEPVScNUTTKduaK9h0Jy+nJCGBi3m/7OWaefcvAzfS/GO1hwiCsc1rp59
ezqHuGUKBapIdqlxDQSPqTw9JtHoSEYEv3y+ur/y0lZZJyAHTLiRQmhu8ZuBpyprI48xVae50n5P
oDLE5kHUIjnqy/PtrYA/A38FbtEVQj3QgG02W9Q5v5+0rPjpyBOaumIjpnNFRPPkUwbu1lQ4Yz9+
u/VAh80TpU8MtsC7l2qrT7sm7HfCqkMNK77KL0SSiAvV1Pwf8YyoLY7QMTTNBogbbX28L3n6Yt31
y2EWbyTlrdMn2N5/SLSimHQufRTfOkaNYz5ZjwM1VkZGatdEV6my9Ah15Xj1SX8MgffKMns6eHKO
84TLy5p+4XIgcoyUbarHUoZ6grm8FcXqOOIfjKTgb4DWBTmj6Y+2WsvlJkQGL5jY94IEP74rMSNX
Z3eUJzNRI0aaPmX7ebkh/5TkrUFz/w4pe2wC7HpdAEs/hwDj8Rc/wngVav9L+bgO3RTwJIgwecQE
wdQd7ZJC3k2MgJL970bnfY/JRKwdAG4TxL6lyaxXxknVlH8P01T+Dr0chNjivJzdw6lrNReBHZbc
ZgSIZOoEdSlkYGBLgVi5VKWavpyFA5dvRfIpVqbWb0U8Gc6MFhRPqUIZI97HCgT48+7p1tVaz5gX
WzzSn0v4MvI6cfOHHDK4tIkgfUGfYL14087LH282wErs4XwP8vHK9jt+kMvACPSwr/udQ4FWpCZc
6GrYx6jRzqJgrHZMXEp5qxahWuSyGq/dcnP2tQMmK9+VP48G1IwHDFMKZWzToJYFq4Rntva3h4w+
ZUEqFm99gyDovc6IyAngd2dR9SQaAcCvgV/ZJ6ugWKW6FRNujz/UAu894Lb1blOnsZk1kNiCuqa7
psbG6M+QZyjA+aoyI5lVHZ4aWaMArjAecYuEpPuJArBiGDQihYH4HjD8k0969VCNSyMPIRn16iRK
A87BljmNG0WE5y+7ZAD8ZnPrgEWFfEsPPI/SoQH5eG6CP2rHpUZVGsY43f6PfrHieCZp+uUOq+2P
y/2JfcfMy0tga6YUwDX8akun8rWYMpv2uaF7eWC0rjcjf2DZbxo1IVZSet2veUkumQKQ71VNTVk/
8yw388tqJIs1vbJ9SDGMGYXeYn+6+2V9S8mSFpw3Sw254edn5mOSTQlpl6LxrHBVzrhStkS+T81y
fS4YaGXIuBioC+WkmS3MMyOSt8blg5pqFIpdJWL/TRrNndr+tV68gVSWOCz2ArkIhMRA0WTmZBKG
YTT8bYWyKfKAJFoehMkOhCgpprT3dDY8zyFXQveg/TErcyfL26eahot9D13DFzlPUpikxPMbE5X8
CXs9gjXQ6vDCirOUmi+s0QnaEnl4qpmbIiuJrLFMNddxnQyR2xBhxaRzMPsQqS5xzhgSq3QUBruI
Baz0T2+Xt2rW+psxfQoaWCk1MZMZ2lU9mvY4P36B/51yooYjmw12DdwG7VruCFy+Kc6RCzA/ZhVR
+i7hniBX0ARVBlMFBqNz2rqL5DOydGhoNdX+8UHFuXT6inVXj8gFSGJwO+tAP1zcQ/eEZYSp8ucD
L7d2IzTYfdYxRL+OdkgXL8I3O/yHsWfoQSz5hdel80oTb0jfIz5gwurvKxXcMAYgppcuPT+AfUNk
GX/Q3zDXHfcJEauMPtjZH1ZD9g9bUxqXkb/ybVKxh/onlUICSLpCguXEQqHFPBMKkhUmJvOkU7FB
DDtCiDbbN7AA8M9H2sgFPc5spArJXwzeQJLAhGVqMth6KZlHb6iIyW9+T96EOKIiMoaYyKDdDG1v
e0JUbKcImDpBomZZl6GsnOWfDaleLVJQm0ANP+2SW2tT7SIeVbw43Zsa0qSHIcODogRH7vBgr3te
SYr/FcC3UdQOg8QyPND8qGFctCfC4Hz9LxHKYV8P1Hc1OKrdKIvrG2LMEsmvWW4bm1TpPqZa3SWV
VIxBOWpEVzKCwA2yJk46b9q5zOYcofCLhNbSb1Fyq/bOqC/BVXSJwJ6vBr2/zBwvUrNNINQN7u7/
kq47yBdLBzflQDOoKTv8C3+/XrFdype6OP52SC61mhz8IiUXVuczIPyIiiFc7U0WUuGrsT3xJ38V
zvJ/bK+0+LqvDzDauBkSGDLyIGohvPWsBTs1QpFbOc2kkoR5kg2MylSU00O8aD0ZHzGRyJa1+LvB
5sIaL5WrnBkeFDlWod8bkjmVAB8Bf62JVA+YucUBkPAcooG/XoIyyl1G/wtBaLlNa/FAYE4ZAwdy
vci5xjcdZN5jSXWOGBVVXrjHye/u4NDsj1RfwkCqSLXHUuBH0aP0XlUQoVyKIBq8YT0fMcocV3d9
AVB2cBUn3triz0gWNBintw2ga0ABkmN7VqRmpEmGktadYSvzzBaO1wX0NoKBDspkViBanpBZ/pcM
PbUrO78txZkPt1+FQnHgA0LNeAUvMsRwkUzv8KN1FRxUr5IHsUcANrsg9LgS2YZMx+bBFz11vxzk
maY3tjnl+IrS9gF8qZY/pM7GHIfyQTMiXtlm23bcVMTESndZDhgP3b6u07QxycgphCk5SWnMYs5u
ayJuDUmWyVEn+nxdN6wg7MkqJmTazsk1l0MKJyDtEOGYt31WtRtNrEKps6uGfEn3kShJlVXYA7By
WQhomQtaPZr/OYWpotPV8QEBBUHMd4aOPpIxMWlG0zC9kve82v+4Ce5PiRnX7aDFdPLrKp1u802S
yZCcPJhg5cHLVWqvUbxybv7WpLbAPsTfB9cKFGb6BuZ5CZNl20HqEbnmre3KaKvM+4eccEoq1TO2
aptlYAG3VFKHYIGMuBOEo34RskkJn/185uQk2YJ+T3lkjUcAsvhiGtKHIfApShA5J5KTJmE2I6Kx
lcyFO3nPg5o/mQiwZs/c6MMFJ/BE0trLW/KB3VvDgj8R6cz7DPM+VGFsZqB9JjPdKjIaHz0kTCQr
0XArf1lqptuoHJpWdJAl0gMNR3FMJNJhb/PFQbdYNlYaa+n3SEepKZvN0eYawnhwxNDdLaNO815F
y5LnOmjdMuEVJyJR3cF5uEdk3CoUlP3rG6h/1TyRMCtOteycs1Oy+ClIxpb5BvQhGYQA0x2RuRNC
OPJ4Ata82kRdkQeSD/2Zqv05GUoniIWbnJpB0ycd8Lgzow91n+oYMNg/uaDKm6cEZnPC31agL+Pb
wx2RvqLkjQ/L+glcSKVwdiWfubdFMZBcFjfiher7na2oa92wlKKg7fMbgkFjVIJ4HeehMrH97RDE
o0bevqbYjhj9Gn78mrsvWiMvd9q/lA0ESuIe39bOpRxJFMYtJFqcWCPvgXHDkx7l5RT2g+CGiWrN
c87NbLn9bEioUDy8IaGm5afzh40Rnx5zfnauRD1D/nC3QfBXtIzsGBep/nkvZAkcX6OjsEfB5s71
bkNSTaGUqi1vBIf/hcMnkHc8QgPPpsLtpC5lzsfyar+oKo/jkT8CEuLPY6RETe5GRXqLpC232oHa
WcW1PD883eLmT5WQ2srcI1eHeZYwbXkipRqURpvqzFZ6YZfbmlrrfiQS5bswvNoM/tv8gSy5dqLz
5mD+3xq+5eoyzU7wRqKOuP4jyArs+I/6z6CpOQXc/0igncgQRjfQ5sZQqBMXYCHTuA9HdBoCGsTu
Mhs+npraEe3hHjx4CwXpHFNirqB5Xe1AicnJrzgnu+IYLv0OklBfdBa9HLanyvFeraYk852nWzb2
sfpTGPcvZ2VFupm+mxwfIkHPBn4fnog4Cm7vuTs+Bvpl6VMeEOI8FwKLNe+9a9WITJ1ScilRvWtg
v8jCG5H8uY5Q/ZQb6SstgAY8p0MdUH+SkjY79W2xXTdk6ZHyRcnI9U+rgiSgWOiAaJcOycLYbVxI
c8pMt0Vp5ANQwjqNVqd2Db6j05D5HvCXv1mmaXasuH32f2MRLnMy+WgszeSE0wxh1IyfYGr1j7Aq
A6RTRhvMENp3IBVOsd4SQT5+/Dg53sM4ZhP34nNs8ecOLLH2D9DgiXETxIH49230mLqAgRWTtHHN
hTcGocOINHwPM5N7hKE5SvAPTJUfQ9YOyTTRKhcuDdJ74iJ878IntX7jlivSDUf6x7UqPA+Can9o
PpU80UM7fsAAcf/a2RoHBvq7PFLIqlTJDsZZCwc0I8sGYQ4c12kY2dD8EykZjRnBNGO9pmtUqS3O
DpWmZm+A6qA93QxVlgESlmMA8MNfirMQzHbknczWvNWG6043gccPCyQjniLM5mFRgIx4divW1+3h
0FwchrlTuo+WY2fyrDP7yjcbnM3m+usisvTJxWxqAgrKr9i8ohvVxROhViTJyWjh+blN7SCiIV8M
XN3MPJBFKbVlxy5SSglz4RR8Jlpxox0IgLb8BEYJRmRlWVTszUmD8XS/1SwbTUKGmgwCjcNoGRYi
iLwejtNPTOBJhazsFd6UN1+a1h82NGTLplEohAfCXDiRxnZiwBLCGsOfznqGjhaK3rvfflMuoN+O
mtdq0m7kFBhl3ASVKi1TMwzmJ1ohdPtlo0PSnGnZdXyWryEEkE2NlDLAucB3j4B1nAn3gUc4vN7d
I3pinvT+F0Kq1n3ogQS7sSacx0iA8WzY3QcN0H/gwYo/bMGJk4h8v7o7ZuKkC+PX+X2/9Ov4IlkZ
YqFVTSAO8pZZmjMs9fcGsd97T5i3OB3iopo9ok/MemSefULUpkJCN4fAyvMuJQXApCwZMcG0NrTm
zutlzzDVTyRg6JFYCd4wP53ojXfMGgYaFwhOqyFSs8c+eU4xGiJQ7/M8HXz6GRLibFUsvBlqt7Fs
qwiCfYg7N6bmrcAHrbFkJ/uAta/20Ht1TkKu44x/JxC9ZSYizC4p1cgxxofmpEnMhOa3HVi0/N0C
gsY1kQqZHqnhmYXsNymh7DsNpFBqirV3mkyVbM2mUCFYn15taIqMS8doW2kRAEZolcJSWTGvwFcz
Il63l63pXJszWwHCFWK9RSQRWpD35NmYDx+fZHbG66nBDSHZO8ft9ZLdfsG24sZG2eB/RQfYcLwY
DVYUW4bMCVaXVqph/fQNTBEUtoLEvQw8O3Y1P1Il37n/8XNNOaqFFkOgCS7SFLBh0sLXbewz2tpF
RtI4elqoWjAa3ylsQ2maN2xjyGB3cZumfaZ6huir1MUNwowDfE36sf0IEFyO1bXMJBdI1HgTkh2+
ExFiWYEZ1OYMf4jOL2PqVSOk2ZLkMjCk3ubDlW6lPOs0JiOcX5vytM11pEKocUByFbxHJWlrW0rd
6zsICwiuKkKgBdiwy1OQArgkLRaIwWiF4UtoXfy6yXvKJk3rXZdMnF5yFZBfW++XVXoy+rpqDBsi
Mytebqs7PEv16ABW6p9xZneYumYBBC6v20oUJbg+xQ1DwlAJSoBhMSj8N6IVi32RlGpNQdqDfUIr
70KccDZyB74QNVMHcno9ChCxzSBLaGCMlx09+4CBsaa0My5Binx/F+sUOAZpi6Hceur58EO9DkvO
Kwm+xtDS3M+bduN+gcG/HPmr9rbJukwbj9UhTY6XsF8CgPopw9gDbfnDhijtpssTgyZ+Ltk4X20p
/2P90uJHKMDy2xDw4lCvScpjh7T+BcCrwAhHPcG+iSN6R2+3BQvY7Y+zp00bs4Jl43rOmOQVbuiD
OM9aCgSL0qFVBAxbGhoHEI7Rg6pnh/l91t0LIEeuh9iXjCFRqjwy82TtmI40VPqE2l59GkRZxj3T
j82GT7ewAmPeO4VQY+aSEv6UQDhbWUsWF/hd0TQGX4Kxp1es+bO7I/7q0RrMWQ49w36QNHbOdTcC
8yRmABH02wZJqNl4sEhzlO+45Zs/QnvShLiHpiA/R/AsCJ02umy3TUDgC5nikPaR1HeSpNVYXMwC
zgmic39oS8yWleeMwfNEoOTSqqa26NYLFymA5PzfoWO/BTGtgvXFW8BzZDtzTB4zcqRn11Il2Ndb
qEyRdanaXlrEHopaSUqjHYMTx1HaNQieIZUrTzLBYABRX+58XCBLuNphIxdjUhHXeaT8oVEuRCdu
2tvFNpFVS+OBqXBoJX98Q0h3oCJPfj1El6InoLN7h3MB78z2nnUxrOoSfIncoYSzx+DI4WSKNd7b
9U3op2L572sSrasc62Pg9xGeBHi2Esp4oWnDgGG/34fNkyDNgiTQslhaECh2peAiYM2CxPZ+QShA
olPAymb5w0Y0qyabtENoRBCp1r7DOISR89rv0ejjB5EKMcPMMikP+fRyFjMeujQ5dQ3e81fvktU0
iRyb/m8r/4Ky/OEf/1X0cXIruJdoAS5bWiTvAejcLhngPivFdipuGpE7XYs7yZkV4Q/B+gVj7S8c
RoYoYd0Dtl9ZoatF4x936RkFz+8nxDdcoNwXtIZRBIsUM8LgEWfe7FqQeJJSjHV6zyT1hjSun6or
0D+QfEcA3uEH3u0BIz3BDU9fjqV5QJ5DI43hnqr0nJlBXjkLtu9VqpsVxHqqVKG7eLSA18DlFy83
7Z5enzErPY07+g7s39GBTaUzEuy1V8OWcw8neODxi5YvtK9P4qjC0xC9iIT5eSiJvIqx2Jyq5Vws
f+Fy+A/BdsGlZEKv3k3a1T5J/fwTFt8LHRXRHxI3/OhJVjyi7K6dShSbgufdAqfDI0mF73WxaFkq
xJLZbp2Z/li1xqXccUp6e0Zzk16IxM4B/tHiYbQChYxRjv64ciLB0e9zizKDMrOTTLrJelv4v0Iw
KMZZN/T19M0mzkdQTYkkazbpCENQvKt1aVYdDmGroy/8Bax9WZECVHXRzVf2E+TKfVhMHLwT5f8F
O2+9u0wC8Ta+zIrvt6nr8TEn4I8p6/8JPpXIDOmIHiW9MPiq6sHp/6VVOIzEhidFWpMgZudIDQEB
mzQ2jjl6nh2iqroFKPtqRAV1FXml7zQTNMQ9v4kR+YvYwGeWRABrPRuvMPdaFOE6rUiOUBZejRpR
GRI9pTNnTS6kw7YhdRnCuKof+RvP/B1wN5xa4WKykXqm05oHEtFbQ+wBMHhxkQKwfgrWreCj1H18
wbVm4n5INkM2dBtYnLpGT6ZIRwryAMkLEBfVrawLNI2HBCwqjZQzYhbcVCJXJpVyYj9aQKzx8gat
2GenXr6bmNE6bWEtE8O/faku5OjVP/09ObCOEcdQNWe9kiOUxkymDKX4gDXWN1QFrm2UtF2/iPYR
iKLmJE2yjROG1abIG8JK1wKHUelFC1YJx2xxBNVHyMv3ymGWEurhh71mcG5o1cANCXUlXAZN1pHf
lErCAIrxkQWnBBNwBM9ydkNBDSt90lr0ldp+B6+QKo5bzLANwnoegqA5GykwiCWumJwetrnJXjkK
f9OQEADx/y1L4P5i+HyWexsWE0QJiRRfYmOlHMDUR8Mmqhl3vU1rVjFu/9C7uFXP5LjmfEnfYJz/
SZS4Nwnkegos33hVqnzE4DWjiI26Xb2dzoMLg6jpg9YTBiB3D33hOHxYcTMZt9cfpDrSrIhNWplk
yWI4qkYqxi4CWIpZOs3PkrYh7bz9fDA5Uzi6JRA45egZ/cdwu080r47H9yDPwEb1UVfCuWGbp7xe
7G1DtoR0ROJcDKOaAFpA1qfj6vhnw7UagUBgEpQuUMvDWwyChnR+M+n/qjer7lWlCXXBmeWHwW46
Pgt8tjn+ybAZSiOYUR26x3+JiJx4NgjYzNHb9WT1s65mK6CCVZK8u8NUb7h1wUVJfAGZmMv9riWn
XcyNYHUpG9trmDsO4ks56Mau2PJyqp+Br0ivrLZPorBbMbso7A+DA4OCrk8r5+NAENiEfT+IDkxG
3C++6ZSct0z3RPkea46VH+d4KlYA8Oj1S9SghLSUGR+QXILK5JnYQHz3gEza8Am0wldAmt8m3hYN
RVcB3XpGvFc+z8hpaAQw3NMpk7umbWK8BKOIVjEINrHjNjWaVmOtoZoN6RpFKe5XmXWjOnTAAB4k
Ur8zyRHxP6UkuVwlGO7o3TAgPwqNeLYXOdildVpYgO/j1g4KEGz5YLzggd/NxS+ddMJUSFQT3IDt
8s61W7S94yoBa6PVcvOAqt4ZancWUJCJ3CoPHV6NoH2sMFKHNIC1cmucy2Bqp+ZDegpzLXX9Mq12
UqUp4No7+vU1cDPnUN68KIr2vrq5zgqzTaOS2wdBF8v50fG6EWkoNVF+pxl0C2MicGgyUkeOWWSd
g/7fRvTFjCoXD0G56O/rVkWl+DvMYExahlOs90Tbs7EdjPxLOvBmyKfySKDVT2E8DBidl0EhVlfz
BFHv0Pes5DgB7KKxIJ5fhT2O1fKSpMDdOTYseyV0OyPCpKo91V8ab2DMlo2VDu3sQ/PpeCVPvrv9
etfydZSJH7u0ekgXZtjPBSO/lmV0awFHahVlmJPlWcVD8jfvWTDHaGdAtAebK7kAAGTJEKt06tnL
Il5rYvRQGYwWtPfZ3fnaSFxqK/hohIDOzfrOUvv2YNxublK5nrO4CUxME1NYr+wKesxOBA/h2JzK
uS7hEq0A0Ox07+Uef4CSjkPPpWJ4jYtncn6LgCLU7pT3tZwrIEZ2dbge+PprdGvwo51ApfqQDo4b
Viq1SyIcvh8ruvsX5ChRYo8vHeALmPz4oxkEvwTS0MF85h5qHQf7FaCQQsPJyl/a3yB/toOAYIRn
a2OJtOWgozunXOlZCwyaQOg3GaC3eIuyhmCMXaF4jQTE/YxwWU5kPBtBEYchbsoM80BTbPcPzHaO
2pmck414yvERevHAX4oks0DYwZ0McBWr2qWaj/I0zZQoug1C5Yc0CO343bJQaUdV7p0ro0sVaFO4
kKw+NLM7DuIVBTkST1nfQDsAfK82yfGjL5FZa8bByPAlWfVEmIavCRbP9jWgCdBMbUIcR1amMNb0
l147tUmXxyrWfn39yqrrqnje9uF7OnnqAoAtca7eIcyiXkvKGJItzDiS3Idet8sFm4USVArq3hCp
qjtX+me6obmU9J8VAZvjTGR2wGY4zeAvzoMHdSRn/Rg8nwxor2rjdvxqlxuu09EB8+5FPQHwYtNv
3TKBnpUsljvUmS/FolOnUJgsHYniNCROQiZn+W4rKXIBJF2DjpFDUMsMTbEO2+Tmg+a4Dh+b90v6
CxgDRrhK9Cr6H6P89RgDNJ1EFG893exx9m2AxNn4n1RQwngpO9Cc8iqk9PCjKOXQmz3VSqLPs3fg
MItpv0uo8BnDfH3EyxgJBqJz0TE+nY19yzDWwq9AIiKtstelQwhYUammlHVZhpuQr9ttAYsbAcPc
WZZGWV7f46ZHoYrPqRVkMFJwt4cEk8bOuErRyv+cEEaWInr+R/OfP0IO0JbDSlZ9Lf55Hc8xlsG7
txSeM1Zbrrtar/Ddsez4zgyNfo98T9BMFqoIhZv+MjIbxu48mucMS+Cf/LSVthEpqTdWCIwjEL/T
zjU7z778Nr1ZvPVkc7iuug7e7TEh4vJgQT5gq1wIIGbXCJUfOD6OcdJHg6uee/HXZgLwS5SJ89e0
ljc2UkxmlfpUCBmP0ngFJkIaeKYiHsKkzP6yKhNwT+OV3WKx0GBMqSQWsJ7P7X7jN2H3P8iIgRGr
Jvvw0niIaKvSqyiVLsWXsG3grOgUsVwp72jZboQf402fNyB26q+lYhpldTppK2ly/2c3DxBdYFNh
uNln6NmP42tUwSYQM59dB5v4Z9pWw6j3UoWTypJArCHoOFjkfXVbYSoI8ICqcDgIDQjKkmuGoObj
oNp5fXsh1LAgxrGvJ+d3A1JjWHobftx5KXT3L7h70FISFcxo40R/CMFmgu7rDwnL8vJVEsWpVf9N
OLEulMcVctAlFn405sf0CeDsqCWx2TPUgmXe+GyoWCGVgOf6VZQVg1NSthCOfqPJOVFET7BRHYLo
6NeA8n+koKU963twLlTgO5N2vOeXBV6Z1Gu1SDd2M4USwaNswixQRWwu5Ouxb8wTqvfYHctcZhlj
MyGaxsiAoiFPKTKd6TAgIfK8hrCi0BjbAH4jSHRDYMJoOFIf+RMi0DLVfVzknqilcb/23QCer1bq
XE2lggLxYkCCe988uJCIgnlGeDJrIHF2ovnJNQwAde5EisfinGk2avHY1Y3DdDVhud3gARlF/nSS
WR7A2KYEv4rqbBRrXghJ7TRhO8+9+mbQCY1KuB0WwE9ZbDqQCyoy6SXNiu7MQmVnX0Ln82Psnk8y
JPpobEAMqBvbWLRkyRmzU8R5FF1GzqoLAWVVqY4MnD98zkyH0LeDWLnUSIXf90BpCl1sONpbfm0F
IZC2W73UOqJsnmkiCmmVagVphAYkqi43OE/L1MHGiYmfrrsrGiOYvcC3dgeKbzEW9aQQWHgPQNs+
qtHKndmFxSuFZqI5PLvCVAAHgt2cBhts5ZvfpDyGeTZDbN/8C9VFR0NdLd4zIJWpx5peg4LmwmAC
M0mz+jAVbAnek6+FnxJp8f784aSBEIMfgkSlIuFWMHCCMGyRCh70mBQFan9o1GOiYTA0bb4/ybI2
UuGz/ODFRaAFR8ZiqdIDPHl9OW4bRaFL/83AEs4rrpRMHdaILu20F8RJfrePwJYF38ZgSINt97I7
d+220wADu7lf/kppWg1sFbz+N5zcvg/SQNYGLM92qqNDETL0HEixScKz9DIxpgSFiI6yD2CVO03z
cuP/MkHrMks8cXvA1GCFFr/N+Ijj6z4BvVtqb3mFVoYvST0TG9zDxo+4DDrLrGEtMhv13tNtDosk
aMzw92sv6p3sDSqwvZeIJE4eofYyij2bNQDnCUZ4C1EZCINWgpxH66dQH/7iwFAv4suouoGgp45b
1eUAewzWMYGloYQejCrtV0/22TrTdpVkmBuhEFsNI2RLc9vCxks81zKa+umnxQ4vXzItsLqxnkBA
nRgFTjzDpL+Msu+3DQ3KPR4Jhcb4MVZiFadyNnWOBsp/lbN5QPyAVcL0+10wEobCbUh+P1ZAqv8D
O1Oskq+ATKqNkBkB9VlpicWIey8QVFvHmeuCVAsH+nro1IUKOHQfF05yqhY776mogNNGkRzOmzpo
ivoG6LcMybzB5KbKguIXzvSq0VZgpnISQdOvLBoZsljTJ+h8s4LxqwQ0saV4RK5FPOt0zbcITZp3
KRvTwIdfvjYDiEcH1fClaNWHezQRCpnVoXJ/As8AtgNigki8WsuyYwg1xC6Zdqpa73NPDaCqyT0B
u9eZ3xXp6aHrIBrGC5jBwVg59h0pFdyuR0dekWxDUsuZ1kL875C1TKjw0di1Fwdw2gyRoCGVqHK9
qcgqHRg/7tmTZrxxX9phQ0H3dshWuJAziuMmqbEmh0LNLsj+vBYT7bSvrqaiBomez0PnawkW2vhE
iQtnLDXiZHFBxmyGIBeeZm/gCPkQ4ACWmWV6roArt3BEA8lPLwDIgFjnwflEA5FYQaVAehz5Lxb7
5WJJLIRa91al1A4I8U5BWbtUXbIS0Sssj7VMTWi+eY+ki3oQtzPnMVXyIJfbp/keKIDgAQ4Eb6VL
HhpEnC801NiQHKUh9/48lgDG4X1XE5A8O0ToTKVoVw0o1uC1vp25dWCShASKkcKzrHFhQCsa9I+q
rJpN4YTgnxhbN2VE/ANTsJdL+Ah1l6Upy9q380URDll3kvWz/MHiQ36XSgdihL0K5sbfpYB7OFBV
CbU1toEaGQEaM7QkYRWB8qwo4eQSUqpxVmRb4agSN864+EHDqKiD707FGGfvSHUecVVOeF8aw6QU
bRbkV9g9ZECYYquV/DZFTx0fVsXU6FWATBn9nwV8029dJBRTX8OuVoj6XZWN09ITObJGnUFnpwnB
rAtQJBqlFxWJMjp42Z2OBhkGf0MfxQq3TUKsaWqfGwyb5JSrXWkyqz1gXAoWx4F6R6KyOawZWwTH
sCS310MdyMm7ZZ8xVloUdYMp670VKwfVGxf9rHdc34txxdNCHRnHxS/ClRhCyb+PyDjPwDmKEUnY
NLxXyzv6hAAPYoXA+lp5CFKtYrsltBwvgffE9puw1u9MUyroVDW9/mMZkkkUhuKcAcYA/HmqcJCO
2qetLkGZk09DwgaAJ2SaMEpFubVEQbnDnlPYGj8ZQVeiG5UTKf6R7UCilsOD0HJ6eFXiP0mJqvB9
PKofRFgeDK+jWQ1+/WFI8zhDUe991nhZqZ6a9dmx/vQwB+52Kg/Go0LbQkCmwWFP7WX5l8iNjteE
sQU5LCpabnlSuz3PRx9HxPef3QnhWGXA85OiGcgUeYU1AtKh9LhIPjYnknp3yRUeyfdHoM1l8NE2
ajr2wTWaE2q5AzrShojguNl6Vc/RgzQEYpBTFscaPrdb8zkbWHQSIBmoaX41/xiyRHBawsUTo8it
iLqCSZZH78Qx3SuPOkldqepwTqai4h4UmQUwgOB0QbYoIbmHGtFCMgeIN29z7Qwqty+3uZ65+dvp
Y6fhcKatHN+OaZnLzQP13WN64SE5fUsFeiCGCZKtZ1NoJ+KUysegMKenwFY6BvL5/y5pcR+A4JlN
HnR3YQabX3uLxEggIe7ZGJVghI5dD6rKxIglaiq497igm8lmM+DKKJyTth4u2M8FiSnnjn+o/IWE
B6m97VmHXPYxHVpdP0zSnzJpqNhLktA3KITUlpNJGwqqsrAxxmKrngMs8iG8vl36fmUcS06HZSv9
7jCEmZxqAq+8o3/NDQgeqRhoAzPIri4nUvj3iRrQ5AsXqvSJ/veH2RJRefqf+1GC81jrk8bvH0Ul
Oup4mSwmGmjfcjqI2rhNlgttzRKe8ZDzjGn9jtxczAkrhxzY+ABhr0h5j6IsgSN6OHZCP20Eo3rb
gWut2aPmTa83cA9nP7/ybr5d3MCyl+kAur8zJ7vvxe/+ozLvOaDE2S2Hl110G8uwiE0kukM6FbW6
I/aKC4CLktySt6z/xRlEO3cB73XLPdBRC0zpEGJW7aznISLKN2I/BDnT6WvbA8HFtBJYRAeQhX/l
l29ppFsOJ5+lVE142GFmU+4vtVvp3dl1souukzQ9Ak6r39+udUfNYpY0Yv/k8wHTxz3MFEzq1Fhs
6EiCVeTR0CEf6hrsarNBut85RO9zeyHAGnRBBEQEExEcgGale3T+MNnsCTonRvcC1FAs7Hb+5DwG
QM89sKr5xV1lO8I/uOPVJUW6CWJpgY3iuC5Aq28uDAGe+DHlAuRRF7pNE3xA9js+NPPx9G1QQSrt
rIrQdDn/1SQABDlQzvIdXsu1eFMBJcjh40CIIYZdSqHfGZ8KwfWB7gIHPODmbvcUGXyRzaZgv1as
MTlFC4bFS7w1opor6KvKf1Q5CQuqvm9wp8C5xo6ZYRa1Ju/TTs1pMcKwY5Fc527OhfE5OwWTt7J4
dQM4dJZLHvPLeT+65ahlSynuj3kmKPrgpx9QQ7qf3763X1KKZO79Z4NEnrop3wxTNYmF1S7jDRrw
B9ltLOUFwo2r01MXGedvaRoTdpF/kMa+MnNRtYN5/NW+sGJ+oH37ufK/5lJxzGA9/gJebGo8dy25
rDTMmZfCqH/dGZFQh98hhO8czVXhYbU9tm07RBIEf4qqukaZKRcNnWQ0hvO2XFWUBIVOuXIN5mrX
IzCbfbgabFOkkbO6ArJKiJLzToYQLe6zI5JeFxyvGLeT6tQL484xEJRoIwXpnfmiiBPapUw6DuSi
A7nAD3D3XeSV7o3aZLXMW/Nk3yhJGFcBlUb9PkNXIsKeU8Uxef7HSBlu8YcoX263fQ/DA7VB6tXd
0ygYCDruUSlib2EUtJCU6Y8t8GUPoNa0aLGfLOrGWsXmXxdgYmxYCnlvXIx/oA/W9KZvvu0rhJ1s
C3Ace3mYOL/p7sztDcd9BRZNKrIOUcut2/QUwsBzhYMUEX/GhB+OTHMea9tNS3J6Ic/5AjmUKztW
MQGDohYlKgdijv9Hg7Xx9bnMxnv+96YI21Plw/dlzz7ejCWsG5FzoU3/6baZdpg7Dxzyyoq/UfCD
Q5CIblO/oSaPyBIfawbuFmdEKkg4iyNOjGNwuLFrHZHEPJ1gwr5NNNI7Xnrw9yypNK7oVJco/Xnp
Tzz9SVKD9gHCWvhyPRZevQECH3qLR9N++qgMeQj+LQk8Hwm2qhZYTqG09bONwj3ihnbNh7UsLBej
HcRDoUvJP6g7kYh04r5/CpQDnXEedXCkYKKHkEOsUw0kbEOLEix5zx1NoVpFUO3t7e4nUm2+eiPa
J6+gDNP9wMOdCQItq1D5EzCi48q3uXA/qo71GhxkX5yfw4/LMCtKXrmghSP9XrGq7H2nskpjF76e
y/Q7H+MCMhec/7z2x1uLWgfFggaR5l7k2OubGcKCBUMB8lENEdkmA1uReIJyzoLGvvktPNb0oI73
XwlOPGc2vPl+iutUwCP3iX0f38A5Ba3MrdQkifhf6z3JCr3CUPkSbH/4IB441LiaaBGAo14zg5cf
tzet2XWWTHZmNoDVFKQUWRh2D352c5JOufLlumIJ2FhbDwcxzh+0El2tJgLSzHO7hCwiLoqjF3JT
lVBfZH3gmSgFNWFCw0B1HV+LHmCbPlcCAON/TRUDTX11L2ygmjBQFt4k2GA9QCrmhU5Gtm/OU5Qh
DSIgktwqok6jiDdSUH2MxAJb1k6225jBI/mXO4DnAg2aDNoymqr7HQ6DKbapV9jdcEifAdqy0xzi
UjvSGRqujJzeK4dFfkFUMOhVyL/PzrtVNXPwP0z4S08ZkeMQ42f9QHNULoSDUR4vdA9CAWAyJs03
Dxvfu/Gts/mf4Sp+sestQmPKXsvyOD23+d3uayWoWeYGTW4j3D9EjGWiR8N7rxoXLjjqZfFq4eUA
FpEBqhsLx8P6oI/f25q6H4Bk4zP2eQxn5UDcnObG2hFXcZoT9hxUrO8N1N5sIwLAG8EHjA9Zudis
NjWI2MdJuTbQK1OgUWFAsQhgdybC+BD0ywMiH92BFu2ECUFlORuSCTpnrqfSEbzGfMJxYrY/YiUi
RMP2pWaJLMTzaaD2H452A5SjTkhzS7pDajBi8Du6wFcdIPTO5s6uipvm2ir3PW3x9iguJm7um16b
WViEwKxpsyL95jQUR9iD5TWdiR83YX9Qq/nvU8di7aByAOBWHkAgZL3+xN2n6lt9gAf4TlIqI7Lx
gsA1MjsSAb4Cj4GbJ4iir+PGcjv5eZN5CWnGOp2dbDn241WHaXcT/9JwZyVsUxe+gU7kxNejI69w
+K7BUmf6O5PvOZOYIvJQ8rb5uw9q26HkrX/jQht/DZVPjgcCZ+sT1N6hvABRpX/NU3Y45nAMD/fI
2bj+BwBIg/KLQ70bTDMXN1X4yxCAB3Ncnt5LNc+39FuiL/PJlVHKzRhQEn5xSFkfb6FCLmvdzmg8
548hwFPpODE31aKRm/3JytD4MSyfNwsZcHBE7ikZ58xCflyX0JbfQ6bfBumfUeDxiwezDU+ae3BC
Sab3gZgTYhuKJM20Bu3k1cmsS4Ke1hw+5so7MJ8hBSu7coHkcYQJL+wcEdw5bjSTfPrWhcEzdirr
HIADTapvO9hvG2wESNdIE1T+gd2jropvvcRFlcvLUO65FU2lto8c65jm8piWGQ3sL/unGd36MWz/
qTMGX2hAzUJOEWmSc3EQUBtnCetjp45r9z5KRTVByAspzEXVK86FKWm8eJ0/UAQ2lfn19dcm/0wt
LFpbRsbJ88jFGyZcri6qUk2SUE54ZPLCxVd3TBG2xoPu3osYE4/6Y3O7aFztBhmXLo6QthhhqUr3
YlApCXTzeFuAMk5lp0xwpl1BO8CGn7kHF5dKxSHYEBfPy6nnPBeW7qgY9UMYKTD/61zCjIf6WBY/
XlCnQoXy645PVcXSfWs9XGoevyVujOfkTZ0kPLKIZII1Zan+t9Ofzwl3b8Xks/donmkPkf2A1xyX
jeDNWMIN+l/tFKwr2uhP7T61dJBCHnfeaDw/oaj2M7jVHo46FRNfwGC8t+PUTyULdEt0ug/JbYDG
gZX12ztW3N48sXhuJ+YlDznm+GhAZYUCUsf+MnQlPxr7pA+24VLGvCU3onvSGihaUc5MTll89RCW
Cag6oNsjU157eBqs3flY+OcCbihJGej9uveW4cwt+pAWXh8BTzow9Zl9lQ7IOqlnwbRqAsYt+iye
ea9mi6kuRW+suJQvLGSXNl664SGiVPq3r8s7dGDLWy/8vcyAmDdPQQZhXA4+I5KzhJ3RM5Lgoznq
A1zuZd5kvy6AnRvdm6wyjt6I07++fp156f1M51r4AQg4jhjCAnh+Ih18FnTCVD0LCssy6uPjVLmG
XKLnqd1/jEZZhlKXSPNPygzDh1k3H3mhEbUuUsu44yHP56WH548X3ueE6tLzhxWh7XLmSCiGNcnM
4QdxseoRkCUhj1IG//YKSQtwaShM00hP9DXxksvu70I6rXZ4XI8B0gf2bpjcSJkcIhHYIy7N8Ai/
vojV85uUKdJI7wXCaVBDiURB6sEY275ZIlycZ81yQbcv4K4nMc85T5DgkF+NshyuuZSSbtCBgKAe
3I7Ch9s4xEfeM5rPO1nzaHUafLnmwZA3dmfOfQA7Blsl+yaihOLauveffAUh98epKqb0kcQ/90+M
cP6oOgyAyeOBNPJ9ikSm0wmpZufuoGf3atyS6ig1KZ3/D6wSgGKv0Ffr8xQw3kCyxUG6vBROvHYD
WH6Cxdk3FmDAK0fqYzjzlNd/A9RgOGzBous93FMdtO2TpAV1HhXSUZiL5R422LtWMn9RJngCJp+c
TEtlozsP2VhZ9d1YhIyaFakh1tUnkXGCl6An69boLa/5YYsQ22FghJPT6MGn8G4a+dBVuoIoJ6Xn
14pOldrYwRMxqQ2x6hcrL9Shg0E4Cn2TxQM2KyzWiCT1j5Sdiqdy5WbvXnBbrZ6RIetqO5oBL3H6
Slx19KkMW72uVpWzNJsXZDclxHQR19Yr/geR9T2DRsfFPY+OWXgdlPjbACjyHWrArnRhmLr2Gydh
tleH8nz38lxc2zTv6JuXkXK+VE+b9iU3kh9US4WoPQcUkR1THONx84FDboTHDMd2GIYGDya84+/L
OWVnDJE47IOoiTebzn9xn6mJgJ71OKWA+Bas41rbwCV3bZ6AGI9KGW+QnTxpggB1oLQVo5j/gUNc
e5WHuQ4Rg+mXDkOdf99DwpFCK6DX2GI2eIYWzVJBE14lNjB0FBjpNhbBfQLiw12iFe0pV0D/nrtm
gH2YslCbNEji8TeB/JZw/KEzglfe1WUb9j7f/Z9QANHggiq9kzpDfLtSzpei3SdsayUDULns9xeN
zqE4uveftghmyzVyehMt+Wi90BK3nKU2kw1G5bk8bAClmMotVx5WfvcqI62/ofwYaAj9vVAgX+88
K8PyXUmqLhU0DyaIU9IuQgwWWVk4Sh1zvb51bAztPTrnuJZYgMYz8u1p9/qkN+xMpJeeLdh9T/rd
lv8P1jWs5VInkjmKMhLaadDHIzZaG5N/PPjYSSwac8NiNNUAWEZE/CQiEQVjzEoS9hQeyzoiduXz
Q5Ot6SYcBV0oOCsiK6abSZen/+5WuD5pOwhx2Cq6mPfab0k+knTox6irg0QszIP8VnBOliA+IYA0
E0YUjq5nzp0TaEFlEaASJTpm5QEzW0z5wfbE+igbgG1N+f4A1kvnSIlC5n/QAmaP7BMy8Wc8YBSY
ALsFcNNZBq6SbVVjzU9JUp1LkgT4EhLL9YM6WYQCp0zt6GPMl6u/5h4O0cX0TMw+/Qy7hpnlnmEF
et9qyMl9ExB4RW3LN0KYuISMUHfhlEKE6UMXlJoEQmOWKjhdzdcggEsZy5/k65oItGamYvvtpGYr
DYA2qOGJW4azuwvVfUrMsqZqiIMIR+7XVsPAS4fk2yECwXGEaB17uXIezcpV2DlkNCvsVTg4OtMn
xX03ORtxt5CJZxRmNx5D17yvoew9ZwvOE2Iv+wYTCMQ81YEx+uE1lApAj6YYPkfGDC2ODG92EnWV
WsjXHwafaMtjlYcJa0rWjnETfZngxm+BwfcsD32ZxFz6PKX2PhlPPu0PZOe4n0J4hOvwV7sORBI7
3EDv8t5GHw+DGbM0teWZ0lBMWYigyYKD37er+KE6bkbRI3wd9zjkQImODL6k/W6LIcXu9l54D56L
IytsJixXGE1/HCrvjN/UqVFsjURaxszCRuoYbQRZwknbSg3MkSKLYNjMBAtnQMaTAfmiWy/awrs4
QrFAzGU0loPVvPfD6gC2TKNw4E542lqUiFXaDrm/Kfl+hECLWaTKo/CR+5s8kyQSAZKO8bxqclOh
ea9+KenOYOCIvTD1SutA14EFJ86eT9ojRqCD2hkJKccpNKgPTkmNEPwvg5tJ3X5XUwsMOlkVtV3T
cM/myNMJE6dcK3QG7P4S0XmHG66znHBo/kAmdQ2TEX62eepIg4gTBJxQvfnyh98UOQj47+6zSwOM
fxzjRwdTM03ChnhqE8pZYP3C9YY8wyyQ/FVCzigdEXxBzffxpeIhWJb5VzZIDtzbSN4/PRCisVw/
ZoELmJTWFMduItvZr6fk9F3NizPhWRJYEW1vayDnxXN5Q0RbmvA2N6v3aOdcK6E+mgGQUuIaTKqf
kzxE+yV/7cpJVfxXg9q7d3+cy+ShnabxalrWKHME9Ve0cX/ksLjzX1vLBueWW9jv3v2LOGwpMA1t
MrAPzfHBUmIjSQCZuPJMfJwY4E2tjUlzrk+ldnwBdL7bafLYMbEfIiUm86tZuUM1pU17XEWxMZQl
cThzH3v78fEKGwa2g1GG4opM8rypLGxmORJP8t1Qvu3pmFogJB0aQrhVGHNvI8sfLselhr+gRt1J
uUkBa67Uuavi6XtVb2wZx+OBTXuk6f6a5onEUsxuaesTK08++31l6wFTo8HRcTebSWxFk9pzlLVA
95Dc8lcJZKmDb28iK3oSnmtwRTg42ZuiB7EGBdEZa+qP27jpAsPaicMdeSUqcyNYsdXmPg/k9E9O
Ena3TCEvtMbyEGv92rRuAMrIHhQVSB+fOJnyrMDrWoB1EO1BKb/wtTx6tfmdHIoknBFMaP/yuCUE
pCAiwLBkaiSUyq/r4yuZE71a/YkAuz/HiUzXUo63GUDyfg7TC9US9pxdMQPUW9GMLoXsyGxmkYaH
9B19mozj/NNlsF7dmF2r5orjok2pSBDERTmvV9kQVjRsYm+SdOSsupSTsQnssP1om/qAoK6YWAhu
RhGsQxX1cNIPksWeYliAKfIEc18NMRjZtd04GftgU+mVAmIemGGOR0ENh/9ZuN5yJdMEpxU9vuO1
lXK5BzxvkZb4XTOTyRWv2B42k9fAY2Xz4Hj+ZswcGS8uEX6FijgobYZ6dar4Z6st6AdT/edpRuGO
iPLnfA1WOjt9LYSGF5uA5vdf7qkD1yP7C0K6f2zrho/VchRBo019L87jiC1YAk1tNBzcA1OO/KFq
ICWZcauG8lSd+eNlydDJzTYP+ySo/SPWRRiHHva6scDEG/N4OfuKZyGdlieMvi9QftAHv+S9Amne
8TdhRvu8KIkNZkfrdQu+hQYDTmxJtk0iUGqlb4l1O9W4drlH1vcm1aFOWHU07uHBwUOSfg0yoHp9
uOqvYqirV1HLqDc8DPpGEXvk3St8KrYGgl11JC27HHWkgALK0YOze8ohrSaGtv4nw6ZILLx3TTdn
zrVFi/STUl2G46wK6iIRjnGS/gA5W6rLjJbywh27E65Tb7TTV1GxoV8xU1kFWAve4Pan7zLADRu+
wWpUkeJvDHVu9LvqsUp1zirveIdgfWQu6EokOSDT2lwKLl7gt/qVUQ14zS7nqpqqbz31ZN3kyOKs
dEQ19aGTt+3BZucDSdwuI+3QPftGcy9yxv93sMelwrSbZOhQSerLctKiJfW/TRvI9cW1M/tVenvp
oR0fSb7gxdFJaHpkJSyKZD21Q8MydioMamS39ZxRb4wXXqYlFPeW1PCowTAIpzC3GCa85omc/ZSI
WxHEO2/i5kLStAZD7dknogvDwh3LCIpYZsKXbS16EiJ+sWXkolP6ENWT0q29ReO6ruU+yadMgISX
s6lC9q2Afwisxn6/3fyMhxzNYQu6ha+P4sFLYsWRO0RTfk7IUElWJve5mLrX0ld7GVgxgmfxq/zG
9b3jIcLGx6ORdpr86JTY4AYc2Uo1D4qJMSgJ8qgawoyCg/e08qBTrer720+vTg0SkrPAh07n8JBn
TnEBFP0IrIL4wa9oRfObROT1N57T+8f09qCqfjLb8KhlUC6kqx9YEh4hTboXOWrv/dGLio0SACPP
+wVVO6zwoqhGPQ59epk8sDOVJwsl+Hk5Qfqy7RWABQOyZynBKUmtm3M0/44l6AcGmEK2x60v7nnV
wcmIehaZ4qBXq3NchQpQ8r4LiVeh4vkOvYG3972sMTCaNc+D9zGPvddzUcob5PDldaltn7iZ25yi
qmSffbv4Ham2rmcKdrv5ZMvkz/cfIAf9/etqf+YfFyeANmBoBxKws5zxN4vG3ww/x7eT1txAA9iT
Hq7XP14WSKGjMcuNkg9+10BvAgAjd4eRYZltMf+9aIEzwAf2acEgaP8tNaSMHcjgVlkgiGA5htXD
+VfvlOZVrByo43zqPJpRdKK5WpOAupztZnhtmjIMbMPB3pCfrhelOnVeHqAgil0QIsqAEPa3ed/h
7eBE/uZDJ2nnG68o+HBITlZVME11H3lsENc6wsO/gGhMzHhDZ8ZJCHiqhQ64RBY+2ZtYZ3lspUF6
oCIFapS+UeN6Lv+Z8oZTaN7ICl5tC7EJKUsxezzyJZEGH5fwWEaZwc+KlQbyks3KSiQTnd1leYzY
EqjfCjFZDkRMZ6SYaNkmaXht0ltLH+i54zpIY7gaJrSm+GR4T6HVg2gmb57cK9f1N+P33tmtS1oA
xjxrJsZTTHSi6a0WTQ0n8jAjj9mbljdc/ehD1aOj0GPi7112xQ3fPf+rvu7o4SaaCdq84yQvkF7R
pOuN4+GfR5RGTzlvBsOFpkRilQ6EMFMFGsLmi9eGUaJyG/SUL3gHlWpjXildbJbMTc/PpWl4JZwb
VhCFoKXwBYQ2Lb2ws9JqWSpPopI5jFBpALxda3ks6yKWJEdF5mP0pQ4wF0up6GuAwXVwr82A4QG5
XscH4RTlZw6RcMnLoZqSBQl3VGrCbrtESqg0oz25ksYYroBZQecDRZgd0Mwa5BkSYOK0tz6GqqQF
bD9UndWGv6uVVyYgGAubeofvWprrLfuc7u0AYqFfOA6WlsspLD7EjAM7DubBhGgJIsVtPTUVhplR
yLoeq3LIR6HGRpkpm5XoKnrw7gwNrmHJWcRiT0TPNRy32ByT1uyVHb+56pYrxHUrKE7HuY3YANgm
qCFA4wTr+Cb2u725e6IaaOSHQkb44/xTfjrBdpjw5pdSG0EfVUXL9DkhxEZMxKyD1PxOnyed7HCk
AOIBShZgnSOX/Lo7w/b/uumVkhEJIbRiQy18+bQCU8Gzd4P58jx2gFnBmwZrHtmjVJXri1UOAOsp
fI9sk84aEsOv5tGCaE9Pk5kmBAVH8OBPAurWyBRt62Yz0FH5UnVPnrp3gI24frsdYVMzDw3Paixh
atP0RZRkWia4AI7cTK1VSqz0ums6WE89aXicsb92wMPZoRDUw4qiX3X23Ggi9c+Dq4uon0LPy3Xx
OG7XDJiEV3YtiJs3l45swKynpdK1OV2bD6wd4nkFPI/fs9Sy6DsVAgOJIfjd3h6V423UoizlnfC+
Ko0MSRSQxW+AodV7pSVMivF+n5LDznILW/K9jQPtpsRJ9W1u9jJabLbOjsWydnoCcMq6K51bOowu
QB52bgUFcm3eqU50Nu48PhNFTU+gYshEsOvy9G8MbwUIFuivDpjEJHjY3WM0jDTK5FOckb5NZMSJ
dLmg5CNTxPkEtmDkncZHVb3sjYcFG16gSt7KbBDz69xNDmOxXJPiIF4mBz7eqnrI7ibHhkg1nVBg
xwRHZsFOAo1en96lvDE+ISsElR3cf6Vmx5wJlSgLEuBOThyOsf2xBYQw8jP3wLEf5Q4MLMq5jcjg
5bs+MrfIX1kxQHt/yUW/PxUOMoyTZGxLM6pMWFrnbq52lktc46WJjPd4lnCFDYmdUZTcD9BYm4Hy
1+lwfebtm4vSDhkGdxEU99oKoLKmuJUF1UhLg0QBUhAUWNJK0iYBcfiy6+eZHbauTwNdt3fH7iVi
RiZNwnZNj1GNJZorPKLbDD9RxM8lQ3WbTtO5kQ5XvHonOM49m+HEYTfVi5f7lwL0zR8TjfQfPPZK
GATHKCUAxdsS3Q732XztZ5emOKQBwV/7kK/wU78qWTQlrvraPswMLQgzbqwCrr75kA4YfQX0jIHL
N1L56appRuSDlY+T0vV4l3lpHWtarZC4hweZUznlAlBdFD2x44Z/T/9oJpv4cTZxwpPEL6ryx4GM
AybkS/UxeyOscvDRz8cXMKRJoO9aC+nS1JiZNUVaHGn8F3sqB0moobzXChUehuuqCbGLIlBiazo5
fFMMXk0Unez8IP8Adk78BPQ6a4ub54lPcdtKrOnKF5hXpv5AgM0JW1ldCsfD9eqsiD4yNNUlTAvg
UD/O6/ae6hGsc7eiKC4c5Ikau7V8x5xZvFWFfyHoR/KHkf6qcbdHFhVFscTaLWrih5ygEx5LoIgb
t2aY4o8RPecTBB4p9NI9UGMnnFLHPBJkJT054146CUC2vhNVyhLN0hmt9serz91hDbIWjaE9FaKe
NdLvNkhfXpjalKa+Rzqb9D5g2xbwFYHz0FzBZrzBZJNUIQ8zuU6VpxxaNYwWly803a0DPpnQqFDC
39E+frOiNZDFiNClxNzXXOGrnd5hTNqQRL3SJSX2LFrZPzLGFA5U9ijtYr0g/AhPdRbYSJesdOu/
sJIu6Mqs2QEspLqj2IPY/FBlaIZkv/UAWARtHNY54llM0W/I72uRIsaLbH6Hls1Wb5u/ZuVlBYMR
lxpl4288bZsZ+9qPnGlmOcUqtXhNgsiUV/EpGqWVu5n1MkYBHYpRaTJLP2B10oe3X8SrL2QVRT1X
NJXd4qgyznb/e/gspryolpKs6u/U3KcDBx23f1Bkaj1HtQXbS9a0mOVEKcZ8nJTRt6VP7xst9elW
y3GWlVPJkmuql0lFgN76KvUP7lz18OftGBNz1AgpJZ8mmHI5kos/CexYL1a01t3PztMxtjeW9krh
E1rWy5/Xadl2uykuiQfznJsGg4M4wXcNWjDprhKEulIRK6kq3qMFEYflLnEtV5cH8orneUG0mD8s
FaCGInbYp2+RLlOUI4PYFI0zT1F07AUV4fRjHXTiLoLoWdA0VHcuNF+9JgMfMUEME32nFv9WL/4q
bn7oe/7wvDA2BigQEOuGMxYZCLcfU2D9ZRmD1xxEXXgjPktKiwcyD3x8thVPzboblT1eirVjj8O0
CiFTXteJhS8DKvAmqHpObbZVgCtbFR+VXbiOLBpCi4DErp4N66kPPHA0aDY8YQjRDrdItcf+u+KE
Q5sSdz8s2RSRwUxZ+Fyly0QEkP3CX3Ddj6hE2/wpj3TzWAlCK8rAC5r+pR3esEtsUsovY+kTg38B
jxPH7fjFWtnBFm7aHl7evQgxa5MzPEJFnv0jq0J8xJMKfOMH669KpZd3PS4WHPOzHOQ+69OHQ8lq
ID76jhBfVASTp4dZO0/V3eN6bqqN/86ypWFMP6IavtOfb1gNpuKRsnFTnvVDA8cqAD1omVw53UaC
tQvUQ1iGKFirxC3V93sij2wc5S889uo5l1blOVABoAP5jt8AFjDLtrR+AOVsIU+fFHuxqlGUhnJJ
nOBc6I8pxMAh1tQPJfWuUgBIhllf0spPwTD5I3BDrSw/UV+O1U6iwrDMGGaT3E3vYPfP4Covyc/b
X9r8mGrpZLSfqspEpWZhhfCOAQNLnUaPoSQER/n3wYpwR8JKBmLCViQ5qmhOF9x49xNcAbzaWQKL
GQ8X33FS2dawJ0Q25QCp+MA9LXmQc+sLaDnpv10PYa3uWIRnDeZvgEmwUiWn6iLsa7LOUT5+XOtN
8qbdklwZCVCjqEQX+kC7+jjLcywmpVzrhfhKSviY2dVaMlJ6Cf8AEhgpBACJAmCmbjVeNbrTI5/s
1SWeEMX1orhyO6jOhpBFWd/hDN3XAp6mWoOiPhF1EU3CMaFFVZWm5fy8BJvZ/DcDlIaUks3KN+TQ
5TQWt48tHFGh15XBuoXNPoHvFPjtiH0qvtSBvCS5nH+nL4afkB6Psu9euOmsnCAJhIUIeOeXQDcX
Y0trPZDmwHl1qQC8y16N0Zvte4zqVQr6LHgdMQzeC+J40Wm22ogzhITmZ6ozC5u9RCugbOYDYM90
qkhCxKKdo3UyzjhO1QDYZvzlXMh3eq2CDUAvYfrcA2fAHPjYb666cJ63aAGx++aQfhSytfuS/WoA
hbo2aM7CS3sANilCMBfP/EF/i5KIIlZdCwHmGI+b/ZYOyK9W6WEI6SF09qIDVAN5KxWvm6aq1lUY
d8R8Ryp9itgydfIcVog1PhukbnxkHpql7vAoxzo3P06/rRlqbUkUT4tWn0vbFhhwUhzyv53mKgkj
lUbhZK3D3NAk64xprEzcjYSTr+8LsLM7MVW6o/E7iBWgA5q6TD15qTiFUoC7OAuzw4rL9VwVwbc3
2hRgTO1RmfvtVMIkzq8rdkJ/Qi94roccXp2680Y32yR2ukone4D8IuBI0ao41pU4qpGwD4DDihDi
IK+OTos55Z2muq5AzQRX9V5HWx+CANu2U/5qxm2ADdI8lIYZXrpwvk/7FJ7CURwJrwkCbwDpO5vS
/0Iyx4GSYRW8kICTs4NdAPwoW9FNPEDuwfuTHSSdxzLTxteEKf+Drh0LqMXKnxGCzrfZoOP3mBMf
y4poh77ebBhKvP5bAgW9a0WS/eBBpkfYPwNxYQwgb50KHKqgR1BnksuhnkX52LoIELXXatA+F4Lt
bx8COm79Oj2vwzhdWSBY+nMy49hwpuqn8bXrVOfVD2YgYwNClLEDm4kULFE2Ubpb75WDifbpZWru
pThDZKvMGA3gL6/Al4/1d9zYlCB1iNf80l0z8vmwXN0udmGPkTl0NigstDclsNUyS3Gh3m4gO5fB
nKdhbo3mIcQ2OoureMKekaVWHPngGqSK4pIEx04UVVsN7BVcE2kciT4SzlIHDU7DjUaqX7n2Ilgl
Xnhdeyp5wgkgzbHWQA+zeKrVM16NkfVBDNIAJa+eQuHrpi9E5VTgqdMbQBMokUCetIKLGhdwMznq
MQMeAjstymgCgNIAKFvKIVE4uNjKIZmCoYFtTiv8TtqWPxxWbHq5RUKaKWmpuU/9Ykyf0s2Kzwcc
tPBHx9sN+eJzq+CBDV0Q5ESXk62XnwivQjPfRuUdBAxGZmQWhwH+LnfArFMB8h/JnEzA0A419916
2BCKAzCIBBsobmBUhsoOjKm1zUcdTLfNCngERLvxHI7yZDwlKHO3NWUjpVMBI8E0i1NxTMYztgdn
W27fSlcX4SLIVFNnMatPHud0GdfrkgjF3BK2CfVjEaTlOog4+QxbifRjyYsXrIjDVDlQD0oSafJP
4Tx3q1T40VWI/bErISFKQhzSnM02+kufz4AT6AlMGHtK1wYDjWHFZZIAjAnZ72HPxewqygWkIxum
OzhRrO44HoiDwi0+EN/FTZ6n+GY8gFYEvWYM88sh3JtP7QMctyOPY9KF8oC/tDNBX0eFFW23neYm
LCEGMjl8Gbz+FM9aez8ksSeFyaMs0IOTuRkUaEQsr7NZL4c8hxImr0epj8HDdz4WSU5Po7b/DRBb
AmhATURW6fVNgGuzZG4X7I13TAG3C7I7agVgsCuqxebjoVtU56F+8gdQSXs/AAG/APQAOJFPTlwL
CqLUktX9AuJ3oXz1OUIQMbOYgGG5D42QHHglD6EBm36ii2VVT2hGLlopUYpcTVYOMxmR1zA/T9Av
eGMTyrq/SBzT2Ojs+prn5fuMeXYQOO9z4uEKaNckyrEGKB4802vv7xyPWZNRwB5fJydsM9tj2GS8
0f+23SJtxLEY/6i2QEZKj7RO7vKK/c2aT6BS5iiYTtphcWVou4+ra0D7InW30PuPkHzEhLJOQRfH
MlfXGOSN9KsMrPT7Hwgv7+N1FiY0mcVZpWWD+0EwRoH3sAPAs79+cQDKzdQcckGphJkgAkqotdh6
zKYmY/efUl2Z8t+XJ6sLdTmW2smRy3f6ffxemhVL+binC8NZTvSLJeVXoL1gKjDEcC+pfuyYL3yb
eKWu/FZjRk1DoWHQ6AMxjhTD7ZnmgG5fHV1mxpc66VUN1QvFvw2D6Uatu5bj/3LWWPOhYuIJO57U
KVchvpsU0BdMrXPXgkWCaN6dpPTMTFoP2157DYePSl+1n0JjSKhx3UJ45fbOgRg1YzplLbgJi+Yc
ILl36traVHs9gITFlRq+gstb98YYC60mKBXTHhOJ645gMV6AaR2Q5L+JpI/F9q/AftkDKjr0+zwR
ImEm6INMAYTWIY/nlRcaxbvC9UjuDfKvNkZ1anyTo4jRVfCU+As39+NpXkvNKregxW2JSqeSw/Ss
kNjs6uAgRDETZDwPW86S00A5rt5VCUZErRpc3ci73jOVJqn+xiCriCQxluhejv8K7rURUA40tWJ2
rr75USLGMREij4vWaLIrPo8BULp+xTvlt0o+7WjoKkjxxWH4x5vPWtpCT+xVDp8FJqV9npP5hOUN
wuJHgYDQf24nFadmP+aO0U/i7qsjTuymQfG9wC2tLdOPdd8FiR1duJgjlFzOCEabdaJ4ODLpoXCJ
4KmcdYEwz7IUzDD6pP4ogMhPa6grVQli81m9yjkMaubpWtuh3j8jrJYWNM/Tt5KiyZSNoajLB81S
2Cd1Jv2Ja0rkC41fjYaPacChjkZyqT3e1kUe2NeQ21cQ+wtpsGJI4qnc4cbuYi0jHUCpHn5e+po7
za+OyL01ztz5Ru14BKcqi5xhG5s63h5Y/qDoSTTlwiRahyQ53YDYXvRjrqFj/gjHJmyfp0iRM5ak
r4SpPkuSVkzet8Bx2U6gYM4yNtMdD3uwIWmmF20Vuj6I5NFZCbSmFJnWF6iVgGmOlygdbYz1kRRQ
VT1gNFIEBN/2Z7K13ypBAsvDtgOwA+dqXZRZ7PIRGobacjmSyQyf6ik0DFnd+SVQOwwTn8/K1bp5
i2zTNfgE7R4axW601eRqJzH78m3wnGapvUtvpoABEeBIM5kjr2GfRhmtPKAkR38Op8/k9dn+MuSw
LyGoIO9tne3UojS9K2CwYfJxZJ08/Yxq2Xn1hhCJ5fNtnEaRhoEW13FiJGZ/PmRJm6yqj3KC6ps6
KJmKJEq6Lh0QENbc8VyJYrjFVKMiduKLlkO3rq6qw0yrCQCrll1bgN95PsAtH2hfnZWR3lqk+4U4
vqpx05POI8pU3oOI/nEgI5RwW/sBu0TNycMCsmDj3G6lTHqWIiypUhOV6iH2PGy18R+FWtt5HNgI
j7dvXsHAYDc5jShRmbGyASHScgFRhlB86vbmsGvi42gUWT8Picip5ZODxbwASPt8pbdiK9XXc6Ea
F+RZm47F1PjhoDY1C9PH56okc0HRgZyVSLB9bKePAdWkqPxpT+we6fieTUHCPWPDua4akfBOutIm
2xoPuFLujcmJ7Udbm5LffvCId/yHvfU2SRcIyV+/eNQVeslSm9lwq5AkhP4wWqAYSiBenKabv7Ln
kBLOsbnfXQpP7ZAcZPFVjQtRLFF+vxYMCa1ICqN+CSHlHSBwl13K3J7Vk13ieQiw5m1IjSUxFu11
9NhUo1AHV0BnRoJqB6tIvPutbWJXpDihI4o4kSGQfULLbLyfMFJ9lh6/PRsUnTwHj9O6rWnl5rZw
BnEQAfZOA7SdZ00dRaF2Y+g6kUo2LTIB2xl/4D4en4+murLtqozGNbDHfyKY6fco5Pu4FV1odqC9
DcRTex38Dzl5YTZW7WRuszmG7UBa8tgd0S/TBdi9lE8Lmbv8/r5JPzFcPCQPQOG6Z5y8tl/DKuvG
KVUrqWmNeagC0coUnTAbMaAIrS8RD3fDPoATPCHZJdG0FJFyrALhcqfuarS7F647p32AGktKi0Ql
zkM3r7idUKKFAWoxSayjEZ50OPodfsLIY1GkYjXv8TcNr3CkwsdyrsqOvY1ciTGBanf08aN5DSGS
7zrktnlm+lzrue2YTrNSHpZ6YzquRC92qWqRUO83t86Ye7sJaWSmof03m5Jl3LFToKF4dTlMR7gQ
QsDk4xQmAFwsBYY0ZT4mJnsXX4YSnXFcfHajXGahVYxLeCxZySz+MGHW6DZkrXcOmlMQw/enYdij
eBjaGij9KwyhI34aBmevyYEOZ8bEkcZiIX8uHGU1g5VYi3WSUxfTV5TM8k30wzZRuK4ytPLhKqBT
IOuq1q7crLOWb6uKvFy7WQHeqH1x8cm7aOqGoHKm8MyJOQd4nmuOuvnABLdfl+nzK2tdxbCpHv26
173aNz2dJRh5KsoqxhpZC1d/SYe+rce8UPOf30t7qIM01eApsEanh9dWxnaMMjDmuLkOZSOFXtc4
uvixAWVgGXY+f7+q4QQgUlPT+A1vqzqgFu6mWCMW64feCz57mEvO/qYBdSribE996Mc5vqkh7ckg
K5pyuDpUC0VStyOVEh76CMIremPSiy2OzJI7rrL79DXoTEoUNtYhWPLUtnRIiBTJrvX8K5fMDtRG
K2bebc6lMdhwW9oHxJ/Y2VOeFLqOntQCt/9WlFC2PXe+RGFaD+LakXHJTlsDoyAZ89vQyDhg8+ab
AHsUwjXvzLky7x3IEAH66RIhh3soAZEi17yvhiu/+S4x6ds4rSzfe39Cat8nurawoWYDQcXxm1py
jNHr8M4I0W6jC9CE8ueZB9i2hPhpX4JJ5uKI2Nzrr+ODSOHlntJr9Qjzlah2AoN+VWNnombjZCdj
VLp4XwKOCd8PKHsCXOQlCU1T4dAluUCQurT/o/wAzlTCPEKjncpdygaCXDz5YMQY32ti3itV9UBo
wyiDCwpO4ZX6krPnOyAB1AAcXbrMri81W2do1gtmhsI/lJVuUx6xtkrl8bWqOmN4lQUXa2mt0Ngx
VYDYGfG1RiXBwKB/CgGOm9lV3Y5YBB/e4MVuNBQRBhCN3ptH6nfL/ELxe7DNYEeTmRdydDObYjz7
33UXzoq2bhau0QFlOhpVk80vuNMXCSw71IKwa2d6uU0l4dHNqDwAn3xQ8o9yFWs6Sr1adzEBCrab
NEYaUcJRLFttzE7cYGpeAC+O1ooaZCWruFnwyAQJW24MUGt5NNAdfts/vQm4Ci59KoqiL4hLGd8x
BHYfQQVyCuM+uUW+m21VzUOsWum15iE7bwbt3TmIs3aSh0wTM6xQfJ7g68E1V4yXpglFGitqCemb
V6VFhmSvVItM010YnU+gaXVisXLC+OBlnkcehpEKnzW7e+LFhOziIHVhOp2xxT9KN5wBxvEiM7c4
ZHFmf/845/WHa6beBtfJCqFZUGt5Mr+OyStpQFQ9Q8UcviGTluZYGfdFSFsUuxI6etvbiBMUK4D0
j5587xJ3Vr//jhjyqY1sCuJq9uRQlaZst5fGPRvqv3jFiNzxbvhN7w8HvaMBAinMrV5gQ2aZhe0k
4pxaY4r/0lHnOoBjtneQ+l/zd9YWfs4ckh3PDfYYxHsx0RgyTQKJsDUix1jWcoyDdGwdknSTKXq/
+L0Dih36iHc8W4jklWeFw4WdhOIvPTjGPe1ZUwBmRYApmzA930dYQmg4INrtenCHpk9yGN+Efo2a
Rem/hElhUJQUDpIsm0Xjs4OWgb2oJq6vLq4U8d4dHHJ0eOQ/hUs6WTwDOTiIb5e2BPU6u95kFN+C
JTSJRfxUXxNB9wMtt5lFBSV0dpc7tfYjrwSS5d1QPIToLBHhuprW63r0j7x6wqOoZL/oOK9Bx1Ys
410cZo/VUAHvWRf8aMTPOKGrmSI5YenOGU5HkLeOJrYYSGKNMmoWgYmMN/u6UM/hTn0po2Uq29TZ
it3dkktWbOpvRiTENgrribodQuugrUeiF1uAB2X2tINlk0YETiSZEW1/2GWjb69xQ/wMZHm3cGBg
iMECN1Z1YVpZ6o8FUVrP3evxJmSs9FjcAU0qFeokgMLGfvETL20c3neAd/GVZy0scwV2Y9z91xNl
HtxuNi3PdA78gwrbfCRNCPw3MYxaxFbKRb9JarEcWj+X7DkG3JY9qP+N3UYM/3KBnQg5A2U64Ky8
y5SVUR5LRgdJt0mtOG/p/HLLymlggWB6jB7elf6GoeFKhyhEzpHJtWhoHdmpz48Kwy1zDjIBkNht
4Mn8422z6JCdm9ERbGwvY5I/cRuNXl3MlYbR6ipZrB9hqParH0hUKaSIg9hSbolvDPcl+XC6XRV/
nsdCLI3E4Ys8tAK5CA2zWne3w5F19aQKrkp7SlN3MniaIXVioOMlhJaW2Hpm0/2PdVmi9FUu44Jn
qZxOYUTPBsBd0CVj/3s38Wh1gTa1HrjtHka32j89iSSLp8WzNEiATQ18oIy4Ev1dV8Dco/FGyt1J
Cjdle4qo23D8n1mCKzeZpc4lNJ49l9l3SvDO1iDrGMI8ChB9aSetZpo+ITmNJoeGmbb31pvs1KjP
HF9409KvPZaiW2KCMk3gcOibjP2GnXDf2VFbnOMPoB05WockRrWNdMsuMZ+bTvmv6vz5IwHjwFce
47gbJyDR5pjvtBBoTfa7goJsA+kNK/WOURp6oYJKdCoSItd3Bf5uPTfNXWxgHV9MQiiM+05qiaMS
T7Vsxxny1VVnfzn4Q8r93qeSK6/v4Q1SD/db/6e1JkZIs+wf3O2qnRPQnEGsl4kjk/NR+cjALW66
loCdRtigmC3E20sB2tBrUIkdd/O/h0zT2QzJTDcRrCXRMW3nd9C3utZah5Pz3HATrzIzKA0eZiYh
VHbhjyu/3hw3CkjXBMv2jTx2Bt+MUOq71J06tq2GIG3gp07TpER3J5pTWSo++W7cERSz9KS/x/m3
ohRSioO8t4QL31sNn36W4JgLPYgPUb4mR8zDMEM8ghFJwrjtlcfPp0Bqmo78mcLhIthHpCsHIMdq
4BmJkBfEGzKev1OV/UcgqAEBIUOmYKQxhm1U/DyKKZay+S74YB9PKbhhnhcp+716v8y2UfZ5G1wF
rLerpclWgtsaHQ1oUEdheGhXny2PAtJK8MARq7tAfl9jLLASzEp2E7+Rw1NQBm4Waf0N/YmuAtl6
Ncpe0tbPF7ITZ8jFwx6f0RAEnbBE59gX/RIuCkP4iLce/DEnLypmd9Bq4igqD0/pP1Ds6DXQSfRP
mcfayw6r/Mo/j1jieJ20+0wWij2YXl1leWSXnjDAqzReCDEdQI16/p/eRSZLSwrR/kK84FoTCXoa
6QorKCODioOz0SrPvQK/QsuOuNg/cNSOSMW0HwxxuzuHbGoTlgZZiwiaGBGORfl8fFJu2JpfIEC7
0MQ1q4+6QkPi+o5R5epK0ugnGUejxoyuFNpMW5vMCo9QsvtdescccL4Vpwp5JjXTSMGO0iTFBiT9
46nY+2I/3UXhGsY2jDJjC3ZveiybVo4xE8b49hsA5c4pBfIUVdtfrTSQbvlCvn1BKZEglmvcjEGR
us8sghhNiHfHLWG7TPRY45k3ln3FGywUe+5w5yHi2wfmku7vvGyOayXVxtf50So0N3lg6DVHIzy4
I/gpgCq6t/K2aR8mCl5LM65pZXqlqP9aiqwcQvesXK4wMSb+yE2ihcUHSt3RstVUuYXx9CAfWb2E
mPz/YDA/DAezjw1fJ8L0bfr+rrXA71QHajxQwq9qol8tMNANo1N/piS6rs7khfD7rBFmFzEUizxW
dFNN3od4gdrDpThcJYW+D7qvNaiN5+FAybdFbd7Hm54L0dHz6uTtEz1Tua0rHg5sFI8R7figzF30
MRiF01lGHriTc70qqi+7lk0dxgnP2eFnChKR43WDkHLHkxsHpAuGqQbt4T2Jyf00ULajang7aH9X
UpmmlcIWwqgf+uVeWp7XUvYJlKMQPLP091HKcDk/ExkSBdOC91taxeN0CPpA7l939x0rAmEcgToz
ykFkvedwg87ATaFupizajyJ7WqwRApwk2kXWjGqbcWfLiJ67jApYUD8JyBwp6zsFEAlhRnRxBEnE
l49ZiVBMWeKgVbLRthMVN7aUwPGODNv/lH6DMDgkyJdtJB6FjXr30yTQM5sVc1oZTMTL0qmXY7Mv
GLktmaBCTmkJH4TBX1xbWh4Cj+hFbzF+BFOlOKscjliHpMZ3IadAW/c1Opqw0AfskaVmp6OXl2eL
kloDe682HJF4FOCGVEvZseuskdl8JsN9oU3TR7/phuN10hr+RLug/xOaQDPJ6c0jv2aGYTAwpH0i
EqO9QZ6chMVcaFtfyF4yuR3cc4w4l97WFE+yqud92GDYqpVAYcYuNRua16NFshm3nxNFCzfoIfGP
Z00CXvLXDUak2S+N/tSjvE/Uupy6qqt8XQBXmthr1cHFLSrhn/7BBkXhFxHuSdC07CHmW3/pEoTs
ZDFmrL0WBf+Mk3d87dY6iEWXVVKWYPYxoCfM5KWQSF2f8PWcLxpko7n9dnsGpKTYmCV9ZR1rHkZU
3ZG2OMZGPn5qId9pgt1B1aOK3txujZRpK97mKxjPg0vJArx+31S5FRlctJrXQwG8dBQoRBNnpeDc
EI1gxOrZaLO3v/XxRBFpSj/vSSy/yXb3FMNQ4KXlcQRiCJGBKroCxYpD+TSy5laoYW82nzVx2/ge
CITVPbEnWFw/B6tLr7DekfxQOktWlICdQc4J4PvSRcT4+YAh4J5BEx9FvKegLQ4LllW3qaY/mUFz
gzoLGinQRmF3KQfBe3gN0vVfW6H8jykO16jYuNycEq3uKqZE9ImiNxZV93C3E+e12ciSX0g/YqGW
xLcyfCdy412KIAC9yYP4gP+dWqZb+i2rOTk5hFirLkC4GuxaJQ+XosT9Pf7mTsJuQbHXOFx+M5zX
NGf2XPZLlpACxzgFTIw5WG/9XtKy+WmZUAIzzG5y0sxRRU8cSATV/C4XSbGzfpjrOHGk4DHQKEr8
NidyaFUmDiIr0LP+ByXXedYRGkHxhDlIvcyfmTqOlpRwhiEXub6xq+K1UCJ3SjTkiNqE/mDQ97va
8ulSaqwkYtulyWVBnIomLSjqpqsHuGWCIPd/NQEIO1GbRrrlo+HFTihpKlI7qungZU8u3IyzVD8B
JhkbRCgkjHUiosNFawUggouGmTNj3NY3dQW0F07K0aldQILTb6W27cxaRRBod9+S+iT5cfnk7OG2
op5wkCWbwtWeLkFRzg6y69c8kfKxAIFMv6hMGuYpX1+xkiDeABxcJSc1Qdf+rfOKFx8FfADmyKSZ
SBiotIIvEbIpR3KYkuvaTHHli6muGZyaTRu8ZmwgrjGjPOliqFrqTTTYSZTyu3Q+MGfooAFRy4pS
LjkqR+v4mLgmmszSTmZ/R/WLU93m9WHy94XCCZ3Y92XSe4IDT23TKhOuAvb82p7aGgHCnGcOl2rv
SPgLhB/ziKW04yTC13NyR2rnq2jQNepfMoRLtPNcZe3mPQMW2wTQleo1iF55Eq09NCjttlfuMe2Z
nyuniG1EMy5Wy7mP6Uk9pjpI8YWqPiSApoFs5smHNGWrxDIqRL5oRrSGcaXNTEjwhGo959msnAVp
MFQNjXKjTBMIVRGSYco333Lxa+Nc8EdRQQ6p1+tE8lVypc/b5YXjpPJLOH+sDx2HPKGR56IAa5yP
QqbV6povLRL8kHweWuOtsd9j22wWY7iTRvgylQStaS/+favU/TDdxFbk8GUUJFKoql9xnUzBs39E
thTCSBsOUIwUaWquIOekOZ8uyTi4+isI3kPxTWpbMTmDV1X3e2oS4IQco2yPWo5lQ9bA9HJRnXZQ
j8CBJUmEcLsxIEjIoi6uDoAp3ZApSMMbREpttfRRO1AylL3f95A8Zgb8R0AbZ7AuwkjKwRgp2Ww4
/+ABRrp9CZQaqM5G0vioK/c4/j2lL1wsjBieWyh8eEVp49VPqkswDIM6fBXNHgwqLFxmlgLcYoRP
JpUfoskiBFqwOg/LlZ+2yQrk4tnXvXGt/XlD1yPudSfAJ5Fbc8hRZAj2PnVW3elhQlc84y2AalfO
m45bzDWcdfxtsQDIO1drXKQSxidD8ZN8YTNB45g5mFWIXvjc3ckBkH0Lca/Vn/U46qT/Zdg8z3fF
IzdBrWbZgp4z8K7VGC1JbrkWpMPwIRZl7+4/Pb3Ft9ccegM+anJ8LUsimI23zCm++jwgL+0qIc1x
Kggbl8yLk6Ka7GEUxzhrTKVWBbGtyEiWDc7EVpqLrf5oLQ0NLdJu4Id/iHlYZifPOxevrJdjCrit
8G+kJvDWLH67a+yI6QasYaVcmSiadFAnip/UpPmGJL7NfHT3lx7XoF4a9efgtZzwVi8lOVYhjQxm
UmshGthqPs6PvoLeaG33TWamuSuRWu7dnMQ8AHM++1X3riTy1B72C+z4fobouhehWsBfeHbmfbVi
l9cnMk2oa3+j+DYPaH4+0OCbDE7R3KHlKY4yMuZgNeUDR4ekiFdxbKEKIDSz8byrdkcbSZyHyE/M
Pylj7SpxLl2ywoIRUsw5vRBS5t0Hvq+kD/NYWdYYkeduVqdUoss/pc75d2e+kCyAUhi2U2rLjeh0
qjVfU+pUziThr2gpsaTUKGQAA7JpjZ1bxY78C++pjoVcfMWCTFx57y1uVs4f4ibmZTzp+wLkNsvS
anFEy6wZ8z8yvPr3Fgy5See3Ogv7U1ijfU+rr4EfvEr8tTBmnhgja/9bGMJxj662aSGU5Xrnwpgi
DLfTIXDH4U7nbGYWGoMaXf/3q6VO/FASu/ytP1SZ3v+PeILIoxIIuiw1cuHePHu2aGjHXHMgSMac
uCv68HWNe8ed+72gUgNrBdXOdOn7r+FDMsBYh7zUEtUgmwdFe48AavvAWuXSc6TRD1/LBdJ/DaQY
1WdYYCpo2F/u7PYgQxqz6bgHMo9P0CHvLLRDkcikJG6hZFAJsfklh62XN/VQSpNzmYyBTO0BWCI/
xkHbkuatMU27EN9u+rwbPTMm+0DkVg2lyIvot0EzuzlrIr55Nzj6gwyt5TERipA7NahCw8GH6KW1
wwgJ1a74jw9z7hxFiSJrBImFOHdL+Iy9Q2+DN4ayCrNOej1018+Gu7xPa8cf4RWF6EyZdk3ceTS+
PWwv93bHR2xlA07Bl4EipfL1uiL9EWGexArM5PF6sfZRaQTMbG4FURowaWmPHuO5yS5eQXi9d7kr
uAjAfJGV2ln/YURf0+7147tHpnGq+df0NzdOf63T1DzHLZ54vebFpYc6IGixwRIR+So6wm82llpB
YfnOCq22LmwTq9P2OJXA0STSbkZORIhVfO9PYTxEJql6dQyyv0avTMc+PiJayGeyiPYK+5CxpWz3
eQmVWE9ziRdUFZ5nZlzzrXt+HYBsSpefFqLIyTabvAsqdMQ5+KpFMmYXI0M9W5sKScQwFU9cU7m0
LuJoq+/JyHg/gVsQS1hsDWIsbyKJMD2wECPvSuzgBxuiWbtntN1K/Tvn/eWYCPRmiMfBXMWX8QJi
/xE2Ql/ktrfnp9bKkfS0VgE9ABESs2KSqpcVBzDnsuq3rQUm5ynyCcA9HGyqcSigj1H0b7ZsfeWd
OeD82G7OIalFKAMZV9STdO3ArV6jJwp2k/KhD4wcTPlfRfss89w/zegK2VhKiXnZ6wJ7DBjAmdZx
I5stUEKH2MeD5LLZshXiHTlsjrG8S5G7JUxzyOdrHSXkbjGARAoKVw4i2VXrpg9/Q/kErVt8DCFj
1q10KeVDP1M0015uw3njSHQwa6elTtL2pU3tCtY3hM3PJAMZpGqaAoVhQ3FEZG5is6D6yqGv3YsX
OUQke/T9MukEZk+SPPs87L76Ff2UUA5Ua9aNLUSw/xVY3zNFu2mIRT67xVvjxaIl7G6NpTLAQ6jN
yfOz/2y7v0x0REc9sCk4sc3emQJQn595+kvcl3CZxaRpRPTC9cT2xrxDK5x6nF69th+xGtoN+sBz
4Yp/EsLyrK7tJWW8u5NhjXOhkdCycl07wRDDJt7m0ihXWkV9kb696zzXrJO/PadBAMDu5A4YGyO+
p9i87nT8m3VhX5DisakLoD0Nn6LlnSeneNDJMsuK7Dccs+/n25VrclL96aQ+2q/fMi8laucbTpc1
81G1xTWbNVyN/m7BjYDzV8W91JtJ/xr3Dt5bpy5X5gtnHSPeid3eCpFolOT3x98c/gePTUMx6YfG
dFnL1A9eGU6TKXFnOaKhsPLvP4SOoLatHvDcc5mfUdyDi57MrizaJlrgKwXR1P9E+YbTHGw8QG6I
zfXb3OX0w4HAAPEOxWIYmczeA0TwJ7JVYWzTSgrvukbRSOhLSiUOSIZjxH8DTyIDXU/oXxIfJLf6
Bv0ksJNu67Rjk1LHyRB0hljbGVzASF9DDp6eyPm+xqhhaIbjnu7LGUttkMiK69ORXrEVUfHWxaWR
MnebGNDNIIGRJNqD9nkLYLUPXdRf8/6Y1psvhCmoX1/R2WMyQqq9CxiCHJUFNuxX4dgzqVozjV1A
d4zNSG3Go1kPj769ibgXw1PPZX2gfCpupypCrTpizdMd0rnGrnzIekOQrkyYQHyded0A/QbdtJY/
S6DNfgaeVipc9ShGElSyDoQx/dTvKA1nKqAjxQ3wCLJOxGrAhEDHjquOR4VFpt3pCXd56lJLZru6
pUC+C4Ki+SC43km8p3/hqvd02fPBtbkvpE9qVnA1/EdP2bY/JQQVx/EQ7XAkzER7pr7fxRf9xQzp
ntSFBEP5vCpEIK53k2p4UT1YZ40V/s8Vs8+bpsZP+KH0aqk+3BJQAaz1DShh3K4vFQsLR5zz5AX3
lGR4KLT9IBgq+dbq6ZaTEjVMh5PHqTKQRg3n33gweCyT9L/VNxHg9lOIvpP9gqA9JemzHfcoe66s
N05YMMAdqNk9mS1nNIk/IawDMfNoNrIofhWxNKGrSQkLhAF/kKqFgI2uLGzTTqegJkaYEdP3p2Tf
7Xpqnn8PXwZlWEMTXrGVHqugPNMV939P1JP2N4fljjEa7IFRzS0Tt+juK7sr/A9ndPF5DCBoc9im
KVmxQ+Dy0aIxUPQiP5niXusJRMM4teAjK+1rbb5djsITAUpYPLS+rtMFa9XGWiS8xYfH3XGir4C6
tcKTg3T/AX/6IdeBdXqaGCBZ31i64hPukKWVztDK6Z8z0YA1XW2EXm3FU4SnEmNQ14I0hSi+V/YB
rmfLip5aV9zzE8FGogNNfEnO6y4QKDjcfs1INjfSR6IeaF6cgxnsdIcJlA+P/x4wGYwicqjZV26f
7sO43rZzCGKc9mpcyUj4io8Ej5UTxoGWoicntMbFvbXGMbmHQUFJb1O5C6es8MaJckwu79xbKYQu
XfhVOtXgLlyMfmDUCIYG7uNlo7U5Y2FUo7X6dYcn4hUa28QiC4pNlvJfZkz8VnhuqedsT8fNDa40
KqwNwYtQD9kvpOOm2Huqn8ANTBfh9nsU4bxfDwuJSwMEvkCMczMeeG2IcYjW9LEfmrmoQO3TddZ/
TqQh8daitJdJ6R74wHQKdvjQyglxFKO0oMoEFl98/FGGzsbLDnt5FavuD9KdvSiYFAxF5MVpnNsu
0+M2ZdwH9IVhxLSmHx3BnqD6RV9xJ8gX7f7BMtSCzQRw8F/STbtjAg13xtyvYtalDICjHNlBoPFM
p6kHASr+1lxBJ3qQe7c48/em/0CXNpNWX28vXQ/1X3iTn6c2SuMz9Al/gdOhyriLpyxlxu1tUy/7
bVTqBls/xGGcW42Q9cttkZKny+4gbQoHGlTbRYbTlLfmMgjKFdYaS8A35q0cz1oQeHLfKwdsC9ga
bMI8/mPC2ZI31GJ+xZ822DewB2y1sYvh1Ni7MaXnmaXx21fGbLZMIVnUT038K11pPQN8kHzA8tWL
4ciyDZD62dTzOK6fae2J12MvajO9+ygHpWTpLMCEt34nDgVlRWAdF8vkmW2ZagzD6QzNeywpvrH+
hwYpkcsvn74pKs7gvCx0CWm41uvSjT2/gkPS592ckhvI4NdwOwVpGvJ052y4Fp3lgmEYH4W+hHLm
fGWiZ2iZETs6p/z6tfju0AG9m0365oeQW37bh2aTD0EIS40zMimRGeS42PkmkWeywwsOT38pVVLA
T64WZE/Bl7AQf9zLg/0Cy8zQJdhUvGqcnA1SM/WlBeLrg1A45RBCLgFTwFPFNb/V1qwO2VXF6UpH
Hafrgasq89BstT1tE7k9KOcRZSha4kALAq2cOj+ddQVM9UI2vgfSRTA8PlaWFKf94u3DbX7swk8X
y+IWIl8eJjsi+k4NcNW7siRAalwRqZP9/jUGG1ZkPjOTpVD0dNZ3IxPmhJavnV8uiff9o/IHMp0c
R2YusQNzNH8hRCb/G9+J/f+Fnrh7U76UezvFcmtIP6RRKRORSgpyQId/zwhJpEkZTySxZEitWwnv
QUFNTgzqiucXK1zgzFdWjgMEXN1GDI1RhlfJ8h1B1NhlclUCsaVtPOUumHCchymVQM0dyzr8MB8s
0lI3XbtdlHG8jjreCaX5kWiynhcRhd32LZYkAoY6V28TpJEBuEr2QvOBbIjlPCPg2j83GKsYpzbZ
bC4jBNGwjj0lYsbc36s3V2CCkOQZcDnVfFyIxvMIemLWtwlr9k1IrTy3bo8EB9jYmXTmqsne5bog
Icc9ptMzOD/SIj2hCcAqRqQay85q0NTDfZO11qI1C7mIujczX7BSVuyHSEnfp5s8LF8SQusgO2wr
SIWq8jNAhZMmXq3skIvKihY0Wo2lQ5SyP2nCXtZAI715MqZUPPjWhLC7jdSzgzNacUWTG26NIt6m
34h/8xvs1Mwux1+cSZ3hsI6FJ17B96YuO8MnzkPcdtbalsTY5twVmf9721q5uOhPwpSywc5a754L
2D3wu6eteodvNp2DHyKM78gJt+R+psw6Gsm3s/mXOd9HXa8dJIQABUPmydYlwXPR2DEnZuS+izhi
9YJXvRpGwUwojZY2pxA7VSPbXKMUmL4qPTKBRg9z2uQRV/ja3rZSsQyNpBo5ZcSlc7HbyYJs6Yef
ymM4NqOy61MeZB3eyS/0gGPYYcjh+WAy7rrB5qLNRj2Y1ezDKkc3RebNFkiBf9Ci+Ckrm2cMXX94
10Hvh0rqP68ke0O8HqeDnx9rd7qzQ/qVd1Q5HPn2exMIES5pT+/eMzFk0G+8qvXz28ia/b/Y8cxQ
hmTueq1Kkmn1bmf2rZexUrzEpFa5oxnqgBaXKjc2cQlRTKI6E3SSOCEa9JTfkiOk7L+Ra02FMDax
k0R4Pso+TiMU3W2/BUg6WWmfnQ5fUhRfo4uAa/040uxJ49mq4ih6GAxg9wO6Y27Tp/p3jgSkHaeb
mrviwCdb/SZv/8YScEPy6rs5vF6R1ol0cngontCcznKrXSO3rk26I9d6cftMhRujqjd+1xMESnqN
IiWubT7olszT8fLwT2iQA4jlxd4pPwBu9FYbomGXWs6DWWV5uUu+VTKC3pSlRIAzvTpFegzh1xkq
lM7mlmNasaxBg2z06LHnw9Vmcigcfma62oO7tPhSSZzwJSxltW6eOoo+jfITlOqAiSpelJu5PVft
I6uJfrgoAbE4nkvLeNeg/wGi1R6I6UyUo3hH3UYuNIePpBLOwARDrpkR4EKj8X5s5luius518YLx
iR/c/2UpmbQ5Rl37EPFdymW6ATX2fYm5CCZ0cLwqLzYewc9/uC1OWpOU2UYQ+2ZvRzpVVPW6blIt
3ZnVQ+EYLKJzpwhTWBIhLmVtfxdwgwOdsXLOZMVQVJALB0zdv4JSxwRv4mukRAuB2CexNSEspG1f
+yNI4YL08CeiS8MfC786tcC1kqYC+HNMIMUnl5xEN9eeMSmO1hV12j6M6h3VeEyAvdJr4IbsJuEB
xpXEN9bm/fvhIxyC4AJjs2sKQMgnaw2cPXfwqgiD+5lD6p8Bu5JgTMhVLxKsx8AfiGtqKynOL+gf
FDLELUEMsalS9wrFdTIaG/NgbtLn7qb9psXENAP1qxCvRx9kobplLeadFWHVb+lu1JhIlHZkTq0+
HW4PQbds8deo9wxccYN0si20vzbsswLMkc1MP7dJj6MoxnFtYB26a9RubmOhf4T1FbAokYqGD9Nk
hHGxPlMuiigIyQflB8QufJfdwNEQ4t6FjDSGE6AUrxI/hGGtK8L3HiNwXw3oVV0Wuv8KKGt21nrQ
q8UX0RP6yUC3WNNY6gf5B9JupY3FOH5KTPUl2EXYN1O2AM/3+gUw4fkEu90kFo1NJpjsAyj+4lvG
dIhm3mdBnYRZ5qa3d1dWzloLP87jgswpoTWuQhM7Xu0nMGN0qLbs3lXxvKpqiPmP90QejYj/YgeN
5Z9PWXwBve5c/VS/WAgPX6dhBxt2ldhh443oylpp7xvj7Qw9H6wq7CTDf0umHq63PbbSiAX9Z8h5
HN2u/MBDVnYXoa9RHIOz4ed/B0ofigaNlFEOlwp7vXYoK9fWT6y55Se3N87dC3py6ECOwji7Ep8c
5xKPesgSuxQwQbxuERFprRS9zmrkaeUlhsesoIpXvSWQNvdqMqoaj4PWFwrpg/Ao14TUmLJSuznB
9ZvbI2XffpEzBC5yqLsUEuoWZZqN2V+23/CUIeB5P0wDQXtstXWDiXFZ9JBBvJji1Clm4nfycag1
81kBvXmdMc9N7bQYdN9Pobw19yQlJXAJ1de/nVg1CnCeRQONFUrEmbhsScBzJE7QScm8tbMPu6gV
4aLYs7gs9Jbg2gdVFSh/smSN/94zXbYnpmKnJCKdmLHBIIEioU4WbF9LELEa0E9wokAWjtbjqvS5
7LiOUDzqNypAen5EqlrLXAVceovkQDBOcoRLucki9zhTinS0zIzt2bjTlOxEohCcWdZ8YL+j9Di5
68Nnm5rZQwx9EWJbKYq6+4yx+JrVlQX2gvisedxILJPdFKizalk5INL5xpCRXQ+a1/I+tz60EIq7
VsFnLAKilNctfkkln8uI/defgiD26Q0JUm72LseOsIHyHxfyotwYHPzyUxxxQ0wQnE0bjvzLl0Aa
H/OXnwHdVd+e33Ww8rPnt3RVku0Bhr54X8A5R3+H/s7ErziorNszscxD7qJN84BvWTVYyH2laZHT
CfvjEd4At9YKTlePoeOwJPcKR6bZGlhN3Pk8QyzG/LF9tE/nUwsJpua7z7XhqarTP8+WKRRFG10b
cOr8yySr9LDHR62P20rM278m2TskTcUOT0kh+rq38Bg4t1LeRv0IlBlgpHo6DSXajW5T+4gUQ2m6
AT0RqjJqt5pUlg4wNZVwbjKOiOS01vZesKmjLLWRsMEKFJf+WKSmw7XOU7Zvg3B1JLMV/vFyYdLO
nS8rBp8vnOgS1Q0WA0HmljifDLpDFDoZwodrSzZxxfXJbKWrMO6MC5TvaQFZ7kk3avdWhhguyvH/
HCWw8KGNt/bO5JacRpE21x02FfLfNYkMo4EIQT+k91kWvFWCxsxRP4RFRStt1SqGMq8CSG4wD2wq
L58lVdt32zDKhN/2CyORXNc7RPOvt5Rfy4wcN8Be+rD10Jd41UyJplDvObgemlyzmXdc0fpho91H
77bNOllqOOiBEJg4bMupejEeFKBaGH+B5US7ZM54QtC5hYlW4zvINOpPtucA1J2tx0sbaPyM1JTv
rWmkiGOqCuHVoQG4zRMNr7yl0Ewqun2YjVa8OF9EHMHHDo1+xUlCEYg0Q5HXha1gNLtXJGpS8gvQ
buJHDBbb3PSdWq9skpU8KobOMrAx7bZ2Jpn1hOoPyUrCQcbhYWQeDHivvqbCYAbBd9vyL+oTbTWz
yf0NorkeLNe7452MmJdut4KQw0Vssoe6wH+NFOOEKPrJUWBBamcY/WOtSw/6nnAXRZkbgWA7UZ63
2voCXtpLWrKz4i7ZuXZnOgeSbEXRSFz7h16gA109wP1dRFchc4TjUTHN4gwl+ODJqKHBm/ynmOQm
H4z1L+HD1G6pFfYiU/Fggev+Md4keV9phr4ldkzH0knqyVaTcPwRaGIOgs5u54uebh5uxDoHjGNa
K3eopfhMWMbFZugFjNFMTZfZ9rWEnhdcrCkaS6ufNQTl8xM7tjz3URc+aQQAO2ixIenSfEYSC32k
FQlRHa/d0ZoPksEa42JalAP5NVrQnJ6Nks6Drb0bCZKsVrjOt91cZfwR+SzVIHyoOGFnZXn7j7O/
ffGQxnBDqRhe0i5+wGZlQtuf0JLn1KWKSC6k9BnBR3hIMnxE/Iwmh28ZPnUETepQJiDBtGPHzGd3
zTPwBrwjO+DBKVqTjzL8DBtWVyBGZFuyM3pFmmLZ1qcJnNhqebr/63y/Ue/IxdAMdzbI3Hirrnyh
rqkznhVHs0LVE7IVwpgB8YLlyAKP5gaZUEvi8aUfeJKoGHx6S9RZAKGu4nDpQLmeSMLRszxUtXzb
BcrmmkRV2TDbCFyp9N/LFKThTN1w3Yg9HP6+AEBu37G7u6cH7udgq5g+DjYjqHqoS0dkXfbbplL9
vIoITohNtrfaPB8/P+Myp13dYe8EOwGCFPb9Hr/THzngOVkeBJut3YGpMcUWUEsWpUsSTL6s2Avd
Dz1Zq06r3si9LQS1iw6nDF/dbnXF5chaTnCQ5GFUecaNs0TvvagevphcVLTQv7Nbc/04Ju/fgwJK
aU9yUaeua9Kb6uKFAnn32J6qfUkANvx2W68RvTVUvIpPOkX/Goy53gsYOwcn3CemdVk8gMcvdL6C
51fAYWy7I1idd1gEKl37D6FTSzuba+R6v00qNEtmZl8UglFjiqXq1NjXGolHSOQ4LM36xxCsN2Zz
mKnEJowxQZBwiglJN14zugCsyJLjw1DrYSgLQikdkoZBuzqurxgsOyKHvjsrT6qFtAg/4/BkPZtA
YWTSHEwu+YGUwsBfmyN56JS/aWRgEqddQw8rvJ5sYBxC4dvfypiDX1bXTw5jo1tsJFu+cD6W4mwP
Kv5hNGev5CT3BB0oUmaPD566wxt9NXQ/3vbS0/5XCoijs7vtDvRz9qc2J1gxk5gSK5Mc/pBBRlK0
CglqTPUowXltBV0LRLQXjgTbHn/kdNge8r9Bz8tZkVmtWVA0qpVV7Aw4NYxZu47hcm22owz0TrHR
UXCvI8YWlYh8ekNrP/1vilIONFq/mSau5OFjtDBAUm77StfaXZBVSdaNT6CSMOv7hVp1gMDx5YFn
XYWUe2Nl4naJlV25k+6qzOABZ12bLasP6Fd8+GJ5kfRb28jKnHHCoHdo50mAISBrBE1U9mne/b1a
Bu/JQI2EiBMOvTWEZ8fUje7OUVziXGoZYS+3IDnfM9fZmOxF3g8sozPW9InTbhnzdCXqFb4EcSDL
ytaNYfWxh4Kqzt4NyTg1ll5b7wlYeSZDqc2FAEAoeQ0a419kgdkgQmHlJrr4YTHh2nbgcdo01vyv
CBJQD7BJs5NVrfvZBgwPcnxDnOJoP0gM42p7S4nBTajA/o23ZyvM/xWIQg3JoJ0Bjor1p+SXkNe0
FvpSFrC0z4o2azJTANvOkzTjZ+H4gwLJ7wJXdn+EU/DzmD8SQynfx9V4oDZqXnqhx5qZg7JZF19g
pmxXsP4y88jwE9kQYXQdQrmoIMukFJOKwu5WDhrSTPCNvsqiMteDlH79wY1KnK6NMUsuMLnE6Qv/
suS4ZD43R1hjWp4xPsuebrQb7m8410Izp7O48u+34DLS0igPkvOIJIEl7jDEmsLWEhXKl7TSlONO
D5+yaKs9HN9QzMkb66pZETDsZjcQm6Y4Y9FTyMRqUhBBEWCgXYHpm1++RJQfpfsnTAIaAYosrKNd
WJ5GOrWiu+saZaXnxtcB8aTecqJEXa2HOhLysIy+x9nOGNHGTON/lIo1cKIR5TJGrWPKLg+u7Ls1
zWW9D2EFPpjblqo2gBitSic7YGfaNO3hrz24jRoB+aadGTlQ1tDuuqHCw94WGyMz07E2lMtqG12K
GYUsOYeM8vrbbdI707qnD+5qgSbwKgDs04qvHfGMg5JJg3jEtPjEVLyeiBMLKkpbE9LE7/1NZiCY
OvnAeQEWDdz/HcqmT+aCClL+bQfYsvCChmRFA+oThly5EEeLJQ7YThgfwhu1dAWVix9Qe/YNMhut
bbAXiW6Tg5tpoleZYcQfehcxHDOIEH44pr5jzXZz7MdpnYcohKv/R9jy+Mq/JALZMe7okpjUHAFU
frhdc24rPMjEPiNibfXY8qh4/3LyvsTtPgK+Muu0uyQHygOoqLDF0DYo3kc698gItkumygbJl/F0
yJMKjP4Os97SRhLEi3zt51AS7FGhh8ttFgOKPBd+W68UrkJA8Nhv/Oc1JfOeZzN9XlMeZSJSdfAR
mvOJmPlETa/oU/frlrl5uJN8jYlus0Zr5GrmJMqCK46D0YCSPRdOCbHwP48upsKFwXVFoh7n63wI
eyoc/hKpl1nf2hXdLYVJcHyunGtSKY3eHpvVs6x6Frfyl98jbScMiAcKnoZgDibub+2QXr2eBraG
iEzgqiUapQABHRHYO5lSxx5Dl7MtXUCXgAodqGF55IXiyaSfoKcp754UrNS0tqSb1Y4VuzGlNCuR
cVwmh8+Hv48CSVodNxoolscMZO7iBL9poRnGkconRzobhe5S+qODENstrWgVtSF1lLu2hKZQPcr1
+VGgJQFU+jVsbUKilm0CdERU0xFkkzF3f0CXXkFg5gGsfJh8c+D8NxJaO8AewtXbl8hRwXwUQtRv
TEA+2+/Yze0tter4eI0G+/bVabQg2iHmHLFF/5lzlowyYQ3b//mLFpPRKCtln3BC6LFtlTriChEE
NJdV77F+oByKN4dZrrP3PiXxfLgfdCzG4BmqRMaYWlY7cK9c45bC9XRc9WkB6kCP9sZSYDNsLnd/
T8IkFkEnTQrYldEyJ4a8WOkEBgjiiI/poxR76gCRO4/ufKSd852VQgPmXEPYMkUPhahk0vNnX+MP
gro8uw5h5sCw6AEEX91mTJBe5sHsK8+BiCiVQyEPCIqNHD8moIgBoNqa6lq9y6F3sSJl9qyUX4TQ
l4ULRxXfqmDUmBv2YuKAypbr9RNqitVc+HLy4mAFlQa8+klOGoIl8CCskGl6y9fBKdtoHQ08uD/N
3uU0mp6cp3OdDPXs+zmBqVghEH8ZqqDGew1Pt7zHQr0Gg+tj9JXBzHQd7sU02ReKIvE5x7JQ6+jo
Tagl80Dfrv+KNwaXJoIa6RZhJhjDrzqFBuI5mJ3U26FMYB8Rn+nDVZsOQo4/MLBMaN+ib0GHa0kk
BIWs+Qw8o5AC+bKTXdT1+6HKgqYvN4di1jzGi1rHtt8sfBSq0crKs2bFVyxtnI8oEsnCWZcn4W++
1GpeCChMwpjVjXHYI6dQAXBIsApGoQSxRS9NZd2iEJWzL7X9jurK7b66cgDUDRg+xQN/BfhzjKnl
YteszgipaOxN6ve9rD6OFueAVgYHR0QCSySyz//PmjzvdQjJhSAr1BhLnYceIgnX6hF0fWf4GHzZ
/8BdM3lVCzswHY/+PUgBv05lpOWdzLeXyxRBED2yev+ZGzx5zYd4WHLc1JN9uLZMrGf552eNAYd2
F7UvYm6MHpbp3DH3dEWaLB5ULyLvhvU5GhxhmVSf3162gY1r3n+eyHaG/FIx0QUEu5O/t0+DO10R
sH5dm50zGwsjKERRFrdVqFmBRt/Qqn/M/YUGFD6AmYYyF3I9duarhjqT1ubJ6CAscs33N8lt4WHL
wztabRBSCiDgr9KcZjAs8DDtnT3FYV1EDi6jQMV6abNk++jAmjIV8AUyTt/uVDnS55QoklE9mPPl
4b9FCGoGZYfrhU+r8DkFHf9rQXx9+Ffys7mhfHCMYcUd4RhCMGqu8UQ4XZrxc6jRHT0ZBjDvZckm
fAXZaafMyTuEvXVaqbWhNhSbEp69qVQsmXUbjKGlwC8FnyMYhKm8gcThAf8I7ORvCEs1vPdc1jQL
GW0sv2Wyzc6psqKgsOWCR2yYTvTCZV0F1+gqy6UfvGju9gQTs4eJQKMymNsXh8Pq06fm4xxBts30
qA6cfgy/lak6Lqww18fXsxEvxr1GaZjooBrmwQirDxlcQqRUaJy6Ud8bMkab58wVyYjYE9EB3mh2
tsAN37ve4VUAJoggBe53cST+Xyudipy+P/VBgv1Nb+2dm81Ywn+UjROKeKmwlLR8Vt4MBZH7YNsN
e90Yt4KgQrCCOurNrKah6mx+s/glZ+FaqSZI1TpDa5UqRl+6RXStAotq7phr/7RoRD+owYi3ahJF
9cHCYXKw90nhhnIKA7fyRYe1TAu19cKgtt27kVZENjB5UMDz7HE376N2awigx0fwOhAy+tTFsuRX
hEDkRkwy8fqbL30led6vz5pjsoyWAKurY2dB+J3TFcZpbrNs2MifiFKdc82GDUnkUMlppO/RNll5
K1g9+94rY/iZxrzPdNm6VK7BbwFOMLaFrYLmkH1qK4gLfQw5p3ngWEigSSAwsjGE5ACOiW9hjrCu
NqejYT3h/yGTA168U/sED8GMU+ZBPhFDIydRAxZCpP8ygsFpGVmKNiS8gSuh8SoGvFKSwt358ldt
6B+Nrjn5xkES/2ZrLhvPVaqyguH8GzJaN1EUosOiSDx0r2YZ48QMHe7xQncQ9KiXf8gxx877CqmU
bjQMMz7hpWqxzJpvCVsTenomGGMthU/ob5Hu0iDlgqOEsZ6pa2i1qTATryZwerDG2zn6UctTICXQ
0ZnJzEqmCSfwpEgK/haHvvkUc2ll5ydGGxuBv8cd+j/F75WMIFn4qczAcU2fNxIE9QLU2UNyJjqX
4NMgbXQb6sz6CRbkwk8iopMC8ahe018RKTVaaLLIkoXUZLTEFMQKWntZWsfKor7DUuB4pxnfX6XE
s8MjxogQZmbFD4EdnBLcxZ27wldDZKhl4FwA3piSwWYplJgdn9coooT2ZlOLTnC3s3gl4sQNynFJ
UrmPGW4wQC5QJHQRi1h54H2K7ABGDLrI6xBfhEKZjx95kbVMgh3Ndi4AOCj7+UcMqnltMsc2kDFg
hqgkrtnJkVygS8MiVdLT/s1/xjd3TN+NsKVgZeVl2LsiTjTHk8NAQMaRReyUmLFzZ0iWmUelNyjP
PexbUpPI0KF73km/AUBaxGIBdeMF8EAOcjIl87iNsE3hIh5Qt26hTupujJ0SB9OUdHxZaGAVd9D6
98jGWEAboqI51RLGrFNPLMuEkrkpQwMuqqP3dE/kNhnUHlAD6STvJ7H4te4G2a4zQVCvcWxmEb5Z
gGaBLYKtQikV1Qsx1PGj03/SO0wt+dUBdbgqRfVK/wu0OT5mnvsLBcvT0y0Mx26OWqup/wpB5Wrf
YSwdD7BDj/gXsgQ5gM8a+MXCHjIBv6sD6rw8ywvuM9cUGDKl+70U4ni5CLAd71eH06/tDdgEgkV/
TsAmSEwk10g3gifj0olFAC4DkvgtDRETflq/UlTDaK9Iz+Gnb9+fZ14o++2GNjmiaTyTwtFy08az
qLyjU67E7cPVICT9AOWVx4yw5h2cX1y2KvI2WVHcWVBY5JJLLd4mTHWpzcDS/Mzhgx3u1jMTBOUP
DJbr/x0kgDOrwquU1pud8S0uZZ03FFbifpkUOlZHb1JpwKZcZyRClWqofX9UFUI2uEuKCO9rez2D
a49hVERyZpI/5o2lKc8ijp+SLN6tmrvs73nObkEeplVIGvxUQcWEy4A46D5PrY7dE2xoNwZzR9uL
nccdPwBcvBgT0s8ibGbuVzpC71UPPBgEy2uOiOGBY0652h1B8MCZ4gR53/2vXQLSBwzmtKIlsrPT
JN44fJ4BoZv4ehJTUYKGo8YBiTD0eQzvg0OBLr07gp1mJWNpt9fZZ1K96G5mptbk0nfsU+Kai1L1
wPeV30DWv+4oJK+/Mm3RXZOgWpsL+kZEow6gOlqTdgBe/EdsfgFmSQozzO4LGH6ArPkCH0X15H42
WTXqDoaXMMm8RDtiSSTYIMCA9yIh00XSgWqQdxEq4jYi8BmLvoFtx5goAzEWWlRN14Ea0dF0ek89
+xIdo9L1dkJgVT2diz0Iidk6Bx3FvaiUZJf7d6LYlNt++DYZ3tEOuc4MTUOSkkRmAjuOaul4Xlzt
nRMj8KgDkZebhD5e+NRa+cLGZeveB4Dz4JkDg6+CU5ZqnXtlsWIQSwd3a+q8ToMzuLLLL21uGWeE
caRcEqWwFJCIeESbtmyfd2sSiXqblJlkL8E5UI1BEsOUs1UzyGJcn8ucfnMk7tbXCLlxDy5BnJ/+
Hko7U+arEEXOttwKURGoCagSP3tASj4qpQGmj7HHX1T+oApy9icjAbbnwPXpxrVY3PrBoiaoqKy1
RkQ7n9lBLEqIZmG+Q+VHzQqoSyJrvqXLx+4bffreSKlFisCSGVgH1oIvW9wRVljevgqu5syiq+Zg
if3KD2kVYdlWaE4NU0+HLyo1iorJL2wcOVJxYAjcJRq/TiqnroqCiju2I3T0BeHZvJA9t164P/YN
ViHPzmp+s3DVMIZ/TlggQZHp83l6m8eYZ5p3NV44MtvyT2Q+5a6P1PQHD9k5FbL84qy7gKjItLHD
SvBSsvpMVJ6qcEm/Y4uljxGKZ6Sq8my6Lmc5ciiVp/Hj3mwAC4bySelkxHmcuVlix1FPgB260aV9
e7SJDsy3PG2fXdkQQuQ1NfYIgkIYnMM6MCa7orzJfLXX+b8y2dYpIJJ6SS5fqlVEdQUe1W6yzeR3
Tpw6x0sVl0GEaktqwj30SE8uYGiNLLQlkdhdAgqaeX23RIWL5eyeVFVtUJsJ9DuKdjwwTDZ8lKsL
9aDUDv1zFrCVVfHayowT98Y64n+q/Zs3NFt+B5dOGH6Y3JGGY2XUqjyod7OSvJlW5tjuUpnW0sdu
EjDSmBWVKWgY+gGIaUXt6mzDV71JplTpZoAeTGFoZt8oPDJemKbHxxkQ683QFVG8hcwTNwQSr+5q
SYc8Aa6Sl6AZ8Jt2pGU4NcIwP8/ByZ5uzhj/xKYQCDfGU9JHNZy38bwuZnB3gQR5sY3v1ZBhMUw7
dgq9xtOTIrG0RDBlw3Z24+gZqWJdq/mv7iSc3v9YNE+tnj/Qkg7Q+RsTyoqe8AwTRUXvKBm86NoA
Ux9B8G8VnoXcGZhs7pcsWhO7RuegwRguYcvoCqdlj6gCc7KBYbscnBdcV5JlIMDpYq2j1uyUoBYy
mz9DDQPE17HUFdpLNMwxSbhqvV10RRFoOYbt6R0+gqvlKj/eaBKeP8HLg0TxFZvEmLs1x2bL33RV
KXzkd3/9ppjZDBvCCoxgcqCXPdrgMgyGpcPNUi5s5tDqjj5FSbU1stORjQ2JVDVLqZY680OAdxnO
qnaFABCqn7mpCXmKWYd7gbnfapEgOO6wBD8aGeL1tAIzTZMlOMLcPJy30d137RSH55iww/2Hm2q8
EDwTPzERH3pa6ojRzwx9bfa/TprdCHpkW9/pH0cTtYkoPpyqM5sB8hRlz+XNi/iI0gUZjHJwrKlW
L+4GitZN9ss1K3MLJhE6JzwUb84J2lNmHCcaU5AeE7wRnjfXGVS1kyCUoSroSWEAo+HE1enejpIh
lrPTF/kEncQE87r3enZx7ywdgByIH7i2yTjhY1FeiYDYFo9YzDLBMvQOYr43db7rTcQZDRtYgG5n
rc/+M7ajWyaqwyu9ajzL8aL9EHiDu8Upxc2/rgDCvOU006v+tWxYFdcJb4fK8uDzs7zWs4/Iq8Po
KRJaeKcu7wfCZhMesW+d4gzFiKAx6+jhmpamt4ElPOYyiYEzQwmETLctigHtk7nOWjw+ZG0vjXtf
oxPqtOChq1/sIqcesU8c5c/vw2nsyY1c6n1HlITeBLFJp+NfBkwH2o88idUHbZQHTsWzOYcYHIM5
f4P6RQ+6CDjojTyoEVspd72Q6pq7Em+HDj3bm8eyYvZLykkFSo6x1pwtQVF3sGEI0IeKwDkJ5WKg
1rIa/UUxoPZfuDMc+SK8BlJ7fRoacDyxNk/KLuLeErEDXT78U4eEpO1+uGmSsp8Pks4yzb9pHfAw
SaptCpdDMCbsXqdvWL486pnlgZMVoFTDwrhxjPoV+/OeYlfHIlaKyiUyXgHPYQlHSffTdxCoQav4
YdJ8dr4Dk9dJOFRgjNqhin6yFLjHFgOZZ+2d0n6vXw+wfbGLKGQtTR0EMTVHmKTPAe7OVn+CWoU6
JIVBR/+CSQqBOLwn/mothOoe6D6dShepNU7J+hkXGXvMvmevxQVGnB4bMKUrPvdDbSFn7V8PDhBQ
K5UoRmYo7td6R+nNm/wWctqQ9FxAoBrnfreJmkxPlsz1iIHNYc4rzfXTAci+SsInbZixwUNRwewI
dA3CD7U3HbfvM/9CqTLGlHNFwwqfPcI5B4LSTmVu6/nVEhjTJikCzMflDM7Bi/X4i7ahf3aLY+RB
hAZvN6kQkRSyBBogIlIdLjV+0QOY0msIPLMQWfxiqGE08TsB1ZttIAVc6LpVnIMDbv5r7cccixYp
009I3+tEwrGe4q2fxrWW5WgWDQZIZA9MkjgQwcbqrkkVK7Qpuckk9waqD1RTkcdLzZsZgCMKSFiH
5S2+6+OOaWJH3+q3N2GaU1kyJrmPfz9s/UlU7fLIAvYT83hcRgYjktt13Wagr6OAen9ZQEQQJei3
BRTI3fOUuMHcfQpGhH8fnyCxWA5R4pKqbDsx7mOGoYEveIqbzMOBN3iH8lw7fVIOkBYfWs06EVpk
seachf+ImiWnEN4oJMEX+GN7F4p4XpcEYKkiOSSl1WJsRAKrsZVulBKm+9eWXflGcCb3MI0u20h/
GQ+UspzbxNPpKvZ7gGSDYExwUPmfpWv9c9T8AZDf7SDz1lx6trOQiD8QmSOo4wjmmQ5ZafsB5LU8
C3S3Rq2PTMndS7ru6RlSPFofTBuJ+a869mOCji4dejyegDPQHnPQTzCm0lfHsYNVMAiRYcqzgxS9
DLKh0SUXVR2q33pVnmnfukwGk2Fp6eV1dyWA4kuqM4cIBAo3uMZT7oOaJoJS+Rj6iy/7IZy9vpfy
6q2vcJX0+rxgPlLZKMgvLOJBxNHzWJpkBo48refYje3jaCqezLlC3JLCFQd6aAlx5keCbxszyiN7
4C1c/xUO6hs7btAaFO2/aa+rmFlqoaNJ+B1d5z1jQjoHL5aN7Xs/fFsSnAVIk+w/EeFt0AC/9kcn
lOCOy0hl0Ybw3N/jNTTFHdAKEA136g8w45w1qy+lEw2IDKWSDTztPm3CVGmBGhO6iQP9SweQdz5W
78WESq2O08Y08yXQm4+dnJP6XqdQtiDMwwUd3pzv1d0ObWSb/TZj7D5zFws/FntV2ySSLUJT2mOd
NRij34FkpoIVkiPjTpEnzDM7A2wofFLLwTLaZHUGi8dJ1PkeHbbp5kLIDINbuUTAtWicGJn3DZfh
2qiJ+Wegaku1SjNZ/xtfd/xnf+HdfDgjrewTDcvzGIsgDW7bMdc64h25iviK/opUc+7l1S0jmGpB
H03NooEx12rKqHSBtW6Te9ERX3dMmfnH948SQG7+xLzBvt1ceS8/utMYz6ktkEEaui7gRXXuawMl
J8MCh4Xn6FFhMdBz60Y1dzS+lsKnTvKJ/f6of05LrIolDsmtKlCEUxoBmzJI5N6M7/TsYUeNwpwU
xrxTm85K9fODRwYQNAA0yB1ugAz9YLmznNaKSVJ81BNY3x8ZhNBxRcd+JTUQyo13ByINliSlvh8H
2Clh6l9HqfFK4HDSchIerZZFOgE8cz9R5WVqfNKw3ALzqdaaNNMLzbngWlHB4b+QTf/tNXTUigPw
mIZkqCIh3gTOzqNm26X8+iaIEPe4KIpaOGy/DM+w0KfDFm5RtBxKZy34Iw/gRVPM47QjKusRkNt6
22MRGEnvMUGB8wJQOYkcsj5FktCtLbQccQr3f8GKmWwjcH3wUhw2NClTL83RDxyndnZivIV8JAG8
aH/29oRLup1/Smc5rRdDekZCcwhDN7fpvZoyxXs6sZBR35u82tUyJ9c9X8dHNTU0QjfUiD5EuD9U
T04YM1COStRsX0Tir5IahEuAaKhz024DQyRI53dfVTsCM0FwYVr6OuIwWLT17mAs3Qhr11IYE7E6
KU/9kfmOerJiiRrvl9yIkV9n4uR/8Eo5YhBX3Wfp3Tp6Gha7qZIIofvLKkySCIXqHzguH9Ulb0ph
Jx3kH+OxrU2S4j+NMxSaSbVzTR3gBxK8+e6Gqt/TmKj0jPBhB0SEEluPFgXAQbDPYAF7f57t20/Y
x9kEt9Dj4grKLMD5n0/GKZ6vSVS4u1rRFsgitIcbE50cJ4rNIViHkMs7ROhvXK9HE+KvtzBBjAZI
FJGs4YQnVUOrT+7p17pu7pkql05uCDhpnIKO7VbLBp+iswf2oJNFVqbXOirpvkKidtFpJ7Q2tj7L
Fq6hU4SHO32s3KLrhLz/LvAD9lcnApBz+5wgWQboZUNonfe3zBxWT2f7YNnCceISREmwx4wgWObC
D14zJeVf3GghlHWNYIJomdFZmGR6/2f4QHr8Q3KWAN3UBZvX1BOxPY4QAUwe2XiH1vvlrdIgk6Tp
A9UM6bbfWOyd2FWYR2LQDmbRWQxh2HDV3rpG/BZ5ujz2ljMNcV8E7J4m58LmlBmhGXHM5ZGFVa5Y
NgldHNxqm7ltNWKOSYH281q4gBBUjKhOqeNwPKK07CzUGnu2yUCoX+eTyunQ2e/T7j3VTzJd5HVe
uQ9LVWsc0/ZZgTxBrBxudRDtFNfK6k6QrUhDyAjApyAhxICB0HKSNg60BjscsY5gk9v+RPFGHInP
flQAeFpc/BKXbBwV7iEUoh/fEP27O4nRo2QofnjTzSipRLWfztenRriez3sCQTdjhrVvucJKqrpg
GANPi5TSt00lCQBF4keLhx5VbGMzH6D3XSXS3KHkaZ9QY+sjl/oAQuupe+GQ8ltme2r2Yr7LQjOK
hlgOVgchpLLFuwYEhpeJ1AKaiP3ywaDS3ye1Qc1U/WCwskFLdtTrfx5zok06VprFWIhdU5wciruk
5ZxZChPXBUsYNRkVSZogiVuDX4/UMSpYLmO+nPXfUT2+JRtnwSzrQE6TrpwmFutnl0ai8bmOMpcN
NqRW50Yng//8NGloODdNij1sgJYrB3igspFQW5YZxL8alDU/k3sO6IQV/skNbOel74iNQ5EmDW+c
1GkIBsrm5LJvTeG4fIA3iWJkhNVEOPPSwOcQF5JT4cuOgl/eIVHLueJczIjNa2xptX2+PElmP/Ay
z8sV6dTtXRT5Sye5W2dEkGnkp1nlLgWmkNaE/HoAyAVSEwdJKroOrXBS/gSMJBiyuj8xzHI6m8lO
oTihJC1YxyDEP+IBlN+EpZrNBttVSmU0lXjhizMEpAIlNUTLpmgN+gGSp14D+jqWysD5QtL+y+DC
uXIFvtWG8dg1kJYPiSQGkDF9kzPAx/qTJre3yqzTmvjPA2QClSBupf5yhowAYl3h4URr2kP/C8g3
1qc2Xhlr+FB93TWwBhWYPjVLEfgVdlGG/wGHtKyt1svNueZnw8lDP9NnGK7Dq9XCHPMCP3LODSdt
YI2MPE+FXoYLbe0qsr0QlP0gJ98T1sqTxa8FFvZhhkG2tsbboRGcwjnSaOhgrPijofbIJ7QBaQ3O
5vrUC8Os10Yi59f5jHACALYtYJYkaK2aCbW4VJjYNSBX51X4/4iDAU4YU7DLhNpQEBxyGO62vAtS
F40qlmuW9v4sJPR6SiKYB913ehMjViTlPMHxjAZMC5KMEwEAVhIASElotApy6GLVsUkFRvCRaOEm
qfMHM49xTAeGMaGXf1qRluzCQhgRc7gfunF1WT85aHSoR7OSVStYiULk4tMb78MYEVS9QtAkQsxx
HSCMxqwajgUoUO4noE3y1EVSeLZmqouxpTcA3iVru4W6Zu+/1m/0p+iGrz97+I1F3JiwmUyLb0MA
qBbp8/PG7sni1Sl7GR6PZ5YusCrGLjYgPFXrQ+H+jSEdT7juZOslTXdC88OqP3DWlMeqvTR7Ze4P
/lh4nNcqelG4JcAdgDbIGJoL8qZhS3iPGtD3WyTumlKztaTA+1CLqwXa5kbxy5Foeqe4MMQhy2VH
2P6/njBlspwtJmtuD6IGjIwcASqGpTLPjYeftpoYsD8dpSUbxqC38emOBHqzgAOLdUFNiJioxzKI
x4ITFCU4gec83+piNOl2/GfOV1F8Rt0GFy3iGcMT2quVYFuQLbB0az4J6tkQ99dc2PvbuRzERwOe
xlKbUk8Sw2FAhWpm79tixsqU0Pl6UFJJ+JWbGoSWkAj57xiHe2ACpS3ln9apT6HijkHhL/43f4IM
vI5uNcSbgiLUt1aUuRmNnuNsCMBl8XVCLPNFcbvQFaOusFHCnCecwRGmtQfgGzYgcgS5xIr4FUg8
rCEtxuTNiKZejcCdVWHbqg1SbwwNztPpt4Xm6oRfqehmLoGBqzDtEiaRM+KycS8UYprmX57NZQHu
EKqMakzd5I7EQYuLNeUuxqXQS+RLvzbUt4HBKNHaAqfta9FUl5KigcyIfCYeHP0HwIabuM3d8DB1
90ScXJSgteCDrQ5HpHAVvYCpCUFMq1+ySKUndE6enScOeKiGXhGRTGZuqhHbMR3SyZDFymtcvlA4
Sh/aXOFAyeqw4acrArZ92GOPzuiD3wwPY/W5l8RhCGt+dCOfb8sluCgDs/E1d92BvIq4WogIW8UL
3gdXHSXtDvu888kzMr8DlrhtQFmU+vjfSU6iGII5/shfpmIxMcKat3bFYe0vEdUbSoKpkI/6bgNm
59kbSbC0svu9IhIe5+VBHs2EWZFWSUph+auIn0t2bVTglh1X378Yje9cmF/7d1oBKkzLyQ0nk8a/
37FGMtoRrNvQ32e0W8b9d/PgTTdIpbEv2YX3JC5O+MiKZI94/zfcPs1DxRgkKeazYqpw+ssICSmQ
4jIiyw9Kx9j0Zmh3vaKjoZJUV5qyJc0tuEvRla6S8rBb6YlrclU/uNIxZ0bXx3uAtxqmfSOPb8p7
qun1V07w8CVbbKpolHalAIcYYIkCl7dcKdhGq0m/pcNpB2KzLFyeB677PGqsdp6WTtVJsVAbr7Gw
yShu9jfHEuOfc8ui86nfor5qqH91aial3md/zhFqE3MiO8uE9UkoFroqxvqoUDImQV+JgGYs1SYj
pfF3Dsxac8eZfM3XqfMR5+yFNTQF3FDHsrYJ0PrVIOzh+BXg0iRUffwyCNOsFWCeXuLFualXNMoV
XRQRrLSOP7TO9x2Yccv/HDmuDf8ksVw4lNfPp/PY/q66hZHjqAjhmsPcYjK0uVJ7SOJmADTnjK3x
coOkPA+nhU8nyu+sZQdPh4FjgtJB5bRxB9WAzJXg+jC6yZED0I/eDRlB4m23yrIfY/j0HkhaZJ+U
tCBNsqZebqVs/WxYfJdPHzcyScqJCZmfuxgNajsHl3OUxzsqMdCERm1srd+eDD3gGxFKYks4Vnos
hqQGKYFO4QOyG3rKZWA+NjRLv6t9NDKBdeL5jPc/wOQVzG0RfmTRLUfCk8TYlkIGofiCjvcfFOw+
4MN/JIA4rob/9ELoNicWU5GpSEfpbSrkQeMHY7Pll+vEhYgevvSCFXAVx4O6KRJs0QSOmH1JENG1
iCjQwV2Vpgx/zB3N39zaEQdvoVLULjNLwNlIzEBKPXCJC6XOKGNHAIM1+QkiuVh6fpRwkuBmLnZ8
JWP8ZiGhAAhxozxkKkiVSY3zUKNzTRvRXUtbyyf/IcN8jaTgXNdkXmmtiwfX4PRpU4opKjrxBWmC
cAdHwKs0Cbkylhsswxkvrau5frkgB/2mVD+AyagukXewQ/kQHwQe0x5kdlCGENKRGT2LtegMAhSa
cV0eeZQs2BlXcli1/7b93TLhe8MFUcf462WJSTCbSHsj8Ba3avdtPF0VBNDs3ClM4FZRCXuad91U
S6GecKpg+RlfHfyAL3/j+CoA2W1F5dL79OZoy/zzKLeRFhBiIZZJaa89Il9+FILaShuFFVErrqUC
2l6A+oYFGCpHQ2dNcyHeEJXiG3SdoARKsL1rL0iT4sbGaAC7awwcUa+XHWbrh5ICrBk9tD8rkpfs
TPW6ryKZ5A5hyLEXNmB+SNt/L5c7trmsDtFmaVSge+udZM1XvgKGPibJWMQ/WqJYl2VtxOcI0Hs0
2oT0gQ5bTmLO/e4k5FKeYZWlhqUHg7jRaM0Nag5SHN4OtVYr3c+dnwvrZmHBvSz3grTcUWGzdIP0
jtD287LMl+bk6zF6zxcMDV+q3vyDTqQarurJ5BllpLD6qpDODWtl/Ugn61rpgiXT3kXpRdn5vXKi
FK4xzL66LRjJN44enN+N5AEvE73BZphHvvdsibih9dpMsgzlLFS+A2aIELOzRGfwQSI2aOsBhYKy
0y65MiTcOuRd+Ot1t3oT3xhCkFcaYD5xGqNC2MNGAgSbXLr/OOMp7UdD4StxVg3TxC+TymdOvch6
R2fxbITBPZ+fBhQ6i6TYCYBHhB/eBWZORrezrLae3CWTrvlRpZH/1e46LIks7WWYbLMLJHhb+WsA
/rov/JIb/Dc11gICbA9k5N+GjFqITGG7UNhbKatXddjy4v/vRqOjB0ecD9Jbyf1xoy9fFtBtMN2H
h3W8ivxbT8Q0MVqeUZWKV3YsBY2xJ9I4cqhL2+7//L7JbKMvjGoGUvIgKU4c2I4F/QUCb49LHJA0
Mxu0QP1KzBieOY4/dbI24Ol2FNzL2RYXNaRmnOBbfPy5A6c83DQfvumWOJBfIW1VrfukSBQ2DFTt
OIBoPVPGMXw1GczDySszSB5uMePNK+HQXQnyP30tN1SSa+EFRLFNousVwBwlnzlZoqSgE+JiC24P
k9vv8ypYowEbJyMEi6WEHcj+gvPOikK8Yknkr4/sx4Y3vaTFWj6LVaaPfmZijro8X49yKjcKXUqR
d8D7XrIKUWcd53J9C5cqHFtIeb9UvyGkeUuP5UxEK4atWzLRi3b8RquimKFGw45TvgeOtUuOiQ3w
Smgu087x261Vdio2XQ6RFwqoTgYqMZZdrLSC5LmuUuapN4is7ePC4C+ZD0iOqbVlnmiAHk+ueqDP
JQ62gu2PtInsLcExIo32oNLtmYIZ5My05BqgVH9bn607cZtOhL/sH1G/2/Z2XmvfYP1MoJIkCDAz
dgCNASjN6d+bSQXAzN8hldyLnk5w9PirzWwXafgDd8cNkcMeW0yrO7JIPUlLnFui4A7BR4k1xsWu
YU+GmDZQwjZRrPI4B9ZJSrbaQk6gPoQw2WtXoITIp/W+Hff5sb2bdzNK9RdbN/na1tXnFlcVDEvY
jBaO0utHSGc0DeiQnEw3xV3UvJolPld8n46Cftd4TAM07AipUemM2SRkqApxemmct2WWF2OOzYbk
5auYSCWjIov5IwrjPswZGDuPdjdGx9ldAiXIgdNhKBArHGYlKI9qfMQf0EhF/0+XM/lBaz2GvITY
Z2DSAd5FQ3XIW6joAXoHTIqpJfz7tERj15dqsRqL0hhpAR9cGV8ZydYnVw4qoDQ6WkvHBPyokexd
jwkXHHpCm/3zWX/jajHBQsSHK1eZ1k886zSLz5VhevvXJZBbP4Wf33B37KhpuIXRkxcsZ+nFN0Yj
lOo449tojAM4QAucNODlAwWa+pHU7CJp+FHJrNTv/tvdTOrSKjG7hL8Qy+rCqzRr1of7NVBXp3rR
rQgpwoJw6t1QaNLsoLIYmiDygBSLxtQ4v8DGuFhqIwpL9YtLPQjrvuPtR+j7AIqCEDdlUQnJd/Mi
wbENuI3DaNdm2YuGA3dD6tmboOVcrvSvAqLurKtFELEZIFn7lfJPoyr2BDlMWloAjkLa1pKwBicB
1/5eKGXi57WG+Ll5I2GIr2LVKjYP6IPsNXm4OXJVw4r3yrRzlUeTWfC53aFcsSxFcWJBtSynxF2z
b46ckQp898OPyJUkei+Hd7ainvHpkMNDHQCbAPPcswf2Wm3OgjowxrBodktNZiBKqN3LJX0nO2IW
6zmOSYa+6Cs8KaJhUYCuUMuApMIPgk+AlLBuG5CEpfpoiQyEThpF2X0UGtOqrQnASCAzree/dEMd
6L6IYRRu2vYGMM1jr1VQpcZnhhCAgp/4nVVeW0z2VvGC9cnYwZNd0OPjAxkaDYimR+xhAw7nBXHG
+2VC/f/Mm+KrJCC6ltEYmHXTY5AfcYiIcpRNOV/bmBlxIy3OJwfTVyIxRvWzCaYO+EH9c0vd8EPf
FYVXh0RfjlePFZNqFIiLvKefuFtweb0w1e6NcOJmOXm+fp2PLXQL0UAyz0QpDPYpljcrMmLAJzSO
oahI2wYY6PlYXKnJsJFRNJYCSqwXHI6f6LNmFgXI4p2J3QLcAgrKrEHauQgZ4az6FCdFuDej+6ZG
whi8hWKaDdJi2sTjBj7eVZMUY6EJ1buogK90ISqEQiE1NXxtqo0eyyo49V30+3CdIMcMfzaNp5zZ
/TeQFLTb5uYbDAhOHQYwf4gR89Uy8x0vFj72GTa9M5A1hAMaX/Z+ipjsgZtQgh42VDPZ0AwJKcgg
XTn4YiuxlApqi32ss49M1AuH/4DzyYsN8eTmJes0F3S4zPTGTZLaMepPlmKwKpQzwF7oFoyexrsb
VMMas9GggjoFX1GUwvO5ZIWrv3aKGyJzxGGLc3tF6O9nZTpNiwlaamvQdvEqD01vEeMSFM2Z/89x
J0PwCjGR0Ni5DbdWl5zbSGr7EnQCu1ydd1k+nodbejjj9j340Sy6pidoEesJbFzQyor+UxSg346N
8wHM6M06+BYGgdSCjAP03xWi0jd80OSMFV7QFux/iWgpe3ZGZeXSNIc8T0mc6RfcI3P31IooVOD9
gXYNThoWVxYo36HwiMJ995y4D9V5lWXG+SjR0Q/E9QlbtcD6xbeK9JlEr0xE6cHJWvC8nKZ+UNeU
La/O2JRw9LFmRl/K1KrIwrLK9QSdPDFGASOTxnZMLV2lnqaFLLZUbm1/1XmYkD0j6VuUp9q3AKPD
uv+MMLdxiktvsMPG/Fxm1Eju5B3G9vSp7LmK40Jq3ejrGCrqiyis06E9CFDB7J5GP49wb3TEfGzB
rg3V6pBvCcX4yjiaMIJbSIR2wNpB8fOfvtieBMTqEV2q3LghVoJrMXKcrGlQiJUcxKgOXOzlyClG
HAHl7vIWE98ZrttA/Vp1T9AVuqZADgamxxKheqWz9D32N1TmVaiwN/mbRAuZlWN6V+nyTTCzYcR9
YLkrKCPrRQ9u6QD9F0AGATg2cAOc4QGZ5OBIxGTV+ubMiNXDP7tfCZIV+P8WPMwp7hfOOEhiBNDB
pU//1KXXI1ft6T9MZv98wkV0TMfjNwI200XZb0VBtody9rGHMyCwcZRW+hD96YLu2gxd7rnji8Hq
FIPeJcGDyTiaiNWaWzZOB6tNBRYY+9t8xasDEq8Kiazz87/Ejp5NnuCTj3DbdrEzkMSZZo9TYvAN
E0zdm0Vo6P0PoySyN8Gd4yvWig6qsE7y9zavI6M8NkDD7ynJECeL8FKN8VrgEOyKDdBZwSqAzcuM
7ufrivvuJHFjs8JgOHKYqW7mnLv+Ojf+QgkuO+zXL7bH/IL3CZ2kOH1mZQZnZ+dgvNU5exG0Cb3P
yLA6ZVShGGuE307YiW4IaV45iY3gPDkOz0568IvZfRxib6hJxoLs7tb5spnS2jsGKcpijlKNSfTv
w3PsgTKGk+TUj3qqqo5rac4m9rNEx5jBZXGuD5iUuQYKZhg8U2jEH+AAWe5KW5xPyBT5arxVD+JW
PTqXn30zG2VzdMdAdoIbLQbHorxhZyriKx9dFFPbt4dx9qjunOjYFoWrEsVB1VaFCsgy27ClY9GO
6ctGsmvchje0/udfMbLIK0yfzLMuGKVlbipyixIEfkQEIP+0yOECn0F5xlDabkzzk98vi5M3RBM4
ldBFA5z23ROAWT63vV8TvcZ577Y6zI0eNqcnu2nEa071aXA+JPwlOQFRFRhTvtlhjU48bSQyMeGY
Wpf+9TZHX1SXiJqNxFCT7G8yyvijAHdZctatJdxVj2rBgrP0TX1YsgDwO4lplYrpTzEBILZ6lpl4
PKs8oFvtIy5zrrlWAPi602ugY/LH7p11pe4uQTs0xpsBk6PCrmtQpM/AKWpt+kK3Zu8f+GanID6N
RsqitsP/F44JkAP4ylMwM7XvXUFTZ6L8ZHmVsrN1E5m7SawToAoh8eLzA15oRBtvIA388GY2BfRR
3YKrYLYjWuJhlD/VKwY9YaCrnD9P1YjwjyspurinFldh6pwqrvFfvVaMeqr0zckMSEA9Fp/vIVbf
7eXuLdjUZM+TWqbMPvBkZ6KOSNOOp3Z04QQJ0SS6mKQqUjG5IUCHIa3rwGR6CYsK1x9zYJn8qs9M
7NV/sZlalA5q5th7B+DAdkKZM+n133D4WaRQgSeR2ehL4CQD7KNjX16A7fuQ+JxgdcO2jo8c4cz4
P0MEbFMk1Yci/bqYMXCIv0PbrOVdPItaQeqMHLRZ2ThOKQijGOgsLOOt9OOScSFVeJLiB+L/rw2d
BKtkV+BzrBIRO2lr2ixU9EILzOwuM56A1dip9dQdf36sgVSy1mLwK/JdesNY5ansHYiWswTc7+S1
mfrvwRqmSr/JHOjihNffIN2DMgm70V93UlgJhgpLP1LGgcHULa3Ht4o6sDcMamqe2gX9ixz0GQ2E
yxQoj/iSMmryJVm33qH99SgBNy3XlMZkmiSR3/Sd6Ws11XZZdv3JAxizz+BMzJPMDlFcR7/8aMrZ
vxn3BcJStw4r5y6ae6dq52ZrzWDU9sEdFHGuTmfO2I1fl54uH2TjroujxcoDcLCTdCSBNaMfQC+S
0JHj6emz+rxJrmQJGyzHlsRV51xWOBVT2zurQxiNsmrjgFGaXhj8kYsjeVAvYKhUZrmfORgm+Cst
QgTBX5iuLIwwpk0uvg9NHnSvh46t64D0hNrF/zxLwL2Q/EKyaPFQ/eCDSyMCMw6OwoTh0rKUHh03
Lhbb/jRFLzXX5dLgV5zMvoeRbRqgRNd7DFONTChSkafXDd7ZMW+W3e+KIHxAB1WIVgYQnWAI0blI
oV6+ZOaSCQvIaKtjV6Z4S8HnBrCwznveUF8W/mE1+qndmQTEJB3pCaON/PfqvUzlD6Xud23Pkwe3
9Tq3zngSU8uVVM9C9ysJhvR6S9UXqU/Wp3CrRPp9xq/APbQEe0sF8kxRFLQXVDNbmoX0CB1CStaZ
9hwq6mY7W3BmqXTyGoPSOh6j+RpZOir6pox0KVCTXU6tgFEWkr7/iGchytBu73f/vqbVpc9I+fIO
YyRC3MPxEAOIZddo0kF3CZZJl2zkVPzClcYyHbOtHEyyeTBsNBR1xMxtQIdRhWYXIShiGZZty8Na
uxvOddQLSW+w4MXVOOzApS+ti2/5kCbCVuuX6nybeYOTlygsYkkI63FMjyluy8YCuyNzQUNCpyU9
jZNy5mxxml1cH1aPIVYKSAxn3MGAbvz0JTN1w84UzYgGgnUxLRMGTSiau4hicr9upK+b8qQyROwS
t5Hjne9gErVnIRohRAkdxi1rxKfCid0mAB0L+76+G7LmLZKINXFUPfPYqU0cZRAoeYDcKlwaIB2N
2UGjJq+l5Zn5BkmnINLt5jpGQdGfmptpLzzgj4hZg/frfkuxXZ6FDgPfgrIE7U6mbm3c4pw3csAu
BkKE/9NZ0bQdSEMra+jE6ztCuIMYwY6pbwZYXzqRfil3KOWkU3I1B1a3M7dcFB3Z2D9PV6hEGNSt
JL6lS3go8j/WDFGQjlx8ikg3NUov8uf1PN8cyMdg/n966uHIIMm//xtuxrQ018j8Vjs0sq/8g/Vs
BpRvnotX3hUmjw7wasIZzRhIXwlADLSAkW2M9cIcdS3GrlCwpUUDRoyszrbDuRcn7yvsp+gndNVk
c1nvZWEZdj8wJ68cQCBEQf56PDsncdC2LaZLYCInVzNx4tk36E8IWviY9X4WKDw8ZHCBzqK7Dl8R
J7nGgqvimi3x66Ef/7sd3FZNdrc+l//I70H4+AKwN+X1oTEuMDqE8VpqEhD3E5tbHGfuvv3KSivG
wnq/wgTyStnF5srLUmtIvuHJGTSkrcnheUJHk2Aq77b/5NwUto5NNkdAGONDI8CXnjRdIFEsaODU
8/yf6efwBfQ0eC6fFDpAMO1UGd0VLIpNVUPxo5QPCCIepmaZCrNS3cfkevh4WKsrYQI65HGXGx/1
lXy6HCuX9XmP2Y+ijHT2pbzllza0YKBJ1J47YggLI/6kFN5xpFIqYGh90KirsHkV7Cf/rWv2Z/bu
wDOHkNTDGHfsyiZG3qbJSuwpW3Q7J1WVXJ8zKuaI7vROdJ9LfW+yxahRtcMZRnftkgt550dsj53N
uave0lNu3iDdYerH5RFf1xWMdVbTY8ZuEB7qp2BdoeygWQ5VRoQBiYlhNNkIYqf8cAXEyBDEzelC
cHDSwtHjws8diKMF1a2by9Qh18iKiBT7BP0ZKFDYuaR1zCdsR7GhsCml+ED9bwlc74B70YBQgSSE
p10yI8r2QbWxRZVJG6KXxoEDmwA6pMWQdFfNrZcs/kzijW0jhfodEqILiJ9gvu05VDeQj4mJcYl2
uC0GsWJaEmBiSx+NI/AmiZ6bnPLUqf8ZEy7J5ElU8WLBMaoOKvYU6WQRWJ4Ae/9B3aO4FM4C4sd2
Qwi9UB81vfmqVATG8jrN+V/95wir7GyKxeWXG0cOLwH/+fhEoKv9nUVW1rEYkL4HDEf5ioNJgUp4
LRJlxgFRcdTAOJsr+7BGAuDuwF1jEwTy/319Z8ggb2fa6ubm2QFvKjLSytGwkKOTzMGAzJ8QFw6/
Okv3cqeLb9E2f4h2sHzvGtUrzFm2rmpMmA6/3br8eSaYqsAFetg5b8V0ReFK7kJoakI0SkgkC+co
rn5gsr1BqkOKfa+Sc2GKrJNfZbTSBcha3qaOwrKFR/zcOseXKO9DaXhz8tEAvgjz7qPDdnw9oEXe
N8VuwuY554g3eT5R7nW/l4Htgtt97BqG1hJ8Hbq2y+LvIS0gQgJrwJ5zY35JCrwj/PwVS4rE6Y4f
TLrgzvuw1+65bOtFvbwrKhqgMtQb4jHVwHY32glN9otbrQ0LzLzDVt5Ug44qvto+tymj3Ne1gI2b
pvIkXuYmZ+eB7pGx3JiwIQqmMKmKsu+yKDuOUlmlZ1My3Xxdj95CO01EB+1EfHhGjlPcdogcVWb5
OHMphZwCUMQCUQGTmb2tKXBjZEJe+iBPUn5poId7YEXy3ZY8Ho1ekBJQ/Bl7nlmIKpMD19Qpvl6a
xjkQyRqypVLTdMWU1YF/U4pEnVeeKN1aCq3cCXpbA7hF23gdQM72f4WzsJ0DHcgAecGBVkB47fgI
SjyaiLtbfnnHJAdkXMZA4nP3KZas/D+AMM2FDX0DTHY6npDRdK+58qL7sBpYO143tdaxWyDeGkKZ
SjNWjSZumd9Sq5AH5+qlB6o/KN3AYyS6FweQmndnekW7F1kcRZgPTxbEdZxEAk9ogCADNa7hCHNP
H6WrO2iSqORGFa4jxzqWsLLoJMGkKtwvIUYpKwOaraCT93LNT6KKjuUtFBSeoBq6R1WEz21EZgC2
VqpOSUP90Nf3PHQBa0nflHf+rqxDb/mTfoDQr3Q/H+buWVN5efIEhD/x3D5QG8eV3yTMLkZUGgWx
SlWvJeWQ7Qv8rGFIQs4pRjNmxtwgEvs1k1xGGsKGXVD3VZ8EP7OixoOU81WlXXdS3LMjkAwBLnqO
YZy0BhThJVA0DJP20g7rPD4cZBNH38W0GzYMmcQpFLrEy7+Dil75uXIlLMWub9FHULQmRUurNycs
PS07X0xyR9P4s41GU+ENOIAP++R1pRGlV1iIumPlJfWAYPzVssDOyMMurIiS4CcNv0iIsbgUQKUN
+9ihKWSS4b+ilyk/kgyxhf+C16GEV6DjuqsMlfchv+Bmbduo25s794TLQg6qZucykuXLH+j5Pi8O
c1YQoElvalRyqno9OBywx9Bti4qQdHIB6k8QGPqXW/DHbfy+Hd/V2WPOLu4KBtsqz8iVYJ19M9O9
0Xfxf/0jTDpZzNakC+0KVoVY4zHYwdNiCYfOrBsEc04P7sKVaJ24YmrvhIcWCZ6p66JkvMu5/5gL
nqlAOTK13ldCNyrOqM3MHO+RlLu1P47nMgAcPREzHT6vN/QlFSUCOZZjg8DE4RlmC87WmvcZuJMi
Hvx/7ZTkG6lGHQNstTubVg6xaikp8cZjjZr1mJ27GQPjbkZq7Jgict7Hdc9mx2ZxSI9qwN6i+cqn
sq5Mp2ipk4jWhYbab+JzpmEoZgjcQ6i10D3KabQePDcEe9Nvn1wyIwvrx8hpMBByqF3RBYTNoToY
Z+oDh5INtDsVslXtfVcl+QJDXuPuUrwxcf5Z+Vb3APgk6QV70cwpuYl3Rlp83AXIOIfv06Q/88YC
munTAE07V5/KRS211AoIX+2FCiAI7MjnGnF1lgn7MEht4x/ZVzUK+oDYy/4bClbRvFUOkm+16JGx
1mdF4xnZ/9VR5xSag83fjycw+3aRFPpbY6JDUxILEcNy0E4T091ZK6MtPQbXClkyrxDHI2CarbjB
JqWhZoCrVyaJt8E4vjSzTWRyypcbO4gHqB0axC/57cfRUGLkvo6UmT9PkJ/871NcgPrb7lO6HYJP
n+8ZbtgNZ4d+9bIj/Ddfy8PBUdhvK46i3/3QLYW43A+IpBAhghlO3vHwkOsjKzojW/s9S0S8doTG
Bjtfz591BP7TEPh9io87ARtzMZUJIIiKuCxyCjAqX7+uZJwe2hN4vwfCutxuALXuf9HLm6xHekK7
jZIghztmVCZyhJyBRl7egzbI29ZE8rOap1FMaRWrhVewZqP1x1EY0DC6QWEisP5Vw0Fn97t7eVYm
EiHNoF9n0VF8reZhqmBykFkbquoWG0F8p4DxHit0FqXpbq2t16QvW+VvYUOnW5/tYpedtUA6yYVA
ewLjpK6wrTgW/HMSi7Mr0UP4/nQCpks0eClHdCU8q4nkEKM/UK31Vvasdq4t8LaNsS6tC6eXCHSN
AFeBmdfY0tGQRDSD1AYCJ51XUv1zy+5Fsj33XTytsdXHwfcNAoH2Z3oU6pEgncArTZDSfbTmdIsz
XwEuwPK+qQnrpcVF1KHMcJFy+KilU1Ev9ctumGT2tDyIDapX/32tPWapudGt+4j1TRYWOR5RwkEw
jwbN7GFI0t1FLK4LWuGnkQMcHOQr7T8kHA8XwzWesQttiujX3ROaHCWnC7uLlblhbnOK1rLeImg4
nCYASPEyrJDSGFOg22DZWcNUMOrL7EN9VECihy1ZtItNbLDClzt2Afy0hBl0Ig2l+5ifFeIUedoq
srnyi2W06jMXeB3gnSx8pfdfBGoP2lzVNDOYnP1cD8lmwlETzVRInmvjQ04gxOyW7oFRHuIfPYJD
RCkXU1YiSqtlHXCjxEoWv/2JwIY1JQQnKcwyvVpdtZ29TZJXKxajYAKHu+4RU3pb/0r15r7EAw/r
SHpnUfJeFNbIa8jdgBIjFyHKLr0r2K5qEv6jy1DFaSFC+N4XuSP8OAtyWZZMdvNqzB2r1Tc8uDMi
ZuEqZkD8+O6laWw+GtQs7g64Xg0cRzi2UwlY354692QYTUVoWLxLFdBadZdQ/dRW+2iFFDvDJjLS
1qZ7vHAIYm9ELXd0Yy0jFJjdeQIg4vFnFHqvdei/kyidEYFXltq0ElrGqCyoAEfBt7MuKhtmzqsS
OSuj7sEA0MRQyQootQhCbbYSHycEknmyQmVhpCS8nM6JymUucDMWHvatxWaxiJoiRVBkGsDe4vp5
bfic+W9ejMFa+NU0Lt3qiwPfnh8jIqT/tJD7vv/SN8aKB+tSJfEv7rjfdIBb/w5gaa3+w4dq0BrM
EJj+4kmD8Qwzb2LREwPRwsREmuISs3d3TK6425kMxvzPTvsXy00WzTHqMbcr1IovNTgq1Y84KM4S
CkckMVPD2S1zyE18k8zAitd/gfgK9mASZcHiyuhyO+nJP06rrAIdulWcBdWkix67hpLtE6sv3jQH
VpdVpWzybvNpBlvATxnYFcyG5Band7AW8GhSolTXyxKVMaqXLCWnSAYrEuBm7Etd1gdN9DE5LStT
fiS/uL9umUzP6fn6reBXGpjRG1cedj7GdomINxrP1thTj0PD97yjM9FhwFD+3K4klQMceL4qJqYO
zlahwISVYiBW1js2ixB8rGjlMQ1VKeu3HooX+Tm6qVXZWKDu1m+4DrEw70rClEXHY5/6MFECOzmG
/G6h7eRB3Ox2iyMNnX5IU2GmR18YU9YMJpFISmqRN/VHDHLA5K1PHX3lkHFe6HlSyc975Fu807qL
/Sw6f+5Mx4fy1219QLnSw7qmkbHo3R6yBAm5RsvjBMRTtAJPwORXXUn8S4ZHCtq06Qn5QoN+ifll
Aya5iIwUiXHj3Bxt3fRPKL9zN+7IhN3V7Jm/Vrg+fH0VM2XObOPLqjaI+2et5fltIrLq47znzo+H
A17grGoksIA1sPFhuNxpKTGTcyDZmHHhfr2RF8k6fvsXLOwPRKGFttS0fZOOHNoY7m8lHzT6EtF1
gFqCubHZCpydjvaW/eJqCKjy8RmkUV/CHOhjo3Es07ZjA9KxyNJ2ckISINhubk4h94ef9pL3EktB
YB8NWbFKqjfgk9FYPguQWX1OO/tcKVsVGpX4ZrobhpWEef/vFRsaujunfBKcYpkrkuXAOJ5MFwy0
CcigA7Cvlq4IAqjAjsHD3NwRB4NIy8vrM7YP9OvzLNjZb0DQRsMWsYq1pu+1WkGDzND3LpR461JR
Vi138/YO0KXOXafTHO6swzc3YYu3eCtQEVIhMUPnGIzI8kdKsq+vbylFTzYE+fTLA8nDn6RZBdMP
02lr3qV2YjRnfFfnCyqu11sXfqpEoUuOjGr0nUTXnmpcTGXv98GJztkMJpr7lv7ESB5+K+jNvBYg
G6K821JocMT/w/cQMJJqdz/XzhT4ePD6SstY5iiZcpTVE1l0EpkjTnxwbcXjwDtdgXgGNn9cwPF6
dzUQYYcBfVeAvKHzTzlMVe5LOa9MRsLs+Bg3EvbcgxakeMhYC9PUxiJY2vc2AWdLKOEbeWw755my
LdnNGeAnfzfRM+Fa+BYKfTnkCcyX2esIcvKBRv9XssJnK9g1YdQ7SAejtAAKjsfoPe2PAU2gk7JT
xzbmeBIz5opr1KbbrjyxURnffrDxCSH/WzNjehJ9YrW1zdTuiQC2CaUbsq2Ph0HPK7H4FntdXi1A
V0PKHmuTiLbs4dv+eHSFPEyOFEqrmGR0a+pkiHvgP0HzsAzB31MoGrYUlN7DeAiY83Wyh2MtP4yS
gDyVM/lhkAxHQ5zUpD7IggMCQcUlDhPuEPQDxPwUI10AhCmuoWXBQNhFcLeKF+g3mE+ydqLU1dRW
LxwLp/q7rZZn+CuVWqlTRds1CxDibjIiRnlBET/49KWgRukXdtLztUjMxibta/Y6ku9NYPFlGCvr
94t8lHMtlu3odSd/bELMsDRQO9ZYstlEBa+JY3fV8Y2DEJyz62s9V0U2Ng92whkCcIy2pms7fEvd
G+rD7EjQh6FgrxqC66m/1yAnGPVy5AOAdC/zz08CNVzVuwZs2zt5pMtQeKdzzYdjyL96uH8oTN2l
uo7R8Fl00zngXeyvyqlP4P5vh+5njHQFRN4ps9C9x26d3zX0fCBJHFKG7+6mkXXaUOXa6qF4lc6N
QIyl71r4AHo68X+3lzqaKTtEtOrWRr0w9R8zuMx7hor9+lcUV8A9585+/171aH3JMCW09rJc42kT
cfFCo3PAhMY6HcsE+BvxubXMw8cFVe1+8M7xQC80TUDUaM9PCF60QeqVWGH0tQTX5ESd7ZcyL5jD
cZzY6TUk8/6bFeCxP57SYyYQAQKvSIWWZl/QFk+gCHNY6Eh1vuL1N9nGqYmPKhLR9BlhFo9z4Sh9
AAChQabKrE2FoQU1ElpcktbDM8aaiYQymeNDSvupiRxf1OgO2b4/hTQwRE5w/HV8eC0RW/6ZE9VL
rJRKA27A0RAijhPXNZfC99XL83ccQ1o3UPodqHsLHycj/XVqzWYC7xF971M/jhri8/nYU1rTxOUN
L7Sxl27h8T9wVBw/BS71ceyPVWuJxnxwpmmllnASWn7k9VOr3tA9jI7XOur9FxbQZ/gto5uVJ/mM
FiGG5vqpbtxvfQ7JPKguIAeNjnX8O/OCzuku2l4tZv/Z01dhWrRX1q9FNKduJCdPEqEPD1DKTHP1
XU+YqEuIhVIgvjAmYeUN+euhKmjzywr0VAShEUJ1zNbOqPJZ9DMup3Se0e5PTJoTso8S2XUl0fUm
3rCWz4/Dpfw32ePEod+NbVLxs5mIOdrjT0J9Amx+fQfZwresZ8pC+j1n6Os40iRTVVaL4CY+IYxX
F+JdFWTcf2DZIgsxt10ACf6gN3lMTwwKBmpfL2pjwUkFa3VnwF73gN86vKLOX17FcPC90L0+ugNm
iIlid+vSYh7/bWpAM0MJXQHPP4HBriuffIWEpcFtNhubVrwaEUiObQKG8/8coRO+kDZ1xIdgWrtG
s4ny4E2YcJLAp8hbv/hXoh+ILhl3q8xfNlizaOj4q4JOuFW/0KS0ktTxlincqb+ZplAFb17k3dLR
Cyf2Ebm3HhndXyZPDC/fwTApTccY1UI3z61QzQKKnnYTS9zTfgYl46kuqiIvig8yRLOiekvNCQJG
QrHDezFOL3bZQHP5M7bOH+DzU/U533LAqTF0Iom4E/DgZ80i7j3Kc9D+UByl7Q4qyutmu7/6UvjL
W5VwJh2nbJxmnmvukDs27M0K1/tP+rry5Y0FN/jo97uIxDLwwVCifPJRv5soN2Ags0RLZv1dPNJv
EAcpT8CozUhUn9Du9rkEe68kT//WkdB3oWEXE+PgTbAaXG4ldUt93To/MAbeBgjiY0+gwKhRMlN1
wHAozHkc4AcchAuemin4hzXMpG0+ygDyDtK9VDdOKwtfSplwUiELHVgpidZippKJsDv5K3j/3JjZ
hj+6mvFa/Lzdi1g+e0bSEADsCgHPO3I8KOD00o4zpD2rxi/QeKx1bHNt02gmrmHqcmtfeZCqhIAc
PSjj9VCmMIPDLDJcufqEF42RfBXuOw9zlzOpYeN9bdv/N+x7pC7f+LIBdWUTM/dZTSqVtwxZRw1R
0ZpkxMlyYTl7AcRMfdlMWsUDB2j773eYCVvQjy0X2tnO+GmIy83CC1R0tMbJzjFNtagLGLPaLWaZ
LghxABltwssDMedgz09IHPVzwztgIxXCB/5JcqrtS0Yj/jUrLK+L2u9wbIm/qi581WVZAvsBKgTe
vv4gr5v/8sZRDz6Dk7W+p3BiA0sZqcnPEWSBrVG1SpDrUUPZhEiVH+WwDBGC4So0SYt07Zzf8L3g
bBVOOz0+Z2wWQKN60nTJbRLATO4p8a35vysGqfVn/HTC9jALqx8ohMIp1pEOf2+72uAqFxMtTEfV
+0m5yNtB4JMzJUo6cXqczc7/OQUQs7CJTKb0XyqCJNa6S4h0ZZb1B9EJWCtC5HFzy7kGWBPvcGum
GPyMZDSrDnCv2Rn/3MIRxsItde/CZ6kOq7MyYb23GrK7DaskPg/bi/i5qvqmCeIjC8ZX0HIumXBy
qaeQ5PbPvxmPrhXVXoVqM3WqFGmlgXvR6COwdiTrM/grybx+JIpx2sh+ftrUttXPbj5HjpdnrHnk
xJeHObRZ6W3voAPq0zcjDp/Z8P1KYaW8YOtXyOjXv0w58ZplyhRD0YUzmJi0zFzBpzYIkvNWFBUy
AGKD9hiIOttdWtGNx8jfa69pfq7C51b9K59EVLRpOjPU8JwGQTGlgUrsxKR0Y83aaoNOv6qWNfLr
7NAlG1oyzseWigOzFSQ2wUWGwhyYtrhoftEiqAi/d21tV0G83XY6EVvv1D5tHMb2PA4uFESG6Wa1
XgPGHQMYRC9OiycFlDMJhxD0m1mUYb4LkJhJyPpyxJBwry/9S0lpB/vV0l6wTXCQ0cVisbFa2cuJ
pHZyFjjaY4gbjf1fWG+/bRjzVsF9ysRPDM+y2v4jF/QbTBJw36eqa5leQij/RF2rIlXwlaEh8IX0
/lLmJrylntFKnEDj2eaz5m0m1pK+0NsYqEtscbpmbKslt8EHV85SD9QLe3bV90V1j8+lB1FO3A2L
+AgaBzZZ/L/WxcO/S1ltny3YzFttmA6AwlZhdkhTE2kHyF1QVHKKB8W8QvcDeuTlQkJ8m9zDku+p
hDAZRiMiUMwFFuXx22xVdJGWd8qmwN0JiVpfvIjwohuDLTz+s1vDhp45pmeTa1kcKN5Eh16shsEi
pOEmso01+1u/HkyRWQNIcg62FRKYraP5u231bfztvk1q1dAx4TmB63/gyq01OfRnBqXyTx9ZuuDp
7j5zVwDgB+4PJ9iX6JrS+OjIDAU6AclF2y1zL42siPtKHHHqx1ISdysCSO734XbSY+p00LW2Swye
1jeP7oQhxw5szx1k94A7dAi4bqNaRoppvoB5+RkW/iyNAe3eZscHjROeQvG5jJ7Fue5WjwFb0H8I
51Cmkb/eg7oZll/WojSBxOmopbLigNG4LmMwVYXPXuYaqEWN9KTNZqyfRW4HZMLgahjGr7gfD4TR
fegBRgtpRKYiV48lVAAOTpnpKLZjupn2N4+B7xWoOtM2eNQAk1MFE0fwEHLxT40+7pMWPlEkMgbE
MPf3KSVVuAG0+iKL6p2ZBblVd2ByGAgOM2MFKjcEKUsvTwptBEILVAkbCgc4HRS9gNfQVBTB+ii2
drNgHbmTQWydnlh+RJtqVyE2vTunfKjlFRpYl9pj+wzl/lPI62LKrvFwOXYi7RFjh1l2nLKrwW2m
AStQc9vdK+9LEJ+LkTDhmvfSsgkgvu1PuJG3d2h5TibpCMOIiVQYio1g2RyHlwqrNQxi26PyiTgk
3HPEHN16FG526dzuUJxyagjSXkeFV89fYM7+Zk2L+a9oLVIll4Mvqi6bS3cbOlxLbIFdZvs2pd00
hMuWsznQIJuFFfyU+Bx4UiUR9GYaaiJlElMkAWC4OonYpLMhb7+DIDilSRdltpVJlqe3XWxk+OfP
2t8YtQI0g9NG2UI2AwbN0qlvfZ2nCBCpG/z5ySfcXjgvd0HXObv86AwvAgl8fHT/Xo6xRwNFkeF6
iOVQRm2yGHDba1A4L9ZHUiYlC02y0ftmDKL8DsC+7tO0riDad2CngIIIVu2jY5RZ+XP7iDH/moTz
Ad/2DDajp99SJ1PPef1FJbeOtsM6/gXh+Y5ZSQJznspM69nSzQ0+fb1M1M17wbe2dFIvw/p7SDgI
cpa8+sMARkRq3/kOkIPs0tcwMucvBPiU3+RE2Xp8ipv6r2vusCmfWnjjB1FFyRJ6doUV4Y9d/8Qw
xZBJw36UTN5FxZxNfXUVShaxB82VZcqxkJGENa0ez9s1UQqqmOt9Zr4b3fR4XjDzDvLL9r+tFLcf
J6+FMtyyZQGnSsIErVL9peDOPhojrljgtx1shuW6Fnz5uubJMng7QQork/2uydgQYRcA9m0g/oLY
m4eF1FhHEt6HzA1Mbb0DYGRJW5hmqzPtlUJhVKK8ykrUfwgCDfaT6kKsNEK8Rc+mK1EnV79DGAjq
2g6C35KKduuT9SGNr4LVvsIVyT3u4DlydyGix7aLQixptz/IrDBa4SHyoV8e4srmauzLo51CZDsg
mVMGlqSS8lR7LtCVIxOia9LGtyfMx8dgAqVktn7k9Mwq9P3acySjkC9k740/iPZNbeZDetQGOxX/
nzTOLdeOh+RxkIL49enTj7iEti3DzwpqZwDENXVC/zX3glybbxRSjYVvMvZR5XNx3DiATg3m/kAQ
sCN+xsfuQilBf+CuvVS3jZL04+hLwKTBwHJC3PmRL07qEK6kua1985lRn9f103rpH1JT7LF1DaQr
xcD5RMKjczGDrh5Y7duwlrfW1LuX1cDTGlhaDG5VMcFbi9eI+mxZr4Ix5LsXFLxyha9YP3qmGgU/
n9TwaKfCwSu1TbEJVl+H8DCSFP4Nv/hoCBZlJrEwxOKjHBlKc/AROGLjOBxTp0tO0BDtBGxQp5O6
Ow81xX4rGGY4sALfQ45JTlxWIlT2O40UAII7eJywvuLWekj+GZL5U6cdofOx2f9uT9PNa3GcKzht
uyPaeS9F0Di1t38NxlqJPYIYA2KjpmFatXQVvR5haRKWvQXLvpyoTtk3M5JOZbYSkpgSJ1UaTKfx
v//uRJZ1lthzRCn5PRBgEICZ53F+l/RnfzWTHMNtxTVmu74NZGbbQDAzvS0Oe7H+NPe9I8sZaR68
G3Dm/pDH33g76ssdwLMgnD473xNyKc7n6jo6ltV9DCE/GuYppC+M6f7AFo9nY/kSpbOYtTr+JCQX
TUuKUBvXyYqTlVj9ju7fCOITp+k33SJJYnrHBTzmCA2tbSHifn/4r+eDT32AvdPGWqOPIJTC+VrU
6MdRxd6cc8pjg+zvYBedZg9MhumRFGIOq5uWLXYxI/iSPfmRCZ6E2i6Ar96m2YxcuKD1t0rFPCni
33cRxcugTRjyb8wTtiladNolI0eDABPN7WSDRIJugWUbR6OsUdLLOnJMvO8PAnPcMd/YhqlsKxjx
ab9axcq8pxfPtNpVAPOZ7FlFQ1uI+5NFbk9jsTDd/T+ggZHsuJyhu1ZyJZuYXti+Jg8XzJ/YY70I
Im7eoYI/lz0JCFTXsnu+lrZ477E37mY7st2nxAev24LUn7rdwI0Lr4wJSQOJOfzRTKivSTRS8ixs
CMXJ6HLOldUE1Qfncga9S6nX9BlWtyL5k/h1ucLkrGDvVYTWdAxXzerhgx83ow4U5d/YlSIwrh3i
oCAb9/UxUrrHmhPGK08PCcO5bH6B9ZBqe5/wcLtJ+Na6AyvGHrTRXD1voL5mtcaZ2mk6+rTZea98
1Kg+EHPgS5Ag/Fx7ntePvy+HLobI21Pv0BF/xtfbd6JvOurlV7sa9uxNqIVMem+fB7Eo1wLEh0dy
GyAgk+CMelBBrcIv2VXMq/sfNLPk+AcU0a2GyNbw+H73+eNf5dTFynY2yh1PktRM9BhCE+IOSSCN
68zt7BIKPYQUj+9pO+d+726DfON34NlkZb4IjZXKBu80fqne1YLDADxRrutLHrXI47PrHdHIB/DP
11wiQXFfLdQpogQnerY9zsRXYEuU5gAgQbaHy9GJWXhLHW1NKbh0kasMZGAempET7oFQqEU+vFsI
1v2Npi3ZiKgaamCbPrcpdORl0zaOurWHC/+zeFXD//eJzNojnwnDf2mWUknx1YmCh0mOi5u5lmy0
LDdswqtopWQ2rVxTOmjp6JQ5h66MaRPzBHta2+adngoOFjXihgMerhbghD3oJfMm41YJ376xeP26
c/gf/mgLEP4/IFuWVMWxMPcQPBB80EslHwA0H7acWPuKM6wH6K4O/HhyG05VLYdfe2caLprl9mTx
lwgieVhWwHeYhyxFTpoUyK3+w5ch2d8Nes5ZmdLUXDg3OceY53o5a26OO2NyBsoeCVcyBDzgbXCm
AYMauR9expe91SUV/3GRIYoit8+M6+Q3zh04Glddm7P+aJ4Xjsou2AJfxQ9Eey8t1hycxZXmKA84
1VbD2k/+ORCsY0obhEm3EDKO+8JVu8gXsLFcYEb0/V9XASbOFVVJFcc1lX8SjJnnqT4ADCq1PCK5
0AHedD0qSfC2IR9B9nFMU5jSb3G6M3SRqOmPrYrVC7CmF2LbLpPoHlCVY/GugxDix4KCgLcZzmLN
6CJChMF8oYcyHTRv+/FF47h1gorZ07GYGGHYkui72rrSw6Z1Tvb2XqpWC61sJq0t9QlH8F/gcdTp
llQ0DyhB9qbbCQYGYWbJ/qAqLZguYXNDG6ayvlOhS2ph1FdIwcnH3tv0qUPee2PjlhyBRCNA8Onk
o7yKm6TLNu+Ze73siimyvsFQENZRbPoSGwtaFJNKLexBLOBaE1uvSBD5Y/ViayhSVpm+0fgeGkJU
l2x8dw2zqnleDFbcUqaanxErqlaHHc3b4Q9z1laKnXhZa8I86ltTtIz7qQjXeBC6QT6edJaHuitK
PuHejeA+IFl6bUie5DrLDryBhpRrtXH1NQfXHhblEo5/X2o8Cij2/y73211E9KSl2ptBwXZ/oFRd
b8MOUv7alht3qImUm3JUf3oxA38sO9v34AXhaj67J90wzvB5ZG+RC53jGaZw0JrY/NW7iL4soPnV
m2tKv2m/o5SYfU5xQ+L8oa0csZKeu9OtUOshht45USgl9js1rteI37ZViWf111B3Gf5hBR0PDCtT
+gKtX7f0v7U7xd+TLjx8qdnEDDu6XBBDuFXhh+FmYwxAPT1ibf7UcFhhBKGdpIufTQMMnwtAwltE
5dBHlm7Ias3aimLwl+yvRGcGI0DRV/J39cRxj716YXIWqpEInUQYwII8M7eJlgoETIGK49GOZebO
5oqFNIjYvickh2iRiR4ZBmrxoGzql458xhCaz/SYb8pfWJU2JTN0AgZxV4Y14SaVzTvchZQJiPL1
1hunh8WaSiynGPvv1H13Tro1LU06xW7gzFamUjS0byQ0s0fjjik8+f8URhNxcj0+qR0cY1/y2WW3
0Y/brqyjtF7FMj/9gkoiSoefyRjanvdB2hc66tl8kJ/OOIFoLcR43H+XGh7cQ/Xlz7O0cg6oas0b
0dTUlRKIzKb7ebDn72tUGAZK8ZO6KH8X7u6Vx9Vp2zyAXmztC0lC7GG0oh+RSZTRex0EkdSW0DeE
5hJSL3gnEq8lG/ilU3e2AEqZqItWxRppcTsG8WMOjnGjXyMbxxHJxFH4vuVG1IdswuDlruNmFx9Z
eL2GL1TO7wzFVMsrnb0ZZ2ON8BNPyKnPInt8tOWkcl4eB16iH81jmDVQhFVHIBvL2wQQKV/Z/6+A
cbgmvc3qIxtmTVCwGGNDBcPuEPtqU7dKNGavqYacEhXlmoalaJOJQX7ichXJAfcJ83tQg0VjYZfp
Z4rFfF9zt90O/0JKPi7UxiUAV/eVbaD1J9//LxvMO4Pn2hPLSK3CCTGhbiYB0zHUjTOjC/BbhR79
BZhzBQ8rI7/68CyyO/sYfvjG1JSHhdlBTwHlNtemDBynMD921k4/8kMy1Dcg99Dh1os1dlwUcPBv
PouUKKqnZM0ulANhxIQy8b4rg2e2+8qCWypDThjmza4eI8AGTL2arMsIwN73qhP+Zy99KJSAm6C8
CkQKyhu76H4d61JsikZswKUtWGP3PfJtb/ik8xASqtebNMFF5syr5WxsKR/HmSNUsI22rxzUpOiH
XFEf46sfRNsaLFY/FR7DRYEUQEOg7OrUNLoucehNlD5+u+Wpo5FAA99mTH9n60umA5FIzPy98j+n
31XAQRfBIng1TM7yG19J4GnNSp0VIoIUzB7YzyDf+UXz4aKqFuslBYAB1eSMBrvv0uQs70R0gm+P
RjuZRIZwUnW0SVUPSbnVOrcWrx+861eptnkg7+i5EGIWErsVX8oeGZiC8JgGHVKRGOQM/b2DjBCE
avyj3ybMGU0AQ6LPnlpewteabbhfcuVhdZhBIzOCi7hLzZW4gTEN90eX+HiBy3G2CryQC4w6zvjc
ol5Ndmev4sAZqKP6bBTsi6vGSHIcHo1Wp1N7pnoo3p9m+fXiSRlTzItxZUtv5pGsU6l2uhPveZLz
z5y9qN22Ydrbs5AnA0WBBbsnTejRV5ufKQlNq4KOVsPTI0iVXqZopJPHVDPqp73cNawfYTzMsTVD
YLUEWYFvZOqBOsU3jCvBELPOAzPzskOlt6u9ft8aLatVip1Q5Nu7dFIQwVuGTo/QtiNZFCZiSGzz
eLLWUsO92hPL5RmrOo84W07C2JdoF8MQnBTwDZfVvNpR+un54f7mdixp8tJysHGZuR+l7CrX2aH1
Bo3Bwg1f7W8lSj+aAN5sQGn1vKUBzDjVDl0Zeb6CJabp1q6mHdpSHA3Z4oSvZUW8br264G03VoFs
+sPD6pVk6yJfxctikIVbtIetqH3Y1W6pzGxKd1LEfRHDISyNcbLpPPjJrW+EGWsYaWoRCbxckfTB
6utH110QfCu3J0OhCa/sUNh8CLmD4fimWJc+WuklEnZnx73RqQ2dW0gAPm/6/4DtSIj5SqYg3i3A
g6D8Y3Y2tlo9uVUXeANL7FAXF0NW+2jELzisvo2pY0U3tuXbDgH1Ql0PHwyOZ9edt7CoIBHOJ8vJ
ZoREjFSAfDji5nJzQuo7HgKEcxsCg0ZrtCpG96H+Df7+AhOUGB8/9RvBnVo74xCFJTkKqMNN3znv
obGWnA6UPTzfj8/JaOcWMu68FgUqOBIZzHzoerk55y3zCQSOtBOp+wmJTfcXl8xAKhjcySY7sikR
fRbxH+5SYJmXHXc2gnin7rH9d7oIkaKiKGzREfYaPZcAloS0e78DLjmGvc3mchiX3zjzWE7QpmuW
7tjQhehKd0PFdI51k++Pj7qrO8NOoATU7iV5qZp7qxm9XpV9ii/6+4V3nBxEvqXTBe0YTxFBc/2w
jgdREN1wimMtFW0XnQlk1iZf+PcUciDdo3GfGiRkco1EFTSriaADCBv2UthMdLWFar6zjiuLLCIU
EA7IDzAOvm7XypnacQx2Cv+YMUUAtGpeT4zBzEsLGt4jC0FD8g3e1IG+tmqxMmvZDCytOAoL8DGB
5qjrBSPvy9s+TtpvHDP1FkNHMfbhFo7xFBW8G6FOYxZFJ0zj6rDaFI5Bih0atDikc/WaZ3zJDFRj
Uv3dn/DJGEUkL15No5TiscABFol+10WkFUJ9W/bgBkHdXRS8qMQ6n/x3XPZkqxDqt3Z1wV8tBgYg
XkrZ+hqp07Pk4ZO0AbumNmQRc036Yj/iC6CAWrUwETs/4Z0UqeuI5XXAu9eZqYT6G0tGtKZW2ME6
kQM18KhpJUPObv5ppXjRMzHL0kA+1nneC8/fqcCktS3O2r05lywavZhF3t9tFJVl5a8pQDIGnWcO
ojhX7wjnhmzvaBb7bnVbpjJl4ld0bRlv8cYTVWrYJDyx4eJKO8Wl+670rt46U7V1jQzBoznOpjjO
ol7nVc52ojIMlMT958h7ImrZqy5Plv7NxUuXty484/mSLLO+byp4zPTEEt1L7FBoeO2Qx413tyrC
qdYBM3S8yQ79UeM7U6DmwyjxFSSc34fUq++nvNhqmM5NaT+OQXiBShNIOVqg7v9ToMIuBPDFJ3UA
fBNko8gnv4uLe+hiDn+TUxMVKeDF+tGUef+8PthabaarUBzfskU8o+xr6OUBVSlGKBJiBjUGhO4o
uQfnCerpkT7SArTV1plt3LhKvLEcWC04i4vvH6v35KR40GakfacylG79ioUFGvIyNSoOz/x8Iw3f
ur91mH5hgHVVfXusmKgpbnKu96m8hrIODroCLywLlGloLYTvyPsmDYWQzf3or+iyFIFppy+o0G0f
qkp79+6mVbUFfgighS+UQY5d4MVzvouTILtc+GCzagSM7PJp8tvTe+dAWpkgcxTA5ylGPuzYBEQU
82g5sFGcPGeQf6wACfMy2PE+BdDOasiI5HyCG6FzKA26Wxdf5xVg1LBvyFSSMyAZk81eJ85UQBAh
uys5co83lLHZOxDMy5m7KWnXf7erp06DVOQcYjeMx44XzxsyTb8+gsAmhi4BeX5r99a/I9sEdv3y
qNbmXpK2qAJIMYF5iSn+oAWKHWpUYuw5xYA8oniHsHi0UcPczd3TQAxTgEMaF4fs9UpwJKmHAzr2
Xpz5hY8EQnWKb64tGTrcvQPT3OlMRzvox9Hel0xXYy0LfSGPuZvPsazpsbCPwR4e0KZCpaZ9w87x
KZcxKqxJM96FRibUpjv2LD+fLs4JZ/zvMttWneDUumH0Vy8VF5cd5S93Hvzv/3q4DUxLIwSQjasG
/7xVr1xIpf0NWfG2f5YLfjyfbo6Iggs3yN/gUSMXJOlzYUlLGNbm/+M8I9Vd8oMIqeQvMClVsK80
QTzjFSI2xBc0XQ8kRyJd6gp+JCPiarK+8pp9yhYD29qIERLvaoPYe6a2C9W11HwM5+4FGBvjlwws
aTGIfs4b0OtuqQzBWezrqdIWyAwnxX2NMn49yYLr7KE6hNvb28U4L6yxtgwNGbkZj65ffXjNKnXd
K0wFHqJ1y6xKwqsp8HqmWsk9ZSKZbyTSLRZRgBIoEsRsUGLOlFceq0+RKU5YFTlSx3BBT4EeSDWA
t3XCnHSYS/sliH6U4T4zuVbN+lNoFeIDuzkcZ0lDtdgxsnbhlMeOJie+QTbfiWdnVn4d+xhAHI4q
M06kqFAIa0/UImW3er/zMXTMnzAfuw7hOQUza9FjyUGXBvaeT/W+EmLWEeAh3dFVT3YMDZxElEC4
PselPygEwOOD7+FVTAgXNKIBpJg6LO214PJpJqlf4dz7v0o2SAMDcCc8D6rOXgTwZHpgim6oUNus
2EBYtwgcCSfxpHpT4kBqNYgI2U7KMKYwDHEICAlzhjyIm1ILNG+3k+uJclZrD/EATxi+BMlRzQgs
h5cWDEMw7Cj5NlkrvSVb25WS36anRHYT56lrPw17weSLUZ5C4xCUFmKXM5VO1/0A++ub9vFVqnFO
NmVOADmArApzpxpsDdZE4050SfDp0Q3xBtnJwDk/0Cvdxo7mMLzwkEgIZhSjhc6amghiAmHXvCjm
9tmcwQE2YHMPL5qGJMlVNaZSBoCyBCNs+fvaZR0yqlnoQ3ck7iI7e0hcBGtt9FNzQQgTouYaTqNc
3QqBiZm8m/Bo3uO1QTiqBSemCvhZ0oDBpl3YTTGAmkdCtKFZYXHMTxHEb3RY0G6JrwOPCXqfdYtO
+FLtencCD37VCgEhoIbEtchDqwNVfhvBGxUF+hjyBfI08zov/0wzAt8EFAVO0PaO7h2lTEmS+JyM
81Mhftr/soT4k69RPGA8TAASTnuTtcM3F4JF38u4lL3Sr3QQy97BeDF+xEiQyYnEAbmlJF0YgXFk
vi0iXj1hBxpL5A4CxOTALbo2y+GkJ7ilrHhUgIej1Vtn37VDeIcGeSeR5n1tj5H91uWzH0gLA7xh
hWt6GgVI3JViO1Q8Is1fWJ7WB+bhIZEAcMxZRBN5tZcGvebDhu+1mGDPhyTO4bMokuuuf2Q1NH5A
vmAyy1nif5lYzGLzP0Us9jkBJ+AAxuEyOWSni28QSq+U03ylLQ6SfGPI1CBA/8VXHiXNC1lbFCj2
caH9ui2W2bsQJKTHTEGzPCiphKQUSzEcGhr6UycqKkgyZ+Owg7Z+VANa/xHHzzgJT0Uj7AUG2YRy
G9eRLJmdVShwU4yZciTvL7mkHCaGBLuG3CygutnO3DpzGN2GGDZoNMktuh8z41Gxt4wFzWSd64zT
w2Lt2HOoACAdKnW4H4A9ssZP7djM1sDIA895k86ys1vnd8WSaT9s3x9pbLtLk9CPVgfE/BOyueqL
hmgM3InF7LP37LrF0LHmYnJIMLsKa9pV0dnjaEJ1nual6kl58OTWOwaEjV7pTWtEQnVct708O8xH
2v4nLqppn9pD2pWGbaK/C019nKstCub4oSF/fZEx2FgX/tIMeQ3RK7duxVkxZ07/TQTy7UP480Ep
XXwOTIg2Jj3Dl1wIquoPyYoqmr72T+2NWdqe9GKTSSyvv2WQHQVjNm6gfM0sLHAFC0+mfbA7Ca5s
Y476ajEr/2Zy54iByz5ys9fDlETrxwHV/tY+7iaKzbxbyeDrr7o2/hTzKwaYkh2lb/qXBPGUfE/4
Kwmwe01uRK2PtaDxXxEKlbwBDaC37HkKrAQ5j1wvZSXQHvID9rXrzZ4d+q//yInCQjXk+pVvO+4Y
+Ic6cFZUATUipUMXpzZo8Sy+5wSuYo68TeE2HTwEHI161rDUKFrrbpORNKO8B3EIH6LOQ6xuCHra
lV4I4YZesIrw/AvtD24spTQbwDGNrAGm0F5ppqdc/LUOQ+O5kwL8BcEjN01plYqge2dLgkbrcDnz
HNjVKH4agKyPEqP22/I5fYycTvbZuEHrzo9fVpFxeY29SS8ug3OCj+q7GfJTBioHejup/bPDs5XM
49aV6IvRGt+BWSFeoBpOVJ8Wuguz0YTWZZZblVcKF9Gv/nMRcuLsADZZtH3+q6mG4ttAg2HvUFMS
Nfm8XDLLEFrJugQpc6YNAUdyanLKhnL0mWMLj4RTalurZttuHKugMs4oJGZOa3TIQVo/12icQGUn
2tdzO4p+wJD5sz2cS4aizjQcqyztJxJ30fAXLP6HPklDig94NOXzxAINRh4B8j3GW6RWjRlWIKIK
nW1/T7snRY/NMbpTjL/eAm6jmTBM0+dyw131Mb9cCb+Zs5Qy26LKERHtavNVuG2jg23l98Ht5FCN
vZkbikNAVNI6gleqSMgASKwPkA4SYRos4apwQ7AvY2XCEm5cyOKiV1A9m/QVaPiqD7Qx/iM+ilcU
/8hYelJH57gs+4Zrf3m9euZRf3DVhwFALbfIJklxsan1DbTxFEvMoCWtvWlWPKGMlbVnSAtgWwJC
kn27BA8pehqTJEgAfZxt74PuEqdztLDCWt+sqkl+arFAvhsfRYaFNPPYtzsDN6y7EqyI5+ZYwAjc
foIXCj6xP5Rthxi9ctRCbC+2Rk6btmz8W/fhZo1jFdWb3Z8E0MkKvHS6voIECtYnb2M500WJ0OKR
XLF+sTZLEIERhyDMlDsdFlGL3fGdAZ0pSBllNGgKwYWSMcPGb2jJExLaMgGbOJJ2/syiOJFvVeJG
YtUK10uEt9R6M3OGTUggfNRD5Ck7CNMG/kbLQLTg5njCZeKXhh5spAUcDC+q2dvG/7J7eyZ7Q+ud
GsUC307kphckrbKRio5qYRozflPDY0Wws68/Ws7MAwYowcdNMeDDCUMEUy3Ty+h5SDZCDVsgSp00
npkyUmnprOD/E4JWEp3Pv8/0XzXNSFdIkBmv/fpvMl2ySGw7+UkTanatxlljwv1u+QqgdwHgRWBh
afxUnGH1Jrr5UTSSVGV5ArqCHy9xmwJFw08rM7HFPm6WorNmtrqqxRW8ktwhXhS2QcOhxF9zR6Q6
4XCuRTjaEolsPd5oIpoEinD1Dq6PxtBVyIedOlmk0NSF6+khqDMShX+s/ZTNP5S0S0Gq3B05gmxZ
+otiAD8CN44/LiwjoWQJSAS8qFa3Rff900eqfoPZ82o5ZKBP2SvuP1hZB3YpyFm3Hu0UAVmrvTqB
8IHIWd3SRPeKfuKq7lyy0yeKSDrCsdoAa17f5ioXZylovqjCT8RbVGdbva2LyIEopFdMzjJyJUqh
5Vl5cqOwU3vgRrICfLlPiJvlljBua9ZArfPL+0bodDB90PUXI4fgGgDZu+9fEZeklwpRYzpjKart
2xWx3mUZev3RdVsEQeuct3QtiD+wNFDmPBNyh6hJSvMxvxyCSbJhI3UCJcYb3V7xCEJ7isKWN4jC
5avmDYbGlGMEBvBJ3EejzaZSc5jMVMZl6AYxu0HxX49at1PTKcG1CnIZoBjlUtK5E3rFI1NJEOZH
/2YGnGcjda26IgTwdKm7OorwNjakusD984onWzaO6I0umEwb09j8rVZU/t8AiCItz+WpwiKigQBg
LUZIjKqN+Bl+VW1LHj75xUNnb9YenoJBqRL25ClBx81FkmmTlKoFd3bzKOQhuQ1qnflJIUaLB7Lz
qRjrrW+Vg+QfzsKauMNnao5rBtQgW7kW06X+tDjqA0pqTjwI29po7ExYvFO645MVmGTKcFQHmM24
zrBOzyPDJ3Jld8tulfTfxT1kNmy66GI3tuGcv+V3ylMi4VHLif6uH4rJDc2hcXlIOCvV1+n9bdr3
vyhl2yxWGRyJKv+ngjc+pPH45HSnMqtp7DKALNG6iVgC4whW9JYgd+7d5Vr//OkSfXP6Sz/Y+JXA
0/e1n+JdBf1B9SKkPDW64RU2dKSw70vithPDzrx9bwijit9DvJDuuRA113DOrQ9HTsoRGmQgBHun
cKv/Ju3dxn6p5KaESReyFZjcuG4C4rdl77J2cW9UlUZxLS3w83feMgi0qf0V50WdfOUVtu7GmNEJ
hFGS+Lc73pv6jHdZdl7w2PtnOP9C8IhUgfSRPeQpJZH0XkdiEm6egNm1B70uQCsFDbl1rb8RBJlY
hUCJuB2ti7XUrT/Ozn/C43QF3f4t59yif+69hfkW7fkJ6nNsVMysoRQcaxgpzGHOB0ahwFa2VGqC
trUyFez+IjxurgltDxNIZ6olugOWEiDWcBzGyzLkTUfcxxD6CkV4Yy02Sb3lhP4XWPm7sQ6CmLCj
jw5HvsetZ8QR7tua8v+jvd7vM4pTMLv6DmWindzlMBXsiWBiP1betD4Tkf/9dow/QNezitIP5n6N
cEX3tVK7oSYwnCziop34vXEFm7kJQqEunv+Y7+77DrkqNrODxq4m/SE8dgtYiHwzvuaTEN9SIDHC
PQR6cG1ANE2vkHZ7rqqaT+COIDIlbEfolu//M2mOXo8oYPvyHULqKgYhw4zLJKJrTTlKezEwA5vy
LX7/pajI1Mhh0o54hM4waUefo5eC8rn5dKd2CouEPM82x3n5Eccm57hueCOkRsoYdkRJM8t5LNcU
O/1k2n9hDAKxJ3c2LcZ8PzXZkcMMgazSZGMBEeJloSfsTthHjjXjWC3H9j3DbFFN2rKFfdG3VwME
p8xxo+AZB2j2wBHbH8B1RyvHpxJMaMJkL1dA5j+Ag4yFCid0zmy0+9YKD2qTxwh3jZm03RLwZU62
YkBrc2aCVsbd+E1xy6g8Ft2MmqnO6RX4Mypg1NGWzPEs2HqRDf5DKinm/cLsV9/kWXEeTc8I3EDL
OBFluVvr4Nl0tQ1HHhvHYXN48/BCJZMwaKU2OvLZjDjoAsvDFPNFaU5Oo+/Dx670ZI+cf0cb27fF
GapcLbLnog7J3tpL06CNTIhXjTjWjfGSTuSYXTpJpPLC8tmUa5rb4YeezazsArVd8Cd6Or2jfaeI
Sz9MuBcu2/RVAU+YeOMbNIyT5Pt3jTCXuNRyP4lHExicX4th1UGqq0YN6Y57oYgDB7F3vNOLIM+P
dWacXj69vYkenHinlalM8htIauyOACEjOX6uv3hwzFRwP+ummTXv3zPkbhf0KcKrqy75feAtsc9E
DrBkArJJCq9GNkPt+pzULNPfnJpMiqO/rWEKiVKPggdUtUP+edpMsymYoql+7VqUevFW5AeUA6K9
iyDN5HQ06eXQkV9PIrrAKXbZzJpxeNVXHQdMams/8Gzch8V1z5uUxm1vH5otf4ryatf2WOwNRnRG
DmDoMqFK2YHK3NmdQwSAvbZEuMOTQwsSY0bCAdpvlOGb0XiKAjciO4DP5Cy8grAEY+ofl1e89JpM
i2NCQPupYX1U7rMs8KuWKz0LRpsO1a7sFD2sXIv8VwAXnXWCzvh+GIQTxFkiepe903dvgnXzDFfr
pkF/Wm2ap17sWrK3daluHIuSL7c/iCGyV6UQFtI1UEwKnDexZY2h0/GwvMS6H0lZY89p90hw3+uj
Ey0i5xaSVDx6IQ6BcSwDY2yZ/87VHGDqhzQh+S2NLHCkIe5ybLqXC3PraWb4GihQX8gZxrWAk5BG
Hk5lXns2HmM53ka5iKQYNu/WUP/CflEE7vx/KH8rmPdnnPwN6q/DSCebl0PUPnTGRq14Fxy+Snbm
8ggrvJIHRVGQOJJJ/kfkrJLLTMRB4PUgYjWyXssiMl9j4ZmZ4PbuX8XrujuJn+1b7/QIB6pWBVsg
/vYBd3ySzs2AfvrMv4HuGvnMgpaFwzwrHQzWjuUgt9ze43gRBqlthIPabEoekdT4IFqOMY9lQjZR
c+Q1TZ5FmEuzGzAOEInTFXYnfaEHILJu47kHBKBO6S+9zBQ06M8wrDsEOijrxrFuzA86yyoIDGmn
hccAeDNEH7PL35dOGM4wY/wQa6mVLpZQOH2V7vdIbZD5Jzlk5l7S04e/8Zs5ABxIK1mumrxjjMgq
E9Qe4SQ96rDBdhY97k0q6D1GkDw/zGIr7IZoNWSrxU+cRekT4xaAxkNxys06l68LWy/vq6ZpBofg
ejwPIgOt0/xCGZ9tt6VnUTgU816BtEuxiB+nW0XWFDsg5HcIZ4WfPth1hIJ5foGaQwB2bs3HiPrd
jzj5Ty16vRjzSO/NWtTVvdRDAff1i0V8wpKEgyGJZoqpf5hQDesNUEoxiTXRO1Nc7Ecnqtond2+9
+StcSPArPbOgYctVltaAsKQFEVYicGcGB+SKXVli8aUdlWqdMAWMRywc+zU3evH6k0sh3CD7HySB
G0gHhYucChazqsilJfxhy1hrYJVK+R1IuPzzlPUgQtxFcWi8JHtQZ4G0pTnda6EPVKEpMyz96p/Y
rwQDG8O0eI5ZQm5yqrFtJofuE0c79VOKVrO22eWRmPpa+HmB/mVIg7sR81Ie0084rZLWSQklqal2
Rj6aJEjQ6ONg1Z390hRGIpXlQ66ceWYOowH9XHFitgqZ20zwEX1QKcMwK4NXZmaMP6mkjV0EJKLt
cMCdcKAAe8pVKxsSjpGXj42NgX/AcoZzVUnA3FEd9EobUmaaKlaEfPVXABD4j+2Yx7I0Kx3zIs99
6q7KrOjYS63NdPBY12bIJkyja/A+UmFEOkJA1V6jedXubOqZ+HQAUPABLAkMAbQf/D9Ambl0U1Nu
b63AmxeztssGmdhKOIQ4vKwwh0ziWfLs7IiN4/ua/e3Tfs2k4+KaWUopTKxsh07a6f+wfev2hoaX
keKj9ygjal2gFkByO0YEpM+02aKMQZh+JhS2bfxdIg/FV8dMT4XLXkUJ+zSXBXSG2ZU6Gbi7I98r
5Az53XKUDWOGeLXjVWrNmzYu2ldrocNWQZVtUA59Fd9Em0tuRPnFiuwvD1Slp79peXujB3j+3Uu9
DlUL9KhKvsVPTBso5TC9C+5TSRSwtiIVarEucfYFvTXl2cSfz/xohxxPA3VMLp03QMsZMYxD92U/
yDO+FzT/vwEl/mN7neL37b2DlP+u+VFOx7QDWkNOHixwQO0spnfDQmXTXtZxFT96USWkdZh7WGoB
Nzsb0pqbKRWxXtCbUEtrbxnc7bLZRfYzkgNocY/QC7hpHVMMGePUfOndBX+4mL9q09pCXSaLskwU
Sr49/MoBxwpMNs5XAyTRd5bPNNSvsSTjL754zO+bm3ZA+8pK3XiELGXWsgKH+MuppElMkniEWcd9
X4cX3IGysQqdDAaaWX0saStrdgHhA/Y91Q3mGxqOJie63ckW9I8lNHeSdnlsDOKGpTxZhGB0M6qf
/n+ef+6xuG2bwpOepjP7pC0h+Ti9WHGgz4UjHGOr596NajhBOUlpW2b+RzzxUkbxDfwqefsIVWZ/
dmgIP62cp7/XkXjmQWpLzmap3h+hOnlNIJIMQS0B+4eeOMqI8/ZMDTBXPuIq8QGpPb4hpRToYB3b
yALR5qabinLHWmxeNA8nY0m6hBiWq4f+/w5e8X8AFLNgZyoefib8jipKhFqzPUhAyJdbzBtpWlcz
av+5vdyd1rmZ4AVVjsKxD+XDL7HDQEbqqEfMbM8a/xVTsQQQxqM6TpEfOvHl0QXfMPNX34t0IWFW
M710L0YbKJZ0YHHT9Xklx9bxkEa2SsXIajqW+8f/8aMeaFGc0ltCBAl/pIJoPf4yKRxRR+Wy4oyS
brnLsQZZE+lRewHfNx8CKG4uRwURVVxUXZmVh1glH1thirgfxChlAS8f8W+S6wO2e8ZIzKJXYLvK
0ZN9moSBm26FsMklBvE95WwtYrTMzrBcXWIJx//RaPP+ADw/1m6eu8vwX4rh7h2Ub5He3+iuE7Bh
ffXSsEyR+vVcbYS+dlZPBJKfNChNt1UuHbtI8+jRvQNuWIUCanrjIXZeM6HZ2RB68TO0O6VGNP6M
GLtiS5gQ+XK3xBSaU8L+SC2CKIx5cN0TRJoQwjP5qUf0PypTZXYL5ZPmG2BfQ9x6cNBKWmW1b8Ua
aZe6gH+D04lh1FR2BgTFqbimoIhyfGrBRGkgxk/O/TwGyiiY9+71/7vvsZ84oxfBtyqhr7pEss6O
dx/Eax9agDiRKgiMocAn9XXQzgpmMxOnrNTKx5pEoDPJw+08w9We0FHPo2jPXHHmX9fCeaEM1O0q
cPM6dJnXtrMoXuR4WDfyq/76xMR5cENyR/npOkANaWjDcqhZYRdPSReHK2dTAR/oFP6rv91wFYAN
Bn2mKweC6+XhbAuhPz5hZGU6OwXtJKHVyamwDchEcaw20/c3V+AFWjy44bqjdNB7i8JEyIix/lOA
9nCqupF7dpppC1uVrK69+/HTUJYl8arLGBE9J+/TyKqdZsJmcNHIsrkKiMymEbBRKi5y7ks7uS3I
bSIoyS/U/r2t67qk55JtoVZ8oMvJ3JjsXecdHbH/TbfQL43/zl5r0FAo5abg068zisaHQMt3lbuT
0vy6A8J0NxxCef8LAzmIgJbdB8g1/JAgt6Y+Eba8OU1bqsiHGofn66Qqq3GJNs5TfTb+1Ps+n8Cc
TaZ2uT86uj+KnPN85v/b+fa3us6d/K/E9BCfmiZ4y6Iif3s1LSp//nq0zN1Gaz+GN120+uEo0ski
eS2BbS+O1bbBxSDnA96ppciphZXf8ChyK9Af/Z9dIigwSwX9yIqpx7QI52Z6II1GZgd7uP5Ni8sb
1zTUH3kytdwDU6bGgXq2r5o+SJVavfiEaYL8qs69ojpjBcGlKkUTdnmNEdV7bVYCyKSzlPjB5RMR
pD7/4i7/JnW5Yyn2UtBKMm428Ll17H9clUXayJgYi9icsG9vsXLMDpLyhak/itNBfRkzgA5sS2Mg
t1slc63UZH/iyJTQGpHkpNPL1zld8g0uRuJCiH5F5kc1opbmU6EKLn1e+VMKc1+6Xq6LPQaUhrvk
6VkOW/2ISQ1U1udmxfkyXh0kqVcvb1b8DwoF23wXKyU32M3o49l3b3ph0pQzE+y6d9xkbKt9gENo
hsLQxweWSNtPbJJq+poWtOqP44/2UMeIVYXIYydT4hxppavOuah81vWcUQ+px6nkd2y5l6d5edb9
l6NN1hLHMVFG702FEmGBNy6rtZcZ/0zMF8zEZmYo+tBE3QRuSwbJaatqU0yj3JqlBro5BjFIqwuG
T4ALlA+jA7n7R9My6H1H79DzkLrTGYnBD2FeuZyPaH4VWQ3uzwbmVk1was3cabAJBfvr3OrsZITG
4D4Gn26W6YZEBgEleZA3rpihC4+6CONme1M2pfF0fgukg6Uv8sDgKvWFtEeRpYohiOcXNgtUOR1q
qyWnGdtL/J9hyZhtLsqIOHs3CSPKd7th1AQoWHojd9pcsuIHgENE7+CWW91Up0JF7O/RVgv4LVdi
5W3PFWJ6B8TxkfTzrsOD1VzRElHsf+/aMwKlozBwYe5//85K7De2t6VERCmwveMN7o/Qywlapmg6
nC8ht0ZNvJdoEaizKd1aeHfnYzeQTW74eFy+RNogT3yHwnSVUh425Wm+wGIt570wzCuzf2fARZtO
oXsWfxBUlwiaEK/wweiOVDakjBZtdmtSG+LYBJWe0lnLIwVXTD59NRmqRof+YQhKfORJEwQGbc54
4xGw7noMctaGNX3OiXTX4q9JkHBwpfVf2LcJLNoKQ4BpcOjlhw1Gnk06dZ22Keapv0Qt+R5SMtKG
Fo7M4Fa3laxsQzXu2B8U5OopT5Ry1/mna5EcP7MrhMagfsSNUhjvix1v3k9SN9yXXyQSoSIJpSDa
hUOKzUq1DLNdtvCbaT/1EaUPPVGIZyoA2C3BJUsVufUvgrBtreZK4tZByUlTkZQBWiyVsigVLZVS
onHkGuZwNaBuV2QVyA62pPBtmZhhjY+2FqjE59A1lSBQHMc1RKWVp0mMlfhfRIwUKBBsxmDqEcqd
nfbOmysaRW4GgpQIWdXMLcHTs9PxDMszkhLTr2cUKnu43sSX3ZvnBc40w6xGErVuUrFp/cpy7K3Q
iSB1RVlSJd8/yc4uxZLwkQYk++LBcWl8hkWvEYT4kLP3/wJPAkcYibm2RAF5OjMcnu1k/GG0NzEr
OOO4CHm0+CXSsz8Sxx1W0+TVANs8SqA8RxpNxClBSbKZGi07uAO/IIEufYS1Q0xVmIThJ+VJj+hx
gv/GCbRkkg5RMXGQ4oc/xfvJOzkAfgVjHCWoIADVdgzeHTFxIPbxoFujhqvx6AbbHbEet3R7H6da
WJN3IbaXpUErYWzhpBGfYI5wgZnJD25J0tAKX9jyhThi3x8fcKxhHuA2MyOFro/U69e9m9YTXxKz
N01e55G0BEFzecccCUw2/pG521T9wR3BBrBqHwh/3yyPPAbMmjQdSp9aSK3d2on6tptMQK8lQrBw
tt5XyCX7j0d9WfLxj9LJVq0axyUFvcgqofdK6DWeN9BhplWekxKHRTv5BQPCXkSJhrwXAnyR6mCz
rW+MCjx3CuF73Jc4eKV0WO/Q8IL2MYn3oVfemL3mXrEzKCnO/EOABbUEx+w4ADO6FIIlZJ1x4q12
ZFA1ylUrtyoY9R4b7G0h+9dsnuoyzYlzU6j0VzK8cu0UFcANZg3Y20SFYPZ7vFYhraD+fAPywFcp
a88vjf1IGyRePZ4r/TphjcYNam2DAf/hc2MlgE36EBPb6BKERahrRs2zk/tghbSs6p+FlJYaxqDC
Zcr23+yBlukz+QWveThPnPtaPwMW/Y/M3we9oauNWWOJIbtjlF6Nt4y3TaO/rsTaf8Y8SLxkrLpi
dOaJOPiqo9UO18ACpfzrCQNUrI2InLHIlXGD5Yu0/oW0BZy9Gvz8+8LMDbV1aeKlWBjCXeqjUczy
32Rlc97rY2JQ8mvIuWviihOnfrJVzd5NIZMVnHJlrrWQ6u2g5OXo6r1kF8YNlrGL5AOKUzeXO0gR
K2J3qo21broVsPIiyORtpUW/E3setkwHAJODNrCliuIYlAoyNodV5cSt52IoqrsKZdVeq+lU0agj
F0Ya4aYrg0TNK0cRqiI+FosVaDpAZtkZ70voQyZMmVkVTpBaQqYLC2Hp9c8qyo5aZ25UAUQZtes1
UT4YaxW3Q1+ycecxbjPU2qoDPsBXDtUy9DrZ7S3n+juxCFfAhiWy2uKl5d9NB2CtfWo5PB8OHC4q
/t+Yam/5D0C6hRzR7GLqbaHhw2kiqiUdczVjlE2FO0V4DovN5I7cY8Mu037a7xEiTkqSK04KCZX4
vgp8TrEbtMGEgD1llTv7q7hwgyJr1mrR2+6by41Na5sycwTHaKMQ7zKDmbJC1hx9pB/8McLF3HDc
YStnBCcMqyLbRqzwtZzRE/yoefUZGkf9qMz4MDKTVdK5fkEs3qOFDABC/sEVHMVjoNcpKOSN/WHh
Mgwgk6Ij2jjAeAI/vF6g6FipKLknlGLVbbubinR6IqEVZ4sqbN+PqWqo+NF2mDSBLxFAUZ7WTAyT
Nt3qcIPDxXNdf2I3KI697IT9TBH1MxNsuNk8gSXcI6ToLQevDSU8exfva9aaKU7pao+f4PETT2/2
QULL4abYhfFrH9kzTpeSqF08TcORjnEEURxtYW10SJ2ImsL+pXPfkjjliWVyLh7JyP2gzrLDtP6i
5UAinWi2tCIp2mBaQz8ykKgibtvxRMBY3ax84+VGLq2hAW0TvW3Z4zcQDlePx6rF7V0lol7A1Q1O
0ufmkCuNwQpuceyCJ3XcCSvQt47HP3VGX+bjYEuC9n7By1OCx+ozfcM4qnZzcpojekKdVerhSlEb
7V9o7XkAHZqgpFhrv9SupE1v+qOzaIzo1LRG0pXh7kT3MKjy/dhZf39eQw3xDgUeZJtZylLgi7rJ
TRVscMFncYWxW0QQoZLJusPIPq2XbNwIRJwLVAWbpErUUC8aOY7e7n7VcnIWD84pzuv+4PKYbCrt
hKiJm9LmaqDlQ2wJ2DgdhgoTdbIiLAy8tAUyRPyfCiTNiA2cG8JOpGM3b8K7cpUVrX00AOcOtQCm
b7rvS6r2RrIKYHLVQkywMG7myFWa8Gfv/HzlOEuzt9Td1/QABKTJo0GaKkWCEg2Hlu8bjoPixoD8
lL4c5gVSazu/Be1FQ8jDZdsvkGer3R5HMD3+ySYgMpYcVhXEJTQ2LrrA7bQdPy1+SejS3QdrM58+
kMu63CisIC/T0FJMK8cZLZGAfR0rs4D+grXT+1zw+n90RyBCSExYhh7P71JhErS+yVuxmXs3EvAy
R2aS5oa3wHDFG/vts9uqcHySygZUi8lf4PDjQB8fyF4sKTh59UsLsGzwcOFK4Q6/NFGUKUrF1q27
cA4WdCcrhYeX5OL3TIr4LDY37o08PH//lR+OwypKONyXwB2xN44FY1fDkjmKYEu3t+LrQsyLKEvo
Du6STWPW2540gNzrL0AQrw1DYrIS9Ogd9lRLamrsoO1HrBzgkNBx9FR5VgUjESxDMBgqQ26MCOdS
7a4k+MR1catiUaVYJ2ynNN6QsAf61SfWmyIKJwULcBIqFE0pbK8s257yE3zzTlFWfsqOMRWkauU3
DW9YJtSDDnlP6s9uAoHjM8S2cnjC5CXDzL1YyNSEY6T02LuruExXqlrjGDC13kR3ivpdolJ/6NWg
hjmpGGSBIGMoPInIPXUcBNNZONbcD8jQFUMLhnf0hXO/HFcSPWmdtRS4ZU1bkV4qKz+ckmRZLUVe
V9bYBCulk+ceN9uNdT8FdT7QgZbBVXaHkx+UuxWlwq09wyDBucVXEaFvVVta4sfEeaTFgUzS8Ld7
dmXPGMYIkJmZgJDbrgb66ctt7p1nOysk7nl3Kmm/eJ43JP3bIRyV0pboSFSQREGZtmIgdiNQSbqf
G1o/TaebSaXIQ/QlSGap7LEnAfbPFbPJ1sPUfuMZI6sQXFgt8icml4M5RwZEVrQJ1RonDdZsCinq
3OU5hRWZoemyzIL1k0RFYpsq6wXEkz5k9x9SkNny5NOLofxLUKoK8p5gszQ/FHmavldqGDiF/CYc
+XLGCJQyO84dHL4iIMMtCqynN6Hdx/FBl3S2CuFaYL7yKqxMEeQTnHQY5JEjZU1NMDPDNy4lQeXu
WapJj9bgX5YhNnr+TQCidcEBsAkLLVpmvqyMG/aShw2ko/n6PvystAdprIpwrZluiuTsCEJNUMlG
NnFjuVHYnl4ZNBgasd9LQ4fkPBZgyNb3tvqF6UXebUdnMnjtIX3yfu1szrbOhHeAZoYM8on36Oi4
7Pjum8RvOlPTkk34TJ4cjBYHHimGhh/YVlxfdsNa/2yh9cf4PbvkJwu5oXXMUv9RgoUeenrqIYAV
/U0VPyQFbLsK/8Nr8Oyt4mJ2U6Cy+cd6T4fSB1PeMxjnhM+mV6y/pdmpwbR8Mjyg0B1Si15KNhbs
mzwB4kvWhuRWEtUDW2hWSOINfreNRKsi07tImSZ4mpsbCPVBgImA+UsgMdm2nWU3gHbelIpe/kiN
1XY3BpW1LhI/u0lNnVH3XtLOq7fuYMfqbJ/8wJvV3Ptk5KPf29ITtI6Dh5t4HGQq9GEWCH3c8p8w
WWZVi2ONdIqN+EqWvzrFTwbQvoZ2vISPIlOP31V3UKQOkwMrHMVBiByu9DgubfrxcdS4JrJMjibg
V0nL0ZX6M9U85wmG1kVGPEVEwbY5QWJaqLJZnHeQ0+OZEhyVSEQt70QErKbCEuryklRHjRcYuC8j
FM7QrtBl+qcbF0Q/EX/EEgamp3LGNzH4/+c/E+WqtaQ1pZ4f25cz8QZCATRvimKEiAyYcEMNkc3w
Aeo5mW+i0LMLqQ4rUWkFKwQwxFYG81H7gLCoi8Y7xd/dJUPlm3kyP2B5DSGLunNG9d4eWrmC4toP
C9eHyVRxrXXtGoE7J1I3WVd9oJFay8LU30aNk7wO8Oe4HB9onQYfAtCTsZmpMYNEypzOYfEkFWPP
30Xgs2jmZy6f8XYnDEcJqATq+RC361WyIc58XNxmNlHxOHIFZ1r5Z1b0CfDCELl4tuB3CqCd67tx
6MZR/WBa4euKT2WI57mrxXB7OoKMs7WZlC27xfB0/T97kZORORwIZg1ieY+Zfs/T9IyVt6P2Kf6k
1tSCpIbGY53EdwozFsWDX+KLMSjTI/RZWxrJ7CVU56nwbcxVE2NaxP9nvej5HVuW7HKkJBk2hS8E
+HnyjeTH+t4AJaee0FmP74uUtPCtf0wDS6qSLc6NrUs02KcNgVNEU1XpOogltzmgy3vtceLlCjK5
+Sd+qATikFTut80qnKQMhWSc7UlVNmR9tT57ksQBndNF9XPDDBDopRZpVygngQgTFSv1Y4Ia16Sf
GRAiIGm6MzmjJZIt6u+gzEN3QRl85qxHRW6+Yk2MAW7cfCX0Cvixn7/9na+m1DArhXpddubdQMuU
nMf015pKycm+2Hp9jWVbsgMUuFf2nhI9QScN+Z77l+jyeePnGROnGPMRhxmEoT2FYdAXOja1/dsl
LvO+nM3EVsqrAQJ2lC839SsGSK5Ssrr/4z75r1wGejC4zbEUup+LPpgiTrCENBZHeYCz8EwU3zjC
S6lMZxJEDogdAQFyfbPiMNwlr8pht9WmZXv4JGNuHVVqX1NlETS5UveQ3EYT2nXA4Pk3AGpkOTXb
VgpMnLjnb2lxdBfbYc/MLfqtJ0pDUlsddzZbhe7Vx+ZbbHn/5hIsCJVwxd5DxvKQ3rdCnYzaWl30
BIAiEKwJy9g2QZgiCaW8zdWnlYRQzU7I1Q7qhT8z6RbKvVXQasUGDvufc7y8dk7ski85YFdm050V
gXjLnmP3IwrLGl55W4TrMInat4fbh5pwL8vNrhMsna7HmCV0xdYO0G6+Ypb8bKRR72mPkuk+YcgY
Q8kOs+g23pmES6XuL1baf8+hrGwtb308+5LovMonhKRuWcq03DYBoAV8gO+TTPvXiR7NRqRkXyUV
xr6S3TLCWkgajitF8neY3LHwgNiR3/wZ9M0OSafLZjKnjG8+xoI/WFVA0+24dhi467h89foMtre8
6bgfXvO4IizE5D5IhXXGNENQYvduBva4BOs13vv5fPax2UcdYjqp1iKzDC4tLIlLCnn84QBcLyBE
KOOjdK5BtGheaVSBUWdBm87s63jc6qhofij90j9coxOk4uetGkZHnW2ovJNgkTBu0OC7e4iTwJiF
jHVHsiamTxwpaVePQU3MJq2uLDpD7lvfeUDijsUpK4d+c7TOj2pvwQ30Z1DgidrIbRdcuqyipAa6
as0+NllKoBouUGxtrc3RYkuUidHPWdPrDye8XGx7PhI2YTbjry9OU3kyFT4K7zX0z8EO//N2MKYs
s5LCZmIwKEcEkHiv1HedrghwzdVENVgrbC+OCCJCJA0rZ4g7XxCHvc4QJ4hVk2YGtVpMNJpB0yyA
tTAXsV5AFmcAjXrLv4SgJ2J1UQF2YrxaheiTsBPOLkVKOlye/j7MLRyZIlFgs4LHnXozjhVnX2BI
vfYDQCL9RVCA39q8FPJpTxhZbTsL6F34XOvEIBKe5MZ4Grn8MX55/LWqF56RDqWQxhbW07Afjfoy
X+hjb9SInoC68df7yMmYyDlinF+3TLbsZuuwH8wC5jo16evCe4CqC4FJGOzOV0wEgUQ/oKt/aN3k
V1o/V7rKiIB5hXjmIJey+MU0hH8BUDqt/tkfo2gDCR9TnuGFQEYj8L3Dp0QSN2eZ5lvbRvKPpCX5
LTNrof2RS4yUKPtxEyP8oSBE14KoSC7idNfMcK0O0h3NPdLdLePgb6Q688uqfkmNtO2JkZ66HjxO
CbK/1CIkXnfoHZJ4D/xzWaSZVadEBZKyaJ40ZQHz/Ol9tDav1z6+rZQyKtogJxCNqjofSwKuF5Ah
oZuf0QLWmfREYl1Dsm5HAV9TooI0H27r8OwlhGxuislNsg78voLZqCiZ+UvW+sPH7oZkUq76zGbI
GdSZHSc2v3HYRNScRQ485UaJ/qoajmRx02EkMC9K69FZm72LymGu5w40n5+oPeBpaiBH65tLfAu0
WiYzlcMzR4j/mOnSbRymP+kh8w7v8L629l+Q34AmMfl43Xpmfwuu84hK/xTOk1BHEI5Xv9hWAYzm
4/nXLEis2BiKshhCdpj+SB0lURsoDF7VyB07n1cxoI7hgX9Yd3yxE1qElxS3c2gWr7I8vQRvezo4
rYte96qQWU/heEkGmso8cSVlC3JTgENd+TgjFWBS0ScHSVqhIgsfJmdYA8IXnbPVI7WUMRQf22Qf
R97gQJgpLTbnmLSTDUVjplbEzxbESOdxLT04vtJ240hxiz0Z3V3apk9HiaYwB2YcYbuauKxN9yQI
vFk/eEf5Q0+ZkTcEFDZ8o3FsX2jsvAbc2d4UrDVWaYrq24yQ6P3VUVhexbbpEVhjt72IGLWQjbuA
+sJn2XsiU98nsfXIoQglf2YKUMFqs4OWeNXyPlHM1j1Sy5Exhaj0fyUINNjKUs54Ftx+k+KpP2Ad
pfK6Ff4GoYMu3QdbuG3oT47Px0OEgX7AUErFDkllfBMunbT5/3BfYhgOVtlyhE32eynvVQSkm0KW
Qv7ffYFPLAI5/PnJY7yvAsD2ecL0W9tnxYU1q2tHAkRP9SvWsEoTqPXCC+gar/0A89DgJAoTjxQc
bneIE9A4vMDWgv6b6Zw1tXiqWyG0z9pulxbAbaZwRDmx5HcE0GVMKDp/lxznzQxPEJ4b81qaF6xl
dMrt5YPAWAXeXDVg2rHYcx9RiHtyrjBvn9ziMn9p3hgGKCw+FnratcqAGPsn8Nwz5jAFDqhz9NwE
OgUVWSGCWM3VUXUGm10RvpaahQ4w8quJBwD43HY5pV9PGXZ8sdCYguaS4Kv0TatvpYMNg5y1c3oo
9mYd9Z4wk2xSbboj/kcuZZv+/G+OUnxX5yGo4yMzAJuxcNGlMh91q/RIxYVPJAmRyiFWSVG11jGJ
4WDDT4BSLHb3Pt8l+XIJvF6x0IaCLg9gOog7OxLtRLpfCxIb7Az00pYs9bDS59pTwokkJQC2sVD3
4jT7ai4RRs1TqupbIwK5L58070fMI0UVVOxHAekSqIbB5h3iYjLLrkbn3ap4Fmney0GP+8Ia/02O
l9lxyjJP9L2cVItJ+KHxRkSoMsSEw4mV4sURLEbha/F++BFiTdfxr7kfZ+fyw8HOV4IfSoMVEYl9
AtWQxoqIUgkRGBL1l9tqysKf6mWK6DIHcsc8FXY0lYUDYC0fRTiOr095leVw9IRGP7B7q3ZPqKmS
h7zavV1liALkr3GcR1jSAZZyRbDIKXWEsl9O/iDYzLS8/FPEE1D1jc2DmrG9K9yui3iAdYFZD73w
RF3rn58JwSngvIq8Br32IEhBPIw46iKltO8eZjXeEJLOZnBzUinqfO8nz1lmCmlexRjXIk2ZvPxU
TZOEFFBiR2SLll1m7xpCjg5SglT9pQVs7yItwxyQsODcfPwpVgbrPFTH7dRSbHDnbhZv3MT+/0DO
YG8CNuqQq+RDEFAdi/sitm5vjes+66HXUZrbED03zZY5QQhmfVWjfl+p6rBrbvjTeNGkFp/XPmsd
bvXBvPWuCyHioUn8neMONJYhwcSsCYghKoQhB6Y7JI1ebq5h0iTM7bhdEutYB7lajHQ00Leb74Ex
1RAVrXnAqf2687o9j+FUei1J2rFSAMim2LA3A3V+AO9hClM0uxDmfcDQGvCe2yb576LR8BPwfuAe
PoE1u+64fJr8jjzVuqeScg/SzQc3i4kwF9Qg0jxDf9EEoWbkivthP89+EkINlEjLGe1VTINlIIWw
v62cO21oQxcDWIZxLvYipCrpVyur+qHpOUTubNJ295izBlueujIKag74rlSD6lSmPnzlgxOY0zzU
kYL4BHjqIusVHrM/euFwFjqBF33rmF6ysvM1ubyGf66pte/TE+ZSMITIzOInoKzlP5NXu0wMjgDq
vHskw+8W89K8pmuJVyg+shncc3hCeXM1q5p0EnbpPfZHIyLV7Koee48en+dyhK7DOSZV6w8ox6NW
LwwpY1HZ9XArUWiY4Jihd4NfCAo9IjfdqgEA/zlHrucbgDNKho5uw7p7eQ5kVqhIWgt7/uRJ6dtm
M4uT7Rz4fLT3MCx/SOVJ9wNJupq0Yvno4Jh1gimO0Wbf1iCzjODMoWrkHene9dpP/LELlbwNVSjy
5wZkxLb0ahmtWgiNMCwLTax3jRehvYqeanb30/gsTQ2Dotg0fAub0kYn5cpVLq+Nw2uwrpO1Uxj9
xjr+L9AOV5RiH8LHQ4Apjitp5MsFweKMIc0M+fonTnId3foYow9FGTQWARhYmmu1XF+EXsC37nOD
VVxwgW3Qf5HLVxuxB9PTLe2Pq69tThRFu3yZyx/jXisvhKLU88NF7zBlD8qEYFCmyeUnER0LszLD
FHBmHHESOhB66jNkqQB3PH+2kLCyjcjiPaztqPzOHQGzp14foDKxhLWtGAdyk7/jtO2FKxKTx06l
nJcCvgGd9ut4/RKy8PSjZwVKUl7ilQlVZBclZhlgEuci88yRMwK+5HqpYxI6xp4N/C1amnmp11mI
Bmqc3gCRAESGmYdzWPO6LJgPnNyUDD0UHewdi/x8g0TgOLKpnXf15+o9jxwVsj2eOx+OPqgbQSJI
SNyHhWbxHfaKXW9XZkm+fx5i+M/FXsy+FcTN4eAFB64Fm5GsxcUgOsOdmheHNETCXUSCLTW8TSBW
xc0OIbLBw2NnxRjZKvn/6bBXo6jrMotD7dAzL3k8cb1bWyxYK5j1IdTjrDTK+lmHAAJ+aELCOu76
ZDVs8KiliZbWasMa6/ZwS+DLit23zKWnPY9acas7fKiZ6rGhyKXaASHVYlyq2OFX0VtTzLPyR+G2
dQqJ49Pp9mU391nlja89oGHutgkSUkp3uDatkMRWKHfZ2R4XD+6Gwafc6Nf5OFlD1ArtBWRq/Am6
7owBt+7dli/5j90Go0WDZa2nT63Owh1PUTLP0NGlYycVH0HP+GRpYJbXD4rVCmNf4HlCrq/QCyZE
EbKB0bxfCyC8G43tEibiX812Nidotf0WJuURkpozD/ScV9jBd6f+/EhGc+mW6sS9SJVQLJosmenF
2Ux76Dt9WlGeop+rTs38zEfFWeoGcn5WWOmIBwlCKRx1ICpwrBukgga3gWTwc/e37fZ3Kd84ZB2Z
TofYPJ5NOprKygKIhvu5c1Q63osLnvuTRMS67w5nOmvlHkO+vQcHuFST11MtV/vyX2SkjTbd2dw9
D4HsrMuyfxkgqxbYTCararWFor2koAqQRGUy0+XCuMGSLSAf3bzlTH2Y1zHtdgBmxm4BpgbpORpW
pFn5lfMEuM5jgem8/KTk7GCw/EvexDNnEicWgEZzWbL1odHzXncIYRhA1Uhig96EhL/EzLjILK2K
3SkMVQzaTgxqpfsSGkc+agcip9F4wxyN1DNRfEiFkU6N8kP3kRacG4Pbj3npLH7REAdY2P9xawZn
H8Zbv8EXGo0SMbHkSgonol6voew9syAFrq93e0GayZOdlMRwpiL29bkp8IolT84msOwfh7w7HnRl
dFt1a0U3jMCypTduHsjnKRtUYRUrSXEMPhfjzC8YUM/7u8TQSnVyZdU60oNTXLika6/DU7fsbsgy
hkXDLsnGy4H1BZWEP97NGGmCoonf250RMh4LcfoQZJluR++YWsQGN/HN0irWlfNc4FZjArhonCrJ
T2hvvX8n2HeyTgMiJ0hcznOU4pdyFamjRpNfCE1ycw+4JlhDD4JwF7WCVKhctMCquc3hLvWTjLrE
j10HlhmOIXKzdTtudqpwC3JOdobBC4sPVvpQOmdNWjIIzy8fIO8x58kKD2sVWxUJkBIznrzzC2lX
D3tGQR/SKrHVfHRcMXyg0Uv7APm9URWI8nsZRezbYpZVTA+dpML5vZRnK5DXLa4GEyHH/4a3+9rn
l0HurPl/rinG12132C5srZpFRLjCeOdNMGvSbENq5s6h5JMUCn5IYh+vuTRsZWmwx6HPYZ4qPDP2
et4XTrs8yDet+CbyGyX1Ba4qMR+GkgVR5kAKq20XgthVMK0w5pul+M2B1VVrxK9QoLPY/JgS5XWD
OpWCpyRlX1oXbon1yKpjXWPe3OgsQgFnWXXkYXu2HHt4j8Wc6zpPR+eLoq/P3PSPkbItrgmSZ/Mx
AFA6nrjGLWf5iNN8DuUcRlrzhxzMcLPw1ioU7D01OU4P6ofQflV3yKCuTu2Df3BPt6dwGD9kRrAg
M5d3EQOs/0oESjFv2HioPzpzg84giewuXx8pgHVtJA7Cfm1Z88xnBks4ADorygoxJ3wOG10KlYa5
MzNh++HZ9p20Vm8KB7iw3vMVsJe0pVRe1GFcvcRd+j4gtCP5Gr6A99/ELu2eMuw3psY7mBfyXgS6
dvQ8IoUshG8El/mAAvJ9mM96aRiJFaXzCPeQf+Dsy15OwvSvUOnHH0hDlSqHObYvPbdlQ4J025fA
GwRkGmOsV2qQaTQL0Zs8mlHxJNa+xjzCZc4PQzLzUznj8kTz4aqPUBjB9irOQBWPUkjbw9qVSzQa
mhzdDx9J4ne0wO2dYKV07mxFjxwZqvQZdty4rAG7NKk6x3ZeByTPODB1D87/r4CwmGf+8kAVHcIo
PMNuI4Abyj9b5tHdAUuAWoVwk71TqhX21uYn+kpkKbCxJlD1EfFcTgYBcqEZK9Fxh6zaBGRHOyCx
QS43aom2TONBW9+vG1jLh4HdwhG7xb5MwLDBK4NjAh8zAgEv4bh5KIR3CFpmdnrVRH+YV1qmvp7x
BpAjISwZWR4+bxHjhajST2DaM9l8YOX2buGvR0e+FX/E0ZuuaQuNsCkRMCxn+A/jgnVFi97cR9Nx
VF6b0Xxj+9MFS6MbKxv7baaq5/DzmBplApOPqxNK9X9jBbRJ1UcaZ/5c49/41xhJEa3paW2I2MaH
kflIyKaWvf1/6+m0J4aeaLkvY+aM6hd/AuktNVqX/KAs/oIdBh05pbrfFt6oVC9gJq970/cewAXF
pe0MKEZ0Sg+snO7lR9jsDpG3+3WsLPhcYfEcczXmsjQJgb0mONf+qDh7bzY6xwp+n+btwQ1b5xby
91HVbk4pQN8H43E5SDYqnktWhl+tPG/WWpALAImaHpSbN0+ABPVsnRRqs42WbBKe0uY53A8ntJ3G
LJRZ3bfMeJaKSLQUbPj22fnmH+yh6ikNXXD0yDoT4K4sPVOnKkWFnNveaHOaNStj1HjC0yCj3CCu
AJ9CPY1EHEORocH7+35h/GqiE+k5v7Z9QJJihMfI8gCQ39nZqKNBh6c55w4lyG9Kk1WtzUk3jg8S
QJR8QMf8E4IDB1miAyaG0lnfynRVNeBczukRKuASa4YvVWCIbtYo3zNYjj1s44XiCk3yPvpFmEqW
KIX/tUtJ4rdVCQf7oq+d+xsR0+2AI3kbNsgRmjxeJu7kb6g9Ex40/OC6pVbLrNN4fiIVHFjy/Fhg
v98+zD9GdWYwEwFrrhIbIDl2W9cs2HrXURCuTBJrO9N6oWLT4Aq/srIrY0PnkNnpoll8BKoJYGoY
fd6dFKdaBiuDlWDiBdTx0dpgkastqnupuBNg9V0xLiVph7W0jbmCviIgnWpr1K+ANv90TS/Jb0XI
QzWOo0nIRkMBp7aDHPFyKqVJGbTIG+Lojnwk2q5AkNGuTG4GRhb/qriGvb78KJJw/y4+4WVZClaJ
qcJzJtySqlNeo5gPsoICxcnMvCccV2vlMb4DuO96wYhW+N7RPd5VBO7F9WuCaervYwE/kleebwhA
ZWFCwoT4pYJi/z99fuvsTvpEIiPKDbOgKOAAvIm4C6boYvTclw0o9VqzKIlXAAPUXVr4Xn4ACDfL
O+qWXRLyROmh5dL15Y532sVjKXxGOZNh/9xVk1bvsFvX3lmCaodm1zm+cHngVshH2tzfRPTYqADo
hpBxlOk33YlUKbs3VH1NuYIKCWhMoTGbuN2VgK6KTsawsEDFmhhhCkBUFmTzWHQwmQB46JeVxzuX
56jS5sHUyQSqtkKouINoxNfEQ2oL7VFiWdrdnxe1wdXAFIB2aFy8Xi/Nf8fyKCc9psNhokUWfNfb
7bD88XidTB+fAsudGTxGjenO3pw16eScaDnPkDTJ2xP7NijLUlvqeTT+B/BMAu+qFM8z8APnIzET
UE3OaeplC8Zf0CWJ5hzO6re1RxAu609PF3nlVqBGCalKoFKI7Pg7nl3/z8RpaJn4Y4LTfzCB9BsM
mnzZgLd2dJ9od63Mt4oaMgtr67PIkmx3wLKCo4ZA/43xLKfQNgT/F6D/fYDJcBOhrT3kpNBHeDmA
wH5/uNq9tri83lEunJMBkCAeuVkd0OZDt8kZnq5FlVjrr8VwxikLrwdA6U9aJdu7njvFjA9AxSON
yqy/gilOSer/Vnmumg/yV2H3LN5Sz5i0KVwCqpQd12mx2ODqVSmJo/DL0SRZEmJ0woUBve5q81cO
E+UACBG5+syRpsJL98JjxG4L2+DABRHRjuLZ2E52jae+f3XsgT/rLql0Mq+qURcp4iWPSrn9TMiR
EF4Lox7o7SPb9Z4u8ZE5/Ur6ASmyDI2wtRe3gPk7b9XFm3UDUdWEJMD0IkXzaovo5QAmwv4ZDlwg
awwVtTpcFrk7h0DGr6okoTvVoSM+JsbSN/kBC1cSmmC624UE+awZ7Ma6raWom017x7839BPa9m6r
UiNVmaDsgZlvAYv+Dh1bBvj1YwMSRUG8qSpaDj2PcM/YpWqXRaWPIpek1XxlWjkNqP+/9bctO+vV
S5+TVRYlYljFqFXOKbjFWVYvfp77EknKnIB/ERDGKDXAL/hGWZvHxfPpvIvV2RdxSoP/bFY5Vgi0
XpXe2DZTOEFtJsCRG/6cHtErWntQAXFd+UMb3FPOncvkWhTt7QJvIK5svzRVJGPiX8NfndQLwTW0
+6ZHtMRtRAdXFeqcKccVuOmLJYR58r6FwNwGUtuJ8WeXfkQMBq0EWitc2qKmXnHPlNpw32LekD9Z
IgGBCcL98OPeQJjh8Wo44Q4IYlcgy+NqxdLSOq5Bn+sQ5k/a+ngD5jipqkB8AArzLqHa94NlM7id
B4TZqLzsn9jEMxSLdSuhv1PeJsGee1BYNw3lccddfCUWq7Eeb8ztLryZOCGsKhHtubqGV3AwR/nm
cNmfIS9PJ6cTKg/cgOSwwmUQVqR5hejg19wzIUyWw/YMa2k97EfGAEUriW9ARLeFIDMHEq+5mY7s
4I6gTwYCFqFdsufDb99DGMTSlwD6A+47iVEhzgJyW6qIOrSPr121RN4BBMMQOs3uQaLWozjgK++k
sk5SokWgdJlMR4R2rqhBmgLS0AOmVPWUPA4FCa6aQC4gtrHxWR8ZprgOovK2fNF6wdaosZXF8jiv
k4NyH4yLlJ2w/7M0P7khG77raP3jzEyODq3wamBet7Hl5rBzVZFfIv+HEMsN6rI1prhDxzsSBXTX
XC4KsIvg/qmj9EU0Zv+OsAFPFOK/g+HM90XQo7ioI+YjsMuSU3cXjdCpPcYPmoCQ92H1GGVhP4tu
SA3bESnoO2T4XgN/sUXdJyaJWuu18erlDLfqnO2ENtbKXQOLjKaxxmazeBYSnGHC2SRkXjbd4BaH
FhSAUH3+neyCwgkLR2zQtfoISZkcm7MUmwog9AWRU6Z3eO/Y/o/lbc5XgnBZ5bKM+0LcCq6QmqXT
6sWlqaBW5U7YZ38YNrpzMbsRP5v9j/XUWrXvg1eVq3ReMaXnyAizFFSj3HbvVYU/ayD0/Tz6vNEc
C3IGgNMj3whVFqgnY5B/hgyisgpJ8WE7xmohJ8cyUT+l2uUtg6l3yRme0aTqCloTswTtdijMyUZZ
Okw4GUcmOL5aGmiexImDgZL+wt14/QpUEhgrURjyZ6W9u3Ji2HRZs9xT0OUUoF1ZMaJ4bInMce0S
GwbbMWZhlRWi+MDbLvv2vLnMmLaJJF1SYcAz5HssOaiwuHa3D4xaMvkSFCsNN6EiE8Vi6Wlg66x5
++YbJ4r1ZyLnDW/BVpn0hKn/+evZFkjXLsxFOogSLNCV9IxCvAgsXh9TjmtlPK0jPHetqZQFnZzR
Qlt4MlfG/imZ+FosRdgIN7hpYiyCHkZqtw0QYSUuRa6FWDMY2Kfvp+Dh1XN8OmLR9jMNa0Cus1FG
zg9S9ZCvKwMjXC9vVBNeG/FEJWMlWCeGQI5sE7h7/+6WJPkgglS90+kLjtVLBdgJY4fJkQXoI3O8
lbgOCqemuu1UYPng8DRwM43zyIkEDv2MYJRmZOWv6edBYP0NhH3yblbCTKIiPRJqvneyOBD+64q7
FevnWyeV044Y9/oi20A5jR8g6uQSlQeabXm08fSJb96w6iKqi/FFY1gL4lEZMC6n3EWcHaiG+/H6
mjDpmwCOdxAgB/WGTr123YlnVK4+361ObM/2UBQ0nBrfjv1cHNlUOVwyQcCyr5bNKfnJMhB+NHQo
dXieZVSRjh3z01SYX66ubkfrwsZGthVp0w1+b7sMO/RI90GjpHi4xSo/6aUyi5q2VFw/REC1gETP
aSBGyRRSKZwF5K7M97OoeEHKQcg5CuZhGSzbxvIC8UHGTIWaX1Dl3IAKatFfEh6MCH1gl/AC5DMt
f14ffkTEz7IRxjIvNfsYS+jKBCqVBaPWb/I3rjRquQ/pGUDCZ9TlW81/7gofYBQEMNBdwSJfY4fJ
7PnwQ5G+wYw5s1CAvGGWVb3Jyj85UaO5BQcZmiWyiZyk9+o+ubE15tZxy+a/dnFoN3sTMzwfJ2EQ
odK6xiHlAdB7k/j/WwnG48pDZQrUOeS7vVRwTte0UiE+t9T5wIXfLLKgQevSQTsXp8AyO158M5bl
bA+NLQ92OK0GwZS9+SKgilbl9kCMsFN1pJ04qdQqXBYLM43idIONmdp6H1xetJuE1Sq+NhjAwYI7
W9pRLJShY424dgX04r4TsrwNRLK+DSR3ms7/5I6nMD7saAqqFOG9kRXKbu1g+00ItfugMB+WasfE
y0JBVrdSqttW1InXNxEoDsCUJMJTdZX24hWed2zssbUQsDwts8w2j/P4gQUuM9SZpluABZlGaSzO
QUv5w8Dk3bVPN0pk/KzpjEImaiRet9fZotVztWlEkEyzHg6MoQxKDtyKN/mvBw4BcuWU/eOssBA/
DQ0FclqWonxaTvxUH8fYRMOgJgYO4N33UOcYvBr1UiMBlS17xQTVRQJL1ILwmcixnU99vItoqone
Yot46NJa8SwvrM6HNkO1g+Mb9zggC7rSMD0Nx3f+EhLQ+dSTIqK02Lbkq4on93RcgmzLmyGQ5bbK
QQNhsntY8kfAwBEbaoNUoV9RTIeNJXMjbV2eRI4TAp6oLWs0MIIk+/NPI4a8SVT7ifXemgg8akNm
5HuTwddDue0F1tB5SGxEuT9f7tg5I34IMyjs1ji1IVvRISrJCFEdtKstAnKBfjx2yqL1O1IvkU2A
Kdzhq0mR71yGGYMa+mexeF43R+3gaytsiqDXDcL7b18+X+RpJaIVUqKHcKTMPiqb/ZN4dCIjC8cs
/Nisgcd7hSavevUKbe19aMrMUhUR7Ja2LrA8StUwNFb3vqLijv6W6kZuPN1JaTfbEU0wW6p6mejQ
vzUzYLh0e2J6WSpFfgbset3cEal2mMrSEg10upQtcwb71mpNhsR72lg8V9cG3OoAWsFekpwMoLAJ
09ADE8F72nqSlQB79cj0Qfb9RwLzaw+oOcft8Zx/LaLlG98iqpZ+sPZu2OCJhEOSk7k9H+M9nDHT
q16fRlLrGuQfN/OYrbwVVMbqEL5N6CEjBZbKuR7OssU+zenyhlpjQWghIm5gJMnY3dIqPsZMBkni
Q+mA949MVCpZFsPyx3BVLz1xWbEr+x93aZmeM84J7/RcJn4hzm0JHhEgPiR1pD2C//NnL+2KlWUa
2LZVgEI5wqx0wpptu2WVIIEmr//EBPEn1Cnw3vAu/58PCzVtcy3VSMqQ7lrYVaJ3M+AserFH7sAB
39uyU5LZEn7T0jOUOWhJ8osGH0jYvuDgECJzHoIzas0l7rsD4cMDgTxkut5NsZk4YlCODUs1GqKj
SDENx6t4ZkxAXgR3EpRF0FtMjYd57dZJVGQXaYpeQ1PSMlUA8ARfO1cNLcJzt8Hb2r65Q7FTrc1e
NTvmWxL4jq2YDXCnjRh47v6lqPzYF+Kp0WGfAEkzNppo4zGF6YY+MiSlm7L0avkOFHqr5X6oMQPn
kT3cfxur0C6FXkOGAzWCqN4AlSVJsvDmCJ5dI/ROTw6aYBB4srmNYngNtfxRJFOxkVob61BeP4oE
O3zMdMaX1qD2WpwbBRUUpckEmxysvUdmOlHE71b0bCwG39b0W2OXpqU4lE45e+AncsVLsJSCNRyk
sbm40VgggA63NfKjKXojUBHEcJqszREBhOfe68YDMVKsOFxcEbyvoSWfulwt1C6NVdsXsCu9TkxJ
50Jqjrfsc1ql5dLrH4IvbV08YSSXtk70POOtwKBXCzZYGmtqcuqJU2xj44v8YNicH+OwM/ZBU+s5
p9QDM0w6lrN4C7d0cySHDqRxx4ZaN3BkQLsErfHLZ08KNfUvExf7F6tjTcSsgqMZZItmV38XOJOf
mXCXIxjJn/1ZvnF5xM6wnx9tfnfqeslqFlcKDBeM+ELoTkec5Bm+l5r+mQjMeH4dBSyjzknE6KiX
SgZGX/DJ8nia61g9SvzQhBvAdbFulgG95ree/bvVQoRbGH5PRHzsYst+udSUKofWnaeG1A2pNJYH
vyicsnvnXtQYC+eTSOmlOkUbpop9xPcZYn9FqgqQF1cx75vX9rhU/0aFc07dzo7SnROwsHzGKSJV
iMqehjasZU3NiUp9xsJm7HQt84yjnZY2uobRkYVF49UzWkTYOufI8iJtovd37BzDR6r5iGlCbvem
bhH7FWIeJ2VN7Sj1a282dQFIwphrnSA5EjD3DWsqA3o97tRREFjsBBhaX2+JECCVe+L9jA4V7r9x
/Fxi1brQ3AoIj6jPTCk4xONJimBiK8s+UjvlEnZL3TZ9llVlb5bueVutmJAuVxRegUSH3YrgtgXK
/KjzDn8NahBxcljCZBYNH8d26e2VFiC4IQWqGnr8qnOyGh3MbmOD0GZ8xuN1dI5VkPXMVDj03K0l
WUqqjjhBa+6wmydahH7OycNk3m8wrF49eNV5An/0yLgy/FIP9k6FQVq3rtg5vW1uN/hKR7DrpPW+
K2LPOaGrni0d3PRZkr5t+jFKV2DoZn3h7wRb6d21FD7oHR1kP+z4fvkNje6KNdVHt/WiEU1OTvZz
Rc65OLM2TDASouZqSKZhhD5NpfAA0GY7fWTjeoutB1ScKoPUl2w+ywZ9yhUR9DO9H4gPOL/0Tmub
HCgD88qYcZcWSvSArd4+zT6DyXqDO73d8OQ/OLEm/eqA5A/aoRZZXEy8EaSG51U2hiDMHcVWfqoF
YgS1SD7RddtEhiYs/YJf1ivHpLSfeoVniESgTVV5wakl9/xTeCKOQ5AHPt0wLanZdUQgZV7ZoTIv
iuXcc0YLALpWeGJQygwg80WX/0DcN7wPglX0DkxZnu/c8BUTwlx0cboW+yxOeXlFyGmYPKUkNwHx
IS59tMZMWtgcpGXt/p402DuaFA3vy26ePXrjzdEwJsVcy9S7xJudhWvdDT0yS8Y2xfbw3/lQgN8e
URbqe2jntKCEf5uedGKEgd9pMJSIJkKR7+IihdZlqgJG49X/+V4V9ex2YKtNbLpjx3w4MmPqbev4
BKIuPCZPI0FJsyjxRjZkHbVxWYfr9iW5K9aaA6yQ9MJumdXHEtS/ChPAsqHj3w4MjGUsCJc3GsLr
mSNtjSFyzZo4LCI4CnUcpTDlwdpdiOcTSvOCUxFaakQDiCce+bgYWQrborINEiaNGoeNfC1y3qQo
yJNGL3r0VLQPfjvqfnfKSqgbDA1lG7hqRmzXJiMVE7FWfqPBsjq/HsGenJ2PjKN2mZZSeyRBFd4m
So5rNusBciR4V7nDjXHVln+fwYAmQRzFU32x7SCIVIRYF9bRuK8Eoq75QSGO2qbYJcVAlRwQ9zDU
a/CYfYzofFSncQxQvZX4fFJ5wopbcfa/3SOCzg9NYBUg/per+MXo3OlWOG/VHDz1xjL0E2uXj6PL
kzBsPBzH4WPCK+ErpMPoAR5ynyOwVDa5lAzq2OTlPUlYaeRsAqIOxerexJ3f/wY7Gmut8ZXRhArN
UHRNs8n/5foP9UVhoNFXTaicEXx1Xqh4CV+DEYkx0N6mzWFedCMFgEsZSiG+7sxTdo80LbnLdNxe
IiY9upGccVDa8A1OQwt1WjHqCgXhF6UuJgqU/mj+vlGjsBqsYT2cMrgK2m27CmhK8dtaNK+mIY6A
yQiZ6UFu5CPLKZfax/5tpbY3StM8filB4nFw9Tbi9SIaDUu5EH+7hzDU0zJmsGmHGvpZrx8FGvU2
RPdJOEiSh+Xwd1zzwyptQ9TKr4YvB51DKjxLKC5/6NGv7D6iAPk63ZrI5mftz2nOsHrWqxQKSz+t
8ejtV1x67a1f/hJiVlqEuGlvJ2EqYCC6DjxIIzhdTbdQToUXCWxb+2Kgghea9O5Bc5cwiD4gIjR8
Uig5BhsHSbJQJp88av9d8MAyoFW8wRn3Kaqs010GqWZobQ32DF/IolOdqB1gr+ZkjvoHCX8iiVvy
619nb8o1VVbY89inVOTQUTEzS/C2evYOR4R9hVpvhcpbuiA2blUwBgy34KUISFazqXhO0rsowkqZ
qcDQVKLNw2SuebgOiyR0ErwcnoNytz+qp18NgEUx7jsdLhTupcp+MakAp8CU0pBAzlzfy7sicxq/
dgdYdFaDmWPZcwI5ziRXfUPm/+JL1dK77Wb7p2cEuBHa9DZzr9jllov5Ce0P4WsSSZ4SOmDkiHrI
UsAVQBgYweHXXKMXcucnH7GG5zLjrnwTJv8+IPvoiYfErC7KdP67jEhn/dsrZZQ0C8KgAiAyff0F
5OLbh5xRGT25wbj/aFrpedHl7oXT+zGG22H36H38A91WkLcnjiaCyyts8OG2HoGgYHlm6CwzYWUj
9EWbdiPRSpTDOKKPvDAYW/JGXg+SCkFF5uGkClpgP9KkiQaLuhlj0G7RGwXwQq3Sha9UDBxd34qX
u1C9F7Yc/VcnhenOJmcMOP03LYQNGYYnbKwlWx4Z5auSB+Ly3FvovOWtT4XQGy904VjXaxlucpze
cGgch/yid9vdffe4n3HhW9nvPsK7OrRxBlCy0FE8bvGSMf6U55brUg/3TdWI7zk/XomXaUJvk51N
+jkFP7XgZRThlZ01HMEyxyHjECA97ow/cjHztphQsHXSl7XXyX0w01KLRlBehBaDhDSIddYvBlFO
71ljnKQXonfGjAkAAdEg3XLdJIhvuDY1oqfrHS8ll0JXOPqhyKeAZW2dTsQcxCXHS5AndBd3Z+4c
HQj4vnOuOklCQ1xlg3eMAp4/E5iTObVnTXyXKYrEVY6BRLlOEc54YRZ2r2hLMqjfQf/PbSFWtpAm
xnsDGu/y/Uz7tBCKssaHyFdhaCP0Glorb4sqrYIrvwQIAWnXAv+6TuOmDCR23k2w9LD1bXuo1qIM
8CilVIaUJzl2hbmgdO1m7IjSee9PNh28sLzxli/JWU0PbRwwmwArmctl47TsnQl0kDKAoxMZ9vQk
B9cm8YEF3vHsVGZcqlWLshmOMqJNtlYsQmdk16UykKa8VJpVQ1s/EHAfH+aAHEoG0LfufjOby712
pEQRmXGa64pPVUIBEfWRvvRaK1fCnI3fR3XxkC9yso250MVPxX2A5fIqjXTAoVDsWlISlF3FdcjJ
SwGkk3GFE7VKUlQKydF/Ls5CwUqGFcd0isGpPNUlqlTIU7AQjqpa5RzIDiusLv0AIfwYeyKsGbTA
/8JNUgJbRALT2/7mqOuzoit6Nap9WiDkKMHY4CXDEdyobz6NL974iXOkIBKAodm3H8WotdFoG6t0
qH350ElkriFmeK0Z6lebv9H8jAP1SE79+J28+rop8qX2uVmGB/q3jAw+/TPsHVewwyN0mrCQvxez
f9MZJXrlMOC8xeS67NIlhdJaiCTvyXFy/w3CniCc0tb8+Z1eXIgRjOPAY94vT4zh3wqlsgD97viX
DkAClu8VhjxfQAa8pOHTwHyEJuelR+DAXUjJCd9YPqraVK8G2ATrBTNB0d0SLTo6zqyz53Yn+RRJ
F95XOvNXkEqTd60GWLHfKf0eAYNyx56X6mou8DIuPwCgE3MQEKUozzKGooBjDi4z4vakxTxxPLMq
wmN4GP5RNVeEgdR2EsSziS8tZGy7gJt8HPOWTfHbUHqRAt8ActDYsfL4JvSeU3jyh3EEodEF73qY
4nqQz25peRTCI/Q0tkJFMwpYvTxsBQxnGZqgim3zOW+0Q/tG7TpWGjvOPB37QfMN41ZKZBW3dZK1
GC3RsOaVqWReP5cC77ZVfUv3L/G0h7V8PyB8atLmIJMrcFE3XFYkWYHE7dy4zMrsrp5dnxqyUl57
QASrCdIYSBHEm59oY1NxCSeYchxEBHGuS/VxYZ0nwOeW/bTFMkmgSjwlVqxpinGNfYfL2nx59dC2
B4FhWc6PlYMZcOjZg+mgbhJD0EdDViiAg66XkZllloU1JvImjNoWM2LyrWxa4RbAMinDWFAEzy06
TysbL5BHnZasP0f3nbp5Hr2rsFIc9OAT2on72jo5tqKGmON6dhVbpVvHOn3iYtIlfvtuvBs5TARZ
7qtKbdS2sp9W7mNNQFwVu46ZtY2TaxV3ZhSsKK0Wm9YksJGkyqEdRLBCB1A4geD+Ji+pXxl/udWJ
BpW7SSXK7qsxgFOjP4rs31bKfmMe/oMkahboo60ssrhACLtXgFmPiPCAb5KVquTGfSMOUQ39tUJ5
H1w/kVjfcf1Z6YrhRLefi0rWaw2462u5kF23gHRDAPF2ca+h85rUubcMzygt5bXETcizgQnHZbta
ulQW6ON6Wwk+MRo4UwZEG1XFsfKdPJebjOgEaBwtAER1Rjm9+D+26wyuZ3fze15tUQ7ZusAGWyLF
yAZErsV43VHFLI72PN421UQ/FnNhs99baJofuL9vbXKvWBzKGiTL59op+XOEwRIV7645kn0htmu+
gVq68xRjwfsqRpwV5fnk6Nr9HV4Bdl3KPGIoWRa2bAmtkxD6m4JlbO8XKZ2PD5sLMcFMGxLkLVNP
hM0vtiecVzcc4HT9Fog1S6rJpGZMKRKe07iuOiTlBmYJhHcH4HkXtuxgP0DSR0PdHutqr5nPgm0a
1Lo1NO0iRtCaljBa386mgqe+t6CUS8faLQw52K2jWZ8VDGaDOwxO55AEw87+sMDhF0Oap05BgUv1
PIB6j73JM4qqedwzIsS9+HMnh8rb+UDzNLNnpqOcujj/Pp+6UGKAsGqE5pkvH7r/EUkRkoi0nRQk
6MQv//WyIIYi+viEIVFq7ZnklVR+dled7BHfW221muid6VPvVPOulvS0cu2Go1RaFrIw4cMjrxH/
K0NO2Qq2qwQLNIhV3UylBbabedEwYrppcjvixedgV+KwdO97NgMW+flmDLSVBKlAMgTwo8KeoaZg
uw6aPz0OqtGX/qRxPrm1PKwYhnIsmV5g2JLNlc3RfANTfdK5GtTeMB/buUkUHG7gvGYE2bG4jQ8w
8EoGBkaTyi8rIsoNWv3gR4yKx67n/6VdYlz50J+dt2QZDXxYt+m+SicHtzQyRK9KIgqm/dkxuCwY
41L6Sll/8VXpCD1uorGvJNiJgkiK+APmMb9i1G4SxhPRtbPc2/kLOQtnNGQIXjS68XFgEx6/AUcp
GQjxCQIaxUYIwm4LTZ/CkfFbUW2NR88rcyMmEWtd6aw+JTdEKWzkYjoe8Jz5gjrLpatNQsd5BZgC
kjuO27Dra878+0PZxXG4P8OrgOUH2J5HT7pU0oHw+7AMzfjfRs/y4GmTlU6EcP1cHcTR7k/JEEcY
MYjhRUJIhaP3VMxpO3+z1hIUecJ+CsgVwOfvAwOMmSBZQU/CasJrp1oBbf9dNxAFhm2vpvaMlZzk
w2rZMuZGikonDO1AvHqYnJZtHdvV10obZ2Gss3olIBgvU6+voEevJlhBdo8V/u7ubAprvAlysQib
iseUjvDdL4FR4MU8/WoVfI1PIz0O3N1DSLROkZspzrCAp3UX/egsKJssD0PJVcsTGEQpA9b7jBUm
kopD9XwghDuDGPpiqQCDQDrZu59S4mHSd/VPaIi9nza8UGbIBOuTIs0QU+30p4+l+7Q1qAvPrlhz
DGyVagcjtniojdpSbVzK7LO2q0NZOQGxEo/OD20xkX4d69bqLnWzpHiM/g+3n7cjX//RzMjzYX1E
O59oZdGGVyGLtfwOUXRh0hIPCDoKMyf4JG1Qx1AizAfV6rOyacyTVuXG7/qgMFkOsE4XSU8mIEHT
vCHQ21RwadlgqKkhPWHqaF/6Yeylk1so7bH5+GqgoSoNklOQF1unhEng/or5j6cMFo2UfM7Il2J1
d2DUw+9NLOZ3gQ/Yt83FCATGX0xEZfP2zyj9DyHtLruPq3WMr48CMfizXyjALgiOaQjZYZ1nGweH
8My9nzqZ8SoYmj/8G8bRhdt03aw8i9vF0YFewsNWzE0CwR7ycIn0zQcmmZNmJ4OE5NKM8lUNp73r
0GLztzHN9DkpTaiwHvrKwa41f10wQjRinTnxpEUN3b4NUIso/1bGvgrbBEf4CguTKmEKrhxk4aO6
+M6/9lSIe9U4bwrffIfjWlP/gerE8rOxQzQZuuq+XY7CbjLnfOutTSDS4X1B2Gcofw5y6qgpVHnw
2+zzALUVTiC5uKb1ezWMxJBpfTMIjAsXaMMApX9q34ifQpZ0LKb1cXwB87klHPDinoNsjVENbozE
B9OUpl3IW6KPF6NFaKquXDSWzvdXGcwX3N37GqWPQz15HiAf3r/BUY9xzgP77hFLpue2Mo8LSNI6
7/Loru44hZEfYdbY8cQ/kaq7fBaRJR7gtwLJQ2Yf1ffgFgVu6LxutEtLv44V+EB5weahH/4Ip55I
XbmUKvfElrl1qygYcBLgsXuggHQ9flaqH/csXIBeJ6JY4/ClzpGs5mp2z/2gXBHMcalyeDC/V0Xj
0lIYWfiKVDqa6rZ4kwMbf4QHuBh1iOtRBZu9tKGHaj0hKXWhr9RrvjHhzkOwjF/sepZ3UAxRoUQc
t6eI4M8UnkK0Kol+D/9sCSUqWi+HJCs+TQFGVW4TF8w2vYZPcp29YkWETlWtUmdi3sG3Dvga7Ee3
rQHM+X6wO3II8Gx8Ef62DGCfwN56imAbVZ2FPqqMQbRBH9J+JgWHAhQSxUhbspnA597Se5NNtZr9
lV26pxorDxxt3IJrwum6o83H6fYTdjdiRe4mtH9rZD57j7gCOAcEb2oCJekp6Xcw6srk3MvXQLhK
fRj0rNln0TTup+oC/u1cm8+3DgQ8Hx94UySgfNrZCAZiRo/fTroGgk1vKfV9hTC9vFIWlEeQcBJK
wQ5iGeoReDAAivhBJmbr/GhsVeuzeRCe6v7F9SFTiLszHcWWNJeUHirSrgrdFXu70AbJi8r+kPBy
Alvufg3VvtA6zJ9wx+wQTY4eKXjeovpef/gbiuZdqvho2Goe2ML9WVb3DrTyTLD3vCvvkTcW9xdC
vdLJ942SoQ4/tzlUU2RrOujPYeJny8Z81MQcJAqxN51T6u6FrGOzrKg2EDKuLwIDGLx0Zpbv3eJY
TtI4nO48BpQEbRAblTeSNBM06m7BHlg7ohRduDNytQNsnxwea96H+Bi0qUX1M/8oNvGfRems2fQ8
TrcG4eCHAWL+c2bgrdHuBSy3SMeElkXoJHTbBxIjdqwUBOAV+TX7pIotqYj32lk3KUSDi7/iWhxf
cVazOchRNVGd9YamRr+Xq2cCFVyggwmW81AVvMcdWpEO3UBuIRI5vQtKTIRdq0qKjPTgYBtUuu8E
hnHg1cJX/XGRK9totS3ZTMBQj9nkwhC9nePDjjtlccevJcnu7zevmrWqcGKCC5SbMSCybQNJ7XJU
CKVBAnVTdlqprxiLvENijPPGTenkIt/yTrLplJuBQaumBzdw7s91+bCkL66mA54mwa+eygho0D/K
J0TK5xhuXqOc6ATYKR07H9tFovZV4GNfD0No00wujimYaE45jl6H+NU++DbByZbxaThubBYBUjRo
MD1yHjtUlD2WQ5xLwKZx3EgjiKm7g98eEbhb8ihra78Z6O2zpeTS3Aj5F3mHJ2JYM/+/HswIkyxy
QfoOaWGp0UzUPQc5M7Y9OwqIp71Ju/9iDKaHwhLWrow52XIUWONaTOQ1fi7dVz0fyBshFZbU9qyM
oCROvAhK5Mh6aiyMlnSx3y7e7SO5Q/Glv1HrqxYCaNwSc3O0FO1cIrpvDcpPn4r2PVBK/4CIoqPZ
mPLCYnflADVI/J9Q5WnA4Xioq6P2W97RKotovrAd/kgmGMKymfBnmDO1FJE939i+IH4dwEuCpRd9
k5dRQSELSEGyPc78ofl+BU1l4lsMBZNZUutEgdUwW7KYqYLkmZyFFQtxkk/oKe1vhbECWz3fbDiF
/6LZH0UsakpcVLXFyhI1WJ1oKbnhqZHORP1PXsCrm54jTkyq34lYKnJQuiAYErMMTAZzsbFrehUb
3+TkSLZ+x+BHy2iSdeygg0zQZK/cRbuNEllKESUU16piLX9YroXlL1A6jJ5DSwRpazyN7bBGDXS4
n0w1f+el3Ctm0wPYmfXAkjTPh53U9w29dn/TYUYkM07DUfnTDniipmt9+UBOxwu652pl8ux0wOEr
vMCC2nKqaoHbEekf/GSLflBARxuCfCwaZttlTw6uk+EEAhgMD3lJussnzgivuVuXXd/uZCnBenIZ
U0fNckf4WykyWXwNKU3/Ilycx5a0wpShM/LdQ2r/QuD+zye2uDseJxlHpFDeU5AEfm7ekgq/DQoi
80CdroLKY6APs1HYxAz7zIV03/9uHQDf4qC+lUO1RnA9LpQmKZH9mZS25bsnLxTrKL/Rt99rAQVR
s9ioieFMyCkcEx1qPnAvEUoGGlM9U/Fr79iRDEVod62v8ciwyiqYtAaGArw1WHgNDKinKcU3hR5N
Nq3SYn9bcFSX47KnYg7bJ0VCdOSV6ac1Xdzq2/0mm20CQe14WwAxHEoUn55kS92/XjbFazgBOvln
3lL1NXg80PJCUib8m3ZGeGyY/2lxRT8KEPfki2e+qNtNVLlQFae57aVk74y91CAx2ynN/5CKwMBR
bcxNGiPTRRQKoUJA6wUpWSGfKLCg8F/F10EIByuPuSZUY+WnwpaKWbavPyM/fKgomTd9YOSQcuLk
aVFoUEJWLzfAn0wFph3cubhfdTxSrTFHF36rVHzj2gxNI5EsfUpH8vbGDUjYgjUp0K7eB8vqop0f
tVIRm3iRLqJb+VecdjL4mChlYN+y/J/jmWDc6k1ydD4bNbpmYwFdAyms3uYt3AnK9K6MqBngmXfH
sIYxfgauG48NjLZih05SqrNOPVUtQGK19/aYlqGa85x+XzLT/OTa2TqlXGGo27C9VnlGz7ydBAXA
cFZ/36sDjpWfyWYVhAWkPqk57UZ6flvcnCJDozoIXHLfSd1XdXMlJupQTLO5GL9YWis8dw9esh8r
bClHty806GGxPanQ76BPJacAZKWvSgrQvYc015j0p8nL3move5hRg9ihaUB1k0nR0ZmQAs1+xSzW
AGFhsOdSC/2Lb7UvQ0stMK1CX4tbSliY46jCte4iPaglwg9MC3GAdaweEB542lCmEPuBDbwSW9/q
rq1/bqsomYXrkE3fRGwFsFefUW13R5aUV7EX7BcAJmEfVzDhEKXCLH4TnT9upBB2kF2hpieTp3ek
k9q6HvYgqwWkjXmsKzkOj4DS6sQ/GAaC1Rm3EpM4hDxCT9dWHkVGOTkpWZSaBoH8pVow3Y/FevDB
67JCDT1/VsbcYmlnYr5wqfJpGfIeistvw1Gcc+QJOCdjmq+zWukMzgJ7Q+Kp0l2bWIrIRyzI0Ulu
c+zNmKM3tXijjMT57lo6wrQMxbImyTLLRJ9AeR+2mJc5Lh8YH3GqlzmNitexGiIDdEg4hHqipUp1
VmGNN/+jiIegjo5VYuDI+fzSZNEp0bphEqbVQzL9SlngOEmRU6oaWpoM0RNyaiXGFSrq8TLUvP6X
fztbtD3gM4Q9En0jIBvM8Ff5cS/Tl1etXaYzrhnJGbXhgrJYg7mxIdhcpfn1M5M1KyQuoOkZHxD8
IH3HlgizmgO0QwiwiKtyIADEdcoIxgIFr+e7lp0X0LJHpnxS8H4/jEYdG1BGSC0b/yTqKGYUu7ao
kXPVVpysLjk3YMSzdfPtiPLUQokmbZ8QaKy2z1yRjocLF/+Cq2iHF6nGnVsnTT/eGopb7gx4ooOK
z/hll+SZCTXfD/TJanjNVZOXdJbjSxtPaPzWWDoJQxHHDSRWovv/oQHgEZFCQjrLm2ZJfNikYJy5
Zapv9L8Jo3gnf356w0BUM1PPzZ7dUtoZVhg+mZti1yt/6/R14H5zcRqFJeuJTLdqTXexfMorMras
TSnDZ/9eqp4L/YCs8Nb9ljLQm1HCjIN4vake4aU6ubxBFtGMJguQSX4wXZIQMqpY/E4/8UeX0kDi
67cbFQU/38hvxTrrkoo4u618UUq0U59QALIeTOIg5Mq62U0BDXhOLsRhPcXfHHZ3P1ZmoLjyhPv/
4ogXnBUH1TlrEBQWflGIq4A8KE3VMr0JGT6z1YYy8cye6IlT+Mqljc3cpy+74mBI1aEMv+UqRiX1
f8/sf98+NEMCCX6TuwXKlw9vit5bXhWB2FsrebTPCLkgHiXH04tbL3biJMHjAG1HHZpygFeaioOd
Uh+r0ucd/uZTVQW+QBw87ptZ9p35surF6rK6j3NWFgjA9yidxY2NlFVsCCIsq1GsiONEffmC1nj8
r2Zh8UQJaoZ64Jh8oXYFqykazc3fazv7gNKWv0K7nVVUKQgffAAXft7IJXg0VFkaTNarSIiL+ACo
O3DVCIqjOPjwGz+6DUVOQWLdyFwgFNPb20DcOtlNpJv3QW7XwyO22i4xf8q8fclZZRT0UuvriH3E
SIOOc4AvYJVrPb0ZNo7o6KmLGiewUWij1GYGdUVqPOdkBZsy7ecelyo/fOYRbGxwk/A5fX+pRh34
7h0MEpWLccVZEF64bwpfWq2ChJDFPLj2rQ1S7zHZamAoL6o2IvFxE0jtJRt0n8uMnMypzSndMHZ8
48XF1jgY+rFdqZl492DpdODpDLCyLhpzun6WtUKXixKUGmFIZV2TffT5aAsnbw/XZJLfXLLGnmHw
ePhoD0peIYTMVQoZwO4y5dWor3Q72f4o3+RSYnvH/YtTdLFLjrg4pdKVKx+lVlHSNBPcH9r6uiuC
E4EJlhEgpJ9o7k0if/+HgOMwjWoSWIuiry12T+YmPytji5yoAtthF+HWHYemo99gfm7osn1kXoYE
EdSPWBG/CwRptJ7FB4rf60KDQ+LjTrv0WyiZ5prQqBLc1rg5FnzodB4brR0iZsOR5Glh3gTWMD9y
BhKeFszJgQ/4H4sZPnXjpRvIBpeDGrGLjiWX6wCZoHGFCurbLwpOZDzGrD/QtWaZ0dUsHeJWzi1a
XgeUwDOpxyBoPI1MhdIhzVolcWSJb4FcZLoYVj81txMzGPILLMAqrhqMu3NG7+SenoRDI5QDQvP3
7mKhb3CtLQJat2ZpnxBklbYBy5DsytneW2ydoLVD/eVU98dYmb4TgI5w2z2+OuN8SIAS3nzD/WSY
G2yIa7DArF/cTb/97UTu3+Qgu6RvlgdHq0jlIkMbmxCs1YJ8+H+d+aQfQm0geGzs8gMFh5DXN13m
jpd7A2P4ZAW94JlQdiayKofhr6VIURbpuYOouFA0gPf6sNVQSZyJu+vG22gBKKaZE/zY5/CSd0hk
RZ+nqFuL6PAV789bsw9cy+9X1GR27YtHpMlQHwuuOQwd5rzWvoIKinvR1jWw0qGTxoO0x8lidGGF
pfSvGZsZli9tQpha3iqa2MXGMXNOtraBTNEDSnA5bqig3zHqLa8o6euX4EGxez1I2gTRcAgMrzE/
wjgePKm7NZCdBAykDNcauyd11wc+rL81mU/CU+iM0wkvkJF0weLv+VXcfj7ERMPn0QO8UVfmb+S3
7sGIrhwPBW5eP56P/GFmLb7aw0ymeltYO+tL9CYIYtZEygaLJnEaTUgvwurE2DkAVn8qF28uPRS6
SEnTOkYjeIpO8G0yXAFQcPE/SWzKNSFFSJqKNMHkEpGRthhdkabY/2EuVRqfYAbtfoNz7IBU2gmR
EIb0o2iBbOIsHvBvQY+QVJFAJ+LorYpt7dP/TorqcR8//s2xiOldNV7SalhiFF9SkNzjJ/uc534D
+I2Oam3A0fAuwSlGGS2zl2eQUWrdgiCo30iD+xJcWxrOKQRiIK8QXTkSphDZGVT92QikQGii6vuq
gT8NiK3AO7RD2cu4c98C7IT0tjI8Yt0Cp8OiMPFg1KIGQ8p5yXW/I2wnZag7VhKfIZEs3byqLWFm
rmcigMNUEB2G+zY9qKewzYmPHKLgSfHnPRt6rrCF3RU8hNpYp380sLFTUCSPgdd9r/k0bB/Mc6jj
iPUscA9bmgVtYgEbPdX8wPykrUIh4niPWLQxRO3hRCzmt2QoRgKtv7LOthyGLY3BUcCLRxjA9O0c
Z/il5Eq8KHzFga6ztxcepqrlGmR9coA5DFTH9mY9EhTZTrVRSYSxVZy3Dm1Ke/FwYBE16sDJA0Up
E0yRzyHslREO4yk/QEc4yDn39e1vUBPlGDT8nJasnEXPq3EYaIm3785SCCwuntjuHeqoUHSUV1y4
PS4J9SzJjW9YRuGQmNQpDZdakjwhXKrQNFdwxr/fXaepJlp4FC4zQsa3cIs2Yfj2ntkalcC+F/Oe
am3qY+wKi9n18ps03Dmm+ymny0pku/VzxRMoBYrQH3RrvPfG0boWTbwYG+0FPTbkww2mA8VxoZbX
tGen640Qd2SkHPbJuQxH58rQ/fZ16gauvNasrhGAZC5qdJA00uO+WdKBvjAYrqPFIpebGA1tKtzW
XKNM4jZ+NCCdRhHVqbHJgbgh7XA4JxvK4vSC8ke1wbT0nbRPu+AZpgC2TAQzJYz/fG4Lpw+g2bcO
vn9c0BCMpgwlmk9MGUG8ETFl3SqczSWlIZu3dBSTm7f3UWdAl3+uhcZm7+6PMMwGVY2GjbfXD6T/
xNdUPkjpVFqfdn+qGmBgC+2qn8gb0d1jjzP0EOiDJCqFWV9lyDJ9kzCXIibODCJl7riY0mclT/9Z
HCyvplmQwlRfxr6nkN6WfRjBORRleK8b73P8NCN/0FIuECo9dYGpf8mYQW9PVwlkaRyInfkWUBHv
qVb5chMMUsTlTqB3/o8ib9hmTfhFLO8jthpx4MG2e/Fp7bfTxoXFgaCHOuuPUp9yy1a3+9EMdnMi
PFoGspCrbtr6on1av6McsVsqqhj8GuFuo2nV11lkBAdo4D8XitJ9OC595mY+hKF7WrWT3R3t9ERT
P3zZnfdwMFsWrlhLYQNWgsgMx33qVukdOpKeFj5zwiq0EORjV/W5yx5YR21zBhQ8i8Vdghdk3mWB
kG+TX+MwVlpkGHDCbaP+6Cv4+3qhtrUgm0QMS2/zVJ8sW6Pz+gdXv+7uVpFnFWXsaeZGcIkKjFe2
yxsXYiGKrQYsRiuQU8VDmhT0r1/Q73Qhp52yzypFwQopz9db3BgRWmpvgtRiGvrN7Ak7D6D1gqJZ
YRHWd/37REbjGMzcpyZEfHtaOqEKHFvLdNoQly3xFLyIC1IyKlhK2oZdZ4P1trv1ta8n6QMaZIId
ltQc/3srT6w78uaEIGlJpu9vIKXWHk+hagRsDfx4sNYW2K8Glt22KIRnmk9LcEv9TRpmYxcppgj7
RS0CMb50+n8tQEIfNCHBdVk+VqVwa4RnpQCZ3NVIGESdWiBNs4V7/sqxSBYy/7tIH1UtBp1vrSAK
No4ce/N099Jiei+nhsFQZic2RLzBg3QnSsebJSvkPIABHgBmh2gL5kU/roibKmT+D3vlfsSIvsOg
KydPJM0k/REgGLietCsRW+FYF5+OuXCa7M5NayxKYdRJuEpqhE5ZOSqojmVEIxW6r3qyP5yHnHlD
86mhG2+AAO+N7UwBZ6utqOiU3lJnv3lGAFno4nyGXfecRMPiNrzymxikSUvv5lA4/PxkON9r4dwH
i2qsw0tYrIGKt/TNd3tCtkHyfYVZ++KL1i13fDlsWIuzBtJfqFn8qpL7YmkzmzdFbto/uzvyHYsK
ra/3udTQi7vHJXMbC40aKUixIORi2f9kJns2/hagOXh/eHjHExTE0pVwJKV20hHNumEd7Ysr4Csg
rDKpResBvuilJWPwVtqvql3grt0OPj68CUquztiOqYWgA1j3RTpjchiwE7IblMzy2Nr2pT0nZBkZ
JCmmuSwTZqto8VZFOmBNNP/RH7w2Blr5teCUT9FOIqfsIIqTxcvrSklMyqhhjDHOjVzRfPnHZOs6
qpvErTrxizxN3oeUqeApkZLuUJqaBqqt0PC+l0zEehmK3QfyVRFEHH5xInCAoZWC+y2H8icJTB7N
SpvJ/j4JezHevkLNwn5JvLPOw82NrS50hQqZyJ4xuJVagQdKhLgUKk/fuN0L2ZNBmhZW6/nW+QvR
zrmtDembw3M/AnecjxYR8NduVsHRSjWHeiO7qQY5uQfHbdxz5IIv5cYDm9uzBQa/JlnC3lN2hXwy
MqAtIJ3W2TIz5EXT/Ab/HO5wuH5ZwqcNLGgM9NSsbqT/J9UUmTdIQl6twetS3Ig+rJQzA8zFfEwu
2Hu+ss+7xV42ZmrlUZXeJDAf+PbO3eJaNeHdiaWMnrxMDziXtZuAa8I2F/AJLfT9cbce5tz5XNUj
qnIW46Kc2/dSn/gCcVVmajqwwhLm4LjfYTueCQg88A+K4k3bBJHw2ezsySCJuV6NhIP308JUYGkZ
mZ/ftP7oQhpAuGXIO9REh1ZkXsPnTn8+zN77rZwhdPx/IZlkSE/QhQ2BzlaPRdHuZger+6dZxD5G
m67usrpiSVRuJ0iLxG3q7lM16w7Jdz78d7bGGwx3aGdkcigY7TGhyTbo5oh3LxDzpaidCU3sxXV+
vpvTr/FqNUvhF3ITE7ifuq5FwqiI5mooxWYm0HlFEpDLMoMEK+o2Ux+M1gaJT2OjoH2/KC85wrH7
RloZuoqj8xq6B0j5bdhnUlwFxsTtVPSYlOEwvUORE/6OSHjuyXWSJSqsjCNU7eK0TYCUcslfCo4d
iegSA/NVpMjhauBGjqTtCVhCBwZGlzQ4E2PjR7AS1A7ZhgZmFjkZ6twxymQWlkYH61jkg17D/+AE
kBQnHS2oC4rZiDTu2s2A9QISCcQCQogNfIpgcahTYx9ZePQQIpdcbBQFv5TvNoXZcYwh1RzhsUhM
0ankUNg7gkH8KUwiIdIta1yaXsVy3EbuvyzsxB0cf1bHxLAcaQPeG6CJ8RYLkpMPZlZLW6l+/yaM
VJCyAUKkdH6IB6LrzaEsE2IW9dEUfx3TwGCaUQR25NSp+mPdpPAFa/Wx4Hfv95iFEzKpehwE4Wt6
nyq0RfENpx2XZZVVTll7wjcUrhGN9ugKTBavbS5Ks1wLI+sq2/14FJTe18PwK3XLMfzSm7EEaC6R
ObsT3FPt+nkKY5v3dnTP5dTeojRlYP25sZRcjob7tkrpr5eT/pR39W0Yf2s8Wz7vzJewqe/kXvA/
3V5v39a1fkI5ps1+mGLuQvwsXAV4ePePF95Z9/NzSPMvbTJ5KH6NaOqZKIfo9sYZyP0ZrmhcCYe5
wFlIfRAHZlIDi6mfthiboQV8Sg6W3ycDJPUV0j4bZkNmUxNVCS4en9NzgmY3tQpDXwRVbqCHqKRf
xYAuNW6CBhsrraOnOBWzaC9UZpwCBty4Wt3TliDO3rl/dVGFlLu6kLwaSrivNEVH4/XoPaWYhj/3
dqpdhKqQxojbMm6uuQXJMf5+Rz3gvbMt80erKFWk+5SThYUQkqfLZnHV7Q1b15Bik7KMk5GfWp9D
omgO7S56a0QPjfMH2MG3gdnfWP7hz4npoS7PFyUKI0O3wpOUqnk0OEWE7EGIuqiCFb+u/iGHe1hy
BO7PG1pDZhXfloSAR+sG966oNEiL1kLWnnjSpR5TEHDeKn+K8glLW3p7M+hB74drzthyjjIu8yev
RzVGoMeBA7qtA1dMp7+2S3YIe72O+J/B4v7awdQXTFgB4qgVFtfwk6A1pGJkOA46u6h/1xMfNtn0
aWU7oZrtMC2jJBC4kZdP7TJUmejvzLJw7egZ1sh1Fw+O/Npc2zL587pj/xrenVcMc4AfMAFYWSNU
OBwjdXHtAiTj6LQuN12Fw4MGIb+u+q6wk6OVq27E5yyUhnn3rK09IaSYeW2LzaAHdW9pj6+6WEch
Sw58GtH6DXTPgZfegZ6HtS7cUdMKIDXG0jmWY/aWz8/O00OWZMnPPKsqZIyZcRG7Zaf/ARQso7/b
w/mW4/hp0l9BCHeJxzTq72kltXuOhPwIXkinJ+Skz73bIJuhybUyD/i1Ief1ETQ21LVhMdUWH1Ei
bNrHSWdpskIwreMuovBfhQBk3ljysH+Rkg7oZtiChJ+3/cC8M+blPKIcNb133ehYt9BNsdv8V6+Q
AkGowsKWgW5NEA5glK50MVSLs1mvPLfMZ7YU4aS1inn+680Ib87vR4/ZohXnP2Zvm7qDVRAhtL8U
V9IzJMxuuC6sw/HpWNFMZ1TmaKxtQu8jZg3Q7Xcb9M2U+Qgtyw/H/wxladjwSftN4dxXJ7yHoCFH
I2YoKI0OxfTP4/Ql6FdXHvK6J8bnjjsJweNitePzGglsCi65SAgYXlCuWaIZUPx35wZfftFpOWhR
dRDefbYV9+4+vRSoxvQcpyzP3SHmkTT/GDK7JO9mSOggolLkXVTtVHeEs+278Jc1VH6mXdrj/rGg
+YryNYgf+bun0s5u+cFwl+RStky3s2Lp8WAtIW7HnND00Oaexb5LnOappdek341WSIH52BkVGO8K
m6gvW5ojZ7JGInXZzFhx3ljuVq5q3piiJwjmeKO1emmlltsVH+8CHa+UAW7S2b6rfrCshIf+m84Y
YqnbuFkbQ8EuvDyAd139AZYrm7g3wT9bJk3LhkubWziIpm+HMx3fqfSBYTzaCnJe7hdCsUUQl0NM
pT5h3Jh+tQpBsecbULtvXSMBV38sHb83YFtdB0D5Jlbpu+J6OQjfDNt1dADtdTGStON2CZaoEZex
5yNmsZ2ATDjuH0m/5vqz/zmco5H+QUmhpTn/sS0Fg7qWA1fLtTO1+baTfAbw/Vd5vpDQb6ue4Ocg
4Q4+bRfGDh9pORI+e3uGap7G7DGtkWFNsk+ymdaOIYiww6a9wLHtREmSFPuuOad2djEkLUA1N022
+ngjXakY3aogjS3aBwclYI0mEvnys8rnEAGzp8XhmCBpYqDFDIt3X1xqtc6mwHcfMYe+Ja/Wlg+0
sdj+zThApXOu2mr5AB4CF1q+iIDy331LL9a1M2Hj03ZPEIIlWnMnkE1lx+YY3WmynxrTqnvr/jh1
6aU54XArqeNY9PVNbK9UR1fsFbsYm6rF2nScQxX1O43fhNdP/OHUX6oNSyNhFZVfg2gGiz9dpN1B
8lo2al8qBBfMJWZ6j8/Mw03qfwP+4Nc+lJGEnukTkQF4LFabrJTH1LyPhlyyqlihhwQcignP/dgM
MvYAniSmayvS5aB8lpFrLPs3ROq19z1H1yTAUs7Fh7Fiao3Fbj/u2W3r8SvAhqCES/WGAlSkO9E7
RlYv+pXWRsj9y4aL4aFOEdn4wVUUAdOtb+s81D3d2E/gy+4OGuQzwahBg/ZkOg+ew7WIHcVmPXi0
bt5y3bieIUNDOfpsYzrxrIfBR8AwgxLuzdSvZGwN155MmAqQ/PLwOtGIb//Pj6/4V1EVNS2pAyZV
QEkRmuE9lLfMhTQC3ryicurpkvThq1cSGZHQha8KrAZ+aCC8aLmUH9+F7EjdDt8zgaMCQ30/17au
6jyB4+fIOJFGWgZxZKAWckSKcA4d0axHAGgKQUMf5NoGf/PQH8fq2C7BxANHN+V+WoTgie/qB/me
lLJYsG+eA5FqdoYmX/IH86D05sQF4NSEmdvXknzKvgNJlhoVY1i5UewLzKuyBpI5cFx+pE0Qv6mK
8qbfUTUFbj6utyvfCNbl52ivFvC/LsrMTi0fOg7y4uPEsHvSZxZzV76yuchqxYhR8TT2B/KFxyhy
smXE880344YUNFJ1HiD895v6G4EKiuygzxrb/SPsAFhIgXGn1d6tVDo18unF5QFUcUQcBS88v9MR
SiFb5W2zEJklKgDqcA4lkIEMngdGBHfqD+mGkJplLFx4z6xelEPl3CCaLLK809hBx9C1Xc8Kbpz5
MB5lhwju2CTePRwrsVd/kn0ffrkX/wzExSxXgxH+HLUhGi8ZmQhVqizHYnIkp0wGXS4VGYADu6Jp
NRzh4g5Tarf3n8d4ihNKqullvVpLv8rkIATB4hMOvAizF0kAAfS3veMHg6+BNohmBYX75STzrnEz
bXgP/WHVexxWMX6RG2bNbQxsbqX9eREja5Bb9uOsKx/PIzJwY1k2WxoQ9yYX5z/AX7xsiEnaGitC
680vgDHkdL4M0ONxuPoLCGUTExjxDTZie7MEzSS921J1vQX0WwRNw8SFBEKoGTztMWChzqDlX5rF
7PpSDayQILHdjUNac4oDO1htv5247XyIcjdNL02brBR7P4TznFtSeNR0Ah+PQJtqrMGDAyA5/85w
oZtDOda2A5EnmIK0r+BzX1PvzsLIjxhA5jaBQEIAxGvz5rx7207RFc7p8rwqSVpn5uFI+IXSm5ew
JTSOXfNJTFVietDINrYaoGrnevKf2/Qk6x+GL/m7avrNeat0nt03ZLTgFdVJinmvJiI9/z1tQFVQ
0PBosHrgtDLDA6ep76wDjYgRF+cNSjedQQHu/ctE/9S+HUZ+Wdqj2ty2cnGVJrT36Av0+0ZW3QSG
b8pxKplVtFBq+LTSDhfNsFpVpJG/PmMj2m6SeFSQVCwW2ArGvxpnbxH10qrHedQnoq2B3gjyWLOr
N9QnAVJ7EZhQWhf99mlWKscIpCEKcDTQZTl3KPIRzZrIAAvAbq1hoBZuMuldRzoxtB9jdlPpG0hm
CGTh3hpRGhj+9WkoQIkvmmJ+osT7ynUQ2dgn/Kb42t8uRdd/VDQBFZyzi9l1O5lLdgyjLE57ALjR
vSdyzwRiqgG9FByr5oj4UFpKevgBYaL7ksMHXUHYxmf2tnpqic9DZ5noZ+uR6oq6myU2PJUpovL3
GhHQTYTkjzsECoE0wEUpHyLw7sIvNk3oZNgY8YCBwV23fgQIH+OOirbzk3DKcU7lcOQzReQyOZy1
pOXxKAsb1Tuo0mdNT/EE3H/GGnsvMtNmZzUGguyXL1HUCp+dJPQ1DL3g65hgaassag4iXMtimqPB
4aSimXUZAUEBa8WNGPNDz/ysZdu1IxRkk5A++b+/0DaQSzsXbX91OsvqSIYKlGOR1ShVipZFxNBz
kvCXO9HBsa9opprvEuWue1PHc/1IR1V5CraIfUK6KlURyY0Mg0lN/x5plq5VbAzNBCWlyvOp43UE
Qm8pJGhkefCSyjbv6q3Lo0XJGXwh4eu/hkV9v6S8GjFV35mj0BvFDKb9e9rKgj5+piq+8sZp8Dkr
UYA+k0COlFnrw7Mhu42bT6IwH+H0z86dU/6cSx7yL6i5bAeSx2iDZ0UCtp2iOIoOoIb1jUgRJrKS
2WWl1VV73ONk3gC6xeXOlVeHosOrm7lpC6L20U+D6hPVE1XGNpmJcPqT+ZMGLCkbVinXfOEjgTf+
hH7UlkONLSv1gRB3H0OKxB1igh1FhnDFGiGPEvd3h5Auq2D4z0asJxKHn3gZqEvMwrm7tJOarPhg
noucQInAQ9SGPcKUNMy42BgtAM6i/tk0xjZ5xLGi/XDZdRLZepmpV+FnY/HXiqO45WHIQvyQPYl2
tcEM3tav93XZr8AYblCtE6IIBWA1kP15MksZqy9MnLsY6M77uVnrS1QUvC7nKA7+qutvwhBq5xrn
sNJn1i+jCCJ8stD5/vzzhRrMt7ayIJOSo3tfUpNRon7kpq11IqVAl02xeYX8y8ZwCSx9fo6rtU7z
mbipHNuo9eYZ4gckm42aqS5KpOQSvcXs5aZuEuT+HPX7YHzcryq8P9ZYTAt1KpgNe6TcTB5kg60E
SZ/olst3ejQ8tVXBQuWiqXAGdbBKTB8gw6aYZCBg/fCpfaI4R+sI8hRPG6nyXMXiiPOFCqxDzHMY
0bfoOY300zE/9YbqpT6glrAE3yDvFzlG09cDWuqiwF/SuniAKLWp0ryPw9eDjqlLJwlKNA/dRMXx
P+B+N7lkJj8T3rin+74a0HHtiNuBJ/ZPWTGCQFLD1BRalxEWfBAMiOKmUG+QtaXqLHHZk3lIhrYf
tmrx4up7/Tqj4VZVMbssXEQoUI/phJEjMpUrNywa4UbAdsOfYs80Sd5NWfP8St4GFxnDv+DLAlC3
5g4ZkG1K7CKwZ2KzJCxRS5gTABeJePy8+T/Zs0Em9Z5XZ9fVPcoon6ZX58S3vqemVsser/VJtV8k
czJw3By7D5BBZNLtwZQSDklFfRVq3p73uXREw7dvEWn/1991QCvh0ncOXcrzED9T5/G605p+VWSb
kXIs1tYA65AwrZpidHcGIq9FaWtYnApjuELhUQcKWM5xgCdkFO6yNcBkwtz/WNYKmaeDo3G8wsNL
QE9uxH8bL4BzPXYdyj/DvGhUoV7r6zyCFRlcStM8QykMAxkx7jNCcwfqnSHpp6h0R4PF/26JQtAU
FRFZNb7jah/NT1eTX1u0UUFxekvj7t/bTw4krlbLIB/q01X1AdumtWanyCDF2RtrUoZ4gcy+aKPv
q/t+4vm87cmrVLhrRanqZXQUu1m/jGy3MIpiSzi/ZWRxCxQvsipL7uEWuCt3ZyH7+uKjqzRWeWmb
ETk/P6soiaIm2qIEn5jmBQQA1OI6j7EKpBzlLXWmWMP/SJWf5Y33LGZ1CORXD1l/iuTiCbEWnm4E
e8f3ubBu9CHC+vKuRVGYaVJ6Po0XHQGh6dItwIa2wTd9l6KFFvMX2XnZe9s/o2N9pDBs5VN4l2jy
fNdjUkrEyDXSZLO7Vfvd5keu8b4QbFQnjEjVEWgtzQ4xjKLL+/QtHjkYrqhBC7/JuDvttzSMiUOc
qkfjqOGXw+cI+UTelcQz2vduYvi0BjUSi+rcf7KRDasWDb3ZQWvWUveT23U9xhVZEzO6vEyWZKz/
nNoW9fv3sWeF0hHZTr/JvT6MRBM0sNJmi/0HpVIv84hUWTTI+Etw6E1CBRZCROqGOg2HXFXH9Wrl
QlhW6SnxxnxironO0GRSzfnfnc5QN8mDUa6RjTjEiWXWX0VatuQNIE/iYlrJ/rbNBVEuWQb0iySR
+s4oA1sc2xyk77TrCmjTYztNKaYMSnCVHcglgCUvp/fh4Sz3jN85CbyQ4v+s3btfbxhtWpurlAHy
Utoq1EI8wj2XWWk69tilc2N9FYLueL/hAwfbGqzw0x6AclxkOIC6OWzyybooUzYWb7zM0OvE9aBs
u4LoYJ8a+Zd5Rcgk7qgyPvhlE7WZrLDpRQQVIIZwEvneOrIPwRH1rJi3aLdx8ISBhjLuk2kgny27
e8b9vZgH75/jAbOqKiAqX6HWdQ7SwEcfoTNHEF42UWfP3vrl9Zh07CnxyMS3JZ3YOL/pxfYCyelw
ulXEQjRoMjSqs6mgxbsVWKwTIJQD4dTxexZ9GIL9MTefpEONH+9PRJPVrZua+9/dG4hxs0t4jFCq
YuhRufCumrT2bcddsKgSdItFP+bCEXOLqfg9N9CQthcBAhAuW3l78089eV+5gCSHmmroR39tVwOm
MON+ywG+GrUZgg5WfdUGwegKEs1srp5USeveCZqXCBtO9zL+8y4OmgBPu9sZPM6dgdD7kQ4E+C5T
Yz6ief4mJlK/fLq1INZCQd9D9gw28kCptTr2IJR9qoaMJrjCQ+U+6xDmZuW5JavmLZn2t1Cx2OXq
lTTDYwWpojW+ew9r0eNbGX4kRijRut8sJ4RBcSq5q65q4vOaCzpB8IGj84J+G4Y9JS8zDNe0NwOy
ecSCSZSqSN+D7PZEYUhqSHATODtxSOtVpoUul9MOJ74NMZMZKSeyViHNdmSdY2dJZvu+74Gco6Ha
2fi5BHomUh7gsAa+H5MvcITaIXu4en1BblSTDB3jOFR6gYWzJTh2d3oysoAfpM5y5nr8isKo/v4s
GD0NctWAT0zYrvIhJZXoTQV1TiA+CAngPa6dLnvkUZYPm70Vw3Ge+1+nuqwU5r7yIsq40bwgX+/T
ld9IwhRnq7dyhCy+wW4ON3iz/kEEi6lNiQdnKgnLZ/WSve5QUQThHrJ3zFwSvXe44/bnjiAor12r
n0fVYgg/N5KKaaD61o3xNFkPlhNN+2mBEJTblRmNQNX66N3hpMgvI8xq64w8WS2kitOMiyBbJb/n
v27m5BSxOkShAKycxezPtF4u8BMDiVXa1smINorYiQD8w+DGX5eeAJzoZYgTB11ZoT0FFRYd/U8U
B0bOqbMyMdq3nrDRxi/pcTgRWAKl3qdJzBFkT3RatiUg7/PMy+e0PDciEBUYlAPiI+r1u/D5D4Xs
FHGAqTaDLFv96bL7z4fmetfX4vh6J4D66mEPxIFmXur3hlGsUDy7PsZwmeRl/FUlV6f2gtQsjgq6
8oMkHXEr4pliQVvp/UC8pgSeFcOuZ7Y6c7BiIe9nSAYiZst9qRMkH1GriKPPh7+FKn/YsCVVUzq0
xKKx3mtkeTreUvwPLB2AZn/FD9YWig/wTB2itIhZR86AocA8YDPRbAbYPADxB/H2fL7tsmi8HdP2
eYu6972y2Vl5fGg+sFoXRO2V4e+7KovhOKxQnJsN+PpxbS76J8hWoyaEoCG8CxifE7cKksAbNpkq
Z86R3tgQCR7q2lwzj/GZ6wo8RpszlnuToinUSoM9c4RakxsQfKO/j2Rvvw0S9vWMnpxWJG5eNBwA
eDfS9iKdEMgBDm92EUf8ghbo4KuJ5FJoXqzlDAmubWBHu4+Hsshug5MqaICBdvCv1BHs0msIwm+h
e4KT91JrgUcuecHIeFLeUpu0pLYFNt8ISkIYkI96NDeupgfz64/vVyURp6SDMjbOWZ7ZARS+QdO8
KnPNyWR1svb8yOGxJ4T5OoZrKGfU5VFFR6GMEBYyVSB9m+vpTeQK0Pzd3nr/o7123ifThzcwisYT
TQgmSXXElU/j7AhPoI4rcrjNq4KzlbAxdMhFVJB0nJxwODduaVwjJd86wzuMNThhh6eL1k5+poeW
o2z2G5dpXoaiNlmCIzC09iwUwL+RQMCZjtL62R3YJaT0Tf5nBXjL51dDzBNnZvzCL/4auIMpW0rf
8DjET5xTQVEE9p27+uFnL4FjI7bMJeR3T1fKhF56NQr1RDtd36R5HRopdaF69hZs5XsMORIxRSNQ
rhnTO6D8wLyFZQ4DQUxGeDnimmR0nqIh5gMOCvvDCoWJnbhStrsWNwBSjPsr3+iidiv5nmkR3KQi
4ypUFhmJ6lDCU0yxxHBXKB8h1EWK618z3fEyal2RqE86xnY9szixNHmQcD7LFhwuwJxth9DXz1Au
Y8S4xHqCq3+4ItraFp4HTcELYbsfwehDLg/MqqWxWv62snhnCiQ5yudCw4wwoUuT/HnvxD1q96LE
MRyC7YGtFhiEidCuNF2275/P191pQP5DXmp6mKnZPb6aW0BRR+X3x4nr3IUY2dyItSth11sPkBYs
02lGrRvYth0gbYVxX9oh2aK7nuHWhE0ydSq2eKNDVuRvGfeUFsBxfo3R8jY2rzCSL2OhlqzWggsS
n801VnTXNxNbmTu6d0h+/6IUDSfER2J8+k92YuOK2ZlnFsMQZ5dkK8UTZd3N4QccjdbnTDmRb6WM
63Ic7PgVVB9abClihCGJtKI6F1FVITo1VWZPgeJwYhvCoZtwi0ceMG7/pQU0nexhND2yA/iIUPE5
MqO7QFw91cU3TnJyH6H+LJ/vScr/hMzqCkCX5+9jc7keJ/E3ZorKW5LOojeC6RGjxT8t9COedTXs
ZNKOXYbD3x9FMh6iG5PoQ+XLTmrBZWXfYi3B1DD7U9YxWhIl4NGWzkf6PDZJ9HrCTr/mdiXDqNa/
sKVyqxc0qGNQsh63tyeOiW9NaRVDSmYm0PxPbomrf+0vNFbnz1/eGkZskDE8bbzjPyBUFr5Qz4FM
2/FU0ITV+Kf8ukIKoj+iS6x1MS1gGZiHSDTCLUG7qttBcgNPd8KZek/kbDVdlOb4+XkHvH91nTU0
tBee5NN8UDh48DAtXDe8udODYzo4q3FYm4GLDpaIiDbBT96TQRlqhCg7m+xr9XQ5UKscKeaCrFIZ
uMQRKiG09EsdlSpfA/i8NMPs3EB4d/IVgPFKIPd2KQkCeC8u1otymagHvCJDkeA7Z3G/Jeykaylf
j+ahxaSm7XZXdIrJNWlJnjbPG+p8QkhuGvh9qksKq4YQj2Iyk8hTVOneBGrQOMvUENAWPwy47hzv
xa0mh16Rh7aNTPjDB42BuXN3VHaDYB6+gq/gzWusfamqabVxyx1XmFaGKArvQG6kD0glBlf/LDgc
V/3QVKsI4VTBudhlslVfu9hYW7Bk2tjL6c3G2ub5LaP7H5OfTrP7XVu+Bj8fVKb9EjJUkAg6R6V2
Y43fjV/ZU59iHmbumbm+41yuxLcri1+lMfY2/BeCIzkfbNkM2jew+kxzrVE8QZ/SkY1A6/XE0p5c
3NtioQ1IKL4+BIS0fc2jx22oXFwLSL6Uv+Dwi/RG54ATfkd7tBcm1JzXUqgKCHxR6ppPMMv7xKka
BHY/C/0U/1vMHfVwdXsd5D2MzsxabwW7K4LRDahcshXhdeCP5N4GWTyXqOCbI8vO94NB/xRdx9ES
RXXLr5lwaIZuMeg66gPzk+DyIBt+28d9v8FCmaG/FXcZCY8UJp50PAD+KcbbB9cRuaBQ31LzF0CE
ZvAyK6D/GNiFgTr/xS3Uc4hCM1rDo1Zbbx1QbEGjGifYOt/k5ISNaUj0Ll9AF6cZxwL73E2No8WF
reujeDp9ELitQho/WI2igTh8E4XLzTxMPI6d/d2XlcnNsKiH3dmsCRN3dX0eDqFYuZY/XMOPyJ2E
ruHmDYfZ4/ChHQl2OmNRKbYd8qMDKl0dwjdmY4K9svg4/KwCw4ypZQSxkpdXam3WdsCdnEuaFAZQ
wXr0/YlZJMadwvMv6+8YTK489ZE8uwi37TCx448cZCh3iWD6VKG1m5lFr37S1AkfjHqyqV1NelbN
zNOo1ogkS5lWHVg2Ni5c4lERvmMzy/ZHmhu4SNCOmrkvKCafZX3N91p1tBz7rac7YFH7nmmrE77c
Idnb4jWrBsjp/Wly3Cuo9+olLwNALiBhr8sxfOPCiKjLIp2I88bVNz3+RJxqVHtoIlCrmvlRy5tr
jN7IHjUA6ZRqfw9Mtg51LmxGYN0obyM5nmZMTni2bhyjyNaRArhSPIDf+u4SICSuG02L4kMRO7F/
O+3riCaTOBcvhce6eX3MFwZMXjBvjYDe/CatQE1K2CmbDfyhMFmJCYXkt8/U4MGagmyn7D+LMudb
WT+QwJbDXVk5sYoRsj+ceA/3EeTKbyXwLO0ScbrR6J8QpENm2kQbqxUr/JVdsUl0bR8ThQwrV2LV
WX3wlkQiJIhi30B5akTCU4ZY2v0binqInt6s4DGFU5nQatPof6JhMuLoPr7yZSmIkazB8yVszycb
QKhBhkL2Gz0uxRKhLQh0yobM4lP0Pv/xHkuqQMBxrHsAfKQWXvnPyAzxcB/dM/+M6nx8m6irpLLe
itDqZNvBoO29Hje44Z9wONT+FEl+3CE9KyNNATH4z2XK2bZ1irUweoKJjvpo4O28mWZhBQZRCcqg
Akt/feutoqv0Og3xDApN9GF0fplbkIrFBaZFzH+nFZGtY53gr2CNUK5O6AZi0RgC7FMxtmsWQ3Fj
3W2BOHyQ78POv0lx2i2ketfInQqWzdEu9MZKFFmkathqqeL5a99WnTu8SUimv64UrPFsHBBhQjBw
3VJWbYhrxyHZ0MRmKmYyOXhT8L37l0IsAm6u1CinL92cihcX+XJJ2HLR+vbAKMzTeUIfcuH2wXQD
ScHAAnihl+yPlA2NcqtO6ZNV5vdXAld4viojAJuFkI7x6fz3sQafNQbODFY2KX/kV0Qt1X5Tlues
DXh+QuOkL/ckE/wRjhP+oycujJrBcnE4+mbAmRpwx45o33JulFk4Wsv4FDOnbxzwE2F3tkIDvON2
IXKAs5AOCml54zr/G2VHvXAojXtHWiEkyS4LQJzr/ONgQPqk0I3ObV6ZbqGwwNI/SQTt8KeavP4B
LqsO6E0l6o0Z7SBnv8/kUvA42woc5PMgcCEIzAJ/BttSVOFsRQIQA5OeeHHkN7Zw/n8SzvvbPqMW
tiI3o+Am0A7zVxVnMXcQLd+eq91cL/WBlzobwANfQbblY3clHbHHb8xHRzXVyfebt3M/8f9AJJb5
7E1H+WGRLRPuFEzv7dR+y/IuEMedxBDj7gW6C2LBJwac4Gpi99HjwsMXokTNwkG6aH0SpS4upKEz
exFMm7K5NoMx/8wxyDkvh2vv7APQ5BeuFH2nYVO2LxGT4Q7qdUrO9iuBufVvZZlVI8gLuG2FjzPQ
fmpRBFK5ElJ77XgSEpe8lzIgyJLi+1RTK9B02tYTyoMPsi9Qc9RT9VP9Ju7x0olxijLS8Yu1tXnx
2HF7OJEfY1nzMst4r5B8oJAuhDSZWwf8NOIabrxVVGbR4k2ZbS/yR8Ri7XjjvamNzzaWFVyYo+7G
/Dsz1l0EdzIf7TLq7MKKY+rQaUxYh9/mUTwbtJJeyu6rEVXU/2DPZUPO2S/1zBmq6b5f34gaEsnC
NBMDUDIIyeXkNAXspZdKsjcKZfAAA6gzoH4iXloIW762yCXdPnrZlOjBE7t5ZI4hBH9cgzHirS1/
2POHwZtA8Yb9+Gbg41J8Ix6nrDlzPKA0dpOvG/gKMrsC7m/bwIEzk0D8HytNVyKCL6qGw3ahw1n8
cHUNN/e1GMOrtjZLEGKfQ6ArANPXuInjEhSBWqO4EWQN45m9sJNHn/z9D80BjObIwKJsll3Nb6H5
P/OhS4l4+Gw4qLC1Vd1aoNX53KxoG7GsCKHMs23HB4XmpXhxxUe+jG7hx74yPvClKU/JBabJe7tq
fnV7mNnzPXDRRsSGFKVG+zKJ5d389V1eJrUtTdd05rY3l2O6zJF22VF5GhoL4Rn2uTGfTokGVitY
aGIXtJidAhWaHOIccOjrXlwZS09noOIU6GZaXVzcFT8+TPRu9vNaU8pP8aTGSRt8ycOq+BuU92ik
fjAM4OyXMZMl0IHVBrTnpuqoA80hO/JfYM5AdfcPSLYEk90M44ZolH14ygmtiZPOZVb6CLEvcX0O
4G8/ZL5ElkVZTC9wjx3xB7z6MwW55zLQyEaXoKqBpf2wdrDlmvT3sqLirKiEC+N5mW9Si4tisC1y
2aI0Fiw0SBIXocNzlH5Y9pkD4vt8MJ9knWhEvGyA4vjrwhFDkBgMwu8thfc6T+6BVgAdJl1SwqRz
jqVimkpZ/BEdrskZcNNtFKAKyrYaQqtkdiHJEK3wuPqqcL6BwQnXiED1Vppu0W1s/wPxrf7mqgVM
KtVEWayfdSY4thN7s7c1L2hDqyapouiXCgrfeJyf1oyy49hTKFPPuI8kzRQwGZ/WOKOtrsy46R+d
2kWa9cWSWc1YgeXOfE5lBO8F3MTgpiGYiMBq53siTPCHMUmsLRvCi0F18t+N2gWPBQRMaMsyeiZF
jloyndxhej7hPK40S6IN6WmWtVDh3euDFv28nYRQfOhESkXgmvf1pBb3nq1+FAIHXe1DnZPRFWxm
H+HljsC4NdvNgnhC5+HVgofxinczZ+xLF0gkY31wcb1yYvg2v1tZXQTjcvHoX5oUiJ0APHlLECIR
u/o5Wc3DwSP8YVJJW7wyW7JT36SgkyVa3Sqvduj9k9C8Vk1dv0WQrJTDTv8uJMn9vk+BPH0bF0Zw
jp0al+6uduRY4LPWRbQmlOLYNVP3iWpb/pmNR55HeISCtZ5mnmffkFG75otguSZF1DjabJqexeEU
1wGzryJzSixjJSBRc4b+3kXtbnq0wcK3GcfFMbRcCQNx+bRHot+vxZfIzypRCe9IRlb3oOhIYtE/
Xxo8kIJBvcxfXfWRwgjQWDgR9uafEP0aQciQaxE9ByE4z0cLo4C1EBrKy7ofg46l72ODuW5bb81T
/qYhK33ozICt/+iC4sS3KnaIFJAW2T55DuSZkllNq4uPwwx/6C4nTGvypO0gTXre7lzQIqkGG8RV
Int2XWjSW9THD0VeRSBy67qfpQReRklSh7aFKtEQYM2wGPf0rD5ZMx05NPRpqGo5EuXCKUslN4lr
a6aWmP2hS3wg2OZavsKkqkc1WxGmiflgl70/T0nFU+S2EQE5o3rnPuhRgh6FxCHlEabJufRa/bIQ
YngR3KfoG6730bc/SVeo34WvQmxluhLplLNxRlbZVRmGmoeof2IDCGpwqVi94BCuSoCwXPg5+vNV
y1Yvbtq2CMBCT5rIsndVpHKZJD2/ADvVyi19cR7yh2jxufwRsycIirLoeSnvvCZxx7Tf0/GAEHgm
tfVQJ6CtXUwl6oYK08tbZ9Q++XbaKj1NtmPJ2PYmxN9XWe/G5KafrGPwvou0z1HT1EOD1eMExGXf
SlTcWtn3SOjDxYyGbCGOOpY/dMLRZusUuvp4CRI+SCSo3fThGaGuZ/MnMrFAu92g1gq2mzi24Nyk
2ZRm0XPfriUANMMLcW8mg8k/DlWH9pmSE/qBcdRvZd5uDWWUhmpkfsW6S4QBwyg7PKsI+6KW+28r
xWR/72SamcZiHmZLSBEUFE/NAU4FSScNGvy4L6ITdIZjHO+oqRN8CjjVw/S5ui7KQYp7ka0cbBkO
xgBkIWikSyeRW3w44YKpd4nFqDoJsGMi0RGxLzQMbcDTFEtIq92YUXSAcltNoYPJ6Valb+eU66Jf
kGkWR8gRBiZsV36T1t9GZbUphzK963scIn42bA5cATo8pj3/c7iDrv18o9BmW4l57VtmXXxkAc+4
3hruvcS/rqPFFlcktaK8SObJ39Bf0kRi3MvaMAGHVbJO2TEx1XagRK9MDkmJjPm3tlV+/mMHj12a
FbXILpKkCk65LSrdqDxWQ2eNeuqQ50SsKpOodiUFR0sL36UbNe5tNLxDFAorrENLjP58ewLdJDjD
DV27t1BUjz4X+4QcWzpxeH3I7OiNJnlJm2r4uUV9Zdr3aS67yKX5RN6OzzF+GlPiX8XDNHbMPnKk
jGF4EHm3b0HvmKXBDbTCKV3A6ai/18wyOq4RRWu4sOJx2Df227ech7/qXdSQiAjJYGe5M4rX/aXf
rFIw0vYFbyF3CdSCXq9DoF6/eokxdK+jMDFfpcPQH1XCHq3HXL5LGciEo+Cir+7TLWyhD91MTa1m
fgjqam9YD/p1rFEFgaOOduqiwuZFLwE/213dbEmGvgZcC2HQ/vLuoKx2TQESrOM92zCcmzyoPWsz
KipX6dY39J4DrRo9cZNBp2mgKdS6A+Sq6smJbsQUd/yTiaTiI2QzBU5u9lCFAwYPbmoS+gIeW6oj
Nh1X1Zu2wby2GIxTION71vvOnMMmlGLZGiFl5DwRsZRLO81k/iPBg1BitpKr3YnffL/zB4EfYgBl
R903/BSc6Kqf3f94vkMHgltajcGB4e8EDw8iIHGK8P9YK4dnABcoLw4b/QOS0NhbjQkljgJmImmV
XinzE934i+MiF5XbP8VlntdnvvoPjYX5Sp9lry2nmXFnsLfmglwE4g7WV+sPz6e0yt+6ODvUkMCW
6mMDCtEOJUfROcrkVuI6m6g+4ThH3nRzcujMXH/veeZOOGJK/680bkQofJAnOLviktO1TSVBrFvl
b76wtdxSS4jVszmxgDwP3apOI8XeirHvakMB/dytOBLsan/KgLIO4pijXFu6E4+JwBklHlgeKBSV
Zu1Ci2cRJ0QLjSu9e9RK4GDZ64kDUjq1qvDS/T88l3rqY30dJjIXE65cBcO7kyedGTvVzeYLUDrx
t49DYWtG+0hz3IFCp/KEHzkjt/sVSqMMbnXkPW3gQKrvODXsZmn6SZ6CazyJT8hBegCYjlDrqYQ6
sR4cL9h/L7VDJISxPf98epKmzYmBQqj8kiFuZEqUVD8tJGd0LFy1etggTq/rrwjbNATBKn3XCo/j
GCbaTCFQjBKgnqT7DgmMbtLKQYbOhE9KCGXy8N8wz7GrFcNMe+HVsrpWtXR6g1L3gGvGSrH9GkCY
kh6qVXa2P9eOs8tlvXuoPzmYmnQs6W2Dm7A31mYtIVowUwyteMJVwjlgREzsVoWYTpLQpMCt2Y27
K6mFaYKr7CPU1vw3HaMbO2lBHubuitnukBOHh/28fusAIQ+LcG1BHnhejJ55m/vQegweco19WBlz
V2ptiJrzaxOdRWpOBb7/RRK4uSL4bZpaIVE2zbrHk9meqTGoWIZ+oH00j+X7nFsvTscPTNlJ/znN
uF0mcKIhFqIlB+1wHCzq5aOiE197QRxANp9NSxpIPIzi1mlcGnx1GTvTjTu56JgT1LyNU54k/xRE
76sZJDNSv9ijVKa2hdVBeZ21nvPFxdfwpUaW3qtppnHHP242W5zWW2TbM7pMg0A0CalOJ8rDahW+
Gn7+vHSGJQi7xeEFBlLppYUJFzCC6PimZQTsS1JbGuzdS1jffJsN7fkrQpZTyc9iCHz0cnbiOQXX
c0X2stZci5CizcQzAbr8LEesaw+5eQ3ijdjdCwuafwPjc7JFmoaBsmnnmhC1ABEY8amj+JbD+tgH
0EXfdCdV+mBkNKMsukf+4zTPGSWvmmegdXu2mkAoXIJgqw5IpF+re2AcH0t4/ukNUfK0MUPYMz5M
V1EYT6HS2/8D5SlduSLEnZFLTb1uuIWDDjlHEdOQgth0Qyki8RpQxXdbWF6TazIlmzJ2QxaH3+JR
mx6b4SM1Tl3JkZ51U91S+QydlNKbO+sZlnIZTgy4mCRFim4XvUGPhO42+m48UFS8iOW9h32ZVzbT
nN8mXqizk5pCGD7MLtV5u7ABv5n/BG4sJFwAxCK+n58vBTCeXpTsPSlNU0StOGo7FOyW4nKLyseq
2PYSFwMoMmK3yoabm/eeGgCz7mAvPtY0xWrmssFDJdHI7JAo9+XEq+xsQpscA1BVr1E3RwrtrfV5
z/DQH2maiYAeixNjEL5NO+ofSxPy9nwzXVX3sLHOwJC6Y1pFOmcDnwjTCLdTp1t/IaNiwtP1Q5xV
Eebuv2q6fQuJLlcngTrjoKnq79qKBl99Jz70AMZn2FNwHh8fL5tpu3tjdlEhOPwUIbD1sJ5a2iNd
BL55/GT2dq2xcS9xHOhyF7CJdXbcMeWkzrkSP0vzkDMOKGbYIPxsmAEvXuYt/0fpQFwihLUG75/Y
6Kzf6CsVi12tFHHLGba1vZ6K6q61tS+BtgW65gtNk+h1P9iZxxp+K7IUM/3xf4PquMxV6abDREU1
TSFmRa7pAdfkrXqZD/NJC78BCZbbWGEd08vxtZDMWMND73A2Ql+vtmPntMkLHSiM8GEUk7zqHAtf
YQe8dlf4KkY9V/s/5k0E/9jSUTW8XWaCoZ97K8XEf4GCLv5WiVfcT9QWkDpMGl5ktpiBJDYqwX+M
UCuE7Cw1xg8RjkOH4wJr1DRZcgZ5zfHeSaYhPqQSXG+BhwhT+yH0tqQt5HA7wDypfAuUx12VC88K
fXYzhMnG+fSIohxuvzYnSuGhAHoWo4E6+ehrQlofrBJ9GmKHz31Pg9npsa1Ixgp9XXFUkSz4L7+I
H7CzGqPsvVPW7zk+ddx8bOG+Da2kLRD/urr4pYD59/abAjnoKCJ6aZRYQvbDpLpHvQ3aAXhv0Y2A
Z+gkjC/Jj+/X/ojO1CY7TqmHTsFd55KTSisbCiLi9TtLZgzccPKC+CoG3TgTSgp5EWpH3SspRQLT
WdtiqCWDOj9CSgdZrrJIDmzA9GRHyhRvvO7XI7WFU0XxHy+/yJfl6kskXzeEKAFU15L7Ph3YeTT3
wTPLuRP/9T/co7ZavlyAeAqJBGF/Hyud0GQd1Q948K0lvkaHTR7x7cskaZ2W9C/dtafFW3Xci1Xz
skw3kxhwCfMrY7NjIwjX4FyvBrlZdK5M1n+RINtQPgACkOhwUFiV2HA6pdCuqSH6+Ww97YDsD3mn
jV0ciBGVDWqZwK6uMShhLrf737XeL9XXsG41+qo9fNV2HpwT/+c7pvhufCEQ37TAhoyswRJebye8
Y+Hlgofe9E6GJMWcMnegDRPocanusFK2PSaH8IO7ht7OybJnAEXXUXEtKjvopgUUAgsamRNNoFzH
cMScJGj35U0FicQ1ZGpJyOkP8q+M6Lkum+z2MzXxJHbT6yWV3KK7iQ2fpVI0yeiR8C2Ebsnpf8WX
y3x3406asEWXhIjQHKp+JerpzUdDoAXzJxWeI58DQ4iuq7mHlN48EwiKB33aqPxGawRI4XyDXoNU
7rb/R3nn0dwMsCoE3YPEF6tLRfnqTPVhyR6k1rOy/SIF5bnZRf0NVaTIpEsm2rW9/XGbIdIsHmZj
tZg6DAV05gO2tihHR+IXT99UDdbMXMmbb7Hq69tnDvpSQW64j1T8MNqz2nPXBBOAF5SPjAZ9nnZO
K9eOAqAtsNjAn0VNKKX12JeoKJ3+fuklnLftiC/3znctPejSxD36msIY8EfWaUAlkMEQKKE1pLCw
Q83GAdxSphdeB/M2mXfcD8b7NRPD8v5E7J9gV7Sh5eWLKcyBkkf/ECzZt3F7EiPX+z0srWlSIqXy
GyxHGzrQSmFVYIBUR6i0lkhz2Cbz9g13txILhSHmQzDZySaBQzC42mydKaYsBoGlNASuMpQDIw2M
5lyCsAE2l5VuoAPMvgY1U05ZuOh5n0DsdPQTZhpcqVHFHl9qw6BJm2GhfUUX0Yz27s5OEeXw9blS
YfVCQY5aXEj4G7zHVotammu61l43mi6UNqkDrBwgkBhWWRzJ6ZSkerNk63zvbzhK1awBY7YT2VMl
y354WQzd23+QvTs6041rNLfaqfR1ai/H+5W/O3jvJlr+Urc2rdw+HmJvgLzPPrfWAM7TPA7nsfLy
PkVowAOZ23CgNzE1ElFEqKNsj4IUv59RwqQCgEH1VTl8R++VkjyvLZBiqvq5V7ntqppAqMm6jcU2
FGVk8kqoP/thPr+hdzxB/eSTC7C7EHTO/EZJ09aWkmHDxiCcciJe2FE/bmmqfN8pcyDexxuvjti3
pBN46PKlMSRDUpdsNVBgItS43HK5VVKs4RB+dLyO6W3vG02twZVGC4GWvuVKjJczuCoN4qunMyyE
Xd/oGQDgN54a7tpW3qB+davImHK7g53PBnLX8HAKB5jT69IWrrabrcdBvHFWJJaFkeZXu+jRGTOr
vh40tnnXY/D7kfx9FnHNXAItEcnHE1b+bJQbbgZ0zixwLWrIk+R8qjA1fqH5SMXc1Skn2j4kokpx
S0/wrBqGIEY0YBdicOG5QpMID5oRuniqIN8xPDxxw8RljxmOIM4WI1uQOYgZhGGgfUneAy0ovHtG
J2kfAniRX+3iJv5o5lpUTXENPTMrbSiI8vlix22s2OK8Pyfq8e8AAeyETGRQvg+pQDqeu2KZ/pGt
F0TaYOI6nFqmtQlXxxsZxMXQ4pmjrxyuaZwsQ54W30r6tcKiBL6RFnLN15eE1RV5EqBm27gjouoA
AhQuRWUOeCAXkJjbBddj0vcgXXxfa6caC8ZNBW7zn5mCnvt/RBe8mMNJhtmj/Ovymrt3G1JAYOJ4
lQseRkzGW2s7Btr/VUkDvqdziqeaiTpOyf69/jQ1BVc+Xd5UKFUUv0Kb8EbK0ODRqv930EFwwo1m
449e5/9IbQlptxy6Lp0j1twO4M1YvAaFT2QgF2AhONSY7ENEgOl8SOlpcwIhQ4ZD6xJ8vM1pUhL+
d+Wh+aoO+5nHSac8XkudJwdCBBE6aqLhwUWIjcwMTiesc9jAhGISKJzZ1OXqBn0RsIJ7FnYeDa1l
EPgNZqXTISlKQGzoMs380rOVq5A2dYDuxqEMmioqbQd4o1jqq9xnvkFGoc1NPuegDLPH2TliBaoD
xMYXP/iolAR6p7nrHj5Y7pIue/Q4aW1GkU4yhYpaNMKYqgndbD9L2zVgVwnxZp7VYDDklhEwicHp
e5rrT2x9IzFkp/WlYELmir4Mwyo6BWLJYLG/bJtvKicCxWPSpUnrGiGFVHN9A2h+lLQqmqZ1Fdf4
XaRZkKvPh3/9eF69BltksJFR/I+4wSbthcGsmcbYVFVCQx/K8AhKNSrQ7nW3PBMBTEaV5fOHcjcH
QihPZL6+th9hxgdnhvc1X0DfB8h3PwZjal+/SjVbde2ZU6IpiWtYxxUXk9dIVbVFnsiR4MghW0Lw
IjDoy95FBkDDW3lBQpsoUwWjh1Fe4OZ2B4lPzANzZDc3gc/28LvPhI2wEwPzxjzV0TCUdhL+zlfm
tdhjSXJl4AQyW/2d6OtQMe27SrOjqLYi39hJN3cNxHs7cRIX2TtOEwWAuERXGmthU8Oa17STIDJ6
vytaeKZQFp7E1nDR9FyUrB5K1L/QUVQVvmGQNrjk3wn/fWr25K2zU2VDucGmHQL2pjIVtgPK4pMC
jG2OsnaOsfXYcyhPkTrHPtCS7oF3NdfYe7FUy1SFR/96VDu1GYPDBYxvAW+CFeQExBWhTkUffoSU
Tb+qwb/6st8VMDSrT1xL57KvSL/9YPaBDwRK8OUdEYeaoZVNlDpxYQ8FU3brnqT371n+VYAq2kMw
ZuwkLqIAkF97dIDllBVjTEPAR8Vp9Z5bLJXqUNidvyOyjVkzf44llqIuU0e9mj66eSM28F2YK4qj
0ZYRt4ccVGcaRlVK/VA5z4/7GWjIG3OhPkDiL37vqC6Bxws91C15uh8YmE2cRDDuwLm87nV2vyjZ
ByVBKbAbnohAbH/92KPhOoPWNtfNebE2ydszQSz1uJM3+4gUbdjenRLm4ZHQ1AczQUBhjyikSH/9
VzTz7kZW+MwRhZqwlsymbHwglTHX7iXaxA7mKkbp2Qyw3dlYaaIn1f7rzEUZGyPVntbxQqAIvRwQ
yVykX1NKdqiDFb+XUzh9t/LFnMjyGgPtezMa8WNWADl0x66Q/yPFHyeho0mDd8GgjoGJLpqZNaK3
rqf616vhAgMZhk0UDiLzsST7hvu30zdWX7dBeHNe9eE9rL/k0u3RsPCXFvRWKKNN5+ZTt/J0xPmq
pxyZmCQCZo6MqFD1vPnZbZ44gxwEEjfMXeABDrRwgO2EyhkxF1aXmeKRPxFwegw7DuPkv/KfvIUr
kOcHoHqyPnmW4jfcPoECBCetSaK3jhHGIUe0zjOESmM3G1CtFm7sLcWOQrSfN9W+sDXZJTtCU79y
E/3Gi1CAzJBavD+fn6xrX8MWUQvOXEPpcSDNtRdwuUZtMInbnEhYNu1+H+GBpfV+hDyLkrrn9SwW
SuwT3fXKKiWwTKwlLv7FRmcqZFu6aPUdCZji+758QVq4EGe+eahYPPqP4yQfBDfSl/zKA9DdwWGJ
b8b6Gt6Xg9SRVZAft77SjbmSaQJqFJqLU9Ppxs4Xn7FMtsvZUy8yG1svTsRAntLuruON4UUxPEp1
fzYPhgvxon68d4V6L/t0IPUaJwGjceacsuQi61EEHfdV7QDWV/8xgegbFB3/cSee/LfpJUexVlFi
3QLEGUF5CwmXfYxtObsE7ptHYQugQkYJBQ2aBJ+M4ybPW08fXycm8jkWy3EwPUeiHTX2fkQqM6U+
IYU15JEe6OZmXhh947/6xXrCuu0r16zs+23rWMxJe/PIgvsmWPP+UgjvNRGUoeG4v+GixMMGIF5t
7E38rXIc5iRBdb+oqzD5WM4JjySohh8kCDuelEsecRqdi8tqlC12scaN2EbWYfejVJWMakxJS09h
2362umGmYIBXqC2B+CWstJMZd1z/+OeKhoZLYQ6TFCkixGdQlA9CLY66Zzevri4mZpzAWwJZXf9n
1DhIvKROfrp55OaV63dnepmPIt9STyp/hEl5eIKfqQObHHZoiRqXQEWnjPLV1TIPxKt26e9Qr8rR
2FU7aOa1RwxEZZpkirqCTZdwBJfOsct2yOnpu1Qnfx0yYg9NfqwJlljl9ej6McYisIrS/Q5e/o3x
5VLJbxwGOLY0aBR1Sj1yPA5j9ZlVHEF/K4AOsuHxeRPSlNwmbPGmKAl7P7BWYhUVKokCL9DWHEXu
6t2HrkXB+ewfiuh37ibiy2u6omJaP9YgH9l8eSHeGc4yJyIW7yauh44hp39ZCz/+zBohbJP22+t6
36j8Zicha24hb2JMcDN5xAtXXk4OwY5HFrttTPhmlstRSGGnGRH2NOMYvIn64RkmzjWckwotc3Jx
0pKSSeqAKC/I5bHupRRHNPhuxcAiL0MIF7YCzXTj6xegytIdfCEV008Jgi2VGugs+ssgEEzX3p/D
ZXF0Mqha1Xn4tJX/vOcJMccRDD7g1G9E08njNe6WRhigEs63ZuPTd2pJtaZhPpld4tOP4/7CU9DA
Jy9oyT4DNN9RMSzAFrqbERfE96BoTIlZRBYxFPEOyEz/a5i4H3m5Pyz3203MWVFWc6esQsYrjtMg
Gyt+fkbRZAv//kYPaTrAtk3lrYCgdI/eADmhkn8jg5eC67Y0uyit+flDXaCMfFQH+lpocBDZWW+o
XOwGyCbdSefe48USru0YFmAGQ/ii0GFPqafaqRICsOTfX55A6inxbEHHGB6++ZWUhbBUcng+MhwO
spZiuFoEN5OxScKoMMdoCWefF4vzeHlld4ABr4DeXkyNqdedAXgJ911e4sIKN5Xb7NRXmPURh+UQ
Wa1/E0T23WBvmM+1KZQeTWcWhhSq8lOoo6ZQi08v4TzIoRofY3kVfB9i2orLcmURDC4IkT7+ZvHN
TeXAwpXSWaXYdSPOBTyeg53RmXVrthjTsklbWyXC1phiPQHAgH8UjNZO7gifkdy2fg9QwKefkkeq
JqGSFTx06+tRqQYlr9S+8CCW3kyng9CDfqjCDMF/W/Ra2Tpf46Lio+sIQfchsO2dJ4C9BMljfCeW
gi6EPvUzik76hsT2rmDE1lSAGXDg1JSkJEY1gHho/yOK3EZtD22dFp8ejW0uWv1/ehQcMh1e9kAT
p3/6Y0NeL3H/KCZEoLsgqllfCi/qDIoyVIDlWCo0dEPlFstDfOggK11dhxOeJgqzXvCtK+PIx6cA
D3szvYJzZJkei7UdS9q3neXcuYALV8pGGdhkJLWxkIRuKUhX9V9IuvEeaCdG4KOBSbFARo84PdSD
lMlxilfM/csII9u3UCFtB3CtSoIJlL1j5HMDyuPH1VBhqJzzdVd2RrJf7xzEnFAdWXNQRszojsph
D2RipuVxg/mO82DzbRu4izHiG5ZaZ961BY/4FAyz5SifapI5yxtZn2l3lAfz0MONg5wUiRis/mOD
8dIRCnPIdADvXJ1b9yhUEd5ul7mvlHSVViRRht8OU28ogureCBzajLEUC3kBp8dyNAutIZ48bOb8
T4TAP0ApXEBTk7TX8YFcUG187mPClys2T1ZyJM7IUJ8oax/d8vcLhPHMzWcixo56vzAOktM/nh5d
1TE7qASu0KJEXdRWpQ4ew5c9k7A5o+p5J0JYKhS3R1vKu+tc7lI+HhDg9/HiCqxbv4igwIVV52a4
F2Q90n250FWHEQpRbOYM3ev6PIoKWHT6kDnOqfYzsTrKyxvaK3vEC0FaLCAiTIYu599Ml/Lu3s26
nDNm2/Fvgj1FNnY4P7pozUjzMIyEcku+JwexVufOVguINggZAPt5bl9i61UVqgAmvaCLLViiWrxM
w+9mf4vlo9JuXp69R4P5EDNlbBMF6zAdWp3VKevuJxiOdkuJg4Q6tJirjDJezCeOZ6cILjSNDdPc
k3DUZTs8ErQVswJW3fS7oQki1WeDv6vF52YHy6v5DUpSxXIHnsr7tdKxX5Ldwsi7D5nZdkSPOmZN
V2r6rEy4LzdiqnzQ8QiCz/s5G5MtAH7YcI03nKlT2WKnyAMZcTB1jwVabQJ3SZRdYQjJ6s25wFyo
oBJjkga8tPnjKA/MS7ZQOhCC8wh7V/ktJPrHDmonH4nUEUY1SL5y4gHUpDzRb+Ejl/q+tP8oXHzp
aHV+c7O9eX54LZMlruw99qPUk13UhXhdxAaqVq98e+1lNEeQP5oPRLsNIbeRHQA0CyAiqZhV485m
4zUcGrpYONI1629d3qwuovG5UjK//vXkk8TgFZKcZwfR6IKSf0s/Hdx2sqmmMHMhkb5a+THw2hcx
IWHMBDry5agCCRgJnDMqvLVVyH886W4MHNyjLEO7KM5TUVaCV11ufIziACgIoNBPS5pfbPcRTJmV
8TUiSiDZ9BbPNVhqi+jOEND2vMpFrEo1fR+/DtfcJgFMy2B9zScCVA0Bir0AUPYxvPglDAyvcVHh
4KDSs9us9rxIsQ6hQFLEUltcLkQSKb67w4Q+HPjxClF2yUeZQYtfVWVwyzfcQ8UJNosZEaVZealw
pQnfCWEatoqM9ycF+T3sZj+jyLJqEDjyhNcGq4SlY0hA7qXYvPjjh/excDDFUMKUEDuX/fGLj7XN
WABysaIwqsNgNCiNTSBTieOvKlgUXQ2WnTAxkgSy727e4ZNzg6uBKSHVyxL4roLLYNdtGVcwxV13
VwTynpjsLZ4v1ru7m0yz+YxKLk+6kqj4HZeuyiunZqu1yGUMSNR9K4XqTAtb4fX7fdx9SuvTy5Ay
8nGOb5aPcE7GN8c5arfMPvdox91fw09hnkXVjRaSOYrICVKHvHfalW5ZnpDioEWKKWcZFAnj2KQc
PwdI4fWgSSraz1NHXoSgetvAiIk02f1MymycaNJW2WKchWtFmuR2hqiNivYRl4M1MtLCHONPmmGu
Qmy8UBXW/xe1rQVh36QCw8jON3O/mXy9/1vG76got14VN59pgJ84CP0kaiEbTUYNe8H4cx6YA6IL
twq8pu/3JmF86gWIu4ua+uRC/LO80TAYEPddN9iJG1XhQez0wzvNWy4jNw7EoSC1jmmNu7/I5Y66
6A+1P3jWipYqz5y71y4FPtJz2ihP4CtHH5LzPy0HocaKC8s/sZ7IptKvhVqJQljBBlsyLJhPUGR5
g8uTshXiaXyg8Et+HcfSLQ602r4R2u3xTlvVZveb2taDRKd+WOhDPH4oIEywciV+DCIWXwEo6EMJ
SgSxuSF5h/Azq0bZ37D4tpn8ZRx3DN1chWH0xDr+k0XC72QQPqVANd+XBCuWTVHo1Dfd2K52ubSN
ryAq+xsvqWzrK4ncLwRM0TIp8mNB/KU7wm7Ti6bj5Wb+5mecdZ8d2qyQKcsiheju+sEmj+Zx3j1L
egN7CeH4rSRIcVVMTRj0KX60EP+I+1WgxXmaMbIdYLHjGQR0B8c6HPUWLWeASTKcXkrj5l8VoyoA
+IbAhEPcF8QCVKho6xCrqM7OauNhj3jWX2fk5qC5Z74hgdFSlIwOPzhA+AjcrmuKmRbPiWc8whiy
Zc3HvYLGFR+eNtf9geq7w50+TWkbnSSjg8avkPiZKiB38wwq74+f5FxxZNfEoffuikQ0/xlzg28P
r7vZWaLSzo9pdAJMKSl97RX07ZN4cl0TqrM2R7cL0Z3HM5UILOopBL4rVDImaZ/AHEKL15DEVLdd
ftNMcfT37cw7TQebgkSfhF37nb5DcTD4XbFcukSRbMANUEGCtn1F5SIO9CyMMoEWQ9dJdBAnIFDq
5TIBwAYzlhsa73POigjBhkR9d3A5W7/NJNc4Kw7YJSVYvVZ/MTa9ppENeUVFEw6eIPATL1gAydqh
tZ39UkCfL8+j3yCUZzBoEDl2Bwy/mJwTv47DF45GKuM/HZk53hyLfSisUhqcBug5ttHi4VBZycyI
pjNfqgZXEA6RMprnhK+VYAVf1eek3mAfTQ8m90XkJg8X+VNIeXOsog2rNlvK8fE0dWU66PV8jCDU
h2Fy6xfRPU7Ge5IzOAiFBYqrQWpix7UtiRWdPcWxjy3XyOgKWiUw3m5sO2ZK0nYFqmJfOe2EJaZq
WIRGiNmRVsXKLYZkWMtu73/R35EEVr0R+yVUpaHtBvGOZ1i1APid2kzIGW1qsg/d08s43aMlwWpO
LqNx5EEtN6yafyjsH1fN75eEc1LID8M3y0T+IX/IARNzjl4CgVB7LbzFr4oY4FOkNc8l+5Nq06jn
r8O4Z/avXVa1BC6mdsQC7rQpjzWmNqpXju60Kbrt4I2e4ZESakMTLOdZCpBKvvDaPIk6l5lAGrVm
Ho0qhKi8R7rPUQZdm/WTkgE+2pmTSeyW7ucllkEAA1H0sESmiTAaeN/e8kzy4bjuhqjkAXs3zg1Y
m3W5eT+jGKaw0eRVsZFfTdxvwdeAYr1oLRmz0WN0Q3egNoyPQDqrVOnM8t6y+qAMvhfMmA2MbO6u
VgTlrXu8NoF1RwTF/9lY3fbf15Kp8DROovjHWyrdeWleZ00xqvc0P+ImVyVpU9MIqqu5S0SU45ku
8/QwPETPOT4cl8UZluJFdpQ+MeazyR3N/ZulH8bF1DqATJoA8ow9GrpdSN/PWgdRYR2z13rnIE4R
kIdRXYjl0iDTPtg7lo82ZBO5H2gNTkdNhrLewVdWywAwu6MxabgscmuwHcbHopL9ilQm4biQ471X
6YwhKs9/Gb4abeEzdW6rMhab/bh7mJ/bInoPKvdGmIeYuD5P2/m0B5lFN5h1OuG7Z0JIPe9P0gUs
azPo3faBS8ifchMc3S48/vCzM3Oad8uU9MUtUDQn8Ci6VsyULKpS3WopdsYZ/byPkb4U4a0/QMds
wUqp8uSioRa5pIqe2smbIO247ysnfxbxkQUb0mLy2d6Si0QpFd1G6+G3wSGK6s50uuS4QmBQDfbI
ny38L4udvaguES2T19WbTGqA6qPWcY4OvvyKwRS8FWqfSp7z5RxcxW3tuKTGU4mTf2G6rGoqD2Wc
WtrYJY5DkTQCz4dhjYPOBoV/CoagP4cz25GBkg/P0nLFCaQR6LgiQBo/c1ywY7iTStd5/5gkRBvK
lkaCytEM+JzmdVp1QL4ZBmQn8LgvcJtgU9OMQBDlpLD36kHzgShwGQI+AxLJoGTyGmdNFVYgbcW9
qYl50XkQx6vAim6K2sajAZiMwX8Ivr3KSNbEfUzmhi0xwFeJSg7p26Uo+nOf98NW8rxIUiAac4/l
SEyVNru6S/YVJ6/uadSsBoqJDQZ+6QMuRDxKDNU8RQgHYd3dLgarnGX/LDDqHpAjS4F8b6j5Zx7V
bdgi1DKgZvHbb1hH+lGcmycAV5XEFSO9Dtj5sPDhsuU2N4jlN8DRy3CjPg8xsz0TfLHs7f66rTHb
AA+yPnRFPrcojvjwzJ+IQUMqvxrJdc52zFwHH+LsXuWU7WA4HuANl+dbh0IC/h+Q670DHZiKt9LE
Q9JicsyFgnB3AOlfjvumaOHV9VLYoUtEDmmh+AjmJXNUqkxz3ZGt4eFgvMQ2UlIanTG2OXimmYnf
gGPXHkHtHb2wbTg53B67NThSnmQu/O2GmaXn6zxP4DlGdrM4Ze4MAcsT04QsbNEnWFO4UILCsd2m
MZm1OUNHtjVi14KN6IFKTjjGaKU7I5MZdWcEvwNtkzqe7ToqT7OmyiaNUU9Z9JNhhCTdGBEnzDNk
ue6r2ajTfkHkCqp9mD4dMhkypFKkyzZVIpv01+gq4huVCq6n9ScUbI29EL2SjRDRs+LZCMBNIT+E
+KwgCB0/cMauKEpw9Pv/LnrzHAJao1CDEIrVqoxTbcvzKXcjWP1ca9kzY5DiCuu6/yLzd2p7d435
TAXyu9VH8j7R8mFRSEssMCEMvUfHGNHzHTAyQq3Q5K17psMSk57oIJHBk6dJfEgNBJhPNA5FKCDE
cyy9lDUf5KfJCxmRyiyIKCcyfLPaCYFaLFAOpIAuSlveDRRl1tspqtD0Xl0/RY8IhGYQg8/VX733
RqvqWlpq4xqXUIpm8h2XcwEsU52eWKC8bJHpNUwuha433GGm09U361gu/3oAWokkC4+q5Xla2MFT
Fx5wnv/TwAUo47rnZfBcB1elqMZHWFdWnAgG2HnWBVkdumftOnNvS3wG4taQhpdzxwmicfffUhNm
d7Fh0NTl0xBA+MQYcbLNlmTC6lR4DkDkAtLc1YlBU8+uZivKgA258tJZwa/nsLuDQ+H3VBXdy/uA
LdphUIGS8BVHVERbDqieAMKLZbTooDKPSQBUfwgqO1JmY5UMOQFgKxnLm0KbS8af27rdkjHq+jSG
9Q/LbnYqlWUL312JYJW3W5wblKuGO6X9jhpiLfh1hdWfKFIAxUVgBxrxWfVy0OQSthAKuhYrm97H
XRnQrArBPgPIUxz3w425/u3FvN83wuTVahOUgGwfkz8TMgHa76TU2+fO2xq/VILD9DwIeCQQMNri
oJ7JAcIusyiTcEBygY2NUMpJEv5wBpJ1YQW6WytdrwLNFaNeWdFwL4OZwg88cWsnDazm5Dc50gwi
qB48E1LS5ldeTb3I6MtPubfR+Fb7lgEmKW3ZC3A4CpYnHLi7pofpOUrSHasTuPMZrZbZINn68P+f
fgTDAshh+03K2md2szUiFN7+ktVLa7pC9sFIqPJT7Wv17XjZDMwZh/e+zuggzTeP/RW23Nf/kNYx
cCKaZRMU3+c7h9hi6WlLh2UyjfumvrZo5d4xFp+ulGZcx8Jprws+yD61sm4NlJ7HWwM1jjaF65g8
SbL++76IFML2DudhxB/NGbEhHPivewteeTj7Aox+IlVfGKR2kH5Gf1i/ofnzdgVJPLBtlkyrfHDm
bmV2RmG3qU3HbsY5uuQ8VKnW8ZGhwBhIyqrHfkcL/M3WmnD5e6Bm2tgfBO/o8wDdzHELGtv66D4S
EzVY8H04RmWvNVyY1wazd4/GtWD9E7oq2H5/TRIlR7Z5szyZwec0Bz7lqpHaVu0zoHDzm7oB07Nk
vcrVwrUvLgW1Tp4n74hUJIogvXFLfRpoDV1hBVt53XP11XJdW4SO9kaDWpK5w3EqrMaVqtlUIraR
b6xU+mRPqz4Np+Q//Mv291nJmXBWshA2mzPeDvt37peXwYXyAtFO/ARijJoe68U1IoDqr+WSMxKf
OJnYbWUo9uUKQYRRVfbSGKpX9Met4+wKkAyNs+45zgFp7MF1zhLViHdTksf59AZKRfs6RQQ3qMaZ
0ZZYIKmbHedE7fbDYE1QjyyFl7yuuKiuGJVzlDTgsTU7R5Qf4SokaSUCKpJmb9F7qCaEbQHJGDV9
QTR9+y2x7N/HDq4TMtOvDIB0ijyhQHFOwt1DGVJKBXIGrHUOwMsuA0ktsj0bsEBo6/2DexUFCOGh
nOLG0eMItJ4aYB/s5EH/Rd4bwLXHxNfKGxHMWQ8eZ5SvQA9vwdex2iW2ZAgKpogdu8Zhg5G0ZvO1
AbYs9XDYJxAnfTvq89m1qCxihWgrUXU8D3t6LnukztcqB10TnreVYrdpvMZ/eLTyBtw5GJ+hNd9u
QxoMZuo5W7b361IoMZ/9eLy/tYZj2AdNlFV8devRJSHADwU6Ebc5VUq1Wj7EI2Kmg5ax9FC4Q2fH
oVYUsXzxdU/RP8i8S0NDfIs6QjgfNI3uG4nl9fBgaO+6y9GM8KuJYHip6XfkpbwnBz/nTTh/knBM
YvXlC6sUxnfxYDrtFVZD4qltJk1fN8ZmMd8FGOTB/t4BKHooH52bPgUayb7DG1De3cytWPHef5fa
ZN1NC5JajndaCKOcyIRU7Avr654TlCDrtqNMeHgZCEahevqwNuG6srtN27G7kdgMWjzi+iI+YT/n
oNcCkbdoivQpPBcLPdSYjCedO4JKfK7jSRL/4pftt4XtYH/3XUXuFLdQfcsm28IXd3quAUvjsiFN
1kCOPxmP4vg9OKMxoSE624yss7yLF4c8zzTIEhSh2+zP+iw5vlyz8P8NsgtJxOEoHRJk0WQR85+D
f2kuRk2m4JkkTuRQVNhQZDRh2GlnuU0+hiLyRVrL3MPM2WF6Jit0foWvFLwQZXed0v0b0dDIv2sS
D1GsDI3vYeFCGqF5b27ntX6WlLli+E+tpOmeAjjDQGMDwyjgvAUA0sP039rerkOLl4KImrWaGT+2
oCmRckmAqJa2EQGHtG42CBaA4fSkEobmTabZmRORlt22rDVQBzZN5Mx1gjTpeAY/IpyG811Ve3AP
w5dpQxOAf2O39SZxodgtoI+J7H1tOEeLPXT9xNIUTjJ67SwRlzfStcnzIhZs9hMRk77apRoRsBX6
9h+RxdV+Xag+HTYXWneUY5B4NIq9apD6/vUpgQMSYFdKGWNQRsKFeCDJnAxseNW1692uDGsYdRPs
5ZY+241DOWoY9wHnS6WNETRnQvh5z4BpTU+fXm1oREcIt6joKNnAoPO9exB/AOaEWV83p2548zQV
gNpc4Fxdj+q0fsGOmJW18X6rWGuiTAvDPITmzpx48ej0gAQjbRS9e9AmLHCSwIe9BQoDBy6/eLw9
jBy+4B1ipu2ESgk4c5HyaeWOBd8lWGh6saLsMRZ6FQeLPYMlahePGGUNSdsRPo7XSVbEISx6olVK
nQSP0/Rg9nduViVUbmW8lL2yaSkOLMEdVI6VqugZXsGUlN4DPfm7Wj+QqRmk7W5Z3GIfuvMgK76n
nxT/gxUbS0allPlpgBeU6rqhEAzgbqDBpB2nga05sWrTvCYrWJDLZsuvaiUTGyyH/bf6o4+Nw2F4
xqqEjXtrm9hT5AbS9L+jrFAtoZXLmt/+5esQ5FBLVhgejvAMMn6x/Rorb2/EdafGEo+/qn6SzTbP
Gy2kZIPuFfQ7cYLzG5w7CLEu9gJRRr5v1yyYyMGKlf7iCCmTulhsVYq4QpIsfQ2nTnkBbS3EY+Bo
4JAzMRRj217syVFa3ytVOXFd69zZud2n1vjuVYJhTyDXjflRENRkbyF6QeE7tCcGKcUJG35vpQCN
PBcchuKxXZ0cV4Tbh2+NW9pknqhVgabMgxP/gS1a+SiZCbXleYS2WvAx5F22BrOv5oN8e6uHxKbp
zC0n7bfxfq5qmaw0RGNES8Q2AkSLgJ9pBVQWEiLXoY20Vww3kUCOBZgZugijAYVHbCmTsTjAN4kA
sYXacnKGXHXNDXhybfUdxhvMpwAH6nD1aIweQqgCRy0WaT7RJVQVbwGjtsorGQU/Yf54ew5XHAs4
ZiYCkHwEDzKAm4CxvE+DzsNg2c3UYbPGZb2LUEaccH4qdlREJjilR3p5z/7dQ5qriPj6dZ61LC7Y
DSt5uujVJjR2HlTj2cdqOrSPmu/gfHIyzgM/b2j5+74UNh0vtAZQm2KYwG+0tlp7/LZ38hiV+aBH
9djlV+whCnC8Yu7JTRIHqx0EnWoyDlJAQmXLw0xNxJEHJHZU7QIWIeprX5TKS8yWrHvklbMJyxUQ
HcnMnu0H1LYP6AVOmogLa+sMFwQIeAVDP5dhMf0AkWsHSSrTdhNUa2Dzz5dvnpypluI9viugZ21V
KoIT0Obwe7i0EuVOINkFQpb5tCVYentZaTEENa2eD3QxCWZKPGIrbadD1unG479fTZ2LjBxoa+G0
A3F+iyvYCLizIh0mBCzx+1IEH9vUisX7Rp8u+p8a8LXIC73YkLlWNF6/lk9pdXbkHqemwybSfNXP
QkO1rZYLeZW7rzDssUP6d43bfdFOag6xq0toAxaog5RJHnUm6F+fKzlLGT2k7mGbhZo6HyUD3GHs
Tx7chpqGkSpTOmR/syb+6taVAlRMxztApDzoEB+X6mQjuM+wp3NgxRxN9l0KRzJa5UwRne82djiR
gCUgbaCSF6FiMMZONK0SdN2zQsuQe8F8OOo5EgGFVkHtKRv8bvg/+VfrTmB55K32eeMTyZ8F9/yC
iOkIPq0mmJXh30DCLfpwzeomB8NJwK2xLSSI/Wx2HALDpJ2XZI/h04QeHl7KUIL20BIgu/gcr1qq
2JwT57k4kpD5PS8rV1MtFPTRn8yqkYEp5zP6kXzf/BuHhsXFRqPwRg5JR5oSKH44ivladRmuEYtk
55/oef8qFIj0Nwaira/X6WDymrwWOzjTNXa4DlGRmuNYLrTYiGQPWt9OiE+RfO5zu4OvGet1bwWv
APUEi94Ko6L6O0dXeeVeV7/8m2EKJ8wNcUgevRbH7ZdyocKlmEqobCoRmEFtOYZU8cgFiJ2rZqOY
hsBkObUfb2qJjFxi1Dfx+mL88QS2OhtKQQZSsaoF57QN6yNYEKUrAm1wlH+45we0H/fmj3fxg94B
vrYKOgscQul47KpP4APsi2trinRZ5du/PLJrggOdsfyfz7iU+mjv+dkvCnceoRrAz9neUPexkcVM
TlfJnK7U1Q0g3FJGwZOt+19cv5U5wf5PXPUkcz3g9EyPXrSowXfAj5PMU8bQL10Gte8xDDv9ovOh
KHXngVza5qsnDJXiqsgaNzO+JtWcCIJNQ3ap7hKWIrcY/Buxp5JcSAziYAeSupG4z4WQd9qXLTBd
NLgiQDocr0L3E4xne4WqUpyOpsPwqCTZICJ/gaYROxMuRA30csZ0U5KNvcH3pf0eC+KfnQz0tc3V
e5GSBQCshv6K1EVJxwkFlDBqSt8zOpdM8CPgPWKVP7z0swBL1l8Wf9DkGVj5gm0d1z4CAEY8HFo6
pmLhopOb1kARhs4Arcc+Tz0si0P+cax9bIGB7LiemnTyORzd3CrWrkGCJg0jKCNd+CUA0E9RbZjo
mETvjTQKs7ldrjc+OpajtuOmhlf7w/5YV0tjOcp9iSOd9BnkqIlc51c+0rXXo+flvC+2vrAd77hh
26ETz1tESDN8XN7MCZEWuXSrBIYcz92I7jtLJdwrqgfqBOjclCegQNd8GKjEsrIRnoxNIGexfjT7
sBfdmMwzBIa+9IHkha6PpvO3eRFKPSmYMsloMrQFDSMYdkoaZa7RqpVRaArMrMDV9yOPCSgjwt0A
oyrbk8Q+ZO0JMqLWFFU0MmsczlVUcontwmnijieoITJJ5CIR2oBXp48ZIpp6IE0ZcbdOwhrQXKsL
R464IArokqjsxy5LYfqxnQo8mSf0BhGVKku+gBinKKM+xl8N8iXEU0svtl1UnxkO/ElISVOsSquC
klC/Wa1RlNTERoVAaMgBGE0LMpkI+QbudZMC9jCAirwJcNqdYg/Vk0wfYD0Bf1N8YuA8XLisaJar
BmI4G4vYkHv2SmdFqiqG7+dqi7wpUMJFYQ2Lc+ZBxnDncFOnq5S2sycZB3JsadUIUG3+a5IOqCDO
uu3m8vfhiCb32gpj6VCRXnBRg9s7nIqZl3gaqXTAR8fyX/9DIruryTSNqTtyCZwgAdZ33vpraAuv
k/O2ZgKswc0XcmV2mouIep7TYEvUz+E1Dvf9SpDEYTRiIjNnktpcGrkgEgiQfIDbpP7RhBaDjf+6
C564rSJJf7tF6BpFUBpxWXC0XyTljTJHMRe4xfLbgTht+yK33xadXhocGEu5mFywphkbmVnsXp5z
rCVpEO+JjoaaF/9crcKsKy8MZXhoFGj4RMq64S3YD2YZf8JxyhdPTafwMQLKTuiFzUFiHmuK4/E2
LtO43cFZMKsXhmiZL8aVdK2OXRjbGvdzXcOHrK6Pcx56MDQIQtr0AuNtjea6LhyWim0CGWxTaN8Y
hJwJiZ/uQ0jv+tpLMVg1O42z33cgPrNYD61UdGIA04LjfMQYdMIfA/HRJMNe5QbH4okSxZpjj9uF
js/ojUwtvF7VboifiOO83xU6fZ96kk7d06CQ+2o2hZb8Knts+uDVWbHtrIiR3Zab1RSZya1rZfro
AGkC/hToYZyR40A/SRvrMlDztpUqOzohyg9qBv0OPlNNTig8k7iY1gfmoyXvxg1OOU9dT9CRKAiG
w+djQxvYOguUqMvVMOdF8v5PKmSkVcomc8sGy7KuDfZ8hiSobXdQbdYdckzVJaaFsRQlIva3KX6V
+Mm4RAA8ZA3R97rTFdAuS46Ic54Z5LwQbQM9DZJWK+KfdhdDkFPwofvY5JP1fEj1VGtdLa9NrK64
hlGth4ZMDVf/4EHV9JLzgTxKkQHt6+A5m9ujDtlJkfpla0KyjllyFuhDQb8T3PSoSTHO1zT+5Msp
SM1fIJzkSVnFh2UYJ8tUE295nxRpnhd/TVXrKjhceMLK5KQUBO3v7ezr/rU96f6kMk42X52jlP6S
GatSOE75lEm7LnFsH5qgTxcgWlbTIj7kTr52Rv/wsJnvb3nPJKCbrgiqkgkBj9JPLGG6hmsW9ICO
YEYrkonBhC2V6/gW30YqJhHphJ6VPBBLdZUdBAc/AjeBRMhG8chhLhCrjNpxhCN0wwdk9Sa7TMo4
Z7x32YiwhY22sfJ6bmqZ3rrGw1TqdYfrPpyDzEZCpKaxHSNUuCgKZKGijjy2w8lR1EjPEJ5XHMcj
jXrxh2dOE8EROUFk9Kl3wdJDGGP2jfG4r29LKBxnmt/xfQwtrR4oP9ybNFuB1d9IQlrubcBaW52m
QmUnuxdJAB1zWEmGav9lbwW3E9E2+mB+5Y/E6oo0nQVrHuJ73fXTkFF+O01dZjHDEKkHHRPGW4ge
KK8P4n8FyD5z76F3FiKXvHzOtioc/GCK/T8c0HO5CM/VoLTy29IT87MQVUg7NAyDEu1Rc/txJQUE
e2latSK5+xV9ORN6novaGo6airJOqKyEqBpEwZZnB57mAYgwZWjihGeuAkMH6QBI3y4nzTLZo7VS
eAwouKCA/GQt+FaYgWN7U9PZZddUrJze7LLRaLIdJeGBhGkVEjT5qb64smGxnsIh/NhLij1Iq2Ax
fgi15++flSn+b5UzXaer3ogdNjTou1dqrMaIPgtwqaaUEuIzU8YN+BH5m2K2qwt+WDSsvbYZ/YCH
r7GtZ5AwF32Gp0OaJq1Ox80BOBvc/ueW6EnzFiY69pSPYE8GUz0Z1RZeuQH/ecz+ggzLxFgJ5y0l
+rApVAVu6BDp3AisY4h7EEp3tWWxCb1Zxp7ZkcADxATda4GU0Z4OheYRYKq7uxFBi/FeRqsUdE6A
zElXRi4Q2rJto5kjZ2EkENC3nnW6KNtv56MEZZZqMUIpNVMNzkwvZENCbmxYfH7AHkU4/NFepJAd
0Si64u0dbwKWCpFtFyLUFfngp3e55WLSW1iD/shoLNGNOaySHYQH9IirgZoShVVl1OV8KiPMxUhK
+jf1h7EL9uw4n3vI/UPZzsGP37n0l2787pD1/z7T+3U+CaC6SOc518+dGNTleV5vtEVIDXk1V3rw
VELaehAQsTscbSs2VpZAfgx6pFO7MeJaluUKugwqSDwlFka7xmhP5AkepQxtce8JnhCMVrXpTYIQ
xt22oAXOUIhIBdt5FlyPVieUB7fScKwkD+GZvEsh0V9UUm2ogqAoF4BNv7K+udMTvDWX7aeQ+V0J
Nxyyt/WKXp6+ssUM8q88qMAgJQws3h2v0g2RanVOYjiJQqCHRsBgSS9xD0X5xYLwo2re6kMUO7HS
gS12Ii7M5Socph5fgnq3yUT0lObc33Ft4Gg1ZbXZUxWyRj+C5plZjR0wXa3HofbiYBbT4IJj92mc
+arubxHGH9JGypHfm+reg7jrWbTs88uWzYxK87IlMam0jr9PivtNrVS9D4Uj4n2oDr0XS6vwI595
xN2RKouHXkJieSz5aCjyzC7DEEBeoiR1aHyIbY6RkQuhHLAWWLIy0z3+BuWQyWlNx1K/uU82o5pL
Tin73c0QWWTCPKx9vxTqyusAphClN0QUVCcsVoFIhNiRp9oURj22vFig/9LXlPq9wsIULkFX1EKR
WqiSGNCXYqKXiSV6zHKvzwHTM3SMT8Ofg7SUSxl908EcWLBmCVxeTCrAInUOI/JcbbGHDCCv3L79
TBZvMJhSuBcZm0YXN/PACiTXn8VA5fHCu+GXTlVVhgn4m8s4369MqFt34liLRMVgZ0RlBx3S6Dua
x8hv2qXw4C2NtdV1ktU5wMDPLK42VDxXQ/RvJRP1a+dhhkSPwc3OSKaYkgbc0wScRGoWdo5DTgLJ
LlFmxuFmqq6nHSdgFug6iTSC0S2SQLCCojKV6wyPosWkRMAcOq661zXZ299kwtm2/FI0ASJ7sfEm
2hHcLd9361ox+GArru/iCPtI0CmfuKkFanLzgX0h05ZRetjRrVPCIdgCQrE4S8G+52MjIAt+n/aa
WMTaWSyUK1Dc0R/g7GW9l4Hqg99vCP3szxn0PIBi85FUeF5rsV5cN0mxh3HqczatLW/cIbiV4S37
DVOZvfmiK2j96g1EZPr/+YeoAtdyDvmMnJYWHZlx0bgJn41owWW71XBcEQN6mjU5wLDJ0fXwYNNQ
wbUOwGtT58HwaawLGghPPSdCgRteDTZZ+eK3sfeooVyZcaTSSxHMhzHa3+/SCTQh6Bfn6OnonkBV
YPUf4fjwdz2jlekZ2ON0agO9bP5XLiwBi3jViGgkSn6uNNbk+lTqxnnGBHCiqvMI1NSd9zuJ5GgB
2ZlGsMO5GW3EJIPJW+fZyqKtYhWRC0Pf8BIf6luMqE/dmKryvq+Xvd3y15UmGfYDh1lL0gnYAf33
1mfcIBezFEddl8b/B7wT6qTZYyfu5+h2i32EsBkc9ZWx9OPBfPjGiv+qslR5PbvlYaz2PX6NGeNh
03e9rXqRKUvX7m4xiu+JfOxbKujcs6d16+6AM9jfhFBDnlUHxkmNHfkwDwAtu7YMGuLV8a4joyMV
+eiHNoPqzC5WrmCmHvmtgE0e1GbF1VD3+lmo036Jw3uvze8m3LGGX6Bd+MxMlLGcqiW77WtYYDJf
HUs3XDWnjvwqjwSpI/0Jn8awzw/KwQ/qvVnpLmYD7ADUgPrOc9jiphAka8ZQYJ/QwgsxxuJLafvi
WOd27ydN7HHfQR/RYrqylJ+LbWxo85/FZX7iUPfh0FWofmTZw3aH+pIHgDAtaWsFsNnH7MZa7IqF
u7nZ83jJTFZrFcImqClGEV/+gCt7gANNQHVcvCgFn6fMF17/Jp8Xrhhphd1Szi62AJYWms2QvQgU
HKTHZVIxoToZQQrnvNNz+Eomxmlb9Xe9+MTSvZt4S2FNk5IoMSIFHvgOhhSHI1IXU0WqlOPNnQWN
f9ES8/cTTo6k+ZdJT2ugrYp9qFLYbDtzHAkkEmD6/e8lBBywZyCDtksQmlt0pfLrrsT8KEhjq5a+
moG6cl2Z5nEwXpnM422Bh4ZmT9OBXHY7AAIGjm2yWIBFc/hzN+9nnqjZfbs1gtwxj6geky4tVgLz
ne8kLquA7PHS0IE5x+PvAezayyLmg65KaAUshz6Z2aWz7Ejnn7nrOWY9sAvZMN/UE8YVB8KWql2Z
hLJpVJ3eMG9SThnQh4gYGP20/GsV+Sli9DLmh5amsGJSb+0nrdMrDwTobpVqWXVZrRnGLi4UrrDh
6avr+Ehb9n4D7Qm6npY8hIxzwYXteMzv3vMjXvaSJFeYSYHAlkMM7w8gkpF8WmLY0l0L6LAzN9v5
qxVWILre2Gvs8XblEZmKnnNZ8VEQ04647v8EjB7Gv8SR9HM8gHyzVLOGvuOqcYyaMic+JoaWzNqh
dQwngldzi220iCmlh2OFHo3mDC9zN3z4P5cJ1vNuhjxHDTBtf76YshAktzSwaulhuxoqOdT2QuUK
QlJaiKamIBak3EdSFdFZcB/43KcI0aKPxqd9FA83QSBFaBfBMRx+mOm8dkQOuKMW26FmJhSKC64o
faShYoONY58uhaGwQdFplhSAefsjIXwmv4oLrlTx2SuCuNE6Yu4wP4y9P4m9AldOQRHGrxkcRAqS
5evledNNisshOQcvsniagDgjO73UxhJuYS0ubNVa/LUKvWLTF8vfQtiDcMrMu+mIb8vY6ResNkon
Z3ksme6CdEAnJvPjQ+sVuozBJ7fOYp4jE5xret0o2H3LyBtTwkiKu9ciIZVSCF/B0gVvsgLstzDE
FcQLbbrzWCjodU4SEuAdVpm5BY0OCeAE2mzXSLlOEDbHJGsnMcEkVGETEiiMcHZvhQebLTiYQn1V
7U6LTaIxs3fdiuL4Xv519cs7llKyFHVxsFFVTqHILIsfm3t529VHKzTs2pT0N6eocDpwW9AN1wgF
8VpRvF939MY0simQJg3ocAHFLFpgtQ8mjHnez04ghh/42XdLVV4yNVlhoO5gdrKwv8vr/Mhtby1D
Da6Lo+aAMfFk739YmEGi1r5iAOdFA4e73ER0dh3hU3ameCpp8bA6TKqswlVwwDCKff+zlmKEr4q8
qshvWwOl7AsxsG26ZXIGZOq61+HNMV09c9icScRDnftOIM8P7jmKmKaRz1qm/lquIhXnQo2tJfCC
o1Ae0g03n39H3NpCqFh2WMUGpKpUfpoQHsLHhiz44z5sRDoueD/wNwqC/Cvyo5AAxlbfyLD2QFtr
isQHQMzb/+giWIg9C8g3mmlm5xipf+mKGugcXk6JeP3dL7OQCNWxCxzyssFQFki6UcQqoWzboecO
HMoTJpEdi8pXu42awqDZ1jnBKvruIimchV+3pZVU88EWvGPZ9ZdyuCmhHm15H5AKxjCT2tFvR786
7/baU5CelDjxJ/wx4z176bRc0FgyQc3a5himEYSy0DCElpLpHDsE/q0+LyTgH3pyvQmDi2ngxKyB
mfybqziZ2J7QzFM507pgXHrr9B5rAqbiMY78RdzUGjPm73qr3b9SHka99mx11cIyqwpN6hDr8mEX
gjLkHfKvYt6Cv+eYpdgwuW7XXI4z01zgWIMlagr44O/0z6bpcZvKcdb6P5Kk+hJfeov+Ld+7NH3H
rvYds8m5/OUfwBBOOdQ6SigVt81WlfMmGKGh0DsReRKtKYaHnF1p4Q5HJdeMh3yllvFL5WkxH+QW
CslCUbei7xg1sCbXrwKFVREO1PHgExHpDFekIAqvZNtppjcDSA79Z/Imw1ECTw59I8XWyiMAUIIu
wr4zhNz1JciAPLPVWQe5f3fxpTe0OD4EEWxehmvZ99Ocs0Krt/m/+b6+gWRl1Xtc4vLJNZz4BET+
4FJ25NrXLbbCrZrR9FacGt6t44FmC3yBfeVT2FjKdCCcJ/NOAnftsqYo6HWLefq1vMGwCAMHKEI2
5T0BgCLZAhNpOaY0vb8Y1YQTNF20gbTbnuZP7duPebWoOinx+clJzifkv6dZ4gsewh8Az11/xamy
s7xjovrNoYhO+4hNXQhJpHCkf474tM5Bb1481EI/QakA3s+6KFYiRlvuLOQ52NDIhE9s+jF02y5R
TEs8/UjQRMGvXwPCybFP8e1g/B+Ad2SyqJcdRH0wZiZKO6XfTyUHcYerlqF6GYWDG1jSdIGwZElY
XKFyR+HEK6qupfR8Zmf32M7y6B8O6nkh4jIzMyAq2KbM7bqsOBlveSb3aOmESS56xrkH9havUngq
9h0JOem7VzpLnPEkwAlis8H7nhXNfQIQbNNGPqSW+4hA5r4ZS1+xx2t7Z9j9z4VSMdUEa2q6mcc/
0odWmFYbPxpnpOIq7ldKp7ItqpjxTtqW3fPYd9XHXXDpasRagopcQUTEoisucskInH5zf1M7GrQP
3Vnsd+sF1kBnn1aymGDKSvySzaV1LOPRmM1H41LzwSpmKHV4DKAFe1yeEo6I2ABMqjcGef2JB4z9
T0qYidqYsbZzAEeoALxFnlzTepFeCeFB8h1N+7pgVVqMsGempJDA6ifcIF8QKRDUgkaKtEKvV8ri
U5mA0H2jOvDpUcibQjgX5rCo61KlCXVp+CUdR+qlF/1hUjN9BKzX2yQs40Qvxz0ExiMV9RTUiOM0
Xu687c+a0p4aWYP72ZX5IRq9kJxpPBIMkbRRDfcWjQ7Neg1Grd9bwHpdwfj7KTZzstK4FJSI3OuH
jr1wXUvA0zU8LMUyKmwUOACNygmtMzWIYgDzGSCqDk39y2vBRUADNChrBIG1YUyP5mL1Q1FVjqcI
YIo2dPoIMOA6WBSz2e6cNjjkljqGYPmu6+pc80jCniJU4sj7Sz2xBPDEwxSV9VucTtYxWPnfYRlv
5iBn80/8cJQd6qQqg/9uhQl1EnvddwJRppg5Rl71kedK7PlcU2vlUl0EUS1QBhywbUXe0U9mR9t/
8XVN0Qq8ka+0E1cj3Uer9BWSJO4PGl2dK1OXndlmSEBazvdCiIx9HYuFFXxe5pfjoNdH/4T3TsY+
+QxurNGlKFocEKWDspfu+gb/U81BqtwmU0A6ypU1MdG6/LHanurIKl6K9qtYFBVarFe6zxlRM2ta
7L+IM6TVaHzBXaATgFJS367JGTUd7WW8N7q0JvMtsvPlZlJTqGPDuMo5sQyhsu71tr6cXWtaxKmf
oWwSUTOzVlb9zZY6mXLMuXINgdQ78Ogw5F4jOUDEeDVZqKIr0AOgAloJR4aWh4jqGU9TvX8ShWQt
EsnoklFWAcMDbL2KjD/qihZlfIhdYddVoYG6grCAmTk21uy2MYjDdestElG4n0xl2f55OD3gqUSG
Gb7qIF65I3bXD5zH+MP5jgvoVxxvXQzXWE0QlQJkK1h09wQx38CXO3MaD30Nsc18zBjWfS2KyJ7q
PecvGzZpU9hFthqxip8wo8sez/LqdapAK7DcWsV1I03jlDhRqsO1IcFEogbKQZGn/xOb1rYrjmac
UJoBWejNYGJqcLPL6fbr+cY2zIUbuOHnlspJAMarl0MHS1frON4XsQJENvxqBrJ735onUTjjt9b2
ZGVgzfnLRKUnvCQpMGxeETPFlw+Z9gFiK1X6dd/LgPUdzPfSzWfcG9/tuk7nh6cpuIowk9zggM/H
DCYzH8X+EA1j0S+xAtMIEG37oCxN1ZtnoF5JhxbIbBjT/G2IVru1iOq9zP6Ii3Lo8zBxxsLsDkcM
7ZG0pktktSbm/8Jk+zDx4ZwDcbYB0w6cDSXXxLmN4wgZIwr1iDTnXX/zcjj6Qqsr0ARDo/2fputD
FeVKO+YIYqG9sgCcLzG6hrGQGERwcITLBWJR+BhBjcWERlH6dlbux+tYKaiBzHXJXKwevPGhdG2P
JwjN1HFzNWCEp3G22/kMdTGSay4hgDSMt6osYUwOF/ztIfmGkXiaTpphXQCT1jh0SzxWiXiseVyO
Qhx1/XGBKdYvQieIehAPP7LOWoKRT+2Rg01Q8fzzuVrZF+91/5xFR6G8Kw2Z+ks7pURgF5V4Nnza
9PDutKbyGOHHXMUu3F+PPx53x4lYXcvxO0PdT2sDpmfwe7ejAF2Rxs5kSQhnjSNoKPOC+XZAZ0Zx
87fpSlcJqOHPcf7NoqBeT9wXBM0pLgSL8El4UL8LQHJHvtlal91iHlbvFgpjIE7Q+tcREz/UZICC
MEBb2yjHbw6A1qdP4ftOhjJcdVHChq8J3pNZVvtPu3oBzCMurDb0W1pJH1t1vyBctMP2wUD2+Y4X
mt7e15b9DHOOwgF64N7KGIRebFubEIJwAEDjHR10bv4Ni9dUAf7HRsy6LDSmpuTaVLoP/IIy23Ec
Qxbo+gjjXCYOA5PgAa0M6Mm9M2xPZgGUxEN5mt5XJ/NNgPiPs7fEQ0sa1lXn5l4bm6Qm6BqjB6y7
ZUczzBVBQyBDhfbWWQdg7nzSN1OjA6EyV6Fe7hPy4kk6wnUGSL3iJPeRpx+D4krwJBCm3SSM5YoW
jQ+IrHXN55SpLEr6op91I+TiCKHIM2JCecRpzh8czYCTS+E12VTVCyhtBMHgv2aR2Iw0AfSdl8yZ
kq8/ekJwkhcuC9DWEYCAAWyk37w+b32qYd7ps5B8b1pa2TFyH7u6fy56mUN4i5cYfy4el5+Mk3le
OyADzB2VHeKPLh4SbniiHq8ZcAjO+fT8grsG4lYWXhVH6ju0OVCWiDi8jHaDmn6zLJtxzLR5uZfb
E2aIQOyEJPy1NNT2f+TZ4x2KfiqubMtqSKXvdhGnyVgrf+E5JOTkehw0X32RBJmE6jdyEaiXFkhr
3+YclhzUMFAeIws5KGVLJrs56+OyHql84pWOKhtyH6gTRTWTsVs3VZVveR/drj6Q9ppsPD6pSFSs
ifjB77usBFFsJJ4y4pRhz7Nn4nVpW/En+jLRph0NQ8jbkHGhPXMtjwUQKB+jILDnhIU7p21Jsp4y
Y6dFBsH4FQ9mZwuh8exVyxjTi/G+pIItLUrMBNfSUL+w1H6y+7c4LN1Iupm6H0uourNonKq0Qcu1
l3RDnyFafRow5j9yfiQMeZXeux3QPZ/7xepZmbD866TViMEES+VFoRVnqnipEi3DyKN6r+Cov8ud
CkVoL3G12D2ZW7Bh5tX9e1lFDGeynpLuCINltqjDXmmGRd6bxkI5Klg9cpN/deS+casfdnN0jO2w
F2MxXqD+NvNwytof/CJGbPRcyFyuG495qPZ3jcZrjIrgrIVNo+eDJ6oEBtOV7/5ymHGBbpBlSgvY
P4kYoa3kJ973AQ6lgFRQisn0aVYwMnX1ycLgHL2nKWdWksRzbrCRlhSh3DsyImP+WumRR8VsOtna
ysHDyn6Fo3NCv54m4U41QeL4LiUrT8n8FvoerbgdXWno9O4udfDT5zuxtS+jiyBxQYROetUwcAWU
aNa1lD7qB4MclWJNhOFdPgfB4a7FO3kp7wxnyQIrar3rTy9oRgY4R5pCgrCvkA6Qn/FHyn9zKWJq
dYXHzuaFZxIaZoPV9DK+159tK/pHfYYpsDVIxlPSFXClPVZcddALNOa8UHf2+9rWlUsMc0Lv6/ob
3gmgw9LoLFLjGk3qkrtRt4FrtUW1MlvblNYqGBzQQ9TxR5tVJfoFEzEHNko10z3xZmuAjQdyJ+J7
HCda+sxpbezZntcRtb0pcq+Qe0dmpdg+xXeSP4wLsKQ9BPwOkAj4MXUYw+g2Z7Vjx5FEawsZNZ21
Vh43qMMTfztVkLc4tTKsQk5Y54yjoVEmfkGAzj7U4L4vRJDU/+9C2/NPTQAZ+JD9sguQvpopLcDV
TprtDl4KpyuZQfSK4HOc8dCkr/tVypSnq8KPXpulYt6Hvox+2unT2PWFaA8dz2/tpwQNTLndWgd7
1KtWYO9eE6Rpzr2kMd9iYWlokdGB3IO8JfIcjjEBntUSOO7/b2MgO2S0ld4QloHvazfaqTpjY2Ag
bKn71EYLEz9mRyxHK1OzstwkfIlcV44T5c9IiEmgefxH968ZBOvmOcpooWE+7UcctysfNzpBd+Nz
4leWqOnFhcpJMjFYJUA70fLqsW02cwn1m66CPXX7SIMnDaa8Zc9PiSZghmY7QO2fGvkwM2B2IDZr
miHV16J+BM1hR3+R6w2urxbqjzHhn02D8HYDNYTtHa/6mLB/EyihsfKHwvI17Yz40BjV59nhVnIF
XW7lfj689nubZEnvg9KRFFTBxXioHp6va0zOCTMzeHzmz88PoTUCbMWCQFKUivtzg8jWSh1Ep0nM
4Og6ofPuMFYMjXhFQCTS8jfNSLVdFvN9uJg4hgULnfwkq1bVlM/mmYxH+fRuZhaxbjSvocIPTg69
FpKUT9gv5vOo0CnUnMk9deQ+s+FivdolX8IhyjV90DvJHiBfuefM0auDtlRJZb3ADamjlF35sk6k
AgPgmYoI5kEbtC/wXi+tkHYEivRvW7LSpZtWA6A35a/jxmZv5kkZQ9b9PKYKuIW/YrNXBjPhzSc+
o3Pwh33jcFojdHgjOMKeM80Yo/baGnZj7SkNd2h/BBotzk9iD/99NgvKc+9o2Rtzk3tJHJiIbCKq
ArQmjsAcH/a11ZucKbIMMC3El/3UTyIUmzhisO0MJTol+DK2RJ4oaDkmBt4JK8iQku+2FVqsWMdP
zg7LaTSTpu7cPioEgy1Xt3LgFjUrqG4OTmYDYF0IewYDix6wxMbIVu4xjojrHMAvcyQu9SkFR9xJ
v/jDXqhkZa68uv9eKAFduLSWkXl7REcXxrq0MzjFXYz9URRF/X2KaAo2Gme78ny+lhtTjUH7GN6U
8oO/Sexg/LhIWsuSqvBBT985R3whDC1aumdfjGronZpJ2pV2FENoAJgqMoYrshIUVLZWksQPEgod
+hqR22NwC3MTuW6ZzLghHhxYiGViIe0Jo5blTh5fGs6GyHxkxbJ1nWOewa3Z1o8ORwLOzyWtyB3J
V9YoOuwsaMlL9HNuK+4W8MIkfWAN5rFJaS7zJkpwsKYpCmfnRJBJtDReZRioytXk2fcdLmYKA58M
ZWM0z8jOJlKM8H/D7tHpRLGJ6reF4nd8dJkExxD8EJjz2FNhG9D3p+HCvLiyhHHW+sEvNOJP82+N
NRilaSTA6hqRuq0ld4LzyK/8V7onu5RVQvAbwUBMl1recf6fv6n3ZCeMrcRFUx2TH/6k3/DpT+zf
CxOr/fMAWr1iKYJthgjBnGwUs4NzHo2LasA45HzUbKTI7oOhzeJqNunWZvwgEFFTIep08Z9HOsPi
1RKnMexkxqmpot2zxq14nNv1j5wxTzMqeLKt6HTGjzBhmrDLEduUDknwWp0CeSgAIB75gJRsOwLw
9kUXReKZvtzCCkSXNkDueUBoqbe5FfE5xzIu4lF2+okeyh+rlxiK6apfE5i68uzCkRIvrwVuk24i
2aT7XgvLycz/Lnyh7qK55LlZZgaBTV8X8sk4/iht1QcpmmOeF7HoSPkt7ftemMwpXg4COFKdvdK9
E5rdE3vfQhv/Qm8MMmTVxNZhNuy8iBgFiawbuxJpIKpZ8BYi9Kp5ut1+jQUFXBzhvOwkpF22ZT9Y
XtrAu/GWicRPYUbTS3F/Ef6OH5qpiWVdBmPReLBs4Jx6C8N2b1Iz0goTwZClhIgGr0i1JLWBdKj9
YOfsFpQAvt1Zcaltzy41djwcQbzntUaSb2NK3fTNENw8dZ1QuuzjZh1iqGgNaQH48Z+nKlQLLexM
zHIq1iYK7yillgdRArtLmL7shFl6md4rFmkchlgthnH2BTUfppuiVq+cPRsvsR5qpgzo0JjPGImH
rDirG5YUkn6Yhj8KaQFoQAsz2tpYhKEgIdTUN+WICQHRRIzH071s6oxJd1vDcc5EDYouvFtAbCXB
6fCDuChECKIB8+o8wqHhTYcloUSLbZ4+jPushcFltdz+RgWp2gsHRYvXP8+Om6geR4dfRAA04E8g
Ya7obPkV97jqnKph45E4LpUNGt3iDcez+JFBegBTkwtTkcVna8MgBzXMxZ/ZDVBirUECVR4lK0v1
CtCAjmgqt0xZh1Np7hK+h9JkcgVNET1dQMHN6+LBvdkp1LdNx0Hia6EILp61MaF2oSuAwCG4UXJn
vDZnAU08AB7c528nKX1Etu9Wh0f6HL5W9i0zZPgnPMtJ2ICLKs5xfoPowaWwe+6dooBAI9XxRLts
ZoIwg7O03tuKzPmTlmo72ikEeqxtKPdGncqjz1yNhqwLrQ+8kh9EW0i4p7QHY2vWfciaFiaVCvMh
kdOqOOVwZRv6E6/dMIp7fJI7pCXtOCpaELcMn+hPvGzJ70A7jDXhPhOszYuKjtsPt5vTuxwrIgqB
ZuPzSEqjf+wQnGwLG/I8Hzcn8FQtj74OKJMwgfs2fD0gI1Gyp24SsutN3j/aa6sFNuBtMerRogfC
6rOND2YjlBK6aTimSgUXRwX0WQn8jqG3BEL9RH3s5hLSlgve9KLBMDj6YFG9cDMQAo9TDWBkQi9R
Ff0sJ5YELwM5V7/WxtYc/d+SuOb2w4Z6rSRFbcaNaHaUMvGApLT01eBmU18ZlSyAMpWg3gHuNbY5
tCE1TMu6YQvCYE7vN0WCUURzg3Cbu43OXAPMGNn7uO2N7vmqtAi9/V8DToMbywM2BIjNzpMjF0Ku
MLHAlvJjfxWvTnSTfVpRubJjZD1/bgx2xZ+dpQoORwcj+TGEyD49kMpObVh9ZmXSsbrg94NTKA5o
+QOo4NJ5OU6r0hwe2pFbs/JQG+L6tAT+4ptTkQ7oClTJvDnvPrTEqXEuYL24zvpmpoUJTxhfn5Yb
XPIBuIt4VUGmS73USL8g67w2u1K1Sas06Av2IIm6M0GuAl8Iy0pEW4o/qFu2fP6oZLQ/6EtCCBaO
Msw6yiMgxT2An8d8C6x5Wn1TeKNVvbWHNF5yDb502VXomCkLltzRQfVEo82aLR8hrZ1Y8wPUojSB
QP7Ar7cM/lfzJPpOo/BgKTMJVls92MMix2Fo8QOcQo2KmSkC30GME0aLH9HgV+6Y/UofNE0T9MY0
K6CCAsru+GcePofXD5V5/wgD7OhAsFz31s/iUIi19+TiWAw5i4RyUgUnS/ApDzhLyNjgeSAhbr7i
q9ZqQLNvTNJpEMt8tW89utLkTxtEg26jdmzCepv3iCdLHLeidw+Dk365Atur+WvSREiaDjvh5MOk
1ScpG/qLgWwSAe21wkO2bfIzDk1CnnaAxFJ7vDErPRbwqCvvUGjGP41QrbF8mWDYELZ00cjQiPUz
o88Ha4Fw/xbgSVBaPZOdgbNTRgrocqT8tkrDo+3dIL/k73VA7WenbsqXzll226k8qnKL2W+Gsr9e
PCmZ9frEKSvCsvjQOatonbZ9fyyUY7NQXRl3o0rg3h/ltgua8xWxacB0eCHh4xexJl7P4ey26byg
+S0mWY01krtjC3Ikdm5JeRT+O4DkZCEnQosi7n7MnlDeezuFUqWrhntFfKKwnfQL7tY8btSWS7Tu
ott415hRroFq2aoJPhF63b15k8GMFlLlBJNyEDnSeXJ69qozuNc6h3v5oJxqmZ/h2z6egNXXuJFq
cSP5WHyy8go8e7VFVjnzDS6SfJbTSieikWy3kvFQVBy+UCaUvZVUXwnGciy7ZiakayNFCpFHRPK6
TeHwCgYhFlCoAgVdklalFM+r6DZ2pLqNOIjObAy6RqQ5NrxjOzKXLawiKmNdx1ot0f+3QOlJ/96I
KxHnMPkmie4F6mTpnZDj/ut8UfkjwikiG5QeRs2undFR9KbdN12A383uN86G3P/Zx2TUjai5qFUQ
q63FwEJF3hY2HSamHEzRl3wQpIWVV39eTE+jDh4n26n8cE12ZZXSraCdB6B+dBR8K96dDUzAt17Y
JoL/89IlDT+uEQbrukzAVBJGxWdfynAye6SSaElsQA7oP3PSQowOgTASIcWpzSfRfuDW/6rXpbGI
nbE2Df2zPW5FIVlPFtDNQPpenDzIUn2pdJLCS5Ipi1OdIgJsx9oP8ESsK3A/Hz36lftF71taVTDk
lKx4lnirHLrEM/Ea+KUXQXfjIkqVSGdTS5ZS6PtfmeIZxgFGKjHOTh2hWo8R6clnfcYv8jotaBBY
l/oUElTByOb6a9qe1q+L/ekFlFGzb2AKXAZPxmQWfD0lXACYK24lGR9UvtGnviBiXZMfQqlIiv1F
KvH3OoGb7nhXd1cYFllb4FS/jfWGgpCFq+8CC8FRlSv1RxZvE0I+BVSFyUEP8Lphlo21TUloi4o3
a4zsFRkY+INL7hktq9dbVsYCXXCKXi5R2nlY1r3sLQAxs76K25yHwDk2XeNLxX9tl7W05t2evaUC
Ai0yJ0tSd4Sf01YsmY8K2clKsUM2dpVv4tE8EWTmeJjxohj6H9SYRzmtsC4c2/B7tkqGHNz64hHd
YqzBwxtda/LQ6flvp5Vz3L54Lz/7fNUUyYb0PJsMI+XsSIBPNJ6IKx6EvAKdGZDSGlA+obxpj5SY
62MJCN0Y7kYun1RKiWOHLsvB9wpmvtrqkxyUsk/Ld/U5KXSEA0I0eekBtXXANM28aQeIxE5g8RFs
84OyXgdcpwek96FDYKLoQeIUiD2BU4uI+3LQduXE0qmDwHB7HbavFTecHb8/wKOuMUXbD6ayEVkV
5CO5BJrcz2rxlwqVJsxLzZKZuwBGXkXQ05UAHZWEHmP0ir4csUSyKIPfptesCSw0QnWSRy8KMDW/
gFC6HrxdZCUtGyg4HNH6Gh9/q1xps0RkB1MtE38QA4VbiwU9Rq7utB/+R+V5ErqhevAGEY2xPpv3
06nDJ0qDYzXzkMU9TDmCvabAbkRjnHLICUc8rt8eTF7FAFNSMDwnHwoN+2W1FG9TWZAKhtiHL1i6
EM+KM59/mMvqhUJqEUQDRIk3XFkyXuzbJBAhh2ymgNDh46rghxByRkX94TG8SFlkDAZYeWMBx9WK
mL9VCqHlVXgVxu2YGDP1m/1dTtXXalDuWh2Kw46DD2cw2qbk2TowXhw+RqzO64zWowq/7uCITIpU
7LKCxazlGz3ek/KgfZTiBgF8Zt3/ZRlDswHjqF8QOnaBlBx1oYsQcEvHlLVJ9L2ont11+vKGsNeT
JQWrCEX+RFqB4TG74SSvj89LVVUnpOIcRM425UySBjL7tcuMyXa75pcxFwLEaps6YXpmKuCoZ7+p
LcdeBitzuKURA+A2GLmT3LEMPzhCdheXXnaOR5gYITBHeivdQp5CiblQ64G8ZEgd3XQAVV6b4lTU
t+lrUwXVwhg0a5D/RnGme8dK8jJ3OJrjRC3ljYznc40inGiKBWFIGprngfPlB7PMEpF6sg8ZTGLt
3wFuhnXTEcOxBamjvYI/1ODKQbFK0HWYnfr2c5Ofl3rJNhnFK9tsgRytd0GWuAZhOEfL66oR/eMz
m4nyFhFy1HiyWpWlvmdQ9IP7hA1lBLpsPfGVxPbQIXizyKCfKZTxddqt6G8thQCZlEC4Wq62KC5W
iSID4XQ+kjrrWXNek6hu1GSZSF9tbrZnyhXyhlPUzV3Qibf91DztlsdHoxyiPD8gFE+XaE5XD8YB
EaYHOUkfp8SbHQ/34ph4jgbyGZ/1LZK03GgGxF6ioLAlcT+bVX8ENK1A82PZPnVOS2qOXDGySx2O
XtUfEWyxLBkZUxtVsmJtWHtKnQ2dp5tbklDj2fn0Ue0/HzJIIdLaWTT2vBMeDiQvKu3brLFvQ5BL
DXorOlyfimnKwoc8XAvW58InDhq46s8vgJiwyQT4HLJNG6jyCcKuPUQI/wdYlFQkqlwBvpS5ehFs
MBnt9OxhQBpdEh8T8X4GRC9OAjzUUQ/4Tef/uBAUZpmGIazhLqWtQR36WBTRwOmq2I5N/TGdNjB0
yMiazzy9de+l47+lB5UwyyPYx3HbHrG6n/r4zAJGJA7d6zchPqqR3ahDV1pRoFRY9334HJD6V2Ee
He9aZSnZX7TIITizwiSKcLe1+EdM/PUenfJ8wPr9Oe79dtE/iZG833WOeZ5HdYEUXmDm4VKo8dd6
vU9oHsrP4pqaxyMMEBLuuPWU2CJ+vgXPL7ono/6DabCRcERbvtKab+vTc23SBcNNBHmIaiySTR63
17p5+jizkSNUViB/vy9MFc0aetYrIGWFvxgW2QneG3zh+9Vd5ME6pug1rXTk3NA1gh7J86BPgXjr
92c8ttX+cmD/HkvicUld8pFhJUM8exWqN+z6DgJ2QVvQ0uScMPS7LcH7okbu7RaoANdOouNInrBm
5TfAkCjhFfZuq4nexj9NB9VL1zPqs59ANIxgQwR3qZ+iEioUQLZME7ItyAPxo1CR1VIuczC9NGRO
L28demUCFczgUfkozGapa7K9fQuiRGC5HQIn4eD/Uq+y2eDKc/qkKK5hTYQDYCEbcUXWxT1hBWKU
fYOZJVJfsjydkrkN22Fjm17mY4Hjd+KCUgXYD1ySuwadt5fpko20igm3KcUWubEfPOf5G/fcAQH6
eDt5Mg8vWc2+jacidRpKCiHehv7jq+5wlQnmMOYz8c4s/qx7ltOGA93pZChYE6i1QX0RkXGuAf/v
9OWwg6RYW7BcOYdiw/Ye9ClBAgmLYfIhKinpNTRYRut8dbfvqwAj/8OSvB6t/04u3v2wf9TyR3r0
bhOwSJxHeMTWxN5ACSwrsDFwIsQpwsvrd8wCcV0fRM+FU74jzGPFZ4zeLA0QD1qCWO4WVAlczoU8
xRyRivpcP+tHqLfyWn0Zcg7ir3eS/88MCfjhXg5wJpmUu6w/g3t4u4HE11jzkFTj/qN6Eo6+Dhae
+BuDGyhvSg8q9Ic2Y1hy2Hgrc3/9Xxeb23JnJAeM3DbbAHB4oCQAjDeaWe67GMAVnjL8i9x4ey4N
u1f5iWXdjRiUkcXkyheiwK0xANBoJH0rTtHcJnZjB0bNbT2nqLSxt/Jzl3vXWrPQnGQFWUkBD6dv
X5okonWz9C12ZJfaOCTcxkMR6Ic2SYtHijrDBwI+txfzX8lAx/ONtq0Oo/gTf3ukwdba16ZqWA3Y
AIcBhz+FsZeqXQD1RkKtv72ldpuv/tedvBw1LZm+jkOV081gAmYHb2ECWvjgnhe+mo6nNAzpS7kh
pFdetCfnNXwjj7Ow3Wo3X5kBKgpHkK8TrFNWpwy7aFOyWr5gPeKa50BkUMuie6QccFxNBybu1K3x
HTtWky6WgS4yMYlvenvaOmtuuA6JwkrlH9BUhn1gRMUWz51leReRUv46aNeUJpvfKvRznkxrk781
fETH7FaWKH8sUpuXBScqUDCiHaoCt3yUsdhmVHUuyviUB6weL29JLP4ssqUNn0cANV/SHgdp9csi
MJyHXXJbEkFNxPOiOtZTwhcflES2JW3KH6O2fFTgv4Ul6TjveN/Ow1pnjQ82OaHkXDF4avd/rBiL
T9vSAzpzv8Hfx0ccLDcC1Ayq53/SyDY+ORX2aNEQHVRDEAPJUJinXPTctcGIRtFnbSYU52jcJtUq
19ICr75Tk4APRyKElNSnPYNxfOxbQdA6PfuXnzwu8vZ03H4qtCE3/wVALg7JK1QI4s/B5M2nwXUt
YxuSLt/U6gL42K9llK3j0x90hTuvnNLjNirngQhqAyLlOcpLVosXYo5G2IBQ2FA9EFmaPEHOQ2mL
FVLuJsi3yiJr5CUi87Y+HOxdRCCESvvuvxur6YFrqN7ywf7cuQVWcbObZwZyC6aM7vobkoqhKeYI
afqMikdxSwCK4swYGXTj5fj0M2PALMPqUtsKgnXjpKKLY6+ppA8s1oLjf6QyDTY6mhwFQPT+Y58O
eebzXFnzHB3mh/UQVw0ecFt6U2T0coHe20mYeDGgtw2PDoG6KnFOmxvXTbBsq4bb/JykMhhJAOEg
SwGk1OrcAQsfgsIXNoO1ysbclzqzTr4b60qAOjtDNOLY14CBNiptntO0v1tkoUghL/imj7z12zo7
vUCIpj1BVXGqcsFvmXYzYAUVWXT2+8cUcUbraSqiB4ZWptRhexGXpZnOmKQt7nKuoNp2COSjHx8V
Oh4XCSYcUiacEXQXGNZ8yZkEbqWMl72YI/Ong0O2aZEdE7n/0wXztsWTHke9heAYRHi4TLgAwnJJ
fmPp6zhoP63yg4Hz6kjGL2tn1cWvAk5ccOBXasrOhK/sg3FdaauaQ2iyev21NYFeUs7eLccA0ovv
5yg3pzwM1BT8xaVfbalDC9m6n5sItvOBx+BSR86JrM6CO7eZ+jB5aYb+Ily8S/fxUiXCA4o5r8xL
ULWRZ/hX3P8EhG1K1c9CnA1ki3j2xtu6qet4njS443028MU1LSABV8M4/0ujHuxtT/8WPXDFYVp+
TLgwVsGR3LSFlRcA7bPcY9QDZ9xq60kAWfHHEnomLgOlt5HmHa+yFcMcBHpgum3DyBZWs/PjOw6+
t2jR8eKK2T1Mu/Z5MnT8LH/gcVtPzyllGtAtgE2TO9UDJvLT1ia0AWkHl13EPCX4o6p/N5p7sRWs
3pBBduxHN2mmfxACBhZxw7aXlXTjc88ssDG8yfMO7OM3OdGSPYNun3r8UJBpO67l1pPQxOAZv8ly
BF3t7CLOHVhd3cTIR4YZmFe8I3wjqEOWkQcKLkL46YLyfNMh+Nb04KwhVBMu0NejGq/nrRjUpS7m
IGDGX1ziinHB4VmmhHPGz1sqAPYbBYJhB1EbrFizQFamfP5ytsYVhZG6iIxguB2PjLifgsHzDsJo
EXg9fqZTq/L1Of5NP6q/CbF0nAzoFbJDDUVKyzU3DX6pcnK8Wlv4eHcKwfzarARxIJw9wLIXoJxT
oRLNdFIcrhxZd8VOG+H+4eWo0MES+ISS+gyQSX7xBFSvo1vL0zYEu4Lh9GT+uU4Gtq3dzehdFNE8
6jerMKMP29i1FfkOKVqjYYDfBmCIis3VqmIDgJjygkoT5f+zyPA1i11Ncb12RfYXKDHhnZF7rnQN
FtTyoQDgH5Qra96Wkt9Gb789I9oTWqTDc/cfXkxp2QU3u3YoPPrU4LiBgA7IwM3plGO/ajsHHEEd
zcDbmi1mvQodHp9xi/mC8A49N6Dq138/KPYqskt8urW5x9MON7OXIF1yhWQXlt5qN0FB8EAQ0tER
eQQgVsYFu4snQTCgpZHdunJdNbQ57I8VuVtlChwReF8WIExwwame4KirrP+UMZUsT4wzAq03QkqJ
smb1jEft2fKMhl25UZxjk86GJ7kxNOV47tiCNje6dFelhYzzBmsekUDMeRXpuizKF2PtBbAK9Njm
hvBRNDtJ+YOLByKSOzs1O0PuU3vEkyXxSUeOKluof1OMi0ZWrnD1pLYdWZsZ2XLdcUl8GIlFc4wd
fn6JqB5o8bJFc9WgTfqBELCUJw1O8tOO60xybSCfboUfKv5wIwy670BDLWx8Bi8YKM8tp3EuPTQi
9OEVE3yyB8R7kNZyArTtMLy1diLD4mWUJrhIs9BMAEeUhznaW8chhA7NSTDWFLXXKOLt2LZFJuWP
HmGIaga6/HtyLUovLnEaWjaEjc39G4jOEEaOEPqNiWWR17/rj1J3OG9g8Xt0+jq0iapjvoFVXAVa
G+U8Loecf9rOR6Ka7az8OI7Os9GZpq3mEOaRn4+Ng7EKoxzAyY4ZPkmbzsZ08G1RtVox6M7Ozbpr
zmoU3lf8mquNgYleW5FaVbxkCIz5JLVus1h4mk0BqcM3iqCGuTwQDRIzFhXbe6wKlIIHPQ9lqE/1
kxXwRVrLsHGHR9pLa/YY7dlVJtFbDOTeGm8GvpuTqqdrP7fP0+LIlps4mHfTKuAyIYv7BQ9J7lnP
o8e3smdZO3ZARMapG2jynnEfA2v8DqTvwLJQswk4bPRW9Z/4DQjFmocuJG1izcjnFZ1I8tBeoM7E
4AncPTq4zrWzjbENM6YF9V6F/fBcfzfMMDIK3WjmNyo0QXRr2gEL/d4emJVRpTkqywFOKHkt3kGR
yucNj+i+qQtYGqfmkfbhygI0eMwk39UeIFEtMRsDvPuMAIDRcH3feQU0xrbxOC/DL3buYvLc1JB8
iA9ISBAKaTLm0sAp2fgujIlkmo9Dxdz8j8i4eBcnnlO6hBEtlceOXco2gyX/JDYlNodbyJE+sY8d
7oP9OPk04ENNE8AdyPYmaSbJAoliQ677sA+r3t/2EYjzrRMABeItBoGi1ShbqDFuWy91tC6yJngj
T34cs4u0bcwDOvtUpdTLlud4KzbjQ8ZtJ58mYT/2mmCbSMigX6K7k3fyaKt6YHLJaO9iqjVl//S3
uc9HsVyJNK52aC0xBfhcAx4LdEhr6+8BdtS1CLVBnYI8ihYv9HeOPqsJpNwFg9fAJKyvWbO684Ra
Ly7H3uYManenlNhsnptpG5mkFhU7hqKXgLwarpea8v6YeapByY+jMn+BAcCnetAWnY1P7xEr7/mV
Pz6L4OCpmvLGcL2RkY/dIqQkIfv6gsMMrmUFFQjnuvYuFRGp8kODjFlRR40akOWrNkl/Vp8mGpn0
denrWDb+MHgpr+4gKKUxDzm+vOXhw77A4foD8Cv1u7N6RTtlYeqZtgkT3ol4DITnf0kXx3a3DnDf
o8CAI/TePXzyHmFZthxkAmY+vGTpachGDKFXy++7AicDTk7Gs58ECdL9OK81ibkS8j8nkhABQDff
Cw0yB9lOLaJvI/ju+jXcQ30W5hSBaVUiO+y2DUIfydg86zHHDPbfnDO2iQps/1V5D6d3emJ6NsxB
gefPgWE0PavZ97lkMo/Llglj3sUb0qQF4X6X9PuRmJU7kBCGoec3hHP2gmRv0Nyf2qUbOcd48glj
mKdB1uPU5X9NGGBaSsQNOpz1xlNcNq9gpDkdbaAfC/P3csHSyHSCHNYEqkDGDzDoWllFuXEEPM83
rHgzCU5QzN9QZ0pfAoQ2NFLEtZ8kT1KCyk7IfRwW/5uVNt3enVBgJkwBUr/VqA6BINYxaCGwXIgF
iG19gBXaqF4wCkOMGpcn9X/EuD3tAI0wUwalYnEZhpjX00OFH8kKIQxzG2IG+WGlEEDZALEtnA3D
j1cjQV4l46rFh50xHislNCJkm4VrBdc5Oxp675reJ3IPHuuOquxvcSJrH8oitnxFgK5uQqck7B37
x5c72vvDh9OicjTYFTbYnOeW+8BCC/pnbjXXa7vpYEYryfsAXiV+21UL8K8r05O7HdaqACcteBA7
+IwYApF1iy2eunxsHOtzo9sHU0LMIzXljXKS6/u2Z+NO0rUS8xwvKlUemstkoAIQTU5ahYyXgJyk
7EoGnhXNqccd0D37dWfUH82f6JStRI4k8RYv7VABiAA+sVejKKtmcwuFu6lWqhi2u1hwTcJNKWhv
vpsyYGxotsOD/R7lJbBrlRTq72L6CrHNEAj4srClE6xc/u0LH0txxDZu2lPRFiW49LoziVC1WU6f
GcZJqrZZfBiOVK6cuU36or9I9T+eyQGjpZixQGKmdAs7rHCfYLdmos86z34jfFSvWcBflIuwge74
W68QcBYG2IMYmG9aip27Nz27pFHnav9ozSSu/j9UVyECE9qSwaYMGEdta41Uy12AqWuElyv/SPyx
5ENV5h8PDW2QSJrlML9MaGbaHsmo+OEpZEM18+FIbMXsba90B56/Z+27sRJzrZTd718V0osa9OrF
b8L5Myo0dscZO/2SXbW1fl3oXNzsTD/uMKUTmhTiEkySlwH6f1HSlK63tV5GXQ4lJwr2AN42rOVZ
dcYqiX2LE6wohPsWTe8c+AdRIcjlGRqRHKeeatWBs4/4WClnTX3FAFfXTm29KXKgYvyv07rH0NGH
NS8U1J7jjKk7tuLo2ImKOcTjfC62AUD345noA+WRdv05FtbQ7zu+7hlfiV4GdFyrvDjPDIfl2FXu
R3mzSaWfYgxOniqgG0kRYOUJNvrmbae/iIijFwVlei/Z4erEsKJwaAjfp6fR8slZA2ZYBaigMSlj
kXNT9N/tE7VfmLzeZHWNWkvQBLsGHejF5/iVS8iWdmRuflNZlSR30xt5a+NMq66yuOzicEzS+lvf
oY80nsyUw45WIN6hWoLn17rNel052cdfavlADLmQAwKUU6fUhlZ8kpj1+OVDNTwYEvFjciiZ2wDq
H5bD1rEUqSO+vYi0QXfqa4egQmTcAIDcqdN+cbF0vxatmyDhJpE02MJ672HQooLhM/BvozmQqjke
pF5bZmSsX/Gx2fCe9KH/9nssVAs2jnrM3RacB6y3deS7edsZSghS+23FJgNVsjJac4TvbBmX9WcT
qft+4sJa8HalaqyJxs5bxqVAeK3x1M9Y0JHYza9ebc2Tfh/w3b1cIBKrVZDuLC16nG3uFm8076mq
Eg5ysEzZuvhaLbo7Ui1CpVM/H0Tuc3rrlYhZJqATmTtQNYulpE99WDZIo9/dw9RBkHfOYJ5zp0QX
TW9MeUnVdmku4sVc+v+wdsnkIr8pEkypxQT3ndLn8RjbcxJ0zecgLAUIqqDxYda0wtcfzd5IhH5W
R/W66u8q/mwxYevCkjJNNcbe+96cHYI7jBgDj3D3bQxzSDd6BXgM/rD/G3G13hcOBHP6UrwiP+Ok
VfpVpN2srPH6VCLS76FXu/hKcGJ79Hgar2mA2hg8UJxy8lPfHIdG+AdAF0BaTZcDfRev4XlX/Hdr
dYblsdFRve1AK6vLlahIdngl0sTQV7GOkrQ/OliWAfLPTaFpH8L+zkz/SwKhExxhq0ZRvtg2NERq
2Fndh6gFAnUWTISLJGt+jnKz+nmopFQXjK/RtlAql2Rpv+VAKjZNO6xnIQDTN7gp6WcqR5rMco3H
8xdRyWSJUcyc4sJikenUv2wvN4cuKY3EGX1Ojcs3vKVhOsxDCbd+lS7qvr1nfjqwSOjo6iMPJwiU
f3sAl03di+FYwB2sXa66EMc5Yfl463kCoWtsQZYw5JrwzdPtSE9lOB5iNVLUVvsHKozM/SlUeHbX
Gc3FCN6hpxwEDRVAuEbWLRqXT8vS3JAdD+aVgdrKX4Vti3Kh+gX62PIziFwZkxbKfAW3sz3Rw/n5
c+v/gBauTd2mNSoxwU4lrIy8TjMjQ/+M78vq8zqGSFZLDlMxEti00098KJmODLZz3b3S+B5c1PbP
5Ir2KSfeRiEXnX9k9yF73uO0tyKyyDl0L4zuj0E1dPkOkWAGeudWS+noF3TcYxvrYDSwuDBDNp5p
uZk9ZKk93Q8HGySU/TrYGdMHBmBQWsQwIxDqi7NdGa2RRHTdZ5MxYF1V1HDk9kFJpY57w3+vtD64
59Eycp9hSoZAUmYFLv1M5y1/UOQjR40XW0r8mKJral3CF2SZ8deGFXNfGumBkkPswZNxVel9bwpV
5KYCflFeRCLgaoa4RmHqhqvfXjriJ/0yEEUgdKNQ+K0g0PIlKLADzuz3ln//4WBkevU0B6uB6+Q4
c/xvy4vXujExU+8OD9aYRq58LKRi4DBi9sbQqev+mJ5GtCml7FsU6ZvPkfNZZM+p9NzOXe01fTc+
xeLh4/GzQKLZjclAyQNp/f3AvBgurBvISIL9EsTqsr1MvbBSGn4nHMEMIlTTcbqUavUUmbIR6KXY
h1j8/ODgTvZfrsqrWmTGUXH95UIBifV4KWIgiMqHY+wCV03CD6orGEJvlkTCTjJ1tgnj/teAkrU1
b2z/imxz6L3WJTRyqJ78QHURcEUM/sRXkEWj16FySZWv2WanrsXvl0IR7Bp5uJz2O50ZAiL3PgXg
VfXLYNmMajy0FegenTcuvOOwIEsgDWqndWP6aJxgh9SKGOrD62HC2PTfcjO8LkuLwfgqsuPYI6em
3mR5zpJ/mXNyu0iB75YAvGSPX56fPRCY/XD45o5THy/9MN7hO/qBwGz3zDyMcJIvqDoVX8nzDOFM
QZv2R/uVbfjw44wTDTlA7qDWbmGwpDiAVId/d0Mpzs9SDoIjJ5LDiDdtis6rxv+2rT3eNZb6UG0q
GGhlMHalkqdKbDFOoml92zLdI7F9z6TDrg/1SAiHTjx2buoLO5XPHvAgUgADsVRpGJIcCTeww5WU
uhpaVb1pNTDZHqaq64PVg/4J+mXGetqMqBSXBaSKePf6PeFU4P6bUfSi2AWwUmVAPTRDvww9jizH
ewZ8OR58HbI210pqbf3xfAMi2U9V+EZp/Lcuyutqx7owQi/JMMBMheW+dYP36EGCMNNc5ujKic2v
48g8yHxbikoSMndhBlGP7wK9Lto9T9zaA7CErYJPZxU3IN2ufysxD9EOZ8ox4pVmrAyBljotBHQS
LuoHk3DQ3VIVREulj3/nvejABz9wM8bwZs+WWsaRSoSuCjaiwPm9BimO+aA+uH1sal26zDgA5/AD
5o3HipGW3qbZMd7gW+JEmdsGdJzuu/BRMCsnhfldqKcVPEYt1qso8hQkLNeNB8Kg1ShAs9Nj6W9B
L0oVf0Pfqe6ny03V7m9SEQXCrBGdx/SoYAj1gqQLQoLe617DveRuEyZi1cVGL0GBd0aikhLT1AVG
wuq+IF1VJpxz/bv9p0gW2mmT5/jLriemuxbD5cPynLkmfQh9CfR3xmeKEIDsOrWP4x0AsHKHPgtW
M7yfvcfOqzpzTgse0G2PGVa/HZeza/IOLXm6ktFyAzHTlJ9wjSHMFVaTNuxQ6PczLoGml/YufnwZ
4+uEXdOXNj2dwhOZxD6wK+d8btq0U5uFvkq0vJdShWXl38q0D54f7Lt6OfqUI+Ic2gTiPZKvjDYQ
SYzhuAy6QQPkQblAfdSffVpgopQC9YXwYbogxcseBl0aETb1qr+zAnwqM9Cqfefy7F10DLRzCX7M
DdEVprNaK37Z4+Qp3fA29WNAO7ifwlPWDqOsBpoqq230N5PPY7oQgBZDrhlW5LA05CZFa0DLvyyQ
g+XsPen5P9TLlIh++bHGAm140dzp9RDZvduazeL+dsvJgQwegi6vU21eSDhrWh4eOCDxbj1J+VJ9
QYV/EfrI42ObW26Q0+j9JWWNt30VZFtsXwrtwAwyH5InGkQ5utmQnsq5ytCe465uAITmcrDf3tOV
94yltjOPNvW72YtiQHyOf6hgECWEItdewfwznqXpn0TB/I3CMmqw2MTn3Msk2t5tB0dLxIXAdNTu
YW05d2N/AFBrkyOhiTx4aru2OWJuC0ZTZoPR+5a20/h+k1TtV0xznZ2qsgq0PR7pHDsAh6w0IVSV
QlaO4Yf+/eFcJkYBsxCCp4vWCvcBo81Dw2jITBgKmg3up7z8pYw3+W2ANCecYRGfgZXOQfQfQ2x+
bdQTg78slH9L/uP/6KnKtbgcwR7sApJsnUhOwgTR4olSZYlXCeUlofnCxo9qASCRMxEZdx59a6wf
KlonDlTf7k7jD+HXTIOhmbBDbhneU7R9CnX5NX1ewZPc8qhgnuNR9grjkhNt44dPN+AOYaucZWn4
XXxdSgM71R1BAbGuNmDI5gc55RSTNjt7CkhkN4uvKz/wNJ3lxjm8CCGptku0F1dbDu771YWxQARM
5ajB4bfzZ8p5j/Mra6VywjfViMWN4LS0LQ1yby3rXep1heCZd/MCAzhxrS9WX2jLATqhByca3641
0C6epJXvDcZOfPQc2zFLDJuwRMVKBLoh8cmorIsVGowX2pveH0Ozqi1ddIsDpe548ZswKRDzHc8u
1ngovnmodC153/z+V3HIc18vxdfgC0gAxRwBrcj8xhQad7DA0FIvL8pCjEso37ybW/hYWF7sYUzu
nc5zoHhkxv61+SVIpSBD2PvfJFaD90sLrvxi5IcIW9RvvhFnQC7ZirwT2C/vxE7xYiJxsKRq6JpS
3B+zs7TgWpjQAk/GP5tAGTvnmUEJjGoWJK6H9UhVOd7NBGuGqAIO2IWqXb7i5ZtDyE900YnvUMAG
sJTxIqV+NuJ0kP1eecVOf7zCIea1lKDh1P3IE4k2yPQAfK5Y6wk+ZhStS3LqkHbNrvm4MOWUFCVg
+Z4lrAsk/WwAtfYBmUcBioBnaIU5D0Xt11oqiQXcfDDAqlMW02iHvrvHMntyPKxW2+jRHjNSVT48
Tj7x7gx0ku/irllgl/Nscb5lmOLehzO+kiXoFyrocQzUp72283jd8Kqm/Mlo2KtUVwHo2XzdMuJt
/x6KjScjGYrjwaHkUEpQYRuwrBjQsX1gz1/0J+aRjq2emDbkc6aT62UhCFyWinzkjQ/yTtJ7wAOG
TgYTi8biIjC5VTTDHbkGAak3ZL27f7FPd+50u5mkmVTeX+OQRGicBcdKb/PBjctjTQyTTT5NnW+e
ItlmOivT4dJx+br6s1AXaIBlheuDXWMKGnhWIx4vWtyaph2ThtSJpgpXdDBnkIVeojBzUbMmkiUB
k9BCnZkAVvg8mrqAbM1y/rWvhCOA5dpXXdkcinv01StgH7xda5tL9rFOnoAuk9VtG4cpl7bo0GW8
o7XuD12C2uML9CBxDxYwjlbIYQK1DU0JVzQo8yP5sLRO48fYl1rPhQRP6Ln6CGr4eR+b873cM1/c
RtpD82RdV6ApkCOZqokRxDYBHSGtAbaD8cXFCQ1X7vNTAmQ2mKvZ5ESQUXkYdzReQqK/vyAdLN05
GG+UwMwjBYYg5XQnBadiu+HsrCAd99iQTIzXOTEVfiAksAflm4hJ1Tt6+ehVYafc/U+am5E7YaX9
t5dDmVSboAsH7Ijn94vwswFtmj9U+HCSuP6ZZgzzlqqAs83JUumtNgP8w6xktCCFNg6GM48o43cg
vehZFaSYrSvQPEPsuGsTqMgLjsNRZ7K/SeE27H9gadmF7zU6/baho2kx3J7hmr4I4nyivJL1C3LT
m2GuQ8aamafWF/22140qAccAUp00WKjEno2ZZrJOi8e505AfxeQ5oQvCbE9BWr+MrYkofLEwvzwY
GRmYOJv9nglOFyvd+rIUaBsF8TJlEejNthYRDpXiKqu1lvYf4u1LIASYGwds0kO+Tg0iHyHDXb6B
PeflfzpRsHtuxiArXYtYhbQrA3JThxIC68reaEiQi+S3SgCnawiB82PYTPE0BFMa9x+B6pYm6SRX
lL8BVP9///fVAzBkcY/XnehX41dbICtGE3B+41hwjLXnJNhepZVj7ZZhwmu2OGu02Tp1740x9H97
LQk+2rw+lnweMB81gu53WIlkCI73jLDUE2DKuXO9CejksH7q8jd+tGY3i9ifSxX1f5fOUEd0K4oe
wolHppfpNwWM72OXoM78Chge8eBksj30wac6HubNmBWLjqNOOWORNQcC/8geWM7Pl6nL19+rXBBe
IbhvyhsD4cqAjQLGRa09YYTskklqsAIW3L28Hls4oS4Go2ZvtP7pUPWKTsY5/dEQNXq29FIez7S0
a00abKFgracmdCd3yOVcdG5r38Vk3HPzqyh0RWGTukw54ka6bHBC6psqAi88kPFH1K26UpNZIjHn
tC+9PhLhCVKiW9m9o3ffqw9AJyx9q2qHhlPFzuKheYQRrQoUEiCArpVXsXUWqf1cKUIQmG8DiaQ2
0uCEMPDJ7ZcvUCBfljV980yoWa1q3ipVGwBmhr2AuS4A7V9mZGIcb/onKX9Lm/bxvFpqqJuv93T6
CfKqUXiY3qc9Zw1y1OngLY4TwcSmaLHnU3zvXPIPahOWT4rBhRB/Xn70hLNBxkEEZAbx59E+IxW5
tyPT2t3dgAruSKCBaPufewK2fkLQo+OTebshY72WEWubQwQ7maAainDPy4r85SIQ2/lVp1G7Kxoa
tJrL4A3BCw5gvRViyuxURcxp3GctXT/QOCBhsUIc4ganm75mYnQfpepueh5Em8ZwbSMB/Y63jOUq
64jnW3+L6aVFlTZMcUPQo3SWeZf8aDW9VeRNihys4OlwJwjY06tzRyU1O0BwhOdkpsxQvtFzwfdm
jlw2qFzvw3+5hBQXyDVTZ4o90O5svGRemG8q70RrVGUWXphHh8o2LRmwJOuzzRznOeMtpkVWTdGp
9UnzjdB9opzevmhKEkWHlZS3upLDo1J7qb358n8xICtyK2jX0LmXCpqpwHSJwzF1jteaz5V+jaVv
uO+LWY0MTMUbc69UzNRemwoTFl3yutn5Wk0buIylGIgyn6SRJzGnLfYVpVOlHzdPc52o8YTplW5B
ywJHa5FWil2WEhQUDHB5Fh5Z5+nKq/GODXW7If6iX928VbfN8jXiZ87Enlav0P8iNnsW/OstWwoP
AZyhHZ0qocsOVzYMeirOtF686rFHu9fv0Xg9sBWHON9W/AuEIe3bdahbTyd/ONnp3S3A7tYpSb6x
tmDT3jiHLGHY0N1SXd90J2hLghM6tsdj6xxWVuphcWC7BiXQWSqE0tc9vYmaVmP+eKUcimpWqL/q
6JUsWoRoF4yFhsnd3perJ9hMt1gIaLbhj/p2k0N5bxdqpI4ghkkPfs1BoPz6NCd9qZ6ydYLa1UDD
ty1x3dWyMvK2J6GfWRyguQ1eQBB9NzbRqB+xkn8ZnjWg6mqaatJ9bNGsdm3pngiz048xCZmGCf7i
jEPV3Eu3+/gRaPnge8e4tyXMI9aH3F8DnFuLDi2LIKIGJuejaQQGpS6qMPY2NZWxQwVPFRHG2g0r
P5mUTqaXWF3acrs3JVej0re5NLRdEjCoY4zpQTZk6Y3pjrzd/SLytmR4uGioMVVEaeICpja8X09r
gLJFEh7Hnx87fMsxj2PpxumJk7zzhio1m7V8wmO8/X+roZZzRFaVzgW900WjSBIOtxoXd9x/KkeL
eR/2QquN/wzOC46dqSqxfN81gidurTQ88fgw0Nbq/nyFXLhJ84nH0E/Gvigo4HEPmD+AW1OrMZi+
ma5AlpgeWWr/FpfBlOWJuxZQrJ9igcRp42qv98Uhcow2syNzPy5P5KgW3S4eU+h3wuo0WksCrmJi
uloyk07F7BzN9xcPahCUlmrS649L2gD2WDHwNnLBXhWoxP51Hk5K6UHSe6YTCxO2UswGaF8gefiK
Wc3uDkZFLnGqpAqEFGjy7LnSrv6q7juy7QykJV/Q5m5tDDeihnWnTXTchuLOlnJjZ3taUGUI1s5C
pPruy63ken7bHbH8gwwYzs9Vh05MgfF3TOaanIJXRrUkQa1ayuIHxMQXSuFnT6Vk72yTw8p+oZMz
xpHEpYReuWMoTQU4g9ypnLiPd5R9JYueJES5W5FuGToNoE9PXP+YILR2GUccCkFDSUfH85397Gzb
k39L7Afm3ADKeXgl+xH+IcAR2Gf3+41J9xjgDhxfH/8sarJsQKplHSceDkCgJW7xo2hThbhRn5v7
NdrQ+xqr9VSqXPPfvFBqV19jhtW2sUz4yy6+Ytcg0Qldi9DVRA/4HqoNzTeFPgNvbpRD8giJaxxo
ATwVG6DNSmJz8ye7W/Pzqo6HFRSzScp2iV2N56Ecr94vEeQvU5BjvKiYyv0qq8+1edQxuNGss0Vz
OkjAZjUqJSRybG5fPe+Z9hKgO98AhvhFJ2/O1iP/4ARBfXbqdfqUcfkEZGWt58c373mZERCX8+4F
fSrCnk1HwOzdubZax7nzoKoJBtRu7TI9N3NmHloesFp6pFEap/nxkLOUbjVTlVH9xuU4do9/WSVt
P/GNHzeJ0lWCqUQwZkST/mF46jgPwzIGMk/ZoRuTxFjEXHJRhgeLBHHi0DsSE+M4XJT0GjDty88q
iWmdkc0F1oYyX7pJrefK9cNhgeWykisJgjzgx4lMXqdIzj1+JbiyLXUudwt4XtCCIbceDhsLQAks
/poo7/7AhHEtGbHak/ffSaNuRXnEtMtC7qB2Ji5Sfzpg50F9zwqwmM37bhG63uYWAro68lIjYEfs
rQYswV3mWYsqZhXhUGZfP2StQlJXMkm6POR1My0NWVA+JDsvyjtoEKj67fAIjZ11ajbHWZFRTO7s
xCztJTmZ73xmyFnMPIeCbvmjpZCrJxuEn6ZfDxLtavNs9CjVZCAIYnHml/2CrFLG0RffxlNK5L0X
Wx17XtGMR20ZlIMNBkb+bxVzDrRmyQ8peBw/CT0V/8ap2U6I+fGiXIQ18y3GlqB7+z/K36RnT3ek
OimGgE9TMuylr1bn7avKNqFTkm2onEExuImdwD/kC5HZ55SiMoHQbNhDJSdxzJm5ZBFROHmnqHID
3ltBGGAWx1cWFbw9+34/1w0GcYT+B104Ij2/8FMJRo6bkFallAWumgEjl1AywFEgCbpvATVT1R2N
tTEypd9ksqJA2nKJ595w2oxQErYbtuW67A6WTGju3YYTAcUJQMnelofOwsX8pt5L/oxCvga+fHhd
YEqC8zxJzwLYFvch3tjChIPw/mM/Mjy6cno+b1n9r9si2nF+SFm/upH2Nw4XKy5tZXHMrw0LNbxW
36nswziDdX+OR1K9zwwIPTB0Bw0hpj1RcFWDKnNpy9vtUAgtgqExcVgJ1c8LLD36f4VXBQeywz+i
p5eyOw9T596klFoPEm16XnxOq4xaZR/x537XzM+VrwsoQkiSDoRUFuuWdFuTv6b5DfCJ1qKY0qL3
WrrXJhvz4TyB8Phxe/agZpWqlxC2uvMkGidhljHhcJEkEH8CCCFqISSy6/4R7eLZCdOcVhXCVmlC
ZTg7mIQfM/KYVkr7VeepbvWJjN2ZjSFjULBQ0+AHkUieP475kBjUn28bjYnnGmfxW9D9szvjL5OH
XTx1qPHNvb8zySuliFNgUYotOdtuIU+PyyovswosuqDqKqZ1QM272ElXpiyJtafjKiOUyPuQLMkt
5LPjuglxKMSA0Dcvgl/UakIQtH13kBY42VmAGhPbKB8yT9tYv+roGJlqGZtLgftRxL3ctGHURh92
hVTwDpPNiID8LE6pTaT1dAjOfiMbBdDX8YFHqshYq5rG9z0UTp2zoljcegWXTWhpMuZ1X+yH6ASe
POKHHMsfO5vv3GwcD3dGpWfdI6G7bLvoulDyVH+dXTSFsdgzsZOzHBomk/HFoMWEG6Mkg8RFbK8z
cDkAa5wW7BxZni4UOWl8Gq7B/Z9NAWNbmpPO87uAfoZTjFXchHNe3LJdUlU2F3UBB+OU6NfeFNiG
+OrNWuo0B+gzcxQGZ5u7xpsYVRiPObHdlfLhsLXBSL6eprl8xyoCnKFrPK42yZr1/nHM39l354dX
f4l89nSUY4jC2qa1Zpsu5MOT1S1L3AJ/fEmojfm2QK1LH66o4wBjPlVSRC9WiXRMJN3JEOc4X6nL
HqB8deh/BCC3qpLp8T2yHv+iaEAD3FZI0T6uBUzc6ta+5KOMMtO8a5z8h4y1B6swmfILIWwvcL/T
mJlga/iEvuyW7giFx2IHEJU8BK65g10D+S35KieQNWnJQNxeiH8fFBfrkv/N3a1DOlfdEwPa1Jtl
HEAY0BH7xLG6J1/Be3iJ2VtE7O62sKjE16zn5/XUmyz0AAgZsXnot/5dF6l9vOA3ZQ+zR0JwiDAi
5YnWp9XnXbWzeJBSOnhAtUxZr3quXkCz4rR4jGHouKwLWViZuorXS/tgoDyUinyoBlm5MWWRv7SV
eVCHjNEZhsNNfJEHuvxtdgP1/9JplnIwsHJQTZnZ6sqhb0fvtkaHtr7JcVKVJvBUIYItd2Yc5w13
2jSdnyr8Ko9JRXZ+YghLZVO0KXroPUWwoUREF5n7ee/hkKl3v28q5DpC20MJPMi31gV3Rvt/Ours
h8gS1HMkgBUyg4Hhd9O8QrlbZCnUbAwsqd4mRn4oUqhLTdjAov1f00NnWn3U1BQUpp7kV74gG8V6
/MLI1AReZomqB/UPrbttHgtOE4DkE9lNOO1bw+2zrm/QDleuUUOQwj8lxBRTgIxfq2dh7L+7+Y89
DiNo+6WFatPMX/BLoVAuu+EqPUdSY1/5vSHtZMyKJOpLWJt/mRWJ+tntqHG4p57mQnoXiNw4oU6r
dhsPZaVSGU+Hh4obPq3HtAG9szR2qHTWFuKwsbSBen9KIhtj0gvVTnLyc74ZWEcskjLeAxiQacCh
JENgvHBe8mWplO01NcWtyo2PMixgkrf3AhOrg4VSHV+n3HiWbzalO64WEOozBVGZtYyngFlv949S
93+zOwU4CinSAkEWLZBLI7ZtJUHcsI88CkY0AV+aGd86Pp3pTb+2tLCUPHKHw4HoTqVNNSOFl1kV
uSMs5hkUsYQX9CPTIOkQ8/25jUul4lP0JIhCDYKCOT5Lof8DCcad4L/P4Q4JNjM0uqLrkRGgvcfo
szkCP1RalxLhsjZaedBa7xJ86EJgTZw6ZIwh0vBl8mZwfWMLio8yxZCaHYU73wCCAVOcivoYRO7m
KBL7ahZsl4Yb0IN+0BhGO8L7AGUABleM6XvzhvSMjpduGxGh+jOkvgCc+VKrHHHFxCNWdT/EgJD3
QzlwzooioCydcCG1XezguKI1Hri8POsYctaBjj0Ew3ySqSh5vJspYSsMknq+7NcKA0lX5tLP39q/
wLOr3NuueJe1tRIkFbKcK8g5BelnptyIQ5HvtOWrlmbEaKc4uEjTIHANOP3Ev4wLpBktsXsjYYdh
2aj5jk8uDOoqFbPvpUdBriC7QtbBbJrWTGrwKZQwxodpdxr5FGtOuWWFCsKKPVtlUb1FwmzBZR9w
gVSwi01AhKxV0a5yCcHjcw1HBa4K7G2Ww0eEKv5x8c3rG+GnMLfIs6lEk13n9NIC83QbQfiud7TA
jYangActobBZJ6W3JoO+TfrU7kUxLyUNJyfXpdB4bep+ZKHJsC5D1plSky6FWXqETMm0vqIhuvtH
of5wycJECIcIKmhTqMx/FgMf8MxhAypMITH4SQN0SAQ/ebYhn7dGDYJ0z8We9ZDJdeE+xz+7c2L9
p6tzd3vXo2kLxwHR94F7fomR7/LA2LvShqg8A6WrPvvXOcK6tP62dWcUjtVbKczMZ0/fxvmiPsLs
W1VedN9QzBclMJVpMYa3yGVOfyyc+jeY5lwx+JSSyw/s5MPepoCzGApX80G4KolQM32MRycNrF1I
Uyq+fxqCkF4hJwbzgddqMEEHSKaZscwoqPg6cIDJ0PfgtcuPU4U1lw2wvqbi8qUSCSnBHNTtijW6
hyS2GY8RNfQsAd+9FiocHdq9AfP8ZQygspxk0LOgjGjB7aKYkMa2nEEQPS4FXtSC1SIDbl4KhU6H
MNAltaQPlef8Sj3uG/gVJy7YU/jUYoN5Br9dp4xnjSqJ7zCIAq6NNCIUSomqC0sFqcG/+p3xNomo
PvzntcW+QdG8Z8Alv91R6RAp6nY0PbxpOTmGPBrJQOofoA39oMzTZKyxqcQ3y9Q7ZhZNmoo4bRCw
1rGZOjLogsI/OWIysADiSYUo10a1rFn9omygQnB6zhHhSGtDClCGtG84RQ/rj9wIWx1FbqfCYzyX
nDvGWc3NezEe0kS/1dRoHqstcOEdQMlzkVY3EuYc4VqwO2qrfUJ2WwknhARQlNvK2QTPytVRXbfc
dOd3lNrB1hi550whBG28fyZ7DNlrUoFG/BfKn+fV7XZpydmk/E+VRwVGyA/chV4Bv13076KvMH6S
p0OVM/fdFabA3o8kHls4gcr4Eki3zN1Q+xe+tuHF0LZeoWHlL6Mm0TUj6VSDq+pgsKpmcpKEh5Zu
XxqEp/pC5YOmQC7TAamNmuDjCZ0vG9c+jerOUDQ9sc/SVoQLFUG2oSDRUqi7KUaNsJ8mHGPUGUXx
gbh6d2n+Onev1nFDkdKssyS0vtO/ucLIXwAOK6w2NZ+7hnOA++IGBt2raSL8v+swHJO0nVt3+DvY
2j+/0yIWh4jF0unmTj/VZn9eDz4PHpIKvGq+mxNrkoBWHUh5Du7XaNxt+mGzd6v6Y/2eij6w4NBK
xIttZSyP5PLmxNaxxYsN7cgqD4Cz9ZZ6jesp8ew/VIRKXWFFkB3oRzqnAXKqfIMjMpVmB9mOjpe8
ld+h303swaMz8GxJY9qqMA3Eubg0jQdZxS8zAKaa0OsRspZ6Ndco9uW8x3+mwdug/0V6nAlA/RGs
TT+XOagJZnnWyeEifIbICpjO6Foeoq8dXyodhXyH/ln9/8EiueRF7hu3YcGyKozgeWqrSRxsjGzR
uc1xzg4i/Jqlu52xPAJnchAY/m1tg6rAId/lq8190JLri/1mq5nbTbdXE3zWPUHIaJIyL44dtYGH
AHsx/IQ22yMcEloLSRbm4efwv/jXySADGlmH/ciIPe6mm667njQY4RX77pN0H1wk8+FPIWBTgaaf
Et39j+K2UKx/shNy5WVLnVuT2cAKzRV3e0JWePldDFzeNCnlPO4zAxKNB7b9IwR7cojJrDRcETai
E5DAiVHm8ATVXJSesTWX6SeYaFhEJWnHJBby/Njleh8qkot71chREtNXvPrQUsheKk3UyLGVFmnL
At1TC+FvgXqSkWVNw6MsBRuvzhbfB9o2S+yDQoMzrHHUFGFw8I7PGLSykt2xKOhHOQlC5QTN6H5B
crV1GDIZvZDYVQyScstPNzXIfTMPlxsMLxA5HL4w8Z0L6cjmSNEbaKiblIWmj+5JF7sOQ+uFT/tQ
+sCYYT18fLfqR6V7J0lqNGZe/T6OVevcJCk1Znn/rsLCV4FDUEjbU7Pde5eZNqCkS8szmsOrND5g
EhEzBT5ZDy8G9GCmHZRBlOYUoSoo3FGpcnCXYxI3T9TZ0/lV15itv43tkLOQZkEHUe8r7211GU/s
lf01tw4pOdKRntEqRAHBr241VgmrwlZWdVk6+InrSu3g8H8EK2ZAsSd8Mu4JD6qB/LsZIslESiVG
4GoHIPGbrIMVU8bXXNin3RMzPWHQVsvbt8SdlgAuNq722oMmlU/zKJx/WkHUwPQ5mx8blZXtBhhi
8WEtVod8ShGYQtXr+ejAud5xqHCxASfgIa8Sts19/yivOHVvPNASIP0kxF3ZtyY8QalI70H4ihj2
17wMabuKBK87rdpDBr1rRtyIetUTRiyCL7s5HX9cA7OVR3c9Pd/vAT/NLP0vaA20ouP3Ul0SfkKp
ZTVf5lk453p4vde//yrlSJfjJAMuj6165G8rCDfRhcLKXaDJUtZKo8yMEU1GujEjKuClYaATiD86
PJ9Vsi4RbqZ7X40kjthQj+ZRYc7TLB6xth8PAji1iXEchCJubEKuM75g7jwQFIavWgC7W8pxvQNZ
WbrhnqD7LCSrLJRmetpkIPdZbCd3Pd7Qwdj8e6GraZO0M3a08JhgfnFYdL7xhradNQ/qQg840Drp
f/V0xFtoCzN/lWKC/k91j8Z5Ui+u6MEBeigdfxBLI+99UCg3VZQloHRcZLjq6Pk1N9i8nBct/Ecq
sq4k2k5prDcYOkGPlbXm1co2foePQJZFdC/LNHGroCOTLHykd9gTGD0BIb5/xIOuRM6Py01t4jbz
+5a4dTLZ1hIx5d94OzxxdDecuYKzcFTMfwCVggwbq/BVWH9N8qy2uH+thONSvsc+7KN2N5HwPjIm
XH0q7X40tq83bFDfSAJX0ILbHYI1i3UZws3IENSarTvHmkQx9zrV6RjtHhJoUcD2SZkQ8QKC8089
WjnWts9k+PQdmRUI1SShVxjNj5vsz2Q6evREMjbQKQBPAPPZmwl0G2cgkYWtuHG0OULeFDhYibjV
sfdb7Eh/sV/CMSv8mfaBzF8dAwaJLnFQLWZRpHfuWgOLORrEXhSwukd1wyegE1g+PTSPbJJUNDEs
2Uq0D5SWbDuVMZHeJXUO6Q8nDs9pZibl8Gm/rVFNo4tgUfEnDIiU2Soyq8Hj7gj3WQUDBzrzZ/HB
vnYKP1eSeP9/3oqFngNG2HIrLU8UWlxgZusmyJsTPE+8XqMeq1Mq+ZOY5KnJuWJZHPMLbIeVwjbc
Ax9PHegmUyUmDxcuyPc0U7T4JjrUgGpJCDcT819fQl7e0ctv4C2wT+VAvaakI33IvEwbrpbU5rpA
GLVOoznqiAlWy07R7F9y5v/fWvlyJO+Xtm40yGUCrGhWhniFL9dK7Kz8QUZpOiX/lEQVzK0QN7Eh
fxQmujtSoxsasVhgmr1V343vy4V8tw9r5WLLMHB9euOGVY+74rpFbSl8THLpXWTYMWwuHonTuwS8
GuwHnDbdNVIqfSs/oS3Y0n1dt6+2x54Jat+KHXxUZxjN4ddXsFJIqEPQlQWsquxhRqXZv3AdSkD2
PV28IIIDnQOa0rz/LTqCSwgeL+91ZWQJREAadz1BmjSB5oJEHGSASjZG5wJhEqL9JEagGzZ1y5U6
s9C1wVhgCY5JtTOxAi++gsB6DrIJv7Ply7BBGV7E5cB+SLzzgNZluMoF4/V8p6pig5hO+z/uytgc
fmio6rzPJtoPVYKUkDSdGKvydV04fejbPtGO6a/gLr3bhMHFFkRu7lno+yJKE2T6v4LL83Tm8k/G
kxtdqgaNzP2OInwYOxWvSxBUsEsowQufp+PjS9XcXQ2qayn/qngKysI2uKGmaSak9Pz2+P3pjEQp
BvycZgBbrdCExFHNp7JPQmOLFsUYhx+JN9HuK8EToUGl7yICiBade58tlJdWD9TSIs6aS4r3/0d9
691BalaKY8evNAHXyGLGlSDPyDzXIge+1dL5PwS2H7/N3PKSNkDGXtfRf7UVRcXK1oppwsuDs5QD
W5Om2u/1DpaUfpb7fkuTaBXNDJVSrV9YLs/1btjvREtjEQVf8piJW+Qh4vA1dYgK6kAS8iuWcHt0
k3guOgSG6SH3xD8vTrB7ljoGvCOZ7HJBKmPP9dJUI86EIFn6PxfTG2mIkUEIkV/YT6WRAFea99QJ
2Xt30kZNOwUATb2W0uiUfB5JCK23Aj9v2iEgKSa+60pkao5lwlutuo9kWryNlS77FHh9nvghB7Ov
hW/vNvH5oMCpdJ5JqFkAO6f+pN0ag+gAgJ4VpidCTPTHGXXpVjfUwL82FNnv8SXOXwlsw5Ke+7Qx
3Nn2SG9eypmgARxYz8QR2HbItIdz1E3sFdpj4SniQfbp/mFZvindtuQtkQL3p+NPa5t9RayPl0zh
+rqvBmxE314M0ELmZdWAHvhpOeAOjhn2jk6p4p4YFLVMBSRz4+UEdnLS7+ikoMIzUCFBVopu+qHN
DG+tTEXdF92DW0zZZSfVYCd6ZORx1cLUC6XpdJ5SIRspL7PTnn14eWskFg9oQapWCN9c4XElJH+r
wJzDTQBhZuT2yy1WJe/muEXDY+6XQjGp+3ugAAo/RqCOLI1n29yk2jY3RbzPSd/VO/Y++Aee9605
YxWfgiLQ8lOLnwbFK9hqBGVWXI9quVO6B2nHF+kOJw9c8dgqMrrs2e29d27SSzwm1/SmGgsbVdfD
sFV2d+RrIqMmbidQt7eH1KnuLKqzTdiW6z+sj+4o9dIFwdroHr1Exx+RJQKWuCFYMbnudI5tocvI
zCAdrwgTYm/en2YNu0Zkuiptz3IdduYKXL3yIKCx0ikmvp2CGui7ceMDbfFFyjyEseYzzpb/RHd3
Ad2Kvkon2yZ1Ewwn6g+lQG0Urz4dNKMUDi439BGPTzQAeSslNocGEEVxUxbSH4K/UwrhLfCGUNgJ
Nr98qw3q5d1Ca7DWBihArPq6BVf8AFn0m16nUvnKWRG510XAcn8iAaGbLnF2KpzDaMck4EQrMZm3
MTN/thnWIN8sZmIARyYB/SChZM+d1nFDq8W3NlNPU0cYllzrTk5GW10o9PSqvH++An6WLJDjFT3V
n0I3wIAeW3UGrDFIotj4u4/jFeK9mT6oQz5E+s8Yb4+VWNcXVkTrCsYEqBu0cOsdUoodACv6YwjH
H9M9jxNyeOk3QRyaxc9lnl9E0RNCUieFc9nBIVc0m387wjDeKRKqBHssTliLqaSD2AR+fIQo8YEb
9Uy+BY4RVaZSRgRZi4Ce+DmIjlyXxxX/9sgqdkbgEBRJ5y55G2nQhFTxXaY0KhIoQyBnt3MvsjZu
YT+45ukYb3B2OVt9Tm8PZobgfEbKwTSAyYkxMdbnAjMOLMksmYPTv/hyfG+4PdeXL5R7vKLNEHua
bbpDQ5BUXGpgLjycdQVOX4ZpI1wrvt8ZKgbCUFDNqCTlM057927U7AOjRvQheQxNEM/Qkk4iNbbX
bkferre+gxNM29/Pfs7/SO9b3WCw81bsRvyJf42G2AznRMixawaGAUgyhpt9ExGGPAQ2V3ayGVCg
hDhd75zHJs1KLJg189hCo2FpLFCylBwPXsVDhmtBEK+a5GF45whHJvq2hghFIP3nVPDcDIEoDNPH
RLXfZOJXdo7v2AlQxfLw71wCkKDVS4YEBvXVK1dH98k+1Y7Fnrqvxn3Em8clrRCHCcXux14gZwcA
QXJOJNWB9tMejJMRrmlP62n0V/q4325z2gRgdICv+oGwLuE7SAaG7P+YKkFDmxDFrIcKwHBH5hex
99Ephja+XLuCUUaiFmjFV7EbtyEQ/Ber2Poi96N0rpoafkUcHxEHaSIW+dp/ZY0IvCKI4Ja5m7lh
nBwneqpeV4GPMYVxrUDLbMRc6zKx0f1BIeRB3XheZ/4vAhdwX064Y5p4oZ1dCOvMh8xPlCDUD64T
pLUGo/yozrCMEb+tWucF3WzdnQ5sx1R1rvhhm/H9mpAGNv93XEvP3aO19DjebpBGBBBTw+EDRH9R
5ynQ85A5/Kv5Yl3WW+Y3+rlOZ4cfh0hWqgBrLHD4wSRwj3XyTB/t4s0MeQbUpWTefpvJtsPrF/Qv
US58rzMQDuI1iCIWpuQtrAZ3p9dbmaF8rxfDyFh+Zs//gTJZe/kAZWNkbS5qliL4NzWREtd72iID
fcBdasqFzcYjhmCsSB3fvAqfkbzkDytLOuXWWBrUvBQg5Cp+0PjO4+qvRo5GT7LRa0Cn7OABcXbF
4VQjdnoBWzRXsCtVVhvewwNR0hNYMyLBhZzuZBILo/cDrAYAyt7tC3nkcgQMQ/MU0juzBLDbFQvL
uGvAp5BQX+C464XyLonD8Z5XyOfIeCTnCSalH5rpgcHVLstKIBjhwxCtblsmk4cEgbSp0y22yTBu
VA8eTf0Rc2F41IoDTPbgQ+CGa8sxvQZjy1y6uPUi1C0PYYbwJXcVPNxCot3A4gYx1teGGGwm9Rx6
n1BNCPdc+9Op/XWp5xw7DGQJx3W4DPYHlWrlqGBhNKTHT2FY/RsP0N9nxZkL5F4Tl9me3i/vYUgV
Q4Vq3IkZ2MTJt65GawSk72yILBySqbAeyckaFFfrJFaXFRzM+vu+D53ZujGoqgIt56brl0T/mPvi
MijTao1TP595lj3w/GySM9e/ykvkXt5UR91g5V3206WljJzyVBq/0S6lBHun3jUCkNVYXvApfzF3
4keYWl6zdClJp1gu5HydNhEWODHB+eo/J/tk8I8HtyiKJwIQjTFKPiGX5lnCibUV0lkPx4mzxnRN
AaY6RRvvcgdxFcW+UWtkD+6IvAIR39lCrMzpzWCNQETQILzszid5nFqn32EPwlHtbNnncEWnhT2r
Mqyo4Ja+4C0JF4S+x7HrElUeTwZLOuzq+i3vIe8sDyRLSoiGm7nSR7ui5JFOifkzUaJBuafscdWe
mRy5NLqx7Qpk/AGGZInuGRTD0dO9feLnPo0UWmea1796M94mvJpSJBo69eB3Uj8LlF5OQvMfYZgw
plZgXReELsWKY1d5d+UCnTwNm7cwQwDLpR+Dw9fhBJMoJvSBxhdHnamXRZyvoswwriBlwpk+kc9o
faw4tcjorM8NMpA9jJWIzYef5GH6DrlkXS5sbrghpRm7+1xEBQFgWpqkGbqYqiWnXrnbWve3XAW+
LV4ukL+G8ehyLEFx+4rplBijrHK+X1MX16ZYc/yHF9Avdzhmc+LmSg55qP2CvGtGUZTQ7nJhgoRh
UOrRG7dhN4+GlV+Alva7Zndlf4on5SkAuEK2caRWzSNM/0a1nlljcm6aG2INYVBpdGLMC16BuTv+
XOJykOP0JYRqdUcUTgwH8GBOulSBXGlR+FLp/ddkB8xLLCumyXqZHUheRnOfjEdTMRx+ngsTYMhE
/0tAAX77/+cmnMP4qYAjF7C4lhfwtdkmb0ZqMaTacS6sWF3O8bcvK128PxS2VR2Ye/4/Fm+Fvz/G
6xTIRJNHo9S/zCK20SvhZQ9jnjjr3zIh/zqmwKEQC5qQhCgMqi8+4qDdmmgA9XdV8i4Vm/rF/FRo
oCptvTyIG5ky84XzF8map1AhBD+VRrMYSRyKLtRGBz5F0WafeMzkO/T0h4vpgM2ueObwLEhDp31T
4fLZ9a1CbxJP+VZwzBK6BUVgA0/aNvfDGZxfHPZG5prwqxfYd+DJwatBqmF8rwt/MucZcup1S+qN
xPmw21QNgrpC69MlDJTrnl8SrXGYsZSCy9Xd1263Porh+WzprVGoiMqvdk/zfvAKyFOKRg4AtCOS
SKPje/R5JCOUQmmhtV38qrafD01JOKCBAiNMxKdGs6sr09Nk1BiN1EyLsuFDxWzXH0NloNiQlFED
KI81Bc63QaMq6c/4Bk0gKSDffk3e36J2djUmC+lobye1C82VgJ/iVdxFjGCT8OHB2TqxI6t28u1u
nkFOI1ykozD1bUYHezD7anE3zCU2FuMTWWd155M4xAFSgLlR319UYTFqYWG/UYZWqI2LmA6KWXHm
Zb4Kpvt6pnIL49nUetv6xCELGfq51G3l8jbBr148uE4VhXWbmo6WfX4UERXDHv7xzb6g+kFj27tK
4Du+tNjlqp45PylTP8zYkVB/MaE30PK68a/ibdRStu7MM/ugzpkeFn3S/xEzRDMX1I0HJA/Gjv+A
dqMkUdyeVWmAswrV0C4GKHMN9HOZLgpKLiI0UACXbB4SZ0wJ+F0WKxNNcmKpuJI3VmWSuUbspNBI
UlI4hQVLQ5OX38u/TwKIR29Zdn1YiB+/mUY9KPgY6BsoTjmVU8OPDYKuW1r0yozc9TQxkBKce/OZ
NuV4IskJUc3RSzflw0MAxSkUjKsA2Dax3ZOslaYE6A1TuWQRIVrZJMuVR5JuY1wBWkSvrqvRfKK7
cjaUbvf1W3IlS1/YrG4sNaBJJXfUB6IrxOByuZkX1IY/qK6MA/8V8GUgbuneidgMoXqZAr7K48TS
DXmpPnkxwYhocgm4TF4EqTM8LMlSRpQlTAzZu9361XZhuh3uu9iod7eBBIJwuR04mdW2L5MWfRbg
0mJ8KK2wQFHfvHOTDoCgwDHpfP7vBy725tIAZIUiFtlV+QafZmyTFhwdGAPXKADGopMMLoP1CEdi
Aqz3NnA1kPREIsfpHmyR/rTp62NCobMC0Ft52yEv2XrkFvUm8oBeTZ+LL6gkjB3Mom21/eGXbKiZ
Vyji9yCdSs+hB7tcvobzsETdRJo7vf+v+mzcutDG1wFGRu+MVmjsztyKMrV/OHhuBuK5nOB51Zaa
jW2dv5txqqgig9A/sOYuMyWNnB3YtD9mhOdN7DlHm5pOZpj62lfv/oAfavkf3YWgziFqPW9OSNgM
yFwlJcWDQYDcBheQxErnVM4xzfGQoySSwa2s+zmSt3vv/XUfS74oM86BC6tmjPlCHaCzLE8Pb6Q5
L91MWvXhYdTK/J6tkm82CL9TksQ/RErwwQeJmpGQ8SDtznMkKZC0lcPFMiGf7pBSZwmoAcEK77f+
DkajgbxirprJPQTYw22YXpl1NIWeOhL8O63klaB5UPoq9Xhl6PbZwrAZTLmzPm0SlBNYzRGX0GhR
jTMQoBbu437sQ89IinKkJRMWl++C3gu4I+HFWeGVCCzhraJKkFDruKVJvtqbxwICUc+i2Rnsdjh4
YdXd/6iQRrSMHQjTGVVHwh+SGZ0rFJXUI1BYj1rjA8027ccaaYiReey84iWCVllGWpnSG/fZTjVP
4LEdY3tBt7nePlf+agxHD+IPwA7XDGKtRe77ohSA5IwQ4Ed//8ZtA68TNyzUpbxStAWrI/u+fFgh
3bR+dqN4/7vlIN0UZZNqpb8RLPQiknOBjvnSzGJ6wwfOBHsIa1isn61vGOijwJS8u8bJaRYPbsaP
jJrYPe8N+HG4KcYn+8K24hqy0mzob697wdjkhkg4w9pjOpITn+f7BZ+coZz3GZxC/Zlcjzb68kQC
PfHl0Za1OTDyYjuHk4jn3yK7/LlP1ynv6bmoIVwIndPbhvqwcgpYmM83s9dvDom6a9vYbr4Rx/LY
/8X5r17gqk3qBw4kwu1UUVT+7IxV24P/S8PsptTBGrRL148uk7wvTHIel4wLiLwv7nIAm77gSDQA
bciTE99zeKbYbG9nemI6wT3ndw91X7G12hs8vx7D3Y9aDtyq1xcOIHP6nj3h8nulIkmb9vqoIH7J
dzIBtTTR1efDnvH4A+peci6ZSON48yN/f2x6POBqiMGYJ8DxtpOP1V7BLKk5f1sn/DcKAV9duKFf
ttuEII++OIT9XWji86+SmsVYxHGvYB2avmGNhIkzqpcCfDyWZ2U2XSjoN9yrY14ahLMnfJvaQy/4
f/K6vbLBa0jPF81qy7m54qzKe2Drh0pf6g0umnuDG5xIg8ehzDDGTE77OWNHryxd9wO5xBX+wRzq
flqbLJYIZhcqyXEv5ginG4OGs2a11y0fJ3wa5Peb/KXQOmPqWLm0mqYDlXUXzQBwbV+6dTU1TY2v
QlW6Gu1QmWqGmZZcBf5ZT8LGmzSabwLriVDvEZOZvwHcT1zp91/hMmstUBfZWGOJjsyDKs9mxTW+
eaKeNbNPQ1nyI+hYh6RUVn/9C+dmVt9MxpucG5+spx4QwZxRCvbku6QC3HYmSMFpzZsLe+Aakqsj
pCgLb7G8JjmAYBJEQgYEIQkzowaY7UKVxep3RP4Hp8Fh/jrXAiCZEUyc/ruO6wzuW9jE9B7VjCw3
4bcAJReYWjojZFDE9cagp+UUZj7TtR0cw2H14jcyaLUU+bS+HteLXVcLJo0QqUNagJbBj+e22apt
l46QGxjSyoYMz9HSofYVY6vjPeBuX4jmYiIzOMO/nek2rtaodj2V91poWVp6pnZ6KrCDxv1DS1Gl
NvwFSPA+fl7qKL+M51cLohYoxT3CzzMV0sAtbuLtLGneFESckdPmEScibzH3btSZ4I9PbvOyalpg
lSttEnDz42N7nKwuSZ7rKe9X9QNu/sp/+17t2WObvJ6oRyB6fnUlBA0+gOdLjJUHOKs2faNxSP0s
1ioucPAEtpRieWv5eO38Al1Gwu/wlIC6225cUJmEH6Mtixxobq5JZKCfEcaeK7pw6LuoGxKd+jcB
DrIHkM3dZ8cFAB0QaFW8i0G5KKPruXzVX9MHizazj+7PZJiqgiCPSp6DrDLGCN/lFoLD1ALGImk7
kjCULTH53NfvIe6Iq52w3wzfn9QENIRq2gWDh/4uuCCH0ZUB8Yk/Lgd81C7BTFuKm7XC6Xss4Mvn
U+3pkjyXhv1UNjj5rUpIcgbsvI15Xix8Kr3/6CpZFlyb72rYUJWv42nNrcExK+Kv2BGlISUB32+V
SyFb8raCFXWhRb7GhMB9H7+wqiioAalM0ZSQFXu75r68bAtkfesy+zQF5GcLT93rpv6siAOmxPBt
EX931Fm3OQ7Z+7TuU/ob383Rqn0pUUgXJVWNc5zTpgQY+iParc110aVVfd+GbipQovHF5jsW5SOj
wYw+2cj/sCsYPCnle4R2qWR3oDwTloRy8wGNZUXskQ+8fFSHKgKfA6MzBUHGIwBZ4HSugpWy3xj8
nvA3iB71WLyO3fXPQvBdr3QjiBs3YyCJKVeh7W9xZoQGBWsoMeiDc5ittCMXVPvp0COc8Kbdunkp
GRUY0sWxx/hlivlwlAfDiIbL3BmmuPDBy3eGV+XSnZn8vWyXW0EWJl1Duj6xEFrd8idpF3ypn238
oz5pUnPDXgmq8BhVumCVyz8rsJ+IxZCiBLHEjOkUwqI1FiKEqPWqgAsZT4uY98wQH5khmnJwXinJ
hReSaieiqYeseTFkATMkO20UH+Y/qEz9zg8HPPTFD/qbdNtizBcQ3XV+l3TOb4GwK9tPzvpua2Po
l/YEAep9HOJBGGBsBgivQZke7TQJylU4CtWRKqend89pu4zQzILkQ9uAHB8qJF088X9YaJoWtLkP
qu4A1wGTzggczwRRESTvhINuxsDlk3xsqwjvgYv2bSzZTbzmKUynLyqU9eI1yfKWWHVqi2l7i300
gRJ4tRLngX/O2o+ZpJSCjNqNmkCfUvcvYI7no7sYPneR5GGmbDv3eDn7khztIjkWuGtkg9yVauL5
NxHGJ0W2ZbNrfvzMVkfimzOtl22h3/EIOmmRda+BZUY/Dw1Yd//GJlcxn9MHq+foEM+teBeG8rLh
pnqM1MYm/VfgfqWYNq9l6IkSQ+d3P2+5IGkGxk2eZxtf4avx0ZZVPOfIN/aljYZ0ryKBJI4Wt8pr
nyL4kisIswpOu1m/5f6c4kb6OT3GLrXj9+tVwl3rzXgzj1HgRoxyRXskp91mKAC4dJGFDL8lg5nM
4ntjdeQIg0GByE0reLjP7mfhNJzrGN2JVUjkM9u0u3nagwVNBxGuxArvr3TD/KKr5nYGWa+TwmRD
fVq49ru2ZyQ43Nd0LCEv4+VgKiekCXME2K5oZfM/cKbvt2n+Pf23mG68nTKAP8i8lAMQxE8aCXGv
0D3JfNJBqM8pln1g9/9g9LsY1k6XY+rV92K9pfcYZg3ronmhFZ+xwxvO802s6MZKXdJxpq9qI3di
qFOQK2cD2D9jG9MmV8pAd49iOJndSuRP3R3tG0s5z6NT4B3QO+Ae8QR1bozADnR/0/pytSr3DEJv
azvjfsjFkpEtH3M/EOR4rvJYx16zatOKdiJ4gMksAfiMTDWoWhVOFC+W+sCGpWhi4XaW34UPSbOI
C8ISSfm1nCNdbksJNdFTWcZjcjaD3OrMU8rQ+bAWmNhKuSW9xgjFXU201cwnpPLW8LZDTU+ycVNH
6HG/3dnG+i+rKSReuj27to0SVdK4XMqPm0QNJ0ZbqVBDoAF36Mq8nt0IrZP2MODVAhbBWrX/1IKH
3Vu3Lum8l5NzyAotxMLMGx7H3T/9HytkFzdotyrULqKQQuT+7nMNIQ+MvPzfhLSOSch/sBaR63FA
QUeKxzesP0foaabdi/uk2/3OA3VGNZfL0bSDe7qT1N9FoZG88Fi03A/jR6nPgWMRr/F+GZjm9L34
a9UV8TNmBmYoWBOzB1az+Dg0dYC2Tuk3HiagHXkOGxRtdz05pE2oG6GssBQHUx8abDJXX53yIJv7
eTj/SglQyn5DKAff3ggPOdnE+fMvPYOUsJHkOBaLIrbrNW0Qn4dyxPLs3u8PuP76Yc+2yJQHd9rN
Q4ocPXkEzJabyHilQr3cFLw9Pe08/K/6Xt+PTysew80z/AF+GzxoXvD6MxK52qlEKrUTXnzOvYns
x3PZquTN3adDUcu7c7NxeU2Y4iiB2DUKZ3Wc9YjT+etW/IZhRc1cVGnxarzXCR8eEZCWCBAa01Pf
1aGLUuT+Vwj8A1xLd8CD+uA3AWY4e5GrxE7UXP20+8uy92RWUrLjxySW8IjsBAM1pANAsIMIO0Ue
M8eMvLZMq1nDdo29JDcC7resm0msgm8FLRWOb/GK/bE61GVP6fve4FkVfPRnAAL7qoYyvMHDXbIK
a+rwAX/n+EvTBTga1MBrhmaCkiqGBn6HLMYt3IwhkNbStZv1g7cxkjxHXRU6FBTen9l7l8qOWkOs
DGpOytDV0SQbLO/qLfCUABkvHDIIeGbftnGW70vhNlUmSGCi7ZYz+gFvX1usXR9qDkxpETz2VSNT
W+j+L11pwUoYYbCmjF4HcdCehfcjEo0bN5ttCLD6SihnV91LJINzuHfOlOzwr4IAr9oLWjMLJ49y
goOUULoEQmemwl60rUGOooCn6AFbbLTQkNxkDagVrtadC8+lhujnGTWpMFlTIsexWeZqAbc6A2Wb
Uy+fU64O/84Mq2ERFIQORbVM6QraKL2zJ6FpzwHNrPmICp1Nw3e8eE5XBUuaRAjVHgppVJNRSG3R
hPTKqYh5zP4BmNPurE5PJlBQQwbFfqisB9reP2M+laHxVDwA4aPiGKhihv4boUirPqaDDELL7fI3
/7V/gW+R+cpf9M0D7khjV24r+/ouepfcV2/rMokx4Cb15oJvLRblvRxlye+qv5NpM81pIfp14YPt
fS3KHPwujCQl3cfFyHN20hGAf2cgVBtshPFfTQ/+Kz+mGh96IZeDMSOovHMgGgFcfz4aYeR4Y3sm
qvnelm2iwya1RVN/boSSSAL03M2jhbBiXpTtgOVbJk1ofCi9Z+tANN9XXrFi1ALx3UgLDx9nbrXJ
O116GhgM2pLk2IxtSrmUeS1PgBo6/0oEkyzsWkM7J9b2L6/mKfsSPz2bY7gQ4Ehv8IGGkUc/EhGg
OR8CcybZu/E2s3uQHabgsZZQn25rkW9pG3bsHJeLGwDmQ2JkX/oqA+Hl5ORDDqr2AOlJvOpgJnoL
jSoWo9N9QyMCY6BBS0mfx6WhrWttiF7ZWjuzRJI0C6pA9TzHmlmlv8vuAqQ3+zXgxXLRl0ON8d60
nxZ37Nyz7kZJr81QuSBGCH3p6DgnLMcofKVt+LUsK3yHrYIdHVUuHI4UTL66SvX5WAh6XOjtNDyl
EcbLw4sqXpOWckkjK1x3DCezUIX7E+hVu7fgZF+tgscHoeRxi7tGBf6BGKoopoC1EMrI862I29vM
Egxpa+pj6cPAHr3bh1WB5hIbO9giYovRLZZ1Xjf/QYw4R+mMnPcdca4UwYsxQb7Rn6ghlk+TXE4p
ia48Ib3Vg0vvYtHVxLquIlPk4D2Nbz1g79Jy+BvqwqX7jkQp5R+hxEt2e8MBNf8yiAiRuXYyqiMe
DUigxtB0OpeWvS3yh2rEd2KGqKSoOihGoq4DhGZ3QIlvGLrlPDfONumc9IKhvOSzmlBvWUD2htEG
NyUnHQ+78DMR4Fp5HW59TXkdjvhoz8Hz7it+xwpWZk4QbXub2XqLwyLRZyK2yDSw+wtKfsrDADZC
Jx2IDtMnfmeyU5zuoY9vAVDMqaRUSoEm4Y1USHCT56sm2vfpXN/l5OEQMGk5yWq4PTH0J8JJSP8R
VcXDuzPL217QNy3f48k63TrNw1Uey0LrBTs1A70Oaw3daq1ecugGm4bCRaOQJ3JqGmeejDBbvImz
z6KgMu/TqW0uMLP5OjHIQ9JxTZi8BH+OUn3K5kNp35dgJSLpJLyhsYFNTkklUhkJp4H841d/XJSu
/fxY6AaAP7zBCpoh7L79aoNItoIglhP8tovPjsI9vbWMv2Bq/StWv0cUtUjSVZ33wAYjiCohJUGV
1+2S9e8p8AfO50p2b6QW1o4dpShf1dIXDCEVVPDEV3Mws0ocOnwDAXe65dw2z6dMgfBox/x75Uq4
sZ7gMpf04FTVwtW3940uJI0gDt0EKO89J7LAeAYYhBbwOtKDkRlsguhu7ysYkjU5ctAqF4EToVFc
saCKV8+3B9OOv3lwerzbDfSq43ycT79fpPup1Qgz81dMLNkoykmFHFWLen4gB3hV43acI2lyr14i
BmkCwvuNlmW9YbBes2R1YpnaJRAqf4mLUF8YBkVoYigU/SWlnEU4UsYiLfCA0JD9yH6b4kjqLsNQ
tMfZMDROYCg1Qqek9GTPAY6YBzHl2gUHaTmnf384gJd/5zfPriGjfPSmH5rCxsWThvfv8nV5Mj7r
PyO7GDda/y3WL/+g8JbwV63E1c2XDL7CjT6ZFJUgDIeKFGb8iahM/L3yGM0jjDHDyzI//r7wrmH6
ybd9sAxO41WXPGxn5q0WdgGTBw8ztq1xrhJZkU9zd4lIZO/G7/Ow/RW9Pg/wegX2dVW9DNI03lbj
8z3kIAdMar2irunray37kOeeUrdop0IXz+6cozVMZDu7oy8C8HyPQ+bUHr3aX8HkzOUZ+Rb4kY6j
27SEJVevO/yBSd8utROezwdegRCcgKBamue7Q1H4mXskUYFclYa8Qc6tX8iLqlDv3/hYqpk2ZrqL
AycKzciJ48chdkmcHHNcaXtTUGWszxeV/9odw5zNW2HXAzFrN+r6hgRpc8UukoXd0oYfwanNcNRn
QLRf78rn7ghVLYlHUtHkNNFJb72FLf72ERLdo2vuVA4tIYQhPKedpDe/HzBkxvLWCXGUF9ifSBfm
cQ2yx0Emn0/NFCK4W+svIbgSyk5LBHHSCvnr0jAi8yTzW9YscXmFrYZwM2xrUE+LkTQNmRbHfBJq
zjS9R3YVzDObz6BEkAVUldAJ1UcC53D/8RAx/tGab/cPv/4OS7WdbUFm+yWzqpIqCIBoCEbnve96
zQLEhzqJTEtlMEE7zpGauiBEV2EZilvPOTAnfKEN0Zqjr9cmiDw6qMtBtclrHKlxT+1LFvx6nmF1
4svVQwm2C2wg9e9Ohwx/G8Di8b+hKm5iDXPYy7k1Nt3SBhmro7Bx6frGDO5Qj28RnRzuIOCDHQXz
fH22JkEgqyt5hA0HX0rJ3NS0AzSEy2zUxz3JNBmqSac7+vNMCYBt/5/BauMqgyDZcWuVug5pdoIK
V1WUp/p1xulYEcvEo12kCZpllS+6cpggk/99f1mXhb2ZilQZhSl2Lbf2e+4JQiy6Ro54ebcGbhWd
qNURyMnUKFnBn6cG9kaOohnNQrx6XM/KVUF4X8uslVBxRkMmJdLTGttiV8Z1Kyl5/ytuf3p07oKa
Iu9hzTwgVZR4kdHtdWtYDRg8iNfQVxea+7Wo3ZB/x94rA99BdPobZBGtHDrYfgclqKZj4hpnCS0b
l3a22bTzh3pF6yzsma5A3+hhTWSxxJXbgHFK0N/XSOH7Q2S8CJeyjnkGzyf/rQLNjB07XFAFqdRT
e3fg9YpIsXmrcdoTv8I4jnkz1x8Hi4q14h07KQYWzwRpBJ+MJUjEviB6MICLGWtdpymHnub4mxAY
AU7M2Vm8yhZNRc3VvRY3MNztN2DU3vnJG7SVbyX5aiIf5VoHUoNLUF8nWyoi7r2yPaAhk3MBrYFN
Li1zFQG65TrV83uz4cpN61zsn0VstQWNmKI3/QPmWiVHnRCU61RbJXlEkNND0x/TllG3J6yPotD4
ZCpuTwtyYX/gf7EDPoPjlKBXfA0ONUeEeous3vxnJfGKPVZu/Sg1z+HuWymdJTsIHGm+o/xu9bTh
i3ErfC0f4L8qZvGHRrkORQTDqwNp3fpMTfrtkNmfLmn9YqMfaQ7djBp6o1MYfScKY70WI9v7sCPf
c9X6DAGWT4UpXshqpFXG4QAqkNAlKFRpCJfzcuxuuJZlC/wijSGzTOLDpCCHfVqmX2kovQDHp5bp
pZwMak+CLfLYHauWD3y/2cBp7geKDJShVTGj5d9jUBrSP7bYBjPJ9/YgDn1FB+A73DVbh2KmIAbW
JXNv8rrdaj78RwJpzk2e9vAAXeSbqojw+70PobNwS9FaAUGOyz9zvWGX0x8HL7776XQYi1d4upKl
v9rTRJY4WICY/qzMrL678sFhU8hQk0Rr8XKH5W/dBjKUJazH2ZPijBnt+wl6gd18eYMR0p2dggC/
QhOQATrJYrd/F7NmVpdHD778TuBCQRItZYwgjYMM3KopyZp3ECHahH9dW6cgXLmtxenyij/SZPUV
A5gNt2ouFp1tMHhMYFfQB83p1JQBShpe39OJ8kRdn+mZszqbFYbHtLBZH58Iu1iTaUu1u0+YV00k
KcQkLob+zOG9ca1HVEAq99O/jK68FKPTwFaisbNAQ/clzCOeOOV7vJHrkpL1bXMf+ly+TzB1JBl1
RZEdvnPS42Ogv8AXMwmFiiEEgdqLMM2leGgaBXxdkh2gIosVcWdROmX/ofQ8xNyv8BzXBcP6aGa8
ELyYdfZF92fynzo0/JKy91v1Tl6pY9s21679t9VW471uiByauIJTSpzWGS8PvZa0zWUHocGTjwrH
kk01f3xyKBR6EL1vaRN+t0azdnn7PbHbHH56srFawxUbNiD05c4aHu+kq3qNDruKuP1ySXc45JkK
7KUqFB8ZJUcrChCTFThtddVLxrZNNN3eDoq2NuSjAKXCEdNZ9/RseALBOznmmVJe6Z6lsrY5l5lo
qqwyK9ow7x48OPoTKCk2LcPYTgsxaL2VaW+6SCYs2aQfsB3jCOPNCOViJi4FOIqHCWwLMtiWX62/
ix1HcM7K4yT0rp3xTZWIGzgXXxjF2NEVEmhSyVfxsPSBYyRWfh78yEO1xrF30kPplI00j7CAlq+4
8eLqxMSqK3L1YpS8g9U+AF5pqEIdDRNkAx6vW9rGqXtiIeeDmLHcKajEcDJJ18jan6dT9v3N1UFN
SDBtWpTZeDtu/3WP2bFM4V0FFiY4oJzHVvgQblSNalAbx5o3MQ1vstLy3ieJjdAI01WJSz4IPDVz
YJQaiBndQPN0J9mDEeUCkgJwrYXnsS6tPr4FcCNGCSDdtE+yrd4yPFlOqla3A+BHOmbCBOuUawMz
2ZP993U1LBjESqWi5Oprofmb1kKxAPJamSPv92VmJj6V1e9Pqwa4lkLmy9N8/es1k9X8cQQ+s0n+
9BBKikhutJ0eNsu23WxAeCUyrHFnzjmk2Iln1s6QZCrZMyaxjOP0/v800wUuZLf/DLBpMemtQNYd
rkUUAU7latT7VVlOcTUVwKkZw1G7U5U1G/qqErgX+5lGtNVQ9BQxXBzeEtXmTOzrjly19W8jg69x
4/1bOzLjOffh1mVaogPeIfpVPjU5iFnf6KZnj/1xm0Cu5RL6mwWukfdfI9ZN3NBLTpHk5HRKL0sQ
P1XmUGDWyNmWmfg1K29YKh4hLL/CqWFA+vnfhxjlcOluE50t6xxky++SnsT1wKdwqBwPgkfGwDgl
FDwQOkhZ5g7jP6/KjIEx8fOof49pQRSwO/iaWViYiYmH/UBJ1k6sbCLzcF+jzv2Nr6FjxWrzAhTz
iM0tSNkwd4UXLMTyI3lGj7GSnk3HDAPuSRB0VJQAyfeCTcSLdV6koNGGzA6lvRannjJmr0GmOdBn
haxM7a3BIuGcGWpLqdnGqv0uBFN7X7CaCQLj2YJpBo6fDLCwve5fSSxpyyBVVP2gglmP+RbxocH1
AW2oOtzbKmqufwtQh+dOHftVYyZFcvAeLyJDeDRG/JRoWEZpDQ20JCWjYDJj68vobhq0Hj76Zm4m
BvioqGpM98tRM9NNLzIbtt1boy0G03Iz82ctbIFE7QDJvUBpBcKktPH8S5VjeG1fL0ZrpwO+sKx7
cYN7LX7CZ1rIsawSOSzgUtMnZwedk/FaD26NF7HPtXs9jADtzTkhTHFZbX/yV1g6Kf81r+H9ilCj
DTNzJW0bkYKnu3OIkFtz01oI0WuBk1EcqxZV7RGlgpZ86QP9hAIr7OXo3i1fbdDr1k7uUt7xcnfW
CX/ef4MCZyI8vn487MVuFUjz7ku0WNPX9vZR8idrx508o87cTtA3yv8nR0gtW5ejJTu76rLaYWgO
hHbgR0o/W26BPJok2unSlIRN7TM54QrxlqlsEQu/9YHExRNjESCxAywqpqcm0k0FMHCI9E42+cIc
Z399bbFsVylIjvdf22jUpf/mRmsAw9ulC1QbfifT1ArtlNNNT56V59oUUxtVk6XRwAzSCrP4k5MK
DsAQx1s5m+JSKsQCSLOFn7Mzk5cstheg5MQIWrt6cqGxyJj9ksbVhy6BIZ4hUieT6QCvcS5n/5f/
znaj55T7WIi1t/LjjLoFS9NeFhFvvHDqIdQmMCHPCHlgDBwlado5qLRdd766/5Ob5prqJln0V6X5
BZeCYEEvcov+vRJpSLJWbdaS184nPjHt98Q9LiukTvajrFHMlKq9YEeOkjFxUfH9jhEuRq+HTHWa
9S+Okt4kUl/tXtQrlItMEzxra/vPtjQnvSSCruJTYj6ddnB5zaejftKHr/YboO8B+ckFBKK2wMRU
WDYOprsOgTZ82cTbU+i44b9IhSksTJvkSa27YSGw+fWe7srV4JHtZp1GUgpA+tkvSWZSCnkwsLpx
S+JSjUI9C+iHka+/M7OY1ZNDa5ca1hSqW5uzWpXTykd3HD8dBfVBwB/LUlyJj/7mlhGnT+cp/UJb
FBtWXpDWgsIle8Jv6ZRDRve5ZD/I2V8abmri4lnfhZtcaLLFPY6XPCz8RvFtD6ajLhtFHbG0dwAA
o3J13oJ/0E8Ji3oKCyjiyubIwsB/eXXPGAFkk5pwmRfBorfyt6fqZjCWaNg8c4zl/N+niT17o/be
kUF2KsRo42v7SUwFPKPepuv79mOge1XH0PfTcT5Nx/iiZswmbokAYZ4EV2R/zEd1tjbudxkqCi6+
0fSYitUiOuVhrziJAHRQ+FGmTyRnaWjhx2r86F2EqJvmeJ/kjNBZvZbCGx/G0sAa/JnKYf3l2lZD
CSGZabbvXB068XASVZGVqzNpTs3iBC7YNYlZmWwbU3lrUDlNyGW8uLykFLPAzeX/W09GAepz9Cvm
wX6ROa3THdq8BGc4NdiT0sHBKnnL1/AEkXpC61ebXndGL90ijSSGA9tSoz83kULDenrM1yyaRI0K
JevWUeesnHpW3UPIAhLPifrj6Mt93xwWoMo6G843n15WTErY+95x163mcwgmr3zm4HbiISWRMntP
yIHTQHBC4TAu0CdzP0nKEJKnPbNTHzTGeOCkCOc8OP3rkTyr+7N2ozl0SODs0l/Covzam7UafJ6u
/PfKdPPRUriywD2fSmw5UMoVqg05yni518SxcscDqbKaoDc1BK8qgiybU7E3LSeqPY1W/s4Yzps6
t066MrBlwg18ROt85r5bQxi5Guqp25q56TDavIduhQKV2YKDRp9ydBweJRDGzE4Ezja/oTMVMx0+
3vG9wa0z+Nig7cpy0XKQA1XQtfgeJ16M1dKuSRWKBKGakSPqB8Ggh6WB+LphHq+9PKUxOYmzOBz0
dwDwYpZz0rQoFMtH1gmDQxkjWIYKmNibyTgnW+zmh/PmI3PztMdjmYdj6AcUi4RVO47pJts8M22Y
3IiMv9hLfpZzhs9VFCz5EkQc8QDt5c9wQhnpQLVYR2rOFsmAASZZ2boy6ZcENT2UkKKt2yLuL3r3
tsE/Z5IzRlKE//K8bTjBWto8L+bU/wj39Iel3LgdPLMDqBwuvUeF5bMQjY6W8QLERPVgaVGeQ4YI
HaH+ZrQ3hGbJp08Pobm1kK+IpVNhu6sBj3nRVNzARH6JHpKnOqR5PznH2ge9PRON4e8PqnWiEF1B
cFu+K8TVAwdftISAZm/zNbNUsFDkVk43G7hTBzVpy5gk3H2pq1oUiyv9UNzlpfnBdei8rHk8znWq
BSafaKwP8aXbgUbl16v+xZ/bRMxblxedzXtygMq2pCyVdXRfRkQCQjLhFrckQP/oRFA2ibNcY7C7
aTyWFu+B2R45g3eWrtKNo+FzznI9S75MLSILeBgtD83cQOJWa2lwBgF/2EC++PRlDZjC23dwhTFK
JqynVaRKlx41wh/of+Ghm2FewcO6OgU96kHt1JDMssLE7oEkORq3whlMXDH2VlR2SzhFrVvDX0Ov
57SRB6BeEWKfyIURUFwqcLcJmlWinUyV6UOV8U6by3rglS9iFx7rb+azi9jaatsU37xsKErgR3e/
Mz20pvspU+gsMiUxG3N27nWQ3ANNSE0p7A2L1Vc15GtjB48AQIZrzPvEyA/ExgHdgEXdsspeTJ7x
cL8LrgUqU9/Pffr3PNlb34+/0TIDiHLYJbuXBamePX86GKT2UlPGc4Ck3+Y+iv1iP8ka4NLnmytw
0jFKEquYYUssDhHYFCZEfY+vvrWvfjuHiqO/59uVm3WsK7bufuj3Kfs/651+F8OySK+LfZoYthsE
9AEApeRzDu2p41O4ZxL4/5AeNeNrys9NvWfjHTmGj1USfTjTI1JzEyrnhwuI61MNmGc6upa+1gHe
TcNWjox/REc4wjgNnby1ndtRprwh+hnv1DfumpANMflVYSbxE7EZMlkwaZ6O+fy3cFcC6RK5u0m+
hEv3RlMDJecH5D3yd/JxXHQ1QUJqUHN0+4MmEgCqNYAyWtmHQvNrp4OQnOMmIU/54RKFbqs70GFi
uMvk5OiHSb0Pkq/K1ELWNN5PUNM7hpkOmQqC4ZMlKgGuy9PQMVlF5+tSZHomzQ+keufexZhavYIA
iS2WmUUByYu96k6UGK+NVUSfcUF9CRrR5YLt5v9QOr3EdO1KKv+4Uc2xd/j+r/SFwAv8jQdf2JnI
gMBcC3+cWBLxx34BrwVhFz0H6ZUazna1sjWgZ8sVC+qPaWL4TinEvYbJhKc/cjZkbDGfPS/CVUYl
gBoiLvj9sdluuSScddYPyqL9w6wh35WGqUpJ+i7AIB8h4djyl3/BlrptN8Y4CMf/x927L/LIjEKu
gNiod9N8jBVH7H6P0+y2NRUn48ZWnLx1WIn+6b7ZhUlko4UAz3AzYBHW9UjdqiEZ0MFN35fEyNIg
NB0b7EFjDYwJmftsUDHbB/gsHuvklSWaoZSlmL7xM3bD3Wnr5mjxWCvALQ9iKeNGh4V5GZwAgxrS
tod1uF63Xjr07DvXrE5vEZnu/mmnlsI1SUzcJFNlu1Gs7gy2ibSKPehSjEK84Gd5ILCYjFH6D8ya
EZ7rQmqfQeVL6gS2HQzoWbbTAaiTXAz234razxU/C9sGMtsnm2du+v5JgxI+7VvYizUo2DA+M2pe
OWNdIEX1vFPqcJ7osAcAVk56gBCFvN3v2WWLwDEuhjiBuBfgtnFJ3Turtv/5YLUxcuR8yfrrnDl+
xOtZEM4KwjCy8AEeQ8NJnJi4SINw1dN9uFesRI6cue04z1QDGRwnSZv1ebQIvpIqUm3hcAT2yG4k
QzK2FOIxOhj1G5UJRUP+NIqM8x/r7KjnBoT0+RmWyU+PkVIOmbtv9QJNj3+ih8ZMHOo4BC62HJiK
o9f/94EZbP+5pG1Z/+hoz4BMxKGggowFbUwqdjHDPty8iBatZtrcKs1rISzPVECvWn+fKbzF6C5y
I/89DMSKRFM5SP9KJrmzeioRfcm37PsWG5RZNltBP8q6XFaE0GgzpGRqrwzPYvfhugtcqKSGQVgO
HqxCo9bfQx+2eRCTj0/9bE8BRXjYSb+twCDc6H1jygZ+EbocSGo57A1RKNKhPld9YoXW8KW3plVr
Xzh/YR8NyX1mUS2TUjOlugjB11d1rwUE78qvDX1Toq08dLbV790o4GV0WQ6hY8JseFP3YElh27iU
22xFpy0uN8/cH8BIGM2uuHI6BfWMHkXhNDkD4yFxqsMPIV87T5Ey7VlNbVqMlFpokzECxzMKWiDl
jbU/dnAvb2dIKQ09hNrT73dqjzVuQEvUJROJEykRsnR416ecxy0CZbLAhznxhiLLcY7q1qWQYpVy
gE9WDWDJRwU7r5VZcCaSfRPsZcIiQW2FZl3+SLhu5GWI9BxYfCnh75KbLF39plvi+mLhMgKiA33X
zh/oMIwlPirn1VyGNjiOrhrrBIXEZNvA2fxZ+lKi+3zwEF9J+6beigMMfmJp+s2J3/gC4lrgfbEC
jMXEp+bngbwIbiehwoU55UXqY/chAAe4SybkZZkgbEg5IpYqtlybI+5zOoUU7wo7qwBvVjNkEVyM
qUywA+fXZ9wtUcJZgec8v3KgdgbbO6UpNHcfY3fT8UUATRhwfSkq6cyJNTSbxeulyy4QQwtgldmk
/92XdOEFMwKkFdlY9XY6sSifG5wiZqOYvAkyCbwWhTnw0pAsxSJg1RZqQZ+tqZRftDvWcMCewtjn
B0CBjNLfB7grgepZwZ9h9RTgJpfA9/xSDqy6oofcRQ+ixGqfX18WK2nOIqoD3hXWRM1bJSGsxJcE
FqLATFH8PNWg8WLjhOJGrokyMEQnvBie5xzj/4DHCb67X/W+ggiynDGPNxBBn1aHg2t0p455Dezi
kasctZ3kT2QJB5HRxXugzaoL87pKdzn7HZcRunsiXTfODQ8ePu5cKNq6RXmxhRT5NzRvURP8rU3l
o8mTDhdtuDCA9xZ7+7k0vHfxUBnl/Vhe5h6NqRMXKdBOtpKkc8YZUchw7is/jQ39m5Xb/PC7EZTx
KXc594vkv7eDVAtRbiXKbMWOjZI+bWRPmEMjtKgL3FYi69OVRLqh189GPqZcfjE5dNaq1b13cygY
aoUiCY5fo8cxTQdni+wQTIqjDMxFFiPdNPGC3rOGqTFmNb6lO7Shzj+3+2qtL+XS6aB1gFzOFS+I
LVZt172WkhO1sIIA76q3duls782u0eAx2Tpib9hpE8GpEp6Fjzkgx5+osj/g0ux+XFYev2RHqT9Q
iGg5pE70TM+bq41m/YShHp4C4laWODzLy9O7XJqUau5YYu02mEpefJ4K12heACkc7/1eogaZ2V2j
zeRv0e9znhmIbVcEokoWeI3w5YJDfCt43b7CLQs1ENsorQ2WPNixcQKh45TSDVdM0h85kabkKO+l
J/lt7fFvlJokN8T9Ix3Bn9f55WYZOwq8EdzVQe4UlqH2ehUFIFqY74zWDwV1tSRloQKvZ8WpfGky
8BOshbUdI34G6iyNOlSL86fhg402r1N271dGMqX+JdMCmq3o6It4nxlp5LotBFIpw9GF6B6KtO36
Yrd/C0Z9fb3RpDBLu98qG9or0p9s560sICXmPS6k1TlzjCiXyMwA33tlpLOGu0GsSwne1zZK6ip2
zPpqV6EW5aZHmdcEsxdqiHVaFOMHk+oVjoXIsujGryldoXFrBKWorIcS4QxDWTeiFmCQnRqliIy7
Hymdc9SMLogj8vpsYCnz9XIPB8CwWGYHrea2NcYmSsWzALfdX0yofU9UbVnIAOUTLrX16GM5N3WD
R/LNHgCcngwGN/DtP8i5NyfnD4sz95fdLPqIeXnzSWi6mABHmP0aICyalbJ9xc2zch8l6eBO5OlY
58NkTAACjZc9jHnEjXj7cMsQqn9SmHwn0toZPwRx8mnN2Dy2wgTw/HYLt/ggODFKb5aZqGXsHoQO
wDHOdHgFhKoK4/4K2Pw90E85k8usfOSqkWa+KOdqDX9yr4zODw3QJ3slXrRmnnY8B3DoX1dtVw9D
8KiDuEay3pyUXe3x8wW8qPrKh1a2fdFPULCWs+GV79DMOYliCCYD1f5h2+ux6yL7Cd1Db4YH8vJv
M4jIfCfy3bqZO6Hz9ZK87C2mBcDdcN5RxmbeokaBTXEO2gpGnly/q93PDfpn08oI9cImtTi29LxV
khI0APbSf7MV5mCFjmSze1OjCqzOgkfjLqVzCcaBTatZMUMUcGkXopiusN7uBG3ec7n8bpxNTm3/
SCrQeT7+W7vezKCflNkLnFeV8YWqGN4pakeQpjd7b3xDzlDA1ftg1AYMhD2FqSTIaRfb5yCS6buD
T6ZZsbJnjekeehOoHPdi2C1Oh3zNIknssUXmXCmu51WSCy0a7tZDiGT+RrQwlzztyCGARaxQDMG7
h3g23MS/jwjKlyvHbaOyt7UPCRqwPA+Y3xfzc6cC4dhzVzgIFAALzmC3nvz+lxEW4RakMIz8dM21
1x3moECm5hVkdQg6cMNk6SgizFsa29dRuaxM6VxrsxLacOhh0h0tJHm9KuBUBvjxYDxHKfpA0EFl
vEw9n/8yOsVoj9ycX6Aekb2GLaqqV2hjdntxwIHudRshWHyDK2/MMqubptOTwIlqmkvfv0rIL9+B
NRuqPWzVjrBFC3UVbbQSrKChYk3T/O9IilTGrf0SFRKD8h3ddm6AjQ0aNEHTutXlf4X4v/oZuAQw
XfwHJabpajC4ft8MumFb3ilidfxNQEYMP0u384+5exspB2EPvqzRAjlDvr3o4Gs3AkgTXgbW5ASn
4NzMD6VOPCQ7bWrkji3tQ0B8vwM3azHuCHoHoU8dUU3tqGGJH63vw+4sXgZx55ipJSaerlp6MJ69
B1PEWev4f76TkHcKy8hSgQ3lXDsvlNjXIeV6X9p1kicdFAd74CEjCBVnBK0xGK1M4tsswGrshpJF
i6XS0fb/czLwYIFG1GDhU6Y5RQVH3Je1LMZbTPbN3KIflSoBmkE2H/nD3Rbf4gUC6GEE7eiiCPQy
G8E8dHIuVfk5Bx+3NcjvWZ1bUb+naG1SMs2ix3RrgtUvBe4dwuUcOWAvbpLDV0qgSMp1GJZbOQNA
z2WA6bGA4O/wmKsL+zxJW2nUUMTcvpobRposnc6BZE7BeF6MnKRoHz7Ktz5s3ofgEroFZlWokSI2
t5dHG2zXtCWpk/RAKv3X/5Skef10I+9dfyMeWWoS7N2p4PBeRYVLtYoP937VjWRzNDwinPfWnty9
68SlMndHx98PKIlDM36jP2kCZIpcWCvgsBEJY162T8zaUGyLoYULU+cWxendAkH1BHx5fVqqDs2X
ebO3KYhe/y9Ok/y8LUntGaEZqvBi1+o2sievB1YRomw2EeRfL/96LvQ8yJrR8RLH7x4AHJMtDSma
VlBPOjUOlE3tlESAzStjfCbF6q9JjQCLWuIui8EzJ5tcL7EJXwgadqvdrtjulWD+IxaSnadYCEmW
ALj6mEMa0460orv6Bbfoo7SP90FVq99jTgm3MWS4X6wXEC4B+bkvdlfkiOZOiteU+Jy/PqQnLgAo
eB4d7j6hZbxVTkODg4xlDDzlr0fPAAEkjYby0A+ExEtID1UUeknD6UzpClnYO4l0l/HqVD3MRpJV
X1M4ADEMR0hXneMEhvwmrQvsyATsA4CPIXGk/II1zLOplikpi5BUHq+k5suqSEzOHkvJ3cYZyxTE
/90TW4gSoDEDydptaXyIrFDOq4okiueGCnFZawfs7O5NnBF9R4oqLMjkF7jcOJrSENU0wiW79KyR
XOOWNxsnBDnpzm61hP7ct6xWO6yabl0/Vlxc9Zfzs70SJE8En6fxoXLkN3awI28rpxGBCuSWFizN
qew7+G/gZabTBl/BxbAQTtypGXXsgoUJpME5HSGQRqjo3Juc/pRV/RKXT8Ik61eSBQxPN7K1rlo7
e2rc9yd6J4qfsWS5K27twVuvTSRuMRokdMQgTIhfp2zIePjx5dHhuK9kNlsLV0fK7S3fRcLdg9Cv
XjJUC3eK3J61hvIPWVaRooZYe6A6N053fYnBoZX3S8cU51GssyQ+sLY7YVSdMO4pwk8h3z5OtDya
b/RPwpGn4a1UIZs3umbg+4WlzTCAA9MtChwNL4ddz6Wbji3SMJOGisHpnb5iWz1/vz0FZUIAcw2m
DIOYpwRRk57rrooQ+yUtq8UQ2rpFZfhfrWiJXqdb/Axm0Tn1Q/4vZOEYqBLkPkKSBB8x7s7wJCvX
V243PqpH0A0LU/LmlB8mSTbi1U2Wp+7s3BLp6xVLnY39oZtGxvtrNmEBVRDsvr4pxmRIacrdyuDp
u37pMh2gp2xrQy8vjI+GPQn7U9844gx38FmkOQ8+gjwpVDwYn11jk2b8dqj8KlYXtiAc4a6vjChX
7t1HiOSWhN1mqW2rnHW7MexH3xqOrRbg9m3PZ93+OQguQKoQtlervhYxnfA6uOLNju+mStoFvqcl
IDWEdV7lQu9c2mVlCZjNz5DLJI5KgTI4Anq7OrVl1SUTD9wU4PMHUW+2iX9/5mCLQetOZjWNI3dE
AaSeqBDoz49n15vDo9xMk1ANkaA5w7hJFgdRTeCt+nReYq0tJN5WCkiVCcugFGb1SCepEmgB8kaq
rfwVVhPdKnRckDYBWL7iY0L3h+X9lGBPq3wCGIDjUqlP0ySYmYZIrsppc9gCoeIidxQe+QPstDtg
+SQETRpS1NWAx9xHFBgNeoMm5YW5t14MBE8g6uwf/3FB3aSoXuHxRMhJAj/yVW3+j8JrjzkUZ2rB
4qY5NhYwf8fZuYQlkJ4dRdTLU7EIb7ldhWIArFH2YfwaSgRQqeKIEy3DwhMKEWNHRGJScWoIimpk
hlOvT4YRJK7qOjW5RvFKA7NOdCe+pw/WWKxr6sO1c6VdcvPe4SYluZhwrrzEHAujSP+cvXa51cbo
rKXB0oGvUZ/0vjA+YOOxyf3/TeyiyjGhy6q/TVwJ/aL7OXgLMDM9jOpn6ARSlaILP3hp8YDHfl0V
58x9a4bL3c5IymR3yS2VbxJd/nyuimkuDlm60laVQNUYJGzkvIRZA16T7RFx6NQIUNE+HIbFoDdy
99ujozGn2jqC4lbAkVluwMulebRKiNuaMabH+nNDO3bUicRDrtrUDDI7Lr3S5e8ymm51pukVFBc3
Fjn/i0SXBRo57IWKjPYzmsesxSPBoH7xd5iFCW7U75y8fbh9j0Oqs2oWIKPMg6BEdhKypHDew7Cn
La1Zk1D9WiSl4tEHBY2o3mj0NCtQgbeKlYiMLEPCkB2Ar/NzQ+4IKcRGC254CAWvjoubX/zt7w45
kfXKOEoxoWLm7QhXmzHtruNSTKS0U9sM5GGpS9YXRS/sxr4pvJbHQ8VkOU8wF5FX1bCwDyRPE7L2
xXJVlvBuWJ3hdpxgWFvVKdLSfOX7sQHExNMEpoDfeescOn4sdZ7zxzwrobD0AU+s9K2HFNKzEJlz
bpVkv7OuLG1g56qpWj2a+1ODFcttFD7Z5Ybsvvty9vnUN3hG6l9OMgWIJdg6/daJrPMijzSowDC6
X/o/drGJaWW1+BfV5bhLqGpVgseWuMnEEsKb3hrbMJ2dNyE+F9T5JILy+VnT9QYbGA5ZRVpHbzsN
NxyRNvfNoGgE76XfpvmPLMWlzJrHz6d/BLAW9HfZVyT0WM68BEp5ztQy+tZHc3Z8Ql2D2SzDntsm
g6LBZJBig742aaco6bGfeeOGDjrGXo4NwSFcaTUXix3JX49OopCpBBXTI5TM4hz19gCpaxWMG5dd
mrOXSE3wzS5hoBx9fhKXNv5/igtqwj03dl3TiqpeNjaZqxjWj7FQBNjvBQb4kVIa+oHnvwLxLeAA
Ar7iWjCMC77heGbUDfl30FfegtOzO+2gcxutC+nB3JlirFOSAgYRwLOwbe6vUfCeqeLUcuUv2kCS
onlujNztDdReukmOS1pAaW81crw1gSGGc7iSPUk6b2zeiO1gJGPgnq/ODaGLKPK2ukuMMyhGJmwP
T7KnHQaMa6pH0xYzMVIcFj1mC2BRZRNCt/oOJzJ9At+/mp/uL6D4+LEVy155MrXytbJbsCwOfNAR
2HnRfDov11YpgWiJnW7lNscDq5tKaajf5Zh6LwjZHHpb60Zp5CmrhHqkjdy/prHzNMSpYeADHr9M
Kji9vBuCxZ/nTtUeqCDovbRnbHlW9MozeOjYUvQrz+7H7ic5XPhB8Ikjq045wAGxibuM0A8dEiTb
A59FO8fc6fEv2hye+A9Tzcs7H34Dz2MjS7Zqqsy4AxxTWbMDvNVfUslDI7xA0dQhw22uqQ+SuAE8
T3dNVsjP5NJH6Vlxce3irF6yWBuHogOhINiinnFK9bmlwTXRIsCRA5+UqSlavhM6ANr5abD4gEiy
Q9wVfn+vJoXAJZC4s/lBwCFNjkI/I127NHz9GlRUjc4qRyw2ieklImqO0+VVCJnKwjmQB7AdRQg8
aG7t7ATrR4nB9QdUTpv8lDUUkvOinxt2dQelwfzEYwCRgF5a46YRrhFU0u5JPMclfZWTPp27qRQi
7iW29sFb4Rk8hvzx/upLgLAx5hoHJ+UzF7RRppLBBamkAVkrHvs8cTDPnk+zc+ixRAKuohXp1UVb
BYJ3/tnxC2otdVZq7TeDgze/nvKNEirOeADWkU1ZvvqdZ6vJqLZBfXKcjKbo6zAG6+7mCbA4MUDm
HumRBxp1VCzPilskENPffzf7riUMQN5re7wQd7IaGG3SKIUUoIm6iaugj7p5LXI30SnFZC0fpMTn
IOGcUbtzKd/QJv7PgmS8OvNX5UKXF7u9r1FNNsbbHk4mXQ1sNLnFT5X4HszUrFxKT1V5a8uHdS2l
WybDUKCILhq6NL5UgPK8/w2ORToRaF7k20HV/AJM4p1Azb7fnUKVy5cIqZqsMPRT6fWb43cs3E5a
fqIoXVs71JfTQa1WvS4bU80MjJ6DTDLNY7bua8ioIfrfta6hpU6L0MC7HHTmJJYsvg/1R7rdXzQX
xbI8z5lIoDM7eWq+3We17jyiVMlKhHW1nJkNuA1xYBu+ri+QFgw6qo2SuhQZL7cMPZkhm2pdss7z
69JyfxEMJaKngOk4blTTprJ8ElSNYSVCM7UZ4Tr2uy87JDjeYFLHwE8nnSdcebcW2ZOV72rxXnBA
kfxeljO3cyAumylIHb9F5JEIS5xqZdsijuqrcGLig+rCdIfJYtef1hyjmIqeDR9e3G6pqrQudEuC
0vdw2a90/kpkIjnADatHUlo6kul+fflB30No6agn0hxgff8wcgfI38GDctHO6PeN7mHaTltmw8bC
A+oe+6VV36aeQaD0JXs5Su4LuTNubiqSFazkGbhpiA+tAihP9Aok+DD78zELl6AnLF6xRMtcbQ5Q
B/du1YqWwjG4nRdzdpUa6PuXijqh3V8r/Fw4ALeTy1sJZcOKwINK+NUFuEWjTOEXI4BiyqOZpTKN
Q53S7lInVECFu57F2+j5nSbaqy8BF3lnizmOODJxe/4pTLacnDB1E/M8rZqbheIdpVqzi0LikkKp
olwg0F8taGpKEhFjZe98UdHNAPabe52mgB+OnhVtClDoI7a+ytTIPLgHNZ1P81XPLVwJG6puyHPF
Itn/THXVn43Mp29bFf/2CeP35QJqUS7cwR7Vpl4gOMlFsr6y3j4HdFZ8EclbvWPECiJPorigRcZW
SL7exreDd2Y4BT6WyOGcjPSDL8jB/ZihQSWc7KoTExhaHfOEnpaveQ6QN9mHzTvX+rwZ+MAZucCP
UTpJuBOjG8ekzR8vGL4gi/8hyfHA/Haj2dRKGfJzWNSQ30Va+MleaFxLWy9jWlktbc+YJzDkWzAd
GDV2Bgi251uzg+zuzMI8ue5m5/eCLo+zwMxvyoAnfsZKeZHsIFdbokyGY/owGTWNdzUquzwH+wLZ
8AnP+60YKDvvxZOAnMsPuTjFyXLvRRqPtFw70i6H+yrfe4BJfgO7huJyclqSZCpnLmW5BbHSKOYd
S45DL9pTkDs1KOsrxy+B2jcT9HuLiI2n7MYlzNIkbvjGjVj9T9T6Ijfvgt4OhbTgDyl0n98kXltx
cVLyk5WX4ltHo05uolFgFW9Bcl0OoCi7oGqTjqZKOUjfzYdrpKh5DFbMsi38soguutEio31Vv+kW
8MpMeYLYHnRoikT90tkJqXEEBjZz+Q9hwNWfRfBNnAAzwEZf90/mGxZSXezbadCjC00nvoMzg0hs
Q25szL8YlmIjZYyNJWNzMy9qe9RJwyBb1iG8mtV0dO3CIh0wPPgn+K4WZnR4gNDf3CKBqnwcW1Qh
3Qkuj7JdJN/5P60vruo0x38vqLmYcVrVIXscniP3PUb71BDlV46lv2QBzVwsteRfYDh7u42xm6ts
+86T34nhjzyrEY1xdTfQu0mnl+HkcrvUiC1IFnlaG6yGUw1TaEqNkp/JDzavMgGd7lAZpBNTaje7
386Vbrq1LZ+V/9lpfwh2Fp+V5skVJLqIhu+cZOhtRKY0VTOgIxrWDURfRzFrX9q37fUJnSDSzXvV
WkGzvX6O5Yi6r6KBvtxet3oz94s1dJMLkMoMAAM67y6SfYEQRavutCPzEvWZ4I4ELEpWwdAE7QG4
Pu8Bbp77lOa21EW9ODhBdZgJFAtyoECUQb2nZ9shQIJ1W8vPfGNFvDPV/WIu8wS2DUBNehwFGL04
fRPAiFm7v8fdurx87J67Z0CjW31jUj3+kr2VonX9Ntw5BXjJawhlbNLTKft6lPL6HqWZNSECl0Cp
/Z4S0ujxrKGddXIawIwMg7utAADuP1VECe62FfLg9OI1Aw4D8J50ORQNwhNlnDcAVdfKsz2ZGsuG
w5/zGd1//eaiXIriEUvcU6p3N/6XXK4IPHcg1afHLbzBLHJNc8AHw/EAWmuC32OKqBhYRXdyjMh7
3QOdGGAvsjJR+WiWbQRjaThLSxGOy2fGHX8AjR3XlBemiXy0X9e+sjjtxu4or4bheyp81mSKXH1U
Z57TXhfSglTIlpD9n1x/I8NjX+GyiBM97kW2zyfz62GsZTHdeZd2LVUkb5qzsLGNYL0TPC/1o7QX
p4RFUHPkvxK/5qTH/0GY/IYIlwwtfDpk/7H5kxmbZNGv4fD0PWwX+MkvQkiBi4tCL7LxsQKA2GNi
cQJMNL2x0C3l85YjBBSBukO1p9iDuXDjkcsyJeW9AByA5ZxUBLCq+QgXwzF9kQag+QKMtuBbIera
HSoo9JymegooHh7+0VpKCnjLaudwqVT3NQsR9rRmAriAGao0DtQxNXalX7AjQT8VEi3qndnmcZMi
m+CuNUDf4THrcoUnlK+GnGwahxaMhmjmcMS6ucVR51yOfgFtkfBKrgmWisoma287orbybIp+FjhB
qOvb0oZ+clK6UnVNTH/o9KKcCztYJE5Ny0XBQPj6A/tmSuKg1ERO5/W0+MVDuYRAljzrFIBVv4ll
nyjptWPKVH9Zpn/MfwHhQQtS/cXB7F+k7Nxk9hyd6JoGSyns2BArHNss+xGhp0c4Mw6i9d0C43aQ
hRyKJxbrZE5cNpftbZi2FxVn3HW+V7lsahFp/xLMKcpU26JMp8RWPd7ekKeKvELLdReHdSGzkZg9
i3EPgfInDx4WW+q6/QiUK26BYqjd9/pOClN92v+BdB0rcU2NGDl4yVcg2iEk31MKJCanctwYJ6fx
utAL02tOoO6fbbOo1CbOZk3ht5y04h/E2wZx1ZRRTetc+WkNjPYfRf03B5jkM/N//MT8Iz9OwtC+
pE/4khPLDkBeruv6rze5EJ1Innuo5FZUXmuY0xDaRplHAFOJE0JFjRrpdopgQPaeTC7QDFDsDwwo
rNF0XRP3HZORpU1YABqomyTIW4MgWhlvug92cStuoTK5I4VxCnBajzxz8cNAZw9wUXZhu7I1YkqG
yW9rCVuh7/gZ5THxNgZyPqIGVkBs0Fvr0bjT9pDUVBHfhmhl0LwshqDPfj4AdpfWdCjLOma4nyWQ
SWXUwDmZm/bwGp6oE+J7iQdiyLsCwFsS8EhewKtbSn9t018QiO8vNcGzhqkmKNCZpo3AtLSkMt2P
tsK4g795prT3YlsHk8/fChB7ddYoeYo5Pj8/Ib0gcPMdmXiCBXPGintNt/EsnHwBd3bPJselu2X4
wlikek3HE112JOT/OqG20/7r2XVDz+lyhGbimNweATqW7TQUNbDAD0lYunW2G1c4/un2ljt/1xo1
3Z/FJstbrQFRGbOfiAwgFPipj+zMCZpNH9f7iTZordBquvBKsKaWLyfx5u1e0VMAHeTPARwah33K
4xvooQrN0DovOruGfqYoI0+3EPK0ipEOK4kzfyLb0cSNIRsY4YBtxWCygqnAaaaGoiu4njqTs9AK
bGXRNOTMMnEcUVlJixHKMdung1gI2+8uxBlqllT+t2F5bIoQASq8bDkc4KQSISIZsFt2e+OLvDqE
nmDKLbTABBT+nN1SK2k4kjKi7TAiLZy8dTtaEbRzA0multxqZUtU+CXQvUddNuwjeXDOdDM2h2d6
K7u/rIn1n0eUFGK5d1t7c2AXouWi62jo4xpXyPTNRQwNkNFprSSVSpRMqgIgrFpZ+ht9Z80Gwr14
i/Le6BKzz3C6ZVSmT+Xo2SZDToIzRPyet6O2rmTUviqu9ki8ir0iI5fFB8reJ0BaZgEoGxOGBxOn
jIIDaSTR1auh7KpgNJiSJLVFmW8Yb7uHWV7PBUUal/686VJUC/XpnSrs1LP9C0KY5mCvoaLqVCoV
PFBqI1ZksFdixLrDDZtLJywbyHbELKT6RWYSMSCq00QU/EtzHlGMwy3hB3nlo1kZ+k2p2oKMhyGV
T/gnFoh1ayf6W5kNqzwxau09diVZ+FKxXSvQMrIWW3ix1guVEx8in706GcuzaC5a2CtWg16f0a+B
cFXnRt2ANw5QADy7iF6X2FgNlYUWnntiFlekkePin0/QaGDEUi+M6JGPGQFWl7dJsArveJv0G6t9
dry10Na3lNuKyDibLGxL145Rq16WwO4PB6LAlSJZEqvMUv1tDTeQCarw8hpwhgvU/P9q8Ozc48mD
O3ED0+evTFVKfEzA083O8XmvWeJmSR7WCALKrv79oH7Bg3H+tOP+XOo9PlPu8BmiExxyZPk5a5LQ
HAYXirwe3MapHAs0jysYwi/dRjWRCb2dDDpUzL4A4oXnT32QCWGlopBGRd81Rg7ykgQMsu/bDA2s
YQ2AwzSf8CGm/mUsuUGD+ZxpP/weKbbBtJkFdufd3LRqAtbb1Z0KbLQQuPp+zXHEYvIbOosZFQfq
+jKh7e6342Vi55ucO/AMxzcVo5rn7TVoG3lNME97oaZzsJJ/o0W9/BLdkAtKNnSBHVtmfX88N595
s3ThPYqxMNRoywL4qgz9UlXMjrjmSnx6ZvSUuwRW9Lia3Ukh2bypywkTrxkYcHrnI2GBiFgn71qj
aVcNANCKVn3dM1328txpmKq9LUsJMeotSXNKX/iiu5zgOJNf8vQ+7y14yqT9sce0GgqL7LDcoHQn
pE7MAxezIsWwsNNjUCdwqhJZCtKV05U0AOUhUXez6dwyAqbvjE8jwav1bD9D5SEKkJTjdau04j0n
NiERuSn361yA/rVQnyJr9Pj/o9xyqO31tJ5Vq6myMnseQaZbo/D8t+3ARSHJ0NgnA1jRa5Je6Fkw
rH6jH4JiKhBSSdqx043JHjT8d/QOMklTnndh+iIpp1/ypj+4fPQwNY1FDSvlCgKos06FqavjFfOY
+lgMbogn4Ua8N1uc6dYN51kbnOGkZ6cmUNQldnGrt4SLYiwnjAqIuwrWLy7pAIs5pT5fRJ7QxANx
sgdjB/w9qVdz7m6Z3DMc/CReNlXrBWlB8QFRhtJqjpYdIlyPHOwTUeb36XaLc5ipHv2OKlkOfPQf
VNt7wNhIBY7PwvDQSj42n4q3WeP5RIn8CCDMuDeMrJHIKKsf4hC4dTotPc+ra2B+yQFd9KSn4BEv
IVJj8vUX/xG74KrSGpKVvBs4mEC/RvhcgAFzgWwjW1SRv5E6XixILSBx7tUtZe9SYZlA9Pd6GF5K
m48hU+4wIPzuR71DF0jd2qydGJcFBmSV+7nT2f427g2GbSU7lwpfkZqEr/y+vq+vPO3g3hNttPm/
R5vzmFvIeu9A/DHaSBSuAMXGct8FzLJzg15UtfhCKgPwJhm3rY4ge2kb7ztwTe3WJZ+8RS3t+jHA
ojDq3KEPFZLM169sOe7O1TYEMcMchSAe9ZclmTLJi1JoJBolE2JXgaMKHgXYr365cR769JsB0gVu
yz1SF8+j+JkKOGeebBMiILYdF6y5WI9MPLCZPdPDSLLaZzw72Ha4CasNIALHUOvNGiwT5xCSXSNg
RV+QnTx+98sXM2oKkR5aUq3aQJtJdL5+9/HyG8NpMd80msOQzZHPMVkFtgyG9WYhkFKrZDgFAzCi
tUL46HD7rNlxep/rlu6AaFgICC721klh2HZtDALhqFIgenPGUL92zBTzISJI2xMEgbPs5CwMpBnX
SfuWFoN38OUzZUPzSs5aUHYlf0gawspy0pnLjgv1Xc9s5sfsl/UanKpzDu9jmnXrC44wJflawkuh
SCP8z4GYZlJW41gBVq0lD+ZeHkc0BJj5NSWRFVwEzX5XKCTN2SFUVt+z6MtJt4bIwu/6BY3zJWdV
9MJhxn7RZdtJbKNP1FGlUpDTucs+JHFufx+865PEpZ+LDNOmsrIDdfm1dq9vk2IUZVNsKyTYw9FX
18TXLUQ6hXmkFYunqpygkiAj4/1NDqiETLxRvFI3iqfb4IE5StDkSJQ0sQjYrF5W/qv2YkDrRQHo
eiFDaqWnWcVBKBke1w68cJ+VPmdOm7NcNL+OLm23vT2h3cRd0H95ud43RFQPLGFrsUsJ7oKwwrEk
zGQX6QEP+U5UGua4RAR30s14GFX0AnLIiyhLl5tiFbZdc8FIadJykYbvOC4g6RF1enIXfikhmQC9
OlhPxUUzksRUS0XfMUg0SyQ8fMKNOHGVSU3xTHS/KAIRsdtKeEB/aQEpK1bs7n4mj0I6ExwUXJHP
nEb4srw8Pb2hcsGoRNFgKv9YOgeXNmAR0arJAYlW7U7zDketgMeI312YbgPVzrHjTeTQykY6EmyQ
C4Y8KkqAWC1jY4prkxLxHFCe+lYD1dRgw1XyfWwTbTHhy8DlBatfS2COXdCUsdbeWfPXpBmM9vYK
inRTtzgsKMFkyzB8XzkVVH5N138cXMqjnhdcEZzdFU3QPf6VCffpNFxT6wVgATMizTX5vKvlrfrn
EgN2lFVqQqdfZk29gh1vM8UzWoPy9dygtsGT3hS2AVnxBn0GS3njmig3hIo+byO5L0InyhKFJlab
Doig4BG6CqTqons4ufrnqEs2CxA8TnCVKDZ0ptm9X41PSq9pYxEEEZ5L/bMVhSw40NalwiFqgrvw
o8qucoURc4MfZNwGQpyXCGONqtUqAFSWNWVkkAs3yBqcX54MEfsHqMkcVcn+hBhS+DiLtVMcbph5
uYYRwYLH6zS0cuEmC6idnFTfnE85et89Ls9DF7AEXqrYMoPdvaKFoCGUgzUD1qBbRoh1HAOgLJbS
UNfKO3v8fnh9S7ODS4AdoD/fr0eI2rAMOt/224kQ5gTSGCafPLc3FjrsyOe8EHe+QeApFF92mAzt
mCoj8KG2bznRZQwS2x+y/lsSWhr0oUJFw8/UkOfKxyiEFndJB2oWqAchginFf/i+qCNlIbgei/6C
tWKrusmdYF7xSEI4MEUjdZcKxPmQr61FQPLZBMqIcd7Lj14h/kkChRviXtXuCh8ltUAcPbhJvcHN
AROwHID/Rk+eKY05oqpKh+hLqr0aqStraTfHucZi0p/kCldUpOuO2ZrqpYYfoZy+VlY6KT+DITTP
eyPZm+jJSGDHRsdCiZTBo0MGBKj0+nnA9YzbHyTZzXibNhbAMPlnLFgKTgiYayTy47RxXAws6Wai
RobhFyag07/XW8OUk+fDU6VQLpjgfSxly5ENrBQNkvjvn3QvwdIjWx5YjEb2VCogVoROmLZMl72f
dbRmyDuRpvtxlSImLrfLIwqCFF1a0MJnG4VkZ2fRs75hDuO4z4+XA3H7nZeD2M1XKo7S/aHk58G9
xnBLMDToh1vy3YcvCRXPgrpUyV2/CYjaeQst9fw9WOKToJ6Hrk4jQogtgdjYubhuBc/pzWq8NG91
T+k7cdxzQNn3oU8VRUAzgL+REPVT88nvIYTyzOjx297GsAqgwlbmhyfge5KZ2WkX93sRyRNrsNCj
xqJvNH24+qsuViHwKCZAM//dFtq8R+eohUabTDHF4XuKJ1tMt9z8oHtwFa7rgUKdMNmpEEaU+7a6
wi5RLGyoSlcfvRKF/jaNFJaNuFzsrvumqr22xC6vL/DTxwGIG+fSflz3pqgzI2kYN3CZqseVYx4w
pgsXLHRbohWk6f1CzHtS2Qm1PBUTDp/9p5r4rN3tavrVQjBPMp3ItYeH1cc2VrEeMm+VByA6z5NI
ZhCzfnZ78I47zooIb+utWskAFm7DUF+KrtjLy7GeOhoOVAlJTaMo2cCOnNvWkNxPzk5UOx1zVclu
+SuHGYNcGmpp4/tARUVt8fRd+mEQl0BP+6snRSHHYm7skMRP5dTUdvc9plMLLQ03muZKzpvi7eyT
bhBjfzijao/ZoVdQZoJwBADBuo5n4i+yakGRD6CgO80QKG18qv9GtpMkFza3U9AYYJyBmX5Co2zn
by1K2Yl3TSs7+738gQeOrIfrT94Yk6SKTsa9bNJyeShAce6598OjpL66hfz+vh6cosWjRLrkJe8q
LX59RLsMbhleZm/v9hU7Hr8HbnZ5+JS5qOOqe3pxAzLx8caLFeM/TywNfq12kTpmgQIEdOKIN4T9
krbNycc8sSr1GPdC1d8whdcOXDlJ6U6FIg0SdDAFjBaDswBW2fh6dw7W4bS4puLoMW9ErdKQuIgV
BNBLodOOf6QeuFQInAZwcxnUqS3HZKW02ghH7GI1AaBXUScHwP10WSCP7kI7YdZdWmrs3z30eVWD
32K3cVYkJgpTsH0oYH5FLnOXc/LG/J13WeF7oXSjo5GuO6QCGG1rb/8hIl2+8DJgEqe/mgKnSgzQ
rwHdm+/9mgV2uyi8jv4mDp2JB9T3qq7OTmVfyCSSCCcLOPXsGSCqsPsFFTHVPSbpMJ54xiQjFyPf
zxXT7rMZondIJqmeXb+2NIqPgv+sqelnWyE/zYr7qBcyFtB/03HOIXp9jyIV5XaJ82J4MvUSbjrT
kuH0XAglcY1IOKg5TpJmTxBMjc+2+BAmbu9d0u5XnlYOV7Fcbfm6AY9KQ7L11HpqwkmTpStPasUN
WtnrJpIuDV5OvN0IZ928+dAqREAvdGlTgUZ6jVh6lS9QYMBmheyNGMfHf74/CVJ3cvkpjsEb+MrS
znOttqjJPw8GjVAvsa2DO9T45uao902J5an3Jg2SJXoZW/e1/3G9pvmuu5x4QVkXDYXrKkZkt05N
zEmOKKBidWE7ihvkgERddqVkUyBjdJnXdv/AJMuG2eKixK/m1jnZarJ58UXZJxltIImp4SE8C/Yu
mrOcZQPnAKL5Z5VWQXY2IlZEQ2P0Q+UbEFCtnbhTnDMrpHttYcQ+uq7oV4ZHah0kMCl0EBngDcDV
7oGOqoveVHer0NdbApKIPgdAi2zOAHBJmJY8VN0FXSIaBZ72bBEcvNkSznhD6Yxn+vi0HSvn1Jvg
jn1PekbS5GjS2eeTip37fZ+UF0JupSTpBZmlPHGzQQC37BMjginJDqmkxpGyd8SaFxrxUUZ2JcUh
GSg2f5EkkB3HaQxkv2XKtPDgGu/teKtPFPUjPXaLwxNpAAJEsmWvL3fH2K3LfUtErMU7Q95koZF9
qqOpVNQWcZgkk9U79O3SYjqv8eZ8m2Okt1qWFRCV+9VDgDfDEA/R3btRFwyrhCMZeuG5Z29vyLN1
fsCMKDBZCn90JehdnhST43kk2m512WPP8g4WAq6/G3vDVTMnMj2VnyXnItWfPtdUOUASdaTlRim8
q7a6R0P7ue0DmIAcFp78659d2ZKtUIjhw9ty7263kLji0z2Vp5aJr+hPDTVxzpoTbbVFsh0NSskB
40Rv8C6Pl3+OoD+MRLLMooK9rM0UJy9h5yEGMgmmLJojALdrSo+5FJroBjW2RUv3BwyhonuQ1dqK
sBEhI4oWPdKo3UU6++UamXJvjYStMqcgZhMKMEB8IwPHlMX6ZYKhFJ7Z3x/JozPonvyPWkfEa/Ik
FYAWL5YnxHEVUXX8zBG5NfI/baTWOLr9FdCq88yUI1h9WAN/zuA74y28keZZVv+KSFCvJzs5qSf7
+kqFyJWIBe5lFLSdgjPG4opqXT6W+43lilrGxGuWfNmvbneRKxPOoDt+4hGT3B9JJ7Yfp4x2Pp8L
17TsKY5BU7xnYdkpW+HZgX0H8tukLJ5tQISa93ngQ1Rx6TONfZcaOBgWESfVyLREQ7bvyF4gj6q8
i842jXfF36xSFspolvAsKLyJ13rZgGtVwRngpBPnoXZf9Jz8rvJ1tUn/Nxv9O4nRq+umuh9+zquF
nT6MFJvS2lwhF59gvHc/rH+PHjpNqXh0fFPKyFMXNSZMr5CgA2I1YiF5UjsYAgglUszm+Xcszy6I
fSfjCtRbD+BJTDnZSugWnQsCKp7Hcb8RYfKsrNOaQ6mMmD1kVJq67lOjoULjST5kTOAyfXvmKmcF
6/MTjyY/fVTkUDOdjQECYJvAt5Pk148GvOTCnm3tRQ/NNSakOoc8lalgI7BL3im3p1OujRwSZvNw
4e24j/vb70WwhEB783kBzQCgClUPSVPUR8iLP79gFArPvBfwR+Kovpj6xO+5KdAw1MOPJYXh7H6I
1uKLaCBnzTNI6Uk6YNp2hrYvDGTvJcxtuqHhOmfkfYwbmmKN4bTjKvVEgQwA85L/qp9pcNBQB7SV
HiWWyySXfjZOCxTIMuSXPtoRW7hp9n8DqAJQt7EmQ2nZmbZQlDLbbP9FGawl9FPtVBa24yBdMca1
Otn7Z15+dr4D+NU5ka8oryFJhV34OdgWXXCh/nw3LO1XYXbmcD6nt4yXggTqYYrMU8x9JcQKz02r
F+WDyxwciBJi5FZpKD876sJuYPd/XnE2ezRbwpQYrtwFR/HUwkuJ6kqWgLPEcdzQSCmlyuQ3V+Am
kaOdcF185vN1ZQokoRka08MX+8M0iB6T8XykR7030iHwtSr0oHc2IDEa0JhqXQh8GYgUcUGc7rNS
UuFkxmyFVB/KJHHwJ5+Z0mGkeJcfmvp2LOjebCPan/Qt+t9s19raaXfUxSCJPQojzlnIkgeRIDay
1swQOOUPlc3VEYodXruhnyBHDDUz+U/TSi3eikphKTCwYvnGFBqj41iJzXdKAMmNmoGUtbj7cbB7
vxRfqnkHX5UNblVkhp29yEECGyMVl0lMnrHsGaSG/k8nM17ptHctXx499w2RvkZl0qMzqwoxLhOf
Wtb4o3nVNmPYzS8rzjy9HQUQB3d5jWf/EOUoo/3V1z3YQR3zDcZ6mjMeUfEhuQYbMnEdy/knMiCo
9uBIIPTYMuRks9LGf06lx8X4h4kcZtT3KCdgMfeJ2CPRwyRyRO5JtoEOtr37ibZlml3vpbPkzv09
X1zUImBuzGpW1Y2lGeUTRHTfyo04mwnZrtl5bGrXuqBWpPNL1mHkx3gtsTTPfQWF9OGCJ0gq/PQC
2jQz/FwAWu8eJOK8vtziZqtz0C0AqB4CeP9YcsMSTdPrLHyVSzOylKrydfLHCecEkeilP9BQ8oPl
ejGnqIDdJM4rJD3zMyZrhet7pAypA2S/Qhkj1uZEfoojgnn2VDXRUHeDjsvTmCgoB0i7k4vhIE92
Li+jmi2ANr/FbJeXR/drQltgWWGHTQvUnok/EdTMO78mMv1lKmDv7tF6QWh5Ai2mpDhTHGrcGHjh
xqn2NUnruuB4CPtefH87sgEn8EPGIo3vWrQjK96WRW+GXF7YLoVBL5jkoxRqNypAIK7OL1clVD/3
kW7+3TYTT1hBeTWk8jpc1VtR74uP4WfKnyAZSdoNipRL52N4HBJ/F70E9izVC55seostZ2tpavxB
34TsnYiUQddpC7VfVOTAQf3wMDTlNT1Yc+5rWK5bvEBZL3QEwO94I4SFO+RYuuwvbkVhBNTpOlot
To0Pg/nfm5ZLFzgLuzpB9doNXN81Mnr+W4gD5vLyQJ4kIyr9IgQDJhU1jwWinhdqhnB3vHzQY6TQ
jUhRpdxN+vNRb46TR4FMW1u7riOdavbeiyUkwHa8O3h/EeZo/wL0tMCaTkUpra54vDzskJRXXYXV
3tvupuVsRICa0ctxnxWadU+9pyvTgdzG32ZIP7Am/xA/7xQUuKM6AnAgV38Ek+pltsi0Dwf3ewv3
eQzeaNFq8WrtCcVUmZw9myKmHPjBIKQYd/J73UIDfP3ul8rp+w96bV5JyBHBWvZUhjpnRNEgxiq8
LmS2WoBlIrFRzGhtHtX0mrdeKGqvzFTK4nF4wB1R9uMT1oozNLq2fhdfXPRkbuC4cLSLzTUib+YI
UIwlmM/JzojJcLG9pCt6gXlYjMY9jEs22OyXA5D3K4DBntY3R0z8ZSc8l2ZBCxQNRRP5TTFa6cos
yq3isUWC8h4WsBb2n571Q4o8/sW/BjWX/r0pFiERpaCJym/p0NKq1QuMHY3wPPe5i54y8T7E4/kl
W0htBBruAiEIdP22//a0J66+Kn9/+u+q1/iyqnP54/RtDM38M4y51wiadIqhZtu5Osui7XbhYyiT
y6IH9qSe5zKVkaOtHF6eP50S0wKxCJhXndz4Igtey7B8LwyfAsJuhsQU1txX4dVEhO0hlri8f65H
isAsSE6Axg7iCeRAN6g5nV9Pb/fYm17VwxWTI9QD3zMVJ8vorYdQowqgA39boVDCzwzvO6qPx14a
7dowveJmnqR1yuj9YbFX5GNPKI8YikYODogEeQEMmm5Xkf/2MSA3Nuzs8qkrcMa7PToywwFXNAdV
MTcQQbae1ZEB79N//DgYHwqZdRfosw8UEL6D3iHkml3paW8BNBTDYDTalgS14AYZXBEjbcTkzPXf
N44o8Swwmg8tcElCtyke+ffexfgEWHjhfljzVQz3aOogMr/foLcIzWLqWiqT0EsCzuOj4vJuJqIg
qZL8p/RxtimBbpGcOIQI1p7tHmLC9odT8zoFNntuufdD2LQmUBpdHzbwR9jNyb2/fjte9mXoOxzz
XnHg7pGahsrgyAqdqKkMkgDkhuZDg/cYED3oefDPmdIAsUc8TuI/E1GrZJET3hzbqwpkJ3gxStFc
Z3Sm44gOS4rB+qlsF2bpa051jUYdbI1Q39FYiEVubpoTtTvHwSEAP9WPLp5G8gLbuDqwubR0F5rP
Hhuot8ZBQpLbrWjPl5sP8I0iofInUjx/b+Yr4vimauY392AajzeK3d5De6rpgnW4dxjZWRH8YpPI
YE9QY+yeQ0m83fawhgaILXsyigGGjNDVLBNmrqL3Z5yLO3pwBZAJ1gxvCW5xT0qqhhxaw61BpaNl
6IUR/f+Iv3w/muqdxYDkl9gabfuKW4uoQICkGKyIby5L9AJRjesjIM91SyncqPWB8EClTja/NLym
G3xUq+OoVsB2jea/Smptm0RFTtonWr2TfOmofWcCkon2RHGHHQKpl0DY0S6Gxlq6E4UZPmrVFKBe
U+hl28bJpeH9UZEUWc2aFz59GR+JUjCnrKlCAvDxbqEDKYcj4yX1jesMU6canM3joKarvwwIftww
0jsX2tLcykvebquST9CwjraA51vxsfCItKB6Y8u2dN5Qt2XrrUXbHn6BDBD+6fS5xBhfiqjfGGu8
biBdOTqT3NQZhXo/1vzmmvit60QDfuGx2vtlum5nJ3F2YAfZtGoymd2//uabJOIknS3ULwRqQeYU
muZI5CYdm9b2Eg94yC2XBQY4W1H99FYP2cz5QBHzhP+6fxsvxYJF6YAllgZlDxUxdRkE0i/nG1ZV
5thTs8lkyeojol+LY4ODcE52uiFSlsUxUfEf7WPxmhcTTefWCXDeJC3B+8yaJ+I7kWRcQbXU4mQ8
Pb3Llpm9h2ET401ii3ZsHh4VV84SxqbQESHGlc3RhxatWgSatmUfFxzB1StLRfq+yyEkyrazSLiw
XLD6OqiAcnpxjH0Cr44mwKVL1I/rQhMa74L1kdufE6vVfv+PZYua9GqwbLpFlODZ8XO3Fwx5eLJl
8gXCR9wSfDz0mfXp1YZX331rY+Buw3hVeV9/TWylBJiYdNHwfxuhCrHvoWiRF+5lzaX8Fz3uZBKP
GSVadWX8GT8SLbc9GRvUcKrdC39giRdyHNiX5Vql6ZQqfV204pXP3XyHa6mA8yBiRyoDWlnHz4NQ
5jXbZZEbo5If42gB/wVpQhuxnMtVWAH7BwZL3RDk+wbjDVysh/MbE4ghAQfjijuEAB4JTt50y25B
hopbaJwfQPgS21Ik01KoRTAGP6qinLrO3heh4Y9/tAYShHudWqLJtw28STYwA9UJUsv9cOBo1QxH
qx1FVn1pKfRVnSSP5stz9JYqSTg2b4AndhoeL0bfL9uT76JWjDUUeVK85td4bXSUKvBgEDMr09Ja
BPvb4n+fecV4KEYBnb4Rkw1+Sb1w/exz2E6QeIy/ggYklvGJEqygFVMVXizWq8tyzdt4locJ7Qhv
hl1ZFwcng2ASiw7oV1+cmgIhMR21qhlIFaTCIBGL49QN0eUhjOtDWDRUNJSSfUYSYCBEJ+4kwlpx
1V/MpN4sxMwNGozh3IUFp7d/pmvh+FZtuTeAIFnvNEQrhQSQ+hHq/qHxU6uoz0zKHkTVpOoIxZqa
hEj9iBqDRAzu1GizJr5cl5oUufnwoToHhrI/xznF3NGdtTFav7rC4MJO9a75uWyIEw0NUqZKhMSF
gWDxrZFZG19PTNZNBB9Z4/ue2Uyy1kfxrW8tqqK5h++4Xw0RxrEjv82/b0MMsl7SHWsCVgZRKghQ
fRmhi+4jQmM7jcu4d+A2w5tigOU786jQCEcPV27CLLzBhZNa2N2eiwcxE3SFEVpF31xDKmq6/k3A
wgG+FILvoo9AFkQSQXlVSgjGbwDY/zRGPS3sCABoIAOJ/+X0kYZrriBKaolA02GuheESbNlkd113
Gy2QsiT0YrNELpwZ/vbd45jFgV9JoJZi1XYx5Uv/Bs5Qw9sVaPyVzabdUGxUvU6UHFPj1/MT1A1V
ZLp7vJCa8yUXidLvg08BJEsTT7DudE7HdY7vJD+l7dD6FqU6U+wqIAEmUZV1vA/BVXWQFvK/O3AB
lMZKsL96hjiE9TtDK9TNOqL2nD7YDLEkIQUR9gPNyq26s9SDdH3NDLxmwuk2+iAWPBeqIJ7N3snW
Ul8tKZw1jXQ087+vgcTAwjaz4YbiQ2Zdkr0NrPx92AYxJYjHdqWa7fJd6oQXMvR8yFqBat0ROno8
W+kLp4CHtPx10Rn5gmiPAar03du7jEkkulZfPCu+OWbNYPvG3Zi6shQDP8Kk3MgFgMNOrkam0SKf
LH4trhiyq7FHG/Zoz/AamLCRPoTRfr1VXN5VS81E+dp1fvdP8Iixn5LYPOwmfxEcdZwEUdRtSxId
APOQKfyDLdgdCxa7bCho7n/mxiku9XUiBrihFZmJkZXeMpCwmmvpLUzD2cD3TOReXVb1iECl2l7R
Srsp9ujJlwt6OGBVrZZewaGkH3I3Xivzwdp5s1qlZPBv7JFuDQXRgz7u77mWAKmFBJ/BMcE/YTRx
VIk0+YtNxjAfX93SVPbDFMHD4qphyh5Agl6Fr+tdxo3huhFHVHqAS1b33+vZLkIG2mF2+arrCyIR
jxbdCkTziyjm89U1m3DSwJiyPMMV6iFtVc65fFs044e4XlW/TB2tVVQZtUcgP0VQkhgJTexPYXVS
ZYKT/c/6mrYaC/qIFXZ68p9Qc8bIuThL49q9yCex2Ml3yn2dkNetLtCVAAZtkw5cbGjSSGKj/l+2
+Y6sJd0rJoBxOdw0Z9aW2khJKelkZI4nFqBs1j3FvvGsIRigEnM5c9efyWd8YDC6PEm0Bl9DPe6I
A2FiDvVZs7hHec9ZFB81fKOvL3Ikr2HdF1HgCOQTPGwTWXqfr85E5s3czW+HUN3hLakAiA7Mew2c
W7JjVauG7ALcHAzDPnxp2eJTP2PjPk8wWPFIBMDzOycAkp+0xPzUXbU/99WOmpCE/gKHAFUjaB6S
dZFqLoS9M1mDcNEneX2MK813NCMsTjamMHfXRhxUCULuTGP5VU7TxTgKON85oi9GPojF78hkPlah
Nan8Vdj5QJdn+pv5aAOba006W5mYJ7a8i3Nf51EhGR2YMS1KR0lf03yDX6fhlDfBhqp44JW8T5Ht
CBpqc7p7ow0DPakuWzTOyRNun6ckVNmsYR4wB/vm7HUxzDAPO9ZxbG5NVw314o0MwEwkQ5GeSUIN
FsQC3wBGwg0niuFcjwfZleH1uJhyhF35/NDCBOQL8SZjvrlClPa07L3ETYyhIyPF8sb3cYt6R65z
flsamxh7rLv/Rzi6GPC2PItZ9KXEx3UYQVBYUDRGLSO5/ov2XWR+WH8nyLMc1kic0NmbAEJ07sVr
DIxBA2oP6g3lagZtomqQ2BVcAHqz91u005pg9qw37Du/Y6bGSmWWR+zPoemqHGrNxQpL9L2pDcey
+PVOAnbmzrIge//ztVigPGo18geE5OIoDfhkt+kJqwn6TYfkkIFSwOS8XdEkDyQr9A2tCxO1zcyc
ixt1/9a9XXFuBIR04EwkQ+zExJQ2OTWUY6Ww62ieQYOAdxG3c3KBtRvhJMUY1iuEbaVYaTtYmnnY
Q6nPiyLpuJYgcFQN53GFGVEYMgzaM2O+UKN0lZpQPYgLz34Ng6Rx+LsD0iGPVILxQvFL9TE9nwPA
yOIclEy7rO9I6SCZFnBf1PxF6xz9HYDGmatj+BdBGGyKiBQPniQSWeCgw1TJP6vY6ySS4pNU+Zdz
Su3y2IV0uiqWJSp+yBDLZeVzpiYmC0K7LlsQ1Nbo3bBema9kCztw2gd6p0EL3oGG/bYIGX4NhcKO
2C4B9ndk4BokL1LcJI1+9TvuRgMdwMslVTS8mSTWAF2kV96RDJiLu9vwWCNSUiVUdOnDwIuL4rFS
LEeu/7ZYO0izQWsaz+JYPzIVkfrh0viiVoivkC7QhqHEoJ+f5GubfUbEgOqcBcoc/likzGGNia3U
ZQiB2SBN/ZhZpdYXJPu+HAd7K4eGWP3/UM4l6WhALdHbmQPiWXpEtawRRKhKlp6Wp/PqfnT10/MB
07IfJ53iCJSFQEbAYP8NWCZkysNEpHYMJNT0wXzsCMV/KRJ7VfJJ9DLEbLkJ39MiaJHqaSHBJQaq
WdCWynU7D3eiagKgatm9hBCCKT/dTsl7JtT0Z/A/tjBO3HzeyrHw1pk4yHjnmeeJFTojEue4Juhb
CZ01UbUF79viD9HgwsU0dSqMeakGC/f4tXkBEeEGRIA2umG208oGvp0XyqH1p5eZorNIWUox76oI
Hrsy/44ZqZh4WoWcgBerv73esDjqzE4uBufUKdrWe8qc09hf73/RbEpx7YY7YJzhOEPAANbT1aV4
Q+fFgtCk4/pfNz+NAzNLUn42cBAL92plBaQ0qU+yGQceaiNvfc1esIOQ5Zn3lWgy7mTFiLuElQNZ
SSJRzoqfn0aSnUQ0gPiG1U5egc3b5rIPBKJe1yUKYM6zakUbqfKw4KHLwFHQL2binW6bTtZ7eri8
NA00M6bjiOD8KgxBUtcsn9ftfnABG7sbngWiWYv9si7XsUpfIWg8nWsJFPeHwcPbDVLJZSQ1yuqz
fAkKG76OoNzkkr7kxlPrpqgU7VVBgGyEfRZ+1gppQwk9mQmVGxr/v/pOxc6XP0pxCsgFf4bUjdnR
kVurBz3AfHXwsmT4D5gz6VGShb6Emxq7BBbPqb/lLXZonM9u4O+2kZS3mL+IxDCJ/bNC2MjG7LnL
mDDXC//QXmid5xm1EHi5dxksm0yk27P28mbLMrgdLWNYtoJ8/IZ9C/iWMQKh3f6LErk7ByxXqFj+
K0k72Fe0cFBBoLodRpvxKV1UNmHhxm7AHjgB52fp/MawvSR18UUb6sgBmxfD+Qry28sDQVhFZanr
1BM8D3zpDgOD+S9d70ggHqBkmQjSSqOEonShB+5QmshHma2MFAZe1RC5exdm0kkVY9YXne4yBxK+
c7ZKGTrKpY9gwoaJZbh0a4uQaQNKFR+vw068cWP1lC0kTgE/T085Q1hcy8ihELjavZTfiXh9s7QI
9m7eN9qAucJceFzAzmAHzCnx6RKx6DVH05juNZxa6jS2bbs36Fuki7v03UuP0zUL3e2Jfaxg7MSa
OmSpsxh6U2xq09WbTrKzemSCNwmE4I41hqmIdqu9nqvECByvgnW1CJSahYgLN3nr25pzKhWHH0ga
EDCdHb+2OYwz+NXELOYLHx0ikReAf1sHJQvBdzgkDJOYEC6tbZlhP55ulJ7UQ0o/GhwIzEssT7xL
dU1XCWh6agzefnXA0TnPWrg3nfWfTF8BrJaxf2NT7Pc/ggamhUswNeJAwPsAf3p+JYTmzBQm9gGs
DCYTqV5uOq3W8Fv1OTUUA31n+mhTOfzpz8Rn+OfO7fuUNoEq6yX9HTop0blSjCrMhtzpJeDS83+U
Q2d3p0/PX0bgT0DZST2umqbJ6BLta/uFpNhMTs3f0s5D9dJ98J9RzkOeIBS8ZhQ1Ko9MwUGNYEuF
Mr3ls5S/7oQGS6RYs/n5woglrp26+u+84VCArI4OLJiHV3CTXoeQnh1S1XMm3/auQOxd1M298rhI
4360qLJoXHGg3nQbhtQFiort3kcI8Ks4T6HNekl5t+kLSRktsdlJ3w4hoje5vwXatUI5lOPV/hfH
KcYtfKhNRUDPmX9x+5rmK51P3ivdrVFB+7G+tJMWbJM2xGTxyH5MpRXuDkUxpkCQF4WjGxB5GRFZ
i8xbIHW3O3SNphJjSSaWLuOlqy18aZctL88CSvuv9tsiV4sk9rpH9cuEgRfa+14tYJrzbEyK12KG
qhAuGnmZpcjse4/b1CqX58xlFW+j928RV6yJVRCO4yvWP+91UqXWj9QeqRnIoDRPXo2++mgy1AO6
5iZnERvEaLjb/XCBhyx0kH9sJBHFoB1Vj/n6enK01UWarN0/PH/hUKtYNT0fxPKwD/CFMY0AdlEk
7q40/EV6XsCorfQDeouqkMCWoTR4IOpNrkvnQJkf+KF9A9eFEHe+eqtTfJGk9JAjrceHQRLB4aEz
XWKL3aLTdzUSHGbbnYsvc9s9iMjMPsRJ5LEhrOWKUyd6sZ88M4TeORgj9au+7BIYEzTJ6KpaWNaj
jTD7hWGWprV7zszBla07NrOsIvGAbvd+gNtH8KZFIFJPz4mTACIXtiemeafybE1hTqWjme8hrgVW
vhNRZSaRLxH076bCHu2kiYyiLTr92+0LBbKxMf1dGrIJANlIpRPM5jkIG1/txUTmso5+AM4EPq+x
ytXsZTEbniPaD47x08XFwObBSNztvxsrE3P0vmmvE2T3eoda9N+jCqXGYp5gbLmo4AX5vJBYnPS2
DcmlHczkamKOuJyUHyP//rbaHernP/CBzSfhLdREfsUk3PwKaVDddLaJLh34+mmcnXA5LWzARSGP
jU1uVa5Xs7WcmDOtg5y5ZQXSqM5sUa54ZK/Nd+lBOXsbymh38/w8qRYrtmqJlGgqI27qFwbFX7wZ
F7B/vV7Z+xCuqTtmbyQpXwxU5Q2ug3KqV9uFjvwLNE9bAsHaT/YYeIzdhLleOBJvvk3z5KORg+fq
Fd93kEP5hmkfHzH7fHSqm1wZ4w9lfch3Sdc7P9lvG1nvCGtemzF3HOAUS7LYk8e2JZYBlKMOoe95
Sf7MgVJCzad5eLLp+3w1Q0/+xid1skTWZIy6AkpOoHtBV81TFQGTJG+XcYY1WENpRDO0AcwpS3xH
wCns1AU1BkXM19aUKmab591miCRIP5jKjpe0SB4hXKL0pKZweFszq9a03+YiV+urBwpz9wYcL1U9
2KwxUiCCzpouFrgZSp0suyOzWnCHEnAz6mgyQBcPtjcFGtNkzHTb670EeqoZv/LjTWwfngj3B0RL
tVk2Dd31uH6EGKNXt29ct1bHlfYF14hdFMsMZJ/BTJE3BqQAhjDITrKNIa3VE+54z2Mh4LXFfycf
tyKNIOFxsvYlgdcqlLcTrYmolgu4sEwWR4hoEKdFLKNe62SjlwBY3ePM+wvZsUb0TvfsCOue96aM
EJ3lSRkCA2lTeOOFd2VHcwN7ruNYA46cADiQOGT7qx001VlE9lAsCrMehbE5DOSmNbU4fXdMS7v8
gc0vNenf0i+b4fSFltMqiX/evsvilFd4GP+rPtF1N6hX037Dzt/t06YULZm8knpU5Uiw1NijUdHz
/rsNJglnfiOEk7YhdDw1Yru4WD6QIBCkWuof2rLBB+euWNuUcd0GmJbhCqQBCCD2Sdzx6RD7zF0A
dm+mi8N/C1ZRG8oQKA2hjz8AThUBb7RzvRCNubpaLwL5SkKBkI8waVvhnk3e8wmx4H9z0SKF+rua
vMFBAGm32oI3QFQfNghgZc/lWlLDjYyTg16uviaiQixzAmRdOXNbaEpZijwMzmQukk/J/OBsQSa0
PHd07M4odAqVP/Wd2UE1kedPAwMoetdNhpvr13r5g/qhnGzAB7HWC24+ejB6pGl1WjPFRZ7IcnpZ
9yMMD2UBvOJZqbqlupXrHLMEHorb+afHHSOpSf2MKaKOmEBkj5YbRHtCkwmBF+UC3RJbWGOV7CKs
OkNJ6Po3wEj0FTtSOBCTbvH3s4FyS1fj+KsbctkHYcRQXvEgJhqmpFU23r9OKaTVo1c5wFKZulfX
OVGYkpyX1eazRLR2BYQZonnrH4rwjeU/jWwGOwGhvdt5ZRWp0QBRPtp33cL2HFJkyzTlooG7de/D
i+hKBMRtSG6hE5eLKk21ue27PJdJ0BZUQ6CmDLS/85pW9idQBgEPUnMe+om8CoZxdooNl7EWeXqN
/KXY2wEMdBkMRvCUjgBFK5TXv7qI4I+9lqI1GlPa5YPTYTG57DoL3oR4Ax+n5Llq/fl7oL8Q+x7r
DH8eFomZKmsgo+Yql1mBwA1X9+qw6NsLV6tRBoy1XdB1uvEFOlbYJGH5G485uGXuODvDKEK5bQ63
gOMa3Iqk7aAUY0HuJrQORHHkrJLfzeF+uucPT5qSb56TH7XFykz5yGfCcKLVnt3vPbk+F2trQ6LX
skTmNRBvIZaCxvSMGVeq7f36Bl+/ZLUfH7gGzaVRzkcKMgQ3F6LionnJh/DHs9YEIl/AyisGx8Yk
Qyu4dJwwigRdb9qx73r9O+YevFJOpgDllEVklU9+SUwu4PqO9pDtos/tQGVS5cd5Ys1F5MXf8MfE
91IEdlX+JiWwanS9oS8DE5VjvdYniEUj5VeWNNggYnAMQvbz22ivCbmt24mH6kKcvs5s9DZB6mrx
BdgqewAyu83a4yVND+SPEDBhNNzUzxiEc1de4hO45Rc1MuqGqKzcBVlav41NYJeBcAbWZKQUkrkz
yPPDO/YuCP4wMD4IGnXL1zD9woB8DhYDTf6xwYadjQ9DmD3wdLkyMONTGAMIiH2/agnHFyqXt4wa
oAb1fcWlC9OtpHWsfPKpw8DylRg/wEpCdR8Pj1ydVghn7AitIz9spkThpl2YPMBjgDheTBfMnYW8
zrddSolAu4AlK2Tk64u2h6pS5qpEc5bWKu5M5Uj/qLRWm9vK52q8vvs701TTytLxfPXVEi6BanlP
DkOk32e8R5F+f0NSB8hgXs9eG6ysV8Nm64G/RHDKyfpzXecEoelG8VxHlNkO7eyDXTx6JfzxIMk8
8INLTQYFUJtbe+We/Y6dMafUiNv1FvRFS/LaOYQYwGZgumVeRfc8bLO4XsNYbok/8aveAExiyA98
p/ESs3VfTdlDBZdHBVBoRaWgFXlGwLwQW/ipyKLVd1VCaDfTlFPUcSwL455zTEaq7Kq32cWWcreF
zPB4oRdOBQdc91SPaDh6zbxAIJSi37rgbo3J0JOXD8NRsTwmDUoaCjn5EC5VB0pdTTegOBVJdJKu
Nv1wZoh1TXEtmxXe/++bNC/ua1BKi0vCOVgUAEOtTndp4iNwsawLyUAsXzcaxkitnGdrM+IHfVUJ
3HBOwpzsLkJRg501+Fqb8zldWH43vvMbBw0ZICpchPjpaU0njxOgFsc+ZFGfM6P/fnr9XwCtw5NL
Oh0p/vGDI0/Evhrl3Scn/MoOpK1mnHsgjiaJ8QcxcL/mX892Jyoi8imQskvpatomLvXkk0AYLSvZ
Ti4XlwIjta47eCS/QHCHREtiFHlkGL7O7cXxU1Gs6fXqAJfxEN4uPm+xlUX20tyVtjhY3p9mRnlp
bQTfe3Sy6eXkuup1JuZzN0Zc85LqZVYdrz+HVH20AY7bSJehGfVEKZymbyTJrYdIBD3k2wjXIwRe
Lc1M0bIHVNTrjTOiWRUpTOTWjMRxZ7CnczDJQXTNqZlc7RQyPlW0Kz2vIHVU8CLma7ir/nxiGNKb
djNtd56W/eZ8fQ3Wf0NTIzoSuzz2hMvWy82ci1gHDOpnj+NZ2zlmoEfomRZV+gFkUlsnVub9gyyc
1GCVzWzWmpkGkbyOEPFhskd6eXpurjgWDbvPiudKLcGJpxpvr35LKEZv7X0pbLeZFYaluE2sy6Tz
cyv+JRD2+N7hEiHG8/JSTsDLUz8lnpYpuiMAlATwzMp0FvvLR70X1ljCb+F/5FmYmRPOxQLQS/dh
09xj515OkPEJy5MaG3xJm01Ts+8sAJJ3Lys1ba0vVQy10qS0yvgKTNZacaNvUN2+Z31O3ZvWiowr
e4jwmXebreccsVEvNXyfF7vHUSLhAffFJ9DfNiECIApA2oOjMJYZffHqY7g2ivADr6FaLjGNyJxQ
tOtvNSDz9ssFw4s/di3r3XVphbdgNGuE8kkl06jLvroUkIRnRx41syU1otIJp3j+WvC+xHvfpqqv
clRkW3f+z/bIgpKsxOCRN4dkaJOGRGoPRaiyjS8Cr+ntJA8fh0H4jW2ktT7nlMSo+ZX63yVdU8iI
9B37q5wAylroGGW9uKjeE/o60vUD9oMAz0hAB1e49a68srM6wFSQmMvL5JW5mMz5djFC+wDrMBFE
rYCeWCz3xstp2t4iBtTrw3m9Tf2Ofvh5r8c8aQQK0fMKrzsB3x0wZqVHU3zy9lpFwzGrQZUExMXk
cv8pJ+yRdcoD7L4xDbD0njAiUxQ0VDIkHDa2iWNLzwKl5AZj4sjekhkHGylIvZXktg/IJeUd+hAu
o7lCVyMIWj49YWmtzAers/fjsd9U2BQi7QP+2NCiWEgczYLjdOda8n3+fDvyT39nokMk5Dh4q75w
v9+Vi5cyHWFTbTrmcJjalqUrj4iB/TWmVXTclci+e26AlyfA5ljVxFvdXMoeSrTTayni943kAscj
Mju6nTqw/uH7qu8beFmjVzGCoNKRiAsa4h81qSR+eU4YAWqEnskJRZkoS7cWL4+kY1kgcdQnM0td
d1hLt1Slq18HThebXdhVguEUI4W6WS95++6w0K+g3++tqI/ptwT1ZCIQ3GVO5Z0R8pul34Tjx/qb
L74ebl+YOhYb9V+mktTO4IODJMqNUPaCeXEtGOA0n9faFBstPjcSZ87aJqF+Wcb+G2GN0A1AM6Og
xTujmDcgppSKpkhFkXEA3Bbe1WwtvrBQNmK4C14hQcxapaiZ/zhajazqPNuNRZbiT9CokVyIvKuI
P/Kjr7SBvyqWOgyxkHQ+K8P/9z85O7AYaV5mnCEkp5Xln32VdA53ZEcEiHcthuxcXbrAiw4mb/fP
/9k/eZmIZLN0UMVzMePq1utH0CRC3L+OBaLlrUMW4z5Cy9ilPJP+ZVR3kHLulzQmReNHaBkgBLoG
zkn09E2i59a3vCSTAo9M42W59mccyCWmWy/ueZzyWifHVSs07B5gyihLRgooxa/+COH+j2x1tKhD
EYWhr6QZa7ojJkKftACjfiS6Wv4Mc7pMfZe+Tm5ylMSMrtidMYL2QbJE9+u8XvC4jMWPXeZLn5Tt
Y0zEPuQhqqeG2Xn/Qc0S0xj5ZLwbo5BieILBx62XoxBe8LiRQl/7LfITPoEqeF2a1nAyARkwgxJg
bWfhOw3pOigTvxAApflT5LdTg/GwyzrbrMHD7s/bBeax/TLBGNmkyPPtWG/rCx+mhQg7PBJD5e1n
EcG9PsmtA0lEF6et+YbLux1LFcp2KFgg9SmyXXbZcKbYK3rl4PKFpH0emPS7X+SwagD5fcEQG0T/
ezyJ/TCMJO3wg2j8UHlvGh7QEQY7z+V6CY//cPHup1rPZVMZQNUCt1PMcOrcbCGxEq8vjUVN17pz
SL9x8dyBHQAGDkfSXKaWD6dB3TyzOaTWeEj4MHDvLw8B9JEoCKKCBbi/AAh9IGOJmGxDkbdWr1yz
rH/cAMNHJQ5mV2uZGGYELE6RRTz6F8LpAw3V7OIcwNn9jTTQVWCsD2eJ/WD/GNRmpAXXRBAXVSpg
OqKi4Yu7qLV5gxw1c0lUcz+yg3IUq5VPkaAy1TTjveSsfiaRw+jBmW+NFFtMyK3fK2cwS522nNAQ
WzfEqsXQd90evq5/uHQZVN0uvyvD9IscfN82bAWbiNHVEAJXwH268lFja10w2kniqGJJo0Pgn3F6
xyuyfgBmcx3LlG2nNhjf4IZg+at9AOpY8wCZG81Ucb7xdeiFPFN8mgr4yXr/rZsX4uIRVSXbGF5x
VyxNiE79QFkn4WTwP/+vMZBK9+qETZTU1C4R8j7C1LfsLih+v90KADOe8lK3offQ2JfVk2btf6PU
yVvPyq4ZMmHYlN0+aVZ+72xwi67crjONXGAjtXfwopDc5u3TfTwhaC6FUhTmFoTMrOyMPmohiEqZ
0pdOkxepoVEzEq+mPGtk/pN1HpJa5j4n/VPRrOvN9gyAkHkJqmhAE1wNqXT9HrMCJUfL8YBQ2jst
O9nluinjPmYOsohA5OQ2V1E10NUToahf7geDtqP6+qPGsc+mEiN/aO/lLv5UZ3hDfPzkWKiYEfaN
FR2ZrpRTFIzRHHZcp3ZNGMSHQeYvdkUmvxVyMlOIyqnf7QAGfSoxPaEJOBGA9fwmIsWFe/V6IFpI
CVaVpV6alxKWCIsnc9+rFPKz+BDh1fCkrkHFK9BSL/9DK8LbE7VX3v4uYh5d+L3r54GaNo+liO0k
2R/gnk0awwChjSn4QZZ6rOYZSKW9Y8/H5phEK8mC8lddm31r/84BI8TkLID48yRIK739G8xgYGGS
ZgtS60+W8gx9Y0uUe47VY93YvSPr3/K0zPssk+gMC3kyTHwGXyoX4c0DeVtzp/832Qq5AuUrZS05
Phn7u6asYlbJKxooqZ3Pn/DYxI2ZEM425u3JC/R3om5hnfp2jgYwSMoRnHgapmOnBrLSddC+Jji1
VovIEYvda7n1Jc8LNU71FW+8+yigfLb+f1VqoNU2JKKOIcAf6QKWUf+2eglCUZ44qGSDNfp32lgP
WzAOKioaJnptzyp7RAYtgUoV152E6aSgY0CRlC2neKxKURLPINgBUB8MkOghRJ4hjY/btwZEHoyF
enXnbbF3vdobfnaL5/4Lm1bf5kAQLpx9dVE9kuPoFl9JMRfOB0Zj+D3B4maTUqxFAlgK/Ogjot7F
3V1ZkDte2SxKx9p/+Bu62q10t3FJ9psuCSKD9rfnmuUVBKCbY8LJdzVBXwGQEsmytV3hcNreWwBT
WQ+JOxBO0L5bA4q7GKcM1erjQIuGmLO13RjIVBL2FGJQbqsm+MdWXXyOJbv55ZDP6VdbKNPchvVi
8AZtV7f7loULzisoB6V5xfBWkxW6XmsTq8zNoEmsdCYCz8p4khcY4jtz7zioaOl2tyUwoMoj8gxH
/T2wZGvmis4D/1w6n+POZp4gZwwbTGnvUm6pXzpnnzKJgOidhiwpkGZEpnyvxyJERcvVA1MZHccn
NiN5fLo+8yTVeUJGc1dXkZjSSHoT5tF1Vjy4Xv+wcJyKEmc6kwQQ7BcAYRaDyWHg6+7hbmMGGrvn
VOLeyu2HrD80ATxN02vK9cw25Z9b5GR28AIdK+4ypLUw/xmVc0ocRaKIwHvC82qm0VLJN0TEzOiM
y9RKXgZ3yBgSqcywutY5fmjprUoyPAw34Hiy3TWpGbEMMamk+y8S3VcTZvOxdohxHAFlfFhcMyW6
tmVB2+P6jZri0TBnFxybp+kSJZkY6Oq2acpV9uzG92cUgkzEzSy+ibjXKedRxabAOLvbc3iYvDJ0
C54gBnbLL22jUCdx2ea5QANSyXwPQjo/LoW+s+8+t5rH+ijHn7eFTtsAO3bdL5YoMbu9qcGn/QEl
9RcJmd9bI2N2hcPo+V2Yv+V7WuWaDI+UwVzAlQTTY1dX5ma1F1d50xgnYJwKnhjMqHC516C3McNQ
iDmAApq9gg4iaQf3RQw9aTB3riifW+qVd/w1v9LMwQXPyXNjkC0JUmnGurmpl1iltmz+09Wsh4Fc
0EIcvOhqyJ16xGL8Hv4CuBaBnelSGDyEhXPPgAe3VtjdUbsDTpdsF1H3BmFwx8iaWJ3krlXLJXWe
3huKru5vlW9rF1KNXyp0Mx7YhVq8dU4kfBvXX1CbwJf8T02XFpoYlqVhCla+ZQ6OjGCV6okkDYM6
pdV++ATQa8Cg769/S1hM1fnC9AtavxFruEyannQ2d8RvR4ekFE4Sqw+xMfwqG1f0ti7JC8PktLP2
VxNEKYnnX/N7A4+1DqewDdvirbmeEn70NMA2Iun60T0w6uf5/ApIZdLrEjw5v+6oPfR0OBvQkhgp
qdBGNik64bGHDJtXOvAdSX1KjlQgK+r6Bzkf78+wNGmqYKes2GSFpIQNQfhlkViP6K0eGo/m7atN
BOKj0o7I4LKru26oeJC2RedCrQCtWIbkFrmlo4OCLXGlcGpxFAc7wW/e2wPYQKZQNX3sLBv9h7mx
wEKFGxN6oKjTfKwH2+Hk9ExGQ2JDWVMXWya8LerA4egXmGM7HLqUl4DRp7upHQEnwD2HLiv5RH3q
o9/v4+hYj5X3I+q+m0ZPrc3kYq4I3Lly7fq3ndHwB7IZ3fR/v8pgXGe+19Bbn7DMKGuBBLhsG39p
mcKfa6fo+0IIe/75oX1CIhqA+ECA9mmQyWXmxJ+60U9EJ8mGkg0/7n3oHHoTie3o0pg/4IDFjN3o
SkpvK7XZtA0cnazZ6tVoDbsroUW7i/ZlAjX+gKiGx1UZigWlzOwkFHZk5/wOAHaqnbqu6rtPlqk3
xxXu9az0YZS/27iIv/tvsSbTO3/RMvilXczQvWAig9vtOy6A6hQLZa9Jir/D1cWfYEj47y6xiYUJ
u4F6iEQp8lsprJruDYD8BBuOpuijAgwTj/Eyv+viYzErjK00c1ng4LmX34rOuBXnlF/CgR9K61E5
Xa9ykVEn9wOSUh+fMPpoPiNOyoi4sdzt3ZADVP27Po50YFg03/IJnNTxKtYMg519DjSRYkYt7hEu
7+jFG0tzwCY4tOdSYwFHblUwXOq2u0Dc9SRhjeWx2KGf52q65+YQmaG/MYG8J/RjkmLb2DU5IBhS
aH+SiXxNJaLCQT0fQfMOGFBPwk8D05fwLYDKwgVphvKTXSVF6atQAZrumxKRjwdf+bBNu1HuMFT5
LZRCA2ehd8g2Pid0HSfyrNpgfkc+9MOeNzjX/uY8bfNbmL2Gqp+D8cqiAtGK7gkagJuxPgdfOpKN
MsdJLUtFZlXFrfZd68u2oVJmMiP1qkl17KCXOxirSOiiVENqutM9gbO/1YO4pwBbgRfK2Yc5Dzjd
LKE61qm74c8vJrsJk75a+mnfJjMNnoaJ5KpaYyHqqQoTQrZvu9GOJb11X1beTjlZkBPxXUtXGvbX
4FbNF4qQccEXF/UO54CP2K2RgRwWMjtSKtmpv9FQRWOoCNzug8JwQ0OkSWvOsRILo+Oe37LZ4NxJ
xVpjQv5yytswevep3oFhU7DmaZ08UrnIoSfahzqfDaKIXFFWt+ANYEIXqI9wETV/7lEC76mXhZLJ
q6o/iHBnqCrbb86aM0LQevXCOFW4CgUCoqejyU+d1Me4nBkdzqCUTtpPNPwoz0wWZoSEQtoXB4aY
01ZDdPhnDhsrDj58HSGcg3j5Ti4LPQ/6hXNIRUVgF8pP4JWsbDJF7VnJ4zn1jMuVn6FGSmHaF29k
5gr9O5ghYKiKxdEx2MdCcXDvY5k/n4M5u384ShCtvsldLXhAWeJsX5V1LCjkv0Y0p+fOaHnAIgHs
u+C971NcsNX6+a+6TbEFX3hhJONQVZwO9STqXetf5W7/OIX2dOwSvIVAJm61ojVdujJNZj0dnXOo
btA5fRchgsazWEQ6DHvcqDe4ZpEUq8WOcv7yekdrsdOKRSEm1f2dZk6y9RnsjsDOJ4WFBARz7gGi
J8rqJGhKteSqyjrtGVz6B/+cxSU23FhDe1++0ZU6kcFgzxEJkRN16p42VwMr9z6m3q5TeWGa3jUH
WW/eLiFh1PTJ5K9mnk8EIGtkSYKbvlUzf/+wRQtwwTxP0a32eNqoSm/iluDYe6FUcLj6UQ+j84VO
iv5gHb2Y/0g/dm417kg5GA54VhnnKzu3Xu0j6o4XcCPCbrxxO0l6B50Yjqm9p34KFd4pPt5uOids
KJ1cKo9ZURfJSnWi0gSLMGHAjPUxpHZM5oEh1jfIyJ3aSNll8R9t3TgDahf42oC5KHztNpuW0vXN
H6XCeSbH1S/G1JooQmpPwCjc4JfMJ9SE4WEy+6T2js6pbBDz7rnh5so7trM9kwazOxxOuvI0Kjjc
qlT0P/laKTe9hDcvYksYhnVvYEl8i5xqADP7z25z0GLbhuQB32QtFGbEQvTUzz2wtZBkagSCxkmp
IK0cByzFbnPnfWa8fFIv8LXCnzyJX+U8Gt9Hn8QAN2HogTpaFdA88Idqlie67m7dZ/Ut0w+/NcP/
1rqLh+2fEFAMBy5/YikI4Aim0UAr1QCp9weMrq5SbEm0vLZZ7g8HI+BmTZj7ugywL0FIAmI2Ydqc
2rxYIVKJvJVsc/h2JiSXSWUFt8PMr/pHztt2KHDJGzb26Bo3dy+oqI4YXDX8xANxaF8rCzNj4DDA
l8tezgHf7hdvocrdhJCv6VaQ0w2cAAc1TN1GormO59EgTSB++yHxzLk8Om4tj+EdyIRpnQgghYN+
r5S2zoZTQEiXvP3ftkzzAg4nJzKGwGfWpOEEaUxj3Nu/so+nAoHxHKZ3XZyLpZvTqwpZ/PHYGgMG
0VLcb0wYlc+3v9QMkVooKf5B9UHRzIVWgG4+0zDMZXx571wZxbnWLRG27UCBwwfocpKaUGbBVssM
ouK00nF9OvGHwfIL2zf/aVIPWJ+ZWb1wm5jYb4+otLBt30a5Q4vBraf/5yUpyf7NlDyPgnVK35d1
QPN9HvamXYjoMYoz4AtCiYBnRkPIhOwaOUs+pL3aLTmX7Yv14tBJuVBhNGz7s3CfzWFwuZHI1QYg
PEkV3DaDPD0GfmXzx3FielUQHKjdeOxsG4kJc2wvmXBfb3g+o1W88tWE3WmVq7F23ym1A5IPQSkU
bq4+I2bx+cK5etvXmURHcZNg34qxgCb/lDPG7yK1Y3tx5X5oFMzIOr+99HIr3iFcX4xj/EYkHqEX
m+Q+cxM6JK/zKDXhb02Gn2UlP1j6KnZm8uPxcepKba3Cp5Mf2WmUf0MCCphkFghEc6rGMeiEL0ul
uw3XAOor9eR1canJ/Zy365CGSbD2CbBuXWxaGSoqumtTyLTc6yYG7iU+ebO3lmCA02QoeH72gYH9
WxPOV71s2KJvvWQREDMrOUB5GbbAWvOgvm95qzwTrt3kTUPpvNoagEslQW3GO2sy1roo6E73i2wt
kTX3Sko0/wTQB4VVpwrWVGKULrQpiSn/2dGjyofb2NOLFBe/lF2J2km6XtLnrxTyDsLIfd8eHGAF
8BI/xNr8oZdc+OVHLLnwGVJ2CKcmiWBfF7/eXd73700hbBC0k1kN90lSQUx4BwsTNCR0awHHLxOi
6HetWEMPdFKFgjASemvRSfZcWqloc3R3XSzdwzPEPVnLQ/OccH+9y3sxI1MsOhDASnLWWDYJXxpU
e7IbbRk4MeN0Ob9yxdwJKJWbc23HyLxhUd5WmUR0fgyNPh0v/8NeF80GHbjtLGBd2urZ5TIQpvrT
eMwkPzwPUJ3LPPzaNK4GtIjS1SIQFC9kpPP/CLzkD3G0vWrjE2T18M9V6gUJDQTg9RhYxbJJ70Eq
ril+Ej44P1jP56o8dKkhmUuIoxD+4vMsuJzMcIiDNFJhApAI6vpx6r7cL0O7OHdofYJGRdLcjaTl
iIoj04Ld+dp0ysdE+XURxJtkdKbnapJ1rOW04bo7FsOI91mln110jr9SRC/5GaFZxOuSACuD4cds
YPbcoGHVY6XYJmSfXLbsvYyJtspsu1z798uIHMgvLWUrS+3uoM6F7zh/ER+leAXadANBme4qQcPg
Fgn2xRW9519qO2H3rIEncK3LGgZKid4VO9wTAtIFC1EXxSapcAEqewAhy24QSHAyze+d3e9Fv6ee
LDTFR8v7ni8cwgGwIQrzQMDCNyOVaTaMg9a+1pVb1h6Pa+Ql9MnL/BYf8AMgYzpJVQagkjGk60fO
BsWV+8vAD4ZphDfKngFmcGIZmDvkE1GWtOgXC/8kmOpSA7OMquuwJYKD8Vc4SEszxvHsD73yRvB8
RT4q06cWLDGJPGfosXtBkYLoD80s/F4A3NkjX6W1JecbVpCSq9iJjh4333dqVZvLCHMrJpv3K5hj
7uIV1c1Wkl2/G7+bbzu3wU7QFD0OvDIScerA0nj7c1zVe3tWIpDMcr9wqGUtVt22YaNcWMqqG2GF
fVltrlAFSrqY4OHqqwBGbYHRFVzznCrtHQfzegd9pjjULFe7eLsGhKUEu0eZ/CIv6f1JhBxc6DR1
XB0v8pdgupEMJIbKw1OBMWCiSnb430Q7GF6Q/znuW10ag5E/jaiUIgU6mOoc0gkUzgXIHewqHLsg
msYjxa8T6Dby9anA4FImqmvWhX20mUohB3LFYBnI8dFXNo0nilXAe5v6v6bIjkLCA7BCoUoJ3Cxe
ZI+KtJVz4sVkyOuilPEKMdU1idixidedATr5QINJmfGaWsi/F1gIKDNLfZt8rTnQ9fV+lESPfE2T
Mz2Vz8zJV42cWNLYVWRz48a/5iYmhj4ObM3yomjLPTJjB3V6QODLK0AHaRYVQIAiW/AiBt28Ogv2
OMfS6LGAmlcmdgYir/P9Q2cc6LSN+E27rQvcpdHRBxZnnL45/AdQVMjEdo+HvFoujW8F0YVl84s8
MUmD/pFUpuYWRk7B+nm3wI7nNvAWh10VngcBIB57SxnmIHcJH50NVgioIr1aIuh0Ef7gtS4EZLbe
bbumdPGJYIufLftqMx0E0eogS7maDBLgAdJ/S0Ozk2kXae1rGy6mUA09X/zvUSZDDFBcZ+dtmKVg
+PhfnME4Y6iDnnXgm26AG0rvSHag0aVw8j0HutIoXytnLtbzSPqEeqeXAzb4Rxot0qgo7PcgagVy
NLieWqC3wJgS/UR48T7CGzH0KLk2Q4KoZHkyrDqaqj6uoPKq6tvk2nUWBGEnkmUDEaov6PpF7fkX
HWiNjMha0qqOOjJRjTBKkOVXs7qXNbIXxASjgMG6LN+2YniERxfHK8LqZUKOg9aAHf2R+ioKA6aK
Q22RNfNBOOwgzS1k/rnbLU1D1ApfLlmXhSFIH7tGMzaAt22mI4UnUdrBLlmlEfm+Bita68l91xSd
+j/3zdIyJZypr6KPQ923s6DUmzSBxzl+iOxpyF3ifSJxSLs0BLNXwKAZ9XV/JcM1PPa6j1pJpCcm
VJ7ZzRvuZv6p722HXij8eHdbdmWyP5WMiKVQht+sAsIQ55TSlL7IAR0KGanAa2i9Y6lmitgv1lU+
hrU9sPEix/WN3elO9tmjiFgOfTpBaiAr+MAXC+c5njzRFrSexa9BJfAOyHgnpALY3WZH360oq/O+
NDLW8JBqQxvysVtzXJg+gSbdJFYVOIgiuGYqczxLjrbgEVsPmxrm7cfuO1JEg/V3WFx2kixvq42r
R+v+JVV8NonAOFWjVs1duBsMTYQ6ytzEb5uo3BvLwl7wcRTo8og2JM0lYlbMkLxHq9NNp2aInbm8
SxONGFUxAP/C0SHqSUmvzfvog7V3wK6xbIcXEYJwteDftTnVK7Zv+EkpvoeWe5pfv5l0R41+MixZ
mvXTkB8ldL7MENno3bDZ/0x/CARDJdbjt4WHtrGYt63bu1/SauVzKJE9cXDuO4Ch1nXQz9vUmEKB
LnQooL8/cQtYmRh/q3Ja9UzMxNfbNyvqbO2fyIclG5b/C6ez6PUsjUpXC/xYXqeFyhScafN673hj
7T3WGxsuZQ4zCSd0/nh9JFH8lkN2i/M8ZZr9DlEiMgLzPmuJKOJyfbkdOduQ8BFxYA0vpkYz6cwt
BBMRy4B3zyzBdBv+6LpepM4X72ZbK+w6kTiXvVgSBs2pH+uO5ld+rbE/Tj0qV6pDWSDR3WW+4tJO
ts/QFlNsO3NU4DLLzluVkubamGbInB3VRtdSSlVrQCt/sbePOfl4lxvtRmoAkT7RB/To0+QJatHM
aUpFCs1pPMsaeZmx5U3m4vwnYUJDaL2G9coOT7nTvGmwGVCIMxItbUYrcT8xCtXb89Fq2y+pgySi
s1UrwOxogOMkAxE9GAc0qRTMUm2+OPie5WQGSdIG6Lm/1K4uxK4bvnrUqfVzFynaNhBrEoTL9R0r
UXWZES5VTVvngsZK2UBNT6/g9Ns9s7+/684Br70jTBlPnEN4Df1YXu5r6Jrp0+v0uR5IDsM0Kivc
7WaK0LJXSgeIALMxyc5TDuu3dbcQR2TttfFIo0tAnu7/yQz4FRTmi12ZHdhnQE+7dXliPKSb5GXB
CPRi9EIVy7UIA0P8Xf/mv6EYhHYlg5TECuUFkqh9pzjzcUDnN0uy7YsObhobwu9upDQcb5vAwp5Z
zg/KACikuVF7DsRJvMreLGaS2es5zgX+ZuDKdQ2A+XFHWOldvy9j+LcSadxyQOsEcT7TO+204W+4
MQRHs1ziPEoudn8gL6SukRgLB41UcrMDQcceEVYYnHYTHBEO8Md607DQOkfe6hwc8V+Vu+xW8a8d
QPmxWXWWH1Lb3oK2MQ27XNmerUI6U3gc19oS6QIVmGKqydMM1fORYhvXDFoMWm9zbraYIBl1QJWv
3KhSR5z8VX0UWAhy6r27ZnAyZNoEipbUeuymx2fWClzYzXe8RzOa23G9P9TI9JwDKMlVypU4MDzq
uYWhaxqpPkIMf25GTfIsTNiJ3ihiHmQ0JBTry5+CGjpPn0/HHLlJX2cfdMql8BA2kzu9LWz6qe2p
ih3WtKzqmOaam31yo9XOzf3hYA1K86TEYh0Nn3TRglmhfu5DBut0atv7XVyeRZFdKrwIEHLusLxH
tFoFlrrK/3Mvl98D75ySEMFT7Ol7AfU2opZ8nOCdyrJ6CRoHVMycQLZ1i5b+7oG9AnyAhpKNP0sa
r0OslXQd0HycxgXyL67OcwROehDMVLmanXfILCrYEyPL3eCcqR+NKjBWK1hi1hrm8uRE6wbIXAxz
TyZ0tfOdMIy15VOQpzDawj6qE6U7+IzG0qHyX6aDnvQY5quTwFcdIn1ovxY4GQXsPbvlcYhEcbuf
kzoG7s53voaYw5Pwga1Pq+aU3ujpf3pL06+VbSG3i//HrE5kGKnfmReY/9X329i5MT8NlsKdTJ60
ayQ6TU0agsLlP6Uu5axNmEHBWZfD0DsesutCZ0v2zNAvm4cy2XrZiOjEWScecusiRLjfY/AfKxlH
f876rkZ/y7xXRrqxZ0MWxPBIs0GSWV1VEOSGrYthO/DAPXLMUkr7VYA9HX4wpj6E543WNlqcYJQ3
ZW4RG0g+fbhJCieRO6yeDBuA66lZeEzhnTL1eDp9mVh2aGR9SxqOBCtyUZOQ09sZdIaDUpQP+eoM
cc2B3aoCkzPkDg1pSqraSSCAFMbOc6Vd8aM2RBIXD+o9us3mtV/7TaT6454xS3H9QhVc/N9S1FuZ
BvGzKCb3zsUuTQhFMIFQHhl2+joqqaqzaBCaC0PvuzaqFB8ItWVbi+EwuVrykcisrG29DWa9pAHp
S7YKxmskGiDfhUZiD53WA7XxlIRM5i0/zawFMHj+o/PQgO7vrflPBMoVvRkmJmjQL14J7x2z/USt
uFBmoLPZ6DVmkuqVYyK2uTWHoM9nE9ps+A/REUnGrVWcBN9TSN2g0mgK4ihOnKy7s9NzXLleMkhf
6S1e9KVu1FR+P8NPCw14NFQmSvdl6F3U2kKMks8XekeQzH8GWCd1+MUbb6ps7ekXudiWJvEu6bUr
s9mOvvlXXJT1YMIjHBEWpLMXri9qDpPi0kiEY4wIFaUL98DwX08zAeHXnpssp3uxFARw+M10wm1w
4AY/3oqYR6nc9pdDTrf5edQQ+yHxphLFeuXMZ857ZCdH94YQTYNYo+1zs1lCoh2UtQ290AFs6aGd
ghlMOhjuhhZmNL11VlXJi2gQzOlrvPgBUke33KuLMcGq7Gh4mBh0hJbqvNQgQUG2UZylO+mrUm7M
VhiCAsHVrjZfGgxePHDeb/9+M5+9prgQISeCbc64+bgZondf1o0wtoTCwnEZUB+YUuQOkprYC+Nv
xXswpvAmcwUyD4RsP4BeqBJBydW1gISXTP4x3x2GHIR3wXHuvCvrDiZWoRGyPMpkLub22+dklb1G
+lzukxWhAib+BHP3+haws9hR9vAisbtjesrYkdIoDxKUPkAdmcXWH7JNhimB07eDqHak++kS3Fjf
afvnIzrB5bcutVQC44uvY0w61ZvTDx+zXyRRfFif1kS6WHp4voSeunA8oCHtZ9h5fEBVK1nRdDj/
CMScfy59w2qg/qE3J2NZa0pYFjYixU65onhWVkQTCMr+6eRCa1BbqeRggMH1A34zarjoc+HjoGbz
8PAUaW9dB3qBtN86Xy+ew3o1wxzAGrq4C+FY6Vefum227NmvL5kBezAk9q39ayv6krLDCAQv0rWU
tWlhKDrE6Ze3nt/unUOBLrsBwQlgq0MdMT29KoUrcqjiz3kQDlJ64yhNlHJ9lcN8WHYk+QTEPWqv
M9mQi8CTbQ1VpoAX/uzM6SWNttnOo3DvTLHdjWtn5s3VANc6sKFFin1IsylWUCKkPr+Elx8mA3e0
3vZF59o0/jrJNmlpYCqxD2MwWLIYIAifo2f4re21mFk6D32aQgkJk9T+9CqEaPJPPmCQRV40inTt
jfMCDN/GQiv0l9RheoZ6Ae0JqSigcB+UmJlFE8SYx89wtKeWnl6LJixuUkCfGFydNsweG/EWUKHB
7072Y3XupkAf5MqF9MbWJKJstXVvZc3WSh9jn7iBwQVAwrEdXG09LGP4cwB9WF24zlc848FQSuXK
1ezpC+FbjWYhIEKwS4vOtGAIiBZ5lnn3E2C9FeghKvviT89Zf9nR2ecmNkE0Jt2j3ynvw0MP0SWQ
kT9yZEW99rqzs6Nwqsxb2qZrm2GIWabQIrw9YnRBQDKIFAlgc2aXCWEnFb+TIx9o9yA5c831rWVZ
3UAEE6sizcrdaTyHRxWS/9vXcO26y86MrGt04sniQNuSTV9PXKjxOLCIvpH7Dp7yLgaOzUwWoltQ
HMleNpAq99V1k9cFOxiYQZmyRJ0wEiQ+ycuDRl5PHrLPZU3G+PstqJrhaGeb99ionKdBLJOdg3pZ
KAy5j/UXRO2zem0aKu7WLplQ8/XLjGpUb7uUa7V54iw5bPb3MwQGRy/MTvQryp0YKgAVDheVY7ch
SwrBJhgRChf/Vo4KevsOWHabi5Xel4tCPAoYjgVxdMBobqI6KvBxf/RHf6QkkIjHepfSW2Dp3q2y
N1NS4Lv/nzDIYfAp9pu/PKyNys5AQvF6/quGGU8gZC5+Z9ekKxp06rxWrZLvPKusP5DINdusd62t
NbHZXz/b/yHPLQEmzL5QgnlM1rTgmvf0ccEye8C0bWOnOzElkRX4612PzYM5oqeWzoFfRhhNfwun
7DvzAXV7ru7OoHNocY6VQmgiQs41Hq5rJpj8oGffH2Ga1KWlDjKHmNqik0kEjKFEn/CC42zPTtaz
TiKqVB1uDDYXRP1ABmlqZwFca3mOf1Z6kfOvKLwnV9Rsmv7AwJ5z6ipIUorKVDOzUkI3+NJGuC05
a4WQe6BIR2RqDrwRjhACgCWcDoPrw7qVnA8HBvZWfFr99kmbxe+zerT9A4JGv8egG9X81fCL6/Kf
JHesmwGLIQ3odC3wgExXIkQs/Jzsi6SQJxdgvV2xfWqnAyGx1NUymVZ+Wi51RuaQrjGK4Ikd5Am1
b3+jHAy6Una1dE7VumeQKObUlwUlkAM/gItGdcEbKsjzgkA45vSvNBT8dZYJCzs7rSStKMBLEVtw
EkaSW0uvL+59qPPk0qYaGe3V0BZA3HJrQvA9sCrMWcZJXZ5Q1lFI8GCKZ708q61aACdu7qNoUfGi
9Eb+968b1tYhyk3NJftXzkcV96hnVfLi3klYR8iW9/2uPIYLFHbody99D+fX9l/FcWyk0EFxji72
Tl2BTMJqwQp2t9Woa9H0JlkMph+QTbVqSbx/KbvxEelIbggU1O9HkEnsDbVFrTtPoH3D/V9rnwFF
uUAA+TexedDIkyX9Tz+IkrI6nKgm8/BIkM2UldUDlfIfN5ZkWf0MKpeP5F0Qlwhwd5Rj8J5Zss6P
zkKQR1tjljnB2hIp7noZsr7O6EYjbayQJOhZEtCTWQDmKEQOOuwyBKOfe2BzMbiI3z+SRF3sjKf2
xbypgElw0Uby15qFB6GT58MI1ml8vPZgWshekRtkpqSnJ0U8oVAHlfnmwJ+o/XLDBpQtwUSNvgq+
qjXCrHv53SPLszsJsp3q9n41sG8ZmyictwNHwzA1V3YUcdyaiuzd/Xi5VPTTW+WJ6Xgub6qoFv9L
1hbHBv2QEke4xhDieO4rZcuA3XV74qw/mtfdhRXEaXJUkbGGtYCXG2fd5r6bhhg5Wvwthh7LS9QZ
RY4TSov6C85zJT/KFd9yzIXl0x1XJe1QlujDlX3422/p9Ql/dloeJfSt7u/78Jfcjm7XsncXBzK1
v+C8U7bX6b3/0Ckth2t2WRANkuP0ZNawQG1i1mf7+ia6dWHOVM2ErkqKdaO77iSoZU9hQYmvzu+A
494HydwU0cDaA5BaDjXJMtgQ0j5xtkwxOo78QT4YU1KJ6UTmm2QsxOj5BeUDsY1av515oclPUn7G
In6GXYvBhvhYD8KKT/kIsq8LL34Agu1z5vIoEOjPTe5T+iZdZSzWIthIhMD3z7CmiEFQlQgXd94x
8y4bYhFGsRFKpnFVZYSv7quZZxZWTqthPQEO9GQoBDVoRYZXf8J0m1qHFX5wSFGktf4IhpQMWsiu
2vkx//5VSJSNBSQtbCxJ0nXSNW2T4h5KXdRJar36azarOrk/wHzLKwM5mEwEKnl7DTrM60YV0zlo
4D05YmdlflaEjM9xt+31Ns7r3DrgCA4jfn/9khXrjgtyhNFRANnRlTOFiBARfOCMTSZ59bz6pIZK
J1abIzwuUDRtrU/ORVdi1Hwfs083TQcLzEUQFWeC3VT7RbRDl7o/NPEXeztzMjEN+1d7tRuhbSfM
DeggQWak2PB9u9BAUNzKkmX6fD1THhm+hYaHf3Xfmbov9XqFwPSGzr7KoODdhNJ5ljYmXSf044NE
4LpHQ9MJBWG1oMHNvz245QvnRlR/OoXjG+wt5YeG2+oqLnNc0Sh7qfyUAqsbIcQPOxemamuCWvMC
7DSlSGyJPw4XSYm2S5EdqUmwIznkxYDuCoOhDJ+i1hk153kj7M0HbZWGOPWJhYeOS9HxStD6CVqA
8KpUoU/NNmEeNRQl6c9M0mZhzE+uLVFiyk+WGXIY440yjOMc5/n/mNEPWio98aogSd0oYAeYRiMw
VcbHbzbkiq5aJzxcu5vUOGnKVqH+k6pVraQOoxDaz7w0lpPsbeylTsKcGEV3+3bOA2GR+0gUsLDv
nNLDbs8AdJQs4fkKVrUtOIVS4HIFb+CZwZ5HdZeHeD+VE10PcCvKSeIKn/jjm4njjcJqpXEWxKkE
kZdfuUpRmZiGIC1PrKyCpyoTrI9/jI5JM947+awTCHTvmPQWN96SqHxsz2ZmDg7ozpQY7byFbhWy
XVBYYIPC0dIe79hEqUHkXt8SGrlHg26bS2Hf6fb5Vgj7S487+n1/IJFbgYB0Zqd/O3fEQnx8D8oI
CibD/5NQK3Gp3EM89Cx707DGmtGaKgn9CzeOaViflpDiLk/voNpjXEbwaFwwIwpwJZeIaq8AzToB
vNfSxCNT2F1rb76qaORPFxNvi1XSvSpfvr6n43QkZA0CVwpayBDW2a6JI8adCP/6qoOS9/PZyfWm
UqjS4rJ5NVjRG/sb4p7w94XzzxD5ncQRKJc10XPtxf0MbKo3FrKqpSJBsw2TdzDnWdW3m4S66OA2
TsrDJt73SJ7icVceQE+UEbJ9RIy2qbvFLNdvduhQNvee4wRn97jZiEev0T3RcOIgwz6sue+IKOnO
N+U3/hbysb6/RwSoedwMyi8x7e33Fn836OZMjnDieJ1M8e1nB1Igaqy8gCwidwFjvOHZNucilRnZ
zgGkqHKsdgDtA9hTWGOhnk5Hieb9Uct2wBQ+iyf6j/xCwmmXwaonMsQnxvK/yLE9WkcPko2cj5Bd
MUsFPW4qMUWYpiL0oUuR5/aM6UV6/6DlvWtZF8v6f7epbrVo7ckNf0jtIXmX9NYnl/EHj4ogdro/
95+o/MX7zOtB4FwLkwvxuob93lNRIv6U04NcDKIj/cQWxgxANiq59jSyAYM9j7a4ZBIjEuWzDPDy
g7I+VpANJwt+gzLBnzBBNoX3D4uiGv09DBsHUoLAss57qMvbxOrLDx3CR7NOY+LMMO9qAq3KsDNl
QD2dFYnfLDqUMYkWlslHmoEWGQyDUI8ygNcV4vQ8CwoVVe/8izF+hOVrTZIofuA52WyP44lp4xeb
qwiKHfyDuhNAhYzuTKEiJFHGZv7XdaesbWiY5Ch+zuHoNLdt5HMhg2BGxOoYJ9FVth6mrw43GQUf
poiKjdvuHC5lNk/GLbItXD2GWm6O1s0fOVQ1ztwD4OwHxItm7ubOjh3392Vh+99FFUG3L8DpoZNX
Cp9+OCET2/G+fiXfmT6E+ulG5+UaAn4t6qTK0CJSWmrBjyDLnSs1kJesiJ7yG4YGtIh/rxPmqsGI
KybiVmMjIrwInbrcT51DHG4yyyY0z6VZEbvF0h9Gy3sT6TxNwppxt1Z1p7iajnyX7t6X6B3YWCf8
NVJTdpKQF9NhqtyBgXhMj1ri1Iuks3UPdBhsYQbyJB8BDqVP7ACCPMWjr2TDP/dYLvxKowUTBlXc
+7rtYdRsOC7HjaFm25ZqpIxCCfa6b4/oanh7qMWTr8cPgol6Bc37vHBt4MW1Rd+KIpl6vbn5X4hf
0FBlrQmYzzXSrUZDPCRUw/K5Iv04NMiZuZyhfx1HZ8wuxSgYmxDWhP6R/ZmdyrLasG5dOwfvC6pD
1cx5YLMlfEEiQlbWpikdTFNAXpfWXpCrD0IgCTtDVyv9NvSOfN9BytQebwN+avdm1M7NSuBZYTSj
qj5D849TAHhP7TfH1797DJesRlnHSCUpyazUsYijWflmLLRyCt91o41dvZckn6d2P3YgCafxc/Sj
9SEnZAQ2SsJEg45HNUgyJyQ5JNFfeVJ7beLNsBondkz0KljdxnCfKEkkIPHUO4cfQ3V93Ny1UK5l
YoXRDV1+Ka3jH/Bfgf81veuB+DOeKSJxNIhAtQ594sfdWkk32MZoceHfc1iR2JoEzw6zN1oCho8f
CS4Ic8CTj/wf0cXS4kYC0TJqt7EEplSDjkzcjlHynjblRrjtp8W2G9cC8tw/kDgsqOhjB83NZQGT
9NHHAtDRVFbUan3os+o7BJbw8ZSW2nZPkuIq/WM1/zi5mAMfT4yPiTEyXt9DbMSE6ymhrrLUp9kZ
bZ2w79G/oZoAOTBOBBw4J7RRsM/V4dGMtKdliExFSVZYzr+jkYd4gHnflyyWYfUSyrL6AYzB4q5x
AnlAlMKi2dJVDhRbP4z9y0tK++SiaphzOYxIMBE7ILgHs175oML9If7l200xu9wCKDP4XhdV0Uik
g3IMK8VQJuT2WyyO0cv6dmvws5sGrlI6iPv/1N3Z4P99Yt+2kYMeeHBvchqT7x0Psu84fvInVBow
j4ggRkDEnSGRRljh6VAnUrvilMIc8FqrTs0icYnGuwS89xp6GJCgyRMPQ1HcWqgiFTMsrDtFUjUI
VmmBL2sRdFJxMYhqlhi5QGhtcuBeNAn+oyqouljP0kEBkXx+BuvRvKSBP+qG5a00/pPjaWc6p3E7
I05L0/hnxztZMXkK7iti0YenQVmcX4/WmgPcZORxw0zNGQpZjA6zI6aoh2fFk4U+nCW9h556+NOe
jlW/PPNTy70RdnmAaDKt7v3DPtSEUdwW4ZDtlQpq1FpHlQrWMk/eeDQ3g5J/uYdc3pRa4mXmHFgB
qMcrsawNwpGkes6XRiBYglKvgtI8zR7I2XK0btviA19Vv+AymSZ6sBIonCbF//d8STgvnmdWRjio
XFjf1WwQREHwozcHqmjEOxAIeuFE/uPtaZ+7U8ylHiBFhEQtrbmxhkItQ5gqKvomErGjWBlQ8HtM
D/o2tSqf2PbhfJtu7ovVO76hqcdEoRuYUuhYvqa9MpeKiDHErr4B65eT2fM3O5XsQOIH6gHs+i5o
SLpznqaxJ/G8CUAChVxyz7V3iFiZIzB6S8NSQ1sdOXvA/UURRlPNwH+wxG002oOzg/Wavm1dxY66
A3KXHnavaP00WSMm0CAa2a9Y3AFzhu6a9RIA+qwk3ArmfayjEAWp2U8/YAnH+vkCCdSSD0N98cul
3HveOPU8RgijxFD7WXMPNxiJHW+fdnuwmxKpvd1B1xW3miBo+zw4DO308D2Xi6oEDCzidDLB485P
z2By8BWQhtDzGritjdq5qGu54pQWsXWGK4y5sLXjx92noIHNrTajaWVpW87lTtW7yuvsYfPkK9u5
93NYOVasYnThRzN0LK+lCIso5uSWe2lxx4esuaN3J7pHqWjON2l5SiPL+AwTpu6Vo7lG/5SQ59aR
KWOzie5sf2SccIWiQ5l/Frce9CBevc4Ra9XL8UE8tbC8leMle5SYgtjzJYUP0wO9IxGs03Q3Alo6
DJBSEMGaYaL0BlYsrmteuydeZK2MNcgFNqI9adSsr8GkhenE1WbWmSTqq6KoTgsEGYFrUyYPRNGs
gpEJ+SpOtOQVzJ/0jq6tw46g8zQRqIzfEIf9VklnWQhorcujIYT1w7t7ev+2DuFzCJcHd+geB11L
MagtI6m3tLG3ELyDDBkBUJq29Jq/pEAuwHkD9zTzVsUSyKWATuKQddQ8WaTuw0qnKT1d8aXYY9A+
40ARaHILTBFa8oR2XSci1//4SQ3IpK31MVNIHSbp61NvxuC3tqxBhdciY+a18eT5UIw9S0MEVJgJ
ayNx5S8MYBC4hvqCYeC+AdHVtULaCZUySO/z68AiHEKQ2hn4eeKlM39heNSTe7pZwsqlW6ejCHDh
h6Wic15x6lfWJF9LlsQbMIBpFLuaiTOsIjmyZM9NPsDMge350EZ+2RXVba/WTzSBI07UD+NDxXi4
1tZq0MwVum48ovz2aKZV5KVLwrqvWBdVXMYXjhgxOGrzXz7U2NTQMErExoWOHa9WDR1eSHx02+sn
F+tUhrVYKr7NLBY8h26QSiRDjnhZvV+/oQYP0PY/zuZkAnaZgfVbH2NbULq+85S1OdKDm3cEi4xK
qfOpz/pLeudkzfZG82QJ/tYoIZzANJ9Vg/vsHEbB2BfN6hd9kfrCIxMVWsGyKSJAgR6eW5an3fUx
utYKbuVC6W0+pyRIYCKyzuzTSvewo9re6T7Mli9eDlubFlo9IBgUw6NXXXeqrH8110nexqt0QRf5
x7rc51g1y8vXXBy8kvL3TXJTsHjIidVMA0nXaF9ZarAd/+L9h33e7dbyrV2rNSGkJTueCvkxgh3S
5lg/mJJMfh4zUm0Y0mMpVNqXQyO38VuO7pag8zPRP8zrm9wbw2ARIor5Vp92K1sYpqEP5YPF0hZ+
ILvQfLq06PBjJ0CU6TxrYEUQ2ZyTIxDKHQIYu7ycuuhbd9XCGPZk+3sbEiKE/JWdqdCwZu3yP1dW
t+ZpW/4D6MQ6fqRJig/umFAe+B7r2IPxMw3yq4H8HrifyNC6bKQzo9VEoHP79uT6penauar6XC/P
E4BbZkcSROv9Uw62qIVfwji/cgX2vaeJlWKFOZS9nveK2tMxB/qT1pCkZXkJ0THwF+If/zol5VB3
n6Ihx/Fxz3HTz4MD5nrVlyEL78O5BEnX2Ua72hAF66xbExQR8N4HK8p7nXvK1sMysSLk2xnCpeeP
G4UMxeSKPaoJOEf7qkuCeYi8uvLiSEy9Do/O+sQpcol169gXTrMpceEGsS+aZaNn2kllCOHHjb9Y
62zeth9RW4oqhmjANpqhZ3kgvq2Eo33VrI5u6Wazb7GzCDWkSPyR3ZjE1CI24INmJktqRz/BkT6a
o/FK8UuTva484NtDYJY10xXZ/N0kugBS7Nm+pFHXWKeZXLDfbvXOC1boEa4HV0hgekWtVaIRJ93R
l8J2JAktHO0tzAXrtv90A7Fhpe/XffIRhOvGYcAhoz7+udmHJ7n1AwjmfE9ktjNUjjDAcfvbiblg
6et8nbxMkpux3PQX3O3YebcTk3cwAEoxenS/Zf01RMlgRAmAR+A9CGuq1XDDc4v0M5ZUYSivGpfk
bxonLZv63K0fZ04wVYLHD2OQgB6e5KaMII7wibG+qh/hmRvJy26FK+ZSY64UZ4fyBuSKvjSsp0o/
lEPZdq0EFk5WT5wQLL2wt2AxHmJmCnh0N0bfbM9HBB/B5BSA9hlgjE2qC3ykNZWtNGG5xBSCVb8h
l0zJLPt4DhXep6RxI1MDwtdGB89TOqX+OBciUqeT1hbiUMldlWw5LaidnydIXqhdNMeBMKWoW3zt
1FgI5dYZwDuQXOFXfFNuoCBLs9IT6cj5nHoF0fqGG4R9o+G7dpsSGe7l4fCg4fpGHbR8h1by4JXJ
y72idfEMRf35S7bFa+18ToaRdyHJQXLUqE9Y5Ud8coV6rWb64rtKrhOsth8SImWC2X7N7oZ6fYaK
IiylI4a6Xky6c39X2QNoqMKnyevwiYcAyPewYON2la2kj2VqzZ1fSrRRzF6vBy2tyQMdilF1VqGZ
FKradpO1VtJs6s/GEzgyWjIz2t3wBjjX800km2T8HHcR1HgeMTwG79s8uxzhoU4bYurTiFhO4DQt
UgCrfBu2Pv66cAHYJzHf8z0PmQTz0GPa3+iZQp/+9usyeUvQ20aSgbT+DCo43ZCj0uzymR2D14D/
FWaXS3MBRw7hf7H9bTL38Pr7K1BINYY5cR7YY6BhK1Wtfd710P/p4ZrXtuZ3dWZVaGwoWSEsq+xF
eSVEW++Lq9tnUBHXbXaxxqN9w7L1oaptuLBaleVJGd2QzGWBIS71VNwZCnwRQksXz8lx3F3MV34L
6eKbMIh9wUTG7uh4DFgyYx0eyARdr988f9SxxYQXOSSUbDS5uUa0Oyt3kVYw2nEgPNyBZrPLiUc/
3708SVCvNtPd/Zg8YQ4i6gfTLEHwbSY3qd6NN0HEpLYrC3SgiCJnVHD1IMks2KhHuTV7sQa37XbY
lqSIYMJ1p7L5MXi8istkhj7IQNFZMZlHnb7Ee6ZvgUPrSj6kjml0505a5P6Cxr5k3wKo6I8jNxFw
1lqK5NiQ2+3gbgtX4U8OByvPOKzOf+8vpmHzzR3waHULON9x7DUlkUm5saQPpsLUu0HcOVnIkmvT
tTh8UatCCwgzZV34jkKzG1s6HyEot19AQBJTc/ggZSn44XSsdv8/cfprrbHl21xktpIX1t5VKfWh
JI5/nUr/RNr7MdAavq3943+Y8VyBOdr+J/uv1+sjID5qbT5mg72aj9r6EGIF0UdyAw4MPb+z1oD2
xF19dps2toX7DsADJ1MFKzoKvFvE6v7j1f2DD+vpVXdK3p2XqGGI7lwCPmExbnanH9MsMGqVQta4
sdXMP4phkhBBaDqZwC7tP6tfQlPAYL0mrLsdra2xHeIR0jrUlVi8BXE3dkyyjsIT+tmFg4CV0SHU
ZMgmvtoBLPoeE9XQS9MTYrwJEMTTJKYMewn4BeiGb/QG2YSQhrr7Y5Q0A0t6MXjH+gf09UVeSwux
gp+6kWCHE3e58s7/nplTEoSz68N+bEA6X2bOveRDlvuYaMi0euRt8c4JTqBJ+op6p0Hm6gMjqYPc
kokpUNQB6Cn3h50UCM8rZpdYaUzCBgepx9HcKCgWylwr9ZwSOM7MD+ARzdw1Ndrtfx1ftw8sKqCK
FZ7aAzRWhUDDMjLoC8EQAs31bTr92wiOlTMgFg6y2ob3ZSy7q27eDgdd/qKhw56iVMms/05UXbUV
4aC6GFZUQBq1e+LYWMXkXPHzkxtXi5n7ec+fO2EhRK4hISR7xRD/xp3th3uQVGtha+7he2OdUs4v
R1XUUZ7b/zegToyUlF6LvnWVEFLED07Sc0G8fW848qntuL5Z3S+UhYid4hw1AcD3RnIMMczuT8Vg
AEqVFhTrECa+kHTE8j77pRZMiKWShGMJt2sHqAeAkV7bKXJF+EmB6aEpJ0vkmDV6fBtMMzRs78Qz
pOvWeZR2yFp8wM+eBizc3FuIYsQ693jZteKfPrA3YE+Dfu/4v6N3drlAmsO8hh5LxIA2bgP/S2qH
qTHj0GfWxP8QJTJtXMzexJif57lfLRg3AHHn0uIhieoMjZakZu+RJCd0ayXy+9+O0OXnjdWW+vX5
jnvyIkFeAAuoIuJZAo5I8NI+CjkVBtETxnGyZyzzj/uC+4sFBejR5iPZG/RxGTD4w0JcWZ0BaWsV
lOW5I5GWBwaLc6H1RUPmIlapy+GrjKLaAXEznvzK6rtZL+YgH917rK5ctXLPTQloo7Oobo+0UZwE
HFm1LcD/5i/2QZRMMGErRuMhhFAwUn9ucpSi4iPqI3bMQvl5/G/na6jwm21hCGQHlir7vKbvV1h3
n5vsOF7OzZR6dbItY5dAEFLzCIBgVBauajLQO7jV8ae0VdiWSbRc2qxygP8yXFEbH7SDaGccvagp
PwbGqvhNSJi/TDOyGUf/OaU3PJEXetn1yp0tbthS5FvQa5jZXSKPO5p3EbhVBOee6DEF7K5LSBVW
TY0YhDEct/o4yxmmwq3Hso0RpAx3CToJadPh9aiwb/fKFSTgA/eHt9iaiaMlQIWzcfakiqbTi1b4
kNdGgxx4Z3uk0jJOx80tzKF0ndmVGcP4Ca5NcbCtcRTtXiz5xUZC8dBKwbImXMDPPS4kDUvT4EN8
/kehkG5QNNFhFMtvtlWpKmDxjnSwHgCYeomcHeSwM3PCPMZXJDeMSiXlrmowQ7fL0iVDEuEr5q5e
DW6pj0WtnOd9u2NxH9YhJ3pz3YQJHymoeYvFsxjBc0ouYN+WPkIkuTj7erN4VwAKdJS3RPvcYJ6H
54VaOCV2XojlPBZKGttiic7AU41BXGSf9W9ZJOR6jaBY3riNhPbNmnyxlOtDaJkUkcUq8dirp7N4
gwqX1UpbHRYBbyw4vIPyDGlIg/5nghBvcOP9Mr8sTI/AMuzCvVAWnra0nkvaX3zMr2dHPUFwTYnf
o88Xa2TzcWs0wLmx3kbCUSXyG2R/vaDoj/bo0jlJA68aAjjx0J2hoEuEhXnuZA1Lp8IKEqx9sOf2
3WFffEbteUnS3OZvjSHMuitH6bH1VByFRNdQJ3jfgXAW29BvHf/l6Xaf+nDM2w4HgSJ0Pg/2IWRG
7q+PA8DnzNy/k9zlXKz9haxzTLBv5/uKPwy9m+Rv5nHln4yxBkgJ//+Sj80yN+NF7/lymqm1bNDJ
VSUMOcB76jmje1qLoJ7qSQGlt06YLmnfYE+kgzTs/t49TGV6rs6dKacpXyJzjl9AIC2RVtFTCS8y
A1gWqggBTeOtILyi5LS3HNR+bCVJRZU+MI1vmhEdFEWil19aMTKNPWTuNqsWSmCmBBiyp3vz1W1Z
pFMsE4ybunlNyW9fVSqiM1LeF9vK9K6eBdx1IK+YjNupNyDEh5+cv83MVey2RuZtCYvb5L2Wu+W3
MRRywfn58pfB+B0geny5DphYkYXx5uKuWw/FIL+EPNF1328RBwXaXboH9GkdNwY+QB3ZU7wz141F
y12cPR/lRC9liKVmWwwaPTEBQX18dBz+l4lifYz54VdWH8r70FvZOdkWTutGLEcNKWHZU7LWtPTv
CADHCixL67sQTQDGBHG4onVywBk+7azypd4G1/tfdFfH5MGNYjWRCX3b+z4fV3yJwFJJDZEoWjm1
kaCglFV75M+tc97le0bV5cm9o/+/tnyIJXvuQx53Gh0DgAjxNFOdKmgL/oUHpxSsM05HBtRXuzUk
9Hy9PjGVPZC5a0eWNdqfW0EZ4upcZtMMnNkyppDaYFWB4gkIm5oYeZkD0fkdXoIhVRiS6mMKAZeE
+SDJ7Mly0n2Nmu0goGqOasI93QEuAKSFLl9YAR15Y8VPeYjMW6oD0hbH3L/dqL7TMPxPwd9uidKr
TVKOB9iwcrUF87O3dX3WAarjmROJ2H+Qozy9sDDCNpKePC+udarN94RCywr9+49AktwVeBSBr7kz
3buBI4iEXYFqoIh7WAplcZ8O3NND7z1ybD6bGXXvCSlId4sWeFdVCU4csscqB47HUR6UPAFs4i3n
QedRbx0FfZEKpzSrOIFANhlc7X9w3TBS3fe10JIuV5M7WOulrWEUJ5Hd05dcs8nFjKzAHtm4/Kzh
PG+TKPfE/3BPD1uqLw+1n02bEFDTAW3wIqeUTngPWIkv0sPEnxZK9YyXU0TO49GGbVrzQ3gH8dDU
5KmVYjCt2jjyutkE89C2OJqWOdtJK/Lcg4UMH/5ZiWZfUf295StEKD6Fdz+frcZSgtn3unqm1AFi
GnZpChOOs5TeqaXk3FNZtWkMh0YWz2dYAKnZKqK251T8iepGw4GpeYPrvWs+bhyWHXFsErqkJ4Y5
bSDk3k/ZGXd1txSn2kQxF083eMCagBq/IY7b0QNG5/bzbR6hkdTRqhw6ffNEPba2UUYceysLb+E5
rYqeS1V0w1PwbHwXP9m3n7/7kqbOru+wTwOGwGl2QW1Q9WNJE5o6XRPvbXtSBGCgQLhdiZ3gPySF
fIUI26QZSzKiQl45hWfkpmSf7VhT+3coCRGXzPkWNuPfhVswG1VW8d9CZkyFrZfZYhFU97Kcr1HB
cbOtUKk22ZHXTEYVeOH089z3jALv3Bt6ALablNrCFlNuE9ChRWQejqUIjPENa7nXw/LYgS6H6QH8
fQXzrnQdJ3dYDq9K8j9LdTl4vbyitIR0+or2vWEat5yas7e4xyQAAEIGiS3qgdNOJ4MOUmCNLl4c
VxNlvZenL8zhotdOCLe3VMIv+1/2RsubXuSKPFGpCrZhrJvhjvhfGC6dtWoDy18OCMOM//OrasBA
F/Hp3gTEUgZj+/aJB9oumSsSShpAa/hTWj50g0bieFs43wiVC1GpZqvbW1bmKMRTwSzjeIef6vd9
AwsYl/Se74lFTsRdCZFqBqpyS3qyLK8mFxAXNFPwTdQldKf3S3LhT1KSS2nAhOv2qVW6byiJis0y
7c6uVyIc3c3ABT5LfkcfA4o1jeuaanX1HYXEJ7T8bBZOEIJzIfixavuaxjeXqMu5olmxnPretbYO
R/3FOd6RXIFRPPa+qGz3Sa2+hzY1IVwzx8J9ekAIbVJfUB0whZrg98U3rVz1qLhuMr4uN9dooKH0
uuQytBcx5qa2xTaOnxLUOV+fRSw0set7EglOJB5HY7sJEQojBwwVmRJmWLvv/zw3rabYQOtdZVrJ
8ixuFlCH4zHWmppoLm/XFjlMQbMBU7zdXMrykW717dVggYX4PJ1YcfSLyy7bbJoCuVfSffG6QzaL
Ro1lAs3jt5KqT8mWYhN5dYNADR7SDsHqSQAsX/SNoDpizuZE1KsL2jwDW5SSu0kbw5zx0XI0fEgC
MliYJ/EHXO9hHLth0g16JsSgReixC/vd9yUDvjIKTgFhGKB0vzcBKDDFTmj3Z3wV5bxZjqH9B1V3
nhWvy5wHwy5fmzE8Dyfklj/MDzzRGS70IZwS4VF+mqexEn6h1zR47EV/zkg7AGoIRKPFmMGwMTGU
YohwosTNJlKQbd0RMdMgZmtIvpvwn93eesidEFD8kHtLYDZnAex3JNH51vovBrymdlVMV9IF28aS
Umx575fPfHNxwph6LfWN2LKKql2xppZQtciyX/ASinn8Gnkztc11k8tqxL2Y0YcPZicyWXO8L6H4
HuhpeRhGVAOi1DPhza6a9lGgqDT8lvO0/kKPN2UvAlWlM/TrZNxX5fHz+Vea69FNqfr2tyI+/ONa
DJZiWA/599VI69FePRhZlAU4qUJT3WVtlEronIMqlrYlrnpjPHIVAybT+wIhUEIQW3kIcPBxTmCa
UeoOOiz3wGcOGTJcvGJNvqb6PX7UBWwmerCiiUZznKm4Wj7X72NDI9EaibkNPfRswQIsTBImLicv
XUKDqjfyz8JV1//o9GUXcRHZbiVbWJN/KxdReMNs5H+haj9l2pR8/yz03Iz2BdcF6oEHpxT9wFBd
nyeKdxIC5BWvLao4qtGQZGvVS0Rru33eb7rfh0MUEOSPNwzDSBGn1UwrmQvqYQflTE9l+NxG0iOl
AXRCriQu4VdKOhTwbSq7ZkqxvFRG+6VDO7XIELqIeepcwiggaSvRBVR2y20vVXyKkzRCf7kMkbaa
tnJs0rX9vRiQA/KWUBxRvfenL3+FJiBGpQNOeU0Hy1XPYerlEoJvWAejzYvb1TLsbqSkKdq8qJZg
vpSb5qAEmlztffg1ibfgbw+AMXw2/zkISxcF1ZM5+2EOL2tZx08Of9Fj1XkGjOxyxMhfHeLXDWXA
Qv1sjNQGcv2Gu3TNPuB2mjkVh3JvabXk5k4RfJKwOfQLJ6wrc7fk7DiWLmPtI4vipkPqO0bMYDt5
eEY/1RcMKpnMMyeYeBBUMoTAurahP9+cCNvPGrUn4fSHvdmaBdrDzolz/Shs3eb0fPgfQhFkUfuc
s89Dmhy7lK0rAB2Tl6ZjDplXfryX4Kqf5ZGniAj5PH/qSrIG0U93SZh6RaXh5e59CXOpaU9ClzUv
VJVRFPODtWTdX+IuIzUIKdk+aEeOnFX2idvV+IeVBvQ24UDng8lxf81qvzZXaO1rRPvRCy6LJJwf
QO9vr2hPMHz34KeXYTV18y3K9niNSuk83OePbGb7951+lSydv1saYDgyNYsqhp8G8R06di3LcNHT
oES1n/VnG8xF4g0gmATGNSzm1jfIuGw4Ea5aouxxq2Nm5zHHdQOwKO/qtVQQUPzFhFShutvZi4Zf
Ik8rdxR6l1NxaH+duIPxbDLKWubSewpleyhBCQLKBE+Mz0onyaFly3fUH5CxeXCAX9ekpng+vjIW
M/I74xa1hgYbAocgHm9OFcFrtCMYxQ2QEUROwqQBscKxY4voTlcCI7sVoKWExCOHBxtFSvMiJvzp
Fgbvvxg5BdCZQAshSPts0Z8RKrLMI2XexKS4rVen/RPOXEGmjUJtvSOvFLV8fT5DFusSF/rPidil
45hFvut5PqL/4PA1yV9xetVpY+lLxZz6Qzya1EY3pHV2REjqP6YzTu4pXLPkxWpYINjDVlEtkDpU
5/T40qefyHci89ds5TRzcjU4UVbL4ehkL0kaCuvTbZCRHSed+2n9ofpBBNNsulVwS3jhdBMGIq0T
tUn0d6zHQ4zsEDqry4bl3qXlXBs+sCf3pdeScAcfYd16xphCTHesYH1vYIrNiBBRNTOC24yyjpkc
NAvxiyBXMgXEj/Rk0YD1Vx1LDmqQhlL+zgsZo2SFQBPthSb0Hkwtq5AHN/OyeNhm2/nPMO3BigwE
WiBgtBTJSNEUaeXkJ5gQVd5C1CeI4B7QbqR+iBoW5TfSk+KGea0Cim20hGrekedppCLO+dSOXDCS
gsDUGSVaqRslAy38RvyO/gvuvwFK1+MPxLeQiNbUJpEW7gm7NzWawEGXeflVrK0Ib8yfcomSML2a
7CqLl3mmx7mHLbjjlvoWgRkvVJeMqm82UAkGQnSaBxuV9kh4MO+m8tBt2qDX7GdIIoHR4QC+sYHz
nJAMWHrO9+mjV/9MJLGGDb0/K1VwOHPYewjqE+LOl6BxkP4dnFqBvnXXkWDx70KeeGj+04lLEmV+
YJJnf7Z8uO0KWEmxduzUzWwPHOvCf2+K3dw262XwxfTnY8PaesQX9SqDNc7RV5W3q/aBy+7SDsD8
ZZk4A7DQ9fa/Mr/7VJch0bOLmjvexPoN8KZh6Qy18rXdyGIPUlTxNuMTxyLt41HaDMjSNl5ZjimR
7xr2l7kDcrXIH2g1s5YNoZ3nbM0R+k9xAMDaEKtH/viH93R/SO+1d1XGyL8WtA4V1apYBH48IKJ5
OJUeUNwxhxBaBisYNMtS737INhfT2EdpsWJk2kJLx8I80vuYP5TFQG9zpcwU1PJzviOoA/yNdX1C
0TcQZ/IJcZkDXa/iBFpVnewSxhwrRLF+mhG89jNconttI9Lgnver0yAhCJwBAXiDrNE4cz0Gflba
35RnlF2UHMduQtw7FyYFChyy9tEcDIeQJ/DfGDzj43tVffHT5JjAYckKOcNzp4XkhsPW8+9yC/Px
uBvZhBctnNAyJnNgMqFtPXmBrDQpu76jS8aOz0tUZif9AWWNmIl1VOA4BPZ0EUSaSVJcaIQEKNhE
A5SQx15EtgZih1kO7Y3EYRY4aP2zfOixosz1ymaEiSM0t1mIIuZvrbTULwFEyLyb86G+ypgCGc8i
s9/f64taReFGyZv4rmegcDju9jGznKbohw8B5W0qU+C/KqUaw1ycguACFHcFTk10I37wRL+ah3IB
dVzfTr6nAtk0wWGO6urbTxSAcppjuzJahmj0VgMwaGxGV7PsuGfLk0AZ8GlkqrpJ2QbeblCW9jLz
vWlvUy+1p3SqeKXcH0XS1TBOCRxOcA3iJyE4ZVrJv760d2OAJ1EIT/JMd4eyFa9gmQZ5nNmSAaDR
GPvLL+i/WVPJda78v3xf3vdt+1uOLHZQalwrxdacA9gULUdmMRYjzEysJS64wIzSA9369u/EuZBA
8PrNwFVmStgEs9KDCECbQqOe09x0k9bU8LaqBPd8VmFAFWZiylUX8BiarFMUR1+SaDoZtItHCX3H
9b2eNcG0P2kujCeGNWDEv9r4Pz41G04SmrEFlIEtYNtkhZffuyJTqDi6lv4XEUnFynU92/F2D4L3
YQIbVu0AUIqu7WlAQwqUVVWAfNYCJUBVO2lJsFiNE5cR9DC7ArhlyXwqnbkpFJf3SVgUI6GBm4IL
ynwP0yQBZa/aPEslMAaKmdQkYK8D4Y8ubfc2hPGzXhKIfJUIS1+YhSW1aZU0yFhMoxUVqEz5e13B
IcH1ATNRUW3zdupF14Urve/xkLVlAJDzmPYK9eL4/fsVj3ulymmwE1xSxOjPNssKSh/A5/Wc/2G3
wt8X7kjmEwTkJ+rzcCPDj5lWmKnn/dlTv/xlPmFNCfjJOrRKK2ONJ/Hdane4LfRWsZDRs5Psq8J0
Ms7k4UeXEXxqztpvhSt+XfY/Nf99w2NTghlu+rVsF9inFtQSg15/jcR6rEpHzqpc0bk86Htk+wxr
M/8nGtr1Nux+wuoGIk3gEg2W+ozkYnklGoBDGievf1UUtxVKAPv/n9nonJ1h2A+Vo1tFwSLk/9Xm
iqg1OR1VXSfGUaenMcx2d6vltC3li8m6kFVYB/JXU9hxuzp6LcayS8p0Dy2ldLnirJ1VKvwEdssw
o0gQUOrZWf+vXNeNFNIm1mRuJiwfICxqxSQzHBg6k1bUCYQ2b8y5zOsoMZy5MO+7DYKLgoedI1Rd
ssmwbQ6HNTIYHXU5TSdLInTvCnoYVhN2Wtu29bfAF/v5O+KfoR6v9MpWb3SgEp0fbWqqRSei5I8/
lqYviTb9PAnUbH4nmj7Qq30/+eu/kR89phADtRqxcNFD6UYpFD5VKCMWzpLoW2DrYRqtPTsBpkDc
nRCjD6VI74ALfkBHhDY5IsUuVkEBlPRg92eUamIlEx8eFqGwbYIBnn5pxbD96fpkc5fX+RVxaa/Z
AU9ZLbNudrosOzy09eJi7xsJf9nEs/+VQh+R31PrINY6ouhUrOZzpQEc9wVVOkF6qGECQGyseLhX
RJiSSRHpdtEbJZpmQuEIzv0W5zLayLKfOaM/ZZ8Yn7RhHL/A7NzQH1RHygMzU0dtmzXPL3Hb8uMT
CMMsIvXTpBdi+orgolExgKeNOSQf6WVNMSHYHq7zVkqKjVbKOzOH/o+lMqEJqg1d5FCslJ8dEAEv
veRqhdv7bYOSqWlSTClixt9dAh06Nj3BlK6iZjx5daeuDv3BrOtmYyMu2W92Zkr5HvwdeBmZ2Kjd
gv9glwR+13rxNvAtM2m25C6hZC+LGGh9B3kWCrg7EoxBLXEdF16HTEO/rNh7Ng+Ly83olg3u+9Bm
lqD2K8pKWXRK62EPeLoAef53KGVkRWBaHMPwHCxe9f0/fj6zu+H3uctjB8kFKk+SfB//d7QGUS5X
9n9YknqXZo0/AmRxH782oVr379J0keIBbpFPn22bscttJnxhNiax8jDIaWrf+AIbOprq7a25xWie
oHBMMjvJVyM/s/G4gpW9cv2MDYx1xlhvZiE8a7i12w9HSUKeUV+mU9EZ0BonH6TNdAF9bm5bYJ8z
fcQap1oZ+o0oetw27rXH37UMxWCMts83KAEBhhH+BQXHsYFHHWfHYEYqG4pT7It0oNutyaQ2mMLB
2bwUOoDs6ZFAHpquSVffCc01l9EyWN2tlVG8qv4TO6kmDTXZncPhA4ZaS3eAuwwz3Xm9qdR1Drb6
DLIVmoNdtw+hZVVlegnjm4Ix+1QgLD201bZ04ht97KNxyAvZha82JJVBgPRrJYYoQcj0HrhN+MQr
1qLe4uHbAgdWh+k8koa1+F+52AMPQc915zK1jpk9oqji/6sBpggKZuRCNX9pq/Pi09xmiTy6hool
usMB1pjWPWUbEklorHkAGN72jc6B/YitR0PX63w6MLz3Gk2zQKgVdsHeFZLD9EpY21b/DUHxLbdf
78+cwielbYlE3KYaGROJX2cBVNelb17ZI8uySKB2XXHas4gicqoVREL2HZI5gAUFc3yj44iXXTrL
so1eEdqLWBmSaptuDKODRcwwPluOOgcyn1cSNEOh6MsfX9UYmbdnlOizJfel0ArvancWR82Uv+Zn
Wsxge42WhybxyAQWr15k3I0RNCsW2Pz4alyDpKVkyOkOZ9ydWheo4M5rBURGWbhGsD25KhfDRKL8
9NXcAauXDmoUS4erbvxIdYpNNFHEPfi3+s2nAo2L3BnzkoudXgu+nlYOnrQ+NUw6WYWCE0CXFzeC
1orPQwM+ZmZu2bHg92WUcyCPPXiWqFVxb/nYCVTM1U4DW5YRpF1k9cbF97XaP/HwWk5coDHDhxfT
DTF3vygwk3zWE6lgY/d8WcreGU3zd2KfgKCCw239MubAR0MvtRySvtvhZBEdi3Lq20msoTbqwfgJ
X5JQZ53A3YKJin6CNbnUSETltW80UHLO9bCFtnPrd5fRIEUpPgoVS0PEEiZU/ozv0n4tnIAw88Xb
UT6lbqGx4bGLpc+E63J0UB4TX1tWq9T+uA58xK9uB5Y0qAWJ/RM8QaHs8IQx68HbfxDZrLt9C8fr
P0mlzN2RNbaBs39bj2jH4/mah2OraGJUIydVuC0fER2RFTYPXfnJ4uk5ybCZ+LvZdbi2n2leOqc7
N/3U+JtkG+wttVR0nKmvu+Er8nzFBiPPCkhYZx3qxZEHtw+KfKBKsl0p1c2x7PyU2NCzl76PYMZV
ckuA5Qg4fUIbrLygo7+XxrI4P4Vcbe7g39sD2lfICkjZ3X5kNEWIeD0XIQoi1bRzmcghV5xuyrKx
m7IyXfZ0UBJmKhNJYYb9Q2naiIMh88GDDyLzL4YGowe9NyPffRKVHGRT2mlcqv00KPc/XsFYsoH9
CmobIiqVMJZu4u+9qfY6tKOs6B6fW9ZOU57W5dfK3I2qAKLZ4exme1IisWYgDacoZDTrOdEY8RB8
ARzlln1ZOVShm7WE0GTsNL1OIzdlUAu5/P/uUVmz6SjwRBtypmrv3U/bfrglSrpntKerAajpFrxL
dqHMF8gDX2QJZssc/Rm1CGN7TlGh0wksxw7InJ+/9ZADny4Jsu5IAOe+IkBZ6R6yc4tjwFbaqYQk
cEoQO92PXxAccHcYkzOkWXAeXSYZincdf7kCCoz2i/Q+hFvLAsHq88Hl0VgWc9Ah9ASxcFo7CuaW
PCF55wXWcPASYMXZcXYN3WQPFpLSIDz2FYlvPRZ0y52FCgNTPqlYXpyYX9kx+enSIZ4ML/ABvnHq
vuf9zkfKFiLI2qV5dtvNrZl8tKoQeZqBl0frUtuYLtkrdW6G34l4i+QwaWJVO1Qt7WVv1YB7LzMA
jauJY4ndYQi8G3VCTsbbX6xs2x7cqjdBOeNgUWKFvsGKpIhUr6EE++rLeYdsmGmsS5CO6lSwTi1l
iTuVDVJVTXCayWoL5jMUntWuCX8tSafSAFkSEV5wXS665fxyFm+UQOLLZg1jhoIn/hx4/NmC6dx5
Rms0m8XknO6xRuGA3eBWn/K3FUIPQbfFenon4YLkHrslmLrnrWKlzd/sfon2RqnBUAbaotOYVuA7
xozobIZmJgkArTdLQqtabOOWH5OGmKDAFfJdj0PcPCgivklNoApl3/txZvrKQ1FCNQqqjp3DJj16
LmppGsxsm4thZ/lswEa0iwlC5kviLL9yRhuEYjMMrrwEhG7Ri4hjT0NZOSda2moDITI9noapHILh
aq6WqwAeHKMlQRCYuvpOYn24IuykddSnMet7EcNuhaiGJUA1w9DjCeeS5OKorCNgopTQYyBFXR0L
9JILHO8CboYf2S2HXjpQn57nCOGCKIRVe8bWLgV01Eq/XUIUt9TFhRWB2vhzPWJQs4ujblO4E+Oi
8q8G/Uc036XfZzslkl82qVdHkyhGCnQWhH4sRMrhKgVrmdjIg4Jrn7wp5zpGI1sEYPMfIo/1dpus
Aqtb8Dnwhfh+QxTZt12ju5ztOYzxhlwU+iQ0EmMVvUKLVSWwH1k32UJl3/4sMsl20hNmjnmK+Zy4
rrdVJer6hT3vbzx1075UPC7GrEJHAhGl93dvIafNYsOFZdPw7OkqwgRr4NmgdvcRrA5uCHajSrWJ
bgMjq9N4TPKYpW41h9JZUS3kikiJl81xKbRcCyBCei5deEOmo3JEiVofhiQnU0VI7uUfIRwwcjcy
4AxNiEzcFYegdesd+bC+bQB4t0irxfmwwYKMUKksjwAYqMt2pEROZXX8iZYqv3l8CjsxAD+jvzMP
Fh0/LeiAQEeb+WHKGJ/59zyADftUSWHKot1EVwsYG0ELSdvRLs3z4699SgbR58h9lYT8Ovh1JoVC
obZ2EkPktidkCcUATh9Z4AlBwA3Rw30MIaM6MEHTu3iOTiik/QwQuKBZg6FgrFtuU7v1nq2LSPN1
PQqW4FDf9Zq6xhj5Vnx6JGeTQhJNSZj2gDcjUezUtzJq3FSp7/4F685ug6Nhr4w8rzUmOBz1qF/o
I2o4jv0pwVZ7JoGh4SHrUNkOSyCPU78xCKCY/r7Gm87f1OGdJ1QUaAQrn3ij/mRN9ShW5RtTukik
XF5NRIYuxX35EidgFvnIQlGwzz9zLsKQxMwT+VfuSY1mr9LbLn1qlxJUU0yv0lY0mdHSSb8qstWt
K0mg0/x/X2Q4kbSZjSxRveGsgqczI3DM7Ewo7U/gUUNJRFp9cI1f1Qi9WrwO3gVTH8G13qBZaBid
5ggDOt9Bgj4s550uMPyRQoKfx/yoT8eiaGeZa0I7WpwSgMzqBOs5MCsvEkCl+PoHKmuATZ9dQL6Y
ebsfJk1Sd0BXM9y//vZFy7bZ2vh5Dz/Ygk8s2QaNyGaJdr6RcLLW42A7hW1uEHeub/2mhSf8yKoW
D7W22abD9fDGI+4+d66fR1U7wKur/PWjsO/u+STOKdEXI6KM6FOLXgfS07x6OKWnoaajBh+wk1Iy
BLDbHkMUeM2cepPIdbFDyinxAgnLYlN6caLSjz5i4j4y9NKnDNIFb5XVdJKzeQ+T5woymmK/aOdi
42hYwXiAqlXDVPvmQM9UVYv17zOWCeM94YBQDILWdlUPeNx1YGqrkhKWodZ4W8TkUniRe/Zx1U4h
5o2i+J47nYSuTmi/b83f3FfqG+6eaREDlNCPslqwdKyNpwMwm9TiPqpy2YaD4umvVZqSImbaXum2
jjPVdrfqestJyARfnZMAmPSMDii8g4sK2fN76k1XjEMUXglbvnZ55awbsA1MutOYetlE7gM7esnx
PPSzSp+wQkZhZxZmyUOfF0xl/Vzi7KXEUMTYzstcoPbkHpFhO+7Ex5PL2YC22jxGpuuL9MQRl4uE
p3MfxWt1DDVmGGSqD/ByUIu6omMIwuYqL/+ml9w5e8M/+m2Y9RbIg4RESNXJ4Uo3GgSWo1OFGAH5
G6D+4wyGpW+Czf6U8vCyy/nljcr2iWrTTVQ6BXSB7hQF38yfkqqVS/UDVJsjR3g/vFJ4aZdIab/n
zEoo1WkY2Uz1q6zqq8pHgO6MrPTbTP83S03yrpkQpmoYejAUo5Tj0woj2YPccNt0Iy/Yb7KSIiX/
R7bOpDAEmUpRBkzYsx2a2FqKa1lpjP0iiUdZFOwNwOesQ2x1FZ9lFa3b/bOdyAGn3/QWJDnYL6yp
NyFM2qM0SQ687u7OgOt1vrjRmhp2K7V98+5CvDBVHH3o9slCaBFeUgWIV4A4UDZfM60Mc7uSNEN6
+ECnE3Be7Bxv+OA8BhR85+AeOyJZb2xdAJvfaFiipf1sTCjc0zca5c34M+SuTURrQfsAOercGYPR
/vBC27N3ds03WSCMIyRXm61tyjItaRTYGqgSSbeNuW+rWoQtxHP39NVhQQ55BCYakI0Ug+P3B1HO
vftS9NAMnMnfZF51RuuXOdnz1AE8s0tICPQMTby2l6+g/EMUTk1tf0kLupJwcL1kNwlbD7r9pxll
l+Sv/wMlH9aYu4SLlsZ4RXHZOYK2raiuL5GYHBVTf2JAq/697nJ14gHmRQBO/saIgArRL6ndYCUk
zEis4fIq+7pG2QYoTZVDVb6ftasF29EkevFdmuWAeJmsTm3WuzIwdTcXsLHTseQaeCXksZjw1n6z
ivt7bgA1Vs16BCB7L0ZByFL38CbXzi6/8soZ1cr2fyw+7d7paimyPa4utQs65h2lerO0j40BvZ4G
0sLrGnYMbsSuAwln7mT46y9Dsgh6raH3hqnbpQvsWNSfEMs9TVRO+GHDs/+EOcGAk5H5dOoDHK0J
z8vk4EGWuF2U7CBn5eHV3/BFUWEKhgHrVqe/ci5+T6I/Cic9xVvPPn00M7oKQlWtb9A2jP+ZcOyR
seKJMhHfZ+OUJzvBJqfQ0c8EBVe2gC9Snn5JmMtXZuDdFnKnVfDcWMRrQ7v0fe+VZEIz9LnEKgX8
bqgSYHTHobAqN3F/jXexA3vvBJGIyQXz27bjLjniVNQlrbN8pMcXdUZkCH602PtRa05ksit9xL2Y
4OzpE0gBHzwMFHm3KPlIeU9nJ4QYARvBcIDIDjorwfSM9oH508qa/990LWgP6SMgycETNRy9mv/p
I2WV0Oj5GTQvcWoD1Q7+TCahxm4udiTZEFtXOqWe27MLa9NOK2nPvejLgKjAFw0MQPK9JLnRAELx
QTswKMzGQr99q/fSfpHpylBUIW0ubnhG+o9ejPFynTPxRVALYC3PKABe6mCtgHQgEwUWfTpVSPZ+
zKV5pcqUdR73q9pf/fOC1MBjkCixVNsA5ZivzpNInWOqL9gvFMo0KBVxNv+j3g1Id/JntgG2epPO
LRy0cFHy7nMapajrW86UiLa7HQF4WGaNk7KnXZpstMNuxVRAP5tHL8a8j8oJw0M2YZPk/w32iaZM
vPu6itfE5cSIIHPIxEM/+VVo/4cwmIs2o7/P/rFwNAYC8wGHTpbr04GTGXXizSf9BeipJ51sWnKF
REumr8PsCvM7fmS8uqc9ZbijE78l7Z/Y6DQja8ZNz/ysmt/C2QbjL6wZTH/p6VHpJuS8+G+qp+KH
VoK5g9RYoF2gbKfS+GZNET2mfo3nyrGmZo0kKi0vhzVIFploQqIFIiY074neIp8HOGlbgjZI2DtS
vT7pOKKrjfBHVl8dDp8HGceDFxBB7OPYLibpCwo9YDsLwxuN8KqfhoGWdNCUA/LVcYdpGNtDF2nJ
TwVKyUFUs6uxYt4d6E0PYon3u7BJ43h3QkVGms7k0IRfUgZrmQ6ygB0+5tsBQFjVx/1/NffVqsQ1
xij7US9aoWUVFMIqhvoVSdIy/LveePp9HtPa6L0wtQ4uobZzgXeG/7Em/DQyfJ3ntE2AqDxUnZfJ
g8JtVSNjux8sEoZ/T43yz/1Za3+s8gsCqajda8HWhrHBivY5IXKlne7R7KyOkkBLzPq/N4X0oa7Z
PE9xPyw7jR2DLIVc1H2A4A4+IRIjf4JdC8fKLuT4KDrhveRiX68b3VTsVQCX61TJRqveJFnxWKPX
eO7WunP/sJjGq02lBWrg71rQmJTbN6234JhO5KlXzavDCseliqBQvKp/Hx4giJ3gPr6orNcGnI+a
m4bYzk+0c1int6EI5O3ycuDGDjrYFm6bdjpNN2lubiV1tR0FDBmabM0afXLp+D5BfuHg12Bqf9jY
Kam0BNM1hMBHH4XtqqcaxbcEmXaqcPpCI4lBUn/8HVdcAQ/v9neqsMheip3JKfADzPVmymb9S3GQ
5aIUtMWjbGKJ9gcsHMV6/nDQQvI+HGW+zO25qMpNMtyqVrRCXwkyro1HiJv1CYUqVZb3HWYYQuaJ
g7JioeBXpLEgJdE+RdG+x9EzAyggiSmzLaxCu9lrPZhH0q1nz6QY+559nGNJsX63oSy1o0RHbIbz
68JOd5SutePhSEQKCXAdvKZjuTkEWoqfG4KRx/9cPDUTabwZj/rSvYMG70Pmu37DWANjCA8sgJ7t
xkanyvAhO4+ub66emF6djxfMjrsrHiPw6iexbJqq/0qSWEpEsHTV2WT0WjKxnR41Na2nbS91+Rc5
kkfKxLovh+3hFQcasjYNHhasbWVkYlKofv3i3YvZRe+r4HkZr3Nex7MTlK2GCLp5ObADxTnprFQV
JCRcT3nU5iv8v1/XRXuI6QUnA2iAPZpOSP/J633y6Nb5b7XbY1XORYIDF9OO0n46Ej1y5TX/0v/2
jEBzSdMpkaPSl1UKfR2rIQ4p3h6Eh95oRYnmL+lND5EIJs/zJTKoKpSj8Q7qhi2kncV6Ukuokcvh
4AVJVTFouCzlsACv6JKbUcHAKOea6WbSHORXoJk5NjVvkSp79qSTwWKa0AWL2TUqUCIAjowICVCf
oEEaqziGwwnXyAXvfgpM3TR48YIscS25dFvFuN00NBuTlXVT65pTVMSXZC8MWWsidQeHVcoa4AtH
AoFj9z5xZB6S2u1XXlu2qVNb67bwcz7X7FB12Hge6uTpTr+bWDJQs5LqZRXacKkqHF6lv6/JXjHV
Ijm/GK6uiVg0rOFaTokhOeDPqgkvAaojNM0M/5eQRYCd3ZuXvUw636QmfAQbItltmo+0V9aJjdli
rean+eCgXUDAomvMOnFnWy/qKQbbeDKK6N0iNfBqMTrZGW57Ky7i21UU/NYD/pok5W/XQsk56nFp
oCyetZVcw2Fb/H67xfCMispu50O67Ie/N8sMwxvGVnwyTl9Q6kV/aDiIoGoYkYhv4xWRwOuW0drg
Rrwcz84dxWv162km5k+sKHatEmajXW+F6I6AxkFZ2h7yjUDPx+41DUJYwuo0aCblF6bBHEY5MjXd
Qt8Sh55Xwj4JbwtkmRBiFngCV3jgxaiIPmwb8wPxpTfZBXnVpImOvdevhTQn8MyDNfZitUTfksIl
keEk4lEVa6pYBl0U+M5T77iArLINUyZ5FhUl/tdNECgYhMNc2Y+126l0r+0wgOHm34wo5xtxArqS
0sEkJReQJdhANqwlD0MNEk8GU+SvegxfBbyh52EEon4fVc72oNjJ5ai4cEBrM0LNuaXyvbnzSTly
W4UFopbXffJOEqO0OrfUJMRI5+xATZQL5te5GrZlWW8e32xQ9kWEQW//r/7zT9lbw81KiBbjJSz4
lWGNjua9REgWILqGO2b8IFTVm32rHZhk1QZiYtA/gEnDViNEGZCsUzODOQ4GtFyADE9+/IDZPpRt
u8uKomH16bOVVft+koeYJA4AbPVWqYtYhbZKJ+ggKR/MsGl9L6tTpJvmRNTS5CIAG3VtUwRbHser
Ixrjf1btTrmCbeb8qKEbfx6qHhtE5NqIY0yisphH0cyxCWdFVvoKnjGL8UolWPerSVR+Xf9jIFfk
dH6mp9iVUnS2bi9w0ojP7iOlBKwmgybHLmErslVyXN6rHKRl0Oz+Go8T5iHsWflQ39+lYxYCZdrC
QIRQdnlfaoKcIChPhvX6EQJvwuWAj3Jppea26h1R4rZH9leXuVejPqncOhvkbkb281h/B1kjNgtB
ppRxhuqcOEFDD+pNZ5pYTgT0xEBbyuoLizcVh4gnYVzbUTEoB2goaob3Xru1IEKKnn7jUqeP6Rsc
6tM+qRZhReGWmDwHvSqtfrTgBXxepuxR2ZlZU0I/dTbB8lkfxPHLTYQtdUS65hNc3iyNV1lkx3dF
SI04aBb68vGZtWSDMEZoXKTQl5pxb/FgdMO5rS4bfcCPrtfg1x6WzoL9Uzm9Jj++nDIHcToOPqsd
7J7qW5jpVJf2+SMGkk81oximQGEwUbJm01j2IspgHMOZHzERnhU29Y3YLD1UyhPqEDpbVJtBl5Ur
Svt/SCTfR6wCZ9LjzOTsu198tfrmO5oSS+7mEhTEFMst3VNus+51IbFyPPl3+ZXlqnwc/k2PRUCv
VM2PNWCBjzJ45EstGmPiNtVecvkuhOwQ6zP89tg2GXuzbq3AJ0Pbi7nIxaQ1RFNfA92QOCJ54avl
MeaNDMto7NYDInzkPmLIracGZfp2YRA//E1JzUuyTQnEnI/pJdsLfHI8nbKo8diI+/GxDiLcrnFA
bxRuUlmj1i/C7q0cwbGl7WdYU0i7D8B6CBYfY0m9kCF+EoPQTAmHs/VIRVquOkkj1RKmfGWeMr9X
nb1igdur1Uhi4DYH0rmzUDFl6wgLkf8eVe1oLVURILoDr8/yX2it5va3xqfkbAemJ60ZPhfR6rGP
F/VRNN+tMsEDdidTxASgH2QnGO1j0/GCX4N2m8IZtLo5YfejMFoZ9iRyUIY+nVl6zDHikG8c38zm
rbah9trX3S5HaCi5JoMzrjcJGpKKk81iswpDLDV/JU+YELK9kap0FOCfyMh3nkbqprbUnmlScSH7
KiPJy/bp1laHAl/a9GSLdRK8PkqObkINkAjrkSOzlgSE3MIsub/bB/RxzS6+THAJcnw0/god+ok9
pRxcAeUKTaYBFWByiIds7vqZK0ovWxsUsLh8mxO3x03dAjJPoFXTaf2g8QGehgsS0r3CHeugecq+
zXUNKiXKnk5WVTpJFu3vqBwtBNaBojh/c/vGXH7zHjqTLCX3yxdajaqXhP7CMjDfDOB4tRn6V6pe
3oG7+0Xq3+sv+0jhOKcQHiwoBbXhFk134ZQQKQY96+cW+NCGy5ZDXpnXvmSfBOdnrD161RMqQTRv
287Cfjr6NyXgCQhK7RY3luMICXwjmdI3AkV/Pocs9ou2r+mS0Efndvnagp9HK1Rp9kwrogGhmsjz
etOoqI9XaDO0B0V+sDHQU/xT4vj6VrvYZDSh8ht152CEvu2YCfgFz5ZcR0DXbO001P78xkz/0vQw
8qNxYD203gqSj3M2dVaXrZkOrNj1+GOeI/opecQOPKG2+rbKj9t6629ku3qZFNhUy+4k+b9ZgmRm
ZpLAR6sc5jVP2gPq0E4d8FoJP3uuBWUz61NGC6/+fT0SbZTU/N8hNe1v/JSOObv+FFSPYTH1i5ri
BNCpltasWSV597nn7DpGnOVZYVubZ1Wv7MMaYyCAxLjglQuZeevwLAFhDnBGz06xfWu/a5W2zN1R
WgtezzrYxRfKpaUApJrd/IQIupptg3cSuEF98xSJxMl7P4uqV3yXHox+mHdj3ZWFCw1xz2Atm8o1
Chx4Z8VH9C+Rzf0fDy29u+XQ3iu5a7/HdwURzwpXXn6ppF7RPtRishUcKOQAqcilOBbQpoPYoQp1
Mr5GAl1wv+uOadbI4NeMRKljOUqIE+4f2coGGVG3jcPYtwTeyuWlGDGiKkQZHn8BI9FFNIyQVJNe
dFcHvtCLHksBjPJ7246rKOvrWQ7zBkeep3bxBONcbNNmV6Gkx9n8Z8zROS4gORQ7eVOLhYogXd/y
FqGIKsvbZmolXdOW+4s4hFckQVyl59RmJuBK3b4r592Z3y7i54h2DMVBBQKEB7FwvU+bFtFLcOP7
/ygml9YGR9ucUwIph1FN9kxyMjGhsVVMDxksfOr+xTFFazxCRFw5vLpcEps0Bqmt2eNNg76RUJhm
HTf37fPWMQor0A5Uy7+ULvmdhxgTvFjouAbEPmnBIKTMYwPms5L6dqxPfBGG9Q9dkI8P2/zRuCzU
jwjH5SNkAe3I427elIvcHRJGUf9Gp32PVB5acscOOSbb5431MD2dNt9M651GEU81rJVnZCgvy98w
KzAiYC+9l26arqOv9ElIB+SfgK5Gq8p8wqqi01UBkzEh6kPCUd3MwrX+1pLItjVGYCe1Xmzr8Qmg
kFftjSrgAGSNnpF+MdTDRjONzFrIRzHM3Vi4Jp/AnD1IQi8ySo6O7L35DTfqEJSkULozoHMewi0R
j1T4c8Y/XH6/sxIzvuWXDpBtXMIssDd8+QQDMmG0eIM6VHk+wbHnC9Pkd9Cwxx82GTYIWzQeg8cV
eTLvz6IsB8QYwXqZdnnPhbhkh8GJ/M4wOXfYnCYvL/d5z222xe0FiLd6VDbBPjt3JqVU2bsc7quN
bSB9tGfgZZzVt+XjKf+7KJhYslBiDYxtZ3F3kxTWzXCnY8bB21efTL6dRlone80HY7japtIo9SYq
JS8jcY0cKURQb4SVzRGg6TMWOxd+SjMZpBuyzboaCyhYzMJBRo39Z13qUxe32TogKEjFU2XyySly
b1sUZuPX200BZtL+PChrJGoMqJpxkSIsZApd68UUSJfljJsQwwB4ND+uGdOZ1XBB0BzWmFdB1MeH
Fe09xjJxFqlQIIDeb7qT/Dpjh3/qp2s02hqC1eR9O/NFibpdCizxqSzJ6BLPE7TXacpx6GfjWGyT
GAQ1Q5JN/uXRY7scjWJ43pTYM6jo3Nwt9EbyTCKLgJTuDmnP6vgFsBywLmjjGLvQHGbKrAv9zqyg
O3YCxLcQP2L0r1Sb9g0uF3d49VNLVdiM892wdGE552gCC/kGx36rG3Crmh+rCDDQKXrGqh26/gHU
dY5khhNc3c6DPy02BJlbvyb+gu4ZhMffYjgZGciTOB5kBT4l+pHmNlNUDMDNBvNFqBMnR86OQwtM
wQlg91eyg3XKTXCiZMNARchEepw0FcGwnPxOrmB/T8ODYZ4XFN3g7m5dKb3Ww4Vykw69Wpo9ssWP
jwE8Duvtf7seXAyNSKQtK05BCgvuv5dnmRvKsyE+Q1FYib1HylF9AMlhW0UKSR8Kq4mSbZBi3QQF
cIxZu4FyAYfFOB318nic9tw+dfc8xH4GX68PpIslPQtGJFsrkmuk3iMq/SDMQZMLrg6V/YUmNKrV
kxMp2Fm/zwP8GnyE6t5+xfHnvz0p0jAPqrgQRIGsxSxJ1BWNQNb53BzcKBYcxVFoGweTySTA8CD9
87HefvqSMX4FdLMEx6oblUfI6pJ3Wlyvc7H+jjUgawzDkFpcdqRuqj1HtgTISZzYeRx9sG3Myrzq
3VL9K9QnAIsohCFqpMc4HIvVXYkMh5PRACOn8hWhuwucQK76XHBPw7et0V8qgV1dITb7Jb/1scUF
KwfMSBzJ7Mimzbrzhp0lPqc90YQCPUAltSybXJ2HOqejuWO8bMeF8aA8UxCocDxOuomXbXrYScme
bWqPOT7O+UQlFtwn5Yn7of/q5LGKlRMw7EUE47a0PExE1gEBJ2YqvtugL09Vu7sSUCHY3K/kLnfc
X8OEyn8wZgvH1BP9rsfNhDfSTWUhCrnFkD9T7BXJoPmjP7CGbNGTS5+dEO5U5IAjbtxTjGTtivtj
D0KWSh/mOf9cRFgRoE3qYVTXacfMDLWZ4Masd3VGVgy4we8DexuShgcM9GKVMeYd4CS70RSVEOFm
XpuX3pNBJ511gfKio5wk/oJeNkpgvCMBVO8dYtjKX/28kqQBCzR3kQOBMTi9JZU5hjictKbKCNZj
puAjd7yF15pLRO+h+5UkBTS8ZZ0g35QQYserXZbWN7eLORaloUne8fQRHr6R70zn6T3qhcfvdvYJ
7CecY3sAmEU+ckTjn4eq2OKUD636nY7sUblGkF+21zLcJbVp5L3lEA6m240yX55J1E8btnpwtz7O
HS1XzK26oK3d6PsOgBjtCQO+Q25bRLB3zADOugnMVNUtbcfN+ECxQHd5JGegurZMZ1zXm2G7UT8j
nviUkldTFOWtb4vC5RrZWlvc5BTdLzPx3VG7tSXKrYRdOGMeM36D1wCA3xUa69DkFbxXiJDIB4Q3
KdBtmwnGAmtagHHfEPCektCCzwo4YTCW/CXOE5FSb98dL57rB/sLCgLd6YqkwHsQ5T1OvcAqZ1L/
pBVPVJa+6Tqr7qXs1yJ5fFxzSmmcEuGjSiQMzqBO+d3tjHL/A5rxoVvLGRVNMydUFWtG08CqdQrj
3MkEy7ppvlvsgdwyOTmC7hsGMLuW1lVhE74OtKybr4cDFRJD0L/RIZoMVSqS+OABPcwIvc4rVMfV
0/zEgCWJSUU15WSzLIl0ttBT+DBfVgV9UtufPmBNulg3u8t2ipdIWIocY6u1hXwgrisgYY25QbrG
qWm6H06tIHZAckFayV56j0THIjsacVFroxmGJPr+saal1SAly8BNW9a71cRSqpu6kKastSVEAVGV
5botO5u02NQQ/pfNKw/G60zaxoJc0lKKeyukPMRJCeVvKnNOMwB7A5RZkRPlF+PMYm+O7hnDVe/E
QLEGhxiYkKTO73xkEj7sePs81WEKzv0Z/Em49Lac+/18HvNkZ8/gjQ6/r7sFj+Dh+wNDb6D7EEO5
fjUIJaU+05cPqHtcvoSZZH/f0wy6KGkgl9KCttf7iswvEVYDj29PRO9/xi0R3D2qAO44xvlw+2Ry
Yzqs7H+/m4A1fQf8EalTx+cXy4qQINDZ1LBBopYfbtSZvr2/t+6PXRaKhXo1H9Rv2uYrGamfRZ7L
fX6F6mWJnTn4QWGRFSzGxqImNiTHf3M6E4m4hkr81Sq/x7b7ArIkfaWFbWzQ/epDwBLeJmganTCy
S/2EP61P1e8fAZCQbF7JN+fID6ku43mn/BEJZ41oIUbw5JV5lyDNl5kcJ2nMSOJQV9QLz5FZhGxu
zePDWXzlXqn7Gsh2pdqSD7qSqgyOED08fkRBtvRz9gyeLuEmhH/ASyjfY4kM6+4RF7MGQ/mMaFJx
rJnuynrKGkOsNxh3/z4QOVzKYwVWXtLvBGbAHlMvfnHv/Ig+J5Znxa/TNCEsuzqy5R7ly7DRYvwe
3MlNejAkmIRo6ekFfK8xWrmg+01qzjIbIUcYln6K9PCIMXqwQR84jMtuLaC39WwCnB/2W7G/GloI
jWBmqNT48jpexZMll5kHUaJxkKT1a7SKi2UfbngbfvJSlRR5d6CWmJnixCKyK72854xyNUJwQ37P
LYkT4W4Nq5G5YUyLDqynIOD0R7a8aaxtfyxb3168lVw6mXhwx7c/S4HEdlmjeN+q5SSAr70AT45/
2fKBUaF5sMznj8wTncDbGsgtBiuGUuU2kFxvtrPqKHR7Zpq7UdU/0EGFgvP0+5OoX7xJByhbJS/t
7vMgd71fm7/dbQL+ptGWrDQkhI2LSJms5U4la+iBAhCo833w+Zfvh1BOhvSpl5EfvlXT+uL6pMsq
tydFv5tuV7Dbmd+/hAMx3nJGMKIuKiLwp1sO56BHEH/0a0BBjysy3kzneW7vPno+aU4d5dbUQlk7
z4Sv/yerIiAR5fKhZnb6u1Fl1uIdKZf7xxw05XAaWak2d1uehR//fzk4qxopmetVfk9evZGjCwq5
zvj9+f61rA/37ARzSnlI/ZQlADbihKq6667m24mWstzP5kLsOvdAP5n8Aq9SqGAqyaUccT9dW59l
2knQbEXp4fyCrqZGig3UBiQbLvDgZKRbb/uGBWb4koV6kokAdcg/TN0a+vwfYv1YkHu0YhGbDJPT
38k+97QzPXElBARGJRYVpRdfoe7mzAm//MIUU59Tpyl6DCi4Qi583mZjE7HQUjChBu7b4obm+ylA
nodJJsT0R56CwduPFANgPnR5VyMtRkv0lVU9vSbJqlimfGmkexXfslItcdnLr47ohKcuOQ9HVh83
QTsmi7gM16ewRawqBB7i4wFt6bNR0hJPR32AiOv45lNljCUWHj77JaRBzCsHmTv9YMQprXq2H68a
xUlwagPR7vhZUpLt6lUcILr8hi2BKiGWE4ohmfpmWVo//s8BtdSwlM8+pvMNk8llUg9psRKGsy++
VmQVQ5dhNKRxEBlMYDI+4UBKVl7B6vrXTLQkktFIwWHKErjxukZ2JFPPkpTMqrWBNkuM/OGK/t3p
ONoEs+fuAQFPQ6IWEug1fx8yd1efBT0FD3xaAU2RCjl4y4Tu89SphPKY63oo7QpNHmVkEJ9geh15
Ux4N+7k1jj8cZ/fVPnJ3g0sILhf4Twr/JAFVsNMWkli2xqsFqlYsWpdG0WrqIbBBoZV0PIYCrcGu
XhrOvk2dOw8uDG/h/z8koJ4CQyKj2ZrK+JtujxR9uSGGHijw2eAp9YiRE8jBwD3fmOwcj1ICL2mG
QIV6SdDWTrUUZF1JSGRJPV4VUldhSc23OMqt/nl3CN4GpJTqCoXmTLjPQfaAjGG6Pz7E7xUzME69
IBoHR8Yx+FZxRNFV1j/7IcyIf8nvtb3R4EYKThfa1eRJ0JyvnG8HbHrh6y+iqF6+VTWXuW9yVtUP
bkr4/kjNBCXD/tjmyU1hOnkQUwKlX/qk/+XGCF5r/v4lNK/a3crhvdTdID13Ea1+5ymQHcIFdkBX
oAyOGUyCV9xIVNkwWOMvcXEpYlDUGnHi6wlYt3A+KPsbCcthRAGXIFSGZvHJzPqXDTvpycKag2wV
KmksfZdIP/6r1Lzmdh4WwGnNPAtQhk0NV2Jn93anmRNEBR1ZLq4BV7Df+EvfnRiW8MNVi4GVQElu
xpHor4ByGeklZPlY3uiyNFfGmx3+fJU5cCjtYDn/ZMgtcP2+CQatx8kBE1u+UY9RpK/N4ShrUqiS
Ptv+RHwBudOIjKNbvIpUhRoYaQdlb+y6vJVMDACeNGcnevHw0PH9E1A5Bu0bwWMHv2Beix23q5y9
T9Ympg5K6ShTKvYa3JzUGfyjp6f9kvW5f3ZxgdlkwHt7hWrW30LTgdHumgTxntMJ7X5Qy9Yy+zCF
9PapN01tvITgdpH7nv8jUeYYkr/snHUS+r2oZR24CnppX72vBHFcqtpvMOmuhcLStdG1RTBEqukA
DcKDQM84vATwbLvJQqLe0M1mXhgqTgYFJWjCJOuDXKZvbRRAfE48wHw5GBtSHra0q4LCiIVMosPY
tXB3KvAVLQ28KH1nQgaZRAcQX7V9lroEZwuGxUB50nPDol9sqIhkqU7J6kNKiTno3pP/mD35YCAK
J58x+DYkch28CwF5a86NVAFMSPQhHhKCnVDu1re9ngKsyu/uaaa/F8CZT98bZ02PUqL0VkoZfv0b
msPQi/W5xhXiWeWqhaDVIFAe8G5nVaWIHFyoC3seyN5px0jswvNpoofnZ9onHy0Juerma4TageIk
Flw7nNr3BtNK6xWZmuBvLz+JtSCgkYnQeIoYy8o3yB/6WW+VehUGmH+8F3WZapmIVQrJtj1gQCSx
WOaA3Px1VTEfqv2UWqoIryJWL+46bSsDbgAXXrCfwd++fH0XeSDaSITqc4uqndr5ewoODtgo7XbR
eulsUe1lO3i3TyGKZp7tIxRofAdUDbjTV+YhUx/a/Wkv+rApRTEaeuIRXUIoTwewGzpXYnvjT7Tm
qYhIzg6AmMP6yPhGyyudDs4GdheEvAlM6f9WJ3dy9pGkXxub2HzCHvlgGyIETIN/uThw9A3DzvKE
JJOGtnH/+Iba0J0LElGX4e/XnCmOkznLRxFgBGt5j8BGRdVsdKYgv+T0je6bSqJXJxA6F5bkrTed
zKCud2NdDKs6aBWaBgFdP/ne049GjShIjnh85r+E9IF0P2ZLgEmOzsVQtYzJ7Z54gNdnatk0UkLH
ulB0JDi9VXki5+Odwk1JMoTcNw3XI/iSXZmw/zT2M2/o7C9VvJOGMBWjlePCqKpQp1cxh7Dkk5wq
qcZMXX8fjIoFfaREPzHXb48m95iolPto5Az5lbUCl/7IPAkbnHJEw7OipE2b9edrhmrR3ikloksP
18GLNltKlngttvwz3cCvLigzvB5/bQ4pfqo/Y1OMRrc4ISM1i31h9o3QJ8bTJyP+qWWwP99y4iGr
vF4+ynHiYsEqXrOM6zeBmRw/lk1omCUn1SWChj2Y7NWxRx8EwiMhFhn99sh6a47StF8Pa8jputyl
WppNodZrN/1n2iVWHeeOJQy+Fbx6nxSXmLyNI+vE5BaT26ylq7qSpw49X9V5ZTFgXCyubxLey60h
7clbmthj1Pps9s0bdRpeSJ32rvKTHUsYQmKAuvivrF+6UhlL66bLLThENacWGl76FvJVHoK71ty0
hYEsX7S9UJTNjSFrqaSDnn4bBBvbo/+VBXriCNZYv6AnX0dJBwQY5zXYuqJi1pvncicvp1KkZQoI
5vnA54buczzOCE1APW0j11iA26VzN6vWhwX5MwDZU/TyhaihVLurFdJvb77RodynxZ0AXvWTh8C0
x0/NPEqHx0ctbu/iCKLoLXeRB9BcXre5kfRw8h2s6nddPvLWWdQQR1UETxUfBviXPljuOvMd+aOT
LkOJ/Yq02lLxmELcaBtWRHxg0yoXF6rmHG5Gqrr2yYk8XuJbWL7yG5QGCVHycNk2C+DOuawlBkzc
IC57wAhd+ajDc20TMmPNCmz/EL/POsP621NztrXHxUq57prDeACNbmpfWgwds3V2VolisBLvefGg
dOXEnzA1ROh2X3dOcBfEQ6KBHjFMSDF0VJ8sWLftlwFc29Lcb6QurgZqnsaU+ovFsPuw2TBLYX3h
QPXCE60ShKYRWT2liImIzdisthN6aN06anf8gia4GCcrbCTCFjXkRjUE/LqXv8OOoFurNqOUoRIo
oXdONq+tYbfOa5PKIumR2oZvwAkQKJafogl6eKlUbDjlac0xNqlupcLGcEN9ZjjJPxdG/CvMTdNH
BH6sRU2MJOd2kj9RAowy0CqaYazH32DjA2HcHjKt7gcaeg2FYVApfFe8eAwkfR5CG9/uRqcJzeu5
XnbrssR7cqbk3wlHFnVUR0BvuAS8pAvYBgOJwSxh7XEbL3wK+xbjb7+LgpZSAwxbCydpdDvy3cm8
2Ft6Pp6PuEl2LutDRzSBotnowsWIIfI+ErN7wz5vfbyuS6Pw8TK7ce/dZ0NmKKOb+yhoqysiiXDy
kbKX+KDx+XR/3aHzTThyDz47cZpLllDdyVMP7IL9lW14fBamOeWCOIpG7M9LJ3eIYXLkHPl28s+V
CL0CB7e7C2kv1gC6/DxdLvFDGvUV/pq7YoXmkXuFfWCL9SjJwyPVUu1RKfLmMF2vF/5oA1K8carA
PstOdNvFJLyBeru6fRZk8zIoIV7BELXhF2aikwIv2bSfyDkUakMqRnRiKCAHKIgssjWrbX0cC3Ns
eAtN0o5UGs4eU5x8beAD4PI+RSFJlcdu10BuUQ8LjdhvTS8Xw5FaM9tLhCJd7mCnvoyQsJKgnyZS
vVR6WhhRLv/bQFnJt83QZf0Qc5eD0QQYzkugvzfRw7Bfyl0lZTvuQC860w4RQtDN8tD7p0ZqMBoR
pN7MjHj0ZyDiQRxVX3ue6P7rnyfEAfsKnGOjlukTO39hVhtWqINnL4SiRAXzsnycV3WqfiQoWzH7
WlafoDjVIMRLVB9ECWsX1zCXBBTwF2h+fRk7JJGkfd8iiz3Of8k/JU/ztlStZdsOp2ltXB67+4fl
mELk97XXri24BEprRUR9mmoZeVzHGoAu+KQxR524LkXgoWayiMTtzrZvn0uE3saDVLUgs2FAwn5n
l95odkmgmwaU/3OkxrrB2MlB0hjo20HHFInIMD7/7FALIl5er9eihujpQSRNeMJmR7s2rl7T86u+
ppgNhq0T3UUpiEiLMQFMaRW2d5e9v4whah2qngaTDUFY3hKdbgwP2lmeTYOveKWlnkVnjZxDuO7Y
ZQ5l12YQccY78CohBVHbaCCbMuqB8yJr2DMo6c1utMvU1UGb7A1Bpbs7SIcpigBNWOK4CjWRDVMF
rz3E5gswkPyvbAEVS1gHSBEYaPuQuVvGUN0+WU8gTA6DtAbPpUQBDlIR0Ckwxn/yXPWZHHeAYOIk
qArkXMW7q1Rc0oDoXcOcb5L698YnoFLRrJ9hRsfW9L4t272FbSrV6KmwuY0DjMsiJQrFgZO334i2
PcD8yG4t3oezxGNuruFVlIc+0ZiqYPXGGBbz3R7COrcm+H/4q8PI9SHobwhqO0pT0hGkG2A2ii3W
5jG+GUYHxA/kKXzH4vshjrPApo2OZLGd3KE1+gbNHKH6y7ERmkeEBIL8IeqV0ATnySi9t+PR+kGv
K1hiXTZCDP0a7UzXisup1EigoxYWho5iXBXa/N3ILDg/kfLU1tv9G7VAo295+/x99FQ/MwY8owyi
DN63bn0aNpTBFeQG9yb7mFWzK3iFZE+wEwzuzaU56NI/JBFL+QjNMTBpPqqaIvSTYuY6r94/2Fzw
X1xnxSdTkbd3RArmes7FIHRYwebwszXrAj6T1550uBBjORAJrmrHd6RQEonUaUOktmUpvMreSE6N
PLK5OK32YiYkI5PJQOB+ZOAMuPMua6QrT/flZmlpVExcTV/xaEJfLy5a0Qjj5m/40HE6wxcXNTy2
U//McnH00y40AE50bSwjQS8tHije05bKp2QopEnJ4NmM7SJAq7nn8FflxKhImj4iJ3O8cEccF+Mr
GAy5VfD12X9Hr1HujIgsnsOPcBi38sfE5eB/u7PjrwxaPzJCH2C28JkaQ/3ojUCH45CtaAIvUNOS
spvcGHIJc0ybJN3smsBoA7FsjZV9l/16UgE8dxmwOgpcRlkN9ITxFCmwB27InhiOZ0FAwvvWiDUF
cl/WOhodPTyEd4H5jfovS/OoW0gJPftXEYVK0rxkBsujUasVhc5B7VFmF8BZVNefRqfPEvOFpflZ
Tbv8IMunlFha5TTb+MvcA6bMtI9QGDbmQNssV+gbfunT2MtAl9H5q6dL/g553DH9EUBBVvqRmIKf
hqs1Wf0Mgv1Y3wdu+4mYfrvtIX1WxfXaQbyrmfCYgLTP/B/BShmakEvTpAVYfs/eTkjumQXoo82p
eQm6B3R9d5jOflnXxpzFDp3FNk5j3DG3FtwgUdBP3VHFYabdLdCDXydZKlI7s3ynmtwuDzYXpS2D
fcpP3JOhR8Iyfy7x5a0nHcnq1WqE3sHZtvyjAq9haGxLn0BwSUgno+C5d9zq0M3SjQRFgzejGTQ9
vmCBr0iZdtU/2V92dYfOsILOuGzOD9tZBzxUbsb0p1e7Xo2zSz1yfuDgIj9kAeB5ioU47Lod2csp
oXo1LkTVMjEjpEhYsi7GJOrHn19MTR9YA7/MGBQ0L0rcXLow9yl0/1XDxxlJ1RVCxCpQSZrkpSEn
kYoAW/JUw3wBafLTwUcGuYdGSjFqVVioJK2rq9nPUGXWKPdiK403RdaMdvoPZQVkYChVRpgKqHsj
JuA1dflokfFtIkOu4RZ53D89WRrsxJBYjNkesyfXXfs7yh9jEDwVNE72g7igBgrohLZ/e53NTFrx
IRmk2xJpaapLUcZly63jYJ2Sia6Ef+DrtpYdMbLLP4mbMHlZuiaMhIuaahPdlzRJGBcINrFvuP5y
4F+HE5BxBJ4Mq8t19Nq0gXe5uo+Dtg4WWc+NcV0up32cp1Jv/Sau8BbFmb3vReBjkjcXuRq682mN
9z7qZJ4YlN2JWvbktJmIin2mgVQ4Ysica+AQr6to4bv8cWezbCKuMYKWS4EDtF8sk1EktTKLrBU8
aGDNFsFkAjedAW+ehdQqYV4znUxHA3jVvjR45eon0cXDlmI3GP7FGKnzVSxujcRkKbfAwewCiC5z
dKLcSfg4ajr7bAa0K6avBPdMir7Mnba0oCeB+clYkqPYezfdtqya7onpYr4WCheClkpDWotu4/0K
cfznbInToLKCl3xoWSd6UkvbOgLhZQDMDhVVgvewgG1QUc03ObhUtYivNdbuVUXy62EsUv8rQ1h1
1LDvmrQCfT+VNkjFA9lR/NWdBAqgSDHcuJFvh2sDvDqqWV691pg/Aji2sTk0ffMDHmdKoZVmaufS
5k5k2FoBAkw7bkholcqBEerYvhFQ0dNBBu24hurR+FjYAAlj1QtloyphwFdEUx24H6Cb4M6uTO7a
nTnrU4IMSbyHJ2v46Tzb10+uqJ+PNFUN63JeyTzIvqtMZzUc0uJ7Std3+xrwXrYAqCYyuUNVE1Bu
898mAv+FGlgQESnms6N3Wp29NZXhDwND9Ip86k6Z/mN7zoS2jyBwCaqAVA6uyvdXZIRMIyXxUhvc
6+fu1Zr6rriDuJ5rU5mDd/T25jDQ6lkg/plY/RGs/kyC9w+8Zb39uK22LSvnjy2QsqsQig7HzxZP
ctTTYwLeFp57VeAZEeGrK3UqFYLaIRlXKSNW8aHfFlUMHm+7E/3kG1uU5/AFNOkydm+VgIl/fmoO
aTUS9sr3oIHa+bMRzHnIA3SYJUuCbW7jUHxBg9KD5ZRdNhzrer5X/Oa2erli2tsyH7B9yOMcJd6+
OvEN9nOFhro9fNSQJlQ05kNfzty/QBLQWTcIY7Rn2P32T5CKcRtvlOR5eDqqTyzEbqo8560fo6Sf
16yjFNxRLnoZ7wpQAc9Iab8hnwxbhrzD1zAshzuaTAgf6dREq/Y6VEQuC+KZOa3zP2hjMf196j3Q
smmWvjV3M0G1IU1pquNtcZ1BYk6PTktMSMOTpr00jQzIJr2OnH73jsHqwPvEnK8X03SYrC+914PP
mLXTbN2pbfYD5qf/csWmEx6D4pZrqi4dZQwG7UipZ23e81pEfbgbAZP4ZxLSi88uC1vOY7aSHg7v
mH4ujHpfH5u4thY+ZUImYbFW2wJLu1h8ZhWfsZdAo+tC+mIkl/R4hOE+tr+Q4z1SyShstiYYQhVE
EUKGv4C9KR0EkW88t9H1G2xy/Y7MP2zPnlvj/OvEMTPXLOveXT8M1Vk+G0DA80Pc7G8VVTVMQ1+Z
DY6536MvvwAK4nqR63YbUgrF895zpTE7F4J+U/sZwhYmdAYCCPrjjJ3Jm5R6d0Kk6amqNvI5o1ZG
bIWyAybNP3BpGVOpBuOzynF5fuMAZS7Ito49PYHS1wEHa07MAdr6+19qaQOPICnUFMGdHeaxbSWP
2zS/JlJYCoIwJbKTJB+ZhAP6V0a/XuKR9l5YPRyrvcmLBX6xFBSbAFA8LDIEAzjF769/WcNAfHs1
0rKoy/69wH1C4beJCdlNJ2xQq9sDNahihMz/l0zvAqfXz4Z0YOwsuMpA3Ubs82NIN97dXyunv3n+
tkY+2wKzYcxYoVAE+VFABNU8Mx+PIFALimkTiK1y9pFeskWxKXBuB9DDcyvdHbz7grdFdXEm2zi8
3gHeRvAMTertQtdhBMpYRMz7BGgNHtyQfyPaTGRtmvnp1MYT/WqxDwU+4nQ4VQsxQmlVJLWxK4v+
A+VSeJFb3HLbnikSR92B/xBZmF68iPxYt/CLQefVSnsole0TcIQPVicU/plp43uBww0D6ABMyW0d
gHrT4b/pYTseyH/TA5S6EWriRjiexf+B9ySYw+9F+67QGUj3/91Xo2ntIvE+3fUMEGUM+dmRDp2f
W3pGtIY2Hz3bSkPKQrQotTrmdFfgYJ8nQCX38BPlYnqjXL+47epyh55smMf4rYZ392gcJQbAue4w
KI6MoRPt8C5n7Bywq2tmvNwnxz8UaCSeiZDR7LIBasTg40C5TZbGTCcWTp17wO/j1bjuVesmaA05
d9kdGcHEF6sZKchoiyY0/SNG+4rnEt311970PQm3MqCfEa3IlCcyc8VjXyMAgyrUYhKj8wbm9Lv/
QCHgQuz4oPA0S6c9dpeO9aYpq8oLDKanUMsISefIgTs5bPB+wiSw3h4P4AnbIl8TW5LhUWD2i0Kt
7VeNZsANxnO9e85ugwbHz2yBd5XY8cteuLpGY3o6c6LEKvUgw2XKHbD64YtsHsGza1unEFny4wzE
/ezk/mNZNbKKha6dIvHqpExOYMM8y4i0EiKSQiKKg2MLA7QBXmz64PWALHYipup4//I6wGFWJ0u4
OkSoOB+DF/E1RGFa19HQGr7TAs/ONfACEOaLf57wl+e/bdWBEmRGWcXteG/E29ibXCdfDL1biPs4
8iFsOLGO3lHdsD1c67ZPc2fDIikXQWJXrQEiXr0ncgXyaWmxAfiW0+aYYdegL9HHNnJDUytePB9i
JIeLVBZjk9XLCLFmN1c/nclMvKieAEav+UHiSR2JoybVFpvp3+FJhukc4p55E+YBWpZxtEEXIkFX
EMrG3/2RcZrs2abKVWtelni/llUFdjDS2SidOddFX/v/IP1xaP5J6kjqyp6wPIWzDgtb/3vVMxg1
25ldoAIVjhCNuxlAdcBeyyjWH9uMJMrHAlSFWETISuFDt2QQWAV2m+kQSEBTo3zGUCzNYx6mZjtI
7DsKC3MXh9JjEvVnwarzaku3XMaF79naFkOv4YWTDSbTpZ7kOmA4aEusoxFiGtN6Mh7JNy1Okdxf
coIjUHt1GUZoE+N2yPiWdqtqpGQAfnVSteGP7y8vJtDiKAY5urnOLb/osCHCTKef+KnwyPwBAnJp
Sk6sJukKG1enuubMHtFZTHoRimfWQe5FUwzQHCJQoOdOU90QIICbWbBU06fDfkZxY2LXyhcgjVxx
JW22TQL8q9ncsVqw0fwP507+uBBCojvnYNLWcvOc24vaOOwE/KcuE1wGV3js8YH8VlWsOVq7HUOq
WEtqsPJSOb8uupAFWqhI8bOO+MHpxhRhrGp8fRAKdg32Vg9/RJn0mSkr6rD0DoIbZW/N3hoOsSjQ
c02UCOQSmdOb+FvCQ3MP50HOhHAzwAZbZsTLPXjuzV7udUaoUp9Rw7KTZ0ffLF2FetEeFGu8WnuQ
tDJG8EZJ5nSG4u8OpsMhzQC7ZSg27jStMU/YAvaeJXus0cWMAFIURzB2a3Pjx+EjT7thcx+qRujO
kXDAUWsWvXRlD06v7fWq343kxpmKt/iarpH2fpsoezFSDJOxr2XvpCojaS/dpGbjQpM3ZShQ75kh
eK7MWpD5IUS//3w8ihpH5cFvnJgsb7p2OB6XM+NufKYiNgDw3EO8LIyMuauRzI+HQ0F4+Pg+ajqg
F2qwIeAUcmVlAmfKSuMScJ2qy0pA8ojYWJezNnkj9s8slzSESLkkNoNaOxTur//ZYI1ot8pBMVrd
M7HY912HNmdsfKSkbSM1CtSK0mlDM8X1GYExaF1ZIEgT/xq0j2Xs9dT1MAGX7eo3r/qm66t66p7t
7QyBSmRfrV6vLRCaglBNmUQ1gFz1onOSyhR1uVBxjHhQhzYXv6XsRfr3n6J4IQWMGdNJ3TSFJzyA
mdNv6BTooG850D7ePcM5lQjF4kyk8AfrflnwX7cjH82rt6EfYwk7qhcV0Cc3M4ENktEsx65oFfi/
uM2TcaIyOOCl9NAXzY9hsN+5kTDRfxBVRQ5lYK5wZ9qryR5hQ4MkUac5PDP5WNyJkLt70z3cLCus
cyV/EYnGcilz+JIjruGi/8zWR0YjcR4fGDHmnxZOt3h33g2scd1FtNesCoreC9Rjf2pyCbRSVrsY
78Whp9BMho6RUgPAhw7L6yQa7yjdj6ZYDa9RABnLSfRj4odZTV3d7z5p5AEO1cF3CN8QQ5HjXFbY
qU1ggmLn/WfXfHyUqC7G+h0xlU+V+Y4nGzn6wwp6UdT4UwNJRkdqF1+HxB6LQD2iw0osEAA3d9kx
9UjmiYVIp+FK8P33jBSKywE7/aC9y7dRGQujpdXY794yG1yDOlDVCn9lzB0sFwcVFmLRTk2NKjli
4RESSKm2Xh7o9yOI38vAvoERp8x7Q9j0B8KIi7estWVdPpqHR+2XfT7h+dZ/JUz5DxjqG/Ckj6ch
TQiEbHKASBvLkwoTAKgkzxregpxfRqOjn5QZEP14q9k3Ywz2P3I34+LkK6GVbOEVl7GxP18aYtSP
rVL9VMU8PTs/o7oLIF7QEKudgy/PiHPRm1xhCe4ZUadB2eHYmByOXBVZvWNkY/NTIrn7BaFpg/g/
nmaQIh9tMSc2y6/v+J18UbdRyGhed2szfmTnx6AQxLI/q7fj3igZxuxL1SAeunkZwCWF7AclmT2v
X6pjPlUKUyHbbx7xba2lHiBEXmJvOncYuHUHAHMD+y08kvnLbWYtJD8E3ZYsjL0vpjEbFlrax4Ol
5zWl8wm3ryAT6zlRs239/uM51/CT5ZUCFC5M84zeXpio2NravCgl5/7d4W2uE0XcYhW6XBTFcgsJ
2J4kC57iMoZScLyoNxD4c0plFHh88Z+S8NoZZRpjg1g/WTBTOr4I/RFatj/RnsoRNn5haa6VyDIC
6NzUOjQWRnkuUFp/XzUcX5O4HT8K+UMJh85+CRBKRyI0yyuGl2pnkmp4aZkvIrLh18pbOsv9APT7
afwQj86fbVofxYE+qT05U7RbxYeWRDfklHW+J7lziBHl223zrwZjWrIsN+cE5P04B1ttlgs2ibt1
PRTF0cJwJNy/+30QDRIihUSr4lIRIb8xOTFREgjlt+CteA+Rxvw90+qYaX9L1ole7iAoUn+lakle
uGdZR3IIbTO7QwuPNa/Klc+Tr5oILlij4QOlzuvSk4fY0TIKl+v5nMPeupRDkqQuKttlY1RiWgKW
BLY8G1rJyKWD9U4k8eVOwwRh7rIyMEVUlrfSI75y7+1z373gbXtO+oM8AFXu8J46t4+aghlUzv8X
zOeAO3s6A6w8tJnK4mmcWo/YAglPGPNvH1WJnBeRxyQ+3zyuo1lWkdnAuN0TvnO1e0FjewjPu6fy
BoP2yQNuzfIFdAIFekcPKr4H1gsRztzkGgTWEmY4+AygLw862Fm8kpLNt+AcvPfIOYY9mOOsBX+A
Sy/Uvs0rgqbEd/mBV6M700uTI5MnEsAgyJYukru2C75NFgaEaVrmyRZIfJzed+VckZeFGEXW2Gr+
cJWg2MvRP7VJcEjhbJGU2WVkVUHVJufZJRRs3pYef1RfnTtc8ZoyU2KA9keautapgOqiw8Sw8FjC
tvRl4IwT89e8ZZN9BrriP7s7JoZ6wGjfoLUmcszb4V6pzOJTAqGGhYz5JtSIyRyhxsg8CSyyUX1G
6G2h1qwjaXpniywq/vvUdZ8qW0C6UhrlyDEdIUy0dZIx6H6A3xWC/dnu6XMqsaGqWYe0JwQ6Rl6L
tWvnsh7PvawdPYzetI1rBN+Tx7b6mAU0pIUEjr0oxNDS+hL4Qb73IZ9UGewsIflVLcnBVZZPdkQ5
O2B0nxbz+wokTiS05JSQuJpqu8xc10GIM75WoKGZEeacGkSrL3ULqzIAsCzTTrxPU1HWtiC5MMBY
obA2x6asBgc7Rb4trxQC9U7qXaxvpaXfphF7qeaPJRZth/jYUIhYOfuZwG8IBeqBFK6P0/WGGFWX
L5cMhRElwTNam7hurb7j7It3Hw7PXw9bzx9YbXIQYMm0BpqtUdBm8k6xJ1rbvZNX3nHSiGH/6uZ6
3w2gwoKsX0RxEWUlqZIPxtns4vg791PE4IafBggMuYHQr7CDlTxaj+VZsDJYXnqh4HGYTe0Njhzp
fxwJAJMdCGihL8jSCnw9+a4YWkyox9M40jP6fBKDCvVyEY4fVhLYAyyFBsA8NjtvugMarpy5nwry
kBO6oOSIzZgZ7FPPvzUTq2YwL+IctvwU70pGjoBJuPV1zYO05eAZ5j/88VVCLnfD9AbzV45w5pLc
3XX5XIvpcXH+yqTzZ34PnjeLECqLm7FiRN4RGtilNz7YauBRa7axKbQDM2UI0u6LR8myIa4SdKJR
+7zdAYjFnfK2eUEa3qtJtL8+W826ShueNfdgg07xXYuUhKI7+W1lA4S5GAq7mC+VGW37JBWiTgKZ
XFErYGPoaiSj+hpVq+jGEJgFsEuqP4/C1O6lXck6VqgBcT2rFirZvSLJC59uOdKegZ157k4Kd6ak
TyZkyIsxE1jfn/LAhvyoIV6zJI5h5zOxI6ERT3p3NRjvxVvIgHeTFx+Q1mkuKTniBtAk6UHxSfXa
eAru8la0rn+HA+E8co8Ey6bcz3j8JEzrV2fAHK8Wlmd18zcK94HSCqqYjt8man29nC+56LpB8J7i
uIGr7N9JXimbexhTxVsRGjcohBXGU6L3OO+VDULj7TMsYnyrtuXMv6j8yXwXr0DBdTFrjUDGC6fH
nQX3pB5d8OjO6bcGFeuAiuti58mwONZAKl7Kdaajb/KyuKUyD7lTKm8ILRYvkbKDPd5YtVQc3cHb
g2uPt/CfmY41ylgq5CqQLbBTQ3lBiX7KSlTgMU3xjDRO/fYZwHmus7EM67l5iveY+qvDohyBN5f/
HaX21WzpAC14qE1NXZyVw8ll+pZs30ineShUK1QtNRx0u9oa7oAQuKKIPGICVOObQ1rAM0R9NFAj
uMwfNIUmoaLTj3dTJyEbyUhrIMAM3PHM7RqbhYHb+MFdmOdjPYrkWNSNwLHBhusy7/Lnwre1l2HV
IcctAKHde7vF4TIma7ztAiSpMSmYPgFU5sT52gu0i7PGOP+zxobBzL56je+UjciVjEZbch2FOiKT
02dFek5mtscCzj3ePedyqTokl9HiYK5C1YSsDbk/stzPSmMvoyPPxIbsjYs+I8IWMwp9piGLavn+
I7AuwdpX/XUnHEEOnOpfk+ROXVlkIc1JyeiulxmVHLpeQidM1gAPumyW+BoRH1rJ4zu3q2SK0xpM
DIUCnqHJk/aYRFNGTuDlNVB6iWh3ODz7QvAXKrk5pWyS8uZJv9z48nD6iZvDObRIlFJXNNH1g5+u
UE0hnaKxQT1bmmzol9ZA3RhRGYmodhsdC8SCMEuzyLNQtYyHXWO7htkN75mDzaMOLZYCEo7/l6Aa
Nlne6l45+zRW3d/anJkHLgzukzmlbpEcoeXYNfOs0zUx2SkaQttUnxq2aOv5pCPOo9ndrOlDKEZy
z0+BvYbKG5xuToBDDaMyDppO+uctesjhy2DLoZHSqnEtdcwAbTlmXWb4j+9Z41IQouJLGYydVarB
5C+i6pNbawRjD+Gk2VenQ2272ugvI6NbRc7utxo1LVOd9qWfdC5Z83LZXn5qNl6O9sYK6l7cWYSm
RluS19BpDVLD419WAk+/qiCY5LfO4eWY/yAef4Cl7Y1ezFom/RzdQB1vh1vkxdX7F9jHcahXnTHx
85Q+2g4+pzzyrHJV6qry/E6cNhlyWuNOqJ7pj9u6FoVzzgpo/R4vDlQmbhKhnhPG/grHdNAei4TJ
H1Gm9MdGM1SsKdnlui7+/TfvwAB4rWRCbIWEXdOho5S9Bn91n8mvB09NJGV/kSyImrE4pMDeSx9y
pdcG0JrIkFmQngdYjQwua28N+/g4U2sWpWglValRAYQXUupS/Q1dvWc+vTq9hMNul8JJ2WtDuaB4
dYc1wITz79WwATeqo20h0gDTbAAPz9ODMxbZIzvfBoP5Y7rx1iUCRZu2rdNLOxeVCetecAKsdw+6
wes9Be7SjJbT86A3OoGFALYFjSWx9UoeLDcF49dITNZ1Oy4Qes2iFtY+Yac9wDzuI7cKFP21kCc6
tvyiUwidMsa3XrSy1srenFrHMPytCGkrXkLEXik0gNmGCDLpcahkgNyE/J1fllTFuCzSoFzoKqqh
hQAUOMGzTuFcJSv22kD/vkhZnE7vqoiG51ktp5UUfhssJKY2R5SM+Oq/b88qGjQT6xvumVNpUm3k
Jx75fA/UzgcFKg5AZSXaT4oMYUJkjIaas4RG8qRLsLlJvlXuxL57Ar/onkoi4XOvBI+DTymgsLUI
8Di7De+74U6awEnEKdJrm8j05zpgAghnbVjqE42qqmfhVZUX6zbycUZ+qPWezOvxSJ3cBocz3IxF
WOcpKcPaN42BYA+SWOvF3M02qH9KFWLIsM7mywwYUVdppl0xJZcM61YAXakXXQStnNfqn9oipN++
ywAX2yIY0bUj3qPGVN0Fg8+8ZywjKyo7a7Iaju2n9Nt4emkVi3nnlWoyuvXKKozLmnUCGVHif2zr
MHjAsb5FeS5pcI57q+KdkQlMfuhZHEg0/+eCtzJG9gUVB82u+P7EkPMLAMNuRuoYK8QwQKc1pG1J
klFpzq9riI4wSunypjnEXGu6eEDSn9TzrqpkLMHz5vEOZFDX72abUYM42ulQPQFK+KNx/yTL4uEE
AxQ93JGUvfUUjQlm8UZnVupRQw6XkPJLBYRsXK4VNxdOXyqm9VpQ2o5NlcJ4shW4fH958nB1hrxu
vixmSsDA9LkwJP7yAFavBCQkRqqzGyE6+BPw6vfIwVHajZM7FyS3dahu5jk4ZgRsnwkravxEIvS1
XmygAoV8H01Q3u/nh2tnVirJT+0RYtQS5NRD4y31r6VgCK9xNJGbMDOFem/lflirv7C/6G7pj523
dPonmXKPsE0rZeE8oPJk+9CYtFE+5jfb47VPXGdzeKK9NN7/sHgIJ12+Hx9QO/vfLq7lUaTW/CO+
uICPlJT20SmxLPE76TwXDKE/j/PobYd8UPnVoNBlUSztlekc1JxbNql9GDxtR53NkhkmQkt/vE7q
keIYpP7QbccLA/8Tk7KMdk7FpCtJAjx2Z649vY8xTJcbwZYsXpchi1nFL2VZoyAXcUEA81t3TtYc
qja313MNVYmVvk2D7aSA7giaApbSABUOFIk9+bYi2VNs8DzcYhWnzY2GNIqbn5l9jSOYoyyc9zFU
mg7yfu5EYczzV9ndqm1KpCDJV7jsqN4v40IowAyU/8nv942HXgF20T1uLOWQ6MkaF4/VpxXmj/KA
/BKrK/bFEGY9c3UgCD+9qdu10qL+WMetzPc4X/6jbraY25mMUQM292nCEjOHlj4u+UESKVKbuGso
G67afGCQWywrA32oumQZWKoStcGpM0h5YqxMD0DldVUetpEO+oFuZR+maZoTAH9zUgOM+IMqX/S7
NG8P3tRlbJWSg0W9OD+tvxky/8+fuzxoQ9yCuNiIRW4QoDgamkjI0OY8zoAI8cQOM8o+qH8mKgNk
V5knHCvQXDZSdUesz0V8UI3owUaC8O3CcnJUTM4YG/1YZW7VxwKp6m8R4CzT5+EgGFf6EBrDEXwo
h1zTApP4r6q/x68koYN1S1zQJcUQc9SXDBjvKz74In2DXmiqx8tr19D3YWRdpp0NBPLUC+XeTMWC
vRyfJq1yZF7zfK92wFzlMKlh/ze2NbuGMmgyRe9E0gTCiq1tXj8S1HF5bSs0FsVaPzwFHFS8JgT2
wHukPdGSuIRyydmg9aqQ9ZXsrw1ls2bHhwC6MrnGKLcer3bS0SymbqKe9u+a80RgLO4CLm0VLbzN
hQkJSm68nf5s9jYr7WBitgm4JMnvd4choNtHpagIG6kn+QCoTSiChH+NyYRPU52lFcQscUIlm3OJ
CvrUht4Pz/TomGJjqXKhDb6hdtGk629VDBVWUkfdj50biTJvAJKl9SUrCf2fjpfeiVt1I0PQemOr
T6z/GiwxT5MYtqHLA6UMeVsOJ3KNhh0FijEaT9eNSJRzXaUBQwUpyzk3bJoMgCk49cp9fo1+xgu9
RWG4ekucbSh09FlI9gmzt0UTOgfpnmCg8Ud257J137sRl/gnkJy7VgqY9Adi41bwJGfYw2c+oHun
sL2SWYNYdBK70T5S7tV2pKKEmkBg6hE4n3afJdSbogYRwbEb7a9uPYL49jXrJipFPXeR1UURqG7g
s+k/ukNU3je29WiPinRYheB9h99UclCdYdjZBLhbuGII6ddMSreirJU1t99me3iuBvM/0pEri5hM
e2zHitHQeOr4UNe5VSc4Zrnubmuc9tSnmdTSLuO3a7OISGxEXmhLLbc5EEBv/bNth0yBmafO9UF7
IX3c3+fMSabqruukNsUZxkF5kWGjzWCjOQgjUmwyUbtMb1gHmk9u8relqtjOYi6mJguf5bSFuy5R
5Yqm1Q8ARliftswrkhDJkm2nA1J612nTfeO8Q4gI44PV9AHjuP4NbogIGWVG/RQTbx1MyGDlXBKk
HZU4lHZ0hNFaRYCtXzglAvA2BxUnLwCzqhfIYSG0kXXXGLlh52NgW+/pxEhXkSyQ983vGl+OcB4U
N85zxE+Uk9zg3mRgNxDCYr9JXVsfj7hHTx3roRhUZU9g4j/1tB8DpoXHoQ5+k/Wmo4Q4gX8FK2kI
RBEh0ShmUb+sd9JDAxpMXzs1ihJmsM9zlQJoDf9QRcklRtadNqfyG8Icjb5i7/a0VmHysiW16huu
b7TLLnCoO1Rsjaw/f02WopkCDHxbLSY1iVc7Fh3yIrXuQkNKNeSU1OECUHPWkz7u05YU5xZYqb4L
TLdbrymDvIvtYbSsYvVd6wvkIvkB3kUQh1btScn2e9n2glACj7Kp1R++LIGtaM/7S1/4vCqa9lbG
mPyWJOU1M5ko09iPF/MZeBpEdxvkAsWBW7SSgxYG7SsDXQT3BtjtnB97tAooWxyNmbVXvN6R1Sqk
oAnckeuleHqD9cyZf3wAYLIs6gxpK070K71AJnvZAmzkgubgYUpw0FV8Y7iZl+Gm14RvPJVOUYMo
jUjKfoEnxoJWLPyI6bdH17jrUW0xSzUW1HphcSWpXv+4d+xgfwuNZ2XXkvGgw2WqJvH8ZGf45a2g
IaZ/kb+RqpNZt3s5EN9yBTyJeVR/F0kGdmP7h3jgmycJf2uNRcAMfrGol6PjJjv4b+kiTvT8o9YK
RfUY9DvFOiu0rw1Jg6D41ZzYlJcdl6EmhIaJqCzRF+J+vIzOp4wxbTPz7TJ3Wgl23DEmvToZq2bB
xOWSIPW5nvciEGhXkH8Flq/tnIrbDQA/Z03dSnoNAelknKsBMepdtMHpNr35KaFeNohA61JVm1MQ
9rlkV28K23qxHykL9+8o40tJCM6nkVDPbYgFWb1GQeHzHmdN30H/CkcFKTZNJxZVYaoL/Jdr9MrC
aOFDMvxNg6igZz3M/YgJagzFw5psgYNrAP9z+DsLjrrfzAHKQPJiu3FU5t/OxEMVUEUW9OTYXbh0
8Ap6OTa2ymTmaHy/oxmCbgZ0xiVsJfs7v1r1/ksvVzRJO7+ZXc6Y2t9OhPWKiP4SpNcAMcEhvjpy
dTGolNL1FgWCFHSziqrvMZFJ+O9rVFJXk9/vvv497DozMtYUVVTVc0ioKpnGb2pWdFctqtVjgQE8
iC1dlkwpbHIPDJwleFLrdgqsxfEgAvLbpAudxCej18w0vtlLVr5MzGr0m1MzMUfg6aXolxgw2zT2
/MN5M3N3VDhsHFBOvUSRcdecDS+CYiOcdxIcBAIhzK5poKM2rUFP15OcBVMKezE5CoQUy6hLRlM9
ZLjfWQdNkNVn2/R5k9H6khdB39Iujl2GBk8rETiS0NPb/L/0tYmwbmBnwI1UniQB19SYo4QP7dj8
cIDLFB3HXxSZcECkQhPajLaG6FaUH2nmu79cll+R/NSEMshVOaP7jmnBtYGAe3Eyoy/ozcdva2BG
jDpJibJvz/Kke7W3S9EMkGVy86F8JVP2oIiXgLnjNbYruhY3F2Ae5sl0ELU4S24jomjKBSga4aKA
Rsp+NpwT733DRDX8GBTKsF35OyJvKVza7qIZR+uSwi5uvCn/SoGy5sum7ZcEM6vqrLt4zpTMd320
qS9n1XNxDCRlPthVVQBq0ZEwiY9OR3+dcIkQiivF1pUUkc4KTsgJhfyUPhwGmq/m80lqND/Rtgu+
noVPI6u+bvJPS7nzcFzW7jzIvlTtQR8CaNSzC6/evaXxkbO9fg7cWj8D3nCqebtQ/fpjPTGSuuBU
CWPOY5e0sHJx79YzuJzBTg8RYOnxbzTCCxb7opn95EmeyKH/xC4qpZvtt1nhzzErHa3o3Hw8Xxnq
lAJdum30+e7VbhNYr5Jl/Ppv9jrXNmPG0RGGy2+HXX5j73cLkAGeD/0vnt6MzkZZdRk0QfCvJCa6
/hZh3k1xib1DdpR2lPegYl/45RM3t7kib54w/63ghPc6JILDd7see0m9LaJmnuyQ1q0TJzIG/yfi
zoT4Y1jbWRebWRZIaPjjzZTPTbMIS7aAWbFGV+LqHJz2O9Soq1ci+Pn6YlbV3lKtQ1RS99UYoKLI
IHNucMbECcG37X8oJnUHZQb4cnDOCqBsxgywVv/COrHCU/ZTtY0aLvQW0HlcFxamnrs1vouxGe0n
VVX33U597O0LhcCqZEC6CMbEfL5yxkT+qFr7ypctcP0+3OJ8dv5XoAQPTWt/7bMeNVKyM1+coyYC
HQyGcX7pA+IxwMFc2Bz/Y5AQvz6WCSPBIC+dtkKJOgtYnrLhRdvIuX7laW/RZ8uR27llJUIeWLvH
GwH366Rdqe9Y12HAcbhUPPyJXFjIdcQ9UGp2Ma0RUl/OGYEb7eZSg+pMQfEYFbEDm7d4/Oggpum8
HYwMs92vPLMngP9p8aGYx5Guop23pKFDV+c9cOMN0vWoEeVj1oFc45+gIyjI4neWvflPbgjvGpvp
yRU36P4F6/dSeuyHSF0iWufasPxj02M+aOJhZXQcklJszv5tPw0eF+WNv5wK+GlRnnlm0VVxTwJH
NqoKfPK/YsGF6iWVvbeuegHmFWZAOUdkt7bkOvkARdHHP3wva7kv/ZO6uOj5AIfNqBYvnRQhA/aB
oBu9enQKLLv6KKhKArJ/0FdU01c9vtJJzSNWmGYk5ue93RH93stXvzDaV4gXa5mD7OHzznk3p1Qc
BgBT55nDQKA07gytLQJFFgKxrd2rKPfJ55is50vWsGuYRQelZcM/ETC8I39nhmxYjNia4ISETqIo
wei9NKnZr+pLJSWOnUTdncxj4uXIP2oNngyuxD7mAKU7LUK9GJyKsOvF8KTkUuEPZs84hKac5Ox7
UIldtsiBfzo6cH/Bxc19UHG8pcHtQwI3FIEqzT7lvGN9i1D4OBvXuiEPtKLz9M1La66UWc+0ielk
+HcBhfVbmF5BrP7xZ3Slf2R7y5OzyO7IRbnE30vWtCjqaopDmHsB/tJBS+9eEBCLuZCfHPO8amYO
futmy8hcqXaNu56BnE1X97ppm5ak7RiK0ByO6y8REimoyGr5UD5KtvoYLVb8lu5gFm9lIuKpWrM5
QU0YHaQF8MYcUn8u2IAC343kJxjhehgbKuXUx3qyDXktc6609UkTaNE5HtFLk0IQSoE6HwveTc3d
odYAF2P2djWplm49e9Vng/pOmIldYrvk8SyZuVDzM6XIM7ED4cgTA4D4BeqIkMNcJ99rjzV6/4US
Mc8PWkSukpzM0aDPAMO6qimPkDBj8b4MN8yLrTvWtMU2JsLkqHFCBdXoqGSi8rwbz3WFMcGuS6gY
g6OcS212QGS10S5xR7Fgz51/kp8ShhgHKSZEGw1tji8/IABcfBxqvWuY+6gUi768BqhmVu6Nydif
8eypVr7KMevfhyt1PfwtzQUvTOrmUG9a7n8aRIwBI5rsCDG09fqCdblIeWlYDoAXXLg1dWdHPlp7
NR28j8WgDSexd5j5WSx6ZJQZB7GWgEIR1DQFTPc5lAXqro2yui8DYc83J2WWW+PnPNPWFGpml82u
X4ISu6gyiqq564oUVOUjOwSCRG/G1h2C2AY34SfvS/XqvbJWRaCea9T9MjDkXwej5PbbkEpjyZl3
uJeeHEEuVq3PjW7YjR+sE+DWBVzAmL3K1JYJNGYv4QlAz1kRn8vO8J15Ov/cXts/xgmfPMVFygR9
O0MU+uU1mNoY2hK7HaWiG46tOYXygFsyOmjSZnwpOu4RQzZxCGQkjrApsSIGXH313JszCQLw+8cW
HV7+006gUEGkgEP9DKn7RjQv/78vSXj2d1T8sZMtgdBOEpq2GlEl+8ZPmfaA8hT3AWntkJ8FnOmU
4zx0UMt/wQ3d4LQENSBAXOEnxnWCpc0TdKK8ucrVHelHTQo/168sYrhIbaBcTIp6UBCvfjSNQ93z
h1i6AWnSUJnR0LqaWmSZkP4yAKuEADbyAXF1fe1EVghQuWZREBwDKQVdcDySOwqKU8+8A5JEgDQr
Ak9OMcViQL6io1fTyhDEP9iou7UfTxSjYRMoEUWe5QciibvU04TMJk0C1GKdNWzOy4mjl7gYqr9G
9McVcEeXb//Z3v7bVMPOJbb9WK/rtx8crP+ikAyjY0Zf+u9igNXZkvKPQ6m+DxD37QBH1QuTaZad
WujlH4fncPiuFixFyvAFNizZjz9uXbaDfTZp+ETuEwfJ9tEzYwROKI1MefUdZN4vt7/4m8n3T1rT
16ftBbRLAytson87oQgtlY52EnZF8fgnzQKffF1j/hBcZjhtPRpH8IpN2y3YQKiCQ+YrMUfuH5hu
4SYItPEhAL7pjazj8O1z41OtbMITWi8IUe4RBYULyP6VNNZR/su13sgw7W96X/OoAN/5on4nwye9
0k+I1851WllUaHwBCYpAkN3Z69mZ2XHxAJW0ThbNiV3p5VNpTQ7AGr84+OAy2s6lpizCNlDnp4gJ
O/USlM2NrByZeVLoq1BUGeqQwfeBQOTVrKYHFb3R50hlm8sMwgNpxJQZzOG7/LZtrC2wF7dFW+n4
pC1C2pTq5AcruGM2mAHccZPN6JFMW90zpZSDOk7WRuLhIUMgjD04Cy6DSdXgsGNTZ23UgR6NX1FJ
dgUWr1nuiXwRIkwG9Q++SyGkv8quShm7AxS6YpldqdiU7rBkfZg7X92aWkp3bzCLEYRH2dcwV11R
PXx5V/d9MU4cdXqA1oexmkPybl2FLvYIBDnh2hkpwIMRYB6kpzZtLFR3Ow96hA4DH8MQy2lPoAaH
PnbDmM3zdXu3lX4UTc5pmR0ilcnCIeEfU5FiphglpOhgDVl+if9Ydcrt3JdYIF3ikgmFaYG6T1yE
idv3x26xIirFlpZ2afd9bRTdi4yRvb7tDS+bFW55sC5XZjJDQwcVY2eu+Soa9fsP+ys69xJRr9tC
9DtfRWBhWUGOWUDQmWkbnIj7jvpTte0WEb8wKq7mAo3dqVhBgPoAgqwfwncYI+lt0VaX0sQEYEyW
Bvw5WsYa+LFKP0UTt10MbPlbbUd2SQasPK1VBBLZsdooG+ifKcgMKppLlkJqBXb4PFj+kNYCyb2A
q8CS99rhiapp6Vk16EadlaOpMx8InPnfEbuyCDQbHfAr3dlV7/A+Q61/2at9HXCYh0z3uRejjvvA
hymeXARBehLZSPQq4AgjEGR3lc3za/1PJSb82HqL6I5v6vLEg1OVpayAC8vwJg5vHhyciGKNZJla
7LzPO/aDiZQ5Dwhrry4wOrf/fl0t3su9qJ+9WDrO232aoHRyZb6Aw/jJ7Eo/onTSP/lMQytTcW/3
dZ829Rx9/m0gkuev7jXbffXc8aCPIqCXCLkFERbGa/nEapZfexrXdxdZW5vLES2SW5VnuPZBGzpT
hXSRdcJE0Yv8WrK6S8vKkL8mPyvIBGfBWVkMTSoqyBHkDtaVrBvz1WV/MKwBGwqDg2MJTOG208+e
wSNd3SaofzRu//alWSslmCAQMwnnjmVToGmFOd/FCIDf5HDY99XWLXArOzBJOpptvj281C8VEv83
rJxO0Z1GHfvabIOd7qPICpFTTsfkjKZ31eiB+xfOntKDRnDsvizu6vr0HszWLChQQ6LZd1MiWDod
7nB6fTc8gPwusffZ5rtaM3qVgcresz8p7Gzo96v8swHADKG+x9X8K6gdGvJ5bzn7dPPmEc1HfIlT
+mj9YEHQuJoOyx/fCau6089Z8yNnLMadvfdj7i8h+Oacn1nFeChEZ8J6bUS3Vpmoqkl8iPve/QbI
JWsp6xWiVAyt4sj5OrjokAnbYjkQ6fI6J0BbSrWwofPDuYkXpKHC63moc7Kmc5ftasrncybz31a5
78IhNTpeEm/VqMzcU3eCvkF9ApVv96IwkHWlP4Hi+qwj22cTYUlAP+NIVVBsQTuW+aa+WnOvjbcs
kci/LQprSk5xMiHNk1v1/voz9upUW0D2jD4o4/+32qggLDJfrM3fGZFrOHWGk4yQiaLzQCxphZfi
S7sETgUF6psIDNfIgXqvmAeEpuXD2bSzLB55SzNURhU65DfKxSpHPYSog6q4LoQWVrXoRUI+bAzp
Ax+0Nbphd9LRZu5ERDp0KyqZnv+Q66ntCCHCIjLRx7TTH+NCny2t4BnhOlBjZiPOsEZ2VzNC44OI
GBrnVdf3XguiB8s7GEbxh3mKfWhA2l67XE60GrYRNCVdNgixG9lD24RZiv3gd7fARvuYQddDI9EQ
v9fH3nGmyBEoMCP+r7StVmHQNdYbjf/FTLSxIuQe8q7tRXbHjo5ZyMizMp/Blst+WCMB/40/ylPd
8XP2bPxSkoGMqTzK3oo/ThV9S7VqQ5LZ6OBM5gDQbEjtXSAbcDZacgXGA/L7txmokg4scpFo88JK
EmuoaA6Ufu2e49UxwBAVa7leCKofeptt4E0Z/sjm3279rpajOFjiR61q50TNe3kmZTh0JyfnpTGo
kKJMX/W/pdqkdScwZHOfBmD9EuczaKxT5msmUD9pdE+hAxqH4qou/iMPU/6O9UMXO3tPOydd08mS
+Sa6cwhdFHPtwO3STxPS9/mTB+tMK9j3mSOfSl4+6y4sFysct+Uf5PsEzV5bBd6dwk6tU/3IFDvn
IyArWAjs82cMwJ54Rmlbs+InxaUyK2BCEk7PKrxlBuE1tbCoB2oMVQvn/FBmWbdudZDAFQspHsnT
zUPgADoR3/AlmfKU0x7ry8cuV28nYlXwoEdnR+gItv1yvLKBgl93v8Xg3fgo0cvUOEQmKz6gRU4a
MwDrAIbQh9XpmnpxlHnhYNGQj1c9vJ1bZ4kF/nNf66sz0tNdV0gCtkZDL6aV2cbe2GptK8k0/11Y
KPhBBZR/+LkWtePKIXCpFpLaTnrliwBwp1kMv7I/szZ6lVSKkFrH0oQhoygxVBqxSPqqFl6Hz931
IM0MCQwsRMjyJaQsra+sJCSVux6hQZzDT3FGcpTbOtVheCh0J4JPuboOY/QLWyNF0jXtkPpzSv7z
3BNoXj8euOzASEFW/EByu1OK/CH4hJjOrQYByIWC2wFJH5x1ESH6kTW/5MIBWBigKwARA00DY1j+
+vzWj8yYMD7moI/BeheW1tM9g4i5oL6U2pyfKLakoi8Nhn84NVSxlSdlRnNuirpi453xSQBRPghk
JcvuVGaAhKeakXb8jy+IosT5/PA9I125Gq+y+D0yrEUh1Lm8rG+1S/yYsMFprFioa0dfZm/owj0V
DDosyH93JssZT5RKnLAIHBkrRuzJ0MRVUWO5HgrVTJFK1oJmjL3J1ZPnN96OKg4Qw+7EPR8/LPd1
+r2qtyI/Ngl2pXTyzkw8vAAUM3OaX4UKaoO0fgoWzObHEi9BcMMD5aTJeszE1xGctdLOJv2cnA62
Klz9edPM+SEFM5NFhCrzncnBtDqyWACgv8nyBJKjuDElIftbZELYmVbk6A0LfZ1ZuwNHMep422/y
1NHl868pdDwJiOsdUxxIrVw6TTFHhapKhTwT9hWuTaqqAjbyw5Id2NliuS1iRROeQmIlA79zAIeC
OxJNN0EO3RL3anNVZI6NiCGUw1Wa7y383wD8Coy+WNW+B4rlunHHVVMqdxaZvFckgwDsX+VWVe75
JNyPyV9ZEPLV/RQFaQjjrATxD5TY/zG0lWOZb9hlYwe6Ox9xQGSjISXKI+zB8vdxFfR0O49LX/wb
DKCDIqKxAHKKQKWdRgOpNUOI9vCkIQwAmrNmbDVzI8edeKhynWuq8nhxCcbiLIvTl64aNyCDP+Nj
hzqGiYHk08jt9CU6nn6BnOvrMs46WHTjPA4ZFvcgPbP2AxFU77lW8abFBYY561d6NHFVZ2HxerQl
tWrrSQ6rpibVdkBRjExgZm1knpxluyt3txJ81cy5NW13yKZpx+nsX1Ji3dd+HXSqlZx0+BN+TpzP
EMVVppsGeG/Razl7upm2ZRTgle/yxzhUdnqnL+fa0Fcx5gZ2UjayD27KwCOeoKYPUkgWdkNkEb0A
boKyugWh3L4qHGOdfYMqjVsGoJfheKVhoHbyutBS+3YZ6vgCNWBt/5Ym3ZAEK2fKDKncH+5LLhwI
etIA8TkdVgsjlMSxgL9eJz9XUZtzcutAUk23Sz3Szw0m3QNdtmbRp/fI+p5IbVJBUi3barUAtOBR
JTUlX12Nhprxx6ln6JbDeU/N/lxewPrgpK/o0PJY7LF+aaz+/FUikkpJSsNLuwwMqELEhrO06KKg
ZDvjYDJZoDHIaovm3i/ItFPhXWrDTau+J3jwNI/+OIq6WPkJbK2pRknZq8NyNXErGZqEfNt5v2BI
gU7grbJo5ktIovBz/+lJl9BEjUl9IEGrsG0qX/E3KJ2z9xHaXxRDL4cajiLeeFmIlylVGzX7e2Kg
zHV+hG6zg1UGAH3+0THP09gwq2hJBuc7dqeBj+Ml6sfHtXvpQusz2vW+Z+8RW/bVd9914XT7JKkx
ABr4Z/UY+ffwhoLkWqU/kDcHggRky3RsNFCcWuPt9WB38ejm1j3Hh9ai6Ieo6xYfZsWivAOFKLAV
/vaQXqHPmOuxFRONooMkBeuZ13oTJjFxsGcZxvPWC7s569Oq4boOYCkItUV9cx2Amka0kocCa1Py
ouFPOSKot9v9lj3Fb5OVCzdb6GSUAzX+ZCPT7tgqKfaqycbCWCPZa2UK2m+lOXIRAOSBe9yWeVaz
ddbAnERrfHcgGZ7OqwEKxucxQnRY63mFESPi+OvozqywQMoakTXaNjKO8ja2TNxmvszcEECYbudB
Xqbivn4+S7Mn+4CxtlQVlk1pd8t5fELhNEOPYz1qZgbz+sNSqxO3ezr4yn0fexIzenZ26572Y/t8
8caZsALLsOziB1Qf4huL7wgrL/SHTC5gf1yyttBxKGDeVx3PDsTek3Cw9yJXY2H5Xllpe1NWjF4B
2RESXt/5DW1hp4gxmdDLCovJx/JzznnC4XheKMgI2aSzL4cwTbHibRddo3IIYSGCLCuMd2flWpwH
w8GgqUA9u8OI49tMwJjIX2E5pRuu72cymvU0fsZi0QZ10GEoTa9ugr141KErB024kmlfbIPp3IfH
D/+xh5vUD7BsC/zAJULBYSAodd3Hu0psV23dUxhH5sUzHMLHkt8aVbzR7H0ecYwBhDrFnGwQLfOc
b5ffSZemBEF7LJplgQMVcyPhTxBUddvhMijaHkQxD2dHpdfLIrrI+DazGRx98TFkH6aFtjA1fuYp
LivUlIDdBtwc2SLg7oCJ0DRSRO8p45TOdp+Ap25OJeAkn7tMPJY+DelaiFGxP+0zQbAu3FLLbcE9
6zhnbQgGMjv2UToygNWYl6uNJSZL091KIqXcA7zDEJU+nqXrwm1/OH/WN4KoTJKNi8XNqU43caP/
UfgxitAOJVluvOlzyDigAC6G0UnIUsW0WCqYUtJOFnrGsZRutZJjPnZSCHJxj278bQq0H2GdDsyr
VqmI4p6ZnNiupvuStYyHpRHPLCfIJQQA4YqHi2Hh2lNkQ3lgVCuVcAXXe0bXO0hkkzn5BekPJqOI
yGBA3xKQXED9AJCVlPaXEIBOGEJa8KgeGk79HVxZk1cESGl8YHjZtvBD3Qbp3RfPntJGKMkBZaAN
Yjx+8ZSWyUKKZc/cfVYuCn+Y+d3SPbzo6X7FtrC+SdbMkyZSYjweLmQ0Fo9ugLfWX0dwY3dq97Er
6YdOD4e/OuL9E8pBDX5RxUtIDZj4/b1nm6OqTYgT47MRDdMJYxSYgF6d9Qu8hBHELxLL3gqtulsl
lbY51Ya5ACYATzURFGnXcY+y39zcS6TONgkA66Z9bEKbrpwX7O4zBU0KyT0Hasr39Xj2SIhitX7q
nZjeZAP4/zurkaNbDsPPvlCWf8RvbIkEMSiV5RWQxqDNqV8mOgebWIQwoB64JOFg6AOrCO7cbf0l
a6WSSr0IiEUZf9lw0CeV7r25/jcbzHTWSrPgnJLj5xeUlT7/SdbHgpKPfgHvILeoqEcznuwZ1lk1
Bi5se27uaVMWjtt3oh3RO+8xIFYSV0MOPYfNLbgcMuTdNPMkT5xxxiQbfFQ/3dnuB/GfWTNpW1m6
LwRuZlXBWeO074/U87IGFl4ZRejlBOj8VsX49VDRD1Qx3H7DNFw1GuUIDBIoDul4SLD17C2YQMqj
fgO5F2w1lWOhzNZs2LJGk3mrZbrmflzgw7WeGyhDWnyJHi4vI1cKTiLJ2VD/8kzHEOpwm1qElrb9
oQHOlk1l5W5DzE8VDRTla4maNNH4MJZczEPIyEcAkiCpmnG3owQqQh2+JvME3hIRa63u8y4TFZxy
vcsU9IgoY7Rbo0VNd8HUzb4IdOvb/o6LsA9UmU5wJ67FaFweZhIxaXsbcYMsS4uK+PIExS60Dw+R
hCh94dhjilEhTyNwfKFKe2eOYrY5Hc2sJll8CSD53Hb+vbT/4WL9vTynjIJp4PG/mBrNjJfZg51r
0umSL8qfynwd+03TxgwTj0nwxsrtvoK+dEMg+s2xyGkq/MQbAXj9Grr+xmJ4AFLWuh7yOsoJiCW6
uDR4FbpVpxD2W3AGuvzHKSUKErGIXaZc2X8v0xGyheVBHGfJXhnyv1aIv1NMj9G2yGna3h1tSXoC
sZYPnRq+LwUja4gZ+LzcfPQTBFe5uWw4pP/vdYvCLBetL/GeNXnRfQSoaM6N4/DB7xtAmXCrispr
uqALo5yy2enCACsoVgpqT6BgGBGTI2jQ9TGYf2SxukFBQxei+Iv96Gi68X0Wz6W1+YdefhYmEapR
exQyFd7yan551kbNhtb6KIGyTjIguMlJsXQ0+j6UiZ08kdEQGJewjukw17k7h0dZ0U2iXgJ6Z/ea
VUvO/AFjHlnO2YG8oI9qNuAosfU9oreGWB7RFoxxoPoNRMptiNmVENznHTyXIfm513t1BL8X2xSx
dNiJChB5SQc8ZdPWjYIK6WM+o9J5XSlzOFi8WH/etrliuZHNHUfgM6GUdLi5cDw/s9ZX+gNcKVEq
zU7Y/t90MC6tYLIrLDPkAfW39GcMgpUvinOZG+RleOTAQdiCfQ2JJ5JgLE2tYy2npGhRJx9t56hY
EX4PntyxZQjZgs3hG5t8SBYuj6d5gOG4IioYSoW6N2L5vRP1+lcLKW8dd1+bYc65B8h5HnUmpsCr
2JuFiynIydcxudUZ3JOZu3S4pFzY9YPib0xNTJ5CAGVLpJE8pJXa8p1Jgy9c7V3ga9arvSWisYqt
y7fiZefPoYRwmb/8cTSTy2+FJymDMcXMU4I/+85OF0jARiXD2D81vniBPgSunLeHYWubqiYIgvnF
knMU0EfmuNsoDGC4s2wruV7PjQj8URSRiEfKmo9gN8gXd63m8jvRHdg2sJxCsDwN3d0kfruggLyS
Aj85Luyvv4Vc+7/3oUxMiMGq7rSt8szkNK4bwMx5zFrkVLafT0BKoNMUKTu1SBs8piRkzzCygyA1
MftekL17UVRACetsWUUQzU/Swzq3hbDKKtrnh3xWBpjYLlp+UYGacyIL2xAVtQ+F4E4Oq0a8IsyA
8ltS6/rT7DcDyoH1WNxI2/pQUPyGqreE4HuHs5g6O/VHYm799ZL9u7QsNf31QfJzzzeb6OulWTxE
zga11pJ5ZGinm9r6b3diGc+hFb+WmNJfxcAtxMRIzO8eQMH8Z/iabgFx9pHJC2yKQTkA3FQ459Md
E7SI9vPw3gCTwkawSIkoyspKw8zMCVFjIAmEeo5FwJP/bnKDwqYBtz+cgrRzs/hETVJh3CA98m46
212SwGzvmYNRHtESoVrp7V7U4qDCvkkFkupXipmLvoN+UFOXkbrTB3sax/czJTKKTb4bNey+KV+2
SDmHujTms71BD/leNKlWnw7VaNVwr5cyEAJs8o6o1V/SEx8T7yn1KiLF1g2XIbgIetCE75UnF9AH
GMI9ojmZVgstq5LmXtDjAsJP8NEDeLQPEEqD3GOQJcx2/+aFcioVqzsZgRt0ltsin8NqrTQDwqIn
G24HYIyfF4bX2yxP+sN0MowVr0NUqXhWtljVFOE3pqmtHipTG62p/1AXiCKp/XK874nY7zS1EDKf
zfwdVniBbzt9Zd+czxbWDEe1kqDLEe6Bzpf1N6aaYQi5/YiTv+7p7CXCUtuzOJOofhmzD1PtYHoU
JnXoWz7mL0Lm1yojAoDfTUuWF8NiHEjmwxoyRK1AjjPIdDLMEsuwrp71Tx/uHOqBaO3qomeFktEO
ZkyHoEk71TSUrTEFPsZ68sgqwGUnQ3yb3eB2pczJ7lBTzq2pVt+ahITGCcivFojfLT3DIPLybN04
ERmtt9tl9hClWO9f90BkcSj04uF7WmkpIqe+HN91wTyhx/odwoYWoK+VoVj5sJEk6OrkoTxTPPlN
zKO8K5rl2LBE5BRFMMUjf824ZBgBEwrrgP39XDl1aaeMKdklvCHRxzV4/yAxxhO2KM3TG/YGIXxq
q36qa2K1t1P/Q94xeyseNfcTVRUW7mI2eEeEYZIjE7SqT7+HbZkEpkwJcSe+Lfvb+k51uo263gmw
YzOclNvSA/vSBTIQQA6tYoE4bIBgo198Yf32TwhO8BdyOO5QrQcQkEWtnrl1zJhNuIJDaxJK73J4
tI7Mq++rdN5rKm7ERdPlp8gcjszb82yyRP2tu06PTnIDKa1SZHXVWdHzBWs759HGBK2IfvQXcXBq
JBWzkEvfy/SYI7UQa49Tc51LmuyOrMYf/yjKlXVDSiQH+1ycHfLmcJx5FR3CBA7ZP+qQs1ZVUrry
/rrp5X4uZVA8TXtjlgBSl7QD9Tpi0DZXFU4HwkU/5bVSMHoSi7SnU4iVqYTvAZitCS70DfnT/NQO
+5U4NEb4vRkln7jnrG6wQ3VAEFD7QkKprZ0SNF2Nm9Qwww2JD0IIvlWdN99FZQOJDUybG3XqNnr3
m9HXETPTCudn1hi2Vkhd5hTSqP/GvLJp2h3ovgdoEnCmfcfpW+T6nE2dH/Qa5xvjlF85erBZGLH3
X3F39aYK9qa90EinRLZuZs9mSDE9aiXGx22NiLJLFNK998t/hwWaMh56rNLETdtdhze5HghDomyo
jJnaAB2A0muiB2++et/liByBv//DWpxvAKKO+bcoYz8FEdYJRuQ9skISTXcYv/wvS/dGBOSKzzzI
ffNgcDKqSNz4c7GCC5Rj4lpOBVgzKnKkpxihKwg+vdyxeLd1lpZzi9J5QELcUx9N3VKwNs+KqjhP
S/SRAYncpIobSz5o2++PCYATCZSM/KR3Eiqb6nJBEbtycXi16B7vc8kYeOheCUxY8rppyn48z8hm
rPibhTmp2+LKakKu5b2WQifKkJJmUkTT7tpNEnZ4UUa/7/4gecrJ9Fjoy+x3KKBJyBhA2Q03vUXB
ft/iB6ymsfepqjpIhDfe1TnG9iuWiLXgkj/FbLyJ6hTNYBZs46pioM/vg3SGyjztpIyi6lYkrdnw
Yslw2nFOzPDF7pD3eYPZowkayPD3C0OU6rE65BkNJrOhvo7Y5kkIdpNKJ7foL8RKOC84YFqCrPGQ
6FIiqWdJ6tJUOijeV7+RXuYHua4PFuD2QsHqIi3OExur0cHoBdacGc5ksVFWGwQW+eZ1vD70tO+t
f933De3cB1DNGxksreKqLEcAXAlvdJn778KQEp93uZaVd0HXeRdvi0t1o8kGCdaGvzoJKcbr68vm
K1M2paWhYPq8uBXZoJtz5dYaFFRVxxU/HV6xNKLL8WMUIhMSuDsJwhsUDzihaKbsYRdlYQpZm82I
jroTPykPrmY6AsQQjEkqMf2bulQpVHljYvS5E0w6iDcmDjPTxDjMTAl8Jru55DPGKivbZv9Nw331
hH6pRPWh8dElL2JG75Dauy1h2BLTCgIzaP6y5XMGZEXuuy0TRoxAN+EX9Mani/V4M5xcXmeJKBnV
eOa8akmxTFdF+Q7KM8LfwmNM4PEIwD8QVs+Z9DktndyBPhXkLHPGiVKX1ZU257AqMXvFJBB+DRH4
ed1gb8gXljfs1XWs4ecGJiUueBUFQM5gFhG0GBREtuHDEbfDgI2J7Id/sgtwgtlzi6EaS5Llc0n5
A9gJ4ppOIrtAUOQsI42SkAOemUsRDlre+ZOWpBJf78d6yA7ZcUJcGefsTv1XO6Nu61S0rY+o6TCH
fmMZC84urP/wl4AAfuXm2b+sPyhUWknS56ZpX4SDGEpC0Q9Chchy4LR5LSPSY7U/KlgB0azGFqOe
Agw/5mvToJhkFtzsxX4dNhHiSDznc9Ao1yU4Mzeft1+2y0ZZ2OhoBHZ+UlHpLvnO1vYJ17QnXJDK
H6KY4WOxuGUYrD8E08GkjyVXhxVGeDpt+7DtZKO0qpMtFc2xzQ2hgZeXOm6sg5kvB/X9FpAladJh
SKzYeFYHTp6xHonJX/r0ii4nWi6nSX3TTfAlxOi4s6ZbSUT+eQ4HHqHHWRn5xISfuY7FNVYjUhbU
E9Xg4WFxHZNOOEmpcRuZdtZl6DfEd4q5SkajugE3kDQkacz3lVGtjEaqXiMNj19KXe/dSmvHzQc1
4azPE5qLko+u64upmFtRhgi5t8s1PhwUlitw53cSBIcQ2v7nmeXeFEn5n0hxARgUckI46evF9DMi
WTvFsYMdnJ5z1xh9zdAit5n6OLtpymusvcataa38ja7QBsyLOeMHT1gFzIxHt+x2WK9G1aCSEVWb
6+aPWEe/tAdKJRCn4sNN3GlE6iwS70FrKRtToLUhl9rsmhe0oDCCZQcQ2+4OGhS41UFVEfjORsd2
U1luHG6KC3F+oXVNrxn8bePef3vTUrj0XQXcYfY2EPbMEgeOkz53Min9Xx1RDWKTDtRHz/9bxlOL
hUMd1jvvP5NfOtG6MblybF6T16rYCzdU86NXWtigug/0EH4buFBFFtAJoBSUMY8B8aXh5Wvq1ynH
csw6J4Xp52lS+9qLc9oh/y+DKhFFyMdg/shAy9b1NemRcDyMUdsbVU8G4N8g9FEyAgqxLfnSWxZH
AfK2/iUrkJmVyS24UBKGg64wNNW28dS3zECbNd5Ou5rju3YjUrGJlJjZ1agVIoX+2v+Zw1coYA89
7YJbY8hLz7jhZ0JRO+i00IOemJtvrxjJi2cDYOb+on8K4tLLy0UHlM+JrHZvtSNkVpgylQlKm/VD
arbZuLe0yKt2xNnrN0jrT/Ey/VGyVhQNiTBOaPZgMqraKG5F4F0bc01G1gJg4yMgPJ+jmSaZdv5P
NXecppM++YK9x6ikjsBfF0o90FXL/7WAO9OeZJzZC2Dv1qn0bk5V+Thzrz4dSJgUWffI0oTP8Rui
SzQckMJQnfYwyjDKjxvhyt/Mre0dUKdgqEESt+EhC/yckCLz2IE8JbLI23WMNxN1Jp9QXHaDYPgt
EJJlLNb5XiCnmcHgezB/O1aEMTO8kQhtRiVvDN9cOFC6+Oy6hSErmt+1mqwmuSIQjdQO5eV1mXLc
iH63rqU8nZtAeQVEqtc9Ncy9ZbHwM1SxepvUjYmDz+KIB39l8VMG+Ht1RMSR56SklVCvLWJDQtj9
0Wo5WAQQufp7djksY50ElX9+shzqjA1IODkxJdJs8QbEPBwKWKRLwiK0Mkx5QwnI6yGQjhKKYAg7
njVya/QR7f5Vr/AnXz3kNoMEVt++fj1JtFdM1EGnyn4J4rqKSkMPmHudtVstGesWo/3fr0yjsU9G
oQmDZXGA3vYHGQ82ooy3oHTNe3Q0r8sKhpkLC2XhySX0bzUU4JWgBSpPgXK1+vVnlKzklG1tLbMR
n854pivFquPTkBCg1fttiIhesgdffIRo0hVwZG8QhDEk0iF50t+mCcZ8xMMBoFFVZh9M2Pdk3Wyb
hPQVnZKPsduvsGucmr5q1UCSs7xjcHMU+49cylJNz/wgt+LDNP32aCNsWnpd+m+sjdiS0BD5iGgg
GUWQVUyO53G322F7/fRPs1WH2zZmMVzfX4TUW95KZhohb/GwnE/xMvGx2AyFEb+A6TGBfsuRHATF
eqKcgLjEbaMfHVY0HALkiEJXXQ0+1at7jSsWjqmBaL4sYFiBIyXjF5V/usGmlhBnBHDtxvb2wslL
3vFb/h8+A8YufHNNIRjy61RedfJLiZkvJInCAehWqKa9MZsIseqHi/qAk30vN2s4Eb77U1dLglI6
VKqmAfHyU8lLnMC3epu0Eijctbe6ufW4wYt590ag9FR0UZjXAQc+oXDsWaRMzmLhdJMljDV1qJfr
4ax2JarbgYfChqTDUwaK5Q/4yYl/BJ+NnOHJYOVFgyx6uGY8ePSU258Ejifbkn1U3tzLtDow3ynD
UWTWkfmMk9Q2pRA0b59pOlMDUUdV3nYvYXRBIPTk2LZ8Bi3IhPNc3pr+lg/CSKa2BwUbYQ3I271v
vcVNyAc7G+vXkUkbK1LYDbmPITPgBnLZUErVtP+mwFoA2GvMTAt3MGzLa5npXyl2wPr+CoY/IryU
f1apZ8z7ejojGHCG3MjLK8I0NZwCXENlArX5XKZCqXnwaNqexGneq3cdyyWBi9XGbFjjicFLmkVU
svwB9SAu3aiMTEUi9yxgGjhDNMw+nUROa/e9O+StjLDhjeFv9cqOTrS6dqmosi+exaVx+XmGXj4N
tGTHFpUlGaTKEx9hAUbfm/b2uHdsTicrOqm3gxSpMmH6nObZsAGj0hiWjbUObyjF0d43NhRdZLaN
pwaNp9AfU9FtTWr/1ES/cQBR5P4H+GJv6OzdKjX+Mie+Za4GC9ovN1nbQPWVJ0lA/b44sNIGIU7c
Zu8WiwSmjFKwJgjYfdDXgQ2PaDhEpAmR8JjFvc/rTf+TLKY2XFFqiSmsZCqYXbmaqqJRptOsd7zz
K0yPjwm3aYAdgjYSAJcblqv33CpYu5gxzVLnX96lFqt9QwIF/WwZQJmj1DYYUZJneylfOH9/vq8f
E/9gnBL5XTENtGeIrd4Hxje/90M4VDnLTXPnrVyMlwHovEuA4QR5FaZhF6As9exl57GfdmfY98EJ
SD8StGhRUTYiuWJeS+3jAHrfQQ4N1BL7QqxbynBKUlAdTMkNCAbj5crRGPPkOoZSHcMPJEf0ZbZy
pS0AutfAuCGR+6H0vVeLbO9eBeKt9qBzSRA6svZ+zPSBxG90+UA8y2F9HjmzxkATFXeRGikEl3Ph
TBX319ug+afC+A1K/7uH47kz41TRwxIcpjObuuMV1RfBcrzPLBavkDH9+WgAHEH+5oexRRZlvJna
vf+gfpl+IvZUGTaXnRwHt3MlXuv6mD47sZgI4R4hftygBeMkMwc1SGvl2wQ5LNS+TG2eQsrajcfT
XUsKTko9KRZVP/pEUEh6G3ij0OH4tzCSPtzBLAT2PS1sDo3Y7ZYslJ5gUykD7nSWUdX3E5LR95pa
h9XAQ6dD5ET3aTcghK+RODGdvYYJbMps4bB6V68q/pkMCZa/uw3oPTiN9wwwucfyzSPe17Ea3YtK
YkwKEVv98ILo2U/yPQz5SJ52IjNWOfqnmGqvGSp2rxInQXNAiDl0mGKs9Ia15xNsgpxoqnktBi5V
tHj+GY5YJcABz8+uRaceZ+4CMMIuoZ0GQ4B3j2LsWJT5AnfOgcb9fl12fb4HY7DdXYHXMr562g68
OnDgebXaHGWA2Gy6OeAYHvHX6eKsJOU3ktA85EGjAQ/KwmU0urcIf8eYa9lNIy5A39C7Fkp551d4
6Xzm2eANDOco4TaSvdw452dv2KX2xMueEmGqUS/qv6s1h1szn4fwdkLGf3TODqls95ReRdY7JdRN
zGXY8SAozDxJH9wUYzNUCOfEG8XTR8U/1uIZwcyeOhklrBUMl9eQvQQ+5VjR/NTNI7KjVINPy1rW
Dc+KyFgqV9n0Bs7jzWPh0O00pO0itpdCKxMG8q9rEnrJs7eAmwv0Rc1B3vN7lFDlZgHOlLSgYB38
Xk9jbLpbWlxKOY5aQatklj8WvSHAyTUpdY5VXLvqY7oDZXFwjvhbTZFP3CMNX1M1PuW/mJmu8XT2
5kfZPWGOP+d8rs09xhYZN3s2YuUyAK4elQ3pITtM3HOYI2A/gutGtaSnud86FSNZpFkDmqQEp3RV
6mFfmOzKsI7BdsWkFDHClEAvqeo2QJ76h4TCX+8nqBLH+aLWDOol5/tObcuI7wKRdvMMeUomMzNJ
0ondkyZ40daCwaUhKw+h4QApZraZeZNMWP5cWcbbC2yWObGXPaM5S8LjvskRFg64ZfNuyHdPjEah
rndnEzGZJTe3ERtqIJULFC/TNcYMRyJbLdBAqtOqJ975n4Lx+SZnv5mLqXyf/ZSsSkCxA7EhhdWK
wlUe9Xq2a18NJOhp43cPWWFOhkLEMKzIJQN0YtFvjcUqGHNXb8kKUAi6viMHAZen0sAaJRUQiw3J
QFHAyHt1avyF3OAI7XSm5QImZ30ZcoanYiYkdZgvt4KfvnVb+Vnq0F2K792h7mdLRKSzOsncFpZg
uRxr9LbaAkmbP/Oma93GpfRCPcP1FkgynartA5GNcqeSz6ivmt+PA1prmtNmgBD21uqMNqnPRHiM
mMOe+UTdwAfONewwx+32jzkCeb7oguz9vGmqOKlqOjqUxqgSFYpvv3TREmw8n+LQm0iDIn86WdFD
Bt1ig8+kUiQZJeCevdl5+mnzvzhmgH2IRL4OiNwSOzXwMmHRJ8K4s1vyuI4G5CAX3LJcXvxp0MKs
585qv0WHDZmrgKRDaMJdXGB8aDbBhrqQFuZaF16eUXvJFahsrKEkD+Qldmyn1X7Y/Zck+Qb5HxKD
tZiZSHsBhsFvfatY4C4Red6scAGra9TAzZ3/xnRDZOIz9CeK+Pgiq5UycfRP2SsSEp7Von91e0ZF
CIc6dS51YNH6yxK2AjUFLlPWOB4gtiRX1nMvdNcxwAYFMTikMY8kPyBTlUs8gdI4QqShv6vjMsJn
I7wzAxqLzF3JBdZlxOIu+bj6K013XbqpD6Mxvh3NAN0p9yh1CTDnXVYcTST6Fs8DScbAYgFPsDTm
LjD166XzAAGYjIMwBmVSZkXsq5VQmciq5k7nCp/ZQRnPJrdBpYpYCikO/AA78PB8yASVsoapI826
o2mz+NFXR0yxmmgLonZI7GNsaVD3E+4OdwBlITJXr4FAzLup2//e1qULjZSpVztiQYxc0+ybFo0s
XmZHBWTYaLSgFFiVh4oVyCAafeMDPnoMBGWNlF1zXMBWrZFvQ+kvvMsjo3QLr/J+RLbqm94ZbWLX
+h/W/1oZkvvrXQcbgkd7FHBwAUfev4O+MuwvE/lddPqjD1IchZW3U+MIOSYdrYE2kULyFTcXujN+
BBOVh16mRDEGCYAZFUC72r4AAiXDGMPlz/3jRzMCgzHPxOQDAYGBbeZSaFUpDkbxpRG65Ztu5Z57
p5udmMw1WxEbbdR0iAGXIyavS1n1064ObY2+18qxjK5RNF7vj1p6saE6s8F/oOQ+cAapkqy3Nf+h
1Q1XHWHA9gYkXB2XqnmGJj92xYGKsukVbDU5holG0fZfXAR281eGMGaxioNcf+0g50TWFa9iQyhL
yP92cAdn8YLieL+N8iVOSPxqjul7yhkshWU+Y4op3oaoOz17dtk2e55q+Y97J8HBrhnrs8XNSduT
sRL5kLIUVoqQc1lJav7Pl2rVb9vD/0esbPP63O8DSVvegq+9rNt6yv0/+BW3bN0oIXin00Za2b1v
HiAuydcfKB6pP5ig6JstxbfIsy1H7vvApEY48j2oFAxmKGzUhd7ZbxA21z33QtG5E9V6QzKaBgey
o+niV9H5++MkCTC3SWK77IFf5MF6fLOUAfC/p1YMGJsOkTmJpx++AA1jqpdu7TSsWCqiTSt2CQFZ
URQk9Ck6bsFYoQvyXSEeak6p0jt7QBa/r/E8xemPvE+xtnJZuVUyMIAN3FhwFbgsJqJPBDpe/IL1
yDAsf8bYU78dLvLtj8RDArR0wK94Ym4ii349+VyWrvcvtlGbXGtl2avgdtNAMKM8T0KGqzxrH72Y
L6FXYlgzlIs+IA+gWsGnRGXHRnYewvATPzgPeIPdeGtREXTUip2a4TIUmh5JdvJHsQlVbSjBvv99
IQeVzcsntzSbhL7sPWNaqdai040TfnWlFBtwn6CEPxvNQhuumMmhWbM+Z1j5a+6h2n9BPb85iGqG
wReJqtMAG1UjvdQFjBdrG4qrCsJ29FHL1QRcWwPC2T8ixLu3Tsnpq+/ABnkQ5AHLfjUCpdAPDbio
vAFh8a2nJbGXLtvXfMr/3qJGp06izEEhRtKBDqY5lo0/w3kTZXZ5lAN6nzyKmp4Njmk5MzVFakWF
seNpAc4NCsnlEjh28qjRNUPAi15/FUs26i8b05bbDPfKJpxoFFiVlkXSL5PRJ1j2b3/zjn2IE+TD
loaGf4uOnqdm0eVyYLwk1Ac+NfH73VBZSVmq6MFkCJLAl0BZU0I7KEoJkB0/z76zaUR4goRIVQ/J
A+d9cZn/FId4Ni787R7gJ/AIgoAxSVGNhCVieXJe9KVrYJffE8zlEipYgqpmWuyIkCjnudC206SF
7yWiCtltwDaGnikYJRfLVUfup/+EBlWom7icDLJcaBTtFGoPjgpATeTQh8O5j9UAWRUXYnrWt2U7
+C1daDL7hV5vR+MrC81b/v6Fa4Rg4ckj5mFVCGD/iV/YKuFIYtkMIlD8F6pZtCiJwWBmsm8DjI6P
sz8VKwv+rA/7BUcFrMj+cVlBJwYFv4hDzC8kXdHcemEN47r5a5WupOP6gtm7Bb9JqQieDNUtmVuQ
+Inj+PJNREwZE10ErDfkvQ/gcFCcG0vMSqiyikB4wQXmw+SP0JjNwbwPIQ56/7MYqO9Kopi5wxXy
ghmhAnK6b51qafucXrP02B+WVhwOECKCxHHxotA2kPGXPUyjIfocm/7rQRWfOwVt40aYzP/d/L5f
4/PntacKNzPJVRRIMSxf7EkUByQ3JqCePtqjgAaZBUTGS2szXrQ5u4emKDenBpOh3uUGE8KzW25M
pf1yT+EScthMcPUYOMVsjrz/M67bBdoS3aeaeHq2bx+jRdKwHW+2UdRBMZXHgVq+JVJNDFI6xJ26
g5Vi1dr1KIiK3uB2IJQL97uXwzytG5rh+acPIYqk47TfDhIUacmk6kv1CdpzFmyWUaaN3Li/pSfZ
088+cV+rkk28aG3GMlTAhwaIRoyy+jXFIeO/Zw70taCxmPJFkgmsRCBgqSMdmnivX1YJbHRJXwxN
9/GUQ4q/3fuQzLE8rnLAqU7OzXmuDGy/FZZV4pmFosWdTZBloHlmA3tsp1WtpcVawpS5GFpd0oK4
I56Z5gTOdK1G1IEkOgPhoF8eb+cl2/DfvPG6Ti/jnynsYxfEnRcOgtJ+VhC9nu9j6/6W4GbHSTMN
ylrotbXBAalxcbbeaHDnCn3pwvLhmUctydcfPDDN1H7dmuNTvdtViwWpeltV6LJY0wSTKSmX1nqS
l/ziE299nZoJQS17Z+GHkYDtb1ZfmQa8+3haWS60Rg1RmFc1HUFF8C9sTknpP+iIn/OErIlvdfSH
zH72afzQ2HdckHSRz4iFxr5Irve0zndX7HWdGXlgoZo6Vwf12mT8UhATIZBnR7D9BWhLxxHf24mT
lBfs80U0e1pXOOJUwL5hTXEevEYLhd073zh2pdEisieu7UMCGZSxl6MPmuL511E/1kWMxP6RBsNA
4dmOilTC8LKBZes3jFDbwLSx0J1aDsA8cuM1n4lliTQxYaHTDvNfLJSge5L6x8rbz3UTSYPu6ukh
ctupxJR1hYexeP81VR1uZk8W93OpPkLMBmYQyS1wOEB/c09yPfulM2OdDQ/+y5DAU+/+idqs5IC8
Qt1GtIpKhCzbcTMbtFnjanA28VMFYd+c3Vout4nELCJjOjZRMZEEmOfzNc7K9GcGm8IGc5EpXX4n
tsQfvw7aOSHQAwgQarQfj/v42576/8qrEy2NK/OzdwyrXc3yK63HZHwj2pQSVTFf9GaymUwU5CCj
EuMMryLDnakKF1T22Sz9tXRuuQuUTJsFWNx2tVibtVDS8dWaHZDuggCVvHwRqTtFJJVv3adVXACb
A30rh7nImb36HZsORRMn+xtRsCF64+o6AHHR9+d8PkQi60FZzJNoemcGalQBDjcYzud6WYds+/6t
mpNSa0GMfIOs0eCBQhcHS6FqnSaCEwhpgdhauXuQ/QxecaUQqwqPItEqD03B+dnqY0rmaos3ONW0
EsioYIXrGBMBLFIHYsnSMpEfLhnOOMQ1lapL8RvAopfgcBVGQD8vlG3mr9mUr0sM6uNbzhwPzQbB
kJyfvDH9shzDC6BU7UN9Drg0Kg+Kyvb0QB3rCedTf/myWRUugWHt7v2pWxQGjk+chcc91xqnXtYD
62MUZZDHDl7THdw6VkmC4IepONXyg9Y60YF0cmY3+60iT7R9fJWXH3WG4XDGGM6+tEbQJ0EvMl9s
/gdE13kaOOAI+yfgNwNITdX2ZdZwyo0FgJXxXEVRYLJjfN0vFqN2gGgmGE8mdg+5DVvCLJyjJeRG
U15IPwZcL3SjyMwxbO0J0f9LMqmVhlNF79CB6zMJk9XNjKEz9+C9q7YvLsIg6yqHxiII6IPs0vIo
x774TZdkzoisIwCrbXLobOeduEmiwT4r5rlbEdxvwcWRVbbY7vnT77vS9oaYTPdMUwiI41HzfM8N
UmqTH6jrNgshVlZw0CxQD/hXrC2Xv/Cmx4zKUtpkVtkqhnc3/Ste0SozKehmJst6mNp9adQPbmWu
XcGduoDNw40MIdDr77ZA8EFIbNfyQus7UAhjL6P8VeAMCg7ymWl1FvghOZfnHYhCrOfPMAEU0/Vf
27pj8fTmFzWw35FiO/XloiXbe6e+vuLkjWSGFHaEpuDE+ELbKDBZzRuSLGOkl/XNZ5AoZQ61fW6O
HYwwuKV+Q4eN5CEsNUydRH6kjy7zxOlyaKngwCYjMPvDWFr/zlJwf7p68Tz71xk+PXaIoZT8dBK3
6YfNgLZ7fIvMfDyEkWSe0/r6HQzZpoWb/tLrutmlgShOn3Fo3ddDE3ECDO7RaZJrnSGvKz8ssmtd
HzRCy4MCtLKPyotN6LAp35rRHIbCWYLNSbNHQyCPbAwPRJC7K5ZJF6LAAsajQA2bX0S3JMF1duix
59h1fUtSnBk2xyVQ/6222jBSI/K3yqJlWlW9seZV32gqMgcfJjbHYNuZZDODMHcWw7IQ6zmTeWX4
tfiXHNbieBexS3HDNFqVtp0EFmbFcLGDCJcDQ+bVkiDhDeQCgo3aeslS+7/fh+XQ3ce7Px/CMC67
CUmAHtmlWGIGebNcpjPq3AO2j+bRMxjVHJ4rayzzDzj8NV5/J+xShOKDJ2PVeuXwoJpTl5u+YzyG
0f25ZInl9/L2J5H99x6Xx35vAVFcVVCJGwrA+6GjI+BRP/JNLo1phiJbQ7dgwuwk9uVQfbwdwHr6
nHWTTR8QudwJSrS7BEx1HsXX/um/N7dhtm36s+0t9T7w0LBaK/azewZANS2a+Q0V3HeaDn7e8zzx
2aFQHNvRNc06xYaYm+CfxnHMPcbrjM7WVoWCxL3/1+bfPX6iEIQlgVMIhI6nhVb8r0SwNrlyVpIu
VkJRwjdh0Ysaj2yCNHw7t2zUiHGuJ/UikJ/Et3ysSb1WDXiCyblHivxQ1C1BuKZMesDzA4+I6FWe
EWYPK6zkbSaSqOvNCRGIbKL5x/amOpHR9FW8Hc/Eud4c+eoAqT9w2e67+nn93gP/szAJp3E3v4Bv
HI5zz3IL14eFb2j6QgbHmfro74caMdbfeDk5wgK9RIUvZD88ZJDmWyk+HaxKXnrzfr7eFKGuTFR9
AoZnaU9+wGvXfDoPTdfrTBqY/SdN02TVfcSW5uJHPxuy4DWaCs5rZPArogVpZ3sSSxYaMaahyfI9
YzfKQ1ERnJdyolSnoM16Mwfuj8bQd9cuKLu52IuAR7XToSxfLyFadFGsVZM4xpcILymIRtLJLmHX
KyT31CqXGlvJ94ItS4YtgZgCH4exbtib+uCfDUb1yB7Y4RQ9RUpG1aDaMM0EDWfzP1pOfaecvVFi
4Pf4Dtp3h5fyKgmlN/9cWUxBUdjZ/PUyghdGhwvKNHeqyIxNv14uml8hmg/J58W6xu4yLSJxSuDe
Emygp+xiExzS2vzYhRVVIzreIAslCSd7K/7drbqxsqF03c29Ka0e8ZQPysLmdevN2IpbO/qIaPxt
UwxzuRT/aWnAnSBARA/FIzs2O8yNeeVjdjSgGZFBAOI0eRcte3k33aSbGtcwdtJ8tiS0Np78rPP8
S7eEUu5SSM9QxQ9wsBNRZNcehL5sOU+NAMDhjELFIc2cf9kAs0qLZZVG4vAUdZXDrDe7ynlff/9H
Y6gypRUmqY1gnww4XNWXbDzAxMwpBEvTyaJmfezogkWB14j6v6fSbHD4sBjBs5ywdvVulgJLlyPd
DFzAlw2xpaOdJM9qJAsIh45CSWmIlbACgrJIMZ8eLyhlV1XrGdQGw9btvMipa5pSy/oNjgTzVjex
SXNAx188EozVOR0W849HF6/4X95snhI6ClyoURtplYDp1cvWNkgmkZ7KT1/rhIZHcaJXvxZPJXWp
2f/lud7xhzUCDC2crnQxGz1tdHKl5BOywch2hujc1xcLmXJ8HvcoDHY6MBvkFfzQzA8cmwNJlyWN
puTI/TLi1lV7HNmZshUIKvr2InQhwh1NWVB4TzVaiJJDHZMVBtbUMMBKNuW6SnhzYZTRhIA7MrK/
2SLHqQXKb74kN7r0Y23woBbAs0EG04DN69DNmmT9/YpQbp/Tz/uLJZg3wcUTMjSBrbp7+oQKcupO
cz6Wg9p6JvskHsywWJsAtQHb1DYPzgpX2DBgQzmmbp11ruJxWZuykfZ80SWW8zlxVb3gy8K974AM
fEwEEdL84C1wV6JF7bwkcuMBu9DsFmRgDzTrX0QhVzvSvllKhlSuhaT2EyDYJ+Su4qAfTvZSYeNu
nqmT281MAZCBRzYI+ub30+7o+/gqCr+icmgnvdHgjpZLyX+KJvBhuMQ/YNSTkhYiH5Y7mFZ3fbnI
JRIJQKZ9quOdm1KIsvxYISC0cqm6t2REQ03IE9JNqpMbzqetJmCVeh8ynZ5CXT0KY1+65ok7iWZl
rrr5Oov62EeveWm85XUzcWayi0c4qi2ZrSE//UER63cAiA1M8c+Ji68iAhXvBwXqHbVewDSOiKKX
/ETBUQ0QbdQonRhZbvK+YPsRCHX8L6FDD/p9dQm3/lYkVCRqyfbtBxRpihzb3TguZBZ0pUe2iQL9
mvjluxTNvxnA99RdKpWNtvMLyC2pQRgMdPmsGp8GgKEqsI9TnCb/CtvVv2zuS3jU7zeV6oPJxsB6
R2vFMmhLI200zvMNS7I85oEuHuCNuIK5aepH7SXJ9G7Qr+c0GHWLxaoPw2cTkWcCMBtHv8K00jpc
EmkyceaHI1cQqCCg+aibUsRXqCIU5PGWpdzHTxHk75uR76fIDC9gs163oRp6OP6+/7Gwloy7irVL
C8ozmmhSCqJEPHvajvlo5KXlqUDCoJ9vyvXgDPOrRyUDl7IGif20g3evcvegoU/1gBZMrxpQYDis
o52zI03IVF6jV2BoAY2RCKebsDSvofcnZDTVouQ1k81CukCk1OnCeccm0mAHwKV7EjPLMiJbzswl
F8EAU+QkBe5NjwEjf39sb5X8yPGtljNZUSzgzCBfRbGBtBkLQRQlYXcJSYlxvXtBTqAzUlyPMIxb
g9mLKJFKNdMMCRC7IlXNyNmsYVGMNYI1JdVM1tFAuKV/1EdlTyXtez4lG4Hu3IJ9dmjgRVZo6fki
vo0v0UaXX+QAbtdMN9F9VoFwotCUUqrROPNvug74rIbKWXQJ4M7qTuxr9xkvh2XH3dHpu10uWwFx
RcflvgQym83lU0Iy8VoNLWNfoJTve+Nk7NI0NBVr6c9YfC+aCI3CAVkXq4Jsfq1y8y/haJzIaMk6
hh/J5rEUkv4r4pDwUtt/S+YkD6bh3LF/aWKKeWA+VizzOqZxbaHK/DIRWezspQxbnc7aneU3u+yW
r/mV+1xow99L4h89aExCWtWSzT3lTTfqj6JPohZHj5l3bL8OvfnADMTj51zFH+ObI333R5Y/lMSl
gB7R+TQjo1SelpjN2Tho89oEjNAnu8w9ObwR6LFOfKmfnoOGF3YadsUpwyggnnvFENnBL6gmKSEp
JodAvjjgFJg90UPTmRZz8r/8wXzqSwtPqd1YlFwf6JMByTMKokFDkDl5JQoK874OvA1BiysJbrdD
QvTk+LihIHtaGFWWWUY/4jM+pRbhTOXjJ49xhX0WLgnpxdtgg4gYo4NGndz+qXPweNftblFnCa78
odGst965PXHhpM+8OagRKUVhtYQay6hK+z3gngpzeY6RhgWlWh9M/LxpX0pjN5aQ/hpu39LBGwoo
XSWpD6rqspvlKVm9ZHyhSoSIZBwVWT2k9JmvSx5BLC989BaF3MJEW94bsfApWaZxSyexqjHUkjwO
hZ8Ax7cVuNRgyJooa90dl+veVXW250rDicoGIxXczlbfISST06kQg4cI1MMGTr/49eLM3kFZWow2
mm1bIsJjMTzgN5Tnr8YsuglnIQ0PuqfwlSPCrxwBuPhUXLVdwAehiEo7FMgPFp9eYdFzSD4zBh8a
zx7tojbaBEI6NP83AVIHH4g87gLgvpRUQWWGdtbeAZ+jP5Jk2RanvtSRp0qkdFAX3aoFB678ZU2C
vBNaUsBeGf1838uU6uF7gpvHE89OjPLAPXpxJZFlDP0Ly/nxWKI0xT0ItjXP/XnJfUsNLwRuuBUB
dXlN5h9K7jl3DTLcjh0XbCNMLELymcbGT8JEZc+25yAufJfCV8s+jFLk7LXBvwWSua3SF/G5+UfE
sxeo8p20SVqrKbS9Xbq8mkoP+lP3sXJmRLGtCgvXCKISYA7w+o7vRMyveSA0LclnuYAin26zCFuw
ClfbDEGghyPASPCCL+bhYy//fNZEMXNlNFzXFF/UGluhhbYRc9YVzZz57iMIlHvWbSIktOdEz/4t
CEvQerqzoQtzON5yCDJO9UFs+s0i24VvsvxZD9JQsh/FGzb18AwOaNEWzYMa5u/V9tTeaGalSMk7
B3cePRIGU/MCOeZgOoYPlqlHVxisTYa0fNyGL8D5+DsPv3ajAZU7gVM8DBLnPdFrB93SWCJMeshG
eIj3vTLgd4LTGdky9z3buswrVtKWxIZC7H+fsiFcGtIlhx9IikS+tVaPUFl0S/9zBDq4JcK3Al9j
o81VXbyRNvZmB2ONrcGTa7X+EsJjsLiRZH+ezpnuYLQkHZ11S1wAkJ1XGAfqh/llTovjlJ6hglHE
VGecHm7BIhAyexDZQwZagkQnFB7JT62pkP1HmQDTbBfB9Cx/cM3GBVRIqmsdHsTJSTbdGuZKxM7e
gr7EuHxc7scVPPnokEcI7m/jukzhC3bxukbQs23CS+Ky0X1nRYeRTj9nysq2GeUqVzFyR7C5Y3Wt
F6lUgVLbCvFFT5eyqNqEZ2Ho7B3huZUywOJ0402cHOSPQFsQ0+Y33AQa3ifSvTrNzw/VTANppYrS
34Ug5PNEyG2N/mKSe947Ljh39ecRDRvwA0n3oldzXyB8GFZ7JeVm8Kr3fL4tgANHspuK0FTpdwCq
Zx1jVNGmirq0MiKiSQTt914lQw+qH5CUNb32beYDbpggErrR0mX7N5rPrdm0jYnOJc16NKQbbjg6
eijbUTb0h1V7JAv9xaE0Vn53TvJBuMhBhm8/XkIhp4Lp4DPJMZCmQZcPYZ38NG69Z3ROmecfgq/H
Q6UBou+CkHXYoIs7RP4h+wH3XoTHsvPUNLKSeSPe7BFbhCKCMgiWdkHcWNhBMHHqBXa/W5gM5TKi
S6C8Z9LTUeLNY38CZIXxX+VrSiMUxjGW00GStb3ijp4U5G7dO/9m74nNdWWdfFD4s7rj+qTKYlg4
pyNQlbkKMtaIHyBXj/g+LgpJ09I3tDP/eqQ3c5VswrKbwMcBLGyFvrif0F30DyA53Bk5KQTlJ8Fm
zfiqr8xQTHvUJX0aA3NUaSNWYWhzy8MMtPjv2XujwBIHxLGlD8F2e+29eBvqeiKhh+WbcvYiaQfY
I3PfjX1Hh7z6PwojoZW2o0QNc+13AQwVQlBO8WGtoORohJwl3wksrIgUU2R29AidAuMz1jGTrLNZ
l7cGXf0EuBAAb9x+uTRocIWloRqeDjP1d7MtegwPwGbQbRz6XMJsXr3Ivb8lKptSPZlMDSdzFkTb
pihWm+euRvGob1kQmlv7R4PFU7GZWjPXg3wNsKzChQZmmvdWdmrTg+RiF8kb42fBBWa+HCKgC3Ng
rka6tKc+jnYyK8KOnQ8Ec5y3uMOhgfDKOKGS+4OGYv1pBG0CgQskqSlxgneHfL/YQVBs55rAWqmM
mChtkb0BOq8cq1MELE7vctWxoDu57AeJPdtvIuj/fILD4PZmJFhHW/OLJtsfztX2CURpJj/Z3WSu
cI1FrQb3u6sVA7ZWXoWIblAS44C+vIwkKU93bKH+rQFHtqLPAeNVwwFTi1GmcLUg+5dI2sFNcI+I
j3QZxcnkBQbY4btDnfbtbpctrj49bg9rRMFEcykO72VJqZ7FAkfnkdG0a5jht6l0iphLewlmEWk1
mwP/3fQV8Mtf/xZFxuI0WzrWOBmffnCfgheyppEsYW4Z7BTQFmmaZlHGdj/DEkP7PJGedhzaAeSB
yI9fo8Fzb7FSvZT9xIHbldpu1h3ZURMOvMe3SOJbj5QQ/9KKxUsY9SuE33aiELos/vPd9M/ywU3x
KAgBdZrDSUZxnrhjnoj3i6rHSt55ztS5k3C/UfRQ/xCzLryIVl5+z4/bcsCdvR5ejSf/7aOMkb+W
KYNjpTm+eAMRVV3rV38pn6L9IC4SxNFU2lQlxYJQHxrNOzazDiknL6QpTmbuJ6DvjU9Gnbyh4MHk
678aStlQc+vRoLNREQH2EXYO8Dsu8+8HlsfRi8SP9zCouAtuLZzKI2figQF6PMr8SqfZvgYXZrPe
r5UTHCIVSaoIposjAszTzeeeExqIwZmaViKrHiYnSFTu2cehtsvrDCxe43l+uykDhDZZJUsSvDWF
MYAliO3zdzi+eVy06Up1MqyDO5/sILVFz0IxU+UGGG9/nmNvDJj3pdJygfhADAojIjrzYQrlGXIe
uc7u4Ek1Flc9OE06v3pYmiRvjTQlyML/gn+9jDES4Nlk90FL5wqwJivEYBF+O0iMGlcYx9xTRqWG
RSV3TfbizHn7ZWKRPKuuvNOj+h4nLQIsvW+r8mq1w+NIUhyyf+t+4Ogb20awjDS+0v8MB/3WhULA
F+r2qKgUR6TBiN44B8C3ec+WDhr1DflM3mupG86CM9XxgNAtgynLtd42PFkP7n1QOuLB9fh/N3rw
kMm3pOTqJmW5Ev7FUIZ8p8F2kmVwOB/dADdM6/F2YcagGy/4R9U86ryyfnLSUbgv2LRik+Vke5V8
Q8fVUDnxXg8XsHAJn0hFGzDCQKIEBZsqxyJuzFQjfmsTrrOps4472L7gmdNOVf9a6rNA5cxUB2ea
7CiSTyRpMkNUpKukGYtPuJRQAPDSnmCpcRc32rliXsQPpd2qrL7Blzs3YP7oRyi/FnrXVuCzwvCM
SeKnJTfISEESU0rVSILxCzTGWDWK9Jk2IPxOBAyvpEBe3xL/vP1vruXGBF0R/zZ/b6F+WSrxjGjZ
lYiOy59i5WfbJPvrWbWsMgV1D8AWJDMtOVgssyyXbk1W3/e01/QXHUA5b/3gmdVQvq6v7eMGdWi2
5jYfS8EkGuTy/oIGjG3S6z+Yhg4l5SiR1WZ2c3okEMV7/SHsGmMxy8hu3xuAs6TEDcReWgpQVpx1
/VQt43RjyIA7KW7NHoFgS5fyYqSRiITD0wn9y8H9gtYHHsE0vVtAQu6ypxBAzKfsqx4IHmSGl+IX
lr60rS1kMpqHGle2V4B4eRzX3HOcP2a1iMGwMxi+2oFAlbKMw9SJ8lb5SQ6dIMApSttL8DevPgdS
FMinf/kZpexIHKBVy6ERuH72R9XgVcEDHDj0SRkGVYvorRZ1L98sFIXsy67low+YvEY1Vl4GQZKR
oZFHQHWBGRLtdCByPHZ9EeDBkkmnNWcXBZN30IwsJ1ppwZSbhjFLN/B2oLHyuMRzR/p4VQxYW33F
HtpIQW4X8+3Hbwa3VUpVIbbE4w2dfHeVOoyvzumM12lQ+a3cjNH9jTiuPPJkOgWqaOaP5J9dtAhO
naxxwjHxUeY1M6gjitCG4RayI+GOG9fYaKUmDdL2ld/Phe1eX3yTcCb/lYVbWSTtoX9aYpWlyW2T
QT/u+dNvu1Sb+IOT9cgMfasvo+FCCqrDSmfgZRm+Iv5J8BrcGaeUfKdX7+i//oO5gseqp8AGJDnx
eR/mxY8QGvLu0oy00odZJP4jG+Zl3eSlMbeLcqYMkzRyAXoQ417aDvaadN1m7FTOZcG8lPPCKUx/
RyqoGC9MgTQogbCSYuSu2zj5FBzo1PVfI0nxKfqcNTaUUzIW7l4TVEYj4NWxNIstcBeWznVgE3Jo
gnVW7hw8hWEhngGopkURi/p/Eyd45VDYhFOAa0QggQDqG90Q3xE1aSXtHL3Ms3mbQ3hUNAAAi8zt
cH4h+O0WWkt+OBg/nTIYtovDjCMfSVISal0PKSdSv/pNSv8+oUHbOD+9/ieTxY5d+zb7819Xb91t
4ZNQWfdjVFEktheFv6HDigUIvHOH2IWPbnbohY7WO7ESW/YdDkOWp+njxya7LwiN7vfs6sVKEk1d
zi9L3dWU43dL2rDyYOI0aPO864O0NPUOAIij52ds+H+eP0oypHmf6oKlbzU9thgvRwyrHzZUscc0
6ru2Qn2VFWnvCnAqdHf217Dx0djk8tzW+wymS2VTsapJ25RvDcXUuU7gU4HK4lpFHMY3UktAc6uJ
d4mTK1OyF7BiGiSr1++CjQaVs8G2e9TPiHA3GXKXHMqYLIJX+71vYCqAt5SXTeL2n1zo0LFp/6LW
QYm2OwqYp2gdLSlAYE229Wf7uW/l01C0IAH0zMv3060PtWsnUniIlKAJm+7ewbsG8CblusABzgVC
YRq2gM9AQhOINzR0xw1Ix5UDqizfe7njmbb/fzG/R2doJJnWKxFiePp2/TVQs3dP43H29e/TBv4M
xoFLXdQleD5BlnZk7ZC3YLg0XoORE2qOeA3o7EVQ57kO5ZeZJN5oNlLKLT0i3i3KygDi/crjucny
wQ1ouopAfNh6q2DY6wc/3+Upw+l5NZYJl4TAypX1PAUykHIw7AkiTWjKR/elCDY/JrCRdfgLIEaJ
HJVuWn+iK9vmf0GdD+YtKIaZazIA3wEB805crWAdqiKDRQPJUJ6rIAycP8tCzLaJOgpBNzn//2Ir
EGhyjd4F9odJspOaTuhBzPNjGy4k8o4o7YNYZZnrQ99XkTXvVtYct3HMPdRhzZUPESIDfxjDL1iI
b1kKLk+hDtD+0g8rtqgqzE7PnIj25HDh6RppXm8OI9DUY3YwgFv9lNoTVnJ352FuGIxgSM8PwVpc
vo+gy8UiEKmcDovecxJG4HB8M4nn9f3X2UDZUcAz1txOxCWddMZCsigkaL5adLaMpGDHk10JPfzS
wvTrvqT+GRo8ghmKDzgHtLcRLxDHHR9Ce1w4meUhHKfiJorZhR6wWzeXUVwXNE1JxvD6WZyPOqtV
8OQFOaEJcwQJLNHvE7BS3evfToFzH3xSwMlI60sR51zWyl2OcWzJfynlq2ACzphC9/03KteZrtmc
I2NVeFzxcjdLHQccaySjdApTevZwPthH8BR2aFhmRmHkblF0iXGMlTfKZJ3Luk14ASVaqIxlgIem
/YpaVLo+k16YrgirKMdeXFkHZPUujb33HX+GsoSsStCzxg69tXwcLCPNCm04hDjArWzFtaEUixEA
ibG0W9rzbtL9TFOYOmiIeMjcCzXXZH0spXFHBvc6j3OBPRDGkf1oM9PcKtv6pvPDhWwNGHuOipmI
ldgY9Er0Kyc6YU3uH3fNMJuN+QEeTUE/wRq8G2oQLEsJ9L6mKjgbOUBRYBAh0Xbmyl7LHkKPRlRw
ALLyd7NSRET9tJrV8xAbwoqqHG6E0CIg+OQBk9GLwx2IxfM+yUwzL5OC49AyEjqx+IcntWxZgZqr
Zn/EBPr/5FnkM8XvSB6jQPWfhpEAkoE33bGjijdzUHIv9u7KpeVChI+gO0y0Vg0eP1FGZAe4jEJE
GBnTLjxqYEw6ZeaP2Jw6ZSogu+iLPoMrq6f2BuX/IaE02QlnAGJFuqBLtJjJVXIXasn0VMF4Mnqf
BuKl07ZNwXpqUIBKeWOtwTeVDr7woa/EX2NAzpljKLRsSy2W/KugUM7VqvXZg3rceSXVfrPfIVYj
hfMhl3c1yqeRzxxf4aBC49pLSGzwikFBLED4sQJRvipO/iCsWeXayVO761U3tEz4qSpcYpvUDKRA
hVE3a/wrHN5AP/uBBTmgXaiZ/mFi3qnaZTp50iUnd4k38dvmqZYAdtlOnZ0dl+Lx90+GdFpEsUuj
A2f0VqvVTgMyQpA8fsXxeMYCJhNUrifFrNo1Y3fv1rrm36su4jQBcOlI5Ot4pnJxOcMl9BrDktnf
IR0aTcxPQiOZVGzdoezzukPP4VysYZ1us1SHb8lZvLtA1e39EhlwWCY4fyMcJ/OHWrraF7IAVUS5
wcDI/Za7CGs1YUAD8CD/DTDUG2XOXGOGEeyRQ9zvrQjM0OHrDsQ8gMpeaocbVRCLDujCkA2hRztc
yacIPwRjnyNCJBPJz7OqgKPNxV0pcYstglwg/3DPzC8ESvDCFsw8Ix8Wa+qjv40ZwSUzqY5m8P3u
VoQuzdC9mxjXWKH4B3DSQ9MmOwpZ3fbgSTPoVwt48AKBXZR8rd0/vKoCaag+/ROXBfXtzrvz8qDT
BcDsZB1qrHZaWis9lfh4Vm+YA5bguNjsckfe4gVnmmmF50cQXWcb0TC5Yb5UT3WsJEk/qnc7mUMD
ra++wgeWV9/93DhUfKgpuqf6JFnhdfb4d92Gwzq8F7oqmS2/v3sVB3FFB4XpRu8Zfw2eeadLaKn9
oJy8Aw7ItwOG+2XeSzWIko8cViNlgXnEF9kgW7HL9QYMcBnmOqMEB4RjhnoAlxtrs5EUImUXnXgF
Udi9cuXwxvBeqvY0B4UxhSGqUwG1OsgxGDM0XIueRFSto/NYcXymTn2UIamCbvCoBCZYG+hGWwZp
ha4zE5jfEKm8C+sdKV9cLB1Oo24RPd2jWpXz23qYEFyi1DyHOjRz3DU8/dzgwRGiYP81tqKM3Bzp
duE9Atl9HEFy5oo6wlJ5b5BO/vldl4sbx1qP/vw0dQxfevphWbP8zZ/jyJZS+XtDtmg1oyvtwODR
y3jp/0EKPO/hiprsge2eaQ/2pBz2DPn43/2PUDwOv1gfwopyBhxhMz98QvleuTh12FXa400ZX/b5
RUIAhw5VeU37I3VS8GPEwnCeFP0Q+SsH/P2yMHg1u2P3U/o6z48+CNyg1Dpsbe2VfJFkuc173y7A
DLgiJxnL6jUgqFzZWPhIoGZ5M+hJyx//yNnDo8zxMIU0jj7uS6o4t3SIYBDslmcutTkASLSrGYSz
U5gCakFlf2A98wMmETPJu1OeTnhlHH7ffit+q5napI7K05UpyjyagOHkdQ3Bq3wTe1ZNuN1OxDI2
Js192dUrZg56Y/zMzANEy4pUVUzUtIwcFwEs0niphX2cJjyc0NHEalzwg1Nem50c0bJMnKQ4bQND
sqCEtMEz/Iy3bv+xqwBaEpWh4Zz6rPECGXhze7lQZ7XDg2ScXYgjzXim9ySmqqZj6l8HiqUJq2cI
SLWEi4K5nduuRwItqJIjM7kK5vtSpsg6DhdHZnI7iMHLhIszr6IUpyjaJm/AXzC02nhU0/alpkpJ
7cSU9bCogqzkUnikr6dWOh2sBUABA5nXOdmaRh6MGjU1T3GY2lBBm1IM8XVA1pJLfyF9ZrilwfkK
vvw/dWWhimtgQyA1/eA5s/ke9xL9IoAGurN4kVfNr4N5JXCejzh2lrjMPuwxsqcq59TngfGZR/7b
1kCBxYWCEnPeS+yLTUZ6F1O6+kxr2nndWqSxysknQ2acPu5xffvEDFAxfFRS5EVGTzWrpday4bP9
meOAr1igPawCWc/DOr5sWSzL86CFGeh3pbq5SC5Yl6DpECR+HOGcSoz3m7N2aUainZE5okfVf0GC
owkXfXNuna/dEc9Y940gzeCFn5KESdzry/T7ZV+52jiCtiL0Pfs6RjXp4Yabdyyh47MDg0/AZyt9
GQsYgANaPCt3QfdAc63Jh4LpfTLNmx9E7rcyCKMQcY/7QtOQYzk0EXlgqdIWB0WhfNEUHa3JDtUG
0bzsQjAPiu714HwOaneH5PM4Kq7NOVcq4/Thg+EdRQRLFdbsqygMzls2Tdfuj9IwEUhOebX+wjzV
HvHMehhBahtd3zruoyBcczEZYrxwH+6TqMAc6infP6c1UQ8Esmnr+hSOc7lWVOkLiXb661Hc3dca
WeiZnzFnpYtx1D90PcQUPQj6h1c08MlZAdq8TgQwdxNXNlKmFVoPN5VjAtFfcBxcv6dNvSZCFYXW
jfvST9T+cWqGMGzNHeRC5K/lYHYD59sfGdUR/GREOviYpYqsrE0RLrY4NHKAhtvlA79FSCsOXOw3
lC/P8hI4ZQwrzIPkz6iZKT85NaJ6C0tVIkDZID8OLLHlPSqck39Owsdey0e/pJnmZzurqzd9hKk6
r4AT1xz0NGZ5rlp+/Sznff6P0pt5YFkM4I5+HR6t+Mh8pPVK0O1lSOFrdAX1XWuy1XmfXxI6Nv3R
nToA5Na+2GP7rr0cbnb/XV1OBThR3lmcVD3TDZCICu2Q0byYa54DAQ8q36tqWCkzK4bjl6bgaEaV
oS7CZz5v0xFr5yzDxHtxlaa5/8OAT4v5YbfYQpRX9KgDEHNKRV9BZ9T9JbVYCcoTwLbVkC7GIrBg
H737LhizplLnqwOma3CzOs3Crwd2PmP8oRvaX4j+JOivryOx5m5YNM878rI3dB9AMOn5gACKicUs
mxUHX4e9g1WKG14nhEP+jkQg+ZBmDthQ+3gobDet0r3PFHTDKhuluAznZl3/HJa4lUbF38ByJf7l
/5Ceo3AJtwOJqhN9B40ySEC2Sxqyuh9axU1CapxfCkfn7hWFOIBkXZzw5H66XVDxJeX1Z0Hh4LJs
AyXt0P4hFDnPw36n47Rn5nOOTImZuBJNMnudNTejqpwqALWbKFJFdx6+ZibhOdFlL/oh93CEkiE1
m8xfV7Ftrte2TM61Xfu3561nhCIQgx8qlFaAPH3f/5W7s2CCuZC8kWCXxG1Ouud28RnqcXzWRjGv
4Ex+mA1VA4j44M/qCYMqgQVGX/XKTuywTtqQqgvMJF/GFfpAuxtsB9ajQruiGmy+ffm2lCjYvEX3
BaU7UafXOVbYIYaDnV52K2n5MfS8tR9vglETXwePD1Mr/jY4b8beAvnQWnTqGaY3W0NaA65lE9+W
gtf7mrkHs0AwCQAaXcgvUIfqwVBIq+JUEzZNi5vAbzScbCMlaYl1Mf5cPuvfdp6hmfDXozr67Ozi
Sm+BNZdj+7y3mBeFTM6S4dHsh0HtdMoHGGYCb7nU4t1kuvuUb+qXtNM+irV7uJflqhiHoZQZ3Lsz
QHqOYQlFpsFzp/88KKB12qnPkLGBFkZH6u9VkuKf+yewdx/buzBEr5JL8mTrlENNAphivaxqPguG
Kq9U4EphsYdw8e4gutYP4C8N9PyVjfcm1NesQ1zLZ8chDJGB8L25vEIl9Jb4msZa4mOWizfuDEzL
XXR3mqDBHD2+95RkhMFIF26iOpn21rc+L0JIMMv6N5QTmXAJrATXNhkQ1vo17DdUsYTX8yCM5PWx
Xe7uCIFr7vgyTqxd9kVeIWfdCHvAbNNIB+C79qTGbujoJarVOHBrZQM99I1O52jl4CDdhmd3rbkL
BIonuvx7KIMuXMLTXfG0UJxPR9Az8H1ivb68sINNLxdGMT0HIsNlgiQyjXgzP5rKIBo2cwBPNbQ0
c1hZXXQBuvLtcdwdBdMFN8G4KNljsW7DXw/OoBwp/TA0SWp/E7fteKQP4cBiKfZ97cIlHHcVhSvr
bDsqDAhKAaqpiFvCoqhNg13Ds2mrDFdTW7Rx19gN5d4zERPJxNbTBTRI1SDmMgFXTNQCVrqgiJ4h
rAZgFlgvBWUSI8z6Mhhp9qv7wtatIeCtJy7qjjgbuFDOuSGn035NbVYYgU7T58mXuB6fvEN6M80P
kZjv17YaHGdx+42fzv7Bd976sYpE7uzy6hIERqGz+4D1q9leFzk+OPygkQXQleIbrN40HWTTFPkL
KysG/Cukv/ippmnpv9FKW8GJ80ZcMgJ9hvD4o/MNCdBUhEztwCAIk9/VYAutpjnAbcluKfYIMnU0
W8NUFQN68tkVPAoVoWIe4rfB4LzOMKwwfl6oiBI+zpAiD4VjGoHSKiV/u2ofrJ8Z9Lpq0eB20mvv
ZH/tjfV3M9r0O9vmObkl8zCJuBZDAlK49u3YWShweCRrabjqGLY24DfyELUD7nGxsWoRokGUe2lX
9wP5wEQbspoAuAb0BprnGoBxphq7JpH9tmLs2uVKFXdiVaNXd8O6l1Dbnkfbgffi/839C8OuI/Hx
Zb/00llZ7vw3Ox3VHB73LtzUd2azqVNoQLSDfxH9uhYica0uge4nsyAEIcYZujqBSQ8cIWsWGlp2
Mk6JjFocKmvP3LxPUlSUwQL+eGg0hFUdftHCXDLDwjIv6FfTnA92DI6yFsgzW21FIGqplDX43Q8k
FJeFzFdHVbplXLCawtPuEr0bcxO9wx3tT6R7b/ZhdWGdmanYFkIRZjg7oXOe76DZrM1lXg+CY6CW
MVtb57DydnTA4ubT6iML4T8i/xcdJFjrlX65hPZ7mmBXKrlGMzWMew4vBJ0VgfwFnr8oq0mKnF7D
zDymcyNMHld+qQ+vRuiDd5WVCZdIxpIxetqOguJpmHX6Xu3Jt9IlLtzrrFHtDvD3k/Z52tlChAtU
1LnkG6zLY/juwb19FrFl2TWTxTMQ0wveZxon+a1hgdK0yvoHU6KPdynQtDcIYP+qnr6uVqXRInmY
87ivGKq1YS/t4xFv/KrDjaIwYyKu2m5m1EKvuh5/FWNt9OFsLZugh+BYrZv/5r5uypHFaursSpZU
/UmsQUSmsRIT4wpXVQgCdxkMfoCv3IP5VL42UUX/JUKCv8Q+r/vQpe/IbebhMGOfg4whn+QgkeRj
ddk88IA8Exw9oqCSj94WaH61GFbKNqUmXx4m33YxxCvv/6JUPsRSF4Vypzdfyr8zg/HmppGHPK+8
eqeB+tKndIYU9VoT16CjzSrwN69Pvg2b47TFWLO3aEhHDo/ehhj7ZxzPXBA/yQ36tqowHhXlx1gc
akGXx8YzO3JyOWI+1W4DI9w/F7WhRjiTr0XuEWdm4vZIFSnoX6zWKV6atYeTjJJAeVOpbLj2+NeS
OI1k2b4AQgTXXgladyLFFAF3um8iBx7tDcU0hvjktv34E7BbIUbRXAV0q/OyEG5rPd6by2EpJvgn
Bp6F7lx2ampSfzPDk+qxBrYXJXpjlGz1mNOqTsmfdFRKifWZm1WDLvhuYZSfhNx5JWGvYcy3dPs3
FrAILPnB+7ywO9q/mBdQN3buxGF8GVguN0EvThnuu/vvaYgInGV5uk0bU9+E3ohTGJQnA3aOBhJ0
866wu0IF8+VueWumE6cFoWyF1of3fQhr6bsrKiU91S2NtsQvjF/BhYSH7eIBxkDC/BZW3r/o8/Yb
IG3Xx2uNUub8ffXPdsAxvjernUH1FTQ327/V5X+E8rR7ZKVayjfHyAKyKUmnYayqOS9wZhd69giP
3LzceoegaIjyzKJHadISbO1W8Pg6OUdIGnl3m/NSMRivq9U0hcbadEqBczgTNUDhPbMEqCSSyMBQ
pc/yx4JawIKxxY5zsgpuv+qlhGk+EOMWODGrQAdpKQC3nF6sUVjBGUE1aeZ4j8bhKOUB+HoDVMeq
pSKleoMeUTJJ9SxuP6RGFULzQVywQu95o85AGoidH+N96ydwFQB4WaBp1w2BH9SJUmX2RTvD1Q6D
r9xydm4tlOFZlgEGghZGrcf537sk3+TstDQdXtP+ERyIirdyLowjyWMtinsPZK0y8wgcwi82HaUK
CTh+xyUsqXvSeLgoHTbhrm6bcPtyFvc3kATE/Kzvtrcws78vKBmuWNz9LXpVjqozUVOrngsmaGRB
d3gWadnmrGxLKDShueTi3eCBxc3ntEawRE7lce8d4KL+26om225BBC3bpqYfyMsiy/e9PQEVTGHv
3xMiNxzkGwbncnSygdFFsxlG8lAGpXDUs3pTawA/e2YPbp9Q6S2HN/bcTTGF+GW7u1JPegqjqEr8
YKUjhRi59AI1qGGqp4NgPMUFz4HmwhT0AdDNNMAIjRCximw0HOMKJD5Pd+ePnO8IKoHNTAJb7wP/
BtwFUetFsltrSol6PB3NA+2rnbIiybYiSJx+gfX9Mm8SYxLS8tWEdXU0xyyAlKHwA+n6mrS4mlLm
56dFsyk9U9Gzy6Gua4RLJhsSdpVydY/juiK2leQtaYCAyxQGYmrRdr59LdJNSzRuKSGP4F0t7stX
cjo5BB4EpD4Hj4ZrS3ZPDKdHvpPueAPnf94h37v83RDyRNpFp0OfpY0N0z8NRFUwsU3wvQQGk41A
Q0QJSFEXkPJbiMBgGL8EbBg4kwmGqstJXRdhwCyI/eutsb6EWGsgETJTGpbg9gtuCWH+1NqPYH73
t5i/4Cmg+b94IKZFLswcN2ogWki8Wd7iIXR6KrBAng6maW11v97iFTtd4qQZHyywTtV8VZFUkcD4
kIB2s9nfvr5uN83RRv5RX0Uue0X10CHesayHc+O/Hv5fKaS3buYRJFunFAgYEuNJ+qg4/GV1wNsU
hfVbfB7XkQtBgfqJ2RZG0MX2YwE8QJo5DWvTFws3xZNKLRQYN3SGg+CNCF3Uzw8+ZVvkM8+uJkjH
cVf221OAgC7b0wCgKD0Yu1cMmTbDnV7ha4f0qhhEVi9UBHzxBYunXi4KdPAkiCirc1UDsohAKUyB
CMc8WkibIXBSjlbsVjYmxYh8CV4kTa4LzpZQCxDYorsEXP8qY62On6VthAbDc4XYV5346KNpklLE
hh2SFwOoJc3Fe4khC0L4kZjGxh24njEX0MzwAcZsLmieliRuIjA2q8VhpqpyfucYOKGfnaf5LdVo
7KZbQ5XteI0vhOmD+kRNomxE7QaEiwKkPsc9ER3qZNm+KvRaC+EmQJveja2YuHaSaeyxinNOQuXM
cd3pgQtPgYzNZlZgoAIaDc2GOXqyc9Mw8kvgLsqlIay0fQhQ3u7kQ5jGH3LDSr3/H3QSSN6iiyci
GLmr05O7qAsYf3t8qsWAr/ZYK8lT7WbW+4OZ9xiMAYbxq4O4EYXwP1LJqbnWVw1dd3+tkxTdxkNG
yFnE5w4egOxoD1U3dk0t8iHdiGaHPz4ktEVtkDHCup+i56X9VeaGIQWBlzUnc9Gn48ibXJuEh/G5
xMAFnRO7hnOSP+sujnspTcOJyNPfL14Ee+yBbw7Ybe7xeONZicX0X9NcQh0C1DC3VL8VL1nLqR6S
DwyzHIqKa3GcvTvPHVbohNd/klBVRyoL+1KnmQtTV5Mjdr4jYGRjvrInw7OMSPufkU83/dXD8U+k
LeGk2RXc3Jb8GtQLL+5XzYPv/q/H1k/TnwJgaNayEBw5oE+7KmOseAHsAuHkMR99oNosMEkRGtj4
6MJ5pv0sX/VJcGlQDch++UgcQnwgFwRhdbaVv68bSa+pSn7vdwEMMykNlNa3VlElluzVtYKonxPE
UvfFpzq3YJAxdlv2jzR/LEVBcPV/RxaaSf5MET2IHHTglNlqd4qW2ip5j8PA2to4IB3cndguEBlx
V3Rw0Fqwfw1R+FrKdQ3JbKWoON7rSwoHxuDPDFu2XpIgU4FgKQ0xDvaFC3ZwbrI4xrx7ZMjMlKSB
rrK1tMVzQx72sku9gj6Rc4nxQoXd1Mdv99s0hQf43rnx0AV2tlgKdpYs3Q5s94IMZFj9hqKU+Ml5
7rnxM0gZGqDkOhjfsfNNJ+rydsbOKR+Ay/LFh09utKqL+WeEB1odRAKWX+Sf6RjzOb3F0H1tD2iA
vxLI+dAxEAG39rM1W8bSZwLKMH2U8OlHO1k2FeqKILrx9R4ITvVSlLYB/k6QB5gyZ92BHf/my5tb
ijwf3Bl8xnNcrlqvDjV846oo11H9rammsG40fZDzfEemONTjGVsyWuObP6OpQDNd2I4OfupDjL0n
8qWNxxWFXp6sOv6p+OlQqruzaXxdugUb9022olMkAh5hyVb8BdK5RjvyXhqbwySLUVDXmeTLd2nL
KjsCHn5/ysn0F2rD/naowe9KdLOk/ecyycddJx+SzFAvkkADpe2FS1CH2f26zr0n8pXSWUnV4fEH
U8vtiKrVF6lUL0jszuKskCgwekoIDs+JxmSyjxqhPh+0nwggtvtKEpAgsNYHrLmfUst8TxwWSBkb
E2TfcsvGH7uldqeLLELqlRRxk1Tjip2yi9FS6l5W8bMAjuqSQ51wjrRhbGqQYZVoUrV8/Un5saYZ
4Eq1SJgGn5zpHlrMmVGNlm6Ofo7tAVSKW7/3O05CJFqADgS0YUgzs7DmxbIDjD8/1UmHC5r0llB1
huwbTN/L6rjoXeHYXZEaMDyNHrhS0Qsy3i1qubXiVwZ6S8RC4gTgngasGmD4KXfWoSuBOaAAXpwU
KkqOetjSA6TR7Lx8QFPQRzniIl1I0LrzCb6Gi/S94FrlHzCYhnwqvvspDWMadNASU2hcoV9cwmlI
uk5KoS7dbNaU9Y5T/UeYZk3fpDF7APxYqwXnfrsg6zyv54ID6eqT5RLLfi3WsM2N3a0y7UMRrHr4
35KZ4yDiYIQL6c6ACktIPGFtyKLxL1Og64EX9KDYiENvpB+Q1F+gvCOcBQZ3IvPtD7NuQ6tfHbR1
rpaEOE4kTmW0mGCuqKNvudhC8BKH781MnlFWtjh8FPNAvT7Ji+dseQyk4iTikOW+mhFbGtkZMesr
3FS0dt5UQvSoDUT0JA6EPvQ9XvdVeJJOJxhSmPtV1Zrt0sI5k4nOAGxoCJ8JQJ/dfBwzb3+Bj/Iz
mPtHHh9NGqyjl7MSSgvs6Hcg2BxFXA44Ys1ghASDIzmuUcQX/kr3qa6lmt6KDoM6ci8QURmNsFSy
CVw3YVVaEXI/7S2tqethvl+8gEcl0/Rm65GrlANV6hlhXtcQfJxzu+dHWgLt2ycsnxIA3ibL+xTh
ZOzEhehPgk3veDVv6US0jS12+whEO3LsevChpzqnpxIbwnHTPIjqSkr6jUmK8IA4DEqOhV+akI4b
TdePVSestv0hCPpLmyYR+YnuX1yDCJO1VA3f2j3DrxSUjimwUeRpviTA7vWQGry/hgxGD01565Mf
eAEYCrHJ3+zZIXWRCuL/Aa6SKHmXIANe44KsXhV41EXAcvA15nYaE07mDs30HfEDr0AWt/a897IT
8YG5rUZgaO557D5hkMgyKxbTx1KKlkRXyIuuPvBWCNvj64y40OneDXc5DZZWXM3vAQqPDNBwyTtX
TTrjPIudckcg7G10xLa6GP2Xd+9sC57Xv2y5ZDmFP8AensIJFmV8AJc6ec/h7cugUCdU5Mt6V5zF
8VVwdIzUGVBJnw3bVV4TS3jHswywkP6EmEDiJ85o4NCLQVC0FR4g1WK2VrlxXK3QiCUpjCTEv/sy
O9eFyTmMDTMwJy1qs67oSw6ojnnYi4yJr2ePASeZOpyQ5aJmN/KqS/s1jTqXSrrK4B7U+gS9VdKF
oyCmZn7DHC5JH/1VqtuIY0NgIQbc1YQ0npTNa3UkK3gsMV3paP8jeqY9FARTszJ0fDVoIMUxcCMK
QTfuSaAtrtFkFmsMw37CkMBG9/XGCGl5ogQOEWRARBJb5J0dBJ4KFhP3Wp+RWsahZfDJZzjW4bkH
mPbP/WLWt391+XIcYZzY2wuND0C1VcfM9GPyzELKicuFm1O2Ed7pBiap96iVVbbRuVtZmzab0ad9
z2+Ye4NNP5BZ6ye0np2HLhGLjqCX2SBRtGCtV3vYmYZwWR3PpiVybQV9LNYBaStwshjrwF1YBYQX
KQC+VvYpHDOlJVv9uXd1ro1Z5t0lxmRdQ+16GbJUMXhgIjEwmMmnlfNazEUf3E1Q5UMVo+fCUhoX
37J9WRafPelOb06J9YOtbVAg6+ZFA2aZk2j0+h4ghbDkkq7GuCmFdw6sRtcAvXySTVWV2KECipQw
OPe+qHmoFB+9CI7IBnP6F7fIG1gA/7jwW3Qi2lyPU5JtMmZblPIRwviyQJKGcxcjmL4pYo4bb5k9
Hgkm99qB3miCNhGM+bRN7Xone3EsEumao+wKiqWOeWN4sAxDSgR4f1zF2zzTKmrLXohAiq3i7wYB
S3iy0uUjiYk2t3NcmZrPQw/tpHmvf2oNHlaXrSH7TIoFXZVw9HE2XPBakAhDezV7naFyg78LNzbi
SV6Zr5Cz4OvfpNHqtUqFXvcuVwmfEELtOxJ+Dez2MyjDn0LHwn/n+tqIRVN2dpnnxZoMxfbdi3/w
Uyl/UtqYC7Z8P71Y+DNvHthyyPOUfftD+4ffBOYancAC0OQ9bqhOFkmsoR4veyqCQd1IzPU96zAD
WkGjzQqgEqVivTfVXAEFOp4s++vF29461jh6DGFQcr0aUjQGyR5vxC+XRXcTXaAolRp124NLZKIN
JUfM9zstqRDpo6WxiC6mi+eA5Y0xiwXzkQDxUI7Z06zbZISMvn1LqeeL9gqezHpyg22ZJ1Ga6uWt
gBxCkOYzBxBivdaP+BrJOhaO2z2SutCW/dfocXmHb5VYkFbtji+S/j/J/H9JxHd0BSEycTdRvhi/
lcpFyyz6WMjKsqd26odM/9JddT7ekTVkp7KTy2+mN6UKAiLsQpDQcnAnivMN3TtWzbldztoRBb7h
vi3vD5gPUjeJ8c64kB2GdTIKWRRKeErXehNE5zvCurjKqEP8dPRse/nwVTnbrsfF2xNQHWl1gPZt
ILy8FBwEuAPf3kfEhuQXWe0Leo3jgA2QSbhUu6njP3j0vUzcLDlGexLL1lkiD2Cy63WffIk3xTeY
ylJxqGHpreD//Hz7IJHgx7FR+s7vY8DuDxIefSlGlkLl2Vonjyn40iNvem0rD8+hRTlnuVjgfTci
1X9d25AX1WEikWrDCrsQTKNdPZbWt6XGAKqBYvbZZxzth3EabNKbMq0gzMX2IYlAlInpnemO+ZW8
J7bFdorb4LZh3D8F+m2H65LrF2C/+c8XdR72se1w36+1/o0/VacjywEGwgIB0VtXrc5j3MlAjoP8
D7qirGczoDWU2JtM5AeFjaeTgo/jo6yMfwbdiKdR7f2LjoBMBw5AFntoQdrtMcq8DQ9Hq55ooXkJ
qd61aV0w9jXOgx1JK3IBPVZYjR9JS3zBimIjqL4z6dUmAYecKVCVE4YHUnhabc8cNyTiI8NTnHCT
UeYKUisjbS49FyiyCEge9+qWulEBDnxsofcGSqXgWOct2uywF0oPOHQAWuEruxJFr4yWfnV2mfe0
Qsr9i1eytX45k5OG/gKFAAKy4WS9frQyYiYWtURCm8tUXASwWJKEGoQVWLk6exnRBsFRcbq9vYFo
/M5j73R/pn4ZSw6Kz5/26PURL71w6kD0GjCioXXGogdT+6q5/iM79M4DfYGejlKa3rzcM4nhstpm
Cj0w601tjCoFyR00ILBI9OBoM0p5Fi7SFs3JLuCpj0AsaRzltAiOUcQm5xaosYtCy1JtfttaimVl
OZ6kNTdC9f/QPNRebF2XyvCPURtMr6ibtHAN7qiuqwD1LrnXR6X7C6u4neh2bYu5TARyO9pMaDmZ
WtvPX0RzFn9fuusVW3TddCRm/yG1mEsjSo/T3v/XShoBUeRaQhPoyEvMa6CAsQ2RAtxbzJDMhXba
4Mfg8zLiz4xUVxAUaY/NJJMA6KR6cq7xo/hxa/o309LeQML+60WDmrLeaqKw67856roqciPeTqrn
7RU6mVx7H9MCyTIhL5dsJhPiraJiPiHqb8P2RZ63bxkP6wzPF4opmgcyGWCu5IYj2uVMM9UXUoO3
i7r/WAcOBL7GmMfpZsdlOsg+XQ3CXccQk9KlAVp6yq4Qsd0DBSdpZh0aezc/uoIjFtDZrFe8dZVl
KeQAFkP1aRsr1xCm+UUxx5yylCqgVVzEEl5BL5eBIcw2h97+S3LLUMk39/oFmJoZvWk3VYIgacw4
+iJwlTLjTiLipe5tapIr6z2t6YE63BddRJ3ZnE/CVQdYp+wJy6hqaZO2nUh/NmWDSSEl+p5i496F
VdMA+08uOoS/EZdKAFvKnvbtyD+wP9WV1IWUT+5KjhSc1pW1pjN7vxI4qJWTXDfgzrUJdCab1fju
tFZaPie3pAOWWyW70KTWUt0z9qpkspVsQNq1R7FJU8XMTN5+1KkK0Vm42jkLV+5L9rwsSV6HrUD4
Zy5iGLA+DrVjxI+X4nVzNfeTxlH25su3V+0XNcDTvW+wMFMZvvX17imXbkuLw6YK9LSvzpMQURaN
26HukfAplacGRhUBa78cuPDTxW3JEluxy6zUBb3XUHnEZ7BnV89HtlI514/FD6+SqfN+eRC4BQUR
Ur7crcx4EI2Oyq5UUth6gJjhW1xyVJ/BTHCJYrI3rJPZj/bhMEEyrv+EJqGc2KT4eXP8sM466MVT
STk3PGSFUVBmud0ZW1drWnYgIrMw1GReqjE2h7FM8YRfRURGTRV7huo0zvRLOu2tB0JmcFVQMVcv
vWYNGGrpL8FqzC4JVa+iE+9g8HsGAKXI9kOzDClssp0nXFoez7vrjUSEt1OfUFMSBMRCNvxD9s/g
qze7h+2oE82shcgW2YP2RgdPpTa1ZQ9rSB+nfBA7g/I4279gwmiTHml5zhtpy6dQJUKJ0xuwAeoH
GvqIN0S7cbT6krUfOlUH9JJ2a1JPP5fHXMjzEuKytpSsE6WBq8XSuL01q1EvzEnC//wW9NIa0sGX
oeqRxNMW8kulldtiR2Q6CkLef3FNIdteaVM/JX1inbOjqWXc2zDB3g0R0Ahqg+73oaEfnM3ytMO3
ir+ffSD4o6o7ZQh+JK/V4kCjWkD6i1Ywr47Lh4YVlL39llCTwEIuD15vromWGUGVDnODPSpHrszZ
Ph7DbOgubK9vL8zyWQ4VPuJ4tEZyIv3NnkFp/Y5fGSHArxP4nK7R6nPM0OjGRTrM/CLdUbd18pO3
br4+2MzWTydYsBvfo7rMLgNvTriRLdwpWJOVQlGs//7lRT/KbnbKBNBknI9EEFAgBKH1X8XuDpDC
HYzDdWFzcvngiwr3n/acwIgmDC1pjb40u6WUqrw07zvgtzhSxiWxW7e9AxVJyYnCsULT13DQRgD/
Ct1qDZ4AOze/IgVRHe8+hMjHciynbTFCc1U9LwDVfXABl48yo1QEHq3L57ne/4VvjpNnm5P/Ju3x
g3NwcvnCIXtwN4mFIANBA72efS9HsPMLJYjcQG3rQj34ezwLIdqlJsHUoCi2nI6JG4i7OTrU9MAI
4qVLEGILehSZ7aJ1wxoT3DIi9y+lIwHtc27V5FWadcJsuD9PWwezC6sM6Me7MGR3dE+cHjuPH3la
vd3gP825qBWON7P956JwEQ93g8jItrS18n4Kdg48T1zb153dWZWJpGPVxsJ914765XnSnLCtDbxS
vT5DjPKsyMbWiVWhy0mKWqUxJ0PRbe+L64OpA5JE14RbHljRXsW4mlYmQ23GdUpT2R3NqRxE/OzE
RyJ+WkzEzra39ZWROKv3SSS6dACbU/G6kLMkcgymct/OqwTPTj2BHKzuh75rkSx9NklI3KpE8q7o
4OXSU4PjryVPG4Q1A+DCEq8RHQkCOuDPK97/zFyr4NFC5obK890HeXxHhIPTv+Itwsa3aEhdallv
69VX6w3TYGxD9yGcJ7+UFZQP68RXJ+lH5nEHOag/wF2N6Kbj9qiNCSGTzA0F2EX61rkl72AyWAHZ
jW3eBqhj4sGkuOYa6W5vKqAcYxjibn4jivHXuwrOupSfs3lSVQUM6FWhbioKoaGRfBCiK1tfyh0M
p+ElQBXP8Q+Gdh2dI5XGlCbnCY2ZbpA4DYMxgdb2fYhDi+N3UmarZRNkdGa6tr2IIvRjJ/c22Lbu
CKHUX0bZetzx/LRcAdeYk9P1DH3JD7rHbPYnXybie5JZZMp3IOf9jwXTAy2iW763X7w6rLJsz0L6
CUBtAnxWjCwhBIW6gcHKChgA6z66lc1DYIQHfIpqhE3pmNfhwnqVnjWLKvOKLczDbgXyvqhDQla4
iz1bJ/XkCOSm+7qWRoYwl+c/lTi52eP91YGZrKBLReZUXSvOpIjw7d8QyBehvVMBVu2m06uFIIbY
VBErUg3c6e07pdAF8fxh0g6VJp8cfD2UcZvmFDM81EicG1etmgjwNtN8UBGFiOnN64X4oVpcRbYj
fmaV6fwTWqSoLPmnXir8nY9ldwbjccZg/FwbrGaRqMLT2uPUqqbsVxrJypyi5GF79sAqo08a5w/t
2GYMTPEsLbkLEozbJG0o66F2FDCGSScC2NZSB+kBojatmsw+tRbVu9qy8s6A9XfDGYlHmnWNLrau
0+txgPr8e+VJKz5wyGw+kodvNHzBAZFTQ2mo0lCpbN1rk+f5x5PghDz98CMdYFA8k+O1OraJkO1u
P67G52/i27C4cB5escj5AsQHlyYgb/LrCgKxkNUOT2I237lSAB4KfCbWaOzLqfouGMJyCU4Ni/g9
f6lrgWKktoqDf7EhuEPTwtM0S96fgTQW4mdL0u7hcrkTf9UyJ+ciAH9EH+Q+3StU/nWOuw7qgrAX
+5i+thRzQWtN3eGurBdmqCUTfHK0FVWjbKz2MvHslX3/qOBCuDEKSJPJX7RuVbzfJqeQoxMH7FmP
c873mt78mcNcIO8VOwQU/UjBJcPXhcCQ0AJ5xi/JmvARmcc/TqzWkhwnJax7SX2HEcCqRkal+VdW
3MOsoRvoWTF1yab/5PgZUgM6/UkvLcLzgpNCGlMHnxlrSCA4ln2nJnT569WJmrrjZXm4lqKNnDu6
zpCA6GnpWEYUs+W7tFtqS60LGznMnntf9HSii7nJ3Vgn8fNupIt0fOtKeO7uETUn30Ky9Mb/pAT0
aNYgS6+waM5HZ6LdHvPx2NAIw2RAK6Evbx7xXpml5yS4X6UC3OQWFcuXN9fkN7C1+mNbdwmx7Azm
vsJYNEIZgqoVtC5lJLu2pDmipe2XMkIq+Z+HQUFXinc9s8vJGVCbHFM2KmlMco7PvVRP6/LeT/xc
SBhJCx6pCFZQ8LELgi2o+XNbICVt6BZYLLMykQmUaO/HKU9j4lEheCginAxAROmGdZe90IHTPwAI
JdV1mH+mnFE5RiN4IZJ9GvZYzmQYHLCX1EF5O4tzAhqPEonpGKf/9kNfZ9Gv6kDr3BW79z2vpszr
H5V3lRgiMjB1r94LIQZfSrwZBBPgUCYE0yu1sbdF/JOtqa9Xo1YgKYEeyxr3EWYloZ4j/22deNsX
6g9U5HMLBCiA9gbJxqsVGaYUGqkKCB3YdotDYY14RPhl5mQQKrIgFGtqdV0v8CKm13s5Ui9KjYCf
+XwleBN23wkWzs4F9UZeiyobhCEqtYLexqGjG8YDKYlnlYAm4v/NZw06ElULuwfRVoUz0H2yDED0
FXWY+FlIQUeM92xFvKSaaptQ4kAAeBIpAS3ZoCPxsT9j5HlWB0w2K4KPQtrpwL59OHe2P5NFNq3H
x20IEy5ZROA/v8MQwUBQfXShfb9NjTvMQJnChk2geKtQ4ARm5cvplTi50/7vubhBGoH2wiEdUsoT
oDlFfngXbxIfuXHPQT8W29oBdbT1lmB90G5+0mdDUF3HqG5xiqL+E5aGP833/8pZmPU3Zjz1TbvL
Yw77aHHbq9coNt0Y3DHeOO+f/dke0p/4LngihReNiAx9o59pLv+dJ7Je07J5jIRa1B8omW2ikBOA
KvHwhssnbXeiFW4c1J5V2cXQPSJhyX8Awxu1WvlwEwjsrywNZX8WKRgx/ynuTZxCk3X5NRKXd7HO
zENiPbxmuO3uf7ueDEe9HGD1/Wi5Eyx96yjS2pwHmsGxpq8GPUHbl2BCt6kaYitl0nDsMHoHckh8
W0Oc7YaZTQ0npdcwaPW3qp6FS0c4D93Ho9uKalW4NBo7kNBBsq6K3Th56ASS2sa3PkE68zFwBj1X
V3KHfNuciMahgWv9zWHQYafiZW+qvQnRxTUN7V8g5yuy8Kif5Zvo0fYaNcXvSW3yoLw3zKlfox4p
nzgp5WeKpydRESAoR6HQOUd4UmtIIIXyNP3m+slprOTAM+trv9r1aKIxRafLvF190RPXO2eYYAYZ
9LM4WdMvZmLp91KpfqpIv24w5dZtqV/MuK5ciL4EvXTSXYXnNpAPE2yMj1UbbmNyhJkdVjujCi/g
Etqivz5i6XLhCXYd8/tOEAmKKPcZBCJUAwQfboi39fETb4ZDC/m9YDNAAJ9svgX08P+iOCGA3kIh
5AZ49RK8uTcX//Sa/HZ8Ql/lSmE1AfRIDD8Q+Eyacdv50vkOcH3TtA5IyKac79mKy8WPgEXqZTeO
tiBwq74JA0LBpKxKlKzxZR5IGmDjI51O6u5WxT8zHaWmxSERyr8dWmS2SEjSDlsUu7Wm02tkPnQ5
Cbxm0ntncTwqAEfeQO/uHQbYQJK/Gv8Ev9PiLITwIbPXk/XQiVkaN/7KFjqpNg3loIL3i7uHENdE
8qTwrcb/atcVXAcWJ8ZmjkseC0MaLygy8h8xOyHqEIzuqcdIWLOFKxp8Smh6a8YwIZ20/S12oGsM
t4qkHvsPnHWoIqzT21m8jfQEYt9knJYESTI550HwJY8XgwTITxNMOL7rOOsztKNDTbEYrexxzI4d
gxi38J5b61Uyushvj3e6TavqOkHzBRbHmnMafZlOw+hkclCQ+psDJkidn+7BGKjWpeU7xPW6Um16
RxSGDCsvAKUDDfgJKiKEF+azwOQ0VHOYCayStlY04Vpyl2eWknGDIc33t6PK9ZU+9z9htQGgej8O
NktpaLQIxvuyrZwuMHqC7BHpYwX59NrGo7wwwvceA/lTbzrmRuEYGi7rbFDweYbGkxe62OAJutOG
YqnlRhyZkK/m8c1j2BlL2rhAID7uceTD9twB94yIev6BLdRSQzfYCdTuFRZKuy/Vo85p+WO3b02l
yscDmtNUmOJKk8pf/3Fbwbo5u3258parMabJpRFlWMhAbpZAvcPPixFFg9NxvPBcfAOvWp9us1F1
JwdmLSLaXZeeLwya3qQtHME7WiEqdZdkza2WtBamXdAD+MfG1EGOjgjdYUkhzOmMDKbB4+GhC5O7
UDMVZKzc7e23EG1dbN9xFioeX2BYRs04sD8AyumfMdlpgnSy+r2ZB1v/HBGcaxKiZDO7dy/dfIAN
jMfhsPVowzNx5NZwg9clPPhwSeABWoEV0HfqAquBsNrgYY3kOJVHDy1Ynt5+oYibh695qqW3VdxO
t6VgllarTU/k2tRhVLhOkfi/PUxBeK/fYOkJoViWjikAQ1w5K7T6jGOKrrrOq9L0omnS43UMTbNS
d2QFuQj+hK0kmojq3/K9Un6LaHSa/cZAD0XuvKSEz+seJEdnj6WGbTF+uq1I184wZ06pUfGTZ1Y3
3Wg7YeVExaWijgODdrayt3foVS9n8g1sX4ZqR0OMBx41igvuu2/8k3ftIXyCCaPQOKWn363raApJ
AocmKpP1oEHJApeSNVdold9L0ZMr2bqPOCDhzwtdvtk4BvZGUXFBF5vqO5/Vrkdd7WpZsIWa5ecE
Y97/xSbXD0VE97qHOD9wfIyEUlqT9OYMSIy6A8R0YciwSNONBNfTB+FThYGLXTdVC9SnHIGJtIa+
2e6fkky4EtHhM/QI4w6A6IgIlP3dTM2iB4ZB6mIAEWtlxkORNTDfOCPCEVDa/jX3pEyn1OadJUvV
YiIqFNphcHzmm+YjhBevkFEyARPc7riMUrMxiKujt2JpAucR99YyWWZTOnIJSbvS5PWniJI8oqE3
HW/hmSC9n+oRTuMGsYF/4/D3DgG7iMnz2+iRNBFl/OzJfpZrd/VfNW9MJMO43qR67qL7V2tGhl2i
gSH1Q5jblasvHN6rsOo9xUaehDyDov5CLiIJiURhsa0x3qnbdOJaEU6/UX8r8JGx0kyXiqRMf8ci
Xp26GAxMJ61VFdnB4H56wuE1aZkiwD7cInYEYfaJQHSt9pY6yYnTKEiTBdu71eS7Bm+bia+aoySE
PZnxB0aUz1Ir+LBGf/vFLk/b44l1c/0Zp4tYEVXurL2LbFC5cWHKEwC3e75eDahK0hgiRBkTNf+6
BEtT04YSgtRW4fIDSz8k+ppZ11AgeRhILkn7CKQhuhxp5nw98GfteLoUuK3KdlgwC/kCuK6dbGOu
6TAHsf20441Q75hHsXVArYiLf/S7L8noSQWiimNOT3wYJ0f5xaA+fbv8i+Ng6luTo/HYbwF2l1vJ
lRMdi4ZlUvRxv+oiRyIenscvuvYt1AKDe+RvAfsy3Ja1U1W/GneMAD9mekiLPK/1rUKJ/21rVv6G
0YcVOszPXUgTEXo5//e1FJPVB9b3XSX3AUZji2/q4ifWsb7oopwwKnwaeImKuLDbQJkD26FiNWDK
JYuwd81/2iGW6hxpy6ySQfczMSxevuorN/No5q0IhwzX33CYK9Xyk2RDzWPgSBNau3YBAUcM0Btt
E3xunTGwfE64yfDMYEKKCu9YrA1Dz4FhXAWN9MoUqO8Qw+COjO0w73PAxSTm9O17M7QUpuzdk/He
RlokpjissXWoLK1mMsqV/dv8I76euzOfLeB+4xnz238cx8scqEIqY+nmOgAI/4IRMOaaZoZs9iim
mkZvvInAnu34NA8qZySipUk/0zK7ZMOYAGbP6Tpt4V/kr7jh4XpeQCuEWbeK4SOc0WjEzeN7zKwI
RY2L9cBe9Se2x3PxbK+xuTicRPmXYjtbqHKNS4ymKA5oxe6KH0efMVjXcLm7cdphfPIq0KyPnwSV
Vuk+oWtzLZDCMhRJBgzC+x/DpRv2ss83tydqSWEqjS97JufEJLnkwAhqkISvHtpVZiFsNo6ZRs8Y
a0ri7+5rWsP6bTM6dyJ4fIL7du4tI3isomBJxI6uj2LypFscVDueYwpRhmi1hsHspvHPgIwVDzap
8mn5JZ5z6O5r8CcUm8PsvPdC7A0EHuXy9ESbibypRxBq/BBGTeMyfAonP1+gEfSyW60dZSPwv02L
ZPfEIeUtgt29Jp2Koir/v8zuVz2eRtWlqZA1A5O6qicrj4lFskvcxQTYd8FO0mp5OW1xt3kiKYU0
ApE+pa/R7+jK/KP8UXzYoGDA47wJ1D40D1FL5t24lKzv+ahfocJRc1OkLe23eBwESrSTv2y3KmAk
JunpGl02lYEVQdTGgJiObD4c5aVRGdSXM8w226/yVDhIsJ8qOBqh1rYwjAOL34r7ppPHxCzKAD0H
EOJnVV1dkm4H6ejTVOGIOrtPEMoriPO71iPATxuEswUf8bY7R56U1jGZ7fHFVWg/3QRJXbbeeCnR
BcVWOXu9DTjyIGgNrMVr5Bx4ueHKBT3MyWMiL0ysQN7St24Uv1QIvB52Sspkl6ruJwIhoS+i5k7c
MoBi/1i8I2FmCTlbC/eTaSwUiSeDwaWurp4pFjHZbdn5Ki7zpP2tjt6hTPu31m0szQX9ZYIF3tQB
0P826j+1kQofk5BlZ1nTOoN2kM99IJ7RzHrfwLSh6MruMZ+SZ4gPC2niG0E8zGpuydQ6Fc97+itA
0HQxkHttbBk9aatRM0nNahyvHwAuQ4XP0IS4pUJ+O9Mg1pwX6+wsa6YDq1PBCyiY8BgnHg0fezWa
QQhZa+Jk9DE0xZJdqoJyReF7c4XFqou7qNlG1s0XR8Ef4Zlh8Pprhrq9QNu045mIzakU7/DnrJbD
4bxGtHLVfg7JJZr8CJkGyPzp22I9/jgw+wWLWGVki1RZGcnMrnuItd0eZfYovEGjeks7qmCgNy/z
bzFOdjudDE88qWO4dWKoCekig82xUhvyCfm8ZtRbWFE+i0Nvs/e7Isbq4mCuo5gxapV/o8Ji+QdQ
CPlC+DwN9DXgRLNMvLK+lZAixunE9CSQ89Od+kWBQ10gNOTTQa5dvdI+8Xi46vS+KwGfRjS+yINF
EGD/yI3oM2zi/D4pMRD8J9MEp52mHiip5Hzup7JjpflAcio9exEnv2L01+I3CyoXlc6YK0lUwUKj
57yjytMSkXUgoAtsAO30zf3cJAl4PTY17oVaIauJ0n6r0r6lfN7jMRGBeSJiCD4uJkFIUq1u5cL9
rFFCC8bnJqXdfQqsfEiWadj9+LdxZcKdcVXu1uBnTIxjwsAV5Kctt9G2GeI8c/u/rRZExr9uyHFL
hpyNI+OP7pmqaMsBWSUhlw1EJ6ANVS6G0bRfjBq0C5S+GgMRKiT0U3nwKns5mecX+SSMyt5gBMT/
3xwhNLR3ykXrVy9icp1ZTyVam5HjxXRDJt62G7GrHXjvUuoiSnqPCkyHlecX2uhRTOfL4Siat9Lx
9dClocDAV+k4fdpoeGx7YvEKmgQKSccQ/Ib3CnffTUX1VzTn7+H6R3tNoQ9m87R4akRb0MyAcPhI
X0TcETomNKw5xCObhofKx0QK049qZxmGBrfza2tFvC6LHJ6ymG1Q3DTaTdYEwqk9J3NXIdC+QZj7
ZTOta1pqIkLy7q+Mf/Pk2kMbM/BTyPTc9iNrT3hIG3RlhQ55orMJ3KN6OIPP0m2C4S01ALGJaMXF
9TTejAG6xPAZzoo1RkyJa5jtyWc/DF/q8hHOa4536CunRWYazRfKEv+Xj02UZ3gjrVWEoBojrgc/
w4YKTEqV1H9pys0J9bTBewe1fOpS8p+y+xb2kQlGUWlX3xnW8dBjdNQjoRmcsuEVUGz183dlCiO8
6QV6epI1/FvFl+IIgTeqNhrM2kZuDOCB81g7ucqT8uMi7HnOXLh7kq2Y0tH/0OaFIBF8QzIQw+d2
kOqMllQE/2Rf07MFhVHUaRDSIutyPsR/xBTB2KjLVq8L/kfMGckHryzEmFzzh5AhMvTSeBV53ASA
jpUBZt6A8ZuTZFGjg5VWeChx6z7MOXyWCK4OHae2WOOsX6bMSJGrfKvuNpLGESljbvfr+Aqxuc6F
knKQ15IM743tc16K4SZwCAgbGNh1zNzb1DT5wsFGVfC4FyeO40TRGuq3cChrS79PmSBPVSUA60D5
j3JjoKH2Qx9KglPwqm1OSRnoDyl64g0/EHEnyf1meiKJPaP6IcrxYxvbLyh7z5/8GWUEKshxZw2F
oAEMr/jKG0Y0QRkRZ9KfdJT9MTIgbPcMQ2efSTibGJor4L7OsO0hoQAEGv193GBniFu2UvjYon8r
FT3hq0m9TDMUQOH0c4C+6YS/eKQC5WiQhl3htj9XLsmDFDXHplHXuch6lC5t1xo+KW4m8zcBT/VL
paenTUWGrc+MxYZeF2ZgqdKqoglj6TPSatltQ8KJSz3ShQW+zXKVXPaUmFpyPNrISNhhOfnrMPtB
GNGYL61X6SFqK4WxZZ/K9UqG2lKta7qSR9d+qH1niqR1MNSn+xh129s1wFqmtVLupgFujBjYqZVp
k0CbX2IOmK0czW85aLUw9hIPoWnx2wghUhRIJeSTwjMd+xHIFnoGKGJi/EId0eEFcA5/bOC0wmmJ
DIe2sJA3l/LyL22aas2QVEtYEAAn+mOhtd/tnNqonLQ9qoLj7mmlkvFhFDW5N2U3ryfAiMcdMQmP
T7QMgdZlAzqlzQKCtx4vYAi1fI/9rVs1EvRBOpK2Opx7q+kW4OoKiCz7rRK7NJdFtfZLsQY00EkS
BXH43Q2a2SDOFhlydF0PSZDqfGWHNBo13nnG/XK62b9lWzCW4L9czbObGFJjeqhE6MACzkGdyT53
E69L8kDvd5ZTXgpbaWJx4W9nG9I1vkkNzMDBVrHSLOfcHi96fEQ2OBrgv1DzW0TatPp/ONRis2Mu
AWGBz1vofDYI10VxAHkdYvtZbz/9ErrbFvcTlks0m7AS8nQHP60nF3TH1exfh+796t2DQWTv2enI
sm5SX4yE4xOVEbCLLDJZQQLnTcxwgX2Sp2krq8NLEjA5dE3kjMJW4N2kqSfONhuUm7Ni6UwDMncF
1HOSSmNYGPA3+utvHQV2G/+TMh+jwTaMnDFQqEUL6kTOWSqyCksZoca1KCAtJjFtsO1KIOvPG4VY
6mj5sFk0BSbMODFSXYdnSYr/4EpuV8e/oSASY3/CctYWEsyWy1fVF7SruQg5Hl57TULr0drhYAj4
7nXSgKk9s+ECzWs9nQeEKSdYdAXCklO36eDwsKNskPc5czM6bahXhjN7D3hENranIb0jhxqguDI9
FUc3zuFo/jROrA2jVD6u/8QpgG72S6crC2Aqjk0l3fcsUIHL8T7DtLyFgR7XvMsHUZ1NhpFoZAiF
4p9Xg16CVUbG1hZ5kpowFtas4GRh+PqKodKHWJFj26pM2/qxJTLXfBnYD1/FG/8qtMhscPDhz8G4
Kv37SOzLIJYOm2fr7hnt9eELCao2En+m06TVeZY+Vv069VVpXOPyMJVnp0QmCCr8q0rEMmyx7DNj
t1RkVlO8PfwPzAvbA9f0ZYNhcpRAPcWmBqyPRdmn2F85KJE0KZx6omZ1IkVzt1DBFcfaV0GH3c6o
jF7vLKX8OEJ7sBJgtJind/lOXGaL+l8v4xXokO1Qx1LztJrM2kn8zqtnhINJwS6Lc+LiajvbJ4C8
3oe+fEhTorxiE2FxDE7YnAPcwS/QzflwnUkPAbsbNrhgYI5Cd/KIXFCKHmGzKWjs46T3IAOLDpek
3m/cfCiokCR+eayb8/rMc7NKtrWqGuuQ7iRoN8Lzlae4QA/8XUUzSuwNrS99P2KmILvdjtL93E1N
lNnN1xm4CSfF+VbmQfqM4iPhK3UqLGxCJcfVkvxnOt0uOl9l1lcZXvIl5GG5AfhAk0GvYvfVbIZb
s97Zusc62bEMoy2pvWf/7/Tga7Im0UOlAWFo/8mlL9KJFx7NtCO4LPNi96/smtHx8aH9fsoF7s6c
7+DzA8vlmXeRhF+z4aA7j0IUkXmEv1E9dc+22sEwqA4Jy94VB7q0ZRTePm4caOqM9k4mv0WMEvOo
ASjNRFY/rnR/rs9cAkNfYoyWl8d0xg+kLHmonXSin9i/ICzTLTSNsCR6czLUylkcrEGC3dZvlLu9
nzGSy1KVQ3C4+/wrsPOQHiVQPrJxbPiDJ3O2pF/c/LDUmhXWicJY02iXlZc7j3UwUh4/u7SZQlMH
kZQTq5oI3+vDlMSSgofim4UAZ1Gf0ce9T+U8IyaF2nTIpPY1O2NpYNABbBipjmaft2O0QcjMmorv
BvC8sFrdFAsEslf/gI+r8B83H30vQstMcm4i5zayLICAQiU4gQ687P5Pq27Xy3/ZOcs6Msl9XmVJ
MuyBlg6ciOCJ2+wrlkW3CeAZgB57vZ6hwbyX2+5VUopVkm/eqLZ+aImW2YsMN6rjJfccyxumLb+9
aYa5JQIwIqKNm/KmlmY9TGS+9+jjrh7T9h8N6rksv0cE+dwvkGFzeqJTMbmGDuLp3PC8ZYQG8rRN
kxJuC0CtgEKrWOK8P4dZfrIB2tcZc6/4MBfr9qxhXzzaQOBjRUeQfcTXfXYIpr1fhz9R1VBJHCNY
EtRlmMptLu9fmqROGQheN22nSNWXOdRYL27bU7BWRssgshnkZbXC1tNxtEtSXfk33BDLVfsdJmZ3
w3ifVV8YUM1pM+V631Hu2NUdFwsHpjzsP7CK1TJUW4Ec6Ntpxc7KId0VA5JEfBzkdu/YyBvigTXm
EOj8uGWZBYvBX9cY7AwONuZr3/4eXIskx0hhKqqrELxObtgsTIiRdqTZIXpAR6chrbTFX3M5VDaq
pAwtmH5TD8t0HJ2wA7gqLYPF4b3Tur7A7ZHdO/PQlzzE8TKh4B33QjpzsktuzzTm948kjyv2fcO1
IipuAI9axskhVd+CM+LmUVQF7wzwbCjjOg92eqUCrwGXbtO1vOOj2oDxO/PualK7Z69WfpXlPiS2
lFu4ZgwBS0einydocWF8e3R6VCY2Hy+nWjgrfd6Al4g+ZEJAYc8Zpr/cqdWaziBPwFY9V7jcz979
Luz0lnZt6isUJxgPgHGKInUq/Gb5waV70h2WOtJ0o317H1dByW/Reuh2qAadST/umQKJ7EmVz0ft
1IePJGwAqs7FutBiCwzhKFzsiq+5+0JgUNku/GIw9xHgPbqhXa1uZE9W4ZdEOUlwKB3AwR/ijPDJ
tU9IeU5LF7O88B+L79RFQV0scAocR36CemvsDZrq8sK4LZvc/WnS8CPdO/qhUgu3ffcD/uc2HbXd
QhSlAqt5H2DgvQCOzjDW+0luoQOgmn2ywqp0pOTCAXOjAEDC+Yfa+GmXKeWAKDc4UQmwiGufDrvK
ilXezf91C2fYEXSLHYFuJCnbufibiyLWagjMDdlBmKnwqKysi8PCCG0RLRsn57JHvt4pW270ymeb
FvvFH+7yNTMbhes46Y/q0fccjuFnuaNzpRyemOrIu2+sDJBXWlttsyJOpKK8raEQQaZYA1mQGNZp
xgMrig1sX6WkuOOdMgk9GA2G0lS3f0T9IM0ptvdpVU0glksFS9MkdPL6HrnPdW+Zknq3jC0epiEf
JkKU1al/X2+3yxfOBLNZAG8GtQ19zOdKgpfoh4VJyyHJl/2vujy9vhiPnB0b0IOfnb2vIPnlXgLZ
TPfPH1Va6C3zhOs/3PYyzlSdOZ6W61DYqGPrEG/PNZ+Zj7tRHRhc8ZPKAlPB6sONBVGhY7cv+sRy
UUmAb6BnO1TpW8nsCrhpE/SJlzT+qpoGNicCZy6DsGvMki8kumiOiFi7tKd6s6L1/mtsQGXuowb9
9hT4Mxbj28F25hhGtjyjQM66k8+CBPDGZ0IbmKJ3fpZcFLoKRp6B7+F3q9MkqFnNBXJMrEaD2U0o
5p5Zp35MlP9F4MEtbNZkXCA3eKa1gaBRYdxRV3jlYbJ2K4mdHsAQt3RplRbCETwG1vptIcAd2xGs
rvdAmmHg9cPU5pwqhWQ9zdJrv7ahGMtGjjLw6Z4qzzSoz3iXKkSEKCqG+4Q5FZKl9xoF2D/dwBKB
bM+kpG9Zja7W5GyiO4nYN2VZF0iIVyTqoC51O1dQ4d7WsgiWc/AjEYW9SHEANAAP9F5EOrtkZuMM
eMDosDE1OfXNEh+h57wgewPl3tHnzrc9HjyIYeHZ7sAuQrYWIlNWf8gy+AFU8DG/KLqrposxS4I1
CBHl2iYg4HPFoLeI8D23V0imK+li1OHe/ELsxKFuPK/tVl4YDVPT+Udt3TK6cZuNd6qSgE6WyzZv
RMwWC3C1zni6nyegGOwiSduGOlrz1sqC+ZVUuWX18k7GJGPdnkMtRGAZw9uT6hQkRRdUR04WqXt4
itHbCFwlmN1avj0n+G+UsFJwkUJ1pEWL/oedsWbICT9M/qvQ+05owByZ+IPzjtTRyM/HVuBjTDTD
zH7H2AtN9tfrskSAAa9V2fBpZp8gBoOSRR+8gQmC+fJNn/BqIP0ezhRgia7tTvyWWwrEAzfyTiwO
mkDh75T77aeWnINcaH5xBqb7xjMXC2wpmgYmickkUdsDtntdt3lUm69tgfUo272QdI4eCm4N41rR
Q35W5b74+3+bSgm/IB7MBnpQ/CuMRv172ghDB88EoxRQdHvGbYiegfXcsvKJ6SL/A8cENqoESTMo
u1X0UPWltlQU5FSMIH76O4FdLttPj8bv6MLD/RYRBCtRBddcIKtccKXuZoij4zxjg+ZrIa79y3VK
w2T9OZGrA3sgr4EV9P9KnLsNFdKJBCqTAxGe2ZdL0N8UEMBCq5WFROzRMlA1tun5FBtNrwSksDyL
tCcaWnx1YTMrP2G2gmUYe/LP6i47SxqqcBaSVnDHci8C/F88XYMjyVmLQbwc+X4lcixbfgOTyvws
uwjMXVrSMiE6KZBKYkvA1eI4F4quTy2lHghf0lJjSEl3Ovwd6KIfyCd87oSAtiQabtQ6GWaqcsJq
cwfPYlhVHLNa1OkQNvSY68pBFP3lgGs5fnvqBHtRDJHzAr+YOF2gn/y6qIIgSm0VBeFAdx0zXbya
thJz3CD3UO6rBDY+bNsc2IT5DzJb2yhKdAEk2YaSLWifveUuCi8AREkEMpvESr2kWLVs341rZl9k
F9S++Y9HiWjkq3TLArldfkuSc6mJpIV3Rw1gF1aBB2jp09xZbMudz52qWSk2LV1yCUdN4l2OOkvL
ixiy/kIcaSnKYNc9UEfjAqzE9gRRqp1UUV4o22fMKjL8G+DXUY9AewUisA0GefXwML3kMSyMo2R2
fMSG867JcJOAWM2/xD3phthpXRdUE81Vg5uLHttlIEwI04hQPEhnZaw1fLJBDyup20LOerG4sfqd
wWDE5eG5VB1qrfOi5J9rvJUY6SU7N9B9qetl1zuQuCBtPMHT3C32J8kmN24519Tb6bIF83WtdxHR
NfZvg/JvqU3Xskq6j12VI5JJaSWyGLtIzGYqrCbiNVUOoMmD7jCvSQQwfNb1a3FqSyypiRDMeyC5
buVhRBjUHWlO1qTaewtLhwRtwjO3Cn6rh2Ys2neMAXT3GHjiy2DWxjM2HolgSN3ukD7/ydKE61f5
CgtKtmRmpp2AfMJi12ONR8YWst+HdX7bhcSHxtjDquicuP7d+IIM+QLx1nN1PS8V6lU8cxXl3soM
u+nDQLD1crJD4pPuMUhxMjqXe138bd+dT6swwpWYi7PuTvewewB9/hTioJEM+TKpE+GPLRcrT+wS
LYoMFVvGXa18iruqXGH7OzKHbFTEei43mLb24H8q+sodaZCIyVFqZUSDYalZSrfT/w/+eFaZjQKY
c1fcDfxBTlsPOGaPGNfoOQFR1x1Eb6oSpwQKOu9JBtCuOlqBYxMV3AsiHHpCCDD6YWizw9vHQ3jp
820JLHeFM0dwwOaAV7byb9wmBBBTzuIFfuAOS4smtFmnFWE6cVDZAQ13Aih7AASspfdPWNdE7fiB
ka99P5EZHNzs4jhu0Qt+HZTZqlv7NW36NP6kGo9hdRZnMOZzJkSyJGVL8taKzm/ZTb3A141qywGW
P6FoCzy1GHShwKFmCwiJpqTwVfZZoknld2HOwQi/bGWsoOTNV1eT0d3nxNYdQhAhunNoGKl5spOT
HQRV9I7IepAMFZ5PtrqCTHCzFNmd5egsBslwCLWeLaAQK3rzAYDFeIdIVpeswt0Gi0wFCsfb7lIJ
kIBQeydUOiU2pSbwApOZa56lgiaB3xLNYwI/xm+0hR889bAHF1+JQ6wY2qrwe/oPYlKAFgN9IY/P
CWfvPcXvHYbNRXw0Sk8HccFe2H2dM+greU1kLoFYodGa6Cpxp4kIiHtr9Yhq/QzukHq0WBYj1Xjx
RXl9WFyyvmwXvLnSL+1RqZ0ztTFduml2BNAcMbVorEFSBzbfqbjXFw5jQ9xyIBIzr8GV7urTiDAU
hcduVllsef1Q8gfO8LWmKqnH0byf8GZKvXh1Ki7mzvRD1xgBuvFf16F/VGuWMWqkuG5XgfiqLh+Y
Am8tfrmXzHQ6xWiPgcm9j7jwSDKgC6ieWgNoeMARQdRlCqM64rd9KSYsK0LyAbwHa0PyYmF2o55S
dw2AW6L2QcAgoflRzLzWo+C7JxL2ub43mpUij8LKLyK4KffBA3MCt0uLhBJHw6dv5mRv2VvMI+bu
k9EgMNmPJMcP2bfyyeDrisbIpfgVEOp5JbVYBQDGWM6H7bWtylJtAKmjXQhApdiB+OwG49rqOGRr
WpW3YgBt1u3YGj0gK5kkPGmhVpLYEaDYE0GHQgHD8cZZbNq5MMd4lg8ZKeKhQlteXb7hpGcCI4mu
Rv9lcEd7GSTQ0DUvUvgNx9XqkhUrO8t/q8AYUOxEpDSWbkH6CIBkp2xwrpsQybCTN5pEA9ejyZMB
Ub7hPahzwM4i8p2otRI7BfJNNuaRrTPfulH6Cin0c3278DUJKXqEYVkSRs3Fav/rtWeAoQCe305l
I0Tsldugp5nX/asc6MVZjZ9bX1woRLKpKVpOE6SOSP1nJbeIaAfJAhmjILpfbUmISQZ+vxtL71J9
cWVS4NQdNeZQLgD0b9Shd08u+Ottr8cQIRACOt68B2DUb0ngfsMNnzxro+8IYDutRXkoteUoYJU/
VnSjQewQKeB3pJGXFw7EaYQwauT9PhRpJxCFOQQtQzIevDxbJddTOT1Acf/Md2s6u77O35v8PRmP
DfuGHUqPYpxzaf58Yy11eflMIKoGhwdwVLddfeVK9vqkg+fr5dXRfLw/QXasmvsSNm95sjmrx/cE
xPpMbldJW5RAQebBG6D/AIa7lxjFpLH1HddFd/OrIIsDGCBzldJxBdq3vYrp3ejQdioHaRRPfe3T
5W6OrgEyzBNsppae59elk98LnBdm7HObfjkc1pKF/PIVVVmOG6XJu4UzHuZqgQLM6kXSwF+mIuwr
BnrtCZTFm2t6/5fHzkvCKl2hciw95nS4qUO1vXA6wLBdNE6heuscD2B7JJNGKI9rLTo+6s62bjXv
v+ozyPuxgS7ThMKKGdIrDdMEBF5CbsscNW5w+PUpy3q0xUWavoVShCdd+rYH5bDjcCSyxfGJQFaQ
NlwFxeKDkxSxiEc0VLNRHARn6Dl14btlAB5HG2VmLaGU8XNbPy5G/DuSRl47xlHG6PdEiix4wxGz
D2JleiuQaOc08re1vMiL4IeQasiL/1dlLkDaE9e2cQuhRRltvwXZUT9aPziWSJ4ygveuOzuzsMrR
JRQi7mEb8UN7v7xsTHj8eFs/iS6oTRt4PJTrSotXUu6aKNtauyfKDsOndROxH3azGmXWXMMuCWXU
qILb1VBnIJDl3WVGn908u50PzbB5hPIqLlMOPPiClPfYvBdSML1ZdhR1pzKVW+esLDCNV4zvJ34X
iGdQm2wZ0CN6azKZOIToB3M10e2JieJ9hqEcdBM4fExQXYz2RXoYiGSYOoP0ZQ0maHG0IcWUmL3w
RicEJXf2RaJTRi3yRKCM5eV7kUwZr6tzTKbM3sc7EeRIp6ehHkTNx3DY1Gex4vNi/7PLvOiv0mpR
qgdf88MwXyKbsKU7MQmZXkeK3sm/0ZToE61VLtSNakex3jqgkYg9OY+fq3EcT3mRS98+zR+lyELI
7jfMu1UMee+HzhbmvLF0gY2YZs5YrUeyjM5P2xPqxexI/3kx9G9DTiZ7fGgc5GP+Z6OF5tQO3ufT
WqV0Rn2YwI0ZFnicS1jxhM/LlgxDBEyStMmplFL7Cy902yRm+eur8q99UOMNLdyHKC+2nFDUHmv3
8W5xWAnWh8VJ5D15+yXtWixj4byz1TzLKhgFhB/6Z+lc8rhE5brAeQPXjQS0DFGXGMq3mKNhX0rv
iMxUSUlGYBeYaTw3EBQ/uHZ65bxT1PtDBEP2xC6mV17pbukKoIst6Y7nwq9hr9T0GHxjIy+LHCsw
Vvp9OyXrTbUAIna0zC8+2jCeGVb2HK1+MIw57qqAuNQobkwus2wzqFhmsw7XiJW0YHXkg8ZVj3GV
Pkyw0Fg7Jr6aeANafV/vkY9rxJn7HvlDfzosCbXMe6wgQJdvX3vXtYmKEfOdZYkCmBMoPXaaayVr
Wc50SdmqRDCRG2+Blizx83w7ybH8IsMNXbKlz8TFZd4nSMtWEzwGTR4vRroBZ84ROkfmgMh7jr38
LC9QXZhREquEZG8D5KdN7BGGEqFgUMTtq0CfjONBfR89HqU14L0ztsPbLGxX4bUDNBv0zrN0K28R
UGlBBOLN1xF0OXvKg1FjtjwLLMzep6FNrYTDnS04zWoCDAHemhSWgU6REsZQ6x6kHnzgqI/3zrTv
QDt0TY6lMyUQhHUNYHpePSu8EIxMOj8VHMOCQ+n8dTQPxoJjraiVv7iVdiHS69dUpHyNwHSFhnTR
uDF1/dpz593sp8crxIl79nAdgh2bNTRxqZfXCCwaPtlH17+4LL8WDsGJKyvucbQyg74mReXdc5Wf
PDVogeKBfNE+QkTjDn08iQ4BOHMmTKxKeLT5vH4YGmsCSyl0erf1WCzyR/A4cPQBcKEOJXRL91mt
MPxkL75J4U7Y3np0D5AfkqwQBj9OUm8Xpk8+nTrTQNChLihMwrttH+fVUU70wxv+zp3RkojGaje+
Lr0Uc23caGfkln9cwwSWtvq6xjL4RjuzW9HnQZDS3XkTiEItZEq0aa3eKzXO8XusqYmIBgOEYDUT
JeUGEJXAlfpQ1OtmAgxeSPu5cxtxsBXwZlpTRtIN51hvLpyLDxSI00DPWzEKDM4Mn3A6TGkaiwap
ncvc9IEAUsX689WQ0hW5lFqUEi/30i11TqOgywEbOUHhhG7s4L5tda0+Ug917AytRM9XM2+QqTny
doHAIRUY6VMTBChUcNx/B+looW5ivMwR4Hrw0bxP4q+msB3QO0wTe1wYgq1qH/wpXwUJFG7jrqs/
fKhn3JzBaT17MWB3vU2wt0UsLZXJTM/bvDDqiADqNpBz+GEiwOKxpFbvAWUsmdaRWpSbK1YG5USZ
rDvsIC5zlUwMsW3rlb3scgLHH1KeTBHZY1ogGpAyl99huFAh3569AFNU/zv0mdTXr5koBdJGKGTG
mVSX10v9yvCRTB2ncQmBLaoVPRPSufJ5bt/ylLr47mjJ00twNI3FRd6aU/WESOuqcw0bXcm3/vI3
2sMXtaqkK8nLQR3hbv9UjcCGrQYeUbJl7KkQ5HbIkwqUftcjDmwfpLyUPYquSqSNiRDgLtgOeC0+
TTaGn6nY+3kWGGTF/M0EbkVksvxzymUAtETwiONonn27JOBQhCINDdW0/jOm9yJkcdxdMB4LuniD
5WcC1aeoK5NSC0sLkN3Nfx67pXrZiijz+0ooIJJjT3UNJL0jdBpGBoTzpKw4lLknEMOXSKp+zPyf
WvqwthcyTZbi7csOJBw9Ba+LX1hAHBHayzX2OK98H56ZXlYzPDKHieTc2TjG9KS+Pt4ZU1Q5/kfi
+vQKnV/ubUzBK2qYXJhQpqmtt1QQ7mJ2x1h/XazrEH8MTgSHtjL13yI6EEE+GQdEw6vovY48UvEu
R/nRpP/rWgAC9IdlHUiihR9+glZ3Y7kIC00PQfHL4UcrP4uw9rr554pViL7dbfUDhdjDAZyurzui
GXM6ah/Ji+WhcY5CrhTKrKIQrIpGTjnaFkOLP0iGFaPkilLGZmSEoBfpGrnZ2qrmoFH+m19sYg5d
8w8uYlEASLMrjKTKpVnwbmA+zzkcW0byZjgoV21fUFR8shOd+g01b77S+4VZHVTXsYGsWcXsBek2
8xYW/Wgz33+lGkfmj2fgupe8CqJwe3msDeAf5NtkpdPOcTnvtR3+UXDJrJjC3ATs3ddtfs7O44n5
NglTcNxSn7PZhfDCuQTPFF99W+60w1OMyW61QkOem2MoIwQZ08e2+07kk1PleiiVOJnblCp6yBYq
JDCMN7EW3cF593W6PCKycW/bcSaFBmGJSdUuwR3u4wSSruUJfZZ/odwi9RHYFLTe78z7pWxhk39I
4eUXgoBlgsj1w5v/p4c6EwnyYmNqhw6L4jo0ZAgbZoK5DBpzcGVTguEv6n1vhEnPrSmOwZmp025J
zQv6O3jATMWsv99DyrfOuVZjsmJHtvodalRE/2PbaCLUEHNRpYKjpGdGzZKELWvgwWJ2WIfRDrr9
dGtiiOXiFXf63nwp+0Cu+IaiYACABUIeuts1Hp123Hm8STe7cttZN6nbFdgxp/qwikMgC3oiTgB5
lcPAmtBNABpzQsiHJmMvHcJUK74hmQyF/ot3Ih3MGoEFsxWXLB0WzTNBPEp/K2Xc0v6ZMovZgMC3
6gUVHCcXVruRh8/Fb9yM64eVQTXWeVCpLJMCdX04dZ81gSswnPKYApvy+AstyFrNa7DvRBVYaHPk
rAcGIfukY9THYG3mXNXzzO6QcqIqfn8kbllpGGw9xWDEg+fGYJSrVocrYWLbr+rasSjJnr6iPrg/
gEh0TTFLcE3Zmf+f/PE6K6kThm860DqH1PMvM+5red2lwGqBD4PUbJ733KFk5o6Kq3rYEMRVRkXE
cjbLR35t6XIU03c/55tZtCwaoFm4lHM+XGCjlMZ4CLJEpdzu1WeOoO86VMPls1ZQfMs2esVevzrj
Ff2Qf4zezSgp087isfY52ukVDcAVxMBTMx0zmhlCuTEpYQZM8YjvEZRuv3O/pKZqv3iTaOBaRR2M
2EBuBwjutJNK6PFb4k8cq2Yf+rUMYRz+IcqtYMoVDtVFuGrY3XU9QYA9w6eF2DmvxefnU/jb5wd+
Ig0N7Ry+GLXcnB0aWzuztbKr7Fp936xhRqwZOjPjJPWicIIxxg/88AYHSwGKZse7Ud3cVOoQ+5Ve
ANnJRDZwJeYDcq+ecKz1FmSa6TIb/yWmpif64kCnAqIUDAFRlt8yER7dqJR6lyHYifOEok+lSnDc
o22nezBow/62vcXemdWfoWQl/mtys5OhPgWGHsHOXNs9lLu7mHc3g38Lq5gr9jjE5vcIyBNaRP3Q
1bkevjzHwjvJ29FuB4BT9of2uNXt3adCIfDOHX7M+wYYdVCWgi+d+jgdKXCd1S1OLJ9+jIRZ4tdd
4CQfTLt74h9BDFGme/CVQ7XZhyFn+n+3nzibc1alYfkIc1GfJTA61XlJikeasydr90XJV+B64NpV
jRTzwWamCL0TS85KwCY1I1QnspmKkQGKTS6G3Vx4KjXaJLMF1CcFDdWEuo6RjahmleG0JxnJrtn/
3Du3vHmzKXaKT4HJqaMBWSY4yaBC7Y1T2gP0G22+mnlvkfTqDbQ1nYojRi/gHA0tSYk1LRCJSQlB
CPoTjI45ILy2oKDyKUWe2gzplpDAyc+tJb4Ag9AmmTBxd7QuLpgwFZ59bLIUB1UH/t1pt+mV4euN
Ei33AdJjnt3A8wGxREhK8JsENeyHyIwUBgHuQkeSOd8TYx66NUy8lx03WPbLknfuNKMVbdCrESqI
xi1zzIr7Fm3bLtt/LKbfPQSGP5wng3CkbUi0CIla1yicy2HB1kIn/Zubut0zA/3OnlSREo6lsrN+
4Yp/Xfkmo2UDvdb75jBSkNiVmKkHeCXVRZ4gUq7AORWURtHIFhQIVzpZKbVY1EgUiOYsBgQINaDV
uLSBkUgfhQN37hafz5Q+fzNeV5J8SfU5BRWrLDmoA3E3NZOrcm7CIA6fNHcY4hDcJpKnxreMRJFh
FnZ/d4fzO5yBTrTXqdexJ+sstBvPzNllZ8Vj6gk/Z2INKK/CWIa3Qz9UwOogtfxoypYq/0Ga7pEX
hzo4NfPRwwaPPUS4X+ZRW3igxUIiwaigrlGXWeO02b8ATPPlDM0gXjEDC6R6Y4erUYUzs8TZ3n3W
/bWAlbE2xdP2/bZAsp6bXQuUTarMfUcgDDd4vvy72dGEa92qqx6JTecT1/Lcj3qoy0Df0BvtULm8
OnVvY1aqC9CuwY4UtPdGWN0hYMgLXxLD30rCO0dfxGe1Q7I8vpJPin6VqOLyKU6lSuRr5BLu0Sq3
quEynRnAGI0SHnLAG+QTvpcSZEQCOoniXNFsRpyK9xKy5PH9aZgxZ5QkywJuUSVk3jLy4uQRGVM7
MAJKOodpts+YqFYqvXb8Bf9Olbu1liksBw94Q9tH7pZ/KVtgoVOUUw447SVXPdNrbPV/TKPjZJhJ
YY/p0nOTKMo9UdmLDSHsvDbjBWVjNLEXBz8NT5t465zRwe4YXUo66GNqhokW0Em87szcZVKQWnPw
OwxFzO3md16mzZ4zEURT5ng3dZoY4NCqlRPfTBKM2qJnvbvA99xZpjSwtS/CYfDetjn6SMpL+/qd
JKj570c4Mm047q/+3/bwoGWyqMg4jLQ1yEl7Q3KlCJs2dqYgngYpicEfg2EfuBxTmRbXXleHqldq
8o0nC8C3CO+newK02RrJwq219PD01jIXuEaQm01tOMpRLZheODpNQoAeyqW7KndBR51QCq2U6n1S
sDx5FXehci978ZABL0WeVtjGA2G63ZyKSZ7UKsN6y148fH2wHuK2OCyCE7jnC0Ush+oQs5SlaJNM
+WuPBgxjibBHEgnqwH2dCpmvMfVuz/wyLCSBhueto9XwsfONqxmpNR+6gjSffG+EY1XiWp8y/Vl1
kSWx37/Yi/28kQPn0tgw6+N4P9O7pUhDfRT18Dves3gY7LygX6OY5NrXrsIHjwfQS+tDSp0Otgl9
F+PyK17i5jDn2CvU/dUBQIF/dkmMkd/BWnxHtQf8gebflHu9POXkpFtxA4os8Cez+PSnNDABdPom
MwpayqjsUtnOEiYszYNAqPp4M1awbgpdIqH8EIgqqTBb/5ARkHW1FAWE6MdZk+APFpzGxX+2H23k
49MpvxfwGn812NLq9+A5tf5BdV59URU/P1c6nxSgu/LCurA2m5dOe4oGEMJ216Y3eKglfDSOi4gu
gx28a/cXhsBCM/7lnVKY9wJ+B7v+d3bgdzxCQgYW4TL4BxB8XmmW8jcOarek5KXdqEmxV5Cun6p+
CtD0LmmBuUqF65xnDvq1+EIKEgLlyeH8hDkK7ZZncqx4ZRckxR7VMeUvIJ5vngsbCUomc/N0OhuG
0oswroqjlwQ5l3KPhb4amikQKHLHpTNY5dqgQpbt/7hOsYYJvrSVrY2G+f8U6owWfDA/+iQp/qN4
biprloP6cfyAJjuuQINa9/H9CPNCRwalsqcENeHI2bE6uyzvpb1jao/J7/GvLbi31WmIP2klj7Yx
H0oieKqUNv8PhvWjIHj7ps3mh7EW9xhjDr7yDzh7Y1Ms21zMzGVh9tmkofxQbobWwU3Y9EI2l6+h
I81RMiN/RnqkQvKjHMHmwLL9FlWhTsrxyHfir0W4S/e5cQsZWW5es4THFooyfYWn9joC0N9C5zJr
+wYo20Yn29nLbaA7WOUOHb9S+ygMHqzNPFOkfRzNyHmyTcw5oUuu0W15d3gKbUuYcEIpmhlaSjRk
LrG6letD0KdRvi+Mf3bnePIiLM7v7YCGmtpyaRu5Rxwro6SZMkThC1B0Js1PkZTm/zvtduQIJniL
ye0EImzL+F91fwR62WLl9YV2VN2WzRJQw5owj3Ygx06m3/wly2yXmpRPnT4/Gp8EzgXR7iYLED/r
AbqtgBtmnJYT2XkabUk7Q/1p8jUM7w8mNMB+DS+C42bVFIkdQkLH4Q5wkSJ4ftXB2lTl9vGQ8ro9
49HZP6EiOoXeya5ymQXhMWtPH7IkXG5I4CPuXbXjPi4CY1z8YQLIGsejTxjWnXdMTSofN+6/mgdE
KiVHyN6XIoECWuB5PfD7DXkXeNNVnlnFl/PvvsZ2p1KusimC+qkS7kx7O6jGVVqHstfcivd9i8zf
MtbdochTekARzIu8f06mHnBhnP1Ky6XiVgNVuhhgEyeHxtwZOmykqG8FWNyhLnLcXI68AGMEMj97
XFKHPoNADequCPDDkH3FIEbwvTk3U469MquILTp7N1GMD87he1QRywOfTEbE5Or1OIiaLFjdSAaT
rmpadMDHEooonEVMeBilOxlB2spy2effpIfaZXkjVCVXMGMFQmS/WzteQGY+0rJVsmr/PTYi0o32
LMgrHcoAt9xSZAqNp7wIRd08/j2nRkkPoxSvrkrzv2meFs3cLeCxWmtMrPkislZtIvVPQ7BT1tTa
LkZ8CvJjfhF4voAqnCPVCOpHtCB/RZhAzpHOqKQoqYSKnrzpEbKkLaMLa+xA5j5XzmblT3ZJfG00
lRr23vTXLPnjVMDHkW4Dkq6DQLhLUWqTtNMwHn0I3ScaliroWFGP7Uinks7C3T3VjrrKpMbeHHbj
A8Ik7kmcEBA2fuw6+xCNJUJZXDM9tMkMf4Hz0dq5scpwbKooUobjA5OwY9NZCKDM3XmE90Ysn1Px
DYdW9oxCHok7/90u7gwd/UEWvbcmDFcxW2kdgbD4Lcvs7ZEGjguM7wV2AaNHHd0gzxIzz4A1TPvu
888Zs221iFy5q0eko99WVXEhxLLAvnjABr9UwaPY5NrFlSZfcuLPkr/CZlsr1PVAnUBmtR/hwl6L
4/L1e9J+yXD3vV1d0Y4h85uyUD+M/a0gI/Ez7NeD+bwObE2paNwC1RBkxa916G/3lZEYSVmJKI6K
y/PWL9OxljCx/spGEek202sEPXUezw0wLh2MBQTQbDIhYMNBsGetaeucaG+lL27BItmsQTvhVeog
NYdW+EBSREZRPzPMTFZggwh3UsSJLrUYXg8tgMQyAckYU8dcwncbwho+Is10rjQ4Atq6FXtehcuk
tXU5kmUf3o9D06bFtqm68CaBRQuANhL1YQ9QbxXVLo3W9b1NHwj8Sf+fPQMxIdM17cXiZQNE50rV
WcMQlNANzxRDtWM7PCn+2Y8MnRAWCE7Owr8yifLPj2zt2MPl0Mz+eUCAuxeaAWKpM2Sro9tbthai
389lCa9o5QJd/Jljw2jKIzPFyRgqHzcmCF5ILtI2VHxLR5sKAdE1Qtl6W8n6KjxvqOmCyXLvvnz0
8B/52Xdp8GHdcXOpzjhBUKnGGbtYYLDqfZtKMVcj+4B3VOktKKTi0RbFtqPpgjaRFluYiQ2zq96e
eGf401WY+9aCQdiD2M0tC2J0ykxsjAeG3A7uQvlhtEirJUE6yap4HgJb5qHVDtlmCKVEFC4BTEcf
3VsRHtXIL7D19MeLBBN2ViPeAfJ9BQz3aXkKpxzk54XCRl4fM8SU4sYWn1BAX4aWbYFJYffXzXQO
Lz1pWKgNc+yaqfmOztVcfyyeYtJ3xwVaFallVojlr6SmcAlntsHddmzrthGFcFnDd7xW71Ps7px0
pouFPA6Kc5y5GUEtMML9X4jwicGupLcvIE5rC4fPbTe2ypVHf46EYrEg1urGrNsP3bX90m9P3+pc
iVfIZ76G7D2DBABwPvNTepCSHYyz80SYkiauEoRJ0PHTHWASCYtVqVoDGi4DWToALDQ/pyz1ivJz
g9/9fNpfq2lYhV7BE3Bhuw6A9tXW9uowZkcntu9HVyOOpva9La8/96SU6+oXJNKQy3i+6fOh3ERP
zWcGsxYaYfcMeqHoV72ymP0W0cN2xiLQZttXny8rMGiQsgr2y8Y4hOxBuW+vCQE2Xi4zRY3aRVrf
+zK97xx71VZ2mnlj1Fo81PtJ+42fDmKEA2areOx27EpVYRcn+Sf87FTDgz9Wx1UEJNoTpDfqtwi7
Ukj55WEvJ1cB7s3UbqAzPbsC1JJcBf7jZYSNsHJObmJvYQCyTme5bTLHCaNt3eWIl7aZ0YM0Yq7f
F+JbpguzcvW47TDdyb4dA8GJjgU0gwPWNfrAN4lkbqPXT6rGC+muQ00tMdMkUeImZ5KBZcb35rdc
Wue1FGnfdNnRLNaKQCiFtWCmbx71fPgcxfUC/neh21O9ylQo1gSuZIlQyY6eKI4kS0W4v7AbEDIo
mmOQ37H4b0HacYf0PL40rLOElYL2w6obhETntX0SIVWDlLKfi9HhELlufzZ5wIi+957R2bWdkl3n
V840TE+TjN0BZU4dDzOmw0GFyb47jv0jjd+gpClQadUqSzn6NllPR9oruX9inpIIErUQyPm6Edoo
wb9jOOB5MYhJ9yJG5KRRnXh3Cl1ncy/JnSAYR5luL4804EI/RzWiyaHTllL08KEIF7B1vBgbIeVu
GthbAxIu/cKUyN9JtRwpRGJ1QV554GeOV0srXX5rnwkZk4J/TZ5HOUKMK84T210SdDckBI0dxf1M
WDT1GI/do6EUpUIZjff7Tr/Qw+IBvXW0SqeP7o7CmaSFQbEC4PnHqAJTQYIVnDg24G5P5L/sXoZc
8s7Th7r6sSZshrUeNmp2/2M1yJulpvAWbitfJqg4c09i9FBxz1SRgMSyQ12zLBXtoNB3CAbO3seW
w0kAZOi0VGPUorW0Q2A0lK4F6vmNmypR6ZhNdZ1KxzcQCzfcYhsQi1f5PZXAULo3IwJFnpu1rb2y
Gvd8UJGZgPkC6LDv/xBWiGN5wbfn+vWVnyoRdJMv4Lv/MqniDfseWSOYCx/XDI0h9fMHaIiGS5F4
1LWBY0FVqbIULJkpDtZsowmdUpH6BJ1NltUqWWAoZUZCVL/Zr9CQmY4oAFnrl3zPNyJsnci1cBGP
Dq5+bCn7/jW0Q3lvmdnzGavQB35yC3gtMXi4rClkKS1xbLU0Xzpgou2m5DkqA+G7MTHnvP2eU2ME
ViQ0ouVwHuVF5NvTArJuppsRHeG0Lui1vWwQ3riDcQ/pToNZd3ZbUHTSqU1SSizkFCmSnoVH46Pi
DmHNm2UPS5r+BowF9jOFARchMfCfR2BNEzVRa6QSQ8SOrZ9e4IAs3SOwRqfwPQvIO/meqX6n2q/t
PuEKbSjzSC3DYxBppRmu6YCvmQ6xkHPqxMqoPmkrNPsMEq86Z6+eQ4AwhfPgW3bgZzl4JjefBNEx
4rTy4dClh2Q8G1C2I02RKuqVTgfUAi2zZ2E5O8CWjnTcR9+Psxl4QPSfi08xXgc0UXUH6Zffu9gU
qzHxI5+sBoH6wSnQWRvH2l3KmCFexON7qG3qXwmHfgGI04mfv7lsmmhc5MNwgv2W/BBpyL9sNFPP
XCxjkHm2xg8Pc2rgoeFXEh5m3RInUCCDx5czcl6JdCBsm2E299gmbixZGoOnW1BS4d2xGY1eEtdP
mUe8JLElELrroeB2vrOw2CDvDXfh/g/cQFtUuy/UGvYr3q1ZdM65aWHlaZlxKM1+Si4unpNRNb1+
9DiqcbvanUK5zh0RwbTS1qcMl+I/CVcbsKSXeGud4Pz3OJYlCVjTacfnNKum6jiyMEnx59JrSt5F
tVi96fzqzks18B66p9ZxHWAAhwpwB20zIAHIkZIvdrlCF27PmPmy6xMV2ppGybznXSF1lGN/gOd1
i+BIazF1UZlcQ8VMCm0n+WO5psKUOM/W9N07asHZjX2yc9StuGnglN5jM+WukiNmANzOAlbq0IsK
v+O5YJtajMlFlVUYg1FNK0OUrLLy8jwtvEC16NTu7dW1Uo5TAPzaGdxQ6CbOks1cCqSuKf40CkAp
nS3JMwi0Nzno1iRJZ42cLJTCnP+OBj5/IBRAqIUfex8F8f6O2cEK5DCzF53+QT1h73YiXcsmfqN4
kBYSkHcksyoZL5t3VfJqHMZIMhDOo0PcskOmwLMPQq5d1Qn4lkSPUnFayPVYrcYcC/DnPunqgvFz
w5RhhwpDYMCSCfSGl5z/+WEKd/ysdxcUAr6rrrhrSWgiderqcvdhcmsD9dTm9srsebuDPKdSJy08
nBL0sNzr1ZG/Ic+Ri3l36ECJRtBz+pJJTHpxIduIU09Io2Qsk4aS152Rw7N8tdOgnfBs5ExSDHsP
hr+vY73haCcKByF6XxjO4E90i/zZrdvGsty5yDtfR8ocZhuK/jNTCOMsPR+9QxvR4ivLuel/VBvV
+2k6lG1x8zL0nnnUtUHddKNsboTBs6apbeU47QEkzSPZwpnXVdp2EKEHVZtPLw9E0suF8NGuRiUI
sC3kVx4YD1746Ok4to8amjjbJZ2n63gHnmPIAjwdWKg7AAuq4NYmGOSDWI3dzWapGK0Wbyis5qgL
hox9ov5wsXY3BmdbnQ0qoX2pxU6rly21KWKW28Yq2t/aILhI67/tq2yF34agYLpX3JYBPLHo902V
WoVJLah6sY9ZlDM7/zK58P+CJcI1Z3EeQvys2OR+fqUgXJPacee1X50T0FWIFARaJo0p8uc0jZC0
wnd9nFEk/miPExHlE/gaE4lqnBkDHWcBaxJMqy9jFDFhOtXg8rvEQEnwXFTANt6XNICisNMsg4D4
pIDdjt2jhlKIXBEb8jpVOdShtSV3HxlMeu9bxzWJtVt6/Y+kcH7LS2NurKrRtMEzZnPc+NEg1KPc
jl6snC1x4qpbeAsKkp+Q8QXbr7XyNK1JBeiaPhiKRqkXX6OSiY8sIX7gluXH0yWnKXpctfarFi0b
CKqSZpNWvRG6Is8Vgrm0bHBTonkp55LKREj4+XOKw4vk/xesZJdCk7mj9XI+b8bmfV8OfscWUPw9
Xnqq3WGYSbK6RiADmdKIvtNGe7hnyS92UdXmR4tPkceLmDkNwVFyTMzjYslt70rxHbwVO/98wfHc
oJWQHsysMf9+BaAjImqW5gAblWXNYPcaeEd5AChs4JiKlRewwAxq/EoTTfRiqswn7FuexhAs857a
Ki5MiBRGA1c47QGYwCc036F0pQABvicqJNrFIOyYRK2nl2f0qYpeRSZCCHD9OhNPKz03LgwjoLOi
V4X1/YBqzlZO0627BWKy2BloZ/gR3VDuQNRoX1cCjs11yXwyecaJVLXm5OViqyKRWz+htVrSQDUN
l7EF7KcmZMEaO5qxAnQcB+qkm/elqNIXzjmoHBvtZ8cS5WTyLV9X+rq/UlC3xib9AqcC/kH4H6Sr
Cr855G4QdVWliPyZtaUQ5uQwYyYYcK3yePnxgxsJajB/FvrXsIsGueN0SwDddjMoOmT+l+1xYM1l
9itjlfy6Cs4DlBmJRyijtVi2n2dEgFtS7RjqZJPYG7GSqiv3kHupmGU4vo2qqTpBRYWOSmbVTb1E
KPVf3hx+OWeF9BLP1UBLKKStxE+YAJwJuPKSnTU4Cv47p6DtEUyDmjtXO5upZrXLakFKpd/jUsX+
Pbq+Pv+yo+C5NYSBUlspysqhRzBQYiU5AAH6hpJ+c5gZHlbW2KJIg11CPlKZEN6EJzxvbmzW5kXM
YShI6SZaVrxzGN1EzgWN8xswqCZSeMZzvAGKsONJAcFCxd+wa+Xv2VImKfK/XQrxX/GJ1Uiki9n2
Ahvetnf/x25Mgjk7MafxGjq/MCAYj6BrUbwSPbS7d2KiueffVLTNbXNwZ9vUMSUVP4icHX7Eu7+e
zAxp5/rnrdQC/dW+BJ3bWofEmB5YvNFbBJMG5EK5eLLOaC2ysN07FSzbu/5yERWMI9LuOdnrMBmU
2jW66bCYxzMN/ryi52NkLKrLqaleFoa4zw8ji8yygb9Ldub0NgFgG+IE8qKgP1Td6Muj7MxMrTeP
l7fYrNUgTcMUlzks5JXV/X62bwfUPUJFqXHY/C+w2djcZBvPhRqjTyUaEcRO7N49RQbFUb1UX9Ml
ef3qZhZErpGm5X+cx2jgLnKV289mm59TNnFX18GCRB9RaYaAZoerM0ljwKHq2x6vO16RcEsBG9+m
PUWaBwZU1k3Vy8YUorXn19uvAqTKIjCqUyncO3AYQGkEb3Hzh22uKdMqHefVZy21FkgvQV16Dkan
JOe8OjXpEF+pk2GCeIu773b2CCUa8532iVsgoOXFoaiEp19Xcq/lTKTRoDkB40Rwaeyb8zfO0XOV
SXbG3pI9LtpUl3GG7wrxuACmBhsO65oMjs/DloUgaXCxam7jar+fmc6Pwv5ieK6GRnDPRWtpsRIV
ueElTATzuMRDUyabqlQehiBEKYUnjv/IAcqVaiXpC7tuGqcc/cJvyG6KEd6fhIGZL36CEuuhXLxa
Cf58MnM8Ue7IRcI8Jrn1FeWDCoKqglZf0+uqXrWlq817LLJqMxbByPw/QfJBWgt8SZOwP64Zj/EW
yd7NhshPXqc61w1ZbipTInG+KDPWLUS1Wqmj6opCtYXSRqbJuI9rq7ebzxw+fJTrwSd2iUMmJTAi
8UKeSj+2xH6gAjGkKV+DE3jIR36ayHsuP6FBNwDa81/ysdayu966Fey84wXhjDZyVvyYUmjSNbyF
naLNDhjn17pJ+yh9ZaTEj1GIABpki2wZpMXslA9xuqA/1T7+DfMvcPtryVtHbHk1zGFseAZdWlS3
l7NhXPpNxV2nAWJXtz41XV9CvatfHYhP3mA8oz0QkCPvh8Dxh4TbYUzqC6JPaGWsj7++4ibzzQyX
1yhXOCBcU/B4KVXwVQ9bXb5V2X/dnxBUL0AI0AZIN5x289xdeWQVOHT4NXCrVS2aihobz38wQ64B
UCw9cl4n0PIVQb3aamNxn1/mN3CsMdh5U4QLONB0QshJMx/5JFx4LnmlmdQeHXFEnAHaKFq710w4
mVJm0njQO3LMYwYCau264STtv03t+wpubdZZf5egxbPN41wO+rQMbyDNYi1IWTFa3MxbH/XCMeuV
VqgGMpfF0Rbul3Pm3983Wz2qP66Z52sCWIlCOgrE0EBYDmwUCNlDo2x4BwCQqaHZZTAM8yYWjnRP
X2/PxNRyY1R9PXSnS4m3M0rS5dmuNxUebl1kV/wF1YKtx/0+L37A41zXS1hSZ9s/EOzyQX+TwKfd
GATmvVeFn9rCVJL/kGE48zrAJYlS4WctOc9VTFColdYP5rA1v9v4TE929rwk94A7nZFsB0Hzkh+x
c7qhOC4kIVpGguOHdv+vTwg3bsQVTcg3xX4Ng3/vSyDgPgqf6+5n0967mzBWaFL3NIvZnsdDtZQa
FbshiO+ozCSJD9Qns6ewpmV2iIS/xJZ83spAz1yzBf2jnXr+jvBvQd8Vm1DflPPO5Leyct8XFYSb
JhmBSJ1nKteFqhPh2jMe/3Esf16PUqOWvfZolu8k3qJiJoWkrEXIpb578zwWTw7Wwswi1kbB42X/
bVHx9SrZPfYLztwQMSiS2AHFCwrFXzIPuubNKQSMiF5fnYTrA38kX92BMRxyuDvqWqVi4I7prbYA
cF/OjGWHFv71lx8IKCgwCnCw+M9L5aiEtYtLRR5rIm15dZwQZpr5zJweGhQUX8NtdRr1+hOYAmX3
Kuupb2wv3PUPFk6f/qUQQjXIopIOWcln6Yotl2igUx+9Php0131E4er7DR8E1h2FakJBb5KUIv6f
ST+C5Uu7Y9zyn3Z5QM9Tsz+w1voU18Pqzabw/A8AYEvVC/sIO31VwZsJ7bqDQNqCPa1l1Zs3l/Jh
noWvXlp+7IBzs1xps7T7CuoVIL4780f17z8JJdG2TTvL+0GAI3EGOSsddpPNxx6RwHE0Pb2zkgqN
EbS46iLPjTGrIS122MzTX/oLvfHCLpUzqhZOPIpaJ5xNaJLBNXD8EwjMG5SZ72n/vFwfJ5g54bpQ
kodqEyrImAIcKoF0us8qd1NKUQnFT5SNmY3KPtdsH4zW+5D9BD+W3x9Z0EQpYiMEQjknjuJ77CJf
faQxcbtqlmhcn1w0/RfG83Iev/4dIAUBBEiQb1RzT5S2ql3Ckxm10Thk2IvyvUzj4ODPamtM+C3I
aBhZ+SV5j8CcZclNF8MF4mpZkWVNTROwPfO5t2i+V2LugfFs+cUaGIF9g1WeHDgyzMqPm7N58OQq
ut9fW+/YZ38gpqzM8DMqovrROx3FMOqZoOKcogqOimWNqwxeqOkO7NCfmsjS75tEc9OEGU2LMCIz
nvMW3364XS8SfZ6tIji4zOSC4SE9mOvb0lqTqlULGGf2lqrhbaKQhszpYWhvYQThrCJRMHrjhP5+
d3k7vqNgg7Dl/1MtgMSFd+fru4ZstUbgZXoOjj/aupZ31F6vsphWQz6aBwxFz6RPsWrcosFk/zs0
bx/MPHPeanG8LYvpPPll/zVrM7qcckWg9QhmQNhCQmYFkfJ48EjPns7W913fcQdNwNsmGHDK2OcQ
gYXok82W8SXVriyYyGvtUT5V+rpMeYe44Aeyi73BMgtVjMqftpN5ClBfqnn8CYxDcSOm2q20wr6k
J6RZa7OWQcdqucCqaOuSKDof0K399z8n2wAPzXGm4TQBWdCVRccCxK6kyOPl7LobDg+H72Gnz6kU
62mFVz9uR9p0kwP960GW4hhhvlPt3ODZd9iDobUmGwBkatJ3InhhPKEzOsjg5FS71BKoa7g9zv0A
n/rnoxkFaFV+z87nxrYiFMJaUktBhyFragyEzmYJxJMOnZ8QnLcvnB6J4PoCV9zfC2Uwouhd10c9
Ot42MTtLQtTL7/UIlV0LIzfyyO3GsDDB8BGRSApF6kHfKk9Yvoqcd2/DnZwF/KqboRc34K+1kzRw
BCQedHlsXJphIRVvjFgZivbmSsuqvHySjQeWTKHW/3+Za3iDqanudY74CEx6dpEvQaAj9X/m51Ai
ezVH9J92l3M4QmgXS/k+bUc0CN/sXDrcylYm0/WLbaSc0+7KmcKUxwHrg1SvwtXOXG3mIpL0Xvqf
n4u372pwlotulkK92+h1ekpkvpkOfFShODDEfAQiqdJKlflY2frbNbRKJnnq05zzKK7N0m3UUirV
kPtZK2rnkm82+eOyZ1cT84xqmtd9qq6DSNTNV5JS6P47h10CWg4BS9/9F/N3XdwIdYWIxWsNM4F3
uh8DHl6OEkVJioLbcXc0jMVbegLMrkGld1PIXswW9MvkBTyGRpWdwcEmjesDfeW4TdueBiRxObqi
DVZgykQwmwHe/Y1hGwTswnsq8xyC1JUiiMCPI0WXXYEF0q76+HMbq6F8Kb2lzeBwcHgxaOo8zZEM
/ozN8OnXUjgyV4TbWIWuxSeipoA43cg5XokVijCK6VmcciV4qytxASt6uBz8icVZZ/MYvg5DnWlB
Kn1WLlL6hx0mHwnclctO2n5nVwV74X7Vq3pePzQMXGXWMtl+g1yP7ZVrFgTYazOdWm5m0W/6S13B
RjeSn5rd4fH0TQNBLRBC4Lo3wca0dE5D6reVpicAXBdqyeaui2iG8sU2JUWZN2JEpml87TsGNTnH
L9BFMniwRIlsclwIpAwHXypuCHcEG8Tb7GgKqJy2oVKuxitfMQgDf3hhihyoPBqTkrJTJOug8ClI
+nj3XN6cl9BFFekvVmxNIWgTwMCfDIjYPgR+fEbdAWl6EoFQop1Sa2gMEO0oYS4PmBjEOm1Rt0nV
zkl1qC48nnrUgctEkVSJQbLxcpE3Wzts2iFC67cIFm3k5X6smQx0GS9hOhEXBat94ZWCkdYuBvUA
PcMJKpPE07zVRhfhBp3Ra1Wd4udTxutXaeAHyEatlkKeCZDKx1h/01yAdo5iYeq7kC/BPow3cvTk
VvUyRxThd/Vu3iBVm5UCWyevLB6FXhZUovThyp0TCHsxcoIHnFVy6djICtt6yVbTGVBxy5KX6wJF
WfNTL6wPzhSxo+bh83vlC3yskDSPeH4W+w2ldiOLqVMYdtzviyEC+XKCuzHRo0xwoRJYGisLE8E/
nFwkvqnCxXrrHEU7lSXhJBJBx1JHuw1Jhn8dtDgYmjzrl1uwlfSAQhAnBFxMp/3Jt+lIJzQ8+tgI
cqlx80yaHbF5hCu5CFXnMhX4ja05T5yMWo5kfdGUweH4ryBHvk/TtS9K9zePA1rGUNHXuufLbKEl
q/M3ajgMKa1h1I2UvaydvurQpU2tOYSwXgstRJZ4ilRbKrvp9I/eagIwtjr+RkZJc7cfwjvizANq
Ph8tHQfl79LPkL302hnhEdb/3cNUI6lYG4gws1WZr+BZfLdfbbwFX6z9o6xWFAdoomSCOZz0v7Wg
p59v9fzdf9xM9uAsNpjrt6rrislQW8FNkH1qZVjbHjytUel9J1pmlontBO3VTda87vCygpVmxk1O
0Vx3XXRKm1gHiytzvu0DoWbHEzQyPlAKqfkqZBgf8gm2t96F1JfEptRtFo4s7C775qfeeBSw+OPN
c8h1/zBbzwor9Aui25loOC8d4jcMZnsFEwJGdkJyiT19puLSGptSk0fwuN5jZc4SX7woxmxhz1Ao
GF1ffM3v466hxdPWgrcVkqql581Bnqruw5+oOt/fwriUQfXE/XTTcSd7Zy7r8GawV4bFwuKgH22T
aYHQq4YlruQSio0fnxSZ0aVXlYlDdag8pg+11sYt9SnrS4ss4wNhNXMpmctizhnRrMlpk6awwoHA
YRsfZ+B017+J8wBSMjCoW0B0/kJG4a6RFM3OV2oOV/swfsq/9K1y4f0xxLVkqj7hCd4aIY6DPpZK
B0MomHGXLt2n0yiTSNmf7YlThxGPkFpXUV9nlGyeylGEUfrSDa3koMNc+MBBVaXVzk7POzxsLx70
DLigDRQFVE5Qf+9Q1qjGIgZDGpzjzuKBSIQUVRQWvehZOJjLIYBn2WX6YgTFxInv2fft+OVaelR+
jqranJEOvteu6oEvaqGDtAU7jFMqM9gdufPf53kV6T1IULz1kfxxw1MEiIWznMwbW/K/YECtvKIJ
t4SZ68wKJsY5sfEx1738PGH3nmFUiwysKNvJvi+K7ln7qcknkL/zZNNVqxfjXqkKPCilQXeaKlh/
a+D50+XT/IURGQQaBiaEy8M5yvZBxXs0dKcjuEbwH8FcGJFLL0FZAaE9PqXYPla4lAs1eR9kccaf
dPy7KzvXO4xZJlLytj2UsTEt4tGaTFTX6vw5xB29VpAP1x2C3HskU3yua0RA0ILffHQfrlYfki0i
8/axYqVKwBm4p/qn9xXNK344p9fNRHjMKu1lnAMK61Jy7CzfyznwQfJ9s0tBXgHwGatP4cB3Zyy2
/M8y6kuvsn1cbzqxI4jnWUCzeRqCaU8hGvZCgQlt1WJRDIzd5aGj8KY1Dwb4s9a6hbJdxWpt71uS
AedIUKOlsrsLGk3+kyVz4JHjPwpWm9HpwntD/G+T56IEfxaYRh9uttCVnfqIjDedxlUcbESgqy42
w8yuCL0L67gDlC6eCQBa6TkKUzUimySSrYtHB3/6s+Lv1Dzqetwmf1/ojP4hKMzkFh3GT4dLmFb0
/29diVmwnAB3p5LIkxnEwWYI4jtgDJFNRW/7Uus4LQGkWuuB8pWeRhhqB6Iotn5gfHqzwQs8MXZs
cifujCs0carRw+740S4qihxPG5yrGBiACDhlGU4zYKCL3B7ub16LbGJL+wNvMd61UKMxSFJmqtVz
4Ya4jeOsJ+ZCv7c+RTRZWS8dYQxP0W8Pi8Kl6dJ9pPiIJ0hsXsuRB5mM8Kp/H8aAzc7qgTkQv/Re
ilfTbqO3qqUkP5A479NHAn51n6xacW+nWwF9ipn+uPW7yzKMrRh5gRcLXuC5YXFAhl42VQGxvSJ6
1DoPYOLUgUdpkSmvL5YrkmJS14Rh/BqUXl3c4wlNJLkHtjlLctlzIZgiaWroXK5opUGCStAHxqHf
jCCUEi1GK5sZ5hfSIQX40y5bDTPL7NPeFZYLA5E/HS45rgXSGiFQjlmPg7hqmyRfXlf0YdP0mki8
ax/8XdVRpDre+o/uevHOCVxcY+zh1KAv9CiWi7Nk7kJGykxmWVZgH0P4CD/RiN3pQSIt92yJU6ib
x0sCv9dqHbXITvs5ceuOCIzVySpwhyE1NmHDn630Gb6Gd8f1lV5DkQNJJIRdWl+GwP3asLI+j6kt
/Q3Hpenepx4HPJj07QrauZ5jfdD+6l3vfurhicRT3POyAoyhJcAdse2tEjACMPiLcGlWyvpdZMMm
auAJ/hhtbYEirLlrO9IKr0NJfgmI/heA7WWybFvzZPUpBo9gXY4GuSU6bac/uodI/ab/4i+s8l84
2qJbIYsiXnPlkApYxSQ1ilU620OB7FzJr6IZ8lL0bF/W4YfSulVTnEzVCAc3fN34I9D6u5X56es3
LMceSTMfJ5rtrzk7KH3fkTTvyAktNDtg7q4rp11HFQAb4ChLNE1ZB0TEN3sqk7ESA0FnlolJy3A4
6FV3CtVtkqQ0VJsuF/uEgG8J+VccD42NCcgc+HmkFWllMADyNtRgRQaMyhkOMFLBUdMhZPC4LXhq
cBdHq23GVnvC4cCg2cHGyTI3S8pRBYhILvb06NNEEQAb03rViXOLBVT4eCjG3nyQUNPRrgsvD1qi
mtFKQiYftdi0mHgHQv6b44o7irtt+2YjOgeP08T+tert+CSo+Byxv3V4d/cE2Hor/KtQZp09y90N
DFeauQp4w1mF6e8ye94+m/BvqYkkITxIVBYYIjYy3noEisxQaSmiqqx06UjV8ec6N6mB8DjQX/Ge
nh+w/5Yt7LP1oSPn/WoQBP2bVm4H+C7kaSKJnRhbRB+TjNQnxhQy0KjkTQ1BMx0IGZL3ID4+VpXV
/LwWktEI3Dn5coe+kY4athZr0jlYVF6uVhXQWu/ROJRZWwWzfOQFoLgug4f44MkAVZ9sgJ4sYAGA
Z7OvzMScL0Tm0ao7Gdga+cTC459QlKBHIqXiRlZXG7A+oGqZDXhvra8fsS4c2t3J4ntQ/J5BBOoV
36prb8cjtZZ62XU9ibfKVjGEzOzBGf3ojuji6qM3qSTYGEK/wTtn9flRgj8LC2O07G1pIP6H+VtP
CQ8BsU9/6mlAvxCGeURk2UB+0YdfnPSpIMrvlrZYF2Rjn+gh6cTRCSYPtJO10dcR7MI3u9Oh+m/I
+fjVJoNOSm3j5OoOEbY0WtJJececgKK5lA1ORabexQ18+CDLsBT5SLYq9IKud+d9y7ssMaIyAK2r
NtP3kZwcKkuXeSBme1qUmaNcHBKbezm9Ondc8ix/HPvdi6qqMjcwmRzbl/FmPH/LmuXsSvE+fRjp
R4WebKr+nT8iX+W/pL9aVNLBiN9MI4m+r5+Nnv+JpK2bBA3H0zlEhHPSRhBK1/t4dJJIQDdinIlh
tjHY0Z5Ri7QrV1xOdjPjiVkJunh6yZRU56gxUz6ARKuuGyvrm01+tPWOYqAmUSDUXDGp87btC5OZ
Tt1mrtX6LJ2P4GAMJ4rnFTOhMaZ/fvEG81wYctOFwqQFrnPeyFkVUaoP7oJesY/kxaL5hX+YC2cN
mV1S3Onf27LsU8OUG0FKXJuJCjxWP+VUb6tM4DJwBo5cidyZFJEQOCRYMBxV7h9L2mqciLcdn2Wn
MdKJtbykpbspYGK8B8I10dv+t1Docak9y0Vcp9vyfBVu8Hs4dmheaDKBkEweyWKlR1MKTdskBsmh
f0Xuhyx0Jd2kXq0a5ge7aD4cwHy/NRArOU3DL0/IlCB6g4TS8aPZEZ7SlbEBi0c3X/LshJVnSyBq
2FwM6htditaAGreEb1JqVb/aaTuWJknDfm7wkal9f+BK9EeOr4jlIZABiKcZHqygs0n/6Rt7OXxc
XSi69zibcbGFacZYm3mqOHKNHeWX2qj/Etva3MaeVuGu5JJojdUFKOmFtVUoFN8h+xK8nWwwP9e4
5IDRbvlnBpVAsnJ5/8HAWVdVdmFcIi7Nl6XY1FKEVpNghqx3l78NXH0dVm6WXjPEyMuMDgwC5Pbg
RDEpX2yE9XGL0pH84SoCAEHGxHuSuW0sdBB4NKl9+S+PzbEY7gCxQui0Nsp/XVaQcEy03La6RUdL
ojERL+sUS2/pYG55uMLswBGJCamu3hD3SDwoPZ7QJKqw3a5gfGLG7J66VOPnU+yWfcG8G1Hb1ZRF
8uwN73tAQwOZPVAn98UYTsN6Ja8scBJqs+XKtLnbgxbTwBVgwwRuAfESMNoJUv5xXDhS37iDKT/i
Q7LX1vv0rKpRqiCryXIdHIBAFD1dTQEzDuNQmvifPum7xGAMOpDw0FLettX8kLmW/kChG9e4Ro04
H1l3G1stssfGV0PzKO1XEDwKWQK59AbU8SCVS1LwNczJnRLawYcUkpGzqDOylHU+CNH8fvtr9j5B
oWUKdC249kEDHIMW9ptAi9Fb8NZuj8wHeXHZjytXIujyuntIJDmxH4pkSd9LnjZc5Yy9j0GpzL2g
5ahSuPOYL5bIXjCHqaYDksPa4r+6jbviKZrWXLDfQTJRnM4ERnYk4+vYA8ROF7MDnaKldrv9RUIJ
j2pCQIyrhf65cQi4MFBXzYHLuPEBLLT6z1ADkkBpggk5+RXwHd5/69uQY1KCcSLby6gYqloqOJJb
hPL1N8/Dh0kSxjMMYxiGoBnMeVdtDHyMqqsiPYKA4uForRkP8vaKB9/9cfgtL6HLc9e9TwN7gASy
5v5iEIljkkGc1YaGEYSpJX3xG0xqu/KmEUXRVUlsRfKJrOjRYa9ZzlHRagnEYvGX40vwEr9D5X60
+CXIBMxbNwVE1OSR8QTF6prZg/RfT34rUWTokCY2WTgRs/cpu+Tib3UaootjGa73Oy0wsMbFZfL5
1Xi+6TPHV+JMQu+COaLSgwV2mrZFTnO+YeOvV/FhvNiq8r8S8ZWGOoZhqvJItxGPAZKQCdljsn1b
lsoQ15djr9t7hw2innQn2Ws7LOAglie3zhwRBHf1xxmsdFDxtY04Ms6dsM9edNMCGtKmppS1HFsH
HQ43h7XFRjTPoZB7xNS/QpO8aUAIJvsW1wAlvUd9AECWmwqkCuNGueLLVJgx/KrO3jwO4NOWa2Hq
M7qkiovi/XTy+0o51x5LZH9ixCLWxTBvy+DkVbyJSWhdKNpjHcI78OA+NZR2W1TWZq2LpU7uc16s
CqIYlRTkb4Nh
`protect end_protected
