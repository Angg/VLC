

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
gD7l84kB+WAh1ATog3H36h0/cMgn9QL5jGe9p9PjvP7N+FJAVvGVlrxcgBw6dZaWDNZqNANQuRFv
ZSE8fsSCFg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
YQUcxim/tlzHeVlJ7otHN7u41KO3Yg5DFb1yF4GCsbXGLtUvWNlkFjY+UPIlgYImR4Zo4dTHJQ+j
3BaUNSUOqAVzT9CfyUelv2YD2ZTfAtzIe1Mboyb3+StKnuzxnZmIhVPiZlowdW5lQ1r7BjDPOsge
ztxOfUTbvYcTUE1ABIE=


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
eu4MFD/NMz3pssr62VCh1XDd9mthYydX9VaOq3lWUwHi5/7e5dl2SAWHtYwTnBgGPY+jCcMycJhy
WSlkhQxVj5BsMm2aAItwXFvH2mSbjlPggtI0/+DNGQ4x8LQSFLTDYnnQbBrHlJymsS+/asMkXACD
SJ2tF8LF5tMhAlMPZZ0=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rNAzbNlIFUMjdhvgzZ2FokzvR4AuFtV+1AHGDKa9QgeBsZ1e0Fom48uKbJ9iakvqUoUcKKAvRzeY
OBkbx9P7Imx0gvIgzFsgiVw23cBYWOhbhSqVb7mef9aKx8yeF8T48n7gKldUkwBHIPeqaayRI9/Q
HCZO+k2+HCjRZE6L/Gzd+IOdEVUFOg3NtWFPk2JFkfZkxs8X7Vg/xxtvH7uvp+/EbVyiMbnwDT/p
NSqOyA+rJwBJYD3xRIPTFDI83XJLCF+1i4E8hyu7Y0F9MtjKugqEHwAG+JK3jde00nzNNaeLVUQ1
OfFMZJpkk0Cg66d2cvJY/G11oPkmvTq/JZ4+5g==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
apuTRT8aJu0TR7Ciy6ONiGK4AT7TUEiokS4gFf1g+kDg6PdKk9VRun4HKszIadRtahjPQo0of9uS
yvu3GS4EQo+Y+T116wnAIXnZSa8EQaEsDkziOI+rCvXv8IgaPYN8Cq0aRlASFL7IHOWNI49V0c0A
FIG/+5U7ZyNQFCVwuE4gCgK/pA6apm5kY4FGJft/EdZ5YAbR/nCTzK4P53+XsKHrtGfw+/MthFWz
tI0OtloKqc7laKZWKOVFqWq8Qmq7UL6utFODtxEQqzczH+q+Gw4rkUyOosIY+cbB67hX+GlmXXEF
jMwvUcen9t6c+wiH6rmBDcUIiuUHHz6q+jCwJQ==


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dfDj35aI8y6zqcW/IHFxmCDw2mpyex25qQAUnsL+tIRxivv/85PqpCOrf3b7NWnwUKMrsxtw+JBY
mtlPsVxQKR1gn6VkaHwbEgwxXXxFe71Z+1nWQhfF8Nt55jGvq1joWKMrurSV7Mo+HkvHMSszXj3v
8ElD0S6sN91oml0nObejOhxzHf0ybK+sGag+CFA7aBr4k4rYglf7AzOYrPl3nNoCkyrFDQFa46/w
SXJm/os7zUHbsDI5GGUH3BU+NktHZV6GK3iyhtHTwrMgDtpGk6vKHMKULM1Gjv9g1/jp9Ao4cUhr
bCVOXM1v2e8A3564rmh3if78zTzCKamPRAB5Ig==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 962560)
`protect data_block
716GM0+0QFfhRz763sNyjXBTQYUJ9ggB3XypPcp8NV6yKYgX67gSFLWxShcTA5+7w+lbku1Wkteu
QpDQoESUINhh9tNcRNIA0Yd24teuWiP9Q++ZBR0F4oOF4HLx/uEbnWAMjgryiKSa/L1+oxan4SXx
J4XqpHzH2sDSQOBtY6ZOkr5+B6b3v/WOF2behEuJ6Opi08qEaBXiubLcgX1mwUetczXmoMLsd4yn
C0hk0vmnQY4NNzmInbHIAT4kfzsdeFt69IM8p5bJPQJ4vka3gjVz2cunC7BgbwGvo/qZyL+sF45v
+nd+x4Wg9GOA/4NZz5EXgo7a1xTkGv0QqkmcsKeqQgaOukUazza81veLCZliNLKtTk4Wa1h1Iwwv
Fwxd6xPXz2mVfblIfmMbum9c43emtW4bmB1df+bbutyqUwLF4TQU8qmwmjibEj1KUvSPrrYkxi1h
HIzl1Jcn4wH3MSBPs8sXy5yF5g6NaNqJoCmdf9/DOgvqe42eSpn8kmR1jCA73U6/8RXa+rTQ19/x
0eeOnmOrwpEqc8+81UfTID9e1Nv2PTc20pQ+5L4cRp3SEzn3IV3XCpBylM63zgdC57CrZFtWwU9G
7KRIzZJs0JP9431YGNmmhB3vloytqy5MyyBgRhsJXrUt24xuGuWqJfDxES8intmvfzNemPLekg1W
XNHbOES6UV993l+zWGMg6A10H+bGOY82ZnWRqKy69lcvNHsin2DfbBv4j7omYIl7QOQgLYpEpwNi
423G4CXA96oKmp3NhlyhqV2FMoIHQVEPgmtLLemJnfw0IdV4LDWcnaY8YgiYtSNZrpVJ0tLs2Vfw
ctd+LGY4iZssv0tYa1Is/KBA6XAQ7nezZmjQiJbpHiDHrTpMpbPRuJo5HjGn0SErXO8h60ONwMlG
uERiU/ZwYfISxIefLmM8pM+WxEqYA5yDcxd/NmPAhNQg8I9eQU40JNxDE8iAILYQTZlw0jPT4okv
8UCgBgbRNO5C0PkENErKFKAg5B0dJVH2CNIsXcndKeP+CM0xL8MxEMPt0PjOO2AhYS2geHOEuB0o
5jwGx7Uf4VjvYiLnCPy1IRPd2Mix1/QViHthy2CQuwmvfMsDABpWL3MsFOBTKx0p10dHBoc59aOO
mkeyWg+TxrIOWz8g3eBbsYZu3Vw8qBVjeACMPwgeuXnIBkE8how9iCJctHIokpA1lM5HU4Jh8XHj
zgSFrGdCbD7AxJEu3dFrjJ1BlaD9NF+bZoFBimoEWq28Gd0iF6LQ0NkggYgBsTgwjzOF2AwelgVD
Xd4MOHeM8kFtfyfM15OaQrgLvNw4MqXYTfBU2IZS8lfbfzWxD82ZbIpoCjjKqnvN1X8oZR4k6gA8
Hx0t3fF7YmsNg8jSN+k4MK0qJr3ylkMUd/ZytXrkYyu/7oQfYr/wdNt3VMfZ6ogTkKSJ3fx34XLq
VQyQQMXj33FZuULOPwtE2iv+u1Jy4zbfHsKI/EKcNPiyQbIsVAVRSEZFj+h+0VZrVpiErzb7LBdD
CAPnf5ChG0QI9sBo7EFew19Pt0XuZkjvnmmzqGg70La/us8eYvSq7JTxPNPpxWSP9zoaXlDwPcAb
MLBljdpWx55OVC1xhjR5StLr6efLLz2KUE7tQ2uZn5zFa4+oUVuqxByCdsI2iw8C2aCA+agzSyCl
lsYBtlMVDcMCCbNB6GK3pgPJ9q0yBHnKWVUV/1f74NWrROpin7efM0KBge51NPGb1s9eWhnT5Trs
AqjVpArKVsE2n9nFSyRhoE/bqdbJHBFPXIc7tpJcDBomMwkgWRkYgB/w2t6h7+70rM/hWnjF9/h5
a5thCvG48Uut4HVSHKFaDWq7G8JswSJUQSIPRPKqdjWXLIgDWZXpTkyd1pH06npA7iHUr1Skx78L
Xw4QSb5CYzSqJ+utIXIGyETAP77rShtf70acHOD6Ai4uQXoubP85eHhWO3BrWJSkW7kexpPV+wJF
HJ/bgWuCXpiH+HmW183l6eTAOC1KbclZS9qRtbarcuWwMmRqhl2t81PFRajxqrm55USGhxPYfK+b
72VC0r6j4xJPBuUVL7RdWRH+7tkaa+f3Cn07nqZnXN1BuxRnGWFJtcqkXObD/LbAbj0BSSxWJ3OG
2MAXt8mPeuspZTdc7R9bh9v+ZExo5md5zjvJvfz1AYDrrM1lpMNI8qjRBU6vxDJJO2fA5dntjB5r
xMUZ5HbDTdxhQvNAukJwik/QyqJTZXfh/zoWv/jn+ookxrrjmoU1BAK3CHp/ViHfr4Vv8tcEQ2+A
KK4ve7yo3Bav8VDV/0OVMfzBSUemPOa1fa+LVlA4oB9kloPuXHbsf6lKmjBRg3XHrnJrNJ4eTYfY
3uvgVJOAmF3sSHSGvT+ZKx43d+iqqBSnjWsUySbzEzlbezqILMk6eY4XSmEWJhlo1EPtRUORQ27E
qd7AZhHrMRjM8edaZFg1KF1fuQBznNMNE5OtfXCohc9uFXOyBwSGTW/PLCYUlmh+8/kyvnVE6iN/
eYkLYXMstTY0XWzFa3neJpp+wuNdh8VSS9lMwaeasCMXvWZH2G3W28ouYBbcFEVHFMHcL7aSqswu
Tc0k5IepVZR+yxaLVk/yglyCXdzm863rjKKQBhiZQjmvlMcmmhsFa1HTc1aVsPifZMKjVc1H2Nwi
+Hh4mupGVQzgBdwkCvmLNkp8kjlx3Z1/sjCfkcmRCAB56VkmsSFIz4qGeh0q5iwGNPEvCwvEoQf3
0afOQrL0BsP6BIB7sPBl2QJFyx+DhvxzSFKK+XfQOjUDlmpXb4hUtUcXmOBTlfsTQvDxR6kpRGAr
64KwGSQ/xVLBePrIEL87VdKLq9/zHPWraoAS1gtvfiEOdkZCEqeNcQR6AzDliGyHUBqf8sibPDuQ
yYH+ZrFSK86trQhqYP7beS3XN9emrrj/BdomyoB2aaTLInB2B8daQGvES3GccK0pKgE6B5R2qdeD
5KdoqtU2BbCLqyI1zHMC5ZThz4qc4q5TJR2Sjyx3wI8BR4TSXq4Ic6IXnFozTolPENMn63xUNvwB
jjTMzAX1O30d/oQ73nH9ri/WpfDeZK+l9UTMpE7qiI1gewqBxfOVj844YevwgfiLnG+CovD9nByU
99zLcpLafGgC2Vuct5PD1ENcSefcafb/WFjnwO4k80WyvSNPQvTsO0AINMqmj2GPSJjUUAFmu0lc
1fLHQv+i0CQCGnmHp2vB0zop9zCr+zkvTvPmOr8cMXK4the5cKaQWIUG1CvhNVyT2wOUhD+N1h03
+P996D4Rx5DzEfmTAh88T7SZsqECD076f2tC1jt7dqo+AECTmq1x9tzL+3DyboCL5WORrFNlI0Xw
VmmOQ9dz+JonrLI8KYneUaejaurhPQUW92kijMD9HDnkWJlx2jqH3sdFd4sJ4mqO7LQY8AUuSiQW
1z6diWNuMvFbkwFaP/XIHFhRcDDBMH1FTiqdunakBOSMcSQkO32QUA+zNwUARbAdKEBGNdN5ci5+
iRSwE4lYf0AV1kUGquvduU3tOqYuGXBVFm081sKdtw8IIVPIg1vVpq9XSlYYcBUtD2YGQqlOsUKK
w7zXm5fqRABZtWxE5MEMmaB5Rbq87fTiq0qP/UCSi9rI7wShWZtbLHpXfPEU5vUaXt9tnPtaFKEY
Eo0Fj2o+TJMr5/UMAVMP80mYZQHuVdzXuQMnZg19nTUzbdjUVZmzckI85aqWrH9L5wpuHHJuFAIt
04bVy7sA0roslsDhaApbkAStjLJmRq0th8yGjpB9WF4+pMei+lljPX0PdVPmBrAawVfyPTfjrmVR
qe0sa2G1sCTR/I0mR/jguhk2O3RJCx8Kxd9Qm/NftjD+fkM9LENfmUblCE1rlRh2JEV8yAdZkPja
11KyoeVk1sgzgRnJ1g9s4/B5bFV8CrH6P3GY/MorXyeqqJDcujQvJfoLLRNiXhXO9/LHDnXai/Oq
14AB7//RU3JKfCfvQ3e0+QZgfoUGHo+tWo/bYCzbfSohonLQEonTKzWRE/gaG9nOwA4SPXDs3HMw
xT4RNhDWNei2fHCzR4z0DsY3F0OX5w9qfBlvR1z0qsPt7FMIz1YfpyIkBSG1vGGxCd7OmIQjLTtb
cJr7ddMwTrpWDKVWiRugC0SAXMc7adpnpWEW39Jdz27eN6jh9/Jw57awIzHtPE+Ls8Cioz4iI2Kh
SQ/kh6mKYIJ0OKK9RLBDhDlPvIH/pFCB0JsUqjxjqVewz+RD5EvgTJtnKRbZjGWla4JLfLJiRgNT
Zk/WGZgnYOIxeB6R+i4PnKs5Py8KV/fI6pSidBYRehUcd1gQrvixNRcau870E66it61b/+S3i9M1
ZTC3bvMdiKMPyf1IvukMXWyXogZVficcOJ6LzSf5tF+Cpzgj2uaubTcaOtZ1jz5zzyj2fDr6Y5bo
WbFOzkWFimPRX6S0RjXO8P5hK1lOe7amUEiiiGRfa8XU3/ZhtVP7vIa/RFzBU1Wl6Fgku2YOEO7f
4faXZeAFgWUjhYVUxBiM93jZou1Jwq+Bsiehm8p9ZoeG++Ixmmj4GtDJNwl/zCY/mCTlM8RGT+Qq
2Oi7TW0T4aqrZGB4u5tf97x1CeTf6dP6rAWwTyjcQXBY27lCilrCYkNYN18HnHAZOjYieBO91e7K
a9tAHZ9BDmSSMeSlpi+ttkqao1GRz8PtbQd8jR46CkJxDvUc1iKFSgJG20NaYyDqQvrDNx1yJ3Zv
Tj2gzRMRvQBy9yiPCwbug5Z5ATrBytoCMW+9xbE9zIPpr6Vlgm4p1j6L14OyfkvMIorTTkdbZkvl
eE37CpfJT/NeDp1EnoSSMeWkmy52HAStyUoEbbYbp3iWHiELEZTi71Wm/MS2MugYt42JrYA1Pigs
mhvD3Hcj1UY3HGTO5AC/uudD5z6KQM5YIcoPbV1DfFq2ZwXfcZQd6QP5k5dJBelMgeD0uQRSEtbW
F9VljVJsFMCWeUh65XcxGpO+S6lhIG5YQ+UEvaR1nWN+ae5gdfmLIiDktTCC15Y3BudStewEoGUE
MlWLnU860Z/27Ks2AIX4ev34u9u8ZoMJMLKAhKq9R3alzINo4mR8QRqF8mtIApYu7ugm4lDLA1iT
0e4a8S/aF6JtDo3LWtdW87ziNCZHMnghp4MrckBiax2ck6QEB3Cu9OQU42IyWyftTMJy9A62v0oN
C6muGryOciMpnSvlNSf/NP2pv69BIsg53tdsr7Yk0cM6frcXlLzecUNWncEWVPP9ly/HoOd3//VM
gxLVQtlta9rCs7h939ak3foEfEBphN0Sn5XrLRylf9AKmlDhq+ZaPJxAFUgdtz70zDtuVQSJLO3z
8nrXDlmp569kBQJiEt7vio28fq59+ukbzNg337LLrsph0lCL/0rRnpch5GEN4/+4I+YNv6yzt/gK
vX0j6Dnub2kmhY1/T9DK0D4euORXN/XOl1ubStlHPXZGbvNKH5OyUspj5aKC9Tf3fLY5Rsr7SmcB
B7KiKfydxLZeDVMjYPWseQQ5RtPhVOKjpHJpXjkQ269u7A03Ef2ED3Gx42XVCKpcUXp5ZdRDd/IU
IYXyRWmIoCJnAOe9P7Pb0Ci1LpN+nD+KzeO+zZirRYz0pG9zcNeNIRf/5a3iXqubtHUjfvp2lwnw
v9g66k1Ip8F+hdJIGhuTTyXpeCvCoaIqmlh78eVQDiBOxxEoUi9jJDBYriM3lHh32KUrAcGy5hKg
lrNhViQm9E0iu3nAufLaOqdJ1mwuMGAS6CaBYwW9dK8VrCyEZ9ljASfl6Tvtp3AKOzIuX3XV0TGk
yxvxi5Qt/maTxQ/mlRJD1fRh1TiKLsaZAIWiuPCo8vbJ3eqe/VZf20/ow2iX271NzzvGtw1QJf7g
DAhCzl/Js03ScpiLzZRJxfdclSylZjEwqJOPj1wzA9q9mmfCkh7T13/Ujhg/Hb7tQVJPqgP3a05t
xRnfhzEm6qe5XsAudB+RSfg71+MXzrZw63b8r1KnQ4hqZHOGtbzN623FBLKJsIfp24dsKTST4wrr
h0/Q+sKUTxwwo3sIC/gIMXOZOyJhwj5HpoZMGB/Yxys1eLcZQCe2/6W8rlL7olQkSKnB0Dfo/rwr
tTX4sljJIqwJtqS0jkk8yF7Lp/kpB9N3QxCk1ciBahQjak8Qf/ZzJSM2j9GNYumUMa/QOE2R+q6t
eaG6l6ABaFcccZ9LJbbIedHStw4xd/OtNbqj3kbZXUN+2l/eZtIqRF+mKEbYCI7jluecUhPDtgJE
wM7urlr2acsOCbAAq16YAuAVaf2h0HweFbR1bpqhiOFGl8smCOSn+Qg8J/wlMPEMqdlGxe/C6j2K
gl1qpCO3ZZO6gHZz3iJjRnPMbCyRxMePuAvCYew9oxMvm1bIVGXuhZH7cFlO9q+/ihV/VI67zHcS
SyphbEHgK7F+8RLsKFxZno/CJj6k/sysrnTBMXKQDndmOMtw2wepJBLkuT08WJbuf3MTHaaU16kT
weQVciEoFGBBt9756T/h/VNOE1MWL8KlH2vhQkZHT3HI1wgkdvJMqE6HDWCwT025qDyngf8Gjm28
6DIhWQX3+4JehpOaIxwj0hBPc2cA5bRDFnmk0gqpHPa5wYnqD90iU8YhI1QPD7hx0yOcoBuhDNMj
iofZq/BSOwexvUKlgADSu4RUwySdT9dCxhY7AfsEsayuTCi5x+6MLJqVYaITb/1Sk8uGXN1fgb/c
GmtHeiuDvrLTeN4h5qKMLYJq3Hn874H8e2QjhPA7b5JbjvRIbN+E98MZZJfAFxZO6k9Q5a+6owE8
gbfr+fj/qocDuATzjB6sLhukOzLgXh2ePQz8b65bpDH5mNh8x5WaO1+0AwXD2sae0iwSO0Yydno8
9yU7RLefoUvn9a90aBgHfTJM3DHQUbKfQ9/1/lVcuZv+QARiiF9MOl34Si34JG55/zf78icEEkAn
PFDEJHJs6CNVtw7jxOgl6OJCemKiZ4rwDfi3U8TvfMBqFpKgy4iYHO+/m8xFKtgK0CsB2eVdASsF
gyt2qlK6ZguEULdKO9q3rGRstg/PM+CfwpwV27IHW8pfs4xzHUBoaTMP34PnHCY7Z9RWcY1isWh4
gI0hkm+8JoUHkGib5P9+95xjOZOnirKoHAykT6oKINTldD+Vpsf1FCCT4jmvY7TwjezMkU3vQOc6
mEIqGP6TcJn5mdryU0DSvCgoZqIS1PhE2ulAFFHPnElCbffCQwi0ovtL1brt93wHCj7aYBp4AigP
dAs1tdlWyNIDG8IsiJ4rbS7eNmrHASFjRscPoG8+XI1fIzTNw96ANKTxBM1yDz+KRGGDZ9ZKG2fC
c3jhtO2a/cvh4/t5ogSPeU9iPIJTm1Fo6eJJIjDGmb2Jjv1psuerP60UJ7KZeJNtxuHlvQlO1F9Y
taxC5uv3NSrME0cUHTAVVEsM63xPHKzgu1NXRqVY9B2MVcoRSnzWLPuklonXhIliQ+ulKv07uVw0
EWJpRfDEL/OSPcVvAN7mdomG1H8Z2n6Y3JzJIMR40fP2NsZPXGkKLtP6QGo1d5uj7lZGBARnRCzC
Oo4FVrLUqvjQ+BPXWcCQb8U0kx69SNPoT3glyXnm3YSCj7UAAuDSeYRy2R+H1sAjcOTGUH+jk1dB
x0LbHC4JmpU7W/alBanSUZ2j5LNO0b9B9Km0o3qPo7NNf10TOEF6SQ1T+Lg9Uw3oSH9y8zxoumgI
VcPGKkqiF214aDj8ZaMK9yWQ/sToSqgVoUjUYCrH6G/TlkIwMRQyYnsKndKw/BkiueTEHkwh3hpx
DU/u8YppUhGy4bZ7ZkdJtd4Bs89IcmqFXfLPN2VU5G8l7U50RjjOMVl/lJDm7D+zyL6J7bZ0qtfU
NA5MtLod1vGLm8lOXW5oTFDgXQ9ahWG0F8J7q87wmuOA/FRZEzthtjMOLLsaZ1FDc3absTmJPxO1
Pw7yjJs2F4IlaYHJs7w+H/7ciHujyTEHHDOPYuwicMHvOheInIQS+ZHmj92r9Fi7lYy6fLLuwjXe
3XSALTTl/MfnWw1f3S4tQSpgBWRIZGkfqHLZKeilG07MToOECnFUaW7yISO4RCZ4GOLaDIuiQXu9
V/4nzmzcTmg+up8WqDmECGvwsIXJgEm6/1vZyKr4kFlUPE8/JSXfqFkpOjeaAw8s9C11DU0EtqKR
Y7o7iigjQszv5AB5vSBLZafXmD6NjUv/w42nLIjF8Srhqqb4a7uUEE1B0Pdt1SU70G8snRUyvjHc
r5Ceq+qIam6Pj9U74qG+xejTdtyHvYVlg3FF+MKuboiBxgb3GC2T4PdCPr7fJ+fJl3SKwzA4/yLM
K59ZMw8yombmKw9wT7W86Ebt78CVwBXOGTPWRy72ltv0metdG85LZwS1BIX8OlXj3ZJSCFke+nPi
rfRlfUhtB0akHOs1MLJpjFl1NJYbBBIp2yU24X3SlY1nmXFHVw0cWDFDFj4dzWccVuskXPv35y8h
vW/oLNHmGJCRExNJLIjnpLMe+b/VWO7g37DJcHYTtD0jaAEbJFxMUz6EQEFpSKBG7ZZUqJa54bkP
xE1l/1zsbfQ+5jbDJKsTotEh71D0FCTDHvhBzjaSOKMkmOtfcBghfBYolte6yVIbGZRiO7ToKE+K
MfOL0/YlxAIPzMkFtHRQAVzrqlaA4vzgz38bBeA38/PFo18CEzIupjsBjtQmdnaSv0XP3iwYZdXJ
zwTz7V+/aol71mFO+onWFj0R+Z5aP9A99AOvkw70+TZM/vleiRpP4VDS1ICOZ2U/V0ppi3QIQVFr
C6us187weAie24RHHfpnCijqFTq5Zswuxr0R/nPHY5xPNnRYdKXDNS4rVEsUgHM/IYDTJeqcb3m9
8GBkwZphyi1vnrMcWZSH3XK7yvQ3aaGM20YQR1SR84py+CTq/0AGb2vaM0IQzmDIV/uhLq72V6bp
nMla8my8qbXNfwubJI0Qx9tuIoauRBqGJeaNiI09L0eZ+zNi23jNRIjVsqEMlZUCeQI28oHP4MAO
XmgiQD3UvCxOpkCKfHWVVHyVLfzyxii/+8pNMg5L+zU68pj2G6xmBW6z7xe6k7Kr72CkFjMcgw0n
LFAFENkiobownkAYhx6tx+PaFLwR2Z8x9H1pkH5ugPbAsspIi0hEi6aN1cLT+1gTeu8xqF2oiFNv
5TboQWI76MyNfuhCuEiN/CLhxbaluSOYI+Nw7+txh5spB7O5emdX19f3xtMUWziOPfyF+7Rbxoza
nObDbyCAsFVb+I/gmON80ZuM+NFzkXhkq25Niuun5tpF454Ubeb+ullTrl+llyoywvmfah6BSAB/
antOOEpDzJ/J07qs6fP91slzFltvFxKE+SL3NQMqjWLitWq49qu0qBzcwGYRoMQRWx6dIuV4mUtA
ce9vjHDQhrGnm+ltw4fTgzWt0rvRbFfRL5YKqhgSNF3u6snpdBqs5ngla32AXIv4kBdJUaGLlTij
KG7M/oXvn6pXcl5j+pnB6n15sxcivna4Xb/rVXqtKn1QHaVut98vKQvTMS4pMh1UUHK6VwOsmVkU
TQyqcB8J0wP/JMXsHY/N/9j4cJJ7+/GD2YQry3kcAqEQnjjbmGKZ48o+rvJnO/TgifOS2U2G0edd
bju7yZJPiUZ3YNbLWQCJcjpml27rBTOt+mDn6C9o4RtOkXHg0zLLYEuy6uIAwOihxovluAMAcGo8
jI+L/id2tqjvIxpD8AMQu8bd5MRNgJfC1js7IL5jeTitUD78cogeNoTAPWq2ZN0dqewUON4Cxiuv
+mSgQkzZ+XmlG6OQ4W7IkByZPPNgUKRfTmGAGHzDS8qpQ2WL8KSLBlAU5rIC5vngMyckA9KsidZk
VhXsGm1Nqs2sLCu4pSQFhXJ5blFRQJC/KSE/iX4npRuKdBUY0zE7vw24FH63KxsjcCV4xnacAX3O
PjeF7kmEMLg5VY5xXojW8uLZaDyShElGd5TBVchSu4IaBWS0m3q6BoH2hcSFZKAxqKbvqU9snNoQ
HtgVmIYc672cwUXdctolBJzXwHqJjXFEPACwNAVuBTB+zl6YLP5eaCu6J672LBk8cqtrlSZ0Fa40
qhN3CPvLepKC5zj9UFxxLsQ/vd8KeZpPUirWu3/gWLI9pw382B5NLjvmtM0koKQHwucegIREKoBR
udW2nwfrgEKAa0yean0BI/RlBcD0eG/eq1MAZriT3XPVv3k6sAdX6qk23FFM0GxuOyibyDeYw9fE
CSlqp8DepOhWZWFyheP2SOFNULvwKK25v4E4X4pZS/EU2MYYP3cIAtZxT7crchAKSXdyjm9khWpm
0z6MGRoZiTpA4fxfIC4O1rw4krV07X/7tj+b0f5Umc5pSWphs7sz3ZyNVERvD/80BU26Zqo06i4q
T/bBvv1IQ1QbmTr5jpP/5BMheL8PkKTIkKD3p5iW6sXsXs2rpHngFkR12rxT4Z32GHVxHLJQoOVt
sj0LwyrofAga3eUIyyuYuMAw81MnljfQFP9skpmmHQDWFeSvd1oEIsRdn+My3YqQw+P6aDBm1kg6
6Ns+KWBAKPIWOcgzOWwO5EtREZ7Azz09J+fyr+g+ukF27eRVedVj2my/AL1ohVIXxriAQbFp4blS
Yr1YqN0tsl4xMNDzngJArdL7eMY6pSICJOlqQl8f68SsuoGJ6i5DIkHYFDA2QM/FxML1Km75jLGp
YEdfTJnwvcdq+ap/xarn1yOrMNrs37NUV6SQRCKel1J5UI1nXyk5yS2e8uT79ChH4IJuJhkhzSlK
kYjQF+3s8LPhcShM+TE8uvmlnwPlOhBKxp0LaYN3N1z9M/fJakvpUHbreGdOVA20TLy+hTH2DseR
93LvpR8OQzvzrwSd4lqnS114Fm6IR394pZ++f6kCacDNoTKWb3lyatbqYcXiFS1M4Ep+G+NpHPBS
6vdwc9UlPAsquJFsOAiByCL2bGpDhgZfYxY3lwDnBWSXQiFwgi1JpAf0SDiFQRqWIHwjxItF5qzE
A5ynCwqyuFSHZHrFTknA+s8qukm5hEk0VCcUbg13768xIlV/E8Dd4fhUw8StFvSyPooBMMASBEUc
w4fb0esHIhDHfVhx0u+1RlOG84dD3QpnPzBJDPbPGtaQ7GYsWJprYlg+te1WFrRwkUsbQt067+FC
oYCaTgY+BrdCHkU+LerJXMruAruYXhKHWyXBGv4WtI9vTAYcbW+xyM+9qfkkFOzeNAEKxfgNonrs
bg7U1X9H9DySKwlymDCLkusW7APO63LYGuWGMrBR5evmrhbB4kSfjEBRgQllDqatlmen6Gq82Mf/
jaTx0d2BnnlLnXLvqPh5cDC7pCIPCPwis6YZ2JxNKm3LoDjYfZVWneU1Cm51W7lAUxaCiPfKKQ2f
18VxMZyzyggHRZ7T1GoENbipP701y8qksSDNEaSnFnwTFG7nbb3agGbxTOTjAbwzLfzqeXL/bVEI
TH7dcfJjppqnHxZuUBia2EGdboU2p1YN/FN+U2gIh8UfkARk0Gf58jK14fwrBgzM2bALPVLaKEdb
uqUXfpG6wVN179U1lNKiOA7G6Bu+arHPkqykpWpk+LuJsxE88QYu3WhfXkzOUPJrmMnFbNGnOksP
B8j2po4o68KVi+/wG7JA/iD4bToxBVv/PLiRGBZgGJ1BFzRGwa03geh52nwdgg2mIm5QIbQ3nBG2
uvVq8LVU90tPEctf5rKgRa91p27V4HN2d1ThUzFRAikLaE0E6yGcw9wy8OYyVJ5tO4aE79JXLKOn
aWkdJCqw4gztZGUezQolAc/VbXRMPDjwTFIKLidR4djiSNtqQmdJRIXKrCv7iRM9izaD5nmkWiKn
IVsaaQQLZHiEj3fFZeWXR4f9YDU8RH+3j33rCk/RTajKdJLmW0W0M19C1tw+YhSTFZseFmCUakZr
wNcocHfkzz3SWF0VSoqDWANXqJYUgp9PNgWbHnsBFinWDKH2FPkzwZnVBDi+rxYj4c2v8qgZD+fc
lhUPs2b1/xJE8hOLUAGgUxvMbwDNoF1U+uXNJ0W/w1ot4Q1me4yWTbDM7VuILFPtOcoq5XlN6fCn
+1ODfaqyaFurGYNFMJ5E/2cgsnCKSSdA5j+Zf8o6/2t0sUk3MjwEjjbMpLGhCy/0VtZRTKrFERtu
qcE3Z64s13vAJ7wlNTmgT/yuURSIxbqHGCF6KjNJjPeH8ALIJIloQ/O/0XzE4687Q2n4lNtynheW
mh22ngihfMrbVt6hABYF7eeHFhznWAysrhGAW40ivis5meCC4mym5nSxHPH+LCb74OVYbEM80Knf
2sHzXdVi+Kw9cc9A7xoPBO8CgTUGtsgOn/7HCe+LC0TbuXaxJc/1TROKMeerhSCrqULK69pZfmsL
FLckOzl4FS7OI00CTg/TpzgHg5fG3oerkWmT7SLF5cGSPdDjwrQ1gCMiQC7nAW9p/X0hEwcPs+tf
ypPdZtzlJIRVEfXnryRwgs6zTpvD8NPkz+KN9mYMAGnRc2e9mfml69kkO9dGhoGq6WbAmflbK150
/HN0V8+X1bGLwyqVJNnMudNlZe0HBsX201HQrEHmoKKUNQzkcFtcLtBpHKSI+YNJRj+h6LZrmRKM
oCJDs1cx1Of1JIxu0y07/NNXofrPPj7NhkIaGK5/Ymg5bWsrIjBK8QWArBO6JneZ2uZ9OKOUx/BM
/6A1XPQhaB1a8phnRl/SpENPLGc5Vlm6zW5j+xVrVQV8AJGz/fVum/EtvJjycvEoBjVXBY23LdpS
XGY1gwBH0EETMfWjILk98lSfX7cs+YmJ3QTG7KZ8rEZbd8Ojin4w0s8PxaTZg6fuUca65CmVIWbu
i8/tTAFUSooeRtO+1SccwOofU0pVXF9KPo9XhWAKFetX60UB+6JXisFvBAXL8bBBdlWJEzemBHls
ZDuhOKL2+eEoJ0PEfSMX7lyppAre5S0taZTTXYJKMi71MUeL4VhE6/gGhaNHpgYBhyNzB0geGseg
Ww98+LjF9dSttZcN1YIVGok3Y4/2V4zaTAdCl8tk7mC+MIR+KfN0kmW1YDfPDWGTcj57XsxO0BTT
7suZ0bOfvXxAnKSUQn9ts3P4u2XaHqCTS2lyg2LZ93eqXhEtYgo96GwYr9ADHFHgE+Cn5xCiPZIi
D/M/gnm9QNVnpTUpoWxHMyBaDfxECHxCmiiM2QR82mTOB+rNoxVwLklc5oldv8VDcmkH8ryJWAKY
yBYvlh8lOmMxRzlmACFQuJEe5+Vrl56XzYTHtZUld1zlEm0Pj5xSrqPLBnUuJAlnHWJGGoZdge2P
X4dJtXwgnpbTB4hJLVIlvFuCQXBNjV5heAxZ8LqTl+4PCXbRJNgBfIB1E5AmLMAR24u1/gcCg7dK
/lCAdNG4XkNC5lGipvkpHk4dR9SzAUJeFcqHSs3LPMsyrBKghdwKmuPkjDyZZ31AcvoAGh0fThmz
m1UN0c/R6yVs5BX2DR4UOrCnybC9ubneYXWs8yLzukbtpjmPKt3Jpzj7CcaYASWeLEQ6sqLoZLim
+bXqMrV+AsPr87SlJbGlUVa8ZPdadsnkNzsiElN4faRquV9DIFYP/qfNIW9xHGD0wR8QoQSMZWfk
Xh+7gNz2b6T6op8JnLaUQYUZNqNbHp/EzNmzd6qfXQ/aO7QG9uPsJ9VdlV1/t41BQe44hxpdKLHW
AKj/ixg6qN6p2R76FEfXE83/cXigB3UXEOlXXS34ZHUvQgltRXgbVvHyn0zKx7RRhVGK59+uLb9B
XoJcIgbGfpPswaTTCyZ6fwlJeiE/p3ahXnTNNChzl2yAGZHmigR5B76LmcadlHKdvHuF5Y90vfW2
jJG/Fh6Eb1wMwQ85QkejFA9UwvMqkHSgV2v9MdLbf+/8G5HvofCbjUmlUydGhQZtYw7oD+euTnKB
sdFCdZP5MKb1B6TZ71Tw8JhnX8g16nRWE5nvVM/hLf3gUOTDxmQm6QEhZPUtbF7+dX1G6oUwOo69
DilDUZNkX4WP0iLb9le8fn1aPtX34HB0keXTSJifNm+QqeXoy+ijPJv/JhN/uSvxGNsOrEgnkiqR
H1VuHsxCYTxmkJDY3/JkisA0MkXJcYfHbIXr4H4OWLpTqIQrsdeEZt9hAdFpyrVn6pbIWLIfSLjK
UmGZyLkvV0YO0ulKZcRW4eaxF035nyuP8uRLz5zfxoMMFEo63tGqYq8wEY5rXgersn3pqEiuOPB1
h80Obyq8mhoSC+JAwQsB7owYbvdGwxkX2qZyNT3wTzWqcqEzoqqVfh38PbXkvTKeF+zAX6eXcbxP
3uL3pfHv8mK+m6fiZkwcaZewGy5f+UI682Zb7hNryDqUHJgBZJ6+2W2wN7w3+2YttBxPfr52RdaU
wQ/C9oFOrQeEakB7tCCCtD/ni0sop8+IzCrvHpSHXd906gWydpG5x9ge/n+wZlaDMGhJfpOkdYgW
rOOYRK3bjifTZn4JSj+qyN7ljwmo7OjR7Nahr+9SKS5Ltx6oxtpz73ankM2rLl8kOW0AJluekTny
mBkihG+3IPi/aBHXce6XeG+sZdOA45tkHBagn6W7sM0DOIOEI7GF7uo8cGw2hQjgyAAp04nmEu+3
YKnmxuzfBTg7JpMnTgc5TG0qhrc3aiPwki8GR8QbifwzhaVveQvuj06uwfwp4C/BrQnpBY3Lmcd8
hAY8Mn0IWGQoAXQJKZv2il7wFlEjthoqABwyzXYAidbTHlaegkAEzOV4t6SaYNYKOriTjuvWGBx7
Ci/LRNwXMlqW0UCCKqBISOFZf7jBE3ArYU7oHZanAkdlZYqgQKAiKGPlyEFLrbCIJcnOFHLtg1aB
JNgRMXZYEm1rOW0SnRYA6OmYP0iTyjsTy0Bbd3i3mIBPP9AVtl/TA74YHtdu9sqsymi92eir3TYw
nIC7vR1u7ukU991Wx6x/mJEEVL4ejuR3Xi7yONmw3U6buerUdYM82Rgs8xD1doRfhz+WYmChQEnC
mTfKNY/QSjBRa7ZzCewxLPosH/J4IsiMnivtHMIApsDwGyC/7BBJYHQrLu5PbABp2v5Uovu+9HGB
wOHUVpsZhhRKGcf0A3Wn4LsLZJr1R2Ertfw+jePhHLMIMUNZzcqOif79ED4OVPOXSkK2ncAWAgsT
8ZQJm1x4P5p2Kb+UVnRvv7dDDxnLRXD3Uor0ErGgkKs+cx8yFwYbMR/qH6HOAlPQYaEL9IElPUh6
epsfZTequGlDXKRHiUNYTgi1ksAI295oZSlxKs0YrrkG5gGMQItIySgiJpuobio+lC91JPbAQLFS
Sbo16SIQKryj8HtPeCAxeCwD4OcBnNKdu0ub4A/BRiu25Q+ieJDsj30zTcya4rJvjqO8UVktfFdV
4niVREVpiCyKd7EKEwy8w+r8vNqCcZULXZ26c2N7Xl+MnIODRmygDuLCgHgdWSW9vvlrQdmPevxi
zLxCmwUhwH/K/W4JfphiEIkrT0pJbBE2aGaWYDuXQyp10FmK7uD3htJKpr9QduU4AbtWk6VCsZFJ
lbyEd8bGnsHWl8AJn22jxogoXIOVkxvNFdU1a5I1NcCkJ7RqzFpDYI8h4hdUh630qzFBJuZQZwDr
naCtMTtbriTqRrX0eWT/tPBQlkoKXBdPG0kL6H9hM9ToSSUh3GTHYjVYKloZfjEkR2ggI0b4yS7f
yvEZXceClfsJ14XXaFuDbvEH0T4tXBERfp5HxekbN1e2N6MKKXwvLhzt6zZbk1OjKNfVNR/fdtVg
FKaaSq5ZBdtt3/5Myv0UCSoRMvxQ7EPlcUbITTqKkKnedVgNGqhOCj1jxSZxBp5SKGmB0ZtJYGDv
4leFo9K8s1UYdK0q2OpolO/sWsfsWisUfWbeSWQMYK7j+51yX9y0MZT/q0mpKMXx5q5F/a1z7uY9
0UmApiauuKugAkSvn/G/SRIteSSpz8max/ncsFNFk7jRywpbrODO0lJLg08GeKctERagfXi+cmqQ
YUTNcHTPeMhKrh7DDuVo9i3yPvFNSCDuYewrN73WAp6pJChLESQNmVqYlvB3/wjNVw+fzBogGujF
2xpY+C88TuOBTjGGc4Y7zyOaXnSPfzOu2KoiEsGfZLY+/bbBoDqOGUAZdvgxNcuErKPdpr4nivzl
xR/GR/GTCdx7zBM2sBdyb3Wb4d+8+Wk2sdNB+W03x68++YXjqAxJ8UilJ1c+ouuLEilWDWZgPt5N
5nFVV7D8Hfgc5aOfLLLHfa0iwu86wml34iD/hOlPi6N0nw1ylSW/s8JsyBAPuvTe4z6QIzzu0plx
4IJmXZhE6nU1O+VWVzzFT/wSkKgoTzDzW5S1t7lXKGuD7TiSsdm8/olUOd9cC4BeN2om7DRQZKLO
NmWcOiy9iydhNT7JnSIAxGF+Sn+EOrQQZi1VrQBGxgy+iv8gUXelsRcHzl5cnQnMI3+HSWom9EzZ
kP7GDP3Uhkk0zdx6DeqAJ9lO8kUCTF4p4esJVe3Gcl3LtE5Kn2SdwZvwDn0fEBRYmvxG7Kj+muWv
fAqVd1q/ynZ8YgcIyzWJrV3h2qXA+lR9hIw+6sgVTWi59JD/jwXmmG9HfcQLT8zMS5P1swXXWVsb
y4YC5zbO6u+k7ekyzzxkRbjJlkh1/9x7cmsNqEt62gezOIVddWTofwjKiP3igXBKUqqjqi+QAIqW
FDGbbGG9IO5wNxCnHya1/l4C2P1UmHLyAzawdiPtgGDfjhZsc6FgoQduuScp1B3g9Zwmo5hJz2Gu
xyUIhij9xwlGnmFuF8epMTZdnb17J7UQvD4P50jtDOq3vSrpn46HjJMTs91p09i9iaiUpLvyK0vh
+SEgqRR3VEZDTEXHq0Ohsppx70iRxrPZ2XhpOat6grhO4YmGDq1H1AQn2V8uC+eablef9nZMEmwu
OVuUueBmcqEhdxyz8fFerkCP3/id1oBt7Fr6rFHO2VEhVqpjx5CT63h8ZEPN2WeRfP5/HW6QFFpj
kIdOWhCiAaTzWL/qOKTA0rDf2w9Cdz0qUWeuku2OpLEVPwBlBYzwkyytQpoJUWKJ5i605FIKNJke
rS7BZsIBEkhjQvE0WgMXHmlg6NoNmThsj2Xx69JrYmkMOMqHq6Dn5m3v4IUV3BHCvx7LcPqlgnzU
Tls+A+DGuBwo6/Z6A5H3xDsMySdTYKaBPimptgOv4P2v+HElDOAscO9kbPo4/NhmMsSoUUUky78q
pNSFc0/GJvS0ppdcqVgP7VCtKwN45D53pu/6euI7vWic58b+T6gsxrAD45xAeNW5/ZEJ6V4t3N8P
avbKZ1DeqpbLtk0PxCOnWCGDV4EvYJdGRSsWB/Pl1jRz0Gb1mClWJLlT/xYDG1XZmf7uRK/O8MwF
b8fkEG4PJN+GZI9Gv0h9NrsLCkFfQZBA/kd43WHDWa4hAnieuzJSFDytXDwsMH7kf/23WBvU0ut2
VCrj4h37+gWIp3owzesJ358W9IJRdQx5Q1jHI35I26EXxWZgL7lj61VDdsqvx265zebdn6rfc/GS
rIg7sa0JVAg4cFtuSYkAHDQPm7IlA1ruXhtztRzEp/GgVHgCmwyl3q4Fo9rw1DiEOrzz7rLqo0cd
PetS14jbFW/CHC5FSqcLA9htVEMnk39rOjBcE2a0L1AfuBHPqD+BsuppRDCtMA4hf+v3yyfHxemC
ld82hzuxKE78S5ReLhtmlgqFMVU6NkDmfcj+8+P/Oon/atPUXSqR2hOemAFcZ49hQ2DYEn1aNum0
xyFqRrRrtlzvJieeHs/X8QZvE9LRQI3pTtYTYotscmscoIgnW1akL8neGM7aqBbimYHg+1r42Qu6
YA1Y8u6X7qJLl0Cn/UATOo20aprN0X21e/rbBsFQ2fMiml4WHtuwHwsLBNk9aYieSJsEGicbqEb4
sJqsV24soQs97yAKHltFuenX4unK3bQWR8SMzPko5Ob/OZYuHqdcZNcwED5Idid4wgYb3NJtifrH
Ec6f8D4IuRrkvQtkuwJXuxdn9nYis+nuzzbHqdWjtPM1RUl8ibTmzXlqvDTRE7F9m6W0GrL49pKG
hDYxOhrUm+gdOb3WhAiGvSrIhYS51yg8gyHto4bQvkRKobAPHB+FyQwmEzo6WNRvh8tvC/CBt5so
8KJNN9hdmt29eNOiXzGqwPlWmH7wNbA8nGxV0ghuOqZpMTi7HNsFVBkcAPJqhsXQVavVjbL9pdvY
5w4GQkHYiNtPkyGelHwIFTJw6om/hg9HSp3VVEt1KkPjl9yG24A266KQXD3aHi46sMFItFYZcuHg
gaSrdBrXjuek0cWC4T6kmqXk3aWUOEgiofSh9pRL+/EVioveDBZs/lUZTK17clngGHYUKIAOr2Z4
ZMO6+Wc0CDXeODppnvZzcXieeDye6F5h/9Ksh7Lk91GpkIc7G6DIG04Zn6Gfqm6PyXlqy+USim3M
OfHIHngl4XREuZYyiGbCSRfl39Ef+oTl7txxHldPnv+avv531bLWgHw11m3Krwo2dj1Ruat9HbnB
YsW5ABJpuZz29YRISLIAh/ynkZ6M8JZP7jzSgidZ6i417F+uv5h05syy0YuOaESLh7puS+tHe2Qe
tpEksKOHUsZkTBExi8BTOmEWeQ62AsxhsQ9Z1xscwCx73Qo8wZ96C1gFv6L08hX9RTKCTa03dufw
jH9Hd9AZ33epHyJetygqpfrM6NdBbUrvyYtPrAfEPsca5dkabryAJPmVZGmbp2lxtCc4FKYsW+Wq
Z4X+6WkPtoxgJLE3ZEuKjStzXtHDkNsrzWsFcSvPnGAiZYRCo4HMgS7MHvkEMuPwkKjL4kyOfLMA
M0pAtDDzWk4XqvoVgf18BO1p8aQ039DzosgcLRmFPKVicB2ypI9BSEEDwjFEgrhMyTvfDIeMQM/P
kzFpx+tmn9Vb79NhN+ujJkapCNTMwRFPu36ZxLyScOwfuB8v6ay94uHNmJuhwRoyEkOujJf8LVZS
bGIn6+rOvthVVXcJC+aU8bjJQmk0U3T0WZZtvfc+q5pt2BSRAFpnJvutO2gIeA1+YWQ3ax/bE1fK
09UdgHRWgdlTMnJcLnU4g3gc+vZWKhy2bnh+ho9XmCtUyzVmuYbV3nFljP8VSdaiIsMzrm9fDSqJ
bfpvUNzBEYWkjOFNhj/h7Fo8x/Vyr5T+oF8xD1ZB2xEYP4DmzlxGMPQxnbi3uukLDESh19dGSwW1
GJEJhMP+ooYUmnH2n9aV+I2Hpf8RO2SvAGizMbNhgXqyLwG0bWNv4m30IPOsa4RS3PbRBWia9BRQ
YHYEMbeiHU5c3G/+VfqmTiCdEersesNoBGBY0wXqhHArk4KH4LZ8iqHcj9j4RmrDH7b9L49xhZ1f
TRWhFduU3z5lMHrQ9mnFY8nOAcJYznAnuyLQjMBzJxYzUMrGFipDmCayiq5uwAt/KhwE4nnHdmem
s12H9m6Yjj7LzPyjpVZmCpOrXD6wIgCBlFU5J7FYzX+eJ3krlhoP8OW5nsafitE00nT2+UqEkKBB
ucUkRWt7xJbX/1BoizdrOVA+N27vrE5e65uJ3RxrCRL08VYj/hHNhLTCgLr2oYkJ3hB/TbyaLyEh
1g5uoSxQiau9Ps75IX+yCcAYQyzHzPWVXVjmCF0lqJRC8RE+sAHcX29t+i4DP4cxAMJWQWewX2Sq
1LVFqcMmMfk063CwPaPovpzyASK8YL80Kdl7HiTp2XupfBWQAwwu9yjcZ5GYUFQNuYkwm7O0469F
b8RDzRlaFGAOsslTCQWPu0BumHhTpYwu3avPMVi/OPIqDHhRZcFw7toWZWW+Q3gvAAXEeN0nPIfw
u4y8La+iwFQoc9FQHbW5A5eJzYY4dZzBTcn5ckM4yTW6fP3b0JyeFeP7l/hdOpaggpjj9eko6pHI
k0ORAS+lrBgBoUtKP1WJJdgD7/cUpQ1DVi9Iyi3T1cboLOWpv9bSjOJk5i4UwdtH06Gv58Z+X+IY
BEEBjQ6zPEzdrpb779RmYOy24hflEezRziQZe2HI3PdvHmzrq/H6zQ+5PnpJGgETEqmkghNdOyq1
j1+Qy9BSnjAIcMOWK6B+Yf4cJb5vJ1ylxDTcdRAkmInWepcp3GE/9m25jJV1sJ7UsLRHB/5F8L2k
Tzw5QxnrvLaeLHqfl225Otc1MY3ICbUEtPV6r18mr5ThbU1j+g2HpD4ggLiNZdvefxbsEjGrpeqR
XYWEm1jiSkA1H7i3smZ/LpgEdqRVDCKFkx7j5NKWrFLc8D2otBwSRJ4mnh93A8191nMV5vgVwtSE
tv1MZEVh2xQNVh9o+55hGYVmrIldsnlny18Y30UMtLiuB8hUsgPclAFA15OD3cvHMknKhwk/z7bE
V1te3Ie9CKi4/Jx/s80aB3m/wJvLHJ7Wun6noZ4njGt/SsDo5oR2UFW2V62+vO0Gb6Bo601jtbqu
gz8phAnRkuqYxTTn9gd5DPhg5TQ2Kjvx+R0WwL/rXJ6gApdRi6IE94+zoIWbyAKJg7B0ZyOzPi1h
dMR2FHw7LHBze+3/QskrZjRZDXcpXlo4dDuJijskC6F/sVLhRMzxF4ZZgHqUxbk1sIr1mP/y7e6U
auxPqTN7glF+B1RkTdKyh8LR5sNBAbu5+ksyizQYQFHlMEcG6pW61+y0J+wEp9qi7SQbQBrOUYqJ
3RSGsdJcqW7/N20nFoMNfXC8rN2wFRO81AJq7857qCoNjwiBMxtkEchGfE5jHbWcquiT2QU4+781
4dabP/B7pYZtO17rraxGeKoDRUuGWw9+fLUwSoxgkjpWYkISmVY2VAoyqiIHRPVTTPcdXmvy9cFm
dntfE0bSHYW0zvRUhhfVJ9G1wDcobBY3shbPdveIFp/gITnHF2VualKngduIKp5lsjUxJOq+jHOe
5U+i9u3aqWYMo6hyr5y6z9d8Q38KDQ3Wfald6Dwsjfg2v3mITRbPiYNi9X26PdOA3F/fq8R6qVJ7
+itu6KANqlqgceahkjcsVXj76zI5uZX9rJ2x3N55nG/zKRwuw28ZD/y22lASLJMKejyRDgn+Ud1b
rKhH/uuyMCAXx7sYvc9vZxDmnYhFBLTqr+shME7UbRjxtjnQyykAuc9FoKD1glEefSHwIwv+SECE
xeVJl+wf7XLs+kzP57Ui3Q5xy61WIT3Iu8O5byVRy24yd2GnjkDTPLJKicDa1h0OMNJcpdT9yzv6
FsKxLyGkXwJGO6hdhCRbFqAoGsDLRBOFO6gmikFBH2YFg2VljwlvUouJ/W8dkd9q3VFg/rd9USQ9
5NGgR8iOxdbBJJJmaozdUc8vdEuknyG+zU0Y10lyqk/0T7PKkVLG5+Lr/8fZz2Hx5Szb/zbz3Arw
rkF9L6tQ/Eb5gR1UbwQrAmgD4xzcx/GvcRt8WtRbMLp91wDSPsNoqNvZjcpBJ8SN0xvZTF/HvCDB
m163bQ3GJ90vnT7dqMa8SyHUy1v4zjVKMAdjBgTZen0xXnSqHoT6Vq5Wx47mKyTTZUMuu2GsOyR/
4N03wQKBxTuNFNIXGyoYtXJSlOgsUamXXPQYiFM1431/vDY7OiGX7tR90Id7Ssmkz2OJCT6eLBUm
L3ET63GDktzBHHIhxpO+M/vWk87og/xrweZ10SyRf4Gxumh6hWphlca1VAfxr6mCUQBq2U2RS2UZ
ETRxH9AXY4aq+xZQvFYuydMxlWQQy9B0lfAFeVtYGspB0yDUh+Wx2gSHt1d2RupQ+NuKwLv/g0zB
uMaBhy7XbuJYDY4fDiQufR5Hn2th3Q2g6Y2vOW3hdbaI+SaWf8DNwW7Xo/p42DOtIf0MMMhO0XZF
gLOzUcw0sf2AA1Ar2ok35MAAlBokIOc0w0rxeh0hYGl8DlvpXjEZSHcPRAaIsT94GCLwg7akPa/n
y2zWhXWFpMnHU6/M77TlRS1TYkCmpQ2Y7rYLYum+7RdxBUCKED615KBpo7QAqBlGsNymplmLHGtX
VdARLi9z8aePqpULO8PfhZhq+Wt4/J/GZXvDkjOIcNt3dGk0Zp2miljPgKbApNxRXgHou7J/OQCV
kq7L52uHm0wjWDaMPTOp6l9+9h240kGiK6UY2/2iizdeZPyzT3YHWlgvHTvPwMUMvO6t/X+QqM0y
y7E3lUEe88L9URV/9AjnNY5Ao/U0kh88pstbeXWxhn/6z8gSlbYprn8ssQkoElkkCD7cVyYDHaJb
EbEsiLp5kc95mvXVNbYN5/l3xdp0A6vG7yx728l5M8HnmwUHoJuM0PLQdbcxyuxXPZFIr08jgCoG
Q3/br8xLPJY/FchPZwIXWfg0k29XG5DhNWXS7bjxL31tNCN9wqkkzs1ymtzOR1Qz2sIx+BoJS081
pSsDKHmtomTQ7iMDSlbYf4tDKBIvtRVJNIEbjDX5RLY3VO+dbkrgXkXBwhv+09a8ZQjORmraPPmf
X4omu/gIhznThiLoP3iAfYzxd3HngVmEmZ+s65lRQYpb/dRlBUUJ8oWo19UlAfnI19u7PF8eBQBF
lFeWToNZRcatBAIzWfY91maLO44caBzat/1ob7tcd/z5pKDbnh5PzAXy04xB6ZElyqX+G4nF3rQL
NWnjQ7kdTVnbXSBlWnpZPWoZBTPpjci4+FR/QHiMaW4aU7u2ZxGnXj7jl+8nrOLgudqw+auUMhfo
fqCXnyNPS9GDhsjmdNiU2upxsjv+nMp+TXmX2d1Tyaj3j8nBoAMmuLHu1mUWpmuhgszJroKmlxQW
yYPZzihWeDCX1ISI7Sh75YrKioO1y5r2NgzEpuLzm9w8SVEIvVXlLGH5ygpAltjjv4mXpzn4+8rH
vUFDp5HdPdvrBxbEZ0YMehjp5PNSIysOACXHQh56FSd3+nkgDQf1Z9PN2bKQigRFVA6Nky1HrANB
WEGmCADPedK9gGNZwI2raRk5BipVY9A4nRWOZKYH+k01r94KhfCtBdo9a3YGRaFtM6XTtVNblD95
YzoD2ywENxtPNKQc2KMt6KBz4mm0ADYU16iC+k6Y/gLK2g5Z2ty9Qb1IcTavHO07sBGurbIZIdYO
UICwYJhV5EBmzqt96VQDNHxC+hL3dAXaEpmAbAJsloviksQV3W7n7MM/F5HBCjnbS4WBTX3sxchm
z+K4RJDc1juRzqLsB2niIAitGY+3R4KU/ph+CEfpiWD692jGlbn7We0w/a4IUqu+AwI8iBIUep7C
XurpuCkTGnLI4RT5RRQsz6PWZvbgxGlXinMajN9gbgtRBwrwOr3Lbv8Eic5WT/X7vbL02VA2TL3/
7fV6AkD+aOUADZdbqyL4f81mKChi713dfLswNI0phkjOOjzYbq73lZdilP4Tv1pb+tchvJtVAgNw
DH/gQd5s+XC9RvpK5bmOYMVv25xmCqeLrGqGvf4yQRju5K1S9jIz1FygeIqlDmUjcVyWlXoykCLP
eU5VP14GNMzTHmBumHMVrHW9mfxkLb/Motgid1mWV8S1R0YRfHn0jzI4NMkaIWLNi2b2OLGdbIFK
SJPW1Y/N8sNyDsmV2PZ4O+TQJ0gYVg8shQsYICafodsXdXaLls96934ZAKhV6XbmJBAce1tQYhqz
yEDcKYbSqHVSsrR7pwoGUBtnhMRNuwBDp3wF+kxE/1th2KPhPslsw+gkkZNtQ2OX9LHKhv1eo2PT
XfSuZprBOSyMQNoy9Jpj87FivePN/2eTEE4njdr4rj+1vc52Ha/ytSBpjHi5gqZBoakszja3yKmQ
1kgdyGlr9mFVlCAvyBsj4Id2r4zQjB+NQOEYSxV/sqLXuJ/C6qYdjbPkPG6ocUE0SowP1kjNlTFe
T+8Fe+jOVwkpHXHwxEHUqw7WPoxNaXb+MyQAvp3y9RwFkm11lS6IcT4X9EAUXeJhlAU8XzEcLhil
3iaX0n4mjr1YMsDe5+d82vmoBLhMHYE1JHLR4Gm03DGrcIFZyoSxs2u/udX+WXwAMJL4E8KhVtw+
nOf1NLHian50iEYzKIkbcjBAum1el3LER5wnW7zFbkC4D0oB+JIiRUFCDxFATJvO9EAktLtGNJwR
qQ8lH16TyB6yk171++zSHUxpbPuBXoehUDYYzv8PPZGGvlyHtNmSc4HkqZF3uqJbSd2WCkKBlZ/r
w392RsUT5rKqp/Jnr4I45bemqrfjcs0adcm6+qlbjqJ+AteDzM7UEsv+znDd1eVKcsBgFxfvz91M
ARiadQOEZ9xOiSs6qXrH9K+mWNhC9ujHNQk1W72/LtH8s/fmLYJJNDCfYWetYRLR/BU/lvgWvc0l
F4BczqKk3kXa8bDtuV+3hRfHRktfjbWCGALsot8EVYsVhp5ki4syW3wqa/00edNNLA8zYUP7asrv
Q4t6ivy8zttuksaCkVKisqWEfvAVF+Mlno2WM77ZH0w9RSbfPcPnmOQ0VcpvKm+8KXHTmN7LFuGs
QyQQHKWnyUIfayCo1WtWgA0vEaNpFtIp08MRsiBL8LbF0eYgw2aIWECEcvZ/4Hz0B/i8Wj4vGjNB
Q4gZPjGGZ2eQ9zChTVNBl7377aZwL1Tnn6xFX0HGqerafGh9BaBFKWl4thS/oMDr2bCf6ROe5wUZ
MAdrWyiEAp4a2kWLgtkWUxnWlyvyDkMrjbZ7/EvLN1XNsFK2gXYQuxwXquoLfxCVF/0yN1by2Lws
9CwdNGxe3MIiRca1RGr4fk7ThC0laddQ6CSm80ahZsqvvrQxr1bKNXbX0go1oTvEhqYXOKoudwsK
7xsSQrCeI56BFQPrL36PZ0q/XWBoua1r71GUfbX3Q+18xBLU9VusCCEHxv6n9VqPnpvXjunfZiLd
0qBf64QESr9xhxdjchUkDDLCgL+cUV/s86+o0rQOw/BuuTCkYLKSAv1tmzLV+L+kVYGxN49u/ORn
Cwbk0TU4mflDPCOTYeAMiObuRheqg4kTgziVhHZxr5z6rjjWeQwBh1yOX76cv6j5s2I+IjxcMoBX
gHahW/wqOFWAiZJ9pP+PZr8cEc1ZYHlkGbVHeYO0qWpK0aeq5pJhWAODXf3XpiR0nACqq9SLhTPE
mcDC/3TpjZXt2hzL+eU7jPmFLmwxG2bBCU5W68P7a7UauaFC341UibhLz6cV05IzHavmPrlyUXP+
Y3EouP7O0uKWg5Fu7vQkcyk+67Y/ZNNvjJpk6RMnQgcrkPTew9hT/UaNZVYMzCnXsBR0XkfAWOLG
na7QMPQk/cNmGahxkrJsGP/K6BOfoOSB0ZwO79BTHi91sCvcX8t8kzsCw97hgKJVtxjQCMBv0wFP
QHBhLLW9oGy0b3xF1a6NQkRM7NSHK4y+QYs79lqGtRiHeV3Yp9QSnEY9HfIX4L2x8bxNIiAmJ0VW
iXNPkjSWtcY2C/S2LQDSs4M/13q/Z18saOAbhuBFbIpQgHzAu8sFHLLfiDu4f1ht5XtAmig5/peE
GCiAAsBSsxzjvSJ6Qw9wfvBmxudEYJCLVxnKqJ40FaLdn9iA6pqGXjY8w9XSQTY7LuFmbviJfNLZ
DLQjq5ieVOYYG3zMJF2Lt4tROoIblgAohsKcLzNFJxIwyWqhD9s+t2kHsO74iPJKA5VadPpuA5Zd
09KFCnPKZ1UYV+hLydTuLu0Sfk5GFe+HbfN++43ObEcIQ9h/pK+2fH5Nil00B/hqzZkuaFo3pVpX
IJ9zCIuLB1p8svPEiFRaDFVToLVXnMFBehd7+5aRY1yfELhrWYRZ1L07dDBCWB2nSWz/vi+zz4Ki
OSMHAZrQfGvAz54YpUtJs14dfHrZ5KN4B8fuFs7AR4BsWr6eY6G8wN+mBGZfT5Zt6oe8cR70GVmp
J5Z0kSWbtIWIJ2bi5jrb0YfvLwzXVTKwVjV/3lkLunEOf3fvxcw7ndi3Hn+lTamX2rQQ3G80TbmC
Rq4TSxgn5UkFUZwRFxY0VOrbK6O1Bm84Zhm0jt7PR3OJWDJ0tUU5ceUz3pS6xf/L00lRaS/LXlSP
4Za4VgUjC72EKeDKR8UCcT8P/+/RpLP2Wa+BKaO2zs/QkDr21wOHQejxUc0tljMfs3hqElNzxAYA
IM17wP5mNY9dJCzIwm/GK30slD1+Q5Shcge/OIifMHFO/kbTPoUBcdlXP+LzAZy0VKe4OnCO8RH0
/BZNCbeXP6FWWcFU5LpKfBQG7eH6dwdxwvPs79LVRwDJJYLWiUcrtvgz91ldgf9Bp8ClZqsqj7fI
4IlKJOvS4gvw77/eDlddvePN1qCvfIiCjUQ8vSmK0Kikc5mQVEQtSMUQMvH9SIR7ojTIB3v1VfbD
MIIjIUS8Sav6NMX8ouJNZzEVFMi1rEgcr/KN8kDvHfIoK+T6uySgmYcR6xh2MoTQZOiph/ojEMjC
jI0Y0rkuakSsjO9e6l56ZN9WiXMx2T3AlEIpdFaHhz2P8TVI089DKyXP4mRa57+UP0/cLxf3H+ut
PBIGfvyI2En3NJBx3SyMQ3qkb9Ec+Shnx1N7H4crQajEEEOUSUrWuh5KjPEAUWtlzqOJrFF+2FDM
pNYA7ziydHsvuLxAfZo+dTEo0GeBdVzJFIpuZFPeRfqX1jjekT6MbCG0O0fvhSIZQiR5KJvA4l02
vJGnCwujuIn+et1jyirr9K+cwpH+fPzS9AI3wPXxy2YPOXJ1r7obtpMS9vtQ1/SpVlLsd5bdYwEU
doVUzh6VTJlu78Qb4Q3LLv55sD83fOZU+1JNnGaTdqR8OX9FU4r0uTAmPqanEHqiqqvH4bObCAN2
MIG7sM1Aid5NcUBJbpRAVdSMee7Du0HB0llIxaQH6J9IoZjvu2yfGIAxism6ebKD5UW6tZ7Tu+wH
AOx77sLQIB5P7kbWZCO27EO07CiZA4V8SEED4gYN/8xWmYIGi5x9ZRCyDJaFLrUDVz5ee0ObNCbx
B0VsXSVNbDGp//FYhvUxV5oG2tjd3Z9OnfKq0WYqOamu2mHMUXT7GlstojVoy9B6dt/c+M7y05pL
Wj8z6E9ZhUHrp98lvEKgGBmvkOE1GopWdmBVxuJ04hmIIPw0TaPPkcre+hek1CcY9U0FFNMIA4i5
yngO3ybPpoRhsyE05vrL9OdYIIuFg3VDF+QfXt/RLKzHrAnk8GsUUckbZd9I+bjIeRIL77hsuAwD
j59Hstz1rrzUjX6H3rTOlzKHSYmLSDRwnRvfChEmDr03ZcC/6Cmdf7tO4vXhd65pE/JQNUXSAeFa
eOJV59kY6YDAXuGzDjyA1lYJLMb88TDykTlDkerOG90ZCVAGVl2L+uhocQpVhPj2CYmRRDSxsENa
v0QE2ulznvCYhbnUw0/sBct3rwpqvGZhuwZvKRflXVU1gCFCrc2gzVz6/mRpT3C9H/f2YQSB7Ptj
FHYpozgWF6J0nTpbRf4gmYv993IH9DC77lDCH/tIMh0A24jK6kr631XQNN20amXGPY29FvpzSpdj
eOmlNFcKMkkeBGIU/kvaROz5/SWguTsNks5GfE/xpcthvf2oNm7LnzxY1StZkvgMLJR4agsxeh5W
MCC0U0Wnh7RfYVc/3YjA2p1AxyObEZGlpy/w2906g+b98ClYbuDaH4hJyrv2qXLtmJY0ffwsxAUB
9bieNB41gTMGpK4IkFDVYA51Q4oVbPFGxZRw0RkF0VstKhU/C4R5I1qNzByeIPKX1+7Iy4e0Bz6e
x6nF0Ae18Rbv6pRjwSAigjH/abLatmp5bKcaqrPSpkA/AkodljmxhBobrGv6sMNlzPEWxPH1yWle
KtyQtJb+u1vQMq9tDzIhaGst4BTHG/6ftbrT+n+vuus1I7F4m1GBMxC7scoTSlrf8SI5J43UkXTC
qIyrtrQPNUOi1QOvSeqaHbvNcOBfP82GqwK6iU1cw4TBqgd4rDUvrvom4trBJM68SZUq2CwV3eki
Q7EfjafA/mF++cTh+5rscMV9chawbHDVzZdz46L8NNBUeLLswyUTTxS38NNCwWSIUMFo19RDmVgU
wAxu0zQyahEMdR6MMZI4DL8raVz6kscuSnbtT3zXSuWs8EeEoGsvWPzY+wAFh0pE10aHXZB4zBxW
TCsv8IDeLlFlAXuJpgnpYr6nZPBBo8m3g/YV2hXDUmGIaHRsgWHMldjbP1VRWveCGXmqlUln9pq3
oynP+8FTfNAN47IdXKeSqsmc8+HDUACcI6PZa+HjTtt30JcamJiayMv96Ycpzp7WvTWE6V7n6sra
c6IaExXgVEuwsc7UQqQFyRhGQNV6Tz2KniDaZnebRwZLz2Kulj6l8S2AzUiYg+oAHYH1W0MhbYNS
jTMwNwqXA8uACq/s1wiK+7vCmUDN/5idX2/km170uVfHoDwW0Qozt8AU0kVz8rvLyg8ivMDPRj2H
x0Gq3UIhQfWriH5DmMIB/f3WS7MWhU7F5bbFlsmPHjPwc8r1zQ2wnufXKaQZOQelQEBdeKB5wItO
Wr8WDK23pN0SW7mOONSokcF1+MG1eLFRHoJ7t7ojhFfKtiVA/KSFtOz4mr8X0jWRznMFqD9fu54c
Ga4ifamkPHQ9L4FoKm5vkIjwDSLsvWtgCgE4LlbdO4WLvQdix89Aw6yTLLdfjVxZnyHZVlaVjoo+
o5LLOdCLlMisccJhlLZpJTFRGcFJlpEDL1SbSInltiIol7w1YlhW9uKJco7ecXo4HPbAxbjUS6Qm
n0dFlJs5QWOAGc6IArZge07Z4FP0H3Ui3E+N7sLCAcijnK+98SD+H4ojOCwOJYWH6pP7QA2SrAXO
azSwY1RAOLk+Pci7qBD2KzAUxt/mQBbOhMdc15X08alcy4fSa07JqEbVvU2/hrKuFmPX55srjZ8X
g8bPr0x9IgcFAf8uF/XexWd7tKgGIizrJ36oXWt9+Ki6xUGP4QkzOEOUD0Y+g6snxLL1gkuFAyPA
i3deyImr1QsF+KY+8+8z3iOuZUrPxx6nglw3hDP5b3FaOASHw+vPgEafLyvjBR/drel+0aYLxxxg
II/gYmmjlkChke/yMIHVWR4ccPdIbF0+2UVPRSpg8AcxKG7qtK4ysvAKPWHae+iTaeIwVbvRFf3X
JercySQMpJLmhfn++53bUluu2pinOdVHl7l67YJa1e2+/oAM2HIqvYUJvej1wMlm2/kOZpzoNxSy
dkx9cEWw35RXjqSTB1iKhOIn1d8r7Vl607EmwHpjTP2Rv2AWzQUe13s0D45PoPAFbGXCzXdj98Ei
KbLcFgLipZZVbSHwnYDHk+aIzAGb2Ut0wqsDo4V6IVAxqlUGTFf12+ngJf5pgZBYskdB/SlytUUZ
Dfyp+HrhmdMVxTg69FAFgo7KX6ieAz/11jRfw8KG1E3+GjS2tbiJ0ENA4DTHGiVIMkegaHyYNyky
V/qfaRnypS0wdmXnwwvoBk/Hn4UtF9fXUWLDPmOCvX6vnq5baoZsdPZnXCaG9b/ti+kLquQ29d0w
EvE761QnfZfnUQO0p9ro+7NwtI2QxV/u5whGbH3UuG8b5tG4MGEd+CsEc3z6p2UyBQnPv0GIc5iw
zTb5Fpp0JsM4ebusIjjQWsckx8oUSbkP4epzeAfLKUa7HHz7b6K9svq+ew/Tc0dyEzgoZmXJWYyG
0X9Dj8mnZLNtdDpu3r9n8Gb7LtOf5pLlLyigk7ZkPlTnXB48tq/jRSJtIb87OnQvoR6ktqxiO3rw
AHfA/SS8/sD6/ZIOd65GqFOwFAEjXsbtqYNjPfoMHwF8giJWzc/UH+syAIM1T0BuMtj7ht4S8HDP
G++/GfmcCguNaYnCrb/n/WS1SbOkjO9GQWH0SRXYFKkAZ47sXBGOWbipju7kNNiKIf6cPQN+uwRP
gtZ4TsLhhRze0FbpyR2ftwyrIm/YMotQEs+WPo7nuwx+s6fujkiJEB9VNsjZAVpkIP3QAfwNSlA7
7i/IV8EH9OafK2uu5t2gdsBV7AKbKRAfuxGUPE+tz6xillTzjLc1FTtdupzyuTFgYF9f+NphXNlD
nrBJnkju4LF2xvNys3kL5lBl9OM7olGPLWcXXh3Gzo5nHvTM9iia8vxiSzw9yEjrYKW5zzHlgS4h
vLBup6O9gYsNdNAJ/oNFpTxe0IYNtjlpkcDMnuRSW8FC0fDJBJw5uuNJGepYhSA7MFv6/mHEJ2/Z
Ul4dOkPylX9gabozPVcOM7UdKaJARdm43x3t5O7EzTwic9inhI+wdz7OO0+LEPlCneQRwqDfKkm4
UEPYLzGH3QNe7Bt5R4jOCfyP92tgbatMopJe/StUwGC23prtEcIp58Vb5B9Fccni+hXdwo2aUrH+
VcpA69GD7TQagD8t8UoKUBG3pZQXVz0HERnl9zsOsXmayt9+MHTnFyPP3kuU6Az+w09OjfpyMl9p
qDD6iJ3ZoX+uGasELVtVTqF4UDZJ6gemaJj79chQYXNAPLuKc4rq/coF5bgfkVjbGauFNI4GoLbG
W7B2HSwcLuHHdjGCi5GWpyG0/r5AbGmUeO0klYRo1LHE4ZJOgt7VS2YnuEIjj44HzPj8q3K0vyp4
gtVhyGgaXVYlz3Qky6HSG1IW2RLDVF++XPQBIWphDTJFrXpmn2XEhS+35qAHM8/8hU7JkqH5G4dx
ii9gB0Xb7cNN1Cc5nRU50BWAvcRtIzuGYtrRIbPmruwJftoXrWeZYf3HurFePeAfJfNrHYR/jSMu
iazaBwEkHDGlowP8QU+gUCydXBY49hT5USuPP3LzR7u86/kmpHdlRyAMCLWzi9eUOTYNlvS7VOqU
V1oTgniu1ttSmlTQTSvjwxINcoY+DfkPA8gLfFpYYOLGfgn7Lcpn0NgCZW6fTIdqHLziA0oR8N5o
G3HEu2n2+iJh4wi5qB+fp1iSG1KNpQdQbrTFireKI0OFIhmhclM+OLzRxFuErm/N7lE0wzd+6Ht/
b56SanI+ozqGTvyaXR4hr5OWf9aPEUgwDtTPUJmLczmkdbM8r4rRgsZ8R4b2clU89bSHa7YZ+eol
yPKLcyoeGmaC9v0+CsvDJFl9GVqyKvm3CRoHi3Z3ShyeQD3Q5W0OmkErULiz6XXwYvqSg1B4t8i5
DRLekn9hEaBNMICCEXdkuiMQ9B/uiOzslheIOcKhJvlHg5OwWvGxNDcKrm7hws8xMY9LHiTlFIpv
b2BA5v/MNnQyAmFA81Z7/zxeEfitDyXF96eiRS/miGG0yo9QorabRakWy4fGyO/oUYt8qSXm9ydI
qdyB5ToQSDhnxlKhonvzi9SsVREwBhmgSMNLXa04NLUG6DocCko3eCPXXiT5jGFZMiyd8ReFWDal
IM77O2BLTxedwAH1W90QpbjYj+fyWaT8AINJ5ri1r1KLV+VLL7mLLnucD8vEC4TiPVu7FnZXIMFV
ZpZnBr/ecztfLIFjJamWPvb1HCzZt1vZAHxWmiE/LabbpC8ANtQFUanD4CtZMn4uS+sc83xZooXO
NqnqSun+cxrhRTqdf9/l2hvW4Mh+A8vlqH77CPj5Lb4KkBAAhbLMFseK46yB7fec1PQCUYbyXZRE
/zoZNwoSib6+z1TROiFJvr49YQWY7kNv5VVOsW8+te4df7+ac2QGHhFtb34qOK4+beSuzAIbHHRw
CFfvOb4dqF95kGoeSCV9nvDGxlB0EuE4Bz/2rssBDKCLhHiqom54qBs6IB4FG3eXWNeBXQBzjczL
fNcIG6aMUG/t86eGjw2Bpzv6ZoccGBP9GaPVhnkqHEOTGLA1MBEu7EnkuZwKdBkd/VGF3dqo/VTQ
db0Kq9yvcV/gvGdb3h4WM7h4SZL/rDogxoPMolPk9IN4QjLKVx1JaWKGNfP0mCmrbErsIbP9DSs8
MUnHsGNEdycywE5MnIt2BmCNuW3GmuH9ro262eMXwWIMZAHorkNE8aRJEUKnFH9qpnjvIoyr8bIw
3jPsEnXH9jQQfAjkZU8qLsCL7ZXSb9vzuuL7wW2NPkQGL19h3NMAtsZAvaWqa1GWkzMvCrtjuVJC
ZVZh7iHOKU30i++gaG43/hz0U+MOaG2n4NHI5jkurmudy+vkg3Lb9anA9VRkLpH6hweqionMvTZ4
8Ez7gFQ3AvslDu3aD3ZFY1JSY9USxg8iyiK8vnJzmHnFy0YDTE/v98wE3K3ebDBuMmbp/utK+3oM
zCD0X8jn00ysjZcTWt2fXmbeu8Uqk0fE0Id6/0LwtQ42LmiZAc4Q+6UME0I77ZOFxVEz9cA+2vi0
s/anMc9dGgos03pVy2c3XF4o4fCm4wJk2fop2b0ij5taGoJ7+IGREAx7KUcySoQSi4gPYzF5Kp3Y
TVqrcPDPCtYWlIzwqNzDBxEaNA73QRGVDw1eFKcJrd5QbEpWYvTZRSX8s9eb4Ek+UYkx0q83AWyY
Nzxc4gZZ3ETQidc4N5alV62FuhjQIpCX7XOz++2Y8GBo/N/6aAuF/BgC8d1nOK0pjSTKUUz4rg4O
feCe/d0I/QrCNUuFQQVvsTBhkFiC+PjYvRscfFFToazVTpTIKB3OhqCPt1/Cf868Ve2ZAd8qxyXf
FzRNsvn2tdqBi5PTr8R13z1POXbw7dzw92C0Qbg8lwjXuGm6+b5txvBMtldVvZClQjja8xQFG7sV
BlCuYgtMgFYHctuhOFeOq+bhwjnVLuBkoSd5QBjBHio3YfnvsvuD/K6TkYFdliyl0Yz71pH2fBNa
X01W4uwkeuYhhA2OKsUeTvWRWx1OvKBNHr5JJSo3I6YWlLqZon4MnT9b2ljxyl4PEtmnS2e99a1e
2qt6atseW0Sz+XmFXdSar9m7Nb0iIpdHVeKIJ0+E2/dOfXKMnIgOLvf81q+lPi8ogV5rEG/1wP9c
8SMjfw/DPSRxLyc5TgDkWNo69MnRl4mVVAdiqm+CGi+mVIN1xxIzYq31yIbHvm9ofTbs3A9t6Tqi
/4kiJ4QsONCVaV2hEQDGG2YK1QwR+kGCdMp56SK1Ghonxs4xt1CBnGt1yFIhJ3z19w2ITZIf9TFW
Cjds9hGkQuu3do4ysgNtoZz8EB4HdyFTS5EVAltwE/NVx/kOwnzwgbtDDXxQe0cddB+w2ed7MRnA
Prl5+Oc6qJ8fDBLBy5yXFNJK1dVePdv16+y82rd0cDk994Ph72pIzHijxuXfpUpVBq3sHQBwU/vS
2FUsxuWbBU22nAv4p0UUjftnXmCmZPWmWLvUnpxlabEwrCPifHsxOT36yb3pTOCBrxQFC9aCXJTS
9J1r74czcjZHeynPvbfx/fR3dzHjw6AnjPCIMctqQ5sXdwXB8oRJ755KNgg+Zg2diqYSY8wy/dOe
u7VX2PHBV7IR4y2OlQt1KOZEwkI/Y7iZ9Okvb98j6eJoC2sY+pq9hlgGfVN5KsTlS8yhRLhUzQmH
K05pzITgPBSPRYoIwIaXtXdB7+ogA4JfakVQcMN+yrP7XmaMg96fbngpaqFklEuPrXoRZhEKwzte
tu4Ma5AKbQPG3Kk5qUVMq9LJeQAUC6Barl7GuFEMKcPwAaOpG3EO9EPy8annbc3jfRsTkgezAViY
vPkyEgCfu+6ZPGgPVmqUgsBB/s4np0kyDKQ+ETrBUnNMQDof+ccqyxN3xjeo0eVkE6Mc9Y9dRnnJ
UlXpcWGDeXfhezJCAUAwXaYKQJONXyrh3Rae/SffzPtC03Fux87bcg3Rpa58gjWgno+Bif1cwOYG
0Kq3ZB2UNwFWKVS9/FRrks4EebHAdBpjzm0XBVRBTU/bYFeRDpcxARr7iaO53mDM3pnsjYeyh/3w
3edvl8V+UuT1zypqvzB2Au+ExSMOUgUyI7FGbB8xzsV67dS2VL+q/Bek+QD1uUEu5F7W7zoCyGDi
I/HdN/QuDcIN2caehJ+l5RyEETYe4qYAOsvh3VdXs1Q8IgzOZF8VB8ZJ6juklHyrfotUGXgE8JaS
tTIWAMh7yU05SD5DwvW4WEsEa0DM2/lU1PQRdKXGXGixtsZYR97xb/AKJ6DOsVeMX5mhr5TtnrO9
+1XkIbMDzwpfuMRHHuEx+sAru3S4GetDwGQM5+37YxLJeQbnLEFwXdwMcHudpzFvrDedidmAytSZ
dJgXknNDbRkHba6hkJDaLApWGigfWsGMb/SloqePOiX8v5908qwEiVVa9C7i8RaWeupcnKY2WuKM
W2CxDQQYsIQ8xkZ4Wg/NYgsigPIo324wB8ElKtB+zqPi6cFo5HSrEtFV3M90dJQqaWb4npIBTh81
xutbMuzaYDzuEseVASx1mLv8SQYkmEjOr2RDaOqIvZU7No3ZRwgd1P3AIS8QIY9PJ4fC/qeYLquY
4oeeCzCm8/+bCCfWPjtgHEf2fScQH4myDBIKXrvs0Q47zMv1gOC2QkdXBGfDWmhsgi7v0jtkHIPf
1h1kNdlzGYvaAxv2U5Qa+8zGAB89TU02XrcPiqSc5AdiyuqkTAylNx7bN48iK0M2oSJTjlLdTIn6
w/zrxIGScHUtq7+nwQW+cKtA2rG/cgnqClioHp0se8FRJoE/iz5tweCoDtNKcL+Nfcb0c4een4zW
APm5jxUsd5A2DjhXTSDwCT2P6wPe49t/VtwCJdMN4eD5Je9CfRiVl1FOLHWruncNj+AgLvFE7htY
5jnWlijuZW5Cma6onbiFnmplWKnywq+djeYNKbasQbro/90I8xRlmhuly305k4KNL7VJ2LKC5qV/
1TrTpV/cbjWfMhixYP3LXYEAEWjwwHuU4dENTqG/cph6EcnX1DIpN4jlSmZqn+Mqtyuxg6yNgAyL
BeaXw2ZZphL5K4ecpa0PU2GrXYZT4XVeL3JtrToNl38rz5Cdi2BhorJIz74F9fAAXkxJtK3/WOdv
JYh0T+oibOmdZpzykdoFsqRIjD42zH9Jd3F/vTOOLCYOzCM+sr9zWROIiW+TmBNOZi597vQV3XLf
nNLuht02pDzVKBJ/i3zMepZ1LGKUR8Vjk+uOeQaiNbyy51v6UU9fQFx9Sm6oXOX3ikK1x83HpClz
tXNYbRtURBloZCTysIxIKF5CILR1J9sYOUWwBYVwjmviJofHUM1v6lQHLBWlyJqsjwEOSVF7/9J4
Fe0tuoIp70GyDDa6mYMQbMZouwpCsC8WbM0cFTk4kB8ThVLqNKi7NHYP9OQC/LERj8IxK9p4HnuM
3kHdG2bZdE1MSJVKhvqhGvfAWN//2YBT7tUwnmsqiSFMYbG9f5zOPKoOhsgohjh2R2BgTNuRcfcB
QeoHLbAIl3g2mU08MKiFXYmUwU0B8DmP0rFRohXl7HXlBOSisGTlT/p7N7t0NuZQ6b5QqPCiRWfV
ClMAw6cEdPNKZxeZbzMMIN2iS8FW0HqL637w63wrWbIY6GNxxFf7sLjX59Sq1qC+fTyfjy+C2BSV
oMI4fa1fBU89oD+KuvJtSBXI9QhhHIV4KJ7P4BJ51anxlGsfkR7kKBMDMSVAJRuvkHU7A0wJHXZs
pqENDqpMlEDoQuNYEVezjsZCRDqLsaOrygRNxGQK72rbGcNVpRtM5w1vnZVcyt/rTEtT470XwOnw
GRCtUz0EfrmbnnWtlqKFGKiYEc2WU6iKbofc1gTakS7iQpPcx7YrCRUiFukGZbrw3spICZGDhl2L
54/zyAesZP1wgwe5hQQGq+p0JSd+q+8BRXsjI+vKQWBVw9zLohuGNnE5Lte5U0ywEOdlWdw2iGMH
ltS7Xok3XjdSQQbJ7cbOUXKFu43gL4ODpnbAqT6nBHPeDDpNL7orQNj/mIvicRKKKajpZ4m5z85g
9YtoDq9zXj7zhFoFaSAdOYYSvHSdugKJGaSjD1c568MmNwkr7RavJF4Fxv0vIJO7q76+PV7gZAom
cwfbw2wol57y5aMvBJ0u5bNqESA5m9QM0IG8WMzd+MPfgDn+RNXjpoTOPROAspgwzKH3RooHJHyF
YLlnXCkCsrVsJ3gTdIm3XnvXiJK7/fkPp0n0SBoi5naUlPDA1piCAXJxEUE3QtrJnZzfbKmqCsmg
6BhMPiJ85NnYr6H0yJ91Y91sryFwC4a4o1vPbYNzYIsw3s65D2pJI5/L334U7f69Pk3b6GmRDqFZ
6GCUav8At5nC2DkfQ4IEQZr1pqfH43bznlCO7JEXtMsBTjgq2MnZ9fkeQpwQ9g6ppG1SpVSEBtVa
kuDu1xge8RUegKQxHGFruB+I+THiRfuRRBpirKUPDapbZCuvWZ9k35B2ByfFs1s3b+Cq/14kP4f5
YGTPqWCbSYKYyHWRlmu8+Kup79WI1HNrgo9LN/wIPy1iMudWG+wMgCCFZNTl1Tn5NRfnPNIgcY4d
pSMl9XasGEcWI1HL2Ke5MrJqHsQO6CXUD3LecZ7LuTqU0b6IqmEN0lLBCCLrbulkJXpJcybbHbIX
1opP/urhBdufrFuEB4PVYKdkGGmAT/VHU8J7M/3YTqqjthLuKTiAdw3yloeM85Dy+WwqSyxPhs0W
7lyAXXfOrVhqJLYNgzrmgibE0mq4BE4JHYu4v7ZouaHnR/q19OX6NF4q54RI4nRWGVo2tmMsXxWh
3rMCRr7JXrnkQ6rLp423LRpiqcYiL8Lo3XtUMfczKbeOEES1SzZiQRPrcbwxd4DFDq4D/wJufUjF
uReo/edVjdLfKYmJsY0e+BE32ZN2QLzBD6TuryyYAw5oUGKzNxlKxROFQenG+wHa5Y2Hewqlmd35
9IDIpgl8vu+S/wbdrsHlMkCGsZkesM8ZlhJn4XVJbrGWacWiH2PjY2+LKLUeInKwj674rgBZo5sL
G7ZwIPUeXBlfTVgwFKwJ+gOVJxEx9xHfNxbsP3ANY23BqDFv+c3PpfX9/4ld7DfOyG0E8f1xv9RH
G/8HM6zU6DoOebC+ptZgRaYAFV8vItHi76QDMUJ9NJmnFOejjS7P0PQJaj0k07Y6UL1+FJUrAQGG
KgqnWZLgq8EMVgosJqQPRaXMNluhDM3KiGNSI1pbiRa74f79rMPgzThVaqYmdBMXKWlhFXtqIpOc
FjPr36IKwoyFjayU7F6FCyQd6nkQkufGO367TiEKPfx59EzllnTUBrX0a2SF6wtRikXUovlMdqTA
PQTnYHsvlNSpVv7xbI0vjIumgfRZf+22hucsinIl+PspIm7VGcnQGQb+urUadnd8JGqKxfFxLHnf
jghcfdSg1l9rFNEKsLHzLHUKizf/nV3Bp4mV9cYE16iV0IhsYE1MdZolF48YK7XGpumYtZXiRJym
Y+3kpNESYSHa4f4DRhVKaLrU5NDCZLkOkPZNJs6k7nkUWfH+g0BgQW3z3ouLqL2A3qhEXP1s/vVK
RPgwp3UKLx+cIWsAiy8ocDXN/m9q19EXO8cOglAvAdsSt6p08UHggvEbwZuus4+20SEuH3YofrTy
OgGMRlTnt1/JHz2uegMsJ4GCYZ1hj/BYXInb6h+oFARw6Mje1EH9CeoOfv31Bd7gV2aOrvV2q2R6
GfK+ON0RlUMilbtHhgPuxCrghVvowH+cnS8TaPtColuMJMTttxqhvX4oNSpsxIBjLu0Kx5gD32NN
9YsmKdXlzLzdQPo7tdYwC2fKf8W/JiJtp1aHw46FcDMmkYY98ipRbymMc4MzuVze95N5vadrKQTB
Iy9RK22kwTsdDQTa8vURXAfr6V9PC32jNQaVSWyl9i2FSZnM4wrrCeKmvBlJTKrvZP57jARNF8E4
dHmQecAW1UpKDi7STZnD89fyKElTjfpXbhuoSohLEGalNs+Brbap8YlmxpMkxWHcdlL1emtY2CBl
yZ9THdJ7j+JrxJeMnoH70X6yLiK1DvBvnGuackEVD47qUB2vIjU+4bzxxCwEAzgR2+qHsrUdRTf1
c0MHhpugAsCwPq0VIVEXXisO8N406AZGfEaZzF8MOWAXzVhhG8otE2Z4KzANXTiOvSNxmA1AJbYI
FMiAByyKO3ATxa0bypXQJaXA9LTgIIE2SB2bBUdb3HY+vD9AxU7N0hSDXrp+do6pt+N9biY6pkiT
P0iSJ0sqrccChrcOP1+9ZjXdnBYF0JVYmKDPg1MO1pXCMmPKQCpPTUSxsTlP/fnYUNqXz51rrrx/
vEHfmdwcU9Yv3WVNRPx2RbDY54nWjn2gCeg3/JURlskHHkcrdLs94ifJv3HHYMk4MNAnYNxzpPrp
i7/yXPv60S/7t3WKxFaroG1eKOicRf9cih77PpySIbeY7Kl6petiW38V4/xVUXI0r/h08rH153Nt
53SpwUNNWzII3uRZWiXN61suQ9Tu3CD8sly8ZKqWzbGSF3eoSExEQNnI9zfJD+OASdmVeHh5jNoc
FTArj4DKEq9UwL0Qg5TP3+pOjPq+ri9SlknEPZdIYh6rdBAkVCFqqnxjwnrfu0/txs6eBjpyTytm
+soNzp13bSSND8iRpZmz6lsbfMBvd6X3A5TjspcT0lIo6gUyqzdKxGOv3tD7veN6HWFTMYBAiuqq
5//MCOJG4OOarYVsOQ3T0G8iNISsNafaBgc40XalWscri4LwP2qqXePALQuyAu0Y8JnI5Rec8ZV+
2a7FQz+E78CCLqpd5Now3q6RRwRxOEHFJu8w/toSX3u8sHn19cNpRml/rp695GMEMzw8nPGhQl1u
bHu4tddA6f6jxmj8sr6o6ohisdw+KbEgKWFYtITquV9nePIuDXQzuFzpXF3r7KxMB3/uM3CnJa+b
Y9UosxrNnyUp983JOKxusPf9T/QFrGw3iSFmf7OUvsB3DFsJhstrxkxxN4L7dNiBtJNfhh2kb0aL
TqJ06OLdqAfyKh11MzsCgkX5npfUGOqRrILiFpnyHaXHHfWgsrATHwNMuqXWa3O1B0v4jrYnmLPT
sWvLSFAMNBBz1mxjyJZk85c3bD0sDVpKcST3FGLOdBq13AY2KGxtDWRN6ae1I7jP8eTvyGmWdZaF
5WVp41AQM9/9RW5ApOO+o7quAjiACUEooFCtPMZAp4dkSyUS9wGR23FrJD6Sel5oj9T74CkWpIn5
jVx6ktmBuLOgTE90Lfy4WtpQQj+lqkrbxNARVCs891Eq4gXX9KXl7AetGG9gQh0dQzP1ggH3Uzna
QTSBzSFr3wNlAmyL1fvgJN9/IT7g5QObm8NrEvCJ3JOTxUATzStxiDZySbqed7Mp1BNp3l3T7BVj
2dluDD5d5GUZ454GZ14Ila2uWoZ33+z/Wnaa7+KxS+H2YZ20ThPTjIjfaeYLoUKDDNA8IWPrNP5M
Ygn7NGIBTtrGY1GvNap0AfaiS6GI8gLKmI4th26HnbYrOEwBve9D+e2cKLjkVjIwD5j27nQYSZNA
hh2q+Plve7ecnBu6ht+dT4/QgaF1/MaUETL+V3DM3xY9zvNkrKVwEYsIw9pw0ZIgNfg/BzeNgpHP
nkT3bx57JMSCb+7yA8hNYoKjsRufMwO6PTDgRNVBGePWHBeSENq9MDrZ6kmNz6yf+zEb3bOc1m76
6m6aRUvTDOPgTtaqgWItG88IsbMMui61CQsUtkUSOQdVgrZKcU0uRnRZQFKuZBUbqzLWA4loNUP6
LinKIS0MBAP9/RtO+rwmcX10dfgfpNkgtZ4p7rx3iKXKNjimfr9XIgmgGHP0iQGy5yAi9muhxreJ
ZMfyvxzw/I/uKNn6/aVixC8U0CLXza80P37G1mr1oXV9g0q8BVLtIWWfZ+ZObTd2J6PTP6ifV5MT
KLczWNectCo8rYjLDT8aPRxQ/E20KNDtQOLTLG4teSMQwLXZFitrsc5Idh/GxtNLDFi0uVKDsaH2
w4Ks5xNxK5F5iqUsmZbcUu3C11QLGFFNPDYTvW01wNIRd//X0Rcvavl22g+Y1E01lLKGxSviR8C7
2lk0uA2VAadYINpa7ulds2FzGj8wYdTRlK1eGkNDe/EgmCsF/vqPADSkSo4VGrjMRsC20PGeDfpT
0bwE1Evg5Uep3vMS3ZnvkwZYEh4Jx+FtR/xxkzlVSl6XbWxADXIHMOqNw32/qAIiP+VYu9Td0Jdt
GedEeDgHuZiDs3brDswO0lVnXGnhf41L1ODnDyJvq7wLxTj0oRjAtuHyyW7Dtfj1wFT6j4nbKqwr
1dLYL5dSDsRA823AUNfg4zcppsz2QeWVz/sDHZjCRomIl0SCwPcPtPbK5MlCS5NhsfyMiRIuAuFm
4eVZMhwwY2g63iqJHmWjw2MtEl9gF8/6656VH7i6LksAdmYqn5IdGZu3snQfiAMM02MjwbKApGt7
iTuOalrrFOg429deXm082DiWfGuHdajs2ESYJ0DsUE0TWpHY6ouh42zniNGMXbSjFn3elirS2jsT
ODpG9FmmUjkvqYQGKoQ1PEqLk0Ge4ve+9IuVJAPpwlk0Xdp2Uc+q9uZdT8n4emb5+htmzjASM819
ELQAgzthB2tnbKfGGVWX3qFw91lxwC/PCJ9B79X5p3ogsjEsocCtd88vwp6K+zQy6gqallyZXclX
02jwDdKWvoYDD0dVJaV23IQPjhO4AI+k4bVU3O/68Wfj4tphtVGshDQVAE2kslvDFQLP94wPxd9/
DIpm/m4e7LjcF/+XXk4Zdr/CJ346a2jpFfTQrAoTj/Y7Onwu4OVYAKuhb0tHAovzGmU8+YDPTwTE
yBLaRLN2bDvVrvKJ67yiRbf8zBCH93FzcmbrtekJ0h0ny+uI/EyvK7Akf60rSBVPxV4ObjzvYOKK
6m/ORnolvUZ+lg/MF7WRvJXpT27M/cHmX5Bymq831XRFZYM7rITdwOJYjLmDhPKj1JomlxJzTbF4
3HIMEP99MBNfOb4l5mQ3QhXCHAh4XoeRUMoFTErCRbBtMnz9brxtKcjq4av3edPx/S6mID0ABgGX
IPbDvdfGOe2fGZ9kypzilEeEFilytjHJ2mUoGc/yJG7rsVXcTSj51AU69gMGouzwuSsb6MJdGG4C
KO/uukEOh4C17Wj41iBbmB4dvF/MnL4PnUiGJW+454Tu3/GzW0oKPQqoH9tK1myRZU6aKRbcuS3w
Q4iC3uStImhi9bHA1N3f0gc+WV4imjC7mXy6qbLy635GZsDnzINElS0At92h1tAZbg1EZnYBwezI
D9gXH8N4aLype7c7LVe+eoSXFvKLw5WAQXpH8ImAhNCJtfyzqIl2YWdCUoj7J2J1Sl0/CE5LqPj5
LaWVTtoF8ShJLLChYr9WD+e9mHN8h7Q9hImeSaEYcNmEj27L4aSN3vLhRMy2LM95nc0CRZgEl9ZF
5++r4nTyVhmrT6BaCh1mhPkwoHG7zN5aRHom6n0DKuI1t6Yg/CkOzP+nAINQ+3OLSD0CsGQsVnI+
tjiKml75pw8Cj0LGgkh+CJuwl3JPX3xHCsOThv+KNzE16mACiiworKHZ0qzzFechCdYJX66xP1MT
8eaKD1kZK1yzWmlaSfz5i5LmfH9iqckrjGI1NLIXvW428+N0McFnxwKFFihPjZqMWUpWFlLFuzLt
SyLfK6vMMjuYF7zDsamV21+SXjy397ie3YN2Ekueq0UilnNOqEYWxltibZC7YAvvLDtNYrRZw/Wr
LfJFYqfLNaGR42hvEBeM6T4WSOs842eX6AhveNCm/xtn51k8N2iW3Z4SVoXJIXAyaC+u22/R6kOT
FpXztHBsB64ndDnfsnqwayofMvc9lb51u3TEqdGjS4Ffx99qyiWaycav7msgJe9nd/yqVTHAGG2n
EWgPqi7gpOtzCk8S46Ewa71VqIwJwJd6BtE43p/qLjcpeeyXUcEguguzobUlWXF4DIXsgG0F3znc
IGtNnKivEBC0pY1XuW83ppf0V4Wh3hNvV8eS6s7EsJO3+25D/K6KrmFqNkGqk+mZJuk6xgt5XLTR
aOEWtLsy3dilcK9IFeGl1ux2khXyBUMcNe2R4z9rYvCXQPzX8Kk+oHG7x2vqTlBUw/Z7z1y2zCxi
htawddDGebCn3tIkJtdfEbm/lUu2VkwJ3LbNyu5u6O7LP1+SOsBw2CmvL9L7VlnLjigQR49lY3QM
uFNloWFBM380oYi39ZV0Pje4OTogWRaIKDw4dGRwKsGsmEgcocy+IlAdUFDXej8aNn+OMxWjYqKu
kAEP75ilqKoMNcubvHPP+j8hBd7B1fTszsvUercDIOh1xCc7TttZ1VYRkipIDFdgex55jgmCwPEK
YlRXUMHbOjCVMBpZRI2BUddFUeRuLEdN4RdPXOxngba6fqVw8XK0dK1mZZSvbP4Y4py9+AZA0y3s
keMHm8e2+IvRSZH2F3LC1IHyTo0FBtFS02yZr8sJEWBIQ9Cf9+CohGtY5ksqhLZN+Lu/RiKU+6aw
z+diZymgYcQAr+xPNTS/4lOoUHOJex1RRHHiQzVFlipvGCTrxzXwt5wi0u2nqAXCXqSWXTZDXqul
Zme+K9lfiPSlJdM7qPqbUKZSCChIcSR+htL2sz7BjKgpvpdME7ypZqCvMXPA31r+mNS8V84h9HHo
WJLA6mII1eA3BOLE8qNTGLiS74+TN5/98THVKbA/cT4mtSuWxB/nhFoft+0k1umHSnJR5TL4PmnC
kMek+9lW1JXbxPXECu4IARcr3In4e1Iz5G9A5ktFGhFuEqg5JApuCz6FbAwJP9xkhEo2rbD0thXZ
BLqmXSoUQDpIcRjVkUKlJ3Jq6cyxozKaCgkOV4F49Mzbpi5/CwknUdLIPatUqp4gwaNRnRJUnkKW
0QYnAs2JE0+/e7Os2cfon1crtLAWvNVG600ZBGYdNTPlPnTaHy9hpWg5xx7BLt4MVkTz5ZuCRqgK
aMbkbV2lzvQu68VBHg3MYrSurBKqskLfrA5taBAUNUH5awTl8KqGIht+rsYffFkza6/6KCzryi1t
xqIntb+sPzElAn1Y2QdU+8pXxHe1UcUHmLfwpPWRxVnst4pPqgtxsWLb5eqxJEzMM59wOL4tA/Hj
JYfiEe4ktAgbs24EiRDEvGpk/WO0mEuww0/dYGq7rstnr5ioKleGHKNP+5LcWn6uf1c84jzFtnsE
QOZgQgWSQQ9WbW3g4j9CEktY46SKUQ84sN1UIDS9IME1J1S/EyXJEoeX+7KiSbZ1D1wlQGIU+Ea4
6JljLiTGdNXuDjwu1r/DX4cl0/Z0r5Dg7KJ2nUb9rhSPUZXO55gnJamQIF5bPoGzoulfAT9JdQcy
LNxNLPXvALmKjGutNWdbCWtLv/WFTuVL8T6WS9dZ9L5AsKysP0oeFy+HLeyKQ09cF0yoMPpad8rQ
sXMU1IbwM8M/7o1mZ8cjWTbvUIEzI6d/Hqqaf/88TLugW1LsO0lrRFL0OdFuq3jfBxG+IhM/4wIG
vzlKVho5pw8V8dm1uzsC0j2L3/wN5QSqqSv/QwiUBPg45VJSkmI2iAensiG5Pbx7UrEpipN2M2UA
PHuxxDAe2wN/ijch681HHuUkQufjgrHOYyFIhE7kOaNzi0vkQfvR+utTFmuHxVzHDcu8YqtINg6X
2f7GEboTLMjOV0FY2idBS/vHNb7gUI8frFVxscftu9eKMys69q+nEmzv+5ZP5EoxpBDQJgcK/Yx3
6TBBWdU0eHvOtfbaZYmLuJem1wBx3DjZh5nnjx+upb86fLFFfg4Xy7S/n+9hh1ZuRp3CVc8RMO9v
g3/33WmI2F5DFh/Y8fqIqMV4cVXBSjA8y5Pr735/J1lhqBjujFhw3ZAFEeB0tEbPcMhL98mJwgPO
T1HsBoghXawIGOMkHoISc0wEWf/enf+LFw6Anqv+ySoi1paUzxwMo36E6c9aqr8uSk7ZQ67VxaLp
Vmq8p65w+qDmUDPVhT8K5JxYoahuM76bzxv9mJa81jq7pDE4MMoH8wmVftaZIfV+usyU3t/DLpET
k5sswD+/2eebBqZHgxgZf2yEkxYIjwhrFAvQBU4ZUlpoCS+p1pLjtAngl6EQ4XjsPt8aTD4Vu9iZ
DsMep3co/8CT1WUjDBTP0K9/uTM5PdwDLiPniGq9zl1VGn6wUMWx1WAUP7po6hGrcS67+e/pO8P2
Jq2V6WAkYHgg/9fRGSXUkbEo038lSTWS3GXaf24qWDQ0tWAtcodWhWrwHsBA4Mih2VcjKjn1QNq2
HACU5NZbrkhjC75QKpBn+cuP/u24rOHuHhpOWJh0G1SIr8x7HaLtv4oeRcB4gsOCAMUuJkJOtmYY
sHD2nN+d2umxJFDtBkVBugko0Ru/+3cjsvBpiEAfwnUae4TW2yeWi+axwGt+5omDIQPt/g+9TA8b
3IjXZjYXv5x0ssBjke/WvkIe/hx8ybeI0sZ8Q7p7ieev+oEyNnnn0LBvv8u6C+nRj38K3337e+J+
RJJOdlTP+0b0iE87xEq5v/Ao24aufjm3uOZnQx0HwhoCBJEXDvbOJfVM3YX2kVkwutiY4Clo4M9b
62XQoESBJx4oimcQWRbICf0Aoohdthk4fGBRzKy373d+wwQP8HHhDnSf0p6uLUwvqHKrXzueLFxe
E4XpJkbjMnKjsoTfNc32t+X6gAhbVO5qB6POAobVXd2Xudh8bFFgnvH5XZSY0JhnumlNCfbUQjRG
bXoL85vBIhJcqBkPAAFuoN2h8qgoa0q1Bppo6VB3+atqA/ntvW7j1FKAkk8gPJD2h5mJnpP5FnIR
gdnnhD/CPxXlF+xgHVBoeNjrr4amcmuqu5HRUokqB1wtcOsvXA47ibhTiQjIUFS1Ejet7dhMJnWp
ezwTUDkS0PGeTRNVNiIG2tSnQrbDq3bnrExZVuIFs7p/mmH95KndjENO0v3sdgzgq8gD6gYHQb4F
nBXpLiOcrhj1pEoDpKTe7q/FRQD8gJpHBm8GbwKPOIm3WeTo1y/jAG76x3z1cQviIOXF29mPylZX
i3qe2Twl1ugOqSpThG3bysEAHBg2WoNGsQKygerblvmlmNUf/fcLeZ6lJlwzSkPq0kdZtdkeIrj5
oWahxtQtjVKtjcJK76siANXVoRBBbBQqiku3Dg+VKlz230FlmOFPa+jQkl0xfd/OhLSW7EPnfKyr
xaJXnizDOP9jzIXhnUa03WykmuzQDI4KE/syFwIhrALEGLaukr5MhKdauE1Eg0mMtpsco5RkJliM
WBz2PpLgdZjU0AqcZnWmbsSykKSb7/bYDmstWzPIrAbQPuif/Nza14O5izkaWS1oCC1tV49WjIn3
iu2Ua3mitsUT9Yq78PpFoSobgims/RYWyIdZnoD5lJLLFGUkfYX2QDFO5wnH1Rbb3K/40dQhPruQ
jy5bLNTlrz/WuF7zF8S2JVxqphTzzFBZNMN2qklA+ZMVm1Vc9eKeeJsu//6hpCLJD7fEz8aa/y58
y4cBlukGxXGlAxow5OjK8F024Cpvr2tsjTiVy35RFk34zMMQqDFbsrN/aduT713/cOhisijOcgh7
oPuXUtm6ox+yrgfvYKUY/T6O+VnTrW2L1IwdwfsnFSli4Ekw/y08HL/7lu+tZoAarpGImtRFXHaf
GOrPE/ZA8bgnu7bgjFaIxuk2tVuV+yVaDl0TVQnfywnZFjPW8PX6aQ0fcgxl8YgSJZ8KK96a2h/W
Xq+mTUWNARTRC5LPc4eTDDJBXbMAIP/NG/BS31zJzIbJ/LNunNf4JADqoqBNhMBUp+jWQFsjPNOq
k6r4TAOSFULSMYhIRRzkfyqjuqwuwKBxOZ9hs5XuiFzYDlzFe1gE/lxyNWxEInXfpIIMkkdTC+Rf
n4QxToMjVOuDHdbP/UUjALk00bSvV7kvMUXE2OQkvyBzi+nt2vRmg00h9R/5WOhkKnIi93wpi5bK
qLJC02a9Uvj7ZBPwEdGCsbPgAV4H3DHV5oSJYR94+CiIHlKokZ2HgY3ZiKivoEzbUN/Xx3hn4Ouk
+4gUQg8lso2FXYjDfoA5Juy8WKKw4VrwUnY7mlMk7sNhdVyRlaCcCpK4YUuxxRUuqHJHWYvH71OB
AxnMfZswcR+YN7o9iQm1y3EjWCQxpoAG+aVrtAEfHz/snJaFc8azJlFVj7LlKdQZqDKERg/9PVWq
ahkgF/SGB1BtpSR0oMDb6237ecPaQl4zfCPcmx/3ZeEZc1Fwtt4nTeAO+My/MsVYQGdO3vRRZ6px
59E+p1JauWPUjY3EJeLeX1r6C8gfO4M2oBoyg0Epdgn4FPX34tYdWQFu2/yjvutlghm0xta9ruDl
jZ0bTQhVebRpm6A5PTitfKT/QQ87+4QNM4wLeNSbrEcdr4LUL5W53FXd2AqHkoSJc2Pi+fqTrqeX
Yyao7AzDYNXInZwse+u+GgT0mR2bjBPOFZLD1wGZkdI8frT+WFcea0Po/0/LpRAXyDu0n8B7IUTN
SN/pFf6u+Tch4WtTrYEHVY+yJHcNwp1WjU8GdqDmzmoiQqBTGHMnwk+bRWG3sFWETWAhzLP2xAzP
hC9hCvb80G7ttb6uFXTbgRNjeXDDNG78exSxyvjzBYlUJ/3P87DIbt36iSPUeZ45/j+MILuNxNq0
nTMEEgt6RGeKVX3R4fSc7+PsST+/Tx1Z9wYLt1mgZeMQuIBVix+nw2P8sr6hdV3F6zVaz+xATJgZ
klQ1p+trv/irO6vxqxcNujJwFIum4m1N71JtDVT23Dcmj/OnnNi5uB7UBm5DI1HUJbNxFoiNk5b5
wXAkfwxHnFW2biNTznnj5apab4Sp2vwks3vT4HSywfPF5js3pFSSyJ/xdyTQxTW0QfgZCoan/Cdb
ROfr6j0+CFFxd/cMUntpmxaz3P7L8WbFGfAFZ0ZR2MxkMBGTWXBKAtmJ+Ol1NWaNb7n3FoIss/5p
sW4TexQ9gW8pJKWSPQv6Yzs7ctXh4FVKZav4qdMzsRTeqs7D1ch5b9Kgkuzd3/KV5rVG6uF2iw84
WX9yd3QqymFJHTR/E+3QEuU6AGVgBmc1St70BYOv5MJ5gG+kGLHkFNopFH2x83jC5tPuhU6Apz29
qe6x/5y6jaAFO0w/FmoqUZ7V/OWa1qLrPiUyRVc2eFVwHGTj6Q+p0epuVHd+asXEz0fWUMyRo/vB
1t80fHOXXCOWhDb7JR8iXk7uOy8SRd/pgASjb7p7E5b+bd2dwlVoaKh/440OwSx73grMcs9Ggi2i
ibkl2EVphOq8SaPagkPAG0Zv60LppnTiMzsyNtBVoXocV0MVrKy1PufZH/qxrSc56QP+19oXb0qe
Xa2zA5ZUlYziO1bR9w3n/5tSBEy40m2RNkl/eI/2GQoBF+RHH7vm4Y/OVnQnMCRm5wmzbqh7Vptq
JDlJca0p+eZE189ZvEkBTsCYSLJUqOgsypqSCibi173M42pv1zBetRn3+2wt4p2jhMvjeVXQQFiU
5Ptb3k0Dk50nBCzUgclLZYIeb/felHfVtYOBkTgfwFB5B1lOpjGFK5V18NThK4CtpcYCcw4Q7Uh6
7KmA7jBs774UFxp7E2PHTNkNl5Mcieb2ajwyVt+V/Fmdg50MRru26NuneLeIqobXwx44jsj3pRou
3bHR4Kh+rzwzGP3IRqM1s+9rnDM/PhvNRjIsnjyCFXHMrQR1de/wqoqm4XF5tAYBPeIrbI60m2Uh
lyoZsX8Q7dQo7jnApqj6/+1h0ZjCHEUj2Kf++3dO4PmL0uVx87lCtyjLXgwDLDprVeDFy/G/R2m/
dbpOJRHOixc26fCQWZwlXSyIOoSwAsPInp9omA/gjouB1Kxu36ty/VDlewA3nTW+kltdmFePvDzC
0LPJIvnIo2cgOoecawaGo7Yo3PFcikNZJ57tarZuwIiJek03b8R/olO+IY9E6DXzcYMtjoCnKEy5
y+7SeyYsscW7AZ9SGVLUG1rPs/p7OAbts+qgU4m1wziCBg7Oqa2s038LnaqbhBBXUQQUTpm23ofS
8sWxPzXnND0Shn7MpmT2PQkg54n+PTYtAYd8dW6qJ7S281mfDBRNpmoqpValE0jN5N/tYN7Yb/Uh
SpL03WsqnFXALsieoxf1NIxLMyvyDhis2y9K4c5MVwnYhAuHff73BUsgxYQo5wM1JgB4qkF8lrs/
Rl3p+s8bOHq0THbzbNK7PYtt5I3qvyp3JzgdH5Nxl6UIM4V/c3nhIX1DehwzP8/FTKrpqQIQdvgM
x53kMJAGczEbLTz5CNkMQitUluPNhms+OEIh7VhaS9n9U6zAbA8Q3QQ2hwpg8HM93/NX39FyPNfs
ecUF62LO48lMQl8zokndhvWKEqb5RbQuj9IzOZ4zHhjyN8Ve7xQWuRThBnV3qGkufF6xGLFlxm9c
49Iqu0UXj5xNprN4OVZ4j6yZupOe/S1jCdTMFVTMJr2dr7S9RCz3HV5jBBgsUZdqtj0sqh7jiCy7
PDC6eoR1QNK+WVGX1ukIdWAUNarBHlVgjZNOFEJgmqG0bUVuorJr2AD6dbFNnR3MfqzD+I4CuGnk
ZSJ7nZuyV3u7zaLMNPqb/Mxxg1z61Km3qcZx+OanTByGeK40AlYqCKIdl/tnOF8s5Y8pQ4X5vc4V
g1rwbXso9T+ZCp8pAkIt9QrGU4QJWv6YwXvFzFzTROJaDuksVdLrNcRcj0XRntVqBtCdUPMo7TXW
Kn0rkXIzwE9URjprQnIpqzfpWHBM+zkZgtUX6zrAT3STy8Q/sUbtVtDOYWCjO1uAcJcSI2NvFRyT
5jcmkLl8IWsIsdqo404o0D6rKbVoXXw0ug5PZayJwWyU5TM3vKMHlrr+HvejclpuvnuGfkxtT+bh
pVB16yy/XxRSU7J3zGaISicYsYPXfTByjM66JkbXlVrREMajeaVrxv9ZWVB/XF5MTBn1Ws5xA6GD
fXlbR18NLb0nO98MakWm4uIo3RX0v0IE6C99aIGD4tM6PG6vJqJBHF4olIyjViBEtFHNPcg/3PG4
OlZvm27puuX5paQbOD0g2hpJ22UXVEth+76uoloqzvL+cCZyTDoMCvSnMLD2AN/iNRjUZVO1ZQpw
d5gt0NVbvLwTzXol2esQG6ebwFPaELa/c8nmH3mW8pu4PU+vunpSBNZF0oF2COB0ogFsOiogL8Pd
jaJN5IESfmk28y/0CKvdhiJFk7FqZVJi/gqR0wzbLBfAWONtvEmZvYgew9wZVujmcmi1reFtGxBK
a7jFowcBQkI2OrTZ+mwNU6+WbNZoYSzbD3ssvTtHQzBP7f/XX4QN42wsnjsOeUqTRsblgoNb0t+C
pb6dIPCBdDN00B4TBYanvQQ2lbrOBdeWzKCcP8Vxy26nPrY9Y+0avD3CqdZMC90hMYUev9lXH/jX
2rjo55Y0sSb1BLzbAK4sRUPPEhWe3NaJ6/XwLDRzHX8mSQRGb2yehp01Ea173Mb/NlSQvMM0wBgt
QODQIaIWu4b8yx/eLneqmLG4qWjE96zE7vynhzHaoaSJx3JL8IsERR5byHPWhXhmb2nDmHHzDeFb
8a8cD4CVhPWySsjjugTzIZi5Ap/ZSEySw+p8ERgRpMbM7oY8Si4aA/M8Zmz49ms4iFXZKTDvg+ke
s6it45h8Ri+9/utaydzRnS5ALjcQoAldcggtCA22pJOXBrpzh+4AP1iJ697qMNyRdgx+WPOjSU/6
41Fi160pa/q7X9si/9uwjc3wVqIgE9i3QpqxBfyMKaCX7pNrbTAxs4ShL/FMckSFkNxIbwJty4JP
0h5JYCfBf9LW1oC9jVnyQ5/LRbG1YsmBtATIti6EE0yppdW5CdiCTHAS0pUqbwL/8D4UnoYtCkNs
convAysph47+MimCPbAy9A+sf2nn7X1oP/g4JPHLgf15sKC9QW0V0OEAHiXZpNZMYNdv2vJ8+SZu
YKQ3xt0sE5MrSgHGnRQbThY497rHQHcn3sMPwF7HtScvXmfLsZg+fcI8mawxnKdxEOC658WNu2nK
p0OvIVIiFI9FX9WbP3bFjomFRkrrApLVFZruzG2Kv0zGetCxMYApVJnDPL5Vek+EBwxU1iqX7OTF
AX3RGsJE08akkSbRQQkmlwFGCa828UPOMTrJfKYkgiaA5Sw6iMOGo/YrYUq/ACl2A12EonzVBr4w
6FZzCZuKDUM0Sn+KI7spuAeIumyRUkx36GBnDMW7EwF6b8EgESqG5LUe8PX5dYUR+q+v96FOqz1L
/7ENCMqNtK42ZkZmSiZg4w7dLUt2JqbM9rww2tGKstv+TrGlkUc8VJG0fXDu0DasMqdp6n91uuak
q+m3bmHb9UtfBY4rgjLZMh8ajEhOgRfBj1n3Ky6afLAWhfWGAMzj//vPDZEkoUDu007r8VVjUuxk
Bou8eKy3VQxJwmmdxgZiHCvdEg1TQ123OSR6YVLx4YWCm2kr22g36gx3m/NBOnBZSTcZK+wxfkop
2AWdLT5Fia8l0qVt05LPXUlFP9+ZZUeBrSe6sqB8UeoFyWWr/lvNVdH6s5N9NqxTyYmHOsQDnVy1
P/IfUPCyxP1ee/RH2/q4rkk0ga0C+z8fMdxWtCE4JB4Ud+FAl8zr9nerT/Fd4QyXGo5T/qq+c+uw
Nr/et8AFQa8krfXA6pK6Sf1FP6zxyD8dpnb6/pwqJuFFGMm7KKynb5nIzsJP1G8Ld1unJcDoiQuZ
FYXX+mdz117l8eKwgABL6C3E1L6x2n1yR3hxUwHDin5NeTxrz/7IMO9l0H6B/PbCZfshlsB9lEx5
MMeDCaVV2bqdcuNlkGGiLNHDKw+hkC90qxKVZkd84SMsFG6enysWxhbB10wTQzKjRoh87akGKbaN
62KqBnBAsLPqmUc0JoGR5SKk6qhCkR+25wEc/PaDw2kaeEfVBJPxH/M1Dyk91j16KNtOAeHA/5pK
YZLFPPnRwgddJCx/5S4oieLURwoXdh38zWQ33RYt2Sv3RAvafHbU3h0nrWpTWH9x7qMHoWNc9lTO
2mqheFgCTIktlvkosV21GhGUrGkjok+y82WAWdw+We1rPNpISo+04eP4ArPzicRTCAix9uWZZgXD
0j5lKoPsPaKGVhnBddyaLWGmeAj5n2PAw5mPXFkx6M3d9M3ReRICq59slt+RDgsTK/AOoEczzpqF
feB4Rwz0XkghRe9Sp294cUg3S0hffWYL543u4SWcCXYqkgq/oIyRMNP8g1GGldoAAN6NXmIxJUU3
F4LSDCq9FAfKMXlle8fNQUI6i5smFvs1uYOYpjex2XQQ4NIg5jvQA7XxBI3eiPrZhCbibIJYjUgJ
PEw8/PckaU0EYF24Rj2Xwm+1mI2kdt2q096K9uALpZyce46x/3ojn5nAjAjFdWlIaFjYOi/y0vd5
qQGGgcBEdIGrsWuhCTrm/W4JiYw0Dk5xG+KtHlZmj7ItSRs+njExqKim2CkwO3SjAIpybysYK1KM
NvqDEvyF1YRPRA5tHSBt7HODZZiZArW0onGEAY8/urPuulbU2TaFqBOMsH72p1QAjRjC3Bi9x9AO
iiL2yLkt3XjMhCFKUy3ptoLOd41NsyOEgaTrDUxIzNamZq3hO+KdRB/BlrKlAXJIgKH6hbOIikd3
hXXYSGoaWG6Xqpkv65XyTu9QqzykIbQ0uGwT5gIY5k9keVtB5jmVBshzbp8ZgSe2GSviewNkl3Rn
5Wf+yUjUbML1SnBpY0Iby19soI+yBhvGzxjn8hCIgBvklY7ZkMO7McvoQwZ0eearYsCPNZMYC7gg
/tUFgJuc9tCdkyA8mAfVXiwWXQDfwc04U9fSrDXVg5H4++FW0K5rMePn8xth/04mWlhG06qKorGa
vOAHHSWXhrpGvufkpXEZHs+WTLeudgbsxiVGg+HkmdL+2snFxw62VpwA7xKopbIFQWQIQeB2Itzc
8i17PTmf8VcYYiJr8Q8R4pFNoiwRWDw4Vxs4znDfZQDSn4ouUqlVTdLHTBxfRn+kEDF7E8DGtZvE
QGtQRfz5y4FFdEwxpzzJNLoZLnI7MkNMEhSzFeqrDSF/mG2o08BOOgHJESG74+nRffNzp6rG0rwG
wDvrTwBIZRxsB9hB6EYcepidQpA7FsgUZIoJ04vWkCYZkgoGGtdP+NLTx0U9WItDHMC7fS9MBmB3
zUuLAqLP7AzTnZLQkutiP/14XN3MOLIqxzO9bvott8iirMkwmsYhsN3fghvUJvttwRVXWCNRCk5j
S+KoRdP7qMXqyQANvDn4PJy1qOXB0dZTASFsFcsaLfyGHbewHLrqlUWg9P8F6xr12Q2NGxHfPcCw
wQ5FTdNencGha8KuvX3C74pJK2E3v474IZjL+/4q6RYmil5bxFpULpZN8lofQFtMGN56UkDUSMwP
LRWzFD2Rh6kOChqmdhkC5IlliAlVwKto5py51hU54mQ7o1lv9z2ND3HqQAsMNhSfsV/7pcWm1HAC
c+xiEXMURzplKHhNEpsjISO6jtrhK7XzyrxaSHJeEhGSXJWfFYBCzN4rvNeL13qc2siyL3S/5Pbw
S4LGdv9TK92Rv+DG7V6ychM602I0VEsbs484JiWCzYX/1DJj2wDzr5KWHPZ1nTf+eJJE04yM5Z1e
vhcTd1SEMxPgG30Ec9mqFEigL3c+LBCjL+MEulwZnIEorkIRINzC0TMdm4u3P+Hp6TwjipHstKEm
WNTnf3PdiQ8QR9q6kkRa++XHkHKsvOnvgszkOHE0ZqfpdqkGXVtmie8dLCv8OiOJuXHPmksQUy3i
0GUV6UZUi6mGl7ulrHXX8db7UjQRg1ZmNquYV4zy1AHWWugFN//xJNy065Vq6DGMa41cIR/EDC+N
wW6WSgHAcenjigugueZ5rF2fbBtf/Q75m8Bf+xPJkly/R7rXhD3QdhmddU7qVm+eZzFw4qiWhLiM
oOY5Qix8sOI2fgM1uZO/rCDF2WxuYeQyu9q+rp7Yegd1q/V1zQOofh7U6m6SvRgoP1xWOm7NK8ws
I+2Oow8GAjUG+FukXPDGsMACGzI58tjuMip9C6wEtLvw5l/fhMfJVWRnEIOwYlJa5ZtBHbSC+54H
TLnJY675sPzwT1TCeqptf1yGxIKyNBGuSTafHxEx63EqNx3ZAgl2ybULPwDv1awpPy2iiUmji715
7eeg+ULC/+3bR/XSPiBPG8ZME9cnjaRXd04E1wfdpRBoSld37Zx0HpWTCNlZwYYAN3ThZ+lGk3oE
ngPziuXpngBeeuCOW2MUdwzspSksZ2XZKUmf+rvtQ2gF3S+3S1ny4gtlTPvV0tdah7ZDu1eAEFQQ
BDCjev6O1bVvCGsgBEM5G0106ec1SMbn6hzVWwz+SCMvX+4bPIlNtjcCGTwASveowpDHMQxfoZqN
GWUMly7D2VycIquBRGEIgt120poKwGdHUw7cPr+4cJUoPaE6FiSCI7YgkxpF6ew3VZR0SNDqt/0a
T3ExUbpx9d8YyJGw/Eck6kjRkDWhsx7DDuI2WS8YTQsYnhla98A7DFTrOmTXCg5FfKTtB4nCCNxV
nGSh+9SKu6W3CnmHAETVHL4vLtPWysCNVsS0O8m/Tba2taSuWLjwmdNcJnKgWt4l7yc0VBefPd8F
NvOEW+EQp0q6t99OHlwGPXXrXYMhvOgj7Jex9r2fwxIerkyeIPF7fuIFykZKA1xo84ZgF4dn0rCn
PT7w0o9Ws+bxBc5A46idyl4Yd1cTTZ0wihUQFG/lFnipDJTZYyEA9Mhz2EEKkLxN6Y+MrlIPUyz5
m9PtrjGkpE2G7X/MJq7pRLubJrBFrMn+LaWsuEkeN3POrwz1v9IYP51d8O9Y4s12+In4ytOL3WCw
V7ob3PQetGIHNQxWcH35B0FQIIPxTcXqxy69sq15o0P+91UuP+8/bkI0V4jmf2azS+EhjkWWuujE
fjEnP+6ikM281tm80JdEpDZkL/HIR2x/SDmIAMn1v5NpL0519c/VgqVwuWMe0Er8kS79qkBC7qhW
x5ZwWf8YQRMw/7D5KpIYt03kPYCroeR3RxFnfVWCWpIw9a6GjuSA0jeffCMlBZIz5xwCiTk6WFTj
1W4qWh9Up+sIFRl62zXHW9xYr/q7sgBMzyWatVj/E6xt0tVOMmASu6tRT20pixIg3LUY76kEDvVV
F+lkf9xEKf7WTDSlBqv8rXAMgRFY5M7M1E2UROVYJgHrIc4WoXTQq/rKEhjZElVeT7EBiU7gL5Q+
TM1PRWdteC8SZuz+K5tJF+MfAu2Bbese8lhJapUbtkZyGdFtO2NimGiWkZopCGqppEHVvHz3Ttgf
uEhE09ThfPsWXgm6W6IQL8DIcZW7xRwho/8JyEukAwEbweEXO7flyEx/ruZQY4AuYqR2b408XfVp
htxl8KhIUNITKZ2jHQshtGlgqZW2umbhCx6WNYNhOXH2ln1oqPn7CD46tjWAVt/5ojgq5bpaLlIH
hNM9Inq2A09KyojfOEZZBJojhpuZ//EOfc1/HTLxbgE/8vuFrgmMzRRTLLXwg36HJ9POeoLxTJu+
8Xc49U3Q4vI1vg/IsgTcFmz+iAPzXLp0DnxPu9BkQlYG9TFRBJnNj0oPwddnZxi9XKqvIxWKdTot
H7SS1dbvzV8okbeqp7ZAWmoKIagczgb6M+c7ubZCVKYUiRp70icMJ4Z3XPvhbdu0Lgn0Hlbn7RbH
6pPLwDCcIRzRijTcB1+L1wWM1Nui13yz+3jPD4I2PTzJqqx9ikP1MW2Ag7ohWaoEirs8ZSA9V5wX
Eg6w7B4vw7IT77xdyfN3PHqaOH/uhKgw/lx5ok5w70Hr3lr0fhJkHZSBtyscSZVBPzf3jAZHPSZC
BljmSq8fg4G4/9A3JpAcBaqaNCcjYHqRs3bsN+k+Ff3uzvMNnt8bcAE23jy9IjiWHnu3NFxBcJvq
/Lw5Lk17t3uEW3TKqcSN3F9bw11ET46KDlaqAsE3Iw3ez04NpR9yJ46MtUYdaHQN6o3iT7ejmR25
2P13++tddu6uLHXX9bFs84PwxrunXhYcGlGYMGhUXjbanY5HP304Ox/Lz6wlfzji7vFsLLgtQrkK
mjOWMDeXUeq7FKqpCw6f+ni4WK6jn7JxNFIFdZaMWdT11xZcc3Bye2jbg5V5U4zoqEystS4EJ6jx
WvnpU62P0M2EHfLm3k0Tk7IHib3j232Nx+uirL8FztvTIwWNVfK9xNxUo3bgsCeZdedyoIJH89Uh
AVTNHbHlID7BYbYY98hV/mKe89LBh3M3urKB8JP68kzN3tMrJcMiXDPmkvkYF7nZRbILVJ+irjW1
EejiBZltfeufnc6dUzaXztG02yLyuCUh+rhwMceLzkGdLmwMQNSOw0u+zZPubf97IpFABT+mPMnl
CaV/EhfTGcsF+rDTfHbot/bNBD3xj5CfQYq6OoEIswmxGYtCPlFMTn4+q/ae3hA+NGVaylejjZVU
XtTA31Fvzwkr/1cA96TeI9xhA8uv6t37AQIyujynzDKEVfRbx1xlxT8SUt8pinY2rhWtV3NlxbSi
HvJbvHaokkHn5VS47rzbv21x1lNMBYy4BgJbIx4rjMo6JoilLFtQX6SzX3RW0bcld3CGxATHfOKW
ESB9sEO+K0m4tV+475NIFpNGFbmsXba7q/VnUMp/rn3abTlwfcHmXTmSXq8zOgCJFiqmaDa9oXhi
GHIR2DSYB77Vkpib/1ap0JF/p4WhpLZYJNLQDaLL/QfDw75+CUHEDIA0XSjFonHhC4cQR2NJVCKG
Ihmy9c8R7ai2hTA1WHshqUTFD1bIilm6bIDqkGhVEvBeS7pcJzYI3ZSh4StKfKHE3fM+hzJ51wkV
ScMFBa174sh5i5RoZdvLpFeLI0NZ0BNyTsdSiqNjxk4YxEHdK9ba6CTRdTeUFNRpe7MyegDjwn4a
habAU04uOy3Fh9HIIcXJIVsEsa98B2w/Vh+cP3LqwPwGCpfKBn9MHhX0gi6kQJVR9SMGAYTRVelO
V6NW/F8mU5vWaCM9DjeDvG3MB6xvkj0uptXZMFiN7ZWP304fHIOAYIEgdDy+loe71sEwIPGvrRKH
okyzViu+hIrmEJiVUnmgFcQ+KyEu/ajgKc5SPIA31Z3VMA9ZD3ZLWaoM04uAqqCp9/xCAon78whQ
E1ZCwAlUfrPpvTJQ7z2X2BopyVjVlDaD0NXmWQ0RA8vMwhlzS646Qi+qXyGu+H3iQ9NgFOdH5JfX
+t7vto1RvWROW1UmC+i8cyya2cOW3JbBFHP6Faawcq/U8tNFt5pF+oH4QNY1+oOAlwyyoPUtb9Vf
i7qKdMj75ZMrOIG9huE/zOasRe0bAxTV8sVPOElHP3fVwlr/lbq6N0PaXptCW1fJY10jzBaVSO8v
//lAEqCV1ynV/4mvECn0mtFZS5ttK1AB1wbAx4xZDYy1HvOz4sUSlzsWrLJ9wuJnm4Vx9Rzua022
RSdCk7MFxkQla60q9HpGoHgc03TuN1FELGReUOpWy72WfY1Xz11KdNzSQePhYvBZc06O+4fhz/ne
zLdYvztu1OBQzAB2d07yvmgl3VGT1bZghEI+ecK34+LogIvLTdQKtAOUR7rZKN0NgUqnzn8YFPnK
RJvu7W9YUm9iaWt9NtkIzVzIPNQTIpk4RwPf66WnTR4qGXiccLB0K75iRADc/3W086tJ9VU0ck9d
OawA739qlXOK9nWxC3eLBQJRMp5ympvPade1pfBcyGRe/fEG98INnUgnhHlh7Gr8wIv2PUwyLjVu
bqruXhBibO/+TuW5mIV4L0G+oof9S4X6iyO0p9DWzRKmthW4+nBIn1Un2zxJHziMxEHlImqnNV5h
wOIM+mmf2lUfQK90H+/37oZpofatTlQoin5Pdlxf+Jyy174wUeHZzItEEBf3c8v/L0bSOfWqOdeC
PV1jaSNGF2dDPXmCf3qpnDOzclqjpjIyXtoHDntD2GVh8MJSTo/KyHomFniv0Lbrt97sTe8FM1io
e5Uk4AcG2wwwoIFhemDbWmSU0Moh0Bf+ghs23p5zCfz+WXGKJ15AUccjCfIY0gJq+Dz/zW+IaGHX
bUhRtZfzVJfvMCm92VZICGSz1ZnzuVVsvwUeJdPSqZWtAATiPVtSICDC5Ya8J4XBhAL36eX5bBsW
ACWD7OrT7w+aoxnEn91KI+CQ1+Ydu1qflAg9nr+gAu1T3Vb2F8vjmUzqB52HcwBggXHV1uUOBpk9
JITwdfCS7SkIuA2VbhdbE2Um87v/TcMeZG7uuNpQFEZrxQ0144z+JOtAw+9QY4C7OX7QnVouJKNb
ZO6f0IxKqSQpPguw+M2LOuo4x/DzFtS4cbAasxLYkYDmSsWzJ3otX/TVLYiA7eJ1NOIEVGYtqSPu
/FKKV82jWxsC2eZJ/H318j7RJteGFmuaZDNEuWZT8wI+hXgwuUf/pxcWJbpVZzOcBkbIlRZHiXK4
zBj0h3FGG7hfmmvZ5C/s4AMm3EQU137G9+mNAjYp6VkFGMbTdqvqfdIacbbqtFknCYlTHft5aWis
ywg5/rfhhqlqr8GHgiVO8THxDUFdawTl+g/HhmJzyfEEwo4aVN2cYfHLfnZQQWrepdc5gVFObRf7
Cr5pzeCBwX6tCuJe8UIS8RyU5eJXB7V4ZD89J/atBOarZu7nC6lXiorXYSYnQ+iutzHNVlp9OrYe
Cbi4sR2v4P99ltISkXBcI3813SBRTGOEg/q5bzFCW1VZdKcqWDWTZrbIr16wf7zRJb6xgpjlRZKV
m0BsCUWMh1ui0wboC930lMP1OIoJ6bUdMMwMOPJztjyhLf1BtM/At+c7dDtpKuv096cflx04bbbn
i/9y3g6YqJG5sX2EhrCSe1yCCzPuAfGbk1wpvJZvIwVkc7rE8G4DTyiPF7j0rbYUsvNLTZLINCyu
ZH7eXWnFuI5sBJoRr7qb4dNwewolPjMeKpuxTa1/TC9NhjKBmj/L4S36Hu4QSpf7dJ6F9eyHxQs1
6HTeRVVZ7hBM8oRlqlqsVGyIfU1arYM8Mx6LFQEY46I4koT+mIjbHjFtGzEFt7TRaewm3bZWeV63
6857cOugM46wocpIyiv5SWz5L5FbOTvbz5iAU5v/o6chx/l/ShIxYkztsqGuYSL/NQaq8NzhBOTB
VGGrKqdCdwgJCLCeZx5IkT5XJHlKZdugBnJrqrYiqGEjp2oab/qEb4hS5lCAc9heVjZETetpCD0p
/lGqu35vn1mI8pHVQWvZZKzaqJkZNLkTSbQ0e5uH2aYrRIq9cpbOc3Px/RrhetDRzdUloJIfrA02
je2muOoet226YBDytY0q8L8340j1QtFYgniIXBOMc2UA2wXEHqY924SJt/M8Hp1Jd4IeFIOq19JO
os4R0nX9Q92WWqptUR3aKkTBgCAru7+DXwK7/BB5qyQQAVMcSGgEkPtx4xdVc3Ubmn4M1VaEJe0f
2Xwnz5RLeHBDKPz0epFq3wbdAeHO0hOntuhnD0f8z5AaPmGqT8D153FJHu+TAokgEd6+TEoxLkAt
4iI0HEhY7Zj2bMo5KG0Bj9zymAxjn3yCwCVIyO56kdJTklAsaXzAHL4qKGn8wXPSEzH6bKSi/HMh
khqcRtSnElj3onIRZ0gX/FR8Splj29DcAV7blVL2LotSt1CRhiQQst52ycJaaI4kjuhMGH5Kys83
FiciU0FKwMV2+o/QimMH1XuG9mbDTxvYcsSKIzNAaFtm6ORex+rqTnv9fZCXvpn0ZunrWlnZHw3Z
uSlzxtcTCfX/wSUq7ps7CdWeyzbrsWXnR3qmtzlK7btSNkK+I1VbkY0yj/gCgrXR/m3WV3ZtjkQ2
1qc79ypyE6OknZpAPrf40CPyLVhh5Od781KQ4J58/TQM8133Se4zNdCOpTcJKbbOQd4SgWleGQQA
SmvIggSfnHw5rqOYGomxVUQLmvqGaj79rHJPlGckiQnHSqljPHidEjRMfTnJR7M3TAm2uDHkoi/L
kPmbR/GFOt5TBsdtMADUBvsj5aAyi/JKWkmiTLj38Voh/qO0m+XlhpPxfZex+mD6OuEBDYDSKpgG
2HFWc8PDa7p8PS9+S1ML6LEjQzXRSK+I4tINgc1D2ooxuCgqmCtICaFHlH2WUsxt+y9BCUm9PGWd
tRo8zu+atpazQsZVv77CuCtFnn+qU0iQyeqAF7b+SRHBjOjWWgRQ1s1lRDmQAU8SZXwkD1VkpfeW
0V1nMjTL1PhkCKC7jDaBheKr98geUtHeKHYn6G4LU+EEcq50sKTcNGcdlCJlKQzv1soD6yOb33ny
RY/Lue9w6jbH97GVNXEmrKYs22aClFuWV3jrm9LtKJonGH8tUUBFDIHgjMYnRfNJ4nIlulsQHWyk
2Tx1MMvlmlbn2uqnDQs7BypWt1swfRxvso71TzzBLm4QEbM3yTrepeVPpKyano7ychKuuyNiGGAc
m09z6ZMFZbCMosdJybTWNHwOkNiwsILlKdIJBnMmY/zJT3XNEgU3RvIwAcO1oeVsTMmbGzCK/VZW
emqBe/VvqbLK8+Pqz0DAlIKFTrw6TPIsCZQafHbT+mlpAs0vc7hNJ2+tuwTORo0Kr3po69uBlOrN
K+7qKHZJtP1OeoB1FmcxtfcnJKKxIQzBcmephS3BV31fy/K6nZJJspi37iy5usA/gbbfoBRENM1z
O2gZLPwgdvKY32rUKqPmZ+E68cGSHsMfPtZAMXSp+UPIyBGzwZ7X4GiJbWn5ho+OvAmUoykKziKC
2E0UtaSZ1b2r2Hf3jAb3tndkhJFZAg1vs1IfDVVI7db9GSRmmxb5sfxJtSwwZzsWT87yffgpcf1Y
tpy1nxnh+yazW1pWjKByndtSAPRg7uWbkCphVuolkgC/4XKEOVEWa/y0klXFPc1Kl3FyjXCCFyz/
i/8tyN/ScXM8s5c9+sCKqmS7mo60+NpIQFFLSWu32docv5pdOHqCohi3oSXVJOotg2KzCldL0y3C
PYzee2g40rnNCfMVz29D4Z4kbIH2h9S7ElT7s8DZcGxcDa4NSJJHvhVS5jT+buXb02t4kVTVFtvu
1hVNKUV03YZ0k7gXkOdjAB0v/czJraOAxipLsbTBe8VZIcgOu6COzwtc/GxBRhIZtkRyzxAn8TXH
JN7VgSfdMVOemNpAZql5EF7IKgsd8zcoBrp5/VJ8GRQeZGQT2jqfpnSHwnHmvIhRb8S6EIjQgrit
571FCZXUaYFM0p9E010Ri1ru4OeXGMcd+iskp6fZruDZ37V3OuZf8DifSGbUkDEAfitLCfzEjoF3
opA4gMNAQs6CBGHa+RTPxYh+CKB/KaSA/cgQ1UDy6b/m9lvQNzBbSaDorA7R6wBZ8bq7laVKNMSR
w77ZcoHscIAhAWsjCr1mfzDi5OwRY3G/RdgULKQy+ek3kl/qsZNOOdPkIn+AQBAOkAyG0O53bcIl
LkxCmBmwYwtr3jk6XJVMWJd0DPcnTW+JNXYpDAF5uumyMqs9rtQWmkNVoKGr6CZQgEKfQ9ICW+f1
RCzw7yEqxXqf/ZXgmDLwCEwAgugnWgtAgYHdwN+afFLWIzzd1juf58Vq5vQeFV3pjuV78FeKjpNg
lKTm/77K1k9JMkKxObao09r3a55vxKCbqenijYjz65BBkIdZd90cjuMymhxYK8nS5MnOvYt31IJ5
IKEDfmND2Bd62kCWejBfkPMsNz5v+xuY9Aw7fqMTqv2bXr6S3s4i7JONH1WRG1e2eJmf8CjH8ML1
0lvsR9KMfEAFVxDCDA1vZxNqpaW7geJ8nOJWRstqtAM8yZ/UMaqPth6WOAXEtkdzLiAhvwVXQy3O
IIbstVbIL9dzL4ALA20pOqdZBS4/lnsNq6HCjaqOqNrY0ZvYqDQ5jflj9zynFCCUwGkeEXml0K4j
a6vsqs5tDYkyNg2Nny7gwew8OwEv/ucNQXIiRVTdrsHwOsGrBxjTUNW3OS72fb4+ZPhDNceMGkGq
RQm0HR/JLpxDWkrbkoJXsywpTJvgDiv3+RYKLVQBKqT8uKm27r9GSPiPFeMv70SlmoRuhA3FrKxt
P7YbwuVF8akTMGpCcxavLwwhiQIXOq2X//tvOrfY805lyI7+E2grQSMOxonrZ5qLndz2MG0pu7li
iid/ar9Wjrgcrhod0EyIPlnKkjTVprIFAlhUG7w32GDTxbEOhMbOWsSXJXGJBwTIBRr72qtq9hqQ
EIF/9qqEPFJ686wtLUhSA9XSXHgnNnw8krC3w4OAWdBnKdPOIrSc3qD4gq76Rrwh2VEszW9L8zKy
WopPMamREoRdDthIq6uKzyIy0yIoXLl3KPtm4QbDH1EyE/thJ0T6cynurbZsF1w/C6pHZk5gGO90
iE80jTb34mKAvdfVpj8Sm+SbckuAWXeCKEhkZeUGEM6d6HiCmoLwr2eng2CMZTYP34cv4O+7DrHa
Wc+jExJ5tPJCl/u/NZh6hXOYiyAOwko5UQT/pvWYQNR76bBjsZUHfypPq7FsXNbA2DP9+ebSFngP
p/6pbZW6Yi6mxs8tCpS/VX7XbRI73CpLxnR+/n9ucBaaFB3XXbYRFUkC1lxJEMlWYBJg616S0jcI
h+N+9bAd2cbP+EVGeoXrF3qeHypkbnmc2cAubm4IoORB+kg90xUyNnxzO7JXb/P7LCshlOTgSJz6
9FmZnSQdAPql6/tVJE5i5+Do5H00UmtmP6AKJYf5sQBht2Cq0dhnfy7u8Bum0mekt36p/KE3RgUs
n+v6BVdQg08L/tSgeFfhDxLvFOUxfIzrWPztnMkrw32jblW4r58QiA+QFchVqsj2Y/5M4AEvWiYJ
uZFLkI/qI6PIGe3ar0QpMXfv+UD/l+5c97PKjWFTLtFc+E4YJJ7XaeQmcZP6BlRbPwWuXZblrNx9
Sd2mf68bVgUt+g9PamlmDtUx7ipaDkRf6zFCndGrtE+DUeRDHZ8/BzLtK/BRR4BJ+MG3WARbixNk
q5lJPcghh3cgp/PbIgzfOi1kzpUjxvlB3FmX5vqhuOjEYvE8osO4XsOiDAHUl1MapE+T4vH57VaK
YRW1xmu/gKlO5Sq32DALCDmLrHYGyPQcCKPJ+IG6/6rWPRc7B3l9rm+7mL4RHbhMrU89eXZdscqH
EuSAt+cxkUH8JC7pFvA/rG+7KL9VVG1BKYZdx9/quyaMkmSSnFz6kw4puJquJssicmP5UsMiVRIX
u8Q/8QlhEDzqcJLS8uVpYpS3GNe0i6cuXjLv77b/P/2SrPH9fuIqKQfQX293ezTFCZ4OQM3IqZKp
jyY/rmqlWsWxEI2xWMr8aqAvzPG9D/XX9furAEkl5c5asTH3UrzluvtB1TrgQGYFNgPjZsqFE5cz
vUuRSlWR5uSd/xOxxi9EEO6gNRqZmNXFyoycjULusdeKsFUWCXXiQvutAcXgHNQmIR8MZjIqVlGn
DvuCNouGDMjCItQSSMkoQlLLAxEAqudusD9Lw723LZkJmgHSfrLiC169tsZZiOQEys7K9W9adlDn
gmOe57HBgxtE0wEx8DO1mECTYDnwYMez1jjy5vbj0k8QgFW6ebtLPDjEImXUlE9Im7Mh6jysdkTv
9HdJcnrGA7IWAgaSBLEHwMitampJ6zWuirjFxhHkZ174+RDbvh7g+VCMkHuTSdNzr4CQRlScBf6i
Ols7QXx73zJaB/lOyR/tiYOn2xiloTMd9EgJeGMtfSG851FHlbJpEVQLEc+QqXl/QHmIYazpdSUM
R0lAfNylUNHJl+xiX5XKVZtzWD1g/5k8NgQvZMAKhvobS5InusLl087N0qXaSfp3EqlMauQkeEDT
Q7pMu5X6zbf9M4ip5a8KK4HuBZ/A1dmY4am/sWDRW3tiKpbIUuToG7wpS/0d1PwmBAgIKGDFAxv5
7R6WaNrgXrVRGm2bS6xK2uJN4KJTRZ+DgKwVGo8NB8UiCV8vsmqZkhyoTVBXQOQiWOiHxAL3jdEJ
/cjkaohe9vyUvCG3UauIHl/MemjX4wbFPLzU5d14Hkt7oJ1S2MQR+1dCL1vVf+jvC7h2AtGUO4sl
0iZJ6hp/lWe8FV7J6REG3fRg+P9EMY0o4oJvw/SktgaAew+dCOA4A7iN8PLmETGo0+CmdCWC4Ium
bdIK9lyV9urHDZ/EVPfJSTPFxMKnhtOBKyxqrpMX1eoOrHtQKKsSEuYqjKYBYWLlEhvh3S1suLGa
PHH7XtaZpO7SD7K6yaQyE0t8C14mBRK8o26aKMnhDNZ1sv3gLJW2vwbhtRs5miMBD8isnWFB2T+M
eve2ADAJgH/iTVBiCamMCjD5W2gnKWCrrxscJpvkbFyErDHO2wJuhMysXZIfQnpIApEAEj141v4s
oGvGUFuwG6I5kaj9qvzNp9C3QmN65Atsm75FTqbg4Dan+evlS5/3doQbMZTKOZrWIHHwVX/+JfP1
F9ZpW8Ms8jgzfVKrf/nBJ8XhCE4fwUWGz+5uoTFovBuO/UXWZSs3ccREcJ2mAGZPnOBPrhUkHwhX
aHkhsHyBoVtEezz+VAMpiy2c5b8EbLXLhnU9fnBRFYIcY7yTuN5+DTtsmlKnMuSwrKfji78agdrK
3x4Dfer1nB6KfGDclS+sjODpK8YRHfWWx7c55F2kqC6gTZ4T/JhnKwd99uNuV6AGarSId/U36xmI
f6YJ/ubSsOxv0kOvHM06/EzOiLfmGthn5vp3zP55CO7Q4Dk2aGt9v+jokTvmhlbXIGOzidpANuWn
22HA2mOIpQYldUaRPITuB3namA+nIV3j1yUjI9Nvn0rSHmEUG11uhLyPugYXEweI8UZrSFDdnZvt
IMalvtJXodyTqWXda3SfPr3b209fqvB/HB2ObFw6aD/2mwyzW48/Tqrb3/v7ZYeNutYhf3B/Bmr5
19YC5QALlgYD1ioMtf7PAuatwXJmItkXehuEnoQGfmZVnBP9m+LvyiXdF+kUe6w14Q5gzqcTEVPt
dAMAWfBmess61w3T9paJ+Q+H3CsQsFc9loWRuHgsi23GRmYvNce/zJUn8C+PY/Q/X7S/QW8rxRV8
0jZ1neF9fYYNBQKqd0wBCeoRJN2gJmdri24alChHSxhhaAPI45pNPOtBIW5/Abjm0eqGx4vhshOi
R0WU/1i2zURqYz76OI9xC2ol9csy6Eg42I8DjDWXqeTW9MojqMjhRacJ9Phmr/V/1y/4XdfCwMmQ
4yOT7fgoQk2OERJnBG8iSqDiVPcrY721kzTsHwMILy8r2h4PoV/dlkcX52CHHPF8YMhjhK2bAwve
eEQpMl9oO4eoZ2qIlsPtquVO+prdvh9qxzYXv1mQekRrgbLbWbN7kI75NxeY77r9hvsWTbuVkqk4
4lehtGK4TOWF5tlQAtrpbSBWHVOB7EC/7EaVe9X5hsdaAbG0lgvv3mRyxwE6i3Vn/H7/Upl6YKie
P8HjdtCf5zgmZT9mIANvWSAo4OlBIq7GhTBvU8cflR8eX2JAMUyjl9ToEWwLg+v+EE/tSUU8jEh8
zL12WpR5XbNFQ0axSj0E9CDZJrg+DF+x5PVQX6xyAdP1ln7myVnW2D2RDVtoCHv5ZGIHvj1JfZLu
5fsBSMHC2jrmmLr3Ylqm/9KKQ4deoIglPxPcL3SZYseEdyZIEhtNO//mPdo4+rvQBaWhInafrwTy
hDdGVC5oxsMpWdFJu1mqXt+e/aIZnZC68YrPAwbJoPijp7l0l70tpRQ7A9UmXw6AkWAEcLK/kn+s
lrDNJPpWup9tV00Rlgl92+q7zbZD0ZRTjlbtoFm3NrQ3tLcHv6XcgD3/V+BdKJipN3sQI/A3Gpli
xLUNR7+X/5403kMDeGhYeA6xgpZiicJkiPWvpuyqm/DJY1sRVgFZuJ+7t34lu6tumaZz2KaI6eWk
nEHyEL8fnzR8K+CyZqEU7X7nl5PBrJlQoG8RaUd+/+oK8K7GQthYVIE2jJoC0P6l+eyFcqFlK+TF
IOWiLYY+qZvu5M6nhUkWGsNYk4LzNBEMzGysLqWOil0ZHgQ1haI8utDdAixBQ4WTq6n3Lj5YDbNH
nmqFZCofU4jl4YDmmf4foLra7D9A/jEge2lLsp22VX9Oko+zMBmkBfE0mIXEbwYM2HW0ze53KjlZ
AC0kuUYelb+5R6oXfFR8a0u6t5btj1cffR9/h6dYZTy4qgWpa1ayJGdBjP7zjzNS0y1hVK8Hy1aN
LjZ5KbC7nJ++trfLCv08EHl/74Bdr64yZOth4i6ZgXMXvBr7n3jEwybRxNUViJFtaDCU9PXfUTkY
Bu/gY8MczAy2pE+rO4tJat56rs6QGH5k8lLzG1zcfJfX5WiCvLBv/1fLGjITzIQiUy+pkJWfg1Qn
Azgeiv8B90YKf9M1pwQyCWewUqzJnZFMMRws5Uoby3QLyG5oG6EiYxHNWxVbCsfsbaRtaYzkoOSX
T0xrQv9fduHLzbFyj4qQyPt5UZXs4ZzkvO3QLPvjkcjx3IkXpjJ97EcWydCqs0++YEXVnYmmEnME
s7U+5OTnKXEPFkvtbGWRjfR0KdOTPN447rG25NykNbCJEYhYY3W+M2VvMOwMF2tnrIAROFe2Am/s
pXmUr3y2XGSzyN2MMaY+8cn14hS4+Ruc2aMbHitbSolH0XTUe0Eckbhdg6hOReSMaGAcG9EuAIsN
IPh7j3bydmSbJYYzEEupM+MNtWXRzjoydjnFvHK02RaN8enx1sUFDI7fWEooN1KdrAzGBz1luYkN
NtDf39aiSFAwWAOBbpajhC1AoFo8P6ljXcR5TSGxOQ6kOvkYgJCXb3hD9qh/7DMfOHHOSKTqAsDO
PH85wbgnbtG1kPeZnU93Mkvzo8CA28KT9Iwzk0iKmv7yf/BQK2JRVTKKj4RPa7SZcAboVmq/2+Ju
MM2gC2qt3RMl+lMkq4ihQx3OEkx2PRRZnYEtl3Fq//eb1CC91tkqaAoV4wgOwGyfgwBXlJ1zJ+Vo
7h7FiqO8MeHQ3MQBCwYS5yCLkVhtiZXe7tqZOwp+7V5ichmKWvF4h73/FFrJKVcLKFWm/pqUcWmM
nXCqrJyeBNw1qarxs9j+/ktmMcvE89WDoAHMvWfM6VO8H5GsZkBvjH2pkOI+4i4UrhQdFZfeld2O
5qyJ6ui8E+gBAZEFNIwQHsokjFor+kQBUtgxrEDtWqlaJoXZ8t1OIyrfzU/3y+2kIUZ1tv6BF4E9
gZHRDTOtO4R35n0LytAZQkkR793x88zeXxqggPrQGdwbWKSqHIpQWJ6/+aip8mF2EYHZTtdNUKhd
SXACRkVV7X+2mlh3sM579v7UJqDe/5pQS3awicP2OyBKrYA92Gx9CqB0P1YuV8kZYaWHHE8d9huV
K8CjYDL07YjMM3M3n9Fy2W40jizicLZc8Je2e8Fcr9F3WrDwUCRHETGAbshbRV5maEEeUGgnLoa/
SXHsogu4TudjWOhqOnFtqaKWgFwp2mKBBqVXdeSuh/mF+kpSyEWPhzRAZlqUQ34yg/yqlon7b3EO
Z340OnfBxGeA86tFroOBDJ9I4pjvNuaE9EiJj9++yJh3N6wVuwYzbuOzhzmCE6tbzX9wCSOx7tZv
8C/qYO9hcuulSPD5NCD0K4Dfn+M+TCHTPMJqofJjpcn2Te/TYACuDGmBnk3jholWL2ryOsVjaZeT
jCk+x4m7muuI7VyxztH5iozvJNZe6unC8UuFdkasFJVLZlyrZeswcdBd6zMhHtc0wKkdapwiEKK/
PrR3wyjYJS8RaSYV7bONMKOSDpAdgIDmw5/276zGCeMMHImlxfQVhFQScRp4TlI018CWTvlLa4fi
SrVBKxqQyaqfjZ/0RQlIp3pAU4td2UOBUIuSM1O1eGRJ1DkhJyG7OzRdO+zP4fpDCqpKine4qzx1
+voBxpovQlk9fMSUNR+NvhzDssv/hcxdkMzhBn9gdw54Pxqf00ID5WNay5Ex79nmxvFpeJM0sZT2
gqHiwkb7/3zEwDV92OR34tDLrDjqkdbBFdLHBZAHHU9k1IobQ1bsl+XABXezpWk6cMM+67u8WW8K
SWGZhexkxKa+WGWXESa+nvldyuV3wI4Vddb2Rf6AO7kqU9HOs8FiZdZI7gHV+If39/3lUjYdm3Ow
9koWK6m67E58PYZKc46r/ufaeV9J4PnbknQuMGFiyAgAtDAB7N26uwble0CRlV9sN7obASBUrP8L
wzsroUhUOGX9FBneRRHltr9w/iXXxLP8czTZRunOw0BscJvVWwsKBy9gjVMs8tdH5tfQR0TUymEM
VPKAUI7HfiiyioK8sWL52DMYskAdFgNAXdklU4cmcZkt3+dqRvld2mAqMCC17UW4t4LkTCQZ/aup
Id6qhsDzBBlHW39b2Vnu7e3Boz4qwIc7jIkOgYJxGcXtpFQ25IUN6uOxYy1TUJ4L9w0Ly9syAa06
fpmQlJYVV/mbIOSCTKAO3jEPO13DAv4rcJyN8bjpExBz4nWepqU0jeuSiFPnBLtAcOSGTF8qbdfn
VPX60rmTdQNk5m0ZftKbrmiOsDFgiHnmtBVDDADA419PsxWNtPphjbsesb/q28nCTH1yq8feZs8o
odqtkKxLkmS3p50kl73n/Hrv5xcSxZ9itgvXH8ZuWLnBtSGhnuJTMqRizhq9bqJ4uskktt1hIXtj
cGgnX9wbwZERW3wrseA4N9oHw4Wb7+4RHWOtc23ngXStFjSiq6GFEBd70bl2OLedwT6nUWW5YpRH
ZzsQGNnN93MZNiygRSOD63u7tl56ObazBU8Ti/KijU3CZDM0VUglmYSDRF+ynJOJQd5BRrvriajs
wSwFpKsxXetfDgQ9MkmVqTSdpijwfDZEN/n6adm1xttxUt85noTw9LZ73T/oSY7oBL4NX8PpIA13
tWccmS1EYEF40wZVrIdapsikG6Fe+NXbfjP81hX9udM7MmrG3h7JYiqq6Exn1ZQFYjogbeNow4gc
r3QgcxMOnCuimqN1rWRZkxNBtaXDN2+cKZ6R+MPfOQNyNhzTlRkZJQ39aeNqAVKnm6ZKlhW1JPIx
FrUzCoXgOrnA1Zeod3vB3qh7Q5UP9L12YLqgRVZ6Wcv/cLSZSIjoE1JXY/4bO1kin6IOAAP/XN3E
qo+LEajXssfZx7Mn1vyy3EFyoRnx+MWao8FzKjrJZQVub7zvpz3Gpl7q+4JeQq8ywFD8AIfGN5rn
PiP3G/L3KONs7b8x4UgWhgZ4X/s6B+QKptNMqAPGDUcag5REUjFTpdixhT3tWWTN2QpzVCZePIah
Ams1Afxy7+KK68D68/zePYRG30QY/yBHiYBpSswcfMVLpXFgGYUIu2Zx4tvD/KWXtq/0+JJKOcL3
aRs5l7owMKrFxwIbrVz8dMhYmwv5EHj2VeRRUrGCxkA/kRW3FZqf5nMcAeWqI26WVS3rSlxcKHYl
iXbxAXAixUM2Y31RHu/SBiVwjENmExqLk6K8RCp94tWwaso+sI31QoiwmYkVvyYzNafzrjdft8nW
v5J4OZdAvD4abWFqaCod/4VSDQKgdtb/otVGjnAo43/QEdA09sZTxYJmLkejZoAvWPBRM1r6JoIN
xz0GxRw0lmSRNdWBwtaLlGLJuU+jYZch8+Tek/PEijqikuG8vSIFvo9ifwypcjlj8xx7rCycVDy1
fJwvDWjVX4k+1JtmyyNjBL9RRNZpczlh9B+F9hIQ3T2rtOURb8bx1Wl962kv27NU25yRVZsv2ayr
mrEHrKxwTT1VsVLYtGaTUiwcCiVkEz704x6PEQQUHsk+DeQDSGfzzmCvdQjm7rctMM7CPSRoZGsS
44pG5ORg3/oe1wRQSP2k7BC4IEE6UcvysmbK0nX9AISnZxs+ZOhRjVziKjVXtmiq0PEEnsQN6ScL
C0TT1BYHKM1u7Wjj/BwyyPwlXKkdMJNZkj7WTPS0IaXA8uwplQTz7gphpw4UF00CAMDiNPjVSyvt
SqR0St1jEmdAHE0G0mkbfYYA5xlUphkgoQ5HVJrLVUZzUoXcYH+CJaS5au4Gcu6O70Q3uvJKEcSn
zlrnX4lItMYUqwb7lQNEtH4ekyvO+grhSsNYYljCpIBYyWcwGT4K67LQ3uW9B1XP4bXFW45CZE02
qFKkU+bNuWEwkOmRVCbB/ncAAsZP2+dZVdinwt56b9JmA9pLolxjgJYFuvTQ7SAFwQiGL+J2ifH0
Fl2/BU9Mdm9d1Bpoiq7Gb9D5C40f1K4xAOaNTDicrMJcXCnfRbb82cVHPLEXv+r1wXEMgmXuppEt
Y6+164H4DNh5ZzFXT1E5Tto2GUmKl0qwXJAVjYxhzENTO48ilgg3iQvnPL6BPH/k4Wc5mQ0sOoBa
lAVnKUKln9bcbBwOuVQes+PhswVeGOZUKv6R1JBiUmhRZjwERGzeKdgcLnhU45sYG3P3M7dDiMq+
CBDYvu8b/IaAXBCHyxnHAXTrWVql6IyixrChPbI6ecQmDAR/9fprjajnUTDXcG1WVr7oydeNFMGA
9lBS9FKEug228ozUKjpWwiwMBENTisib/DrxVXwi9ThKndQ6Uy9wavPPUaWzK5wHfMX+tR7RDUbP
eNjbPZy7AxGSkH3OPGYUVlX6DHJYYbBwjHlg38sEqDAc1lKs5fsPXMRPRoCrkv6yW9AKzQv0WJDn
Xqfp2vb2ucy7w54YywBgCxttafAI9JGsqexKLeFq5C2oxQDwd8c8diWE/SDK3ZomrS0yejycbhJP
o1QHU/Fz9P04al0hTBpTIoj8KSIg9nG2428cYwNKT7FvbfdArVNC83c0B4nFcz7R5Kk/vTRdYzse
+8jRteCbvVBTMAshQehfuC8rGUoFCc0ueeu1pICbgGq1LyrGcyniihkDA86bg/Hr5T5UTaNnDZUY
2fgsY+mPJwoaPTq6V2SQVhMEhL0IVB+ZtkHGL2GMoWHszvihoMxeO4e0yaD8Ffz7LZyOtm+bW39u
oYuey5Q8bpF1DSJYnRtSjY/N4XZ5QuoI6wZbGn/8QdV7Xp3Hd3i6QYhFNmCbGuf6v2ZPx144oIX5
1bwb4ZYVx/ChyfV4q9sbbtD1G89Ov/FtIIw6KXz17o9e2yJUimm7L13/6JIlQJTrEPwYH5n/b6Zd
CBu5yc9eSJljYiESH6FrbklNZ5wvX9kvJZQBzQe/J4SaQZSvRsTapnY3GZzvjIEO5VQ5/jLDl+4C
81JJXK/SNHuO3FOtGO+EsEZpxXz+PW2p5w6x/1frq1wUE5nVKB7LxBQwnGOWsXgq2Ry1YC1yZjuM
tDZNJI1y+JgvZgButltMfiAUNhe4HHbNGHBDe04q8Btq6lvub7ldYJasegdWHZ+/S8wWZwzaz7Ie
C23akC2muGghFcZYy7p44hZ+S7HOZ0pqUzW7boqMlGI00l3sBqf7HgVh7G6SQX9z17ZyQ1jl8X1n
mx6pm+42zRmhvJ3HiVGJSoy8eXqtjBcNgztAcMySAwb8G/EAOl1QjkzFN5/EgunxVOta/oFqgiIH
pkF6U5DGu9wC2S9bz9aJfwS4hj2HYwcydbt8zE+2zEzDcJ0VLdUhD+ztLqRDDGECxj7OZZjyXKMV
+qgNFot+69TspEdf8XenPNVerd7E5sSyU4IYjE5rNNo1IsZoxor6TqJ+doWz1qQCGDM29jPDn8gd
tLaRQSNVMbiewUzJNk7792GodaGlQnJ4AdGW3HKyQqoqagks0NmjWJJpdCkz8Oy8oHhjl8iFoeym
YfTBqdC76dLtDJ2aN6e11i3SfKeQTEmA+o4mLcTGN8KAFhqj44/TpILS5FIK6kl/Z4SPRCO74lVu
h5xGXAx+4a8EEtbaqs5qr/YrTwesQmHcT6n5VTI/5keM02TWXlFugG2+XegrLGZVK0xIPm5qvGbo
GXkz9zi0zEZpSjTTlWqjIV7YgiW0SbH+WaCRLG4jaylbPY1yYOQYgHJywmeKw4O6fbAtqUb4ReW8
ruYoy7Yj/RBkX6wqdYrreMWkkGyaXdb5aPQInCGjWULbUBsZXFQQIBiuia7EFXnq2SzmR7UzltKQ
IRr9lXW6i0GDJOb3FIhJ4Lh32GLu6RQi45W+a/JZvOhJ5bwkdToo+Q8FDh94mdkCbWw/axYAARgS
dEhwquTKaX94mMDSt+bfG3pS+9dBs4fvb2UERsWLWZKB12116G8a/joY7uBcki5qIcsGDLxczzi0
uydt0F2FWafK6NuWWtH6iwe+klLXnUu9uB1GDemjCSmtg1oCkdiebf6OKI1n/fPimiVn8wbjQzRr
MnPT1aGyOeUltV6h1CzQ7PYzjRTuT3dHzX3h4Ad2ZpQlCheKBO/ggM0RkYIXZCsJxUBQtIDukr8g
UdEgyFoUGJ90y2BTHZ8sYVxHRnx+qSg+TJD4RhTUa8bbLIVjf5FQ/UYLyqOI3crye2TdX4BpHhfr
cwnnFk3m/DsQZkt7iTc+Ggb364HCW9VbDRaE0dNtIKHuT+o92I1TNJ/4Y7yd6+vAof2C2lCI49Ct
L9gSenkaeCYLM32vQMelJFh2oxLnmZ8z1jqWILU/EyHVkUJtSHQp7lyjbOG9CRvshNSLK9Pn3HAN
JGJxGddEalc1aPKWHA85hBZhp0oRdX7Ds8N5HsryEoUNX8WIP0p4JXjrfiYDpIUkbays58Znxc5x
lDFlkS33PQTqcZCGpOQa1sprKQrMEWs08PXdtMSy7I7NQYhEnk0xakPRpGGm+uiadyYbOQyIdlCu
ZVONVX9R8KbRZn8niXHYHmiWoAEaZwO4zB+8v1fHfgiVpfUxzJyjWnlT28jQfpslKOyuZX0g0ZlR
FF3pF9audoWHJ0/igJ9WVpI27PWzAz3JK0Q6uXbSLfQ/K/8+kbYgjE9XLbBsVB297Hwiyg4Y8Sbj
z1i2DVhvX4UdvO6z6fA4nE/QfWy2/qNYOzX0uJlsp2wxMC3CRQGZf7ms6tXVaTPKlwKS9aG0Bizo
s3wkKp0uI7xFKxzVwrSYNW0Jt96CjDIDvcVCfAl6gzrmAchIzMrOhBANCFuo1vUtTSBjp4rCgE/U
pCojMDFaHPfgRRvcGg3oCVwe7tX+4iDr3Jpo99EyePLQ6a+MiW/0SAO6Ht6kKlZf/4+6qvTPt9FX
DCfSD54VVofm4PBGvgfesAm2MBMLE1idAAE1wMqWZMRtXkcWBY9kI3UeKqCBg8fJwfQtuHJ+gbVh
7FZ7+7twCmv+Jfe90qAgtmRHnAixxY1+3wHCgQGMd1vO7D/Ls81oz0mNnmA43tXsiWJkGGR+xB6m
2SygbGWap6ai1niBfPmdtxhiW2vUnYfg18bmzrKCwcEPCQyuM2mSCQN+Q9TcyqksGOMPfHB3dGZM
YNoCsbHqPVbH1fqfM7WEvcg0DnIx1f5Qi411GFrjmm0kEW7gQI9gOAv7ptNDXz8QG8flauWYXErP
6Wx0Xq8br7ZBgLgkPdK6Dk9rct+G5im4HmuFD4uihJ0OpwWhgI2kp4MACgzLTI8fu+B2dgghD/tR
Bbfek9A5IAVKida/wQ5k8Tt0oWtqEvXJp49aFyNFvHl45PAjukdNGaMUatAndMa71T8kwA0wTP3U
CAjV/MCGj5XH7ElSGFuQD+Iryq9R6eK8uK+B4i5wyqAJZvPoSw5hR5CbINefa3JwxvNe4/C43QlA
msoYm8T6znEiOboucRtZAciEUdS1GodrOhWJ3JYZmbjEdFpwOFzwP1usskto/lInVQxUuHspErrx
e6AIVQdHey12FMCtz9hHuoOoDOJpgMRgsj9UGR7Jto0M5Q5ASFN2RIzcq12s/dYMoi94gmEtFdna
AC3eewPvuqAQuozblxxi93VJP7P8KN10Zv0LAqIwykAperYnJp5pL+nVDXTgRKizUMKPm65U5Ypt
YH5bYlvApWNqnuy96kyq9yr1jc51GmY9InhNmtppFxbbVh1KdwKsBby9kVJYfgRUo5b3rAYRqc58
CzOWBd+q4n3/xkZXVRAHin96PHr+NI/Ndgn+kBTjEE1Y1qI0Ae9StqI+6luM302PzGgCgE/mYeZh
sqo2gE/AglBkKskCdYLXNrQFZJ1+eS3svmma6TkpFlzu1mnCVD6zGawJq2Q8erkQc5gShB7NtTIj
dk7pJPcjlNoNtZAnYcMJeKoHcYrPB/F0HneoiKqnWaQ9WGOLgaSvdgyvVMz6FHdB4RB0GWm+c4/z
NInig3Q7Dcx77l0gh3J1N4mdnqyFaJ7mcN0IpTkTX/a7J7byNpQSQ5gANcxbMzCj5+TpZDh/PRTz
2/HLA/FzwLA/eXTIf22wmknBdwOyWbCicovY2zARB3vKjshOz72q5CMeeRQeACrgdslfZLhScvLs
OzKRLzUUqSidJAkxeTu7ntR29ETl3Kk3WV3xzZsKT+z4bb6LfWjEDuaNu4BjfGRFPMlvGNJSaIq8
yTfSzTh+vQYmyruBL8bKfDzftKjrflT16JmWx1dhxGcHosdcyfohTVCYUkebXiuN8x3EOFnd9HjC
JuiAjNfzPXuvB8Oc8mGdE1Ke9TE3jK1z0bpnVvYrU3pgPt0DHMS36MZ43n+OPq9nZJmVTfdiT8Hz
Ubr6IORyVzIJYr14LZscjXfA70H9+dG1B3SJUagO8RCJ+J/imgp3EmDyZBL3n8XQgsL1hdiob2sD
oaSJyYSZ6R01nIWduBaN0PEg+xoznf/rNVQ5pRAAjpKPJxZNg3wQHwGqp7JNKUW+Eu4aLAZzk9Mx
rK/5R2VRDHw0trRiNO7xFhc4doezxxlgY2Pa579AwY7hGUn39ov5qQ7LDKfyU2q/XP5pcfQdh+ms
UeDttzh1Bb+Rd/s3XfzOnc6hLzt3QlasTN8pfjGjlfKB6GeP9La+y61JGsL/UeXoIJP51SijIQAe
T7cBzFJscjvIkDFaxp22R4JCstS4WQp7wNJxvyLRumej+Y8eqsr4C9XfocWfWmfXrH08YkgI9J8l
/99cfC1kLPK5ukuqspfK4tX3IKlW4dsAJRzNE+KF8L1YhJqrX455uH0UldXOk6sfAcDz7+/VvRDE
US4H2Qbg2D6ys0AiKJBQQahhVFAVfYUnTVCi7bheRGBEx4CIN+heALx6l+4z1GY0U9Bo0Sr4CA23
VoRG1D28dUS3EofrEAU2bHGyIftQFaUEEf08M1HhZ6bCNrl7MpYLer3m1loFV3fEAv3/+omeWWwA
zRhuIsR1dIvCF6BVSsKXwrx8A58QRuBU+OdnNZ+d4VX3WAWXXPc3nMU5svTwKpDjfnIc7VEkwcN9
vL73ydvT0A9VG0ph4oO59mqolcGBpXLybP0GgGQxn9HsWQU02OPQQgO/4Y8BVUPs56+4Sh+qORBZ
Vw8J/A0mCZpgeaq9l2/FcIEUmyuWtQiq78WR4DWE60UAJo8KfAlrE07+J0ddcy4gkw3Fhtz5Te0W
us4Xx8BAbl6SX9RmyOPiypN8Y+INWoayad/rx38MkmT7LpreIAUoBLqDhcxQEnn1+6fb8QjfB5ny
pbGcBrHghzfF6CBZbnujaJXbIhKCnnk2jgNTaCKssaTU44NXp0DQb1BMBRUPn24D3XA90FpMNHrQ
MrIKbDbiv2cJXEVP+c8rkkf5zg178RoMETfEp5+z8/jobl9qFt5yxjVl3uACkC6+L+L6MbKi/IVS
c6dQrn/rAN2LAOyY8uWvXYtr869lkX8QOlALR/GE0hlJPDbnAjhNpiipZgtK57ca+NC/x5m0Sr8A
jP/iE6hbfTsHAOakkBrvghZLK5jmvhXs/FCTS1jP2xFg+z3B/zEbKs7DcqZd+fQw4XrnrAdAeKr0
HcWm9cBngVXbMS2h4vmR8aW9b1jujcsoAjOh60WnZkeXMUlD5NQf8g9pn+kdvfwdTpwNCVDTfZLU
5Cs3MiS5WDTsKGzXz8/3TcCXIkUEB6GYlrZn7sTBCzPrTbm0a3snNnbObxFrA+Ej+yt2WiDKfeLp
ipUJXVBfaH0ftM+SMV9WJk8VGQ9WHK3CaSj7NRJ3q5qeJ7ErNPQDxQKqLCx4g3Hl7K/1hGSotRTt
eqsPB3Ozs54E+lmbAuEQd645vbpjhFi2D8SMoZRDe9RtoZUurjuDGe/WxRsMXzQidGBUQBg5BAxy
k5ZTT2oAo6VLSrNYafkBnpguGNn1Axlq46bgxNU0pv/XE3JrFKp+uZnl2ZB1B4udsL6ZUtrgPwXs
drNyRvsZKuudhlid4/ztk45xQz4sdeFgYJKZFwGllBENi+HiGtPfO3Q7BHQcwd+ZUvKEdaPbQ6Ri
6r9m8pVKVVM0kC+/Pu1I+E+vP3fPFdhG6h4h3Id47Y2RnydKIvVPipBHeW47hjXEIGxYAxvibFnZ
qbCPS5A6MED3K1F8oZoaAfVN/KUKcRTWeHfi9U991GW0xESntfc3YUsVTqYG4VCnX1EU8qdzSvm0
skbP0UGAPEx0111i4RLycDyzqc4kqQ/x5VQ0x5OYZhQaXiFuBGfu2JeMnvoGhTS6HgAi4+nS1H8l
4Iz0yBWwRU/GNrUKEkNr+nsCrY6r4Opi0LRnfP5G786q++e7m9eF+grX9SyCakPOx6QiLknW4h40
ka+u7OdXME3947quToIOyUhEzQId8IeWFr2O9TMX0QLewboyjHzVqoa5hz4brKU0csn7daUAkj40
U0U9mY3HiNaGN4gBf6tVmuqsIJzStiO9zH9In+sKbqmAQVeINSroW5JuTlcH96SQluZiL0E8ng/1
jEL5kJHeQex4D0a4Lq3tfRM/EQsydSQL+JhepbIkJCjuELhVYNU9qoHKYN4xmSsebUnryX9wbNqc
p+Xafp2tjxMaAxmvrcqBSn8WQ+jbdpcEWZIfJkDdpVhyAXnRofCyHVtrPQIeO0h8TZfbo91flc7X
LLOqrdkmUglQZh+vwEhwllgJPA2eL/4QpnU6cwQpfyBpmXWzOl2oL+dgp9b2lDj6hSbybaQWPliN
vo8VOa1H95NnNotphQ33WyH2yYi/cF27Yts6OzCflborKQ+sKcl7gmREcwVbG3bQvwfg2D7SW+hw
+x9AIKVffDG7MUY3isjJnEnkYa++F9oCl9YSnGzC0+ltQNEFPso62UGijLaslzfDPfkM0diyb3K9
KGaBVBZy0Y34BAtP1ZEQm5gCryGL4ULoT97lOxELDwx/L8BdT0cq+eGWjCC3B0hi8H3C84PqKDDA
repi/cQT/H3E6SKkR/aL29RQc6XeNfTRcz9MdEfTrfOOKBD5cdXewaH/JPVx+/pU+leluxN1stRO
OJOR5ui2lwVkKacN1jyKuTJ53bu4JH5YiTrpCpAfjQd2ssaLR4Yz5V2OghCkAYEjZQo43AIUOz/S
Dx16BrP03AiKqHgENNfgrOxcwtg1Ga4XpzFz2C+q4Ep0SgWKFBkjJ6F+LH5IhwytTGDtETcpr09x
1UjrpbIqELhb9Rg6d+uO2Uyf/QZdS0d9pvYYzsWkL+B9whHWmR1corFTQuHLQmfX1AyJcxxgBb1z
ivTaNM3ar45jmQGrRmIavh2lKbjDk4Dxu+1FnUVewSj6pyXImTeIVpzsgsA3/RY1KOUNwGhY8Jiu
tSYkeGl1eY2uOV+lWGdnE7vihgmZHjE5zSClXwUREms6Ny8tZfAZRK9NGfgUnWQOYWQAo8lkjEnz
6wZ6EGu4f9l0CSyNPOTsNZhp9d/mVBTzmQeYzvzaSdjTa7Ga6sBgeJKv6mkInEIlUkNTulXVBjPl
3ZFORWaDTfsqb+FkCkWGK39KwMU2voICmrZggZG+JEe7Ed4wTV471LwmDu9rCXmyl5gYI8jPJVwZ
/dEOJyvwIPQMiX4REtmKUj2dp+cPM3AJGmlN6En2jNtgCKJDn4Oby2MjQ24QkwTM1CCfKupkJKIX
mXKuJ7XFloDcrITpbyuv+mUWtVRyBaKaJ+a4N97WYwJayf9MUTQan/fVrKZtQQjxj3WoT+k+GFbF
lxU9Qbm/CeTAcvYsHGlpe9E4hkGhHWfV34hjO+b+WVIm20zrzSz0gmCWiDseDLs2L70chL8QGrUi
cRT9HMSnV73PKlZQgi/QeF2tPAewStkKImcteFlTpEb3jK4qD9W5fxJTYSZjDzkbcWCFU0PqFg/6
xkM4uIC95MTTQhUGSh3HeNwZYDf/XIEjkJ7DtpbMcQWlmzkaDz58qXOA//gAUODas8Jy9pqWm+DU
A6arjWg/eVkcIgGpsKI5jq7TE4z7aMZnk8Q68ik/AaaC3x0w/KCPLE1HQZRXoEJGCVkaaqs8mier
ybsBhpmF8geDzTaUNyrTvKu/jUCQSHaSyB9+rGCRTZWVHW1knj0HJ+W405MDsrNWaOKTj782EoXn
+1zK8A7dT2tTZjRMdMXC45+w0mDfI7Hw1GTq5RkZXaShCBsx2BsYX0CUkuUHHNb19/Dr2neZ8DUy
veDbh/1rrG5AWVfWRKNFbpMJfpDSkoIkAub5QFphuGrm1KTkH/521aqGQNmuf2+UymoHNByGMnqq
CtAcO9/ppJ2pRf8s4Z5/Uy3QuI642A1a6lsCXtMy28LentJgcitjKoIM3J8Y8279CTWzma68icPP
pPqYfawDOVqJ7pj0qlAofHXy4zM5KbdtNDncXP2Yj5BrrBEW6jVq5AUmAKVUxDMJUhgz0C5CiSnG
wwEYcD+nOfOhNie7mbaXnjCvP4wnKiupxXx+SuIWFF7WAxftZoetrzV+Du4h45KyNUJeaJsd1MhW
uWiSAk4l4t+MU83HY57MBDjTHm1w42QoENCsfRCa0X9GjbENeHwbCAW3Iopxe6MkEv7pe4gmjnn/
AgpkazRvW/QQ9i6NEqLa6NCndIFvrnzpz2ILdIw6HhNQDevxdtfyysGzaL3tHUBybh8zg5wXIZMT
R4it7jzeievT3YeIsu2dkx1kblBP2qz0SmvTpdvP9a0/g6dIxfCc/4q7LR+L39Nh68qd9s0a+JC7
1jzXFOoQGUbrDRLz9FqhQv5hchg5vYC8rf5J7pKKiR61sH6rlNcZJ1vERAkZGC8p8BxDOMo/9dCO
mpP5J897WPofQ9rIEWPk8L0oO3SlLETlqQ5kuQUUAfW22NURIb0KIxAloH8RNweX7hgRQRHBBNVi
9yUbPQnGYha3WMnVrKgPMliLIcyR4HzwnKIrq9bxnioYlIjbkvRKJSD5CX2UsxqMDCMm0J6gT6Hn
3W7Sedy56aZOQYVzffKxNCniAaTCOp+MDt4k4Tm+1W3x9lWH3rwQdFOS0oCwqQ+LRCrT8oVkpNa2
By2VfgRaRRJSf/Q33ohgnmMf+/j/UGJcEjp1KEQ2b3x3jZBqWQhhc15UpA3PSwghzOyEP2lGVGEO
TeoxHJ9aasmvCcNesNxqUiX5FyNjsj3DN1oi/GjDrv7AIo58lER6ivlhndGF5mydZiugwxfmPrF1
aly5vqfzdxzayTIqsUuccNF5nIr5KFh5sqbYGIrtQlEtKR1V/FRUWJLBHeH/0cscpiOW4YAHQFKA
PKIzo1Est9WHdY+q7ZC+K0/0SRNj7WWGmIAy7waLLzFpVkYoujq43kAfMYqN3fvnsBB6k5dtK+IF
lYMZQ9orfSPXFeJGLoCb7kgeEzU0WCbcKVjbs52yeDkV8ubGItBypJq0N1geirF771Uni0Q/sEih
e1Ep3DuzExCsW1c1TpzTMXIa+bCuDeMEGBwRG/BphxtfOlkMA19z0uWeqk3nzaJqloI8hJ3BxIcG
135LhgmCQA3DzK/bV/ycKmXj3fXYKsWwRmykBSDh2bWrln+gAB3vTp3cXNDCxNPDPfgWBvBt6DNc
33QaMI89nb/MGKf3CDAMoi6ya1JzO1LtRJ3HdS1YJ1X3+Uw748m5Wq4cJ9nlRRWOI3YdAaKIJtWM
rijBpI9HYuORLqB2NM0gmoO4kceFgrvPLERVKB5nx65MTAFNz9fUHRp20c5DUIXe4/dGPBX3WHns
/D8GMhnMP8A+Yjk/Gbyi+252f3nxv5/NvrbJtvcsj8TnxVyB9Hq9fUFRGGRDasT1F08Mzerl6qkO
PqtBPRT7AM4ohbhryPX9An8AFFgz27hhFGPrsA3yUBhKdU8PDF9drmlfpm587AaMoulcG62/T5LU
+/RKeBwojJuZfr4xXxNE3OszH1rSGKH18BeEdqakENkn+OsHSDTd6pD5hmZZemWnE+/t+zZrUfKs
Z0JC83hnMZsgaw8aOSon0Owx1fUX0Z3VXDfN6XPadkWVNsLD8/rKqONBUW4GvVvPonVUrbyGt+U5
3s5/rpGE0N255B3cRqQRxNaGTiusT3xnBHj6Gna7DnU8SlD9Ss7ncWvlYrhxHZSD7KBR++eWMUMM
G3WVusinD+BGE8uu4koTNsh9+WODTWjU1QnF1lP8xZVBlgIDLIYG48xJ9cjUSVROHuxrXP0COK87
5Y4gWnt7o6NnaHyypHSTIYYHZiDskDtDy3r124LHqITFhMXD3OVvwF8dVukB/EA5kYBqFOvROgr4
SLJvFOpFgJhLZhQ+7wGClbM03s351fjjD+y4OQ2qbbvIMfRZkss8Ir03xtlNX658MftPdq+G7a3d
uHmCJ6m+hltkGiqa5/hJY9NPi9ydTB5n+X1BcESq8bE7UHgiJZHHS7gbH93eI5C98bvPbfp/FMAZ
dz4rhK5G5IlNtaa6kvavJ2IHa1a/THX/PXH4nCwOA4yb8S3QIw0/+ZJVaW+fU9+tUT1NmQsUyLPG
RhQzO+hByjd6nTfefGW9G3yWO0LmsV2yTuxE6CsH2Y0SfZsDbmRajoEpC+Nh/rmpGOEoFME0LXk3
UNoEJSbtPzwOucUVN+qITrztLt7Ejt0hn/vJQacgva4pCOOInz6Ay/X91soSK7ZVID0iOBMLzU7e
f4XxtT+MnNCedl+GntMNSaPVHKUwJKxykXa/g7XTlL+NsUDqR/722qys6nAlVv+31ne49ZOhaa2Q
z2CiGAPqfKgGiLTaiZxT9pdC+xDkcz5sWrkKTnpwZskfCdc5qHiw9lJwEwA/w5+ABXUCh87KgZwW
NkDE0an8vsWeMbyW/4WvodFzHYQ1EQ6MjCWAZI1vYfJB1zHXIV+7/SxQ3bvy86fO02x2xNWMiZ87
1MnActwhasVuu2eKGBfXGRnoMnp/7aGiuoXbmj/GIeuEC9mhGye7/IExhcOObIc8CTkp7plvIppu
KcptoYSb0pJe4hC/HdmUJVnA0NZe5lSQ1g6U9PufRW2MR6Rfd9zzgQUBacqFOdy4FIHP/9iYgNBL
YjEbqBtlG8sPa9n4aGCGhCbq4Qqe5KeMhoiKV99fIJfnGBbKViHVEnZhubAmPDIKJB4wZeKGWxYU
pUM4PVUQfdW+HPg/QcxKV5XOfLleM1EM0wJlEW3IBnwLeVkeuernVlS2bsY5qgpGJ/gKRbJMaO4c
pr/10erKOCBKHkSmUV2UUQSdnvb9DJ9b6apjH9xUBEYjo4y9AP6GOF0O9f24znxetQm/UXG4Ks5J
Aa8G2dIzNuQs8VFy0ldMLaN8zA3ugOqEUEZeKaLzNdmGm8/Wwfs09XB8OE7snQmwcTvhNdgVhbKz
T/+DfMIlGzwdDcwLsf6XPrlPn4JTdfb+p5qp+phGBp4MdlyxEZc7xjP1u4A113PA6svwmfULfsAV
8Rhcol/E2yzfm/DYG31IXoHgPFWQiuo761PdQi+fCT9uUMY1dSd7lUA36Fn+vVQyJGu3KfuDCOzN
L4EVGvVv9wOHXPkMnBBJpWLxFxnXLrIa0Sa2vHiazC16/zu9US8YwdJ/ZPcIXoDyaBVNUFexVY/X
H6bfmQJy/UXczECKub9QFFu7KVgtWmqyYd+o/jrNWGZAmPL+QKtwUHFaJNvWIU2iHWgoV9LONvpI
rntQp/mcC1fJoiI9NrSCgpV3pc12JVuIWOnuvh+I0gWIJzkJ3g/Lgd3dG0isjf9GGbCicqoxU5qd
lW97JS+n2TZo+RnUsykMmrcdKiXEOCe4HY0UaFyFJ8FyCvvCmNdAS9suF0NtbkAf+lg4e83qMtxL
QDKBiOUt8ZbASoCCv9+RqfqfPNZ7KtF3yKLHgDiFkFAWveVwXxfg5dQKOXZtuwRrbcsKPe/fj928
FzEDuyoVlg465dH69y62+02ATr9Nt4i8QkB9XpqabQ6SlB/HGUj1ccB87biXggYIvnAGpzmhRMfQ
6+IgYgCmYeFMYFDPSUrWnTYcGKPPdTsVEOPkfHOK/TKgPyq9HdNQl7QsADo+7wYZuIFAWGeU3swj
IsknxZUPVstlb3uzKvP5xl7PYEen8eM60DW9NTuYh4JPPx5SHjfDHQylkCp7mMsMsYnsSBbLA88S
mTi60g+x+nZCRbss/44ezpA1cfV41LX9GIHjP2rWyMdHX4lVJTgNegkuMRVEXkAVAGUTsyiILR4j
N5xxoISTs55Fg1tvPugreUQ2Y1cC37Ff5nVlRbHgrg400RwUIE4bcxbRTrH7sJR/PTD6va6tTX8q
/d4ZQ86DYucsNSbeChNWixXEPIK5tpbgZpPRWq2CNDarPnVlfo0jSc0YmvlOaZH7TnlOhsDyMhWY
LzcaCCtSOn4HzCVchAquRkrdlOPtQUCCAmQ2INDwkeAtGoxYw5P282Zne3/fuYJSwzDvF0d2/W6x
PJdB7KlA3Xfzcxah3xWUfRUHG3SpQ2TGvz8sUR0AfJeXd7y6uug4KN3ErhpdxRepUGXKybO99OxS
fZCmcPfz5/JkxxUyQsie6KYp+jfEH/HzkKWROBy5EEPgf3naZiruBo5RonpMOfAmfa6gE3zERqSd
CVCC8ZSpamSZ1qLCDshR3xtOXhsznKR2ah23VCCd+PPXrEBQMkZ0ZqQMRwHluAflG2q7UIMAsjTc
W6qv3UjlAznOE+Jzq77HwRE04EixsHE5KQR4pFUtP9aRv3dMECDSXzvwZTKCUzIHu5uKjHzjGaGg
uPyoVSB88j0A83nvrLPepfNpLKFt/sLMnplmz89cx1ZXLu+67MRPUXPy38HBPmJRvSo6r8HLDA5q
8Tq4J6Eem1n9peoQh6r6wm5DxkzW6IRVk4m6tREnoYY2k8PAFtno+LtbP9W5XOhlYAEsG1JcwbVY
XQDz+NmoLvdK53NIIRmrMU+YNToRmXgFS9Kz8t6reDMtGvtkJbHu8/zJkYeHAD5fk0M8Yxr/AtAt
Iffthzz22lSApteSy50Zf0/n1l/cAh6wUkr6S5yYlg36eAxwN0jfm5hxeaINQLLrWF/4Jlbo1a2l
Y7PxEqk9gxJhfPvkiH9PLrlepGQFjLNdlbMoba2v6RCfWGMMWZuXA03JFzOUA+vyPnQubSNpTUUt
neW1tkrnO/FGr3MjujOAOco/80qByvNhota/PsDiWi/odKUWAbI9a7RNdyDf94NqGmnF52mnAsOS
J1yusiPVpDNuNHExw3wRwZ1h8d7Q+Mm7z1M4lzGxTS5tKJaICQLkuy4uLXahePB15nbEyFpyT2u0
B8UU2o6opSwz8htJEIufhJYo1vDxCK4fGXVFjcL5jLTexsvAYRVZVgNwxXq5URtE4oshv3IzgUvM
QifKVDVLfwxkt+Ox/BFNKwI9c/XlangWOF6T9Ku1wrBYyr56KZ49/PD4rjnJ3zA49yBoKx+3OXmd
aXgtuozVODarykEvGGoG39rjm4JOwENEN3uYklnnAoxdrP6SBWXjz7TMZtjqB1GAXj7HeFQbjwLa
hiLZvB2V5E+XEKsPjBmEdN9wd3GA2pKG7aAOcnEulqQaUkNzN+KL5DsGrpx6tF3vr1Poq2PuNmAv
5NjUbktCImFJVl6VnpWW2PogKFjO99hUlEaUxRFnnYbmxxIh80jJcV+cbx5bViiBFFcMAZe0o/p4
j8QjrOBI4X6YV3pVAS1K34wOMfsiYZtee7fGUyfMclffQ1oVV3qahgWqexT6E6UG0AYi+tyLlb7J
6cCrCVWeudQOJkZmGi2AbUmSjPlDtMmU15nQSNdXU4uZJYfd8QE16kU38HoQiICfA/4ZWXRju4Tx
Jd8x08C/CuQRiVYZ1tS76Mh4Od51InHb3F1FgaR2H8K9xKIllF6vGp8d4UZzjdBMRL1Eg3Ux4UPW
JjoOjmbvjRtkVkQSIyl1SlgeZ2hL0GIL9sXWkKVbQBFQ4oEi5V5UsE90Ol/wTRXx7MtziwDQJTPn
9GwXTkeTrcnAmzMMUUG3iUCd7I/7kpQPtESTqGFRR0u/1EZlI0Rqo4wXdcHJ0bYJ8uPjenJTcCeK
8hzGifyMP3UFX7MlB+w8mibh+vSECnrKtMC+JqEo85XcRAhf1oLObl1T8fdgkTx/vqRdL9lX12eb
jFX8SOtQxmBlm1oB2FDN+yVUsVavkLJZqb709IWueScyj6dQjoXKYOgo7y566rQPHiQMG0z0Nu5U
IR+39V2vSExA75Vz2NYSNZJ3eltHRqvLi1DJ5vnfnU9ltt4cmI7wnKPfgCZLlXhxIaCQwWFjLB7N
HpIEzHV8ZeuPelrhUbywx8JOKRe/Lu41ZrGF4Ezk21z5kkS4wR4Szi+LUEhpxF8ffe/eQ5RAMVrc
uVoI9utRJcpgzK+WX242/gEQtA9sJ8YwQ0LgkJHCZ1UNST5UxYyJ+JYNcfenJZl6+cvkwi9Nnz1R
In3asEVqO6gMsasvBpRQVc1kVBiARmUGOrg+DhQEMMnSPOCvc0o65nJvIdMwJnewndGV69aTrCKK
jFMXKWq9rDhwqiqJD95bUYD0DWj05vlnu1T3Ms1MRWJfnbbxebyt2QpXwCtQw/4jivep1vkkIZ7E
bqZTXbi4nVRX+TZ2kwrUnIAkg/lhBUKX2FZl2/+77qBK01a7E5zpOy6/0d2DKLKmlKWNW9Lhpmnq
+eifCOXG9bUCvkjL0WQjDGPJ1i/hVhRnud0zQ5HibF1Mgrx8PN9laKktbuRyhlqklmx4SphWxMYn
9TlD1LRwkMyLBK3byNeJ6YtB82jzuvAueBtRf6dx86+iJZ8AMguSH6EsGGf/e5pPx5Dz5i/lBs7a
tWSagVIZJtdS9YMkMuMf6lOu8ri17AyMeyThGKwkh4TERQLI6FeVrAeecJCfJ+ITtr3hpflZS3nD
wvyWuVrSktKl5qyn0N+wgpWtXH1HnZmda71yqOV46p1a3yOD8+LJDt8LxPw8isvKRn2s6VFz0J7N
ALmHU0+CXlWR1F0jJhkHfQDjuektrk60Ad230/WwfTJxu07aQi/+q5Ei4slgWsMb3KqEjP197+S5
5JOSFC2kNAGPa7JRCE7HAVo21evb3ZqU1EUjjb7M+Oz9/0Sq2z9E1HblmXeyf0Kr3Se8uqrvoE/g
N3OXu72/0z+FnyxvurhiQ+6/zYfUJGVMtVFd416ebk7LDya6jebOVHFs6Sej/YRKKZ10x433ZVv7
dOy0l23jJ2Hx0cYejXgkk0ULIFFRsPVIq4XHSFfx1ZCCIDHYVXzyLtkAVKyqqx+CmCq/B+OgcVJ4
HdPYKBqdpydnFfRDCE0rdr9ud+IW4JejwbndJBkBvnM1Dvdsxv2PYwYDCsAPJyI0ZTN+IcaGZflt
oXIjPkx7gtZKded4P74FUh2TiXaLkKlu9XuVOuPOUMPj3BxcSWvneErkxPEei6wzmzn44F+0D5nQ
J11aYPjffFJVeRVrcQarn26P7LJnqc8AVhpmme3+uOi1kWKpKAXrIKMO6a7B+D8OsNgm3ObETXsV
alcyx6TExZC5mh95f95RXNav/yIv8Fc6oDIxC/h+75rw2TP+do1oH0Sxy2/fBMu2FB57zcrACD73
/1m254KUjo6cED/o2Wuky2YBQHxZg3oIVGgfkKRwdwnpOgUqBJb7PGZtpsjrOgLG/JicNCIHzwj+
pzMRIf2j4vCNJB+7QRiueX/lWaWYAmnwGyz6rcgnstXAJhcgLbxrOQmGK+2ZfQGjZM+Ii0Ln8E8G
9a/rO0iOI/wJPsW4x3ILgF5nyfn5d4bjiwk/qdpGYgOgSGUkeGvu27DAWqB3A8aKgTKqWShYqHB5
TsmSjaTW5Qb7cD3BfA9HTPbXmiNav4IEz93fq1ORzBvgsEfL43M8yG6fVOA6s3d0sThuOlQIWV7u
WDG83wtqZOmhO5mlf4xMZye+MVwoYnp+01EfQV02M/r2ueF7rm8GcNllHjVfT/gv9flgySZmqqv1
ys5kZq7xxK3kormrRhurdut5+FnbHyNlosg2/qeP4Vpetk1Bn1+X9nd98jxCbZs0Th5f5tcd0r62
ySKw968p7N1TNUN3ffsxwPH7MWtsejS05bzh525eKA0ecfemPJpCm0WaguYV9/sNq59UrBNhJe5B
sJfqsawTHsH58qfVjLMRC+cDqAq74sbSfbkJYVZW/vDgzjolUS1uvn80EuFwcl9sa8IE1LuA6kLF
YYwkdWB7uCw6Ylle4b5uC/tzljdzy1zn3M/2u/bFoMkO38S5FXuYeRN+SF8T/NTuEVKeqUKnAWJd
yQI7MCA8bxWeAU96QZivw7zkSr77N6Z+utmjsvUui4iZOJlAgFse37dfBJCYMwyuezU3RA2IS4np
smwEy4QXnjDFfhqAed1Zv0bZdeIUWWF4taA+LlEJUPrdc09Q1jpa68C127UkOW4R4/WmH9QmYsHv
Ms/MBLjcS+TfqCcaFCowphmIVGaeodT8Ix0qY3LGqm9RDia6927db3O4SFZzt5cfGCyLNjFeN4wx
VoRpaMJ+mjeMEfWZ8kbxPr/XiKOWQ9sRGRkBbKdE3LRm1OL0AyGttlFBRrKHitFF+9LHy8q/0kh+
mVe0TTe8r9okCKpOrn8MhXI8nZ/j8UmHSw86FQ0CT6jF+5Brie5q4E+I5F4sbUHUsbnalj/DwO3J
LgxGvW+dYIfSdoRZpyGkxj2lEVDlce1Bx+F0aWAcYgEQdUZz1ZbI8D91ZB+29ebGiVPssBPrTviU
PQ6jOf1vwWnTum5NidafFah+IiI8JdhDT+LR5mPvIeZm9uXJ/VLkZzjqQaXt6lGNI/+B9rp/B9K1
F4pd8ySPLNrkLzpuIg4RLkdttWvOy8n6hK/ObWzhUeD3594CDAk/DJwBYfCs6WiXDAjlvLoCyaQA
k8hHWidwik1FSC9MlXP4SOmWSRKsvWuq9fkbRKSq3ni/jYNZfBpFsd224iteVT73Aq+UyO+/zSm/
7MEk85ZrtHBwe3KMTXCsHRgy7gdcdM23mQMLxI8FB89W3AilaFGjYEVWamKY4oPv2Jrw68ecU8qB
AhVAVPji8OlSWIgzMoGQl+cNyhCVZHD1rHD2JHjWVbVFlJUEnW17lZowrlbdevvDf12W2BDDJktS
2kQ4Dkpw04UJI8gRhaPGMZ0IPWcJyry7/J84OkpiZXar3mrXlV0zP0H87V6fXVup2Ssuv+6vSyKy
fLgCXrbEAuY+c47FX3il3rZVJ03TX7wkRDSLf+8g2nLJz02EGQBFCUgkehzgYFIUrFArvfDexjzm
KMaTzFD5dsM2S5fz0np7FYRCFDMee3WeuH3956hL5xRof0h/348OkmyMD0J7jdor1HTZvhMHrlrg
bumfZtd7m2h5rFMn3rVNBvYcixH/UsD5xuOzKUTBTFfvILoGTzEiLuPq3S4tXPMnKkbb5Lv/v9fc
881bAZc0AFkFyOr2I+T3g4Fp5gcWyzvuWKyF0bx5FY9Ybsuh+EPSsHdpem8sSJmy56npnZqH03fc
hDpNpLprRhFouLyUdbU38I+bHkBdqhFgQDHt4Q8pO04Zaleae5sdRqe1+QB6rP8l9pPtP1WO9HcM
H8bZa7/xi4BJu8ryhWwz14tY4JqlV0h2TRIsuKzALEIKo2U6IlRFRZlowEVawCbDeG4uQO/3XjvW
VOpDQx6aZAbMkhy0Wzq7r+HyYdbDBtTzmbSXr9REz+GQ0C6l+3+VRGfIOPgpcc6V2Ulk8ba6+71P
bvVPMYn4LdfpP5fOP1YWHQOI3nvXWMuG364RYd/+pwEB22ZS98chT6uS306Fm3CypnIBlAul5GfJ
jfMiy/uuQAKXjqkGGezu+qZeickCSGyqnxuwnGz4V6Dm45BC/Yk4nCcC5TqthN+f9vxPfx8w8zFf
+37lYRJyxeXIpOIrCoCrFsLznZosebWeFyfALRcmnE8UrucOYjO9baMw4BdOJFAoZWZrmHYYFNEq
2dictGRIeKmu5ZP4YSEJbyR2muaJm5Fhbtcm6KohPOF9almvftjWVwAMVGIpo/njyOa9CEiRM5em
RLSelV+o39cDZjdDB5R4pvw4A1CXYtr+hkxmGnJMK/AYKprtJybGoM6ZsA6oD6EpprP/91dJ2nRl
9Qsb98gXKS9820pYh930d6TlVm0k6wNbTe6edooQd020aciqrlne5CpcG3FlCqgkDidv1OtfnmyH
iGNiaWzUvOOYAtHWLdPWIiHsim2wzg171utwEm6wMiz3fYP/QeuNqKhIA58YPhmwKXJGkfnJ1jst
P7yxLZP0lKiojsRIYbZOVH0tBue9paL75zak/lJty+ID5hf/9WYdbUfxDjQ1lIWStXyDPYslTXes
fBAZmRtqkoJAUW3kGpS6dKyCuV9OZYdP7+PW9AvWKdqhXqQCKC5Pu0rYvgzM/LnGX3RIWpAjLyjH
Rp6FqzFV+jD0CsQRrYc7jHXHwny6OlDIQpxl6j57lmEawYaEhgk+7nE74o4LCymaOVu9jM1L/P55
GUKcXPs4A9hDV1JiwZFR0ptZlgs/lFCgTLykgK8a/PC0QdGrxQfFA+9/9rC6kVeAQ1J8CGFjmyis
hDneb+jJzUZug7mIwqUYsZItS4dvG/evBSc8wbPl8xKkBvgfnpzPJRvfVP+a2Q114367/ZE6Tzd9
UkHKyAlMylq6sbs/zxiEnTd3tiqbmAjSZLb4HOxyvucVtO/XPP0VkC+iQt0Vtl+tbhxBJI8W3Odo
0wNbVWhaqyIRnlcf4exbRUo3DG0vqDtlPM6MDdeOHuuuAN1L4+nVoF/cqeV8VgGh4k6HU/Ta+1Ec
v0V/BrqO+WPtWwH2vJW54CEjh/83HXr++ft4o3OcgaxtkMM78fLD0wK5eCOQG/1z+xvyR4mhxj8G
uld252YL19l4rE/S6qbsxkwkfUxFkLR848BcdnZHjcc5XbzoGNZr0lotyu7PFFxSG6gNTlyBVyvq
MwWKFG3TGrcZCgEyIb/TYA4ysWPluHyK9deJ9XhwxEaLrwRiA0fnfuoGIy54DvpT9oFYukF8+1qb
kV49L0ouOOi4X2TG8RuWpHb7ABqvIAi1ANkQBaM6jtx0dbxfopwrTd2LVTC8x1C+a8G48Dyq7Cis
CtEgZqMxc6Xc8TUsgOS3qrSJgPTVR7M3NXBRvjTbcRJWtXLvZoRVJVRb/ITLOmY7jFgwiSxuCoGA
2W6Rub2XTzNBqX9+lzbFZqVlgfMOi/XXM73ntLKgD+rNwWrcL0P3v6fyyk/ssMkiQKwSKJ566IkO
swZRmxfvdSfSbDLF/60EX1ImPMGAMCm2BbbfXNHkRZkTFBx1rMToZKwe0S7k8SHa/b2k29pfJWtZ
ZUUe9f+HCni1wW2Wt/uUXkD1/5T3OL2BP+Q/BX1vVo/MEbvAjjw1mqxvMVk+Iv2GdSkSv/CjCmDB
1xOLh9k8i6B2uuGsuIXrZ/UPsTu5ZbYZy7y5mk39KkIufEh6V0Yh4SKtNTqoBlZsSjqV72Ql07LC
Z49ZvI8TXVlVq/XecxTkSE+MdHeIR1tYGxMaHE1kfTUEp0LS85QM50aeMkh1JVEDBDCNHPXMXp1W
AaVRT/18yt/btf3PpsouRGSpdT1Zfqw2p23sHwEwPfE4dMPoX6FaGw0VSKdlBCfFL+st5lCD/wng
+7/IK7EhvTdgrebVOUqQZDE30/CrdVg7uRGxNPYXhBaAFKtnsu5cDZPHpbX+sS8l5HW9cLvWOPiM
O/EXuoGyHRxK4K8wTAY5g4b6mu27uTax2xZULXiiprUSnysnCDlYSbp3NEiSLjP2WrS1siPQzMrw
wdme4THP4/w29wDCtEuKTSGRB+5i1wC4tiLPXZAWMBcwwxttW0L4uZfeJjk7xQFW9hOACd63Wl0y
LJnPyO+vm9BRhjIwDDEbQKgmJR39G8uvFFePnfXmtBMf8k9mM9uRZHBAPlV3LASj8wQGNMC3uIaZ
2WRGku8+hTt72PasJozlAYZRDJCObYIzORlYDANpQ9vPZuU1EaYDwrkQc+kNjle5Kr5oQjvSdDHn
X1PhGyBzXw5ROdCljF2tSvb0kz377L2vMVjv/hqnJUHm3ko7XJ6IbR+J+K2v865yJzueGo0s3oU5
ZTnBqmjDUiJCFgqmSXWYaWQW34R7nljI4F+gko0+xXUnxh2HC2RtupMY5IM27DT+ZHKyf8iyUdeF
BdLDmAmBxaQSl4K+dmOUPy2V7Cn4CCSTd1kVST0YcfXpeBMj6LAO/GPAU/+CMoNRIp9iZrU+dEik
Pm8pDvyb2i8WT9d/ueRuwrSXXY+fhN3M77R2hao5nq1AOZPup2ww5axRMJzIbuYVJ6qgM/52olUO
pXY9/K0pkUrB4Xoc4ti758xjMY6JcAsIACKdOj6iufrgSoKI0wEi6Y3QaBgnc1TndnnyXgibUAPn
ocd6ABb3Y0oq7arRC/AwOwur0BD0Trenwo5gvAp3gl6m3rS3PKZ1H2UaPYcdqG3Um/hjbEZEreMa
OAqMslpA11YDGYV7DMhNuXtjVG2A0wY7iEcL4tMs4Vk0OvnYIwWg9ff8UuHUj50TxzouCi0S/4YP
ddJwo9DDj/WLRRiduv0zKqsJHGdxV03UB2rnPHeiDQEhEG6Mi5B/vkSH4zOMjCByl+zbQdNtYUSu
wNTPuGw4v2TDyGfVLkVC27itqAU6zNF07ljMVjjwMCGyo/6xnvA41yARZs5CFOS4Dt1OGVLa27YQ
7q2fYIKGgomjdzfjRjz8odisQNSzRFGrASJQvRHZq3r+7qBUUjr2klT6+mHeFFxjFJp83+useZ8+
WDsb4xZ3p9XwIdM5LMYLwwmvfDvhNTZBPhFb/TABbVKvqRuF6lpvIveCq9lQruO5TE7gmoEn+29H
1jDSJzPgj9iVYZgWudfxwOROQvhpq5TRWV15dSnxiR5E38YCV/ZA3/BtZI29OtBgfKVxtxs/Im7i
10WQru9dvPjOOKLGn0r2wsAGBGf6t1KriO9mG6MjUU5fzpJc8RiKdvRHuMTL5y4SwUpuVjeLRoa3
+MyNj3n8dYeKVMtl7XIawudUzPnvbB4R6Dcz5LNSrNYQovAB0Q9giVcw+XswCYFqQ70UqZnrzaBt
Rf3aD1h5Qz6Awcl6Eqb1Wf/jCQVUUi+MZc0+ZYOg1rA7gx3yde3xkwy3Pcbk8s+0Ed1+XNBcveLy
QVyk3QijWHSXBqeQLoN4n3qjF25F4NhUSpE+FugIo9rHdsP9LnGb+pnoLHjzWswUk0Sls7JNVnq9
nmz5uNrpqe7I0ECOwTXv09kIqHBt/Bz01iIO8m6jm6aue5oaQBHvt7+/v6fzlqk1WL0tCk5y6uEx
tpDTGml/drzx11zs/FTo78Vr7Buh5fWG3aBn8EMZMlFX4+ydW9sPsY0MBzDgSYDdpD/Elh2YmEhr
KkkLHTDEwUxWtV+BnCNnVkt1mqhaxFKLXRBc8RsWgzJlbzTgwCpPrqQEiovkAVMf82r36U/sjVsm
HcL6IWMi0uyKijG40k1wXpuJvrmGTbYOJvUz1cMwOPU2z2uvlBUigvDl9iI+lvgE/X7AIFC2LejZ
vEBvcY+W3mkh21ib40xfHKrZbU0CSaSYQIs9YbgYy0pLHdPaJm6LLosyw/76a5frenI0N+tqgHWY
HzZnGJOa0CRfgqrD/89rno0tsMxGX+dY7Z42ixOREEUz5SbHlutHXX6QaAkFBgXSlkT76hvwmY1p
h3QIG5AhpFNQ6+i/TREq71Ujz2neWuI4IrbymatzRZOsPOFKrWzS7soVEXV5Ea1Oe/UrN4gpUbf4
Zo5r3mOp7fAewZQG82aHyn/YMDXMR904CN/YpeyT8ugZhXUpE8AcJkTirDrDJSErUwu4x9VfdWQ9
ql/ZnYKTenOPMP0KheOP9G9lufMtnfTcuvS9f/XeILebyj2ckpODzPCS+iRIopXWgkoJKbTADsG0
QNg59OybzBLhGBvfF3uup0c7kWwM+gjGVoTxPoj2QjsVb/bfaNeRbfqCEP9hTUiFYGyIqiTkUCYF
8FLHw2Vr0KfEy6MXgN94qoXxAkADpLNWDXTdFgWdh2PpZ77ibmP565565X4aXL1aRH+05E6SAkNB
CIJUFScVek52+U4yHWpwF2hMfwn7j3ALBf3rqs9NkAyts4BCzasomZUhCADk4l52BulEj42kZ7B0
hn1DH7QgJ1jnfVT9jySty2TaOwTPCrTMA0cLSuFIma6yI9Gau0D5hUUxQ2SV1CvhdrgomtHD1vc5
EF2I1HpCb9oufxkXxx02uft3j4iW+tnoH5Vqi+J5X5+N3lMcRYtrR6aXngM2XoVXt1xbvqo1AxCf
lzPPdYv/cKbIe4u6nUrlwnXNbjhkUh3jkFiMQ9XdPECxmPN2/DnUTjxVXyzrwD3VmLxzafmazQeH
8PrzYKxJh1B8e5WVGwXWxz38z4lfdkF598L1AV5X0No6sYex6kwjSJ4jQ61AIAiHb80rVpgC8DVp
c51DF8M0HhStb/MA2FFiQP7LB5i6gCEcK28TPtna8O4oeSLhn5IJXWEzIy2NDcCg/9arWzkIrxYD
LMX3rjHlDaP/WToTlEAzFOsFWrAn2CSpyhvMnHM2O+DzWAvSWHQgxX1Qvadw/siQWxB9ZESZnqM9
KbOE6VqwtiwCUW/DXjePyvI3ZPZohAKRH1Ym7xGq3e5REdug1RlADSF8QguD4xFkGHypvyFPxuVI
nyiR4hv9Drm62Jhibs6Z9y/p3fsBJY/Wb5UcJu8uI/iCA36FjyjP7Wx+dtuvqtLkLY6BsBses4cS
Bwt/Ckn+W3K7oqiiooQrx634mwY6rvHU0BI/W7sLpa23a8XrTASKFzyZm3c9v44Tr5F7ohkD+xNv
kdmyC7U23tkF22+/Zr+atILd+AF1EMRcQAUrtO1B38gWsXoZcwubmM2JqWoDj4HgZ7Y0kFoYmM8q
IrDCks5e0L8+hwNPDPRZTa6IMpIyyZeW5K6VNiPl2lrDM5a2S2zDn/yOfSD/r27U8ZeNKD0PNf3U
EoPy0kpG2HNcvj+L2S1l+Gocy4tdUp9xVLa5g8s/KbQj9NbAh+XKfaTuUpc4TYsS3JYM9q97hTI2
K/52+Z2TwSaTt57hHu8Q+Gs5nq4WzJNKnk6NomCtguuxst+TNgMfNfTz+WCI1ltjzuVgvz4RJNQA
iTR08nxlv6guvSL2LfxueQZyxv/7sV5uitsjfSSz1XftCqcLMSI8Q8FxrF68u1FRQpgbtkuwaum1
D2NHyiDgwG4CI2AMl6cs0WIb8TIKh2GS83Vy6YdRv3gr0awujQGL09rMayjArg9KBiQpbCYeFLeg
wus8/ML8HXbnuR/n2jCl7igAFSfylyWpVWg7088YfhA+icpiO+y1KBl6tbnstztIm9gVVghkG/Dl
mhvR9aoQDKqeHak7i81cMBp/74uDJqlbHOLRjBNc3C2qBG6K8huJrWM74MXZNOBViOzF0ifn8n58
qJtp3FrxF6ae3rucRRwIi1BBMao1H/91zOx8m3YnYEehnSUM2jBxwJRVYXhNXyqAZdTYZqlM9y9p
JI3cpsAbU+MzyxrZ58ar15Tp+kACk87Ylu548LbMilRgp/6vz57eVSnHrr5yXRAw6VuXFenGpp41
ab7J/A3xB/uKsJCbYe15TqUXOlZU7OVbWjMdTdfvYccG8onIOIOmwoN7Xb5JiEqVtJnKixtp3TAO
KmR+R323jjTbb8VVrpem40Axf154XGy/bCT9EOnUTi9lRptlNr9E6mHWLolNdm94Ir+9Hpzat+R8
SYHkcrFc13ZsUWzpNvNmudEr+wJudPQFfOe6QhQSdXrmIjDid8gH6/oEOxyoXp10y9/hPLWBMkMb
nAQrT9WfMmKLPAirLrZd1d63f7LJfpxdDDObPJ2BK310+VTXnu0RnNrt1kHGDory4c9L1V6/S3LU
93+f90yQHbjPa15xF4UewHX5UUjSKYjfg2jq2h/vv4qVNh+O4G4/OqpmX70+VuNbGrSyz/jsBa6C
zCiZRxD5KHJSLYoeM0iQLTWmWZhut6xPJEc0v6LRKgBglSs+6cBxRpvBk0+IvN5ng9Om7++zYnzX
GKUcyDXAgk86gE1e/O+D4VDllh8VXz8t9zO6rpWfCOip6s6q6YHPj5AnLq5HZGxPklSmAlicfhWp
27Wj0FJsCb+cFQGp/1NmdBQo/HK7kMujTZpPGDbjyQvflWrVVijPYmb7rLA+kLew2h7Kjhyo61UW
2VQO+WARK1AMRAeNMO5V7X77mxWGhkgtyn96YrCjhSG/Es/FdCtcXF+b+nGp//vkkrm6o6jT8U9d
hl2DX1Unh4aQY2daFW7YrnayzpAnASypAr4rSiWSzdLVT38o3aTYFgnEW69kXqBLIJ/u3bZ+rlbn
9o+I+W2NT1qA3u8VJOl5a1dDnL2hg0q/z9ZMXTvSUfAqJ9584UV7w8TlyAdsDOXtiOHPsIAPuLjD
9UMe3wROpq8eKQ78OGOTWTmu7PtVgt7prvZwfTQQ0nJjXq8UxgwZ/1fEwEw+GukVULXE2m13F0SX
y/uQ6iMyXYhmf3DhlrPGHT4mkpkqC5cFhtyz8XNY7m/8fK38FWFJHFZvp9X4OexsjoW5q06aQgDy
3K213MK6QolYnFs/TrVtUep3+hGKoNZwuhlH2XNYdTwKsdW6aplgHE+dl2jtD/SsrJ3BTMN0yzV/
z8+CDXXiiuyLf0UYX7zeFZm8q7AzFHGkQyobiz0cV2Qo3KT/lhjX/L+/rkHW/OksTBXnU9Eh/150
o5scY4rstpde7NTzxlYEwrN3nawJvNIjwBSd2itjwD94lcISFq6WPkmDYcFC0c1xkiodWqJvDtpZ
a0WqEvSdYdBhVVQOwEMkMRJnKzUgIV5SCrzOCj4BOcxZ9F/eCXMetamieS+haP+z/EX5cPVDUBi/
sF3kuF7fZiAiJ3Hh0q+cI4lmM6X1bJ9Les5Bw6EoWt534naNH47ycE76jjb0ieBjsESCwZLq3umV
xijLIMuqHvflUOCukiRWkK+FlyetxX8/91Vx6xcQi1PO/lXDcm2k37YiCDHkX8RX0Qb2Ja4P0pD3
4yFr9OrcBAOE0AiluJSBEsJJDY2ZMLEbT6Brjcp8jGzDRMmLDqQxhkS2+pL2INM2dPqFy9SblIr3
ywL4ujB4lKlpmwCyiSwmD55T1fnZnlFI5sb7bsnemOvMeXrdgpu27gqgH367HUWrc98g8hFZyldU
XhK7KoOxtAqwGPrNFkkpACv5p5X9pdXhKzL8wykvod3JEfpfxcOMvoYkCLxgw+Q3EF2abRXYzZVK
YHyrn9125JH08jfF0bzfvJ+QOS4Uj/cGJ3dri+UzOSwG6iA3I0Z+Fo6ay+eEwdEUqDGCyavdZu6p
rFk4CJaDg6HiWrFt207m3QBrInGgvyxlVoartVyjOXJ88T2z0KVfM5j0FaVqBsoKKbOjD2bRZmKa
fSDHyX91CaarmSFuKsxlcbAx6bwPTgvLBfgsu8FYf60kVWLiKHNVjle2s9GlmF1eX+34Y98ioOOB
cXvxZqXB/nX5rY5xuQhFameMJ2R5V7nhB8xUseVnXIY/5v3Qru6UUP20nAcwGb4/1rDmc0as4JEp
B6yZ95c6MvMCH4WoYbketcrPUfx0Z0LnsspSJ8OSLjaP3JVclsi88pqwdkffAN1SkJxxPqWGnpPm
w3KU7U+lwqb6Ds0TN8ofbMuBg2JYNlkJp4WLHsTRHTOvF1KIdxqCgJqa7B6DraeUzdjuq98tnGho
r+hGFg34QmlgRu4Yhh/FR3zCKu2ydYAwX+pGmp+mbR5Z14aNvImHoNfVq5g4vNqOvxEtUy+ppaJB
6DZ4F0UQWakg7gD0nGQOMduk/iCG7tDWyPZdBHCLaDIzGQ2PWwjXmPQYAEVJRY4OhLBhf4oMauwT
cpA7oEcO1J8wFNL+QYqu2imnQ1B2wk7O5QyxWn1eh5bfPgbypcOtU0N57KGYLNtBGaIrBkyVSeUV
sQkw09TaMucb7qAIKSSMlaZpL78q2kSZJSWsd9LA+nD4ZvDJIU9ny7rSp/kkzrvAeSRhg88fV7AT
hKphs8XH31049I3QWRLhykahjVs2k4idh1NrccqZYKKQdr9WOuo+MsiQ53oFlFiTzEy9w2j2KA8n
WJBeB9i3FUcTi6RdFYhhVyJk4sFdIzvahfIgg+e3C2TEBAm5ZN5xn1Hw7ux54AM8j65pu2BANhqm
KgSGVBYP09GGbo8KeQZHE7t5UocHwm/6Odqsr4k2BMIwMgXUxzbG4ccsJCto2VKcz9jt0agLHY4C
SQF+I/xs5/w9uqTVmaTw4YPk8OaqvyiwuPBgUae2FvmPff+4CYJr8ne4Wcc+W1TBUy3HXXr0Hckm
CwfB0gmuFYbEErMcGobAkA36JzsMNbieFsOtFfoJFLKwV7i2ZmIhwh7rX6HDfrUjfdNYl7ZCzXWp
hS42IQGVjlMuU4xQx0lri/6HAMcF6Sa5b4Ps4nYsm7juXAWlyiYrGzzDzUbtO2YBwGoecujfLPAr
XzCRr0Xh5Bt5PZZiLyMPpW+8RAO3Zo4N8ND9AvL5FkYlmoByPEUwaNVk3oE5BPg+bGp5XLZ32pGu
QO0y8uKl8HqP77fcxFcEiWxb58GcXvZZXT1e0Aeq2uN3gVoioEj0pKlnvq3Sem6YFmLktlFly60j
5kTJ/8n/dm8Itlu1M/tLDzF4+jsVfV4Ezo6uo7NZAYE++gICX8sKrzaTS/YBXTQHcUqEEC5EHLxG
Uxn4VewWooZNDIh4CHmBe+1IpOe65Byx5QU6xjZJbQFiVBlqlE7PYpr7P2qwBwdACbkdsfESaelU
bk/A1bLvnW47X8pwk8vRmtA/i55ZxA8L2K3KYs1kqaektobgAVgWisy8k9uOwqzvT64WcqnGO5zn
SYZ52Zx/zzfvgH1958YND3uiJ9dsVzUsEaQGWhYCkCTeAKxw8jK3L46FgXu8XhNEEzzMEChJ/4KW
JCXlpHflpfX4VkcIskrOlpv3TTTldJD8T1Qn9P4/25wK8VF/7A7HBmfvkR3nGV3AO12g4fgJFJxa
xD91DJcuC5l1kRm7rkleurtO44lGwjTrbwgSoOjeCYsClwjUj5ljykjcP52RWJIzDYTtIDzAjLBz
HkrX/hVHFLc0Mp6lGb+zkqVnuByMoh+rRTON8zbyfmH3u9C+8FOHjFP0OPT5A+juN+JF4bKIfRqe
784cdv0ggct3o2hY2jO2ouQEzGRfZUGzeB8WSkn90UNvLLA1UYm48v9q7RXH7CDs36r2C2At9vGt
jF/iZQKlSUaMmFnJJP/O19ytGp3biXETplCujFIMMqC8R7pQxmQz2t2uQ/dYsQEk1Ai2Pcp2Slf/
ykJiO8sMEhKEXZLbkoMOi1+19YWzctY6WMSVrkfzNHtwY1RGVLygzd5H+betXuX98JeL1cM58g2g
Qsw1L++sj40ePfKEiHY5gQ/lKrGFBWETC6JPbDbgKRzHVIttNbJ2vasWWWq5Jd4ZpUoCUx5g4EAc
FDKjx1OuZ0qTUbaJR8VaF+K5aZb3K7MdOJK3DdFW9bcI+16bS85lhthwV8RpQ0osvB+lHb9OHQve
Z8aEk69eAHDLMI/wiaMSs0k90i7lEYqjULv9azpcZeXbDS9klVD8sMBa5s95Hdtweo5ZRB48UUYx
tUNX5CYYx8xXJ/nwKDFEC7674+MbdU5w7Q6Yc1L+xy9k2BdJqEIrP99+9UdxD5bpAjDN64fWGhIj
c/659w+a2I7Kz4cuHzCn2ZFwdvwE04MTflN6sbzfKkeyan4C+SgaRqccgOZN6Nqrc4ufrdjhKZ3v
oNOugg55kmveuM/0hghXXqNHvpT95OcETNSn0xG9jY0O3vZ3Xazt+3nrsJYUd8ePAetMWDPr4FyO
GWj58xY0vTwBvsQw+eBe2FT6wqEGFqkXgOAzdPvCLSVpXIZI4+noolg6/ivprzIX9+NzC9U/aZ1o
IvFTjW7FjomMLkVEsmTd798JD0ebQeAF8LQ76MoBylH9WOju+loPwJybNo02J87hjgLTQPtSYoSp
TsM5BBSGA3xPe9nRbFXFG2ePP62u6QUQOx+2MeIeS/NxbCJkIdOvABCCq4Tw/jYAyoc47Nx4p3V5
QnU6bF3mC5KDGl8NHF663/xj0a9l9TxQAOvH9vcfLXK595j2czjomhyVpHL8xHsvKZRgdX07W8Vr
OWuObq35Sji0gMhTU3+CxsBa49uAxG3/fihAJnzghYnTOq9RRYuDXRFymfeldh4Dx1oYgASv2e9m
JCCoUFjxTs2jcKyA7hf9GHWAEw5C+2MZYEAtbZxHMSoUbgzR4s3mP237LNe/EDKUy7lpLnpk+H40
AOnCO5mQ5OZK4KLzNhjtCXoTq103yocCBjKjaVOWL7ai7c311imjsX0tcFa16mSYpWhjzQRP83np
MDDK2Elh743iaT+CGFIfQv0JRJSuHoDYKz36Mpnhv2kdFCvUDieJcK5aVnrpBG+gW5ZPZJ4NutNT
6sDKrpDDKhpXJVhYPaoWW+ICvV1zizSASJ5OQjDjBemnjpkzh0oEXJIqEz9ClNunaalYCqbo5RE0
0TaSTeZEEJkibxhh1+EJ+8YfI/b8wHnF60cqTsQDgQic1GocVDk6Zv7nOw/hwXyIYloUpOqendO+
vdWAJcQfIaJIwe1Bm1dwwcxVez+rvd7T6DlEosodsH1XRcGMpV/ycvChNxdYoyzVWu5FsWYisACK
pRgND3jlgny1YO4/ygQG17RHBmlhEK1CXfO4vM6NsfyC20QJep9DEtoH+LyZzT/gnIAWlTggXYfk
XoMqBT6uuAoSzOhU109V15oSvHmvN0faZ4I4059twSLTrsTcaXpNbJhYO6N2DuCrL7DJUsSxr1gU
N2B2f0D1NzJgSaCbOYbi+ubkz5A0d15hhtmXHRXZvXnT/K1bL1tQ8qarWn1/IcMuYcXUTNZOMAOo
aaUUHjdpvVAC5MuHo6+FUvAErkxoNkxsrhgsQvFY5gkRHQeDRL6yfIUUxLYVYidn/nJD3hMt3/dy
vuT4rL2P5MSs4kAzV98Ao9myJrpYQXdIAujOXu3LiOFnyurBo1mUmEefTXdqBId4zuXTD2ncWxAx
W5Wlkzf70OuNfNMNRkMrgtLEddUlZNt8d6zkfrLH24odVCOfElF03asxYs6wLdEIaX3vh2lOL4bf
K+1+MCZkS8ReQLxdZCO1K1v/SvIK6RZWw4fJIrMY7hxUfdOhvwZsT+/Qmx2eGO8OuEe83ar1yWg5
rbMn33xbeuBcvi502x2tv35jzmvg4fDmUa/IjQzSj7pdUsUkrrnzJ0i2oquFZvJjTNlxSFs1mMxZ
k5dZnYnyrm3vBu1plUb7lRi1p/DL9cCaMqgeB/cc9oMbTFF4fdmWKe3bb6qViX0eeVownU9O2DF0
zy//aKK/YuOe+8GlI9piynpVeOFGY51rKn07UMKsAIRZh7A3Sr294X+PbpSBkWahZ4QN/tg4ejmN
CoTZS+pmUhUJL+jshi17th9OoeF5tr34nVHEBUlUmOfuNQFW6bpv29TKmg5R7CXevSsgFuML5Qpp
G/X1qWAq/xAGigcGaOM0nalu5kkX+Nqc4qaN6iiFZk4txRvCpeAI39MtpimCA/V9bnVIZhdqgE42
c7Az71qrtu//M+S49TatIPQRB0WEpITpoLsMnXYE70cGj0OOvtIObPxAeTK4I6AS6hTFQ/FCP+RH
RW3dbBcmaGgVFYBdc5t6InnivTwJivYXoKGLlpeElJos21duhLS8YohzTq11S4KK5PFvObCunSfW
M6yRjluGhiIC7Gtb8ux7zZQ/VsTH+lt2brKzAbN2w6CD3E3Rpwehv3lsOSbl650BvduMxKkGHcuF
5FwPQYo9XSMnBxzdIN4KvQEKgcUjud2zBTqhF0BwXGhmewCXmoaKhSfZzNWSFuFTJ4Jl4uJ5gKW6
qyi+EXE1jQx0FTrmVdmnUQZf2Twy2wA0tR1wJJ2slrEaZ6clHGluuYm4vlo1mh3R3dU+e3d9JR62
RiHLTiLBSPF6Uh62KmLZjx9IUDJrOMrtENBUeb1uaT41i4CgB9+yWOHHksZ2KLw+zn4w/Nbz5CFN
PeMq4dzbjF0/3fyqu5A478U27FDhgrzIbOoBAGRcouzLYBAzwqi58OAwMBMfLxS2DYQ+KsNojA23
hgg9yaplLlCW6YD3oEJ+ZCng1s0MXL+vaF6ZagbOYrcKlmrflPIohrkgMofmYPqySjYpMLweEczZ
TGlC0GCh906GPXy0qkv5bME7PYpNvK1Sohwl0d41E8Wo0Ch4ZSQ4ggMJwj0XdgjGi0SIIEfM/NDm
oHXkXLw3d0hDQZPK9Inta1TV7MNjS1/veEmJwIZ6PFUQSu3OxLfQfyg4a9BCwadNvw4r95gnY2ZY
7yRjVfabwVxNvQqCtA/jgXg3sYAvDz5+T6NQ3cLluKWIjN3p+6m/2nNnKP31YZ2tJo3red2UU/3c
wKlsWE5OqNoIYkh/nOemcaS5aezAmwzsl1Rj4sOEm05kA+rOVl46j+Keh+kqwXwxad24fumrX0BH
W2/cplVxN/t5Sd/ahUfVVqHBHoGnDacpEebK0n7vbPEWSFM5Wd4DuRiSPewjNZNZntqH677y5Vw/
ymBpppjPDTWTwMIeJNKxUiEQHx7/QVCqXAF9kXJCNFelIAjNncWZk1iCnLR7Dc6T9Bmio17nWEPO
MJQypS4k8Kk7/g1apxrp8xPADap8rK7HVEEgwZ5EdtHUg884vxal8/ySCiX65XfsfQlOo4bWCg9T
EoashnZLFKjeQE9N1noK+Q1mL7ZqHw6Z71mt9VAiyPI/rdphWp0eowzht1jrlA0T2lcL71gP7i3V
inHPAWISf5SxcRQV8+2e7IIAVXHeGU++z3MQZXyLlVbTZ8oeJtpqTCiQ0cMB4sAR5XoFVY4mFoMd
xvyuDwVJr+XTmbLJrLk7N+iqf7tGiGQYo5zHkgoUwSc+olmOlmkG39cCXtm53vxXTTptgh6ZX0AT
osXvoaS8mHK/cv9j1UaJIZye/qjEy5vme0mAwPaHshL+PDZI+f7brH6S8SmiYov7wnL9bSpKQenp
9vcud2IFrxZnVs1awNY+zO8ksiXI6n8+VYaYJXmCmN3Z463z/N3ktePqsrP07Jjtms65L12KUj6n
96Lxb6uamm9dC+BpdYKYyjg+dUODvQncAJ5LxWO0h0IDdSSOQSEmJfPGKkcd/PuN8HgN/sGsTCeV
78QEc6l1nkZJzgAidFo3jFK/SpmjKIAHlhox7vroOkb9sBMb00GeJB7sxHnLTMRYLa4PU0nwpJFP
7FGlmxORn1g05p8TXcjqDhDZx/1lYMK9R86VjQgh9d0F0+LPpDduSu6np2U4fc22312+4Rust+Q2
08G0iJSAEMUfEoO1lMyZww9znvfaI0ZkYXJn7R7FZ386h3t0iU/k61WxemzF28d15aJZKr+72PKH
vh+GSTKtkV52jD7D7Np9gBNQPGJ3AuRhYfndZVeUS5GkozmZsxrefXphsQ+IThz9zTNiwugN8Yb1
LA/WhquG4BOy+QhCx4UUNV1QpZxqs3PwUpAw2vRtLg/fGwK7unSjeabI7U2oAg8frMth5Jf+fcWl
rHXo5RIOiXsuFrauPPw7XQNFhHwmipgSo6jSeRqGJ4wS2W3n9CsF2nCxMcZxoG6/t+xBvhyU+9ru
DopBfndNTTJbI/YWtgaR0u0VKiH64ZamSmbitX9ICtb3YssTsef65H5zWK6RuVywZayDVGL+TdZQ
0mXbzTQwu2SNnkFJ0sgzq14/btcKNZZ1py59fsNH1IEUx/eD6KLCx9kIUM3gawWQlndBB70vl3zx
hzianHGzn2NPa2vW6pel3GvxWd+fThFNNaSO3C3RUriOw1KzSLXCyE9qcm71adbz64h+Szc+hc1Z
WAWzUsKkoEA1LfYaJinm+9/TJcApBArWnxu8yUIR2fuVd1cGyavY+sOkS2hwn9qVmJEE4fyzd+jt
cIZDJNUrDqpb4qZjmQlHIFQbSrLmF/bz0CyEouExclWHuWjJssHGKiHT8EwN5sIO/r+RU2lPrM0y
iawuvYz6qd0744mCDjElUVJ9tJ+s8D82/5vCo7OVkLO7j1kfHBBHfwxCR45eDm4qSLA4AOpI9C7i
itpZRw9Syx1zjJKC8vEyCXNU8gLZFivV5t6Iw72MM2hhb8hPpmeYsNtUpS079xDmFrNeP2Ww6spB
/EuAc9kHa+9Z2tTp4kKmAzIFPZG/ZBKv+U7JTXQ6nf7gs/ScBI4mkHhmIUrr68sR9XYt9QZ75CHT
5XvEa7FUGhlsHevYk0sAW4pQNtAdAIFBC7Y/dhTvmDv2g4oVY/v/7J/v1+0seWu7/mM7fPI4CzsA
c2At3NL11WutLepGohRvq0ChR9FXrqvA2qPDNGJtTHQEfEkrYqyzEa+v4JwMAZfFY0507yVByTW7
LPziPp2SvC8LPqvKP4Yk16P+ieRXOuXqs3QeU4E+ODXwR7dS7dt9/B/LXlB9OvSlXFUL8WjWzHnL
0T3Gi91PZDTG1XLEgiElQeac8Mjx7ZIFoF6p0TDpKy6uYkvAcU57/VnAknXMCR+rgv8aJHLrg3Ei
8zmHvr71dVhBFAfwGEpqoDfj+mX3s63zgg0+xyOoLJmhcrMbfV+nslJ5c0RynuMflln6iR0kxvHr
DffFM7jGPuLRF++6xAvfUVyo/njrSBwmzvbrJlMRv43ljLGDaV7E0XwG3kUOXDjob1Kkv/gFcnfb
GJe1vGHSA0pNIOOFdW1MKOqimk1mAyCEVMDBYR3lj3ytJ3LP7Y51hLyRqwpGcEfjZ3cflx+pg4zR
AZWol54ASC6cPj2p9zAlwqTZ/+JW6xD0tVniI6xYwCuwbJ8Big9reGvqFPsCAmGd3y8Zc9Zfvtf8
FCSaNX0cgBSZyXKWcHx/rHxV0bAHIovnvif01QC22oVV4t1H2M0bJRCl87jjTaegttrm0F0m/cxP
Sx8fqn1rsMWNhNWSbD4z8F15/a+KFfuM7LnRK1sNSIe1sm5rLylRs9deJmgC3eN3cBSNSaUOPUsU
batpHN+TlnCyAKVzmsAjfyr7DzvJxIaR4aATT/CT7ikq+QhJ75mgDLCBBQA+yod2AF75ZWQDkc8Z
4cDPiD7RlKA5POiJ/MRspTrwtdW7w/kFzGzsS7tjR+cFWhE7Zf1EPTA6YOgM2QA6rv7qCdn1qQe3
9tl2r+yK6kSHbsP7HfrpEYUd5NgW9vPrziEUrEzp/IEwTPucwhdBI0pUALZys/ICVqIEqoxbDS7r
kCsefzrtMVOKSyNYCvENlUgdIh9xAbZpFZNbEtSH19AqON/icY2nrqPLwAONsbziz796V+24HxqU
zhdDejTqThZCmXHvwXcIM0v+MH9htMi7VWRu+V94LdnGOT2D9z9SdnJF+xJ5V+6fRjqxYOMfy3pz
2k5HnaqG2ZQjQlAWXvtMWhBLpkxuwI0uVDMrt5f8/0bz7eoFn+Hh1W4uXvP31xVburF4l0hMHc7i
Uq9tDi4E096hJu/Mi/4ug2L1EpVyXaR6J22one/lXkP/QL2pHmBoD3Hlt+88Ko9ueQr6BbRDAwmY
NItz4N1OiUbcLGvexS16X8b9XwWmOeZn3E69vtcQCtIMSGITGyXFJm2az0GWAlzAQRNE8BaXupyz
hRMR+KGGKaX8AKxWlHZLDes62JloVnC/OkLRL0RDLtUsJ0+tJH+U8j/eHT/+EFd6OJ7lg4dAtoQw
Kd8m44y3AyMqZc4CKsKFEX2bfhtlCt0QaF+nBURkZauvYy4oXoDcxAHyFyTZyBlsXbf69cp5FKaX
qt6K3KQhJAUBVX/UrSiHANuHxz3JkHtfyA8826FH+A32gCmZSbowUJGV/FnfgADw+DnFH0fdHPbk
HF3sCG5Ri8wnWefsBFojBezdXisqR7KX7CZ21erX904G5mmW8/NOA4O13RRrgU3ikVQ5EViCT0Xn
sZ+3Mk1OGunrngXksg7iJtnTZk1y/wYN1enqtu8bL0PlTj8l8UROboNBDe2ddENlNqOoyghgAs9G
35EqT6Zw0FgdlcrAcF9DFxXCbkrBdm+jtLWFQU1QieR4ZuE5OsitOeozTdQ5Ta96RbSHdzFHZPYh
h8nTYGEx+3lz+P928bkrZyEQcpzmoRI8FqaZxfVmawGUCfsphdbGkkq4oDhBi448eM1L7XdBdL8f
+434Q3txnT214oTVDm2mNxQwN0LtUW+GXFaBMXWtC1EDUjrSmgJwawOu8gbAGz6nXhTyeHXuV0BN
7datteh8vA6zR+5afHur2JRUUvt6k2SS4cyJv7x2nctI/ZSs5KcmlTNv4OrUZl1GaVDYF+YDnPuL
uNsSWwEY7tZoOXGhxnryMErJl8/K28mQcZCj7s1udc/l2hkSywLeoCWpZy4m+xxlZGl7xQxZi3+R
5FVJTBNs4qxu1GnE6Yit2grM6EWaVWalmkg4glnShI3gcAvLqHBE0KFXKITp5WGJ2rPIPZ98YTG8
3xAG/e39Mu76mkB2azRlbn2X4AMzUEC2+0B9ZbuZaxCgK/pOttzfylVOEgUqPKSpAZ1ud3of5nAR
VHTL0/VfCX7xzfi0OZdUn8mP2SPAe3jplQhzgql0O2uc7mnk9HzhZnjNc4H6ithmlU0KlMhfqJ8u
0Jk47Jr9AXcdMmb5JyPbHOomdwvJGLkMEt0EWABf0u2z3nWUe9528uvgV2Xf2tIIofSyijbHqKVQ
15fAhKT0hkRgTGVOJvlGNqM6a/PtYi1BXRb7Eu2SDDAmpFtF+tjJVnkg7gv2BvvaS8/u/P4Kqudo
TnLpZ6NSXO5H1efHAv0K9YhUzMcpV/Y0PO9Aup19bvRo27qMsEjHdMX8QuSNCXd4lcIWqpc7Ap6J
i5xTWzUcpDFOk4UhTbI+6P8IWJNq24ArQR2C4oOCgf0dYceczWIjV4vedhVFM+7lxIoOCOHKpaC4
Irx0WnXfZX+1eOIUsamMz8SV/IcFksYYY5UjcJkd0ONgIoNC0iH+/KeisOK6FfBv8lEECbQ4TG1h
RuOTlX2JBkzsXCRlVJyBGsvbnNKqJq6vNbQJMBYgEC/NbPPa6Tr4hWKLYUybxBtcUhsO/lFE3h66
YKgEdfoIVaoIQ3F4yAkqMD7P5jRuneyDuGLUSFEr2QBaXRenhFwBCxdXIx7UM4D5CLFPOEho2/wg
NA/eMilKa3dMCic40SYjY1OZwHdFNuJDT9kPjH00XXsgfMHFhJ12os9jmRlCdLtzdJh+Kmkg6nlx
gAo2t9RrZbQ23T89+dLm6tYLbxU/yBl3jUxdc37/q96Jiq62ZShTjUNKuLPJuPWzk3Py/WJ1GVdT
wLoabPRGXrFkzm595+yjzCTXDP/6x8InQ3OwIg85qmckcJVyav5i9OxK23ChaqADSPuSW7syDKA5
dDVvLNPoOvaKS76CkOqXycqC/jA5ZlJuVsQMQnj861UrXc1lD/HijLplovccu5oggkmH5eea+TdD
fDgwkXZeIzSTvPNihaql+aiWQ42s2GxmbLvS4TLl4wlAGulbw6EEeQguIt9Qhu9Rf8K+4B4fOdEF
fe2UlKXSLLFaFGKOO3nfxjCyogqJD7DGIv2HU+6H9ZenjEY7zEUqe5iXlxXWTUgDwhbAt2W2MMLl
KU3XfI8BeySr3KFJaQuzO/J24eavh9T89ukokvxSLTJk+3dNItB8vWkoOK2YlwU4ByPAlL3XWIIc
EIuHpvs4Yt8j19o74N3L95/9bT9FMljwAke5glHx91G4lzDWt08UZgh3D9c/Uq51FZ7VcB8ZHNOb
BasjV0fJi9ZNg9ItlHJpsKjZRTbMJSUU02R5PDd8vKCQs3s1NHrXbaoHWDTID9OERaotXQEszqMq
D85Kje01WlOQ8qfL/reR+ODtSZL7YBHbU3YJlZIKF3A/FcUdLkf6HVlPuUZ7cK8zfiD+ynD9Y7cN
sidVKZf3/cxTrZKAc810Vkp9RrvYKQDbKFtO4JhbWtNvrYnJ6kUr0K+VMt6rkeETPEwFbTQ9n1vS
eSegdI33YhNCt6lhkBXDLWlIEATjNTgHUOZ9mHVc3WLjv6awKxGNjYkR4gGA6L4x/AqCgyPimgfz
iBjOKTnlofs7++ogqsFJEQCAyNux+AYYn1LJOLawed+eUBZIibNFYb091JpUs4FKBMwfU/EI1tzp
b9WRLgPNb2AyFILxxDP1iDc9cuxVfh5Dsjh0U09/RZjezQ9aD+Jg6y6TrQRpi70LTJK2hwyNPPaq
zpRMKaR6EUevKS6zt+T7sRBkIH8gqyrOWjl1gtrSVbO8D9CPNO7dN5MPjj56H8YNQWYgXlRzaSXo
leSOvCX0ByfEmo7Rcz6dlRWE9R0lNjNW7zbklo36Wst9C48sJKWFPk2bk/viTl1ZTNYMroKnkLbb
/4IJjUgLx4OhVYiQtB5YHFLDN/qTdnsa9YaVq5Zu0sIYAHMw7olEMASySXk7tB5VXT4NZx/tVJnz
UJzy5m83qCo4AT4VAnz8NP1RSGAzXHJyya3zlkuKaBgAITrJ+rchI4N7HRwz9eMK4BZuIYujgi8s
0pIgG3ZkUNEjprCz7z0MazY5VHG7vaPb+I2aAI5n19K/0c1MqEcNLRS+wOk86izfEVPYRQx0XqKu
JVfzoQEamrLW/KYBLqrfBraYwbfI9HpRbWFlFWSyCt4AZwdnMG9Uvxy12ExsWKk1cjZVROx8Ia55
gLE0Sz4685KYZ6QEQodGirzzZAXz+F1t4FUTU39iCl6OoVFScAUH6B3B3qOz1okCqvTRsDXeXe4o
X+nwexjBg5CNNgPs0fEMnG6io0D/Q9uQ61serG1wBjOcEAaG9WVovBAHvtjCZ2a19QBB18VDS52R
+r7oiMcVW/DxY0LmqbxWKH/PWkVVP6WN8ueeHy00lYSiKYnQsRiEDYzRj1Caia3cX2l7xBaWC2Tv
pS0Tr1FoMnkZYZGeOU9o3zeWHatDPMHVUJXoDbOlTlLjAtQA+EM4SXfseoyiOrfEOrADjLa7jOS1
2ydTCVXKHp/+jdwSxU1/wQ4jdx7XxM2dKiglLfUGhdLz1gJmN6E75xOjZM6d+8iRb9F+/UXwSVJV
n+dcPeWko3YH6VhGJQjKZiBBomxjc8fRu9I93CZT1yUAb6V5rL7RGj7+r0lJ5Ua47ImmlIo02DSA
XiWQnU1gYilbiwckEKdcsEPCybxXRem2NlmOt3w4qtivJzBXTK3NgERFlrPlxHN50MecVWySaXXA
teytx1w4RFt7YRRt1fYxugsjw0u4l+ElK2DRtsyVdKrZuF6nbZIGycWubkyXpfDIe/7f1/IsyVxO
cx+LCayl2hIhy8rMSF6H5endL8URponb/MM+8/O7ER3ZMZ5mBmcRlKnw+T6fcmH/dKw2EGmqzc+c
6C674qGUQP68IDRQNp2Rwi65RULMYLSV3xaa8AZ3PKBnV40OFD0/vrZJgBSgugkBOCRoPb4NRtbc
RQ7tlEi0QpOTCJP+lcSx2BORhguT8lzaOK2CZNeaCAeJUAXE1XdE3Qo+VVl7qYH83bDUmRsF8wTk
F9Yq2cp+0h6Gcbw9Un+T2rbw5Wr8BCgiSeo9nGFAECVWcddraIo7xuifY4B5j7BU3uV2wuXdiwT/
2LYchJDMEXgEyYsJaKxLh7rRdfl+yHwGGEEkCipuhA9jYbCHeOnPy20UVKeB6PaS0xTWZ6XzWL53
on+RJ3usDChonwZcctDBV934BeEYT+dX/KzkvJkx+uRb5T29sIscgj0K9EMi8tHri+PCOQXXNYRW
W1e6illKM3OJZb4uj2cPkur51ytOXe+8omAjy0Tx6n9qMwDuMJXzoZ1BfCAnf2wWrorzTmv3IM5d
2PXlZKOxo6eMqZZzwHcVT/v5B5R6kNsO+UPdbKulLn+Wv16cb3eIqqkDYEwyKYnVCd8rNWCAWAZr
79QtQmiC1Dq2e27gEcd9KBYJbu0qUoDvSrjXJCAoJd4Q4bf86Cp3k8gXlaHj9aI5RvmRXi94lgjb
Z+gBcNkP7D/zQWqyEnxnuSbDonkSwXc0JzHDUqiHMDULAgDNv5Y21wrJAzDuR2CN+q3WdIKYIRs7
sLDE8ql/7sFlXjNnhXSuHXT2R5V/+VNuXnG7v5NKAxyVobkPyK4pZ8xsEkZNH7Mmu5OIBhMS0aee
XVbuFg4+sWnmcQHyATeRnn9ty7yGWposXBjsW/UtwuBFuAVylop6dgss2yNnIFskD2IdW2I2lLXP
8Uaf6gUyUacTrMyQiEEz/WbMJyaqdxvo16DQ0/EYrY1ZBmtOoxbNuE+lWMuDtd1pAcDdGmHYUMwr
JbOcLRVk05GJIaR7Ux5teqrdW/ARDjpfnCoDAVjUNPpbaPMLujzgW3OYYhoP92QMwi/jv9zThNdN
v4JQCWtcXI8keMD0NipkbphY3L+kwNKhkBCcSvejf8I+1tTcrr8SZXBENXXhFq9IUng33GM0i0+Y
/CKPeQl0I1qisltv0C59cIiPJKVmDgYazNJdXIGHanfQmYCeXJQJPwedo6cah+1e3V4lmPTp3ncy
6gxm5wWQZMOnmkKywf9Uyqk6VKtGTFTtFhYQJ7VXMHsu7qytURLbvgo3ifJvXx1OO4TTg86zaPSu
/pLmxqN+542IZSpYkw9RHHOumuo75KuvjtcCRTFvhychjMX0KbWaAWHpkVxM7cRknjGrgdJrsUDh
qZWsAKJhxJfky5h5UoNl9BoZZM6Mk2HYC/qXRqtG3B0MLDJJ+/8STgJIaGPYPAvr5MT9TVSF8Yft
2KJchDqQy8RUN3mynbR8IG235CkW7C7r6LnYulzDIUGsfJql9Z7+jqILwSwFC9tZ+zwbnU5GNnGK
etNyfxzvuFdfdZaunQSYo4sCKbRU9CMDsrctTuhGVhvEvIw1c4JVS8e6oiekq+7ZMiXZc0mPKODY
t0Uy0fe+IhJGcFPG/k/idOELJX0PihX1aImCMaez8sj7c9C13RPqi0KL4QqEDRD/mEp0MMVrKAJk
/l0hgVwgESjAjxa32+02Qu84UpLX9iaO5BgFcFL5hNQTeCyxZev1VSQ/oNlBHRfFvaG/i7jMme9i
LyWOb5npj1mrSkXdCCcEpodeHvNVFqW9Qudb54qfEjNHwcSqNbPANeXmfo21JdCMKrEYB1BEEXiT
8exRfPuXGZpC4yejaPSlSekzUgUo5kOdimjnEgmer+gx9c5w/ll9XuTUEYqbwM+kH78/H7AnHKiE
+eJ5P+AOlpfMLtVWS5ibLvS4cwn+5YBW8C92WX0ea7LwoNdTpF7KykEdowUFUqsela3Xvi7cubkM
3bkdwaJxeJiakc0H9Nnz9igg5EfBKBdMywqU6dKOjfpk+R/epKow/GzRib0X2dujhQtHbDTwI8qA
oOCG9Yutzqn/FUZfHhc9D1zmZFl0Cog3gj9FQyo+U5OyXODCBrNJyiXpaje/8iTj5s5OvaMTC9fF
Oh+ddz2q3gXXDhrPCEDM/CAcIopBOJKdTYqd+E1Hhl8scwpcu0gm1d4eJZATQ1z0saW5VWioikF/
KqAc+S0cWjKdX5hCr71ASKtHRa/Nvr1hTW0mG+pEd66cjOkMQx2Q7jBxVCRP3+qOeAxvW04pJab6
T6pV/S9DSlFBrCibhJcv70peas6iH+oAjMeB10xewTlFico2SuWMRH2jPz8utW/MbZqNWqxYJcAv
DfZUEI8jE2HcfKkeH0+6BRjpqnhz+GgJkSgD9rxkkDgWaPwV5EPwKyFLvK5TuYuEL4zKaVDSGohI
2tyAqOYAEwAXO22px+F7X8rbUN9sBQI+Wt9RwjFj+OeGNEAWmXuAXndOK/9td8cdJ/YjaG4YiAin
rEv1kCRFcGbNsygrBlXvQAnmyWTl4fZD+m35VucSVXXlVBn/dBvca1v+g3O+/zWp/jou+p/ygiLr
SmU7NKU2Bzd7pLEisNkG9b5tILlGIbMlpjO1PJ7NAAmOBA2+L43S0VhU1yw3QHtUdgSIII6d4PGF
qfdBUIwr1tHK33AbbrYLX7aEMFd1/vw7qB70BDkvPmM9R+jT4U/lh0k9gB0mPAau92EHq2o6jysG
Mvs2SlfUbp0H6pymFTzcroN9fOnvjRDvXCiczaxcJg29xivGrYYp8We/SdfRECoQEpEncoowYhgU
JikZ3rKmRK3tQgSz8mLlDIzbrRx0frcaBaX+P9izvK1EVTOBS0OIE20yycHICYunY03OGysw70tI
pOuFJL+Ujh/c7yMom07MBBm9F6naxYrvyOD8BdmTc63oxbq4nqjYle1NW55vJEFkmI0PKDyYrkbH
jpqDzjR57qFK0X6pPEBERznEwBJe9XpEZNMEXiB8Rua9M9npV03CiKFtJ8gyqWDtosBanr3GVKhi
5PTlDcUlPuQCjt7/EGIBcjpFO8wxaziEDDqb/GOsrkPazBBVacociUgcc+Ok5UkPaxtDFvHp4eRb
j4B9+rrUJOaj3HK3Ov1ERwRKOGHka5OF6ixGNyoXs3GRIOGtFRPVwBww7AFLpxu8sEe0Cgi3gX4K
M+Tor4VR9rvIsRohxPRec6NUcjzt/Mt+uoQIL5YUsTLQ6LfkNXvxTGTSM4vtjT/GeuMoP8uxH3ak
gHbreQAA+dsbGutk4PnsDk9JglOcVm778Nf/GLPmRYCOOIbVj6i/pFOghWAb1Nhoq72bCA41sBMI
XlWOHVjN/UvoNOYvbfH6/zJxvQdZJiE7POLTce4ZQhlH/beeaLZMzMPlC+FiCQwrxx+HtjLWObWs
9Ns9YMvWVrqiGEdWXFDThRzddVmPFFxY6SUV0zxGzyZGJD8GkP16nuvMx5pZSUPKRgEVhQWH01zB
fZltuFXp+BW+nHItlt1umHur8NOLfxDM1oj7GA6oSgIuCT7jrnfIJ+mEu2dnWrjDkL69CLt+obXc
QN7MKrUlrmHcslCrw7dDYHr7UIqvh8DaEB1PGEdNXI66uh5FRN9gIskfC0kLrAABFejPVHMbNPEL
56UH7CmM/nRrkFfRV6EgVr6HjlBfZii5t8BqWZVp8J9Hha2W7koJfvHwHZ83GZP1k+I5pSPc1k8e
7cxvT1rPRZY0o9XZM4u5nKHkuR9v9q7nrD6wGQ4z9+cKAFOgTi2dU0ThdiU8Pjw8Apgqz4NYVgqy
grWbZZRTEs4Njqww7C83bpHtJ4hdeizs1V9Lo0456ezNC6VVcwkCuvOyjh1vb/Dg9Ne2z9k+2lct
rwwusFwi87cgcgWTBQzvxMqFvoXIanMY2GJ4pil/vVcALhygh+uBqggilpRQ3OgJxiAvCzR2SxNg
z0HFC+E9VKr7J5drq1VSWYt4QLaX8F2bA1A6CULu7a+FSMfGewFpjge7jtekCnuYjyShF3JLMpge
M5ifzxCn1oUjoTAqOTnIMj9SuOekD+ZVzZllyQoNUv/Bs4daPJp+A+JnfRUS/3UjZBzuXHpeQX+u
H4LPzqtnidzbWijXOg5z83lXBOI8LE2n8/mO/dk/zO6BZPvGde1B10fAsOIShwS1AjnRWTLuHShg
kmKEAFD+JYmRRO/SFQcbDZM6PXKoJOSTZOI0gmm/KjOYypk1wk/WKv/pv1ktAPxxv2zn4dm+S98P
HMSikbGp6EGFnZVG3EnaE22yavcESY467EVQC2JWs9yX7PbhZmmzM6H1kt1nQoCEsWnUAMaq6VFe
9YIelYKW26/hMZtLot1rWbc/wdxRU2hPlx7GVs5fYz5CsKRr5aOe4Gl7YqtNQRz7pi1nA47vzFdl
15eeh8ZKDv7Vx5cRUROk3ZD2CsR+Js0DFv1CXbUPYUnzgQoXIiyx9CCV7fOWyJ1ajRKVWNHjEbcY
2sRWOzTAHnkE/eZAxbZyexizcARCm4yOFXwyhMCNPj6T970lZz71rFnPfo5pTPjWKdbq51SWIrC3
2OvIMYs/s6SFGyKF1eJ47k9JP8netedQnIfVyDNQ7ajj7nFzYdGDCueG8uz/wGvmeKStiHJbKV1w
WE9zzbNZdqLWEmXjHc9WpLp+e1yYrrqzW2qcoqbAJUHujb05Zbm3vvBbkuWXrfGnM9cWw4V9I4cq
l5SfJyg1vGbP5w141uhRoqNxVSPGkfYYBE7yrrCFOVhjmtposBC+urby/FST8Xt4OuK7FAxN305D
xg0MwR3cx0dnmB4S5ruJrSc59RctaZIAm8ODRbX/oCvcWHMSUfwG9f8XiFcigEA3YKSwNDSlexP9
uUzSvbcTgqV0GwNFvwQKX91EyRZfVERXmCSOWQ8p+1iOgCCn0Ji1jyEwOA80EtMBoMNAG8FzOwU9
LHl/suOs/GnBPER5RBLVSFYlO3rInHVqu96dTDORMldEHsHz0YrVwYSXejjddv1qFwuOHlQ5Yepj
L6jqqE38uhC8I1efFjNBjQF9ZE7oCq3I3dM48/QY5fXGQ829y5uP/QYYgatFTUlP/bNrJf6KI3fB
HtYo8POt2wMEsPhj3liLutdAeDZ3I9hKk8xCE3kK5Bx+7ojZm+SVTXpe1KR/ai2DPnxU6FLxB2j4
xJYZWuEJIuS3JYci4vHHn+dPfgFjIVJZTo6SwoVOfcOpCWq0c2QGgyke8k8IPu2bnHeBiM8fH6TL
dFrWaSeard+JLLzLPwitlXX6QjMqE+6CPCWlp2h4B5jd/e4brl0/C5kAGnl4oQ3p0ZW0EY+hFuhP
w3ADiNPl+ZWG9BMtg2RscCgWllNxYv+L/cqdBeC97qqhbyXr8661Z47qVfubRuDrhnSl37b30b/V
qE66mUnXJPHaG4/GraatBnRqqi5UW8b9OT3eO2YP+3cExlATylJUyGWM1rTsMzCCYMd+gPX4YpTh
EbZS/bJknyB7RSXUG55QMaObKyR9HcB7/Qcxo7NjkRcbfJfW5DBBm2hXPsBtsK6ONvQYLzsuCsyV
M+yZKkstHZJ7PUAluoJx5f7FEVjB4KO0fBgymxQoJkRs/6aJoWsFm+rOYtzOoQFgAimj+323ghUB
Sfh2rv/71YYMxbe5Gxkbbvj2oD4dwqzkHj5DK2Zi1BaznTWTtgL8xLWZ0aZMVVzHXD7726endNHd
d4w9B0cKOHucfBfEDQMTEbpoAbIj/FZ42BNJC74ihdC04oxDPboNXasC3jRdjiwdN4Ze3zjOUrwT
XqG37im3rPX6qKKQZOZHZWcvBMrAauOpfS3/y8Hwp+DwHaqIZIeuooLYb273lXHnsdAY/AbG4mYu
Pnh/1hG9fuRHltY1REq9iiC+XGVdvuW1RaG6ZPskFY50/NS24AViwUPw46IBM6cQDETpST+iDMqk
om4egmqczCAlbnMx9MP1slV/H2hnUNZOFyexhNW3jnXJDUKksRJk8kg6cIXFnRU1Pvj2foSWSW2c
NBNAfbfgU8jABiQI2XBRedYauFtJW+r4V2wmNBEIJDHgPBq6qd3oR5rU23cITOEeCKW419AjBQUV
gE2rmzlDI/LQnmakiyxi+lnvtVSrxmGuHIQY6sJzSMouiYmdpsBQUzvgod0J7scLCTCdnrQ836tp
0YFD99xn/cHS8WN9XWb3chNqP78cYBcN7Gk6kFFnK6t5Q/E/Sxk5fexP/QdWIpQk3g4loS3TGfpB
AgVv2pIOEzqex7cDFJCKr7w8Xvlj/BSVzkPnFTuPWbZh9sJXWAb6tSPNL4xweCl298oN5V/8lzCe
S+vJPqbRfHGJjH9zD/09ZM8JKQ9OyFi4+uhYW6/T8lAujWW3kIZz64WJrHT9U+bmstkX+IV0ApD/
HcmmKz3+Q+cqRvmfBo3Tm8Qv8SLE4/Q4JnYsRPRQC2CZF1Bw5nFd/+66AsIu7MT4Lvp1Qprzkc6w
DykLwpOFgoKJ9+o+6Tvnjnwc+bVhInFnEZzIqk+rrzgYatT+cM3UG4rZuIfAD3NxXdyZCf457cN5
38HO4BOGG8I/5Mp2m8aYSO3wauUhHyWZ1gzwXgvCD+5vxeN6240YNqdsdt0zRKzZBARvm13dIYXL
HMEPp1G1EKI8vMcGWgR9OzwXYedrCIBCAHAqw0cPVyuaWjQfnyEWZ1bGf+QP6sRrWPQdtDwmwTdT
AH0amR0hpkP4qEjDkqkzViJS6QQzFTA5CcBR+ooIpM5k36xXz9XZN1FqLaQ3mQq0rdhMOFk1jyLF
59KhwOt95d5vLm0fKDwFGfsKKQcVlDPR3dapaJknrAAqJV4XdWKHRsxWIma4G5bWMFZCpOjxWdqh
wBUb9X4xY+yGOrd73AxRULV47a3KUoqZsVfLDp8S3LpRs+eSGWXSVwFlvqBOkdKaWOndcD6gYILo
l31d/F8VBfK/zCQ8FttNQjIUWiI+RNLv6joEaKD8lysDLRxSt2jPdcq1jz2bKj5U5roWQvxSzbDo
SsSc7YPq3JY9iolf9mqNdZ86Civc4h7Wykr1vPBzr9toPW7bniO24Kq4kjvubHozK/RxLw6DmNaT
yvt+0oPgE1Qi2eVOPwJUn9weODhxuP19ER61oemD3wH5EcdmpCDUcJOsv61KtnQ8TSp2n8BhrVx0
fdfrAaatOm8yaUFSUosJLq+XTEXR7gj3BYH7u7YHD/EDJZOhINkHAOz2iJLG0ooucLdS78VtV0AJ
ipaa2RvCaw7MG2xpmXrAH0HvhG7gw55EyUk+wzmNen0avNa76KNyAKyRKN8cifENHPPnf7MRDBNE
R0hi99UjoCF4dhScCGI8dGt7WXCZnKb3O8hOC4Hw+lXb9jaogJgBb5whAX05njkuUQPKya2buVHA
lpn7x6PN66PVP/ae0472rhLzYeLVwVGxI9YEeMw78Gn/2OWTnAlrj1nS2Z472KSl3wtF8lhUcn4G
UunEYnjKf92laiwA4oRQynh+u5Wnctu1LAhRHkftSMYyj79Uj9zgPuFsgi1cy8WxZd1rcxqW5IeI
ChEQKwuJSV0KTfB76a+eacGkqfwY9FXA9hl18dQ71qe3gBxGxu0XZF1rV85dGh/cjPmYOZCr5qns
wy3ohvnHoWODvpGb9EuoWvdq5obW2ybxT6CsvppsvfaVSueI1v8hWN5NhlXsh56kVKbYufXaYzxG
A8lNmy0lI0moOy+tTO4L6xAeNNxlvUk1fvMIm74Z0ZqBU93hvw5zugLg7AAbmSJKCqTUNdvWBIVk
Lns/8pI0h0m1hnRDXFjprgRD8FEp5BhpP5Ruy9BZKuL4q4k+zrZZrCjA4c533GZSHQhyKGkpVz/O
BbomaM9DGXEufrEWbOH7sUvNoskesAjA60gaGpkGoMMcE2Oa0+0IhNjhEmRSp+vLruSWzXCm4lU/
+wmfixebqW9gJpT9gQflMG2TN0RVVEEsJAJD/L4Z7W152GzWd7M/Y33Np+5U11MaP4TNtdi+47Wy
xWQJf88xJ4iHOHKCHoD/hDhiJ7o7kIX4SN0Uu8aW3r69EFIzBBfH9l/9d8O3WYgY746JLVCWtViX
eYlSDDZ6iYGeRjZgDnZYLRbwr8YpfBJE4mfdH1ZesgAndgfx+BvKwpgsCVB37nRus0xbLrmEiB8w
rN2bsfctCsGZP1U2VuKUQ+9BIzXWzV6II2IEOX6TZzib+HQ112s1ZsCHxPbmEx4+GVaJlpoDLXtb
MkASv8Oz8PvHO4J2bulBNuuiOMJTjhGDMv+aObLCU5SiC1zaSQOoql3Kn2v/jmL1cWp/4mZXilAC
vLFdkHVykh26HITu8Y3bvKH4ZBQqHJwoGiFk1qFz3Xy+qFhVrK0bUvWRy0oWORSR4X5DXPxO6P7v
po4TZ4V6Ee42M6NoLFrEMwtl0sCpTXNpSJosLgaph9g7rtDpnPNoAfKsfzteYc5XpnvIJSrA2be+
8bJ/KkezduuEs3XfXjQ+QBwaUSgJgOrNL5VlTgD+A57ltaHG7Jgv5q9I2khS4mcmn4/ezN18FpBQ
8f0GBjb+dYFadWszXLXIoWoMYbxZJroXmlhNf8kXZahil2OLwqLW5khvZ0l8VoGHot35i8e9D4cZ
y6R5q0bDmFvVYM+4r1iv2xf8cbz05/gtyS2clHnp+nIkFEtIS3qd/T+cyjiJEutaIqy7t5/4HllJ
3DbUA/LeNZ/PQwKzCxr+bDjT6VsLpCCJfVmhsZoz/IrRebv91iDOhgr/p3mwZDEgFYcLZmOE2T2R
jcSLN8/p2I563XFIavcFXzUKlfaHcqHH9XJNFwLzKwamN0VBVnb99h87c8K7Ir63QorspHgscLKQ
OlnAWH2lqN0HxzI4SUKRJaHg/vwnsh2WiYptEkGPtXLpfTxe6iHRfnZ1Jq079RP6nLEUAevns+cG
3JsFOHf1l/ZTBRtToQrOnXSX82ovBL4D6nfNre1SGAzqkJJHGoSqEIMyNb19DinQbE82Hr4+ZYxa
aSNmAoS6JOuwTehoXvvkdTM43onvB8e2ViJsZr2N6zGHrGNTvUYR+HQ/hTS6hIaZBukC2HxblcI7
z9w4rONILqpV3V2gKm7OUexOCypzVFm7fivWi7uQNE0Yb9p6RodHBR45s8cF9dj6m17jDG4nY29k
RWLsssmbDohcOiRldIImmpGiNiWqJk3VXnwLDE5zuxrXh/MCYrayZ/egszJBfL9tqCIzgPSuEKpm
DJ1pvK7r7bdtkxqzXjajB6sTJ+aghS9C+2WCPIkPTMHWwMoKO8668X/qHfQUMmnTrgcg97g7vDbD
NNXawTQW/kIZYELGcU9dXWP0ZG2klMcOy4JUf9mqwv4g2knxsxE4FxmbXL2KIICDZkPWp61K303D
6bJP+bzgMvSnh5LqBBMVa523UTsh2XEUoiVY9tZyeRW3i5suQZ02usaVXqdVT8wIw+hGMMcYNBeu
pNIFzR/bU5LGLJNHjGnSCkumDdQc7/kfiJtJA7tPVufy+Y3a6D2DuBRXvLMil6yo3gALkHkQLa21
YdAzdAWIZA0YEEGMQbs23XzglYLeWO8MTfrr56ruimRlTMMvOdp8VWeT1gcuMSzLO7bk5UO5TkXR
JeOaRnylVNpfh/WWnSe5/L6nmMkTjMyK4vYxL6boKyF66qkq3XhsZ249fzf5bh7BuyU7l5NU2+Bu
odcne4AgZGqRdb1vEU27Rt03bbLSIfIDT0GeztghzffcFjwhB/tovwwYwBTlSjfOtT8t0thyRkJ/
uo3tJJErBnsnuwLHIZn2/VrODpgGLNm96KQg/9vz0ud4Y2PYhyJQ0dr0zkixfiXMixLpJ0CVIXVE
w8NLYQ7pgopvZPythhgY8shOZmPu9d1LpyT+msvITLNuFK3nvxaXC7ogUtElSsYOA98i0tiqMyxW
OeB/ckYuGdv3ROnqV2EkySPnGlmpdVV0xIKqvNqspedLxKvA+w+vNNjlpZUkhyHfX7gnE6yp5+VJ
dnHaTgiJ1gabgOs8KvC0i7t2c+pTRWFkLFci2RqLzJEVFrkpTw90EH56KLVm/EC3Vq3fxg397n0i
70gRbdzKH/TK/t0vVWkfGGU0hn8PM7n0HFrQsQ1NJLwuAs/farRx3sJ59QUmz3JpvXaD9cuPqvpS
uyOqt0c+eJnSYfQ3A37nXa4JC2uyS9M33T+E16d+Lqr9zhMP/8KKOYJGBqbXjeeA25yx7kV2aHLZ
1NFzSpJ4jGJTTtnV2A7uk/nhM6xGFo+trFeMLfk7zlsJt32NLAQPuSweAPA/PtiWjFAOpW2Kssce
3rnhrThTVitNO9EcC44z+RwCPSLMqiAkav+DeDJLuGrfy9lRzMBSg7PPRx/Ti8qGgDQspxmYdbxN
/m7pGGY+u0DZaKZ+EP7xht7fpxdFeErqrhhg6QDOTmIZHkrLIMfzOydtlOrXEf9esmaaHYcGSgM9
TjgEMuxYgJRJSUi5nNZ3TOY6HXEK1HV7i5j6Y69rsxEXyqh30XNAJhGlN2ZOXrtMTEpJIK3a24bu
mrhgebzd2yTDYLnII4cJaAeEj4FaYSyE1FDQUEsfIBh9XQlRu5aX69xtdNqxDINYIpF4k574OjWZ
NeYGwu1vSs/DvcKXujdy7KgH3VPdgATREgpPXryfBgKulYpWcyW6mioTawfhE964IMZ8RCAZiAfF
Dwg/3PA3ND0PaRtRgWceTQfzCi7dnutvUNb65bxxM0KPWlFCYv1gSkZxE5l7DuLU0SjHifaFfzrN
pYlt7fpkFjEJ7kfZqTRcyN3uZZEPYdwwKiSig6avZ3QEUCkEfMFiqQWcBgHwDpGFNqhZBnVA8FX2
2dbdcs/Gd4IxbLpXJ3qYvYkwiojXDhTzKIB1DxWb53PGlDkJ0nCBKgW3UP+JiEsGYBC7mR05Iskq
mBP0qL7D+9OUlkkpuzQSYSSjsL4H08tZgSFx6t9PRnVtCoJG/6KPrklvY5k16qDiHu6XBBoyO/Jf
7IqwNYRsQ4g2ylibyOIj8PDN+Zy44sfFk6ia9e3bxlhpbQcK4hrzMqAWUaJE7UqYpQRjq85qhHzh
vM+uxOqqjaG1c2M5HbZik6tkTLmHLAoo5lh5N4PoIkFfkgE2XiyVn7X2t9Gt3D394ir6+pN90tSi
e4joDqoLfPRfYvt8C2seepO/egVKWNV8NZVwPg73+G+0tuQrmtJK1s8VCREhUoNzcoo+Vc17mlnz
ougnfmFTZJFjQxrMrq+CawpnJAc4Ilwnd4lTZ1IB/zY9Kw3aFnsE/SxRMuHHtHJ5VTeyGKgKt4HJ
56hYxNyAPLsrWu25mssMbKgvWeFgbNvrT2STH/xyNt7CCyyXqH7/OJBlWaUe5xkG2bd5Hd3Twucz
Y4mf9DkNUTpbQRKY+8APagI19H0GjGH8PYu4WJlJz+VIVvghZKqfCvdwilsuFNWYIdcbtZ43XOxu
HJ6s/cpNWQ6l9w0P4Wzr0nC9qarBa0GMAUPLanRqLMNNQneJcLzEhRaG8+6cmEvw7aIaOu3jCdd+
KEvMz0K2OeF9OFXnd+qJaGkQvIWsNlLZ1wfjDrpQomegwodlIFHxDtlDPI8JhPzS1Wb4k8nyEPY5
xzrnC/e/kmsYvd7WXAk5MnsPpObisqOLcf04D3HXdEtcpiKt/JHaMYuYMM3TOsmyJ9T1e+nE9lBB
qYWfg5kAM8vfIWuYl4Tou/wvYMD3z6vVkLOfm8seqObihrqDGbKXS251d4iUu2R+hT1tTI2xqkfL
pFQmDQKDa/SQYprR3RkN/+zGJQkffAFNqKjH3FInQKLiIfWiF1VbvQkKOQpxl449eeomMQQ6wUbl
L7oyjaMgx6gANmxeGDA+s4vHjzH2T+wE/R1xr2Fh90SvVQVVF9I9z3NuYIRLnDCiZSjFMbWU3z0Q
+P+fmH8mnALeFREt9rEfvCNmXcXthB4o5dLlZo2UIu0ZB3mERi4VjK7ANNqXwUE6tNllG7JHFDNe
arJw8vzBN+knWRIXFNwqLfWjWjwn/sRsWfuLa7PdQeEXLf70dugkBZUUlrjWqSrOW0uqYSWpB8Zn
TzVS4cxvXdEwL4IuPqfrtGHpm89RdJItTf6DRGTQVoJ7C8u7ER/NvS6g160cAvnOO2/qXrwK9s4Q
y9P+eePTxRyfNUqC+oS4zDgB1R91F7M8ld71vWA8+99/J7P30sXV/gYrxZaPlYW7zSKrrMPXptkB
+XN1Nt8tIVBX5yvFaMwOKTiXeQ4fuYxwEOzNQGeGCrwu3QcXDma2iNtGdJfc3rcACHLIEQ9WrVLw
TqtbzH7fRflI2Abvh7FsHearGBqqcH/4motEqkMf5aIOtNpJ8EFCKKtTWUCC6YLuW47RfoHZSWS8
pR522UjcjRreBNjoxgEYXiRvNhVwiKJBqn4M/hvYY3Scsvgs3CtzBkcE4SWVnzDbKaN1cFPMuGs5
mz7EDILKiEqJWma4WYU06Kj8Fvdq0GT58j3qfgv40pTgziQvlHm2cjopUT/m/tsfKtdMm9dyh2Si
Za+B7/V2zXoWt2BhoXQx1Yo4yYGm8d8e/oflr2LGNDGE8xD83acFD1N1nsN3HhQIPpCKkQ4t5ZZU
PvyYQcr62kB9PwKCHARBlt6jDoQnsxKnlULjnmSetms2PCNvFFeo3qAWXN1zM4G+/UtuPedqOxGI
Ce48DNwEpJ1qC0NjC8T+DNfwHWFiK1tNpQ/xiSHqhQ1PatWSFBLwq/P8Y3iMaALHVbVpLs0AQcXO
k1wPfzZGf3G5KR8NFWx5NwpznJ+N5A69xRzu5WTd2U7wfzxCndSh39a74mBv23LdFzLCbChXQGEm
fFajgmmr7xF1KYXDUknE0HYkhAsez4WMN3k8ebLkBrp0fP2PsT7tSN3YAA9gjilcW+jtcEy1XnNp
Sf6CujwU7P4/JJ3Q0rBo7dvZR/eUMH0nIZFyTzLcOsFAdhL+Lbt8gOq7VnnolryA9D7SL1XMN522
d8DXhHm60dqLsmURfpUmED0rZZJgPSyXitMBQ+0TFBWSYW6dQ/uJjfVMGs1TZFqbqp6WW1+Tuzjn
6hsZAsjfKbDgnHF6NTA2n4d/ucHDQpEy/IybiiB9jm1clKYM/JenCMopnZola5Fs1YTTZ8L+3S+u
4Ro2Vn2WCHQRh9Pq1sd0fv6ad8hoVDpCf0jlzlpCn7cJkbaKsVZemj6ftrpOO0E/h35TYbvhJJ8j
9AYHAK2WjOaduDQVXLeU8jYGQbuL9tuQROIq6ynuO1CLcuV1L7fOPxK3J0QKv/FksxSYIKI3FiX2
C0Fqqqcl88hFaFuI9ji4QbKIoVYCsD4oEV9abJj6IVur+ghAxy3mV+2N+a/BTIgGApkdJM+2g0ic
KJVXT832cdnQN9QaMYqwcluvIMSHbhBuRlQsDDq7jWCIjs8hBgzRIfXLa1cn/mue4OtuNoek2I8M
RoTeP9kBFKpf/pXHGD5Wdz1jKM/0fyKq3u5Fk2/Nrtz8RVpKpXaQ+qGWhZACy5gvfZDS+o68iC2u
18aMQIGp6ynGPUF04B6GnyeTGo9PWhDnkN1J8OhgC0dikFMnx30gspVgJsJPSgmOVYufDY25q375
tKoP5OtrVqPGfLu6dfLWVl2/A8WDf2LkMI3thiyfss8Xv4PbQVjpO6sHbOfCZe5qGjc60xWZXMdW
5K4V2uxWecE+ThYvlTRsPGMA9+KMwkGtXWso2Hpo7jGJGZ11Wm6tZEwLHwRcNCGUZ6UE3z0phDqX
/EtQHA1nzWEOVcj8agLJg0a2dstdduezTQYrB+vdv2upacrL3HMrKMsCafFgDPB20t67O3DUOstH
DG76/TaoRSZc6sBjksh6Cf5UTLIVhZIpit6LYPX7PMdv2HcKQdgsWJyseV4PK3MN6z96AibXmxBs
feodHf7tI5g+ndhrBlL8OuVpfuCU0qKqjJITc31x58HNd1TWtFShv06vhvIk/UG4zptA/okz8xIz
pNikl0MskirQoTCPnE6OS8vRZM0uTFiO9SkOq4CebAwx/1qNd3Fjl227CTjvuXxGzZIWA2IXOd+P
YIEpW23mN2v+8T84CSrsdyGpiqm+/inGxj7qYsZ05qqqZ/+qiah5aA4nL8Y+Od8i7qWKbY2buEJd
GW+uTz6lCSYPFN6BLqunN62nCqzo8HhzEc2ZB1MTaPY8lMF+RaJcr3cuw4Sl8/bqNKwE0b1WWybT
/sfQbyr6OvGXo1+c7WjNcWQvBcyQE6j78MEsm3ZFuWwMGUQc5tiOlRcs1VC0uc7gYshA/bU/bSwX
tSMQSxijS626vGg15vQS8RdFp8pcknHnzxanc8e1MXNTvtqu3UB+hD/jGheJRIO/oJQDQVZ44Vk0
anxDa7hzqhjLrmKL3+6bQ8wW7lJhmfta2wANmB3DhXbuBMYRbSJyH1G6JzsTinIfcwcS/Q7jlXbc
YQgZBfDa5g0+mcDs39JcZMk2kqbyl5jRL/71/vCBo+rBV1VdpTxuJ+kpy1z6uDKK4brCwaxmUdhc
7qvIXNBrtQt3pZYeePKDRwmwqvLbkkGCANXRbNjuBNG0YEEv0+W5ECzR8fuzPbO2UJifKVVZfifC
cn94qlceMR85whKBdnYiouJIvTdCMe5GK6sE8nxqIYVYXkrtdHAqpvw2iaowxKGdSn8v3zVoPRW8
mduEaeskdFwZTjBsorUTC/HQu6E0APOg20GvuOSjUXQ1qb2rnJEcdpefFWnwfYdtxWsarlHfKayd
BH8hl4R++GfRdZjVhJXStQv5ddE18Au9RG7emzZmpgO7stJUGvysuJ74viH+Wc46dzJiXSsFUfDL
wcS8dgirvOX0OpA4afQdmd6wn/a0bJm+J3cBAAAg9Qp1xiHchdGqKC81fFo0laC2UOR0cZfVxQ1c
8XWXTSizC7XOb/Xi2PitzQv2sUz/loE+FhSio05WSssKe4y83tCLLUE3k/Kv46I+rFuA6POaJSjs
ikL/X05FPLwFwB3xkQXbr4Hy4tkorRNPdqJQKG+VjQixDt2SmXfWXlHzMM5xl0k9I1tD1/l+C/Hy
oG4VD6I/13QvO45yb9Dsgw6Qmn6SdN6LO8jZT/0Aw1nz9ylVajOmorpOXTpvp2exFKzFiXx2wmmA
bxAlBbVNlOqNHo353rhYReVhFNDoFfvCuEicacSZRHETQT9+wCLWCUKJdyAylpHp0Zz9VgMPKjKr
GvTV6ERgByKK7iaX6LE62R2wCcDUGkBVZ8XsSjA6bHtAfesoNvJI6Cgq2WTjKwNwD/29Z6dTplq4
6oHR2PZCluyWkXIXMKTWSAEkhFhX5LCTxfJbaIbG0gupkl8SRrwoqiBPYDVSO7vVYRiF1W0sMeSe
bSbeNT6iqW3n1mdcs0pGWZzGSgirGtdFCSgYnjeiHNgyRJXiuGTUXm27ciupUU/KrJeJt8Mwe18G
uJd/RRXgfmnjG7cvetlkZP11k21WcaNcf6eT6hy7+dR9Zs1GB+JEmBTYaE45CD4OoaP/mmcob8fR
GOLHTfsbXOTcGyQrCZ239csHEYr/3TahAdG2wXDrSH8MDWHmO8fCyZ8kd/niWKmSfRIDUwC+VaWh
T5ifNZyM/HGDnV6mgbiwHY/7wieFje077BYZx12DQKySAY77ZHnBH3KG2z2AnjafGr548dakzGI9
52S57g/aDnCrItw+2EYDuyTGX6ZXcSWnL55f+hAVWMfuBtxUNyUj3wTSNVBdlgX+gpMG4BDdYelQ
MvIFpDT66ZF0qjXjegqpeeaQSheCkz86l3VOSywajnZFfKzw0lJUaDYC7M6EOy2VwUCgqpMUBgJX
mqjp8Z0I8XRs5dssIpQCbieRHaoxvjYkPMyV0nPkoxyu1GrGt2Ydsrb+dNJKKPV7c6NByWwSfIUq
5IQP+r31k8RKk7Ynb7gYfylKF8veq08SEpARjOZmL1qaNbiIu9XKIBaoEYhARBm0Ud0/cB7Jv7UX
MnMj8eqKafV6pxjw6Zaiy6qzZov0uiae6gf/PZOjdv1jV1o+gQ8vcLVuLy8yg0Got2wHeG/GVHOy
yIkJxA5awM6UGtLWZRu2IW7ZWsU6GxfUvZI8mUWnVY2r4Gz208Af9KP2cXybBNXMbfrC5H0zPl+N
NJlA4SVsuVUuDSuI+EmW76FI/z2ZCbANBZQekMk+mN60fFRSV/Bjx/XKJ4J98G+57HtvaOtpplXN
Rv1hOeDWgHVWy1ASDfaW3wYAgI3/3W7r4UeWSJZ0XEIYrincpeknofPS5X7UThIXMFaVGAkta+x4
KNY1PWI4bDh8NJgmRSUafrKmNOPjOW5CDGnEXGwiHg1Uw9derpnvCOzcBawzDnEUwZZbh5BHxRoJ
dl3vk4cfB48GkNYPggpjGBebKvl9Dzmwhykka0S20rTkvQ8su+fyvxc/vIUGkWuZtuBJtCDrmAy2
+rTyM8oi8jZFIfqLz0dFk4ZCOLcEKIEe6uwoGLU5vW0BMzH6RQUy/ljoTqNwBh1ZGBEi55h0L8eP
yBvAPm3R8JgBc/n9Agne+80pzHKpwVzEexsvEVnbSs8UhKXJITOLdxZk4v40+I3Ci9NPxLwXOiKn
Vvq0O20KOjtrmRFdPHoNZZ4SFaUUvaNf0KGsO4ccBxgQGI5M40btjPQToMkBukHunx2c38aAZcrr
Z2pPcu9EuFPDsuvRbeEyVxjcO5apuUjXjy1XBstNx/R3LfGxPjqNb8LKFrc+ufGa9cWi8Ocr6DOL
pD0SXif85bxzscXsOWJl4hLmy0SrORGHsvCjCmNjGHzimmKKXZNryv4BYyYHiPsKksFRegzZnBX5
0Jpve9hS/OFEZTVwTSEzSsU2hdtDQHcVU5cuVRJ0Bq9IhH8PlOR5S66Rgt/WrtSCcyNkms+D3XMS
dWM3//IrT76II5js4DphJ1OOwfJ+CxF85aooTl1Z/rCstnh0u/n7mV+UtEuAvP8tpS/wiDkf2e2e
7ao4K2FR5cK65hi2RZa9R3vJlQ5kFE93GvA8A5sP751WvzJCfw380A4qIMgCt3GnSI7bZO2gJP0L
SRq/cfd/HysMaRzo59k4A+CKi376WNnoEErLqgbJ7aZDgoSWFR7OMj8aZn2U4R5v9RBWrQ6zSDxL
F1KIRNGXcDhMGJxrJRLJIZ7uNe2ETdOGMRV6K9XwHQ0rrJA2XWmki4MD2TBFKw3P6nkCXOJLyHvO
xytzT/6cFoZ6WnQhYgkUHdMsoGkPzrTyYb0Y5ubs3dwqJdsPeH4KJmRb1rv/jOHGXjZ5mcQnTaCu
yuyLqcAQMS1hf3FAzOuS+LtcSmD/nUm15GzN/BZ239fxOqx/egS6OoSv6qLdybNz2pA9V6mwFpMg
5n/oF08IDI/yc7ch5NpxJh4Avie11O0/gQdzYFD11AJRtC2oAJZCAIBQupZgB+zwilCtWAxxF79I
Us1hBJN5mrOTRy94jyL6+Knsy3FX8mk8/twdvuFjVO3HwNVZrUH4ZHLPzr54IoFSGcmQd2QFrbjL
UMV/5bXdpxtNgToOg8VQ5voz9JDWf5cWX0CR+XpRiG08GMKoFVW0dHF1mxwHjnk6HUATjZEo8u6W
P4k2+sXR3g8lvSC0wk+D+nx+KliSO5YKtALAvYIbyyy7jCPSOJBNER0c8q3DQtwj+hblSa912GGF
iORVWdEnU/8f8DBcWHaX72kfbEryloAHXYvnFFvihHI/tCarVAQ6dJlAYcyfOy3IU7fYx5vrSnHx
GuHcxbDStYiR89dO+HtUNWnKFkVvnwyzP6ZRaVCHOq+JxQmjB6zu1/tDb8q+fRwYlEluQkhXiSMj
7bFit4I4Gmn5nRbsI1pLjqylFcdoT9P4YkyWldgiVa1IZAKl6nXjJy60wLZD3OZcvvl2J0t2iy2L
rlPTaySD2e6lRcYvJLWGPny5PMkvVVDuFxA4mXlPyRpSfAFoFjwHjm7lcwNknweqAobx6tsBg3Da
wxR05qKbhBDnJX1vfV6DjRpmA1MeFdUx0X9MZAh2qP6oT6rianUUEsEVGbQqOMZwusqPe4iouZ8o
BwjZW8gY1D8gl1VXReK7ligYGIhk1cEMRs5ktC5XsuDii2Slc2R4iibfC5Y8izCnsFI4k4Dxskm2
PWJvZ4VrDBH+nOrNJM/HUd07s18dFcSfEquXhP3/2mMl9HHXq412UIurjs5k16qNzI+IgRDaKw1w
Y/fcMZVAA6BxMfPNldpWA5pWe6eW7CbdR0485VbYoqvUsQeQq1yKAVE7RHyaW0IXUrQcZ3/2fLYl
lIwD3M/moNof/m0C+87r3uzY8I2Bps56MaE4ZgJbzCvSSA6F71MEo3huksAqZCBIIaI5KQut9Zqm
VaxHxXPwIj8xDBlZ2nLH0Aw4plcbr/ofFqZDcjuh6x6QwhKVXcBd6RI4+Dl3gl7YRllY6nZgKTe5
CnhqUTimcBkGX3Xhk9LP0ONBEfFva+ZTAoeEUQcq+VqQLMMSpmTZdGvEfv5+ugdJoLxjWRuIIRFr
RncVF3ax5rc2TsM+cwTcCikNN3Sr2GJgatm7IKQOOMJpnmI3atPt7vv5sVZABB5SrKc00MG9Mj1F
UlxeH2umLmR0uemZPvC0ew9+LozARrLCzQJPJ3Tkn3iCN3oka2hfUIs3JVbmUVuI3wwY+0YVlGwb
HDpVNO82DGc7oxLm01o+DF7jU5DF/tJN6e7sIubkQoy1GlRp090Ko781QjJRtUD0Zx8V2Uz4nPTf
adHLSPTAvv5Gan4s3cPGbKf6MMRFBl1Q4fKtawGpBx49qOiaV3vMnDfhB1fZy+6MECuPqLqAFWYt
SMedmPkjEZN8Mv7gk4eSScE/ASjlLixVvI92SwovPxMao2oFd1xF+vhNxcb059IvModFESKaGOfB
dykNWb2Z9Nh6lCygsEciFwp2VL+VKPJOCpHcVJE2dFjmNNVD+PqXvLJgtsyfI9HSJexl4rqpJURI
pikzngj8KpCowrvIaBfsZGqiw0b2ruqwK8EQ78Ew/PiSRgaf8qtesrjt1IQDx/Tjv6N4PoWT4ptJ
LdTO2NwMvE83wWRvDZX2ADg0FmfeQATNT8ZgL0uP2+ifs+b6qXG5z9dBOAyx1nTFPYYrR948LGBs
f942tsWa+3V5lZi9AILdZpuPSvjvrUrD0QlnEBZiu2QLK2CqK5mLiAXhjgF7GhBEZHKnKHrDHJ01
cCBdniXPiLtXRck80zryJ3xsJNZ+Dqvqp8ljlAXH4gSdEEFCQZiLXwaHjk0gYbmnOTlgWPacL51t
43DPJN459u77bS3s6eM01HoC8C7bu3PNPR4r0D16il4rXaDcWFJqP9Xb0uqxsGCDZ26q6TfkVT4A
GX2W2WFW9UdWu07XmxOoUnAYeo29Y7BzkyBiylUrpr9NY6ydDJiy7XaQ9li9pIKFk3BcGka2qn12
i64pe24PhorfnQH4dpbqCsdAdU2vGdSaDvT1ljtmOTb4eIotMLdibS/7fNWmdXIVPdDjXcGFy5Vf
y2wSXfhT4W/MxGh9PLXYOQPiCCnqjCdG+U5xJHwVQP4QjLQDAOpStpjHdYie8NY695FrZXWEQwdi
HzGY9BjiKrJYE1n4YfqWe/l351/qIFbg7chnmvdAbQ9CSxENVTtqZDbbdkns+lsaIWzIk4mpuFx1
r6Ckev8ug18GiuLcZUHm69tTuczwpJTQFbQ7Sv0/OwAwFnhlDAtQeO/bi+5w8f6xOsVCy9s2RwR1
5hJoLeOx2rJEUJipDDt58driDY0n/fysYcKNYw7WFSSp3qR5lyQGc9z0ZntR4gr/ZPUO75cA4IgO
YPbIAtz6uNJ6cW7/OpWWVH0tyib3s1dA0oAwOvEry8UruOyHXIn+lc0Yew4/4znfvwKzOELtDHrK
G2F/KdtxBg8Q4QOutQ+/JCwk/UcAicy9iZ8INU0M2MRdQFHgjDo9rw3o+n/vrTPZ55mCFocnpIRB
9Qo4ftBsD/inquoZ69TYb87B+h+2hb1pCviiATPhlN6kz9L03nwArU/FhjCbz1hD8KtHrGDGQndi
CVT+9L6SGa7ujd6cYXhGQINs66ZSzE/YrXt/tncgfgBPjyASD7zcQR/HjSvRw6+gBtJzxFYtoIp4
UrE+935MGbSclapcWKdG0N89PXYtWJPlSz+/wjU/3s9AE6yQj3xbcU22nqnIio8vH6t0bXnvwWUj
umRCiY/emWgBvd6tmiDUmLgbo+A2fzT1j6wM84V39JS8kzI3lInfHjPjxXprybAW22ZtOt8pfjYL
YFcsEY2GfuPgvnZZAjOp37wHQRmOVlPl3jJEjKCQeB4dmyz9FPUpifF1bAXxxGVkFEVedNpSzDQj
JxyMc/+z+GphoUP76+xus5a+hx4WFSgS34pmJoXvgk01ItfI5OPvfpaj84FtMQJrKhaDUk/Nw5Lr
lsJr+ElAn6VdYc85GGe56f1SJOgUjsCouHbQO5TZldU5e0j1ujIsvdG1Tfy3bqvXHV1AE6d1X5T7
MtNJnKHeLuQSGn7fmDquOZl6b+hV8PndQHJW7c12y1hFFF6eJzzWdNu50hX/TJAB430WxtGyvrqF
8vVWaZzMxzPz0ZTogL7tQvExNbqu1e6s6QDSiKNlyqW5nsXItwt/lPRqeJM52bfa6B4vuhX2KDdJ
IfSUHGG70YTDBaVx5fd2H9IjNZceggvrk1tGaJQLQqKZV/7i8kz2a38/RUpxqFqd4m8lT7TFJzKc
a21iHl5xVTLq1A+DKb1xUjMFWmHKio3YTE6tAAjDtDkKhseIHPTKG+riWkQAJdpf5p0uZ13+lvti
k6+zIahAqjoxZ2VUx7lVdwZXAJarDD9DktlR/VBfbpDWbrLZU/ixu6fVVcCF2nl9dQojSLWK/xIl
NPAOie6z0Lp/BOvWMM1+2qBFzv6COTIZ5HLIFr+FGzr/cB7Onw/a3YLzZG61hiNBWZoIKCuOh4xa
4UVu/LJGe1Bi5CVQlILxdaCmwOei2nB184xju0h9CE6Zr8ogVpQKvcdXVcUngjWkwPbF36ubs9T1
+Sw/rK7a8lTskCpA2K09EzTQ6H3tcPYswAFB7s07lgsfexSENawP25ZcAwK34DQwgdyJ8Bi65jaD
QM1l6s4eH4EDpi4qNocd9qO6lwK1hvFQ8tUjPNgztslX74GG9cs7yWcZyGRsUi7G34fxj4e8v1zi
5i8yklVRs4Sz0PTkwdleB+/0zWXsCW7iYVUFz7QZgOg+m+TQSB5W810Njm6YMkra1h//2wcZB726
2cyxqKi/AvYA5I+UpLNmT7q78H064HG06vaOI099XykPBdmgQU0WBo775NeYx6oLdJmJ8fbWxoZp
JO//pyRqmaCE2UzkaYceNNJMlTY8CzUZBDJzNzmu+9ngBROBRJgeuE6kSukCBSsElw4taV/32UIQ
1B/H1Tc5d0o9oTVkO0HUQBRpChqLajaCj6z6722RK6xqb7IuL6nazp2jnKksn1NAmtzAl5M2KUMX
2z/BI5lN7h93/Nxzl5EH2p5SE5GbdF+fhnfJ5fxU9+vl//DdEGhzrq1P2j0MuFipO4V+einpQyZ6
YESMvNqzQZqhFqbR1SQXOmtuVWpjIpCFSj6lD1pE/FgCO/Q+ZA716qTbZQi0Yj6ltEicIsShqA1I
7KxuK99GpIl/x/2tf06vRxgUIt/pvQBx7IetFN4iEEzQCWLTzrmOP/+qqj+JEUzDVpZiE67K9fvV
EE6QohPdELcB4H+ttdnR3ruixXvzsuHZlxPi6NV1eA8X1B98LZFiSTSkUhe/P2wJDIRzKOMV+rMQ
XnXKkA1r4bdQDggUuMfeYkDvgyD0x8QsoJ+01qfFF3aJKa6kblleJo897UP/7Z4KIBn3TvcQZe3u
d/2IMPrjab2ysrH7mZYUrC9C/AhotENMiMkLTJmm7fZJ9eVuRLwR4zHxnZvRwg92bKgy8GNdKmZy
jE34vTXLDRewD6eks5Fd6umEHp6mKyBijn2AJQxUlC4ERdFBAFnfGmZS8yhIliJ8zU+7nNTsyeAf
oS45T1pK3PHuRQa+B0O7Jb3AktRL66RHiv5bllMr6JsoyTQeChtTtd0Lk9hcfzZfKC7VnShk9cZx
OdqyxOLhDECmjeNIb/wPisZ2AZOHjznDbsp6Xd+QGCIDAGXXk602f8oNbgsbOPTUmW/tZwS8Ur8C
y6oVLZClMqeMznbns2/CzfvJga1zozdEQAy20hQzEmxt3exK8nnOGvMkm5r5LyGxU17I1eGRuZaQ
PlroIWy63eheL+M2biXShiCaf50TdS+DepnFrZG5ZipNOq4dVwwrW/9ztKVqjHvrL0nNInOTuUEM
qwb2s6Qj82BTWq/htL2eUsYON+uo6HnehL6cVYWuwK2pQG/HlUHcuT8YsN4pjOszvMFyG6btQkbb
nP4uPwzdFSqUjrN8GsMDR4Yay5NF1IEdgROUHc9FtWVvlk5o3z8tO2cBS7KBa6uGdz74/O+rgSOO
kaqtJgu0UCfZF0ssy1EsARFXeh8xAO8DkifXa5U0oDuloagV0Zo2v3uAriauhhR+FDC8vwg/OKCr
S5DjhzncWwC3cBYDFUcMyiQJ7Wskq1+X8eB/DnyIUAcymjmj2dmQhlUbcknsw5ayaXOEogvjTX0q
SMOBXGZsdhc8BN8T9Jlo+sJkdaXNBeEqMzk3Wp22FtkmiBYrPBSTPOdoevsuwfkV1gEIiHpcT3/2
HNF8Co9echf7wkvoQZiRivZv9x01DjejKEePy24UxMdYiZVeM3UxP/jWcOJ1p3zKv2fsr0EhC/qN
H36YIy50Jn1wdlGkvSw6JHRzxZWtCV6r6vAu2t2/nHN1mZD+jsK0ThKzmtKA2A52wsd/hn3/u/O2
9u5PW/tiV9fcasOiVadpLMKTI6nA4nXZUZTHkLnfPseSSQKnnwInvlEKf86pVSA8ViUTKuyz+5dc
s/fCTejmSK4wySMN/hOYAQFQIxs7J6lnSslIzkHzRnToBNAuSjfwLY4l0iL7dj9g2/ILbC0c/lpK
WLBM9vdyAXPokTm9jcpHkqSrpt/0NBwX4X5kD4qlMDeYjB7b8zwtVtE/A5MgkuZqfEkvv2FgwtdF
YYQWNHVQHDHjQCiGEPTyHPM/Ec/CQqID70eOF41UAkXYkW9Z/yRWiORXl5q1iC5tqGDsG5KZyr/h
+ka+lMU4p+anryHN2HbEwjVsJWSK8udjOjCTkSx8R7nmM9Gm53LfFvdEwz2/i86rZ3pVDkQiN1u1
tvNi2ah/AW7xkB7a0dwXZbINBm4NO2OzKCA6JRh0OnGA+yD58sGGQH0FKWuL7RGkXPsaqmABHzj6
U97SMNOnEMKzGsmtzsZ/Xe5bDUad3L+u5AlTuvNl3/uvvlDbOMeFR+tsXFs6ai/yXwoRMB8m+nai
ah9znQI0nCUT6vR7iwlcljsIi/aIDLnMdyG20LDu42fsUlC1GzIHcs1moQs1JRYh/GbMKIABg6d3
PH9pODYDjXLZO2R9kKv7dPkwMU5KKQWQI4xdtVWhUDrXqc57dZ+kc124SvdFlVUdlzY+sNTqjwAt
GqTU23AeigTy5eCwup9kFknw2U34NX5nY8BsW44FwI97+0F9KUYJhAVz30xP2GfM0F84XOGyAFNJ
MF18CTLc/Wr8Xu/kZ5smTADlY+RKHgBN55dzFKiojqSxf9843D2+Xq8yUUC18DxiwyQfrFVnI3uC
T/vUALgduiyE2hRKF4lMHu4lS5E0Vur4bmvu8yxvywC/fHz7gAyWa5UGw8uQCRCoH37InoCWAHds
2R2N/vPZdb5w4VOBnTnKu7jHMJJqQJCTmLLRQgiBy1wchsNfmFTySXTOL0a7fNatZaHJ6xBgxpIY
iqVaYxm8/CWZwfp6shqfu3rHyp904rt5Y33cCZ7fVlGwgHcZ+C9u0ygw4GNSi7DtE1lpQiQRsFli
NyEr5lNjQQ8TG7s5UuOVZ8jizQzlRW2MiLoQKDMozbRx8HBNIjvWm/pcBsIz/wfge8cD3ZJOmse7
ILffNg5G4MoAhIKtd3FFtdJ7LJDtOWfV0p3qQ4ILTPFL8rp/Biyd9LXa3oBmYZYB6J1/5GZzZchx
tMN6N4x5p54pwCH1RB4X3MfX9pfthci49La2zAYXepTgnUS6HaBfym2lxgFOL2X3KL2KHlRXE9KF
BGJJ4PQk1DU009q3esRU0WtMTFwJIS1Nmkl1CJPYHTWw9v8RaprwVUoq+zN8fe+10Uw5aOw6gh7w
yspd3rf0s+DYxO9k83zzT6eNtyvFTf1ZKN7frIQ9xlIzwOOjhYl1uPTFqi56TmaQWBmZ4hUPBnMO
0ha4UBhSN2J9JYenWs6G2ZGEjzp1cb54leiTM0kaGNlMVa0LZDRpQtVV0b5fMfb+zbEOaoWHtPxw
O9oSIqUVUyFOhxdbLMHOh07pmCVvUfVWS7DafzyoV5dD/Ixn52EupvKFwL2/L9s4JfQ3u7IfuI0Q
Z3gORvsT9Ovc5XY/xOlfbBRRQkMKEzFgcg9KaIbvWodudmxAHhfSU40DVtHe6V9V3md0xcsURQJ2
uznFsl7iJPkGnfhAc4KiWC86dbWv6ygEr0ZqAoHodczAwXIf7E/NDmtJ8Q64ricNk7nFPE5uX/UA
G4ee5EobxxkD195MpMCh0GyvmOx22sXthBKsz2i2hiFyvKlv1KZBZLiRFKeWamarGGxE4KTVbsAP
D/O80OnFwJuoEY0LUZbKAI/IAgO5W2ma2plGL+Ezf2JVR5qkkdBX9O62+5AJ/m2YIKSA3VUVCF2I
yVMQK86Xafft/YMhXICvwr+C9yk3dHVrgSohYGEcZELUzgx79Wn/dQcrNKgZYdPxKEjMGc+FkCY3
2PgrSt0PLH6o6IpDsiFr+7O9gPRR4PXdwjZ1LPSksp4LFJb/ZqOeQFa3dq2nqTLGT8U2gbysgYxV
k36wmFNqbQxMHknQTmVxvT65L14RQB0eTsiruCOMczGT+kumG7mS/z5y7EdFLyK/o9+LoXf5qQn1
DP1+D3pKD9JmH1xdcek3iNXGDcutpMITAQAHWISPenC499o6lTE2anYG2bA/p9h5xGF7k+Hqo3bK
3vhameFPojDLwI8LDs4umPY6VLLlBeQXvBDFPt29bGowT5ixNoiVmGEV/ZtPFascrjvX60GHJcPy
WGqE+Z5pL/0Py4dADo9LZprznczZSbUz+DXchOk5nBpADLJ3AafLQ5fH9rGZDQShIND+z7JkUzHL
BfH9dY5V6r6JU3CB69xmllOxp/5U5wE1eMdjzb2zasmfrSnhJIKKXKzau63disopzE3/ifF6lPN8
m//p5A5JfZFMmIDI3p21JP3siDLwPCuQL8eE+PglPFZ3vlXeOXSa6hFRk8iv4mbNCN5cszpkkiHs
V9EhqNFbgD2aQbhIzhbzdaUfQNDi0y40Nt66G/dQPbuYw8PdMtqiqIzJ0/QUbZae6ic+Px9v2avL
WYhSw0g6yC3HSEh93NoDRfkp0R+O2eSImZYRcB38oEc0hC80zxAvT3Zx0jl/4sOKKYjWd7UBB2ay
LCEsOvOVCk/sVDtL97th50YE2T7yhgAqFexPRXoge6luGJqKb18wmBRVWtVgNTpm14vgqjPw+XY8
6JQdd1POcNtsIdiexplSGfbYJu+8Kiri2aQAwvHQpkvyXvM0pl3oZLv0vf7vW6EtoccI9h6zElrk
lcnf5yCnL2SswCkJARSF3yghqYgoDAnRVnl0bAREK6QdGq0Ok3cbht7xCcz3wQe1TOaPA/RhMZ6r
aTpkt6PQ2vj8SoOW+Mm6G9ety025ptQmG5cLwGj727ngp2hcvX+nbD690QM9lijDlesdYFAY1L/z
SBD1XJMq8KQrPdwUljt6QDEFvel1lFBHqptstqmMf0tzFa6tgzjZiIcM9qwm9CIxH+aXlG6Rbd6y
xO9KSh/2n3CynbfbtM5pmterROe4vvOwLSQT3tdTkyLCpL4osHY9JIe3uWey26c14sb8Kg2up+ff
66XG+YlmnexfwWEnmsLwwylNCN3v2ety700jnWz6dQGlh6JcKuLUBPo4iFxUOXlzJ4NePmcvTJ+m
tT/3/VfNoOeMzU6L0e7+qzUcJxsYGCe0iU2FFjpN+yBNST+YcvxSGdVupYrw+SIemM0VmVZxc6z1
bk1Ja1PCpCFh1sM1DSVeK05WIV0hvvb3cy2FbIKr+GrmTGPNevKQn5AT9SV8pvO7a4yUAaQZRIbT
gjwFvbGrgxCszNQTn1vl3wR33p7aantFQRi6564h7fmOpNsn6A4etfI1MkQA+5JOpoXL3VI0wS0Y
Sn8i0q60AKsRpsBSwnvR5kLvbpWJ2mrtmKi7YBtn9KCzxrEYchYqBw53dGRpdYNusF8UB1AgBz/0
kDT7ETdKq5/fzxIHcew0SOSeFAoBBB2YXi9+0m6aKe5nY3Hq0XPdXPitqXHoPs5Vk05YU5M5C2qn
v0vOpFlZoKpgBxdJNe31myno5UgLATLX1aTy0vIt6xYMmnXSTmXUavki1EJ8/DWCRGdbmIsjq3+L
GzfcgvX+yn+SzrW34/jcWX7pU+FjgzDopMg0C43Luh/ClBd6aA9qNCbNg09PBsAemzdtYrQ2XI1q
AoyxJFn7ZYiH3iCEobZ2eYBduO0zS/bc32TA+/wMlY+ic+mntCBi3ig79OcgRqILkc6B2A/yJb2m
0H6myS/SU5vZdU3ptlsSFgNCeUupONUsNCcffClcEBTceRM5DSCdutdh4UuBRWkgH1UgjG6i99hB
1mxBrFbJkgijMn2TTudNcIe1YnwJZbW/FD1KEDyKnMX5HnJ2lQgb1TqUz8GiNlb9L/8FOHYlMEw9
nOBCIJEO2NUgnN/klXQQnz7icHJYJb6EWSU1a9Dm9LvhjQeDl1Q+h+hQfmczrHy4N8OdiRt0+xow
INAyqAH4ADzt2Tw1qUpLXGjxDoJg7aHS9+KJQnpmr0amtZgNO2sTIEnDTiaaYmQAQfsuPWORmSFw
mRqCUjwIKxTigbnLuwIxAOpEjwVGchHcjQGWnVqDstHoI3GJQft8+SXwveJ1ydu136W5uuAbxUX7
1/QYlDFdHwu0npsVkqvfWLfikPo8jnDo6R5n5m+I0gcqiD8FMRyTs93VelizbdSGkOo/O21cbZQU
o5V3M4h6XL3eYns/RadikQOgXt1RzAWmcVhq1J0+ULANj3XTJgJrpQaWn3o5R639Od0BoY1kO/dr
XCgbak6ITddahMXBYPe54AjtvJQ4lZj0HNdgNBSc7HyOqN61yKRT7qJhRcoHg8z2mVz20CbVDE6L
ULq6taCOeW8Ih7Iy2U+HLJq/lu7ej4DU3BQqja2A+lng+ibzOublG4K6B3uMpaZ4LKyGrEGsa5Et
dlKoLmqKXfCSbMUqIzVW1Gm89Dlxc+LmEMMCrMYqYHjpR7EZyVj1TQfN/l9HDmrFiKg7HQttnTCM
p2fpJQIQxBst6eb9UcSKpavAQBr0dIwdgCs6o6HxnGi0LvSklaQQLWgqxiQQW5GxwO4jm4vaDBeJ
+8ULwF6QIsnnvsKqkR3G5EfzdJOr5AGJC4YUKYIjaHkIChvhfcIFsJxMwHtAaI0TeekvU01OVfxG
vMZ9RCnf1iGgza5XdA4K1YpqkNPMh/yk/4EJPKymsZI6CY77PJ6VQA2VJlgivYcR6lyFexLsHucZ
i7u/mhiigV2qrumSgAn64RkyDTLUxIRcejUZseu16E93N+49cjCiMAxCPXWHBbja7dk+3v+9e/Tp
Hzu8GfJRAOQzI+t9Rduxf4DtV5TbwICG2oVPvwJ/7vJqvNhR0eS8y/ylO0TF8c17CXSF2q9KfzQY
d5aVBAEaG+YUY5SPyqvofLEVmU63ZkVm0D5p59iCgCpedO8uGB8YZ5IPs7M8/ZoFSWDHG9/d5sHY
sema8xo9gJcQL/5DzRnApZ52oqf9WrXoxoOUT9fm6kpZBXCuskd2oiU1/zSvdWq8vcT9c2VgDK0G
x/F8EffNzRPVzybYBxhQgelfFS2SAiFFoTZ1eVaEgMDrFSrtsHIrvBlDbZK4o+lVVjM8pj9hscI7
jbjfaNMozUm4CVg0Uma1uVPKaeY6rpQcvtU0BJgP8f6aqdYSSND/ZWHXTbhp/Joc5ctJn7kxQpGB
zCddKLHSVOEwxx9D4siKnTwPohJ+npTXS07nTgCg6BYhUTuw1nZJbG4+BbtcpNufxKjQlNOWbVQK
vk4i+NzlZZSWnfwD5J8UNCjc62vCSRJlYtQHTkNofhuuL0cwitn4J5an+v1+T2WK1UtS3VbXdZy4
TiHHluqAv7F80ZdGjcET2siATBRUCT1DedA1yeZ5dwmcMkR7y0NM1Lk/FhUNoF4Ddj+Zi7FGa4F2
IdVDk2A3HgFsHicQm970Bj0t3V4n+orzHNe5zDgSmX8fAZ3yhvfi1WO2u1R3IwMcg2+pYwY1umO8
qiw7REzZCF84coKTd3qIRWvjgA4A+hGfSqbk+uMOa207fwNqYb2bSHfdwOoMnytBjkANb+Udfy7R
ec0jwlbjmd5Y1SPRKoXmdc54uOcmj51/87Pss7gENDNC4ucgZJtspimNK9tNnDt9yU/OfD64AJdA
gV6xhZs5SWWgIVmg7ysaEd79JMuKZ3I/mFGcD39p/xdQQ3ew9szP1GxUNOMwXCADHnCNVmnx5005
6VmGTRUtukkRu6MhJlf8gHl4ldgBL9YPbBdXP9dS+lZ/CF/B9i3VVS27b/1h8KV2joIXQLeKFv8u
o1pJ9VGWz9GCDvpp9kcGo47TxsAmAJR3Pe3dul2PND2vCwkchLrXGIJX5PfTcHzDHN3lD3LZTjny
+rNVV5a1AoHcpmbWT50FGq0PoG4AtTB6hnIRjomk0tH6GHhzK9GCxpMeI3w37VO9pXoVhMXtbkCG
pYKHs/eB76S2qgYUAKm4uRbNiWBHqi9YmdD0fALI/kcfoZisa/5xXzfCyxWBb1NIhs0Y8LNdOPAg
i4msNx6DxKB5f6elM4ms7d4Xwkhm8zWkMmDHra6GdFh989PnHH0qX0krwc/tkkYTNtsgod1NypKO
CCjqEB5jUOvTTMQKoMzyG0Yk6EK8LHnQA/R2cA89B66yhwIb6nZDTW+16d+LOHMfL1C237PfPkQE
UHOEEadpYpfV3R4IcUE80TpuTolG7gDIkXHY+okp1VG+jCJSC8MsmD+d7wMQ6Y6JdspQdFD43dlV
fxX7kHCALEoM9QX3ix/AEWZPkXKe1MjUdDjkF/60o2djy5oU+8zy/mO7K58Pk8yrekZdw6OhFMYe
1WTpPRn63Om+0Oj02To+K8t0x4X9TxY++rtpxN14Vg+ocU4guExBOlOgeYcsYzGtVDwN0aiMf1+N
CAzAl3LmVDrHl8UKmsCpYgmp2CyHNmlGWIxJbo3gFH0I7KD96n8YkzWiRFIKJTImQirHUQqP/6xg
PQfTT+LgNJDrxvDjcks6Zlv1IZ08j3Bk3PAh0gj+oJ96DgeJNN3qMfodYhmo5Nk1OThP2UuZXtxj
G+IVAVFmmZC9Vrygk8BOG/QwdcKR1k28H405Nx5GOD3wHLrFGZoCFtO/5m7Re4RCXCkGQD6HCb4T
cn5zcuzfB6dQbXsMc1p2BO+nqu/8uPKpSHIy0vQKv9y0Ltrzu6xiZkPn8gNyHuMPTPTcESQkbumR
y3I4RBGPCgzPf62a2yV+HapKgQwEVYVi7AD89+z444O+Bxili9vb8g2cVhQd/FJu+513HP2bZuPP
CHyJjtH0MAJYoDCVw5nZDV9rbOP2QdZK++wxASYHqPLG9Spbzf5/U37EXTmuFvykfVdHkSNnph3A
kjJkwKheRa/cOxzdIbrmG1LZyDYmRAK92O+SzjBnuGVmTY4BOVTGwSnpPqqzGSt41fZ4N3Wz181V
saTxHxRFx0pwkX8cL+sglUUoyhS4mP65HRAEDROvAwDrE3s+86qVwes18vTKCqX7SAoNS1GCF05d
lXXIncBRcQnJzvEsaYGez754PkfvK19IyfovOju75PCHSqa4Ty9FsR1RPGpTIKZk1qQKzPdWtGtM
041vMEn4Pl+ZEtnh+AcgfWlbuGQ+Vzk2aIC8712haMSLod5rxuXLeXUEHQYSB3IMH2ReehtEfNdu
MwRVV8QVoaii90Jny6pefBvQPCR4JNehUHWtMlF0OqyuIkB5VUm0qm0yHPTSKc0wLOHyn/GopKGE
VO6krMvQ+PZS1BeLaqmIRa6Ss1cvr7Vn3Dk+XdXVtVmO1m9mklnGRmarCiemUjrqZzUG4c9qSVX3
h0eY1ajGU+TUmJy8CrcQ9/8sWzbQ73IvW+hqB4lVJCXgVi1KF0jwqeQ3iUKbZYQbDXlZ76DrHato
HgxAjgg9O9BC2iATzYA0dZvJfGiYjvQwpn7KwT/AqOM815ryvIV01h82Ljjw2ZZsy5jyDYSxUc0C
dj3qdwq6IPrJgEb87rY+/mcMDQowIKzcnV1PqSBa5T7FF2U6zU4ryN0XEHrnOK/WNQYCdZuxEkvk
5kODUK0WARgyJqfqajlZrVrehNCSoJ9jM1KVypyevEcOFJ+2/Yt659l6XFRkRBNqcEXLSZzYDXj+
a5fYj7KlGC6+bHtPWYhl9SMdZgMDgpc5c7Wo1Awlk3Lth9ANltgn9jdAqfwC9HO7UKDxihgglkVS
QVWBh5jjkqJ68yg4/K7CFaeIUGaC14f/11JKOMJnvSo0pvYgQEUUrr0l2ZYRN0TeH2DI83aQ2cl/
pEPTeV8cmqwPHFN6jdZV/9MTN8BIep27yHrOKdmC/2TQZ/WfrdwQU+cCBOQrGVGQcM8LnYJ7PplP
xSme4eSiR22P5tJ4nau9nIXV9sThJ5F4EaHVBOlb8qaGU4wZWbRKOK32fvkf1ijzHTumgR1TxHpZ
mFA9V3EvY/42MPgIhfseGt6+qeP0ckltdDcQSm+YEgWM82p0p4oYLLd2KeZtJ2KuTg2E19mJU4Op
mhJfsc0uxhwQpLzbVwA8Qciq3c4Mv9A+OrHxC/NZp04pDoPAzDh1DIcvb2Cub0htU9xCXxd9scl1
t8wUtsw8NPKNqSo8jNsLwMomONX4eBaynj9yy7f++ElGUlg+A46FfY7UoK/6QxCSHwhNaClm1t7o
7rwSoyRZqwoS2LQ9dcSq92oSgTzLlo7vr2n4dJtRn8JRmAHLetOKWroz6sJ/xDyD10UbFmYEodhj
+GsOFbFD2uo0hjh3xIfem+E1Qh3rLaAMmUtZs4fe5CGX8qncxPil3hLh/3lkHmNku9QM8O1KBAV1
QRpNLEQ2AJsmTlF2+IhFAJ+d/N/1bTPCAJzBeZz9jzVB3qUe+sZXAgicFjfwUBx49Hq+0F0/Q5OZ
4mAnEpbLizFtEXwnJqv3yqblWIMISMCbo92VnR0G1Z1XA45DYxSTBXGFGvd8oXS9shOQxkkMCvXn
4h7ghqFl+iiaC8RDrJNaB0zmmadn58HB8k8VWVu4wUnN+831A/HzjtOTgrSSEgoCj+mNIflfEU7y
HPNefbL8ZkoJ1WKokwkXiIQzGgcMmo5B7alncclNpi4eZFHOqB80v7ramOBsF39iIgraSm5uhV6v
jGM6IOVVoqAeJFxA1NeXvbPyhtVHMNj1SY6S/m502P3nGYHy34tV9eZ23cJwTOkTrzDAy7nssTRM
xABUS/+DPpiYxzpovHKLQqVqgC8a7WA+6o7DDlEuGGHbO+4wkQKOcVoiURWsm61FD5ajbnOIKNxq
1w1maaoZcnbuh0cJ6d3uz7A9I9KuSrg8wofulrALM6i5R/q8iba6LSBD5/qK6okdjk+PAM4x8FuM
XAW6QCldjg/aFLTE1myX6DYrNTyrZYeAzDy+hUDHjv/C4R5OOo8HnDagmbHdS0GCtbE8Z8bXHrNb
f5OqgOfL4yCnRpy7pjtavCw82vb4AmS9QOEWsl0Op79ILwwOw0ta2HtQTEm/c+Z2U1nKoSk2t9q1
QjluACkIBGdKiQ1wSD5orif1LQknAYX3XHccmM5b0yyTGHJsAai+tcjhA/tJIV7CUI/1DBjWGqke
5ca2GV2OZK4gcHpuGgZ4ysiSnb2cyQ5TVZyektVmhPdGUthxhbfEYYCxcBRuFN1CbTqqb9axXLzp
E7hPO3Q/L/Dk4DMaVvrmy87r7DwgC1s+vFqJ7MqYsrx4bKOWw/QzRsApBfdNvi1NfZfVqEG2XAGd
J/xRIii0QCN46wMzrZfkp15IN3pQBwhqG74Xnn3CE4ABL1EAJrVYkdMCBcWQAz5ShjuiIZ+U4kSH
4jT+sW8fI4hIDbtboShPY1byBuu60wN2WB1y3AXwvi/NPCg62ThbF2q02d9VPe6obep7NzJqlxls
eKgqN365SquhkeN9Xl6I50tzC/ztW0+Bj/uvqBM1/CL3HkSUXO5EndG/tck74JocAdj0E+WMRgqT
rf66nFqZXMh0wuhE304W4hnfwjVT+cePt+P6r52SLib+WnzneN9c4e5WinjFgjGZFb0pg/H+3GKT
bvcFMU0ejXqwaTXKX4dzViGEVWAYiOrESegZJRn0YrNxjPFA4595Y0NW88HB5WD5ZF9lopzGZhTY
/F2EUSUOoPaJX/SD0n560KFv25QDvkqvknZoMBG64+SklDt7p9VYkUJzjo7sHlkl+z3lAx9LuQ/j
J0OzRk9QKdsp4rBSZ5yJ2kkPZrJ1VKla/RAQOwY4kRIIphWfV9E+A6s9SWhM6ZhKI2L2iszFApLT
xkxhu1BFw13SGwdJCH6frkRVqj7LAPjIlypqX/J64gRG41WNIMQdy5qG7faUJpBWN59QFlZHbLb5
T7hEoPKsVI181aUFNYvzsjXLFpGEZeKRUjM/pZBqnVPZ62zBd6qwRum8raSMvltkZonrb1lqunmR
XfK+VDz+eWheii68iCpp+KbtE78CA7i2rheWoCCCgk4P2H1LqYzH6wB5NyfPxnUVFrIBDMSp72DF
M2oYQCYpQmIcIZ7MVVZs490Z/1j/V4bQWGlFWimtZAyNapJpnRFLe/E+Y0MMzpwEoQcfRUsFM/f1
C5mW78JTwiLIhmi8iCI/TZm39i8zR6do0wWvjdR46RATF9nxTXGMZ+K5vsc4+LbriMY2r+tWxcC4
vjr51TtfdrUrLIlX65NA2eewWRydEBWDHYlm+ZKTFu99zpw5rvXpNKmwN3uNmJ+7aNQwFE9tQBXG
bP9qoi0r9Jx2haSpiP5fIjvDPtKPpASxLvcxVodLqBJxTtoqlG4uvtPTIvLbRN7PQge/RFnCJGId
VxLDWsgCYsjiLG+pa/ASngPloKa9S59JocU6P3LPbe/TilQYenV4VvFBSgTWNOVlxRSdoaewm8Es
D0veia+di+aQ4QP9ISAMdgMSi3idTDEpIx1ihKytPayFrH99Z7sD/FE9kucdWQD1Okbjf8//mVSC
OslrZOrSa8fHfP03pLQV/nfHUzLAfwmmkTS/eOmxhOcTJyRCl9NPIOLNINKaNPD5gAyu+AMt7DI9
4oNZpmH6JAyhUKmLE5UQ+TkXwj9KROVU9kS5R7dLA3anmPaFwfvF1no8Vx5NSe5Ght6MpJSxJ8o7
p08p+VJTWiTFFm7xBe2NTT9m1qT0cuhy5CBQ0khWY9ip1xAGkVDkmGl+UTRec99kOs2Q6jjyqx1+
7vjVHuw+libR0mwNU16wp4RsAAiSOAgA16HTfNq3kZaor60zNO7LGooTwM9qPj861BUf3pNMLb04
e5vBz9E2r1qC03SiyVADegwis4e6uB1XnuHYi5oibgU1iZanLcUzZ065S94+tQAp6C0BTtArXeRZ
yUvVAdYx+m92rFOPI5SD4DCytmHg8a+cOJThTq60HO+PiMq7COuuha5StHpUc4KrLRhDs4sn1JiT
0abL0oUjiE3zZUtZ35QmQmxKB2jphK2e3Y11RftMsUqGbRjzTDiyvcr9mu3rG1zUXuLdTVOuQlaB
LqDYytAAwsdmViq8tkIJKeMOh4MidylytpD2BRBsGRESuq+OpETEF33C06xDwvZpB2exOle6J27C
+ZNujwRsfdvSK1webBBJk9NgYTVUIkUpND12YPIOburi3VLjqR3kwsqkYj0+rxi49VDKu40hAXOG
ZLYoYpB6Wkn74xIXHZHJ0wMn6p5JRxZ0M0IIgbzRfzCY5QsZ9jVyT6XRq5ANH9gcj9Bds50KBBfy
cWqdD/rdxbU28X1mz8CI0UEF+2ViGrsPgI8ftohbmI/BidkqpCGQwcxRUYfVIeQyLzhQierzfakj
n+H86a74KjTL3FCM0MOtCoA87y6HGIuHQPodCYmQUJV8pzXOylE50u9kUjOcliK5rdq1ULYLYf3H
MCseKfN9uFF8z2hLmXAaXtVWa5qX0hrpmLOF/v9bZvcuSQI3JhHbwvXHiiqT2IpYjMN3D9TZNtUP
te/lrMeFS/nMbOGoQek0vcSg+dd3b4DnuNyPzgChhKFRxT3DhWRoRatWtSpX7RYsE7g5ddRDmOrS
vV1+vtvIOz3XtgwKusj4yJc4k8xaeZncHws+nyTSmfbIfwCUeHoC0bwOPSVBwAM+saCA7wIXFbSB
BwTL46mgXEpISKsEFu+Q2nZvztkhKDrKQzME5Ot8Qt5nLNDlqlEkNjf/jcAkF8oflfH3yub9enJY
aRgmTLh4ELtFEvOX4RSdv5JI9zyGy9SvInwF2Uzdf8oSO3emsqblNaioJ87V6OPgccVlrJ/V2bax
WXV3J+G81OgIP/WLxUz/U4SVbBhDtkh7hK89DOO6yFz7Se8R8tk3RnXD9sNjV1pCPlY2B+GJWMr9
GPXEKWbSyerZOAJWNPOccczCIcxoE11B/bRTnYBwWqyv/7P766OAtFu5MkCwe/zSP4Cu7kmVQQXo
xE+P+Mo/yLTuDPh3aRCQ1n7etR7ka96K7woGCy0cYqnsFbmVe/mfz8DfKA0TIpSFSk3hcey7TWdy
1WFv9V03XAo0dJMlzIDRqR4Gb7vyfLnlADSTMlI3Hd/kuMeh823icD+xN3cwxoFv1Md3Xdrtc5XX
RqcL5JBVHMO6tywuQ54TGJYd6yB6G+9A81+iS7ctOXScDubpS2IHZGWjlGs+T0lgyE6BTvsbXjcJ
cXNBSiCCkRfbBA91cJ9BQIrTgJvuJBg1t9T9BpV5aGVCcj5q5gP4kZeTzmTp9lmQIsDg5mt0r8ja
VZwKMYbVaPKQCINkvxRRf0n0Zhl846EeKQI+6CwXchizxAE7ZpqF/l4hGDCzGS2phHKqaTfVJxMA
aOXXWq7LaSHj9RhCPEHZZT296O4lnQ78QtA3Ihb55IfrzdVSuwoSQftL0iESx9WOJl40lqmGUbPH
fIBRVvER21Pk6BhtPN5ABIlI6mabye8p422xBNL5YxPfsbUESKdCmtDdRgUWzbgVPqVcGg6SBONA
J/t45Z6qN3gTFixzS8sFAXRWQPGpgDBkcruH8EgjAuGpP47ZQaqilMWYCr8XvBZesKlGFoBAJWYz
MLa0D7tEFi4hbRy1KsDjseSZQOMQlNeWD6/s8df+YWDzcJGO9/925NDbO3D74/im/W6i71kpidmh
0DhcaJLU+U3zGQsCNE6xpxIQOGjHwj64IX916qAVnuS6VouiGCl4LPTuq+Pk7jmcCia4tdN/h5YU
zfeZHjLxbbtFl6/uXd/CYpN/0Cyt+/0H9GkcyDBc4tTRt2Ta43eZ8duwY2GPTSYjNFhR1y3Gxf0A
1prSUXVmtf2OUO44nDEKJXUGOx9JImYrMDwykjNy76el/WBxuI9bpNfIuoMAg8+g57T4o7imV/ff
DoBgXqovanD19ptCB2W4bYYM7awjV9WZ2DidHvULrt3GyxLVIlwzjAKVectOOtSwqveG1HYSSptd
w0++A4lRrZInrMsDz5j0ze7DikylU2Jdn+d9mSTNMfZprbFvJ73rWVv2/kcIdJ9kEynWxRC5+E0N
MseYWIhkyXi/x0cj/gY/8m0vvqbnKW2rn4UTuDWsmgJf6ow3YGfpIY5ohu/vWTzaAus76bO7d/Lr
ReNu1CccZPPu0sE6sjWf2izcYU1qWVYiHmg+PngEIpAudZ3SbrbRdROsmtC88Ud6EbeXEnnK1Vxx
V0mVpO4llVJPjyyi5iVpy4w6Ui/eXlm/v8Dlialj20/z5XqrDtRP9O3Uuxx0LAc9S3PrfCTKbkDG
zeMTzvWk8AwhJT2QARBiDXbCY8Kci4Zrlin9TqAGDeqocLYD3LAfEMY1kInm/dAkPWCUU7FT6Cih
LyS2O9LvrLHam9hvUEGD0FfaAM4C/NBWL3bQakT6KDLxppolveq3kZQIGpxyx/xPeuPexVZVo+oa
GPeJemLfEJGKku4cLImJA5H9G2AFqItds6TVqc5x63nlUGNJ4dgoYar4DgCgE/tksH1fBPBp11md
/yoxOdzQQlqLWL/xT9Hw9unAFmJ/8IErOSb6aiSwoygeFVzKbOtaDtj17N3ZqKxEG1gy4tshQyic
v3CU/Oq/d2G9X0yTlcriV6D41jkrsNkvNCfGxyz7mvqcq9Na72+wISY8tW9TbiTQEECHxN9Grw+n
ot+rVdy9wgZuMisk8t3HQoTtPjfzEFVBn2fDblb3PozDpmhOUjLobXUOWxVqFVdHhLb136QjvA1S
uO6VrcfV7RAXbbK51sWAC/WfjoT6Bz6Sf2b1+XmqV0PkDELGIw6FrSqnEh+41GjZE5JWqF1RxrZM
zuvqJZ3LM47u75XW1gGzC1bqKic5MOUYh5SADbAqKZrdMLRiqCxCouXPkmpj2RtV8v3djsiXlJtq
zrMh+qtuFwifuEsIk2N2IpLhO6m8aTc9aZx60IRlrxGZcvgXd0QMpSkUiqnNK216sU1H8xd3/si/
tZ1WIzOCrKbmQ/IStq5FhSCxwZmzfBiBsfTRreuzRQr3sr87kDL7CdNqtsb4D3wWoSHdl8RihU6e
C5e/cZbtjySUv/je3oD4TolFb0/m8bYGgS4XciYVHz195ztoNwL+fDZOazw6ijw4Z/pYn2vdSGsC
t1jHQnNEduViBoYrEKggqY6eH9D1HIzLN7QfXzusKZ0jDZf62MhFK8TKj+Ziq6MyGw24VZK1EcLu
4TGfPK6xSAKxiiNCu/6VHbEEhFeZ51uKVNOollexTjPwOXBncdBvwOvdhtx5W9qTU7TB/lMjI1zX
F06pqFhXQvgy5bDGIVp5h+i8rVjqnwtrJDi4Fv6MKcNGEh81zlx/yl7E0Z7IwtXr+1WIka8v2Wfo
lLRyt2MNxi93GspGQsMtiOdIM4kLRHriMRP7seZwuKahmFfRdrifBxI2Yf7OEAXb39jE3QIgHfdF
tbSlYPPE4zPw8wMHLgA3U40r0tQCYWDV3T2TjYpntIyyJ/5cuaGK6VwS+gyCr4HYPoOuQRhlGcFM
Rck1WHGch40WQth6N8KeP2ufqEry5SxTRk/ymlzfSrXMxbkK/RvjGRqBy+MHFH7zZcrsdMbLKZdf
/7GCPWt+9nrxlQTq6shcEUyrJMzKynTLKR3ZYMQGz+Wx7gVJprq+7NEeWhPk/XUUzYuE4Mw3+fTk
haYH365qg+sd00JrzMX9l/IQ29+67ilS3n2acBvKlUGdOXlDEtS3Cs/I1istN4A5Hfp9fngySLO8
GoPyOnpj9cvW5H4kBQpgz2Iuhr3ieewLoVZsx7TF55lxclzkgNnJt6XT8TxNtQNpMUrDS2lQxcC/
zRspgEkZDHIy5AGHRO0tjsw8AR+JW7a+Eag9jmuvSC9nWNFRYBH0iz3zWUViFitEovty0Fj67Jhg
N5d4lV2II0zLm2hXuPjxfuqViX9RexIAuBvDQmC4ySda5q32xSVIW2vV2GFnUWuZ20fvD/Ul20da
nlbSL8C9VvusspNdIzKIwVWZ7Pc8D7cZdiA0GPKozOrSmVEIE9JXt+yFK9bdumJh/iCPLbtK0KPQ
zgVqhcvim3WVlME4hADXfbsFrIRrcEnQKd3puewkii6dpwBKoZqQeVdf22KqUB7lZ1FNiTxID7jG
YrFxAovFOSuTKttlpVk/ZFILqnYT/vxf/SVgEiB/nreR7jqvzxxzRG87D43uKpB2Hp7x8KHNqkJO
tyul9oOh2PN5bbTtAvIMNh7mSa+RXrX56AX5KqCtig7FtzTAaTtq1WbBJvxSpQP0JwfMEpjabd0Y
tYhUZuBsVeQsPsmr+uHOd0y3SiJBbomIfshGcwNZLhujeSOXR6TeoQXfDBPweOipKCCUDq/GzX97
y3QHG9eksSyqR+30vOmyVLzb96MNftivZv6qgadrYR57VBPXJADFZ6qre1hGO9e44LLAXmZtSADU
sIohbmWmDDctZGuhnXMJ7We9mRnWC9AFD8HoL8D2qdsf9lsNxe7uRRj76vqhj7YDYVWvEWLJR7FL
JadzVT3FO1V6ccnuGcb/jH7JFVwycVf2AIZqR4mpYU03zdUzODu0jctbB3poVdTnWciiPJzwWVtI
7JloAWCjaKHHiNuuSYNINgDfeR/A9nlA6EQ8JC4JwK7hYVYNIXK32A78xd8XhR1/frgoW6jHKRai
GRRYVjQILo37Bs7mvBWZpiGPlqA7XxkWUd9mIvZRAsG5c0DVicLB15Qq5jOUatttlSzHyqxi3TtK
+YCWv84zq9aEz/KvAM6yfi9+m/bttlgeaepzH0jdr8oHw2XDsUSS2hX4FleA3FT9daJJPBVI8TmZ
8jVObk4eSE1RbcYo3J81imkzhPwKozmAda7p2JQzXrRtrKQbY5dV+1sOpRHoEhXGNUm18cc+DlU0
bzVwbElzrsRG0/n4cpxsQvRfVY19fmZnqIK5RLbc9KtctJRHEybus6LBfvUXThAgYesd5q1qxY9f
mpeD5HqAiplz2RAmDvANArAB5aHt7ONnJ/f0r+uILd3SmW1BXZqs/cGao+ewkwwsc53VbYU15N1l
JSrBUK62BYHmfBd7zIuuBDP4EXzviTDWdsvWamdJ3xXvkWiBBnASpoGjd3/fNLjV4WAG80LTopj+
z0i+eqgEuwSksQQQCCBWSn0Rhjymmd3prQPqasrf0o0VicYswvDi0dN97BvvXVBfYawsgSEw3s8r
YwIMpO+FiVS17EpD2G9/4X3WPvkxAyUJnHGE/YpGunp7/WdouqD8HqyJSLt+VZGo3Ooi4jD0r8wk
AldYXpUmH83ncyx6NILQNMfqJ1RXmPp5tdkO9QoM+R10JUAJOl5kqfY6IQLOo6gYQruaQZh846Ll
6jc+lfzGQu0mB0WQlUgK6/5bVbKPqy6jF31i26xwKY8Jb9u6B6nt05uz14ziI99+JvAoIx1ykJHH
+Lm0V8c02WzR+zkrAI0IK5biG4y4WopVqpQycFcdwG6aym1uM7I9h/UsRJf0eQX/Xe1mSBjai+vm
9DrcgheHlrFZ4hvKa91bM42ImZpdcsreMSz6uSSvZzadtFob5sGA+NEuzD7JSejj8hLRO/oMSRhj
nOax57qCc2ITX7bRcdvr6mSaAP4LIZqe4dMfMG3ZFKalHz3dCuPj3IhFqZIpdU8/XWCZ7Vmy7Prm
jyBpfk0svS8TUQfl9Md4y+qrb+tNYhhUNHg/gU3uxeW5ezl4d2xliFoUDSoeD9GktWaaezXFw2Lw
Io4uIsz6hXL+7IBL4NDq1ZXluo1T49Rr1ZTv1UbCQ4e2rxwRWXlbbwoEYXtIQx+nX792pe5edilP
TCaephv/lkZjdEVunwlr38yG+cQEsXKmd6ZfjlTyzP6zUOss3Uu/zlEoOVyqWxS+ik1Klr3YGuq1
JIf4N2w0gzhYkAY3t2b7X394Z0MaLswvCrd2HqojWwNC7HtrNG89g5IpclTnTExlozxuC4JY8PHD
TUcctUJGjT6WZd945GMMFP4p8tTW/lZdqvHa8wng61LiNIbqkMTgmNBgb2QCgHIGcsQ+1z6iWUTn
3ccH6NKlqKrcDbW8fAmIlvW2RI9r+4ACwz94ZbtcQqUID2ms7fWfMxByvBE5hSGBfghHyLvQUt+4
QIHNAYye2pxgvf3cgtnLXUKnBmQMDi14m7PvC+C8Ui/rj6L/t2GUKon+skb7XOKs3G7oNcShiJ5k
/nj3iSSlu/XAvm3LNtZd4bmdRie2uc8nx5sXKmwNK3mHI2rK44NVtJoKXsZcXnd9jP+b2lNbz9gr
LC4hb4pxjD7vrPGygh+LdilWRLCUWaBsin+K4D1CpWLpEyL5XJq/DfriDSN87RTbEgDaull4E6UG
SciMc4AEoO6gmU9jeIqJJ08YdWJrZlhkCwP7BghKECGjKg6tFEIFzrfN3KMHazx0rPu4LgCedLjO
/WQxxO5G0iwAMfiP3MBaX3ZVRiBy3NUsXXxBHJQqB0hKZQ2WXF/Xl6kfff3Xvsw7u4WpFdSLmjho
6XKgsA7KANaoQWZO5Z6sOYnB3SjPa8LGIzH5JraThV/FxTaELMmx/fabqHkl0oKDh3/UBLdd6L2i
UoyYM+uqlwH5wQj6HHbOgOZGJuthcSHhSThqvQjW3kQZbD0i0BBuk2sluVIuyCg1vSIvRRxdvuhj
iibGrS7EZIKeG0jekZQQJkN267wpSivgdkb3/zHMuAiGRsyOUGT/Swm/gktpXYXy0PHkKLpY5NYS
jfO2zynim1nw6lo5yZ60xr2X7mUDdDLHqFQJAT+g/N3fWvu95o6QFTntm0A23zpWrzo3+GrKgvNT
s96CwjzuYrK4CSd2k3s2I8a7KHsa0TVhrjrWC+qka9m/pGIOQjnM7aHFIlc4RXfscIL6KMq+buYE
UmRDb7swh/IuYQ+JLmPO9fcBSt+eh0u9d5LX0oaHJAriqv2GQ9+CB/vCUYUA7esu4jn8f7bJcu6K
weLHy1/YojaoW6m92w4rdhg3eMaNclPDinOiMqGs0fAmHCyDuDu89ipzkTrkK/e8aOPkipVBjqa9
0xFIMstKQbOlqBzdmp4DTmQURjdceh8AbRJX9erH2/8n1TRXDChaGblDOG1QT+UIWoYzibFE6PF0
aY5ZCUzurZO26q2A0W/73+M4Xn8t65zNZVlieNAd6ZVS/RUbYaVSCc2XW5v5n3A0TyGPBkJij+gy
LBrZZcAqtywoSZA1ohQ+UfjXPlo0x4w9SuFjsRFsAjOEoEdH8XZrXkTvpWyNTEVpZbYfMvk8AvfB
LIQJEdOoKxy0nTpIgh/e5W+cO5lYJJUmU3kFenUFXDf+E5RvhnCJCW+iS3MyMW9Cx1UpDQt4XvYv
kHWkgj6I7hD5J+nndIQU+QCuDvPMm7v8OVh+cIVuDqDQkrt3J0XH+5raAVegQnIudsGaUTHXDGSu
jPUoddYTFLySENFv/5JgwWf7AtMbUH5xUI2QOtbu+hQZ57dVlJ7twToGu/oY7e/dAvctG3Lib01d
QKymLZ4y6IZ7HIMNMt1T9FdPnJnO9mDd1pf7yXyVk4S2QrNTYQgLQ78Y7of7GnPaegeYdZ46ohug
elszWBikjg7DaHXSeiwJbFAlVawviv+LFOzTQEq1T390ox8omUiVqWcts9YHNt0LKlT26fYYaQmG
gTTxzI8zQpXWQwlnxM5FdXqAomRh0RE95XeCBL4AxC8VQrmtDKgBjshLbXLrb4gyJN3mb92MiST6
1kmHwbV7+jSA8PirGqrcOB6wq43aWNqtT6FLVIisxcWiuqJWi+n+sT7ifUuQsWApeLI+tgZ0gZuz
JkW5WZONRqOnCPufWzkk5UDj9tV8CUVfGatyoent6OO3DHStRnZXqKxOh6GFc7peJpfRq4aVNGUQ
4+umAI8DxvFH1YirAhodQzrGvs1BRejAwEqdHeXu6mgefa00dwtNFfBPDs4s0ZLWtQ65AW7OCm30
wzd2Ao53MNiilnP3LkcjAOEpYaDNVQAgCUuGHRg5CY+jufmH93z9ouISq1YiNhCaZRRCaNfuMa7/
kKZ1xCDFFy6LMYDIO/V4Q2cXsnLsnvypbDocr+S+YB/Rm/X10lc17+spuXhTavF0nuMaKSGaD3Ve
nqa1ZVbyv/TDGy/kHAHrobMZtZW5hSg8EYhu0eX+Y3i9q39Lld8+EKMmpUidSu184bnABmQkF5FE
a3dG+kFG9v5ySmWExuotUlDW2WNIzb6Uq3yACsuaWh3o2MpEkGyirjMLX68YlFQBK9F1ts+vpkMl
ihH4lrIslC2pI8XJVnwsaO9XMcl/PYnjmotVTy/EW58+VQj9ulPyCkExm4bRDuF0PdZupuGFzYI0
pT8dOBNEOvdpzNDLeFL5U00NxGmsuOzqN85llwdxOm0FfYw0ALIbd9pSCb0zT5cOKHoIoi7+7MvF
IWqWhwZ1XNIgcVDBc3ZQwiInGmq5/FEM6ylPSq27yZ8CUeQQG1dHjV2btFBWKhRTkX2wdiX36oJ1
yDG0MVJ8AQWBS093AWNsBPzz9jq+y/iXeslW7FC9qLERWZ2mr8NJwtEx3jUm5Le4U/YohCVFllO4
B2VkAoMa3AP5sj0uL1WuIN+Z4C2zgpCF9MCQJeBUdZBlMAciu4ZHi/G1KhmxciJy5hHB5ONeHHYv
lCvUXt2TF3jhK9h5e8o3tJMnpnxf64fywUShnoG9Bo5OtvhpRWx827IPOkqyb2DAsl7qe6faaDmG
ECg+z4UFv8ZpG3geZu9kHDAZ4l5w/Yn59e2S/kNm+O5BHwkFhZJcy/ZvVbuTTUTBLdrg/iE63Lqs
xXwHl+AxhbEf802NiYT/vjecOL2JsAk45VjuGR+RiR+nZPLWvQ6C44BySHRPG6iMxe496BJSEbuy
ku2JqC78GYBIzt8ErusNYJPmQGfEXbHyYe2cbtzPpjIiI5+XRGyfqdQTXfJmhFXShGp5E+XOWA9N
3oyEQDrPeFb5hRw1mCmRG6+5Z6Gd/308BGK1RRCQ9gMgDoqUNTWIDYmeaxxjYiukAc7hxaUi4dNw
nr6ny329FDKGVbe6Ws2Z7hTqQdrnyWGTxuUFyBbf8hUu0oIF1bzTHb6TVwaGnchaFTQHjp1pE5nO
urxPoPz/SE5WwL7UNyXkQlJrSI+cQfMwDf7IGigSKjPWzPEtdexxYvOCnHVn1kRQ5bPfIUIJ8zL9
t3umMP+aZtfce/TdhDNhBAE/ncy77fwEs4ccuKn3uON0MuzrMhL7CE3mSPEH8O3pYYcceW0aIB5y
HrLAhiPTfOkItFpmeLg9mykkinM8srflof8amQjbp0O3wbVrgrjUX87UolAz76kuyNwri+8vy8jE
OCcDsgE28NQswxEPT8WKwGs8GuFvBfU2UWPPY3Gr7/nuR0YMYZEAPlkfWLA7ITNNIlUP9Qv0X8v8
gddV+++K9TL1vbQRNnMRCsRI/JBWoLy6Z40TPDpgSgRoRe6Zu65zsvKLQ5/GDp9mk5ESL3vnTH7S
70KlUIT1/EQwt2rugRK/QAstLQfxYGuOtA3t0A1uBvOOpjURhp7708w0HzGMOIhObQueAjdkf3zn
/VUIdcphEWl8Kw9Q8Y3cs1AN+dNb2bHSZk5MFRutFa7iKPG4U/bo7mi6FV6d+nQthq/FECeapQf1
1OIUrJ+ND3oYomG0BSaFgBdwu2SF2N/60KSGpBYmIbIovJDR9rgK9nKW5cYAMv7YD+Vk2ZxW5G0/
giIbFNXsVakfitFOLwtI3kugQr2YfX6HXVg8LV5EW+DgV1pVa4cQ0gy1bgtSdKj3ZvQe08QgrkFi
Cpk/JQGhWuASbeyEwqbVXbip9pggVPKJmZYm99CoDxhWog1cOtC3IvrUIFuTLjrZfvKWjB3Ifx/u
CAl5reYe7g1S0QYFt9cpMGFzPtguI11HbpAYZuUzJSnyJq4mjpzMWrRgb8GW8TChtOrfgH5qFiz0
ciukDjkJgp8d/xBifXiZ1ahdJA/VSBdZobWyVG1UB3Hnn2NXY1qugISSNzxYPIEhF94T+FQMk5ql
RhmiSjdFTvkymt44glpIws1fwFTBf4huhQqtsevO6dHS85vhxwIq0uEJpq8aUt8pZwJwfrY/QjLc
qajfiX3/+7If9AkeaAjBFURsKCSuq27LkWCQ/oxNxQMSLa/x1rd6ZYsXWw99pi4OP6Jct5MgLfhL
Bi5S0ezck56fkHPaC8NlQKvZ6GDfOXusPmOEJLbE31CEosdtgVwEIL3htiapuzCUNw35fcKhKtDN
/jWztooqgTnaErfVa1UqvbLI8UD6fu+m8nTLsITazohL2Mu15n/t5LSsa+w7ceUxHx+ulEQNpLtE
git2CB7/diO1BBhOhN19DvNECXmNmgsjmV4LI8tilnm7e1ghRSySslj+Z2OHGllCmCHuEJTfQpfJ
OvqJCMhHhlle4SOljm7xXyjTN7O6vLiMEpMedV0pCED3EptDSSx0e3kD+tZJQfEYyOJIk/w0Bgb5
Dq0+8CPeKm76Kl3qpOeTH/WsPdXVh6xUtN+YKuxQym02qNpfyPYBpD/PQFdafN5FCOyjnURdA2Qv
fTa4m2wXIZphK2qIOj+g5ldtuaIuK2Ko7a5IylSVtKOS9t+zuEVdrnUjgkP3eerCQXUJOAvmPrQN
T2Y3WReFtUxkTvI42aOi01YtRVryvXJRSWgr3VL7sx36n4+VlpGME+9AjKELQtNbfDf03PfDcr3E
KDTGiSovfEKnvFo/d27iHXGBpluDYZtrwfOT6cu68/tZX54YHtZD9flpujKZ8rbCLZwXa7FoBgtF
S/30j4ygIWGcz04k6UxgfkRm25AKpJr3b8nIiHOsIJejxZvY+mWveCDyz82Xx1ArSgLZjha1IuKm
Bva0wlqE5PR9gwA5nSHcubYb0CEMSZVmiKSgWHfUru+pV/KKzayPFgQtnMjURUlfTs/7xgou1ebx
r7+UCWFFV0JUl9crXdV7fsffFHTcP05TDBQaCfkL8/XAZjlz1kgBSTMyLb8db7w049R8g/ytkypf
sBWcZe8J5dShx/T4zHpe+lYb5lumNIadWF9/bvpzc/m47x2505elDNMCIR+w91325WH9MZobitvR
qYeBHZG4Xdw2JwQDDVO9z4vXGgYJgjPUybHaq3S9syguZbMMoyfv4Q3Zx7PQ5V+lOMgm50H3Gfu7
7frB1+eRXpIT0nhpEiOukyrakNwvoFg6Cp6pWwjQgxLklv0zUqTvMUx4nyivv/Rcrps5pSO+uGj3
g46+dLkkf26dzGFu48VvatpDhrURKQyPINpCCQ2VKITnSTmIWTkGMh0Pb09CN8LpP4IzppnsExhX
wXGKhGKsyPKMOOf7JoslXiw2wUW28pLOCKNkQlvbCGLcje4xOe/Ug2WHhY9400LVcJSXNdTMUbQT
yIALo7/xgp71yhrcyoslyyALvHq8UZMrJ/yuYK+N6wCvledtIOblJIS9uP/qBcpJFIdTuyFffqgK
arbsqfngeNWwCWj36D6d7ag4qZI0elyBOaYu7FzWSgEOZHN9w4+Cz6ES69jnIYu7n2yIHx1Nm48M
v8DyeowtNVaqVl63PGMQSvqvIEBctsgkuhl1afVTC8ZLnycMgdnkgxXTz/FdJRpVCEBwtxpop5S1
n0QyBNOtuMoXfTLeBnCFfHLuCAOLghD8TVs0L5guC2gYuG+QK4xXYvPxW2aTFHUXPvrehWcjM8jF
dscgIFDhnLdxwCJUrzNJAu13EWwZmSZR2Jv/R6eIj3hONYFnZtb/bc6ETJM3fClYUQnVqlVSUcPu
ezDY6n/aDvC6QYmoGnnCIJyJtCUa5gm25p69ft+X/3noetfLH8Jh6c5v32kK2V2w2NQSYjKxGgQD
Zs3dI2D7oFuqlUGzycPrVokG2UmULHuHMuZIVtRxenJABFMZNt1KCtfR24DMMuLJp6SerPlBlEYN
BCS2f9J9VNc0vcCtN+6/d0mb9q8OfQ23DtPeFOWjUGCoy+d9SuRNw60wtna5uSCR2M1WaeQsZXps
23sVRfhXuxU3vmL0ZU4lmhwi+LOp7eJMNzvkl3P396O6sOQ1idIkYYlB+i4VHg2Do+Y5skDm5c1T
AmyCRit8/cPAEqa4GVg6GYl6ke0z/aSiWSOtbkqKewfHx67SEJ/sK+LQ7GdiKRz3ty2wAznJUBh+
YVm4uuYH2MZMGg7+5fj54dcR8ejs7ldWx9DBa5gwpwZesrD6L5EQX64Dg8x2IVUxmmbmaZqbrE7V
oVOa81dIlkfHsXTMFzDkPUI3jzU+y/vlkowlJEBEnSmfxVNSbN1gU3C/cwDG0LL/vq4BpREfdaiW
vbcnIj29iNzVgL0af1dihfyTwtu8Y+DCUZv2nTu8+KRpzurDJ2/9atpuTd9VT5GP91e2sFpP/UFr
wAJZdNgfEUfUQBKqYgCqF6O5OuQoD2HeQROUcovdm4A7c7lQRn2FfEeMHGNdkofRmwfO7orIEW6l
sb2H9xIlH7HkqzXDwNnvM/Z9ypFYrCeNFPvu2aaWQmToiZAO/lhhokp/wcAAdmwLybLMUkFFjsG8
zi8eWMKM3SAZXwSVJN7ZutW6M9nM+QLKVWaV98gRy5QLMhWdszXLsnGw61BTKMkgUdQh8zH6UMP/
IU/AY8zLc5HABhiyG1A2eOC9nTdztK3wk8KQc1KUglwZDSjcTkc6vA5xb3DLv83toFthfjTcAUKp
n68J1RDZpInEENKyGDmgr29YKTTbvnzdg80WeULd39rtYb8oGcWAtAuPued0mcrcX/QaMrZOrH7M
VVS7G3P1JnAIdu7JCjgLRUPOSTqhOr4gBnKUL8GIKoUtcxF7R/Gif3lij3PvGRRyEhvyaAfhA+4t
4WV7Aevst2s3A2fdtMy3blSIuHRWVfdajmGRkX8UNCXE6pzWVNNCg9TCmvXLt3UPl8YNtpP74f2k
unfZYvFaHBMA+sHn1jjTFWVO165aStAxnoBFpU6lIQ0dgtRnqjNxkJxjnPbFPG+4CxvcdW4iioCr
0fXmmaamyiWB0+gyaXz2/RQMNCS1G8/Dv7DFrooGEhkgwONECy9e+R5s9vl+ScAHTbVMui3D5s1b
tv+fsJUVetDcojgIP3WpsV3nw+EHbsffhro19b1rHv3nEgCgy/nzeayG294+4jG8oRT3QlpnUYOG
bEx8ka1bUHGw6GDtl6wp4uXT/kfxHDwBagy9+WdmeQ5yuhZfBx872Jy1rdFVUtMcFSvknfSVMfSR
If0X+3zQKgOTlZC1mBMWbpGjfpg54X4w5cd1jj9peqdWxOGV/DNaCrvGEK3pcIsF6FpQisGPcc6Y
++mCUzgglZMngGcJCGhpDXplhw7FuvFus+dPh1T7JPikj+Ycb1/PK3mpKNhlmKstcZKyHvAGgqLC
h/zRobu8VRUXlHzMzDxdoSL3noiXWx9tU0dT1h+gZDBucU106CvMEvgHRjRY0V+MJFnMfO3abSe/
zAv57/KTDvJ7Sd4WgfgjleKq2L+HPuqs5KmHS54y6QawSmfHLyOgoFWgCUxVL8FT4FC6OYw6+bto
KFARAob5gioTOfosWrvUBM+du++Vv70cJEKjlGHLQoFh5UJ7ROYCNlqWBGoJcZP6YYzmeldFsfuz
Ea5fR+X0AQr853up5sba8CTTW+r5c7f2jQJ+FAXHoW+cWKSWVQjNNpDPlnHN18YilOp+0eBOgzvJ
SfTpRUc3bRrQHOjNHWPvF5U2LcTBkF5A9oVm8W5yLQLisjmParGiM1RZ2N3lulSEpSblLc9dnBqY
gYyXhYPzZZSvtTGH7O82xV0gj1lPAbE33C8K4UDoi8D0PmehYLDtarPi8mxqlpgzT5rhGV6L4p1d
Bwwuc7fhx+ANP/M+iedA2vFhcOzCYphu8O426hh2HKOqRu9TaKipp8OHQDcHFm7FFOigJosmVCta
/siT0BOOS+VyueUiT3q6R2zqkQkqSJBAkuLB5C0QNBynw1phplh1sWJEDCRzwll+lGmBMU5IYpe3
ZJcTl42gOMUo3s+uIyis8yC5L+DmUP7lpo+1ygKhweHeauYkCQU1p0j2xVESYXmki3WdeXDldzpV
cFMJlvOCiknjb94de99mWmOzcndyUgi62Ii3HnSZe3QdnCdwEZgNSIcTh81mICPfyw5LWsZeYGiS
E6UQwm5GkNvNtHYp01FKfwGj09mOLqSESCc2kpIjqGJGJ+b9qxNacVCvYjkBDpDHv6p03sHyjLlZ
nOrPrpGhe816jGAngA3YkbSd6c4pnS6RYsn8V8jtg1LfYTNeibjZ31LSBTUt0TPla1VxInGwJoX7
Poo3hSLQfko6utrSpMsNDxMgv/yspTLqDFpp9M89LuE4F4sispNiHP5Y9dVIo4eHr1zRwK31rqFk
6gS8LzFOwQ+9EnfQue9+EHQweHG2LE7xKvMMbj7oYXsU3e8Aw8BHcT3Ny/AcD5iHRLFmBpM7m/I5
V42TO5cBSKjNE1g5/aXdMNLI6bwylqVlKfcBfLh+MaDP5TTWfzTbt/BNYkaTmVnYxs5muvwlYHoc
Lygzb6B7XAwfvsqoWHR6TcCZdyRZKjKyFHaJS20uavLxxhr8yff3/6s+SGdi2TAUNHTq2mqxL3oD
XFquiHA3dYn0GcC9B4Vkj3V3655+KXvar1V/r1FNsIhV+LqPjUwvMugjDwYxKq5quz4x8/yVuIw6
fdIvgVV6r7Y1POB2+D6Pe6dFS4lv5tIZsn9RShG+sajlcT2CAfyFGJU5M+69WNPRBDLi9vhE+L3I
3ax2kp9RqiXi1P6ghCWKGDXYY49p6Z2X1dBaQTvV3yoBPbNVprG2EqyEK+GdchCuRv7gqrwHI+E5
0KrLOknsDD7EKyPYKlp9K5+1nCVpthn+dQBJgkWzVUMrvmLQ3I1zSPkmyEI8INYvcb3iuaZHH5aH
Kx6ybFjBPbLbWjdgzoxy8kn3tRJSPYfs7W09i/xJRnklXgoooejC2ebpVy0eW5BikrVa+jggy/ke
dayYgQF+CwIhONdBaxFNDP8rryHdDsqQspUfrLTBef8cpJjrzLMyKd64xS8ZCm25ZG8WIQswkssT
1glAOEY6M+8xohhxqdFm7wXceu/Vk76mMuTErYQGCR8eMXwS8rDQoa3SM2NBigyIt3dt0znK/wVm
b6MMNXNBeOgdPB5k8jO2yxcPje/kpaYHKIUvoWGYq6trBOXkeki7PWWQVpQNuC5RoUMoicMoK3Xr
X3yv9wvGBCjRhIAdkxJnT2//DDsLuXSS9ApmNY+sjAGSf7Qs3AKsHD2+4qlqfj57lfJDswjve0mW
k2rRMXz6Tkk0fDbcKwBX3+BgcDo+2pNsdgNIHqr7l6jFeoA3OSV2G4byqiahx/qzfKXlfxHzF0Et
VX8kvIJKmlHXmoV0ViIfwIOjgKmSUU0Kq0Bks7VPHegFOGeL9bU/7QWxJ0jVEHuJXjCupJ6zJyw0
AgJ5RUX5CnNgbOL1HV/DxVs40W2AyI7KqJ7XPCU2LcWZQnZ9Qs4hF8hRcxyDN5VoH59ua8r7XDJu
sWlynI+FAhL5GzZ0Kn2hrKJa30MM1yhWXSZP9RbUmdIzXkSplw1f94GPtAlxZLyA61wAFoXsllyd
6/N88mBQtOV9OcfabJDeJcSwO222VJuy80hVSlOFkiZSsUD7J38QFhNwOGHH+GmF0zAdZ9BTtk/0
XuOVTIDzQqwvxhzOIGbM5R4pbAcMN9RjlCfjSXfl49tGsD0axyFd+ZNuhrFF0izMhukTEHwtncvo
GOSt8ZkTajSEtvRZUuLgs5G+ba4DyyaJLyRXuyZyUJy8EnF56N0iluXkZ64LEAeeo/rTUs/HOSt0
1l3xQcRwB9knVe1gTYvSa13qBRiNFzx4Cqowa29loxOYTCsJdGR3R/ikJrfmgjeC8BdamSsRZHvb
IKc/mGfgl/tOlavDgztpNu2wjWsUOyrxS+cCrYJzatjGAUZ6CC/cPsYS/KPEzDxWnJKnEWND+iWG
lBgwL0SGJrs1FaU6hao7H713oJTG8aVcdXmpPOx/KEVbMivfw92tmZZpxoFN1gvj2rlVvXVgx6oe
9k27PfKLBQ2AWDU9K+2NefmqUBzlIxD3VazuAF66BOPOKwCH9yRsROyzvAIjqU785qHzvV8PfPGP
dsOr9EGIXY6ScH6akszaZ/hUjOJdvP8d8ZjJ2fA7AcXtylXW1en0QRJ2CILQ2Ma3a0tWwtGX47eW
ESIbyMkJADoPk+jWoEEM5oBErvDqBeZHsIg7QGVRY3lu21XzJtyq6P0h/aTolR0Gboddm8QeXPtw
JgwO4OqL9ryrdhmJxpXkcvAEbSU2jeHio3/Ho4sIooMUD27CfKs6KdmKwJkHN77E180vBd8pkHma
VWwCMfOSk1eITbHx+EKDBqBw8M8z7ARP5uMaDnlFlNwfyG1fY/ZJB7ckm2RwbZ7LE7UASZUgqgZq
Fmnp5dDQhf8dM5LH+7p2+DqezMJG0ER3yk+b4z2gmFIK4CyjjX2ETfIofqJWW7ixD3dnV6RMI3Oy
XpRg0NsHm2a/XC984ws+cFMxYyd1CSn1uOLPoMq9sUe5c+xCoi/rihMVGBHrEcjrq2l+Knwjvoc5
wlKj7SsIbpEwElrpRy+80GfI4eL1dv3DlbIMs6SCj00BemIXrVARdyA+EwNXG7e1rrUWnQ8DIKSb
QkhxaGbFBpxEIMnbEZbunKhccUKKHaR9j0Zf6VyID4umAn3WwmlgzjFQkixkPsylMfQuIYweEtDj
1kzPUjCxBgSU7aRuuuu+agC2OLBSNYbGUCipwSKY+5XvCRQYMaDIH40oMvdFY8VUO6mYk7eBggXZ
PiChpsGV1uWy3YdpMFkFpchkGH8qCFlgu6nG0nEo3QCfDH7tRpJ/8xUpihV1GTIc7UhkLMJkXiWd
0pc1Uj6HI0yQkwhCecABZF8BqPbRrwn033ExRv3lc+t/fcyWUAH/vLEC66GaAKL+rABbdnOG7C3e
LhzvjK9SonfLelMH1JHiyb19yC0pW+cDVYWIe6E4IJA4Mmdm+M+ypIOv5JHCbJkwntR6IhTjT5DJ
MwmLg3sEpZZnNLAag3bZ3Uqg88nJlAbeqK9PTdF1PdTHhzU/9KF++FkzzszW59hgvGGi2ijRzVWg
CG8KqZGrq51OVOtLj1d6+p2pp58ojJacnr2eKYZyjQ/EfbfPYF5P8NH7PaM0ip+AXEnsnbsPIy1k
Kabio9+rozkqrrp7RXro83l50KJ9Q9N6ejx6J++8qvFPZuz1+aHHY1Izn9uHbCaGeL/O05aJhmf2
xBpzEbZFL74v7n23asVsC1oyAxA17/G8RP2OEbNl4goqura3pZ1CKiKOs/wCKWCNvahdP5DM5xDs
0nBxOUxm3XkTBPJbQS/TjVPHQMLGaP/tVvoWK/LrUvQnSz0YYiH2/D+pOrvd4SzLYvlX9EUbB5QL
1LssoKcjV0zZ2+cIWFHJQhhVaZSCAO8nKLRVb8LU4C1bY6XlIKu7A+qq+oqiYyHoiRikz2EDyJmL
ECODAOsTHq+liVIJ+FXJV8099EsJJdIToejZgdD+K6ebDMCteZ1MWk5PL2oaAmWA/nors7ovUT8G
ld8QiSWUAOgZ9Bh/qrDuci50NeRdFauDXAU5cagDY2Uox9EWcWDJSfo5y/x7mq4ARBY12dCVaz2/
n5IujGW6fFKv4FwypD86Pmc1+X5LS6rykoDZM3adIdiZ2P1+dbjsqKYcS5RXrR+v//GlU7+yaZFQ
KxYn4YIpfekBBlDoMuE1YWxl8DkBkdQMvyFXea8dfosYt1kwTp7DhjnIxf/iNvm2t7F233eUImlW
9mnbhmC6449KR1wZrvK7VZhQpls57cAoXlP/SghNwbOKoNv3o9vjjXLzfmU4gg43JDF95C0b0zzf
B0fx/yp9MDBlRmvi81d3TBjf/Uq1hIJmB9LY/4UQ0xDxL4fPvidLwzF4EB1tX/DhRtqRRsy+CJ69
tqrNzvm5PJZegUo0s44BwMFio5Y8t8JA4wRA9+JzsSLcAxgnjylMzwjw4YdebRGSgrUGwgcucVpT
6b1uCXEnC/caKxvKDCbF8CG4DSduJzl2KvDj0Eye172KzajKL2Hdte88zRCYuDlmSxskxThMK8W2
s+F7FIN+izW/l5pGXWur5JOOp2hrl2vcMYasUG5k7OWKwdVrefbrxdSRfLNgDGu4usIYpZqUaN8t
zpYkjzls5781Zw7L8OvArbMt5YHLjg8a4fgQc3dc5wz9nOAhU/2QdsFxm8cEgsKCdqJ6OKwIdNUy
PB3f1qimqFIsTvrqeHKZGIVEtb5eSeFwAE+lkvJn/dLS6XeI3xf8iqibVyGtaEKJIyU4ZuM5VF8T
noV5nlhWbsbOdYxaJFq+ufe0V6cLaek0n7tEyd6mrfPa6Zt6UtKIf1tgwNUSJ9covbN/iYJnVXiP
K9sGx8VNp3/mjo0QHpG7ZMDFJ/hx9oYoeC8WMpgfDkK3/2Q4ePlj8MNHQ77SvlphU76FCQtoQoCg
qnM9JviTkwfV/LOFp+K5h9i4OuRpyljupEkv51sZ5yyzvLGVu7v9gAH0fvOhvKQP6j7ZccTHY8wm
DTFHJF3BDd6rub8G9pYAZHQmJm6k6aqkOzPhK+76K5QBKIuTXlkXUkxP1olkOL3toStLGlg1iHsi
tO4hB4dTlZhKEbsGqFXtWHGT7vvXE9/IR3tXXxIlhXnpJRb+sAwmgExxjPpDCa8hmkoUqCWowr8P
sgdvFJ63dyarxq7SBFOuNk32fi/4D/YahGQ6YaptED3ffGptHpZDw9seXugBM5IDPNSI663Lu9yz
fNoBU2+PM+Pugnli/XC+vRJt8hOUwWvVQVRrajCqQCZeRyxzHEk8MM0YrQnxjNp/Gf8heJrxFMac
lt0jvgkp2QR9/79Uwu9L83bDmBJefOzQrWS/lu4t37TVDQ9L0hcEDc0wL/75qvny10m4biMXY0SS
/bcOlr9JuDkz9I6TzWfXNOJNZp2ChWai7Hj3g41Lp6mhbwiYNwRUOs191dcSzV0YnIgdIGu31Zl3
VNIH7YUz+UuGQAr3bRqDRHXS0ooDuK7XoQWNdeTChgkpNbwiItvSCAfiedTDbEFnlguEvziXTxQo
qQj4O45cQlX5lzPSdIFNTkP/HxKr3+ZaU3F7KHKoTdayvhV3bPbbjBTzurJtzHg2oxQ82LP4q0fG
gqF7BtUfTQBUl/l9VQAMv9ZfNjmYHE7vbe1uyiWBsIxkkzdBzDYYgl3ZcxzoESFJ9bmw2rxzQouA
MAwtCH5XeRGLLSd6tu48AJ6SRwkDGS2TVfxbFI8qrndFXY0Z1AcXwgB7pnHqtlnG9j0oe/fRS/pc
WNrfBAZXltu0cpHu1RZTrCEB7oMEPIdW14FZl4w/+SjJDiBim+Vil1QO/xTFfrg2u8Ofg/OZYk4i
KpZThEHzgx9KWBGhC11nU7ZXmfLmtLyWnUW/NsTpa8TgBnuflPPEihqpURXiCCGz/f1ePQ59+Bor
c2kBhDFrqpF2EfvvquWjKBxyTdUSB6h84JjoOLO7yOH/pRDs6R1VF7qgPN4iQpzfJbmK7dK3f8ON
0GD+0tDFO88fWU0rlPZtz/WnWzhV2MMscYkhg39bi0+2bprRcnW0Hy+jE/qQBcq86lQ7ho5X2rzz
pnoNA0jpDvp3uRLl6C6OGH1yBTrVgFWbvhGDSS+NqAmDeiI06IPQi8jmOL3P0JBrUBRoVluQugwm
Xzi4D+MjdOrHydopqZVRMJMdVZxQbXTsLb8gT/TPYDb9St3cNEUnTvZoXWNT16b62O3v/kF8XUoJ
zMws9Fb4Fii4Q8xlPhKKdqrRUgbtEpMBUl0B1Xv9S9HrB6irP6uqY+9/iN6xaiOwnd9FJHmFX9NC
cOtHPxm4E7KJcdD90clfvu42jbekaQ/9dINGe6djKB0owaM80JBNfG9KkVgFgN7xl2GNQm5nnVRX
rV9EU5MxYGE0+LHSlKZxjY+Oy1mszwxWSj1HQpsY6vzwsDyx7Q0ntlr5gtY3K/vh2SE2iZw6W4kd
SqwADh02TzF7ODjZ8P7HJaKIywJeHyM4Kcv0Ihjm/PIg/b0n1N340dEwwYIbLySehAmH0V8i9YlW
np21s9gG2Qp10LStk1Se/YBnIifPjgntZdMhaJR5jpbi4jMVzJ4q3KyO2XiSg64Ec+vB+UMcS3sw
NRMjxYlSD3z5r4f15wi0oW+2o6MpgTZu8BPwlS/LrvIbDVXH9FXqs5hcwHwx71QSuaWIZrn+U9i/
IarPbGHUU797HVLkjLy8HJErdopTtXYzKlu02JN//mL9MTxuybGDcl7gxS9LAkdPE4Jhl+F49U1Y
euAc0H1orhfWhgBj3U3C94/RyCyyOwtufsBKxdnmj1v9lX2DOxaxpYJy6z5viBfEvBsTtkQZgV+G
2VIUhlUukXXieRUR5dCewirerAiSCMuVJO8rZgrSTYWW6nkwRoB/ZTVbREykP+xObJduC6LiO3q6
t/yF1ft13jNEjI4r3I3dD1ibDldvjnwBNDld+MigRDaSACBpXU+M1Pynp1uNXRmCTQfmKmMVCxX5
665F3f0TeFA2tnGNcwYQ/hg+e1pCN09/3DnUWbUoNGOUEIeIB+OebWn8If/3SjUcYpkeQVLsqtW/
LvKTesGiPMFiou5nqlcuiavVzQGcBKgbExf6A4oI+9NfQqhrEtH9I8sCiIk0ZUIQIQ6njISXosye
zxCga+WvBlIyAB6U4rJ4tL9oMHXxJUtpKAqeHXRpKWQQ7dBCXSLN4V4R1JjJEUsd3Q6XcmTWpKbU
AlF9sxyIPWdtV/nE1KGBcJnTGiUPHWE/lebpj93ffx142w/3ShwfNO/aBy+IsWjF6Z9Cf/AOIZYI
9ZxNVgh2MAcGawcLweP7aCwhin0USwXYvCa2C6AwjBoGTnn9bFm5dh2uYYlqkNvU3onZDzOF1PAV
XXmkkRI3ITXcqonHwF+KCkmJUfRVSkOspq01rPb2O6Z7n8hOQILvIZ1ZbczFNT6Tu1Qb5pu3macF
Ls/9yNn2SyKPlOXm0MqrYwGD3PlY91iq44wWaxepdmFS8zl9ryBwGDGeFDm+KzmUrKOESXwrdHri
l8Gq/YYGixmlH3iNmVQVUA3AgllovmBt1ZPMJV+ghTo8CgjPfcFGHddFC8zH0pNpErtXbOp6QJif
RGVW9o7x1ougJ6oOqjRUXPNGr1UfT86oSnSZJera9WgFStKIUdgVPYm0wBkhZU3xYBswWxzSEqKi
/HmmcB+VH5HI9UZDqyNblU10Srx9VFjO4VPNvjqbaw7vgpLESnCloYbFMqIJiKsefe6oOuxUgErI
87i6t1PyWbIqu9fk0hboJRaG0Igtq0Lkmk7lQqbZsj9/o06Lo7L81ZqSzQGQCKZornPXWlgueUe7
jgj5yRC2UEZq2fEPro2lMsouO553KadR4H/p3kA6scY9inM1+OTxCPV7CL05DryIZ3S75yB3B4bJ
rxEm5KcEZL6kfNy2Fn0GStla9wHT3mDow8qZTzIq24jb/RxfHYmlLHb7U+KHyNNg6L87ddUhkj0W
7bZh+6GPihtQMI2aiBTzwciUdoWKOaB99nU/CObeEx/dydIftThmSNT9ARlGYzC0XTq3zfgCOfgX
Xy/WHCX4GN44oLoPm/WBvHrVuYf6tKdxjWSXpfs72FORSEAxF2qc2U3NxI7P66bXgcOQ+VWZ/VEO
VCd7FZJeJGEnP/I7zEweIHhpkS1bzLxuIXFLTJICQG5WRP8IryQDORN0JFz8PQ+gpKIuCTKPkPIT
wxpVRZC9HRe3l0zWN/CC5zgRyUmw1bNMu4PbDn7RfDUFRr/1xq6Ky+DQm/tCDC+UroKPcbg4g9Au
me2xAGG17KtBxT8E7SJhkmGp28FgLfSGvK0IBZcZO6IoRyIguDJ4M73b8sj4mveS7UQaInAdhkVq
K9Br9UL6WMqSBOF/rHdQjNamMhIbkvPzIplb6a7mqZhU3yRmO+MpKogu1Q3sQbJfSRCZ1jeL0oIU
RL3hXz/G5Vr1oNw9NF90/RT4iW18l2IaTTuHjcq0ecZkiICC4ZsOUGcEs5lwY6h1WOYslnjPkzN0
7Srz/9xgf5Dmdj5sDE5AWHJX4uiurH/6JeebrD9stiVyxG/jY823KSK122lZQ0dTudav6rL04azr
0h08GnzC97jIMFtDyXJWjli5uJzTTByaKaQP3OLJpTyI8r+tH/o4TYnH7vVM2P70EnPUpNVKv13+
nioEsany69UpI7uH4/Rs+0uMSE9kKQMGqW7XxWWk1f9YPxsoTwhNPpL+a+ijGWGicAbY6rVKJY4z
WVf5v9Z1PZXV68ajgK9aXoLWezn2IaTyY8A0rW1YYaNAxXwrYqPjcqYLmiGefkFGR92kwYJaOmZ3
tPcApMOs8t8zZC+A5VlIkda32n0lz7sNCC0RyEeLOteG4Em3cFTVX/q4GIyVdLZ0UHsBWPRoIcJj
Dh9SGXy3bgjQ+Fu5oCI5JG/kxF+Y8g5D2ChMcrfuWIr75YoWIVuxLvNjmo2hsZ9RSmyg7Xa+jbQa
NyHp7m8FZhyPaF+Zf0Vkh6rWdQamhlAlxLlkeb+R7prNp1zzIlJCCbz52QXAYDNlFNqlcwoel6FC
aa0mwj6uEv3SUgVKcfVBlYY/JPCs/+XUKFxUan+1Md4T6lam4czem2F2LEBPYLHALOIqO81VtPlG
+oU0a1RpFn6StB0R2WzkmSa9W/OC3jFumH61IA7CWC7WR2LIQaIVSD6goPNfzdYM3++Bll418gQr
BmvzzUXkcqSvRxOJjb0lX7UFlcPnDPI521LilHT0NmFi/J/c+fh6XeobzF5oPM4YjTRy93d2+Qos
7mGHJrBIKAFBplCbgnUGxjxZsas4jW4Ss1QroXmEFduDlELq8gbUVk+pkCrAM9JznJE47kmVdjE8
Rc24FU5lFqb9yQA4urqZ8FYix4unE9fiTuy7/p5aGwSWbh/VLHIcSXtDKTHy4MpXFhyjun6KtHXY
qVq5YHhndSfXB+ruvHlzgfAHnIJD+ARlYe+El5YcwYcHLhguhPbkY1+Sq2silZaXz0nGh2Od2DGI
eESdoJSwWdTO64XrIKxAZWUps5L6Hmwr6huKYgRDEsHU0qseVGmuByrHSSitQlzyCk4plIF0Y8dC
MtF3FEV9Hd+RZHEugw/u1hL3CoJ1SYVZJIH8sA6R4DvxWLWcPKvusBaHq6mMXncFBmPglevcns5x
7/pYiYqKvxF3vjir0cnDqbUHiVBVtzG3MvC3OLt88CNFYxXX+aWPcwxJ2hV454zu9eWyEkowhFk/
srMAC3+h2HE7eltYhYLhA184i8EeP/sJP66pEsHCj4Gq7cATLHBXSTtqx2GLe/sg7flaWrNqYSc4
Zzy8tDkYGseAygpEIwwEVDzgxFM27FnnOuBU8BLJEX9/iaMHxc5vp0xaSsk+m82FgCg3ckXg49WO
RjggP3gybUXMe6otn0JRLvM5m0KleKUyqx2txbTJUJSGya+hCykqJNCpHkjg5ZAC7EBaf617efua
998W9h4QEW7Jh12OyWVfmoGSD52PDog4JevJS/82+xwuBEanPOwseqUxDNUyn7+0UO26ifubtQ8W
FGRHSt6SlrKGO5IupciEfBUWwgcsgaK4fKs5jYMgVQCsD2wZ7gfpVV5eREGizlclakfymkEAFe4v
TBzusJ4aVuIv7U3BHCSGvrCRBdzUD1T0vHGAqebtrmO3JF9+VZqRgFeVZQ8MIpWHd/ZxSPRxlY/J
3Y3uWwEhiv8KP/8XYir3Zofg33zWB8fDgvBvQdpI8pDNgfcikSzrGUCtEDicfeQ11NV9ownvIJTO
WSI0LkNkzp9Vz3aWAJ6Eoh5QS8ml6HZhKdXOTwMy9IsVQWAnaTUSCNq8waFkod8gEme0pWk5kOXN
NBQUwdaaKuq8Vb1xPAd0W3a329ltBJyvPO/08J1ZGdvdsemyqPJWpUwPQYtfJ9xDywwzieqIg+BM
QsCWBnLz3rE6DPJN7fUdFrtowygqsMI2F4K/pDZc6AuFwNqh0cFZ5AInqHih2uFCmehfHdlmkuMv
Ujye+7dsFiwH2mLtFoWdqhkLj0zEmMlzPC3BNyazVVPbNpVjCzkJw5pqkaIx5/UU9YFmp8vqcUcy
YMpAjsVx1ebsc3qT+gTOQLfUjHgbiFhyME538UZhnUxBZBJtrQ5hW+Mn4T9e8AeCO623kgwx3fGf
GyP3Cka7OVr3MHzJWVCWrlLnt1Jyh18sdn+aARE1JTKe3Zs+4D34XD/raT/4l+Ju9m1m6p3JgK2g
lFYX0nEuH4RPSG6tvh2a2WBtDVq1FlYQiYiPN0Z9wCXcbaqMO4mxh/t3zZkL2GeH/xUYiph5hhxS
t3xs30OhKdN07sNw00/sT1t/1glnjWmLWUqXqBqvFVsR2msBRNApNjdateeUhDUgOcoVwiTMB2qB
spjigW+RRrDPI85lNjdva66GUgUuAMC7LNgHjzwusWu4HBV+eRq3w0h0V7K21BBc+oqr2kpjJHXt
4qqVJSdRYHkau5eaMbTY9gde03FYkQN0JyWHSR86wtpT1AA3CxKfT8s2AI/NseqbYLZLypWgPTlu
MqbVy+EjsqjUjqmwSs+FczNQ2nDP1+8wN4nGZltORyDtQGfmTTPu3Uv6XaHMl/8mXB5Dzs2voSxB
sQxdZKFqU3TGIbzUBPtM8nmxkxHvPvMad/RxuQy4M1CQibzbQomyT7KUE25HmzxGaL9UVi22qIw/
6Nng+di0MCI/xXSwfUplKF2+Wj91HuS0Ww4Q3+mLkzBMVjH+lsVaFXkOp9+2CPgL9CwsKpw/K3fY
u3WaSRFv6gUmHfMI1x4eCijSyFbIPmJDShuYg3lLADl3qBv8R14+f2zPBUxhM40wOxhZm6cXlSEz
d/whnBNtp4OOUIBJpJo+KSaCEcFTywSA8jfwb9YS4d1amiwEbBJsi41tCI5GqxbIb+mVAN00nLAW
2wF71VAC39sDMBpFeLe163US8tL30dHkusmBoNPQlFDxsDfpkLiXaRGWyeyzFjeo5WV8apQgZAix
mfbrf7hUPjNuYvaoXEWCFHVQBWAp9cgeDJiN8UE6FHcsLMmVc0ChavC1V0Nt0St46LpexIA857oH
U/ZKFHgZeI9EOYPNwzW+KA9TZBmCbwaM9apjtIlN9VPKnfl502Fiszn8d1o76cjC1oDYh58yfmMW
Bbx8T5I+TE/dMASf9Lednf5/7xvgQT17Htct1gBCfcvMnj3LOnaICcgkFZeDkmF+ZmeJTTn0zBuj
phYunxKl4n5FhrCVvBTGDD6KqEL/+VN+EK3sEZSaHwa54RmX0n2ILiC5u+aDcH011ap5bwXqJ+tu
+Rg5ndtlkm19idrZaGzuZknqTp99dtCqeorosjB/S7mY4zcOO7bSKDZK8+hBqqEFBjaFmDsV2Nxq
Jn8RsOO6PTKt7Wke2ijSrNAH5ZyeMmWgQMeD6N2yy15LnAVsVsn70YsC6npdMpsHg18JWbRF6BsM
tr0SufoFZZzF5HSrIbFfvCAt51xwpbbMVMiRqCRsvzyauc1f48bNEBUgyowGB5RMgUfNRfGDMbj9
DsE2Otb++wjgVPMP8JgE63u2U0jhZzXSzwJ5uWQV4sMHvGemHH2ht7t+8cmLDsQv9qrghjjUvxzI
AGkA8RqaAc1S2Z68LPVLZ6UCFnKAO1aYW+AAS2Gj6MUOa7LORFSdyTF8i6b6MmKv5Yt8wG48LxfM
EAyNC3YMsD7LhVadUqj3t6ktyDWlY4qRvpEJtAG1yB6jUNEJ7J+3djGlSZYlrfVwVA5QXSQgLIt4
gbTrjioSVqptAAwZEPCxt6YtfxDWFPV91WBGnTaObFHia5gYlyRiGVhRMeT/Z7GGRLgaRZy8A1Hm
4oHdITE3apQWNeIW+iJmW8TrKxYTp3en+bQU3PWnau0W4v8zUKbl6uAUoVsSuJRSjN42aY0V5tWb
bVKToR/IOgib8ARFKoFn6KJwYqDJuoDWismOQJD66xk9v/zcRbnTlW+CmeFD21Y15ZpNRqSUhcyd
8vofPbe0xTkQoFNM1PfrB76elAUJBRIwmQ6w8OXTX5JaUC//rj6qAGTO62ciQO5cx52jLlnHB/+P
PueJkEh5yRNjuCVBzIl4a79MIBmY4WP3VR/QVXOJLyvXbpGp4UBlNKtmra6FE6x2sLP2E/mvX2U0
B5X6rDdh8YL07jHVi9YmdUWCMPb/doqekgAaRqb2iF1scRpVFTLESTK8jDApMvOmnglq2fOyoixF
0qzJc/VA0IrRlcLiWmDpm1t1JhsLsWZB5vrvXjmw44vZFezvG4fXsZAdJLLThwRE2V6ncGdu6Lpf
Qut0d91Gd29/JWS1OTglBC69j7h2AlsKFW+ddFIftUjqazifODoDWle6dC6tOS1Ds7vAaTNZc89B
juPTAy1VAwvXyuB77p/MyMtCcf7Rekx90RViOjBJNkvebj3Y+/C2tX/QtZ/CQyUZQWnFPlhZ4fL8
SXKllZUgUHHK5INcCut2I+Buu8Ww8DVxEdtpBBkNKS/HHL/jZ6keJUsEX3OsSuhygl7op0y5XtNG
nuVdoTz5IV+rPskyLUmlE+ypwJBAW7+9IIiFUcl4td3XHQ2SDIwH86ZfMN7zI4woWspZd4NpZKDr
oi2vb4j3Rf6Z02jMXf6DN2+3zlm7rbARxQQI9BOb1CvfDNkZTCZa+g4qgk40aP9AZPqNANGOOiHf
QaE1THnvBaJuNawgz3gxR4KEG7OBWewjKccayJ6//rEEv4U+YfDaMl/eK28/OMYdbY/J12YrTXZN
b0OL6Xq6y/MZuoHYP2O2EZ6INtlFS+ynEvFcsty0X+gT6Zqu8vS8nhJ99T6muOCJl7QEHVsWyo/U
gwlpzFDH94jkjBBZg1lTZekeW3MunbyqXiwBdErv0U5kfhs5okysfFlbkFWI8jgVTz/nU+oBYwFk
OgZMSzXh/rzgJnJ2pD9qS6ABB//7h9U9FPWrlFAV2pEEDOGp2oFBpUXnYUbSsnMi791Ppqsn/jst
Ja9cTh9o4D/Jca3qaRiEQxZLbwaCpCq7GcqHOQpRtjWlmN3qUjtT3Dw8RgrTrXUxnpyhtfTHoQ21
hchC9aZu+4ZmGERh62L5hEAEdw6i1glefiUhzeyLLnbJuyM8JKy+Ht6vjOkx4kC/Ipwy4J4f4OXZ
RlgYcgBLmtzZxsJNpVByxOODuuJV/hce1tR75ePLStym3YE0kYV/p48m5kP7P8efFtFFgQJ3VAOK
UV9YXQmW5ASKZrrpzUPgwig1BlRYKhJGb4A+A+xwffpGZHM/l8KwOOzQbS9VM4WMu6k8Mz+6Fhya
gU78Zy4a6cEn8hkWGnd/m4UPUcuTsWHM1Y6jp+oeiGFGOBi2Ivyst+a2KO9zMuuvwLkTE/xQLSUj
HId/DhR4B/hjLuSqb7idFKHZxYKLbpfLKDMrfN+H93j07MVxa26iO2qZLUpxBBTpb0WnzS3zkbhI
xGC7/e3JYGPSBSlBBZ2dfuuQrnk2qrj9eH8xozqNZal+9QFj4jcx1OBEL7q3sQX8auzB9IMfwYXF
6MXaJDrrzw8AiF9bqdhZFXk5V2yTBsGd1aD/H/V3peVBQbv5oNccEqO+oVoUuNZNUhhQYprF68Qq
RdmJ8jiOpHZiXIS77O8qbPLIZKShbmnYz2R2GM3ZLnnjhDdl4n/JDM9cj3aU7OnSL+ukaoJCm9Hp
55ho5Kbcp/jYp8WldsqqREHROa6Kw5arHqtKZSRNEOE5mZCDJzbZYzUAg0U+e+3ch7ZSGu+EYktQ
nxCliV9xAiCgCCVl1XOkc2fUsVacigppl6suvY+Wljaf2Ji7t3fXqUd++/nl/zP8sY2D9/ez2zH5
0Rb2fYsylE1/g7E4QDT7/pIJfLrzD0EhdGhk0DjQ8g9DSwn2qeBO/DpEWgq05IjXX9i6YtWJi13d
g52ACAN34RgZnmYYZGoQWKg2nGDQQSPqqae90Bc+Xnh+pZZ9KOB/Roh45Vf6AUPIP18cnLnTRt7s
rbcrI+SqBq6xZpajMPFOZ18n9Z4AiZMufKW+g0o643Tw4CsLYfVIbwSGs5axA/L040iL5Sn78Km5
Aqg+jqfLGyaIncLWHHKziMnIyQ0vOOq4WHdjvVA/FrUOnEW9Lf8JheFAd4LXCyIN9RTS0pOWxteZ
PqkKec4Zd/ulOLnboIp+TVF1kwYo/gLJAMGD5WOm9t0wCIq+rVcFJ8IaLhZAS4Aw5evJZfrIwlcV
0H6ZwbpRRRjmvqiF2Yog9pqtoUAE1gAtBWBNCMSXZsPAP0FfRqqbQPmgMjbSHK+ACl9Lzcn72RxT
URCSBcmNGkFhbVkzWr3Z8hLgA9lfMopYC4AEatEIaXBa9/UpaTgfUOJkPVBs05WQPwBEH5CRV5TM
9vkfcdi9V0EjvDq692famLQhLhGyqKr+1h3eFp0qW9YRWYaqg/uZA98br0Kkfr3xN6HPOlay8A0/
Usk145xTLQNp0j+bzlEox+55IavfNDRUmVb8X9LgpG9+RZKij7e+slQwGN0i7ZySHJ4r8jqe5HuX
gjIlv1tr6pTq75Y5e6M6u4qs5kMwtKQ1wKBWi/w6SprnTvF/os8xaWYumBnw4ko3soc1hFhe/O6m
UqR/RiE1O6tyZg4kxVg6g7O/MbsODsfq+2FJzkSZ8Mm1K7TfAAdnV9V6B4rjfqlTjHDeqO75XHwg
1Z6Ha4Ed6Vx5fHcgqROTpSNdjZ/Dc8IOGLVizUcmfaztqO74or27ufP5yQZng1aoEXU+8RrHiT0N
JbsluXzVbn982nXior1tJo+QUoOj66v1SPE1zdwrsoqajXtumrmV5qfU8aZyiAV/4/0RA4XnbTtc
NIy9fFRsSUKHCzDA1f8m4LlAosVhdE1TruPIXzym0A8QZJ8iVvNrL1/+afwUWe0Ox9PMCQ+QjqXP
vSnZupVysMPvoMP+Tduo9nzn2hdzKNnnKqFxCgvCVoY1cbZd8fe496bNiguTz3yf8DNOASaARm4M
ceUCJ7/1cHf6rkcLnhZQwA78bgOqDarn9m/eq/+5AJYOoXPZ3j4dkea20rLo24J3AekYplvKeoMr
qmZX4MqQlc/UrN9SfopLJXkQLYfAkfbN8VGrNBUqLIYHYmm4BSK3Y1Ta/zPzQnZoHoxeCoJfHp+j
zVU5dAQt2AQyug1ETQwWGcqMJ7ozUO96CL9JzmvNKQODKl7ezc7ByfqPU2YP507r9jWVDmS+bTD1
7LsteOmDYjHg3FgsDlvau+THcq0fz2361HO0lhcPzbg/UvTWbeAcDXn9c8UqgUq6Vuac5bI7BGE+
qO80zP6vUiq2lGRyDIm2CyZRoJEDPPaBbJlCSYS2y6Rjg8S46J01xB9vIoCZ3CTOczyCtEYPrdzg
YBZNU0yHL14ElmKgvux+WUkXCfRD+2YPEYvWoK8av8/tq8H2g0idYlh/kCh6hVvSiSgWhxuZjNwk
kTiVYJpmzoSaklDMcNDaRNT8cFMboCn1R8y0gka4RdeeICfUmE9+dMRL/2Dy1LrpijW0OWAqW9Ye
K99/ctISzAQj8dajE1lPvDfSUeo3NNfDl0LJt7gjXTbAFf2l5eDQ6YnijRFApVImH7gZk5lauHu5
3hAukW/d6wEMTMzjjLGg4PV67QmVeSsNkNRnw0/PqnDyUlxt/Xmc4VIVfmdehp6+/MHYUWcenfqX
K2cI8QTftK115vA/Ns/hQkOou0pZHqOqbdpXHhF8PIy2bJyBVUNAf4FA0g4LCi6R+Eaa/9pGrqJJ
qUv58kv7ACGD1LkuUJ34gGG2fd7Xj/CQA3ArQHcau3hx10PcWFgXkQJ8SCDDIOCeCul8A1f8z4Qo
On8B8GlgdOfkcbjpN8zgj+7lGjNzRmxaK1KtzJbf/Js59A1nfNuZeM1/3/aHPM7XHxSoOZZX+YuF
MQJfIl43mIHXfM2Flt0fNRsA/M1+Uv6jFRG9k1Psp9W2j+OdamlxHFBrWRgm7mFAO8MZ7uk4Fl+i
qEuc0aP7xYbgsevnp3BrdKXmru9LAqJmfCPpeNd8bPKqWa3wGgKFCfq2yeub8Qqh8+utZ2CRYsgx
o6tCe69iFhSSAbCccI8h5d/CUnEh2GFO8fprQqbJbtbLxRCR+CZ2m/5l4t5mwqlkj/0PCDqCkkXy
4mA/stmb7cpqbvOBae9M/PgHmLSo2jpqmKn4fLyZi+Zc5OK0rRXdvIaTgDlZkEKgCRgSaWAENS1z
XqOSQl+gEOVuGv+H3bxYKLXvr2N7+dgKaWycQSYBV+sZh8qcigtjBB0Y98xJPfb6zLc8OcEXxp95
dJu4Fnsy8IglCxsbksW6QW6Wja6qhQpZ0Yu7yH1wuPo600lAUeHiFjo0NHwXUge90IklcN6zIrvl
8wYVG0sw4cNrZ2nv5qxG3mS/LNSRt5VFIgnVB93cQOvwWNbtoo+rSl/IliNLrkIFiqWqczatE2xu
JC30ADj5vOGiBeFjszwtAr7t06BBaO+j0I0PcqqsaCZj/4MWChHWX2iZ1xN0KXsPA79qZ4fNC7Jy
CaSjRePvSpFojDDoSzL49bqqW/FJinSbWdwiolx20JaaQGU4iPBVSy1UqJgZcThkbNcnbcwJS3Vj
9hD+JdHBv+7MNbHb+ikLSah7Ids7R17i0x5k/tDigmiwJuafUVvDfXmAZ5bxrBwWN4eV3jYbv72O
eTZa7ytWjfsVCc/vmjS4wr3jF0lC4gxQTtUb5h62J7oG5Fh+8qXIkVzjvUdhivyxI5YXHzv5x5l6
G/5ws5VrAwqPGA5p6SFYoA70ph2PgBHgFcUSu09JqyTmO62Ioq2C04DmvQ4TeGIRKu0LITQ93fQs
qNfgx9Q+hw4OU9x+Cgfs35057PsjHK9emEtWXt+HFzFl2S6HVX1xf1T4+9UVJkaXRxPfcHiK/bWM
r8JLrG1Cl4GZoToPUJIMllTnY496utJ9K0zIJeaR+06WLnqVlgFAXIxPCsCaZjurYWD2ujPuUqcQ
BPWzSYvkdkwY9JSsZcCDK8kdHQxVCzvBv+A7Tyx3fmxN2Sa864T7gBqV7kaitYzf8UF+oy9CfPN9
De6NJ8kca4gTiq4Z6me2fGpVPrR2alPeExdk44J7p7NBgRdgevEculL17wogrxWIDOyt+CENiKJS
ifRq5lCJqVbIrPka5WKLAtoqmBhFGpMER0IMI/oLDf+k4cZSwvmxDCnXkKuAXAkcALZmduliTGz5
L3CD+4uCtU4kwBV7+vJ64gsKDll3mNOOwC2wRj9UwBg7pftjrMTkbcikpiP4lzwRg7vjDJeNtt2q
Dpw2dwTDr66DmE4mPTjx7sYSpsN+hIEGEYwbxD0QG+yOOezrIORaKGZgDULbc7TGz7NBeStnU2yV
klwk78H9K42iF0Hx0Z3xpkeSQS0xZ9WlbspMJgZg2IsOSOQDGARbIU0G8qNf2qMHQ4d+6L/kLlKg
14DNbgiGu4RImY7/+K2mcND/AtjdlB0rTtKmO0mAgQY6JEiwd8+ljMEY+wpiamsXzMLeXGG7qWhf
1EDxwk+O6fhcbcS1Sp5Rpn3+3ok1waR25n72IK/r5ZuA8unYyde7+vhgU32Xn4N50dMR/ljZQ6y5
Bd1FTeUaoCuAGR0PNrElLcTDAvEcDEWksAUfKiuZ5tqwI99EXQRqkSG818xm10YwzJJmnIxHlpaa
TWI7Sq6QNfCt0ujqJ3Y7uo9vcMgelHJ86X3SmBGRvhZiwEgCmq6uDx8n1ame84GmP4zCIqnsrd4B
CCgJ0f23ikgwUVvj3cLjX/5NurS4dmGNk2ba+Ilr3VlFQ4ovaldr17F0lwCAA7EEucQKdKkIflKk
YjNOOGlK4qKfWD8luzZ62YzmJaptbR7hEOsw9W/c7Pfp7klVpUYbhsEeSSK+VnXrK9H77Czqz/g4
LLfRMdGdETVupyA7ko9VRak383tU9t7rOGHTo4XyPzmECtQOTTKS1qo+PXS0yAVyUIR0mn3K+aPq
UK1o1l5s5MSFssuQxiBos8syOoKlbRquSJMGaN93pomWS34OTxL7rf1N2DakOIkYPZJ1+vlmC7GI
4GomH6S6zE8RcdM5SeCDUpd4Dv6c9C0wS8ULPxb+fMWsKZnhwga9PfwqYztRvN3OzlFHdexspgOO
oSvHNDCQqagPkQp4ewVAa+yEUgBWvgt5/zeiMYa8nFLw3hxyBW0DZd6N+/FzP9Gr7FmREQaN36zo
J9xiqc/WywhWJPLcsnEdhcXspyCsmcCsxTDZS5Rlzy1+/FNMhRP49+tadCxW47vnqcuIYA26Eccz
ZIjGJdWs7uFcsb+S7BGL9Dkvxi6kgk2ikNeS5g9fgl4AptwIBvn+5zZVI6X3dB0PF3G32y/m7I3b
KVnWxVZey3zoH0BKMSitvTHy4ENe7lblRK9jXSaPMYlMY94WL6GSmlg55LIegACkbsKj1qGF4uVs
lxRbJDrtv9VOChyYQRKREoSnNxTficvMZJHHzFLE4HXZ389dsvw9juxQP92uAuLLzJ+ft2Ja3p6U
+jI5afhuH6BZn6zBgXnkfEcgTDih8t0bugK99k6hor5AC390yCko8KN0a1OZS1AIDibwS93pq9yt
P1ZuHYtyG4hQ73cM8JdDj/xKBPEoWOwPkYbizV6YPy1H0SveYi5qykvkYbtSzGtuWcY+bdPrXGsa
Ue+Hs0zIiUiaD45gdy2EW8j6IysNvu/N68tmn0su3isdf47+hfYQs1aT53UixAmgYtNvj5cIYM8y
nIYgJnB2gZH2VBCNzrQQtF0z0CiKY5NfTFUUSKCrpYjeeveJtK6RTg+IaFfQgYmzv8fvSueUEJGm
aPF3hGn2c12FE+n9MStjr7eD2RNawzZMgnZRrS5LJxapfq27+DSrB85sd0HafpxtPKLAOIeRBAEC
e0BuQEKU29UhPIOuUCmtYIEfKajiNvku2jvQhhR1H5hSoppaan3F2j+pqsVbfVGwMrdvg5X+72i5
DvKL1kBjrPBqn86Ldh5YreucdohY3B/JRM4EII/9lh1dJI4VezkUFknTlQo1orGR9Ta3IOwfUBH0
PvsrBC/2SO6EF0EgUmkIT/35my8AGxEOuaDoqvjeulzZmHZIsUZCd2UB+Hq17T44OuTVz7n1dyXE
UHfiLGguHICLTfTCEjBcS16KUw+f/ZsiM0thpGdUXNZr3TXh/FnYSMiSWWOdImeKyT+S6yE1d7KB
Jixt3ly60qBba7znM5CpSd60Fwx9BXmUpqsedITYs4m/I2Ac59WgIc8pQy3Jrcetj6t36UZEztcX
bMLDt5r/12Zc7FT++LkFQx+fAZUo/IVT7QfKtTu7TRG7E0U0fJXsaSDSlLUIi5SnrSZxVltlD9ag
eDkpDAIOq/13QQBDxH+K25yYDHJ9+ztTibyBe4+R0iwzWYoDoThdaJ9zfmYM+8OqxT8BuhPayxOw
8DUaZruGY0uR21qbDN0gHj6hJH6fXj7AtYxUjBhxsjxHxmecKyZORLoHismd+sZHwlbHXitViQdj
uCUucyTW5i97aOi3nywKxTskBeQAkdM8aUmYYmkFsFVh03zadoFynGJqRx6sfIU6uQUNjjlfIyVx
TALywbuV8cPL7lFpZgUNduCf6AS8RYAWP0/bbBF0ZRc1lvBZQTKbwgjkdGVaQbYm1TcddcY1YQiZ
UG/P9/O/Ls/PlzymUTagMi3u8g7qUCJySg/O0qy0bFYcUczMze0JIZMdZszLCFItTvrESh3e4E4E
wEmK1zKFycItmxhMsb4ZgHK9d5ewadS5KjERm4dnKbiuv0GdPmGENP9IQ7qnWpmkB7b/mAs81ucW
OHcOVD6ke1MObTSid7s1h9dcU7r2X23ZnkA/TyMr8ZxDr00oSnRXyGaHV88uigCiVYD6iJ7dyIpS
apwflvn0eFl576mK2mEfyimawk9CuCuhU/cqFo0xM4RK/AIs2SQDqjJ84OSXFRh34i/iowTST9Lc
d8e2J6Ox0CmRXkDR6TfTs2jMsEglGIR8WY0ePX8Q8SKlFjgS101fSMTQZS1LelPHJp/yZp1kT/cm
mOYUE/+bo3Nuz5aa5AgIGUJG0IkDDpInk4tGl7VJ3kgAN6LfGSh7ZD83bXcqX3YAQufNvvA9+9up
TEwEbE6hqAWeLFjBH22gTbF1I4fSwWmEPQM0gwZOwP+yWqpDtxKsZsB3HCwZvitVAt93BHwh6oLL
em35T3TG9ElzpCDgfJcFGLse3Y1ViHA5RtcTa+uzV4AE8IBXHcgxTMJwVHNwTCPVX5v8stGknbSV
EnwFNw7WS6Yege8Q3HYxDhXWOc3CDovDsKjSMQEJ9K54sriqNYHOWAcVDF3uqPHG28FGu/4iQhdk
lZuAOxeOffhWg4Dv5hdRWCqAmnjsZTyvKInmOeq+wXMGUGaJkHCouZ3FUBzcFzVmmFNoUFsFhHV7
1gzOn8NGBer0pBrUqTbsg4leQjLWmRqYTXZhmX3j6NRS+JkupUwnWS/a0rXYx9YlfMnrfEvD5ECk
X47xhsHhFKRoq1thg9qpkp8+CZuGZxofYTJhIrsPqi73OYM8/K25or3R2W2epXxj6ognCL/enuci
LvDVU9M1WIkTTZPohVrRivr0LCTsazixm9f0LB/gzXU9Yo6hf5rbBfE+qoLDe6yAt9l4m/R+U/0A
tvOTG1H7l+eW7kPl82JsoULDXeyKyaGbNd/zlFZfXQ51+0aHVk6rQtBLGjRngf2rke7iZ2Mkvfgp
F3p8jr4p30pZISAk6wLkHoSltn7EXKCT6Ju5EBgtAJsERIBgQgyGFnjLsd8B8vfSxXdC50oaSU6x
y8PXvFlU/LDMRcQ9UW8ryc5sKhlY/67veSfPpLTH/SLt5BcyDYkYCuDuT3vP2gTD/x/o9KS0a53M
yM07SQilrAAO9ZFpScMPZJU4A6vaAGs3a1TZHGeXDioNGoFT/HpG6oVaVB6zKm357W5rCcaZ1vxq
n11X0S6WxQ0+p7nriSNVRwj0pVEuOgDgzq7msCy2fSEEfRLQv/8LYtI7ZpmU8bSmTmCWC4uli841
meyFebXyvPU/FhN0SCR9yh3klvqe6APyh4lyOG28yBi4/v+FSOHoDVCnR5+gA97LQG+G6uCSL0JL
NQFhbk8Gb+qqg54PUHaEHy7g0rVy4GQySqcZhpKEwLI5Sh6oclByv7whS8TOoQ9CIYzPBTh2qKHl
3p61p51CvB43fyKmpH6SHLx5mxBCIMDZrRBQIDBql7HHlpWS7LzZPwPWTBYOGk3lGwlxne3EVr+T
XmUshocLWHnUTCMmPKcDMs66IHgU3oDb4p8HvzeDljULH2yl0AWz+0unt6OFChQwPOhF4+ILQF/N
NIecAiCkLXkkkbKqZSSjjOUcTszOzA61NIQo4Gu7e3llZKiH7CUtK8xddVTKhXvP3o+yTnZ5Ys3/
h80ljfkiqkf+XVCXEus0zyPnKfqlcmxLDShURdSqOZCZ2pZD6Ll2RMkZFdhZ3bEt6mw1ReHAb7Lb
g6lcnoJgrwPRCAXbp3wy0QDqvCWfGCgwyf/I0a7tZK/DrO3Q5MUxL+yzvE7uTLYaYa/QUcEmIbkQ
vMBW/UHWWz9kkS5rM3O35iba/U5QgqyppzBiTplK4igEYYSgdEQl5xK8dX223pPEj9OOLsRj0lvy
1mB6R83QxN1IZriEwd4ENCu3LZn/l8oXgHutjK9gN2twMdWDJniBpvZuk9aJ5vTq5zr2ZuDrx3sV
EmqtMd1cn1M8N2PKCwuuTTaEG2MWC94OzIHgTNWfw6+0/GLyNiHZZ6OI6HjZyyrX3vHRyX0qIAmu
LpnnvJpMbOr86you3fJb1yAajLrHGYGn6KowK+Lyu/YdKrSANJpN6/oJDAIvtMpdZAWWh9A9FeK5
vEn3FCUYaxFyCojCxsNElj9xtR2NkmL2+cYBTV8d1p/aqwUHTxq2ajMbWUM2URtodMhM7z20maob
qSI8j8sUuRdcokZzOy0oGhxgQn/jHP7M9koxFH/kGxmQ11VaPqlh1f+IDDWY/CfG5uP5lzTbi4CL
zaFbrt2/kPWcWPAQ7LF6PjNSf+HPqHzNg6gRCCSCSABG5r9mYG+63IGRBmbm/77J3ruYSzwtbe77
tRF57LFprc8cuQK2LHB8mVEiJY2utBSmN5X0cnYu9JDvGl2Q3XNyvErUK6twUwUm19TEwFOS2VCK
OuJDiwkXVRmMixQ90QeI2w/0KjZ5/Q46sfEFAvHo/ZnES8z6xQyCRH/01PZJ6TfJ50zniTfvVTaw
+bepeDFs2nO/k5HdfjaAlzrZRlby19cQ4ezjxCRTIyJY+AM55VFXMWn4+LUUB9DqrNS9NHouansZ
8d6zVsDMOzLl15cvLIkXPDyr8A8SeTKw/dp5tI+Ehh6TEAdJYKfmeHw80xE6NQBe0E5E28kXlZRc
Y0uJvK1fq7Xbgg5fM+pjdt9yI+SVRhF9HjsaXMrJ7SGICrPFhBTQ0lGOLVTBTqLZphFxPvJDIEBa
bBk0TzA630pKJwz5JcLTILPj2hWYTB+dZyo6DzDTZ+FFCyENvyQFMPQJ9fRQy/S76zr9LfCQRzN6
5A1/OhzXK/VtQN0/mfdeK5lWJEFkvPVLI9UlgXfS3zD3QNQqrumytcsuB/ZbJ5qRj3A1N552GInh
3KEsca5/8dmfU9PKKD7AUNoqIh62iSLm0GunXcVUdaRIYPQN1qX4cAQWZ/E24X2a7TIj2us4Z66f
boLMH/jt+1O2vORt80vuwC7ccwyHDkMcDwdwhj0juzKS+o0qbiC46daa4Fbi/5O8YPuM31CbJ/aD
+f7kE3x92wg7Xf1JB4BsIR10Kyi+jDB5SSGZC9qRFUh8nYhPggEOXbF/RGZrz2pVIVlsVXuVJbMW
a4pQuFePoyPNFgu9k4evevGVknh9BFwUUt1hxMVvvZh3rU6IO5hCGFz1aWcsWbRprKrhhn/a5twJ
NE1FChfK8GsGT5R2DFuL5F4xW8xyBsQoTs1S4fc3qqEnP7sLJXpJFyHafd1fGa+KARaix4IzSB4T
TBjJHe+RuBtPAfM7H1jTYfRo8C65cJjVybWbopoRJ41I7FIyvKyZSo6PiVjsJxG9k0viI37Oc1rc
RQQho7iEzwRzvjX8OgAyRo2RbMAXGc3Kgnj3jRlcME3oHw3vYwiH19kT8I+gg6wPsihPSa6+viTe
PpQ16kxnAKI9eArhgpNa5B7KFodORvrTt+dJOZytMjexv3D7B8TlerVO7A+crOeadUjpzmSVh07x
QfXV3yc4M8JEB/XJnzAHVgUAeb/CSRZnlVNlWx9582x4/fZ4Ewyman6dhXT9Z3MaxKAQuZde0/e/
i0VXfWfsVlWF52bEtzGCYMz5Cv58WOfTaMWXM5IFKlxN0h5PjhmC8x+JM8NQzF5XgqV2/EbBNf1k
WwbEx1rK6BrlfT5V/5z/s5N7FVrXcN9Y8BlszrpCLfMH/MlH2H2j8AeCj85HbRd6pbdD4fQRjYv6
8pXCoDolx+DesdZcb+B6tvBj0tASTVEG674KIVMh8RPVBZdfoZCSF90NIZD09ip2+jtvpjrqz3ai
NVUK++QfYItjA5FeCzY1GNdyYfwJsF6aNwewtkN8v3VDgMPZmsFpBU1bWGNJE62vTOlUWBnjBhSX
KDoaaJJO0jTy8XA/qIwu1hpWGeQFYjM7qK4xwGMKMbRcv/rjPg00jGWgy8wa9mWVh1LyqoSmQ5FF
mAA5UCBqxyUGkgbpmpZAi1GwIg1cVOKikbYCv5NkuoykNqqyf0szo7w+iNizN1c6g+daLX0Sz19y
Nk6oKpHUVFboPQm68oPY52Aulpe/XCyOFxyKtzO16AQ45quZIb3X9g+A65DvV1uO+w8WdUuQUJJf
u3meOgVb64gL/6GRbjBrshCmoYBOKpSFfP2WU3Q1biaN+Qtced3foWttFLMbYYWjr+NeUgNt4fgc
QO2+mk1ybmPZql81lONgNkOTJ+bYc3JyfAPredvWJV4P//t75ERCup5AU3fOxbnCXsct9BqnFckJ
Bz6PNUf3+q20jjZSUlj4mQKubMPL7rwNecbHnYSZbA38BhwKPEaTH9ecfwSYrYvFUc+pwDheH17S
/hIxBap7t50RE9dTLKb6y8wyGRMq95VADS0I3XmUFOAoc8WtwrLV2dcPKu/bLlpJPAB4pmmCObk/
JgOsGnxOcrpukF6lpdgUpw9IVSUBTtyWbGYAtPtZG98rvYJ10Uyed8tOXKGcfrOHtUA7nds5JNp7
HVHhkF6A9avjPo05lVjs2Oonov/JhtTMZ0kuArac1vnXbQwwkKNDiSY0WDYo8FXNOTXs+tCC2uhb
SyYave80IKo8SLqBfK77vzMkcKRYFirfhThyhy7KYIU45enDdQuxxc4N/CytbAXTxxV6hFj7IixE
3LtRGdP9rsjBLLD+Nf8wZrRITjVKZcbK7IViYW0bciaUtPutzzoXYv9dSUn7hTTM8Y0DMJAPfCBI
Hpli/jG1pY+lMH8p2RlfLK5efrxQOZh5iSTIIt0NvpFXvDGM35ZMyr2idwQSSlPE0uUdG4dXqkC2
Cp6dRWot5U2UTn4kUlMXmggkSLoWiumeOc+1Wlw3qULjRdtj7fnl7nOkOduRNY+WUQJUp1DAL7gL
h7mpN6Mcn0sBjpKm2zDAhZNDqoS6kTKknFTpjPgucb6uqYA+J3KZ7gYxn7JM1tcdqLzM6gWCudBs
i/y/YZJunzRFXsLL4DQmiVBuz9YqDE0WpyVFLqszjPX5dPuNjs24p3gHLovPG0DEnilig4MTHBGp
sx3nuHRUL/YnB0eRW3KNlTmiNgQ5aP9WJa9N/W5l4i2i24luopvWC0PD/l2fj5PRzHOtyh9XL4HD
XokBeekJa2txKHQsvMxa4YCMV8xHX33YZDdz4jd7uW8h2/SekXXWBjeaTBPpyGCohi4dShY6+C9c
kakOh9ConqVZMsTA7ZDxA6vePgs/+ucWo6uZlDGydJVg12thlf5YxfU9q9/1PqSoL3SCclIqd6uH
qagX1zTzrNJOrmWm/MeWejCFr6m9CCpAS6qW4SLytGvtWz6MwhLiy3NuwU7BryWzf2TamSiiYXkS
rAYuQ/6RSAarqAfqkkwg0dGagqbSpPL8YrVd9L8w1E/AWFzrcPRWWls0H8kG3em6AgBk/3m+0Tnn
kLmS7A8e14i00W8K1LrI+rdTUHx8oZE4zfoQ92bZeYz61DDtBGHAcn1DAx6ewpOYrg5Vb/Wnu7zy
qx57gHu8Q+p+ltAZJb3d8/6Xe1PENrZ/gE0v2yilif1G48f5zUW0D8Fh4HdrGn+12ftTN9hyI753
6sHByNaiFlbnTHy4N7qKOow+bX7YIMHkVLZrOvm+kyuOsc9AWqoQRYFAMfH6QTEBcYy4rr3JNTC3
ZZFFnPzCQLH2WjT3JOzsP9gYFdsfL9eIcZajMVlJinI1vgwQUtzpKc6RRDAKjfrRTnPDrkBph1/M
Dxsls1vr+6onETYxE/OHpd3xFESLnYO85+YGz27IPikgre/T7CDqcKGaCOOfa4knnoYJyzCznjLj
0jAjWZAxJkgxhSb+PoSxeA3e3JlblSJ9OA3OgcabfdO2WW4r+Vp0tmOFCrhgquSOFfNeyBUdBprx
CKw4BuDqZd6RNAxFWOkeDJdks4xC4WVPIlbSxZJjogudoJleBX6JYwj1wO3cFYHxaKbOeVJuJLqc
R1wW31o5WQgUH5uOEAOCyeKFxI8wRDnUq4C3mAVAt0tgt9R2FEJzG6MicoqT0f9gqZn+fNaDxC2b
AYZn6h9XpS0dGcU03/fYFL69mVpaZ/OoaQBlZU0slI4SrNI+j+TNg6WOtx9xXSO0OxxgdnF4kzvx
MOHLPj5A8/sMnus3SeVRrUw6NeisMvf2Nqlxp2glV6z5JP+cD3QgLbNj1c051bC70CWkXuDvnWfJ
WZXvdzDxhtvayEex6TagHnvUX+vVN00KhXzE4b1KnK1y7W8qYAC5AFpT3JlViD1Z6p7//jRU6VKa
rBPGKDBopy04nWZRHOZfEF8UNGOks51pXa1dULhkFOiAcnyvREo/efCZ9CDgWweG5TbbVa6Lnham
gTD+16A799a5QThvBVlWHWd0kIHdrXfAaYc3+z1SO0MWlqLsXVV9R+7aicoOf5w47iiv0Q4Z/XvL
vsZJn1tLOak0I154avqRrk3ud1benkrzY82z94dXylcyYlwXou3wrgwZABFaoKoYEolJnrrU0J3K
of19gYrZjrkIj3+d8SQcxfTqIFn7FCPVeqUgGY4FOw5iBqk5wEvFFO2zFbSq/g4zMNo+kW+eNBrS
3dAQivtw2RpK1v0sAac5W2hVbfF5QfN5l5y7giE1foPsh+7rt+M9d8qQTpVFW8xeKCdVJQDW2B9B
N0DXFKlAxWpq0W2vPQH7pxJl3yP9gsqQCNQKnuXfVIC+ymzm7Vgu2N7Xb4UDSfFA19Drt60sLUEa
Seyb4gZCuQq1f6VzeKohkmCsITRaAYCtmOgUmVWBcOGxBvzWZxX516PiGdik4by/XBcd/qojRjK+
4W3qJDDnwMDidQmNVUjt4SYKwx1CrCtIdJye85B0GhuM83Bj0+dFQExS/kNTk0ju/iMjHyi3lGQR
Qeg7zeXai15pFh4BMvPUoHuOYoGok2DiUCqFvQ3hCe5IRqshgs/RCpRnYvgCdt8fI21NHVHnyL1E
l2ZDE/Ota/qm0cfL3Y60bQGlS89ZpXuZxucBuhnac9SXsejbXDGeo42ALK32m2E4ounvPmFJ2uV/
7Pk0aNthv3Z4/6FjZCPI3fnEG1XqVfOykqjaV2RF5nuNe9nr4HhPAOKqJ7ycWiv1f2buFEOrNsz4
f3NB56CyQokwxtoq2+UI9b81Z4Sh1uv5wfa4H+LosHa9PPq5mw3kBmKw64IsNYX9Si+0eJYa9kp0
iirIGyPEXIviUhxTWEooBTpnpsOuRNrhKFBjINRdiOXstHhugNK4XJTNWRS8qWrzhPdw2r8oIb06
zS8UET8F2+vMu9EXFqSMByYsPqX6+Q77KpxnhToQiiKwJl80woAvnqL54PioQtPcU5NkofgWF/WI
EoTZmmVpP+1aRTCQtkQ8yylhNr7eOVuy5MFAC59kvNeKx1CeHd8BHuCkFN3DDrcQRZa/+W2EnCJg
h6F2LBbp9BQ/XPL2356XPgBpdMXuRWUerpsFcjcPLYOBwl34YvjNdOquyG7ELFCwG7q2bjOWhLAA
WM8FrbTgPOEFrlu1l3J6ru6AiUCPPMErICdbjLAR5nfb8o/Q/+0NsCgmvjvNj1drmorxHuBtw5G9
pWnl/587Z1H1FcafkHD/XrKm5RwQp6uaJIE49Rq4J/ptyBEWQ1XxqZuSE+TZrfz3FVC674FyRm+y
vAmOTcnDu68TyGw05BGRb9IRS7pQCtImYqq2jQwzwul/eG8bCASqar4CIEtT1noVCTTJ6cCWsbH/
lJT16M/UD0aUCJZCrT3gsVKJDBLRevUTvMYa9KEK6Hm/MOJTLV4b8LIYm+u29ZYsLbK6e3usNli2
Hop2bkoWdBfONgvTeST3PQO2JgezeRSKtNPlRRZ/gthSOzgAk6p8rUcI09pS0xUSLw8oF+MwRpqV
8Cg5upNzC253Vfxe1sYWmpSY2gJmKfK0xVhAW8OwsvjR6hLmqk/NT+6XNx+HKMIEgV8yjM2JvuHy
KgAxvnUwTLfBYKxyda9mES1mwxwtyGbAVEYQ2j8Ui+eCFCWqSiF9EOpjlcbOphvlms3cwEzUYFQV
/vAjnzEYdH7RjQQ4GF7bC1H5dI+GJsF8gFea4/TW4yiYHA30d97ZPnynFAmYetCwYQYShR5XCrZJ
pcPJk2Ajkukli5Fl7UihtlWjptQ2/xB7CSm7Y1/iZ1O1S2T6QjTI/PfhZNbQ827tVnxmbHhqsGdw
7wzwAEP2hqKbTn8FKn6EgX2LWga79BTJ+6jzYuXH/6dwhUtn0K6IJkFrqrupnnZL0Gx27o7m0xOo
znH0Q8vaGp5ZiVJSHZAU5c7j67LYLmSwrAK4PPNV5d/hb7UW6V2c29oKb62NTS8Am4k0CUnW8elC
K+BNh5OTkVtmNsPCAdABBf78R2Py8HT4lvDCclU1JIBxS3zx5pQ1LBIrkP7d/Ce9PpulTey32RJ9
aDFzbgnKSU9PNa5WKXcfv8fm7TDCaHbWPIXi1knGpLpf7aACWvsY2h5eVpU2fs2M6vkHoh8531w4
HiME2OWRyM1SMBOykKWYLtbxVSmcquhv5Hut5ayN2wsWMCA8lvstJQRWDSOVMCKhNDVONxnODuEy
fLWoEClV6D24a0QttNBjPpdBVSypayvR/Dht/asBI1kqMAkyAR6bRImbtRZcYSTMCNYsDHuBpQR7
gUIwSElpeqpXaSqZQD3n/V+uRn6WWweEx8TrdSMZwTTjhLx+vY8oH1vI4DTfxivexcwD+zxF0xFL
AdB44rDye/nzwbOnC7RZuyUz/hVblPBda2cEeQyjGUb5jnIgl0IkNExVwO8IoEbhfwFkFmg1DcKy
0/0FnLe/n6RBm4bO+okXTIMVHeI5rlEQr6Q1v6A3Xx3auXlWYdUfN6OPO++sm2fajXy9NVI4E3yc
5vvPAr8pNstCGtOF/hriOwgM/f6yrIfHoe6Sjg5K/tjX75dGLmOXKxpys76A2Pu/SbmuAoqDROi5
ou8MFIBJBpKhpSx4wKMyOAOPde1DZliIzlVMDh/bGSn6bZ/um2xvL2azoycq7izhWy2ERKDrJvlb
jP2TCXc/H1CqL0iqFTMIPA0B0au3IcQk0vuWF3WoLobQkD04uAioGmv5lRksfv6enPmGT+4zRXa0
SFC3EgNuvAOVNuDWfzYh0OT73Zu1PUheOGOEkZzzUL90dERdi6Nz18DNtr3IxFyjX3gAAtYKmrNr
Os0Rs+GU9rew58+vzY7N2vKFlECGt7q9ZkuFa180SXjR9Y/mKQ+chP+D8exgpBJRS5wU50Z4dRI3
F43ZZNauYUryDIZbRee5jjTJAiIbIxzjQuVhO7T1OZQOTfSr1ma/+WLMmeZKWn2BMktl+g7F4HmY
TSUpgkhmcZgg3HOROWmRF5jRiajekA/Go9JktlAiaoQtgBOx4yK6VQo1LpOOjlWXQH8cT9MgRwTx
RWfLfTdYIBMN5wL9qX0McQC4GYbXziAceECy40H0jMJlOAz5OcEuinYijvXN0wQ5gEi2O1hkJ5HK
dH9Dyc+huo9kmS49VkQTqT42zguTMrozLELTdcMwvyGkYu8lXNh+9AJzBcjhsIuhPzJ+Go30hXLJ
PlSrvQ27D03yxBqkyAUK046hP1p24QgJWytZzy9Gk9Ysc9aRpi6+bnEzczfG2JZB7vzCqYi5Lkrt
AhrxsRdMB/45UMq0oK5wOE7HKZDE+BIJJuKwizn/YHk16u7LDUwpqCoYx1X0RqCMAtJDPYYRAoMQ
5F2ndVvUqn2jCjmwIDTBowYXam5rC9W2xIxcsN7lLZ1fA/oQSfwKaU3lwR9mP4plFN1NrCBmHMb1
EpABH+tNItuGSdQ9FBtFVtE+wScsg0ipKh2rIQ7D6P5wOGaFsRm8CThMrBuLa4NPJL+DZev8x1h7
f++FvXs+7z9HrVLmWBsPY4wyX+yw3VFwSa+WEtC4EBcaGBXkuLulQnGUpQYxn1866trMaFPmmtgC
9qL1SaPkeW5QrhIoAfTvKWWIXLA+o0fcaQ0v43J0JWtcnaMg11My5KCceTiujSMJc3U6Uclv9KKL
qVtLLIwjSMy29keMIaz6VRSXMrT+lWbMkrnQWhyFz+H+u9nc0PwU7STTIiNW0yL4YmLjaxijeWIU
LpcYRi1FrDR4hVJAmvxfHZ0ItsoVX+SNQ4SI2aXfDaBl/1Fyk4Xl7wplkDzXFsL/giZNiVXyYvt7
PBTV4EtudRW5vdOTfRKnIh0ZuIHvHW7bzu5GjqISQBGyHv8B8h3/qE/Fl3sFC0/dlAMGDHHvas+L
7JQxddz4yeU0KS8N5ONevahWku7/HOom9xmLEQScYe2vGQg1ry2YB2NamWszwMkAdQsBD2VpS7YW
yAabCbx4pSP9ujKG/jmL5QlcdbfmBaoeT3dYfHCPG6wV49lzxFlFMos9s+FFFhG1hkpVmHfLZ6o1
3K8idCihJB1RKC+p7WD8E2HrHazZuEbH1Mab0H66iQV5rHYs9gJxITpLWBVzDWaQcZK8vHBzn9YR
i8tRM7f1+PthhfG4qBF88Atqx3NEFQtgIRSKtnTtYIy5Q8wrx0vw55gpNEMj3HPpL73XiqS58NI9
Vzh3FDWgkNFQOAO0tDnMIoD2eqZ8C/QSG5dmnr4L3IrQ9PQnzvH35ZCgrUpEqc2omII9YpbwRdqo
t5cc30gMM5bDB/JTKkKJNsYpQIYSLIg+b9KRRKRIJKYZnYUwv5nb6eU7O4eSypVZwzwUs3vrUmG3
ekewn5B3d4ckjK4I/DfV7Mfw+B8uDeIOvCNj84EqmiLZ/YjDLaNLSZ8yflRFqf06jE1scjHE9+Gh
h1PaPY/9jAYsOezSi3fMiIGkY8xqf3XzSFkoNIsdIUZgUNnws8X35Z3oxInTGl53Bci33z9msaZc
sO4jIIgq627vpwJtxmtkdmtKbLnWLpLdbgnHDPu+a7K1ucnmHJTM2sTdPs6cXU1U2UOgwbRW0xVl
ZO5tNCVEfMbBPobjWaA+qX2GOWsjdlwzacTjFlAGpe6hQbdLrFXNPWvt1IJjFtDnCKQOmY4SgTcY
et3hMrPT/YSb7mRN0mEpXDvn+Y/9JKs0UHbsmizE8bnkly2sbrkAuHmVshdPGW8Z5tujYbB7aLAp
BdIpanv4RPEYKhcTYiz8/Nw0OC+NAdthK3Ar1m359np1zeyX0yRumSrHTXjDcvVca1bFYbtF50SW
A3JMsMpQoHW/y89uEmRn3sK382U/x50EB06oOkvjPO2budmOaoZzvo/dY2aFHIyJd34c6BBVhujQ
+G9reYDKbv1KUQ9cQMTvX/WzsV75d431wDBee5tnxD86iYy79Kak+PJPUuQwOlBEtHyqVCJvm0Fn
4hBqG7TvRBXmOGMPUhPFBoBN+mtdDmOffp8gLL5vstiSdptjr28bPkqIli4f8/t54tYLn52yb4sW
LHhZWESYd6P+RZ8bVK0IMH9s0+sZyX12WCHD4mVfmcBfqKt8kkeLBCLuN+JKhbYCOrWScOpsa2Mz
lOEkv4ePidm0nu2YAV72PDmfWh2utyLNx/9wLIivUpJyxuyC8rdl8wKnKszSpKvRTEJ5fbfitFc9
e1aa56EK4KmojjwhxtJ687KWackmoftpcakGTQX7mhUnDqA0kMIlIYJ5nex+egEtZsGgVWtCaEEa
ddJjZlcCah+s4LKCkGsRBT84cXFteziFwQZiuZlJJqE+0oe3TOzFxJphkWOPrCu0H+YGnsiEefsF
r4B4Fz0r2sBh1bPHjwCBf6OnK00Sw6TP1T1tUcs07MZq9dt0BSaYkcjccqpkkBHTCiQOzD7XW1bB
gpa6ojxHppC+S+ZiJCIUSASmKf5Y9/7n2dKl7WBi9PXVQdDS278LipQ69Udj5pBtJoijuYFai9Wp
avL2JR8gW8dlf+RdVuxZGDuscqOHlJTHeqNUS5QhpmnJy1GUMWfBGuW1wPB6I07MaWLydQzQlE0Q
/iPtr3PibjJLHBJSyRnfDL4XoCyvEWhfRzTDcMFKkEkOx+tHAMlzsX8nj34asN+5Onusss6SJMPW
9lOwooZHkYlEsTp/RA6mOe4qZy7rXYZJibe7BbBL/FvK9AucoB6fAnhiEc69kffVnSBs4pE7cckR
1BHyW5EpQL7z+eYCJN+xNNCHDuZ9+28iwT83r/U0PYuqBExl5qK2Xa5W34QMvT71YmvH59KNKppr
VmMs7JEkxq/NRgMzzBrNRgLS48JqeMNHsf0Dj1jsGbRENC7cAU6opIbX3AsxKzFCHs0eWfxG0sxH
YWsulXitUQ8yj3nCb9BfW/6khQjDWxmZA0r2RsL656b2i+/kZviAOa9VRpWnXB2XhgjRceACCrY+
5ZinkxnSt+ymXjnjp4lLCSynZALzJOfimRQKxL0EAEveQ9DgpesdulVnXAcNz+KgzOlswNYkQ0FP
p4njLVyUH1Lqu+BCwPJtXVcdiBZG4zsyi7idnHCwmf7mJ81GTlv6lHyxcAeaC/pz9zrFrisdHXfr
8ZoEqmTnttIbq3WArslU/5tBuy8P1xfky86SZ3xeL9z+busgt2YpOigKvawqspe88P29AiPQSr23
OAJz3H58/PGwu2b6HY4HfhaC+y557BYnJj2Nw83n3TiIQzglYehbD0sTUwXUlZfim+vrSfl+xsin
b8eNhcDlJOImSq6MEgHa/tgRCiVYMdbnil/DfboMnr6qM5/Nw2j+RvKD9HYihT8mBCyCDOAlmASm
c6nNDdtlirz6LNiCm0IJ+gleowDfXIpbHc112n4k/SX/Bl0Q31gkMz0XcamsHpjoSzzOPFqEAc8G
qo56JVOO2Eq3UifmTbssFttt9FuwyZooVvrhZYeohohih30uZXlKVhLcqFV7N+DbfNEatRdAN/ib
YpRbCUMzWo2qWxdjMNx52QEFExLkfHccXoOOeksW6vNQPVPxOdCBMsCLHN9vCCx9lesgHpMxtfy/
eEen2BzBBw3OWebuW4FiguJ/fNxWm4YLNLjYYHWza4wJ4JIPxp31fuZjqupice+Yv9k8gmV2+P4d
5SjZx0xueIBCXpt1cP9nhWvWalgzRawFeZoZwEqdH6A1K052xf5PBw/V6GqR3+NEwdRbh+rF6E3o
jjTnK5vWfub8OUYLo9Ap7LEYTPHkoc+WbW3YZnW51Vi+AAmEZEDYGmGklAgaXtymqZrsjZ8BuM8M
D9v6MgryxQtzCgX0y0Nm+P+pq8WMDkmxJT8NWc3aBYoA/G6pwfsfFwzdrKtOLg9drGrG4gD64znD
2+VcBENee3o4JFc5OWNejFvFFBOuHKzRZ+mGGOEzdt6OyRpZvkyrNr7JzWare6k8N5n8Dae7Dhi/
6OjM1xs66vbhYXHDbctUaQ+shlav6oE3dh8Ft6QePhlvOdgbMKBSTUella6sU+QfOVxhWegd/cdx
AvR01HigqeSQ+E0u3Nrb1TsXSxdQzFkrWy/D/NRlqfE/yGmGjNPsrsIlgAKyP/WEZS1soXHkDYbd
c4yjMzg0FUWaEu7RZIZifzYeqqzAwrtWxWBN0C/RWH0P8POPKU09e0N1aeObWqnA5bkJ+xFKnSJP
RZJ18v4JDGCHQlN43MwgqHqo3Gzis/rUGG3kj8pcC+JRxVaxsNByFYl+P8zFKRQNd9A2nBlIl3z4
xMIlnc8TVEpL52nzi0JmAeT0Csr6CXcyJ63+vcWNewPvt49gYNiwHAQlfhoykg4bsEUT5luAyEp8
yUVlMb/JUjHrI0AzZmc735RtylhuvMxayRxKcM45VOl1SQbjKB2bECp0F/joOGGRDbFBL+jxcGlN
5LTMU2oFinJ/QSL/OV8f8SKkoYwutENZU2611267wT1daGQqbX3/ciu5zkkFU9wXBOK3e2mTMGFS
2j4cCW0PipzMADcxJe/aF2nSUt4oGid54vzDnJuJPnuDU2nzxUT04eJPm5SqT8watK/r62aHuCg0
sS8l4Qn82RPsjmFbGCOyy5o9rjB4AI4r8pob83EYOiMSLychzq+ke9PdHx7WciGpKdeScv56dBNY
uMGnH0AjBdjkbtbZCmIbrnaQ1lkHxiV3BcMbiyuDyEGlSXCP14lN2808RZhhk3fmORjfXnqF5jSW
GSnMs8wBP5kGCD/iP6RhuzI4fFx3CVpCWMVd1zgo14W3g8O9dg/XoChjEgaBbeQAgQuH8lLuw4eH
x8XTDQDHtYOvprcUxZ+sHVqa6jZajII28V72KsXW6MoisrfYphygpJVB9zkpYvxPL/aLC2l6B1bA
7PKZT/+q/EqWt4Q+ZIsdzpk8lue1rQzOB2m2tQinfzpwJEzHgQjecdud4V78WTyh/PKq0WDZmK0a
Wcw+V/a7JP5ikFUEXTk+byatPHSlBFjfQiBq4JYLSOasUE+Sicq1tTAsacqUlTPfQk3lOkbxNg8u
T77pCtdppb3tJD4Xj9vu2AYFTQ6WRPx03POOomqaB3n/AhGcjX01to/KzGH5PLQ8kbktocdUvgUo
B5f5XY22yqh86uUsgUZF5JjuVix60eeoDDV58FB7eW1nFb01LDnmxHT9PB9HZmJhTJPgfFJ2KTSn
ROcm+LXf+j3WuPfbzH5CkHiAE2Jagv4uXfDVsVqrQLFbKK/SZwPUCX2f+vxjb+wYhgqFWhyyz7qz
rkK2yID0e3R6mtc8veVIqNL/jlhgld9kWdm3d8Xo98Ko5P0MHuzSgGjBC1oFT6xLXlAbHRnWDxp2
TAy/b57qdlAU7fbv/Vcvp0tkJfTxyFBPkJVX9lRIGxhdSL8f4u5KJo/26j/W703AJuY3FbvLZFkj
nR8SYFX2X4gRPdfnGe17YDRsjKaJh8ch7tOtIf7YVSxcJfq69Z4KqFvIBTFsR2ue7RaHSCsVz4c7
bBv2XW+H8mEAqdiF0RAUdzAcocIIgmtjQTu6Ual/poCfiie+v0IAmLXfcZqrm4dUnffc/TNvLay2
oNZnVrEQLndlQHh9btKWt9nxFdnAssX7CS/VbpxLvXObT4RCeZ8l6TGcXnBIH1WM6F8Wb9/8lH1M
mGhIHpGYdDuHAo91D2oc00NXC0QZurzGuSM85iaecx5I8b1MkoKYNl4xZvswZtlBaaC350SfKgLk
vBtUedHf2FTbMD36to3Vbi2w5fkPMzh+QET/+TRhQUZETDuO0KQkF+9a3tBfa6fme5BTkR3MAP8y
uklOtYw7c0J6Z7Ow3FwJHf30LLeM7Kdp5osFlszdjE0qKOdrTUfFmabYXDW8kSs9zL+zAP13BmDI
ic9jPXgV4XHomCpsasAnqgHzZb61mWYDOE0CSPpUqWoR9Zq/UZsLjfStZsKX2X7W1ea8Oab8iTBp
CCE+0kxaipwJhc2i8axWSvM/lIfv8+SjHBjOZ4a0HNE7xCss0PZaMhVQh4c5n8uvTHdqqAUJ0hiN
aY1V/VjgjN3tl0M5HJRmrsDfz0+sKu3oThA7nM2fFjcsOH4oz5LPyU7UtCz6IU78cnUSiAcKOcJY
2AiVV7+x54jboqIqdQT9kWXHvOqKHQoQtB1EVCso4K0KF/Py+AnvdTVIkEf0QsPa19P7g00gycOI
HphWzMrCrduaWNrgNCGLfAOBHP6G4PcIkfUiSWq1iHvRzyG6C4/DVObO7divVARRpwKUu2EJrgpu
pjTbmdWbzvE7WxXH9JeOdiprr6e+6nOCQeW3yTidE7Q6cSOQhvNjo533vSQPdswKhBUl3Y+3zqHJ
yDsKiNj45xpEIM7+jfaz8ghWpDdFKUINi7gXZJo7CfACID0Gljdcf1xHysOp1FTsqla1FhGpLA1K
r4VdZwYlA7v/cp3uvg3x5s0Qi7v75e+hjtq0dRMhkHy6uY6zUu94J30XhmHJBci177YG1sACi/Xd
MKIHX/rgZY8hiKX/M701P1SO+zcrwdZUvpqDdj+4l8TnabgD+SuqRK1BIYX8y5SeyFGNmSX7dkBU
LnmCneQuZd/cXUgc1xtSRDIQ5dbGxyLiEsYvbucP1sjtOjkhlzlWiGtEDxOFvjUW1Y2MSrYzsFsO
YN00UEYRpjsPby5NyB+nx9iIi/DN7gvkG5uwfbCcHrbhrCpcXMEMKgLSl4qousEXlWWR2ZFbLAuo
i1Yahr4ig6cqdaXqWRK5Cf9t79qcyXY1ZKXrqTKWqw39731j/Vq20tbwYIbxgaPqqYz0KeYMMJTO
S8J4GnHn5uLs1WyftsBYAUv9hxV1vuzzq7zK05d+drFu68uZN5iiPVwA4GP5OHv8icpa3Fl7FEdl
2mQKHXZ931LJjjJ7VkM9ofUfF1kQ1sKbnaTPGtjhh7bLX6T31+zz5Gi+VLXi8XA/dbc/UN6aopl9
dnGC9A/gaTM0pbHGYJR89lkrc8omJ7ki38JNCrax1/iaXUpYIbrEAXEjLxzBmUoIwBDhngC5i+fq
DN8a8kLIrInEp0ZiqtcpO4+slwmXipEwlHXNE6oZz4UxGNEiF2Z9TgS4lgh68XjICE85pEnrB594
y0NhXG4VFoXDBcdr/ZPtKM/2MnhXG9LxDoFUJ+wegSJi81D4kPKGJxiJ996VYBTwrcXBcCcy+L+v
wjbJ6MSsr4IJS/lDRp3VLnM6x1ANFcNCz8GJcOaY/6F8pPBJyxm89ijS4U6esxY4Kl7mvpiDwTQz
GWJxD0kYkO+XhhT0GSO5ECxOM+lf95oqqV0SeibWJk6SJglFKnSZnGBH1xbUcmZ1ATv3MC0BlT4P
8iKL4MGDBufImsW0Rwq4INmdIng4XwlYjHjQ7YZDS5S4I3E5qw4DP00V1/9OPm/4ZSr50hEFJkjT
g9djMrCfz6EDvD+9CRWYHvj4FcouesJVF9MoZpeD0qn9sQ/3OvN1OVL8O8exFCCeI65foGhoMz4I
RnajhP/WigrtLN6UCyEGglsi5bVkK5DfLAtC4FdFA2KILa1Sg7RtaehsF7stOlsu+cXRkOvneAzJ
s41vzCiis6Rw8Z0aQgpzbFi1aMtXrWpc97gxkGMGMYFw2gmmtmTzpsPQLavBRM3HibRdTYqZC75G
Sx8xeJj0Zw6BgfNiYl/fO0jSfhAW4WDGD5/xjPgHU9mdKYm7lpHE3SlbqT65182106UhoX8CFJEA
1CDTyFOW9Ykc9lqVhWOoJwgZvdbqgV1tzlfsV8bX60biFwkiDEwn/45hYvTkQEXpO8iJHBoUL/FA
Dv7+mwSFqfwb5VonCvVqhSfFIZDZ9Fw8/BcBAV9dgybV/ucKyOq6J6w//aejyjgh7Iaj0tlkhSU/
q7bFk7dwxDwuvlc1BZt5Dlzmziazs0Mh/eaf8ORg9jQohswT7wSCotDjzJK0kJEvOqDKeQzmOYGP
F+Chck/LUO+rNTVyAW6zBWtiTP8vfXIPeNCWmdoLdsIgLyIT2gr7VC4pSiHZx6EB3frvSkb6TomW
pqQLzZppR1aG/t+WdP8hclabnktaryH8t8+VG490ADGAI7tN+UxlwF10R0z9i7he+nK3CDltgoTa
h4WeqTOb8Rk4MUyj/i2CgZQVYPz7Ikq94my/+gdgXi6Y7zowCphKupqjvn5xv4nW2gR9ac/N+xVv
MQrDgy/7eLCdMUrBos9rI309c7RVbLZ+d/SzDLO/AUyNBHYm/L0DsSKKaok3jKKmilniYnTM3IhZ
/9+ZU/+mLuds8eAMP23tlQ5knYZFeCvj4CBw/WFiiXTMzey+VxR4J8+F7aZnZNXSFIMKv8fsaifF
Dtxy2bpqgwQyybLlBob2Yi55hBpXWGis8rYCVyZ8F9B2kPIm6scr1TojSMGOVSZ1sFEi0CPjqIdU
wEbn4DLrVb6W8Sz7MdcTOlKG6bvQ60f88glJBhCYd84GuHU3FCsjneEe90qsXHp/xLpFfdsia5CR
rdeUypoI6cdwX07ttS6TCJqaAK9Ll3NCsR3CbBYBMdBrgIXJhx2DWBT1j270aZSZ6p0LqVIxUpeo
+2ghJhmBPpJA6xIDQe+quLomS5fcNXUta4ib4e+AHddlPn3vSt57rJlQElbVLY5hSMH1uHVa927b
lbc6EMZ9xBKA/rgYjZnArEgJoi5CsrXDDSXxcnHNixG1/wR0JMyCSDXqunU+vKqWq1MgqW8Q1mFq
aKseduRHr1qmAUA5ncoK7Kwtz0HexAk1GcX5SzZjMWRoH++dTC3NcjUuBYoU0gCZ0Owtgj3T/Pl+
zmwaNwZ9FASUv5R8tSgX6FOCaA645lsr5dsXIRqlY5JXrUfRTqZOfw1WsuHdXRr+la1tykliLn+t
ao7oWmbqpuCp+Bo5QyMHZshhH1F9qXZVKEMLNmuZxKwcSC4tfOpyYWeHweFuDsDV67jQvqwgzohL
Xkp0fgeH1S8P/vFsy3Di9b6oArFOdJ5Zurbx+ZOHtF+dAZiGuqOR+t8LhzkReWVI5wVC92uOxhXS
dAdfz+uEyWRsgIKzvLf8JsLNJnJ0thyvKcikMOLEa3Y16yT69AEbj0whBzgAVH6gWxB/0NlQIfHI
GI93CrgNx0gYQnFjYcOM3aEyZiFSkX3BI92mqW6B0nRAsdsNudMZh+ruXCbPxOxOFVdNyXmic5Bx
glbucYqUVzQ66INgQzg9pF/5Z5/91AT6pq5B5xAExd81RO3EsbCdrnw+jS5kkqvIC8eHA1HDv+bb
G/BI8Cq0iY4FQKVcx97O8QR16hUrOXvnP0aEhMPnkm+SwDwt4AEq9Cg35sUzZunNyYsLTQ/MENJq
dxgabOhPRMjzcRo+Qbp92C54cuzQQIOM0gl6eqthtc713cEsHsGU7sdtwh49uMrLtaRE3D5MZ9ZE
2bBZY2nsdOxF225oXphN8IWCyn7nDP1+Ur45d2ph3/ezCpX508N6T6hfFSHXXZqMAA0chsHArVA8
qVhKjL7FxV+pIW4KsndY2svAFCag3kxaxYi6VLju6WZ1q8Jv/HnVariyq809h6xW68wXTiPL8nAl
RPXi+WjFn6axUSwvU5vYDGt51Q1A2oNGvCze77gjGXviTWCBm+D2iLOs1KZNd2tpBj+/AFHUvTDW
fjgJCWYzvEjXOOtn4dv9DOg1Pyl/hhL1JBJxZ+Pl7Fi8+IJfW1Jqp+ocgrV9ZAsHjIGpEp1fp92V
BZEP6TwNt8NGEv3kHU6l2L9H2SPL8XZPA5vyI+hYS7qG81+g4js3AEBBIh+eLf6OyB686pMoufWu
rIPvSAZagcLELq7g0SRbwH+d84SBZvcZL53wOOoIl7goheRDnltOIykqBOOTJF0fNknFfQYHCek5
ijN9JqfIPQJ641WuahLck/V5+H/nIsxG4Hve61n95Uzs3yHYdMBY0xOOluIzYuEwCr2lZR5gFM6F
rjpdvypW5iIXoT5eDKVFlARzbJYGPKRxZiBSjwQCF00Zf9K+uMVbqa/edoiGORJQsAgwqcRxU4Cm
lTItgujrv0rNxlsCzdmcxe59GW+I51dL/zN33vr5d5wKV6xk+IvxDHBtqPv5F9d9ECH6KFgQ2p7o
Mwq5aioPq3yqGXdSfANAJOQuimkCir2Lfuup1n8mHYvrssVlGn7KmRYwjF1NylgQmnxE2wYJoZ+3
+SPAnrVxFSWB5Am3D6DkFyWxdP5rBn++y6u973QGi/c2Beyhx73bMavpLsNOjwLQkgkYzruJymDU
uI6cHtj/B8gBtkHESz0xQdkJupas24Zmy7VSz/uqbN+zqtpRcU2SBXUHayOIwdvt7y1mpGpPygar
12eTEmbdRa36FBwtK0NVI/X++A3lnXFxgugUZ0hdZjR1LH2gLfL+JyQTWWreXmRSertTF8dE3Uza
/bH4/aSR11HF2p2Yr/TIhTu9Gp3PHN3cg5PUmMKxPc9jBTMSXtXsKXubGENs+HO870Rc/ErV4HTQ
fL77p1vbzXquzJlowTYBtz6yPkOpJYeo8sIK7y0FOGY3bQzX2uwWyUTw+GvLoCqle0dFVZZdpcFv
rzhMuv5hD79I/UkATpSnbhPado2UQJt3Zk5wObmXaJp+wVw+eRvf1b18Th5s2WMrGMiH8PUmgr/l
bmTtesDcMJyo14JYP96l98Q5rmQhHvR10epBYrb/b+VuaetpaCdBOUeCKcX3tW92ZXMqsi9/wvws
tKpdBBUmQicxWikNEKB6xeqJBB/rHpY0xiL6FpTMONjqxdlDDqPulqbAmOIKgsXF8YS8Cn2uZrCC
bdHFxNRHOEh/Bfw1Hw3P3Arer7vfbTXHS6nx2HX6z5HT5sJSEQKYb/dPTvM5Q2AiSxKfV0PbmFGo
r3gl0xFvqz6Knzb0CW9QypPnB/wREIDeNBg8QtQP2A2/7boDVgELQa4S0Nu59naDV6igQ4FTKPi/
Z7J5iTuBwHe4xQOFbStM+4kWOglZC9i6Alqc83gwpaGgbqxG9SEb8UrDd3N4NvWkqiQi3imyv5Mn
gB9W3vxFYjdyGFlOzxPp7pgUdKSSr1yX1DEqOGK+domJKgF0HwqI3T7l89ss+Nkl29A5AoKTF/tr
JZXBJ1iaSwVdBVK3G3/g26hBLrO9y1AI0EMpFgXbervglCvJqDvRdKFwiUa4ODT6E0NS3/qQwR/s
q6GU4glhtphfMH349mHVWwSdN8lMGXK51l2uAhcXWwIdW0eMJi8L+PCDU7kDq0tptVF1cw2CXm+N
drDFtZJW3fuvy6CKV1UxA6tUWuzzWLihCKG7otAxdzMCypOpGuLuat0C4aRc/MzxPrFBi6RDLUB9
QrqCxYeOzo28huy701QSAyqFdvmcfeOgkvLr1g9C8xYuUQZhv3EUl67yIcAmAe0N5PPTL9F5gGNs
KoRvW9nwrR7hFrWKlqwfuHy+LHy16ddewm5VBLqhnvHziOHfbHDWko89MbbMBAOilrI66oaAmB3o
dh2+u2B69nM5GeLsUUzfPImyDyHysroy4+LcFNjFfaZhAR9nTxXJwJMGMN2LS/burUXO5Fi3ALyN
Li0xLbMsBk2/eDQvw4WQrr9D5QkBywL69JT7+zT0i7eZIjOz1wOBg6DCb5a6/sSzn10yzpcglKcT
QyRYMLJ2Pf9CYMeK9WhLS0oJPNaFUhMcptyRre55t+3TyhxLMXGjemD7gZtGYLlWoKaA0m8s7uR3
FFmSVv8a0xkOQHvySts7c8zZ3PylDORZxVbl6ZBddEL8K2e8n2We6FUIHUDedGTqc2dYefVe2ZTL
N7wmIn9GiDdg2LPqHqNNTgKHeDxbAFfdp6kCAZkdWSpTyhxEhsv8eqLwyi4AGsdTnESV9DMoFYtP
3ytasNQHlk94PFhRNtg1hIGEIzl0gcDbSq05GnlxKh/A/XnMDtb+by/b1kWp79wyTvNy2iTGCK5N
4FrPIafy1A4PPQmZrheFtYJREOOVc+lidQeXu/V5Zp4p/nYh48Hbug9RaBaTZk1Cakqo0u3BEW33
2YKn1Hc5vbfJ6QIPG9zMzybgHvT8UqPzoZ1RqC9nu4T7KqMi5yCIpRJh2xsnhekjMsH176Yc6rd4
feqm3rT0kQLtNXP6EvuHodDOC3KM6DMGLs/5JkxykmCInqZ8BVRFMoBPostjMSuQPQF/ASgUG6gf
p+vnJ1Vu1giup12roqtmIfYjIF1E+sMzPpuBeEUt4YJpxSz2ARpo+Ta+pJNhgAV5T7UVfHKOwkRI
DedpOcIkflcpn3MaPbJcaLI/uoLzQWjKvOyly+QqSfaEBNFhWOXvQAhxI+cdJlCn3uBL8L239DzT
T8M+4CQT+k1QoSbo9LVyhastX7VV51ek6cK+YB/TF9Tos/XeQzUAuNGhePPXAlccYrMXzvAkaW1N
Eb3UpHN+GIPnqfEUK3lA9+QnwiAGZeMkElmyI3ULBq9/ZhHTY6RkacHhrJ0IV3W2Q7v/jBFjCPXW
QHTjOO26OxkjtLlaf95hsXTklF4D6xJ58jnefHAlo61QVZkpEW/LoBbLyRgYNXzmvLvFZOllplMq
TlwR97FX7nUrYNpAICCibIvNwvAhql82E2Sa0R6PpBggNpvsadFlpsnsGbHPHOuyr2NCfASPzy6N
6c251QrgoK3K0GGrNielereXAvXggct2KDa47A9m5iIwKrzaFbwYAcETZaDq5rWWUWpUv4HNHVaE
qSM9o/tbEx3SxOeUuKOMkLXA/Ih9mZevalbhYp6yu6jgSN5pnkfTMmMw0QNlKT5I3Wza5jW500Yf
5UZ1j+wOvK1Nm4Wwf/bK6umCYkujqGCam36sqfhwPbv4zmT6snLiYN/6PXmESESlcsB3uLPxgnTV
JjW4nrf1/CGpEPGLqwhFnOH+8ECoSWMCltBahSWh+kxH0yNyy99I5/GY391/3FbcisfUlgosZJ/P
z4BX29jnLnp7qFnoOBFY4CDivUamn60RzXpYJBLptVlXwoglWxjdvQRn0aWCg1aFJ8Cf3Mj4Vhov
ieQ4wFTANbwAuAJSYjwL2+aNxugEKxcIwyd/KRgtVdHhNns2YIEjzQrmMebOUlWWn1NkUn4SOmsR
yT58plGzNELdvMdsHrmstkBO7MJ35vfHpJLEDsIncGum0hFHNrpfXF59SkBB0ppSJl7eaCE2RCKC
i9nGdU/gg9r7BMfwrmDAKACQf0pGXvp5ddcQJ4KRG+102ICNhm6SQugNjscFBs0IXU/2wnKbVh9L
aTzq+9ujXUhsvHPkWbtXrX8acMvRipvKWpvBnxiEqB+JB6uufAZ/x6Ro4jfURBc3I7oirkVcy+t2
stmJvxk3eUpMuZK9vjGlLaJaklGMBeECdr3i8Vat7D06D8VQcmSkOkoh4yd3VXO169wMT64oPqit
+5ah1mgvfgrrQ9HCX501Jmn4SJFaxXdlIC2t3xbuKPjlG7CQWxItRpyFCbs0HYUjKYZ2aqcDtmmT
sC6tobH5aVca1wAkVN0Q0KZbSEcyXNtg1AN/gy9Ku3C+K1zsZJpkRCS/EuVxewiMy2Usyoafaw3T
VP4walpJvMEU5GycFBiUDV6AizH5wbQ6Q0hV1kmyJwBI0K+oAwjjVAnQpUQ0Q41r95p4RQmeXLWI
p7dWjcysw/cQrS5i9dA5UeYLxNCPUWyv4TtfmZuLRhY2w5MfYgPj35aThkiN3TbCaluWlr+ATpzZ
jWFI5EM5rwaOHGJrL8o0VOK560AQKKVkwOY5lX/yZ4+OSdVUekWGh3XXaaK8UdgI5bJLcmtX8PoB
yzQdeiPZETUe076XTqTA1ei1KtnqjekS64XpOzx8h/WmELX6srOLDUHBr5odKUbSyw8Vb2ivgIFm
9QQqjt6AJ9Inxl8hDYDuFPNrqaPBJEOE3MAP7qveoT90J/irRHLMsulsvU327uF8nqE9exEbY6bx
5ifiF2N/H/IMIUlOMEOLYOT4L0p2qvtxITbT9xh0oWvk3fj/VFwyqryu7fEdTyyPANpjUD53qsgI
ogUJIl1PIA+QswK7G79RWfVeHK/Zsq5ZNWcUyalc+DTR1TkQx0bJmsFTAh/AoaPJzKnp0ARR5FAB
Nrza2rPj0TDcEpZ2IVZQ7ZBt5h3QCU0uibS2lj/zuPaWYYPWbntFErxlNN0fYVsu/D63aNEhschL
Bck33vNt8JTCQW8P8xW281OQNBpS27hWC9Ehbih/ERHmlnaSg1/VoeRFXRdAJtwRoZx2n//GztsR
gMp0S3eCioe6zHFITftDPDDWa73nT0NfTidrNw9yg3tBjSyuqzbg+qUeUIC0ZVbUqRNamK1wVDAj
ioKO+wfgpU0+ctTw2hO3Zz0G3s4sLRdBGJ4a2p+erOqxV3rsY+XqbAIs/IVd+0iZvDthSZ9cGvfC
QE3xffco7Eb44UDvV8gzxs8nGu3VoWQbeQpPt0q1kx9EbAxqTMZYCb3tMaK+mWVLAi27s1dIMNOe
qKIuyzsUkps5b4oCSXODwi9vIBz1OYtFRAo8DsBFjYwmbrAMmb4euae/pzxbp6YUpt7VWUJe7u8M
udesRIukzn5E+vAaEsSjsNmzY32m6sK5XPHZP+uqLDhPxD61y4jBNd6Jm3U41lG1PH1l2BOtt4nF
ockoJbMAzXId76p7p/3flZTqvZ2xIWPpb1GqOGcmGGkbZH1oRShITiDfwtATBks3oLwO9G9qdGfQ
yT1KlOc8bjYvZadG9ltR6vprWUXjiaYuGEN4bZGH31QHZgE7MY7oYbJSINMxD2V2bUrQN49ykn+t
r5IKEJdWvS4vL396b27oOT+9Q2onspCC27Aka0U+LvV9bR7xyvbfb6AmJ8saXj2jAX4eoeNFKym7
SU0XdKx513Pd4VTJvlT69sdHh1QUMK+1YVUR7GNha6SyFOy0w/f6LwUPBaYlP7eGa6qcHM9KN9cT
zm3VYnDM69nvseVCZILbeDfZrDAVcLdYy/CUlAnP5qFvBDnWE4UvwMAuPIlPes11SufG1vWEI2vE
wuUjO7ihfzpNa+yOYhaTRMJKbt+mC9bkhVn9Rmstr/L//tf+hAHA4/wcyFmuF1Ajj2R9lFYpQy4S
Br9WesZuDVTDCs9qjTedhY2B5Qg2/Tg1H3OX5bNRnMfCIzgqFE7tF/Yo5Zn2loDTeUn92FPPsGlC
aK3gxTeQBHRJDARQOI5dyf4SFo+bDCdc5MoFMbEd9tEPU0MiHj2vm40Bn//wFYNK45LGmq0HuaGM
pL/XRnF93WAMTpUnQS6FuZ60zTfGZs5SOPIOVmZuQL10Sgy7OoFX694C4k9M9qbwjRuAPczU9Q+w
k900KuP0wXN79ENvuN2uvE3MdnYzCqL7gmueUsrRtj706C6vHzqOHYlvHruXbOHVHfZwFs5bONlQ
Wur8Jf5lG5azVylfCjkiE2kD8/X/kVQVC5us2MNJk1jka+w/YmJLCTDYJ0WA3iUbDMZEdRbdonpz
FY3RgAdZleWOzMHG0T/Vu/eKg0DQgJ4L58zhl83xgc1a2ht7Z80O+jO7Mjz/iyi/EIho6r8gBeiR
p7CyMYqIgpHDDkZFfBKfrp5SIIaTIq9WMwQxB7jYyMP7fAIMH0A69jHftFQo4eaOt4JrNLc0it/s
z8cQYX6+S+xdolrlmReqsY/ueZ63p4NRMABNiHFgQMLbbFVWdCxV8iFXbQPAlALNse7BRsTT8BFV
cfvtDl4dBZRnpLSIm2b44+aV7Y0g5wmIeUTprakQ8t+wM41t/nBlc8x/cGeKsWjtifPLhc724wOU
qd89GyVIin8Mxa69i1wYPbk1DjPQK3GAZyASBeChq9Yp8Q2H0WfXCKXjxcT28nAxVl6g1vloXsR0
RaFRvNQ0U92v3QAbv650Sjz7eJXcBYmKj2eycW3UtlpssknJvxwJmj0TbYu4t5tLOBEjC+ixsJp/
q8zzK1eLuaRlfp6Ir+TL6JmdqFvWkZ2LKBcf21fSy8EdSwkhqkteMMXLe0pD/UT3qvC7cVL24BWt
S+gzJQb9tLhxGMYlghBGCeIKPA5oZM8N8A+mPzgI6uaIob6gFOtFtbLoz3GR0S+A9m4hM1ydBLTf
YS3JanCB3d10iBzABa4MsU+DJIFTTfjA4NTOQ4a9o6qjqPdg0oTVuQhq/AJejc6GX6xJ/MX2fl2g
NJFyr2J/AK5ja/vPpxnfUNyBnPyxu+pEfOC/QCRzmzpIUdQxyaEfp7kYitsvkUup5zTB0DTH5J4Z
OLkW7yuyfpu8Zg2j6TGsbA8mE2mAawatuxsVtS1ESRFntrUsu6SNYyr5BIDxUNvLDxNw9Pzka17R
YtLDV6iqIYh10WK0tPwjuE70fL30XJwdksakW6RV8X6kxo8hYAanhDpAjdPz923JyREniMeRBJHG
yGa1xt1uJNvsfSdQexnMTTDWzEjwbbixV4YvKSUgH+PIv6hqTwe/uRJX42Gpufi8u0uInM6/AW1P
PRnAg2y9VpyH8ccMGfsNGmqGXtYlo6EUWL9vgtaaGNk9L+6xcOC1X72Qj363LWw6MU59hsAzSQNZ
4SHdtykiXuCJDyhZRqDtH/IM6HifdipM5fUujar/NVwenQZYmbp5riLAOa5vQnpgLSWSawNdGLkB
ggF/T+5s0eJhI7ey0l9s933Z7HyqLIPvqsvVw1RwMPRfUHt47wt2UZQDEEIMhIN38WKVN5D4i+3L
G2ticLWXGTzQ8uKYWQ5TEO/t3tA5efFYA2coQ6LDo99slwCfDPpWO+gBwxvFa2X1TeDQTS+nn9YJ
Qp4tZP/0mESv5Ae1iDEpHtbx6btRyPTTc//XlolJnKhwbiA94L9QvGJN7veQIiyGUkwkJ9uGPvwT
wJmpwZGPQtr1sqBr4V7nX5QThU5ojDLQL06E7opPYogB+pDWz4V8gdI07kVm51+4A5JRfq69OFH6
twev6BEYXXMGdV+30HjDNQqCqavnYdvuimQrlZDoK041L2LeqVqNiwXdW7lvTgwEib5U2/TTm/6D
J9YLR19WTYw9oBktOEWGPdo0I/Uykk1GWZiONtaY43C270+7Q5giyF6PIr/s5WN6qMprJEbgxa5Q
3DVCySW6vO4kb1ep/T47ECPaATpR3wX4RCH3Y/ZdsrRTi00pUilkERwuHfidCRIzhzLLR4qO84uN
b/rGEeO7pqMeJtnWxUMMreGeq12boG9b/XYClKsA3en/7dFbkRiL5vKhld439wbTV0sZcLAjAkox
jOyqHcq2mua1ysz6kF4unDizITlgYAHLIDdmIU4bv/PgXN231fv687plSJ4xlp0w6z61MSZr8gZD
gA7Fty/PBty0g9MZyqkHqMpSd/YUeqqbm/eSSAlwAQOjsoYMCA2A6B6ycl6hmiPts/hK5TFK7PwR
TLNduMZ21NWam6tOdiPDK8yNn19JqCoxZSCC/8nHSOox0vTqJFLloEjuX9wR9FjJwAXI8W2Rp1Qm
WPpypve381CEGRFay4Om+h8VnYDksGuZfaAusUCyeU5JY83bkW9fQKnS1Li01JFzaRqSOOJa8ALs
qDXJ5A8OyzTmxMZNbuVQxGJf5X3UYFqU6VGHiTtVgDCGuAUGkaZw3xkuF80oTfv2G7JTvlBYetAS
Oel1MuvQLd0dST9RkAfEpz4szBCFvAaBUildLdhspxFnR8xSLI1mLJ3+tb79+l9grXGH4PC6JTyT
5ZiAOb6c7rZwOsM7I6FRy8SsYt2r8V7al6IKmQM8KqxULko5DEreHFk6sTruK5k19scCpYdxA6/x
OeEWPRlTw/fyUIYTUi4ZCajdXi78vapqvJl/n7bXn7IzNbNdIexIogiN6rvX4pudrUx+3ep/uuVK
qmoct378eDjWVPqK69xvmmKoek7HVdg3oIuUAbkSTnCymxVyh/k8RFxf+MCkEUl7G0fCv1IsXtub
ZsvYCEareyOt4de8/P49SPUKSWEBl+ZmHDbyDXjDB6WyxJMeYtSWHdu7Jp9GQ/0Upys8qZNua5OL
fc7YbzdqMo5tOe5n5lq6IW6ZP0dYhgGGduXwML3ioa1FvJrBwMbncPEiWrDpegYHkoqOKg085N/t
z5PidLF2iTEnblG/upXnFEwA7xq4VjcyfdwPTeJMQfmwRsTy1ESfwFiZmxf8YNZzDoGHyBoGUdDx
iV9Beteow53MJyl8Vpf523eYJbegTo1k2kwxst9kmB51cYdHFNOjw6YbVB/tK1svML3h0AFiH33o
bRmCukzPOI9Og/MwZn1paUuWQcWPeVTpVgQk9fePe/b+q0nbZRHbuXwf+niACSHtiRmGWV790Fwf
I7x4ahRZS3XyQEcB7iZJfOC2jY8h8jaKpjAOUkJydB3MZ8JW9PQ4N7agXSIW8i0bqUmYSrdeAb/V
uHaGhxmN6Y+ylmo3WaaDl28ACdTl8NdK1tPWTeCrxuNEUm7kvT10l1TWrrJg8BPTexhcBo5s7/Do
Z76LiMyvh3Sy/BSRJ61Z60P2VEbIxkeicZKxZh2aTk4IGaSvnZ2QhpR6Oc7p/wm5UX8uMwTYWTyT
R6V8A3rJ7fuTfu0+mYOtF3iVaDSIS0WXbBHg4BRVO18OPGYGjGTFsQq+4qmOTyxw6D+pDd7JRFWe
lzldyWvWh9fZjTwwSlyl08e/OIIzAzCAbDRwQfMjsoW3L7MmaDfNlz2V2CebsgF6kfC6+eiKkSzZ
sHDmcnjka0iLhoi7YJMGsqpxTcByerIYSLwWJcSBXdYeuz/aCkLAFnJ+iPMrjLWKSDQtOw6gFsk9
pvtm32EL2uAo1tGHNCpMv43COSyGAFrRLOlZyNgd1x0wj0TX99TZJaUBVsxQNfhskIDkmKMvwehk
599EBcYK+zGGhY/dG3heugGr2qRn5/CQL3PzVhh+QrFWROAK/XcwjnP5RfK+NkdSkNOt3l1PZlmq
iWsyXde+3+x6lgotUhEh0xbBCcFG++47Xp/kFobOqY9SNOOECHTb9KI50s1DagEuY7XuqgW4uY+T
E30pqleEPn1w3KASijvUzuRfUhnSE+cmGWvaOg3LQ7kmONyORWOrvjOFPi0znMY7/593hM77g6Vb
JuXoKOABxb7en2sj23N0aPUHS9mOk85a0CpRT2B9cj//gzQDA+7/RuO5KrEdwu+THrAwvN/p/uPT
xhsNCLjcqhRd5KVOYBvs6cTF8yFZ2CjZUf1o+oFppGwnZdWPLk4HF8VV+/uFA13tD15vuk1fR905
U2TjqIltzoZ4QdzOAasPnVlBeD/2n5FwlW8sJZD1xrXHBz3oT8jgrJV+4nBWbNJ+ehZUNOfH3ywk
L6il2lMcPQstHK0qgOJvMVSvsG3xpwa+GrZDo7otXtfuiNxRvLVF8ugGQQrJEVfmhuCujENRQFDb
kVAbVa2RVhm9EGOz8OCzatRdPnVGuO5XnW3yaPlKHgCJwp16Lqm6jUf6wSa017Q4jiXmyJ4QsBDX
WMga13DE6yuqq++lgFiwu9CV/CmRSh1BPiktO0SUutQ/opcjybFj9sDQmSiy/WWbpDorXyVK6oMl
Hz8c6DWTvJeuJBTtPB5BsotLqsT/jylA08QeCz74DzgOzz2k3HrLsDWYLkoeomD5ytAqbrV5DQ2r
ljXyhSzgUaEGW6CuaSvnuBGQCEUjfM+Paka/G5oScdVbFI/8x2hXv7KZxo2newyNpiMf8zzRC2yP
lb0tizX0mhv8cTKF7Jtnh0X+nm1GorZNPTAs/E8DWpij4AM2UnGfWuY7jVcm7zHZAcfFabS14ol8
wB5W2aLYH6anP2lwzooiJP6PnJWYhptaERQ+tD94vfqYLRAhEatpw5tZY3Ek/jn4gpPrRuNPFeUh
/vVDwwI6d1YMJMhjz7A+GaK/lKvCaidRDrd8S0BxVMYKey26pD3xJtRFh0mBjgYPOxiPBK7HyVQl
zr8pO296noMQ4ntWnV3Af/4dfU7QpL1+PO+JwaEfYThG+bDYcyuPWPGFgIYxs4cFaFes/bFAW4yj
1W2xzfB7hkNSAB/bM1BpJQO1bLs24JqVjJ8zHsrP2gu0VFoxloH23Udvjfm9MuKS75ABTInl/WSX
U87MsuJ5E74q5Hj/uQHK+uCx/zW5CB/J/P9z2h5lOPgEtZwTa1Q6Tharw9QV7lNbQVkcW3ssrhyc
g2DEQCeISjYoTzqiJlTSm0KDEk5Uf3qes7MJtbRv5ChL0aHyaiBYp76v5lUC5Xb8kryAATBnAW/K
y/wAy/ZnVw/jq//Y22KbFSrVCXL0IGVGnvTloPDFSmd+HrO9G8cf/44lcEoiiFLU9G5x3BqKEwwF
lIqUSt29VeWqjy24T/KG6hYDTgfcbK9+fivZoXayxSIZg9ybLQUia11Lh7D+WxUgUoTK5Rrx3pAm
L1/SQDrSqHytc76LSgdO11Z0DdmaGyZbuO2OAvLuPg5uHIqaOLbzuMhRDwlc9GtR4/j9zWCjSQmh
Mm3Pm//2IQA5lMqx5+E972nCPgQHsMSl1dIZU/jIIaYiOZAeme7ZGi9w2anMZkVN9vcBjrjb/8QR
vjZ6PA81Fx36j+cYRt+pVO9UTBjiAzAtq/Df5iN9jGH4eaIZhQHH2EVKjeIEw+HU7EGSgg9DaVJe
VcjhDvtxnylAPS+dMaZv6oRDlnqEPfFqa6Sczdv/tnz9Ofpqt7I5k8/2tS5OkQ213VHDHtd8VmsV
jKmHjnI7ToghfUwGom0+8zMpzzXWv24OTM6JxwzJidkVZsWIuMMWlmDtikbeSan/Ium3plGQvEBv
srvW95OEjqw5MWgotUfhS6r0aP8YZn+eojyj1rDgY/x4I2RyMjWjbjCACKhRcrD5WkDZcIkMtcHG
pgM0uXY6OaU159sO0qOZ2t1b2PMKFyOYqkSEtNGO5MTTumx3LXlj3MPUwq5eBkPy//7OR4sIvE7f
6U74AFY5PkHtflrKxl86q0wiYp+8q5un0E1LDKSWZizuYuQw0SboZItK5hIdXMgaRR4S1qzUx7L2
sa62WpzsgnbZTcoVS3wFM3FVhO+vu/gt0L6MSAuDchZW7Y2L3fseBeuCWZoOllSF6NEjRg+3AJQ/
nbI0hHWmi8d2fCW9r0Dys5DkLll+3yzOx+9paGkEFm1mSAe3xTUIXhgT2FelML7o0Ms5uDtJQsYB
mly/54C3A261cDyFGDcl1d6kQ8dD2E3Pqy/C9blfWA4pQX1Ov+d7vDBTrXTPS6pFO5QmhQXpMdPM
mhRM8IPuZFh/dLOBaC4NCg5t9uhNLQMTjgyblivQ73qtGQGVnoKP8qr2HIExstroqI/UFyURCFGO
F64r6Md2ZIO995OFFj2xNOR/UUy8bWuaj5QKzxvNwgTzATX3IGRQrWMFsy//pDgHnh975a3zBi2R
xfyxzu4KYx2idFVkkXBlTPK7Hld+wDr1Jj2ZPtLxh93AM3MTjiUWCGzHuEv9IPF6dTsrl7Sy3jpk
1BdB1uuyW43gYLttQvew22JAmzinBGlfPa0UI82qQ+fRy0itKtgBEZyYwFDvN1qFIYA/1f7T4WuA
NwgYN98mqvoQyRpYkaal1GTJsE5OVlrGjwdQtLSKQPny9SWiihvh8qlkFuexCFBasnQvAvZlKMJB
kbtVKmsCpJz2epceNT8O96I6m5fomcM0uv3WMayeGEZVrEixj/KA/8CYx/HO/BSrPPlLSv082Avp
kVw8nUA8QfRb23Vby1+GfsCrwOW+DksjOmKcr3+1JZGaPVCwWgIkqTVTcOEwtK70In177WoB4F0/
3Dyk69MGZ7XPr/yoswbpE2EOSY4f27VwTEq2lsxVWyG3WgbculY8js4ZdfylJj99jn5fJxbYhYoS
bw7DamJYZBOIW+RYqc603LPaOx5YG88gegOWt+CGFI8ZqPdVxfDG9d3hxcJFj5kvr7/iOCR3KyOB
vh3lIfRa8ge1+Fcz2kekxkg9m2LAzNTI6yEwFGm0lxFOZTSVbMJtojQftRLbN8+ricTzaZYT78rI
5+E9PNV6iLdPP4uxtNYnoFAH89Mr426TB886tPAgJzH9Ca0H+SNdOhyzVn1whihT3iJ3RVEp5ycQ
5yFh+e8mS3dtL+DNvbBVRjTfBKHzKyRuV7PtJwjFc5zXZChMc2LUfvW51xERI36Xo7Hw8zBi5WDj
bNWV9FxGtg0JQCIYa28Fkm3aB3fQxHMn5IF0pDxvQ49ljP+wirtXjnRYEwz8NArgkTFxhbpEKVqm
VT3hpSSCb32eSkEslLcWQUAfceIRrQq9MI7AkrEeSmF+/OR7wGNPNa+b+60e/qHEtsDdpzwh/SeQ
+gXc4F+9ukrFSjJIkiAuyrriXA/XLjENsP7miUmYpJFbmhjhEeZpDlfgSH2gQwm3lX+yillxO8iz
LadQVDGZxD08xznUX3gcriuboO124kgpThdVWMJvgrcXVfkG+i9Hhb01YECqWHCWtVqTStuXCa7G
eBrXirlVBkzXItzds8k5z8xrgMYw46+taaibUW1YVG9MImKGDM1JTGhsPYat5+ImTIiKpHl33qxv
wDDapuLjwwzgX0gGl62fMfb7Wyo8w3f2H4rJbX4EFiQyoYYUPW8clVc2nD9nKtyABXfScaojZq8S
eo7KSmlgsO9eQYB5RXLAwsHQQXA2XOnBBgdbH1HS3MC58NOfXxqy8t6672g2RTXna7W1hG+2oklb
BjBNiVNeWPmaKjFd1Zt2fIoApcdETmgceQmXtd9aopJkqXbvaNOTlEmQxvg/ye1654aWhUllvnGq
XRf7HkUBekRj5TdmlJgmZWNzLZSpLGUSb0rIYjQjBb8e6iWfwzgBOgXLvxYnjlnxwLaQxhBellrx
BCO7SukcEb+8OfS5Aza+4MwLhZdTZss8WJEwgoUOjNv3XEN91+a0jhrL0dvS01DV5nlmg/L/ENUo
Y+b2a89mvvPTVO1kqVgtkgqb1Bt4CRWv2VfTpNOxm2QodwK/Dhvs/4VaJ/rZWqcMJ67Yr2IarySZ
vbprcUVefZCeqlA3iEl1C/4Jvk1Fxb/s+bjbQDlOz/6NkD2/EJ9ymqXagd1MU1+39jpKAnJ3LnN/
Tmo7/cJ+ObkFyeznOeqWSa5EQxtAdabYXSx9Cor5wIjY1N93skHV3Igg3s1oL2+obookZHf14MwK
oqAPv8lsBD+Vjlu0ljz6VmHO3IhnYji6oWmmEzZ523kLbsiduxmPGZBXWLRzawGCED+HWdFcDvI7
4g60MvqBrC2cjiwU36mhAL/736iteF44FmuPwWb2lucp7plZ6bpEPDuoCHQiAA2i/oZfKZmPtjT3
qz1Gl06zpGik/iPwEB+dwHsX2DNPVxGKhUhuqLcRwGoY3JL4gyXcV7IzHzHOS9y1Lu3vXzHthBMG
y1WDJ2PdX2odrKHi6d1oGHJpuRRnnQEJJXYmJiu6L+mybuKOmnY+xFB80A9FyPQuO8SF7MFqCKj7
bq5zp03vm/KR/lxI/QfVhg3/KC/v4ju0NU/u6HjWv8adXJgBATPb3KVwYpBRUhVBUgsr/O8k9UKB
+N7K6cWE2b1FUi3CbPC/oAicWHT2IFHtyRT5YrcRqxad83HWmuO8nn3IUqnzIGPNGKh0sdg2HQVh
t3d9yU4yYHeVPeV+gyesQA38x+PqNvxCG+l+Cgdiu4a8CGzQ73ezt/S8yvyGqGUoDZUHG5ab2MR8
UW9iCLEVfZzRxjQwn547108qmZDgMPwjY8XDBpFPsiuPpW0dDZoOu28dCM6ZqPH/yi6ept6dKIWk
BwPJGFx77B6H+hwTY93USXgz3eTtrMruFgVDauaFD+We/svwlJsgh6VMDxqHuy3Qgt/xX4DcMD4y
wZk8e7dh58NWwUCoWd7oGRGarzSl9ReJpCUEoCi4rYEFbHdJxSJ6yizxfz+on03BUgesX3FCT/yU
JPLLNMKa5IbJIIHQ+orCBP5UOF2I0gIV/6NvwotQe0ZqEObY9s6JTE2OIQ/yxg4trbr+yMyKVqCm
lA9bL6xvGIhiX2IEISdql9vOJ+hI7YSKg3SY9v4te8qbWFZykNx3qAhocUUXE33mp1rBGx4+RLNa
DJcWm3f/QcIC+Bazr2bUlZSurmfN/Yr/DzxPMDzaonsFyshjxYQ/mhd+CrLFTBEqxG88gY9mcvbi
XeQm8TCUIiZ7pveG6SDDdqYlH67L7GaWW2HO1H9VPm0JNo0IqW0xICwgszX9t8/7YUvNGwn9kIAY
c5sx3Ll9ZbQaRwkdeNogPbd0D2uHGua1FnD6obla1wmzZC2hn2rxmH3ZPBVx+SDwLzkTd6c0g0hb
K4bRK7fUsLq6ixVVPN+2nK1J0IIwIh2T8SHmQ0vnCWLZpPRbG+gS2FWhOqF6EUz5lqn38k4Jn3n5
vQedSmoc4+c4CkHBhA6rdEA9D6h/rOaR+9MnW5vkpDgBQPnHhAKp98DJNy9HHNGQaluJNBP65pFA
SIK22p8mmcrYdUogbYKZAp/80CkUUpH6WNDjCqIbXpNG27WCGyhyAot0t5C+cJk/RNWAwv6xX0jX
DadH6pyemirCMpcOEMQxCL3sKazafx8hSfnx4xr+1vctsDWqD4b8LZAXpeZ8onu9MuZBmt9GZlyr
k3mCbJ/l1R+OMwkGmenkG0vLQ3pQ6iz2ykVxsLWiQK52vlkT481suJmnTfAuTL5a99ENp3RKxxO8
0D0MwcOEh8S6m4ntkVxzKNLmFeIrbirtC5MIGrv4zQO4w2s94YPpR5DWfSn29qBuS6Ow6feSlXNP
mbSxTY51MlZo+5lWzqYgf8zCPQhG38gvrRlmdJRpr67t3WC4gYzNThLJrfavGivpJYyDtMvua8qP
glNiHzdYnKKcKjgfMMpir4pUGbpokgeZiHT6j5VHBz+uhmW72SVuOBNE3aV0OFPxqTxQdFp8nSWg
FYYV+Di7cW9Eww9w9SgmBaJ7uOLYnVL66/qN04CPXcTOaD34dqYAvClfI/N4KeAfs/hrQiKBiH1E
/1e4wPSsc1uilyQ4ds+XBc9U1MMeGDSFgrC4t6QDInKGrIlFrmBkpB5zKq6kgdEEy6JROA4+Bl+h
PcHmGjchC5mZ3j+EFyIhk1jOPpWl6tf+863cUXYBOsTG+wjgobmk6J8qDFrf/Jm/BISxzrCF5Ynl
zvC7pxXt+2VEN+Dy9xwr+CFqMupP3naltOQm9PkyeZzQPPCsim+Wojt9tE5R4em9av4YR+olzg7l
SaPAsO19p29HUZIrZoGlnwPlFeueduJW36Rc0ScJM85G8oIXd1smjTESzl5AXZxEV+ezQH7b4HVN
De+z8aD8irI1TEBr89ikjRv0F5UsZyt2WD+VS7vzYP1482++PuendetBm5qQyoF9XdKdd6FxkoGt
5zVy5UKgC+ZqCIIDQGL50HlnE4kHE5EG6KUES812TDdn8Md1RPhOV7H45XVcKRf+6dmxMd7lPBVq
Rp2xjVJWObXiW8R/41lKDFNmiZNZRmeGb5W5F1gkPR0R7p1ll8oR27v3RVujKTwhbwX0O8FnFsGs
ZReemJZBl50qDr5DbAzxqInN1MQv99lolPqO4zPQ+LwyzqPTJcYm+vRql9JhhOka6NpHVYB+HQYL
9diaUMnoVUHhu2aQgIEn8EYzcgPwDxxSLGoV9WG+ckp3QsHpIcx7bzrYQIa/xm9DtFOvFvQcVdmC
JWSZfk4eghYzBwb1PzM4baudNHCvrCgm4fyUHpDqotMaHDWnQL3yu3ujBCC603nEM1PfJKtYpmqV
yDQ6C3QpSDSHpIWSHTpcyNNFlSP6ZLBZ+vzWMxI2X10+nrrj/HIFv4yXXjQ2cm9XdGPxJLtEeIUr
4vhicTjMy0UJEHwX2WxMDJF7Oc2F3aRQligqlnaxemcwOoZ33Mi0b+r7FhfjlEw7f1WNa2cKiAwc
xdsrvYDx1B5mZAEqXnsqUgunyUNO/40Jtzdlbu02cGd8ScdrtvLQzCbEvyx5xITwSuwLdFE2n08u
0jQlpTiDfCb2zzHqLEnmYuA85vLzW0rErpcHZAuCpD40XcFZmnjg2M/qGxOI5KSX4VPin82VNCKp
Iu/SimZV7Fwp2tzZi+ESlmxG0Kyn3TzZakcl0KdehMeA3ULKjXMnoKJYOQ4L1YtCcV5JmOCHJQQW
rm4FsqRqMN5jPX01Nk5MzC0H5g3xagiUnLrb5jY6MEN1+PIOEU9wv41uRSy7ZxLdBF9/LA8tpMBb
AQYWlqb6ViQbrWD6XgVLLLQ07P+h48G8A2BJrgZJ14oxWSTyZy45DY31Fgl0Q6dIDXzgyTr8LfwT
EDNk4Uk63BZjIFWz6dMgO/q1Mr+pNzDiAlwqFTzTqlq/ApGD40NbCc74ReNj8bSDNaZ19FupMkt/
8IMJkLf/XSDqVS0yUt70ukEe9SkfefHCC/voQjR8/BHp2DNlztgufxJ4I8NkhwokSm4BBFyxlATp
RnouZ3fSEwvAxYCseLvJMFLbP9rrlxoDJIsZwE56iV9ej9fVVGu+7v0SKod4qhTmFdfQGv/tJxlm
m9MHaqT1P+spx8sje96C5JI4x1fb8t6w9q570eqIPWK+/HBnDV6uF0bkNSWHoeEQe9mf33e1Ok6H
jIJLXztOqw3igN62kWgaGWphx2cBq2TKz9bS+tE5Aw0C/AsTAtjaDxFBrq5xYnyXQ8AFf1X6P5hz
5J8gdjvqJfSDi2BMOe0gZUN9LSiXovESr8gAKGKUN+Uo2sRzFRyMc6Z5JRaOpTvohwc8vSzsA2EQ
c3kM8drcv+kkL+DpaycwrmcUP7QkvfVyl7A+tGWOEz+ild4kCeCDleQgBvklOkvZCAmllSwDajuN
IGnpIqWpl/Z+feahjtNdyVlI34kvZXxoMDRqKQQptp9/EKahvSFV9bqz9PsYkwMvRqrhtGwTtMpe
HVTh91RRw2SXTzkCYF9LFYkKegz7koHZRQfQuFmZfMbAVn3VKljx1Ahwvc6T/S9QJhQOI184um4s
4WzN766YfPj4GSW3VyPCeMRpSHHEQ+VyT21l9Db30CmKIlXKwC1ELGJi7GTRe3rKgAyxEAzno8Jv
522H8TUSc2cIaLPlVAr+IFzraGVQkUZb4Um/YCv5gpEhcxg1iMVTQSHagEGHUnSyJ7xwQqYzZ1ss
UVSFhDInsE1BA8Q6ZuVQSe7GxF4AZYuI/G5wecNw7H59fSVo3W9u/At4qVWV0HwRu5CCREbLpTXb
oSwNghjDK6U23X8yVzjFethWdn//cXJzgZEfRM9rOmPg1Lt7eYGyhyZV8++yqKyiNmRj/lS0ZIxU
Ci9gXMVadtJmfYvki1GeTXT3gCkwzQyJzGU1Om26Ab7CN98sJTsc6HMYughLcdCTrySIfkwTtWPC
qJ4cK4pCzkUk/3QkshH/nQ7cxdAztFExdjVQcDghwnmFCrz2jsvN2efXSV8BDygJ1UrR6fsQhV5/
1N5SBiSLsOIIJAaUQlgJfzyPExH8YXt9fnlwyTiLEAhtN2BixTlG8GPVYLuvx2oWQzRvL96ITkeV
YUBqrO6RP6pFr0w0bXeuuC2u6IGLUYY1SFNdgjJDYxtqq5Ho1eBABuDNZ01jDOExGoTl9n23J1zi
a5X2rPD6TGYLb9YCFCTC2yWhsXCPX+zGxw5UDMfi5O65WkcZdcrLyF4j6Rc7nFeOuQLs8Exla91s
vpgD27usYhEL18dQVqIhebraVYi2ActgpcDKCEp2x86sfir/cbo6O3rpGe0BpwEqVhTg9vLWpnOV
WN1dqqG0s6liY2MUUx2yYgwJhXGDteuA11R6acOTTnFCmQ1S42P8f2zmuARc3UXrV6huu6Ma+ImT
nEUB2DGOvr4pbmfZWAPnifBvm7PoGFY0spbbKKDvnSYwHGrzvwW3CjVQLEjBu0zQMftLkGZsQy/8
9Ggt+9r3QrT72Zu8M1PvXCRq8za3LOz94FsCUNTFbWpvunHQCOX0IuqBFIPeImpbZ/EvJr1yLA3T
7KN5md8a6hCBur9IxgRU3IaWCQp4MqjPymPRgKgOkYxuEt403o3VHPNM6lhpd6Sq2rbQSaaiv0SP
tPoWh9ToHiiOi15z6S8t5hDCl9NXTo0OvdhUXR6r1kzGZ0fo94C2b1qQa+dHrQscPfAYqxxBuMif
CIb87D9TnNMks9HFxsX4a/LTTZgvZ6cSuu0i/dyup8xPYFPUgXUX9/d2yAmelW60et5cnuxvC/cW
t1xYBLFNO+pKE9p5gqsq96lLRP7ycIL3SCzJnM6P/8u1ONcSG1Q9hSQiAApsOt/FqCS56tk5e3XS
gStxbj7vP5qTxHR4rDh0rqKjTWI8mj/UUWpFChGDEGm/w8hPsxhAP/g2mQ68ZwC5lbDlBgeoLs+M
0O16V0dNTY77gWB2fQbKDTAWexwI6ueRySq7BlZG0711JCnU1uRBzpSdQyplF56Fk/yE4E4F7dtV
5xxT+fqbh91WqiRG1KYBp33qHfvWtb6nJ728XXYwd5E3mq8DsHQIEWUnFDf4zGkixSDkqsDGwd63
G+1Vfxv2JM74svatwU5Je61J0KMK126RCcqvHRE2a8zYA50JQavHzaQOuOhdv5+Ko9VvdzL/xpbX
2hPhVoi5oR14xAHM7Z6G3glOIxEY4Rtt91Q8CtJBBaaEQIRVWhPH3qgaWyEeJVZxXxZ6Ukt7wmar
VjGVELFYwbZn+MrlgfHiEYelbME6C5kf5QLA43hTxYuR56944s3Vv0qAN+wmMir2obbWjHzDElSb
UyfM7y1q0YcCw62Sv214F4LoDH5eEamsLE/gQQBX2z1doJnhlXKiHL0P0dgNBGOtkjtlgf8sZsGE
mTa1d9OA41vAPeNDIBf4QkVKb5dwctLZzvVNmCwVXf8W5CWEM7DkkIQp883EGvrQeMVWc0gn8K25
wKrfbdCzHjWK670Qelfs1GbzGI4dqZEgD4qQDKAAgYZkW/0VJ2uhk2lWQ84lvRrzKn58Dnrdg2zn
tMK9WOTI/4iSSThPEG/uxI4k8D9Ipk2WEBEEMojMuFz8qi6R0shVSvG9G1fwAz/gSiaCmIg8mMZj
MGMgog90pVfMg6d7DojiVDCW9AufECznvDR1idJ32yEqGQsrANxDfpxGeFbmm3XEscRUk1gR5UjV
LtdUdxx0bbClarw8TrUAZqSLNlfOeiGvNxxy07D4dyIXz1sirwn72FQEym+w8KGEcs4GUnBPSq6j
tV+u+x2Qw23D9ilVUAbWN/CJCfzLmpHGpVHXmLkvCo0zOT56dJNkoPptNssCuilO33VHIAe3uGxi
Z1jmCGQ/9CnSGkONzrpXpwzNi+A6OUpYK4hxgY/485BHtmf7EXd9h6OyUuCYJPlDuYg+gZvE/jS+
zYXeBRLRc+wTmVnBmpfSkd6Ktf7/GuyHcQdR7QGzhymCtII8a4txbYy6NWYELCP+698BzvCikJ79
S+5+K6ee6DGB3F9SIGs9qp4w9xdrSLO/Qs78H0HADnFjxRViM3gQtMBJqDSNfJWjtFQmM6ZyYi3m
OzOP3hxQuzQ1vGVobNOJqqZ/7ru05X1LKjjZIptCDaQ00fIxHam8W1OPwqaaK+rdriWNW9h8Mfkh
Qaq5qjs6uk1J7KOQVHRVnYpkgBbHmEkNx3MY2XgYSrTG91VzQ0wvzKTV+TQ4k22cZ+lx9Dpc2too
AFUeyoVtFYELet6nZGtUSt3P2c86TDUaQp1khu/SCQ9RoKVYLkHEpmUZhfmtmV6YiZqFPUit+4rh
2Q40ejHGi+OLC+6nqwt4aEbppKnT5XJuE0p/B1zPb50iWCfgiChcEgTFB/NrYml3bAlXgeWl5QE+
IAhyYz66O4oXwf5Hdtcx3NcZTye9kVKigUfN5gRc3t6RotFcdNDMnNaerUAMYDlW/zktGCWTrPwN
qXKHx7x+MSrIjHIopWi9GG789ODnzzZBMERLfBr2g1A1A1si/iuZ2AkROF1TRKJ81FRtRvobCnVO
yoCXWPFN+fS8m9htUPmaWDn+mFNUFpSPmkTdW7sYPMF7+MvGjeIzWAIUNVghA2LJqxEViUSKK5t5
Q5ZJHDZ2VAITfY/GYN+ZAU5QJ/E/HkoUVKYWhXHTZpildarHGJDWwrtnUcnShvxwOz4j36/Da/WS
o+5J84/RgUw/SVK6UgWNaIpIjgdic18kXW3WpAVPuFLtm8T0kARNJrYC/10ejfRDV3rDbWNWOcXm
ReCWzGOTtzFxvQaaUk/UmxUw0Z6UWqtGtXXFVoPjHBdkMSrCjAzeTffageD8ZM8aylmgbinrA2+l
RN/y1E+TLznSib4xpar/BmnB3L/FaQ2EwZYqURagKQmUFic2X2pLdfHQcqqQSF0NqdhTIqllyyFb
KDj1YNV7bo8Qa+dRiYGUOpvseMbbtpb05yYGv9TP82d9JTm/Ge9apFnzB1Bnvx5hhuSd5peWgVSF
35D0bHrQmAeBcGARb46oMJ6a7Bp+BLCoFA8GS182VQChBRBn50Zerp49kVE9LDplo3NpAmscZEtU
LKZWAuY08h+NkHswOAdhln9QKz9GOvvUE1Pigc/NqjwZWMw5wXIC7N3Pn9nx0DtpDhxu7VuCG+xU
hJJXOOIO8NvrKRwcx2Nl9WSbC5s2EEHS2oDjc2ir49W1Sc3xLo6Vla+K5aP3ZaBi87zqA5gSKfXQ
x5Sq9PxDP9s4p05heT8nXKCpZiPJ54Sifowi3NT7sUldEYeXuHnDjjV6+91IkxlhEOXCEh+iAx5M
9E1TI34kbLLYtDWWFl7GZLQ+iMpeitPn+p8TiU06f+k55xS3KdB7WHFgqiewccisnqaZnhp5n7wx
+aSlls1McSJpoNo4l03lJ9rK015xqPJM8DsK5qYEEK+YM2DcSyV13UMEcJxEltbBPDqcyrhxjQh0
QYX4QuNcRtPE7eT8L6VcljIjMeptbPez70dRnJJVPS+Ph9s/L7fEb+VAbTCZaTpE9Myl69m6OGxL
qjQvYLxC5foMG5kbp3KDZ7uvLzWr2TlWoPEk3vNHzPhHhDHbF7GLGajAMOH3YNpMZEwC0YRWEyLN
vML7eL/a1h3ufbsa+iE+u9SxR11aKsznwzH72n98/gTeuHN6X0WnuT+/55LAsiKVSr81evwKhr0d
MGjhMkC9jXL3JRVZu8oLV3bQ7rS2Ap2N79U17amL7a1m/z7gAhAHNrchjgU/PRmg2x6wFd+uzQef
NHL5/J0wnYuFm1IuFqXhu3MIY0ZLIzpV3O3rKFK+5MJPhHI18/GMnvHdDKaVh4Q/UA/DUxwuzNaX
LodQIP/Gkbovn6Xa80oTi77wfy8dQKEY4g8x4jU/Z8m+6m6xzzbt492wRqFX9gUeKWbsxl6mQcgD
G6OhSrq+jvfsrZBvobenFUPeSez7GYN9l+Ka9UXtSn4PQR5IVt5wk4S310Nf8LAC8ykwbb9ADEBX
Kz5bU2uoqNbQwL98YN1CTI6VQnj97wQ+3F6cOw6Jus78am6LCZWgWUo23OI43xP5JCLxsXAWUEC+
wkSTOvZWUiiw0Nv3OSXVRMdmc1ODu7IzgyRuZuXHGzzXdG+Uqz6eCh0TbCwewMtPsgX8B8xl1n9x
78qGwHMKGCHs4jXELwHNFYDkOCMn0s2MEo0le9pDtgcuLySwKdKERE5U+Ronn5vKMu1PzWIYILJR
env6sPMFTirStpuFYTY2hF/HpRzEbDZqyPvldJDA1uNomUhFXeF1fHDaUZH7/oRbrT+6zvoH2aYD
N5ANB1fn7IHMd1fRJNJBIMSGcv0VHsRr1UbUGgTVoPzorJXfTe0hClBsq8llay9dqWHFqwX8s9J+
BIrQHrM1tHI1HsHU2+u9rczvtHuj4NMRexbx8CGGXA+lslG6xNPny9hGhU6TyI0WIKpWHUwNw0Rh
VT/mdk9gPnJu0vb3TLVh3x8RMSgt+pbXML+cmzjo5I7gRcg53yCNti6B5Z0ksm5HkbcegBwOkKoa
/YEVlLPvACMSnzsADBk1hLipYiNkmFKV2MQkc1O/ClJT6/dIkrz1iKm6qDIHFtttOT8hUe4rs5GT
tYbFMnsUr+mUAhhD4kkTHdxVWJhYKN3LbZ4Zj20scXn2FZM1OtIxi84mQLm6toDafHgAIn+bRzTT
q6cZ16cEkbXzdGTuEw9+3Okl2B+2eSH+zp42rU0IaBEzbIc0Xx2HFiRxog05ItfarbEawqFGuXRB
g2vPlqzPwLFscRFs0My7IovHvb3eKo5YfxFBjsudeA5qVyQONEw4azrffFtMGjiE19tomOHqHeV6
JhihfsFctzW8HoKgZKYOTGPE3KyIo17lWn/xhx07Ka5dOWrjDjbGToj7oqF2LrvAydzRmlJd8Q+f
UAHcyjx8HdEwi4oU7x37i835fVpf7eGiRfbiKAgtvDTx8wvNb2l8s/d5MJrQT7XqHtjUC9Aplkzj
sF8X0Jq/VMwfPWKtwBx+abSDWOm1H/5VQLk/ytdzZe3tLQ+bS2T7Pfhq7lIpbdsHcGe5eqUt+ejA
PE9kefs52NMfO4+ox7WRBeJhplJg2+RrkBtpiV4k/nz1AFt7H1S4Ql2MFuaxMecpmDpQfsOiBD1k
M7PPzlwpmXb0t102Yuw1sf95i84Ykq8vZ5VhliAnrYpcaKb/R7LxD/AbjMv7U522ZHq9Un6mFQfL
e1sYDlEh0djGqLp5zHi3UGIrg6zrsDGwEQ8Tf/Yrgf40KHv9x5VsA+NbXcpxx2BWk7O+ImDsJjiL
4tiPIybNgy5VSY9C6/ChdbySYP2csdKmlTkvUIimt1tUw7mIktHbqoPQV0JK9DWxrcy/s/jr3a7y
FwEoURuV8kD5gOuRnsQJ/x+vMFbTVTKRvCkH6WTkVSngKD8P2ZqlvcVUjZuu5R5aHq8dFLnp54Tq
FL0Qqx2qas5OkHzOiFt2EalpG/kpXlzeHR6L/TmeuH9NqV8mIRyaUn5bq94P6+EMsrn3iTLqtHnK
OlRjAxKpE6RmMOsOFFfLOdVoyVMvHByAnp3q80zmXEy56s81YkRCu0MYPTro1lrQeEPaIoL0VwzX
jq1YS1qt4zf9PP++beulqKhXlEOAwtCmp2zcd0iWXgfuvADOq330v//+WnPutwFdI/uH4nXCJJZ3
rfH/jocTmeOesDQuroA9VZv48+5NVpFurdlpx9Y2+ZQ5XxwXVAJBDGTguMCCcnpQ10RujIQNRLFp
+8aCzd070hXBC9RgGYNQMFuboQ9+E5FC+sFs20jG190cr8xxu/R8TC+jvihVIgcq36uL2eb3A1jj
fA68AsL3CPGgJRuOiLnpy5jRHTqVFrj4onxSjS5mkFQvzLQVGPYxAovp4o3hgFDXcOfGWVj00tmi
5HlgAdjxyeW0Xf3jtPTYCts5h+sDHLv1zkdWNQC+HWdlKX0ObV59uCMW5zeDy+HuSNhQFi9adQob
Om1LY5Pdz5hsgE6ijE7eYNodWY9NOWJj1NA1KlrCQr/lOoAL4OctsD2oozzM7hd9LcrbaDIoSnFI
4b/dfga/pzeAsZ6d8Fssm6ivzTgeohETwNfixVQxR+9smT9cv5STJN+GxOvigQCY5kNdkfwJvyHU
Mf27brlloqClZH6fXc25YX/RSQ0GA1v0epRzNarAS2Kjzmc31ZfdXDH5L4g3r0GWm3Jer0eQKDTo
8HDaSlI7+Om3+zI9sc1vea7Fc5PKkmS8I8PQnAhFxYP+Xxr/ZTQ/XOC1VSiAHlnkXgJbbYbREeNn
SlpGbcRc604FLKCCZ/+i/T9ifAZovE/QCKFsaLz5W70BE/Dv35Sn250SY0rzPxUhkumOYwKzrtGZ
GYQZGgwsJuhyAKRp+ePRXMKauEimR3xsFqJyZYxBDSgS9xKjIlv345jr1n6jiCesoNr+y9DUuJNj
6uYkwrGvRelfYuZdvX2SkTAYdQC1ueA2oi+21olprrtmkgzrh/J/7eyqgW4RbGkSX0p3QNpf6aPI
LTTRD7rWR60AaBoFjQdqSS3aPE305A8IiK5sGC5uf/VTHA03/lRGYSPZEK4T9Njds9h9OZzIux/+
OlSrkSpPpywKnbOyqQJyLB5n/v2pF/ONKTpITmDfxhvuhJjq2mkpTtJSI7hLFvabahi4rYfUxlYR
irdI4p6NJ0sgbHgAYs8OmctL9HbTOKpAywbgtQeRFz7Kf+EpYq4LOsi7NknyrNBKO2A6fYC9t5wL
BZRS9JeIf12ubBolS6loaJrtyVbdFn6iaC239AHeL0iqPYCerIapdo7oFjZkoKAtaQ0JzxeKYUq9
2xbQIeO97TGSkU2gsWTWkyWNj9I54/7pA0B9+OrV23WFf/sjlDteBf7ZjDVwVG34GyyFGdt33ee0
8MKSCkPgAFowTHE+QNwiQMj/PtA9wPqrFekdvltr/BhIRcPD2AHXb9v+vQh+fvY6rs+BQaPf2pNh
v1vk97XVIjvGDqtjqCs9zUFiLAFh0fZOWeJK3ZoPcaY6Ks2Wbiv8diS4bY0gh50FfvyYp7zSR0Ck
jwW/sq4itZK9ZnSt/oHd/PoRgSaj0k/x3KAIFCsd+EXKCGnAkqk2lHe8r+WCL2kPrTZWfvFBwrSX
pomtH+Jexiv27kL3K/iow0OOFIFbsvyJJhzOHCp2YR0BuxuEwcyIwkaWPx8Vldu24kHsZ++fCYSV
sVlf5FAlgJZChg2ug5Bseqt+Bb5SwoyB3Qonmqu+gAjbR6E5htH4l6RGu5fvDAOwuDg1nj7KZeB1
KbjJbw3dza9xofo8pQPbXcxwQKyXKhv+moG1x+mWyzADDFLwGxjzlc2juLa2ePmpIXRIcmuWiCEa
Iy/WITzcSbutnVD1Oaq+DzjOpN3982k32iheI5uY8L+gVfBlyj4gFp0mBSFQLZyOA/BQmXibBVJ1
P2pB6UIMrbSR7t6jBpfFDxACym4DY8KFcPp7i0zMfyRTn37aMwCw4xnZ2Oi9Q5pFrzQ3XZdzZpXH
LqisTfpqGWHwibcl3nzLzYOtdk+kl/1isujja+WlxPVgxrae7QEcFjYSTOBVQDqLXxfVd7mvGIlK
PE7LUy+nwti1u9Bp7TaEqxk/d8bhy02HmOfkMVP/dYtho7rSs6dDDtzn7L/Es/VybeW45H+0r3XW
YUgjy9pNp3ddRvmSLP8OcqhcKVrJnSaMKfsDPTgGKzx7crZJK41dxi7T1MriiKY0WAEyxBV9K8X2
CY7HkqtZAeFOpIYsPxHqR2UpPRST4zMRDcT0SA9q0NT3oeoOzQIh/kjJKIc1hTGH7ycs+sxA+cf/
ql1Yo1Lp7p+yrV5VfystJMfC+gKAvRe8DVnxt3tz9BU7dXKjCw9UMI83+7bwjsb0VfQYykx7Rb1z
3rn0MXDdUcfDI7Fl23RcGc7gfS+ypUctRS82GeMWl6n6B3sKbqRMyI8LL5p67n70G3h++e1YGFDU
/EwMk9utYDN3T3swdqp+nwHvTs1eiYR06toEyXTSoRiEH+lGZW3KxKjssNxWEbIMHo7vS0Zi3SFV
Rl9bf3j+4P8hTtfLv9hh3kwxkLgdOQ0daLpjMOSbWgVdpnMgJRuhQzgMJc3nETOu8wh209dM71gZ
mPBaaK/z8jVCCj5zHnt6D66vjS3KKw6BY1JoveNvr734LV12NTQ59YQPyfM5XebJb9BE78H26c2y
bganeh2abdwkl+aXzdLiNQ8u2eEtXNT7U0l8A/QG6l9SixTSe8+N2Z5PAmy6iyHH9LB8KrG3FAuf
mfdcVrg1A7zKluVq/FbInlivg2we9Tkv/+0At9Fxri/FYrW1iP1CrpnCfQMz4uKhP1mm4nKFIx6t
oVUbrUW82QaguAPFYR1rd1g6Tdqbt7an1RcfERpDPjvV4zWsDIN/sYt+LiYhR/RXP4EfAVayzVSp
2Ma5Ydr9H33YgDd9vnzVl8+jj0qPCsgH2Zq/dIxhYoLjPGh72B6kPHTFcYP/LpEwpiQVzgxA1WRU
Rcdc1Y2Uadl9OIiMwslKBHDgbfNmv0KDmG/pIX4F3NoOr5QpoK7RqNEHM5QSibEm6SodvbpGnfVZ
XcVHjBzjwcmAR4dp7QnPL447Muiw48ikF/K8iZW5/40FVLFn05fUqn7b8zxLAcGvFQrWt8Sxsa2I
FU9OiPv99lxyYsPcxmAOx/ftiQBxWM1XWm/bXvrrMyNjuNwBuXtmxbesDC9A1eOfdzpglqoC9gqE
oN3MyGVedh/oZe1NCZWXMlHsu1H+35txn/b1V7NszeXdFKozFNnvd4QQA3e+nw4YMFGipsBW97P2
wrnpMbyHQCx8zBOfY2zoRJDALRmf8Ytdu5IEMMSUMX/3hi8HZZV8zFxyp0l+6vmDDZaG0HkdiW4W
QFLJwZYDXEh/f4OIWysA0VK/OL8HvEsx9mz5YeYDO9EeVgqJl/408KPSvwEQrFMGutYBwtlFXKe0
6pS8NQgTY7/l0T7MY4TN6SzweGO7FxVeT9iK4dRC+LneAe+oM1UM2YHqLvYHzGfRVwyZOtQSbgUC
GJKLhZJS0RUHK1vQjxydYmVBKhIlOL246piwSYPIiMkRJ25E3VeYRZna4lqUSuBA+2c42QFVpV6E
3VgoNIOzRtjBua3qkfGfV+sylLTrcPgRaEot08CxqYVbr50HkvomyyzEKGgY7ZBdM+xm0Nj9pZrW
4d2fieLldbt0f5p+RNgiXDZhA/07gYlLCjKY6mwddt+DcAFRwQ1y7dB+qB3+Ip7g5SmVfcWFgvV5
r4p0MztsebxGT6bLLEX5icr7s0jP6MgjjqnbxuK1Qkk5nhdA7P316yliiriPnBPaech5QOOhTiMr
786GZ0Jr5zqXOBw3AbNgVGozmk9DRk6wk6N3uHXTTFWjWCqlP6zkPvC+wpZA+rMfqxumeGWuD1P5
aePCBWoWXIRdSC3eBZURCVQ0NJQOL6fU0HyJ6B7BWqsG6VYsDbiOxyiPpyQwcR71YlGzFEuG0Py7
EyhImMGR20fReHDgHzT3FKiYUXdIJMR2/BKg64q/201twAVCgIMoNpCb1SDwPLZZlhE0biX9Mp3j
wf+ez/nIfUjS+hoi8Dlb7qmdM1vSnNGL0Co/zi2FlDBTKCZNmY+H5cwabkfLwIofqt9ba1XoU7lO
+iOYN59QqMBW84dTlbGaD8w1YiPpdw+1bBhrDpnxvPd/vkzSQdrzAKjws1/xiJM82mzqmcI+8eRY
N59jyi4VkvMdYQVZyjZFD9w6S9H5ezR+yLU1tbCYylglUvkMrVPecv3rdbLmvpcOe3qhevDygbyn
Ijih4NjzSuB28hGJJJ9aGQhxeyubq/yXvGqvDUNsvkL0+oEBTWKLemdleaDDzClfnrdl/bktTygl
kv/7EuUbXQeeMDnD08U6QdqhST/1B61GzmjTfmYgmej1zgq9f40IMe0yRI4h955SULsQ2b8W15EX
Wr4+urcROrNF03K9wTVKgA66ClHRZPHD5ZlRph7GGaAQF3g8CpNYJPJ8ZZcqzSwtRLLKwXO86z8Q
EvNZT674obSrIUNZA3FmCV0pWw6AtV74ie5tNfvJtWLu1ZjxMOXcKYVNmaCw++IsTxDZDtOV1xjy
ntvjS88yP6qEKWc96UtsJOOnJZp0CZH00cwKMAbn5xVCvgA+Qm94EwTKEUd+yQEPQOILM6QoovUJ
u3rhsgoeMgL1UVUVxKyztJQNbhvn2ERgue/1LJBCao8O90tYmScl6E2ULXsOa2uc//RxidYQl+GD
rlNJbzjFtyZX7mp5+Hsd2a1WeJCFnzRXgYYaqub46rySS7R2pPmFnSeZWBrVquxMcJHIN52/2o8G
U0G5C/WFaWqJ04nqzeVTAm/0/iTYb+P9kDDPXWvFKgvRs/usZuYAhHFGYK+IjLP40ZFKDe4iBP4g
opE7k7h5YdzCJ+JoKqM4jhtCVav4pfcnBj96DPLdGFDXc/mSQBDXIXnq4VJ1NF1jBHIuwrX12IVG
7pyM9EpAeOeWEl96u+DEEnwlH4HPJBD1Wvv/AzWq/mCjREjn2uk4znopVTmkJ+rKUePhcq9CSnMJ
MuuNPEmtZ5EmwCw1c8r8HSGJ3ZhiC/a76tdVsm+Z2vUQyaF5bp1ThX3NNskskjrwOeuvfQ/YEI8e
QVsYrU66gYoEjhQvNQey/ZbVQC6dkx7GNTw6DC7vUtuLawSGZ5QfunyTxMe/Lk3tgzyl15uNZ56o
32Tf4BzK8jVkA5Xmp1qNAHmlJoZ/xkGrUHDXPqA9BUuNoRMNDXC5qOdS5u0zttqFHtbVVdCdsBgT
f7WA7BTHLCqJHxKrDp75uDD11g2h8bEACos2umdYbR+8tIXv4hgQaPDTzJB9jae3ZdjQ/UuBWsQA
Yys7h3yaoZbRaZaPfurDKtA81UjXguCrwEYPaKXjLad/zWd+EXay7xV9K6tK7loT0Gp29kjdVcmB
NtdZZf5TXZKQRPcZ5IqXTHr+cKK25Vhb17DmKjDKNFKncg4L3AxYnkHqXkhx5PzKIVZhdmAGiLAp
VD1XG7m5CEcWPML5YbCY5wL1BjyKeuN1zmOJPXopTcnPwApo8BU2d6o+2qLep8lka+FO/ZR+44TW
CHxbIzs0qRt4/1IHlL6aS5gbqFX3cEp1SUoybwlyXZ/6kXN3HhOUoRoRPOiPhR1xkIFCd7axWzEo
vEdpMFhODX1XWXGPbpVgb1zzrom9YgCwCLEu5Akr653iAovlk0Qfs0/AdiRcMpKpBUZPHhzQnhG4
aUzzjCic5qyfhUQbA/27lS48yhDsS+1f6KqZ7Vyyd8vh//bmLgEwkOgsXi9XmBbU6STA8mgZn/uQ
/8oU7/Jvr07k3ge1eHoUnSKaw/gSqHgd47T7XzMzkWuzktQY7TxqvGwbLrvw9HVKaPrEO8ECxLcV
mXal4nxrfjC3OKxlOeQJkc5330mUZjyuAJPFiMNjOgso0bw6ZzsYwZKJqEaP7bEjDlf6YJDzbQqR
hNZxPCGd4rS5+69lmcadj0sAHKPqccFkCPUsFaclEPYlEuDhEvSJRYlweSimGllFFyfUQ8pd19ho
+R9ClMpemKC9S4BZ0Q4Zct/RDLcvJySJXWWczcSG8KVl/MJuHH7gW81+RVWZCn45BSq53r3Dm0ue
+mzsCXJdHO/QD0UtboJ0e5f+8Y8Q3NMp0bX+p77QIQSmDQZbPv/XGT8TUzH1EyXW7veVfixSTLPP
JIBlVVpXPuhCEnIMyHJJ+04ZfCwemWuEw/UMYvFm+kdrLo2G0U3+UquYkg9l38UxWHR2ufdl2t5I
gRSdbfK8cJcAWjIp5pXY3y93gnmFL1zaixpgcRi29KCH5ymgUSz4Fsye8R448SlWfaSv81z6N91m
He3YO5euEUPyeq4V49rPpZY7J6iI/ZExbLfqgcrcGTj8io4n1w8O85IX8KapFhZ1sIXcYoV0X6eg
Ww1tvjc6km46CucgWtrc+mYKzjwL9Kehv24WAk+20+w/p7vwzvuKMGu921XiJt7c14DsEFiUMk+/
F1XF/T5Cgd5BCFe3OBMMJq+mDOSvO9Vx2rLpE+HVjrH69t6JLdCoYmhutpdj8FioQopSMIU24xPf
goUk2AuowbmLShKoFpvDlMxciMRxfYQYIkduwofzCRZL2zVxFbTMOruu//64qTld7jvXweyjGoV9
EdDevrursAW6bNemeZiMRqgfCvJ6CjwppgAFisrCGyviS7ezjP6cpehtTDE7h8zE9/FZx8UvGXeF
S8OLxOw99/3t12qfhAcj/6hLDMQBNDl2GDf3rMKS1Shosj4DLAhiMMXkRoxSO0g21hEaj22uUYjw
42WPcFJEwU39aE+QGWCl/cFoMLHo6w+ju6kdAzbzE1xJxTnZVsb1c7JKpY4trOzsG9oMzAt0hE/P
0mLuHf62EFw7SXFvAnVM7Ii81kiup+3JRlclguw3ht6pdCw1pl3ru4MPBffIYpn4jatqitVDrev5
zOwI1oaYxrGyiil9sOgxDNmMuI7iZkyXU1cqiiM3TVh2zhyQhIEFCbqPSitbJd2BaRy/Ua97DOqU
1/j1GMYXZV+MoZtU1iD13wfEzfTrNCPvB7kjIiBXr501vk10oU5GPjWlevsuhMo+3shWyPH4QtkI
XhlxROKfqnxf+Y7Oiz/yqfAG84wvlBW+eEPrVSDos9W3uaqw9wtXehJnUq5KBuK7aQGLJNH3ZRG/
LfY9IiIzalK/vDBM2x93mi8S4SKkhe7CdtMZNkMVpHBBvahmgU6AKdiM885OkwJljiCUWqOjiUOT
D0uSd4v1zEWVGkFFNWU1D6C0E4RrHTXGG9FakZdvbDwrUGJ/fN1MJuY58Gva7PoKyj8ZdlRg5vr+
vlnkp88jJLuQo8hDC21SddTTU063Ljoe2XtPwYyhgeE2RZ1s4NsKUyBsTgdltT6JuzbduYrNM8Jh
fvh4cpipLA3Hf16TEIVIIfRnafLOCrlW9nDGmFL0eCTkC8aeQh/7KlltuH/EJ/frqqqtlu7b/uzW
U2kY76bgYXjoKPBAw0t8jfXCUavX8bHXNr9M2brIYVSpJ8kjEVI7ahzwHEYs2HHrEb9XYnhMzBNr
UBXeEN3WrY5OoiHUNbugZ2zpZeMGuyLWimrcO9nre7tEfLijnk9p9lOPJzvrE9YccT60HtF7K7V3
waX7ks2+8mhVs/ICGHMH8CiHXrUo4OgXQYQ2L0S63TUrNgeH276JWZVo7xtYKfkdwEaPwa2FYsrj
fEkQanKy4D3qrQgKdPPlJAFuMjMHY/HCgqigMzV2YQpigW3BW0880XwS1yys2OlxD3s716A6FAWg
PrarZFLq9rwW6q8lOD5eXED82JW1y4Ojm1VE/lm0DgvQ5/sAv5oni8bT/aaLvIIPVzpaP42M8/si
CHLomnrodAa60k6fvrTcJYJ+VSOYLz5hm1M/u276yU37wmpLMJi75uClD29QeZPN9TYPFwlNXvp3
Y+3YNlEUjIsOZ8fbAlG9agvbceLkCSMRpc6btEKJ6VShMZttJC+IBJl4X5d7fgAxX9Lof2RtaWTa
s37/33VF/7OYXkG+BN+m1ARHpdXSLJdlNJ3bCHJJDpwCq1Nms+wLdJHeV8dZmYuBUTEJ4DGOGhw/
RfgPta+ByL2zfAtYlzKRcIqctYPohPJmxbX+61UwvYmwU/7cl71rKIzlsTh7OtQeogsT16QlQhgD
1f7HNcUIamXr2vbBUz+LJZcBjMRtyTAw8VdMcuaywHYzwrtq7+YBqSG0V7RQQacvv3M/U+ZEnBsJ
1S46q8ExbjoHJ+PfqF62B/O9IT35gRp0BWRA85y0Ue6Wbyxv2B1HvCBUmSjrMRXbySPM7zNHnkYR
iIzKb4lol7ZgBrAfU7XinpuW4uZypun8iO6HEykZ7fCPxz0v1ikvoCveI+Fsl7CKO5Dj/4J9f2zY
9A7cCs6qleben3dpC30xodhyNKGJHZIiThI8CU0H8cHasSCnoaNAE40ZGsS6TwowYMxeEZbNmR02
rYrUZMCdJEhTjB1mbb1L3JL7IcygmmRQM7uBfzzAoGAHOECHivVo91al25c6TYwiXVvuw7GNRjF/
uFbkGPRiNM/48TLgHf0MMqTni0OcP/bKbiPYPgnqgjINLe3BbccX5hCHV72gTE/VTAieLUImitWS
Ma4g6bqr/QbispHrTaENMFLVr6WKq6HBWNPb0Sz9rnsai3hvdkFmXAI1wU7ZDHMWCGo5icrAIVCo
RjN3+9VuxkOBk4ovmNpYvcRZBUzcnF8JM6li/8yHDJ6zC6+BSV3HIpwW5FCyYHM19TyBqwC5UQrW
PTedcaAdVvu16ibfWJ91vBLfQ5Txwop16HHeB58Z6ai4zDSTZu0Zr6UvmiM/OS76bE9oVT6f+TB/
zXQsY6UloNk1X78PVSF1+ZYiiIN97jgTUiAXl5JrWjPBOqNnBCXstUYh3cRSuNW6mDtp8wwbPutQ
tnudhD1JIQyKIsxv1Dmw7rt90RdnS2U2/IC43JA97Vn1PNNU6f32Uj+sCefbsJ+Ffk0xvP8nsDOT
rxqqNavTgBZ6Vf9MTlCl2wTKQf2Vk/sdt8fNEDDzbNP1sau7ifMYUbl4/6EiGQhf4wDGC6YNz7EU
8/8Rh1vYe7XY6jF6wZkU0Ib48rC97H6D6olpg3QuxIcOXKLLwoTizNi9k3eJgqWBOFn/RVSXZYxl
jxfevh2l86AdWmcdlGRvm9Pm/fBTo42huCjSSoQ0cYzRZFQayYrTZl0WKfPij7k6bCXEWBoZt7Ft
66QZd/Uq0gMqoSaZSLeFdXKhEjbvO5tViymFQBNkXs1+ZuZcmqwSbpUuQdCam6Ukgb4SWgoANJDF
xpGLL19jfKPXTNBNNZgnGVtq8fqJP2vXFAwxbNC47Uln0222Q0D4He20CHfP271Eh9mGGXQdF0Af
jl26OOVdczkuRrw91q/KgeEH65PL2OtXFRbv5zsv2U55ylT6BCn57861qMjChUz8O+1BZEGhkMI+
KIfWWXYw9B/IoNghJfD4HZa0smM2qMCZYXb6OzeN8j9wW1My0EYK+/xWPHyUMACSSyQnfxmdRNrl
dAasIx8Di9nXEj204gJBh5mQNx6ZMPvGx0O8Kk6UHYdObBJaTDDHjcz9FOH+l6yHx+5K8ui6h1ku
/rIJgcnViWRITyxaJW2G8q0Sdkv6rzBRJNfktVsE+MT3wAHhzRome5b2XyAII8kf4fuq/7x+XNf3
zGMIK+9LKFU5tMehS+yQuODt/QNzgu0V/vx6HGA8lox7dZPR7e1cce5P/nfSlaD42rDeIntLy69r
18OZj1PzuAU7QTfEEF4YvjrJXqEAtUETDXXfrXL5Y2wV7O4PdNUtrBsIByQD6O//iiOU36+JXlQc
kSqNKl4UvAXODN0YXLGSVW6gClX5loUknKwDTbKCB/UiOYITpTeiuM+bsbVnWMYv4lu5jUPT1Yqf
I99kpgHPU/89JmJdzvIQQKWNJLWcjonG4JQiJ1IiJN3Bc0tWAAYZZNWWZotZ6v4qVxdIuPX6Bs+B
uo2GjYjY0kSkXjeT43bHzvUOuEyXTauxl49vgPniZUinUnhpHWnN0vs3HJoqZM+v7Q3Gn0+DJfMS
g3GYfAebMFY18fFn42J9c47V5S7dpHjhW9dRMgXHG6mLBObi8WJpOKph9fLgs0NDN4nF68v8TJmZ
JjFQt7YVoaHajnsCKfBdMpyNlIIMYz0ke97uL2QBOm/HChg/LHZjRwJF9K7fPQI4Uw/ImDX0ndaM
KI1J44/UX8vaeOFn48A1E0P0HRQtJgutddp4uYo3PIh7xY+be24lWZ6tLWKG2ukBZiuoj4RzATG0
NELZBpzvuhF2fIJzdz1DXdj6lKB1B0zpXJEwnSbVwn30QjlZQyo2kY3t4WDYqk5mesF0T4w2wzFw
9jNlk+pgU0qaakapFOEaQBIcGfmps93qZ9eTGSXr04AqmAPaBJJRlAhrpSabbRJPazZsWJsgtjfP
KCBMEK9GGj80hIk0qJWbPdIwyiH/kXLwfAtblPJc0MJmQDBvQkevZQlJgLAjsQv1gzoPI6pj9HHv
6ss9gktOfZqsPUUz5tWWXNBdZHgKZvowV/RgviQoIMvbepenJVEQST69zqI3/DaJBGeBE5QKR1Au
ren7sCk1XwP5wnUIXfq5DcM6fXoTKYrgEA8V4VDGKKYZ+HFHzT44ih8V2vG/ZY/kFfwNuR0CrDNV
nG1VAJIE2gHyLr1744uMzRsQbpJl44htrCWmT91I3rCiVlZpj6fktITWOadW+KsB4YlG44/PFhih
I1g6uR0lux+6FoiONx1n5ChKZVVvIeQLXJ2XQXnkdBLu9BjSd0rW5cbr1sj1+7VueWvNo8dMUEG7
vjRJj8Ys/o/rQpmZPLiuT0HqG1edwqIiCabfvN7sOVUlOHS62aWMpNkKovRnOnSdKf0a8lOT0ZOk
vLfUuS1WHGj3TNWJuVsdgv4thRWBo8RZbFJU3OmDsa9/oa4DSstoEozJdptBQsifGG/AWksJnMFL
HxA86ZT9kttKi4blR8LUj26enHAlgXhvinFf764hWyER2UvWsrqI29YW4uMwjjZl9oV9LG9gkfZR
rt26ZCYmbPp1PM2M7fa0yMmWaAx9htZCW8YBSOsw4Rq8tuLlih8XPzT5i9f23V+V6QCBlmTFjQ/j
5KBc/8LS2tIW/+VJYle/7eaw2XRntRX9bJlfQmRQHpP2wL2bcQWXEb6CmjcJwE2CVrkj9g/QaPfK
bFjV9FKZ1wvyV77QWQ6iLZRztbiIlNlm1kzTiZWkwdpr3ZCMX8fz1KyDJEPLwxJ1x5XCqcYMXBzD
H0lqDusZyJz0beLi90migE7iFJBuHlHBpJGVAIdvPSu0TYhNM8LGEFEqTEwWSt4UzA4TzpIOzZUf
FrYNK4/BM6JvF61+5bev74Mnt3JnbPYT8bSK2hUkKXtDYQaiYAvi1e4rp3+jtGPj+A/+107Hlb9U
kXIt94nHcPOmzHPthiHhg1hC8SOfIXwO6G9I7cIT0xZeuM6Qr7AkS6fDscdouBUBF7TTXXF+JWBw
xaJJ0DVg5QrGzb1crwE1eHiOKTfqoKQiNnkTD4D2xqTuWrLQTJTjBQgFYaLlsSK9emW20AwcUc4Y
8iF9kf03Q3I1a0dDjdn+vmhP2wseenj5NPMPUQzxaMzgHk750cAVdbLEwsHYPP7P7Y75OUPASlHw
Hx0LDU04pkAomuMM13cD/xkKLXrasac7iSU7DpLHM9A9pg1BKIGRgJxYl6+HfUtxkMgAcznqKUft
sOI4rEdhL194xlQskVvZfFeAieMKcbFcPOeXHDBYL52tmSioto/jFBPFNP6Nhq96uQ1Pa47GxCm5
9SDep6QOFHEEjugLfqchyXIdzHujoO9COq3iCJuIHYG+4YeEZcTKWEmJMJ8z7566uoRkeCPqf+ZX
MqZY3RcKDNXoGGANZdXEVqrGBB9jmJ3pOo8LKSMptsh6S/8KVyYBFCvTmfrKGwcNaTDYoSuUIHJg
aMYlzUZeMXXa4hrmZ5NE/xFbFrNU4PkgebCxD5va1AXPGAHfTUguC9CARk0PHEmbiDC+g1gl/BD5
6oHJFEDvOVSfRwxpjdeuyBN+PZVy0/jlcLR5oRDda7WBOMp9HWrVRGpeKAWL5o8VGfRvPw3VRqKH
rgqjfEja9WcALLdVIHgNU2383opHvIbIPe5B9cMfw1GNSTxeMpM2H4WUNFjrwebaMKDDsEVa49gL
p7sMMeFwTASh2GdmHpKMxgbMYPhAHy6cnAYkec1W1PsNWp9QTLYoz8IHmtqt5mY10PITvwowjxQi
l+TjYMbJJgfj7Yty6kd9vuUhpCqKL9vX5vsunhpELm4CEuW2RWduBsyQ9BPUFS8xrTP2cOKWQqo1
7N1WZP9OPzWUHQcSQe+PCjCcLRgB8JPuGv5vrmbEmlvEUYlG0PKiXqbOlfqlU1E8f2hzS8BhB5Vf
5RFhjUrShGHplCm1bJ4fJhsquc5EnJdcGwwR1a860N7sSGW5ogsSoO4KE4sOKs/3VYqrmb34GEB0
lbA5drRLbKNGaK4D96oatz9+EcTMOVnT5cdVGO2N4JPtwGue5jFjvjHX0ZiQS3Nqx34l1Q02LztB
kRSs66OQRqqjezz+0bqxN7FiUoJdHGmiq+cNQXhn2cfyU5nUMv9LF1qHriDnSRLqDq9QNBtM5jZh
8L/B+q3tgDQDOV7mpJEpxuMJUJ9YM0J2Ev7RE7ydIutNt9tP4AQ5Y0957u8M3fguAbfgkhgQm2RO
ivFgtSsCoH+ApjWUT0keBnhCJ5cNuR7dKLahiAViQEKjtghhNbIsdNgfXkDsIYhzr8PQdfdhr7H+
DqygG+HmqKMcoxOjrXxJXNgdJhWIgaoNy48uMl38yDy5FtC63wkTuTCjBECnZeX1MSLSkQel6d8A
OrVHalDG0bNc4N+aJDUW6CkBCSGYiU4qm1fB0HaZrcR9bchZ4L6KD+UKoBBGTOX2M/MXnJOGhEEO
lW7zYZAzA6k9gEhnxpk96B0ualzS2MqsWDWwYe/dzXKZynXHg9YI+Ga5rRuwB9pXeTRttrS1p+MQ
DN4cx6KH7YDKXhnKc5xXFCZx80b2GI3DtF9Qw7umUTbsBwNnK3RQHTTLfv6/plHOzhJHXOHKvz/h
SHS6wtY8890xP9ND9m3CVIHGVk98aE9Fd5ExoZt+fXPkHBOpxQ/Eh0YSCKjH23lQ823vbCQBbI3O
ONgfqYpOivH+wl5FmfaQPxfsOFQzGnLr2q6frNO0IazwfzJJGTzvQ2X9D5ac1dReXB/8eep995zV
AZBwf48Ph/j4bNBGeLZTdCMi4d/6Gngq2Ol3KI9EXtEF/5LGTIrVyEs38T4LPxwX1LgVB2x6IxLU
OSIQkgADa7FmCOagGNPU/+kQh7wN81pWwUM3acIQax3ueUfTxeLxoDnP633orkFstx/fK7vTA//L
oTayf2xsZE1cC1AnDf+3fK8DqQEXhJWEUT9gwbgNxS8xpCq17HCbRRdYjIhSww/YJa5SpsdvDFYf
sq+1TOg/n43mjWJmnJ+yBsII1DVgT3dAHbr4RVj3xXEishE+4Xnj+gY6rLdmJbXnlgFsRESJ8sbB
83Mt2HGxPiv2vOqxhyddkzBl+iXrUlhVT8imNSRmDyV8fhui6b1fRqeHBCE9tVXiD3hZbafWzUG/
NtnL6HyL5fpHdoPIf9MKQ21YPVIIkSLgSd5B1IirTw2Ne3/T9F0U1qntL4QUS6RCez9KYjAupMO3
JfiQ2pMOQp8bmkBlART069SuKlXNnXaow4mYOh/EwC2x47mqK5SzynBhPPnIVc2Xi471IaM+3rkm
uyMbaPpHWDzUgwvUSBxqFDc13ZmkAFmMf/GfyRSNuP2WVXFmNpaF0o4Y6HLQhImX+00iErUgqNy+
HpGjKN9pmtDl2y9Q1iXMhCut0K3BNvxqLYeXC6/imPP7Hl7EhdQtJLq5dg3x8f7Ok59tBHm3+GP7
kfu6P/+ptT7YqyAxHlUuAGyyrUHTMZ0tRmFWl9066tfko/dxLOOuqXQ+S+rEiYGFAuLDoYXYJ0j/
NFqMjtuF9STWQI0Cj7Av+5IuBaQX2BOzvWxfBfPtJQrK8HO5MEBuWxC9JJoS8CXQ0gzwCjkQwIjU
qBPjHyrKWedKm4EN60idPVk4MugJH78q3icI7Iz/88Gdm207oosoDufzYJvcR86vu0M/zMfk8qpS
REUMujZK3+qVwcG8rF4pGATR8o5NP8OPHLfkUB7tX3plU/vQktMYwbkK4oVn4PhBTY8xYe2NLgmx
bJ/keZneBY3IQ4CkboQbMg94NwhXbPkBIMzIEp3kd/ULvso+miFU6REs/ahniOCFm+FMJQu/F83t
vmQxNiPYhhPand3HtUbduGx80YecRJ3yuASyeEFGLpSmyanvx0R/Qv7Z7F0kE87nmZd9xqZu7+0V
DSyQIBDTHa9ZreOCLKm2jPQ/OY8MlI0ltPcoyiaX4tL6jUjgVLG+2Ln3OCEf3gSxZBi6pdwXrurA
hMa4MYxtckM/tLknUHWocjlOjilaqKtrN3IIowwZ5Qks8IVHMdm1Ma4WmjADdch7TrrqQKi4/+OC
dnSRa0g8+kv8LgGcBSai1r2m6+b2Rx/xMpkQoOS09mYeQ39dbnKkwlGluXVgF5FnsikOGmYQSLvu
a0X7Yad2abbiqKQbV67HHUHUWKZpB7HBVtknbng0d4592X6G3uG32uQGjytpDpl+oerNEMFTcuZ3
+8y3oTKck9FAeZ/Y2S9WqFffyKJNLujbPrrrhtI5WEKpQNQAn4SBK8Qe3KTXJY1l9sB/O480y7I9
XR6eDRkeklmyjc1PASV/yH5FFpqbFsubxR+ltUvTQ3JxIxpPLXTWGpbGKtwtd/2NDgBADn9QvKWE
iQgTHQDUlQnbiHgxLHk/gtCXLYnhHLpA+tqtOD7FAVyPxktcBlcoeDXzjmUkx8yjRMGaDFrDmfXL
NcHB4Ol0PbnL/lQ8i76CDQUA3yQB7JMmCvSCRMaGx4Sx7QYgR9sXMLF/jI4/FsCypH2usThOqvsj
RPQkTR20GmwA84bSgQogjFNS5kuRRHP5t5Xj7mVsukG1/3J/satbJvauDTMm444VViRDKuGP0Up+
Bpo8iN9RlqKVPr455FRK2KSQxJ+cVZWaiSwmwkqFo9spxp2GtX6IgSRjXCh8B8EOsZ/YWAOeSwUQ
eTZ1eoSdUSIVJGscxpAUAf7KnDC6ddvmVl64lvGIevZ+vlAbw1UaAT6/Wghl+ZWucljfOSseuHIG
y/b26KkPpCzNXdcw+c9d8DR0B2FJ1GjEN2WA1w6T4vq5fZhOExbnJjN8T+cCIKfS29C4tAwOudj3
/kZS+PpQ/g2peU1NjZMqXCZbnAaDetXKYmMjschf9Y64rOYfcfSXve2L38IVDykK2OzSm8fc0jlx
BGkrfNnJG23HzAuFE0zKJgSWGfhjaxDxzi6aD3NB36uJKPh6AoqvIx6XbXspnJ8b9Je/utGz04F1
70oOm2J5jKaF08L74uW/P/rtPKLQbqNtjcKQitdsQgw5iuqqWTkVWdfnqV6Zbr3jU9JXL4tlbCm5
rMVzvCekDUTdIk5hl9HRmc4NcWubyGbqCPS0glmt5vVQsIW6Ep7JXrdX9R0g0QY6KPPAZu3Ap6ye
HiQEj7Enk5qGj9UosNyNuY+wqaJZerUkCnShZPXn5T2RkDaLwC2Yt/fWMbUul9sD2/YKgll5zDc0
vroA7rc4duL9yfSPELntabjstYz321GLtslE/bcrCEXfx08VibtYhafDkXzlBHcJVsrX6Pc/97r9
GX6apPdmw13pKbqZJcb63L6IhmJ5Zd88V1LZK5avnvCJbi0X2P6rB3tCK2dbCJXvkbdg0O4p+QN6
5gC40tT8iOP1DOpLeLLGkuEzJkfhCsBD3l9ZC/drqcZ7gkMH9x8N6lqGL19P2ZmTmVR+pwNgwZnl
8+IzEKoroncJHIkDC8Mn2+SmF6IVSWHnsmKg1QTXNtaLDsxTSYU3TT91FQP2FUoAlHGDltA28Gz9
r841JOgXFHiOEnJ7QuYbs7Xv3bcoy3C2HZELnTMLIgaRNafepQJbQES5l/KNHPNkGfgen/i9fSjl
TWcy/VbwDBeb1ZwtNAwImitzJzU8OINgSPMXnul40fjS4wPBI6j7dcbhmFrtSUXqA6rjYSPGLOVK
ssXjUJwvBSPi9sokcL5XtDdNIr2rOZjPYnS2FiR2VD0cmN8UozeRYE28XhwGKxYKoiiaG5v0DNMB
TrcvkeSizl4B9F6l24MLLTutcdXzv4vO6h1FDBS9hD5meaVTtbAFE5ttQk+1FVPZdOVS7ThIoFDO
0gVw7bPW9ohMA9AU+gO+neXxuKoA9EtdF/upOvrKcMmdGw3ZOYabMQWUFuxivpylH86XTsASPIwI
TXtWeWkJt6Ckwd2cUUfHb4fe4VvY30HH8kjozpW4LAplhXm5suc0oWFCDqFsLQFPCig/HA4f2Dhx
XAiZ0aOITf+O2T8SgV3m0j5qwaWV6/wvx/cg9xaCCppzPJojUy9L4hW0ivm7ws6NT9+yrCO36k4G
XF5e6YHLYoDCezkC8ZYGxnwG5U0SA54c+p10XFTJZ2WoHXuDSFLWzCKSe0Bj6j/mORWFoPWIaGW7
0FjpZU9tFoNJDq3tIILVrntwJu/N68AHvE/Ys3Cmz9+8tBy/c+qTQdJ8xauOSMwYIUc+6qEQMh8t
Hy2906iGe3C5FZH4tzOr5UfMXQy5YKCjmDk1UYZ86LKndz9f8Pm8SsxVq5khhGTiSL+XCx2JI1lM
Q4Zt6fpb4JHLFaYsyJwOUJJP9eOdPzIuNrCdop/XMX9x/t5Y3mc0p1YqHbfSOoz1wKzHye03T7/y
13yMxcxgAj8O3vKzGksxNJWGhdC8id1l4p9OlX5+P1WFN9imTc6nXMbs2vECKTwzKv2Rhwo7ce7z
vlh2Vnr4mbJ1leajIZtAHyPRlX7WYDJ9aIVLhK8MQkNBE6uSfU1N+2qt5niD6b6sg4wvxXg47oT8
dlhvZ2le+jWIDGjmDUa4FhCXdh+NdWs1J6Rto/wR/5FxcI3/z+WDpn+Mlv/BA6lxYjqMnwg5uek1
h0XZhknSzsYBc68nJKk6RVibaNI9i7WcZpsowJaM3CDSsHA5Z7ceeWmn/ybTUSioT83F/K+vOCF3
JDO8Lhro03MFOE8fYWff/zrlIkVzjYEgaB8awqlCFy9wsEdfHSF4sWTfvJTcqzKs+2D9EvrIts9K
3bOhQqrAgY4PhNVQvGsmeZHtBWZ2v7dyR9AalKyjFerFgl/19/bdqhgBcDZoJRQ0dNUU9Z4oXgaq
QOAlHSDUBX/YEc5IunYgA14y+X22k6QWv9B+ijYwSJaTatJjswoVA1GqUA2bpUBjlhZD1XRSShif
GhkSS1dZh5Hk1wr9tR7ERU/Kzc6X8JuoxjLXUzsVhQxupKMQAA8faEOSmYMrA95cdrbGAuSP//Lq
OIOTMTJFdU24CxWDJ9KhBHfxmDsIsRWrAUw6e0IFzbzeZbqBJWp6zZqpGXgN8XGEZ7UcO2eQuihz
wkqmzEp75tkhCVxgmioBJmiNFCc9CgWg/Y0wwRzDBtp6RfvBPpKppQNy+zcv/VDWEBV/YUuC/2DQ
IPtnTLYE+yw6RQZ6JqfwKuBn53unpgnAcTXazpVFTjUxmLZ7Bu/CwAPH4oZfc3Ekp4fwrRU9HAJe
+XthzDh2psg/5cfRJi4mkBs4w8q3XxNNX3oPQoy8E5CnhCSpJZD8nGKvsgGQdNyb0E7MDwxOoK9b
pSzJvx+oSBEmqQwwBRwWzsN2oczNx+EHg8yfMuH3SqB8MGEzftF1TGJnCPICvK0YGB+aXhV0Kahi
XsoStylTgqoq6u1fHXL1iJz/FCODhJjW7zuogin2fNpka4dV8DR5SrV81WdpASK0Dy5l7jwdIKDb
gQix4LGATCszPDWvWSNl+Q38Ed6qeMNYdWALywv8w/zJeuPK48LGAavyg2laazasmGOswC0r8/Jd
PK3SnHGGEbP8UkbmoRjuqa4VeT/aUS4jdF4tM8/QlX9cO2HCnjMnMsuWAjcCIlofvj+SAeaeRUQ0
KndTNPg9tWOH/hWOZ0r5/uQBAZ44wEkg9q+Be0Mgg7IiqxW1fSZ0mdeOQD2fsgOC4B7sAdht0KUn
jNm7Z/aIrH2GHF02RyYSz3JRSlafkCSwQvST5o/CWogQU8G/UoWwxhuMn+0svAR9moQ8lysFp9ql
fYFfpSYlu4vxWnJqVdmJwYCKM7YODswr0FVAjbfHkHlXLXgMY3Le9FlN8LcE2kVsYxa7rlxfIn1r
JYTpI47ezQnihrXetk7OzzRslvWyRfMqALv7723uOAzlRoN/c+zvTZLNQ6fSnq9fFoOSaES5h46r
idEHZx8CJRabWfBhLMOSbItHiaN0JB/Yg91TDgb1K6ZRYFjhl1FczOu3GyO7lox3t53J5VMcyqyM
U5/SH071opOZokbYh6JWSInuekt8hEon7SgV9gix+KXpEmNiBTT+FoPeTNd9nT9y8qvIbk/S07R3
gOWBXhKkifQBdUuw15DGPm0BnBrbUQc3R2fS1JihFdTdaWKp/irCQtnhvBXLk2TrKDJ9tDMJod8Y
cbX2b68iRtJGFcQFyx7gtQthL19WlfQpB63iA+XN5v9N/bTtPWBDhzuw02mWJrYOieeffXy3e4Tm
FQn9IrnjuXS/Y2VGFYqUC1z8qENnbWr7nGyddKk9NeqSdofFEgfwDEyO4c3QngAWbgyS5RaJbPOq
BqJWST6JuZ+/yVSO+vgxhUsX/VKDl31S7m8a4vnuSito2o97MiKtlgKHL8kJRN/uxK71lSIQ057/
nciOAcPge0sEl1GBiE6JqDby9kLTs9yCLDnzdkpwe+WXd3zRyFfEWobR1S2cDDJLAFEJTLtSLMgc
G575oxPb9Z6pGnhpN7nLd1jX7DqES3+/uTSRQx91oaXCW3PwSRIIRF/JR4beKb4JDWrhjVWzeCHN
47Ov4e3Cs2WJr189SoXxnslLJTTIsmeM3LIYJWO+Ags+WHVqV29TTYECewdaYipJmkLpdaHvj/Ql
tNrLeip7qSU4aDnCUVNWDZ/5+pqZxFBqGZUi0PG1nWXUxetmX8Gj9E8WuI/Y6JMKAlMnjpwbrHUE
depnbywD6elkLxB3jGI3dNRtKLegTNJBQcYfo060IMiRMBDF5Lwpmm7/1kRSZWx9rlZ+epdO266f
yhWDK4qoV1D8dMXBd1Es4xBvPOP6Qia705/YDus+fUj6S15dZGYpRfbrg9RlzxASfBwMBP0D4rmM
1Ift+IM6Sk/ZoUcq+/GxJJpPAc8N0zcRWbILLvQuEexUIHa4tEEAU0O5tgsr4V/9kZGyc0iGqL+H
IyORHbuBNh84EvNCD0ggiZSmnqLSV8HujM6coQdIknXKaSc4wPT3cb5fOZNtt2xLje/k/HHXCx3J
KMaSUJLJq9VFQukGEbuTYHoAPG+hG7ak6yPFGX2GlcSKI8t50ES8HhJuN559Z5VqWvbeRCTWmkSh
E3khpd6hQNEql4GIPfv6ruTDtCGZKxawBou2RpZftVr1skaIRfCcyj94H5hQiBV3ZjeZuP+NrnSF
Dy3LRbv5BpQ8Y80luybzpw1exJPEAnrlAUHMW5cIR67dyppPsPQKMPu6Ib7Tq+MVMzrpmJ11ef4G
f9M0vvRe9FPzxZuTNvhm+hCeLkVRM97/EMxLH9tkRgoVbWqoHbLtGpb7NGTD8YNHFu7ki6fdJWuQ
b0KoFKKOIZ5JvCwZ+CanvCcLBcpojU1HtTCFhPbrvh4FDtgfNPYO9vZqhqbmZEkl6BDNb32wDUmr
Lvzf/sJMdMCz9/Zkz7bv5Rj09OdYiR4g64chZj5yviC58mnfvEBhn1gjo0JObw+xobctMSYhaDqR
Niu8KoWc/1iHXEe1iSWY4SFFGrvcdt3gxhmRxhcW2mFT1b2TQ1l1W261NwgHvh0/4I6quYe2yM6d
KnpDNDLL6Eg+shKXsHVfQzjpDkRb6IgHwcu1xM2OVRQ9yKb9Qx6JujPENBHZMyYRJDfSK2gesfIt
eTYgeEdnJ7TlvzEI1MvVucGCXbJHAgdhB2mWU/E/3mS/6ygmT6ZmbQDgmLfh5XkkqVDEoMerLpWB
OeIlhdfFZcBHk069uXnpJByIwSNM+okz2BHCd8Uz6YIQ1g9nst230FH8CriQ14VE1vdjyBoybFkx
hY6O6Z0fCaQtANvRAqMik/NFevTC9cPBO/PZkmdvja/jgj8iGRd1d60VxcEsO63OxCl+7XWO+sNW
umOUGzSBk0/po5cRYWtJvzuATdUk/ThwmRDI08DdVk49nXd5cjJWkoYf/AzVs43uwT7wqX5Bdn0g
PwwMdz96S/VKs+HzQeyNhx76+oE91Cc8fB8jeK3+PL++5iJpX/4/Efx3129Sk68VPecP1gxy7GN2
ieXzaobvWu//VfBKuZXt8WCJvIcf00y0VCfyp5BV4/HREh8phLij1x31yyc9OIUCjilD7puatj1i
UeGarrTrduvI72xtRKYrxJXfMdVrcaV+ivhdytNz3ymzoVKXOv+zSj02OoELdKjKa5adAw1GkBCl
UpTWk+Cdj6SqbsOvxw5/aD/p+xerWFZiImKbUjlI8ZkTSxSLro0yOhWx7DwAc+NvpjNHx1+OUhY6
j+duRqdgGMOOfobxyAIdii0IYNl/sSrlHDEpIZlKgJqcTZCTUpeBiDw1KrQMov6RErcIHo7jXnUq
VWRjjT+4hEbfRwv/qgHHPawXsiPuNwPW5eFSMKjZhWQkXJX2+C5zlKQCLGxD/5WxolxfKE/pvmSf
psEipfI5xsbCkh/02KUMpx1LyzhAYHf2mcnGQJSWsjU/IpHdIv6w4PtvVlDvSGa4DAWjXTnxBMVz
Vgrsf52cAjFWTvbxA4etA3FtZ7Q+QezV9sOgTQBT8fwq1hS9f6+eod9iY/FsRKLV2m3HxsvCOPXG
K8/HKwhGas6wtibMJv6V79oOEPrfke4HxsICJu6++dsFaVly25JnxTp6VXe394N5ijDru/2gWZiW
QsY0urDYldDOM71Lh05zoDUjJmBi/FqpwnHFfY6hCQi/NXJc4axofTNCFiQafWF6nJPXTt/X+mpI
KW/d6WbZc9KjMwr/mFmS/0eC/1aeqG65yR/nTtfkZAIm1iUTXyhLS3Qkc+w2Oaf8vdAUwu7yhMhv
mVmEgDsZkq6q8GVtRejA2onTpnzOEIXhhNnW76SEYkIiCUBei+aY4ZtgpRnw3DQAk4wXYCDk6DQh
mh4doFE1ncASpu/EzndakW4y7YbkMCJp9GE/vd6at9AwVPNlsfk7qFC979fq/TW0nosu/86di3w1
1rLuLkK1jW+notYYIl/5Dd3nepDEepi9D29sqwkEP3Ver4bujOWpYSS/uTobvORlb3bahGEcXuz2
ayvBykL98By+mvH89j+zYCEnAoOoNIFqhABDHi+gBsQ5UAW+UOeutlsJf7KfD13/2wuHDuSn6Uw4
P9ZLGkdtDQQKXqQTKk6pfF4YrhiHY8DRteW5UH9X0fBNZI1ZayBjjPtqTpOdltX2wRXRksOlGdhV
e8sOOpsFLoLFFyJ3X4TDlBXfPg7lpasXNGLfc3bmS7WZZ8vIW5kbU9HIi7geDLi0lNN0eE85l+nQ
ftdLsatqMkK3AMCUMeDavRQdfAjFSAulLrIoepngs06jbetp8zTXERxsIBPqNXPWk2tlGIVCFBbL
3LlKeKv6rzCPqjldc66eYh+MaTVtw5c4gigoUJ8jUTgcQUUhnpzFOKvFp2BIXXN4hIXn1KEBG/KQ
WrWQnN5WCIDPLCQE5HEaOsyBpqyh68X7fMG5ncW2jDM0TF02QuLG+aEoJr3bX8FRdSqfSwhLe5Lr
NeCCzWUb9sjeV1n0staiMPvlyKT+FYTQWhUkpyn37CVYNjX5sMKzGXryu3jTYTf5zeeNjNN8cmvo
BlGSIKgHl+WveCIJOuQDWxGEr/CKycLQqqInmh/pbg+L9RYwPg1eRFlKgDFylmBrVW4G4750MGBE
+ZoGfDDwA9TvQ0FaPE3mkKM/pdPJnjpegnhjvqsj48twLh6So3jEio0534jg/SeHJXxcg7+QZw4+
vT8k+rjhzKQpVqS67rqDAd+LzWk5BUEZuePZBuW2hoN6BOhbSoGceN6HcfovDowS9zUw+BZPk3kX
3eZbm7ZOrbS3EZGQHaCKwMQ2bhP+wikcM3utCRjXZ6bxNKjXshK0mgUqLVGmxMJRFibUcIDDG52V
PykcjU8fpi8x4habzQXpkVooc85S12JmmG87x55Nxgf+Eav89eRereR4IJIojRjqdIg/92Ub9ys8
0Ik7u7E1KsHoZeYg4AfPy1B+h0CuIys/TjzvutnKxSFQOWamlBKY0Av40zCduEb6+E0FMUjeNSnm
itiXXGy0ahPCl2rfT7o0a1MSqFVTUU2xXpOIPcit4X4FV7uvAcZFaa/nZvAHFf7FjvM0c8DruqJ/
vQz2OtjPRDpYvhfxs5uCflpG/RD9I7iHLeJtV61qSDiI8EilQwyDLGSFV3EP14jrSyb4A/j2DjCH
2JzsHwNKFbIu0mluSFW/ONDn93ID/3HcePKNFIsRMKKpqRO42Y0NTgGcSJAB+8clZgGgmU4FQdFU
g5bR10bb+TgOzMN4O1To4cRrgm01C6vzanWW/EO01jR7hZyXvZO0Kt3xpxU8+ql1JW6t9xejs07M
WFBq0JOXefotE85Ndc8sWQco7wDTgCbAYstjbSDdIAVCGdV9OG9OSIwsVCt8X/ilO9T3nBAxANUO
D/Xxo8Q+xatIM4rngusUur6rA/Zi4vrWEa7e7H57/+9vfRfQOzVci99Wr3zHl77UngaJUOU8Z13E
XCJeryoFJsw83B8siXjXj40AT9QmLMD6rqlXt1qcXnJz51oF094PA35wrPAVpjMd92mdfgwphzzY
SPhF4od9qItWJskv4iWIaYfQOvcujnvAQQOkN6kn25O7M7FoXSdA3InGu3sChlG1pIT8//wEBBKa
dQ3sR/+Oq/kqyzkiGcrQOGIZgRRQT/LRKKkWDTtbauawc56W8cSuolLoA5a88eIsomijNt2/0tz+
th7qsvm4dbRxltfS6/gXsz0PW1qfQIuVxg8WhVFhlA1+sA/jzMBvCI/HsGFhDmD8XHSINdmzZzH1
2/HkkmFEYruIk4VL+cFe3nU7Ttprnhr9OFgXMVaTa0XhOaXRTq6r+UOh30OJ+jKrxLIu/ysL5l7b
mwQLPaj1V6z9FP52J+f9X3UAVfGr3viNvV8i/nzeOZwTi5ey5TpZBoH9hAuN8VtEivsOtJjWI6lw
zyzGeeIIMD80nAHbZW/5VPZI8YnqHGTUvvhSZrwlur2FNPTS77HYX9qd90oGZSDX1KbDKdO3Fa8W
7k9MLtn4lQMjbpK9STRKZO/dTvt4t1uwwY23w5Df2C+UOBnmojNW2TvUvgYIAWahYGFFQLq1Fig9
vTfph12QUBKXkdpt92/bUF+4nv3zlr8u7HSgNCVzVu/BALstHTzKp2RuB57ny8TyYQQ/XRQcOrd9
Y1m7n6lHRJsfwjEKItsnauxGOWasgXzcKhqWrPnl/CvfWB60Tnk4cWQRMcfYpit/9Pab8GBsyQrb
DAMQzZj8cldw81ny1BPDgEvbTQuUXmhLIdnVUyzO/2Fo9ThGf5emuZ9BV9vC4VAzUTpB14fyk00N
GlcPI9AKmsoT8koL7JGBJnT/9xG8bQ0XriiEbMJzHFzHVWGyEQN81oaG4MJvFrjjJUZkZWoVDa8x
8hUiwlIUTGf+NpxOT22z4rypjYAHP3aA+9OUqT94XHO1zGZYPg72q+bxQDJsPbEs6S46eSyjAvdH
sMKW9hR4sBL4GzS8zAHZ+ZYvyqRgDQen/dFFzaO+WRHKQDzVosUSfQD3eU507eSGf3I5XMgeVaR9
Raq/jEX6NuCV/E/WYkZpm3EJO187mQW4KwW0wSa3COLW+SoM/7tniLIMItcLsOaJAdMQVjHrBb6S
IWurrYZlcC2lGabxd2agjs6uUcSX1ECkV1MGDuAC0I+CKVzXpYgOl+sxW4heCAMx9wHql5m/GBIO
DU7Xc8c6dOrbtINAN90K+aeRHtXmrPsX6yySvximO/gyZjA64EA3XI0Z/xQMaEKba+BMO6ogc8GU
nnzJt2yUvEJIGXtJbnT86vV7pONMxdJK+VlZwS9bMF0MHiNtL1ewP2Dxtl4U1r1rV42CIuzJ1Wtu
S/pjsj6xc6kKJxbIzwiBb3RNergXf4NaSNGsF2Tp0c7BOzakzNOO8lrtJAvLxexYREwYN1MySKnH
yUb1jeUAouDIKOEOl/TvgDOLbF3E8GwiFwgBfJbBvZSj0tWIDRhUKk6s1cMY1TLHXpVaHgV7R1GQ
+5qvl5ac5F6hPJYBLn8zp/wqowsu2piF88dbR0+OHvUcfQ42y29NUrJ6O+/AcefVBld4oXIHu6ab
MuO76DtG2P/Kx+5pv04DKuAkIUeKWAOqFT7f9oT8Skjcu65wKxq0gBk2BMUOkskKRbXJ9kJhIgGy
6Hbb+A2m0hoRQz1YcAMTTvUYhNwJD+Ml7pouT3c9yT1jJHT2VgdJeyO4gn/wxz4+bHmASKEl/aL6
TF0GV4UY+jvWLvVCXfjMLD+2GbdjH90TH1WIkMo0ika8WagUTjLAUeY/nrSONqmrOpXyLSf0mdiv
iAKwHfOcMcHfFrKTE6EClr0XXsHdPyvxkCS3Zo4GrdBZE69nT41EDY5Y9J5bCWuFGp0hfh5hOkan
nrrlSjOAAgoRRNapYrbxLfrzzmPuK4/1Z1f4NvttS+QljFtq5Rg2zsrlZP9HXTJRGhBN56dEYiWy
+dnJuP9v06BhN0zy+nFXk2fokh9OOLtxPouiIRk7l+k4Xayx7gFj+dwHc9gd5nniaKP9ogbXbS/o
SYw5BCzZOUtnsVUHcaNdbM2uEmOcu4IOA55SCeY6uOTWFaEreKvudTFAg/UZE0Am3JQ8yuYastgi
ShnvV5S3rKHucxQZnFJWoRVCHP/UMNmwWjSALr4RCMSpqlzJTWw/JojpVJjGlHa1GjXIgIH9cwun
joIE5G9t/Ts1I5de99Ro/bQ6VX+ZfBCbOn7yczgYqSmgr0W+y0xN7fJ5yAQa38siOJaYbrh6RIDh
RNUDOYuJdLSwPzyvIHQx7tkUF+ObEweIjHToJYHhfFBgKpvrK4LWpEJyrytGyT0JPgLgOtwSUZcT
apmX3vhL3Wzz0PmKvGdLCcLaDksd37iMJswR22onh1/56C6ueC0TjQFL48YU9ThTAwFa0PjTVG3F
OamOYAlDHChEJIWkeUrtE0Swc4At4X4fRdRtfGFHANdqt4jGmZVXtACwsYoJw2e6eh1c4EDgtQEg
/sInljDlERuKHeHpSh++ko4J4mMGXsM4NpIjDWlA+Jgsx1EnIM4IW1RqmI2joNkSf726cgZNFds1
y/fhUnaWyyptqFvtAVf0TsKKWN6SdSScAmBQE5MhTDMZ7NewfX5stlfpr/1mdSFrbxC+KzaV3kU4
CesQhg8iwTjvd+CnSVPem2FJEHl22sYta/E9XHq2lWIG0d1jOkXod8YmUsKBbN0xo17Xk1wSpGME
lopOFgC1cznFYz3Bp8mEh3+lenhJ/YxDZ3s1Hrrv7+a8i/TPfm9C5hvIWF2ReWj71RZ70DEPT2+S
VPt0xsdhv/8zKlGi8Rhl0GJlcLMfRz+lBRExGv0T4SmUJVlsKXYzLWb3yyf4p371CRrm6kyBXZDK
ORAuAl0njb7JMsSCY9FvOd1/uvLBlLrYO1GQE97GCp0CjIHfWwdCus6kh0//5vu5zOdlkkz/m3eO
OU92GBTjD+MGGu48QbQDegvzXhmLNuQpPjG9IsckHHip3ikBFfGSwS83CAZxhBxmY99zHiCObM8s
PaHb7kClH2qFdRuliwfhaFIccD+0HqbYL3poN8XNDeA57pKHF63ISQlmiJczni8KX4+/pX9V8UUn
fI58TtDqNokDQ0ZNkP69+9NmSitxmZuJYdAxHEwikKZ5cGs15bWexqM0zIFLUg4Inq483vwTIrVi
Q4oiVMZ8lsPNFmgg9Gw7Jv3Sy662izgNSWSmYewz4Lc5autO4dTwsalaWiJM/oAXFdn2hAMRYFu3
KIV74AX3BFP0o+se1FTyHodOjdep2SG5WuAomDSTAIWTfe6UVH6GKR0QfzWNq4cyFbQBQndlz/lv
d8ASAyExDkvJyvHXJTUZ1/SozerXSnkAq5MEPReZMoahmLGwFOiM0xrqvTbpS243PXpXdVz8ogFq
r/HdhQS6iFBtlV6GpHUUC6BEkZz9KDc1gmGmL6wfmoeARQXYF1ZgXZeHA6B+h85F72TKgFa2zMv1
mHhXPuRNjvKsv8wcTDOqqxPjNTe0hAZhyYTsEbco/5FirxQAWz4upBF2SZTDJs5L6W1KdCv7skPi
aA27z0NKfgCRw7oKrNaGPZKlYveeOUKMHy919Xc63VHz1CIXawDEL/0nPyVpXHlbxMWrVL2nzLuM
ePRQJYcReFEaIxPz2YmbDNRCCOtzhJrdjy4UvNNNQjlmmNuAIIQ7e1S3zDTKbBQk/QOZWN4j9UzV
G5CVgXnaBKHpI+FlEItauGVuKUY9k1+KPtAf/C0UpDXkpbc8ecgdcr13l5WUB0oyBsNH902oKkk1
cSsbw03ASrbK9T5HSmtaSxvM6biuHMdE7IzAcDCH6yVHThf5Ad8i4Qk7uYyjEXLl1bLmdrDFEUC7
eGbk0BOpenB/DhjImH8JMdD/GASKIzBjiw0PFl1weqWLTJL6pj5rt0bkTNfdU7zdU026Yorp4QC7
9S5kI75Prp8OJMRIRa1VYbyGcGVHiiEXH13Ld8CzKx98UkVMy0PT84OAM8V1sFhQnVvi3FiOc72R
lYC6EfzcXloCyOJkTwpd/0pSNzxPyeR7jm+NtZkg5dcAJNIxLgHsOzh7WHY//H56Vu4vCs2kPZ2G
ErbOPvBOt/lf28k/CAYh11SPpWw0D92PvjjxLzUBU3gJPi6M/Vw8xFXKZnOIHqjlpw/N6v0fk3W9
FVcSWNY7bHwu85F25MqH9xMfrIfMkkp/B+fF9WRmHzSaMDuN6YDf8acednwxHOmoKs0pNPzHFUR5
dBaIFNCJJVN9McD9IROC/PeDyShW6wZVk4hB3HpAlpE8xQ1EeH9OwqiFUpUZCu7uMX8mZ9/FKEt1
8S5T0hwdfVwQgY0UH8bSFfnEQs0LVCZ7sXFmJ+wHrvDRDWlyZp+MBn80DolLEXk+tjDD5scb+nka
BCprDXwYUq9s6zLf43OZZGkawQmHUpZNNQNNP+Ft/uljA2uD38Dno04FWEFdEFPEkSib7+4JsaB0
rle3RXkj7Yo6ra/SFYoRZPGmf8J450vNTiKvRqXJBt9XUK86JXrOr1P/AMEQEyDVAkwdnJgho0Z7
TIKXB7PZUag90E0KthTrP8W0K3jp7p8B5F4hqXMMf/4BeCkr+SbJC7z9eXzhff8ScnvA5+R6EJQh
04/n2S9S/FBSb788Pe+BtCxspwYjOzxiaRwchqdZR7ua2yhT3gLVXGQb+qTdd4JQSSj5koglcQTf
tEIF3qdwX4HY+Y9I7F3kvXoyMvkbUlape9xwSZ5DKgF0NJp7yiow24vCh5BZo/z1F5TjilMLhKE1
y6joULuvbhbvXwe1p0nayCa6+PkOINXJ/DHHN87rjCg3s/Tq7zHBECRm3lLJhk2HIm8aUK3L+szH
lS7X4LVeBsfQZDsUYdTy1oS44RNEwRDOa/niK2Y1RWUJfjsn4ihgnA5+fDytInoXVpeFwo0xwFVR
OZwrJf7CaauMydGjWVGQutODRGUCZiQC/kCPjX63dXKLAayLoyItOIXA62XwgOgXw70+FJWTL4D6
Z4coYcMvOjcVMfDXKiaks3lpUrr7GmByVdNodhYiHyANyMfAjNfTxfEFcNCOSl5+/YD9pWa+6mJC
oMxwcRjkQAx+t5UwJJOaMRIaZYG8awQZgC/XtEjGGVPg+NBbfK6D4+BlO+BlXm2A+Ij18JQlujXF
ayL5h2EpS/rwKpBfZXMUhtYHSxbBALJxKniUgeBF/ZXNRWqUa40j9PBtZ7CbOlZRmYTmDBUNou1X
82Uu7hDQGaP7yAMG5AuQIPGCzaig4xSNRWrCHDOe9etGssSwvPELdxhQTPi9HBwviiloZ6xFGqmr
8OYHn1cqIeex4gw21mZMO04pXp3pzM94HRGcyI+8pjfYtX3GydA5/YJBXVVd48ksPNQTW/M3kgsc
Ulnw9vZRbGAwvjwFyDpGxCJlFPgCGGOFtbDH0fuZdPAcek18s3g/ly7KWMYau6nw/mh2HwAF/yt9
blf/iZyCEqGNNYFLPcQ43XuucaOp8e87dA1sz55d44lVAtDoEC33NRUza+67GRt6/gIIznYe0vMb
CTLL3zyZVjs2QbXxpP6aZbusUKT3qqGq/31vdSW7QAQzc96DG7JG9N/GRgSoC5BS5HIxEmqfv2Z2
4AvoqNJN4Yx+jvG6RzGgq5t8+w0mX12NaTu662zvVtUgmyoRWIY1ndInSePtQU3veH3dwuW6gOQx
sB6TVfsuKDvARK9iZ0LJVWx3AXDIG6PzdUCywI27VLdwivDD9GbnNcy0dAY7MYXjODLEwIGHZszp
CjP4Tp/vdf4Gh8u0FF/N/gaD2oLWdZ3omnaP84icDdrI0FVoBHjZ9vlxXhHO31XZ8psh2Tm3QUOI
+ZYONGeZqroZ2OJ1DVSsQ5Wo2Z8bC5jIHkEoQAwk5b1+UGooRrftLv2HAUw/oMzf6g/ermdHBOC0
wl13o//IykWbkN7OONSmaW8PBKSGd120JPPKLghcZ9yWKoJ8QfsOoQ1Ub1TU5DE1HmjNnK+A6aPY
CWm5oxVUNPlHMB54yBblecYsY7eGpn25j+F7WYDrk9rZ66ufc3y72jxWErBp9yj04eL9JjxoLUGp
H1tdbaeaug2jSf+dt1gN2Tsn2OF+Pii8sH/3PNRP8hOnO8wzJUw50ujRT5EM0/DsygXYj4zfkL+a
UTDFDhHUIfslCf4XlD3TrWOhJXylVXQQuMsrvYHgd9tZJubRYht8+U4M1Yon+u5FKrqTaY4p14MO
AyItf+P4n4NYIlu2ZDk1XffmLtAcXamW8ZMOo94YDgTd+X3u8kN3ZLAJHPegjghB6s9tUyq4H6/E
vj2rZc29LQahevpSrJ1kyOGuFK38gzMy4FnH3HQG6y1UK0b0ylLImnB5yFIpx+MgjixYGbJa1gfb
awdqkcZzZdip1c0YeB0FtCdh5bt1u+Cot5Isp269BTih0ywfeGjsRKL8P6kIm/k+az/zH6A8InXe
aLzNgkmPm0A+GKVOtgieF3wxQ74FptkEma2tyKeuceF9kIoQqfccpZ7B2RUpxJW86jT4BCC1WVbn
va1Q32eEVzMdJR7nPUImRSAXoQCX/pMOpcrXm2/E+oL7Zzr8k/bu1XZeGFzH6MpapxbFWGY8fH19
MHkjknMBQiMwRf82sFe+KsVrlPRckUdYcsB/f4k32lUF+EfOOGYGp1Yxni/tQcwaLPRZOClZ4ckE
1iH06ce11OXI31YmMYIS5eq7XSsrqCmxGsO+E8v6XFQuVdER7Eut5awo6kxigGePTME78LorZMAe
2EqJpE7x/yjPOtoDixY5SbMtjG6a5sQEHS8CFRi7CQgjV7Cx85wGPvP7IJENL42MDm8m/xIOAcag
5wvC9tPWGV4c22VCu1oZrmEWgBfr2M1lS4T0mttvxosyLjAAdWlEQL1CYqEhv0PgTJR/VVfiM96X
Ej3+g9LdTSndswbKw2a+RckrjaeUJrIY0ypHLeT2lUukgQjwjE0SWZIf82ZdT+t2GhimOBh96roY
eNgg4yyy+tH+Kyk9PBqcoqdq7Hmn3OAp3+fFmOdW36i++shiF4Qh40cNk3ym70rvEHQ8YFTvLu5i
+NphZWM+7san0myNUvhb7kXRwD2iXpPVeGSxtc01VLPO774nPgEAE9FrQGbXyArdgR+H+4Fc/YJn
fmfAwVSzuXR/UGV64TZJuL+lPSSYqjMAd5r0ucYfVaWjILzzgTU0zQs+HRMCS/OrC6UQ4DyBoBmh
nIjPfGec2ZbHDVOOn1BOuUyhJh5+I80kuE5v4x1g/uZkygC2Ny9KNYGMpSzYH1AN0uNkG1G8BJbq
Ab4+FQoQpufe8b0xIIPLlxldXtsgnuQfDKmOOS1Pq/F6x1aO43muk5TZhNcQ6FkDkXXj3TPBm+Mz
ky+deaWuFnBvYOJcq4+dLQJtLHyHArQhf6UYUTzNTrPl99o5J3Qn6PagiNH76D2V+Y5SgNOg09ky
XsD7PfzEJgLM5zHe9mPrrEbkOuu65YRsmsJNUXFsbqU7GO54bZyBN+2MbgkD45BoTKnwb3DraPab
lpfwjDjLYz+4UOlcZ/f0djlw77aku4kGniQRaXHmuFgsj+IJtAK1n+cIFKUl6pfy0c0m2Nfndgu8
zjcN1qwEVoiZF7+FvUlTpuHZwCKj6ITEO8x3BIuErBlOO2ALRnc6jY4grGdKGCAA2LUwL8khCYIK
zUI1K2CZTKw4uSYMySbVsKtSvudAR0EbY2U872eUlJVCu4/B1ZSAAJDgAFwPghMDwBgK9raso209
jPkpN2mQOBXaZRretVX3dyjEmPpl6q5r8Jrn2yN1eniCzu+WjfADcxiZ0+v9fStidxYqIXdYCLjg
ebIybrBl6HmBbyGK1RH0kHUKW/ObKMO9VYNM67Pf42VBUKC3d6E0xptra0zk0w8cYE2lNahr3J5i
ZhRezqQTEZ643jEUCQl+5wWyvmtuj/5XfVY3m6ilgyLrZ8FQKvwF+IpSASd1rLZwLrfdBrsN7mZi
UuxVWm50whIeFzTM/RYHCuj+Rd4/aMeYNV0oXwJtQT8/WLR1vPm0y6W5TrtzgB6zSj+b+x5slW0N
3CJxqr1MG18j2BeHe8qNIO0mFrNjPV2IHjuwMcwYFoZ9CfbYtZHC3S3yCVTvvjiCuHALY2pp8Ki4
laAfGR9byWQ9XKtCX/ZX4SLaYR4Owq3rrSCyIhnmQ6/AG7Jd0zhpuoufrM3IY869SwmvIHaGz+HS
n/R1V2n0UohTkOMU/ZknRvRiSjuf5Kzef70wrK2nAepFoBO6Y4GmDK0oO09KSMof6/CbUjnBNwsH
qPe5V5OLinz0lAg8jXZTJms5bAKHt2jtshTevjFQeIqhLxaFJXg6p10jDUXFZKNGXkASq+6IErnb
Q+HOAp183UjYIFazkloLmSnsR3WSRC1N8UNIimrpsVcd2fmWfbynLSiGw+h7++o8JzaPXXKJMZZq
64P0hS0alyzUkPjz4lOVX1sToKhTRk/jPgs83bE9IUbwig9nkkisEtziOBEGayFr9wh2JdmSuc/r
NyUm+F6POeQXM0F0XJYTMd6eDGV1MHrEZ+w0UUAw1UdtD0i1l1DY4NJN9KQBJsaxRSC2ZkePdyk0
E0zZrVkAJESNz3/aUegZtxpXzFQDwe3GRFljofrSCYmOdSRtYh6Z/Nv2s7y12TvMyYJSyrYrf99p
c+3DhCrL/K0MughpeFoCrVnShTKiLCSnDIdd6yZhe2/laQy9ElYTniWjDEDE3a6QQOO8xBJeW6Kt
WnM+8hV05meF5NLf1xbs0V1qLhk9t3lHOSMqBTyE2dhBebr8G6m2bVDegGIpMEHr588LvrmaanRH
QTEGvuX9Qwtnyc7+LEKf/n0+opBDNoWPaPpUMupiq/57G5XTlWlRCb+siur8DZYzUy84CtpiMKcg
30ZZgAAE/ycZo2VWip2UnRIBJZtz5Va7T7HQmn56IYQav/3W7S2G9ol2hsSIxUVey+1VJu801lAv
5qxGYPVAa2AKodck5sJsVND6NAxW5f8fP0VpFbC2uVN3905a1m5EtlV7MWTwn1M4226o/bXYV0yV
XJBvKhnmmfwmuoU3A+wpjlJ6XjvLatbiplnxet+1aY/MRZyTCW3CO949/B+NvwmLHAvEqYrP1kbm
+mKIC4tFM/iFz8XtKHB3QV3nKyZt21LOfmdQNDaSuhr1YZ6QTg8n5f8YKoIXy6cSQiRKclw7YysA
XOo8o4LFssPYVAMHI2EyNr3dRUN/0MT9rCrN58H6PCKpc3/eF0gfv//9o6ttZLP/WkyjSO81XaoI
rgFIias+MRYHLXXvo1n0oQQdT6FswmHX48NayrEheITYlvm96cdIYrjoOCEjQHW3Vbm6md3qb9/T
SQn3OKH1tW5iZGgJdYIwdLdtyFKkaRF6CE6XITlddIjsiiUvFtid0rZ54UOIIAAoEVxuThCZZVie
e7OGkIzJW0p2e9KtGSeTjEOCbQpUWSiTR2AmaZkc9wYeUwHhC/lSSGbmyaxv2wAUPZ9ky0G8UH/B
Wb8o3zeI9My8ip/+J8Wk9bmo6jko0o6c+EhLh3qft466iGT5XnaHlBsNXGOTu/mt7Ep8az2naX+2
sqDu0KlqIxHvJPWU+IjW3VEWbnT9Gm+2Wv0W4Qz/YiIXPFF/eVyXtc2ljBETjIdPrL63uR9AfNEA
i8FQzNvBiNHXkisXxjl9u46WDsJCvPseaDhr1pZ0GetFUWNw00i841G2zGdCGFB95aSzRU2QiBPM
l0ZWKWb433U2kXO2Ps4s3EYP7rgMpYzHNJ67cMfqVxb1ZowumjHWU1k2RKwAjeI2eT9zh74rvG30
Ako/lRgRJ3iGrsd7MZPKpGtW5WEUYSMAUO8HxYlktcEWWIXUBbUBESbFzW4t5rvmOyFQnIESSO9q
rRKIfxviTKDeUcixcNi+5z8k13LykCj29JBJ64SdsrVxxAQvthhKttnrx47gf91hDvt1yKznAlw/
uV1DqMsS9YUWv4TflCQ58/U1V6CKFeV09l5AYTMNixUO4Q+4hslSxbKKa5HH1cGBxorkT/Cj2365
GUHg/emmW6Qp1p4qmrLOeLMLkaqjzjG8cjEwAMrwBec805TfTbEfphNvNMP8UEIxB8HsI42usIrL
ScBDg0QuKGa/VuUo/jkbhz/oUyxw6bnwuYHSKFLbHdZr1zg58avrvF8wHOYFwvmU8nfhj9srFXai
Ajdiqv25KqDszEP55HFfZDQTF8v/AIAmyZvx9XSqAr6HNBjDbjYlFNn1AB4y8sXcyMqDSic3RJwE
P/XEwpnCIB0pZsi2yhzHv2z4J8XZKh1KY4rzZKtvl/QyuXZb1gLCEhc4PRyb7TPTY4j1we7L8Y2B
ZuX5l+TEOxjRTca76JVAEjPYk0AIP/AR/IyTGAE2gp1kYDHs94gKvv6oE/YHEPpqlaZwhpEy47PA
jwNhhBjDD8rLjnkeLMnFINtdTtk0iFUsYbtUkC8iOScZ5T26HzEM+y69t2VE/+5nXym/3g8X/0oJ
l1D22Rh9v/YKrilVXu71t4cmTJD7JWBt39TfrkRiz49npIC1+mo2gtJBhf57//6x+breqy4hUNyV
zHcVz1/6qVyq0dFm04uQ3JQdaXxg8NwbnqXjDRrUhhobWRFH9r3GP9CvHY13bVi4blErJH1fqJPB
jcJPP0Z3A/zwDTvZXfaT9pwfRlpIDswgTU9c3wws4+9BdLBfAWg628aaqyI5Ilj+xxOZcQW3P4BG
Y7kjRWHtTy/XVuy5x/ULg323ubBiSjGKr6ItHterAbJu07lh0CZd9Ei1vlFSnw7mfg1s4qJwdT8u
T/Nht0qY39KoePADOv6fVbEoC28abS2QBb3sAZGMg2PMei4mOzp7TnPaPbWoyj13b9D5uu0RzdDd
1fcX/V5lYFup+NcIW7lVOdWBG/8Q/nqWjTDJFaAktfS0P9LaWZmJd02v6kF/3KRgMYweu2WshG6k
0erHhcTB2cpvo7hgVj8Et5GsyXdY5o28zfyaaM5BQE/pC+THBuIinbJ2keqEGPx1TqtOK+K2hc/x
nXnpmEsHE4tIyRQEaIjwSFrtVyITM9npBO5z7VPtY2r9HqD6ZcZ0POT61Rhi/bKDeMPobUupPX9P
FRW0W7rIuQYu3v+TnUK4tmo9GwEHpQ+CerYjMxPxh8BhxguMnfcnT+MrPLXHwZulqFtyrYOuZqYZ
b1SfN8fp+mRA0jmK5ksDGLlzrUZfmAoxO9cjLbhNNVs7veyliCVUPhbPkYXWlwOjtC9PKKHH7G3c
k12wgwyv5fKcYOB5BPaX7uW+I3UCrvQVdF173U9EUzNGCxnGbum8B+MgWLNUlP88dkBG/6/8WGdm
rj7z7cqyLTOPDiosk3IpjpcqIBekJgYeTiUEvvuAz7XCEDtRikp6ymmHy8jqr7DkLcMWI1w32wJf
pzFmNTj/mqkwfLxxaYxMZ9aJCKmI42PYlaTOnrjUnYid8o7D1ltBp8EtF0hP5vhg8U2yka6FsUFo
V4JEfUkrZzEsuSd/qQTCsqdoeoO40vH70bpqvbBeLDDKkoF781b0aJV1kTA42nMC9zKGJVN8HVM5
c7yRsLsTHRMZ8sZm4K5Y8xK7gnbxVlXG6QQ2pk46MAMdjl7acO8c7QJRzePZjtFoLJz4YGHigFK+
PMyajtcMk6Poi8O5WAp9QdAn1CE+RMEn2WxRByReJduqfBSNjKe1TAdANxkDJ0qS3b7DsW4/L9eD
RwzVqe4RNh3YViY4VfIZ6uIaTlr7xemX20jctWZufcd8DQgoCUR+V3aIGTTTGLHunbcHPlpOGGZi
S2hhI5gBVrWLNKTaqHUZnmMgolSE1zVDrIIOjY2IHd+GTjm12rMLhgesz/9NKHxLbdrWhrpOCPTt
7krKDQxblNS53voaLeW06yia49HiTYbj7UPv3o4obDy3KH06YXnE1vFMiS06nI3kv/yV2fwnffy3
vmKEehm+N3XPJFqsF/LSavf+ATwtgyQk5rzvRs7P+Th8tmxTjKJ6Mvz92payZZpGLuTdCfdGELpw
2X/izmBowIACv93TZ8W0t7zfHOF1WJax8WOCnz9sx2bYB4r4uwcOhDqYu5Cdvn7kvo7oJx7ZLj1i
YrlPGnfZBFq0mdYkdnqJDZi00Ox7JBB+wAO+tzq7yy36AJ0+hdVJxl1kDNDQTInBRGCmPbGkmPsM
GXk/Ggqm6T2Ml/Fa/CnumxbZHiJ+hqX1VTEl4bc3HytCdYoXpiS9ibJsKJ1OymZMnL7jUQFm0TUb
V+a3c53uO12v2pC+ka3Z+3ajGxutOg0lJRb8WUrWnI3Ij0joPVHU7vG6/tp1ObTE6NkpWTr2q+Rf
2SO83Tz8aS5UveS/tLb9xzHNMtowiE3cXkHFw68PPGfF23kuJlEuxp76r1lHbQiLpEpgPhWhhVJJ
JjBum1IMLtr37QaDjRKzA32y4Gs3fr/TzRSBt+xSfBVZrVysQM30g899LgbKHVPqqGm3iEsO0Z6B
zF4BW/UCZOtVR4gTR+HxER+pjtKCKQnW0Aeln2gXy5ki0bczyXAOLK+we5a++Wm4ZUJkb3uTVTKN
saegCQyOs4euNem6UKrIrGdk0Gu+nGq+2JEcaXvdpbIiOBchsIKkCMGEj1+lBtz/Mu+Js4lOi4si
iqRrwwU5cwKa4a1oaWs4Bd1DuzZ30DMskCT7FntYxsIPR97TrKuvOWaSLav8TqN2LagYKRmBeRDA
RKXpnLPJl8nVB3jYMcokaUWh3gpExDqQEWQTB0SELge86Rq+eeSYCdyVAvx25SzwNtteiSYT1H31
Cyjm0yMOUu6fwzVUrcWGm8VShwgQr1nZBwfHnjeC032eybtGKKjQRTms6/rtvK5q4uAjUTg72dgu
IaLU63t6J/+UhObt8IQuUX3+t2Ah/NmalN24Ak57ZXVICHNfC0WgDlaL1m9WpX9IYD3wQiXo9pJM
uUe66awkFwmBw6v4XfzReAXhoh5keS+e4l2FCflfBD3RAkl5Oi+q4RCxqaZ2vb3NcqnVKZkcWliW
Idr9Hmze5aPO8snLSKJWGtEWJcEkcu1Qt7QtatxWUo4ip1B8RbmaPQa01KPoGfpigbI0lvhrOIES
N4cVxzvSdMslmHo1MTsCpOzSk7aeoHuxGIPcG3I7naD1suRxrBcmcpfFK2xj0DINtC//TSAl+cMM
h4lLDP7heEvEfK/W5ylpA6vM3QrlO4+ueC7jdtPqWFbRxvIWtylug9EgIiMX5SG52hDO4xoxMWI1
bx9Zg/c9C4wSpKDChbMCinlTgIoKuZdlD8C3+C1Uvv6WPvkH2GUHwS9WB7/nu9JYeMFh8VKWHW7U
MWK+ftP0Jc4vKom8SI/WE2yHbzfwL9sK8eGGcB5DT/icDar9SVqCW+l+8zfeMbyNitR28egS3OPM
q97ukEBtlDGe9m8ceriZAlipUmRLfEZMWclrob9huLNuMQGseQZihmUpq//XRlGXkjSL0ydayCte
lL4NyaGKR8ACeBQw0S7tUurk/ymwfIKqHs/QQiQFE8YRgiXSevrDARRHa5MoFgiqpoda3GsFhNsA
Or19yGQv9OpFQJKVuDxmnMoCiKcEMjTdGvwvUrM0fnB6YAtBJRpbouLaYYW4nm+cU9xhZryqDqPv
K98J3VY4MGm/1sIgaT6VZODSC4yS9UfChEs0FYMmgbOxST6J+KnPXub/sTAuLCRZms0mZFynH+OG
YjkUdu+fG+mclgRiYNiUODCE+4Ok6NdvmNiadivyWeHkuM4V2Z/eMjF3VEE61HIf1PmrffYgt+9O
Ef+jwMcIvwjqO9UpWMuCQcr+sw5i8Zg9Cb954oeR+aJUCkYvFvMix4ese4wioHavhEW3YLfMRWX/
pISfSc4aGDxjaUF69zJj9q7ukovsE6ygVGWGtRbz2OPmob1qWEGYDgFF70epOWSmmMtgqRxo2LSV
513G+WEpH91S/5nXb00WzwbXKx3ColLKRqkos6c+CB3hpp02IexMivq3QpBSx16p4cMBUd7J1PIP
0jUxAE/H3UwVYErTB1Usn1NFhKWrVO7LToD5Wi82K6m19VL+ZCSxprlEnJ+IY8kUyNO7phHt+dpk
yjpyRL+Aspc0Yx4dqxVTK60ipNB68eA5kZtlWJFTb4GA8meU1IfIIljm+wvAz8A8ctXh3DlszpQK
GDej78ZMcYzz9mVsOd1Pn4z/VIP+2qcXzlKRxVHMNe7O9OwQKaVTrmkBOwWaJe9TKyYZzdygk5wN
DXY/8K2mCyPWygCV+USh2jOgQ2ihKZxB1Y+mMz1Uf3KIo/AnN+ftSMyh0b9pKphA/FXjA1TH7Q79
wjzod2ndGvnNrZDpYv2UU9pz4bwTCdUpnl8kzPp6qTZCX0K+HmfmJ13tjyr5YLOrnt+OzqWlr9hv
YFnuJoah0ljf2W6ft9eDKx1QH8naPRK1GkqRQj/FNUAs+mnhFm2Fq004FEWSDDAW492rDJ1qa6n0
JklIH8KEzFtKG1F2dnAhHljHyXbde0X+5uQlIGPixjS5BGtcD1d5wU8jqYsq2wzCqNBw0KzFv2wl
Af08wuWrtdneuKhflpX/RuzYX0lieNS5JkWdkL6KM3Ho/9gQuemLQUeMhTIVYtwO0+mPVNpHEYOb
PAPjfejSNHIv1gZkPcfm7faMP+MTebxu7B6YseLEBJUq9ulI/JQEboXp+1ori678vUruzuP84kPm
WQzvuN4OvsLB2USGFLQ5cOpe1n6rMfi7eHejODn3h00yYC+4PNS6Fbi1MnkwizsbQSD535w7Kpnn
ua33u95kxSN/qa0l6JGTPcPZMnCo4k3d/CVdPL2bIuYA7CgV6hIlulQN8OHRsfGOK/bqeHQ1zYzV
9G6OKPyALRiM0Fj2/2kPcWvnGgpVYdWvgQPJd5mF2TgOQFm7KBKK0DR+5cx2MsP5I+SLUC1eDnVQ
a2toWb7D4gPLC1IinrWuBRi8eAvNIx9+UAwMczeSWuyCHDgWlbcdLZftdQbYDbyUQv4hARAGkwkX
FHzj5WiVX0hxWB3bpA9XhpTdePIuSLw4myPb/Nk+W81pe9jgPYddDXyY2tO4hBFL9vE0tDzPOqft
5CAblkL9Dr13P0FzTnL9W2qklxWsXMP00LiJlfPhqjXEO24DxRZaK18vuhxdGFYbtvSSkxWx2/np
9b7ATPBP5qMssV1U4WAT0oPZxtWp38LU3BhuV3zIgqJguv2rcSRABE6rpmY9eiuVGFQdrRuulXBb
rfrCDefk1QKNZ2PXF46W+Ucfw4okWnbWnRzLnYtLMv0PyUwu86mb1nmsueRViUTUCiMuRlm3Mk2B
qs8Vyxs5/AvKvalUWgBZuU6cxBKR7BoK0LnXUgQz4JiTfjxgYSTpSLjmOnWb6t1z0IVO85aAvinb
LOWKtfgRYMkvouNkg5vyiVq/IEgZC1lGbpoADb4hTSPB3noChbNUNOjaBULQbz7n1+bLX6TbFVwZ
maScDZLme0PwnG25im7tF1mPPcssopKa9rfguCgcWFdm60xxcLnyvyDykbrQ5koVyJIyaV8fwvOQ
dIOlbV6uZMSeU56qOVR5CgrQVbNv5lx/6Vq9QKWdKyjZg104vPNTXuk+VJORbMb3S8mLw76HClhz
Rxhyv5nG8tbXLwGpLC05NkojxRFNmC7Q05WoqJmi7kZa5rVrWBbsA9VmTbi6rcENKBmENsboPgUK
sbWr834AaHt2IyC0Z90hFm48NtQuIEovkwgs1huNf0Jk2iDPY1LKvY0h7Vn4rt2rKA+eAA8BbIRy
Vey1h2R7+xEm/ogsm51OZt71GzEb7Xidne160M41j4/hj6Xywbd5whyj0WwDqshPyvQ2wqaLdCcP
kyjh23LZjXxQaq0mR7kyhjXhcI8GhC1PUEFRYcASnGvXm7UUyiubBZaHFZ18OkzygxfsWtz3VXpv
TOdboKwsuXJOnCEGN8b7eQiDD0iMitqW7Yn0IIkJpgW+rn4ME+ZLK6AMWIWb4HVdW+U38B3KPsqN
P0hvrXpdTayvWXTAPokSOJ1gCczbwc5LXQzoqynPe4h+MzqWJsPRBV6qV7ejpt+1cDaq8MNSlPc8
/B5ER/Y+dmCfTmI13CNF1dmZkm9GuUG6y5M8SRTabayyjKt40Qx4Tn+wQsQidSTIbzW7rJTYYoAK
mRWwJMjFGuOe48KlYSnr2q1NX6fZH/WKw5n8dtw9TIP85kTJZR87hKxDdVFy7CNM8YLqd75po0Qv
yOA6oln/WhMGTFbqYwzpgb8+2ElH6jOdOxuXxwr2ATJx2DjKRkHQB75rzTjhWxT5Kbf6HWnfvdKY
PiPOrK5GElM9DbTeK6Pcj1/smF0wOwnvGEL2CxO9RzeW1NJVWmINjUgY/lJ7I1jWbWyW8P1o5jab
0FHqHlbCF9G3R1xNnp67KqMCGK/a1EVs1IYCKzN9l2MDFdeR+XNTaiFfFfVa0VAnh85zneOFiql+
LsDMNHlDV31Z95Ap7pcJtOsfWSx9yMy6cAaPYQUCUr+Sfd3xkVowr3NiwQQsM1Ug27QZb5BhA9rs
gLzjYikGhvQgW5n2wAuVtJBJoTRZMuOJxMQ/ayzXCX6MTJYhZkvG6evhu00db5xKOeoLfdHn++0o
LIPpWE5icZ0VnPrWdpglaAIJyRiBUlZUT/QYQ9khVgb2/jhzCMOEOoOs3AWcanAfcOoEwks1hdkP
EFsNG55XS9u9rXVapaa3gml4/3RyruNP8vDJtwSG6SjX66CGMzXQ9Vg2gZUwV0vormqgJtwXgJEt
4uUARHjcHYPzbmk7CX3sR1q7z9njl96NXabKqlMtLIKSzBWW95IDcbgyH6P7gBOVhIo2cMbvAkLk
DKrDCU3ILmBC1zlg9f5e+Z/F1LyqEwxUmd6q3Q7+9N88JaVemIzDSsmg3bRHwQCPSDlPOV/BZK/d
bJkvcNgX6qMAsZ47uQRhvi3ALkuswqpKPwZAOAZe52jG1ZV5YKTcZhH4emHqNihHeddviiKiuOy8
BcvzRizYgVwsxRvWxdvAoFs293RDVf83LJq2JsMCNpTHaRm0L+pzg4IKdsXCyv1P/zO8AoxEOF/P
DKSTeA6sCxN+i8Bu1bUEVMyHyjJVVzCGeduL/IA/dSoATjF+/ah0mNseOiu66/CcGBk+wHn5I4Qc
pMZtQ39kkoEVplXvM+EhE5pKL/azoT777BnuPJXd1mmn/wydMrKMivFcssaEuyqEyUU+z+WbZXMR
RJZmomXNteelj44+v2NUiJUs1At8HVjDPXJUrtp3HCYmWLFHDc1UT0aKbADK4lW9LqcrJyTRMIlP
LF8Mz6d3TqvrZjFEe6ZMUZq9Y8Lvv4s3Kfiu7cGxwIkRbDU3p9oz3b5dtailLzhNg7RKJ/Uo2I+0
myEgfQIO1KU4Y8IVslFtTqqCWoT2cc9AfPGX78JoXTCLiSEmBmZZq0+yIT+mQCGyOhak1tUewIUt
x6BlFBpMDHxmQFzWT0/TNMWqZhRFY3GjrJ68SxtrDaoeMqHoIj2NQ6c/J98+roHhJn61sbHx56Hk
YKU++3ejD7X39Yj3xxncLyxFIcR0geE8MwRjgIcSEa3tMLf2cvx0bEfJXoYPfLXc/ccKsXLnkdzl
LZWgtwDrDHCCHKGcVqlObRfsLeVAxwLKI4HrJ5tnT6noe088i+J8XiHE6TGkjXph/TkPtUOv2o0u
Ms9NtPIwCykjh+L1PrsNOLEWJcB+PNQQYzct4od1DQqeqFGOu3S+/hVBhI7XthL+bcb8Nw7OepvS
0ASl53OIIvWyb2S3wLkRAYmCCxz9Fh1w+JwndivnQNnR+phFDdbuZfDWsYFnN0auRX8IIsN2wk0X
qfDnYXXeuj/3qaGLuzr1Y2V6WDatqpSWdQ1/GNdl+CgxB60KMGR3DjUiYnh+Jh25DJD1MRIquVlw
HxEwMLd5kn5F5iTdolqyE7flogxZcqBzdyGy/GJqN2dEdpu1cDaaxBuPSr7SkmCy8iIuViR02ftX
ei/cXPfxWyxHag2USUlzV1l2xZxPDBWgj5au/5KyUSII6Z7qPmI+MxFUjNSANgC+WibSnd+Qfee7
Khz5/zyEaLwKiboFFY9hCas6AMh9ZBsHDjiUkAookZ9/E3qRSZcaQh3VKoVtFPm+xlh6VTXvLNrx
+onbGtYVwKEwO3XuncyQG/ObAhyDdsuEOIzWEJrlzNhKmHtjDe9I8uYq0uPcH+kF0BtmXCvnK9pF
mMMVy513m9bsQaR+kZNcwmqLBC8MTn21Y8MukET+H1ww7utTZ6aXmO3cMPV41Jr2lpMjSh0UgbLA
ehpwcS9l+DQYwK9J2WdtKyrqy/v+YUT+UoY63NTXEDItk039QO7azsAa1NTxOjS3dojdOh2oMfkQ
czSEvCnBh4Q48Ss4cqPqjYaTgx3ftHu7eSBKq2BPKzzDAmaLgkIW7dVkdVulwJtwdGyUp7jDNKz0
XGWVh99BEs5Y2XLuUuQemRPLmelifYPozTr1cmcgcvdOJ/bHu26UmH/aQ9bI6/3BC/S3mW1x9cpf
h+2aq1dDsVPkLSS6QWT9KNKw8uP0rsZDg/BKfESntmkeV8mFLsVMlRdsC7Mm0smm35W7Gr6LHv5U
rM/mPmzkemAZcrlZiTlZoU+6+Ksz01zmwHGBT0oNtc8131kAMT6L4TETBeDZzM6V5FTIdqHJYv4F
Gq3b4DVULNuLRzMTbvek6eyQU2Jkii0eLk2MZXwf8OqWxbUoMSXnEy9SNucVQeNDKA4R96y6UJyQ
O4GAFUw7z+R0Lo33w3h4f8EuIddImfYiao82SbDeBUxfKwtVnJo06kLex3EdmdjiYw5gvhB0z1Z+
cUditeoU5ChItfQ55WmeRFnrrtGDDnhO+5tYoEP1u1TKD6dCHVQ7dCWbVKQ1Yo5t5lxO7b00xkco
bd/LIwCqQKZc9DGSRt6V8mn3sv8N1YnSkweCRhN3Ky2BO28xU1J/OyjmuW/XhqyKVuHiBw/pbDOI
lTE//2b0YC9qH7ztIN3ZMqJhuUZgexLOPEvmPphyu/GfCZtQSacBw9brKH3GXQvEpw/0c5GaMMpa
5+qtl/6hsWJgR7d+UgaHp9O47MF9rRbmRjwyyuh7i0hxD7F8Z3Evik62knA2XIEYp++7ufBTtoAg
IBXPT6TyLVJrh9lVHgO285viBZeXovQXWKXMMZ1tQYlpEkFdzxA3Z32zbJLG70ZmPqY4WWjX1bNj
6HgL+jkwb0WlmxSp5MsPPfjsK3XfbHkZiuw5B2dit1DlAW3icANmoxRV50zN1FK05ncno/9r10OU
Fzg1a7ANfjWeo7LGI2VzjlHvUdtptzGAh9pAmyMhr3Pc2mR2LCbKw5aBxwzXXoEh0EjD0Cv8d8dr
3lmVqJr436+vaffTdTGE/VeS+CoS8Jqs5zSfc7Lv0oFsoRugntOR4rYZVJcJaVbrutMeyMMdJ/EZ
mh2GvNNv2QLnrnLk3itjleUAuLf42Pad7r70VmcHylNO/FO1PQ1fz/MX8089OdhU0tLUzeIeDhYx
HkqZHL9H+WMsBepcEduYSs9KQEK1bQiYl0yvv4m9EhzDI/98qzuWV/O21f9q4LSaseKTvyJMuczg
sdu4b6ozvgSLpsPRjC2O4PdBzFNu5kbTffZN5wzpWZyYd9uXBwqaTbzbWR+ZmtP0cB00ptTJnF9W
YydIfM2Wnz1vzYK7X/lx88C56gkA79jlmkGbhFSvcbusutW5nTZVt7+TS0iv7IufQ4HQ2Iyb0E5S
Yh1BQdGkmHZ29SqOHPbql3Pcg6JaOSKfRSL99uvAve4Rzo+p82R6w4mVzrFXr6aFsGT2co/0qNUg
yzBNfc149Jfz4Cz0qyhHExH6aWObk6vkLvqZEWe9ngDSkEg9v3hTV6m8/tNRKBXzcBhmzhkqfxF5
7IGNRJmwGOM6d7mFdxltMoGLqSLzSxBrByu9h4fetloK8RcwmZcz/h1soBgnEt2K/h50cb9gNZTi
DDATV6ifVqzMuDtfk8c8Qg3OJ1uq0zRVIlptTqIgzXq15BBZhpVH9Sdhk6e+VbY6MTKgbYMOkpYs
jvjjUFBA0xveU7SFOpNywrkJJrmUtAKW9PYWuE4xqbFGHS0lGFKlmcBZC4oCDceS7BuGVjzuo47Y
0G2iZu5zjKxRYnYpeWwjDRyHVd/UXsRPVWINYpKUOQriBZ4fyPA9ynQBQPWCRj4pXmlalZKxnlgq
IpvcnNGuaXFvs1EzcoDnQYqQyHpLSTlP1sKl4JrtfuGfCO9VW52oNJGGVvMH0gDkykX0TydF4+Ue
uWD5Qj+tP8mrtzM7knDL86zc/l5barhjI/3JYaeDjXGhDaXfhZgq6wsj0VOHwwIDuFdWnDeFXEL5
+VlJ9gi1O43j8b2fDA6fFM9O3lyVM0YHSPNBA2Eewgrq4pjwfsDRGR4ulcDAslIseu4DgTlrPaGR
epk7k4XzKsAaJkxxCYu1HJzsf42Ih/WB8zT06yXa7RDlMcQ7NDyyQrQqx0mNr8eTPLyCkg/zOYB5
z3v//XA8exvsf0RxKkidBE/HPTvCxZO6hMq51B19nDm8vpGeo/HIWkIHAp2NnSOQS3ZIINKJyyn0
Rw94cats04k3aluLg5QhlTzVnRnLlr4d6Gz2wFE77kc01XSIk/dpBzvF36HDzU2AKkSX4luqYhCa
eE6mjLr2OXRId2Lu89CFplub9ked0nCNIejouhHXviyU9eUYUL1eGGk3O244xgZU46kOLXUSbhEg
VCfHaC+V9YYBbwSgdQ3WXnhOKhTsqHgsUkRXnRkGhKcN+218PKjcI+hiQ7527HaCgZ9BAAX5209I
rRIekacjZQeTQ8s8o1dHqnU43W1exhlMpHUaZtKJWwDBOIXnq6y43zaq9WdNP4NXt+TwWWMCXdpU
ACiOKM4nN46Z5/HF4jbZ0Nfs9/0VPtOvj5YhodYGQtbpDlQqCoOKwJnMVJDA6mZSU3xLWmyJvn0t
5qmWFPWQsLd0aYiZZUWRZXQuWeMDGDSsXtAReFQrRefpvnpYuU3uGXKwKTpXcC0GzscKwP72sZbc
pK5kp31sRPrZDzn4g6Uaw39Q/2Cj01Pp1r/XF45IcfgrbDLYN1k5eCYU71B2floU+ix4ZnfgkjY3
vhH9yciuMcbvJ9soAeJU1xyREybVtuCdy/WhlKfAB1R6uXFWLlrjLQbnz3wZcIIUEmrom8HkHhM/
Pl3RuiX45KeLNqA5E8XbJTkCKBXxGg6HxaEnClqFyQFjLiXGDA57XAS1iDa6cjesA12rRAAMyxQv
Urft/loxMNq7zeWnngQ/4T3GwMnWlTklgy2Bu/PTL2p44QLfOrWoDiYfOMflmDeT0SOR3Luvhjxw
8bWI/kGMCK3FqXisiutWgel7DU+fRPCF5nxhiZrgaJWb3c5Om5DYhQSRvjm8NlGkryF6QMW7sbrg
V+zbKniwv8Kv9eC/WO64wUaKtPgqx8ilfZVDu7FPCGZqCIOPBmiHjl2oHvp7skpYagO9X8DNL+P8
mkaT3VLWfy1Iw+9Vsih6XZd/lPNVrJoRNWh47UlaXRkWlTgtj1eKYmWvdPE5vfcihjoJTvDhfFv5
8ocbTwqKFJWznqZy44h60cTVqMPBy98OdTNFzhRtRHue96UZQHhNjeZTxVNnQwp33ESDDWkorN6R
BvCdLBWXwSUnSPseDt92WYrTgBhZ75mBgEYpYI+T6vQ4MWB+pLeHbxR2YGEOJ4A+WTOTPSWD1s3+
C/EP7aLB1UCyE76M+nViXOatTmnEvfRZcAWOhTELFuZl8gP6krAWqUo6rchbPtxh2dI0zU7LMbgL
HqxjJTwZcpYFyej628yOTZ+pEkOEQlBbJWnNle1/nGtqi4pqHRBKw1pz/PuPEjyG6feBtHg5BJde
AJCpOR+jLIbM9um+89Kxv16G05Se3lb0DCvZLJWf4FC7PjRmCaHTp8HCPJPPvPMeKUrKrxwjolFA
8XiVbYt72tcSuKXAhqzbCJP1E2UUbchWGve0ER5EFzTQhhEQ3p/2OL0i8XCHA3AJrgYn+mpgW9e/
0X7sYDL9jTAe8Vx32N5womxmaDUcheEo7pcOplaFGxwiDTfP2YPwGaYQx7RJ4U1+6qJg0uuYI++0
b2Zd6MZTJAewQAuxKoeKErMJETKbPVY/UkuLNefdRb/b9AZKJgW1DKxB1zwFKDz0s7UYa/oWJs0o
M8JxeHxvwBpx+tOkPBayOuEGAWkd3WtTe0KEArkP/bMIktuOOqXpVwYjcjSstF7KQ9KKU4HG1xTv
N/NKCQuG+fK2C7UJdTlxNx/c/ufmhYN5YWMfiSg0MWuzsQPWqbYW0Ip6IWM/hCh51XcI29EDrPqk
wnYsYwDsne5qLXHKSIu7KkbX/gIZJRevP/eR+b/jZs8KWzdmbAZ3tXwayRgmi+zuklpS0CvbV/Yc
DgXecuuDApUNBybru4tMqtU/u2DYZForp1gjxf4nus88YmmciA//neCfvmfuqraH0njd0mo8CAni
l16tCZkbE7yrq+0qJFJc6ys/+6G2gKG7xG+R9WohyqPoktPi1Oad+tmHDKj8RypW8ZWGCgTwllyt
3lsceAYirWDvy93a1aBd6kKSP4r9YSUustYpib8ORa9gogBwIdo1QZJGudoPYDtlEH4jZ333XwVg
Wit3tsZ0ZXTn0TTot4h+FlUUD7aF9xZYFaRwawttV5n88s3XlUTLbZXiX60vwpaWhbZ3HD6slRh5
zVEf6Nn5Vho2pqja3HwTR054Pgr+UTRekEVrdIgmj39CJ1EyThv7R4qoR/IKDoQOzYKcJufQX707
E4Q1Ryd4ukpgX7VTfaBF9cnUvk3zBYfoHiiuTLcRvgUWex2Dmgs7zj4t896N2ZWgFXvaJEGo1HfM
+QZxttBDQkfeDAhnGfhBdguGrqjRLjFrn+HIABAWVPcPAvLUgR4hATKkZvc/WaDv/6gMfHQT3IvO
NEsV3h7tTMr9O1qhHUkATQ6gSL83hNoLgrwhx2UaxbXJRif0GVJhLj9tez6pc2GI9a3jGmRbMZl7
m7kvb/i4UBpItlaWLjEhZxt5KyZs6S32g0ixUo4Z248BeEWel2AssxC8ieX39QzvUxcIlUxlxrsB
JIub8bjVtgEh5VjgFDrB6LjFcLXxpNwFKakcXD5yLNBoUpQh1l2N6gRMoKmPsn4c/MhUE+oTVhbw
YfsVBlkHYOpcKHpfOIzBIcfc3w4EdrS2SJfFctj2xHMDBPgmkFp8MFf+n3Kp0m2DpK96+pyanufN
WIwQhgs6gnJ1wga0XKDQwWVz4o4EFrhN7SPYnFklp6TzIOoGTdsjMJuTHz/7epbLm5eNOQdcjJ66
Pw99EEr/Mwmgg0a49kXNu6ExLdAZ8nVs8ffv8gBSqQbwoUrz8uHlZCtIq9IyojSmTPC4ULgg3FZi
ySLOp+zFsq0OmoUE2VZ/+N2+y7i8U9hvKnh2BJkQeNTUKDwZ0mqwzKranUADnW0jqEzgPNaCBFV0
3TNtBE3ur+kRaUvfbcJzt5pE1bpZ2sqKfqQip9zlLOWR52BpkZ9ZWFSh2Y/0sFi+y2EtNx+RMe54
54tGmUYL7E7V5ZDAR3LrSuu9C9UDaSkMu4zS3o2sU4Yxz2saT1tywtQk8UK99iWQ0dEpHRSUaqpj
6Fm5QNHBV3EUxQb1dfeh2PrtASEbp7qoQa/Kw6OZv6HViUxqdREeTtvSwNHfBQ+nTSAA2fo4r5fZ
d3r7VefQ/Esbh/BucQG0Wi4uDTdr00sRhPmfNE/yEiHeRnJRPvCgywe+D24fegcs5Qk6+cf/b6su
uZV5saDX2nRxj/rsgIc5cNp1uCPgGqs3/Cktj93V2+/jx4VEF4n82l0XgzpiWB0SyFjY6K9WBhLB
McfqCLye25k/tSG1XFHLhDMMIhUhoh7gPMu/eKgMNynAIZiWLt82DRutvHqb63g079uL464IEvFn
3c0ZB6N7kGucy5F3SLqMgesYn55IG1RPfe7bdbp1kr23SHsLwK7X4ABPRgCeO2ZxvZozjOYe7kr0
wwR72o1ZMPhMfXEg3/RlrGCrrsNB/k1ibbfhWNLq1vXRM7qonW4hN3kcYHB+FY3qfS4bBz0nECJu
ARp7kj+umvGp/iIGJJO9duXBxg3kd4u8YPLH68183BEdY++YYX8QwcxFxfuzB0zbxxa6+6Gwtpij
LwS9LRvz9EYYMES9k+ld+gRn2FFygygpjYd/m9jxVIXYcnZY7Z2U7MmclLYJNjqwVM+rt/wJS+vb
6eUnNa5TPD5b1KcZgnM4cN4MZAWSlRaRcHdX3DX7pFrBaOUNvOFWqx95N9bB2Uz07HPvmrdHL//h
jN4F/icrwXlS4OhhkL8G9UvrUg5dnQSHJnGdjftTFEy9Ntlx8IasOzVzv+zml8MRfINYTGE+k9Me
TrAwJ0k9rATr0iyrkRcy2JUXc+tutCTvZlXMsN40A0ONFgwdQJCRLz9lC3fAYXSiVEkzs5DsoLGX
Eh8Kn0WJcdvr9lL5XTC38heF4GxhWe7NIjXcKSmv1g/FDv9zwKnGFhFYxTqfr2GLOoKex0pC6ZMM
+7ePydrA+cab9eTXq/gM6OR+NgMSKX4Ir2Z93Np/HKdW5JX5vsG7gWoUTxEz5aDx0tFwD6gUtDND
ZLP8HTp3QS4d4zHWReQHxwzflNeL5Cz4WKRf8y+tRoyE/zXlQnMRFGHwMokeREcWjg0dxpMjoZ6/
BD3sIF8kZnU8Ch5d5uIEAv/6XPTQB9k3imVxUwlevfbr6pDW28PK0FsAmGt54/c5rAJWZ2PSSBdB
CMGhQDPB/EtOUPU1vsoJ9ZVLB53hnjkbloYIDtn1rl2AdNVad9V4TcwycuJj9M/58r4sgNt7pDsv
rnIrgCotnFouMEiIqMBDuZsFawwWguI5nmdY5WsjE6QKrkTSDtCpMRj2V8rtWH1dwStABqJVNGSt
snpAGRcfvLl9kuxa0Pue55QlrJOIRz+XbgBPCwdym/OD78xf97vkZxyncHQYMGPKMcYcOXGKAciZ
ddejiEBw0rfsONLAtUFAQBu4CpJktTVPnc9ZNJ3qfCRMMhyLV+rbGW/p0Trqi48jtwRKgcXvshdz
hAhJrAxf2x+k0S93S1fXgz4kpeE9nZtIutxhscX9hrL/zAlTz8KYDPKt7BrjWTDd0b9YDLR18oY0
PPeJY/mDMIBnyGHBRS0ZN1BLrXIy7rO2YPLRhTbITAMI090rheQbF8JJS922UgqR8zTCK5glaDpJ
nlJgJpYca9S8I17P7ZZgTCsmFRs7ir1f8RbOdvAsadoL4NxxXtxwhes8fQqd1rXGyBLjuxBixr6h
yDofyaD27MiJ9FDWpISpmt+NoIJu02HnvyS1j3pUbs/sMR2jI2bH/9JDTs9zVwCHNyU14Sj/3tt6
/Odb1Fo553QULFbtqpjya7RIkqXYaAQ2N1a6PMGpccNWVVa9umhldxXbpHxiZGxl1eWNZm3AYqMP
KkkQXS/SgR6MFQkUVhrotAwM6azGA+sgvEnRT9W3a7NepTM4CDaMCga4blGZolc46/dkDAFLGDNZ
gFPU6SCBhRk2swKfdgqJDTyM5Nsno6xIxdJgFEyxaPswtHrnc4S4304wAjeKHfetyTscdWY5paAB
gNoMPWjDJSAX9trYM9vmmtLirY7bvTkvSVU8s5jJohr2yfj2XF3S6jHBwUE2fkdkmeitss0q9p64
yUixbsGbAKxhiiH2chONq9FhgOY+byGmm728dfj2igdJKKb/7238l9WLPXF07rzyrLPN8eY3PpFO
2TLOQ+J1S4QoKKtEuwNoa0ijQ8r9sSoNDQJqZpa+m8wwbsrnFFvnLSx9lXln9ERWoV7qGa9ACWkM
QJdcHa+L21DVNk9cnsdxtdtlmN2fx3vLCq7ESMydsJGR0Aq/JvoTxqK2wVnz/3w8BCB5FwXEXbLr
bUvCASTowGYvf6aZ8a/vG2pzR+dn+zNQl6L70s7rn1x1b4bsUF7D4O/vfbkYL86OpJzvzoZQ2Ibl
rcIG/0p5oYlC2k1luKg8lwFYiG08zox9OWTIPzCqrp7TT2uNmgHIiEQdKs/TRulp874qJsp8uv7h
ogjgtnSPwvAgkjgRgYiuF4lnSftAyf1EFvw4YQJD7GM15+9tPATA69BMwABevpYlaXx/VUDkJdJT
shcUKzMe7bgg/6if7SN4Er2s9m5I4KW0F1FFkwiITHW0uktSq4fZFkL39E53leRhErUESLH2uMyW
yePcupZMZRvspfdlvjHr8EzA5yN3I0N8f6FDxrA9PwmzSD60B7iEWuMw9hqhDEUzNTF7GGuR2TRn
/4E2EKdPApKgKr0zp2CvmTqoVMlsIWF3ZbWZys10g/jPwxrwMN4RnlE/UTYPvhWnmeY3FJsaNPJX
zD6q1ckuoqEZWbaJd3jlvduCiNSZUld3fu3hv9HiOCaUjdwMW7zMyejZhA90iLl4/qN2W1DCTuPK
eXAQg9zIRXCxVwuaBhiFSd/42mGMPAcM+DIMXYYtQpxbUV45EVJFiLc5BZUVCp/gA4HDodHTGb3T
Z88r39NoUwyqzdAmEjOhTvAGoDKhOH4KZkrz7Is9wYMqBaxR35ZPETice03kyZbZwB050bQK5E9i
dTa6G+9ps8vmZy0OTvru7tqU0N+30B8nStYK2C6dPYoUV4Cx2e38wKSTOKirCeNuc5M6ETgk9cU1
wo8w1OKU3nrp65pcD8AXB5esNL6YKzrU0nR7mJhpcTXGkdGM3MAUcnw+qh+Qwr9WxxO7EmGvpP/q
6BODhTQxnUuLYo4+tvQN+oqhT/+3fivycG1vbXN7cu/xf/Y1cELVpgVunIgMAr5f8RWr6hRh4Niw
4T0lMA/wkKGvFSX5QNj5BwgTdVPyxAxUAu5IdIt217iOOS2kSFEiRF5Yl9YQ61JeU9ntz8UCSasZ
ipqw9UcgwrnvhxW6ghFcjh1YDVzS/cy9LXz2FwmsS+ogaXu3ECmtserGJ5rUf/mi5fYKKKYJ15mN
VVCLct1uYfyWn7cAenVJ5b2yfgN71EvVtl0twpWtp0WqjueDc6di+Z7ueO/vXRG6mQieypAZmINj
v0GBOnvOb2kD6Kr0vJNNoL9brhBcyDnmSdfPIsa0bFf7XOvlXSonrq2Rroj9sVdYSjff8sccM3r2
TNd+K3dAvgH3GGcNJex+HyH3ZqUKGyzqCKLWc1yT9YoNAs2MTNHTetisJHLZEDMSQzi62HmDWutv
+lwxTyfbuea375ZnFY4Z6kyvX5qyt703z5tH2ntcc5lVXhVg3deZxo45T0+uncqrLtPxiTK7UcA0
admEr0esKkU87GJk6Xf7JLQ7GQSk8nnLUCvhHn2E0i2CtXnSuCYKbDxfheNkIW5NS4frwat9NqWl
jYKobZSDan3sjgtC03sMs/WAUGttDjUrOfKY9Ap562SWdHEVInZ7Ndg09tc7T/FcRA0lyw8yP/Ux
bmv/Rq7/LpakcwVJL1l0R3QqOnadNd7LCmxMQTE6ffLxoCoWv2/A/ccY3l2q6BbgdbS1gMI7Vwea
CM8pnoNqFsq51FAlVxKY7Qd3VgQDMwd1ZT/0i0XgpFbMny7VSgQ2kuGZPsNsv0ZV/dy+3+4o5atQ
6evQUnQbpriMXrvLj5w/UJ6VAhOn/hrNAZo3JhizapyetfRB/2p8PYv0sy4Olx4GgMxVwJmvMUZE
O/cDvPoAnhCRLQccscMOo4xEl9l8e3nH9/bLcu6N0b7/FVUJRsKRCSPdddEjr6/PDhON6QJxtWnr
P542ny4hs8BYlwbFr8qzjU6BxCUr+nDLxOojNjcXGESK4pphmRKayJyKG2WBy8zzrscby/FALfSR
T0x2WcfvbqMPJ1ycLiFVm5yuRSgJHyysgQtOC8LmIDSUFC78HM+xvSdr+gACWfmqihlrRCHaHrvX
yX3mbiRkX1YPZep0uXQNzAxgOFZl6RUUgvvPBFCI8Fx00umUfWsy9W8MRac1bIPKOjtl8lhEQEZ1
/EjX/f/ie6zGRR0387mRcJ3cJBfSe4qtKTyu86dJ2YT4BXBZ9/Iyb7COmgtgNl63XlFbdCMYPTV8
WBz5ZrnKoouV/5d96lV0Nl9Aq/ayGXejhCyEoMLXoUyQO9lxwrPVilBnrWtGEh7fLilDBIHf04lw
qAz0aqNXH0f/sO4vGITnPWjgqS7/YAjN109gzECKGuowUMTTvI6INZ9D/fIBspdZmnZ+sEheM98v
qhPSYOU33hg5WA7QENTuxj8sVzIDQxKnxw5C1XmY82n72v+JwbhZIvzo3HZ2bMr6swr7e3DrnZ6Q
7zAO3PQ1haLe25vZarLJE+UxVrHj/qiz07xNXjU/wWMnplfAotpOPAIs6mjXeh1xlFRaijfPeS4B
ClBzT3YTFsOFWv9YRUCvhmdvbfbHEVsD90lD9HPRG6Oul/ak4B/u7YBIjijf/F4bP1tzB68ZdIEf
PLzG13h3XEwwpcGk3ZbDcyC1Fh3cKJJ+qj7hoMTXeelBmxj0geze2FG6jgz4nYhHvNUkWJHYT2XG
GMc3vlZ5fbHKGCO7KNVxDCS0SEwnxHwh2iecSdRDsoDUaI+xOzLTBIS+UqRBTqrJfYP1QXidqx6G
1yJDxLm5eBoiBseg6h4EDa0JEqfUl0c7VUkv+yUSlVa26H4OcDjwbbvSk+s42qQhQWnwBBYkW0hq
rIXG+QkULOrht6oqhEI3ME30nwxMrPQFT4OOgHXSaxqJ848irMGzt/Xsbj9wj5tzMZ0fJBSh6obi
m/wRLI7UQxXOuNA7Y2G/s3vW/tcdxMC4iL/yq2xwVPD6qqG75sos5k7wpZLoN07ws+M8CNt7mcpB
6l3CQ+o+Jwf1RPdtJ01DBxSWvZrD/iyiLZoPfraBw93aD4ZVHC3rjsW+ANJd74oM7ZnXWOK9gv9+
8Rsx0rf6cuOstHz2WGUtYPLWq6bhfz4ciFdoBw4jpuPVouWtUQINAY3bFs5cXmRgS4x0IzLcoGLm
mqjm32HRgRtQrMMeTGgTWlHD/rKiMmiNGETnnqCXmlpwKX2oH1gbsbTfFK7mVoLhAxILPYRTvucG
ARkMvC51YiWwJh1KqcJ/ilET/TdGiDd5cZzWnPkgc2Ba0HOKP3SQeBEKma+OewviFaESIoHzcuLn
w1WXzIGw+nXtDNbdyuYFFjQIHNgpBEvpc0nqCcgu5LGnC5Od4zzKRQtEAYIFfle0CVBzJU/DkXU/
5kUnh7cGORU3IvHy4Xmo5jymvX+N9g3cf7lzB/Nv2YaWwEMerw4Hav6UrFP/e9hPjXuUYx6WJILB
0TO+0nQ/X0s473Qa0pWLyASkwUoJoWXpvWzqYoZu/B6UtxgSRkeIPs2F6zbXdoddaD8+WTWRKyQ4
z8HlpBVoe2QXonv6XUkMNQbEhruQ0HTGeFRzDN8+ARHNVib7tvDDZ4KYxj1H5RNrPdywII8Sa6Jp
dS6irggxyCvcGKdIs5U318zd+kxfwiI1vZNZfC9aRavL73LJdTxUlTYEhmeoFy3rWZKwo25ycFeJ
FtSVzaINVOylAxyO3BzcSeCZsu6vWoAEPJ8+DmSwvLj3r7mDPZm9NxzpcRIGQy5xUKiErL7PyIpb
4uu47CN76DIlnomYKsTEiBSSM/zdZbGiH9wR++2W8lJCDxj9hZNxxMFK58wwWZIKur3vgdxxlqFt
5AaMXaHcwn65fowNcKqRkk82bf4L0PncJOey46ZnV2TJzgT7ormwmonIKtbOE5RKBpKNlscg4TME
3Drn076ktH0Z+Lq1xlFBn8p5QEAp7QQOu1REcTaI6omQ8YwkEZAIefKmePMRyYa8EFL5PPr1bGNZ
5dNfMSKM5ws+fl4JpWTREau+orvw0Ynf3loP4Ahbqc5xlE6xLW5qdKOcYIBoCLOgmXq32CT8eq2A
nl6NBYMDece/uA8bk0xEmzAz3RZkaus41U2y6ZSDrwKq7bAIA5MinnsiDlfuN/+tW4Jdj2s/qA7T
8aKg4T0CMISiMETYC/0S5P2vI6PZ8TReJA3CYolGA+pUH+d/6NHnjwEWmuri+iMVYSKh/QwWEIDK
WOo0rxwWF6J6DHRS1By+q6kD9xYoE2K/p6fm4di+8M/5wBtg3Q3RvvI7fNHn4bmSstps7EuCYJPz
x/WFnv931HE1FxFTk4tzV6II51GpK76BlabvE7C5RkhTzGYCGuySqRtbuf4MIaKoNXD5KBFqlKPx
GsdCFsDckq9lL7qWrS0WZAKdwSADjixwokUeBabjpupZ7aV9A0WPtXY4q2Sxw9f0U8r3Rvq+dg2m
RWJ1W3MAER5x2gLK3KqeUzHlFT5K9FZH4kh3Mfq7xQB5NVagml13wU2EWVpotRmjgZE0Q4MbLpGQ
iwmCg4r5hSfUDZAu5LcNMP4KdHP2XsayjzfTEbAgqSOh1X3G0lj/Y4irfhtuJc2pqcI0ZOJbyPXS
DHsrYfyIfQfYlsAlsLysZlO+gThT02MazU/+dDDt9sRBtNiJspRc38o1QStYPEOEl75UOnH74k2j
YhGJWuZ80lpta81mUZNlQi63tVSV3tPTUYeeGHfhjst8572vhvSUpE5irq51wbAoximubQ3oRSCo
jS4c8D0+JFUNeWSrpDa6ZxrGkAOGmaVHL9yER0J9sutKUr10CL9SUD6QR5wYcnVAPmZMIfikK5xQ
yp+Y4WwN1FjjW4rR0BbpiaXp8NAAZoyyvC1MuA0V90NKTa/dLLCV/bFo0uX7VMnxPAs7Vmh8HTsp
MeccrD3ffuvLJRS0o3zCr2xC18lUDH8EtagbPIXJ73CynsjVMy2DhO8BSztFrwqxdTgV3g52BeQx
aal7ywP2BdyK7d+CTK+Jm9bmzcw6+EDCprB7gvFbBAyokTCPHmNdlKZUEQv3+JG3Vc/CXNV77cxE
YGJkt3dwru8hZApo2eWfFG5fnP4UwMfjP0SoXNpB3O3teSk3irTQINYlC++csB3PD/epAsmvn4Vx
+17v7v02VUgPxIiEXag1Ejiy6oF11Fy3c/M1cWct0sr4oCYZuLHMW/b6o6MpAZzVV0v6M9j6aoWN
LnSRTYS0qjjvSwGvoTZ5oOoB0KO7trqQClF8+HCOBTMg+Ajx+Plpw+injGRdYicVDDprpeNmVLct
H/0NtEw9ZIUM4jMgbWo64OG7oRXwLdjMkbxwfR5LXuSoUx3XrfG2gsBSOMx4H4SjL/TK/L4uSiuj
08PwrFgjQIsNCWPl6gcCilrWA+jx/HVffSmhPBuGeKOlqJ4/FGRPb4d8JeJdu+kil6duiN2m9Ibr
8+Q3s7SDCIShG8R/xm5MQnoFvL3wouTMeOMgg09HgfCDNmvzndrqDFf88MscBGTKlmQwRLaLHKXX
3WbKs+ffdYUKTY4tvx93uoUaQjnUwrmeerBA6Tet3Jw6v7QlxsF4x5B/S+2LbpyhRjSFuyxTut+6
I1DuVYSIMDaKFNUq9gqJGIPyi1VMUqWNcUdSqQZU/IvLu4ikMV6hYZzjtLY+qozf701KC/7Zkrl0
9yNfrF4md17Ma/xo3mK5/vRi//dsxeCdQyecbsJLOReFJ+/Y2TeWsLIhXDpe7Cu9hpetIY5xdGef
XDAJ+TTQRPLAwqdOYnUl1AYuqKs8NysyfwWpaaDGcig/ynbwPCCjuOBtjOwfNGXnNwHET4AlpvCR
AEamqhly8+ZyunLV9EYSIL53F6iEgkEjm3nc4XMooCIl+fiTYKrwbLboA6i7WJ3MIXK5GU80UXck
oS4XZLopNFS7pl2BxMJWW43uEKEqtz0+bjJ+DK+aqsBdN+hWVhWx62YwoIm8nBHhIb0aAMwl0cAx
keLZro8yEPXMaSDEsT5zWPiMX4JeH6lkGspWbHR+vuF9lXWCybpNMlEDtpVVc7ODP1MdzNYSJXy6
ofSfeYUnur21Oo5DUBTsM7wRYReC5ab5ScMEYDYQlRkfbkXQUV0T2dYgXJRIw4b2a8018CFs/ong
w1imlQBXjrthoMS94F2Wl+wjiRPQMNie2BgvHi8HdIlv4O1+kMxiEaUoaPX7uTov6Xu75H+uPOry
laDdp/jhL7keGc+EDhvAavi6fmBdkwkY08be6UomEr/UGi7lP/k+9/8fooyMlHcLoYID8JA8fjBR
izb4oUF+hZVPawK94U+c6ah2mtusGQzX/YS4xiNe7EOBtFPHsQvKWZQMCewMkYo9vcxnK9eXtMYn
OgZLyC8b/4JS2Ia2NWmHWjTv4pFljgzEArn61wHxGe8U8gTn9qpUmpU6kc7gYpNsOqietuYtQ6/I
6etcn0r5h7VVOPBpGCht9yDMTyO9XjAGrBcM8um7lUopxYv66ORWxfwd61mQkOpnR2Co55pTh44z
8TkKnrArRfLE9lrpZ0zpReMCfdQGvC/Gku2QcB4X6pJjvMQdNHE6Cee+jmp3G/aTl80Dx9vU1mEq
bzIWdYiJgUZYAYoruTYMF8ziWpDEq0xJ77PTP3gIGJcFkujugYJMUkevCpylqA70m8TLwWpNeaPE
F6yp+wrq8lmKcczuQlUp4jw4DlDWL4T1ph5TqVUzDdo+xFJPCJ8+yNr59Tcpg6Zu4h9REJZHPAxK
zGzX85UlbgzNapjV5J1MLMbDGIUe8hp+wSv8tPtSSMtsErU5C61FbGn65BeMl9Fa3tq0Eaz1PYki
8LmwhmhEMND96vXIEzKWGeaIB1Wj8XfoPgmH7k/GsumRr5BQGbCgKYY5UhcsVukI3J6Yv3uyu/cZ
wPFyNsWg5Udt22jMXQtFocANowA3tWajyJKYpVpTDTntsl0h1KP8U+7s7YYUqDey+Qi6nI8d3QfK
1jbdaRwBrotTFEuJNqnTHnSGqxDVN6xNuoyrlOLYacGxzigFAVm+1v0l4JGip/vMqO1WYiQcOHFc
3K5Sj1r8qpym3W632UWO7NtufTY7gYKPt2b6LQgASJbAM8b9xjUAbu8/o5UiJEWllw3ZT+zsV+Gi
7i+rVB8cnDh8KQQQyD3bACZKNWgH9fxNFZjNWt2gDmMfJHg12WUtmGy8NoJcsG2LXkB0CglDjf65
l+rfDtR5WPSmqoO6a9KSLeaFi4bWjTanKbZbSwZc/p4ykULlIMKYxgXYz+K2kmW8ywxcs39RBT5X
gBO0amtZM2wB3Su82shqsCEGonl4uR6lBFC0P+ntI6WfPwIvoch3eYOVBjzTyCHHP5lVw+UKCsj2
L0qtCLkBL3oeqLXhcoL6MtkykAbY+KI52qQdCx1wHnKgHOwnfecCB5NYlWiqxhtCAJTmBBoUL+h8
B5GYUmPEM4afi6SOL/mO7LmDFNtnrCiIHcdIAkOMaOYLgxgyI1UIwzpwql3DMm99z3803HPUoXjN
/XIjoj512q5v4yvPpqg/tecVGqg2j9C81Zix0q5KImikBjGUUUD5E+p2VaOix47eDDe1/zrwj8/a
sjXpqlelKeQwtTgdJzhX0tms3eFW1GFbgIV3+HsRIPUGAH3/3f994zTWpgdKnb3vO/tbeXCsOGpX
zWSopbpYy+DAHUT6JvGgBRuZg8zgSqbI5uvIsF7WCLcSFyRerbUpiDxiEXWpFZ1BiHXae/0MI9d7
5dnrVwQTYUS6seYI698lVF4x8faKvTMJCLIuHH92XhvNm5huD8tIOrdRDfEt83t5MAUj8UrL0Gox
/K/aq4YPI9xmkbAAdgv1rO4VcuHsug0IPYv20AoIOtQdoHTRwYkvLOgPExmM0Ua0uUKtzCJYosdi
IykSJPEfFTCx1fv0c0oyIo0qBEGO/zr5p9qFMlG7xarEQM7KOYDtmyDU9emUnBjk6YGdpFJHa5YE
KcThOmzvNgmyKEeiajrZo3o8K0RDWVpaSjXGFP5ttL7vkG9ltYXR+9HheZDTUZ4HiSmI2q80Gx50
zNA6Mti2ODQRmMZLUQ4nMemvl8r3h/hQ+7Umzsbr53gxezOAh5r1dBj5+cU7OiEpbt/G0V2NOdvA
NAHKQDMP2r9ePTbfkgvTVsdmXw/p8xfM5Yq4qmSTXFV2tucXt0rhSLv3z+XYRJQfmkJIQB4Fi92n
YNscfOZ8+pAqm8K6KGGLwmVQsKps/RPMjaMUWEZUo0QlpnssbcdMdQ2XhRnHgggqDqNi9bcTEw5D
0458Z3DeiYfW9ypmXPXP9z/gpkharatqyaSGmlF0TvEbTpo7QVL8lQBxMzpf45lMhjX6Waj8Cf0J
cnh7W7JMTTXKmhOKzi12TJLlZnXWCduJ/pWDQfTwdxys+GcHvyi6Q+eZ718MOU102JnJXwzKssoG
IMdEOoDpTRQpSfA4YNLPv6/McByFQMdFEbTWd2tqB4tr76frRHX8kujqGT57QV4gAiPINii6PALB
Mnxbu1ZNWHXHlhht1NwyU8iw1X/MVNGpmkwHtVN4Sr4zS/54wWKUwqFz99OOqfFDXuQWam7CbRsp
UOnHEw0gsoOcT7TUPbL0It1cVI6lRVk0XVGt+cIVCBlqhMVCdNRbEPUo46jWALKvzbMjRl8Tbdi1
7ADvSsTfWuYwgcic5cyLp+CPXQM4IWpPOeiig7d+qTA+lLNe8O7qmsOFHEcHO2289F7p0RMDQbhq
gjRBCuGGOQiWuf5r/JFhXg7PyN8wgR6MPHWqO9H1LGVSRke/401lw/1ecS+7LndtGvH8VxPmxVwe
VqkfYZEEAhnga9xDCtc8Vl7kw8fgsO8eY8xiI6MIaqvsvuasf/iAuTVyQCT5VSoQF+Qd5a7A5b0L
yDGziiO95uepH1mtFZbODZwMOvoKCSqGN2xaA/4DumgNZeakPNPdhZ9Akrhw6OJKSQwdOtA55mKT
jx5AjbGRyiuiugD+9kc6sLWX25hjO4YHS72usLG2WfFQS3bHoQ6KUT0B66pShMjKDB30r3CLFLBa
tQ9kSC7fK6PioGemb/No05As6DxfDgA9PL/zlQFxYFCv4l85yL0lQh19lDEVdFroR4rqYEAGzwFs
k3KIdP9lRcBOaedhpTnLydVKUwdqswEbZqftyegUNnLOgxUvmVKZEyfA36RJTEiIcH+hpvjoGy+H
igSz8fX50AeF8E/1MiwIrTFYoPy0gsAnVbxnabHTmtR7Q3/GzPvNrxiQ1QwCcytnlH6NS8CKxUXO
DqzbcifCAyuM2GVS2YQMzumJmLdFs+WulhYoZFIJ19terHTbiBravFnnvOaRSEeS6yXuCUaYAi3t
PeKOVSYNMZcl4uNWLEhVu/fzL7lmQNK+3H0s1pD0SZLsugyHJkst1GNd7UTc4KIOqwYyaf8KVfFA
MT4j+pYd7OzlXbuHG0ad/41VBA5Nc7+2Hz3+bMwS/TWjqsAfQX2EvWLQ6pPsN5ydxZqstoXT7lfp
4xCkvKaAfT6T8rDcTepBjI23dCJf/Ga1lj9eYbPYWzwIKUtSU+0IZfwTeeM5Y5uSEvKEGlLqNC2n
zZygNWX0QvwAaI1II+DbbcRgFtxjxud1TpJWEQKoEjF+QAsbR0KP22hgtTHKU9kY+Wkce0t/UpVl
9TBJ2AiX2QFewsTWkWdGvt+qmUiUdDRtd/QtOo2nnMEjK4Tbr5j3HCb0YdAr+Y06EIOsxirIx6Y8
ajzbXM3ojymzPL92QUX29V/fD/P2Jsg2hcI16LEKraQueQqc24eFqp/YcQ9uGJI8iKWRSvLKR/iR
uPMQP4FF6r7/Z1DG2ByTHRBA8zeQEe2rNvX/XmCD9cuhxZEg9d25poHU/5+lWA7hvraUXBD2aMyg
h7/p2uwLNQWArgLZj0r02KgILAANBvzkDEYAVnAh+UJ7XTbFZ+aOEXei1WR7F0gYOqZ6gf/0FIPZ
EegzXqflL99rWx2G3CwYq2vM9UofDUJI7wbct2aY0CC933btMPmbdHG9xD+BbFUgUxz91f2sYh1H
SyqL/MUVbSDkSOErbZrBXCKfXk41ZUziSzCsVv/tQwblh5snY7Ey1b7RoKSyDPIx/mx0LAgu7ylF
jmggfDHRM88IYVkifGJVU/2o2lfPR0rTuVEb2HUsdNVYY9Lqv6l2LmA0753PLJGPjSga7wbeR2xF
8BupkvgcNKX2A+QirD+Pbsfj1YtJ5nh7CHU3Jp7FRyxyeh1x++pRyUvyb0OzvtwZ339VP7n9z/ZK
S2TVJJ66XMN75yl5Sck6AJAJ157iNgNIQf+r/sT03QpaC+8EmXWOxq5w4Z7dWExqnrp1HjuzheGh
8QGW+fLbgCBZCc1W51RcGgQ9iIYVzLt1hmRBVKtAr6d/g8VDkp1sUu36Hi2IntUSwi5Or9Ht1M/w
xSSuEtYBUI+feftv8vQ0zycTarN6b0JHcamAILrAxgX/ae4rRBsEn8qdGqhg5vkoRlgzGnCHcBql
rSLVmmEnZaodX0hvbniSqHwVJgVPGSwLijgrZESKiTzHN028E3YRg1n4pgktsaQV1vA3f2TDq3Dl
yfVN/o5Lw3mZsMH2kIVlA0OvAFVVcLR+IHgRx5T95d2gfm2Wd66GW4ygBV+cbKNcYLXBMwzcZ7+7
svsL1ECx3mjfOsQjZVGppEpgs7/Qm4P3DMNcVBYFsfp79mH5K+VwWs9NtkspXCHBPVAaeoctFCQk
grZRb+OmqGEFd67EOymANQTwX/KqWzf174x/FOEG1WEtHdoeY/xE57t6QD9oHQ5GK/d40+F5Jf/B
RH8tbjVrtv/0DHplBnt0qAxXDOu5rHiOkzMI4osjKf1EdPnYAotIEQuvr8J5emxq5p+g8YKeTaEE
gyoFeoi2XlsbcsS7IteYE+czXo5nMv9ZgLWM7qyAUrwTNnoa5RidI72thHI19biMJpo0d+BWnzpE
grOv79HldzGETxkT607emwiZPPWZ8kNswsl+dVcigH235/CkzRQuheCPs3kropQaLm100xXBrMq5
HQTvQ9nlYgyOABWmun0rQF4l3clhX7qv3RGv8J4quNWgF05qRDNySGarUzsEutbV6oXgCZ1AvpGu
+i6v+CPg7UmVyVLIT6Wz0M2yjcBWyQY9bbyuszJZVQRQcWDtxH2yut9P5aSCHcYo6mET07BDmHAb
eWnKIsINGcNNadvqaSo2pOr3PlONjcLTHHTGpDAbfBW/NkXtb/o2vDnpAKjhgrnHaKjOkjotaoIt
0hSpdhcRnafzqOQoDsFQaFGfYjlBEBCsERIR+GPDfhS7Dyi8AQf4PeAWnZMae94zKcfC+8MILhAn
2qF85A12c7SDx17SXrBI1AMtHAA7Z0XJbHS0dDEMXEjK1wvTFUmUhmttz/lUdn1C/b7H3DnZvt42
wN3ZxE5NxHREGdo91Qxa7M7v7BjOB5urVGoGYh/WeGhkP2f98zg8iXR1bjVsbi0RsLjBvaTf6Qcm
Tbpzc7ihyqYWW5YRz9q757oFlZcARozOjAL/1RsyHoDhbuF8CZpOz8+niotl8/fGajCogkza+x57
T75G6pMXbC0NcqjKX0b6XuOLaiJPshVol5ZmB3ANHnX5MFUAXAJT+l8YSBLm/zFrqWflQR1hiE37
oQ12gQ89oImI0n/ZiTSGzPRxZGi7FjJXMMOLjEgdU9Z5BAw0uZPbWAfZly4j5dn3i/j7ZuW9cNti
eNWtUbGpV/I+C2ei3u1l4NVLQUwHbG8teBDBILBM5xL2cVzPdroJwO5/4tZ6eIVXIEu2QOKr4eWr
K3Qwpdu8m+W3rr8kWgRQ8u5HI+zUxIxdAitLxyQzVMvjGCMIYxLIcm5DxMJAoojS7Q/9Hl0lvB1m
ACg1qphfKO03JBz1DwPCdmpm5te2hrBk9rLGig+RHPxhE30aG6x/J08yYzc+eBcKSw9cd0gl9FK0
4NMoIOUT90g/oN/W+HNaxwUGKWI6vTS1mIETEsO3Pjss6MVOe71kXN/8fTWaulGp0J2+0es0gZss
m5JucJl8ImKI8TTqTWtr2eKjCwlXcS0T9aIUz7ofecFfNi4IkvRBEyt7cXGUv4GUK1fLt3kcY+TX
U4HRssuNy+zAtgChBxpG86w3pZlftHf6n10a7aE8sD3Oa6rx/t7TzqO0qs5fhhBqnz9txD6RMjIQ
Yb6YI5srUWk0VX1yP6gn0Cf9em3j/qPK/Qoazf16oHbPrYPnoStlDafQGp0lyw2IzX8d5tYaIuMf
rmzu52lfc7Y6xefpglXKeakL6sWJkQOrgl1YMScVNjV/Z546XCWPEzYV9QF4gi4Y35fZWehBrNLq
ynqXHM6LkQi26s2Y6ud5A+aeXElzfyujso6MGkUmUwcyrrs3Zxoi/gwnVEd3u0XsTnbV5kJkWQxU
kzNCyAnd7KfOnDwcMD2ljq9mMJf1/TNPds/Ot4Coqzy3Zq69eoeY3AoH8cSj0U6Hxe+/BPlkNXlO
uQkmvd20/nZYXUbLAb1otUVr4VQtSrUbsP+hmrl0LddUH4zoNJtHFoHZuxP618gHiI0hAsUxA/48
S0u8AFO36gobztWjBP9wVeB/caOX2BJUxsoN5m9L5WnvkbQTF85MfxTwlCG5FYm/Rc3mL/w7BtOG
53UrDGfkgdua5V9onL37enqpOlw+qM+VjLBS5+p7ioEeejeaEb28BbP2vZvsMic47FLX7yqeyU1v
O27UfmyZxL1h0/fQxQhfqC4ItydufG0JKpc1Ne3VSPYHFQjsl0StsAFIwfQhkUsGQwmw283y0yBY
KhlFmZkriU4JShO0eck1NWNi7qTstTOL1TqwbdkkcbQQx70P9WebNo60jhbi91AxSwY7ESRx4ia7
fofNcCwuAxdmwA+rQTzTAJFqhmOoMzIo7irUM6ykkII91DikF1reTwZprEIG0Y9Vs+XDjtsS/FdW
MdCPGl8kDRylu5g3Cix3R4rKLQwDcjvXK8D6wI+Ek1p9E9QfFUa2yfKBOpb+Yn5cX22bJ67u03Vl
DMFk7ebAniBP7eD6x2d+fhQOzYqpF8v4el4XWzWhZrFn9rJimgyaMHLqF2y4CgoIRediSP90kCay
0PDAEx4NSUV/OucuOnAMSjbsRh8T14EcJ8tikO25f0sUoaFNkeI6PZ5PbL5QTYk0Oczb/zpKGrZj
OvZ5HZzqZctxpkfcAJ/xFDgCjNPTE2IF1U3oygQjQKwiGLVo4nGmxl1yFz/WZK+/6z60gIXGD3p0
I8V+vyj8EMEBvcIvqq/AAoRdemXibc8WIpWS1uUKzWkb7gzFfbhZUhKpmKTtk6aUk3ekDpRChPwZ
0pBgrbcOZRLeHkTUwOleuFHbxdUogMHemeOAQW30kTh27Y8FHLBohCGVXEK2dhlYUc00H4I+s+vU
1l9Npd3bWmm13J14LEOfFT1Gd7qKOl+QCqD5kJRJ6X97lAYW4v963LqvB1jgGuntabKMVdnq+B+t
ueVQ8gYE1MuG1tYOj1lqPeADrhS7eZDHH7dQigrkFJlWgi8l4HnMMAp4O0b3MZStiqmTtpC/JDkD
APk/ridNFP5GOqqy8tAzlHW78/VU3PnCqyomJrBgdNVVw3BVqRZ/3jGVVqu6n2KuAdwsBwh2I2fy
4B+dx9JbKOr8OhTUeUMN4sVqewP6n0U6xaDOthfDzjMlHFjtOSjJ4DZcdbD4qGSW7KAeajlsSQa3
fC3PJuH/rHYZBycIye/82Ivjk6nJQOkW8G0C3ZgnEJKOKzdq23A0Hvu5QP+qukLuctSDCI24Q9wh
ll+M++rVfbDCHSa7j0bAUWDqVpJXbg/OvPLv3JktgRLl9T/fABjzRcjp947bN72+W4P4UwtruNE+
/VGXli9Ouai9PI+/hnUeUdeE0iED1wBMQQDM1Ouifr+JplQUKLRvRqlBlr7ZwAxJMwdIR56PSW9q
sIcS+OIWyLxLCgxGAW+9ONz6Tv4sJoBGye+EwdvNBn19Ybp8oPjHqibPrMPDMEOZmWeXe6L6F0U4
On76qndJa3kH5bciFccDxD80kJALiV5xpoJc3IBUprdB8woZP87x/spYKkAEoTYjwq+B5CwK66Zm
gFQa9dNkXnCPnKG9/yTZazuaMP8DN9sEBHBPtWj6iPzu95BdVncxRj7Izlcziq1tTMB+m9k2WQcT
Dbs0NgMorOfeS9AXAhkbFt1kgqTwl+qRU8kw2ty3gnVHO9zElaVY8UraiBTbl8IM/qvcvTkhWs7G
lVQlahvgCOGzhL4+1HzkKa3/6jcM30fUo+tA/Fc3wLYbN8HVhwRck2rSfTHixC5+7BZ4itPkSv2Z
BwnRi6Y2Bib02PNEoVkwkN3mrKpI2udEopeo/zqv4v7B+iaIfDbccpPkuXt4J2DVPcUfA4hyj+R1
Wzs/a+s5PPX3r66ih9O1SWIpeTNbvAbRIrTa6ShRqVpZ2xjj9kVqQIXEQlTe8Xkv9kqYMRbURYAP
WVjl8E8OICJfTJzzhBX3YtuW5zda6j/kgCyfz2va1k55hmBzDEpaPXQ0Wf6PC3GHWbbKS1JHTq1+
UDmdJp9TQPEQalsaBeYx9vtiLWDgrHY7NQePg2Sm9HviSJPyJ8kDGwls5jL8BJAyWao+PSpOpkfY
9w8tbb1z/GjlTeGGdNi1tlOLnGbXy2DBvmQ2jDlEcrSgSxNIBeMZ+0+qHD0ywr4iShMwEQDUZoEB
M5nXs50uAE1mUQ+Nifcp8w7GGPkLgSpsrWO9ywvskZ7ScrjhZjKxKDR5/9CEiPrJoeE/Nxxsba7x
wM9tJV2iK/NiWBbA3K68jcRKxeGeVuVbg9yER+j0sjGcIujtD/s6GI4gZoiUL/XZbYCEgnllv3Ed
QSGojlHe9Tf8VrfFp/6Dh1jzgw/t3OQnE4exTv1UtHkpROTZyI8pfRNhnWviWADRFwyubNOnLLQk
unzR8o3fJCHlNr0gyUn0LDC5s4YqTyo28nsXMzq8rfqfuhNYXKUCHEDBeUyEAnktGeh5Xrv7KRya
qIZJu6lgUclUzp3rRONQamsrtX41rBPt3kQkTTifGU8pHJgn3nLU4zP4+gbwHOXPxP/yhFF9JKcI
zHnxbuEqMOv7QZRl8HPl+RrEJCexxFT11dlmCfQf0qI0g+2kK3+NIqBY58AD7P8GxrmlHknaDnuO
bUoH9ZUFRIobL9186zT9L9fsa/id1kq0IsryvM4wfdbOErkF4/YnV9alpyfQfMwROTb36FpV/UdP
TAHT3Z8t/2i/jfGFSHSAsZJxEq4JvdtrVbLtW58TZPwuIqgBCIgauCiYcYVf0JwRPV4YXBYhFMtr
3zOPUKGulEFf+pBXahmUgTv+Jfjk4+e6o2HRXhk86A87nLrJPdoNRoU5HatdI9OKFk1s7FyhTBVe
eIbly5Sf9W5uDnGJha3TQscwR2bxP/h9lIVN6E82nWl+Rz06KFXIAHMqpFtgYhvnXp0F8fJBu2kr
0QI9zscEXDx3rOsywry7BgJmS2eVJooPunQevQBtLfxk/ef3VDHit9Vn0Ce2y8ZT++Wkxzc2+IwU
GeclLNXSRF1fdoFNEillsS7FX4roL7LszRo8jYl5/B2ifL3Z8aXoGhZM0m4IcA7/7UqD45deaPmd
maGz9IKwWRhEb5LKX6dvX6nMnAX6aoskISb/hoE95tYeNnBUIVAxMtWS44WmO5AVLP2BVRytjFsY
ou2s0ctCIr73TwZsyfoiT6CZbMgnxbM9PBwZ0rOSf3sf7QPjieGxJOvI1yx6NjPJ1pJh6yAGZH3Y
i55jcaaYtd54MTBL/tLxDR0KoK69g51CxKmLW5ld22K70Cjmmz1ADo65byMIod3v+toXMxSVUiox
krDFxvU35uXd2Zn8srPxXwkHclQ0We7Urjrl3pJsZ2jAXTR0BT5A3ceBv5cupDExsEcT3XstcgD1
Hfi1nptYNJO4NmNEkz557IFkM8Zs553f8sLb8jKio4spsy2iqAQ/QyfNmIITwREsS5omXtAtCQsJ
VyGbETTVqDB7YyD9tROSMgszkYAg0nDViO1X4l8J0TpJWHUkaw1iq1wXrZd7yBe9toa5CYtEH1Rk
RTbL3GEj2Rqz2/tFXYNiE5I7EW/4zti9V3RL8IjdkQuV9+nDQ+R98SjpW2gqgTOKRqgteIszFb8e
HATZD1Cfv4wn+V2s6up1z6cI/uELum6ffnxq+RTeTJWoHwZUuMTCohOT/1nTawQxUOIV5kRF4Nbp
boJ3gDaa4r0KGa9nqPOhTuJ1JlhWaCZUwsh+aaqLs2zOCsTGUhJr5uvRrz2yat/25VCgIu4X8G6Z
XcKCEw4+HoIi6pl7NBPuHaqkWKYVMSY2MqUBPXfcljdnhC/c1FqxSmg+is6OYynnE71K9knEsyWA
e1jcF7U/vA8pSi4PTQ9Io/go7ZA6jJHIVPRU1aVHLty80fKEkTm//RqZSzEOLWOoELngCFjdtGEk
0Fu9czR1TsOP+8e5uOi83lya9LbEOQNgzJxeVvZZys7w3gFfWdeWwxrjShJKx8kolylRQOuFNBj1
a6VFYCLb1Mv3rR8QQsAGgjlF/t55d+dSjxMc1ZS3esyr15XH7VJ/UgzQfPCrohWYEN7dRAkevQ1L
j7xlokwwITCWruwrUIWpYjrmsuHUWNF2UHdLhNggnuZsYf5KScn6X0aofbUWFtCTl939GIry/7Nz
sh7oYl1duBk+IoqUrAK0cI/h0GiqK8h+iBAbrbrexRAp51GNnzDTxS48nBhPDlxp5kpxtCK/VewI
F+p+3wN595P+04TXHj294vKWr4LV0A/PGjBf2BDkaQkcNWHbrheLDq5ufs0N9Fj6Gn76KYk8ihNV
2quuNE5AQJq+WyUEMq/Q6tQLSqg36hOtDaa9h404v6XJPPusEsvROG8eCwv5uNXRlt2CwVOglaBS
smKAAfCDTCAWc2rYvPKk6APpYRWQija/K4mfwVeuB7i1zk73ysUkeoTIGzN6hSZuakrcUVbdfJZf
AICRyx4f+gRcP1VfDt0rFK6/IIAFNNYjZ5SoXPkB76c7scbM+vV9sl2MYeHdj6+e+tCi9J6ROKui
PH0ag/MOFRVP/SGDkPtvt5bYLzT6kt+PdWp5IErZ1hUExKjxkjedHhPUYACCNPP9E5j97iYtJAOg
JEGJ1YMFno1PrLUVBvn4pk6UgZFvnZAZtHwyuQ0i/X7Nu+CxmMxPXu0ig/U/lV+M6IOpTXNL98Te
XPmmXxPFDZlqqJKK3yKuL4Ro6ieYqNaipb4rk1MfQCWrCRpNe82vU2+GcKqrWbbssYeM7xUdg4ah
CjLMVWCDtNfRKfeqw72Y7J4JD2YKTdXAiu2B6iy0WChSbFcG7x6CDvIKymdAZW+g/hPL0LVKkE7r
kXJdzuaqs6rwF+SOpwV58QXbV+WoKZmjmJxGXujTU7VUScbxc/ai/kfVS0qpPuJ7vnXrArH5Y8Pw
vJgsXLTyTHZTAymO6JNUDg6haNxO6cR/IcpDJ0Wpt7S5hzLs/dV4OAFK9ElB1mwSBh3C+vI9o67U
g9dON4DJElVJFMqUmXznrpfEvQtdfugI9XjjiJoo4zkNu07xm4Yxk7PDTkfj3k+cFP6FIm/JhmLc
I20Wd2BqQHHVpM3wdTi30+1E0eMnl0zLBrusP0KuWL70VsoNIoHhLUTI1+1jr2bBSCda/nZeCneX
l1WcKOlizn0U8dZ7C/JSaYXaYvqlCXkkA4FTpfBx38K9SrUO5j43N9XLsqP3SP+rb1UcB7tuDxku
ZQhpkQ387AXCRW8XqHEAt6jCEFzXOMKZsd1ePzjw+nPvNBhJGoMC9azGbS0EhoA5BpIEA8pPNvk3
0YllD6UgaOdoIxojQpy0K/raOcjBleinzSrsZYTiPuqqwnIOmFjYLYa/sUQcGekD6ulVT0w/gyd4
q4z5vt94D4oW8U9y/2en18gt8zx08bEzaIA06WoogpNPhheDeITh20JKU/Te+exIl/ACwUlh3tZx
kj1ZVnoE/FKqBPU809UljEGH+5GTrTT7VGl+vCxJH9ftC95OVcHC77EY+8KKSQKIdSsjLeu0FT47
WilTqefYc7RjQTqDwn9XUedh4Ihl6vgbaANsS7HW8tdIbUEXtWvxF9gzJKnHE3HGiIxOxM0NPMjY
Boggtk+NTYiMybKFmJ+cKn4UHyHXTk6EJyFZorNpYnuaMUpG5Y+zv7Al/wEZR66XUa/muZThECVw
12SFSrBva4ISDQnjVlZCdqqGMEixupV6WFIr+QjLGF/PkE45oGBJMPJCuuZ0aLsvQOIGGVx+cAgk
EzrXD3WqNyJtw3PFNsw6HUugjbyILsZwqrAO+N8gNOHzrEsWAZBk/lEUuToZvfGs5h64LQe+Y1ZJ
GYldashpsZOy16N7V6AhcU1HsYXR29HI5V2wUkFM5jVqy5FUewtsQHlLgynDPdAA/Ach6vXNtyLs
K3yrsDZAMCyBFKdXdKDg+J+/tZ96lcSgV8jfn6s0JX2joBUk395cuRTn9zQaFcdOQaMCNVVNNOc5
t/QO2pMVRkFAlsmEnHcKm3PR3dYuurTS3bkuEFqgBhvuU2OKbXQMMqdDoPfn4IKUfLU3EPx8Umrd
KPlwQr/8QdIq5liV6k9ExaVpsz+bt333oFLbH76t05VXDVphXfm5vM4XHaQRtiRVHlz6bqrHdb2Z
CKYt6c1eqjpi+mI94b8k1b8b6Gc8hcQSJ5/7veWbb7nOZho82d5CGth5HW+hcsaijBc0jEk8pUjf
XPSgc0lFkKUS4b2IEmVqvoJ2YmsTCfS9BI3C7mDCbnwp2b/yzWaX7fgrqXIjZT/G2F7eyzXcRi0e
yzrVGWhfMsG3Ivj3F4SuC2SDfXTIkgtXaPVeBJvnQ9fmmXH51UJcTHRJ2TD6ChCkjEeTLy5vbW/j
b22FKHe4gBl1l8HHmDQYbTm/eB9POBwT4qmcUsQ2mc2lqgYrl68f+D/8LV13VZ8PbAW7M1lf9KQ6
D8MmwUH4a61Qz9wNK2cge2RFaXSPM8+iRCyQfqwHFkZhTUP6jWr9n/bj1qbcipY1yItJVXxR2bCY
EVTvDLqq2qRhsmkr/kSP7wXKeZga+IMy4+wXhhiWmRmw4Ix3dhpv6JQZ+r8GHul8F8tQu2246Rlf
3darhse130hmwDf21wwRV/44IrBvZ0JDEfXjN8jC2iQaOJwrriZRPupFWtcTP9U8UHt+D8BWUsU9
GODvtkWYvhF19bcdSGsp1NwIU1yrM1iFfrkDEVXUHQYf9frsEfYlRGYqkXROsmfVOaithB8CQEk7
1uImzouymN/3Z+3TgUYw+JEQGy52ApCbrZ8BG2IgDrTOyBnbisRPVsnu65skvlZdDxhsTNXfdjrx
imnw8ZclktkJ3wzNDRL/oXuzvwUEq9PFfxukw/g8CmUBNVqOGYpH3r000eaufGUeYHnvfKl/bMgu
9CZxA9uTJc1U2yfNwuobCl99XzBMM5GANPmV8cRRPkmHxDvuKAIA8jzlxPO4lQCiIWUfXhEJfeGF
ZMJMQllsZPKHGjgjJSMjyH7qVciq4qTcMaW1VmGw54AJ2SrElShGcBI/9uoewbGU8Gh/EZ0woR8y
FkwAyCvWza88p7tYp7a+21hk3D8pY0fy5ibavFRUl0asmoD7Fw8rp9OEYovavyRRtixBEsD8FzMD
AaPXWQqbkuw/pJEA5/m0BJff+aNU7rtuBC/hunmPyigQGpzgdJq9UidI/HJhbUZhqhMLGeeBh1Gj
k8fcWto+v2/+StikwMC/WnSgdoEP2BhIeG5c099KjkRtkA5K4lgUo7/m2hllRthG222kf/2jl8d2
V+8T1pPKKWaKMzQDw1Aup7I6bemy6PnRHt1wd0Cj14iP90ixHwvl41mWhDzIVfqxJzBB1lZBWZ/q
2GvC0WNihpHfvuQ3bdAYZXbrNHIlY4CYdFO4fEasnmm23BPwnJBbY6+ZUkGfM7vrBP3bE6SewRie
c6fBFU4TsmpK+uNeXc7MPAktJXSH7308GWrRvCbHnMUFx1YlvTJKpuhdw5lU7t+0WQQ5Vbqg9jND
ids7sslSXK9wP8b8eVMM3jij5qwJWxJhvkqMlOCTlBY/HtAZIPRx+2JigmapxralFLcl9fUIFaGP
+Y6+KhJkjqxheeV5KNYZZgIBHloQ1gAZexsDkheLUqppA/hxbIrTKuFoTv2uIg+Doc/wn9ejy3DV
+h9kkVlUwfDFTM5J648LQVS3xCRewIKkZukcehnjLCcVfg6GUVve4YqyJgjgb/udhQbb0k7W3WFW
exhkhaHXDqT8HWklKIekLudWoj0hEvxEYHBCimCorYihkIu4PZUej0yUsVvMmvk58OCOoWQZZDc3
OTPJvUigBKU11pRXgbYEfbau57wDoWRIC2Es8tbF5ID6DvKjeL+z0USo6KJ4KjIKRxvY0veUGVl0
NuRZ5qE/Dlg0UiEmniENRPzpXBv2mJurQvqvSIbvYZbDer/NYExtfvOj4cFkJiEVgYJ1KkSEpGM7
MWsWeuU2jLcfMk7/w65zGohAqhi7WAMYwcxJ6i/7DO7uPI5mk5XSXY4HMGRyHcuvYC/VdAYWqmq5
SLnG9R/QhAWS8LcvMvq6vuW4Qx4jvq5ZcpYTcEpW2LGlDGRkUMYIazmctqUEA/iuLRuRNJzb33q/
ZInjdRW9CRll/NRI18gsaEHXdCt0V7WgN5NzmhQ/3qeRIE5nS3kJsevnjZyaTb22agcCZTzD9uPF
I97sWNN5EkDKQPdLfOXWKjqWg987R+p66idpjub+GURtgN+bOX9fLl+LhndZU35NjoEi1iBcDSE4
RUyDhU6wxkve6f11756yEIzSrIvoFfznxsM2Hs18dEiLRfbs8+0ALiQfV7OzKDs7IWxez1RrFZZN
4PRSSpfHa8I0ENqbslzoiIA1VVaB5UEPhi3EQl4fFs8hI+sdq8QLr4oLnBos73AZXZcRvsMA6Rtv
98tdFZDAgGRcrPnwjTT5y34ZlZzt9gvFdeuKR1PiDrjxf0nnVTvF6Zpw3mxlqScSNGhF8jWCCky+
fxHYLNz++6bzLI3vyVgZEPOGVRz18hT1UvSB1ndJZvSaYOKhwv17SK2p9RbyCqG49nH7Yc4Il8Mv
ky5rKYoIMNYrReytvn8taKA0CLV8m2mQFp9NOWM0g+rBlzvbg7PesLPOE0evQPuLQ+vjA9JI/qJY
OyqAMy4tdljQm+fUQK+dPKG4GdStHchLvTAY4ZMF9W3krmaVS7I3b7aLVtBAOczLcXgX53LlfumA
bHAxKNjqKFLFqCzPtRz2xqO1Csji85WAdkMz2ODzonQfKLltjSU22SfjXP7Wp8DMiJS/DI2KjTMV
B9+Qp9x1sryNjaJoPEMgtSzC9M1fdiY91ht9hqokpwrNFFZ9L3zvJz6/JGwsq7qxHP2QLC81Mt0K
Fs/jp/pZvIlRiH8RyA/PIh4K0BU46qu97gNwOKlxmagSN+sksS+0mp9vYBif1x8aRcdYcaFvn6Kb
mPvw7kKWMi9CYDnEIb6RnWXJzzcty7jY1TTw52Q8IDFsT4SDCSCJLSgqRTJnLlv/1Ew3mK5Lzppd
fTAja9f26G7IRp3yu1h5EzNC7r3z8enJT2uqBwux+DsvCVcQRI9pHo7vDk1oWDlHvIMVIsfBzJnP
/yQ+/t290UkmazkGPapaLda6P0ueji8K5MCjPjff7i3WXsYKc84iKJsJpMeym8MKrUQY4n/Jf6e0
XAEkRh33LbptjBpfU0CIpxqD52T4orIB4EA9fUcsSOn9t91xZWkzM3VoFCd91IXTuIyvmTVe6oaC
RzeYJMWVZSk89MDXVbnoT4GO+p95/n1Gtju2TumvAWDFqok/6J2POB14+f3sjikUO4/RExi2KtfT
rWMpl2EdrhEQDGtmqahtodngD0G0TpxRTBMJa5lLE3o8twMopsWd6mNDwcnY7JGjd/nJKNoGm7QZ
c96vX+6pO/hsr/jONotf1z8L+9UuvVqPNKp6mc15INp8Xh/l04NIJ1jwmpodgrN+n34xzzRQTqUo
tEqm95VDgUE67ud6oqM2rnWwyPsOW+oschXaVjdP/MYHxCLZLQkZCxnKBRTxi5VS7zF1TDqwVaKS
aiiW8N+Wrcio0OFnC7hZNceHLKyhcikkp2z78eMgTJgejf/zh/UoalFaXgCZASrs0ZhcMQ0jxQ/T
JOo3PBkUV/56GB8C011XUiD/Lco1VRoX18IQXL0NN+9bijCXZUev/MHAqmJkmvyu61NU177bWhBq
jtxfS8yiXWw/vTH6+FuKV7muwXde86FnhExCf1rSKH3hR0W1EyqLteFCFcpoNFe0ZpyurI2UEZlK
TOOXdzPmaeDrWZ48LvavkVnLLBvo7ejQDjb9Z2gQkvap6oVsl47E7WGOaSsprdWZHTYJxGNbErJU
xpWC65YCc7Gwz7vLC7nrmzNirXmiOKxEwDxvWkGElOkzpMPOyVA5nbAR6pjQf3BMooGqRP0y3FiA
UNFSWrfnanPXUI5ID5LmrCSK/GgFzEltIKsMhnQBBiWZhLbqiSjvGa+Zykc4LsgsBSfbg60zLQkX
s+zw9tubtCP7iC1t0Mj5sCOyrMPJOeV0c10Sl+8VccQWOvVFbkJM0kEmJhCV6kO7RqwvgOC7Aj60
TkfGNLEgl/7Ghp28NSVxeEm6wNHxoCTqy6QKkWSa1rshli7ZdLKzk4tKjPzsE8I7cEkw8VqlCBug
hvyiobcTImdZc28PhUybEv1QwhORlWh1uwYWq7wGqS7gW8Iy8UudAxXg/uQ0AOrn2URVUN+ei80a
KG/9d7qYbc7EadjL3zTMCNvyxJV4CdkTL6Am5XXlSp6f4xVDUvl8g1sZ6Rj7RIJv/xG4I64J1oYG
7nXCESahj9b9WiiFqEHgVp1rtKpvz+mjwAyEykLn/fb2ehYaJSVYL7F3/5IhdTbX64MM6TtkbWl1
iHCctUSnEmjmuKFkjMw1ihYg23/pkfHrVb67Hl9Hs9xLK0zORkV17E7vsqsqsYJ6lsUynZZh6ON6
wkfavuJ+T1VUTR5Nz/BECmgJRfRp32Esq/lpQAaFJHsKUk+l+F9xOFbRu2Ly2Uy+tuyA4DKT0Wm1
p7Rr+NHU96J09ewJbUORIGZ51IsY5Sx6hTc2Y/qUi6iewajzMRP9qlNcnmLPcRaYL04/smKCV+cM
P1dXgESnn5h8PJz9HDClfmwojmHIazfRsencMb2FVmtEYs7JnV2an7pCDr0CCXr/Oui84gL0YHwO
HEETxEpuLbxbUZ1WwFXnxCeOriFtW8/uWHFmV7l69p827Z0u2FmyK9O9DR6Tp/Z9XtVK4onOjUaw
rKwXydpByNza3lpbknb/RYAGbOvT0ugCOZglz85ke6OT2wC3rL5Rza6aXeiYRQdMv20FRgT+IgQO
hem4cjyCymQDUg6knaWqPg7oRLew4AaJNGictIxHQMDw8FFnXzPjYCIkfuicMSu67sCIN4sZLV9O
yxyR9TiouiwRNBfnmrq096/v4fSaKXqb7ih1nS96ZVcLK3rJB4W80h6/62QkMkWH2SNsCLwOohhI
Gqajv0oTL2ffaBCZqkCNz60PnQmNg/3f98HNbg+R4CooAbO1rqBQa6yGOhBdplGY3FJ7c8Thc/uJ
gYSSLwhpU37NgsJN+KTXcCS82R6stZT2Ix5KMdUZLW3fC8SvSNkFxs/7rYKR01tQSAWy7Zmo+qqf
9EfatPoH8bRktK919vAWG5+I0kqDoOaS59LamiHYmzBt6px+YcXCZ5MWXz7u4+Lde1TPZp5XY7Em
V4td7As+ZTs19IZwREleZRmqeAaJ6j8lneb90ux+2/RTxcXB25j90xVayxyE0w5s81/XSa03LdQq
GgbFIyf0slfjX0NsShH1tGpZnk7JR4L8v/vbJ0erXztGIug4seMEMfpSI+miiLct8RmIusm1v+zt
YruzvGbq3tCEwJvv2fptEFPnCHWJ3HaC3GQDWc85OmDIV90H+xnzvH5/SfL5BmqZwwvUOrf0arwJ
rNt8CrarZug6kbu77jvFHFQyP8mrlathoDmtKto2yI8Wwrn+Y2FRCis/N38VLQK3fT1ONgu4HSvr
0eOKqtIg8JqEtbL2B+Ac8+aTVqczFWxZFqNR+B2PFOJS27N6mARDe2/zvuiOeukXKLrFgH/qsfIm
jze2VmPK9frPxXd9ir0dj09Jqr/08r91Zxqb5FNyO+Ca/sVqXttDxVrs66K5/xL8fx8nGqFn432W
1PvAQSh0sYFZcUGQfZjTmxjhZ6eicgrfWtcLh4MAP2/NHwND2GsGOyh60jWvH7KGURtwcyfjbO3b
GPb6zG3rmakX+WyRwryqAf2nmqqIGe4x5E2h+7shxSmyehMjxZSr7uVInEvFMukTwpk9Uf2uM5c9
cXnh2tUQYKQVaPiZEdrh/thXO7M1fgpFT8zEauLwPOp8HnWBh10KD5gY6Vvc3ZOVO+Xh8r9LcfYp
yFcpQW1D5P7IhbfNQURbckqigPlAsBtPDtv8MDGhpp6qRDyNW1Ya/LkXjsScpmcDJnVUWD3ELuJY
5q9JA54P0WuiaGfarCjUJOj++Wjl6lI+mqZD1yCQQdsRPCGtHBU24QoIb4jjpcbqT4Az9525ZfU6
aivkxeYVSS/9RXDzgifU5hJI7TWhL/Bbpfa2/vt1yMDHxBUifrzPphWjwJa10mDZ6giFvjcwpxl4
HL1FC1Vu8X97VWEPTNJUnhiAM4h8FjirTuUPT4z6a7OseJdTqrl6rBkc0BHCJFN89qoEjoKGtNn0
2WVWng1qtJp1lRi2G7LisouHNnhF4jkadrH6RFdZylwsfIbfhTV90GtAnipq98aPC8x+JIssDdjA
MnSmyxTEoV/qOjwZKNq6IXLfkZ7Q2J2AHPrWzfNc/dtUnWLoe5qCtn7vSw5k04rBRX9Z94w2mrHm
YFl0q7rG/D8b2AMjk32OQ4555GOcHqjcft7ei3/B0rcaDLWSpEpU0P96Gwv5pbu+XuSv0qhatLF1
I+A/+6Ii+O6/VC3q5TZEM6TXIO6rwLlVAO4PafFujsJZ+BZn3DoWXERNJYG7/XabD9YZV/B4wh16
FlD7gKHKoKWOmEFHHizF2jmHVfzJc46il+igC1XyabYZmrg4/5zKZBlJrFgVawqn0GXDMhp+vPUu
YeAikPbWTB1HMSl/Q+g9S9iASb/H38fARJLFQqQNAk0H4Pr0scLpk+yeWcTlNh9mW1H10XsxQhvH
e08fylZJVlC3jdpe5vRsI5TSqtrhhwhQKg7ZKud7Kwuydi5KEGPmRfvrS+hBYbV573zEEJtekhYk
fvoEORIzhNqxw36qcwYmpD/JYMWc9lPxDHtaK/MQawbSJzbXkR/V/4N5anaJyFLhBDUdOY/EPndG
Y7V2iZP6u46ZNuSHSQ5cg+jMP4ylwH9mVOZD0RVcoVxWvI5ZwURXUbMVXCo7pYufE9277qK5gjMM
FFiROgnumcSumoWNuoazsFSldQO3Za0Ikl9r3b5oUFDeaRAtgDI4UfBsB6DdPK5BKnvkif/w8Xrr
aJ1gY/2KTa33Z1rCGRpljZR+wJ4UhiNQdfr1r8nGGTaY7MAjdSNRaihhjJFP4erV164l5Bquc/1s
4+h8L4BX2D2MoxtQ1b4+ZKvHrwMC7yaDQ3pE07sMERIkOjzAFiDjmyPmwTtVg/eFi77wTQ4h8lpk
2wBfVZyPuZUEPZ0BC60ozfd4IEDeTiyLWhdo2XBvz37TvOv7OWyIXedDvjV2cEfSU8n5E1jQe6Ub
mVnDEbyvq7QEdup8AP+LKuCq/C59yeyER6KY6WYTiVo8h5T2+w0TtZrk6GE1rfaXguRs87yDKGdH
gILndqlzb6A1nTzub2WHJcCS/nxEJ/8SZV+017wpBYh1enP/98npIAjpnojVRw0PWiGsskyt5SaG
mlEdPRy+Rf7ic4SBXg7FvpmE/KhIdbLvaR2z9K/z4wx/I5ZTa1yUtBI7fKPHDhUVKqte3JS67wjc
bctJBq1mRTW/qJ2fC5PMBBTio1bjwqrqg9QqQpCzHi1pN/uTQKqJYSh4hT0eyIdQvRGowKFsgHkT
7DYJyV0XN4YJCmE7zwFbhRiWdtA6rrwUiTrXpD6Vl/5+69tVpEu67NrgdJmfX/UrmaqKbMImKijF
0qr6XGIpqUglGMUsF/M0wVK2INKFYqB1JqZp6bZTUpv5beqlZWau6udQJx7swpdRfmhCRLwKjtdI
qMm7xa4TfanKfqYq/yxGgkMae4oRzMZEAwzSymYg20NxTjYN3TwjZCMVDmyIegCtPWxJSc6vhJON
rLZsIFYbh2akf70H4ceI3WiaX/GgGZCg1sEvHALDWZ1RlHyJ1wq+tKE/iOjFlg1y0DWavkiIzImR
NZbEUwrjk7LhKgvaleRkmDgMB9Ydk9SoYa8g3IeC680P1/ZUjN1jHDj6tFGViCWT2iR0fr+BRXoG
gHURY/eOg4XB9bTCIJl+QXB01qO4XEUW+BKod3TsURQ0nGmg4z/ErJmQS+wbYGkmg2gXQx0ijQoJ
5CuhcYwEFxry16Q+T1h5IbtUQNz29mKu4PeugFzlsu91Bjw58kTiZwBdbEQzzMT0UQNMV0gROlvv
WeUrioJlWmJaaGXUKbtpNArCEX5a1HoGDUiQj/pNNFoi7sHMuIZ9mpLogyFlONcZaTRI/mQvTIrX
jZbN9W+FXir0V9iaJWApvJOtGrR3babZHoKeREraJmegmukqM9SlllRqh/kUnkSeu2RGFBZobYiL
KgpmSi1kE9ny8A7mU67oVjPf5XLcVAbTd4p3hatdUj5VeqGppG7MuVdo8JiKGCDvgmZ0q9EqoxsS
JjONsVDOkIpmmUY8uf/62lx8AkV5+sfd7njyYR60xJ5lhCwe4Nq3w9SkVMRriHHNS4cz2PN4plN5
0NHovpR59RvxJRNecq1dcgvgkT+ZtnG/WJLQdb5FjyL8R1vlmzFGr8g5KlScZJvxavGGrENZOO3r
93NO/U1bTJAHaDiQEAv0CM/PxtDLBCafvF+AqKpwt3+oTO15YqKyix1S7/cOtvs01bAJj+jZvEok
gelcVEESqWY1Pk+LPx6y6vn11XHbfHLGN5BI2vrX7XjuO4GydNoXNne43C242ojYBV9Zr+AeekkF
cjKeJN7OE4lZEmKFS4Scv47OiGJdMuE6EUeYP3pPk5t65vvttOWU/hQwPT957/5p7k0SZymmyp4p
a0Bfud1nV+tobM3DKjZkDq3m27iUjuMOgXZMm2S2tzaIXq0FcfNxEELfvcFeUiW3dj8PjtLbHSgH
e/jta/Eun8Zo0zi+8pVX88v11L/0qsPcdLEwKnxoxQ1Rum2dtd9jHgj9cAlNJiMTXzZMZ/1SYuLF
RuK0XtNRL8uv5bhw1qg3SIQesx1MBD5Bp+1sUY9Tux8R7Km24aujPF0/wBzk1fPVYruiAOCiqwNG
nYi3wgtrvm7CTp+pofrVGfrDef0cyvVRTYiDiINvLrD95kwDgGfgW7u8OmhBUcG7Vf8Cz6QlGDPH
Rf9xBcg/Rbev/o0gpKtNNtXnYLe1rVQLuIsnOXMmukI0/iGGB99q71LeNOfS9osMY1FbkOWavNeb
JmVQh9ntR43ZtleWaYV8HWmtOkG5XxomLWp/HS5uhpRU9Mb6gN7HP8k38TxWqqUsQ28m7mqmdMut
qL481ABLlo4ZOrWE43V/2lVy6qQZGLaYrOBgputwDAA2E9MELVbeLa4VltWywmSW5DiuB09Ir/1y
Bh69FaItn3486NhePuXKQEa2XljJNEYa0L76bb75ENeZ6nVxWSoQODFxOdFyfh5j/EGQ17X2hHYk
EJpx5Nd1wX/NQtGHl9EKHjJqCVJrKIGwfJVjy9TcF7SXic3IoXZQ4eTr2WE9FkePJFHBqCtmNFG7
imig3tbx+s6jXxiXnYWUoYtXJ7GHMyT3GKcwT1eo5rYk1QpFAfYHH6tVw3GRRKjFd9M0UxmNxXkU
1enh6ip/+xEBuXXoqFb4eWXR+sLcxY9s+TyWseuXhl91eJ5ugs/m8sC9TPp+NqNrLFDzjbccwykl
10mtRelv1+Qnd+fau8NgX/pRTKKj9u1YFFiw01sY5FrdG7/p3j/VQRwDrlA2K0hMnztG3JbKrDjm
jrLBJq8jqIJ09ApkvkSwh00lEhUnUpDr7EVzSkuvjjHMliaL52S9Hhd2us86TPrMbFznBxy9t6XG
mhFObx9OL9Ztv380fAqNlkQfa8165+eZ27e6TyXK49zbR+SuF0/IylbAUD4+N/PWdRBHj2SayzuT
HLvPmTR+2ZP+2ap/L56P1/6mXJFDScoAKc1vHwgswYQesmC3Ngz6PVJm3UB5IappqTlj+kHkntrR
eGw3M15Wm+0pmJ8HQCPIfj79RtrLMBwGidqGd5HrF5hF3LtRNOQRuq589u/xI2cgMoLUGLWyHfOg
SiwTNZwr4LqVeCSAqdjQ0gHHgr1FKVtczay7zQ1P/8lCLeI2Rd9nGeFjy2oHM/urrQHGyCL6qd0p
3A6wS34sMESUZjpMVZQzKXbRWey9Z6Clz+OP615VfF2akdixXoHuB/d2gsJr3T4IsObKNGRRpf8I
IvpfaD3HLy7vCJMTKULKjY3X2o9m2ZHK2AOP//bj6s2p3MH3p5BTpguWvnA6jU4Qen0uhyprLoge
5na+zrCw149rVt7Q5P2RFf5p8tBKpZiSqyfs7a/lP6GOMlVnN/TOS9dYyo8dFQwd78ZGtXKteTq4
4EVbi925r9UxTMLHOEdN76O0jdN+8ehmwK5XRKxoODFW7WNFA8R23ct2wW79F1/5kNWTtJFcjNRn
NgOA1YpSQ8JptKVXF6KB6EqY2HjOkEmpEKS9hew0Feseb4T4/QDGPC6ehZrmSYV/DdOlfyGuoftw
tfowY4s9nqbLUCayd59OWv0QK7trJ6aIKC0Sfgepbu2SKObRj+gXy33IbV2N4rAiild2fSfVjpeA
RqTJC2xsviMf5prT4f4rEz8UN9yO6+04AwqBODdBpPMghnDtbdoNSSRDWzStBy9aRr7NcMUgvh4P
3WQj8CZLrQDd9QBeLbZZoQ7w+VKkezMH/0OTVwzfy4tytqXqvukTc1N71bBLGnLT5KvtUzf+Ui7l
aWfHXHvGsE/RA3Z9ZXgAsrbyBYHSIEAlHOMyFwbdeCae5OU+jWsR5wt/PYGRbiBJgE4oLnau0Wif
f/wVp/YGx8hj3VESHvz3MJ1sG8UdF9gFA6eZA0nX5l+67kWl/mRhCepxnE1RQg23M8IK/vO6QeLl
A8OyceQLG89NfCz1EdaBRbaUeuWB05/6Gj5zbGegjhH/J7O4mBq8M5Pq4OG5EJQPJhhLGB7lQeXg
5IgFWZMIwrtoIDCiHd04yOGac1isdEnhPST9Khr/5lwHOSppXnnVDzrFJNWauhKKOlmqcZkdqyBI
PNeeUh/lb7u4Tl+YqbuUF1ikBhUpDiixpAhszOKRMIxYXrpD95Y2VTL5qmWMFArG2xlm7pVp0Wa5
EG2xUD8+PVJP/jLTaaVMfsbhBdVsKZ0+tQ1ZOq2m5dRIBRoITCuftLCc1EnUlFisehWLl/3BMbHn
Ybj8XiSBwNs20RmcO5PqDQ0TE8EwUHpSUYIvv+Gix55mKmyiapfaqCLcZQn3GjwgnxOsU6ATJMFO
jwRXbukvZ5GiwRDrSlxwQhltvA2Jj2UBxRZ+hfSxAtBGbgPjspSS7ZJIGiG95Cn8qqHxgUbyIs/v
nFOmDsVCAkPXU874D4bijV7H7wDr+qzdRfKrJYZ3C+cgxPPYzBD+JEUXbY8D0UAGPhHrQk1+aEVf
6CFfizhRJsX3Nmym5CaOaWzy9mFKfnOXavb25FRPsH1f1bovA2LJ9o6X3AC5u2AnhtwD/oXNbvYv
oXkp1+Mnlk1dJWZgL4v3nXUE8WRdwppSLiK2DH95phxREqwQAVpU3TjALiYePRZSumBFz1VFZX67
V2tsP+C8WTXIWK3Vac1kFFC83KeaFHbHSUSDFy5teD8YG8HosoKOASCvBfxylGdAXPi6zfJyhoNz
8GJp02/qeGn1RzfH0adnOoV3VVEuNypdpjZoIu57xxmW8F2/FCnBWOAonnBr4/Ji4ltsttc+dJix
X/HavTVRzjP/zUwGCKwZHLCyuJ57KmSTw97dpPn+doBP0Tfsoon8nRxKyYU87SuTszKI52kdlAPH
e122d9CvI7MKkOmcsgcKxt7n6K63WlNlZPhmDm4THZ1JA9HDcLKBPYB7u+Zja88SrZz1Hi2qgCzT
O1rikX+RqKb4BBv7qLhj2p5rJHZRxZpBD5wKZSyO8x+Dv0PTetezVt0CQFnmtXsrMvwgYX6tjRgQ
+pa1k9miTjGSLkA3o6H9Pe83ohgCHx7FydBiK13vxxH7FEaKRJfTh0Ll4QWGXwNjdbp0s37gOMtc
8uJHqTO7iQ2oTQ5wPJ7Dt/0SyjMWvS7MqvhqPf0ChGGsgdOoZvmN7lanDjcEfxkpgdo3HDNpmDwy
oU3acmQY6g0/s4PZJasyhTKm/rd8U6AsF4Ne/ZYiuWyUhm5OIH+3VyH6KMfexD0v9f9xIVKLX4NJ
O9n+lFBwXRI++zz5XyTWFwWCNk988c9/wmb60rIRKwaPhDSrWDoHOPASB7lbHBCRMK0l/yoJePOp
Cj3eBBloZfpx8rfArvB7t+viZlDxvA2FVSFtwSxrMWMcBYbK9dUmqtrEQWvsM9N/Rbx68ysoTrDf
e5UXjqYkSWjNLC44hQ3znqHEw4HqWSFN32qYsovxGEk54rnYNQH3CBhMsQqJ8VYju8ARcmXuD4yy
cGh9q4FcFIfPtzpmB/8oDhy+nAS/is7dS5Ef/3awuk+WduInCToQsbS9BpXmGpkog0k8wlRX9GTu
woD1ZuXAaVAAuKiqsuWE/1n0/oqUjRpHFAFATdvrpkHpSZCe3P2/lFph/CET2YDPEl7y2xeJKzLH
aVw28fmOWfNyK6+GAG65ILV/Yh2O/V50RkFIp31PWCxSGBgjq8H5WZcKOFrRGj6WP6KWWP8o8jrG
6shfLyiNqqJYspDESuPIVkUNfNcOxj/3jrKjrNS33554irKMgs/u9n21HR+m4YcmDF1g7fK4rcMO
Ers+z0TCyjtnrOYg2+iLAxrjNoxAEyMhH/eqVegiWKgcLwT6Fpw4FWU7aILiIjEy03kzAnCKt+As
zfZBQcTHogrJt8slIH6Gm+SSFFqOoqdgeQmeeNYYP7DnOzHJUvannURkSc8TbhKs1bWOU7wddt00
cmiDiNS7yUKTojfwOprTMJEpaQR9gkgHMTOqnAevDsXUf9VRqaaW/Lg4FBPtmEn0WXFDhy6rXS57
F/QXfcZOhC2EgNFV49+VtRt5LEfLMjNxFKGcSuBahvFmeTt+jn6UZpKsor6c/UcFOWMvbo2cWWUs
MJEYjmNSKXerdi9NO+mt0M7UNJqbAXOB4TKYLcoVAl+CvvLamFIKfgezNoj68af5scne+KraI6as
aA0V8wc4D869r3hngh4RggFfIhxZ2jQBu549DMFgewvK9CrHG6foWGAytlwWcmGAkY6wZWSm66LU
1UayjGpnNww2o1/PcWmZQbKjkoJzpOqAqTAEyLWyxuseBAtsgWEjTdTMBuwAaw5wHyScM3VXoaxo
yzGa65syY0Px1H1L2p4UZzV3gBhvulepOOCjraZRhdUTLPSmzZpqRif/N8EGN9dV5luYfcjbrvFM
igqI3WfFFXhlyohh0eWg6Pjfpnqsz/AEuSQrSgh+F/PspP/6M9zXpfblHUJECccRYhGF8sWEsf7Y
k7QcTvbqwBr3Rrfl0zRFAEuyNYFlLAcfIAhi/h0Nuiz6xWLScYC6cTZu6ROEgfxGAY2t/zPh7+BT
KsTqJOyA2NmkSRKEe2YRugaObL6fSOAxe1Cd2XQhfK/wNJeDbKDJ5W2qQ9UTEnZsA5J6fcc/oQJ6
fEyEj+8by7RgSA5cwgSItEzHK2vGM5e4dHhAhynfomXHnFOWHwUUyjznm+q4OlGaI2/t1SkQIvMe
Wl1OxeeM8JejhUk+ErumEkfNcbRZeTTxmWfSeNnGk2ujQGMOaGW8kSFdJNk6qbgA5pTI2qTZ7iYt
ZKIcD+gnTXRrTWqIRM3Igg13ei8QvPrrR9/yzlJ2PFA3QXQiSbphXLwXgnn3cv6437xocGBcnk6U
o1mKFVDi+FwjzmooFVSbWMWVyrt7HfbSrEtG2mU+GojwZiqjCGsOYwDD+qFcVkZtMlho9es88FYF
zB7ihiFZ1wD9whhTelJyh88EPBvjLCdrydmXtXloUAzJNYETHvvLjyjxdoAQpo/4JdygH8u57JW4
6Y8mUq9h5E3hjzaP85ZUG2QNQ3cC+cJmHtEF0qPfMdgsRPVW8XO6ZeZGEFFxA5hM9KPIvNkXkE4v
ln6eO+uUkYkOrGXvy/gcqfGhar+ke1YoW1To27GOeeTSWbDQHFmYz/ropE6GgmT3CS2PvX4/s1cs
8wS2wQRkTUtzbuTEkF2KyewkuHTvHnSoe3Qai+QmLfKxs6pdrimHjA7nm2FCf2G7z4wvFC6mN4W4
IGJ2AjaMx9sgHVtbF95yEBDgY9DdEdpPoxo9fZVeBbH019u5gFDGTDEGkZNZGRN5Lx46rfXH9ylQ
dGNnczejFhwv/Ed6wZbmIrV+HpYxHC97pCPLyj3M4IWeGKnVM2kB4h2bEF67YBeO9eJAnofvRQsn
yBaEH/DcBIUyujMVvKgF7FKqUdML/H2YEKJbJJzRxNibmw3wWF7GksX+HmiAhLCr6rPp+N2oiLqe
2BTwoFSmU0inAvpMpxH1S/hkedBT1IXVt7dYJsWIAA3xifl0G7kJFZhUZemTrG/sx6rHXACPILWD
UuURUjPcpd8u43uzG9il7RoFnBHCgeOFs6OQlxMS0heRp2YOaPtus/jr5rUjip//GAPoFFVj7v3+
QgYFqZ0j4EV5bC4X+/WwPq9CvbHim56T10doedR38tFs4LNblJycwvA4JHc4MFT3Dd74jilKq7C7
51xfIr2yJiHLerBF0aSgCQOZx8rEZ/FCdzc1+MbdRX3I2HOMo8Z+XQfs250kW4FdwFveW1sS6yCX
7nWR7d1GeP2sGMazcD75JpSuRqHX8WAAqbmZ/8/rDJtbAYHC4HV4om0JokocUJBEtqGBGbO6GAvX
GynqUeHid3+4VmxqvqLP026LK+Z/hFfAXHq7pTcILN3iNyAzgajdNIlLeSyM1hlrIANmKkGKb20p
8weH7Pc1aXJ8OD7zPO1+y/TIeD/ERFH2A5Z/gkaoKxUPWZCZ2PRMoFYhQZIuHQT80jYngpWXv/lw
Ir+y9VZWVppbiLBBmK1mkn+NHTKigpwoyikTThaCcGAKzu+ek6If/q9U+kKQb3rPoB67fSOpgSPf
vo2BNUDs3epyINrygiNo3BYL5Y+s5RkhwMoB/IZRJRhSHKAik29k7qwSJxJu3STvxaC2inXJknMT
b5NnR89Gm1B7P1HNKvtTbFbO3TQivclUeRsqLmSubXilHw4v57Qazgs8hkxtJpQj6xsAWSc4MHjf
gRUu2ui5Rkar59Ino75JlxtpXix2JPGNKA9ovKZvRWo4samGUyMzxgyO57OEHLFTaOo6uIqbcfdE
CmOgZgE5lO/oR8CpzA0madWRkx3yK07FVxrD5f8I4E9GqiTQVJldfCHt4WZb/EAUhTq8qWFLWpiO
z8i5mlSt3dq/bw2jiOx7BYTeyHUJ//lf+3tSCchuVBr6ko3pWzbZlXJaolXFAiN0B79sBtWJGJnj
BR+QU8158kTMhFZWx5gNJ8nKCll6VSQxMEqU2j9/fDFU7q+fWu6dAScpX1hFxE+zFLFPHRbJFrS0
aaXP+6FxpOrniv9sY2G4GH34l9S+pCdIkRZncVPYZ45pdBZVpm3i6YlgkcjPisyxVVGiCYFtlGnz
1jixGOgFueg7XyzxXt+Z/HXGgCqozB41c4m1z5XdoMpVWY4SKjRq4HDyMR6MkZB7i7Yw5gqwb0CL
kBzRTXsSK4NzMB9UMjLCRcJgqaK+J+jkLsxxu7d1TxJAPL21zzofi3l+QWg2fkoXVQuyOi0d9SWY
H+SVdy0uc/IOkJQ5/5I/3UYUnCYc88+JXjDen8/eX9ncaidLNHlhk5BzE+KupW5lwuMLmnJ5+Xh0
g2x09EfOT9eZwgzwvfKlPFpUQ9MnnFhuTAXWTmZo6girhlfVJ3zg6V1KmKz6BU1TVD8Ant0DRIhI
N2buNzh+n1QyjRnz070KBMUNKN2QoNUXv3TzVmNvEPu6UBwTYybEb9so1NN5I4qmLby3Q0vni5PG
rZkjizGGxT5j4EmstZNMuktw9zZVODX/SjeJF9inPMYQBu1xHgs+DxQGR5Q4IZwzTPn7XMOMSOst
tYbfv3EtpYZrMY5ZP7QLvfqAjqgbQD94XwzBlgobYNDhy6OAWaIepeurm0rMRAeDYR8XY9Duy83+
YNIO6aAKTIrV9qmkJuJvpQlCEMRnYlYdpEoMcpUCjoy+wkHHF7WPaIlMPdJGfG3ENxZ6CC/AcHs1
n2IGdX5E61ME6h3GWf/bJ4IYkyKC4IctIdepGb45eDfJOd1Nu2efTGlU0PeDyRH+9koYZ5tn7Nz3
JXfasj5DMOLcHvgoovOII+mrBdTVkvHRasyU+EB85bMAmWRbU7Tkx+4fOnakobJrAxZJzyQNJe/Y
SzNkh4x8sBfkkRZ2YDx7o/5DLAGNUZpbAnh+6zIFRZE6+A8x+6/4/TTg0FQ5pe+nvb+sESYOtHWf
tfv6xRKBayUfaUtrx6FyiItLoAA011yVo0OUwonu+L8nPgKrkVwIyo3zlGcpuQgWRGolb0nwsPWL
32+QoBInQadIPjxK/dXOrnpR0jOkHe3hpNa5HfQb5g+mAOafvdtwzEOxNNz3iBqD82NkhXF6A7aM
LmLjUO9vUGL002aBLj6YLCBXJKCAdm6iEye1M8zoI/pAMri0XAdVLXr72hN9TRpmvAkq9AE3wU9n
bB3XM8o7MpJKNy5lcOdnvH2RlL1eLBfhjXeXXZU8w0z85a78sb0FoLXQs6IEiqyZE7kfTKjJkCM6
3k5/wqBSxCP12DX/w1l5hZdL8j76h3Y4XF6r9PeecYD6vzWSWrNK8AO6QpaeUYJhqBXgDPp1CMvW
owcSkRwEoG0yj1aI+LKHYnQPa4B+DGPLgkH5VnjkFBoxOqJAFdbQjh3/pxO9wsluXliwfWNc89HV
pIWG8ANYAES7EQJcP/dUsMW37msGncOOt61e1m0X+m5MWU/MlrDWq+mfdvhjhsQWGlH97ZhqGT8d
A6b8bVkdmO8zJ7+KEa39AMqYVRTKnZXFjy94JI+EUSrsbgq/1THhLLimrJyOJSgjwS5cxeFlXfYu
lzhmq5mcY+EQlOec+YCi2rEI/mZK526IePfmR1mSZxsYf/EvMs64K2yhVYTxQrc4ZyOj75X1ObP+
4QN9/7dVFKDOjg49IDifWeffOAQTzgdYVXgqwjx9MGvvOJ+I4+0j62j9iuNgtuUPUx0/JoWI7scU
cTt+pEhxaZDKoFOoC6YEu8S1kU7oPOx/iHwIItANi/RASKrVbuY5mgywoStqiDrd0gcI9JOMwvG/
8V26xyKtKhCuUozOGJDjDlHgo8T+fX49I+Rw8HrvorY26eo5x2KELtVa71ywTMTYmuPnRdE8Kj4q
MKH+1xS1d08RydhEilKCI0p08aRZpsP/xnP7xxoWf9RSrne8x8eNLjIpvtXj8S1h2UAj6cMIZs39
+9+9YJ3PxscGJmBxvxx/6RG1E+r8qYEsWRs9mix7vqAEZXVBfAyCLUoJAAxlLwAIBd5BcMQCyRS3
l9izZFbQryIMkgbHMCENIyV8YAAL0FohCuhZzzAA4Mn7vKZhO/p7vY9fXBhOs13Dk1LfC3LakBtK
PeAl9VEVJ3+G9xzm7KYMlEMfwEaK+96kOQfZ3gnpZmVLbWwY+RcsQPTvsBkGhOoqPFIiLX96CO0D
ahjiHnSE53wI/ulCSdOYBtWFeOE8o4VoAOF8ZNTS31/ZQuccwli2j+Sf4dUP60MNSgo2wI6hjlmH
JbGvVElJYuENO9waqKqEOwX+ntxUdXtXJbeiHBJ6W1X9gPuLc2m9qgA1jGTmdCfreLZxmjTiEo//
Y/Ce/QyE0KJVTHUPrko1OeJJ8vxmFLdE96oV9dG/OUDU39lz2/GosFvmNC2A1QIioKpz4XGlMNTL
H6VlazMOwS3e+ZMHjqbpcKRvVeCTWp7Laj4ohjGiotG1u5ujhyhjMBCr/rP33H7rikEu2nWbz8IH
+QZCZU07/A5VXOpyMNn8xP78YlvPDzkYfg/cFFls8DZynY+/jhMa7K//Ev2Eeb9n1LA5vUBYuSEe
jAYsNmPSVhLfS9PI5cB1TvzXiGaAH1NraZ/cwUTWwuyIS8sGq7j3XqfSglSP90BIvYtBg7tokadg
5Wg/X7KJffHIEf0L8oln+qk04/jMETMflcOZfLvzlxQxl7bFc8gBDikOIsLRxPR82sppDE8O9XFX
JMIrCoVRYFDiU0rWJj7c8KCuzaMD5t02Fb2btpGBzR5POdrfoNMpLQTC3pyTjZX79P+sTQI6c15I
xE3j2Prhwf0vY/LnAdh9NfgthDu/9dhSwu+z3+3he+a00XQecZqjxqPCwz6H2GVoVUHGts8yIrEe
rHZ8h0L7QhCqwrxFHHK41mLcpZRHTe5da0vdMvxwtpT5DpLHLPZ+It/qsWTDpXfC5lbdkMqGgxY2
XjXrkvzHCHpMbJynnYJ3l7wIbCGptDVggw0Na78z6081YIiLuUfsVOFDVio+xUE90YLr0wN+KX92
wYTUlYs2A9TJkIMz4HTPRwHHNZRq8GLx8k+R2EYJYP/bcyiQNQSKQjpfkXVvTCOsy/B9HBpQpWbK
gU2Bq6cMPfjwwHlXLIQKZW65MF74FJxL6+EAXTd6du96gwdHOOpC4d+1f5JBy3k8iluv+fNNmPsz
KaDgaasuK2iZ5mGZe+SUfWFyjxHidRp8OeDGGiOvSr+fwGNpHge5LstJ3NfxW7GtBqLg5pkDZUKQ
wx992W27RmDuWpLHn0xMljUzx5SN/E86oFGGjDzi9p0NJbXmg3CPZ+Mx63oQYvSmHvSnqm4e3Y3e
QMTETraH+W1DlBhG/UHJSqURjBP/Pn4PHLUwh1NM8nw2BsVW8lH26MriObfEvSD40zFvduwywI4M
/1Vq41UUbVTA7xzuUaLb9G+G87sEBPvbHW4ofJDKXio/e3CqF5p+wdXYDrUUAbFhnSqgLz58JyHs
97r5MPl9s423s0Q5jp+ZCMvlNS2ihVnyc0OKiR2HNNnu2jr0GikSAECglx6SfnJc5gkdRzv+IQtU
kLxeFum0Z1T0bPNU4EKx+wj4thXwaxD7DU7mmZu0zNbpS54NB8a6H4f/S6LjpqnHxiNGzYGVfJJ9
2YXX6FLd09u6+/gbbFihnQcSBCP+obTfn/UlKI9fT3HqwYc0++JejWtfpAKf71N5jsiza5x1b3GS
oZh9XhA5jeZiEw8nTvBNzkgDtIn2YCYuHWELAkvVIwGX3frbOjEn4pdabnRR+prLxV6uq5YdlbTv
Dq4Pswx3yJ2cT6zUd+JAqO1qb0tVgjgcElBjIO4gSVWRfG1xNydAOXyBBVBpmi1HZn0BqEkySnG9
wMJ5xU24ABATDFlqLLr06iAgFxateW4VyUc3342ePdrT9QeGSvZgtmx3bUxQz3A8s0EhjGqq5OgQ
8xw8uGkiho9Hwc+bPPYs48Cq5y+onsA6NuEPmJpjXF8UJSs3WObqCetyKgUzhcb9jSTCrHBjXNdI
C9dX4MCZ91mBU0FVseYI4vEhcFR+2lphuENI7tbs3n7DNpFhXieCeC1hyFc3a7dODre3J6aNeCm6
THQ/+2JI7X18sDkCwGUsSyptp0r8rajNvuSBSG86BELI5l7D5d3SQWqxGLBXqHZj2nAIadO0F3DE
l+bRWyQkQg7iwGAfmVdI6TX0WMPiDDHJ1jksK2HQ1ttWpcsP8gwpZfpkRzOZ6sXfLy08g7iFA7Wg
uuSyoRZAxJ73miezO87WbBGh2s1KKSs9ij1bBg4Zctozb/z2DpRYV1xOhfh83IQ4lWPbRT61Qax3
W+I4/w8bk3QVNOq3EFhUa75RD8E8F/8qIhdAuJdohp89tgnIIUGs1jKSqCe7SsERj0vSkej5GlEt
Qn1mjnOjfWG1++izUdIhlrhAS8KeceSbAjXe7oIOdNG3Y8Wwdv9H0KdzA2MSiG0AqLvXe2yS5SE4
UipHJ4qEPO8OHxGrMWxy0ChjmtgRCpL1RyyMk58JSnt/JfQyBuSY5eejSP80ycnFWnqkW3/CgCPB
8YaqXn3KrSiKsyieeA4+68vlYILnXxBF3gheGL7lrSYeS4mNyLkSgSGIr0MMoypz8vtdocxDA/pW
ZlA7ZkCH8YnrSyEGGIeXhAnzvvvmmvAoFupccFDvhXC8dw2upQ8aRyXXzIdvUzxeUNBLa6tHfuKz
CyC8e/4p4tduleUwCzn3BgdqifM1okH2KCMsnhIhSOmmRMwPnbxS7z65Wvtocf0/GFZN/RR4wJAP
sXpl81bA81Va4opHypwpHRuln2iVBkGIwGHTRXDlACFhbBgDdBvbsS/lKPDgv8aVmWra0fcH3dgt
0MzwpoFecIgivLQQ4FCR0M9nk9RfKsHZErfIKtpRVtGdPPQ5tX2Jk350fTbutwQcJQE4ghC6tZz7
sesxjLEkihaNme76ATJBBulzZaGP4PwZC0Qs9gLSEo2UaDl3776g5DNCD+qzObvnNqWB2CJ+i33I
8sqTPPlX5lUKaD9D+rwvi01HXvqWz30RcPhLB7dD/vaoh5ljvYmUKALHUf0gMayn+aT9N0iU8zJ5
TK1Oxgcc1khV76c0HWCPoVcTL5cUGxjgDF78MBkFL53gv5sd2ycLW9d5ZtJFYtv6XjwrLNKs15nW
FNy7qr8/wf7Da2HVfJC9t5Wbvww+Cce7yH7/7sZ3meVriscN/RBxIZVm6Id+EjPFROhhErohH29l
UccE/BSiWT3ZZxpvoKfSO8pMewBCNUU6kBjmCjsw2lX+V3WYjasMJmoRH/GKTj0Py2JVV6UV5Mco
HcUdPbmoh4rQaH6yVly5tXRNz91T04uVFpHfj2tZS3W5xzeMNVhGf5G+GFYEp6g7HbwKVBfR8QIL
87FnqzV/Y5vOYT8pN7fGtS0l2BZdRWWPJIoeW2CbqW4aJCTnZJqMyXVpYqyNYIRsN4H80ubaIcUW
M3nxNwsFPIB6odQ1axhkq0cHKKV2/S4mVA4cSIKOEnInuZv1nljSZIqSSlDRNAJWdyuKvBLKeeOU
+2Man/H8gF5S1dJZmnyxorQSJ9EFazhD/OoCsgpkumSnEG8SB2Kp8j0UC/fnvQyWrQR+9z5nAxDe
Cbr0I3aUD3y45bQl68WXnlv5a5R110IH77DvZiEeTwh+cZiABJnYJlgEsSA0LvjixvRNRsPj/M8+
zqIw6R/BmOhmX0poPU+27l8dZdcQ1gEFfE/AAEWWrzuMIcCC3aOs2zbYt7uzjw/dpZlgr4N1/Vvk
wkvoMUaI9CvIPoimvDeUtIKSyAu4e1j9MWBzZq0H8bioZP8ICmq5Q0+xLVGOJIe0rWnsgITD0vpe
ov8EIm8KE7REef5Bp0uJEOMBKnkCCVfSh1YD68xyrLqlwHGPvKPBjpaNnW+Xv7MwMjrUUz/4cCCN
nwzJoY73dk2Sqy2/FWF5x85JyECYIUV1SolVgVaHDnPY78SQGVNaHrIWWsYZKzjZ7NtLFnLI9F32
cpOFq4a9aBlpEh8L1N2Zvb/azv2+AOHRgC/HgTvjPqIBEO5SDw4A5gu3Gt222sxnXbtQESMv/TK/
D7AIs9mcPexvfEyFFkuBQhjH87hgCcjV2a2+7X4yfO0iXLDWFHpXcmbH4eT+7tLeQVXwKX0PnrKD
1caPpuE+/gR3WYylvSAilngq9ljIamFlOrdfqklFYf0PTszSQb53DPmi4d+zcUBIP12wfQD5jN6W
jQxNYLZjqHt8nT4L6yB6ui/YkeEEwFAc9Mr2KaPSicVNa6K33vi3bk8WxjMhfs+lRhuieDOOl4O7
qTYclGuPhnc2+DXZzmxs1XnYrBlj/YxowMG3AbpTOGSpkWA6aeBWRInJ4JDm0IT5vli+wpmUE7/z
Z+DZrCM1CpGjwaMAaQaVjAbcpS3vl4/HGl2a50yzbcGk3fI8GVNt6ysnKvyl3fkUCzXNTuozbGe5
pDqaCsT6jQacATtROvyn+FXb+5ENxZH7WQdc1iP2RZU+OWAG6WQvl3GDUP1hq5qmSYqHlxWlncOx
VldGKkoQY8MnLeDCsvVa3JeeKWxoKnWSZjQluFFCKYvXu6ZLoNt6Fd1Drt2nVU7FTQd9O1AH/Rg/
32bBP0zaAPUv29bik+GSPqvs8ypssY3D/IG9YRlyYaTlsei++e/f7U3BHoo9F59L8UExjGXmZ5S8
oW8j0uybqPW3T/HrKZRaVn1doSsVqCg8smu2lRpy14UCC5WhUzqy2ffNeYBeoTBa/h4DYniwNgcS
tG6Iy91ZNzo7nyBZUr5kX0fj4YIk+/pJR2MlXiSNuhloy1hVEh5vVX0EiHuovhMwJnqKtxlJlFVb
8Qk7nCt3wx/JNX0UkaXrl5SogjEQR7ZvBXFFzvc+W8JojJisDoT5Es/H9pBgOutX+g3hUXyET+YP
nhCj5kDZJ+Gp5Yvyj6eN6tz/JNM9B2CtHR90iX2GAo7tOGokLGEvCtm281PBgBIxT/OZrh3mnff1
gNF/knXDQlKD/7u4lLuEGXj+imboth3bLSKlG4p38CIZnwXW1lf6yr89KOcsvfQRtl8A+5vTYGHv
IpyLYhvVy2x4GVQ7CCQUo2CZVxrLQiKgeiV/BkAwuifKS+WP53rnaj3GuXNDFsJL8mm7gSQb9hRF
GLEIoHqS0lLlTQ0prSKG0sCDl+JnewGFyKb6SitPv+yNpiHXZxRxSBXDR9niytumZi5iyriQCUDX
79i8PEaoQaO9rd1m9FnfB4sJoJu3YwNlNtXXddSrsRnjvdKXi4xT/YgkaoU7XYF7Smz98NrsSaKc
AK2dZN0xdeFW9H1g0nd8K3VN92OajIZ20Pd1VPRAlLWzfou/muZFpvKXNXXXM7z6QfvA3983FTIy
U5ft3oKKM8XjHCVQbVf7DkKLFZRT8HDNDY476KW87DplKFyXn7ZKg4rDqj2SgnqAx4AHGw21vPoL
ZRt+4aZICvU408uj0jVuYfZi1R4suR0q9zHVFKAAS//GYfQXJw4HXSiUk3SZN5WRah8UKkzUJ9Tb
Q91RUtxjElM9SyoFcYKL6wuK+d8Zt93qZ/KQEzZmheeC0wX7RN4itedu3xwX2EzLEfAD6TzSivXO
KizMLeLG0qHzVepWykEb2ohS6iKicQ8NNah24A4mPUoQUHUkYq3psgRvnXe4CfISVsys6v6zfsXf
Nh7cAAuwQaYfvzgCH3uXpU2fAehtsQ42M1yika95DVmzkxvT+duH7cRnN0MnKlPnymOcKwAxPEAC
ZAlw0oXIbHZlN0zYjc0eO94/4uV90j29VNpaUiR32ipSW/ZjBri1ekY6qZaeZOuu1JgYra018Jj7
kuvYBp2LBHsbVRJ9PvYxtVmbSBx6z1oiimQkzYxoBYAdl1LABMAxdf1ZpHXgb+oSk+7kjsFILmFD
PVXPSpJKCKSPUjdqyx4vvChkjbWINSyJSwjpjaea3kMqRxKkd/Fq9Xzs2vTbPdBYvIqD44f3aMEJ
L71xgc2FkUc+dAzFG8vPsfaMtRLSJ5Ua8G/+MVVCbAeCqf0rXPvKAl5QlwiYhmcPmAC9cebdFyF1
Arcn9butuQoM68USYKZw4+5Yt6Igna5o32gQI0pTYQGsUDWEwxDLO7MiEwVir9zrl/ZrbGb2ZCWu
MVl9oVyjLZGx65Lx/Y+02YwgMDPUEW95EbOWs2IfEKx/xDVb3MIJqgjHZLWJth29PQeNTNJirB9U
QL5EVd8a81wug2sIKNlAr5+NBvGtlqU4noh82rXVm0genV1Hzx4RhDmKDUTN8maAmRgN/k5sK5mC
Yd5BxNrKBvsGU4I7j9w01uRLXCPLuPBxn3xSQ9NkvIjYTEU+0vYkX8VzNTv0OnYqVFBRNuVV2aNI
oE77AasY4RfZ4pgVnfdoTkmjS/pMSW4RtllMUgb7S39ZdOJRjnMrfS3YLPrgbSWpe097/cAvquyC
C+BL7NwAuzhvXve64YERqSKFZGluA24KmAFS0lc+h2ZhbhhZFSDWTEYYEYXUdPVLKtubIoCLJ9LW
CBothgDsfTmzfXK6c5N2JxhnSzVSJczN7zioCQ2s6d++nHeKzAeK3S/b/brlbxhUjexel/j+zhr/
/fEtsgUCyMzPOnhy1K/ZmFnaBoenXhay9Coj6VuqrJ1SF7xE+Wx1dRpoKS6wVdr2uIrHyQJLfn1T
SLeII+jQ9/rfUaO+yJkkGNxkQIrRkkbI4Zk+DQD9qgrTCRLAgQZKlxOW3I7UgvwyH4iAyvQ+smlT
gE+g9s9JTNVt708Bt/Jz6bXGDCIisGA0mjGGGYst1OOfIaChxYJWvJjqKVEw3oTQQdag777ambuT
8DxHSODiQvDS5eo7eJ+yX3rD3vm+FxLyj/Czy08pPqtS3DI2Z7pGH1+ufCkmTmizDjaJXykClmdq
GrRr3oIpFSStox0RDb6rfnM0tdb4xkLv9UJSOQJQBhyZPHgkFXs+M+xN+Rj78sJ8+EuYdkZb8MJp
3MNSh9SMnP90rWbjWISy+/cNoiX1N1Mf7eqoUeiBqIDKVj1EhtVx/NLSyxd++PYL0lx/xtFCYC+R
RtfEAsUaL6dJGrED1xxJxRFXeS/IE2JaeW88lIKYpnxe0jU9Etjj3hFfPnLTUjbhkanaZnDJ2pih
ACEaOp6UNh5eZd2VrMlNL5Eg9nEMqguTD8EqpY33EEMFjHOcPDl7jGxqIyIgyQ9CapOTvOURmDe0
MpCHv/klVLyzFhbq3WM0ZSyX5QEqyBtMY6t0/S8g0QGDFxgfXexH8gqyme98iqUudY6c1uAnl2yj
9UWBAfMNKwAXGCVMB8tbVYYo5XdmcNOJHsIJVM+gctAJlYpnhhw1sFcMU3nC8jf170uWCReolfun
Srsa30CbguqjEOuCI04kcUgCpwQsUrDSFvg9rV95WJKvO2MYNe7kqBujaNUKFAx0dzOxgc09bCBa
XhDn2YJb9FS9cP/+1p8lVc9gXZL7vTjxAF8wRk6CGTWUoA73MMWvnD70AzQapmXLeyYKL+Lp99jl
ewxV5vcrBp6L3hWDhRqnBlZZi2ZLklJ2gtsp/QDo2oLc3E/NXYs32dte0iu69LLpioZ1coWPYrOM
ZdnKV3i5qqkDQH9b+YQcHOCTs0s2wBjvD/cCN8tkfBmpcW9+GOWDzenvt9zS015fcilvI7/RHLYi
BnPAjGkYsoea1WL22T2P/hc03bM1ESC9N7hbDrdzjKSqHwOosmX135VAkd0KnCDmY2vhYAk68guv
HIgLpkvKoBVjPiiPoajWB2cCflL4jsVwZw1WVIjZwIMQXZMtZH2H0xzA20rx/PJ/+rWueYz7CtR+
+7BwqjCeE7UEcr0oIQpAUWb9vaz1Lg18aAqgy6oCZ/2x1Cb6gp4BPkjhXLvEUsNAfolFm9ZjpGHb
RWPxj242boZM7+LRun9OpUpRLYheH/xEFsm5LieK3xTRG91++LV21bZg99ASqdEg/kyKKigoXdbR
KwJWXGo3Q+2q4tHzgqFWtEb9I4Q6PQ1U6MPoWc+ObgLp39QM12vfUfrdg9HcIvTF7pnt6jdYtJMt
EPsbk/LQv7eZiFbx49/cN/tSuaqTwuqf92JugZhMMDNb6J1bzYcgxirRBZOU8O4k1N5/P3W2/Abn
qUALyFiHLuG5EWesZTit22S3Flr1a5XoKo2cQB1cS2Uhsc25y8RGwzgzqPPEGeyd2rHdv4q7LtRG
GcGP4bRVe0P8UV3o5k0AzfOEofgtB7TcnjXb9HSfB1e5sTnZrnHL7dTGq+oXwCPIIedNyzAnAUsS
AU6gVFGlIiJgDTWDXYyotwwAaYg3hRfMMaV+bzdgz1LWdlxHbtkdwNNWsub9OtuBdX3QTneqJn2v
VDZ7Tjj+vZ6umjp6tPNUdKD1bOujbqC+cK5BpXR089T5uoccWuECWhnzHwTvlfUEHfEUi3BNFvrL
xl1YsthMf520OJWcra/giZfrQ7qc9zFW5qZc69UGV2Kf9XX2FmcVaasONaANxaa2WdOvpsLIjStx
yebSnfBoIes0gtNeEk9ok81pfGNHCvVo1xgtJ4jn6y5WawZLNhsqMusno0F2ZqzyDmBVHxtCe0Cl
kfpU1p2uOOXSWamolAYrUid02sNBkGa27h94uWHinXflDbt6IP3Ha21Ozj1tu1FRquvSSqUHCI6G
gMAYiQpe1fvpVPtfi5FiqKIuMnc8Q14QjMSVNcnR//R7avD+y2dTfdedDgxsrHY7XGRHcXKft0Mx
NqtXdw2CbQM3rEtB6+HKgwLW/pRue83kk2sKAf2NFbbI4CzwgQv2Ab2E7/zU0+rAQLtGjGXphA69
2pJhwimH6JBVmlqOGalogJYZ5BIL26Kg6hBR2Nef3Q3Pn7bzrpYcnRZf1HmoaxQf7wQJactts/vK
QHxXfuQ+CmHzpSdMskcm4lLgZgCa38w0oKz8/vzoIlwkx/t5essv68AfOPbUua3/7BZoTXDlY/Jw
pWjXvnIcsZ3ROGuHN3jpCuStBVkh/IQu8AXRspSlFLlyijflGFYvscx+TaXZJnFLJH0JmAVTZuod
+oY0hLkxohgqDkDpchogiWkkuTQpI2arzICWSBlkwQd4txzThDzOXI3CxUgEsSrDhKU9v4f2ZIsx
HhwDpojoE3cE0FnbEGtia9rd0bOYQvkoJcEd66oyMJ+MfdfPLg+EkFQ83A2oMSC4iyU7kvC9Boix
yl5LVQKV5/rOgG92D2ZNTDZ5Op/NOhFnNT04zAoPASGhVf8MxA7rY1SxSRqSaborO29crDrJ6Y+K
wlcRtxL2/aSJHC68eNF0FdSguNvXTolBywlioeUXalWs3UZTXCteUWlCegn2gYBb7I+5nW7bBx3M
2bZqDTX+AtWhDJOourFbSSD9R0CFUvLsuOl3WczKyZzmLpvxq7JrWURmCav0JYBi7H2jvuS23sJu
7pKL/FTzWMzZ7fD9uyJCzIKQBrGp5bz7l1KuKHV5lCQyDj5CBXdRNzKdXMCJ6B+ziyuuzJJBKYEh
9m9TMCqioXJylT+MmAorTyKbivWYOflXTNmrVBPHiSOXhvblSAt2uhlUrKUHR2DAT8bRvXsLfDEA
XTjcED/dONk1tPJGU+/COJkx8SoY54F3K6p0OBIycxhNevV6mgOifAKYSlsP0bTkPZk8WQ7KkoEg
kVqGouzS2n4LE7sgu1fWCQaDxE4RVMiOhmRDwkSxgzC02DAk6qMokRchCbqUj/0oPL1E/rtM8/is
WsbaqsMHfD5SO8DFNpJ6V7BSSnNv6uOAL5g+Wl0sYPqtBRGD7Z24yY5HZpWNfmGyLvMJqWJFqh09
mAfyUDG8YsXWT2TFnq6XLE2j+w8e9YAsxCzVwagydNqHWVLdHjr0sn1TS4LxZUjw2JHWaONzZN7c
ONaJsv5h8sS7JSt6PfwUxbDdiLhOONuwOgvGv1DPP7z0wl1lBJct3CGBZ0WjSmtDfxx9U/RjdFRW
cnIkvwhh1p9LfH4KgE88/xBrsH4i2xsCpwKYvAc/ycr2HSvYlSYIhK4PglREbs1KNJhIhpQ2LWOX
6FhkPocLVejVhgBb6OJK+KSXzQK0fdaBrj0iYr3XNFCuIvvM9fJZuj3TtktzqFgMIotB2CwkE5Jh
oWeWP4q/gRLo2NY+qTboFJT0lsKKDlJox58ehNvxaE+u6mXRLgAtqN/Ipj4cSDbvU2GbCEAYGK7+
fFv6ixegmas8Jx7m4rbzrbZt/4HFUoDxvm5F+cZ7KYo+1x7dP1EvRdBg3XtJ5Dwy3d55NEulabFI
4Dm4oH5kZTVHirdEIdfM+kMy4UNubR6rM4mkcMCQQkaV7wDNvjQpnymRU2hS4DlTpGr3HoSyu2xn
BPZaX/M56Hi6Hidj8DAZhb9v+Rsx2IpZ4PPcfBcvvsT7bI0ZbbJu2lW162hmVMOl1UW7ly47OMX6
q/O6AxmNg3WulB/x5iUmBU/GJ8uhiq2IIA72Zi5ZmtezyJWbY1yuLbkTSJ+GDJCveGFpXDwPGUnb
ohjxOr7tWEBtT2acGdb3aFQ6xVZpJwD+vrRlqJgkbw39oPXMPxY0+nwdX4DTG/T8nHVtFkKj6hxp
E6tr9MHWm2/HXxibSKcJPZOGHmqdkGi6nS/CaQyfAwjBci+zUVVu6OU4tC8e4N3sXdJqUExXbNib
wZ48hUUF0oKz/L/pJ4H7iS8FDTMi6KMdGhBPyldk/fRzmTB3Yff1O8eka69nwbYQSOr/cJKW7zom
3b/Om5EggIfKw4Atsj6RGrmLBSSdW1agjVBTzY6NULpN/b7xkLbyGb/FKAJP9E5Y+JTnkEp47/Bg
3blB4iUTm4E6fN4qPcg3DBvoAf9/+uKkuP0Boz9N5SJIN3nQdYpGCWpkWpBz5UVCDwDecMkpiMkQ
FXgRHkmmWx99WkqJ1dJWbcKLxIIBWAGxW2Z+Dbsc2iivMIqAG27tQB+0Jkhu8v9p6Yz0wSpuhxgV
BbvzO5o0iMLHzK4TlOg5zTJpTix6ohESzM0zDCg0aYng9uGRjqd0J6KZ9nTZxnB0t7zTkqYRyKvJ
JHhXnz1xpFdNWrslg5hBEJzqNBt58muPRu38oja90VPz9iiGMU76omrLH2bwM34WTyV8PLz8UfwR
Wt6a2/FojeM0rnCUnbUG6dwUVtbF1n2TbuE6BBjDDZvfXkO5QjUCrs6aylr+nz4CbSLSFYjtc4gw
Vpgw7ESde4xVnBemF+F3+fkOjahSRxKPjMIor6dhrZlH4qiu6vap+HYmvtfUMZr+NRzf1Dfl/Jqf
V1PgYHH4eSV4tRuYUiDME1BQNczG7ze7n9p998f0P64qqIyRd+2ThajA9VS5Tutw0M2XR4vSnbfZ
jTjbvXN1KckbiH3Yh+mNkKbsgR45+U+YZyzWoAFkfVrGB9Xk4rOYm3g4EmlAvYkli5UrWWNc4dX8
LjCjpo3XTNyva59X35znTlU3/gZwlJi88Du+2wt/0Swg5+vrUByOmQ8VI0kkaDet75yHCi3kJ8Yb
HvaIwNA758St6xtCPeLgxNpLXW3kYXzZArAdoB3vJwxst6pMEDJ8l9EGuWhkTQBom++8rCwBTSL+
1T9PWV5IzYcipggG/FRpMa8Y8JBXQn+Ap6uUvdNNqd2R7xy7pCkvr4MGure0uLdosSBOq/T9Wjx1
YR1nkbk+TbXvfrUMYtPbVtDa24eVy3hIzuXDoXMuB6Rya/jaL8T+Yj1kPqTjZ7V99hCg4cL81apj
8/QOeh/IVh6r9BKvE0+WT8vkhALTRlmuX/femj9TaDJ5pNCcxW8lUGEvyvkS5xRnuMth4UnRMlY9
Vg4Fb0LO2vjx9VoYRYSn3wE2ihOoJXm952pgX33G4jp6dV0to4yecz+rg31QV07yHQu2bKuqZmn9
TVf/dwcYpg5WV+G5okGsuflimGKkAocbDZhV6ah8DM112ZJt5JBbMWBFde+44JLtkbYro6r0cMPe
hQdQgCviR3afZhZ4WeHzArhdJbbQalgCyWqmbd3SS3/nTBvibrBLfQqwCtNUr6jLFbxdvGbjr+KK
oQURAGuGC5/ham14ndz4GA5UoHGyniTBR6aTaBEbZkx7tSOpy1ufxnOtt27Z/VRp1IaH7YLfNm98
jWq8S6VSqrXU7kAapRks87mYu4yLbT6nvHdkSP0C/xm9Xxiy5g8PR/AG74PaOtRjNU1AV17pmmA7
gxEPtCbnJ/ZGGRIwYqhAuzEoOLPgPX0XkRDJ2+GsRPZwM13lj+SnJqZ9dUSKkzEbN3KJSI/NJWnG
BVodE0A3tE6bVRq53azbkT7ofVrEROcF2DUmKa35a0YvNi/k/VPMjl3MVxbG6AUOtTeV4BLW12YF
otnFmh+TiLASdQLb1cKZ1/yPKYIcdSWCUeHOUxJDKWnjSJS/vNPECK2D1a8y5340C0HyOZ65s6HB
AeAbZaDMvYA7gCh4QezKDqrq+vP4fZVH5PcieY6MbxWEQ6k8gPexil8zSjz9eYo4iImZPYgeKyz7
5n6KKPQLxxD5OBG002WSXTphQeIgrhooJQwzPAANqD0PdV2XxW5aBtLicX57LjxQy3nEj8SJL4Wn
Px75qRKWt7VoTiRBi7BaP6nPtJgVwdBMMkqvg0c5d679Ka8tXbex54jn1Ie8ytZkQq6x+FPUuMPz
lGZFlMV43FgS2lCc/RYNanKci1MCMfhSrnP7/ddGn8tZVYIXqDvjjQFGtCUDBiEaPyDThv0cLnmz
agsbpfXdsGP8yLDHBQlVvTJk5z/0bDBjBK6YoBVU/U1O9DjwPjRWFVAVK8YG70zK0tFBm+irf4u8
C+PLCwCUJ0sAT7O5J0uvoyvqCkzlvvJhEfq++KfJfsBW4cyEWtr3QK0VL3GRSnA2dXYytGuAdsWS
OjrTuLvLHxuHogBZ7EhO6wtrWtL34qEw3s0C4pVuIefpmPo3YEssDvSo/QDwJqY6E/IfVk0sK6cc
ZH3lnHQ15ugTU+9vx5z0S6oJWAjjqXUOJdId0GIsCNdIyJHgVVlBLZei+aIELUdIJcxY7Ifpo43y
2broEY00kZ3qJBOusDib+jpRe5J1Kl2JQGzO01sC16r3E3MhSpOpo25i3ibuAZ4kVEeQ6zjJMdUm
FFyTvOdf7Uh5JQauQb+jOZZPGBtMKB1EWoXNrgXZta5yOFfFghjpMaTkhrpDkxj6GwE78J5yktUw
dnmln89EyIKhIfmfu36y7fDxYkYK8j32XIqCq2CDXGc6G0ebKY0tMSZFDuuT/zUWsOTQjmjaGUxW
qdWIuZNuitBYoLCOxlHbjjn46lm5otDLmCUi7Dzfqdvkz69Ec4MdpsX1Eda1jPkzPviW469hIMlF
GxuH/HAtShBUyaR2VR6G2gG59M9MSqwp5eclV7bsiOX60HndXLC1j/xsAVlQ3hzWg5NzicZXTrS4
VVz7wTWePnNUvLtXDU6zMzl2LwtgFZH6adSDxwpesK9kl2kwntZdkcjML8FXQez8FZFFa+a2P3aw
TGQYqGcuxXQ4pyuoXgTC8gEzbuiue2B+8WFpt77sX+HZWvYzR1lVyOiKunPFA8eHQEdfi1ojWx0m
vcdC8tfUoKf540T7cpiRg2eR9dFS4umyWPu7FfAGoAUEgdyYPHF9HR5onQX3kat/pXWXXpXVbDWj
DSPqtOFWDpamK6pFeHsttVHyXDTrN8CFUwxBJRTDlIszJAOPw49O1Y7YVX78fJcK1ti2rbRDXljc
DRuaDzqLoZ3fdx9fTBx5uQJxSx7BewpKgvN3BfSQrQrY8foNHTLpebDKZbftvcMHZvF638uIaZVw
l5A7YzwOJp4yJ8LDeWuhva4rc0lB/PjdTj1LYaNutySfmQ/UGcHtsHlnVsWn1j20aTuNmILyJpFI
7NquxC/gPE5ijsHFmQ8/zZlTvAQpYobTnkzNfjOfuyAcbY4ZROsPQdEm7nl1lfOUlEUUKlq3TPN7
Ju+8+mNas5+GVOpyEMo0/Y2pMJhZETUWfplpsUQ8k17yiX9VQt59IbVjq0fT6+zTt5qyE9CbS92E
umaw0zpno+IbvK2yC1BOCakfA4EkXE4TDpoq60Tl9llm2DQHI/O2oZdZ8MCDjkOKs25lzvxinHh4
LvdYoS+/0dWFxFYmXHGc+oRbjfVNlrAt06RfLCeysGygLWF1/oSBzLOxc45uJ1VqaEW/gECBrJFw
XRZMH66b5E3BTfJU0afmoq2pSzKwiozxO6EQKpziDZBuOekxitAGfhIBInmjyTvvAvzk86DkTU5Q
Y4OCBrtklVO5O/NLHllnrLOshlaBMspqt7Op5iVu2oSVECMMxFepGwMG/7muHMc9wUXvhUkQJd/4
ipB+YN8wzk1iJhcry1gC2aivu3ZGzj3ULjciQQMLoV4hEOLCRP/WAuL8dNYBUGq6MWWm7QUqS68V
F9tM/lF3IPo+MHbZXwoRmi7bieLGBJorDj0tKxARStTsDdXK7xQaecqdPt2w1cq6oNq3EJstESnj
0P6Me55urgcTon3YNsDMj8zR2qPp3aj5tX6eE2/whTiXq/fmt4yIVkYTUfdY+mSSDk9q1orptT4u
FWmiByb5fpThL/ZHqPxLKp9qjcEzUY0CXMha7KUYhg7Erha97v6xjufZNP57pFx5uG3GBealVdJH
P6s0tyJ9OVWjegvY1lOaWhfnJ01ElbJtQeJEP6csdrmjPtBShdFV/uK0qJtzdXM+spQuPZnY0TEf
HcdpST3gRrd3WIB8hkfdXePaamuLMcuK3UYIeBVU3eexIwdJ3J4l7VCJA5C7vNlGVY0yQ+tuTAL6
PwCaX7krs+w+ZuczyZtLQ4K5D3W2nY+kgrP9B7XtlNyBv7h0QtfeB9OYPri/83wCHKJCwiGrMXG5
/Fp+WRUCqwxFnCEeo500Ct9G6dVd8JQ6Jmdf2aTNw2DVUqGF1YAoz9QA7jIfhpBVu0immBWTv2HM
m0RqdG8Nd+atLFTT6p+jaGuc45gkwIAHHwwutv5VtfixDvgL0jn6c4fVcgL68ETnXFnaLe+3Hcu8
FTSvKpcidlVeF/ztrhv0qvqhG2zO+vZWVFhJicTE5RXkfkexVMG7/6yWCwcO3aOgE8MvJCXImh/J
G5FwvGTIr5w1uVmqky79KX5rg19mJ3qOYJWVslCLiHrDUSR4c/WgWq4k8ODABjxYmoytXlWxlCTL
HmS4e5S6mAr/8FcQ6Wxarzk1cxBoyVrh9N83P2Lscvqwrj/C6NuKG7wJJZuO22p109gf9jvGa1Yl
89R097xFVCBmK/vFYpb8baOixLE6oyaEgWBN5Qhk8Ld3MIr+/lq7ZCM5V8g0zbJxfal/qv0iQWg2
cRxs+5J8oY7OF1bM8NgaVxQvfPCckb0qZXN0NghVZL05N3SkFvjN+1hTHJmpHbLFEZDg034AX79X
ru8lLNzdim42EqgQidwJj1MSe4TpsN3RSkV2+EVxKvKnTM3ALDyydNswowIP4dYrRctaGfuCyiAO
mgB9WLV5VUVrkBr3SCiyPv4gmnpYLW443UUXkEXGro4ma4/YDU9UPF5aYFuzbeWzbpyk3YEmERCv
HlS5GHKYPo/Xv0a722XcKPBEiwOtUUWhHT8siPlgE9zlOYDUdZkp+/ZmWYiuAusnIsrnTUQSvfSs
qJkA5gcUCWuG08OtlagWluTdbgRSJHpywURb2NBbBFbGBtZqXBb9R5bXByTxEgdkbwYF6Dn6Ugvt
aL8y6msPV4JbLx5S/4cWnCAhQq8rpAURdVu8YWn4gK/5W61nAljG0ODZ3l9LsJPemOiw70CCj6DU
v+IAqRrk/+zdAD1gX4dv6AI2dICoa7OFn/rOqHM9jCGBTeKMZx5rJ/26QgRrCTZaP3NqDud2uJA3
LJvLEuiFOh80qgj5TgBRtdGy5GQHc45ViP/eC0hcmMqXh+KR8cvFMbWceDnKqnq9iKozBSmbIvjV
NlLOnyWqHkH+TAtd+VVDlwjcV8rHKTcDxeU3WzSHpYe4apjH7KaY3lTmJQzTeefhxMm/D8SeLB00
dFXWQsLNZGQJstoI9vD/nodwxja1wvK2nr8fXyUdDvcj8ykoqqGCu9H4BJsG3RIWSC8pNGTivXtW
HANZoctPIiHbVCAaer1LHU2qcsy7MrmGiSM/Ja/4uo0MUoa36qfEP+jjXBHbpfC6aKni2fcbkMOy
F5lTInQXXXB0JnBlGSxQInHw9YJbYXCBn8cXjpW4GfAXm6h6GahF3NHZeHAAOOgcx4kNTukpyHYD
O/bJJWJw1NllHctzLFf0xdZuNt9YOq1GxzyrU4afy9hEwxHKmxjJ96vkuyDbtuB2ivv9T7H9nBIb
Htek1T4lQxJfU3wyt23QMy+7ssYkft1QkVw/S3HJD/mQmEEQRYHkybbyvkwVH5D0RzIYQseaZRsg
WGtVywO/FRBLrUebnN0MRRZ6RSjE4IBM4U4UkrPNfRNSFrKppYz2ZlR/6C3zXTtJaP25s6yNQ5XE
OIGjjVQGqd7aF/THWbOy6v66Wlmx5hpwtr4pWT9bvLs2oYgrPJ85b2s8Mz/wRmBgCbNvme04yIPF
JBc4Tm1xYK1501m/7OhcnAYyDFRla9soFX5dz8AiVYzxAWmZo19Gqnqa5TXoXbL6rE5HereyWj6B
dxzPlvzo1JJefiaUGD/y2lo5GvoW0TN0HYvbB76TF59koArrgyF06SNO54Uz2JCL+4E7dWar0DaZ
GlLPSNFjVvxS20IwSCZrgubRXunjrWQB0qp2QyCz9aJhAvTHUVLZw7oEq4xWS26xnR+/M9FNxruZ
tOJrRsd+ehVYGzVh8Huvs+fArWp+IGlEwDOM/K1kN9V1fcU5SCdEW6v+PRLNrUUKYckizsdkRPpQ
YCVZjucXw8NKS+gSxoF17OaFm0h6Ydzv3JAvNXG409bCHJHUjz2MhuYcG6gn3hJ5hpmlmU3Idm8F
vECjIXI4yCQaeQGa+N2UM282tRRvqt2bfbrTpHk8iXt2kD2sshvgiTrsBEcQ/9BclIFTAAP/dlkH
kSZ/vmw9nej1MpvAJr6OW4GjlQJ+JjGVS19giJ/4wCUQ933AXUcl7yt69pxURZiwnlT41HAjGVbt
GWpab3inrHVSlBhABNIimWanSkJ6qIg8EMtljOkrPpyTD5rl8uENAVvA07Q+aOHwIr+T63dGafrM
pcTcc+GpTCShOlIIRxJh2TM12qK84d/KViYQ6wc1/4gq8XK+ryLGHcc0Nq3Z0VnibFjYsKuxoijE
iVL8oJ2rK7jgseElBpwuyi9muYW2vkePgnAkW3PxfaEJP9irxb+Beve6a3yEI2h96FXowftcKtri
/sy2/TjdW5khmb+xIPa+AGG5KHP98kHQQ+LND9pzd4w2vry1a8/2sLxEEGVb/Q4vmy+Thb53E2du
QtHHRo+Oi7GK6baC43WVLuSrrE5o0Zgc84rmBz5sLKahLEgEZstotAK2+AIfpnc8u3qxZep5ZZ7C
3cSTJLJagZ7IN6CxDZ50jfS0YvR0AZKC/H+ovAwARqJ8UmBK68/tCPAMw3BIRvLC3Y5P5DsSaRR3
Ed9KnFhKnzaRE9Y0MzbRobtj76WCDu02gCgBcYW2h0/Y0mQ/8vXIaUmkPFOdnlyrgJamleIcxClN
IO6kwLNy4ewr71PxiXQ0kG1DrBUAE5xhmj9Px4eSqhLqAUelUdTUL/rKHwNFA0D9F5kjOTaokifs
pL8LTtLVSnLocTHytycPqU7InOm3YwosMWCo9DtuB/IyB4VZsPnW6QVp+O+ah+LdIID6rAytEBgT
204sbSNdGv5GcBS1CTbNlR5gQqGfbIe5Pzc7bEwww4ycYWe35d4ayT+00Rg9kSJSAcw29PWYgyU6
dLZPlqgo1rQtTZGbtivsFJFEnasAv4WlenScsIZja902fwEv/IO0enjTwDNgoIN9wD8KBLH1tZvu
d4Plmyn/1vpt6kjpAFeAW77IFFJpWGpeyZIkOWFQTaj3lL5WQfJGqCeEWg7J9z/iD2o/WLrIQKVq
vMWboOnMbm97ALx6rzJjsxGHG+W2c3mofPh/H49cAEarfnvCfsxF0rJWhQjgtNigeHLLEzM0YTWi
66QvdND44dIQqwvgsZnqNZq8PpglL3JiDmA0RK/hrTGLxiNq8jeXz7vvd8/styHjFbSV2050wZBk
Q1NeE85mELd+RQn2yQ/1XGotceJ2OGnlM4ecY/EjXLZuJXs84Ml1qm6zue6HawIIjGIQw57Ah+/4
Ge1jvlPx5afB8okmT6VjSZt9W4ULk3YUSfKy93qFV1tO4JCI6xDapVRImbCEO83sqbFMluaWsvOn
zXHaMBtsHxNpq4o4+hEc9ceAW8TbNJNRrjcAkdxHqocJaZhKGlEXPl8uY5AWFajzZLf3SBt+lsl9
Y69aULOPvmG+cUW6JewkPY5RqWWgb+uXUPEAjWkgLtPfHenlImOphprOv/mfYOcY70kRbbiCl6tH
asDv1YqmyqB4CXV8Q0cAemWQ/8c8LCajEpHbU4IMIsWjHUoEisY+wwgHLrk197TxJEeUvkCvJOA0
UCPsGvRyytKID2D2krHoNAnCYpZK9I4CgRpbvnR19BW3fNr3dZ1M/YsTB+/9gyITNMwpqqwpXYr/
ORmdsEwP/IRv42pTpm7hTLlO+UhYbRQfQ0rFsM20IuLYW/0HynBCJ33KMFSDV3OsHeKNenXxC/Fh
9GGY6EfF1Md3nPUgM9K3dzRLbaRvXGdFGJNZoYke/1m/ub6XU507hncvH3gTWa1bDUuuTJdVvW0F
YZa7cFmEaNd9D2waUW79zWnfQ+YkL0B96xXwogRND+HNmN7LMPnKvTTGSlRgaRXVg/n+5zlxv05Z
saS16lgs2pkG4Vs4+yxGx0OQHmTIXA7Mjj3t/vCSKBjWFySL+CuA/UPIpanfscefgG+KeJuGOYfi
/GGwO9HFaouFK7igcWK39+l/8po430JCStzS9GJXnaOuaVtOVF53JKGS/y9Q3iP6yopLzF4OOwxD
T1goCYcFI7+gKMfb2nQhXXNLDwyhRdCZzlyPCSOtkjJs7gcQK+ihWm0QVzACwOnQF1fBK7DAddU+
LDwqDfaz4w/Qkrc/emTGtOvNsmEeyQ06DT8gcpymQ4iye4o2u/Upj2pHKxb5UI809Qm34gKXUkPM
625yospu1U17sYuDyXXOjbJadjfPNsxk4ZssWCTzhLQDuboRYC/Daf/Ut+vP4YHmkqHgrxpgspd/
U9To2CB7Oq2+FtRFGFaJT9RSRgWau7qiIPBbh95in55VB5X5g5tX2H45wNqpr9M/CxdPmo5kH+XE
MP2Ft9SxYiiy+/KJorrqAEabsOaWC8V+sVw9BblV6Ypa/KOQfs4LrM6JPNhp+0KN1C8sydH+VOlD
jWa0GIb1GmFVyj9sUok1R7U66+6AzeZA393tHhCNPBxqdgjQJpj/CXaleW32Px3Y93HSEinLUz3j
Q+6j0+GNZBEr0YnSa5XI6QZcUWzGbW+lM7Mjx0x6SG4I84XAG7XplWTHw56ufkrD0Uf2jH5O8/Z9
YxLa9TkT1ymtLNDL23X7LYHnYQMVP/0JGh7Ml2xNtf+eLLZz8z6z9ruipwN6i5IHqfw/h7s68eHZ
KNiKaKNl2Bo7SdQbzCNBhOE56cC6i0LdvS4EtO8vxH896MwKzubZs2V9UXlRZZxmuaiHF/YI/91m
/LMDbZA08KNslsw9rtVeEqBvIcniBmvootzFfq8yKtnZqb9x9b9cS7Yt2Gr/fT0YpH47YzW8g3pT
Oz9Iv0buECG65Ct1tWW4Lfz9uWJcGB71FYkOfeGQb8RYpqP0S795a8Y1RGWYNwOtZ4fyas1CGGqH
yU+62rOoZ5ZIUsGtUHy/dgLXeEYSQV9FdgBUqohSDjyaFIR/9w4ymdGATU85zvBbwc+ndWdOHC8i
YhyJW+jBJdf2dYXUU9LLIHpWiUhw4+kzhOKShcAgkSEmpbvMm1hMd6IbX3infMxm1CUqdP/Gh56G
bhOI/7UWdp5Dn1Wul5Ce/cc4bbFITD2C7mujhBn26hnNapHNIuSUvJL8lGVRTQgY8qG2aqoBNNAr
WwkJe4INjFbhVoQvd/Z9/j4wiFcP+2zW3j3PEPcHP0GjubTimNuyPB8OP0hKwZ+wi8pDMfvPp17T
z98UPOQnG5MI0vVpS8hhtgho4j3lOn3YDprrvV4S0hS3teA4IEsmaP6wci6ifrhY1MJ3bDSlPXjV
ufhBm29b+4ZAve8hRgilsGe+aooZmW35PyBchz9gMDdd1XElTUDQ3bnL1kIk7/a2I7P54XD8ujQ7
k4hi2bp00ZDNvX0NgPHCt4DwUm6yLn0iDKq98YrPChUL2oke3PPRH6mV3eHQPfHXnZ2sMCnkjEFd
1+vz4MXFBi35o/HmZssWG9Avwut/vqSPpnycBfEadmp5kP9lXqNh1prWJBjCrdn00JxeTrvkGjC2
acusv0K5iO0feFxLNFOXPcm25bo/Pod7787imXc+zXldXIx5ODNRT7T8q58WEc456EaTJsLIrCem
W98wNGsFj6fXrQFHFEDgoSf+UjokvRiH2FEV5saQfVYO4izV4JgqYOwtwd5tVXOd18iq/QlkaioF
Cs+7GGAYtybdL4Nodf1ESTDiSxk5XaH1xY82c/QTtr8Igpf/qqqvDXEB3XSuur8NCKHKN3YA8Mno
0TOGf59aSlLT1BjQpy65jVLYoaEjd0owouv6odgVYq98F561hUf9LSxmBTnzK/CeciVhNQE2ndk1
QA7ul6uEiGYbUQWWJRvRqt3fsuE0muyD/+G9UltKFI60/L5jLIIwZ84/xOuhgoyy/aVDGEEXwuQ8
WthIqBJ6IUVPBCweCjsb/CFb1y7tr8mPjRecblDZzFLq5C5ua16BrlDG1uDGHRnMDpm/DeOkZP8U
Y0r3K29shsSdej/MPQsK/qUZkwzC381vTg+yIsFxzje+pb35SYHOzWvLSSXPeaFxo/Pd+W4ZipQo
UWWyjR5o8NmES0Hmtboe19S7uJnvf5sjQyrWt7b0FUgGSi7dST4RICar7rm/Pj6sYOOYcJX+RYL4
dCfK6Cof/QuCJ+qB7BmTuDNB29v/u4S7ESmSwScwuCDpO5IwcnzNZy9EyXhLFW8NsZ24auBSzLwX
ocaNtvLNkyyJbuoq/YwOGhImtH9qyi5sF7qkG9gmIIz4qbHi9h75vkj1jSMo6G+RM5nNzUHNSWjT
84iQhNFHXM1OPlEk13a9gFkk9UmohTgFQdPw4ey9hAvdrg1l23qhMKQmnkQ90ZSoOTZwD3/qCFVc
aiOQoKfFSt+Oop1RBsQ2Q1RPq/dJuGHuYNedAF6qOzklVIQP1jvP/TmHvXRlRpXpg2IuCSOX3I8D
dnOl+GWgyuEwKL8V9xoVHWKDz/6IOqfnlsHrCwkHGZ/oNwJjTHFZDcf7k0V3uHrUmv3+BMOGUi4E
OkqsZyDRbZCSjcASuS8+y8VtjSiSF7pmvbRZrHPV/psBqk0z9cRLXvNMxfxkq8FthxkCl3f6X4bM
N+SgQUx0nFzWIQQOU6cY13h1EiLm0S0zsrGKubYRFtJna2Anh9sgaleuCyfo/8D1P1LIx/mAHTWy
ZYc7wT2MN5I0CMvbPZPlrYPEtAm/fY3RQ0YpD6BtNy0sh54Gr3va4WQHp92qEtb0b269AzBIEALT
QqQ2AQY90ZZHJJmj94+CYkaEm8gLx+UK4v1fqZrulrRAO5t5bcAKvs/rxZesGgSSEJIS+CL1Auhc
syS4uqcFOON3dhBNP2I9osXb4zk+RCHvL/0M73qE1fsNyQxV2CRjC2/mcNyeujFzMk7c6DML3cxo
FRA1zU0Pgg/BV++YqrxNBLYKGjK33g75FvavtObgH4IPFHnLGg8HHMpEKZ4gpgXeKwkhQJGtSw4l
d9aN0JzGfKxElTM60V+PNgbqraF9yFmEUXibzC4zZaALN8YU/UvJTp8xkBk00FqQX10QIcFEffaU
IqKDwfFkYiF2AO5JbLcwzp6pyP57pb6C4RfpW9NepVftYLjVPe3kiGHlnQk0nvQjMBkS516WByfv
gHZDUuchwhN9gHC/Vfr2BoCSGyNcLjXGj9gWcFqgX/WS41v4Z6Ph1osi7q/MwgBuDxDTSX4SN4Ju
TNprlVrLZaO8Ci686DkWMXgeRNnGkPuaaT9osR1nLYdXZMGXCG0jbNB6qK+PC9CNNG4TyaAqqiLa
SAX4ZGnmkaWpZjTeHNUL3HCTDbcOHGWSk/S1H8q+Wb/AGDlhDD26NgLeAXX6UjKyRf0T01GrtGxL
ombFN2mRWDtLpfqGzglU/cD8T77ilkc2XOQ3IhauCDT4CogOZBzPXbt0wBRnxXbYNU1YDAr/C4ZC
CWqdcuGgw+aa6XPRdzVU7rrdua3Vv4X3OvFORyoq4IpR0eXdiDE/hyYFNYhh+r3Zx9xAc3wBsELN
8AWT9jFaRf1qShgFrLq2gMZ4EeFq/IUfkzvWKZNZUTzQIwpW5DIp4h+oIAmC1NAMshUG1GxXsEqZ
bO+/YV1thi9xa4ucJr2MzkeivCP9Z3LdBGpiM1nvmcthJcgFDd9xo0jwXPUYlc6Nwb4YQ8GIf2Rz
Kdj4FYRVAtXC3mvGnRgouMjgxYVaslllTBmEtoVwo2DtMmpbG3P124PEEBB2Kluz+EBeyXtxgo8d
wt9MQsiocEHwjJ/RpnZtnFEVfwjMwsElOfHdbvZ0Z0511D9smSB2SVBK0PHzTtgXtbE5Bdkr3/XX
p5maBuR1C5oUEQayFSzFN1pTeIAfSAaPSfAmZDXoCk9udfGafijFs2hP1DByZ1VIcbDUDWEjOvfi
n+7Fyf2+v20pQbG7pr22U/5OrLKD8nWSa5jGEG2ts6Rq0W+VoYOHaKxOl0yM5nQdLoQEY1W/koDi
CKep8H/wcgDNvxRHXvg1lzvbytf8xjJKb6CyITfbn6ovb5xkNSNUN/pvO6z7380ZcaVGpfL/Y+Rr
dth1yAoxQ2L5ORiRThw8Ue2HqyvSSTKtfGWzBR3jxbj1e5OimGLuA7NwbFqNocHKLNr4Nhx1qhyQ
w9PWcnbXT4hTw2AfLAsVzDUbMtk2GQwZ7/RIkIW45AdnP4qWLuSJmu12M2WXE9MSnf+v+/8GNAA+
BkD8Ool7jH9DmcSid03XmUSNKSohlhztEZ6ki03Z5dZyr1RjJPulYi3CJVsZFj20IbeumTEdoPX4
kpXqBQqrlj02uQejh7klxJWgO9lYIJGdp1thJKy7/dKGVtJH1dQLk+/HII2/mBW7KSLA8J77imMY
Iyk3D+khB2WFbnKVkLbY4D6a3nH8KtQ13vPsvSD/ohEtZhBNGSC6HW0us9yiGUABnVoGEqUdm8NF
F4F6r4LQBudlAXYtQ+8dd1gsl3WX189OBRKMD5aAY9T86VWRShcnSLGyKwUJDSOlusVj+PxULrYR
dkg6cJK8ZKJmUffLPVnFXAzkZ8ZNVdrkPENRj4uIY3BEwpVqhm+QpY1ogF7Ky4FWtxn3wTxAxOnN
4xwB051PuuMBieS0LV8UiApuhtH1BOObvRvP/YxMmoR8y+I5CiV9DaNpmNgTEMsh/UF1JC0l4tTJ
Nf7kU3KIDxbprES9pn3l6TqZiXzeenz2MMEwenBpyYgicVrs4rb++w8O3sQ4wwKwvEfLU68kFtBC
/19PUBw7gTMrbHnMGmwZ2JHJYGhky2Le9k93efomHlchDiOhr1Pl+PqkTndg4PLd5jrBvOHj1Qv6
BrBVmNYgWufgDAQaRjGI7tKk3IoWxo/cCGZle6lIQYlh/sJBqAesCRiEdfN/QDMUJMpBxdF5Z8tJ
R1Zswrvk/iQdv5+mwcHUEsg4EvnutuH/CJDwrlxY63t/5RVzLiKwiENR5s8lj/ucHIm1vXqavZfU
7SF0BPwFUy3nYdWCkbYMIE7E2rn/E54HoQySLidY4wnAgyKxKC4vavvnuNxV7ci76ktskpKvwYUD
PPEjI5v/npgwemZvXBduLK/ny8ve5TSEA4UUB6U9iJiwnSYIabuZgWgLXUzJUKh0lOOdexZ/D/c9
MaUotOG2+vmCS3YKIiqr46wWpnQPzGIlwuWmbKekyAyK1H9MaiDwpq1cC5Ge29HR2NWACzNTNmaS
4TdDBSHBvVXCOoAZ8SE9dwfruG1XTgxChZDZa3kMYGTpkqLkxjDVCzyFgjHFe8pr1Es+qIQs2pzx
DVWRTkh+QBfV58TituhuhmB/vkdrYcDAiYbHwe4Hyq1O5LBVSB7E7B9b0v8xU5GraOmNhNdyHf62
9SEpzZKSMJE3jv9eUmsIm1q1CxcRzQrawj+oIOXQrkSIlOf0rSXzABN6k9PbQq+Qf0+iHy9CFBr+
Z0cbKFKm4Va8ZXVO2KcdQUSE5gQr5byBxErZBQtWjzG8gI4wCRSM3GMe4z0kwTTEJUqN9fJKA6ek
B6o4k+1G0iI2lbq/xLicF58aub2RtmmCkwdqN1E6iPgsCX/OQIIpgrvNg3TdCzqzti5nYY7gx6IS
wueD2LHxSkqWbS2WeJTM65IrruT0oJ67EYFR350L/aBFUrmFkCRtfZcj9MqkAlrC9iUxvOHOTorQ
ywyVV+yNzPj4sbdH5n2hnTshFqEX9sGMr1n0sKVjL1XdFUdSH89bEADFFJH3BFBmZ9+4VEA3Ze2/
qOdBX/igvOnZ/LQiOfSuBU6oiSHJaak+/5anlALrU0oIe+0Z+wV0esofjx8G/L+p+GQptO7lkEMQ
jPWPwdXCuy2JYoOIxwobSxXV+kaPh9pjEhHkoBPWYJrSy5RsC7KZFq6omlSMMJIsaimaKXxVSoX6
q1zXKRG8Gi/OI95n1k/4/3RWFmv9ndy8IxZwzxNbc/ograhVqnWeJSBUlDioU2Fh1q3nhUsMVpPP
uYoTHG5LRsgG4wJXnD+1g0wEg+Kc/5p0bRCwy1IQJPJuuqBuAc6T9VKfONrlZN3FJQub0LgKspIm
NN6I+gf2mp7bVypiccRlVWNDMmKvmmJfHX4KUCOG1FWEY55pw7SkXXiWIK9dzRwTMT9Gthg68UfV
ikkLRwVG1J8Yvj1xJUjU9R0c/zatfVPs3R0PwgPCep/PZtG7jnrjc40z3Y7pkgVhXlscarOU60ZT
it1EM1ZP1UskQb1eF4AHJRd+LzrImJfaJpKP7/ZMPScZlI9lP+iMPSI4rC7/8uqzRuz0fZjYnduY
YFWgtQLYt5jYrWFCRzjfZ/OVzRf/XJpiYVUYIsoZmDeXbqOCp8GstIblgO9vD9a4tq5Q4LUUWTyg
nmYUxblxd156ghPwXK/kE4HSSok/3UZrLyJTl35z5y/K0dulWH7rVtodgfCKtLKfTfVwhM2Mogx+
LTjAMHR42z+QCw2kw3s5BmkKS4/fqk7X+KPX7L4pMv1ddgmjuKD28XLCshjEZQhscXCyO99X8I0s
zy2w1GCr3Pnh7oYLwPnEycjPOzG1v2XKK6cL0fAGulJzrw0ptH/oFqYDVtHwNZM/JqlsgHVGtOef
2Me1wOz9qUVxxYUUm+QPTeNAP+blN0dVtmKLtPeYQO9VAxXF5iOaq4XouwCU2wRLbQAOLhtk02hL
8k5yBgnGHkr+JZBvsWJq+Ow5Rw4+ottqZMgdubUdhI5jhJnaOVvzZ7eEIG9jyizi/paw8IZrfU7t
J0t53zqdf/Vu08wdQtCoRzuK3zgmYQBsjdBzdVu4dQG72QMlOiYQfdwCnYM7wFxw9QdYaUAWM8Ox
lULqfA5vTJLww0OnTTApQRmbH21+i+3d7UCQioJEL86876HdiXEJ/R9h4WHs3OzFCG1laJNAuiL7
qvgM9+AVS5W2Do4Kx7uJUXABzUnr+HhSfAFccU6YOqSh9cD3Oc2Wy92wtlgs61O2oyBaGRl64Nc3
o3Hq3gQsoFdCTacTEtv2aKYNCti6NYmDv6xgKvZ6CQFAwCI3fkG/7sRCkgLmj1ouRLLNDnn7BlE/
hejlRaYps5Vu0vT9j2rDcOC9RbwB9m/WPvuR9XsR6A8c7web29wI/KlE007CTH6ZNch4s4rZD8m1
74QhrESkuCn8zViNIFe8VciTTqrqwBNoU0BdVtCaZ52F9YNmLFyxwEQ7wP14KBA/JUq83pB8moWn
EvTBIr+kJdDa6HHk1xqYNBglmbmQZBRdbckyotkIWAlBmCebg9ed0Jhpltimd3nszwelzRroyOYa
mFheLMU7qtDmKIEZRWVj+2cWPZ791khKsRuRJr58WesSFWKvqofbNVmjwM5Mw5MwNqIPLDxYZKpG
qehFcPsfExTX0hnzyOXxZkJWT87DcSpYenQPiOa5vJNTWp+SPzKlXBcDk6oV0xq3hpngdl2i+fDb
08qAwodbUvgKZEuKP2Qcbp4lEexzhzNNgQiRiDmb532sbNAHaGqCTqYG/KWNUIWy8VdL/EQ0Fk8p
7WC9ytmh43cy84L0sbF5wCu1yIAMWtGHl7K2/qpCmCgzlztoTy8pLzMCGfigOafqsK0WCEWCP9BE
yIie9lZN1eM27fXeA4wQ+oO1andRo5mOK6tv7Fz+0djUhsomGBxNvFJjOGYwy7xCZd2PEjNF816E
Wj7Fw+PmHcJ35Vl9weXKpD1JATkJHtIM1K4kd/YaxSFNKSZImLGMQ25mcaAu1wcHrdKvS+MjAlrZ
mA1j+B/lmEtlTOGeUTSDQL5oVPOpRJYCiz/tqPdIsUddFvUAOrRzgU7sdhkxf2rDS/6Dc9Kq5y1e
i1XWx1ElYAjAs69t39saKqsWh+oofGz3OIC4nVfE0gMX+9x84wDiSDWsgegAAlolnLcCWYW6PtaS
GYqdqu7QEj36kLvbKprdBmmzz6ZUngZ+9pll6SF252z48xToqczaN6zgw/KFic8hyTtNsY8d/jny
dzqQXrBSAMk6rBoEaACX4YV1RE8L36/MSUxh0Efh3fCjp0F0e0Bf5/SfZM/fjxWWmIt6YGJF1SpL
72dQmI1aZio89yrhXGe6/VdfrmFPuxBKCJmeDh4gvbfB9ZhdFWdPVWurgEKmsQWFwCGOXk0qYjgq
9nj/KHc9UzpcmmMlHzMcOPvKBoCSsEc7LVMNe+aDp0gpwyUu/DMa5J0kbGmsPylbw4HlGUNubkdd
NamMEKYLsoh5t/kVCYe9a0RiJSaIaXG4Xg9zbzUS5WyqMXNJoV4Y8wBpH9bLHBrHnYcFyxbRrx71
916fjd6faOhcYP76ZDFeBBEDjGzUnnbhgFkjU8uE/MekJgxg0Tz3jzKrnPSUNqldjYNSUhrlEMgY
mm7b5ImIXeVZRVf5uvrWMLnWOjgN3NZjb9oNAQPR0xSTxyZgQvv71z4TB83ITjcX3V243Y24ufEH
rPeQi6xtOKsoJQ+Kznmw7/w+0LhOsRD0I1hfCF0OLG0hB7oL0qxVqW7FYRizNjRYpe4DRyDR+9d2
IE/Wvh/2a9LfGKQ1Ork+3UOfbNsq1zI5qSLZyl6cLeRPpA/N9VaGaTpQkxq45QN0vq6kbqdA9H0G
9CxfyjYFDw+cyKl1irqwU9bSqYtOyH/ShNuO85CPbDpxF71IWwU/oysF1uLpVkfFFMdxFE9a8yd1
uyzd/OYfUT35wSYLzm529UokI+b1HEm+CKP/Ocyz3J+o2FcB6rZAYI3HSkwcgG6w1WyACophQEuZ
bRfJrKAil/5pa9OPOfXm4ifHqHbQGAhZh8ym3bf1dJtdt6UmDcGBfBdGbjTlPRc+bUkwGD7Z4M1I
PjsLHeA0GX2c9856QgaJUCbVs8rK2FzrWbXuHt/CyvAJb7q2vLkX29FnORBGLxyhI83Ij167eC7w
ff4Cn4Rcoamvl8LZ0MFSkjm3kfPkKTbT35fivQT+1QB7HyBt0wFwBuFRI3QX8SS03R1oMHQbKXAz
MfhNkJBphcMWqlPkFh7vpLNe1bl7BPyY4+WzTIBdmGiZ7e/gjDL9oVozS0m3ZdRjc+lytpkVVgX5
XNDWYaeAq7bF458kkdUwoKIaDQRgM8ZypSZDzoFmE1mEH+/WRICS6XbSqUbf/xwfcLWSdQJ2AafE
zr9HHcgUzWbieKWfESVHF6K811mlSJ4pZOmUFAGhvoPVir/mDoqFrPGSwiQTPTyYKcxmHeekM19Z
jDhmVsqwcAHPV0XKIuPCs0VpeJdRehlWizrGA+46Io/hwm4G5guzqfF41A9zgDxZjgj/SE+Jg0+5
awzx8MZIs/IVO1ZoguPFFaPsi2eC/ceVjaspwddARiA8B6daAeL5/kXX3fMH8bScSTCuB2Yi49U3
LMQ5wsNGVcF7J8geNSWZhvjtySzOcP0L0bVRpGL4ctJwwUo/xqwhjRpAzw7OAGdB4fRsDo8i/0ql
q2etd8zM875CF1DkfxHHP5IMV0Vo5llL9sxt4LNbDsjE002+0nWpSw1DKHB6Hm5cNeKShiLP60pA
MVw/q91UHgyLcyOt9ibtOaafXaqCfJuljZ5HaTVO02l9hI2uDzmn3q6FVoz6Cnd+HID9bVW4LHKb
0/7za5jdrSrs/L+e5GyiAboJP32xHkv7VDSRFhBgbmL4LktaGDu11c+v33dv26Ou1HdFsJCgD0pP
6jY2rRfOCF1SISIZvIBruNolpgTq6h/spmNZd50gDEOqXwKOx6+O1EFyyl/ohBn5cWExGj8g1zj3
AdcCltTVdY98Qm2E+9OXpJgvK7Fzndgwb259nmkGAarYDdgglEiP+/YuGxFcalN9yCBuCrSiDwEP
ZS6aaIi0F+4TPtoB4gqInN/626hZDLV3LvQRIwd1y6kV2EEW5xXyTYTIzfotz4ZQYEV6whN56hsP
4O+ESpnJ26SZSxEWxCbIEThX0Dqlxwt6xtJpcYJdlK9zcloxdKuaPJOQAiY9CxkIYFvM7d8i46yW
IqMdFLVTY43bntB4vWDaFwMuSUAkcSa3fYxLv476Dz+xafhKNqL/P2ZWagu12QwK3dxIproW03Dy
u9O7Gw+nHIoTn5fzHy+RY6zy2vTzij6yOVJ9kt1XOF0pNOv7/fDbHQp3EBEu3YKUCX5I6+O53Kqe
iHLi/9wozHznkf8PlOOsrE1POXJ7apjaghQdTyivRur43KijUWc5zZwuuggMGt10iPFhppUPYxd/
Bfj3G68A+FZQaxF50CzS7+WEsFeAmZsD8MbHlS6TKlzcsGly+BhkVyOagJiGj48ZHjLAfTc1Et87
jjO+LSnfOShvETIUqjrOY/heffMNHaukU4XxOQG5sCxc1c4SAy1JeYPWg0eV1vGjd5JOgymlhaeb
ZoWPXYYJcaXpRPxc7odPNdqM698LBVKZZFiWyfc/jl7+EdmNw9QmxT3tQl/bdwj9WU066i/ba6cr
0OdhcsNNGh9qDk/vOhDi5qfGJ/ibVyFGwQ5gti8sPK5BE+uY8L6oHPobYI4nAm2A5wYvNIrmV3Az
SfIQQSzgPtYAQL9xQ4HNZkZYvCNuFVsoOUp33yecHCNypa0IQGKZmHMfW3bhRKNyygY/hpb1n2py
OAqakFpWoisjOrg/nWUVm4+XC7f7we8Pv7zVy5CGw1FPwTV6VLWN6DelMlygGOSU5SUqaljk+0U5
weKcVPXkfDbXdrrX96Vrj9HWBbysEcyHIK5Cz7IREENe8JjniEu6yaVVm/Ex5cAfLeMQ/6JnzFbw
vSI8V6pHQxyTvewAUj4ErHhI2Rwv9MXFc01EbJFSKbroB91XEcizd9HaI1ootWeH3Qo9CPIhpKiZ
oETyTZscv4Ix3pNXxYJDWIVlzEdLdIsByoIpstVesENGoxut9d9ABcAdHhaG7L//ajk7mvqe87QD
5GF8J0JnayA6znFHE/sQwgYc7oQ57sDg0hPiJFMFKQb99x9dKpYMePCcSlqCz0N/6eccYyNZF/pX
fkFnD95yiivoPSibgTPvL1svTqmwU+nhrasgco8RXnNJqzleB7Dz352Wg0uh5agsw+LjH9Dw1IwS
uTHzfUt0aopwpBTeMzTHoA4gmgVjtXg9GorHCATR6sgOw+TBGn39fz4zcGLW8d1QjHiv1wYNWvit
Unqs5KtLjfJI0D5Boj4EqVX2c1Z7kuiJhpME5GrhcRZLBEzisB/d/6grV3mTIRPiTrjNj46rQ5Ea
gxDVTmcDe5ffOZKsYmvC/Hi7TvB4H0ixaQ+3j2p6q74XW8t7EEx9pCQYV6NUHh/VkMXOVVdZab+g
nf7x85eqleSoPIxw9hxNDCiFfBO6SMex391H/crqprabtVTN7r9pvvMAjNJNMQTLq5CLyAKV/aTH
a+1S35y/F/rYuiyG/dd+UVTvvv6mtEBbcu9ZUoUX3jIEeciWt8pD1Jjj69p1Xkg5Huky+D2kjQhS
PniTdwQj1CcjL9cKUlRX0339gS+SN47jNaPUxJX8XFObCfFh9MP8XfDfWLuY75s5ADKsQbXBW1vG
hWQQZp3TppbOiIbvun4p9SvnO5jVT3f54n7ZQLYJhC2tWMgRBb+HvpzGzSj0hnAkVO5TagBqmIKw
gQbZCmcLdcJRoeVSVyUHHFmXzx6Y8b2gH1z64o9u2IM7CwW0hHtf0A+PTQfoao/3kirXc5SMLjQb
r2pKMyCxuG7851C+71HcyYXLVsv1j5fmZolsU8hQa1s5vXDd5NK5lBsQAIhU0YxELaZPzVVuonpZ
5fXUpyya8bd5dxZqyd9p+JNedEgeY0mu+ftCHa4LhG9pY6Mfa6rOURvSvUVimpdlZgRibKaOJAnh
kwCilW2tStVUQ2arw3V3FNwqRzUmyI3e9JgEF2mg4wtuMJREOsk8gUNhE/pviM1xfAcnYFE/ffi2
rjhuItwJhNu5omjSZNurFSzh+QYVadi1dVr5BqncAuYWFpPJH0yDcDessNXlufmpAFfa/erVuhqj
rMru02fZsAYMpnZIuFFGwEITKUKgxr84D2tw66IMM/V0oY467g63b6dhGPrzm3btziOdDUxQYNcW
lzXdgePF4gzxVkVjFFmEsyuaV2scrD/j6o7mlHlAb8gA/bClvRy3zW9wiww8zKAagJwBVjmWEhpg
7/g47yVJ7M8j4mzkge/N1OyQzLaoG3doEzBy6EXJCEbIp/bABhc8YeKpzH0HQcuUE9HMx9gLG0fO
DJ2axNJWNb6mmeKrd/LAl23fIVvtxMrDveWHP+A6sDgbp+0J8cWqKACzuTzaIyojxP51pNrau169
a5QhCG0Z5zjGpkzFbKnrs46SisOMzEpqooANH1Bg45rihMV1eoFTbmmykZkzc17tRC2ldoryKIzZ
cpTOQ+tdcBo+hk4H4U7iW+RuZQc8N0jkfnTj9dGie4rHgQRv+D1TnGR0YWYCzMasVrZWVQci78Ea
YJ4uYoF2+IdF8aGktA0GAIQM/fS+QdXXUikazWCt8jM/olwNHxDBuM/MzEtbL4Zz7p7QN8F+8Uyx
l+QiglHm5unCkhljpMyzuC8kpCzfHZLaVcVGH+eBG+JKANyIJY2L1cyAjXbNe0n1CQPCWVxalBhB
w/X0YCaQTgFRu9yHdh+xZfLqSoEujrasFC3ar1ktRO081B2y397ScYUEUeY8dEvw7cDymKPe5SZv
JcDIxHEh65Y9DLg1BvmogfXoesNyKJNkgG9pbW+W8+32qajOwOtGztUBWNk/+aVe50GPFIEa5riE
Z+w2pxnGgnGatBPfo+xxlkl8LuGFquDDPCoA6NHuyNceQ/BnbQJujo60MllP4yf5YUZ3jyXaHziM
QJ+Yqau9Hulx2hyxF1sMVPrpVbhNf/HdFzvtGqFDMsFVjxYSDlsFBAYH6VIAxVWF8w3luGHD43gD
/JU8+PXWXX+kkqRZ80sTxwlgpU902SQgXjcUSxr6yoNIJx78HatPEahtcLw5HA6TZ2K6OhSQK80K
Hl7gkyVS+UTPLNIEEcjO51B3diB3R0k2IYD/mWnJP4suvDAmTYhZXcPP+6UIDYmb/07BrYpYI+94
ItE3uHF+5EJApVzLTLOzxQ7vIEDsOfCOSi+l4uDyQ/u3jQuABTEfA6Eh0R8gsd7ih27e0O2r5t8q
e74oIgLMXihszhR1pRBugfZDXpZtgrR3V2JQYGTXFhIAfsYCYfOt+/f1dPv3+sT+xzsEtYRdRvgg
dxP5p0APFkXA3nVcDCyQvqbkXZeFOfT/CtP8t4r5IsfBkv+Ir7DnW2O+ctzhP9JITeuypktatKre
WwPkolJz7i/Cw+Fax+qQled6wfolyTdJ6fTCBBKnWoA+pzk+1pbU8rQmqjOhuc/7VgksKV49srvb
vt+TAxJTLK7n/bY7xChBPZH5kJbdvzepASlMyhl5SUvxluNmWcZozcb767Kk8/V1V+wFZDWfw/mW
q1ex4hggkJgGix2Vrvzi8D6/BOpwBcd0Y4ALAaorNJLkLomLpKlRaIGwNWn2SulrfoTStnhwHia9
uElnyBGzETwh9zo8F1va12CrU42n+T7LR+URpMV1CqckEvT9HvtFvCzyTJ7RfmgEcL/sxkql2kwJ
MB4FDRB6Mz3vFlBXKJ+SGkwEUgEC8Hfh83uLBsv0gEgFO6EyH2YxCK8rC3paY3eW8gbw1kW9fLDO
X2sBb9RB87wZoYe8NqNVWRLyYR1lS2SiU4WYdVD5I+5VQ8i5TR1e+koSpx/3WB+iZkrLtC316ZPU
EbUGaBndf0CGezLPDx55zv1TIXbeD6PhoTyuUw39QdnYGkd3iu/quknA2N7ZSyHrGEE7HnsWMGPl
toqVA2+eZrF9/L41hlDX8a7H6jKvNFPNcJB7Fs8x3TBDB9RVcf91gh4cDPuWuxRXWol8cgd+MEKH
3+jM5XMragA7YZApV+LxJSm0B53hz5GfcsWFljGnA7lGS/317vd+z2l8XXPjQFu+ka3p+9ua+Jkm
h/oghuqSawQWdzte9+uVHXrWv2GONufZj1hjh72BTUMQAnxttEPyiGube6EV8czA09/vmF8Q5N42
UASmkwxc1dUf6n2yvmU5U2lU/tvE5V14ESuwZKzZ2J9vWvr+7xmkbl7x4Q2HexdlPcXk2k8TQ4qi
ns0BaIwCYo86ub7vhfIyJS1YQOA6sSQWRs0G4VSnLENrKA6nB58+K13g7BGpZ7xEkzoadRH3gLTh
NeQmXRr/eBiTIQPneFF6Z9bAW2AmthYSIFUdQT4VL4U7cDUf8BYqeIWkBs9R2XyviHMgGzY7EHEf
PW/1nyTNJ6xiFdEO/95PI0HHKdQqFHFwTg1kowQHZxiDZGZTqyElYjJ8oC/sB39xQTfUNt7YQMEn
Hai/GpT3WeSYjEShhWebJhb1+YxEWn0nIqwOpr6+qZQMin4E172C0VXdyWo7oPwQxMprU3+lC8OX
53FaI/B0IWh4DxvtTKSSd37NKM3oY1I9T7e8N90dQCLjKwKxu7pv/kpwZp3yFaR3K5PLAv2s3usR
D9+P2IiOxmEDHWj2hPTLTfKQhluwYhuQHxLvjX8uUiTeOeOqllNywKQJL4E8DhOI9XmJ8uUKz7ek
Qaw1O955ZyHK6LnHK1MK0XniBUDgEBHuF42uDpW4Kl34NnGn561cDDxh3OjCoyI/x4DyJWGVx744
mYezxH52vgT4YZmlo61agwTEJsrPDkfxhNr80eG00Ii5+fN6uWk4zRu3Y+0B1gIaT2ZBSW0XfQmR
EuTpgnYX8A8PC+6M09AspBBX7dOjS8AMiPZoXTEkPUhj/9OXR+3Q7b6f5l+dAsgvyussNqFPytka
yyP/Y64ie+ntQSt2nsg3nznbqEqvm+2ssxOWNCmdxF4Xsg30DkrAQ3BDlf297gl1XLB9DuEu+1k/
PFOdrs5YlJI2mbVJHVRJXjXHsgonAt4bgSjfYkO5iGK5UbT8X9HYrn/kavpB5du2uCgTvo1EADnC
fRAP2Rm3D6InxDMBeAl27DWP8oKBBG6F1kp7m/dYbVwwl4Pi6bOW+PyP1XwzQPmwUs6IN/qseA7x
Cg7eaXGWrRN+kfIJWlSDj7sH0eSpj9CU1rTNaCtiRb37bS2IZHxp3MQt9YXymJUrq4+GxnmIFL6L
yJT+FG6G4hIOCFyFYlrSELdEXBk5YeSwoF+Cec/hjSTbXEUkZSv9ewQtUb0QzTEshX6kt4esMbJE
PKFm31Ihm7bfG7AnWBeh4Dl3Kp2UIOzFBfDgkzvln++3z8Gb9JqRogtL+qrLzO97osCnP3aCv2cB
eYrLbJc+U9FH1L+T1Cv2YW8bWlLG/wtKuRj1kfRDlrWhTwp0KkLYfa0hHdQA1SD2sS5DfE/l3ZDg
OwjTv18aAXE5F7r9uTiTTUcRu9X1csPXT3PWNyjI7Kls64SvAX6gwfhSN7T31eo0nysvSYSL+bs2
I7GEslhN5sgFzAexxwSBKSyyQLOOTasuITt70U4iWEAzNKuTaD9Oc+wCOmb5TM2lHxbp2/IKJn+v
ApGfAYi4jfVDdEA4Ei33stgIWYoF6dNOA5w/+gzzxBhaRSEQh6O1E99ozNMmaeeeodr5d+qhZko1
CkF7UmMIuS/LyFayd/gyY1E0hteIWLcBeO+AqmXcHQjrSrj1JphV3U3LBhTeMdqiAPrnGfpouNzn
WOSuJ3vfepTPM+sx6MJrtulxL4dvgLjbqzd3lID6UDG/2ucNo/WQ+/Del+FGdV/lCd+Mxm9ZXdEQ
ipUVSYhnozfNr++Lij92yZ2L4Xo19DjeLMQqiYsDaaptdfTea4sM2OBjf8WPoa1tD8ofsv78B8yh
Ndco7CfX7EIjRSPajgOaYHH3fXtwv82bXWhPHIjjifD0FO39N/WyoHahppHPkNeozKuCKG7j1cK3
z9oaBSTDMcJcLXxf+G0hwEoqqhBS0B9mZrvDGJKaVdHkc6RxFUKakJUrvBBz4GzLsPd2grJxko+m
lNy8be0Goblyfc29eW8hDR9+GpYa0DmfDjNOza5bxSgMoUSSlJV47aDtAr2QKElImtehCkOgFy5e
Xkd2VYAHvYxuk/23wfIrXL3v6Ov+GYwr4f29n1HhaL66/Zep5UrLGjUlH+gLkiVtV+t1JrV9P8No
9To6rPtsqFyeZrrrkfNljP8uHfXgOHZE8yiJn9YiJjF4PZzzxFw6lsfWs+2uIi3yUOGeGs5Qn3lF
iGEJzMRO5afcmYxhJUN7b0md1S+lhaumBt+COzl1dva27drAIgHTK0wCmEKrkhBdDt+hxIP77aKu
T+2f3YqZ1Cr1+8Hn5l4bVhC9gP6g76RnZGh1KLm311ZhxUfqp3oEGggWHqnxE3h0bHqJypYRvT+n
MwQWE6Z1/GlmyBb42Wp69LBqSHb4TrqS+BpUNhRtbbiC/sL+g55psU1xet53WYx2+C1mCaANuRMW
Xe1qYI2Cp2uvHEn+PVvrkafghbEt/h5V4fa+Rl+RsqM4nlItpNEbhDGwILBld7bSI8Gu385fXNpU
32303w/wWA6WwZlJWnAlDAyCtxdaX/AiPNRWLXJiDOuoZ3W8vOmZ5YBOV2iZcDncKi7c0L7G8WvO
zTLNQE4Fymr12LqnHQkdRtVF11tNJKbTI3J5hmUoFNscJOIT2wzTfkGyTgOxCTmhWrsQMEfJCVvA
LMe/bMVnAR4I5O4HvlVWUkKkRWir8i13Csq/kGqT8gtau6yvA7GxzDyjYIOV6D62ZHEW3xYC8Vyk
dPJUkcvTG+l5FSRK+EpcjSg9dccLC8DvL1rSnvayPG1Z1jHeLXcYtLa/ZLeFQiLu8uZpOYTq9f/s
i+oL3Po1wfeJ/3oYWpUTTVAmIzwZKJg27rPPQRoW5UQjrGBsBbior8y9zGI1vM270s9D8/m4dqM6
y3lAlob4VLaFWZZS94Ux6isNNBBm7qCrBCPrNYOCfp3tLAWTE327tIdvPm8uK8nL0AXfOJADGETj
EwbxrHYFiQgN20Xqo9TvgWHcOhTHgAVTvLgwrS4NDJ6OLR8Jghhq6ONC1mA3U+wvWyfcOKJsXyBq
NLIZDxFKxHz1PN8fzKJEBfy91XJvvd2jWsHecWcl5+F0piZTcMRC7852p5l2cr9OQNWPoIno+u3u
MqvKmM7Ulss3SiucLPWcpLrwlH3mql1iR6lBLiq1bokirUqMlTnaporCfJIkgN/Z4w7e3qvYN4sM
AieavWlCC6qQf28wY791q92Q2l8z2E7U16/pmpKiNg94ujsFfxeU4OWkyCOlGD+wnHv7v8v0F7QX
/pcpE7D36jSoLVH5k2LVxDzR1oqWsK7YTCdm5NzQ6bkPEewT8ykKQtHg25+jNXSiOhhkhBoUDPJk
OvS+OQ8o4lkRXKIcKAzfiOd19g+LS501w2yUTO28OSX+UdXNRR5oH8J3Eanul4D0FNsSGTxv1/h4
FXCNG58YI0qRZEFsiIZAA/J/ybh824u8J4FPybAdH64Sv80WtoHykdAP9b1jRkQ9ln+mgJQVzrsq
Ib1O2sEXxvkGFX0seQDgXv4B3VPNo+Gwp1n/K2cdGVhz4xcR6kW0yusw78Fll0ts1YWvMWDvgwpI
JIBARhos5tVQsOivryRR88yZ8Inco+U5Jvfm1IcekRFw1qVZeJMRDRUBaGxjpn/tKWv0VQCdkGv6
Qq1JjI+1K9lmomMULp6uaiNjpUBNpP74fjHgdtOrZUZl+mGpc/9gRRVC31EcIgV+6PpafrdF0H+G
iOYVZAVBuueFMVmZjYbmI4+N78S0SJgQN2oe4W2MeWmkb4bu8OhlYX6AY9O504I2KLtOoB65oa9P
WYX4qmvyZ8Vw6RAny4jj7LsEFyTDyG+JvYWbl65IYw4zC8pSZ8MtMqHC9OujMKIdzUSLUm93xcS/
I2t59qRjyB5tt5EzmmxwNct9cNPm+wVFgkChAyL67Le/6dRaPBuAhntAyU7v+YezKkzkhuqKHrkk
vqwqXfh7/Csh6bs8j3+7jmMCC3ChYoP4BPDCN8UNe4Apn1vuzkesi+ReMAPVTgr5dRcbPXLPoPFg
/ti/pQGB1UvnFQEXioySSLbjivzfDb363HIeu+NC5Pfdt8R99uTPfJRCHPwLpCS6yP15EeIpW+17
7Pb2yQ8IMZhTic+/qvqVI3NXtfUFiqnpXm4URWej3u9EF5LVjMnDCk2YfSClHMqUu94qPAZ5FMLY
ikSszgs5YZsgd0CJTpEBtQzHYyn0doBlBjZO9xfDnVUkkNBf3UvpuzxO8LdTj0Z40YZmtaZmk3oJ
MkpuEjQT1Xv2K/pckNMeIdGKYMdjFrtkRLYRXATDqZZJ4Zt/Zz9GZox7dxgFD7L4JfA+u1Egtaps
1+Im4s+ob6Buu81A6CAKPU12Vn+osh+/zfuQOKlZPN5S+nWf7IZt3eWsHzyzui4+P8Zwx+PvmnTQ
U8YtkUJqKoNY7uTvSdTo6ju+WHHTmNYlpXPF16z81OpfCUtci66iYA9iWhtVd4V/rf+kHkcPiOU3
W+gepVHQvlB5AXaQaimfipdQNwGVaaIKjPUeVmkh0DNzLiOX2clweWp+twtr2t2hHtJGW8vLGrHB
MppmozVAAotuTC9rGPaEQm+ax/1+VI1gUFUzeHTjDMcamBVF1Cy7s+s6/2762+w92H4Urmt0HnBA
7sAsJQziCl7Ioq/nHCd531M/fZkVqWrPXJe1RdH9i6ewWXeAxKSHjYSxr3GTgovJB/m2vTxk+yc7
+93Was+t+ykRd/Rcfbv0s4zheF/mvI3HNvA/RSCnpCXNaPF2t5XOAmZxNwsusP+iL699I9HdMaXS
mH67Rhb3HUGkqbcNhIBTtd0L+3nzeE6oLkpTVFoNdVjf5y7E0i18ZfPikSKgFLlyM5LslBeWMr3G
ohGPkg8RydO+FIrNlmkWr8CF/y3HpLKQGflOIAPPlAX6HMUFAoHoDwVRI3pZDWaZIegCW8a2GE/O
2qaWnubUjbzOjGDHdQHECA3uvHW+rQ/HSGtdU8XLrhoh1zZmxwTJxz9JRCydZxqZvz+7coLRTeIB
wWjm5nuH6YYAShq1tSo6XjXksF6i91FVC4YdPaVrQifpOe0DNeiP1FxA8tOejdalo8yFxVj/aYKk
zY9JOir5ubh5Nqsp/HeIal4dA5PX2gS5wENcfKs/sQlmY+SRmPu9zpv1LZZFJVN9DGEJQzv0fcHG
KzUXHnYuK1n2uCQ/UPH6ADPEIG9EXORLwT3oCYdZ3FijdhBesIxkBxEAQpYF5B71wOE6Xzwe82wj
FMn9mgCoM0AW89aNDYKncbKcLSdW40qmSJykqWQ8kaFeuTy7McCH3wZQAvvN2+Ue4ndeAHBu748j
bgBmPM5reToB176Vt8Pu9VwYKJd+TXvo8eU3GC9gxjGz5rTHt0wMQczy42R7r38Vn+Z85dB2fkvT
P5DOnIjDMC26INZkbsvgwjZgpXHSpbrSTD9Xl50cCXxIHYAgNErwgXRnvGDdsho1hMSt6BBBQRiR
Ctx1P1rf5BXvqfUWjDskNd/U7ZGrRE95lEEzWxy2OzL5Dv18/fyJTP6FM7z10hDLD4RHbiU0WE3C
tvZA4ygBWORQy1+XYYhO0Zut2I6OZ77JCI3npbg3OotyKuERckBzqVIcSE9W6METLJwc2nVXhAgx
yd4apswirtulPnD12u5UAta6WcDSZbzZeDGHm8r/ctt+qyqQeXZUsKc6Kyge92V2O7CNW64AfzSm
RgSbc08jvdmLlZ0AMGWcvIPPWiXoANh4E5IODd7wlNw5LscQvMaLdKoW2Lc4/xZCqan5nbpFk9CW
rsa++3fITi8u2J/Mu6bnI7jJjbphhwCybMy33ePE8FsXrWkbMXT7F+p6X90nyR8pKJitof1srvAW
6zqsWUnrG8MHUmXD/Zg0nahGDVyBG78HGpPGcizGvuvRnguBT5nVdbzdOGCJIy22sgm/X9C8LuvY
9aTXp1pLVXFduZZ60zBMmg6A7WME65MGPfaIi5EaQ12vf5NOVzZ8fNmm4eSJP6Tvxl6tlO57OH43
bvD5qVS+FUiDmG92LULW7rVMmq4IECXzrwnBjiq1jGopH1c6IguUC1IRbUWceLGKq38wRqyxsJTF
dZYMTejnB876WGgBPyRQG4B7Mmb5uArLwn6W5iqF3CfuoC+KlkMZSL6slxmmY4b1LrlHK1rCl87H
1HVP3EjVfpv8KI0acTSrle2eHiiqYKssKVeLYlSM6X3ccBuEjXqol48qHPMA2FzDGpJRC/VcA6AA
pvtRiXHEPGp0+MPBTbCdeYPy7VdyArDK6oVZH7wQ0Gi4KwsAb8O3CvGsd9f5doHrR+jOJhyQNNDm
E+hFjDmB6QV6if1cjCXLNdI6bdFwN2BaPXGFfnA8sEMHkZDGdGhlU4VfTnqQfFqrpmU//rJubQDH
haLfmCrmxISJFfVU74GzRPjxvEr/aRwrdLwxR5KPclPGUCx7ZKZLwP8udhUSteNzjq7sJkpLusE4
JeJ60antKex/YJPyKO5bVc/PTRxguoQ/3wU+GPDZN4OqOq1hWPJGeP24RYXF4VSC4TxQIH98CuGL
2NnTprDKx4suFT5OyFI2WRvukoh2ROJFdxMKfCkDlWp1lzFEtrDm3Uvsm/tAVH2mO9c6gxkY1x1z
wd+4G75r3s8PS1f98hNE90cvixIHkEU2p9qltN62Zsk39wFS5Nhn9iZO5s0wtfztnA/nRT8zqWED
UzkMi5FZKtrcx5PJncVRwRPpDYS+DSIPrEkRz21N22DgEoj3YP3Xjl3pCDX7ybE/kOnWvrOyj5WY
aseWUi+7KXkwV9Pp0P7fCpp6UryuX3TJI/+Ahk5YFykrA7Cw3kvUR9XfajEtWjE0aNUlWFJY42dC
Y0yn1yipwotgQZ4gVykuZLEZnrRKyJ8wGaVKN4TS06wv3bPqVF1P8jNcLiVL4OHi08SxSO4Wdppo
pp7VMfaq9jH6sDMAsV6PlE5Lr8YNZTJEFyQRpBGBSm4d4a+yJZrT+UWsR03seIRc+75gR9PT6VMV
N0CvKaRehM6KqHThyKEX5UA9CnMbj0d1oQVcLPctUehIuYgEuJeOtrtiAHUjM4Mk/EUujgeHW90i
eYSnIBSFNu3SuK6a6xfngo7LIa5QDV+/Cw0+7m7oLsjFNki/F4mzedfA+6FGXwDTXwxBenpuVBZx
6EWem2NBWITB16odp1fekFbvCy7y9jfs3m24j3IKt+gPtAQ+qYA1CxQ0S++kwTjSmszQX6CwLGsh
TddkaD4Y1dfU/DwNKS45r5gcTxrtlKvhd9fhl5VsgxAzglOyrXSdOs7iEnWGfGhypVU1kBPHetB3
RAS8RWoBhS456Dr5C1bUE1jeLNDE5mWrINJso/oDmZb8iPiM8MUrSnzp6kG4/DERfMTdyK9s6/oY
CDWSYH4lb5Ye0J9lo0kWq11ztQACjfpTAU1dJ0ZEKoZpWLs7kwmSzF14XD6pCzY8CGDQywZVchpc
IW+/jhcJP8gndWOP58oJX5Mw9h7O1dIj46qDsU9WJ8KYUjYEzUDjtSIktsDneO+wSUfwoF8YniKR
OZXqmNZkKn2X4Uny+1DuzYJ8Zb3/wwQWsppmgBwrizBQex0riX8sTtjgw3jUhNzXqn54IulXNlYN
PctryJm6TCrbi7/fpL86hELyMPIxrptmeecinz8Lw2yoTCXy3a1BBNTPUPrzrX63uMLfuk+zGKFk
/cF+kNGV2C1TEN1d5Z3hNYCipZZURQ+8pK+pNkBgxJRT3b9Z5dt7iKY7Gk3GgNMyQFFq7b+D4DAu
HDf/U/hrD1dENZiBsepZN4DzeXCSPRWf9q3BkLo4wyHg/BWTFAXzLQqM/FAH2LREBJe9dy/JMvRG
zCJRaJWoiPkYbENcJEYb9vV76GgolcIDc8RpI9D1djlNYKXVAsivXz+5A8nNdM5kXcbswoQJC9UK
9/2OIhRBbjLNYMQNvlw3tg7KcOaoHSfnXzrd0ib03yAuz4ii8pf0cd2yeT4PKo3Z1SvAAKCH5zG1
Sc6q0Gl18LdSBveXtWvQGCVf2GQ2ONPGDD94NEL9n7Laz/lw6XYaklnWPtvKpYLvYZ38vnugSlsZ
/adeMt1nj6QzEPTrERvL/bZ3xUrLHq1f6RmI4/jmy0VqF9U7ZgPl4AbFcDfaPYyIc10NksFROsaG
YipN6yDbUjm1OugX1LRXE4IIkRzd64dgJN7GJ1cce9valQWPmInNF6nbPbTKnoHvu1cwcMst1f9m
Tpx2wBWlOPUmzzlwZuKONAUFEDki8T/nHHTGg039ngpEo3oXkiQ/9l33gq6gl36d9zVKnyFwdUFO
l78auYOExJhsQB6xxY84s29HSUzH+J6Q+kBgNeOxRj/X1iCrJ9fxpeFceJbSu0AGAqgG83uChQRI
4V0TJ6BTizIYVixh1DM9onpD1nBqXW0PVhP509ePYlyJwBnc6reP0y+JD2X7NpujiZm+8/ZGjzIl
OgiFLfYrKQPh3IVI2Upgj7/N8FbwuSzH5RtI4zb/Hi9lum3WXLqSzrBHnOTu7/eTRE5gOZoyHABp
YInHnd4sB453HP+bF15OB1+U6YcHIsRWeDg6mEyYO5Y34oRn2BRXKUcpMzWhHAE/DkyfgZCQiOhE
dHR87JgspYIL/9tf4aQMI0XxytrpbGsYjvZpjmuoLyD9z89/J870WlaE50yLxta3iEI41IJjCH+7
sZNHNGyR6wNGk3yEfc8NV01PPkQC5g7KXeWFMKGQcFGsPY0tbW9AqXQZJN/qA6ZjGsO1ARdPVDNq
jwDW1Z9Mdr9WHJFN4Uhjkku4OzWWz+5MA2Kz0w0tlwGaxn2MB/Sd/4CsF+wJL+YH4NyUA0dM5fob
NaYXLxeNCupCZheCN5WKTt8YDD/SGMKIXeBUJrQqhaellFmVec3c4K1T4gFKh5AF+ORpg0jj+Dc+
RTUeQufDmEX8gMavK5xzrRCxFePsnhZwu1p6ybEExTefLnGD48MSRhH9uh7L9TdQ8hMZPZwzUxk5
lobjCmapjLO+XidKHYAhE5u4HoXZna0G7wNjmTnjcgX6B0l+gB0ypdhby+ZXCLg98lxiu62a3qWG
yhNODpUymq46C93DKxOonZDChHGjs0fcFihWejPPAKIQaRju8Jo8H95CoSzkZA3jaqJeDKR3kIP/
C5txoKQ7asqOT8sYQLbe4uuwaNu1cgkCL4snzwmqEtHeYII0dfoC88wLIxL3wov1VBPnGK9dj7fA
tRuM95Z1HOAjRmvqvlXNTkv1C77af8TQifbDJC7XpWzmnO91afk2pJZX0WsWuL7eKl1+jIC1X/4d
iddzgAwjtkyqhQr/vQb6lb2fIxHnRm291rC9gVpVCw4Qg1bOFSsj9iZE9bunLmitT6/+8xHQKp5W
wPAF/niVBOlqQ4nzdwkoNEzxfPq++bB2JGBZOhu8eI/OO1Lc/JO4o86MH3LZXWHmbLTwCIvsQrk5
Ar6lfZdUNJaenWLLw4mAz6DBygn+ms2AAfkROAiScxqRz9/GS3QgAwBVvTiKiCdusQfUyTLotToR
H2DWPU85GoISEoAi1Rdq39PJHY/AZceGqSLyKJ9+Ih2j8ZOwbeTBKBSmCSSE5HzQ5Dajqzv+QPgl
l++xDGua/ih9+lJ7vuCGPDfStd3CLI3YLh2+NKiZYCuPX9kJ66Atz7EXfJ2eM8EhZaLoUt+JfwB/
fkKxxBUlkSbWlvqSTMwsnXf8+Y/eY8iEXOvgUH4DbGVsIm6gJxroZK6zK6+2Uc9pUDDSPg9/x2kz
YW9Cq+m7J7KzhfkQRmZotGjejtl3EZe7+NwQDnN654wPgYzKqfzq+v4yiiC4AFABgMJSRYkrvwiA
64Xho+X5QIozcUX1t8hyR5Mzsnb2N8CrHTyzCQpA/GoU37Etws1FDODCoc1UmiyKw9N36K9xSvup
fX+cRPy8IPyapjOo7ZlOFx1/3nj/f2lO91ABV9CK0Qc84nT/rCAfsI861CMjm3GdS767v2A/2CF8
o3/ZKEAaKe2QVijGCmN+ZqH5me4huT6QhagNA0Rkm4gZDh2j5+vOqcsrCMuZM8ELAG3BUiPZIdHS
thm7PctArcC2p36hz0mmYdiP2uZkFhA5WdT5nTyobVfrWjsqv+8ea1s1jQYBcWCDSKx1lBPclMCA
rrTGbVqa4/2lVG3Lg0LKyvo/v1CLYhG+aKWB5IYu68nqqrRlVGX+2+ZvllSNcWHIeshdTN6IraDH
M1p5maCG5j/5D2atTeZ7eLOVcRistmzO/0sg+oh146qIMXqeTUPPNnqH0NBhwPdiYq4j7ggfBbQq
NnRNhihTsDJF9ubkyXUqBNlF0KMCxsYMcVPAEQYobfTQGq6/o0dcOnQ7cLIN6O2zYeVd1H1ATzki
GZq3/BV00Rm8Aidl6TLVix5YITWisj9iJttRg/9E0ZitTiJMLqB2pdjWaCbubcKueQYtTV1OiPhf
ZN+JENJINfaBWI6pdav/dgcnSB0vIpi5ydbkCLCB4PHhql6g99hL52Wdlw1bRQYhzsGRIa24pc9J
6wX24imI/U6bRjAzeGJcQ+0mhvzCFDpI1kUiiYgniVuRkNks8mmg48CvC0hKTu0bLZSQ4nhj3XYk
SWn51UGWpOF2Xh0P1eoVYUf+jawUlMZTHgCh5ig04Ig8i4O9q65NpOitpuiLKbMS06Qr1nseCGVI
OcgY0nmlXeIR51kg0LJinoLentCeWSN61lZPSp8KziWR2BQvFZefH7qoelhTqjK7pme2Dj6xjOgz
1xjazSUqc9ULHIW3d3JjPpPj9HZhT1NifQFOaj8nponx+DdVEig3ebZOdKT339NTwqJYsPMq2S5T
iaTk6rmx0p25w1tzk+QAirYa3zCOoJR221W6CukAJNdXAy7dnz8fzoac+dZsI6Tso/+DTUGQouoz
ktS2SXtfMJWe6BgMqoFg/gt2FT/TlD0UaKADDndouKLa22EJltJWXMHbDXI9BVoi8eijQ98OMoNN
49o8PPDl+r+x6zhiCDd1HM4fmpLZIVGdccIiViNvBGXx77vtzhJp1W4UlxmlbJsP/nJudgxzC3lX
emEnax7a1rgk54Bj4q7ws4bmY8XolnQ8WMVIubjkXwoQZWSdb9ElzqWyC5Fsh3xFjz2TR7/67/wt
FUYOKMEOcBXLrXYTiz8dwYnXUxrymnRUUEkKzXOJZhvjwvPeOphlyA1KcJ1yaOMx7QfAOjmhrhLB
7WpLJslncoXg7TFaeRWL19ij8ICKzkQ0PkRCtQdv/RmHilLSlF0HIG4VkYQ2ZgB/6wJHmtXQ4rF+
mToXCKbUZpprkmYiGNZCKzRUejINUrhCiXN4kYg8q0/IWn8KPuuMs1pZ/4z6nnmZUdUJzq0drmy5
g2tjBY7CtAvCCUucDb46Uknhwu1Mv+p5YoLtqPbLAv+oNAqGIvg2+Aqd3nctOgq25pLQYJRPd/vF
uGvE33OVBYw9gbCXI65FcOuoF8XSPIGqc3LeO2tf8qKlQdDJvOn4faQerV7S1ItFWUjd6382HfQ0
yUR6tV0f6QJKUvl2bUKICSj0MwV9I3JIF+6KzSZa1s8k4xWwhOjURQXvASrhvEMtS0POasn1Nzhj
xOY3/6qXTTxXSEsvvmmdRHc/DQS35kqxfwL+V8Rt6GKt5trM/MhLhA1MYAkAs8HGagOPbPPUJN5j
slQxPfaIfDWTfIbjZ6KrZO+SpeLMPJ+ZlspQlhWdXJvuALEXQio857aQQyrL0N7lVm5OHxrQO+h6
l5q3TxZ6LQzXrPr8dp7zIHD5wKyuB+xDT4u9R9rH9akRGgS7IvMo/YMU2fjLbniht8qKT5Dx9bF/
N6KEBoCzN03EQxFUl640eiBChzNiengI/uYh4A6hOOyLR2Del6/p4yjjBZnPqwIa2w/e8fnnrLqn
wFOlJOMCa+pyzI4VNTqesJ56eo8XF/9DhDxhQfmwaHVe6ExtR1huWkuWtEOoPVlHAf0pY4Q8pKnD
yN2tsNPJlsKcehsCfrXTF1G0FL4ZoC9Tz7gdzKXMIUUSMDZPbnnJltUH/NN0qhD769a1/uK7HFrd
TrFgqqBI7q3uE7FtooLD5CFAR9s4P4Oq62yMnBdC8dCW40REXj8/0kjmxtu5VKhWEjlW+d6zf3s/
zn+3Z4kcF/MQv6iWpiA/imxWAsW++uqM5a2AZV2Tte8UanCtg8AK+0F3ul/0gdFxCjCZI0wo8bA/
b/H4OyNsHQK1ub3dd6hmCiv+T8Kn6/90I7kCu+jxT8Lq5UlM3pwR7ryOjx/MfYTaUpkRqHLvc7YQ
8Jf1wOJZi+n4Bk3QznjVHoorDcpkrDQ7DEPE61gv9RhKaDfZNKxCp0HwydiYA/KquqACj+Cjssr/
bJWEKe383ivoA4RD5LcCAVR7yL4EjhBcYYKu7aA+qLiE8s+nf3w/LANS3UB5d3B0j6z+WsUY8Aj0
xwN0NPtN5Wn1ATboHPyIAGjZnQCImLP1KgnJE2Fn8aDmxHHeVbMB2Gsd8Xypqf/McsidgHv2ctrD
JPQw3PHDNg37fKdRTSScBea0EA2gvxs47o1/sYrrNKFfmw9lFm/QugTroaf7Q6HJyORgZUC3j2I9
Tr/U/aH3PzEgSjo6AtfmSU613MpJpnzWWkPEm0iF+RVoUzYNUb5ehFymn/NC4MLv2p1Jy00ysewJ
vrUPIiXm2uuIO8SAV1HeNkO12bPMwIdmStn+XB2vtR19r5HhcnUteebmu3jumzyg2Btt9nwmZGc6
ncya4ExW24ifvIh+yp+wyIC9SXzImE1+nvvRdNfyYKIRcPsTEBAhN141Pu1yUrS1Ue4atLq0ZQhf
MJy5Wx2iPKab8LaipAdi18gkQLxlYg2xPt8M7jFiXtj7k3Vn4icBMUzoe0bPwg4lbPlXXmeb4Zxx
UHS40d9OMe4Hp0zfX50TBSK1EmqcGuamT4kVUhUA6oV2q7yHYe8FjaPRF/i1rxu1ivzJDZ5wGlX1
6zbr6YGr+Z3af5xwLszIUbFVJnLBi8ufUpjFPJhubZlwqnyn8esZVMe1G92rhUamWCzYwtTRoaI2
+DoVrvxKs0mqpwz8idX45yQw74hHdbcCJQHhbGrJlcjQyvx0fsCwjgXFKp5tCPqWse5nsbRH7ZBs
wJP/x7Qa2sNRf2I6Xd7LhgtD2+TBSq9onYs1yfH+HjSyDEkXGnKklbSKU0c/Kckr5fB4lTSxnj6U
Xr5W2sYFrmAUPtb9FxcJSQwyV0ewh3xuPHkhjbo5NnydzHvmt/na2NjXZskmaXTJwe/I3FaOMe1C
PnajGKjmEYVnZXXBL7c7+ngscG3my2OLtcrxB4fkrJZulX7fVJ2wMd5sp79+Fda/lU1/bCqs28gU
imz4UR7tAaVSjr7q0bZFqqzW9RhRL4YcSTaqyL3Qd/uSJA4nTdWYf8Wyxvr4GfGEqsOeuYF+g9rN
ILsawZAp3MXr3xOoXfsYHPfYPdpJgTWB6LpMtNDg31LxIc1MYTHxk0lSzI4+b1G9GsRbHavgDw7/
Lgnu6zJmjGCmkbh73ejkVh2L98cPsXC6YpiNdfW4XxX316mAqDm0kRAzwrzCR5ywWzMESz7MnZmp
OUl5TNmLJqEvkI1Zv1BrPFnxd8bHRWvq19r2BxnNeTXeCUykDxveIoRsxn049/PM3mLrOTFkq8zA
GNKcH4Kz59fxTDhCdqfFM76sL8VSt9ucfqh/TDM8VlZUy5j9T3Pjlrmegnpy3tG9zDawUQxbEfXM
SAUeMntPEasadRZX8ZkmzoL07Zh9gt+j6A0vJvJsD2Cabb5tgakW+AVVV3lnnw4hHFuXJB511qlW
Fgy6Z1GTnFY8lnEtKtJnRtOmHYVqsoQLYXU3tiGmrXkQYEVhPG9IYYH5tXDYj4+5PEaOKDIJ/D7J
lTxr/OXqiqT7C0kRiRoDeY3m3XaT+TStvRASmqNxcJfe/xLwVUTUoOp0VZP3Lt8z3PARNe0ty/Rv
MGyIqXsqXOTOEBQ9Pyrjz9rkL3NQjCf16BFJQm/8sNzB3v7EXL1emTsg2Kt+CN2DJ18VtEGQVzYg
17R+NSEZPBATIwEqVNVjOKfn9JEI2n8zZ2TDMvgK3V+eS01SwFNCCBaNIIvJK3YIYlML56nXEuef
ex2NGSPKfAD7i8xrFptyEMF7F6/LVUechQyeSPFaWJtcBUSsbfjtcowecA3Fqh9c87vpXgf/FWEW
dV6w7QzedeI1ErBWIs3I+u65Jwj1ejobRT2XDw2qxFkvFda4DSGO7L4VDPViacSuUvQRjUhv27uo
7O6etG0K6eQsSNLuXZw7zcd/r7NGbQJ0R5vO7W47XN94MIQYPyx0SAjmZBhympv+ISo5/XO2mJPz
e/54GdjvKMMvITPbrNNB9dnZCyafzOSErHk/6enOtjjn+n6ZOtmC9ak49M+AyrmTWGY+4es7NUaa
9owbpADU2RpZ/PHJnC3ajWRi5Ec1Mn6USx9XN+ceKudgnW2WeRh8JNZupqDzL5Q43+quijghKvLE
9YVgMWYEmk6Phmbt9/5HEs0Uyhcb8mS7rq1ooV62SegLot1YEMChkinZDFYcCPDDy3ZtoPGCQ79V
x6osJWrt2H3ANIJxIV5tyyxHlMg135yINYbnozI5fPG/B1LWNugBbQl0s940NC4tK9Je1KwN/mAS
vBrnSG42FENlCSDzCTdPIHtasw+CLPNrPhR/IAZ36mQg3zHCe2C0mUsZOpSSPCdr8CWbTcU/a4/0
bbLBrJP/4/lemmsBxWDR+kevtIXYqZuSkvHkZI0vlDYcskfs4wFK4aXjknOD7BSrCrtP9aavXR5Q
oUt8//a3+iQanSbniCBGWg1lbzi06X70xR6PkIk+9SRmPYAlj6t9+UknsSiiYPy36h7z6UBP087b
rAB+QSrEWqAkKmk9xr1I+gTNveYA2/FBI30FAeWcjdNQohq+i58r4+lcintlvInyQ7oKTSGWr62H
Ls+7gLbi4ALQk6FHktLR/2DLNwSNbm65Mg1bC3wnRIN27Vj8osFvG2mLvfH+jgyLlJ/L5zSwHXQ3
vh1rzxw9rPyO2CydSoux997RaPqCJYF4/Wo3oevxnlBmpoX+HmImtFpfZiCbeZMpL3XB9HTOqs4K
a5cOh3BJ99ARdlNua2btF9SIUhB9w5qnF1WfMnzupi2Zk25UA5WpytOlA57ZrOA23/fLiJf7lNLr
9oN0AV2TWwnGvi4nqn71NvTEZGFnGn7C61PwHN9+eJsXWOah5YSz27o2vq2xGuegYV36wL1aDICN
J/VmDHR6byyGBPYS1/lzJKnayaMJJ3B62GIeXxGFvMmVi7xKY5aqg3AdttqvPZ5U4JHySmA5QNP1
tjMXVkoNU/9FPo//8F4NzY5mD+pEXYlZhp7QAtyiIWTd5lWP1zQD9qF/pKBZar3q0hFVGoYzIxix
qceQG69d2x2lmnU6fOtTHQKfLS3qX2HYY6oW8fFcqVE90XuMPZa9lcwGnUIDXp5xvnhDV3lY03oQ
rjkdnDBPEkYMQE4QJ16sBo/TerCjZRubGE/a4RUIVTQxMLhhZ4s/RtN3z9CYC8AAhSaV/092ISUE
bfyhfaL5WPBQey3fnHDwK1v3VMBMj1o2yB5qVGINHhM4Q4FwD8bvas1a1v3hS5JFQjnM5vOny0Us
qGjjPN1dQY4W2MX+k/+u88V4qnFFyyOfv4zkNoj8zYB3CLVLllTpaNXPNMXxsh/oWGeJCD54ToE2
XOaQyR0CswkZfWrkFyzTDjUzzA9kY9eGGKtS5Cyf5maG71Y5PR4B6Jwv3yx/+uDUyAB2cQPr6fJ+
6r/dYP6umygnri5pySl1Q9U2Rqy/ABofBBHffOvT1xS0LZ03WiAvAqIS1xqmZOIvl/OHQ3N9bh0k
1g7nfNujrIXuQxyj3Tovl0yRqNcIsAdwPTKNAb72lNnYxjzXUn4W/gQSTgnU0DJ7GXotvY9zWb0u
kVO37FBBVjVfb5i+oBAOrDwDS3tn/Bek5SxbXwDzPdU+sO+EaM9yD/KyStPko+cRguyBx7TFRnQF
+KeCn393bk5ELB+IpKrVfxPGu+qrBZLqZokFLa2VYyqpkfY5a4zraBMfakT9zLOkNMW2UuC6OAGm
kDn9vrZd8K5HokHAHmAzcWQu4DNK9fqELkEafoXwEcxx5rZSx1nkdYfSqJkbniZ8gMlYc7Fn36MA
RoCG4EzolPSvZtUOF1t6tj3YEqtN/reBYOa+AgJzzAApZvbU3L/ZkJGBN8FUuGb3I8I4OL+hc63K
7Wg9BnSUxX+SLrNCr6FSNNHAr9hDF2FhGMWaat3Hi6dOI442pH2yIHWhvgq7FtEDUU4GVQ1wlQvu
DGckCup0EB9+8xcZiquYIjCYUMLO6o7MhIpzbU8WLmTwtW1HQYCUX93CTOY1QdQsceml2i34hGF2
ZYnu+AeqsiW64fV79g/UP830qi3oumvYrn1MAuFUfSHkp6GJRobsn0nHXqdwLvWIVYgOAB60BQGY
QtXGf8Br0cCNy1nqbTZ17cqIvIeGNasCnOhnhDcVKEhjKuupSIPN+4KbFOhX6Cib9KdQYz6+XzeM
XTIc50y8q6PxrPgt81v6DsbjLIZni3hH4NxaJFGLAoo7Ah+L8flJiJ4Rk9iYDsRP9QscYAcQJTgu
t3iyDdEoH48w2FnjqlcANsqJOwkG7LSitf5wmA/IacrKgBceXS6UTiivMTdPHwNjbM5hCXDiJknL
fPDMXuNgh6u0r5CjjKC3BpCQDd+HHVNKzr1HUn6dDu3b4+pSORtPHmOLlRva7D5/ApmhP8tS1d0A
1ysLlo+Zxq0wgD+FqxdYMfbb5Wcz9+wnHHOzPSJOfpEILWXfQWmCtusR3yqD54pTHRMKFMdYs1SQ
vxW9JL4H9Ezh472sd0PE1kLb2IwSiGJY3KYCw1mQwRl6gzHL50GRvJxI5lrpAaT1aovDyKRIZBs7
Dz+AFOOeEUeF9GbhKIZ0SXVArFfCJYhYgyAaJ9FVgTHo2csoy7SWGU3AQbJAqF2KNryRXrnxMoaY
tcQ9dHJx/KM3Gc6wyfE1XHzdkfU1ZyaHKc4t4+SCCdSc3vGUlY7lRgVY+Ex85CJKIX7MCOMILlrQ
HES8JKfGEUVHplw5MwVq+Xole8zIFoOcim07j/2AmcPqboVieKQj99uprgEakC0SL37csfDMS8KH
QtlhcW5BPreB6OrEPdKf+hQ0rMtnBi4V8bAdD7JheFZjT0E9xd7HX3EG3YMT0NeFd5gM6m/g7xXz
bZ5ei9zndvTCdTbJKlQxce2h1tDIQKDX/o8OPpZJxxz0N+CUgh2BlO6D23+Q9NqWNJGcwwV2yVTQ
9EeX+jp4F23gTKSR7/yakNkOHxe6aP0pHDpfYnM3wB4A0V1oMb7g61vZ7TO9gh8NeOG+8pjpEnTg
9Tspk3WuaBFFRqhWPQJ6y0CC5vZlGKyl7m1abgqQnH9gKcUqd2naJt1PJN5PRmktGM6uqzpb5mYN
+Lr9NWfnpUEV4Qz3HFNA3P1x5E8nxxB+pF2gB4mKsQ31tQOb0C33rPQd5SRiL6GviP18uTH+9f5m
GtCHa1+ZCxBmT83u7X4SBu34gawZc/Cd5RfNXzmFqXVUjOkOpAuYZHtHZ37QHLxf6yRUE5EPJpXW
FT+RFpBwzwSZYVINw9gtRT8GkJoDBYXg1tuBOqhGQIbXCGTy19LGmdhm9S96pFWNknbvTVIT1NW2
a7JjVJM2A06w+5/9C0wwbz+EOdmVDLR1yf3uSHHebJRIMIih6gYnVHSpAZYZ3NnfCp5AlhViGtte
S+OTJtfjmN+UxC80KH0vmHpHk54mvSKbGQWQijp7g0C4kdFxEeEPnxoQZWdXsFAFIS/gCgd4BIyY
YS6pzt22K4sbtiFkzMKglJWiz01QjSjocQdNZzc3TX629xkmZW1VkVBXZwPtPl1sVoiQv5hiUlEl
+QfM1zlQZ0oZMIGFFqBn5KdIJlqnNA8RkQcnp5e7VJHatwd9mSIxWmyoZBWDgA0TuIO8FINp4zgS
MbmZspb+SDb2/Kq+v31JYoTpu0195s52/2+tXjqeXFNfSw24VoTJOWxRUhC9zbDpRDFspYcSkl6o
/r/3wZ5SzdqXl8oX1qMpyxgz4V++90iHfrEdb+AD7hTnOrkWvlw3JZ3tg8/kzak9+dJN5RT+AkVP
V70XArYMKybpwop/OS+YZctXbfkZTQ/0QCSNboJcPL2yGSln/Ory6z8HzXsF/RHdExBq0OmLSlqW
2QCPc8qxQdtNMSiuADMFI3ivMn9bmgQj5lNBiNeM7uZsBdNRgLWaVUooYt0UTmry4IrV4IYshSLB
7ZYG+a8o26oPf2g29MDF87MEVa/Bv4IbQagn72nECGh4W9keKHgpiL39Kp2t8C7b4DRbpEvIfYFb
ypGPQkUyp0gJiJfrUum7j5eQV6wEF6o87XH9XiEKtQWgjBRxBYjccppzZWbatAWE7FhHuI3W7GZX
sZLCp7xCV24fPhDcYwqpu5bbACk0RqvQgeTqyGahNIxWLvaImve11p7O6RlMaDATpRlRUI848GQD
rmcB4ua8yN322MaraFv08qNuvAIHFZDEHLsM1FUQ6OCfJHIyArTfw5+y4S6m4GIJePjEz+9EE4ed
rzy96qmSWqaLfqzqBtxx6bfdsmCTvmdO2kTMwJgyisxdY+eILsMnQ2xmMpc5WvAYC00kOg7vhzMs
EoQeoEWkmCvVI61C7CLD7BdLR0JqSH579yfTcEJWcw7TxkD2d8MILRpJQapCU/V8XIVEoILTjXMh
qK824l8Z7UmDR4ccRwcpMwAtLJjk/5kAQcUPmSp/SUqpXxs8HYhB6ppPsmfbyq1SOeIEbRwO/N5j
F5ydNqnhaC67m+WIJ22K7B4+I/E8v3eNdkgxxeDe/cItr7s87w72Vxb68aYosI52yZ4lG7qXSv6t
yp2Qcc0hUd6YcLaMTYBgUO/+aBDFcPuty/cnmeDGZ7O+wzZYKTz9XDHMwzafxN9hsBDYjF7nO/6I
N888b3CR0c1Eb1z4ZqAzt60kM2BoYzUusGoqOPGGaJJP1Lubj/ePBv7ig61GdR54XwcGTV0pyy4Q
khCl0z213P1qtdgsmrbpHiYsKYONLRh3PgvTEdtP79MX9jyAcq/ijbBCNBSxcGndK5EhTmYEffEb
NORGeIlgIP6AVo6i7PSQkaSvGedhu4aj1mON3DPu6khOQr3oKoqYV9p1ETb6BictZ8dnoDBDJS3F
LbYOC3Qbpd+iJN6d05xMk5QLHomK5usgT+lhROJjS9lH7wGJdeHfcjfLbVDugqSch19FUKt00SlB
ibXsqwjNxLEtBih1XYImMn2rvbNPUE5ZcYnv6tp2/gqdoISMeGMjuDJlju64fnjptPxRbPXTkFbp
TY/WVm4/1BHMvLYOlc8KQEW/xb1NDCQXDIdUqmf2mYGHj2b+costm7wlyI8xIRWet8yAiEhq1Rhh
/Bf2VPaUCB9TFNG7ogx1A7gFSiMBMut0qqnf5F/+Kc1o0BpKemAMOT4e4ViOV9uIjtgGW9DBLWTl
0JoxWUXCtPiSojLuwolTrDHpzaX5K8AMVfB2/vaZOglsCQ+GLfPz2CvtiA4Le23tiTzObdUVP5lm
Q9oHhjDkNPxkh5pplPQZaL7d0gTyE25NrUGcKBu3h5S563aydCMBSZU7If1xt2409UsvPTOnl0r6
pnRbSflDIq9X1fCtENfjkLbNRMF/nFG+SnXEEJC2A22nTKIZPENif+C3MVhyvkIYk3W3HNPoE1J/
alIeiOWOoDyA0odVzKStrW4vxn3cyKBmfhgvsxRbv714SfKAwJAkHcIV1jyW2CG1gcQZ8SAa99bR
T0K8VgZs8EE6k9W0xJBkRmKYrK3suo3eDETWXLFFBcqRW6tR0vX9MoXcsoW2jJywbQN8RWAlnPQO
8lbbfqdu0TW0tjOFyHpebk323F5tRrSKVlhnNnGf0bH6dXX6mKr18I5maRPWTMZ/D/QwwFGWshtF
tvaMC/1ZwTTar2ig8kdV7xB55TyMDkODVjxsGEvczf2+id+8+ngZVUcQ3TQz1j6VDWyNIE/Hd5bz
K0qiSweKtvIkR2/tfyg6jLNVdPpvJcI655fIaDLCUXWbZCJHXKhH8Y31pcCCzQn7FjsuFkPo6pe6
Scdbiaxuog48s7xykg/b3L23QFolr0tkhrBMKMzecGaGUrdkziZdWGkBYRndcQQ9O0OqIgj+TRs6
xxTpEAva1Vw+QPkaSHOf4lmcWTCG01BECSp4xvRFJ5JPJgDk0+mQQNIrPEN5ifImISIhL6DmcSJB
Udt/Y0e3Tjv7p2ew2UgfhV4G4OX3ArcHK1Ap9xQW5nV5OLZK1od8tGdk7yAVh95o5WV65O8OCoWY
j3Nnt5BaD1CXZHVxZmMoSx/G8tc4JhuPozZix3HP1zhJ+9J/1xIB+vPW1vosJB6x7vI8XloiHpDy
DfAPZ8VYPldytqc/z/5Bathx9EOLyLPptpvV5zyss9RypSA372h4Ys0dTu6HY/D69BSzSl8MIkzl
oJ/N/Hk1eBFxC8sPvI4Ot/t4gXPUmfwDMK2z23XhflEkER7GT4kaaxpPnwHb7wZPvztNGJywUbQT
ixC/SBTphIEqYNEXSjrlW70vlxRHKRVuHDJSA1+5cak2qeZie+LjRMUEsWpCHeheAncqoilEim+s
ngKNdiaFXD2c6ObIimmuyPQTAiz69mFtvzF0kzgbxmBEAvFFeLKToPTHLRc+ojp0ln33b3OzLgHH
peo24aL5hAWDY42rsFN5gEDBu/KAdUdWnhkT4iBKn5ai34w2xTeNVzTxzrSZwuOSnqp9y3Ppm/uN
Ds20HAH0rkKU0pBwHxVSkbdFKEzvU9K+4EdGJ8OjMy2/PM8CBwRYg/+wVhuaZtMY8C7eU5zBaLnQ
WIjHOrB2g0tup94ioaaTGenW6RCOZjl4jA2FnfORfKv5ML3tiBzPpsJuT3AkfIYwvWdf2ui+HWDm
IHqKoddgdqdoQCWXqcSJ7cOxgnepiHAsP27/ZCDc6cgkPBGftG0qeIFHUk4tUYWrZY5+KsDW6w7l
prrfhem5jLo1T5Ws6VXi4JmIC3x4R11JnIaP4fr4eQTNszq7mstNtLlOs4AGtVtilfjFKTtm00KF
6Si4vCHUILyBj2PZ1OU7k9RGRLUv88OKKcqnO1ps+IQ6WWRLXr1HCfHuYxktF7Z4sPLJnIiXOsBE
loTkY4Xq6hHaSNNqOR/m8UVKGDkIpMFfKnQ6uhte08id4swggkKvL45dZhsmobjTaX6KUZguOw0c
Ll/AWB+fCnMzWnvMllBNoTnVavIyme000TKIAp8ClZYBSrFcFS/YeGyJyIpsFMCY9s6lCOUu+bcY
ZNl8xuzZ81V+6dEBbJSUD5FwZVLqJruuNzuUFwkBYKGcDMTpG5t/aDjk5XOXfOlXjZSMvIZktH8f
mhBwk8zr3rnPzsWPD/Fon6ex0u41q9gpcZuhu7EjCDIGPy+iLzPm+UxCaGD/2q3f9/zU7BTq3OTo
MYOfUi3UJYKOF4KP8tDXRgDlgf/ZDHxz2BvcLyRMmOMA8Bg6JcqSGBENoYKUoGIYthW8IJ21c3FE
BIb7biuQFdqTDDDbuMZu7AIj/itAp7YawEyCNTdVvF81OTISAwd2mp3EgiTBDzvlD4CCZT9So4ZQ
v0SJdW9toV1+LyllcgvFV3tHu2P7BbfU8V4D05B8s5EfwxP8YFqvxqf5FXKyRxLNGWVCZQvcuRJ8
zaCLhvPglBJxg+2awWVwVzgPGwr8OTFiiwL2rjAlYaOvfxl4DbrLvN+Kwitaj328zb6YFJ1qyDwy
2TH5FHHD3piPczxkfW2jpVfWwtgNCaD263N65lVbCKMe1ZfwYDgn9RpgPLo+dgWvvTSptzF+wydv
1nvDutlLs5Jddqjcu7w3ajcjPMRxmm62GsFAdbAPBBKW+EyJziVm9Y44vk5EdI6CZkV2qtqq5Obx
vlz1O0JTZPc7Ln1LrVg4hUJsbqPeqe88EQGKg0zy8SV/Bx8MQBjurmoEhKYGHk4y+e5xexKDsQmo
SmOmggLtZomO291fkzXakQRY9NRcWP8N89PYmTu3amLME7sfgbmYGUGYbLKDtF2mAkmJ6zCb8sMA
rRUdp+o1E0y9SXOkQ6t1rCbaw4wQDWkQWYEv3CIHzDp48w59WYx4gEuQ2as9cSYhx2MLU5rvG9Ed
2w/Q38qBfprOMeXwFA0OUr4ePdX7p9oBVYqkip6GaVsuGW6BiVdu9LYvp+KOfJAeMuDkXY+3h4zE
7i+ECB1vpKnDYiKy5mVaAJd+wjZi9iG9B94QHpo1rRezdDzcb9aaBFYqnMigiUUXyQC81IWwwkMq
Msc1EW/7rBvZz7HYCJ0g5YB8eY6qbHQhuRGVesJXz5F7PZUnwQZehtomSEcq+zchTZXMlm84U2dD
Y7Cy8cPF8xh8EQyyDTFo0QZyuZaxnPMIcAQNAYw0074Wf5MqbQGfxDEDJHniUL++2L2W5wU0gfYF
q0ogeqjtncuUv96mOUDj4udXcWa3vuz4GrRqt9gjkf0NWMnabUkIkCQRExAKIJYiajNHzNyMbAbB
AbGpHjF/8YsYgfA7LKMn9RO2oQku5yCpBYGS6QHHptUDthgU7yhrvzUYaNzzCar/pSAKkc7E7xSK
Gp1GRizi2gDq/4g9XfRuPG6m3Me5XNuZA4M5CAJkUJclB5lWqYgGb8XrhFDC3MQvZUHp/7Bj6c56
cQ+ZrGHBjdA1ukuZUXEqh9Q2mdfPgpbL49CJhZ8VqaXhy+AY1nyPx068u230VXyZdDgqBKYfm+9g
2VolfU+Y86w7s5ld8rYu/mj369T2XC36uZHIzC/weka7drOfPeOL9TzqgxhCyWTADa5vo+oOtwQu
F9waKyF6p8f90qGtscOygjX49+xWS/A7bFc1/qFdZBI4zFkVKdvcQeurjxwxP47KDHThpM3xoVtK
iBXFqOzJjoDa7J3u8mZoz5JDFlPcSaP8KmY0tdHRDGtEg34dh0TCn1hDuQVXtQdvBjmU7ad0bgBN
tn7ESi4pwQLEaHqzsgfLITXaO16tUCgX320Y3kmj2EZZPn9M3zqBfI7myUlAGv+cnr5kWTqtsmw9
94JyCUd2Z1jF/flB9OpopM8U2Bm5u9Lzea5Tp4EB5yEMzaTFIW0Zf69znCFMWYVjZB9rrBEK+mR2
wpnwH783MmTR3YyimDCyg9eq5cNh5EoH8Nhg8LN/usltG/QKTdYNHdqRlhqTX3D3r0oZrJtnX2XU
xrjQzJ4qbDPjAoFINubArUH2sOeLBTxU/7NUfMjyNjRDe/Ficl72sOhKT0o6Bvhh/hBF9wlTrwKl
ijWuN2GJLkC3eWXNoD6TsC7FSeUi2uU3ZMrRbKHidE+87hGhrjeUJmRlR4sLf8miKGUSIVyTMymJ
+U83WUjFMHL3LZG6Vh2YfICkDBk0Us69SjccmegpTCsGSfcslq9JBpgM92MVGrXW1BuOO51BWN7c
2v757sehXaWhCiv+vcfxx6Rf3s7kZI9zaWAja8kvvqjMVeHzVJ6F62kF2zTjaIFptrxN9HJr5Ksh
htUbYlsHJKZv+6lgFq7GEponqyJNkJiKS+mn4Lnq5+UXbrklMTQW8MgPNpFlrNi81QHLJkyv8Wrl
FDEyNbryFCjdiB5iA1kcu4w6v3BT4XGrUGL3+zZsfCfr32bNJ7MTyLfQk3w4Lt4bzU/bH0Jcg4c4
6P4UIBwf9qIAjP9YKtSm6N4nTsz7GlG+hVP2alM2KNQP4/CeQb4WxsZ2Y5XAOo2vl6I2cD1ohhPt
so+GtGkhjOQ3WkTE7MHwq/310kZWT4OoklOpOmq9lSx1un6tITTHLtqa8Lux+oB7Eg/1lPaRK6KX
ZGdJiuuWFnYIw1bmPcosApNQaHgPTAm7EPQxq7BlpsQeCZIaQio8N2ERqUyoJJ8+PcQSfwK2RYGA
DEvAQfls3LxwXdqgHAifQrAKkSpuKfgLS/CvPD85xCDK3vCrcWmr9MbN7u6y0fT/leKcVWeh/R1d
BSFfIg2rjhp6DHREOpwJnYXvg8AqF+ALmkUTEFHWi0n+zSwEi3Hkv1hbKDEoAgCLfF4S/Si98XAv
tqIgZdQV3ElgKrJysTy0Q7YfqK1tJAcRRKp6s0r+4DYpFj6S8vEnbLd+msPZyDHLwhV3k2ty/WYy
NEy4zA8Up6p4ZIW3BdW2hMD/tl9HmWalBNMVSdEW2nxoMATq70gVoLQjchkLW2N1ICIXqOrlkGSc
QocB6mjGMpVjbnD5vBoxNyv6a8Dl7vEFlcxUl/Pnyasy/mIYGO3wr+1mHoGZP0TEbPYVX2vmG2d9
aoDXOKxpeJe9aBNPmt2dRnQIRhYZJKbLl2VJmleR/+yrOhRwwKczCSsccPABiQfyuinlB/hrrEaL
n3koSfp5ecVKzc4AeFuO+qOrMPxpjG9apqMUYfHk1GFSbS4i9lVpL5f93bb7XhVKXookpJf7PS2h
bAkcB2cJJwmMJ47L6VbR64nPoKzj2cLSD9PxyIqaStpUFYiXuT31u1Dk+iNBDx4lfynDmNR5sgh2
cz7D7AOWzThvC1mDYXaRwB3O2j8B1guHFIqmnAM2jXuAHX2P+B1wtZmS0BaiHZ8r4DTAGV+iYVNJ
NxMcoBE2KA9k3c+tBnZ0H1FcCmEnniVapNaV5ABQmD+dOkdHG1zCCNOoSBR7Qbko2ngWzjcrSL1x
SHW4m6lu/BrZx5TADYK9ueidtvYEIHG+dQ+gJGi+qV0STxQD0bQJGZO6FDt2qca4tC7dLHas2IFb
YpTpNg3AptEP7ysF/t4vi7uzgUWrMWw0ANqWWT+p+1y738OSu9Xt1gCaJlJwA3lADYFvLaz5Cgfh
Qs2P7mi+UdTUMV+YXspTO2z1l0yrkQnHnPdC/RYUV2eMWj+r7WPztABLMz6gQMSo7S0DoCufinYc
LOHon9MydZynsA8HDIJYPFY5l9FurGNl0aD5Na5Igc50Q9WYt2DB03/HyKweRF3vvQdBO2ozPC79
8uMhWOS2DrEIY/KmLriU85iiAqkZr9DlxQq2JqThpg1fJVyS8O7wdOVGKhUTgBlbcOo9Havwn7dD
8r93Y4eeDoxA3VwraPikVFfeE+nrvWlezgDSrM6uttiV+CoOs6WhkGF5q+8TcaApCApzUqt3IBwV
6hq+WBkWDZDGUFlQcnJL/nKOt8U5m5acCdUXfCVl9def2NzRijj/HtZbSMp4yN+j76bEjMfN6m5F
oGvMgwdjEvxzpWQgnKEmgJK/dV0tJJvqB8sx5gF/RcvNzFB7FaTUaXdqgN0Ws+M97AZlahyn1hbv
KzKkMCnzGe3o0ABZ7YhzVjfjT2KO7PK6xBt0vrBdulAmf1L+YfaemDOPX+Zms8DVJrruiQut13Ze
NmVFLhUhY7djbtdOEQbkOE5/fRNxmH+6URERIXxnnFi7GH1326sX/0DExvMY5R02IYfy8RTCq5wa
gM0hG5wSWmrJQ069NsBt6XlRuIAXKH20dEmxxq6UEyeyUN43RQwqmbGXSsqBpbvuOSl0IrhSzE4+
uEmv4FnY+WXjOyedjmprljX64Mu2YZHB0RjcpLQQxvvxuya82tXxL+vAaVhg6UZfXdXFK+Tvyhah
EJ4I5XjW+GXjPc/ROINx3sSdgWx8k2u7iEEYgAKFChcckgugQ6rWdhjXODzSekwBL5Ei3xM9aLeo
35RQmSeBQZC3porASsx4ql+57bN5r41oItLc8ZOgVf2Vf+aaEhRsrSi+xsQJcysv80BZtckvQGJw
YUHVLb8iG42f/b8gzEKFJBHyQ8SIqngic+Bmp0RUODM+5wNQx4Al0mbfKQ5XAWQ72A9FgsA+VR8A
r6QoLUbZi+suINUBdjEz1WgtTEiPs7VFlUtkWmDPg63+JtZnEw8kh0A7hVCnJWqESe8BtCXm1frd
1yc6pqS/O62bIIqQ1IKQ6NISqkzKXI2AiVbbOHyY4uC6/5gi1IKkCXxMbnOtEm5XQ4TpcIsbC7GF
2R81aQbhfdnOo5D51bDEJWJFO1/9x2y2rVr0Y0v9Dnte5/wvGjfemq46s4Ocwkwb8g/zMVXLREtA
DCa2BQY94yjTadzrG9y4UT1M6hQKBNYrs11P1PKWOMKHnbEFGysSgUi3g3E0OfAFrfnsh0uH1LWP
Ky5k8jZwCutCLcSY75RbIK6Zyp1ciGXzGpbEVrXwL8F38HxrXGNQykRChXnie9LlW+S+TFJRxAyp
ZS7P61ZpwqFEx+tqrnxSmhevXv/PCAs3sqh6D1Z5RmyIG7ELwpVnZ03A32bZJFzcCxWJzFGAkWxy
20R2GJvQvFsHcOSgLr5S0Z4vFc/Cjv+gv3wwJCeiG3KyVEDcDXB82ygXJdcaMrVuSOqZChI10lO7
d+poQTSQPJIMF3SERECjVNvybQ5M9WMxsrejJ27gwoUn8BxwPQKp5VGriEP7Jka93bvtoLsYz5uH
CTk8vrQVTOIBgEWrMTIzUUoHxa9/WMbERYAHiKCe+RNHRR+IZvMPVmYFvYGr45pRyr7FyzJu+1wk
VkKHdOZlwBwmJKqf2LkqISXJ+UbZOVQNpbKqkbJJYuXwZfyGQZcyxHVXQmnmWI3wsplEonR7kQqT
CM/j3ta0/xeGClZA6VujQcBTp+4JoSv5nB9S8v4Bn/J2NSsavZmlHqZ9yVO7dLFuWpRMU1G80Nj/
0BWkqzaIOXhFcIQYbh7u6KljNMEaoVFUztZA/2s3S8RvSbrwjFL4yU+oCyC1BnICQvQJMVmYofLg
meYHcHp9LD3twmOnHZqQa36bSMjazeU4y73rRwN8Nw3506nNJafIkJ4nO4HS20B8ExK2DjfDw3B2
Gs7FI84eRc7zuFes4OaaLgzwt6wQKtZUNN1DTxBZNWFFTKV/ZxGOeCjLDAknCSiIJPOdrrHWFdY6
5rp81yxcVNW7nQYrsuHP0ONgGT+ky0QeiOmPKBKXNdwg30z2vw33xjsl/ZY3axXZ7XaNCsDH+w2r
s1dXZ4qLmy3CwE5MpJ2wYHvtFoENwyfKr7m0B1Fu4haUHR2weki4iRrGpLUNdQIO8E9dtzMIjemy
FjTiaFxRwqHcdPMU5Jq/+37IaPBpHmaog2Kf/UmuuQJqJaOuRR8SRMF7cu0kpyHcu7uWP35lcdLp
z/vErLiim4fYc9Md+9ktNdQS6BznWmfIHRHMSgnrIKPmUavsLGQv3tIwe3DP7VzvwqAopzt6L5ZH
Qjy6QHBClPW1T/yx+lbepaGnGQI0p6TYgtFCtLAKNZ7H+rhXIEjvi1sXjqYS8FP4/FzoQrE2U2jP
1m1KYB5R9vEJdxcebzHYjpN6CzUnuWaC2Y/yiyPsv1vPI+fk0gsOItTg5WT40qqR06A0QQAHnsWA
HWo2rzzCxvCcYysLRaq6EgoVgrIgTOy6Dr+8yjcAd3mncIm7A/3Wm1m0NqJZ5QYt5PoaayJpaMDQ
v/hsSaBHzOvtU3ZxxDBXKfIInSKGyZ2s8ERmw+Ko3zeTaL4sor+0YAO9Wj4U6IBxsakXVwYCbPtd
7JwYGxW5+3V6NM9FiRMBUJCD9fgsTukXJwGrDALkrcOLhO2EG0Y8XtNOPBVqvNjfNq/M3GCTBKuJ
9uf//YeRN6YWdIVKK5aL0gk+6LDf4wgT60slY2mbsPdioR5iCG0RBKiRwc32RseqkvA78+veMmOd
C2IIWiQ7osUNVrIXm88TykbpJAcD1G+tRHeHmV+T6i6UZb1yM+KaLhdmi3qfl1mRTvh0k8Q8n3N/
33y9abBgKBDvtEsVakllW5YMkkVHmQ8tsVlnRnm3beMwnOCtmE7L4VvfdEqTNGnFNcYlRH0w4dhn
u8SfYuJtt7ioGeosVXIGu/hnyCF+YC2xtCJXioDuta/m79WhEflag1apQWntcdoYEBBsJsAnvRjJ
l8gAuI8YSj8fxUgVvBVomyqW8vWy+FaFy5B/GQdEcJbhEHJJXPksMvpJFcd9nLYk3ZpyRpP+FRh1
5DLFAocR0fbXH9ygCMZ4S6bm0Y/mhgBIEvNB7fzAQNVQ+3WYmklpenitC07uHp8yk1WVz1v0MDE5
X5JSF9sk+cVeoeU3VqNrDdZifr1XPcs1rPpZ4tDdXOCNmF1dmvZRyK6wJ20DawqckJSlU24OhVVU
3u9sVmlbpeJ2seM+5T8nOuwFLvQMMQnT1F4np3i17PuEf6duWVby1gYO+V0eXaBnBAjAn+00IpS3
jXwMOekQ+h6ZexYLFaRtDAOofiGFvPnDKqMRoMa1oGIhLazw7WatLuB7UXnZLPhAj9SlytNtleIP
JoOrGrW/QI+gKPPAnNF1+ty2ZhhoK5bsQzSUwVxdb0vuyxbQEzW3JaszEN8rv3P1//Ef5FvvH9p8
UlXrkECxL4uYXIfeeYA/3BilB9hSlM9tXflz92XuR48UHOfnC9cerc/o6FiljeeNdNGk9lw6KC+p
LL1NPlTeOAbOHnSr9M5CFpRbwPiJO60dHP/7+ZPM001cmhFUZJuC4Sk6tpX+7q0cexSu3hliwxWi
CiduFKgTdNnzPCWqlgiufnbD9aFRExNR89qkay0uuxBOZUgnpRonlcvNBgv60XzLglHyCycQsQEs
1TGlbNyVeQnRO0W+gW2ZcBvQK23ZYEEIj2DWY/puABxYB4ozn8AlAvo1SfUdZQufwTX/pLXKv3Ra
RXnVh9J5/JoN9BWLHLq6I6cfPwFxMNnweM9uI+D2s55g58uM29inOEqCuX8tcIj9anyWRzzC4X0f
QyDMQ2Qzdml3k/YnPwYJJcBdS+1Oz3TpFQJmJcKLTwZDXTIOj0RA7+tWjNvFgqi22oTtB4JkauPv
c8IxBzfA2/CjmFmWz/KRVBjFnfDU0N4zORA2BOY/lqmB88YR3vFjR/WMGV9bY0b4nEcQb0RaeRKO
6qiXEpOaak/S0vs0Eu48vGCEy3+/XA+OSCAf3AaQtlBjrVoQayM8BYjcf9mdhWmdpLgVNkYXr1r4
6hTpKdB6opaQkbCkc1XAbR3jIAn8YpNBvLO6CzWyuZfsVpvoyO0xb0e88KxqLlc3UGEU+V7j3fAA
4w+NYP7244DShRlwyXmqU1cHcFv54CzKuFtUVcCAWStTVRrENmxDedpwQICCY21/U3JkrGp2wFz/
wL/k5PahrbrlHuwBYMUx2GBhL39CCoBah7Zg5b+dnxREIPGamiYGljX8gEr5OB/zDxIJDy/FsQa9
RqzZ9yAMdiurVieCM0p61/SnBEhgN+7NNRfRDKIVFWpMc30esi9zhy7JdWZIT9YH+PDVK/wv+IE3
kclBNHIOOm2rT4ymIgyvt2EF8aGMvo35YkZPH6vKnpeyULZUo+9RGoVUVNNdum1ywuikq6906ii2
VMOynL1X7e6OqwkHDfaQpMropSrz7Hetl5+GpICgyuYAv0xF7lq20OnF13qOvOIMvNu1Lmy1tVb/
Q3Pj3LuxoQUsMLGYS0PUbCLMLXlSZ1SPL2OqbZjwRAHo2Ps7roZJ3lItMp+Ncg3Y4x0h24Kzjfm3
9MtslNaEtDOmOuGV4MZhzEY1NNrjE1UfriKh9HhuQle/t5T2HOpfe0dyzn/QZFyp8qArE5SYkfir
G0U3gP7OEEL5MA3G5hkB97Cf74CP6P12zAIa14Pi/b6k//fnb6KG5/OfmKdFMk8I6RUqjKQtndBZ
aKoFBnfSR5OkOt+WpAuFBKpodQHEa4hxZOhBoLTSZDPY97Ogd38woz4IvU7Az2Jh6MVq8nFIKfm/
BvKGNSRu/ABWkezLEZ23tScIzjY+aEvuzpBfubqS9CREoeWGzh6F9BKixsdFpaIR2mTABagxTtrJ
ZMn/Wyy6Ozp4YUWmsFeDyz6VbLBByodhA24w3yEs4N2PWkoaZ5hvleHGF4xIBGh/DuLCR3RjJxbY
h23TTmo2s8XwCMvFbYopKVWy25i086Z31bepIjWCI14wQcagYSgmt8P4tY+BBwfV24emsteWg3Qg
mflkUu6P6CZAbgvAEDRXS2+50OSmXfasZIewLJ6FVKXZZAreM4UwkRCxB5NhNqPJWAQSEksayv5h
xCjWOR39REYf1qrUOW8oT9AvnU2aL+f2X5LVrMeQ5ek2iEYLc980uF7T8Jj5glhfkss1mgCEbfmC
+DeDTS/ShPmIGFIVTCzU8oe2BHNk7zfG40kNhHngCwMrrPMTwhHCTbaQ8kRhzIam1NWUnSLm7UdS
sfSYE0YpZQ2giZNDyFUu8IFFOxJ54aeMQu4wYkAclIMblGBvP16lLc2QfDhF64hBFTAPoKlCNU2D
brCzNb7nlmm13m4xK6UQlT6VY9FKvBC3KVNhYZrV5idNEAJ8SjDCXf+Naze+ZqlYklrSIERvOGKq
/ozkExoJC5z7Q7mXfYUnlQXJiG+c+uqptwi0OfhS9g+5SJ4e/FfykWBN+uqVMzTeP3tQrN50Tm2s
249q3o8HDPSdg8mADgb5NgQdkrkp7yxn92jTN1vriscogl3698QQ5Y6gu5X/6um03MbckN3NiOVp
3FD2bx6IEF8dzU71N7w3kj1d8ZRxgxNTevEY2WlQfrbKg2iZdRflecLmFQpzg9PcpOkVo9omGzA4
EJ8qyVR8OA9Z6RHkApg+TMvFtcKy2TmNGVzn0U2rktwoxlkhFaXylMOE5HRtPDujcFDTWdZnCFC+
bpDxy3JIaYuuWCT5fjSrXohXhxGjQQb19SUa2xteXJEEzugmTH14vePn8jIjOhdX92z9iSFENA1f
S+neuF5ASxbbiOLQIm+TeAxwtZ4pFV3RSwetHzUQNR7Ff1miO2nPsgwrZChc7jE7e6A1p19kNu+m
JbYJaurjFa8ON92sVtoePmgD8nkEG5F8375l/ij8dog5/vh1ILPTpbs2e+G0HN7iXm9vm5bIM2t9
WXCePInAGhzxMSy+E2BuOCcMiinV2FmdmaT+ODeFEfZ9Ee/+54u0Q83UK9Ej5yuSnP6nvn2uxTHM
Apwj5adFxRu+CzDZwPtgS8Fzh3mLLhCkssgzOM/bgBAqgkOu4RcXACuud0fD6syPhmGox50Tuh7x
V1zDRqRXvZai5417yRR0n2IiUOvk18pneSn3StzIey230hmbBZWG9/6HahSsLXJS/rUjFxkrwN5U
QyGnYUC/k6js5VjCbRAo3q3UTlpJRH128ozGRUt4wAxkH8agI7uDR14Ko/teyO7AyFzMTnjjRTGd
1EqIIcTLlxKHDpDpS9mWJAAvR046pY5HaXgUobNwLwBEVf3v9h6CR6y2T5jgYNdBK4yZQKITqOLn
p80yfSDMO6J+QeFTqPUK6fHybGSAxYoKmfwMWiSCNoJtyCNm4FvRTaoB/Ve5I1sCw3/BSdV9UOGo
dHn3kHMUzhN5qqFjqBYVtCnVeJlxCXbVSOg93xKs30ushwX/JwvmiaXAmMMIznWpxKnbylyHf2/X
E5nzyABhm7H/PHwm8f0YFhe0yYqlvRtloPyM3FOLGQlh8jTdszkYj1tT7SidnMG1NVsrTd958rjw
TBqTCskLwCvHyeRdv8XaibGLdzL6LPBeaqUIvmobiJv0dtzJC5IN3sic8Qzp86czx7kBDP8d5q4f
0BCPsy8eG2KCkslHx8jSs08PkiO1fx3YWKyTEnz3xMsOcRk5973dDuwehBwy+409tQ5AZjGS1k4u
VW82rIpCaKAjd6X8jjvJCsYhD9mJxhtJJBTBJ/9uBVSFNvlWldMwdUQUn0577mQz41R7rwMqsYHQ
zwIP4A6YfMr3pPFyFiUyS118RwhUEu4YDCgJyziwPRvbQsTFweWPUZ9eOIkLKawfBAjIoOsLE6YG
6C4pPB9+dz0s77Hrx34MaYYAIFof+UQmzn5sGwV9LLjvT+GY98TLKhCMjsieiXsh2T9qnd2jX7hW
uQ1jTE60nlBFiz6biqQUC3pjgzoF65IQJGvfi5hvCQESlQCtDzEBsSmMegyZJM1kGRZPWD7M5QIO
iG6SDQieSrJ8N9pXDNtXg0nv/JWNP4egfaS6JdXy003gWaU4tDRkqbJBusn0I+AielaCzEfvg+Ly
BhCTrSWuFoBCwiYnK6VmMb1QKhU3lBPzX/zFkRDRmQDBCJpDuRBR+LcQrDZmu4fAghDNdZnNJBk2
saazQ9LeI4dcKFu0dLphro9AZDaAqP55ucY+kkLfTiG8UgTEzViHZt+vPEQyu8wlaypHfzcWT2EL
MYV/H6Wax3nckK/LBQcVG/jgtOEo1AChEcWyu/Bn9GD7fif9lMBBGApoSJtJHZniL5Q/pwv3povB
DmfBMfQj641CsbpoLeaBjq4ymATcn1ZirYcjbtbAOMQGY+2LsH5FgE4jhWS+ufB9UhNBLcV29Taq
muGZ7tiBDvvV1onK1iPeShVxsluGFrxATtGuPWG9+80G/XFTV1y7nTD2d6VXsqwb2Ii8DJT0BikC
tw7W4ldMj9aLp4JcaZIMKpmat/UsZa7nB0CemTrbREN1bhzusaXMxWxTfpk2dCVdCZoG2ecjaR8H
XyQwM1d6ini1nOZkqthjaqHo22s9y8LIHqH04JDeafwjMRtJpoaVRoWeVpKcqAQhoj2lltXazw8S
CMmj1VLQdVfRxJjbP7Z2Pfz9wi98jnEgRDY/5ApjuzVOpRvm6RuZ8ayr3LK9KifTdcDEqyGrKh8l
flMeSH1hbBOJcDIc4iQNPTUi1/Qma/9FqWdF5xmIdVSAGt/ud/sbj+GlhJPFgj5yE/DFJljKXDnJ
uN7mQd/SuA5yjSu8VhYjULo1p66znRXZK1TdcmbkBLfIAVtN/yLXw/kROPKftYhKcqaFxoY3In+N
1Kjo3O/BWb20ifqB2wRAdILUiQozzibH6ykSt80reBEYG2ekOoh4AaH9G/uZdI1Jvdg1UpX7eD4w
Q5MDw4HD7qsW7UMcuW6MVXwfSbJuJMeVfClYqcFKFLPt0EOo/PBqhziiCkR7XpbTsRyKITuTxo2N
FED4to6EnWy8JHPOGIZ4a4TKffw7yGwwigfF6o8lkR0DHhDMZVDpbYUC1q7w1491Kfuo3nF1qw4C
vcll4GdK4rKnwIkn3HGLdlBPyrEQCdFMAjlhdpS0iNnD5QD550KfzUr/WMgJjP+uEqiCRYG53ByD
qR8q0lKP+KrpSUpp2HMQNbqUgKIZ6QvDHAcUhzVo2ZTGB/um8Y3Wlj2zbsKTyUL63gifm6tvuyS4
YnvtbWXvzBAJASRRgK547JZWe51/VUpfeTQzlaZg+rVwDWhVibJcCC7cd0LzWiBY9+6r1BkNRZUa
a329/Pfrif5w6HGX3xLHi78nkErySiMJ45QUU4HCfNOsuyrfHyHtiWHWu/0nsWPgniCd8G0IUNJy
WlUWYFYpVTfeqE5nd29XT4g707vA+mROoW7Yekmhjlyxtkej6O5a31U9ZA3XFvOwzgZdLERoHGCY
o7eYg0fQyTV31GsRboqp4Mq2fxBC2tn1vg1CLOOSm7KNo+OOm/aN6/jEfRQJVp775PVC7n9tmkDB
PIc5w+g7+xP29PwlXKxcT23Oi94FU5j0DNRnlvnhtuJ2yIcUISAHMws0axKEboCPCN9EO0oj8BSI
Y2Pt5ME4chpEa5mxk5Z6oGQMjZGHsKZQdaxhfN0WB+2iIEJaxqn4F7HI38IXAc34yWmdos6BXaJb
l9bNH/zuNphYCer+j1GDlRjGgB6o3/qIU0CUnvqXgvUdsI0lX9lL+HENDCmwrFC7mnwVxHSfwphy
G/ROBxhca1Mnr4qtNS6cKfmi1W/IbObzqS3RaEVA4jVAOlJtZGJ7gwpkltiWCUw/tbs5EQILq/Kw
wgp6+pHp+qh59R+bZzIdV6Bu25WO4j/QeBeJ25+Kwhn2QWHKZhPavaflqJa9c8g6kTvgHZVsNJkq
JwBCDdvfwi0Qhn6HXJ7DCjl8viodsRNmWbsG8i+o7vYWEcOAToXQTo3Ao+lvqJlAQUDC/YCDwcWX
ucUGFZHObffITiN+rP6Zn/JfuQYQ2F8zz/7fnDLSfU+9Dg236w+F13Cya1/qFl27s24GTCrpTEGM
dcMFld09RH0xLW2ssVG60zVYReQ7tEXS9W57gOrrnvNmSWVGRnU6zLDEjVQfe0DupPmZjfN9wvzg
l3PlGyXQqj6gzw21R5k2aSyft9iVClYVA8wA6wdNCd/ZXelFF2w4osokS5oQA8m7LOn2+4x9DeFY
dfCMv0XzVDR/2iwMzK/RSvprYp0cO+kEC/Mx/OLcFy72VwO+yWkDhIeBZkH/j+Dwtq1Kg0BCSI6s
3WaCteTLjNuN+i1Jh7SpaNXy5uaVm0uJOxx7DmIRiVBBRc0IDnxUfXPXrs31t8enMan+nkUpHRP+
wsLIKhLX1f1J4C2xH5bW8movszOFQsTuGpIS1og6S86OsoMRVHGLdD7H1mEq+PQYqveQxDaHtiOH
td6UZAHTeDo6qrGnzYfRmJbuJ8Zqi7aZVy8N8nf+Cyew2ag6+x7bmrl8LbJJ/2rSIHbUTskBcTvd
o5JTg0BnlO/y/qEDJU3YmCbp72paMb1ZPm6wUIUnm5vO3AHCqvQaK8oSN1B9mq59g9pBcJSF7mVR
s88yxRCQbmgXBWgwtGBW5/bTH+p8fsEn4jk6QsTUXghd1TNBlzGuGR+OEN/FWFNJoZPFm74Xy9CB
HXr640CMXKo+EeVWs7cWIGbYhPzjG8yO/ntdYiYpkq2+CJHG0pQZnLr7gaI9v1dovbp+gEIl3vrZ
1UOjZMCLJnI6CiaAb+kVf4BzUNe/8UBVpxtmOGJoHU/8+NZrj/SuXhuwCXtwaWDPSnPOhudDvzkx
WgqM05y0UmwCt0OSFs8oKPezPVpW8WqXPu10rO9Z03OZYE4v2QpZ807krkgkTfAgsZelz9vvy/b0
VRE1Y4mFAWQHp5hBvOGlmfplSfgacPpM2cwSDrm3BNjBZIW8kCjtLn5u1L/uKqErhApr6nSd931A
WRyl8DltZN5GwuXa1U2wu+fuLosWSij3QWK0smFovO4ipkrSfQDsUs9XLmgzBKpBY3SwDfUUaX9j
LXJt0fmrh24WxnwzKn0iW0hOhmxVjRA0tS4ZmU29c3sbp3QweyDIinvflEtKY0/Jir8uIX8xhvNj
8SFgHEM6E/xJozsWBBDKer0QQaYVsRWyyjXbJ2NtVjzakBETOlPQw0wzfpioyg20lYURWrLjVi22
2MHKDvRmxzAa3/rAt8kJMjSt+pZafea1wB+GRrNmpdWntCQB0Z9OCsGBKdWi2YL7eF5ujYuyYTVW
Nriimo426X6eZ8Gja8W9lQr9Gsn8HU+g7TWrJN97G12TnoqZ4tTETJXWYAShgDXl0C6I3bmGcLKJ
Y4lTYkKwDUe3UYP30EQptHHGaTnAglYxne5DeCZjrm1/ypBMz1h7d48s7KvxWZTHdRHDVUAb9gGj
djcXu5bAIZecuSRygfVes8JV8D8lLnYoSQvZrugJvRGlWBwZn8SnHSpZAw0vud4pV7tmw+9egllo
RUjxLiBkNw8HzJZShz0To/qX1dL150VjGsDeWv7ZR1YuoFerV2aCtNAbnFzKV7bBMM9Xf5+T9Sl+
/qT3Kd91B/KXiwirl90BbiKQG52GN7ZkozQkU30oPZ6cb3Hh66DQEwUpEzeGM6HL8ktMIs1mBe+k
yHU2HUDA3erHb7cd/OMypvAUMVifT8jWiMQ2KOIxerI1gRqYfvSxhOErk+Wegf1rTXfvnS9GUe24
AV2XtpFliy9Tta0K5d2afT/NIN6b7cBrbrfL9HpHC0qllEqZ3lB5tX15QqqEKUlKo1t77WshUlUP
F5Enqva8MSiyfXKxQivd6ulvymPwH200US6HBuToYqCiktsY3HmKKxSV6nnObDMuivcSlZ/x+qny
5fJU3n1lBsGUj7YuuQE53YmgR3c3MccvBc4DEvdyCdWzyu0hnesZ2Hs7zF0vuN1xC5SlF/ggBMLV
9ksV2UT2bJcuOJ8D3OGh+ypOgXssD+12EzAc8byW2nnCfP7JX5OES2NSiDA0TOMGQbEUoEwLsiJE
965Gz9KETVu95Yc1k4lTjMfHw+FBq8E6NMPTVWN1BbqI/63JuoLE+QpNbDpX6cjMlGc2KaTzQrWr
Ig2tbtsIWGyI0nOBZhpJAtMNKMJf8aZZxglXZTvYkoMh4Zgqok6ASOBX9vASwLh+m2Wwz/wIknfJ
oahxfL/bv0/ZZ8nHBxcybUqh0Jx56p1lOJhk6eU432ukUI4Z2TVaMsIT6I3JXEskKxDxudJdW0E6
zKIGvvIDDqNs62Nfb5Gcr1R4kgJDHTTN8nsZIhM74iR3MmmsfiCH0KXnkaix7Tz3po0nidU4IvVQ
cQMfirva9egjyZIiaMeY/p7MJVWwFCrLk4/mdBNslnMknrym0pjrygAmI+84E8j/W+hcjGXXF5HU
P//o4UQNiedeBm3nL+Fp5ljG6WhBXHuTfvmo0tqEXZLiAZqxR8yOUiPpEEovO/ThVmeyfM18Ayd8
D9kkyYxDtR5OQLTgYj97aI7KdwVrZ8AtIbUyz//ph7qwviixNgaPDZAZEOrJ+GgAKMmXNxUNbzJg
7H7eFP0b1kAvup9zESgWe99FtFvG4qq3it+Etfl3LM5S/4KLZO7ot8AVfHp4umMk5Ov5CwYVRXMH
ozFhLhVyAhQvC1M2qBAapU2ipWCvAd/TyTCcyV0SBwrR9h+lNbGLNyr00a0AoHyB6zx57YhCWDAu
xHH6FRUbx9GsSqujKR/R5FFbpUc+4BTpheLHXAEqtUVK55eT14mo6lnmzmkqUla9LY2afX9rDw4z
GtcYLo6mBItHcC6thhhVOmxQF4xM2ty/YywqbAIoD7nE8A8NVBbAZMI6cTDANS1xA8GlnpTpaVZL
Cu8qq10lVW8kIlFWl9onDfSa46VArSJ2nxcUrLdgxbu8Sj4rHD83ePYn0/7Mvoslbel3ZOb8RzYY
LMPzBL5cLhA+DP9TUlStuPa0zHtQbwsUlc1QvUin8I7xtBMEi3SQwn6nJeI3OzrqFE5Ph2DICtkV
cLF3Q2Juq5DXhwh8gRoeK9Ay+IOGULlNLP88Da4k7orHnJLzxxaLy5PlfieNdcfw+nyWqIq3yKrQ
AZXSDDp0hml3ijhI61GZ20M0+QveCV5TrxC+zGZQXwRL4/75pZa7ExWTr2wUBtOTYyEgNXLnDPLg
2Fs0FACcPddJXYWVfOyhFFYpJNPMpTqDjCUKT8jLtNoOTH1gaPeYE4JKxL1tP31jP6lgKvGVshZE
4f8o2+FY/P+YsimGocai7snfbz6YKQ/Tgf/Mmg8PuHoDu2+3KyHv8oRbAKmuYFYKBsn9Z0SZKedV
V6SCEjrbYxX/X2KEI6EKXXl1C89UgGYrZX7VMUtj2BjuMcYJ2i0oU8F1zFx10nxdBF30L6yM3iZn
PE2dNI2khkcBrCo79VoHsJKXGOoGN5ysyCZrgSeXBVwwvFT2oxC00PKIYRvCnsunIYglzFZCMCn6
Zkx9LZEe1TpQHTvLBJXZsNn/NaCNEopRTX4v2PtPPyOTtO0QMwYu7vLo+75GQFBogDzrAJBSbPBT
TQ4fsAgP8PkJxFeMCdJpBFrlEZkIBAXwNKJw1hf3QX/dZMaQSHE0eHO08PIWRqWp+Qp8CcGQp49J
+Y6IS146/XOCnxP5cpouw8psWPlJ1OH2v7mVgPCrf2ArJjdHS2hFGv+vYgy5eksLwPymS7QKNpqy
v0mF7EhtxuDRyzSgLXTPzaLonHV9SzYCKi11e0X3RBcFXWDLA7WoHSFwcMg2lm0UZZ9zBvHk4RCP
fH7lQtdGjA/rf5ye0+95FPVoRu16UQDpxFLSpTk4SGeIUuTW1Ets5P52DkmtAETjOlUvATCRVlQG
9f8x6IslMTr2Gahpypiw2QN8Ufq0tPZx4sSv37FRHe+WQhnvy+elzfucRFQS6k/kH3H8YFCdfsvR
+oqYBzXxk/VfmlLdJw531nB0J74eiyUpoe1ai4ePouZhWvh6/TgMuwmrIuxctrDNQPlwi0Yw0pw2
M4WZ4/JNuoy5WOP8pGSe8k0sKbO6XZel5sEx71U6vW49DgARk/W0bFWkVENpX0EOANxbese1U9rT
a35gY6nZwnwv6ll/Y62KfRSn26fc7tPLlNJ/MWBZNgHNAD+Yhea36c1F8K6O/q4+kJHQG9/dme6y
od6tZZVNM36VbFh3Z0ae90YZvW7lgC9AUSoDP9fp+XaFo3WIQnA9jaiC88rpEF6QzoZZYPgqP80N
1Al2t8CBLEuOYfErrAeOxVOksOYzPldJd1qE/cW2F8LbQ0bcqET4RR/lEWPPtNH248PabkJn3ojK
LVRQwvQhOK1WYTQ1xwt+Z7L8GCUoSk4bMPQv56g54TaONy8R2rIyqcYyKjF1abRSz5kKTDdVbdRg
uRxJ8yRzFRSuE5jspoykL8OB2k79Fp1mcZ+mltlJm+XZpiFL6GO9FzZOGKffsS8GQUQo6I2Q7c9n
VaWB1mWcfL/PDDvXQHL4Y25Tky5gdGgTAOeETo2tJEy6xSxS527A0/8FeAmY6XFLiTEdkuhVzP7w
UWgnaI2z5wgSy5y8Vx2g4AlHGOiZ44Yx4kH8hiRxgmTdnC4E3AL7+hekghMvb8TLaARkqTtF+pQh
zY307GRHvf001JkHRIE8oGWKVMUhJpXeBC9dGQmipADBPbSjQ1Y3PvqE+aPlr2GVpDTxzoRZmUW+
dLFOU5JNh7OA/1TyGzIooeP1JyiqSeM53hwSUMtiDwaVA7u+yQ9bG+YkeYRD3LFPxmbRpoOheQOs
ZcMXbmxEJHXaNennR5MYyhyI8y1JLv2g+4PVdbhgd8aI78zJDI3peXP0ThyfF+1oR3Da6/Qiku7h
/ODVMZzXZpucSuxfyyrDd/8T188M44F4tV85W2L3vptMs4RrWVXQoqb8sFDYu80V4tYS/zMWf8aM
bGDAy9wP2U8P7eeQVfyPNqgomxLp+792qDbPFHm/jUpp7I2P865bmdVr/p8kM57Ly5kwQ+7RLtt+
SzxDlrdBZD5dWp8LI/cxzGNVCHznjMDT+iuwT5Dmr92NB9Ouk5A/AR7pEk+uGwt9qt4N9uJvgyum
D3mnHWPq1RBEvLFdstdr56iewGgDU67ayWQhW2WFhf5/Gk1CL5xr0gj43ufU9GZ3aDH1YDhqGIQn
za8/AXuHWVaCPOf3z/XCcdHq8sbEb8oDGeKasmn0mDcsygtEoMxhTAFkKBW+StrZ2wao0MuFziaI
sQuQ7DKlRmPgukw9k7vi8RgJkxAIh0mtkZiCSPS/SDjo2qg3+5tuhYgonlJEPoO7a8FQWcDF6AUt
M18Bfi9KEboYu5JvXuekdrIArgTGaCdlLA1Ed+F80XPe0vwRkSKlGIZptuPDjjDiufZe7V5aon7A
1ijATOQWwsOyiSP1W+8MXxl5eUBKzKXWXXxuzqVNz9sB/DxP2FvZnCU7trQkaIBsgOqiD5wtdjdT
OI7cvWjKlWYEyEQ1/3LKFXjOk5Q4lWKpv60sP1SasgFj1DwZ+h+/eS6IRaeB4un7BjfemvCYauMu
OhZtMsgydGnUjplo31+Vu9a4r6oQzPfu8syA4hGGIG0oj0MeLmL6mBLlSVMql+DMBJ79R+7nJiMC
sWUXBy9s3wLw4fGOhvs/h0161Rmu3ZLAM4spPVIokt8XjqJmBu2DUiLpcwR1DBYdL9fMSLyMEH/4
4JAw2OobEvJ7yRI1w0eGi8nWsU9cf81fjdQAuhAaZ7K2SlN78/7pl2zwfSCJTHqC+UyjKRKSnppr
g0QUqklVh7f+I+jSX1Ty4pCs05wi410oX50heRrrAavacu7b5oaQtqMLN6K1T5wT88AHvhsUcJ5n
5Fmd/ofQViUWksnbDu8nPn1y1N9GOkEOpobnz7SUU6XGWw9+9alvh7MWVfjhFaVObaQvD0XNON/m
GSGAPN74uI+OJMPeA9NyjRi22PK7a01eHqbrgZ2oyaIzAysVt6QLrFyIvnTrX/Qr9fr1M556uPg7
nNzyclVBDQilBYO3FF6rdvxJnLYSv6DNCEMMYNqPFOJgsnCpCH9jjkP21LC/d5R80b3+3tHedi5E
mh+yokg8UkF+L2g7aayelFUQRYhME8ZrlmfDgcfCPfw3o5Oy0Z6krqZj3rOw4W5nM/16Ep3VH2Tp
bhz7jGz8ijJYlbf72kVPMb/XQuKxLGouOh0v+A0ewvQjQjgxlMVFKiRk+vcF6PtA5sWIGwu09d+g
0/uylhgg81c3bAIds98jcJUVh9zUC3dlzbFEmKRIVuMU8bbyGs4Wz0kk4kIVqLAhgxVGjTaMU2VO
TiktOcMhPC8skQuZ20s399RKKTaTri9EVwJbVAkd9oq5XUdRdYLVrYj5sOp+bSyzIOrUXnVOlfWe
WcIedsBk5zj1u8nnFdjckKaPWHy/ekWR+Raj4IcyX/QrTdGKZPd24Lpe5U5NgHkVCmwk2xw0HBBL
Js8u0fgqK5LptdBMKw+pXvVsnM6xl9sJ8QpDOIC2FoNulh5vG5dhxfH2EC2M/tbdsN4jtOREY7JX
IrEpTsyPixrFeX0fRE9owmvP0RJbhZnbFCLaN0Zh/crKQijfEeEngRTQQnTzAcxQVSgdEFRXBsU9
4sa5TRHPvO10b4jh8O5LYQlPizQssGjOU4bdzCZcI7dMycdnDKCQwSaUj7FWwN0qBhalTOrII62j
UryhiZJN4b3F6lfshmtRSYTwOp3go5zKTzI9WZRZVwuP1feqZSCnhxJlrAEDI7QAl3lEdtrf7qLX
E8P6pWCjEc33JCogbEM2SiC79lj0eNP8y6V0kLyAYoiLj1GuXw0NoSKZjosd+5liD+z0YbvL/VoT
IG636zrj6qf74tfJPa0+bTk/Zq25ye0qlw5zIWBdQR7nRjJ6KrfYZQ2ipuep8eQJqzXE9gccuMqd
s2ayd9bBrDqayvy0SEEIzQTKPY8vknkZ49x82YmN3p/2oghGyaDqgtxXVtBOUtRLDWjvEQ15RPpH
9SvOL1sGDg/OdUm4Kjqb91LtQ8GFX1prZwyCgGg9N4ksZMag3wj7VndgDAgZegrvOUYf7ihLkCi7
9bs1wiHgeIoU3OsQu8PuoLBkAxgS5ZJp68K6WvYBTLl7xHOMPHJVCtGqz5zqCAHB2Vp3f/dmWqkt
fo6H6l1GRJiZShAVXktz5u4QYRd12Py71H4cDWDPJvXH4EX+sFydSMpvLKAiN/fkjrjXZWpYDiWK
xHVti5D1ao/gLb6xoPpl2uNa11Ee7NEVx06LZTjFzf4a6op/8shUWVy5mYt8epe5NUJgtsQEmAJX
WzZIZYpCDQtWuZ6g9mpk4FxFhHjP+S58WYW07SFgD1A9jQS0fAc9FUZukgP80CMv89lJ5f3bEWvc
ClaLekeYEF7uGWOd7jY7xh75XojBMI7RVkChgNyBDTsh7hRgkcvzMTftYlYDgigHTVoZsL0aNTrn
Sruh6Orv77YDJLolO9F12FMsVflV2F6VEph8zVKf4d1Mo0QOjZHx6+9NeK9azeZ37Pi45WZgspN4
18Aq7Q03U2iZEUCmvyR3K4lM21r+5xTnmG+mWiC+Ex0RyYb17DVrcHURFi95cKCaLlKFinlV98e/
83eDnYtqShcpmgTZOAWcWBVC+utyfOBlgphjuZl0XchF6ibRfOvmD0enFE+5Y4TcRA3ME48DEP84
dSnaWahfYLnivPYFGb5j4b5MbrgtL3U8lPetuVocB9yxphEiA48uGuYU8EIhuJufnQfWGCp+Q8Ok
4j4YKjftYLF1KHwDtUZj6lYa6HOvl784pmY9XHA5Urf0fJ28dRsNkvPW44t0qDieF3ak4jG3b6YL
War8qFVDZVTM5dJszfzcGqGMoVyoCCiRs/WodXqBjPpaTVi/qykyTv5el88Qi3IL1FD8k5a7RJHr
3u9QLI+mD6UjcLMy79Nl6q7S+r6Fj0MPFL+Egiug9nChJiBUHxVR6IHsyCACBS/q09spAdkeZlZZ
CefaB6Kt7624nkqVO5tENeV6b39BksdDUTJKM/GR00VqO+6Neo4BxQwb+/qLZKGYZ2Aww/6foDq5
z1Erempx53BLZ6L3bv+ZO6Xvo16JkJHIOcNTBzSK7ym541W9h9PhBIKuDGYybUXsAAKRUGGhx32s
Z4jkFdDBQ/4EGGmwJ7RXmqNQlG8N9GKeU8ivWrfmr4vOGFjoxJ4dz4Sw7UHESbYJw9t/kx+pZBl9
gp0z207Bg5f2i6EndHKIM7lr5G8KC1wQrvE6IDjOVKasEmlEgsht+tdWspMvMNA46NsI3uikPx/g
JCtsznFHJz5RThrEGB6os7BrsdRLvjy64F1igUca1pqSwVQwhLlC9MBM7WqcyFs0eYfp9MrBHEVx
ah5auWGVqoefh2ERcYBfSQZGWNwPcJEo7/8zvmVJF6QogB2Hwgi8vS8NVP/36i1JnPIvNpU0/jxi
0O11R3nMAw83X9k72OHkMVkUD2JqSbxB1n9HqFuyxIB+x/3xcJSOPpni/7S5QPu2YI5YwWWt0GbA
TZcBjX6r/hB3V0gGJ2odz+HTZ/RhfFj2XP5otu7kq9dh6ZkzB+t/74WCoUcunu+PMSC+0WkEij19
7sZb1/U3uPcePuBLdx4BIJNnc3CKCbH2DpXYSATKgqqTuDUO3JCNjEuCbTbOHmI77Y0NqaxMtUZ+
gep7KgrHecK1fecCHo3q/djidbR5EuJ9NwbPAJdndg6GGEvQabAp2UXZxFRaPmYUomHOVnEJL7hc
7o1KON1Sujz0GqLiz6KFij25qp1L1NNBfsdF3AXjCEupW3JJ/O9oqyJAPPY3wOb6ffdurlua+77q
CGsRFVZxbq4AmUntyRcs//V7Pzya8SczsWfqNE+RkB5iEvtj4zEDPRaXzOgwVaoO+pgclpxvgupI
CZ8AVl/d99y8KUAlPM9c76y0LBVGySAgaj3m52mwG8jg/k3B08VCi19aUg5pfUM45DXsimAf/poj
2zOwb4BBkITInulUxNWEcM08Q92TjmBYsnOeW307wKl0qCKMoKJjDGfZC/5Gnogl30MTIMkDXo1E
FCw3J78uV0oS7Ao+x0PkweG+8Dw6Y9FIte/tmnopl2p4eeYH2iVnV7qbc9sVzBxuXwFxcMBoB15b
tI6Oxm1/yktY25DoVOO1SVXoDXYtOVt14NbtQuXLyBBPPEfpC+ajrQtkv4B5NY5lu8KQaaYD5732
Ev57KrIcdrGUG2xNDIEphxnNecDnxPY06WWq1GDnMKMHwUQg0LEi39DOodW7iMfzPtOXB+XIOSoO
AHIsaiY2HvIRE8DAu0FiBG5tp5BBDoJIr2QLv67eXQbfPDNXF+IIDqM+5kI5XKUJXypjCoGsMTkK
TGCFlSyHkbnZxrCjP1Rjhr6UyQqhGr2FDnlpYANmFeuSi3dRvs/v+f1jeD4kEb5+H3WXfxWASTUc
YYTtOL7ZSUFHAV50EiPxndd7mZOIaaQzpqg+2VBWHQmFFEjQTyyul1zNIpc0kU2ByAbObKXlBHlX
JwLiZz1p4kG1Y379xCKYH+hJfyyter/XlSZ9Wnr/YRV177lmGarkIzNhjXKe+GMszGGhiq+uzN5n
16v9nKG/SY8gKHIxAjQZNPVAi7gByVh9qOAK8em0QVzTtE7M6rnLzKw+C1S9SLZxKPV9Tu3+aI/B
QAKeFfYeVPrZ1vUz5JrFqjmSYkAWmSrJPF1d7yZNl+LJo/DiDD/lFASIkBaubvU6oDl2xJ+APll4
gyTV+tpWZd5rGxuUkWOMBTOFfSPXhKo8SU593SoPVxYPiwel099JDBQgjiQolJsHUXbJN3Fxbq/Y
1HJpHlidIKyQComYHq27rOldtK9oOG/gwGIaL+S56aqlVrE8VKycZBmmSHbNx1adlUooD1mHzfEq
s++ZvNPy9Vk96MANNjqBmDAJ1VO4SsrFF7uoS0T54z2jNtkMiYW0ErMVbUFgCVKub4E1IKSBym40
X5EtdSZMgkq3rPgV+0geozW+iSQG7a2oLsY/NUYkfrzVPXHVfqKu5kdCRrrJiAnuMAk2OBEXXL3N
Co2uJ2Hsz+9w6K0SXR1/NcJYMfyZJAzDi0QwgXF51YpSnKj8ladvyHfhq7bck/gynJw5C8K2LEJl
U5qCH2rFP2vgGkLfqP+fgpsKD/hG9KGKLemKnbKIzNQS7FTkAS8bzkLj2VQyhSqrS0veFDkRM8vH
bpkbb/ZeSlzFxBJ/mgVKVsjsaaStKWDfs8prhZG8NeC6u3WxB0J3urMoAvQDd1742HdcZ5y4GHcv
J/Te6wX4EQMHddQJ74EKEeGFJnNSgpEDPO6b/Ppb3Fl4mCVKcStLPJcuC0Z0294Qv1FNpNg1zrVI
asghQ2H+cH2NOJeIxlPjjPbra/FUUpGYpga4IG8FzaqsNnPRxyVvQ1ngkYXRSydTZ6PY04ZYodfA
6TxeQtkosR0jnSDnJNkb7/JBj1+qVAOFVwqnq7y0vAgI4VOfGwSNMlJq+M8HjadwMxfK3ScDMDWm
CMBTNiQ/5uj5/y83/+z28cCFQUMUVrPRavFv+GZLK5EZBsu4vo9UxmqvemEF7l7oABtpjaSvzWOy
xx+Mn27Tm5QU16TsX4s7KH/sfRYwD2jKx+UskDT4kdoQXNaDAjQ1zOf7ZDWtk3mzwaAB+boeKwJm
ifpkztkg6CIOnyJpmZC6q0Oxl1K4lMKYUdo5tjKn/tYSaxPDHB14KUCS9sb7mxbFyHFhOcbHvh6T
82Gp6plRwqWXKC0HZIi+lNNS+k6QMvx8/tvj1WbDxfHw7eIGSp+8CU64n4N71G26hB4zVAfHga1o
Z4RLh4EP6uJO3pFtRA62epqCNH4lEINMMx8xrMd2Xbz0PIr3ik5A628c9X2zibww6UnkwzlIbkMU
wgRNsR3uISGE/yMDFJAAHq8fGeNIhRmm/otSTIwY12MMrSz/anEm8L8hfZJ5xBewB/G+1L+anJ9n
O0XAKMk6mwYHyZdv/xHBCZ714BqkQdStlKnOpP8Mp2xoHugO7MwEedfliPMynVnEvt7H2bDe80H7
IcoM9M2wBPecvHDJb5CITYyM7tZ7baQXdOiKZelLPXxhO1O9symeHNL1AuQS8UNiC+hhXwxfoxtz
tMgwCaohDgnUHhLUlKWcp21j20J6H90ww7SwOUCD3Orb9725fqoLNSez37cFsn3/nE2g7e1zn/eU
u7PvupvyPkKEprxUOuKt4njpRt5aSLjj8wFdMJ8nPXoGppW4i1KRUBq5mfRgWwar5lsSRKv8KGvp
HMnRyjwp0myZObTqhvosWk1DOfKUiJRoxPEZ1De8413MAn1aJcitOsZJbqwRtVIo7XWe9LNra98W
/RUNizybEVYzBgeLV60fLki6hrPnmd64tx0mFlP5N7iooGBQTohiPK7yB0MC5T8MZsXBAaCw5Lcx
n3wkWNsnGWjysEaJO6USBlivGLK6+untn6l516201tHP9WKDkg+Os7HapY4hYw+aXIWDEQTIQzO/
bU3KpojvuA6ETXno7S+Lrkr/Pt6x4kSPnDLKmpsudeMF5VJrgB/PEf87RoqEwhc4FkvPvp5ypfD5
2Ud0d8B0dlV9LWcGz95c/FtanjgjqKsGKIj2/D03X3MP0kUAgio9kFRdhWY+wIX7JUxIhTFqxgrV
N2Xzj4boZHIU1PPmjh6YosTseqyORVwQpoeeUr+3WM9+uNvVse4wzFJ1s9jWBSg0vYs7qI2eEMdB
XL5ycy2m1qlMvz5NATEpePNQK56zVF3YQP0ggTLftH9E48d9nShsI05ubFP33lKrWqjZw+ukXQ3c
Rzccg5ZqJ6dwRpOgb+Zejw16DAux7+9UeBvrvIdgL0PFhzoyyH0AYsnDUmG1rYxb8SeFmTnS5Lns
/tjzb+IoX0hqH6EJSblEEswBFGdFiFepECN5s0+wUqbL8k4otMi8oyCS7Z5YhIqDtfT340FV6BMd
duh+rPz1qiaKzPOn6Dm3A0Gydt6e7/zMitrseRSdWXjnVy0dBJxX4sLCF6lEWCOaL+ykz6+aitSP
T5RfezquCae1ShJ0otiJ1PpAYxexym2Tctq50DcjTQyXndv6PkU8F5SWxATNa12iZ15fp77WRpMZ
8ZFH4Nm18UvO0vmh+ioqT10IZ9q0rQsz1m5Dc7SWGWphEUzReIJWbonx/41NNYBeQdIEh5KB7guX
dqwSk2+gSoYv1zPO0a0LD9b/wbctpryNzQ2FRlEYiYb/g3knfYPjdO85ogaiBJsKGuoDVyyoYV6e
U/m8djOsyPWwPUf3IP19SfR7leGOMvomoXW0hrMH0zWcyADhbowHzQQf8Z4KDonW3JIChfnOB7+x
R5Ir43QfNH5pIqmnfKDGvgdFbxDcHvB8ETwKzoX7LijD66/IR+0YfeHaUxozBDUJzIg/8yzYgpG5
ry8UTApI3idcdxRFaloa0ExobvtuzI5IIhPtu+MvH4pwWuuUOzbrGN7rZ9cq9N/RCyRKd02G2Zbn
abyHBXtmieBE7McNlnCXZG6tHs7Ug3GSfayzAID9mMXUEICmPU9VPDsVFY5GgKptYWSuzVRfEjmC
hgnwipBoNLgYNmdcuQ9OHU4ZbylFPSP5tkUugEt+Ml7gmJV0z68/Yl1Zm37Pp2qxu6AvXYVRF/3u
OMMp2TOdvDJ76REfN5W0rezEeOaEaRfZigfNzHNCmi1A5sfkQFF5BJW4zSEs5BHR6V/oR6QaE2Mf
SgkVnD0ZGfBzMVdvt/+gWq1MaJ/nkHPyeDlpjXa66YSLGYI7z5N5BGNxmCeXb5zeDUsOWD/Xgdoq
Od8i7g0m7xtbr53Rru2PVhp7wMROyVaRNrdINL2YD5o3InZ+KyJfPgAxCIZCeeYGKgc8Y6htC2ro
qMD5te7qJKOT+D0lDFp2rgeug+BTY+ZF7E5Dbil+ZB1hkl8AGEB7xiUT9wa25sU8ASlF0WjbOwys
+lpkdckmrILs+mz4syWxuapZ0o/eyNA5wINHWsvOL5sAF+iHnn9ChHmwNQW+xGqX5syzQLYZoZ2T
PcRbTeYsdGhL3aiMFQ9BLAHqkfaM+nhV+vhjche0Us9FzrRf8ZcFJ6yXxT3sXtQCTtWchTWeoqLJ
mpvKD0NzxNf2Hswz+Qwx20Gx+w/LXeHD/fklZSNcd7ljYXhVCB+q8BBHlH88+hoULNlXI5LuhvmN
SdIQLIiYedIs9R9exD/3Brt69++38tlgm9VIQBTDtXIQfie3LxLkH2fdHwwtjviPXDz6K63rLpuE
CQD+Jl1oIzeBNs9dIali9lX+x8g+UgjbkLHi9VvdTBhevpK9usLrEmA0gOYTSzW5EiIxluoJSO9A
E0E236xYK+Upf62GGwibDf+EAjW3uDFHfSw3jjW1USV3meIxZhzMorjvbdi/FrWxLF01LE3XCnWj
bJX/clGs+3ECNWBm+2kblv7nP69I5H6TtS7Lc5lGbVYBLNmGIrpSrGA/FQx0vWz+YeYL1vlYG9Zm
/8xLUYl6oJbHjAlH7VrnK1L0AyGDqA82ZPpQkGuatlEVJ3K8jB97G+T8jrgU0DEH2DWMXCP/AgY+
Lszv5gnxa1sd3mKwt0IDFsuv0eaeIXBhjVqJ4i6LQ4vM47YKYWTc3+WLNZSeV3ECIRz9BLh61lsv
n8kUhV6mP84G4x0RluYJ6iNkhQf1ID4CeV2cAOT3SM+aIxJzOH1ySVI1ecFVHK4E9F7Oagi69dll
2qQoFDkqgQC8+lrcCw9JwvFh2Wg5KddQwAF63TveQWNV7B3pViFnBKYPEmtxJ8mPkMC6G1PDeZ89
QagnWed/6af59bV1XAgz00k0g2Q8FqVZ743tlPzDgXCGiOJYeQWmpEXwIkJOS/4DpT4TqZrqHwD2
kFdoiYlpHAJ0xr4AiAP74KCrkhhOyZ7rDWNhcbreefuWAPVnttQqKTUznqaxK+gb1iGRaHKI0osk
li2idfmXSC+72d0ldqaL3/mn0eQpBXzyub+Bqoe1nVMHLrjCZVJpmYMo6GhBwNLyNeJBl1ZCCzKL
JLVvotaMwxe/sUv0DiV/5JmHoXBsBj/OWGfOrfUh0XJaon0W1GtPQFO4oS+EJsC8Uhu2dmeCkN/x
byIFo1CkAM9DtLuZHH/eEbheyEmWvwGdaC/yqSZy3YnM7gxa7ts/2+vlL3k/lnNMBfnH9YF1YL8M
g1A4DU55WTxyVc+KHpScEf3PoJZAGi/uVbFZGN2349Hc3kOygzuy98Ya65rKp2BxjV9lzSAAwKsL
dnJf9I7z3bwD2akMdO3Y8g01wQK9ZQERRLsxgKqFzms+wR3FIWGxX2YHOuuyqew8KvkgSYSnvwVl
JTxoQ8OHpj94PCe3L+0JOwKz5Sxbj7U8/BLRVvnQ53tLGRtl1iLuz9K49Ohxq06Q6S0vlw+swalv
xR4Aojfpm2U2IqTa+XxtG0d6NOiGUje0c9i1Dc03XX3qd4B3h5tbpSic9jMRUnndam2ZdBOTUdZh
wHC1HQi+/VvBIibCzeoBVFXHgZs2+CO6TLfXOQ4yoIypOntWA93XLePvCwEdrd3jSPpjnD9cUOsW
7FUqVATCZtxBPEFFGvJsqa2+umt/NXMsQRG68E+U8ctqz+SfRSwhBQOMS6FnZLY1LjSiMyiH1XB6
tbmfjPfih3wHIGaqWNFGSZAA2gdn26XWADxlB/oAeaFOaj2sbjs4AN7ig/i1ObT5I7GbP8tsNeha
l99JpHTL1AHqFloK6pVY6krNku/wCfxJz4lPKisWOxbzuSv9v57RvPaZVFUhjMBqXNZBGRCQvldw
/ILKqhHm+sMU0VPXK5yPuQhwjoz1W4yR6alXcDe+17GWaNhXBRy6Rn5IDq/djjxTPznOybU5ITHK
QFBaQy58WAZk1WoOtf5zNRONurNgY/BBeMcSfNI/5s4xpoUGZ3coDc3k48FSYnuN+r4KGYR4LvPG
XGXlFKT3obYsYs4JQHfLA2fFF+txi2Zc85LEbX2tUqHH6c5mLtonJoeYEyrWP7IIVmfuBr7OUsDm
NbpLTTbZsIOIpWjm42J0Yv4IS8wV95rDsM9RAi596O1Vx5qLBzEkKRkrKqFRWOk6do9GVrdXvBZB
x2ddcpImobr8WZ4sws4W93VdqykQLUH6tmjJM1J6G5tqxZEgxfgp1YWtXAcIDojPlGJLLbd966Ed
4qDwRAZcKcdohEK0TrCaIwIVrYZYe6tqipA3vmUl6KzSIW/bppQgAVZbSaBlHyqqxotCfGUA1Juc
FHb2lxSroJwsWLpbBmOtLTgK6bLJkD04vHpBdGeORKaQrs/XaQ0dVw5CbaLn3SpzyACEY1PPVG2s
GCmMM3GmZiwfQP9WX8CLYh5HusD+X0vtldsjaVgXZWGbj/KZB+RSNZlDJ5DMTSk5x3MWjnVE5lxT
MPDENClQkFjFR0obION+yMgQdbNGXzgJSmKM5gf1P2USvED7p+ALV/tLexLr7I35iZPD9fvvWqWI
KbmvGIYTeY1sRhLzQ07ep1JY+R4AkXF7yNKJFwopdMPglc0rVc1gw25Eo15XZmk8mJq/Qn6fpNCj
4dYtyEF4w/a3J9x6MGpMaGgDl87aapEFe1U14Sso+/+ZWxxftO9GBmFh+FNzg7GT5yASVpEwp+vE
cH7KPLyxzqxzB6X3AxMF0hCyO+4hNhqYWpYbbQK89SDMR7fgAMRWjXExUt5DQ5Hq8IlINa4bW7Tu
u7j2YRoJRar05PVbAEus18Mg0WMJUFsfqH2mjnjJyBdMafHVCTnPrdeBiJNCi7byc3tIuFdIq+D7
gmudaTyubV4w2fSajHBjEIdTmdV+N2NTUK75lioki61rfkPC0EDUDFM+8SDasQ8ENVCiMbSd0yPX
6tkCLQciVeV+hKSShsT2KREp+lw19cy/HwAs9oF+HAKEUpGiUJETPBVvpz7IK6YqlAsK4zd0TmW1
bTfssSjCgJ3Dwqr31NrrhJUuzr7GRs9YuDLSd+Z1CH8sD2YlB9IIPRQApBHczhefoKLHcqvK4U00
IMR0WidrygfwWUE2464OHIQns+j6+ki+mdoSXzkTMbu3UkKSCE7IpBMAF3h04Y31tmqCqUkkxzwS
9JZG2ula14JV1oyn4C0hztTq5F3cEyn7sMNrwntE7Y0sgGKE28Nn1Pu+plYw26r1tZNHm+BkOgap
XkJ/ZyJbOxtiOfQEsg46os0euMzUNVlcj6jtZB2AmmKpqBJf7hOq2ZHw8AMOqPgcUTQrkRJr5+Ip
5EWYwFfNY6HAFIV6A/6tPfK8w2Bu1hA+dzMYhOfZQrEQgBBX20GM7exnVqn9RPYny/SpPK+LaUbD
TwLq4RCsPmE3DvzZaZsMQ7e4G6oz9+tAtz+QnTma9+RbfnSU1Cn46Ok3bpF8QABBJHmFWs/CRqJp
6L9VnHRY/rtfS1lKs8iNGs8HGUbPZYBzLO086WWy5K6VUYbbyDI3obLKKGm1clGoF5+CJGLjeO+t
olhguano3lI1gAWkzgEK13YtIAWylxq/MQBqPATTBMyzYQn3A9ilFL/cGAw2I0+m1WQzErukGOzY
Kn1ZOGYzQv2K4pTmxjcIkxewQg75IiWI75Z881vgNy9oNmqz953vbEjB1b5oMQTIukbHDn+xqHwa
sWgvWYUEgQOx9f72VprCXuraTeeXr1FPjc5fOgtP6dvnbRiN4P4PzJ6Jc2YUhyZ6yebgqLsaoKax
QPcU0RppIC/xKQqnlH5goxOemZVh45U+XDYzte8wCxGNDKlgO9+0h8l9VDyXZEaieq2Uov5wyERi
M9jzpscY6/EreVOoCZ2Ai5/wNaVmynMxHjNcjGbtS2qTh+h/8X8AgOMJiCGvWIAXKEKHZNsIFQh6
r/eRSZk8YlkChNjVAdsk1ej+hw640UYGGjApjknNljusMMIHkc1VCKP81rP/o6cuds3qauzl03Jy
ThVCJFDuSGJ/dvsHd8USsV3bjQnGuCXBUEnPKguoYQ6LrteBr3zOt15elOpE88q4OeajoGV+x9XO
Jp/OhguKdJJyFFe8Civ2NK25mAujjNH5bxnCV5VhPGwRGrV6JsO1R2mps8/S6zwDzizH81ugkjQ3
beA7gc2XIXpyLkTsTFLtYWC1y/mUwmmxc9e9jcLi/w+1Sh/0TLtry5pqmjQouZdYN8eAs2a5dM/e
vfvY0Jus+/jmF1gWEx5Kx2MdHWhGTDdp/oF7yK6PhHmOxtHtel1IvLj9H1kSbkdqHINRfEj2SdIS
BvLwGhTN6Tw8AW15jlOXQm8mUqzRZFR7q30QzO17GF0qA+7cOTW55iitftcmpbbLmWrXjxYXHLIv
SZjTyTs13dEgdGmilXEHLbGmK5Tlq8MRKCuav0Af4OJ5NqhbioFE/0oG0k+uq56UUZGBn04OsxLo
wgGFiEtExJzNt/LpjFyQ67wmNKOXHIeF3SemZnpIDcjW84NayznUtD+PZ6qBiIpO1OECaSF01Pxh
CMv1kHdSIGjqJH7TABCrsyeRUA4u5H52McunFa69DeyhtIBH7dyHhngnfUOR9HShcndFKGaBys6p
7KuNiOaARMsZHe1ZVfYZEVkDvcjGoXji9qhIWL/FWfHgFZrmoS2n4+Rbnn27RWujxf3M4DOV9z9O
NeoBsw7JK+s4Dzf1c+fWQrJF+YPByY0qZ9oTHxt9OtBA0lXYrNSDSJxolwK8/zXbEB/4fPweXbt5
rfWD8HIU2fa3ku2tGsApNrTCkr+1tYf11nsMP8l1w5d+QmwzS1tme6O0TC3AqNlMbahNkX54Va0S
qIQSR4tYpvJNzs7Rzr+8uoN8KysB9XIO550u5AMQUYqeKJLduGnDZXymeWV+sFvRzITnPQs8/AY/
oyyWZNHf0/dyo0i/G1gKunymmhAw9dTaNPIzL0JrBbNm2iuuXUCTNmERTR4RhGNNnE9nfiFZkVGE
45l4CfIhfRLNy7JmW0ZL3TwtuywA6WWWXKLHN1lZZVuRR8DIvOIuf1oknjs6B3/MlMOEFIWPp0qK
CL8B9HyLnzIgfRhl9ClOftf3atVsCYc7lpQ29HPwUrgnMGyZ74gP9q8IQyqinnma0Stv+qXdlb1C
tCzesfo11hSEc0A4x5kC/COj4g2R7Jm/P+jbYe9CXHh4X6Fs+t2rHLQvbR1VKO0L+dPpSNWTXPGX
NITxzGYGgyZL+C+bTeTfqGAolVz1cjFDPxVKIDqgquCfog6NqsXFGLDe3R46NqMFY9benW3D5F1J
fdzwA47A+7oqsNEZrsgNyi4mmDA5s5yOIu48andSGpAKEcUiz5pCPfZhY5gkYDhoVdEgCuFTjXef
EQNWw9I1H7+bwtG1CSGK6Fs5PXpDPxCZhNrmAmq5CMGgydxii/5ba3C5VQ5in+KNTuOsX8WqivXy
EnNNu4L4BhgQtMDK7cYBaKf2Q6wjKvPns9263w8NcX5QruuLo5/sR7+cNtujxGA78xUWUcGfUr/k
EFY1l1Mw6/gAYJ0IFzi72INut/SNuI0LnfDDt3FCQhLr3r65+rrgObYHi8YO243g9e5xzlnXDzWQ
dnOeqq/7CkpYwrYI/Wq0+NYrn8yB2VpVGRMw5pvuocL1iKFfMkYM064G+r08g2tL/T8Gm1GM7aQk
+uLZEEmv2fBwyzFH3MWADtBkZloEx/kNrJbD/MmlOaBNxHdCXTSQqNmDDzJrWBG7KP0b+t4AxA7d
3OE+Wz9T7VyJPghcd+NKJ51GsG5uDFQunqXO1i47rt09/bU4YL0bF7pjfaEqnrYkRF6kO7MFnHYX
IICbC7ZidHaMqS2/8OpMf4a2ox++J4Bo728dgSJU7gNom9jlME5hPLoIpT3MJT52jjqBZqiRf+1u
0X9NT1+Pr5lVw6/Byxz6GCgoAc8rwvQrMhZHDnq4Z2FnQqHT+lO3h/62wspVj//mItbq43BYSeHz
sip3VmOQJHwmDeujUGiELJKrwOgtHFjnPssmL2Gaa8CkWi8nTDZnjA7oEd6CUE5bRncd9VvPAYNB
aPGZYVVnm5x2S8n6c+bjxIItU84rZeNHjzWp4xbP0k7KViNPxt0u6yPs9K0q+6N2hblBZIowEwGE
BZ/EGP76Wyh77YjZUhjJE8EG08CjvQa9PA5w6S+XiqNcFWsVa8K/oXYCMx4PVvg1rijO2TD03EoM
fxZe+LE/5cVXeTzHYBxkMzU85KCWVhN23+R+sVhry4nMVRb0Ac9K5Xm6pl1VT3SNz8EP5SW6u8Vl
0EhutEhj056501WembCFij7jwnltZ57qeGRIoOwmRC0MUK3xH4ZeyEklHIqHYRSc6m6M+Q5o9oYD
wSMFqW1bXEuXzyujFNeK/vsiQ37qb4FPv3q8teyH+nV91+aStjAxjqSxC6rsLN8kAsa613S9Y30T
RSQRQVbeySHi8RBfQlZi5ndh4JxDLhDYOoXo0G1sJMIX8YAt+LAafqrOorbjEJMJkHzrEKHq3yv6
sPgjF2rcGhrwgnLNTMIsOKREBE1sVHEalAOLzAJRm/4MaQhoxgEWqupHeh6rCw0fJw8NIKCDbaFp
Cpbw93FL9+y29P4XPjbzf5OKwSQJyqyFML2PwPL4aJbtq6stUPnkIglAmu2fZx6SASxPdWqJecXj
Ez+bQj7D6xnhVReD6BmsYJV5HUU/KJfCiYUS5y7OxgX43zCQCZEatgAG0iCvmeRkUAT/VXYvtDew
ovJpxF2UrLDRmyKcfTCub/Wgi+cpShaVCrwMpkCWHQB0ppTEHDSZdzp3ZvNxv9gAKSpgLe/UbYE/
OxKtjOCv+pSUFvGKX3yAVhbXp5TdtUwRD87dA3s3VgW2mDWazGzsYOCwJRtJLzi99rU9c+OjcS38
Gxu2BNUTN2K1jQCxx05Rg5zRkhySCc4e3ACAoqJ2jgmOOqctWDbfAxbS/xVP8wEXUNEQiDJJWdNt
ByR1H5WF/SPjRaeARqQs+TLbpQu7sGBRhwStc5yZI1HwvYIur2AuJ/f1HJL4QSpEtDsEfjWmrj95
78Cfd/O4vKHiBiCEEUStKx5ZZN12TIdqgKVy3ThEBC2ibLB32TyGhVSCksYwJARG5YHC8+61s0Hd
kLiH9Qy/2A+bYeHvfLsI8YVghpo/fq24nquKfs1kD8+Fm0Zz+Ps9QyaltCRazWnxrjGRco3qCHwC
wdYZZ83dkWwKjkt+IpF43nkhCRhyMncOSIVkVuMoTWKJy7iB9frib0fnvp5wxUW3pg3a+HPIw3jE
QN0Aoead/2uMZQJkCElr5p8Ow2cpe7Ndk3yG64GRzpmGrXmS3S4Dxu8FnoVVOGDuRVWJ62z5wXu3
hZ6muxtHxEzeLLw82ASQglHvUNGl2GNv/YzosLwnJdwaJjTXGHZgbUb7rocqyvNCYbAy/iko+EDE
8etvnDHR8uqOJ8+Vsz7NP9Jxby8JLRe6dk8PoitFumHxkefMe+7/ELrUFP50315gyvjLHbnsZVjF
MYSrdQBmYJKaxDoeaECfuwGcFCxmAo/2dL3cDugsl6neZN36pBRnbt78i4F/x8M0LR9KO/v9ilo/
Yes9ZFW2yH6yhKxslp2sVMLoU6pfv96qplTc5h6H15C4KBKqRhwDwCeFTt+w+luAIWFfuKK4z1Xf
SBM3PcNAateSKHSUwKZdY1haGhvC6N2HxPJH/ucoFjD03bAOf/Dqa9+P/C6Pzq94X13Avu9nap27
7w348Tj3vYWyrpBmlhvL2wKz7OAhZdRMSskYapENQ2fFg5tsWYLtq4uS36GJ/483n2ihevJ6glnS
hmbZJpDohvAA2mXcgZKCcxNkTmnk0hvYcsbZQQ0hLRXLOaK8/s6v/yElzwf2Lc/BjeCIIrimaRjr
zEE09jr+WjS3+sR31H/i3caBzA54BMzxeNCYSFAYgFaf9j6iS6ziV6E5wjGmTM7eqxd/YysDNu0Q
yMiMS0/bY/ZFcbSirssbWDiFDiT49+8Eu8wj7MhYYV0pOocNd+31QSvdJC2K81UtVmcgs9S5JNKm
HCfG+T7iSvykxJWlTSUa9W9DGaaDTt6lVxzO3eIBLnFuJmBeCHj/1LCPJyZIAewN6AMwjeNwZFiB
/qu8Fp/VP1/ygAr3r6vbaOuKVFsFnk4hUZptTDK5MO2nFovHJ/Cj9yq6qbtt3zDu2svvnjEyoZ6n
vdp3uUHN/6F6W4cn8gR/MQ5tiK27YfNvcdUC9YZHb0CqY0ofVDGlCTa0bCZlaAba0m7Eo70XN2Ms
2mIANHR8fkOY7rzB28R1Gq2fl2dWtkTFzgZiEPHSsOL9pubRQOd90bZdw6cMUmQi7+AwXeTT/cmk
0F4qzv2F9X0YVM8iH8kiMf8X63PH0kOZVA68LN3DjMXALFE+RsMfzyD5uj+6+HzHZu71aF31jdrE
WpcWj+UYXh1qMoE/jRdKEUVUwo8zD5a79AC4GfIgASpLL/AV7bWOGvS6OvJ/fVGsqB1ci4afsnAh
iS5IVpRAnNJYGaG08/fLHm9xbpOANsIWXhkAx1zWyGb65SDKoGa4j51RE8Pd+X3R3gWnaSclARHF
5PwzQhMHN9b8ydNrUE/ZdRRLqNDHYjw3LDkteif3ZmftoMOh6bjMVwHR1ekDmysPPngpehaRl2hq
GVe/AalPOoOxtFGpPCSQODqpTOLAm1ql5pm3dXqBKlsRbt+gktnGlIHjSmWSdXYIs3r4fFbzKZEV
f/9nT/Vs/Wu1/EeuWYLAYLg/zj/hKc7YnoyJ8rKESMY25fBuFRtVY/ooqAKFfezPosx4OdJ7nku+
cq+OoyCMZZaprIe8ZgsUj7tKmofPaXY2BNcJRdvj+4rrn+AJXwfCPWJmxTzC8dcTB7igjGCTp1pt
AtxnpuBZQUmapj4otTqQS1LL89uT6J2rpTsDdZhv5EPMPvpHMynPxPict9aZl+1zHwHWnc1fzUkL
mu7gnJMVVG+tcEi5S1h4S052/4cTvQj5ygRVttspUwkYOC/ZemBmR9YEwPpBSnQd/Jxr8TCdidEB
R9uTk6+S8dxtLUUAlhEMOlKT8J/j8e2TC2x1Mu+VOKA7jokvPZQQDzp2/fTJ0gdrVhOLFPX/EeV9
p4RDj8ADpOxe8aqU0u2Ws6l3j273ArCWohO9Dsfa0A03vIz2Ps14mzKu3J478eSabKSSKyPCD4uo
QERBrFX1SmavwikPXj0vsKa7PC+b20RpuxykkuiRDtYNlaHuv8Ebjxf0dMLnUQFr4crCE2BjhT22
8jlNqjfUhna1cvL+2Twa8Fsf+K3o+ciKDSl4Ic2HWdS9Oa/HvxL7J3AMBk86wLHYbgzNLp/nah3+
m6Ke5DmQXT/HJOgNdfYNzk+RhF89IYLl5ShM7KYxGcbHE7+38SmttR5qozbibpgbV/CoKpldAkp6
9f4K9SNd43dPdcTVtPNiqK4ns4rPtvD280Ip/6qDqLw7O6yQJ0rcDOhvYA9DM+AfJxbI+hBb0Cmu
MbtCUoTmmPzsWMICJMWN+rfNZnCGp1iAWb5+lueIaYgn1bjKSiM/qRBLB9azRJTnQn+lCKcfO9Zq
Dy6mVzqBwTVFxdfDP+GYvNR48miUf26/NNybr04y35CYMVExi9AegNhzdzW1S7hd6PiOHgSK8vFO
0bZsflnCsHFwi51SNcu8mt0XyxGNfK1egmSsD4xkDw99D15KOm4UAnLkjWWX6erdL90oPrCTj14y
0zsE+eeh88MOMrynoO5FJQEy4R3TzfhiNeVf1dw8Ijlu7fPLfeq1pqjAYr2gR3jGCXTSEIn8LzIU
jlB6D2d3G+VgXZA/0qYSWWheE+A55QB4DkWl6iNdeOtoimNmRsu0HmBfZyuK7CvDHYtJLwgXOi5H
k7jrol16tLC4DurizGOgun3nPyFSmVVKHUHitAFudkQLh8LhTpkPsliUPBWYIYaDYSugyF1t1Qtt
8qTBNgf803HQLuBAwQa5FOqCPwsvBohmDv5XBshu3u1jtpWmGFU1fQoMbzSLlrHk4YoI9V4ATwVr
F1JHewWCq2HXXwFo85DcMqKhtCaC27OEL/kk8r8gYk08xF9dJOJiOHN1vWl4ro+3yxRvgZLbmiKg
pmH66H+vSRHWNmTXMOXiNDFhy7tq8gUHMcQKvv0+IbZEX1fDT3w8gxO/37fgUqlGNETq35bIECiW
aFfLY6E/KPBi8dgUFE0L8A9b0k7nqklQzlKr2qi6Vu6OLRxAjdTRNQIodLd/AFX27jdT46wuVm5m
Pq2iD3HMuh/uymUlJFerRWqFNLK+dOR4lVyOXZ9gVaJn3XtqBuw0qji35AGXQD9KJFus9QmFnUqS
ikzLIBsQGK6jZnibo50wwrUbGEXtcQj4tOzRAAonrLVoj1IPCk7K1aUOqxPE1rD3KEjzsbxBmFKt
btGotUULHYXZaTimcS4vy//XNmBmpMJj6tA1h3Sk1MGvGxHuTB6jGBgz7dKVZ8Vd3swB1aYO7X8a
RvY8wycHtQ8kteHwRLJscADlEa++5UcVuaSnPPhBEWPFW76RGhD/1QdxA9qbwwkFBaTUQJ85sZdQ
C8OnlzM3KZEaI+PB9qPLN9bZv6DqjtmK2VWwDRlO4zHAUTBUk8asVAlvT0oCIJSM1ZDDLLRkiBvq
Z7i/aojtvqVLvFLTXuxA/mIGozxiGc8355PG/YZ2VlzCx7H2OBkxt/ivl+y3zEUV9r3Ns+15Yedm
fPkxGu7yzGg/Pa2H7+CqdZ445fNyzYmiSQgiZ651jYd9Fdl4CeVoghqO7E+8aY4vjW6NapAjLnB2
Km9JDCuyBsrY+T8RQmwvHcCk0n2HuRKF2sKJO0nFZNiUSztTuhg7V+p0yBmdq6AK3Ghf1qqhG0Z1
pYcTdbUmZXRVpG17CB6924R1SlNOIHqeR/ePac3tHVw7xN2nXmSVb3vJtd04kNfBnkhMzDcQp+DQ
jlm0EoVfvQvJ1T4WQX5DPbwtPCTazEjXYSaqy6+CoUAKeX70Vz0MqCtZ6JQrJagevFAOMxukAPSn
LedMOB+uTnQJFOfFhUjiFM9mXeYVG837srMby+dLrY24S0EHbxh++rFqYYdRqLsG5ywX6KrxZ5Ro
ejG4hGrFlJhQcAjWiGmfzvEXoyGGpHXCsoP6kaoBBJ2ZvCs1jf8/52MEpN0AKEKVBzNI5tLBZnKQ
PuSgjav+NcdKw316KckEg+eAm1Nhwg1hgvyfRodeBeYZ4RW2Q0oX/Or51+veMakf6RtkqOfHU1Pj
f5JGz6nbR7zdGO53C4L4H4xiTeR414HjgBbjUKTVxdpxEun7IZjNlVQyB9KR5si9BG0J8Hmfp8sL
94LQ1Fy/IYumCOdfbEt1TytAmcTjpRCHRV8fAyS0/Lozap4royy68SpIDuUbS8n0rEyWAJQ1F5+C
xUsuEvNX/WfUesmSwlfTyxhPPH1h6Y447hzPQ1v7P5N5kgIsRNNIibNJEcaBAsI1QSVf8wQiCzrp
eGKWU6/VDvJJt6JVUdBqF99zGsgSukfZXdyNOYJTqFE0RvZCPD1O2AHzEYsnbLDaZVZQNWakI31l
OFhnNOFG/yqKLlEnE43CZcZu4Vm7E9liIUaBD3pTcPgStL4Mv0avw+BSJAWtrVMdbkQxV0PEOW12
Q9jmO6rA1QuPCwBUoVXuzBpWm8HRoCSzf4MpswyQ7H0ntOi1qDhE1V6UFjscZlxF3KeKluKZXJnl
wXCxAv3SiefOI+spe1TKhK7xLt97nUG+uHBeFN7cReVGHWqDkgiowK2UX68wndAdRUONNfeWl6Or
BuyDgSVm4QNNKOv0xdrGH7A4j8omH35I7xpR8vfbW+L6oRLhl/sVVKCd3SZ4dA4yHY7jN5s1HOVj
MpZcOjhpcck4m0bgnuTwAcEZm21fah4Fzhlb6x8xjuU0UL9efKG173h6lWOM5DBUp+T/I6VrnQiW
Y+PAr5RG630eKXOuDFGRdqENeoW9NDG18GvuAwOF3IfrHU/PBYemdo0D55iPZ81Eb9E9z4JR6e7u
zMXgLiPB+9pOSJV+z4NT1xys+Pgs+TLiHvVxFY+kTPxhxVnX8QK3AYEHUY6pxGqnh8fJ3FzJxK5R
E4x6EcR3l9Sc4vXZT5tuAbxMa1pqxIiM82ZGm4703SnhK8eCSn9uGyT3BhWBM2AuKYpvKm28tuWp
X1jkpDE0uKpQUVv2p5hwvl/FO9e4hw7+PnDLDgt977OseLNfCa/Ejga4hgbxPG33TkFjKyIw3FAC
dSeFL5Ki/u3tJ127ZvI7L4nMxL5CFBwUq8QfDbYblG7iBtWB1zG/A9oNO7e32hEbzq0SAhpWV4Qe
/rDhX0rL7nfVZp8SL0BtVHGHw8iuAtk8zOh9O/vY+X3XjvtkDG8blnHe7e4pYNDIJba5WhQfFMOS
iPEanT/cii0OiMRMKS6W+2dK6mkMjVdiB0eSNWmecPqMSl1n8rWMNrwp0iTEiSX8nVmgSlc1lAPQ
BNWBEa2EjDQQHVyd/yp4zLbxpqKDPWRtjt5+f6qxgzQpHOi4/a8CkIjChSxg972pH3yaIKUSLTm8
/5nnDQSsH+II4YwMpbwG7mOXMM+bPrzyq6VIxND7vWe8uq5UbscqTLIZCw43aQiLRu0aND5LCFkg
kP8QMtvH6hgO5IW8VD7JSA303d41hCiI3NTbNvUVGmc2Sf/Hvuq7DXKi8w9JXowKO0L01Kz6nYCh
UPp9LCNsRT3IGVR3uQg9tO/Qwz5CR63TS/75ZQh7RY/9TMnugasbB4VLeACIheXmwEWawA6vXqe+
L4qn2g793LGLJtueSo4UavXdzLM//6d3cR8+lduQhIlCh1eR1rLp/VTIU2A05o5uaEB/mdvlRmbJ
s/1g7sPxdC2RrlhkU36gdI/5J1aEhRWtfqH2bRdYKkEsv4xOFpdwEleIH8+RstX/b96AII6ElVU6
FMzYHYdvS9bQFKq/32n5qTjeSV21Jie0fYp8lcEpSy4plRklZDYuExtG1dEPwLRzINsODl/0C3VB
SlzYZGAMwBl1YbvQ7oLabK5hhbmFUHmz2EYstnQRXwBV/zYTUTZqYOYoxmL19bJaIWWAVAjxu1hh
FBqdlaHTZ9M2yw9c86k1N8O5tyNwNt0sKLtbIziS8R6vl59eDMpYpEd5rgOGgGpjlEYg6LLXvUyL
5tUyjNXOT9/u3UlZwykRR5Z71IjMNmbG6DyeCUIFmYe1qoNRusXBH1HQt9fYnBnRALxxgNRzvUak
wXfKrGAruM6l3suM7958w5MCQZ0V0Pl2jwoOO93A/2+eILLWZw4yhIU2Gxepd3zXPQQdW7I7rVRl
kncWQfaZIcEV8x+gYKSXPDnZssDuC9ZD4XA3Vrhq3RxCy8Eyq+wnEtZBVrszIY1fTl+0VreWEShv
fv6o1o1JyUij761D0cRnhh3hBfkZt0a681HNDS5AQy/uFEIu0nB38M5IBwHJ30mlPtkQajXYQ/oD
1ca6snOF8Tdc5esxTsaiABqvG205Nw45dGgVjEQQ4vHR3MkhyxaF5ucU58EnsCc+hzWEOcdqWI7h
8xxtIOSvRnXMNuAdcuKmJkmnTMLDwZC66yOxhLQJi4gv7piGQtxX9sKXHD8UGj1XNjxlWKnGr9DR
aNNFGU/KEuY+ldoEM3A4EDXe/3yKL1lwQdGr3NMjvyNQC2WA/s4EGG9QfuRN0efavGmVxlACLFbG
OiyFahLhEgRdedgWDSjGUk6cEfbrgCRgQ6XVUgROnjrzSv14zsbIHZj3pRx/cLXRE0uKah4j64yH
49H6aXHy2N6GhPHOEGm/d9/QNbCJMbe29rGz6GMmW6zP3qH3TvZAnj7P1iGlDnyCKQs6oYHRQ/mw
iuX25cfUFGDk3X0cj4r3l8cx6VpDU3GsXS5hvWP/veNGXK2ZhAaubaAji9In4xwU2+zmI+YRaPv2
/sJ0LBTb0bcQQgpddrDUJiF3gAMOWqBG0FHWd2vW05aACyRhfaoKp3tbHQh2ZOKyCn7fbuvMsrO5
t8wfaaxgDGVCibztwwhzZx719xvGKzrrt9cwudgVn8/Q0TqpjTpLGFhvuBhgj+ogvykNN3DUS4NB
x9cA31vw3xlCeRjV3/9Yqvgnp2MO2HkNH8jfatXJV8mxqYe3qCezRiedGV4FGyDWswD5tFiwlI/Z
FePktAaFP8votYjt85KoIDSBbr2HU+5e6NSk+SqnvDQNj3fMiyZovJwXvkOhxNXyXwFbSKHSPi/8
dn9KPBOYyFz95jPs9BrnqZ4ooBq9FyyGxqFNYl6eDW5RvZR0TgVQBOTxtH/Mo6C6r51VzB8WPc7L
ALyC0OyM/OkRvrTTu3+As9joQw6zV3gD2az44JV8wgM6h2G2O8LP85dvTapLAwN3cilvXPxGI7tr
yo958rwZrnGOu40FV5YTQgJLB5ZrC6vXCKcnyg3WEMfh50EP1+ypxJGX4yvJR78rTnJ5ZBjx+A4X
HnGx2SYmM+k1s7sWeY02id219c2CAgyiqTyKODA90DNdLhIYSGNxdEEAStxN+Os+K6zog+XLukzD
4QMfIpsYXw7QZ923BR337hRLsZbGLKfxQ6LfklAdl5hrj2PDcHg8bzk+gRP/KXlYtxdr4JnawHV9
a3ArP7y8KUqvAP5myLOqRv4Ljf21yfLiZfB5vF8fi/wcyUJkXjUS+jClrzxaMZK1cR/Hob1FY/nR
ZerehpW94pojA2/E5JRgMpKIURGB0QPBKcEtt1YeuhugBKnC176XcxCQAApImt/9S9mKihlzoDCQ
TzZgtlfk6rXHivoVJtfCI/JHeV7JJLctZAzUJN0lDGPMu2sxJ28eG4cBKQS3NFUh2S44szhS4WYX
80CH1Djy2WDxBu5F0d1/f84a7S2cdDApr566OzPX3+wnQg/LKsgRcTgASCmwKkr7Kkq9PfMk/ZQS
/+ATvTLjELYK7uLwk9mEOQ16tHgUocLTXz2WjeCtD9qW7tBAJVxlHHABQfmWwKRtoPCrgX7zpUyc
1aoBPfnei7z4vLYZPTVHMi9RoGAV8wLverocmTPleZDvjWILvuNA21MnOJGvmHjPDY1G28S7K9kl
0eyF2EWmsU7ZAIvHx7NLqILlq4Wvq37ifz1UCKu4bh2sTi5T7/w/GdDIkOuBZc63dat7MDhCGgGH
f/R+jzRYStZ6SSDwerhlyzo34FnS3V8Tspw7Xhps7gbL3SOJNjv1PpigDluBCJqaPrRM5cg30mHf
QelwpUAnN9AdRQ/w3wF3DbuWkVOsLloaoIJQ2r4R7zEtIIY9F9pT4oVbovUwT81NW2u+rtcQLJtf
ns3bEOo384+5zJe7X+eVg3yU08kr+HmZ3dVin+/PbogsGuyORzFcUt1+hGI8kdfKEZMEq9UWqmt4
WlQSlJ6SreRiejdRiWSEX7WmKgz09VPtVv1ubE0O6zLVlO2yHZCgtTXraaIeQQq1O45UFnDPNJMi
X4iI+EFx8JuIot9hOHGMTqoIx0BhKa5enPAjma+MFnhp0DQIF9sxzlklKKkHB95zi0XhpXL9l80u
sg4HqVuuK4EwJ6a7GPTR7Xi+2bIv3mdVylIUovwnetBzFY65YfSFnkomcLPlTgL62L/n+GKEGPCd
15VBQjIwgNL1twyqWm2pKbmzGLzThuqEfVd9AF53TL9bUfrp9EUxR4Fr4AMEEVK4veVRiqJFOKB5
8E9T7s7VQ7cUvf71wvibPa8cnfXSdi6aT3PRV3VDxhKI0wbjCDqxcEkTfmEnq+Fgcv03rvgxYO9v
2MdfxXukXBEJ65XHwCjOSxChMlLO/eWEhJYxSc2nz3l292EsnyOzSQ5tyM1slP0x2qM5hw+uRdBs
cI14B6M7fefKLWSDaps/Dd7c7jygN37qqD6366NtlMc1Tji2ebJXFCy2tTT+C93I5O+fxHx43r95
GsxRBr6X5Cc6ChSpr+9uwOTTjihO5ckgTgXPg0UM2qUQTnXyxpuwWEcaxzK105ytqMjZNpqPS9wU
izQInznl3qh3SuO2y0scDU1V+4Ki+4VdI/dzPZvyKCAqPnAe+I1Dmb3AH/ISUazLy1N+m93PtHMk
O4dLRtdQgzq4MUsAQ7Qy9ODoh0+YkyqNPuUhMLURPDt1oQ8cGN9oAauU7lBpDJRxL9xjeVceQ0/x
OR5JgvUs1A1tRUSKaI7Rw9hjAaa5YnUwbnmZzJ1IODUQeBE5GNX+KAt1t5ITggBkHEIE44N6np3N
XlieFrAsv40QZsilMXiOoir+v16qr2fBJjpMJ0Hc24tvTjW0P6Ko7JPXm2IsvYQ3maFBQ4giIJwp
x7FRc8BLjiOtRzTjjJ4tD442q3y0dvOLCxmnSAPBbBjlN91O7yX21ZHUTl3z0yx2l1SkNotySaJd
JiPJ5VhN4Ep1cpPtx9qdGDU7v8GuoZs0sOLuySHVHc+3G7TsgT2jP5M6D95jyoY+CxRyJgB4zd70
e7yZHNkBmAljgWP31xZ9aZ5Yht0JmQ+RvDa4Vu+l/Hc5QgvLSHcdEJIIq9WONrCCXIfSFVj+05Tn
786IoH90087vF6sgjC3vGa6z1HgzNW8SimAq0GBoabdbadFbmbMun3dJdGcEvBY/hJCN39F3Uoma
hJplue8WNu3J1K0m3yzdfyPxFcu23yxq0fXeaFWO53VWm9steJoNjl0ZJOvANaAFQPmJrjm3gStP
eoup38VByB8PBdB9d5ptJ+hp4w325lrcbhfPKRWOexcQneC5nQyUfaLqvYa35CPuszbs6A+GSTcZ
Y79g3NS3I2Sh876XKREWLjgoBHDY1Y9ArENbmuxeZaxXhH6iZAqgxYejBWqwXXAP6GKIoVa8mxHH
34S4zQVwgFxAxIF8c2dp4UdxYSzSjQGDabX11Q3akw/NX38AD/Jhu2tJu7AVFi8UInKTXWMLse3p
Y4+CNTUmP8LCrXLcIwOlmA1gMuvykyVzncZ5k+LO871hYD7TxfLBHNpM1jL6qUJLhJZiotEBgeFK
maw7olLIYSmyf3wJqP4UGlIVwmvqQa0VllNKvG8df+vTufmq9FAh0JPwdd5cclumexBgBLiPma3L
XfMEZySkOm+gGu7mLvkn7R8cLxpEKbWMNXfa/BJjfDucIep2ouSzFShKUlBb4HZISRBPCK4VvrPR
iRO5QwUhIhk4/N81zOFtnMPo4WLnvyjfQY1AF2h1WLGHcY+9mcB9x/dSkY4UAT8+BWEqMXZ6u0JW
avkx7oyqbiqYJ9KKTSXSGnHaZrZw8xS1+hjUgHBSPh1aWHsXoMsdfZEi6DxEOp55NDa6gR7Lt0D9
BmvpmfWFl086/a4y7wbkNjXajBIf+/zq2PssPJ0hLShe2sWyi5QfGGmDV8t9OaA8haiaAG7byfto
GcI72m68YihsXyzNheyczudKQ5xLS/3xaWSM6SdGxALvoeD4xHOR/oOJ7EWxo5Z/p/xgtY3HYO0w
My6tIo3QeYpTmv/iBVNcAoAyhReTGM/kaXkekEeUcFi+gVamYie4vRaLxyAqQ5dOb3gVW7TFH2Jv
I1E9VNx/VohESENML3JKbVBVq1nDbczYsq0/iV1fcUn+S+5eu1LEqUSe42Shk1YRVB7xgVnOytTM
PKzia/Ys66JLYjj3k+t0ff+kikm8FNUfdwWgnKJrtyFM+awxITxZ1K7ysGPpqeR0grLhZ0OBHePg
nReJAiShNwoWDWl1XPktbjvQNCHeDGQonaVKCui7L0S1o/ArTqIi3j0OAQ/CGdSVc/211XYfSw3Q
rFFqbIjyFmPnB4VcxPg+R0safDIwobrAwYIYs6xJcfIHANvOqQXcEtpwPnix+7tvjt3v6V7KatRK
qhn2WHX6UmDesNiVMLKwPJ+fAsBY712qUEE877hJOhAHG533cTCynYbzA+OJFGwbRXhRNE5wISl6
DOJHbcvK55cDpozZbU+pEV7uvyIyeoVZQzeH9/uza8p07GaXkqZBBVO1SwWEsGeZCyBpc41PYx+1
8npO2dZ0FvkuRSP88hpKTZ6fXFpqVjxXAoQw6nKOZuaer19cfRoq7/Qpl9Q9PScbejhCz2f1vFGS
rc09abetKvVShsnFQf9cOAZ2V+IdK1etjIUzX2/0FnHQwU3RfTpM1pkCzzLaj0wCrrgECi2pJdva
Y9GPWPeRd+idzGKSKjDb1VgOLb7J4p1cOT+VS6sEaWJ9LNKjKnt3SBvN/bEqQNalixvEPGSVGaN/
mSH94UsicMql57PC0gLXfpqP1wXS3VUlti5gE8kvZZQAeuUqzU9rjpBHN3U8wOGqx7Dfzzpp6YHM
X/obEhpXILVC+OxoeBJB4DpixH7IeN6qM0BZPJpFNuw6fQK3Bu6uWIs042oATBoH8EN7slMetHgt
v1GrVG5k3FJuYpBekbMMukTJSQcFiwJmz+GfJtpch/qjiryqO7lqtcluR5YP7tXw7dMNbEN1pdBr
T8n87DhfT3DjzSI1OJNtvtOrJfVAcG8wvGI9TxGFYF5sCjlm2u0UGgf5QcOCsoo3vEQPT0X3Ffro
XCb69MBaOGxLJd6JS1fe+3wqh6kNj6dxbfdUkjlCfj+U0moGjGRJbiKzXz4ZAP0krRRNkOL0Pi/8
B1eZaekP8/fq/72ovFnzkXD8WQRBJ2fI+tmbUVuBnc96QQbdPEgfEOivK8z7zRoA7IwSbqiOT18P
U6jd/yfzkuafwHxndklsCvOP2W4KNTMjG9mVWKp/05U5ED3ZUAXrJ9Dj3KFs/txBSL5zd8F7+2zm
M/za94TrV7nnuVwBOxs8Uf3TjNRFRQwMbbxs78Db82mecPW5aXS7c6GBVGeLxavwCaBWwpebDdwB
oNZ59ej0u8Z6KC+PCQh6nih0UPqhSrry8jOShOmAfTw8EUJoIr9naf8h24BiyGSrj9AbL20NxtAo
LYxnUT4pdvaUPrxlOpuvUKEdLD6m6UmQcuNQX1wfghyMdx4TFSFIkm3iV0Ag4i3fHyOzkp5IrT79
zNV8dfSVVCQdUep7gkhQ0fySJnlqj60SgpT50NuoegRJvmdCqYizfgGLgZJrqnve7eZgFFFye6Dq
hnjEn6KSx53Z2rUNnRy6Z6uLVzkqREb4ODBkzhVpG9AnPXjfUrKF5Xod5IJ1iP1TjRQ2fFyCgBr9
Oi1tX4oDKcg5bpYcqocaxC2Em39azMpc18NNOv6kKbO/AaDGIbsTkiDhCGH8IRBHP1Y8SDXCiDdr
z8B4R1tYDhAISf68A0o/JTYDIsIQROz52eaKrPeFvJTyFYqA69Lg09haB24BJfik583lE4fPz/AP
/B3Yk8zBZwLAuX31uC1JGsfZ3L4GoxQ0s13v0f3hA4aeMWB35VZ05wEG5ZMvfl8RvAJzfXpi1r39
kR7gUEiMkSzEm5QMd7OW0AxQA3Q1Kng82Fqy76RsWOF3SdFqit9H02Tj+faiDKMtyfIq9gkmwKvC
0gQg9JAZP7QJxRvJQUwwcYQXTu8WFVVYJMKalT4BRLPYf9DmZfu7tRAlXaLs5r7nQlSlCpyfT8c5
Nuny3gqp4yHMHxqg4RTCufi/hX04uIKYAm2hTkCJGAmYUP1qaf+HxgtV6YKPN/DaXZYb9DAJHM5l
8n8MPL9v3GO5bGhYMrGDNTMRPOtXRCJFkoAoOiHfRFk3zfishX5FLig42PUiz5zUwU01/gJt5j3x
DIHhcx8ZAHeLZq+2rpKVoFY0xJLnFm7SyCIXiq0qoLyztP4RnZe/HzFZM7iFiOIZRVlX4UK5+V+1
uhZFAaqUkUsE0bjCj1FRQicDdEoCeA8s8ZUj+89s1XLlbSMIF81SKto2o+mih0aD8CJj5VlSYXwd
ubaNi+elkFqTr+Q/lUspSgUBOoICM1nyvNlETl6Tfzg3MC33SjH+Qz1Ibj8dPDWPiFHuZn7K8eYE
MLlgdzSbtMmv7xSSj0ovOHe5mHi618ZOk1Jg3959WSwU3xz4yiehvoFgPSZhGU7f/D3SyYXu6uCX
S24+RTB0DrOzfsTjIhbijTqyTTf+rjXpBSeZcivBCsdfKipxgO2YAJgBpdkkxUur3FAt+lbhrmN1
bj/wajJ6Ns4Xwq1OLBk8EPg/a1fFwbPFGS+a6Yi8g8nVWyH6ddNz8zdozklNwUaLszreQ2KQYm9c
99Ri+9TN5CRFasm5+ISlncJs196I+7LOm9NCDqc7vgsIbF8D8sGw+UCtURb1ciyHOZ9kL1HtuvvR
V6vx2lC1R3+VTAW4d+MKRHspVTy27ApO3hIUonUbEgsHW3+4l8bn9PWVbwRtjjHyBZK0aPxsuryt
4SZYWfG8T4Qv5CaTCiIcIDu5aln+mvXZWqSJ6qGKoUV5gcbxiZtCzHInOG4IL0WDl5z0ORMrDIRx
KlrIe+jae9jwgsrtEvnCHkgPL3GdwL9PvGLzwgTQrRMAADY1PMdcFXhM48LcwjJPJhyRrobWkRP8
Gt+1eMcgM9FE7ERmlv57P8S4FWHy00On4qgJs+Z3kEctONBG4V+NxzHpZYz6L3unUk2a0sbPp50A
V404OzgdMpdA/dxfjjZ8aXuMsu5GwgWbTgRFMIQNcVXpg/7gMJfnFuC2G6lBVBV0FOKC/nYTSuSD
stV14W15wVY2+vN/U+PX+qRGe8ATDgyINRbbEY9QELBLt4jlpORm1QzsbnYsgZNr+5qKt2+bNw/w
arcWLQAqzI+8JXK0CO9Way9An8Rq9t2Hz7vq4O/PxFJ9E35gXQZldfusttM8oWoalhLNV+kWLQSp
jQlf6ZttHn+wtQFPDhn14UkrF5FDohG5TNx8kqrf8nyvsBj1+8cFw7zrnbzO1X1VsZj+6yUzWM63
3kOSvcGlqgY/9drQM4oUIOhnvTOBtMhaFyLlSOBwxNJSy8R6jrtwDuwIqtfnMjl7fxmbpQE7OEDd
e4gDL5j/mCEWTR0NdUdBe6De4kCAg803eNPwZWAEWXievs5wM11weG/OOM3+rNFMFg0Q0VPJetid
NMhw7xaOoR3iEEo9m9CoxGDrfZt3gFdYzKfvjKg5RiWApi/Q2S4qlXPIMmZOP0+wTvkvwYWb3lut
UV55l7QZwFaufMl+Boj+yoSHMBkh65jsnAmKE+AhdECm/m3ylvymDA28g9VsBqNiiOjcjyw6WeRW
HYpdBDWqPR7GhlHrWqzR/edlGiZNzmKXRFdKIiLbjQPdZwbwZGqmdkwFS0Fia3Xy9I/vIjxmY1/J
KRy4A+E1jtykD84QypFAObQmI62pDqA+Gv+tgfRiLkUmBShmvulGDMdpxgvNxgymo7fW6iPk5wqu
9M9laIMWMsZRaHfRSQtXxpEL9AwADhWk5AhStk3bFeROUmj8ri0bsLtMyJwxji/PcBhEbJmHalIl
2F5G5JvX7SVEqI4OOHzC7s5uVcg4wgyHRFHyepvkWSRBBFt0z7XJRvcyabLxlJW6f4vy4QHskytE
gWezYUiU1RxtPfq9NmO3gxOJXnJ1X2rJFCBzWXsBPpjyJUjJ3rBoetVnXGf1aHG2SJgU+q+09IYV
1/2ukM8gEQsXAY4rCZRQvRACWbVVa/7jBDdua5+36XFvkv5TP0WbBVH/k9tqUKlKpImePJ88WLwK
CAqb0B1D7KNnsjWyUN+8ysKpD8dalhC9TmXNHz/WBBux8/Ab1RYfcmO8Cv9oedu1eybD5SaN6xKR
IfOHDt2wPeF0sq7nO2fToLU0plf0HQgmfzIoX+InRGWkPO75WI2haXTjjY616015kjUkndYoHZpl
VSbVVoxE3SOJ+PYthEI6sOAbO6J1wUIZvD2BO3NjR5oKb5jQo7UtqtVO1vmLewqelpYwf9hqr/bN
UiSjiLqm+3DwlJnhDROApIO0r2lgpw2l2kFsYpS3A8pIK+CclHdipQneWLuC8k+Vk209Yx7zL+ll
eh0CF0HU+Ec2ibslA0e17iDjaXuSZFUTKCnloYb5tMoO17ZYvV3V0oaONlxSs6gOs8wkCljWUYyb
LKFk6KZMISagXh11yFN2vNOHHdQrhvZD13uS+MqadSsSpomrhtsEyi8iuVBYaeW5Z/33EZtzAEqe
ZDUWkyYFUZqCTP5cmRqxxMveNRr8aR3Cx2yjNTwtR0fbvLXkADc3HYoeMs8EPY3Kw2M1+jVpNdNk
3KJQxGw0BUwMDxJ6Udhhtfr4k9JKPE+N5fpUi+lfA6PhL3cvx9YzM3bkBjrmTK1oGhxIALIUo+84
PEyNxTQ3OOaMnvk090WJd68VYfOvbhRKBZL5Ui5wFsmYwMJ0rzRG321TxXo65KfRQ7JQ+hz1T5pS
dEqrA26Yi3X1rGMlYLSm5izRvqYOW4uw4TKLEN4cD3gEjXYDB8uP+2qpjZqc7hQeBSZPELJf1x83
n5dfn6ILxdY/QMWDwax5B6IG2Sbiwr3ziqrFC+N78lWlOvNnY9TqXUiABXSs7ynJBkxTlWi9g5rn
0IZ4S/cHc/XE2Apy4EDPiX2jEzRPFBrMCEC6WqimKdMjXo1Eq7ZEjhupdWhPumy/FB9tcmrnv4NA
AgXZxXzqheNsVpE2WLMojj55GbWdwQaD3eHD6r1z9R/VrA6l2D4ZHhi0ficcu1JeuOt/Aw4vrALf
c0xVyVErooYjsx6m9TYRtV0p9qT5O2PQFuyDOWp6lJqaOY9grKT1hDYUqRJYzQNFUCziiKVRSJDQ
7jP6yDgTAzerXikgzVLbYSbeaGyBuK73AaBsdmnG6Ue8qfAsquY904gnX8Bokl1Q1fKaVlBHCNCI
lpJt3P7k0oBDbqIisaEaUvR+OO7fxkhrYxPG8JLBYNLQIE/OYHcHRxbZcd6vWU6w1EdVMbIXE69w
FfXF95eOg72sREDoQJbd5rKkhp2zhPDnhzC1RRBQ3DkNgrGrxFmmud5zz8LrPDwgi4bGs6eF1AT4
UK3seIq+g7VQhxIP5EGFvDRDPaRPIV10WAZR1hlZCcKMbub/fBdraODXKP1FrQ9TJwDxU+EEVxpM
KwdqFgO1R+K1vZmspi6fbzbMvuGe6ib2yCyOnsKteXD76nFreGny4fRcnTeUTlGnKXk9Ggr82/Gd
Q4MwMVauq4b38+4LTMVU91O46FSr+n+NlNOApNLjxK1u6taZqcZrNxD5xmNf9gzVRF2N32VfKqFj
JHv97JE4pOEjnsW0ADA4l4Zw2k+XckDV1AVado0OHNr1apXQKQyFUeoupcq1yfDOHykWIo5nUZQh
BlzDXbSsEcJRD3/m94mH3+9/mU8JGAvHRc89l1puqpA0AooM3VOiCos2AvbGG4YrvMaTggDSnoYc
dW2D9smGoeVn5uXZUL7Gd0Esi9yFOPnFcJqtHwq1Qt/mj/9eoYOEflCwZ2WqvRVViESRm0YuQm0B
8R1Rv+5JR7wsuPzBuDXvTgvuooHqS/C6juOP6Hffff4K93bt0+dOvqx7LZkSadmoo9xg9wDl7rsJ
ajq6OTORnKo6hts8Dh08+aTdRb2/bj/22L9PiOUOgRoy3UyDL7Auoum+CcIn4tmedvx/zKIOB3u3
djjGsIYPa+jU5YWKjBpNBMaZw30paD3h847a9VOAdIinJ/DYpcA3h47n3QNzfrce+0KnhfBS8bG3
Jm+jF4MXtPzQcm/GpSwduCEKfZtQCF3tLTBUtUb97zCFDYqvmW61NeMjZqGq2NUibgy2rn9c/BQS
C14lgI03D7MzPTSKohKwyLCjQ6gWdnHRvmKYi9H06Q94SnLzkYCmxbOirjjIWyHNMuQgo8WyJ7BR
DNuA4fqxzGQpU6GxnenEYmsJM9nElTOq2zlfGf4JIhKjjLgj2x3kBCK7VPG5cEoMghC0/o+weRUA
/QXin7RtIt36MdN4prRfv5yamiN/5FnBYm0bh4J5Cvo0bQaTYC5WGPs2Tuf9rGacSO1/7QEOCLRt
3ThIK3IEjxmkG47ouvzTXczLfK0PN0yWUmP+1NnPkaI4mZCrdjudyREMAygkuSEiRFB6wf9YEc/U
IYAWIHmKmX4TNSWcUEXFYKg48yVvTR5Ut8whHEBtbLbmHR3MFbB35AvT6aj1g+cBqLePjDojB+tj
xkcHG+wcfuEwVtCRVz6KkYP5yDJl6hKiKHatQr/zYfvVj2Nm23qt8D1NXHYpa8HRUT6kGMvaqp1l
h5/WAnK5ZUx/IFBZU2fuhp2vxLArBbjZl+mfzA5JYHVPxZFSz5WRpt6M1pWllwTHmW8VK/3SF0fX
5BoXRZ+eFcYt6eYo2HNw8i3kexKEvNomaoVUBhv+z/mWwVP/EYnt9vULnaS2VLvBsTHdL0bMd6O1
Qx3cTU+oKc/3y5D9wrC6+gswCQaPSlasPyuMNNjemnabKIJSDo7QwTh0R1H0hNbqfJzKE+T4gCYH
8UjecMDGMHYKdlb0vWdsQYAPXTZt96HhGYESYHrXdZgrUDL1zx4GQPfoKKbR32ctRo0IMmiuaGJX
9Fa2xMkiWbrzJtDyxWxkEZZzNr/N8uadYe3THw3fVM2sQ4zURRW7pxmr0cH8yoRuLvBCppC2WxDH
oevWspc7PnB9Xdq+ir33QYZDUD1QFQhc2Yppwlv/9pF3pfyqBs+VkTQ8jBv7neH5LV7l42yUlhSj
84kDHLrzRCLum8udfWwahclMz66ETcWzWJBDvpW5vfhCxees0z8AAKVY8VPVbIk19P8GD5EwxjMH
KqSjb73Lrrq9DzVd4RMo7ICpZDgxkHHKKmorKSpw9yl6Isw+ruOmd++E+wz+8d8dPGyHyQsbq7z5
/dVDZod7OkSHQ+uCWfmzMH7TuZQJ5y448xRunN+ArnzhpsyLneTfQsLcZKfvQCodbccKzTkw7hXz
59/dNZ4cTYZefxk4nJhCUIVjX/ox/xaP8Hwi0HQ07+sXlyjGjND2RG7zsS4Sr85liSVOc4U7F7mr
Wz5DqQArf8BwrvPsAkikYj+kvxcJ4YIDil1UjsDVL3S7yBd+lOIKfL8a2YgrLncK4vqJikTkFWjE
PZU0a4eAFXvcGHtXC0Yr/sVoSJs+Bkl/afoa54P130n5I/+QUw7CghJkjQCZ5ITwbez4Y1R9FtYL
E0f65+e5Ed95LvEbULFMiJB1hnanOR9nStT6TZGN4Y/MLjbNGReHzfPiO6MXRTuR9rvflRLSqD2Y
afZ3RTttfH7ff0kOwx0GQ951ZzlPC+iDd1BvMkxp3K8mUSTuWmawy2JlHB+mrO3h/b8FpcwnvWTa
HyAp1u/qvMCoK3oXHd5m6aR8/gVhRe5pIRX02bkFSgvUd4BxtLBmwNIPOz+lzjY1YaAE2RHZP7PL
L9Ir1mpXIFX5Gng1Ij7yxkRiFq0BhU67bYW4kXcXo7hNJbwybzjqrrVzjlk73Ys0r31dr7p0QRGz
m91K1w7wBnLSRyhrT2MsJC4Z3oynA1Z2mLtgEdRFg8QmAlvmMJPQYeJKus8kEbq0LE9Hc4Hy3ho5
+vWiRQi+rPlOGdtteZwNm/ru/zd1L7pMzm2LEnCRduyMXLubz+AUsROv1Aq7jNuzx7T54ZdOj6w0
8ltHmTEjEZPclI88K4nSSMnyLL3eOsoKxIaJYJjVqkmsu0HwAF8uAyCndAU27aUuwrDRaha4kTbg
Ng/n25gtKYyO//xvV0H/0A2s6ztcuTs2p37Y2vYAAldhJUPIlVV07Id5q4nVH+RWijmzBdaU4GKc
xu2fErI5rr3wuen4iv4E32qqwAbslU6igQI7YwDbpMGcnGm52DIBsSIMCip7ECCutt3XmXEjubVu
FZNzWZ14GVJ3WZ2ZQCUBntwy57QP4RQj7EmS7S+PI40Edq2Wgl0+bqVrPuwRcSFqsRvxQf86F/zB
s31w4USvMOOoWhdkZiGbOXiWL8in+LqkLjTl79qBHC5EUIvoVMMH6OGbsmLFcjGA6m4b4iIOB98B
mztU9aInQNUVO2bkCXoa8t4GeZOzh9kHj+eEiYqZSbHI6CjfqAcMXKbn4XyxsAgNE4cAi8rsl/m/
NKOrx5q5VwkgH99NT6rRN92v/GRRzQtEKg28YyfTwW5jJXK4KKuI6pP60KApfG6EwsrEiFVhHjjg
zVFhBMYbGRJW9+F06ydg3qNylBfjXrtOpkb50T77IzwDo5g8fdbej+O8PThG3MPnnB5xUCAH6nZa
P4TxMRxkjeYETETF6znILU1v9FN+heWpCrlnJygCZ72qS8uKg8EjbF9kzWynNU9i9MBILqpQvWgU
mUMHezL3b3IBoGmX0F+8hBdYscuOVSEccNPQzTS22zR6fbAGklSDgBKDNk/Zyl41cN7ve2hVuoQR
pzoFoY5Jk9LzchUnEK4+dy4f5K2VkEN84TQgGYwlk8M03CQ/978HZJ7+Ei/jh3j7ODJVjO/E7c86
sytH3OmRSoZB5RuHLep1SiJaEdaCsMoAfnS1ooNjOUdLPJrcC6aFrCovN84lUvVwJhH2TUj2MbWC
tlXZ3dsuKBSoQgtYgG5gFuGXdGxuO1UOUNv3j5QJdtFjFvZ4ekZSFqQfjFgeoFAOFYLIs+tO1tc+
dzLI1wjfeskBDuIXOnNlQFVIOtTc1q1FwcnS7N2mLGZOBv7MfB3djD7uNNBr6ePxPw4YWoB/Zchq
EHt9njEOkbab0KO73/4B132F2CvIqeXEyXC8mAkwrzyuEQIYXiYnHJR0X5i0xOga5SFcpR32INap
uqyTeLEskA965JV/uRwj9W/k/I8v89iIAdRos948Nzda7yK6UMY0GjmlDbuuC5wJVuqHA2aszdw8
2/nkzrJi7+nuG5GIOA70/2EbsxCaST4ooVyuEQnenvK2ze8iwkoh9uSEa/xGC/Brfv49uVYs5ohS
uN9yvTBSliZGpYb7ZF/uovT5wakXkLK+aGW0cDOK9N4PXzTJ9bJZdWRrhHaZXuKdKwCYs/eDy+hU
JAQ+C8Y4fV1wBZ7+02GPn6RZ5kbL69nrHRuqDsoC1ig2b6ri540TzH76s9PvcAlaC2V2t+uON5El
1epcxLaCDlOP8pCdfU/NaDG2VDiSc1VyToAQO1Deusd7yo30EK3ASs5bc1tAJ/QRqghMhFGWZUXa
Qt645YVN44agFEilvaNozWPUR0SY7go0eVIU5qbVFHGexFC1Qk3/au+EPVGw9yYwujPuFrYVyXQV
XI86BLXnUR7O7Lmik2pMHK6zalAy757lIFfKxy86bAsXr7cJgBpbX9++VF7JrSC4rFuKeSi+cEzP
Pen6wSvkg7u+bin6yWTz3KcVFjpLDU23F9DmlsGAlHr64+1kYs1KOWLAPQEkzA5dzr5earWRkuVO
u4A/GFCxx+wwT9LTvGIz/m0zwwbUeYWF2ntLC2hI12Cz92K3+ub9SYyozGBn550g0aloYpFnRKkK
LBNsvPjolIrCKluQylcNmZ3VOFXmzD5xOf+RR9317ty7/Avh51pi6muPiFAPVHgKesLFpTDTGeKA
TTfd//HEoClt02C84zsLI/mjrKX/jYbAJ9fZDrBfhzutwIQkmoGKhYbxIzs3F0+tZX4dTDO3oUdZ
JF5Qpwt7KYVrAw5egAqxNcNHPrVm02LAWCc2zW5XUfYmd84MUPQ6y4k+vVg++tSY2cPj6bRk5pjl
HUzb1PbZovLPUY9hIAOwP20vczOjQ9vaQgvbhbOU19sU0VQl+399vIXX5DV2XdYRXpVce+hvD8Lc
V+DAEzbGNdOvS2jUz7v8CLX71BaOarFGVmVxrw+GU+262UjeVO+SEmI9P4Hjp9dxvLaEwPBGbJ/y
wFh2y3ClA6nl9O5tFJUEVLi3tDKvyK6G6bKEmhwdQINmv6MUZw0QoqwS1EIsm/S5BnYfhQHSlTRJ
xZ1a+wzOkgOl9/dxD+Y7KgA6kmiH1SiVxYCr8uf+5Ubm8WH208MiaJouQSpIuOdCxYph3uBnNEK/
qzXDh81lNfIoJphP1iVWAC3OjsgE8JjifVHgS6AKtpr78zxn5SrhnPjQ5Bwu7NJrXh/iwFW6eLlr
f8pCZOFs7X1gnWaf2ghiGuUpZqmx8+TsG9Q7bvdY2zdm92OhUSdz5LYdIyJB2fUlhjisZQMMOvBs
AfeEBhuj7Y3fUSrv2cjm/VYRMxUu9PGQ9Ez1QUZWdzFAUl30+5ayF8qZQ9bcG5ollAVgFMQKLGd4
7nzVeMVBpJetXH0wY6rRpV7mEVGXXiR1LxbK8cHMcLbo1tFt6HsMxwR/6/I2MXGGcKgjBYYiRhsB
Syie1y1Nb4WJBSavU8lGKqOW9cYiEcK1enSyAZIGa0fDBvQyq1K7R2UDoMalW57MBlqZfCNT1hRP
oJbURQOqcchwDMqyRpCDCGvLGZv/tHHRqjnFULl2p/k5/dgC/9DoXt+7qVT/1THKBDn+q2zopWZk
InMZwevvtjv7Ho/uFFHTKT/u7amVgfVNfbE573j3o2kvyT8tlnGITeo5g2QYfye2JycdYG/NCGm9
1ZxFil9mzJEiAy3kbowuC8yncPEXgXx92DoT1J4e4JgY7E2Odqou8wuODmXSjUK02kRkOrVgt/Ud
yjKNHpE2ooF2AW3V3Y0ycS/IWGuP7SZOvo5wX9F7Bma6WTz4TE1KWxfRKW5pkOuLRagJYEewNBzK
0GHXhFkbbOsh4R0Qk1M3EaGiUM8EZUQeVHbg44uWnHg7dtS9MjNXCP0x13yiNc/j4tt3+CL0Lu3D
fBg4yhb/xTlKNZzNoIlxJL8RhxrTU/EkIL4OV/7MJBFWedYrmZ9pSHRdLJSZI4/Hyknq3vB6BgHR
Napl5ypl+h74VJ91R91HF6RXGPHYHk0UDwV69KqPqqkPHTAMCJSuuzKa/+OhIXgbCvFozsui3iAV
M9k05f0tKWU10yDlOnU43ocZm+K/2AaUkIRjVxJQZ4bPkRi+CTkbmCDLF3PxMkl4taLrxKdqQXd/
5SSwmiPdAPobAR4ShXbaQ+5ARP4YNhugLlnPILKL0losFLD6E3jY6s9euOLWsjRNgHqIpSx2T3/I
DwSflwK6oKI2gdvQc0fnCWyNlooeA4+0ziYuUHCkTtY1u+xKCzC4172C2DZGrnl67EhOW1Ud3iHG
zMGFxZEdETxzycG3aZD95YWdWs4jQnfAQL2gfTt9IP+hYWxAm9KxNzfeNq1YTr4Oa9aD66ZlbX2H
g+GxPVfNfS2tltB9dSKKrKP6RJFNNv1c7UcxfmhIpPqzlQJDDpmjLxqdMN3xbXFr48sJm1vck8VZ
7dCmuJmR70WhxWB7bEqbK+ZwgZtb4shV5MVZuea4Fx/3meDOKDK9erupp/t35xe+nXu8SO+JLn93
ONcRO2CLPLbHD18FKrnXnzRSHK54BOngfWv6EFsZ8897jhS1bnn2UWSAgEeRPn8GEEVlJLeQI4Jz
01aT9niJu0p/hhRiXaodz7fMscpr11qs73AuMhe0hSPE2St6hWsGypnKTowGrwUbLqYdk0GRvXbf
uj5wNZ/lLRwGluxsP6r+8rHiZEQPmkS+kxBC9RHJnclFi1FIQOQqnMgSTGoKTwEDC1XfT6+ZQCrv
kERRO8qPmtptkMGEwHjXtzXnzX7YilLm3ZHSsNIrye3NEj6TE8fFoC6PJWzvS7FB/9XqFBzt4PQN
Q7YlYA1Z3PJXGKMW66MAriSIVDT0uMXInPBrmf5XB34N3E/IIQ35d7QoVBHuYRHXSsMT6XZ7nxWx
W3FDrbOCzfoI8OXo+l75dufUTjybZrZJmtVIdTnbty823WjUt2T4nW8NP5ydEn0FUDIHJI3TUL2p
1+sFJY8memqSpiS2eD1zg/3hfQ9lkswYSCbgoiqi63XQuLRqcg5mFDAJBAIvPwphuP3X/Gm9Ic8P
eS8E2mGJr4zdjtDj9P73LKTCIHjGdV/LflP9GZAeks61VO4XQ1iHXj+xi7jtPiYepFsr42jT/5+W
NLyxssu+aDiMZiA6lpR+SE/blo1oLAS3NtXSkH1ur0bbutZkFHSVBlzJeG12WPy5y27cE8yk+qMF
9jh6ox3/7/U7stiedjaTGYAW5xpVHZdttl+FfhLjBnvo0hMQA6u8YUAJVyhUz8ia4080D1IplaHH
s/Ex72Mp563aUi5VYAI0ixyDE1IMSfEmEFgHz9Nd3Mscepo+YnFF6eDfPJ0jMkcbGAKkc1Y597Ig
fdbhPL20/IAgQrdFnp5VLDXMp6+fErR8BYmkjoOwyVTI1driOW4dhvc2U19xJXnjcBWPAhaCzpap
T73wDMjpdXu5W9a2r9ScLP1HvBxSf+GQ20xsfjrWSCbS72SGD+ZGCvWNgKT/abK1azSHQLXa5Ax4
rD+2JUBUUmEdhMor5YroqrVbttI+/7Bljlruaaf4lJOMU+daAs6/9zDwrJ7zVNSjlqiXY/WXJbel
ieeoVfmvfKXREMiUMNnBJE2tm+iXKQRvWZho6ZlsLhuIfjUtUj25n1AmCfPzi6I+AqpDKx0J54Q9
JJXVFBIB2PiQLltk72FFCtCv+e3JOa9Kwt1zdlLgKI56cFf/PSSgAcNcdCymPm/rRYtDTJCctdaA
Sk9n7BXvHjb5ZXX8PE68wRN08v9JTd21hJgvyZB/TsMkVcRdoWvGMdGtJPaH9lduJjQF1MnIQN5R
TYs5JrF9H0REmtK4bz2vfFOJnpsISBfEG5TULVDSzFyYtz8tvnzzXU59rtdkfL7+J0lh8rx8Vo1R
tm/0hjPZUxOldMrk+UVXs/5fKxqChnAze0WYP4f1fs2d+JNPrIpx+JZF+m6XBzARJe8HFlxjsE0+
/PiPqqs0vLIJNPJN5gdivRg/b+b6RIST9aCDg7HqMAVu8JYI4yPC26gg1KTDuHtYirOs3CabGUFo
g2DiIn4zMLsSvgp+nGsK0p0Zi9Vr/e7RAbv3flAg06wAt/jZyjnk+f2+6qtEXahNyvbqHpz6lHRv
fVyZR6KsP3gWemNP2mRFHoODhROynbsF9pXLPZ3CincEwoBBa/196/zld5Sebvi6cqQJcWSUYqS6
vldVW86229N2kaPc/YAiiDJEIHvynqc4BOdoK3g0mlFQCVZvqp36djtsqT4UOrme9wrOtz0i9nTa
MQr+vP3+fo4kQb/Ubi3AyDJ08adjLvBKAWbq5+Vene0MbpfoYU6fKeLWUw0WaGDYpaQDzKEVF1qk
YeSYlb6kU6o7gDnU0gShfr0l3RbiUWCXeSzsGsZuA590xBAabTQVd4Hm3J3g0LgnVgrt9p+/Y2BG
9C+NliNhsrv56qdQEjN6Of5G8gmJMVQcN3XtEuTW8DApvIO1RgkCaH/D/YsaFNX4bKVxIQpMcUr8
qGBQmvbl+/rxss0sCx8FJX17+exBGaVYmrOaTEYrqDmgSj+4SgciVmCDAZ90fqTwsdvhXWz4r1YU
NPMYYZOIsKykWcWmGVSERVkNnX5lrzmLh1RyDCAD1VPkrK0cgGdXRHNX0lNU6gJmiV8aHTxl3Cd2
rWCnhdFaSN9kyVQwoE+LNfN9idap9q7ccU4YUP+2zizyCidpzkbzk3WeTfgq8jpZsm/g0AFmzrRJ
16YKyd5LuThszlKFxB/9KWipSKN0jYOTXHOBIj9PkEUI4mMyeQ6EnlxiFbovmqcPrMo0YBdmPYVY
1BaYBx9FnojEFrfOgtOmyacMcMVpW7AY1s/gaImwU/zYHxdZH46q9IEElkHescNyvQ87QkSbOCht
jEn3bKj0SEUZ3/3VHG8bDA9YGeoeBlcB/6tEWvI5Fi6BDIaux14pVq80TPmfOTY3AE+lvzXoGoVQ
5yxn0Yn/bTaxAkjTYE+Vid/97Sbtiw0QpeA92JkETkAEBT6aPq6SymXvvX/IjsmkY52F6CyDr4vt
7i7TMgaZQ2fT7UREEdf7KwxdzfYWxTaF0ySrVkMV5CkQmBLT16FSRnwD5/wet+p4JViHnrcyLj1U
SE1lP2Pr5YXsbhs4ao2YNkYFBX/GMoRdj/idAj6E56pMPkf8fLkTFhv4OZyFOpFUPYriT4DzzgmG
JG6HtmBjAJ6xnNX6J1AvDpfBddmqWALnPpNwXMP7rn1wnYx28lV4Zod2sZ6F1V8/bCV1nUuOuIe+
LF0wuAko2xkYbt66kLq/511Wv2amOiuPCAlJklYhHksKxant1t1esre6sMq7RKwQTx4YUtkFHs6z
RTJE/q/ks6103SK7LmKj4/cT0LBi9AUP6+zCk6RgkelJpMik66/10oz5Rnh1k0/I784KDUMTuptg
ER1sZs210i1R96KxFvi83f89ovg+lPWwwU8DgpydzD2N8AkvA50T7mWtUcx75NdTwOwC5t6CpWTg
UYJUz0LYFfGpFHs/h8XBI8oAr9S859thL568pwhE972K4awSBievAEzaDqJmLJ60r+z69Tf9y99U
qiP4GoNYditXJXuCz8ChFqhpqjcfnntM8zqMYpyZ+nMe/ErvSW3xVEXFgSUa41d/bwI1vO75btFl
wuiolzU8lTyzXA+Uby/p6GEB65ylETZRvKA0HwXKFsgCEPuF4y1GYTl+ubX1LL81+MvqG+Z2vnE5
iVuWqRo+uEJRPgDKdn72UTlStnMZJjnqzXKhi0drX7rLyfMaX6DsJqdM7ZIz0DNY2btdaBUNmmWR
DwEoW6AklPgPVTQ8Jh4A7NcvG11wfLMoFpmfy7VU5WpoTiKaNslMz7JmkMTy8/QY6Sf2CjbY808B
7gO4GQ4pbU4O3ViaZ0eqxPuy6s6lgcQYAw49Z0kjHC2Pj7FK1+HPWKBFBziv8fKkyX8vV+pKl8Gh
OLL07iO88gGjaqKDCOFxEbiyaXLr/+xltKLZOYIr31xru7Z1+c2Op8JmDiMey755kCovJG3Sy0kB
AV/IijXRCsbR3Q5+mpTZwpnAHqitDRERqLqcU9MAW/BWvwYk22XxlW+t9Yx9vEmZgcvhEECjbC0f
5SsAXWcAMZSciexfj38/rJD5bkeQa1P6kh1AHFUzz5GNiPd+YxidnSz1+dMt211WNqeH5SFAdBZ1
emmxjnVu6hcG8w3TYLHvEgLSvnQBaHAgpxTTOgwo8zfJGgyVS0MKL6UVhtJ4VkRwu29nP9wv1y35
RpVS/Mtq7puTmjNKt3DedK34LtWz1wzP2sNAnD/FwftShaXnxR1AF4x2fN18WFc4Odp0h51g0+Zn
+9rwXZQLTe5ief38ARZbdQyHTJ37DGBcGVagO0AxqxhYQeMinoTfpNCGETLbeQNNg+lV/PpskoBo
lf3chn+XxSiKU6Pq+WsUGv6o+/Rj8/5Gsr6Mu3bJtLtarHb2a3tCAE4MffDZ+yNxQIOjk2YwHv0G
a9PfQMgRMYwu9irym8uVFi2tugFh+uoOfF8w2caKSR6DaaZsbnxnIVmgbzLUaaMLFGRtgoLL2Sb3
1qpzbRA0mB/VKO6hA7KCWF8RHIN7FzKP6aisYUEGgHcMUEIYfRNAqvIReO/rtyl1Zi5GAvf2TY8J
B2tOdLBKk4Zczo16QGIXq2i3AIHtxlRNdAjOa2DjuI8GdqUZ72Tlz9O6x6KaHY4LjRmV9RVuPmnw
lNSsQT+iOdIKskIUcPYU0WV/SLRpPhIx5+DHNtCKkHXhWV0ZBjL6pB+/wQkVK2r1JSWyTnEnLpgw
N20oRofU2pm8z8WTFtZeiAGfF/pLfRSa1/jhVPeXJlY2JwimICdv4YlEX2ecGIjqEljFdsZB+8L5
Xq7DUOJ+856qcVdHkDwlC4akYbtUg3M0dOAOg/hLd9kfAB9ZDdnsAfP0LSeCr93P8bASjJ3hVQH7
Otuyfhp9PjcJyEw8kcZIq77Zi9BsBTF3qNeeKmdbWCZW7hONcad6CdpI5zqRv7FUH97y4lrYYeJW
2h/PCDT1IxcvMnqDbNtV2vPJvbjAC52NcbABUyHKh/KE0EjZjUPpZHO1LPwXj7q1MPQ4uTX5D+wF
jKAPS7Yc5c1+7xx8T2OmnW5WTt3geyRjxEsKFtg+ietqElYbE1/cZWYY7/tRIcXdoLfMmJ01BxZi
eGm3shFgiyEVlo4f9BnEJMEbI/O9Lg+/loLg4fk0aW0rZwkLZB3S0OQrcYHciIjwwUAVYyfLP72H
RRPG/zlVs5C0g/0FW1kiOqM27qd5I3q5AcxGgnugSkk+A0XPVSmSdD7NfU8FjibjKw2iN9glwv/7
XFK1AvFk5V02eAu/nfzu8nMhoPnFo3qEIKPtritorzqlMsEt/A6j0uxg32HRhdN5IB6ghLRC6pBw
SK73uE63Z350o1Fh0wwgRkKw5D86YPNTPNNhkah56udPZdgAm1SbdPtB7D8Xe2oSPg+0Dkq3dUge
NBe/hXfEWqbQ4r8xxasFiwn2sKRvyhJCEWDi3utr2E4PjNgXysmxZXLrOwUDjl7Bu2jE0lnUTDsT
N2f2m+3SWhk/1mSvNrdTktfam9HoDTWjrmh4KB1+X9KH+8NU1ft0ip0V3FZ2HToyLupqsEq5LzuE
ODQW1TxN5INnvG7id6rHeHHFdBxIgJDXzFP6n3WAtNaE6v8teipOSSjuuznzBXGr1LSv8UwhRIpx
pI0Vtn4XpBJ5yNasrc1DXhmUFZ0ph2UjVKrZdsxBRo+JsKiz7yf0LqV5lh1aMjhGbs5vu6TJu992
TkBJMCsJkphHteyZUv4pbdxd1Wcdjj1MwkmniEVRxvb/x9yQ+LFuYATZGjcTUEhtw05YZsVnuJZ6
ySTyH5Q/pUwGbI+mnOaitQMReTd/uaX7bI0uhTzvs+kJyxe2uHhRpljPCRYjkB7ZXiGgfAj/87Cn
orDALyaswdLA84gcW39UPB2d40MBtxnZn1NQuhkb5jT9uFx9QWdiX6t7x3WgkBGIyLNymtObUCCj
k6FBSmyizbVcjqMAiVzPUy8LVyJjSY3Fsy+lbmhA0m7vwrS1yhwW+ArQbVFj9vaqlOnxN/NcFS60
knLBsY7PtQotF8r0D/BYPaf3rsANXOpimA2G8azGmx68GCU3FfAktfHIdy3xg4zQfDPPd7mVNI2C
IYsL1p+ywspdvHfhwGh5IEFjQa1mpFQa0sUsNVupsSYDb9O3ETV6r8LaZEl9JTw0oFewjDZl7krB
WIwozEC0OROq/xReOokH9iJjsuyut3gYOa7373G4CQITYr23nxtxrGpVVGLTiUGiWJsEgeRk51Je
u3a30UslBdvk5HSDSVLsOeio9rlJEV2GFdcfNH5TkJrKab8z/ARG8bQjn9c+5YW/qSPxcHnyB5HA
ePjRW1lOPxdjUKx/EoGKxF6xH2gm7fJkw//JJA8ZXNG4JMaQoOZl6HtX8TMfkFiAw7AVuCZ3DcUO
YJVOsXQNk6TM8kxsTLeCeInPmtSrKtl+MpTfHzPqa2nvCUeRr6WF+9HpR4C8FvyyAG3tm6o8tdSg
l1A8nVw8EzFh3S8RAFXNWuCQYyeSZ5WM8bKYJ6fEMQIFkkBRPtMGFFZM+h7Z3Ct6dnedTl0TDjC6
ru0KGKM2XEGNFk34JWk/waiAr7KiIbAGYUipDA6u20gUNU7oltFhjfUKm14x5BgpCwsRzdPWUW3t
GfwBniT4FJVniTgNyYVJSvQQY7Gcr/Mh+mbK8KsioP99JPz4Hzxgp9CAsfULXMMw0ui8gIWfqMdm
NDYHFVa2N5ZkoSkBGcGYIkDk44jyLiazN/jILSL9UuhChT7sepmcNwttuAUeV7LN1jQ6VqBFyznt
Z2FwETwe7a12Fz3kRXgQwgyCTj3U9rAgLXX0QCauc+zqEkkR2pnBc3tU2ekl9PikotC21NBmjvst
UfnYrQSMnplDggNU6f0wiCEi6hMe1m9u3l+f5U6Pf/Zw3nMRfM5JMonLxvToZZs4A/evS/Adk+ur
kD4eQEWDbTD2hl7/iJwGUH2+2EX6I0D22hDD97gsWm/4l1ThMi/A8HB/A1Bibt4qupzXsFHxvM5y
s/z2s4Kd8ZnSWrTBHG4ImtIKNjJHcqxnv0//aiPSxknOfLQESCeQ35xNzTmclnTcw7yOQJnGgOp/
TXTEDIZ4CKKiiOF2RfScbSqbfX5hlGx8zoEemuOu6qA/JCm6IZGFhO7ieeRIFa0cZgEH7MgtTX/H
P6fXbBqvx1niEWHhG2dm+X9Ti1WVBrCbjVvCYkVqd/hwXvV/oOe3ZJ2+SDhhHxUMUxB3JH2kX9Z7
YORttvcuiTiPeMnhhh7UYzNXEisFCklSSBgIqltzaeHi0S60D8EKhTil0S1+KArzxXt3nqZqj/+d
+M8UuoD4fgiBvARC4UCqhMn1rDKlocjjalaQhzq8+J6ANM3NyjuLhwky/cYhiaPruqDQZumvKpoe
VoZ6QB2KJExJJUdykJemzqmJYbsiLzPB5tnwUsGFBuDH+ig47UiC+8ZXJcWKmAS4Z38bNMKC3pYs
5pUtp/9iemi4XOxDMqeMHfp8ZzuCa2ffJsKMT9AlQ4DruC6gGfGnabJwiVNlAd9/sUobmtlPIFKb
ql0CAWTAYnq0WUUUI/MuRF5klR9jRq0wjZHS6UDy+Wuna4FaLOhq81nxdI/uuzglmj+X7Q/laAsO
zAsgiiu8XAlq06pbWVciZqdQJMekBnOlLyuYIcD/cQBcxcjo4H8QA3igy7T8YyStE8IU9C5kbHVp
qGlktEBSA41fjXo2AmmKk+kME6GDoDIS+FjuhFvbesePlbMsiDaGlCZsCyI2Ae9CGG/LtUUqIJWE
g8xDWYifr6gopb7ZPqYamalT19+xGmLSZZ386EAyXZQxiKWX/h2r2ywA6nObXlqHSiKFp4yXumAh
JaUuZd1JdsCDM5zjs2coP7D3K74tZ80VM70WMJXn3bCWdcrR/4+/UYaETYtw9A1qyIMcgZsqEJV7
EbF6lYmVxMMfXoYZG8kcmidrpWZ7C4CsOe+VueAv4m6sGIgA1wZ1vIETNTjUoRB86l6btR9RkHhT
8904hO5S/Kh4MTbalpaf32r5KpneUq0s5QzD9bK8/u2/HIoSqe7ziWtLDGTrPketf545pwfDAWiP
vHuMigJo84KpUb2FF7f4aF885PHHxuQvSfCGDKwgEP8hicMg8M4CIXLKQOUEUNxWcFnsVql4gFXC
QoQbgmLWNQ+LAA8MqE0JoSQ2A/1cMG5uBZrLNmtxjFrBXnMN4kdbXX1dXf8MIed0SCHDMwivtzx3
o07h3qvvDFRA37zcix69Xasq+/t+h6i+qsgotLocgTbQGWPbhLByXvz7tf9Sp4SD+cc9CydYOMz0
iR7X+M5L3a7uClvO1f9SI6e7zqS/KmiE3yOzhiRBIhozEyEYGJoopMtB66x2EuSWrw3f0OUPS/TX
OcvlpybNYcrP83tOr7TDF5v5Wo7ZK0Y5kO3B/JdkmyoGFuP8snj/9p3L2mH78PCzDouWXuTvxwMF
6Gb8oGuHzWdJEEcw96eopuImwV70XcAilMfIZAkoUAsxmoZTW0081i4lxfDNWOst5klRLwUB4wx/
S7VZWB2hq+x3K8cV74QTB+eJf6KxbjJ/F2MAVVQ7KpS3nHSNJaInXsYfZjGO7035HzF0QHecV3w+
bZVBo/FSDrHTU2YVoz9dS2d8tZPKG6TQc4NbZN6tPBFd0ZvKTP1J4tSgz7IZAJ0abTU4yfsDGazj
VFTHmcLFvUXlE5Xfc4RmmwXWzTO7JlqIpm1Kf2AZqwIRYVD7VtrWmhvJazGt1G30feWFYimSyDlL
v/9D/2adtL1h+U2BYJ9cD4/wEfeVOgV7LXlOugJequcLEHsE5sdbleePpSuuSS9FxOHpV+dHYK3d
VFcTUB8iF0qzzeOI/xKxtrGI15xm7/ca3dMyDx/kUHOB5rYF6aAPzCGkhZZ2keX4+uCUD6TLYfbL
QTpVzBTXhm4UHFV3hJQFta4wDb3ZCfNV7i49nK0Ww6EfPV6G96Ei1AD4RZWQS/easB0t0zks/PJa
RmT4QeD5xwFdYGEQd/WkIlNq+QRchPaF46XmOgcuk/fDE9iUyDjvlUnU7lDWVCZKYIH0NVhyHCZE
LJVzGSPbK/GtFAb5H15X6iDfISvH2+kx4gI1vaCQCc4sPopVx0dCD+s0hLFFqfEfLL8tHQRJbDLr
CWSTBmbuadJiarW9IWgiYo2Q0FjJLE8gYqbujf/gpSy+Pe+srXgfGR5V6i75QTbrIWw+COu6/XeH
HwBX0kSe69ENgCjhqRA61wmbZTXKmhGwlfU/6Rnv0TN7b48jflmF26cYcF5+3fgq3mtmRIHso3BD
ez7Rky3zuLVUjr2w+VMvxbrHMaU5+9RQSY8zlG0ZStmKITfdyrV4XD7qK131/pRstYb9OnGhLgQG
O2bTni3l52I3b0JS6CVXpK0uwGwPCkFPcOmlnq/18mTE9Mel+4soMtSIBQcrjL1MsmTlnJ78JWh+
7/eOJ4hZz81nK+mQjGefAkM55WIf2pOlBypozQ6pcM5t7S6gfo8YP3WGZRq1zxqsSKcVli24AVZm
14nVAgvxZV8TtgOLxYwhUKX2BTKq02BpfYWoopk0s+K3R0gWYwa+8pna8puLz1XLcjmpm5nnKy2O
N3rRnQOPAka7ewoVgLeJ87KpKA8YCzf7IhUC5Ejx4T1DqCJPkh9LWnGA3dKqWXg8YabXqK8LXo0e
4RBbSllGlCzZTYLK9rC41vzL7Cva2meuR1RLchTU4ABH7qyX9wGlJUP2tgvr/6IOOo/Er8b4s679
sNyVL1YERlTYlqO88ore8yc1+MxyjgdrVYQdffsYzrafLxeIdehyFPc9NZvDdE78qAXASSMpwCFa
5TzhwNuwXBvZCn02UZakv9lFIT/BrAlBQXlr7rSEu9mJAs5bkZTlN+jM/eaB75gphKJaBf1wXb8+
uxSE25/X6xPULdmvznybd+X4mnXClJEko9nsAvHP/Ffzn6G0tvfctWmgu1ef8xqNcCWAgx0Oveho
h7bXJcXypLxBPDh/TsgdoauT+yZs5ijkPbvtA67M5cjjpnAxABTO1dZdHm2WnGSaHbiOX9lK/om1
dlx3jrX7sm4pAz4UnadVmuoIZKG4KRkBCKvYwo4MSj5ffd1f6kDEOB0vPQrWiy7rSLgJbC+IgHWm
oIJdTxMZlwwdgfxxfx5XqLTSpnTzZnYxISwm+OpVC6wOEEQiVkEoICH4Q0GpyGxxFI53fytQ72zf
XSWs806fSyAcSfNTBTSM1axYNau6Sbg3aj0JpzJ/5V5hb44KAFuokzacAx4uxSPLNcww4Ahp1C4i
nVcKVRLlu1cF1kKh6gIR2FEpKFGCBcqB1FsvdZXC3O7ZoItQrasxzhC7K6oCw/tUartJkjZI08nF
n1hkxD/L3r5fUL+VMyGidxIvAY8e4XRSYiHfw7v4AO8dEhyD8VzZVCy4DEJKmWCVCGsfH8EXGZuu
xkKZgU6Ky9Ld/wWWmf9G16OZO1GhpvR3D0A/2SNKgH12saQqfCLPf+3Eu2FjRA9gfDDkt8fSZHjh
wDfAUj+OnSJXylv+VYnxlUV1iArYeVD0rAa8hpx38JfFDLtViN5m/V24cPAqcxHhNoGrc74eXz8s
5pT7LsZ0hw8tAEDFDJkKMMy24jYKWKMq+VuRHABLZagSBwHkaw6oHppvKJEYR0+tP6tuTESbGv8G
Bne5fTSEch+2KP61vPAaJWT6nSLhQ/jxo5LWuL8DV5HDdHIyv0/VmX9iZNEBUd2XpqU79VuDvqH2
dxLBOjCx3UTv1xpVqF1JN3Gh1NxP68dRt7zSGihJNTMkwOYs+TiAA93O1ie1xGbB+sPpIl0S/DcZ
diKTHFbRfCwGQyRmqOJTnfe5INR0OMs3AhhYwJoJ6tNJEG3ASAevoCTSThaVO2cPClkvsyuWJMjx
MZYIktfFZcLbEttUadqcpMrjq1jhwjAoHJDwgueJa/sq5Q6mv6zHuas8RGJISm5TuNHNYvJkS01E
9Z3TW81cU6bIkVNNYl4tR12Fozoe0HI6RB58Oe6t+8I2tNMM7wd4X+HaBlbdHAtIbungZLIzWNGG
3lOnb2xalMxYoQm+CL1/YDtk5bRvu2QY3QnMI5Bb8Bil3fLSIOQuGKxTzjfo6NG5PGdP0wT0P0Hh
rjwOJ6fo3kUHi+bwov7H0Mpg88wsayXWJ6K58euPLtJGoucbzz07gMAGLyFD/ebKNHPAVB2Y/7+z
O5ICFgHTHQJMSydv1JaHr/SmbCqvN31XD9vsHXZ9vQbrVIr2hCwz6KalRr/j5tH0AsilfNeH75h2
NffYcJstlHEcaq4EZwI8rUJjtBJoi8f1wxGGWfYS/OW2nwrXkourfzyY95ISLArs0AbZtVtADiP7
p62PDjm60LqBvICTLeom1JzWjLl5TAHSvnwWl/7vDQqKTl51opQ/AaPHYMuA8S5JK+575WTGNqYz
Io6bBFWFExGt7OcI4DYaejANXCnCm+xkt3/oognQUjet1XpWRhx3jlc9cUMzGRE09fwo/7qeJAEO
X5l+X3wngr7xd4viYKawSCPPvikn4cG3cOWANIcUARUm0+Pa46f0T1HRLjiT565qn2dcLLAXG3I2
CeFPlnJTs9thF5k5xoRRzwWUsxYbAbbvSMoRgBgDKFwFp/x8jzvk1jA5W2VzEB0ActuFkc3OiQPT
0nePcQb9xmXXAD33t+BpbKHbFo+FW//6Tn+OOjz8oqRB+5D+DjIGS2AB+1+AAJc+75zXZa7jhoB8
WDgfl2bPngcS8ux1e0f2A+hpdD0b0AKIYjkHDdVd5M1c04lYzmF8LjRsJi1jbuK5Jowb9lJ7Xjjc
UWK0l1EOdegO4i8zhDda8Y+uHW8H46hHi8fyYbE/BG98WR66NlGGkIEY897pThijIsQb4jQVTP/Q
aiWLCAhXgt+F61rq2Pw3Fu7jDqP8nif58bV+nnTxwgJ9fyD/HIeQA2letYa4IdjXFgcGnJfIs6Ff
ZhFbYoyQX/szSI1Js0FFGndvuiTLIa1156XO5sPaIeCSLHhumX0igqurtqyTeERHdm0QyKeSkPqk
S2SPF39FqAfXT4gSnSBH6IcpOkeI8qxbbQ8OJFDhgVeeCx4jlP663jTGN5QlKwhM2/SDrXt6g+lV
Tcy3EVKSmfh9+e0sjJrExHlg0LD+MI7uLgVf0iDxXTKAEUtctfLxvc9afdyi6sybuIiJbWfNmUH7
9hRymrEQTNfwRzKN4P+OefhKpi7IGpLTAxSHEOrcHQxVC61P4RUKGq6wj7TxoT2ao1nm5w9dWTLw
bWh9iHV5rG/W1D77YrEE25LbqH4M+UDIlrUsCpg97FjpNqOJWWg5aj0fnMKFc76amjC/xN4NDetT
wUU2fgqNOlApiB5DHxlyVnuBVRicSTFp4nnBM3F/M2cftt01baGEtQTMaTB+Y+rqGNDgW6PZaBCF
usy6B5y6BAQDGkYjoWhveBF66GywQwYM2SVpO77y+HRQoRQ8pNVDC3AvpjSt8CkOOGMu8C8+uhH7
xVZXm5hblt8CUstOrKxjQ369Hm3WLepQ4SVygszpwDn6SiG84UDfw44l2DKO/ngXb/xh3LOB//Br
8vkhSjadFQY4rwgCdHWE6hL3c0fn9+DKP5Fpb5Af1dtsOuNmIDtGQXOSDeSt8V5TVHr7s5dFMHRH
0WebOf8Yc9RqUQyctZYCLiZmMWCjAbIvsnYyI3+6i7+5bMQIRzmCFzc4tWTU45O3GX3vQh3+oRlY
TrJisraay2HmVXhi0xge9ZCHPv107vU7fFEQR5X0hqClJYGHhxsW3Gsz00jF85qKlpkYCjVU0Nel
yMY2aF2T0I0MXz+zxzyUourv331dNMvwohtcg0FmGah+pWa3nhI4BGldHe6+yGaMwxBtOC7c+YBW
jNfEPuzc3tva1J5R1k4gODhVyIgi9nn7Dk/CDRfGjxAbp3in6UwY1HCZFDliZxo5gMJNulN50RLJ
tgqYla01bBnBl/CrDlDGLJT2IFLDDR+N1PBF08+G1JNRKpKPT4KjLMh9Jeykxl09uT2dZPT+j7d+
3WdWzgND5xuDc+NDO6s18ysTH5U6PjmD3lRjgFHLMjaI4oSbjrzOGdbzGoRWM04Fvq1j+T5lZqjN
4o+5uomM1gRXBYNTDJl34AOMCHsV4FYyVXqyhAlVnGOJmaAMWXZ4vNC/yP022K2OXV5vdcgKfe65
1kZ+ze3QvPpZxZcwkF5elrQhY+LeI7UGFJLEe4sjEHb81/237TS+m+E0YIHKtbrDqYxHf3P7MkpR
LdNyvt6U3YmY8OkCGuMDjbZ2PFtal3nfv3rbnlZEeqPnexyuOyL5vHvIrFrbUVH70RM1G/7lBp73
P9cijpzge8ONAxFxIUJL7DILQmYmqFLtUhCDRnUswYBZ8P+VM1CtEpVe2AXzi+0hfvFWuiSMilnR
5GZ6dv4RRQ6fMwrmXuuhDI/GzF6cFvYeQf8tiC1TKZrgPCC+qzDZDm7gzXlKc/eNzVUcCxfQ8vRj
WfUwk9msdQqtliwvmBZWxTrQI7m6RuxWKaTA+RhqEIQ7gIzGfwoLFcox6coHpUE5ghVl19qtZ4V9
vaR7rGzZX6DVNqdgfI1OYpkVahS9ZQ8VJjmoJZYbNzmrPREwzhzFySEqZ4pDhfgvznyMqj2ohGNy
UfXi7P8eBAetLwtHOpRQfFoWi9Nm20q0G6s2QR/7aQkglvjDHM4GEhRg2mg/w3UGEM9kLbw7RIB2
g9qCpg/9j+gwybL3YZNr4R6W8DKqWayIycc3fTgYCGZOF/fSV3+oE8b7WUCr1uTcv7pA2se90Fe3
7DKZp9I1PPSvosYE/Ld2faEyGqLhMU5+q8aFHEU7BJ008vTIRfJyS2It9LpLmF99o6QCYqSYLKWd
uS06+XFceI22EmBtSxI+053fvBw/NcbKZx3P7uD8Hvz505GijWyuIWXnwCF9jLUFVh06uVc7jBZk
FSbpmj+fYBO9C1+UrJuQ/75FPZ+p/0fJCiLe/i8y2XFOSKL09QfEfztYTWbvEVcVQ0DaMsBFP6h3
4Tw0JJ8KDx6fn0haxDMqIx7Ly3EhgLWLRYOeI7yoAITX3NMtoN6rbH0I9qhTKceycKA1fyIakkaG
wI+zaoZrUrGsxU6XHq0/w+7ufTB3emUbKxV/fq4FhTrXka2mrc4tN7oWHTkwPrSdnOoKY4/Fyrjo
IH9Hq1xenqkhVj3NeOFHjU0LpdhdpwgTXNHytAsrcxSAqU5dMXylYl2Z1PAkCxU62lLdrgtjdCxC
xGDHgJOQs95FoHvvm58DX5Y653cr3W111ZAQpWg+oKVCvLe6BE+yL+tWF1+vYB3ermDnHIF1VJDn
Xc4us6qF+qDsrJ9Ugw29/T0z0qVxmLUvtzCVhoK6v+V8nxKFfGyiJWiNi7YziIbSJd1w9vqAEsDZ
DosBy0L9UrVW3NLsUWXsmXvZeINpryk1hv9BpopOhjVmPvOxOO7h+av7TqYpJJcY4bH2DTLftbOX
YzlDwIQf3YUqyZO0Wt/okNyw6ExvWyai06h3Ho0WmzoiIGE79ix4p8BS1SNPNinYg1iGWD0FWo4H
qYnFE0P9sHNyzt7f5/3tAmJSPnZ+iEecB4MBVdgkJwknYNi0dn3Xf6bgJJ7pzEt316iXJDBC4M17
tzYvsxV3eZ/K3WXPNZjEDZ70QugS0CH8AxTmryBHJFKp1rrzSgED7N0HHq5VhYoiev8tPbcdtMsh
QwJorLjk5hjNcBIfu5AqrwQWHGRKJLk+KD8O4PWjN+CSTAa/v6tCc76sYKNma0rWJ4pKlZzZ5cfp
/y7jEBKXEkjMxNdsHPYAprpVT8at/IoNqODXMg0VbxWv1Qh+CGpEPn2Slu1QkaRZbw4ElYu1kBPj
WmqVMIzXmb2HhbE7XhJ22vYALssHUP21YKrjewLeZxzrLIgCGYWjfu5JUWUxO9NQgcbmiPwJ6Ekv
wzgalZWETibBB96EwEd5Z8FlEh7OQ5AOZo3doXFSYKCL9+860SYTaV7n4D6V8qXrv+QZGi4TSLZv
mEZQN7QS9YuE9iN7Uv98bflFcy/p0TbkpbKiueplUULLK0mywSXC5CUJI92UW/kwHnOqor8DBuJn
hFvJwSiEmX57INFnS5BO8Ef/wCUUITDxqiBBYFk62K2smJP+a6Rs4Pp+ELh+RTzdMOpJN/9UWhbl
P/ypQMEMMlyUnXM8EYWJ7ilz0wKUa/6H/czwz5iDEFmoaT3kGis9p0LjLKJMNNyOXhlokjlABI03
Je0IX9TTaBQr2Srrb70q4WanLYoH5tXminCY45raVBG5OgODmbHuqDYNw3YdkRWDCULzSLjcEd/G
zXmVUczuH//bxqBFZiARnmoP0zYWQ6RuXG/CpR5xlln/08gF3sZ0vV3j9UkcoroTo9KYwPwcCf9v
jQCSn+G7i0tfAa6AoFZbSPyOPB/4zLNtwxlrlQ/wrF87B3YkGz9Y+SxBkvFxj1vdtQJReM+Chxdy
wjIU8oKiQDvCO1oP6z8uoYR/f7o6YK04kV9qzXolul/BeLzve7GdVTCM4dbdhZUlQKZf5O+rdcsd
5cx6xUabzjQz65MGMidKPeAKgHQHw3IV81MAwZuY1Vzk1p/iGZkUipc2YfcgYp+/BeYomeggyjEv
uxJ+EJZWucyQAO7E3kyHzOGVmBjoHXZQblycO1vMkKT6BnxdKMa8wNIZma2OMINueVASWG1Oh7sp
dkxlwj2l3NyHaglg+tZ2M/wuBuN1F/msiN6QYiHMCRlwThOqO0wWcqwYWXBon0N63tbg9+BGXGAR
3pRs2MkMip63/qIaarI07yWqi3Yer+mp66JYoU2sOMYq/8jS3+yXSbjE3xwWK3x3LlkT+b8aUPLR
qALvTW8tqfIO4GULf0q7o0s9LeySJj4ltv2W3HlJQl2vJXAUN1EihJ7Aoxvw7TUB5nSsNpiyRjbr
2S94e5WLEZh4NtMXiRGRucqrwfdlIT7bwOgatExsmt+kvqw5iXZdnDvkVEgDX3OSAF6aXIDiktNr
tIEKG5hdL8aNEAwHt1tJWTpQQ54zh4sXtffrubzYcKu3DAJyn+BcK1Q1zjFJgN4Xhc1jdf9aLRa3
qfTg+IMexjPmNWhM8d0gLWILEDk8eo57l0ndbJywn3Mm/PrmIJHYbivsbGCAAr9+kZbi9C+2Jck9
g/8WSbAY6prnmlYbtWUMO4Inpc75ufaQbmlVg2pjBGu6wr6q8pFcPRkbknNn+g/xEO08az/eKt/E
wl/A7fhsuQQfFAGKzvD/x+eFg9w2PhMON7nGINXlHJuFWNOlrPQss4VcGHUot9z7yYnWXfCKEXww
WwbToLUtwpyLmL7JeRCGI1frgBZvbDRpoAGGLrz3aKfWsNT6r95sHHKrPSd0x7NnVID+A6zfPBDZ
uv9sIt5JlsTyIpi0ExoAjtmHmxneNZ4dkv2q6fLfITvrW7odDYJiRrQ7mo3TqYOEUIWsXbzeyKJV
hy/57ZBZ+6lkvpFyfevhDHaEM0s1fD5THXZpdHmAcSbxH7G88gTSROqZ/vXOvFXNii2HYIcmRDlq
MnPeg8+6R1cURxp9h6KY7ZB120gFhRrwnCnwNts0wodMIAykudBzIo4wQ8/8BM89yWbRPN8bBurC
VEiS0zwmKVTgUq7zXfCnWpP+lCknsymS9vbclZbDl/5mmONzZ670arvVSc8QsnjVCczVjtwSDSUk
izaBtzDoJeNiOskDR5v3W+9Z2sgz8rW1hfZv5OgicTCirUvD07EQp3U/7BEMjbjdGRGCn+iCmPgz
sIGIUVUClzDWs8kJ1v+qQ5/NxslqYf8SZ8wHhzOFysbt2TLbsAFEotA54zPLoZ+y0ERWCmEYMrz2
WzwXLsUFkxxmSVnSQgdVN+pkYO4/OwcMSmecALUC9fiRc7OPrFsR3Kav5QMxP5Jkk7QZPFZmHaaN
xfglwbTpouebhXKuj2JGkgUd8G9kxliYhA4SmL5oZt1hKw8qqAHmC/HqAU8SvcpLy2cHnujEMRr7
dbf3kshANJ30Njo4GDjj2j21tI4tNrbbMzhEoytp+8KwMK0gCy+dd12zmWqUqXHtRvgSzBh+xPI+
naEGet2DuWnIGqwP+RHwlwhshrf9WoVstlQGVc88KF1Fg98LbMluirJJKG2gbPhDvlqtaRnsu3fk
+Ijz7sjX+UlQTN5t6LiTBCfzTDpqA9wOTrYZenZGM2UxAbwqfBO6rZOoDjurp/s0sRH9C9G4d/rw
Y3RJc86X1ifDww6iyHdedIOua5bwd8mgQdHhdtACrLMl6PxFcK3O0jH4vLD1bH7xLFz/AfB1Xhha
SKu+5zDNXNdaVnTiZzVeMGdLbHSf/JoJ+c2d7B80HBEyCPLv+JwMVKjbQPde3fcu07hRP++Vjt/6
PcCAdNCB9xv3YgFHP9LwcQNJ/AQlXtRRiwnl8owF0P2Pf2SdkP4tT+JQ30eWr6GvDMmHwMcrP8cf
rIcLw1cbvgXlXmRM69Y9GqaBCSz1VQzQOAyBGCqUDHSaZE/1PVG4ezw+YUSTnmTMAZIDjJY4m52w
09hRip5+HZe8b4r5y/dXIEAphrVdsxNnuEHmpyY0HtEqXDx2c0uYwwupG1NlGUtBWQHZhwOxywa9
uKvrDH5rKgh4vqhhM06NSYo0uFP4qBDLNnlEtOM5ABhG/MtIzKDLsEUg3TWm1tSuZYr9oFGaJCYY
Ilx7m/9b43Fw874hwlCqUd2CqRnjDUy6jXbLMx0gSfD1x6bThNwfCjWrlbuHBp0yY+CoRMLwkPOc
g3s5qKJZsdlMby2Xp8ZFY2MiyQZI0LBGhkMuU/Y8Fc71lx0bptKs1fNpVdmnkwZ3zEI4lYrIov9D
xiz0z1CUFIdSQmuoQcTlpikkW9rhnI1yWlLIV5JYUtsbqSV1hBaDdN5sa92BiaRseshg3Q97a4IJ
RMg/8BLX7mun1+JpcV5MfU5aTUp/PnPJ0MnposC/E42iYjHDoBfwRhlWTchmyPpa4mzZMg0nBU7k
+11+U+oAJ/vxK53/fCiPC47EsRTVZOEe4IMCXPElbIYIr4Sd4DFITrcyl0E6qT8vPnXoVnssIdU9
rsqHTzUcR2iFvakGh/n6mHLOdGmLLRDZi7T/vouAcUxs3DI31YqoKCYBQOLHUa3SQYLKyu69Pinm
tLLqfBXDeIANlgSuLGu4rULlB5xPpJWfwDwi/+nmc1o5GrGYmUdlAtEQxVTF/UQncMD0RIGc4tTD
FR5j0u8wpIKm6A5wgAconC86gVeQknIJNwgKCYVLnrD8/IJ1ijzCrwZgh8g3PxrN7dyIAkr58Ikc
41GCyx/TFKF+mGwoQB5kt03pn66KT/7R1FsIUwmfoxTLxi1ThhvSHgMmXoFmO1oIF/fIV5bA+YMJ
zFcflbL398bPteCzs8olAFUZE1v3mHIkURdzqrlsJjUFI3hhU8db6RraMcaX2zLjvKMtVy8nwbWj
QdMj9mIb6V5RDnC7RbyWGr8Q5Cgbr0GFBwo4DZM8u7aMMd3ClXj+KiKwTMGoeYAantYOLuGrzgP8
lwDoHIZtvAokHq6BnhanhLNP3ibB9hjz58icVwHqtyGC2W4V68F5slJuZBmgKfUG8xm2iecEtxNb
zAWTWhnMbBs+IirwtwQ2EvUGNFp33kMqkw2mMKgX7obR1py1Yi4ZOu+Wvv99aT/LdzzkExAmWu40
dtxX5irGKnVzTez8w0XGe/92Yr/v3n7YISZXw8lyNR+u152FrIxplQBxC0sT7ynGiHYO1vLvJ36b
Mb3SDoH75QuCs0dhK94wl6C2NQnyQfegoZoWm5RexprWsBaiDLHMIFK22Sjj6Pgpe6/edbGN/wSK
JvToj3VHTY3iXD+dAjC320x4OE6bw+zPibES6TPoEl8i/CayRVU/KjS6k0pfSyFFVjfwh/ZbbmRW
wubVbNJN3VeCCZDfOplyclGwQ/dt1z8xVn1GrxYZ9qn2FyM4ZLx2D11lXsyf1MHdy7Egp/gcdb9g
nYUWnCw3el17HqMhB+wOGevlfo9nnTBtygbJyqGW016dw+4PzOgXnvzGsZ8fdoZNiAU9hNy+K0ea
EH2OfhJ1dotTyL6QNnfUkfBjF5KIsbprXDFI5lZK4fQ57FFj79liwrEa1eGVH9Hs1S6FJKaxIs/d
r0I1em3+fyf1lstb+O9TEt9wZBcgsdshsDIjSIvpS1ZDssh7LkF7y8ROl/4/25UeDGPIs/bA/14t
mGqQGffa/rHcL85BxJJwBT9tltdpLguYA3++JEDD7r8XaWJWnxpjSzfKhzipiPYnyfRSPOJ62noU
45Pbdifxq8nQn24oGHBCPsM0oh6Oez0SQ86nNptAxaa4Wx4MXuD047im3PRqnpmo8AYVmPMjiQhl
N+hcy0eP9+zoyhTaaD6nPoqSq6mqebNUoyl4xlhUcyHTe1yAGNhwHwyJszoAmUElF8zO028kuzaK
dZjo25tiANmKlpf27ULTVGbdTJHGVewfJLoVBotOAMczIYrvQqaWSncnZ+6ic7Sps/NiNZi0ILwP
fbF625S3/CEKcs9Gd0UPju8S1UyretHzxHKSNocIWkOMz2Owc3bRT9iLtXwTONHxh10YqqK9+9GF
mBN+vnnHWmIZpH6GLfpJqwJFUKkfaVlOPQj2uHwlX6Ekj9Tl7O6XPNg1pnEH9LmCEI0K16AZQikQ
F36jvctlRJ1uOntgojdJXQSWhxi/rEtGgRGgSYc7jPFYOH4Q7ysHIpfBqT/V1rcDUA+vKumFfxo8
5WOm6Xrh861NlbfWUppHPUtsDJFKj56ydaKRRONMMhjpQGHUWQ66Cyv5CaIaXZxAyyf/JlegzZBM
dkH9nj8nGO4QObK/gTDMfE8bPcsorAbNu43XklYWkAQrpxoT5ey0RKT1rQXlvmZfQyUk19otRU/B
tHjcsNGxXeM9+LLSEwe3SimeT6Pkmec6Pi8lfjCYF4N6Qm+IlRDxEOtUnb0H2WmiY2nSqQ0eSYPw
h9jryynVvntamyrERROQ6YhjHL8wiRruX5toTsJ6hSfPkDqJaFDR+5/ANmxb1rvmUXRRLRaBFe1/
DKAK4kaK1/kU4pnL/mY2Z3Ak6C9V2uglVEHj+Gad5gKrQ9mSoXsqS/nEJLXHnJPt/f+U+Jtqpyiz
SL0UlwMPAjGCfgotN2BWelcxrcZWQEQfGCVdws8FW8KJUoIB3ZZN/Pyib43uJwpX8jDuN77ESRlK
gP7VDF3nXFYwKp1ZTrHfuK32uWUUNbvJa+SLaHcBOoIem4AgC3M36zAUXudgpxozEi6XnNJHfR9M
Mejb4Gz/IodJZHGSv9ORiW/Rl27k4HImoWj1LwZGnxNonSyGHZAZobNZ8tQjl7sgSdaoW0mooMnu
r4MVXAKav1xdI3EcKpmwJ/2qQ+8XBV+uPoqYxnmwYpuic93qtDjT6q1Vl0k+8WEbzztHH3j2TsnB
UZv0jeSFGDGQv29jHknVG+ERGzfgy2tSu/iRg0bzIvpQsKQW/KIymMcGuaCNATyznvYF/CQ4x0Rm
ix296B0XSt8WTfWndE4OWY0xnVxWGLxDJxwsfLGn4TD3WIOXCFEIcN5z3HgrBlNQTUkQ+8XRu1YO
sJHXrDNeAbMC2CkjU1lm30B25gvCcneqIgsrqf3+q88gcg0ne/s1ZtOIYTcmlndUjPc0r2+iglMm
9mmNBupZa538vX5bR3PPsQ9UMi6lDBGb8CzP6IFWOFtvs6Y0509IxI7z0n+Jg3uVFpt7RjfO0RkJ
bP99J7RoQ3h2OrEojZ/tbiwVX9zO5AmxerkoITjnwQKmb9nR+WQspCLFPeXz3730DdEfzeLGai5D
m0Q+gzqBfNZPlDt4zUP8/dc1sWpGwWtOtowda+0K1UIVa13Ory3V3RuEU/fXdm/92jc+Sjs4hA40
a8DPFY//smJrcoE2fTJ9ZW17UeUEREjGn0nMepkRpG67OGCG+h9q/h/MN3cMVARZaDG1vWIYDOZE
SVhLUoXzyt0g9PMwukiqqmGpujc/xfxj1lyOt1BNyC4TqdO903HmM3phjxyDwAe4Pf28AXNzM/Z0
LkwMBbDmWV9FZxUrGMnZQ3Rlufx+svxtLv9S7hkllzdaGBwALt8bizp180PCrI3Jnrx3d3ZNrMtc
+5LpreUaDS8SY5D0oVlt3RnQnF/BxJoKBOyVamCMRPQhNP93EioNtKn9s2NNLa0rt6fWh1BbJSbc
DgIAGVEBen+FRK09Kiy42KujH6TmrqONyxYAGABb0gC+Bj6dntSIM/GMQSalN/7pbekmlG0/9v12
+Zmty6sWEfB27jb5LHj5dKfx8IBWNmYF9xF0B70GuFLElEkhlqGRKHZRrCJH6Z882axuN+hUGAwr
94Jpwx7ITUJrTmB1yn2D1K0rea/zavP9xfKZ1mMGDn7MbWMwDv/YpqmT0iF7mQN8ATVa85ZPoi2r
zVM2PGX3emHbtbaCbwKHJZ6dbgri103R0xO0WvZpVhU+DPr86S2cnBM9ytX9aiHBMeHn5QK5iL7r
YZdSY44Aio3qO4ESQAG8WDo00jbdCBlYKYM28DL0NXPIZVBc31wG0lGtKH7jmgLOrjRm6Tof+X7K
ScMbZ3Xc/U6Nu144b/sRxkiMmvdLOYZWUZrgyBriL6KmRnCIAx1+m6YeSfp2bAyl709TG7jObPOZ
/5Q4x+HwCcpOhFlQ8yRf+dxqcEliuu9OMwEUyCqUin9mAUZZctMet1kOj5hlpx8YE7bOJAstZmku
ITLT7GMDOaA1InV72kDdQH4jY8GI8zToMcAo8z0EI9PGt4ss7A7FxltBTb8JaQ3lB2cVHby8aquR
4RD3RrVECfR6UZR6mJcKwvTfQatp+kNFEx5xpnwW9200hfFQn0pb7xoIAhXvffmTM0HClYihIbP7
DcvxoGm6dKp1pFkw1JPRON0K5P63WVbq6NQIq0nlMN3HEnhP9anjmqGM0vwVwD5WKu9lP+JHXr/R
bpiM+fd+p4bKW5DRYh1EYTRwHc8mzHQ2JPuAim8wIZx5VpJYXpZ0mL1ZEVCM0GZuEy/7BYBiUKqY
gcg6BUh6aU/7CvncVIUtrPtZ6LwdLDEdY+UdLf1SF1x+/jMk51mC/NJu6WnkeGWUZnqn0QGNpve0
QoQn7YmnleeKwfRQoiQ/+wlmX2QyQVvr0h3EcDQf/83CxS2k8xg/hvHaqi+yWMVKedMqCtZ8DUZJ
dzC8DxP0QXpaOo0iG3Wqmq2z8HStvczoPvOj8W14QH03PjNyLr3zrCQZ+6AFe+Nikm2WTNbmfBP/
on2NoEin0fzTJy0wF7UQq8Fi4VGvf3p3ajrqNkERMXK71gsOn89BseIpk3PZpzDId5OnHewt6O+N
xgycbG5em2ulIIv+I05+Szug77P603FnpKqGKfORxvXcZuILz/Ry7IE7MepSFLciFRct3Gtv0+yr
mGJB3Y79lNZz5CoAPLfsxLwNxJV9f87Z+vacKSD3AnneXSZ7xMDeLY/wFzr/hi/aLf1flc91wsIY
c/1X/x96+6ZgM3fQ3V9IfbRSNQJD/AH1pMMN8tSckC4kakeYelnybwyUYh6OrWZ2j3pkPBCTxI6r
6GjZhS0G6SW8gNfzLfj9p6rbSHYBWQK3NPZ72taX48w6UoUzDJPSCHw8w0W7kYCBLJse73Qm74da
GFLZoWinnu68ksBxMVAwUaQbJ8esxvjgQK0+FXTgmsIZ6EJRBm6Cf5FnWpNy3kYxWei7yq5IFcxa
Z84NM5TcD31LZKBM+936THDYD5oR6qLelvVLSIMJo6GPlDWCubD6YC1UiUavl7dTcs1DrqVqmAqU
XZvBlHo0/i3O9JNSYGp2zwerv69VEG/ZZlHe+pn2EoCFyxs+B7bnlfLzLohlp8F1bfI74v5XYrNl
GMY8wFtRHwldEotLS+x3phw4oR6kloR40muomtIJz3wEw8PXwk9NsH7ZAf0MQrIKDQpm/pbUGUfv
WNFQU44NDZjMUpjPDyx7qDaSXmuDDnzxJzM9WFxjUYkdbtpjXE2Eh4OMt2EfcjC+deK9ax8QXKXE
z/Inzly/y2UbjxHvuIDf8BtDkrx6xjil7KJm5wkBNQZ7whRlwgHRVtyW8EKI0ToJaP3Kmdusz33Q
weMcOtWHXi/0+UC0yvSeWNoZ1OEx0kks/QTdoCA6VuyTAr01TuhihPAhFQdmBYegoJ7hHaMtCOxP
JIV3C7yNTwL2OxpYl3tY+ETmH0iEh6O2Op8JeguqoxMVj6+pxVkar9yr8BLhyn7S6/oWuja87Z/1
umraZg0OSxZpXFq+WpJdmzKQGUDiuqnxEnVPpUbksV3hgMlBOf71pieuTDghTWhTrUkgWVPu0w8M
WLFKlGhzcuLeEqKektcE6rK//bpQm6NKS0gNfig5CGW39Mg05CqfgUsTLOBBCKoAFUdcaN6fv9UY
tQGJ8qXaZnaZ2s71YEEfkp4mxnty/bKgbOgd4oflUSgkHBflRUXX0uMuDbLyFDnVdDuLpT4V8zwE
H+4/tg0NfkML77OYuHN0of20z/8OK35yHtUle3TQ6YehJgX8pt0rSOuvO0stnJHD7WAkRWLa5jPL
9x4Cu1Fl9Zhtr8N8Tayi3/OIs1mHOa2xD9JHACKGPmInK8T9zvPdzvh5w0nBH6vxskoGg4BNFzaM
we5a8g8H4PHni9vqNLf4T+UBStnHqkftaiWwmjdWxMCpt72Y/hAulbDIHnY0dvsGmwBQngW79i87
zZRBwYH3Lu1HVepScgegru1EgX2vslen5VVIQ8yG2yKi0DhLy4+4yQMOZ+YnaWCrxxRh/BU1RxuX
63+Gv2HR0yBQX2Kdu+WklEVTNvGi/BOmAPauKG1w76N2xw7qkDDmsKB310m8qXRmUOt1DLDUrVa1
BmoZdorD7yzecLwRzNz8f5+R/7pjXYWzZy3rEJ+i89pAtVC2OBbwBxP3KlE55ppmWckwUcS57xQo
yUJymFmwkQB54bbF1diswb1PURGFgtJGlSXa0p3RlewMdACuE8JyfSb1FPSnBKncUX/SNpr7woUH
4O5r2Oi1mKlSKTM0B1HCNjCaf4Re4rkUfcD7yY+jk/G51BHx0gTVAMCoylzuzDCjOrSJJ1oHX2+S
apWNo9+Lw8jC/rebEdg+EfIi74XbZNlvV+9MVivmDusWOUz379GmLdQ1O7b7Kpdkyk0yiHIyvZnB
psoWlU+kPLILiW3f2zEVu0lpqqVapNHwqg+YiVwj85eNtv3VQKqhyiEOdplCGdJFjKEMGGPAhF5U
o/LBw/SSPQKrR70+iHlm7DMW1XHR++5NsztfLhk1IvM3YfVJkpDBnVnixBjbbjcpE2jd6D0x+pSj
ZC2RQFZ+C4KjZUSaYLs9FK1B0b4emaJOEqu/wsiC+Pf0E9ifjRzTEM9fXBA2tRbJyTCLflc/RsZQ
CugY+Kffb++G+EAbsmMuO7e+KAKYnwYHqqwfWwEBO4IKcpOaD6RsLVpBtdtGoYEFU9ir6pdvt1BW
ndpAdCJAD1qLpVu7Vy8GWCvhPrZOFKixNYfgsj5ZxTdnNK6eyCuHEhabSOxynvCeedLpSQ4nbWP1
HkkJU5FsI4d5MOiAFw/YLVFlrz08KVN0R7FERlNdvf1INfrIuhFQMbDuaaxSQBHvW92awc/1GJt1
aGS+v8m2AYsbOJPO+xUeGII/EFwvJtGv87wAONtqBJuXWem6AtE+Zds+a4KwLXp9fF3r/m+ip0wJ
bZrCwkAAaAd4T+Zc/k0j32TH7Ff914oGT/zcFKf2yGXZyRwgMYdIqwNF8lSvmoToFXmklK4EreHO
CwH/kLN7x6rubzsyLneRRjHjgHPjMn9TpXLy9gI/ZOHzelwywFQ4WVr1yTVor2gf1GILkKEPFDT+
hVQUfU/s0JcCWY9F1LhiJBrf3bwfiPBEoH8P6U66RIgtLAZQPlU2PSK/YeZrSPBI9mKA7tsy9q7a
1/1JFcTU5Qaa3hWZzs73ndcC+RdFobIOg5zBgBMJint9YvYgMPap8ZSLZiLzGr5DBzRgA83zPP4b
lJvv38h9bOnvenAbQhbD9siIP48FX5jARzyMcyDGFXwh8Joci43KbyIWFXeOFAAYxonYPwxD4/1s
hhYsL8CbZF6NBilNdAZ4nkPB98EDhYuPnYCmZiMdI9eo6aY+Peif6zWO2R/H5WJcYzNx7pc6UEYt
dtaAnxRJzDP3LXT/GhS8NEDbsOW3a6+GZFF0KPGOQclbCUjFgGaIQNNxTaBSAu9CHHsk6AZUkagu
y1AlvDmEXso3sJ8j6TpAl9IAOQwuaobDi3oefzFWwTkc0JZQfqx/cLTyQLVRQoH+OAWt9tudTxGl
Dfbc75aaS2N/ZmIWygIc/XMyMRHPz8RmMRrPaEJ3jZl0wcfS5HLzJJXpfFnQbqKGI31m6qy38Crx
FaV4P6a2tuqdrViDW+85wF+LnQzIEq2BFisOcAAC02NUhWS1BiL9nvrqkVWTTBfsjtFlI2EYKjOE
4Tv+h9B1zfQtDeAi6pGdwsZUcuc2imqL+TkjXuS7BFpE9J3AY5adB0NG1GmObrWTwhsPHCuX71Dy
/Z1zkigjYH6ufT0coYGkdtD7ySh95OuTi7/8C+xyYAei4/H/gK/eCDBO0jSU1z7+7LTTEQnNN0of
1hEFz3en5hS5OlL+99bf4myqneissNOGSvlYMHmMGqlkt8gs72U6mEYsKuJncdrPRVD2ZIx4ipXs
DX2o+TqaH/uTUiFPiTLtqEkCjFD6ajJQOQSiY8UVXfz1CMWmPtqsqBkdVbhDkYCWveUOf68AQJ4K
s6Bi2hYy9ggjeNfasTfenidNVa6wDuoalgk/K5EvypdiSQf+iyYcdqxtnNkQrA+9E+ZV3kp8bx0B
MV2kdKWQoFFWf+BcaXNJOek1IZF85gN86KDkOvg52DdI9IEJKJkq24dOkpuKn2Y9T/bLVDc/tfAb
HgrxkSuM4/xMJLjpWoa8AKJFsiIVMGZdCHuriMCH+FzWyTtrMX4UMSDJ+wWmmn8MwR519brQMiPm
c2CM51Uv/U4wr0kHWWgvJ+pl1Y2a+yd2BivgUFFq7DVaf/2hQWNibYcLd4t8VJtflOA+BpU5n8a5
JIPf318BaZA/LEVgYrSDX9x5tRtWd4Lz6eeh4If5C5rbHrw6TqTqa/RbZdASs0rY7UZo2B1YewsZ
s+rwDoabU4HYtJh1e6ojA7JTH4IikjPfTN6qN1si1UdmOVsHd1gHvAXrsoTX8CF9XoBeAXFEJZt9
FJbHOHBG/cYXH+5kTZvqhr0sJ4UHf+JdjfFggZgGGtlKIPsl5Qa97yOh1UBnPxTLbfimvjuUHI/G
4BhSZkNvzNSqm3HVYns84i/kZw9/GBRJqo8o9xuOWpmhmqnvoycoX2SQJ65HQ449/rZaxsyA0Fkc
MOrHkz51qXNsJzvOYCaIOaRozmEUkVMUIvGC+t0sgXzLAeFhmUidQAD6vGYFPTWfzCz/BWwewD54
DwSz9HzH9KJ28oi99NfcszTtVPVRLd1XlQTu+gBprThEysJProwa6sGdKFYZKUX0kIcXDdKXv1Zk
+LG/Cg4Gd5pXbfemRsSbNJ69+sdkzbKCZJD2kfSW2gKiXXJNGwYVqh3HGtUkoRDoUJHZyzpbjiGX
8HAwm9ZHoToDjVpwJnZLnSdyfZ752oiHdpesNJ8N5jtC6zjYEmEVvpaT+47poUfy8hjSCyh0NYER
uDPs8FGVCj0q5SCXyDfaBSfSzR+jVvLE8XatHBHXDviz5NGa4hpI6crcjEihoj/yKc2dD0uJXEFf
HoXQCGLFJjUNLd5guwpoXxUiKfGqK+6KV8wE3JxNhOr7ifMHZQFcdIVwRia7nH/ceY0gv/WGImzP
kjIk7XHrA3i7Avxpawet0YBBxuRBjYPBj4/vFJzJLWUMK3HkYgp8TQ9NTel/R7wBV+iSIjNRLvBQ
w0Lu4acKIQ6vcNfTq0bKRiAFEkuqNl8Q7gO3dKZZEdWrKo2KyqcQSOsQ0YO1l9MSWgnAKkZVN2gE
qEVRZoCfkyDtJzCdQBk+BfPchlgKCvvyEwrG7PCHqUhjnNcBhoeM+UMSsDAusPM+yCZfuKxRTpaE
bT42HXMFMI5hVsf82vgcz9OW0r8FyfjwZqBqv/5IoClPZ7XtEh327O9e2UvOfMcfaGOJ1IoHLsru
Y6H79Ox8VtDObJHTTS9wZVnsx4ifPw2CU5LNqAbQ5xOgnvPB5T9LYVGCOrMWb3UCUqOIBBC2YSRj
RTnvedDfEwzxhuTnWA5OgSW6Y5IoKyUDRUnHZ1pmV3R2SLYBFmdil0DIPIZ3K+zyOeogAdVpy6om
cTpTXv4wUjDiGQHnRVXWaQ4E8U6WYoyXSzDruNG0gGEHQSNK0siYKq2I7qP/5Pwm7va9Ya6T1mFg
JFPXCoT5nL22QZCdkHUdsg22XPmYJ5H1ZlC6hhiIFGrnJGC2Eswg6Xn/6GqhrbRQPaKW3/ZH9nKI
T+IucRlV2+N1jQTKVbXl/xOVC1TnAJCrdo8xbOfk2Ce5bpcYmfSUBkjFLz04Gb9hQAV+DynUDKn2
cOAYySZyeAUbke4SH0WgFVgqYu3WHort+9DA4z0hlPXiughrsV6RoLwJlw0ekddzyXJq4tg5KRk2
8Emyvp6E8GwUgm9DLbPZ4EmGmMFWH1nEUwBeD9kq0ufxMp5TZn1M3sOQ2RHwiBiTT9GPRdvR398t
y+P2NmlxEVWeioMO9OKMAGz/YiMbJU/MpQP+MDb7buvqwvKtponREw3A9afKJiBN8V3j4EYGMeeP
bThKPBM9ExmqAxgpk55zrQ6+W2Eohq24A48aiHW8QjSan2AWB/O5NzeffYkYcYd3uO60oAdYLDZF
P8+N44nNybAaOiox93/pEu030+whjOP8zpTtZD9R2ny4mjLSctj3jt5sQVbL5x2zt3SxlVQ7S+ZI
oYJeVBDTB2en9inu25c/6azKftsTqPgyaRAjtc/1bhNz2UKZWoYe6kPIa2JDaOBseiQ/FYo5vf2Q
su0bJodYcKx1mPfgyeJcgUyUi9E7HFALmZmhdLOnZN3ZrJOz+mYcW7Xd1iFC0WdHKKz3IUVdkHVy
KhMx6PTHSJkIr2V+MCK+n5uXrwIxXJWgKYvuA9fTQdLTYg5xOYiVDqgGTWNuBXc6YlP6G92Vp7UR
9DtnQsI84Ye3KCD3N+FQ7jeVoXntVJTyeLhRaAJNDUY3ryGP41HyGbqaTu/yK8kFr/G1M6axruqX
8QPI+zltYcxEimRJa5vXUrU50/VDg9Xqz57s7QRcHHG2iyiqZmIDfQeKr6pnf7tIgBs4EUvjPPKH
JI/8GW1GM8qB2dIzt+80i2ZUxS9UIKVKwXVd3bgthLlPJdYzcvwUkN2gYeU8Btsmo9XbPXEfkCSt
GYi5kAnId19aEl9z9RTnVxivD6ZRCQ6DAcWxGVWdlzUOrnh84SsukkPQBanXsjtmgElalpcT3Q2m
h/di0vO3RiYMlhiGwwOsQXoRd1LZjGWUiOW+b6Wd4Np+1SccER/Vyp4/w8+4NeIAZr6rX6kkPZ8v
3cSmhhaNPQzzlqtKKGYVJJ6uhg7FlD0H4MqYWWMiJ+9pVdE26ElXd/qQRATl+EQCnsILSQIwdxvJ
go7Yh0JqU67mQ0oLAjYUHXMym18jruGVyQEX1AjSbI3uylzvCcQZUa/nNiRfx8FYX6F7EbjMUAzS
wuheVGmDvB9pjWVhyoAAqUC+C1sOWR2vidoVZwmchAG5nqbRryzgIdQD/BnEFlGbxzKaeLSYZSwE
Yi6XzFfLtPr9U3A/60RiiAm5bwZq6O8ev6AQ2alEKFdiyXiutAWmZHAyal9Cwtje/hg8/uLG/JzL
uDIJ35TjdOUhRGKxNztnhMuigYq6iWMLiUxO/yZhlPx/sJMH64Gi+iBY4dCtYkSpkX62h/7hmzys
wl2fd9deWDh74PF/f5fpVUoIl0GL0A4Q6z0a9DdHmeFaXU4j0HCJG2QI30gPEX3RelqiCXLgDDO/
wsdPILbu+yONULBZ9+a9t1Gx9WKm0vP+OfUtpDUyLUQZNIecBiXrH4YPOywC2u53zR1GGH1a/om0
T9t/dnQA1IsNk0vUzVoUHKckEz+giitzVhqM85jQJtj1e0UuCRyxAEg7KdDlnGKqapiiITDFya0z
nWa9cJzpb9JQdisYbG7esIrJ86pMNJ4KrDcTMtfzFPA7ilvF56oUSK9V9VllaSt4DOAIYCRE2+D3
U0PykzZwqcXyrlCThzhbJ4cFrL3/zIlRV1bHYj7XXlQXOXdseOm23ZTLp7LT1L+/6VmWdQVt8jDt
UR5YkZYAeGVIg+IcyZ/wnq+xgbDAKfZx1Uh3/W/3XtJLfkPAHxW7mEpUfv9NUTP72YZ2S2CK2SEn
GYeBzLiX4zF/9RWoodKhcFDOaxMQsZ8plOzGqZOVMcTt9Y032PS8fZWU1vgamSbCGG83aW1WMzbV
pMNAb7GlhUAx+TIe/lrRHlHGXgKX/1kWFiFxXqS1X6x0Atkv6gjZX2zLhPDv0i49NJ9bR7eU4/WR
N7VEpiwNvcbUJwCIYa4UlYBFSvme5HAiCl2PKPkNgGH8rbw8PtLKy3sMwf6NrN1ChXvymmFNzYgQ
0JyyIDwwMtUXoSWTswDEwpAVEaVWWL70w56LL3dPzXWvZuPhH2elxFGj8G6QbmioT6RNYmmKx+vt
cYheVBozfRx7Vh6ysKGI8Mb1P+QpNKbxsfWPfGVnaoa0YDy4MmK1uGOBKACppJQowtzD6A9Z2Dcc
pALctrLAQvucFeJS9JhzLLjt1b+X8Yvn1dJdOBFgzSzN+LL6UEo2JjZbSifyHqqTbp6arr49FBGN
umehNa9++XFV5dmE8aKVp6EejbiuXo+/vnqWfeYoxRiSfkwdoybgJIYmSdUeOtroA4RCX63an6Vu
iINnNAwRP4DJ6jJIYHsAvc63AsD5Gp2kQ6uEPVWvUvQ3EujpT+5iBZwmuMw2Ct/ADm7FvQpGnQIn
O2Gqg0092JoPm/Quu8TsrnK2cFMuezurB55q/SjkNLUcc9wCuTmquPFjtn/fLLTGji7SIuulpZAo
R+252BzPIO7rU9RFHCajWF6y/9zT5ZFWMRdBKzjidBgzgugV/23zQNSeY1sUfHUGGAixHZEuzC/s
/Xmv9ItNoztJaILAoLraRulM+NgUTHfPYHnmTz4AgGJMW2lyCcnnY7DaG5R93hjc7uPBpM74DduQ
MegKoIarTPb0GMxjZfpxFKPIHFPoZLXz96q4Rgd8G09kGqmfhhUjukLYsf/4+5v9TPKUFCBFuWu6
ccmLMEhsw9cQCOTshKRRf3EeEQDNoy7yAdZPtHdmePcoLG3QvleOhkpTZopZbkp/mmIKMMTkBJGu
rEpOnkgdvHdTbN8GwETRuagAsDehIKuGcrJBTArhOfwwkHnJhE08GtgRmj+PlWgJwBh5wRS9ck3S
gE/QRjUO96dX7k2CGBiW1HHCoR2EInV0IX/6/qyaSPDDuMhLSbsaXsUfDt4c9TOnDbYko3e/MKCx
o5UIj3GNyg2huz8ycSW2x/Vu7HOs6558I/WUFtkspzAHEqVIVjy/4rBCPmSXPSHCJrONkZZW4cgE
fndwY3f+Rs41Sfc2mJ6SFL54Wlikc8j9RQWuEvQGJHQVQvPeHxIdLmR0SbrJxFl1LPiCLneZ1yGc
mt4vCpFbHzoRG4/Hg+wxiqtM7aDr+kPtttuzoanB4XglfuKT5hmMvF5F/FrEoq2OCf+LK+Bqacma
szWZuRQDnM5A7ad0YRXDFPqdv6k0l/NaGb88uxYJu21aRdDWTuSaVSVK7Qw+TIxF041gATTjhWYr
hNCoo8We6ZlqrZGWi/8dR9PAVctrW/HCh2Hn/znWBWlI8kxZZuDDrsgS3XAQMTLH/bAtGYZ1niEd
/BeU5izcdaI9SwQS7RDJDAgPROa07tUNMPFcdFSElBUYuDGSI18WVsETjDVoGP1+u1gIkmMfE5dp
fPvi67brcTrS42RXrDFcpceS2T0Fw3LfItY2F3WCjWwvx+osQubRR69ZAV+O++sEmqzG9E6Z9ZvO
jzMoycbfAVsImJTS//sqc6mHyI9ZGpnb8ILMpoLFsgmR2R97bRNJ6M4hCU6Zpak+CzpyTm18rejo
c4+5eYGUIbqXHbvI1YxAGF9ZJbIfSK4wNfzKLgZK5IPeBelCvxiD/vq8KkSfNvguT4KaqQJhwdTl
36WbZjILVXvYLgQwyq9/NuCI7W1IvAIuRtxrmeoF+aNL53sIoOeekxjMPowSIsQ0I0SBZGLh6blA
17N/I1URsyi+UuSMQo6UHHXlFkTomuKlNkDcQzVN5S75ejLF7MGHLBX/+2B9a5nmPNBBe4y53Vmb
DwKMBPOXKaIlVHsUJJYQlbDRJWM4N4G9fv33rMzNvrkt/JaKFsQNDVy7vHvQ6m1jdDOT4+AfKOxp
gIut9XfPTVH2k7zNTwd+9mbAp1thdf1b+9RfKjbYfY7R5Qz+sWby5gQ1Qb1k6Rj3fmYEYjguNRpT
GjK/T1GMD1jIq5zjj1fEn3KpdOOAzE4sYA815h4yQ9cTiFb1rXjberH0rkU2oDRn7NQQOW9+DOMN
Tx311JrKUS67lx4HObADr66me8HKLmcK5AGNrBfTINx8Sb3V/EfGp+mwnDhbsAbJBGhOXpmldSaP
8aMkagBVPtUANDEdEBkhcfGt5tqtN2/XJO7u1sO0tkl7KJjErlZgbf7mb/rlyk0w+7NHrqmetyml
tFfxuCSc7+a7u51tUwSFswod9Vv7Q83Cgjp2WkHFH9sNRBjqYp9WE+WuUZIU5AJQYxUOSuD4kIqi
geV+CEmoZSB2cHFId8VYq31zy/cs3+xZObf/Z53UXNLXVUWfrf+YaXSnoN1QzM31slx4g8hfTTFf
WyIgXdpPgjoHkqOxhmrBcoXn0jyilciXYaDVvhtUbSeex/zlQn0z4wJc8qr0mt+BFL3e1nlXa20r
JJ5KotX2UeEYIPnGtIDTG4z+dF2UBbvjzGoRNYkwnPQitiv4Beu2ppk3vHd9oyzuXqQ4DoU6Nt1F
3t5ykUGnMOuNnJxwcB+Q1zsdBVdHVUHC+IsWc3VpQ8HYZ4MIEItfJk9DMktrOndmo7g/ouH1EbF2
7s7BKMkRSZWCep6va0fs0AQ8KmM8xmxqd5MjeRpPWbMX/9UVE1PA4jo2pWl9Q+SY5G4w9E8oq/C5
JP8QKlhvdwZ+7LOOZBMfxW7qb+6l6LpAGgZT0nsUA/GRMnQZaM/vT5S5oRYesBZf2XiFlwHS2cht
IhDZ5x2wNoPB1Esfzf6otcJco8dnhDgEM40vRFPjvZBsRCXDttbjxwlBtnf3ITIlAIUpVVnqCY8I
kFKQ1Qon76keVmfcAtFSKIOIBUE86gqzU2mAOSSjLjr59YaDq2rV0C+P5zjiQFZ3L4aLVwXFBfWN
Z+tzvbwan607Aably61BYGfeaahilE6bYv8RwEG8VqTiZNZnk+imVR/TFbbCxhEgy/n28AvVi/KY
wmdLGQw4ptKcU82yCjm2q8tPBSnqpNNYBD4K7p55JmYt8FYg/9Bn0DpizEmCzkJlOTxsQLaOhHs7
4aHUDnt15exuao/9PekA5oYgPLi+Z636+ywESFrNKsB3YH7MS89VAjt71VorRB+H+vJTOx+CN/6R
jXPvKIFh26UVkHHfTGIfV+bki5T+DQodU097NAnGkssYkwUyacUqEWiNcoG1FXnU7AsYael9zWjh
YRmjg2MBEI1BJ7xk6VWXg92z4Et6Ekja9vJN9dDlUyreL75oXTGlkGiZII6RWrGxb4zahtvjWw79
9ZiMPX+//K3YsYpEPGQOPqeEWCE/KCG9/I6qDuPSc15BsAiH1FdzY64+T9mNxluTwox2PhhUU63H
YExHombtku8JAtCOK4cFnNmsD1oG55cK+CGt29ZakPhy6/Ghe3r6qs4gFtElkEfW+6Jz0e1pDuYO
e/xaXiri2aTyegBee9ssV0L89jBM3RxRFq8qnNgkRpT4AHgGqToEyrFQaJasEoMi3Cu4StUBqe6I
n3J9Vq5jPYx0c860clp/95hAfA5v8QxTXM5g2wXKZQGtM0EG2oeJewEQCDy2pS7xnt+XrM2o1l6w
idzJz2D1QjHlup0KiwXHpPYXZlCbb+svo9+vFhaEZKQrbwei71HjCt2iVJLEc1dZsmeoODLmqIIG
22b96whFXGWR20WJJj6bJBax2eV6KgDIxTvtRB7QKfvbkemaW2Q1CGXFgpjy4Ad7kMZOs/5LGkV7
SfowQuas+burMUVhWhQcwm5F7OCDnAVMHkw2Fur8lk1XKwA45bubef2y0V/ikknhxbBiJ8YBYru3
o9dyVO+Da3fsJ8eHymif7/PDPFVvSCsVaV1/ZhdwEe/mLnPFdpn9u0kN8jivQ+r3igwOgFHPgHg9
U4iy/d+eT0QrIqs3MxGi4uHiDA+r9qSCzadFjuZ7s4nukw/6UdD7zsd+z19zT9+H48l/b3g5oDrc
AyngWdbxhhGeRoTl4ku/uAnY9RmKOPC0wNb6IG/jxkajlKimfZ0Zb5mvF/PSAA2y0zdv1vIsLIKj
T58CXVPcskIgB1VvlJhmsFidbpmsYAGHblKpxhBQqMqmgFuaKc2Vb+aNu9yMuBHe6ejQ43Mq2w4+
h8OrJUNqYPiL6fGfV0bXia2zIL86gw3d8MagrpAoKWMBXM8pyoDbWPHcVs6JgIfk5SV1SA+eU6ht
8ssaC9dr1o+1H+Pz4dRtOAW8Hbu7xtDNAny6Ovkq7/oHW9mXXPm8xRhqeHiS/QrLzDqTd2FzLZuz
7FjKcN172xwwzo2tkvgZ5xXMFOziYaVVSy8tklqJuvSHyczhivvwKTK4IzsixaEKS33PQDdVglJ+
Qls42Lo25evx1eAsFqmFleHm2qeqJWwontRlUZZw0BhthMUg2/TrE7O4e9laUpxwodBY9GdxDlhB
9GXkpOIa1kO6aOAMGP3nXZnRlSNWY0wfcXSddrSS36TzK0gX3KcbnI6xzuCYISNzBFeexXg9DwOp
ZobX+mvOAZlCprBq/vQ7HGommf5ZBDmxDz4xsKCKNV+xYqvFDiKa0JbSjBH9Cyf+mZJWTogbRXwD
Zs4i3mE5qiI7KZqMEetJGO3WMbenA5D/YhLoLuJpA+pqpl2xhswJzsEsfN8TY2ZpL/SeJPLmO4k5
UITOqLY31UWkF9IMT1dIobgb7d2geHToxPBMroLKT7k+DQcnSprGKUl+ASY5QB8QA9IxO+/sPQDI
lKG2k+D+W5IREXtmk8jki5Tc3HlZcHcOtx355LMVvG2PL3cBf8+9RfRSG9eCvE3Lo77fLWwkqSPS
T0Jrt15e3fM4rz77aALzOUz5g0Jw8r/lOX+LwybSvjLujt2+psAJfeKJTJEUK4T1/p8WyMQ1m/h3
tGL1MocuHTddNu6APj1LlJKpGwKm/2LdRw34164wbk6yNMrDSewhl9j3PnlCyB3LkyaxsXTqxADG
NDxY/h/HCXPeA7VXREbjqLm5RRstjuRrlOACGXfDEajHi6UpMVwkwmT2EqWdy/bsYaVa4ner+3+C
mi6MGUqsnAx2AIsmlPOJxJ8vPfru9nZILV+2xqQT01f6o0AscNuHWDs1T4ZmeK24BIxE7M64Oqg4
xpp+Yn7VRIMQYvwzRkouJu2l7SnvAoXyiE2HkmGRDaGRQxBxrC4fczTWRPrMAwRjbNXwJ/5z6X08
LVgDaWoCdQ0gbakJyWDQ93z3sPzX++0SNRFWyNuQpmdG6VwKpW2R9shfRa/hisFR9Gk6meogcejH
AUSiaqgfw+YHJY2BrHtKCZagFo+mr//qgAUPFwDSuXZp5OrOBoeYko1OFkx2Jvnkr70kydFdNAgr
vDO9idvIwd32FdcSryASqHtppvjiTu2jm2Gu8MMHyVWaj9HcBuy4DhB6JYSdSHxOlnXAAshl9HT2
lgATE4w5qoKUuhBIzlgkcFDBcq+aC54596ebODp6LrEyCfrVCiRFKObe+X0vlKOzcN/h2F3Rni0f
PlWAdMJUqJI5VDIxkWDWUvJu59jNA7Nm0FvNEHdUdYhFTe0zQVp+ofH4Kw2FSRJgNYcrqsm0S9ej
9Bye/e3lLZxdLeTZakIAfXndC613aBOAddrIdzt/Af2OzS86lCZSwFunvn7XMgqJFAYBwCT91Zon
1soJ285rA34emPAfoJm/1N3FtVJK729S+LziVpuZEov6taL8JvNBSjcIFacQ71Lb2K4qabIkGWq7
cxBc7REPyC6ac15HGJ9Des8n/6nqsJChlMzwLo3hWfYw+ghwlANCN9sS0vNNO0j1tZ0Klz4diU8Q
/UcfDnYIbJpFntU2SLuQtG37MsKWfCX1BZHu2Y3sa0H7kRkRe1RJu+KXcPEQk3sBr08y9gyWjDHW
jDtASPjfSE8JGPrpsIGCDfkBNWR120TPtjxUpwbUBUwDHQTMm5ey0ZB/qEOKP70J77Pj2A7l+hMy
Y6dj157wg7Kg6tmvr0XtHWr2wTVzU+0wB10fiVWWwYH9hI3IUmoCGoTZ1+XQ4E9xl1IxBqkOoQmx
fOayYQkEf1O0x6nOVbA0P+woLVOOAjlTHcePcQSXy/Q0V2B2GiPalaUj3+66kM9de4YNCZRCfYt5
wPPNjjvRPXCO0jBQJ5bOubAKdtHuBu6zFAdTsLDA8H+7Y7JhP/OrwqnWN6Cl9fvgi0RfCcjFApWP
A6I9N8d435dyQUeo0o+P/0TXB5czJBSxpYTJS5nd2YjmbNJQWcue6MBm5JOCO/4n/bD2ZBr2rAUG
kGGmUQDZGeWksHwXrmVGjOPVtXF+mAk3LPFOq9jedK8Gj+q8wBIx1IGJ9OxoezxuB2OEYpI4qlzF
TNi/HsTlChnifi7I4uuNKu0Ij4d2QZjk+CYdJIuN51CrazR7FNjcGN63QMk1PKf7D5wVEBNYR0JN
CiPEx3xd5FqhZNAREkR8hRyY2d75/mparJVHbd+h0ZUrfDhGMIB266q5dIQikYor3wAask4ll31f
IEsC6Icq8GrPXuRbH44HSTeCbSUR085dls1/uCNV/7ggd8khGf0VdI/U2vRy+YUv/TLUwY5PEGYr
xhAZ3Y63EPb8mlpYvj6UWKII+AQIYfzCENW11cBT9JoRekTR1MmBwA4q+qLpfifEujzYbCSCyRYw
xb38z6uc03Vd9rElnLUVA/B3yh5wz915DCejQeMHA8WJ5zdCaobZWVo0qonjW2yJ3+rk5cuAhuFs
DlnMkJiSux8G/F4BvIvE2g1ptSejXL6aY25u/4P3Tz9A1tLdkMkZJ4vu5t6EI0cu4vNFS5If4J1o
aqdo01vtmhyW/yrIu0CZ/dQ3Upzdnq5Dmj9RvHokUxcEWa/KERv3mRSC9rCbInbY+UlXImLhZiu7
ZDpoV9L8GBUXwo50mQR/7JDnU/RL0bYrZm8Kda9zhkU7MfV7Wu8WhLQXVbOzH+GvDZmYlCG1I09K
/B5JHkyei7C34awgTLFKaK5AVhVeHEDCcz//qIZmivEDGlf5oLgCnQWHeovRWFVuO/vvKkofbZ/v
6FnMYNIs4vAaWN/O8U/HZXgzPyWG5yDPvf/oqgBo1BnkScVCBfuiKV7xZkR4fG4gAZLZH5RqVhhh
x7YtNl7tH4qWzayp53rECua8QssH4uaAKph//6E5BnsHywD0FrrC7py3pQUbv+lDUg7b7AU6oAKl
6S0PxLsfcgYdHPAs2tbOd8+B/Sv5KZsVIHq+r/3caR7WDsXk6nLf9BtXiUzlC+C1i8xmJXOz1DEP
ZRdJteIIrSWxkf99+7lZFqDDP5jGkkYm6hR1QzPvr2MfHfPGBM6mDOk1DYz5N34L4Wu5kVxtTo2F
j8krl+5KAexloDao4ToB0nnV/2aFJikj31Xd+Zxa6qhh2Ial5tX/x1LEaSJnB0zDL/YmZ+U9Opjs
FiPoHlZBPdh4+yAsBqbRrKyQiJ+Jp041rYPJIRsqBxQL32H3SuIbQTKyIYWjN5JnN1aFY1VOjBVl
ynU45YFlbQqcbqO47+yS69ufCX2sSISWzDQS6zBg65dA7YHVJVI+gviJKjvHbMQpbVdaQ2DQp/jp
vLS9Hmm6wTVqn3VJ8delxima7M2YAYxBrZFbIO0G11ZJbOeQnxV+XC37+hvtuuTpOBL38AVsoFMC
IjgCCqWHai/IUMXpmMtWyw6AtVGBf5RdCJBUoVkDkMfBBGZtKdZG17fvV0rDE9eKUoX2aGQrofya
53Yy/NMcOuwQQu+tjaRHa92DsmHvHtI7kN0/36S64mtM6AJnGgdBKD2WlJt1SAPoXmyUTj/bfkPS
GHDBmIESmctWgEEq+F/KavO0gTMnz6JVhRtrChsqK3DjCAgVRdLrOsMJgUjbMFKWS9d8IHFj/uxF
LUq6SiaKk7EPdR3YTPzQis9dg365foTMEhVXVsTo0wvxJFrOsUnixxkt2XCbBvB4xR3HpIGJneOv
ptYiTvEji+BoVPPFdqlH4NX6EEtlBCxsrd0nki5hpQ6Xl/G65Dov6THHHvS2QzrWBN8efGvzTT/6
G3R6iDh0rZQvrBUPg1Um5vrYKQiuswkdrjkkGUbQ4/l8+erJjtv8dkEJ/yhpfIkBpe+p+vCUWeLz
lHshYBDJdyih2kkg434okrmu1zRHE/ZxRGuxNIHqD4Gu4JCfZm1cASRSLQpeW+bgpl2GMxLBGqzg
PN2TdeJH8GnBQDp3S6bb+nZ1os5xOC/BlmlzB8dtavi8y6Kts6Fwvq6HLclLzxXEEfQJdOnGI90A
l4BrnrNox6yN81myf40ayBCaX9fpRqrJXnK5GHmBNH/HLxAxHxmE9tjx6+GHHU4bXapSE6Q9CjCB
ik2JCE77fdhn4xMTKj6O2XoTmteA6cx96mJZk4UAoCUNUrUFYUuxKfUvdhMMwCJY9b/WV5UvCyQm
KfMq+9hufNfadKJRH/iWh95/rcIwlr+m1hMEhuBm3BAeCsEE1ufgWtvAQMwsf3B578doaJQYR5aw
wudJYnF9nRcATLhZ2vzH+PjbEToGQgPABmQ6Dn/uJa6Ce0CfndpsqkNceBwTI/+PlqyWFsG7nlP1
ueHM4h/rVJSaxtYLiWLiw3RHQYegLG3Xq0Z0OxNjdqzTQOtj/BLgbURKaJYSrFtCsC0zRmZuWnT7
fJEi3ZymQBOgNQ7x8dRkkU6F+gkl5HXBQFRFL/OtHy75AvuSr5LDkPo6jr96Q1KDg3BjBz1uMKIr
FWwBeUEW0Pt6FpWKKGD2Ek9J5Ed5BJ6nvqeBr7FmP5ij3VUd2DJYtOj/kQqa3Vn6753eWc5eH4ve
mAzMibRJ+T7iwdxZOk+BrD/9foIS1CjfW5IejeG+9DewPfr4ECFhmNsM7ElEHRAysitYsPgv8h8Z
TkEbiqDeuygMEBCBbAq+zQwk15J7gJotqLAtC4vE3T5xRCXVTX3XA80ARByHIXfqBUFCh0Y/MSHd
G5O1FoBzDvf+5LVmrmRxEk+bURAX7FE1GM4Z7xt1/eRVDeaU3LoH63uJdhiEBvIYDBkJtU2jUEE5
KB+Ro7ilpt+na8hVYCsWl1iSN4Le3pATNhVlsq58g4mZePQlAT27FpjEdBmR4i9y1xkchay6Thw6
9uB9XHOr22JCXfD5JZpYn+ATnPH5bJmzHigq5LGq69BIYyYy47h0ze6X+h17COAq/bCdVeoBTjzZ
118GQS3lg1mWA33Pxvd5Dc363dO48qhfrQH1v03QbzOGHRSUUuR4qYWvyZ+2sGJUUFKGFmblbNrj
WPU6c3yaly8azDcluO9lKe4BM64jSs4V1me8wAfOnzZjAxOH3ObWyiLnXfrLLZmgcgox5o/dWZZA
V0SfHxXvBJKLK/q7zwCJ+4GrBl8JaD3SunHqFOTUOJfvHnzpisJzbxip10ngI8rjnmvbtHLHa05K
msURsEZhCOTN8zrSK5h0W2u+5zi/C7teBDtzpNodjiIq2DNWVBbANtu6x0Q9fYLfiB67sLq+KTcU
jp8E4aD/9mSr2EVNTZzxJqvImLtfGyMkjHxZtsOtKsHJ60fb4057TeHrdIeHkB2r2ew/EhEX9PQx
vAMZy56zAdyGEmcdqNcwXtHe34HLzPgzazXrP5Mj7C5hvBtI3+luUueCSTrmhqA4KijG6vpi+TbA
mPlkKyu0vxJU4DT5OtmFWbsd89Usa4PjJXSX9U2djgQeqbMULgJ5mM5FVuR1v4niAzyHPkiphQak
0lGpH6wSX7fhPgeRGP/d6qOSsiXz9Hl2lf2KipI5drlYR06r3mTwHlF9rQEiL1zY/iEcJ4U7vmzs
XJnLr+Ythsi7RyVKX3HKdSSNx7l/9hW3cS08WAtDCQ2FL83HIlPtvG3M4cfmxFJeQ1ogkXTjsVNa
gM4igAEQc/p0nhWX3K61MmsX80CqqJdR/g8pnP4eO2Q6aYYrZ+cnKuAbAyFdpYz+ceINWeu68ucg
FsUMnPYLwf3Pk+PBk7wIgYpi7KOD/ZQIH3Mm228N6fMWfHdclNz7rV8RpYU2b66P6kJE5tRZ0k/Z
QBcZfqyg73a+puXTwzS/F1k8fQHY3uC4LCkN4uM2yuwnuOjDBTISwvb+1UAz6VlWsB4taEpEEKd9
PBxOYDo3qvrLS4Sod7uMGC5RyZHp7Nve0vnrQV68K2EHKde7ONQTeLxLgVh96hCVMuhEii0VOICq
5G3C0730XWm1V2PNZhSyWLEGJ5q78aqAfnFj0+99Tm5pD31xHDgnsNIWtrHFMaN6WNi7XiZ3A7zL
ltRygo1CXGB4HJRIF7kyohgDz3DP5Os71ZSGeJAF9kX8wzr1Y37ZuKz77DWdQ0OKm6AjIBvMvF9p
timHqpiRu+yhJQHhpaOMJ+vVkb1teGtmH3M2V9Bl73tGJE11mSwZJ7vTIoP5jlOA3g8VlzcUfhW9
IkFPFArUGwaWCk0B+v9I1t0gi7cYm/bCpfpUioUmkMkTvWsGyPig/JM++4hmDj4UdGhgCbu3i84R
jeeOo1y+fcrN2Y70GlrFujoj5WAgyPJkRtPPfGo0pUyFQsvWAsZQ3E6VBwCmNdxmkJunf295wwjd
xcUaEbgtDh3hKkhBmedFBh+452a9CUB7odT55dFnV/MT2bW7cMwYOFZUGR3/Tt3T+jhezWQMn7Nv
BEdXEPkeY53/Yrm1RptSlKPo+lp6KvdzsEOHB/NoDvaPxRvMX3AziOvNJdxOVzSCcA6BZw7jFPUK
h2Ea2GOvyn+5keV8LdVHdf+6izF10mSnthSSGW0411OjFBmY14aN0fMkZUqhhBgC1Vtj1sg5Tzis
+qpKrfRbhIAn8SSfoJE+bjAex5aFjlBoWKO3RuU5dE2IdGekNARM35TadWhNgPV3IBi12n7cr45Y
Gzc95s6qpLuVZBKrDl37HNBV9yyEdbPnVHDFp3Tpi2gAvaLDas97AFL6GWl6610z3RoF7ZTZnAMk
1K+YpkgCT21D2VOrX0sh0PIpOLLVuSajbu42vRsETxueqkKAFhUN1rQ1syVdJuO90ncZ0C5YmKtm
3ECXot0YewzEa3Tqeb7EyNVkliOIw/Ke15KHvnCzM+WhlcPsX2JwmxpKgqSZJXDscr0QqgACiqnv
iuU8pwA79zmvt2w6V44lff2ztOQEaJgGrCVdizjMp4vEfFNwSl1l75t6BREUF3YqSZ3hUoPsMJZM
W3LsFBSnHizRAUBQyN1dyeE1wWI7BvD0c647jliTaI1v0Ovimo08zazxCDZ1W0uzlbWTjhAbPbss
E5S3T1JAlpQAp4Owz/TIZolevoiK1ZR7061QWv15r9EGGrFk+HO0vDTnQPtu0lBlPtCXTq/U06rT
9+HaZHMRQ9HKWbblcyFnNdd4lH32VqvR8/YgEZVAOh7KsHLiH8DNJNkwMzPoFxFuROb8LFEyf6O9
Zl6J3IXoheJtuYpGQf6rFbkQ3i9JgufcaguIwOUs6IwK8cAIhoODGVPYS3TCWcXi9P7uPHpYkZHm
YnWAbHmx1G9qTXeAM0NkNl8XI7aiLq/jWqRc69G9ODI1e2CzA1MZIK/Mgkk1nlVyXnLpNtk9zIPp
cbvmW9Snsj0jczq/o09yAf6PB9Lq4VETgwiS06wTqRGSl/PuRpxOnKlsveL65ZI2qUvB+NatFEpw
v/VSAB5BmbC6cMvZ0CoWH5DboJcJjlXpflIEneASxgUoRWp6qiZ7G4PotQWzpnhJXFvw3UbULYAv
ps+8a/rx0bqe5dhSkFoNe+SgtcjMog+AMwq+u+md9k4D6BLCeDoxvE6vcJ5gegkAx5uOt59NOoXO
/XRG4+u++5h/B2D/kFR94Cxp7KkSoZa0s9RsAM2NWv7YfIJpAR4onqZydev18AvQ37ipSR305vD5
/ZKJfFbs5UC/kgO+hVnatXAu/4jQn00zvvRuB+1diQ3tES5RcK9qVPe1+I31l2saGSx7LyRWkCu0
hVzFGFJQipxfoTpQY6mCS0vdxMPRe9qy2/3DG0s6Qa2NfeGTfhp1toZ/gQMUollUmHdjrvIaAn5x
6WlmSMkvyz5RKNO+YYR56o8eNg9lrMblm0Ir4ckEvwlBSgbnf2tmw/8m28FhFiEJauEvlBcN+HvI
UX0pek8T/Lv86YetdvoguTpNxP87ECF1apJXKknmgGLuDOW0hnBkwzhBsb6OAR4gK/iAck0STYlj
CPNCrzU7g6/0+2AgzKApiiLPPXbX9lN/otkCbJmfn6wPmGyDTrZdHbjlTzhFo/M9ulMorXa6tpyO
C8wT41jNB8x2p40AX+ekR1sE5ORkCNRpIpi/smYAg83oJAIUpSY7VGET2Qyv710Vg+QF2+IvRvwe
RYIBJ95D8VBAh7LDXJMMGACNvpShpCQ/gXunp3B2YGyvCEbZOXtjabnShA9eWWbHOgMOMoIBv9iS
ZTSxqPg2A2jech7o0/ngWd2SRBBUqidn3xjk/vC/DrXuSaFeuxXToBGzBZncIxvg34cE3opgN7gJ
qgx+ERp/+eLfeRJB7IsO3s4cqIJNhOuj4ov4Q3+RXQNzpGyRZrBcFIZMIm95BHn6FlS9Cbo7FldN
iZDH1p/78IjUqd0PVgPzJM7WDz9i79p1bjM9xdrQ8mVEUXsLumA83Run4zMcqTjlhKtC9Hcslc/s
S/j7kimIrtZkE1IeO9d5R/9f/O6BNcnp3N66wTLq+s17sxKUvGXJFUHnNpZfJnFeag/HDo100DDn
SzH3ccUsGJ//4MO/sYbVkYnTgYAsWGfFna1PID3n4n7FaUd5khlJAVXD+NlFGr/wMDtYhuMxqQux
EN+9Ry00oAhX7WOfoMkeWYo8Ct0GeGVXaHyNZ6k7uVA9E6mauQoDhjXNwG+Vgi5J6Bam7T1oIlY2
/xXVmxbSky2I4e9xFo+ourR+iOxiQFLua0OleZYpLCpGVw7eMzLq728kXlIZoL9CXbr7FWmhRVkr
HKEsTPTpZAtofhhM+0h4nghrfacZDN1y172hXs8LIW32c3S3lWZVK/VNt26TUpWOkwJvrsm1fBYt
AK7zihCrIOH099oPgg19e4Pxh7ix/0o65oWpy9qkGujArrfj7whtINVsgjVJ56loJmF1mW6VUSdt
Hbxrlx4nUQGVKGAKuGRZcc4DkKLaX3xPWTHoYL/G6Z8nsSIQIriSpo6ZUfar+ITu0yRD1gKYFQDv
0yExvNIHvUpxof60P5XJ44QIbX9WXiyambNCeFEvBwQGXr9wyrBwH3rkXmcMf4dxt4HCxsjICw/n
QRy7yHr6byLF2Bi727V8zKdmoYJRePYQJ1FW5lx2zwabeJrvMa3APaiJuvsm66OwG/UwTOMai+WD
eLLCsh7MkaIxlAxybw1eIQE2qQ7A7xpEGXaBUK9nUJvqGNkcY8IO4ffDtN7lYcPmDhxbXHwVr2iQ
A7YYLqf5b4Pr1P9qCJUY9T8TxkvZi4Jpr4/7P5W0qxA9Kt9UEUXZsihcxN48bNhQQvq7rqQ+E3cN
JxSuYS4hi7RtB0MF55ByQMjWFC72Yk8ElthdbyJW4Hpnue3OJ4i5Ee+/5REcyGaqthMMfnBZFfYN
tAyavHV55TPmE65PjbpWr3IqSOsw+yJwN/3lstxhbmrDVnZdjkPZ/8xyluHIcVgqMyjLO9c0jiOn
0H9aL1g8zi4VxZz7dYCxPBg8EUL68G9FDh/fz8E6cXxNIMLoMd6NDHJlxg5J11sJuJOkz+UtBdid
+zp8kAIR9mAPpjtCmySROQ77qgWoyQYG1RZtgFIqcH5zhyHVH8M9iTCLKuV9F8tHwQz3bKIdl6yG
RhF304rXu8zNvHWPrj76+RxB/URT5RjWkx5zJ3Xp7XAVKfESWX3FzGo/RkX3yT5vVPxYsY1wgN5f
6Ky45ScP/BC4Y0YPygm5nKaR8My+84cT+G5/mStMXuNh9ouOvcGn22JFKaYfII2TbxdcpSzDmaYs
/+SJMyBASpmQDd2MmhNDkoYrxHjfClZCCm7MLQfTSBGHyQ9VSC2y7Fka3QAy+V0eCRq1D0KIWSMV
lT1c8PTh8MPbBmhaY0NdPd7rjJcF2u8/PVAdS51nY22uEPSNdbQUipAAloGWlCZKQRuTR1ejq19O
p+/Fbk3cm+QXk0aXB2z6TVw30TexIQ9fkALsLFSCzBVyh0jKiZoQq1zktmCjgcBRQMpugXIwdEkE
jqPD4iIDG0EzG8e/DPVXQQLbjROCe5UPJV2XAfyYJ5l57y5TTot9jTtiAbOa/ygruFcaBSEK+SKp
NB/rWMoEPZXiVq1g7D8z8erUx7UqMTe2CdCWmWuNVlVKuTdzxT5Ny07gPhnAnWK8AaCNZg4Xa+v2
SCfEy2N0CN87NOrOtj94qMm4eoZnadb5KLkplJSquUQMskSROoMnSNPZriPxatoDLLvYQIn6rJTx
2JH9eB+ozBVEYN/8UOmDXf8s4YohtLZmWPUxVg0vLHKon/HaaAKPSv6FRZv7lzSti/y/EMpS6eYz
rSYzcJmB1N5GzxhFSY2/qxnrBOEL2EWwdUTJFU2NHcITc3TOssdb4iUDhBqp08NHcL4XvXIP5cHu
LiTqpBldS4hbG2y4RyT7oD4neFQvRM14VHdmU4WxzsWP0+knBQM+ZPh77oClTP79VXIk9gatmlw4
L0sAVvM8VOa6LPtERR/RgMxS6BgIUKlPMwkQD9zLTUbH67SjSaaCAz/PVoOCeedwGYs1ekjbr4CN
V+T32RqHAtYV8LEMoYSn61Gr2NUX+c3sAbXTjk6Ckjh2bMro+rpVU1bfvhdSOE56tHSNbjH6W/uF
rLOalvu/l2nXIdVHEEHk0x5O8Y/LWMDXKAgCg8Y3keTlhKZu6vIOVbmlQjcLd8SMBSY8Eofgbaul
6mb1EthVoxpyX8mK3korsxQ8FzmrqMZlKah8i8zCFJKg/0CYXBFN9WNkxX14oxITscIHAy4Nl0M8
HftYLGSYK3JpUfbNhQKIgWYX7648tMZtdZjSy5y6u45hMGT1J7oUrubwU9+gEoNsdyUNNqkRq3r8
n6BJoiBZ6TPFiOdUE5MJb6CV5/oLeTh18Qm2LwSH0NuyzhaPFjXY+H7t2ZO2D4i2jkEplcNmdYbI
LV3EdggMntaCNerEVAPSq5iyrUq+lKlQJj+t249epZszESCoV3aJLBrk8gWyte3ntcgmz3QV7mZn
3ISGrga+Lv2nxMAursFyXEtcJ/z723A4Cvrv86oiSPD3XXQBo+50MERVtfY5Qzwmk+7yspI8hGLE
pycJBZpg6yJ6H9TQ6/5X2+YoDQnfWZbqy6cuf5ot2Q9WWIu0qPcf/DzYydgNhNR3s5fN3V2mYJie
6tH9e/ERUAaoqw8G/3Uh83+g41lBStyc6d40zHt+9SM/Gdci3fZm6e2g88cDtCHiAQIsYy8h8VLT
ZuEXn6I586gvR0CaBZ2Hq9mZby1OtuJV3jYNDkXLSIuO06lrbMfuCnKoiWZB2jss8GbyW0qhHZPp
uUAJ3C2hRw5bdhYp+/xPHXZL5Ot/8E/yo69gZWB8RkRGHh8WaM4Xx18IsUCMNwcTHIt4xZtk15oa
oNwxl4/8Tn3gBEl69MH9ZkKRUUTNoMiHgETZucTSwhrzRM4tzyqGQt9WjF+2jTDy7G0dEgg9fGM5
RdT/Ve6ooC793EeZ3nxAtgWht4PgGwRPPZyNuIGhQgJ8gj0PIYqklfJloXdc43OXDxEyPXiIV4Gl
7x5n/7gRXnVJ/v5MSueOziV+4d7N8COR0zn0FhYS/1d65zfmSxw538YOZ2vJt1TDi5dF1clcGoKW
kdU2m+cBjFxPONs3P1RR/3doiyFPE+CnzAiDTPyxoS/mGTVtg/EAysL5fDY2GmYNEAruMbylrAJ0
J3PUnLSvRVtlRwyA6VJwQkwXaoF9s2UQxyY9T+FL/pYoK8Q3MR6tEEGCV8ewL+5WZJqPc9EgqYAL
72+6anz1AtxWkbe3qK0O9daxU4uBLhAxsEa8V4G//PJ8BpEVgqDe0PAp6//VeUeQkpRiQNeHkAfq
Ohu1Xvbrha2VrA0v79ExGedKOizhrMT/Uo1X7XHT10j7PcisF4cBZsn0Gm+n5OQoYm1JBFAXxTxU
L418duoS39JGcB6xPIq0r+mPW2RvxLU8w9ZbfjlVHiXlmbVtbjuwKG0R+50t2gNi6Il/AoNa8N6l
2g0PLt31PLFtPRdPn2cDgDSOSJAauWtL7dqPIJr866EkmKpH4vFecAFBEykphlecxKoXvB+MRWoM
NSFHmaYUu+hU2xDfSmsTA7yI8V3ai3pVum5tTRxsDCwxf9AaFPLYpwI8tsTsXxDbkwKphUDudTl/
sPeroCtAyYmiNHJ5i3M+y0d8nJcNLkcU3ArNEftQP2iS6Uou2sOA+LAxelOjOHy0Daxap6b2JNCE
NbCt3IcjV1o4L6od+NgMZDArwlSmhs246hrfOEi4tTCcHE7k3MxwAmpF6vpj9wcLGuGSEw99NAPc
pTD74yOpymsS0hooZlD2eKEDvsDuTZkAgpWjMpFxxgZjT3+9CLRSyCQbn8HjLw05gbGZh86ZI/x6
ViBsdggURQ86HZ11K6ADb/kazneGy0Gbg0Pu8znToSYUwxAV/3A8b+dRoLWHP4EZSjrlQ9hfjyG5
8TT5MHAINWSfTBtUMrKznSTgkoJ5Pwm0P2tsYBQC1x9WDsWpOIWwdgEC2dli4rvbNbJIydwtC59P
PmApHYCFmfayMpJHk1mi2Ugm27POrWwi9wam0duVpBim+sx3wuP5NwjQdIVPQVaGxzNhDbfITzmH
PfTCJAezPntKXgcBbUl3bgvXpGqGVooJpDGfTwXEzqtQgU8FjxPWFESmVxkG+3KKsp+SJCwnBDq4
yTiWX/brCTRvAgvmhgY0Hakcj5D1ZaiPZ3DiVMia+T6eok3Sxse0FkJigdJ5rg4eCmcBuU7s72rJ
J1dxbKD2ZwgIPmdZ7Q5FlgyHl4TBJVGf/wmDY91JLOUOZLBpGLPRr3wSkEcxsTmZMGVhLf6aOfKc
A66nAyRBeOcRrgajpm9j3VBHzNWTgca83xLk49qjJKsmbMrz/vmA+mtZ2ggevLrwfPeEZAYqBFba
uz7b6JvMfZAKZIz4wonDew/C3O6mAjHujzEoXNpw0gWHW1OhUHzeH4toqcWuIOALamGujr7eECiq
44hgwK4AXEvBNMzBsZzmIhecHB6d1UZMjoorKmkMftnS2GLOWzHcZ8NG94R8HaV2j0xLkJRb1sUs
buNxR4uI2rODkyet97HLRHCOOPQvC+ZHHUB6GK8LWwQj1BMDn34oWtyVj/gKr+lASpZIHeD2btP2
LplfQpS7Ciqbe8XMUTXf7hn4GgITVDsBH4KQuxGeRdRAaOO0FBDXkcwTo04cpcVsOmTQropU/3Xo
oJK+axl5GzhrKzfVWv2VmYAQlY+a9fcMoHColjzmF922449zntns1mGOGs65aLOIXeobFA+QQODN
Rdc+wHTEwJexewy2E9A/Mf0OdNkiYUTPffpFL1B5DFkWS79DIdQvEWof664HYH/I+oCR4ERYkUOK
aCULTlXV6a2sQmOu8m/D15Lv08Z6PY8to4OvrCWAr8LjaWloJhdBlHRVadAUMv3TNyawA1qrvVEY
Eo53R4JAXe20/eoeM+VKVW71NWGT9x4smmhmOuCx+BwOwPOoGvimYH16P0gUfVwBVm0ibXcHy0zC
UGrgrQgbPj5zyWjlVt8ojFIZJljgx54QYD+tdZXFd6FIQQ0U2Rsc/KWv+6ACP/1jdx7cBZ7PZCyY
4YO5aJj61RnlPKMCRlhkHV+t4i0nR2U/UPt1/8fRR8KFecFEU8egYIEshWJw8vTWm4J4m7Ykwc7V
gaWoP3vNjTDaA0YAn/rBLonaG1WpJkdgmYFG6vkLkGg+fYqNdQeJAPGiUioH5R/RWtGqn1n4YUfD
m63shfQOhulkVL56uAHQ4unAkI4/T1z06s4DfgRiy76bwpSFEI7ssAhi6Y+B7/pJ5vNL69YrPtMJ
lJ8sKGKwUn1GJ4PWvAMYPbncOlMM01HS2L1kprZ+s6W7/ICn1BUYNha5I24UgL4jSddyesLJXbb+
AbFWe2UyusVycTB6cnW8NqsWz2RwlVH7ws2y3yOpNpoZ8C6Yt4qVedW3hNK9WlQEnA5jTLIcHshJ
vSBY95PPnMFyrCFFDjlMoKkYIvbjpou5MjY7NRaVEhwiqH8tGnGQDYPpFZDLv1Bln1qEGH/WxTL3
YDzGYbH2vplWhz8Ut5UVvZaMsT+JBHy0mRGSmGoyVIr9Zi+MvZk/vcbvqQ7RiOv/IMq1fAgzuhJh
+zoeA3SzWiSpEKEWwmVwyClB85AZJwYuZ/qOrSHcDamQ/1nrokx3DHwoK1HBsZs6I31rkmjKvSvz
lNHEfjJI2wu4qCTUX2PfZkBD5LaikHYvdY8jB5iejo4SlopbFoo8HZshmmDnKQS7v3/2dBoScp3H
euPMvyeSbUyzeVjLjDrWCif//DurVmySgOuA5A9EUh5qTQDccFI8Rv5ao5WGoZhbGWs7go8a1wNo
zd52dqf6uPyl5KOfqr679rSgirLZy+BWZM+5VMOW60XjXHGlo6r4JlHUVIUeRnvMDKrS2Ol/m5on
biI/nRHJLXwFKYOSeVH9HcjB/+jKYC2yN8g15lSJvGFHHvNNVNBQYXBNIkMGX5/4DkrP2+pawOml
v9wKttZd3k3aCBhl+kXZ5a2fKGVMCtxP1JYYky0Cx6U3c0ojl1OZs3wH44fcuTx+OnAPn23J4JdH
CgicF1MzTm+qHPgh4/eH2hnfYWgxYDfLFR57KPehri4ZZ1PhtWmYeg4hYR69tRL/NYRVH2F+C/pd
fQKJo3SoN+ygeFI57/zusVeSax0aEKPs3bs14Q60c0CPEBEgP7sdpM2GVeAPm6qFxInMGyQci5zB
dMdSI865pmHqIzysn/CsH+gULxdNjrF8RuDjoSycQjwRuV0fQpHsL8trXZH44PD/Qu+KhVycTOo+
VYD1Kh2/zM6mMGYn/Rr71EQ0EkDGgI0hyB0bIm8jNEfI9ExD120gWFkdZHG67AWS4lqSlZ8Xloc0
/sz8uPMp2Pb3y1UVQa6RM6gCDIk6sPetkfFz+75ERfQWjeMLrwFVuSOfDAXC82/JHcZwJq8Fze3A
cH9SnJsqYFB6xMdU4WFGo0SBwjncUww2/pIQF5SR3oJVWGlOuJgiDgIrLz8X9HpAM+cAHVMf8Ja9
xjFVPPku8LGPHiBLRzijHX3fPhcAf9yLCVIWwf7avHowPzsVP5WVZdcLBJ2NGDzd+id3DPKY6GMT
ef88AfSMDzTZXXfI3lerlZYf0anQjAAewGPh9a1SvShMhlbr7leN2IneRPmY9X9is3w1qQf0ZD9u
7d4RMtOabwU1xk3u94ebM8+lxhrQr4HdMfZG2q4CJ7fZUWixWtmECkkxTZ6J798W6dZCm0kIE9GB
ioVlJeokdPUakjxbZa6nhXR+Aw/m7qpMZ0xXhKzMwiz6p1pFyMXecnalPqN0J2XHWVwNyeFOOeYp
924mdglaCnL2VPsMjPEuaPIR3BOdGg4w1Ulv1NvB2zqhYmHtcMjbl3bT5r0Vf0dx5NmVSioly3Eb
ETK2xW1V0qj498VQeobA8nD+T2gB/rA7iTKeF5YWT3wWhGrrPb/Xj6pS+GkWkGc9zWkUaP3zOP60
w0KJL4nLyIIU0HTzSGlycsunYgkPXKwQ/Mi1jP0XlWa3GWvf7Toe0ZQEJrAJG6v41qDtHXM2HTE3
siy/VYOIcBRv/Kl0rZb1jmf6eb9pKtnhoB4tVPzDIr41qWs6XGUfE9mMcJEAbVaD8Xv1j3CQn6OI
RyGqWT9GSV0YZbCU7QVmMtgMCdnsIZCUVEJtT+h5aIBg2zR1hxyJwNRNz5BvUsQr6z2eT0Tkzvwh
rQPhDVdfkyR8zLM8S/QAhpbFHhoqDAX2O43wkP3Rq/pMmAHsxpEsCOnkEN3Q0Hb8qQx9zsxH3uQs
2zIMx0S/6N52XuYu14xPofH5Mv/n/Am7C8y7lC2iioPM6DLnhKl0csqruMGbdHfDFqTSgGGC28Oj
4biXPOs0c63FuvXAsba3JXF0Vbp8Dw3aQs5eD/BWERZahKRKe/jKoYNsVzyFJS19LuSkRM528MQZ
6phvxVBn/LDgjx4PKrHq9rZcQxg/avrySghCNgxkD3OzoBP8YHpeZgvuVGtPUonM41PEATZiOt/J
WkhmEOeBn7zB76M67y9zDYEd+98Ht6VEjmW6Lk5pWvODF5UdpEEDofpjR/Oow9Kf66ff6afgt+Fm
FTT6MIqRhFvSuulqNoNhoz1nn4LPbR3aAO5aBBiAdF0PPynU7XYRUq37SBPgebXb7W5lDE6unluo
uw4BM07pHtzrKCIhLm/nxuKWpHpU/gacbbKtg0IrUt2VJhx6UqsWlnx6dwTrL1N6YDbiHHeit3RI
rowawkAJCK+OyHKjZUd6nIQPI6wFDgBzE4nooyaqpNQGoU1aEg1NP7YcAbTYEnM9I+d6EU0ImGpg
J3CTF0SgywhhmFdiL+qek38w0gC+a1lKKOsPFA4ZEyL/sLXLyvWgHpeJVNECUM7aEwVFPv34DTCK
6ep8iVfgN9GRJjbjXguHzTw48vWvNUgQMc5wsgh6beiEIO5igd4CTi+XszGTAveuwoIsqbAfmYTC
rA52cHHhVV+Yb6QZN+cHMk6lP5dLoSHCC24Vj1ukZu2baY1wyqjKIeaPYOQYl1hED1hIjwKJJWaH
H5KfcuNTbR82Y8eVY9PPSjYSZ75YyWjLFmUc9SghMoBlIWQ/gJXZHMKeHUUqoL74qKaMLG8Htob8
RW8nmTXE5gSW35rRtH9aE/b4Dcmt1KoVLqZ4ObundjN3TSNHqOMwZkkJOO2tB7mAN6Sa8+jdLs+3
lCj9lBOibTyCC38bVxCq1nOWvSEeX6WXM3VrGVDA+KK7YKvM4HhKeqS81JIRLJKS31RySCMR4EqM
unK3ZKFd3Pde6PWqCJN1QvW0v69OZ4N3KSebsSfnyILsUeasYSeU5CeyONb+5Rqgd51G8vgO864m
kjam0669SuYAcCalz8h8itsATXrnHfSF1OyaBRQ1N5dqt/0asFC3R61/itXSF0QDzpWFbCX9uHc9
Cn3Jr4Va3nxg/qj87QONuYIblaBbKgLqliuhDPvZCkt1aoyXLp5ehGXALmd+fQnRQ4OcJR+E/ql7
vCtNGgUMfasWk2QwPnNGP5PGXB5b2I4PH9yNFxhI/YSM9e+kEI3dV2N3WuhP/kKSzt5PmrS22laS
9uDxwXVXnTJIMjqvYfdOY3NLMWl5ojPGcYnNj6mvfKMzyHvvpgrJUuIDZxXwnwk+ocAQhyHnBO2F
Af/ewd92xpg6I9BrE5Bu14Ffa0nlzK9LPSN+TwQ/CQ7B9VWwko86LzT58wR6raDSuactddBG25H0
jTD23g/HaQBMpXCG4xBdIDivFqwQwmTIIM0IL9dfiQPfu9H0twpZ7KRM3NSMP4hsH9WVkVWA3xw7
Ttx+eKTHti83gy9dC/n27+ebc7olBGlU9N5Su/cp+H8NXeF2BXt+7e1FA8hXS6EWSklpfeCssx2s
ExRcZEgoj0zv2eJ6vtXV4z3Zxwk70i+oVkDzsVqRZADr6QtSjh2NWbtWKARTN8wtO9YIiE5JocC2
Va9k6LXgkfWefBRfCyfxOCrvYD2tItI3PqlU0i1FWRsrVTm2PV1wup84Gipsq/javjKdui7EIV7Q
P64HMb60RFVfA8vxyMAQT9VzNSwEZrxleXhFOFVbMLErOFFQsc4S6/xWZTdSrWX2IIThHOBd4Noy
Ol4efnyGNcd2jF/Ek0SMvGPMBcu7gWOlstpA487yoQtrZ+BdwNJaY9y7q51lhBiuoHjmQahYAjap
t1bQYpqYSF8kGmcT4hweIv0XDPKOZkr5lsd28VWhy9iDO6pEw77o+byLU2jIS2hrVJq3v+Yd0+qz
waOqZPkRA+xrZd7HsOlEiB5qH4GEDsoI0Lt66tglXTGQctKRBFykIcT4AwV4XF31PdNJkWiWXowA
paN3HDOLtHDlpJ6jlxsZNY1eo4uMQ9XIQD9U0vehnex41barpqxoqKozesathY6xnn86aJbpHEXk
Pe+nrl+rmn/g6Odr6K569NJlOlKrpTENoQnu3IEVgSJs/ZKeoYGrnvG/vQnwyNcIvCesE7cnrXib
guj7lEuAufcyzzAEMPj2yJ0hkc4EVqWEaTRHQbwfsZcJePr5M9MORyNhTyNQwBAeU0aesPggfsug
SRXAP/4jFKMQLSO2RSZAbqp3KfBcHMUmkFWUvYbunhtnKhJFtpvpTaKRvO9GDOz6GK1rmXmmeIVN
MPPZ4DQxdwWxkiGTVgyfLJKQkz0yk0jwQbdMpqVx/vQdzekRPee5Z09EY+8MgtHy4EYu/7z6C+OO
eMDpGo+zB3g1WnfLxdQAg0qJb4ldK6+TIrO/lMj7SCAL5BFOENzXvyYA/3seuYgp2GxZeju9eek1
3wMT08Ycj2fE1IGfDhe0/C38NZTS8EikutYb5XpSn0+LGhSS5CCJ9dwfM3FvuJ/TmzlMyGlgINzU
Kk1wZ4l00udEXO8W9JJAC8bCsMfb2iqJi8My8IxlNuKf3vdV8NTHRbRzbDnw74GHHiQQkb52YOm/
PAuDYCMLKh8XuB/3T0Y4b6WgAnnjankuKeFuuuOgKcN0y94cn5qH2bgQ8zRRBQ7i4oF0nj0dbedf
WDaAf6cgA9D/8kVbbOZ6xGG5wbvA2WTRF2pw9F7I/nJp4eNI+ynM3EeOCl9lUsvmruu2GS8RGeZP
NWKMLz3lr7Un3BMJ+MM0FGA0EnAlO0nILxVB97CZYnD4g+WcScuSD4JZ9Z7Ri1KNF/YesN+I8rHF
tYEzLONN/PaHl9QfS6UHKqyVT6jQeSNnf6hzpr2mVZxSmz0EI0QlouDBuvpFsgz25g3Qiq/PT4EA
wmVcytpsqyA6njxm1D7wa63N5SMGWf5lGQseu4MebSPQqNSlM0EjJcyASsG+NG+uIShn03mr4DXt
UD6dsp9DhGlkpv7josvErm8USxz3739KVXpkD5Pia+ZydNGLqwid22XYTtjKZSbnC0rJTNi2ZmmU
RhhjuUiLEv8LNzRfIv/rwd9R2bcc7DZmFcjA4nd19bPw/Ykqqn9D6TAwX8F2kw7wpqwk13Efrp50
MlSr09J/E+pMcEek3JGgMkVPZuMIT3zuln1WuTjTTF7XygCOjyQx0iSCqFC9Ef4OnfQlijhL0Hzi
HRubwMvVyrgB9qKJ2pGNsOlPSDqUAaTeN1BqVYZFN8Yb55Bn78EbrinNIrd56iR0+KTtmyQI2hCl
BDIGo0HOjpOk9S9XIpf+maFvIMowaVpWlDIhCPjs/6mejP0ElMUEM8/Ugk7tKO1NGr2KmwLh4leh
XGYyFDIXcoENIHEGguETdhSM/Ubr5M2bBE0GYqeoeSvX7ZbMEYvD+1fwebA3ZIDFdT371VBBnE25
0MvONZGRvUIzfEIoCBf13JwBFWEns9hu4eEYekC2e4pmXaQash+BQwa2EGT9s+CjFyqdTt4GmlNP
cMpC3gAw6tQcjuo3YFNHJJ+0U95A926ywyxiTOhdM8v52/JFGW2/iWVs5GY+xzCoIseVEB56mtXn
PCg6ssqtX7aT377Y91/KcjI0TXKdUbixIJEM02fx7YdwIWOCyfLPlXKMV3j9l53wgVbAJgRgcP+M
fubhNw7YGBYS/n9GZszaMo6sVQo3nMTbCUPnOMquOJdzErssQB0CmVGUjvlQaQd5kB+iv0oTdvGj
zHUR6suzzVXqZnPcUwlo4wI5XCyJnVsw2ZOOugrKf0UiI4PZUsA4XXLi8ojvvBePcyTNslk2RQOk
w/lZCNDxwcP2ihHWkUwvmQS+1jbNO03RYgIevaniBjLMhB7BWD11iS4EYTKE+icMVmGxdYSP4i6z
wyUHu25ZwbI/LKQXYu26xGWQnHL0Ac/Y4QCEa8PLMjilX6I/D9qFyyc7ihcH1NpUBFXithUcegeN
8N6pk+Idso/ZM5lgUd3Nbq3nfagayh3AmHLlcShYKqKUzt4kZI3moHmsSA8ATlZspThVRLiipfhk
/4Yj9KeGLkNLXdTiAybk98AaiOOs19krSwI2gY1SxMftJPgVZDJDEFZ8nublGuiYq5ih28aNf3Hb
MO3vqBVSTfeEXycKcj2Z26z6+orKh+HfCBf5HIBXTT+8t/iQ1zvXKjpNHeMCZxID+XK5CIl6RBCo
kRBf/7UjMHxrxIDvrBYNt3kwyvZZdv5EgV4qZkl+FOB7gLGinvyoLjII0QyUZiM0kli9g2ZMx1sE
YFQtdZ02Mp0wesic71Be8wtvELGJasA0AmPk6jZlrJarXYsuJ/jIwf15Bx4z/PdEtAR3NJ00OiN+
Xpw0cFbSlTaGmnaoC+RMv35Wg1204yLyOuXgxqL6SpdrfkROYhR21NEMZw2Hhjn4Qkcc/59fCfVR
NekqT0ezlFa1JP1L1VsSYnO+TSJWtPxOTLpuDdRMCmFXEX8u5s5b3ZfwusKogeoo2dcmrTS7c8DF
ebSUTN5Ppx1jMGSc7eZmYoteHiPuEtPcA9Rwml2+o/5azWCjipv4LXPlrn4qcUHH1NQ9vbflzh5c
KXh2T1azi/qw5I+Ii5D3d361FdILE03z+i40ZDBz8pKhFzW0yvMVRg7h4MYL1H8lSxpDA+M2fPLB
TjElDM3IUIg7pDxO7iM8xQOZMKcs6yMJRGfkf3E0UuAuEMgFjyBqZKWp7eYmPop87yDzP9VlWDOi
ZyMhBoV8qjBlBj38VnEsOCAQNwh1JUYouekEJPyNKveFzWJXZ2+T4c5DYoq1HXDZ2939wNUSuQT9
hSWKD9sLO3zpM5GVLgGdL+WuCL+kVdTc1jcr7dAXvuAt0TTOoOz8ArdwATMT0gZ1aiiGi1Q7kfS2
ydxOQFcBR3V/UoDL98RL0RbPYZcBtvwr/6KnAaOmLlR4PmXcz0cIMlO+37JKvMQPSSdJPlwdYBXU
wU1zLfBTO0903drWzLYbkIwIx6pNeOOBCGr1avTWlz0fwYMzVuS9b9XxNQ+B1dD12v/vSOBLCyIR
eRNqukgRb4L6q1gTC4F4tXbYYf5ewHCQ5APVuUGfVnJ90x2T43B4xmYyvBTtUhBwtPSSJMYpbCk+
Ecct010GPWkpuAhvTEdUXQpLMilXNaxTIcKHlvlFoYqBahC9i3zwJThbIZhxQrJ81XWgP7MrVx2P
K2NCD8X7Qk22UeOeUhhtYqcvAu5bmf4ZGEOuuh5VpK5niVkb2TUYq+gUCMCtBDakPmMi3DaXpWef
VTD17G8hKP48P2DuvaZcHjRD2VSm5mvS1GzQhWlLnO0oirm5SfMtBQk93rrQcb9xHUIhzhenuOlD
okCpK7AxKd6s9sfC+wUhw64VRsfUwPM/MFxTKBFdd5N6P5a/uNCwvKgyXkpafI5qJuUKu6ERBY4j
Ifn88d8zIVQXvhH8dcrHDSfOUkR3OHpz9aPy9Zqm9igPxiDlinZCD4xmO0ax7gFOyuBTEy6rN/0f
nBdes/JAezScEAeiMEkGHUclWVkTl/1cTW1WdMX87T7AgDPKUvQKHcKfGfXMiVe6rSlaEQ+OphYI
gLFf+3lVJix3sXmMcV19MQdve0ppr76yUJ8vIM5y8PHg3TRoCB+aaUF9nPSDmP7SKrmNLCblmj/+
1mQDPEu33WSNr+Ct3yuvxWyYAXWT889xguLrFKTP4ovkDhLRX3mURg6cul4jlOAQqkJtrb5zQAU+
lHJaKS8F3epU93UgCDlD6FXcO+EE3egd0m4ZQqrikJfcL5Wt/AKuCaokblLhwPwji2nwanaZcs+s
ra1FBSfxkCwPprwPSYaN1ldbtgEXDrnTyLH3i/BaAPiaScJ/VUCE9CqaZ0vZvbTokvKbwRrYs16/
MJzbTRhPB17CLgZS0bu3PKoFHSgmCG51lCXwOmWG6xtltmywYGOw/YUYUaq/IJpHZJZydYON/w5Z
6+lhEAGG2YftbSWWaJbAGG+hBkI23BCR3armyLk++sdKAD9Z7kxbcvrZ7VABzdjagbGyM047VWfg
kkSh7LGBpiDMK0yNR+gzoEXnmBqBnjWd8mMw4hfTDw23fGKVCh8KSPzR90UJimJ8ObSksF0rO4a8
Euq1Ubq1LiWBIAJght6n7wsQ6moyxL61N79TvXs6MOzlbKxz0tp/Nb6oA2PI75y2MLSpmFAtg0Ht
N+lPJzl1Xz+zR5O/Qmysy88R5ynfN4Rh9/FnSSbe+lLhUOWpyr+y7QIzlLCVR4KPmIA0MKjeN4N2
S+9lUVJb/TcD6c7ISMNLHI9meli0nMmtOf8j3ghTDa4ph5X6Xe2p9D5xfdtlBoJY+v69bzAyOwwZ
iKHyDyzN+wR9boOP9AcO4MyLfniZwVrox5/kSm6X4PCOARYIP3uSIWALuqylWjwyXqgVdbovGvQu
ixG7gbecRO03hatHY9RrYxa4/c8UDIazUHkBR/uiunKWxoi+OcWPxFN2iCET44oYCuAcTGBce0m0
/qGT1VI1kcQfkbKaywR6DnP0gcuvdm4mNqFamfiKAPaawV6girTxZ6IQG1GeXbXd4E5OrhHT3X0E
qbV7tbyT4E5Ap3ZMLsLfaLyA+jcQy5og1d0x80VRHgeA70kJx4dRRXR875cFTqLcoIOUT2SJ1Da6
Wtdr2BIKzz/EVr/QGZo+5brS9ASqbu0lpZm8VYwRjkBWGiLzTAo5zB+5v/PY8fffl4i/bI6UrcMf
SIGpHG6wumGByhPnLK5wQCq/Bl1jDrIs/1/8Ovq0DjWJPYgJjCBNqoCMM7jhwT8NPrX7ExwVrbLr
mTbXVuMpfBUcQF41vz5eZEyiIzvOeqiTSs5k3saC9/xDshjnt00iEBiv51TEfkmFnHavV4VOdCq8
Quk+7OBFGsD/KkedNbwMGe5NcTzt4cPcLeMjbLWehbo/oZBm1NDOjF3P4qot5dELXygYA0ePU819
L4D2OqJdNhZOJ1qjsvTR15orignaJrs/hMp+eflASmpAMAd4zcl67Bg0sj3a/5VxoMbRWF7WL133
KA1M6ICFLSb56n1b8VJ2n1upeAiqaaLmzNE2rJ/PRAL8YDn65G0B72MQAg5iqrLLO176xxMc4MIs
qk4p3AVfaTgxf7EPzLb5CsT67/kCRE6DyHFKzMr12j3A6ftqj8rB1R5prfln9mW6brePiwZu1itC
tmX7A9R0dPhzjSSvaInb/XudDmw93lXuyXXLV//MdKTJ57y2tvxpe6mx+FpFfNNzRxWtlIdjskx1
AM2vVlaUnBHUxA/dXwS13OxXvWL6Ug4JH8lKzL3RQejsespDvPoYJFoFwKWyHHZWC17C09witBzv
eHn3eUOJboz5FpPYzPnn/NiTPltT79CDcj1HJuMQaY7/kx1IKhDiYh99BgEiX+8bYzhzx6W+yBS/
iNCz6Ym1ppay7krobPierirlJ6KpGfoUOovgNXxvXT2ufZX4twVaW26LBfAa5rgEONQxZpi5KrPy
NhId8SezHDjJEak5t95F4bCpu1rYl/X8oD7GVjOeDJ1O3RucwpTUl1yMo2IoRRi9sL9AoBSSZ8Lh
cqz4KdCHYa50LEeGaY4wo+/DqMQNCyHgy1MAbidD0C1KdlXZ7pxvKXXtbofHuuVJTqaFuptRYKJ0
p74CxfXOCytayO0pWBmXCyssucQD6u5sXbV2RFd6TbPOCj4vxm7WryV5kyd5jl33Cgz3dVd7Ipdj
qhvngdcQx688ci/hxC88muEmVNgoYQWAsjJVBJQUH5WoA+a2J6VDTyIO+Oud2Jv3rZ8W3dmga5Q1
Zx35A+1hIhOcycb8v9F7oi8OEuX/DbX0Im3uvuy8HXCS6WHUoZ1iI8pR5WLgC8jFcDqxsGFDFXZZ
4BP/URm/9k57ltYA1vPvLj8UADVXPyV5s0WimLldEEWFB6mL4omy5A8Q+jNtIWjqRT8zlbxhNaGX
izByPpWXObVC2tCpWzgX97R8lA1cgyn5gpoklJSSpgP9E4Qk3I0blh+NtYXhE2bIYDK2pGbM7EaR
SLnpm1Kd7aQui8Jnn+ms/hMOmfSS0Jg+mi5RVWAaAj5DAh9lIiHR+0+fOGsvuQ3hDy5+xq0KlijB
PMFsUeYiK7x8774hlrSAXYZqvzFkbfDRkyD9O0PWABI080RYEFv/FJ9ltii95uS8yDGp10WdkEG5
d3Zb4TUnwtBKf2vQh079XAjpQe39sNw+hZYKZ1LC6bUfMDFcQH4NBiuI0M19qrJ/g24AXGHVd8j9
+XBgAVo4wqeuXpibtPnokE/LlhhQvEeHbwnlKPjJDiZS2r3TtrO5ktW/+6A8QesV3R+Q1zNa5Snq
SrPjxyclD3OV93+mdPMjGGhdX+4w0AN9Kw/pppZqZS00pkXJtTvWxrhx0y0ixhcxbVqf1fRgnrfO
7R1o1y+Mi9UG3EoZ60akWz5WTGRWp7O3e4pwXUDn4oleRPVBRQe1MPNdkZayCEV2rJs7gKknbrED
bi+vW/YOkhaPqRkm0liAQV9HM5Kn2lmM9wV43pBjGq+/0zEGAWxPJ6nHXSGvDoNXGGE5R8b5EtJi
BOzT2UvbVULL3mLlYaBc4DPp38B/QI3+sBlgjU7LBA4XyxFsOCC/fiELQJZn3iABSN3xfcNOW+Aa
OzV8RXyZfh8WnOW1bZehbQMio5+Gz0QCax+LiIsqPzx+bPQqxVuB6jyU1J59VFYPN8Ya77sanndz
wF0TBf/HxwKvQFz4Xzc+eKE39La1T1HaLDA9DXTKbbLTRZZf/k4C0xYQW6gwvMYT2TetbjlvhG1j
d4h8DNk1A+f5BfGmbuRXezswm9HQVlTJY2plE272OpxkAsizNKGE+LDCMSL7evls4f1nDeG/8iZD
PHuVcjREfLN0Hf5jl2ssjTX/dq516ppkU1cVXHjZn1DZyIBq1ljq4kS/nxqMZSo9ZSDcmWo5R0Zm
o8Enx2vRw8otzY0Co9Qko55HOJMIFJky0LpUkn6PgV+b9U8I+mCrQsoqUWMHzQvkB5YUGlVLayMN
5FBB5JISmtB7PrCb0kVXLvaBcw+qoLD+g1AOo5G9ldX65Z5WkFBdpG+pdDWJoEVndm+jbTG/hSXm
u+zwnbbrDF14ioq0WiS+BquyT0y6wDTwT1kS5hR/WigtfPMblSE0/7a8XM6Ih7NrzQ1k891mrfky
JfYXzU4Qyhw81DsjcQsjemzNLtWJEEq5N9nvOgL+RJ3wYLJCMpGeaZWbTutVyQ9bryqwCKgrTn1a
Fomaeear4mMTWRf1ViKNjJNN5FhITo0m9nIaEiTtF2p4JXsIK/Hp2xucRJo02t6/mnan80K1iv7h
7dmo8snucS6e3wok6uXY2XI1ocMMkMZyQVTW+B7pQVuUtEhqWNAZdsIhla8pbfLMrcgZrdgNpyxU
JhyRF3jUFg2KOh1I8kFTkeMP4yDSZe2gWs4vkCOAJr06yGq3UOoAy1OMEHPVPYPflTGDu8H4Aclv
hL+ENmxqNatqCC4W9OY8Hfj95S/MG7RDGgm5jWb5A9Z7l+qSMWM4mLKg05pVt+4xrHXj/r2gAj5R
7Rmlk5SHo/iOeYVVx5znxWYhm1hgKM7nSdGrCtbsxQBGXyNy4oim8K4MppIsehJu5SnRR8izlnuL
on7xooYCaE06EslE/oHcSeA08KB6qXMxzcGLOPAomqtSDXwSK+03I+gfu5ucKWTLSkpGg9xDqlXF
fcLkgtZ3pe88N0IR3dc8a6/KaqA2NIZkOVCvUv8LN9IrKa5BPv6TcIN3yEbVRXRGEEemm75x+rd1
Yo9+lKoqk9S88KbiYOAQZ/q2XedyZ9QqLpLaVYSW1o2BWJF5J6MS8nyl8dCkUxvQKdd7BC3ku9EU
e7fBRe0ajMkFrPA5L2PIppXXyIKvt7nx9yXY02MHUYItsIQoTUyn6zIiOwjGbzNDy5kpgAH+bEFA
iqZHCiSeAH7qMQwpS2Kr/b4DUtfUarEO3QCwS4r4OohMOCU9RvQW3wZuhlxnhsUncqZCRgCPJq94
A5vLDVDGF5DRmDm7GpssFEufeMjSexwaoyU9Bg+qD0mv2GGPSEijDuSQCyS9bicMnl+71wkE4fsn
vJ7oKytndElP+B2dlnR2muwU3hED4IhYMWnTM6SJUjmWbQsA7pR/VyiiV2dwyBI6ICq7eJ+hxr6j
brGprDZCqLM4fRH21e+sg4I+cSjaudpgxUYN7mko+Qcgq9c5j0yZ5LXPIyFrdW7lSnGSPDxWYH2E
5kMmwlVeRBulhrn27lNtvK843mrcbM779L6khKT157KNcWiLt5xbOVw2lOhAVCsvUAeIS8nVRBpt
8quwpdhQ9i7zP5rMHBhaGTJJRftkDMhXxnAJwbkjWH06dLltuNI2hBF4TO9Dzv3tOBoqEsMWPUQA
Owyca+h/YYpqSj0wwDMEZPYXMWXuM23vjSG3XPHiWqYMi2OCuzZxwPUfUqNuaq5iNOjqba7hijZa
Vu3MvDZhXWnnBK5DZEHIfjzqaQV8VwGpHMkvh28kYSts//4y8JTRiOqmq/BQzwFZA1Z2ULqvmnCU
Pwu4uhzbchE8IIKzfW8J39Hu73SJ5046DJCAp/eYs3rNJja+l1GxqH4kYtOazkShGjHelgsXrlEw
dPQajd72A7J4ou/4MdheHHzWsc3e8sXndql6naxOICzp4CZ4Q9qV9k1dm8O3xdZzoDGMuF67jNsZ
zsiYM3kHbB72fhx9swNHCL9p2jjDGiIjObK0em3D9RSpIGfKUjb6nsHxhwkh88sKdIEhAEnCZEJX
sF5Y6MH93WskoeozIAIERHxF6Fytuvpqjx2PSl1RSXCk9ess++cDtYkonKFmtQYyCketL033JAzR
Agnsfe6IuqaCCk5RG9ShLlh5Z5VE/gFAkLSdXaq6U8vTD2RK5VrvOVfPESwXV84r8VQEjREh4l1C
Kr/gw5emczcB6nsU4SZDU7/BAyzTP1ZH9NJx1EHzKfDuSEiblYqVZESWg0681KfDWegIkOogdUbL
Di2Catc/5//2D0RP04MG7O5oCN3QrjKql0N/+QsP6aBU9RHsZzw1iKJA+gAC0s17BhyjH5sYddl/
4eo8RUn/OdEbR8vxcT1gBrxbB7QUToN/MT0suyyLsgp56kRACZKKrYE6LQE2gYqTCQSSi4QDokQ1
wi0BzcutDNsTifqMYYTJdE+CxrABtzZqAmgf26Hu7MvjUr8/psgnJgciEPp7pcXL04LtnVVpCSnW
iztjIBx535Dw2Fxl1CA4zAf0oLngSTeyQijkljM5t2/4AwNX2owXe7OMJPX24gHsqL+zxln4OMU1
eozozjoqUGfvbrf6r7l6YRR8XS8kFP7yvXDpSvdwoXnwUOSiforyVh76jG2EyKhI1MYr9TjrYnjq
bRWICs5js1TUFwHABa4S7ZoU9QnhGrET3qP0qa8RpsBxcdm92PYZ1jlplBxqXemgXR8VbncAD/3z
pEKelc9/PczMoNmy62FnMayJIfRvVPgehj7PcQ5/82zXzRF7tBHOkGrgaCXUdwaSir5AYm2GPNz4
nWoTyke88BZsQ1gDOADvq7+ANGpOpZIW9OmTx1vTxYHwZRwkI5zXrCysloJ6kn4fiCpln0vjE4KJ
+m99k2XT3ppG2HoxQ1zShEhOzzsDUih9yZPh9mWfVG3R4wSLHFJG0emv80euUlqIoEjHVWUleBHe
JVnzwg69adY1TfSpst9dcbXVwHm4QahwUWgt8e/Xg8A7lf7gvNI7GoaBUNv4H27ij1I66c4efD2D
JRdwgW9IcMkP4hx74aveOabm/y7g+ss6YsbCsNRg0DveQFI7FLlqBFSf9c1nWbBIrJ0V3rEatSs1
v2eLzOLcCVgI0S1x/xWxhiH7EKpVR/nxSfrY1Yqp9lI+X70HWyteFkCFYBIkqTqBtc4RM98HJEwH
ovgwhAB1IzM935Lf/y1u+R8KS3YPi8NYzx8Edt3/V1aVmVGwAJ3tqKk4IpLIa38rxeVJ8+H7/5/b
BviZu1Bwa/Ch8ZXzibB8ogN2JsOtZRHtrV8hVb02dvcXyF2jQimNoFCROZwielTJ5M50IZVnD2Dx
qpbMrq68lG/WQZ0XJOlaEDgAg7ny50ly7qfquWNdObIFLyvCUG80TntDuUXL8hMv/NvJPlKuQ6S2
lHoQBZor0pzVkd3etrE47vlFhhkJ77arAzPpAbbJEXl6mX1g1D5x5NPNVcBN44oEEUcj65O4iN/c
zPXOc9XT9rjGRt0fyS/v+e5JCaH4LO40bHcQBjuvejEMcNGt0T2+15bq7isCW3vzVeI6eNfFxYrF
366XPYFv0LNWy2hq0t98lKmYFrLcffNv7Euk29PWrKWo17RgdElGJpGp4b0GJeyMF639ezVL/w/8
rsnm2kI2z0DFNcmdDNBGP+Z+WYoDSCI6q7XY7zUIc/KJ1CQHQ2MPDN+VPNk7WzX2MBtWacl7mApQ
+T/0sis5VZHE8X3FXi1JPIF10/bile/ddBqq5aVntQ464lY+89Xl1fse9kOcHGAjp1bTnilHaZmQ
ezeOKkmGhocY1qpkQ1UMlHnfxAsGhIbPZtpDIAKJf6ql+YvRBCqXtJTGQoXT8TaCmCR0SoTMW6IR
2xOwvpZkWNpOgUQJgjN2DDkOjAFHEMajboQydATA5v/9xlR1aBwiSTims9OxhH3XKF9UABnP963X
uiT6tPIP2Fltj2ZV4IhZlE8CTPEvenHuqgqa+SfYglRIInfRtrLHeCfxLG6FHv4823cdMlmmt1wJ
LPZ1oJvv+lbZWOixJlscWS2+RnktcKxGLqqiN7ufDKSIm3z9momcAAgyFh8iWE2BmLFbAQgwj6V4
M5VfHWdtVX33ez+Qntk/oV3rMXI/1ZhD5cjyMzRho4aSzZeIMA25gjTXygqjPAsiRzZjknWEDTIk
BrDxaLNrHgvN+WR/SfhUmumENykBCqEJ2STxIlH26BvXseKw871Ak22dYT0rrGFQfsekySuF5U2U
OEg4CNYgITVrE0yCYF46tX8CpnRa8AFYEYhgHdAo9SAdZMDKlPMTbHD7hRYYCfsVMFS5iK0ERwz+
umL/iSeU3qhS2uvF/bGIA8Xwr9E+QTyWe7EGv3p0WPQ/RxYzB/j7sNA83A4an6A3iNZJlGO/okRk
kWqYT3ZBOhfXEkvx2jJPosDV6279BWgqCqbd3W0krxzPrBDxYZPQI/aO5JW8jNPT4hOxzc7MdMWN
7CcPQupqbT6udyQZDrewfnV7rimHClOYz0QUShclr2hEkMkP7muxcV/wDSFQImooKEiU8KU/tp27
lYevSDrY5DZwfyVYBoyHzW1DEgiKUBTIWL4yrAPVKtr3vSe5ZBDT+JX5TmMuiW5EWkmTM+LIa1Kx
JH/GeLbXdkoZCyBGNacuGpo4JqEvq9j6D9ImHYxBYUpSE+mfMFQB2i9eYGtILxrueh1a7GLN4Gxo
B/Nu9Hw3bgN/gMjBRkvfOxMDeL64WUKydeN89GxNRP7xEX5KA1al0bKhbPIXqXPul0dxrN4lNty/
M2P9qF4CtBORyKQgsh7/gyTPJH8vuOfV1i1tr6Lg3GmSOeKtfqZ/3OHVavJxU9QWr+rDFIGnUQ8F
EBbD3gnQNFm0dIEOaqmOnBGnDaALvGTSFuk7FH1gxjwMn85PxscjDb1yMZdHUx1NREvwLG8y2PRM
tGraV6JB+5oMJB7Jf+a1FLMOJ8M+Qes58BOKn65RR3QWCuq0KsM1LpeOrWCy1tAC/HPWQm67ShqZ
I0lWRc+gCY2tpC/fYLynuBEjGOfFNqcSZcnoz4zgPKionzuCUsmWzphK3l1Nro1WntMISFvVrViI
4VCVg/QbVQOoVji93itWw9AwkPZKqcTuvJOalq17deL5dygr1Ivl9kALO1tmWCmP/zecKZhM6vo3
eWSVDGwbJnPwsWEX/KNJ+MdYikcU8ZNMtl3UYIXb8XyJt0dSR2U18crj3tr97/fJVQq2+5JhG3I5
NFYV2rNS7x5GZAAh9SIe+H5bLh21DHecCQUfsa5vl4WUvmIQbw5nXUp+N9QA9u0nLl/yrTRpTWIH
X3HOSX8EPvmt/rHPSlPpTVvV+GEyggqdYPX1lVo90K+SJyVQ/+QvFjyjf7VTDHg1PdPRqtDwdpdw
u4zh9Vj0/MDpDge8jkQOiUHEScNi5BX+FqXAI+4EvMPBPErj52xaxU19s74jQr8BI03KtLpFV2ib
rMb3d8jsQOIHsa7JLh7Io14eVigMZ3wQCXqLDu2WesDDghS46oXOnuvCeXVy0dM9TRra+b7FnGn8
jCb2Ig98+kAsFZMPpCKCSS3ipcSpID2StebH3vmdW1QL4ZbJM6Qo9jqlYpHLWB2Ucwah64inOMm2
knC7vpvxvj+k5pdWH0yUiu+IOyFW4DPrx8hEqJ0WvfjhX2bW0v/N8mdQpUoBE9u5i8NoNQ/CMH2u
21GV1Y7rB8JtbMS0PFRr3u0VkrlBS7/8dfHW1v6yF67XhS2l9tWohjdg6VGosxoLQ2rrbPEEOZqh
pUEPCDmfXjLqxWYhlurKaCGofJBfnwi1FMPp9bo+aiuplJW1wvW74CZtSntRibtzLEDCBcBGCEhL
D5aWNdL/6wXCfuv1H3FFki30XnvGlu23ZmADOYdEk1Zfthoh5YXBhFHbIMCow4bJc43td46gGLpd
Tji70Qy4KVzbTv4+4TMwfP4DXaD8whxHcSvQQXBgvmnHKvc0JJsNsGSNNhf6ZOBLgN/KSPy0g2DL
914j++f+O838Yqda+LJ2+Nm62ePCYmZv5YDWoJmADm1tOmGngY1fDdxL29gMdy9NEndgKkdR9Ivl
/ttaJso0bAcwqPPWX4ZvNTYVz0YVmjZZSIhzvSxyyvqeHWq8VRyz/hBlrUD9BoA2viSRDDzSktJC
5ia1Vtz6urN0qvakbcyJz1P3boBKAA/ph5W9yGljnwCl71owV3xQeq5E9VnvS0HpHbRszoJTxEBw
2TQMK9Vjap4I/PTNbbb8sgfW6gE6co5bSvP2/BhO4soOKGYgRBaTMAt9X9So1Mj7r0Rd+pkKv6KE
XUMlid9rnW0dQvX2Ag6pYse3A1Oj6a3v0WU+QYSZQfdpwCtYj6K6ypFMQwhMQoR96LdEK7pkZlhq
sgQB9zHz4vKAZYP3gmnNHDrf3eyKwcpASJgcUdk2a+xpFxwb4NYquDC+SUkAWvPg0LBYhj1YbrmC
fm0qFVm1sGncq26rFwgnWHu9W7FjRvvqsQcS2sqkiejBi9oUJEVQA6IV+tDaRSZy6H8tddpMAk7V
bpp20RJt1dJTAfzUpXbVF9dCp9gcMmeuTp4PmUCx7jX6uVpvFG/nFurz2NSE+OmYvhsFEiYQ+uHo
+45EhscpgWa2JOUkg/3PAtSprYw9QXK/zU1D3eJF8trTB1+0QOkKKFIeK8z/eD7NicfkAWF5pf5q
6RVulhMqqmTNgRgn9JphDWHUBfIiSj7fXvJoq3FF/nz/NmcuLLC1vQDfkBkWnrRUoRw9jBFhBaX3
mvKQoTpNPKOs82PQ49FlP/x9tnCU/C/fOWKvqN7SQOnfHGkC77yu6eY7U32WV+9yidl+26DVN96j
VkFpaFuSmnMKFN1YJF+ZaGALmjduV9yhjeiZFccGatz18IEA2eJbAkUBRCj3j8Pg72kQiU3twcjH
cRKLPFHcvqJmdsBwy7e2s1QeYGWAKjMEDB2J0BLhDrjLaDjwqnGWw9i+yyAGWehqDDjiT6IJ61nY
jJ3kCmIOxLIA4MCm2/BCrb7Z6HLOmb+TPwcljd9uk/xxBXcqgIspTwt5OWQzjK62HasX7Yxl/dKZ
kVN8is7jy9BFapWeWm20KV/70Df0+nFrg8ewrBIS8u+lG1sDIe0qECs9PUw9rku37P0NsXaAqGGt
kLlFbam0vlxx0zMlDH8bX1Kw7EpRcaKznSDHlC5uh7Tbbq8KwvhGHnOsosGc1B99xxepWeeNMJYt
JOdxcUnjMDaPnJ6bpFtseZ2ycfizF+UA5C4toH02pGTzPuFSxZjE4uIOt3Cr4Jh4iftX0zWVuuuE
Gedohl8HBny3kPJ0mD4zaKWGAM4tNPYM7lrLqja61ip2PmYopp0FQ2FfUHtSs4t3aitFbEWrDhFw
iM6ybMQUW9X8o7GRmaMeWyTUzD67AwioekPlDw6APqamOR9RmD9pnOD3C1CkDmvsLA4qav7ait+s
svtsRmZJI1u2WkLU//2aRJrjgIV43LwnzKByl8yqZqoTZDHMU3sVpBNy/Tgi4E2C3Rs01JnzMo/2
h6j4o/CxbPq1+SS1CJsVDCkkogKogC52V9+WkCP2XYyIPolY/LnaxNy2+zNfD68c55WXesHeFWSW
tL/AvvuqUt+wrXeVvfKzHj5kGtniY4ctBpcvc8Rz352URV/WbJ0QM6OXXGAQGzKEKX5Fuh5YDCs6
vei7C5T99hpizTPxrR9aRmPYsOeUoEq1w5i5fimRlXTQza7WOQETelC9HGc3oIcq1ql5Jaw9vau1
m902cKfNHE+yX422uTdaFPZwdGfg6I7tq77PRLPhfu7djKQbQFcBxrR+HNmOD3QrPtyAsvqfRDsb
2UluLnRRkS8eL3E3JflzM/fagVsiOFmVvKmRjDVRf6fnhz1HhTxks2IfEqMXMoMrbfvszh8JXLoz
6FCtARYGFgXb4xnwEju/Pgr9MSbgOC7HnXUpARDKCoytvwe+Xpxc7VAY7BhTzzYo3BxB9kQBRxd/
2IyyRMBLfxry/VJDeli7fpBsK6yX7id+p5DMDTMaXkIMCKqR3AT3KukekkNnuPoKH3vPl9hYDDGQ
yur+7IY7ZkewC6KzG0713dMjKNY5pVxUPtqGgt/OVgjK2Sbqs4LhRsUfiQcqXWZh6MiNF6FRmi47
ZcaED2CXNUuVnK8YmKycI8hpF9GjgRY2XZx2VOfezTS78UaxA8MZvezgn6+ei46TlhLTDbK8tZWz
rGyNCZFORns0zZ20rxiebje56GXA0etPgPr+A54pJ5UJoKU1QE4Zm7BL1rfIcSDmdoV6KJH4KJOj
oItvdCvWckvVYi4Gl0EyaZ7AH8tnrFst1tTxe1GppD+tmZeCWFpAriH1/bM/3OUGOTdXMNkuTB2x
kguqX6gAbBLSc50zNseu42Q/WD2CyoWGRUXXrSf/eoUrlmdRjovTJ+MYy0Qo1vcgrYp9LEma/4gd
3W2wVHF1ied7p60/edaoAw9nzVM5xjpRXbNWU+qzDnrLdjCkV3hm4PJpgBTIiAX0+iFiCVS+7tum
wp9UsAuIBELJsSw3RD/dW464WW1sKz9poydcrULz6TQmg/w5EqOsfDCP3u1KB3LXc2fEXWTrmNM0
gztUGLNFi0us8UOn26sSBrbW+94FDo/UTo3DEEXqMzvp/PqlsXDP7JQqylI5Smb0lwgtuNqwQZI9
oepGhiKIjlQfehC59uHx+50msV5JoGfJme3NhAVUl/G+g3wcdThWjH6sd0a19h0RKIa5Ya6QIGMi
/n6icValcB665L9nGuVMvKFapJtOiX8HYjToEUj2aGRtbkeBzlkGSvxftsqjYR2ad/EL1Jvjf9Fd
DLZ57cVMjsheGR4pGX6Cc3r4vfH6Uh3kUxPvgst2vk3QnZmr61D4Soc9mu/ldAa1O57ru+8KGL2+
xjp2n5H54GH/QFTvgEImBc/OEE+leKxkOJTO9oJCN+cQb1JBjK0zLlFxn7YnP3uSND0GJbyxfY/e
RROi7Rp5Lt8elOs3yCMK/RaGB0B1GQmTVVVOtNL+DzLXGEbcGO5EGFFgTfYbGrbpuGQPvJc5VDQk
MgQl8M81uoueiprkQtzWTmvfcuaYJwAaTm5rsU5WBT6QlRvkA+ordAsajla2gNCTfa5ya6Gsnaiq
fz7TUsglwO/UCANOSj0MJFo4ODHwM90xPActXLAdTxUJrukWwLOOkhoxWfI28gjF3RTAqgU2G3kL
FlmQzDzGtS7C75yuyhiXNlUz/yqLeUgiLdF6vW7P1tF9ckmn+Vn0BqtgI0il0Ykw0qbcLb6tuePf
aYFGG88dI0IOKoSOEheLx+o79Cnl1sVrddq2jdXugCmZMFzmiIayLlgFeo3D34lA5Nh90FlfKcDx
QzVuOsHevndZ9SBNwO5LWdehR8dmM2xpupsUODVh5oHsGLceyAZ/I9l2NDcssTADmV8D+8D5bgEO
TZXIZUan7pv7LvkX9gmcQw3z6tMcmJBk9wuXFZCAoyB9m1QIN6pnPXrVBH2FDe+xJCOaIMSdF1ul
9jfRXATlr3m2nmdG6/UoVYCpLeWyxrD0nB79wuVSx2d71jG8faVvy/eZRlZyuNjIeLwIFpv1xREb
jjY28mQQctbOdUpn9Uh8rF8YFi4WYHFCT6erucC8K+X3i2FAXJkf8tfOO8UX/UHzcVLSoaSHIiLF
SjH9JEiMieqBpIN6q5GaVC1nmmkMFyryIAIpkGwFTpq+ITh+oZ3c43mipjq5u2ILenkeB1KJ65Kg
O0zEo5LkR6s1ugxpIKcyQYK1GQBEyTWuCjpI5in7C6pSaXjhxjnWrnP5hxTaaYlpT9VKGe1XS9or
EhV7m7shez8F/Vi0JEe1hSNe4Qn05HeNSipuA6c/sI0br48o8NwT8x2aGtgJoCqHJao6SxQtqDki
FSz+0SGOYZQymo2vl20DtygtFWjDb8ISqmtTTq/cAKCftSOlH/Ie3/vLYjgjuzPb9RxpioP9+/xs
Vn/6kZBj8RIXOIq5dY9Rruc/pKwmnzGN8+3J9MXI0dLSvSDGRQyK3OHZ4XhzPlDIBwMtsbQe48W7
X4UZGGQSYMCoHLtKfnnZ9mo9eSIO7YOXsIMX7qPQ0a1i5URVr0qzkPzW4BvzIHlX2C/mDrZq+fWM
S3s2RcSMbsWd7bO0RPZxK/l4XVzrZ3A1ubrf7JqbFe9bNaqlWccMxZY4ef8SHrK9F+vUd4CrhQMW
qC0GqBiDm8rDucfGao1ZSJakGWxB4LGi/WWUypvcySIoabEH0pv0QHshMRuPPBITNGeqb2rCF9Ma
exrNhtDBzmQjIkVm23HgUguX1d+NbRCi+ojnxnHJvzZW7Ds/28sna9CDzgjUTH0KkERkA0JJbnGs
26lmzGdv54wXyvXU8pB5ZSh4P37NW/K5GtbGvdBZcX3e9auZcUZncJAT/59xjhKy0BqizWvbkGki
UYw164iZoTIuakZzgsB3YDXoW8DdDpSDUON54PlxnPpXyaSodMK2D5lwci/cZ8+K7kdhsg1zGaTd
gftEKNWvIGVjGpbxoQ7/s1+mE3FbjIvw8fey1DkdyU1sODPjObUWMXNcZuBVDhBMUXlq5sFZDyKp
zk2eazepnyxSTF+sroNogODWzo7lr4hBNODxItcTN9YlN/luYM7CZTZ0mXvd42gSVUDaJCSknARV
CDFqoGxEx20tcGDvKJL6atcQaAkUh6wTZVCp8+gTRfQoc35zPCzjQ30pIW5DGwQCx62nSHBzFiNJ
TlOImM6R6q1R/uWPp6pD9EfJJO4nAX00fBwsnFJ3qq9ZbtDF6MZ3fAkO/yYihzt/mZs2PwoONYH1
WyNDV2k1fwJNOMY+AGn0WvS8Glu5eSKC9enGw1SNTIi1zV0g+DFJJZwtWVkk5ydW6YLe5RUCtVoi
9ZvTYjyERfGMGnwjDy0oRgvBeBGR7Fwg1M4F8WPzosix4oORDUJXCjvAZRN0/3K4hK66h2otRuTM
rNHZV7Z2hHEOtOb1TyzZZaCHCKhuAXNkd4Y3LM56ARFFWycR661OEad47KMsMeWuySH59/o+X/bJ
iHfzg2VcqxlKaEV+6q2lMzM6dH2Qf6wh5MiV+tlLO4MtzofMeKSMVKHDmbX8gFsUZ3bbrbszpRi/
PFNq94OB9OHOWGth/5D1JrJ8Wel7XbY1KQgzTQwYVP1HCMuSODRqyTYztR7cqH0m+a9tjfK/M/lK
Jd8lHYrbgzyAE9QKgte0Dijit1P5oHhcdGJG/AFeCBKraiymHYFdXPwrrDjepes1r+E+sx7mKfn5
4JRjOd6BEEiIA1+MVIgPfkv4lZfElUpgLcgYRMrty4g1eF//Af4ubHKW+kpSsew6Xr8UoT0udXv8
or7/EVMQ4u2uuVHslj4xCsDnqmHxSOm3yIiGqrsWZES2aHxV0R8f+d0nw/WZHfq0e3ecQbGz5VZB
joiiaJoWjQ3S0lSdHP3sU6kf2KDOIKrsJ6VrfrbFqxLoNnhRwPERe9mS/LqMlYdMYPoLRDNUQ6lC
UIrywd0pq4PALqTx3+03Zm+CGHKqI6skXP0dV666naDJHNvwnXR1gT768VDByJ7pLYEGwaZfM6x9
50OYMZ2pr1b4lP6EjEApLLSZf1GibR3CR0tLmrZcXo+UDnNth7N1FfvWeaxcJFn/cC3t0xf2P/eG
kJVyrfM9qqkgpJuyY+zZoRqoJG2r3n8z1Rpkx1tSJc/FZ5dJHM4HgYbuPETQYw1W5Cu/yNP5cHee
RxSrK/Z48wDtR7RSoe5+WriE65ZmkKPYEGCtRj2HIROjOMKZ+GGPSQsEyqdBpa6q/MtFUkXvW8Zz
sK8lWFhsOH7BSc8iAkEJ+46e8YCpBD6UsBAPr2ktpt1AM63fuRsR6wmZUD3ono4eeS0g5Qycv9Mt
Jwi34FoGvg4cDwbj2qP2pYJw/RlUZsIut5PDGstVMrBVbnPImgY/bq/42JCQzNBORfXIudc5fsJY
nHLAgc9aaPnVSaC+V6XdXyale5Dc2JG+QxE62wupRTCnhI9CEhr6Kb+wAXDCrPZCf2UnbkIGJOc1
eLK+7r7A5Ns/PxEAYCC6yPDZkIL5ZH+9guhV1r7wyWI1pZ0T7AJDSFCyEpJd211cttJ4a+kkjl+z
jEJ9FWNMp6kk7gzk6NSOLXOYhrQnigFwUL7OxIwZ4DPyGMQ0+0CC/TZ61EtvOEjxnbFeSr4i0s3i
9B1sa4WOlcNp3D6kCDBdEPLPtkgDMvpw/9t1HhOjBwEXQdzFUXipTJYLKYnnXWkcDjFPBv7P6tZ7
5yKKpSfjJeyHXIIE5xPSrw2o1bcQnqIwg++YDEU2RsqURYjAH5kc9UTdXX+PoIptDGcrvq+ueGiA
4Z6VOMcJXuYkfOyZA2VkKEYKQ0TjUNTNBUN9v9lqCCcmEhVDXJHiwHzzKvx6pzhEfClSy2ep+e9y
1ePeQseMLe8vbH1CD7KdI6r2+thFwglKywmWQj7tshTvGsgQqHIhiE7OajfWOnxiTUzltaQdUwRR
JC2yAayHQvf49UCpNWsHWHh/D6qA/9hph3mDm2xJGCfI2VMtZwJbiQwLJxTkviwoATH+SWkBZS1o
yU4Y8z29a/OMzbZZO/4FvXKHns+muwrN0MnZtcD+dkLfhHh5FFJ0d6QVHwcuSAiY7MaV1nFG8yvc
vaRmZMT8qnrIU8gyMY5PzFwjRhmLxhzu4xUZdYL7D/DKksgYXPXK4InAdI+wm0oQNszBpSpoZNG8
nd/oy9AsI/+stDZjoRPiuypdxBVC2aLz2Axu5YV89AW5sAuMCS5tqA2qxDRwPINQK6mmspJXI52k
lQ4++7bpczxj8blC6GBWt59EULgu7UBCkAgD6mgthTgyYry9Finh+xuoAQH9vBws8XOh9b7bQuWM
eY/aCgf10WeKdi8Wrw+cFpYpgqcgyxVc/wOprumG2O6NmjKGRjxc0xvvhhnYwKM+PTIzIyCXACwi
L2LlWq1gtbSWFAmkCT1GzIcHE75pmUJSB4jJ292aDmXCJfhf6+AlCHkw03VO1KS8dhj9t2xd8QDe
cdNyXuRLbQuoAbQeEKYLfOzbsSCenzRc+p45tSuxcZqXSrtWQujBk+EOxfOiant5lXTmz2C7vmVs
KZK470gptgX4R19ia40BG04btWmPJDyjDcAoFoVHx9pMjyPXglurHQ7XHOF77OCHEkGzqG6uQYwV
Nxrh4PGdqdKHMidjZy9UBOwwKL1wnBoZJRVpONS8N7aq2cWeKqbK9RiDQOriUI+fTCD8dAs0ipmO
VbG5D5ZhWeWzWTR2zV2cpqnCXx/JUSevqGwPEYnm5xgl34R7vjtQnxkPwKEvwQfyX7cgvmZlJzSm
UkDy8oOQbbJ67kDQ5dsRRLqgwLu4p1yZie8XbjvoNemWHgk9lylpAXrLVSP0WASrMnkgjGRbRIbq
rEftnkWhqWvIvZ9zTt11BBulN8LDP/Vww18MkjjCHW1XS0MONCqq8Ca0rcLXzSAN2deQxJmsmVLj
MZ3QPSBWxV4p4rSc+x1Sj2y74NNdGsWOF8XcOOJ0EMWr/lsDUNenmK1IfZ+7/W3eqkWqE7AFuKaD
ZOTa+sc+zLsx0mnBp3QAt9FiUJBTM5+OaGeGzfciBNw9RIqSeIpzWsskrVbv4+E3DGE1D5/7PsUF
G6wgjvBaQ3C9udPnXYl+MCNMUGhv+0NKePKDFU+yKzrR/NcyrUt82NyGQhnPTFIzFTur/2Cyh+0M
Vaxyn/EkaUc0r8AOW/mPccHMJ8BcxViWIXeZqmFO0z/yj/JR2a1QpzMqc3et/mOeAuyLNuaT9c86
R6teVpP7gQ2DrrBpp5z14Fpag1Hgzhg2YXavnLeryB5NMkiQZj/xrRNtVUCz2nUKyegEM14iPSVV
kw1ddMX+J74tIn3qHwwVWcEqCkz+03lAlpL08cMVaAplGshAZ1RdkGGsEy/uuI2tpHKcciyv3TfL
STYJhk1XUp5SJnjVChx6YSFX391LWFfJ7lg4f8zTuFn+TJfWlElkpkIV64v7RqJzxyXMO3ySqZMu
7KMGqPTks70bL/uGNXAAHSI/Uw0JK3vFaDQiPXNPnmmebyhF4/I2HDLlcIxZoNUSNy32Gqltc+5G
OaO5gOCnDNCA3fawgLJ3WIx+4Dhsgr8VLRPCo1LVSmrdn/f7ywad2k188JSAICN1Ja/Qcdip5j1d
dMgvkO187oI1NqDJVUbdEL2BWlMgYGwbFPhiIPQBIDaBD633gUFtoNdBG+CCjmasejgQ2d6g5XQZ
zkgKk5cmmGLLspe4ZDLIKgiswbNv/fMaa7Gtq25FVwJhiaSOZog70Ace2gjPBeRa63cax/OpMp17
4wvJHn9CcwEufU5SAp86yqAOmUnxKnTnDrPTxTT49gBsjM7mKEXuhDWstBPZStV4g6sPa8GhSZKT
QjJ6lmbz/xSLD1gSJ+Q6hq+3GF1rqb1tSal/LF07f0Q/jLJlVMwFWQyVh/k1Y7MStue1MZIVxT9/
uj8cx8jeL2cnufkkk9OTHJOaM64o19eaG6qd8hIRtnQgZjGsPFE3VgWzzDUrnhiY22dKpBFLuWYX
PUBLse8A1HRSOw6zvkcr2cTwhOHSur91+SWj8cLaV60iFjpGhpMejKD3CBs3mKO3fNVq7p7tTPFx
cvM6PKYT1edCPf5uWtb2WdDHAl5qISCYoek03MWqJCJUW1nlMq9OVIXU0dL1dWNc5c/CHIyxonuO
AAQUOyYVRl1Q41i+4EZvfQguUPyUpsggX2JYv+kEwfRh6NANNtrcglATFwgP/3qx9oePvMAaXdMS
ofuSNUDDHmG1SFMzJG/amQWxJtVFvZpfV/bDC0jOnC/wMAkvWlWBgXF5NsI6R+juHrCwh4/lfxqZ
thMLebpCQFF9d5D5DFV8C7QLwNsHhMLYiVwxjRv9K7G8z+UeSUxD/mOEH8daZK/Rr5AhxWi4sqb4
XN+Vl/UtLo6FxKLBa+2CWDPQ/jzso9Qrmd3UZYEL+vW5ET/g5C330xAXrzilauOld+hU/KC6pCle
Nlg+Hqjpa3dT4N0c7oLrRWihVPovwQZcbMSRdou+glNVNAvW7FHQOo+O/t5tS//BlZ4MSnXwTZ06
0ocoKrL7WWqOsawvnB3JGIdFGtD08F31hAlUKIAFyOwyEh5p/y38tkjWPvhMAcqlwxd7Djb0VBhs
cNpYfMMpM0w1TroBKju+ITxNOsRtya+rKUdbi+SRafGqPkB8et7cz9rJucq4ks2BcOCUPiMhzf41
EzbfsLUAXUM5bgzzzxsIVt2nsNPqkFvcJUt9xyoE8d3sI49Jd+XgGl8j4vLLCBnYu4RNga5+YuCm
KWURzck3Fqv96E3gkMJ/7LKoaATloVOecyymp1o485q+Obi0qwN/Fx3bFua+/JRDi3gAgqcGxR/J
IsOjG4CtW/yVmCSYoMHONyrxiLDOJZtt5hq89qDCnFAibnsewpRmOlZA81nLTM2kK97U2QwnYi0e
uLhzBJkd+Di5Su5IcuU4RUinMDKPsP3PmT/snZK0Dp/LBsPu5EkGhGzU9vMyaFuoUur7ElfDTx7j
0P7FSyhVIuuCXqpzHmUGInafhIaCK5n0j52izXC9lsXf0SZ2D8Kw7IBY6rC2TQy2TFhCnOeTYpSA
sSX5jwwEY8WoVEfMFXeH9VDPQ49sN2XKFrBVrOd9I+Ji3rsy9ckRzZrZHhZ3tHOyb+mwz6TZjxdK
6RHW127xNX28nSDR0QpTlOISl120VRQcUhEP5OJmlMtIXxnp67dpJEZO1IXJv3hCOW45mJ9JLrCP
aE7mrTTdyQ/NOFDeiaZixqxM0w6c/mkKSS0Or5UloSl4qKq4YkvjG9Q73LcujAETDTU0tVZrjpgK
TMiqQOojpQO5SK3L+HziwvRFqJPIIE50OOlxsy9fx7ZS+MZqZgtKFJu6hP05BJeej0qeODGSHT1F
uHyVzMPP8KBTdejNqiezSd8/AsneX5/cmqpQiQziluSiu1rgxOSO2RPvwQZYxR9b6+y5o1qH5XP1
rUVdTIQSyrtsna1o0MK8Zb1ewpBNcMrUmC1jTuMG8Dhy4rVArbHx/q5IFBuBpJEn64YYQNK/Fkbs
FiZ5vzBavKUX/UDLju3tcwcllbpwV1UERVf4Nj9GqgC3mM8elyBOOQDk6muMakitzDy0uEBDTNC8
UNtXbRyr822zrbKn6BhoTulC1yQpWa+CxALWyz4jgO3TihoOPz1+lJAiupk5us4T8u4T5dTmGmbX
Slv3Udvm9pu4t4G5ot74yn+O2mdWXtjhwN6XSYrJTfDGp/mUN79GoEgwTMqodoa5hZlOPqhrnrlj
Vme/V+zYw0duSNrC8omtXqlBDVoDjqp9JigKV9Zunz8mmGuoR93yf6dwZpx+GTnAyeEPKC1qw9M3
sfsqedxob1oANIT577ChG/0Wegz11qGOTXGh98kBhnXVYkijBl52Yq4NbkGeUkBUOH0VhK0aq/G4
WgKRWjMGr45S3nzn8z7MjCSpk5Pt7DvR220U/C9xPdjF5g4594A36vxnmfRqBVhfD0IUqyQPrrYj
hTXCdBzKNxAUuOsn3XrkP+1Ahh0kMPwqFZPYpsup5BnmKYeB7jS11GFevE/1ZFokG591v9xjNcvQ
hgTHni17AeczHRHoZoKabLpu4QoOeR6fmbz3HWoaqQHPfdACFWXmFyfabbA/MABWeHxmeXv8TwOx
/vxtkJlXivGE+te/E6+34R7hBXImL9JRyvlI6zNOKsYAnIMxnQRiwwNMCmRmh4ILiBVEtf6cr0I6
YUGHHdkfveynN/IRK3avG6hAbK0NB4pVD1cszzLde3AxbJ4a5W7v0W4JJhro3L1+zzRd/ZbesdW+
YhCyf/p+k0MTx86DDxiN/9YpE/kylomgZKnHx+JMSxbYcQ6mepNCpWBBOq16QKGQS8e88bWO3H3K
qiDZSR2qR5ZiwWTSPp7UF+fSl3Jgej2h7NyuRQbzHogr4C9tflPQIKOjKBvMhFqOwxcY6us031zZ
edJZKsWgojPDrBr+UBeaFiC5GMPXnYWMdKAoHyB9uTiwSeJFHojyRz5PKcGcIDKLwMOkl9rSOrxm
4s4FYAgy/umnkJi6CWUARctpJDCNsW0KyhZ1SxlIcF1TEvU1Bu46xqq9i/aRREC7RckRBsVLQkZt
fC+2m3OkOKUhdDf6vij7YIFYN1ihXmoFEBGqwcytGMGZU8rzwaEY/Omn2WBxyCevIjn/ECVn4pbo
RlJqrjYjyaECuSkCX36xYBwcrpMSl9EUSW1Eyj/ukoIHFYG9hSR0SbMUIuewAWPLx57qXYb/hubX
mU/s6aQ5wsMK8ItK7x3b9i3Wqn5fGoPxfyRpp56QrTIBaYLa2HwNWIqMqkf08kdWXinN9Yj9PNKz
Pgd/GeabT9hKMTKng0M9gtgU1N2m0r4NL27lLQVK7xf3GOG1smO7kr1YNlk7UyigTj2hBNh/Yqw+
4926nVLl5++SgktJJbuAOfoFA0381p9F5qbD5H3BRp4Zo6oLjObBhw0J4g+nr1FC0+w+0/SOyLXZ
VmjfXI4nxRBrN7QTJFWwkd3x7rJ7xe6lNY7ZI0FCUOpdQBU0w8GiNoojVehGwtRTKcMY11sER7C7
sk+fIR+t42yFTcp2JCU2qgnfbqDZeF8t4MSLUl/9mmkUDZ4mawZP3IjAegprlvpvgSTESxpDcyKg
bRWwGX9/MTlhmooI6TXvXiN8HlWc1tHXurwZSk16oxjlJAxGOLVa+EtBOUUZY0NgSzjciS20EpZV
UKeCBZVkkK+c/E+Cw2u5JIAM38csiU10Ww26fl0DDOXH+vIKu41h3UJk79JeL+fYkHKJQ0gjBj59
MvVet+z7Zgf8oNkG3ZsMqzF7u5kFiE6FHr/YqOeA5oQIgG/XqzrY3hC1mY61YXTsuVo8V2f10/To
NTcbH4u/LnJ0focnqw5+PjUMfT6/N18qjXYrVjL8WRDK0lX2VX4FjSplMYtcZi6YWbkS3W6kmVZG
UQAhf4kvIPnCNjQTGCRg77ZXKbKLYtgEbeZsZnguzICYmLZKcIRhoeKKan5UeCUhb4l9F2u7OvqT
H6VTtO1DkexHIP1W8IGOnHV2tucS8mHFmM7X1UgBET+AvBePSNE2qXPQvSK2TC1E5HKAe5bpZyfa
dCC2CYlePcI9bL8VMPRGWkd0xemQRv4+/CBXo/Ws8vDmoX37qsTa21vHtvX4BtgAldX2fXwkO9DT
HGI+KfmDD/3fUwW6IlSjjthahaThcTtne90EaJnpnSvQXfM4Mqmlf/bUK5lk0RT82e2t5XQvQ6s5
2sjd7fEgNo1d9aC2yFiNerMW7qQo0m/F9ZoaQMr0iXKr2tweI8LEatIkj6jdvFitvBPEzS7llm+N
4sd8scySZViiue1maKPbdOOX2qySNw/ALkJIcAJ/E5gbSHl+i603SobO6rDqsIQINJ8LNJvvRIIy
r4M9hknsH3plztInxXT7YnE7NaQpTCpVTVmnHrweZzf1bYN07MRI0TgjbCDrEqqgmuOzHqcFJ6cZ
MOsPJZ9Vi/z5CCPorWx8N67c2X76w93br2wehubgnHr40sMh1zEHKO8XtOsii+NX8lSnDv4usW75
UTEuY+kozoNKvuRY+aRND6zAbGKw5CeyJnTwV7Acgulwll8/0LjYcDdSB8DRvSVLXgp19JvjiuV8
ciEDuA0k19YN2IxXtN+uqfSNJpr4Fbj7d78KvxKv8A9Wb8AqOWb9wtiKuIcyJrNgY0lMR8wPJ0vT
BgoejdCkLRzOx9ApRlon1cZocMFi2AaGQ98Uoj336D9taUqdMnfqZ7+TGWz/infM/Vk42+R44zn2
8pmbqKFiRy8xrlLLEKiqAibPxIf1udrtopKNC2AW4BAUx97FNLNpY716QiDjyLFUs+0wED8m5FyE
QANdRmnlbTQiT9B6oKT/xcKIQaxB9nNiIiinRq75h6Gio+S6SS02t10PWTuWGyo5onVjVvUoAbY7
USIt0FRm+aSpxDSPRVPvg7XU12HgJfF/QvnVAiByw29/uBBdR0t5izcsDyvH0BMIAr8uO6SmVdLy
SHMKuQVrSTefj48T1Wc6KUWKh16CqCqI/r6/cpKVLE8fuZ+Uk2Q/ltOeccT3BLu2hBS5nwf7U4Rn
WD/Pn37UNc4AXMi/A9JZtw8hTkTWpn3NdszO3wKpdNdC7umy7A13HaM8Td3nkQi3bhyW/JQK60H0
Q9YJdiFA2ogvYb5mjFvZPQIt80pw/iL+9kepejWgapVzQyWOk0E8VDzNmUyyWAMIQo50vrd4mbNp
J+9DE52BVVqRu+xGQ3cU3ojgmg1gNjiv2YDWSFoZLUS2t6IsKE9q4CM/5C4BZRlFw8m1q/D7zi63
ds5VZvmGryqEzbwtkfrmrV4SI/mwrourLYJH8eKB2gFyRZQaImPIG+/ogF5Z4/y659QeOlJ77HLd
EX5frx6jIoHdG6CT4RrYY+aY8eSLwIFR1K+3fAwiql/nZ+Iz7E3kO5+G0v6te9JIFewux/Dd93+U
jUxyq3AoqKkx2SEvhJ7im0i8EcwwK92A5ZfoURykr958tP40+HfDCs1LRv85bK4cYIRN6uLHLZkw
mMLKO14rtatMAgUeNd6f+u3mKSxCFxzHamgym5PCwAoo+RiUI6SDtY1neWXeXz0JfouuLyo73k+7
izVHT5FKsKOvKZUR24edk4c5bArrm6E0sBhKFO+GBWWkMzFypaId8WW3ng0kO+wYBCTtlsLNmmeH
NmWgq9rb8G1hxE6b+JZ/om1gGBtj2Qrv0z2PC7a7PRnsz9jjaCwpeD2rTfCM7OkxeLeXX0AEETI3
38SYCW2jQCOR9r/A0jVU6xEfNaEJtY6wY7St/J2s6YnBiyPCTnQrjPEavP4lvxCdcrkwTj3F96Jm
4fENAw6RV11EY/1BRldtAOOxTDJ6htofTrhBVZ3QiAP7A/N9V//oxe/E9iB/4e9T9LaaMlk2j7+k
DzqoP07/jBrRETZqMqUfCBaMAadQtO9tf+Akx5h/75VYuNEDPn0TsG/p68EegEhAICyS+bqOVpih
NGEMYFSMgom0qiesAr83y6vrRmwblCfI2n5ZlmjGkUUnf2aAAGRyxHZu2hxFSJkVr9k3q1Qiqi72
scksdXX1FCu89ugxrohtm+OQ/EvECcGRLmx9fPBJOntRBAyQqmSZth/6HDglz4CBqY5XczWVtk4J
P2m/0s2sNxmBH9v5MRur/i+B9F4ZL34tzhfJRK5jBPBdUTKNnvTR612bU1PcIccQqyNYxAm6Ba1n
+k8sEiBVqNDLX+1zoQc6AVWDsC29HVXpykECB26y83tgQJMkCO2iH2hbWWySa+0XVrlolIzLxCgv
AzHI6HiMvbI59vuY4cnpdo0wv+cAT5ALS8QsweQwFhbbn2RZ/kUA4pQ4kxrjZ/lkYZAB/KIaCw3R
oQwBqEYFwzmk2FrjoefnrwTC/lbme3s3Gznsdt69QrL5HO9lghxCDpo81tyQdMoujqsNHKX+BPuM
XXae3Mg3hIXAa3ra/FYS2OA2Wgk4g34jFV2DhGs3MmQ3OCfrUODQ4x6W0F/u+nBjPS2achb16S3X
PXQsPOpfeR6om7J6e28ROLrSjPG9YwS40tNAkeUHcmcTKaUjvxpYVO0FVOHAwXqW4G7J8h30t2O1
dI3P29R6LBB6DgvTJC58P0XYB8NrSji4/VRBmjYIUu9JnjpUliG+jFNZ9HGRUg7m8Q5o+hvzootx
lkKQ7qkYYnjOgSKgVJkqt4+6P1IEIWE0c9sfW37MTHfVCtpACnHQEWilM+ipAjNF53tN9O2If4d1
4lcgpb0cd4Vq7pDT+SF39y5dwpjMEedwdyMfjs93sqPRlIWbAiOKs9JTInm5Kk8G9j9FS6gv+noN
w4b7jf1embNMi6Rmnmqq16cXXlqBEd0kwnw4UvhUjRN/5/Is3QITjgzoh7YeVzm7tIAqQVblqhVi
VE+WLKv2ZDpXzGjPXhHejI32o1DbHw48/Fm3natr9KpmqyCVrxkPFqyWlppA5W+lV9cwUly/fC+W
0AtOUqhV5f15UGHQZKpmYnO3H7UoqMYJl0JG6ceAdMVAjcNtlYfwtTkyywtvFGWd9XRrPOYuAi5s
6zcLuBhLEo8gtZEexzJCTjJEi1bepsbiZ9J2odWRu2Fsq60pWvj+As4b6RI2Ew95MZSKVs+8ATnw
ikvvMCNZmtz/V66fWJafHJjJkfUH85hIDYYq0ZcoGstpIOkzuwj5P48nkVVE2HmuQrMZ9CljrHDO
ZtajwZ6TzxL1yvVu6/NY7Sn3oBXHf75PGHwlcFiZBAI96URmScqVXlpxdK2uKTzDDJiSN57f1uqI
CTleoHff707YAsmhLsXEDpQPpcDScP9Uc9EM4TUlg9RGd18m56QSWOlxxZ3M2spEHsHd6UQ3joKP
wRbMvGVZINVizNtipl+I4W0vAK53j1R1x9MbYFhvlcHiOGQECkjErrTgLdJptxKrfZrYB8gX9Ohp
dr72Yq1vCQzfy5U++ed+CUQj/KTnWSywSi62GIKmzZ5nHD7Fbhl0c6ednbuW5AgwE65q7IsbdzgN
V7AFUQlIIxsdJcdiwbSExLA9/CSVYU3XU6LuIiD3aejzLbTG/O6h8qXHmo6vyVTy5HKTey73eqzR
Puypx/wtWHybuiblqsPrmbPjkDK7i5Xo3Zs2v+RJNHjag3FWtHfoAX0lZGaIboT35CVnBH0xs6GM
+2ubgexI3myh763OxJ69u7wSpbdds452rA2cliGxkbpFIXpGnJgbxrErSMkO2/MFFTW6VYuuwhl1
/eFImQ63cQlmDdHRqb9idTqLHG9661AwDLovnaSBiAshQva75oWAMM0bjo4Wtm7PlLSzv6x2O77R
c0YlxZC5RD1rI4upCyUG3nrJVTlnNdG7ekh2cwt8o8SU+XU6twmFQCv97U6y0NL1ziaO0ME9LnHv
lG0rJ0fGsExfv2Gj8xc4YPhRMiyF3S4UDPK057HtRgFR0Zi+HiJt9V0dx5dJ+qlr/n3x0d+9JTnG
MPS/WoRMCGoHxeRcMgTi9lZMtZ7htMhJIbhkcioOT4ahNWLW7rac0Hdjqv2t8270OAmiKCNzRmea
g3Da7m9CRpz048Owi3M+wNNb7jPt8+UEfI7n2ZW6+to/P6kIot1XTV60WTaHto9b+bAKgEEjKbdb
IOSJnnfAGjyRjqcNa6U9lT/kvEQ4sCJae7QAJChckQvqx65x/ULotQD9NC7A+RFOq5C1m2J3WaSb
Wj0TCMJP4pehfKKJVcxwVj6h3r5fTgrH9tmuqV4wDBwmBekzLnbRjI97UXaBcEil8s9otn69Np9N
wTpnMnXoA3X3n7fGT1C9qj0mTc/5MPvL11dyywCh6Xw1lIVO7zLgsiTjmj8SZumQAJpTQCJ/L4os
eG5lA2QWOeIpfZbTLzlRbaX6w7C3FDk5ksIlMkd3LEDol0T8LrKTu5r2o0TKR/Uk7r6O+eVz7t+Z
Lybp0f4VV8B93jp+/pgV1SDjitIEpBSCikckV5NufKY4vN0Rk1FP+Sa8e7VyQluYvcr/wafgAf85
zTHWFjAOGrsaqjK9tusNRRCtZAW91Xf8wtbWi5BGkVlesYFZIJ1FiQbe2ddT7VZdiNtW53Yx6Tz3
gj2jlJlK8LugPOlfEviGE/RdQwPmsm1BQfiCqWZOy29p/TfW7bqirSCHGaL2VAzR3Kni3q1HAkLx
pUjEuxpNuWo+9m0CQy7v1YUf9vg8rOIOOmokBQ6Bh3bOa75n3jrFbmRPCT/Xe6yP9v4nHpN/eYWv
oj4aaR5QI8/4F809Wx1Vv0MTZioTYCbVCny4Ih6/810QxX+QlPp0qVtKRFgpy4TI+KhD59W8MO+p
pdJuA/9AoCExaa1b3B1dL8tWIg7dmiF1O4+281d5JVVh/mufENIetmMHjt8oyX3Isfs4opf35X/U
S9Ukn2n3XUrM5i0xjL4T8eIR94SQOkp0fwRz8yX1v+OYR/75Na9KzJ2F7pf0fyD/9/raftFeVWSw
JKkFoeKGppM416TgYPAetijmpuHHdINgYRuvrFS3O+vDYxgLTyK6j8PDLR+sixkUT2kR0OuOj1Oi
5Ruc2j1O/IBpII3koVZCFxhFIbPA+eJ2J59DKy8IwsVj766v2dbkp808e6lRpDWSro7PdjPSmjke
Fnmu7dJ/k4rBG7uI3k2FZKGniLpoMCV5GwK37Ijk/SYuYJ2jyO6NQd0GvVPirHZCpgzgJ7rxPBuZ
gzejPtc8I8isU9JPX2aHRECDcPae1rmgfWpIsW+c4ZmF8xZ6MENZwsBcYvqe3Feb4K/1vKWm+JvJ
v0LIPjV7uq+mL/UmZLM7EYMZhHi4vl5IHzATF+SEF91lOkMnA/LgfInY5XK77TQlMtJ2gqpxLUPL
/rJVnmGWFuLqW8yGYLkHUguGFaN2DRDre0GyuCcT2ss3RJ81vm3GdS2MElCFiV6uVMuip05IIjcZ
X+t3l4+coXyFnD22js7CpTiF/thE5VjmLXxgglpr2lxVyA9gdMdXmM3mvBBwvQCPWuSj6LQowh9a
N8mosCD2GFHggy3vfmmUMaqhXx6lIsZooanaDmLZoP3nrNWJ75acgZ95zC4Y6W8XBA8VwTYGRh7L
syldiDU34yJT3Ob67EBNePos8JNNLwN5KEUQHV962xzA3esdYbIyldl5bB59HnttmE4JTI9XB6CY
qF4KgqrO77Izb47LNfLdy3lBny61AZ7g5gLlUCMvkjY6tY4g8sg/PYlxFI31JPfefr9S2Da/+ZtT
wShT0P+D97QssvGH62dKWLarpNRUiH7IIm12Yb3Y/BIQjO+0B7bVymeT3gPOpG/huZxJqX9b1lrr
aKUfiruLqHZrz4FepFCVoekkpghQKLJ03ER9bciTozfNPH+Gp+mLtuxGLBcdBodATGrdqH263avn
fqJl1xMGraCJUXud5W4hOkic19QYyr7bD0tVNSXdktmB2N66fyIRZkIF/5j5uU8yz52GV7erbPGN
sWiWQRtmBDx3cDSeNsa232CLpYi/Onvc0krHAZ2hmQKXjfC2MmSybcjDxoIaaTqmC2HRhLl7Vjzb
DFEhhtlMA2Ds78qgpaxktSu9nxdnz4RhsRw7MF3RQeRlCm72DFOvoKvbg45YxOrk6UijvFsUHzqV
LOcrUBjg3gMZJ9t3ApmY68q0gT6shmvje5YFCaWxPkR9TGh5P7qSp1b2oWVhMDUgfzm7jE52s5OY
VKi6YzJvKy6zdXaIu+SaYvUTR08TsclCzuS7a0tpCuR03cScIQSIKAcJtEovU7t2uqnnVbK0VVa/
+McB8eRjlaIehaM0X6kelj7VPwdm6gkPh/0vrMeH0RyoJ2I7KVT0rlD410suyYy4AKigBcZiQsly
G6PN6uJ89aQ5dzN2tPf8rmYdVcAvdS9kVSU0zsYT7OIaeWBP0cT/6vTIL8PvyiF/LqtvX1EuQnim
u31+qxA2dCTgDGBoKWJtt+O7UJRSQ8wvyoyFOOiWaDTpvlrABIE86JWEvlflJ+JHo8IV/DVSQaQo
syN7SepQL9yoW2AyEJp4K0vXnOnI7vS/tiZMf9uzhpaeA3c0wIVxMviAdq99JlIP19bOWpwJr6Yf
9G50OnOLLW12LrPJdFMV+nu4c+BIvRJBoOqViidrMsPM4aTt2Vh43u4kXqwdF6CXpVOT8BzyCIBa
tjYwqpit+LuyVxL82EeuWCxFMhxV1NuCaoIF6WYaOSym6mYTg+cBFjg3FT7h9KALJiL/s+E32/rY
BSOl1efs0s/fgnLTU+fM+89fyv1NS2yMqMFvfbwQn+gXZkNGqT3D56c2zf26CU5CYabq3Fmg3QIb
LXvt8lyb6rb3mjqO6YjSUiMu6qiKHVWQAUngZOTQ+GCrMfZdQxdKV+tkQmu1bi2y/wXL2Cf5VRrI
PjyJ1zKAJmSBIAFX6NqHUy6RyImgIfO32DWng6hEUVgf+9veXJeqMMV4ftatlKzZL2wRXj7RLC2S
2DA8EJoTOD1V4qbg4aiWcO5qrZgmNdQtOctQNRulED9jiw8KgZo6sOgvi/+3cffNqDhgu2rk2scc
aIPsYzQ895oOaNd4tU7IQOLUl2G8qu2gnTFwfcY/I05sP5tfq3OXmboHVN2vIwO/bV/KSB1o/wZU
6YaiLwnZOrEP3AShhINyDMer+OQK3sPwj7JRAHLmgYXMMJv/bmle1LUjdpq33VO9d6BErUla4o8N
DRdE9bHdqJ8SyGqqrTeSk8WLPx4NDctNg9j6MplvTCk/02DAZtQpvTvuyJ44jlULNskumOX2XCif
6A7xC/TZutfwkY6IPAuB9xbXp6qNLUU/kBu7ggNbyac8GsMmWt1Bgx6Dnnf8yMoizLohmPoL/H5c
E8fUK7UW2A7l8VpNU7/jzGBtKi+48ZMdyQbvIjgqTmnLt6X4aJYuj48kJZvG0BZ3aKaJqG26VqLy
KgzwYNb/5eFhuQmT5Pl3F03eOKc8PVGPAcOLthQi2+kk590vNNaQa7sMXk3d8N9Bs8q00ptrMNrA
lfY6YrFCTzZiWZrsxJ8EQJvqnlmNVPs2vXHZ8mMOOFUnbWkhXGjAwCVOAF5A6h0+r1WX6/umRke1
6OoQ5ggLptqNp9soU1iMFIdq4uRhOIL70oatpXpKzIqiIEqj7adUXaHD1s41t+o1cQIBGPR4AorJ
3pLTJoIbjEzAmXwHLHvI/RFrqETPtMG1nX5zcjNJJ5beGQg3pF/h3TGf43u6DwnWDwk4pV75hLQ0
A/jWpSJIFB+wgF/Q8+ZFtKKB8U5wC3kPLhmEPJvHOxlox/tmgLLOuoojGOTku6HpXDOTWmAsH+iv
k8nOubLxt95P5ArVpPtgEWB4+B3JSYmpPcgkmV78lp1qwrDFR5Tqt8JJ4dxh+GH1MtyKqYBzCnPJ
8PeS+/mmRzqHm6QK8DLX3FfetoiiiRAeM6R7AjRt0z86+bfvmIlWeSN3p9EECo/IZ4zjF8zUZmJ9
uPAdtzQKw6Whu2Wo+nAQKi6LBissotoaoH02Pfg23il0HGbTj7OGLJDXPvi5J63838auFfkmJU66
n/QWfMNWahvHY/7u8k9N008R7s2Z/sbff+2K3klLW6Ye12jMG0ocVoYYhtUud0BCkWX4mquqZYNA
WYInZyuloN6qgffv03B48ZbexXmHlhnQsEWdni5xHVx7thKT9qNO9rC6dFSGujlSSOzbdh6fS81P
o5U+tM5hsFKOkMu3nd1LvMFlNVy/WFCWu4rjkufaOHYC8gsWlBEBe4cs7432S3tb9tfiQpTQH1Z8
O0X2SvaVvT7rJHEv9q1/L+0Q9wI6tm+Oa5TewpOUyQAEvkRUr4GF3j9BbMZKhexGjOxxm2Dx5EQ0
C1kjx0jhONqByo130GTMh9BlJWNQSrceC11D0mJWhuBoZqME2hHefGQN4H8osWuuNxiBrlhVoHn6
cYvZyobFcIbDF8YSQPumYloDdeATx3R5B95JRY/1VNAevmPDDEkYdiK3oaTO+L3HRPjtgh/nCEuI
QdszSmyrJNgODxYZKf7SoCt3f1eVFT2Yh+BpA5zJr9hv7zn3Ptji4v6/9JKSUB75jKnZWeDqvdwi
c5Q6mY/v/jPW9QTS+lV9zCEQ/Hfi1mWZqzEoOtSzRukA9wt2agVFRNl/kJKqCKtehJ+e2vp64i6/
GrzlMz45dw6PHHTnQtjqOBxT1scmoxUxoYAilsQcSe4Yen5dKD+KLUtn4RPcfrAvkQK7vjhyxIsk
wHQdkpuzCa/PR+Rccbh0LaztVWbogQ1ZQzj2ihM3UBREE67JSYYxAumjqwM0DQjv9pcYJyLSKHDn
xahKaR81sNgKpaXPcrX4LWRu/SHkKBa6S7gnWR9XwqXC+9gkMgvS/FNu3xwx9VJKIUxg8tQIcNqw
KExlSUtb7c4Xgq4N2C7pHiBTA3y3tURht/gP8hEYoReA0GPqo0Fdvjymon1xWRfVAWn5hjxnLwJE
E84hkuExXH5oh7w2NQosaeG3TaK9Dm9RsYsS6JVbpM61+CnEpMxdvVt0h47RlbAmoI4OnaRwcORl
erpKoXWDuE+n9NoauMK4UV8TiT73OGhUAhowadE4vSDsvu/2NrqnbsMoR/CsYwMi3BtcGd529UuU
jqGMzlrA4uDQlSJJuabKbOBbbMb2JgI5xPpZwAh+lcYnjOWoSyxkI/ApBg2nRTJI5r+esOHZRCGo
De7sEkSxbAVH5jDr/qNaWxSM5krazUs1vuyOakaysX54GFx5uZj0ciySwOxljS45ie0FjEylHl12
LD6gsGsuyFpX4/KQar+EXqZJnLhxgVdCX5nqZlwZzrMhpB/Ds5S1UHHuCcrVRdByk48Bu9TJ0XSv
hh7wd7SjM+18Oj0hkkK3udWWLptsr6XLhKQ0wzn3citPeLoFSN7RnBViQalL6OP5sqCyQtih9VsJ
U3Ie5Paq/33jLNymENysxANMg+mDGeXGekhfuXhfVB7KMF5bTqEW6CTrsFfvyyclbQvEcnRhcCt6
TikCwauWRn3clXxZiRpZr7Qy0ck5q5fM8QbBriMbv351kKwu5kk2TCyld4/DrbyAaDGRNsKA5FAr
hyGm+4Jb06VmgofcDvDSYI0dYS7a/d/9hV17JcdWu2OspSo0cnlX5elZS7yvpK0yoy8IVCW4wYi4
GvJzeTud5WEbulXfG8b4x2kbTjnHbNBfnvqT+2kEXj1ulmaMvFi4CdaMg37D7JNC5nimtDGQ5jvL
n4XcXTMVGEQc/Z5wupBhkSR/q7fzKfo4i5SIg6E7p/l1U2CS1HWjlQjijiW53OD4Qmu+F9svG1aD
vs0EIkm4QikFZ6qctWYtEEU4rVX0mPedDHy/H+G9tesIg/ZyYnNQvziehS0c52Xnr2d2mu+zSgUP
oOREYJW1Jgo6P5cKSoXBk9rNzklSpwIN4C1jdY4+6ndwGH73X6OggxzxLx2UbtBXoQngQKAX6XYV
L9261yC0SoWCgi2/UwTsfP2LKbn+scIsN5dpbb+7L9Ko8R8tahBgip7ZoUocby3+o64bqZ7xM5X8
qSpKALTl+kTHzdONjv21dSDPAKNkbOV7uEwNUoMZOzZjf8vzDlK8+3N3qf+icAyOg2cCUQDkn6Tr
CYiDpXQ3eLXUGG6+WOcx6Ztgxw6KWP1b1rAflOTyZhJec1IqQCVlHkfwmpTTuicyI7DroYVvlHjW
djxlP3LcOQoSrTlSwUvIb5j/dm6gqoSPuHR4SYjCmkxS+7ORKOMVBjeHfpf8dXPzjUeGS8YxizDy
F4f/NaOUThjxwIJWHhYp574BBTKxs4oEUr8Hu5drZt90dxUOE8hKUbnafES4jhp9sueUzIpZfHi4
jl33GRhXLbpudxnQ0+wARQoE4MjfY0uXBoBQtOWY6pEdodnGcvFKKhK2XThMypSWQcPyXc4nqrNK
yIHFeVbytxOQ9R8DjshBUVRyip6TcqcYrtOgzdTxbqIT8qFA1a1yUV76AtflYdmjynPfiwJytnUo
nOkfb6LY5+/pcNa83PpZTBIlQ4q0mtPcBg0PApKKaq3SkEEJ8LE++HpS+FBM9U5jQlPrSEJNMTY/
LlxNONa0FuwtyZeVmv2Ihutz910PB7H8CIIZ2tB2s71w388R9u32+d6cwKNsQCgXf5Hz5rbDobgj
lbkVoU/nGj+x6MIhzDBdZS/ggJIIdCHj3BOMgPfBETlHJg7WRCwNrAap0OQvFyKAlot1s9lrD1BI
kft9pUulLaw5wfPFeCi4z+SSfpZT0KWHr+/PSmeFGZp85jELCiejdiSOfMyPbSauEfcmdwj9V528
HLnkWhngAQGm5Rr7NCZepFuBV8c8hhEKTtThCy9vdIn+6JdjezXSk6SY5Jmfd18nMBNXLKofK9mH
a+XZ1pB+aZVn7IdyLR9uuSIHhlf8e3ZlXqk9Cidnhekyb8O+boncrLe+O6T3aJRbibCwzlRXKQV0
OT/d8DKXbggG5WsC5qbTSSkPL/bhsKjMUtu4ghpefAWaQNzeKCNf1CtBKnl6i6ktkdifBiBWnJ1P
C5O+FJ9y4eAHLKYuAnwmn7uCMf1X4DMan7X8vy3ngPn9NLrurdJ7wkAnCBKCtNvSIYiWEJcCn99Q
+txtCXpGF8gtG78Ak/BTSaxrfHT8J0Lapv/CsQ8OXBph1cOhTNVu7J6mAXEStrnk9YfDLpnaQYMP
di5uvgKbN30EIh7YL5OPsfZA+RriKcNrMFtHpFfVtK91JK/56AvN/drR6r09erC+1igOOTxQT95p
Reu06hQhJQmGkcUvNPcuckToyy/X/ue4QUPaWOEHr2wxoxDtvsXCUcBCvmH0ZZ3zsA4eSHYoRNAN
TR+kKS24esPZsL8VB+v/5kqXkzDnOd/sBsCwtr8nBFjGn8QYBHPAQo63S3Eg/CgPHIeiuN5Q1oYR
6wVKyyT6KGFFRedNbSXIEvid+BrQJjnMFK3zrJtDr0nyOSRkz4dIn/TLO0CuukhM02Jeby5yZCsz
Fy3KCjbC2pQ+1paKpdb3PUp/D06CL723EhzmOjkzmurV3uaopqB6pze1EIFnQ5fjA0LpDUklBbtO
2LZYscZ8GVWJSrr4lKBvDtkLsGoDFfpO75K04nSBS9WZm1gOvqP0NGZ1DLLIb2YNSiBdgX3Ollr/
YCgaCUOELXj4N1Ryf9gHA6AQisSPiqbK5sFaBYxW7KrzhDH/mkRZrVvd9Q/Cx9hKJWnaGp6i/cz6
c/E2YKZhtyZbxYFKmHXvrk1c/04j6npyANBYkFUB+PwegWfGOdgQllqOpPB52c+HWzmxQ2Eh8/Dq
qo/WxldX0P7gneBNA/qShYANpHuUpvDoGmNdlSTrrDV9l855ajNDfuTddfNkbqphpzgC4UM63pt1
YL2MYHTTtJX7dXTF87OM0Bazl7uhXRkOFqQobzkts8oScxI1ekKArU56WLlDt/8qJcqUXU1TgfyG
pi/dJgC9v5tUdiscE1gnlREQeN6Ffpz2pxM4Rx9fABpMh/gygMiqBN4vuFXM9D9fk2BD7qw7HeFh
7CP+qJOrnL3jdmcX6q4KzSp2nUU8jBREMqwX5Ij+Kv/jwr3z10XMVsVXkkfefoVYZb91qgLX9Rv+
Pugqf5BFvk1J+QMNxDQ3G7Ac/fpiLzbVNBCIYINyYZPv8JbVP6HG50md6QFtYScFNwaKBqrsv3C/
mUzmUSB+h75QbNBM0zMNV5gQ1q8rZn6cuG2rreYaxwYpcNcpmZFdd1HkMzZ/ITUimUfRcqRi93Wz
Xf/HPDY8cpk0kkVgomyvac16uyJiIAkf6E+WDEk5bkIqUhEXz/gjfaxm+bVV95OYg+HG5hJ0siQg
VNTsR4lDvWdzz/eryc199aCn4XiApVjFWmMcSAv5mp68tIVJKKzAPddmlykjAfYwgvrLayb+rTT9
pTwYB7WGYzrQqFuEP1uSDTrh7Z7Mj7k5kx3sEhVLztE1GYcpniUVLNfdJ5PwDj1p5AGBGJQpHq+c
E3bFcaq1aIUCx/95wXByCwpCWirQXgx3yT4tXxm5l3u5uPTueNE8SCD6Vo/enL3dbGJFtmJPxLRZ
6TqdIygDDBdTHzw+xNmuyM+/WckmT81VlcMMybE1/0svhdCMEG6sGSol51lGkJ9elKuPEKdM6xz3
sJO3wREGVDuiXQPVJpsakKPhCr67CMzPasQOwne+y2blIg4OJJc6591UtI8G8RmWUni3tWjO2Fow
yi6ykLjhpRxudsjQXQSoizV7bTJz/oH0V+od75XhdGAGel7/duFNyuzkymJNQ0ZM3R4cbBiu62Qr
KcP7mIQrA2NSSGIPPkAJDG8I1kXZWKUCIEDuAbemcb+KTbm3oK7YMq5eQ0Awvk6ASnLWxKX2CR1l
T9BkczF1SwOs4ErfvHvKtxIu+EItPPrJwcR+l8ufG4/A83cd1xacvaRaQu6vT2+oKLl9UisP1FaM
z4cdk7u7mDWSWBCcGwOstaN+mTkAbTRfrxwi3vGS/AsIpznNCDquNDhE7XR8vA7ibMnE2WDP4T9v
HkqO8Pi2Z0eB9xOGXewiAJKtE2uN4/KeTG2whunFhmPlOwsA9wV6QRBk9d0oB9ILIZa+oHMaDpbr
u2d5nX/OvGUCuz8jtFCKDBpqeIrbXJ3hCbgpKDuT/5Z3rIm2uxicqEU/Q+rkTgXHHBVSRDXZPDSq
dmQzHIq/3k+Q4eRWJmPk0mL0AmdqCfOYDkqLIwtCaf8zRZhpkOyZ8KyXceGA6KgJupB733EleSen
O9QZVLgIHmaAKVeffziF0l0SvbWk+Ijjmpi7j0pxyb2Eh1URjE+eOlCPXN6v1ZhiJPrji/QnBAYX
WhKKK/3L5pRVOzprm+A4FFkrG1/9PSR3bi2/d3uzFpqKu/NaWskiVQt2e8S46Alt82NQxvS6FuFE
peEkCr1eBGHSgHQsaz5gOxj4u0D+dsN6zaT4E9/MSMXmKhwW+AVliJQVg4kt1YsR5jFdFBOpzkIY
Gqa/zB4sLGAdhRFIBgr3pVJA6ZFkYqCNzk3XFPyG1Sr06S/+QxKzKmplath/9Um5RQHPyG8/Y3wL
k+Y+jtRzKeeNXRFEf32q9Rlx1jGOxaZ8PWckl+AzVkQlGbhNV/ib6qohZhAWSGzs7va7gGWx/qD8
p72oI+SD/FT8D4/p9Gm6P0qr4Q1a1+yqQNL5znZjFMo2+IRt3PeuLQWjZowlcJwHPNqrJFf7KIww
wMQvcJ5kb179Ayos5F94szWvwkrEAj6JObnNxcGGTnG1PV6e8/K6X4+GRSRrzbu4qkFOO6N8JD16
bcLweaRakeZJJNZEzjdE2/d7CDvwdj4vkVU+mgZac7UWdgKgubX2xCuyQkrIsPC6+tUWinDJG7Yh
jN7fKZ/W+ChiKA4Ehv30nFC03Q5ybY9AqmGH8W/F1+rYOiwuN7c3JyIC9aF855bm/FnKQBWInySy
pQMN/XxSWVXvicisiPG1XABug777dwVtqiJFJyo9GY8xLaiIZ7sffnz9+IubVS5EECQE/wE5eeVL
El6Q/kiDMMSQjCO/sloE+V52eMwCN7vbBTNbihzrbePgVFuX3P4YCse5b/aa4AlzdVA/5L5kDWeO
cR65YdWX4LMSX8zFZhTZHPycgJ7pp/eQKcs7WmQGokNv/6OzI6FkB1o4Bkk5jWV0+IvJk1+9QoqU
IHzMV1NDq7eAhe46+Ek4/tX6fkE+SDYAViobf/Ki6wyiH63BvJIj0GH42x3aL7rz94phvmNEUT5z
w1orycIIcWPXxp2yeE1iwUATEdAjkjqv/6oTymD6/1QT7LlUdeXpIkaJxkPYxiely1yQTkERS6Ub
oGAHqz7tRyMgOy6q/HE6omRth/gqqXPoGyvK7wf6/WjfF3nJFH58d0ZEXn3Y/zaJUkBvh72kTuoC
dBt4R4jPutVp+ZwWXzuUKEiLbkq4eqAIkG3bk8YWLsb+vd8Ri81b1XA4Rhqk8axiN3zxgx8tAkeq
3o1DLvhm1trdI8A/D8mIuFQIOpUMsY8cgqzTiJkpEuhqQVl8CswN7oOouBVGs9JLn73zQwmGlTb4
L7o8eSodde+itFOUJHBc2Cp4QWsLLj6pH2qcDhPcNgmRZOFA1zkzBemJ9dMSjT0Xrvk08LQGt9+N
DixOibcm/FUxj9/8mgB5HUxUMZoHy2CCpCKBmScVmlNG1uch7+C2Aeub/VssiqrviMM3m9QPjaC/
STDoN+ge1mHphU/FIzLuhikVC3h7O61+OFaQEbnk3oTillJ4k5jSs1uuMzzIvmqJyDHwfh+ctI6s
a8ytLKX6zTHVvuA+82EPgBcKbxE7WxcwDHvMxPw4qVdLIiqqhdma831s9ZzHalcc3b0e3CtEUD88
Yy8VFSbIQdNEBVi4EpikhdOqTYWZ5ViLmjZW/PgVcQp/3dVd/omWYsxLemULzbVCLH/dH0DHM5lW
2aTavjj+hMAA0UwXPX06gBH2Vte8JbKFFRHYNRKMCTibH106eNE5l3mSEwCxdVDSa81DmFp9xdIi
1iTfCFN/0fPFY+edPsRozZxOLWbf/UZdfuEa7emOyvFJDqTnqHGSJ/v+n5s9e2EK8g3OJgDhIuzR
tp1biKJ+EOQDefIcfO2b1bb5iNKG6ZPlgGS1gumQpSZ16tl9nubj6/+TIYNNunUPpt4yRmkDJbc8
ywrA0PPY5L8KCgJnYILzzkH+C05WOOJkjsPoh6NS/enIt07ft3cGV7FEZWf+ya87AC5sZe/W0h6z
pv4fcqRpdlOd4GI/qmNxM0l0kb8eTgYRAM/fAYr4bxR5R9cp1Uxy2V3k76oWbOQjJn+jEf54ikKv
LfeC1WdnbEld6adQy17+EMIk0GEBXi0TCRPUr7tpKld9Ty22wJ+z2IFrkqLQs7iNRTPf3dEN3B2F
xNvo8Ps1cc29ib9FTYSoMy11CJU2/qy6PinXG+fI17QIAOUB8kyTIHQ5al42KRZ7WofAKvbugtKV
N6e7Qy5zve5EfeH5NKdXYeAMBrjJvshxSkSa8J4ES1ViA3kDT1ibFTJ/gMpRa1HDXPoytOACZea4
KiZjbmHZnuatZ0I01v9AYNMq8rHCm4Px09u4ACkgcshFIU+BmvfWqjuhoI9NrJNBnNuTyin0HOzX
3U7h0M6Ii914AksNOhyx/mWHi90zJTE9CR7yoetU/la8hcmR8Y6IceVerHtOh0Dbd67hXY5P46s7
UeTK6Y1R7+ZY+8Amelh3mDL1Cvx+drSS3uk/Z/V+dkmrhnZkpi+HZHkdbOe6UkGYvWR7trIceEQN
ZovTBGA0qkdbqNq5LOqDOYx5P/xHl0HNNy/y7anDd7F3U74mGiGw6ezma9lmQwhToJRpcgHhAPsv
uL7nFzhzGOsYhykwkNH4T3lcFl/cKlN3+OBEBsfliY+PYTov786xV9g6svNTfpRjbVqGZHt2o5ov
wFkmdkw3zutqpSZJgFnGy8bliMN/aw2+9xkW/NoF6+9lb7ombTH0qSEldLzmuSjM1ff9Ta4+/YPT
nTDNmJFdu7wzkzdx/QDLxwnJicET/WOLjm9HRvxnIbEeSwlwVorat7YRKgLxLZ6XzamkeaKDqPkL
e0qEvt/T+nJ95h2dvzOZ2F6LNqJM9o2ttOLTbYyHe+lkg9pPNwu7DBZScGnRHwc6nJMZioE4fSl2
X58OIAoTGgQrfiZetOBqZIp5DEWfNTy4TjpW/vnA9B32oJvOdL+MDLj7lwUy9hSajbyCYpCG2Q+v
egki9cIHjgFy97CtQWnMWDHOjMou43IE4dxKgt9l586KtOiPEhiJ5xBhDnq1Sop5RVT6TiJCF+y3
UFI4hnuKUTcYy8fhLBhGjraetvEJCb2UrzxNsOOUvZaL7inPfhkArxjHr7fCwPf+c4h0e2j2i0J3
eL5TH6L7HvyPs7Srs1SPy61yvRjak/S6JaVH/kROZF0nAZ35R4iJwgHdm4lhOtgNXAyroVlsvnHk
BfmdFTV0PFpNwV/2cCzTIgt04atf/Dp/VRNWHxAqK1DKWsg40FcKFjHx8XjBMchWzIMEa9zQ0IPi
dw67eupbAouumEVnX+sO8zJJNaW//Vyxhnx/vB5ObiSXQlplfqfUUVveMV25GF33FFj12wwK4VWW
hdPrJnd/Cf6yzbDaHvw+08hO7rWfA10Y/5U23ja2wHZ5sC56AUQlFgtC2Ja+bGI0BMx23jdA1A7q
PxLXGheAyg/tGEWbpLLW7z0lE6Wg1zhTd287utDyKMIOrKCwgAhjzQo9DFH829NveHF7kmph7017
rU213JtMpsAGdB5K+DeTIm6wSFcTykbWneitAOpsxDJ1ih8OCnp/PyVFh7TirOBkvv8kqSU5Kgtf
F2GrpGr7UCXG4EUr43FfkuHoWWsuWPxyf1I68q0CKyRTzPQKnPYEPOOTwR4kjQBHPqFS3jO72xPi
KuPm8WxTJbuv5rrCftI2gNMUL+TN6Q1Lggcthyzzshrhz940cRaMFBSNXNsKQrQ0NZcbHWd7pdpn
c24Bvh62nmOkMtPZfwOslfbzfoEWJ0P2uRaeFd3Luxo8LcBZSFJX/qYfDJdrAiQGxDetHAkqeBd5
jBQ7OJQ/LzK1rZs3C3rBt+zy5RXJ/p2kXuUIF4AuaIL6yh5eGgeBlyyDAnKKTSppNCcjXhP/tzxG
KFMdkZ5HU5NTa+A6tEJ3DdGrMWNuPicCIZ2bTVCz+z21VR+jGvYV3fhH33ef0p+bh0UzsS5RGL0R
X3Sf9h8zPQu9NWKqfAsMwCO0nbi24Ws7N+5C/jOiPUbb5YCs2cqgphAcAP/iGp/R3rdSdpGR+wXp
noLQ2N+hrt8CIO4q1Lbg4UetFB8qfsmsAxFd1UF/5ugnmE4KewJ7oYB3H7Rpkz8YhCbcewQPq5HZ
MpX/7wpLHwuLxHUwFhl/ITS0WbzejPtnyfPh7GhbiqtE/wRq42Pz26cHjOTJfq+ewZPE5eiZfe+L
a20l5ZYPxsZvuX9J7RTzXhdejP2nsT4JEAn8coV7tmLYaLhOQMj/2z57pxPuTo19TMDVapH4H6Th
ERtOOogRkglLalLYY53Sy1dImH2vwlidPIkT1Ii9hen3ZUdIZptZz3gnLjQ0Gq7G+QLhsS4LBlnr
t/+qGGcE9w74menGzDbvw+fkUMign+qdJp8oY1yviVLjVwEjTOHCHbHkE05TXOQyPTukuRXPW5K5
UERD9MBHuv8NXT7B9eSlV1I2iSSVRTHoNoXjP3rQKw5nHCDG3Z7P2jb/fCrl7OB4N5TD1PTsgcGN
vQAwcwaCv69hEMgzd/cfw1SgRR1J7ENcWX62HLwMNTkXZq6EQe5I0OU6aKeQSKmjQvSX/D19hoik
gvYs7tl9/NlDtUvyRKtVE4YhnM3a4SpkvmwVg2uM+t0VTcarMZyI2HlA4tUYjYaQmBGVF3Y2d8yK
Xsmfhm17uhajJp7fqS+Cu2W+cc5B6MSJrTF1Fm32OgkKmb34ciOyDgUwWzxMNn9sDPb7Ay736wdS
p8L2mXbubhsQGkUI+78ACH6qrSGibWf3gdjYvS59kT4c0zqzUTPowzde1q2KT1XiYN/SsS7W5LxM
LvTMMOfpSj2MXi/BYiqUnJ4oQgYmFb8ppiagj55QVMgiQTZ7urCOKKotNorTcZx469+W0P0Ay2ic
XzHVMuCXxff5/esKyF4ib8vorKj290Z084ax309nHIANsG15/GgzwK4Vt9Ama4FozkA4BfZhRPwi
Fbz5FsmTW2hVndhtyf6W2M8LS6LqkQAFAa+nB7YxAkTOF8yj7tuqbnbpIdZt4kb2gI/0v4PGGVr4
EDhuxSDB18CBv027Cnm69CESE62pGFUm4aFNeyDOdDYnZDtfscrwLbl7Cq3LWNf5uSreeVt347du
Z4JZByfelUJxzRy0dgluEH0a5MWfAn1OvuwlcOO9DFTbkNejbEZZ/VW90FMMZh2xD+9JKRLRYhvN
InAtSbQmB0jEFoTLOtT+t5ezgaBIpuLeNxPZWSTZ8zX4jW2b3GQc4/2JbUHj0iRML8uKp45QuJ07
U9q+ApUh6qBXxnVy2qqS+kR9lKOp9LVAgafruUV9AywAWrTN9bTuhOm9J29Za93oGqAUt+NNyMia
WsLvUjqzOlASLXXnsVviK70fXaheRebLHYm9LjD074YMCl0iokA8/NcgjejUHYaruxfKvj+f5TFD
CIsjfFEFcgqac4APXddBOYaqcGXhO63XBhSSHOzizfbeGvo1eFmGxOQsW1hXSRcgGRcLSZHHv0Cf
BbhphFxJHKkn7F2AhHg1dLeG3EMYoM1TsKJxElNfGRhsVTzfdBuDq1Eg0rI22B5F1NcnTLK7ikho
pjf13YBcXR8mqUCh4DeQ/3uA2N+MIwHCFDnItoAKS57lira3fp9q3ClXgTV2C7VqAMwq38GQDJgM
UgCOveqlMg63tuj0sXS/Z2R7pub2vtbtIgoiEtVeVDwUXtUIzI0/9aXzsb7hV7ol4e1SZIfU5wI3
kugyfJZAL2Ofhf56fxptJCtidJyhmRjmAO/z9oBp/390+d7NKXadrfKq802FxVfpCEiaYkhcxRcS
GvtXXpM38gFlJHKk05jOiESrvLV+T4N/hfTpBLHa/88qk4XpX3j9nwnHWLos+zQwb9aTgMlD/Zg2
pRNhSzeVIJZ3k3iRTo0pxIkqp3Y9vrOH25nIvhzi/0D1tVhgfGJ2+ungNjE9TTCdxAcZoT/hnE0C
n+lheXNrorlM2V/LaF7buQGLbQ46zw5ly53FKT6LJUGuNOaYKC0Z/r5231nS2pVF0XBMWbex4iUs
faRWr+UqIEH5J8XR4jLI26Ht4QOxT7qh/EtZqQKVGf2wxTgtJHPH2zUA2UyzJOGBHbmsB8D175Pd
QbP16OIgKAwv30tCrOBfO084t5Dyc4vBjdqh0hU/4GsCz9isygxvBOp4tw81QaolaivG31QoZcE6
fZ1FB0AXaHnkDiwbcFJhvjKLRMol2n7yNroepOSM2Sdr1Q5sq7YyySzLQzTfAFuMHi/CoPZ/BgM4
bW1oBAc8wlgzy+6zrjD8l/ZukKWyXl84EeirFysaniOSnEhIsjqASL8ru/QIOaYvG572ZT3AkbfV
+D22EgehEWRhOY/2KMoYuHWyqhe1vtA5ZVItGxWLz1MkIbIa+rrrNggfsD4C6EYOhl71npyp0pA8
7wJndaYzVn4xNxxE/xHov6CzExSwwZjchhobuLy19HZoHd4M+CrQFohiQmnGGDyESEFBZwXEPHvg
t/GxkVs8sbHIpc/jzrFf4gi5t+30+9LKIcUVCNuqSvV+L+jPFOlL7V1h4QlSN1pD7XZvK50CJNW4
VsnE0UHFIL4IK3g7hMmQOynxDHVtnalhzGksdCvGUIz1sdGAt0ODz+PGQXUE3bHv+Xe1x+vXSG4B
3cX9Yc0NhZmGiwzaL4EGUb8VQBkbHQ3Q2L96S9MvkLkAaBS5F45VAbl0Ob9BhJEW+sk0FMxF+Gyo
0qSZXz3ENvq96J2RR6dfD4TQ+R8h/qsEGlgdUjLn7D1MPHzBHSxzJFUoN4Aoj+48PjJHeZbNW+ro
gfD+cg/+6Iys0kDGR0oNVtKj6d1OkU0HnlHKS7nud5nMUJttcYkqVM/GCQplHXmcDRt9VZc/Ds3c
+/h+NyT/uqiPsRe5aeN79kO3See5kD/cvc0jIiXj5+52DVpXAHgo4pw0O9bD6Tur5f0PffKNeIDD
s+ibbM362I0rcSnvb5YHunEOKvQIF85qgrbEyn0w8yY2AgYQiQq4/BW7QkRTyuAiWtp9dSt0Npv6
BmsRHgh4/giCzMH7VIpdZgjNyhyXdU+88xPnJlClMXGhQYtSHPjjGvxbsXDqP7/Ac7odRr+lnqlo
VIB4pZL2eQM+cjWAJKk4VTKQu89r6Fl8sE8s5GnrJc7FWjMA+KejfxtObskPz1B9T5IV/AI2hrQg
SRoGn5jNXrciiEFm3UXTMTDAnI2WIo8fWxE1I/jqc2Nu/50+qTf13WLXYgP/iYIZksDo1WRjyK08
8WfeR2OwtYzweY7oVmr9HFlGiGOZGHg64Vb6BZDwzq2mSlNkaqvA8IzbI2zwgOk6yPJzlTj0CA99
Hetiw+6gPP6FvU0w5OYIJmdoU7CcKUjTpv6FAyri+Iut/PgcqO2mJT/2hE5ImBeqzr24kM+ysxQl
cfk0DXCHXa6KFuN341u417bSr3zK593ciz/OqOKk2bjnWLydAXjWC3hKfLG2aSB4zznRsq7sfy4Q
QUj/ZZd7SL79uVloVp+Q1Oz8W1H8XsvTBflF9sQV+FAsJ9bfk/LOibuNuXqvdUDmakDFXy1gXaHL
RrYiYuSp5ImaKL+4bwoecxwutGarh1RSS9J5tKjFbmfp2bcYhiZ/O5hALTS5gImQR69ba3wc2Lnc
1ct8xJqlRLTTVhYcTHC5ajnuzeo7qm6KoCm9rsMiWiavlxCd108YD0rRKZKg9i0PnfqQabPINbj+
ngvI6q81SvuN9B6TAuG71DwVHqp5XZpcxAQB3PSvbbg07IrihWsJLH7KNjEaWZ7dJWvld8DTxU15
zW1WqalINm4XPVZL95xly5yiIMlgq00/T4phClRJJ/gbMct+cp73IlrI+rrtXdMKn+RknJK5VE0l
l45N9+szdmZVD4N5VfwJAY9KRxNPMKokmCViCxl+2gYQ2lvps+D/cBAMiPhKkg6bnTjs1K/DEjVb
BBstgyCA20QY0R6URJvudyYKW5LsR8Lx/xxgarFmh9xDgb6VUdM0IO5sY+Gkpi5NcAvrapGMkrru
XdcuuGVNWM0SeN5W1C9FwuEqI3NZ5FmbD+ddaCQy+CrN45WvfH2/BKS7S9dWM8I8MG4ajdVHgfFG
HBJk+bV2DX1KfW4Zci+8j/kwSTIxK+Ut1BsXBQeAGlnRQFUpmBGNzZtcC/8/zp7OyfBESl7H6U0Q
BHSUtDNdpfbmB6AfH8URvEqDYm42gtkufAKsZPCyuXQKNPHfhBXiY2+hhRk4+/qLmppolNx/K03L
KzC3cA/DpJnWE7SunjMsLcjs6V95bGFaAGM5ymtK1haKASIOhuP9PgBFoBfsNitDr7Al4Ru0/BVP
o9Zf4wicCc/mFjgu3yeDc1gKdTYRIByiYuZDXqR79VWQnzgiKc9qb9QHQ+pxdN87RVC7u/frf0bG
oeaDG+3WytkQGjMA2xWzlD4FsI/+2lFXORmStDI+iymREYSAbZiINCutbgHA8EdKejCdDJpNnAcS
gv6fqExCLxfk6H4loOPprYG6JyzWqz47SETp+8GHf5zvBIts8vjMwUxXdREUvsXDzZJgTapGkMER
G2gcSyX+lwiivKoRbY/1B+3cROOPZJw8zpjdLlJpQl/ge6TkFroi5NaJ7fqX8uT2UtVguZFpI1r3
poPC9HgVnLj5Q2Ek9kxa6fOqyokFqb7vCasLyX8mf40Ld44RE+NBJZ73b715A7KM9C88A02iTur9
pGT/nE3RDO/nJpvGBu5ommGfb2vAfeKMUG2SjxA485fKA/7K1EkBJaZQOz3Kz/RKkYRaJq2Vv/wJ
TUjUqEYOHbmppRRw6G3RlrZ/lKV6IL153lFptASCA//e6YutKjWOAFNpIACCO4ceW4a6eUQaYlA8
DqgzpjJevI8YbOtFqu3UR1D7jLoFG7/ifT1XAf114LfO06p2fndBjD5oi1F1teUz2qZzkC6b9aEI
SqluFGF3QmUcF5dm97cLSSbfIZ6eCZIfz4qO5qIa6fwLYqjpvVPzyjIYKePlyM+5Mv0jpLG+8aGt
H0pl5vDUT5QUKhLsHLfywHl/GSNYhFrhVpmUHVJaLQhXRKhKKxJipV9S3gP+aIIEcAUG0gRUaKFU
cDENstebwjMuM65J1hb/WlEBTNlyFt5wpdDNZHC6UiKsOBd9gi+sdO+6FTXuLVrhtJjzX5ixFCFP
G8Q0IowDKcg1mayAVdqR3+r1q/jFsV9XRKazHIAMo5jT2xmSfeq78x7Un3LmxeQlZBYBYceLqQs5
Vt8pdhPmxyxn773u4Leo18C8CVnptMKzyD+yzcvdR7t6SHqH8cPft3hDlk0+jxYQxgq+mu7JHIuc
bVOVQ07tkVrtKMsctRGhdh0Af4A/ADgkJZUjMiTHL3I5M4F/rAmwlyqeJCyF2ooqoI57R14tUYZ3
er0h85pt6oiDmmYe4G3kFloy8kCwb7ebx8Cd3WLkNbuM5k35GE6zz7j6WwHlwsjzCneN61r5XfWn
0f0OPIQqKHS/PQHmJPXZp4EmZIk1pg5LwmrwN7fDX9OrGt20cQBc84GFi9JGZGvoNHBYp4NSXtLm
FkjMyDKq8muFN0RAvKmKhfa6Fer/GiAv/irrxr8rkAjeSYF9nhNHhI3wqkT5r2Xogm5AwlXYmTyf
V4B2XoswIgQ2V9jn8a9kR6jABZbd+F0FlMAS4Ek62mwMxgKKjGGsuR7u4GckY3v9IGedQSmrLOAm
mJGiKhQ+09Y73QI0FD87WesKygwimRQcCUdGgBLa1B+CuVd3WAmulNlEuWnTq0BaDmgR6n0mqZDW
6rguulL85TOGXLia4FrXIMYYWfQwd3E0TFDomIkdHxP7A63oxdmy5FGSgU39hzIpmJAbonjobUU8
uJo2bsi4m+eUwVK7JkQhr3jLI6oQvZLM/LI+8IoIPIoOyh4uFtvE5K+maiQFGdo2XgBo6Xb0c9nt
4rHBwM1LUHoCM+Z4m/ke7UymL1BREHgEK2kmvKk/xd1MXQK8A0h6LPDWbs+/7LlJRLlhlOXNc+IT
CvImT54N8Rt7lSwtPnwurhBf7Fh5JQdTKrp6ZCSJOhd/UCCncGvQ13W+Iej1Ok3az8z4dndWq8JU
p+ZKadC0C/VDUTi4Ba8Cl1k30TL3SiL/d7ibn3+i5LbVf2QM+KgqQDhEZ1WsSFo5qDQHZpmPs1Pc
BReH5YFN4w7wY64x8xMcvvHDCO8EPbMJGTSP/ToeALGXg8wk4nZ4fsusj2x4wBW+2jOozGqr31fB
kxnQUgNgn58ZyptqUYeNkD6+ZQvTxywLlH27b5Fl1cltz5Ehe3k+ClQRVdBhIKfca/VDG9KqpUhR
56Gc6zHIsu2JnodnzByb+ECFJhe9JaMFMj6GOAD0WzoXyKcdEXRf0vKa1p9EdDSF0qpoDTdpvG39
5bK0p6as5GB/3M5HOWKBXjWdEBSaBAihjhonFZF235iVbSznW0v3HfVX1uIHMITVhyUshPZNwG2L
HtQPoDEcRvRhWpGzz6JOht1fWW2aLJdW2PAkGAsXnmi0z8/gB6uBNpF4YgUAteKKzSRu9HYk3oGM
iymbzwEJmjT9O6CZXpyDeW2TFQqIO/ORxrGpmxWUzhv/Cfe6qL/Cb8xg4QRG+U+CE0svQkaR6jqn
4zg/hokNgotNIzUnjEvJJn5CYY+CHTIcpmgGpdD02BQATrbYn+6HIjhn0VnoYIXls+c+426DkmhB
kltkLOd+1foz59gfqmZk2C5b6IivtTVGi7QlHDhOMHp40pMD0QP6XUXRsFwG+XT7t/q9qAJdBIzK
go+3420ueg4ygQM80pfTcLBKhkybh5atPj4D14qmi/d48uhfXaR2IZFK+am+9LXjzmLfg+qJgpsI
CXmkwlbJzSnsi0m7kGsoPnZKT4E1aJTvXN1S59/rZO8ZCh0e7Jw+isHPLN0hUTGkk3QW+2cceb0Q
j02rVTFnxW7GLNUkEVB/EwuguFHOnYF/I22Mg2N2F0Mw7jGfRqo0PLiYDH2pTtM/txY/lCkZQbGU
0ZtUGcPD1P4f60mYqaZ0QmXtXM0lKVwTbeQ9Z9dWOzGiTJhSfbuprEsd7G1+DD36VdhJXOGEyAI+
BI38Yt+xIRL86bkkNT+CZfqLU9p+ipWnqLB/Weat+3WV0RKiUHyNA6HcnKHfcJmIsHnWVBZeLe/c
8dK+RkjsvLLHChGAMWZxhJst3zhiY+eG6xkn48DW7407+BnNbL2j2XSFpbaKr5jSIu/lx3rh8LmB
V230OZecQRuUMhP2rq07uV/nNmXxYk9w+brzDlxIZSL4WgHfV5T1ULaKtaIN5rYr0LpLOSm2bumm
MHy2LxVWoaKjc4/5lbSTvwgWhKj+qE+uHJB0pTc0mG3d66V97rm5Kj4RCDzrjigcOdNf6IKlJa6Y
IrZUzV5P9GsjE8ic/TlpB8/mbCvZ56svfdQuzRwepoImcEKWr+Kj+0bIn38zkwQI8MyTNE/nqbWH
+rls0W5qIPGN7+LWsJHquVw7yr7bngwEznDQHDYyZQzgUP0aghTLjNrEJ4NRjPU16aHoBnmdUnml
2r0U+sdexun2JGuMjrwbWdyzLYyGJXjfhHjvE41JwV4GnVZZ2r+nQyLN/QlDxzZnHavu35MwxczN
zxtBdBy8S5wlfv8H4mIzo6j7je5FToRiEYerdTBW6gX30sCtoPPED+wk8Fv5hrR50o2OVpjDsmH8
GoFoxhoi3i/T1Vkjx5QbLupwnzjfPsZlPZhN5o74wJHH1I3moYSnD/LQyW4R7RrJlCk8EZO+HVaJ
i/KF2npGbTvoqPubh60HNBV7lrVxX0piLi6HiIGByG0aMrhD2l2f13LzzpRsr3AOkoNOEdAAe/o7
YhOWmvioMvcOBVd6cM1U9V8/Cutv/Tqr+L+chBDSsTlJPhX5mBDmySdQEN6Uxn6QOaTfYEQETkJ8
MCM4HibZPb2fWQUnwHAKEeOC+X72b7Uo0fG3hTetuOJj3TpRuE9fxUwLe/azvii5nCtZECjaE4fm
2xtrhTbRxT0FRc0VKA6RT+eX/67egrtmvtVW/GxOywDupcTArMdkd8qoxv36c41Gf6aqZVQzgkb3
w5EeR/LCQbetpvT0W2PkN/q7aI55YjfKzeGfh2sMyU87aIBf76kliI4Bn9Flw5EEmPmYxBX0xDVw
B0U8Icqz3VH3ipwQUNqTkVfGuks63QapxchLwXFAXw6j/J1MQb37eR85GdLyJwwivcY0xWqFLQBJ
FmsBHVqRoqGF/w29212xvmp3rXUtwMlEtrmfIV5fGNfWeJ/g4RNAGJuMQkBECVol5fwKJi7Aa2Cc
B68sf2B6xf86eeaOOiO3y/ExNr0pMephl5TaTE5tF2k4DlyBatE10/W+rwpy3UZgP58UIfi7LAHE
4GzkG9OLawq/grUpP0btV594Xsd3ibO7+gE943XRH2Ovpic+tBGgfjmBigx/MI6PFlflLeL0wBFO
hBVWorSRPk95JZ5/nDcazw9PmvEp1BGF6pDmyWN4/PqWhcHqUEzXha+Mka36uoBCZC56zYTbWRP7
2+ZFU2DvA5HZavG2CQ3hq76p7L/Rs6rejl36rAhI7xZyFcnrKEovdqtaAJS1vKMpGEWnRUw/J/Q5
kpSKvyGkrXVktPR/5sUqSJ7m7vpo3xw6L4QbBMo6uUgFwgnKhDPL4f+byQKXv8VB2pMArz0ZN0vO
yILlfEpZihskS1i2T9QtvCMLtbnkVYIw+VxJG8eylrp0zW9sLtFu9EFW11PLw9B9XN/vVLh4TAEr
6gjIlXOR9v97UhWp/GUGZZWTlXhd+Q/aD2ttfs3mjqwsipK4F/Z0sAT//blhMEff2LR74NqqhtnK
+hE6pVbfiZ5CrRPkeS0QFGwqS6eb9Rzopsy7SVzqNuIDMb8/vnE1BbcBlB/hZC1muXOEw95tJiTN
zCmbwGscpXrt9cL0oTH6lRVBMsFnXgfZnKic5R/ffBjWRJGpgf5XU67AJze8YuiR9C3Fy3MNW4ub
npDjdo+zADuGVAnlVhqX+jBUM5tRFfEGYEEFeG5y54y2kwBLAR9SXgiVgJM2SlQ19zXO9YeFkdPm
2KKasAD23wep2WN7Giy5uJgRGGXEXcP5JY8PqGmzYgrxcrdNVNGUS8c5nOG+J712iJAB3Qcfznaj
YjLs08GXjp5+Q0XFWHtNl4DSRd3wuHg3uL2P2W52ylawwMA/shzPLQg5rThF6bMXWu4Oj05gbeDE
SxiXNumxsSXpjPyE2+LwdHlqUbnQoDnfDDRrbmq+7k4jN0QYFKuWzNoox/vTSV64FQzavARtBOae
rarCXtIFiqlgOus1ToQaOX2hxlzRjeAcu+dAsi15sczWblD9u20J4SZh2cEsGaQ1v3F30Oxda8S6
XKK9WpN7HKRAMYfTDdujLHsbXa+69MhHmRYLscyeFuqMsmnY9ZTv1e1S4K9hMDVzemRneJZ1/O3t
J7+CuZGjDYMdvgg4q9ow5QSueY+RjRXwYPjyiX+lSNd76F/SUvLCZ9oTJiUJvw5fLx+U+ErPD0u/
VsH0CDFi47KUwa8hfUEg0BugcvM+tHkC21aMukm+RRma8Aq58RESS2MHph/rVEvtxlDdlZfq7nzA
lMOVNR82yVU8+vHsoGc9emcIUNt4vXlr12h/JHp7TJO2KCx0R3KENvjsBuw5rINZzixUoEkicJYH
uwFySXCC7ryP9AhlprFYHQdRJYVWggORngNWuJE2DJIhz4wfhzNTM+pfUBJB1CEzFnNLG61Q8+SF
Ff8p+Z2XkzRYp/lYgrj/m/+Z1qXGXfbmO7b41GvRUVFaPV6IFH86JrmaCldFvMdvtIjdvMoPeWMw
BgLR+VvOecCf7E3XgAVvHBC2pXo6nnYhajuuzBbKxXHdsGslsXun4VUnEValQ+FuzdgIwus1fUmU
pYsMoTsj2PWohTWEGQK5LbWIdrxqy2x6rn78rLlI0xeEhHW0bYilqMWx2taDmkgQKoB1SlOzKmMG
C0Y/pfN+7mK+h3SZ+j2prNp3SVv4GfWlI7EDRkL1Z1dTMCgsO/n06qGsiVGHPeqo5zRkAx3FztbR
pJGMG07f7bT+XH/lGqTLDm1mOcqfnbusgUJM+0z/fOtXTUWJbbYphLjY/cA08DCGhpEpqkXXorpf
XwDCXGcY4hoAxCBTMU+OgMTo7W16bOT+jEyQM8dWao6YT27RmG9T5DsI5k0BOJOT6k/JFvDP3RkZ
rbS7QuqkkLLxNJ3OeExj9NV8LQQtojW3oMfDYinwXQPJiP1cbbKZA8R5V/pGwXNjIJ7N+mhxDTbB
Z7EL+BRwCs4Zg/uyqTe1TKYYBr+0w4ojBLxg7fqvwb0rHI9/E4RMoJhbWaHW4Le313tty5DigVA2
Bvcqt63zjhnxZyko1GwH0AK8jfmXEudv0DEI7u8AzM1ZnzOhIA2uSBrsTxAKMI3rVE7aWRCEEBYD
UhXeZ6fGCoC5qqCGQFrwXNhchoLqz7j2UYt55M+kctPDaZI64hy1JYgfMpfeI/Mta+hsFVsFkUPP
KDXxIfpajjQJagJqwBlAJgzSwimIra3V1f+aKBiRAdDHawgVLvibHCxlaiHo4czeVP3dWrk8uMM7
W1xQiy7Mclks/HnrD0JOVk/3Q1T2ZXBY5e4w8X6ztBQDH6P4uodAa9jjTz4wg5voADcnFDNfduby
WbQU6LOSl5fy9fAbvmsrscGPdzghdeEe5lTvjrWKr2jbEBlhHnKNO8wacxnsaR9rqggIRwM0y60U
nfqVgeJjfxNIs6YlD3Hfibn/QdsELQudbEOT1jfVYAYGh7Feda80Egfg3GOv9Jb4Sx4IgOWZWG9s
Y/IBp7okUOT2lwUSNO6A4tAYV0j8fid+lIGnnj9iO30FH2laAkPXH0zHfyglsqco65MmN85xqi83
RXO8HBOExr7W9RiQRLwUHynSJJ2c7eulcTrA4YcBazcwu53Ut9R6yyvQnO7LKZEdKdCknXaAvncd
VWwKpK9A1hbX+brZSCQ1ZALrdE3ILoOAr0qYxOtsx/ynPMMbyxzYfG7/xQrNHTie3+AeWwBS+xj4
9YhNUJ3nFHcQbY8+PhyE/cfq9W1OKjAOgLbijzohSDUO07SrkMkoJuMmv3HnZbo3jAPBDWw7Uvdv
XvHuhHtMi1qqQUf0Zez8O22S16dtCiZBiB+SKl4E5uEAN+CQjB3pst5GR6tSEhMNW7cgeak4xOll
/k+ihucgV1du9pSSIlazY3WoGpcJyUaPljC1PT8cl4A+8YufnPEBpz19bsDUViOjXJ5gPimGnEDm
1tKRf/q2vgyJ/9n18mg3O6U7fG+NEmVPR1Jt+6An4yz2yPB23CLwPfkbiTTZvTBCVtIrgNN5Q6Yq
3/NzVBCUejo3zjW1koYc3i4yj2i5LmQnaqwTuugvlpMOO2QrloA81b51PcclNuHWv32fJa0sig40
ali90JOTpXk6a2MrcqYGu7XOKqVu6FVQGm6TMMTS6bdP0XO92Gq3oAXHz6zeAEEoCCtU+TCfGG7r
Mw1K3Z8aRTI0DqIm+i6QShhtiYMcZTCbJ1dElXqzQp45W1fhQYAX0J0gKR0uvIxK28cQ8PN7WJ96
ALENIs91kyhCx0WTJOg1NjfkghONFGP6y8xFMhGbqDkwL4vCgXDA3hlFFYyRQueTnpsoBqxdv2Hy
NYPPAOlIKjxPMPA1R3RvPE1HSAeTSOHOmuLKsfyjDZ8bGLTw8ns/GqVAsTSqIbuH7qp6TUeoLa1c
yZWVDQMadiG/hgbSmtdhyXFQj6jDZuufPX+m2hOUk3uY9h0solub/iR2SKZ+UBgQBQcNRFVczKCu
MRe5qTUYepLPr/m5hI+OtB+1bWbDCuYTzUkEV2IKFQnc1tk3/eG3FfYbHjNlaCqNfK2Tc6E0Z2pZ
2M0vikZJWHi1HtUDkUtkypCsaaOGEuHDVz10jxBi4S7dhkGd9rH/EOWb6r9HDGwczjYPhu6ghkvY
6tm5lN89D4TCksogwQGObUO8gvnIAEnGeImA+EWyjtfF15BgH9uGzdEQM2B38mQsb1asWNdJ4iTc
PPEkh5EckIBybK2tnxjzv0RDhtJHMKKePD9C18MGxPa6QO0kPFkVIYQqB0uHuWDtYiAM62+96KTa
kjEwnY+C78nFZagG/gV0yYvZCprmRwLwg+vJg4M8ShHEzAFN/ZZkGw15BHSFFx3V2Tgd+Sar1GJL
/4/liqMJpxIxwEHedThBx3JMTPRx5MTsz2sBiYxqZoyKzEaF4EzXrcQjTxwlBegEPX754tZnSSJS
kD8yWWAgByDPP63Enk+lfQOUCsIjSOTibG7lY/QbvpTlu1Vg42+Vg2FHgesBPrqZeWI/2iyWJcxc
0G2Ves2Oogdtk4JP/r5w7AHhwlHAYiNO9Re/TI/vooQudph3U8ltTte+j+kgKs0W2I0Gk0hX2X3m
XKtraQHTedrRWY9IkdjrMUaRaHOpG7ZbwfogEjo6Cxb3ad3/1zHs3nz+045llfV5XnuYwocygss6
O39UiRq9zSYIGGZhFea6C4C63TJMQQ/ml+76hIuzAJggwz+t1tjgBGdpWtmrA9mjsJX7AhnkI5c7
NZE7SVHj9D5r0G/H3kUS6mFoP5uM8dWCcVDDL6lRVtW85gb5n3V1ECvGZvmF7T7usKc5BgkJDxq+
UEcGxBIyfbJzFgo4SFfOFog/N2AiG7jUJfJhxtacLYJtnfjD2b9Ai0A044RFb5zu8kMqxkxdNh9O
Arj89eebq3Vw1HLjfc4S+HTdckAnVIdwMN+aDqUQJ7HNao11g4ceJTr+hT9LMMqP8XXSGGuf/deq
9nLcT2WxdO2IaQ15oJxCPEC7yPl4fANHAuvrA3NDcHozmSNLs9e51ZtJfykL8lleT4F00UEWCbw4
aheD++43WKWUA4Rmen/p5H/gomAoZVSGJ5fPBPRIPnI6q9jxVCsUPC1N9XWIIg9+6AD2bIKhSzDq
G40LrCYxCgjYc9TsGwiAoU+Pt16WJrjdeqBHcCjAwazyUm8tJFYFoh8DfKGtP/p9nvqipobaOM4c
Nl0DTibkTF4RkwWZXkFDEoHKSP0euJLgG0CUvq4kZ5R5cElGnVINyTQqfJsQ9GinVdQHGzjV0Fq1
Y5ba5b7wRqFF1YLnyWx2SVHVjy4PNEpciYBgZzZcVV7wFYTVWLzGktvKSULZfaNISncbwIVzxN1Q
X117XlWX7q1Kd/UkwliN4mxYVmZ3YbJx0XlfiicbVo+F1Zt0hWnXixlcB8aFnbbngnDiIUXaIdV3
Qr85xhH+cqXb+H3bsvIeCHUOfjs0mq2AjJHfYRdzr6cfGjXHdsWpgDCQGTiJ+FNcNkQioB5EAlvI
jFC8U3A0T0yDu4aHZtjfbJ1MAoiAT9zvQUBioo89vLzQgJ41k6mFa5Gzz/nciJMtYoLquVo1pJ8m
9ie86w9VhoyraDNvp8JNPYN2ZLWzd3iZC36wvfXlxwCzqEIdRfN1Hql+B51nPzy1ATlhBtU1zOnI
LUX5ty4Ph8z2wM7LO1uaGhXLk6Q78runo1nbHk4VQVaI/efauw7rZDTHbrNmrIUccJKTNBLe6C75
lq1CEGo38jGQGVtT5D9GZ42Kc4HiPpMiPuwX3VyGX/IudBFwHKMxMqdm28LfzE/FwfpJ3iBVWpzl
z0tMhbo38SKr9W5sjNSDPO5D9L2KETomslfpqMQcuKnANtVzmorbFXUkCEzqFyvw9D2KFwhO4L3+
eW4wbQu9DREFDfzsoxQU126EUIsAJhU+qvj2FtYYUwQiSH8oNpXdd2G8ugvMcI325KMJoKnTdjPn
4cER1bf+5shQySgoFSexDP/J+rzzW7JnHBYBqOCJ+X3dEiZQMoUUBK3SW5B8L//YkeUG3xMwelGo
++0JR9aeXiaA4O+Kp9aJOrmKD58TUjKU0i6B/ec4aArAwVWuBaQjIV9h5oadmQBUwZ9SMgOlDGAE
D2C/AHfAQ4SMxUq7vVxtqejpacq5IQxHH8jRtZCcciN+903CQmw6FVLO0Cmq/udhP3Kk35pJ4q+U
7sFs2ITGpNxKYgqhsO/878yOdqV4zZaUAjr8pqHBfNpEI1kdIYjlmtJMUzXeFG6NP6BqvIj2bzKK
7DjakW0MvtJ1d5WV+qWCpo0AcNT+Hq5SDCUQTy0u2c8EuKm2agQRaA3c8c3RsbNCJ5SsBV/ynzUf
QuB1Q25QzfeIDzsYdP8IFD4CyIqSy+KvH7Z2hfIGY2zeHcfg1kcIft5KLxwO/o1Od5RoftuiEpJe
81W6KywL3d6OUdXhyQy51ZCAo300U8DixjjG9oTHdcevvcYyvkNgXcwc8HGilHj3lQhjbM0h7U/F
VNBm2Gw3uA8InPJ4P0HEEme32GyKAnJGzCp0okdtSlv4SaSsvzRxg8ld91HpuPMIlLPmZGfuiRgg
8vpL1uCvGxTi3soJlA4OF2h1V2xuD4pD8205r6KRd5rKw6JipFJWrfYtKtyeFFgC27NL+G1a2sBw
svRV5WwjEqCAV0Vj7uDvMfatAGVNF7mAxalyBH9VSLEQTyo8P3DOCpzHHmJCuu+4x5RAgg6uvXov
e03gHoBRE5xlcYPLO/vH/yH//5NglZ2hk7HmEYp4mshX3DAwdLmMOhuQ/cFkK++PRqrm5rWroCSV
OzXYg6dxuXOdfFL2c+Xdapk4IXIjT6LjbPA7gPWemwslV99S+6zqedEGHnG2xto95zl2rHq6ViC5
BLoKbFqv8PAY2D1PuolGoqmUqQKNPqWWVk+cG1YJ5kH3Fdq1GfySlDIUPEa65qo9xxFF/+URHNKd
+WawK1fleeLt3wNY00gTts+0JrhPhM9EDrH57hka386bAnRFi9sJTUkHOSOJcvSGfNB4zV8yiF3v
CbS5J/IAm/zwJISXZpkMbBWy9cb3296LXzLKhsiWS+eklIhAlhx2E5R0tL6R38xEkXGAaKghkmuy
LfuJ55AFm6s4YOvVREAgATRHLRFm+DNGeJp9wWScTCsm11ALj+Vc/Cl501VoX1fRl7Qyc7peAEQU
Pg9qpwfsI3yD70oIfbwmw4jUYUcLlJqcblT7fR6YA2OvOnY2COip8iMXzcW7to2cxEXB6wLPkMHl
ExnyD3GrfHL/815OgUpL7voIHx0WqDninFx+RPLeFsf0p8KrwvQaOpfrxLuSQqhzHCPlKeaWr3kL
y/cT/N+YaNT0yCU1EMwDYnPvhsC33EHz4JousUm2Oev2eXZxmJqiVz6r8RioOF+iEiNTt3UI/9PC
FYxJ1KmygSJ88CXHChqlMwRop0WW5ODstQGzk/e+yvgnIYMYYkF5loNAYzogfzMY0F21GjMGvRTv
Zd1nuxvjJmyGnBb31wiWJBB3VakDr41qhMJFjlsDyqUqCHOW31GPo9mscM72hOwu34ZRuJR8lr+2
SvGRNzf4FAz+4Itm3+lZ98HUA0BV5oW/DSevFHeI9QiOUaiBL3tuI2/MU7f/eENVOgSAEmjsw1Wj
Q8lcjc19WtZJVbiKjqOu4qYtqZwNbHe33ztxZCkyOguOmpJLTfGvLUylbJ0AHvNVWluMQSqDKVGb
5edJi0HKg3nOqW/n3bT/mgLTkrVpiXo6eB03jTFtkxDYJ+XHenrCmFhFtpWlCkYm1p8393oNtbQR
xStTniZ+Ey+TW+J1/IGsw1oX/a3U2nWJ0ei6YEd4pDpsaT6sr6ZLBW2gjhbT0QTKXOZYIaPvqonc
GZbP259bYs/eHVdfhjlJC25P58xH87C92a/cfm6OHdLumjsHv82LY2EMRhsTF1VTGg9r3HYtPXuP
Rh3HpNgH9/gMTnLkN6cIzTvnxRrJgNjWJ/CCZ9R4t99pWTA3ww2kvvQ2hsJndcklich1wjg87Pe7
UG53wlORIBzZ9OCvBhq8NqdaVZqfXwK3sHSyYYmPo+38sn6zsNFeAzVvopw6qY4ImuavCQdNZa9S
LEUK7pZMWKnEXHY4Nx8vzUiUxHu1yWFWyFZQ9Iol8iYGt8suXlCOK9buewj3YPn8ef0Wqpf9zS/8
6urxmcoKsKTMtjRxI7SUTWgFpsNnLQgG+5bONWHDzwLFcFBacS2pO7GAqmHHjtgCDM2i9ETA1Efc
YuehtprSQ6Q57fee5qryu5Gtq8Yn7zTgr8YpNTIWnRIM0shF1NpH0ma55Jft2Dxbs+JrF7swv5gB
qLjJ5ua0vILA4ppeJZvwz8wk6tXJGRe68nNaPUPq2RInrqCYktuZPmGWsrfUOVbfnR5rRCylwfKa
S9Lr9E2dYHt8wBhvcZIBvRhXGwWP3h1pCKo49HJvib0r8T5E27UGTR1FkwbRAc9M9Co4urj3DO+X
vAk8gAXaniQ1OtdnXF3i0in9tgJMVXriyBQEcpYOqfrVirXnZeDNFTgNcceL9tgOx1I3YbUv9Shl
PXBpTYztrQdH2xfqC3CzGsne/z0qvGlshUTd3FOLaEf1fiC6O+/UU5BlUa9auylupMAGQZLXgyL3
Ljj6NDiLt7ODAZ3F1KiUf38n2H9MHJVuvu2DdEkHihFYMxcyDt5eZlyBxcu3Z8bHYs38/9NwkWyw
KTNFbhFDLkwZIxHQC4PEg75vwBl3Ro+pLBuGa7PUnJfTZFT0qWqFFgae9VupAAIBHCwEY9T++8tE
zi4NPmgIbTTTVZ/U8O5D76y1SzorMEp9nvcABg22bvSCZBD3gjaXZuYV/FbsFQfpdlThR6QtxVsB
t1kYfEUmx+AwZPT/7QpSpGJLrGZI/2FLDNrW5E6fJ9YnBy6qy2hxA/zCbVB84nww7FkB3wT+XIJ4
m7VHOb6NSotqBp68J4Vz3/mDIBhLgw00cQMCNNjwhBvh/vDk095geJq/SOdFHo0OMyNvUVqLWS29
uiMgVAcHMaOjkX77JFZPg/zAHQD9SVGBmS44sMCZba/0trHIXN7iEgm0W4RUTVneYRFf4F+IQ+EA
9IEtN/JlsUPWtiRLBjxhqA+4bosK50Ln+jd89lodybd55f6hiDUNzHdig/12+PuynqljDnXNRyXm
r1oRtET/e+A1q1V8uVoXZxsknXF/KoYS98FTJhMeqLlCBPQWYXqQFosDBsZPCQu3erQDkO05l5DX
OwJ7oFySv5xZRDVFW2yAEK05/NenK9n+q9Woa1CQuMCSJubKfkk5YnfR4I4LWfyj1igK2JUDKqs7
jjuNe21YhDxTrXGuOmn+YUxCZTCrqrzI6qvNCxLLTEy26mfr/3m/7SZavRx4Zc1yoH6rApmBHhcP
uKLIsxqP/3TN+R5gYvs7QVR9lZ84baS3ZnwCjVKQk9AGAszFVuitTooFXrrBWoI0nyCC+6NKdcFM
w/OTUEPT4wIYgHNp7o+Hl/7nRXtqchgExlVaBnrbjDcYcwcAwYvOxGzbgUCX1dYzf5Mw5taGc+64
GSkFgDocGjybsPKo7m7qBh6my0V/BRoQPRYRby+DsmQFVkCs0UD5oM/t1mCMT/ZQCp+H/nj6yk5L
/vVIb7RWy4TsG8zcD2yaJLI20jtz+t5LVFmmmBkX3Tm9/Z3828Im2NBn1eeMVZGz7jitJb75N+80
Bz0bSKRhvaiA1Au1aO4/vYn1Y6z6qMx4A/Cr7TIJmkXieT9SIRfoe3Zv3ywz3EAbrfuZIzvPBXux
vxK0RSZnQfEnss1UQBJBqTVQvnTcM6atIVo82O+1ccsmT7lVeVmq4FjNzomdNtu6PvfKhDwyNvZz
Hto/59AOCdrQJilsCRxfdFC24qElpmrsbDWRED8Uzo5Ag3c0kH8kKtOw3xDq9yohYA1qc0ZyuBQR
ydbCvVhbmmJNTgACBa/uWhf0pCpa1Gk401FxP/d/IBShx6WqxmPl92YK52EjYjsehhvvBU3rp+hU
uq6mpJ53ckMXjK8vdg6bKyQ2c9QpwtPQZ84tZXbxntV0cKZwZZDap9kaK+YwPj1k6UDXhcGvldhz
nR6ZAQcY5IxwYC5AvCyLE7ARrX37tDxIKz1/MWRGYNieOLIlcxUjSaMCnLwWDJ+Zsrgnv06WMTpk
aBxtJykCDIzu2uxeg36VgS5CLXCmxc+wsOhY3wWAbpzPKo8q2ux28d48TqYUzGNegcXmtjQtkFTU
ZhF8a6hK5hptWZMeFUydAQ5l2URiPbi7XKMyRE8o1PmSasvLX5tG1EE1qiC4vVRkwhaq3g9Rg9y4
coB67iATRQG3PjqAXS+f+jt4Wfix7OESmj+q5KMDdhExGRd7EjNOBqGFqt7rUP8ElTXgtIxdmrVM
g7YOcGuwTN2yrTfI1/2VjWpCu3WPfnCCYM6EgdrWHiLupJHCA7WZRmK78nxcguzaPIANAU/Y73bv
DXBLzPXB8ZhQj/ex0m+6vlek0KE9AEE7SJwpmf+ar4lGo4wqzMiIlvlQdqCnHZUagCi1FGsWEYi2
UXEAQ0BUQ7hyDKlj2Te2K5GhmIhOJPVBFFP+DNnvbH6ETb7K4XpENXrtoDNAOjPgIAshzhxDO1u9
GMFAiiSIJVMeUaY1JszBI536URk/DzSJDxv4NDL8MjdbwcsgEZfFGtDm6Ef3AVTlv8gDQFWoKARl
Sj73psMi/KEYE+Nmqti3pO+WABd5lSY8EZ3usIlerBmMjIc9shoeRfFg9gGA5kb/9mVlPcZVf2ok
MNktNLk/ft4yMxF3P7q+wkHHgiWfB3BiXkrdIbYhjdPj+T6kupLhPvdZqsQrLE7bJq5F1ZXKl7cr
QBQjN7gIN7FZxKn14G7Vv+nJTz4CLOilxxpdcZm9YFHFFY5LDOk4uALfyUjo3vkB7HAaQZc7uEoZ
OBN1xFpYeihl4OSahp8jy8HI7cuM/b6G3UQ2Ez61zKPxJdWB37Z1Oe4tygraq8qtHT6XOPk/Uy8k
gLaPTWsHw5ygaT3kT9xO0cEcCrxbHU7k2E1H4MYcz8lvP+C7hPaypwIUdI54Ut72lgiHF2Jpb5nF
K6J4ZiUaKczEwZOkEg+EBM6pwPQmfh0QGgV4BCdNF2kXNVD/SjkHVsro3za2EBHC4mxlpEsmCT7N
sHLWR9/QvmqqQFh+TOwnFzubDi4mMZNqbA8nNbX+Zqyg22E4i7WrAqPspFTFMTxl+1Epurz7ol34
pDnkXiajWq5bOHkkwIEQNffFqlNC5YMtD6ETS6tDj42CPSaupJ5asHC8OkmVBQYkG53lOlwb2Xx2
WCRJaMSCMSRpbj2jYzpgGFTeTPWxb3FJ53RO6V59kN3eLNIzAreqlhOXCNMXUjoRhutOxLgtdtsU
9ZwJFtwStHopTSIe1/REcWESbC1jXZ6CXEDOtwzx1odJ0GGJEDOAJZK0x8IT53N7lJrbsQAJdgXB
MunrGiR6jD5N9ccnmynmfxX9fGifrSc8la9zwZtnTeVVl+JFLDxQdM6mok16uPiK/Sz6CpcrChNJ
f9DECMiLKnvT7gFbHH0E/VY6wlytYTwboWf0xO9WOaAR/R1ULU2n386HJ1rvD3GP5wjHSXAmIiB7
ZxAs9Meolb72QfZ8I4VrQeqY4w9bCVlITEJMQxF4zbvRVFrrzOBA8zd83lEV6eYDDmI5Z25c502M
0w+qYTrpwfBzfVjlkka91NZN4D77dt19Y9dKGURZrSqJTJRUqjp3GFr5sQez3Dj3x3oKpw4pwm+W
49aiESbRlOiMy3rVfoW1FBiMpuTjMtXOoLtZsTWiLlF6/Kip+JGt1mTSIpAvJuABqwa5VtiqcWA5
GraeoekXWP3rjqqtPAC2ca01feueFd0gcsS5VTZZ18aBtaxJaCkmSsp4EU+5DLu9P/B6qolSmV47
jDMZO5Che7S5eK0Gz7bw03uTBef6pbD8YZPbuYRH8yNPetKJGJ2BhQIMRS273gffFgoPt7t3XHm6
76FT8ArAzbS4blIrJZC4pYRCCCJEDdKqHM4XTv26VB8+6h6v3YUyA45ZWV0v1jWzYAdYwgGFwKCj
w+rid3vKSP2gxR99CMqf6LJE/KlSntfO/mrVT9KiIKM8cqA9MT0QfEkI8cLLlZZPoOXGmQ29x6Fm
uuCs3Y/03aelDCar8H689xARtdb4BGXVYx4u/X1fDM4NupHi39JkdDbpcqoDKGhJvoXVrr9nzo34
22Tf7TGsyfCbp6OubDImQdtypEQETgRkF158d8CYCi/kL4ZRbrhlsTdOFNu5hgl2awIA43bOYgL/
hvf9LBjqM8HKhf6rt8xzFReEqRcakT3mEMb6ADD36irzd0sja3bitltyBjNRcmUM4DLzt6gTqDFu
pWGKjFA+79JrsfRNjztsSIJhKXWYuLeL1q5zrHONFBTDNJa1WhzS9+fMsS6v6LHQTIf1n9gbhPmb
geZkNW+7V7TtAzAx/YYNNrAthorJTwY7o+UI0j0a6H3RSsw2FpKAY1VA3/0w85c8jBXeGAMFNeRN
ZGzeoizIRJIy28yVBz8LlZyVd/O2L8nis3fSnTubaYZxeojibfF5WrM3QEZpcDFCven5Tt32hiKd
vmC7HHJydIK35XN9ymrzgdhpbD0NKosJtpx2EyxwhO1pLR24tNI6In1mPB/yJpqVKtMnIpEomGGj
F6e4pg3CdGDRgu3fhf4Sz8TREMvw9IzHX1/U+ERZ9+UhgtvSwruI6+chVMdN5/P2hJWPFIUY6c/1
FO99Z44yKKAvBSFk/zNfy6qXDecGVahAjSDa8P5osTMzAsmSO4XzC8Ox8JKOPm32Bm4TZpKiyYIk
zZ9F0RZyIIODAnSMDAo5DChhK730pu8c47BOUS2biHklSIg1ykLp1sAMIBhtRS/r2prSUb4cjVT0
JiL2PuzmsM8C1eOuUUU1h/81vpe3p4vFdoHbn9kIer0U8wM3opu0qnXUgo15TqJQWC0emwZreEIs
gQ5RNtmEFFMkD6H48B3FZ1WvOrdLYFkwdoeOtvZwnJvkK3kp3D8S/eZb2/XI6wpLFL1qq4lUWnsC
kGDnUdH+4fJF9CdEUZfiEJ8lOwKQ9Hq+dM9BVu4HcqlisaVMEMys70jqJiBQ5GZBPNIZy4udY+pM
YuCIxEAotoqRVmpGCvs6ctODgpe+e1pfJjN3XhBG+YIajaUV4BrHErnpFnTZq5wStwyniC3lxlY1
yGOgq6ME7LaNCD7eJkc5nRTdIDrIUS6oc5UM/gad7yFigv2cYuk49jaFXEcuCwHUTKMi6kaZJ0XH
S4I0Jw6SYGxsX3ZFqc+iEOtyjquTk7SkmVS6Nzt3GaFjJ6Uxzyn48LJcXDlL269z+TVysjHbfMlu
+uf+8tyg4h4vgCFTb0n+8c7mowjHn+QCBRoR5UgiCu7xJQRFvoVKBmN9R6v5AXICxAu0gzpIx9I3
e9EnLG0XlTYDWhFuDmFmTsuFPgX7e15NdquYlNF0/R9WpV1VQTtvCNoTHXc6Z4VtzL/NawnDmTaa
gAc11UJB7zLsG4hVqPg4nmYg94g2vgf1YwgFOAtaPdDwjCkNxDspJHNJrHlXLWMivNAarFcgXkvA
aF+ZkY1Ttc0uSkMWI34i4v/5FTpoSB87PLhhCLgtWcFwfFQgMd0blndyiUc9p/9NVgDkJbRkAhnM
OaPdarXqj558UBz2wIttJV6C20UQECZLJv4j705iodLtHLPs2x2/ox1d/8S4jiWQyYD9Le3f1aOZ
YG7kAiisO/2tS1TTDT+7BWhRSfGsRihb0EdJkvB3xdaeyJO8UqGJMmT+I7qqcnV1BFHjXphz3cTu
wOrBYcLW69ZD1ZFV/Bat8DFX7stTOZfPFQAB7WuNrE9hjm1g1YHRLQdMHNZU+eOecOY+RYAlWJGx
jwUKSwr7NsZpvsE9DtnTCv7WuPvq3B0FziJNoyyKMh9uEuFSrqf0ZSGkzmEYGV+nURSU3OZLSi4U
kRSIgIs+4oYWfAVixBNQXuj3Puf5PSHu0J40FMY7RMnmW0/YgIlA/pjp7nhVNBBrhIGsfUfe6NuE
61iCgiDDQ28LIOlvO2X2pld0X0SGXm8q8wwZBGu7xvUWVtmNuOX3RixVUntOyuNYkw/AYArLyVei
XMF0MzAm9sua0GTJYVm94GHr+UJcNR5Klca0ufApDCpS3gpprshBndl+ZW2si/quddlCISVUQphQ
Jh9ZfnyPy7caMCrvVPWMaknvZznvox/SAnWU0aVInQGpDoBCNdPh4kJQzVds1i4wkFe+H64AKtJt
WgVLp9fpFsDgLsOpPLUQ3tnt4jAqPleg7Rn0gGABJMcpKG7hgOv0Silxz4lgpWmgD8nx4iBXnBpW
sw/yJtQsg92wpW/7A+qBGCHZwL5NMoUHmHQqCiXr3d6ZeYgO0b27WAtSUYY3MR00CsIBsXKDQFIE
ZDKcHjlbPrJGyUbbjVtTCKVwyBLDcVBUKttZ/PSNiIAqpcdebR1ATDeEmbgVDzCB3GIzUPiVHmPA
ObQuk+dB1oqsMWPEF7IvHFL0cQz3JMxWjIqi12COH1hQdET6ZBLKAXQwIZqhSFqBxzFPGl+PKxop
5zDcCCjS7+65+n7IpqRTHsdtbBdGOhkT63pVuk817PlrwH+b67LZCVR2NgYXLt4mhlMdKex5hUKt
EEW6xdkt04tTCLLYKecLfHui2mOqkwJEbn6fr5aKpN9peF1btyQAH7UopdGv11wADJtM0JJeMhpY
ijNAnZ/20TTBrtBj3rx+APZp0LoZmmzLitA0Z2Xff03ejjl/iYb/lr4EYP0zhZGvEc6VhrRgtiRP
mt2ofLwMUkYZVOHX5GkVkEWDg7aHi7uBsup86ke5GQ5/v+7HTwj4EjffEW8iXSuiWCUZ0TTTNBXo
f+m7bkiFqsEX5rHvCprY9OWqWX/prgYm4n4N5qoDkUHDi+8IHFMn+CMiBAD8sv/q8dcxTzJCZaz0
06Jv0LxnP/MvW6tWnosm6zszu8h228PO+hCVuMmahEoXdAKduOZvYFDm2PXBwVRTMlML3qDuIERx
l6UvyHxaVL7C3ZA655Sz744YqwFqIuQp4fIva/FG5naxhKSQ+g1iTY0woO+gRH726XLAUXLZ0QdY
HiQUyiqV751IYUswhJx6RydaE+fKQbKVxH9Vx+OtQ5gznRQHw7NCrXBELOQfpmbW0vLbTVUmmF4g
ZcrwfWwGvxWAfWsAIJGKkAxZY0ec8E1uDjtPv81w9OJEze8C49WKByiwCVCsvSrHpP4fAZ9PBi6i
A6H8xx5uI9YvXuLhz+SlZY0Y6eEgdijen5yscK3dbP0swNHB0HPhUFO4K2ooOAY6U0SZz4vpuaQg
fX5cQb+SZLdSK59LPOyUqUSa93BqP5PJopZtlsm9qTRULpvBKAOff/F9KnmDL4qYCY+mqM4gpGqa
bCPv6PrM7gpyf/9YeXNy5cKufzHifhJH/dc14BmnYqPgqdYZERNNsrZY2KRxZgaFPahlVG88Phf8
d+Y/KmqPDRDd0fRvlqDWvH1poaPpXr2ZugLvic5DrKFFCcWRmG0HP+zPlSphM1me972LYifj8+gW
cnB7ljGZeK8USlEPerG90lIUW1x0YO3tIWJkasqXKZW6f/nISQ2jYsRNvh+0HDgVbMgm9fy/kCRs
lTL6LKkFL85QdzPo5edrQeZbPn13/sai9wiLVo8Yg7WtWryE/CjfEpnGyfWB225vGXWMOiKOQYKY
D3AAztDDaHzbhJpdrQSgqDEC+MllVkafh7g/C94Qzp0HCtWx7wIGH3zNtZVRj9T7fhcxRxJOhbJR
i1P5Xgp1VGctZlPBu78JdAE1M1rm1BOAutf5x1K12znn8jOo4VisXCxvEJOq/pT/N2qeqUcofh+5
f7Y7D3jdEPWi6pAv3+uAqo3bbwnA5Cba3f2Aj/fEVEwskmLmUcdqvvrsKPCggEJijMfRlMfRZTxg
CVv3w/vtbpOj1is6XHhN4aTMXsqU55Dscau1mQZ5gMqmlPkQLg8uPaONiLXyUaSBtRS+wPmPOl56
oLpDZvN8qOVs+/rm1q5IAjHseMeS8/wUpf/kArDr/gdI8WERfx78I8SMfcXZcS6nyy7K4355D4C+
uG2RD0z4StHt2pHY50SWJ9AYakSPavlOZuYVTpITl8tFfkY4AmOqtRvWdVzqyeh39Gf9QGSIfMx0
p18tSKegqhKO7QtfkE5kO6rNPjcP3ucawncT/1s5qo8q28PzgWdg0yo5nY3uQCJUFYzcVyNQnFHJ
eUGvTzHwXy7O7nWLC1ddtB8DgkZ30yTkLpMYvwnzUU0liyxGn3evkj/wBo1b+Y4WhKtNQ7GRmfTY
ZbvoI2xmumZInH17XxStZ5gPFJXYKW00HJmSug52Tzxx0+ClIHPxtsJQzcrD45efJspzWiwnU0Sd
yhScOI71xUibm/fUDU+elLuhBaBw5rY4zsDe3ONRlFZkQVHknKSv/kYV9cvzHL2YCF081JdiaGCT
xusWu8VabWfdbDOC68STXYsk664KpEnXvmuMiZho5GDBFQ1tH5UimaAxvgMmiEtloUaUMbEEdn8c
rHM/3N36GWOYE2lsDKDVxBEG/MGUAL/O8YxGJ7VgzHr7pHCtSrpvzr7ZiXa4MeZDkNWgIHiR54dL
B1lHySXhbB2kgDYXhXGxGyUONvPVBFStUitYwvfIU3fmR1JUsd8RplVzErZcnL97JYbo4OIoItLj
aERfy/sdhbZ8CyGwVg8RNI+46kNwW/532mQqgO3wJifvqzYlPRiLecr7Z6srpmHi0aDBAQl2gCoF
uVyKNKtwXNSYN+pf5vIEIai+ckM/bcMuMG3sGeiALoI7Wiz6hCEJ73Cr8O5HjLEjmho+G6+XAzV9
teD/Crbr9akG6FUXYDMS/0KTpV/mqhv4U9lEqUuE+n/a9MvKqRJ9nCojFsyhi/M7rm+S30oHtf7q
9ZYrNSFx1nIDHevcvoSVEyR4tawNXkIGTH+rq7z2DGhZoCwFqzl6S2jEGbhoDETlwPuST7qCW3n+
MJzba4WlrzdHaYHS8PhUZxyI3Nsoyj8PNJnVxhdffHu3q93ig73kfurps2sjJVDJEOMOronUmtzr
8F0UARH8ZcFaWHJMKbsSoZ5415qOsuutq3khe5UaTcDuSWMPYbOcZ0p+kMXgLkij6+QTpu0fYoQJ
PixAv3xxu1qjC6op/ti74XmfI8WwkKNQ1xYGNYJqjO1Ln4bIPg6ur9+Szdpa3O9kOblZgVKqApJ8
vf9El7eoyiXI/3OxZSlvno4IU0TZpFltdDhwvkKB+wxMutTQNfE3F3uAWHYH2d1KvlMyJwXNNKWv
WLZN111xeXBZ2KQa6H7Ujg0/SzmWSj5ly4t6fHHa/6zBTtgmU0yZblAhdZrnkqQ4uKBoIj2myS6U
AsDXZkNx9blmA2nbLYIR626tpgDKusYR624mLHVBvrs2PiS3weLNotEeh+wVtcx08qpsvbZlqwNZ
YRnBDXlLCi54476SL32V1LfhOt8oCcq3cMlv5LOt/vKcClrHGkCmAkRk38WuVhCJSdZYBo4rEPnb
xWKdCh86FxA5nzxdNOJSdFTBBwiuMKxwS8ho1qEqHvkCA7AzQSGnISj588C1MY5VP0enUCbXOlPd
3Z0k2v1z6xmEhrnVwJK3nmMIDL//nPbbx5Aiah7aIu+aMqwxFRv3MQYmeqrK+8ifAw/R6W69lj65
/udxKerq/SwCWRmj5RkvE3r4lCK7aZCFDYBAAlp5qrRio2nuiPutprIfjRbZ+TZ/5CFobKMiRvGC
M2uRl63bzsTLvKcmcBosiBTb1GD0q24RFXVNUOYGFJak+ZNF2IkFvtcHh3LR9LVZ+puCucGvTAXv
UICOs9FNc4KhgjjiLdsrBIMrHcWuu9V5RuwZcE01sYeLaIVk93+c8QZ7nO8OTTPOgXuabv/3ap5C
kDuPK/rK03eTSzMx9+I1O1UL4xH6Tzi8lApbiPH4J+Pvxq9IrUEtJ1etK2gLzphUwZm7UscMeKiw
nc28AI18upcPlJUO28UzZxHP06iKGMXBT9NOkXxpTwCPKcM/bLQ6YGoOKyUExmbmUJ4pmxWUB0an
AbRI4PnNs2u1ROjd3CWbCgV4XJ270YPenLyOT8Yl/7m+lBLDPTFKWmtJ2Q/jyU+dZXXTVq1J36Tv
4CokE81Yy4sklW+DWjH7hpauFFWqDvjw2roSlOSWdFYswFOC4L4Tn0qI1JVJEcjthnS4WJKCjHCG
Z5iNYvFQgB64kJHomKcqzIJWUzDCdgYF5MtjPn+i6huJtAxlaQ53m5hNjfMbOSYnOQ+PJWhWg9ga
WAfuMk0iJCRRWrk7iwTq2Q29b/cOJ173JzXlcNpfj/6uQFYZ9ZvsRm6ZnjK2gbjTHEcVkMa2Aek/
mtF0wZx0o+cAkEDBzv1qC0xZoMWbQIgmP19p7qrm9DUFgVc9meEkn9zpUptpgKrgCwGl9qyO1Cvv
wHrXUIEEnXbdXdOSwhNri89qIdvFZYjI1W9E1/JtU0V76Q8MqkoOE00Znzc8t2J4h0uvEJo8pUg9
kWMKmwTdfe+yP2LRhA4hm0Tf8k9q7qGY3HcAnsGClxK9QGIGAP3b1O8BZMt4OWbVhD859G7KKAJQ
RuUhgTW7Pg+BXoP4SJMYFOEwIucMSzQp2f6roaZTaw08FoTxONwfC5JV7+VpXA7YG5ps7xA5+XdY
Y3VCQrTyKX6b7SmN5YsvVhCvAjBFsEJ9DJQUlxlFXR5Jl+MVlZPnz5ynh12xfqmjASmb2xM6yEa4
+MMuA57M38evJspmhuJWsmr2GH53r76R7iK+8zYoHCOQNWrmQVSFMdhxT0PEaiWos+fzNX1rsDmi
pgjUQlB9TMm5EV8OVJiKXSbrzLvXU3+qKl1LK2hg0XaZYjT9hZjOsjwsPxpyb66vxvfBpe0BXpac
hfAfq7tmDyrr4HjpEKuyvtDiKab2g83FjPL1c1CvSZUrCcBpiUu0yoWxvmiedYru3uJ4qy3brep5
X5h9TB3o7LXgXtUcy8FYohbnwx1NztOOURi6YII0mjUnBz5Sp9t2YalNCqhdLjwQDaIhnN/SLSm9
epZrSPmE0EN7zUv+buVTDGDPxYOVUfjqnht6iCULgk9UOG8X/aGkRptbDvikxLNfkNfnE1z1glKv
eDNH1s6GedNBz/PMrhAr98tsyiAWdGrbCegJd3vQDhSExO3aNOGnM1fGAtuNXHRxpmdS6IrK/liM
iE398W1snhnur9+Pnli8DLcjXfnYmXtf+sa/baNGd4khWwLqMv+5KvK02c6dfbYH2ZeaF4OScQUt
6v9MMcqxabBm0Tk8yc6QH1ywFS7fv9IGaIJnPBXdgVLgH0IKuEPL5z87WKJxrrt56oP9Aq1ru5NP
B3aNERqsM+wvA7jiKao3BaUXIwJSmPEPoy/STqZOK9S/bBQwa+fWih3wHBmc+/qffdJ2DdbLgTlK
oNvwb02YhPz0/2kQFrdvaDnXdQepSTaeTe2NtW4iIjM/XgPFrA/t1KTb3jxN3d5KFzMZkSbaLStp
FcMaBu266+ax+E+w3SmbvEKXaSbcou7EoyN/vNuNaPZ26k4J56sF4xesRbDI+sVu6H99NtjXViUb
ttN0QRAgBvDpN27pppOy7QRTZrTqMLNfkYmPdJ0Q5ZiWBiJL9WIBwMcctlp2/R9X/wFDEmK4jN6h
6Axyw8GFAXkHRpnCCWuCxjwUWUqWrcDyxfblIkFUbkOBDaykQOcES6JHEZHbINY0eyFDo384qwVU
Tk3v5w+5fNVfSNdfgWiICQ1tZVVOFPyHMoBr2vY/oMSGLNUMGN1eOAXN+tGxjmrNRDcz6qkvq/ET
HPlN89t1gi4MgRys3akq5X5j9iSJ5IkTskkdmzYGXB8Aj2dtlmSaszZWVcfS533v5GxIgKpdHGCq
Ir/OP/xXRVjIrmy3lMQWVIDOon8+4ZkKLlGreWoCld31C+9VckuvuGnhr3wB3gapstKBHdPrd0VP
k7b4IsmGFyf016YS4143Vee3YgheQAYcOdguSc7jTcZfrf8Qjf8jbSrgPqCjUmEC4rLQ8UJzIOOp
uXaMZwSHe/YTxwoB3PYjl6MChzOZPag8wSL+5AmYfdM3EiG4cQnek6Qld7ZTs6rgEwCvVG2Pp5he
XKGIKx/CdtfFlxUkgmNIDqvl09cmI0keTQcR/qHwsbfCzcsvdltHth04A6/kFj3yzvODDbzmYQPQ
p98rEdOzoT3c59J6tjZQW67egEuaitP/03t7poBzLLuLOBhTMAnjgcBdv88HB6uH1mZawV9QuDae
IcrX2ZlTZ2Oj25Vsg+OeTRR1SN1Em6ixMowMiq5XYcAeNHXowy6u2EEax5e+j0JmqZ/lcm4UPf1X
TY4fB83/5ktU4SB7e5aS/2XlVIm+ASjsLcgobhW2Pm3D8T1KLPVDyuCBsPYsp4R5HFH9mBhZgu0U
pVxPiyter2pr1ANvUr1RL6gGne/R5S7jYjEUpC1ATytK9cbSZ8JVvCX5veUsZC1rERztizFrhg7T
R46yenWj7Ll0DcoBw20aO1Yd8HTMesc6radLSY77AiE6EgzeGyckMxQKdpaCs14DUGVSB+Lp7NiK
TDBRnM63KTwaeuqQ534yS61FnvoE44NR1eYDP229sFg7MgBxjqFk2/ar8E5HxZNysO6L7oDeqvmR
czLOVr8hJhZEkYwibG14ao6564RrOz7yPUDbmnUDvSruiscJTsMSDOmSmIVXoNSfG35XT/SEFiuk
941xy5ywTec3QAWcnq/+6Geu9jGcjOr23NJnDJpcYEy/QSy84Ev/1WSWnk+6eckskbH7FF7ANB8I
fmNkHlOLyfG9IXN68r8VyWzAWJzVlCIu5rfwVfiybeeRsXwmSawVOU6MXl7MTb9MC8msuon5qs2l
4CW9sMTZgU3RwgNyjRzZeEmc2QAfbZW7i8ShDtj+Kvfn+EEmO6pT0hA+2m56ylcZde3q1m/mIYDx
YPHsp1QufFe8V6AzV6/LIQCnDmlp99xtncDVPtZ8sCAT5nVgdhQ945TORMeZ8W+W+k+J+OS1q8iI
WzKw3wyHn5PvaK48UYRq0IcG0faG55yY4YyI5GvuLGeOO+fpDC/3o/AkYjNXP2rVZ7fYy/NynP8q
qAfEk4udSpTobDSLjtxpw9QVviWi0d16iWzFrsKgA0xKvdvX8NIkk1+p8s84ayWEiqVGSCH7zZOX
nBa12qZBDvgLtSxvvbzxeNBUObOYL+340HFoeLyspxGkQdLm4NviPtzSMQLpNcF0fU1FO1+ul666
qbpuXhxZRdkP+AVsql9sOTVrWdSkG2pIieTmDT8se429ITpFRYv9MyRnE1BTOIMYhj2DdI2TftRe
2kpWhCVnWPIY15neUN1SBdmhMn2aP5HcQUXMny5xQ/rTMTqnb2kyabELxZaJt8mwwF6aqfA/+tUb
2bJfqdcLzZ0kFIzXqvw7rx3h+aLKwstHmDf/ERx0ZHCnCq6ivK7FbtyxUNyqRDPpXBtAVuszU9u2
cwBBVvZiFkIZ5vUMts/SPpLzlKdBBcLUKJ4SZQZfnX+k6XEUAsaE+1cfagvbQIbjLKHDrlLe9S0R
qfwiS0j2b0dOlhY8e2jNp6gAhCcwHW/+aIZZpnw76L6ZdFSR0Uam1CZMoQHL8GIadLinDQ81KjZt
El+pshbU/tl7wxZLR5rlzm5Rgc1HjN6pSklQrKU8emLL3cn6SpUarHKhdy3tdrbonXNYZ94QWdHs
LGURkmqZq2CY92sf3CdWRYxgMNXPbcHU64X1IWKYx1g6NBYoSFe52Xx2EW26RhEh0hxIwgThp82T
9JSFSo0qJVXZolZZToig1rh8xNf5MAJ1bSNtHXfVkXj8vxOynsE0d9CDQeffOCddZ95dNirE+1+J
bSWidbp+GGj/BWeb/ew3Ul0IbKasGP4HkWGrvyw/XlMN1YdHS0oKke0gLbcOBNStbpMIr5utwEJm
Ak7HxllmfofbfpRUEM/dzK/oFHsUrFinOcj5wSsWqSc4kcYHCXjucDA5zE7w0R0iQj5ESAd1h0Vs
v/Hg3HhULb0le9cc5EKYVOM/0DOvtAur04xyClLL3enxph6kHSn3W6ggCCpv716/oup35v2bs0eI
+nzC0RjjIyLHHMkdgaGc2ZBEv1HK11jXPN5QCK2IYO4DMkHSZqGWnjJiGZ1W5+taAZTQ53LEyhGs
1sANPK4nzzF+a2JP9ORcpWDJ5/f2sSxPeR0PpOQ2EmYQ0kBrSX5TwLaUbcFhB3Xw1NCiNfSOEYYs
m6CTQLoKaafuobijP47ifAAthW7+YukHGajaXkowDk/wFIqLG7vhtLhoX8t37gOy89FphL+6ItBx
KAj7op4u+p6Rq5llU5QgMqzkP76i9Oi535ikKAoMYizTPQoSRbPnYOVmK1vJVdSbC9m+UtF7lLJP
WzZEuvFhJC1EXgAg5fNgB10+HDK29NItgiW+HXzdd/2waZQ7xb0Pir+jt8xh3vClW7lT8mV8Pi8L
tY7Ns7AYWSrOZloc0W8nvxrzF35KUfKp0x70DzILjdEJbQJEHk7ZcbSwvayuMlVgtnRoQ7X6DM7y
9xqg1AX+qyRV8V5EOl92tcOdbwt/Tzu/nzgzqcsvkQbGlyjjeSsuibkPIp6NZM8DkWFU9FeWl4pv
Wj0rMGa1aFRh9nszLmoa0cUtUnpjks+gKOFF3hoI/ywLjir97ddCM5t3NytbtejVw2WG12EnmsT6
ULWvtw68+b7uAIAhRJhrFAYjOvZPcLzlnuVmDeCq2xapHvK+olGU3kiliaQDSkO2vvi38plP6TO7
04ipuq62AifkJ1JeEuW0u/4z+yRFiD/Dn3oaCCHCoI/4adHRNbJ4B9nV9pswT+0Ef63QQa4zxP6a
GgUhNoMkPStb9+oR5ZlVxcTSU0KeLVZMD5zg0pnh4l+uTNljpT07fI7twy3HS6mL4dpeeNKkkx1D
Ajybvy8wT/PgZHbklrpahX26a0wcG217Ln/qHSwxNcKp91DszucjydI/dCyZ8X1APglRvUij90Qa
ZcnargHPcKlrksyrA4D1QTlbvP+oN69wZ1Tb3MubGn/xsMdigaJh4y0UzSp++S8eEg0Y2x6WGNzs
UP4gnzZxK3VEywz5aOmAnLXdIivjpcLndTUqglTPr2ogCmnBg21K2Kii14TC7cCZ55HKUzEM5j6f
2AsF4gPGmTbvlTNiWzd6WgN9XQ7C064orIuFl8LQiBzclP7vHYYxyoWqZPWjoVlezZQmD8QmyKeO
Tr/S1Rpw9K5hOT71gCVTzckdtJiQKEcD0+RP8alvY/coGgtNJooH2/rNGI+8f26gwo9DksQuA+7e
wRTURcv4CCJZUAwOFM1je6JynlBes46VGB0bOny1J7eD4Of0M38YppGBAWFDhNTzJ+Bn3xh+qPpv
TuPrhzTxC0pJTxcpS/I/AX+yVBcNZX9CJ9O9kceUWBIsZXkXYMSboe+BiPr/5YGnZh0cTCEgWzct
G5rmTCjCkmqVIaoZ9WE0h7s7jikP8OaAfF/aNLGEd6g8V6QIUBxF+uGYEhCwAMNUvda+2GpeGdcp
QNlV7ECc9i1PDdEz24GiExXAdhvfnE/+Z9tDch0SmLg2i4qGVGi3HqgHmL/psiNLUcjnHgsIG4p5
Q1gEJxccwkqI1l5D1mrxp6KtJCg0I44PTO+XcRt5TyeGD+HrcgQbyNdfIFSmvMWR+IXxOTwpRy8b
zuJWH8rWgol29rzT2dkCukLk2aUKieA5xvVeS1eCNJWRonBxdtYGt76p7zHhqK6QXj++rn/nXvs7
91jug7sRioeGHndtoEV/4y62dzwNoslOCkvyVNDFqdFB7jca5M+L/iSHCns9RtESsw04prEWad6F
JYlItUPCHz4WHiSZaw6JIu/Q0BI2Qupgu2TRhbnVcH5b8qVICV1LJ4XHMALASKyASSfDXz23QKnp
bTLYmPh4kq/iJNr25FMvBMY0/DwLACCtlu/YJoqytaUP8A+ns/zqjobh9CF5m1RXN0SgrM8MuoRf
XGu4TMyUqqoF0bmAC4d6v/bfN+ISQO4kNdZeRsHio6iqmgp2AZck3xqPDabOEpDL+8WZhOOdehEP
ilxWePh0Org+hb/rT33pEDlbSlAh4KKn6LHJZagFpIDyyRO6chsO1ET4Tmzb3okdl4n7FOXtGcSS
6OQc+hFpB6/Ek8/iQB1ZDODDnHHgs76q8aHj11PJ1Z2Jsw2rTIaJSz7oq5JowcZ0koKseJp7yrLW
MlW4Z6UTOkgRI4JkPdEgOPJyHUUQ7xYo8pxR3chlLK1Z94Ofxxt3qvLjy69nU7ynlwRp5EVfi8mK
mCwX5C8i/V/T0sNmNSB4UgX4iYBUdmWrrM9+kacnhvXsfsymBEuAXw+4BF+wRoMlffkaYR6tT/Yy
7O6dU8M7ZmtROpe/wFo4uIeJieUTO7/oQ7BqJXBrfeS352up947SY0IME/2EVOZRW6Y8yQQSuKHA
lmdaos0DOTrPZ06w+0IhALmUQov1Uqbp+Ktqk4n3WwHvHDOTeb1TIX/PwHomksRamksgHWNrlgRa
ml94zUz1XkxD5gytPQnJsWpPVsGBmGKSckxYZYfEw7W5Bh2UeQozKP5LWJs7L0m6JinfKaf/fekd
mcAfnJf5Qs3Fgv9kp6cBAAVU7+zcX+pr3YscQ1Yz0a+c8ep9Xkz5lGBz7CQjZEkxwuZyZdpYobCx
JwSUItqaSlZ8awPXe+yGBYUjhe6ogJ3KptB/t3vmejZKCn0ekLZnqm5Fs7lgmWUbS/IpqIxkZuQj
wRSN5uQv3QAJsiL2tYKLY0FetJeIpR1jhmLZgAnQj0Ozsgk7EavJag3jXOnA4suS3z/xDeBWtjs/
88fu1PCaDSZi/yCDFQX+m1ptvVx2P/8PzfaNJX2UtejK37sAjVEMskVN7JvJ0c9pDLOcDnQViZih
6L9nd6xlGJ+TibtKshcXx9p+eM3Tyb7XncwvdgPiYT4HZdzTYB2EFuXMV26dzga5dFIGQwgpFqQX
fVNi4SZdE1XBeDjKUikWSszaqvxDH5m665IowBkQYin8HuSgCm0XzyGlBOk+K7MheXeXnr50j8zs
lTPxgfjmARyNzKod3i7S2VLLJOrtLxhMsUM8+E1IQnVp7TYu4GrBWsk1GOj7nGlCVUt6Favt9QLy
/6FCNd5y2IdSrg5mC+3WDvjuSSyJbIhWXZslkRkhvaoJ2sq2Bny8bYm8T5ZDHjEKUQU8O510UrSD
CuWstdX17Lv5tl23lmeEkz81BJ9aw/cRpe2b0os3FI2IaefoUOkli5mxfUKbR6zfSoqzeLzNIYa/
c1n745EzoqYmUAlL5lcWB0+xZamJQdhMAlp/TSuw40kr8l2zwTiyCHgdCvwVZEC0wRggYL8K3ATE
OZugYdScbAKEulLvkUjG17wsZOqq8z8OSb6ka2W/oPJp0ZSTeUzwaI5DZfcgKvsc00N8GyHu7Z/w
Z10w7CfP7qrFeBRZSeJSVT+n3XKOdgyTlwfBPJc4DUH4EJvBb9w9hZ95X1NiHnTs2eyXORPPcb32
oNQmfq1wni14J7UCB51JaLuDYbSgUcoNIxDeoVD79pzI2kAE0HKLkGhpMrPPjEVXdQj8Ramwc5j4
2pXOz6CvEE5gfZ2pIVFtMqL5N6TF5bKHvlmlQapnBs5AenpdxJdKGSLVC7QYTHStqys4W8XmEun0
u5CzfnuLPu4BeynHSBQXdfazlSBZMukldOWo36NCVty/pMfC8cvuY2pImHn3aGQjgOlkb2TTCz8Q
w2L9Y9kBHP9OoDwCpUwJD2TSyWxdm1fOdfnyCMY6W130mCuHkG5xxOWF64hTE99ZSAtdYCsU8TUF
ilUvwOKfAqjUJLbjIIpFM7YYTw3vvn511UXo3jKByP5R4+MKXA3XiRdYXzttvX013fhsg8Qpx9dp
6OiblX344SwQMHJaocyqUKdyLK/Ka5p4os4IcTg8wCCgjKmjWo1S9iMtNbTNEP8RJvFTwajbH59k
VlDnGDimh2fzBtgW/SmQHPaA2rW7LFYokBJeGhliex8LEYRpNB2vaRvtnv6DSew1ifNQS/3CcLWG
K6Hqrdedx0WxWpUCHMy3fqqRBYBauX6YDA6++7iGebTiwPgJekJFoC5x6I4WoNVni8zwwQhLeYtH
pV3MpOAr/0Ck1j+Vx+YYzw2nC5T0PHBIkxQJqbofutHU4M1yMcglboBgHCajexfEG/a7j1tsB+4Y
GNvXpxLysthTTgis+6cgODBN7bXDcyPXEymcJtt4UOMce/mXivlGzFUvc8h0+wu1MG+RQp8VtPK7
i19S5bCGnTTMqkHVme57Iojg9s3VA5syharH22riwQyRRz9vgephTqlpGP3Nuw/T22lt5wheGCkW
IblQRo5muUK9WDrSQEVa8zIg5oQUY5hiGKa/JV0SUmo4ubL2qfMsiBNC0z6xMdQ99dD8jp1tZYmr
avDy1T6Ezkv58A5PcOGcWbCP5bFVQhACD/VPTjRuRG5fMEbqFBLyV4GicQauNhZ5ahT4UEA1jARR
ktsOVKL4/MrPf5XE8svaKfkoTanb1U9At7xD3JL0onYoSzT6e1MrQ87K7zA6/ym8A3p43JsMfcTZ
tRvKlbnTKZmUBIlnT7WUNu32RsZUPNPdrCNesBY4T4c9QhjlQEwZzS27t2+l0SbXJN/DOEnWgFCz
WMqSvU9Bh2fpVbUujLACTIFBXooAiPQZ1Tq+NCWXqWF0tKk7Kwz0jzbjHujp229OIhv1bPxsqDC9
NWNVZ7BeNH6a+6x8fvPpJ33GQR5L2O2rKlSYs0X1MGMVTO/d8X9A5/viJsdEiUfgfK0mGCEiVX/C
IVwjvfrpFlG4okbWWGt4Tph7QqKN+G04ciyFq0DTvSOM1GzyXDi85vmwAe1YaMyDa2GfcNdBZAtv
CdhRpQuQwhWcvIfhmYJAdbkbBqE/Ot9eV+B5kaDq0BVUZGUDvIBB3acoEhmruRUmfEDtIAv+Jzxi
6+AW/rP4fZ6JiN7re+bQxA5I3rAGyO5w2LWTwSblgwwSEUjp1EHRt438PNi44HDGJ1km7qTE4XEM
iDsfDIpaiWUxs77YHoz8Q6OdWMdQYEs+ZGb/eMkEI3qlvnbEc/OU2qP3JV1p21H+m2sDALM54PGf
oJw55dfeZpPs9Nmq4GjBgo8I4lcdlH/lT3DsEcgdrUdZKcinXEIFaAO3Fuwq0tadyB/fDZhFj1vs
AeJ2v72NXOzWLxxsrT5Wm1uuRAuudolwaTboltz1l/TlMGOM1lVZI+KXhmgVikd/ZUdXkhHhvzUk
tKarNCwrLPmgorm9en8Sshkn2qoxQRbJe/bipbbZxxm9DHq16ZLMjTvY93iFVrmWoK0fMR/QJvmn
I8igkybGguUBJTpo61RRIc/492PI9LRHLONHp1UMY1/tV05N6SDQXdDulVGpGpJeu42e+HlPZgRc
IKUq8MVaE2Lu0iDeKWiH2rEXu4bXApjf+xhGB02c6qiEc5CFa28I0g2LWsfg/ZrQuGbtTJkHqU3J
xcaCZ2C39+Vr/47sdUd9O8X+2D35+GkSSbbSAuoQ+002YOoFu1eyxR815/1l/jQUXrnM7RjMK1X/
lKPjPPbRjdhy9i1llG9YLgeCbsGr8oZyGg9lCKPtXKyra96aowwRSrxEsEbElidQ7Fx8F8TVLUVd
tWV8QnZzTDnQYziHqbjXI9WCnGo5/0UUr4n8g8VHALgXkmLmxSJGT/eh4pOsXPRpP96lVclycv//
qEjMrPmqEAtsVmBdHzyoSXz8Mo4COoexkPa12/wtC6G55g6Z8b/9j+X9hZRt2JgoiJDipdO5hmzy
/IfRdP4jP88UtViCkdatijGXO3UCnLRYR7vgcYU+bM9zka8vktR9IGIMOLkvv1a8xpVNzY+4zO1T
MZ0mpqezBwGywxnDVcq8gaa8PJYyzezqYToY2O5B2q/LojJci5ri8UxzhHrMiwN5I8+1VQ66U2NF
R1QZDgCivieJGERlSWN7NYUBbhfWHFYE46oFwbMBD7GPgMrBi0uOaqMxuUu3T7T7HTXkV3w2rqPS
Ou+d8mJTmv2g/iebBvTK+xHXEb/1PoPWn7r2mLKtqCZNXU520MX2w6sbHleX/RFkEFojzWBF5Khu
3B/G6Abp3mOf2p+SN/usvcA0HhlSLYheyNrQWf0YBMYbytn8EQHlb+ZiistHMv/DA8TLVSM9SYFf
zW1BGTS6MBASKc/hY/h2iLpAsWKB2xNQqDnYU/pfc7z07ZY6Ay2pcn9Q3YjdKfMm0HcPzUJr4X/T
V5e5MudvSJr8VUZEz121uTnuB8IzsiCn4uehF8F9+SDdQZN67qfqiFZxRpQvCBAdFZtdIuxGbrOS
q1HZXU64CLycp1GBHZFomWjlqLNTUM7TPP70z1ReQua/s/u+SGcvMQMuemW7bj7uH6KP/umz0ZRs
Kb4ISGJ64lUuazTIgAQgJ4wc3Y4heNz6E/f1owyekvTtas/riHjTe0cVaEUwjmTgO4zScNGk7R9L
wXfK82N62c/RNfMzlVjAZlC7yRp9etkSlbXg+xniJBDUHnwOWTMAZoP77dj1D/eWEOm07np1QMDS
5uzAmRePZzS7KVfFT9iSUjR4ViInX6ZYO1cLUCJSPZ26JXiKnQdL7JPFpRLK/5FMinRQWDMPzu/i
ZJ3c9r/UssuovxSXhhcQXoDbH+H5EC0WFRAasmMCOf3CNdZW1ACLirRRB1SxvzL3DxnRYw6h2RgW
PfYYGFcQntDgyXHwVblwJyRH0i8BDD/42bkiEySMv28ddJw9FteJH07LpiOvZqlsYCZomju/YQs6
4ZJQKG3N0j2PDQiwlJQqxZZJ/1J+43kGdejJBL3NONW2JtEEDulpD4Bpr4l4yFAn5pB4uV+n2ZEh
RMwTjV57t1YowUeHLBdvOg3n5IfSTzBWOJlXYamkHmZ3f5EP8j8aWSjWuusToo1hHHDESUFo9h6+
M+wTBJWTi+l12yuv5GtmcVmfMUncOfoscUp7Un8uS1Ocfd3IW8Ata/LB4PmYF13zju5IFS5YDnNA
K20L2cY3gNsbNLXFJ9zLBYJ91AhegyQre9FtN9LiogWe5O0AXQ21xP267UQRAbhC//CdTaXO2tsr
0rZR+TU3JRnwoHr/epsRjYNr7rh1cnF63LfSM8rcgtbXms65+aUAByNQU5qKj4a/x8HhpCiBwnkm
uY4YV0u7W0NzLOo8HK/050mIq0dCvGRLs3IFOHQ8xUiB7j9ACuiwELwSRgtXcg6SKjXT9Gtmymge
sCP0V8hp/8bstg36VwpI9/ToX9OAzJ8rDNWnM9O73EEhakCS79Vr5LmprUcg0ZNV0SaDmy/TuFQD
i396zvsSkf3951rMojaE4c2fcNqudG3ddGNJMHtjJ1Wt9MYUGcu0usQGipyvuAStMlg18eyErBdx
ehJMUjdoLCMOuM7eU+SYK/qdGpucTX0DBbacoYp3uRIMJWtwHHtwv9w+F+u5haZ1sl6VLjwW+Gvi
NmIaR5GmunhvC0PTg6LpM3b2gfxVhg2Ji+3vWhWEVafGAqkSspmPhzbaFnljbt1EIEz9FhUA3mzp
8lnw2Dr72AOOhmxA+nntcFG2LuW4v7Gg18O0HRoU8VA4/PTxWo+X3jdMhgr1VZ2YVCa6aX+JqJQ7
ca9wxr3aba4CoBxnhe+leSWD2p9N8AtdGV1ZVcy04PxJM3tqNzK06GyRxagnuw/yYm13RN500OLE
2iWENjmdqMvAtqKD3vC9p/rXELRz5479x3V7BkxUlHX3e2jOjPc8qT97X9DtPTg3Ogr1/4Rxl/jk
9Whtz7STyt2Q99WZwxRYiWDI5fjU3OeHTrsv9GXPft94OkwYyJzZ51D/yDKRu+pX3tT5WKIV/tqD
lwFeuj+0JKANsW7pY9zJHegmQlYNje2/ypTu0FLvTKzzzUwOkYOz9V79u+6WSSTh0JmTLPK4IB57
XU73J5hZvOFHvmrzMWAiJcFD80gkeGSgASGZrdfaq9WG4bJUkpme03wY3VccUD8dHi8384jGIkMj
ryfaxcJh+ttrJ2ViAND7nhT3S6p33eajK04XmDAtbT7OpMiDqGbex5D6aVBgDZAL9E25TRM/XUfs
8ZwR/BkLNgBH4wjjF1Yfbmy8VotHu5sgBCrwqrZ0qrlVL5FxY2GjbpcfazK7VmJbebP+gDvqyryY
oDYvUN/1RNb4/V4R++GDke5XS13e4RKfnZ1Q+Y1LQiDVacyJIUcGbP9kxgzOcul+eypk2kjfaAmj
ITX+Gn1QW77bATr1NFcKTMHvHyh3NlzmV/NNdSekYdUEaL2GAL0o3WbkVpUxzrJkCwZJZMJ5h+1y
YL18GT3UW87oP4mwpHjbHuFTBQuZQBrTHaZRIzZFQCiScbzxbmAbPMXDziuvoiUqv8+ZfGg4DKu6
PAyfnwNUkTKSTwN90+tM+ZQdSPMiuXvXkSpbJ42SD8cHdvUQZYzRuYSuTa/hKdRn+kY1PaaLaxGK
wfTeQ19v5frmQPWcwxaE/7WGsVLpexoi05IMFTDPkrVj2yXAXaSsa3au4jVclzFJEJJEb3x0dzxK
QyQM20UQr7E031+vtmg+YtYpLCo5rTajxtKegRV8JAtcPdc6Ak56W1GuUVwY/G4MRDqkE+V+2Uce
vNzRVvey7dAvMz2J/seEX38DRMR/N8BAbBdWpinNpPdFX240I4/a80Ve4yC/Ytw3IaJUCdZP2zoj
faeGP78Q0rYjmR896Sx8cKz51dQHK+SmRowixiGiNvbEc+cAwQbIn+U/BjoeB9GRnloubF7PVDqm
QzJ31GfgtaVzOQ4FKsMKi7g8vFeU3qDHc7nDg0V3q3EMtwJc75vbt4wP145fDy8pa1Djvd2GZbES
qY78kk0GlrxGw+hRWNofm7ceobx3hyOyLb2ojoItwQBKkvRYWrxQDTeu5O2sUM/zgkB7p5Lz/dt1
CEkBp8tg//AGEpEP0Ssy7IcMI0GsDhD+5xek/9MfqL8fUOIBo03GDi01NO+7EqtK4DZQ7oKGzmin
AYuqQfPQjfRCgq5k7CUpBXM++3/jJlkK43gLv3mC/nrMlb+107SGjYt3hSk1xl+k7f6QApq823AM
Bu/ter8tL9gYEKyay/aNecoaYMZhE/2MOsMVl7EVqPmANxfo0CNi6M7li2fSECxnOdUsug1PQqqy
EuXFS7SoFrZtnBDGqLmsBri4GgxgtGff+6QkkpMrS+O1Unb+jpdvx2KvxUSDcKQ37UF0UJ3Ke4FE
olvQqjPhZQshGjwddnOweStbxnhJxSkQrhkuCOxcqIjjVCEijbGBMkCrsS15GH3HmmVAPskMs/Qg
yUIqou1K+8QbNXpxHNogKTxX3GjxEnpPwRmIXoB8fJ3zARm22NtlEw1qFfn6QRCc1+80a2mZqlg0
/1BH5/mSFqIHBYFDZFWEPgOkYqi2sWeojj+OY1p9PUDYoszAdGWJ4PEZBqWXuWBD0EqxGgnr99oZ
J/8K+IlPOpVW9SGpzYKMdfBdld6iYo0KfBQePx+GxoHeoxASz1j818YL3h90GjDWa6dMktJD/Rnd
FhGNwmQ0RAU253pEuwZSxg09y0X6JuEzN+RxBInuPA5KdvI4xbOYJUor2WxICLM/+sJjhWcLWNge
rVBiuEKwGtAmrFZpl/hV9Dm2M+koYEUGntSaw2/jZrBf3rypQ4zYGoE1CAwGBTH8mGuAwNHrhIEg
eWYrSwAP5k9B3OGMFlZnn/oOZ2Bqti+aOgrBRoaz4rJJ8GB/gjqTqIqSs0xM9qXdOG6xoFikjvNf
2YyHWY6vHTnKZE7Hx9jjKwnYDyxiQhNOy9g50U5b/GViVIMySP2jTI6KIODQpBIKuQSKkBgiKmzm
2jQRnVowqsk6esI5zsBuIzKIkwquv3v4ObBqnBX7ibtZwiZarWknFRNhnFtsqWuHihETbJEdJ7C9
NE05d0WICloBbbkX2x+oicQdDrxGXa1BvgnrDmctojzhb9NOI8iJWGtfJ5KXVz1bs3PI1hk4t8tn
YovuLiGq2BR9HBUI/hRPTfQ8C1/RoEF0zg1p5jB7EiM0D23IByDLPhnIKp5sN0Jm1hC+vbcx2mmp
dcF+NfIEp2MpIRVfSmH0ImWE9HNj7btr/+VX+minTL1beHnlA2OfwQytWpqHQEBnaX7W1bmH+442
sn8nFZlLqcqOZEqTD18in7DRPqh36TqARTCsOcwhXPkJbvrqyU1VahCn7qkGKjFZ2oDRb6EYT3F1
gGfDoF2BeMdRTHi4DsJe07qj/9941Qx0jJyeRID7XLIyubCc2FDeUCYnNDwR5d1DSJl7+qhbZjc7
WgQdgOtD+JLjVBaiL5FCuIGqCtcpJ60uh1FgTlsJUnxXigIH+qONbEbOosOG+Sogl65mmhuvLCkY
BL8mstQRw0wy30bVYXcn6UN1y8aY2LnNM13KLX2oOuez1LG72pkA6InoxQS1A6DJDrgubXUpZSkK
0EmRZwADqcMazG6qJ5+E6Y1Mx1nyTU/4qktsD5U7Vxiahi2mfrgKgFpTjIXUx7YIPxUHFF4AUQr5
oQjiqN/qDTgM8Bdi7e5KBl/EDwfNyPaBrFSRrH6ASLhhL9JhX5BwyjD4aDEvHQDDTrM+LQJVMPJT
9CwD5bDDsJC3JrJMNK+hITbiz6/JIA+EZigvZYLxEmjNuiZ/IvGgjODtiygcqIXZDs3A9UPkpTMe
Bm//XnDIulmzb/6q21ZKD5xg37SluamAFOztOMM9yVd4GJ2Mwq7zyLQQ1pHu959rCUOG0OJclJCD
dsOgw5aQp76Wv1UJZMVCIwgv1Sm5Xj7dvTQT7liY3IlrLWdG9B5jOjolcgKEk4fxhJWvWhuT4oBp
uStTskDRiw0fa0QWz+bcRpEP35BYYjgB12bYrUdvEFPoYxGj6EIUqt4OljEgNwTqPOAmOuZI1rRi
P3AedyPeCLpxTajJjgWAmFdTzMhSsTbJbNLS8Em64b4zyxF0Bo6PIP83lg1bJu3vzZJfagkImWGd
w2mok/SEIgYbIIpw8YiuHBE3mH3LDHMh79mT9FeuWsI+ljwrP+uvijIbDfjneHfTR1tx4zWCBdcF
E1Q7uHNsT0tdCjwaBLn+OUEZ9rtqGRAhfR27T0vJiD+yN3zJ890Ird8+oG68saIziYDynhfZhZ2m
Utz/OWgPve0GlX1DrHIP/kUZIqimSb89Ebvf+3ZnCBaSoPdaFlN5HTK6qrYRZXpU6mkYNyw6Ax0n
yzuaT9Jnwz3KB2I/JOzSjDC0UracVIYHAdDuP5Zd3HFUCC4q6eV0oPH0NR8LQeLDAOTvtB2uH/Lg
9AlbbsJ5FESo0hAbmiXlcVvUWnNKjc7UmIxDZhKqWdyforUxHWj69SSvvcuBMzSEJ4UjYjuHXEmn
5kwQl58ZDfABF4EwKbE1r5uVpSBvBsvVoL2OAEo3zoLeqaG3k+VdXYen43llshDtghXwdTTPUaBQ
mdpTDA4zwBHhm3Q36qh1rE8oyjhsGPlh1MfR2Wi56riWdBZ+abUMgRjnTWayCRW5O5Dhx/wdbwQT
OYjIJrk6CygZqa1FMhlyPZDdOVZkpfKZyvelydFfuPT0aqSrQbxZb0vUDY5oLmxBsnhdbl3jPOnJ
espjkB3DYQzsYNHVWyc/uaNAdHHQ+Ki4/4/nTpbbE47iT4A8ROFE5tkosLofzJ5V4D4rM0j0ihfU
Lfvrl0UVgDrL5I0z/fi3c+P0Z3pfcFEx6kEIKpPU5hyUmQN1rh+9G+ieg9sQX0zCZmqJOu7Bzx95
WPrImydiJKynHaoIr9q7B56dUmfxpwEnNoKclwiMmxkO8d5UQtDyp9w1CgZj/J519bfT2WBdv/t8
QKKluNLFst0U02KO+1GVxiLIA1UufUWQqY1Jupw21Zh2EtA4/GFw8bXIxjEeJ4Zs2lIjCA8e92Tg
9WwyWvYRrpLa75DXDLJSVYgyk6/xplHbrYILiC/C5juflAEd+p+S3YXv6EWXTsr6oh9Zsnh6QAEp
32/mgpLk1NSNtWboZW4yACan/+T6kWJtP/wNwh79n/VETWm8KGNpgKujMSdRieqrgH8AvdNXmkQQ
rGiWsgPJERWdrJaLwJS+F+ZrZCZ5V7B7A031hC/UBP2xKSxJTAtmyDgtlAYLTFPQNpITxXU+2PkP
q04n0WJ6Ekum4HDOQWK8N1eWnOoDPuvzauOkQTL9q5oOsPfWZPDZ4w0v7XJL4fbCmlGj5mS5v7Yv
k7pfV4r+pPceID7oIDTuN1JfUaRyb/5yJeqzDJZ1n/IL5tDC7H2rwG999/ashoFWcWW8DP7nckXK
WLsr2Uds+S/YukBqtAXGjGny9mxXirIPYDrGzi+9NjZ9wH27hPTU/s1ZubPaUfST9t9Rr2TMcDnl
Ip3lD9NLztOe5P6ogzwbXT70J+x4Z5IWtG4+Iyc49ox3eF7hpUwYUNJie4WKXHiXbDhiVRr5NsJQ
VTucNUg2sTU15W2QbOW2DMVOdrUYXVokz/uOPqCEvsFUzBLXCw9Tx2cgsgT8EHJBhZaVCpfBlPZz
W5PoLCSs1VonMB2DX/WXGO9PQxyT3JmGuvZ2stSrcQRBl7Jkyrpyp0F7vc1h8Lz1pLWmCgu81mgT
y/YIb0FOj3jsexCIm2juC59gUWUVSihejtvWDgvAP9xdXmABvybzoWlqnPTJCD5fVM2HTU2wtrpK
mBg0/GVkFPEIMe0Ly/kdaQ9K+L7xvAC/VPTTzqb42TfnEJXbLO+k9RSI0tIH45SQMITCqtlTg1va
cs6pn0zqwOH+FsE4nB92iBe4YYb3FsMH9fzUIQtJUfwhSdiocBnAFDfsiTo3M1P2baODLoIEaLMh
VrJ5KzYusN0tqh5GGdz9xvhoJtYQ8NiI16aN+vzLLtRuZtFx1LB/u04vhjQuEIV8xlgjBVbRLxIQ
/Q45Ueri+XoayFfS2K8YGjDNpAcw5QmMknyjivLTUVu666LfhQGlRh9KG9ABezJx3Oldv6G9GoP/
UjbctAJYeLWZQXhy5tlDpkTNgJporJO1qvZGEYVAxz3PZNGWxTblp9PaKiKqTlJUMZQlBNfvj1f5
XcKtG2H+pjXWeLzI+9GEBLNbASvI3PCTgv+IL48ied2C5d1Rdw2kS47OD8AxdRmDqwYaZRluoOek
aVuNDgrCSFCk1AMUSzbF8YPRXk0AnsYN9am86hBgmEM5ogfhFwCqA2wFfCzHQYQsMiLseruBMrX3
uWjWofYwjmNoIAkqEj8apcN6ofZH2FI9jSrB4PInwuON+0QEX5K/XhB+mSy839nvQ93ZJAUvcVdu
o8L3oyxdveuw3saX8Do50deYRwKfYx6WX2ZZQtSQALN/Jofu+/0HgVdSuf9pDXsrbqAwdPOho1mD
Cdt59jtRa3Eu3eIQtaZ4X8J6lJQHV9WSASeEMry3YlIozP5akzg7vVcRF/J6fkmcNCjiUgEFXoMq
CLEv/SkWFy/Pfh3IJbkXFlPBbIqWoAvqJwNgmmcT+0rnBIvM7e1B5n88xJIoTcA4fr+YAdhwua54
VtUPbwcvNQ2cU0iwaICaH+9VkmXfDXSVyd+qFhIDSKVw12bEQPmMsb9Ik8dmpl9xP5vpdteTa3s7
1BLd25n0bGwvssZt0roWvFjsEODxLuReSMkj7LA2/ICXESPanlKShwihlmstWPHn8G8TAzkQIOmU
1GI7ggIKgjfqwKTzeZ/5r15WxQWgXwYWuXGIFfORPMzBgc6tnkytUCPk4K29iRbBe7wIl7tly3TK
OWPnhnifd4PrGZ/vTFRKuxvwEaiF/SCQu/vcZhIxRmFGgyMlhf9J2sMUyFxxxxIBQWCkxaM91uDP
sHgKzWyiUaqK+/2K1VuZgCZD9gn7Ii9CevI95ZfvunSMwudQ69gsnM8XYbi2lsOMKEJDA6X6S/gJ
5MQKXfQt3rQVmUO35juZnRPBUMk/Musq7ad/81RVhm2UYrhDPcgTok1hkCAt5O8uf7WeE5vAT7ND
08S7bf9PyP5MpW4khO0pPlA6sDNfYICGiUcNR/qSg+BIgjDh7Ya6B+1ViRNqOD9bKuJgNhsJYVeD
JiEszCD3+5yb+zX1q8cS5x6pomRskFLS+5tzVQWhxh2ArP9NuJ47zIW41ztiedxTqAPl2ZxRwKi1
iDiR7Z+2uEWzSIdnpeyHEC4/Pl/IJAO6q8++qjdLskjU2p86AyV/wCANF59L+eOtMN0/iFkYVWvL
UGHuI/k0e8S5Rgi0prNW96y2usg7LSumxonZe8Juk5XzBW7WIbUDCudxnI9J2a7S6czpS5RiRXL3
YE09/lU01dQFYmyxONVJqNcNFd1TpKt0r8nEUOIWCgHmy1YRX4pZa3heMU+NfnHtcDftrUFQAWzd
yxmJKQiy/2qzVDE6/N4Z5w6ux3Puiv9ZuA+sfsdHEZOE47E1LQmGhBFB9dt+chqqXm8FUoZJxCLc
0auPPh3vJWyfBlVPrFYRV7ZO0TLGCeJp8HNO5PGLIpf0en2Ao4lNkEORqusk5klHWYnktTc7yv42
YulYieu0NpTpQsrbaP8CQgoUOFH9JvblztO7kQ7wsce9Saop7Np9b8D0S0iL0pzbecLAFvsXIoLv
qFXYnO7TeUgMBMAFMFuhTMWrsL0XcdLj+E8jfF3UbP6I8hobnxtjp/ZCF14ElAnz4sLnmZ1/nVuk
DiH516iIBe0wawChSPgrUWz/Dh6qZImTD7PCVjfVVQdh6fHydOd7in6bNsG0rTvxP7+C8JxgRRIo
ROMZzN3Hqu159fjI9IVWtQcJxUwI+BY/Nj5h/702+at37UaDlkjDIMBPlDyznc8RjSWuezNAkabC
xc9z4rmnVeC1nzoUv4HQimROwjAqe0Xg+jH4rA6HTHFt9sYCHtBRXhHgRazuwaU8sYLhQZQOVFYw
Puby9rrqEptyqTkrou7hppgaXRzJZDVU63OyhSy+8BvelLjWpb/3LLxjakRthWHw2QFktZXFUAdv
SNJ7G5xFLZv/oR9Y07vWQrWwm4JJNvPNzCRHxUpS1SkPDkM7tDLs8b14KJ5boR8f5rrvSlhPU2AJ
MZevfmfU18t+6kQmO2Qhd9tCpeKReKO9sC9XULRMBMExQyfUZVxi7UrEWhKYPwqUZHKe5Q4h4xFw
taSk37ZZskbw3Au9lUIXhk6KLY1NMCac7ELZ34MWlzzX7Z5nt+ZtzNBtQKqKeUNwBt1EdimtgjHt
0rgiUsERt2KUj97S3rIu5e+GMKSzeAWRL4PEtlEbaEQoTEn7xVHsbczKP7Rsusd/GkRBat9bnVjg
G0ze4iWyLPzCaMq7MRLDnshVl9uy4tScs5Dt0JKqQaa4Wogqg3Dkq7oussrwTvFnHbgPSPh2twD0
9cHv+4tkrTTijAZ/mlckyya8WTkU8mntFKVU7PwSpzPWLPrru5TTTyORVm7iaBEzyB+u92B+4WgI
6yYex+I4VjEOJTCT5OOETUYRNXZiLfUU7yumbGS5KoOtll6NAxnhUtgjDyv3C5EHjf8tYc+kxU5v
8vkwgfKN8LMqLVFjZ+b0y5sLVNX/itq+4zNqeVLDGyVEInf5/Gej3DUkdmQXTPDmkK8UaxPM7LXk
HeGR2uMafNzqU4NCSSRDtNxSMZFXm7SpNMLTtxWl48X0IaXgfgaHaPtA/902dZj4BZktIsthAT1R
FpajM9jX+dmjrYCFM/mZ19PDB0cMaOuBRXqjHaT+fUQ371Ctk/f+35JFySGx/sDWvk49sqnJIdrd
HOQjMxJayq1Me1wU92qoXiRxuwefgvEXRVC4Nw23JW5qVqkDkVw/roYXJru8SuKmHXcndiIDummC
YuF2/CmGtc0Z6YUwJLAy5yK8dFXpNBM1RjPUHEY9MUPaylvnpq9pZxajv4gF8kC7Kj8ssvMv6n4B
9dsocrIM/RIrTBqo0mVKG8vynzT3tatPFNePbb3bGV0fW8U9eMRViJXlgw4Oet/rvOV7v4Dcx/ZH
LaRraH92S4qmHY9YKzSpdVNJ6oUw5KOjKBH5nAQyuO45Q9PCLhHiXP7Yn9kTarDVHIDZMaB1Um4v
VCMUkznmLYPBiQZ4/Htr1x7ZrldVtU2Mpqn++wzKtw12FdZTXYeVuEKBkc+lBvcaXfo9jvpitBJg
bUymgQ4uxStApjxaIvmy6zVw0avVxdNRKkKAXh+5oOKj6PJmVQWXiOOdJSmrzO31x5u5gvGXDGkD
FPE+1kRTMJKJdpdhalW6iGaqgJ84vU/85Zwq0d2/tN+OhJL+e2MKB4iK5RAMLnvfR65qbPl1nbot
YoiZIRDjzTTYIltBAPNAusHR0hfpKQi9tOkH8aVd+2xzoZJBlWWJlhGnXG0pMzp/KfkJs35SnEbj
wuPMnNtCw6VOA9Gk5n21y4/7oEfU8ZTCj7z5yLBbSUxOIu00FC5zw5cB0piqeeUYw3Qgnc+8/wcp
cFWALO3uPZgqZkPfCclq/t6cDxWV6baVYQT/pha3Kxm222dpjeibuoHocNDEUzAjD9SdLit9LOFt
B5YXFRvhAQy48ENdN6IJf0V9zqENJzlurE8mvv9nUNiH2vTWnQ5xVk0Em7R/Z29iQJOAPhzaB1N+
clqGzxe0qecOKeyZ/c+w99tC5a2u038hdVcQwRQ3cg+4YoNx+8D2WORXZ6yqoww/6vHR27E/ZI1A
MwfDyluv9+QSJucvn6RR0SLRw7NiEGVAf/wmy2g9tNcZnFcRUep5VsEcJklt410Mr4JVZqyqyMEE
SE4t2d7P2P+Tc4CZL7jHU8b30tRWo2qduBtSP4pQo9eEGt/Jy7re8zttiiLD1xZhuJpOypKcSh63
EOvxebendOMXmyTumhIisPemuthOHKR9SMjCUkjSkethWiP9M7dKWtOx3C0fSbf3xGoeTl3108HG
OhV7+kBbV5mDxvBAsKgGnKGIVs/GyDGuDbqFFzjLQIKcXv2F3haT7ykjmfhPVr1ZdEa8GSgTRC0z
9NIgBwToZ1pRsSKI6XjKTAfWgrX7AcOYDzr8VnWX29RNSZYfGPmsn2HSLVua0L2uUSejQxG40Wd8
VePQe2K00N9lkIbDbgbAYavgP5BuqO5b4Dt1C5RiDTWf9pk3g2qrjtG3AZiiWd9Hx6nLfWpTc5EW
NnhwZ6R5qoubZRDNtc5VAxpwDy90WPErbnK7Evejibfsgz33gAxLp8Ku/gFXmq5otAOud8oPqwv5
7lCchPpb0wW6hhe/devCUoo5fp98eOhZWpT0Zu73KOj8AfWLZVaO8En9UmHFxlzMMkoPD2zDkC45
7uI5Nl5uiUH8eWaSvystjvPiF2rb2MMlFfNntUTW9pcyXvx0lnJgCzA4Ki7esiVxmnaVDzU9XzdR
U+bkga1aVx8HOWPSCFCTbUpIvVUbn5lhwMMbLTG/fDjN/BN8N9bunboHCp9hvDMA3M5JI4hEr0l1
qtMrEyCMgD/LYSWI9ifxYl0xnJNRKZXMeHVSgEIcuuyZL6CMZw7YcdoUBhyNtda7ZwqDylHReDV4
10jbEgOC73usmrnaTsukWKDEeSzJg7UqeOAFKGbGP+dmM8lgSLjHm92rhq1c27wanVp7P2VSszCv
poKxU4uS1MYzmeT21BLTp3e9nWswqjHrG7GHCER/TKmz+ZPIarJcNm7QsVeDIaKNXOQVHqsdcBqE
+WGp3m60D5457I/fvsouMOA7z3unm6zhZWB02g5A1ns3//K5SEzCpTNG4cVJ6yRukIMGFsW9rUGH
cO3NBpGNuxmSnx6vpHR4B60PNJgS2PL+MK18hiHKGHWL+Ezvoe+5nLbdPp5ypdixyTX0eeOzTgnj
hO8lAhYbC5VcHXp0BvWsdo/F590KqnIx37iyW8OwYF4UF7FEGhJc0ECyM02CME9COPU7Z263kTCv
8pePivc1vUUe5ah+B1X+74c/1IFXr3yx/DGH/Qlr97Hx7SJXL+U+G8JPjkGY3d0+Qp9iCmV3O/Ol
E7aq3QHdCZAdWVymVyO4tr79onK9Y9NELhaF8yiVsBheBTawCshL2MjmPYvW37NHdSq2iWmSskuo
2880ttLKHJh5wE6+5zSkxpEWQSvEFztrlk9V7YtwUfjatJjENu7HNp9MZTDmJjTCa6xL3EZfYvOZ
PBES+UT3lzjrtn9HScObOyqh9QwAb6ePzmym2K4wA8JZ4XdOjQ/Oc082Q3xlseNkOEyTLC0rQBVC
Dp118GM6fPsBdE7+dL2U6LA0WE37/BCsqFd3NRMx5TIjUQ67F9IbYAbk3np0KoaAxRdZNhLSgNw1
VdH1CmSKRtC/UXSLQ6wqKSjSbX3AdhtwJR7oYp0KS7Q83cqXcUZ9ne8E9m5HjoTz+VO/QF6pKrCk
v2YDgOtCWJKcadQjGyDFIKxIUXDhu85hqq8ImKZymar/M97SWoPPfSsfI1XX1WKSwfURg38gqsvO
esEy3X3VGTuSRZ6/URgXmyQSvMMYTHT7pvEf/9F+AOpvxIo24LVGqtZRoY/pnOLaQWFDwgsD5z2e
40QmS1NVaTYEKEAUtVV6DEQz6MpDHrvhdkcrlB/mKfKz/V6Z58LqmkeXpB9d9WA+G9QrL+Sg6NW0
hbV/mQQeh05gPndYLCkx9mCYw8a1l455AKZz7LHnkm/kya1tTLLG3yiodWzSUQgpfdwIItro6/6e
l8DtOmNTgES4xw8GBPuahf2xzlartoANnuLr7/iq78uk0PpSTa1ZDgXEZ4xg+swPhqmBCxwOGGqx
TjnIYNxGQd8u2wrJqTskgYdpTJGhSJSWfcLNkFK0qPWNHSm1voop20epqS0YWOJQ0UMisAPnMDcj
wVPgw3Yf0GkRBAkexV3i8QXjUoOAAV52HfzPq68/DujHys4o1XLC+nJHk/iSjN2FUGzzKc6wmnLV
yXQFF/hm4is6yX8vZL2mOA2BUgijQqCgVTUTFYF96XP/08K7IyM6kWJa4J73Evwy+EiSeqsnRycV
2kLwWbDOzpctsn5FkftRX4mkB1/NEYXhwt1NN7j/GRDEabtx9FTlEoc/KKiuRzCA5vbFGFomi4j6
Z0igZxavFV6aiV4WcDRGKxptcQwNMREfFw7XfKxQM6VbzHPBolCsRQoZvUQr/KHyEPzl1+fgaUvR
erSZRT9PgtlJVfD6vkv8Gxx1DAPW9B3ihqe7f0fOmeVqNW0SBzUGQt/wCED0/upPfukzSaAK/wu5
/25VD6QvXjWT1ETn/MlYh/YuBZYeWYjxEPZYJucNDPPyKsin0cZypN577e0r2mB9oMOGShfchiQs
lw7YUQGfpRKDsat1+BLQ8EjDn4dB+GQpDFmx5Pq3Wjv1VUtxLhMdaIxtZPRwxtDJiyJl77EFp65b
oGkYS/6b40nFnfJ1yuY89DGuNYBU/a7N/o8mqOKsXDMzmu9xTkKly8r5ouyH6FehgpAc72UI1uvl
kXFLPJ+CDCJOxIVnc6i276HM/ity88fOEtbq7tu2fJYrw9gLJymOCZliEmiEFaPvXUTzwriIrIcx
lxQgk5z6NVgfSzjG49qxJKyFvRJyAO4O51wlI5PbKppYg4wEODa2nJJiaKSd4+tVYpdBIb0w2aMm
384erA39s+xe1jL/4mrXw7TgSnx4kBM9euW0C2hUf6T88aZ/TmiHoQURguJxkW5Of/O3FsXgjf9o
5xtKGDCK6HQVcW+z5uj0rkecPfFTpWpfBvzLxwVe0JKVAzXfybVyjl33LuifJPSR/YKZtEhC4/8H
7/UhsIpjtXOro/7nys9KSHyM7cefVSh7NMOiTgCV1GbRKs16QsboXXFSbqnfILYdHAbjYY1XjuMV
1EjT2rY4xd6aHA9VAKRd0jxQBRNUcfFCHzoFhoS6sf7TKDifzmM/+naMUx9XcHrYgeXxaJz6XnS7
SPwidJVfBZB5cpBJYBsPgDjbJgzJ8vLiS/wSbdFMa0rStdFsJ5jU0k8pmflqrKNAinS9IdLYpWiC
J4MW6ke4U+aOsufUq8FAYcmOOxXdCXhPVn4xxx8eV1qodWjC0aHtSY+CfN0e/N5idVLqALNKK0Xj
i9Dgg9lLkp6OkIgrO+doJsrexkYu4RhiRJY5imgS6gp+JoFrbmT6ccXV9ToP7jPiiBoI453ismbE
ONOfvgMUfrkYgm8+tuYM6aM1wQi1bxWyPZ0snBM/CU3QD8c/2z4GMLQHrwtT10AMoo8Tf2h7vZar
qdvYdoaOmdqPqEi5Ozi83fSvIOByChork0Vd96S6LQlrfCOYuAUAyBo12LMlbP31HU8mYod6RUK2
ziDcj5E9X6U5cKbjs6ns9Rm+xd6tjM964mBf/XAfE4rliWE+sug4sH+ASqttLVyIvpK2bdw3pvjY
9ln2VH3jMEqn0SHSQmqd5jzlDq8TfTM8leyCz461BUaApXcpf5b8jzWZnWa+FIg340+Tc55LFwuw
7mHXjtsBTI+JtDM6yOLXpceu11HiblI/m9dOdndt48DxHj9InQMMgdKXcj1i6CDpdyhAuASaJjlp
Tk2GXDNDQabwPENCyiGlrouV9e3avZnl+xTKO2x/SwferUto3gtA40smLK4SvmmzIEPU6oQxZuj/
eyIZuQ7HfSpqQy29N5MZIrXBd5XNaZq7HYpHVoKOKBEWZT7+M0w9HobkKvuYWPNGc/9DA5JVG1et
tSpWIVvtqIMvGsfkcuaI2kH5wMESptqjIWcbyLktxueQQG63k7RSINoKnpD2ZeALNiBMZfRTdlR+
19QBrafs1eYljMPZQuCB1w85BRwh38VRlXhOeYeWCshxVGKT7Ml2nn7Tihqcb3CmBCxnJf2ZJXjv
GZuD2HE5ENp7H25yrcdRqdU6xVq+CsUKAXLkaN/fnOwvkEgzJeChM1Gs9A11IC1vBHAAHqgAnntm
f28FateXchYuxrUVbbPNT/XPyMgtr87WWixavJFLapHd7qxf8+6VpjOTVoDNBij1DiJuf5lDBxx7
AqLcnWAsSVdhLqXegFTRP4ufJLNwoYXhemI0VXpTaGF1CW3uRGoJ9D1Emldr7KoLeGPFz8lr4PvB
YFPgRL3Omfct0czAhsjIi8x+5W3fglonytti+x1SJ51UDmgZpyLQcW5VTK6KAFvkC9qVnI5A6VH8
oAt/+0+h4i5tCbAjbOVNeU+QvdPNEVORzq/Z82hRU2FZS0dTHRHrDyo0ahNAaFhop7vpYbNB0fHb
I2pFPVZ8oDYFdAJJ8r7YJksTM0ZrUgMDMOUeZ1KKWD/NiSJ3Gd0VExslKdhmf+szLXEhnayApZVH
QDlExZaGwF+17GWHdQpyz3CdBuirvk4I76pSiG+PHk3J2awBhmI3gawmI4T70DGJiljPAje1P6C4
sLNpooxM1PErw0dSIQ0A4fEzmUVrG2d1jKIfn35BSor57egN1gKs9+dC6cOmcl/EKxlCpDDz7hjz
vV2Kt43wrgrak6t5KWGux74fVQg0oDOZou9O2+TlBzUPwo/AtsyvclhJrT0KmXjACW89Pbe0FGEA
4fXtk163WlotLkdJhdrhOeTd0S5KFAJhVOZkH7s5fQ2l9DA0YuqrHssWjaB7Eaj4t0SELhBMlIyZ
MDOeCu36AGnUjEMEEeZYQEPpSYMGmZCsVdKybBJJu/4Dl4bUyk3tyZAXS5OdrMbSmsUw3MoZIyXU
6kRM6NmdGi49r41W+CCtTgnmtD2HQhPGd+m3AZEvJcAx52IZW4fcB2ZzAfF/7Ol4hQ6Zi1rTLOFx
fibhU7+tu5kQyD6F5dAucCnpdOhVH7bH49Lsh+YuNNaLuNH2fOuciF8XoZmnnpWzGa1+mQ8vpRNm
DB4fJv2jq2x0jT2Z4/Cd9x3e9IRVrTJDof9FbHkLur36+/7ID6wlYzd8KXfM64KvrqGLPvrfY40U
1Ili8JWtavtfqXL1XYInUkZpajnujfkr6N2uyy9aDP/Vi6el5K2Yv6HwJId6EKI+7TKyPEQV1wk1
VQtoK03wUGtfzhC4yToEhZgFDQBeK6/4YXgnQ0IejMFEeE5DlnlLdovCt3IWst4O/lSoMzK5/hun
rYTI/UFMpAIjrN9LAInjbTyu0sarmTQs2qDscc8mY4ZesX1rmhro2K2l7K66EmAGZrkR8PS7AMEC
qeN6hbSpHXBurCoH9xILkkGKsPgINr6QHmgAu/driDZAw5vreeEAzYROzsSI+3iaEJga1+ODTuOM
Ue01AosGljsRAXHC5RgdJtiIu3EYsAjl78EfUfBgEXqVZ4KYiQ2Q0oeWpxTWXaoHmFxB4KW7nFVO
6gQwkMhkQVoqFtXtIDlXRJwJn/0LvCutEUs4D4dcUwLzSIRVejM6MaFtlBjRlip7Uais3nrlDxFq
1FVfTaCuYwrQ0gkBppR4Z2hmsRow6+kNmuYvFTQ95nVXaBvbQgupUZO6sz3Nhs40t4iF+AJPn/qf
l3PjlpTXo5KteWzGPftCW4gSCTajwgo0WwH+KS0oFWR1pFpKQf2wyzh02uML4zTz6Gx4yDHlDm8u
2KDDI2vaU9n1a5qPRRweyWGwH5b8wUyo21NUs5usLfapJUtvuwlutGxGV5SHwDPcKXlGL/MmcAJ7
23lQuZhCiSpsPTmkSo3J2NBNHaAl9GBLvyUXwPDSEXTsizW2vVgbf3esRTCHKi0EtydkH9Qm4kG1
F9qK9srsP1j88B0zzkHHzbbD9ZNvRjFd588mmWnYZUXUAsqkERDBnSJF289/y2HvJ6aHN3Jc360H
lQuFSj0FDLbyvaFNSPiwJi4N1Dl4FLTccEKLxF56bNO30HsgI1qxurBWJSsfUqTJWOmI/dZV6Ubm
U/5tWWJ3w6bDyoo+cK++Gh93CtvssGMNXRDlqI4Ey65tcLVtTWgIuld9+gHpYGlKEraBqSHhCbSI
5VBEKKYgPz3ZbB/As2h9RTBkGbpKDefNOOp7/O1UrwWEhpBeSXNF3Wh8N8aq6LXivDaBonVZZY4Q
GgSIe5xtonDPCLhVurn2Srh3+9ofkC9YPRsEsut6TVnsFSfbPmCqqYEjjYj8H15rFGnibq7esn4R
aW4i8S8tpIyTqqUq6sddz8lC44w0sGJX0gBq/L0Oj0Fewcq4ZWq0B4xCh6fmEjkNAqcPPTZr/82w
d0cjjd5Mj+gxxfI1isM3gjAzlQL8B6lkYTJt/Dd5kIVfht/lXZCDeUI/FEOMtiP5kElsDPPwjcKo
SOlhyTErL9wCCbKwg1Ap0Lmbu4C+L7KKRG7DEa0gr+zFUMrFmoV9JUw6ewEAWka4DqCpr6GxMwe8
UbfVr3mG8qOojHQetuvoGrVDM+NTgyugU53K+uHSEOvu4gahGjkUud0p7AHfbrHrBhkTb2g5wX9a
sZjOglqsNvCe/rcTNysj5CUCqmwU/sXMieO97PWlsxkbr1J79elO9eaRna6LEKK47ujfpGatu4yd
rqAn9iiuNyhsIpzLVw/TsX8KgNXR3uRmd9vLWPso7rvgv0p+d3j64VHxfdybyK+CJqNkcxM1oY+4
7yFt6Z8UYCJbDa/zvCIG+msQu7JNuODaqmlXSmSoRnE2BJzEdXk0+oyvUuAaBoyZy3PX5S0KWn/Y
3qd8vwjEI2ccdQWowC4p/5woAjK7OKU9Mn7e1aEjQptd6YovJy4mffuK5YlS6scbeMG3GEyu9zRb
c92wYTxu97tW+1215GP0Ww770RyMjfQFO03fcbdiCPQr8D3cQYm2uLkdBteOZACUajYhUEcO072S
8HwRnBG0N4O58d8hdDkEDuUu3S42tMi4jOVnoeu7z3cCV/t27ACZI0zo8rK8cZiXztJCp7xQ9Qvb
BPtbzcJEoftL10s9DMP6M2M0Nx3wj1qBUsyMQQdp5H4c0aabZn+7JbD2kMePctD7mP2eOv6XKda+
0G4kGSTIGYYeVWtKzvE3v6o1fICdV+2eZF0pjMPgEdligkoAFEj4V115L8rNHiGbBi29OoJLXuj8
DQpO4VlaeJY0xkT2b8tWZnKMhTtGc0cU7tLkqLnXW28KlYYcO/WEe0/FuE3LocUXGFeFaMUpj755
x5v5M6w9r0iLlHhp7czoBt2kJaN467jBKJaaZOUyd/fc99BGi6rKicuOgnKUjQp5/JkkzTsza0Wu
9SG5TkvVQwMuSYDhjJjgqytAAFRscXGV+kitOCxSqwhJQD1F6MsbPO4VACJPLX4y9TsB1Jsdioq0
zLKKFOmTD+qfoiIpCz/MuhOyVvPgr86joi57elhMCyiYKD0IMUYtqnEKWnqYNet9aHbfRYGZenjs
SsLWR7FJgYgRyLvHv6vUVkn0Rk+iuX1yPwsNXQLAlaPpyt4MeH5Jw6pxnNAEDGBp1IdgpzG3EUUN
0CGqXLX4juhHd8ZQgdZ0PykzWEHvWJ7EUvoH9vxSdo0LtwRDZGOF3HMX3snN4IOBePvegsooEiHO
5ctvrOMGGHJWpBmvtrpAJvDpLCNRsk4+cJGjJmLVTgruYp6N49vjUwFrVuAq0f9ZltQfga6UFQo0
w5WVTzEQD40AweshOqkeqsLADju7ihTdnjkeQomRxQGGVzhz/l6jiMTBmvFII2333ajDs+4wI76/
pw1NJlPux0DQn/4GxASi+gdM35Pscu8JrgNDZMc+dZq8RZOCC+9wQlIOyC5VJS/vyeNJvE6tPWiV
IWzLmZBbLCtnO05Xvoff17xVxYyOkr3Q2AThsB4L/DL+N3ZBxP4ToPCdS1RShKg1X1ydL01A3Ufr
yki5f1I3r2YtTmSQ/Zgp1kFUFAk/LoKlNFSVb1MQrMe+9VjP/SUHS/dHE7Zwpz3Q/mhAoInWhQbx
jCr+GG2ZNt0NHL6Md+/brF2k7Ujbi34tKeaSgHrmNWoWcgt6EXPb0eL14yU4dZT1ucbng44kFXc0
ygAPEpxnMrkNbj75qITnwRaIvsUGSa7bBLfzBwaWvCFCe7XiqjSr6hqMw1NuwpxbfeCbMSJvtkhv
QhZNVds/K7ab1AkbiCZgmvLB+VJjwXlYyjkEWDoKpIT4H6J6eyDM7BG4fLLjPBZtvWprXjVvYbK8
UhR9x1q96t3oGQ6hC7Yyn8pmcDHaD3I5wRTMgoi1rws4HpCw+SRbXnMsvbF1LNDEb+7LL3J1ViiV
nOv1dlLYmBExoUyvRm/F9lycrah6/OPKogibfjUVjqQ+lFsibYPJVFgOn0WO8Kc3EfM5y+Ai4oyp
cA+kn/mv3RgpLQL1Qus7aGHoxDGJz68oOOkgdWWSwvR3CcG/GAPGs6lTckNNnblvsI9sBc1RyxCS
c9qTLFfsk5HnMDWulwLfQNVGOD1Dozd63w5aT+GSYFqy9Wx1+ypiQTfMHuRBrxjhGMXz/kyC91pX
MQnSNC1OhnMQcTmeCNuBJaJOIn89aCkITAzHUc45HTw7wY2ylrkGbiJObkh3AE24hewvaS7yRAie
M40hmGk45La5+wdHa5jkagsJlCYJaBCF5ak6VESsWLxG96oNOlgU9axHW3aFficeM+cpf2qXYYVa
raCJDeRHI5ZQHHiPANlTNjN6Q2IKejdKWaFdywn4Bhy1DVPTTY/hx/vfGVvJKZU8+OSGTORQp4Da
jfEwc3y6ZlXFuo35tQn8dBRL4R17tIor2mb3mb3p7Axp1aBmKgopMnnTuK0NZTRxx99VFjLvtyAc
0X38zVWM+jApYPPn6IO5aKUCAxZJXUw9CtNHGd1EB9m8hL4AgTepgviSCkgEyU/bnbuXcQOqrVD4
QxxfaktLs/w6bKRW0SRLPHcCfB7iXseIShvVSnz3GuR/Tg9KdOsS00PSODpNmNUdsCChX7OkkETq
sWD9tm0GZmPI2eD56+ZvMOJlPxETCAqNUNOmmBa9Hrc8VWpY5Okpebr8LSqCGnlZwbgav1S3B1g+
qI/wq7BMY3EkjvLUQNPKl834kJk5txdkbx10cIXWTg7Pv8+5hbf/83qvpoYv4sWfe0jqIkA/2iSx
yiUaQ6TcTmsMIMzfn5jDMpB/gPnXg/REal+jzkGQKcQvO6nTE+LljIjF0Rhs8eZk5yaVJWXD8GVf
U+AAc5OSn7dShg2kfl7lbuD+05Ufkp78lmHQXcZf1tpCl9CH1ayeI0t2jnvMlhAefruXnGyPgBgs
rEQkbsyzUcQ5Oi41aA0PoEqPDucT8q0wBiXpHBfnIHm8FPrvuOsWyn0cw8PU13b1SJpXP50jkMEf
hy3KcLNNGplSLGy4WPRdnZ9d2taX/3IHMzpVapyl9GSGWUCXN5hK797JwHeRsBVELbehYV8rAoum
jATq7S2W6bfUgqSafVVLB+g3oOS3Yiy9s4M8r6JWiOVmIyh0hRiRfQ1Chjkiooan55vlzr3UGj6U
OUET50uABiP0y/OrOA7xh+5z3pSp3w/6qlCqmMydbPPm0u21ZxR1KjlKGRaa0T3TCM3FrF1l17Rk
WA+us2ANIoXfaA3KobJHeTwj1hTJcm0arUPwXLHAK0dA+PbWVBe1k3lEFX6rGun/N/7uEHd4u2o8
HfXkNcGakGw6CjTHBJwhY2L8NkVY/Pl8ku+o0EKGJvbJQ425ri5H3LVqcDwgXOZDpo3ELXCKI828
FKT23X9K5/UYY4BW3zjVOmxABOJHY6ML+h2wTzWwC/Gs4mGDNvMAGtbVPUsRMkURCYCHCaaOXZpz
trTM5KdupqKcJQQ6tKxBytoo0D/7zFoVUecnINVQ9igjO2PdkOrTE3rLpvoFXueVFBOtn3SdXVPt
/mecWLY9jMjR2wq2ngR1bWuux44dfgmadZ49t9QClnfac0H8LU9LaTf2Z/YRAesnoLBcbEqcRPpO
zlpXVEuXg/SMbskbtbprJBCwnyHHfl9XSsiWIXFU6l6BXsmFjc0elPX0tWv4T/fez52QvQH0WI42
G04lGqtYx/xjquyMZJ8GUVMgNsV6jA+c0t6uNWBnnIheRpOGsx6erQAFNB954rpvf18loAyJz34J
sJy44zi0FY4hwRPjI/bZantWhKjlHgAOheDRTUzT/CnIRVy7kc4wl+34JoGCWCI0wgJtZISJ9v1K
XzekHj27zmHW8SdQabXp9bGNxAnP1t/T6ritUCSX9VgrOdt7YrYIS2u8Hs571U/xKosf4V+WXoo9
3il0s/60/8Rl0OwHVKIZ7DnNYOnaYtqb1GqJlIi4zh8AMdqDaQFqpA6pL1dCBceB/3BT46jOeimt
KHoPkwKAZcg4I9CFJsXrZJMLgY2SfrZK8IJ0Y1i7drHasXNRdrFNbRyFGrwlnkpRbAlUFntYp9iq
LZNHXjZ8lK5sEHnHo37CpiUQ9tEqlnYv2kzu8oSy6/N90WGGduXgTxs9lOPNriQrFKaYZSD/OenB
uyYcywBhi7G11dNprkroqG6XFVNQjZ1Um76N3WuhWCY2thW4jjxj4WCnniP2hBTlIjVolQ3R2LM0
xczj/1J5dREVFfNMpbnQXRTT2VS8xBD7miR+c+iIpdalDvlEvCIqeLGIdSwN4QyukdyEyCDR0VbM
TkHTFX21ltoWCeAWxYQVF/cQLpPZcJbVAtcqn34LcZMW0jD/C9eGxUDECwrkk+sZKuAlDMxWrLzj
SQcV4kpzdNx0nrclByeeTt8Xm613Qh+FJqg37knE2aIg792X5baSwlr0q3D8m1dBIx6de6o4CGx4
9h+vCdg0Rp39xeHWrZ2N3zawOnGxXEsPdQ6aG+cWVcVqdrSnrMwMNAvw4TOxJDQTFbGLswqgss70
7AaWgckPlAcc8ykGtHApVCU5XALmDFYXmknVRZiRvl7CLAzvVQUOOiUiPNZY+Gz2xzgfJ5efw0O0
8/hWqd9+iGHJj0dZkWf9H7cugLu5jBtfsNWgeM5kmzB/gLy9pJO7DKTAKsL70x0Tn8N7QGt66gSk
8gQEe7Bs5RZd4dafY0gjkAM+RSf4Rl7aeJ5FIwawN9/sc9g8Sws1bY7qmRXx5OmlnSCihIxzZuu4
213LGICiOAmqCX8EK1mEqxm9XcgCbm/4lGZ8YyneCYvyWSkLeaz9O+U6o+YpMNInCv7wrcSDon4P
I/F/i/j/j88hwBJ7GPZNZlJ7BEmCAQ5tReqHC2F+A8yEmJkzLBmQrnrSIY36KWCqvs8lHpes0NUJ
m+lruCTZOfxoAupXMb0taz6Mvkv420Lt0OjBMbp5ArYVy438XcOTJZQmN1E+S2whZO2y53CC1yb7
qr/HPrd7ONmperMMh27QETUAjQSpekaFJNWs2UFY7fiqhU8tM1R8A0yW3NsG3qBq32zZ8U3iC6rq
zV8scu67T2fadgRtCk1R8/RM3WcTLGryaF7clCs/LvyS2amIg1ayX9/qBqxKtsp03QglCV3P480k
Os0tFhkGMna66Pcmk7CDxV8nydPs8EfGyjBLN2/fsjnNmICbNrFf8yspQigQV/gG2zlW0NjnaQUu
oyPkC4374krfYhZvk2jP1iLkzAf4Fs6mG+gVNOgWLdxhFpoYBUfQfP1cIirjKCi1ehiGiqUVe9qT
P3h+z+Tzwfs8aSPjBuOhcs0/aP09cI73kt5BOhOIrgtnNgD1O1AIIWBZpDfFIyAULDvj27K1sUZ1
LYAEfvQEcSho7wpu9X2NIhFyVlrV4T0qg3p24/KOA4eVgOXORaeVBoB0pxBi3A6qXVqDVhuuTgNF
bKZJ15VVNEHMWtnhf/OsqNKA8ilyOjjV8VuiDpoDcdS1mdPyuhijK/IeA772m3moncuJRu78P5jJ
S+FBAa3IdBzoha9tLOrXum0pjOKbAtfDOlCW80eoUc2/FGycK5Qt/BNbgJPhhFWJd/VFn3d2HSHI
gZGPeT4MrVQSl18RpMllUdg6JMxXGzOcc/+VpIB4zc8zR71383BrIjMM0nngNXXHYwYbLNDcW8xB
hXKOn+yBT6+MkeGZWkEt8g6n3G05Swk6ncbiALCrXHGq6/rMZ7UUuEEvJL+j/LnVmDj6l9mC/7mP
3aW/2RQjJY2gLD+U/gqSEEj2Up9w8we1m8SxCmQvs1jIenjRfMsGQEj1aHxmfXjw6wJYCqOVR82q
fJGC+Rt4KYWTE7kggW3Pbmlk2/YMQVg/OiggR11Vq+BfBFC0b/kPE8IfeiwQH+PW5Cjnziji2faD
vHVFX9zvQsnZsgc7ofUxpPzhJRbaw8+ko3HM7NBJdAV67bu0xQN27iOvJzrdTLkrmYjZziPmMiYY
Ltn79EUJ6oBFU1o45znFAJQVnOZ9J/ZIxKAu1eGDjasSmJxSro5qOikiPc3XnjInGKGC0Uti2EoV
ZQe4RBqIjf2z2LyG/ai2XFiTAV5+FAEfoZCJ0sSIDDkS9ETxCpIHC12YVWCDyusZPQX9NOT9+ZHM
gcHSBcfLojlxy7nhimmvCHI9bYVnN5jP/arflsFpuwF1t0eksh2mhdodbkmLWa9dXxq2wii/zN1H
rs4nFykic+P816P0o5UpnVWFjPhadshP2g7UeXgLcw12LiGqbOHwomDa7OayNP1PjQNcXA2v+31l
mrK4I3rb98dP3n4l+VWr/7rjiqLLClNIzlRXPh/BCKlBONlU8KG9pbnzEE1pV0zT0esvuYgDEPS2
M53EWOR2tbx3msY6Z6meMJK1FjKlwbWE75GPmwCy6sPZ0x/hOI6Rkg+muHoE4T/41HLhVrh2O1YG
+JGwYiXzHzNUtkJgqIrOe/Mu4qYAYHtGwtlVm2uWWRVvDVpz7NGEZFn4HPqf1+wnJ/8zPGDlI0WU
YWbWjRxTR8US3NCm/ZMJwmYJL6GMm89X6Igd+4Uf91pqmmXkWj90S17vf+8m+wThUoTKIvL9c5sr
TZVcWlsZA2lqKZHXPN7RefB+xvWcWAgYvZdjTPEDSvx01tTAOLZs/SG+f5ZnFCeudxN7aI8BLk7G
wLftK5X3FHG0WuwPcJoxndH1vIsYTIDxiS24mvH/QFtdfi/YBuZBsVrO+TSQhOz86sKM7CkZw5cj
nNde/RMOJgWtPrJ6kxZH6AWDQR59iGCEAYfnLNgaGKvLsYpkj4VmO4yeSPDOUvM2EjLUCs7QC5O8
NYNcYulUW5ObXkERiWaOKGwVLZK7aY5x021QoFEX3QP2xOwOG+nizNtCKyy7OfHSt5x6fXWYV/D3
3hOUpz2p5ub0OfhD5x9mJfBAHg4esRkuYrt9vJzZFbmTW19or7oXpboyhO2I5DWz2xTdhZE3j5bm
Mu6iuUMltKnDhZT1NfVMH9v5QCUfUl8bumjN3Zb/GbRIF9dZwyvXJwomv+DyWANfQSRgIVNJAkTX
qoOoHoIcpAJYqnDqQGBTRioP5C0wG2zWvvkRP+CYtIbgcJ2w8WO1N+CzzoKucizlZ4ZLEMbXCXVG
r6OBIwhVu9EjL9OkImO77Ep2Llxtp9Aa9gBpfrVZNnuRYH2Jl3F9MHgBi/1qjGcWO0wklRUMd8Eg
O3V40Ma/K7uHKgzf69HLWg1NSMl/TqUoeNILjW52NHhWaXfIC6vsBD9OTyqokO9SsfSQCSrdmPe8
X95YHZl18t19rhgTqvJ4AkgJ7NgsqyL860YGVIVWPVLeTHO/LncDf0HfTHEo6NL7OzQrjsGOWUaH
NPd4qb49G4JLS/Idv5XB9ag9iAT4KDpcgsLbr3C9Qdkd518Ojkz2Qh1cKgSusQiqxlBuktoZLyXT
YnNKFNy/PywzM7H3jf8Mh2m7K5+qS+BtEjtr+Pj/akLbSm46yR2pe3IYrWrjSotCH/jilh8X9QRK
AySOXQitgbUuqgXob8wVKOyuhpIQeFLQyXz/rMxwYDAeP2hxkpXfiZGAAssmd/1CAkfuZNeu1WkS
8Yv1vCfmschxbYDQsRFIXriPKvG7Q68UD8iuTHUAtpZ/8PiZOtWbCMArpOOqRsMWuw1Yl+TucI2y
GQgxtjhcOlgk91Y2oG5zSNtXPHB5Kp8bK4tt585BGFymCd3u3ToYnxn2X1nAHHiOfHbElGoPhmqO
BDDp8/i1Qh/xo1xWXlLh37sc4nw7JCYL5RNi1nQAg5FEz/VxC1KtxJdhejW3F8fDbLZJnwRZpJ9b
7CBw7uakVyepTbFyVTVkbbRyMnK3ewzRIoT7nqBffsZguKgxW/MKhAvPljaWEjzytOEXZWhkh7T1
0deZ1sGkxq++94gLZJzUnAljIm4lAL6ju+5RxddAovgECZ1T8SuzVvqoe594AuhCPDv3Ydr/nwmA
m57gxgTqzcG/arTpxDUHc5FnKFs/coYXmepyQnu8Ya+sM8FpPw3TMXHARkv49kMpmXy4XbAe6Y48
DxVX8NFB5qUBpB17M+AFzgn0CdwDMClgRGolbgb3vc1TGE6/oeL8Ybc7g3lppFWaslrd8s7cZQx0
LDWkNmTjxmUsHdtjauEwmdElaLaFy8MpsKtI3yJqvRyVKSLt68xt/2IHG23846/rnMovM0xRnYXT
VAOyZbT4jwskKIMmKlVRFtlq1gp+TDqYC+aStD5GXrivLJQT1eZodEPqGQSt3uB8kjCqucxz8OOS
uXJavplabLmvs+/4TVlmRwcihl6wCC4LoSj33tS1hHew3cjs5s1mGPiESgNal1eeNt15Cl60Ygz/
ycL17y+Y8xRQ536OeRVWqZQKrkXt78DbGODxVtDepAglA3MnBycxuzT5okO6QZYNeeKwu+vSRedu
MtmajjbLp2TYrilmqXmAfDuIQE6BNF5d8NuDkmy/ValQIDFNllBZzSDKMKMquPXwtHFNMP+PKgel
fBj4w59hCCDRghBZFpomdyI/wjVA4ocj0XPIfLKbPmsjTlbVnlRODmsgl8MASsaJDOwf+0VHpnks
5cqf+C8Xmo8jG1/04eewaGxh/4HYULQykufJYzX5w3yzWGixvRlZ0KNgurSResgMGYNEfrUCoEbt
9yoqeR2UZe1jOcHipOcPk+BoFWfHyd/Bx/XDj7VzZ5SCq9sS4rfurEreTIKKWXimx7B8+ezmNbQQ
mobpW7zwSFY8YCzna5J4RpgsR4f3ideyIap2Piz93+vuoPMLgffBRRjkNCcuYJXI0YW5SBfgLlUo
DH3QJH46/tzALQIfXY5clpFuy/RMYsBiPQzGXq1kz6xYAVOLRSDTH1vuO30U2+gTV5BI67dwy8+e
8hZdKGQv8Kbg5r/y8MoRFQh2GWnI+E6sjLXysHoVBA4Q49jvcAMbVARcOWo7V2txjxllJsanPDeH
SB1CLRx9xi6GgFMmbcarC9bT44PRhEVhczb5n47+Qm1v1sV7/R9YnDei8UtKlC6RQvlQ3HhFhdY+
9sRk0IR+F88ZAaYJJHueAjypQiJEfnUX//lnDG3LeamhWCgbKkzc8BeZwX302OLPnjc7laP0n/hb
3APW0c9rswLr97+0RXnZtmXGXm5ERG7VGCfhEsaIzx53aFcKpnxeKqCTRmH83tZrxy++o097igKn
B0ekk/BsBV+cIZOg1OuZTgXt91XE5/KZveTBH8ByHkoTg5K6BJJTFykdxiMuQ6VZeCPYVhp9uC1u
h4b3fiQSiQaR2csZ0faWcepfxm1qeKdP3iWvMrM6bN1223BK0Xw+mwM3wMLe3cqSuoDGSOxbaW/B
YcSLAJ7u5WJiGZirtXSrferFDbd0WNhdYRHgZKjclxzyUhRSns6wKIHjkUBOsGkTryxHUpneY5I4
bvEtU6EaeGLYZIsHlAM8J034ltXcEbmTeCdITX5KIWI/SPEUWkwMgoJ4w0rSRP2eYf5dM1YxnZqe
c3gpDu+aRVsHMFZEmp8A/SbPFjSlvY7IrVuubAavYcY+Un/lViObQx9B1aizCYREmu2y93UVW4CX
lkFp9nttjh+zxnmFKQKfxwFkBosm4cNo6/vHKM8/CoDxZ+wpDyz9Bfx74806B3LyHeGg6MFgZWLb
G3Tuq5KB9a3kNRaBfHRv8WPEeWrnGe/ot3MMct+tBpRQxEv7QGdRBv/9/F7QS9vFmJ8Ea7E59/QH
Dn6kehIpr+Cey+9AERZEzXvzb/72E7v3Nvp3qQV9Bepj8mof9wFNtqCQKasgQkQMSTmAkCrtMkcp
6UeEAlRlxgUWDZrhPxX9uZUxBCJ5iMw4+BEYsZqQkIgnQ3VitNI0vKvuvX9DJcPXSQAIKYhknxq4
7Bs3cX5JdhTrvPoEg76pKgaY2h61tG7jArBlKmDbGb3x5y9b2a76+DUF2PvwH/xmupU8qjMQ7onW
6OfEdxp3v4FuBzBgNyEmqk+JMzdeVwySB3cpXWLIfz2N5ScxXUS3iJ08U0+E8jD0is3p5yZQdB0e
+P0ng9uuwJC74quM56M99P4chesb2aMuZNQzrmeVBhQw+JUhIeYuWmOwRimAVIOvSlvkbBzkLTbH
V7qSSbeyfD528JgRGhpo+hJPc+NEkiI1jBf1lgKAH/ZAhSZRPd8tC49v09gXEi4qMLy5St7dmfmY
5bmhoGzADYVt9if9mF5b6PcEf0NNk4yPLSHhqy1/xI2iQu/axhEkju1xO65PxeWioWjcKHQKrss1
oJvk1oqO4+de9MpKQprrfVPtDhhW7UXRbiiQiW043+t68mHVKIU8aXVVsN00GUgoZQ1gfD65pJkd
4kMFYk7ufspQ7j74hVYvkj+TEfp2zQ7NcKA0Mi63n91KCuO163XNpHm2chODplx/ITPMmFQFIAHb
xkaTdXclhAfe9JiMKlpnmcBRvmtWKWOiU/IvmegOO5rX8Z7NMRurNTmLl71vCWe31NpocG4j9wPN
IG9CIpkGd+HeySNIc2QnB1n6URPFIB0s0fsNUpJnT/Huz7dGZ3lYI6IlynDa0RzShL1qBzkiDxLy
mwZQwrEs04DPPJhJ1YiU5qti3KW2Su7S6yZ0l5NT7UFZtfms7kc2k7sbNgxG54/eJosnLYyHwwei
xnIpWU49ODCDa9iPzUljGsb7ePL4bjbrfj2T/JGIIcrwR5UdgEkto7V3MtnZXsbEU6BjrS3NXO32
9mvr+iwdWkufNb3tS9KtX1gdcN3h1AU/OGAAlGhjUrhhylIjoIfFr1Uc7fGcT/v6wEN742SVRmv1
N2FyEymcDfjZlZLTYeUtQXAO/uQad+L4YDZVIT35iOBMmCaPjUf8uQY5MxgjkTcbe6KIuQe1uO2Z
V3mFrIXiwngJIwyvktWUh2/QjGhVpaRxrLkMQDG/Gnc/dtdhmTGqVIfQyXyIdVYPcKmduvIvrGad
eAKJ1G6EZt2qEtWhvCIQb8Vrf3Lzuy26qp/hVkEWduUi8mejePu6rhDwH8LOQls6DRN3YfJI0WbP
iyzdDgpgomQxaW5MF2+RKKBM+ekFJy08oOVlzxxiOQywasnby66Nrs6CB2vC+SjZD1vgyo2U4Cpu
R+7RKh+xkIaqThxinuvoxlB/DMrdQI9/5XoC+Zh2SDyt0NNxJY3lKnx78Bd9AZLMPsu9FH4YJk4p
dSQYR29Thpv22c+Wcteh8BT/uOnACpVsT7TVD9vil6OtRAjzkAXhRqqX9vHROaaCDcM8O577FUNu
ZBTASCiLLj8JNewQTecJWYXKNpxMjdLE5bQhwWTVj/sC31virpvKDJYJXd4aJR0DvWWIqCfjMCbm
tz+l6sdHDmimAutKXfsfMJGvX44abKHJP/3gI1qPTFlPoCfYUQhYk2ERqo8tLleQga7m98KxpYvp
AoIN/jefMOAi3C8M/JiLsPjZkGAhgMi//N0h50/3wtW+3hljntNytUgmjg5kv+CRzv+acpCth9zR
Hm93oNv3qJMeb3RnftE+qpLNRBHw/7NaE9YAxeSGwBOXSA5kgJtLz25JqkEnWthgaPAHo7tS+1xQ
UwSeDq0zU3x9DDpyGBT/9T1xXQLTSf5xFoTKdCQwDqfPmTF/l7+bQlrhdUauDo4KAUFppiaw91sa
f6Qn8+Q7wpzOcvcsbibZ5c4jVUiQ2PEmtnBQLBuXIkgayeNHfwpwbuxMUYHWd37bVsVvdvlxctkc
UGCOGEQ0ilRCY4NcMS+khCX6lC3S4mj8oufwT8nswNRAU2dAh2DAe2/91ZOjjdugzX+D+eHlsvFE
gD4Z4O4WrvrhGSPlcjpYLGFh/ij2nyM4jfw4eXlZZdA0Q1wWBUn3i6cCcOICEGrP++z6EXev46te
sLH2JPKWz6PdIHHbe6f3evLwwd/qlgzKHbLPGZC115NNuFT5F8MZwwLub6GrkJfCY7zG+pwvXo63
niAhYNjpeBUHkyGj0N2mK2jPR7HnyrgcOVL2mR2eXU2RDedKbGORH4THPOx2CWMByS/o3gBrJjBx
mzp3tgOkEfPUw/4Fl5B6yyDM4AGB8Ibrvn0Hji2aoYKe5a+9lSR1CSCZ8X0tUC6uGfQ1g2WYe2y+
Dze5x17GPp0vZzjUyrx+a/mj7YBPU/rz66FA/mHf7OgfDxlPDfHUycnUaN85bDj/Ar3gX3HMhIOd
2aW3YUHvTQk8wDFAFFAm6Tg2CZmnmYMem3lTUAyeqicWawAyz/a5gGWKj/OrEZX4SYaJOWHCq897
TqYQWsxxX5eeOOPNk2Azi8q4jCRgnmsZIIq88UmTlTkWyRWYAPl7znez+k2Cf1x/ZeetTdfpgpP7
P/hSy7qYI8JvAPk/M2W87I6Z2Vc1TN6jPSkF3pbn12tKVM2qfFZ5ccXd+kHz01O83ZmzlJZn0B2x
FDpujJIZ0VOS3sgY8ScUeXEhs/T+y73tF7h8GogYqlf7Y4xAM1b/F4lbxbXEVnd9BRqrojivXYL9
W2nDyzDtIRHnllqyJ1B2iVDIASQOtN7DbM1XpOdjOxOFq5ifPJEn/mahXtH+sexBrnVvEsuKCWOu
hbU0AJBrs0eSUDNEIQDPtCpgcEoQhlIWk4tV4cqdlaO7Dg0t0CBXufrDxtoKngNg3SgrO8zwuwj4
5EEC2ScbfduF8zNEm5r46kSisKJR9RayBLasNLAZSclMarp8mcGqllKjAuhtibFXgmV99/x8aOnK
Xw2pN7/OmE0Dzubr+0W8Z3jdUXAzl42mYArRwuzzyNZ+OaamawNvMES1W4otj4tfaqJHXfWnzJjj
ejAEgHUzpGLsS4XkiQzW4tqp6HU3FgVbj1BNVCt0eHEuXpKQaTaeUZElUF2aXCt5/O5lr+s6Bk9k
7ENpiMD30Glr8gZMGi+GAmCU64eui586shwtyKv2kwRQz3nMquWncTzBsFq71RClYy0y4OiGTNDR
suEYdskT1HGjK2y2YIRDIHT9hCe08MmzxKa2sv2SbE0/kF6IwrWiHBmnBAeemNaLHM8tvG52mLGD
w5n4KAkW00ExSIxavlioP0SbM+tamIQF8bVcrkC8Sxjie9pg+6W2XEs4G9bqLfcqGwUarKmFydex
qazotGOZ+ZewZOk/Kk2Fbf0hBXFwj7faFCvyfMHK3g4qh92b6/sFAmL0ZiIjiGO+7PgQqKg8qwiM
Xr4NhJY+BfWrBsmoQt91s13m3DiWrSZkxUHCf116d/4VrK9269sNuKYIu56DtwHEQdZQi6dkqGuC
m2DRWsVqYTO8NA0H0opvdxprjLgJpfto4aWxh8NUXjJqb/uLMbkJm1SNsuzmeRx/q+gVacsLxC5T
YAsr7ce0rI23/a8UMA7Nj4q0akgqdC90NIPgGDbpbkm2ppSh3HDGoCmWfhGAmTbWB2QKrjLw120W
lMVwMyvbTe4kHomVWNZmyRv0wRFODGWI1M8icKUBdpAv6srX8DdkC4IDE830kP25BDLKwPtkUS2j
74E1OVv4PpBjiLO1MD2/VSHi8G02wOrGtfwqWG44b8ELWveuyCd6b0RRhaGGMppaWiB1CPOtNbBq
q1vRR5hJzUCctyKEHdJslxrGKOqxkIvEJ05ktHHcFxWJBkeG92jIAHNzkZR2s9jZhU4AnDCyFJX2
9DFsHwiXvf8kFUT0yJKBOzkY9V4fx90HPLDVn+R/SOXqGtGZuqonIq60j93z9onVYzrRbRffr1iZ
UIPc4X/xMZ7u3OyHjh5AwIWFai0KEV3FlIRmt2WXnWNm0FJRQk0E6RNT349DcAS0JhOtGzA+UwdI
MFVhYuire8QBeW7EWbq/5524afJMB4K8h5hz4eVGG/PILEJjxnQtGDE2thNsoERm7lL3tQ7zcvH1
1j79UNdQUcUKqN2Xr+hCjy1emylNOEGr0+Wrn4W6ooiy7D3j8ht04XL2xxOca7Lwz+TAk45RlJZ+
kQIUYQqiPg4Ix/rLHdKjUckut7Mn1TgzNtxMmq7okf4EH/Hcy0ry2n+wiiq5S4J05RSXLuedP1KQ
njP/3yGAocHr0Qn/UbsBkXTR0C12YlRn9J9CpnyvkP0FCRUw0fFJ4CgZhFEPXTCDDz/vrsL/ztcO
1RY47ggwgTlrEPEpJK2SI4Ex0BedWmNPhz5tTTHjTKvXWlAivhiuQwET0zv5OxfsJPwBLAE1MPaH
G3KE2mFdrPlPWI6aQ4WZTkkGEg7d3kKmdNJTfOr7IZ4y8r6MuGPrRoIIgFu5JZzTvbAhKLsou7U3
l4lqA+ecxCUfmUueeb1F+sywgDWzOPoeXT9q0V9nfUsPWJl4DLr8SGEh7ENJY6DXYKcaSlY9LmDT
zVtlF69CJ1Ga+hQSa/5w9DC9cz/vJZdSRXu0DZcmeJ6AGcZZ7J51ymCB44xcrhcA8wizZdps5FZq
BKz644/yh/uRiKchA/JzuKeDo3z6suvcXc4YVQDNNBkPDPHbMfWCUp/UI9PkL1iBkQMJZfqTHY/Y
AToqx7ea5hDrecv1LIENIAzDRQFxUrG+O4u4hscX2YAXciXlem7W9eak8bsSigVeVzAqu/6MklLQ
4NT05kNnIkbECfrq8CIBNRpzvCZFhWiLM9LwMHvVfEoRIDRmMpmRRytfyT4TcjXrRs+IIHs9jQsb
PiryE1dO4z6gsnZbC+un0lUkANjBPez/QngsYApvr7NKa1eS6FjSina8io/x7tT6Z8uxnTL6qlVj
kihxfqI1Z+rk+s2C8ptmAsoKp/TC2m0uXGzWtCByTwrscVt/WximkDc8/vQlYJfOwEj+gseOTfH3
f0FCDMAyqMOPMkHObZvFSwmEe5Fst/P5uQvRRGYADpZysp2yOtCg0agCyAR5qESkyW4K9VvFoeYQ
wJLEyjr/RUiieUjCtEH7ugsG6BBa5xxBVHv4nnQK0aRPlGU36JvPT8dwheaARcfqFS123nE3zEfk
XnxGveBrc9ZW3HtX3z1oypJzm5v/U7xJIfPHeCrBUc1K1itXNA3kD+Rs45CKFpPVTLhzlKceHooB
EjxR/OuC/byn97oYlSZRKnvgyowiLctaKfhFLX8kZyJ4Vid/vu0v89XXU84SUunhon4Y7XWKHd2y
dieRfWHDBjcmGEdWrr6Av44tvhkkdYE9whn24jXcO2uMsmCvwMBRWnb2HJpdGLYGkY/NxIPf42QE
l8nEuSKcr2h7Cd8z5xowxMPCZhbgTVmV6om3GCuq1FvJzxq+TveeJjFHRNyouLIxJex943MG8wSJ
9LPKfn8ZLAKEPmeteDNTl7EQvG2D3+dGvzfFqUmKduxYr3TVPkvxtTehgpBLnuJtflhbYMoxNeiT
Y0jOGDIT4LyeMwha5YFgk6R+jhwcTefmPOgQd98ubF8eRVVnv/eRQVgA9t7FlIJz99XJSEZfPRAL
sKpofTWKCSf8O7PZ2+qZau6zZH8c/n+pggoFiW1NdCZftm2FqeSokyW1e2vHcrIW8bJR/qGn/x1U
RkRIVjgkqPeLWiZ9vdIbQzK2BN4tP1mLqMduei9uObTS9bQ4NrTs8rqpZ5Z1HfK4fdtgKXZYADiA
+kpJH8CxgPlJ2hsvJnKrcg/t27Gx7n7MfdKl9xNPPGxk5axW24wvTUppUdUrGXYIdXy7/7wZAMwu
fnRTuzJmqOVuRi0S18oBK94yb3HRNfs//ROVPRzwJ0hqMuUf+MKuRGdiyE/u1+Wrgr6yxWsMm5v1
/IKZBoT7MSG67ukKEQOZV4aKpSQaBN0xue9UILa2W7rZ5ZqFUbneKSeFyjxbN7T2GZwLt31qSmSw
LGt4iQyx38m6z3ruelE1q13tYob8QCmb2ha9XzyPRde+YdXoOBhWPn+JIw/FsbM7sKwQKqfAIG89
4wU3GuN8iFSXHnvgPPdnrfv2WAeXjKb3GX5pECYgrad2S0FFOEnbL8+ksb4P2dkve/pdcpTqtWZ2
3gbHVi8SpbXaZ7RZ8Lp6b2BXzfO6sVK3uT2WYXmcvp/eTTWnKZpscAyz4+Fj/uXLA1c//grlONhs
gL3a4TQiR0NxMbU741IQd7OSXbVHFhuVRhZ8HKHp03dl45ws3EFHRqZbk6DhPsq1xqjumpj3cAGd
peW2AocAwGZG0NmccxKEFsaFvCTTIhv7Ak+jmucdafNSZ/Dc7GFgDxngi8u0DV6O4iTZj+Kcsi1o
h8aamfzJaTfDeIuQJGGeRpBS2j4ls5X3jBr9PfoaMzXYmKCgOBdOQAZG877jor8TaRhs/brXV1VK
h8vNXJK6VPbfIXj7YNLAAoJHtCFyu9S6gtA4J0VSWnlvYNI6PToxvO2Ea4KexFRB1wpJZT2zmCJn
FlAKiQMnlSqrwYkuHoOCUCbHW31ByZlPy6wUklI6j7Utp9wcaFI/QDgYRpHMWZFyqy0BBV1W5f7R
fLjEAbx5VuY2BcKH0tYQy08QXcS0ru0oACGBK542cy+694vWZsI0bWPconyytoZgU5pd6EYsPMqO
AK9RtClOeIjPiJ0/mA+AU+iNWUzdwmKePOBNIxMValWj++r2lc/HC9GgH3VQFjdJeq6YZDIKIEmV
EKc+UYefrn0Yu8Cm9h6WKbmTpBhE7IPa3viCgg2EIxVci+Q19l6NDM/OwNFgZYXR/GH3ny+6JffU
7ntajx5eeU0k4EuvWwwVNlCUgjM+QwMPwu6qju6s6mUNqQZz7yk6q4vxNl7WBbT/hLZiyzCoVOM3
GUm3MwVl4XH/4Ie1culLfqtv8zNqI5VwEWhgyU0puqGbl7u5Q8EVZOU059t/b51V300daRhQug6a
gYrfCd1sYtzCJBDM7T9KRmL9pxf5ctPOwVwjUYPAr3XboJn6lR/rhhGV+H4VTKHwq9cMonuyAMgk
DcML6MNOOfKKDRI4hZFh7QOTDlV6NJwwRvv73zORYSOLKDGYoJZDg+qMB/SbdCTN2sQpI2sQgTEE
RmB2EXoy/egN6W6Esh+IFm1NfmjFMX2+QehAxt4l9gBXXR4Lm9o2ceS+JMtB57BsF8a8wAlmECUu
XyeHSrmo71/7k2iifdOY7Xx6j/lMpIZgy7Cio6nzf6TA07FJnOoiBzS90SsELx4SeyVvpJ80NtCf
e1PSXnEgaAvyD23bVy0bJB0ye4p4PUxJm3n2gEJATe7gsBWJwfxMJQsRIk+/FGdSHCOyJoCp3hBu
ELpSMhZdPM6n3znDSeF2/Wcjo5f/NZEnDUNqGmsaELtkiegpzPPX3pMGR4hr4PFe6CKbk0+5ZlsF
/dc+DvR3IAj4rbvNuDb8xi7pUPNL7sQfiGRI3dMamdljGA2JI6jAqxUZF3yN6sx9NrHhgNpSl2yK
UdLyfUb+c6MgZC3m8I2/NmcNiXYWdXfGu2dc87AzgUclSPnGljdqbxkJuwpaWpCPYkymTxaypzj/
yfJ9TwgE9T5XMP5p3nnEfSqk96ThFoBNnkOma6hkyRCW8XuNjt34x2clYfU3qMP0wQuCaqR8Y4yN
D/VhBmpYlIC5FrnzoXvjdBUAoUq6Ev52EWQUCPSRylRJ2cZ/Mh93AxU9VvblbgPa1KwdjXAqfay9
fn0Uxd6VxvGoH3XOz4qZkdojXAiKN5mRUknyaM3Bc8QmtFYhWu8SwAXA3Jq0klTTeO2eqStLVKfG
knCsJpsRN2SbNjriJSgwfphklskxnjeoSuSLLafWElxFlnS0d82ErIVrpMTKeIS1FF7Ka3K2ZnmC
ebbR5CDfQmjw5LML+iiEqjAADRjDqalF59RW3SvWsMJp2FtJkWLTSRbqNmak7j/4Clp02IVNDERU
V72PRqdtqYfdybFKIvELT4k3evUuNqFeaNK/0jT5IJF0xBMYC1CVnEsYzvNO/urczFT0O1AKylMA
erQLPAalDCV8C1dd8+DzXLXCkQSFC/xFaY2jacTcPh/qzOKlpncJMxVVIB2B0212r90YObJI0wMw
e1m/QQY1NrBRi/pSMdVPepN1iqnHdDeyyYARk4G1w7uqDoURxey28ZQDjYb1vlkEemfKp3Fb11Bz
aEmcOCJiRLjrX3f1Csw2z8dVSLTgXf7yxKC7qEM9/4sZcSlTFGGGjqYOuBjIFkJOtnU6ywh0oh1V
p8w3K81sLs5FWwz/6qvPSNsqPv4oDJ/po4ViS61tIaJrfeemw+yHFe4Yh1wuVgalTGBggXk1sU2V
NS23Y+okmk+oMNOhEvk1BiLy2XErou9ZzH7mBdJCF4RxElpJR5HI8jIZezIrStsRj5X9xbRF8B3t
/o6tPYte7JIu+3zcUiMQBqcue2fdJrOPlk+PYFqRleZIuePFtDgPRG9n/4gTDJf+71RKJ/LAH+j6
6SfynqB3QneLSeZEqRKdCuZ2j7ko/ns4g+Hk/nsCbb24hhQA6c1UJ/OuDwi1qzlSFeKsMjmV1Wjb
94LzBtb6Nj+X606DMIxbEoG4ej2kAjen6koTKK/7P9RMKsxiZIZKq59m3GuYZeJNhsrFU1pZ4uZZ
OnnmuL4FC0YDpE3P66f5ctC8HzuHZA5V0Oqn1/YlWyT/0nfLO+9lJ6lakHPrvskU/RnpngOPx0SM
7cOpTicPjsD6tkvDNKFfc5kNXQDHtw4jXoJbHwCW7QRoOf37/TybhYyfXogSrxuy4eJ0K/BuAXjm
H00muOh1HMYD+hF6MyO2M4gzySl8SP0BMzYZOSYxntwo2uaK0SzFOtz/VsKNnnyLSEz5/K1lP2No
Xjq/C1rhoBlo+Mmq7YdNKv1aZnWbg4lrg5JCt0ZOvnnO5hHaaYHv5mkOk4o+RUc0KFOcMUtVtstf
B0+qhBBSfgp3nqG4Hlwts1xbHZb65qq6WpSVMX3qqlXNIiSFl3cjdYT1xXViLoBH5CG/4HNArhMJ
IS3lmQxYzXetC3mEAdpvXfi2Z8VJEN72ZGR4i+wo8dx9J7jfhVcY69ZkFrgCeDUfj/0veASBRx4E
qPLBs3Rw62V1pcUqG0yOtJ7F964xLfOY7eJ3zIiuh70HQklGTXO/2QIULB1R3qVPNDhU6YlXy8R3
9zE8dwW+fGWTkHj9ts/qiYcgCkcwNgTBopJX2wBBHE1Y2VJXnMpIauFoE8MV6sEsoXzAQuIFkdAQ
Mel/spMI8rnydV0TZQ3L/GQZHJGHWjt0/mZ9G9eRp4baGC9GSxqBggdrQcbP93VbS6WIDmOiELZU
uITDi63nbl8+QZbhDTsnMci7yKQpkagkW1Vyc0CpqAT4Bax3X+osXQwhIRujTPdr9NF7cIR6aLdb
5m8RvLokDTxbtgIGd/LSfA0nnQo3hIUyo2LxC5HyVB6F5bHgagIArpgigwMwAtjh60anHgR03Ouy
xaVExFUrrMCetbm31vY2dHpICsU9RwWSeIEADbnIxf9UGShQrJGVOVK9QYm1z2HzuzNma296KzVM
cpT+tN8Gq9CKkztdiV1jHXoHC92cLS8qMuRvVepVyYPEKWvKNVEVZ4a5pOMT9KC8piIpv106NFJp
r1z2m5AFz14xLmLf0uY6T2JWNHYbAKEBl6VoGKLHNit1D7mHCUREK8l4Ao9/3m+5xsJflcTnc1T0
cWyxCKyY4M841sM5CANjWkGsalDm4VmRsdu449z0YWMY20rLqf31SkfHTsEPI+Mb30R0S1Vh1H87
uLDD8Zu8Jt3MD7V+igaWvvC4a+X5UpK7m6WVG6i0XoKpz/mLYR7TjdhBnv6aLBDd5vwmpdPSinqk
BDQjsGiay7IkWKbglQETkpGXy5J1bfi62cchdfKtbqv5LdZyEv8s7MlRSOv15YE/bTQwwrkkXHSe
Zzu3NrrR6kh6VImueWZKtMF7VtiYp4L7VoDm825eA2fRJ7CBQohy4wqL26zygTcBvI0S61veD6/t
5crIOS4PXCBrW9KI0KOyz9RQ6xcybrkXcdmlPztcI2NFyOUtDjyczfecX2I/3V4TB8YikP/Yrvcm
1mNiX+Ji92BWx+0ckA5u6o7fmNfnolODXEQkpAnJq+1xz8K+sZOCDLQfmsumXSSt+44hO+R5ht1A
sI51kzz6Vr6huAJz8vf5TM773kHFYKMRr+/dSQk7tkGdGWjbrcKWDHWZXA/2YuixcXybr+Sco2g+
m+z6lPjubPQqpBWVwpUHgZjtX/T+WcJ5PFB0dOcPOZichgzDSPK1TCHZNaAuWGRKcvKV06bQCvNu
T4la3HEWgwN/MHAN2MRh/YPLC6yC+0aQMfnyUh/qsK1aiDtiMh0sMrQaRO+qyT54a8gWgcqCCu6r
qOxCqFY8mV78AEnfSAapQP7XgNDmy0fzNcjj3BEOMNxKtg7RKvvrmx0N0ebW/bTozEJX0vhFJ7Yu
+RmTg5V51v25xNztGNhez39aa2Gt7JkFpgz4sEPWkJuMbkYgVwA9mDDm8+iDov5gAj9MHril2zuy
OmMoD/CYXF0DOAdWUffdAcyBUY9sipZ403xwX8QfY8+XAEwSZ/mDaVzJBUwY+8n53zbNxoTMBSYe
KAEDBxXHYFZpwA8qoGdjmnFYeL0QSs/3kErslTa8KbkDmaqIL+0H23twYdys0/b321rR/PPUSyFQ
0HoPzrLNvmyUl/02JoKJE/sXWuvCRSXZF8PL+QXdq50l+15+Eq0bFTC3D9m4peSLodfquFNnDTCQ
E6hPtJYmtQys0ueMK2V7JmYaW+OvtcY8K3PaBpxzIv2sdiw6DTYZ9ERx2jx+qxenT3kSfKwJILwx
cBYfy85MBzbskbD9thCtCbZWzC5M2v0FpZUX1uhph2DVYfd0K1j3UgWjnCg9ZNMKuBRHigwQsQ0u
wWyWBx7jU0YeSYOeF6rok3jT4JjCDyt1Ou8zoMQJI/69Wa+I0aS3lrrfJVMjG/EWeZ0O57C4TXxk
Gvrf2AXjgBqYpP76M99rYiWRqqIJMJsCv45Zq5njP8L7ZZujOQS3VfXL9jIYqPXnrvcbtelm3Hhl
SZfUB1L3zJaGFcFtAadKETbd7c7JF5wMGCxFwO1A5WsKrt9/T/t7iaI9GfgtR4e3I02MLDJyr4ZO
F8Je2+i2TumuATjgzs6sOqyDjjGcPMNuVKJFjAuqC4EZ44yfadb4tStInyfEEN3VeemnhsHuofBc
fHzP2N2JTSmT+HdPJvjGZzkwXY82+bwbGsqfulpQn/vCmNbqRvzKMEo0tZNNS/FMIGfuDdjsipdL
flY9LUpYt1cfJBpwtoqCOJdgtDgdoEmgm0TP4ndZf81sKL09nt+di1pYamCnICb+V75plBXQ4Z3y
c422HYUMqj22584W3lbgi319ezbNBU0SdyP1CEvcQF6YYZOeId2SFi4hr5lQ3+11Zmnm3KlTxNfx
r/Yjk0XcQW8m9pLpOSwYGSG0YJsOgdiguXfurfDLBqPkbdhcdM3I5Ms8d/OKgi/qQJCkd4XCxgxF
4hEQoZ6RZvTScxZXc62e47Qm34qBAVaRTNK6r/wzy76a+bxrd6lt4RIPh1RbVXCTjOtRQ+20g7cJ
QTIzjAj6mZF4CDdlFb3W/r5KuO/is+5ukr1hUiPalSfOZlj7jCuG1gvB6jw2/yPg+L36DYouiYcd
s3L8M770U7tWe8t9eEj6KQ7o+zjkhdzTwI5mhrfKidsgYn7Pf+axlRYzxT/zSScISmSMyx5QJcyd
6FIVgO/BcNMktGTu0EQ/R/OD9A1mrhEviXNgOTdD5fqP8GhioZ4kqzegLzOmJk7ArjZV5mmDxurt
G8clFNGp2ffiH1QDWEzZRq1m712vXtuVZSsXD6KSrr6tp+0dPuI5Trw+uy3oWGWiRELnw1ispfN1
vaJMcChdV7Snh6eukydbhwsn4QioUQ32vRSWxEzZgh/zSKU9/GHoAryFLSsodwtDD93P758UBPxi
drq9y4HJSiBTAEk45JNsMM1g+EVFgqV/NjJYubf7wseadyyAW2eR2Z6F8lmuqT9qka4QP3TGSqNR
4RGpx7K6EpErA37De/eQ5M4N+/D/y6W+nJW24+Uq8emftcG97XBQBtiOaSJlqqx+jnrWEbr4Cdou
eRWi61Rh3WQqbh/7VCmX69aTJI3EAdRxS91cE5ffB0OZTBjAi+pBj0NXz3FylsMwkERlOFQwU5QU
eKtSmAwZJJlTcSm3aSCZPWFcXBnaeMMM4Vf8KDP4NEwk1nu31rJ3NRGovG/UGeoEYHLvFJ7v3aQw
rQMWkyfTgpzJGcQnc3NAjYRGB8B/WEq6F2jinbJ0NgCpcK0wdNp8GQ2kKuZVEtWQ4OOXIhD55N6j
jIIvP5qKIOKB6qVl4K05degNshlcrce9OTS2Kg/fFNH0UOyIIQsAMDc7faLpzabkXOrx7abNbP7K
QLA6HpBQ0WZXi0z7T26p+OChReqYxmosDU00pfKJ4deeDJ6lkQYzawqF1WLHWqE0hA/q+RL9TnvD
el0TnS9KfxGsd1U7MWkO7mNIwKKeBCsAssJRy5Obc6HuWWoMc5N2MVPsNqwUt7a3xUXV8rz1Epbd
u+Vd/G+Bvowh3AfZRg8ZJDHnGEKqAUy6Y4rAbtk5gR7PGsEEItzmz8KHj9A5xHIPWxx+1/YeYKK+
zVSkbVP/Yvo3/9c6Xfh6ivwiaQFcTbZQXrdk2HqFUEOj5IC56pDm8fB7/tWrtUPHGjWXdi8/ju7V
Np2ZWiK4uObgIb9q2ijY7OIaoIj7jO57quRTQzrNNIHA4yv3lW8zMvrW11wNulf8XvbAJ5nSF1bV
+Rfj0MkfPUWH92cSkNAt2/brpjh6JApuqmSVRiOn272Wn6YK5cxX5DoWOjb95X+SsEbKwHexd8yu
LgPZTWFot1+DnVrtdVJAbat//SZfwTHvzGh4pbP9Go4LKdbKYY0/b1Vsx0qluKN1S7qw0MwKjTNp
2Z5f69P8iWl1kjhcCts6r2tfPuVtTgG9PNZHLR1XxYK8iHrBi2eRXncbvNfzLtDop4mPuoSc5iFU
QmuVh9/FV5XzYDLjfVc0unJHxzpgdM7/ySemfBXSw2aEFdEE95laOTg6ZdKOxbQze0YKfLw0xGu9
jdLvtw6W1jgZhVpUdqK3O0I7dRU3fsbRa+FocFC+s6vm220uSUy4k/TRZJbgD0hAkkKnpioYBBOs
DgmwtAWgzfytQkj0/KYcc66j1rXPo2Apy3oPiDSXre2/cthicDUSspGdU0Zl+4rUzJi7BkcYb01D
GqK+w15qYGpdo0qU2TRiXVrKBYXBanjN9dHbjvnwdP+4A+Cih7iUPcPnih4NZV4K4QpodO5xD3r3
XWrQFYQP88FRb8XEjfhgRuzZCynQFvuV1VxnzRJbArQVBv/mTcKznS/kxuIBAlqftR5hHK4Q36ri
LQGCo0Lg1Y2J/lsRAArJbA2c7tGjagTx2g1XNLSGOzpCLKPT/3Yanrq7QdDUy2SwsE62p5VeQv7x
rpnygeKEb9ktZIOwEUsezsZAsnLHvs+YkK/lKJk89MFUOzYz3+R47q0/uB8MNPZ3xINByuYcxEbx
bqqxnlPBzWV+vc8YCdsF2G0GG2TcDSvGOQn5+52njwd4sTOHc+7I9mpAM6D0knTmxZrOLmBwHdRx
3VncaWQHMiNOR6J+vS1JJXw+2yVBC8LewRc/OZxrdt3Vmpvn7YsTOjoFnZUP9MlPG+u7Qfc3zqzX
7ZmhWeK+uuEhltBet673eTVcRdymSiaMUKaYJZAL7qfVbfrUHIif+Es3KfDflkoQxl7Qb3LGaz/k
R/tHseK63L13m+VWeTC8RB1OrhlQqhKUCw2/M9yupeQ2hOsXbc6VAD3sMht4Lrt0+8t05vNgQ+NI
pfxq0pXmbm3LwWKabIr+Y/WOvpi0eGvVaTMih3yRZLpIE0GvRcanccLXJ6hxMaB3q/t9tBDikwq/
Ub+YtoEEhxyxnEEcccNgKFRBR8y1lKCH+h3JXEHKQ4LFDEK4vkd6tPhqo/dNz33k3Hu+3SbCzfhc
ZhtNVdTZyo/pNreQ+P2salKX6Nlrxklpoj3wK3mbW7/g897Pp6VIqdb5NDgrfboux0nCXu86mdoa
HE8Qq3uzKPjHAO0uGXsfXc+nzXdsBtlW3vio5upHIWMC2Iwi7OnTaHQtAUPlRvZjQQSAeeWHzFf8
gS/K4ZjLi8+NRJk5Uezb4+cg8EqcNY4sM5avTTBcWnZzjZC17yzVY6bQaRodnyZWqi3/Uh2BLqh5
yDqV8us2cjc75bCxBwDW5P94AoBO+nXlRuFWEeOu0NCU73xml5L3LmXI/sx1hPC5gI5iQf5dXvWz
gJvKVqaaQxqD0+FnkVnnnhaStmRaYe93uCQW26oByTCLNV9mK1/tJB2MwzuN2LpI1RSdrVz7wOyC
4AS2/HvncG9GzFCZ4EDphGhvU6eY+QpUcvxw3PXwW92psl/Hr9/dNxG5Y8tBlAuZXjm6E3XFGihq
Pg3U+vCcQbMM1KFzeF6mP1FsGZmhOuRI7goHq292F5eU/djOBvmcpWQEbxBl/vkoV/CEoQs2wRw0
mirXlDgd9GSb7+Ey4+eLqKtUkPlPeGqrznZChCBoW7UWQH+wf1DzhKWPbnBqPAzBwXr6eifzFvK7
2omV8bxy1DLnZbVTf/Dd2n+lUUX54BDGPskcyg97wr0cUmyspNr1IEiWTCbJ9Mr9q3C5320YxXpk
eMwYiX4uOtj0omqZUi2vFNqWIjzGJL1swm2G60ilmD3Qx6qbVvOJBvZI5LMjoYdV93iUVCyITmpE
/yg0R3XsljlEJ+85F93Mm4EOtIlTvP0JlixDLcGGvneF2ThuZkBeD8AOtsCKwNcpk8BU0BeFu+yz
GeCMpz73tXBRdi+Rtd3PZC0zoMBcwyobjbAoN2Z9cUXsgAzcRjjY1YCz0kTVx985oheYbwnA/wvX
3DARxSpQdiGkzaumBMHoq6uSX2rj7XaD0NLmsdn63qI5Xfs/2PBNwSHYhuP9d39vkZ2CCs1rNG28
TnABM/xywXyP1C66yaNtCT8ZYnEc14NdWwo0zFIAD+GqpUz8h0/Z/H4tmG6zOjXnWea/QlW6aHvS
CnA49QIprrzTK8Cro333nlRZ1xzLaFrH9TFHnnHTPFlddzxgB/4dM41pHy2nfGxQeTCStBtBMVoM
7bdEaiaok76Q5coxz4mTdZV10FcodtKZwqoMqMaM/FLKGypgewt++uXK5kEaAMU8ot7OEAhRrGCe
Y3U4Trs/E1+y2wUFFs7vWQG1NUAXBvSqpKJDPfIWpYCrOGF9K/42Ne4cyv1ZloKu4rFvKnadSFup
U+LgiLc0urHS/UpaWajVpRC1iG0itYnkUKa2zERY9kIa0r6wzOOLgDYoKq86bHtiHzrVk8exvxYP
Mutvh3J5/egBosFN8npxflccC8dSQx3+YD+vAvjhdMpNjiICrXF/e1FtFiouUFH3uhqQgcYWmimt
pOQEpZ+eyhIqtdVkYjN/c2d4ay6yRuOuz2J1803e56yCX4GqD1nf8XMT4vJmx280IeYBq09IFAnt
bicInXbrVGbEON5Wnb3jTzNHgY37at1yDYSiU6gDM6ITvU12RVlTaHSr60BwcZiHgecZfk/H+eL6
aicvlWYJnmpH11DbQnP9hoYhOYr6I2wzgAhWbhrEF8AGa26WJWE6J2lCCp5xvWELpCxY4XDMqB06
Ivz9QdCr4csUp83xiAvjNjD8pgl9ROGCq5BXNnsgnZxR8VemOylbcU6AWbnbcRzikOzxefTGmmD6
VN4qjnSfoHVvL1CcPkKXSuzb/MFFWour9s1dBiMjsKb/qkoznyADE2elKFEuv6D1jW9rwii9f+CR
a7ZE13WHBZauRjzhqLvMGUveFBXdK6ghXxbwW1hmVHobfkXEyeaKcI8EKAdfJGDS0vSmSXcVPAFv
otTH/3xI1xBeLtNcV6HitDjiOCaqrPzGI62z3CdUcw8McrE5qrJCFQXXxHQpgcn5yIgjy+3A8DG6
BZIQlTZgEazGgYYx2c6Z4nVUq/VSwvCJYAuDNDqUkMmNeImiQxgAgs+OeC2I6bP3W496Wp6CEYGx
QWh/kfbOJbvoeDRbCR4yudroZPQ6wDgFyQbblAUnG1tdJKFYr6HA9gkAHKREXXsnAw7TFb5RRxff
F6KTwYhDQ3HSdXI/SdkR/wS2hxwNpgddkYY2URR0Vn44pg41Hk/f+9Tug4SYyymojNMrXHkLCBmv
T/tP90cW7PEFcu3p1pvpuNhG+wv02F9ILHLboxYHtH+Mrqa9sxHh0XdEbTqn/vzUoKoI5T5TyfDX
7guakJIgZ9mjotHFTKC9xsnCAASmWwkbfPaf6oeO6X0POOJc/Y5svUUKL78je03GKkW/xvOU76dE
XDMsWij9cjNAtYRczMk2iBgcUQ4OddvQQpg3jYxSy2NN067EApxcT3UHDCPEhuBiE/rAyUGEzfel
JmcRaxr+N7zmI8CYVCm/HxFIcKZpylecApt5GuOhrapdTXz96tpDUYVIg/DE0gvn9XurP8zQmTQj
U9f0ZiDNyX2Y3zY8XR3sRrzDY/wUXZae650eftYYrLm37CoOwKHTbSA2iuuIp/MoGOu1YXVfYxxH
jKLKCSYXyn9Fr8idcE4bhDIEnhwoYhvLn9Zz7O0ZeF/sOrCDDKZvfJC5j+705tv349TzVqmha8zB
+A/Z+SbrP/uFhyk/XRxOa2FJu7MxX1e0EUDOxISJuXU4AYCWHk8nSetBpkCefQuZxsuZmwv5WGqf
VJ3zYNS6pZAtPA8S4ab1Tn6EyUIzqmZtp+J6ym5vyLMKmrYPG5T4rHnxE5dmB+t6HGBpxTmBD31i
ZotBsyqNBVbXmK8vIkEKSNBd3SrySg61itFzZ4wmxPHJHMwlXVCumQwYDiSUgHZ0gpUiuRPgDK+p
sgBKYfmpei5LPmnuz2CCt2EFgeoUmsWtHTOOJMZsNziuSoYn6i2P9fDYRlam570MsG0pyA6fIROo
egEZufHVEROHpveU3LFmcfEV9jmtvgkQV1iBhOCrcisHhDRGCdTTCmABR1AffEQwJ5ZkYjNEtXkN
UlvfxwtkGRCH7HOA6VVzEPMJqvW0WcejBFJK8bpP8W5leV5fFjKKJyreS/zuSJtP6eTajZSCgB+0
qVrPPNCw0ddqDysKaqNY1CY1jHO8N3jgIG1lE2ppEf/+fo4tJUIpzUxvij1s3XilwIP/DD337lVY
0mD2QYhk67USzMLyU8F8ATymZHC24ARDO4vRLJwTY2LoJub+xKM/0LYgKPB7lNzB8XwMyb5VAio7
3TXN1+ahdY+FVCimJuIuiC36WyEx26mQWgnhWXCNFgjFuFEokC5S0Cv6I96Q0n0CdN1kD553FZdE
qEoAuHK36NUF7VN7jv/frbas5JqKSm/NL6C45k5Oz+YcrqDbJIDUfOxdIMCaE3HGy97OZt3MTe1C
osUIEjwQGKcvDjfPPZBh0kC/PKycVRdba5SPQerN/DOdiOL72pt0gXr6YHcx69HZV4kuyMT4rkZl
MlJ7MBfjwQjfIGbZn4jBC4cAgeZ9Y046sG0f267YDAYjWTIVda6TC669NGBHwvGlvpz3Kht8laXd
T0vyOKKRP1t82IFG4OxhrAXBDZKnwEg394dVw5c0XmUgwJ6nRA5t85GLOs+H90WiomB7eFW+C1dL
Amj8gnWn9HywaYyXlY3Q8FS8QKy1x+oqwjjGMFpd8JXIabNVTuoN76KEGWgvOPOyiH9B0/OAarf1
hCMo5AR65sgnOMD13rEzlR9OJHbwHs89Wd2+UcH1yKDHSlUF77eIOEjHPLMgqOg41D8mazWfZPX1
0Ks3JxjAM+kOJRzAcvJOYkNSegzehp5JQoEorFJF4G1QWNfGeLYXCnpO8lUIrAu3GxbnfEXSIvAD
bU8WfigQ5mSkpmtaMsfM6HzoBgUdIRlrypor2iQgpFMMheZ7M3yn91UvL4nIAZwNgnp1jSd00lvf
pnbAs5l6yUnZiUDzrNpL94+vsdys76E6tiaKVcHXdVkbxal8oO1pmHHqtLoboQKaT4fjH2sikLje
fQRL3gfAOjhOYr3utbzne28Z/whRccPbCFK9y8et0UU2h7ovsASUEtzLfzgoLkecFWe+rVjwCgtJ
JroHpYNSikoffJO2mUTjAzZ0ix6I4Pwjf2U3rn6tZWq7QSXCpPz27P4MkpSJVRpwUjQ+2XBGpWzX
17WBK2eASVIKtENX/f1IzanPizQWG4a6XQnSXXcZ9Qse/b1LCWKgeNvESORG6d2HUWSCumtr66cG
C5zei+4ecCOZ/WvHdcNVG4z/8uT89B4gvUaAxvIsmtMjxextJQrD6wCDgFM5oHur5qh+D6bXDG3/
/3F/tphnBFctbyyM2Bzbpq+Ik0ohesKJJKUoInmfPHCMn95Pgas+hyggwrUUke35WhZBqUdNeU24
JuRCrgdlX4h9gDDeLy0RCp9mFsnQ/QyclNIcMKL8Nty/WLTqfg52NQH88e+pS1/ah+UX1YXQLrAT
XLCFgAE+E50W7IAcoCvG3kIIactRYxgkd4TbDbcSDAwaT2y2rrmcCMh3TG2IGrceRtzkSvMcCO6X
9jkwBNJFTN1BgpLfziCgedJU8bG8Ixt6nZlUZd1N5zNQyVeeaSNJ3d3gFQgAJPG8I+tfEN5wqzDU
shoGZpr3kaF7EuH9lG4X7JZF2039qk+vutNGUsDRk8qMHFDkypdw5v39QmQVCbJ+Yw0zTCg01uaS
f5kF2PoFBP1hjAPbO4DcHa5yNgyOcINpd3Fm9Clrg41bXOf2pBfl6hSgCfKjQW4kmXfkC55oxKE3
ukpnQzQ32+/UQiTmzcgd3HIZkMPWCUc5tleMp7cvCPA8qSDwwVUBl2vLau8HU4XEHCBYbjIzgbTp
amecjxmaJb11/dsImg0Xyq0ibEPXyeryyHPtLqVtIauSS02WUiQxiLZWIAGXCBu9s7hD872H7d4T
U3uJdxqtJIgMrbMEqttbLkYQa58lUGyLUPopojSOiJbdSB17m6XPZKqfKCUn2HOVQWQaGcjSUVGE
05EooCZtK7sQFvqLlAc9iTv7qSy8SWbUZliONzfHiu8in10Kg/w10P0FRPyQFcDD4DoA9IgAne4I
siZAZ+ohZp3XFOjtPxlNU+vJqqSiI4+NaYukhtjWNedbearRUYkmMIIbFPrwSgiGdh1YMZjaXQd6
SUIF1eaRoni09NvHzxPZJuWFzVKzuFw8KChurf28EQJIuTKUQHWM0NBgDfVDMo78cU5SBW6k3ux2
Onlk01oZlE7WrVjmZpNJFvkKa/cOlzeDMqcaiYLZuzpEhz+6z1U8i+M7dL21f1MEib5/1MB7E4Ys
HYPthiLxUOnLJDIGGzBGgw0UHUPrPV+ksBF82tEbiUyOkfcLEJR4PXv9bm8U+VfXB5t8Kxt6Ij3s
06FwG6dTd0trowntsd8epPoMxq3GXvbrNZvLfRV9lOBVvqwC417nJf4gE91x2vyTiSIa/KgFjPfR
m9jahX3sEW7EpqKbFnomaZRaldGC20c5qcECpQGJ41aV8iq1MWjwDUotAvF/jTB2xayw7MxKzw+C
VpqUMWbQ8UU9/FGiY7TbvJBjeBd6bVFMHGtyfVQECIaG8h9r/3TcLaigx9WtI1m3PsdKM6AnMoae
I+gNuDjknb/tKIecCXVC/f4zAyOTYnfSVBZyPROjCAg7V007iFiFThyYAUej/4+bIHJscInL53iB
PuEZ/Ds+rgZ0Iz8wAXclVa+CotX0f/FrwD2HSrcjltoidDPVX8o01Ml2/cU1617iNT2hvjK9lDSa
wbxF/TUfND5uvH+knp7d5hST+aXKzdGdK/ylD/qcP32gjOqymzuAunEO9oOGl0mlmmCuj5GSgIsD
NPvG9XTxdugN1TLl8dOLcgmRubNN+z92t+lmKix50emCSI14+jVDVbhbHBrV/gECvaguGX/isAVn
m9xN6ZoKXUYiAdW6tyOU5TsOp/c2Y72xDRt90gcirYG6JiIIrOA3g046YVJ3t1nAr9iJL4yNDxWM
dZJqDGFton3cTOYZnkMM39ZKLUObXVKsDgqxJrK6iwBE3AJCU8yFzlRI0zZ9ZvuYEcMQoD0TP6Yv
/vCv94s/DT0b3uKkjDWmsU3RGomHrCJjGb9zPW7pSvNHKb31IuULvdGtx0PPJMvgnC9Bl1O3AUzC
RYrmyI1iQ9y1dsHOfaVPe8DF5zdfGKP0g8rwr9X4KBC2zaO+gGr6u3OO2XvcCBXu/FM3m+ky+y8a
1jGePQCzixB8NWweS4ymVBfVs7Ooj3GbebjKKkiqnVzDnA/zLGcYQG1xX4pB0apXJ/A5/cfGcwr5
Dbun1FHy7zIO/ln1t1Pr3NGbZGbUU2GBA8V7QJn9IHz90HLtJvRt1uEcno50jjapMtorIBT95SGR
JCK7USoTrmLBMprI3bKNE7V/PFgfR4GKFNQBiYPiAKIYWI8nfxjKn8lTEXmyaMBOHmQ3vF4cU4P3
efNX9B+hQxv7PhKHziCNAc1KzIb9U6rNtIUMrftcUnmVYI2yPjk9d7414hRe8K/K9KvIIELN8qg5
y7xBFULRRDVQGS7LJzc9uQgu/KFZQOqkOowUcdsY6wDypnvhLVa98bFwwOMBuoOKM39MyVZ/TF3G
hb7Wz7FfOTnS6QptlscMYFPrqyJB8e6irY+IEL+bDHsg9bfGa3w7eTymGZ952jv/kxWbAeY9l7Gb
bONKstZoxy3SUVf2Ub/Q39CQx5gRd9Pu21BLDVZlyJh718aDFbsJvKPY4tfnyQhMlhmaAfYsPul6
rVWyByQR/LKb3BwMa5DFXcEiN5m5BLz/nZ+wi54rZdbhMYFxVUkP/X/OXAi6mPBs+AwdniBTsM/D
76X0yuWoGeIry30iDx1kIm5Vifp5lMXpQhh7s1Xfifq4602+H6g//lo7L49E/+/S+Cec6Ygh+Rgh
gbgCE0uF3R7rF2J5aGh7pMihdBL7mVuXmMpEm/0YD+xqwp3jgr8JtlgS+47/Iu/WwD+0fEVYJdKL
c0q/DXx6/lnJRKUVrUf7Lc2mqwLXCIdct78Ezydcabz7neSglwLiKnaB8Eg4MojhImhilvJPLeEt
8yvLfQnDpbwhL7jJ+YKbW64P9m2mj37QgeBZb7G+XzsFnOp83oTtCo+gcCIT/KN7QxzcBaENnATV
zhBASYNrQjGwbCuLuQZYU/WtcsPVtLPoAGAYW3Katp9gO+4B9UlGip8k0TEe4uRR94IPvIOXa9RL
Mw6LIdTJQsoAs8U19Nx+M4cmEuzAHxC6GIFY4gXGwYyU1P3t3YtqGTU1f2ubD23FGqEkkeLujs25
0dBS1i3jTwBez1jwCJiNQPTDyJpmHxxbqMClhewFqH9lAXgyzXYo1XDfKGKq7RuCt9LyDjc3MMEK
6AaKBnpzfSBUqKfChnNJQcfOg8T6Igdf3MLthC6H/3NvQXoOcpsMcxapmL5XCPwWtJXdD8BO1nBP
oESjspE3mfGn/RhzDJS/PQNtObho1CFV4DrsdrYDxZR+SzX0LAK/3qbDGhzUsYmdnCdAHEembucU
CgqJKHRchkaw/VtSpJmpMboP7AEa5f0vkIwkd5xtfdDAPagGnVq5qKPSkReoymvlymvcsrKGstau
wkllF2swd+7nAW5VM9dQZOEdW6Iw2GwTMpB2U1bAzz7bxKv0z3SMlJyCeCfFdfT9z5a+8SsXyYH2
FaW48LUNB3OgGNjniB3v2TVhOma4j+28Is0BuY1SgnbTu8vjK6tAxv8I3lN8UVaht9HOient1HUt
EnLczV1G5NZ1S/Z0PvxrgcfOvJLbfuxdzkVyz9eQdqaD9p0f+Id3o1pOgXhbot24be0eoDX18GQp
YYfun8Bp+kYXgMzBzDdBLP43sBZwi5em8lnXBAHOhnYNQNzRip6ZgjkQAiM+gKVPynm0jEiIWVBq
WuRPKswlwk25ohsTxCPHDPg/bNySB7xhQMAncxTzhNYmD0tMmn15+5aYwIhNDBBq6wB2VkzoRwSy
XshkJpwaoAoDsJvTgn0ouhCNXY8COLLcKUmTyhTi562T7x/1AAqceJFio2xl4oZpyKgA/UoYioZy
GU7AZCaYJxI+KZNFE6le62dshiODj6NGr5Z2ai3Jq0fTQRGVZKFqfvJgIMMWIqxEjHStX34f7IcN
6WYjJ2dt0BnBvZJeGHXjFUb5FtuUflDEUJsURakcToealehmIBOj6h1VD3/pkXCX1ZI/q12g1HMN
Adp9PAvyGfhtJrYinZxCaexi3IMmh3/fPHF5VwwLS6mzqtojqBnTGUIHEmgkVqo7TR9DLrrmSSbC
ouq7UA2Au0d3qDyA6Mim+1wMaTn+LYryPm2rfR6N2JnOZgoIbv1u1aIMu+mSQ1Y/nibEOzx6S1Jd
M1KY72tyKUIM/CC37uI87Sd6SOcfRvtHsSGf7c4+Bi9sbUr2aZG2Ej2sB2eAO6htvkmsorvNoVTe
wRt0u3J8B6DjJOVYuFK1pWxhavMCI9RDENpXBC4M+1s8r61JaoMQNm4ctYBP2AfHtqOIiHA6Exg1
J4ZHmS4JH/1NjmtNnw+AeqV1F9i5AwcDdVHiY7yWArgNolBqg2JbTkRbdN+15abCU4dNdsTrq005
toKd9FFtaDsU9x4Fw3YirbwJn6Z2ec54Zm0nPDnYOtnrA14fBAPXFjcm7x+s6ycF/CVrft4oHAVQ
uxl1oLe2r8gVlYqfHP0nkA0589IOe93owRQV7TAQEc64h+Edu8r3NfGiRRyf5m/XpV6cvQAZclgZ
Nqx/hY/LSsS/VMv4OlgFTc+Vgnt/8nZA4+J/x0OPEa9wYgBK6dPQ0A9jFORdaU9+5TZFYdPuvRUu
BUtNiBbzaNeuW0alHyqvz/86u/nbK+1SOiXRysk4mHRIVIj/FSD+3+kaMwfZejy3uuLdyaPNHJ++
6YFNO271+jcfTKUNsYfDog6na5mT73aOVHdPLeA48JDDVN75dtBK7ShvL4ErOWwLI3iyWyAPOlmy
ZmqPQAC5dKaN8ANidmG00c0+K5uruBwLA6nhhTXQ1/qi4ez/4b6FJw5q0qha2aLjwZUBmL1wvQj1
Saob+d0BndNfRJZXjs2DXV2JY/9WVQ1oWcIIswHjFCARfVkdjaRpf/+iV5Cw8zQ3v/U1M9aX7nX+
vvyo+1oPys6WtqUv3/8eo28eIVk8vbU32IcrcLK/RawmyYe5ua3kjZkSzJYjED4YCxGGMe6LKvoG
MTSWREJ7yRCeiDVbjEi7fd6Abiupq8TCh00AN/AGSllo6o76IfVijdNowbNN7bG5+vRw/KWpj5sQ
bXvdcFO5AaRU2s5ju/4lLXCIjkrewNgX4WTb+4iYYycp6g9w7k1x3vlhSbaplUabuRAWsFYZZQiV
/UML9Pjtni9hm/4+3mB1YgP3sBRX/vpHhnCvwDu1kqmpmMNYRSBnAchT1rRxvWv4xsqpDdQnEleJ
f12xIYxly1Z52/oejguLYuW7dRPifu35YagDdmoGq4lbJkJQu0Z2R9WLyTX27fjvVCg7j9gw5aq0
cRxGPDqmkl2tf36TZjZKvOs+25fpsoPYEvmguonQBzxL+vaMbgfKDY/LNpv6YDhn8tAeQYlndzp1
jPot8eluWlgE35Ep6I5fSkGDsxjv/B/LpKEOQqWjqIMY5oZXe0UOCjoiBqpKuumrWNZ7FYpP00AM
5fMSl6ZAxjUMt07DXos1Llup4kOYaMoY/5Szw6MZFAyf9PuYxY04Sut3GhlyL0pTJUN1uB2V1EAi
u8w6on45boEkgVp7b5bQ205bVOCF0aQ5aOqJ7txXMgKYjqgQgdAh1HYdPWytOu+DOO+fG59LMNzM
dhAF0RNMl3vpjmY46AAztCy19kGv7eysl6pBBTwi/yQ2ypSAgytFplcw48gpuWfmVAfLDaR//M7U
wfE/YRRlgwPvdrnxogLKKTdtQsSzUx1Mn7jCAT+7/4PZ7hWQwPlmUIUCxUqK2ax4gGL9igi5yuLq
EZNXUkBTIy70hh7EpsLCsGPTMs0ZKYAjJM42+TnmZq05wtLl2lXXLRmJ6RN0A0ZDFYHMXgbC8Tus
tkCqSauJIbQPvfq05rC8zgb/wUVluKyCWosaeCLV9DZAfaDF4MMV5m1sapq6lUs4eplQClN685Fr
8QVDK3EKahxkeuiV25mvgoT2lREXhE4QLPHmDJEuUzS0UdCPR5FRkNX8dvnBdOFMHWMl1Xdtc2A/
+dlM2jqL4xl21opbJysBDZGpHR8YGrkfoNIvzMyDYR+G+yDrNdKIC+3V2gh37k2ZxPUJgUZGiZfj
SaTcql5OBv+Ezd25H/tpva76vKoZCdaJ6oXsHFsTWS9LYdF8F2536q4EvXQ+0Sv5lsCkvBE8JS0x
0Nasi+5ON0NQ6gE3UnfpenXwN+OzvjhbCnxUYtInc9chHmB/Ng9nJxAl6z6WbskTmRHo1lRH5YY6
6GqkGesIKPTIhDYv/nWgCo8KGh76xJlkEwK+cHMpIXLoao3wEjqq0mxlNp/CIalGww3ZGOkHgk4f
5+zEM8rR57KBYJV5otbZRBEIzjJgcRwDogvSM6SRqoOCUjMsEfJ3mAIRUE5EV2ej2lRX9wAJ8duS
N8Pz6wzXIUdYkW25Pq70+08bXGb4LgZTp66rW+e8bMddb4K4PX/U4OZT/7QCqtNJaMsqDtHoE5ou
8eznJzrK8uB4hs9gqwkSsdslNgFov6MsZPqHZcYS5Zl7J7XmyW9xqz6QEkUSknMYAnoeISDzda9y
F9tK9WBT4VsFdDf/uY6Ad/JxVuU7lvLEZ6dh+TPI7WVYIq9h4EZfG9CmQKkzrkHTJaJHaCFGHdxo
fkE/Wfd02tIZ76QfB3Z69WeEVBtUQBhqyY/BwVy3HxroLKY5lvYFknnDmL9JY0G5Fb8F2zJSMnWV
fKq6JaJnIAfo6thNQW4tiYQ5j6MAhchu1HYS9g2b7UXfMvgYpqhPRRQ5OXMiKV8es8RAaasrfey5
zP6W+2A5VFlcGMPLCjonbn0ZcWYeeSUa/gs3is+Fxa9lqGbNxquMB5u/Tkf/G7hIQy9z1uLrfNcl
Kpax4jWaJN2yhv6MzOIaahJkjRXlMHOp6cJvb6vZ7hcvhJuCWkj+T1/Hi5kgChjtjfX0qgYNMG4J
Ap+gyuU5FOHV9UKWUmQCS5CG9tONolM/GTVf70OV7uLHhn/bgMu3zXqCMGs5TCJijjUvDeLbtA1L
fjLk6Zt1Lz21tYW/aSIKllQF70fpP186IfXpk7gUyLZ1Z9Z1HZt0jlPEfgT0XGYRmjsXsZQCc5Hg
mMH5Wm0PzleC+uQ3thDqHLgbAoN6yn0SpZ7GDb8Pg/PxzicW5kjdzAvUgyFLw1WsmKQj6XkbZ0+9
Te/TxIwHNgTcZMQd+RHhy2l3bduOxWdN4IvByzDZOiKcLKoqJco+EBAoHOx+syiOUcpV6ARUR0H3
Ix+cHfa9Dh1zuid5ot4udOKyTuK2yqDwvz/E+fmpjDFCywlge1Mp46DAguQmOiqMCIzGJs+WdkTz
MgjCQmktYCneYMhjh62fiTXCEmILCA3yg7GXfJPyjIkFyX5ejJ/A4m3rNsMf7lyMoryVGCDCWurz
agQDRchSRRjDRxPk7uygkWq2IbnZqVOZ3CKW6ENTlVxGMlNHsVwwHzQ99L162jzmt2GCyX9rk6bw
lHOa6Gr8FacDNHWR3IJDj+L8Iw6hmq8PSeOl5p7HacXKJYe8IdWxh6/ycIG5qWtZsseKBoYrW9Qa
I2aVBJdTzz5YYLdbilvBqlnbhFXt3qfy5exTa86MBs99g6wCXFS8L9RM48q0kCQ66AIRsX+BebJX
rZukEbtCf3nD9HbTfj6E37UPmc7GPEQUTquSBfMCHwjLv06Hzx67RcMnRB7hn57EIP2LyfdpCoeq
6d4zbAQk+HlbmNt+e0o/596BL9Yvn4VmBNYD0wyZ6btNsEFhGxPC5RPHk4kvADGachZjA0hIoiT2
AfpKo2JwI/TP1d2Fv0xt18zx4UzfQ08SDMTfbfJXs6DmtwYu0kFfwYvB9mS6h8aTRokT13r2MBFA
Xn0YViVL2xaTUpEDNdv5xM6hLMGX9+RZElt64iZFHimmwIwOKcboWlKYBkGCwFZUaEac9NxoXwxr
InPWE7HoXa9fP03Nz8GgsITrNt0LhmKUJ7LcwAmOHjXX7E7ImvczoUEAZKQisUw+o5QqysX1f3sy
rh5B+gLTyOm4WrQWVz6ikPTcP5E42a6b3WoJz6+XsDmRNOPMfw3Jh2fkpfj8wOm5JETZXMhpqbwK
MoLv65GFkru/ILraNx60ZP6E+K6qthh79kXfEdL9PjvRXR3ZgXAGSYW1VMGDkyQYhuykK8N1M5Gl
TdxUBGSOwwLgfO8pxfVJenWRO3L3O2h1Gc7hncfyVCcSDK8JgvJ3R4w+zMAeUe6mD4z1sucPEXBu
dbfFjm6E3XPKNvGp6SSgfEjojDu7Mje9/Zh8Cu5kOVhSMgc263YzngScQfGwo6JLq5MvDmTKNPv3
SJPYpFtBbBY5EhLKYTsQf//QZ8b61JQx9g1cWrN/X8Nh+13in6SIEVrNl/HJLXJisI/HqvXdBaJA
Uo0eo/12NOd1Xl8KBtXHd+NU2CUvkoZC/G2RyHoacGyZHh2WTs2XnXw343dDz/1y9T0GnsTxGqb2
JDnJrcaJ2gH32WOSMj56P5Qw2QMRegMb+i+ewpizZpisuz0cHbkhFw21NJ/bosQLajx9/mZ/dbZP
VJmQik+bb8cLwXmVa35qDZMRSoTJjuQdJnHyLktzK8Z83hhSRnbdIZ25KMHNoPCWwybkVaOZTCgT
XyMtgq+lcTm6mdvuQRRSEu7tyGlwFwhA32vedl8zMbcqWn0dRRKPMEUPc92MHKf8ydygGvwz4wy1
noVmi9MFMtaZyW/ko5MDh2GJqOKy9Q3VBv25qL8VMWLyXaG7bhJ2mnDiaYJRJrcEDq6wqFvOGZOh
D8RT3M9wIAVJ991CTu45DFAf7/CcbhiW7qDdut3gqThmdWDSF7/Tpc1n7PZZ8cbmnqYR8UuaS+KX
s2gncXoZYwVspzJbMspgqZU/VYGvt1Dvq2ISlZDZrwoCMfq57/K0U6ZITxJCHpdWVvaKJivRNzZY
5zh3wg8MFBn8z1Aq/tPlQ/JOXPhHGkfmBA9VeETkWb+u4r/OB/U675DQjkjCMYpkSW+51UBnXMtd
GNPVT/nicy+h271rZtatWGtw4KjXiVWTHjeKXdQ6tYtlo2Hgn76ojccQK46dXRQXHm6j7ivRISvY
A0Jc9uRarpaXwJvwFkL+LQWVLTyPbO8Ji818UWDBiIQtL0x8cnR1Etqvh3BZKi+3eP03Eb5A6jMg
sairE18o11AjrdMCALoixh3iehGnhklm93JP3Nr4DoqtkOcx5FVab+Oiql5e8qOvXzhtKCF0TB9F
LhH7sImN7QfsaoZBDhThVC9EC6hd7kv2Z4V8YtxNdQPR5nSBpTwCruquq8QTGuWF8lxACO+Z3toc
5+Cisk91rjRRah4W9chi7G2csiBffJwVygu54lUKoTs3dXeA68CR8QOl5NjS4M+okJ7DAT8s4I0E
mkhlXExsmZHMEIibovuZJrnbBMVVdc212XTBpVfK0rsUKPgqQmjbO9p/5bA5k9nVX1lr0MDoFqGu
5hiNf6mqQ00ygP13Cg/wjMO3WSGdEYsZtAdJa4Sfp2Dy+8JfSP43yMTGR5xGjPmRbre9p8cqsAHd
cVUC+xsrKKH0naK03Bu1KdzIktvAnG7v2hywVPnyqewl1EI2ItQFnhX98cJybBPgo1FgEQLcSA6n
HywDj85vOt3eDkv6RXmv240YbczMgYuL8fD6TlOQoQULIoEvKMnTEB6qh/McUT+8Ez3IpJsDtYLB
iqUn2vadmNtCZb1xwnhp5pgK3EXXCv9GyfKGPWKFokeJUVCcT7Z9WGRciMrpNbgMtDXg4UrLq8Y6
cgJNqZmgZQ7ghwmGKe4CHjyiVnoQtMl+C2z3jlGpy8uIerUzD9V8vxkU/traQloqjRb3aAmEWkS7
2hqrmMmsqCp5S6dqz/AE3lIq6VO9ku5rlSbSLUa5gvRJiZ5z5o+GVLeahoo42tVjwZt+ZTxPfxME
cbvRFWHRn+5HtA2U+fMd8gXmvf84VC69A02Vp7okJ6ZRpIn26vBzpzBteC4iIdXhM5D2FZTl90+l
9e4mc6o+WDXl0R0Ox2Dg+P/sQlJC4Xm1fIOk4Cso1ACjoNgvFqjhukmM4XFSecvjg6saV/0DIFCD
6NAE0tcxirqNjotA17utaQmxT0tLugNqe5bKFRcL8v1SQ6CMKMo72lc/joaT+vzvATPD/VeW1nU8
GnHq+r86Z5QLKTF5TUFpFMqEBxdWfkME6W00ooCX+8RI0RV/CWbmYmFsMt/haN4JfiQFtat4Mo2m
6jdBOHa1vHaehAlUzIAdUEi49pOl4P6MyCtN94jHZkIrGmF1uIBCa4f/9Iq6YoC7DDTgA6nj7jF+
3wVJyHIqXrD2enU2XZHMTmgUwVKSdKPbS5Lb5L1klg/ZE0z46ENxHbsSXGfKnu/6p434nDdMCYac
O3GRvXd8cuIsMqX6jAXLvwC49gq3Y2ySY73fSUDPFwNe41CdOtorqE3iAfiG0wHrII46DD/pcL4T
dOtkckC+Gz6jsrObBBtKepEU9OTtyjqKZXPlfAYOv7vfcFEuj6oZpgXNanYnwyCcCBX1dIOgyWZI
oYmZg+sh3hfzBv64Syqih9VpGRpZVRQ9iAo4X0vNVR1/9LhMjbzmNlKY2mi/lXg1WyPO6mGFAzit
FqojzEP+EQ2wEbyIy9/tcv5op/1DB18pJPT7eq0v8bxf82BXeLfuwn6cUDVz9jo38HuiszwdAhyI
jB/T8VWraE2JTUhOfiu8++wTCnYekyj1R1levI4pO78SVaUVPSicUxeWhPxws9GO/6VHxSxwHO+P
90FIvHFBYYL82JRCWzZGGAfABUlo5LPiAYDfw1zmGVbwSkv0yqf0wa0wO9eN5tu8VmE3YI9f7IYD
vKp8TdYEaFzlDgjha/UsAjf5tWLP7XxhMUrfcCj42SscbqDYn+AMhRW0sjbYbR68Du0rOci6+Roj
cELegMIUC5JeGSvgvfQIjuqaVP6wUHwJrBZVv8njrczGgF1aLDHEdpCUKugft4giuW9t0L8PibTC
8joh5lty0UbgcTJwv2qu9UcUKjQeBO5k8LuuyAqyMgZJphEqOhiQZXrXWdzO0DGh8oTtMHGavCPm
gpeG9jXPVWhQ+UTw7r//so1zplt1NZSPiuDouyq3nlPNilu/p1iwJXXQyCqGn2CGkAjneMVWmQuU
hFfGi6rigdhzlp6DSThwY7UQFzL4Uo+FPq3FdsbIjx/7anhmo86Ph8Lq3OZcFOM5u8Rm8CeTeFhe
lgy7e99si2mfeIBYOrfGFVHcMNrY5FoTAft+vKZvEcmqcapTfH5XNMiCXbJgH1Be1eDHfAA4WvFn
tzhKUtD0g5KYh0ByTbmIVjNY9x53fLqCYFonkpdszQtjSLIgKAkpIVL65l2ItIIbB85fTHQOsyEo
12mApAop6CLcUEudJ43T7fY103HbKnSSClQYUPN4ZgluJqVqLFWrvjvxOk+VfxnN5/Ha+7u/vkT0
acERhmmLLlWGpgo2rFHIIGjB2WHwwxRuQ+3WVbUZHMAaRsrH72rkKSHefvbuN+/u9/c+YXotCudn
1wI4BH50lulDm0UiNoPRfjFa12/nPn0K8WhEUSnD4LWqZz5pm7qTQ6TYu2iiiLAJ3kfKaY+TJMAs
1ZlEaD30aWnpdtc80DwwIJCB1AwCSUn4ew2wxsfG7g4pNezryAPAwasJnxvTjpWezxYpU5Ni5xy2
5X9Rn475tpMCJYtK7urp9dDBtvxwUNloKNjgF2ZK4n0ZPBgV9zpi9UqiLa5CL5Hym7X1uhrysEC4
q8boYJYYwjEfUPd9MkKTi5e8BTczTQVaxCbolrUiynIXlXN4iNlZpHQbn4oBsEK8BOcC1lvEPFv7
nbGPjWsPC5ELBTLRT0jbfnUaAZEZhQznfB4q8EJfmw2gXB02OpJCgP6YWXKsOcWMK4hh/3sUj9/M
75y69/77Ivnbyy4m7Sakt/XHO18IBOAperteAsaRtGZG2RcNKXCTPl094SScYADnGjOSWCs2ClDk
4f4i7tbsNyD2FYHhALe6fyNm2MRLYDiY2NYCdz9QQAgMhYV4+PZ5haVbveAKtVzYTrE315tA82gv
Uy0w4X6sWv5weK0in80QLfmFccSrdv8D5sZJSzJedZRQHtGiu9JXdlXGuCyTTFTEhOPElAnp6r8a
ZPlf2PBcv5fJSh1UhhY1/zsNx6NkrOegFwnKtksaghaO7Ymi6diARKMuDa7KtYhChxi+Gl1ew5vL
my4WhI9pZPoppeQfwBK66MZ4i1nWEqenjxc2ayK5HyGrETMqaXUuKXm4YN6up33Pwp+BRCAdxOHn
ZeWjbFjzPNdw2thIpbS84h5rY7tTBQ1BvzmuWXQnLS+JZ7aEjAeRoKHHkvFjliWyoyBGL1ng4eXT
zlcyispZfou4W55Q13Z/3AKdsK5Hsxku0m6DkRsgISICmGyRAhh1mXS4mpxuMifmcl4VfZMSVWKT
TEPoKeKObW95E2G0QaWU6EooWDbRrDLebx8Zv/52RTm+aEad0eKtwI/JV7amgy8gOeMBS6Rvfxc2
Cq2lYKFye8JtPYNUPsM2L3PG/dl3eUuDd5s+9akU2JblIQ/6qwJTxxQg338pxZoTu9RPkUZKWrDJ
QecIGoXY+nOgLGhhngxKSKh30p+9CTt8ZVN2NWxkSIYSWs/MWEV0INhVEVPHe7VmTxSbnGXs6XaX
kGb149jcSw935e3fW589g3q9uH7XQcs1QkdjKZwc1VO4o/dtjQdMDXxEjXilw9Gu3Q6HIobeBWZ+
5BYZHhFcnT4x4UyZZzHNvcwHHDB52y1ZEAGZE1mhoSHR+1spRCsqvyaEuFaacX6lPLAYeZJle+K0
HRbwFJLMx2xI9U54jrK/muh4xA41lw1mEUs6zJKdK0H/f/FxDhY2TvcWcWpCkTSsc0P2ldAOHPEy
H9VMukRtmwPu2zg7gWMPOMacKb2HQng4yuXEG2vON7Dt+alB7mitBqKFsW4QNsuvNWQ8PYprBSzp
DoPHJtaM8/TbEOVXM7MtHJB2JAarCvDNAW54Jv4rusJCr38EP0Ok11eAGYJblMAXcpsHzYmTy5tU
3Hixf2+NhmUsPSzho9C5tJ9HTrIQ0HaKmz6o6iPN/MFHqSYag9wildPR4XajI3hLnytpnz2dDgOR
X434AVk2HHe9Y0fFB2Bcd2Cih23KROPVVNPQnO8dTDOAtEWP0k4nCnBdknfxkEdsmk63U3Ltw9SU
pE0/Nb9S8Y5N3MKzGuBWKHZYqRsstiD5Fd97n6R5cjXn2WEsAgrOxBR/2X2+xjVJQvPBVXPt8p7w
6rogzEgzJrtNGNvdxALlhIWIVaME68rUUbBqOEIsl1ApGhoj0cFmIdHPtSRYkxRrYuea3fISpw4k
cDQKiNBcpUAxoz54po+WLgf+XDJ9DVKD4G73pF9sM1n4Agt3/glK1eWCrWeXVDpySFhdfX3MJaC0
ByAGwx/X27nvVNwP42k4yUOumB/7tw3vQKdKvga2Ht/4tOH3zae+wiNkEA3JAzX+GTZBAOs9WyDG
uYtNuhdZ3B5BbMkx8bLRoZlU3tUKxzC6S/9lj57R6ekWRyw1apHu47SQbf5lK2WGCrjoJNqekG2f
pdzih7QSllzUIW+tfsSJ6kqPpqW3hoYbuADwGk2MxZ61BC1mYi/NMWCK8B7cUKGsbJefj9dIOkvQ
ik/X1AeP1+amvXHmgk7laxNdjiKoe6I3DkqVgfANfO3t0o3onQ6Cxw9+WCfnjmD1o/x6SvJox6Vs
1lv/WysHPGmKi0hWuQliY16p9TKrR/oQ37osYZOYY9Zdjkz3dvUTiAfqo+DKyIDYs14Uxv3TpY0e
5qnQjmixonVPzA63+OL8zQijSBOfxBWIuy+eikKgxYrXO0SR1eS9OoZKM2PiqBQVG1FP34viiBbN
dX2Y6plb5QDcQDWQuQIyX6rnEBHHZVeRski6MASGtLT7NXIUUXLALj5+16vo9rB6SUvD97tEqkx6
haAQRCnyA8AUhuxsQ77dnqwn93jU9rVvpbiFkG+WjUscvjbHBzjOlT1mQCsGBfuLM3e5q6akLlhf
1JCdD5ckhIBvQ9nTGiPf9UXIJEGGZABzl35Msn8qpAzw6CaYbIjm6ND1lXUv2kL+JKer8GAfFZ2I
AkrX0mr/wpFWmjK2kUCtGfk7nQY0IvN2DllytK8xhNE5CZmVtb1I3zIve59aY7rOp2CJGZ3DBpZc
LlU271iwJnMVxZDlNEx/WQdtlPh+gbNP6lU1MhDOg38Jz66iCfyn3XHrSp3/lamOkjPeuOSgpjLb
rp8h4F6rMBchDcR2UN8zQVJFRJ+YfmcKTS9qKFH7oykPYlCdYRnzim1Qf3+y9LyTDE8TKw0lEf2s
9DQixzRB8xo5gA4u7NRZ9XOiT/9inj+DDEic1jBxBwyyrToSeglWd4hCOZQ1CKwGl5Y1cAuIngNF
QpXfFX2h3R/SEnYvFRrgUcBgYE0FIumyXP95b+EroEgYX/B2ZyCxEfr1ks6eIr7c28BCdPBwfN32
2NI30uhbx4pUtfC0ADHOafh2DphYTCGkyzylQ1M/RTN1/wlHxcRniDNt48itl5gzXRpFW1/617R/
8BDTTj70JWRtP5PYgW/8zsTQOjnRHW1Ccg43eVG1vGq+D3gHOLarrb2avrECGepsm9IcxE6fmCq1
mufPhwhmZufrgxVXopIqypFgRJHeMKNbtrHXiVFz7GL/qvku1JwZSEDFPYhpMDuicynK5PmE3Sjw
PpuIevma84OXXaxpiV0xF9HMbYXyS3bEECV5cL/loKfOp+lT0W/Bf2A2hPhIhNCy1d23AqPKOb9h
RuZv6kHwalNf36RiohzjST05EOtGKc5D1f/sAJ2FV8UnzkP/eYsmuXycjFOG6pRmHVp5BeLhNddF
2YjQjrLjJyWT63mHFlPTbRGu+fEgSLH/S/kwaVNnMV+QuNruSfjnpknvHPXoU17LBrZwya4LiMpq
WNpzlGLbZq+ycurcLdJ0t9hl292v3ntU8iot/u5qpVJ1f5Kz1PVbr7Sezrk/8bCFeu91w7wuhgj3
1P5V/ml4PdKo6/m2mBi3VXCH+U/iLf69rOm8VHI9cRX/63+2QRc/oRQ5grggTuFTmYomG1w9Erw6
kkVzKNGIwcDLmVRMeI4FqV80dX7XmZChG3sOZbBCMXj2eTuixVBjkNWsvDIch/CHc/yUZmLzZCix
1GZKFOwu17+40A0ECTpC9Qtv16vcmh/iNg4LFzS6KzgZdJOjDTJCnhPzad7Gwj6AG2OnZ7r+lAug
3fQU8PXQwC3JD8TOzkbmACizDy5pJL9DsREtSifnlprVlgNrd46ac1gE7au04aVa9ZHqxFqPewlN
LMukHq517qEFVFsg/huxFlA7Cs93wMCxXAgbaJLM9nRBpBuEBk9tsyfo85TCmQOYJ1dzXQVJ9Jy4
dnbI5nQPQ0EO0VEIe8o2eyDuMgJBtApfLwDQ9d8ywFa1KZC9s/wID7aJWQcS7M4SGs0SCoCDLlfN
CBxyGPHW2XnLA0RULNIy1E5R5IyyFPpqJls9jJ2rp+3p0iOOXICdgEshN6MzvP5//RdWdJiCn6l6
v2T5cED69aQ2qmU85FCSs8Hc04VZySWELXeGBBfJryIU9NiaYcpiV19FdGeo2XEcjGPL86WZqo3f
TGPMfMr0fDY42fIVXjF93jKI7FyLJelMZGUaAsCpGzNIFasb0T+icMpGXW1yHSE5m7cYxegrdYOt
YfY8LdSGR7t/ywEcMmf74zFCdFFq2OsXnMhrRIiGUDrb7Tv3Ngw60nkmWg8nt9cV7Xq5kxFA8p2Y
EoC+yZNR2peD0AIwWZWSS+0wUVbozCzPZG+Z7UWoluRHfKs6vN6D74iRrRTyilIn9lAu0zAguWMz
gOQW+2kb03aMQtf0P4Qe4zFKAF1cQzDB563THqLovJJkEbivaFBiAvqi1FdQxNROyLeWQgyg3hho
4PNoJm4nH1P6WcvnQtOzFSMUPVeMvRbwu/o9GXTzSS3dul28gsrlL/j3u3wqGUSwj3lrpyI84g6S
qhY7CvUbNwBg6qp/wqMwRNM1KXHWVW8/+LpyC6GbX8TsI/3RwcFju24FDcldK8onqEmbW3+ubT2c
ssUPjE8B33bjETa295XXekmwD/ySyaa8LaJ3g7SKeIDCiGwmK4912ugMtkr86LRx2dTkAPyqESVh
iKGLFaP76UrWofiajjVPywaq9K1u5FmbQKRponFktwgYqBauEQT33Uez/ZNOekNibr5k/vCFWcu8
exNr95xMZPbnMWin34f6jIAFMP+KZbcy55XLWbFXf7kLRz+Vr3/svmMcM8HfZ9a3rL/F6vqQ4l1u
HaoRadUjiqhWbxs3A8VzbcbGkfAIT1VwKFXTFuV/rrAqil1HuM9tEZ7JvtwDg3qOOxZrameH340O
IF9UVvBAKPsMD3pI5zI+O81TE73xQmo+isOOuzMJVKteeZOKXl5W07SUkySGGgXEtMaU/1GNDUrE
U3OqQhu9LndeidXqFpYnbjiMHCSUGZznVBN2Qc0328VlGZTcy+O8SQmbeljKgpqWVHIhqixJ3Ymi
yuq3GF40bG5OVqImPnoauHibcUa40KDAtBzCgdolVs3SHcUNY+X5oWEyZ/OYbo3n7qcq58a5ICXI
/+rmy/1vl/uXeMCbZVSyXxVOFWrR5tKStlAvGR5Wfjw9lKaa1vGMNRrWvDTe5BpokPutBAmD6yaX
Yl0sIX/Hsvl6ZD3abvLmp8kW/F55YuNQ32WaCtjI/+465yjdyDXfgW9BEWpj3oJiIO9UP2fkrqRP
NI964KLHo2jDtICzkfZiwuclwL4no0bUJqAYIkQaate3XFqkues/jW6AH6YA6eGB2EADr0+4yEgE
2Rmvd29qPCJn+hyaB8HPfU2SKU4sOeNOKkYPIpv/LunblU1inEOiDPS4ZNSS+ACUA59VW/u6rSJ/
XC/UOv6OL8SXQgLm43NCQepIGYxPmeDFN9ii133NWkyfW+ooJCY+ejulu+h0FRo9/qsMvQEsJJo7
CLTmMFfNbk9KKEMJJGJPf8drW3NLFq2tP45R5e5dkBzfTMzaypkFCgvrtQOPQGbeycgYxOIBquyw
wib30ZkMUhnKAqzc4UnBqJY+SHPPTXJJVPeYpemFoYaUNpDCSXZU/0/sBWB3Z/aXSJKCw+9J3lrb
5G8Ot0NgPQ+1s9z2CpF+ta7QixNHPUThT5P4AeJPLxe1LgpXP9u2PxPo6sse2ec6c2gH1bXMxpPM
3RmMfqXi4RBliCM98InTCPSJZdDNXZ9R3H5g60T7k+DHjTKyb6cIDNC767AZTjRf02UiooaJss3N
o9iq891FViGZG31IucH1sAjBlBq8rRixGlDP6uPk/fWEK2+57K7muQ+zqsU6c2yp9yJ+IX7PJury
hxiudTHDTFOu7cvo7+/eoeXpe6WfWUaAW7k7T01DL9u3Ws30nHKiCD5vLbtCxQ94kbGNF3uA1MY4
6AIcqpEBLZIPok6y6dTTgqKPCGbdNww0P/TMU/9E35EwPPcheeAUMdwwWWEdW21lN4AfPeNapBIT
dYFVgP2/nvlwKaQMgGs+ZNMIVNDRcfHGNy5QFLZbUAVko2aqTznvpNYZoFcGFh4SqKCH/89wG25l
CHbKskmaT//IO7+mI4UTCR4QyK0x49bN8dz414Q+5fqIMuzlRCd/DDAUXUAZMCF0l0V/7tiM2poe
VRHLH7omnWraDGiyj//5UUFch5NcMwtfnpJbdy+l87VnUQCOVjMjLJrKopFoDAmZ1WDu7DVBRqG5
9djpwiN/lwsLmTm51vMrb69B7MpIziEPqL5U/u5FdhGrFf2Z2h3oO6FOLHbDgNX1GKHdpcIbuNDG
Fxby1CMYv7QgIcJLq3JSImzyeWLdv0ST0RMl2zV8fVfrgztXmYj9Dm1HbE/AbGUEhFK4UIde2w9D
5cBT0IfTwa9lfM4W/+9FPue9GEHaeuGP34pJBLjCgHS9FdFvx4agJK+sf7ybW+Ld3x53/8C0yLKe
aUEy+f7XWCISPwDsBL2zAD729MkdkYi+xD1W4G4hpgEuMDAB3c9OQvSag4w/VI9qaipcwc47Vm99
Hp/9VhWnMv593/9iogGbXTf69Z0onzCKWl/bOUmAHLIeS/+xZG1dNuJmjWF9a89D08gQwFCBPeN+
+/AJvJCF7DB+yfS2R+gkNrOvfBo7dg+B1QHj2Sv4/sE0HSEmAKOrc2Db3s+E+lmOj9iL1uH+YZLO
vvQD3ns3uvz4U3L31zqfn8sDR5cV1fckmkVt8uV7aJj3/yvl0Dw4CdJmC55J5HX0g5+Xd9WhvPA8
7/8uPZt9luMMNrTwqEvkLNTkA1fA0A35iVKIjro1irZKZ9mT/grkSlAeL9qqFena1pVWFNgqoVWB
TkzL2e5lRAw/iu0gzA2vlWzGjBLn7IYZhDW/Rj5wlaz3gji5lsHejmbuTDJC3NEG2miwdPA4Rv7I
4RWKW1qNe78xNQ+IUVnpLQu3QgEr+iCRCVH/OMFDQdkXz/dmM/Y6eiya9QfqNKvECldbuF0eE+x1
JvqUuS2lrkZzcbL0XZxF95vmA54hCqO5JWdzd83mUdCBNMLAKzJuadWq3tN0XfQhzsxPWTQeXXel
UHjsx11HAJAmesKCVN1b/OSRy0AnkohibFgQ54NW7XOX4wJZziCpg32OI6urQVQMnHPed+wZcdvo
cW9IpR2sNft5K7r3OrabQd+quZndbx5lYUcoX1Y4Hx/1jW0Fd1XQOzu/UOKbMpWoaSJszIFYRcll
bIAo+umLbCrNuNFjJQGnafSL2oxWbj+rz9gxMFGskw/gPbBu/m5kNCZOa2lbadqvRE9dgDd75mDW
eiDaIjlGoaoDEQRhPqT1gS6YfvmyLvn5Q1DtcMhN/86P7nMYQ+uEK2SBgIIzF+IijYg+xYstpOWm
rc5nA0l7aROR26DVWJawqoN5zZ8H9m+KtJmKu2UHnnq6QoGPdMZTShjDvtgae3gHKYOsIGwswWGW
5geDIomMBA4BEWDR9+vcT8B2RUr2k8lLjX81K/g6yZyxdFwPiOiezP/xnu5DqngnY+NqY40FY6L4
OgP6xs8ErCkIguORxjprczFGGRTKdYI5Gjvm84WBFT7kKoofksT1fBA3q2XgAC45mAgU8RHbPPGE
jnAz0WEFHVUL+feXevzDdO0DrGYVaPLZbFjybEzMvJLRuSb4NoWprBu00ETQbrUHiOKOLLOpjzQd
omXWx8CSDyd1Fx/dmOUcYCGO/Rq7khzifTRnth4dHmtVrSWK+96O+akyzIA/QVFf+/SjdSgDwSSi
po9ex893bUzqU1D2/wV2zC947azglmr0641rOEt4h/qYcavp2tvNbRLxN717Rdo27cQfICLDj+VO
2vQ3qJFqhYkTdPqwzqLPZYZiv7vAFWIoQWsl895Ok0hUtsCuF5FKd0WYlk4l4Xf4kKiKeONw0WdC
t+WRWuseLxWV8Sl/gURAG+4M9yzUYziq4iq011+ZMVBsY+F3DSCYtjj6yxTuLcvznM9QSVcKkNH/
AYk0CojMCWAMhg1tg0GXEiUC6FFcWwEGBDYzUKb98FtKekE59xjs7zsIvPhXQhpgZVKZpGAFspq2
Khgr8H9ll+qXUvPO6/3vhtY3AYiBsUJUct0g68z9fty0cSXdckTpzVy0h67fkAG99M4Ltuz8yjrf
wWfxf1lgywoKsRby1IjbiPEJAev7+aA/cA6/DhD15fDNefgeOahOxB8m/xS3IRgR6E/qL/1WX+1U
J2M85E5Ir7LamKFX4j9X+Ze63slffVSkUZK2UpfJxCN7VajNYoXNdo5BhqWygAwYCgD7lxAiSkQU
MAap2NH6pC7i7FHwjLxvBMYNZqH3Rr9t9BM8RZHsTBxG/ob96mdnKeLNR9BODzy2hLXero/DXZau
R0dUAk7eGPRGGwWU6AT71xRLUSdyJKPRy1aGwXNizLhwgl8LMMQT8j6OgUGqDkwybOZhhlWYdoVC
S8kzwHYDH/aDFdGbgtXpk+EirnO18JMalkk3ZNXT7hh8HNuq3H12WNtE7hqQOP7PSOA/QxKBPXnn
vp5HlD7obNpT9iSMIPfDQo01Q0vRq1TyaaHNy89yF5N/Mlcj5Q782zIgjIHi8oq4zYxlQYLUzSZB
EoJz+yMPjK3MLdq/xRBiQG/m+9R74oghUwcDGhTOIdbz/lKkaLXb7rnmAjbVeP/fWnrlSqEzoFAy
jYqDCe2rrMH7chLemOJua+M0kPEg9sHYcMQmoNZNHaJvbY5W+ldLHG02MjD04NudgjwJYQGEcAfK
OBR14CS1+M6/CoyxrGbQHAWTEt9skfLNAta5SV/4L1++Cpk7GtqeedF74BGdL9aBtvn8hhJrOIyN
cql+3bwd1RPOubksnKhULVznlfZIU8oG2JSr02xEd0OZ7RDi7dTM7DDaDecpVmtOX4SZYK8ji7OL
dd7NexQ/KsXwcNdW8EPyAyPapt2mD7zch2tGS8515/xOqIHP/KEhx1lfjuFwEc5FoOaGYzzLoPa0
4jR4GsG04sHDmPRIt+QYnV2MBPQbesWRKiFiEPPQ/BgN/H4hwvlLIky1JxS3YZmbvA5fuylMaicp
njCGd40Iwq1I2PbOA1RlBL6LCBuajLQJSXDj829uuvA1S4nfklukmkKZTVRm97RRLXyMGlYHSAGg
AsLcv+C9lN+xCQccI2zvYm8dv6VOHXz/ivK4GKeIeDqq6q2o4xjDspMEgQSG92Uhm4xf9icK9Rlm
RF7mWZOsE0hC/2XvxL7rv3YVMWwveqDeFXG9XLUdqEUj7xh9JWNaXGhvzR5YkSrT7XPW6Ol78ck8
L9i8TSwMW/l9a16eCYH0DiZ0Srqt5MmETyPSNj9mpAPUPXAP3/Vrfbrg+VgZPSTt/PN5u3/L9Lh0
swwcLSiRqR8nnrYqJd5WirpxJfDL53IO3MN47VaKhB7YUP1ygAE3H8LpGxFYYcaD2cF+sjuwP6C6
0oB5xy+f5JFl0hF77Qz31yyKV9tsRqPA2VO5/aWzoTR8rWr3AM3wUt5QGnpEvO3gyQSCP+cHkH4f
kU6lzw+dzMg86l8d4vgtQMadeKVoe0KkwJcvJwP5VLjSEvW2DMCgpFVXnzM32vQG7Nfi0e7mRcx/
1uMMzTG+YIpoGt5OHmq8NcJWF2gE0KUoXVTsncUJpafsMLrljxaJFSENxgp9yZ5oy6DR89Mfj6eJ
ilXuFiekDsEPmtToyEeJarLvGz5ZIzSPOwPyFJ0+jiPA8fSES9EAStwDjEe7VlvnWD6TCxc3NApZ
odrK8hB0SoJ39hcbKwAPJlU6MPh8Yh+B17RqcHsatOVwC2n9+0vEQM3hIqSHNlqT1frF317JEHjD
wdEXkgI+FyC7HYhDvnfxLlaXWcq1AqPFQojhFrgNK0J8YF7j3xvBNPU2iitgwtdHhvRPAp+aq6vM
KAg0z2kuTJkXhOLT9SiC1JLiguePJXC4LBa3PDhA8y/MjK4rr5SiILEJxFjjbjL6Q4hRCTWx59gz
pi8urOHspQos3yuKEZHH2eKRGpXCZv4DBXPK8usL0VudBef5miVwbfljQvb0vG3awE84noNhgBz7
EZ3VAUzmm3uTQ8bRx2ijwheurhDHrOTeghXAn8FKCLANTg+NhQgrFfA/YybsIHs7v8LNaLydvGbk
qaW1znOm8bzUuVLHZrszWIt3EDI1b5nIKI0MXQS+M8I8v7diAV42TmQlal9vA4qLDrg6tEW9aFmE
6hqN6l0qHL9qBSYkSgoyXz8ULhzcT7TrdcNiEvPhtM2uQNEW46T3dskCewC5MEHRa5BWo53gVvYE
SHjjgVaF9vsbOpfTjtmCECqteCTjEO6fOENWkIxvZFKPLCBOsPM+6QyG4FAPvDGhX4iZ8d/BOhMK
7g5kmrkxeqQKnI4TNQUNYMKWtSml0HuFBXARSeNhfMAgr+UPJetx7aH6zfHPZkU0TI6JJWos2NMx
Okq+VqI0/xucm73gieU8h5Gdr0BEVrOAyFJzIr6BczK7KCJDIiGUF8a5R2fl6h+o4C4TNYve2lIP
i2EBC2Yi4VZMWa0XMQJptvG4nxQuZb6Uq5D5q4hzBkCOMV6qzYMlQnd4Ux35Tw86rqM821WrfFs6
cTrv5SA7EI8q7nHkKu0CtOUNm0aVxY9pnzxwfiZIXIXmpeuYjpbT8hHlNeHsTw13+XJ8v7PW742C
U6x4v/OUW61GgcRJemKT8r/sJJLZdDJB6yLDfZ6hZLpHXh0QYKBoJBypSpwqEudImFhTkq/gZH0e
iMXRtbk5z7VmjtvU5ehQ2qbBjYlLK647ZsRLUeui6rCI3s0iUfhMG60QhwWlfi/IYLKl6++PXTn5
2/kbTX+f7EJM15H6rlIDMSNtIwqNi/TCaWMLkDo8Tor2QNs2kuhkrWkDBqKhpcjBF2V1vl8ey5rK
6DDEQTX4me1yh93CbiVyyj3nHABFiM1shcX91M5fja9Y0M95ruzUPeuPMoP2t/aERTXZdL0SmmEq
EKn2V5aZmwwo8PQnxIenUWbtory9bHtOsL/uQcfRfF2EV01MHIzO8qPep8l1pKoZZp96TtLwcKS3
C3ohSH8Fx+AwARKQGzJ5LDUVoMFnfQrKMLp9zOVxIuczinD+bbl+z4Jc7RTdqplnX57u8vocN8j/
hr6zWIQknyokPmUJCLZXl4zzTJjcE8K6x3tbA9GkzEBccqXYPOPOCgnBBnujABpSDKru8RjYpW9Y
ULDJzEay1Sp3SP2u4hgKO8hNAwtcL81wAqQ7ZsWgP4VZYwg4kFN7Nw6UmALJ2TS3mDKBdu9jQhXC
v1t2PMrdPt0lfmDLIUq26e3Y+7z5/wKwlDFQGqG47cuHTl53vzmFWojNe2SPjLvHhegM7Ewor2o5
lT5rOag0YCix4FdP3rSgtDI2DIFUuJrrQPZznROvfCTEAtNUTcdILnd00m7eXJ8a+WSES452SIL5
ajZ5rhu9Zb98RS4cIKBR/ZrRKuTukhVcEGon5ZGFFx0LNFjanp3ILXR6x+QufFZL4tGuei3PLK3L
LGnP1JoOXgiIb4i99Mj/0oFqnnWKlYHcHmD+JtlWPfEYmUoUXyLrVkWPlm6Ue8SE/YAyY4rVR9uY
HGgRhQF3HYZEdTvq+PtjYFV5Yphqyyv1sDdA5sY4YBkwLfytsazkqyq1h8yckHYKk0LmPKNU68aX
5Efdbgna4fwYU6MRMCkbud0FsxOiY2Wr+7/AISpfsNV2V5ANC9l0KuiMm9VJjEm2ncfIW3jhqi6V
km8Om6jrZH7y1N5pDNp9W6u9gbodp79U5dMHJAVWULZ5yQ90pzB88FkawurpBrLz6RQaP7CFVJUm
fzp+7001J4emtqUCPTkFOigwhD9/t9TKJX9viKT+NR5dA672mEL/QaUbIQmDPNEmX/13F1/HNkyB
mHXnBcMdAsd6sgnskeY1zaesY1b7NZLaSF0KSY2rulC8YYkS9WrSE8sIuyTxwUhD5nK5Utfp/mHI
MnPkejS6CvI6ZLNBLBnLUwojCvo8+At1A7BnrFkH90jcMEVUZ9GVlbc1/+si1CJCFc7XgE+OzFVU
BpQI/O2WAwJfo6IGfcENKR14gQozrQqR8LBickbmucnwNODsVE+oR1awyElKZnddLbYoR0MaSqbk
wcaUNTuYSGpkjakMYHgQ1qVL27g4O3UumjWqnzTnRA+IJU9R10Kh/GSeKIWQf7QzDzkya3kRgYys
bxTZZbpgHFzfo5unWc4wMaHCfu1//7IrJblgLUiJ5PRVNg81oEMH7ZUzWUNmALGUTOAkqX/KKN12
UN4EMVF4BxmZty6LeeT65WTTcSKv/XTnlyhQG6JRacNc6ujCeAYuQBTeJzT+vte8gC5/69nx1nTM
v3eg66srAE9oOGA3ImhC6YS6csw/mzeWKQDZcXlwEHGfU9nuO4wb1eQ1ZWy3xUFi1Zz45YAfDSf1
vhDaMBEJ5RbQSVThh7QEzxmCGQWW601R/GwZPkQ4Ttbg33OSXXS6KDytxQBjb7PIuEz2sDBMm/6L
Lt04lIUCuqRJcKlcjDezNywUh9XL2V0iQ34pb73S3qP8PlEk7w/sqMtwO56o+XjC3jcUsfkz0LcY
wFyulMCc6M55/sC02U6GHEJcOuZE1JVG06OyEFYx9+nj+0B3vsGuT+5zVz0dMeYjCmXH8fO8mlwt
1uT5LTYHPorvH3c/91BoOjYvaynvf5iSkqvZ3AG4h/ZKf4ygeJ4ZKU6tC7jvB41kiQQl0qcqoLr9
Ng/A5kiaewtJfQ1qoXHHsg8Mn7t80PGWKvwjtWwyvphkaaJFb4zBz5aWveCPEyNoCCBjaNBBNIyf
O3PRfZoitbUwBOd7VcevDccOF40UD93ZKvp2n6tFS55sMpRD4KePH8PEjhJMQmtyRepLk42ONYaD
x3e1I9ncR0zrGAiidMUTXff69QHmEnE9Af9XZZjC8qmuhLwCsmTTdcW7WahuHUGwtfoFuyf6PdZW
8xowbspX3UGesMFLPx+Z0JJTUqwdcjP61wsVja+Z5zBtMsPLwdl6OSOWXWouD1ryaHzoqeE+5yVS
JYIacu1p9Il5VocA3LRrwWj9C7HDjjepMWAJ/PSJbB6Ex5fDKe8GmwcY8/RHxIofUM6laK5pPVt2
lpB9xoreNZPjlGLB+L9JHRRojs5ZVLX3Yl43x7cri+o1Jj+sb0IoA1AliwPPumM7cBfGkMUyYV92
kzBIgIR8PRkDZ7+h06RM0HCKiSlfIUNpTYM1kXUBZbAwFxRDnksY+5mqIhHOeqsl2uDT2LQfs5JF
agxbp5/h1Sliu8TaiBerAVpYic5rlLEspLll85a3sjMbUgJnygYLlfIwu//nQwCEYXUqax6ynOVh
vf8SYS2T6zacgaCnR0df8vhmXaA+IW9NhmM4xgzdywXH9Rnhq+mjNaxgguWnoK64jC8AWkhJ21Zm
+byjTGqf4ftNkwvJOK+KCbrhwVBMHEcJLQHrZwzEEB1mLsAW7oqqypfnIILXSEG31ywDqvphSjZI
Nb6touHfoom6wScCGvA7OPKUapSuaBlsKc7BUUJXigbJg2jCdUIV0dkbXnrA1inwtvtuTy5pWUbR
uwJzCHexjZGt25skrglPIe542ZI/bmHw1CF268gXBRZjTp15bIHKC2LvUBUELICU8To72wIiEo0T
ZsHzxuwQ3ZF6MkY0fSBJistXfSte1YbDDKqqnJrmcnPaAkcxa3i/qlQ0gIhObgCkif7yI/cL1Qcj
+Yvmxt/ovW2E9wDok+aqBTm8y2u2QQx7W7uC/KFi3GJ44eZRF+ZO0RPaW1fjQAz+gIYi1dmyK0tu
MPv+JQXC3Dj1N66Xu5+Z7PotE9zBCqhr9g6levuqC4WzC92QJ/HOmBQchr0f+QlkaDaZIi8ZwIti
nVc0hv7m1FAYaAYenmyCjXOJEkeSeoH1vHu32+PkW89M/RKoseR3PGnN2u+BET56jc/wz4qGd4wY
U8x1PIaSl8t4t+2rdHHIJTUmOPED8wYS/XIHdiO9x8L3cvO+pUf1KpFrylq1/xU9V706HvC3CX7f
kleQEMVlVpKntREklZdfvNmokjGYt8Clz12WunIuEMTgCxG3APcZ8zr1TkHmKv9nh7eahQEurLsa
eg5BXZx7oPTMEQ/heKOclLs/RgK+b2vmDZEapsxwLF+Uev4JUk32wQb/bWdwnCB9UXcxl23Ygq1x
3KhX64+Rri8sHIG4iYOSBXre2funbkpUk27V9OeNdp7mgCloUxuoPnPBf1PgShSGnW3f46vQP86W
m76+3bUQmQznLw2sGyGmOJpVyI21eHRWtQo95oCl5tPwD8cApXn1ta7ShJWwGMAbh/JjnD74ceeh
39pfm4OvC38tu8eF9ThMxLetHJxRtl+XyC7MmTEB1qZ80MK3c3DaWf2u2CgQGQmbOiINGWdGsr9N
+yKrmycOVl/jAyb9VsxqwWVeE6RLztoPLQPvIBpxbJzTyqSJlOx0RZsATzxQXE05tCwTQ4c6fxvI
niPJNtzmZtglFFV+Yl5shiL+7ZvmfDra5bQkMNvGaMTcUiCzzep9B5x0KwP5oFkGvU/UOG5BvS1f
GK/KMewUjN/dKLBwkwwe0DiqM5Xgw13UdG6LpwpWo4JA1C592iEmx9hJCRP89P9Z4g45OHif8xz7
K1Vzu+0EuB5wYJQtkdYvtG0O1T26yz1+fo1Ltr8nQ6ndkaeijOZyIJ198+RJNsAKOzAFRxBMdL0j
7C+fqvNOYGYSW0B3XRM1BXHezI3ahxGjuj29cAW3364mVryBpG/jSwnzf8PQWN3BfsGuOyXkBhst
FQlBuiaUzAqC6xdcBx2Rdof2NAVTgPb5y8XZY0X7iOSfQMPhwFRnmu05pRdO/tZL9sNTKdV1LQt8
C+pxkCL4bo8JsGuKJBQ/iVWR6To8GN7Vgqh7HFr/XTcyGVQMQwg/HTLMW/dc9ypQ/6sGzmERmtyL
yq+ORofSabPjSp/J6zGroqOKPzrpZRTM+QB3CFvu4SqGpL7ZLpbQDZRsnkRBmuaxfptOykVXFjWu
GA8QPDfp2/9coGOo17j7pal273R+95U8Ff5awNCZe19Cd9IZ3UuT0Uq7YKKvlg4GdM+LMUL5qRfu
PyNdu592ELX/v09sHxLa69UWt0MmSgPdM5ihQHbfbVvc+dJax0Qe1BCbyKru+6VZSBXYa6IyEPwG
8hUcqSeLzBaW8Lw9zkP7hucvEac5upqEr5NZdjR/jrSY+Q7fRdVmlPxCUwVRBTbQ4zGyZEZ0H/Eg
1IdYLsm2l3wzk3Nj0HctTbtVmnTsoFKwSvS96DYWLgIDsdCPptjSMgxmJRKqTGZFgDD5pIoC564I
P3AgilckBOo7GVTQg1AQQF8PBrr7usWdA6k3F3dqdw4LoV+p/kv2LJKa3sqGmXXH7AyJwePUv2Ha
Gf04RAWdYG6o+O0VTYn+Zb+xsM7Y8+IQq58KAgVJa27HXhNDnWvmMdWt7iLjkjwLILAQPFCv4yYS
+c7cvvOx1nryIDHnJVfKNeuDj7nzH7ziazXtAwnJEqqIK1c7Ykd6OUxvq8paRdYVw/IMssUthhrV
kJPWXYARHzv3f9IKIjbVkHOp7Ebx3DYgmo7DleQbrb1acus6noRQfgQXBSbOSBnyO4vqVMmdu2Ic
60pS/dawsigGjyh6laVK434gHiAWsuwbSDm9qO3H9Ma6WMZZ1/1UUrV6r82KeeLOO0dBgOUcpXJD
rUIDJIQdhfZOzklyok59kkF0Nr6rVLYq3C31xC+Lpky2xezauCs0tKAuuNAMj1KZ2cn+1miRSbmc
HxSMn3o1QBY0ZEr4zAOXWv4l4z1X2L0K+iQz9q9jvo/VVCzGJo1FYNS1Th8h/ZWTw+0vpMHTP9LZ
2yqqZm64pUCYwk88yeWuLUlDbKxqEtsKQbFS+PGT2trLoLKyaUSUgGb+BqcuzyO7KOz6ZMvAE52O
f/jEZaSNRW+pCYbVNWDwPbdkAEq04G4Qxhp2I2Ue12cl789/uS1onq7q7LkKatQmnFigySFHBJtj
Dfo5wAqNCQEQwgOaS4CZT6GzZ05l+DJxG9J/TpuyKvNCpUxr3UqV5m7gpIpCHyNZky5r/1gtVciN
PnLgS6eO4bOQiFYxvMED4BJU8QuUwdZDPrXiVTDDrQeFxhe2uVjpBLu0pr9rSJJslJSeEezRjN3n
BTpOduLTZJlgy9wPQnfMY29Is2UVo5aTZYsxQemWYA2sAnygu3TZsC++BT19KNV/o1xwkCM9nFQW
iStwUBxn1kjsjEJSh3GI/06LzCZ0f2h4SLUg8MVn8XlvGRrl3q5qraP++9hkPg9xmQLIPtyOap8+
+QV5ypKJknKtc5ykPJqfV3DCxjlT0Cvc0Pht5JMdfZXO51S6RCFdFGBv2HukUeHqcwp+y2j46Wal
ZzgN6MitEJ8ZTOyvVzdmvY4H1NiqpNnx8wIBOKFKWf3TyOvgSJrVopj+dglsWOn9ONksJMmGkeyw
CysxTAvObBGBQyy7RvhYgsj7gG8yJC56gbdK7uKIuAbxCo2kuACYi8g5C8fec3HAjnRsP4fwoOHD
Oga2gsKLz0+gc30hLC6ahsr4vKjmJ7yrFI9xEiJ7W+xRdVbs0fDTSLEidtZEfW3KCYpG5IBlNC1A
xv/OK2Wst2MHxNuOLZHIptxm60Em/d2iDqyrHCL5jFnr+KDF5RZc5pGa4g0CTNt3RIBFLCg5KRm2
9Sy9kIGqKBrSXPxNRsX+k+kYDi/gmQTkmlIatNh8SmqdKBpQoe7NAZ9ntCEHZ4J+1QyVleXyBbOF
0KvvPDGLRM7Uki1kO2xF7LBQrG9IiZSAjiYLmd43d05OvQYkSS0bFnQnEkeb66cQUfJ27f8rSWKl
1IndEVriCzzFfFgkvGF1LtH7DpVI/AOEMt/P1yp6MMzsdBu/Zlw2qcAxJBRRQYbhCG8KG38pxKR5
7n44hYmEHMR9SFD1OADnrCWmhpoAfn+iY+5eOZk+w9nUUEp902E5V46UXrVGjavl3AE5wsiT3ZkK
5P4mqPW/nrS0J7ZZ27NoTqt72OFk5F/uS7qJYZm+sE5RvXU6CRKkUx8Z+bf/D14m5jtpFmInbkc3
3dQPdagCPer18d5oq14p/yMz/oWepZyiqlSyQ8sUCudcNeNC5Jth1JtdW5QdvEH5xHKlpVbZuH/S
jVYBNISio8JPYJ8kcOV5M5F38JKFFR+dbxo+nQQqsaluuC8RSjmq8MnUGmkZxSEuEIlOuWxIXV8C
uUR8LBeYKo/3JfI0Lhlo/FZQ1llwyHUBX7FXLb/pfyxtA4d44g/Xk4BZgj8mbpdURn7Np5+n7ERc
5m3vdpzqJjV04zMWPWRKZylOQkiQmdRN7o1j2T5U/cbBcS+nXCc8DfIdYPeBM3z8DmdceBk3BAuS
+EviDaUwWLjtd2SWt016+DT9hBFI1vXgCQRteYV8rMKYzmh3hFpS6+S1eph7/QDpoz9g3kHGz+wr
UIYNnJpiTkdzSfR24o1JpVg8tqWz7t1Dmw7Ff0ApbqofUeNpPHNCMi/jd45M3iTr65gi2K64aRg8
0IIKeR9KP/YbJNZF21T9RQNGJVxBT9/8bF0XWG2Zz1/I7SeQFjMyRN0Hz9tZMBFGloEaNxwvhjtx
aQ9JgXEyVya2YOgh4x822X7i8hBzqZEkmc48wRJsc4lgGPhZBJMOmDh8BrLn51COORL//YCuhTdg
j2iUc9YqykaQN+g/oM94sydx/uXqpwdyRW4fBEm5NYq1MK6ZdJcGjZAzoRVgvViPdnz39wYbtatZ
8V3CCIFUGk7t0bYeZRrSIVMpRknzfOOgNkW3s3mmM1PcYXL7YLk1nCISN3hPev0ydSacI4o73PeX
gpTUsKU8scc2J1s7fAh0UmjM4c3GzO9dRGL76lxtX+TRWq5mBx5S8KabgoN5nGjAOJbpI4shyfMZ
usjAKwpxaqsX6ux6Own9AA0XN/yw72f6Plk5fC19CGlWCZfF5Mn9+kDw1rdTPtT25muPIGrjYgMj
bGpagtMSySC3oC5PQ26+YCGFowdg0yIPgnR4dkFtfpujExGtk9hLewNp5wwRuhFq70t8EV/dJU8n
VdilnXsau7rWSNz23A8ASgKM4rS+yKgZc7yDJVIbHpMiF/wDdH2I3gWXShd4N5uzdkAi12uY/xnT
qRD4GWuXdotiLvkn2MuRsqbH89WgkulDXOKtDk+j1UIkIPyyTswbxR8L09T2TjXBoByAUYvTTEEf
eqejZv/Taa6ePpT9UYxAymirA/nGwKYCRc/w4ltd+ZSXeaJF5i319+zLipea+HP/DAbzKqPCqseW
7m2OEzpKMycgOfmgR582+JmyJYMgRpkXyatuAD2atf/lNJ/u9fjiQUQdAc/bseTz0mtMZfTA8YP+
tZEAiwhZx64ufFASteRf/5MLSx8O1ZrB+d3icr9p41VEeLVy57bMFkhuz7DvWDFeDSe+jHsBg0zO
Pmed8zxpHzcXJzuJ0fXCjv6NI97o6PPkjVGWkIvwRNDibNxyJVrzid+1XiMkXBDYeClPfR8q9HkU
67QixwdMwAKuwimIDHQKI7GlYjII0383K/YGIXsopdfN+466n0NQxpiNXpHY+gVrUtEFXK5Z+AFA
6zdK8qSBnzH/sB0w7bh4yWc6J5sczPR07w5t9OgAVcRbWFTOTi/TUkH71tM+Vqpiexyt9Mo1RSC5
ySBmwhYkIMenqy1sHWeNcZdJ/4dUF0FUkRRY+AUYugtoFTtsTUFKy5szaUj8jmV+RynRZejrbJnH
tQU1KBuv1AGMPYNqtVwOUpq28RUvzAezskqq5We8IYbrXc/tfHj3vFprrJDPiv5dlfhhwmKaHPOk
0H5Qyr3dmlWLn63MDbiY90IdIG9qkZAp+Y3c4hcunHM/Rzvr+Y9rEiFUrB/AB8p/UmEVxjC40r1w
2aK3ukOYp8e7iqPF2b0rOcWUbzban9DentKOiUZJ9zGNjDu0ccv9RMUxpIUi0GMM1jLtB7lmJGnI
1NnQwtIEgG4t/wKeiYO/BWtofHPEE9I9C5q/stJ0MzV8qbfANmjFUoMHtWy142D8b0CNxNz2vdis
8VEh9Q/wubxXPpoGjbnM2AMO5x+35jnGhJ/nj3mkD5ITuZBL0ZMTT76nsH9fpn42cn/ymyHp9+er
RIT6BjbNes9OTFiKokTTPpIBs8g3+ec5y94lHdDC8P4uRSUbOVZiHbV5N6hOdyIgV/4wMOMA3Oly
k1jiCYwJdBxT64ANXKvD3qLW34lDXhfiX3Fp3/7gXTYzYJ5wxestQzKbRA6TYwVWXLvNnhe6XvMg
cgaa2dRf0wDQWaZQhmITXGgzFIaXGQg2VewmosVKMJVE2/07xyRplPArGp2cPu/L7U/fNrON3qp5
uPUXOo1/qxzbnpB3dcljg6WpvvkwDkDzWVA6iXJOMT76gUHsgOQD06nXmp0WXpgESsQfc2VLRmwd
1IqL1iAbw8iMSOzokCUYb3dtMlXOKBV0QwxEDoU7MlQ/VGwWBSuX7AzDm6NgaHyvniChqvEQxZWa
MRNyhYwtoelkTIugGkDoj5siD0zTzYDWtVosMGORd06Vb4GIv1v0/5aI+DAQuSW9zK31pCDj5hex
LA0QNCLMV1yyE6Hl/bJPLY4ud1WsgUwFCYb+DefotuwUokX2LPafD3w5txFQnNWS36ZcbO85ufoV
9XPV+6KaK9O919fVSk0LtyvUAQKHDmkpCzeu3LNKurl3+PQklVTr113wZiBQVphc0Fdud8Oqj0lO
FOtzanxeuaVldjE420qS/1K6e9RsJu6Y/QyTuBCau3nYvkMVAWerJvWRDFL49msNqpZQlriuyAIQ
p7eWijeQRTmGcg5nCe3zwXHo9oU1DQ2AaadZfoP0XPXVeDXOxz2QUYlFVaoMAbDkn0TfQ16pn6eL
hGb16qw0pCbLR0h7l1VuTS8SQHkDQ08cdREeAL1kjzBaM3b8OYdUrzuX4gZNnTfZ21MwMObKftPn
5uxq8rMTSmFwG69a+kt+4hDc5IBMgLpdTHZ5WoLwG5ecXLjPKI3B7F0vdvOpGrFhJKPF5eRDAHAl
dxtPBWL6SgNPPmnTEIAA7FKj+j9zv+uKqxU4smvCzMqlevfPlWyxREjcZVEZukTIYq9Xp3kt3XJi
xbc1f8LpQO6FxTYQEA2teFYFoWC7EKM4sMTaxe/WN7sFQxxF/oLlkYZC+sEtm265RAWXysOA8QU/
7I4gLkyfQtULXPd51cjuvoZ9Q0/aGuHks5jxgiOQIzsoUwOAwGPe6N+rKVckP/90ce70KjMkLfMw
GhThJ9mQ71WPylo0qHykQmwefY6fMjKgPTlIgItnLCIUKRwoSqPoxSdRvewe/IZbQMayDVIf1zZo
m8izspsXuhgcx915/pgYaGZucs4uZVYGRrSHnWLvL3JvJAsUml1gOvZCjuVFn9Ywj0wyshfs9vK8
hNIjcTX4w4xqyWUDVFYJMsZ9s7arFU6THY3CibXp9LFbylMoxpkCmPBvqrjXHEE4zQM0nwMLiAYd
M57q7fhubzZCWf8umdReqV1FV8DfzxvPghwyO6H/Wg4wF4wX41JtqrhH+9dRkzJxSRvXH/a6ASE6
m2g0b17DZ/H5Etp2xQt7CEJ/s5KA4oxIXLXjoQ6rKDyvj+tmj2dM39jbJeKF9eQL2MiFU0U7hv2f
hyud8GEbnObHajBYpkMkKKH+HL2iSk83SO88zbQH1X9wgZOjmDWMmCLG+DCGoHHmVv/AvWIvDNUR
k3/0auY/cKIeq99TeOjJqliHW94/P91Oqzb0/ta68DIKxMSdzg7/U2ZhyUEz1Sgp0WaygNYghxTt
ezMMjPKg/rsU69sh80ohkX4SLfksr84QlqcOxdrX491GvP8SXPepn/6Bft8oo5UQ1USU+CaoE7iw
d5sE+/22BJyGJGWBlMPThK/MCKKuasKzWphcN6+EyAbDGWSyAxFSGv4r01CD0F97nHxZPlBnYCBh
8F4fUlaD8+FR9+wtfneitzJQIEswhtA0LAOMRgiM09eGdFBTXDFdP1ByrfbNzJMXVzZMvlLqdoON
+XJioHNMXx+vmJuuO2v/PcHq8GWV2KyjHLU2BrW9b7IkjaoA145DgP3ZMYVrbrj5V5R6mYh8XDnV
KX+wbONDScQHwzI2uhc0WlsZcF6OOX75YtsvFRGqpN/bT4B4+pYQZU6F4yh3D/AfBJ8M73F/z9eN
nn8mLbsKyb57wPjg/XEHGwpqYUBXCp8b1LK5Ywu/NLa1gb752NETN2n0pKlAVw9gqoOu79TTuV70
9wtoCFHOP/6h9McYuKOGemdcuX2TMU0xHHEIjlXgRtHUkE3FI+NRFUR+REGOIpaXuV7aKOoT2N2U
aKjIF82tUnIlYSik8bf3iJ2UDlKKr2BKc/CEEOc9Br8Ey0zK3I0dk5ITjimE+PKDGgS+20QMFGUE
0KPSbXGDYGPenYpF3GbVCZQvbGm3reSOfhG6WAn4xPTipPXaREOeaCy22yd407PL68nhz02eTrg4
mcw3pJJFKcIJz9COuDLJjfqOVDWGwBOcsKvz83NJ6r4YKJlucHV+tvOeEwWNJ25B/39UsX7l9Ehq
qNKEHs3YVfTiJvws+ej9uORRW7nxnCVpxKrLGFBu8ss5ZzpPAmct0qn3rYuZQ8YPE7vNQmYk+VZb
6uUIgec1o2ZxZX1ULyWQAYGf0EheJenFH0b2RJtH6s0eFJEYqMv3Lk7Pp1HKRZcZNC7KtR7xTyGQ
DzdrRDL5PbTnYl587kjciOYNpllue6GhnqfCicBcJirKvZ/aHnQTJ3B/0nBbLd0IDqB40u/xMHUQ
HEhWUXPXuzCcs622GUz7aROWUEBoKYAoS4M5JQx/ZcVisv5YhNkFiBR5Vjd99QhZztU716dqPUoO
/M9qV1Hbm008W4WtfeWzrXmIOaA70bZ8CRLjf9B9Vj0Dx91vEyCRVoO0HAGs8GdD77bsHGCF2RUH
Rf1hd6tgsZJzdc4aSQlI+7SedMP/uUoi2Q0KQn8B5ubkYLlRPE1g2nRJjg23f62bLFsumL6mVgNt
zaXR0uSIv1bXR9KvfTy8jbNS+2R2jVkcv3SHCp+y3XW9RRw+Dwg90WsWCkv4F+bs15EioWI2SPFR
fN4Q1ZAvMtH7O0XAjKbZ33ZfdSf1OfP+sbPYupCViVp3eYEm8hq303wtf/zIwR7dEj12zmfFy8TU
twWGlk5Sm5bGCMVdTmpPJeJGTaPdHZ+y2Kn18qdgjuCUtqs174iDpPDPEhy93Ca16+yzQE5WkciX
rAzvZ0KqOtEvJbMV/O9ZSdfruePuRz5k3/3o094Hjs4qbBnRAkvajPCWxZtsPikF3OxyFu7ppEVw
sFn2GpmBcxLtduEML9hP0vZi0LuSLEZ9LJf67cL86Pty6kCklqtmuWYVtnKXmHHxJiDOfzSrb0Mv
+QPiRL6ho4nKJ/IToEXOAma8b2t2BCWFHzef62lOzxN7u+r6TZ6ZNi7aLSsZdbCWnBndHRJcmLKX
rNRkLOJwKaW4zl13vzRDKFvEdwIbcbZTgOdM4AV9i40pY3fgPr/75QIxGPDU1fp/XvXB9UR1Gn+6
cveOjfyvXxSrvSOpq6GcnXMGtIFpQtbPO94AThtpPoqGRao0j+o9bSVJN4oO+vmXkWPU68fSVlZg
ipXt/GdrMg46q2C8/gBUnpPQgFgzhapPU20ERXjjaY6k972Uynh9BXnwFCaHWGfBPQml5wYvdtWv
JV9cXjhrA/gS5lOOh+3iJytIR9Pg2nIuuPg/Qew5D00oDqX6PpTJGfYQMbcfWqhx3L4PbCplur/S
bP3TARCNgv/uOxiIot+mFbaZsG9ii0FJQwXUL9c8QJOgebb3OxluGvyEjpeYP/6aF7MEJ1jNTf6M
VAb+Xiy5peSX3ZokrYZCb2t1dVGBU9bcHhoEXPdigSt77L3oAIopK2r/efaiM660/psFvrQyUBy8
KJEfuGRvhlJuKBAi2C5nmbKfKfkLVrTu/PntfA+Ge2dnVIR5DATcB35DHrFO83gaefQ6BTFhyUUW
oGlriwtH8Nrol8oNA4yaGufh8YTzERnWJ6JdLurgwR84P2j4Feddpi52Ih+Yzy4AVrJh7MxwbJZl
0dER40ZANC9jQ2OOo5GVp9WV9j0xfx5H2vV/wKlAblPeBPUlSCSppQ14br1H/Zb0uc+bP1nMSSyF
aSDt3d0ajQ3zUJjRMT1cQC2MtaIubmrw5kfG8GMocwCPFTo9muIIdfSwardFwQq5n6nKKfJlQaAY
pLESdWc6QbN558y243bnlMu6a6hE/8a0eBnyZBJs6rY5yj4v+P2yRiMHozIlGdGnXop4MTiumlQp
4XCGFjB1LQ1F7L5Xyx+5g/CPOn4GcCNOqFtG0KisWAJQ5z1X8tTl1v7F3ub6SbufZDSI0mNjYF6I
omvOYCsDtB93v4pgBuNzBayApd04ChQmxhw0jI7Z4cBjvRS5DopHo1m+euzPDZvM4mxN/5L58qnx
3qStNxbw62H9ZJxoR7v3cdDEPmqe8Qso/2zxN75IqsKvHaC63qn6efplEzVtGrZRcwqO5HjLoT/C
1185LMvuU2ERJxZfH19yAiAt7GB3jnaU3W525O6QsTvGmRr5osIL3JVTihs0yIUX8dWojrELycW1
cSNzn426nbr2lK94DBF4JS0U/KiDGzd7c28J+nSW7XmjpE49Qcrd+wqspoYaiUqz0mR+ixuNIapI
Jb1QbZHuR32Oisg5sImH7CFCOG+dBElBWdZxrhyzEUi/jxcQ84UJqx/d2+qqDj51Q/dR80U84GW4
/r1wjg0heU37K/lDDuLraWt+igYMLvmPB46pDQas1zXjJbAxh0FdcIzoeg6hdkk14jMICNKognK7
LAa2sUkiZYmV2Va6a6QkOSgR9lUgZmVG9+5pPsYQ4ns0TWIUS4hXraR10ePphmPnog6zkR0oPEVU
IvV26Gy9XCMuy/XWJrftCeQKkN+cNFc/hZh2932bw0aMgbmMBsDR7tEUaae91FSMlfj0IONpC7np
dYEngXo3OETziIwYsZrJrZY4jMcsgNdaoZfAS/sj9Cg/OnlzEq9osdcZ2/MpsWwtDs931irbPqBh
IAL2Zvp9NSNsUSWvJLyFWbpnWjbNgDoZfRMAFSSitgwmTqS93JmKe+zlqdrfKY7YQPLfvjRjBJTa
BvsPOVU8u3gqlvmDzlFAVzDawxLN+WKWWD8IMcqI1D3mOXzrGlZgTTmeX+mL/JuVqvdDWYeSFZ2l
Z71UzB+cczJTSvdZx/ji16F52zbBODHBWUvlaQJauWHKo0kVqOq17+fUnz7vwOLt8Q79TuYSaN9I
jc8fnZbZA0NJdHv6HqwBoM+r8aT/KJlYV706qw8rUcP9U+tqt1u5ILom9DyI5xsxHyUboi9JsV47
flmqUNqokez7/IfdaLFZbDgydhtd3/QHJ0VopvTuOzzcBWDTEvb86DCGA3tJXcqzrYdgLj/4/4o9
ZF3Vm6okkWlTiX1L3vdvKQ0j+vKYHMVfnRHYmmIRHYhJxMZxbvcDRuQ4aLzw4xHzZc9MaafgF+47
wuHtvSyjSaDx6zPMCS4kM5fOLelQEAEO9oP8OmTp53DiLDO4mit2leyIsPVj5TnUV0JBhRay5k5+
u0xLoKVybE2Fasnvjj7tjx1OqV8Bopju+a2053JAP/maKBEgBKWjKCIqwYm+lanQrANm3l4AqLvJ
Q517XLrg0GNW02rlb/YLmNrt5QWSg5U8PzttDO2hpRYLbAN+QMtxXgOU+j7a4P/nZrffzvyyIl8Q
IPGSzMJRHWpLrIMMSvtbvKeFItH9/RTTs2GIk/B5OvR8FFbD28q/HbbdY/P4yB/I2d8deWNcqN4V
gIly/K07znjdIKRHXWiYoHQnIidR96mJoRX4s1r0jJttBaeT1Pxjwis3ThBTt91iEg5oSoKdwGM3
84tiEJxsg28YlWBGElTnz6BNyRMRHaMj0tyJ9N5ICtA7TcyGcvZsm0BzG7iiwaDsvRP2+W3KxZ3Y
wtSRE9ol3o6f083WFYXOcsVo/4OeL4+euD9qLNRuN7icMRBLmJklOZUQwHttkEGqDIM8/EWA1jDo
s/yCq/0QrR7lFJcxTIaHbAip79nYsqeCnVf+J1fsH1BzCWpomZgPu/E3VO/T+JjlYkpsbCqQrcNl
YVAK7Alr/hyn/ElDpD/PRJ/8qppCZgMeO4qC1MagS3gl3V/tuiSI2GwsnEvevGkpMGxehKrFRtCu
7+HpnBM2kcHyDFU5fWp5whtxreH4rzsQHpklQxS1zePukpk+y1yo0DJ1e6PvSWceN6AVdDXiZ7Pz
xbs7rnUytQVkEAZT/jCjlYUemUkyHzbTFFBHvMlLLNcXNK0qXnMfOy9NRzXWH8yGl/MENsv3+La0
S8+xV53fnqdsAi8RU/ngRRRWWtw9pXpJ3J2KHfrSlgIKYvzvaGJJBZQpUYu/kxzWQ+6Ga0ffgGnH
VGHhqCAE7IOZrWRAjlJ2lb/o3VeNLPPrtItvZ0z0jvdudFfmshuig0xNMjRCDmZ2JUM7hStVq1yJ
SHIfUwnZkEbWsJfHlZOG+T42B6Zn/hdBd5V7VQYSQLw6tLXZh5maUTtXVXCzBdDPfwWoQkSTDIp8
iNjcavLnQc7YM8ZLd3j91J571eI2gfHs0yfOBLoleL5t2FHkpLebvnLg/UzYM34Qxgr+szLMEx2R
9ujEp2bp2gFdBz2ZpfUNauMxvoiPBaVclMVrtsX2nbOq0G3EqNHmC8J/y8chK5ObHtZ5E4ToK772
gGuY/X7qZd7XEfdDJeu6oPWAA1YagehPGDDGfTqUxSqohK/QuVjN0iUqV1MROpEaEJg58Fb7FbKZ
NJ0NSjUwAxM8kWCCkocuz2wU+dR+d2hxtzJ+F6tR2YjDMlQ56RzA3kHCP1QM+46VxdT7sUGxzTIm
AFpJh4F46yQkmYo6HwsZha6wtvtGVi1DM9MYHvEFxFnDDeabVElzyA9OWANRw/eoMkevKN48ltBq
416qPhq+U4w+dK1Oh+i/eyiQPFakVdhZf/05b9et3Dm5zDX8gFhaECsBPsDNuldj/279ZAbRJ3KJ
4qBObQG2ayiW+yq2L1brWMjuF4ZxfblG4ubDHfvmLlV3HQ5P4TwQHMXTzxyqy1P3usSHkc2b0xF6
tgS08QLmIF4a1dlIWxCjuJljfcawvGQ+e1JgU3t4i578B0rXj9DZ5uqtlhg5Cs3vnicLc9R1R3nY
ZseToMSQ7NlqhXR4ybV0TamQSjjjDKWdq/GNb/SUiLb8GqmJw8oxAvLcJPczkumiTpnwE0KFtouo
mcsFT1m4EYMF7/+y/kah+nVIUJW/3mGj0kTEFCB8ELKqPfWSAilkB/sRbQHdPHmMLKfn4Or2vTL1
TFXVPCXS8icfB7HJV718CSmEvV/An1cR79BScE6CAxxtmtcfGnoOuA5KG9o/LH/s1K96t5QLI883
M2fCsbK8rBzpgiSR0eX1T45Cudk4yOdYRbAtFXIrc7u1s8tOyl6gmy0p2XbFhmkbbCQp7vYp4xwD
OuGotW0Nk+wucA2ZXzGEJUsrDoAfumyUhpruelPVJN+fGR4rAA82dFpsvU8SNqIRmResYJ5Mj+rm
AkN5LYNwwQgWDgZm0wUXRb47yulRPVhtVn5KaObYiN4Efgryb6eb+yqDKO1ywIGNY94NLKSA8WS+
uW7frS4gkzld9DxcMfa/YXLdFoc7etP37w8/uf4q02TpKWpNLm72ue0zN3sqe1/S+7/Le2ogVuYs
BygMWhffCUCWqKp6gByT9LGyWIh5U+mNwXYTKby2x6GXNXnZbStRe7wKRlFYmN3pmyHanKIqb1WJ
XPUf81EWN/Q+2jShHSOa+Z8AbRrLDzcILhMnWM1Gt4nHoRlh9pJEjdmf+QCBAdg7NVa1CqDKmLIZ
PJREYdleijIJrOzGLhCu2l4F0PfVUX3Pl5VMeY9JgsayU3SFmx+0lA/WPX6+7l07E0cVChPZSXt2
S/ymVEAWVaTBBL3w65y00pN26DNUm1zmpSwbpQfpBec66Im/3P6jQ1NE1ldpknGhue5ijj3P8900
TnPe7VHM0cyDynqP3mw1FjVIAhYnBUMiliftjLEh2q9MqaV/WI8G8BHX5o8ey+h2k3As46+yUPOY
pw+/yxZnAP1h6bei/jb+XG+TV8nThn8lWRJ6S1ecFwHGr0rIYYKnjWwqHhBKKGrUCW3Gq1ACiHEg
Fc8va14bB8PFfG/slbzeQV7MKAoeGBAfBrUz/JApdExQHwkQt6i6ry7q5B5R3uoGYijCVWHVa3QG
15qDQ44uUTiKofhlguj6D9WxdjJqop/0PGpI1YxdDvJWyKgLpblrQuWQXn6AhwxVC1WUJQcn+01T
ravkdptKuUFSGnZ9qXvQmpwuQy64ebWiTiW1bMhmCdaTihEyPZu4rOL4KlLDzVuqPBHgj+OdUBLs
o/DfxfRR+ye82C/TYNMiYFUR6W+tOrprhPPgtu7TSqmHyet90v7q0Vq2IlcxZ3+hCa+S7ykXKMgB
JiNYkTVuGB60C4CX+wiIm6kT2ufzGsLFyGY4S//FCaPi92ywFwEghy8S7eyLyT1xd+zUTvYXGZc4
JWB9BCiueiYkvLuHwQ6pfCT59Eg3UkZBCGNjluaufIytYgZGsPdUr+XN/vaU80UJTz9wofANPjKm
9M0ixQaWuhVjnFMSRO5fvm0StxsIobG3ZQH4hDPOpx6vJ6Qs8v1qWWfyBt2kbLF6P3FNypI2ovSd
Fy3gZPD3PiaThh4CDlSySE2Pr+4OSxn6WzxxKHYtdVAeTDVv0GQ4eYrHvDBkUU3OSMc1zMLbK47x
ztb3tIfGNhzATIk3lzcosR38Y+a07DWbjPlZPPs5crPOSkFsu70XGMZ9p13Fx4adbUaRbUhhvT4T
yWIz7SBNkngyz7k86AIPeD+4Ng85rQIRFe6lRoAca72BIfQeTAUa2IwHtFNovcnrwLRGoS9a+L67
Y3wfD+MqwfgBtuxBP9X8+V9PQd8MnxJ70Z80FwG9lGtmStVVtSlS1onYphtqYcGM03EI2AztY/IZ
AyZp0deVi5f19oOrBAf/ufKYbEqKmJX3p8I/V/Y3fYISuIryyvn1HSutXVB1vpbfu5xYEeIy3OIq
eMknuRYYLcJIxnm2WEvANIi05a4yzgK/e1Wm8LlqGT5ZAIKWcXquNyRvbRLCs4V5Tm2vkcPd3mEc
x9DRJY5SFSx5mvPssl0zCBeG6YIkCJAPBl6Ff0321Q8CoNATfYVoRRfLyw/Gi733O4J+SUXTOVLh
7MmK5Dx+2RLNOVvLfUy3W3EruvGkySyLgKhie0GClhIr/98iSnDYgQXYFvdqHM8PjApXHaBt4G9v
X6R396Qs/8+RtLDkAphSgF6zfcrpvYncpKhCPkla9s8chFfl7uX+LtKUP5Lt9It169i14Hx0/ClM
wqIbjrtZSGSdZyZSSH931YzZqONFZaIO8RXbtokc6m+CUx0xqWaZIRfcKl0FkavtlEzP51f+BR9H
ABtX1rRifo6i59GJ8HYGz7kU/wRKcJBnPBmge2dnmP8gevcTVYFJtto9IsfiYDZsWdhTOpGlYXoZ
hivfDNvjIhU1APlf1oYc1ozSvOEHybFOQTH0ghzo/5cI/zHhMa1QJa/wfprOv3QEjShbBR1tTBOa
T+zrHc/2+LdhPlTzmxglfqiGAkEOrsWNQ9/qTcF14VUR5JL1zywcligYePbJBzY2dTZPZhMoiVHF
yV718MWFws5cjWGMA4+rYAEEh1ijedtAMQ+PKIdKDzMg3S0naYGtPCmxJkoLBNKoM7Q69LL4r9mD
mCdcEpqz/yNTraY6KylVhFkBp6V9BkQ0PNg9askv1pkirrgBO7Zb912vy01IIVf6MZGuzis4FOey
PMWBx0SUDLsUaSpfKp4ii0T/GpN7yaLwUynVsT/QLX5ckogn8GHt1EP6j094jCHAoFx5aUAOMG+s
tLjgKs/snZ6E63UV/hFATlBCn8jFn8zxX2zJdcpTT0ElbdfpgTiT+uvq/Mnf4tbgezWS5+jl6l7L
0lbiizjH2ljqkB+rJ3h333KLDqBLUE8kx+vI6iKTXM6OqUPZmxm80LWWnpnqwIEQgOpsxK8rXSnh
VkVtTLinAs8YpS8Vhxl0zn3FOQ2BiZ6HttIFpxp3NXchSszYOrox6K6Xlzpu6I+WkIv6G6/IstuR
WK6hQYJ6zwwRVrlC6uW8jGNL6crF2zUVd7XZSRlSrBzu1NJi41F5JNDNJoQ7slDRAbek9lnG3//Q
hIZsCp1nyjxlwt/b1Kc4bNgin4vxZ2+kGQU4cadIGjJsrPxBFfPbReooj0ruqnErDMx2ElNTLm5y
ifnRdmh5gWoJVLYuuFAfV4xviztTxC12OlBHy6oH80H3EP3aQ5SXQm2B1QpPZM2+TlbCr4YanBIw
EGJ002yNjePRx5uB75bxeg13ck/hDiSOpZkN8WnsSTW99EO/Plrn1Mug9AtcB3xqw2AqAb1PBcQt
VyP8ztUSitLrLKrRDOOoe8pXfeY44jdkqllWvEcQ3wjv3CmBZHznNuZgkQlGLCoBer5keSeT2Oxn
kM5Gol/RCTQN1wjoXoOonFAqHTOm8/HXwfk/nDzYBdlPQ/d9xk0+sqIRZYVsYgtx37r3KQ2oOzhK
yHrMExuVPc+HHlBLqF/ebQ+cn8JjKx1c2OnzsDGvm1LXZmSV3BHTvgFtTcR2HotS79NExs+E9+nu
EzVNmwPP6BG6WyOb0QmaZSWtGzDWPJ8+FA2FCX1xvtqrcNvYHWUkDr9jaoOIuSlm4Jz3Cux2Xb87
yqNXXE9ADXg6VH0+TW6+At6SX8NRuRu4fMVV2n09Brztye6bs5PkLKDGBKKXwttgpWwW0LE/5348
uQsl/o9wpXpKwaW6T6uxd2205lZh6PrxIXNmCgiouL5wRxwtoIAb7jAeDmTieExmFMdgWJVp8au/
BW1TMZMnwfuxJyBJH2Y8SVwELUFJZ/yjYFLjl7bbTGu59P56Q+oOdCztuLD6eM3DXLxBXBza49vJ
T7u5O3Cr8fgoMTEe+kYm/Oa2h1Am/Ez2ZRg4SY0kMsA6NZ8B7d7/ZGL+ZNnP9Cnl0YKEsqoy+l16
HMchj2Yv0iePcvwKkexU8U291mqsAcINy8+ZlCFytkZDTZj2h5vLrulclguDUIAGRZMVKl/ukbLu
/nXMJROH0n4NhseCe5wdf/+ucgSslShSwH9i5l08HjEQ0pryVf8Y0t7FDZaY/AwHl6yeU6+wmdBi
6hIuVoZxUpPlrRXiuVfR5yXacp9rlXG6u2ozR2+pkhcYF0IL4hIYO8lDlYa6bazFZZ2APdGfLeoG
ngIi/2rw6x7KWQJfagm6beWDJVZSpu9JbjSwhSH1kMMABU78Vgo8OMO/fw5bNaDXoTYiqfbBFKdj
yNP2byvKGH08LDnAxseQqhU3YqpyEdUJp5py9DQ93mcPDfAMrDKOgY7rb/uvP5vN7oTeHyNc+2iJ
bxrzXN6sZ01PKXGsntg59g53woPwje2mHXvF+xzZ9jtQEwuXIx4bNBtkyo+aNeLT9jI6vx+9m2Cx
F30dE4/pMGA4we86Vma8ppO0JHkKTcutN6tZkEQ/+TfUyQrQi9ZL+TFixlYZkr7kIOAqrs80KDmR
dyEH0kW44W6hzw6dxs5V7rttL2iOHXnNK6/DpZ3XO5GIfBWpUZwErP80OXR3cnzRstAK+5Yjy2k3
Job31/KFMtAlgV9jIkbnSMGvPVXDifdp4IOEi3uRLwcrs9WNLzWSlLUT1d/Yy4pcL2YO3CbzCt7C
3pnezwrYf5p66QZm7Jmjga4IZp5xItKqGhVnXQs8rTvOBRfcuKMUlXTvuhrqHei8z6mB/IvW5f6Z
Ut4nXMwGsw2qODaoZ+uRGPZjpkSuSA9NJJsB+tEUbspG7DTBY+o9nSt9WzIzzqsQ1kJgpDdWdYWI
tKiLif2NmKMUfSfCKbxP1Xk2vr5oJiJgzGYUTSbsB8jtaVpshsbu5IaNzN8uIq9LtwXyKAnGzbiw
RvEGUlgnpIqmJRdNCzV7BjrPbLlJ4qv082cEdUR8YS+lhSDlZ6o2yP8JvFnNOoed+moL91RGfLaj
GkfGldNsH4XH0ZyaWYqCuLWus85ITtLudKzAuFbP4oKzxm26+yNEVT4crih3BiN/CIMnnFEXDmHN
vUHLTP52tx/wnsyXwHZYIIPv3nHcCFIHMXDm+5fzj9uBadEpmhl/OJKvPcQyvIRolbG41LnpK7wl
zWK+X2SlyDeL4h5phk+JtWH8f1suNoqk8GnT+cDu8jeLoVMht3tWzylpiu0dhW4/ug5bq4gSyI/I
MzyZKOkq8dwbBiozDEtNI1zO2szf4rynKizl0ltnxS8uPgb/zUSqtZkEJWn5FJNI56NZXizW2i32
B7hDzAM1f+MtFRPMTAt+NT2qqw4oRcjSLfpyJ3wODSwHvS1RPhxZ29n2JxN5uT8X8c0lvt0IM8Tw
//4b3yZei299iDOfSgVONQi9ejMlkAPxyd2xT/v/r0UfkdNZgDnxzMdvzBU5DtjSqeM5EsuzWdC+
pLuQmmA72fyLzHTuQDv+DFxobp43+FocvhyvOpDiy4hNAUbzxWk8MNm3DJTw9QHxlctvs/0QYJLO
zUlXpKBqki439/qgVSVvWeOrCpBVp5259lhfOO/kKaKxHToBXJkdqIrqv0rxKYDQgS8pV+UWiDGt
prbQ4hHNqAyYpyhfDSGQzTIovp2RWr30xSMgB6wNofx3eXQrbtVBMGYRiaYWxD0BYJDURqntZVpO
9HCIoWftK8iemperjjynQU3N+F3v/WGaP7JQGhpPgd8HdcGS+hV6Wu45sZJ0Umf9Ma4G77pjbA1z
BHSgQ4Kp3U46k2Z3MohWQh+/YU667l0zOSlr6pEmpQ53CbCHynZn9zjE8izO1Y19h1olkbGLbymJ
qaIWoikJR/QP+VzwJru60gRmxnqUbcCohE0WT440rSkiMHloXQL/9OJ5re9ce/ycnpc+5CiTPcFC
04/2uwrJTV/W1ysXTRnrFTBYRoqXY9wZKtVdUOCv8MIPbjsv3o10B61qskwAdLwl68lc5ETSvNTb
Yy8S3aWcPJ2xUbj66+byQtXHDl3kny8xd9ftWFVwu7xoQhOjCLEf11W8VMuNKI+kLhTi18GykrVy
WE+yVEi8PSPpQgPOHcw+sXomDM98P5wCgAoICmWYbqoNqyYJVsyUElxHr3ZA8rwzrJQ7P7YRHwNb
z+G2cGxxW9qMTDYp5cq22EmnEiFzrE00WZ//pWMyyX3uzRb80FsuS8rOABOb8v25QMUJVx5k8p6M
D/V6EUje9BRp8q+M0B6wlB4DJiyRCaAOhYXtRarUlOUvI13WdommfPqGbiDGYm+Xdgode+NNHLj4
xUYH2Hup+tQqq31GQBoTb9j2zUyTqyy/8hgAw8ShnCOQJ7DLLIepEUFUToysC2LlLuNmrJGex63w
wwbAO+5Vx9wQo3Yv21iBiIjakvPWj2aZzI/M926efPEYw4hEGn5j9XN5sUeZ0496eFym9TaJ8yhb
OuG20n7nRQwQ9sFe4GLWhrorMpbltldSwWfOS1hww6+KDuHXPhn27v1LVwMmPKgMf3B38DooRspe
UP5QR6ic9ozHsK5RTNI409X8tSSx6gcnmD2Qp1P7nLMucDT7dN1sdkz8lmLyIHV5Io/CFtr2+vq8
w6FEM1DO4LOOhhSxJDFPnNC31VSUF2uNzaIEpdovcK0X3YMkRCKRSuOfsskaNNsuiVzJmpsUKnl0
MXXpUgW8lHISkeQiH05I4HH31bTysnHs0a7rZVrdlDQnz13iNoA3eiFSnWp4JtsDzgHGyJJ+hoAx
MVjJd8RiOeuHwpjmacTDemKZ2YdIMYoGycV5Zta59iMjumuArB/E5WOQxPg2MoWaTQUhvAOP31cC
SFW0kTh/kAewJr5nH+2uZ8QBt0w/VF5J653MDEdjNA48zej5u3QD/5mn4f0wd1UlVJx/fqkSDFPL
tjGhNFiUNisSMT6Xk4CJpOgH4tFVsI/OlU2E+Pc3/ba8kdMIhOJTP5apBcuQWjTBZrEpj/tngx6J
SyugaucHg0cfIpaq46oHcj22obV/myz3TizbrhD8FvT0S4ep7co6ZB4BvJu+H3fJM0D05Iz4D5xE
GlUy/CaAzscz+JkpHSEuF+3fu/N1U/tzYxX4VK8m1CP4WARBnY8LOWihiglYmacDEXK6zujpVJxq
vhDfmW1LWVqaSaRiUhQSJRKMltpR7M2sw1Y3+E16x/GjMRC84/9XKJTwjSaerv1tVBfPg2PGBCFP
mUCcDFe6t343YwnxMDcfrqB/w8tVMVUrd7ZxUYOUe4lI4Y94WQqTp4dU1SNYNW22n6o425Evp5D1
Sfk7raptEiM9WiSqCH3YB12Mx2ygl85oJLnl8632D+XUdUcaCpAW1C01bVS2TudbWU9pcMLPvjGA
5fFh0lLNqBIhPNYZXH/vvnWKw1/vx+pfkfNv2Zt9erj5TPfBZyr8IFAixM/mBIb365jupo/kJkYH
SEVkKFdGlSqhqanhR066aoeLLDRGfMaLWlVE/nbSHIAdQ/1p/LCdBaWgiod3X6y3JlI9XGi1ku8b
7yHOQpgrgwJlghjPC4fsDkgLxxZBUevUo5aGhVxL2348zHWHKIbwPVyCxpGxsjTWVGrKDMmST9/f
Z+95J4crjdyNk5X5DsgSp3l7Lhxuk8GGMH74Kh1y0xSCeFiYLRTIJnWU77UEcJqkcw2s7m+DjnGt
a8qiS8Arm7rX6K/wLhqrXPuVffRmVIPTh4euZWyHmWZ2qpzHvGhZOHw9v7V5208E38aykeW9OQUQ
MRtlxx2U1NADvnXcXrxEtShziKZdaTxQ04pm+ZdIDrW2EDMe1g7+maLqwcwEHABZDRr2Am1pO1Eo
7QI7ZGI71ekfiM+jOaCTnzRYmFuESjnZctNaFAw/k+nTk/w0kwK6vF8AXYLa5B8EwlA9tnAQFcHJ
kA41VtURUVp6D4EeWxX32/khx9rGdZ2gEjNWB6G/9gJYpPciFzdvXfZvGyPiUX83u4Qs14G/H6ZI
2bZla5JjtAmTeHf+ymtP6msUdVEKkPESKW1vvJOqtBw6mdlMOjsAmvHEsBPTwl4kB7J5u++S1bx9
V3cr8gi4Zn2jJH7TIH+zjjajIuhAxOSu0Ek0gvjqtzo/8uN7pyei/hwHQ03rO85uTkdvO6V5h9YQ
gyAEOCgse2BWUJ1L2ozdhlGvQVDr/mtAXDc4oIqHDGyhfoheCn0Sl/8O8jzuSFgsAsGO6S+nZZGr
WMi7HhnopgdVRTtbuoTGBBSqblqrDc7b9Mxwyq6q6fOC9TM5CcZM21BmrvxOM7hqZ1hnb6htLsdC
/LiUG0EFX7d+BKbYj8IvkgfS7jVfBPDj2aWI5Zd/P2DnFtv7VwjE5KD2BKY3Dw/2df+fRY9uNmhd
q3ucBcpWRKtqfJeuQufSesDXy0MozVKWcapD0rpjz8xFVzCuc/arxRFUBd853GiiYW8GASUHv8Hz
/zfiJLbOoDboq5CWAoB5Wos5P7I26y18w7uEdNV0Jq6FytApL2BjdiJCqBHdQmiWuvLo5UFnTRFL
qxKk7boNJTt6gIRy7SiMzLjXBWfv2B27wojCn37g3up1pDzpOeCNpw8UpWvYfl/KhdRDyAaJ1y1j
E9gFK1eKl9/DpdPUMboXhT7soNG6uxZYFYsiHyvl02ZCQyu5JjGijNB4hxeuHNya5DAHxh4y8Nd0
mj2m5NMVZPjnxdDMz01SFyQb4Vd8AtaiXqA6ulDGg2JdQ3fFPYhgI1KgSCLBU5Tli+icputIoJ6b
I0qZ3GTJlgIVF7ZVAZpPvoumzlaqYOoJpunq/5gVZvv3qcMlgbLUetWsHDPxWv1ZgScD19wK7/0q
BfztrUXoWM8fmFD60Fg3xOg60pE0+BFPlejCbnbYss517kVV+rxB5UiqDuV63nCY5HO2V9r5u63o
orBcep+joUZIrKvJGl4UZqs32V4S0cJ4pysmSkYaydWbKf7rpSI8f1LPIQxB66i6Za1BfjrF7nC+
DgSlhmSTmr45ovlp/cI/IFvSIatntWz4PPgWBRvuFJSFazEoWVP6h9/j/jN1x01Qy0YUxjlQuSUV
eh0twrSg5+2eWJReFPYehtpRbMxYDvUxPUTAA5PUSlDT9oZk4j0/IF7L9RpkKjSvZkW8n4pAo42/
ALf1qfILjOBIxbvEeHXjXoR2BrBwEL7mhdNYW0EJv9FEpcEELzV1rjBn0LRFMI4vSePQN6JIYtaT
HMnYwzqexZg8/ZB90nfGx83RY4hkAuH2fk0z2sar/hVjL4ROat9iIpKEk+Dkxv6Tfi0+xpiDq+sq
VUPLORVmMrYBP3AUgx/8GKoXd2Sf07mZNEGyXlugarGIwmTBfpjvE5YHpCfmhu7m8Wo9sx15CUDJ
faPW3X9P973j38CF9lZSN7wT9p4ATtvpTgvaRqzBvyrw2jWfMHZ2U1Y5G8818OX/Id6NW3dHKf/z
8Crdp1uKSz3852Q25bbW9MDVQdCpyx6Pyx/AjJ4ZxlBl1wfrSu/WqWAlTC9DuBw0VUwUM8YeDZr/
dQuzFxKuJWcwR/xfezBv3VILVFvowV7xslg1YeNTEaEQpoe4F+RwPHE7ziNAu+e1x3KPqSrh+Vzd
FjK5OU2JWqFKpN2xQFJUOPDYjHnUFoscCpVsSc8szEGjnwlr6T1BWXvm8uNfnjXbcjkUCPLLTa8Y
kQkads1FyDOf3C2HCswyIMSH4ZGL0OUVEKjV7tuoL5K5Hu+snG2PznND4jPEjMqxBB1qCUkCHdJv
r0knajvcT4nYQ00OTDVIjJ014BfdSscAKsXR/N6rPhiKHDVAUlWOXgWc5uYGvC9A68+IisU6cdzj
4+DirNgfjLNzHo8XZUOhELcpccQmC7DCROVFgE3e4xvzL3zjLBtGUqEQLfS5OTluDSuJqKUeqLrY
B2G3rZN01YYRiePrU7F0dk2h4HVSkIhtLNsRfk8g2kUY9ILfq77vzyTU0LksQ6QhOdW9Q8wZ7O5i
OgoBHY4Z9j9whfTYDwHPXEYg9Qm+8ICUAQ/q/vV6ATCYHYVqJ3asEz76cr+CEMjhzFA+g/899bEN
dXz4FnWO5brVvs/tFilO7u+jOAci8JHSO7iPfkW7bmiS4xXlJOW/gn6fg4Axn0P9WMn4u8+lzrxW
Rv7Hou/NFTjqKDAPPBwxamivRjZmG7ykagWvx2mHv9CFERSWd3cuzgMszkFA0wtdZ+FyMQA2zqaw
Pnx+YkdHgLqTeOEIUig4XyDAw2fhm8Acr87IoIiCiDXIV3DJL4sQbw+gTO7AF8TFk612hKBA8Kad
0IFKlKSicjSd0tCKpAiKOpM7fxST8YF+7/mVo3I7LKiPbJ1Z4N9bxvWpkLTODkEQTvv5dvs1ybKb
GfQx8DgCZARUP7n2EO1YZcIt/DRP/dCZDsafn178ONW4Y7vGtKbYCqOGL6KTKA4pKJqjArrNPJTT
IW7/kCMAEjpCzShvWMzriDI0lCxU4OM0OZWt6fdXHkEWkHKHXeALP2wotgEckdkTVK8sUD4WLpb8
8dzS83LVB1yhLvzQ7OGtBFWSsMCZWlCmh85BpFD6s/8318x7NFFNQzoABjzBaBHvoR9Yf9q0Tkww
2wa9s1cV72wOeg9gs1qwbDwzK+/TNZ8u/ALGnn0j8Hvqqt0vgAtALO4ufFJF/DMHxjOR76Boytw5
I0/KagsxZtGjI+j71/ha2aQp7XYaIME6qWBrMCVceNeAogQw+9RrnzOn/NrO1qjq1tgXPB1TDsGx
nNs0p5GjXkJU4J8TJwpI+NxnB6sP+F5G6hdm1ly6aaTSSuwnB6zp1d87ib6P03Fj8G4eFJ6ItKcs
cLqstQpIQZ94Dk2lyt8na7Rr9L0C9jFGaUrReHATHaxieR7lcL1d8EGoNEiHdUYXw4uNTMAZhip0
rNGMszdZ0ypcw3Sg0o2alPGgVG0+q099Txlkx4m/Ll3Xhliltzrung1Nfs/89eKRRZFRkSF9gEQ4
YSqAMSDddskhtITNtT2sdLNWrOcAuYgoO1If7U2GIpYs8KrxYlVBNmzTboY+XYE1JKnJnk++3oQy
K2aFykyIKlpAxi7z6tDdjOYGuEyb6TLTje2bULYCbcExJbop9ptvqibewj3r+uyYsX6PJNQmifmy
SGj1Pte2xmrRSh1zWx9ZwGHHE5vi/jiQV04JeSFSVnqrKVoOvZaQe/yv9kRsg8ucSssJnHKs8Vc7
IlZJc0fWOOEO4NYglZyizBrAGypU4D/b8f09ySvC46U5gnZHydkmR++gNRnlAUHAEnAiXGhf0Z+G
doLw0yiVwmYRYhA5gkT2LgKjHSAq42E7Ufn+yyoBQfyycT3pxPakqSp2A3jkvqPKuSngZTGaW5oe
xnfcE2vqK6KUNa4ylJhGtmSNiHoRaCxG/SII4gys8AUA609j51kt1qj5pdAxmeojxT2f23qnb63M
MrhXG1Xk+Ujzhpdhf4fw/kSmOfjwTVTYc+BxVGLp63QC06JzLXnzr/c6qVQh3/1TcWSvhbyUBcUP
qyT1f6nmeS28fCCBnGqaPZX0OBDp+sV2pWHQxCLyx5bIhrhrRCn3AQ20qZIlbv7zv7Ld5SBB6rP4
xrDvdoMnsTayfLdOrR34lwKeFK16q8gYT2+/5jbUCjLXYDng5056E7HNZ6nRP5igUZL0AaDJG8+g
b2UEJqPbCJiMyA0nbI6D6jjjuVf7x13Ftu8thWwonZt0Yk0aKxZwdmjVWhVIPlTqeo5uSZ3kvbgv
MihrU8Vv0f3AVNSz45ldmmKSlAcJ2axl2eWXZfZV5x2rO61ZRZPMMaO36YNfm+qeHRV3OVIXK5rL
FXWi9pwSZvG5woxRIN0+H3Cy56ExYP+Bp3IMT97F51+/3ng0cTlMkuo4o0LIaVza+TCUCFfh9kyc
DHoiHH6qK5bsO7tYt0H+7Jv6CIOl3822kOm5KOfE/v7Oano9mjjjYUKGi8TXbLrVgUJ0CgS/z2/9
nGOVCk2ZsCx7rXlARkBDsWPtII5kJe8K+mjpATvcbgW9lNL/8aoprO6oBpTiu04AiRN8yr2LkRUg
sufMk7atFbzQcrWtb+h+QohuYTLeQfdDRnCJ1Wy1SwtB/44jenEN42Dg1CXh1QFagfeb9VROVhrE
sIJ8i/0Eh7z4DchMjXT5aa1KPUykyrb0Z1HUmqkykB085nFxXB1LRi9byY8GzzRdVk9tHpNl0oIS
2qOk7MIDiWSCqYiQZ0TAUfaiE/rO+NXaWa9woySar9KmhwavA1A0RjCPriyp2AplLa9OWlUDHAKD
6m4Hf2eRprTE1T6oxWT6y9le96hfO1yp6JLmu3rqxRVNjt5z1ySc3zBztYgyleuqecfwyp0c6Kpg
K9ukiDis3cn+ALBQB1q31JjueBkZWA4RiPRr6i+hiQA6YKXf5WceNyPRRaB6k6lvtVIcnzN5Xu17
p2xxiGduA/Kty5gUM+pCUorVvrMJ+c5eFq+Url4ayyKWrQIdtsHl0pfZUr5BSAEL81EFkDL3jCKI
hi+GCydlifAWHeUsZBuChMFzJArGs5oPrhMC4HqdGsFstBxwz2nLksnLROvBwKSKT2DI4Wcs45KD
YR3CtdqCWdXNOwYk5+xLBBAxNlC2+cwD/hVvzhQ9A8fixjIbEAIMLR92DF2Ln71oUMWfbP3PC0Fi
G4BPTQpcpCB1BeB2MrLJARFzhT4TNJNK6mt1YltbuXUDBeB+CNfWiyLkIJHMmTkZBKdpUo6cgs2n
QQpyP+egT/fZaz+k6yEJNoWR2zwpC8xr9VpZXNF2Pi7heocODzEEemFRS1tV1mMVVV73wjzz95l7
o0W+WXFhb9yi1cBuAKOldO6k3WzspBm6TpFxXVyCPzUXWooW0ood1DmTIkWzughC0CKN+dtM+7xq
aVGRHJB4u73D4HaJig7AALCvbI4e8G4u0mbqVuAZrkSVqsTesEigJH5RUP4POQdOH+NoTVIPWAke
aWbKXHB7nGeJ99qh20OAylTimq8TbppoJOrwv6NW6aLe3NJrz8WWGBgM0FhmqWKeC+sVbyxg3Wo2
9sPpL45kFKpBrAmqodB7wjdlnDivMxntQUGrGwx+mb8vsxKA+xx/s8tTPvZDoz+DsC+WllI+Jfrh
5EoOC98sCTS/ellLq2Opl9kSg+a7iB/eTlHItVSrGTpjR4ZtcOOh0X0KcNh0U8Nb1+HIF3PG0Ezj
/MBDX+2unMl5jzuaM6XTfE9hYSPCwq1+ck3zG6v8tbcbfc5s4Dj5Z1tBpphR1vxDPTxNpEZOcZa5
vvGJn+VynIyfx09ZaKy/gOwH/6kZsiGR20XdVvG0lruG4xHb3rxMJWx46e4A1rJZdTranpG1YH55
VLy0s/uHr7xnuU2/g48q0U9j4lEGri+z9hvcHqy3gYzn5im4xpiK7xPUok3pnRYgHrjiOYinTqeW
7jfriHAZPH+7waFPaz3U5wDFVUKXDxDwYKh79Kn7zedbNIX0YNrXAouwX+Hv2y7+5vfFvjvIBeNp
klkFwPkqMandDPADBwYyn+gqb4kM3WzEDjqc8uambO1FVtovFgI8072oZJ+N6RXIr02aW7P72Osm
3o5m4wWKVoVKfq4F6iYwTAC4lZnha7U4HBlS5iYUSKEMIgTq/3MMVZQIdKeAPpxmvACfleQdv4YD
ZRFNmxtMSsl7xTdxpRjMhWu1TV0E3Q3cvtHzDH05W61o6RLoODMALhBIDE7Voj3lE+yGfMQvATLl
U2mfjCPf8ouGBVUTMVQVrZUGw/glA4zHUNhjiqXU/Mmz73pFaOM1GnLKg5kLlVxQ6GVTRxROR6K/
FyvwcUkd/pVa/UMMeYuxm4NIgyhq8fTM3WJ1EJwutEicILd85ivgkg1W2iedu95D3NELoMf0kox5
xQtOVvbTgrhxIiDraWu53EbO5enIXdtZ5FuwkcbdSD9gr/bttAFyTovb5Ap17rcf2VC9sPXNUF6m
B8ejFFMabWfPsfrTH3f6fW3MfOIyKybQp3V7j0LM2FwqMPeKWBH9B1/kJEhUj2X3YkuzYjK9L1ja
kgoh2U9B4s2vzG81eWFf+QRiksk7L/zvSf0ugttDYznBZkJiLwNQl4EEv+4rfBEZ5X7+c+soNTQl
eIlhCy4Ab+fzCWPKhF0GLea3vqOlOHI3q4s0Ewn5ZHRPTGgcy9MtYu+ogpj7Mnn3tA6lry+qNewv
ymXo59obHJ3nX7G7d74vIcjEnNC+14BGGRR7Pi6pcgNHvwPuBYQ8TyK0L8wD2yQEWRKSEA6IKSRd
Wxuf/8rxOFljFs6YWwDWKB7+ei4E3M8AHA1euqekuHKxkN81xjgmsMGmEHzzx5WfBnxCCvC4uw/b
y7SSTPWnkpuwc7LJOk0PB2WYr2+LLkMBg7XIXpCrKlBjaY7fzIi9YZg1uSR7ma2MjEcoz9tDIeqY
YW+GbI0LTLCPjUs11ixYmJGZKql0iV4lKlaGAk2d0VH9eIvtr1sLOipCA1h+iUUcDkiK+CfJVdSK
otXlzN6mT1xSlny8zfSmn5EOUjKTat++P9sKMFgr/XaCbxcIXWfemYTNm+ZSvA3At1jrgS+xN2Rh
YlSPFxUfB0YjIqq7SlQKGCAqJzKyP+dpwClWAMc4nE/6m81UhzHljjyr/yAUcBj+xHAf9rAw4tbC
9nVsTPn/LBzXkhG0teoBRwwitWaw6yOtggBx8ejPk5dUkXwQGiN2g1/POQ/GeGm01ALzMM1jxk6V
LDBQPRIP4wj3FEaOyS8kSbunR1O4PqhkNChg8xn58AVFfG9QiuvB7bHkgFGVd2xJcebr2G9P5TFg
8OEGXFSB1B+zPtvyXZTrGa9eDlgoL2bP+M2tgCEeT5ZRb6ML7h5SEJ+IBnpQViDTE+8CEU77IyDJ
OUdOEO2WQhCCfq0deWnHIL6kPnUrSUwLHNlrR5xFZOBKq868jg8nelRlEfEIC4IOtYPgq6Y85VTH
c3OsLSZBta7G/GHLEVKlbxGhE0ZdKq2423BBUfzkUuuklTVB7WfCylXs2Wt6VAgH2lXt1dbd78ji
Stq+TOxPgRhG7od+6TAV+DCuBt/PlXqHKJYlfD4IxVy9W39fF4Gm0gUo4kYt7H7ApVBiWXVN3bte
TNaM5gakLmGM58ZSDGHMO6OaU6+2PaNYT84UY1pFpJkxi2w3ewxnX75WQcJGfYXm63ruJPDEPWtn
GB8u/aFXCikSIvpTinQPY8QENaEGoYIKlfHbdgAEU1W94wKnZAYUYe+e1KRQsTXwve1am4D8bPeJ
einAGfQsgdJPY677qJEzgpCnIwsWQNlGmJWo2K26i6PS0J99HdMKDrEZH6quKVcuNEKN7mm5clLJ
EnUHqtdyMQKvvlBsQGyXfjKj2TfjBfb4w1QkROhqA78xXaM+q1CF4abjqzvLisDDjpBX3KAbr34o
FGoKGy4VH9W+ZDweq8X7T5IcIfnvG+/pb9ny5yyBW5w2QSaisB75ir7Y8hu3HehMkLqXUzv3h7EP
7uIu8bn5g6dnplJ7mxpBqQfe1jx6khN8u6a+FzymR2psn/rni+X2hqRTTy11IC5hxaGX+3jp04AJ
tfxv/AVC4p6nqb2/l0lmVLRppdrGekTAsSOIjj+Z/Jh9xajaoLrAErz42bBX4GZ2RvD1oeLdaD3Q
QhDmwXbmcvvDDM/XwEHGpetCQuv6ny1/nlspsOFJO7hB9u9N4UgD7rFNktgS1LHtbabDdGLW2lw8
7KaDulkuHWb8r78Zmv16tRmCk3OMY9XvzsAxP1hCNYm6d7/9FC7Tg3/jjp9QT6SvSk+LKF1Keoqf
Lf2nnlyleVekkPFF0BRZx58Uxnr7LGxMNVkMU/MyD50mN1qCUkbp1Z6NkZqWeiek0LtcVI9D05D3
QV7qB3RAs0NrWsr5LVzrSPs8PNekHPp6HK7kTZaHHNu62elMf5DMEvvjcVbK9KOR94qPmQrE+pfy
4gcQRc5zdU7cWck58hDurmW/o2uYpwzi7a88oqzCUds4VyQyPGsTh5bpn9GvHZHltwfZaDWPXV66
VFObj598j9B0/Q1Dg2HiJakY+WR+aOaON0ebo+IdM7fCBRzwrWg7fQU03qd7A6gHFEYLVFRrEaRg
fAp0kVkvGUa2z/XVdsbbgcifZHBos+A5xedGFXi1Y9HIwWHNirNWXEoAh5QUbMWj8zM12oTj8q+a
ppUngZ9tu0i71UA5D6titBN6jvuvEl33Xuwo7ZKytnAAyQlpSgX933YeT0tWUlbzZp2q1z0Sa+N9
h3ClDlRP8uhMbV248SnON288O/j+ijmbvvSohD59drWXtw64VyOA/qnL2FGxIuKOq9B8qWaODcMO
CV3G8SLVyAmWs9ovCm3NsBvduwRzyqmgxrtBZwOHmrGrAtw6scpBaVkV78V8H4S9x/qPDqLWdxMQ
yvPNljP1b90xIGQ6PhUWH8McKKDrzuJFYMiB02WyCNna5JInqDY+n6BjWABR9nj0Ibocwb+OFQ+C
lhMt3OTo9UnYOnB8siXswR4sbaDFrivxIH5v0zehRdVhnrrdDqXFI8ZNpyJvoHUKEbyPO909/rqL
PwdbLx40YM/Lbgh18hmUKxrAgL3j2NNDxOUNKHHB2iIz467v3kQZZ+IKSN11BRLOWfpvucq3FRUG
TcBNpV54EM8HRgOKTdEXQxamQa9nOIaeX6PjRhH4o0mgJaBl7tOav5u1JgLJEIx0N2g6Vo/51Fhf
gMRXPyyosp3kcUZhQYYSM4meYashjZksLt2wSnkBmI+CBWvCBY4Nf4DmOe3+qPMQSC9aT2Csi9jc
a+fDA18gBUUPd8IBnGrOGocPXwxoNDc9psXb0hWjNwB8aph2A0IypIxE755SnpuS4em3R46nGCSA
LUySXeyPJoQqgM7MGU0gC975N00bj3rt5vDi/u8oGxj6FrhDxM309+adB5oY6/G9rTFpHQKYRb1b
WqI9vDPAPh0yTtQG9KUIfVb0s2haIm6FTI43GCmdxwOVCeGL3KAqFNrzU9FnYKR3tkV2lmA+oNsS
caE0AgZ5sIbJrshLrqq3/4DbOYMxsk0EQXuMJ3AsmuzoOTWAjQaK2KCJdcr32cegcwRnJfb7xeTc
xm70kGIiFHmba7cIXoTMbywZHE+7tiD5aESh55FxuDYrwBHLvWT4MkarO8CLHiODod2ezLxZTw8q
VBOtRyVuTWAxEdh746jMvEseNkhC3IQXzdaiAOwbJNQ+yzDvPMcPuBVWCrJHuLUt/HgEZAFKtHwf
qUOaQpkZ3qsnjGVvvIEfQy5IPUDbNs4IQ8Q3nbt6yl9NYhX22i5UyP57rxMQGWvFnZqcS/RCxfpc
QSs5pQt9U85/P1FHro+nOTU1sDhJQt/d8T/AK0PYq3LMM8MHfmFBcwzDwPbOSaddA+aAcy4Uj1bG
CCcW0Efc5JOr70DmXBrJ74+BoaWTKRwXj0YW9psW3fwb+MV5lvrqdR4ydZTPmi9oBVTY98OzHdpi
3LzPCKbxXE2yHLwzd2xMYoDURxu6v78nYubaKpLP4ghXLDcS/1t5iUiktx8/s41EWW6cgcCzYB4V
/yWCV6wIBqmvB8EySWk1pqq2WkzWnyx3SRTEHAWbFiNlg9nJb6SFJqabajxQMK6c6CjqEcW8O329
bAT+pkH+LKy/wgnsz4tgbVgdMjC4mzBwEvnTjyQn85hdEttRIdGNRyEENbycvde3wmflQyfPzD5B
qcnHARLavElpnpgM/sLzw8QUWm+phc7DwaOf+IjxdFL+2LStDBrCIPu/YaxBCu5Zo4u7x9FX2YH8
JTSTgkguS63yNM1lPfLZfGx2w2RSQb567QqSNtTo4fHxhl15NSxYcEa34vYyK51IkjjRaZhz1Ow4
CdnGAuB6MCYOzhgazaM/pRrp3DqFpUNtMNtWixAK43gwsfGwJKDspEguMMV4/SLcc1QJesw+5RoZ
oXVwjmvBGYRS9lak3X9raz5/iU/tsmOyU54Wja04E+ci/PEYwMxHaTeojFb8fFG3F2ks1L1Tl4uE
kOO+L+HDeFaJhd5suCcodTDCe0mb3I9E3PmgHIl1D22XeFdUXaqHnh5zk2BNX2bD8mNe/x5pxS+8
mEBRVxbYQYnH2FdA+mOo6c9Pz6gHdvubL8u2KfAKNwce4EDU6uMBxGYf8Itoo6VYRVAWO7s2onzy
8lhQ8KoVGURxyqogantBjI2FiEgc/1rcAmBaZXAbUNWbzO+3dvnLXBPl7HplvIo/FuLQY2v8k4RS
ea68AKw6ZbaaCAgEWdYXaQsZzp2qCpAdFJzJA6eVkDQkz4YxONd5X9ddi+lApO/CJcYpQGy2IZlX
1PS/uKJ8XfYF/TDkRxD4DGCIQPSbjb0DQpbb+iJC6XTYOrzB2gyC1z9AjK/5+ArotYJz9i51fYMc
UBrf5dTP8LGPiT8hj+A6IfebuVTfwq0C9OvqI7ECbH9wCZlsjlfjsKQQ4oyfZcdWASUeafml273Q
wUwttLCwhiOY1QcFxzBfLHNSWuASYOYD069KXM5JxQbZ7jxDkuN6kcoT0/ppck8zoAqE4Xe61rU9
rItiUKTsJY5WDaksKjVkKhrq3w3Oc+LTSGU/YFSLM/c2xdWjjHfOLAcohQvkXV78eSinJUZPzd7r
x0AqqMsrXLyTLAa+q+/87o05mT5wL3z+BWKAIJoA3QFuFkaFl79FHDeeUeuwCfi1A/S9EnV3Himc
Pfdzl2y4BBC58U7zPE2DPGaL8mprh9+bFDcsxYpE0XtkzsPPC+OJRMtDN4bLQ1idErJpFcGZ/jBG
ULt1/xaitw7+WJTseluajrCOUrbnUqwkDoJNRoAWqYjyyc/gEs8KH+ZX0ZD+SOEEidbPvRJdBFGq
EmP+zT1i72Ji72qpNqo9hGEdK/ZfUIHUQ4EvV7l5xs7xDEX31qN2EEwKN6egAh8t17cLiQzY6tNJ
/O5nMpNZd6xOPQfwoz11eAeAAo3X/X9SRLB0Pttwmv4uD+xiOQKXJNf7YlBkKC2oJXvhzMOywNNx
Sxrj1DUBEgP5CJaAv5fZN1hfRIhSPbnbm5tP7REygkbCSk+10vpUW5CVdjwM9OdQV7bv9n9h9TM1
PCpbZWzjHO52+1uHXtfyTLHqptrRvTvDwYEYGABRh5UEh5FPo4tLtxpMmY/3yUmfOzuTndFVLbXy
kpT/Nzl3kWfifJ+hLF3Yve/xT1/Tw6K6wwYZ/Z9pZyb73Rv7phJ89bavYMinGdTY42q8rUsyKEE2
QJ+1rVaZ7Tqy88x8/PTxuQS8x1wKvWTz49b3Y8uZTE+rnPp3gW2/klY3IcGQLLsoUcUjWZEVLhla
gyoVAE+rLIS9mAdutqVHj3CB/Kgv3pRTtNm6Zq9xttqTn50X+PRV17UkfS0FqGFSDjhKJP3bHqH4
Kb1zLPQVEpnWxX1gaM156uq7RyqNq27C/Yxar16MAeOcr+bu31i/74RW/lfGnxTTOd8yg0gcqOcb
gaWLCDtO8BykKiAiJeBYPw7eQpZFgGUZMdoBCujHmpQJTIynDQ8+IrEYZpz7c05iifH3b7RG8jqS
ESmCI4HZN9qfOozQuxeQdEL4o3cWD3537VHvzZQTksxMjUG/nX11JE1HFeL1Orx8AkmzWLmWLGnx
NzItFkKBGv7jkqjw9Xfy3Zo1us2Tg5ml3eIlBWfYDlTWrihTZ/rvsTNGURnzleCSHsW3wOm97E8r
Q6Fx4dt9QBy8hVvYLUvHwtG0D4/0/ZQt/QcmI10+CKA306OlbQNS13PXhCC+2/XR1mdgS4z1jvp+
KQ10qlFfqR7GNSD6ur24XIHgPGlpPImIH/uwSY31wg6YL2gzAdgH4i8PLPR8CvJ3y06FyCBU2hLz
C7p1sirVS0ElP0h72+8jTSOzF4QNKcXOrMlNfXTXRWNUky1duAmhNFPmO2MOpb9yw5hVAu5F4VZJ
2x9w3DsU6996tHmTTSpluMpz/ewZpJAZbiDSIIg99rfHzD7EZFsHtFDM1plO4QLri1V0g+fUiuI7
qjl+l8nXMUZb+OYExf2R/K7J+2+fWailqLVSF28zm8DrtCkhUSofzcvFCOxx+mVNB1H5Qk0yuHTt
pw+K0mKUE4OvtotDC3SXX9kKbOnZZPwpbRN3sX8DGgLInj3oFHWcGsyGrtb8k22FvPIZf70x8EE1
jizJOo1DZSBA7Rdk0GNyxuNpivSK3SorL5aw/C4Kp63wQr6fBzRH0/FYHjOJq9K+4Qe8AYNxkll8
gq9ljfOzPNGDrvHsK6+Xr/34ME9Yt67cESN16UfK9hu7EIt2yiCyqmIq+/xbLwV6MgPJOf5/7nQ3
ywuM47JGbTPqrCzRnpNQZBE1h1pktrR7iuPrsGaM7ZFg5837nrecuoVLNHBrSMDG/yj7z+0Lpc3w
DOnOSVtXsfsfggcKxizDIuGNUaWrFbp+EHJfHGLIEx3Gdh6ZLBqvDynWm7aChoPiZok7hn1Y+cpy
U0jND3yqMdI/UhljmGtUr/yrZxsXyPmpC566Q2OtPWiWbCWdijJQ56BNyHa+8UbFvwRL72wIRJrJ
yW3XrKpRnLzfnT+OBWJAWU0t7ntHYjDb6LEv04l9OaAa072i5ag2WQZLP7QOOGtn2ANPOrUJsRG9
fnStehVRTT7Kho6ykRqsJtwRd7wjtn36NvOSuCsEtcDEQ9wTFRtY2bkeU2Z9155ywCuFhyQK+mKz
EYoyaDjCxAdiDQgMBBthANzE6vxh1gYKLrzFyt6H0IUvQOPHrCUzDwMj1rsxPbBQQr5GaXxAPP4D
mJ7cyK06E7OCx16rXzUBlpH5umyafVbqLkas6+g2DU8kB3JXvu4/p2jUgEJHUiHBRBJ7GiCBLtS+
IQNW4wbTfWgP3TvaY2RAIH1xE56LTIOYhMB7gfbZvFQLA8INSI+hB+cxSILoKZMF5UlcfNssoGAV
344RISDmLMesrKSpqA+Dimf+1+AZPXrFG3JMf647HsMh4BHflvXGk8c+EBnhy978p98zNCXmyf4I
Mk8tGGvdRoN3H+funQ7cQumW8Nc8kDEG85SiselppXKE8uRIYqA1LafVVF6IyHyzgTW1E/65eiiD
ySWZhne/NbtWRoYsveKq+aSEA2BqRhiowFjtWKYI8jwdGHJcQYf43Kl1uQ2bIPBcdWAAm4z/PeHf
58H7G2wWIg0PpT2HyghUt/L87Mszv5a3m8ynviwCXyckmVvrSysWNtY5AqhC0Z1g2hgTIHpUg5mF
0qevmPCLCtbTW4SHgZHYYFYY52s7ndgy44s8uxBM/7kxZrBaGzerT99bizcZ+viLzZpx/bvr0oz6
vzTo++njWKvh1PvWTjDFmaPl9roVsXPZZAcsYC2ETaQhA3sCklD5JLD+6PNAPOfxqlXfSlbwRqAH
+YWoYPAswTyBnllQwwePKBBJXUAZLrbVi4AqWlCJljg7JIZZL0c2X7Q+6GChnFqbmWPKU8MNk6PW
+/6+khosFU3WyYKeTF0HdfGg80gmjVkleF2LnGwivqzpmpPNdgr1CIc2L4g/pfN/lVbojcfi8P1b
S64TPzJ/m3wVSVnXXHxLYgz3CtiiniAVBT2fZseGMYMVrmHwTFG9R5oaU+ArNk1fRTpzAN3sqw0g
001w21cgVQjL9cO6G5GXSumL4mjC4A9IdKR4JwcN8yCK+Yit7qWKFJJh1w/cY9zdmC5maxnBB22e
w140UtLE4i0XrcFS54VB2shvf733wYAzQ7LhzUlQ9m1rJSCqM1QF5OtbhElNeIclpo2KqFQyXwJ7
uyLtgLAk950jLx8j2/eZ4/+Wp+puTwymJQXIy/7CAnL95KIz7MfT3LdSiTMpQLHcVkq952G2x2E+
M6Lj73Pi9+gU176fUHwIE0ArrDOfMpoS5zPvYqw35Zp/rMM1TbR85RYvVHdAqJMJyBiNYLtP6pyc
fjJE8qnHJ6XA93qCv+gmavN37vA+4tVgm+FiMI1MeoT5VWWFtceHqgM0RDGolacjhRH/2VljTtCr
0mn1elkgQBWCIx8x+FdHt04CxK+7/2kAlV3xAWGr8s2pgdkKJbKhjWK8vOKKWZ+2SekSx9FsypKG
s9e6ht45jQzNjvgBgjvtbNMOK035MOq/dkTx90Hoqi5teR6mpASQjttdBViu7awp4DPk0j3jtlhV
Wa8ZzlqRo/6BmKy1rqmvzzVGNXJ25+5a1eOGyibdYGSnbQjR+fvS1tU4vW8mWPAs+1LAPek4PXZT
vPe/UIjNuy7G6dVw6KZDigJqLmn5yaaATSATAphc6geqa+Z8UEw1ROnsgb3Sun2HdNQZYjjH1lqP
Lty0kPItYyW5G5ZpBBximqhzKKqFdXK4xwEIcSrFsBD4sxp++32QLcg8ScsoD8qwk+MhIjpgLZb8
bat1YQmP8BpLPL9cfpGisEdEsQms7O3gC+WTIpaC2u8jufol+HQVxM/PtG/4eLpxsRAaLIjtOnyo
e7OZjknQkc0ovOgt0PcY3iQnjdw02eowyJL+99DmDqwPiWRz8A/VO8xzDyr4cijP4I5mc5S+w7j9
KLS8HgPvJ4UE15YQz9SvVuUAJ6RGaTvDGfCUgf/suB5Z3i01dQ7jkkiFR4JVfTIvwNlDhxhIXOn/
xNu81i0hng/gJjQcv1G7dGHSn5SfW1FKDs7Nm9y0/8ZufkqBrmDLuS0MpGk4Trw0krXLNqB5lyWq
MA3z0zZ/h6WJf11X/NY82c/UDiTHmxxonfO8561jCtavEvoqiPwxQrOOVLLxW/nbSG92IcHKVlDi
KK3thkgOFl2UlcwFOzBfc83c/rbxIsOb110OSMPAOO37FCJpDHbKbiRBxvYT8zSyZb+XArhO8fbn
y0i+h1nSnJj1uLfc2mgOEBarK3w1Zoefd5NyEUM7K2cBJzSbWvCJOxxLcSViyosmBqSfPUH2Ej+Z
zgGpmXzZKTmG03tVvnlkfC+6rOMBGRzxxuBhrOkEPYg3NmVQnpnDM9eX+Y/rcCpJelLzyjCG490B
Hp5rJGSP76hXlXDsP/bMv416hEl84+7JPo7cSoU5HE5abdo8YgR7HoFiKzNPCVaCLGz+JjR70rDj
AsO7mQLL7jZXUPdzjwC/HRB3Uf6aX4iDZVI3jXGJdKxpFEyds8VNWlmTOMftJrzEpP8yCo8/ZjG7
X2g1YdYfRdhBYkKkzbAN4OYvY074dHNex4lUaF5sPidvem/wTQtygDSeXpDv1TdFEboCEb+fiafO
j01tkD4wVJ1TgUlpwKTi/jxhx14jtHbijS5BhOZbABcxa2VBvHeYBPaNDmgx8XJAHNHFAF77FqwP
Sa3bZWZK3ocn9jtDVilXEc0Yib8hJUu/72ULH54/1t/OkUFIlWz++51Co0nTeZNF2f0GTMroqf9+
FY1grsarJc+nK3DACX3yt4z9vLJfGA+fx/4CxOTaCgRuBPQrRoUEdTLt8xf4MLQBccE0R6fmO54L
eQbgIJu/U3FJqZjEvmHNrispOy/P7+jp1nn1xDes15+wT0gOs9rwh2Hw+GvLi8Xc7IGyPOpTlSl5
98lCY6hvPt+hNKGS3V8xhv6DlRZv+rYKj2DDaNRuJ0QyFaTQdS/3lLUoJuNHrqj5BOi4GM6JoD5i
QVSXC9Df17sQfhNHAm+RphMIayf1aod8kISPBkE+ILu7ZvMJCRs2BUAntl8rWObsDD8xlumQ4SEM
V59Gwjd3z6lXAQkmPux6evOrSpIERin1YuDjpopIOGBwPYfTrP8LcPnOPHKnBBR2po1t45y8zXtK
hv5+c05EaCvwbjNUAGWGYOKhnxTF2d9pu8vkg7a0Ba0AnSv7vZEmoh4ulzYwyIJ8/td6UosDUg3n
pnaD+mh8ipY84+ayCzhbolFC+rEPNevwemaM0/UQlS2oYf9u7p9ucGyehD7JvX7NyudGPpkdZdga
E0vHbOmZNqKCLRNBXAmFgzQjldLpPcEUE2LyzHSZkCTtQ9v4IPv5zfkbHSQQ4kc7F20PIh50VQXr
oYZV8C5kS68GC5V5mSc4HQyjCZqg2VkVKa3KT+hyowqj7UuIcu+0ayLY/gv6j7rTu7BLtysvNnpU
jUK+Fttpt4uoFn7m5pncGylP2oLZo8YPqlxVe9A5DHWzeQw5FmoQZgE9noovU/CQAYEHTI04SVYC
YzTRuWlMweJ7wH3ZNdUvHoaxwYRxLuduG06KDMAo9b0h/S9u4JYEXRMpLa4AemUVNzfrr+Nm8pHr
EseSnyWVsbzq5MfQs2yL6PsnkH4gJJhYLJ6hpSo4UYf2n/lsPG+jdCDW0COD/xbZPl4+WCJwLuJo
Na9tdPYu8z+3mC1HMlAZ3HqK2xcM0UwhRddoTz0fhMTpU6vF+KEDN7NczNllRXd5dv+wpwJcGL8g
iH7FZIqAkmVM6IBLbcAh4kEKwZXr6efTkrVPn3H6mCjIIZcP639cIt6dt5121Tp2RqA4+at5BK84
UXbs/XxiwSv4QE7zpWGuwAY0fnQn/MMm9oryKtZ88TMOTdOoXNWA2e7T4FzMtQUZ7ciZtJ3ZZKHf
y0LuL05r/t0I+Px0rcXNZGyjjm3j9/jONfAxsg37lcCaWLqIRfPWjokm/fjutB9q35v2O1GPYmb6
WKBp5NWoCWlXyY+UTZgb/7xO6qoErnJQQBsQYSm7pKjwGqPBX7UnJ6QV4dTjnmYO/6zMFQh3gOcJ
6AllVv3rHaLk5j9vsa4Ox8AQpWcnhKxALEjevTjHyfHIcI+f1vFrgz3JmMYsjwVRmwGn2GAYjtUW
2C8Xeu4L+DEMeFKe71NcH9UB5XGHEVNZv4ZU32MGSadB0m/WFqMY1V/9SHjtuhExrzSUe1qsVkNg
wqh9ZHKIUV8/DEZ08MhzEaZ8S5jinMIOrb77cio3h06d1BuCMjmnKx01ZHa4lZgIZNQqU9BZQPKZ
T0HieRQ1NiPtfJEwJ3PWaz7a3oUgeRHSmf5bmlYtRBn7Nn5akoB8wjs4s4uRUA5IButLbuTFwO8k
pmiz1pkaNaKN8wrdaFbA0pm47aiimoIKspS/72qIsjMV6ckVJsFtHJVU68G9GOM45z7UiP4uikLW
M+F75kXXMjLk3ltvUIV+pOA0MTe1UuuWvooOg7ABN4OmiSCn6ojFgFHKkSev9VER6DGjhTXia+Fg
JWXFEA9KwNWPnsLx2kV6+/j8Uk7LWFyzxFWkDVDAP3M3SuweeXbJjSMOmceePdDY5PO4agb8BenW
BUJS/RHnUA3s/J5tU0u/z7+3t41aqILDtTTBzjxh+isW0U5GtXMA4jfsOhh/8Ad7d9AykkwSSMx1
39ADKK+idW0dGMk5zXgKGS2kqzDTvQYuFjHnuzxjRD230deelF6uR8TPAlILsbb5clTEoBZzh0WE
7DBi2vy1QAjuKFr+tVXmlnXPQEFCb/CruEO1TbRuWHx34gH+xXGPvK88IkNlCz7LtpQHXnSGpUkP
Ap5yU5jw6RsCrV0i048ZorGiK39jj2i3ss1bLZY1vvM2tibL+NPiqRyZv203iBpSMnxlm5R3WFwt
lZhWfhRDJ7j2G3CvjcEHLZGLiUPrDgCV8T/xtpJaoCEvP19TJA4SFsDEKBJoagGlPClm2dD9qPZV
sxaUFW7glRozme8EOKDZYuYzXMROFLcKsRr1Pyszpf1BMdII73UV5SU26JAhmOV0dEOIecSC6oMg
n0WYe7KQLiMGyG/k/q6Nz9hiI3Q6hgF530BQ57edKQf3MfLphp3lp5kJnpJMuQbQMj96Zy24xidr
L5XBSRKxkmKdEQgyj3RWTmWyhT3x6U+Bz1p3V95X+QuenlBNgyArvp0kMDkc5MdBHhuIgT0/6Kau
sSSkTQptRqZgWe0c7+u8jHq/zprUGRpDbM/+d9AV0itGV7qfb0CdB/FG26573pKQ+GNiwfZ1lNEK
tK4s2cQl4LRVsHNzQx9EmTaX4CtvhVjJdKWObRkZFwBbfr1nZqTEi4vQjfnzpt4Z4MBiJ6QSS+29
vK+0kUcunbKLzjEdWPPTndJ9RtaJigv3xSHWtNJZUjQxBPEDiqzslAQhE08hzgGl3sKZSpL1jSn9
wN+X4YFNg2xzPVqqhrfvJLIVvKRoN+Rkj+67z01R51dm7/axGk91xaiyGiSKuW06R7PmZ5bXBKNJ
UCLT2nJ6mzmmMJYr2ocYUUpVMng9IaDOtFOdW/+BovGrKjrMLL1JQoj14Zd+F1jvBi0PoOSCWM/2
s1tvmQf9TIPJYDu049TPfbNGNSnL2U7DRy0TgSlnLYhFPLSoOOo3IwZsTqWXUdcTrAqLhO/spkjF
72ORP+7h5hfWCslTpstw42vorMrY7IiI4SwWHOTVU3snEKkB86l1HnzpNc753RNjRh4Y6Hl0tMSN
SAQhP0zoM4bvGOAhs4sBNiPMznh7K5d2YO8VnpSTtii7vwD0ooVaX+aHNv1c8vb6DBrLr6AUAG0n
2nJg/TMb1HfYN6oEyocIUrUEg8mXZ5u2emxngK156p4UuCf9w823HQb1u9dMw8PZCX6LOibceD3M
YcGGs85sochgL13cnVxT0POdtfqnlJNUqGoIYuQnwo5rnWuFkCdQH20z7Q8QPUOac0aIB7+rRfXQ
AtSNhnZquLyo+HlVwmWjXxSle2EcJTsjznibcXJe4N/481ngKky/Ef44Fo7Tow2U1R5eH5TV0Q//
QGQktwqvyuxRBReObDOzAmhHOXyjTRvDnrhDbXhPrBi5KCitnRn5f1wcGYvtDfAq0qhGflKa4mNl
MQY4mdIOXun6N5sghnzGCcbjzHOMqNN9ttmttLGpYfmOxdXOiY8+Z/zDsWxIjISFRNJgO8bJvzvX
tbOnDmyhK7HgwBwOKb8kINrbm1+R5HQyYKRzf9DQIPIXWAAqK66oA+omRn+I6zbMisY30Q42Zm4p
LpVdvaxIIxt8Pa02xPYUFBDLljH4krNN0WOQhJeTBB2mJiw7rmz3BrJbMK2mkKIi8ducmNC8bbkh
SArQJCqTIV5iV/BTCDbR5jwBh2b3/tNQJCJEHdaZuw0TK5b0AbhmpE16VK7NRAcGKsndy34SyS8A
CANkBp775wbQ8PL6mFYCzNY8AVxxHcgDVWsygIXvKREvClKg7ZrVnG24dnyjpVN+CgiiGfwm/KEv
y6SlT+Rmss8DKYCpM8DeMyAMAYSgCS+G/L5CQ2+RQUT1U+sMn3rsaOxU66/CxNHdoVeXXqWGmQpq
e1JCR76O4N46TQHtaXTkQp9zmJGXYHEbyDPCuLnYbW585sncfyK5KEiGwlVUcWXbegEXRnBRAkxT
22UtKTfFo+5O3yz+adazloYQwl0IN8Ioj0bszm3VTJLQsSUZldxpt/mvZsN8S2NFHlN9SMjlaukh
TgaWJdmWUCfEQbDzMNdWoHCQfKG7YJc8B75+ky2CxMjTzOE+8vGrvoQ0XGs1to8myLbE5QoFRi1u
uhj2KahOcdhxevP3PlKDybv/sFGdr7vACut8SjtLzViADR7y+81CzicekQlSV0R5iZY15LEOMYOA
oz2SB/KzbvInsW/DSn3F2p/vj3zX++dND31RrUAcC3MgmltD4/2n1fLyjxpt25N4mg9zstYRQwyn
ERUYqGNIDWYb6IW0gs5lqvlj+0c0+SxGvQf646O9ie7TLv1QQhq42ENfay4//P3g4E6ARHJztJUb
SApzYb/8mcHsozoWwFGYVCD6gVz/K85jIochienchDvE2dk81Oa0eIqfra+LqaeeztmW3h7BX+6I
tdCt141PV9/vWgpA64l+qDyyl6lSiKB05DIEgT6MrN72oz7CwfJDNtTJ4WCV0aJb1V1X8pd+yKKB
pKK8TJZUcZ803ljGPQaxCrkIzlv6jrhyMqCecpFvD4I/C7snP/GO9Kn0esC8qRsC+1xq83Ph3ycI
DlCTD92ewYctj8VWID1fCLnVAmizMb3dmD5F3HmY9k/5G75oqaU9jhoz81QVuPuD2iV+inUmybR4
y04sVZvbH/crcFZEqv2p4/cM2QSnDAEVu1IQxP93YVcrRG2zfE3bFJapIzvXSEtNBugNAjQUrn4m
GwRuApuYttGfc57VWJF1P67Iw3+cTYx2Rh0XFNk/KoPCGHcOQxEm+Y0HLxxKoUs5DmwVv5z+5vPn
wXqi5QbVB28zdJg4UF2Kbkw7gvPEMiYsXTo91Y9gEG3L6IVSz+jCekYlVf2WxWFjULReKzVP3hqq
NCuwBF/BbN0UwQAyEmILR+gkVEFDROcYwQfYN44Meinx0N6D0gsx050150u0o/NRshvE/EkZyhNI
4ct98MVcqdXRd151XBvZLezQcr6VnoKLwVYKGEjI/fUbbvpFKjBZINIVE3une7T8oeEegHHFU+u7
RnS/d2ysQh7OU4F2CfENxv5fXB0BmCTOvFryrcF5UUtdXahuZeMruG6ABPNa0WFUizJ6B5QonjHa
0kfDv1TGSzIVC//ZFoEMMfO/kNdSJMXB2+X22z15i2kwFD4RzBNbrO8ua7KdATz2RW/JaxSkcSZ8
n1EpAjBHeyYmOqi2pIRaF3BK/MHizufCdyum98lvs53bLFq4SO6HVk8sei7WwYs+PvVNd/flfglG
fzhi9fW+66FMDPke7QI4vkOlBG+BBHh5d/d1ZSWwkNWcczaAxPnxrBfjWAgQF516B9Idx30T/ClG
a4ZQ5WuLM9q8PRf47/vdnESE0bA2RVCtQIWBDlWHApBT+WOUWWUSQTZ8hiE/HvKnqs0RK6ZmZYtW
p4qH67FlppL5I+pZBUj5PukykqnW0bnfrg5oMY8YJzGGq7X8KFZwsk0SbgbMCcBsFDjis1P8GBPh
4GKq19jzyoXnwFRgixoSBtR6J4kmC8lSfoKy78a6EkARpjfLATUDCri45g8X/fpAgfpjyMFeseg3
ieO9jAtSahpwlxK/xgF/aJzqrFPzrTLECjhjH2b681Qj5jRtdzwoVSx8geBdcxwAK/PX61K5Ieab
H7XKF2VbOqPBYkFA8zMbpN8wrsy8ZxoTDSocrhgqzTNkq47jvWaGXsbeCTwy5NFDAstdiRFwPY0z
4XREV8kc1hUTd8eZpk0MrTiIi5n+7mQk1XxG4AWo9XFo98wQPJlhYbZJXNE+SrXshW6/D4ADudCM
99NcDbcn9cIZamSD9sc+Gp1W8ZacIRHk7EUnN1MYW4MdDqzzFk7BGFT9+lmz5yiAAsjYGtq1T8lY
LbM4STBomVCWhh4yeYTL+j8k2xF66ntHQES/rBxtnoBCSCZjUvBphrGj4+HN818vPB/RXV2Ce9KH
JSDV0W2vvdgN3P2NN75xcuy1vc9i91MxPflbhEX6NoESau9C69ovnJvAXaNCOLDPwL+Kw1XpCLxy
cX5AOJGuXto2FWowHZbiZ44VinU4VOVpZiQkpn2p0vixQUOifYp8sWkPCKxri3Q6NnjxJIlyHaUg
T/BX533aDvP8HcaIj2PRuVGwLvEEauig39HP5fp8RFuIX4DmcC1DAJ4lzndAOGrE54tz+XWZnP+m
EqqnT9KkY5oqzbfiX3DZFL2lTx2seaG9admyNnIUGmRUWERAHR3h92XxlnTBHXSAu68zwf6hEtMC
kDxrmXxFr6MeKlaZMTxk6GRq49SFudd9bBOjBfk2/6AfsLh//yRkc2rmaFydLwihPNXlnyJv7VW8
79niI7Srs3DYaDPYQPPHZsKaZYhGllDHgL63I+G7P16XNS2qwhk2mzHzAL49HEhYZdz/8ruOk+Y4
FkkpnD6Yv5doKjOZOpTM2wxdJaGnalbplfQIdcrFZiCyZSeGHvcay+RfbcR5c9PH+e3fiHH8OqL4
qNscTBG7LRupkc5kEyZtLdb2EoacLVbY0QlrvBDterFOuHQ8u4gJ1RVDc1C4f8kmtk8hZMK08fnU
T+WuxdTqV5d6K01GYA5wmYxp+XRP0JX491eJ6im3tkOAc75MPgK+macJwy9G26G2WHseizVxP0IK
R0aEdgt7d9e9HfsNNLdZqzmZHz72wBSBi0L+Wt320SonnVwbrfb36UroFosZUPAjNOovL2ahtg2u
Ia+XYRnNP3mF8SpB7dk65gFub2kUe2dpQS54PR/MvKxs/YSgeMFsF68aPUi75jbvZWYVUZ+TRd61
r6vQaD3opmHRD3l+sBUaEuhTta3tJCxBxY6PMjgb8oZ6zxlvvRWj2YUXpX+E3JxjRktev8ncPGtf
BhxCX03tF7iT5Kf+z9yfSe+YGUxum/tA+LksX0NFo1bdrcVuXWfoHYi1JYeq5DBhMfSyQXd/5NFR
73/1R+0DX7++8qJa+VBK2KA+C4nFQksZ7Md3Y6HnutgtZe54rJhG/51ZStdAkSAiwrLBA4uDeScW
PNb56ypJWPJSiuPZmXC5fSG4hIe2Mr5hx0djAeWFLfx9Slr2L6EQ6TxFR9zeQdJy25mFuId9N57+
xN9FCMZJmNXDZCx2T5CN3mR+MPhDGgrok+8ks4pn14g+z8w6Mvuso5FQGdMHiIeh79JKQ2VWowPh
J9sGyFSGnFVlIUIQSl1PDQEF/MgEQ9zb1c5aKhhIfYtatdKl/meHv/6n4pGg+0lakSHi1fu/y84L
hg/xABp4hpNgMZjf3hHbt39607AcGPQySEKz1CQIIp/F60g0MFAoKSSwOIdxoxcEY2K0MXK7z02X
cB1x1OzgSbquF4fQRrv5DGP6VGK9ErnYH7lV8IX+BngiWJ+HzyxPsD1unxt1QxQP7pPIxcq04fYS
Z8tGTYmwI7qD5P7i5qKYExRSiOKKpRDp/pSMakW3SPg9OG8TSdlxddZlEJp+g1F1glV4nsHFxMgf
W707qs50pV6cnndt7bFQCpfIyzPYka8VEEuLWECk4R2ZMeupPD9xY5WdEWy1Ej8BHMHBGQCpTndj
Ip557MmqSGbkIcBmJVbuqCNlp4cIOkXLC1SWGP77xPzhpzWEuaUq0zu4/S6XQSBRRSyoKCtI10MJ
Y4PxL+WcYzFp7BlZMA1ZtNKu9qN9QId1UCrxZ2/YDkVFCKNOyCCMle6kstrle6tZVI3hWpUFqTHa
5v+WZShA2tS/HF061QnK7OdKa5+JRMBHiaIjsaZbFIOLfxfWnTK+rmUomi0EqC/MbbNyCi4SvG6A
O7rDNLwqBS38Z57q5bMK7vYP6CfrIYm+tJqEF3wBO0Ukd3SMa+RaUQ3WAL9Jw9WQB4ppSNcEPoXj
Nv6+99DIL74kkm5SoXblp+sbaNXyHlEQyHjW0yskYBQgJVb9HZu9olVM18ou18Nc+9vNeuk2d3eS
cWjRE6nxrHtqkkAzGXGmIJtKHEAzBAGxxOpOecMSfgEOmeZsNbbnYupaMqZ7rkcXYt9b8xcMGO6V
qdthZZQAkRd9QWYt90FArFUGgB3DntIu86LXinEp04sFKTy3qYvbxxp3qNsX/Kp6QbraaWD//NQ5
UMgZfByOyGlB+yiTaEAeN4BtcIdfpwQ0eM1F5QoWbLkiwB1oOcaI0rZGQ6mhc2oDc5LzSf7bWk8p
chb+CdwkLg8gZiQDHRfO1TxXZBBlSG/At/hoE+qZffiR0t5KMTvkhK0z82gbbla9xOgCJ9Kpm5Iv
4MWIDSQepGPknnmmeTGnAU1P9S7VV3693jB7oyVHDshjw0Q1KEcEg9Q1Xi8BUVbCnLxfraLXKYI1
M+mpDn5z33zcj+nV60WolU4Gee0MkaDCE9GQ1XPzXeroceocr8nzra/UO/Sz93auj48RuBbVrg25
gxW3wGUIFgo9c+uiNiz1cJj5ev8utU6tq0ece06PiQIteHgYzuzwNXAO2v6ON2ODBTgvodDS9oeC
6YXposDuN25k9NZ1ATtGV+1zGlKusQA+nkApvRmEP8YOotKBG7GldopiLBQFh2W4/q9gLsxwd4mW
GVz1XNIAcqlBCpw8u2weSVwW/1Avt1VyT2Y2YL3oY8Y22Gj4yLI6PHrZ+OfouU37xGB7PqogsGRT
FqD3pj5B1WCNjYu7mtcTq2zbiXIoHMmAu+CmtwznLUTqCJA4qAyQkWnTpB6GBcvj1A3gqGhzsYCf
PQ1nAGJvnuc81V735d6rtTBvlIU5GYiLTHgI4yuoGtR3bby8kdSJ019AK0fLAFV8kt1T5fkbp0Pm
/DsduGZ3iAEwmH9gRTUPVd28L4aB+dh6dDvDn2OIi+tPbocJfcLBwGDZkXrkwQE2/jV56OGuzX6q
saKPwvc1P7YLSusdukplfh/fAvWNDIq5U4qTGXm8nmWhdbjQNfe2qGLzQFPqmjp2d82YlQqoDQtZ
ntDLhIIMJKs+cJ7okWlkWzm7Dq7bY5s16+g5Kgzpb26k6CiXcVv3Qc4x+ST11MaDMajZekgAlp4C
rkuFTeFKNlVl0QarZCbvvJrl0Ez7fIflYkMjBeEaQiFN1/c8XMNA6pogcCPDA9vVG3Tjg/nv69eE
izqMorAZkAufxNZQX+BNvb4UPXdBTWNYx5cHcnxxEzTDgtCJ32SMlV8ZCw8XdLmKSBUrlr4OtVBT
K0yTk57BHXH3adl8xc2b6wTvlfA3FLBtvjfi8TG8hoOIVRckKmV6zyR8JL6L5DleHrBoWuSvABvQ
ZrCn2ikAvlQCTRGlPDVE/0EK9yfV+pEPQCnzmaX9VYiXJ0f4nm32gcqozNrvd17Y0cVylXAGKQDe
ljUatkEvgZ3cqehUFRa76KKS1YW6nXhww8hO70glA+O6L9jFXaIuUDngwXPMMemlwlwnH3emRNZo
ijdXX+SZpiFlNHFxR8NqgwQEq2X8ldPg1gu3z7sp5UUNmN8xcFUB5m4wFJ77ayjp8RM5ffEQnISi
E2FjQVwMpfUXKOAwkqnRvxrr81Ao1qWloPz/8EDc1eOvJ8IGm32i/6AcwQrv9ygypvmP0wVvrvMq
sNGJ1mDqqfhOb0Z987TrbPzxfxw+sIWjTBQMJ/HUln5XKtbQkPi4K8HOCKbyqZX8/AurBStsoNXM
NSd9AEIPMWb0BGF/aKvyBmNCZh8trrU3Y7CdCHGEPYlVDM9rt1bsNz4yJFsQRuZYV/A6fuU4vCpi
7B+pTMeZdc3EcQDwCyKLmHEUwckMSsoin0OXKcKOqNHCXDfY/B7D2QoZNvZs6+L6DJp2mf5guAz3
sBtqtN0mX/qlzgQGBU5cWAfFJAjrx+n46wMUAiyWswfAg/LK82HeyDgddd6ejmEhhN4KoPIUNeTW
63+XeO2yRvU99ljP44sx+xrXU1rTsCifyQMoPZf/PHdBZqGp5ubNbz4zHGhGjPmuJhxlh1a3jRNQ
QY0xx1vXAVjUJjHRvZVPaTZ3th9mFFo4D5gpc7M6imbFs1Zxq9bEJlrTPmV2l2IFgNyqR6/hIHK1
iDQQUxorm5cTaOyHKfXqeRA+umW4jXKJ8FBbC14v7xaEwankPXCBTRbCmAOLauwEcqyQEG95m8zK
gIg/AvQxiD7PeVARwlanHvHhWtQaYx82PSn4uxLjcgUWZEi2UpVxcCl5DDqJRz/WeW08uyEdjkUw
VnRj4lgjDek7xQVot4r0IvFfnF8vLksJlTbLEi7Fr6BzQvGHUs+LyfI6XhS4PgkWzX8lxhJ3T2h3
YMr6ArH5AwOA4hnlnr9LVlF8i03yQlCPoz4YyyiRiidEYRsL8HzYxaUbSbzjqIFc0xSHBdvIZHrv
rJ5I3MNxis4nwasi3PqQPuYhKk/Utyd9HihpKCgvoV4RiyYkLV6JlBqhpNpHttQELQZZFVEUVEuB
BaT2MUVtXFylt6womyfzqN2Vr9M1U5EbcO+SYb1/eVobxvxqbONDYR1tc0rLce323kRQkwG5lqJ0
Eg3tKK21tO6vWd+y9XEAUD6Np8iu/g/LJuNsaX7EYn8PXnuP7DOXAxYJvcMhBIpPhp3SUXQD4KZK
9QCAaSm7LiSpCcGRpmfxHKaUjUQqmF6D6PQhCPW6m1ccoevB7gr1+bPT/koqRxgarC1wHXJvJ/LI
Lg4DQikMv7VTGWHz044TPLJ6EFt189UwOjgkFFZTWET1r7G7x0SAlh/MotD1iHLiXX5sGwBux8J7
zZwTfwxTQT3/sDBKlPNR0NEPkIxUt9J9jlcehEhwFEKZx7+2Tqku0KCOZ04BAdAysCTfZ/zlp1JW
tG30rMsl5EnSofB1YBYI+3OzxQ6YPHl+sm+dgcbA7GqmX/5muPyjatxQG1SDgiBQNUSTFPr94dc5
SeLlYu/9EWJBCWf/Qnkk29VFHSEiQhlodykJkjQfqBKAtX9ZxyeSGtV6+e2OyENyv9fH9d+bXmUr
D/EcLm8/JcG72MHfJX25Bq5x/imYIPkdC5YECrnqXuq9MHHar5Fa+9RljWhXrRXubA8/sDwAMs4l
chxuMU8qYAzikKq+jf4j7neGwUaOpTnO4t/927cNrnyVIaEfCURKxeZ2I5HRy2/21D9QW+zJbQsM
g0nUxD8fLarisLFoHes1MMi7aG5azWapMxK3W381SKmLxmfjy+tYxeNqPYYq7C3kXDGWe1xt9P41
xyYpIhTpgT0+k6KzKoRoj/KKMEnnh+MwkGrJucvAn9gWfzDl+yUTUh5wIPv09sN6tquai/eZiiDs
sMSUdU1cMQw7OeYlB+Xqx8B/1bIP22BLiFM0UFDEzrZ9i0VSEdv8QIDR01WwuzjO0NYUfL0QlPCH
XrRcfveERauqz4+2rPGUYtniPeRhDhVzjhQhFQIgdcE7APwRRvt3vC4LTztSHpNZ98031QLU13KA
Ry1dRnF9wbMQH5imnhdei2z9h/bP3WGMNl+KWEvnPetCq0PHxLnab3GhXrChP+idI71AHoVyQPNg
zloTNtD8hkA2B+77AnftIJ9M3iduNO29vTdJV3RnnHMLebPIpJS3ReStFHQJa0ZMokupGl3l3a/U
UOkYSD6Jq0lou//jqgGP8ggXhblYS9N7CgIUax1ugWxGjOtNWM98s0NB9wCwkEQeN94FOh28R5QW
8eDkjRzcDYgwc3K8p0oVgWsASLMGTM804IiYERtbLVRjfpZjKCCf0URCCPioyXTLzZJtC/nUxQnq
Uf88EbtEG/cO7+YoyaAeIp5yKIFvg/2TA33F+kX76himUF2THU0iSF6IEfo9YJfXK/XQeqSCn+/j
SyhSN5EmmSGoKd6ZDSaaWhhGmeTqE3yz/fcEijolsaqhagkhTHXYHBl0AYKzqBdggJMZlKhlnT2G
gkGHwayuaAncNLYYtaqfASJ+tGPbWEfhmT3ckZnBLRd5cWQWU9giQTmF0EXapf3apALszJ5M1laT
BFVW2fxwHL4hNRLYu5KlXxVrB+zWKlPPSIbGuLHg+WLywsFAVmxg+NOaA/DXUcBSjwENxK4MOUbx
DgAp6EERT8Ma4k2NAzZx2jFoEbPqKzzWoYwHY6XPJUcNEnM3J4nadTixsd/1L/CELqUs7WiICGvn
8BzDaYfHzq/hCurW7xydhHHqbWbBd9veefR/6LSKHtW3/oC/7yMK7L0cEG88JTwVW+eRsssWu97I
NZEHVH/tBh8YIDpjHpqTSLj+tRawN/wgJSO0sHzT/bv/a/zRM9pOXbURLoHWzUeJjHhwz8UMk0Ji
QO1pfPrl2x2jrN865WLjdtTG4oHTuhPqQ7CTO1aVW/c3RIj2WOoVehN4i2C0TWBR3ykZiB9HRrMR
WsKmfWQcR3vBNxaau6/Vh/sumeXRhHgJ9LvWAeoD8uDlX4fCwPBVDNQWEPVQRWjwipCXNqxA009P
q+73zeM03bEbWEyWGjTwFk/YkmDs1NJ68kYuvJNvm2MiyPHZ5fi/vG9Woar6uX7cQSwsHKwvPsHl
yNDV0j4lRS5UwJaZP/0sQaeDSPtk2kKd8UAiHWeT2TnypoSmc6RDbHKiRhLVYPTR9deFeFuC5aoL
e3ooMLmFf8/LoECUjjej95gDURo4F5cyu1c0BA6vPCmFj/V5mVzYxzcCiQMKKn/6wkoJ8dAGwz5R
heBYZElzMtFNo4BcOZdIGpdnWJJBZ8XvXQf3Klkiwr0ABL9yZaT/5r5X7iYwKqDT9Zv7c9/+++S5
43XxmAdM5oULmgDES2nmxx2GGCesA45gWMmJJBEija30unNgLgO9k1iTNS8eAV1G4HjqawwqQNY+
JuIPPCYWsI/4CotUfx+CzUGh9GLjx8EWVPi8valC/qjjNLWY5XdDWt0Bh8qphoQc3UiFWfGDzQHk
VvKsSrgowFqc9MQflZbTFLDu9M1ACoKFAILUrF90VKnE1VciePTL5LAeiLS1H9J4CkkTGFRLPMTQ
gvGXOcI1UCypHVHPVv/d8UWADQWA3lB7570tVrDce9I3MpKcNTm04qR9QN5fzPvQJUM0wAlnxurL
+WKEt61ke4EMSmPjF4b5E/JlJArRoHAG6VqvSdWgrAHmEwfy3UqgcnAjoqxZA+ZOB0+o0oESliN6
zBp8ufxL5jnKsBWLWq0gQ8mnA0495kKY+ybdXsGCugrImYrdbQapqDOyQAXGJf+ooVt9btPjiqGP
IIqChYENdCjwbSvyfOj3+nS7ENNRui9RbqRHAIVjabKrBxLJv/pfMEufFIjw7fSfb4oHpPptwUHr
odaJkb98vY1Q90ptkcm/gEy2ukAu1AgYUyea3oiZLEMJ8xwZxjJFmTvMQTgT1PerbmC3iHRzuJyi
JLteYam28ts6J545qMHMq232IBUht55vQovehkv30s5L2b2M5T8YNd3ZzKAJc9VG/9utDXO8CU2q
+3kl0qn6Ul8jgTBhf4LGn3kaYTkehXgLfzu+yNKq326lshxZGxiFijgFf/mtDp+0EnPRabg8Btus
AGXNavG0+f0MOijn5lNN7Krd3uMHgOeXuy2o6oQR1uOiGo12FR8ELx9Dd1CzElf3Xa4cRVdBNVNw
/x8l6Y73xAyd73sKRYPCg0S0nI6PQ9ItntN9LuboNpPC7ZsNvnCIsXkQ1egSjSWMYzHXkfUTrkZL
4nTOGou3Jj7qt5tzcOzu95maCw4/bXG62Okq7joNexzwtevzDjSBgyIuYWPxXXyEatLwO7BmiJvG
DOFsVe845hdFFPc4CXQonB2PuD2aztAhrCYO898jiRfyjyvrDwU0ezVK8ENB+aTLPe4PO0AudHpS
+bChCJ3Q6Wzmz/I/wUUvmpUmL3waz2VaFVx8xLdI72sg9bdlyspF/x8QL1uEO3eI7Y0ujLEDLShx
vviJSs47v0+MYoeznWMN9OoH5LOFEbrNtmhF8mtmGUAy/d7bPPcCVA0wx0+TAP2M2xMF56jAAFgh
Iva8cYKVLWYl4H5QOOuxebQDm2oUbIClyKdkuVXWTmKf+UmXyVGd8ppHxq0s4h/zmxEmhCELnAQ0
8vTe35yLzSgvQhAGa7xzPxcY3dKJhQGx26oVXtC7D5WcmrSHOxzXd2RHQ553r65JL5PJe1gn2RWn
1IqBqnY/HNkM8VXZyXEoLc1RP6wzRHQTWSBgEGHk8gFcs81WDgf193xp3EXP+p65YDS+WGcrtBtZ
/cL0gYVRo3CqU1gsa4R/ZD3Ogc3Rdqjqoe+ENQhrjKpqh14YAYGZ3AMnTjmKmAo2gOoEowfHYwYJ
BXAdgIJKJ+amXfryQr+e1Kxw6p/juQSUu9EMMPprRVC28szPuUwi2CU9H7Dfnp0NSj5lYFegL/le
6yVBHNXYsp6xE9lTXY50umvDUloeKZ28yceXBd61Y0RDC0Rjtoz++8aRgE0YjHejP2pIRYh5Ryat
U16VuY4lGtICxRfhvaYmjcGCqrVKXbniixnjccsY1W7bhVtbDw8aEERCX1H/We2L9I/oUwFOjWTZ
wHMQI2GFewdcSPXsgpFZx74rIqIIsObEOBhs2wfgHa6TZ1eaujOs23z5+dlflFVjo/LiPU3B8E6q
WVyTTRvq8xE9cLM1W6jOVDp52B06qpbhZH+h5ljPcJcfRRgl0dUzLOmyC4jMTKBNMPm8I7uEQKvL
n1VsJxEBEbGLbeBV2qjM4Y83lLkHK3TXr6CUMcDc+l5TQLsNTiOyALn5WLfhUVQvLMWGaQvMYMHY
ZRSdkLMD4YH0nMN8m+rAvpclsMntuMLhCX4t21HxfByr/Kam/D6bOx2NnB/uypjcyStnmfLpuRnY
V9oEuUPWFMiv/coyDmxR2ZWli1bRDnyzPrBLSfGotSu6JpbsG7NLAjawJuVw5hH/U4NlFU8iR682
VjlElsKsimpVNAyDyI8uWbaO8BuWXsBrbkpEtOyQNsFOoA7yx7F/OL7x+x6/bkpctdK/ChzRqoPM
7vU8Vey+tw42I005bVqstKxpP5CV855jrrItN5gG8HV3y+U888mVtCLPbnZYXY7yRhwC2KSFF8NA
nkE9Aibihvy38oW3ic0ehUx+dATnL2bDtcitfDU3iNN7P6Gchn5LzHSqk2LZ/OFyJN/Z90QgeQou
CibgMMujY557jqXesXw9yk42GZPGTEohzRw4tcoLMDR19tZz5RSNrul7YKdvVXkkRBVyd73CEuCM
oO8+yn6DP+A+qAE1CQ2zdxgfBuF7HU8HYr3fAhbYhEoR5b0/nxSMG3kgyz6EFtYCtJZgzCeLSu3U
XV3XMsKrGT5yPQNXPsLnmDKOBNnf9LkYManWxbcc5ebuwehCNNsx8baL7YfHuSpK1lAoKaWf/Fdh
zGUdhIpxayDRYs+/pfmYk15R4WRNIc7F04eUjQjgr1DP121KTQ7BBlRiKYuoCc9MM4My7nFtXu0v
ldrXiugQwak8psStcW/Yeub07Hbug8sqfi8r2GvZOYD8JzQX5vk1lijJr76/dlL0A+QTMKFdlXEs
YZJ0Ilz6ryTHvY8JioRA9apQ/G1GrYE3I/0s4AOWJVZ5XTGAPpOnAbJBQZQ347NqgecXvQYaTU6V
QaIDgOcD9YJeWGk8efS2IvPgfEFrtc0/jdlfmunGqICISEqWmD/2w/5kB2LK8FN2xiP2WfDC8WKO
6LPmsZv/PLtBP2AjNhjwmYAibhe1cEUNZ3gFT2+NR/vddoSkBrnc3q+z3it26NYRG2BtIMtMYNEf
A35msqxxhzVeRimL6GRyZN7/rKpYatV80YBFA+DejhWd3jWFyjaRTgiErWFyWxzbzPooNsEhTFPn
LhVnxK2JztJynwD3vjXtseurID0c+SqnrvnQgIrF0AMPDnoy8EQP8dYAVjh4F2mremrtYKp+DYvC
xafAQP3X3MEM0Cq+St0CMOBfpUzju+fzO91ISSFG3YXRjpYu+6a2pEQ7Drmbw5g83pfXrIi5Ewqy
T4pieYfb0bF5MefdmS1qWlj8TQjNzBpzkwp38UISo3i1o/x9fSk9VOxvaWmOW2jym8eUk9KfKMWJ
5Q1EMotYXlbKJuiBAw0mNvzHhCkd4KNtVloq2H+jcb77R41XpQNNMScR/Ro+lmKtiza5yvzjxpyh
d3l/loIywGc16a4n7qYduMVWgQG7pzqgPc5CpM+ZAG0vclv0e37s5kUxESRFxF4rCR2j65nPGrAV
WH2N9KQioVSsakz4uR5AZXnSqxheyvc1Wy690+If1FJSjSZx8/3mqsyfwFnORVVYDnkEDlR564uk
0o+U3SNb9AbWw1wMy0QIrwVPl7XMjjyAqjwiA8pSCxjF60mnoZ2qLrh78/Mwrxf6IBTLp+G/E0lv
blLDdHFPl6W86kPFO2D/tEckhpF0iTvXnfNAlgHJpMDXzOB+DRsZluElOhIKAs5GYnkQfbCRPLbN
oUxDsg2SH1sz3oo2hFax6R8mHWCjIr+1mw9+ga5pUh7Sdu//rTXX1OO2W6z30fts4pM34B/4rjUM
uKhEcHm+SkRMCzaqriteBuwU5YhTldk1/QR/NwGRXUGIlSH2lDvqj/KZrf5vmLAW1bqc98dxKfPa
hIhN5/vAU/3UxvmQyCGje6fwlzB29rGHXk9zYlL32qqeSXr5+WLNPRyJtxdqdSUSJDsUCmVI+mMl
3W4HGz/M1mYKYk5FFZJDeLLVRjG97CRhjN1HzeStW9MmrvZKeBhncUW8XXAALvh3h4Oi0e71lDix
WDwur6QzhT/PQBctkH1+lipPnciYySSe6acla3lqyNt3RBsMvB0ssfrrkJsHnCAH0O6Dhp2b9wp8
sIxfIOn47/KtHXFa3NFtg1rOao7uU5/OoVswBbWTpddFlob/SUHhwOC56V6FrPYDYX8QwyUa+699
UHfTC5wpp4oC4C9UtI5dr8vAE1j663ufoEqK6Fj1ZOtw6CB0g5YliaizMnAiMYCLJiFVCEksev/n
zNGAk+h8b71/VIvHrDNQ9Yj/I/bUnI3C8/Dzkk5z8c7lmRMzdKnjrNbzISzOu74lJavqZJLmk6ZI
4jAVmjuWvcp7jaCM7s7/UA6mTC1LYOHEK+ums6Ld6JedVvKaPPROT4IegOd/f1hYnqvXBnQ/tsp6
PqUJTO9ZCoU71wfkHu5hvWhnFW0GzdsomfeMPjtrBnED4/oD02dhYEXzRyk7imEiefW73JGxNLmt
dWiC9LKvW79yFc1TV3VWnbc+hnzDeSbDALgv064VKPNjc8cH33dDhYJ+4vylw5rWviWHUKjkoA2L
lKE0uOV+hU8qOM1Ch5Tkk226i8ZESqdv12OTT3/2AR+ka1EabCYZdMor0Np+BS5oC7hUo9rsbP40
kdWJgqgt/3JCH5pMg/WKiaN8ShfV9/2TwTduIN5SYIhkrOuB/34/fk/1ZSiUzQxGh1mHksO4rxdb
lsdncOUF+Ij574Obi0rsD7ceyGcf6RZpNeY1ZOAPHj28R/i4B7CYdiHl5JqnZzqsXu5GaVGTifMO
DOGONRnrJzg7NErFjKM5JREO9Pujli5qyB3U8+VN0TbnWRBkrWyjCqDs4MS+Ihhcb56HTsiXrze+
VuU42mf3xg9lf316KLVHVXzGg9EH5JA+i/XsrwDZ51uKETCF+kh4O22BhFdMjAW6QH+gg8NM5Fk4
sq42mxuNDo9u1FLkRLcqfq0/NLxNOrhMs1OtQQ7+ZUPsYRFHND/9f09TCSMbfRiN9QvuMnPp2jfd
BpNAmS6OwbcyS6GlHBRoVMZaWhHmllE1rRunpTGQYYpG0lrT4bPI2+QlMnLSrxp+SsJYKbBCCRlq
NNvptOzw+5X6mwNLtpefg+ZdR/bwOlZgV2syYin3eckQj48BjWHwvkUNhI8xYAqM52VYzu9rMyS3
F3lUEdksykS0SYRY6J8ajYxSplIqwOmmc8ylb07HAxJEMkJ/OYYtOX/cT/Efu+rHzwIoJY2SzBzL
7/ArqHXGrXUwi59wO69rxj3syhmflu7EUc6Mhmp/hCM3TOZ8Wz4hVWU5brl5bE/C/BSG1oYrpXQa
osDUb1g9l/W2p6Lo/POR6oQY9s+aNOqIIo/fyQypW/8Rav52CKXv0dCmCEOyQNXeB7eN1ZfiTrCq
DOMtMNLDqo2Hno4Ch2bK8sEjkZ4HOHkwKJtEau9aFsyYceVMgSaPm+TbCv7yV58f445TQDEKY/m0
Iu4VwpwibQuLgGlpxEjYE03tHQhQmvDFPZvARVR3bx9UivG7MAxpB6kCNQaaWw427dGoji9ENVLA
K/MHpQ0pbZjRX5i/UGqnDMPf0WEAKOHrGSX/Qy50+6txpJS04ZsxNJuXtund/C3S5LBcTKgK65qC
qUpDraK/wK7LRCKKDrzpOuGvMUn3hh/CtXP3y5++44SMGDVd9/Dp6apJhOy38uPFlX/QW6Aztj8L
wEpveaRSU+PKoQyFO1S3mFLZlz8lUL7LXausHoIAICztuZ+ZEVsoIlhsAub4m8MMOuclMwBelVuq
hybeC246A6Qd9Ar9la9EVf/I+ukMuda7nzHEiTZ6FeK3sAF9/LzCOREM+Ry1KuwS7T9to0ojTm+I
Qdo2b3yovfH6HPoNs4Ip2Zs33GhaAuTBDOY6uaR9XkStIIsOWhVcXsMMswEofOxh6Ib7jH12r6oN
nRrxETWucZChntio1WtSSbbqxC3FKdTGcqTLxWslyIfD0q3iLI8p64Z4SqR6LV8C8aGUHKmseoi4
yUKqgf7MtQa/m+nCTIfvIQ++rOAXsJl1svXGzBIyfI3/6PI9wXlCZkqh3du4jPydvqr2PWqPGJ7B
4YxOg+KIIVEmG37KwuqCrStfHEGB+xPfKqIf700GUGj8SnxtGGgKUg5jP3lhCBhcShtKhRLOba7j
3/hfgqwl0V4SGFL2SDg7TwsMlcRt/3hC3kgelqEF2nrqaOkUnWfjoMvshyMDWaw+AktgeIfe5xge
PcygBxT6OzXVSUbsLtGp8ArJuWHCePVHe2qDJIpr6ZOkaGct09xpdC4XIxz4St8NIuo3NHSuUEJd
2HS3+Dsf2l5Lhdjh+Zh0hY2eX+MzDgv7pBbQfvVyNxkweEsIKNK5+q2LcBplflsz6pOnYWTiZ3CV
+lVEybDCQ3ljZM0rxL4w1Cxm3PnSSWqPzWZPaTB8JzA9BPg/1mVxNRAqB11zoEGtPrFhHzRicTfH
ksdIPXiHh6l/QzhS/lHCp+p+YHvRisB+x/77mQDgd44cl+AGCn1G9comknwXEjI4uDTaAweWBvfn
nNu4K250qu+Ov8VOBkCe8Ln/Cqd7mQ53VfXuyWgkVYm2cd4L+BUr8Kx+IrGwW+eNrrLuUzQepdmy
9S2OkCeTnZ/9QhVTzCKQ6F4r7AI4Iv5hf6W1KCsNbg64bPSWgxKzzyj+lvFs3nmL2T3pdABgHAz/
rfzJ3CJcRL2aD2hxt/tGUZELD5V/D4GMTwXhfC29weSPKllGDvgCOaNCj6iOzuDFGRoEEPzjNC48
pReJ4tt5VwPv+0nhVLFW/bcB1kgZH1yUthUpVGW8R9prTZU/57jArUlw/Xq9VwxD/j+05bctJmmx
BNcDobSWNLIvubUODZ4ybEIPUrJ0ceLAmBQz6y4gQwr/3IroX20kQU54rByu5/7s8MWV/bNt++Be
ERTWW3ckKtKT6JJ83S2BNfq/ybA9PgAb+wXMLHLmqI1wKFXZJJUbTfonT3jxxC3X6otPnJ7Y/t8f
yBZylw/FFWxq3pc+A6Z0iB4JmlboOmt6o2rqXDhA05lGavjbpKuQaso5cEeSFbd8t06JvvjSi0CQ
cBdA48sKPKExIIhRSvDUVsauR2QxNEKF0vZfoKQgryYy9FREcCYzAc3N7doFn3v3DFvrsmQFFsGy
msARs5D5aYhn4HLC9QtNq0K6G6HF8ydTn2w89RDUeunjKhxeEV8qaHKwx3h1t5bNiSAZvrAH9/en
3U45hxqQRBzr49/HdIGggNj+cqWdsZLdF/5cg1HyYALvIXrakZupxm6iUEvp4cBb7ROAib16OxSH
IthTUmRHx5HuL2F83uAtT2gmz4c4f1uTv36DvBEtGjkrAXp3ZmAwIRo/xkNYRNQBionhAYpYsdYL
PZyhY0+JhAOmRPHmL7HptOKynDG/lPYg+T/ptK4rggtAihhQaUC9oXEmKaCMzu2+7s02tuZx0B0H
o+DinY+lsE01I/dsbh8w48nJzsbGZ6QZ3qJfFCR/Lt1Tr6dZSISLSGGHLtxtJyBj8iQYExWxrkcy
C4BGym9FXLyHTk8zZMrJh1cN266tbvIZcoaeg9mOe5G/5Q84F1FyErbtXEXplTES2zBqQthFi539
CZpYIFW0DK+gER0I29xi8dWWY8CiEvcw3vbkEjSoxNl22k3Oerzhx6x3SFXQzMXPYR/2XCRytLtc
YRo17Wg83giYmimEYqRk9gfnX+HtC8Yb/gNfDv1oNygxyQbd9CQlhI4inqsy+bKm32podq+on272
5FgpTecgr8QxNgnIKyfk3SG9CHCULMZgwO2+vWA2l7ks2h2UgTebDU0e6tNLvcK09MknaMEKXSEN
UcVO6nafGVzGVfdlbC1z7nD2UJgAh5eRPx+JhItXi3vGg4YcCyl/3wbMeEIpaQPwWyArIe5qui5I
KovzsUF+J+Gr1I3EfOn2rO6l+KNkZCXepP+Kuzdd8lcJj59jiddAKKRD0irv6qcOn2zXP5wCtWg6
q3PprvXad+2TS6m66dA3UbSAHawowapfL68U2FJBzIJKQJPdTuwpeFRzocUiAXJ6XjfjtUZlRPu7
430HHzzoigFq1Td2Gm+HLpIRe5fmo/aRJlpGJ4OOFk/iX9VC8Or1etNtXxjvFU2a2pxL1N67f/YK
4+nlRG/f47+dTYGd2k4wZbQoIDHLqzZvDgaiBz48oX04SAMHGEQCoteNiszFNGGm6BHHvM5EEWTQ
UNE13Lbm2m0+2TkVywociiSui0rr9VVZgB4sUXrfO2EW92bYh+o6K3rU4HM8y/o3BQSbdcMKwfr3
TnodSdHrXnNIQIDR2lNzBKWzBBe174zCbgurnBCNBp4BWRg7q4tEyX5JOR5pmRdaj8ODlgQ91aT+
cfhRrArPVwlSsDvuy1RisWSo18Bf3CEl2WJmOx/sgNlDQV90uYT9uQtSXTdJqBi1YAM+GxEK56Lv
foc+pm8HpaRM/aaEZASGqh5nrazsSrPwA9st0UMQnK7AuoFM48WT/oQOtEKfd5W2rPfn6lvBiJks
8MjCs7CoTcEOZmCDToDCdOiQ3NYeioJF/LnxJSwbezQbWUp9C6heLl+igwBy5C5a/qILVNUHVduV
tAQXOJhsSmlXzk5N38/CLeKnNvIwHgqdh7QVc0mOG1yXt9hU2LqbFPOoIQoYseJgSjZfR6OB4ue/
9cP4/FGjB5tC0eVrSY0KU2RTtiEC9iyIUXFNcWQ+wKOzvtB+ioleMOTwnXV4+ZPoIEt6tYRBI5Q0
xIXvAPiP/kI4z/pjCNtqPInmslrAYf2uMIpQXGD+gzhkjfzuigNhiIWuMXFS3lmESf1V527r/W8F
TwNGsWPMhT1FbC5jmShJJQHZAqAzfE+EIwtGJxnA9HfdPfrpGQoaWB8l1yRznwWxGd3iXlqCL5+Z
G8UAIfto4+m1Rtclg9u2GxNisGeVSXZpT//Xj7ExEwDvWkhOXu6kh2/kh5A5QUGnqAf2jfrq+D32
VVHO6fSlrIJ+ksMVd/DwU5q0/y8ycqS5C8IHIiHPChp94+WCTDvZmlgsadhcOoYMXTIF4eqnpDAu
BKbiDxdYcWJhWcqXtP3W+8mW/e4/jVzhN6ov8LTKltWVptZ+blQNLcafDfdA7Ens20sgTZtEUQmH
r5znZhNrQrOH86KsmkC80d9zsmyuO+LnowfpQgQr6YNW9Nz50e/2giKcr68z0JUCCrBfc3l/xXx4
pEfw5N8GH2VBYpnev0bM85tKrl5mGJSTibn9MG0UVZkT5bAbIET3aq7LsLMROApoJnlcjv7I7M/0
LzczYi/HxZmQvgskn/Vo+RIXK3g117FxIPugCcIrGNvnsutCCSozikdvNYHoQiQqLOsrR6yYENXR
jt+Y+MXfUfjpI0avoMpbvsk8ESzUfxPH6WOKFgHsEhyF4cBIdHjKzCiwW4s1WqqqiWiTyXbjUeSO
CCvHA7/SU/Ti0KDQM1bmF5V2fXQT0ZevwSrRkPdI4xL+0drFQjS5KWgXD6uuKBZ5JpaLi2kFFjaa
HLY0HRd+IQwlIBthztlzMqi2y3s1dvI+nVGKH3hH6SXbHF3F55+6E6SsdpXGeyODiJJciU3OIx6w
sPh6jgjwb1Pn+8WjgRCbKhVsoCnXoLdPvPGbZBPpQN8oUo/HdKVGUcQOAfRQDXXBz/KdrGqTBF+v
caUjXOaDssOtjOUD+ppjOt2VS0hypLNESdIXF2VtyqikIoyGgj/h6UBBO7AKWyNykS+3Sx7yz+s6
+pjXFPCK4upmqAtsHeHO3aEXU3FqK7xP1bsvSZCB9sC4FZq5ZCiZL2O61dU37pQNNR1Zu6zsCWn1
QR6zOxOMViW0+ECV3L/xB2k/geFmgcXjj2VBudmpN7SlbdEWFvDEleYtil3F3UoLtPH3FFTTkvC+
es6Xp3MTxmpsFitsAZAA318mCLCEH3EOqxjlmtMLYT0BqOCRdHV2yhzSSRmSGiRfBpvW/R7ekOYf
/m8DAQ0ttCyvbZzJRVLLXwXailDuC2JBlncxT/jCiFIHqzCmjC/okc37K+h/274yAxN7PuJAWgbN
yIZJjZpYPvm7qM2f8HdWer5fc61+nJERhdWIuym8LgZ5pA7JJ8VZuCYwqyM8M45PEBDxfO+a39Eo
uT1VaPeTS8QRraSeOBBZs7nlZQZq2932LmAVfHLL2ppL3d0/pCzNGh5GcwpOn1yj846HQW2v+zeQ
0N3ZnWxu07FSAZmy9v01hGL+UbnyLJUJ6WK8Sus2NhaDitqNeDOuGxOqYebG3+t6MB2W4Th9b0sB
U2dWwAEPURBaSLgsEdb3YlRf4YOwFPAe+9Fo3/XAZuOiyUI9M8ln1U0JPGexumOVuy4ArFlDwOsT
ZGmCKdNmc+8D0ffj9kc2MNdo3QMe0zeOGaLP/cTw+jI/6CjkJMk0ovHibRZARLH3xoI0sUvxDzzo
iTWE60z0xSynDECA1pxZCRa4ztAGZm6+0Q2dkcLE1++eh5NXBi/wayUJydxLb79zYbXkGoCVeHFc
+qNNUncsd+S2eMSg1AIP/9L0PkeOdYX4f/dwgt/P6QEZZKcIjs3H741Vysb8Hc3tjka+Cg77qIXA
2tqH+EfqC0072/xcf+nk+r4Vzg7ssPa6yZN+yga6ZNhUoBOGi6DsNnsHnZZ1GTbJKv/bYhywzJiR
u78/spCm/VDmpeYkyL2GZ47Z1x6k1F8eXt567mNv7ZzqpqYJfI+iWlpf4KDDBmAe3RqBbuO6Q2iQ
KiEsloxI5U6bGSi76mpaio/N3Ld8ZTMb7Shucw2+JXm5CSFgNVJ6wuuPpTmsvjRkyMsEhyGMvw83
Bq0rs3JCAdL2OaPE4z98YSWjaWEpPlBwQC9mQ0ZoKy6nYcsxsy9BhAZ4zrG8FkRfwiYKmb68fqCx
xoN9TQjHybkyzmx+ZjngVXQtZLxA2b0OXdr0tiFVMXE1/VLMtLGu0wpkDfRibMKlK3c8Jv2ZCseC
LIO+RthhrWzrPWv7OHJ0kzB/YEP0dsv7E3Rr6oAa5OrH6vYzjnj4Ci3T4sCbBnZLMjkHCHhmwVq8
vxPDl9rfHKEoFow/wOuH122sg6kXGskmoFGvFWVOcNGMZay6YxhpJ3Vuxldki+rAgi3HLTSXht2O
RLthKow5srzqP6RK9d1HIwaSerDES8sSNhcmhBI0dfNzMwKDQJszsXRQiLZ0ZnRS1NcjMzvwEAPV
FTW5mskJg4AJ3HvtgCvyH6wokTKPQxAypbE5pIF1g7RclOgyUgZXkhwDnDFQ9SF2xMb0utrVwDZk
oJFVWNSstn1EDr/2oblJpBcLPWFBHJhEZy5kCpINt0yHOck2bXZ1EeHv3Zo7OMwOWfj/9AnsVg4t
P1W4GkTjO53IplDazw3GTVzc09PsnXTUwm9g4k8lQZP0lVrDdtUyv1VQj96+ANOdylJVeRr5GDdE
zinZOlSk8EeoeMWmwlNLOsoO0qr0qPeXIoB2dLcyCSF24r3N2u1rYqq65xbqMGADjFc0AfC7oFrs
zIS0ecefe939qE9ZE3cEZEuwn447o9wjptnC7woboE80DBY0PqrqCRkV9bZPGBpYj7ohlS9AuvkN
iQYjLivkT9CmQogfdNefSVDrxvIOTpLAQJFe5EFj0FhdhnKKEfjoWvmdwSLfm2XxS8a8IhrK3MP+
CbeDStkuQvSk7R5rODaSUwTnpyWyf7UAw1djkJjSzBEnmXQUxWX/X6ob1pDByhMCEvBi+2Ro7Ezw
DCx4rM/RtcaGcdiDWINYdW9Bn58QZmxtcGYVYr6P59qcn5N2U8zpzm8jVpu1eH0HEjanSnmL7Gzk
VUagGyjji7oNLXlyS1AY/4CNWDCHvvXSQ4qzEZYdyOd7FbzW8eOc0AO4vvPTz26UYqDknqCqQYOW
58dIL/9awBuesszS6K6H29GWnh5OhStHOi/8VLzB5P/x5C+a49BujBBEirf8cTZAWczBxDbUrtef
0dAWIwevoGIruoqr5aK1ctJ5S4Mc7Z9Vj+dFa20Fjq4Bt8iFcU1Kr7BZ1EeETOk3ZUNQTGM7IYk+
oNS+QrydMLNvMLPv6HZXBODaSnSxmrtA9vItzUYIyZZ4JEEproFM6ONAqr02mPcbJBWddz63TTyR
Hb7K2gZAryqr55TmuQMkqpYIUlZpATxe9BJn48/8epK4PUHHShIrqiLI8clN9HgRHHPqafjkn3xC
pQr0VCo4d3LAz0kMgmHJlSmWg7Fr80oJcQOXeVKZBjSSZdXAVFr3dWoSvGL3GEDwndYj3v8QGhp7
swFZoIgs25a9n0YVr0odyRXVr8LK7DDsriRNgOx0g/HZ9+HAY3pjL9hCQVqHABEV5odXrK592y6R
q6UvOqOGNRX/uv/dZab1kkr/Hi/fQ1kgyDVMaOnlgnQFXUVrsC/p2udM50TkmJWOq0oGxKPxBLAF
iYg8ETaXNppBwQQBIF0M0rV2D+Nk+oCwa69/gpE0Lm6nAHkADfy+eeNYaeSatuxGEhTLL8J3fFCJ
hjddSMA/27OMXVYcMXtLCpNvvt0275HLV9iImaq+/EW7OmaB2F03566yHoIYCm1bI9OBieFdOHI1
q+dSabbnWaMYPfUzGOsP0kPn7xzPATBGMfj2ox/HLnLdsAPumVSzlCDHLMhHwLWx/9i9mdrn36ZY
D0GMCCvRdhfH2ChXTiqQjfjNalcZFDVpwsCZLtG3jucwvrnb0RJlG4pWTrfDPapZz/eJQkNnOEjY
w4k4hZGHUlmTqFdb6Rj4WbiGT6lKWA263rC7Smbf5kxe+4OC275oAGmDQc0hWaalTWBIq9Vm+vtn
ZQeAc6gDKkq2J+Beab/QyI5wWRrWx4cowPkk0lCRgJ/as1fhxCiyDnT5GkJljUIQVjTx1EQxL6Rc
+o2uTILGu+ff1Jkoc2J0mm9Is/iLAksF2z7BTBvsBBRKTs4RZ+3V03xOpMC5vFDT5YgXwcrBUkSi
GGIRdtkubupJ40YyL1wgR8YceQsCtO/CnHqGWK+7AwKiczuErwWTeX20J5HKOasN6EFIOkW2+n/q
PntE95zmzUFewil4UDneGk4WZoZhBvzKnohKg39w1dI8ck1WgX7CyORHu0b56h7VTDfQy50Q+Fxw
1klxkau3RRbwA1Tgq9pRU1K1AUTuW+CP/gBPoYaRiNS+yKp0UFGZBVXb7z330p+x97ysi5aot0jB
jIA361J/rbFSo5GZd+7bFz3biJYDjTDQxcQlAEkAjuWI4v5Za0QU8xhNjxjRJ+pvrW9D5inUAs5v
1UbwwApnrPOlMR0/pkv94i5AOWyNevX+iB6GW6FKBkCNqW/y9K1gaLLCP1YLDnJxCiEaDeidVVJK
BH1zo2vnED89eo01fLbxrcbfMLvffCqHV9phXlirWVy/8+6JV/P//u2i5ckq8sKw/XtSwOUoz6h4
/le78As5MFNYHSTgBoeOzxlPDNuUD4cdmhhAAEdMgBovePJBcpOdNHDktmYldyqC2nBZC9m1MSOQ
QApKfcoTRB30ehn1qU6BxAyEmH+Hu69Lx0CncDJw2rBIBgyFeEcf8Z8G5blys4DmhKWkxVK+VSHE
Sr1E+FeGIGI0A8/Kh4jjxtoLnszHb9CA6c0aq68DZLx63C/aI3ETc/OVaCHi+Vvhn5CTyNnecLSy
0YKOqYkm1ebX+zH3ScQENYcrYfYaJFjhgyK5U4yAGnUbGO64YqcB65eMzwdA16LYbod7I4hFRUUJ
/54zQ28TkXoQwvL44LeqayI1vZKtXgg5J0L9ZNlkPAMJyVmBvGbP0yGgloHiNIw9MkQpHYP3TT8l
xI5G6LZPmc88kvWWSr7CoOz/P2MavNhiRe4mPF/x4YJnQwILA0U9FFttD9Z9gnDUgpzrE2kljBR0
ewloKACc1clR2yU/KD1THjaYepUNDNjHBvfXxnQLYGytroDeB1VHlcuHa+dNrk7QDO+TwRgJhBto
8i0kjN6MDTsegnk+bE/90+Q2Iy1hhzKXXGc5Eo5n9ewLD5KMew2TS6kGkthy/EIKKvsasgnCodr+
36NtLydHBmhUjHxhuNJLTWF518MIuaoTt80gs0WNzD9yOJBGTeBRzceLPZ1jxlOUBkwogWAu8UK4
QsENZ2Y2VHvcALi1LQpOICIcEW3jjbKkTnOP7naGIN3EP2eWsn3PMg8SIBb9fHHLnZ/8MdctmZ5m
WuzKhLSe7m6aBnkUGU53Dc4M1UYfRR0rZ5VUe//NyYcQ2MxOP1xUR2GNTK6cC9voqYsUXWi0a+eT
gIC/oXHNX/r9pfVhHNVIEarTQ0qwPpiOAkeEs6Z/RX2yHiSELkyy3XLamTEkugdJtBv0EYDCvkQM
0GfgRjHAfFEgPI6xCkGJ3z5F/GrvzkUA9oxTIE7AQY5tTuaxLh//pYcLZyzlkQzPaC7Ll8ZY0okv
QVNo8WxXFt6d4Ntv7XhPnpv7WCQ83z6B/xfxIr9NHbxR8SGxE37TUSdAUnqeQ6WdGHKUB0RlI2OJ
gXKVJvloJ4tmk3X6gz2r6+v91BVtLRp5qxPUWK12Y3B8QOYcxioJAGsiPrfPjWiNf/tHgDu4lNH9
BImxxJi0ePNiui+o0a6MATYsHcvEONkYgim9A1TT5z+h7affEIYuyMBO3AqKGkp45IYOtwdw+pNf
1B9viwwGg4A1LOI/1YaqHGVh5jRgiwSmGl6KM22wLJjPRQwqoigY2w5UGKCJbYFZG/uiORLjwzdY
+ghZttJv/kqZBfAZu3nD8A2VpUD6F370moF82D6A47uByKf2WR89CM9VB6LvFA7VZ8ETJeQvGge6
4GjloYDd8WcK2nxQVekfFeJ+pixt7k6osksOL9b1cy3pqh8BbjfuzPV+JvLue2TV10N4hifpX8Id
XEYdGFTNIDySSjfko83HkcNC6WHNZkWdp8aKJzuEupdMxagUX/W1M7Hcp++gAW2SwBYNo/mOAvuu
aZem0SygmWe5zSgmeiQ8i8/j7ygOf4A49AQAgJ+nDZzSY///wotqikZqLX7FIOVHMeOKmotGgpzk
N6r9rcF7zToqe0YCCVnN9qgJlxRNS76pjbUXkLq/aTNTI35JXbbz+3eXWh014qOytcPh6sUCC6rb
jO26yDSjm/kSTzp0TB2rCi6JQgbp6HAWUwzFENjzFFvfHHmXRAmJRSyOxu2F5lgEwLwbw8yaRtOn
aRbT8dsIHwmboWd1kW5KsGFHUWzI3RdqdcCV2AJXLUDGZ+ijjQly/9PV228MJ8tGiCpE4kWjtHyI
9HlAhwzu2hGiqEFunZD3Vu+fEW7C4Uff7F2oqDWUF938f5AUfeemfMWW7rsTiTEYS2GsQTdc0zRf
t/cgMs8KatY/trcFsQw3wI1Dxl0Q3QrPDf4Z/3Ao1IqZrLCYlESsOpmp0/BIoNaohs/s6tb9affU
Jga1deR1TYCU+7cN8CuQzdt+wW6XuZbHPL2vHFw7LPRFRNqWmn3qEpVzrbJ1lgqw43pk7PY4PGx6
caaoxAtMVzvlbE8c310KjJeOZlEQqHjWWTgLoug6yxvIYpr4OTe8gZGka15mtBSy0vWDANIfivzL
U9bWYIStQkzsLFzR7Q30aHpPMJHr1WlVgVBjPFGbKmRjw8Zbfs8YMkqkD2AWROr1W91HFYPhMfUK
zhBsJB4xB5ZFXjkQ1/7jst7EM3+AEtVF2Dw/h0X5sFXyI5SMPPrlYj3hZ3OX81fA5Azg3ngSNaJ5
5Y1XTzy/1vnyiFLFmwjgWLyGLahyk+wMX6RPQEOEZHaQkVveZ1uhkUYM/nYe1SaSYZPAu0DdxhkO
KWVS+YqnSNR1I7nejNUoaHsIxOvN1TmU1HXMHk6aADs4nmIomSTj3uk61PYNgLMfyDT0acDR0Fsn
K0nC7jGtTm+O0Mhf+niEWXJNPoZSGWP7DKU18bymzInSS3Ag7r+pkdKCzkacW0ZiaAIxFUd9YbDz
BelrmZYMW5mNgaidAzOzs9VWrpZYTTg6V1fO/i67nRbzqyhqMPcU4Lhi1tNJT8eJJ79hIxfG0Inp
jMyK/ewhSZgIAYIu65Cn+bGkSFenW+7juaLqdm02Pnz/JWMfpY+U7HmRd/hIKqt37eIrgmLlch/l
844Bi+4HQOS++Ak8tAbKCgEINmnYFnDrSDh4m0B1FiFwJxz7ndU7ZMQ8mIX3AvTSmDAzChgCcQHm
5XPPbFSEU1/sAfdz5esdfCkE3rKXpu2NRZhNDlMQ+0pQ+TNW4Ib8VysDOZhvEkG8oK5WPA5NKEbU
xSJlfPUrwi3lA4TdHfPsj99XgmQH7B4u1IqUcdYFW0RHbAuqnoSHvEzcDWNconmaAWpHOpjzNjF1
STpw0YU2tPz96EKoEubVB3bGP4rlWI8aFfHP59F1YWJ3cwQ8vxLkVuwE4Kxn/kuprbblyxxqb54K
COlbUv5Vy6vAedMJyvesVcpI2ETpVhHPPRKJKc1+THqodJvDjImmLZOlCAHLjR41aBUc0jaodFKg
TvvQxUuo2RotJ4kb/Umu/Gy4Q5tMll+3StNzfpH3Yd771PIe6R2A5sM4nWan2kNBzqYKSHJhv+fj
NWnXQ7PKFs6hHOB0av5xnxLqtfX5JvocG6M4qYD2pJlydn4cMo4onNCFg85lmHQOdgFWC5SzUqsq
Q0JV6HP8LRhBInGbTb1iHDFHw8HuolFtlos7/d6IEDwMw7sFDg/Ay0V5JCRSqtolJCGfHcobkGRw
nhDpM3+T01m/4ZT5G+hD1MSa0OF+ncNDNHWqMPmE8YT8cwqhOBCChK+r0OmDrMRsuHdwu/ucY0JV
JFys0sqkifTyF9fb/szHMf3uCLPQfpb0Fs8fGjPWwlbqoM8WC9oqxC7OcfOB/JRrMncmL7bqZW0d
ekXkVUuWEEwo7oiJ/ojWP4e3IoZjyJoXmo/+fb/AASJ+znO/vMZxwIBzOLTk0xhMy7/M3yAMbLMZ
mB/Ibec9ZCatZ76QKM/mhKzCW//BfIRho0IyCJiXNi0d3QsLbkCGPUL+yOvk29dI6+BnP8kLPMbE
8Dp/YId+61cB5ecujkffxH2+4O/XuouWv6pPED7NAJJ7gBgWMFUbMPpkUA22DuaQE0GKS0ZTa00i
hQFUd0VP1NIKeHX3AO7FDsnwF+1wakd0SbHSIiCyIMyA56k8yIJ4dTu2/S/JO/NdTwbSaFi1Ug1d
cvieUGKIlFJQomI63Al2XRPViqHoSx63eW6VicnI1883HFLVIyq77iHKq+boulHgqf3gFjA8BmJu
4xCAXy20+6OFuB6BBpJhjK2wKJnxg1sHjjNdpOOpGCoKCAhUpRlwiiHf+zdIFF701CoNkLz7W0iP
jq/oNFpl3ZSuii1pJcLf48hurrjlUGHhZh42jzRiKfsNpduP8Gjig/8XnXvIRGd6nZGFyBl8+3Ow
gDDzzyYc6l/Q1VBAhqy/4sy/TsJwzJMpYx6MZ9ZFkddV1jlVUs/im5CgUFK4IzEiuXt/SCsvhyQA
3h2LR8g+AGjr8KV0/W0G2nuDbUpPIoPLpZmcrL6ZoxI09srREb9PHGg1i/3nK0a2DcXhu5tSgO2m
aNThL1y6d2aYHggBH06H3BG7O0Jsy/Sub7/1PeMgEhyD4NxfWfXQnwS3hw5Um0wDwZOovKFQB5cQ
OeK0c3Us38XCwvgox0mnbyNclREuTFaSHhW1JCKNc8MHxuQv/7HmGWX9Dahp8DIEfuzwzmEXJGgW
uR/TLDWzCIokYZ29Hi9h1fEDmFwaaqjOZh75PuM15kJUmJIDDlee+QTEsZJsnL8qNJ6txLlQhygB
tZIhw6Np0jhCmKxCSNAN8lrrolXn2HPGD8LtFa0QANs5A+0clSuRc3A0gcBTz9ltQndJVsTgZhd7
gmcl3CeVFJMM3/rA4jbXv8Shao0Fu+kC5UUaIgGT3lFJDlPj9tOT55y5IKrdXpKwL/xc3H7RfJbB
LkGfEgLOZ7OHdeG2Q2sX7YwPxZQh/argdOmkA1ivntsaNXfBzd1rUrazHHOb15zOIKDhE7kfUJEN
ABgRXfNtRVmvuL5m+tHEzkw5wcRvL3GMeFJaYD0Zk8mVDYo12VGIXL3jPV2wRFXL7/Cj4TrxPArK
XLjSNBpS0fHl4wD/KbyZ8wTAIsYOZWo7LHrjVxZQKsKiHLEJ0XsTc+dMNOs6+6FmrUostd3D/EFr
DyXW9/5B3Q6kVTlfIetvjecPRJUpiARVWcboZbEeNhWtF79qyfeROFpc5cU0NeRhkIc5WD46Pe0+
NDqkfRTKv1q401H2FY7OyaWl8VvJ7izEs0oHgPs3Qd5tB+OLG3ML2//n/DEQfAomCBkZPosBYthX
W6cH12Extwkx2khEfuIXLtz2fT9INsQZLsqmCvUH1uJ7RwQlnrjMVgyNYn+OIv737mBjIdp2T/47
l9hV01WJsv4bXEGbAKwcbuYDAOxQdv7SbHz/MN9Zcq/v9YrnEy2MmEJOfo32yJb8GlW+63TqRj7r
pSj1bNshsr9eccbPCcn353Vk36WgG27siwHcITSePhT5OaDnkHYqjn4ddkp6wgZ4njbMQpofgz+3
rSwOZqIziVRcdmwlJweIiN+cIF3DpjbK/wt4vMFTVwWT9n1V8006fWMOoTYGzfMVtWjOjExdP1Qn
p/YdIre3T1VFEX7/zocrAXcZMEiwIYiOJl2lXScGcgkj6endSNJ8Vef6cntPclMFmb2waUbS5c8T
f3Zqzxudb7rvYgdB8H808tPPwvGAGd9U19nFwBzIGt4/krWeJYKkSBwaxz3wRQk8zroRKw/iwU//
EhkfcgewgAUn+kc+QObjNyQJdAoEhzvTctciZ9bwdzWwct4F14i+Ee5vxkbZAWjC5dvq/O/QUsNp
S/C4VeHBzrrmAAiBOq7Rv++GM0xdH19u4Nv5EP2yKtZQ3s5vpQEPMG+k1GIvx+Kvb0ZAPZDHMGKU
ZNBO2rR6Ki/juWEQ9KHll01V39eLzi2PgS0YhsE6wyfm0RTPouMuiCiyz39jtlRoTyphN9hc2lRW
dgrE1Rni78rhE4bLdl/j+7JY9LgKPu60URqFAkLWzbNjQM9jDHgiju6zxAaVrvk4sUVfIWJgFtFn
dw3GaUjt+rkLzoJrDWGCAB1nDyTAa9zf79Dq5WXWBMAFrFK3zndErgQxmRu8LDOpmAzIQhy2J57Y
dlvlQDR8esE3kuTcxu1we7/BlPBaO7ZbjchU8zZdcTcUFUnQmgcZInDJDWq5C2YBSfVsHlHtNkwK
Wh4AVyDTjhmmgRU6rz/JCZBQU8OYkiGTmlqv1F3ARHzAGT0Xb1CAFFUkE4jjlC4QVPbucr3DuIqj
SxAGn5vK0bB0bEBEhgagDWM+Gzo3DiQ8PniGIb+MquLubp9QeJ/0Hq9HzCBsYXKvaUTP9g1dRiRT
Hl50OAlPdUGBAH2xtMlxsqVP42+2RKvKUlsretN9oZ/U/6Vt/6SMY5ilFLdzVcoRr1iuABIVf4SG
h2LqMSY9g3Ft/KfLhIC2E1FC4bB2VSCnLi6vRVPsU1fC4D3gTubRODgCSeC0EJS9ZrXsJAobB1RL
U4cRJa5uF/agYwUiQoz0GOz4R0cqrI8jqgHQvbHs9h9GLfv/hSVkAPJoqdM0tM1YVklOJJAz6CeM
lxC0MUioMs/NExl3mKAAEYdGwvX8JXctNSjwSYYtXCDEc0h1yb9ZSaqV8TCa5JDHKgtnZeOG6R8V
tN9hz8ln7NngrJRdoyCqXONpuBJtXpodqN77GkZusjhaYCNkC/QgFYmsiKu9Cl9Bgu2NTtuwJ74G
GZCZCnTswWzH3RU2sV/nBptxWNCeHWhIWU8OqeM7xaMHBvLa03cqes0tfob0fOmuLOheL6Nrgyd3
ruZyGhVwY8zTOS/7dJxKXsSRMMEkjS9A51dGZLVpAixqx9Z2nEQzlD475xBPvMpc2994RzXFZOxm
edIUnmvvdao7AqJj8nshRyqF9Y/DB5P4UOk5sqU1U6Z2dCfcGTpFEKUxfQ0AGkiZLPkl/BePBWH6
yz97OtEioPofLGnMznONrsH1Sppwu7hvmGUuZSc8pfwjJurcVWryQob4PoVGKkkUlMik8IY4j8h1
zHr21QiOJMxFQg8m+96t/JC0z5lkKM+zQkFFzSd59HF87L35k+dYj/gVKZJWQZTNy06eDHZX14gE
JfaXnoabkML8XcDVlnO8R7skT1p27NV13mST3ZDcLs3cUKTpHGUPKcZk0qqb3V13ORU8zXaZpdT9
elV10AubHsaKwVz8RCkZlq7X48PukMpug/CubkEwIzum85o9pQsPmrZv1XajyUU7tY8N3/IXbOYs
whf/GxGSBvaf4LFQdO9byuFL9Yrssx3jl2vzXfJdTiS5q4xPOucfRdkrU7BSBAl/N1/ZO7g8K9ro
yLS+dxrX6DN1NtuU2J3lypGtMVBvOP6wYtb5oVbmUQu7L/h+hSPBB3tLWSMJ/l/fVwycTNphKdnp
FDfDyKaLLWJae1l2PuZwXa1tQTpMdgOZ5mAIdHSnDWkAP/hoed8PMyXUO/3oR7UvJUSKTsRNPZML
VL13ahswN7WhokFewbrMDCPWxJ4LRBRDUM4mhsmzcuOjIDmLf4w04PBC4GpjGowAP98AlhA2ubMj
HmHLHkKtEhTgcuWbSiW7WZnNiBI3XWP0O4zyoQX0URTVCdDhyja/LWCLBqJSjctklMOYV2pGQMgh
2m18csNDAGtklxSxyFPPz1bIg76QZsJDHjsb8yYKaClywElFX4j7XD42+eTUHgV/WCpnG0+U6N7q
seiIdxGAb+w/M6vj0MLzvRbZAfzhPe0QY1XYo5HeV5gHGQ3b05sdEGYB5O+OF+JgdgykbxN/B6iR
2PEHutzZvpUVBVJc7SGqT9qHbRMyhQxsFOcMRTszSTEKbV+z8kgyiAzzim3BnCq3FcPzmzApsxuG
cttU/4z9dkCa6VTILNkkPDfP2bbcLnqmJqdeEryeYu7Wp9U3I6krikgAOJtHBMj5dg3nbMHMuvwQ
APr6nMkgs17A9Q0EQiSS/hw1FDrGWQp7b5NxZ740l8zKDGOVtTOwOTG/n2l9/J202hQVa41b761p
flJ9jg7Q8DDnORc+wjITzT3lI3j7WgKPtR3iozTGTekqbX6El2NnoS69lXdLENjuSd5G3jDFDYCp
pnig8eyLLVEGodLd0QRrGoE5AN6m0pM4zrvCW7LiE0z0gYGjhSRXy4DhybL/KO7T12OVep4f4y64
c+G1U1Jguu0lBAYAzw5sFbsxeJOPvmiTsEXA2p7WLnlaKakEVQUMRRaAZPmVRhFMKybvP6HBG/gJ
mY3YCPBS1GJgcnH/E7n4dWgqZEfD28FNmpwOV9hsTIykvwd4KaP3pQW8bR5eqW9HBI2gvrZoSwMN
MXJRcxBHvr3MPAu88gm2QS7RfJZDzYA2ssRcE+SBiMoFSuf9qoe+0AdEXDhk8U3TNDW9y03GdV08
70BtsyHMy5f5qgVOunGkIi2c6UMsH4QhCCoiT4s5sNO7ogWuWw127Gm0AQOzMsZhLbAQpRMQwY+U
7PF9mJpjfS6H2OJn4U4KBNnzuY+pL4XnE4UqG9alYMRdcxBVr+w54tsnYdD3UlGwMEyyf69GNc8V
tbJZQ9jMdz3m+H7kldeHrtbi77lRQ6tlkPC0hrNPElxhxouCkuXwDtQep9pon4SDCCVY1WxLKLnp
mBa9e45R4oyiVJtWexBrmF5/ZsGmt3NWrlyNxNjRCBeicdrJTZmPQu/gPjl+FEbK3NQ6SxRBzkEn
748B3g1ZqR1e/fVy8MW5KNk6jpiPkB68wSs1qXRaqVzs9HctKumOeHoDe0tr+utIGYIJumY4UQ9h
9OtWtBNoRvJ00qco2MOvmf/NtKVjpJHqUssetBqmrp4T0gZXbL4oCwtq11sJG7DGoYZea+sKMosA
4PBdDoEuWdp6NePxc2Sd5whP+eWWZYYlTSPb0bTr3ZZH7MswdIoK8ufnftGyg8EakZ2VNpKWnBVR
gUzomRqY0SqOuGr3ojzEpKD9QjseAwdOCQOFHpgIZji0+ezXTueRLJxjvTRHkMqPfam33E5sUMCz
u1hTAAqyfZMQjMlUddWeXOl8NJ9x4Ac8eZUjJHYEO6mmJDofOAeQmF8d6NKjSJMg/BHBTTjhFFi6
BTBq4C/qgaLXVA+8Y1/3YpYu0s8TV4a1XxCx9s01TS1kAY5N1v8N/0eIAvrJnQ/nkoSHvYV4jsot
DRfQZLesWEyj8GrNMhYjEcsVRarNH9D8QSD1gR4ZoCFrjZmFo1xKicTu4Xb8liRsAcdgq+ks55xn
/Iw3OEMMbcxrD+8nBh6DXFnSbmE/5X/fSymHUd5CNbsfNe5eIAbIN0i7pxkuP65Eqlh8RA3f45pu
B9864PJW/H0K10S1dOnrfmRZoBzjj33+iIvAfUQXUm5ekbGygFKja1j8BJL3G4dUZJZzN9RGe0nN
oWiDxRBYXZfh41N1HXT6lcuGKdlgn4XVEtEVnMvnWSGsti1eM2idfxeO4bI1OB+MefjGNEVPiykS
oD19klr+QFAF+fcEhoWSl6TnqWwnf04Qh+SOn0v6Wyrl/Ae8vD8YWccYvlgx3MmK5xyzN+RNV6wc
DhoucoHFJ9qkStzVuYjON5rm5Za34qXhYqwWPo/LImSe0CZbQQVn2ZEqI9Y9SOvFkRj9JmJOB55c
MOJhXrGYBEakVrrrmKqiI6HKmqjiCGmQ6p8Fv3Ohf1UpAFjeehzFqHJK+ZNtd1fcz3luvFKRJx5F
YTcoAbvFPbwIPDIwq5gQYaVmXyZpoBDFzqIFGu96LLAYE7FfYyk3tngujAmKZa7jFp3DtXkFpJ/7
Hv9Y7oZNwu0c1+GY0rXyr4UNFEdgQZVjhaQ9GaKgnISkCMZwYYmVcrLQfgb0UPOEintOhA4Xx2x9
rNpB7fXjpm9gKx6Et4nMNE9cdNK1/w1azmn2hxKlSDFe/r7fRUdHWEDhaR+si+49CTzgSEFarnER
lUHZO+vNy2p8lm8ZDkX3p0MAoVKHhdksB0YqKDwj7cLN3g/kRaLtPq2m356KFcw7gSOeO59PXA1B
kfNZ1Ikq90XoZ2yfoXppdTCDVt9w42JYux/4joRoSxkzOehXVrv5yMbEJKLb5lIjIZhXEgki5nx0
tog4iIPPTV+sKDpAeZdQ+MamG/oWAmH/bEKO2qho+MUJAnCnMcmMqO350YTUTsqJII9JebCmaXTh
GlGr+6L0X30rYUfsfomm+PMeghZv8Hag1pwTM9fU+AZE8puTX0XbVKrfVeHrxxUgfhC/6VebaaBe
XqN7CgubzQMQdx2SWAg8iPFphNZkGLOMQjWpd4ajdCzMeIxrv+GaGYmn6cuXnJ43hTKirjimYO+F
FU6myJaVICWFUouXZCGctgtSBHurvjG1zwjn74oTDfy1lRau2ibg9IN9g6mvP27yY72hzObS7Jur
bUAyw2cXwf8HXFdB8WzPGCDDWyPTXF/xROdI+IcvQTGja8uwyHyN5IEXYGCwaPGTV+Bjvw+HMytA
1YOshHHQnLBbZ2CR42iXDJFNKGNLXuvCkCBE9TCHuZ8OAe3YseVt8+5OBpzahVL8l/+MjRLGJ+WW
5wwPkrMi9kKltDWnCg0ZRA7ORd45kyzN6Iv+qJCRdR1wZogSWVJuijD3O8eK8vutcC2CI0Tm++VT
7/1nNdwnNkpUVA2oKHckhMwRuzWe2c0eFF2J6+E72ADEDyGkgqwWGqo5Cg5LjCHxoakGfxnQ4adO
5wiLDTi3Zbl7B2hSDExS6t0/VfdzhB0OejdKXQ/2RAOfGSyk1gKsBRD0r1Q69qWetYumKi0x3cVg
rngdSUuOFpKx3YxHytllA471Cl1yKA2b6+clKGM2qHt8S1x1gbhL9wM/gaien8uIvi0rcUjbKtWu
BdnF/sndlvbsiK3WXU+Qb1naT4MpKOwE32oYCnh/U6Ukr4jglNRNF23VPV3JHYkGzHzq2hmmxCEE
IQfOKIsUoKZwbkczt/38FDErYcN2CgB77NcPS9GwWtGdlgsYn2YOwLweStCHRsHS/I/vBqnS9FOt
f2g+zZL6F0ozp25VU8RlHLuO8C/j8UEVgPkbu0cg0q9mRCttxEpusvbzSQvNLleeiEp7bepJxUsy
iQsDb7hBvUHvt+vlRaOr2o/ND2e5n9SWo2tSDaLbcRX3wLE6Mucl88N09end5qj/QcU9rSJqkzfV
NQkQEZnP0YQQpYTC8QJPHXaEfK19PuqgTEZmLLKHOBLTZfUfXTUa73HammgWsV0761zKcEByoXAB
Jc0+qz5j0/prtnspE+bCI4QVRrl3Jn+zdvCeK358N4OQyOPOPu8b/pcDHuPX3JrniE6jVhuWr2ac
V7ZrEQJOOjdRchY3hptY8ULqQQb7REupMfTKRkFaE7iX1slZTtWWukSPXUvRLQWoN0c0DtC+2gAF
0AHUPmRs6EoX0gRyNbdo+91BuklW0mdlKv9YkyPkuBQiUPtK5i81Y0XhTWz9blax9KVziybCs9bO
zqWwKGO1HBUYI8Zw0IHluiKdkEBwTYw4Iv07TWEwxbM1gWcaEWwmeGnLHRLArrRW8lsEruo9bEuG
qGYicy5wTgZQOSXZVe7os8xmO+djt+YWIRRmFZ6+26hGqikPEEX3uTUTGjSvP25mn+3chotTgLkR
hQIrUZK+9qxHhV/l/0j/+t0UnMDRPsSBN3upo5hex3xppVAO9m6kSSCgZ2fOozt+9YELI8a0kP28
/k4Fw5ZUMx65vH664v+NF/zGO/QVYuL1M5tl5/OxTR79UiLQ+T1uaBZL0ohkR++8OOL3zmPNQhum
pYDCpMVLmhI7jCcO7YjJpdEI6r6A0JLYbvO+GJ9PQ5OOMham2wcP2QMtRVPqnXCXbYj6iI5G85Sd
X6gMR5qkiYpGztCNsmVLEH/kyCjeWQwcm8/srK3NVpHUEb0C/3CQCLi90BM49VPGGxgs18dCtFzx
6MAyIdrERBqG+9fd1P934seM6yHwgXxW4F/Mr4kaQE0nK14jHd+mKaMrzUxCq9MN25etZBZOLH7c
xwv6WaablHby5cruZ52UchSv7Sf1qYHCaFyF7e7vfTY3sF20vemAaMvhlgbfK3FkjGy2uHyit1Jh
ScEyooNSyhs7M+4enWv3onrMW1NjgkcBPyiSofc7+0kn4Znp+GgKZaQyMCN2sDy8O8M46z5yzct6
9drxOZV0jGXJ1VEVWEn1XuSSDgigq/qTKMonnYNyKR4TkTXv/qtpkgOPd+31l8KziBBTmEdLnn+H
X+49elPQs+gq852svLxVoHrrNQve3XtK0w8fehJpsgA7uhGC/floKlirNNmn4GmGu1V1YG8T38z1
oiYeekwgoj2+I4AgDc5jSIhoAHih4d4a4E2hjWXrcpg+Rh9LlIiyK8yEaVxqP6XZ/waiWL+E4det
rZ4FcA7r0hw/s3u/0HsR8QhHm5IH9HH5bfaUgPz9HRQYrCGq5sRV8NfdWN/7haJXu7YoMpxWSu4j
69ctG83XshKdqyGGlDiE/weXCNFIo2AqQCVusgcUoWGOdPurs7b2sfYpqPO+jrKsln0XrV7ljIwZ
e/jlO3G2BFXlARQ/9wXzbFZ7gyAIkRk5twrOoaYxW0zTOC/SQCBnjW4gRtYr7Tb/0xgJ40VIJv14
Fh3szx3JkQvI9VtpVeG93N6lsKRDPqItpgxs40I1jAm60Edatoay95stXRmQjx3vId6Sc2k5sM9O
TRUhh5p9r2mlvAiYlsvY3IEg4W4Y7IwnTsuxHdvDg1M1WEv+J8IE5FZ/6albPkZQawphJvgeqpbS
cZ/roJbw+GJ0yjV5nnyGEYnfU6aAIZbpHQmUfoLpDRkTpW50SLMdi9+gkbj3O3CWgZls2b8UMwIj
j9cYChJI/mG0BW/sGu8AYjON8JayG169Ge8UP8uCLNbwusIjTOpwrvRR1gry2hMuEWRdXC+BIP0u
2S73gO76oy6yNDNwWRu7lhqmHFQ1YDOB2bWiK6QsoK/6aJ8E3XyaC1gpC5KPHIKHG6qkHbsWIEq3
w+vD72gbsemb1pbRuqzf3sscZdKoaZtEiq6qDqlXSq4u71mObQMdUe4KQe+RvqyB9GSTyRxjI7Op
D+xtmA0C37O6fNIIUsA81QagSqA9TW71YNdpz53evdNnGtUN7wKQwChDYgRUu3HbGJOXHbP+DSpR
MD8pPf3nDRImGMPiaJ4TMSkrgIOjRurJeiEJpzLD9V4vMJMu2g++hfluwc7Uv71dFvFZXjB/VFFW
dCGanJIkZadC9KWFKTJSRYYDEiAgsdasDPlINF6rGlAcIJtUm9O2hlKZEapMeVER6k5WiNj5gyKv
UFoW9v7ziSqvjdQPGDsGvKhLiCB1UTSRJ98LBVXcY6xXHFvo/QN2THCvO7+JLAX9XBwFWA9jkTS+
MESXED7IWqYoLInlDPp8FNJA66CqaPmWiDJWK5bA963Bq3M0m9NaZKSGWjezmKZRfcpB78bcXCdK
wxyxMu6jBVlr0+1EFENfC9i/CoLw/QOFpERWJg3svVlyMtou/u6V11jjIXMyzo4HTIM++CAyNYi2
KqmnNH0SK75JTrDZXsU9VE0oe5IGNmfsSehkDqrNvYyFojn3mKcat0b2Gs1VbGxHvR3MU9nXbYWI
zVK2MwT44uGHDkGzSyDHdkFcUe4199Q/Yc+oJLmihclFfwogMBHG2k2+Pu65KM47nCwGbEtncOLZ
qHYW4G8/1BvhdTmgswxjBRjnW7Fov2ZAU8qGbiczAONDiPsnJOD2psv/CrEF8zpGMe06hkamqvVl
UZSp3wtBfRynj1Oso1IxtbyrdJAO/m3blVMQTYP+2e1un0LfW0yDG1fQzSxGPt7yr/jqz3cxUqr+
7PGAnj9t61sFIJJr72pACG1DrQcWKnV9XjLX913UXjlD5B90s89QWlI195AQa8FAavZD/17XdSOJ
qaf1QahleDNYolwiz8vhPhkyK2wGrh/AdlOJt5R2SlY7lnyXxN75q30mXAnu8NtsIm3WxQYwlSoj
bSVtO9/+dCylQ18iPRXhbrRtVQumFFf0J9C40crD7y/bJBDNpZdYb9HHHcPvjUuToQ8pQ5m/l7cN
cEtBa4lNDbJ7rtZmwgyx2SXoUey+1ZTDmI9r+pnB3h765m2n4sJrjHtSn1/r7+P3lgwcwUHXFdn4
m5KI3ithy/JtshZ+6plUiYVZsBo5coNSJRmf6sjE9dpUmS99T+wc/42KhBd+ogK/7tQSx+iIaRBo
9CuPpf5BpaV9wBQpayBGJHFnCHYyy6t/z445+Q2mM+6zNTeGmfQDG67m7MZOE2ksKc7PgjJAivkU
+yEnlDgSx6LalOukKfw97FBTaHotinm9eblNQmjf4SK/ky8dKpsWhzYkAnLzHkiDJGY36rEjW3/j
rnQ+Lj+2h/L3+HnBzvlMs7QQXeW2skRY7P2kSzIYGiQA0EQtLs2ek1WFVOZpUD0yxPdprYW8R6J7
OwsDDj56ebntwiuv3uns34MwDDMsKwYFk6I00/CtFo0Az6qzgQBjVLgzLsFSPKAKET7fhn6Hn3IM
qqWboh6xQ6QrGD+yQ/SaBzElLcMtxXujGMqj4irLftNHrPvIzHHSEdXI6FtwULYTpA1msEJzJbft
Uzg3nVtyYB7YTaY0bCiK3Lac/bMbVQzMRUJ9DJqdv9V3t3/91GqP7rdtJThyVx61duz9f8F/bR5D
xL9l4YMyDHsbwyuuaU4UNz2FuSd+DBEIy3bR6b6Jc9CBOy/2zGDwmw6HOLSCWf+2tfSjud4tf3Rk
2e/JzAbtnPO+tR2MpjebJr1aHWLYOHEDlwynhvEj386onLmXVR2Rd0MTnS/btTl00pvfZ/YLEPeE
k6SgVm3zs95waZWM+7wPCvdyoklG1wX175WOYUB1XXuG7PNzS0CTPnlG0riGeyuQhsZN+u53w5Nf
nfnoixkZhyA+iPqg3eSr0vp7rDkSBVH6UC5JrofpxeNt+CO1X4xp47RONWN2Hw02HGC5Cj055t0d
Ex1h0sYiX4m0o5p/49MV/U9lfy+Gn3aEpqVuVGeUF+5ELEE87RToUZ3y2/ZBczYUmrbDSdCMpbFl
E8yzqIUbzfvZn+4Qf2JQv1Wm6glGV2NqH5twWVet6VvplQ1bpEkReGiKAFB4e3Hz64CeCcPh7IK9
MDkgFgSUpGoGJ0ynYnEvh4S4lrc/72cXWXFYCot4oHdWE8aXtyw6KOFSx2ofDyWfGEAdl6FTKh7B
laJqxlOy/0v111zJwimMpIW0KqbLO/etzuc9ps4ZjHOD4/erWiPJhKp/RSLleuL3G426VEbKzaka
03dAUy0Udwb5bzZwOMwE1Y2w/MCVBrXF+okF6CHlI/gb+gA4pD7Q9tE+WFD5EQ03/Cz5oejnVBWI
d7J/kS4eSTFh+c46gisLPFExLWRSTrmtWzWJcM3+knJkIPuOjI2D+Ix+JGAIpH0YW6M+tj0g2qK4
86zbrTwRUnAkeUXXGxrKOP4M9OQEdg5t7Ih79ppSLgA+oRxUC4UmVHx42M5OszanLHduQn5HcHVE
pRyoHcKiDPcuSuZtj9+2hqnFuTeCdq9YxoMe1S1IRf4ltJKctAIJtY+Dv5R7PeVM/6Z9ff6vAYBQ
ziT8XPo6mpWPEH2n4NglOfhpLlwkp5kfsQMoObo2Qy0vY/aQ2Vmy8OKqckeYkQL9ZH+uJc79WzX5
IfA+UFYoEd6WVdSGI463JNetoZxFyRiToy3Ju4rLtFVlRiWyBMWyXJn9cxYDzxgEBwrstGj0OxK8
LtiADPUmJsHbpP+eePGGZuyrnMQ17c87LrowORXiMnxhjyy8HHdM6RGdwVLLbgO4KPXpAV/u7a8v
y1dwdaz8dRgb9Scn0wmlM9ieJygiMniHE7uCtLBloD/RGhIvaqckJhSkeAK9QGrPShhCzqkjbR0Y
m24Gd9mD1dFUYJvHVkLFQFbI5Q3Deq48TWih8PTW+8hI5dUV+z6OWYkn49oecxwySe0zoPs/xpYQ
+g3pVsDrOcbrkMJpT7Ux+0cStDljEEndp1Xi+Ug46XejHYuBimLox+gAR0DmRPsUqQiw+TYx/sJV
pvu0dXmuiKrr3fSLgA2MvMkw0m51IbOwfQlGR/Jt3qchx0wQJd7IMRA8dBET/nHfmuXujJtqlCjA
g92rVspGW6DQ++lPBLi/Bi6bU1+qtgldrUqirzWpDebK9oSME9Iutmzh8Onc/71CIz8XxcMunNeB
WhNQj34aVG1/ptFSIeOSesAPqML1Urz7pBax5Zj6yje3KxXle6EqJTtwdWXY8ZUT4a+QNE8OwDcX
anE6YjQ3qLX9bYUqo0U+m+N6K8oDzKKs6YFhNctQyPk3vivkxBXpU9gXccyX+U+pJSGWEWOQMtPr
WsHzB9dFtk33SKVWkk9jEk7pxjnMQAAqHMKnCHPUbVZqEaLzLG7fBKrqAiVxb90eZb8wSuFDoxg2
rBCAYXsljJAwnA00HJ8M1V/sbQ0ypxhy49crO1QRG0oGzGI02HYyiEt+LPn4cDpPZssKPiF4QArC
NWYHtv3IxxTqOcntBmAHuh0Ygzdtk6u6eGs2worbHXsxA+XbdhsVPoQUw5M2Kax8kIqtrZafX8FC
UJZLJjwt7Eh5BvU/1Fj2+vAoaznner9p1205ijHGGgp6vDmGq5bmZtxb1PKrE4fp5PiRXfpLp8do
60mGxAQhfgINowJQwEo88boCqDXVeBii2YxGfqcOdj28uCJ2Sajw9cR23dsi7KL/8Z0LND+KA3kP
+Lp8or30Iu1+mVix2oRrU+bmUAaQ0nAtBz1/YtdsMvPbbw1Cp4/1+JxlaGvcIBI/6S6r+1E1fW2N
GtuXKmtDCap5O7v5E1PPwuAj+QrYm04FgDO97wRfJJ9tH8clbIMDEQXlawvAhkRH5j1VG6eSHXHP
oyTltkDRNU5H+/FNYV2ic3Wyxbyyy4GfY+UBcqTXaL0oeMuip4TshSOVZYuy/WTaSFdFqN2+8Ijm
eM8DjZo/NcWC/xDQnVOIu1AIJsEpKOiX8DAd5o6heRQDaP5NxOX1FYo6EkVIYJ6qLpkfQcUpuHD8
z2xPAOTl8sWQlTaFZ0/if/8RVDOcTji+j+bxJbOhNd4ryLv4fFRVtuiZrLXCfYzxtuPM9qbsuRTB
bHps/gdPirBxV4p5uqPClVJEggr0D/Ytr/uxfD65TTXmrQicM+G1tzTF072FBa9ohoHE3XdAIraS
9yJWgqebJIe2NjPxBtaKwuNNGsZO7jnMIVqJ8SBxV7dbFqVMAIje+nuNJTdTu0R7fka0wH4zXVGw
xH4P87etlGw722ZKUobRPpvI1+b5jogJKEXMd0MHsSkuvslbS5x+4oZln38BRFaj90jKE3Tu2jSM
W1Itji2QHFfwaIeZiN1aZyvH6uj7YcahCWybh1LwMWoai5XUBVbfaTOYC5j9bcTZXN6Ugbg8j8XZ
6OVIyuqAsOQPCtL/xmInNS103rA9aoY/1diZq9C/NOnHcGT1eAyhhiKDnNNJPDg7eemdX9pjDbiB
scdksFOwBtT3iEHofcKp8I4TZz0XEFX+SZyF18CdF4RICQU+aycXOeqKpag5fBeTzybTmkr038To
RpkC2odOwlUfrrdbl+5R0kUR1QfOaqw76cdRIeue0TDHDbZ5seH2QVLTQKb9+ojRy2kfAM+VppV4
ejrRNDhLhDFmeNQhdAJamgR8f1UppLFFLmLzKVEBAlXKDhOdkqfVyAU8ISiaaKhZsSOzdJXIcgJI
zuQAWfKF+9IW4tJOFtldTS7y8nV9DZOVTJYHvvOxCxfLCXKoODkVXHpLS+jvh0HXhiMzS9yMJH2k
ctyYyUkqz4BC2OqrkYgVFB/9//LbylBUDpfItkGO/7Sau6qACOv6LGFZHk+IBR2aBUYmV8bFYK5j
ZG6BUXJKCQbOvjCeXIbtpqtW0Ab5SHFcw3CdewAtLig0seUg2pVhS/emy5ea+sUHXWk6tTkeutGw
2vLh0Ycd3OUk15qRxarov06BjQhzv5kmvZ9r8ZklqdA0VHXic6FhjrAP+ARj5RXfKFwgidYzIM5x
ld7yQ6IBgoMLZLr0qEtu0B9Bd4SZywfYM+ZJZVIUqPphXXixSLZoTZ1gP/CbOH+mRjRKkzk+o/wb
chRIZgLU3wgDw/L+Vk5UB/jlkRDu/eh3pnLwQPxlI05eEdo3/BsYlRawJRed/bg5gHFptxGSloqP
gbsL6x6yWpg2COy5uNYMMn6rWVN/YRHjALmmM16r5wRmIX3XN/JwhEL6Sia5L76In+iMJh1VayaR
imJ4QCnwaz0IAAyNTWw3QYOLk/air0VJAGgDz1IersA2kku2Rc3rJNH2s0vtM8UglzztJokdMR1V
uzIpwMJD0+J3TBGRmlSopkF5nVbgUem7mSl9cNwk2Gde+8eEsU+zTkEDRW64PyzsjezB7OaBMksm
ntn83evtHyRjF9VI7PovTAf2gloOqlngNBDrXdzcs3FPREbS3/08A79b9cN4MS1p7DGwmY43qhL+
TRWavByJO0qPZpB1CDvhUQdWDILImHQQx4V509J12im9NTGQSoHiI617d5z2eWW8Nwv3sw0apArK
QCykwp2p9Xis0X1XWrDqH9L2koU3oKp0RGpOMzsnNFe9GlsHNuvhd+OKE+hlpxK0LEL555gbsNSZ
mf1ZkAS4PrsG5/QcXHIg/6mbGr1/b/QSxr+7NJaTWJZxnwvu7mSsJVWKxTJOfoo8ckQKYvjHbKSg
SlyDHBe4O692ZR842u2LrZHOAaSCGJMiiNeIHpLUDOCOYZMBDImR8LJWFO7N8vi3n469CmtcabbY
1H8eiooeWzvUYyJXkWOgq2RgTtbqF/nXmw1V0kr5yl8MTGgWay4ytBzVQn7RwC/aRLb23665+FF2
+4eRgdrsSMTSTdZn6OGjfwQv95qFffRV4VZxYlBBqmYr1EwKvLRYrxx2xhNV16bPZmNWeL7sJL3a
u7uOuKt84rxLlhnq7SoPpDeViZki1PtLtWfGs1s+b7UBAsjY0o9mXjD/Wb5weBZ95xBWoB3xUerM
fzla3RnJYKILaeCWuSpBch08BKpOgShxjLXguUvaBFzEPHF3ds3UHnn8Qaz9Gq22dn+yzbOczcmU
QLAxR4XBcxwmefXl/4kGqrK53mSivJIT4oMJNWvCN6+/tKmyzf12uiEUoilRbgQ1rBOhpyrMWUJz
vaNnFwrhFYuxKcYWtc48vL85P4wIOIDXtnjVoRWXciAfZl6EL+CRP8pCkeDrty7l0XJNd96apfrS
cuFS9li3lfhHK8mV7jC/rx3JrDAmeOtY39EWIRz0Yff0G4psTMQwK3qwjG+cImMyURz+3qPSYDeu
w5Sk5CovTGcCK/Haqt3UYPkCM7sSjv7gGdK4tGrkWi9FUqIrfkozmu59Rh7ovZ4oS7HacKjczdz/
JO28+4CQQTT0YwOnn/2MrN0XGhbBJ0NpaBo0eZzpaphPaickmAmFUFJ161DhH16UpzqBxtlOUErf
vir3IRu13/0tX2vXfvUrCNquoeX43N33YmhIkh+IVyGwIvDwT5vM0vM3ctcMddj/xGFGsSc0oQVo
BqRtSpGyjK//GUcHT/8bH65v3mqLk8sHTazImjJ9HTtHlc8GIZWEt2rKvzQ5XxNWX1fpfc93feeC
Z5uqSXoAcXEwkEX7spGeL2fJW26QXHdL7hAaI7snzsHxdo/cELXP0t57c+u88Ts9oknrtvwNSlmK
1e5vBW7GBxhoSzCXPMkw9GLUCAu9qCM1teRfL86fEQUzjgyKWGRE6EsZl9V9m4OphDcXa5YsglGm
UQ8F/r868fpP4Xb0SMOl7q5Ea03FI+gOPNBidFOBI130YUhRDFSUs+WsQ4ydDyyddX1dk2ALup35
1LHJttOKhCnAeSsvesppsdYVIM+bR84AV2crcmrHo266FGbCYA1taJXdT98tkM5JPEgwQdkRJMHb
jKp8cxULdqrfZ7yip0rkMOmIvuC9oCdC+ccWljInHC6O4EELkDWujHU4O20d5YLeCEMG8IQjyNJw
0VluHp4VAmAzmX7Oc52M0MGkiIElISTbvZr0YYGwqjMa1lBzhkBdhklfgsVE+B5nIqchHX7rBeuk
UOJJLT7RtKRr/HsXEnpx8Dwf/MnBqzQ9W9saR18LWVvgutn5f+rgZG5YkkBwKt0hXVeFgPBf7wC9
X3gVSBb7C905pW3f7KZM+vzfUQAFeT5tnIphEIe1wQh2GtoRpk6bbXzDqvDf+2sh3J1ZkzhldlMs
FKck3zMTiq25gr/z2Ews7Pv38sHxCYisXZJ/QzTE67WcR2vMUdLK5Ki806KtKp0/BWyZu6DP/kLT
bifpqqZIfP9d/RrHDtIOVZ1Wd/6zbCOK6roQWfOdRIII1p4JWML3pZ/s4unKggi6KAeb6N8iwW0K
q2xb40AwE0IikHCfHfHs6v9mCiRalej8T8+f+FRpYjY77ZzEqqojzdSKZq3jKkVp/in0zisx7ua3
mqlVwtd5KrP8q+x8EPO/MUdxOrEeTkzuQ+jn58236LP3A139xK2X5gfaDzUzftj1WJmcG63E6Pc/
0FQYqvaojjvQokVe/5t5pr4OWoLudIFmKm+Ea7wv9B0lyYfFzsf0esnDFURv9IvcMJzDneHfxV12
svrukamdTaXW5CPy+mfLX+1PGlo7FDAhyV/Lb7oWWUJFH6pMQsk8NdPGk8chikMhXiiLxMUZuvWS
91pWJvEhsBxlme1JQR+jWjssabfMN3W5j2PGPOqkbdbu75yQLovrvAi3oW2bVnMwZ1TQCYuvo+1X
A6aDKJzmPEA2HkfpuG3nB2VHJlCsOwjzCGF4BZngwhVM0THW8l0rFd21ml2UXV1C94eMVLtSviI9
6bNZbCKRUu5vBhFAiqGz5hQ+P7IimfA3EZDEoDPK7cIPoagCZDn87SwobvedLZ82z8d/RNg8ODrL
HBOvd2wrH2ThQy3U6wPDyn3q1BpUSv9fN0FmB8wsJNWsMwZ0EZTI4nuU82l4zplWT9ahp68/v94q
92E9YsUEdByLEgmJxzUHlQxlleuozLI0rZ9HYbB30LyjhUgbj3ot+KOA3LWzbBN+6aCPkBJCeZA8
HFDrJs0CfxUIxs3bJEzrZ8FTJBvN6g9dEH65szckw+1rLwhDr0+3eNff26kuLDO/KiloHOQIv1Jc
wtz0inK9HMcujZJ4AfmeI4CdsNqhfaKF1geXL4efvDk22+V+KgMUmaZyAbewaePeAAgdeMtQy5ND
FpAs1AKbfK39LTIUsuD/c2pkGOy+BmS2R/05ahUDGxQ9RnHc9Jv1iEQGGv3UjnVmI3B2I4uAQ2fF
oYQJDKROE3k4Hv3JKntq77qijCqe9dC+OpA9afoagHAAFXaJwM4zVb2PZSdF7Nbs1yLDRZmo2Q3Y
b1a1zOElSSo34RURXF+cWKcAoi7osOYT+2cmyZwLoe6Bnqn8kN8rQ67Ejf6FBlNtUG54V4HXR1KT
fFnwDH46U5qtaMZnPyDDD0zX8PdZPgGVIEj2NBqeaD9C5F9sbXzEflVw7aKM4aN8EcGK9rxfUV6a
FgNwwCKjN8NJ368YPSOo7O8tYoHJ/vcIK0DJPbMS0BvckK14msMzMKTw8ezFp7HBtqQ/ba7z5Amc
zdO5YgeEJU/kFxYPGni18wTwS6XNtUyWOzopRcqcLxL62A7GJJkP6bZbbomUOC/40qIx2rkRQ4k/
Kq+HDobM3bYeGs6MMEK3nxTq6OMKmQ2ET2uWH1QogmVFdd8VNu8Hai6sGZu+GCwvt4ziwGHRVAoV
GgzMoMrTd/NNzfJWopU5FaM01i2WShv7rWOY6a7ObN4YesHILCuRy1MiYKzMJ/ee2aPWMY7Dyxup
QXYNKtLLsRiwJOVWudLFdDW2Gr2uqvuJTPWJipQ57qleFBvsJKfzV3oWu8e7+FcMDAvlRWTchmF0
sb5uvrieazJCKZE86TfaquIUXyZ01blkkw5NFr954KMPHw6gJAR2p5zQPzACYkSlNibOfCNe2XK6
Eu2ZaSuKR7tSrvff8MQeKm4AoMXFTEhrlePna6oYibU0Rbu120V/5vNqx+RE5o3ZkrQN/NQ32D1x
mt8HhkTEcVb2GUaJieViYa8EA9fNvCavuXwgqYeXxQ5t7LZV3P21kTx2tMupjCyY42qgKYKV0qAB
uYkFa3g9TUnbnPSyWcxfhsFNS3ejLTQOvPndtrtwwYgzh9CbOy/jgfvvXv5vFjuxiqqygIV3Yjcg
yChoH/Daa5xi3+BxjXXpJCqL6A588mAQZJKnekoLnMdBKcFRR9qWNEGpU4k9NFiBHo99Wo+4E4t+
JMD6bBJw2BUsl1WNh2bc+D6fu3reBDg9dFowt7uRuAbqduZr4WQr0QkqDGl7yN25GN5wdBQjwGBG
kcfo0R6qg82M8GXHFcxEXSpttJtffueQJYArVkN13YIww1vDliKl0d1eU7jL3JFfdE5WbmpYG4Nn
dCeEiq+LA2KE7fyUMIJxeImMokGHoO0954yb1yxQlF7fQjkMh1bWWaX5gAYtk04FQZveREuSrdU7
vuVFVRaCZTZ4Jl3GRKBKUt5geJKUBTjWAexcNJPRSs8vHbQru8XUPEkDYg48EVtxoQ4smhXp5CP4
1h+wW7KbawibrDKAnxdkoGj6RcxLSpoKX2X4Hx0XuNiZLb82TXISk74ILx7vUY7UZC6WE2Fp5Vih
itVaBDO7C2x3Q08SSWNA/fERPZ35reFbk9db6xcmEcPw9Sx9TrnHnC8xwCN5keAAUFkCouKFLVPF
57YEJiSe0uBs4onzC522Jo83JvwEOIywDvZneuzcbcUVp8G7a+/3xOaIYSl6MRAQm5s+/OvAjbKU
Fhpuhf708fa5ntzHCJDPdDP/wZ9+fPKEVYIpnBfuvF4c2IIxzE5HqUcZmPmoWOF/wENdzfthEEJP
mqkdDUs7utWfwNiEvelGcEfxZ2CBNTG3xSkiffZdTAGdzXibzpbOpDDD/dbGEw/rl78ZofhVNQ7U
XjSNKkJ30qLTt8o9YW9Fpt2iVXl0+HmGpmbxNZ3+VXE8fdnntU1bB3d83xokIaJw9TM+AyjA+gcB
vN7O251/w4p0sZJZG8yZobU9KEuvLSLJ73+5ZPNhxxFPhp04o4K+SegP0Bo65Uynv7VUUoS9PNpA
WojOUt3XgPq0BaQx+IamjSb1PBCgavr0mW5LipwighuzROi27Q4YTeUJge/24qoDOvey4UnMq9Sz
cR9x1rB6+d9jK52CzceESO6TgajpLobbH5N4ErxQ14nzy1SKeybXxTStKaLYF/LUWc3f/RKj1YBf
MgjRUDeARD5R2woU6PTbwTgUVe0O2fAGQjkn1jEmFMptsTdf65JIQ0vaqfHPwu9fA5SpVzLHps5b
LaqesG9lyRHRRefmWBSaZYJjp91t/nmYKoSAQoiTOGTv1vPizLuva9Re37fjT8GPBSZjzrrb8dPX
NqS4LB03uQ5ZWCrEGy/mCPWSPaE1eFV3NOPZKk0XsxJtBWrND9kx7p43jz/XX481TCRKShEFuxqF
L6BcKvA3b/d0btA0zdY4LCLlKYIaMjmFwV2zSDHyunQy8Prg4eV+5renRBgmJ3aHj1cH/ASv3tdZ
5in0NGObUlcLBvlGkvPrhLwzqSgfJKMW/g5s5U7x9jDKPHAq/NqHIP2WXXFJREpvmG2WjnQg9Wvn
OTZsAAKgEQ/H32ny6rAO6xX7bJ8BYu0vdAhIGcMOfsYWUfTBR9L9PZnrshm4+/TqiqPZdxcVa9F1
pIG0lXBLqfwcOR+X8OIQzHj1yuAC5RYQvCfI1KSIXKm+ZwRJMPr6ygLcfHqT3MwNsYUqA6d90U3h
E8ZrV+HRa98EFCYJaQDIlnwgdLNayaxWQWAlkY7MdMAvRTrLmkd3hrcCGrFg4Pdep1FLZIlyU/md
LJPx+wWzr74i5SBY2w14yI0jXrzzaZRdfw8KsJJ9Y9MecpIJjcP+Nt3yxSwllyJmHssiQPBSDVfB
JBjcyZtoivx2x51hfVihp/hgDEU28qg9RtmcWTbNCXRXeddqO+/gEDLvkkH21f9boBKFa60tSjlx
Z8xqwLFvtbVRauOrJy0cUorCI2vCk8bELnqW3IB1Agez5bOY9nVHDz9fN0wcpbt+kGS2LmvnPkqc
Lk5R4TbIxaIa7xAfPhjVQnpvLOWfICjf3RFYHd1ENaxa5dJme/RTOj4F/QhK/k6urhOGQKQuu0hf
3Uig62Qp3MjusmbF246fvFFgaPLXZKOuM53V4mI3Xn7prYb5GUBaK0Zj57Wizfot1D8kGsj7qL9k
0NvdtUN/Oc63C+niIoEfK061J9XItPD5FVZQvTPcNGb3+XEdANV2N1bfhItzBHDUaqdt5Ouo29fm
hNugUwfgAUYtPmWyDeU/D+GWs2Vm2wSQEiOweElo55DS40R5ai9L3IyUNlNUAUlEXminoWClMHnt
BrOQVptXxegq0Hscyc+t8Loa/EDOI+QPqvPgHqBes3ggwTRU+0xnx4+FWawZZKiR0PNNsuNRbrGX
yL6HJOQfGBapDiEV3pozccgl53Wb8s342ufIgr1jHo+e4vFopvkHCtr/lBJ2UdPMth6e70QD/vfK
hqTiLk9EjS/GyGgp1geYFKvOj9K8+jMWv+qZw1f69M5q7CHGWIsiviDAs6AyCPFdpf/hNP6Ixdcs
pvu+rWOx9b3CljP7LCbl4pTriQgDwZCNAkiqIcrcl0r8hz/AUl3VXMsjaEKfwNixB1k8RXLQSKK4
1ZWHYG0xoQ7qpkvUoZBo1lc/o4FVn7MDJepXKoxs0ZnTe4md2tRIPXDuqSalvGonpCn1+32FunWR
8nyzLWMWKBGz3rWWNgCJj+ukf5auSY/3Jdxdj+3x4hCOQTWEEwN8jJwB7O7aYJZeKs1erJ9iDT6h
GVZsn3W/Crv35BWiPxZ2DU7NuSkXo+9vI8KKwSg4H6JzxjWzC3vHd3fa5IU1DeN/c0RPMI+sgOXA
FkFyu421IASP/3g0LS8pXWNLD89UL+BJC6KOF5H80F+Jfkd3KflhGcrh4SmqhBkl+Lvitir9nBf2
i3CL0227zuH0+dSZQfQyuij1EC9JzScDV+b4mtwLewrOR5Vhr+SQqLy0oisEciy04WAJDaxn/VYd
JR21txbxhrT8DgMHjcoK0TNXg7u71zoooZGAFRu2hGaOwpARyq3F3HLKhCUXWhCcrHnuB1aOJ3T2
7IRW7K38yMT561Fjboyqrw0p8EErmi96iFyStfn9AOcLVGj7ZVE9huz9m9lEYKz34a4d+hw9wY8h
jMlZrriNgfZG8esiSUECI/oxrUaIVw42sh2IRu7KCsj/WjB32awGvs/erQobkUDYksnASgWh303V
YLC2w3vU7v4LwRXQgiXHH+KU1O/z2WNBmqzGnuoPEi+cisPOTqBhOg337qPMvJhQzf+LlVjPgYPl
kfTPNeTXp0PPb7CDgt4qsz/zlN0NYCzfBYXI9gzJJZZGhyaKQEKucVeWaJJBbN45Il9ypUvHK7i+
j3iYrrW2xOvSXcoSHzLl45d4qFIYSnPgpBcuqLDw/blVAcTiclqRYF9nw13+JxTY/ssFGpJDIKaj
kaowCiRooisJRJTzm+HJYflON9Y0b04nefN4tAunkKVvMt+xuU76vMYIUmg7g02y//EvF2qoNVlC
+DX7dwzMhhWEhloG97S6FLwUCentUVAbewYAoM8DdtG77RT/jauzv0GBkbtgx7ANNG408zT4d9Ej
xYX9JWiA68IyRTgwGwqYrFtgWgZTjjcbZqyZXFNfKabQUkeBZUB9/Imk4ws3CZ9qLJvJpsB8eWbL
WuRZTjtju2p98tUyUeUzCf8EcHXAkiNKKTuSP+NBNIzRpJYp0UwAYQM2n3hlydCmjGqYN0bIDvyp
SNpf/vUhT80VHZRmPMnv1toc5ILLsGvCvf91MkeGu9H+JV1m+BWnbUomOTdDP7Y5shcQL5KnmaSP
xbVSB2TTptx+rtewGSd1Pnhhl6Y1XNOHQEjuJQmddImkqplDdY71l3O9pUEvOntR3QPRua7s+Rn1
y00PgSuagStAYmE/RYtVVysolBuEOrrQtbKYmoeNvU1sRC+GpJYi2GIZjVIDl0nosi40x93OEU0K
ah0T6L9xOxMze1U1QkU00nvgTp30sKPVC2OmS/FYSoNTHUlDeJehSQdJWTNzjrxyOVhQRz+EauZR
Nnf3uqOkYlVO79etcK0FRcltKRCbXNHpj/hZuIFarxLq9nYVrau7i5R+iKxPTg7Nd1OhCuQCu1Cu
1B6LnrYUmCw7rsQT/2bqf8F5czKBqL8B+x8faiEGNGYm/h3OxgPs4O+Qz1fAAjSjo6zS9a1b7SI0
NpUDQOx6cbLieNafuy50lcbVoooz2U1Sfu2m+ErCBBRctip7CYlNZJU7M0JSCd89z3Kil/m/54kE
jWr3mBJyTr0Gm5l5oXQ1VIlVh5O6SxKmAnQFWmgx18tZwaOwj6WMngPS/1DX4sZWt768t5cn5d5K
j+A0QW8lObdIQjz0AbOO2afxGzOCDjJ2Zad0aENTXcp5j0Mhf3zY9JGES99Fjt0dfKDKErEulX49
rmX4w10PhCavy+39ocjMe9n8I1AIgIC/7P7fVX5tOpmFZlOYoS2/i2lpAEJh9Wz91Ptrk/2q39UG
bnCsw3rmKpm3rbpJDONSaQttnLtMjgGEi6qyy9TIIRz+zgCMlqQnGUXFylYlXfGqjSy8Ym9imQ/o
bZfD8uCwLAfU1a0L2KeG4na647Lj40sub6JWrI82UYlHtftbrZ7C3SUkx79Id8x8TZIlUG8ZleKA
1zKIxCSNv7tvZG1QW7+E9ub+AcVM3K2A7qPgP+obrstPqbF9nxY6BX/eayyYFcKJuarM6kfjkTRm
PRRNcqSzUkegtcY5cKaJt+996lomk5H0vZx5QDZrxlWbFt0EHHKgYLLPucKTeJA33ZJ1fZ/NexRN
6NTrQbtYtvBSL+fqTWSVWr30mmlGEsjaYpEGQ2qNrY9luLKtoNTyuU/27OAiBUDk36hOwAA8YAvx
tmL0ntj49mGCAakvrWj2gAsdqqCkRa9iFZj354YJ8XwK1wTo+3BUaqd/s9JXenjvm5f5PmFURunE
CyIUQL3phJwSFYHhk1iQm3j9qbdGnuex1PQMKNqkUSLkNTHIkRdsqbD99PBaC5aWtX0ATBFFpIZf
VXeUMy5kKzfWXCCe8v9c2MXYtK/iGW2ntgjZ7yi4xGYzpIsd2wbNO0EENuy/RRpqCKyqqC7vKiE8
Ncf/FRv0qlz4HYzeht/xxNRr2IXy4B5h8SMYCRzjlsRaV64e5rtJ0T+yCEfXq3D4Xe68u26P8GAn
NC/rcL6bXqPUHBl84Gkycn+BXWGhXho3mYinYWDzStPeU7IgLddzZglp62Wzs9kfbVXlxVztrFFv
zrosyJLoTt05g1humHSWcz8zUWlEemNgU3wBPEjFcRIU2Rv/PCETaj0/GcrtaQkQ6D2L2X+d7iVm
a1Zho0g2K6L2aP/eJaQl7OlA9P0hWd8i7jsKgmY6JUKcCHDjjfXPg+IAlCfqypfibJm91XtIcjcY
LBQOTwrlG+k+5f2/Nw7KGtQjYM79oNWWF5E+6vn5hfPMonOrKp1fJNrkgKWXP166ixX/29UxbyRB
V3iFr4sBzO/QiKQUNTTUbCdJzzBOIjoRgIO2vG+HSEMtEMwtgVa3W/sCUVRPsNRQe5cMTcdSW4fM
0IkIDbqroI3TM3GZnwaAuscI++a7u1su16aonaMMq1F6Hv792lSdKAw/sWZcwFp2DP0hOIbBzr7w
3QWOxgqiNddhAnSLW07sjV3G70xVQ3/qTuHsRyNpk4eSWGYa7VbBiGt5/6Caw9A2UoBbUGqbJ0zU
EjouVQsvsikmMIl3ZxZbq4yED75g2mUekFsVd1ivSk5Ub/1ymEj+pW5hRud0Mjny3iLdkaopGWQc
JLTEXWDaUMa4Xtqz7JeuqsvWORmcz/bAkn+bcd+BQ0Ws2W0Guky3eX7N9ZhBbKGBY30qwCu632Ee
QcV/F1N1lrKGMHpjLPCcZ03x7+agLs37PeeGiNRRaRvAeKRYJmXiY/Khvuf8cLOg/xmBK50OUPWu
YKXxPvNO8LxKeNnvgG0bRDJXq7aKg1XuOGzXG7U8+4pnnvhBwPC/XTHTPc297W8IT7pRmtulwhZv
YgNZFLgBp6+SMDzUIxEbpu/f78tEgufnRetxj3i/Moz8BdBcf5CoOWZCsNgBY7Tbued/fpxG0YCO
5cyrbvk4ImHP5TRFFGjCHr4yq26RiAd/Z8IUilVn5FHziYqa+q4xLE+NWKbITu/ANoEDN6lifkWc
7VpznMJAAqT40G6hy1dD4kUPbGAdFj8lGkGtXkHbPQsw/L8Yr6q5/XLYpprFJWDLEV0Z6kuXT+qh
sGcNZJWLYLf71JGFYbeVke/3R8Yb+DMK0ClABFzDjWL4avFbhmWWA/iZicGJVoTZlvJ3i6tGaXaF
Qes1BRZ31ZlcUQn7DSyiXlMWyPoB0KAj/uUvd9Zij2Lp+DcEOTLLQRBIEclMa2kqrqcqIC2m1iLH
ffogShHj5cwML8WoRIzGLui++xWw0QX3IUJ3YKw2yuuKaxI9lHrvx3ldVuiua3LieHo89hjOLfRL
sg/AhOfDSYb5k3CWVq1k3Qj9MIdbFo6Rp/Z3MyADdoUDdp0UPi9LK+t0l58K4nfIfaFLZtThEm7G
5QxHoZkzmZeicT7tiZ1LSJDFE3UJaf7FYt1V4yx2HYhAnP2jF5iJqKTd1shvwKIrp6eYG44xKNjc
InKfk8ID5hbj5z826eGGDyjspJRBs310r+m3EsGL9/gyMgSk+GdPqls2C14edTSdn58sgE1Bjo87
IfyceO2NUbMwbZOt9kVM0KrUgnjCUnDGXiMOebwKYjHT5GIpcWNOQ1G6coibKn1dCA3jHKh22+vB
QlrspgNeLh1C2Dktaj/J6fHkmCaC+W127WC7FKpKVU5szYx060sbDa6psx456ZoQChyTTX0sI/Gk
P9UrLto5rqQ9SNwbNpk4MfZrKqz4D/rUGrriK5P21eAcJscpFC4owWM0Xzor6D2t3glcHP0VGAW8
acT3gYKirGi17bZGpT4o8rCw6U5dbspooU0LmlN90xWkLyPp4vJ99Wilna3ye4kFr5KD/6Lx2nCr
ZOl3nIGlowdTlOy4B5ImHf614FMAm271r4AQp85Ot77rB/EDInqQ+Njr3BdOh5HOj8D51xw2Keuv
hejpweWgOFXt/8J0YjL4VNshMjdUOxCbZ7g1SEpe5bJUFaAaaujlA+DR7yJdsGdqZG2PMJmGaAaV
aFWrIBJSOGqjcyn+Zm1nGzu9PlXYuYoglqWdXji5MwLntXyuO1eves1RLMjlZS4drQqiSJbLBG58
OpyuFORzzZ9ahE6ohEOl1LIfLloeHTD7i6UhPHZNVn/pb6dBpPg3kUeS2VKAc1gD3kt45pgGNmpm
mlOOG/D7msOxN/CSKpT7cUzJNfrT1tfRDqFELBYWkLZZnRrx3+5htLOH2HA+dj7bA1kFhWO3gB5A
23OjbRfm3uOupEJLuBomShXqkOkc2ZTGzMTGvrS9Dn3FZG4AXb+fy8AAcTdBz+6snr2swq+yRhEM
1OrBQ/hf+ZfZsDV3bUfBDBFNS1Y5PcgT6maor0ocX4qNyhnw/Q+2sT6mk6mHYZaFCG/5g/ZvRuWD
+hKWW+/mpt6LlcEe5r1AAyLlgzCkZlQYAD8XyGzB2dMCLvaiojtGCkRALPX5psAAjpbj0Wl8VsU+
xHrnWuqCo+oTrj+Bgkf2yQwj/CKJGDJAsxTGHWsiNlRIqLCNp6UFwT9IybiC/xst1ppCxNinOLgQ
elPDlTWzzbV8EokOFLlBHu76XH7xyABSvpNPhnhBUTXmvJWc3iQztEGU2dnHcErsbUvBqI3+T22g
1JOp/xpwpB6WFbXjJaxNsHVZElsqwqLRkkO0rjfiEXlrrl++ASehlb3asPJ/Mjvmu4kZuWlPpqjw
2u6+B2kfr2SB1SZ7YMAaLLUSdfCS1X5bOaBZWJrWcRbX4l5j6qAbrwWp/2zkQuIdExvdRMzIwHP8
vC8epgp/bOdZJKMoehjuIpzgGxu9fIeFw29bwa53vwmMyadDxsSKmkU0ot5md14llMDBzGL8g+Go
4eYm/zQ/lrA/T6WdlouuSOCsV4+XnDcojNXuZRN8PmOMHrXVhCLPWZ4MfeZOBG32ZBpEHMdZ1vDD
0byPQ9YdmCsOryaIHk2st3pFffnabDVFZZ4zrM1FtEft/Lnd/bqrmhjQblgNNRegQ8qJQcrPzFfx
5G4Zv58DJAgsMPxtIGXfwoQU6OK68SD87d0X3Z+ImEFBe7XwxPXZpEEbwePs8OouQ4oItPhgJ9Yq
FnNmSpwhhan0fT20YO4c68M6i/h14iCRsZz1lcaFqYdbpIVirwTIGgYUn1hPETZfHpLxLPxwtlPp
ZJ4nTyM6t2TSslTU7wFSgITNnUrcrOTwlvlalJQZGcO6rTU59EFWBjmJ/tzfuRNhxF9AAYfJ0h8d
0C9bg8C5ML0i6klhs3Ft9vIxJ49TAdfA8DdEo1DG3vL2G+eDejh5rS37GTXZNG0z87fwrZ4gzity
BXHiyzBXO3m1HwRtFXHPiFy6qgPUG3MQz8x9VM1QLz6ZE09jj7X2jSnuS8c0IMzbwXJcNcRh7/LC
ObCiNc+iQRHYfJ+U0IqFPvoaKMfL2SqomAW/XYpertz5uOO0rAOdxwt83qrvUv/vzfev6U1pPuOx
g9Kvr76r9FPZlVyDXyX7p5bCgZR29f16KxUtjbxGvHYDrk550a25ZX5hsd2QNWBK5K8dVSClj4lE
jrTaahdxIWJIApfj7lc9u3tZyimskPfULYekBzpHloZCIo7W/iZmS3ApXSPGb5KeGNZseAO4W79c
pJUJXqpOtXy7AP1aZ1ZGVKItBqr61l5VJZK8GwWtvTQwjPhuD4ULEbtau8tli6XSG2pmYXSmSJz4
5qNayQt8Co+tQHsPoe/ZLvzyN+4IbJ7UdnHzxatsFZEmsKcnWPCOwT3bdODeQPs+6U+jwQGKiWPl
Ei2bw44/oa0iYuRFrgXYf1JZ89ffftn/yfaf3gCkTP19eDniIrEsHuqqSvBy9ianN5X5EaNpz6uV
tpDDEIH8njiIMNZQ0vK7vgKryO3uclPwsCVufpsgC4SPGvKebfFtF+qC6bTyBzpgJ7DY4UPSDqB0
DdxCWIYeAhXfNUuE7fx4MEb/GmPWh2Rm7LLzEkbi0bYa+wGvP6H+05LhvBu9jc1j1pyl0VMEMlHN
bmjg/aIl08TrifvVvLCMXk3ZfqNe8Bw6/MXR7EnjOJE041oqZOD2EvqVrM36eR9udQNInwbfuRHf
2SBTKPVT2nEBrUWI88vvCt8Q431Px4Nscp7P7hsn1syiYMarJF97qkw8yliOno4Qzk2ejIV7BNH7
RQFapr4wzYfNANN8xYqGw3xyIBTPAqPqyE4EU/mppZOzQ5fu4PITNkOCQIGFL//e40D02awIkVZ7
cQHDqLuvyk8A/wOl3KWmC0C+A+On2RBF+JDrJZ18RsFs2rqinfTa+lDuDcx1yjlXouZD6qTYXR8Q
/pR9qS5McaNR17nO7jG7u5xajIgdjaQWA0eKNJ9nZRdGb70dOSA4agvWJa+4Gk4W1J4TTW/HlgM8
fcKPsumzz2nr4H/2NbMD/xMcJDLh9QD2DgRFIynGnexYsjXGp7kzOZPEN9pO8pz3bPicVV9fFFhS
mix8RgdzirGEnFzqtRrcD3SNyeK8I1G8Tl0Ab9k2PbhPvMSTrXhLjUBSOSGdNAdlPEPc2m8GEV58
jrBb7O4ackfsOIZa37wsz04nv1Ut/rTLZPoheLM76Z+SIaze/Ar8A4DDACbqIcrC5bZMP6cxu3S1
uWb+nTp/mkthSGa9dd2A4MTv9oZV8db8ab311iL6BN8xocxL3fe3OEz9ghWLQX6KP86MQ95QXRuo
2OTVjQZllhxp88+Ecscs7PkV2dYRCHsD/CKGAHnR4uY8ZVbFHrvNon0eWoXFrvvYv0sju3S3V3i6
6lTq31YNI5usnlTlH/wKYymR9aNo203WIYnIvO1xGyx65KGLyzMeSmPRr+TalEEuid9F+cJXaXWz
oXxaSikgBFEb3ILOWv/BFbJ2YEMK9kxPVVRzyLWg6RsCaihPgGF4NeDSk4+hTJNtDDdo6xhxgJbO
myPvKJ33rsmrFMODyxOPdfr6zUlCdJEktB/9lNPQjNN6Ct8BHFv8BcO9A0qqyvKnniOXuhtoI5rJ
HQqLPtdpuhswRJQ4KJDalyZ0VX7SxkePsTYkxznWRkdzm2xBLkUxy4ysnk5Q4IPUYb6xYmi8gm1Q
NhyEDa7j5cTrOPk1MEQovIKCHDVjJllhj7q+4xUvXIzmmskdHrFvxY5tpz9o4f3bGNVHpFX4P6aA
Ni4zEewE44S0uj8NqIA1Sp5ODF/wzo+6B1MdO5OAzhttO5qrVIxqfLX56D3hUkLGlNvf/V5kmths
SKleGG032GC2UJYre+9Q7D8CpalN1gMlGQjfAaDhlsNy1dbiPgvBxZZKPElSozPb6oTkR4s6OQUJ
W5Epmk0RPQ4qU5u7C6nDRGnKJ2G1I+aNeIhuHjcfFm5DTCN/fUvTVWYZZ2mb/GkWRUSfyW6c43VB
zZNXU8hgyaVre084jUQpRxHk4QR8AFWQIHOaW5KMBIPs9uNUKMs9kSJuQlCVjRDk23wmONhTEWyZ
wWFJu5IXZHKzJ/9efD5W7ylT6fuRb2BaEW7jkIopun/IO+0iVHgad5685k2IzE1R25iuhYXjNpiH
7gWEPEQOqcYlBiN64zHU3qKM4b65RICtormVRuOY81TBWv8yFNBQRBVT3T2cEmN6v/oAc/kFDdtw
Ge/UBFfHzD/3BXEsRw2RWWLGKBMpbuoCxq+/c37LWKjopeeLlVtPAK72vG54212A9+dOV/Fpfjgs
9tV+9PaXLmFKuKZCoQtBiboA600mDPP0ddT+DhpnpqcUbl2yPiPFpj7s6xNuz5yUlLcc5G+hZ8YR
Wsjcl1udbjcE7Nd8thp4UexMMnFC+O8LNIXhuNc4YLcdkYU4QToZed/2p/Rt34gbekMJTaO2vkL4
tPPYIs59PyXAFa07sWg82xizCNN1T5goVjeMcPYolKZGg5sKU3RhmcP/dNBvX/W+LZom3IYGlFjj
yu+IjqZj9emECYnZmbZmYka/SQvmArkhltK08VhxfwB+ysk7IVd85zPqZ3gQRTYQnaDOJ1qIxL3s
40OOyJcH+rCGPUWEzKMQ3rIRwOT/CzcPvTqiOSU9IFajfZE+QHKbExhtYJPyo2xxJmVPf3XBIpbx
nYWaaQpQqsDyTa2Xw2xgkNAH/bFe3Hwk2LClWhiFbDc6vy0M0Rl8jbwX3RSCF8RlklL1P6zMRiQL
iueZMeD3LCJvXFo9wLjAoXYtNJopyCkJ28MdJkZ7N5QcBEKapCX7bTLeqY58vDWXxqu52N7P8GU5
JBczUVjuEIx6AuvyDz+WDN9f0WrW5+znh2D4C+/pQ1v5rvY/jldLbA7Op+kkYewmbK+Vfm4iGgat
VvP5yNkPmUSDNCbku9bv4czu10f2O7aGzwViMdDnr70ygAgdcjwgu5sq1T/1PmrdK87MaaEyjezV
XNGfF+U/EuLszO5r80LqoCZPJf9zS4txStBLncjw8q0+1bKmLAeEUc0vArHph0jCgnunD+MYTRwT
IxYYk3lKDa3CZvqGYRt19yD+ivIpI3KnjLWykaFibG7FxhQd5Gqhwjz/ate9GxKEn3YpNXCECJ3F
zHAfYumOeiEgS49VuoFE1mjWoz7fjPM6xRD2gTzCX7dng4KZcvXX3rGIMfMBYOaDZFK4kcGRTDQc
yFL/CS2g3/8MQ6IpYl1kXGeRL40dvz4yFlZ6RmfP6tplXgauFCghVXy9ShCular8SV7jH+ZI+uNq
wCZLLe2Uo1QTQVxkg157r+93nvyA1SBTNWlTI6uipH7LcN8pygoPravivx9d4Co6A5nvkRazBCzo
UfY2Op6JSJJFY8adnlnNtfMkHh6z4ZwJFqrMdTsfXgdewJMk9hbD3F3lzPU2avgk7LxBsU0nn9AR
LVndD8mKkOQFn1qU/fExPURCvG1afAOwpUVgQqrZs1SjCTB+n9N3lT22KwSoe3BwpngK9eZB/tGD
k2DojLi2W7e/ul88qQfIsHGNiSMBgl95eL3WEURGytBVwtfv8KcTp9gTOT3JYrQNbZFuUhdO7yiL
QD//3oyV3sLXWbTCrKAmQqYdp7I4TEoO9e4xQYjdwNoSsJRBQUQAJ3jZXfEPpZnNvaNnlxp6ijz+
VjFJigfJ8nTgjSUrkA2tyCUuerqQh5lmdna3ARg9ROQJcZ1zl+1QEsues3D34up+ns+ryQO3hbl7
5Pcos3gfeSfHzBAqLLR6lqB+pAhvX6DGU9ifP709vPQI2VJVeYpRJMzjjo4zDSk/X+IbaFVxhe2C
EF8F2ojcB/mLjly4tdgxTDPHCPW7K3+Gb8bcH6pPzSMzNDTeSKbA79gSFyzwGtJl/Fw4TVMDxWyG
RcsDlBqIFgpwcqlBMbBYucL2Mmfiw7GHIU3i4g9dYRCd2UCrxZqfjMCcYh2QCWDXpgUanoLy3rC9
B+C9f2cyNTUhq/TV1bh4qYSCdzIT5dizRRwR+MAjP3IvbcsvplgYNRqYjrs72ftDrKAKHmkJkkdL
CHD5blB9mJC1G12xOveDhoAeMZcuayI9TpB6LXnIslBPKe9RlMwLkB27guvwQGWtLHAmr+DK9eHz
E7TzbVYpoIUP8mbOwoYNQnbFr/bof0xW4KftSkuWBSh1wrAafjPbySwaYkJLQ/YHxa5VqaSv/+a4
roZrYe1ULbGlJikYVTt7WCMGuI/PUSepGeiNvXan9QsU7J4NtS3JVZNO2ZvCLf78YStlyymrzC0T
kInWRp1/refoy8RAjJp7Mp7pbh06TnmAW/9bSWm3uYcLAt/RSp83lFAjcgLG540K17DnJxApDGmp
XQN//kCDCMngIhsIz3NFIHNj2Zu+BT8nfRB9Yh+SJnNWSNE2Rp3B9OPwVSf5Q96qRSmgAULtnx6k
go3VFIUAzi5Xwlu7K8G8kOS6JDyKWwuZ0olCV5I6ogE5ncri9rKgUy/GRruyKT7WyjJOaE0PRy8h
V5zXL21Sk11Qqc/ihJI+2TSbmImPnsWIqnwNgfSwGUihJT6O5s7ic6SQ3y6lNvdUPCkvb22Lng6t
w+1aXIrGs4GCk5SmTPix0g3XEeDltInIIqnoJYrnTNQyn/4G+q21MsX7u0tZ0bGlkp/T2zgUdhMZ
kMe1OCdG4/khbz8QNFusQBaVw9p3y10rzQsMtmBfiMwUxRUygf4OIifIXNI5CGuNAkxWgf0yVird
Ry5nv92XmWX+HSGW/HyiDQwbmeQPUarcb7ScaRFrLt8ZofqlW0lq9oCEEcgavHPSJ6PaV1sm/qpM
LyeCr0peZ1ebik8C4gad2dRb4T3n1QxfQWeoDCblHv2mylAjcs/6GpbMCb16VMrjPnSv43nTO1t/
CyNXaKJnVv3a/w4sXWml80O6g69ZVgjkkFhpqZii9SWLxSGW/YIrQG72jbKLq17DalN77hRffG84
G5VsENB2t+IBdoZTsmFQACCsuXGaMVFuw7n6Lom3DpSeY7gElR2idwm8fi0mWBdsM5hJhLRxLQPl
4UlSpFx/z90XEo3XExXhTER6NQ0Bp/Hvo5zl3Ub5xH1yzPhBmUrz/U+qh8kmxyXJGQVLuLsXvfNC
lV32yu99OdxZxr/wlAoN1HKrUXtE0+0/Sa5smMMWObwanQv28aSgwSnlbPXSsK0ZrkQhob4MJoQc
yon7Am/bYjigfVNs7fbza1f0qFRua7wm6B6jcjt4L1wO3LXB8T7MwY3hVdDWgKXUjCPQm6SYy2Ui
gwDi6REWxkKNRoALxLfdFRH1Om5IdoP6H5OUSxumeFjOK4b02F7StrcdLGo7D9IqIbMCYy7SOi2d
vsgaiPsVtoolp/vUROB0Z2McpSUqJxop7zEldXKDVPylcBcIURAQJbV0Sboc0ncObI2WXpnOT8AW
kuVpOL5YmK76V5qBw6bW1EuL7C+DIs9NiJLisZzbK538QfvydZTjUIu6KFvHLDR5pU8nf+Ah0qCi
bG3RjXEyx3sEJ5EgK3WFqOrUW8xd6OLikSoZSq9x+TpYSQ5DU7vDiT13wyE4CqqPOgQA1fyj5ods
HNsgyGyu9HLjzZf3oWvtZE94IbKQYYRKxlaWX3SsV5Znah0RUPwvwiqi2QtTHMNoOOPVqoriNxhv
Hga9seKXJ541L7V5ttIZXQqe+74I418ln+YCQZk6oyaiUaDs3fjpLIYosB+xNyytbVZJSKF140MV
BwhCv/cppM9ZTFWF29ghw7fzkz8fLMZKp9e5vK33imWXelG4G3keOobvfDuhdgMnDiQUVta27mWJ
u46dXvh3HqhKtsYPNVxsEzK7Og6F/s0tCboxbKNjfM4OLULgRwwoWrou9Tzvztgqtg3K6idfX0Lb
AuRfqv0dtM2Wbv3Fu2aLDufRW79hkx1ubwbCNcJIdrZlx5zKJFhKK9IYb0VuncHVfqx/6zrE7QjU
IXNfq+4W5P8qoxpMJ/7Gr5/T1P43RneH8NS+S1gV8e3uKN8wjglgFejnFeUDPku82fqCG9ms1WGE
hC+EWGeVePKXpzmBpHB35XjQTFTea3NtACVJKC/cNVfOyOeA34m91lvaSPT4zhSCl0oPWM5VPvXH
yvOpUfoDG+TBG0Bx8i4M4Mcg8Y+hUpTsrlcIc2D3ora8O/Xpy6HiXjak/mXpXA4T2yHTQ81+SKc3
izVVzsWXMBY8Kfuk7Cv1/wgfXW+ca+VEI2vFdqszc8EyFygwEdeh+B3+yCPV7XjmN1BEhLW1555i
Cg6V7Bj3E/891ydMC6Ew/f34M0LZhFffIE+fS4OCJ3uTpUPjxDbLZic46w5B/gbYEJ398ET5j2Je
8HbipbNxwI+eIYrJqezwFKDrLZI1JJHSG3JhwOpGP68cz3RfXJZrTo6CuXWAgCvXlqmrfsFmEj7M
Ss3oTHFHcrCIZZuGnCrJfuD61FzKFnvpsTsvJcXANVukKf6EtYyuMrhS8sUqY+Kp+55oddyn1jNb
yizNM+hMTRto7caG+g+zaUHx+nm4AoKitMaQYziRRgCaASofw7OJkcv5MbefoY19UvNB7iU51tjQ
ynrHqxtxq4+ZB7sKpt5Zz7tndftRsdUYjXVaPBO3rPyooQYJGccmOU3DziNLmIUGTTbnWmqc1H2/
j+fCmB7vMJKMrX1QJxpEfLDSVYyDxeLnBRIUyoqIdt54z3244c59S4gwGfdTJbO16Wr9GX5Ahg1L
qieHVQadT9avS5sG2D65Y/zDdqnLJvyGFUA2S38BuPkGNUtVXEajcN/TuPoBOBmnf40IYTk8P1sm
NDTrZsh86MEac9VQBiggSxUCCyHUDjzcuzXlZPB8ZyxvcKOugfHzq+ei6yOgsbcgoVmXRZJ2uJDD
JR0n8iJ+Yxwim0mgKsaBlMaJHLu7aBUqvRDci/8eC4Flv5ENcxURM3cQpfU2JVyPiW1IV28zcS0v
9Xpc/8xUSembdcPcy6cAPjJj9cINn4GVMtS4ZL1FJyc+rjaEDrNoimQ2zA1tFtdO+FSaoTUH5tkj
zbfxEjYBTzL1kilQsLGnzDjrexqUEWhHLPvQElsqM5EbxoCcgV0mBKgUIixCbxURnKYQk+OLhr+r
Y9hMXSkjSn1afv4RGO+UR7FsTFwOHXYx6LSd3vNCWrhNmrn8ui17xHDICKcyCw+1+Rkfztn1Ld82
rrZIBSETw8Kt1hboD/eDKYvlJ9tI9ANockqNewMTBCrBXZQSatjEFyF0WFtYTG7U1FnAmPsfeMKJ
K8vSLHMX0iFGh6VcpMHAwA0NyE7wnz87hO+qzTTbY3epH2CjcKi8So9RzjvXoImhnXIlQelqXnsY
2rE/Y6Hm0o7vg52VdCH4EmCmvE0XU4aaPOiq8DOniLPhqyjbLiobVr2VrqTIm2oYNc43b4T8AJp3
ms2CGPPvQk8/Xf2wFLtzrk0RMuHzwV6hrtLF1S/EtRiX7btcCXuuuKHeFbeTvQ9pGNgDiF6DYcA4
x/j+Cb6NTbhVPNIOfnfNW2iky/SvlV/ehAuqQv1/32JXXiFDnZYMWp2eKGGCtu3cfaXRI7+j5WYZ
HuPKYrVkmGCrLVxRqhRNaBZCnFuGOmklCYHCVEtKiMtXUZHTdH8A0C3VFgsBCS3E7Q3Y3m++Lf8o
WpXmOjyvJ+px4mAhlmU1661NxR/9dFgqdky+gXc112/sXGvQ3P2gSBi3kQZcptfn7xh+gjd1kdyi
A3HZ9/UER7XN42uRhpKTTYwn46N7wTgvuPGPbnD7aGSV56+bwqsXom/zF5STd8TrsVoOn/HDCPMX
wy04z/FI3lPPDSj63DeNAjWIMkFA/RJC01CTMXN+6c19DbrkD7YiN0gtdJvy5tfyOIK1CEQsM45l
rXu0T8xJgYXmid7I1mOjKEnFLPjIi+h3ZvzojuvtoU4VofncQyPxAB7NOIjxtv/M5wWK2aP8fXCm
2blg1Iyhkhu7In7od3NDdT1/EvpmmJ3QV6+i2/plNlCENtpDKPPxNxwd1P36lHbINK6is7WTg0JJ
kzelG+qaDx41AipLviAU7+kx0eAAimqtx2ABAKVy8K53sHUXBHdvuBOxCeL5gIyxR28G360IYwaz
FHEUixiGj/SPkXTH43BAESzV8/EPi9TCmD+vGBR9DMaRA3SBp/RXg8Oy3gO84OxuujWyrWyGxvIP
MKfLJ4UdbCktfk+u6jyFdjyEEl1QmF9zSpawoQf0DQTDajvcVYCns0RXApnVQHSoWcvC0PiyX7dF
v7r6NiZrQkkfmecv11saH6c53RwUvHmFBwA1+qmn3bJhc6VuIzezRFVegLrRNPnBbT+3UmE+HSjl
HMkxmoakanE9FL78YdqNWkf6TcLnAYkWc/CW6YCbATSJwuAeY+sfdip7encWpM1kGlpaVkF/pFYz
sFRoozw1eFJgOPGB/hKhI+GU72AwC+q5f44S5AUYjrxNVVQwGXNlDiBugCM1sd1QL5aW4W0pNmOy
vsObgDW0AhMgo0u9SPwOXXguLjp+Wkr1BSaCsscvEgA2UcCO1xCxnBe3TNHm735XwQtw8rYtHMBW
Ax7LhPPEs5hWfMUGLvG076N72Y/2QZQGipAWdHtD8Kh7tvmGN/ayFTAHHf4sqRZ5ZNln0gnjdKYp
f6rZdP49wmnu8mKBEfWXJ1JRC0HifMDwrBkuKsT6MCODxqnts6iRQwFuD5xWWJcbCbDU6e4eIiTi
k5YXgbg+Qq1V9zQQ60mSMTYXyR58A0/vg0iXA5talz/dUhVPR6Gj3o1DHHWV0cTRHn0UciZBSGKp
1PIWx/iXPmmd4ngHn7jvQ/yr5m6RlmfwUjsYalRwtgJ0BPwS5HWusfxnIwm4B93/IZrMln+9MdEt
vTu92RgUD2RCZa01qjmi8rtRGIobeEsd1so0R/4894ZU2DUcQ/rhJrgLv4tvJo9s1d2eTejbIose
LVjVemIeWvn7NzR9KWw+uRDFqDRVlhaPRlr5C4phiORFLFhpda+qHAhBv8SbdBNR0KP/8gT7025i
NPM/lWVg+X3NWkISNXuIgsZCKkLK/XQ2AB+mV+z9JRasNOkeqMNECBpXhV1JS3j7uD/WaJyh2b0R
kN0NaB5M9hmWVEH/jeyptbpsRjkWYKaHsrP6py/092hxfePTFfHFAFf0RVKQlgfDUURptQkYz+FN
QUy1QGbJemuKIRRdzBAOoNFZ9eLqAaWM27xqRPEGr/CMjEJrodcjATwIinrSjlcUBqAVB3I83tyR
mjK8hocxec6JKPPFJdwpamPfnXT7YeE62mcUdYHKNLeVXEdpwNuZ8PIlgka5hrjeMbtSLEV8Lz6B
XwQOrh8FAGUcHMx23K+FxWKTso3MSia8+dTY6+GwyZg3VsjGuiROI/4/gGkDGDKhQhnHoNe7BTq2
kRAjrFAvvcqak9w0ZICRVjUtQz+rMOmthj4D3SacWnUyL4vv0SEAXCCJlS9BEny6bwGpZqQ/+sXw
P50ue/p2xI+xQpiYdzwMfedLle9iM4W42YED2Nk8uf6lZ4m+bA4/3DYKi7gDyCPiJ46DgW5RBzjU
0g6zllyKiyWabK7RJk/C4VVCad11lGIf8r6EhmFUXRM33833XVVi2e9TY/7LIpHMLCxZyInSBiYL
yG6czevfEUCsAq0D8atJksvOF8CB7ypirFseuD3/h6Vac8QglJd0Ye3y/McxahP/EYwtBUS0wAbq
uyOLrp5VHny7qHrzO8CKqzYsfAY0op1/6BKgDheBg6mYF5NzeNOuw2yBJ8bQdJy9rNv9X/3sWE0A
TL+BMb6+PylLXIh2O0xuVRTYhb+DJUoMO6HK61swsYGGryK6dBVe67tQZsd1Je3qZdX+EZpPpxCz
tXBGxUjiwFM4CCbrtXorMLMzIA7R6BmBB/NyPk9vDdxPuqW3twygByNpZXqkEfhE2G4AwGMzyWTQ
q/epz0epUlq2423v7f2QZe7DaZZXzlCaCvYpkUW/J1UCz0DKAdlqrMqtoJNsJD42rwP0YiJ9Ka0A
DJj+P03l0SD6ms7LfYgNIYGZO5NsqLch69r4lDDGv3rzNuhsH/I+/aHYEgLrbJ9IV7QTZ8H++wAg
2+a4k/0nQz0palcE4kpLVXbC3109kq1B/f/9t0p0cVEPoLHOQY3n5jKt7YLNFjxBi2zIRvWmo1dy
mbUnSzILjBr7ywimdEmBR6YlxvLsgUEKXC8nn5W/dQicVrrNfA4VOGO7b1gKeg69WA7mELgBrkul
Nu9b502uFmvuqJzo2Bwj6//kFaYYAV22/Z9uzFFWGPA7qByHndlsjxQoKAzpESZflC0950q5Lu0p
QCYRhSfePvpGpagX++KYobVWQXf2R3G27JBMSdeeqXRYCtJshSXX93t+7lc5Pj57hs5G+h6V8lvC
Xgi4Mas1tozJMMP2l0KtlogIaquhyO8PvJ5ttnyfpEmAjH3tgn/h4BlIlR1BzgZYkZReZyVF0FSm
M+gXEH6V6ZENcShOPhaWV7NL/6E1fulU2kIWbjVk3x0F67Ll20UPgCX87N33C2M8FbMTME+rOpuK
JWOYfNaAzWOwTm8mbcp+9HapUg0KqleJrBo8MuF4sW27VEFA91udt+fICFEHiKd9wr2kWQsmy53H
nrRwADvEwXbZqGtrP7UDqCEkpZ6kd+KWdz2O24lCecI4R8U5A5bfezolRYFY7mMxclBsgSvgm5cM
OP+VNbc3DRJ2k3kqpmwVZ88np+ydA7Ac0LwCBiOBwXNJUXlMojJiJ1oib54JZY9Iwv3/3lA5UAmR
8aaDgf21FbquYw8G0aAkO+XFX95QSXYcu8OuA+2kZtwkMbPLWvnIulIKPJsphYXQ5AxKbTrhMQye
nyy/S3zQPI4yy28GQ5UAzdIn3Ey5FYFAON+SVCfxcpuSE/nylNASRChMvqE9aI7BR7gA/ZcfvwaL
nf8S8LS5z4nBK5BflGfW5OTFDUBHjSmvuDL9gsnBGFxVV5UnoFlJtLEr2VUz3Ov1Dhoe1CK+3V7+
NfQmh+eQeW6SUX62k0uNuIjj/fE+hHeFNAMyga8RVA5SQaH8yjOeU4Qx+IRBN4gJwZ3L5GVXjMlR
gUtTCuIwdtxNO9PoCctiv+GahLwNG94KHr5VMKh2l7ye/bLY0Trc3vZwH/KfqbKU+d0GHScZpspL
F6jYaZgAWc1l2T56w8v2yKh6pYF2w4uxFJaPV9lXa2bZM8BjMZLK9BR/JZ9o/CcqtzwvHcp/WQQ9
dHj72thC//aoVf4XYFR+KkOKqPYqB8PIwR6l93IDAI6mPnET+RSencJmlX45Mg7exY4IaBLtM4MV
tb7bL7xBnI7jA6ISsR3Dmjy+jEAtLfd4/GBC6f1zCu31QQqOKJicRfoMgoWCM+SgF/uaImZ63E6+
lDWWRZoEAu4DzxNhv26wmAKoWJgtB8l8PSXXgz9w+MLG7hDpogkPFJnqQaY9RHPloSQVsUZLwChn
GPMXAEosk6+uBRljl8+siw/Y/giu36tatzaJSc/mrWq/3nSlpXo4l1G9/A8q+d/H6OX4xba3vADN
q53UznwowqYcFaVRnoqDB6oa8pirdjXy42hgHZsNobXyccv+QLxYgSUzJYOaU1PaUyYMkGW1SNE7
O31QFz0Q/w10mhtgA0eZXg5G+UC5bD4aernZCsaswG4DJ0sKCM75q5P9b5mPmw+a9WbewDSO5TT0
D7FDYtaS+McyCJ3jcYnknhqjUL4wzQLzpOvvvQtxokUGbOJKd2m7OgVgRSh6JRhp8XpM6kV/DVJ3
RHtBSM6ZssJ59XpJvr/zg662VYU+A6coiQoOnKk3zwBI8DbHpUlTfHsBxZ1Stgj6EotnJQ+eydaY
KQwAhYESWFsUDuA1ZOQhyaxe5kUqix5qiFHEDs9sewaEYwsEra9XRQhOk+PgN6RTMc+pnQJUPI0I
AW+uNQMiOj7TE/unc5GNsOSeQSTImzt+TKbLcP3qfnCUxy1OTJqzXa6guqfSMQkwIawXR2Uc5E3V
xPYTaBebXJ1fCJMJqV78LCE+yW0bcoo73dXS+TD7X9GudA0UqITQeWUZP03Mjstw1tbsOK8sLGzg
gDPueqNBWDvA1Fmww6IgVWYGdcMtH1Vzp2x44l2FXeQTJ2Ueyh3BuDNbYTzGuC2/GZuaSRkgmY0F
ABcvP0az83FCNrcIfZ0zNxYvs1u9kAghXnGYTjTBavwdNoVxkV6LNF9qconQh5WtugSzfvypiK1j
g8QQxuIbd5W9GBBw0M4YpqLwET/50fEVaSsDCJ9mASD1aaG/jiljrprTJfFgRRG+MdL35BH3ZuJ8
0uKZtyr+NVrHmBFvl6rzvix1Ijkx3i79b5+YuqmADBOjKtJ6rhOKwct0l6iicTcRQ9Ghk+7SA2Wi
R/oSSkswN+dxScKF5M3+YiPdd4lX0BaKkMtEDMDdmyWC5b6u4qnc3eOwHRfIIynACRnCB87C4lq5
YuqGqqIRNIW9h56dunmKuVNTmfYcIkDH+U9AXCYX3bpgeQJorrhHhCIlNjFOdMvRPSF+ur7r+pTu
yk0B1UrMaGxHnfpQUfH64jtvCyy+EGEG9ORJ5p3NeEPpz95pLvtFtjjGzT8ZayIaELtdO3TB9yke
ltbB8QDlZMlGAmAMr6M5F3RoxXaZzLut7uws9uuoXYofgaWZU973iKf2myyYV/cvt5yDKvEoKRvs
poYTr5yx1av1PDspBHMuYpRmEhIzJVmeV8JdskIfvL5SsluB977BqCsV1OH3zIb9Mf03UZG63k6x
1bZVMrissbC+RNWRKbSetX77XIjzuDy0x8g1az4mk3/4XZylbMw0GCzp1CGlLk2MY6CsHnttJGoE
W1wf1Sc3hl+kEtVWeM5NPUAlXwtncJC4dpVuLy5y5XXP5K2+36SlxOWcADBfX9bio4Ta6Ys8cbw7
hJaOhIp/EtG9fBwBr9wkM92jrLxRtaZ40gWkhaBOviVGOlzURbXkPUdnYUE1Fih3hruAFmtimMVv
eJenSxf5OWC0m7Q+JTxkkV1rU9XBjii7NDk/taTwizZGR3/asbQN9T8A1syGmK7J43gTj5pUNvOj
/0B0iepKcOQwFL48uRUmccGmDORECc7Aj5ZHxfpqjp7M8ioHQpXB5MIuISrKe40V8l2ghDN3i60O
oCeTWavee7VzpkZ6s8Cire5yeg8x33Bjz0QhtDEO6U6SIlfhCDBooPyzwDJ2avyj74fc0z+AUvRI
9tnAMAZUdOp8hZcGREtxHiOC9qZ6xaXbKTV+t36oQT7xe+LcHn0vIRjoiwJERI8mlCfT8w6enoyR
kUiqqfreVwge6aOdOK6XaIGpHd21Tyqr5/MaUymARBckW0lvRoXf8KU6IKcAOZX4uEjL1W2Mjs5C
KdWwm2HoTfN7WEXp7G0oBuE+KNfetQdq8DMq7MHiGYX6rEvk8qT/GInU3a0IYwCkjEQfmVytyy3S
d6OhzSiFh1db+/43xMpJiYyuC9ZBEkH85Nlf84lOhYHYy27UqTA5gbpJcLuHSFMWIvKkalbYJgUS
6S77r51Iy74lOHiCPgjn7gPjAHD+qLNcqEDMlb/sK0QalUg7shaErWSU/AtzC49+u8Q7F9cPnkFd
yC7hRY8YnEjr5tzDCqeimQAjyG83j8khoAtd5uDAXUIG+k8YHSHRLdk506rPZaAMkJ3Lq7ztw5rb
zQNGgpUxjixZsIb1jNk/33BMi01kH1psiNsCLlcHSt78Z/9VwNMYrEp7SeYFGr4KqKXf+lQld4td
jqBhZ7/Q9tPuyxYmeMDcM/VMZMB/v19Nuoa/t1FHxfnOla1S5kZmkTArkAmgOUJOwEZuiEyvISOq
sGUnztwg1xkFQgkxazM4kqJKoIfwo8IrI/1NHfaaBe9d7zQ1wOpja9+F9PGlU66WYsCg+8KI5SCO
LAk5ZXj5tH6i8oCy3JnjJagiUVHuMfw70IaWUi6FaPZ19JIyoAePAwK8EWdtHIf/ips0+qOyx/vF
AUuKSwgPUPt4KwMh+YxS2LbQR+wMd8lNP7hhKKvnI7JCSZ42aKcOSwIYKiJSc/PBU62Dd4NbEIvc
VgPymhYo7+g+Eqc6skiLw3H/JUukSOcBsUm1LW9xHv8JIGBUL+j72BL7glxevtWAh1OrYI98NOG7
iUDXy1LtEd8/2HojO0AC9rDh7qDTRwZlq8D5UDfefewpwZyy7eqBjA3ncPYkf2oMdMaUw5ew1Xlk
G29x+O+AWSQkecaDGExRBjwdriQa28He5FHuAXH9QZTLKOtJE8co+v6BRgpF31KPufYcs0dgHDy9
I7mGZw9OvfTm6w7P0dBQVE7ykHqGXF1ZSX+hP7R8dqsjCqDtCclPXieZWJYcz/iBZLa3oIfqGAWB
MJgPc9qQdA4Do8uM5A5QeE6uphhO+bHSqsd/ibXEyH41NAiYfn5gVBP3VrkQQc0WLDvqXC2E7qyh
USKY5WuY22GY/p+Kn/v1nmOeGftpynnCHux2p864lqSTjteMRBADX3dEFZ7/lGbgof2yoLyNrygT
JK+iIonAqAihekW3kOhJZ8n+WgHXdb/GjEoe99wW610j+UrbYHuvupxSguN7+e03yw8otiBBpdj7
LzQHgA+wjKro7b+TjqQOtMxSUOVN/zRmlsMr5tx24H3a5xw8jC0k5Z+6Z1TuYpwGvnYClcVNetZ7
NzBAYcsMJGZ/7ZcYP5ABwh2eX3JBpVIM4GQlFHFZWpzJxcTlhA6EgXb04PoFM+/rVRBuYb4idF/S
RvEqvhncMU90q1Ebyg2gS6uqp1I+H/khp/Ltz4KOH5iyFk66dW77IatlYpoNMf3m7P6lA5sYOvAn
wMxMVnxVT+E/cpaB8yzBJLsa+MbAuJ4rH9F42BddAFp+uVzLF3oj79UhXTFFHaIN0dBn9XZdhhPl
LYpIvqGwkerosJPr5+Xbqdl8C3n5L21Fry+9vIpDhGke4fAULmlwrJ3OeMDgMizqW6DZljQR7B8W
51WhgPMqp7rmgmtBY7Hpse5n6/sVFJ20RfMyE1P80pnZr2xGUzDeNsyGEdC1EX2RgFGvTLBKhm+y
g1V6my+llQhSxTi2HrIxyazsp+NiAulgmd3q7OwOh9Sl4dpeVpgzHxo/ucSoD7GzmlMQJHkD3sUU
BL7lseCtkBD30/bF0RJB3ywoMcPVW2YUm3KDyP72UWy3u4VaugJn2AnbRMJ5VdWDMeEet+/U2qdd
yJeeDxURLfgfmtkh6bNSFJCe321k+nHVjNzF404Pv3r0fVDvuyibK9gvexHVxVtGFfs7NimOGVfo
6uZlmDF8hnOP4xyfcQ2pjkjFNRwhAFvKIahhvokc/b3CDDlMFI3p6oQYPVbWX1HvNmfliI0MQtpm
jSet+TaxZgbaPiEsCBJj8YFmPEhe4SiQ5oLGib7hO221RB8Ykil5ifiaZegBtjaNMcBsO7uQEAo6
Jvmg3gMkyG0f5F1z2q1poh6CSjE5C6WMvpgJ6kaC9qVCPneTrjWoZiLbNLvgJiuqzVCStkpvrXog
S4iMiXsR5kTmZpfrNtZ7lo8noPQF8U00PBHSK/Xvn99YH6mjjflDmfb4VKsHGAj9bcSLXomxHTf6
bJmV1zn5Y10phM6jHBnr8gZ1ma4PnzG3Z8u4fqHbMQXaZlsbPEa/qy5JOuAr+QIW2ZCIZ8Scrs3q
i8QpYNqAY71zt2ZCK0cwx72XgaBxj1wxp6V8Ni41Q7oI/PlkNLlo5RdC4rEpCo3wgU7vKR10LP23
NiA9MwO7ldsShUyPtninzsE+eeViHXxJPD527FrYDtgb+ywxD0E+eq7B/cW2/EQ8Bb4Lzk7fAv68
HAvSoixj4aotrC8KBgBZFJcksZgfQSEaIA/PyRp+XvNXlAxT9JmECA1BapTV6rFRedWbXvTE93Kz
O2hYUsYMYjsIoFEl/rZV2qy8oL8Lyt1tjMFfVTp07axzzdaC5omRScmaQxyn3FoFH53q8iCF3UFf
N/snQuWtewtKJ25wnuEchWq6uQrNbt7Q5VitnsIgHDmzSlN9tBnXR5U/ck8u5UpiG0F4TxyJt0Kd
U3wEvR6uqRMdScRdYx38i6MEOIhxhzOw7x4ey/L6e6SBeLh6bBz5NINsnAMTBldxs7eqs4+zHTv1
uvZ51NHHHaMqaEtk1lc3JL+8zg+7Ha8EC3Dpk5A/zevuazO0RL1rmExyseeF2L4i4bKd+Z9UlMvu
63o50NUR2O122Xa4QifanGfsJeGV30fPYZh4S2qQlM5JYoarjroEOtUrjUMjXbTB6VbN2j3/wAfv
ZcEKzEAmI68lY2yqh8xZD00m2vwDP1Ud0zX8H07syo1aT//PgbsffWKB6Pzjs5AnNeU7kh+xFAMo
kOliEaQYMTmUKWF5yW0H8g2AvcAO7sodJah8xiU29cRTEV6y3gbPXFnKjtudSbVODKZxfFppI6xx
XEOy+09alf5w+i3foXfJTZRq/3fuhXdwAjWphcrp2PC69G/1rZGcr/T9M0Mzx9atgv11yHOzs/K2
T82dQTvxQRSMO4nE5vutGTezSIe1+bbvf8xNK0lvEax+QJRNxtkZ2cdmvEdEpiqnzqalcve5vEuM
NGJb7JhMKJcpZ+3EwRkuFR3m9R1G6ZBzaru0KtgIeHFK4vt2fKGUN9aeD6jgMFKWhCa7eET+k3tz
+awy5Mz9EDfeiwa4tM+A+DuEcipHZh6hGg4rrW1cdoW8YVJ+5pnDliAg+xpnUlSS0C6mlMN7/d2t
kdau2lZeFI7/3IYodkJL2Hamv+VFD/6GOEwfddF6/IF/D7Tsh8AM6hIi3sPhM6Nl9ejKM+WfDgjC
kMdEfGeEOnq9EQX9HxE4G6nUOKqglOC3lBnIZiKG+gzrbPKz89Ai/PfWk5PeBf80zMItXkXIn5U9
9bbxHlgwOlscpcFsw9SrypydTCVXWqXaC6Tg4kLFHFRl7uyeyCXUxw7jmAT4chB48U8K20sCHjIL
aAaWnC7OJGwgcdjNJdMcVpSPGzCAjllmfR5EC0k58bTwawbxgHWmP9/0TO+qRE/mRPtWMJGTJ1wm
gXCkEKgNMns4jenPDpWRHh/ofe+Z99/x2IYmng/eK7VgzlOxvLy9iZnZKN6Uis4l85dOvkYIbDja
Ox1DrX2t6erPIyiWP1Fs4Gt6dQJRWE87F9xFO+TsVFwKt1Jl9kOYW7zG/R0ifvXx878nLcsC2cS/
Zf4qcM5C73QdkXKxoJEJ7TjITgEmiHKXpZKHt/cmoEwYrKMFkp/UtLHWEqhrjmQJKbd5lGACxiIw
oCFcETYXQZljIotS713g2Vn2kRD2LDrdJ9pLl0CE93QE/AS6GJxnYvOTgnc/bExDwSHkufRDpWHJ
r3zBA5ODb3pKlYEnQWtqhFaG06vtwX9NAmMIGUVvXrBvElmsLXqMGQWi5WtrDcK+X9uQYYsqiMTq
6LtDPiMUEAnl4IsY60MDVH0qwpMaFs2s0FAXoOlx7v7wykEiAtmh4eq1HhYsG3O510VF0ugasOsh
2WoGTAKo9NL2ZPWnceYwmgdapN7xPJ8K4Sr2jO1pR/y3G/vghb5pXPIA8EA8Q7sMlHRCz8E9dcea
VwR5pKBiizNYibbhskO/QQf5Lh/peGe0P66WVsdoXc/4s48wr9v4kuf9tP7FP2voX7Az1instPd8
y4nB29G1qL+vQFmfAjo6PQtmXN2VsEv7CsoLNdoQ9DaHR46K2LLaC1l7vBDHneiwVomZz14bsOML
DCKn/OTrwkPj0lYiIvWPBhntLvXN3XV1roerJ5AX77Qq7PknJoga3RvfijCQjAoR0rGfmjNdHf5x
wBuHY4McIYxq6A+KBY8boMLGnPWILt3mudlmGd/B2VMr4f5OHZS/3TPOYYh4yv1r/EcHQDgvPR6U
TpP4g4AWEfHK7p1IYgIQ6O3cjdKdh5QuY7VZ9HCaeIW5LJLqjYEIhiOPqFuRXioFpt2eua5/xPI1
g+1OSgAcrHfdf8v2I+Tcic7mSiHqgozxlm/pW5xzZar0kVuWT30jquBhOJq/vuILb1AVw0uXPeUz
81Vs5b2Ac2pZ8aOCTF7wFDSxVYonPkImECWWpCHuLcC9LJfOkefsrwe150JecysLjU745YkJJbai
ltNbr82W23/V2j/OecVZaRcDqiaDrDfW3ZN8KSAnP+oq6MkeeoulA6dDih7QQfcA8F+QEvUqMC1R
B5u+Jntigskzsr059xnEYE1k13w1jZDsnc58pf3sbYuDMa2J+TZCxd2Uh8fjbwiLpurcO5CyOI+K
DmpqXvN5jlIH8TbzvqXiIE/m1aZqmbh6Wqwe4Jy1F5pwooMivVyRxVopVRdgc8N1uNThFkvE59WI
DrBbD+rg8QCYY6yicL+yvpg8YIKL5SQR5lVE1HEUXSrjowkFkESqVEmoygAATrn++9YrOf61Iqed
iyKrG74cDSyVq6AcEFqLB/v52NnxUAGq3JU0o9krIGbKDXI7GYeTn19dOkaU3PWI2RQTuDKb5YIl
YQf6uL16ZYWkhwWIABkz4AYfPVfknKeUSHsMzeV6cwkTCjQFMiQ3Qv1Fzj1L2qNRV+79I20ZRIR8
hJW28gmE1Mlkh2xScx701B1HFbZ9wTGYqpf2xGS1dAP7kdZwTf5DPjdmZP9JLB0yhlEzGuSYd8BV
060LssaJXTFQr5kFREbAc28E1AaXO6iGC0eJSrbsrZCCnSc0BU6PWu/6UdQ8lIgeoPSik3Htfet5
1P0hURBq5O+H/BHK22RLYnjT2pAeDNmTl8Sb+CxJ1HmLSajAALmEhCVcqKESg/t6WOPHLNp93YMr
RwM0MKI3kag0KDkxurSRnNl66FC4+7aTY5qh9mxSr1n8Ai7uPezUT6kd6nOQHzix1ilVc00E6mMb
ETzOpq2TFPI6wUtEITfvS1hyLre2H+6BPBwCh2YuzTRy06g8nxUqFbf9wVfC/bhrRBG2x+arasVo
W6VQ2Giuym2J3o6JcLI8n/+VoPSPKfSMvFvsOFZNyMboA48mnXMmtR0+ddCQILq0Mug7Ktl4tM6x
mpKGXDC419FMvGP4SsxRFeQfqGK7HAN0iyumrchl1HqZixn6idZ9SzSAkr5D8ZVaq57CqlbtDjb7
R7uepgH0fCkDHS8Tdpn2G3XJHrPTmsBo6apIoftgb2/nWEqivmWNWYWT2fwCRhDPuN6MlluQE5Xq
m68pmCKJR7gbXD3utdBqPjyVQwFH9NYfMla4pNdz9dRiqg6FJwswsdYO5ggDNt82487vS3IMwl+a
GtGX4PnKuGt26hHnHKSKGwIbMKKGTa2iHDHO2xYJKS4SbC14zZOB1IVm7s9BGiUJizdY3t4PUg3x
4FrVtfjvi8kNbgq1/8U3m9sh4bkPeK27Tr9VpSSWnALQR4rmfulMptEYYE0/ejuQCUW986gBZlDn
XfeYztV0E5Dfn3jyY+ppyExGpTYsmgeL0WO32LkB3VJZVL38PppavvJ3ad2FYlS/4ovhvWeK1V1c
m4XU7gcTkUPIgl4EYDYiObQd8wYQFl7QrSHq447sclNWpdrrgE3EbS287bsZgtFbr2Q0u8KuorJh
2D13haoMHKvQClWWOCxwa7mGI/7nDWBKvNEiKUo2cD36NX6LjPYcEeN94P5pFuccyYan6YREqDdG
NXH0VNI8Q8Utx4KZ25fTes2uh3tYFzcjTygcVrQLI3I81DDffWg7qIYGEgINHL+UNrF9jYWJ6Uwj
MeVOC0rFVlWINR82o94Qrg/ygLmXx7I+xoWO5GxWhRP2oZs1BNFhdgVM/fv0bHJddg7rIeupr2/9
NCVwzgiLKjGCTvh8tDJhgUDIQWZToMM0VpQ2vgeMPV+Dvdv3PE1+XKaBZUh8wB75/Qlf9qA+xLur
9fS12KytI/XpA6PszdNfz/p9zsL3/x3mCpWkLy7GsR3eTnip0SmOll8vvfG0rEvJpT4u/+UiGuU9
en+y3cBiZAovG0y5DzOAMAqyKgvduzzQE5eSiesfm4uibC5ojhFmZ1jsZKBFi6hrl18hechWRgXI
QQoUmcPtpEVcc6NkMShV5x4uC4AMw8c8mY8KHNfjD3n98aIehPRVf1058fOls001AmyIDI3ARxdx
IE/bYRf46fu1v+ODtWJU/diY3tWk1dPA/d5403E6jboJGgqNey+BZYDsHZmCc2ZNRyg3KLB0Dt+r
RVh0dJJMY12CDhqq9RIxMSM1Ql6c0uaIxUy41vOvuRuZUdngoMzehQaQxjRJ/iut3bg25akkY9HQ
WYyx2O2pP5iO2oevkBJw8maNpy5mo1JZ9+yo0xMCHmv74J28LEdaIOoy+x5VQ44q1nhLzoCa+n1k
JI0SAfh/RboGUbO0+lxnFXSa4sWNAkZznmzbF9OO14sYLuJZEHWEVbse6bMbn+Ivp/DQK5+F5wVU
SSGBTgcEqSDgdFRM/n9ZlFenw4iQZh02USmWdBXUvHIlPZrnXKAJHUetOfuYaDbzFCUZLtTK+dQg
khVJWWsTv0hQDz22Fn2yMd89bFKQExvSK0ZZ/ENnO5o2ZcxA2azvbNz0lhRXwJA/eU2Nm+EXs/Ab
qrFzPyKovLT01SJwTtdsXeTDX3/Wj36lXJV9HTuqaOWaEHFm6CQ2MX0adtgSnv6dJF1QFdsRGNRe
rHsDl2EfrlvTI82ZHRKoUpWdsVuMwiRN8JjDchxRVhRM5VfB1VIb20qq7vKk5d81XfdSJ9oKPo2y
xhZgq9VKjShT3EmWTx6ODWJpOO/ELgGXVE2bI+y6uPU0USB5sll2j16dv8SxdYmisfIyG+BpIqXt
cW54bhE+2eeQnjYNXy3lgNKiakhVAR1EYntLfDImgSRFiYF6BUwT26i6jRcrpWxep1FY1bnMJjte
4jMWteOmSaeRqwDAMkOt9VdyI4eJHYDnVcOpR+h8tHNmsgMMpZI3fNyxy1sIIqokvspEsCXt3Luw
TvyymBSIve4h8Xq3B2RYmeIooDt8QRA70tCPCWhMwS49ddSlEwNB4ujNqRg5KeaRlEs8wRB46S/5
3pZUPk+Yp52Pa2ne318/DOWfLwRlLoQSWGBbL9xq1kLfCXadC4kwZnwgTHiCdDTbNb+Q6qXVGsfw
mNLX+dByJWtC2WCaYg8tSizZbN2zJlAklJDDgNY8ilB51JhLVptdXAlKlSq0nrl6os7gVe29CF4r
7Vbs8QQi8Zc61QW0z+GLiCfEbPkdtbUbvidYC5CKbxSRRhLsGhQ3qRrU0OjJ2CJfMN/vRUFlePad
CKMTn4oKBrEtg+JvgXDapNN83hwH6Ny1S5jmcPVMB/VsvB8IjikCNyYVVycS/SkNGhEbhbDAaRxr
1AW3C/+Lhmg7GQ8kIFZyHqUEvlrQqKn0aXLGmmOMjGP0mUT0K3cDcxvShIK+u+5vKzc3QeVh4DnN
7gZvXfHYMnJ4rSjZCpBwcdsDbG0aMm1z/6ews2CkMyrYtPtKLWENqvgusAWJtSysKGst0swW8VWF
TBfLln8ytXeXWDRoNzWw7pQhqTpzJDcWPpyb1ehw/XsN5r5vkvoNvrdHAZvMosuHBfokAL+l2IU+
YJXvWOIgbNwiRYDXVWvkjfgGHSu3tOZ/urAJ/UfWlQz6Y5j9K8/SJTtmNX/otPEcciBoj7wg/n3+
dRR12aupw0u9ieEzUfufYLdicsJaQPPttHp6tE3z5lbCvDIJJn1MDTdSBgMGewPXHAktBwHkd+Ub
sp+GAL/K5uAWZrJh1mjd5JBLVJA0znaikWoC9wNxljXkmd69IIX4CRj5Ckvgo1hqR2e9+G1Cox01
J+vAiFCJd0z+k08zkqMtYSas1hme3IuXhRp2AaMqBTdObn3t05BW+21yVMnTdw5xNQ3ylZapPiB4
W/XBw/I7OE3dsNfLhpK/kp18FLIEd/eantkKkjwjQk4WGyqJsVwCuAgyBYpBP7+FhbXIbm+Gkbxn
4KZixI2NcZdZ+72hmmS1BV8nq/83Yd7yc2mlJYNjVcDV0L+vBu1A9dlwSPLJQBgap7TLEAAxtjzD
ZU/cO9Dki/zGslWPVhODOBEQdg/rhJ1ObOfJ30uwuTKQCs2MMYGdjO2gigv0KKa2GDli7Qnp2Rdw
YCXPTBGUr18ryhTcW3yyAcjcPWsrDNZ/QcqI21XyG3vawRyeOW9s0MM0bQmZOYr4b11rPuVDROnv
NWaJCOtNhGmJvaeWv42B3wDkywYJbiJMhhFQVjlSSboe4iv7ZtusV/j151bkqeht8v8gp+1VuUfM
3h0tCem6fRMbGrMBdWlf2zKPFJllO4pjAjBkMInH3T4udyjHSgU+pRD2O02IfDp5XQZCy0Ozv5Jr
nRCEvxRW8bgeWGr0ayUlaGNR9kdSCp8r45X2w3+pr1KJg54A1OiLN6wrNOVqF6p7NlF6gz1laWzr
DCw3DcTqaFIhr/IOR8iBAiUytf71pyofldi51Xpnvl+LsBxiFDxJ0gKQWgqgXc2E8UZdtSTHFy7H
tu1+eGZ88KKK8sr7C2IWqVyF2iuwir0jt+d5vntAU9VYSif9SOTF2nI3ELJs2SEqGwueH6C7itfc
7UBgV1QJgdggeFhpEUhvWUrvuHYr9ZTsqMNqeLN9a3qPJSfQtyxHCRVOW9UgAGbxoYlIX9ngRvpr
cX6crvR6xBn55YR6Fl9TqTgx+9ahMK/ANJEpPiHQUhFYP9UVkMJqUe3onMpJpFICbZbP1UwYF5we
WZOGSS/3+MOKT52uz4tqyAZTSF2b+qrxUuo6sh3iHQrJyw4ZP6UgrCUGyHLQ+kmGzP69OzJoC5Ym
44RZh0viNj8EwHEMGWdcAyZ/SOOjqUJLc4xzzpjDtFLtS5ADu5G0qfxBnEQN59jnKjdt4VntS9HU
GnMY+0mc3pbVAfFiRSjGMHLhkUJBlF2U8rquNREmp4reYRAhgk+dQ/vRr8scBFego80mm37VLkE9
9+KVVR0filez0Et5v567mboHkxCk6ym4Wn+xrGQxbq6r3OHI4o8C9V976931uYxpJXgBGBj5MBzt
Paxr0zteDTg4kMH6gLmAyNdctfaU39EXa9wQSCF4XU+059Tvaj7wTntI1B7hdWNhCn5C3pD54q+T
tY0IrY0io8Qv/Xv73zepBags3HZrg8h83xTrbdIA/IQn7LBpkdpheaThScd4MC+wIUIn+t4XgOhU
jo4t4bbmiE64G1bIgdB2RHtq0bwGWbJfAInAlu+HBu5Y4vqOj+I855Q9pipGmbbRrMEkDlr5AgTq
ZmvCsSvfQ349jYm5agaHZqTCz8DjEUK1O5kwNTwlU/OsJZbTcGjkhGf9HtSreoHV72WSuwBzMmeP
z8Dl17TlVgKKmcYk1UHQ5PQ4qA/Ok0BRLICstF6BhU0lzTTbgbS/xl9Yc+1a/H9yi9IH1eg3aHkl
yCNGha83OZl/GfvJDX0XJfIyynVGUTLltDjqUhWIQ70AH97RdO/JQenFUVDOJCFIUjjf9d0zz2wD
HLqi88Y5GkGNvdNGQr/1wB0mEOfnh57qORSSd0sgA9itq6uJWNxgLWyyA9F5D9D9JaBAN53SK0Bw
p5Hqj29Tc8V3u6HKRxpadgp+onrplPYZBxnVsgsQ2qDSA0NfdW6oMImGzxkr4g2uDI697MOkAkf4
j2Hk74PAtY7C27rWekqkYNJ4552OExyB+mlMu05iFQkJo/HeaCfAVNtvWF1pSQjJfroXI26WzDBE
KEc0cUsxZp1hjYVyiYIuKOIkl1iqDdKq34rYAcW0mAN+EKc/tx2KZNM1EQaay6tuWcDn6N/kkHLY
uiJE5zljbUNMaS74hhehunnVhh/9T8YsTcwRpLLv4sqdfJyT8Do/9Uf4YOUFVdaMJh3xQaWZbSwb
KIYmdkKSsSIUi+Uu5OOo9JLGohYRslNnYvG/l9SJpkWGpIz6uqrZx+MMuB4wqaRGxz9sA8Z+e3ff
F/l5dVePuJInJndYng6DV+A5IC6Pe6Kfijuhlu6RdE/a6K8//VtRra0M7K3oY+ZEF5OtN6/5LDMa
xEtvjELTCJ1cY/rH7KKkilzFkrd6QZVUMDvOcq5dQ5QAoMfTswfoaDLfH/M2jzmUMhOF3rBLxNFX
4B89kaTSZkrL6LO+iJe6CmAxCCa1eu/ABR8OCKTCnmdb2kqKeNaOvrjfyFojpw6ycuHvTYPZYNPd
SbaJhVUqGiO45/NFEcLvyiP1hBR54Ya3i8Hg3jsoTGr+nCXb04BmW4/AhkGHsVpy1BEzeY7CLnMD
iQvuS80W5VEijIvZ789MUh8jN9oQZOuv9Obud0tV2dI+AFzHBD4kR8sfC4Di5Op8nnYGtemwSJNa
1eoo+SFrrRWOLE1rJFi9ikFyQc6fuU/EdrUJCu/qlQRHMl2FNjYkraeexTCAgz3u/kdyHRjWcfx8
ROqPRC0Kp4mANZqWDi9i2lyQLKEKy0CN0l+WbPfcco3JOGkRSdNzKsM2F/trfV7Dv6xI5UAxpTbz
m3EqMcuMfi35HrLpm0JZQiFI79z07m8/1t/Gzkq3cV5qyM9thlJx0LSuN3b9SNkCsc4TgJc5YF0h
+8mzB5X0RvWdiMg5mQyJzKiDyV3VSCR0hF0oFBykJV2K+9xNP3wlCfgP/mR+QD7jAVSBn5VRD9t4
rbKXZaLPOaQ55z8Jm9WooW5XlNVDwV29VNOChXuj4kQ0EqvTMvwcaGvunrJCiyZLCsCYXwH7r8he
bnP9+u1AyRy8jaGGG+oIp5yqKAYMz3EBOcOHDUojZTPpnZNPnr7wbqWlTk8hXU6TwusfJdfYdeRi
0gmM8uq7jrluKb0F40U2UHID5VTTI63UQ8J43Lkp7CXFpg//l4T/3yepXFWTJngAfGCa3SJXhk9o
VNTxFWA99NN4feYiPltfK/axGk4HZYHHODF7VYllbKs4rUK0yHvqgmcyVI9j1csjVAxY7HbzKm71
IzLbzb4cpxnMk+L8KHB9i4YWyXcob+ysv1IqqaTV26iw08EnIIQetC/dB3gOLE/ytQfQJxXEjiHF
k0JCi4hspPH1+8a2BpuBF52/xYVqrh6nHV4Ug64G8QUGBUS99dSSonqpmyRYE7S73wDK2mS6fhEW
5lXj179VaUA42sRQM8cE1FK1fv3QAelQFFDdblL6uZ2UV6X6IW/7SaDxvPnacJa5t4emqGvdNSb+
314jE3S9gHTyEsvW15dmOsri/yCuwV0DN6XiCjuRxUIEs7DgDYvm94h0wAljTDSuujHVZ2zY3dm4
rWtu4hrUxY/0QhAgtWLzSx7GjiE6weU5/Ewz8ngQ6axY5WiOqkjFP4D9ILMFVYaNExCogJ8bjj7D
DTrYdwGEf41b0pRRRF66p/+Ur2iib/K7lygRmJ9qhphcGUDqzYhOPvFeKND+nbzZsxiBD3m3uzAL
tNm3BiC/csh67JknAzvls/Loyj1ohpuCi4+akLctKTdoqFslbBwf8E1bEY747uc5EZpJDIBcIgAZ
CNI4Pivzh2DV/RcSrbP+NZpBHqVPqM2FCycQr7Em7dx5SvWMI58VRxLMeEeK3guRGQ669qs/s29Q
AF/mFO+iVT7OJ1wCplLEl2Sx/R19AIRLetQE3Tujx3yvMjzOZJ5xMx3iatOOWXZgT1p0HlaRnIn/
HRA6nbto59jrkVjO/iXTfYwZr4fXpZ4SEj17CQXUIbypP1glS1lFhBM8kTwmlc5QWRABXS5uH6e0
B55opgz26CXOSuXLdlGPmDcNmmlhbrWgW14+L5EeHz1skD9dloq0eA9SrLG3ueSMq/lZATsMqy9E
DenQxls+BH7a4BmbVCfRdVP4dgBhqzB9q9GuZLEOQo0mQ1Q+K5S5jRF1GxFN1V8bMo049z3ZDKJs
b2Fo/ETrzgTbj0AJ0uOGy5QjVBLrl0w6z6+CRmUuoBOLtNjO9mEqaXpwurKVuBHQVrkAs6ocCyVY
V8ExhW/ix5Lip41/O0ma9pG7w0i6JCDqJ/UXUKKrjzNs2fw1a6UQLvrqSlPbHSwym0p5T9SWmXvv
Ood3mAZSehlf/EbVy129cizSu2gIsGVvRZKJMRm2yUQIlhdyzA9c6WsI28oz16uDEtd4WldL71nF
PwONcSJdzsuyGbgdifJuhyia+Phut2vikLkeBV3bF/CWlm8mAwC8oMXhLMgYvr+q4ddxU0JMuaZz
5NgUV1olVeJLP+sW4wIRmTSaiOTnrQavDeJ8gmbkdcb1hC7dhGDUhjWbdRdEeJ7L6jFDo33EMOnW
i63qLFRx0eK7OLBynvHKmYytpQFMslz5gJmvvD846VibUe8WD6DCxphRDGWZGaH10h52XcN6TKPF
BpY/RZ7tJCs7DRLoMG3W9Zbld8GluxOL21f1p91JtNTqT8w8a4PViZNH9SPORwzk6sYzpT0745eI
sFqADMbvMDA7H+DK+8APmHlwM7LVTIvcdKntGU1mGscPTMNzkaU5sVcUpbd3u6WPY4ValM7VZ2lN
qm7UNH6CZAHH4eLp+kNSuXQ7+SomVX4CgbvDAKXlGSYuglc7oGdKOkMJAUO0/CfNjEwleflnGNRY
V2S9SoQEfbK0shvxiSUZOBzwYpFeIALhuwKX2BEOXiA3rJJB+axAlP6t0WD+PehIIG2ODWx49QV5
QTAqKvTWmsVVd9v+nilJCFgb+UdTg64j7mmY2Obt1BaKp3LW/b+4pck13o36YMoUSbn7WA2bw7cZ
jHqq3fT13Wa7BR7XYYsNcrFVqqkQ+B3lu+Yt2ZJKt7du7laU726OymxR37PhUAKAkf1eyESje1m7
SDmgbPpD78S1ARms+FWIX9hcziOTSEOKNZc0/gGBWViwxdOyjNMO1CwaLXUH60W/KmhnzxzB957r
TYQOWjx7L0+Bce02DbT+g3+MtO7ehHyvih4LUATjsY/fgPiWfUQwR7Yvv/UKR6YbCjyr0PWvlsQN
xVfmsgEsaYWGigOJrbtHnD7prP7nfVObyz8fULGIyAZiC+/cjg+Lh06/wQc+wTRmElMoy47bRr74
2tdGBrJFP4Vqn4VYMeZ8H6WcY8jkGFFxXcIJIqXnlOM1aJuDFIfRrrMsHEnuqkduibDxRMNFQTyt
4xsY1GJKkgvSGIiVPqKVX/Icb6lVFYBDKvMWJyDBFVo9yvTLIIO7KF0IDhuo6GSan221jJqF4Afl
mpCERxHJGvqF7M5f6Hx+G7j+3sq7xotC1+ufeDVuUWUrHwAQTEP8GVfF/4wq46K4GDQohHcaZYOI
w3LMpE/THCXEBYI+7H02EFWDcMpS/n8scvh5XwdpmkqsvhFw/DUZsCmj2ZLavjhakuBlYTy9LYD3
A2xYfy5t1GyN7gb92NqghRVxWd01KhDM0SMeD/lx+ehmoXzh5dMnODI5o0VzPMs+RiQ4nCR5ojFJ
Erhr4RHzAN8cGrGeaGGK+TSMmcZMkOub4ecz0kaewC6tCUitpmcRRzZP2LsEIhMr1ym9sckeY4Vo
j/krvv3ErV7EjEbkb13RB6ecGv5AJ++0PfX7TDyak/j8PlGvB3sxEw6WOoEpSDpoKcK6txhlnM+G
xRN1n23RQoV6UEtaKefKZe7aIpU+UcuRTE8mUcgBq5L8eO+EHaMkCKwJsM+lMA9nvvwloqOtylFp
DgZqANB92iCGQKW3f3Ax1xlMAw6ecA4zrragxe0C06NzNnvDU4wEXuH5NUwSR0cg+jIn2thwC1cG
g0bmCjMwJq8VyGJKjVvBggMgbbUSXsMwKYCIJDiImZ21DdbMsdCNyFjNCWISFU0BkaKMTNowZAz/
QeiZBit/oIJOc+E4FYT36SLapTO6K392qnfAQ/NwqIUsxM6gkF7uV7c4NGk7h+rHxfks9Rownx4e
22K0hRvlnAbrhJDHzbue/QJAEJhuzbwB1BPuVroEXL526V+V7qs0qT/ECwvkTXJeVjJahAvgm/8y
FGEEkcvl93tPGJoJBRSvTLcpK9Y6NxKs+sEztV9eUOKzYiCDTHDRuC9W27jiizQon0ckHKvMghoG
hRfNiq9YPC0xvxWk/69VTOPwELFzco8KCMLxfVyIvdjaB11Kl1MiYylvPvjIjXM75PN9oGLy7rpF
3lyRfw+sRgf/amxtkqLXOJNB2TEAkBPjZh6BN8WW7Y9bXzsVEbj3eBE63gGcU2f3ZTpQfY1IDhKs
b2KxdHjj48mlsZIVpqtADQ/7Q1ViU6UAY8Pkgw50rGOk+89n4b5SSCxdEztAejEXAw0d/74bueZl
fzEeKg7jg55vFgcRCqiEhpo5Y2HuqYDxFUgfhnhTePIUKOC0bQ4KkUhWeREo72z53JPIICx9QG/L
TkodF5ZGTKlAofp6iF60U0VD9SWDLhhUJkqbCKGJ1Xbz03I6uN+gIwt8V2SpJsqJBWT0z4d9O4aT
0Ak4Wit7153+4W89RwlgDQlbyFboBYIIUq/JVAaH0hznxl7jD0plMM187N8BnI8FjphJsDXRP3ss
9yE6ZIjRXSM9/H5FdoRZqe9YyP9lvBRHCC95LL3VNVlANYzFbAzJ38Js/eGcE9SFDMlP1DROLaK6
CuxSwUM+tc4VTKg9iZMfb4dbc6KYrhggwi0sMEM/WxNNUlew6slpY0YSfL0pxt8MaW9rG7bGXQ/p
PwDS1ZolvzrofZcHKk3FjHUexajz7AO+6HX3yn4RDFSu/grDyIO2LmUax7S5Fv9jpN37lWLYT2GK
lthsmv0RNT3jdvVV2PtlZ6lFsnfyLnW9vCKlF30hoEmdt8/oQR/epgCGdYo8tRb+/RWh9kxgJOXo
R+0nKUpNRlOh4OjAqZ0+6gdxrlz7DW8lJSrJGQSTNK+Xa4u4ktDEBpdlErGWsqE/cmYuMkTOOaFz
P2j1e3ciOc2gqmKL31MENTLVCWt2/NTF6dsjwhxdTJrWEwA0Ec8A79dHjQXy0a8JKsukQZm0SwLI
Hj894i8hkjtkwI3jFroUr2BoiL+5vJ42QETbvbohcVa7J92V1y4J+blURgECyN8F5uvPeHaEUZ2k
fBv1yGsDI/APqC6ErPuHoVSyukebei2kWbZsYV95BI31DH8Y5GVWaBAzTaOfLcoRdk5AL4U15UfL
PSiYfsjBq2NrkbgHcKdN4QG0Py4LcSvh417FRjXHvmh3uArLuqBUlKzid5bcOCP1NAst8iC1k8q9
4PQ5/XlU8gcitDT+sJGaY3Xm8VmLMWLts9IeKA+pyx2ZqMpUEf/oQSOoMtMB9kRJxvtW5ei2rY3N
RZ/UURes8QDjs8UVYs7HstssWUFvV6tdxyMFcH84ErG5vE/BIHgNLHFQpxJuXtjzNiHkSz2hdKCK
Nh/DjpvCt3/VePSl4qNKDJR+FFrQFXgL3w19Kgv5cKYy00HGuP6GrYn8Bf+qacGD/3xjAamkXmJ8
71DSie7unJTR+BzWG8QrIMQbQzxzpikouOenNNgibMVe+2YgQlvHhlB/HMv0RlPSm7Fff+AX0a7U
9U4rI7ecdQTcwqzu90BnnoEDVtAvanAq9v7CSkLPkf+e3acGIThAgDUOuPcXvhiGBVITtzGY+ErT
jfLi3fHFuu1fgWOdWOzztfLIEsGHG1Sc+4v6GXf83XShO12vYK91XdlwETA9Ga9EmS2QfTN5hFf8
0zvizYr8U0oUSiipbSNQbvLzkjfLi9MDdZuLKIrVYWzNUT4Du4iIYJUBPruRSviV9OTOsh4OpD59
DPcxe5/DS4JNMDaByasvfQrFWl3HSgNxE5J/vrom7sUkb444EDsmS4a6F1yWpet5KLGeMQYtxrTk
kBzR/oNqwj6V5RM5w5S9pPgFd4I149KscirLby2FzcWqzzySPPj2Nz0T4poPN6zac7d+9Tja4ObX
ZsDUxAeO0SFJgxNTcMXneB7YknTeJyKpbEHZYX0tMYWpAiDcQyJ5qWb7OAZJAYEDhrRgM5zI62FV
y1CtCb3arbTc1vGcNzIgWeAdSzGdIjHvcuDbqWU0gdbRyKUDZggK/k+zZ50eBp+HLK4lcH1Z1z1O
QqAl1gUuQy6uCPZO+hymh8ueh1IbVvudr3ojedAhzH1niu2PsXYzIxU9CVbgKQx8zYxxmXrPefqd
zQ1/6SyAoZ8aQ8nVSLL+rFCUeHJesMU69eO84ytnm28q8qxcQK2h8/LKPfmu6yb0B0oNQ4IOrK9T
RURzNP9py5Gn1ao2VAntfcJswqzoLiGAYYt4wXpPbtE69d7X7lPwAFUMCnT6H+3p86l1PJtSVfYc
i9N2LRy3fY/URcI2Ulkzf2QHpXVf4nbwvkY0Ji/YntPVkX4AZ0/OSPGUefiDCRn3i1oZsZKeMDOr
MMf9UJ/kyfWXtsc+4D8F2j5MXY6HLsxv19159zLq5yb3lCWzEZWusCVRv4MsYEy7TsXQFvGFbmga
RH3dP3QOe6FxFHhO5QfOoovRg/xFRgPZkecbe0tvv/SJtqEsLauiLp9m5hTlkiLCV+Z+XB2jBB9J
6zUY1vy9qd780JZP9+b3/tF31rhudFWpMiysb3CGAOCKYpJfQ+hzKkAG4RlonmMQplGy42/YnymW
YxhhrjOpD6hD9GbINihga6yp5AdpKQZtCFbARtLOdjZmq9Jf8fFjwZoDFhyRgme3rt4qduNzONq5
aFlJOxthZeqQQgYQ+9S0fn8o9Pz7yxAZb6iAGxtwyLpUcv9NQXgyL2O6iMW1rElHYMJrnBcuqpSh
7XmacN8oxR3AnC3K9vGoSl1ZT/jNWJCXK7ePRm30ctslIqqFj7k3XB6JzLv4aHcsSUyec5favwGB
e7XocEqTa5h8RfjbD0yjWTtnN0m9Vyvx0NwKNUuK4VcHYLisAKXxShow5SkBm0cacgnjTgyKJKd6
5sJTAiTACjquOLyNcgMbRSDyFzNcdWp0mWRg0ynnal6A4e+Ahx7RBS40B5gdBFGzJaCVZ8Le4Uqe
1URMQFIL5bVrJeO4tza3aH+LRS+YJkLD5Eg+RDlQaI8lmtI3J9sdvsu2XIG/tluO61E3/uM+4bFn
yfsfb77tItVIXvGdhpWN6rDBr/qclzdT/bIz0qUVsctcJU8Ob8dmonNUgBhJ1P/BGD3jAHukhzkp
V58V7KGW8FJXzYuNJwOEspvwDTxD8z4AncQdb+MhQ0sjNRuwQWtKDxi0UsZz+w+Q8zQgwCS+o89K
A+xnAb+21iUh8uuVQn4ch5WnYQYA5xDbLnxaE/E/FcwmPAErUxp7VbiIvav32M3ePjzyYg1cqBnQ
6FPicSDgUR7w8xzrDxlZLT6Q5Mtlfy89IoxNIjl91Pw9yfo9pRr4d2+YTihCdDZ1uy65ulDJivGQ
D7yQGIl1PPvioCygKBgd+jTm68tLbNiDMR0/k9ugqhhAEMsfmPJg5ilZqBBWjtpk/qSW2ymjjJQk
1UrSsi9HoLVB6vjdZZlYY0vfXQLO1CsdqKFpttOlmIDRwB6c146euiGXNltIi/lB6+ANGa+sbIYE
XpcoyCd36qclKVa9eZw7/7JOEvy6qzgXR67IYxqMfjisqkDBXIcE8BBD46cGtLWldw7eU4L5ByRg
Ly8P5SJgH97p0EJWEPwVB6SNtRtax+7pQLv9XKwD5MuzFf50kqq5+VYmPqtncH/hUUWv5OOorY4i
KTEZbUhrrnMUQZKrKfyuJv/ZKhyxGWwflg09AjivxRB9mWQrFWrD6EmU090sZPC+6MSLmuaroTSx
FZ9Hjn8pjH3fNJGrtv4B3viBOL+9JUC0M5HWJEXEI8shJsZ50wGm1DtdFRCSkHyBgP/6Qfs5gimx
JiiVAKPY+Z6k9kC0wkMtmkB30iPjiOL1A1TczUwn5iSfFDrr09GRRB4CoFWzpyHAe8SftVoBofP1
gWU0l47KJXUi3Kifro3FySkgv/CKwEnUB7KhrUIkFeoSW5CDfY7EY0kzin8Dka2igD8yRLQQmJ+Q
bPylfVj+26wDbIN/zAaycQs0A1g5Z9kU2kzGSw3OZ+uUzG49lM5B+ld72OZdthnEsK1Sy2Jb4YZE
P5OpEuBAAMeB+vN/hdpzdB98dUm46TW6ahrl9WCLcyFxvkuSY3mIzohcZC1IEi4b7oVy86zVi/Hu
v2QXxpCTcJsKKoQSXpCYsyD16pXSgqdnOFLEpdvPwH2C+E2bQov+DJzqsEQlQL1UiQW+8bWSUEZO
DvLe3AVly4TQUxl3bl5HDQ9mRJzFgNopukZzIgnXQoQR4tmEx9eYxxFAn4itmVlE5StS6Thvo5fN
Ld4aerTrLAewxzP8CoJXsMjSFTpq13xMAWI+dK0gwZiDYfQrIJ6Go7Ea9f5Tf63n7aD82HapPND8
v/fFZp+SyivvNiJHV39BNrDXvpel5rTL6mbc3VqhpcWEhGIMW61SRfsue7oESlaUf9TqsAasYvv9
5Ym51YZb4LXWXlcmcbkEYmB0KPmhvYHykkMluCeqYnqzcAJdbLi8mSHOVWdMivgOjJZlfHvmU4Q+
RC2UNTmr77WmF33VRH4hIYSdXQBaOsSyhbVWHCOm98pHJACuJ3N++bO36DOQCLYRylbOXmclB+91
3OOl8dQYfC++7XJ6kz75op3afDT8M8WNt3h5g+UK2g7LIPd2LX1X2VHf8XfBFtUnhJ9o/cN6bGb1
YjpmK61626xvvYidypU3wHxKV+2XZ81zi7LCASy7ENOefzKqTWjFOywqbchiWfiEQzWwsmqDBvXn
8WEhetYMFCmfnl6xlPLRrIAXEZvwrut1MMjxmvD73dQwasgiDTC3UfiVWa5DXlc+/a/3/Og1fmL6
FMSg92pMwq32ooOycUvXyHacW8Pl/2shaHxAtcjX9eeqW3uvZuS4nKBk/SmaJHmSyY6qYBCER5uj
m/G1CUC2ENoc+YNdVKOAYxSsYOLZLTxiYy1b1h7KXqC4DEoPMs3WCQonshDogS5ESHiWUNAZAOsP
PfKto9DYycowrnlDE202XTUXk2n+fTqqfPSqS16AlcZeXC4JKz3GD92JTK2zBzD3pWQhLbCpsgk1
UuOl4hc5yQHLK8maQzEM7Ua3x0Y/o/iV6dzXlFlzM3q1AZRM+uXKm46uHQ6PgQi1bB5j+z9HDuLJ
IcFsRg40ahcW6ritmB2CNH8IFJMu0rDVUhFbt8tAOCGHqFAas3LH6r9UZdmuD8mNk5MmnuksvS3f
1QyMZSp4d8Vgzd0Gxd7k2eWUyY+xaOKryCQspiCSVtVv9ND5v2FG3Q9G/nrR1s2rCxBCK68S0fok
k0lPmLm3rmJExy7BmNNqd6FeaFvdDsI3T81XIoKmkI/qgY4imUu41MSFpmAXvFIRE6zwRBV4pBTA
Z+j52NO7iCePMTBeWBC2ODCs4hji1vSRgMVnURgqUWFAKxD+8XdO8lNKZM+0/bPF/CFcWOgjl4wS
1FDrNZgJltJ+3NiRkxgGB7Ctf8oPx64JjPH5+nYl/PqoJv8+EnJt/lLEkYMt8stPvuO7zYDaoC/A
FJGZ2LLtGp7bBIrXkGycg0Aqyn9mZ6B1u4jQFV218R3fO9lgBxbPxbMg/9k22o4afS+529iQDRjT
2FuwY2G3CmIhq+jE88HNZMDHCQscWOReKquxAqZ7mJS2Ye4Hj15mthhIZKbSq3ZjWilz/Gz1lue5
/vGGi4MxqIfamoFw0BtweX17/3OW4N3JEiIJyYOkUQjqIbxQZtQedELTg0woGLwo28ma4TmKkoZm
BoQxz9KUnhe5DoOlOfyyUv1jwHGHdbectn6KE0OT9UN9gaM4zC7Z5uobZan4xEfa+Pz+9NWlMuN3
nUEthSj6czUHpyVzVMMMbAQBYq1wZpX50MWX00Kw2lyuteA1womH2kXt1OXadu1BrbXHFvKEGD2w
s6DdQTu+3+Y3luWqOi01y0hcTU+EvSdajYOnAuUfnDHhxydsSWJDcqVwkVATDB2SMiyX6Z7SSy+j
R3ht/KaXt62C6ogSG3GeiqwwgeIr2r7NYw6HpPyo7cMeQKXH4dHEXZvGvs390n1ElkubDmJqIOTF
fNxkoKpCscHftshnRakivSmW6yWzbgeb9Af+mQbLgQhqW/5jH4bvxCCjpCnlpzn/NdO8Asykclku
u/txD+MNClUzWSkfyTv8Mho/vQy6mqYnNOdbQpk0hlAWvriRHl79Dav5lEFLjps+rZ5fWPBjHAlu
+T2QcfsSEoNREB2ioR0v9WqCb1Weld1jNF6KYQyXU6BA8kporAOtYdNVw725ee657lXMRq45ubEE
pJnU9RYw47LdnZ7D8Z3yTJAp3cRwINh7wTl+ogJTxdmoXH+qK2Cx/TnnaA+bUAhcsjVnaAN+BEwP
G+WDFt+vxBk6Poka8NwQZ1ekVSXi/p0OMxv//VSHY5ZSQvTrQL6UGJsBfHUdZmxrQpMLj3gVGTNR
0t42WR/GYbYd3ewC7f/MjIOHpxHWZwolaOBeuL+rUjcbjMIkfp7MFEVSL7uzVgpMh5YwuZ2TUOLx
/K3D1SG5M+6+gzHN9OMWVhtWmCEywobEXT7ENrZ4FH5I+EMuS2f0JT+qVPFLvclNnd2xjBudYx7t
E4huR0ZMpqu6HapsSg3Y0QD12ul7//fu+gtg8nnFcSWzDaqUgfZWf38tC6hiXgxrpuf6mdLXciPP
rtZeUh0VN8WWsPMvpjEyfTCMk0Q+GV+bjObP3K7EvvBPEZI8vdBRjZI6rQffkaU0iB5CykoC5UAX
QRY+TZBJTviXXO8lPMeOVRPf45s25TP8XFiToImmEZ2knw+broNs6wSVyFaR2v+JW46LOSY7NvnN
jwUWNk2mNe12ved8uqIEnDlCK0PBgdNcaKgKxoMFLgNdFcGTQubu3XAmWw8y5hFnhiaCDAISqNhw
L25MqcR/tqUbetNo/PwIZYpwJKdaSyYCZUUka2iECRfIRaYg+M4mlu0RLkNfmHIsqeoWUYnFcZXV
/yYzjw9O+rE2A2WrSD9HLBBtCzuUOtq88A4enHr+8WFsX7iwAiFjcQSmduXVXXmaJMtg5+NnbIqA
nTfxn+HyeztU8/wr5mU03L5TlMM26eF4OT+kkZ5L5K6zyzby1uF46avk7SCbaBEk2BGlnSwrfsoG
KYs6QtcJlugFxK+vujo6WoxuJG6rJ7utlgekLYZiXppqT1xFwPCYb6pnPVos+32JJXSu5xfo/mgw
5PYbufnjnAe4w1yaKNrOjNbDtRwQ+mTNtnJczPwEHNYmjKcvAiJfMqwPaG+33lNp41YFi7cfoXpr
dOFg/MVWcOEEAAk7OawA4c2yhyoICZUhkXo9fuZlg83N6FTY8aY2FwbJXCnnIGCfmWk0DQIXPn4H
qgD9FvpXbZgL/BJjZSWWevw+bRNSIwgBC98CWuEbsgBn09xGFYgBAa0scNXs97CTK6NA4ntCZh2N
rik9ASpg8wsh9+UTMfmilngFzyxZ12+w5o3rSYIavpeU3uzFAurQy6KJYk+Oz7tGYuIfB4wT5EXD
M6o3q56PWuMys9+JUKPf9byTW7GlgYYhgQrTmtfmWFq60hQD6WNs7wDjkDKpaW2adouZCqIaMN5/
FfW0r9V2S0/gg+kmSAN/b8rxp+yrkERM/jyn9yTRt6Xy8z1StiQUzTBG6Gc5bknNohB2CdNsY/7D
WIJZF7mvJrRNosiJ5iZ8rNuTDexPKaDu5SgUEcCxtKpb/p/gDxoDdhVIY4R42MHsg/HV0FqP2SZL
2k0cLaRqJdkju1StDnXUBHK7igZ7JKt9EI/+uc+uhlI+gS9gJRm9drRYKWsgT87gjqyLbjEr5vc2
5jHiwyh3uorG89T6hepLHlrqFkWveZzfcbifzVUbc1nabU589ZThHPGPyck2PWOXhEPVZWcRBIFb
gU2cahkHyLkTLs6YHF6YSTO/PfVMrrqOghIgEpg7k3lH39oGoxJrDrZ/NOSCCAF9ZRwn42Kntil+
NRo5j1A0jIpkESzaKRiOFimPYd6sJ0Wp+2HbMk3CtFAZj1bXxM02tCz+n0o4pxwuFeZTxx5Ofd3M
DMjHXBZljM5PiEj1V8hMygtx9/+qBRNr94GHEVGLUSS55B57nsA54ZxNi3lLQg6ZbUSadChH/26E
l8tO0fFhxgdl+UWywHi4TzffeGkyYPXfdkFRdOoCz6twG08BXhKcaizKZsxM9odLLvfV5xNWCKjJ
zBeLVv5Cj6KXShgp/JkSfQmkB9xdcluofJJoFohcPYB1eMDJLVeRIdtOgn6QaKwo2yXsoMVh8vI8
FTcX8R8V35pFkitCxk4+0vISHaLz8Tyerkx23z++ooGMl0aq+ilH7wiJIKSbioB+rWCaD508Wi8z
b1RqgnDMQb1AJCBvJkPjlO2671pE0P088/7+JvUhNqGS0gfehAFj5QuCKUMOrmw6VSL0I6T1oo+M
kD06A8fgXCdh3hWzr1sHJUvrvqDW+4pPozoM4wS9sKE/Pwt7HNl0VRck5inSJi+iNLpRvo2hDlaF
Em5GBXqDzY9VbvpQ0yt55dHvryUc4GIagwVEd7/TIGl99akBUKlnDt/ktl+/7MnoWzqRQ0F3wCfc
H1dcD8wGQ6hYOuBQdHlWYxbvAs6t5OYhuRu6Bsf8DWOuOlK46UisXYh7MGeYIPr9tanT5wraeH4N
w8087u/++00wa5Jazg2r3Cv9U5rvQLEU7rhT9kmA/c9YcFI5udEQ8iSPM9Btsl4fLIP++z6DlDhc
eLMHfa1w7veOlpn3u7/Htjkut9c2b/8LF4SFnjvG+vue9LbysuFZwp+8xe/jq+ECownb9DDr1cLe
qiD6F+nVE/h8PCfzyQ7H+ZM32xZaCYAdK5oRAW3lcqpbG0z8kXbkienwDNjc1LOvHg4gwdBVRZLL
GV76Qk5BjATmzIFmnNuEt05zr+Kzzvj9F0E5iPQVPT/4ZhfJxcGVWZ00pKCEJIl7NP85eDwpuo+1
USJDUiJk3W8LdMTlnyUEhn46bx2e2MOQerwzpXKaEfoAp1RTyY1eyn+42broi1r3nNwwPaHot0hX
KbczdpdlXAB9QBy4lZQDRVRyJ2cY1G1w0Iip9BPURJQMd4/sT7wQFd7So9/XFHhngfMlOhdt9Ncf
Y4aYLd25+x1m3cg31Bb0+OtnaPsFnlMIwWbopKq6HnYG9MjUcMNbKLtpFtoJ/hO0nhVWMtDjeDaH
md3xRJteXNKM35CyMe87Legy03IQihRR/2eKhNrK4wMoq5fGgYH78bFLyjevV+CSZmohOXTu07ud
Da3lp4N1cPImPhJVpfgba+l7UDlVhuM/+qOaF6jWrtUhZq5dKOzjKiZNXjp1yoppCUCu0GGkOlVB
VHpD0dB22fj+16MTALXGZ4ShdhAZAwdYYiPaYJX8DdEU89Dk+YjeSdrzGvLCixh0h23TjTbt7nRc
Xav3qAuh6ojZ4zRdMP71Xm0O62J3z3ZCOR1c8nLmo8+u6Mb68giU2avYKIDJ4XXBJmzH+97LkdgQ
7U/MYaciIaUlXGi72gYAUiANuUin6WmmXDC5c7BbngJW6n/EVrPKwWEw7fwf4Jp49693w02e2mfB
q3nE4TP8eH20fLWyElCCuO2grFyB7Z7W1C9nh3WBNV9eAJRC7G091MQnFc/Lo2yQMQrzURPlA2br
+a1cfWdG11uqD50AUubw5VTczs0rok75s6grPU3zTYt8PhRviCebrHhxCZpOxf+iFnP7ZpVLjtx3
oDncDPMeoUhwdiOs+PPQn5IQyX6bPyiYI7l6zCobLbA5TPM0KEetEh+OczYvumJVDNgKi1UxEDGk
cblx/7vbCwtbmFoi/D9xcXzr04JmjFpsRH13pnwb+WmjC9w4I2QNYbKiRj4aRC3HunNRBSGln6MJ
SNwlfMuCjBnoKrka/njaAjAMzLjlhIWA6KtsxdGJdsYbcmI4MMdrt0b6JWrKdXAoQbKjcb096j5e
B6IYluLhrYYA5MjtWpkm/J7PxnpnFJs9cZjNL9YQIS4wQyL8m4+2wb5ihQNkf6ccW+DCm3JYDpF1
zQJWDV6rwmkjPftwftjkEtjqLahG4Kg784Fs0164fpgVmqviyhx6YkERI0/w1nvLf/I6QYORex6G
+acEFeBcKYNY+atVtm3rxERej+0dbv7OSFFhGgzes80dgUkLQAgYT8TBpSnx2/DcBQKxOHnJPfw6
I1jmov7mInV0/jw2k0BxKwFsCzaCaDYkA1e4ec9pTmt6LpkBTQLSw0dnU2Qd3PpzXr4IFufg9WTk
AuBT0MzqqFyMDAlxnGiByw+98TpDeGMYCMJQCaS3ZifefnA0GwANMl7XqSRDGDySUVFDd5omql3I
2BNwJzqwTna6xXsf5C3WeHfycpdiAK1CgYTOdDwhFlc8yrDGxooGgVKjs90dNK0vU7LGuZMNHe1U
dOyq1mClZWp6GcdX3QQwBbpGidWT1NQwBDz9FC2CunruVAcIFqrWV8vLORHSQUCiV02EE5KRWNbk
YUjTZ/zI7vnlpclBwA+PfL2cBCEkatzSYr6MMsUege3ixKC2G62Jke1kjKL2iezkSzweqjwOV7bK
OZSoA5+NHKkdGClpevzLG6WScqrxu2GJatsqCmexb7GfAXrm1dFbkHXAI8LmmoLUrm2b4Yg7kzpR
+BAiJCjAtmrJ6TleRFl+mHDngE74SD+Pj2MC+YUvAwh5NR0jiF7hqapnv31cApzNy07tWnsQXjbQ
UZv9aoocC0uaOROAJlMDQDS7ucVGq9UljNLeVmjZk1HhAUFspqvMr5L86MN4dHp0rpTpXJKmChc4
bcQMhMynlMDQFfOoGFT5jgb0zDyRN1b2o2jXO7/PlIx4AMAU8nYSfHt4YcxFIXnICtZbNLFwrn7V
m/ACdxqqZntENSjRoiWF1tyzHqdNFTSw5xdnhF8lesGdkgHhH0qqlmzu85l+Mn6dm1aEXDfOwdS0
6TTdgwwQ4IUAaxwNg39WMLu7txaqtI0K3UqHdCzg0aAuQxxW+5b6kaGIunoJ0in1nGAHpA0bOrIR
QxqZuNKB5B3+PBMUGDBh1aGH5v/I59VxNKdEJJXrLXB0mpXhC9R/ouwERc7Eie62Tbc9HODD5jtH
W5ubadR/C/SMgA5iPJ4onJuUwiHrWmpZxhSmTctDE0q7eG/B1/S0XjCuKj/gNBsNu/hh+MxFILIM
N9E65ZpEH5kn6tY6MI8P2zRZ0F8NXL/o5te4lg72PX6Pj4h6Wf2yeA8803ACijXOM9kW7RaX9itb
6+uuAqA2oYgU1Mw8BtfQUNDkyPp5rvY63RdE3IwZ/422aO46CqDQwPnefR6/zU9k/thaHDRLaXzu
0rsP/En0KyYFaKSHZLvD3NPUIhKOsXkmdxLv3uKKUTNjck2HGdfMAPvtFLSCZJq2umo1dOp/p7fw
bO7BTR7Yr00oQZwfQA3FnhfXBoVQNIQKu1lfk2tworQ5J9ha6HvTS/jXeMJSkWIJRsJcMTUzWvY0
J3uvmzbtbohGPfpZcAunNy5uFFLXCL2A7SbuSQ0sQNWbmH4NadEUHBmsW0d5CmQqzttSHoiTuC9y
Eqq/WM4GQLv0dGykF9GtNqa9fmFbfmedHdyvnfOsMA7x2CKu4Hij0PxcamCwn+a3DkPNnbAX/kWF
TNY56X3E/0jQP2RJvK3GqeDWTgrq153DKGV3ULSELf2XINcRj7wMWgNJMuDXxD8nIIstCLIyOwGl
eG/RHFCJP7LIrlZuGgT8l1+FJxgdAdt0Ipomt1fCiMVS+iHkScwmrl/mcX0hyG0LuPL407YIev2u
9ruXsE+mEEx9U1+kCHEJ0rT9eg5p+L+jIwjzzyadsCT9+nZ8GzQvVhLEQI5rTcT1S7w0xOFIHmh/
eUB8tXydxKCmbP0x72TqlG4vGZK1Xfu/ndutAtVutuWxZRyEqMYVyHqAaH005RZ5GRJPVbRhSTUp
Ugp3w1VeRcblE6fJZzUUZg0+O7zKMSLO0UnHbxf9Tb1BVOHdftNwERtB6rwSU+7KncdzKnX83a4f
uFTAzCcjLXvaGEW0dJ0oDPv7k39jEZfLzVOpH591ilSdNB/Ygcm6SLrNUWNJT9PHQg5yklJVxdSF
pkykCK+a28a0853NfOhpEucQTlzz3Srg1XqMM4AV7YcadVifuSpr7AYbpFkqYFEmAR4cKBes5br0
UlB0uWpJhM2TWCLzpFtP5Rr4yzJpnaazKrLbODmOFJHQeSra99nHAhXNqTSGL0Eij5JF3s8zVns/
vrPoBWDRDIwnir/AWTGWj1z2MRHxi4JHMVfWqKK1lu+Gfa1MScBxI60I3+IfPYC9xc5O+FMLUKyY
l6vJAHGav784eQNhFlC6Q88O9SsjoZjgZFO0GQHAykVN6EkAfNVmmxlRVnSLayAc6n8LmSnUp7hI
jlwiv9OaWoJB1gqpwX2/Fd570kHx+mP213rB4Nf97eSXkC5rdlNX7ormIaOELrdIeY3dP/Y9JNYk
aspS/sYq7OVwDWg15e9CFmifhVtkEO6TGHss0QbOYZrFrP6v7yUj9859Z2LaUa75eJ3hJxFEKlbS
amVmrBhuGjY1u65RSLaR8bKJThquAFm6DeZQEBVQoR1Lq/woUyym9bNP/HI0qf9Qgtrcbtm95T9G
gindndvao0Hy/mZ8zwzYwADTkyodkBTUYkG0A37mFZ81TCiKWchx6yrzZKdDv9BfeR/F4HfI86rz
RQFKf1ZPaAxpBiDJ+vzXYWBfn0Q5NqZcKubtqYETxunM1OO7vJHVVCfsdXZV8g0hUxB3s6s2vby0
JxO1zKTyyRo+LPnT/T/UEAb7P/nyRobPT5LtL1E6XJ/CujG4CqmrNhNzf47MO1VbrxB/9B4lR6Dt
ruu5GcNeVoRnwtTSLOWHlR6WFZdgqdzyN2rAISWXCih4QlgYdl4lcGSiEwRpqHX9TOLw3UFq7n3X
1uVCY/q+9kBJ61Lo10sB7PORY2GgT0uIVer6617JzE5iH3ryrcXDjPBVK9vgGE06a5S9y3PsTdFE
SfuHxie8xCPtcGiXQfbQer1Adq8i4Xnt5Sv440uUGAnHdtGzoexIfPo8yDxUj0GpbUnVLbPQHvWG
aUGLMxq/2mMtbGZbV4wzWToJfbvGZ44GRE0YR9uaBbipdAf+LSVjOMNu0jPe1wwvqEcmwV9iy9KR
NN4+bzCYXwzIwsj4jse7PUDg23pEQK2A/9RYyYWDhbiNNQxXk48B7D6JwqpHw4aUalw6ozYizC4h
eX1F8YVGkUGiCqFPlHzYZPHHbzgs8OsZelFShx7lQPhgvZFTkuSTaKPFmLZan2WieIFYOJv/JRBC
xBwtkbKHZGT9+zdCFA/bONz+zxNNM3Iavm1KqW1X37rDrp/QOlF6z1qi+itAtjSPguY5Vu+rjPyg
08psrraK8x6r7BcOOJDA6tn+aS10jtvVYYtrRLyV/gA1GlIgpF2lvpU0X03bmIqssXPKLe+hzu2J
Q68qL7BGyZ9Jfw3fDMEwk9U61vwm7VaU8CvLE+7OyUuO5XIJCtqS7pNSZsWTDdTzhf617yceI7ua
8NIL593OE5+ZvJtzskOys2fzeVQ4eysPQemMsBIcEIFQ+E2X2hhG1s+7NLepkVR3hVg+s+UdI+pn
AZLOG72rBvuYT2mxNpcDDgPeI092WZpCMXjG0NETd1knZYWggkg/Cwl1LespzZQ5Ub8WlL6M+Bvq
NOEwQ2tnjMF4/TFHbyVX6cHmcM1NDnvsZrkkFkhUj4eigB4wsue+OEu4mAYuufWyb/xNc1IEZG17
E5E0/slNS2fV+QiXhOJiaqnx6Y2NLVy2NqdD97Zbq6x6vdDSQE5E16tdlkMYVlGwqoT2uXDMZkWW
sPLC5jjP3ASZbbhY16NeH+eeoQz7x+XHBXBSPYjXQEANeCEloDKsGjMCgfu/08gNDz+wvx+6eX89
nEw59AAziAGyEPvUsSDr1bhOEjOvvpQdWapuMI1kpfL4PouMHu/xhoKIbdi1kzss73Yh13N21J/N
R4jPr41Y85qGg+y/anUVa3oa7FYA6OcWD9wJk2TdqXpvkLrWLQuy4e6cO2GZVgKtJQ5G8umcjzTX
V7K6UfiA+ERTJjGA3bvq9rCpl+oS+K9IHtFCK7SpHhFUOJUf1bxKTvusSotqn51HFJ6/AUbILCy/
zIRry0O/+0mIWzS9lxTVxgbuHqr4+ImohAj306+nj3+Q4KO+djW5EMtexUM5wCkNbhr6jUNDiOLd
60NHnYIVKa13YCC2+HnS4lTddg+PMGuoEgy4AZtGQsHm3OUhQq59575DTgrr7i9EOBaGrNGVJ8Xy
RaUbyDva4BLj9b+vLt42TeJeEQtXVskjZhsXW2QuFciHFKmxQEtO/zB06c8dzC5ZaYnXYda9ndlB
V0zkW2ANfyf/+itbUN97wG+HbV9DpnfvvnsL3jI5e79muASp+eZpjWpCSh/lV5oOp/O09o4MR4XH
w3kIOdiBBkBmeyeHPb5e8SxlgSSRBUnK8lzXQnbJySHXgOYS+FiuLxQkBpMyA8YR8huTG+0gbg4t
3PkOHwyQxii5HH2d5DqhJmOQipzR+jSfsyM3141oksctokzlljy5oIZiulvTQwCPchMfXtyxn5pD
g5O724DZQF8D/yTH/PwhlPY2VHTyD1RPvF4FGoBVmtt01Rfezw5sxBNXgXX28oXYI9AJuZh+/LQK
+4PIobt6lXLyrxtY6gvmGi/lAhxfkphr7D/fe3KuZwIpqxcDd6OCHT5yxnaCRCLfB5En3D/8WnOV
BUbMT7cr4P7YvEj36usZgg25ZJSmepCC6cCgvjDSKIKiYShN3Kue6nSpUkaXcbX734azbNc26o/l
QVszRKInQmy7JkB6hwK5EQ4HntpT6lgWq0kLbdWiKLqaU7gkmbitDxcUvdGSJk9WWIObWoSiRJuY
vBSgao4PqvW3tBVaSyUPqcdJ4uvhbk169+xktkaKP5hraPb5HQbXnVP/PIsLFn8JU5C0YQByhbcX
T0jUhu2+NhNGwkBY7tZd3rgRDUz8sWvBpkEGKU61EyZvETa/Z/4Tt0OzkIyCRDkkcq5M1ROpz6d6
vk1T1FDjwuMzZ0ztFDamayEcr5OYwbDm/srxSPU5TN0hFKQ6qETG9wM+vQxJPpR2RAvIKAS8+nRs
9S9hjlAzMmV0TPAh0Xu/Wh4/3uyiSS+pGXTZRASomORb5FBBFLj0QnBNzt86hCrzA8vZJupzY4NX
AHmbKGBiUzpu92IlvGnZUMI+HyZigSGLCHrcnir6PjgyeiocSHfjQbG9JK1gf2pkeuGf8w1qF/dK
H24viFciq4T6et6MBKK9mWkMtyCmkzmQ4QchJFRNG0iWL3yihyyEUsuJXiwr3kRmVuSXD2FM932U
FBnA8NlzSXjPnmRTcp8WmaE4qWWKE1xOz/OVkGTp+LasH6l+lXCYSVJTAPeMzDnTzKh4DWO53Xki
0rSypIegD/NEj7lpeuIE5o74on/KvWmtm/m1LfzaRvCeozJRgGPlBdM/zgPX4jZSJkGfw+FwfbXM
hlWL3mE6CaROt3v2sPURjrqtlUtkHHJ4iOs1Hsygh40cR9o0yZcNSq9oSL4lG5T59G33b9W9uCEw
zpjqTQdf0cvhVt55gEKLcETYAZ4R0TPSQt+n1UGUGWDXdU+KOC5VqfIM7wDOMh3vtg+fmCCQn9Ik
QxDoN7NmSohXVYmgP8oaHOhWKtzl+sknU4RdN/9HszHuMTc9lp422pI0edQfLDhxl4I0Hgg5tPR8
qlnFmkduVSpWdriKsHZptCilphjK20w3AEpIw4Ga8BSSKnKj/6SYDt20jIVTZtTLodZKPsVaHDg+
ulnIuDuGl11JVO0YbYT18ZromviNJ2J/RvYvRz/oQZktj+fqQriwrJ2juZftZyVcmgy+tC5pgJkI
R/QRUDrd5YtYYp9oaznFSH8+1YJrrUw6V6MhL3z7QOu6Laj9wOqalzTNs81tGML53e2/VvPzBJqm
3AFxyizgQ8HgmoOJdtdEn/rdkbFgXHk0eqEmeK3RAKySktyS4IPbf5+D0XujfovP6pIbAwD+Yt4s
YZWmLVDqvOyNfNY+GXA20bQ0tqf4ogIJaB4jye5S5k4j/OXt7K63i51Sx4aLudUUiflXj1JfHP33
Be6Rc2xSQrtMxPjcIKKxPaHeS9TQQe+8QM4UxoeILjuPpI4ObqaHT21o66xapvT3bwCUfuEQTs8a
6e/1MN1q7q+Zc5dIL9RZPeG6cwQpievCnG1rvUWZ0EVwdNx3VO9MXUe+wNmZyPxyyIcJX4Ai06lT
jgJorCcmxW1CrpqbqzJsbjDB5aGu+MHLgUny0M2j4qyB0VDPqrpU85XF7obzMeS7WMFQvXa1fV5/
MUr29UT4JjY7jxLVNsgXiYNZ/SAHQLIhAS9xNpozoFakOlSXCte2COATjxNHbe1ClMr+6A6EI6Vb
2BWPuwVSvQSyBPzcF1tkf0aRDOnHw798uPhs1UlKEzenVvR+mg352KDf/UU+eATejurycQ/+m8AC
jlblAk6wHyf6mUlXpazDo014If5pStroJB+VMRBUSlAA752afA2QHulHDtFHowSiifRhfRNSObXc
lVTjruyAL2OMSjxHBmVt3LyKIqhKZXXpraaP7QkmHmvHKm5MNE7ZHsekaEOX8wYz3TBtiCv/3zom
idgkwe1xoy8nn4MTZE+S+k2BMNFDJxUCqUN0c0wNjJDYZgpd62QcNkBeC0Eh1Uac3ElvVas84+Ah
UCMpnPJscLThza4aXHIG6fkBOdQjxRwg53MLwvjNS3Q4839QrAEYGyhb885YmhSgF2mnkWfxlt4y
J7r9uWXAY0hR/DEaWIDkkSj/PiclsNqHQbd8bIzHKu0gyfgSvUlKGvefnm6sXrJdUqHMElSIdtV7
KEfqQ1EGDIL3hwQZPN5xyE/wcQcwVHGXeY+AnX/ndgSTOzwLs5fe9i88qJLmGPwFWLqrbi9mgv4O
eVOGmHxx9s00CbZlbt2QFJwCwcyCz87wRKxPQHA68wIsxYMkXDdtz2Cq91V0GZI7J0dhlryATHYh
Bfk4wjZftuO4D1X/ech4iKnWrRMqTazkwISvPEQpHSfF63ZSWMdZL/1S7Nll79KcCWoea+Eyz4Sg
fQa/F4dsj7SzTYLgovEo+qOC05+TLHasH+IClwcEJH+mw3cja1oTET4UsaRN6oDKrN2TvhUEO4oo
KektKVU/gyiPXvAM+vhUw3R3VUsJQe2vmT6PeoOdNKg1NA6ludgQBhRHTpqRPDxxWoeFcQY8u3+g
Vy4euncwsPbKK7S2pZ/M1vlanMCKwoLu5QGPHoyxd+Qj+iq3mR6Ka2RogbYnwWhLiAi5rfjidpVV
r4x/tQbpCHAykiGHPJc20qgzfGxr0/YQH7vSV3gPr/oNiyrUaEdcEGxuJV0mo2cFIzZpBjSYQJ1o
9TA7n0rj6yb2FLJj3baat1DxGPPWrUdjM0OhBXqUSZ7EuXRQqIYyWoEoOtEQ3QNP0ybrfH/VLDvF
zAsYPsrFhhKS1H4bhU6P91UO6QdIApjDaI0HYsqYqNJCPmd5BnqFOM2ZasdXcX4dz1zPmCqEPW3l
1g7e3cg/df0zUrQP21KoyR0HDrtWEua6+/vK9Rzi2FC2UHLT5jjzRHjkB/MrbYp76mriEFlDQ8Fx
PMszVUYHznplUh9niVlcah5AVmdxEHTLIl/8nG7jz82dTMawDNU1PNYJUvp2Cwz3qFBffAdRx5Fr
hW+PJtHZTuWrNTcpEbfZcXL+zymaPaHqNUczeXjLiVqFc4SzbBjDLU6xO+WA+OpYsOePdpZYmM9u
veJtnIY+TdLCIuiqwyPGoTnl8WQbpXHqe1W6LLowsPeBCHG+OBKHAg/4O/KaJzg+r6C2Uu77T+tK
cAcbWkIRNgJY9LquJvYS/n2C2ssKbnke8GF5Es+AcmUYbWg7cmTL6lecXbZIGXhLlpu2eYD4H1Cl
+Cxk0GLmYJvOZbRs3sb1tCW7R8pUtWptGXoD9II738RKvegfm+A7M/PgqdWWyOFQpUb1qfJri7Zy
ZBm4ia2sGfbs1g8Wv2M4JFIFdMS0YZ+lWSqosRrufKvPxhDoeaadJh3fWMNm08n00z3wkOpORo8T
SpUX48PZ7habQhuBgNQwPjdCRoxatzeeQuvk2oILtvAEPw+EMo99tGiupPLtP9hhVkkXKKuXAi2t
E74gtdmRMTqSZVFJT5DwbWKjYpkJRVa3IRQdYl+Sb1O10UB/PLt+thpgk4pBeq5PVl2rgJe5Z1Xz
ZV1UDnpgXU8JGUGtghxSbmOHdLZbSBeBxZnq3Na/brLcjBD+189tSZGjb2S3t/SWTg6+2GJ8rPx8
L40XkamyAxYQDIcVk4tCjzK7ojBUDp0WScO4qf7TnOmu2Y9q7TLy3hcpfBJLlk6uAYq+PH1QAPw7
qXz/mbVGY/AqEakACcSjREE043reWfrGX0mJDSM0yb+d4mmJOctdLMN78CTlWfuSL14M4uj9JT1r
wTiqkSsrkVo7cq1JKdf+aMeOp1Wfirrk/VjDiQUExgzbK6iB9/8sPnAoi3n2uGczMl0miLAVkxH7
B7jZL0B8LokeCimfx5fYsNcLjhh1+BIaBx4HfLsLv4MQ/yynbxnIzUH8anKgbfIAk0XhlBvpnqvO
lIkJaf2w9MsWYA8Y6cpylcw8uwgOkhkSCu2re7mwIhvH63m16Dbbddegi07Y0bj/rq/SbhQ/Q8ez
4Nm0JfeZHoLGbOSJ/XH9pSGGHyOHN5eCF4WmL0DFxCnJm7+QXnI+GP+w8da//RXkgQKuUxw94L4u
6YsT6SWlDB+/etv1L36suSnc06BAidFjlZna9CASBlElSeeHP0DVudHs5EUOnQUH2Bye5Y2Esqoy
7wEdlrsvZU/NzooucUWKLsUrZG7rYkIXKHwyVV1KJMxF33wYt/HlTvxM6iUXOjh9bI/1Feg/9GK/
lbIuf3oVw9VvsaGquW7RaTeOh0wMlzRqh3eXeiYkEMH1rivCFBtIvRVTh37O/D6a6yg95hCI0g35
2XHccqmcH3WITLr9gAVmqpOGaVIdn1abfCkPRiaVbW+xMOfCCsbhFFT6eNp8xW4g6cgEsQFzuUi7
vG6lelPg5M+mEACs0u8er+v2oRuIJm16bKf84DZrCqhr534iYj+6+F/gvb7388YodXKVIGKwf9xk
+f+O3bcQL+JTTOUeFEYPDAof/RjCVLmzIQJhn8zJyhJ1KJvK1B6q0cq0sw47wLHKnc3AEtXqhUWA
4RlBWLbsIlHyljKwhNq0nqUZ4ULyOoZE6qMyrODlJmKozbhcidnHReYu2xRHJS/XhNucKBxUHYdC
3chcgTYqqxQ1jv5M/oIt7/WLmVqajMAMB0sW/ZEPNCTo0xCREO/PcYNBtfHUw8ujHdFDU5TKgNwo
J9ICoU9LfEJQdLjGh2OytQlAiVwTNdx1C5wo2qcIczSNTQwtOCF3alH3VoBnHMYvQm0hXsUnL6D8
2ZPKOMIR5695xUzGWyUv5Syof581Twsz+1QHUQhqJBE3RCngl7lPMbtLcL/Hj7mJPY9svELjzYdJ
IkQug+sckfCmbtaLpeGZCQfa0O9jjkjrYxotp0AbYPMt7Ihfp3AZjJkekNH7VZQCjUhZHuUxZcij
XEiVefA3lD4bDT54cLSIMDm+MAt6V0No1auPkwKHupGUSQPRVB9Jed8E2dxJU3pY7LrguhSnEMhK
6qqAGNvNCEFPrUMWoYWn6sG7DoTC0Ad2GjK/PxK14sljo+82Qd4Mok4wqJNnAlrrceX5jDghXl+h
+3tXsLXiNFtnVtWZRSs2Azn7XNnzNZgsVjCcEg9LjR2ej+fEyE1OtTiEeG2hTnIPdw8sQMlOFwqm
clw2Pe5Jf9muspX3IlaTbphht8EEz82AqwmeBPLJsMJqV2plwhKS1RfLlgllJGbvdHEf54kpAHNa
yHNr++s19i0jUiQMd2bhO6uW8VXzGEM/qz58r1DrO3Vlr3Amyn8SqDKuWTREe58ynlY2+51AC6ZF
xx2LMHSngxcV4D84Y/qKqEMBjbkHwui0CHVhqo+CoZBmjtr1cxurvLTkEyqMKuKVVkDnWPGH3pTq
iFeakzLEfZUaw0jPjT0pMlCkpidkuIZCxZuIFcfPqHK6ySzzoGSSmm/Az7TLaOHjmNlA1XGwu1Tk
+AlxMx0lrf00l+UvnP2cRL/tTwMC+vy1Wo3iVBA7iDAPUytMKAKkCaPvSVZPG3/T9PLxG3m7/nHr
Uu/Ide5SVkE76S12Y/makYLfCQZ+9FsnhvjgQbR6nAnpYUG4xU/VMjhpBoALsc9WLUy1s9WHU7YK
tcd+keq2GBDmSpQ70zns5kXQMbEp8ezfzjtg//Z4n9SAGK6g+XtEG1b8rXt57TgETkYKLJ12YbaC
ZJ0INhlYuOxaWIJV71OcskpO+2xJCg9Od9psNPo50RSyTBUK8HhSgZuBMZ0IISNI0KR1yC/LhyQC
D8J/EcC835M3YTZsDb9s/aikEIZypE29GA3U9hJHFX9IL4fwE3OaI+fkFzBp2U49WWyxirCKQyRM
5Q/SxBS6ou/dY/VPcv7uD5xj9bYbQcXcd9y/D/i69DIPmB+I1LTP8xd0ROwbZrFmhQI1rXotacEx
8D3eLR4luq5iFjMpdk0RWvC4BZgjpLvslPzxt5+xpA7tA843bTZA7l71HNjjKCP5Kl+olCjNPErB
Qigy04htuPrE1AXKcoY71OJovSu4JaKCB2pEebWNO3Ck0UyUzbPvUAgduy4v9VgShVxn59rpa5bE
uIgboXRih1JntGSBBlRGCY1c3nDNuUbkYf+I3DrzWkdx9puXObSn/l6GfJVHlN5xP/0gD76vmrtm
uaLE4rYOkNJc3P+GtuDbSCp9MqcQjuZxLtxhvO6MprjimT/NYQ58GdJePtXW0b3+qjylmNMyJIl6
PJHzHXQ9RxqPkwjdUU6nfetAtMbEYGWavm/1OkOLyi/S69HV+ZqhKeqttsEcg7RKQ/ISjBMQn+fq
z3mWRlU12AZoNMsciz7uHVFO4rUm1unovrf/aVRWrM0DwzCg1H+uL+9R9fedzaJekC5R3D83Bjaj
HsalIs+YVY2mkS5s0QUJaAYuExLRHQF9ErqOvbgJMDaIojMinS+h0LOlD3M9d/14DL1TN2uwXuVB
BRb+TucPsvIs/K8eIh191m9ljxt54Ib6juGbvK0hJVjzgqoOvwceIhyNbNEId0FVYjGvtCXH5O/T
HnPeIrvVTDtHGl1oMReOJLSM9ti23sFCUyrz7voUo/w5A89GPKPqiutH7tLQUc9OrZh1Rv2ABh0E
HIqXyYJriZ4ILtlFoqMwIwGPPMANpxdI0ho+Fie/ISPfRLgruJKVqZ500TsUph05fycdXSgJDMFV
JLRQkdUiE0N2lsq2sQ9R0ZJNlZVFFAMc5mvGR7IwNuXxQpSN19OdxnvG+sY/fGtViEK28MO2TNbX
UE20kdc9+u/wnECHlzv6K3faFFxPifcgcyN2BU8u/uKXOgMyaO4YBuPX0w19rDU2aUQJc7SOwj/X
41CwE9j+PsbTihwHFCeDFhF8W22nBbaEixsKBPy0XF9SUg4rmbLcasZAE1PVGZasaiU6M6W9b07U
neEY6P76kIdzb/YGes6j/G23d64YvMqD6ZC3TnON18J7Y2j5SyVPwg9tbA3xaXF3EyU1xXEMbioO
eusziZg12l/yBkWso1M4ZWoGArHBUplrarEkVCMVrK08NGzlAJPD6xdkmINRW5pxjoph9A/tVutR
O3yML3nz0Cqkww8M7L8NDvYm9z6maSYBZ5FN0436kqVHtcl+m0JfvkY0UjXdymeFmplE6hNW6KN+
0VTeklf1Oh26ElAlFoc6xUf60cgDaT1R2n/AoOYK0gIbXzCJbnVMYtsavtpv1xCopffWDuZQVCjR
bLlskQQtJ51Dg+IXm1w87kjD0f6mM9i8cF6vj1mWYcixeVdNH5OQZfYEpCbScLGNJdtAuqF+qhn0
fygOrlIpHlTgU/OaoyjtyEiYPJVgW1D+II9bnSeTffOIzHB7HPlZW5FjmOu6g3dVrevK2LqNOop4
zIrh9xwJ8X+CfW6cmr6Vg31ay/pmBVZNK6Srt4e2dCnbQmrwSdeFZe1cUNKDdmzTl11Ep0d3bzfj
bwc7mZV5KV8nkmRI2R7ZbAM8vjiGfgEGcAX0VZlLuR8gkb+b0gvlgxzqNUc9CZmI5L1cAMjuIBDB
7cYLzQEZ8Jb9+cM3pKmBMc3TxDdTzPE8nHZH7UKzc/JYTuOx2VRZgbl/zQb08Sgn+YaL5Cvyp8dv
iRfXCDBHgU4J2J6HVZZkW31JxPtE56HFAdY3EY1hcpxTt6xi8LLsWcAyBf/p+B/mcaCY/m+4RPdE
qwI5zJtmG76hqKmYCr7q/dTElBsZSk8AQ0n6k2KeKRZh4DsMqn443TdUds4LF25W+OByRgKo7NlL
OJS22Sn2V1oQMEMWVTSUYzqqk4fK0LR01A+MLpwoA/bUaPmnjxJyEQC2lMjsi2faM2MB6mJlGjPG
5hR4BWY44ugg+JrE8q+2SB663Es2+eDIzW71cDiD+K39gz8KBUPD4AxdinZXnJ2ZG31nm1LeMnqG
tXhjYjHFsOvo6H7swTrL+4psj5eaiIyLX8+FFIcSWdry4J46MIJJ8whHRkWmOIRTPBas1F2q//36
Crlp25b0bmNK7BG+iNIWzgxFfGBS94iWh+TLrYOGeI6DkXPS5QHiqbLHejee3uhPo47RfHRzDW4g
B24+j3Tv76W/D451/ZHU41lBtMplh7MQH1LZukjc+UrOqEh69pmtINwJi9GQnVvfTanPdBnzoHEW
b8RTKvX2dOAK4ypi7+myfOPVek1eRQkHOOHzcVFjmW1R3tTPG4RIUJHBaq4e4AI8Ve7oYU4a3fqr
mtwA8zaxXAkDw9wDWuEFksi0kZmpm50cZfCa+qSyJYw9076E660dBzfUi2jLjU514919FOMVOnw2
nB/0F0iyZ+K3I/6VFcn3C4sIvvuL1+NA0Br5hXY5ndE5L8DeA7nJ18FmIbCA2J1Ilg9t+JONznTN
3pnltGUvmcru8E5p2zgILLfwOIp/JVrYPcBPooWNjObjbRCaLOahY/Trzp0i5DX9SVlHkaD18Jh6
dogCvbLx9P2X2Vw0qVp4t5A5gVW3xq/02CkLt3Vlbla0+6hLSDKFtrNhYAVmJkFg+d+tXkXGk1le
3l+ehLgherS5UkN27VGXVS8kbzzmu3TfHwlA2z2DicVJJaYyvPExK2bzPUFJnR5XVENau5AUkRxx
+Uc9/gbOZFJHK2PNxy74EgYbksPAozRXnUrKyCmw3AcoD3oiPa/6XuH9wev2bQrHhxGz6bWDdSfA
bf9J59Ly+ItdsEb30ahNOTMF584mm0pEU+XpChqo2ELn79NcPtdt7MNYq0xAfQbzhWo7d/nYxcHL
aB53x9iGGtlsdirJdp3Dc8/agJInzRcCbvJGlxV9hMU/ro7cpy0hVLUnOPgNFG64w25C2KIYYRuY
6Hu2t5WDjpliqzvOMnx2Q0Me0j4REyIFp6ECPsSKNlKfgP7sMVkD4vS58MAZ3MI2Qxdufo1WGxTG
aGwy9RIaqamQMw8ImTdc/aF4pBt/jSv0DhNjyygbxi1YpkqbVEQqy/7ZGvhGBb5IoUqC3bGtvVwJ
xAIVvotHZnFHtWXFGv0f3Kxj4esQLy6JzuMUrCsPwiJt6lw7eZ8qEksK4o9mccMa+Tp2xM+7SOJK
4/WXKAKjDCGDCw9zd/p6FndQ11Ut01AAfuJpl+pLyolo+ZrL/bwc8/be5JIsc9DCTXDa6bk5nfPC
MsVhUoYmkPhBfm5+51RYbMocbzIGUTvpp791WCqUX9Lx3Z4ZJi+XceFwUN0zhr7hIbjgZD+aaJU9
yc/biObSKaW4usvLz4McmUyn9jPiELFpLc2a5Dd5BFeR9fDjO15dxHiessxdpUeOOJXWpQL+DW4A
GyW2J+CKmJuFif1Ge1JivI208hns/J4Sjwx/ohu6D466PvBvqDi73uJZDMocKHyIdlpLv13fv75I
l8QNwq6Ax4OY6GT/rkTvR/o3RCvtw0QwFReSOaP46/ROhQ+z9BLcK05IeQBcyLtL3Xb6ggpUJi4j
22dXJYwLhZQb/PUr/g/bgsGyg/UAoIICDaL5LuaD6YBXy3W3PECSJZxb144wxHvmDaj8l03ejAvw
MYmcj/b9qNQTw2mfxoMp3BgDXercdq3Q/mH+TH5H189gdslYHm+bn3ObjgdVXNECZ3BikJTisniZ
K5QAz9fcpYkLHuKGFgN9RdEL5c2zMFLDm2oP23Vm/763WX9MagVAYwC5uxV8bv3fVNFJ35XvpcNY
9kidNmXWYU88zFgxdwOhH3ev3eyB5tcGRnMTaNU5X9j+atErnyztj0ln72XNJeYguDVzPCRYXHLu
oXfZ2LUjY3SQ0M1KPoPnOtuG1Yw0XSQGf3HC3J074PesEp9MwBI5jmj1AzuGdrS0Pui1qU4hbXSL
MDXHpVqsAjLmxC6j0zVPi9aEsGNaT7YJLcPdKf6XOLsw3iIwpmHQbqEubrrvsXl+0Tzw40Cj8AnQ
4zY43zAereK3PlEo7L5kMG4lN7bleFMEblVmDd84wa7idd2Y9nyWRQsipdlX8y3n6dppy4NcJrum
2etjQjvyz7bzA1W+aNwhvzo6+Ea+DdsPUBZe0s6vFTX0K2QmKL5fOgfrf5rY9ThXtTi0nYa+YKy+
a5YaLbgvi++0V7oao0QfqA6c9n32v4oRbBAf9086kM5ofI5Mlx5mVOl5QzPI+UvM/APhXf7DqLXQ
MgC/MCAt/PdA52ZMIUO4AB8LglHA3lmNCnkWO/PBMsPSNLNyX8M92T1lnvZh/w10A3oQaaejKkO+
B4BQ3Dcal8uo0pBEo84MumfY2Ck00BxMtZpTK/c4YGNvqEr+I/N37+EUhgE+pnlhYUq4jP6I/NnU
qjnhHimqADnubxt79HsnTFVb/H14JU9WgxX0hyhXYMflU1JJd87Wx3h/Nzkck+AP4+G5tCUhOgbE
9DmvaYLLl14RlIwM+EC58V0FahkLNeUxlG3UnUKYoxppczTsCufKVem/FyR+BJ0ly6ybPsyj8Vss
Jr6RLJ073+Dh7QX3v3W3RBrgFuoTZ5eoM6SBARMm31q9fmBgSZCpBNJb++xwAjbuNvD0dWVPR6f+
PrrkVcx5oEvniN7+LPeTI7TYUVg12fgS3obapE4TMblmv+jBJf2J1BCGLG7Hf0mjtslyZqR0RMxm
SWxkdUp7olY8pZm8z7iFA1qJTUpKwwUNV8C0Bbr/UFlEZd29R9VZKjp8IvqtQRMQDkwq4abIRj8e
fiuho5Tfq/Fs7nkXsZrZzdOqvl5OHwUT+YVimtAJ2wWBiuXwelzIN0vtSURVHD83L/77ubLu8nsI
2MzDdjwmgnb4JFmpLn3WCxJtKiUfXuuJa4qrIK6hRtsrUEWQbmIJhYPhuGo8WyMWFSyaF5C0Ckau
rO1Yv/8hINQf9GDBfixjeBj4fY+KaOAkHOcTx+GwsKKYhOYcKcFKp5k1iiVEwY/yleD6X7Kjm6ih
M9/U3y+upNv87bx3aluj7A8vElqbCiPqwNrhVvPqKMG/u0F7Xp1FpTFaimoJ3X8uNPz/YUpuTCDu
KqUfvZBmdvplb490krKj/KQxbJATELZK76mXAVtjPIK3HRvdRNW8erHaTcSDzZjSN9nQW7q1VvG+
UwyNjG4iVu0aAMjgpDtRNeB87vtJeOa99Nuw+FEa680CpvAl9x27rqT44DpS1ZgZpEJ0qcWVkDwd
DFuotnIBP7bWKzRjp7fbawB1gmjiJGxVzkRXGtHFIPT52Z8SNUcY7LGYiB8SOPDkTFNbQFnCLMcg
y9/VkT4D+DgaLhtb+KUnLg1Ef6T80ZoEgGP3E9hr2hn/9pRB7mpoVWJc0MIAJcbPV9cMcGYTHgVF
tsmY+tfq37sfTSKlMB5iHokoROVQba6LRoyNWgDsZ8G6dfbNujmjIj7eJknGIBJkgQmEa3DBuT4g
mER+8G5nkWzZU/YSLY7sEsmGe2/Pe/bzMbCl6T60FtuQK3KSkkMWc3k2RUH1p/LSFLRXcxs6/2pq
h7kP05RpnUpv8eO4OW2xU9GUwiN/7ATxGEpdjSSUh5EnRkOGz24/98L6ucO3NuWPSUS5oZtguv2U
UH3wSIj3RSUU+X86GymJlDK2kB8CZOMWVUsjz4tvRYApGxNpgnq3o5IJoBeOOwiNqPbq1n91NKAs
1zuIdJM4dKZWlc/1Qp/8ldd20Yj2juilP6CJzJTLym76LKcY6euWgxyFlvtmzLJfInyMDABo7+ir
vKWRlPAyUFvw+ksd5YJPGI0Y7nn8xmZTi4M0UrYhNZzkhrx0pY1NUZefN1jMTXQ2qZikoWN7gozQ
7p6IHucnGDgW5BGYSrTo+kgqzM9c3PhUmYEjULVWp0rP9gxhl2L0yoQU+b1Ou5F6xhooYeFUf5UO
oTfNM4VgVxKtjrfUpzhDQ9EEBhg9+Yo/U+epXTpsZ1plNHgvFdpxGVUFixsJapQrxxyEnGS0X32j
YBTkwGX1/1PyM+9NSktONup2L/jk407ib1C/NHIl9tDA8XvNTyAHwMeHpwhTl/UFJ3d5chgkFrv9
8V0bkLGgFCiC1nMRDAyTcynhSNLQV/hUyTpFP92gVQlMPOqZDVAU7DOrutg2ej6S6OS/CSHglon4
hwC0ELUuW9lHsLaLjUscgb6DmbA1V9LFzOmvxv4NuKOLWKNsX7Xou7ItGo594Mna1FXVCCPTEOo9
8GMq63D8c9g5NsckLQHGnUEi/CQdmC9XOiwVZIeIOEsum3bprvZ2pNUI7fAZgGYDZOmhlS8FfBJB
FcTBBM3c7bURaO3oKY7YR7c8m2N8p5xzp2HmsyvBli9atCDgLKT/W+Ixtq+qgHZLndvlcJ7UpaVi
iggRrJyfDVJI65XccIvZCeAG1w+HktAIX9qn/C3x25DZWFxJmwpYYzoyyMExb+xhjFet8A3l15ef
Bj5c0sLBCYDbredLf4IFN9HAp9lCLSMytWRlEHso0cc4w5WqTf4mWcxUa7b18R4lyeSzNtq0RKQ4
5A+1ytHidBIcF/FCJP7hGs9KBg3ByKY4glatLWwKod880YGv2wU1nEYkZRumQuefbFhxZ+5QG9He
5UtLKSPlqz12oS0dI0tqqWkXuQt2NYfynC4u37yh2s+k1TOLgJJGfnKSmT0s5niM3o3jkvx+XXTt
KpDYd9V9fgcroVoanepzVN9SpEx7BfI+aYFwFttaEQ40B1lTFIeASgFRf7zivIveEf7tKd6ydI2C
CMnsK3LIrNhe1tgulW1ENgC8xeBTXvMymJ2pPgjIsilgEOAqMOGliNANKGsgghmRtkfnOioZIlLm
t83eE+Ck1dD2wud/bPvv5Ch1fuznEK1R5ggRAeW5sDEBcYWfm3OPbPTXFp012ucjzgVzHe5ixnhZ
7uYAytqItBR4Olw+K+BCvIGjJYTNoizOvqRqz6+ZcJ2nGp1qtCB7xmBr/LXiRgmjyhz4pCtDd2dd
+zHL9yrG0q3t8V54CDE417ruCrhtRV8hvzu3UWHsCvaahacsVhtC1BYxNVUCWuYXwPtsbh/VCLWc
j8+RPUV00CLdYxrJwapwArUYxdsl5IHqG6Fx2nunIJTWIJQ9sxO4KIYJ7RrRHdIs8FIu1ftpjS/v
tCmZD2bxJh0SY3y78hsMUf4tN+9tYcJTdwHlVeUJl0tDPME8yy8sp6NsM8xci49MRUCU7Dw0xzau
6i+Y3VBY6mFD37AH1+6TtCWiXlO7rpOZl456UUWJ1JIy8hHswa/0pai9hE8bdnC2bpyJkpqnQGaF
FvKvyTIm/8BHqTQlTSqwc+Yewqlxl+NZkoHDgQHkM+B/r6v0yBAS5sRnFMKXvCXFdXBL/5M02NOw
6fq9Fu/ngKmWeNIQigDl+CeBc0zeWwrsyO0YMfChcR4RjJIBHZjHRlE/km6lpr/7/my9fSzKWBkq
MX5HViamv33VjCVFKZrKwT54Fvg1AJxPcu3CCrkAVrlkFKqKbWO4oDrhm370WRvCjLh3cweaKoe8
t3mNcWQ3xGfM26UZiwAbst1elsioGE75a51eVcxE851TB2ubK83e6v+ZIap+HQR/Re3daQ1LwbuJ
UOHId8PgVkJuLp0H3MU1QF0VL4Qid9KoWQOzjX/EvuEgZnSc48sxe8gyFOGWC3+c5VR7gEfW4Yu8
RGqUcQU0hyjQH9vjET3ktZ5s7GvakwAAJmo5w9Jmxatidb+jYOQciuiEvQ+1LM/m2jzuKXltJef5
7CqhU3tJUCnXdSyRJ2LLVvqsB6rjAuPcsU4MgFJSLfD7QDu1Iga0PsOFixQnehlEPu1VSxcw0Efu
Ib50iXW+37ECPaapRbTwgFzOKcw3oX2sEQbLzZBcVDMgjorUjQlrsyUlYhs7e8H5Ma8l38z+2Aow
l1i7LOklCPtJ4YhpRpLfDofQcDguYRvGDYwCi6PAVdds5ygybl5l7bSHFlpyE6MKu8fVDZJihP8r
q4CeWIeejZBfdWTB90A4lDLAQXnJrsVMd9CPpp9WTm1iEK0/NSeI4GoqxtYGd5hpcaKMEFjwrPKH
UnunsHjqbGnTHL0GxTyH4sdzoLexNA19mkpwDyyncIM4aaWyWJGqITwlBfABwqnXoS/4uns4KBtF
x+zkZwL+2Frfrht1rQkqeJju1KYp/L4gJgZFoWNI6tKooyBRHfs1oBKO1JstoD6UD+xIDRRHhzJ8
ujxk9G0fFvUYtOAk14aqt89P3UdxDtu5R+1IwEuwBvLXLbnXpO614dCXb1EC7ETi897lafxoBs57
PpKoNtodfAG37zSV7VTvFia9JIscSwtU37b8icUWS1cGgGr6t31G7UNYixOexx+43pUUz1d9M797
SItspWWDth+J7hIgUVrS5GkTE9ROgYw/h2txG4pKjYKx5yC6u4zo8SDb8rMHc9xFw7/Y/UPjPkID
0nldsoU0P/ZxfL+rALWVuoD6jDqNOMnVVJfGw5O7RC+vyflp1q9P/pr4pTSPHbL3mTWlHXj6cjWr
YOs37mY4jIQK98dt9cCSdAdzcQ7ZBPvLKAB9ZyHVcf4vJhzSVV6wEpG4aSW83v07NOUyNGytOMzI
Hp0z03aU3WGPf0tZFCeJ25Qtwd/HPFp3A0aEMTSDUKm8R6Y9IsC6vq2MmR80Y80C1s/a1Pt6O2or
YQMgOqjfO9LjrTODfJ66SWmNCyejEpNVR1sk+Jxsg2VxEq/VOU20i2lSTfdoB49FdgSAU1nyGR8q
QP+5GgchL5PNCsMEcspZ5812Rl2ZVsNCxC4jBa2iOLTL2s324hZlajuRQxjNwKG93liQRLWzuhPi
P6ipRkJZ3Z89FN+h2INTRskoeLGffYHIHX6Gsjov+yI0xRXBxiZDEDSW16RrjAH/Hhc1pFRbwuxp
uxvR+YsWs+ks2pACS01HE45F4u/KXn6IN/pER6iHRGmd3F9WWRYxlRe5E75CVG+nEi6Ud1YLOu9S
H8gnWtfy4sz0J/I43OLPCeGFXf/HYSNAPYc9hxP0VxhqdKrseXmFkvd6ZiTvGUdhmghMYEiMqJH7
xNIrp+wgB/WDMfbEkuuYOa62+qAsyTcraXbbTxIKC/o2pNqal4OXnjRwo9YGtmxLUif0XAb1W0OZ
NJlRlBsmYPBCYyrDv2RBhMU9yS6kFMKGuurIAxGGhQpsz9lRfb/Zgp/20A1+A2bFlclcM4zUtXy/
B0yksCdscUjVWGjbw6JawILue7H19hGHRghnwLi7EZAg/rI59hBPOt+zi2gtXPPnnpaG0e699Od1
12kEI+Y0NjHhzQXndjK6N5uhLamz+OfuHsm4UDrj5sBk+9O/9OxyXoTOpn1IBQ09uvBs9Sm2VfQy
rOsCm8DN5oLUqtjTOgn5Es+pf3ENIAYZ2CzJT2xMr745CETGUGyHz/x4Gcfwwih0vowuLkc8xLqC
JocTKdw1O9Zk0sZaV8fal7dQoks0SxMTytojjhDDDlGZ23yQnk0Ir92cr5KNr6BpvZ1CNwWM1+QD
klDYhCV3ukCnwDiBSH/F3kUKdsW+uumtpH8SsNHAyp9eRAm+Go5ohRVlSV5QO2qHP1Y5dpcDXBPe
Se138YQ/exHKAzD/QxtYB3VWu/OsltgP8QlV5fwGrKZT1UPEl6edyRkzJywqHMB1eql0oMJB8VH0
6zGoPxxPzDDkYQXBpG9UcwRgZM9U4+EUFSWXVNovyMa2IWfP6vY7Qp3RpnJbwSQb7wsCN/2wQXfw
gFLBPUDPxp033x8OQ1Pz3XVmMJavFqPX/iMGr28iOVG9bVLhxROq1zA20ezaCNBx0JE5vbiprQGi
2Q7cQYDWCRZvkP6/l64AupLubjSsicWHNpksjWBw13Tuy5dvbEiZ/Xqz3/9vwb6bPDiecypDqYhM
l25pQTAq9q9UULbXgrLWGKjfy2UkMij1tMsOuqM8ARimTnPMVryPSsEEfaxC4ZdeB8Ey81a3vBlF
T3mjDpAuU3BUPpiQBjmVK2/FjBuppAD0pGJ3xFJKu+TxCKi4ypThR3GMclvN53jA2c/DReeQ8Gic
ifkfrvZG4VCPrM7/bE8BdJNTgbPRMPYiDY1H+YovGJH4MOiBj9ygyGRvlIhlp2mQAv17WcSQYKNr
rULvhKHUT9FR8gFjrYwidNmbCbLxlogiQsmw5+85gc6hBFaj/LjFlmLJ2/nMKpkyrA+58/k/nFjC
vFlLl78gC3JFL6cUrB7hH7NGcYQ4VHizA04JFlgE8Et8JlmPC/YlC65pE6pY5ud/oPSYBMBGXJJQ
FlG/fQumbCQ6qbuadhatMGBbI+Hm4BDyXFCj3PvwXKFMuXJc19u1euuLeMprfIM0jsWUnOeh2z4d
wIM75uXqH5Ch/VfYpIewzzSnlA5ceK1/2c8Vllcq74vKeLKnhVkJSQT+0Tx0gbwDMteC3AgTsOZz
l7e+06qHes4hhVLdd7JbNzeDUM+mn1kJpugYh2TLB/3kDVqznNTzDeI6v3zrHRjQX/5qNQqlnCjt
ACLd838LuLyJ0surf5vyUBucEXOBumcVQPtAeaKEC/6Z7/9HX4ZQiAkVRzo1bJeNc0UgooZPm5BW
fCXJ1GUJpekRG1gIFXZjpK1OEzn5pxPii2SG78J7hP3CLkbmU/ZTmWfsBQqwUrXEE/cnhN9bv1ZO
19SwukoHnzYwusnBQbx6wDGbhCZ1EkZ7JDrdNRmujgzmJIw9d2nWXSwnCTmcjFHHvzsclhgX5RBH
L2ZQqwI94ia7CNu+IR3lZ9yJ9uNCkfahdZy7JKJbimLFKDE3YPXz4ZN7+kkKEYBU8xicOYH9Qmbz
tpeklsuO80DS88k3PZyDzistHw1JzM6A86nDv/P4xpfmCjvTL3cuVncIokoqQrBhP0UQ4XSXM2aP
kZmTM93tU7fb00ffDtvYxl7FrwtGkAzwFFB44rPHVgXARhTVwld7B2jhm61d9GvgJ6mfSz33lpSl
zpUuL69dL1/tGRfj170UoWPQTgOkfij3p/mMaZWw2NicbLKhDzI4l+8XwPPTG5SWgiTY7u8nprlF
aIXfOVKCLda7SzMsQzE8CFMfBX/E9qrbegjs3SzIz3UfL+JYsfs9VyY8B/R2qOOkVQvuEci7M9g1
oRr65UJpDGuBlBgfz2cETfm0r6VsCTJWZCo1dJ7xDnKAZcfQQA+eEXfE82s5LXpUuHacNy7eLq9N
5tzMaGqL1bARyafRkOWjltcvi8mxBRiyPY85k89T3hBV0IDzHlIWBujwMY2xl6c8ZDRwkykzJK+f
JGfdTIItohOJ+xhEtBkUEo8KkmLAYIiapF3GMhcrq3PkpEvEh3LLzSv1EPTmQGL/dVPCB0BX9rsU
EUmTRokQQRQE9rfv4P1Uqarxm+9V3aTjxpmdcHMP+FtWoKdqevjqHNJ1da+1UM0xh7vAWFDO5Pqp
QmGg4htDblFDaHY581iWu3w4Mf09MiZo8/Oi9uuDCqn3vUWccZAS3en0u4qBwXMIWU/t+CDyD8SG
I6T6pptgyhwwoFVpB+5EfpkaqgNcjR/Fdy1hgIcH74YDwH3x3P30j0ATry7A2AUv8M3og7SCbPFN
TlXTeQgkWu7i2U1EWHMmRCqqHkiF6DP8aRCIFM/LMC69kC1SdlRErln1i4bXn2foP33DUZPSbUZV
ZzjLzoFQ7jaGJbGOR61h8TSQgvEaeOdCIlOLXCsLjZXMYAIg1Xffi3q7l/2fpeUCHuonREu0OK7C
Xf3Q2qKTqGn3sCTekiXBAg6mHaAaBlw87LHneqREftOKFOHSc6HBC+PemRAgTAcJvgJQdKrXMkSL
ujyuwKqu0cQiW9UYSszX/WlWISuH/AOScqlOV1eDUdcqdaLx8eeXZkwP/E+B3uY/vTKey0sstW4m
tPUxPVb0lvGWiU4/XY8h75syEMzb1PFtsXDNMlT9+ZZNOWw+CRHoNYJJgOSyBJEN3fVIud1daJ63
zBk2pp/kYJsdqEDOB9Uz0pplEcszbNdQjEjG2W9Yj4gfuFnCN27qxqRlvBiWDk2hkILAkBdWrCum
xAiGjWVTrsGe/uoHNIZ1r0q6ra0rXdyId4mxx6WYSf+dyzHShOh7G7w1UHsdFl+n5uY5ZjlTn/QG
7glk8eanAV9QYUY0SttPa99gAiHCyrOTMs8nhhbKJ5fgq2hivT3wRyUZm/oq/kRnS7EKT1vPCYUp
nLhNDvg95QL9zwliA+WTkaeMCY1DlNZiCZluhpfz5X3EVdUsNQe5/oTZu8Uq/5DXbqVzJZoftH/z
0n7tkRtL5zMvbrj+6IC4k+YOUL6adaR5pBL4ZUE9imOr6pZN6Ar8CAUrTnl2TK6FCh3FLTDOfNDZ
+T1nmgBOWfbIm/EHFHQaQeiryHzpJkSKugCYE7N8sVDbBa2fVxMzmOBcz8TuWhGqcxo6dOxAih6/
Bo2E6uSR9MWHh5uiaOb1IRn7rkVgNPk7oCCJq0JD/UcFy48/0wTGTkwPDKMRik7vA/rA2MQTfLmi
zD2KamnUvbm2++EF1Fj9pIQlvqp4mlSqpR7PRZCuY4DsT37UDpyTShRQNKK0eGFlYQr3U1IKdZdG
DbKcaMeGq+cXMprbor8cx7Bfrg8YQmgFtnq3w+Vr7y4jZOTi036U3PyN43P4ymXJu9VfAGsA1e9I
B3NRob8pWOERJS5+KV6NVh1v+XpVXQae+rVB1/Fnm3uzgWbmdnrvMrxp5V05F8XoHc/k2o2X+60/
5VwXGrv6BStUrey+gfPLHzFKbhVDseJMkTwa97k3RSGz4QnsFox7xhVnqAzF+qr/2Ws/l9JIGX6F
mvh9l/0QIyVLfItJV4JJi3SsyTVnI9xqz9SNHS30EnwJCdEr8xB0SNDLcz2kn/qfwftOsLZbOli5
SqwH08aMcaBrii1XkguVpogjwZ79r/SuhbuMgkrIJlgkYoEOF49/rCQY9AhgW0zxWQaNbXEFUv2i
9VsdSKfD9U4742YV5ACFxWDGFUpxkTUGgwqVnJisDdRu3JUc1x3BZUSE1xwpFJN4jJIevQSXmy0L
xHYWBjfA7vIYpOvMr3jcPQR6BIW80cttuLgBLtPSOwyIsjJwDNRWoSUnq6xhefPIqKnBASlEy7gM
vK2UIY5LKdMeU5zIjlan8OuH1e1wPOjfHe/KLDskzw3uLeek1gNflqpAKKCR1ZT2isuml634aiCC
3tnIBRfUTAhcsLqEQR3xMgyYizXwqd70vXsxvczg24MlhsPnud+tFzAH3kEwnozeqzXU3T0Gfcdx
oIHWRj7jBcwNZcktP30WY1fslTpzfjgp/51N6tpxe7wzavVpD71Tvmst44Wn1b7jNBAeBbHWcMyo
EMmK2/78nAXsIXLlInJsyXP0bkeB0PZ1Qq70spgoYg4OntJbVDum3H38vx7Vd1UsqX7UqJfFjS5Z
reFVfnW5O/v5S0eWtpcDnB3I/dkqUCk0Yhy+WItANN+2stIReOhZyDwN5x19PT1ErLJ5+Kl2Zf7X
gusxJd4ld9sOD4uTPpeg88n0C1zCtj3GKa/CyIyTnVL+70Wh+5wOFeEOLii8e4LSyaBmfnPR6LJq
zFgGvY7K2cWjtVYOhijqzodgqSFHEFVfSX+lPYT2amB4SveB8xUOBACVgMq04oZzXcSBZnHdj8rA
QbaIfhUnFMLCLoDVHfnQOd9V2WCYLHyHptTFCPxnkafpExEU1NErpO7QXMOXdEOhgT2R4EIjyzIj
c+aTGsUgF5phPrCIX641B3LaM6d8xMeRsVl9oVjrF6OW8Pv/N4i9NoZJPCuVPzZYHgrT3CLXQQf2
1LgogLSjjPBwjJSrpv4CiJkysSudNVCaHoPyXKC2mEEa/Ks1pbgLQRRNuFaAISEns6GmsLg/3GrR
cHPVfKgt3e3sZ3trRKAww4SPgadQUQp6CWeUh1/pOd3rbBG0vBnLPRi/6pBuYcjjWjg83osn2Q6E
4ZD3svQ7euEH3N/sAk7fBu41WQ5YPk9l1bfKtcMRH86a6F21ueGypiCdotrWEIubp/2WqfmKuuxl
fclDyim0CbCkiMx/implgfvzEu0i1TNrc+8D7LwODMa1sN+gj8eJg9/gXaQTBbK62ZMMlPekkZ/R
Dm0wE4QJw644mFRpb7tCXwW93vYdYjsOLjFEltN9YWEJybpsM92Fr00trr4WFWCR6gnODpo8cMNr
SWhoJuHYtSokoltjEszINocojBM7qDWNT/vW05rdTL2P6l0/2cwdnw6oyJcP/hlvvT97Luq/K/Rs
2drDEbB3yluV2ERb+/RNO8pnNngi8cLzvqp1d6JcbNs5Fv7dLGxGVC9esbwOZxqBT923DpovZeEQ
57Grn0FNFE0BHmld3oECLTB2oHfJ76pOpRCKe4RHpq7o3jF+VuF4Vb+8NpG7NtggJZNNCqm+lmAu
eqwd+znTNQ0b2KTJRbLBzpr0BGb3c59f/vLkqeDpKRD0Umz/qTwJQgfHXwM9x80Xozy8FSUaWp2G
ICgqJPgDTgTVGSES8CmPYxDt4vH/I7YTYgBAqAw4oO1S8a5MlfuWDvJmzq7PS3jNWmdYGKOx02fM
h9kxSrEA8hkKe7frIYl5JRDKNf4b0Nzfkxap3+mzCoWkztdBzwTPl1YPEnFiQPLmHiCyu0NMPVpk
NQi/AaUXilrBZo8ylTo2+ah5JIzjMlPGEaE8EuVHmPAuiAhX2wzQuYUZAlAMMdYXCUMAGE1P92ig
XHDzLpMzOaRiY5C91vu6p359DznHB/fXmivEiU/jtNYR9335HJZHll5EV4k7mtKwGodiLWbQZ2SQ
xLyp/wwVG7xUUnZmNOnweMMO75pc4gNLe8W8P6iLzslMhWFW9kxOD1UMooZtWVbEg5c6mLbDMgka
mc1bbUNZzdfpTUPzNhk6yeKEJU0L42+7ne9s1C4+j/vCXHScRo2Yo0ZiVun3EAmC9w9W0WfU++wm
vUHWbCKYmONGfTBmgtlmAiahTo3LJP7Ya8Fss2np7ji1lb+tacBYwmzHK4zZu9FdE0aKCAZDmxuI
m+QaG0bkbXdYgU5Oqud3BRTKFxljyMDP8iW779Vryt40cB20f+OTQbp+5uI85VRD+lVBKVGsV7dO
O9iG3qRDQHRh4A0RmF7KWSZuhjec0VosmU3Kw5smgyYJuGhTkFpjc26tClxqOILgRI655vY3/H6c
g26ZBQDs97gtULl8aYez2fPoXbQRzPkf9emKYRmkOUmFZh1Up5+j5fRe/Fa5Fq7GJuWtNZh4E5ET
LPo6DarCKlr0tTzrKhhEOZmHSGJxW8SwhOPQKmh1bMDlMDjiBLi/r6q92JiJGaItvgQ/xy/oCUi2
JPP0F6l69a5ClU//qARqKV6hsc2PvICuSBx2fYx331/Qd3kIGcc47aDuCFhKeqj/+vaKJwjlILMF
eOjiZWnUybbOK2dMvF4K1/njGGIfUKZVS5IgZdKAS6Gs2abpLImOEHZCW2Xd7LD+l9yzNRCDb3Mz
GvWmJhkBESS6A+JqMFMhnmwXO44zMB0gNLzqM/zGPbTlMTvlE8isbGhUMZHCjBCJ6pqBBVKv/BRP
NtU1FPML+emPv/5tE3Mwpj+irTtZB9vu0aWPdpNBQ314Rp4dO4PJYuc6ncKuVyiK3jR28q6/7f00
bzGpLPXd6qYEVvrZ8F25KAeqZuvixpgtsaNUL5kZ5njVhd/b4q/HkFXmvBu8eAQ0Uz4CZ6Owi4Fx
gms5sfdNuciCOsIN2YlMX6X+vKgRYQvLAXCZIaGPveEIheMAHWYtAaS3VQr6jYCVr79ZPFUbjpNx
divGZfAtev/a2uPJCt9/yu68CG6lsP2LaBTDoWWG8F1k+ntiI2wdXNUNCgv2Cr+GLO8IhKfa2lWD
4HY6jNlqOY4ExpAC/0toJpO8zgYfhwA/G5ZOdM/PqlgriRtBW2CNEN6ADp23gQkGHy6tUMF1SsDi
pkSS9uXAIBjVjvP9ZV9PrwWGF+RUYO5bExMKqAi3+Z+/QDw4tO/sqwneA+3x3vYk99EXkkoV0stA
CE1IoAUGPoMz0VGA3se/z72SR2yr9xW5Q//XbKmddXgNDAd2CT/kSdLFKfGx4d3ay8/hxCoMVha0
+sE6lCLi/c1dadyiBdxS1EstUpUN+oTGpagV4UPYu5vWIh9pYi4Cc8b2gwpQVgNfYEuyBFKtmO9E
zh66mEvO9D7+AeY9mSy7QvnpAQkMUrWvrSQlTId0Mof+s8DCJOJSh4bWvZ5NIdmX4xEgD1dR/GL7
ATR9aNMa9cxgzDEuz1oGukzI1Cn1HrV3I8ZV92j1YuX4MV7J/XOifAx3gf+rMiJ+Vwj38yncX1es
GPPBIHhgIcep80H6EIjCSOyYNorQw/tvYW4lntg5yI8OwOd6DNe42QAj2XTXTCF2Obl38dWKojtU
d+FMMnhoyaELOo0WMec92oVuFiMODesTBsGEfdrgYddHhsX3uNIerY6aP0C5W7hxLA3i1Zoh+zFx
LItObN5KYxj3CvPK92m5qfvp7SQl0s8nSWkrwFbmBoSj0QRGKD0X2B0dwWcyHKy37zQYoXA6LE9h
lfEFexK9v52+tqDMIb0sS86KklO3v4vug7lJdIdwfoIw0z0mQXntRX/wqtBJWaRNBmdcqlHJzV3f
ERXu6KqP3DfeGOLCtFt/GyfLQ1CrJF1rfbYdOd7XstXHI0eWcJGvKRk292wfAA52o4gIxmQOuKCb
k7f8px/KD5a0r+i4mwAaP/+KNTyZXfQeaFliHj/mG60wR7geyJHmo/tyL9O/u2nmykONXcu08EId
bpf2McxpKck67hHbLhNNtkjbVv3dqDTTlKXVP0e4PKuBpBTuyTvL/PK7qrLz3P0PJteKcqNkvjXr
76umWUkY1W96JqZ+FtUiEtGfjdINdd7onhEySJQsSWIHRcd5DMJ3R53BfwOyGf1qh5akpZGMhLuw
20cDDXvOJfb6GwrOJF7OW6IFBLnfm0O4jZ1/IVyRzAuBN8zjDNFQ28j+/kKM1bQh0Dz9Xq+VXR/L
ZSYw51Gf7Mdvu0RDoGEoEeCFub44Q5+tlFfu7HTTvc9Ib16r3udMVbHvXn58L7l1XNWj/GDYxDN9
iOHK/waMeh9Bubx5Ou3zSKxtN+TJdSc/Q+TAUE8v4GOhER8CtaHmReOGpiO41z27R7KvSJp2RW9l
hDRDennPOb9G4pg/GBc7ifvJ4eDnSL+RT/NuGz1/MKghXs6QnDscOwcY5DBCyLgt6T1v9hkQcrQj
LUaNoM/bnAwdbO7Tku4oPR1sHZ08NRXJLXyGDPiNlrH+cjG/JmX5DEk38XMFbEjMrOV7us3l8n8s
mg7/cjU7lCicgasRnXebL7NsUvSeeM7YuDNUxj74c0wCLItrT8IPF83QflEFu6lBmMcKbn58p0dU
oU0Uor4exEbrGZdVUkH3OErWmtI/nhTdIvqdPFAdBncjrQtDL4Y2fXYavDrx3y08lk3FaGtgRNNH
hrXOkY2BJZ9/NZyrq8IBss6kXjljCZSBALIeaFi/iyQ2Lh2Tq7RFB/tMesvZEwXxS50Id5dOAZsD
9FCH6s3XCllx3cHfWXQfqlH02R1yRaV446Ld6tl4Yt2fvZAIZSQHwxOA4ZH+IjQCRsnn31deFZxd
5kxIHRTJ9mTC0AerWLWpU/PgptlHkXQ4ejJsre2sEc5bzIkm9cmN1PjjQPwC9iQXuWERyb/K72VY
3GqzlojH2FjWnIKsjTWI7x7eDrKx4L1iDNY/6czJ7Dn75MdUyZ7xDnH//iPuLseavwWNrVzeZX1M
xBhM+a/sfHdA3fvuFyEw5BoKV8yNPH3Zu4sYfv5VA6Ap+UN3qvLpSsb3IL7w76qqus5VqX9mgJsv
F7xUyULGmDbkRZAGSZ5srbHog71VJhLoniuK1VjW6cczRZxWPVmhvWZ7xMqLzr6pONUPhPv6H+RC
8ZObWdv9rZMAx7VtWYdinrIqDW50BmQoke2pA46v5qcI6GYhRmh4H2vlI3SZRgR0CMwYoE/j4VZI
8uZuIqWsKK1CnkFVUp2ePQpRVC6lsu13tfyrZpZGJkkPhn8Tn+xM2ohSm6KWIXlINA4qocCRcpRE
QwmmaDLOroCFVc9fVQekCxAvGsMwYdo3K/tUFwCyPFvRjTV7asZhWyWhBoJazooEfeaPT2AZcmtH
LwmtJvptTMwXzUoAaTxlECF9xGYn3q04lm4wHmQ9zJljcHRsTAHIRjTnY5NdhpRKlujeu8AP24/K
uvaeUkicibQkeWxu/v5brHRBHw7Nfn1jxLdBwpnUoB1a/Gcf3urq7MwL+0E1UiuZGwjS1Vss4Snm
V8IRYZT9J+eLieNSKhOhOA6a2xEgNj0JC6JDA9t7Oee+Qwr0ROVo36dpQHF6Yc340inobWyN3EfW
sbcu9zuq6I0vRynAkmke9HE0b48zsmvaXMG5Hmsn1Ux1jjnrWC9xeyhsja6Hn6zdmriIIK4F6s/7
FF2dxvNZpIJeah3P3vvUNRPFFPjQEKFwWDTM4onHRZm62+E87QoCM/8f5tweXpryA+go0dAGThL4
dFZr2YbQm2Lhhw23B+62mW0Sbqc4xW7z8VdsJQndwP3kg5HrPJO/rONHcqboR8NEc93Q3cFDWVhC
cGE8n1qViKVzlLOznx83rmf8zysWe10bkOFW84kvSNJNRevK8sNVpMb5KwmFjwfpzN+Hv3nvhchE
yy37sLvH2pnWqELIBNpHf3NeTXI0k6rizFlasPhLT3+fazi3PgPyDTLItOD0z+d6cty05X7mr+pT
+Fj6dI48POrFo9hnkf+Sfs7S3VnF326AWoZH1COIyZF8s9+6Q0PCzbAZNBG97jAcEWEnYVpfYS1n
Rtt8ZaomeN34SELytPsEJALbCarrZ5rTIjPzZNCE1s8GKBw6g3ljuSgC+aDUqOlwlC81Yy1sE/c+
NwTaLZo7DKgGRnta1qjTW8aFJgLK3pcSCYX8Ro3EkqSMxvJrCKQmcUJGXSZBjLzdFlXKjmQeB5E7
qY0WsVEKUYPlTu6kOTGZz1RtioqII5bMOwjzpsL5y0zZnVtfKlzYxS4eLP+wXMTfkop0DAZ6glor
MhAGMHPZL0FDkrgerSWMb/8XNLDOBPosF9ecnHC4TLVtbavSRh31aDUmuL8jw2+5uHGEk6fpXcUf
8kZHTtuHUECMUrD8er4tj4ZewM9rnQuB1qpOf9a2TYgY8i3DLAdrC2uZfpYq0qB1mp4es6oYvTJj
jcm5XPSRJNThrXJna62dhQ0BGGnTRJtvQn0QfoM8Yoqib8APaSvOEkJweFi+Ch5hUARmGQzy3Z9p
7A+GJlMQiVHJOXfqfrBCIvaGAAFspa5Na8zRVZF40cpAu/SF3cpwlrDv4wjJQlQ1rMyIu4sH15Yv
0uKvE/9aoQi+6d/PUgbKm0p+afbCLJV0bli/uZyY1g8ftk8ri6JBXZXBOK4V3oPkzX1PniiwjJ+Y
xwawB3tRBkHecMXyqBZPmVLQTfofHGD4lODKXa761wWZIssxlDBuNXsNEUV/rDw+d6cR7VxEY6we
nE7UEDAnvFxTmDwe+nKvO8BcNfNeVsT2LbKrvV09IWQlI4xKXsASTbjw8BOSQw4zypxsZWU9Soe0
9DmNA/iCWAbpSUCjA6FPiLXRFCU8Pny1AFiuSd1QCa6qy4YmuoQjcDezysjBcZL+/VJra+wPg/gr
+wrV1DWFp1BQ0hIxvKLD3imNjtX4mD3UMThvPCNF9VdqwU2AmTVANY881t+0B/dv9/pC0L/JrHVx
FFSOuHVHWWbrzBjgSDNAZaXrgmOaCHBGfrhfJIrzJFf9Yp3HN9ITqcjoP6AvMmR1oQlwXA+HW+QL
X4Zo8nQYgDg3DKdFCHQzw/RvePyAQ/WsCcoYIzHgWz87fKmKUqy7FuIoFWIFL+8MMmvGh+GyMtT1
PIJvDISIXTGDdoeC33U+ef2tabi8U/mT1kgwxt/97PHJqJxKc1+dCazKC81k4+GTn3PFo/eId7Yh
1LVpbUniZnTFMkNB6JgCI7UXSe3flgldQ1+8HvRi3RAOOo7a5O24eUtxWHG8UHEdpOZexg5tTZsL
qred5Xi9Mc//PFO7tXviU81kmto3Jd/tOIEW1EkbBzHTA3vDYmtrMUbbjtFs8NZ50qCEcKn1MwJg
u0o2hNxETOEWD5gsstLLvSCLNPX8jE6HsXMS95YuXtpFjK84rON+QCIpore+zrqXSKMNpkvpC+Bw
XEl4MroavbRFflLNjro8QzrjoyTRu89K3mVNSgzblmUjLNsBrgiwifiITMpA1KcuPqJCyWIJ7r6F
pTWpOLU1daiEkRhJbMYEeHRjB2OawpwrtjNY1Imymnxu4jboxjP0HUa8BFYdwIJAVHmOjcm7dxo/
+0mipiz/A7sZxbLPHUoWuWi3m62ZQCBRCFfcObDUcVUEAREW86chRE8eZJ2HeWoAFUtISydgoQEt
1ERS6Ivjh4fO+EL36l6okYJSa4gjiHKRAwiDhPypaOZTDpdltCz8bFPqzmfRytarw+w6kZtXrW85
g3OFaSSJs7lff64fuMdMLdm075Hjq3KBl/KEtunrU8+15E0C5e9VXMW0nXTgfnIEyk3bkjUbfzWq
kZlt1phh4rQLx5Mpzke4ms5DLj9IzsAuv11TZmxUkgtEHEz+a3amAGJHun/9SgjHC9TAtuw5/5Hy
Pcpa6Qs0lV805ve+II6Xznn/2mBB8akTKKFPac0rKcDVAquGyMCW0DZrRS8i04lOYcvvW2b96uWf
oI6BXM7ORAndJA3to0RgtvlgThkz4LNvVWRLXlKUEy+WcmhZRXGaIQMPOWz/nilUyMLK3cqWyYHT
IcaKInFvWCr6VbfCnov3P6djwVGq0AR66DKTAb9pxl+tPhE+fICFevhqkiq2FCk9NAWNJ4MseCTa
wLBb/AdkqfkO7zMzm8pR+WnNCepjaknlLgbXAmDwWZE0x3dc4QasfRSDFeyFdN6Z9T5XPEICJmyO
I1/lEebku85orE2w7xVX9E5vYfqbJsZQqcI2AyecgG1Spc6ZWpsgwBZJ3ePf5Yu+93vlqja/bJDE
mJ7fffqCe5VTG8ZTE/lUIZxBOnOueFWouepa2W2+hVECQ5UkBEgt2qKcDd7lZVaL636hfbMghDB6
SyUnbin9xD/nH9kwCv8mnwOceTh6VnEB53drUV9VxUze2Nggoh2e84l4fEhImWnhjrHpraqk0TJs
pTWmKHavxcOwyFEqq2dvtEhApF4tjbF+T+QnyMMZdcCK78mmBP41BUXPoU+P4P0pTPvaB+4oscmA
ZqYNprkFlX+HIFnjz8agu4+hBZApq7e8SkLBLZv90A3j9X6HVVFQ9CLgsj66i3m8SAfjVdYnPX7D
sI//YrmBALRUhsZsYdigYRyPgqI4mQCRl32t0OoFpqmcTRJp8Di5RXJZCOXEc6Y2OFCZmtKKUcOc
+S5KhVVadgR4GSjLB4ApLy0XuZaho33AQBV1Qs+ujDQs8esGmD/EEZBXEnQ+Cz87SeeRl0zFhekm
kNj39AeEXFRxz/FFmBf8z9TMAQD0F+pLk6/TXCbo5bvXIzWp8S0PMr20MzyGze5+qJrkSjb0CXC0
y3nj/+E+LU+5fqsF1prQ5Q3o6/T0jUrPWnb1tmJVUh/pWezZFC8ZuqBqMsVFpOLlOo2PbkNUNXc7
i4OaO9V684oXeixsEeWzapxWcvrzhNiBC8gVdJ+DOGFs50+ykgls7guS9ZO0/75QFY2A5AjOlEY7
xKBlZcVSH4w7jS0DBCmnN0e7P4xFwt2tW8volxeElz1/+HkAtgMYGhwmlkCo6wp6IYJ7rh3Oh3JS
GcXW6pRa5zpw8Jz96+JcBVwUZYCWh7AhZc8JHHUE04CVrzEdymjOzHqJs1O/2nDgv81X7aq+lqHl
6HAboLfveJ2SvKpmUCAJIgJtaW4BtCBRWFUVK8QeHqClj2CJUubsA6hgrpE4QTDh8h7p+4rNSF0h
w4/ENASF55gQyAgbRkYSvaVVVtBj80pn6osFmH/xrZvUNcR3ZQ5pYUNWsbIgyP7WXqziB31pnJLO
PXcwBiTE62jM3S2F2Cb7IKZJuZet/0sremEIq6oA0qcRHA8jsQkCqUr/VevlpPrrzQCHjPu9nRuj
F+wGMRsvFDxZUMnC7NqWY+hz/wK8E1d1J6/mmqacKzZ4uhAxP+D/aX8/yzbS6SctxP4+yTdqzmeg
o/pSSnBJcdHvQnCBLlDciH/UakTOfluSj416gH8m8fUEPLhcnbXF52w1L62oH6vZx/fO9qgK0muA
tRC9BeiW3aCSHLofo6VDZAWBVkSuxpHEw4iVMugiNEbzOtzcsrIiyIPeTURtIVWueSDTkL8q5vDd
E+GU92+4jTMrNznk80CdYsWG+oeUKbLROIKz7dG3nFaAWxfXou0nQG/7wFiRiQj+e8sUzBhVTF7K
1bZbNHzpZsw0kEDmjkMHBWfDzs5DUYyeTPLrHfUDEafHwTwvUYuRYQK7o7GcNnh0BuZQgQmn5mhA
Op07Du0fnDNJMSWGGKNkRLjLmP5VhNn+Y3HPdr9mPezQaWMAbaYZTDfAZndiJfZ2W0+10eMp3g+o
IWeN8bMTjCki+z4ATttIdmJj37N5xmTFzLRs4OZ0YTDqtCa2M2pFH6eCmPfzOxBNMnVXlbFW7T6l
yU/owc1bKK4N5Yqtcsn+EAErKKdyXC85YLMI+AbGbBtrrazjUzaeQCPMeubsPsrNCQr8G/21Bvvl
uj2DD8lYzdcu/IoKLVf6uEX8yKIH5IWtpSxQhR5LLU/arZDIlXgMsw9DB4TnSbMjqsSOVK+dVJcf
9gFVXql63YcxT0UPNBwuRx2zEkHFe5miRoasv0rcwDXP7//Rsj8kPtWmppS3K4BCT3bVEFswjHys
/vfbCUNq4XAo7WXDpEcKANjolxxrYbPQesUmEP6MDQHmSQHZTi1cHSkyWkmufejrJQxTVNDzLQZ2
/zUaLrI5tsgBWZKmMrqcOU5/WCyDtgnCW2d3HvPkjw+Jx4T75be3pfEWtwahRGr8Y523Zg1PyeLi
xrL4juRUN8IwytGFGM6FVCAKYp1BldbZo+PL2TXF4j3w2UMWZXFDufDsT2qt19PCmCEW4yxbc2r4
cqXJe/phD0r85XHBXEXRAbgoXILs1skmCKkYTGPAhuocVTns82jDAe5cYRCEnGfiWiEI60XDMXtx
sV1RsnYzJk1tYTWqCTl4dLuopY9rpdKN5wRWslOzmmZ5thciaWTa7bivw00H51H5YVPK+VMrOzb9
gVtg3zMtcj9pV5R3zFtEr8E60ENsbEtxn5LJWEGGY0LJTthEbSOsiA8lJM/l7ej3aURqdYjr3KN3
x/40p24gSxr7F8a32/QjT0xtC77rP04Gu9tY34nIxp0dWepJ98an74sTSEy/NcTfgzR9dc3nVg+y
wPVD6Yxaotysec4LotLkWnfj5etpGDg/yToVeLUtAksJ6AjpL0EXxOx9nziGgJQUGA5I3LihM42t
isre8kdMa9mn2WYGfzniuWNWMpM6yQgcJcTtwazCvql2sg7Ic+uND1nUDzBa25IuLF/79I3rR36c
gLwVxT4Z1tvBuw3b4ohxOSgXlkb0bCsqvi4qpPsSt5t9ovRsFHlnQ3KzhzIiCtwlezgZzm1R+PP5
KEwGUFKgHN0MWJ7x19y8ptzWigUolmsEDhiRcF5bUpoVFGtQalYy0WwbChWnE7hofElEjgjs105h
wuQPIsHKEvnNIUONlA/lk8oyCM+9jnNWq02lMgQZ+OnpLe1zrNLSAXLxOok4oThoCb/Aiswnl8Rw
+8Pa6eUSx4O3Y5rkpBOkZbvnjkyl94aLTbIoDaWyGFU4ua+qvrAarvwsvROgpC9Og1bt8yhkzlI5
9Klgg0uHAmaLoreVSmC9vIXhvlg6KknZV4+xaTIbnz9xM9+jpeahPhAqboTWP3lYThtq602l3t8L
KE6MDyF1uJLtzFoUlA7OMt8BNDgFnaCn0DbbA7CIPQ/Col3WxRQE5wpkKioHKjBBy40g4z4j8C+T
ek6qiK5ttLb3jf6w0rP8sbk4JXvROjA4WndkIiJ8slHtQbr+wotb8pWglm5bp1DfOTtHdooEHXf9
wjzyBnId4H9vMYbiymE52fYhLl6CtWOAgOkBOsf0uHs0RwJXDIL6nm6YeqAXk+65Z0K4GjkiOwkO
pP6p+QViOZCvCcz5+LDAIQOxDixDQ/KS9znQpwmbLx0Z/wVmNuPxuvX0sjh0lW4NuwmTLNDawqV2
NarmmQf+IugXpzpV5OEjkqQKRPiYNLzP50nud6/JhpMalElsFSpxk9iLkh5oV5m3zBWoHYihesOl
IdgI5XpNDde7QgRb2XPL/pgOju1AD99JZPghC/wEMnboKEThBNEUJUR1U2WvShzpcY7k8Yr6EvDg
79Yarbtvy13fQhX9y3+zwR3Tq2YA7la4V90PHPXlB9CMOXNLvjQs2FCT0ou9x6GmJTelnsKdySiU
gu9r8a6+HNhMgGxcbqXECbXlU5tl7Bf7gBTZhjKF70CDzDrXzddg2xSqedBPS0L+vKC2tP8jxOHQ
0P70v3v9eoA4AYDU0yk55ZP9ErgXdiYrQBU2goOAp1TI6uR2LPB/czl3k4XU3bCnPlEbCaIaghHi
TU0/1PH8krtUq1qx6Ot5vIFOE1l/1E2JjXUywpY12avm21aTOqe+KqDeVTTIs8vO5iyuu/OS0fN9
NOBAqzeMR0H9OF716S+N7puNyBIstzAHWfydLZ5dkZdqPaiTvTa8s7N6i1fD29UUu0/rV8whTgVE
33XPUly47zZd9ka1XU9tmUvMCMUe6uoJ5YqzktRVghQGXtAFpL7dQJfwHqOGL0FQe2hoG/jCvW6p
X0stUlhv3w39b2EuGeWNPViE10o+Zca9zmYw3GZ6VL6U4W1VAav32bPEBQIXamQ870jxIsZPwLiS
gB6BpBu3p28B4FlQZof/WyBStURP4R6mQzHii6qbyXj2ZYoE9JgzXQcrYF/o1DDJ051cCizbgXav
iegToar8nyKS6HlOQDEamR54WDNtgldFE/BksopEis2mZHblJuw9nzYqARbNDe7Ve+3G/Djd5DhM
NJG+ee/K9emWKEhQHCIhQmrerRemhi7hUpaSgXFcEy2uh/SMqltmTFuuDssyxUGsFM9wgzQALt5c
0zGdV/giomGs+lFvNUsDuoA2bCgXlMiDvjPGq9HsRhY69jrmtG8Uvx65KQ94N5tgCVi+4yb6iwTU
p0dgqcIpEhmIi+B30Q+kgSc+nVEDEJM7eIQ+bhYs5jq1BSoKqQaAF3WvRZgfVz9d1Cy6tMiLl+tN
xd8287BCjg1pa843fLyY9yS73uE2qxr7HZIUbt83qtnM1aCWUq1aOZ1JoP4aqwuQGpRY+L3NLiCY
UyFdn5/E4A6Y1Xu3crKaniZxvVXno+A4wUSvMQzDbPz9zxGAOv9EAJllb9AYj8C8uXY0u3RaIH82
Dc+Rg64ac2E2T+riKl42fzFqaj5ZiYdLbKewOkayqK2N6+TTGoXZccrkEPd5PaXW/3obfXLjMlI/
yaKRZN5/CXMzaTQFeW5vHYYDOLqIUiAEa15v4FnnoD5eMg0eYOvax4W1mHgfba5ztzwvVz3+QNQQ
DYxq2JNdFgBXhz+20A57wjMZene0kxm4nGm5krxS66suc+rymrotfoEOt5s18gRILs7MmJ3ooSsn
QNYaLmjCwFpoimvNZtqKVF60WPu8JKgm3g7GYLqdoZmoI4VjHgl888wgnEtnWJ2IC8PDGOlTfxui
3bTxBA4Iq2H9gULA1AjEANpY52m36rp13JWazBEKj9T7WHV0LlOjmrNuHCGfSxHF82EHWP2jKq9s
p470la9bgINRHvP0lYmrJO5hmQvTAJJeYmggej/wtTmHZvbhSv3L0Vcvy73SrmorHeghgmcmCRXx
d7K6I51XDwpQyBtydFctdprX+s9NYPSJzRyHc4m+IRj1kQ68Jb6bzfGmBcbgDnh1y9rDdQtqMTa0
5+WvqIBfIz23+e2I9id7gaqBa1rJQHfRF6tDr6TUVD+8AVEX84WJ9/WiPI744jF2aj/oQtvqfLVr
W/mC0fuzGtRLPmL4rhLCZKL5YZY5y1GevfZsdVaxWOm0X/Ak7qvJY2x11XuIhCkb8/fXwnI5ehfw
LpyxtdjqZyhFyuWHpt3RDl2RgBbIztlcrvyQGEOIKlgVgyn8XyZLZQn61OF68/nsPVbonY7MbAcX
u5qU0lVpfRpQZwSN8k0TtpX5OQ7imRYH9/uZcsC98mWntSdspJqR2/UFNl14EsdKcvVaF06mRhIx
DyxEKyb71eqOgPx5hK0tDr2Vfde0Rv3/vn7f/f+5X4okhdteqpqNRYbHZLfwd0clyBkPzD5tXaL0
wdisE37RmtXUwt1PfC2Mlr+NjL5EMFMxVF7NheGJzXWq/RUeArYBpPzoQ01l5Ktnh8Kl0SU1gt1s
nlwswLMAwCUOci5jp4iIVeQbbiLVVThhpsglvK4RgGGOJXBj0XG+ekAQSL17XPpIfChNZgdUEcoP
qv0F2I71UA0pSnDt3GHWSQym8ugNabw0pEUBIl8JZwj29cYwnccyFCbTDaakhRQiD7JEB7L/dsUx
1rSPBugZSwpDCBGvvrOQeXl/JPtQAqWZkW2lQF7/FBk04mj2oiDmu/4hqYrjZmSj7qwR+fkAk/wt
crb4e7ZcN2G+vHXW/eOwGFWILvU7mqqi5YMjiHg1BbYP/RNXudIGfDa0hxMYmo/XsD7qB5qS0uK8
pVPsLK35NgHJo36sQpJu6n2X21nVnmV+fHsGCTcstbQWtjEK5yn5pSMcNg1S0ZcUydrt7NL0oJT9
lgfDC/vpKcKrm6/EaqBsTF/9MfGVzaDKqPbpmNkuL5EEesZt3P8gS3HLxq5N4hGj265r2Hy6/vAz
4i6c0cAWCDNe1Be9CYodtUJZGXKwb0gvAslVkP7BrzV7ghjycg7e7S3QEqEEMzR6yLltgv0ubGtB
rdg2NgOAzkPw/KDizPXiXVOSbOGhL7nc36FFVvLmeSfHG16Swo9Iwb/UdGkb3xvAsuduWpr0S0Do
Ubwrb+RQpUbQaD1WJuZ9hYYsGHJqPteUNRc3ndOmEoR2EBHhbVXJoeR1hmPecbbWZ09BXewjYe5z
jq1SXCUroD+wFmP6KvAN7ixWy3a8J3wwtt+UHtdjaukCcunGNi2rS8YSfiSt2LrqwMV/I6aD3C/3
FWi179GnGwhDG3nzhw6eL1UdFii5RUHUZSuCNpGCtnnMFkpkSn7ASP+mpsbpqPujZxoDbu1PdGNt
Y6XdsZTZ/h1OdXMASxH43Dl3IavQYXozmxegOuo8gLP+heNzC1wuYvIgLbRUXuiiZniYr5kJ5h8x
aAsok6Lwx5hOl8nNYhA0fx+IAyJ+X0FbaUHbKD992fvKyYGK0wI28FtKZoV0pt184Ck2z0ycANbm
i6WC6BM/6TOmYFFjnqI9QWXZuEjYyz1XDMHhACHAoR1ETS+z7+pXgWh8Wr0KKtTpUTjeUeIDfEgd
cLqMotzuESCJQG9zxAR2xhzAg4U935PbmDmu5tTr7rE7H+X+1xdboOdZdweGav4Lj5UKOjUBk6Fh
9UGUFTK3/VKRyLpd2li7NvJbo6eWU3qzFYaPiTnYpxMtu4VFibmilGoY1Nmxvpb9EdTeiDe4Q8GD
5fcamHUjB6COfpPYcBgouXnJHY6EBtZl/FYKmN+VXeucxJHHtPJ1FuMl0wD7dxUJ5uOSa7bJpVx2
TrbvXZT9YdPAAxQ708m2Larpz8ahDsoBVpG50ia+igy7MNVKrF2V8ggX/x+SZv8k+BV1wX5ZChw+
YRfg2AhRBLhGVTlFEZBC3DEtvUkf3EBBFG3+nCg64JwI0oEoUkILu0KbatFvROy3PXfwlkzignLd
eMqkxG84adx7GapzlcraA3O4ED7S1ruUtaOXUDbdRagOORRpzTeTSarKm1kjC6cyTZt+ulc5imPu
zdjTTu84hFu127wjT1+GvACLdKyUoxXX5P8N+syQRlp9eafypF5pwLvYw/5ixjvTO9RFq2R/4SZx
BMLPbbjhJbXRg3Z08QbCDAVseXeZW17AglcmQl0lkmpiHS9bpNMwdsYUuWudavGCp7zpQ0CRb1OK
UAvy2Qyq9tLW2Ofxhs7qHW2WNRF2kWgwb4k/KNZ8qyzPV6mtr7EogQBVHat8z5jE7GFGm3d9UiS0
XAUwDVyRM6tuxUw0skPpag/2GTTg+G6CyfsZvvbknENCwY1HftcboW7vqy6Szvdst0pQwOcdLKdW
Jlm59kV0M2WMak62j1WayPB2sN7PvlQjugr8ukWFJHwilMNXSHrCzAjbqMTR6AiwCNWZs6P3emz8
ZzKIYTUYG4eF4D4JSzE9VRTU5gotoKEh+CfsG3/Zhd+IrL6ZXCEsqa9sHGwIV0kWJM6tHgOFZHrH
PZg7tWIzWKvVFuaK0ux19vkc01OHM1+25sM18uFR7pxiPaEDMETa2vhbNfzbkNwOzzMAnLogwrIK
cZSkbZLQViC6STLCtzi03rOjPpYQBaP+jQSM7b8HHvRgFS3WRsjNTY6UncW18e7SdVK/svSLClKD
O1YS+Ak7ySjHMM5b47TPkz9593AunBxmU2COxZ6ZV5oVRsPWZGoISQXEZEgY1VXeFe9l40TPc9Nn
pNSltDZCavaekuaXLezlP16EHvVHEQyyA3PE1GdIi338VPgIep52rlkjeUWHzZFD9hsoYKr2LSJU
AELttq4riYARBJfNhtuNP9IMt/wNh8l2uWupLUachCLAA6NXsPHeD6Tx0IvPehxXg8kFHLnSaX5U
QGnopyuKQ95odtWIhxeis6zQIUExSLSTz5cKq5X5cyKeLet0iGKhFXexbduqFuprLaXWPUMVeWN+
36Kapjz+mfaCHNhndaAdbmkL+9n9WCLaOAyx/71qmlXGp3XpJgaxNy5QwnCCM1xgSZ9Zp8QSxp+z
173xYdLmbV70UQzdvV3xQfAd8Cz8uXdmOWYh0+lHtxF/DCSxaLRIZTP2qB/JENTdkMPKNae7el0h
0ZKflOEB41XLB9Vwb8I6mZg4HQWlnY4HOlbFI4xRj04MfLHPg0WBQ+DbOdBt83wDSfpMI4Or5Qb1
ytubQTVNBlUsKqoEuP9cP7SGuPbsy7jkZPHYYbvBZgVs5Jk7Ip1z0uzyJXU/ec0n9oHz8AEdxuYn
bQAH9foIlpjym+6UBVBnwH6knaWUyhDEnpUn25boEHrYmK00F7ozsRkRDJ1d5HZK3vxbOl+26zjG
DcB4z4nEWlX5jdSh+faYW0S9ydHOpm9bFHkDgaCZsp20aAflbyZCcfMVQKg0p0vIrTmsfZfp2LgZ
7aU2dsThjwl+7f2o+KYF4qVPhGqAZVPP6GqS/IvHNkAYHNUflODo1fRKb7q3wUbcGp3trxsXVmNU
rfF658T+IZQ7v6HLSEaauUU+rgWwI73fx43mWw7m2RwPM/SgwwbXHokQoIETCtOCjoV6L5tqzlKQ
4ilYdFBmlcxTcUpM959OzytSveZG5eZcniJdv3ay0pX92+P08bVlovRwggIip+j4OZwnX2f/Xh4k
UHDUnhIQQNO1Dq7BaEzLb5TJSVy9BZ88voOCggb2mjg8rto3ZQ7ymvGZLhXxHCOWEJozM/gtFOX/
/50SGNSCN1YckH1kylOWaA/ACovSWUvUPR3W1VKBq4HC2dUhbgO6AkkZDOfByBmsIfzpZ2YYDXJj
Xv6lMtnnpUN3WoBWH8tjxO35cJaj1XcDoJegrPm5wG5dsQiP58DBfHX7Kdecm86NV03cJZTmAsxr
S7pD9dY0WDVYZ19gCvEy+6YAFOtERRbrn18ZFZGML0kzpiUePVPLB67T5/8JWT0WJ8XBH/VjOY1u
6ze7mt/QAJYJpzugx3PB8ZUQMB2YYr9NcWYahSvwJi/O4kB+SG+td2yvPAB0GJdNUpid1Ic6rqdI
FEvpRUgN/KgaC970uPmZKPmUAQgs2+GskkH3e+aW+hj0O+WMtYSSaziGPU/ePFonGzfZ2a01VXZs
TiU7UzxBSHaseWktfm+/faGrVNWb+cUpuU4OzkkiAHB3x8QJq/G2m2VKAUguCXyNTZFQzV0xlZt6
4ilNCB9MOm+2TB7aa0RidiHdIUU6py30mXGQfoOwfjf/uhwSlWoKICwm3JYmIVxy5cFng2+m+bV5
rXMNsjN9xA3JpKugxtHTrY+q7vdZrmB2KnPTBPBKjrnIfQp+8wWum7YoDWkXwLmnhOyZVGmN/RXy
KZaj/GDqAyJVvmCQlWLmqL957XkzU4QjAl9kwqbl+U+Wng7bx705C+kwvRx3c1b3wFACjQgjAue2
+3NTxPJ+Ahr2Zz9WrjKA25MxTI9AQvN8qdbGjsgMf+x1QiuEbpGpAluQtpUX8dHiQZyDzgpmRFTv
UUIMgHIfgRom3ghAfq/hDhg5qjmu3XgXck3an7O9m66/Kgg0P5oP90Y3DxV3ex4YGTnFGbdJm7kG
E/t8jXEbOWThzX9CpxVbHxOL3Bdn415GX/XXSa8khL1nX+MNmUgkunoGo43N9CINs+yyBKjb4mez
m/hxGZrSLHL9mlhnqYiMDRyniuZTxRTqNMZsiRBfa3oz+7nBNnYUntgNoBxk4PYd4XEzaiIIThME
dSptIyWh22K6hpcoad5lCpbw8YneeaFVkAKb/PWLZ/VZWK5Djwnxa2itY0Rzj8JQgo1l7/WSESuO
Gk5yLAKsZQt3r4MGmoymrZ1dCyLZ33URenMpjFdYaNnSbztoXjSb4BtcRFLHfhOsdSPuG4o0jL89
qkdzJwg1Wjf01AYybiQYxG78cssJC5maEV1mJoX/0v7G/w8dNtW/KFrsEAmhOU2BOsP7N5L+0gyM
yis7+wcT8CJvEFYbiI3Rz7a4YPBVeySqt5XgHgaM4diQZth8kUMxv02FlxVYJFSL2UiW1zKs4YzD
c6+s3nxHGm/roCckilaVRPH3hJnWJNwCL8vrOaj5Hb5nkJFEE3tqvcDxQxIGPRSyooFLVopdxG80
dJcZBTELiHx7prpttObsm9pXFGRsT04asqsWLDSx28MjwV3zMTg0wzdJ0YOV4yOQ6HqzDn7ABNmJ
PdAQnNEZPYsE+h+tvnIRIhKphHjywT0zhOKBNpjC3cH3iB2iQ9QjShzOuCM3AhAFdcbFA/ohMdLW
rIzcMnErXROvkz7xG3P5FRsTcyelog4n2QhmDzsP2TE0r7BOHQza/DID8tftTnoytx6vefQ9RGLs
j3vG7UzsfakAmfdLkSG8TfE1mfsCBkuOSM/uZ1wSXWc9hjvKe3vWA41ckKEtFpxHTuB64DzcRrxD
Wco91Ww18TFT0RHB701LVXln1ZMUNxhLxPfrOQ+UKu5GsUWKiCjX0bvT7O442yesGyNWU2ATFG6o
oLSkBaARQYfNECvw0mfzO45jsT+9dpfNxBpPdhzt3I4THilFOZ8M1YetKYn9+OGYKLipEPCRWU5T
1hEelnugyq+1lpQwomZN2qDktvtry1cHtI+MWNeEOiwnaNkD2NEp0FhoqfwWXzX3iXxb0uUEU7K+
dSMCY7lGwjZnvzRBk/SF23vZPDG2aTsZZY482YI24YqOFC5BoT5cMs5dO2VwEwXEH7eUF0wb7oJM
OUNU+Za80s/jTmRig5ezGT1X/lAMa9nXnFEcBf943fZw+PzPte5jQ5nbdZEiepvnwnzyvlktBQe4
BBL2UHmd0c+IYLO/dsdeehFkHE5LoV4zqqOynL0pXgxuUinwV2HQwjCNUCTfdsMhmvq8eRhVdlsy
TZWqabb5N+YS4HZTXf79Ku+G8br9SX55d8RurVSwS5MXbnfJ0IauNhqXz4gxw9ihMW7kbIhHHX8i
smNVvIAVk3ciuEzwLEJ8JpWcHv9LGs858ypBdt6jQiOTzOmnSvZRZuKaAwjSUU/EqhXB7WV12QVS
82Xdtpecc2QK15l2OEq88f8ZvJqGst/Vmfmjv+ZGC9tSe8sI76ie32yAgPsoMtYarluD6cXJjFdm
ATZw3pePOuG/883UwsZtLP1xZjZjieP54H/79jLW+3nP25CsXoACPgSOP6EpdftvtYmEdrj4m0Cs
PA9k/hx2ecOFXsI1yFlfYXSNgZ++DY0TSlFVf0yeLPh9KrMb9V8PTW8klYuPqA3dRlk10umR2NWg
A3uGD4RTVmmdlvCdHpav4tuGwstDaZkbg5IBAQAFpC1fyG3Jul48KC/Kd/LggF5tukWEMH3h6mZb
CHXhIb6tOGkYCAaAKOtxB6e/Xf4IAHHelJrSQYiyXWi1AhHM889P1kZglMWEtRuLyfpOD3CMPGNH
ZFWvQbH6sfu8KZszQrFW7XfTe3I3nc2ikVM+Hmw5PouBiZ66yGfLNn6SAzZdG9cAgPu2RiMO7go4
MdDS1xDTkm3gbPzjiPuLO0Dzt8s37O1H7Dv0EDkpSxWZBPhQWDiDpkp3wHeIZc/RUGo3pZANKXrt
0sbnzNWP/KvX55m9meuqLagSqeeX9CcG5bwljqAA226Y1Fil6azG3xv3Me5C0gG1lp0mu3opt+fl
YVJRBGblglNjelk4o7gItamsaSzPRyxyEQQxSSPu3LOVwf1B3AYlLj9vgjqWU1az2OZsj/JlgcLM
TSNq5uUY2oWqQ6OKeEJJsragekYKJXpH5UtqpNcQfkhrvPoGtWMOxug1IyM4C1QJv1Ex6ZkmRQuJ
uvZ17TgR9lT9P4gydPl9HpxkJHTd5yF3Nf2bm1byeEe3xXAOCP3bXLOsA4qH6NifQKk76fO1QYcs
8kAbvMNbHPhZCzpwoQIyQG6/V9Z80mvDzqopYQ/zXDMbfPAPA0WS8n5yTadM4/uYNmdyH5IGPmoG
hELzh4hlCDFTeO+gaO5eLQmvACYa2ByBSktJJHhhHAAXtimIBxPmJaE2e2duoWxOc7RFc6WiM45k
KMOElUJfg5k6mxmHUKojPckAS8WoQPNmV8/gC0SStktwXZt+NwrOidCSAhmXa4DwJvBAJRT7pbOW
9PlHUx+IJqeOBKt47To6ttdR3T9ti2R04Gulmkcx8p4INT20rz+jRrH3g0dm9Z6ciBa0qtY4TWTS
NN3vGB3UgvZ0UD1F1jZlB9UfoY0zFHYhmhfHCpvjaYYCxL6fXbNH56NYk514+gRD4+L6uyTVC4+y
3WPEkmMIXLM8t8SOP9Co/YsC+Cm7miSufgbH1Wt5h8OInx39A8sdYu75nAdamBQa1RF84eTm0VVg
ofciI6nSSSyWfTCobxy8UbtVgo3QCt2xwwaPPS7dIxLdUfZB0c+fNXKV4S95wvCDcQlJMePFwXQK
5hXiFQwV5jtmWMEgN4+q6MXehoZwMQpDn16BHjx8CKIFoGCYRohqFmgV50pMm97KcEqXztXLIDVr
7s3GPyiE4oU+dMPEiU2niKGBR+/n4WZYOezQ3KAqWUIYaoXO8xHaw5jimQDYHK4/oAigZO/X+/EB
aItA+6fDFKS86M8XU/kZdn/nuJ+Ujmmcc0T97eTEH97L4k4eA31cX+lnqq9/OVCmZmt76KF4vtQR
sNJXit5fI+MyNBg03TcMl5cvWR0uiWR+Xp4amhvxOUQBf4bLtPQNG0cF9SuLzsPAcx+Kb8jkRzeI
SD+4XXKs55z7FtEZbh5SZsjBX/fSlc2WGLudFybtxkRCRfKszP5y3b9VttIB2OR3naMo7mshuU9a
Xe7pAVHS/0uw9CBoWKLZkAES7iMpwzt2XOs8o48lO0jfCqxnabacC2p8xz34QJ3Hp8MwwIEOt3Er
7mB2fXnxaz3aRoduDYb5JKrt+sx/uKLnghmXSj6VJwdPKC4PKTcAKVNDxqAaDUn9UyDSujHrfl0n
XgYoNUhJFZ0Eh/h/QszotbgJfq2AKO57XosPsN07QEjcVkGVS+Qr8gepxJk/wTXhNsU1uoTTm0sD
xvnWwIPvHafEqRAGK0SzN917jaudJ5IuZPDey8M5JjbHOCyMsylVwv9Jnwv97YIhN91kvtiLA2WD
Qgs9El6xpF5c5an2LCF8V0eS/Wof30G04DxjXkkvvWn6VB76be0tYl6TDvKZHENm8r2bZzNn0pj6
bAD7+cywGdQnVVjcWToa3hdmzthk211XhBZrprLxevt5/8AYOgmaZJWOM29HPJW5pFmG9kT2T+gc
UWcUJflH6cx3LTnt6XYAQfXZHavU3FYSuKJZ+kvbiOLfSSvBEhMiEwcqBofSapuecOccuMrS1gkE
oQWlVLLxIJm1KJXge8blvEAtwkofERUW5kosXDsVb/6+i3uEak6BSuyP9WbQ1TrF1/zbWgbgL1Sk
6HGAPtSAdSMddq3on+N4ojevm1rmHTXyBIkKS1W/TSL0q6M6CU0GlUBvazRjRQgJ4uiP+Z2KW35D
smpFQjbCyuObm/lkBqSNOjkydCruRhvJzw42bRroMhWRcUYWnqaFdI4C+NctjjcobeLiHlTPHZNI
XlBEAykCdtBEOX5lSrvfeTvS8lbvuetJzAj9mJEb/WhB160tlJlh7prmWmz5CI23owS4+0L2q/VA
9xngatn7bQrNmMoWWbelRXXf4HyCPUz2tsPWUtu8Jy/ek6a41qaD5iEVMnDhnY4GDMldnJS8PLIw
n3K788PjSP12rtVH7Nih+CFeWfx0povcWtCnEMVeQFU9RRC6yhoCPox37IaAZOfCkyil7iIuG5SP
MKFQ0dm3pbsz7rzx2TyXsmkPw1+SDapRv0reIFN8VaRlVjcwr7n9hI8C3N7k5Q5B23aUC+mwNMFy
BIEDq/V6xwrYg98hydxtiNg39Zk9YvFIn2aBEp/AUT7K+JA22oooIGPkQ3snHGR7k8tJpLbbnj3C
0saVRlMCxrHArTPzqZAJlHLeYgNqub7rngjeZQpxyV1Yw2kt21MK6Nvkv1EsWMW6vS031uzdSIyM
hcPEMDR/0SdRmzsMiwoAbUclbnkYzd5l0s66voRQ+e5h2Fw01ZfGJEdcV7+al9HE6SisYRwwabJH
BzNx6xAjltTbiK5ylUI8zoY9+Dx9nuc+RuKvoGh35S4Z5b7XM/Ozg0QUag7DBJH5zPGtgcZLUkse
tmEws6tezaJcuP3oS+HSsdNeIguX0oOcyxyRYvjWtzWr7RVXfY/LS05N63hYXkCoHYwKUhiiVsxK
mXx9SYHZkylnVycXgkXrte/9g/S+mD+NbjJ/mDDI70oCikRJJdDbYqgrGhXyGF5T4iUNABOk1KIQ
lCtDPizas1lZrq/GrRbUyWOrNpoGj5rlKQwvLjT3eRV/6NSFle1IRPGnrDlfUz4Psvm4Wyc0b6Ny
mopZcYYO9Z7ayCdZ05JIxRDgckRJfL82j43ki90LsJ1Rsy3feFy6oaL8aP4coOBRMDAI0RcFGZU4
z6IjdjZVlFGvYheK3zyzi6+7e+oZkqjmTgntzogKzDSaw6cPot8N8jGe/7NkbUeLvNPT/4nxu4BI
4l4BtFw5/rrxxQl34wfFAnnUwqk2FatGXsPzMBn9+OF4QG8aq+ygGe3EaGkSzOkeIsrULgcqgnY1
QanaiqzWyWFBuo0r8YDYJRZPF4k6r3Ov4Pm3A81pO8Vw/65nxUVn7wuN3/zxTUjogZExOiYszwBM
MMvUzTPGeUrK5Ow47/Nckj02sdhxFXYNKPd2RaV3BWvc1aSDJKK/+jwjr4z5SW4Tq6knpYZGYCum
yi5nKBZZNQrUqJkzFdiHu+AzeXw5EgmrsglMDH73XTtvM21hK2G8JxvutM4t8YhFldiMfU1hodLJ
o/pU37ac2UkQk5HFyW/lIJhln0JEltwY112LOckH/CcMt7sTW3J7tPPFrRpx1nUU0zVb7A8+BpSs
GmbATwFMJ1cHqcgMsgDCnmq8h8ENjg0CI8LMOiEdIsRZU5COv9aIb2Nn/5UGtE617yaO/QleXK4F
95MhXpFTJD7Mjnar7oblH6qtEiH5MsqpjSVpf3qQ5vVYqc30kecsW8m1aazeUKprQFfj9sT/43dB
7yeNT3tRbCHRIpfLq0DiMSwt2pADkdRMuJdcknrvj65hQwV29UrXdozVijRxGJ2bU238R96yN4S7
F4N+7NVtH5k38vQXRXFmv0sPlvRC+g9aRTCkkWiNmGXU/g3ILb/qoYz2IW/rsgmxCO7AyZRd3Fjd
LNoMB+2m74dtWr6I6OdeWRHrRXROTVvjV8urkjmkXwGo96MyYEY3a1PhRlcyxuZW4Ul9nxEI6huy
v3mx6P0jOX9xb1E0Y1JipydXyjdNlz1pbCuK9wO7cE9RYodtMlvxXMHZr54qakRjc4Jo50JpeYHp
M1EtxEKCvaeVtyNxYqT9XJaOGx2iIpfCQBuOt8UOQb15qSTFLa2RVEOxEXdgvnJ37psyJqLnWMp9
DvAuY/7zP56mtqR4RB1vD9rSLMAwakekJ4eS2nq0caobw5d2u8m5ddzFmxeDbSSBQ2HpUrkekYO0
4k2Gdt3WLEDk8Nuq1Zel2mPnWvillI31L/4S9hKRbJoGfo6Yk7ulJA3XPRsUS9MkzTyxraPRnthy
PzFOTwJpC9MZ3IbbMRHsynNnMgO1BxFTY6sdC7fPOkouCmM89dVCyXVy5kBaFhaHb7C1VpgZg+g2
66BTYkPJL06dAZpC0kicA/U2ljN0XuG+QGaFDNLTqvmdMV3ZkQtMuiDcVoHc0ODpHuIiDe2bNne1
Qq1oeiM4T71W7wukggaAq6x40CivGENBOEUGzw6/w2ZIKDTp2LSOuFCEQ7GGKr/b6c7MXS7il51n
E0WuyFbanfV64Igxyl1YGMWrNhU1iC4fATFLHtafg5aK8BrYFgMWPrqiK6ke8Nci51M0NBsc8/gQ
g+fvk/IKPjJL9qRbtJFL9o3FcrJVEkqHmyHI6z5gcgx6f8d+/R5SPhZcNGhllPtwUDHQhNloq3AP
qm7yXRKT+6xiu8/7jgOJ7o/DUqO8Ub4BOpZqZEORJRVTJHUUw0Us/guHn3uG6lWvo33Id8iJWxpq
TbaDxhhhC/oteprn7LmiqfN/vBvzLWa96W3TXtNisNRYv5dHddklmdqyucN+XoI+6UfFI0ads1iy
D3awrZ6AXgrBGqcAmhGQY2jUYRksoqoCyhOLBNpCXZNDhBPgvpYDwmXZbz+/PeZT2yYgGr1mAZuL
A6T+Z9WrCceEMRej6CMqEX3q6nsPvEjAjtbqByvktc3dau3XJRWUjYtRtVJ44XPdoWGL0Wp22Y8c
MJKjZft3S3PcaGk/P+hJK4EZSZNuwz0cVCzV+cMPuCFex9804FaEPlbNA86w23xCz5STxJQcxs1m
Fl8KUsX8APY1tRcm/L1D3Yklat6w7hydbMWIUpxw7BSlQap5FOtbd1oxhn7JejyktA1GqJzQ0pDi
wwqrQd1JS8ybEwbQmHlpHMvtKav55DEIduAXGOopCc9r0pAiJPwfN5Ge55prc2z+/bZYpvI02lMd
M1f/ZM5uCvsp21DmO8J4HzPXjZIponF9VBLwIaXrcr8MKaXoYGxRuqaTnEkd3GaGPpXW68pc+uoK
fwCmK3qILHahDU++i8EOvfkVC9QGGgXv0Rqv5/BrK8vRFHCJrqo3GYFuA2jSEFYO7BQ+rT7sy7Hs
+OqA47jS7GCzr+hydhvRgkctTxMmIZ3Ue+jjED9lNBIME2cqc+ar5wdxBaiL0Bie2cG/IUUlZDbt
2lawMYEB2gjfh6GJ1M77jF34ow5/UXYUjZQBo299w44WM/+gOtSYUKNg0wFE6kTRuqRoIgxwCJL4
BQYMdH/gekTniZ/ybUY6GMCJYbJUkTyJEDGX72tdVmrpLSqodb/9IDQhXUQmKYhnt5EBqWaxgnMM
04/UgX6eahUl1evgKfGIWuBZQFrm427j3JwLV+9oxt6+G6Kd7/aycHsfgrFTPMqbKWfH/NiVCESO
utOc3VogfI7+wuv3Q9cbaqxxEB3lVxOf5jWa9QO3uUX5z/FQobaOkHUunv0LQqy+qYS2KptTSlQv
EuQSQOzEPv2Zl9cQFgPzoQxCbLjsT9I/opJ56K97vpYllX7BHsdgT10wM2ZAf53TZY9c7iCS3bGk
d1R15n45bdj4QLejlCB/9DaQQAZRQs9rGKczbqgZAdU9MTyioxlMrXn6NeK/ZdhUZae4nHvbe2LW
cPQzOo+C0voz0N73FpiRCeTD7ADYajZkEI3wKSfkiCufYdo0nqMpv1l2tidKDeYGjF5LqD4PJnpU
4l2x3gPSkyQTRVb3CS3tmZ8nIY0csTHyEuinb6QG0R/EOvGi4EbFOZ5WWqPsp6Cv5RA2TwLm11TU
xbdJYwW4aZP6H6296xaGsHzxCds3/+FCA+KxBBuTq43+couPTY+lDUWnh0erY+qmRT38h5rJCmDY
B9qSus91UY0In1j/lE2QprLqRVtvGc/nhHaKqaz8mn3dGmLmP2+uv0tNKRBkZT19vMtbZSlt0yAQ
S9sAGgOexN7exQLIzdMrXhx1tBl9Uk/wC7bfh2ZbtXgl4sHo467JTgWE8J032Y84eyjYNYuXGgOm
qQEOqKfMjgcNpNlnBfyYPkg+HDTElAj5u6sjjps07BONg4oQCUXkeN6Xo1HVIzk4OyIfaoUyyfqS
3Pj3MQnH03FMeFLB91LaH/HvwRFlse/j9FYLgeWovK8tcCxp0ntXU1IhkmadP7jJ8sStH2l1uohe
SvKsVDM7EZqD36XYl50Q2EAQhrzRX++2GeOmhW563GIoWg+xU9Ylhvz8QPy//KieE1AWQqxLGBmw
MHCSAdd09shGVzXbQKX5PvO4BEoAx7BNNA3nEQy+r4L/tqRoo3xqbxBhNYk9bB+7nrXJMr7gWdv/
n/W2hvPtr/jwG+DoSdsjnR0bBJW9ufx5510iMlbn8eT9wm0T6RSIkH2/9LFKiRVW1FleKcNz2o+/
CBB/kqgNkG26cQ8b4878gAg1OWJ9xPG/8u/vnD7eXrRwvLeuFV3mLCj0uzmlMReq0fPwbOkCR3ay
JW4J5BgbnPpLp0bHyZkJZ+ks1dT2rxOjrgCqGyWDuBrWrpJZlsaY8ujT7LKZci4A0M665NEc3pUH
wQOcWLd9FVKqjIHXdbQPTxJrtiIwoIY//Sc+VD9wTbxNRATb67OHJXXwzMNqnJP1FLM0/Me3yRo8
nBMPKy9LJueNcfLRruvksJguAuo5C2suNMBQsjQbxUBwjSSWuuozFvlwy40fSZXXVEKBxNlhqiQo
OvdgUJfYaklmijtma2qB9E1Vywg8SujjFQ38987is3y6ypTfmDnAIuilm9gu9MV8qgV3zXj/y9Wc
d+2YkZCVP4pgkUdlSxW3haQm4cQ4l1vNXirlr3I2Cdp+90Ve/QVMDrAbNYmOCtvbCi40735Ifzfl
dbnwfPqfx0ZW14UVhISdbaXoEnlheOK1u8SdEqv+y6EFCS29qazyPa8HBxzjH9yFUSpcvKKo8v/t
iJ5oz/EMINsjmrGsQVBjOaHMdk1kKJ9XD3TS64eKOj+AlkUq2oKLerU1+IN4AH0q+f5e5tpXmSVi
pJj3juT3EWPp43xiE6HDApSbyShagg6MIag6GSFQN4t+8LYC11UGeZ6uIqEZl/vy06Udw+1jjZY7
O5TeEtLCmi8REY76Nc+onTZzGeqFlQRk2Dy3e6c853i3PsCBhiO62XE+RhBhkNokGw5cEklJZqci
hwIz0O5Lze0CaWkGcxHSt59Jvu+dfYVfrsoDvWLMIPkyjhOP4YX/5wqiHM4Se42Xw85OxHsoAVA4
JtwEJhHKitdpK0txausDSrOcWBTJ+DxxPiB2ksLHt7qY84TCXrObL0gjundIkZEvrtjw14oX6NiC
JTBrspqzXJWsrRwCUN7FfdmDp23OssU5fe/0XjJmNzUn1+p0f3tV0esxiaKr5RkW9yaQZjrOuJO1
Hf6XWjrwK+yzsm3FR7BuUtAtUbKp6BXy5unx/f6WWIUZTuB9sriu1vSN6u2Jlj5t0VnjHvVKttxT
vXdWkF0/SzPMSrYk4/wbtIG/6SDTuJU2z0bK0B3d1DtLxa0aV+0Fq6P6FaIrKIbTyMS7rIvcHqZk
MQ1iIzE7KKQhO0z6EGOmRLNpoYMxZg9cx90DOikQzm5060u2nYeyRMez2andlWSPpQv8rkYKRyqY
l9AZgPk2Q1ESdmL2K5r5LOXLpJf/6w48EMvZWye+H0oYdDJQgl2Mm9m/8qxSGUY7gAl0bCCnLVae
M6TKdr43I5nNee5sCMiOXwif6SGWjY3wvwxX0d7V5qlhGs/wQ3GRkfVeZZvqA2wLiW84byHgzJON
TM4+B3leNyK12f2bYniyZu5jGAjNbODq+XJpCJTHBXy0zDmucO/cWA+Zf+d6fDxvd8+GtEjQyxgk
uGPF2enrQoyu41/vEnLTaY1vCGfPYqb4iIeJt8b79uYbs/1S3zt6VwHbx+uLte4snoV9QaRm6m2K
0YaA1rmrSYF8DiMLV5kRjeEcdDUFUQGaU8urZ7+Aj4XX9XDfs/q9Y0cdKS3adtYLPJTIeO3FlBZ0
Tkx6p+r7MxkkAoogNjMKF6heVcxOgr/HnunjJNv7SY9oYKxhGnZI0CqRxLDSjjB7pdM/g4jLPjkp
FnEqpjM9sTdldYx3jJ88B5A5/lWXd3CvaDgQT1gNT11MVGxZ4iIUE166nO4r+UA/fKay6/Ok9S4q
6It9ViAXZ65aVNCa3MmTtKytQJIQvNDnrhT7O52oMwwWTiOFxf33OntS4tutBR4om3wgZpI1XViy
UGaxMXXgNjrLAqzFlQZOz8VF+cLOUI8sYmCikIKcqhsj4KROepk2IETkyr52rqjsRCN53f+9qEw8
02TLdjg72E9KrjP2IlAkojHHbwo912h0jh23hLmHfGBTehjtEtTKECq+hcvh5DelWL7hUE3zQZ7U
hAZuYpqLpwQ4oriF4uIO8tkxuGKEk3oxzZDdw/WUEn+KMIJ/rmK3RwJZIi4l6oV3vYg+T8O3P9MW
Vjs3vNU78ciU6dfwM4P7yowK8DfyWTFTXIVRFEc5X2OsS4X6ewDom6fE+pcoEWpHMqxi3MYIZ5KJ
G1AxICy1dzYh6X0IHHzEfsDVfQEX32JqdbXLR516l3F8CzzB6vOVykMROxqKYfGjc4S9mz6apgmk
f1PUqHw8eaLNyPcF7lrJqXsU9gQGhnd3bUbNaodJFS7PYyZcsirKms6FGcy5tVIlcnbaVmzIgw0B
t+PT4lTGCycQ/KyMwbr/cxfQfawU0y5qc2UH09Ao5odMe2OqIJerlJ0CCUJ9d+ro7PDRAD32oLmS
lndbwwmBDmquyhJKIO3dw1AZObTAe3kA67FgBLZyPG3lFpTNCOrS5GARHIj8m65KUgZShZnkKp3Z
3i5bU7eTGr5ZgaXl1uuNNPq6+Hx2IDBjtyBxIw1+jLtibQPuI6csKHBIcSfUrd/odVwiB5oREzkW
aV/H40GTB3Y+Tq2rU3htydLPZFKCagm+O6c3bqQUvIaPS0hGGsyUeWJGKvvJP/QmgmMFBdw9Y8JY
XdqCBC6bQfvZiGLn5AmV69cjQ+igXePg16nYEh0baxecq+M/F+a07pckHjE2PI0J5mlgD+v8Mr+q
NGumBnK+xNcD91ivtGe+vqL9T/3XydgJ2LynT1ygg8+ivcVu8PbOcY0+wIT+8SGY0aG0b3d2cJJW
vnPxfaGKhIDJx1FXn2Evu2JJuzB9S6TX7tqq7oQXZqgbol3cXNZ4p7jbRMtIS/f4sgS2TRxTsSu5
BGrqEaY9HCjqV4vW8Xt2VJZ1aZ+kwqV6pFK4AAfntgGlsjv9ozMB8L/5XRBUmlZk4oByPbAhQllV
jjWuOnifBIgqUCBgG77wPG2Vm58ospfanOmznYQeBOBSFMK386nMklDGDncPBWGVbHULqvQ0zRDR
XJSGeFpCCf2w5Rmo0i2OnPI6SO7wyRzn9wiOcSN6zjCCNDeoJi5RQlx3Iyz4LhyzSAHaEFMJYCRn
fChwK2Z4TdMGTDwNoFgkRy/5Frjg1Xrn9KoXi7EBn8krxUtN5N4rLku5gqY1Wo3t4q7wIfW6fo3l
88WKWxIU6yzVNaq6cx6CMClSRD2z+i6NPxsQvXXxdHWoA0xavjE2PO4pnhHNIPO1yoy+b8APZs14
QYZa9Y1WUU2L6EpQjzrvLimngk/bRCeoWqMxHfYVw1R8HjmP+aiQMT53mTWSF51e9HjeKTbyntgk
RCBnUU1Zcfjd5i6yAEow86VoTv6VWROtx9ns1aDB0pKfqfmE8dVaFz88Y8B5KY1M89dcGOqsy0/M
bbR8SH4bYiUCf3VAsRKA6AXekjtwU/+hCMZLJP9Z8R9J/ULsiXCDNCkJV2YQKDTmveoYSSz0imk2
/NR7Odk52UnWripdiDg+DagHqpu6zUz2f4JR9X5DWhmuY1rSLtfLRMnq+UgNk7g4gAUlRYVnGue/
mf0e+N+zFy3KMHFv+s+hBgBLuMLbI7J5q+8Z9X7DfxuPR8+ziYhUKphInmKwqo2JA16Tu28XG2lR
AGxOUDM5WW73FsCL6vKpzlu3oB0WFNRtsvokQ8n9WCfiVPR41I/KZPw8fkVQlnb3K86W3oBT/GUA
Qi6sYSvoOIfW0Fay6zD9IeUbem/yiO83ZMoqanwaibsDokoT8Io9WFhXNUonoTswx45LGf5jXM5a
SB6eXw4W1fo7VCHRsId2kWyHXLYZqQtNJcnYgH2YjW8z0QVN1jpCxVUpGIK6FUY868LVi1RVDnIR
tZW7UBDV+y8OS9E5jlxefQvOeL89LrHWlD0OpyUiZiFGowSDdtLLPlxHCY5MnmwgbLKGhUc5wSbv
3Up5VmThGTlmZswmla17ZXmlWEp9VDsQ8eHM0NvHrZAubEMO5jv/eUFJEneXgIoa7SiivxVandVU
DNr8EdtdEE1gPh6I1dzi4RZ7G3ojX6aLelhySBgxrwa3w2jCm6pBymHArAVLDy8qNs1hPHdZb+du
P+ACnnHZhfxCot8bSYrp05XnWNpe43ClJlSlaVbh7eZdgKXSxj4zJI6RGhfe3E5rLqezZXqKZtth
y3o/h7uwyY3Y7/xtSqf5ADqjBOQztqSqG7X4zkYDXA0wEzIFygeml6/PJ3U2M9U6B/9bjgBkVY1Z
IPyLW2YGsoa5R3ZGyjTLOdydLZ3gRXGaefokOI6QsegPr1PJ+773XrXb+OvntjEDYIqnQ8K8yfyt
uisH3RznMVf8cGICbE9Xc3w70LkRqXIhTmXshE90E3Ip2nurOOwV3P6khIJddG3FCaqleXreTLwy
zFzpbQYvslsmQhEirmD91sIbFkMMUih+rNjJ8Ulga086y4axP7QdQvHEGF0LYKIXehymAXNjpj4/
2podtOzBWSkY6TayT0GvLFDXh+9X02Q/Ohf3sALhgz/V1PpwxfoQnKdHUK4CBlnFcxvsmP0F4R2i
EHRDexb8NVaqM3skzUQBKI2/V+//hdZrKcE7ynY1QvbLn+se+VNNulTq44lpnjqKatsKp7C5Q+Jj
HPBpsaLCNWUoLF2E1d3XFrNEPaedoQJOkFRAj1az3pBWLwLdsjJJgY7VQi0BQmO0goF0753zeD9f
Tu2Ucj9bnhexaClfjPfOR2PI5Omze1YmEtknWuJgR9g17ItQ67EtZLTJP4PdXk9xqvDKQKfOPn7f
GipCqAxIHw+2QGHZhHsbb8GZgDl4vffVLP4ANCblXviamjCiaKXpx7t374dgryb3DULks5zDisQj
WI5oXttvgylqxRzCrh7R7bHeJQvRq6DlMGHBvtpeFmjxry08A801pJPHM84Mzz7+FvSJmHzUxrc7
BX0X0Lv6i+eRhDpJCCumQ9bbhvMyQwnufcdI4gQjOiCsYU1cSRfPNla3flAGMQZhKF8LZQ10delS
SGqSwuua8fcsQCipJ8YcnQxgdxeZKQE3zkex+So+DUANP86CdY5uzE0XYsAzcLpL5r8l8X+aQSbi
/AZvkISXHriG5nutvn3ZFABz9BAcw27/W0hNlYMZBh9rlNvWxGIvWKFQrUPeTPpnLmDGi+hUQpNL
xDkxEU1qUORFI/XWY0ohObk63bPSzx6QTI3ndIL90UD5sobDSxNKw3feFVvh+hr7Hrk6q5lsNwSw
v/eCaHyhC7qhHVGMV/WglvXLPO9JUIUAXvMDWBrAjI6jtUVL+jWoqcNYjZhyRWiAjwtD9t5nH8+l
AZCdDw9z4GKNnAK3whBY1dGF0Dwi3RtvB4rhLj8DqevFiD1ze4VgHhhLMWTiHPTKICncw9da6WtY
Jxhzwy5wF52jRsJAtD/pxDylBX9Hf5nlIzauwewqwi1yFHg3NliggU9yBI8DUOVMH/qI3CjzIHbb
EKswG//CCwMYrdrLqf54ffzjIzrt74+QE6HsUBfbKPWKiqH24dRWzKfIRdOojg7uVZ7F3f9Zkibp
KJTdQVY5FEKs0g3Y9Iw7Yn90liWvoK0QpS+j23G/Z15TbdhtKR2M9U97ok5qqplzkoeqivgY/kJE
AQV+jtIJRGHeOFZylaTCVWLr61/y51FLx5Y6pPIXBHqA4QjJ9el6f9OiNf7PdSTCbHu+N2p7bWJs
T40T1IOwtJ4EnQz7kPKuXkoMxxvvq+ZlQWuxtJkQfGZr8nbtetTgDbv0sqE+LLjL89k6Fy355dEX
hj1VvwHu5rW1n27z3531ryluBi3UPQyL01tdtlD5lfpWbzPQQOXFNwGAjO3W/lbljFhuRuvZBIJt
JpGCGdvyHWlZPYpD8iiRtxLMKsWUGSnN0ljMdqSX7MyRPIsoVmLUZgyTxi5gDweK5ipywxmDRwuO
CtEt0CdQ6QqG9TTnwwAB6QkrHSCQBELNPWOgJOWuCajeJzfjWpMHqM/NgVTOttZYdp2GqSqS4Nn9
iCWwgqctN8Adgk/fPz3T1wgk413HVi7+LvQ7O4bSBXtKXMQhnAI2AWvfUnzNPeXgKA7E7croGLST
nOgPf89/15hy5ihQg+1WQsz1/vpXp4gDco2uWG35bpNTN66x7PTwsM11LytyHwLS+qhSjaT+X/Ih
So3/fcoftcZ231or8v0cw+oJvoZOAGKLJdmuVayn8jeHtm5R06+NGAIxhxNZpCGl4xtW+U+wrhWr
BrVl4GW4sjbm/rAhl4VcLl+VAK14OgLNGyPQkPSvDmioKXaEZdGCW6ktb+kd7kssLCBjngsioW0D
4S1pw/WOk9wZSORqaM4r7WbSiDF8QcRjRz7sh9rlteRlD+1BnmtKvSTXN4wOXZAdoCUqE7osvZch
jJrCySrYPilSc9Wi4kLAytfMxB63yDYZrBVr8BI845/vzXGZzrOdKo5/H4cRVoHLiWdlZsCJlW7S
ee2aYoLI9PhsL4+0EBKW2KlfbxcBuuN+MUmraEbN+6SowxrbgY74cuc0kG2WuMgP7U8me0zkmP6U
OIVYrvVxa+bgl/LI4GDaEXXEuFNpoXtYKVO4R689yYitcMpWbujdx33z0s7OOn0aYVCCdRDb+U8n
hj7dtGoMFv1EWLLv3KhHtCtY8AY6WlU3tmMcmM0Zr4FuAULEn/QqltMoNumC2TJFJPkLyPNlWKEB
cOwR8lVhs+EYc0aXPu1F3R3X4KSfaRyi4TOzvxYLqHqLh3LK8nRRcNV6VzLvpzSBIFpuuxBKRM2X
rOezMGCyiEguIwAYA1ZWlhmf/8rQ0g+PXmWZ1YEiXgATTpHvAHelZIUCLqwxhzdZUaJSZ73Luq39
YXjYXObEnSRMUcjic1JcHM/BSXuWGJoCBdyTk8raeuoMfA2zRTXBJ0zIkMuL3sM75x6P16eU8d0l
/PH1Cp/BhyqkOVJfLGWsqbdo7g+PcFol0vugbl/rzMmm62eLOkBOYsVFk4Xx+bIv1Vl1QcTu5bIe
i0XcmRz2Qj83wZBP9GlYP99mM8fX1E4sxtW73H5J8siiZ5AxuKCAqGJrZEMXYnZ8sflpl/tLNYUU
TPKVxVmUwMZ/LPctDT8H/sSTNI8hRkD5r5tD63ZspT3ngr/Wqko01TXdoNKq6SMZBQc8Nqj32XGG
YDtLcy88O4EsayAZxZFrlE/Xh68nTwgZzSY/A4VdlX9fMx0zDvhNqjSQj/BFweZs7ymOv5nngSH9
VCLxn99m4KwwcLGtfQhbKMVxq95WiajEoCUorGMRy3v1URZqzYEnxCgJb59i4m1XIiX0UjUQN3lu
u/9ltXvWJZR73KS2+X44g0S9y1AcaXVapso2nmeo1xInfrwOAC2v4ArWOwBr4CcEC34LcJpmntSI
5JeJQghOENnHuSRXBQJbj+/iup3gcQYSIQmAKRlgY7b1Q6wydEhVFp0s7M2RjxM0vkX9mU95pgu3
1BPPN9jNsXFVDb7Rbpa4N2GGWx2L/PvQ8KIsl1fpBaP1/vnTBWWg/Tlv9mHP4cfBl4ZYeQt5Zn8x
zTRd3/4mjl7KWK6vHut0dlCPWhGsUrY/OKOhM/NH/nhWAIynoTSQ3iTaYy3CQcUnp9hEWoL6wRbi
Deii+9xMRW9S6M4urMkTiaXME84SMxPBFMdyD2uP6xTgjpmDbSXD/8Qy2QrGamxeslM1HM+ST5iR
CXlNAYyBzI4hYYGxcQUAaTczcIQHgUSdT+Jg/3uFVs/CShSc2R95+/EPgsTwYQUm84Evy/MFg8mm
91eWr/hHIVWdSXKjhuN+f4YNFZm8nUjjWFflECaX9p8GKl5dNmO0uQMDNG0CTSBix+GhKqxsmRh7
g1xDdJKzSbKwVXzU6YyH/gDSnMtlbUz17aTxbXnJSJUVX6Hir+M2fomwkdweL0hEPFKkqtLKFDn6
jU5QI2p9rpjgxnZvMxxKAJZPjihCcSPm2vkMC3I1NS1z4SIeu6pxAqbEHzlGF4w4iwElLyHLTLek
JAsp2xdFLaPCKir1dl0jCSCN8E824eeGJ6ncP7id0GuzbwacDlEbIcr+ZTmgaomreK9CfxagntIu
40YLr0RWMmQHYz7mwXGxR33yoBKIw17QbGdAfM0de3Dj/JSBB5y6Vmh6Vh/fIwKJQjgilCwA8uxl
N3JiFrn6RAOR8lhNr3YCYCu4J7bMAHLYQJLBhiIKs03IZzGQUM6yeS1WvdZF0wuQJ+/Bplstchnq
/X+FgFVjR5M/LPHUhTa9Czu2C2rsFpGy4sfdkZ8p2RXGSMCzOtPKsdE3qGipKR/NwkBnsKJPVyux
189L9zwJVQjH8Gzr6ZFqjOn9fEE1li7SI51SuJ9P+yjjocqXxAVuDfP9jAffnrgFvJd2WXzf7XLC
mO1De1HRqG7RdpwDqxWa2ong6WgJv6mWskdXMCwgQxFEIVjpHRH0+Zvjbrjso+0msEI23UdkYBXF
vowTqI3Y9YnwRo5OSULrxdh7itSC4CHJSxAKjPvWWtrYNua/wXJUVrWJmSUPJyB6CB4yG8Mh8Shf
2EzMq7BoIcee+ysUFl7cl4Ec8Y47Mesz38YpCRHYIsXN+EuyFNdZEDmylpUW5rztp3s6E0w28yc1
sjBAXqFMMhT6JbGBRKWW4Bgdqe/UazaMZjML0tEIGS6PaIYioyq5HJyPxSzgFF5tu+hdCkU7aCp5
IhhjsCgbnvRouZxImb1iHVUviq3EikdKq0a/PGQmYWonItrIBm9FgdvDn/wC4ZurDti/INLAnPvc
q+t5mbBZhTr/NqhciggeeHhUVg7ua3RCW040S6MZ7m67l8GUv0QKjFZG7Jnn6Nb96tvXHTJDqIjJ
XQ6w/tZ1fbpw/rZKoLi1QeXkKD6wph4Lp2DfgM2BkLmW/Nvgsnvup07yO4cJn/POY+J3TDdVcvFC
Tv7Dnf0zDebST80kd2RCZqh3FVcS6DlH6zwSSt6LLes7cu68IQeEG01UJSY4wAtkdEYlsqYDDMnx
ZQsfNaVG5+D0sSaKl5wO7/ZYNns/JNvGha2+KlweGUqHy9+fIzpRKV49qxVYNMDZ50mnWQ4d5pbK
9ZndhsNUzmEHjoOQTHeeyfeUk688r5mwL7xHdIKa3boVogNCznSWskVUou3ySFr3goYNlV+Njfcw
veYG+YAI1kkbmacUWb2GnQC3HZFpkW11+pNKwoQAG1j50lM6i6Zbc9DVpYffbjfnxf0dcPAHSmxU
Gg0Q11XIZIiafoUxxXQJroeAtDI8YSweLe/lMXV+NgqJspBzDkArjS4pDD7Qcnl02DOi7pCHD5k3
9opCfwyEIhsU6jZlThphkR4ouKNSC156t5IznBX/cY4atcuMYTgEwgyDz6b2+EXBXiW0lwceozXr
TgVbK6Kd4kH9ctXw51hEMCG0YF6rTPeJKOpFyyGsOiwl7h7rXnOBAJ92mb9Y+SJGETKDmCAm4OZV
VbdcqJXQ5JLV6V9THvuqRb17Zo+y62GRaGRMkJLHVTHHFLTqlb3kCUhZbSTcxy1suCSsOKuLOWaE
hzMgzqu1VMtBpDl95dGeM0tWqcZONR4RMqXVcjj7ClhZanx9SUiad9Q79IP3XW/meHtfRlf6mxfT
vW9bZ2TZRreF8Sqrvf0qlFQb+PqKGuW+QOTsoqa8sTdUcXWlQXcAMuGpAQFCe5/DCr1/sSZjxu5o
GsKr0cTzM01cw4OtZemHNbKwN/m0VwTPk6s3620dwXWCW90MYxcFBqmuqJ/c2GptMBkD0yC8E+Xt
169xLbPjBmUNqPX6AoWfSae3W1Bwlmb60z9P7Y/u63sjx3ZkgZbl3NVlOrQgz79eHMJRst9tQWGk
TbOHzUzQy4MIy0DYkGr2Wm92g2U1wl5B03981i05QsjNELphVpQwRdVc79lJ5MgFh51s56n3QfHl
zL/+wlkQUzxgXCy9ehgvlm+bf2PJwKCBjfL1A7i977RNl3mz6h2OKkxvEhKLcakPIA0dOpdgeHHi
dxGAagEk7l93U2zCOtvXf21OIURnRoYZ6rk77cEpwAETQFdbH38Y+xMpM+5OjqOw+Vv1f40BL/A/
vgq0tJ2ssWf2PL8PWX7p0EP5QsVQTYAZOiudgUzZD66GwsK7KgTEPjN6WSxxb16T2NLiHEuC3jfy
OoUEArST3kp2UXnoa3wnB8wp1TwIWnPbR2X+G0A5xntdS2ONZo1+YNaXBx9++A+5UAEMHD56/MuS
dFiTR4Ued7KtmuUGYU0AvmjGQpfBXIiBUFpacpXZZMWv/BQFiwEJKY8e3zOdeYru0lGRyiGyXqeY
7gjNYuA7/9H3TP5LIuIrsfXHO35ifuANkBolVo3HQGin9iwCTrsnD5ETatQNVQ09b/x5CcooPH4V
LpZpcsC7PasWcafzg4gqVQIYIV6Kg3jRwlhFM8iujeEQiMP6mpvqGbVSy1s/9CdQumW1+nU8XnlB
A1RcPLU/9G1dVv/TnNt+9PxUcLtnamSk9DDgoCvgtf4kqFlIL6x4qDLafckOccWzhR/BZPJ+lc3M
PrWgosobIJfal0QZUlewxaNEsI3OgGpBuP3L3dM1dyhYqmyE8j2sFpyA5++JfOye6thRgiDC8afR
wI5U4kDusGesuqucdUuF6Ee9ML2JaT/4jl9UZDm2lCFgaodi7X/E1sNRFlz95XEqGRmDJtYgfDj3
R/0yBCs/oDR7CYYmS4RmVXCh3gm0O+fJGVd7Sfez9Wl1TExF051RugijkaoREoFGZn6Ij0+m0ZkM
FBTffSh5TeHtj64VkO1cmR88i8tvmoSFq3Ugv84Dryn9bZGkDcJiHXpEkij52nBurXCLfrlIobc2
acKTVRE0G5h36QQoFXV/eUI9PVFQtqh6UHoP9KAiutmr7P+fx2COlnJwSZy4VTd5bZURWLam2usg
cWo9CQKhH7djsa3o2tjgmvA7esA+1+S/6iGzM0w6Gf5AyqFy139GunGtD3lPBuDik8kCtsDKX0gG
shCify5v2CZaxt1f+Kc9HPXt70XRKogVCazEVqw6F/McuiqMhv8rl2HtqK7AKN3iGGhxMd4W9DYd
JjId7hLhvGhUp9x3uTHRTKRmeeykff2W1qpEVJKkfl91FRXtYSVS/FVI5PDW1qkK71wdM0+Bytky
06IC4GvNe/6Fpc8jdnJShSv5qoitLwfDPwuNtKr078n7tZpSXbLxZbJN87vssHrOwez6vJqEpj+i
rKUz2ZTuhRjPH3OuGL/zCEzc+XlvSdXXCxyP/tlqq8ap2oAAJqeYYam3sEC7hMTHb3Dw3zED5zP3
9ZVx1qvm1LDxT9LVWsBXnNM5b0lPFM6OnRUi9yW8KP+BJZe+E2zRsrteseLachQkG4o9RWZVviFr
LC0fqxRe4ZtvFasVMc2gNzzkgRQDzbNDFhqjDOux4ERoNxgxBm28cREPuegRBH18Kw2gb20tN3A1
PNQ2Kp7qmXfnZ6Eq+ITKC7tDVhOOwm74jRRh878ouNS077H05TbZGoC8vX9ZCymTccAkxLDdgdFG
cGlU2DPb+Y5XgQFovUpZcZt4g/OuLWOPynS4EeeYPpLZZgF4PsjwVhY0knXT4yrWL+tbGUS0o0c8
7OHadD/8v+z9z2jawVWJjNknEX3yphKWHQ2Ep7xL6FfQj9My/5wqiIRo+k6xKhOYtkFG/nEI/XcE
0j1yB9P/guiEdGqeNj2a0Xg3ZyrnBgOAnPp/cmOi33MlV5SgbIXCDKO192+YdiyieKcTiOOuiBqR
CS594NMckzcVW5vxvbgGh+o3UbymgvmS0Bkvs67CnC00biHv6X1yJlNTtuPB+o+QQHX+g1tMOSyJ
izx6UGFaJ70cgRn0UrJ5ct00qmJQ3a1VjcNaSuJqWsiUcRPXGV6csrKQ8+EviKkpnhdu8KxYvur1
Og8XcyFWEOlxz//K1v0CrpgKxtOSxmNsaeEq/ZHBBcedXr6H9x+fxxC+vq8ipIIvhc0QwNl0SJzz
z9TdQe0SLSjVEszhkj6oYaHr2F3CMs3fQMU6vmN3VE3EnREz4TnIox62q0StIRuA5SvqPqPCFn1s
7BUiGrY8HQcQl5sbNwN59OWlzsc5kmRV4Kl4HLYncP1+cl1KxSOaY91AHkqQrFpLbdHjxteULD/I
fZcSJx+2kINQX49QZNY4ht/xvf/gdRpk315zGYrKUrvWU6bvauaUwqTDdqEVZxF8GL8oYjRahHYJ
GHxLt276m7VhfWZzp8l9VSyTdrd5CPJeYI+o21pB5RIDHJSQ32gdMmTs+BKEKwRedFepoGCksQio
XZpBRVtBWqPOU3C28QwVLoS3oFeOPE4fVexAN+dPNvWfLBQH6vHV4UNu44wuAET3/j80k6aTfq56
CZMZylo4vfuG6L/oYnoNb7Wt3ObiCf3AeJ0rvZSuUoPw/KyJJ5ahdZygULBnTix4dUtNGW72cxbw
gRRgsxWWAnGm5avDyQvJibFjjA5ePDuQl93oemfHW4t3aF6dWdPQIDbi+siRm+kNTlGxv0S0L6JF
9VWsVPv8zDz2bpWgF0X4k4xHxQo5ypRmuLe3gk1tl/DLmLtNebtnGwwSBp0PQA8niYBkcHtCd3wQ
YlgEymmHil1nW+Lsiwdrxd8vRJontq7AVhYItCG+pmTHGkokM7OhAsNi0gknhvCU34TCOLR+jw6X
9agAzoPJHrVt1bgzXIUZP3/qPt1L6cq6ceFRNKTzswakofZHlX3J+2NYUC6g4hPQrgcEfQzbxgtY
quBFIRPRUoU33MSlZa108bAH77ggysgoZYyu8VO3lUvmJP898kf8TydN076A/qd+RzXYlE0i9V/m
KP8EhH+mqHq3CB1UKPoW05IqxuDNmcp+KzlCT4xeho0y7tiUx59oSv9bkf80sKAafMsIeeYTJ+r4
p494vsTZp8OSYbDyu/KvpDD195yY14aDjbGfJxrsreLIWTOnXRWmDav9gzAsAliG8BhXjlsk8Oye
Lkzo3yVWmfKBHxOMepQkSZ6R5MIM/JFu7WR83gDuByvpITZrXekn4FzD87aHDBxD0URU9yg01/sB
hGiTuE2GQWG2W7ZCarCEUDEHap4rxqYtXRX1p/znrKW55TPjH+GZqNRkpZhotJMp/IlYpq4QXofq
y7nbWEZS3rC1TfFOM6NmeNfnjsx+/+0odYcHiTkP03m+S4OOmkng6FsLWPFgorE2l15jIqGmWOwJ
ifqCMbb+uEzStN+jG09g9QTFNIdeEK5xvqj8azmOuErpGGFTb0KA4L6c0cjbhBplb/iqba7T8QX9
ISjHtNImWFaUS2XQaxgo6TTVKuYaazxpz8GUQ+qmbkCWCMmAI6R6ZJGkS1OpXxUF7HQqbYS2pYpd
b/d36C2j2EcA/u6T5SMwkd3CRKaDnuThmRRdLQFC6lYYtCxyevKHHcauBadD/DtQzoWUclNOWhnL
8wWurjq0rTw1u4Ki0xFkp5eSI3nsVoFtDikA42+4jaxG1czQXsNw3Xq1LmC2a++Z0XJDQkWivTyA
6APrdC+WNix+DzcVMAMZxEv2IYJvJsnxrdIBhsW1cy8cSv3KJbcFnapeY1iDYJpbf5E3eRCY69+o
DICnMYCyZKn5Qf7u4m7uBrGyt+snF/WoeC8oLuTj6RlaLc7FGa4Q7wwwcucPMCQ7zDSH1jTQkTEV
AH5BXPW3qlhaz2fhR1U8zORQfqxkraamqM6k3ynse61oCX9uoVAxQIPP86kE/PzSegx/nmpcfKzv
FwJsfAVIelNnavzsDaEhJgOaXCneYPyQkbt9/vpwC0ZRdeHKXI/3USKblSsCXB06XD5TFz8ZPXZ9
YjgqY0GvD33Jtunb+du1qWY/7XJ31hJD54WAuvMsWIIsTt2u4F2qn3rgE9IjBiU2U6C3OohyTswl
p54fLaUrIIsgFR0Ggx+nHqR9cLmkyWDHiwAiJiY26xmjKDy9V0xp6Y8uhtw+ULtix5RQXtQgn5pN
pS2p5pyFlTjvolH0d4y7uW9+JjCrA1zOFn5pjoLRYK1C5lJKwccHDudesdD2D/Ql2NcnFM+oTwav
NRh1i0ydgMPWjEz+IeyHGtW+tqXYgEXiqa5Ug2fiSF+Kg1mIVhW2ZUmPZNZKaNjWk4AVjKvmbABE
I7E+dvkARS7t+5bSvzEJW/c9cp6ScP9FXH4CscSxQHnGjQOq4cz/kRREoqtdlmYIFR3e0OYDkJfu
p7XcLC+JqeU7Z6QoiTUvmCRoHcWOSk4t8DaWt1B4huMAWQ6lGVe8Yy5qrUe3aYjAfQ0ADatMFW+K
e5Xco/WZ9YqRRUvMzB3gRIVpQ/o+2d/syWMnO3LzItZiozDGB6qP6f9iwhACHMf1iuEBEq5T7ekz
4zgerllcDE3SeZgbrHo7flbBI2N7XUhOHbPmF+5IFxk7gJZLQOJkFjSu1KJ07KMYVkXrE3vtXETL
axfvqreVkX2P4kYWVcJWEKbv+kg31t0PmUL/zFwGAARfq3g1vxikqdqLyKQYy76qOyqyT+u98oGk
3BA5pbX7m+2YNJsU2L5A4CbHdsLmTZau4RpacgNfriSZuTbVvf+wdq/NTzsTmupXXhWFinzM1HCm
wlXj29U+ZgeKkqPnrsdEXnQXfKg1TV/g118IlpdhC/yUDcnSrCrRRjguEad/ApOa9EyAKULPrsH2
+YTt/jKJsjW9pWe4atmRf4q5Ubv08cQNQHzCMQkjCxvuLfYO81ycD6oT62MkUP18SYwfjV5z1kxp
cGNaosj/VTd4A3+xwxIkDCwgQX27CESoWae1EhMc1UQBeZYiPHrrVPIJrdtMnPs24FT/WgDt67Vi
7SbMe4iR7r6H13OcVw9pt96XSZZID6ilMQYgZcepcXFmL6/9/n3QgLwzqJjMA8o4vusM73beYYLn
ptyfFEdOosdFSGV1YuTYmhr4SvmPR7OYG9XLWN1F8T/F5A4v0bBVphLXgMoTQO3vaf13YnFehyz3
U/4YcUB/08OpzmU37f+abR5uW1lOJ7ya9VackjoviGLBfezgAWBW/47bArCmeZJxro635YmMsvn0
j79p89j7/kqyaalAsydDdcmvZ/ETic9Ilmn9sQLLx/25L+JxJBKUJHpPMO0RSZVqVw3STPiiKh3E
XeU5kOJ+lnWE/Ib+atuYHRF7eHsprEhwtQNlkzuVDu0dMglLLcQxMnPE4QDZZcPuefdFOOJztLw6
NozZtZAXVcnxj6XQtDbTHw5yozrgtUeHD4v+ajc1KUTLOpX1udjSrDHE9Lxi+yjZROdg6Wbgv7fA
WklaCYxwsdeAlzzgCS/QSRZQM5J6hb6BnFyXktBQJu20Z7WREroYs0hA2KbtDc2jmQ4tvYSjyBDn
VGXcmbUvtaZZ9HEW6KM7h/ztGwIrSM2cnis+pI3JeDF+isFVVg2i9y3TShAMwyFaAAsZewCVv7q6
BTZ98l10fn3ICETNCE1kdlTqe2LA+oL6EH2xVWGzneM2KX+uKAl2lo1jFa5SHp0SmxewdSQCClbN
xhea+pjaHOvNOeT0KCe11XtjNi5QmaO0nLwylgChyZ+2+fWTDVO/Ll2j4gS3WurZ10eAnqPNZJO3
Sq7GZTc7JxhNAcPyiMsEqXdf9oENOmp6hXvXcy4f+FxCAJdIWxQ3gYUpgpimYFvU1Ai4BzWOdJY6
Qn1FvNWsvskd9hOyUA6BDdE573fvBexyY/NrjdmiDCyIri5X12L9XxljTjtB0wXukZiwFe83eajv
GXSpKxr1J9M+StgGqt9w2tSDyUKsSH7r6O3QFx4xlc9nRJdLD1jKmjTqfZ49RlOqbnRNZCtBqRa8
RMyY4RZEHdXNHfou3YQiUla6CaA7N8Yp2uWJDNnJ40WyXMq/FSCujvGUBvTgll/wAQh19jIwYFHA
mKTcTx6JG2NAl+yA7HZfuXyQXRvztpPMGIFHo9l1rkgxqyhXck1qW6YOiDUEiSM1WcIgHT3MlF+O
3Ed9ElOceYjPqxxkLOCTA8yUd4rz03QyX4l2o/qkUUzv5hFx/POhuQSlAVIn0GbK32gScb+leWF+
IUfl1y55g0SrIewjWfv+3WJk/VeOJ+Zt81vhUVlIJDzM7TzShIe+2RD3Shkg7jBdvwp4N4gUMku3
6cpZFW0L4gCZGKyz0XOHMY+Myo7CWaj+T+4kQwpW4c1l7SAkG8vPdkzmcMPgg3BzIYmKJRwSFmfk
GLy2QsO7jP7gZ9bDicDaoTa/S6qH+G/rGXjoxMwODI74F5LxdV/CiHd7StF8M1/qyjb7j6mkt6ua
qkq9qabNuIXE+t/QWf2WZenxmLqP2ljQyyF3s9Ys40+GLhyqUQKaVxbffAAQdHNk2XpQWN3jHm1t
caYrRKu+1DAGGuaVXNdXBttuWRIFFQAp6XRv2BZvrkdWr9ofO4BOInGiaoCXz0gyVLMYMgsOyMwp
eCO/nvdilzHnzpLhOz2JeGZhQ36161cFtYOb8+uVdlxFhhvMrImctIPCegBp0Oxie0l3yt4lLaSz
HwsCxzAjjeFCF+PIv2qg7a7LiJp6u08XrjK7VHcTUnIBIdXHqYrSCxz7zB2xP3tyvDTMvyrvpVOV
4qVMB8M8dpPSHohlxa1fIUUTNYyAbvsK3vyKT+WKRVzJlWoM6SzvtpBhjByYCTkE8M/Bz7BSdFKp
H0U7QfpZ53ep+PFOIiZ//JMda4bjIszr2UqQxxG6Cd+o6n8ilzmhosLzPtkJ4RkB2iuah1d00xMX
8jrE7N0iEdby1TeRGsZlFBI69mWoID46ViLnzhpP9aJHZf/famdWeI0/Tqs9ihufeDpVpIijwesQ
AjO5vY6/rF2jDTkpTGh+jQHevL+K2HZGI8e35+txgJxe5MWXCoi78mfg7wCAwnbexryxt3MbbWfn
r2CEaEY3spva5oZJJH3c8b13af2ozUlSQaqOxxeFQZMRSrGP7G3Ycx2ZwB5liAJ3pykE/NcE/oJj
WKpgONDu8IONxilVzV8f31uUnqDWsrfSWLjlRsTgUeP3lwiadGZMcGgIJteysIhbb6fKRPvF0ops
E4x4zvYytaNpoIkOlDsKhPYhTgn2iSI/E+GxpAvDjEsBNZDjeks3LMwlBuafGiwALTRRJzhIHUvf
CA+IRe+rllmYzIEGL8IBNW7bUjLQjbsFJt89tDIFGC+ivvulwar/ecyBgmseiXe2Z1rDrB5wX4EK
HHrX+sJ7psAJ3v1nQ5Ek63gXGf/vJ139dSryRK5y5SNZbzOsbIdvxEBG0WOLToG41LH34YpQm958
F0jv3xSs5JzkxRw1DNgC/72OUZWV1ve2q6F0Je7had/kmD3d44v0CMuucOZBwzXPE54Uz2BKv+ex
6mhavaaTNlMp8NFn+JllkXBv12nlwm+8CeeOu73jmR7og84oVxWQ/I3WNvGQ09HdABJUAPHuOmR/
cQur7UlmHz6vHOfj+9QxbikJ2acjlSG1P1a+yrd2BhIICEodITWR6coWtH+eDUa7E49h5FSvmQpT
UhoWpKm0j8Yt7UpoQdm/HHuuGKJ/TvjKlxlQbbxwXaYTk/YuhRN2cc4pdWrKZZyiF46iJjTo9qSp
YJWm7E2IA9Oioii8NCaeq4CMjR5eOpgV/b0kkGurlGVcXep5lBcuTJfsW2ZBHDJbmjZ9+XEFR5h4
OEy1OPrVr35DyAzVLwwqwsQpXEZ4rWG1JN9U6OJDQ70tl8r173PWy8iL+O8TsyNFDWaHda87ZZY/
py/0OstRIkaAF5AUTOn/PMJCl4jlmQWWj1SNWzNO+4vCgpcvPXCsbyj9GZdytM3hYiwcAgWQVF4/
e1KAqR/dCusZ5bRl2Ajr3r1vqmODOzEbpUJNAEOgCirg1UvlZyrNugb7/MxEZqALOZDSsWtQXWMM
0Q6ZgTTXqmtmdFIcfMtYnSg23JzUAyKP1p9QS+5AjvVTHzcm6OijAyH4u9DW9E6smnnIWZz22V7M
QtMpd+3nl30HJaW3eul9Tzjmacxa9eAqRqXGaqd86UfKLz7TVcQHAJ/7RUnTRhf4myryGe4Q8ssV
b2Q/htJhKJaJVZKJvTvNK/CdtdpBKOkTM/mAy6AqQNY9C4414sh5s7/Z6URLIES5hnM5NOmG7oGb
Glpeuh5F6QAa+SGa1hNdmOXj8fMj3nG8ZIhE10tp/lRpHWefA2sqiUNzPP/Qob0LHavZQQ9P+oH2
QGNBAA+lNvKHCIFJOHmKeVSmR6gDvZdjBIV0QrP1TI1gdCuOrH4qJ5sO6gpSF5dnauIc+6ry0ql4
BwRu/5I6yQ23m7pjidO0WZVK4EfrL8mInfsw1pQNoJSXKH4fC8RNbPiAfiG4sMOXvQtjw7vBT3/Q
5AWp+L7NdCw/mxYNTO3NO8K32hsvASxHDhYMROym6Ctbm4hwX7fiIjmePS/oRs/2Jpsf9DVEKRD4
3/erJUSruxsKLisjAFB9A3hkDoEipOtWIdv4VXO7yt6JnGtDe0iROn975dqEpplH9y4QWS7wDv3M
pXfY+j/VNpsegTIVGP+1O/+ssgaqoqFCB+mKfQCjxWVFu8IL5PFWd3KfmA0dKp/epp3Ksu9Wj48H
/LrctRnB2WgyAn5FQM6vyPc76oRq89OpjaLHgt8rQmqvq5sOQ77ULTHr5NGKH7xjfU4dZ3pSxKFU
BvW77hfIuvGY+747Wg1EEacEPKi2rnzbwyNkdI/72fLUBZMriTbKqtP+dRtbApVYgRZLDeGjwPrC
7M/vOQ4RbIE3ynK94gwApx1sDeb3hAoUucELsCWnA1mQnYCrF/BFhMIoNCKkpG7Ln3x/q2aAZHTo
6KaMtw7rizHqFRMPy8L4vxyJpOL67JATHQAb3zKZQNXLSpKIEYQv9rpZQnqtwOC/q94romlbymHY
799BVWzViz4g5qhMLJA6scQ9venGMEAkT4DNRvTOqwb5STAdnmM6oxxwLW+0WkI+kAVEmC5XiW9j
tK1mi6rqyfnOq8RC/bsqqDh3CSOp6mPzL0HJF+qoOMk6RE0kRuDQcqFtkfFQpyvSmyt+NM5fRjq6
8isJ7EoU1eZ89xg6WHRX8gE9so5u7seUupJ0ti4uuikv28wmF7uJBeR0RKurvp5OK0HS4Xws9G3G
YvXZDj6ILOLECPplqNdqOiL0WD8sXwsV/gGbG1X99YixeYYwIRFuRkpaRZxutTjFyGcupzAKsFap
QmcaYeQdTVvxOH2+HMqW5oWPXun0kM74EXFvOeYgwgmS2hWLLaGkTD2l7Y03wyrgvlSvAXKkByZl
34+zw8+oYeezox5LVmqZn9cJvYRe7J3/ZOdbCDQmwbgkolib3yE2ZTDVCj2j+hASzhLERH/698eQ
6JgsQrDR/mgPrT4vu3xiKy2c9cR6eFUgRJHZ5aSfbLiLvIo7LvalArswWXfEd1w+EXebD6pdVd6a
AYBlkpJImbsX7uotWGOz4uDlkFU2PlUoMdoSgaHKgFEGwecrZQTN0vbE4/E706P6Bex70qbovIU2
0EcPxyIEpZtbG39w7qovGIjx/zQxqiqYZVUIyzdoI74LWe9Rg7CxyXC9OuSXUm8CnGyC9myoxCpX
hQRXyxsh6wW4o+YRMjKA6WhU/80fsDNwRS3c8qLKCoSYFtOMfzyFWn5o9nGlmPYqvCmtVMj2Fk67
dFS3xP/FTKXRwsfhEXAXUe2Tw9xNaHrQqzU79hg5fnfpse2dL9+WMEYiilCSAX+vhqLWilzkwtI8
H7aWXP8QVT2bPug0PgIBHfCUkLlMoLemWa8t3MlemLz0Dh7Zu2dMyOuvRK4CvFW051T73QrgIPjP
s0XYLTE7gSYswATro68mTGplZkhyZhG+Z+KGw479R7Zs8QYvFS5WWZAIXvKQkLPq4yo0gaPjvR26
QLb9ndSUyZ4XWzqzh/9airHD0/vAFJavj15dhczXp7OSMLfmxl4+JE5UKQM2Ts83EW+jEofXEdJR
hvivZERwhyS1iVlzrKhOzvyWcdE85Y+2c9yO8kCItEPRbzu8ecCPq/Wcdehe63tUD+UnLyMnWDXL
U8mzDTsXaKHTHIaCOG9Opj8JD5qUBlx2Xz4yavYBGLs3JaQyXhA7Yw1UoobyPOWfRJNQRQqTX4iS
g+++Ro8z9iYmzKBYGBRUvIxhT3d4HVK/45THRv1sNLka8GF8Z9RhHpvaTj4hAwnX54HBWYJ5oG++
V1+rroMbBl8+hOv4936Npbfa5YiAZvjaghGcj/kf/NIC8k4fa4LvCkl1E2iCPVShrlZp7wl2K7MU
T/iPI91yJfmQhSgbGHy8z1l/bQSsPMY5K+2Ezm07RGSsEQ1LK6v4Lp3hJGR/KyKsri5vhWH8AMGD
pqbm+J56LzGxHW9IogQAGCxTn/esyHRLItqa/irR9jSKkY1Dd8OVHNOkTdta0pJ5gCpBSCDUWzi1
xdGSkcGNDBWcqjejFXs8nEGuvxlL9vu2Vk9/zhnkEFqdJeRFINEaBLYvGDcCof3DOpTug3SUiLs1
VxVZagKd/74R02LEiFgnAe6Gfyp6uTYS2FPr7HXo2WGviwpgPcgsLlFGi1e+0c7aEqpWh1fBxtEb
G8velxixe8qkMJRl9P5vmF4Apk82fArc6FUUz5MgLtfumutIvKpDgnTMMHZ3RdrRFJB+53Bsd4rp
GntYhdbVFx4uzEjXpRYOc5ZwLChYI7qVxPWCQCKl2gOWX9CgDrY+wJjpCS1qwzGNYvstauHVwTWe
6A4Vz6PsDcZFiW174MCV7g/GVkn5WhHNQfDGSneYKxLUlMlqOS1tGvqbSKTNrlo4jkBgzGkUIMka
FBMp10CeCYjSBcqCLiUqZlMmgNInVBF8EjMGYyJi9xfoYqhpGJ939ujHxuInKJ53uzp+rAKS4cUO
vflRDTLebZV69q09jb3uTFtNcRg9X/Lfv8f6A48uYzv23k8NiAiOYHIlcwOMxNNq49B9AZujhh+J
6T4ywlMkfgBLjBcYY2sKFNhSRMO/Wo62aa+oZ7NWtcyS4k8OPXNA+3UOVWS80uVIlviq8M9fh1Yw
oA7rrFeEKc9nrxy7V9XWSpH1eCwp7QsfAGS5Wnk/jOoseuul8+t6OEPLjIQ2AL4M7cn1TAuksY79
v0C2hGawI4P8+0x5JAgkzSMhUfx1ERyo7e1S0gzNacsjDZGtbayDdzGdOCohXci03DJeY1AEOuIS
cpA3ThyHZZwgFMiZJVWAlClUSpnUQwGVe8ADnFjrWIAKDTDXfeESrE7m6VQVdxMNdTHn/LzU5jYS
FqsUnBgav9NCqsFULobp1myC9HaZ92TpxJohU5zxzwfg4weEX8sUDPRnAARYlAgz2MNnaRBvjQWT
9QdAl0/HXQ1hiZt0yHGhgof0bLI/xIq8bCXBolZGoBsD0unzXwdO89aB+m4eaofHtsCB8Q7mwq8G
ng9kZ+3DnfFrsFMqDuVAujtHkDTqCmIjkzLTrcx067e3ijrMKRvrn82k8MAcN4ZOp6V997fpIJ1h
heXHUZaem7DsMnXc2qD+FrgsEBAyy2qYdq09WAtYvq2s78kntGm14zTemGmOHvfc/oBnkkETOf90
wypg7dm2C9GMdfZygW9XNS7BhKopk0n7cmnxzdMSDaKEzt7LkA6ifS6u5QmfFSFHzCSdtYUJit5n
UVIxpM8xK/8OODxo5hgsg6O9lbS7LXeLR0kyKVWhjZ9Nja80WUcCWZ8UqaGfFW14S8kSWJX4WLO1
9fGed6YCovS9pBdjNjT50b0O2uH1c6cs1FfajYOZbkZTL2kVOBXEpW/Qd4UkDWcEp5TK5a7mMgMh
7Kf1SlkxWZomTda2egUiwteXhV7+UqkV+pb1rg5uyZMcQqnVchsNV5Pjl73Tl4OMzxZ8QyttfVWX
c0DGRwSDHMAhcFpFDEA0ecelo700L1MgDz0brC5xvHGgLWf/fI8MOwpyNOaRagfdE/Kq2D/SoXaJ
SB1obHIJWO2bUNWnncuQ42amWa5rUrEloXomSrZeAZirkJyC61CxNxyewBpHrnusDHae6ERMnbrP
bfQJJ/JpkNhPt9uj0Fh7TdMnRDr4l9rf3rUL9FCFV9VDxX2IK3igMQS7AXzbIyf23uVi+0ny8b4W
5Od84fD1HmOxUeYMSDWwcGJWUY+BkYko4QbeJm5bR56uLJ2pa7X7bOYVDG+mc4a6kB/fC+6a/CQi
Kj7zDtGMnMASBjMYxNqMRN8hPofPt6EbALeUhU4/W+L5AIyrhz51p4jH/DAfDYf73V+XfQV57TRR
jOUloqFbjW5X1xWKlzu8ZEbM7p0k6cQogLqwCjUc6UtIe+0h1H3TkEC5678MGxhbHm1nXmKmxA6W
VmCOt5ET2BL1ZiKs/JLvs81oKP3K45QTMWeZ/XoeYWYhhMynd827kRP3gMmuFAz8pcWW7q4Alwvl
iTkCOnjqUoCq8lCoz5uAKJbSpoY/JfIB45by1JHDKjWs/XT8wigEKqE94IETEkqoPa7srvBypBHd
wIwLaZTwrdOZuE1M3o/Otf/YKku4fLvjHHmNYZ0hVy91O6PLYH1Ivdxp46oa0wzScBuaacK1sb0N
OELINQ0ZDS8n5+T23frUkJI3/CE7EKpq3mWiOjVJLlKOCkoNcIeQeyCuzFDDQRYchWFfY5E4Zx6v
IWxKozbAI5uHhnpf7FvvEaC9C6nl6Y4C/HVm/aY5hkZowpiT9kC+40Yd4ZjWLoDoNykpyOC1UYGm
Ft8UGaNq7T5RWcO20EwfX2jol5vmRAdYmb0SHoxXtGWA5D4Taei62YiDdidP9DQM1iIOmPS8nrbn
KdAloYJR3jEKKcLTBqMioVGOohJKxFEKMKGwdHa6pqlcPQIVY0YBUxRWW36JpC74bLs0R240QRh+
j0yp+j49FDHJnYg9ZvyF4Gg55Vnr9HXwnBujtZy887B3gEbxTbU9E1KRQDGrxgA5zNBbOsd+HeSM
s0sFrb5ostcPANRDMqxkVjDnvogjriLTHU96FnW82h6MmKifKH3W1kYiMg8ZhS/0mVUhj9w2QVGF
zUdlYlEQEqqZTa9uGkuXrIGXa6/+2dVuKBKHFMxQ5hF5BKwKLdR6mZNO09qoMKxV6rYyz3EK5Wov
8H6+Wgl/1neJksYh678gtxX37M0ZVrnVHSGx7+zts1EMma0T05ECxMp0gO+DYMMq2cCRdx0NEprw
2qfdzzafcBelSzK/JSUKMZgZ5ET4b4GoOV/ZTD01mYmDaPVpzLlfZsH0Qum6Gd6PdziCMgdDaumY
nP/sut1fH/byrblZoRhfwNBlF6kc/uobq2sNLod3gkuIR54GzZ0NqCOfziDgax6sJt31jh8uohMy
OOu+M0USRrhVcq+oU5KK4wJHSuYmC/Htp4nPJlZkVvB6MUl3vo3/MfY617huYIJ0kF/mzYfCx+DW
Os2X0PCKvQpXOKNysdZRJWsjM09ZmBXXKIFzjhkXYFQbrdj7EpU4engw3rygNBvIl72jBnm2TpTm
4pnyzl3FxjuwGHsNQ7c2HTRCz0hRZT9aqav7IWZxOTTZSqEMP+DDnko4TndceGA6y/3VrBDxDNxS
xqmjjMk1BuH7VNu0EDhWQhjTkdPfHXGlu8mOPhtH/unMWizRurVvKqdINIJyZCJyBjuUo3VCQbto
zIgaFRHfrcTkkFBMY8BYEqVcam9m4V0Ts9dm0G3TQFaTLWPxylgHhzAW6Lq6sWOcdTWE5gVV+MrG
8pkh8dMAnr/5JsFtKqzg5CC0R3j3HwNV3NXLTIigt57TlN8QGlnJfyTkTfH7BwiiSqkkcZETTKHP
ttzZmv7/egu7ZxtdML2IRPGwONFqPP0qzHVZtcizZYY0xWldzzWtWQLd8Zlzp0gk6FWdJX1Nd6Vv
9weYwo9QOmvl71i4GT5IfKeMrF5CbTEPwPNJr1BnJiIyfsEq2Y5O27KIBa4ZJIghPH696np2mdFD
guRPe/9mEfy7/I7KL2rCvsbwiMja71M9+xxrYOhJvIuuW9KSrXGCYoD6oPlzUWpT3QbMNejRE/nu
hOBeoPrt4a9JnzwBaDqYdXF2Z/MKGuCdOwlEqBx+yb0ts5ZjygfdzyvJexSA/VknH0RpHvFqSGm/
w55yKl+FR+0TIwFt9amGU7asVZM1xLgFH4x9/C2gwySU/yDwRI7Mt9NWkh/Ybvpch5lv7PTDsm4K
o8kBmUdfhKSZOeuiUOaydHMQsWrJOH0ifmrhF3CO5tKDekDQmOKsGcSVs2537Q5EqNR+l3J6Lu1R
nyyfVQnbNVOLVzfItYazvlceyJgiPBilcLUVWqMYvgdVcy8QA6kDwCkuczORTmCmKD0gUEq57wFG
F1bAiDMbRUlxqvlUk444SdzyuGo0n+HLjimd1648V6lmHgA53UvYX9yJqAWk3UJzG24FTipIVMOh
+6hq2RoL2lGptD2RCxnCHrPdWjnAK4+7rbmY0Ws8bYsLbL87iGmhHBHRI+7oLxwjIBeZ072GbWFk
tOTo/6bnY2iZIrMGVbh/+8AVXfAeyUWo8jbDANokEUk9Th/+dchQg5jsgp1ZN3h+A24UCBrYsy9N
x2pCv5zFlNMfKJ8KC2dwSHw4Pn727/W9azb1m0wN0HC1CzDBtdBLHHXg4IhgzC34KfPYUPqKhEbm
SOj8Onu653nJkhGoXFft6FheL9y1yPfgXzf5DwIRZrNFQS5Vp7t3oWUgiZqERyHTnsv7o4KqAZ0i
9llQB9STuhkDj45r8O8wd9hSpgYHBr4IvnEnTlTW+9BzNNpDuxwKIsfPOnPx0VNKk0RsI9SSfuLN
fhDs/9ZnvPJY2nUyh/qOC5iBYCfSUJSCJxRkw0WKszu0ufMuR+xaHXhEEb61kiei4sXqNiKfN3w9
W2wMUcFStaHTv8UN48Ff3qjLPteKYm1sDIpadVqRoA2KhZutExp/bzlUv0U5MjwL+WJwOUCftMxd
37vBx/cYfVc3rtqBthnYwp3E10Q7i9i9pQedwlpG3/fpeYieVTe/uPnWMIyEPRHTirvH2dpvrqIK
nj26CzWEynJq6Af/SXxqn+oX30986esnxdgE/XkDWbux/l7nFRPU6wVW0+eIO9N7wohWzoCCw2u1
m7aWYw3VBgHOUHT1WBeCgDfhbQvs3NLFJYAMyB8rCGtLpmaFxbNgvVz5IgVuFNNRlXUqlq5PeKpt
48xo8/6NwhW2pl0g87AspWAAAXppAfIT4p+X1MVE+dzcfeNAajFXKeRFyrzAJZkwsafCPdkVdfc2
Mvrw7SZ7Lax6zxp2UtHu4SxqsCfHFGfanoq1JAz+19YupcpQpBPYbIEtOPOZiTQn3/jg3U1X1JBm
S0w4nFHQ5ry6TnPc858c1GpTyZ7d0nFG2SuVt7N56YcOGq9wfZMKKbXzKIv9fVHRxnTWIwpkQ/ut
FN7hsOfWjDxYke0aVD4SYTamGv3slE+Uz63drSOnP6d/N03yJAJ13d6ccmj2wL/r6uJDwC65kJJ7
5NBRZNf8oDT6qzL86+qurRbN+ocY7mWwO5LB1SDU1+vHKx/AgIFcaU80UPgqdUQlbwANFE88f/kw
6yZqxnZwJLYqH+SxAPUXBLXWUSRyg9LvMAP4zVlFlX2UqdG8V2koYf2tfbdtfA42SxVuNBwgcGuS
O0hiVleo0c5WGXWQwEEMkD97wFIYxi08QbQ6vh+zv3OtlZrDtwMHpFPU5wSRKCzdnTawrxx2X/co
AkMrs/PnlacI+GFcsHuD7aha28OS+nA67tudeiiPnDgQCI3wVj0xkjBZH/51DoOyTF/ZI/pDeLqS
vuVx6KQ/zqxrf7QEJo3+xbyaX/CC4mBFsc9Q3O7LhJlngUlrin6p2jrvYLRL620rKDavLuvdeBl/
o8EFqVe9ieOICduxsqfKukVFQ4CtM2phMYQbN7oDyMVduLNxXS55lmTcHwgxCFo3+B25Sywzkotj
Vz9vrEhFEGsIclVFqB9fxcfm5KwPeM9Rea4SGY6QdZ781DVDt57PGn9GVkG9Gs2EQZU0sIbJLiEL
7t/uwieeZajKYvKMWMcUHApwlCGq4EEU0vf84Fp9iX0geYXoLs4Skaha9hCRZNM+4nWocMapca2B
et8nCvb3aM6MxoDOorBDPXfOlzdF2cw/9mSvKXQohFeQ7nHxQy+YDgSx8yF1aV26R7pxKKxCZnGn
4urvRlhpfcktyiUvTz0xz8e0FNDchUDPdwt1O6DNZLkUGF0JQtJSE8KjQklFdgvOb/j4+7krMVIQ
bRWCt5R/aoXPyU8pwhYwT53CQUEg+brk4JHtnwHo91qyLLYOpjzLKEdTpeJNYPCnR2AgMZ9htS4Z
3mVpKjRXMc1yoriNgIvfJyizGxouJ0+Lvd2bLWwgk3FIkBMPbQOXzE7Btvr9yBmfsMD6N88t9BaU
vBeHazdoPp/XVZfBT5zrQe/NK2glUXpkpzGflNcQiLmIrMyVkM1oFiV7E4DiLcU381FdOwim7OtD
IDkkJkmZNrcOpSa4SvE2pa9S9hRYHgjPj8QSWIxCBISpcvDS97MywuFfzOHBxqw19IY/jN6VM5M3
qiyTaPRhpCMDXkJ6nARspHvJ4BmuY9LfJy85tWYOowkF+bWoYmQWTWF9gn6w95Cp8BGuEbwzQnqN
z7dSNb6HKXqsAXD5w/98Y+HG0LEriBOv4g73SB8b3xb4qeg1a/FQQM9qk5qkXZLdNgMy/+I5KVg6
o5D+rvfV/ORiAMhxcgrFfc4fSKKN5ArZvNWhgFX+UahLpSoLwzp+1dBX/0DlPhwjVlwsaCfbCfpW
Foq0XAFs+KoL7BqOZxWhwpScD6AmdYyhsXrO+vkUJMLc9flpsUJVZ/lxg63J+H3k3iqIREnmd5Ai
irub4eX7xuP2hbWUAh0lJ1kQds6vugU+evNR3Y0vFSBIV/q/D/S5df7zts+laeyukTVqf34wF2Ek
HtVQayR0BU6x1kf3F4URdhvKKGeB2gelLFbmb41rMQdJ75XdF2oe0OSmRts86YDadSuMxYdiddcw
SJJxvtpI78OgAZ9zYMAFR64KX0UWBRYGFxS7vMAXmbb272CpJw+sGSNR/jlalVLl6ydAjfQ0du8N
erIdLY0xehiLMgrquLDoW9zgIqyXiIRzJF9kS2N3Fv0zqqfcFop/v+Ptm1IpaY6o7LNj2Exed9j/
V3/0iWirjTcrYT0ZkKc5BSQ6SSk9yARLEiz5G8EsXBL4xxPj1ynQNA9VLPCMCtHaOtdUiJmR5GNM
lJOUYnZCDnfE9TmEtfbjCSwYeeKubQ2HzHRPiD1KCSrl/lwlDxvtvtlhlJKLJKqi68GXBUm/tL3g
ZeYpU2YQ1hTt5Tbz3KB4qio5nhReVA/qJFkH2mb9KqpJaqZfZPTbocSQaikTqnY/BmC4m67X3+87
ZO9qA9W551lRokhbT8454MrMgsT53qfz6XqoRAqpteD+jVYEjZy1BR+fPZSBi8QLDfjyHGcCmJWn
9YrBY2WfJuJsymx6jmJPfs9FgkHfiuQrBtMvYbGb1gSDw7K/TWPJOC5b91AV+gLWPqaTalL8JQHO
Jfv9COGCQcBW2i0ir4vfvbqc1phwf2ENdl7oVdHdBIedBPkU7RNyyLdvRA0ho2qlv7oOfbBBGrnW
6K/Y3w3ljnHK/1toBhqnUyP3q2AzLZnUoYoYJLUGnQHo+tr6HlNz7Ag0is0uF/3ISvZq7Fcokn5V
XtzGasgRkxw2PKtnTeXaGkjkBVnOlyEx2VsaGVK/jqDgBNDv6WNT3KffiCS3ZyWd/FAoVutvPm73
TdOo0gKyWm8gBxU8VkIBy6W6X3xWQya0jvldZZstWB6LORrjiKwa0hny6JqXFCbDO1IG9sBrZUix
W/1BvnTVPZ5/IJclG+PX0t351HAxOxf42mlfGKhhZ3BF2LfASG2zO5tgpLG1oNUS6lFfaVAfnpvY
O211v9+ZHQeWSSp5BYH5Swi8AftarA7daTGuOamhYqPySISLXqIhWGcjXmws94VOEv+IypUPs3wK
ew+sl5VfqZcisQgPAmsRg0OerEFHy2kpM0nmyJ4TstYesU9d1H/+SX6AlNUwh3O4ShOOc5oXrmTY
ktmsrTxDLA27/kfG0u/Aiw9P/pkX7+QODztzjmJk0LLSoMiA0EjbhMPaqjK08H0C1B/R+o3MuXfX
FcjhTtI+jLZ2mQ7xA1awvO81sXXSagJrr1RdWWS9rnNqakqBSSwxAiAfmiJH08nDB/OROpXueVya
ArrEjxwbh2Uk5rBUk/ctljsd2+vys7TM/+ws4np9HSTJNVXtCQW+X3WjNPL2T3TZVEweB2l/159X
3OW1YA9PqdQxHN8Hh8a72algb2OY2vAGe2bV1DspA+l08nxHoz3OdecSO+XYwQAhrcVvdvCWofS4
Xf/I4U3//P683u/zSeJe932TnDTC7flgIn0uWCVJ7D4AFQOE1RVP3FLZ5c/dQ4dpcAOp+I4dL7BV
hIwNaFvlsNFBn+pFOFHl53/BsHS6BULTnsj1AAhsknpXTx40G4/gcNU14085JE0GwuBimPAJ0Gsr
mMiQwA2m8rEKWYxcrFmf1wOBjNdSde1HJaWPtLiHo4aJ9W8LLYZeKhXb56g7xyg3Z6wqiJDZQbZH
lwIOqW7zDZvyf3Rwjc/znEWiil6V8SFr+aiMB6CUCfkqiAbAcwNDDILIZTtp42V4PwWOu+Khqhii
AD46hDRn/S7sRuBNu0sGwmwif4Anuc92TgYv+Rax9hmVu3ejdIzev1pv+yzox2jXo3cvCR+R70um
twraqsCt94vwzWZFUDPbAIrQJPpNKhtH5rhaz/LsD8vg+l7+n0aZpK0smTHIEsVGR7tNYmsJvCiJ
/x89LoBu62Ew4OjsQ8EBQgI6NJuT150W66lCSudBwig7iKwRaWvKS7ME77tREtJRUUCiQH5Fy15L
fMHRSUJ/lLxO3tzNSiBs0DjgiBG1FGodsZF+heXO+CXgQ+whlajer61LABdUYzqmZRIXe3So1uv5
AMj4PNFeJB/JevhZNP5FWsml2qfnVJISKzadSKXZvYfIokgVRIYAVWi26yPH8UP7rCD8HwnadRUo
EX8IiEZVR5PxC3DoiWB2kvuMllgbMCQxx9aDrEEMR1PBacfzaAnoA1RBYQvpnVfdejYz6VI5JaKT
K1wIc0uVbsuFBkUPT1BtJQsJZSVmKZsS6Djlin8J3sHNgSwQFHi3QiTCohhiNdCP3xYZi2uikMg6
uSppeGoIPAXZ0TNAL4bc9a1aXigEjDSUbF2fA2uLsvxAZviZuZXPQGmRLt5l9ra4Ti8Ko6FlaFFG
xXfiTSC+nFuyNNmdLoA87GjQ/IFi5HQWtcgA0bObfcgE2dzoWhTP1cRwaqGhNHmMgHVHURXgNNEV
3ZPwRH5iJ+1Ad7JD5Vdmk2jduALWYCmBt/zwqFMWKWP4riZNbUwxX1Xmmnx4EOfUrNaA0PrmLft+
PGGS9M6U6v/vJ7S3DX2ALfCvuEyd5px41Um2QRFKyp0JZWH8B1riDMfW1ymzijhlkgePg91OyDna
9dxe7NWeRDWfpyAcDE1irSgd47dKWRuJKmAV51h06ZB5N+6RjSrHjqDhRMiGXnYWaArKSaKqhoJO
FJDVT9AF//RTK9ZbgKOnpmYGDETRZuTLVlMONG7XZWV9nYdrEQvdjUqusdMxsR44w51CWrGsDinj
JHerdUYCk5B+zwO1s4sUUB97LNKkxpUNVumyU1/pnhEXzrsDc9X7SR+Hgq5KZtbXVJTOqhPnlfe6
A4ufhn6ABq/VoOZhFU5VvAbO3vKCtaPwsocpcZt+OTI7l5v5X+HQhaqNWRfBYW3MX4IVesEghf6K
aWWwiYmKaEY6HU8XUbT68Ngn++bde7n7nCE234P+Z9xBYePRmymberU205IAhm6DiD6e8OqZfz/o
E48ToTNYnjuUUUOhvz72JPhdUXEj9+jLylw9IgdIQ/X0ntyy4P/zJcms8GC78Q7/0UmMiVVHKuMm
zrtkutl8PP2L/7F567VccQH92ljAFivsApT++R9S3ROi1J6xG9AWq1/GxdgsHm8xPRouItpFpFOy
Ygy9ZYFUqLFZSkw53HywLlV+mFUaMj1qGpiF99zJ5D8M6K+r+TbLjSI4N1gg3Klw67FekG9d+VIU
uJy/VAINkmScYoLhvlfO8Rad7KYSPN6wK6K40B/0jvgE17SII/tBq/KmZ7G1JDynuzAu9GSxgi0n
OuqEwnQH3F6tnggxFDXXKvvt8KwMUxGUVrgpqZ7cIOyHymlKzkIyCMJxmyW4mrKedZRSZ14MmKDp
RwKRqPKd2s/Hznn/mfi0OJaK9hv3GzdsKU/uSfXncOx0OajZtoArEGu+2zi4LZ/WG4VStHDvo+WG
TlblhB1LTCywBxR7T6c2K2OUBbrr5mJEsv/6gWHBYJron1s8M0KEH9jX55edjXpzOljtY0iKZ1l8
IXvT/9KSuy3v/QwEdzYiINjI0+DQuSzX/aYTrrgmrzTuvt1IDlobSyq80ZnXHRE4XwUEgbNc5AO7
yFB8pYbf1dCJAWlDD9iMyyX1pGvU5Mhi60B12iwLt8PzfZYH8V4MdQqvvzl2FZqjzcm0V5IFHyGS
z0/ZHjE5qlIEBK0zRKL0SIELQW0Gf7w34WkhhQLjvZj9l+tz4Ax5/gVOTSlC9tBrDsRJcI9lVLIS
WfEG7H+qiwmi/KhsfUk0CWa0mCuMv899wOnHj2VzZryeTkjhjhmdWt8Kzfe7c+HTtfhNf/WogL5N
lVRFIH2ZjjEPuenWRtxr6dSc3sigajd1Gr4DjG9hapm5pd2ljGcypdYDUWY/mkAxRsIWyTZrNZOq
pk97N+ixZYQyKJ2tKwNDdTCL0U6CtbwtE1no9o//YzkvyOX2QPLs4AQIURz4Qd3PhjHv9NV14wYE
GXhXUf0QugDXbU6VnQxDomEqzn0fzrn1xb/NedGegeEF229P0x/GFZMeoqPV1dpWGg/6lH05+viA
vzeRYstRxMAR8djsfkErkeEgOVmza538P34PTAUQP3QF5dqFNj3UtcjB0JkvjqJT7Yq534Wd26B/
ngZQPhXZrzBPpijqW9C9qDjWntC+OqAO+uVoWURgznYZiey87GgChegoZn+BRwzOjYcmx/POtCCH
vAws7zZMVBwgRy9+jM8VDrsxFe7fD5Hd/MediqsXcGnoov0o9gVhQQ4CKpTSXvy/8USSXHvG4Buo
0NycWi7ZU6xCiwsSgoOCWbt8y/QdhqGKujSTh56tQhBN6wti3fK6CZB+967agGwB+sn8UezOkVR2
Ga5IYw78fxQ0bBGxa+pwtHu24eN7m/6lyDgF/7X2MjWR7nXvoC8LviBvC6PtVVjqE6USOBmXnCA+
veMEb6a/6X992t6+d5GZd8CSsbtoEe2BeCRAPqQfZNnZ6cExI3FHJ/XVrd9RQoBugAtIEn9OJ6Xz
6L3CNvy6B44DI5G/K6XSvZ4QQEaEMWDQcUby71HmEp4kYwi1qx6tqybdEDQxWgPM6UQeQUP5lRnt
B4c4M8pJPX8nzU8fQOiOE1NWpo7X98JzltM+q2pDGrv8Ry6Kr2bKymYnyca8gFq3/E5orQJU330P
WhB99LkeWpe7tG6AhJs2ijzzqbvDrAjAYm8jG530xi8AUQdEnA0rnXHipaLjFGr+CbDEgZquhUiC
Yy80zqdMkOUzIGmwx29HqtF3OrCSxdMgdzmNSxjCMkfndDyp9AniTf719I96XhBZHuXSMHsAQyX6
buAtFvRn4ZGtVM8KsJgsdkwra3Hq8KzfXl2JlsI+hCwXdThlQ0hrqPUpFL8BNZ8dmOny3f627BTr
FiAYKoGKGuZVMjBpEc6+d4HqP/cGDUicrKdl8QmtQE7DfDtz95mQB5inePfagLX2JQAJ3p072srF
CNfVXkqIWyMpuycbRdP/Va18mosBTHr7X2QCnUFNJSkATRJT2nPcw779X8CGd4EReiWwdL1YvXaC
so4Ylcf1GGlsNFWObkStp1uJcVx8KRn5OYJmlOw8gF0hy2TluHnedbPy9p/LsCINKDtBF3N8qI0B
HspY3UCVneSLBexN5IjAA7tRxP1bLWUxgNPvPGUNY1hgvAES/Hv/N+Pu4euuhMVVYHnV/4ZzcYca
kd9sBGgET4MSXJGzJ53o13ImRlKf5CuH2y4nz7z5SSsYQjpQtAU5F0CJe0ilwVbonDA/iwiuv/Yd
vIw96H+bqm4VhBRkk1eiE3aQ4tRFM1gRdZor1fNaqeGGrLSe0nua1GdfoTr6UT1fdihWXudn7sGZ
SGzlwINs9R5MFGuJxRYVXJhcGw7Spz6TN2dgJGHjGX50c0lXMXCdYL6JeKJz3apL/F3Naa+iiazH
ogXEvVqnSwhryNyAjCFlQBlkIvvEzidMu2lh59qCxPTmUsbwu70y9WIhRZMBUik5+h/fW+wKKDJC
JiXBmIsMnizLjRvfYI8xnJ0esl9pE6TIgBidvActeEhSAdsqf7/rNKWouuBOd4jX/yuP3BgVhhN/
ePcrZMLzvDNYQcwX1P9AabIcXicazzi4c1OX/FyMCRQHOeuSvA1vKyGcgB5ULUtW6MZMMij4tMQg
r8H4HAxUBuVQn7NHq9dI8eHoUQtNcwStXSnzvln9yK+EN1sr6ghy4ihD8qj/rzivcsIpqvouzjal
4EE9L7+ARey6b4d37BX/FaAO1ACxTwDeDNqqlbOG89QRuxDqqQOmbJzyrKv6/i5kSsDb4yQl+yZf
FkVagQfCqy8B9n5tYgVVJpcusFQ9+0173R6k0qPWz/kQKGDGf2vqpB3BzO0IS9orp5StziQ6sL7r
pxMigYtUCfIs7/fibtL21zVOvL4lkbRcTdJnJOB5aDCcjYpjhsBlAq4Yo9Wx2w/m67Nn27+IUKms
tkZQ/IqAGerVeeMa+qfjLNhnQ83SEo1L3jYWz16PK5qn7hQJioHV7Q3VynJV5NqhkIOHyXfnvxzS
Ps4JaWbaXV9hqXraQKf/pWnI+0/085YsFL2oemSTPAcMTfeGAMMXv0E/m3ioR6k4Yo/TZhtxGAGb
Rb0zigW5t7iC/H5KefYiTeURvCYqtPaD0WA6JPnXoh7KCDYLKw8JG77aNGJFNazsErUXWPHY7GOp
eHL1pJWQ9p79r+JX6TIC6U2/TmrDWmJSv4L5Rs5cHcCQk0L81d0NDfLLbMHAR5kpjyGYrZK2uowM
RGE2PrKekRWhaZy+DqEpsTBhorTueyfZYIbVHjGGD/Xq2bvmISMfMn/IGjCZj3xbZPb1LLvH2QK8
JAYTir5Dca0LyfGf93b0qDjLCmiLQEwVGob1g5mUb1Vi3Q/+5CVRtj1CJOx4g3NphtEHmdZtfYRi
NeflrbY+1KwrNfR17oebpVSrpxsP0EQ7HSvfOzuwsyzuwN39yXlqLAIaZ5XPWmoeSLkCLSP+Pfnb
Ipfp5GAZ/euBm0BUiDEcjRlze14seDkP/WBfkL0KAifRLkH4D5/NCykIIF2QYzeEsBAp4B44qXP2
H2EZrcMdquzq1i6V6G5pDlcleoV9Hkkc1NVE9wOw6Ap19zlx56h2qeTYi0UsCJ8Wp/Ar0/f3aigl
jA6DwmIxRZNywdTBk9n+X1v/Us4dtXaxxvW2lt981wNVme8A+XyC8QG/zyXCsq5f2eF0X4WuoIdb
5H7yYAMOWP/1dQpNwlT1pDHwumDnRvQPJjI++uOEod3WgPqqn2Il2O5JrNe4kiLB+tKgjt7PpYql
cuNInp+Hg8p9fJwQrrU7y3siSa2bdQzyWqjz/mkOqziyIvGp8Cj+VXZjqGGM05V6bJozzSHxQYhQ
W43dPM7isnp3suC1WUxQ9nRWOEU0v+v7K/dp7UZjfqR0fhJKj1KlDsxA80joYaCOisR7E9k3OaEc
KGjJKLkHGkfDFaUB0/4cgU43jGQYqylcHuheAzpH+43y182W2ijXg6N3tC40D0pTYwPlsz0hNo7F
ieHE2CVAjB0opDQZR8ww780xKlJ7LW7Ree5PRr3dtsTLPsGpg7kfg6KYWGAzuSeVi8ntpRFM3hQe
+pW2iXPLUAKK5oW7xxxiDcZqu7KRa5vTKyFIrqcGVi/TbCBtup7R5mUrj4qkVG71C/TwoBNZVwbL
mZ+Ebdfjg+8l1pu8bn10xQ9p+Zos6e0qhE/Auz884OxQC6j2efB0C44rDGiMgobuIlveCuYN35YY
0F/Bs4q4K2LqrMnIovTjm9wWyc6mzHyDEozovOwFPBxRzp+IQ16kvia+AP/CJd/e8KbY4+TFt/3s
eQgmcj+gS8zU3lNU1GbIifPBbhgoySC8LeXOoyBl9uFW3RkOPyb4ZoM/6R4CGjHTrRKmVkjxtWki
vUQ3MkMNCrEPLTeFx6AXzrOPm19zYoneLqqJ/+zlGXvBXbF9gbY+DZ3dZW6z1XfUaP40kQr/1CHh
JyM5b/9f+Dbm9ByDKf108ibFJzozVHN2dvhaiDUJtjoVyIEsGtobMcxldYe0Q4ZtTg/WldAxxzQ3
Sr1oFgPqh8oyrdJ+SsReb1p+QtEFtEWdA2zjS14s1p86faGcldUweVrLUskHBK0aB0VHlXr77QBk
dbG8Ty2lBBk55Hq8tOsQziRu0il1WZEgvvmGJ5jMMlSYaFVICet8mnmaaDrVwMER1dNJf52OyIzr
/h7PLsixSfwC8LrSjBuqGqImGL0T81Tg4n4hNELUbiXHyz/0Pnntsv6UXb5y8PW6tWdOm9BlGHH3
7vcBtVJFVBaYFEefqnim6G36+lyc65TOlW1hQOvq9auXl0pvpuOfFmte0RPJ3Iu/6L22O2PgrBKN
Bf4d+gzPMH6L26jtNWpOx39kF2znDZp5ZcVj+y/z2vAN+uSTuwo09poMoL2Gp3rqIDw5LN2GHAxq
QV5vhwjiCatKvvoPWy7SO021W5q0Li6uejj1I2p1YzJ5ZG/fLW+wQc3mCnpX82IyLicCECpA14iv
Xl5dSKn+TSk/8YNXkKX7DfvsbTduClXjMr+SIkQEAwK2rIv0nMdrSWTWVhz38IqFzMrH/7/Cnfc4
jm6cNtsOxCro2iyAMT+Dop2Jd5OT3fjvkKJySQhNJr/1yUL8cbSv9jwmtC/M4Vb3bUJbEuoVLhQ2
UdngyTtcLuDAJTJHtAYL66Pko7ZrJR16Sljjki/Z6AKCY7/k3xg7Z9eoLj+Fl7eGiL7a2v4GXEYl
CNl0pyeHGOmSanNWyVNuASroc1YlAqFu8gHk4c2/mSwzLwmfjBvPNzUIIyotawPLUwkzWwJqWi2Q
nT3FTTxYqr03AomdNMqnTgmq+derVvU/cq9qaVnRINFyplpxwCQVn4KJ+e7Zcgbb1+ats8n0wdvb
6q3TRDO1xIrBUnHcsYyoIzZcCQv+M6xxI17eaqBNFE4elfcOW8VRuGut+YI/LQiWU2NXfuKWVr+P
AMhKL42JLT1NImKmp3c76+A5qluO/uIh5uxjdoBvIZjfPeWDJRU7ZiaLzPU4s5A+4s/kIrF1cEzi
Xp+hK5Zn38U7v8Xp+aTmZGEV74pf1z/4wYrkKA6QmGnqNSMaChwZSI9hqH48QAtneVkeDAcsMGbD
uYi0MKxEb5Eu0t6KyJTewCBf5J+gbJ188v9sGevdLkkytJFeBSt2ncZQGrhjESy5Wwpo1tHlea6c
sm8+G0fEllrEHDZ48ewvxurj/kM3SAqHDmf5upCEFoRTO0t9JTMKSKUYS3+oOIgekxXhoqgS8uW/
wToZBFp9aWxZVosFuLeSAhG0cHwzQTeNKavWrnMmLXoHt2ZJjwhvjhSuQX1f2V3fQe6Fy8wJslgP
AMvEHIT0r64db7fOBrJw6uHmSMtrVB5FDyFuoWsuGrvnnfLVas7Y6zDnMyg28dUKave1Bvbfg/V3
l1Cxo1gQ8RQIoXATsZVNhLjaNcmRPQ+pySpvPLNdM/TXpk7nMnzFtEtB+iUMDEPUwKTyogPkGDlh
oUoXJ6U+NCPDA2cRVZ19Epmwo44owrNJd8cWAoZN3OrZE8AujREZ3LMdFQ/CmhgoGMSmhM6fNdsX
ByjaOTpEpTP658L0nlNNuhBz0LZ4L0eOfqVWJ9OG+6BP5UGL6nRSaKUnzXOAEdfUPiDaS4Igq0jj
yYcrQc26r0UyxY3xXAhohpouVtJzlupyGJl8T5m/lN/0rr3Zy30/HAA+Ir+jTqckLEhdNNY1XQMG
MLxHoTqyX71aQ5GmJrAPRFMFAK1/CNivnvPhsfWFSXjs+ZMe94sv7dEjO9JHZWQeJ5v22JclWlbM
gU/JchaGvgEZzLQQFduCaEzksJORkuA0r/3fVf9zYsHAVYEKlbrj0VI8+n8keb6v8WSC0gaSXXFz
snc26/piudxI4CAKcyvrNOPm3YcoAA42g5N0zkIB6/dUlQ7fxUP6h0VBrC9yaRO6SlzKbGWnmu/g
fAAMK0a11lGjcX8lhbvKlp39HtSE5IhieLx4wJDF3thaFj94Z+wf+X0x0vDwsnX2CzLSidf/Rgl6
4IM8JqZHKUjYgpjRmvAhLZQrSHrDTQXTyR9GlgcAKeJzKbCa+HhPoTTfYPyqcPZjxSFPtAg3xxjc
KPA2WpIjKxpw8HOz0XYEaZRiszBPBFeR+xPqnqfiIfoco1ZgVHim1jRz45D7014smtVwJQbvhy/y
lmvJVKhV+M3NNEdhhafuMZKGzYx41s34o9pIIAtms6u/SqsfPzfP5eXTNc2oA3QkhBQq9EalU9bl
72+DqAu3eCKVU0xBg63RlWeNMEWk1XhOq0LCmKvkHRbPpm5tY8AzA0qIj+cguYAJHjIWMWrsjG5W
k3SZT70BSDtmL/jsbmzBNGAwtNxeceQLdl4vCfsBf05K2W2HF3g+5KW8s5C47L+q/xlvrw+cOhgc
EkXV9RM8/NaNI6JQ87OHh+s9NdoxemeCUtV8i4O3yQG+OgXGzl9RW7ZJ6ucYbd/INyVa70NiLzqG
BOqWRhHpetmm3v7xHc0hV7KuM+8LZzvMUDnPMDHAkC6Tj9BnwwlJX1UDN6DDnetWS74OX4cR5LRD
DKyZtaWNRhMkuaeguODmZ6YlJpEQIxX/dRSHWKyn+94RfT0AcU+xrx2dSI4KQe/IfaUdcGuUBVpW
WOGgA0wxU423fDHPScEKdbK2gE1wpTdOqEdVws2xDD3I7YcHHzq5KLqZEejiy6bsEJxnBXHOqnV1
oU72Bh8ApjFe9l0l+xxyeX8SlisgvmTyK0KsVWzRsF8j51y13UOdjYnYLei/vT9UUzQFgQUD4grj
n0L2tS8TzqwHZdcTQRJFL+RXOg+5QTtXUBpTHZj0oWPWCYDJ0xnzeZ1T6KMRNiKPMHI2nlTwuJbF
grEePzvSQQwzEoppcd75lUhEOxSSrYTkNO+02FtvCSs9dg/EytSmAq5+K73anP8zHLvzY6s+rd/O
kBtNAyqvxGkUc8a0MZOojsyQB3CLto/JHZjkjyBuCnpDUjQEhRUmblu+HxRfSSM2i/CCfmC6q0Gr
QkgBNWIVBKawUtUIrcRiWQRd120LubmBh+8U4kdf+EBc9xcUqWwPjamON4/uob681348EHyNv4TG
0yZeObYUUbegXc9ZZqJx/0NmiwvhpdC1BKSNnOTZCyNOSfRbvuZ9YqFvcZH+M/b086jHGQkS2iTz
0mA20BHnKaE4h7xr61Mf/3Boe5UuJN0J7OC9W204I8TRHw5CJQGxjEFwDIsbJwCS2hv0nM3mjTdb
nfUWeskAP2GtGn1C9d9hqEm6oHP4B07Zx5mJhJ3l1FKXuS7gf9eLDKDrO9e0wStsiLQodO9dag1C
u3JwX+6mSLlrJZOPSUygTm/O8H0gRf9Y6v1uHpsYwkdYELD7CpAyCpj/8wq9A+7Osfzsmgyp9Xz3
LS7N1d6BYBiS/JEBHCcch5s7+NPwZwAfDkaaHRBSgkOe2p1yjxlqRwNiq2oGlE602DLL/0oE0kEX
RacWwhuZp09one3KikKq0kMa/qWvTPpCFZwPU89bbxbFD7Inj62YAuUbMEnMFPn4EcKPHnGRsoeB
yfqft+hJ7CWAYb1R/0Ac5mppSyBlXoWgdrYdkK7Jo0TN24nUdJHTuzzIdQd5F9YAN2SB/DZ0zv2o
e+myw3CqO7l5AifO4npmrWrWb3AAjVX4p3ykg/G3W5zH2wwlgBwv0NWdyzj++JYnYFZqqlkd2Nu4
37vXy2En1S7SQU97v09WPxoHY5IGiMdsy+eZV37toF7+qAi3nJVgU6B6KtqGw3Y8gVjchOhFqE6x
ij1EQAeQ/iky9ycI+k7DpejYdHM3yL61a8G2tnf6cwUhaNwlcFS7CzjW6x/kfCJEK3yKh0c3Ltlp
g44Y/RYDiTdxXSp2A1UPSuNM27SETDLmFKUyhWt1Qe3PvWEl3oehcbl315Fb0LfjvnCxU0Wutslm
yBLZBJds9b986LThW5LdnBZfcKLMm0MfDK5CZIpeqGVkncQ7yepjGvLJsZhqEhwHHq1pXD7WEuIw
mwTW0GZRH4dcgcexsXHXdslOMhnO1EGRjMlaMhlTuSf9FudSzo2glu1grC74hW+ogcSIVso8YvdZ
axsQ7gh5XoofuJGao5dljyAOLwhWYEpABKZ9c1rCPt3EKQy8TNYQTzPQ68BymuE6hbktxjB9mTsi
yFfULjdAHQ6MF1zT/WT6NxvuMC97Oa5O6b9UpRKAjpNEg7l16jZwwehjKUHgmCTqzB/wLZkFwVTD
txieikHpI1myMHjy6MGftgyZNI5zFtztIfQBvwMxZgmYsgQUQlABTXzZ/5tEQ3hVp9HcSO4iyPwN
b9Q/RUCwYAQEEwUvzuF6BbnMqHXw1HPa2pJ2SapxaE1eA6rE1l5qCHItSxZpoP3tR9xS9BlahG9X
KncBHix5P2wnuBWtkK4RlV0LLLu6g0gbzCTkWW7olt+96aLTzbpnj3WB9AxV4jE64GS7hLVtUcLi
lM9BD03dskgyfiJuGySzMY5JK3xqg1lHTuWpkzHk/YKzTenvG19C6PeY0pVwjJk14wWCh9Apc4kR
m8d63a6N1eP0jzKV6gQqGl5ahsdFO+YVPgiVGQjy19x71Z/T1Gwx/2Z1M1MQggWYjQ1HzahS9SIC
LGUe3o3Drsk5jOMsUTunkGJZ2SpblIBTljdwQg+O5LBeou/CzAtcx9emGXpT2r31CfuEw3jA37YS
4zzoVFr/UOAyuW37FTeyZ9ZWtpTBJI8OV1+pOnca5JiehyQutgx+ybjxOhjNXXKyU9twbGtzfjPU
B84den5RNd8eLv4JLjTffKjK1PqVpZ5dV6QnNsUlm4mgb436R8EeNU5b2x8PQSl9pIgUIe19kwgd
2OYTJ2AttbBjnXDjZ3qMgLe2xvczdj784OcnU40WsokRc1sulRSyFyiz2Afx/FlNv+dBCSzRdzTm
KcnHZUOGa3ywzL2lFnTZ4h5u2T1p/BVSyobqRNopXjamVDQZ9hPXRWkhAdhcp8TSj8lY3FDwqluY
6hhcpqC8bpKf2BUqn5rj1IMQgr8P5vfbzNX675DCKd+50DJFyjPF0ZZK2AUL9ZflP/3+0/LgxSJD
nVrFs5+XeuMJ/6i4MYZaHD03etCosIDJlTXr3mmwhZc9he+mCXsJh/4PBUbVxjBALtJVrNSGIggp
2//5aFlnFgIsW7CtAt2fwH96/TbWpD+LXvDhNXJDuqpENTBVvcWtgg3TzDqJ71pPIj24dRaNR2vD
q6+f2wa69xlz8scJKyBGW1C4KmN1SrQpTSvqtZrLpAUjiNvWabdPQG4WoEoyptve4SZjsDO+6YUD
XABBAJ421NPXnUy5aSn91WinSp2thKGAI3nTNCU11dXXyTh7W+I72ku/FchE9cS95ihJ26vCO6no
bs/xIQMJnfe0lBcwQizGFWfH+tzAETfUrQjtvpTqLSu/SmG/zKTv/lqyMyThC4S29PZgi1EImVrM
m6OJqNwQj+cuxGM2rFvlCB5lmY0f0Rb8LR7LAAXMCfILFXS42M3SPwmO6xirTQpQaiUOjRqPv8Lu
I0mpMMEcYfaJbvz7mdS7iHDJ9T19jC76NfOB1tRvzidv6nZVeqlk2i7ajgOaT94EJfKuMZPN1DPX
JBjldY1X8ZSI+dIuAHkxzFqS9D+wRcUdYKHL4PRkTT/2Rgv4Egd/UGxPu1/z3hdawewAWUf9NCXb
pXua9aNgBhLQe0+Kw2/3RFOuwBbZjPwlO15Si8mDorHc6QXIbNO58R6EmgKVvcJAuQNUSJtyPYJa
eNA3mI9/LFBhS1yMGNf5me+NBQm9hEbeXSssMhVG5B4VN6dOVZ5ZZDKtyEzzyHXegkdhZsrX/T7c
6b0vVycvQSi9j86qIxQsIrKU3S4hNZGew2XbuNxxqnwkw2H8oNUNHoCN7Rhxd34IudzwAQO8lFUi
3uSisPXx/TfEcmhswwintL5NQBNrXOvkyw6zHe8FXJaNG3y5wkSszbaZNkAyA3ORMXGx0qwmNu/7
h//puPmJ/nAzjI0a2TBlVcin05rKMqHW8rLCfA2iOUWf3KcL4yZ3ncv9xEnSvlJsKus9YCtSZhpO
sv+2NL35Rgve9SFfqrD+/AcP13k73+NljLhwvVeIRKfrfbzyI+CqWmn05zGzVxCNEbOKH0ITO+B7
vo6wI7ZK82admgeFwpPOEyUOOgTJFV8XFi47+0igkjpdXEAfwKbpqVYshAdrrVM4hHBo/3scnHIC
ml2bm9wkX8hUTmmeZ2HV+8AD0i8w+Pgo/zrmp9OUOC/g0QKaCsAyqA6YKymSd/8S38aYINytj1C0
jyuXvqtOyH+2xFGpsTPRqAJa2dKsWV1+h6qflzcIddbNcBMe6r/vW1L/HhWG5Fhxa3z9TcQpNUA3
zo5xzQte9tMGX4yLUSXRN+MRKmWfdDthsvzeObqI0tAAchJkt3TOmgGGjstpLEFksOfAVfbW6hwq
2pwZvrZ7qyHCi9unA3jmcDOJKFb87lCaHYRvVcVCLglk4jmD9ZW8d6XZa1zPRadMck6WuJ0k+fal
uSj2ynWgt03QsQY+1cV8Y5+KVyIL/cai8tODkrsa6jbLrM8I1/c2vMdEmnqrFrrgMcj6LQPseJmU
tUzyzapnBVIEC3+f03SwiOKqt11631aQHh87DSc8qTNmXRmENSD6lsRq4hXYo2y3QlDxsDUp7fj2
Y5X4TuLZzb89Mpg1Y8JhGuwhZ+BnQ23gtWs3SuGharBcLBPaHIMtfu2Bg0CAbh1tc4m2JS8r8t5U
64wlsstzZuTzccMpeFoH0ClceqQZQe0dTm45b/SSmNZn7NCBIBVi0UhHQyN1sOTOdH668KwLDlDz
X3p6qBfxzTXx6aU4rh5VJO32Rv9o2xPWbcb/9iWAwNyDKZ7bNfs4lMYxmcEk/tTxHYvRoQ2zFdM6
LrEOgL4YJXRw153wFbHnlhJln1LCjY6JBU/FOnj7Duxuclo+C9/ojMnjAterRR606KQ/DIIl2a/6
zxEa5jfnlR+aLw5a6hefZerMI0wmALkiHEnkYn7lIa919dn6KnzoHNRDOUe61BB35vPvSEeNDvMx
6UhV0OR3hIUe5pboJjNYRZqvTqyjA8eAHWE0xIkPPDJn+ws5Skq/X1Wo2+hfHPCJXVdV9OFkWJ4a
XEuFbxQUCx3RWPBm5QUqBADmsOokxSzpY9YUuk1Z4+DUdI2S+cBL6VqBEEIYpduxK/1OpPy85Mt4
fk0WtbpFzYVvAmPd3SplrbEW5VI+ImxrA5xlG3iqcRGIrunBcowUkC1K1JiFKhT9T4a4xg1ZI7U0
044rkOPDnRWUlDVVcB6U2/2eXXb8+4wNEPZjUV+N1nq4fc5JWB4FNwEZxwSDXiLdAR1VlWl/C13k
4EmACMcnobSMZDCDu0xxDI7wRYV6s4blBF2ILo+bVEXGXx7De0psNjXhmhra91lbPDKgmr3wtiGF
TV4oEaHsaBS4u/2aSRcz/2qzKZbDT1m4UzzurjcBN07ObADwWKL+voJ6nRHsvwUu3qjbes+SRSC8
IJmuICRMBI0IPuT+55W7KVXq1wuew16x9M7fLgHO/9eX5bo5isX7KElzcEPOWsTpp8Wi0fyr/osF
fGus9IZpcKUGIlPZ5suK3hWHmi9ezcVG4m89Hnhj7WTaBhmasJZst9Sob0V8ddFKTsxJbBgeI+Qh
rS9fJ/30ZTou/hN5hZFyTDkvm8bPGSBt5yFk7h7LQsZUriuzE/pGTmkNYVYrhfkN2wiO02rDv9Dl
zx5L+E0FQvm9ivyH9XSQdOO+6ph1ZVwhpF3uvAy4cN2mcrAJxQiS2p6EkgYrImkQ43yC+SVL4iqV
GKzT6IOlmQiGV1ZgPijoVu2zuwRNY8NiJE5Mc8bEFoOUWoIQx+TYmafCnpa0TqQ7yHTAIErbpEua
yBqwo5VIVOsUl9q8hrKztqBCZvREg7CEyJnWwqTIeBnhlNX2Hk4iUPlN7J4342V1TL0nASiSPne/
gQW+W67p975RKKN5IXoozJcs020zwKzNC/hM9cZNe6VEfE+iW8BMQrngv2hpeA4FnB57peHy18Og
/DuHVw/oSFWpEoJfzjRjCzGGszYNpAFJUFqfOBM3KUP+OEPvaWtlOqEv9Ca3PqjVKjPzwDr4bwyt
I+E22MHH5xzoyVeJmt6r0fpqvR+B7w4Xd6320rPcm07lpTOePXf63YzVmLKXBE7ptRJ5/lwWWUeg
3HiJbeva1r7qB3RhC4wc3zyf5sdtycmq63Br09hyySkoc7cJGNLXQsMgJpFrcu80cAi4X8Br3qdY
vTrLt06SXayAGc/p4UDAHYQkQrBLQ0qmzu4rTEi2wGj3qJvsDIPw05cTmb9bVbBuKnnvIPHr8weD
jOYrm5PWQTIVKlHxiOj6/sr2eLo+8ID4twG7A7zPg2g5DTlwwrcZXow0Dpupv/yZqNrySW1XIjD0
93BVum4DystZ7A3aaroPeHf2fKqjkh8A7kt7vpnS2T0pWQS6KsHda9XhFEgvNB+dJ8TjivZRJ2hx
wyMKCgRCufDcRZ+mCFIaBCIUOUPzwFfMzMhAgjyeozDyUBl6s97i+5OHe+j2GmK5mJCJrwxhh/Eq
YP8OIWeDY/ct8n4t/yK6rGIRG94Q7J9OaUKchUsYLeF7u0ga1qygzahQIJ9t0a34B9fYP0MRvK1E
zZvPgNSlZonJ3F20bB2343HSxxcYbO4CHzcicU7wqppg/zi1dSFttz3nZIblYYtyJZOMpyqya655
SnP3I0ZKBX7HfHeunKRpyytgV7WD7aozkeQae9o6vDTouXAQR7EiKCQrm5yIskiv8SknMSODYwge
QksTHeJdw925NotGcXDMDck1XiE/bNvu6+5C+1lNEpiZC4XgTsUfzbhhXu4QUps4tGmJCyd6vVtG
9X4jPDw3PGoxYtStl4sNB1y9GSbkPvA160lJNT9K2G/WLu0pdjX8i/zY/0SsXkxWtZ2Ytvew9cTE
/jO697xhXU8cPETDxkCA67zU5OGuyYjYyKpSnLtvCzgf6f8wAYe8rjIY9XR+1LLrfhyTHtNkO1OX
JZ84w8KuuEC52bfr8IVC7ufVSTn2y+K9pkQT0lZP1oLgqoNHT1ki+W40/4MlPVUqeXlbhXsy8+CT
hVvkri/iypLZQoF3Zay5e/uy+dcnBqfq58haWu/FKyv7RQLbKCXfAD5Ba5UlZlspdZfjBpFsZv+l
ZAqlZBEvcKGEOe50NFeH0kyTQxy/kznSPHE2kWsKUMF7cqtlqNO3nQTV3adTCTEasd6kztrDIVkx
MyZYI+SNX6AdFQvLXbUGH+BqnP6JBysBZKj1hKY9QN4tqdQJPpIFUCDo8D/7GD6HHY0j1szgOGMd
WkIj8XBfEemPoqHS/6YE8EHn8h0nSCHr4VzDT7BGUd7NGANfGPd1PTQ4U+ZBilbd8wD/nZAfFuU7
mCtyUi8jM5rfZccXGNqOTIrRyLiaCwXdwR3qPASjgirPY3C6RLGJDoCF9nJRaSfk6DCbPMZpTgeg
V4AjlyXQXpKLASmrXmJbR5NQvbQAu+gl5F/NGnE+3Zt4PwakNp+8Y25nzoHGHEVNvM2xI6FaKr2q
IYdfn+s/S25yY/dlGc9oy/NyQT6z9RcCAh5dwLRL+zhZLJIt56Nn6nEch5ThB/m9vzyLTO6VQdPW
zOC5s6LoZ7yYjWLAD2AhJmvgPmWZx7vNHUo9frQTv5ouC6WIPYe8nveOzLuA51jsWprAH/us2vLA
Qqdv8mZHzTx/7fbogb51+eMWJv2XBdqynAtwHctstri2a2cFKQvRPwKp5j8tUW3B29IqFQHnsmKo
8x+tfU1w/q/TCebyukk1b7K9TwILB36V/vkdGCYhDrkio5jWSwNXGfbpLcwG7Y1ol3v8YaXU9VP/
U+Q6RMWBjPjkEPoGGYGn6HqoSK42DtklL0CMcKP20vceSMIwK4ps1NyzDYxmtA2jNTGEaS6g3ck+
V87yUqqcU7mIMcWiZAW7599QT+19icmFkmdtWEY4q6q/geAhSvAjQrsiNhwXN1TePeNiEgG4gnH8
Kfwcq3R44sGc37tXXuzZV9frhnJJ/0fYAw7408ncZXm5FER6jHHFTzwM4/F8mjhS9iBkZJ51eRbm
Kkdqpz2h0tqLJoAP+nY3RQy0e8SbE4El7LC5SvLjJo7Q11/Lz9ctgf4D5mLZnORd4kc8OXWwe6Mn
YVwSiHEHccF8eROSALYDu7g/lpCoBH55B08WBigcaSB9JY+45XtcHftZBJlGscmNBz3oSm11qW1k
SIE25LxCalL966wVRYqt6oPh9/2nERTuFoCF3JqF8HIost9omiNV3i0Y//1KK/vbeLazM0dmUOvH
/106LIw0rVD4Up2jxPjoTJThlGKbVqNmGST2tl75PEKfEmMGVnQIPtPxjOHKo2wF+aebCfD7W0tO
A2FCRAOcXM8GQcjCH1o3IWvRpivP4fuD/5NtQFrDXQqCsVAJGx5ab20F2C43d3d3SuHtSDZQ1woz
Upy/BNr2y0loTFYZysQzUM0a9oEnNmrSsQLu14SXrNontjFRkh87ii5pYMNJmZx69Rw2B2RAS4/6
/Fd+p94sMC0QglFruHpi8hBvmxO2yznQmt3uZqWVFRUuEIutiyeRUtMs5DwiPjU/KMU9yL0TGu8T
l/0VC3NKrx+Dw8TEtWIGMcT2PAarPxRPRfaBYFFOFNMRTaeiKqmRViBBPiVh0H0HLFF10cqYwmOC
Gtl+Yf8y73hAxeXiDtNVr+e3DD4q0vcLR85TTSARAEAp2G20d8DIIKfiUUyJdJYfNW1TiQQYxszz
WWtJu4MrP3X7AgXkD74W81UacYsy9ltPR82PDqDQXP4D29Kt9tkeh1e1KdVj3hajN4oZZRNzXn6y
38aVmtM1946K1RiiybRNw2Asub+L/yClu2v3O9KYNAKBE6BTBwXwB6OPZDeLfbJS9Cz+qppc6pNW
CYzVXrz7Zu1pjO/sO/eis4g5xnRxG2WSnLu8E0H/CrhaMow/JMY+36Yy19KLwH27Pd/89edUx4F+
GjZrUub6sSanU4TDXKq8Ryki8mDNeZQYHk1YrSIVhAjk4rSdaUvtHFTg9oXACdo1y9lvp2zhV9D8
xfRfC3H/9qQ/g2iupAKDH1AO9J6rteW0LviOzytD22qZdK5FHRAebjES6DqUes0n1e/ml69QYvEr
fpO/GiJtGUyTzlhH5uZtJwp9GLjx8A6nMqoZqlfePdny/oBjtvZfNaegyePAzCOCTV0Gt/HpgAsD
bPkgCplzP0o74XqSo8oeQUJ/Hsd+MgL7PEAOpG69/NdFNLLhttpYbJtijmMBX+PhhWb6Gpu90MDR
58bghp1e657kUEBCAi0ivlUp2Eh/jjJmX3tDdSpRkIAQA8aL3pYC33d7zPhquS07AnpnyRuUyEk8
+rEJJpSzwMKsi7Z+H5kDr8ednf/pHinUwRk8xYRHX1S/FarsX93sar3a9DUbzzf4IgsfFum6ZOzR
5fUPMdQEE4ReWGsGQgRtgVMFghLyqaTG6FHszp9Vao+yQJO4GRqJZNSMbM2JqoC4DlzMJyXPtYwA
kDHjxAaX6aEGqIuppzJb+UrR1NHtoea0esF+gmmFemY7mBZ1BaVQDXGUFZ1hCHc/rm2e3uys9W+D
uyODVJ/c5uw7e52H+V5VeivKvc2UYgIz26dyGWJYsfSALAAeFTy6GhfR3BFEU130KZ+PI/oV6/be
ZvuqHrOlrpYrWKOsVmdreYsXuKb7Q0KJVQYQo1hpsyZNYu3/bKvUtbsFmlu8ATEruGgvCVEUS4ub
5eJp2wBrn9XqiNQBb6nkowRvEhVxzdxuEH1mJsL0I/RwIQLPmVNUEC2FKBZxZqyAihREJB6g8Jf/
fHy/DhNlCoJGYHFF2FseSJbYHSBCXKfUg3Q7fB2mV8sDC6FRb0ynD3bek52pVkQgxX7st0VzqzGt
WNhHNFt0D9VKfthbiQckG7XXqVxPYL1NmmOzwQD+Bog5g6AWsTgAZ9HvVuxt9qNR9yFrG8jHPdGj
kiPFXfs1Eqc3m88esT6RzSghZxRvNc922UMFEksKtxTJcS/CWvJJ4Oe685vfGfTXy6dMmVmHpeTM
+ujAi24GEOBhHHQf2knPi6wWDoGRL+doilcmAB2S7eU9KC7eKMEz8naQ0nkYtsqy+/wVT4dyQv3q
qJ8WVPsin7XIl5Wi6KuvDhadiY4hJuIl9/rWFyfRRJY/rgv/9sS7Ct3YDUG4EV99ZD9Lsu+smGhv
9aSeTea+iEHfAzJ+uaE/jF3a2BW95R5gaiHOObPlE5cYjMQeMd1nnyWVOj6OuchCzSVBit7nViGi
5onhKesLi4qCN9vcNG57g+uflcaABT7JmSTBmjEx/sX4mlWtUhyytVKMzpLfqEi0H7lqhGjF6yHL
FcKQDE9tFHgxxo4bsTHAeepjBs4WmjrJgnIRHBs16mGJNkohRis4Clf2FPQWPPImnr5sX+3pqsC0
f7fajB7WcU8pYd7Mjs48edrxjSZiueTgyRwVfNc+7vgq6ESJbKDiIea5n3EcFt7J/k0v3QiyThdq
PT7PE0rUxrjZeBGvMXwwOUIcqYIDaPWs0GZ0YLIuLSeLoQNtS3JxXpUgfoCYE07QNjy1kDgn0RoP
QT/4NmljLvHlgEDdayHsq5XG2J5OMG7uJfrACAVabSksA4u+xDLVoJk0T5cghfhWTGDkAdtdvd6b
CSTYr2nbQN9540vsE3rmNr7/bEDlVjOzn2bfeDStBlQ/7t6MUCcT/5Sr7A/6FFtMAU4pzcuROAHd
ik3/oBRrRwgGHCp5R498gPySjd65qJGUnbEQYLeUO6rY633rXcv9lygqlW7/D2jS68NCVqvSoSpi
Rw1EckDbp1cIB2+BhyBBMLY4f/UIFIyBAA9xd7OfM2Z7ic3g31ON0qY5lM9mSv/dBAc/Bgc+aK+s
+MYB/4EeLiKVRZiNzHA2ON5kovDqb20ti2Nb3Py8UOYXb782spzkabVQQPyFJ7iMNFBNUnjSfVxc
rsZL9xbIwXwSe2SF+3LkdvDiCxZosQUucqulofDeqjiRmD2PKLrbQm5mup0VU6XIOMUobkIj05lW
ULTIgci5OQmvmpz0qbHM164Tox/5mqtnbkTxTy2v2583sCCuBT+8ZucB/TwtH0VsSZSNpuGEIdZv
7ajLlXeF/wMCprBXslGGA/oVF+HT3gTKVlt6/+E0wjodUPA03okZna9YPTOV+mVaMN+jRR5aHNru
pLWHEzQ2SZFy9PkQ3qoI0BZMTOr0L7SvvKPW9tOB65DZR6ofsPlN5DbHtscmWNM+XAWUcAVZJMGt
PIuLxWG4RzoN6MYJiWqW0mS+zn2g2Gr+qwwKkvqnWib7Ip4qS1oVNJpx4HeD0yZC2/Fd7ncisrFH
UfaYAiiWgG2qC9BO169v2ierc1kgKCBUENvUd6wNdslzaR9dU7vaJzROAl1Cz0LNN2siTaO6/Sp1
Msrw+JnPh/PzvF5jmPzOp8qR8njviR5aOPWC+4tY0LfW9QnrxSQVMMIjGlOC5qASjG5mHh1ZU/5R
/I+sFlG4ibbipGKbuzo9Qm4LHSfN0URaWR5RdaZoRnbM5w5dW17JKcWsCvTMGi8wxNVCGy6lFtK6
iqQARQJpHZtk3C6DXf0/gTwDWJiub03vfy8kjuZfelu794mH6F0tovZasN8QOqTCSwfFrsRpC646
RdTGdFbBREPJl8QpJVJq89ziY6NL4JouqFtsN7FCaWajUmD7gAoVrBCpvz6E4pNdcjdJsRmgP0UN
CTtJF8uRCEwNGVFmF6v6CFHZukLS83YzW+C2HH2pXHxwZqbbkwj7FOD1amnrsBTUi0wH/GuqwZle
7rnzxve1b1xLEcu+SJDqv2uGD1qG3v7hNvqn7VYjXtTfY4iv3WxK0jQP2PGoTR+a5vHFOFk0QsjD
epurEpVhfriWud+IIp3QjwOZww71Z2l2vMOuw51bs8xV+f240Yya3YSvU/PtPr2kvq9qheQFkse5
TePom70ax1oMsPSnFJojdIoC/Qiz/5FbFO3r6upmZG7LgcvPGbcJVzCnvyhW/aIE1q6Rd6wN7wo8
Rjfulann9cVLtVeC6Ugdy+IyG+khP8OLLqGDiGXzGIoMj8oGmIC7bVh760k/Wmf+ldN7Jf+ydm2y
Mns41Y0/hVVmTrQ0rVIs09pFxHmfGh7aSS81yhvduMFfoHF3Zah/RtP68FLhCH5GwRC3XqHLvpNl
8fc6oQFlfWh3Avm/9+IHf7opbUZCMMxUdPDg5QsVwRWOMMA2laATUs1FTzYSy4Kda8Ua2Ei1/U8q
5Nld+whLVeG9dOX6HuU0fti3iswsn7l+Nwsw4XrojTDc0TXOe9JX1ERDgI+peImE8sIBz6KwWtOr
hTDP1rLClgfOFAoZFI+iEpGIF2dehOC2f9QDQ6h0xM+4Bn2u2vElDnZ+nB31PIS0BnbPZyQVvrB7
N6d0rxPhnAycHImbbFdk6b1JatvdD8BXRMqwPToPP69CeOU5bezZfVrwOBoyOTBxrIJLhCmDx69P
OwdIuTlOPVLtzwqVigTi00ATOa7USJete37CwGCWWjeWh6w904ysZS9DPxIXt7krtBRRLBj+joJX
b8DEQ073G66Otn9xUWmI85DMcsnCFDXfBNmJdJGnSXqYgaDDblnW7WI1idjnBZNrX16pK/ascAv6
Rw4mS2qxLMM8R1q/Plhxw5dFyFfyjUS33FqqPJlx++JX4wOCNkIRQcpFLiE8r+D+WpsIaS5ztvJa
BYgb0F/PGxnt2pv64XGLvM4T/fUboRB07/DOZogJOUL7xOifL1H6Baop8fDUdgx+SpJpEo9CXPqT
WcbAnJemqPjD0D1CxH4jkQKxTAeGX3uHDYXhsUxdIX6ZbIXfczfd7uko0/AQCFYz0dlhqRw/KZBf
h4FE0m3OjdONuAsmD4qvJ87FXcZixYKKgE+h0KwKNRDzkFisgPTKtnBn3ChLMFxhzwTdR8f79f6W
HChmwJamAqnFoa/EU4ZIaZHqkEmn7s3buFbs1aw3LqTFTzgFKeeKfkOPN/dsBJbvD8+dHsBp2PwY
CYpAY7UfghWTARyPFF4D7uhxVSEHmyB0/qr+FvOZ9HPIo6hwNExzL3/m2JPWtXGxnEeG8xnYsBqC
ZePTX8EnpIU8yYJF5xnv2c1DQViv6V2kF3QkvEGN1pEC2rzp1kzFDV0wio8LOJSAL523YBrh87dT
zAXognn2AsXLdTmWVa3q03dSygiuoWjFvrGq8+YdvDR6h8WvA1FeH4OKaNxXOJGUWCEh9HABnH/v
ilsBqOxOa+WBJvXDI3Kz82+ZiJMKvm4TmkNmvDADuz2Q3tFOp7penaWdoVu8umWCn2XkQaR+KuOY
wQgk+JyXfBjxFWu5LxEMEEBUiPtONMbHvPikhUHzxEqJWTeBUR0WuBoDns5j/b2OAG7xeJjZhLbk
qhI7Lhxma6Bz7a8zi1EHUuGBODSq6vK9J3oFMF1xQexUEk3aY+AzbjnPh+OBiQxG9daRK0mdvnaM
X3kCIF1NRKnIQg/5kDzgO/zL6iZ/3uaG6LiPtPa7EpEkQ5TkeL+d1nAwlbgEnZNQVnFn06DVy1P0
hfWGMBQ5vwUSQjOFi/EFVBlSsiwEJqKLLlMuDGxgzH/aFI/5Hdpgmg9vtLSbHF4sVcXRTb6Dsi8C
eVC1cyoqzxzSuIV5sDDkNTkNyE1fVehKIpoxh8I29ycp4amxfjNwhiAp0mhkd44HeX9AUmOBVOIs
m60kyz4y5b7OMc6Sna3bANUEzGTdiyJP8Ql97k3YTL2F3ZrMbz9gL4yi2KYLvD6pPwwpxy697TiG
+dFP1uoIuirrBhelwVn07zpKQmWaqMFpNYu76P4SzMLt4TBIIo3hDIQ8AGblF9G5Rgc9n+Kagp2Z
ogeAHFkqgZAXPXcXzwIkpvb2sumzcc0wyDVTACYYJD6p0tiPwV6HDIa9/q02RkYL++cwfyEz5U/7
v7jqMTDHU7TGmdOEbiyRqsfuRqxi4RIEidoViU39NIUSi5jmpAO7iZeFmqNTG+0mO8PtVBksB1yV
2EJxocnW10YtuFpP3w+x+V8ORGN+X7OnI4lpkc4CJKLYMhvy/+Ubro6bdhr2E6ZjmPKMYXnbkwqi
6E1DI8BGsP7kkLyVOjVcRr+wKlswJQifhT+UmaYMruRDH92iDj8UxZPusaApuDKD3HxIB8VTk1Ef
QKtTsxMOIXRm9HoXSzJTpOyul0KEE9AwyE8bNvxLLBW9ltOc7utVBTag6tku5STqj3YL5rFxehC1
GPecjYKxOxz51XCW9B019OLtsYFrvjGCkSHQien9rTS1UF6QkZ4Gd1bqIvAkDtsvrzcPcPiRyKma
YD+r/pgt9xqbSFcdH/Uk/FKxCi8rGx2nlONGfkX7J7n3HjJytJpC4ULO5a71REF/ztIiuRbUvsh5
5hsP+GwZcTsh9jpXRBvkgSKGRcFyVJb+zQCeyKONnbJxCF3Ej+/lqIIVXVoBa+oG9Ljtr6vu5jVX
SDt8zBv+9ERfCBHAjiM5NP8Q0NjX2wnC4bKiAcRc70wtw8SuopBJhA3co9/uLIitxFw9RxFa13D9
tvQQwDXnXeydB/u1xr4Zg2tGEyBTrLiA8vSGQNosdqBKXc2yObFEK7GvVISgMfAwYho5jriwBcRK
wDjfNE2Q6WA7z7V/aU5JowQRG8aivMfd0DojB/pUzZ4UtzNSE6+sY1oBzjiJ2bsChsqqI4XE/W0Z
mLR3SjOb0HOGsZDE+xAnsjj5Qlv0fjEKtF1E3ekm0q910gBhlTTrdysjrfbKVTDzgtp2tJuHUeSM
+G3LZAAdWV8wVwphKxDCN2NHtjMapf3m2fmDgOuLJ33+e3NoXyFYMKy5vJbmW8Wgf2+g9ruWwn7k
Q3PBllt8v2AgJz41S05+N/ibLaKEJKnkXUbPIUFvmtXBQ6YCgjJEGMbB/G0LKfqOIPPpxhzbo7of
8dyAfgJuTccI0Aex/fTBkewrEuNJ1LxHRZP3SrB/2AQkuiPb0FNHQPca7vmcuUtkpZ2WUwxFLw3g
w/a/ylzgdRKSoda5jyaeWusabvpIq3JQ+nhhY376J/Y/9jwAo76hIJd9QabKpcPNyK9pETcPjpzV
DoSad49yV/pq5X7JW0w1VWu4lBCuOE5ENsQEhA746jci/ztPNgQ7yFGcLXcyAsTosMBXSbrYi+kt
8EZaxIq2JIPoT6N5uyajuZyzzRglR/oaAjwTcYXiaEebqOUegLQoXqyix8XgaPLvQOcCubNeOYy7
4TcixMY+PhGf+XCk1int7mvxL82YVrzMZre0BKeaibAKJ8I51mse2EsNOG6Nw5AwBu9lMvIGIuO6
1Sbc2pGbvcT1L3PnAIiKuofuXOGqVgFruDd/qTP7oiPPKFfJs+uUoVnH1h4NmMt/L0fgB9AnAmM5
3tTyt2PWj5MWD3m4gbBafYU3sC/azOMcFs4ggLThVdCUu5nwoCemfC2fUGd0ZAfEEfSKPSNGuZrQ
n8EUGKVlgmXDFneai32FdB0a6DT+fT/1pmPEOqrrFQlhaW8ERRdGs49v+aIcN/BgzqS1upegcj2S
+0KmetCTY+S+/zzPihfEEZLVfGzWPD71Wd1UxcganEQk9NvwBnjcqiRJM83NYoietZCTeAGqidwu
+BloKJ3fno8Nrs8tg+jWqeR9OQO635KZX4zVXXPYYqumAxkpJl4wMlTKoJW3NQ7fyvZJhcCI5z30
0Np5nMms9y7TYgc/i257o8XKqiLGJrcoqDFNyRAmpacA3kSXzMQljJrEXnZHtLcOb+Prpl0wwMyd
GVVeC/vRHsCSvkccZyTaCyH3XbT02vrjgNPRczOHQbDxOkgcULNRzRvIpHqHan3+J97gSZAGP6aB
HEw/CuDCqTxwyXfL5k0uLbdGrdNaI8WsL74t+5xPJyEdiHIq0idVI677ysjRjva/vM1GUa45KafG
J+d0Z6WdpGgJndeE9UXMi11DGpUntP/2vvNMUCPICSTX2o4+wbhW68+wqdg2rjbJzSFf7XObfh62
eBZN4wII2oOocJ+cqeQdZeWg83MH9RUqQK2gRzZEp4HdN7xH1o9hML+cFQOgzlErs6l1u3btRKaW
dI/qntWr+yc63xmTQf14tyiFbqJWJDVx91KS0WApIXsPSrr+kJ+cjRxgdcFJLWPmTv0+1FemxGmK
cH3sMdZQWJvssdybN8hrZs0YhQ807XO88RbdNkPKAA3Xw4lJvD479tqMYrobFbKSUWVcD3IMcnnm
phxLPbOX7v/gPrAL2yh6B15TyXm/S+fU2WnSegsSaAKgjzsQcHbGanfcGtx67TkF9GRgEbOj2c4n
ivNOI31H6SuUyI1cZmpeXABWMPOZARNqyfyzet6xpzTaHQwhPCSLAT/lY4ETJ9CQ0vupepmuJCnQ
6ayutLol4elcgX9kVAWlm+WZ3MHYytkntIKDjzO5xARuXkehKf3SVXI+NlC5+4qLnyO1ewdrbbpG
pne4rhLOUyWmNp0e5l+rr/kRhdiXMBj9uQpd/3EUhK0CLJBOj1fODj086NL9HL3fPP36oMNMjLFI
Sohc7SeJrYrc0kV0m+V4Xmnc0AUjHbrQdBLZYFhiZb+OB6I+KFXXTLzmgAY8F3RSF44ZK7kJiSVF
84RwT1PbU0W7bgxBefFkjabpfS4+QaAJiLZSGUCuwK8txpuD7g4QUUa+RigD2g8toPFqsMiQTk3U
OQzRLgvqTW1/LF7kfNWWa48fejlBDwH2IZD8tIYGoc4Bdvng/+kIT6u1u6R7KrM0HfwXB+UmUjjN
7VZDDmwi/ZeQjnnkqx9Iq62ywkwwh4BPLtnSWMsuorZmBMhD8HS6Peb1It3kqRsssIpywnsBo+Ph
e96BRCZlQpLDv3pDr4sLbDa5cvEJHyIIUsqkYFxAukTKzLRICA3CvYMkUOGG2vCfxNJKuBcZ1A54
ktaKYqmruZbLug9u7P0HVgOOiqZH0poxw072w6P57Mau0yEtcoJRvvmD+QdvvjlWLb+Djfeju0yg
32GfkPfaWbD79iFWJ4w00SQJUGyg40ZAo80FP/Z5JmUEqztdBAJccABjOiKbpkjVjugwjq/sxe6R
xTOrEGa/f6VacEBPWSE3O8W/zps6C5W+3ScBl4Q1NpmFBXODBvNMpGzcMZ7/yoMvbg9FBrJpJm8P
4SyJu7ao3EtKtZGcAszHrOdMKdPzKjz3rcXz7eO3Lgd/Jm0Nxz64TcnaAMO2wIKq5IcKnvDgJSeJ
kqlJguzf+23h+ClMdTaiUr0s/NgGmhVLJK07o9OcC1EEiBn5wGMohtjrro1Q9ZY0BtsPE946mF5A
3IocdsDXvjlXkwUZkTQp07MLXLdx7wju53iaFUYhMHgwpuN2EbFdqbJl67UL2HxrezJaH43b0xpa
rKz4rPqr5Hdq4yVB2Bu22KMIRmhPMeH8o5qoWSR4c91Gi5F54FpSKP7WuckQ138ZudBVY84p2/vv
loQSKwanHkgk9LVgdiwdYIfmwI0LrY8NcHOWj1IU5TBxvIGbCdptVCC8iPsBGgeaSAi670+3Fgib
TZwhfApPGxuUhB0GRM4nSoy/iraUyc2fnZ69tiexpQEMPGbK/ynr6I8SrG21idCG/MiXPMDuQT5y
MrUZ9sa6kHz3qRNDGZvUICYuoWsKP6izoNcGBy89qqakwY3HndjTqJVBzGn09fvfNDK4+KlgTDKU
P2oLjDSZexKEInXELj2ns75WjLL082153W6vycmWunBsH7TG4keEM33vTD9mbxBjI9akVLYDW1mB
ucXF9Koj5YCoLjlRfqxAimedEnezv/0CpUsaRrD9BCWaDIAh+D8ukPrQv+3o3CaCrzb6lAqb9SAk
CkCFjuTtGgykeYIGKJZX55UL0Cu+nl7b0Cd+UVKTbiOHYQo6spAFqiODTakTAWlWLlOK34O3Tbou
QlX9G8E0s3m5Zot7C2JxkBB1mRa4KGiAPmRknPGAC/Sc6I2gTNOas3YkDcVMDj8VadV7K6wp7GEN
LJ5Z5rwnz+sincseC8FOCNAgQ3gUOy/tlBWxQCXp0fa5F2nagnXVksxO81tmZfh/Mo/Zk6qYgPpv
2wTzfnw7QIAl7LW+jkFe3aYIacIE593V7GYDs75bqtEmLWn2jsPl/h7Vlm62zGBRuAKgemQhjGak
IFnn1Op4p0F79ZliQXU8N1lpAG5a8QLHwLr/LeLWPq8pX1QXvSrqszsCnoSA4N9oa6KbLNmfqjvS
9ANeQTy0hNPFmem8liL0S3eUFGYYWy0FJXjqmRNV9zuXXIsIWS3LOxGhM7VCDvzLaCUIKz7t9LQq
7gymfzxcpaTEU4JwWeJ+gNTVxxajwekRI0VQQdHI7WvTOJflXC9NijvBUAr3vG9PyGaxOr/daUBV
J+WJiahpiK4y1rLe//Gx7tp9Qzz0K0wOI+jNAK7B+g+Zye4GT71p2+KFeX7ZkUg4zDJ9wXRw76zA
lfZMrLrSwwjVP5qt/pmKu2nhTO5up8r3ghWmi3f6LOYLD+nLkLmyfoh+TUqZrnAusHgVIvaxZWnh
rs0w5tPhcGEOM5w9BZU9KYK0yb9vvcq758az+3FHprlvqXbXLiyjhlp7YnwwDOvGgP6SV62C+vWx
2u1zYQ37i+BCb9KTjNTCdrij8RcbFuemQGHyB3gfYI4gLk1Lp6SB3NwM5JijVU6guzvBmRt3khh4
D+/g1zA1CAiRuJ77Jh4rRGtgXv+DbnQvdAyjh9tuPJgjdYkCESrM8aLkMfk5ALHpatTjW1hBJeXn
7hunfjnqjXCO5r3uzHhvFMAnDHBcMSKamoKWpJZQIJZUfHzXBX5dajifdI/Skh8Q2yoIUHK8Jyh2
fx/wHA17plxGe4jLpXAxJ19cg+qZmZ2mWdXkcm9Zl27IlV46anB0svv4uYh/EbA5uCMImprW3lbI
Y2NGFf+yf9t696A5VQX5XgrvU1DyemCwgg7wDxioAFmWQtNNv64ow9DFnJk6IPjiQ2TJq+HAg0RY
r8AUCBMyzDl8hmbaBav3yR14AROTVLswOQhp/LuUK4BnXXjuzGRtVifq3ix3rTykKMN9UJOvT8fC
QJ0OAJ+I7K3S/fXGx018AlNwRCFWvVdmaz0SWTVf3pcPG7oTgPwtOWW+xIC7mdr93MWhbhalVaqH
qpmEgF/G8bxZiYxR6u/4htCOcg8+IZo4+dKjqGOjfN5QIoaY87B7X+s2SY0nWVYTdJyqeY/GxoNJ
iyx813EWz0veh9Fdb2v6fm6SzmBk2Dsob/vmEajR8EZg5AL7irkR2EWLncFcPsBiMobxvY2/Ejd4
R5RnXGfNTtdQVvKt27t6zwHdk0D08TP4sttA/uLRJSkGYzQlkly61i8R2lRuGLy/rSJuiKyYQ8xQ
KfRfjsPZ15RrAwMkicwLKLsyjWMyLmWiEvKzqganjQV3ZP60cvM7pgnq95vgV1sXx3a9p4gWFG5o
huQfCIswVbDrw8P59cxvjPuIS5ZYMq3BPkQ4NOcnON7rVSL1zmtiD0WfEruXLgosHEctSK10OG7g
4w/nW/g+w+RTDWU/Shsulw/UzoXZ9I+TfPgxnHykVnEKuWqrDoUUwU8JkvTWtxHC6mnznxlT1UgK
uT7WtyJcyktvjxK7vXJ8sVZaM5Xtx7b7dbJTLmzLPXrk4SChA34+9aqpOAwlx9s9XBWljTQvRPkK
goTMSB84vt+njg2jQ19FVUtdCExjhp3ug6ZcKSz7fqCJEbBvwxdnF/aSvsZZpS/nYUfYTAH0TCOb
XVzDzz2DTbycGaRNLJqOUr/DJ8OBYtfIc3/SGVafy665nIOX70Ppg3bMYpuL4gljgISR50C9ZCl+
lnGMnk+5Rl0XvFMm/gfHyqPL5OiTxqa3XcnxjNEARotVtXedr38xbhOF4Q1OfBPTVyMvmsQlKKVD
FJYcFFgv0AYiPILzXmPHKoiymNh+Dgn2DWXqhH0dLmnngAqoNiT3VmBCK1bvgwpN+2Nw4TfE1Rp6
0PSVHyBFWZOyTTod8ApPk4dHG0jSN0ryta24boIsyhS1lGicYZEZo4tv6SwkxLpYatscnwsYM9bj
rSUtVISy8lvHV9ZkO3AeEUwwyaRvXsNjxKOKvfzRLLWQrxv+rVPTYtQL1nEz+Z07BIarsH4F+D5F
KXQ/C/+RsCO4rmS5BdUwDenMgzkuLOJJipgycYoBe1QxOhxyKnjS/db+eWPkCzSe2LtksduLITCH
/khs8F5jevi3EMrZEXWRPHYtD5rqEVQAvVXn+saDgTZ211mkmA97Q893VnudiUlvmgbmV3Xn9/Mz
oYlQi73e1JT1vSI67wN81lr7hOkjPNoTROyXquuh9sO+81XqmptMnNNBb94vkJi+dUam/aHQqFfq
s0+YtNF6q4cbqKAMMB0znz+zd06vUEbBzPQUEPgVUPO46NADm4i5X1VjfaKZx1Pt5BrAUSatVfu/
IKe/m2mpXZSj9eUzEwGkoF7JP3DVGU8aceeFaoiFj6JF9jeHL2Ppq4tuly3cfRs2rDlkSLt+sIfi
19/y4DK/3ScV7W6dHsw7MCM/nrkRmLWUjd0XaeDE0L5Wn4Vk5oTvxvJlYYCP22/K7bZO4g+dPt85
K46GOc4nU8rjm5m/m9yEZMWIIUJVdKhKXv++ejTnI/3FcW9PO8cgdILZVkrkTzoUxUA66M6AvyPz
D+2U0wolSqAs92AF3v95vKoK3Jl/SUBADTyBRmpV2dmBhBMBaSNL6kRxKT0jbHy/v5soxOskM9eF
noclNdr0MTTjK32EK7CiDAXA7TrrX+3YYi5kefwGLi9sCsc4qGtgq7RUL3MZsQJD8Q/WKd7zGP3G
X2FQwSR0yw08yxZoLBDIHHXwzhsiwVcD0FyQo03dkadEzZkpt7jDgGvHhV9ClQRj7NpX5Gu0TVBa
iEEBcxmEjcRGa1sln0vD4ovSycjX0Spth80J6GCoIJpcGhNeYf8pl66P7ds3njKmHrb0FX1pmMm6
I8pLcqY/DAxP7CGGzuSQlaOdtHWZSKUTS39SIo0+kmGL956hCxLIUyQK9jr7alr54LLlIpoEulh3
NfjfayCK8Y/qlWtUxF3UTjbcmvVm1OpzSj+e3icFMamqt6+T8C35GFVm1AOP+PbMJQVOGo3KCERf
oz9miTFUvRcvh1RvgZWfFRZJMX8G3MbtX1V+D/0Q8laKvArwPM7/K6Pb209gylvn9KHLhtyH0uMs
zc6kO1ReVGQ2HxNAcNVuSQbSeuqI9N85jn5On5WexXwf12totuUwDCxRDxqjMNp6SVe2D/2DcwMw
rb2OkbAPk0MXLtn2P1KvRyaWkFOC/m0YoXp+L34Bm4kxUznVpna+rp3tUrQY7YgaSgWIr++SXO32
azbdNNPW8NEktosd2TIC/wBbS8qylzvUkrmIwedPijiMd+7VyCPqm/5IBDHNxJIUdl6rEMRiYHCf
ur/zDmV6BIP2KkCahTz+EliHgcTq5VQ1vjqk9bvCRT5w8kC/UnCWOKymQqUSCFm23AgTMMSnL4Om
5Ys7J5Ey8cGLrNcNAp8c6b5DK4LwkrZZbj9izCJ/blbnmF4f4UFz3ilo4hJ1tpUSn1bQFcvQMBuL
hv315ygglnjJtmGY9MJohFewM0v0Z6ylShgO5H0y0UraElWi8voK8kDlLPnJQXuDgnAYesLHl8Iu
gBWjIp0LPZhcjEbHG48x0YtSgRPBJTyw9GrGHenROJ78tJ87yKCevqVxiNVS9G1hNnn4Syc3FKQ4
i2U5f64vCAxK2Mx66WTRpOD/8h6HCYti67pKKq2Sf5PUAGNl15CfgIR3lGrD1F/PT7I0umPgqeiF
49zsVNn4pBbTavB4sKdTEQ2bab+4UWgAFlEtGdLXxVMN1LZf4aQWWh4fTmq9GN+vTnrC5TmGMHNO
P9m5BGG1/PnkLuBeyGFEuBruUww1kRMTayWA2p+jtKGJ2U4F5Nj53g4qCG+2yEpYX44+ckiV/qVM
87C5wg5C4eWItEw0t9zDt7q53J8kUc5fpHfd3mSWXBy8tBERXMibQ9JK/+Waj16Bec51wPap04nH
w9SHszESvK1F0iLMp9SBDPdmfzjyEu+/qsP7vHtDRWpT/AI7yOapfGzaWuFbvgNeIc+GjtgDYANR
UYf+kIx3DW3RsUNycPxr/eeDBihxxtqma0ur73ANQODBTIUqM9E7GcC9kA5uHZVmalVE6sHhsFEC
2YECAWz+f/5fMYadt7/qJf63LiXRrfjCTHppRfiFpSFaFOj21sRrV9o1mbHJh272ujrVdrDaxXwk
IVUH23pNQ+k9TDPIz+2h+x1w3F0+s36BAdjy7P8JmtO4ja2lpwUXkobEMCs5CauNE+ZdOLmIrouG
gzsL0bNzXptNC8/esoOBJ79kmLCzbmaNLcWchpr8yE68XhIhqfDcVIkm1zhuRG+5HgEB6QJAaCr1
veIGSHNl+8TWqKTzAFUTQlySKLg1fgEh1Cv0GYhG4tik3KbhBgKqATgyfIRdzzovPrc5gm9zWdmS
7cm9LTmgvXK/F1bmd98KUDj3R3ZruAYeQ2SZn7vuuZHH3jKwpW7HHZW9KO4MOjn7F17o4QZd/nfF
qJETbv3bT1NXEiNg95pZg7TCdbf4iVERH0x+j16hiIcozVX06vEBtl7W+epvhg53GGkolexn62Fl
orw3uK/JR1Vj61AQ7+3DK8z+adGei4pTh+0aUv1Yvz7gxVNigmBuyF5OUwkFgbdw7J2Sl6zUjRo+
EPsUp2tcnz7Fcbr+3UKm5pSDha4rDxSiFtQvQDFhlawGofOQLyPBSaXehHho6p2Jhy8GGiEBw5iu
gJozTsnubF5H2fDGn905w5fhoKugtpgL3tEBvc68zNTZnmP28tqNyzD3yQGCcv7Z/RbMWH3rgkEs
FtoeTSV6FMUC01PHCMFbiNTqcZrG4iPuezWOKjpz090UtCV5MBeLglgCkWO0DEw/ZA9Pr5qfjFPs
v2yA1IXyqB/PzZWwRSnckGRk3tdKW6Kr0gb+cVSg+sYNs6iiuWQ1sCewwhlGcoDs25ZLJv/A++34
rl431MKiRbW2ngepAKnns4xra4aW46rEYSPsLgdIZWWq+yhJKmDMbdYNRjcZw9UKcvtPXKIp4kLN
3/jAbW6hIfR5e58RdeAutQslDOU5mKqT2m5zPWRTVczUXR+p66UFblsssrM+xZByYKELsHHkI39+
keHiGcWBZR0kj0/egoPSR0bw0b+Meu4ZWTm7Dis3thfmKR/7kCFsakqSMxY/LCxJZqPSKM8NEhb5
cCv5gcDbzLactghdr/Na4tczaQG+V7Mo6dFTJ2zAZm03LKGcdbaxiMcDdFwXRMqFWJfFqZIacMu/
gqE0jm25fKf1CHk7UwTslamlpToubTUesFeq/U0FOozb0JQYjAdyOx7nECeZ/J7Cb2b/i9Pzrqac
haLjEou/MD4exkQj2i5aG0gy7e0+z9Y8f401a0CyXBLK0x6onmCqGHHA+bJFsuGh3hJex3KtA3r9
z8oglE1U/RW39+NJ4sPrTTPAUg6zFFa2TFuRYM47CmQB/gMc1ruRrTcOtLnU7H/5j+ioljK+HT24
kIdj8c1s2KLJ3oMknWyTK6vW+RIBRk0HFOmaOLHhyKbieU2djkX27lE7TnOQPGlq/781cRU9dL+w
Ve8RLeF23iH3zDW7USrl/p8Zz9nfk7GZgZvmrQQqznaPODVfKJDdr5dy9u6sLvmxKok3sxQAgEOV
yyUYXoKMOnk2knRep6uauaEYi+Bly5JVN/SNRGLiFIGTPaoLaoX2sj248z6zwJbv8FUvP3P8IR/E
bI8e6oVbXDXuA62gc5sCS/6WYm2DG76McRzlNyjiAqHlXwgqkzuoIOoIU+uK2kTASwN+H8EcSML5
Y9Jd4Q9ZDw8MJ6a2iBSTiaaMyne/KL3o8xNtMZQR855XBrCD3HlNDdTo0PXILbzkx6eflqkT4goP
uLs8+rzivWHQ1C7QO0xLoNPwcK0djYIO0w+XDYWLQAZSJvRlkoIwxfOylzwo05fl1USkIE0n8rp9
l5k7Hm9Mt5+e1fAilxJda4rG1LhlTzWfRr/yWYo5ZusJfw4HlVS715pdPf/J/DlrVHRTJOgOQFrI
FFkSTc4Z2KIucDmvyAsn10RCXEFp83jyWMqJyCK08QSxHXHdZkEZ56Ot/ObESVtxycx76ohdMsoR
BXzpgD5+6fsbl2yvDAxsfrLgA6kTXbQ9ZNileWDS3e4w9El/GG5vuynWGVM9N+H55J8i933xJplF
+vJpJmmDKyRHLo8Bx5O4C8Rzc8UNrvFboyUGzKDSupXymh2KnK8Aj6rgh1AIhnVtR7CJZl3rhZiJ
n9s6z80IjnR/5UWOeVj4ZbyuvqOxyTes+DqrqDLcwhtKtaTW8SSnPP3wICjpvAOcFnM2EcKKp81g
2ew8EriMcItN0P0OxAnbu3cHNkTJrnZwRLGrpCMNV9bHCa+UM3mPJa2iFS0dMbSn7EhATOO1brJa
VAlktZDX6pDIyaSTSJRgvFwoPmoR/K14bo7yUTLaZ/tiH1DxcP3yy7eVJhsnLJFiXvNqlFLf5ehj
Mg5IgsYsHgYRganpVU3D17+iRg9mPWJIwtMtyRX7xaPafRKguxQbzvMg6Au1b/OS7YLrWpa5AfL0
h4Tx705uZWPO5dj01aYfhRK3K8UGJ3PtD/ftB1c0U7342T1klKOb7xgGnindV4n4q0DZnw7k4swC
OViK7Ic67ku7vlsXZg2AWqTNw6Im3aQOZOzEYT37fE6P6N51uFJ8LcPKGqDRB6NleiftGDO3o+hs
TNeeU8PsbgDb1I9jNAgkCFCQNIEsp8bOh0GUiTkwQFTzthE/CL55isn5SrTVOaOyR8y1aG17UT1s
sKCfZ7RA7UdNGRvTakX+FQQOPPnZdBl7YSzTMCr13CPmV22rUrAmpoUwNBrwOmbhmj9tqIkNZm7L
gnAB1bIb8Brj3BBEWJyCPKqKU+fj60yLXlsjCwGJoiVX0rbGfpUm6wI87bc5yTC2RfrMuRdbMX7d
6n4XQKO38DK9UtU8a0FKhS7HkWUhXFwCL1UCKE/R13sHHrplSCxJfQYq8o32VZ7jBXWvxCurOUis
v/1hZfgasNlitOWXWC+6zBur2v/Niz6oGXCNBhgBCuFXN1zUfQvRi3Q7+OqoR9hTIsZpe9r9aRDD
1l1qKvlsy3vduknuaKCBVKJ/gdVOnrVtKoRMviuec8/oxrZEZnJkLdS81upZq00LdMEucXxdp0hz
ij9aIRojPq5OmsSJkoJt2nlW0JyGOJ1l7Sa8Y7xSmBq5rRKL3HVHbnEsWdozur5/BpEFUXrGFWRV
I2kobQQ8HaeWU4ry3CEq183aqt+o3bSl5gB8zX+uCi/xNWZKzywYy0hMo9eREyEZEMEI4uBRH4un
6nyEfbUCxMQ1o4qhE5D8j5Cgy/CSjykWQrmiTNP2IJf5vSCTZR7okfSqeXQo26MLWJ1OtS/H3H5A
NRD66kx1geZcBmbjxLijW7aiH0J7SPti8T/FYN6rBnp2+14z1uES1/avw3OB8lSw8JgyKxxB4Td3
mfzcv+lgfQuXpiT3ko3YR8+BLptfaWyETgQzeKHwUMnKcW7995rr0Kk/T6M7AxWL0ldjb0faiVyB
FHYoLyuJPotNceOEsEEA7xygLoUz05bOxM/bncJVXHl2Qeng3drONKEYpTcPGxDE4jWtyGk4QYBz
9orh9Ckvbz82pZXR/WbtGXweqgXYLV/2CQOuYJlHrVInh5euyt7iS2/lbC1mcgEIuFjTFU+i/SjF
h9wqvPhgQ5t+PSgPFIGAFxfQZEIw+qM2YghSfjVhaN7dr8ai9opp4agG7eL7lXTqwmhz8Y8RauEr
/Wlj7mszNQ4V4G35M0Te4O0ZqqjMvhVvH9SX6Rbq+ZL4kiQbIfn3rbfJSvcQeSIbRI4lD8WCEfTu
OL5wxDdxKwQxS5Swu3jNI6kMJil/zhsUsJhbcvnZHDeLL5LsJz6nSkYUtfqM/l6r0WP0Af+C7Xv3
Z7eviTVEcfcuY0BqSFaYmR3VfPkSIaX32YGtwR4PctR7lVGJd4R5CgC1CaTXguypnLKhdufstIVH
ZJvd32Qv/cWAPOo5prH1eFvkbSASWHX7leDjgZPeJBrbKk/BKFX/D5TzyDVIzfskCF35ZwmClZCS
5DhS/Nup/fDSX5JlSs6WlL9ogiDJbLJsIjkwCQkeskinz43/xv0k3EuZQXCh4yhiMf/yYOG90oYc
f5fQvufwCG4wVpSsisbyr+C7xiYNBXVKRUKxPB+vVmm8xGXZi74VLEP32dBNj53W+PFupxFVBq51
X3I+FCd2ueGMCkvN3B8lECuo21G/Q08mMsIqSDZP+e/AiPzyN7aDIVyaK6rCJZ73e/K2oxNMcM1l
t5b0liZ3cnZJKoBgE/NvyZkLyhvgTyljsXYKkFVmu1iPJ5uC0Rxa0UOsK4jKJ/085qTSRmskhqzN
j6UOWWl2NIVvaBI2oc0XxmfX1cLGTlwwkzTM1VQ6v45WXdUyF2tCumt1MgStaNJmDeo+YsszyhfT
nxT5eYT7wcQeEad8W0d3DtfBlke2urRERoXyGFZRwX14X6T36dW5m5tIlgGNiFn+3gqaMKkhsx04
iHTdn3aD7LijNIPowQe0/5xiynrP4k17CoaC5d0HajCuog2a8Ocd/309ISX45F50eRwWXfc64T3C
SqLEuIVB/k47Ea2BAymbAjRPp568hSBr4rbFMs4IskHLqkJyZvR/ZdeRNaedyz9XxdO07XJa2tSa
3MAJtB8XyoaNxTpDGAMnFXTrtJyOpqeRqivAnv6mBx7TOuqgM24vorF2GtwZ2KBkDkE5AuCtqsud
hiUbmqWQfG0giN5YkhUfw4fcV35YUq8iV2yGJ6MgIqMWiZUiasuDNbdrTD+HHhMc1KNckIIa9i0+
xnNJ1B8MyD31IqoTLDqbm0z6k29x66QZ4J8ywfzDBtj0uoZTqFkXKmB4HmJJF1ZtCMHXNjAZNs5c
8Ao3rwSDHvLF7uBNRBhUTxBQxeADoRgg5JNTLmxGIUWMOSkQlksyYZBiPQE+FDHLbX264oupZ8+C
rclf4UDqUOZJSrv1uWdpu2MkdY9duCX/eGbRShrEBn6s6LX7IS5XwvcLfTqpKyAF9TyijRm8crsC
73hUkP3g+yjqt8ZFfJTiSgylaYyYu5vRqBbP/j799qgrYoh0AoJ7lKmbgKOcDsk564iS3pIF4DOS
i4UVsv696CP71iZT/j0hg9/eXVQGfHCM1QSBP1jZBDcPH4zdR/GAiUO2yeBoV9xSJmDAoYxxr+P5
j3uCQA+xYTJH4FW4FykShc+24rEVZla5VuZ4OP5zwnbjBu4O5VxCXBPtROIjBAwNOpfUELe36rzF
sLdprutt4viVIeZQGLe8sIlakMO4RpHwCWKTk6z1E2Lt/wNBbvvrxZf8j+oiRIBKV3cGcO9Ic4rk
ViO329M5milNnBKtPFopMCA+/QzK7VxgFJAl/llHne79M1hZo40VRs0aEl5IYaq3yn/bWqU5A1oJ
AVciGtCIKH2PBhtJhJ2IP5eEurIc+OAGq5mLkrvyIQMAqAQdA6jM1K6AA8NHj67aMqFK9CAF6q++
n2GDKP6ztRbj28V7iPN3sNNXZNtuUfesZYj5rYAq5q78xNypMhlll0EiKJui49gRYQsooYV9CBSn
x24e73j1dxAiSnvwguxp+/6X/iovtpsY5TdwazGvCsiCAzZt/ZtPjZBeHWV1PiRuEBiW6DKpUyWA
JoYX0KHdmK+Djp0Fd9LcX9IPNME1jHda0W6EekawBCMbPPnUYwhFrj8atz7PwdzXq9bAMwKVGV5b
CPgheBX7snGQnFQFkBv/s9lefSkMzIayrAN6lESK7ejoF3Uh6OGGIygUVvkkmnZNjTo5+vssrSyf
zm+Nez067+bqWN2qtV+JFE8XXhtpnQwrBOTepA56Jgyq71KVg+uIRtfbeX1UsMkjhdtAjwl/Z4OB
3Yu0zsf57PpTg1fHh9cfdpmsdmTM8tVqWg6BZvI/AW3e6xD2e77TnlH1G+2A7C0XA+s5tt+DSfdp
Q6dpOcz440V3k/XX/ptgDWXaj1M7Q7FCI4fIFBXqOEWmtsvUfd5xWVCQmWrPSIJ9W7fDvFfIWYNF
mh7E04UYb6+S9Ja52qY8UOeIw9zvMqsWxCmHtoInPvwdAUfdmJHbVVtggBUv2E7jS5jQiLhZtUDt
qqOD1cn/jqLH40y2kgW3cplGUwyHeNL0P8d7QHTRvLN5p3ryHqtw49OQawKVIpiA+E7fAqruuWnJ
Df6/xywm2xooxOXdSwl5Z9szY8QCP03iuaPQUkE0JXgTv8zXeygbIJZN0KYt2/GxopzC34SyXV/C
nxzHtl+ol6pprjxSWYWqZl/qeO9+UlKkdp7fgnlafnrNIVoDIS9LV6nZBlW59pcA5ZFlQaN/QcFl
e0imCN3hs+l+0dcSkggMIviqchYcjK1BzMCOpHnO9BpJnjWwSvM92bzb0iNspvJAmwbyaHQVTu8/
lOBLgtKLFxs9c1wMyT+u4sobobPDCThKuui85YXb9rkrotKZMYVJ+eaEv8FKJJr1rHp6+/QFUWB/
AoQnndoAHhGeWzIgePXmYIFNh1dIm0xGiCH5LgcabR6oYDZs86WuYVZhCM9cnv7fqCw3IsBF5QnT
pIpY7tWbirrSGRjdDM00aMhfLuHalxNF99fJIAVBt/W++yUEfGIlOU8IG+FelXMduE1Nv5rdoBun
PElcVZ5cFYBW2Zrt8UW+nPEuHX+pRC9NJe1H7GDX72fM5M3LouwhEKWqbbVXJhYn0ARF/cmqmxCc
vmibBkkkbs3d2H7HgwQyJzBEySakDJ0h42YCZa+AT7COgb1fKRHDPrrG3E9CkNmjm3RqmJHj8tY9
Tb0u57Pvrc55z4aVZs56/uGbpAzmHL6DmLAoKqrbKqfIWnTFHMNhFtBQSM8/adoDgC39wDhwRg/m
Yid3ESFepgWvZAed/vx6Uc3wLgilnaZIgJpAnOpZWP3JYxDeojizw225HRuPZDayY0nqNFcD/2QG
+63s2jlHS3BfITMNtwS5WFuEfgInCP2uVWUih+Hkpz6TcSVQdho8LiF5ZL/LLM+G0ndyqBI4MCIh
Ej/dXjz5ng5lm1jqJdKctzrrE185Vp7degpYwzDLomffdPkm5oLb6kWPOyJrxBoNtIGLFBS3tlKF
lpgPhq6WbxeBWfZT3s5WwaF8LldcElspYpnQFEZZIGiBxlRk9CmHTxXWVW1d/UkVkteMfXGVU+uu
UmriAh2X/Uf0HVd0xaCy/M2bK6hb4ksPP719AxWBd6vjZC2UBiQa5ELFxXyXcDE5ARJwqvJBJ79P
aArj2GNSlzSq451afa+X/xMM9Mb7tEyQbpTgaLyadKy/3j6KR7xip3oLPQbVyfCSqM0WZ49VoufT
TFPC1hmwsDIg/eXf6HGjYbKi/OF+Qxli0M8e1TrdTcKPexGZFHJ/fV457LuNGoq+cL5ELGU/XGBQ
u7+H22xijxPMg4VQR7G64+7ZU9uUp6rjmp2QCmaHFv9ioWwuDjTE41p+SA5WRFgTXQzzYaCJF8GZ
99GGSawAeSB3KS5yF4bJgtPqot0x7UqqwJm2Jr6FbvUCBRJFLhBsKfrSd0wo8KRakYrjJSmHGYxW
arvn67dl8Lo/mOeoE5fxGnKVTKt6ESyGIW6GCxeACkno6gLVOI55+vHfEZoCY9rafHPcrezMKS/6
fX5sk3iWlJHqB77yqA5RTLOkC+lIh8pgRy/XL4koNKjoMrAsY7TBtNFIdgaUCfhWM+Hu5AWFQzQy
DdhFtOjaQYNw6nSOIdyHt4kXZECwGpHaR+Uqk+f+pT94r6xM74Z9yASvlMS0MUkM/qst8G343wXM
RPYCPGqwx3lFLGGZVuDSgE4Gm7u+UY9QNxkPJKREWecndnUlevbnv5Yoa5hdBlxcJ4g7wlM9mbY/
vd6oW2WcvzPXJ+XYfhuCt1J//PqMeKUFxAcNy8SL4BBTNJ3ewOZnxbMSJYQlnXSR7Nes3I8auDaW
DffbSfmki8zN/NyaslHVSx8JiDD9UUpoxmdyrJ+IVz/U0m+rdLVrbkg8RCa14eYpR07M1OeWaWX+
zpDTDWMB3/1jieWKqGsShhZrnhXdUK4x2SQ543HgPLD8VqiKVBLgR4kjD0DKpjeQ1ugjt9ZNvzmo
kLw3QUulL2SyQqVdO8Q6fTEKk9MNNgaLX6OOVfdUrfzWOWv+btWZb9gXHe8pJE/4xXWorrirENwO
cTheO+Hqs+m3orrYkRke07d/bfFm0OXbgcJNXXR8hu8smaJq2gb8j1GqUuAmIx953AwiOUh621ly
WUhMRa3BOWTZldS8xWQpKYbvuaKm9XC+YELZ4Pwg1x0g7bNkQPGVGR3WdsW7w0LHGEgxx4pgLKuv
AV7jXjMI1m2VGhqCUAsl9FqcjAEg2sMLfaY/i2D8XlGZ5kYSPvoF0e5SoSesmIDCuQ9J73hgXnoc
YxPU4HmHnfhlb9yh2ZCtLMlzV37/HMVVVZOiyPrT9rudRD+ryk1A5xr2+IMlHdKwoegjZpPPNpPM
PPxtP2RdQlSD2N2Lal36LKvgnZ2JU/JltkETYmuWtcznpnK/7YFnJx2KJHcoQ0MC2BHAKmQvKQ+a
uwlMuBdHk89Kodfn1vCKLG2gZwe6F4eThhASc2Tkt7s2VGep8+fkQ5Xq9nqu02+rs19RJf4Im7il
XXd4Xi57vMFfvyRWBayNOz+XJFK8P90YSywRkVj4qJVaVjBRPlXfIGisLIdDFxXoFfT+g3PYQ35o
RdBBLbh8YUHlwgVoIvkqeSw3FTChq/xCtgrNjdz1NIyEMgmmW7VlX+IK3WXwyNdYXxsRHZN3NjS6
fX9TTeFCHLtflDZmb6bhh+xdVRMsbzxDZJ3Cr8n0yOgTfTFxlTOpYxQIzQbqbwIXw9lfjCSuF5MJ
wSMu06gB0eiltcwygXKVFqKdnDA+am0T7d+yOyam3T/KfUg0Y7oB73krJuy73cLY+dXmnBk6vJoT
uSfBVBLY0aBsM1gB1l8UJ1E/8GKomuChDvL7WhT3iChxxyAiePpZJqEr7Nq6tfsAe2IUhNnBB0RX
4aSEdW/YmBaJQfZ4kZEJzGzZEQLzh2L2PfMAPWseoj1Dg7D0sVJoun74xhMSmxSDQe5ap6Pdp3uO
ctv0yhXBDd56Jw+ZRu7PoAOejKNjPGRy6VSkzrb9jGXYpRKK2CxmuxznTJRLQ8BSiVostQygR7Dd
eCN5UQOWO1VyoosANb5LhdX+MyHJD5IRckzLBcrgqR/tfPAq4AJoZcaQzbUL0jMTino/LMKfJeGM
5Lbi0AceU629wSVDnIzN7ZzWBCfvTB2Ac4wkr/nnupf/1hKZWZGwhAGpxO2D32Or++iI6Dhx4lMp
JxhWuxX/QIubHhPF32L5MEDO2ctaLur6nKmAzPGz2vKJOQNPyI5d8VRKhyn6F0Y96PhnzYeGq4tn
cN2EtaepY+cAMsruWuhzm0uWQYyRLlieTllu/jfwe5u7AznHVbsmCM0O7ugTXRdAOu0X2ThDEPyA
/i4nf8ltQlSsditddzjI9Iy3gGMZ7ObrD59iOvT1bnftKfg+fKCshX1JVvnAIMe8NAU3a1u8ZGSt
BxB2XV+wFV2lehb8YuyhZNQlYAllXruXIG+dPtqx7ml/1v9SAlEmBWGBuPv/OvoW3CwRxa9v5J8J
f9i/0g9UPjyDQxKmm2OIGrEWWGQqh8e7Nah0pRg4tRp+MxdidiG8bNeY2+9oe4PRkAMyNyj6tHOj
o12WUkZI5nROh2G660Aj9U0Fn/gFZaQ2zHHD44/ZO2K8Zbmirl+wL+Uae5JJSuE10TSDfM+8/JWo
ygkezqvjaL5XrtwvESJvAlABj3JutN5al4fmeeEB8I+0JVcSj4RhaMN0NPO5dSgTmALyzo5dqO+d
jJ9StyQkobiHvP3Aw47Ju4S1/cCnyezdmdtbk/M8ox/DR6mDrQN69fhPR514Z8XNfiSqKvn2BA9y
kkONsBzyseSwfbeQClSw9nD74pz/Q2fkMUIBgZGzok9/y1o8OQ1tjQ0MM0IdzS+ctmtmnlYZM26V
0icuuSl/v99MnDM0qe3YHaCYAj3JQyu34vPam+XuS283WffKchasUuZkaOBt2jX3CUZZtUa25/yh
Fpsm6kBdwQQZhv54GI4AXJdX9FeZdUFRU/fqT4J/5F24INUNd0AWNcQLWdz+t52Jtw8RVvIP9PbJ
30thUrWqlgJlHLH+EhVyFVgxxj45xzfEUzQe4FcSIZKlCRgiJ54fYLg5hcEfzdOqRuzN26e7+xpS
yySkybZTolM4o2O2rocclfs51x8BLPvuySOz7fNnqaDcluJeMxPEmfnu2KnLSd5XT/b4YCmrNNp/
WG0CKzKgZs7RbN1QYw4qJ0TUfCkZ4Oq5THdob19UfR8DJKDMOGQsr9BLtnGihD2Lf4zzKXH/tWgD
z7pNLj7a3k3+SDylYKufR+7XR7EEKXdQIfKqfqTJp16PD8AEdR6VTWuVxSzxKFk2KITDzYwDbkoM
Cvbc/DjrzPBUSQGgSakAuwp+sWc8mHJTVxUHXgcNy8v7Ykoq2KCx5CuTDrME4/7RLK9oW0f11HSn
e403YPgzibKmd8KL0zpEc+CKcvf1R5UznBoQ/33pS44fXgPGGNDJbIRSsE924MsT3R1dUEl02rgF
QVUgvXyaD45KTVvqO21BjwXUtp9vWBMhsafeJFnRsGZkQYwZb5Loh/ba7ihbx4hH+zIT45UZ3LJk
NvAJYDZq/H08RRWAF5mll6RVthS6+KgoZDnSJLawRxCaKfYyeNHnk53FrPblyfIv5mPzMUCKSRt5
gqaTV+pRI/rUIjbcwxNUiT+ZAxX1/ywDwf8srHrxBZcdJeNTKOEetveVF35DL7f3x/ZX1EC08uNj
TqKNxI50VxMDmXOo6QdCWDb23xlthAVAcY21IvAYPJWoTInbQCdVsPBkczBA7UMuduegEn3FJ7y4
Nv9oahJ9hnLzFFhm3EXM2OX1H391nqCFIAhQPD6wNqh0Gh3hg0jr+IJ/5ZHoOOz5Qigsr18VyA6d
imfaPkfx+xt9eEpwwGPyF3q9QXSiYHvYN7MQxin7yZi6w9pkXdjmqJm0jRXXSGu9R7etdBK0Nelr
j6ZVFqCAIVzYBL9LLjW1s9MaqPAB81beRZHkHow1I/5Pakn4quPhdnb5oV2sOVumXMg+6EX9bsfN
IR8kU8E73tn1wK3iJAo7Hzjfgj/3qgoa/gNifBfWuivCmq2jckA4fy2qDUQLrjT6tz9O4U/uNYBa
MiHsqmJ5h08CPNpqfRPZR2cfqsCM7oMxfAmcKDqtOeaYUbar9xvK+3SD2Up8pAzGJPODrFueRdvY
cxi5uPApeyVHXckyyhzHcKtHFyzSeAag7EzRzCEKY93yxxafRSmzjOO/YcsH/MpMsGbNXb3B8Nf3
YVs7wDXP86hDDsvODI37dT6dyALYK1XjpikQ/3vpjXYhDSUX0yMRuLAX79rpQoL8fxyO53ax5k6o
EIrcfbg3ubXyi+1DISDjOUFmQdA3hRPg1XLrTmShP3REqoHQA1uZ+qtnNmIlMyFUozAPOR5FjFki
hQnwSR3Wmx4wIx7pED7ylEKcdZvP6HGQ8RM9StHczSBMdMmfoxGHyJMQew7HSQdp0T3GJqclBQR+
wa89K7Tk9QaY7c+duBmB2ZJtBSvs4U1Pp9idUx5pNGJC3a13yCVVDHjerbEoOoh1cmFRsKOk82/5
ofmhu4Zy35cn6HFMkRE7ZuZJat7oKwqWRXabxbSYZvGpRTVGUFUCmuxRVrPFxDfIThFHwBIU/x0i
9ApVpCTl4nPI5B80s8gGO+EkTm2wtw3tfv1yOBsiUY3gIsluqJ6PfAFCnI6ry7CuUyVHCluExrxE
APSzXSFxGMytuY1mGeNxgHOiSSBZjnVljnl4iqXlFO1eDGDn20KKTL6n6F3f7h6ylq0fQGOhZQZG
Ev33+1QhBNgdhHHwRPj8V3Bn3BiewjdyfOltzszqEOqsBEIoLDbVMIrD4b40AbwF7sLWjDNNx/YS
oK2cmkw6umUR9Avwo95wEuCccPte2/ff/13R8Q3SNSo92ANGlxT41pf9XWQdJy/60z9lOKlzuSIa
OXhoxyD7x5lMCkbrdvctJIre/kDK2qkcxNxN9BgEFHn2PYTi8hJmv2v7W6+meylCg+0RdjC1D5nB
4+bVxm8t3iBEKH5eGtCe5ymVNDteMtl2jmra2lXjMrj/lF+AVtE6xsvExFuw9uMgpDCobQjPCOdF
UTO4FVQJO40YICv+KZb8wwXTcoWyzbVF+W32skArVbAkPBWzlr1tID83LuOHGUO2l7VO1ZbDyM9x
kmMq6rLSv4GkU8hBo4EtoAs6lacZCBX3u3PKXtRsnT30ebc2ghkLDt15CQJ3JZhHjq0Ou/ijUPFh
MJQJ6YAGg3SUGUUT6MCmG+KyIJHTg3TRPLWFMrVp4sF+ZZk8hOSTakkcuA3MMsSJwvuhzgrd9XlD
bTi3Q84jEU7dQJCdJ1C6uYp5IDUr/w5PIyekvRMcXd4RvYCPPLZj0ODWEyONyH6lJ1AFBDbgN4NO
vdH0rBDBoSNt7dzWt7jEvFI/r8Kz6LVxQXgcQpu/Hdqu9pfh75x5NwnPRa95uLDGdTPdFRap+0EL
9HnhDL/TWnIkyJBe+BOJ+ZrF1LJBwOS0JYemmpdTQfIl0ZjHK98QG7qcF+ETV3yMG4680bALOBHA
41sIU5/qralwSn4N57QJDNQl2Fom0dAYLNBmBoEE0pRqYjkEul3CfpxGa60WoNcsO/Wpasu6pOrf
eNZ81ydxiqM1yHIJgjJ/ad2a1E5olD9jKsnEU70zEuXzlenEfhosHpNcZeqib2ix79t0hEN811GQ
sAC6UMeHtBDZbw4gWUb7OMuj4hMQo/QjUFmsOjGfhv2h2NVWKV/Z2fU5gIWQ3m8xULrNAUWgVKh4
75okc+67cfColSUyrN3EgBcDZJiUclNhABrunJCNO50usW2lXpu6FsoZi9ULUdymFzmfJ9F/rfBF
UGeMYazN6a0X+5Im/dksaJybwUUaUMv/XMaftaKjTPEo/y29vyNOmGjG9vErMH+9jXwxiPkTwyOn
fbgSYTeKZxKD1rLp8PBmcAMK9NWm8pCqD8Zab77QbaPo7RDFRxoZPVPckbafpcnM2OBCKptMdMCv
oVl5kDgLL2e5Qb1fS5EE88NBwZq8d6pam9umzz0fOuuZry86ZYmlHvBIQhgXHSR4IO2DR8b0N2YX
R2yxC4KnFkskvITpAxyeuUXdZxX++k3B+OULUQX19gvDWTaNtZ/l8F9CqW7FjQLbk4NStKJ8Kfxc
O4D/qqdeJeZO0N0rSNAluImnDuV+0ng7ZnjfwW2cnss1+83kEKJQmNWMtN7/y6woVPLyYV5k0osk
mKyJlrt06k1e65UHDao+qoTwNRP/LjcHcsHAp6p24iZiIDQ/0pztfh7uO305+8e8AmqJWasa7UI8
AA1B3OVsz+vY7q7rEKaWj/rNFyWT6RsVKuPbhoZWSMndSKB9mHMRIw+knMQs0uayQrbQXvne9TWr
0TxmCOcu5m0Z77fGfIWOjq5aYqsDcyQ8Yytwp3FXKs2nfjaJrmGP1zpLd4ss4lfK4HZ55ksgaZEM
KiOn48SDcWAAOwX31pr2FymeSwJytDH1JNT9TMhQKqde0SAwY0dWxI+Raa0HbxeiXrw67FC9xcS0
kZoNu6VFHFXWzLRn91KaGTrCjeXEQGO3Tu7cScP/U1dklCJhLkjXX3Yex0PprwVs5gDhqP0mHxbG
YXMGoqQGLHZtJwrCDMxcOuPnUfAP/SYhUI/Q+FogRFTyffPPSOk9dSs+rTXItUPiPcFL03o7AaFg
nNFS7WTLkHIptXMzTQnEFaCAGU5hFIxClkesAYkCyH8DFrQ9V3cBXlZnfEOAVbyIv3YhYFyw+BnO
XNT8SfHZfVfQE2P0PV9C3JQwWVLss8hTJ0H6VQCTNjJhrwgU2NZMaOcIi6NWj2oK/DiiItEUT54m
ntLDd9nwn1cOQIvDR2DlxlC1kibf6NgxbzQWZzdwyZD4E84HFExPrAhZudr4oimsPXN38hfV1Okl
1yHyYDp/awcCNjp/tA/RJV2truhtIdbYjMPS9fcQTCrZlhE/QXyjNeW7lc549mCRCyHTeuzlvOlu
kU6ZkJgSnTyChrd0KGX7uH8gAkVORu65IBG7jyMiLH7sesgWjkRE6OXi3a10EsqTx1UjjdlznljM
W6SheL/AjS/ma5VKCyqUvNSEIvXBWY0x7B54bJUopwYRjRK5g0Vrw5qcC9/roY/2DuKOGmcgawFY
rsDNYEPMvlKmQ8+Fi/69yHxrpGPY+I02YXupI2hzo5JbRd4ujvIVzPox3FD0BVH8KF8nTSZcuGR+
nFM6f4avakwaU77G2uN6YxR/a/qpXxFES7iheQQvC3KEFnyisW5lbDjA6+pT/+Cu8OcPYTczRRbt
Ns+GkziLvlKqLfLYkInIUQMFO1vNOlH3EsIvbfa+AnV9tZ/JnIyRLzMUJcdxmnb3eQXIyO9bgT25
hsIClaffx4QYmwgwqoRtei9467GITDf5/B+jUVyf9slIFBRiSXpiiwmiNNjLaXvUI2WUrmlFoU5H
F/o5W1foblxBfBmek62pjFLapz9zyNWD9hbJJBXeGU6TyCWBzbkV9Jtxj/nkaBekS8drGJ2q5ds7
v6EEDCbBafA2MxRDARtp8aMkMrPttJtfUYw4YnXFsYHt24+DrbMKEWrr6omJHsOYCcfIsqgPHKjD
s8Z3jvzXpa3jhCutoXr5xtbDtxFHenJiQ3RONX3O8sNL3HVE00/uc/3LH00uCIGz24L9voKPrjUg
WS2GozE9pvpYDWwwDinZj0qvSq/Fc0TF+VgDFDvuOIvUv68azgNKR+eJGfoo4TRrOpRfwokq7r5g
PHjJw3SpDFfIyOwvjnXaJuwhTMw6DOonQj4T4fzBt7hcGxHPSlAEdJdbhfHfYVg0Nz6VsY72hPfX
md3Snx4mshg41CPL+nbNmsfQf1ufF0mZ3Ys7KYOHrVcc0PVjfAXcjlxUX6DnsVtl1RC9gF5SUHj6
FNkyJLIzpZjDyFL8F/8x1P+zOyRtUplsumS+Qh13IEJ5zWLs6adLMKXwzXWXaLAcPDPYxpz4Wf/r
FGdXJt4dF6i66HC7TmK1N6Xc6O7qDnrJioNSS5fmhAih2KTGmNSDOn0IUte3gb7C3ABUqv/0sR19
Esb/DEEKiNrirHy1v6Xpz42vj9hdzuT68gG1u9hDDU8bJ6efrqmAPHq7xC2dfvEeRE45xdIN2Fjb
VqjbyQVko2OKqsSlwtur7HXODp0hCqB+USK/qgc8aVJnFxPOnscq35fXpb9uwF7t3jzs2vvug05J
mKm14GXkBmf/6+7Bk5tHIYXlIT7N0BgkuxUl5D1Q6saYF14v8B5gxlPOSDuCW+sdiVAu00vvAT8I
RNgk7pg+gNpfakH43cki8F26EaZGwZYxC0st3OjhcgWLgmayxatgjSXNFwPe2P5hPsgaFjy/LZmd
FfZzeog4cLX1TMygD6FowGA1kdDYK6vi1ugmGsDI9xFfzZCfsqDdaaFaSgwJFLlZVKe9vhSMMi7V
+S4QPNiiew0EJx0B1/ZKHNX9ynVpmBLtuvd34jo6rxT3zHPHqDAea1Kx1kBVb02IwtfFUnJsnSy0
Fzkmfn1+FVsM0xuAgM+126jlQKSSZS1ifhtrHX5Bj2HYDRGv4UXZhgr1HEygCcDZPPg55CX04Tir
vyczem1NqseOsuEBOMenlrSnQKrpqKu4rlsnYJerPaE0mwEyTqGWNxe/QbasjaMs2YJiVmKnxshD
CI5aZVxvBsFXskpIvb/yHOquH02MwBm3Al1XNqj2Uj1fZDPmts8rqTqy0pxMT3ceDD1NJ8pYr5/L
CdHfBIPXOfIx9khg8hHJabLQ/hrDllV+w6GlEbzu614YkaTqCFnp/YpPiie5SSPR65PAJH7wW9ZG
Zkxbu+LbimHqxv0zE8qRx8YwfKR9OFGjQAfMl5q3BCG3TAl8bDsqlx7X7F6GwGuX4IZexwkZg54z
1SXmJ7AjgqNFliMRRWtE9DpYLlz5HwvyvVYLYfFwEDjUNEru+nxK65WySxNIuLZHaZbExdUtQDah
B5nWa9DE+30yXTNbeR2kQSeKLZWJMogZbkPiN6RftbEDb7pG4XTuKytOOD0nWQDiWT105HBjGzwL
971nIUAM7omxm9oTRTmTpt29sgnWodZ37unLZ3C0H00T7W1vw3l6AJOyGciGb7YeQAvzeOxXnfQw
hsqmb/UaBN8RsXy+6ItC32YVFpCohECN2CAwMHuejf1rQKnyJ1o/RNIGHZgajqtE3SeJBdyU+gdC
d0XFa7IR2e1pbGWjBIaw4cxD5me9ArEmBTcFfa7753MWbB2rmXxEYHUtdHCeBPQ1uLF0EOp3Gkwm
e7o8HnBZJJZ1mraBnvlN781GrUq3YQLa0VxHm6LVglSFO4Cl2J0ntJ8nLrc4SWNaso6WE1iqKDTr
fFAtUK+ai0CuPvl6gs/9Av77nVjztS0pQbw8DNWIxyJKzhYycjkabQ22t7mzj3m0vrZY/nmYfGX4
VgXwyDu5d+EkJ24fXJfztRRa9B+N8W+JmCGPTmOcB0UGNUXZXf4iu2ctj1tSe9gyo89DChldxl3D
B0G6x1NjuviNyspso31GCqR6a41c7lPuNDWeR0f4n1GtJRMvdVPXnAKT6SGZxBxr/+LDBHY0hsz7
ruhvrXl7IlpmePtkkTlM23rkEd/Jzt3smfRcu5cm0VnGz06FfREJ7Jrf9CZ9HOJ1cos9rLdRBA9g
u/etazQ2THwsD9DcZZuAkbS5ooP4aqe71H1RzqRbuIZIOy7yCI/LnQfq+U0f2lVcXADhV2JxPeuf
QEwcgJ88PyZK4M2cu9mEWbeocIUxyLs/0iBQxJgCB5MsQ0CGhkj9sg7yCITT4w1Pqtjp3surPdG8
5G6J8QENWsLJFA3hkxAAtYEnJ2tLGHm01rcy5YY/XGf/i3NfQDdNz5sVsbS0RxKMdXtGDum8Yozm
wSvbAu3T8Uy93J0mdXUykc2Rn4UnVi2XBKVgYX1hYXcfBmFDDnzHMfRadVaUnitAu7DQEh1mQCHY
R516l90BRY/AOdFMCvbTUHdOPTxcqr6ZUHFH79qWaJgDoiBNdWN9ziOloiaUSejK59vm3o41wYmI
+T2s7HsXqgJlQF/Pdln4KaazAM57iyfubvOgKvvb2kdfE92ZvcQIeRGinG31/i+k6HypHKpTuK68
3VnGAnyniYAXmyw5VWZWiJ+9o9Uz8g2oAgeMTf0CA5DgDZmCEThUUlnmYFOEDVfSPpCJsmucKk15
NyJl+UPuo8pTFd11dQRXLvF49vEFb2KHU7Foow6lQlyQFE/AcrrIje+mVOsBTcIsZKSKQbej+17h
ltiw3dqTzDVorJRUcpI/0ER3R5blYCgirt6bUzUqROenef7emjRBCO9NRYbshhQ8XBMIQQSz1tgD
s0/EqHf1Cq3yN+6gt9NetjFoaIQz89i2KvjdDJMeAtqvcoUR+Kbd2lFU51wtZUakJiCzzm7JdX6r
q31yD1LGVrYtxBpV8vfjUY7vxepKGnF9e2ZO+pgcLJg+2SoH0stkPRYcGy2IQ4JkNbS0b8Ul1Uwx
rXMj4ufHl6SEf459M549RtvH0pboyOxXlVZoy5JSCwg22D3wuCNQivndDOL7iorlfB9/n4snhJl7
etR6xOngpTcK8b8+HSHb4bJ/kZD63eSejGr7O+QR5IiEfxAQtx6d0doU/EMBO9uCVp3toV8HMR7b
YPojc8fDQa2HRktZTIZFb9Oyd3Qw2KFBoI3FfUGq037OLZxJNN62/BIPLZo0AgTUpu6yavcJ9mIa
jsS7ruAxRMGDq0pdLUEWdj8uGIMeSNHS72QUoOHUjs9oxxH8Guug2wS/ZLeQSrXsd6kVj1mq6/pP
7ojym9GWhoXfEV/1Pi/Rx4sT5nlwU9x6i9b9sfuFcKaLIibdF/33S9eXaWLL4/MW8OjhUMjGRSh3
pbCFojdAJR0lv6Iw8Gg8XTbsc8TPS5ZexMnIKAfGmIILSbB2SIxofdMiyyhoQ+g8CWTm5/EcLYDa
Iwa1YUrfQ+DqmotJu2tVa0gdOVrt2Pbq2Q5CMvCsa7ewz5jq5SBArZqA1K1hNZ9ZeElJ4pBUflZR
HvEvT8VvFUunvdv7YS7VrjJEN5pTSaUNS421DKi8Ql65bJs1NTiMeRy1DM4/Zw2HkBFhDr2UhWNr
d4tF2IyCG47tjAohFgz6LW2/fkzGP07oPgx3dEENeIMqmgGf49cqAbUBYUKBUlKqXv6gDiyE7lBK
xnlGDqfgEnt1y/+Q4NcDmzK/QGWmb2t1kNn4EyD+AOI+Zrcf9zEGT7brXX9ua4SYrHBMQaRCHL+I
Fht5aoostwAUVz1+8rHmwuKNNHgfcNXczxAqP8U8RVXmjdr3i9PWiYUvKWSG2NdHO9qc3zI6KYdE
WQ62hbLIJBdJG5NMrUJOKa/CvMFl3IcS2/0lwSsVMRlqdmEdZz0Dj3ontGUrktqTHb/Dr248bdMp
LFAKilUAS24R/OaXm7WOlDAik8ALJTvM/Fdmv7GgSArPtF4DX5B9KSRegKTbvkBW8E3096DemhgJ
ogT+7rLOU3kJUeJHip31r1btfXqMUVSb+T43U/kcrbEW6CcjSCdHlUDYeF0tyCSMB8vmX4Fq8zLR
mWuJcOwWaIwRg7N7scIysMzP8YZUjvA6mNx2P0L0YvSsJJcZXTRgqEUdA7mq18AOvs/xvf18Js6y
zAwIdgCaprWl+OBU0Eq4XQvzqqKKbFGXyfm9fbUF7Qq1hCrBR1km4VSB6QgqIiVwSs8jcJvbz2yh
GxrHRY8G+rh7g4qhEt4Bkg5DOhJh6eawvt/7bo4cfip3JlrblWtSo1lEuxmfuqaOQICuFzumOJya
6XsVe4YKxSHfRhEbAKf/wZ1cvn0EIc0JwlzWrFQA0ybn7tSCVBniuagzr84rYp6AffY4U+ZRYxys
u3QuDnKb0xkuPzMsUAnQF+sQlUQcfwPOFFoB+cAPTVikWGA4nA4MUcGgY/BIGKdwks4eKL7p8GdY
W6PF0Wl2dDeSROtEtGAgFjDBd/otV/P2+CA3dK1n6R8hP/27bhoGIWdcgLmaOpG5N1GX6/0Sfj31
ir2vLzjOQBmD4lrDL9PNgKxT6nMXz/81IAZc8sspSkJ3xuqM8UvC2UcO5/dfmcpJDTmDPmj04hyT
VqJolj3rk3U+3oDYL96EkxSJ5jv3sJ4mjbMkvmxaHn3NhQumtYgKjMsAcTm+7dFl6nRXUFP+d9Vd
VF9bkWqvmItWUXebba9FeTyuLZvqFmZLeaudffFDRxlGDKUFCoL5tuicLH+S3MJ1FgP2n2XXpqFd
qBO2m4E+S1IuMQV4gbBG8icZJiUYYZrPFq57bvwym9VY4iNHZN3fA/Wa2aSVGhEwOf+HgDVo38ZH
m93qFLP+oY/ke0EiOLU2VVIMRYdmi75LIq4HDo4oEsb0orx148hjtbrs6TixNIKUUVIKb6WLQ9u9
vExPBViXRJBW6jvIhdfKxOnGu/oBxe7wrDOzLrhfLT8QuI1GZCtVCTJ2R5PhvKaQGi6Ot9fy6DC2
XHwIoZQmjU73lRurpHdGSuJTbik5DjsfOTldUXTxivvWiskMz8Ss/ONMI3yJTKsYtUzlaEQXuNHk
AabBVYyEBtu1281X/zTWkcCFyJHrJZ/KwUvIUGPJmqinJi+iQdd7AergVz3tPFo+zPNjlQ7JIwO3
eYDbKXymdinH265WdIeRbX7q6YaouWQFoQ5y2TmFPEbeEz7oSU8XW4cGzRW9ywnk9Ns/SZNgzA1r
bDM8x4khxUA5rbF7RyZKr68FTvxaUSOIAwe3c/a25LunK69m/bjFO6xdYI1O+/lfch7XjeDzEbQ0
GGTO6B4MftuAKQ/QXX/FhFgoILRK1KUdKlZJiprf0mtDVXljx5w8C2GbnVFI58HwviRsYg/nW9DI
lI0kJ0mZAFafiluqTNBq69+Cfn02PJi7aeasBIZ6TvqGSq/yl0pSTvfBm4fCRM+SobAfKCIWbTcj
/aKqO+aFhjm4wUVgv6KQxX4qdGITQrs5hiTvj3CVE69kQYcYIXuL5nS1/ywL/WJwkld7TmCGicxD
zK+e+ScVCnTN/F6Ylp/No7sQ5zCtnnunRm3dBlvMX5DjlMcUet1GHug8CJcdXijFj7X+0TGKZSxC
OuDOnJ0Wc6zk9mkcMXVhv+MnHlc5puEQIMJmGKqjAl90qcHsMKXbKyvYc4iERngQfgZGVaGB48lX
j3jOxgUby6vQ1TxehYnADgk7TsUBiviaG568UNly4Vl3uSmY9UyhVHGUXmrIPM5blusjxD4jTLDb
X4M+4WPS+fnxtRSfKDdPoE2ynpP8jfzztfLh4Ej7MCIOYe9+YIFYvuT3Hw9rweaLqpn+bKb2t0xn
DCMx5Qns76x0EiH3Lbd+RfIf7pB6uvsPbwB3iqSaCxVZplBG7Xp6JL9f+siK2Pc9MF3QHgBWQnt8
FVOBpSx8m3iP2gH+F8duRXmHR0ibQZ8zy6c/fAwffzQEjZ8+Wza7LBHp/lmFJ4L9lO+hEshY6rBa
RoSwRQwG179ccV8ZgD/zFkXV0O//WQvn7uVmCUgg75ac4pfD8N13+b6zHwduAE/TADBRFLMKfOVw
HtZfEBLf/uAzk8jDkviKJx37d4fbO4u+ifY9TxmG1k/ueKW6JLTy2DvZCcyQ9X99thsQu02yLjz0
YS9NqJoyeroISHyE6wPZVcqlxQXWREieF6/afNMPk8j7tsvnZtR42AFkBuw2zBi8Q131ZUn9XFpl
GWppxHO5JqlmuYgw9XeaTrkP6Wn/tG4T5YhxDl2L+GKRkpRhqXflPs4S8woz16LLmumv3oGDWpzW
rqEQ5Y8McYp8b4xSdL87GCzNCzMjGvIbFnFGu0OCBh7I6csFiDvwpyDVQshRMg/Qs4V+GVFoVSC1
Hc3NBhR7HFXGX5vd9lMC/hk34DHg5kKwApL4JqdITANGtDhmqv/LVbK5iPkhnPQeGLVo23XjYS+H
utu5AiJDY9rzSgc/PXPN161sJ+7vy8KtRv4/G1okBQWftLBSo8cy4ypT9v+LSjrmARzUTeSxh+Qr
C5J43mBQwOSZ3dhYWrWMkZC1+/TrmdjiWQQKNtvZYQvTK6YFscE8qxx5N2qBGCDGvcPGZ72DzFlc
z/l5hS7UtgyFFxX6k2LdDCnD0lPJSlo1ydDoZ+HCZAplkyURLbZe2zasZd2VwZjqFnw+xHIQ0roI
64Ba9quyef3gDlXMH7/AJMU70BWUtKsSUkcgps4IYSKT0swynqfVqfeLHqSLNw5TtsRnxpgI0FRo
FPtKpjJsu/ReRyqmz/r9w42evNgqmANqXUnue95HNaEBUgJrRIDFVv8Q4SyIQKlAAqY2gJZtBUvM
RmNz56VTdW3ORcnaDO+bIU5pTXToaNvidK5RNMlPNeM00X+ZCmqlt0sIuLTOFVB268sHU4UXwgKt
eqLZA8nYs2w5BdTr+ZlIH5EcbkimY5f9kjqxClPfxz95yPsrT0HLj8UW3MpBuY/uwEmRbu5aI2TJ
N0BzVGeORoaYD2YkXx2SZdYVSSbMYAhAhWyvNZnVUAQ/4BuRzZD2bJhvyg8AXQSFw9brx0xPY5aR
YFo26uC8QJ8ChN90MZRZ8Htnb91hleijVbDyAq7QyHeqR5MvclGWwwn3AiwAp/71I/YRqpG8Q6Df
CCLTr99/6raABMlQn2wHlpdnJY3uagjyzdVSFobcDuPoLs/j8K3GVSu2nETdT7DwW8k9xLaP+LOn
Kv3TP4z7lev+iOKhEEuGk44Hyg9czrerAp/JVKL8YZ2AE1OZL1bhCcNoYAFqt2uIFks3m6MGFOVl
3vBD7gsoPnOzL7ab/tXdaslnJaLYLaC3F1w+7sAimHShh12N7NK4lKLPxFwclskWKZ4k+ta6kwtp
NX7tgCXDXiYULp1x51fK+YwiBvz8T/mY2IAkpE+21jQcdJ/kYY/W5irrqRQrp461aEJDsFVTPDvP
n4C5ONopJUQXqhaJCeDpW5IDoFBI+VrzXI73eK5VRdg9DemA1O+TfKWkkwvypodJTIj5Gxuy0dLk
PHVtTWakIgrgLk97nXt7kUuc6YCcjCTUeCe92jQF0MZRySyDBRXVdFC9ApJcuYjxUmkc2I+/h0iK
V+dm0VyJqHuntJhz6aHeWvc6lhdZB7oTfVcObZsAFEKnz+qsAS3qmc8ElvtC4JtuXQc0MRtlkAq5
e+fw7+RWyu2LgHbu9KhLOsq8eLBPlHMJt15R5ibUh3EUfAhYoXWW1aHjN8G1rfa9/m57IdutPc2w
iC0mWEw69tB4ezIajoGKbWQxtg5k6vvDhkYpnuYn1zpqE13fi5kXruj+LjXT43+Sni+7IXtmQIxw
aV9jhAwykiiM3tTbGC0QXGdkGjTmpb1oQsXWYI9sJIBgGhXd7E/bsLVR5yVk9Slla/KbePIhyHRJ
WmtchWFspxnDWZ1J9gf0CkkFwSFB9WyfehL64x/Y212ZKV7bjzYFa9V33z173zm66p4GeEUWuT+1
UkXfxsmS+Qeou022bCBTBskhycepMLy1YwgSxJAxqZnheJ+y5mjdiKOteIhSNFoYxRJj+P6ZKUK8
cjnvk/HUx9rBkldmHRgB9ctJf4a2B2ifZQ92V6F2zJsRyVse9KNIxYjNZUqrw6Bs844vD2DHpMvJ
lKYiBZM1yr4B0YNAh8SN5y0Z27SmNboRcRszv8/A945JzBMTaHy9YjFd/Klwan0Rw2z36z7aSWKf
iw0LABlXAjInKXt/BBQ1pNEwWNWg7SoxIttaSIE6QKHySwHj+7hh9YwjwYezv23Xo0YJcmBS6qFM
aqB3WUf9b4FtMkhDXYORGedD99Fe/AEKU4vRqU5AFKOh50Pz+Dh6IN9A3sIGovyN2L5HSK3LucC2
MilR7GLV0q8QsbzHafUX+ceKZyhtqxp60tr1VWl563nokyNXbw1bNW2UM2/48c37mLFFsLSz0MjU
3YrfML+K55ZXukLJB0IQ5XupRArcwkzqzTsGi3cbFLWj3I8gH6XHH5IuEr5+6UjEPV4EOFd/Ldw/
0Vg6nDQyJccjITBpY6OGnR/CnzXaq5pqaupbCSynDXvJT27Od/001HJVdboysHgnOQmSieKn4B9G
PEF9VQiwIUBI2gV0oLKD6jhlyV1cr95Jy/XgWFuNpalsJEgs0zKh0DocGSIiL4e/xxpbojsvXX9M
N+YQQX9wbQLB8Cx84fZ+Yusr6eEtPDPbgy3bbQ6Ew+YqmKixgrQxbFCadeSbqL49MKIb3wYUGEnu
2dSdrIKEq8oMf1DuPFELa3wmJJrk0JuQ2COElSt2isJM33jvRc441nJn6ffBLGwi0zH1VlSV3Qhd
vKd+I4JUgEM1tTCrJ53lJQ7+GaZZtyBtXaHiERt2yhfBISCE009E2iTn2ArhFQTaTlJB7ThdblXW
Pa9MoEUBql1IbWkhuJWspjosNZff9esrv0hWI6y0TnqRmc9pxiFkkXU4itRsGEktQ2O3YmNaxFBa
pYC5/wrtDNPwrTlPCIWxtgmBWiQ8GSt3mgvKlVo9GSC7J+Jqc9vMSRJVkmVW2z8hNARNkbQpBTct
Pru7rKHGxWzgdDQSt/nv5Z2E/uCVTh79bs4LWaB12hx80L1P81sZLmfxzqVi6k622uw0fFsU0rCW
K8wr9R1DdG6mVa6OsTwBbS35Vj6RBts3mSQ4shUPJhjBS4Q9orJ14R2bEam5WTXeG+bQuF+Et31A
o0tQByjuPYalVHDjsJg756Ox/rR4McyyJwys5Z925RTXNis+mEBtd2RaYO+octgloJDDd9IauCt7
GuNaDngpwifReCQK4FGF6VcVTbLDdSOE1HAfhR9giiUynk4bLqOpcu89J5uL4XakuR11v8150EWW
tYUTnO5sgYRuDRwdN/zUB71fS9EKtxVWL4wgB/WNtagV2Z7sfs9trvaDB/lZQJ6jcihUo4rYU+nO
6arOPSw/cGWCim9DhMPlu5AnzpbQMZQMy1/g2mG3V0DFolXLrUNeYPrRWkgxJu9b7m3cxYjNbV6n
z0FCB7gZ15lZNyLLuvbI6JV3yVapi1ii62+alPY+YI6nLjsLtmMwVQE+RjUgeyt4koH0voZznYRE
CdhVX76kkBzm9hDt93fzgSIT5uQGREKw+bPgkf382wo/4pm572bMzkfk67W8Huvn4yGEUPOVtTN3
bh3/No00Jt25rp7avOvwbD67gWgXoj8wLbVaHxRx9OH4CP3jrc0VMoHh/FxwEPsQQAkznR+ga4h0
WsxzKEY85wsgvzU4Debbz3TqxqUbs9H2bTtlnjCRHj5L+O5rTYHy9IaukXC8dnsbJjWPwYlY5C+V
o8otG01HJodFVC0NS4h/lJRUEwFGbeJSbK8dv1GjM1kyste/BFuHFp+8o3Oi82fJc019UlS4BLlY
iWUKRTnLE0P2EifL9hi8ePS29QfexRlXC53eJxcQCmocNNJRm55jXgl+Nidl1ZPFAKoyQUd+IKi9
PZ+FIzBBy4Cjc7xb5HOHiVKRDgcrYKbvqhDBrtUo2CkEnMQilg2Jjo4rvzVr9lbPA52Oz4jDTNVx
V9hQi0vJq9FT/HsdLYXYOFhly4E1ohUbmdy9MCGP2AlyAbsfxFzodbMqYVvMi+bJyVUoxQUayc56
ZraWMMhUIfujV0X5M/nhccjCuNm2OCyx7x5QgctO66ORgog69CpXQO0Whx74W+iAqtojkHvkLnEL
lcwkAtQRvx3HtGsxdepwgnvoKevTNh543kS1bF9zrxzz84pBLeoBwSeP1cvlPgBK6Jr4mrRFN7Ao
PpwTp/UVK9rYkwHy8xkrnTU3rPwMKilm6tZi6NJvWv+vZbQGdEJUY2Ulr7q+OnX2Cs50aKcVyuP5
moTpy69yh6cxVi7YK4runHp9DPndIJfyFJ1gEEFEg6ngOJ62u+5bwX1X30FHcIBcIJ5PcIjFu7N8
Y1otmY0MGJTE1RV+CHyrTdsB0q4bxMkEpmi1X0wz7ATbZGoUcME6bb2F4xhP+aB5ts7KNiXLqxrU
ywOgCBl2LiMbenmGHqROM0IRLehK00PK/wiK1DKqwYlZLAX/tNUJA9QvFJLe6r1ypaCVGYbKB2iH
+6W7P9nL0IcGm+YttXMM46AWLltgye2HFmFGFpm0syieBHjs7CfKRsW+mLgr254M5DuMrww74EpE
7VxeOSokgG/dJdTaQF2HYh4vzQLrEVrdtK4NeRF1zp6N3LDzN+vvLdVxXaaa+WG3EoK6ZpF+07l4
KlH9UHiaLZZPozcwKr9HBYFwT5bjwOiuxbDBu+5TSbegvILb2Li/AjInQoKvdatSPeKlmszfwsMa
Rgd3DvPUnr/UJCqwrV9pOMIAw4yqnc5iZQqLCGCW/jylVY372fFAZeRO6tiQe2r20o3REJyfL69W
RvsKSoWXAmC4/Oigtxdz672uz22+TMQ6szT6UAcjOT5qDyBpAu+FMcUMl2nT6NwYJd8uGhvo4qjJ
FD5JXYQntOTa2zsWdt49ozkMoDLDiBrIs0LhWWMYJETY6NtjjDLIiNTMVrQrgIc2YB2meCWY12et
zsJ7GqobdgSOo0929bznCdtJtTahasf/b3qAGvZfEpkNZ7Q7NjF2sbZWME1DKt36czB6nRwrGU4x
V+7T5TBzZRWEffwAJZZ0lbCUz1COghBMcXuSg4lnbqa/ekeiDg1pI0c+mOm8XI8WqBLIOrkURnxC
tPYCh56viUUVI3KPmvHP/cm4wJR0Npdxt+hh8Tvph6Dbk3j1cloMJ4I5m8RXZmV50ln6K+l2iJ91
k3G6fQu0J2e89i44RWVtW4ErixUIJ9my/pnzf/68GT8LbP0h8TSKhAJVCqWl1JyOVSXiuzl/HqAK
hAH1LI4Stw/fXJYQgCCEvnBadWfRbVAwNbqXVl7r5EeNVVICBurOveenCLsOMQK5C2zLuiZgrXok
CKOB4U+y4nISFgIjB9dTGQsCHQ22y6W2rh3e1SL4bMn1qOPrSfGKl8+h9gm76isDy5Y8cmB8z1AI
nc9/v8sSA/XLLpG5bHN7Ez2pJHeYOmI89Nvoclh5NLFLYUk3RU0f7O/ENW+SNpKl4u7wNhlYBX0F
iwRZ9FZLlj5b8/G0t5b4+ERibGnLbT1Yp72mrCYCepJFC1cbQT3a4FdQZpCv688Pu2FLIAEe9hV7
B1gFts2q/JQaA8E2P9vhkqVuhnwxp7j7uT/IZmmNObfljL+cb7mdhQM/LwX625QjEkEXjvi6Wu44
fRHwPQ5kYgXJNpWmTIaBemDVGUgJuRB59pATZtCxcmmuneoWDe1Ixi6jOiQPxqMraKqc3fqi41oI
P5dKwQk+TH9sbCU6UiK/ZTJnmGA7YtRZeB+N+Lutyd9SeaetPqgnhjjRg1vMN/MkR+OHrO9M7cWp
30AmCFB/w+uhNa1Y4R18erIyF+adUMxPJyIqgCpzDCApxRcvLKu5iep69EVLKZIdHDSESUAHKKaR
hTFNaxVemyZB81YRAJ8Pedv5IZgBSjT18vOJry0A6JKAYmNw96dEFsoNIQIttSelfgF2R8bGj1i0
IdX9kO9nhKNmHujKTdEbz9w7FkyB2xdTyPox9EsycG6IZb6fah4gFuWQbEFXNKLtUIgIwQyJnc23
5y5ZdxrZBZq3tMtWprll7fTWEEcZVF6vGN1K4aEJoDVGwmjYe2a9kuyJSPUkn6VcoCC+4b/XJcGC
RTRhARPwibImS0p/Se3J46ZxUZDflj77A/UaZnWGSkxDonUs8dkuhlhc89J0lA++YQ9sbGmBVDa3
OVA/Yh+Mk0b2SmOhr9HD6HwWvEmxgdQkfQcVnhhK//jDGZ3/89HDnAxoR2rTVe+KGc9eJ/BKmcJs
shoFIKpSJPNiL10ma3tkqKkMSFeQqMCwFbM9ZJhq68wHqSpx43R8bhjJTZyuse4+Yao7Zyo6VwkY
OMPh4x+f0euGtC8vMGqTHnz6qVzktO5ypMxnlEg3d6A9Ma+U1FAwQ00ZWsqVAJix8NuZWw1VTJgB
xKKtSwrJKsQV6sUHgJlb57AZJqbPaygWLBloh7jOPQ5TXLdlrZ/I5+wcTpFnLngzcRI7WF6QE2hR
ua4ag+HGyoDiyTskoCKX4iSVvVlCIH5Fci1n8C7uIWHbadTwD1Uf8hDjxvKo6kTyqArKCiuDKGwU
IXPffwXc7z0adf9XLNG4aMnoZdjkqW+G0aEXjF8kNfiHKoy+znu4apKc92BOTcVVJuUoLluPP/VU
QPbzhvzOcAQDx5ee5YHqajuFxzBbQTDTjAwWD75kaCgpwo1oDcfzzpO10HsRRzcZu6gX8CEYT57a
qjV+XyL05djc/X/o0fscNA3YWitE28Xdv1Gcezxx4X/dBnVDAAT30QZJQKYyXWrZafA9tlwaCfEO
YTYoWtRCxlPRfZaTRH873RMjx86BUP2cM9oIxAzby1XE8v/XVBRHF2jVZvv+qdNnqv6xNQo0rBTp
C9wdXipS9EunIvuoNovc8L6YBxwuVasSOGBOZdCjRiemmIC8Irc3lVQAYlP6vLkU/MKmzxgr9Y4W
Oo6mLofAM1Bc8M+HzsaAyc6xU3eEiuW3E13Lq1Ffv6Wpt4m+uSgL3313e0wUuaxxzJDx12ckC67y
5FKV4Z4HZftdIQeSSnio/nEKJqoNzaDWFUmePLptFD0CaDP5iIuneutRpavisO2fm1vxZ7/7sy5s
zNiZZcH9nHYzmjEZlpwDAW1lU7zJARpnbBFIes8RLLl7/baDUl3u/XfIF0SVOFz8Q3JMsnc7UTQ4
lA4xoL3wh3b13JwO0qpE30iNNsYPM8QO/gNfel1YtF4MZG4FUj2rt95fPeDoWArqfvMhWL5DUyNM
2GTYmTGh8yhIkGOjFd8/wTbPiLQdCvYZd3j6shClAjT3RhcLVIMpe+xpv378Nr3iEYiKCCjhm3Dx
71AKjjY/qeGIXZQ7u1dxLNvLufi4Hu+xPhyVTX1J2/heZEJvJATb68UlQheHLTZfVLxPZ4Gp+xv/
46P2ynE6RmHhnsBFfzeIogaO8Y64m/zozk93pI4zl8NAcU6KHwp+G+Td3CsMnCXJPTYF2N0HqcyH
pzMKgI6FQwOsi88+qljMzswyTGDR+7t4RWzXm5NDIRQm38i2zhdh4NafwMKuMCFISK0J9sqdMxXv
X5pDwNvyUZbiZMPPfGAV8rL5HvkFaU2DUZoOCUU7cACIolZ3LBznoj2iYmNl8x1gYcwtCjHCn/4A
lo/yDd2RJOsbYLGHUu5ZLs3lQRIE10OYJP/mVMhakJNdeB+x6kTS0ocY6GdCN7R9yLTimJviWLLK
W6BaUI1kf/H5BgeIkih/ul1qynOEj8UmOwqqxPwQ91g4GRZvArcXSwAoUEwAitBSTsyT/S3kGylw
QqygOhjIjKOiK7mYzPYQAHlHL5zya8lV9soJJopUoydDZ+8G6Q9VCyoP18wcbeMWBLBWXax+XRJ4
8TgIP7CcAqCyzIsWwh+eNHfQ9x6p8lZsHTDZHC9D3x/xvkACXeLdx39nzz9WWDUfchAO4r9LMh6a
AWCZILomUd5vwN6Gk/1xZnBkh8WiaSbAbNwDdgMxO334TkyOfQd6l6CAjMjGjZGC+CDk3ajHSiO0
GTGArZCAE/dDn9iEjVW0G5hOAuAV0cc0iNYEOFpqx4HQEEjUF+e2O5/kXESjrlGGJas+gVbiaNsV
+e9LjS56akw34P7LCg0suSuim7DfYMMnksOqxffd8ul0ImMQl0bIbikqZbPHjapxYPXmnKHlfHX7
NwlqdvWHtbSth2NqC46TYVnZschD8bJ+m8d652wJAaDJH2Ciw2g8KyMcbu3vPTR0y+gtkCI78b21
72rZyOFTWgR/PGqi3+YqYtAQyOPgxO1ARdgodcnx5OWVaw/rBSoGbrHdn6UIfDofl/KiD4AiZrLt
BLzZEgtZpV/MFsVNjtTvA8rqHv1XJNCJabRDrkaJLg4na0JUKSbCCkQDQrNxnVb/fQOnJDti5NtO
oZQ/y/cooRgTJnEDTy5iuurljLWqtci59Noaaz+LVWs6THo0PWcsZkFPtjJCWGD0hedu20Cd+LHl
3QlS/GzE193QrpxuIZAGgdne9HcTfaKyfKIVy4Ufg1TeiSB6DsNGLCjsH8wl7qpyNquSJSa1Blho
tBYf/X/x5Fdh2tQ7FzU+9AKYbgkPt0nWMva6S5sAR12gOI81c/l/ll31NKAe9bazpNNa9400K044
bKRjXjsBkKEL/f2E80K6pYDMv8HvesctDzEEvzSs67q/ydb2yHqvO//wb00Q++f0em5zJ4tV+OYL
/QR2GS9Dq2AyTN5drS8E4FZLfVJmxftu+p/kJQuRMhQRpaY9ZsjiemteXN7Au7kAlQBscRbdJYcU
k1LkyQNG0w95cswOWpLkMf7ZgCSf4J6MqLdh+ASJt5NarJitX+Q8VJA62aUWu87ClXyEKF1dH/Is
Jxvn0vysi6aZKsgJuJO2ZhrGs1zQqJt5935I0+18ChRdTgMvkjsREgAYDo4AKfSiBwe1isqJ6Dnc
DnRDQnz4hkOk4f9T6NHXq5/BU1ZOn2y/LYUTo+FwhZJZceyxVdzyT1Ylp6MIoXfQFMqk+kTkbvxY
W+AZPGMkgiWdDz3YjjVVhZdJlonWAPANn5G5WflE6+NU7O97UMS3l41ivtw2ZMWbf5eEy1vH3xV/
LxWHK02E7FdkPDMBAVKvJnmFwCx8SXkGySs5JIpLja/fGSGZPJZ+FTWpEce6u/r8yS5cov/Z0rra
ea5Xsq553T+8A5iIr1fuutt/c/Ny8J5aBt1YaE1HEfFIGCMDKt76//O32bE2ZpmQ6lZuqgWf0B6c
WK/JHm+z/XdsiGnTJcuU3DIb5WtYxnifNmShmTYyFFMD7XoWvyh0BOh1aM0AAW9iIO63h9wtj6xn
FN8Jse7oqIQfpr6/DKBMaWBeB5Vs2LftnABMwtexAfSp/Ou4emOOsKYHHAZ3A1R+L+a4jGKV6dA5
PmHHc9f7y9p5OeewBAChdGul15LHYcwKtjaEdEOYVhkIioo7j8T2RneBGIk+Nz89CuD/zK43qKBA
Xk2VG2AuKwX5rDinDoK0gn9w6hb37i/cJTd7rKnJ9VqmUVAX4G8AuZMcAx37Jks0SZxv7eJnXvBL
tlLFb5DVqziveXLigSOS6h2tr71FhYxEoLEnD+B0Q53U2L1V0atETYB8imqov+lsKzQWT0Ia7LQr
zl6PYFrTfHdQ2m+njvadU5XRs11gs9JpjXrBmhQBXDYDHThjjfAGNbLelFcWlXFzzEHk0ldodCYK
w4CX6DVANA6OcomA7GwXqphn7p/0KlkLgIyuVWASiXWCeMJi5dB/yaTXyh30rlULOL+JsBK6KzPy
TRGsEH/1tEA6MNbMzV8SbfBWwVrPXIYB2mjEyjGY4KPYAq0yaeHbRQ7rkTi2f6YTvtER2JoS+zo/
BC/LS9RIZKgRyQww/0e/jTu4vKoXU/GuyXEDnYqPNgvfkxzrBBSskzILjMRiMM0frJKnERHZuA0o
GkPKhRIXWoiTOOBcSJQZ/OmJGTEDZ4Yrh3YET2D78OAzC6jGZSDl1SerpOd2CEsm7ynnq9v4hp9T
9KtqdqdQp94pP0mOJcoAIlqjURIhSYg61kl7ABzVFGumP8LiROQ0v+hBH2LjccLPVoEA1G1rIwmv
/SD1amROde421UNOZUNH+K56WYaydTe3WcKVdyi8/2NroMd+kmBP08E/AjX/suuuq8ey5h4xQEAj
6uPmCL93wocx16oGb62pezAd0qaheFaeA/gHiQ8ILwjgG4Sx62WPa6bLgEQ0c4YmennHexEwYFmX
0faVby5xXjlEMfNSngTZvpHwK9ka+PF17wczREwWC6+Awq2pfYMleHEGKp1Hh11/zGKNsprGqGK8
dKnrETBVIlPYz33wk4ZfCa0lO2OmPS4MgIYA8cK9tDkv3gAHlrAWcqkXN6hhH0PgrhiPsbG+SUmS
bDyRlv1ynafw7RBgzlaIaxI4ZvfuztkbOwujh+pgx+bY+OGM5DckaQ2QlsIcAir8NcDUWRK9h3Vy
NvpeiReRzRtS/ZDpFL0ykmKA4tILI2ckl2jBQll0IbktgL/YGm/+6ufcBqc3wvoohWHx70YdAS3M
Rv+HMzQgZPKTA2VlYfYBaAfMqDtUTjEwhSCHK2c28svWWvn2Yxw3qhwDjHrETWnaZkVFKanFgN4W
8tlcRt6Wu4mwX9Jg9VqQVpbar1J9eRFNMHJ/6h/CBEMEYJBKMCKMEZy2VFpOVfx8blYczxhiLfIT
zWStcWHbQ6DtrrAQyNP2z6YlyM71YVvUGXsdnBYiN3pVG/8yNHUV4w9isLQbzb8uJSHsMq5pO9PR
nhePCQqEHt1IZBsjhrBVV+2G530jVL/Et6pUsTO9MUKW/T0TTF2E2rydSKu74dVdBqLqtx+PQcuo
kUz3V3PD8wlb7SuCMPzODbj7b4B4R6utjBczsQOK+JGZj7ez5aenTlp4hsN2rQNbJpNvNjVkLOjk
yh5hzbljMGuAXTtU67ZL9yZG0Twt57Gk54UjcW13/PYSvRhAUflIDRShtLMEV7plstQcJei/n/gK
5CKvnPwJopXF8MeyG0zWb4wPdA+G6jPhpyOiM9ZLql3P+rWrjDTSXTCLAzm1uYk4WFGD8XEsqTyk
LqzpM2wnyWViIdMIIYMmZa+R7KHF2VxwoGiGVnsSS6nngeQun0pEbNzzzNWELC2QdHb/fgz2p969
Z1YQivNsyLK5ShUi/5jJaZIxLkjoqCs3oTm4S04KDzUSQcvOCDguH4ELnSOB7sYmo1UIg50Ff79e
nbWlFYlx6TfK9xDeJEaGfLoF4u9u8hIr/OxZZ8JMlhCcFG3UrzbQBdTQxX06BMozJy3gpbKpntYK
2uTTVdoIgEUZnT9LCbgF/kPnJ1Cx00FznjmS+QtC4z0Cs0Qz2dEwj+pJkjL9DCdz1RRe3tqMANz7
rKMzsJZciOTJ3Iqr3+akHTcVOkbOuf28PfmcwPRfSgRyJcfBilOjffcYCsRBQzjw8INdj7zb1Z8D
klqkBqrqCdctBu/VpjOjxYg+M0xyw98FXqJHEShE1JfCYm+NASeli4UNbF85NnK/RWxLNAFyEjI+
QRwE2ZFJmirJy6DxXuNuxkzGmz3H55rOTxPgQ3Z673y0cyy5SGKloUl16rki3Gn10x/6gVPor1Yn
AsQFUx85BhCiEnZwE/tCsY2WxYSzgftL/Tc56iMMuxSQE7T/ToNMOa71cqn3W1fg3j+MAi4LRy71
ru39KAVMVKQf0OD/lxovggqUb0WJ3sWtrMzfv3MMfNDCFi+3HMxSDMNJdzQ419uvKVTBjIHmTt/u
usmhFYAhaIs21V5U6C4upyHeJJwD3WismGmyq2gWIw3XsRt76T7iB3D5/LStAYr6BL4HfVyETIUP
/+Hl7K/QKfN+gE0uXnQXrHWhsXnsIMV2w8TAn54iVe7gDdfE+xWCw5ajN3LEMV0QLQ86DCBgV0ps
EjFmn5OIwES+hbF4nloxU+Cg8kp+sSdGi47xRf+WEAAohyKp8IOEZjsVPiZmCpMy81Izl+zQUEjm
sekhZDbBG1bVeXZh6YT4VFXu5BuzCaJ3mQ/QYK01zVCJ3mNh7/ust+AYKjH1xPLAXAruRFMRCeq5
erqgY5VZc3uCk/W/vmZQcQf9xH4Sfe5turPM0MY6NkH12+qAAehc4wDFOfK/+XZnQ7jAlxX1QyTK
qB++YEX4XfaCObtE3x9eF9AuQ9K0iER83hGGA3Dn1pBWFGHU2Ilgq4jWA6+hp60+kaGce9t+Dqmi
pssuIPIs/xclf6NU4gspry54ujsFH+KFX5kemI0YW+tr9JnoMzv+U8lPVd4y4xOvkDf6sGSC1tQF
atFFvoM6Pe3eh7yiE65qxMiPt9A7VgdyES4fgTqdPYussXZGKPHahCicoN+XPVZ7iPMnZVN8qyr+
jojaxttp1LpO5H/gvUpMdHkY9e0D1x1Rw92XRwwTozDnhKv0E9DZQjRwiwL71sAmMvbWORSDDSq5
R8aXbky6pGc0ZboRJ8qa6T4aoE2xiRAmOLNTgvUj5JDzy/hfkfhczAuhi79prV2epp+vKKlR7NZb
h6NrarfHwlVDR28FiERtXUrl80pIvGqP8yvgUv+0dNm7YvJVXJGo+qRZJCDfPTu5r7es3JcQ//B5
GxM84fsdcITKhPn5754+vKuz89GXH/8bs/sgtPzbFHjwvSZwo/4mtkFv35+g7iO5PrVL+dOyNEik
r6EMeYQw2WnxOn/IJwcxTy2IE9C1/xq+9UJrtdBslra1HXRzw/l7Qu/wk5pSUYIt6vbd1wgn/EaU
Yic+awt5+bozpfEuvb05XjPNWKK7qbmTeQhJtMdQIhzo64GiCU2wtsmdqzsuR306ve0BUuGR5G4v
+EjB6z3Jm4cxMCjdIWeS0VbkpxYOndzZR9+vbDFXkUlLh+7h8FC3HqpQvvGIRBwK5qJB6gvHIDQ6
0K9rCHooW0xWysrJ303XTZ7jaiqITLBECdwt5N387EMaKo3Nli9FNgOufNDLoByeWgNKy94nP/w3
j2Z7LlUosPqp6G/roR0R4MJ3mocG/6qspfolqELbwQUU6PbqVZMsKJ+fET19qaVXRq9T68eTExnP
D2PmUysfsWYgBAn5/eyQNtjvxSta3Tmz5Q84V5pE3ETxyNHagjszyH7hNK5qCroe0Blm8GWtevpD
8TDLguz+ZdQXEDBCtAhDdYFtJnMFyJ58deC8jRwaGNNETKJAqbVIFLOey2hp+Y2OMjH1X8p4YsKA
qa52guDgmuYG2MDRRTI6Sbw35ZyxlptA5weeH/00cha4s7ALujvDnbLV+7mf9cHx4uLL8eZOmMf/
IYlSBPV8DldOEy/Ko7Hk2EGeJSY8cEGUeVFUTGIHw62oqD4/BO92Y0OfVfouOJPA4MgZJdVdtaIf
kJhIrqU0pdU+VhRba9LClA4NvW8PnCQWTaRoYNMj+TeFFqlGLQs182ugtFWKBjbDq5glgBv6jg8i
B6ssZnygD1n10GQbdbzpd92sCuKWTI15fsReRDqmo+TWgzwHrsfsNncGiTTv588ct1+nJ+D19Gz0
ugNygzfP+/D3m0kww+49KWq0N5cW/8uFIeQCR67xkYs2mu276HWCjPwtzQMyzCiIcd5+s6xurAwn
zS1seUzdNPSEvm8Y56XVAgBKoKDO0X2xreLGt54o2viOhy1FdXlSkBGuYTnUcnQ8DlGLowktdZFB
7lYFsxkG2qa8s+uOMbH98coWpRfJpbGjc2SEasgxFAQyz4kxI8BnJFjs52OEO5pPQPMJtp+OujKb
uIg8g3XhRaAcxvE9v7Kc9bRo6txxZsaWPpXAx0Bz70WwiphHE4DaXtmonktsDNKgLONW/wlqPLpa
emyCIKFCeNh9LTBy48el6BR8Z3tnAjllQBDUzWZLIhs+MFoe7sMwspOwmjrHPhygZs2913eatfwm
arlrq7XKrds3616iRmAIKrc5HoBtO6ajfnx1zLbP+kAvvNwsa17b3B/7dp06BL5WZXKLEJVpAdRU
pOWvO0FyUsnQ74ielFq9XbtJ/NFv6C/sF/gsbXI/a3zpaauj9THe9FlszQgnkBjo9CblEHX4w289
bGcbV+oJdIwynlf5HAHXzcC2LAJc+RmJFDpzOVIQOoBDE2KeHchRhU4lTvTASdTBV1i6R4ecGdDh
U3xhalXCsPb4EJtJNinsKUJrPa5DF+wEr+ZdpvtILp8JojJk93b1pNPDTTkyH5eYLQDlLjrNx495
fLY/uiManH9urH5/a/I3pYJpI3xfwdRQ9BEkAzLwc27CxPd/8fU0mbL2E1EnIJPfofUu7gXkRSXA
34+J1P8wtCYySFEPEmu4F6rVgyo/eebYGC/e25FobTNtZRbZTXEZHFVyLOCgOvDrHk0ys12Bo0yA
5xBsAllQyL5lqFZuyoj9xzfvMsJXC+5HI/aBHNLxteEGrTFQMEaMADRZO7e1Bzg6Bc0Q7vH8/muu
pFRNMvy4gRq9f4aJzf2oMnDZ0ynX4p9FdVEDn8/AwFm4aikptrclgAl2I1bxetFe9vNhxJh10Soo
ThA1POE/ABFCyBAQFF+GWiwsTynfVleIsTgWWzaZuSfW4OlOlZ2rPXtmi5Iwt5D1HS3iLYgHgZLR
9MvOL4fTsdoyBlqD6FTMv/yz7xOb3CtdgwB3313rzbWjh/4QOyK+O41kXkJPi+h3wH/ipvHtx9HN
vhH3U/cSKyqX4j1Z27/ZPG9OAY+HgyCiqPV7NaUSksrXwzLz/rm3sg8FOMxuvLn3Siu39u8FFLIB
antO+/sVPrm6KzZiU71rvicmJz4uRn7XlAnBCXWbJItb2v1lx7EPPTqpLkXsJHgR8qFICd0x1xAM
G3O30vr7MGsfwxuyPfwpv8W7cg5w97EVc2U9HdgGn+HQ5OUTZKlIE9EMeb2lmEG2Mr457fmtsaEu
H9cJC+7cdw9ipD5CJkRXCdHPxpGJAZOpAefh/YMG45hvY8yFaaMN9je/urvJ0drYLRNI/16qHHWZ
UwEj0ZXdShn6bWqBW8nEIWEQ7ocVIZMxNBo5CB/SfBZIV9b44LGnkcPY5/C1Q2Zmx0MEpEApEWeG
PnWhIhQ2ATo+WGqgE1MIycf4RHa+K1raAds3BXI+AH2V6aHTbxPA3Zycw6TDJXRYeuv10phBRNih
9VSkN7jlRg7fEjxdWvP/ahrVfzjyEPIyJtrm/9u28UagvNQ1x3nmG7TdjnXvcOFR4nycqharREjP
HXGGewammBpec+FgFvHnqSUOoSh1mSSZdGLq18yifq5uGWMXx/ooBbKfUn6A/n8vQUJBWyCAqpLY
cq5XdbGlCOpqo/HHUyOL7Uhjb+qPzpcJNn+zTjQj0Of/NLZO92cGwGHW3hJy+7fK+yFehz1N4VOf
w+j1oVpHijbSTENMPBC+wAiymiy0WtIOpsLb/bODptpa128exrGpGv9hvtRSz/6kfmoAhWXif193
eq34KjwXgzu9+uk2vp5qtFAgZFmx7EKvRkYA5SGmshmWMeWTh/NckAiNim1kKwiwbrq1JaNAIwmp
kTNI/Ypd3InYTxE4pu95PLGxzmhdJ+JsvKH489L0Rh4/QRtOJ8s2MoU7l5PdDpcaLUSH3bOfIg34
7NF2ONudqtVbP3hsCdVzuOyOdCaLjwGceffnU66JAZxYvWesTfrTXGBKS7OLAyfeQfrw/hg6PNPT
T358VLd+xiPJtcCqKbhJnUOUHzHCIxFzo2SxAxh3g2q1M2xxGZtEF2Cv6LAlbhRZ2+u2LgsXig0N
8v+G5/eX6QS5mWaf9wxdIMgCUcwSUE3hcaVF7vsZhAd5Mh0+1aE+K3nJlGaTo1d4veHg4Zxt6Pr3
Fawqe1nSI0vDfl549V2ptaJvum+CW1ABUh3oyNHByFglB06SXfmxU7tN0yZ+t25XTeYsSel0fan3
274+CxCMg2t3qpuSYJXL1TEiH1XKhvr2vkvf/cHu8lzxtOd1nasjRHSfWwg5FM38L5EU7mtDRPgG
q8ZqnYpWYinYFOaod4rPk3F61WiqQXlx60KWLnMt4vseb0vS5NavPC/aEyDuAYjxQe3SOk7yg879
Wj3OINv+y261Xy1Nt3ymzb1mT+hajzPcOgYHWS3qr4PwvvytrkRnFQf8qP57po7LeTetAsZFcgyL
HSzAsUp/+QZSPYK6bK5lzdFCACcynj6zEn0kKVzMpkCG1cXa06yc3uvposN0QdHmVNsbslOSJBVu
srRoTn0X+YoYozwTYJNH+gTPJ3JpI5xjCNMk/OgNjwQo+h0kL8/TL68N0BGAEdALivaUSYBe5cWx
RwqvYqyehfT8TCBKm840hLdRq9u4RAqwxf1obE4ZYpcrwsMAYf1EwkFsG0g+Z5fUu9kAcvp3PJZa
l1qVg90EzIs+vLMqil8BWqL9wdzJo8LqkkgHnHpsfS/bUwzYKtSKRsSFybgaBbk5KJCBXz62OXq7
3dMItgVvAiMSxtgy7yxfTK9kC7EOq0VuVd7fPTz5Xz07xciPGTfS7/onC3onUDZBl2V1XMh6qYxu
lVOCQCfWMDlecf15LP5nn1A5cVDWr4foIOWXMooGPeRltLAWd0BbViHB9ua+CpdSVoKK9cIwLNOK
WmAXwjBiAryc1iGAgyCF6LwHv09kGMWxGWGiP7QvPXbhfzmAm+jGaNs8imcWaSr76RrAgx8bkC2w
puGBdCJY/xkDxVeWAV/Xwr0ljrrBxi86HzS4DQugzfICjpquUm1+kNA0aOAyDEav2tfK5OJkSr6u
/5KZH0A28M9WZQ63P8B4lVCnO7CrhnoIWLr4Ovi2UnO4dUk5MH/B+6twkRBTm+QzHxjMoqmZ9vVk
DaFvvEMoJ8Jwl27acJ3l4gmea9bS7zN4sivhCcFsDU6Z9wfj/h18LcpVd0Pjc6JirPXEDIaSwSjj
+K8wecSz6UmVJ55KA7dQDxlaaV0ikA95csfnMXmhcIvgmMVxgx+g6OrgzQLyvhkdjkfAwlDkJFRP
kerXYTax78U48BdbFYafjWjSugm0QqBULgyNnZnkWEVWcUy+2FEJOmtv184EI5CmDy8QA+tS/Fdq
huvo+mnATrKMChTpobRCmpjVDoksPSKRAYJ6G1UiTvt8odbOyU9+dqeMGBmHrFXt+0gnupcESmr1
Lc1G5RTuj+AV/RUFpxd1Wv+bO+xEaOXsc2Z+LN2CLTul9mO2L7fjIx60d5GOaYaKvUS0mPSlGSnC
REM/u6VlCngpfx6ljUkUedHdekzNdG8AT88VRGb/HzEbTf6mFRmlcUQXdajcj/6XEk6tQHca/N2N
h6icitpurYCjlvLNjlR81dspFZYogti71cd4L9+s+NSdYArK82S5l+d2r9DaAQKWbuHrYIry/qmW
FPX26yxr5nn9ixGsin0BgbXK5HnRCm1MT+cJ1T7Kvc/8OC1qy5Y7VQmoLqS8GeUNmmzdZ+t5Jzak
ig/YfAQUQyotuVh7ztMvj3febUGWzZQCs4MICo2V4Zul7xdM+50L6PjuQmzNC7Nc2aHEcbVc93GU
JexikffCYTX/3SBu4jS6aW3jlI6OS81OxA4KB1x5FgZx+kLt1ZxOglqpoufa2t1KsBdlIbbvUzv/
SCdo44P/bZqIo58PtZRpdVHRYXbvI6blk5D8H7Ki2yV3kz3+rxOdEcL92SmEc2HfIEnw53C9rsrE
p+yJiWVgWsZKrkfXGZ1fVHKanZxE+Oc9e1kzHdLMHiV+qGJe1ppnDMzJkvnAUM7BGoHYns8B1V5r
g7WHvrxT4VK1GKUyPgTBvTqGukCxOR3GvQcgwTNtywGwEVdW77bWXne841G8WFSBI8d0ySC0l0IR
G+eT/gB/KFxJuqhYAme/0yqon44EtKk43BylcV/0nZIVN4Si6+4nG/ZBQXhgi2vi8vkbhf/e3Lnq
PPoOosGid207Pk+KOPWAGsixceiGDSzreEd/9X8tLv0pD2E4mrF2NhiRxr9dn5lgb/EYodolkXSn
SsH78cp2LoLwa/ZhK7FCtxz7CqQUGrLeMBKEx+8aC4vCfDg6asOJbJEbdiXVZ3lh9H8DRmCdLR38
UhE7Tv8ckrQj442NvE3LlV0WY8JeJxtvHdu4ZaA6/RhpOeLAbGb4bRgpmlF8ZRM14jnpJUf9aOqF
J62htS0i9RVDMJP2sCEk4JBltJqPQywCOMs3Y6gXqE0QR9lx7Vr+PXuQ/xaAPb9KUBsXRrKJ74Dz
bQhT5+kxxt+nkJBY0dpIjP+zY6v+WvycIWm7Uhg0Y3gk4vcHqkSldB6vS+qRUlshmTtu3N8Mmahx
x/v1Z9vZ6DsJ6Tt1XCb4/9x5rXN5XBpK7X67juyCD8Ul0Da5DfAQZxyfc+Fd7PLzLwv51e2c1C90
goYlLdZB1WbwNS1ZlJfhlos/AiLYfQlGOSejEdwSzGE8xqCtermOW5aV5QLP+hR0XsqE8gsCXRR2
kA7VJIDbk7oAhavq0/qfqXv5s5Vn6Qsj910L2G1lefxF9pCV3eIGwSvhs2OKNYvStrBu7SUIVGLM
yabkVi3XJAtvwE8ZU7W062CTxehv1i1r0W+fTb3RtWpJeFGr+xuE/W9gvEJSEvuDJsDcHI7hAjkh
s243LMJN9riobnP0wiC78Xlv7W0aPA2AStiH5qhpqQ0ESHaBFy1uUjay3dUucz5iuAbYYlD2w6fy
OMw6gmbC+v7imXd+pSEjz1DNSOMQWmP/dng45V/ZISfPIdiF7nV6xGRTNT+ob92UjUuENjyu80GT
ks89V5oTvJIT9FJigMAU4utM9wmtfTjqtzAZMIU9pnwYcTVn8IahTWLSHSGrcePAVnBwgqQvQPgb
0OuISZjOQk/uOClX88Xmr1otS1DzoOZ8yxnYLI/YmrhCq2fs+/P7grXQG5JuEv+QoTyOt11CzyMf
zrCtTautxzrJtWalF2IZ3SL8bbouYFCANWEfOgrUhVTlKq1nVFbUVXAE86x9YDAPZdefanYoUH9Y
uyfwEctHXr+1enKlrNDpPnCXI7lm5Ep1XzPOrCP/7DeYNFR8EgHXGWJiDIi8AiSS5NDQfyzv9fAc
nVpf7Fcfc+l759h4TJxJc50ZHLCnDRzcsVI+Hn8+5nztWWq2uGuh4irKRZkxHjtddHIej6s6NKHu
h2OGYOYG9BnuHI0gu40qabcJpw7Sp3ugnyYuP7Y+rS7fZyZHSgUwzLBBM10DqVu5Pi00sG0iaQ2X
RLkUNrTU7MXet+fnGRtGCI+ZDz/1tcgcJB+fsjO8dYvi0P5aFOW7zadnmdZ9ercEzQmUq+0duKBp
ZG7fwfwyEnR/oGQfXlhIuthcvrsjlB6pgDYIH3HBIHOENPdQYRwZO4H4dsd/SywR3/UIe7+aKbMD
T/kMHPnTWWxgPmCtKLU/sefS8eInq0m4VDXUDUWNofWWpbDA9mhShZCkI0zKVCStuDSH71RcDQMO
v1tqAZ7CH/TsfvhzHpjca0AEQXt8EgZlADGdGzcZ5JGCBQ/PTESrdFVUvxihjZpvYqgVPN5SXm4e
TU3dL3oMatR0SFkWwg3bmA6fF6QR//mZ/lb71PuU5/jThEQNfxpLrMSIELOPdUJTbnynJV4sgIWU
/grje3+6JSlUclWD1OmGSajjy3+ZWknd0CPdTln6t9PFN0tL88G0zB/SAaD19mzVLd/a+KoSFNsf
4aqZfa5l5lEek8bo9KyV859q2bgFmmN8ywcOzAJdxbCBBe75/Zp6763/MKEQV1c7gbaZdjfz+NGq
76Gg1WyHbHk2j5Kep9/xufGMyGoSTXjmSlLu8l+ot1CktKFdDq9ysW7eOAwDkBtBJPlX/1yen7Jw
/ivopZxEszxAeeHMiPDtUgHfZRNdCVxR/5C+2N4ma8m3vnuz6lmmxXMQflgU/k335R0JAxbnpnxx
sn+3OzoYxP94RbGoRmSpEJVdYkHwDm+Ee4UZh3qSitOV3RzDWL1oBFDbNhIhc5263iY1mOvVvais
o+7f7EEphOdj4gnEDatJHs1iZd8IxMRdAglGQLBL+YBCMhOq1L5kJMxqym6tOL0YN/MC0Nh4j001
qew6nON/kzP16jTJXpDuUAau1YY3Yw7X8TIMCDS6dQLfpZEpbmAOHYeGTMKDSySOKEW8CrnsvR4e
veaTHA3zyuI85aLEV7dLlOBgnHz6VYNiw7qfXtHRzz9dsP4Cuzi8GTqfBBVuqattbiIG3qOhXNbF
PeJHLWw44gu0ZXMZaFSL6QQGCszFabhM2ERxW1xLiVqCXt3k4P9hsrUWbbp9cRFlUKQPLgMZy5Cq
6QKswiSY7x1qtvtISC7fZLAtAsc8o2H44O8YDhU4FIWi8RP8yEcCwV0CppwWSGIhEm7nmF+EmRu2
tfuna+3/bea4jmDV1DQaIU4VHUstKwTzqwKrUnFwO0F8FKST4vfhSZU7izsKkC8tWN8deHD+VM9A
gH8ebWZXoeoubNWnO1A10m+WCAF2Nq0M/R4Zd+01V0AqzEvjO3lWnhQAzexUEZB30Ptgbyy0UJbd
MmZUeiNzuatEeghSORV65Q4fdgRN4aMaRnfiM15ikZMgnqgXkeTKsBZoWqWF+ezx3/WOp4ERRLZj
YASrg9+LOyCUBePfLbmCGTNNxM/6YCLjpcVtZhW7fJWSBuNdjfPGjjD1LZgnq5tDLTFf6u4D310N
apUUIU5oQwOLmpB5BrmnXkroFoqciwRlb9YcHcvLGCBsbTgP3wcNDWp7h8EJVUhWzTIVSX8fFRZx
/eVt+xW9mLuDbfVOSOG24G2fMqFBo+AXJ68i52+uS1c0VytNB+RWmyw4ctWsxQL+ko/2BMn+hJ6w
og0pR27vaDrOOQ8BHyDpA42dEgMTFsRpva482Vk1n1Hujt/7oG+EpCLZEo3Vh0lvz11EIA8ko69D
V1gyqqSr0tXStrliRSZRQHPPEg5H+BQ+GcdLRJxFbtIMvfi019mEUJCs61vUKGM6+20DMjuOeLX/
5VUQPKLQcxCHsAZ6C/V+6b0LHcXsQhgB7EhysKv2kxQrbDR5TlTKWyClgITj6pZ+jMnXqoaOrcOS
OCa21/XiBPmVNLhTljRlC4sl0PDFDh9R8wcVN0b0D5Sopbdoaafzu7KajF4hsUDkeGqPmVcUYTfk
NwUrEDtnyQJipXQLjd2vo09TRDA7LKEF8O5J7+3byOOUYvQxlAsxAaTWm7mRZXMJk/6LfDK3MzLR
p1A3EzJqa3m+bQSUcv6TFp/wSRIR1tPwuAFlWahN6GkOK7gr26OjXOSUzoxzwm04Kmu6B0bGkyPp
AvIrmcZUjotku1Yh/3ruxJc4HtWoJnpwTmNE1FI/e1caX3b79n7paU7Mj4GZJ9rpcS+eMQdztlDu
m6pIPXnWpY66O9V7BwuGfMuwkjJSmpoYDt9vtd82whlXnOEPrp593rDQVOIo3YQ9FxVsWbMEmgI6
tysUp6nVUve38fZuEjFSQjbTzI2qqzfcQ5GSyQJSyCa0hixmZrIDPzdQ/KMzj/0wNzoQsQIFGmjK
tf0mYjnSHawQa62DlFCe/5KxiaEDMQmaAUaXwOUAj9bD5PS/YNO+uzGKbrMEgma7Z/WP5VVLLAjz
l7NpOCy/NMyiHAQBW5sLvPdMhwGiBVLsb1Z6/fPbondRIc4tTFq7XhxmZRxXBNJ9xiFKq7vuX2qo
281oo5JyIfdBE3W2EVgYLmQBuf/67y/hyuORZORTo9UunRrM5iyBpRQVmGy97L7A7duYReon0agZ
vmpk6qafvx3npm6ymxz/vJhyrh/a4R48ypEjAx853+YZIVqh+JiwaWTZwcrI+KqWS8jSIveezqtq
U9Ygv+9qbxQpC2ZsrACd0oFmRrD+4kyHjsvK3DwaBpVxdF7mbLBeSSGyrusrtJ0xeLPzFYCdMNew
/zLbWD3ySHlJLwptVIGMAfFx/l5Ueyo+s4C5P3oQJqE7Aj2ie9bGyOnQfmKPNXyafTHJ48+bxwDd
BKlagGinOmHWOZOfrfT/RWwsEtv1HzuTyN3iuGNyh4NTP0ead1PCjqD9dAn+gt8itH6XJbOx/1nD
QZ2RRBfn7mqh2Oj/kZC1q6iuBvOjJR3q365oDtwtLd9Bbl7k8ta1HEn73IugzCeQ4dl5cTjNBKic
dOeE+jzk1YqE5XHgZ6MBX8I6SH2qm06ZpbTIpnCJyj+ZnL79yxbLGBdvGVdVsZkBGkGp66fWlwJP
inWHlwqwl3qPFhKkdXXeydLVdSbsrbDRn3PUMfSAu/ut6Ywf8ftOZ06xAbbBSRL9Cctwx5M0afAh
GqJl+Qv9MYypgRYEuSAv5NVKSryQTwYld1AoRB77v+RikPHjnkKu0hTy+XZU0HhcfJx0j9NZkNu3
fk1cDe1RHM3jD2CJVDDNhjSZaiDqH2kAKFyKhuEX06CCJcbKqeEQUlmSnzJNwsMbP/vZS77G9rZH
yfPXf9t9Y5qykxBaajrjJPOLyQfzGd5kJjZuwmwCVxbHk0yvAQXSCip7jiPjUn/4ZEKjCDAOjpCh
hbJVKZlq72dk3PzfDaaxq5Sd7sIxddZwrYOA+5E/xKjzzSt8E+lpqDXDktDpHZI//L+BX7+zyEQD
ZuplJPoe9PgA4aZW0DWBCJeGsmx1ryQDqQ3q5GBaFYNu7/aVbDs2RIZ6kisuDfdOLpOUyks1rFHj
e9jyoDS3eucE2cCP51i56Ay8r0Ld220lPWIgy3FxhwuDN2bVM06qBw6fmvOXKKIVl8PoAsXdH1P1
eH66+0jU7yo2wajFE6E6fec5eKMEMdY+bHaQGdqU7dDKxLjkFTbEagO6S5E0LsKIP6LHUFVeAWv8
ZVB10MM75i+gseeJ9fiQT+alZtt28iFhA1hTcS3UH5TsNahN/4mir8grfuv1BIUlt5LoC5/MQ46h
DDgA1ybuFKgwsGrCKSEcUFo4sFdRNOAUu3Gw6wKFCazLN7iUDFKRFdglhGYLQZgQL9Ueyj0XSjsk
QMIwHL86klHvpaG5aBiq7RyJ6BjE55t7Hns6/8dthe4YFu8I2a82g+xF1zv72oY8RnE/K4FmPxd5
zkUhu8fFnP0O67NBZLXwBnw9OYM+Q4NU1VfodnWRCrPpiUm5EG+ndtjlWJ7JlCTNHxM0tYiVgyH+
skxsUJh69CG1Wms8cXx0yp7GtoDuf1z08Eia2Ih8nfNLM8iRdFwrQzLO1LiBwb2cMyHSNgxikHVo
mEf418GqW7Cj1fwkZLDVUudI/SpJhku9w+koatoQ4eHNVv3kWmhgFx/gN0aoyOV6H9LDc+mR7fRs
Gf7uISWuaSQEMyogaZ/FVmO31Jgw2seKU01vxO3GhXgrXY4W0MsulT+A5cnpSTa+b8EFXb5/PdNA
yNSs+WkRc88VRsg5BlgNr7AO9wSv6CCwdaU1FHjwS7VuGLQ1H/jNfJpp8yJwUvnQY4J3HkvqsJYk
eGc15SW4cBR8Hq2PWBtm0PDlygklmfYiG8sHHt2pHiTup1ejE30vrT4aE3IuevCmZjyfAyxpTdxD
cbRzMKUuYcXUiP3K/QffOBw5yDNGDe3YIvnNHi9+fcvQAaeYR6wepuZ8V8IRFRpLaOiEMaUy/IGy
hggHUr8lET2Ma5nAwITmKYpDEdplJe9fdNcQshDamYTstp4shBUePinuEJyFtjGsqwL3i0SqLnLx
+H0D0Agl6yKt0qr9nqbmTThjcn+O3QVdjpAPH0B15MDISz51+pkfPmVrj6eBNdHkiQrBBeH88st/
IUCxMb6dcztSwwL8VRdXurttkPaLvcIOjqWBnb0CnuC+2PfL1O7o0w9ICagditkSP36yLqdpE+nj
YfA+a8WHBHW6/cFlcwfTHA58FNezz/zEKpnzXtWZaL7bjXi/AQxNJj3girN8ViBW7g1/Hagv0jmu
iQzSYjSl3VbkFFX2YVB+t0Yuk0zfkEfcpPgZFJk5lwWKTTxEylDebS+Bzmcz0ka5/7vsP2oPc9SI
jsQppGUYP5OC+hAGZDiA4yKCSN4VF+do34RKx38+CBEx3T0lfY6rtPodoA4AzolofeN3wG2267Qt
PRXDkOAaVAdWn3S7DLV8hKRq/1bjs7VxzunBFaAHIOygt2touG4URZDaEV5uynU4I9DucqLsx5Af
y4SFs5986j9xxjC59EZUXNbFRQg9dq9/Pr/159Ku90aIqhu1bG01Wz5LdU/bxr+QXzw8tbqd/mRT
T6+HxbtbH8/4NgWB7NkWlrUsAYTBwbZF4vl8QctNM2BOI+UdbpiGXExH/uTlsktqju8R42OtFVBJ
x/N1oZazb13tWp5Lmnpe/tr/rRnCR0/TAdEd7jKIT/1PGOsH3DNQTEevNButOXc+34hwRJlfFaoc
2czqKTOn2HulpKyrmWlsWtDsjJAbyWGLp550Feyf7WrVm66lt9gKfK43gx3wM3pQkNoop9aZBWFC
XZX0xsik2XDHcpH7EFTBxlXOsDowv8bSLeWaXSE1FpdM10OS6rJBTnWlWjiuhs3qawtzkbFGBJ31
JOSY/K3rkGhpdt3kxlRAOwxZcpzSZEyvzucvIzig34or+kx3nSSQGXGjebuXY5zfL/27xd1wXwO2
m1UVWHA8mHzuMxkC258HhbgabLbUcrY/14s6KU75MnndrWIIWyYZ5QnT8eJiMhNlzN2Npg3S6HcR
gF14Q2TkzAeDBL62KDAdGJQ5tWM2JtEDfMKtT8wjZBqj4ceXCZvqUtdqe5ovWWxi46L/+RLKHbbp
iLRAbevTDbsCgpMODMRlgcnpV89oEILI7G8sIVdlL3vu1f/AgK+CpU/lCEmaogP9ax7DgDSP0Clp
uwGNL/12LDKgj0fdJH8kTMyq83d+/qoVnf10HCDcLvwaDop5eu5dnlsftpYwgdrQwYEekZ1dRp5Y
wWUxC6yoXfprHAoZaQ3j8S+pfIWmuLycLTjWq4sfYMAfA1+Jy+qshxa2vD87mmyljGLX5xtTRNtI
bXxqgjW8l4wqBwbz8MSZF2aI8QGhuOQipBvHlrFEAUnGhw2KAy4dTrh0pc7u0Hl7e+c8VcWsDOum
KIAifq4G9X3vUrQlzk2JzI6TlOkHYIaZcX3KwxVEElzRm7oLLSLyayX1i2LDkMtdnzp19yHrVkEM
PwjpuigpgufoRkdKyvm0NU1jzSZUCJ7py9dukhnEQWYQaUqaSPa0l3Ab5DXOfA6rhZ0ktPjtLGI+
V1uV4cu2OAc0ebX+PKUbCOkHhOquTse2xPhYI0Va1NmEn812u87YxTxsVvoxqSSUmX06IkJn9xB4
Tvs9+33ZIw3bCJkmVVda3XcioHLckzZ6x+v0N7DK5JnPOfZyXg194Eg9AH/xu6W6RMJlV2Mr6OFH
7w1j9aM1CpM6InqbVpyvLOncURDKjIh+9UMpMlT/KVwio5pwdG7GEY9mDp2N8BZVhUZH/Yp30WdV
jxoa97Oo+JcAAgZMT92gOurHPb/Foq09G/3AnFzQNpT4SXRtK4Nxr0myJjc+v7A5UdCt1hSwwzIQ
GWzZFVuD1UVrz3umaXvOsDdLZS45SMAItXCm+IEK15Ut5kzT+rUDJR1ah2Kl7WkJcPzXj9YfIkVP
iUAV24eqbY3JnIiaD720Tx4Du8vkjO0FUCJHV+98/2Vjl7LHfrX6D/Se4FMlL6vDuAGJb/IEVaL/
tmNe5OCgXqfJsVZRQs6K6OC3xoU+xUUnJqKmVp5TTgKw4541W5sb6zqzMoEoglikQ4jjjTLy+dci
XrRc7+9X0yi7UqgXDXY+yIv9j8sGD5jbZA63gmL5SFotTK8f3CUwPTq5CQQVAnNfR6FOo/eDEby7
ABK+lZljEt0loEO2XFFDzAd0hDr1xujx26ZgV+V+lJIIuQw0NycnLS67M5Hpk4QmfSityPXbI6CB
qtBw8UBKQx65owfw27g+oKdkZZHxHTxSFQWLNFFgyYIA7ToFbqfEiTS8cKsC90RZYowE53J/ok0m
2XmIx4UUeoX8owrnAlZ+NTFtDX2TG2j2gSs9wOSxoEMxO1vMA8cLDJBEbK6eFA0cviV+r/0sH/eZ
bJNyV4NToIGfYTr6RzQy8WqA/alKulfY7VKzeAtxbabxfAqU7fgHiE2Z+7XBE89L1UYLHZTw5G0A
4KSZfryg8iK3uxq2L5nnAvzFfsRJRc7fLPoNs7rzfCI/gQBfsPs4TTFvkCX1ZEbaHmCbjEyt4S5C
FtmZ+67sCBYgJoQyx8C8T703DWbCMMwF7AUY5Ii3vA5T2usaKHF1MHm4y3U2STzfvRe6G8ftG0h/
uUa+iCVKPi5af8HPkMfeE4YEGkSk7OG85dwGewah54GteSbve1XmzM6yEi8Qy5w+qxrjWyXbfWUY
Rf44h7xbLhOLvoovwK7eWIkioq3y5O8XBOaO2tlNQvEsW1X2tKwQ4QjZY1yQ5b2eH9kQ5xcvVJNc
jq4V0fwXCbKk/vohdUJdyaQrYlbHqy2VKj3mUcIH80TR5TJxmoD3+ecW5qXeQlB8OhBEOf8EAtng
YBXbQsphVjFIxmfGS63nN6Ayq83dUHsIUIW/IhJ46InbbXcM3ZGDkridp0ZAd5kQIaR0fHR7oikl
ybVeUTZ45fpXc0BoQE0WN36+xH/w2Tj36Q0arb9CdlgnC6oXXeO0MFI+2YZGvIWH2YemVIPmx661
gL/qCUtyb6uNhdE/VxT6FIoBxPmv/dumrmwFrz+TAb8N8kwsQoDB2pG3Kp60pdRb/zYPWDhLRsV/
z5wT83eqe6481mUsckGI+XRjeoa11244PW6hm9iyShLIYpxAYYlK53zdRdXilwLDHX3SKeunuNiB
NZwy/qIjLIr36TcPJjVqAS2C0s7atDDNVD3/JUkfi5Mx+CbGc0LQLmY0Y50j4voMpVj6eV0zBs7j
S1zfhn9gtndxvppNlDFO42LUR4Tamq/J6b18Ry1kG3KJB4Daw33v3bT861TMZPab3BJUbkguFA1F
oFPgm+bMMVEGxtNWSZpqPamuEPvGEHqZxURwg2n/zSaKUIARN4BpMh86fIr5H6LtjSxCBz1dYad5
6QgubXCCvnukUGHwl/c+pmkJTpBiM66XBV5yDYEy92rd2nLuBwRKoCDqDB5FfNLqYtc4rWQAqV9D
6QJrB5auEi4/pBpr44Ik19ag+ntRCGqybcvVWfEn/Ql0EFu4KLuBJL4ELVlMxATZAjZAvTZZ4pnk
P8zfmSBIY+0XqUjq9vALGp0RgDtAmIuR5XSjF8iRxzObdxlYlKbIiIg7NUm25F5Rr5dgm4c8qH7/
6mEbQ1bD3dyu0evSnUL2WVkTob+1Wf/u0H5f3I3E+JOh97Y7UTNLsmAIBmw6uoow5cx87qMZTxcN
uh+Z2X9636pQcUeaQaCPwrGPcpN0RSl5r0vH5LJS2bZiOyEqUiEfam904kZrPFHF1Z7DW0nzK2vz
KWvjs1z3QuL0sJluttzg3h4z50xHb/EL45Bheisf8+bRos69t2d6nkPw2nOsJRfXewHbdtjp6DiV
rWKkKYou4mhejTup1BKbDnIDrKrG9nKqBPoswRXYxPLUHiDXFyx3Wmv+DxeW0Dxm9l0w0W7mNta1
8CjIGWBDfNenFjypjzd8aEvO6gTveqYE0NJUkwG3qfDfZ8VhxSzAipAZIJiPkktE5LV4QEhy0EuO
uWvdXRuKwNmLbqh4np4NI+tRVlhIEvifo2rei1/OS6GIcdqv+njyq2rG6SF8730uzK5Zq/ybb0H8
+upgIorE5nRFsgvalc0ZstoedMmE84IlP7BbhJ1KjGAKraZPEBmqvff67dTxJqW3EnhtawvLC06q
QGI76O3K3VRCmjlV0UTnnfo38AMu3K9Gmkeaf+h2kB2oBIQKSWiraf5YxzbZLgUjuPodOM2wllo/
FaKMdwmJVmqFfOsr+J1o/crjUnpJnMgaRc14zrtqJzl1aS//OBTR9IlWujCDNHReRXvuoSUTMJLZ
SUAafGhT54PaHI/unT+r3UJB5G+bMkZltEBGBNprGJ8CYo/PHZRtgLosv2vFr+5y0KO/gg2c3ROH
KwmdwZ/+anm/5c8xu8NG8422xatG3WxQlnbTBDQKnt7Xx/noOVEb2Lw8GMajqVY3Tcs7CoQN/6dS
oBpOqyYiNwhh+I5SovUPzCNs7HlclroEb2ZkM+S7IQ15PZKjYTA53eMCfNm6DEmvekZZor4cLrFY
ka+1TSPRt+gxuz/b9253R3D5f9PetewKVd7BNdFcB4IChJ3WXR5BekGUhNofdBYWB4NrhH+lIEYH
RCjmPKsqajXyU5ehrTlWhNWJMEASUAhNR7ihfRJNOpAOrboqsgtDaTxzrElPoQBixe0kk5y8E1Nk
fq+TpAtPL/3nfHHNWYM0BloI8ioXz1ypX4jnacijdoRQtWyjL6BixZFZRpeovE7okQwkc2YH5heM
jWaR/3qotH9p/pUoYKBU+uUQt4FVrDJL/1GhtYORx5YLevWvF5GnbYKMCIvXdQkYQjAtlrsAnVgg
X5kin4Qxd8jeU2fJ24Xdc5P/B9E8kdhms/36EG2rdzKVTT5kc0evU1xiK55slLr8KQntmLMZiRrx
lB4ngG6OqjmrR/7A2OzWrnj5PruhpkcoDL1zODXXAMgMU4KBAtwQYeZ3D92b4WbJyBRJ7xyBmADI
0hxe6C21bGEXMTRR/p18s+SSGSgQtiy6w8I61X5LHC7Ht4mPA7+6XNVBjiuLxUOb0ZWe+eJY5niE
5/4Z/+JFn1dFhxv7Uq5ckOrSceCiZ80eqwlwfSFwyouzGaiYOcTLrULkHZT4fowA2pK8pslRVJ9D
V6wSuT/kPLhp/SlQi5jCNDmRxI89plHu0RMgENGpN2+1ITeycf0K6UvgpINklSnDsPzhhSBAL2nA
P8Jj9dMMfRaPziEKMccJvM0JIPkEalhtTp3wpMf9Q/1GgPm7lPjzYJUsgr3osZbp1rHRoChJ7ouu
WVRTi84mHY1ZNuwWUXH9jzREXz4kOemDX8y6AuGonKSf4uOi8DFyrtF7wAp0V/IIT9uhXB2y33Fm
RIDicSk0bBulbei5RprGnEQcLiY8EOXaRnSa1+S+2abzdwMoAbN8c+7W8CpoK45+MD1jAlb4YkDm
XSR92oacLNUclJdpR47IWIPOB1Hr9OMlaJ4734HXVamPVYLzKuiH6NltdkNSKemuQlEsK/6P5sEA
q+GZRl4D5CK84nYt2slDR+fkHZ2TQ39NTHNc5adCBkuReCtTsu1TStLiTSfuGYDyRWFDohtMLlNG
e2yhi8B8Nr7m+bIOAegH1v7qCeJy27NL38HkiFrjW/35aiJ8+nTmbrb4Ba92W+18ucFVXaRG5OYw
8XVoXLiEnWnDd9vz9Zklc0ndGcw/FmLPRDtrMEKXb/+mrDlCqLt4PtbWs+G3LqHavS+dVE3gnIcn
pcS15avRclEiIxZzoY4bJD0aSelNcooPxErUWETEy7BODAw1aDujwIoxmaA8AxO01uOw80PLOs28
jd6TTO8SVrXaBhPIHu1bHKhEi4eNjzGWqLHeKBoL03+e/BRI/BmvvJmKUmpJdNF0hpaHMztZ2j0/
xgQIeaQuvG7xfVtx6udabc1lYHYEcMnjhr/4z4fq6/hnzn2lbfUcfaDjhCvERPJEGs+XTuwZZFNI
+iqau4TuS3srWDtSncY4queUNzSUOPUtNVbqwyREHEvX/Sn9HSp6wjOs+eHKgzk37fLCeWdCe5Bg
jZAV4tTIQ+uNM9WsU+GSvmq3O8R6wi7aOUkzHQk3mg1MdB/7wTGzW2ZyLa8YlG/NC4VY7dG/F6CP
imMY7JfXHDt+Ej5QOVsp97OUab1bu2uVVn81yVBxzPv/fK94isiTQjyaIvoif0MonpxBT4Sap9Q1
LC1L3+9Vy5m9NNjozGr3eLwZ/OC0kngY5hpzVj+NmNCk845IdDRiXUM6S2R9StOTTjKHGHFkgPJV
XJFc5rzJcFz8Jvlu3qsRDtLULEgmqLTaaDSQI7IJlce07uuIEtRXrpPrU9Md0E4arnvp7e7dYBBu
KFKoMoAaaKkPemTrUzmqFKAj0izEm8RogHEqH9cWQSQmxo2WHkM1Y3ijEpZ1ssVJtJPsFdykjKGI
qpAlbGeJT8HOrJAfYVys6bLNGXfPfOtCYxsDykkJSa7HdFGYNsSpdiiWEiCdPOpLijYH3d5waT/Y
DChtUiYo/97H5OeANlbg+TrAE/O2krjxtjGYph9O0niCfsqo639jhxAkvqXpZrDmBgXDB+fyZ1sW
S1fOkeGYh3MT/SSdEQPSHbPsWSmXJ8t9djRjTYVUjH7m+qodMWSBFmctcQTECVoFq4soScqtF5qk
gPtUaT4j++GPj2Gj0kIAdU0vBxFF4cpaPmJ8S+zC7nKmDGGIPC6epIQLmiZKfvVdvqIa6JaGAl5b
YtCIp8Xq5gOoluclEEfq+JiAPGwASmnAORcDRkycTeaD4RkQSEDpgHo/70ke7MdS5U3FR/iRI6S7
gM/C6D+CQdZT2SXeamMIgIhRx0+bpPU6CZ4zNpZ7fJhl6rcU/v0wq9aBkzeBbsyAqKSeAycWmTDL
fgndH4RT7TpyiLyyP8hPmzwfDd3K6aNDSh+8OG3GoZCJLmDgmu+S6NL00fPmrwbYY/DZCziIMNEJ
O+2mfo8W7jw+WteAKNqg0U9nlnvVXt0osYLE83ZJAODDubDcqbYaYasgF0FUC/3UU40ZK6O8scyX
g2YTXyIYtSD63pt/peUAVuSB52BmvgcSZfFiI8UM1k0ticHJyowd+0RLpzJJiBW7g9heti8QOUgl
qijDJtAmzgfWvXztxfMKtsoMiSgDWfSurVFPSa09bSdrCwnjw1548TyggbXDdun7lNqvmQZKjm4B
dEHNaOldz5iwz9aOUoE3aQFrA1Nw4jIZJKbzATlvBqhODydB6/IiZ9gBUablHP9Gp9bfIes+qAG5
+YK2nYihFQjD1LyexHxtAWPoQJv+cmlCAONWjDuMciVe6j/zQhltPSyC8GQNEnVfGYi2LGjhRSqp
X1fRe9ZzyPZXA6AwBtmLTY/B1UrKOSB2kkWDAJpKjEAKIdm1qxnu0JsAPOdY8ePICnLfoVryROxu
iHeEUCZXNvSj8JlngG5aDPQPHcwjuEP38ned9EPVNHHUXIDvvPkjGp7GaZaKUMc3Et1RIE74zNd+
PDbUZFtgzGLVbaZsLp6T54+zwyvyLhvRUXmQTO9HHz0VowKrrIcJcjHpIFljN4s+1GnLNkDhD4N7
EB6wUbylKYEf+Z976Mii4LHkM2rg/LNrola2ug8ok1Qtc71/JswEdqYIUPUPhTawhg9jMX0eD8un
EWwx+h9zGZ3VGhlVVIqM+gVKac8t54spBYppsW4eFEw+gLwuqOLw74onLo54mDIz/jHmZwWk9s7h
OS14EJHm+r3rFUVMsnIl9rXiB51NAxpXBw4DpX2mvydTnR43qB0/lAu7Vu3jjlvTOwYg+M9SCLGa
h8DK3eHyvdP/bKoLbiH5CavKYbphApi20xX2643GRYfu+bHwJrGEv6LrqVNjzrZRkCtozSZunCCl
A7KY5iVdL7KNWYWxf4Ii9NaqIUuHRFqQDVndwTqy+v9EWaNdF8yrAnsgel9maZTWsa6ZDCOoZ8+e
1hyTzBu+nRY2CzqklZnHmROsVto+P6VJDNJ9N2ic9942BhavAuL04JjYhx5I790LWvQOH8W0o9rI
r1ZjGhJjFZtKnMrNoDzCTqCvlkjf2eJDvgHk/Fiva4lG2SvJS/hOvX4VSPXF/aZYbzN8bSZ1Kues
vF8a4ieInBcrDjBM5+UCT/0gRLKB96Q5tke+bP03nL1VXAnlFO3u8N/9Atw5Jt4Wkk5CWtXSSHNm
8XusOtJEx+Mo+TxxA5EB5b7mmFwpW6MNZ22hm8eydg3I1C/eklVpmjlO/2cx4FLh0dB81+fEr7st
UTxk9KN/Bwmey9lJf5tl6V+LzlAYQZmluvvJkUDDUmhUEhof5RbLKoS7nKsTxyTHJuZqUA2nf0Il
ShCsM2GyBuXJEewJMtPTzYHr0wfLwT6oTiIwpXhzgZrFjtBf/8bqbhS3k8CAdUcauCAjRWi/Ua+9
6UTy2QpVNosuRklMWe4/TJGAFXwRps90sLF44oXEB15hnP3TcQwx0TwgASGAVp6l9PlrxFAmvnrW
A1UXWtaUifTjDCCcjUlG+bGFR0dwPnkh18tN5gwcJXBTxmC7V51lv3ZWl8UYh6Jg72Don9N1mK7E
oN4tdjHKebWX//fNprT1Mw/j5PkEezMP9+W9Y7PkIiz7QiMR+TOrD2gmMtCNXWs+3eJs2a8ypV4R
qQnxR1QJL5LNgtZwwF6p5GDMGIe/SIGh5pBAqwZPEmTC/4lGcH+xnhlJA6qHcaPNhyjL6VAOewWW
/Uyz/jqloIg1Nw5WZcq1QDWVaDOCLBLpzz9e0uZQY45ch4tGP9Rm06F0W2wljVaYiNE8tMIMu3M3
CA3R2ztgYqlhJs7yBFXGxNQvmkVF5CyqWDIVG/E3NUmc4beCsRhaCQQ2y/METpBM/PCLNYo6H4QV
zu1t5NhS2DFCqTSkX8EMoZptwPCww4y0pJ0vtaPonHPADw6itejI6Icvc9VW28CK7Ql71w0n8rop
sCByBRDEfME5qejgoHSW9pNLnRWgnlFMPJf3KgcswKddcOO6sAQcSOM+1nFk7nMvYPoAKjbtfUXt
PJICItL7W002yI8bIIKLKNCk2+ftTvF33Bfe07O+hCQ2k9s/crRdgTfJ5fjW8OJW/1dUujqijbIO
QMohJFEmd+1azy/02Shcq/rWhkLRb3QFl/YmttQ+TmtMNRJslYn/VFlCzoigcBs2PHo2NJO1xIiJ
mDm2qukPd10UKJQ5RzWyTTZOOnaAKiDqQF2GSv3SvkHt8QDtaafug3xWV26m0sb3xwQktATi3bm1
8/sK/8iR6YSsHFQw05IdERwP+L78KLueI2ipEFu+rR58vTkL08K0/NookaJjtgKwB6C9vbkFUQW1
4y9VTLZARDGVexOEHeCgFGzeE+k0P4KyQTAJ2gCVmClU752GJWukgT+lUrk0gMQTKS/Cvx+Svs93
jFqT9vLny9UKvVXTyjGQNDE4Tv3D6q/DZJGvtmJdU6KkKeK8/+4cj/6WvsFJMbgHZyPyM88P5tm1
qvj9a0CoRqfAqsyCdQMo6Tg3o0otAMKMEIsJYpiYTOfcPOKC8scQviLB0stBzNk2XcbkrVgDNqDt
y/XJVymx5Cd9H91dKYmVOScQQurewQ7TTTNeDCJVVDV2bePdwDCw47z61oabeYoLXd//IZ7avkOJ
4bX8OtgAz2sZ+BfiZ70S5PwpzbewFmZAmu4+1LTyt04OsGuNF0YguZPDGRZbDLb/HnYbWsse4SKa
xbtmjzSiG7klj4ujTRC7AeRfu9Ym2s8EqaWZOMjoyk6Qheh+lgLtC70VHkwdnRmBdby47Rq753HB
uilpmtgWQKCa0+vO3lQ/+s4VY2TED2GYt8X/NA1rlD9furLkiG6zYextvKnECTER71TNQ+/qsToC
V5ywnn32ELMt8FQPugbINEdfjT4rOs4oas1nvsiaSadAHyRgIQN3c9/6tmeaec5e8BFTdgNJJeKD
s5lWvsRRih1ygNrOVxifELUwkYfemDUS87d85piRAOakShj4xAZe2AlGYEXVjYX4XwV/MpW2RGpP
wbjoYU0f5CXz+rjiHWAjBGhkVwclA9s/5mBB5EpdLN3zxIzdg4oFsccJpkFAOUnNz7UOZiCLZfN0
ni8K3JdGZY3iUiXB9Nd14p+/Go4CaJxC+Z3+5thw7YiM6B65svgALRWgafwdoL9Oodf2e3fRy2at
9c+rPK6EA+QP6df/4kwByJxUapxxoWoOw48Bk/2n8xpPFS6SvP04ksUbqlRV3S8kgo+0sPnS+7mO
HbMT+LyBpVOM6StwXI1Ga8wuwQO33wlRsCQaR4HEhw7WukZs2mbIEbZ+SFgi0acI0po7XMQ99bUi
KP+Jzt/GxDYWSkHBahl4RDe2EVlmQGDiYkqo2Ju4jlF7PX/Ss36uDfgw7NJqM8stGEa9/PfP3CvB
8SoDW8ybtMczdZnRrGmYSrRHgjPOo7lVfHS/6FC8VTCvlWTCimaP0L7RhA8ktrX37+FdNY6zsHFH
RL8fQGYpoZRX3ZncW3oot3Fvg+ru7jRqXzD69HB0mDUeHJGfdUDafC2j+5cbsRIK4kf6xLaxzV1y
yFinOphJVF3+n+FzSdlWLsjFxogzW5jn380eBPhZsiJSPzGzA5EdzYkobn6nEIroRcJASvCIFq5i
foPZ4j31tWLmpJnuyYpXnRuBp5gtVXOzaGE8oLJflxI7O5ecQIMcH6te5u0NeXiwEJ/uCbNWAD2w
Fdhlvah4rSNgXjoQHCNP+UHhZER6HX0LuaIjhi/jKqI+VNqDlBN1oaXHA/sB1g5J05UgrILN5Fa1
7SAiLfvTZyrIbDob/wsoxzBmVG/hn+rb9X7Cswq3gGXuT1ZQqbEduj+rGlB3RrJDREeTeZ+61Uxy
l8RD0hZv7K/2WvrM6kYI3Ek8zcuP+0YWZXuGmIypJsFkXLCor+bpIkSpRcXEwXuk8rHWzOTKx2SB
ejdhpQk4+iSx/upiz2WTPM9ByxAFwGD3VL2a6pIxez+PV4uD9pv64bnuQpeJSc57Pw7GxqDVjix+
4VgewviHgbo0WsJGgK8KothbUupD2mD7wQG9WP01q8hQd4rgUTZhBNCE0ZilgFvUYtiXTvsYRuAl
iJawSLOodSbeGQaUJ3yF9xaSN00I/RqeZKNHyDmAt2YFYaikrz4+tiOYYL7ogdj5ZPPsgaQWlRSL
XWWiR5OFNXFm121FgtUZ/SGK9cZpyyy/CVtsAED0xGDlxPQeBhl/39cYGyP584dw9X0tknmitEAz
WE+oQBBZeaSH5dpA8sKhqFX4bdTsxsQQAm8dXMnirN1Gi0QZPvvEPKM7U8GtbX4RUEowNvWfpWtW
EtMgn5GpFzBUzIAFMHg2o+pKmk/Z5lPBLJ+5oQJmIg/84PXTjjwADWWW5MWPMUdJExDkTmzKd3ge
ZrPAtl+N6rK2K0k6tgyp9wiYno9yoLOTk0zsUE4qfR+NnxzOB5PuiBN4qBmYFDxqbxBiuHagozwr
AGW6lvieVnAZUKcEYJ1gAFH3rTQoy7rv+1ItLd3UekEGhGqSH7u/rH/GSlKuPuK2ILiH5zF3hKvO
p9FMmFXj4RBwcP9L/VYlmdSPvlC/l4eDSHScr8WBUsKHyZmRcERQ1UpXq1zVEzYtlGsF8+aj4MPZ
MdHg0Y2NbPLIAzr2fy+MumWcT7nDspdq7Cuu+G8FUJfzsvyUhpD6/XPOx8d17eX9NYK4HezKg4XF
uc6V1Wopx8QOrDZboSaGdFcq//EH2dqOKz6AtI+7oJki2CCbmNFl+wBNSIiZJ8hAOh7wGYdm/9YP
BXJyGY51+7tI6Pb80gDb5iyC749823LeO7LANpM6mvDbAImFb8ukjcnrS9cZH4CBbhu1QaxU1YS+
YcL+XqP2G6GY0ozN/skU9ly+p1nXZhe17rVvNF1rwLp+kgAsGYIWaj1pAtkHtQbHvKO6Ufp+f/sW
+SMj1JAuURs4kQxoKw2FJDv5LU9BuX7OTqvymueLqOgSUa9XPxAv/tUiRYitidkdzn75sm1e8r0r
PWhGiRYNyqcT/0A944YgdCO4/n9Jq9D4zCOX23JeZVwDGVb///Ww5QZpOPbIiGPtVuSLeXYbkhbh
eKXoBRj4Ew3kJQS+47n4+wdAXGufjyqjIAz6OVEXuXwMnRGKxglUUuerJNT2ZD1kJAd2xhymvlgE
xsz+q2FFO5A70kpvlNiqcCQ3ToqMkOF0MXw6oUBUrc2ahZns3YAMzrqnQwJGGx2XCPUnBNfYAY+s
x2edeIs2L9Sxmyu1WtfgE/SQ8ZkddNfPJnRJ89GBxtHmIIKg8oPJWyxNqWoK8PGIudCATOBmxKGr
Yzchmg242t5qlsAh1Z/BDmSfZgQ58h9eCN+wWrm590vitDsXgU8ek46ir9DWIzdcwE56/D0yxZFD
GFTN2ILGY6pf5mRM5PNTUbS/Q9Km5jiDK6IgrLc8qBlPb74KuJSuGN+Gk3A4DbqSnaSVSh6wRiwT
0KXvN315nqxTrbmUpmPTb14NJ8ZTeaBcVhSj/6xvqfxDgjY4rwAYX0aiNhIWiq/o9wofuDFPK2JD
ZC1yYOEIE2tTU4yaqRBykrASgDyu8P6MJzd7geno1TT1iotQs/AivpaHkCgzQhiTK/riFnU2VA13
U+J7EsfbQ1qbJyC0cxf7pZzrv9XFFtauLLqN/Y7KZV8UJ/K0AsSFEEcFJO5qxUvvk7mrjERDrqqo
SdvjaweKEibcdO4PE7DRljDFLqT2ZoGUAV6mbEhhPmxmpox6GNpi9LfyHeUvgZ5Z4SQH7WQ3bneH
IwnVDrGbp/PDB6KZTblZEGE0PSEPeNP62etX3Jxv4egZygDOdtP7xRnkjIP9V9KSCfhDjRf6luvP
DK3iwpawm2/5RLjWN7OcudQx0Wk5x4iSZq+Xoi2AJVXLauxgORaa93d400BQS9X32wjtMoLXBy/R
vyEHp/UBEjLu9Pdjyn2vCcXYZ5U7WV7t/hnbSMeJ2jg6aPe85RNxG9a5sJPaavJVjAPqgf3CcuHl
2oC9ErtAfHPOXTzGh5Bb/vI+/I+6fHlCJsAN7wLfSsRrFhq7C0zlrLJ1mtlacGEUVrDosdBR8S7g
Ynex9Ljzl6qe8RgLFSgDGcXo4LRqOtzS5tCZSBoap/5HLzi+BnP2Cxbly5nVmdVxKgGaOY+Xu9KO
EJXaODabcFdvwNExwA+uJdBn8Y0Gvu0KNmzHi18hlIlV0BJNrtsTr9Ylkw9T4sIq48GgQpSB2nyZ
5z+1RRnPQXxcP2B5AgxbDlW6KJGRY3BG7ee6ie0s1T9llv3bqr9/Hhka4xrmgcJboKH/JzKSWt1J
44M0PyLZpaEgZH2Orwq9IGo8CaQYzSl/k0ximSzRpw9o/J4YQ9Mrg2LeGvQ3WFbRgYRf/0dhhASk
iW4rCkQQwvjY6GhfzOslimsfLv0e/3W+1Ch0JxE3mbgqHfKmA2wemStcgu1YjiCcmXZ85ISLx2nf
EIiLJ2P7BuqZZJSkYDcfC+wJD2/HzXRFMxsp/PRsliif0c3C+1vjZJB7uZmM8Tk2BbxItLDrUo2o
VoHr1oX9DCQoJLKxGpySXf2QxgBBbwCTB0OS7/0dryf6o6RwgOE4+cEz0ZQJbRB4GcEYFpSMWbdY
Y144NZlyCrHrT03QVwJxV3DQQLUGeeT+29B8H4xDECeqElrIDTFE0RkDAmgIPpDGV/5pNKhpqtdZ
51O3nvaRVrp+5Q3fTZ6rBZy0pbJvW4413x42WpG8oKxgTMT2kpaAKXsg/CZjvooVt0MjmDaqPIrS
YDEpe/MPfqqROTnS3+sz/4OcBYl37gPzk7vCH+Ygth9vgiDBhXK9b1hm+V+Cfc3wcxQjc+HRi7uh
5lT6V7k0AaJWE/DvT5CZRGNjNJkMoX+rRwtRC+AVTAgwitL05qYYwLWZnZZoIaHQd7agusYubkDd
Ae1Fni+VRGvfQO/mGP/3rCgspIvprkLmMSLfnzYSlqHTtiFQIFVXjVCnpvSXRxvVuioXepYe1er1
oj4fojCm2Z6+FdgwWtzf3mMCofiUBYMWkYywwGvIA5gVgC39ZgcBUlhr3crq6uOI19WoXtu6x9NZ
D8x0kQ2Qm+E4PtWGAe+nVVbegIGA0qOFDkMHuw3zEm2lODpSA7S7VVleGGz6H+IH5mQjBjiHtV3s
UiAqP7XLAwB0aC0AORCcaalDkCGT/LEGhcClwUwWuVhkN2Dyg9H/1z+F3Dv0zib2Hnbkb3MQWEA0
/bpaI/B3P85ojR1uCpvUXR3F8is2eygumxgWfrxxbIwcx4ryV8R17BqpB4fWtB0zMG/+2Sm2Q9Nl
Tmay1RtJh+0eAf4A/35yuWL3QVsE5f+ZnJcm2CWsnQHzlvY4IsFCGIcqkgJbf7NCuz43HfrsIONK
CyVGy1T4hSh5KhzdPHRMj9XpM8xYVL7njmPIvDlE0K+2jjjT9SwkZJDdoerXXrBwz9ymLEwsOmDP
kwK1cTxid8p0LLLdaKPjFDzX4bTRN8obUkintjynG3MWl3goWjgqWamQGXSs6FLR8oW9q9LPbpr9
blQEK//VYrQEOS2B5LqKZf8GU47H1yfg3a7n4VHJ+Cq2Lpm+HlBo5ZkN7wQ/PjF1DaN4BTh+gUr1
5+lv/snkSk6xVy2kwMWcef2iAT2I+9ZG7qBsmYksTzU6nxZ+b8tSUwnawGFTiyVXuqUvgLKdSObn
DRdMlVIkNXeUNKYWs0PZkCNdxdk/mjXDsrbk63lTp8Iixvfti4Tgd62Ie/kPUYQTmda593gDyxJ7
bhfcYDqE0pcY6sDWOQQUh2wsX6Owu6D19+1WbX/CYLXjyF01k3MEJjQADYXesCMbu8CM5SzKzp94
CqwUZPeUh+fU2kDLwyCbuOyF44JrzztY0LdZ6P7b5x6OEE/DfW+o6ZY0F53Jnn35n3yROT8PCIF6
EPslQU39N8JeUMEfkl9R3VzgjPKYamyKlVv56olkdcZ9hgVQ2qxFWpl+g+k3qxPJQIBqzIpr9o18
dblF1pDc4+ci2W8h7lal/3TXrOZKgq0IcJfNEMyioH79THb5TDxhOGntbD4N7pDng7zr2f5jCDUl
gnv4avXuvm82EDJsNiHVtFHmbAbI8mAmI6vRvZfVW8prWMxlUmoAltE5xeGcAjuOHavHvEvOxlMq
4+bltMM5KaTkAVdRWLaIn0SRBaCncVr3+WXLskNMDy0uc6235i2KAsfi530wGCTUGl6+jAOwkA7G
Z6W/ZNy5WeBa1ZmHViszVEHFH9/lj6S8kOKDHM/SCpQM/IiiJNWzit3wwarDAoqTfMYwUyXbuouZ
jUqVDPOsjyFRRKOu5Xj5z2Uds4hKZ5MHzpcMXLxvx5GGcdTtYgxjacjW/xB6CMdhIbn9D88FW1F7
2U07wPUy5lCh5thpxom1LdipqXYzNvv0tqOq0QFiza4g/nm6psoSR1SMJTD1r3ReMnQgUAtfo1r2
jnrjlDBA4NrW7yr/fh1GjwneWXyV5IXtAgTo3d1dI39hAH0aEnIgcKQ5Aj0boa82kG7A7O2MJBCE
2JjuRJ3nsUcL58ddmN58WQm8+7LxNp3xzkvMbWXSPMVhLdNlxzCEAyYjYoxrR2U54JA2hxygifqA
3yI2NxrBlWqLVVo2eERlq/NsDrLkUavJCyxBE78bDpKd1GWeQdXxKifurQRIkzaEgBIoF+BUkMfe
MpAO0jMDkZ3jAu0izZEHRz3diddLdVcaSw2J0/ENz9ojp/m2A026jz5kKSz+Gom7Y+7BFeji6JmE
knknrg2GDreiIneenLesY0uWKIARMvJO+bl4+hQeh+IDGrdjrZ0Ku+1uB1XCB10kMApLIUTVtdyX
iG5bOcitfU5IlF4OMAJ9raTbiJ8tAOctGOoe9pAGdoGIgx/Xr52idC4+3thA3LMKmz7w9ctqsjtA
Osy6FOSHO+gXefvGfYMxSo/ryCv3RTGhnivA1iry7TVKbHD4HT9lqVUh4M1eFdH+Ih0PmE7qkOb2
GRswEM6S5VqQqciUv/Vd/I7U1CdNgNos31cmfZuC1AMhT/kWKEh13IDIQ/dilBdy1lvRwpTBUENG
wEdWNmhUk0cPVXCtqZDNfvv7xlSYo3PEXlMgaPKnkGXA1ZN5S955hOdkNS5KENGvkTUKhGahc6gx
fyEhmlOEx3yv9Lu0owr9H+g3j3OSJF7fT63eN0Gr5l09+3JVvItD4BUXhI1XEugdlKMnkBDx97W3
lAupmQiucisLyA5/ebnTolsxN6nPiI7Yt1BZMFhia3uN9ICnYHHs/YqsW43jODECXovM5LQWhzOZ
Ncztl+IUY8j1vqkRgcO70iYItCw0VGFDXvYjA2bBWy2gRtsTfEkrSihXvVtSimEzUuEMW2Esga94
T5WuD4tan7kOe85bz8XJDKik0/HOBTON+MMDvJWBrlMP+lNeVkzVCC2nLFXo0wVhTTszXX1h9jld
QGqFQeUthSOpS8XdJ3VAOUPFhSTyxcPZsP7+E+4oQDnHLxfU58oVnR1nRBd7jhSHrkaodSE8E5J7
WpNZjjvcU1WQLkyot+kg0fb7F9EfUgorHXf8vcXDqGgBNpN83LUNdl1Z9/hSDd7SvyYzXrVAV6m3
+GkGQ8uxujmjcxmiLPhGAuzY7H1QKmX1dMYgdGfQCbp/a5pBaD/VqtwRlAVzMQ2LlHV4ENRvo2I2
bdwYJFD8OFpF4afb8rS+1eByd5hS4T9EC8t5fcKoGBgoHWq30jUuMLS83KMNY5BcMya2Fcq60F+I
ghS4IkfTmgNtCitQEdhpIYjQ1K0C4p5Fb+Y6X2XWPFuti8UIBdLCSLE2QEFI6qAdGN+QV6UV7JGG
7bHL4ARMAscDATh/VmbVuo8KxQQL25bezpAJ2F2Ic11lEKk+AqTkB2WSnbJyOtxT+zsSy1Xnz3Uq
rKoZj0veOHCRjjM8bB22F09uGnl/e0/EmpvxVN0C0X5eGVTwsLS1Z7H6IJFfZwVgmJckJ+Wyr592
1bo3JUrT4jkE9XeK/xxvGIp+NdydgRAUoK7qCTnAC2/LGKn2oAEDWK44cNU1sV7yQvFXaxmepjEq
ARElHMSKu4MSQm9TJn7OafWAoCwb6VdBOSSh11JkIR3U5RFfRiP5WtWr02zaHvn5UMbm+apl9dWW
JgzmTyw3Twcm6WirFa3+bIr0ev2h31oJOId4TOtCeTs3zm83zPFAyDKvSj3yQDq+vAEozfwunnso
NcErIB9Oqi5GZYYL2Qt9gvpIHcPUJVxuj5MG6rz5WKUGLxo5KAWR2GjdT2tVl1TGYGZWr7GgXMBK
FGSPQkE5BqxVQRqXU3e3m5bkyjtocgduJ7v9VSNgaHkSqW63fpTHGU4n+M4LgXo1WBkk2Y/GkxnL
jCg5R3hdApkAI1teq8tSAlj0sX25V5np32lSPK9GKF9k7s9+kMJawi001/esfwIsA5WJ/N9aEQgi
5PMRbwteiyHVxzF7tkdtz8FSDRIK76bpQ5HBTM42teUIYZtXdA80vFi3DvvfNGWc1lI5YIikgw/b
HtPvY0FKwtZm7nDzyR3YWUEuIdy1yB3xaBCUcgByJyqySBrGW8cMR6khWvm0EdDywtRatYLDprdJ
DrOhX8/i3wU4K2Y424lx94N2MGREM+O3j6dptVUHSYQ0GIyIzFv8QSJ3DwFWyPiCesFJbbMzEI62
gckb8LLh33GcQwYQNXzd8c05C1i8NBeNKu9I8sJ+WsBjaEtYaXPluyoNZaKI1GZueCNVRfN/FMDO
+iO4iz63D18lKxBTEv4DTCz5L8X/j7KK/pvlywSuew1sU45tlc6Vd01hzA0Ht4ID/imXuS4zhZiq
ZUiBvdLJMozcfeGSYVvvXUoz4LStaVj65qw93K5SmBYNYASbZS14ph+OeQdpuHdUSy8jOfqfpyXb
YUZLwK7D5wE5PxT5U++BOcGkNIZv7BuxWumQQAgj3ZeDJ2lGluaI0IVovCDAis26KVx0s+zT8KEA
OObCzUdXbzrvmJbDyRYJ4G+mFWA3Adx9VtY62vKpD4FtZxPO/0IPZTY8W3ikK5SOIt7ZsVDQzM2W
GEKlVtQN6MAx3fYKrDiv1RA98zL7+yZ/qkU2LTM8pR51fXtBiorVUjf1PIkBJ+0wfagdY1aDk6HO
Zpl9YvoLjJ27FwgEKb/Jtznj7pq6mnyLvMCIlaK6QhqJu+Bx9+rFHmZox1n8jCQ4Tr21U57LAuKz
qcbUDgeqL7fsXj9vDjnhrzdJDhtCwdLvzs2YtMn43aE3/fvlLLxppVaE3llz2vs2MxieuDZqwQiW
Ea3OWLNKk5ObpqdeSO/mMlLzwg1706GKJ+cw3ugigDvKJEEKo4/5aqABCZptdr8pMKDvysnyc7Rc
+lzY4Pz//ubdKU1MogP+1bpjaM+Q+RE6Qq1+swDhfQ3zzWoTGZMPLHVlbjiPRQ1YKzW2SypB1n4E
iaGZ3TOfrjawUh4E/voJEv34qGr4GqBzihyifRSQ09MVsANs/NWHuLbI1gL9eIScm8Cb4FswAJ+3
egUWaSET18/0vcclOQ/z0optLQtHovzkXI88qpJxbYzuV0mDM9fg1EEmx/ABMsmWv5GzZuTYk9MW
saRyMqmr9SEgYdCf1vVeDH/0CmedvZYmpOEL48T9H/Bd1DzAeR2QNm73vTklJK6aWLsatqp7i/gn
bmrOFpS/x8/3Q62OtgME0Tqxq7rVyJUwSqFIs2jOmIvBrV/VJmUiOzkpzNEJexEnQC9N+yxBx9YT
W8aNOVoejIazlrc9BpqCtCY7l+WNzexjbWlrBd13ZYA35+GgqHhG8S0xxzcpZ/qifQ2nVQntkkif
PqqnXl9HwLE1u21iG6qY30ebqPJ9NghyPzz0H9KeiA+3l23WatC48V2/AafezrmQ+V0l1kIVxWy4
qB5WeAxgLgMsbQv/mm7m/Wz5qMFn9JfIfPJej8TYodxJ5p6IX0xtQL/PkZGGiM/E2As9ifWHP6/u
/G1sxikxJionkeO9gY5ULqfK6v0nqtntLYCswNmlv/SnOLKtOcYOFo75hJz84xjU+nxO5f0mlThI
/4BktT8IyWiyAcfUqdGNk0qin9kACKNhdtFvEpasuM2vekLo2br1UPtNmdZ193nIFEuOu39XHMZd
xv4J9DB3G/mQs3KuUS/DJw2B9AK9HAY7XUiLjnFcNtRj3L5W2ZxMEetr8VAJwHFEC7+GmMZjbNOf
v4gixkWwB+qP8RAX9PP8luAdraZuvoecS5w4eoPV9rHfegqdxrjN0SnH5u/F9aqvz+QaqLaWBlql
Jd3BPHGAlS4P4RlbGoUmRVzdQwCTZFenRSS1XuhGAqW1C1KkDusqrBsSxhBRwDYtNl5x+SQdL6n4
vuOIBlQ+zT19tozCRLVrijfn6CPpATym+DioWEeA+8ZvKv6Rp9/ekpAB51Adc2YGC3OAQGBZL2wS
9Am6jbsToT3j0wVdOLjxNemO3sjU7jsQXxg9y7mwS51zM402LVaHmax4Hkld7YsjyTecJujCNzRn
FDKwWajxzaw+SnTo4lfrrZwGNO2fmGbHcaGZxwBSg3Fcd5ok6kVpwSfPKmUbhBpd1yJfbpvf/hPG
tBY97l/7zvM0H1x8xeNCw6EsyIIgc/2xHVtwDG5d7Eh7Femapp5WoaD/nd9Xx068yyRQzXbEUE6O
qN5BJfodoAZ7OGz5mXq32vROr9WlAy5wa9OOP5bSD0/enlUSI2kshMw+k+zasvBKaYWO6cV4WSUL
fg8iy5FP5rUsWuPokaIW/CO5b0kvDSTwRpFDwTIx/ze38TejeAsGW6dqg1YDgrQpQCEMhloPDMDJ
e7lQ+8PIKdO0G5w5tW3XXQ4uVRig2M/RL+oBGVMClo4KejXvC38AEsWjhzqLGI8J/XyUanhIEya3
937OY33oE8Hf45C9vRkSOPaGaVO2gUryVmUJ+6GbuvISE9dSDuXNWfBkDyUqV5hZD7nciLOOuJP+
jcOVB2l8cTkCyB2MVXC4dneA1/0NKzifphxxc7rA1h+YNR2KEO0XJD9XZKg5q6g3v+GGfVTh9xQW
kEByv5aDkQIXCdhnix3Khsso5YAUcEDgoD65VPkhHLQuDlE8AItmhZwW6a0dPdkO/OwAVL3Hulx5
6u/faa1W/om7WAq3/7AytCJzx7PFoFWf6/MawPJHsaEpqdNUK3uHWFMuwgCVOzNdDwdI8ILNa7Tl
22drIOhV9GaXXntK8em3D07PuHw/myt9QrwYjuI+kXifq9Sn7fgW+PeViAoOHKMqwHMrGKrTvXEG
sNuFajAIHWoIOvpLGr45bc+kL/AU/4djlzsa0Cj1OPubld4Gn05y88M65PkQoNHX6ze0MQF+u1mc
YHL86uX1ElUQvK6h4Fd2iy5aQlgHzmt4A+dYKFBpfdrrE91Y6xCFcrdapEqlgqeVlIJgN5yt/I+1
WGPcGjOf7Bvh72ns19gjXVuggwNcF0BH4kDl733ESiDPBquTeW2iY6gjK5f69vqVtLtl4fpJxNbO
0amBzFYv3PnTPzaxW/AnjYshb8n1RQdeSpW7LNmHWSfqigw2d1KtGhkZU2ocCwArZsyk/hp6zSA4
CzrEkp27dCAhLGnxK8UQeCElDMjbsF6TR7Gj1iwtuMUVzimqliw2WPATyP4tHKLR+ySAF80cq13f
/dWpw7DouVZ2Y04bMUeE5kXHKmeLGudt8LL/syXU2sRgA/WqTG7wQg7i1WMTyJ8MyJybfB8i5qP3
K3ugwqyHtlO+UFfGXQFEwhetIhqrE6K/Y6pybcH5tpdiBgPteZBCMgR1Iu9wnntDnER/fNFM71bO
bJMLovgmmx/0k9CrObiASDfRk1avvA2wyyH1+B3T67kNmRxgCSRQ9evmQ0Kia7dEwpDa48/O5zJA
yRpaa4iNashmw7kbRN+jeMayxZphHqA5/VN7HukeTeGDeSxFpyTbvRljjrqaokwhFNdNcY9G2pQT
t+qA/JkQ65ir2kRVn1f3SylxQU16Is/5Qwg28IpJ1me9tRPQWbHcAmbsHgHmAi8moPwXVeDlXpHc
kms6On8w7NwTW9PKs0bIrV0ATS1n7ueFO1Sw2huGz9e0zTxvxaVBBj7lKPgGKFT4E6RcEjc1p0qd
2kDmJpWG5jn//M78Je4wCMuewN7yl6uShplFKCP1ZVy+4bDatqMyA3bWxlXprM08iRw0I2MWRxdW
5DnnJnTj5+Mippq7xeSonNp3JW4NAXKfrjKyskxxIMH2c51LBOqQMq0qLHkaDRuDW8MaXetbMdn/
sdEVjTrObGW2Bl9z6Zz3utuC97vT5NqDbvIzx0qdy92zqQjfqtwXypfNisnkL3Fb0saYXZ17AK27
V+wcDIujEucoRG2OpimeuYpwGO9WGY0C2qKSQdfZagp92PuHiVKeB/zfV7CFDj7nrVbjoLfWlp/Y
hucVj2RCu5UrEVIPJ95VC2I5oCsERbtdryk3Tb4jxlee/WSJB7u7lxpGStbYXPWnNbDoasV4Qqzh
pwzUr/jRdw5LRmYJ1EwMBiDkUJ2bDD2Zqe3U+Ns4xtOJYg0Fiv2MMzhtg6PCp6OBggwfaovCefvZ
ow2EuwpCPokDPe+FURLylmSkvMnTGTLwXnIS0re2bUSb0qysKH52YZ5ASfor/fE/AHliXgH0Cu+E
wGoxXI4MgB9tabDh0zVUjeFQu1Eg8HPCoBQaMUCWyQiaIC8FzZahOOvGZHhqoUMQyo7g+vDmtL2I
CRmnspac/xSDJJhKTkce3gMaTVwSEpDheCBO4KV0S0mbnwATTAZrGV6c6lXWZwNeqW5pVgOmF7vP
fOPOSNp3EhsDdcrdbBP7L+pEHWQt8NO4ValC2YdJEwHB1uUIokjXHswFtsPsV+Yqfw6AOJJ/8RZf
uJnTk1OOiudH7zoOX6+ImaoKx4M8LHUU7wNz7VDQyj3No85YAAyA26lhczfUd5TdFWyHAWeLhFiE
Aofgy/wT/Ih0lp2ucBpyY2n6rAXApVlLz7JTbVQURxp0jL6z1cgnVSACEGi3Seu/+rA28gXzUO3g
qF5tNNc2ey4mom7i+UcbYnYXSfVgMmzCO1I+avOdCP+6ZHCi3u2Z5yce4G3OpGssY47jiS6SjaNa
U7NleNdbMO9luLWKQUNl8atAtDSQLoOoQsaS8GJ9Jo0YLznA80ikaiD7ISfWJqBZX6wZGf5YcKjN
UZQW++0HPDXLCCu3DYFzAvvnJhWv2biI7ZQjYNnAjYdHQiHE5Q6xzfI5VKBihXJ/p2gKUD/YXj0B
yv95AAl6evR+t9jy0cDwMiFAYsTpJ3CotMUB/lqIu7EIMnAGfP2oJP2EyCkmVx9WYtyeXvNJG2bW
wSsqCiSdZ5bcSigcWPaxORiHJYpKmx33LvXilrsVEKlTR37ShqR/Dp/jV6NuVSnyua3O6IuaW+yJ
XPsEfXc7AdsZBcCLRvwX/qwhvow9E6nAqMH2VE+dypmX+pgF6qah9o/BCuFfdTp6ZcUoAyN3cAvz
clCGTq9fDJtYIRsGJm3A8saUrwYE+lszp+Imze3hJES/ZKz8yr6WPNRyCApYU+Nce//EZjvZ5zAZ
FN2DmWg4Ny0JKQLUjhgBYD95NxJ3DaenzNmokfDbbLWi9mV0BKTkT4QGge59LrtrYHef8V0UtxDl
bRecULvF1Dw8t6Y2n/rvh3uCzgSyfQ0pDCwQ9tPFhwAu7TaMlW3ePoSJ8xuLCvqpJDQWmgotYjN2
wXYEpvQVOjCgsJUsiYaMIJj/LrD4750IFnYMJdDpkmAgpg3hNem1BU+UvDg1Cl49V4dC9vknG7yj
Bcl8bCEXHEtsgUgHPAAAlDtWajKlPh0O63R8C0npb6yjrCgwUaZX6VnXTqBm6G472zlVppvxMROC
yUu5rSPrveLbLgQm8iCs3kWGuHVRpoHyABLoo8+P1MKz0LLhBZT+s3eT3hv1EGqp3NtSkE/NLnCw
9H6LDIDHu1mFHk491B/TTJU9XdysU7a3IsE3b8f6DWRfsOBb1WYvV/s1PPuM3LQIkjOuETmfYUsH
seMkVHo/R/aAP/8f969q/9nLUG5uPwt6onvjzxvutRyncEbC9GTEBbAJvlgXo5tHT1JH3GqAU2XU
jnvbOqhbZ2ryi9KpF7xyFbmIG4xfIjkLL7nI3Zig9RIcgSCj0MYq/sHMKfTzmQfnLS2su2Lu4A8q
l35kgXrpPRqWt1/kT4KGF9N1eMjgWQRTQBSPXQxtxElDg1MZeU1Xy92F6dAJoQeldWW3T5jKXBMX
PknhiG98TC0/qHTgHDl/SImoQwCc66x83eh1AmOxT+goHnPDbb7UBzTkvEVjX/Ky8WOTxpFQPe38
7os5bpdyXuZCqoY+a0hj5Fd8nHEy1/+PXrbrnkt0O2iRzejnEtTiyaAuXotmxv70B3SFc30pf9H/
tBIqnj7VVp2vcJgDxrCWA/Hv84/qV/bGIDb3bVOhFuhtcK9TIIJpfwOp2A5jq4rm6ZmRPKWKObxX
Cwv8QRy6IWpoOiI/mzN/cdcEUJiRFF7lbCX24jvYCOBT0X7ecd2tSssCDuDmoSt8gwp5i5YUSBax
HL+C/Wmys7mpjJ00kuQkmwvthQQXc21FjGN1RZIYu+z3v15/Ta4GfQKLiJIpga7k/IATw0UVDz1X
NxWF+p2JRJgpQVWdm/WiPJdWeoDp/jq9ag5fk5aH7trIO80c/zGYmT38YVqiFkkmN4i/LwtVZxze
T9XsVX7wKFLY8ogtDdz0ci8SDPyKCxt+OOLedVJkEHmWMTx/y8zrLr1fSiJjkB/PYzhpeHQyRWBY
2AEgGD+YCxMG3ndeBH6jR7h934sly9scYxji7Z5haMUe+VqpuAtgtKG6toguxDu89hUkWrJ6V3SF
33ySd58QzhkE3WFy1XOAjzrqubEmscGuTwmDkrn47zriLI6OjZhZJTNUGgotpByuTMsPZt/4lXck
HfayEEWPAuSj/F7rCUi78AuWUN5hyrq9QXDIRqf26E+Sm78n5JsC92SSi136t1uhudFbMXp8OzWn
MA9x1GWlBTxp9/ZnOjrcLFYU+o9yPzRO9qNeFEuh4wrFSaZ88J0MGGZyeWGiC/bu4RP1e3LC2BXT
TbuYahdSjeExErl5yDhZay+QmXaoMKWrhb0NTe3lw+RdOiguuVaDrjoasuII1Wo9X3eGLiX6cEz4
Pwe/djqWa8vMIBPC16pRhEivXBxVH9PK3DAL3vkHAD63EFhCGXZIqg4K0j+JILTaBJJmIFan/f4n
KIiwFvGBS9+enT5MSVcD/Gf+LrxDPLwim2q7PnM4a+h5djGWqKZmQEoaGy7sNn177yNoBb6E/5vm
c39953WxYbXZTuuWnwT9oHb0pTeXI+BIMCGX6NrnsDZGVWzCmdFfm8GdDlhWZa3+KCR3sUwDng7z
LCRMzOAriKv9AAzkXEyY44Kpfq6UTohptYVZdV18mVHMSGIxQYnzEwmmw1kzOTvnzibg3MxKKrOO
2PTzr8TEpDSGAbDXlOkedGGiT8UPcToxoQOs22eUvDrcCghdKojNrTFNSdqXrEV/d//3674aYRg6
zaG2jf7Mawj4FwT5DlgU0gUy2o1Is4+u0iT/ZCtfCOhfzI1QXjYq0wAUFo9UGVVk8RR9RFpIT+15
H4YMP2ed8MS2RJwI9yqi5XaVHNweBLwDzwN5pMHMT8qZGrvmvq1XycswWfIaHB4JDfw2mJ5PUPMB
bwMA7u4a7fABfCdDLWtywKrxuy42Dtn70wSnbx9n2WETEtCzyGgaCm84y6C4a5GMa0L5pOeewxWT
AQ6fHsHyVFagXdAoNjL9oIcyQ/JapyBaNiLooMB9BntIONLa8vmi2cZE+5x3L6MCZ5j1ungEgNhV
xMA6clszYDW/gZ1M4L4+2DLA2XqupmvLJvPqChIclKlBe/fJbeKgFLKOvx6t9zWoRzwfTgKBPstA
RpVLxNTl5U5T737fGy0l1bmEYbs7rp8bmXBnvmJQIhTe/c9gPrBAgksXY1WwpqG2L6kyXGQ2JhYu
gsb3WmLDceKbydfXLR8Dbv72gvmJnaVVnSgH+pNFpBosWUnluctznbmMN8oLOp1xkB+LNMUkr1XT
iLNRHmACovTczhG75weed10RuPz0MF7CKST3DbLI1MUucvGRB0EvtjXpRDzO4pFlS2uaGYrBq7Ce
29MMWGOfnyObPmtG9Q908ai5DZGgICgEv0oQMvZnOertRiQ4pSV8WjmQr18CIiiBTCou8iIoc+Qn
XpzDea2v2LZ6XKkbnuvHh5db/XfEuwTBrhWAJBsBaHxeevyUPVwPjcJdidQYzVLPqqdP+oJ5mUm8
ntum5BiEK0ZdZRfNwsexErN4OnkdHVzTtt8FHe2rBVoVRxipWsN5ZThMwf++GtsNOeO0QhRPNpSF
d+s4aw/maHwJUTZUt6+HBrzR51oATvoOBP8DXCAwZBWE+fM8wOod3thKdqWKidS7YLlqk1fGgal+
FAaPdosr075TODjbIxLQ+9F2A+noW+XwZvfTh79NzbdQv+XiFnZ6hNuKjWaDWfZfstTRKczR4CNd
lAUlRvOU4c0VEMnGn1Vd1aCGRdDPXnyMU5NiBe6XznMVvvKyYSYN4tINo9+8K3EErPHKZqUY3L3j
1lZRjk/8hjtknPFnhUWKvcgxyRgtSFCzQfFRR83qGMRA9edBaKYZlWoCenoNXfRsrFxOCLdU+pat
x3jPxpHYSTHT/qEbI/V8WS7XnBRAwcYyavo1jyciZyYxC5yaRT4iwzVBQPdJ4Ezg/JFv1m1++cRN
j6cYJuv1UbGCS9Y1utiYP4nsm3RkSZ7IDpeiVjfTuXWelLIBwGd+pB4SNRiqFbJq2xcsNIUfdATG
qFetBKHikXu3e2Z06eAasq4rjEQeEW2jhzWNjLpSx4etC4FK1vJ9ldPMeVKp+pKBncgf2KRPGIO5
jFa6M+fa5DfiM+4MczT4MKPtUjDJMIHQ2Qc0S+6CPsa5hwRasOxoVAndI7FRqi7g5jKb4+0280zp
PcP5vO4Fuj4DpAaFi6fW6BIxiebF7i1bmi8fU5rYd2SFwO+LoHi78e7vWE+/V5sZm9OLn/i81RzF
KpANMgXhxfBbn1GBYdNMhZLIfcsn6RZ+66HfAKtPlKXM+5pKdSG2VPn2mS624q9fRRRK8WE9Yrfu
xoXz64wyPjLxqBf013DPx3o19B1ixywZWscfTAkgNAFWcEPJqph/c0DT7scy4edbZ3tNdlHviXUN
2BPe9J9VvBBMoIjWPa3nxCsp7FA2miP4O4J3DrgR8aAxd5JG/PwZebasrIoHv1MOnKsekDKBYZpU
AIz/XVCjmV1vEK2azrVDYaJ/85nQcVyVkVJxNWBOs1lVX9U35UD4TYkIacVAOHBZa4PHn9YVs9Oy
+QMsbwL4+IytbUDoj/Ytpuate8y+vHA7wEkFlpUZCnm+kwST9ImGbC21nE9lGYw2Zrnedb6QBc19
Y8DdxIPDJbIeafcH+lmySzhatnR78RTj377l6FG/RmOXxUAp5OAzkE6FGtSCsSl4EZU46T6rXBsb
uQz2J8yansjXohSlEkCCayQoNNGmET/8zwL07pulfRPxcwG29AijToYGUL9oiEWFlOywnoX4w0e+
0gJ/ItpQFFV3Pzgi3mf1P5l8ndd0xP1DARWG7IFMs1/bWaA1AgMJEVIAFbiK6illG1N5QHo/VPhG
tImxqFNFVkN0eRzQ7WaDJ6tXd3/5BoYtZv0u0pncSeGnRi8REqJYYojC2NM2Cdypzu/MHalRtyqn
CQ/1Nd3LWHQdbw1nn1Ve+RZt/Zem5tm7B+5iUibLy7zb6Cqtb5ZKi9KasCZPhE6aFBWd/ly0VGwL
VlFdlhlwLFgx0pOgMg+WBAk8SszI1YW+RvfG+JARw19oyEwZ83ZHL4ThAPR8KQHNekyTcoQrEB3j
GCrkuhUd9ig1eDEZ1hd3wdWyPQtUMG0GDWPHjuDkEYeh9yrJ28IueyEDGsOzct034vnRzbOzUN1G
kZchP7XeCYaYAHlxRJW3fyMoc9+T+mp59I2A0E6nliLGkcdGe+25FECjpVVC8x2chkZIWJhsyQSt
4gFPzlsjz6BQOSldNpDf9ca26yw1GCuzwPDHm2sIcqjBbq9PFkJrNRBvr37kd0VHtSBRPiBCe98S
4bbPOCrHaKdF+Te021Ehiblg9XgjUuep3KW9OVRE6pnTJjTyOExbhui+yIdTuwqjdLaIviWGjN/p
CExJgtR+fqMpoKbKX41n6igz/o1rcpvcEiTtu1kXzqP4KLKCmiutFvFqismeaNPdJUibyK/dwUqX
HxSVWjLSjCtkdH1sZ1NoxdMnu5PubuIeGchImhROctUqn2F7Ac7XSb3zP6g0oSaK7Z1a5Mybkgeb
5ZfnubdNZ0Ymj7aCWfv4G5hJHKGP/xjdbC9uREg09Td1nsrYwto1G33Km4ZdT8kOOWbB7AGCl3Ov
kZdY4K7JIuHMIavDDJGvcl95JITyTSrDKq8po5e+pHz7zJjTe+pk2DgUvPI5sIoK0GmFsEqqzRzk
3TDKYlTFZlFPfjIdUeOTjeA+Y7tuh74fATnSc2VDCAuV1Aw7AdVRFwNBIEVM2CkEZGkZbrLOSL2d
f4eVj8fEPzUqL5XCkmcKSLrHPwpEh4x+qb3puYTq4Op/ufbU/9nBytesgEP0YO5Rj3b8xtXAZtUs
x42J3ISuScWE/XGJ0TRYsEDn4MHnMzbTn5F/vZYdFQuGUsGEUcjpBNEOhXs5XZ3wpWISQk4I0pKy
T6JZkTRZdu1dVCDoazSfX0B8pY2Y/shSfszU4d2dASrF+sDuGAY51JaYf8oLs7oEvO/ShN84uLBz
2wt/mKHhGDGQAq6sqdDLUeEfwjrsnzuQo7ILOQi7FBJ0TOJv8V4YUNbOXo1Mwcfc2vCxOAX73/hf
cj1olgciegAB0Be20K8LsJNCs7jb58e/V/b1ykSigcmxjxwqoSgd9D/ZYOlEhbkXMqRRpvDdE5sl
DozX5xII0eqZiNuCrvEpRdzoD+SkRMYc/rEwMWViibLd7CzciKsPRRq1dJWRCRSfolSwzP/P6fiN
E4660Gube709ZEFdlzVtDnGqQZ/Xp3X4BiT6VApmqjdkK4xJK+6nObi+bJVsVv2mveYNi7r6mLIW
nyvKcie8i/F0DPNFQt4GctuafklmfQ/0/gr5kBkNnVTZHaDlIamYwhSCvJ5IrM8vMLRnV84WOYn1
5PHeO0CciItJALfE4jyIvcUUM7hylu27ppy0F7qPluL4ceJ3cEI9xdChMkMhrox2Wb1q+TzAuLCm
fVhHnGmHVsKKfzhmKVAf8CQ0let+L2FuQvbgQaeHpyabyGo640qMYuJBp3RRvjdtub0XAPc4EdbL
uLBhqnx4kCJ/aMwz7rFOs8frONc7rsI8qtslwIo8ydiiYTWhRLGCAzIMaTbSXxBnJxfJnkP4xx2m
ycAved3wbB8ROHlAnCwiMu+q8i+5RX3lHLsv95cHHddASfLMiSZ33Uogq18rdJwegDzGM+ds4pwb
UMe4ahok8T+qy6YZzNx6fwgPhpo2HPRiNZBwVVFV72JqhgmCY1Qzil48S6zALTBPWjSzPlRXdZTy
5i0kBPNjq/8g4eio9+W0Or1MtTYRltgKZJf0xT6NmrvrjnxmipFGXZ7OaR185unYpep7Rvl+JT0/
EEJbmZiZ/XR8Nbd/FnBYkcCLUynNmMljo5O7Bp5e3V1Q0FUGUcFtuU9C7DBfkRDLVdBM8akivwuT
cO1H5tTXARP59QbZfuFTR7nZEJuzUZLzVIoVZO2d2a69NnmoEQIbZy1GufU0U10/rIknn7os86CR
NQDgKaTzCAjDZJVHe0DWUydns0+qLPSQmoGD3UDSxW+3vkhSh0+OUOPVBGt0h1sDmcZiUG+KGazW
a1Yr23AcQOQOHuaFDG138voTUZtWYOEDof+65bFtrQ/HXh7bDMpguczOW0VsBp8ypvg8M4NhwiK/
WUaw6PH3LYaN/wdV4MmQ5prITXseAhiyMb3rItSmHykWChwkquikRLc1psW4krrgaY4FKtpW65lh
2aUcWXkLuB+Qp1ioSgOKLbYdaPRFVXy3XMKLO3W6buSBg2jA2l8UDET6EOVqndTNgsSOEFcuy79y
kW0UK4MwUSJ5ny5ZX5038ngTdS0PeogEHMct5Xj86TNBqBUd/Nr2kHAAZ91f7+3jifvdYmdKJIWA
21/oCYi2QTAT4hZkaI7njbCvcC9TZJehD/GIflqq4dbzqGvcD9gG2u1DsCdHsDz+2sYAv2KA7B9w
piAqmg2h1HrvnN2jDYKBjmjVp1/hfglrc1xyD+RQh6mwhpXdNmu3rcnS7CxUmzJ5K3IiZAXrZLx9
As0uWw9N5Lh0j2OTmAKcLdMFx1owZlmSjZ7MGpv7i5sCQA4DDYklpkqIcq77B6sxoPIgAbIZLmkN
4A6YqGaGH2bpP3swazxkf6HXdtkgFjEvgdkO5mfcTAwKpsUo4uDydJCGM8rHcF2K/HG1bGOE1Xfq
+XrMlgdxjkk9WZ7usiui4FJkUoJWue2feHorB5oEqJm+m2bqwbz6IrgmMACUKgdFfNt6Lx0TzqJp
zVxxinWyWkVWpJbUydvBhr0nUOtzeQAK3DEjY39ubuCmdSCpZ4d+OCKAx+9h+jun+Yow/qAGIxxQ
u4XBtbC/knd0Oi9wE2H4lrpj28qAevIfVu+nw4GdnoMm2HC3WNgH1zpXsFGpieVVyrPQ0oWVoEyJ
hMXvS/j6cmTWxqDFn4/Uoq3vE1+2NmzzmACAuWavhjstC+P8ozkv0YC8WLbvxq+d3IQoQA0mNPNI
PxurSzD91JUkqdvjo8EWfiNGYx3nBRQQSm+kF/jZ65JJZdJbZRP+Nwg2q/8Bu7VHqTosdzzvWqtG
tQD8GPCWCLaANp5hJG+TfIqAdmdr/oR+ejUnZBEKY/9xhAy3DsxB0p0pGS6GMbtx2ggaapO0H6MR
bjUEhiI0y3M5uPx7spaRiGqVwyrRXjFBSp328BBB70e8vh87Ov01RtzI/fkPnTmxRrsUZLj1GhuK
igw8cCh/AAIUKO//65NOqO0+dMpiiO2T7/0e1beDCH2zh3hEGDBS2TeaBPaK4pgPld5AzFIip15d
qNBxfFC8ICgkOPtr17YuDf6hwFjYksmCM8ew71Ki46WrnTOUhaNYJuHoWeRN4fw98kIM8BxJSUVH
RuFc9Lrl6lmhJ78v25IRQ8oRoiOE8VwDFdJai54Yhxv+yhtvglCTTclS0uJBM5h8rhtCjHKFWbfg
/VX158qks0WZSsQIy78jCl6bR7TcWlXpHgaSEHmvQI4D87NPS+cWE0Ax9XXNWS/xMWbizneLQQHK
M/m0S2sh/exYgj2qvNNM2cYDIx+vV0u0Tg2AMywuHrA82qfqYk26csfv1Hll/CS/ggp7IOVrK0wy
tqi1Z+eE8NB13hR0WuMrIKFWn6YF58A+5cUgs8pSMEbyccvWk2mECrlJtgJjWGtlY62M7uwXguEK
YiLolRkvH60SuQ469/1iqt6qn6kcILCo1IyaAx48Yy1iQEi7sXWJytHSXCK7X/Kui92cV5TjV3RL
0yWTB/CxKI3dH1cyaic6vkxy53wW76o0Q6R1v4bfDQnJHcbhWTo9Z4GUTDL1gvU9WaVxJm5gCdPJ
IquW2+BePj6DrZwIzuTJAdV9Xc6C9yHrQ5dC75rC7pVAWidiD7aOT+ooQa79UAOQFEVfHW074Ese
4axJRj1OZ27vG5r/zTWAmfTMlc/pCOhTVQreJJQoUtVduKN7ookB0nG9OlNbgxS96qyAVeZBMNMR
v4UvkaZoG+lbdNDbqHyXGMEd8kAUZw5S5dnKBRc93GMAt6ut4y/BwHdxJf7uKqgNh7KBkk46WF4C
hQ+k7684hpyMc2j2xMC/MbSmbr1GrqgyWEDNpz78r/GxsTT6bzR23DAI4JC8+lk8HekECwuqN0LW
lTFf3pd+PVCCRvRAdxUgBsfYpt2A1A1quIqQlqrhU8z72vZPj1E2Mxh531F7WkkhWLIpa9wH87tb
L70dbqSOLt26PBtWJbxc0TYC4Rixgm8gFEXsOMglud+TeE5rDmmG8raQk/Q4nD9+8n9xaxwsEb7f
rTak1sOZSClAt+Ti0jKdK8OWhMygN0zLLFQwCO0UMCUQvH6Dfg/5BRBSUgXas5sdG7PxuasYCuBs
NLmJG0Hyi6pro6Hv91QRSV/kLKB5jV1cxSNdbyS+NfX+lahDbh+ZiPwZdrHXBj/HgUZ7UtU6Jc+n
Mu4NriJ+l4UHeONRo9M8vbR3+na/hLLlMLLsRHOKSk94k0C85M+Xf/vCo0Lxyp76L3QRKBajBbjM
GhYVjvWzwj8w63JMP14/dcuczKT9nWh45UG6geANsBuI0nuWoDGtnB0Ye1kdJms24cizxxltBlZR
r2IWr4n345BP3h1COCLofq0XWtdICMJQmkFsUxSTQz3BA2H28hyCdyQoaBoxna3xeOks/CveM0HQ
iW7G8s/+G2LbKGqZbKdHc5MY2lRaLMwyNV194h0GYhfO97sk2rOmJdorVczmIT4J44nthSGf2Ap1
BdZQ7qo5GGLpdIv4BZZttk3lFqc3T+gUGoswEkv4jn6ldQo87cDxkD45nNyGsTTNwHouw3dPSZiC
sugyspsekRqYRAecd9AL1F5a75sbBMEsmMRSVyvpBmovSorOU5kMJ7xzASQqisvj+w53FG1w9T3u
s552HUKyz+T4k/dtsTIWz3tWZGqkxaSWuXEPdfm9D3Qx81ZCpssn6q8uXnbb1gRpayQiC3fT53Bf
25wr1FqhraX+WPhK9lnr91FhD0eNETeEfwEC0jzSqbDEMPVdjI7uY4f+XXcJO+fvemUvZ5hYW0oq
ulLIh06ToQKzbo/w912ESdlDDRKq+but4aqHRT9mPS9YK2adJ/mYc37F/pO11e6p7p7LmuvY9bul
Jgx8lryNRYE76T5GKEXYNlhWB7T6TxuU1EqQufOqzjKpsnbMg+/TwMAI5yDuGeG0NqDEjHmfLLWy
7OpxsWJrvA7pcT9BrwcDgCH9Sl3lTVWc5dOcEvN8OhggCKIaYlK7UJQsuztPgHWzdMSQsIn1sd5G
P4BFz5bWLEWzG91ogcuJiwlch5rErREfkCvEMc4Q8Zv8H0eP4xkJNszclvK3fK8cvqPEZVwfPmeI
JnKEjBqTzxmBDwt/DUDT4cyeAMuimcB6902TuxLlOnD+5bBv/86z5yW/qZX2Z4MPDQ6V2XqY0fAx
HmgGEjvOEpR6Arx3qZ8coJS9EExB5lSPDxcbUPQZwaftPClFfHZFHGHuk2HE7gdUnJfZ2PNleV7p
/19iDa01sk2nVipC3r28Hw/E0uynfa3fd/i//lfdywNSWxstCCuw7MkhAtwS4VayIArN4b7EYYe7
o0Mk76w9Rmxfnk5Igitoz9AtPpiHE5IAKIIfYqnKELtGqdbStVlW9y9UAkAbPRoEnQR8HuTB8SMA
kCLGdehhVJAv6ZEF6Pri1d8y+vQidGydxgs9IvYcrc9H9kIsvd8fLS4gsXH6G25nCAjHtWtwkaPo
1kD6VP01G5CI0BYoxgD5DvnzM/RJtXFXk3a4zVoSpvHB+NsRGKlIyChav5hEPIT3o9KrFZ4j5yDZ
x3VuMPPesPl1PCB2viHOxYDf4fN+RlSGVvph+WX9fBuKfeAzQE2n5ocZwxBPe1pjNYHIoTK6J2c+
u4wOI1wBXz76sv8baI7ABGZfsmJ6W/c9c5JpRThu2A7vgW9YeyR6WU0nldjGCm7CHwT/YrjWfqSt
jTzX9pJd204OXYvrp9YL0OtHW3c5TBBDKP1naN2kS7WEz8cRBzdGR4Kp6G1a1rycTQXoOmAcmiDs
BSTaQs8Ev3QisV8moYtHUI+kS+sPaInjVsl4en/9Hg4R9wblA905o21S9NbP2bdSnUfiiC6XWSrL
0EJ3k+i+PS+tnVjSMWvoRAOP1Na8mJgDD0GHFhOrKV5DjZh84IAnlDmyfnseMZkkINb/6UKyJfdl
viG1t1CGr9PRbOX3Vt1yBEYWUuCBAeULxflHqWz6F61mij1JsrBLxY9KUvry+Wa0ExRRUOZFVPoG
HhmmGaR39H7tL1gI8JomNDvcA1/AofJoKbv0eFMcvc9j5QpZe268sMfhuTJIobZkGuNJjlDg+UCx
ZPH1ajiI8HOgwikiULNpmvzxAxewBItoo+F6ewhWJZy24dFtcL+H465udfrYnoOKV9cluhKqUKpI
hHcrAHgmVgb1i1wPwLsehasQ0xMxeFhhLSR1B1wT8I82k0Eckj3i5m3M616ml/b7xoNhHQgfcZVv
vhPjyVHGLr1HVIIzKkWytSzsKh+vJjpgbesBm7WATQaSdWdy7nrrovFLrGJU3wtAeAzdZFWxqrYh
iUtxNcNvQjE7p7AF0/vyEp8s3shnEw4Ruo6caTUvt/p6iFsfvRIaqxUN6J6lYWVP0ax5mfYy3xdk
6s0DLtcdAszwcp66W8z7KjV8z3YobHqvRaEzKYKiYtUhK/96ckVt/sR5QUBKjCGlln+a7ucKdel8
i0Voywot+tDeR9YDg3kzDDl3cXGqSzSmsA58fRgUxmrPUJBNWradlLNxw5eRW1g0AjXUAzWKT7ZQ
/3QYZjGnY2ZEcKEjem75/isERi7lLDKjquSot+D/9fUZAkhvy3IBRt7VkG2urjHftu0ceZARevxo
EAZFmUQAFUt+BJLcm9U6A6c/SKsKnTXtEgknnT5aAHWj3xjtNzgibY+IYFS/MoUNVejR6lwRndIP
O7mlbP1A2+QtK1OQzgZt2XDoTcm639E2bqZLarcMBhhNT47DGttG31ymBU5K2N5RTI8LfSqz8d73
uqax4oZRFHlUI8/dh2ffAiOdVsi3KRyVtYlP+j9AZwmfJNaCajYcYqWYCWYQ/8lHkEbehDCZ+4Hz
PVmZSsyj7BWn4oz69JvB89hzwjN+dHXG9aeYwn7yq8a7VK1NintJah3EeEFRrobr3U2a1VkzCrds
//emvnZy2BJDmc6p4uOLIV4Jka91/0Jv7fj7XX1Mkdur6y3yLLJuJTU5fxokJKE5GNqEfCX+u/9n
+ZvYQ3mBHQwC/KfxOfQUViS7Jo7dinkmlbnKdkABRDWnmKkCjsEPd6FlBEjaq2wuyBg/GUKnsHrM
CsiSMygmXVN6SeRLt2UbqHLcOgwYmv37Ed/5cEkpEEETLicLLVMMEJNjfRYssE4Zp026krmQsFLL
QaWYs4x1e58aI6fNVfNSSJFY8JBvbBiVo7HLaXt2guCLx052Pvd2bJ55VojY6WwH4ChVaStm+fUB
A/D7kVVX7fUQkblBgk1HxxFuQbWriSjY8VdRX2eS3296q39raoHVB4fYrg5M5T3gGSQmZX5iG7OI
bqR6LrfBUO+N1lcuaszCL5tG9f4+vnSe03i6SA/mT30Q5cCw8MZpYMLpgOV5whKnVj3F+1hhHYWo
s07gsowLCPLKKugpgVDL4hg6mstx6APPYLN+nyj9Ffxfz261UyhVj5U+iXIfNcLBJHEW/RTRgs9y
7Sr0a0KbUoRVP7EsGURj8hb+w0LZWh2qgz4NQrkRY2xepDz0itw97L6OqNtcSJKHH/lMESCUY0bH
YCTjhveG5Qj64ggn6SuygmQaILFvyXqTiVn0gFkcVoMMgnI04agX1mJwSW004OC5jUNaKRbFbqK6
v3AlIJgFFyhyEPPf3oPN2gbIyjn3CW43hBzn+ei+xSLiEqtNiZluSDp8wtEKydlT7aYs83MkZfUC
LZB1VN1hBh4cI+0SmhCY3df/aX05h6V/5ztMeDtA9Vg0unOacMjioB0H4EI9aAwOJyiWHtHKpjjx
hWdqM4sn0fXnwQs4SlxQciyKPyzXMjMVYFNli8nNQV5oYcMllUwqWKyFYiBIYTPjwpR/J6JcYFeR
XWO0gOn0/7hGwJ2tDv1PH7InnZ73yWHmXPGyu+G4b30Hbcuhy5xaP9WiROsN7HrlFCDLs2yHSGVP
7MDJj/kfFojX0RLovAOrQD3IOPT8TpNfppdvJM44l53T976o8P1ujtIAhiXg3H/Tn0M7/q8+2Zyt
PnQnPSXBlUcMQ4vyOGWmgE2VisQR4Blb/k0brhP9k2qteXjM9GxXU3pSxk8NatLRbXOAx2MD4GvO
teQPR2eY7HVxpJhT03znUzDm4spq35YSZsJepSlkz60TgxhxXuvdwGo7sXIHKX82rcThR6xJB+Ze
DOUF7ZdRmZajPzrzaqjM7NgVJnmQFmLCsLG4mM2+mlZ7CXLy0XmTJ5UQv8SY7MwEw2CY2VbOgtDt
2CH/0Lqv/MGlJ57oyz1I0BKfljvOA9uTTDH+hREewo3ylS09BB1V7H01072NMWKVgodUnxIyh0ND
BkDpJ56RaEe2YLHsKx9YhpE7p/YEbKCy6KuerpWTAQztE0OHlTaaU+yqoBRwI+95GnV9T3vdgxgP
Z+TC6yQgGd3FNFqUxDmEJfsgM1khJsYCyiqJZ9dDz70UfPL7ELNGzd33le+tZ7X4v0V3/0Hej84a
qoeASC2lqAx0GqYum87j7A4hiwVSlh+TzapmGWDvQZBzKQFNyXHMa0LJlPDPC/gf3oGojfKIR5OF
1KOtpMyPnRGm9x/dMNIVfoonz9yaJgA18sXJNw9tYXtTcrjmora/zGY9Vdncf5+h77fdyxNsCvnC
QsNvgQMASJl5VLnD7JkUsQ6OxflXC9ju7oe7/3nbpDaFxDn609r2A/292gv4m1pmXCwYUjKfUlrN
Dve/X5SRUA5xL7zIkgnTUkES6DfIIk7MKvrE0S2b3/nMG/o0hUysXsVB4IIBZZN+0NRgbJUaRn9h
zrUrpq3ZjcCmd2uZSXpQnVWRd9sK/Ki8p2XH1cOweMhMq3iARn/aYrB2NqVC3WRhpox+NC3GfttG
hTtjketQBbC7EBeUaYqGNzBHYR96Q/Svb5VIQ10eTIlPAQSmn8tCnvdm36Koefq9YL79OS+gpdF6
CiFWWS547pIpeslAoUKUdRWF6YUJwPWAMmC9sOBbfdUPS4gFNkLoSvZ5Usf7bZPBBcmnE3L7Ynii
kcVP6pgDrAEr/0BJffdNhskkgJdx/w+ukHw5/j+h5U8EWLqCkvTCQgdLBQnp26GOuEiSzOwjFZ5C
YKu9tgTaV5T1tNUO5wIVgnnO7/CMrPNDpxFLHHbifH0Sm2ypw3VzKHD+7Q9XA0PPvot8LUo/OV2F
3LPDMQOIbqA2KxjipgGkBjpIHq7kH1Nz3J+8zuD9AYTvHmlVkPYBEtnYUmz/Z3AMd/Yltz1+hZTb
zvJmm9uhZs94m6WzJXJ3+UCygIvseYpNN41cLWh4m6v9hJX/I3k3ex5M6lReWYni46MyuJFpeVv8
xIfj+E9bkB4KNUCwBrX4OmQrQCIqrEdz9RP2Ub4chWFPFow/z8qRRFIO8NrzWgxosk7lf/SwcHYq
dprwS/lHoy3xp9TIxYAPyDJDpbkCMbWzSnwdo38aBtdngJ73WdvB4cisZwU6kjVT84UTZEnBxyBx
gxk4rUwOwcVuXiuXf897/ZB5DbWV7ZCXl3QtaY0BqIYwOqyCSGT9eJAdKI1HwlQWNVMVwHgto2aN
7yjzp+XqpDOkzKyfSGaAsggXor2JfVJS34VirfGedE2SObW/qXt0Xfnh1+o13IdwqF2VwRbANJEm
r8Qje6fZufNo3yZqU9L4LlEnrbQGLG0gk+5bgQqCZWTB/dqZsF0L9ljrQA1uNNuuvD4vXl3FgqBo
AZbTt8sYtiy12P/9v7isKNjLn0HwpazCkyp6moPLzGvL9VqXDzYGrfWehOf4Msm8a0OB5j+KY5cU
/bx4YUrOoGqXWlqiEd7214StDiiKmi3lex/5eUygbb/l3z9k37mJHBPRNvG5Pboie9Ez6f5Anu0Z
2FfGPlDjShMP0HQLW89x7WdtnEaOa6Pc0hZQX6Bre9Ce0rHl/OuY7vUpTeSGqqbk/z06vmwMqBND
B9VyuWfkzO8lfyhUmCmM1Q8mkCAdswJg7017+WD/83wFbqngyVrius7i8xwlpFLiiUHkJ+qh+K6M
YF4mFOwBR6Nrm7Ylc9aGgxcuLnOzmG43gFy8sTIVG4DfQZbe7FXPfJhq0qhrYnZPtU0m6zT+MNDd
hibCUDlvN67gsSI0KVOsLGDnfISokXNuJvIjM+52gxstY+MHpskyGYtpgrAj+DT3Ey6NTv8dwGyL
SxOBr8/RdeFOvDJk2iFJjeVuP96vPfs39SrSe7vL7kPmLi5D5YtPbkfY4ITQraTgqxbSiWQdX9fD
LsmaqVJ92lcvv+JdCdLCxqCaWla423+zn3KuQ2YANlw8Lp9QxI9C35l82QjB/OCQ8Ux4pp7HCvd7
gPjuyulwW/TH+HBlCyx44OgxHJcX/eRgAjxtlzJBvrtwJrrv95jG76wSQTVAYq6MrrpOKwrTl+u7
Tat4jlqzaTjtr+MWB1wrNqYRoAIYsHsju/v/K2xCS5jAltCMWVqljbh7hJEbEsRXwnEc9hTSPU39
sBP87uG/yFHahnl0w8cJsaztfJ5sIWryW3ItzL1vN9ZOItcUxquA8sF8FYTLy+HOGw4lDB6XHMMv
YnnYp60SLRwzv9ywJocgLsh6YU34xzl52E4cQIYTAmFgDIG0+jats1jONUT+mREfMH8LvYz5lZWq
+QHdkbEwK2/xweFqSLRYATry0vzMZqvJtjvjDCmU5lKxORmNLRG2s8L0IGlUCFnBPH2lxYNHHZRz
CR6tnyEqt9eztlnZ62HYgc5KwrM8m/lHBvXxfwae1Fe4uEtf05otyOVrz/htjjb+KWcbTsYPwAUw
olcPdFAII6CITUDV7/N02Lfk9evtnadsJc1TMyvg428/88Q6/EoDCu8Wc3makByks7tD5bVGm9mU
QAkDzziYvN/ex0MxMkYZ9Cj73LeFmpYhLuO2B89elw+W5R7atQjAAIMKEHYdC5+nBnCkRqjPowsd
U3Dy2TstMUMnuDJBz6VFS7AVxTQr2hNch+K94SJ8JpTg3hPLQhb8F6TN73e8ewlGukOgFR6HNDp6
/gLR7YXQad65kXrm50Hm+gHhy4zhzcedZlqTVNZf5MzQx7pF/b02ySb16a/WFHhB/G1UKmsU7+3V
biGWoEJdAYbuUR3iiXzH8Ps5Algrvf+dOLIRo9TUp98rQM1v0dPj8KInSzuDmAHQ2Zvj8Wiis3kd
6rglGgdl7dnPki/X3Tk3iuXxvp0sj2BooSY0TO/xt1ushBUo4R5Svhbf+b5LiGP/75oTpDd2gzmu
HF47mV+4Lr8CAmAmNps9YK1lDC1K3luew39t3igASH0mGnrCPS8IvmA9kaOuRdyyY/MuVw5IXz/6
5O3zLiLdV514q1AKOl1rpOwYRSe27TnGpZyxitFMImsl4zLMeL9+cNHnuPYKjQEEUU4epndsOfEB
2MymiFfsOGAFWTkhttkwIu4+MEGn7L+9NDibXytJNJw8Togbm5CofE3zG/35if36cFZoXzddHEka
G9mCkkqj2TysfUyPhnRmqitXfKBs4tQOo+JNzvZkWy8/5rf09bO1hlC0dcFmqz1NdLJyTMqSnY5T
IrAbsTYh73pypovoauNB7lIdhWDkY8noLoPD8jRV/rQmcvilzPKXEaX6Lz8elaELkjAjeRs1iAMC
uVcqL0dz43wfyIQzDJE3/KdTTobYm059QNr9Zzh1yuLolYPjNS+ZPZYrTUxQU1GHiG2ee55jFcb1
JnjZpUcZkk+7Msu8Iyq4KQYt1IeQN1DmDUYuoxGs6jp63dQI3NYvqYfK+RAn5nc+IJMMj619limK
ayWr9AoB3+L3kC+9prJH1BdJI9iNjaBYxZku/nvQ1EP0aKcA3a1x2RKG5vu7ysLfNKzeP8iHvuky
o7mkfcImkzy9ITdFE7jMt51AwMtHAgOv2Z36u2/kz2bBUekXJ2zefmfdBffG4+V+SeZ2G65Jsgb5
ZQtpU5Q45D18y59SosVEVoiK73S7Ir6E/tEWMiUV2jbfS510cazjIc1TIwuNljlrq6EoDihFac8H
2oIyMruR54B4pL5wSTb8Vy4X3zqy3WgstTkD741MCMKXjExjs/wdOMYHRY/niH2g7JVJbPHwd5Zs
xQC5KcjPDmSnE8RYLF+Xb+U4nhFafc3iRtf6MQJS6s56uJN3DqNBUj/bN9sLUrCP4MCdjPhMcdvk
h6GOokJXNOuaf/K1neeSZ5IdGIIE4rBO4RSgxhECTKF6MYuRI3rbF+PW6Bz/9wCR+mQEdRt9IUHh
ZF8+RMxV45GiFvKIJ5YDkhBsDQmv0gkpIUfB3X+s/XbGbjuy2R6b5ABRJEuj/QO6ecS+ELOLx4q1
2l8O1G9H7KWMoQIXAjn8+BzSDwgOBxx39d/FGJIBNd3ZyD3U3uFTTH+EbtL8fpRmP25pwuUGt9ex
MRMYelSShtf3Z1YLIm0NbPM3am06mYOQsnmahs/gGEoof0WTHlxd5pnWJxh/yXy9OxT7kHJr36h4
vD7//lxxI8KmIvV5UlF56tcluMOrKg+OMKjjuT7VeZWC8YVjvG0+rBbLScMzZf56phhjOGGvJkru
B7KM0ueV55aVUXbZefxXzKHNqqdXQxcxO3Msu68NSvFKwwEaBcNiy1z+WXDVOLuxcG8ls1EwMyT1
Fde8Tz06BTMFnuZEdrFy6t4ODSIEwCzE7/D06U/yDr8ea4cCn+xVUN9ZTcnBnznvgeitE9GiD3dM
0q4WPyHbQprzcR+1dP+l3yTmRVQxA3gb5iYMmXJ7FH8XBb6BAhKyx45SMFw2+M3S8lNxH3MRNEf6
jO8Bn2coV6AMtBC3u8GXtLL83XVv+dQcdU6nGoSGmcPrFXDc2nLQVMfVv+B9DMu6bA1pP8GaMduH
gBIgqlGYdeSg4QFiM6XCV87kwAE3JmLjKgEkz1TLrEZ4Zs/QhkpjZO7GAdHe6qNDmnQmJuBeA0un
J9KhyS7I58MuI+7cv9ZWgoCKQldWuuY0THLvUJ3BdSeSmlMklE3j9GdZvCyK5PnlGGv//6CRIrnp
+d+ENzDOwAZgXsfJAd3KfP5NRa50x3LcAZ9TJ0RB+NKIeNLIJ9eW0AXI+/vV0naXdO1d0k4dASfv
JmjXokwBLfyMNMhqdU61bHVZub7dZa5Dex3fOqvMTKaUMuEHO1pubFl7nrj2BfZ1gxadz5mQvXf9
lQPPfbghFhqR6UnMXXyV/Ad7m0acj+KLwsYsRRhMqD4oK8/kPacOMA+/6zRewHCdEuLlUgryIoSX
K97JKg97GIuuM7aPsjuQjZDgBBcn4AMGIgJR91bDjWMexMPai/WtMv6vDaiLIimWk4AM1xKZpEvg
rtWozQQRvlBg8EiC3yPiaZ4fmLLZkMhpBkGUve7zAYxj40jqz58hQBP0LaSV6KcwhrbhjAcKo9W3
aBRlYdsk/IDbUtIGrWZI3A7HcqRJAQJqdLMzaHhF2Jb8MB+MAJMJPqX4kymxvM4xPYoRkw/1aMbc
nWzVCRA0RAJuczt5kB2+wCSqZxsh3XaUJWy5puBoQVDRGzkr6jEJPcC5Hihk9g+oATo8da9ynZXU
yydWfih+JrPdi7nuU2l5lCnzfKGgCTw0sxdIgaYlE/dmiZv75dc3VGAvN1ihbv8DY0UizBGEKyEP
ZZ8WGjURCoolqq82zGT8xDqf0z4EIueGp0OIZWK8lSGpdfvgt0tz8twQEUcr9Tv2Vn20jCLespQU
WOAJONz1fNVSG6BPJ64PYXDwtKDxvcT02gyKShRS3cx+TU/3UA5La/yO2VtKfHG+HebG4fCue6bO
S3ZLfGH0QVbJc8xRM1E3cX755O0QHXkDolPVFmjZphhvY1cgSuAfpa7vikAMUkB/OTljYTuFrlW6
jpK1STfbmbjUgxEuAsiYKZgdvS8d0UxaOYaXuf0bGA1usxDFpAB2M/gmQVTxna46YWLk3J8Jef8y
dawmwew5LM5zNg4FLfirjvczDTSZizRWkigVR+jN8NovIpJ6ofeErahhoTSMfZ9BnGeYcn7sSIh8
zU/Uq3UewjtaGFp0rF7d/0O2flE/+tvZ4HdOSwc8jTeIBgSeqcz5TZLD5gQKY7Uu+IRws3ek4x01
/ZuRbh5vqNpjkBqFsARl1XPZmt2XUGD8wRBl/Sa5yC4ovDa6mTlSP18neasMuizwxKaCUN7Rps1X
is0GYCXDhRV2iVufIpI+45JmnyLwRrvgSDyk6OMY2avrOrzRKs+nSlsfvWl/MOfx20zphknd3lLM
ukmd+icUd+M2StFoTySiKOiE6qRlTq/X9N1n8v0ODGs7UHvZbCR1IGOlnMd3cFzGt/V0nwhsDEAx
cwC7Gr5806hWpCvtiGStP63QBpLzmNaMUyHyKCf3+n5tWwsMj+bjDp2wiNfWiveyqF7QOAyEvexg
tmEFLuzFmCK10I6SSIE88k6bWstIwLRmVGcLbnpA8GDushCJZqsHx+KmCGbEu9xrAm2NSK8XlIY9
PHO5J4yJg8yYwhwOxDhI/9CVPiiA5SUwlwSGsYfGuDtygJbE0oOP6N/VvQPn3+F0UvmjB2JW6Xq6
HiDPta+NM4gA3gheCfprW1prM1hfqzUEnZXhlXv4eO9iqSl4jMcQiXSYWwlhpO515e8vI1jx0/3m
9CCKu9RKA6abN8nRgnrX6Z85lyLTYDXBxcOo3utE+GVvezR2BHgs2Dg0GKArvCD+wgjnxghps57S
AA4UIkiBTuHr658YMUZ11p/SsbIclHS4+YgELC6hebc6Kyn4esSWpffnGsFf9MM0Td5XSSjmR3D0
QHlBo0DyGJtWovPs/sTQRA/CmW2+z30PL0sYugJ1ZqEUnVlKLb0259GUPgV6aDLdILhofgUWKFmO
ECKma8foXwJNB7H1d2sLnC3/wnovE+C3wJIbChfdjHJALsbZuiBUwz9FP4Oadi6FS4pvKqlk670q
OPhm5VKzrgSjgItGigMduZouhSUkJaIr8WPwZINv8IYqIaxMQaT91F0xeHZKlRZ6lxMBTtdi9WYC
peqmiIFXcPUFPQILtqXS/75r77rGhVgIaKEN2+BFAAUtX8utAeF41oSuh3BZT1osUrdcLsE6fB32
IHfyAHPLc6O7yET8WZ5cFIGjF/n6B8zoWe3uDSD884VANSKTzpRNvhcSrJ9AqA5AInkOBQIkyIfw
1hUMs6/wkpmtbtK6pypd3Lqg2ecN3k27FqJQRj0LVPhBE6Qv7Ivey1cYC1ImaykrjuC3Jxgotm3W
TNp4IcBTX3eKo14nHGzfpn/vfCXK/86qdMdqRJ2G/wDTVBmesiy+/SsacoXl5usncHc9plEg7F9s
aJVvPY3a1fMv1S+5sezqdUQXzhOpSrIFjC9Nbu2HLhp2g6ei6vQPMrD7nI3D8JaX/LwqNAFI8oHv
CMl82QTjK3TRj6LRb5DNbo7bXQY/GxlQeN9eyUg7aQrWqP5Zq27ACTCVjOwBvpQ4cg6wFzRs4jZL
lewj+u0pa59RODyDAEuaOOCmdJSOQbAi1t9CGpoIn81iPSMeia1zc043KALfb11DhNDFCIDOK0GM
gtZsG3wFxVrr+QllPJUwlZlgPrPoRiDzcPU1yn2ulBVKAH9CcTYXSKkjjGkRTjxFH1i1PfZV+ufE
SNtppfP2iIPWaRz2y+G8uDpMbhpMNjYY9EEFdCjHDyZr7H8406UbzddA4QUrsvDQNpMFyDEuO9r0
zGnQum/wpOk+0cClwsMAKAhAKyKCNLowsqLqvQgbcT4iRdq6kClbl1sZ2OJHQwoSsg47UyoYC7+j
QAYQEqoxeNR7DENhlq5jAszQoTkkBPjgk79KQwOPYSz4Kr+XZXRs3p5kAcnFwp75v7QmMYVsRq5l
C3rPSLCSmY8ABUg2J8bfL+gYb44L/MgEPOoLRKACUgPK4tNHHJujuHFFq5JdaS509KjgXVpHZbH4
M3XGDTmR6hZX6apQ8Ab+YIhamlQYhMPDoZj27AmheU6XoUh526WbuUKnfk6S0Kn7GZLvlrceDIvW
2MVvKKupanCdVCAswxkSU9CdKy+4CcqAv+G13jDGWZaWihCFE2iUF42V7k06ESXOwSfXDwRXOjmm
AvA/bVTLQCihQaFEvlxfQOt7fH8LA4DY2bhlrjEkES42xBICCkxSxg0qwAzG1kHQWVs5/+y8IR7x
XgcYZ2ppGuE/IEP2ZYSmU71UhcZR4DFMha4owIiSEAMowubpcn+S3ApQLZ0WoTMw2WtaZNRGAog1
eS/7AwokwpHTVMRXMshKUDb+/S9coxxeU/ZqGjtl5aSdPFZmJqfB6T3ojmexrp0+8QHn4KY+/JP7
fV87r3SlVS+coU9wR0sex1A8od0sAB6Io+AUbIy7kWCx//jH1Wr9rYMUCe3TlV/nziSM2NBCrjMj
W4zB1VPy3krYLLnCIZsgug0pyhBOJ7r2xoVX9Kwqb2G5vJtszufuIvTlaXtLdhFs3VYufOZOXd1F
+fUfFgCr/s6RlXtwMjnfAUj7mEOMPrjcwvVk2EsyuNqaA7cbFDBQEoM/DGITBGQqDs99wd05obqW
kkUUVCwxQr5ru965mYGgba0KwXhay8hvGp//GPUufNPKOY6G7ST+Bbn4NU+Q/6AIfNejwIu6S0g0
fU+bnZE9oizJ+prRvuU3lnupypXzR9up2mf7tVJvjIE3GSzAQIVWoZBHReu0INhNgpAoA4pcErQ1
WDo8kMtEPZk0fjSLzwGBFGXVwJI1JzxGui62RvkixMXzTOnNTnfgfrbIAi+8dIWijAnJtQ8F7H1t
12A0OICyRyJsq6vUh7SW2eAb6Nba9ZPK3EEuvEq1XXiflekGgHrxfGqLk9JXf1ayOcThlOqMLGPy
SYIHAW/IM1ELskiG16xOtgt2oZ9bbu0Uo/1Fa37bCZmZFsBCebYjhRLDO7WHySMQwb8vct/PczJT
parqbAnu3yyQUXGQP8qRo3rX6UPScDZTR71y6E6E86AlGTdijdB2LRhxK3FuJDnQDK71ahlmDvgW
PWIpFP6DJVgpfdjvRQq0fe17iLRprdqsn7WQ5E3FX3JADGZqYuqiI+zpkAPyiH16IZ/cIJwIDKmh
dnlLL72O8aeT8TI1PAs7iZHTg2nmKkc4q3LB3zntLXNwSzQxxBUe3fsUyhL5I7CUe1/VYJx5//aL
N5qSlzFo2pMcHVpvtwwNsnmfUHYcxHR7k+Gx+GrSeL4sIGrknMAz/TgEjZ03EDVuKsLj50U7rr2M
ds2aOR5LclFCNS1JwrIQRWOUY3dc3FtN0MnFNNuetCsI0sLgjmCxIt9WpNOL9e/xmwtxUUDCTUXJ
EhN5HCRJn6ckJmEW9X+VBWzQRSdgqwii+J4xPCA2gRocs4a3dFDP6hi8gCmRoU+M6FaKrTUqR1R8
U6FssEHGUlVvJBM14P1NNOPbTY4TcsblpjjZuiK2hr0m9rA39STBO/Tb392yqq/PWOvST3cfd3LE
0vGFnwvr3o8tZEXgccaGUgZG5Da7nHbIeiis2SwKuKM6pbS3UcXIao/2QVec4hCivlTNRmiM2RmT
QpzEPJzgGI8s65Z2tt78LSn0lwNxMfsjKomgpizemyZX/P0a4DNiuuinJ0G+p132NKNHwbcpGuZO
nbzLQvHYO+uibzCdqtOlSAiWivaYmpjZxo7HIjgZckJYT2NUekCCZSqz1uJmisTVon1xHURikuad
XlOIV5pqKIBaNXwLVrd5QxKOEyTk4WPkJOC8UHWxdPjbMGHBUeptGObebbGpyc1CZOqDO8ul4mUu
CYh8StlOq9OG56pqigZNGZEj3d0NQcVW8hDVds3ChvN1k/E7LNe1GlLhUkxgn2uGeD2iqNguJv+j
MPsmsLbQSR3gozYDPWTheK8Tguw+Ivezp/PVruuT30TQhmni/WRhg/8GJZWeFyR7XoKRCBnhmqVP
G+K+rLs1cmIHo/O3tXi8liZ4H+zjQeiBZ1NdAFsgxq5uLDIL7XctQ3p9Ci82Sdq3bmB5CLP14W7J
gI7aPEfX5Osn2Vn0XAoy3z405I7EJad7aH876DnlxAMESczRjOypfw+vdHw8qw2gbXhKkGNgALfK
r/fFAn6g3cIQC3DHiutrX7CMLI7kVpZp36wfnzfyNIPoqRY4SWnN2+9T3RuEPVI43KHUeUIA2/TJ
A8ot784dBWMuBWpvweC/7kBG+piknS6Y0Sq5RlbO0eTc5sro35OBC5JlidDExHOwUjLkLba2uwbw
4jmpMQeUkQ6VlJbJmexzoRMm412YCguJaUk69oCwgr7+g+MHyH9ZvLxelEI2+Q+cgNNOh6IvC13v
/MHacR1h0CEu/P94/pcprSrcMxEvJv1OU+/qAVjtZy849oJqi3YQ6IUDWy1dr6F8DqUqBDw8h3Tq
pKsN+wva1euC0mEpQP6nU7kU6WxhzWSo/TxqjDZc7Z1noyJxyl7Qgip71IkbqLTLO6WNyL4IJpKm
kvtK8lF2oasTKpcfxqfEBVDXsnEXRVWa9W3IYZytroc5co3lK1TPOk4G24ztxySr7V31/c6XMBbc
rlGVZipxmSXAWo5MAeEfUq85zOA3YoWcgI8NsMSgLAA2MY4ySNzP3CvciFk4RdgwFnTUMkJLo56Q
mMi2ad+hJ/7gcekjHCyetvLeO17HugOVU0fstSsS0Fq6QukkaZhJCYCLL8jM+WgLblryhneBT/BN
Xhi+XF/NF9XxdGeCIgsoqR8I5PsNeEKnbvVyiDj1C65Q/GwRtqmdIiJol/sS63P5yz8cJzflU9V2
0e2fXixk/diLt/BOKibuxXS13MqY2c8ejU5o7TSmjtunBDpXBGbaZnaSwliQWLePB0zT5Ao59K29
VXJIFQQGaS0X1SpR+0eLTbEPXf9XwUsDC99qprU6fm//xv4nFSemuzrsBS3gioF94DhVFo1unJKy
IDvmJmHIrOODXgjEvJeyLH4rc82P9/LpGETQbUpVWZT43jJuZerw4hjpEnI40Yx5K1sPupi5anzk
+QJKkv3vxhTb+/OVa+8gJ42EzX0B0DBRRmzh3/uZc9JpZ+EGUlAftW/EEnQQ5jvaIhpMbyh9POxA
SRKQdOeAoX4IqmrXyEBXwJ71H2bSvWg67gSuLJ+7eke8/s7A/t+mbvtRzIvPWCF/+ie/Rks95udK
xo/RDNZFbpww79iQNYRUwP+f23KkgyeniO/6poc5n1WvKbqc/37gYZLpznMmE1bNNkWWkZyzG6T3
GNj5mRLjTOFL0TVa73grnxmXfFqt4FudG8mLd6ZWJzuL0szJJLSMnxxbQ2CYF2ZP0R3UUQe/pYBc
MKmPQrT8wqIeMEN1CJM/GFQ89Krj3SLFgW8fnsYNbBj4j2JsTyyGd+Pjm2HlY6q00Kahx+nqPz1m
WaUaupwIOPNFg7MIEgcxGJlLS6fXyeCJ3YzkDYamSfCCH9TCYXG+UaRA31RBowRVsKUmX/rA+q72
4xl1udWIGII6dKbT26i7MztnltHp7858F9TXjSgdjhrmLc9azN0WdIhTxpLuDDvshtF5DeMKiiSF
0Fh/kOEj5vCkSPxWj/e+eFBGjFBtYAG6OtiBX8xwVb12FlHKyYp4Hpri+iMVKuypaiQCMdNW2+DU
hgSsebTJ593DVxm4sCexvrSUhIY2voWiKtCpqd8rl3zuGir4/bRGBbyLNc90nlrUYqloo51kdHVF
wp0rnsD8cfE5rUa4dDBpzP1lujrpjyuhMRAvosE48A98gkfZN2KObpswT7vludf3Hkz0a81h7uTA
jq9WWxjMsZIDSuDaRpPLM0K3SSSO+ZU0zCZ4UPUl/g2jZN7fgPJvHhhOTjATH62XrLHaoZaFTy57
htVozbEum7UtNBVeIceaExNDmK/X4QBj3aiGapbxLK6ByR1Y5lDbHcEAM+DruX1Hg0IPe7vkEBls
gqSu11mBHq68N/+McLlXmwPuBpRugQTtqXJkx7+EJ7ent6O44REO1UfXTTJdUs8Dc+ZhJVpkfE8l
RlqVYME8+rLeOPeBVgABp0iKkoMT8WeFIYSG3xuOnNebwFGKy5LIZgVJO4QtCsDBuqvjzfOi5WiW
EERG9TqQ98wriOC9G04SryoVO7kzPHNJDlP8EG9DzNra2c6dHICDBettH1HdK2urQIddJg4IYc2Z
ap7/0PpO05/dQan/UGg0tV6eC6LWlFEPwejyxiiGEIzfRPw7t21i88J1GBVIWOmTXAqofiR+oflb
nEEVGDF4aOedvmQi+r3+6bg3DwMT42jS1xkQsFTr6thenw+0smXQCQ96kbo8GRS4oQOrXw7FJTAU
fAcBAUwkkff6mJtn2rQBMM8AqGDusf9X0enkHdBq+8wOFtKVVWKyGz9kF+mu3+pQaHAhWwd641jp
io1mfZi9EMbZpbrtBuccNtkqK8238ImKJtT1L8NwtjK5LZXZsGGZMCilsfD9y9FNxfJaOmpA3q1F
pIATol3bS/S3TqV/IRNmH7jEKD20jPLpIKhuHWDsNHfdiEcgo135OV3+mQH4Fs2MD2F/jA1h34Ma
65Ew+wJUtKpvaGzszB1QLsPsTavOasyIUt4DmCaQkrsFiAQBWcuLI/ky1WKuBaIdHSB/JiqnzVvO
juSrKgaI2SshR2qOrxvFZ2AsBThdKqhtQrgo/cSXNWFj1V+xjLwmuO1D5xqNmwmjdra4OfhbLOd1
7WVwZyH/xC5UBQGt7MWUf7Vq7sxCwh03I7YG5dnJ/qSdFuiZ0xAIw/GHkVB5Wt8dNEAn1rYRDhM1
B+wYho3GekAon6bjqHj11t3390XvtGo3gj4txP59/P4h6QrVWqqh9OkIi7ceHs7XHRatJr3xR70o
aY0xSVCGb7wEUqWGjsQW5v/9wQmtYmkY4a4ICjZxUQ+YLvKUzEYB+DvFFk+6PIOGTJn4CbZnzcMW
35u4Ud25RHNv3KLHZNASQjg2FvUDGm8OucfWqq6C+lcl5uAK4USV+B8IZ4Dvgqy802kZNU0TMyf7
HLSKohscNFsE3MYIH8pfuqZjy+C27zjGAN5nsnEIgD1dDeEHIbkluAdg/S7JQWPa80LK99m+Fxa2
puTQXV65829s3u+DB+8+Qw4jROvIVXSu44GUmQ5KLQlpCEH7B6tRc2kV//obEBgnkI1rnwF2mhJA
Ql9nDh30PS+ikIG6TAlQSGjrDoifJnYjD1dD9C32MbNKEGJNBYAIh9lBZcn+2AIYBOekSI/cRkTZ
kx7G5Bz8VeN/QUioM5kNsA+zlm1U9y52UwQ9dyRanvdzm4zkycPl5wHp7vZda+TAu8fnHJY4BiHh
HBJ0Xd5gMdWbn204mr6jt6+OmesjOOfBYpjxn9quywx/2vZNwJU44XXE8uo4XFWRwTZZZAjdwp5e
JiTbgg33DrbSKbcy5fQeFM5Ufw8sJrg7di1q2wNXSM+dxoKArKXDrPS9pRwztzzA2ukSHNA/bM5u
8YIbZrddME/VzPaAk9tI/VxjJZe+orLEAIPKtzccTVKTc68yssMvllcFr41C23B0lCRIhHEPbfJr
TyYo+hmKqYEl/bIp8yh//IdQYhFiuatv7z0DEg+/S178Id9PYJfKP52orLIwDiSESitRVbgG/A1c
3I3NWvOF2VBTRBVcopunYp+IU3f3bjynMOb5x68ALNiMtpeVCSkC+aF1jJUeelUSEyWqRVKbkWMq
RrSq4Ay5/GVLhQHVWaOg+taLEIKrivnVsyPK4lmqF5sEgn74/D8mZXNR7s9Opy/IylksEgwDj6ey
jtxnE3Npqcwg6dwE41995sMWgoqVs7kddWKJ7M5etE0Zg57EIeaJHaYOWwrH3+pg9cP+Err0N82N
mwziughy74u4C1ZM7EPSBwOY5pW2xLcbC6biUr7k7XQFB6/jbWJ+0/kDFZYMgTnZqJa7BxfKcxcO
od71ZYpHkFfG/l/ZNIqcT+NDR7WEUXaabdeDLjLfAR33lEdhnngYAlddAoHHGvOoYATU8iPuWW1S
RbZ8Z/AR/9KUzTDH38cvo+1HbzvrXJ6Z4k+BcD+4HFZmhxPf1LDW95a+6OIfTY2Geq05HyIeeTE/
vypXtTMrq5RqxgxhVLFa9MnT/Frzn/ZAK6ijngCRvY8C2MnYxMKEC0LAnKFWYowVh8L0YRcuWG7U
ZX1H479icmW8Ut3lbk7UTx4x/KKdVncyr3s/8PzuaPS7jVQLRk7AWID3nYp4CbNLzH6oPukarMVY
VwenJJfcEyZyLmOZhn9Cmy326chOc52KNAv8K9FF8hWf73J9j36XLy9tkKnDGaDn6YsR6P5B544J
UQgP/oUAsvoujXtv+pDIVL3sXd+jC+EtpnFMldjzLcTlRSiJFjA9Nf/xKo/VapX2ZlHXR6cpjyIc
O7anrSTu/1Jx/56FMztyp5+NcnxjlqvtpKrjb04sLmGmA13UUAhk51fH52FEAZw9r7I5LdNN66o7
SpnppBQssvEqhF0KX0g1m7j5NHlyxhcT/3eq72+iI5Jqzi9XiG+mOJlR/1Q6m1Ys4gOi+Fd84Dk/
7/aOVTCe0XWyDMUvuEAwFv1FewoSvpkqPeLOPvcrvSmwMLd+l1DFq5ranixOO7qC0lipnXSRYP91
t8eMwwf3t7uazSNHginlcUvctn0PJfKI/WKEbG6lNLoKI8P7eeS23Dcd97FsgdEzgAerGPgt7oMz
SpQjNbpAVB3dcHlNKggHgk8VFP122KqNwf71r0qNAkfMQ+DXuLl5jnAEXXUtlAmxRBnvqili0RgP
6yIPzZSysnr5SdyMoktnx/sQAgnoyGbhRzCtbZtVP8GtXeae2bHQwinK/SWshf5GLUm3pSQueLPl
ZPLMMetHik6+cLdxJP6VWlN8mmKHhvST7xZMpixCd2/pAgdooErs38LqgpPE224XUuF+va+KUM8X
13K0W1L3Y4MrzwnjQ0keDW1VwEyvRya2gQodEdkrbuSOkXcS76RzSTIWsOHsvoqZIa3BHYhQQATM
XuWNJzxhq7ns8jBO+8TAbbpaP7pmhsYP+Dn5MyWTFsyFwu2VQJPj5F3x8DL+TZZZEvA/CD3PB8WT
oY3H9kf3jCb++ILm1psYpp2y78K9up9cDc/NqPMF+ltroPNK+hJOVkyDP2yWQShPWMqC7e55CxPP
3sPFb0OIIdTviDeVwLNn+79WbcZkC8kRQY1s21SFwM5i7s1SHGwplfyuTomyVmBB41j5qfg6RZYZ
734rkCLc26T0YyuUy2somCM3Jx4s60JIsIaFdrlFY/25sTqOhOabExgwqQK/fm8HGuGpHRrmyVkH
0J+5m4s/XBnzrTZPKphCzCXAS7d/8z9SLuXFtba/+1HfQHv5RrneRtqoUy542jl48ewPh8cxTKGP
ZJLyK4Myz3zmGedck56MBZz3HauIOFvaf5i5jljRjGs1AZ2NbIx7Xhc3XO44nLOWinBFw38HQOj9
iubD5t2JN7AxYYtKV7aCK0DJjVwVq7OPpcZdeOdg7G2RACS/1NjyWSKzNsfFVntr+Iva+yprhTth
iXBmJ/JBgD7Fa3JVHHbkBY9HhcGsuzw9A5Kz4dy7pkSPOcfzRKEjuEqaK7sVM893RX725HBYwepc
zLdX5PCF/wxgZInn0f21PjWc08BDrPjVvwwy2HA9GxAODURvHC5Guza18B1NN0zYrz3LvJBaFDcA
i6/09VLKHRDiOoFmGQPF+eusqw07igJSi6onYQZiCPiw/PtwaWMu5+vmtjWGLeAnCUj31t0esrc5
4ZezmlcmJyBYf/Lw1dsqvVtM85pTZyIAxNImSX7252ffmucLFgTjpWFNaEbL1UHjupzHjkcWTwew
ib/7mbi5ZNiSE4NmDJHOsgxLnE53BVBU9PongtmaepBOt92s2V/UuccR5FPzEldKOIal6noNa1XY
bnr6Mn3YBguI69LEF4PXXt/Z6iCcumEWE+qEhH4AuVdNo7iH2ctNWfhiPe2zo1sxHACpXBrAq3M0
ZxKftop/x9a0HHuIQZI31POiDVTGOfZE91q5gY3G9UAd0nNmimH5mvdDZYLVYkstGkz1+l8Nt3lu
IAdYwKErIHqDzDlBrh6oT2APZkwxqkQLfwZX71LJ40TXJCgHaIPUJmHgb9fxgGkDUto/J+H904t0
lSnJgxbzQ+Cl7F/deJeueKiE427jfqHtS0hVboYtr/wALDOwzWy3Qas8uPLW1KRrmsvQyL2giN81
JHzz0HA9q2tHu/cHhvVxbq7BVVu8TibthIGPeh5FoK1TVbE+f8epE3GcBRs7aLC7k/W+MTa3Z9GD
mPQXaLwAijNzAdkkiVfMAgJeNBdSYIeeYuEeQjlswzpZYkdTfoc7geqYVjzNsNrfcHUKbpHX9UMT
pD7p/s/Dp9AAV58Lh9PJIQSwrZOfSe6ZfJfvbLpwvk9ju734u/czKmsHWCAjr/gyDiCueMNfam9D
lGw5nvz+bfRaa08ya47D2OkX/LYeapg5t93RcXO5E7miYcBWKxl3/WToy+Qkqg5xMpq5vmiAui2F
/in4E92X+W8gh7+fvkPatBEKf6yzbI0GcatF6rFIf3LzEM1X5HzJjeCFsYrX2nACZbRRbKqhu/ko
m1q739o3CvjRYS3FVohg7YFGoa03tvLLTkAF46N2+lpR1cO8DQh73KY5EXQqAn7Xuiay+pTnvLIr
iW7rDwTn4geDBmVNLLbeqrAVMGEEeOkToPHAJVjp+nY7CiYG65qvcXGtat1UVbaGATPASgaUNo/O
rc/p0bGF9QrzSIJ9r2hT/S3ftWz3dijLr7ofOMV3Gji05MXF8hCO3r+fv0TbfzJYoRepTy+nQSXi
wRCn+QjomvEZA6doWr8ENykSNXOtXmuZqkOWGiZL50d6tOh5UltA8ObHb1gIKHksX8EJGCfrT38R
ypj0+bVuuBFHvJD+d1YoeyqbAJ/Ra1LH8U6sf6ELpgGCDZaY/wo29Zrch+tiOy5xVSFStjMpOtwp
8uKk5542mGlMYvKymt/YBGtizAOlgw3LaSXopHTvEbJCuLnrLnGTt/wxgwX/+Ewh/BtA799+JNHv
eejG/3t8XRKUiiVbOVq8qg55JvKp0waAXpc7SC0cn0NbbtHEHLpCaS5pmHC5acoX0/gpS66tHFl/
EMVTHETu5J/jmHU1q280RAH0isvzld6fTfCdr165U8IPGMI056R0IRbjsCo7Lz5Ul3EOUu29XFYJ
eQwOqYjQGa1JYIGXYdVzmWMpT2TgxTqs/ZchdCe+ZaKPj9So6ISIpkKLS9mKVu2vxRAAmFhjWdkw
69c19eEXbQ2q4PNZL19aXUxlDVj0L8TCoEZp+eJXOkDPdORYcU1o1cSHlSCpALOiowveuoJB27zP
1fgVz9UBWxLB/xeUn7TvkgHmGHb7mD/5csGkclRkf8rvywFsi/hxKyFrASHU9bXNNKg+YXLZByfH
9+RidQdqV9UnzS1oetDmoI8aJRNecNjfhwJ+ViIYT/ZNjCie/DDqbjFoUm0ShGUmtMla6zso8cNb
5zGBqFoMx6KS7cwDWo/gSIFnSdtRrpKhbS+1or1TOiJDWfCnM+/Lx0V60Azt4sST/gGR2LdSrJua
PKHAqCcZUdLSp82ZvDu3E6xQgrcmT1EIl9ibW6YjDSrw1g1DyJb8pe6QkkbLO/wX+IQym+R7z9zN
lZDhoWz7Rib1wh7dMgTc16bNtur6lO35Qg9FnzereCKgWnxZTUiXoj9Ole2A7m6kvOPUStznb5ZS
ldcMT7JBiWqBLUzLJI6aYNESFodZiQvPcB0idL4g5JB2FlpFNquiykKmk6mGXOWwCSWX+aN8VB90
aJGTtFJ/THWZCsp3PsuUfAI5K96MyULvj7anWAFpO6B7zrpXYkqkyuHgw7B1ckWX+uqn34O3sPcx
D4fbd/oVGZwHpG9vIU0TIcYPOfn3FRc8DhXfGBs+/u2xIuKRicRhn6/XY/FMDAQMnjLHtdwWwtX8
TzjBmk4GfRCvI0LzbKzEPFvz9b8NpFhZUxFZjMpVLFtqeKRXJDKxTsfZ8FFSjVnksuP3HBiZblou
Ds21MU8h7vts9fO9e5mG8iVl7OU4TXKuetP3Mgs8r9npG/xdO85Vh4iFOB4QK+81PqqtX+M1iLK5
tB0Y27sb++TMJqyUIDXg3qrdkd6NHzvongh5lrm0L7DJTKhGmiTqHzW+c3MWa7quaEgMtJmfvW8W
Uq1aLXimYxRorTAd8fataI2OpBLwex//4Xa8Q/f1qqLNaRtY0FLTNPh3t9E2lkbOxkWKRLkYtZoY
OxFkgUcvSJcr86R4zbMnglBtFBbXkPe2dvFYBPcljm4/jnApwo63OtLrbfCPuWotwG+gYvFILjiy
nlH7qSQey5E2vyN40ZQWB1i2DDv7PcBQ5yHwOha4Wln2zKyENbl5l6H5EtKhUUD6j/7grVQOKbFA
JfvgduPchOUAMeLs+cAWx7vT73VYRLHtA0AT+np7w2fpex2/6Qq285diue7SnA9lyxqm3aLj33xt
2wUW+yx/Q8X4UdBR1VMpFZ1Mqsegd/TCMF3EUgMOdEVMgOgcGhNN5NMutkX1D9SesZEaLK0AOFbN
x3YD5w1mRvI4NF9W4dz3CFkNLx/SVndbKCNyDpOTykhfYewBBzhJGU7jYl4//jcAMIK+NrtM9Tbr
jNX2o4rD3NeQwksfuyp2TgVPirziiIJpU4pUSaXq3QNsLFHZXp5vBrtUQ9tiMYtxqaNpAFz/N3H7
oH+AvCBQXmVPuXiDhuziHcFMM8K/qKap5tTi9bbZsOdXmPzyM8cuhbftU5hRFbun4t1xDGuANpeV
5L5VAI/6ZN3+KeZzkiA6AszmM8KdIkaQzBt8x81j+znFmRRONlUhBkWpEi2AuAq7xxMrfiuBZcc9
TNegLGSafhG/zcxkCEuZhrq8GN9FDzNlqJevvgASVZsafaJ06llzof+4F7+R1m3Sdgf7EVX2BOEd
d0i7CSd6qFss7k0aRfRtWjLly8m7ZsNFW8CJfxamXGJ/w2q4vs2iIK3hqAOT8aHi2AxzRtUP/UX9
+wkg1Dql764TIflgZQn5YGfo6AJEujYn1WEZ6rLAaLbJfC9hTk1HkurNNYOa7rT1s492sLRusd1C
JTNFZoFXhd7sMTpeGxAZWM7YtILZ+baqgTim1KIytPYa6DUyQGRTXVGhJrNwwt5tsjk0a6k1OY77
0OMAdlECkfmqBzsI4YHPuza1B7tDTt0SbbuRcDBlJr0IWaygpCjbDETZ3ODYFITQ/CCCROBRLXj4
jv60w/egi0BfbSdZi1JDt7p4eKDrkIeP7XuPvydh++CZTKXWeHOohGRH+V4zOMJGaajoYAKYwbej
5ck2jEHL8XT30Q6c7bBrJYJ0amRnPyG+k5aTtHMnJxwnkJsmzNiAhru+FAMIDroUuYlBbGUbbX9l
vJSIWsdLjM+EIPZD0PgoOX0I/0N40FDN0kG9AnHZsdH1yMWUvajGF80uG0ZZt1EWd7i/8/0yf/hi
S6u41szK+331QgvUnAAaLoIc90U8s0UhEJo4c4jK/k+YoGv3mSSAKACr8QmNYPiCJQ/hUZGZuSVB
nGRdIHbcQTYJANHw7Bg4IAnKCFIA+xZLupU3sMgPPfMJY37v1SK6zPDJr9GZSeHsRh2rD2UTN3MC
loiXxMFqIay6gpIQ99roxzMAHU65KlKsSs35W+Av2ht/Kgr2vGrRWaYMR2u7y5FU8K86hEsumoxY
ZdZz+tZN/D0BHZ/V8Xbd1gKGR8WAyl1wNeVdI05Ykf42YHOggZgjGNRdAGjbJ9tTtDdTEzBoxWIc
6iTDkm3gBcoSU0vc58HJOGxJWbxDGhkU6J2Vfk/FLZjZQHGMIBZGOLtZguIJSPqef3PzYcrkcSbZ
1ZV4T7Tr0zgIr616GFRpRY0pjfHY4QFcVWFyHeaYNtqW1feyrgYd/YrWJEtN9QmeTMnaWEK9WreG
Q6Ydm62lZN21oF6JRItvsSxbIJ1lLvqOieL2jwW1gZ+22vtQ0Ekma7RI/1vZ6A5fwq39POs8SzUU
In4++8JoFSHDpHv8OYZI+c9ivy0bavFw2HPm6U/YE2DpmLZEc61J8bltR6GvOLjv6vum6qGn8rpn
BfaW+PDI9QpshrEbmWUNRmEmX3gxW/Og17Cr3SzfRbFWYp2Uk2UFc+zGFnIVfh+ibwQi6e8EDG9P
AhDnliF/DVDDy80uNMrMWCnTXKWf3yQW//gsuNs1AQgMov4Zyn/2z4bg2Vha35tSX2QNtjqlo4HD
i21Np1gdo7kIMgNaqn93B0h08bru/34hOxxqzOINK/zuSqX+GcW7PNYMh+nQUPv815NuOrXrKNsh
M0N7V5DMx0IE+FekoK56oMkdLivyKwLQ+9HR+iKW/+H21iwXepizPCcWRIvFfdRP/DFiYzEbS7QW
pOZCzAtlJv2PtQWM2UDBuzvjk9k+bFYFUZQefJxNZGblbZ+GLc3Zsc3LqLRE01OczNVZkq14tJy7
eL60QowAN4013I4fWruE/ggJqJl0vnY0S9LOAngsz7cD7VvetDODkLu2hyMBBM11f1BHXWlNsL56
yuaktE35YCt8Jcemk+rYI0o694snjcMFcSSIgy6NH2De2oYI2JkrqNX1q3xEhFlTQwuSEe54iOLT
5Mx7xYV1gz4YWexo2EE+A6XkpDhLpaDP+afyQ2R83lJHkYJuE0Muqgbs2SQ0q2K2aYpYFKEZmTO3
pVK9hRAH46/XQbiYOYghgRv6GwMEKWULbgD9emCLDriXP1muKPyZjDoJt+UJPoGogLviPkdnQ2o7
zum6sA23l+j866MEe47UPSQMIpWSzXSqg8noq9MEqOH6SU1ZP2Ey26yVnaAUAhsHH0eammO5P0QO
BZ7IdWeqWvVIMv47SM/53pyH7p1m6qfoJ59+6IKmqXAtdMr31eUT/NAf4t+0v6X5/AWgs8SM5v3K
EN+pmcUWLKfNiyJUzCrx3uqKS+XyzwOCGwepbG/m3fjBozg4W10ZPWS3g5M5iWqFuAuAAg7aeG30
rUlAL2SZQGo00cuSX8nBm9y2/NWbF9vPSSsv0LQ4nUgA6vgiZOzxZyRBKXWgBu9EN15l6UlMoH/7
s6XrzN9SRLXPgvO15q2S7bHCfi1dWFrnzVvH0oFW7RU4PwdVFvZ/lMkn4nKkRRLGWAkHLwuad8cF
jShMHJArbf15VAfFnrwQ9RicqXIZYR8TL0QsNeYdCwqZlC0P5yPFHHg4J2V1MGfiHC6K+wCxNntH
xT/hetNjl88kAGvHtAC0XbanHD+vldI3aBljEEmnc2n2XrpV0eIQpwEvAVIQBtAnFmGVPHYNcfqZ
k5X/JZVgbOvcvFE3cDjMaWaCGaaHgsk2E0ecM51VAL4T5jTSJdRX6i4cVUZ82jX684sopyjsucf+
vL3zv00oEh0FT0kOFyRv6YLgL2h+qdwAICEk6dbnDapgGqLac0CeYTVwZpGRI0VtnR521LAVJLtr
kmmTguI3a39EKHxkSWxhVVwIFv5XqVbxC0BTjdZiY8AsLMfx9wzy/ybYTqoHCHwBH+QxqomkF2jc
iUMoX+1wx1yKIe8j0vpiuUp2yRduyvdstKJiyrupLNGQH0wup6b692pYddE3FS0QL8yOMWAUMo0H
jnJZBypAmj7Q8FeVEmtrcep0x6Vqx/DsrO7XE6CJNoxNF4L9JVwYGtTzN2Vo6zdfUw40rrPcISl5
hS/XQzAk1TwRhnlCcX1QNZ3L8D8XPbqh4YlNyKRwrVTQuckJKQeuwHjIfcacSZMebLDZXz05gwSW
BzOanCjrHMuG2swdVf3bTCQCncz+6MbwMLhUciFAB6M2C2J3BnIfBSCiEk7JMbIZ+BGOt4RQAZRB
yZG10sluAMVUE8OXbLSic44N+iWxscamEz8eiYtoo+jyqUN/oXHs47mJnZksGVr1IZrGYGyoonQJ
QDODC+GMQ0nvtpXWRfjmWPfBFNbxkqxPcCigju/DJNdEbnbkg+N1JeZ+fLWxZWcXVfz/le37wx7S
AYx5UFN3gfUL+J3KqYe4YoSeniRDzeWd/Xh+FApeX6DWZB1L1N+8RldWdxax8WB9SrdpKfcYZINl
pHHL60WL8uXQGnfkNcHN3i0k6wThJt8WRAwlbReqEi4MYmntfDHqID6sCctbNBqjM/wLeJXSH4NX
/QQ7JeOdvxxc8aJWkD0ItLT0lM0UHsY7cnBiOFhLtmaQnDu5N7LzijBwIJocFYhT65Qfw7kV4IK+
zw3jUaqeAQxCXrmlxV6byiScqy3vlI1nP9Xp0VXzHjiKuVYQRLVZtZhBy9ybUK3x8ZOHoGU3J0Ur
ZOO8LecRZJHSZZPmA9f1O4eVWrz+B6WWk79pLiRL3HC12O5WGhwtTA/EXk23Ir0y+vkhrw2khi2x
w0tsXqFaYeHpqZfI+La0z5+KygdAWTwLg2NUsyanjeLdpQYwOI+khEGVdmBvQW0Fi3nLnRMsYJDn
ORvzVZVLdzbTQCr8F8ju/5qpy/+gkAKE5BAOjOkaK6N+LgLTjmEPlRAPaCMpycbT/K9rLuVe979o
Wa24vxJuMGTiht+/758QImwQtuVDzbcGlVvALw876MX4U05jYsDgr2IXbQD10uxaPQkDyuk1+NPf
wi5xq7LRUU6Y06PAHrfMp8IOqUu6YwmkCVx+QhLuwzb1lZgUKJWkDBMOcwRBLFvblVMXxgkd3j2k
0g70opLKuO1F/YgCVwYXY/EcDBfnX9nT/cKI2BWFwd3Jiu2tF9lhK08DlFggz5YZoRcPv2+dCZgu
rItuvR7nY0KT1/Qn8itlqfQFhBASTAOzNmkwQTVeqJKqjXpsVwoJSgxF9Ni+hbBxixmEB3+xroHj
XaoLA2AqhWmdUH55rkIHJE1UIvsD3/fiovuVlQYqz8NqEKwsAQjIVMzeMklMXhrwGYwFQJ6pmcAU
IFDAIqB9Vf2C9u3NoVkL5jkoBfpLRPLfvuO6Uu5rHhY5OX4w5n1ElaLkZ9IH/L5KZUQKP6lmWbPn
g5kfNqwJB6wDSXOF6jdofm48lTFmuCTj0FeaFpO7xJywCH7mbN8vHRJ9/j44E9nHsEmm07OMjpOT
RdK9a7TtqCqaawxrpJjAC5wXSeqlCX3EEw6wbJlM82sTqTvzn1YzfupWWmt8+lfOZp+iMywvCfro
nPP80Qisfypw1stGxjnKEFC1BBlzAZ8A2HqNBKNz/6MMa9o2FMfezYWBVxkeELpg5JII/Su99XdJ
Gh1+e2GRriH7ytDVrfFED0zImgXY6XxQUITGZw2uyiFoeW4nY73huUQaTE+j4mKDCJdmXjvDqR/E
xZ73LEYVX1xGxU36pe6xQXf7NvMn/3vlr7FkzS6Zs/QDK9fx2kzrPTYweuZTqe8ElNThzrzjEPCF
5NibwXpYE6ngIWMWJ1c4M3OsfdjlaqEXCZ9BeHI44tAUMT/RSM62H+dQkfUtCKFTmLyW6NyH1mNB
9jrBxKSXD6P9b9SMfcq68V6xgRnLWTQp95hchmszNnKtxzsVJAOA/QIYpXJeUcZOu0Db2vA5oNuD
W+0jY2j8TsQFR8VcrwBPw792iY35Gbb4Xy541q08zN52DeDAcHCsunyIdmW4n8T4ZdlJeBxlWwce
XuZE5M4qOAHDZhiZSfDEC8YdKk3IuRtgYHZ3Bn+LJYQUSuxcI9myUprSkLtGrUrBnWx+Nl1MMSZq
GziH+/PbP7UlqVIRNudO2OS+0nEaRaXzcVauePZJ3tU1H2hGY24N8QTUXm32awpVh15iObOXQk2B
0A1UjjZrW30aC7C05kmrK+jCCcf8ZA7VaKc5z2UYg6hrwQkLyEFWrQiZ3IMBA6vfWZjx4GRgHJHo
YBfcWQa6RhfpzqkD5/NJBGrG72gJHrgTQdQFfoKE8yjDstSyn5raM3FvuUbz1fHdqow9SmYYAbRB
um0UA+aZzR7jvl2jZhDPXI4A5Dau+PRkJiEX95EJ7jLiQPcK+a8TpfbB3tMvw7a7mKnBeYwecD3y
LtMkhwEhhXlSCNRUAJjMVH8EVFDKpeoPlhBD5MeBbREWcCRYVsmyH3Z8y0C3HOmySqMc4XpyYjLU
tlyHhxQuiaoenfW0SR8BbbfKvcOdwQUeydbDv2KX9tbU5QZvRCN0LPykYZc2rYzyAKFS7zmybQqz
469RA3vYfI5MjcrzXBLq9m1OyvS1oG7BM7xT2gbECdvp3POad/Gb1xwrKhAP7zdENj9SOza5i56o
YnLXivNvhv3AWPw657Pw/6U7I7bLOuU3iPXhY422lRAYTNNcUOSlNT9zDMkb7WHtVf8/FhZxj2eH
MoHBQs2j4rS3HG8vBVpwnHR+4lOPZrTUpBuJjS7S/dT9tIHFw/QGMAo2fm+u7UliDLDt75QBIOtV
kpUMXEIAZtu5XbE93WQqUcKmCdKa3nD+VoBRfKA3RCYXNLg6JfGb5geHyBEr/liLTlLnWDziTOyA
hzvUQnQNeC3pvr9vGtHWzBKOSa/T7bI0XUJXLHoRq9EAWq4tStqjYoAwkI8y5O4eXzDCPTF3C885
QLM3OYIJJdiOgCaz5XSDRXmgFavZYfC6ufZFjb06OVkUugB915GURniXe37vY0/HlbdVLxy5isDI
0KLboc0CaM4b+XoFGJYzFbkN+4f8aMKHiV+fxzl7633qWz3sBNhKRLHuEiW/guAHGlftBOgQ7DsG
CqNvAdieOOylIPp6UUXWybxCQ3qCwnjcnVtnNafJwlyJctrbb/gfo19BfgtcJ1m5DQQDSstQ6WDU
zn20/8UBijPe3WM24+aoE01T0UZ0f+AliBCrJ36nXR32O3jaKKC5zD5FPJmX328B1UcT4nR/pll0
7vD2vHhA2W/XXW+xfLLNvJehs0qnQNdkYv9nbZqf/wlphEjngdMKIYN9H50n2aGgfXXUEoMQoBJB
tDyI+wiTHiKOZaKo017yR++ANqV0vtJ//gc17dEsN6KTfUmLq2ERnu/xhUjHzBtsXl86tAKPXaNG
IUyDTDnwp7r/VqcE2v91J4jPe9wlkM0gUUN2yb2aVIywVzeJ/8Ii20b5dxS4fOAEc7Ox00ianzYd
iy1AT0ugVgtcbqGt5qWVc6tVlq+WIHXzKZaPFdCC1rBQheCI2jS9zivKG2Pe+Kh1oTWycY30iUv8
21YAGuxDnv9knwlcxJ2sE1uU7qchmcWfaaafwUUHqYQCowy39hLjhvFlSUypDlPXqQJ9SIVlePYS
aQq+jktSMkXohJ0YXTxrYClzaoVHHWGSxqn9+xsdrozf5bEwzKqbBYoEzYyOwCcbHTZDQQ1n/YIu
Ua78gBJpJCv31MBtRyQMFFBsAQTuTFDV7JnHQ/o/Cs2ebqlQebqghoq5Fp0B/MRVTW1OQV4gpSe8
cn0XMO4FWXmDRySJzyudzPg/S5+WQWq1q3Qk8rO+E3PzR1ypDPvlwPWrafNxi+bdln2ZCRUmdshw
ffBObTilMQjSFS2Ok7azGEKsy4KmaxV2C+hJfXGj3W1FgHMHiY7If62jFeDLAaB4LueIbUCk1WDI
LW+PLSsoB7xNGOLN6c9NlhJXECtMpb6qgQFdVRDD2g9LYyFn4MOg7LSCSayStOkmu2VEnV5kgpCL
I2ddnb+iTra4PFmss7dinO9kIiqz+xvLlYuPCb8FqwHNmy7MWMAmdFDTh4pp0Cz65xZQG+7g/5yr
jhFqlIah9y0m7CNQd7MGrKd7idY+HLQhW7Vz3cZ4oS1yZUgjNmrYT8Lx3okg80oqIwvDIfaoHrlF
pcvzUm486s8bAbzfj6s0IW1oTva0Ru0ycK4Tls7Ph2LLHAD4ujCH3PqHiBLDH+dldMLAKQwfqyEx
AAf/6uBm0NBlkjj8+gscdNFFboYkPXTWtrf9AFsugt2dyBDLC4/rfJp+EgQv7L8wfsjrC2ObW67p
mPhdlchz8x/78IesHwnzjy/h3RWU492LyRWDKwPE0Ddlg5XcN09QjDkQ3URuvMZFgEQhYgOPLRUI
QJW42FtgaWiWUCddYbTQOYJWIYXSKdv5r0ZUGXihseNu4qwq8N1K/+qw/Z/RZ/GnfpsTy7GvgJ+N
SBrs7AM7eP+SiUdi0I9z+7mCbbdRQt7G97fQnfko+fQvYm5WsS4kbFywUnKR4hOHolWxIg8eyr3x
cAerslGa6B+sf9KPYNsqvq9JxJoT43WJNbJayZBRWjQmsZN2c+rHCcafT/NjNG+S7pO6Pwqsy1cU
2VR2mw4BbeAJPqpOxh+5pD7hWdxMQ/bnD1OIR4J0brpSnHnBYhkVbRRMWHpCYxqT63+js5kOhucr
t61hqT9eq8krYS6DkRXkcU6CXQkhcH9TJJXwkw6ESfqggR8Z5WuK7oOWAAyDM35vm0qsWB787TO0
D0hKq/Lg9u2eqjbTpDKfVBluhBz3kSSK+dmdmIpRl/AfpdPdJnVYtjlzfOZF6ob4VlEVc3sFWzPE
Cd7kE3Xwpec/MhvLnEdM4eRjQWnC/ueh6IjshduT1OItFyxEU6mfvGZQ5e0KGZpWdFDo1HDN7tEG
h23HraaccCh3AjDLEo4ihWsJdhqzmAZKbs+EgVRqeaM7JTEfF5aOBwbK+2GxP9QrjJGkFBq7Bv89
eUNvSFlbBYn3kIg88SVC1nLAq42t/Rren5SDNgb0E03W9FRd+a5ugydlyYIEyepbGwoOsMekzpNh
a7AkomTZDrxuXqORCJ06Z8srmmk+TF4y/Ude9L2swQbFtIfKLXYNJk8Tz71cHtKaQCtA3OeFzt3W
XjXlp4TYrGTfgU2q93/KE811JHubj9sjrDpPW3JvVhKBV9F4SUa555UxylOu8vE5Dt+yx2s37EDr
YhAuCK3ieVyyfZaTXfgRL5BKaroBkOsOs4FfHzgua2pq7UPWrmwpdH9Lrpi1JkOn4ugfZNDfhpGk
NJKFlOo9e+CU6e0ek3Ty+OPVSJa1ZFuQ2L+gV/gBS87UTosKTNqI219tb1JPWIGo+rH5kEt6ji8D
SMz1jgRnOTTlkLH0kH2Pr1ZPIGM2/gy8SgtgZSLGemssNYeDmjd+Awq3W9uGsSFShl529dtrFDk5
3y7iIkRfJPDFtkAXTmrqIsCV+xqd5WOnCQaxXJoVsRCIL0p7yiepOmA6LBYdwr9cyfAf7EpDJX77
0rdd8lTvfs/0YUXyqsEd+E2ccGS6KjILGPdX4cYjzr1Oltu/d+wR4SYhuuFXqkUslxldxLbflQRm
+POjiAu+HePULKlkeCwVPqJNsh21fVxOR1uWR6L5r1XYwUF3h7hfBKidryQWNAF6kMB3V2J5KbQj
JSjIvZk0ZZMhLmHTtt+cFFYpqeDO+tnSKwdyjpybVe6+UybriZv5I3qxfqIUxjdYJsVZYBDoFaAv
nYiKZdZEDU+ZEXHXBy18/laWBVRpEWlw0cluBAXKltwVonuIMnOy6DNi9mdW50tT79AFcop1pQzY
vjxVmbjkd6baTBlt+EE7xGpReheQa5SxEBE0XNSoslZ4g0Lgg8jKpCM6kOzNmnILqj5mtCErQC5F
gb9iQ45gkhdoM2+iTT+jCW2s85EB3KJKHe+sd/x7mbw9GexRrXkfElC+hOHrVn6+qyV/4Pv5vHoR
kqLBb9LR66X+659dt/E05Y3WN5eAwam7FMeLdBTriI6SXr7SKBChcOP5nwamKFQvzLMibswnaze/
RFagVZ5xNR1YjuRrJGthFC43W7CKOUEpQTXCfOfn5rLpG9N4y/OeWKzCjxO6m5lZAgGeFUqB51oo
zfdIQJd6C3CF/UEAFfew64b43JpxmYWjQh91EYfe4i3aABkd/LE12lfdzht3khT6jcAlBGPMIQyU
d/4ZdFabNzecBJpEM4M7EWbJHWdkcWky8Uc3aCChdqJk9CFXJv38TD+yLmX4YNEUe3uoJV+Cbxl7
v0X/a2tydjKIEzuZ9AubNEJDr7AonfWxfYbCnNU6FXKoTS75P1bDgqNxHLgdvjUA9mzoN2znSFl9
6qjLQBbth1dKtrHm+ni25eQlfaRm09JppRfXZE4Zd3boLDG5QQhjihuHdgW1H/PA4pZdAG/iX68O
mGFdZ5LwL9MSK0iimhVB7Rp5PhqSY3Ew+cQ7n12zNyc2UFJ3NpykUo4gfQm8zhMTGuZOMo9zQsJC
8FUlzhXefiD6bDxV2lAqw6etShe8wLo+PKw5Jw6eZb+OZiDfq/C7Bb0qdjRWIFWjS1lqznRCRCHq
IUAtdOyz7bXDy274dZZiTBVYUZvKRxH1MbDyCozBtHMw/O1ArzbZJxaY9zk+fsygiZdf6VdGRLds
8O05Ia4lrRuXcDctchGb90DnHFNYLR2SXmc2gQi8SEG7mgn10vJq/UjCFUqVJW9jcvlwkfFeBuiz
0JA2QVq+UgGyuwU58u6P1fAb2Kyhk35DQovcu3Xg/VFJ8L+9zYF+0jsbgyY35uYo/aU+U0NGGieV
7gNO9mv+Kj50V2kADv37Aex1Jf6AB00U2CNn/WbL4oCKBjn4brQkWmhOfRd2F3p2diXJqO+YOswm
poK71EcDjxj3Pxo7cFHipEZ9qbKk5E7DKm9vApIqxmWyZyH1bsDLhkII4xKusTpSFBpZItofof5q
cW6YfPQbQInNWagFNhxvB+XdgZ3EgZ0t+ArxUuSm8KyDwsDn/1VR18nyln0yIivneXwEvVWwVmtL
mPmDNhl3BJMrBlBhZU/cANQ7vMPM07KAqPmgtU5ViuVEPsb26JnzA4tMUkjT80chuWI9bMrbgiJg
rW5Prm0+rVA9fq7KzhAZzNNPMcmlU09Y0AeeNMtF/MevbGPN3+Pm9UHSX9A4i4oAUZFYnUBziBZf
016pXMXyWjQOnpOluy50p/5VF5izO5DGdAFCIaV6KmLq5ojwYleqb7AdMfGXT1K561bt6w306nVI
dcYrZU/ZYsTe02eozIkca7ozrw7HbcKWIKTkDiIu6Kww9HpOJDi3CirdxqPFLJ2SWeKHhfSa38nP
6loLKVtHMRnJl9EeBLy8wVySRHlWTQlSKaXeClkAxoFiIP6YQc7m7R8vXYeMQZuRdC+QQZOyEChy
BxuzJm6fWvbdcNrUPtakou6kzplIhBWqbT5g8u0oX9O0FZ1bwMpnMEWa9Nx/7NwOdQCtl321sPQd
Npse2cZWPMvRF2rHWl0++mUtV5HEhg2jRve5HGKIH+321qV0YNAYduHPMLRFUuyBT0eBZ4bfnEL0
Mth+ytFyB9xE0zSmzvbkVxidEwt/SKneyXAReGx0N7LOJKpV3r0aKQJ/EndP8WvwQ10naDXThU22
V/OU/ZA1136bBkI8h2IaYTKuXwvbvRbJWkFJKx1u6elzjEkBkiucHF/nnHRgMTE509l6zWdgSrmc
rMkowWm2aQkZE09/yKG56krABchbsxCELfLj5Amw0SFyHJbLp/dbWJks0l/akA8LYcGeNj3L8LCg
u8gM7TI2N/zcQI3Hwgoyp1dm9OdR6DZEerRK+B6CGeSgMmwRsfFMAOOLaJI/Ty/Oj/aK4pc3Fnhn
hDW/H+g+2jJDAW2hFqkUPVY1mqWa7SP9qfxOufXQmCELuQOy05cNR2OjOnAmtznOr9/WbkiMILWv
sfzFi6XOX+DQiR19v3YAi3GQKKMCIGIXAvCa2nZMoqK/RjDNXSKkF0EGkqEoAow/5rRY/INUmoKZ
bMNZIxVTYiHN1jTn+MMbO3u+TyK9FGqPnnjQULaIZHXrxCOQncn9I8RflmgnirO6n/lbt5LkL86q
y9uv2jji1eNGVZ1U0+9i8aFEuWdZOKQHraaul0Kb0Yy69Wh7PAOOAaPgTpkjY5pHkuimgZrjYwYp
S/8oB2zYLhOAK6L+vF59mWmjqbQzPqE3Ltkg9DcV4yEEdDvarNtUJsX73LBSdhVwWPpUaGgal41W
9OfRkylEdni4h3/V5U3J58yrsP1KfTKQe87M2nIy5muwrzA7Gc6d26feuNskFC5ML7g8te2lCIwC
H1rPIQ5R/sW96LoyAZoktaptjS/nNRkRneWd1O9yKVNNy02OgZebjKQVj/5x1iFaHhHj9Lmu6V4G
dLC7JppOMeTXP8BYmEwFQi514KoQ68RZjmnqVPRv/epGa47s00AbBvqqUDHAtgqQ+TyIyM1+y3X6
7Ck6LdqlB7l/2Nbg/VF+cG4pJBrBaV0PjZb2zDf5CPqzmjlZVia//bm7YUTucF5U1ofLmVoWEsNk
5cWmy+2QUHd/Oz+Ss/WYhR0p3MuBlV9qWdQc0h3WCmS6aNE0sMVJUOrIWFb5a+jiFZ4dVrbs1Tpu
1a2RLf55Fcl4AwfRtAe/Luf89gM/OfCuuwgLENaU0EYi8reki9Ch1HJLRBV+n8y5umckwh6eOdqD
/C0k9bib8W6drzz21P6pRGoXALDejowpY7539b3mf+kqVJnjqSHASKac++Njwjhf7yemzcmrTNO/
f+He7esL0w/fl8l85CdPLQRgsv/nIVO8jDlA3Z/Thd5fEudk9/pEUrNAPlkqeAodrlU4nayBB5wx
6yNe74USw1Kl5TiL/nFZForAhB9dYZHvyVQQ6PTSyNMBX9AUyV1iI8iLb0QHPzzcT4RiBt9QpxuN
fdHVeMadLrj8Br8FelIbrKIW7zqMol3pEl1AbBYz+lqYea6BAssLlhwJi76v1i3tYolRhO9fjvAh
7md4NY1r9AUqmz3oqUohvcaOYWn6bNom+bqdsC1GOmGEGPAmlhxS7R7ANQhiLi4CMbnBmh99nt/i
8jrmA8B/kT457Ch09J5kJwTCjglYbNIj4j47LffiYMF/xN7nbepIOr6iX3l9STxqZGtIC/O02RFv
UxBQtswHpnM/+OZD3M1dbzbkIL07DEzGQCQSoW6mIRTa2mLUs5K0YDGj3IjFffFIFZQCl0ql0iZZ
wpei9nXgKfVkCWkR8wYnP5TAdxJZZVJ9foh8th80P56ZL6BieEjuzrfXolBTS33nYQPWg9sVT9tE
fIYs9+NmsFlJP04SE7t8XG1K7QjiFYtsLW6paulYXkFdSlr8gu8GwDeEMag44DrTtd3D/LxpuS8U
Dh0LyAR/tNCGd1R9inqE/UqrRzh9E6LqpjZSLSR4jkKJgvCj6AyuKmZi8B70ppQ7KLwzIrxDx1gC
ueh/XRoQemm4GWPbo3uZHzer7nNi5ueGWJSWjF467uGjHtW58IDtG1tMMmkT1qo9qGb1NZN/crVY
2awS8MejVa4U21knEWB6JBTwt08UrRf4ZGkr4rWpdxk95e5xZzDKT9VCoEbRXpUFjo8l/3xw6P/j
UAtwSw5gq4SbtlR+nHx6dJBWQQCsVN6usya4x9tpRIsh+lS77utbDoBoRwfWRtDKgar9AN6HK2DB
CTZZXxlMeSuwa4yFD6kLxV/1GSLGZ3k9F9jhs3OX/eOHllJl0WtgJfpbg9HAWvKqfgyAveR/UDgI
4x9mfmzXRUrl3OB5ZOrNoJUh6Ig9oakLSbcqxR9O3cRnOGis7agF21rM6mt2n0hvcT8TD2+11JC2
WHiJO+2D57du+T87kw01xUFhkaSzWYqX/p9RBRAhBlv9MFyNZ4OK9uP3cvACvTL3+UC3FRbe288f
DTG28mqCmI2wwEPUgk8iSOm973qvq0ZBPgk4OlpLwBMB3cVRHngFw5azlG08je1yqVk4yAyo/L5v
qEm2fc82XfLpmMQPnvo+OkFEpUc+tUdejpCtlz1ls1tiW09ugh9XEIC50ncyjRkv4eCFyBwzgIr+
fhwtoWrIyyOPm+uhm4JaMVgm3F/ZqR0QySUlCgOmMzHEJvhnHxuCeq+KGKHr1t+U8AM6+Ll7qObJ
VhE5FRXyQxNP6kMUpTeS0FYe63G6gU4ktezg21C76DOebEb9eqFk6dDzSWArKIhwFLi0e5ghe0rs
Klkeo3LySaV2fXuCE1CmompjYXB5ELjbN0cjUaLrnawvaD5qV5j/07ikZ81tSNzfJI9hImMApuO3
uEtFrjPH5IjTrLuXvj3FywW/hEMtKcR9PMttavmwSxPdb7hibzCquJVK0KBj4O5E6fjOI+5g1K3W
HZWU8kMHz+dl1fVn5ht1z8ikElg685veLwz2HP7wmx0Nd9frGnJqqU4f73kutXQ+orDjuEAQuZT3
dQOnqKl4Xm4NABhTTxEFRyn3mBVq1j8MdHk9oJWuABbrWCt9sfhN/3p/DjtPFtuqM8n3w73cnfD5
Xayy8R0uAt0idlZA0YOjB7+zRKWtrYX6Y2caRVs+00FqycgnLULPijJVCPC73uRSaOFP8gSV8lh6
V+WPgY8gXlS+mi7X0UnZGce6Zwq9h2f52ORMjgCSeNeI/GOxN1MTlOfuAKcGIv1yWyQi54HhOrVt
fi84XgMUzzGXiCh+1FyIpUbpl02S0W/nq+78sTcWSIxewfyr9NsgyY+llhFO6Y2BEuhrcxs8/aNr
yOsCQfoIiUZPc6LM+TNe40ghzeIRfAWtSqp8naze0jQvpAT6ieP8zHg42lclaf6u6S9wdNSN9rBZ
yP/ylMNMMAkqTVU6/TsyZCVh6eQs860exY+IL8Qt2vBnjdt+XXD6NNUO3ejCpozzqiI1QM2Weepj
zR5p3K6wmK3Met+VsYOVpnWVz96iv6102hbJ8CPo/RLBAITz0oFTrKu72T17I+bHrYSxdItd8BbP
lPY9AJvC6wHvtwbae3uNgGPGYASLoFiZYUioxRNypB7RfP5SKtQpv4fhpw3s9QsDhm3mzNK3Q+pe
51SXW+4PbmyQkW8edQ+kcZo3YXr+3JnUAhsQdLEeTsMdC2QNciFPTgfUty1aJNR6roRxK/P9O/Eh
WskFhHuC3nd29UkQZxwEyqswUGUNqRXD9UIcqo7Dlo+1EUEvxVc+hx4ychDIEl4uO7btdgglxr7T
9tnUy7Bc1ySa0riJA9cQmKl9AzMiYtyuzB4cHJB5rIztizsfsJJS+uPaRfgnyJITlROP64dFFd5f
PU2SXCb29E8Q+haFhsUJUdPHhEDm8k21B5PX1In4Eb+CzpAswQQUfaoZ5/sKDP2bj/neMjC8+14i
1FF7V8x2CLikzbcM2n3s++Dwgh+L2l+tiGkMVCiy3sSF2vNZ/WcNVkdPRQo4/tLQb1BNV5xEKdXd
yhsTzqSSCKZ6xiSOeCzFSvV5vc3G29bj0O7lja8BSYxU1YFZAnKKl55FmnU6C0zdC81kjStP/o4x
g2ZFvIknzoZmX/xR1YRhXZ3rgVK9ecA6SHwFftiL0YePErzp+Puo//Z2L8CiL6CdCsXeGKM+tPQW
8e0jhs4+t69LQEmW7dOtFeJ8UtDrmQjP+s7w1WEAp6STjgG4xN1iKA+sgN7epO7cUwfJz9V501FN
JMsgOE476f0Qb+Qab258yJtOkd0BzEAO2mJ1D45H6BNND5G5zif4P7bQPNfqlR7MXORl95/EOTnG
MpZW7nnxht/Jh/ezgUUuUyiePWUubJW2a0gFNjqoX+qupeXROBDxKvROWgikRijVnkXmg/C4rh+M
eGSHySGuAQBokUUPQ9FKALMU4KmrZTMmdcRZfRRgxcXXi6BZmQjAtPVFY7xwa0h+aHxqEtF+louG
7fCrKsNNyc+yrlT1U76F069WAN4l8wDhgl5LNsiI810jcsenwOXkq1WhYtaulsgsTRSmaiVqkJeW
KjgDZfVDHdRBv7EFHcCeginPnlf68Ku/F+/r3cy8n0KazhjXsg4jb7SGw7U8HeL/M4cagOMS2xMJ
tQgRC6FLt2eXnbQVaiRmSgqGJhY+FyRFhMA/ME091CZ9FYZAQLH6kCiIqN8KVf0CMqpZY+eibBVw
fYTGK7yc3JjtmVSPTlPhhxjjC2K1rH4LXrzrwvrx1woAxQ2p1hZN6ZBHAWfeJtDZjkrIVgeWnqxE
875YUeSAn8JWNstt7RYJiucDfH6oJjJOrMZ5EZJX/HqALh8ZNg0vUv8W3TOFAtZhQAyc+Ai25kY0
LWEK9jEYVo5Pw+vvy4vHqmpwMTRbaxPT8nhem6VbwB9NEnmdUQlE85jmwdQIOYNaNq/UlmbWPcUI
FHBr+X1xgkIF7ssqdrgMdgdKe9Qy+6AfPgL2kShoKnwyqHzhDj4A/4jecD0670WSv8PCOCY1RHb9
y/1yWfBPDXQVUA6JGGDokqwr8T8MfztAcT+6KnCIsztrH+inI5tjSlIJQ/RhLmnsMDkjly2vDDgm
SI4c8GfwhYCopqwot/AlAvyYnTsCOcwFLADEu0JmQ2VdWF3IZidsARkaxwA4vh3eo0/aBdIRWCHK
bi75WtEDgWkQq9EXl6beofhIv0t96F9ET62EpHBs9anP4P4oOpo+WC3TG9R38DyReKBbJOMhCMoM
0Zh2MTUsS4mNSD2Y70dmkT4N7CU8GqpzMmFcHh9cK8BBypn+v3oH/fE9Fz5zVc92jmUiFPmaeflm
Dv3dwoPnqqKIKaj7xSNHTIzFfTKhSAEQ0a3OamNQmN0R2BDsr5a/WexVOII4v95FWWPVGnZt9kuK
1F3s4/wIIU/TcImgUl1wveqUGdinop4w/iER5HQ/R4OPvwTlklgYCKp14msZNUfK3slm2i2CKBAT
8Mdj4OCkQGaTrRbmh2McuTu/Myi41tVKTfgq0fgFwHEov5O+s1JXiDqrHfIJ+lwpFMUYyO9hU4OR
b4duHhwvY9xYOZy44bup8HRON75YodiLMyWEwMep/Mj6QvNajuCITqKxkfzf/s2LuVTYfo+jb2aD
HStklfcSf0yeQfqPrdfeG6wLTuGar3utMOEcTf340LL2NJrrLUKfkPBPyDMYusqIH093KU4vommI
6/oM7wM6dnIKDTLxyTpFie8wvpxLrlbvis/54IZ6wRiTOlNNVtuG4zs3nWiMMyjIKKsym34sLzoF
I6S4FQhjYlvPPURNPlBaUwADi1oLfEeHzWXTqc5aMJa63MPrIT7mT5vzO4HYTO7xeQNq03XxL3L7
z/a+l9Ko9eWcSf147c/R2qnLW/EBl+ri5lDBBWPLOLsdZ9p/iUgEWxzgKSEYbiyqazQ2HKKo5jNS
rfabaalqbHRS6qdAbms3retYFb5l0Z1PV0m19c1fvun3YvpeO/uoWrsQ1zTy6lTjVDNSRnqEjZvl
rLf9wb65wbUWMIc5rimxQJoG+8srzEkOwikZw/HT2bnzZ+/86Ky1f1IRNda/T4shHR0l8tYUJADw
6MI7RuopiOP9V2v3zHkDUCPbdjKRtnaZvirx6NjNSU0MCTp5Mhw9gJdow+EVwyakeHAuipBudIWv
cCP1LrnTnLUUwRqF05SBHSAzjFpD5V3kU51oJv377XA3Gh4NTGZoICR6DEa/WvWMlFj28e/RvnQJ
M+Xp8LLQPESR3mxvtHthfm0EM14QVPZ9F0wMHF/7F/+rPZ84qfwiNouHaiWRNeA83t9+P5DJbqnR
BAV9DXeGdw2ssqFHp1HfcKJxaNcOIdihALXMmidVR4PaZO5oCvAdkRM/5vdlz6yUunUE028MqB1i
R/rW1F7XGzni6nflxyW/G5px9IaLmwI6X9AtfUmmEs31hAHrtZlzdV+YfGNu2GnZgGcnxw7q3aa9
DpBuHHht0eEEfCWQytPE+aeO9SXLxSAzF6CgNPAJcOMNIPoGo4CILsDTzsa4aD6miw96/Ai/ek15
fqbrKV41xfSVff3RU2vG8YYmzod2LoLqSQUwSMFTgyrtU05qBMR/vx5wwzLUH27/q7c/NBawGCX/
sElqjmeu1FMfBoGcJuzKpC2mYFtDcgLHwh7fPv73glpQXvVcIulI9OalZ6MWNUQD0xqjskNvneMG
XVxIKar/H9OFDqEKY4RsyMqHns0jcUPmtSx9trj9WKJQdYNZgBrUWLgwSrzkjL4W4qI1Fzq/nyD7
f6TRVeQncN1VGPVxaNzwrFTL2owQMWkZPVnOjEUJVgYuEU41YpL1shbubE0sXV7nnZeaxBxJQPtH
0OlGzuzZGpPFKW8Ka4UxaD9QZKChXFOW1JRo35e+8jeW5lZQx5G1Vw+/nenJT9Nyd9hiBkr85CWx
spuamFjXYTI+0dLAGxCF26jlsLrpU2/G7zsi3EmnLv7IBRBO6bBhKYISvHVtg7HJ4GMBxc1KQhbT
tcjQqaC9otA8BdZ6NPk/ybSzxIhY+Rnqt3JdT73S6dcWV7cgPn0HXhuOocjhQ6txdnBQS0Q9oGzC
SaP/O2i1qCupbvDmgdr/WTIU+siFHuQWbb8KAAyhlW1WF5mOOAkMQpjq6PkDhTwKFn4akS3L+0dV
IFiJi9NfbrzXqWZ1eg/v1r2/5m7uDzBmCOp3jCmCDp0rBQrfegNiX/BjWoCpWvLjhd57pjpwkz+t
BTxlFqUdT6tbrWA5fwpV2TTsrBuzbUw5SqlOVOQdFzEAmMtTB6sn221l135FuvDjC3bufpP5gzY8
rGettah/JhYNBLSLd2GcbcyJUoczyhFe0xGEg+Ao2oAfUmcSrchTJbPGgft6v3sTg7wCUSwgPv4X
9Re0sDGLpiu487xjUhDPbvSfB2IQzigG7SYc4kvqAtGx5bQbMXCFEAJA19aleOe/6dZao72WZjNG
pSTJgSDgI0kvtMMttELjWMyYmFw76ZkTJyFRkj2ux/lYxMLEbYaoHPjDcBKLml0Kar7ecwkB8Q5t
m0A/SqF4Cs3LRct1gU68Os0ynlhRI/jotEdo+R2QfOtZlPTpQg2OQusoQmZeDIoQPpxBNxUfNmqh
wZInKIvhuwyeqRZ7lEH1QaKcaSYvNl2w4/8DzlPmtx5L7sd3yxXteDzMxM7QJf4TZOYIUX9ufzMb
jIpJv5ECRap6XnX1y9wjPZuAXoiLvMxIYyGgpMqQbodFtScHgswpQ7Q2NqWccC6eI/i2D2NQuhuj
K9pXnqKlfFJu+hsHorDfR3ay8i/rZTRAICMRR5XFwx+df2tUHa0pK4R8RpoeQ7QHtqYmewqx31nj
VLfxmpt7ByOCFMu52twF/AQvzeIFGzgGX4o2Nq1Z1kHQHDmFePo6GleiGqy1q4fGc4bxFFnYDG0R
cnvwPycZpfnal4aHmYmYRX0TfxQolFquGRUn/TZghcIBSj0Ca4rbpqkamr6xbv+2O5PjvrWpEits
d1Ixn3zZsEl9w2Zk9P70mS/YQP5rOE3WktV5hMhLnpDYLeGbh+uLscKBQKwfHqfJ6eP4rir+kYQB
Ki4aLSN5VSPeH1PBkBQAR+WEtyRuP5pNXUcp9Z/nEf+rYk9RI6EUkdw0n/osDoSpzT0cGexJ7JpA
Hb/LmpERaOv/TsBWE0pWkvCYGQ6UT7WNjsJjD8uf79eYsWK7iTrEIF5f8U65QPG+uGMYlo8lgRFE
xHMlSmkpoXQHg3zrRRUpHy92rWmHbwnm2zIvh9xmaWqR8Wn4AxYCE/uZ7ziXCppRxALx6qOsAoek
VnsWfjgPxMVkayt6RIYoJj6/uxDJxaZ3SndT/htH0HLKBsF10znjdVrV9MGsU7l0BQfLWAGVX3bs
VffmmIzigLFO4wnowp5jv9V1TH8NyT3wCUnprUGHelrUA/qh9yasTbhUSURZY0byKSlSnNwULY2X
mbwkim26zK1IcPpuywo0G6E7tPpCzJvtwBsliydCX65iHY70RgSowjHPFBRQpzUfTTZsS73tGnzd
BW8LKimutnSO7KE/EZ7bRokGhoMFCQX+5cDzEgTQk2h7Uy4J7Sh/g9gggKIvHDDey6Q405UCro23
rkYGdnKROMdEE3qhzrjEOj/gh2xdU5PUkbbqr3VRTQ5MrpS/eDJ47kgsNXUW8k86koIe0/Ilwcie
/z0nDuoA8tJbNy/5yHZUmuYUN00ppEcPigJP65wJgB9DJVGvldaga3Jm2uhOfC3czFRLyzGDlQWk
nSNGg9Nuv/8mqjffKLnmW6EVGdmZHSwoylMJH++J75omqciqIcssDbP/ZA3cXMkH7IqyF7fbgJgQ
PIsmm7hP/toP3a2VXlE42ULwAFyGE1WiIwrQayn5BUx9mKPME+bIQxiJrjJp25dfQ3HE2ZyMtg5G
JmPl1ZqtQ2bQsn3bwfKK6bEDYi6ifBeNLW+OoUKm2zmO5K8nC5/WFZ21NzoxwVNcNHpQCJX8xw8D
Tqwh3GvK4iKkGZteDAGTodmoRWUeEhsqvrefkTh2zW2yRd7wUY3ANs7gDH2XDJbiQ5eHbEyLRneg
PgAgZgFL6EdrsuUxGgxbblMesrDqnvmbEpc4+WJxe/nv9v7nrNjkcTaogjjS/u5F0glwj7WfwD2d
7Shhj5IPy9a1SvLDvW/1sCCp+LOPiaPxsAgwW+8e93feyoyHG3rlYjbWgeg7CtTl4Sq4MeVJ/T6s
ExhW7+vQIRj/F/L2HP//KNfWRTeFCUqjodm8YXxv3M6Y98Idc7sSI7sKKv8hfOeGJ3BUBK99n/zM
iCYPNTRmnIcoXxQeEQFntAPqn5qfy5oodxQJwj0CcssnCvcrUMDgntsbFCovB0XHfc8gcg1J62FL
/PivG9yMtCWoYRP8BcNVPNpKCqa123esm8kldg80WhQx0foTfn8RWxJYGbecJLfBvufhy5M/LEQH
T6HN2D4xD2x5iIrp/74mUlOvP8AlLGXFxp8uwL19wk1nTqNkj4udtn1tUnVaq1ay9478I2Ae5jcd
/d/aiwz4e9v8ruCHkejP36bhYNTfcfb2XiFfOvCZgPobDPuFZKVZyhByjx/oYDteIQlDOUtsNWTY
8PgXDZzyKi2v/NH8duma8nc1CoqpikTHl9bXPfurrelWHNIJYvcdWvTlU2TNpD+jMOSV99dhWVMv
ME+GPCJkTPzDFT8ka++7UNd6p5MrAet6BqiZicS1JjKryW/v9BW88Et7zi6rrPFPR8XAuFclrisk
RXEzvLxPnFJjRlWkNyBvVy1KF35+4WnHobIPUdNihrdTHwf5HM2Sifc1wIzJFaF2JB1M63RUmRFG
DABnc6TTlsiOXHPWeohDem188m7KoVRlpAt9VfmgKcZNmHtcyL2zF26/2bFCoKhv5i3kVNjSOJ3M
ILt7S6SH/0gNl/Xt/DgMncs7wHtmpEUH2BFBSlPonumeILaebgwtS5cIBV+/0kl+I9Jo7ri1O3bw
0l66ejOmGdYCIh6HGQUS4hZidouZUithhkBc3j8F6VRWH3LNAHD3wUvnPzu2HcdQSPXAriLryMTs
bJqCRc+ovyjHs3wu8F6fu3dvstIQBHFtN+Rm8WVyZGx/+kz1yFesH1P5ZJLBrLYM69ad+o7VNWZ/
G3VgDL/zTdojhyIRLClKNbBzZn2CsubE9XPXROrE0RbGNjQZkyppnm2AWoRc8nlk+a8q7xGpsvB2
8jm6iQwwV+3AvWNF2HGWmQeQ4M9ZX3hT5vxk2CErw8oQG0fCTDKZbIkH3VUjivBeYiZ7JAqrTFA7
VRRDjLQz3EPD91iEAqgkEU5/Ihlg00jFA6lPpyUbq3Z28PNNlCxiqNHdqk0wKIbNzjLhPmIZx1Ar
Qh0MThtPQpigOrPt+OdRJalp6Bqyo9a6L3IMlmnKIV/dAOj/on7pWbvdWFPekbNSy+BqifxZSHW1
8ixnKgYFbAGZytOl9M3on1QC6qFdLmK15AauutGlKtbaWFs4Pro+tmRIjz8UIJPGP6EINZtdmEsj
4h6YcA6rueWrsDSrCRoGlRbqJmPhfJDHryrFN+ZMSEf/gwvIVAfxdIgJTxVilcSBlVIz1fouxptH
ZK+eZYx5h5V3936q84cGYkF0+bE7ChJE5wcCwl7dN4BarE4Ghb0BzEdQudu+shOs4tPPmw4li2kF
+sbLrNnWNPFTifeYndIZZVCWjZBH6iMt/BV9sqrv4bFgU9/KtqLSOMjDKF6YkN7oFl3B1tJMpvCV
O8JoWt3/Q94LM5wpGZC0zFTElYp2Ix+oX+COIFx9V2T/ZWSWYt3Y0TS1yJ4J+lUReXaQglj4IBw9
9X0u49u4Y95eoIGA5Iau4jZyKhhn/DvuNE6AQh8Y1y0ePVZ+fLWCr0ouUpPYuc2c0AayJWMrJM3Q
tNdHUkVJEM4b49RJnYliNW0BP0AdQyZSHxX9HNUzBQmqOT23ip6/boVFZWj7Qi7HB2bI0LbUiqxc
E0EA1oUX5RgdKFRe1kRCLd7aIH1I3cxhzJuf6K9P8gRhqM5wUvC41lD4mOXU6hsFFMFjST+grVYk
t4Z17OE9uNyH+nZQJsVExjnuk2r2PWypLFD05cIoNU8k9Krn8siYZU0hvN30eXrytj1p3fniZ0IP
ThaUnQHmguhnuLtxPW3ftxlvlDyNHBcPcl+U0/OSMbWu89FqLfAo18DU9kQ8vqVOjarmFs8ihdMT
NeJ84eUcMuLB6OgUy3beYdKvG1WnPRyKEyNRKEhlGeJ6bZHrYMm4fIx1ZN0ldZfL9cEy6j+coyKY
MEp74o7+v/OwNHREqNITrHXS6ORx78rzJSZi2Ogcrgmya1dCF77ypYQ+VBKQqqJZAqJJhUWalt+E
akKJpnkzxC54pjKDB3LqPmEv9i6knk7K9YJGgnTKkQYxcmWmLQW1OF86/UZflRR6bVXLZy8lh++2
miEoiPCIS31MoyA8UxtxHiFqK5WmqvQdyPVq07+NUorfLxfxvTbVJTUc5Yz5SWHyMrwpGm2UcfcD
aCTQ0tUC4Q2A5L41Mk6j7s4PbSLIEULSgNFYV8losLtLNMZpK/8WzwQ2LTGZMqaSImjGcyoxXbFE
pyggDEEwdSIhWEYOYHxlhkhzOEmua1OlB9nTUP/114YSCXPkPMY7I1N/yKnDzzH2y86yk0FzOB77
L3fHLNGA0fBG2k1RIdxaOny3xd61ajSfSMgp4OrTaI5MaqmEIdWey7o/W0XQ4FOqFoYgWV9ir9c8
GsO0Zw8aO0wz9qN0Pk7cOjDFr5Lj1K6lM8DhfLyeE+7mWUKNc/dt13YAOKiauRBWbSNysjPW12vw
X8k5NGGGaK9iUIq4ohR5XBqfS2/e0WzPFhe0NwskRtzky0qymcVZpRpMrBo2si/Y+bFQ0SvyORIl
px4uToGQ3qbzZwanuHsat+Q6fNW+IWPV6ZhdZFUplQV8il/A1x3UMUxxnbCdKPqhr3HFzhzYRwVF
/AgkRbpP0IhUhCWhH/dq/pCgKg2iACr9+Jv1u5mzXkDQb3dJXiOOJ7GGBRymQhZFGUWT9SFtj9mK
Xi9brdWuC1dmMpNuXT/CO1ZcD+1ze4rSulNtM5SopaX5uSRjXpmIC2D52wdOthrwYx4mzcKQvOPE
+lWSVQsKKFNWm9dGrTxafaF4LuCZh7yjO0AzRe1CRN3AG5iAa5gm9aVTb6Wi2mjpOekVPcUm2iU9
LOe9h2lwaQ/QQpnCC//enfgBBgz0b9UAZrqf1hGmSl6DrlIOH85e6/FTFestlx1B960cf/RD6lsR
pe6JCG00JW3Dri7EXuGKGUBDRE2Wcutx2zJlrlnILHcUs2z4HWNzSKB4/9GpNnbe9iaH/m27BSwW
IcqoDDxY4CFEiqvjmoaE3u+e/1vOKU/BJ4bExlfWrn5LksK04WrL3rcH5MmQwGpVEAmyXzMBxczS
ifcn4beORZLdQ2tvCis8Q7hyl/l1q4nWQfmUnJTPpvOrn3zJfxXUCpUFyQn0gLBtSq+9QcmOCNvq
rHkvxnwqeJCEXsjh+cAL3J7oyjQs2fdhB2iUEoWUe9Blpts3lMJUX/gBPRptymTBBf0MrlUgJEIZ
1KHTpM6pVMadAtippTB9GC4JNzVltjUc4l8DpPchX+x5oJQ92WHcgAgd9Rz0VU9Z5rWSRSOlS4s6
gqq0z6w9Gr8NtfBUj14fJXF8f4ob1LCiHMM3xFj8sXeY+ekeueFMVKcRPuRPVXUckkwANdLmSeXl
TU5MAol5aFjjgj5D8Sv35VzCXqHtyffDG92tSa+7LewuWqhjlj16Aw/ZWBpui1m346xTvSPw0d3m
eygTS8LZT2Hq1KaKgo0m5F2k4VhntcuPZLXSp6/6XBVsz6Ef+HzEIKBmjQWPPF4DJFbh8L0JXYSu
QReVUYcXQiLoUA+tqdad7Vzt8tK+BvC/ZzDTUylaWr7Tf8hBwHR1IZ6K6J2y/bJT8FkZeEow03gu
GQnVt7kt57Y/jKBDc6GdgEgGKy17h6s+BwWNLHJY686bc/GtNDYtVHFw5L6uW/b+V3ATf8A0q7A0
xGmtJ3ZhRNMPwyPhHTkUvO7m6X1ZH5gi5NUYjDzHKV9dvSuFTj15ZCg9lhXx6JptBc1sQ5sIFKzA
AD6aqtWBz7FXIvBs1rZtY3/3dNsxONhclgAEBHWwfMjzpxEc2/pIlmZlTrly+ue7dQXmAvJvLto4
FFAZa4CbVaT/m7GJNFOslnDDh9kfLPuXaSJn4c3aZS7hPnAx0Fchikjlj2O0m2rsDpAd2qX4RrT8
UQ7U3UhaMj6dqdKEDmOs+hmwNlrDT5+I1yUWvrkIvEfA5stg0IjdxzTf3sOXWRQV1QvoD3LfXdHZ
rQJtPMno7G4bUr7PO40ft+vqlKm9bupAVMdjxDOmVd16mae8npQONaQ8hwALs0GohgN8msmnRgNX
jSIEqfe06AeiGRkzFf6nGoZXUJWCCRBee5IIZeOfNIQVKpiDo4cJxGq5CNJ5x8Je7wiyyBxia8Nz
v709jxMMaPkmlq4MpZGsxgMU0GGcBs5oJbIP9z9Jo1UjD3PajQZ074JgwGUi0TZ1VjExnykwNDcU
2bbh2HrWhpJTzbkLQkKqFDYn3Blpfi0rbfucWlUO0DdbzkD9maQyvBDmF6AWi/poIOTrZZFmZnEJ
96gWWHRkaixkgSadsuL7iXFlYtPMysDlmrg3d5BcedxP92tITw1MDz4SFvaPJlYtu5Yydpc6ErQb
Sv2oX1aMpm4uWEE0UJc9Eo5j0r5XtHzVRoNPH5dN1UMydSC83HaxwcNEPpT/nlUX50Un5aOStyVJ
7+Qp1OXRX4sNGu9yM3MVQ3Zo6wDhCl7p+nCsXIPTp1jiT05gfNHCQ7I/PlZ5NkjDHecMRjoEUn14
/ZkVSWqQCiH+MEw1njufvIyQVouLvXwOv2DwJpBiZITmGGO003bUrMfahTdogBv+MFPeNnPdiA/Z
/MZyEUxRgmxC2/w1SiJ7JnO7eGctyS12oB+XxbL/HDSLjfKQwADuhCpPrLelSA22vzeO8sUeQcyC
sQ0Ye7n+TGBoJMSV8Jn7LV1lwAhmgJ8fnAzEzEB+ZCg+VvJEp0rFWomh5v5bshvtKVkkT4Ecu27D
cBQoPj/MEGFVQMDsYOL1sOdIFzDGIlIJQfxWPWwpKrS5IVvcWRG14yLx1bS7JqsG6gPoB6RlxFcQ
qsr7/u/LUTxEuq9nXMD95O10L3eg61jGeK6eKk8MVwq+9oahM6b/gQdwXakXVosuCaYT70bVPQ3G
xpLMffbvq80m9EEkWBXf2TlrmKLDb2itGn33N4o73hx+6H1x1Pnr+N6CQwLZEclvQpcxGtBkJAcV
N4wji1DZKFGcoigyaX4MPjBCNQU5PeDj3IYM8FpTO5ZB8xmkCbCGb4nsfQaW6Jh60up0KuOUYpmW
MEigvf5snOiajcVKqyTCXA+Sm3c6w5ANWM9KbR92IUdvciMHNeyBcXSW2K6q9S38IfOKszhNRoxW
Pp5SN9PsJRcdpA1gJ6k1GzlBwinMJrYk3sI8TezGav1WwTlcIv9lC/ZxC7GgsQyqP7pd60FSsRzf
UuE2z0OKS7LTYGh3Y4enqyGAVtFPVB7SYdkNgNto1+8SILKdyuEUFfdSy54jV/32eQm5kA+idPAr
o+mMjkRNmq1fKRiiAg9OR4ttYOi2Cgsr/E3kEafAHY3LYaXFBusHa5RiKupefKggk4wOw+hQLcaz
KX+RQM30uNfrTlfkijzU6Bm34h0N0lSdyjCAAF77AvpkzpzWRVSHqIPjmSTt0LD/m6BhnhVCSLiq
b2gm6jrikS21elRAUZwH3ShOqvEExCmef7vU75UcBrG8DjVaUwHipXo4SBXVqKUgv6xdnt7ZSWQL
ZWP4POB/4kJJnkdNz7VhgvllRcppz7KyOofy4FbsyN2sNlQ6S6LSjX1Ki16Vy/IQL+bNtNFB4qps
m7qCrySO88bVwFUxNt2rN5di8zB9BQP1qiTDpIP5Rg/I/AR37X1nAxw9aAudWnN3xkJFSSUz+esX
xAv1lJjzaWMctHlCVpVVa8D7nRfqZlmRv8422Bl4jL6huG1sT9P8tvLXlMv+XKS1e/bJ6gpg1Nyl
QId1iIEjyAsipyOXWPB6P1LMKeZcKtdW9waIIQMbfEhXqZicbAr+vsvCy+I49wrXeS3FC7DkW0D8
vBRPJU0fktEbdFAF/voz0vG/iiLUiU2uHSI0klom+qcB6v4ocQeW8VVyY7WfFw8jU6dbMgpS5lDu
36g49qdvrpdrKl8X5/AOGrMsc8cL0YX53+KD/0/vj2RRon4OPfMA0HyhJRVUaplD71u/Wda9/D0D
2KP4ODcNuYaV2gcwic3yaxJItfJz0Mu4jlq6q/ZwVFeFwRFzIm4N11bxDGJtaPrjSxBCwrYLwNvQ
uiu65EXS621RtNfZA6oGK5d4rF91FOwcn5vh9RRNgesFnhmbCd43iyIbUWn/Vt8IzbRsyhfniAx+
s+EPa2fS+Ps3NbPvpP5aHSsZxZplLBovDTaCjlAy/tfo3xCQNX6stDtE7y+dxgIWFbHE8oNMKsuW
2BHAw311dsz7aa0rXKnDSeQz596fOTZ3AIZXDfpJQgBU2kKCkLMwbxdAWn+5aFva1UmBEK+pI7d1
4l835ooaPFtKX6qv+TjhKTHFTUI+AiAzt7X2Rg+TCuF+DK7+m3z1vzSCcYWe3TAUJhHHO0pbjXjh
6LqUrDWtlZepIj9dq4xLcymrHbo4Vm//oZzvff1D/DEv2SnsqkRKlaGnuc4zRpy0QC3zauALHLCa
33SfqafTDJIJZkqNrXg9K8EnV9SFXtufAE8BsHOolUqLcn4BjKtIZKh3XDaskSa+4ESwzska4dpE
f1uDywpeTX8O3LsyfCNqK0HyW6a7xi6bxWJ2NIg6FtjX5qIIdbP6H9Xdt+suHJRtVlOovrBNvtXb
iC59w6exbu21/TSV/TpiMRao1qkx5aT8CQy6rWvOyl24ejgMXgG/6G15BhDA9r4geELs/4bwcRGG
QXlukGQEIJuIYDUhaTUcpYWjE7imqLxit5lzpbtMfBjjvlfRGdXnepWhk4UGFOcfY6udZ6FxMsDJ
Mt/TTbr7e5V7DPwqD/geziloKbMjMx2qMOaiT12MCws8MetJQzuSTu6nVj3S+W7wkIBz/5U+awfh
aUsn4I9NLLo/S1SJoFfedAFJhyeZQ2KXtEs4NXl9jadWhCG4SaBDneuSHnaXSmNS7xoMpDwiejZU
nqTIfZbyLbtIYuhs63He5XF/InKMa4XQdawQnxvl/btLIC1f27+Ib7WWc195LddT4Rs9cDqdTerl
GCiCt3sGLlWEOhe/j/69BQ7ap1rrQonj14R60ijkQnaqsBwn9Gl58aOQ7zAqij3nAFPvvsZ+nr0C
uY59zD+9KGEp9aJxLQaJdUBJnAFM/dqfLAPi9MKN4MAy1Hb/nbCay2HGYiRW/oRR20YF5IyClF4f
glcgRXLVsbCNqiyrj8Cj+Rab3ykSNfTPv0OuQFgj6wflJdCtPXMT6wr4+mPdWyz58pVy0GfaOeB9
5wH9dVISFgKA8WZuxh/FzAWBKxxV+HG4ujuwHxhBHgl2tZH1ydiNdBAfBNIpIgTgfpUutEG34LzY
kRG1t4tojQSHtIGt3PqfNkP6YhpzdLCH0GD8ixoS7dBiWZNTS5l3NSNztwlcL/TQny1ikfLR/7pw
6p+bdC0522LQ1cVkGUcCttkb6MYlFJAvu/QsXCdWqmojnd9447j3xnjnJSEr+Mz4yJXtCS31oVxV
Lv7cZ7k1jezU5xInlkGHyeLzPKwfze+eo7KoGb6yH4S6DXG2Z71gKG5oBulJ2ceixqjTNUNKs8AZ
kn6BGJsSCX2dr+c2Cvi43MVZ/fJSbJLbqfv7n2ZcGau7K4/i4LncQoezjCvDUzqp6WUNzUM+gyhJ
xTqSi+6Cl+pypP84WkZHLTMkueGXrYTEsalZNgwpmwC73TYoW7wPVfIQ9E/uA4Bg9He9+x6DzdY3
WCS7F9evwQMlFSqASqFu5L7m8/F9FNYgt0NBOdX+mmxGuFs+i9zWuFAYjzvilComScgOGxAmmsrt
QPeZOLiyvQz1LRUQuBDU3zT5tvZTFU++kmc048P49dZ4WrsW5gAVB2G9mJop56YL2vgQctysxI7w
XMDEg53spoDvEfm492FOCRpnVFq/IAjA3vvNObwmI59LsR/k53fHo0EmSWM3GEBHW3R7losKjsvO
eQ/YMfcGbEpUIpprtlarLmg4TRMLSb9beCLwvQ7/z/FeE+AfTl5t0CIAp8NoAQYnL2+XhdKhb4FN
z1LCa1PEMj5jciX/O2BGCYiMvMh66FLbY3PMhARhAx7bcb8ActU/mu+IbgQPNz/nAbObAFUkQGLA
pdoyAQ5TD32/aGAnfvrFzwOUHyPT6/jdejiVi3v+LMnO0sxlRRDwhW7ysBCiimBakgkBROKm3Ohu
iw4mA09udyrP46wzFrLPFubc8QvWH5rTn/AEDRl0KyNz/BURkl1OjauOddOmo7ZyIvhdzfVCHR7n
oZ7xCbTtMRM1dMLuvzYMQnyTJJoXTMpk2Z4E6qEz0hfU2RzUtDlCbbGAIDJi6qJ3HX4f2JA6FJ48
eIITONkOyzNzL4Ma+vN12MeDudVBLM0G2WlzQA+bItWEdIWi9LTFkMWJTdz87RlMYCBp6NTAJF3k
qY4ePuSVZ/pPeS/DOqnaedZVdVEaPja/7zejBjKOnyXqDu6v9nUoko3SX00FRjYTosKzcxXi6kOO
f4Edb6jmZ0Onw5ABbtbtfbXdXPKu1ghBHA9OA8kZ9CfwrDHyBDAMZd5gULJqCQQK5bCCH4+6ZsTf
VhRs1lbZUIxjQ4bTGXj6im0jOuFb5k7zY2hf1lfYdm8mI/nUf1xJIsqmkAUUOjP0Ffqvq809XF33
m2omWUM8mDv/DAoxf5ah5OPFDJ9UIUV7+eE2Zmx7HRySxvAUcPFtiLRNU+5hr4P0iMbiJsy14dxZ
Zh8djzv2qar+uKeS5UZRri3B7Ri7pVZMsFfa459vq2y5Sx0UkcsNs20ydu1q/rUa+VpkXVzzCxw0
1pIp2N9XTzt6V9AYbqHfKzhjg1KR/lT0xuPbJFj5hjy148VtMsAOhY1spOcq5uO3+SOKCpeaF9Uv
jDMqhui9BKd1r3KpMUpfjQOX3NhgteldlJusiF6zKUNSBmDsiIMAr2O6hRiBALKuzLyNLh87Dcmk
13jINW9VltY7qmSnPjIe0kx6qSSECLXHARGgJLq3Mt0AO33vIhSc6tP7HuNnp6oSOsXEgeHCrutd
siQ5eylzz1a5uNPr3fIeIITYTjqrACPWCVqknTKVCR75DxjuywxeLNU6mwBSaWGzAttdGV0UezPY
BM6nhBntT+PD5UIrYfgk1DsWRxkCHzvroVwKMX8hJua9NDJMeE4FMagO1RFKDVY8n6KfXgX/MviC
ESH27EHmDEI/k6gHH0ekXyB49grIhxYk8W8SlnGFv5xSX+5oogJ7nZWKhqvgQ0xS031LI6QNd02K
lhOCzMsat96NBmbDzVKnyY0yq1zmy2o6tdXdpiN5nvvWhktwfPb2Bq2KcphWzFiN9HfWRPm5y9tW
RZfUcyE+bdXAM6epahv4DKSC35mzcG3sYHwZzzHgP3+VZLdxXZ2jsUznb933k4c3ahKtHGToqp+g
k8z/aLcL5FVAt6pkWD0/ay19pnwELvhENgJvgNnRLIVL1P+gRPPU9vpf4mNiBo0saXsS11aKSRaQ
x/8AH7+YRNqfGfUlyhXQMKAhsNZutl/Ssatp5bjEAWfsk2famxbV2KOmcSrz2yVh0VgvIy/C4EkZ
+CPDk2CbpPcnpLUrmlsaEOS+CZyndo9etH9zI/F7R/XFGwgnZXpuIFzTAJZ15aDoBxrWSch2g5CK
BQXO9zHcQWdKVblMDzVfunBCfwvKVQpCS4QGZ1gz+qLKycMgR6C1JYjmgSEy2L7PmlspdhgnXRPs
rG3L/EFu0uHRf+wPMWEfq53em/JGwLI6nAXuu7sZOAi7m0787A64PEMFTkDgFXfqNvyfhIHgA2Ur
xJxf2c53RB1hlZOxwedh8JQE9pjSXhEnr06NfzgqIJjCu9ewQIO0x6l9yVTZQE9EB1O+WPEVNI58
2G6z3qHKWqXr5J0KFlv08nc4a3WG+G4O5+junzLSu/2DRxcGZxo5IFa5YmociuvYPeBDpK4JtTdJ
RkfuWPowSCrsXOqPtsoy0Rtc0bB9xpdh4F+74bhfsh7TPJwxd0GaH7y22Dv6t8Mj5IRUGBewZCMy
kInxWgSt2ARXTKjYw4L1kX88L8tK/ehUo4nyyBe2f9+E6kpOZRLFYudnDqhBxM1L1VzVpqyMZpi9
XpEwBDheD5JOkjVB7Wqej7Bay6Y1NA4ifkOIwXDAiVOdwIuoUEhGpy8vddV9OWjZBNV/2HASxhyT
xuCbKM3/od3FJMTZK+m3Lrj1CZdmqmLkwnwPINX/K5SwCwDtrPP8fc5JiPF13JTfouTpoDAoeNJw
q7oE6ROwM7YijloL7DPX+R/+Zeazb04uCWbNySkcUNBuoNQWvll4trT7qTbwigA/Jt7KiL00vB+3
AAKXIS7FMrq8Oust8bBXXoTS2wGjUttl6VQsfScdPtlpCuGAT6jfBIAazK1PTLNv7OoYCVAUKmWc
ko1haHSxmQ/zYymaSNBeI6g1YRT8TG0O1rS+mmX/CffnfMxuD7E6kP4Ia/arl9fWWYhr9375iRsn
7CClbqLPeSZ+Z/1NjrJ1mCqqlxzeDc3TAVRQMZ395Kk8+IE2AUviJqyJq6cSWIdfp0Rv05EoE9jd
h4whagHRD2twOqpx2SXxUl4FxmXsM6OxLiOaw8o9peVawDj6FdZx7QM1BFViBvKdKQCGnjvqtZSC
TlAwcFmJVVBzCWC/P/Rm6grvFI4Hi0Kc2g9aIEqs+yVu+zcywVPq8SxALfFAJqiIF7+bkLmIMe/T
oq2Pj++nrBqi9/HfRe3n5xIWvjXavR5r48F0c2rL0B47juJqTwj/jAlHYpk7gYnjTsHCCdqqlzLm
qrv1vrA763fPsdqtJKhYM0EfoUMAIYlacn2/ZbghfK+DljasVSwDYkiIGewcOiN6yD/I3UtLEGdv
QB0etfmMXsisaYvsDFbXdZ8tL8+DmJoJKiSamCWO7ZQ06RDqvWBDmhRtIGZJXL3/xwMIGoY/bZRM
g1GXxGs6S/s+erzFoGkQSM77k4rlyWOy82rvHxFlwl4/UrL1t+w4cg6RB9HgQOQIHa/sqDKlY0Nz
mQ7IO4C3C+oyiTi0gdMPDvNFBpqXTtzZhAw9iUMiP99zY/ACg39aVnbaAuTKhf0We0cmaqR5aMuO
zOImNp36oNJY3aKuWng/AyrUXGWPZvlKH1LmbOm1HBRuIq1ZReb2GSsE0S75n68ir8+3sPR1+6Pd
AB4DxEYXfXsd7JnhHDHWcRv015CzEC/DfaLhlgBtUmFSWCmhoSu8cLw1hfkwgmuHme5EA3pnC+yQ
NpuUyoTDr1F3+2hecznIphDjcs0AGQmFO6EbrxZbXQwt7vMF1USO7cqWn/QDApxiGAUZTc0zik+8
KijWNWm5AbqtAHyCuINFtA/qhXGTzAL+dNJ9F+BqlzYgkFoya02CjYtrvPAfjifMERjKSbjCgGN4
uM/jxQW02bYlyPmRjuEqtCi8JJWcdv4umWMLK4Sy//qx4ugs+n+45m9CLr+MMF+PPR1KIz7O1deZ
tBxBzkwTwbkktn2vcthMyvomfpYg2jCscoHOIBl7KqKpe0mBv71xwkyhgf0cSEs/lQxbBlq6QYjO
ijdRU2YyfjYG2hGN+DBc6hoPC7AlzDNy+wrVFcHPuwPd6nse3UOAxCMWa/C1kxNsbHQvsUr1aO/f
rpH8/jYkyerJ9VA38bjyWTZjyVr4IKcehZM0aYE6nD8JJdoPOvqLNn6Sd2cmu+nZtz9PE+neY0bB
wKT9K+shmKgtQd7FB88+3IbpL3TX+1OQ6mO6DrQt2gGIZhL1t9qPbQikpeQj8SIohnit2Tblcwqj
0SXRHG8FXTcdBr58Hem/nqYeOXdzkbjyULn57ADjtEGGgqQnmkcna8ht1kwRRZN5W8aEykhFLAeG
XkixdZcFpjaSKgfPpEdjkSn3yEaAvaUutm2/KpFbF3qf47/II1D3D0e0G1hCf0XaDeWHi6DXxL28
zmYYcIKJSfb486GVivAdu/Bms43XusTtqLmRfxSHBInrwXB3yCIWTZPZCMGKE9FYhoNOKB2SS3h9
oEVu7bcEQXKO+rV530ERw7dCkyf99viwno2BKnlXBDEdlMwCNgESUy33NalkqvExvtzcL3CQupK6
BGf57SB682WyjKeclK6Bxn9OrXTsVsuB63+EdGbocVIIOnhktJiDAqByy7IO3rODyUdV4sMJVM2L
s5xCeTs4bv2/ugLzwoVrt34CEcexVrOcqqxVKANi71fupeo81QXTmK4/85U2kWpgqdDASMTbpwJI
LrwwfPfcThwu0CnXAWwRtuMT6Vjf7Q+M473kLq9JDXsknUYMwXtECzqD/sm+zsHnIBEHITRN4ilf
wyGybUnGzzbETo6DwZJX/Rg0HQ92PNULBhr5x1MoLa024HxkCSFLdKNtxltUiTYPRlD49MNIPFjL
0sMBLI/BrRr6kMs/WxsS+YJJDW7cJg5mO0hr/zXT/4IJ0fZvtKgups84JEpt48HDp8kzoRgHHSOK
YwLdy9gRIAjOZ8fcPhn8hfg7SIcRWXlAp6BEH37UiJ0OQ1DJ1Tc4sTdtqcc2zQilUCNDLWRs2hJT
erBy+p42JmmWFe0Jd19UolLlixhZRMg0HEc1TQn1sDhs2HJ5UeQL7nU1YWU13HQv8mk2V2M9Tgyv
gEUVbasB2NOoJgL8Y8Cp5SspA0tzogY1kMVsRaqJ9VqG/JAmkSW411PK9Wuoln0JgUP28rRuVWS2
4M/2XQr8WnqSGekpsZijVwsHs/YLwx/gEPOIkFo5IGYQn9jnhBijoeAWjHix6HCd6r5RrrLtbu8t
O321XsBMGQTQWaVYByh7tcYq/UhmfTqN3C8VSUz1BXGaMIZkpyu4lE239DAYBwqlyl4JOoilxd4G
Ig1mSAr5TnSZbguQeiACLeWSFFdwBVRu/rjhIh3a1tgp8b/79mPi0n+f/o0avLIk3ctHk6xCfzXO
EGQdfTdccqeiFwewibMzQvHmT2X20aNpQNYp89ALKuBfmrq74maVfvs1bDQN0oQ4DhSViGFjTUWj
i9UeQ4P/eDl3K4sDEzp0KSpWX//SdC3bVW/29d1ZOQ7hAzhy+0YN01TixRpGqdHimdjMPeq0EZNT
uagTpQwziz+mklunx6neULHzTQrFWTsL1oaIboHpZEwcS+zH7qe7WxrYE7p5ajkjhxFQXtD0cUDt
q0lZFaqowbrpMUBZehocTJfupxjmFDyr+ACVtE7SghmgmfTMdbiizsT91CwbxU0zLugUPWBVW8E0
ZDbitWIQBxg8uNdaKWDciWkTlGpKKaYbe/EJXZCiDPlbhOS4cfR6UGkC/oKH5o+xAsXg6K020CZW
669enaPkXB7ngsVFxcNisEgLszUQwDldz9rvytz5X3D0vo2FmPqMTYrtoEX4M2tishQH7ZKfQAdx
nY7IwOrDji4FdLgcbrNVfE5aqDBq5J+uS8+Xe8JgtLLhAKaP09SKpxneFgt0NFKmjLDqiM1DPUwa
ZY1aUQqAlQYbWqbGZZR8Y0hAfizVcPJm64RYGfJaeUpeHUQeZGpQg9tQxmAWhoORWJNLeN8WTkOn
9YKdOG+7RGUJO0oFukWMYIEIbqkLmYWdwFG+VxukYuANt04qwbV+RZJxegQ9fEc0WNxSSaKt6l7w
py4Ab+Rx9ubOzugn6nAJodLjZVel6wkoLG1PbCR1YrUhK3v3qiu9m1iZNUmo0PA24T6XJ+G6Ve+H
M79dpGFMVb+Z9QSYDPrJeQiLvsE9q30GBc0ijzRpjQQ4mSxnGLV2TkAOTUvY0hQpUH0pja/U+ibk
xFGHijNCfbpkniou5RvQ1Kpnp30reU/Idzhza4cGK6XmX7Ple+Yo7A1M14RuR96tR1vjSsovCCG4
SAEEOgZll+bHv4DXjyJIJCIbayjzTOyTGhE5PM3xkLbo2ToooV0LuORs4B3LVjOIqiTcxHWnFRga
xIkPw+dELLQsG/WcW4MrZN6dMkcUa6Q/ldwJ/6q3Jm/mgpe0iKRyX6BC16Y9X/3FWALMBaargNI+
5BJ+HbQyre6N4LQ0gmj3JMENJpwJ5xlBru8Bh7FWUQAIsXBEy8fTBw94FS5dfv1ErzoU94cz2dV+
d0vAhCwO9x6OLASewyuD3JplW12FcfODBD0QcEIYCqzFAqaXTypEjg8F64JugLCxB6BJ1q7JbCpS
QoKmJkg+uhaKp9aouY7rM397tgGXAzhDkI7IxQK9H1FxV3EuRBcTXLDFHob1wcV23MCB4aK025tf
hHwoUYFtYEVzMON0xaTAYvexFY9db2ZlpEKoxsJEnrzqMvSLnBf/NFZ+u04JeGlZm8uJwoCplkr5
vbTB85HciTuxRF9UfIg/eETshJMW9lwcI7RmGf6BV8jy9hspANhqGeWVecSai4k59o0QsoMngTCo
g3UmW1zFznzkY8faZMwcEJt0cOA9f0apT2W7nX+oGNLoSVyytA01CbZ9XCixAX4gV3xtszyp/yb2
kvPU1LxyErbbIhIT/g4+5QmkS5CPQ6YfmLm0bmJXmrsk1wI+ohvdnLxW0gXevqNw7dSyzVAutLbC
xYJePl3Znl825BnrsVM7XN2+vkhAardgBs5pZ3oBXItf0LyFmkCUG3UvjkR4HOOV3xSKRb930RqN
GHepvfhfUzUPSd+DMpECrXhl1taxP1oWrddvIebsFWHtRBG9Sn+BkDdapRVthDdZIDZ81L1PUrQg
lpzOhF58A2Y1YSELzyEy840OofN0u+hEV2/e9CLIOvMWwlrDp/JsTqFDMCLpCiJiqPKlUa9cjjQV
CsUyMMuCqvObPnowYXGnM8Cke4McVz57kaoPAHSYq9kIST+bVbi8T0h4fGGpF1llvZsH3zYZl72j
vIZQ5UUbQ+87wkxRryJtSu3LCj8K6Xw6JHiAhagHTMcUamh3hmiNrmbu+ZLF7GjdXiwonZu5K1Fx
R1yC3kucdpj4Y2AJUFITlcLxWbckt9GbanKapzmx8/2xRGlkqru3uYdjSMcw08HVd6cHa8amNaRO
natST1WWIZ1qFHfuGCKAaCYCJuJ18mkBG869HhuHqXdaIb0cj0XCqhW8S5F++rmv85VyvylLJs4/
Fc3gFskMjSJn8F7x7I2fk6cqdKSGtIXGUXg0Rd0UDC6RzXXEb8C70AIBTpSvDOBCzgkxi+gnIHrc
e6iNuQvuKvDDemhaudGZ8fhKtKMS5kHPDn1/y3ppOvaFdTqL/6j/hvsnBjU8P0LcA9slSo6QDuMi
fBs+3tiD5qS6RqffVl6JA58M1vnLIrBmoe7WQlokvh6hrAFz6TI0uK5h7JkfQn72ybc+nty7D5J6
CJAFI4bi8MCB/UHhHx0l2Jy6CFbVscS4ruP0R12U77qElkEpTRG89LWGmnOk394qT0IemYtOlVOT
7MoRIDOtC9TzsqfRWQ1PZtJ3jozGuVCCj+YYFqdm49DSokv46AAQRR21xkm71IIvu+4uk8vOJLxg
vyyYKUn422r2LkY0P2nwDfXxQX1K4EhAgDaJZK7IcZwFcDYvT2/C0PztMeEZo6iaDhV8JivcWzIr
nwf37BCVEsexy7Iddqq6T0ni/hTAMlZdMGaMfGaor37K9HeXS/DKW2Cwr8oHbsus6JXo9wfpVaIo
pF2p41lQQUtQL5IDjdrR5czIK5N1HChUCC1zph6i2+P0j2W0zvmKxXUAtxMUSlbzSK11nYe4KZjO
Hgeduss+YQprU8FXuxaE6kRt7G1w2Y6e8r2aao5s533a13HvYx3+bgimJ0oW1RL5ffbxqTprfuqV
HxMQ6zY8bK6hgDyPz6MQWk+1Unky5bb3pBhJD+M8kJMgWpNWiVdvbrKkxJcoo0FfnRLZs77FF4tG
m1oXhD6lfvJdNukuY/3kE39Fd/ALUCkFl7um3da9dXLTt0BE9HDsXNPW4BmS1PwoVIoOrHTzPlsW
rHF5RiFcbtdFwE5mYia+4yXBl+GGVDGLBL4DsIXtT6SspoB1+Jqyls5etyU8rT8o00HJrQVCSjQk
I4ye9pyJEGmzoeXfUQHfQ4KXoCy3pehG+LKeogi08AegaG6HFvl/7R2wi/28JvaSpKrFFne56d+L
Dg2Q3ncbO9H0GOnBxBzuBfkBGvnULH7c++Cucq7+0E9W+0YivQ+vCt9u4GGdrLtBVZrA6eMNsO7z
zQPvYZ7vDjoxaQxgRGmsAJPqLetbKlkK19qv0o/SFgCH8PqJHol+AOeDrwSQ2Unmcx7IHxAjFfAR
jtVhXF9D3B6jOLpU4yhH1DHBUnZDgoVKabbqngrzNoFVZQmx6Yei/Tsa+Z8c8KwsnZdd9f1eCX19
9IwmuI24lFfqVqPAHs2qUPAy3bm7fYdqtdYghZWj0eJ9zMWTKiLnyPaVB6xlHV5wDifINLPZSfO6
yIOQx8y3UY89s/xvryuWZHTieNsB551noqkmzLNSF52sTF+2jp6hqIBxf5EClaJXDg2a7S3KV1M/
qtFFgVNRog3FBD0j9Zq1Q8T4PXGOXPTb/QLjLtIgg5EuxoEc9iRdyGu47TKVuQsAWj/i3tmT3Lw1
hJNKX8CZ7zi/eisBpKQV2iOXU7pyexlYEfnyVFIJwt1wel3TCQ/8G9OvG8DNOZl2ShY+AgPU6FLT
mLH0Plod1nTCbvM1sBiinEr1BerJf6UsiNy8op9crwMN5ZD+gIxOUSrdjdw5v7wSxM6B9E/M3iqk
yCLpKCNAhsBxxxV5LAS9KKTospmpa2HdHaudowv8gvZtuPwy71HTqMko3laNSRDc+C/cVA9vNi/+
/BalpDv6Iq/aFMx6TdeArop3aaJ8P3+1758J4dQVAgmp4FvYV/cA4l3EKMI0+SsAGKrnoNSw8Aar
wlb2s5j4T1ps+4xdRuU4YzWpJF1zo8SfCIQmTLzWy2cfXJnhwScWCzx00Hm7BAHJJ3Z9pCbNXn/A
uU8O4PCsJVSTxY3fkaB30ua0M45RnIgysiKgtI5I3Rs6pwd2yCVKGMfSXrsFHZZsnp9TH4h3mmwU
4eVQXl0U4DlKLAglMrVa3YkyJpFPn2QNNhDv8EFYTZ5iIx/Ffwuc3Yam8LryWhfyy/tplwHY/HMU
J0rEhcV9tVii6HfZ2l/9+l8e2dH2TN0G/wn6w/pY1G5ZV5vaEZJE1VLYCUiaCZyjkiHtqu0+cNh7
Ej9CUe2SheAfPNK1S7Bh9chGAH0i3B5nuYs24CwuIf1ZE0WJ0bRHlwZf3k/of7q7DKhO3mptKYHq
Ym6zukvsD1P79man/uQ9RDcYswhHnjRn1Xijfz6rSo68IOA2/S/0gdCBZVgw+RlPPqs7ivNd4wGs
aZz3/z4751NoZmQWOFLOKbXuRQ65vqg114TCeL62QH9vGbrBhz0URuVmmI8YkT3bfOFcHE5brFtW
PWyKWQns7MbcOla/s+TA6XPed9nZkwJO8nOakWG9jRMFwpReAIox5fADh6gtoo64xJQrIEBUuyMz
x7JKsxQHEKuNabtHlb5s1f1Nr4lQ9rEAsTxnpXj51Bq8IK9zFCKvvV/RUkuve2cbv9+7fuhZ0WB3
LGVQS1fFHIGU0Wc3OqzteedBEYgu31vLOWRJkrhlj9XjK9JN1Hpm2Q4yolXYp7KZGbRGjdjGWJcU
hKF2HAJXjNwiTtLwcGDGa8yL8bwDQ+Nl7x6b7zq0h5w+n4RlDe9xywhhQ2xLYCE4iaqdWmBNtkhN
zigkRgJ46D2bud2x6zLDXWoUUALtzR4tyoiL/cGlro5aBxeskVgmUbUYzOxijh89sxQag6+5fseX
hkA52k68IVZyEyIud2DKHQt5rZhYwx6/EEhnVVPqvnA1PvPn1asjzg1JQiLjqvG4p7zGgwhzmOKz
0VB0Di2adRI7Sg0TDubsG3q+tAIhhs1ao++1kZS3Qw/eFYNG81gTAQANVsC/BBFRy30kchGmQbEn
k4s5Y1BWFUxo6XTM/eSC8rlVJqAjKLoBFE8BvxdxNFRCojfAcdo1daopz6RfBRm2HljhOR0f+SaS
MUJPQ4uJKt9yTzekF0m8o6ETwwpSiPijdtF2hMHDFoV4bn8ZnP8+dQX7BBHajiu+scaLo+WewLOw
3kz22xWXq/4BqLJZvNdQ4TtYA6dF883TjGqrTN1PnyyhMw3F+821dpaTj/aa11Jj+mMRcJzb2I1D
DKtGvUyyhkLQQRDoiACHkYhxfUYd6hKjfMQ/tOUcWnK6FJqmdiOtbapvMzEDtotCL08Ad2vg04Ax
bos+iDnbSdiDeM8RX6AmLNkVjbcD6TRx/D1N71K1rNHJGABSCuRh8YD6JsCZRN734t2ErTz/Iehl
bbbdt2mxSdjHH13ph5BkpmIa8ST1R+qu/HT3kDLR0A3RjHlQ0FaPEvDDFleyeHJTVVtrITaO/DYt
m+JScFf1ldLl6QaVWyEQXSOckqbqsGFUXUFx6+0OdE8DtdOaDMnXcpTqIqX55eR7OJCM+phjyts5
TAbXMoBWewPrelraoyh0aQUIsetuBcM/xV/7hC5BGsxlzzOSLnvpNN2b9uNN6RXud6dP3bLzNHcB
O44BISZYfUM2KFIBwgNK+qmsaSYbIHBMq5nSF5i3o3ykTEAO6H0Tbc3/yAvMLX+2C9nC+fo6wwm7
uY+0D41uKrDmZGkIim2VqxcjlkzZ67CRfEKr4Cd3xys1e88Lf7f/ZN+1Q/C9yX08HjMKoPofYO65
7rFx5TjhbPlEcK9rDIpg8i+mhRMpBaGWb7P7y0RZ58hD3kNHciffCGUFbLDxRufeEqOjhxFdbnD+
ePrLg7IqPxBh73LBH7Rb6PnuChse/3rSu+RGkeLcDa79fC0iIeqj9R5QaPg1QNez1Dxruaju6V1F
Lpuwr1xHolIFFKMumUtEx20uetUvXm34pMUeR/Dj4pLhod3MvS8EF06RXzBWajPVjRAtY45yYdS5
Yt1nND282Qvej2D+rEkq1euXUBiOeQApLIjwE3L2kYrWyaorhzg13cHNRC4a/F7FtEgrHuOvvOgh
H1Vns3xKHHP4kJJTT2trseWbJLTQVVdFJyNI0criqZNfdNVxSetjHOsSD5TwFQiF7zN/jTNnvABo
AuAecmuGfCA+oy+PjiRcxaeFbvSLpdadneslGExxVvkj2KQi0NIq21cSqhjRRNwG27buojiPpFjN
3N4Dk1+a57TS6njp29TQtlxtH5K0V60tIeRrVzBzc7FwOXUYLhFOMYo94Klpl7dWzVHi3b+46giW
kPCMG2s0effwvMXwkPwcT2wDAFVev3x7TmIZObntF/OARt1nJOGEdMrrh25xaSs4kBEzXoCKr5aA
veezmjtME6lmCpuxySTAPyCcsWWZaQhQCju4DqvHyHEyLLgadMlyz9mOPmWJhsJ1X3uHAslj2SBK
g4qe5Zm8T7aoE26DF5a507u4nyQq2fWKNWqqFXK4sNJaAR05C8lPv0F0F5a2071ZvwdE2WJzgBXe
HvKEwCaqZ80bmXle/p1rkjAX944+Y8IIac/HJzhjLVcdrLFaGYt0eDUMwo1XMqMrHK2X8qmxjwhk
XMTpI+P6DyP5XQCnlxhZ2iDPOF7cAGwi+lQJl8HbzI39IOzBzZy2Jzh+HjCNjg7JS7uVLzQh1DOd
G9vOi2xbNVhSLh/zxtIUXFsJ/rkknegUY1hMCmAd6AHpCkJpv6jxVel/ZtfymVZfANM70OPrIBKh
c6WLkYrI3q3zoeRmZ979D1Zs8Ri0NvhNMtzR+DcPW3DXpCHLd452qDAYEJPI5Osf3B+362LdKnVp
tkYCIg+JVBxUFAe65eJvdNQQByBGe9G5LdhaYAixvudxfsw5ZZMrhOOEawkjxcrsMU38AJcpAIkK
zUE7UIr7U9wnmQZLVRe7z8iQKrJFa/DOw4ZifcKzLv4JBSA7VEnqR28ts2VuuRXn7btYMXbvQ1tS
JDIC/Q4DEszTY/B538fjZoVfIMNOi5Wl902nDVRc7nCqwQPpwl45tyoC6Qbc7HUuBQ4x3CVKdrWA
4f+jpcH+nqgVveq31rEpVKCV3rRpBhYraJX6ksEn/COIUHLkB7Hrmo3Mn2qRbUZEObN9JGAldU1g
BDmVd25zYLB1/x7dDnDtx2/mr6RPm47SJDW93H6tPT2NHwiGM3A+wBW6n6Mw0H7MwIb53GSa4hod
/PKM/0JpBBic2qPrYqJonJ6jKt/Dy8le5RT8nl0UWlwoauF8DnBAxJlyxxs0dYejpOSeJx9k0Vy1
Hfn5QfP9YIYZrNYCO3M7Yx31Lu7nQyrVExuTIq1i5XoYoToW9sTC3Xu+9TpY4SqP2g04d/KoDNx6
zd0m5jBW9oBNR/wxLMGfBP6K5SXJeazFOuT8+b1nu7AoT6/ne2RyyLWpYAcdbU0TJQnkRH/v9OpK
fB4ipW7fite8JzXPMHPE/WEV2xzjJjIgezFVON7+YQkQ2a6PeAx9XEwBTtfeMMx/RHQDeBDRiKFp
8SKAmqE89Zkn3QaoAu6PFLX1wq307hZz+WiF/OzC60/L7UHDeBkP5ehQq7YsoH79ZIUofxG5X3Z1
wSKb+LkpjKjI2DqCaSXoSgwXCdDUA6DoLBnhO4Gkvr+4Wp1aH5BF+8BIsSIGn8RIoQMaX+m1F+zV
xRruKI7G16WGPiM9N+7Pgx4AF/ftoFzrV4rweJMN80LJq+2xN+U8l0H9/uMrfsspVyissvk6IZlx
0/yePO3G8Y0sIVEidvE5c9EIvqZ3s7oiw6oTt8MgVfWWxqS24YOTdMPnLUdCJ2UhICasz6Ug6BqS
WhBuKMdgN0/k1WIdQPFW8CImqEzOsUyOSYaqneyIusldGDtwhK6WkathD9S2bLPQkm5CFy2NP7d2
MHrXFrtEAX4+kJIt4fM0u0JxEFyXHKFEAzdinnHUhWjj7ECeu9owHC3J1GS44/l2eELHP9hXklhk
LFYmk4/3Ubpz7LhhSalo6hmI7PJ5FbHH+WqXbjmOsyJueg50ygtrRIFDJ9G9Yg525boCRT43zUNd
NFSULgjtQ1ZOyG7waKyyx8macZ/2IdBOgMamHHpWuLOZhSWuteIG6w1QYb/hFzup7zsCJP/KMUa4
V01prC1MuOlDUT/xp5zB7qu5pecq19oqy4PjfcVTCXyrpulPhmhhc09aECUZhvtRsXxJmp3u6G+A
o/ZBhfq5L6+T738VDmWdI3u5iKiDMnHHZONk3qgq3apSbxsrf9iuOwOzodNW/HpI3q8EkCwd3dsY
TEpVtVmP6viFQnQaViOPDj0Tk18o7Prb481k2qNSbhTOutesarNXsJaLxRcCo/IjM+3j7gritSSb
STB7b8nd+MMny3D6aOtawK/38DVgF4VghyZO12+T/BkUQR+0KRF6h14lmI/9dt3YnPpyREgEwl0A
LSmGP7I/fbb8NxX1jMx4LW7SCZpgZgHlP9I8xxK04Oc8qXYF0KRIDLwClXk0DYRIru3AdGQVS38S
KhKbl9lejePMvZ9O5am46QVRcOGgy9oOC8uoYhfP1pgFVrrLu5964jJZw3OXxUcfqgR/NREjIo++
mv/E7uhBjvyPVeDZ/IojLKLy2XRmwI/HBPtpDWBgijkCTJiKuhmoJdP0Rtdk0KpY/HRzUZQ3A+yS
AFDEJKnpuxFJJr8iOzfPxebR6zpHECKNHgVeHWkPqZg1fmuPuHQWHlCJ8hMivAgIVWMKC9ZMb1TG
nKFbs9CLVH+b2D5cUml8ahybw3yPeSX3msLO4risXMKmz8SaWZuWqivrYwK1rHksqXKbZKSnWG/l
kclxNq1ueDK+Unk+Npv55Xel6oEdATDnRokNNfZLx5L0MNi/lGi31jBGzlL8z39rxVce8PbRu40E
+7V5KPuG+YKDhJVvr4iMarc6DagBQ37XEh5uWFUDWf2mqM1uN6lXTuV1NkhFQEetqHppL5Z0BLc3
npwUua1yU1uHGtsRsD6dY0taRWtxSgrxrz6EWwz7i0Rl4vBBkF8aM1PooTtT3fLPmyeu8si16FhT
fmae5Tc1jpEZfXkanP1bxvhXZfWZNqXa9CyilwVMFUttLyISwrW/GYHMcroWfWtY4KP/cOoqy7Se
Lqv9bR6c6LCXVYVUp0tYnhyPM8pgT1f4tPrGJ6GTZYjn+DWSRi5jQNjH5w+o/DNwALlJTOjgIAuj
8VjkdJy90ITH9u2QABTT06gJNMTDH0Bbwr0G1F+ThafeTXoFE8GFGezMD2a3tD1w5OlkHLtYrd81
15U0vLTWOg2df/u33SumT9co6RFQCtOtGyKhWk/yBhjf7NWGBa5O1v7ceCrIWI+sdigvJ3QCbkY1
U3BQYhXOMYVcA8zH8AbbF/FRoh5mLDjZiI/RPf6oZHaOJqlUJTph5zpVd7YwGkxuISDVSuXT55rI
NyDwd+8h3onxjbgRCNH1BZ20KSYt5DGW3q5dWIWYRWaSs+CVebKl8RfJMNVQTpTw6EnKDe7SV6uK
r85C5o9YGySV0E2hfDJCLXdJVzLUKp3a+9Vncvn9QuKqPvpftoCqayqW/xahA6GwS2OlTpde6ihq
UZuoOs2GncAQiyAHmY/lEGVfO+61SoCLZBx7BIvNsgVfLC6q2YJuO8g+wuxv8vuMuQcuiYnMGffv
0Wp3dc21mdN0xaAcUPhpDP/bWTLaI3cBphpW9f0SiWIbs5Awcdp34m7V3WtIhL4TWGjaj+aTVo3v
1Xt9fYWmHfAMhHvCc6h2l9dwYL7QLNJLZJiA+RyDh+94m76rWpT9ybzmhJfBDToLdGs9RA8ees1r
jPHFQWcZY3SUE/lQdDGkSadBQW8fXJFHcLtdorzSkOlkvdFgeAesjJVIAC5DZ9dNDEYYmj5HUXpP
MWZBdpyqy5O9Y6TayKyKxSlQqeiReS00lBzuqKBIZGvOeMcauVPHXT+gDE2RJUlq45rZQpWbvXoH
rc9fzwJCZd9CJF69uJkBJlnde4UehTvX25IF1qegiMaEaT6ma2t2HUdBVlaW7fQnh+NbrOQKnRk2
QaA0ilSp+bjiIlx/z03K/X+l/DOa75amgTxzeGf4AX4ZAeWY//hYPL+1Sls/0Ueu7sdkkB/ybIVZ
BQ1wgUny+nCe0ApMw4cT6aWo+5W3yZfFXnpJxqqc+ncVf5h3BuDOuiBafZTlc6SfFGip7eOoELaJ
qa2MkwS75z897sdBlTDQx1Mz7XHCz2Zr+G4D+TmDkWM8TgwxsaiqN2GQP0RC1+GFt2OznmBewDtP
uPcVtBF0rx7ZQr2hc5B/2Z9fjMThojItCPx120INa9SXCS5RGI31tADO69sT+R+XmZtY2ubr41Si
rleXkXze0q7atXml1oXZl5NKuVDEXmPMAi4I3Xg0k04fVB3Lw1pvjGofDTdxoNCdcqQHLwp4JERK
w7IQw3TerFL6oCZNQV6OCElUVRgQgWhruAME76cbtiYc57GsXFfJrEjgnSrp42JeQuZGPuKvva+A
/foh0714lzqXZ+ovD6kzqfkn9vs6rrAWTmxMlMzmQEu87UQi214MqnQhq9jrpPtYnwPUQlcyoxQf
NzQZtqEGrEoYW5voATKhwydrjRwRLPcVl66Dc4qRFwHKGE0pcgHoKQM/J3X4qoFnOzXS8jElUyhq
l97DmShgujKPW4S+pKkJpwfOdjdzipI7b7wrt+ZMQl6O0GVmFILv6oG5oUx/BgGZPc1THeSUVrBg
XuMbam+iX32RyUue6/JzUvYx/L2UBNHiCTzfH4LdL0yemWHkdxLn4emFF7gD7OYiGJdKldys7XxS
vUfPAUB+4AuyVM/QcmJEMH8kywNkkcIXJspU1ZoYAk8D2v5hE6Sv9wxNrNjTZXzmZul3/I7l2wId
ug1CEsP7+8FWsz04Cy3viF3G7ah8NmhOFmUnwaoJ2zbaTVKUs7kxI5h6m1Eu3Fvn9DIXtCvkDQRQ
Kg4wCjC/Lom7/ucd2oisvAgeOGu7/T88Q90wkXMnVfU/XwkclDSXlM74nf/O/CdqLaPxCAwo+40I
uBePH05T+nk34KKdREE4aVcfkHCbFjUcVjmTp5P1JhYTycgCuBYQnTLzj207Jfe15ZWQeJi2+N/F
Zi9TKIESdrkzPsHqXYwGdp4trYpMkyFGbAZJubM8H5cpUhmzoA54rjbl6lZfnEGRMQ7M74TMuGMC
5CkTCambdef/B0ykxD+b/mflHOuE7m+AtaxhViQqVlsfDuTzVAjJkhKgT4aTPT5nTszftdM8dqtP
sJJcAKIyTzCWoKRV+gKW2M21yytZUJ+MKb3X5enj+uKc7AHafALdKQKC31CHfKWky0m+p9P8dcK8
Ko4JsCpmUKrw3oPOztDMHy9HpjTkj7mr3ZeeYqkxdbDm4J9GaZFGYDBFldMSoGa/Vyp0UtjY/BOC
xoRZewqXU/BDjdyTadWQu378XRGHvM8aPXK0f77YXz463PUW2kurNuYphwIk0Fdl2oQLCWt/bld9
y0WYUrPj5kGOx/r+mkBdzxjOAngsXBTdQbfZgs4ikhvwz2NOtNFqdcH/MAPE+kBYvvuyKaR/NqjI
PMCBPei7QZ0Y9tiSTSAhawKKSBI8ChVYNyvNzD9jADYW31OqZr1wtozQp+H+0S2JEi8UDxGArDed
c3JUjIbn54WKWcHLAse3mjg3jvg7ZMD6BhVGXKOTcYAu0kYUG6RpRb7GmdcVlMycGSWpxU6TLPe7
6cIK7OUek/GuUuReMYoqloLVYmnr/CffJvo6bS/RGrZ6stpTRtAQubpba2YFgK9gPJJG+QhUlWdo
8BIo3mxw2K7G4DvVhEXcb2wz8AOvyGou7dwhoimnCI/9NA6itsVv8YsVPAUwjJR7FD+FVz5NgcUB
ozYbrVDfr+G1wKWJG1gEmKVl5/trmkylMbki3v2A4x+kFWYK11W78NrfS0O80PA2SStM9is6l1Q4
Jl0N321GLHcEbu+MkAGsaZg3+JEtJUQGD7vHl0dupCvEQw+EVA0HG5xAdOCEeKqN6aFKL95R7BhF
YGt7/4uZ/xa8o2eGyexSXNBvrwlifs+jQUz1EiA7vbpsFm/N2vuqsL5eppBUXqLStrMKN4dfqGwZ
FVrHmi025BUDOgS/Nlwz9qRZEY+bq7OUE/ZtxdPjFAX0jMhWzzA4XCGgrmPguOmELp/xFVpzHyDs
ms+cVNqmmDIbQp36PbufDUIV4gBobyOHSonXIrSCs7KZ0gDDjNBTkFQNqqmuOSztfQ5WL5UZmJhR
VLzOlfkIJ5c6svRCrzLDqUsbQptmp0uKkVzE7a9/z8NKMQLNVuuKTqbuCl5FgjY+lcKdd3sTVJ7X
cM9Trxk8v3xh6DayMa0V0tsC/YOTVVj0u28vUnD0ZbNKC8PfGNwUBCao6xTZ/rUnLSaeROKQc47j
vQNK9VI3mnk8rxPCnFSIrcEKKv4m5EyiyIQzlcNwcDIrfTzmEjzu8qWYnsC+4LHmACrts/CV9e90
PS959gitruJE/cQ4X57q80YdmWy3jd4y/S06lLQvO8wdtyqh+dcHiPDEUbjmp8b29V0FKcISSRu5
xwhSiAi8m9+nqs9j+LBKWf6oImv9kb/7LRjlt8EEA6prLh7zLNwJ+UYN7u5e+xo6ysuwtc8SFWCR
aJjSlJid8G5dOzlOrSTCM8nE+jto3aCewChc5LlqmLgpcaHmD6D2Y9JGXAGb3r9WkF95aXF8eMs8
2beAI2KFKMfh+P+MVBELMnwoR1+9ENUoF9ReiDRDP+ZRxOovRV5+jmwyGJ12NzM7qH88qzuxMfA0
CDOhS5proA93Pdbw2b4tO8FCH6XVmks1O6gRWBhGKxPRuKg9+RpnunZOjnfTHfV8EduHgrPIZ4uB
WRR+vUG3bgWkb0jea2i7Qm3Z3p8wAcrPtyVtZ+gfbKpD7Dnr5yT6vhUb0GbctebRYfbiQ8qws9iz
3qN1EN092JUuP2o3AN7/53S+rSm2VBaP+jX5qMuDoDcQ0r8BupDH4LAPJGQNaLs8aVpdXhW1Pukn
yqZrh7SNb5zxA0fsu/yfkUnlpfyiZ4BKrcw6O33JLgfVGjyYecvGj98Io9jarEqXpjiJHfpVcu+o
fhktDh/1yKxARwV7/Ewz/oO8BJcIVvCzycj5BnT0jNgEC7TIpCktD2RooHfyk4huEGdIghOds2N/
mKAF8P4UcGbZdVG8e/CodxuQtopeRA0lPFRo3TlhbqzbNpHzo+dmMp5akbOw0YY22z4nA5c1zVRV
CUSOr5gUyXDEVd8vbNzTFpxzIil+l/KSpPpPj8cYaAuZi4d1m/6LVO367YxQDyE/Z4iPtI9/QGmC
NQNEY9Es7Z2jsad+oq8LUt0qsEqYgb6m+vwlbNEXK/Y9QsWfOH/+M7qZgfxpGz4v34X60iRD+1Lm
wMa+C0JEf+548JWb2qghozNAPs9LXqdZ7FLO292RQ8jIFVawXu6y4xWPDMJ5FJHTXeaYRsP9opDW
UN5PLUmJiNW05RFMODoQoayQ1yWYL1A0dBg+C9buNglfG8/+qLoVOZjEquu38ymoCEDHiM85atr+
GN+lbRJWiH5nbHJqkKTXxDBCAAEdbpXcFtyFcqMy9AUdONYWncJJqESS/ux+pkIaWt5ygh1DBJEm
sDkDF4R9TN2YVaFMmHv28FMEEh/DujBpwq+FJYp8+BejzIs7NtiwQLW075XbWweuQPFAseqdmAwl
uFVT809EHlVgbWs9Un0NEX9hPFzN59cTbnmwdecqcIvvkQ2H3DdZH19qWNkfZWB9fz5tkHQDmeAg
/nVtGaS6F0m48JwsRQz98VvaghpW+LTALmeCdJeub3KltQwqTJNtaDHfqv9/E0w/dJJD5tHr0Qpc
0CGRqvZC32Wrnp/X2cgVr/j1CLJWtyUqQq5hAb5aov6jZaBYLIQUgKOTlWr0ow5MwrYFubjDoUeF
WZKUfu8iafINDEusXG/GmlMFejn5vRsPCyzWjgG+aYDgQx8B5FTFrrGpuAQQjuNHfoS2nL1uWJes
SiohpDq6Xtd/Hkt8r+mP+NzgDYdVDVft9hz4MDIAGyMVMdjbaL6F0+V37P3A/GUVqdXfjNB2kEVV
2uqdwvzqdT4puXbimwn4/uA08MRU8Rl26/QXX0uZGQvl2yb132GcoGUEjfArnxR2TIlU5+smXZxm
V6BjoJ7gAHnBqzl23hRwbgO/dAbMp1mVvGT238BbTCpaE7NWwmYL9VQi5SEa/Aej6QCTr0j549uU
vT7riw12gkDGtkd56n+N/MjxVBusCb5PKjRfZ7A0K040Gdg2ibR5tgy+dVFZrAzTL0BLk4jomWMT
gwQrvgNfRPhVYzwpV6WAbPpD+EbBxLIf15++vxgSBZGlZemgvq6Ovz/G8nUD5HCmmbICtg8zLLsR
V9mcQ1dBiPY9naWJrJb2oUNlknrcE+nGiRT4i5rpla6I53H5o0g7T7xfm8scbQ6+CYu8KiBnJyYh
nKNYBA3SePsg1Zb80v2NWBmOtP9ngS4Jnnn6NfhrDPFg+ZcIQYCiYoC/QGs1sZu34wWuIyvJIFxN
ATTYVffxytlvsXYid1IufmLvHJu7pQyI/yddMAAqy86ms8crniwcfMZ1K1ByfIh6bdLYD+lr1KQ8
6cbt4ttBFP2zxt1EqC5zrJ3/Uk/J4Sali8X8a5+fIETQltnR1bp1OIdYIoBlU4wG3BX02GTP77jZ
id6/I+35W7V2K4G9O5IvZZ7KwDYtRcM6lmVbs4tIErrqTL+jpOAEEWDDRp7oPqUzjxJgT05hMSv5
h/9juF43xHbzFxhBYyWeCu2PMbkdK4eq8SnnMIE2angpI0b+sCPn66DKxGEmheWk13Ig+SLWZCi4
1RhivldwUTZDax232FPLL4w6qN/u3kFCoBQJbSQ9fvxXtLdeqAtZ8k65hVCXfA/H1wEvDH1aT0e1
IM/GZEhkolTrBDuvdg/cj3yahlmK2b2oGTLso2vGtcZ43WPOdYvVqts7gnS2d7FU9pHNz1TpUXCG
dA8nWFprNvZ3EZpchwu/Js/w7VOuSH5cYFAmqyzVZ6vOuM5/vguMkIo/+rf0KEkvSIi1aPnJSrFb
FD+JVodue++x8jT9O7pbhGqa/LENy9BtlwPmEFiKxvuvscafzDAc9X3AcXX0CRtf4SnNvTjVx5cd
cttBTFtUsNp3kvZCyWEvqllj6IHJxKQEj2uPXBMfNssZvLVnZZalx1z/raUihyTZr9zjvZOB0wKc
IsBUBnNc++BuwFOHoyrywPT5vJceCkFSF0ozZUzmrTpSzTlKz6wG8lrjYOPYdLciVub/T8M54D97
soZonnDR0x7FFI9R+JHxoJfRlqMSHbB9sfBiHVI7Nbbr1SiL45UWZ4zCaoNATuIRYzio4o2Pqy4t
3cbpnI2WYieW1Y0pc7+Cc6YhTp6dvMX9g1ySUW626Uo/RmlXQXYNeQi56sbL4gHslgBlC89STtdP
CtBcxI5akOS3RWH3uNoEnlApbadwPfNFgn58DoXULXTWuHQEClUv9xpb25jX7EX+wl5V5G36a6jz
KvkuK0Wqim33PC1GnZ3mr4xj468/rrU4DEMaWb/MPXlaM1DXg+q5MJhPKuqoCtpaFnem31FU6a2o
QjfV28UQnVvbzQnscVZWJ/5DuWaVJUQlxra95m6z2k7t4bX+r1/sahT/7O/95F5GaCGst8UmNenx
tMydkTkz1H6LdW0Qw5AMqd3cw01cHPRpDMV9hJcpsE6X2PjIGEPyoEFcXp/uxhwEO3bjt+Vh+CYE
+tA9DrZ8jXwolAW22KWjd6kFD6nXnPzy2vNSeSQcK5V8h1FUhWaqgmilNAeC6WD4B+DRfZDIgmUt
34VOigQuChc3kxJRShqBsniZcKdtLra17HGmpFbAY+CgNKGYMPXnOQCELQkGyreMg8gGIUhpdxU0
i2s66hdQA5xFuJDGj1TdDjn/W4ovSQwS9RIhODlWcwiSSMMuqhr2rXmcpro15APyKOZPzL6+JO+j
4ViuVCZaKILnO/SFj0OxQh6/Rg9Gwqw7xD8W5eZZQ0xIP1QDtMiEUnTrIXPe5QDqADqtddGNiAwn
9YAzZLrp/6nFDgHQwg1WbYYPeohCd/Q2UbrXSc4bvZnQAlp4fNsWAoFxUAaiAyqdr8DUMQLDDTvr
hDqtoHJzuzRfskYpmDu4bIzRmyl8UucCnTWWUQjeYTYRkzKl4WoOejcmGyWh1otv+MZC4Hh8Xgi7
oqU/jdjzqT/8SO8S4DcY+8mX7y9TUYUPCVbcsUKVrGFzCyDSdi137exUrZvHsS8sZfoUxHCXPcUn
GjlZH6OnPso66F2f+MDFmelHeXinHzAFbqxU/UGren05VsdH/0FV1SXxQOgH46ZO3AAWaVV2wzjI
JeVoq7S/HBo3U3C2rIEOoP1Cmc5prV9Qm/RBIL693LgvIjezvcS4QUzb9ahrizqVXI43+s1R8/xy
byp6kBg/vkdewbA3TCkckHhd9O6koYWx1+Z3ubCejAMGRj39k4C8lYzoZwgsirk7k+tFdPD3aLwb
yo53X3vt9MOju+tj2DKkm5wUXV7K1KrtgRqe30kFs/b6GMwsojGkq3hIAMW7Z42vOZ5PrBizdNsa
2aE6dTXVsczAjZtWWN/ifDSnEaZnCHNWlYHwsp6yfZTw628pFmNfWT4BY/1lPQ2pfpeUXY4kwVVl
F3hlpAafUnTGp3EBiZtOo6KFSHa8Z/1N28Wz54EnQ/R2DHvBv5Pr4gmaC1gqxJxuAAUdWFNE6A3e
Og9WKPZneyBhKqUkuZxu73Hp65KBmeNdnmiBkDsQPQ8gnL8TM6pC/DifIxkPXUEZpBt3tVfWphXF
FJSDlFZxb6Cy8mWaNPg7Xib/doP0u0gutjERqrHCzNd1mePZNxLn8iohoqfdNDEmhI/dERMH3IxR
LVBweAPFhOOsPGjyCp7d9+WahoHDsaM64/cmmj8p8lfrJE/8u5OynnTCjs/oCkUM62239EgmLwL7
BMPe2SKQX4MBZFCNL31/bIoDGKG8m9F+MGxEb1jV9PKLtPJNm2IoBXMwCPsMjAxIuQqrEc+tDkKB
2lVfv4P8PksbRPqIhXUNbw82ZZVwfLh5vF0DDOYLUa8mjfFxAdbyQErYmLgvCpzpmHApJ2hlBT5F
7O3ZUUzc7UEY5B/JpOfcytj/mbwzSsh6pLK4571vArMsUUMqflEbF5K/wjRRJ6Vh6jRmWfQqyPYG
UkIz4FmEArfnNVtcn+uZIoJ7YPG+PL0JqIa+cg6WS7mzCZbhndGNHXiII9shQ7c4/wf2UZreZIpr
OegPcsSFAilA0Bi6W2hZEOZchuBHpfXD3+t42OaIurRiossHo88wOJgM/6ibuvldxMIAHmEWK3ka
K1bkQvFL+LszCZnE6q7phuJhdv2vWzzcIkpWMjDHt0Yc5V0I7nxjsi+TOv2xTwtDKMOvy5kgQlWG
m97h3zJz5jlf2yLqWpn/5IBzUADSg9MG/70IF+6oynN6U4bFKwMKlM8ttqXYbHtAOHoD01DzjLNH
TodViqMhYNyQdiRfp+pmseL9Pn7FP0KpGSlYnQ0JxpsHT6xFBY/OXaTLA9DhRvTNYSM4qaSoUjzt
RubBoIK/Q8meiZZzWw+Ys4aMP3bt/uOFbVr590mLF74aregQI+rtAeUNiQp4t2hzddM1HRi/lu4C
D1QKd/8lMH1DhnTGqrdDtt2jFsfEdNfjewNbBBFLKsPbCnaevgUX4OtmJhTGn/C+mCM6qnmmZyDU
4YuIgqweaiBW8s0mkQJK9JYWr5MN7uX2o872emzjCrMeIOstNgNtcgZ/g6nMvMacPccWB/BjNC0d
niNccQpDjNywCaT03kLneTmLQgp/e/syNJ76dx8Pli/OCSjx5KbF/QO7kBJYlCZu6oWTtFpzAaxS
lN1GR2lNeSyXPPrajajGyQtRGNhFZGDsnABnpL21OJnK2qO2alL4oS0G9aYrjOgWte3Y412WSztO
SfWJ/7LRs56/s5ScO4PZFzvcKVH40uPycYZxs2XVpLfhkLp+ZgGufsFgi3ViFSRAjYAvzmi3AaGP
a62D5cJGuI1cLDvK9UpY9sh9gZ2ZdCKBxl2AhgH7lyitqfUkdt+QjiSu31QbeRgmplszNeJvqzJb
ICAaifE1iO1DtdVbW62SVmHQMJN37OuWVQGVr97/pwX7u+VCRjTRfQrnkYv5Q3I6VfmlGX4g5dmo
Brzmdx8T8upISQO6f4FngQMGEWJ2r6JomRA4vwO97XhtTfFhcF+N5az36BQIMcjjCN4h/a8JaYn6
4jaye4rS+xJCbla8fMYobCr+Lxhej0Xyd3nW3u4gyN55BgHfg8IA2Z2d7BOxr3bgL6HjcSjJQHEe
xHI9l23v1agDLyio12UH2Facioqt2rJtDzpddMX3xHVxWKVvXgTPXEWG6fFAEbYy9ywkNi/hzUHb
sdd6mIgpHEzdHR+5eL5TKk8LdO3HfCzOo4KAaWfERrUb3hM1CGJ7neRbUc6AhBc4xG+6OcmNwszt
Gg/55kwAt+K+HT8K2jqfzluCO5GwisxF4bszhHMY11YO0ktreCUb+xfILbCmHyXSNQQgQydufpfO
Vb7GYgOoTeeI9XaX3pafPRHjgUqHKhDPoQlK8q7AqgmNfKgXAfAtBlcOqmhrSmEURZ3ZLh41UYqo
ugvw+84zdOevCA3LiL0+q8kvYDd9afcE2u66nqPfPVH6qNEndzc9ueaw4gIcbZyuMYOTCXcUdYgg
kfdKilPbKZRTN/XPL93FA1RG91sL4+YmmTmjqox9FoazlC38bS8YYp9Z7U0moKFexpM9rItmkeen
oUCe9N22BVyI5NW/BRTQXo5w6l+I+AYkJOSGl8yQPnnhPvMqgGTyRRlZ4m/Kihbwq6hJHu6ocbSv
uYR7Rv+8Nc0dLshC/EuQgSoEWtO+DbTGxQGBDiaSwVQgugI0XLJxEIBfqz99r0CI91ARW8S9ILTC
BXmFlc4Tk7bJM/Os7L+HVG7CBOAmNmqs1qspXvxiNyoeNHGZjOzIfQ2TLFltKq2Un2PvfKmXT0XD
iAYy9VXt44folA5+FNiOBUlk74GpX/6kbF7n+P/aL3Sa/+7tOP57sJ0Yyp+bZF2oE8FUsODbP9BY
Y++7TEl1Te3hxGUyD8lHr6DWSgVSWtK68BA8O4lI75JadEx56El67B5tm26ekEpfwWk93xZQWkP7
6fj9zjbNtmIjwpPCkAxvNkg1Fiqv0tBZwUnM2OddRGm83aOy9UhgWektDeB41R1Q8U5/VQ5HrAHK
rLFXZW0zyWvrotx28Q4uLGveeE2mt/zhCyntzq1rx3k2hx6hF3sdpLHCEfF7Xv9Q3InN6XzNhK5e
bPgfClsdV34C7DjfW/aaVcqZk3NOSuc413dgVd0jPpeWtM9FbDczgTeoVHRU8MAFSWPfInSrT+MY
ESuR4RTLEsjCMZE7itMpwhpiF/H6+mbSmPUvq5UDzrqA1idF5iOj2Kjk74M+0N4mhugh/PVZNW6p
VwSd1zfaFAlT6Cju+DbgRY58CwRvBs8IY6jgRIWEpCQ3x82wDUXHIR4U/rI8ThzlLvq7ZTc0yZUj
yeASElXvXRGXNbOxR/czc5yR3t9TfX5FOo0wfAvbYyPBatvg8yKkPVV7/ohqvdB7oFX8HsmC+sbG
ko7fzzb1dumvDf19BBNDgjHA6Dtnwo6v2vz2hXBI6g4iMezVojn6Dr9URdk9vfN0b2VcXC37YPAs
mtHz9/RPa+nIpnfJG5yqXWqUGA/Cvz3iDAMI/mjONdY4R+uIJOMdJyY6d/lM0afK7uw+cFxgDEVh
LyKNNfvIVUCigF/t650k3E+IOkSrX0y+JDn0z1KLiyy/FwoaCPNlEI4Ow9RjNFv4mSUZmdv9pT4D
HOHoqwYanWOTQXKAOeAemJZqBcZvxhM53tJCcYA4cLFxXI2rTMQ5ZZXPV8N1z3z2AUMr6s0lSeNp
wxcYhZBGC2ktAKWKhjOjD6EfqcabQG1DIto2R7TTpXX1cs+0Uze3AdQbFi/csUmj/5sDLAX0BZdW
VbiZmI2glXq+uj1OOn4G8lqT8zwegp5SGMlrDldiIdqfDWkr2uUrCc34hduL5DM+jd8da0JgJdJQ
4RqSa0oc20GRrV0whKOf/dsXEuNlI+Hd7yOWWel6D6PlRW7wMWtxp46jbXyEBdecjVb823tVeH28
gH39H55ySSG9XgH+XDpbJw/anF5ETgS50rlJxzYe7NoZ52wq/YfdX4GqT0/9UH46k+YyZHcwUFLz
VNFq6uj/Yf4283SKuKDWL5YZNQoua6QWBmuoDYfY9TMTtZHoZI6P+eMW70EyFGplA8YqJJQ8VOSH
ak/tIKAQ6Dwn42tNr2WXHdywFLAz8UkwjeLeVuKLwQnkR0yKamJb3BPQJIAwvns8Re3dgYi6AIDQ
OmEppWGV2gusr9yFmE30KHPI+nAPIvo/EBpSDObc3BbZXNK27K4VqoQfTsJ3YbZVCfl5FJgMrg7X
Ld0RbC9VTXs/Z7INhBz3uhDwZGScvyLuUxGpzjAM8ICbcZ1urbcG2z0pKJ4wzghH+PkKVPA34xrG
OHMyVfUQC+szeSgNptYyW08lV0BJ3/YKwNy10FwXFgh6Qy2+rlGVh1ma6v6GPaX404l0mCrJriMV
4uZSS/7u6NeOGr2izkUJD0R1u+JeJRCsCaR7JMbhBvU8+8imHL5S37ykLg49H3zRt3gd/lGXR4qn
d+ugu/0XjX4CZzLdZKb0+L9zILD4CMU2chSNTO7J4ELKt4XYlpQItPetTHGAkjIeKhA3Knwrr4+V
tV+TOnXIzG9Xw2DU6SKBNcVp3NPdhH6A0WYNedMowJL7xq6EdcYyqz+dARkAg8snzk4B4dR9LEpN
H1u6mQ4VqIBY5+HdAWZoGOWr7PtXgk20vC/A7kPFnNX9vUOMwgbQTq0LNz+dpzmYTNluAKCi0LWN
3DZFyBgx1h3NextHS685qgjpiysTt41/KTHde6qYcxTKwOOfxOrOsN0/IEmEfLP6qiMy+nnDKNzj
mYdZYSujXQWgDguu0DI7w9g30AJwn10a6Tf2xzd3H7T026m4z/lHlfqnsZGmeZ73q5e1YmvAgP9M
UfAS8IB+ElSeL41GPSf0QtTLBY2cSk21yRtuIYvfEFN4PCXShgmvulZ7YTJSX0h8Af+6T4gbF5Um
TGbsAkXlFLdv5InyW1zo9+aU1Rke6e5ZmBBJ9w11AKOWBec4ll/KbMxYQwyAS1fTbbAiggebmWpr
prV5s1ZilzGdQeF4PB0QWrAJ3XooqtjCtxdnmKx4eQTTQ66yH2rweldHDWuDbaPcvBxPByxzaPHx
/T45WT/bUxWGv9cB75r7HQr44vyUiPl7XVupmFrD2ZUqrY32iTJ0mJUKHlTsK2cAnv8Y+CrcPkl5
kMENSY5nq5s2Gj7F+pnEEeVnvM3HSKezWwMEsS0J5aw3XCwF93ZbqCNUDIMsAwVEHr3nhP8NhK9m
mYahvrZL6zLB32pXpucqp/Ej+txNkJJAdYjpTOOObdnChNOumzHwKo5A204TTeLX1bphmjDnu3zM
EEjHL6YU09p2eyfAArdfx3h5MholxWtNhz0VPwXrOhdpMkkKyu1LbHWP1JMRQvZVjUVBXk6exw1e
G8zriKur8B3gfrdWLWC/xKzTxNt2cqMOJZ4c6/Enypy4LHi4Ggh3ozmM5cvQL8lu5QMBYzHuJk4o
Boj3orJH6cScn9205AZ9bKdCYh1Ruu8MsEMTABL3hPq7rMjr5x8j78FLaX7LQ/0gCrl50UrUUjpn
VUYzva0aL8PQm8mjbaF6KSLthiFEWZVQmXxyksEm0FG6wBucvxgxAUHi6dy6sKid6Ap9RgK3OB87
3dFPd3oY3d6QR8O50G9bzVm3ngcPZCxTpxVJN64wzl7XMF1K8Aj0MZ3JjlGHT9Ht7o5J+qpBYBwI
sN+i+pDjYeogrDiJQOkxawV4oyrhRHjgLh5atQXUOmn3xopjcVSNIHRdKxzYph+1v3nzW031SsxY
k1swGta9LDztnArJAB46gHEx2SN087lENsgpI9kkHW1J5EZwERGby2+JDFX+jPEZAL88FaUUo5JZ
Aj60Pp2nlzpkilzk7HGgoSAYf+hnWahiw76je8SVKzAuKBrlBtPHffPzzmmyXXAiNJBwOLSKtBku
qmr7OAtJ8wOCA9wKl2OvoXjrVsCofV6MIA59N4P19vz/VaDSNUXVDT2SdYuWxES2NFB7FpN1+iNN
07t3joqsBZq52+BpWqzZmASEx8y6OiXt8/HrN+82ihn6jhvc3ZNP7UjgU0puiXs5fpGz/PQFrBwO
YftNrLOoya02GFVaI4h+b/QerADwd1ZGbwBHr27Z+4c6iUEvt8d/vn2ZZNlKftvKZ2QFdK0jfLNy
0C2hGImfQ1JeuifXMyPYMDqKEvHnWIxcUGBMIHFpoFyB/GDJhOdz8K31BpWqWaCNgz1iTmIxo9uF
j7/7AW0bCU7LTYJQzRtc11o6kUfYZNhlumtLgadUotj5wP+Y/P1wP0qlozMKPMehcIVyw1z7VFc+
0KZ7fuTZ2Hkaw6oeJh0XEA45kyb43UPZq1Jth+W3v9HD6+SlkAEvqcuXMwQmSasICai+XPyV6ZhV
PeUrVviSulc3AbEz54H1xKjksMAK0Bo5taaJSFN7frIvegyH0jW6jVHLRnqeqz9ZXYLecidacF2u
31aPBIrJYwcxUMKCrp4BDwLyJytcM2PyRJ4I3B7WSgPF4HNh1es4k4haLQUeWfOElQvqzU/pQMOl
YlKe6OzAPGJsZnN09C70UT8lQlk/oZQWl7aEJ9uoAVycOOH7IB3bDzJ1GLkIILuHkx5dzFzylVGb
Keu9lOiK6Q7MCRDQwz/eDU1jTQf8CsULTVEyj+dG1LlonKp1BHmtDY0SuGaN8ledGUv1OfiWTSuo
L09BHxNK7X1ESn8g0qE5UKmR7nl9O066RAuIuVDb+xImkxi0MG0Sat67Po6tK8Ba2CRAEJLTvRFR
aYdCDsLELBAujoJzlNxSfkpnz/D/gPv8BHALZbKddcFWZDkjOkQ/1TwVLJOSzHZU83xEmIqP82YV
g2ry9SpSnC6jX9YWz03gn7ihy/3os2Rkn6rM03DzG3uiaL6lHKo1J42PN+2tOwBR6MX/BjovO3U3
sZ38GT7ll8VsQT6jq9S83jyeug1ASZ20Rb2braEkgFhnDi7N7JvyzX/U+zQPnYIl6QdQmO9dcAEG
bJHcfGvt6qOsHqwo08h80xfMa7GNXH1WQAnzN21iinEOsbTT7DergPJEslMwrO/3ERI/Eb3fXHLE
tt7tc2M+bGSVfDQZyaPaxGIh5Skeun4ph8tz89Ooxvq1PS6+C0Y6Iflv4EGG3ItKrxuh9igUknIR
WKIaxC4rYcSXUAT6vlzV3iGVEvs1Aa+kwHyc3RC2z7NhzfFINKbhO61g3p211/zR3vyFFhC6nc61
zix7ZCScgU6p4dtRCUe9SKAVnkSLVKq5SdxiDUxWs88kiH+CvbUhaGPWj6aGAPjlRz5GVtFlplGt
eGQSDVafBnu4TPVtYVJ8uMRruZjZcMEyYEoHlA+E7Nc6ql79UiWz7sqxslG8hR7jIZxObJtNgOSD
6+Vwr7OzxUfz/3huJBkF8UakK4Sh8/u+pRiwgejRsqgQCROHeuXD2j/2YdDSmKL4NWhQAAF6oAqY
bfgph63Zz+TD2n55H0xl1FefvFroANa27JGraVzvRs9Fp3llBjFw8ohczDOEflpvjeE0dX4N8Rih
j1z8+Zmrf34AxBv+9Soo61ytcE1p//yXixLRsp+ZaGEE0W8Atiio4HzLZmUJ9qtPAilFMzrYA/JV
3JNZRhK5BWY0HZBO6Lz1CcpjoFMplMFDGddKCnOVLoMVCUqmJn2Mvfcaz1zt5QzFX9xhqasfNkwF
63+YsFOOFZmWK9G9M2WgnXGMrNOEU0+d71W419hnme7Ok04IxGG+ndpmCaY15rWg4SZ0vtOxjkei
gpv/Jxn4SHlEDpm8jaeHezUXaZmS2mxBwCpPO9VlUveT1RCLl9PQCdGfIUs4Wjh1S/7esWmSx+9s
fSRf9tg27SMxETbtrV5vdAexaoV7ad9kXxW/QgUHOrcXlUPGfHXxwQOutgmRACkjhpLivJoGNCHO
GO51fOCzPpecJXwFwTigAFwSK5ePLWdCBJXVZ8u3iO9RhjjRR6089INejqdyKQfaGuY/vvfm+JkK
JjbZLrFoO0daQhaPKvhOW5tNFF/1kTpARq8lOCWHWhVkpZMGVcbl17UB6KBZfQafphZTrxVVChPN
QhIitngPa/1L0F+GXPLA4QLG6fpQVTdZ4e6Gr+B4oesUIzKt6F3Jcsfgd+sj7Hml89J9G40e2njL
3lhj7xnUMNeznRSMVqiCjcOKZzJrGh31jz/RLtuxWtPh2mKUdrMalNog+bR2t/+44KJoKq3+RrJR
/RP2TSzhWstGCspBpWi2H1Aolbnb18TvDg0PzLJd0g7gvyL88oYjoIF+WVQrOl9m53SQ27BT1miR
Ys9caN54UHTyCLPzztb7o3Ibpd6VUlg8RU9E6ZZRgw72bBgkfXlBEKO6Q4y+o5sbasDiOB8a/Hkx
gsqTr2IUyHzGYSExl1H7u+5mfwNW8446QkAdjaGgTe1qqRRtuhexDyjBa157Zklr6I72I/+qtA1M
TiF8Xax3y7N3zfnpxzPHyZHOaCG6KstWGsbueLXCZaKJRcTG/CgkRJRgU8C1oayMSRKB10iEmj9b
1bxYuXeOZMwRO4V3vkBlKDdBO+fM6uZ/qpUp/pLz/vD+UHS4CqER6Hmr492Wt7kqnDkiypQSZhg7
zfj1D75SajczZMLPCrsWCjimaFsC1c0BfXh6AiBMlF80MUfhvvQ/OJRpazlszFyeCacowxILIMIJ
4Iz0nrjCK36hVF+4q0Bo9Y/KKR8lcqKzv2iMM5vcMsafxsNjS/DfYLU4tRRwWsHWk7AdDp4YaTkG
0DOOKoqTEhyWGKf0YX2Pfstd6wGKooyNB5+oHBpD08CaNLlFkHWgXhO9YTkV/VcB0oPSYCWKulH3
fpWremATmgK4GDLYLfi5KzB9cYSBj1h42BKCDkzElkhnoAyIq30C2AkdASyhOJ7Wreu9rMyy8L5/
8xZ76R3M6TCH48wRywyXf3N2YmWQ6oHlyZkWt17DnMiVcBzO+ELxed9wJPMG6RgEuY4ChhVMR5hV
zAZgSkBoq2oPrZChyXxsuBTp2BNe9nEb82jzH1YYgXUv9tMBfDXrKjylhrrNhT+du3p/WbQoJqCu
H77NFOiLRl8DrXnruZGxgISWc+8Qmaz2Y1Btz+pqzrhchbyO67Hf2Gyvq34Vb5Rn7+Hx2tHT9dv3
pRaoPJIl1HRY2K1G2ROaOVuAhBlKcyJNv0IE0cgSWgrGnH3JYP87euXR/Xj26BvE5s+TxO9BDE6T
7BP6XWX3sOhdFRn2vlM5jzS+FwUZX/79DRcGNxHsorpM0jGj1kq+/u9NqiUIDozZhmLb96WqvFCu
C3jvlhxSF8hDMFSqa/xnhuU0AZuNriUBJ2XZKfgaCISIIqXJt6KNcjl2+Rf/Yzi0DjcnwDQ6X/x1
E/Q+u6qlKhhw8jW9YbQnPwavmdKWcvcHOyGTqHdtJojZ+i1HVQfIY//LtjZApDmpQTyGNN5yjbD4
iRQWaaDV4pm8MN8ZRyjpcbn4wd++w6OwstrF1X+skXWGAFJZ0PthNzbyPA3iaH0/h9hs/2d7LFuz
SXHBJIZA/qCEuL361nbqO8GS7gjCggomntOt6gWWac5qVrA1y/r10QHRvFsZPs2WaX6ue0iJREHM
JfsdAdPUF5mMkPh3J9eg8DKKaqGOZ7lt+kBtyQDMUJx4stQwlx/aoLZKIbzYK5nXm7bXictA6W5K
eZ6n2T6HftCT3o8ikK5my/eo0br+ksTefprfDgQkPIB/TPDF9axb9pmA9dVDwqAODYW5qGjj26yo
6nQUaryWpwnLoyQM8NzJM9DqY67otA1LZy9fUnpzcSp05hmj4HWBq2TtIjbtyOR3ax4JIrIiiMei
7KeXYoj1ftfdWhSbVlJtpjjaoUVBPi2lZ9GRBGCElElSy0zHrhhD2LvR7c8LaZb7lFNIWWEiEXCg
TMkKgv+oF0mO3lwcGJ2C3zSkWYgEQ+EEML1wTxwRFXmUUnR3uuGxhR0ag2q2ZtF38UPNED6jQ9hH
szpKHM5RLylH+3rAx4n3CsIsQX+YxVHisLb2VmZHElA18el2owFP3U2iUOPau8EFFORmmAeJf+QS
SKyVCiQ/cVkysxFAqW6rWnB1zbAAl7+LLcuXAOrmd7iIrQ041TcTO3Q2Ft7T+GISAgxfBn3/axjS
70sYfdnO42ez4j2ZuBBn6cxjNdzrOT5QIC46uTnygTusAU36DRmIPFTaxOAjqZ8B/r+XDLXZ9lKi
/CX2JE6RD4yE2Fq7Qm3+MBe2zzSbMCTSJPGjADqXY4APLD4i2Fm3y4VK5zOaApeMVAz63WriMPHx
iuQ/uq/S4kBPVB++5rDOY6ub3I9KSSKm3sXtn5w0yR9rcsWiuvMNvyMwHPuHmINHui7iJh0VlrbI
3vzazUiLEee1P0wGCBp7lfcCv3z4dovZzf5fyyDBQp9tzKIgmyhPqyKyj5A6JkiYYmYJYOHDBq9L
Jxw9hiFtOdKPVuNgicNCRyM3fZToISshtOnEiyemPKSCcIPfDZBw4KMgCB0sGstKrm9dFRdJQNCm
NRLZS5TYuLvygMoY+qwccJWH37//rQvxu64QZTCnOqbH3kiBnR+hxIqiKW0k+wxjQTJ9JDBtTgbx
ebEBY00kVW1k0Pg8yXg5T88YyjlGEsNaB6oxtIcrV/I7jSWBVT+GlU1AtsngTD2+dA4LCq+MreXZ
hjyNklp0mpDivaPOf2G4ElnUlK6VZxEnm/qxtlzuB8ldgajxx4o4S3a8hr/S2sYoBbFYYfn6Hkq8
Q9gwnRnldLC9kr6yEaOj8WiSc25FfFZ6B+w9dUNWWb9LnPg/YjDewk08O5Hda4l5tCm/XNt44A+k
G01x7zl+NzNRcw3XQ5l83jRQvkj47WTXz0ziTnCtdYCxoij32HDXOvYQgdoYtj7ORDVBlOiI9Yrz
ElagKb1FLjitqmdTLuUGy0Fdui97//sCof2yFGcy/PJNR9Bg88u73aPHBMIpwrps3fhEMDi9uW8g
H4Unms2CFletIlxdLYIjUjEhBK/BUaSL96dyshJe3D+EooDEFUaf5Um73c/5FfcuA4G0W2w06Iej
YmqE3TIq7b99itqegTn7kUrZ9XqFV1yGCG5nZ2MweEkhAjg8Vn3uBhJPWF8r7M3VojBRysC8VyPh
CtjFHb9X2omvnmQgpJzHk6QAhj60J/7+FWWJGf6NyfI8IPZU5p5+wLhXGDqBR79aNizghxPoSqFm
st/x690BpDYsRl3bCSQQqfie2ABWUM9MDg57RAstEDVJqwfaLvd0g274ibNb3nHcDoZf5Yr7ie4S
qqL90hmcO+slv0HinEGN04Ksp6iLCkGlyJPtATv9qDfS3G0IbfuPEE3yGELBlpMWOIZEoC/RxV1H
IKLJkhZEEw2b6gQRZH37cOwe5z/y9hXo++xVnfVfrGVIkdm9Sy51yFNAQQWdn6UiiCvMbgHopr5v
roWCpDDWGI51i15wog4huO8RwUQ9Mi86dgU9MVZnypHQotMk7XAey7cu+vh0IzjhtGSIL58jCMVp
FOaDsor0OhfkQjswOf8h2tXwTxNRQpALCihzqA0vzorasIYVfQXCiHJxYOVR2VAlGuoYysIurrhW
UcRXVSR8+cgRn2f5qM1yAqPEWG8gN2Sf1mTn2ntKDqN704IUWPkvNNy6evBWrdZwSM2SlJL6xfvc
kBz/QciLPMah31DwJzOeXNXC1w/y5kUC0bFp4nUFTAukHzEGo3XURE6JJXAecVrOtFexjSMCqPD/
eGWQIPkFcaHfPLFy5k+YdjWwiPeb3duMuyXXWhLky3pLdqWw+LgOZoGD4IRjZ5ZqEqz3uwFEKFWS
006IQEfZwXqjKdZV9LiPvmv6a2Zsa1weI5+6llvxIHuZ6kvzcG93D4cP0B3m+Ai5y9IIDivVI7Ck
D3FS7yBq8ha6jdfGjpl5RDP7GSt0IHEmr+r45aBEh1wugL5ZKZyZWhGaKohTeCA3yswwP9HhkqZm
6djoUzF+ozS08Nr+ivDQJKclWb+KOCtcJz15JHR3zFVutBBDTWpu/c1Z6YgKdeMyJMT4HsCe+FI7
2kah8t7eg6mUvW+kphXKc0VeWyxMKrW6lPd+fuMpbSjRcS09YpPXuLiaN5XSJ+71Xn7hB0NYwO7o
79fCpv+usYc7jVRpvutQIUTuvxBjRNmbPlSmcxvpnT2ZhZtrF2JPKH9RfW/kfHW7O/mHOD1X3P8x
uefxzCYvFRJ1FFrIyucMrCBKUANxy1RwKZyjm5f+BTnnq+oYO+6E3Hl30cG5fIPxFeybQtLJx1gM
0/Y4UEdWYwcrBqvDOcIrC6ezRO+m8bMr3uFi5yGgAVYUcefiOz5yrLGt6XN42t5L/PY+4t3wCoW2
KkrIDzmAo1lSyWiZkgpQJmHs2DFN7ujC5eou/2cUSBs+E5scUomlsCCQfy9nKaierlU+izjaCv+2
8uVvLRam9QU/zC40Vz98A/MFMvqd3QfySZFfxQx23ZO5AI6hjjRJ3GnO0PZmk9eCxUE6VAMHjuub
GJI+6glgQbUSGHUnfLJoHUA1BZTvJxX5+DUzrsC0QGRWND4WjDydySkmhYYmjM/80AJo2/7npIDs
Mc3SnQoCBjVzibMNvtj5S2cP1qzC/88SveFHBcc66e0EjTfd0LrpiDwdnsPJhgwWhSMhwpE4Hok1
7gIbmF531B52cxBMrlo8GT/dG30nPRF8Q2yJr+hiS73EUsGytOT0QQdRZpi21rM81n4Fevjx8AlS
5vTo67UZ7y1BB/mSVUiiKDMPbDjOcaGckZ0PLQBdW6lnFB+oSVzGBqf5KdUVdZxA0uDdZXLrRpeI
buYX/B1HOkxEFVB6iQEvs/1duwOn2J+x1jl++swv0L7P0PhFG5T86+CA7Uwqv7jvFl2AmaOoCBqT
zJA9XYtfC8yq8m/KXDWCwfn4Dn8jzkeSYQvN+HWX/bRGrTWG9vDP/q3qKhQIXFi9E9pGO9g+j5jK
MhnlvefgHu8REAP4c1j8CxyQpFagnUz/aDlRIctPet3uWjwahImKfh1Do9rZPzgZBX9e07YyTeTW
btzXbvJwoXPb3/ZcPUMhNrr1snpAk6GBNM7NpsO6m1zY/eupKhlUphb/iCd9SZ7qBET8h/VAFPUW
M+ZWzYlUrXxZ+zv+b+Y/PeUIC0DN5ijZSuqIRKphsQwipqAl5J01caL5hqQVuHIxzT1PXZzwKJJp
uW2NBt5iOJUmybkK2o1h05tpFMo3KTYburs0pJeuW96cABmcAPWwamceR9CHHgHnoNV+sQTYsQUD
iPQ/Q9r4LOzZh6eRlsvugdKOX7et+dcUUHQFCBTfQH1nYqenDdjhDpZ8727TZR4KwrSnn1j42aVq
BfGAHvDzNspYqHgWLqvn40WNv4wLaTtmVlIrK53N6o6WOgS9BPcOi9AQQKWQx7utPTEHyka5Ih8w
uXQySMVXxnWrA4RjpCNABv+fyifY/bpNx9yDsfdyaEfL279M1nvPIdN6ZOuPce8Ovuj8CnrVEeS/
nJGpi8d8lB+iP5RjrF/c0ja46gPkeNbszfek61FcPe1Mb/caUikw/mwf8zWT6HOy9qHCZavVPZVL
nnBm/d7xSDYpW5OCwqM+aAsvHP4Id1sDBKm3ozg0eF/PuPtI0McDOIn5sKRhewCjt3Ll0rtt5owf
UbVI2Uzr7y94auJZQ8EPgDZuWWN+qqhIogfyHeA3uqPnpN81w/MVbdyeqmiO2Rw7iRRId7p7FaGe
Gl/jYHUSEbh1QEXfz9zqNiKui3PTUmfc713syG4JyHf6M61cUuD94vUED8HEL0ke8CxtlRI5cA7L
VXGVze3mh6vj/73o9v2oOF+AAIweGQXX7/YKpqnfvu+43ckDDuUllJr/DfPeK7Rorf/Bis3EkCIX
hQ3PaEFLiEDerqEKk6EWx8L7QTsNT5OUg8sRw9gbf7+58Gfa5Anaxld3gYRxZs+icGkDQMY8JzVW
zIBkyoZ6SRAeEGBItOJ0C9QJLX5T3ymjOjsQGTZXq9GI3YzFiUysPpjK0op4ZcyIWNtB03p3mHUj
1D5npsEKMNSc1Z8K8rqqY8HDZItBHou2sj0ZHU3s0JHdGGH8uES4e0yQ4EzYjdFp3xbzew4UppHS
VACUcMBI5dmUkk1i2BdtTZXIHRgZV9+bu8rJv6caIZfPqwBBYeF5JTdATFExDg0Y2im4K7GIVQcQ
ZuyWHeJPQnGELOutlxtaaMPFNXIZ8Zeftqdpgz8oHMMKy2PVGZcOjBmJ3Y44ezcaVaQwVCSN2bYu
pcJV1/SRFpuHFgeuuU7LDQF+3u/rWopOCkvtqiAZXsTikOlnyugXBhicHj+gNQdhyQxsd4EfN2PA
aPCubTzd2M0W94KG6DYk9mmxDGk00VYjOXF6PGztMRPOYQXh562n+1bR1DIgPbKZrGFI666iK5Im
vG9ZVkP4zm3YDTOXeajEEzjirq3Xb1FFLcRxtWzV26xIu2Nb+sTlWeSpSQDz2Qr7npGsy63HLzbt
cddFvV+rDfe8zYDZK0WdHj0PUwfclrLl1VnHQtJ0BMl2mv6Lon5PJHRd+B0hkIe6qDOuIoh2NlTp
wp7hR6ySa9JVsELmkXIJyvv+2jsXSBgLWplXLhYfq7ChpAjvUdKqr70ueEScvzV6M2ZW5ZOQLx3P
OQ2Iprd9UHiSfyPARn0teOLjAjToA4lXh82C++H4cYAauZ/HRMCMAtftSpBDIRZ02ra4DzoGi80b
rb4tNA22nuZG+uLR/QnKq5+haRLTQ39yWLXXBKUU9mo61JwXEMjrcVPCrT3z7gOf1kl/QgrdbigP
2qCX8OD/6icCD4eAI3AJcIWDCUVPeaeag0+iXOnuTY7esuAV9Y+lLDutHvRkFJLPV21OruefRx+U
KR44+twEvMmGd/NRMXlViL3qtTo5Z6Do09lxdLZXA5+4IdTHUew1950De798rEI2pFRj1XzlQJAq
C0QRu0Hs930F9k7itjtlcH2c/IrznQOWpzZUImTcP2s/nwv3ccxX0kxMm7bMWm3dmik4Bskt+i+V
ZAl81YI2boqFdU2wl7C/jaJTUvliRc2DvGZKlFMXn86spagHOYaStqssDp4akJe8FsOohV4Zms4c
nIeHJlLKHsoJJJZQaa25tmonAEcs9nVaDIKDvLrl8nz5y5hccCJQkvow0n0YGG1NszF76BNOWIL1
tBTP8cRTTlpNYEBu+/KA1K0WI/EEkU5T/R9OOGVkWvsxZ2oa1uii10G/fpZPhkPzHXxDsUkj3s3F
Fp8yITGqbV+ncHgQbnPzNCx6Cbh0WLensLYde/QgG/ZaejTt9/FavDAjx0CQDs9dlXngd4c0v3ka
6bn4kDnQZngOyIN2kTZhqQbX1jOpRsq/K4CU58O1STWeo4DY740lY6+IvwLPZ3czDezhImWZVfEp
422yUbWJ1bHB5PQ+0kxaPDPI4HTbXeX2lZxowcp5dGehsFTVfDaS+pZ+WtZx+jrVBmt2y2Rf4JxW
nZLIgw7FBIQPmuOq1XYqCvng3jBi9px7RWgFJDIc7ESpmwDqfxwWX/y6c+lXI+pXwj93YXjrr2uR
tZi2zw7h1e5Sah/hEtFA5uVVX5YqLoJ3yYqXAUXhuE/Uaej2xDY/g762HYUsnB8pRgbMDXyqY8kI
oA+g5W/0IqouwaP0vCNBfaOn0sN0fm7jjQLu8FxGtbR7ltDoYP40ajz37+dfsjonRXmMbsveQKKQ
6F83uNAPVeprSoXzUI6ehYOGIAGWoc/CZLN9w7OH+n9CZe+5DgmglWlJZkjSaFKrXMJZtA6Zn7/m
j7byikk3e5AQpjbBbqS3GKPVqwQd/Jbo0WdZU42jpuxMLFOWgG9Jo+KwRfJW9XrIDDoac+gQbNE8
IyTV2yT7zOLSVDywSmUprfQpbH6bMNM6a+KoqLwxMu7fd9qB6y5HwYEjGDrWY9ZiGM9gGyDLdBVm
KTt/XEAJCFILU2N0nC+JfcwRL9XFQWseM646NAMZWFaX0CFEYzQNfCu5ZT53VjsBj+hmmVsUQbAs
/MG0/hnawiHZRDiegd3W+esTPUqsn6i6Q9MuAbr97FKMhYMiRyTmPWlPwgABWSpFTOXwDbYE9h2y
Vm5g+SZSnaaSb0UqTQpGSpTVKv9O5MyyOU7XO6bMnX6OFWdGCqGz7CypiXzwtQHlG58ZifJNmcVA
Uy8HEd8iaszflNSRnMnWX4KvrPW2ZWTgYIzMMuZ3v9wQNBJYcz7/BeittwhYNC6b9e1PZPKJuDGz
dkD5UaV1KaJtzsZLgb+dci4t+73MMHFm8icXA0jt0UuUhZoX7tsghZjr2KhNIrFHPYxgybUIUCin
AFXrc1UaKtLa0Vx/QYIhijpXcoHNU3sd3RaunvxH551+QzzpBUY/idJOhr5uLyRl7GhHy0Pr7Mzk
rBrt8kcMqJUjQHYLV6YRGUjPshOBqBMCkrsWhQLQfGQXv1GDujNFNsD4CTeLXcUAd2XjQ4lfQd57
Y3RieXIdUFFqfNe3ahpdQH9Dcty/otK4jC/ogTWB7qJ0TixW2sbIQYkD8MYX/rndgFMX9b2ordbP
BluOtgg+aBczmEmEvzFs54ywpxu1X/oNuh4OwBpvH620/BSrP3gRbw99Ct/jHB+yQwqhETDXl1+V
/NCu/Sh1z1q5B82ZgBHXsEetYEbTI87zFrWeEk0MF7ivWViS5WyQgAFMwcaUFVcLiX5LaxI9chSM
tYa3SNAm/5zyX1r06rwkPiqj7wezoeDIejBTdPchOZcAJIK0M29KyWbMEbNWFyYQq3sAtfRGylUw
7J5JkbO/RwfJ1bcr4cNKebMJ6W1s5ScGkcCPXeoQ6MMWb4iLZudKAFyLLf1BVsgtIWtK/d7Ic4Qq
JXXAVr+bQE9/fyTOiZzQ8M2kus5u+pdf6lASmCyl8lcoZqodJetYGTmBBVXqRuxosEIceqPhdkBD
0gXmBKbRJoE7RcT3Rr4GvKlaHfiJ1HFpsFH110v45+jhkOZSC0lqt1sA204w2kMYbScix/NIPxcw
zJxye3nhR3uZkeg8gUfwI+V1DGVAv/sLH5vgU1nI4CJCdYFFzNzDyq44RAbNRd4eKU30a02t814Q
en99Gw55ypWkSF/Vw0oA2WxYXD5JHNKaEDWc9w+fiCAHpJUdLh6vTnMeW//o7T2GJJBjxR4lyNF/
nX42BbWwFYHE86ef/c2KwcSgeKLdQQLTXz5jolixn6k59JUGXAesVvXBK3ZSBTJeRs4EDNR4M/SK
yWsTMINLpKBhtE8UNZeNAxP8Nu31tzJqxDKHATdGeXc2sEnaTd9hqv5ajcLhXJ0DC4OIDbJs+Pa9
aBArK8tvIzUliX4m/+HNLYHzWlSxd/OwMjp274vKvlqgg4WKjnPQrVtLqQdb3i62+WE7xmnebYX0
SB9V5I735Ur1gptEMdPtZjLic3C/uVCvUTo3zLaOoauE6GfD8L1t0Yd4Uh4KuJubsb3xOkS59p0j
I6wAGnSkgyi6+k+vxwzZD3w2KFvY3b+lIQxBI89oTgSLFN17yxpDt+qVv3E9Z1r7HNQjBsR4hoED
9idwO3eAq1C/kxBGSpWE08igRm5o5NQHCgL9nA3UO6EEC2wZs4d3oRYgOOFnTBYO2482y/BIauX0
GzeVCIvP1LRvuHajvO5O+JfAhwzRErDPEIRcP7LKQxLJ6mObOtv/M1uCDKEfN1Mxc5aGKvvSxwqD
+0T5kxWkF5OzBd8hxf8sl/ZsMvaUAEUDRI6v2A/Ocs7sTWDyk0pf3M1/CRHkINFb3fx2CotlS6+O
LFhnfRpcZ1uvDQ7WxlFYtYTHSQYuDWL+3AZnozq1HF9htXBB6Smx2Z80xXw4IK4Jh3TVx9wkbM8c
0ynrisvDE0zDSCZ36hu7il7Rc3hUCa3hF/F4TsiDizseJd3wnvqTXF2FXNhtY/OhQ7aiusU7Lfur
gE61SXCNSVvilA3/S38jbMPxtDyrXqrRHhHJ6pSr5guyMPFMzjGGYkE4R5IrGXI0TCiOzPo9qmzc
Uahs96kTBjJAkeAUdwXIUYBqSToDp4stcCVIMc8NdM1iacpYS9oM4dkZ4/BKQULpgrrRWwgZ0eHh
9HriGuEUGA9+gdoc+sryeFWyN/ptJn72xhEZjsrrIL0lqbyQJMV+XELTMyWL8cXCy9a/Jlyys6s7
0CSyJ104LhAIpgTqe66Szee66/dry+b25lRtErYO+DulKW4wXufogi1MQv/R38ODR3uOD2AbQy1Z
d/1J9SHD6UgRboRL/wwarOcDf4AYGNkSDynzGVD0As4sM/jS85ct3k4SpdDjqfLBoREpCgh/LnwE
D/BkaxmLngFEePUtBlr3Phrz86tgWNcP/CGSOOGMVTlqfwkZFl5ldtvWFue9abxVzIjiZT+B8Gmm
6YWo+rYpV0DxJ51V2pJr6RuQcm4zdLXszRBSu7kxYqHZsthuVfxOnQ6pO0HdgHiWVfVSF88/BAlc
d6P0XVm0dSadsXJZViuV4grz/PbofIx37ftLQlAELCXcGj5QXGM560rXjLJotrjtEcD2Sd+/XSz9
DIItVtKIYEonezXNNsd1zkKzB4RcTPdXSnuerh5YSYGX5s050f3nN6cbK1ah59l0RO4mczVcweMy
29iZs+MJF56GAQuHl9W1fxAz4AA7WYxxW5nTciszz6258bSpwoq7k1fpfYtnaUoIXqSJTXgJVwDa
pOp2ppr/sVUjRhwiHgv+5O88nVjg0igVcDusWzrk3q6so61YgiRbPVhCH2Em76FR9MCxDZND7OGI
CdGHbjdph/cyevXWK7/8ri5R4y3+Yv1sCqNGh0Mi0kPEnOWYKUYwZvH1pAPNzWc/VdF8dChP8Z8b
2gJSxylNY1eQLMaeTMusKDqGeY5pGu0jGkjzIUO3eYkRPFDbPRhJnZkdkPl6L/vOyBDDd4llTLQh
NoaowJvnMAWLSsxzSfS7s6AfZivRheytvKObE8MkxksSjiA5UrT9NMfu8MqSRMEbFeaujYXuHz/X
jJfTJYuu12rzIjBP+/+So2eZ/UCucdTdH8bw7tu77xQWpPLNSPCWiyfGVCC9KvM/6P2ZVfI+qBp5
ThhvQ+IBHMbsoxeiSQ5AKUf215NePxr0xhNPFGOMLgtK99oeJqCiWAV+k7hrFG1kRYoxbpfMxVz6
TsbOWR7Ne+QqnKaroCmYKB2BGfshiCWJfU0ql6NH4N/7OAw1rQhjAZeSUW02gbjalEPQrMr8QMDL
GMZ/WDKSyNPi1poWENR0ck4cZNPGBvOLqI46/91D61U1v/Kt9lzF4w5HBJU79dC5yEU6b2X1HTNw
bX1md5yIP90bD6fEIeeL9jYBV2fgLcIujmS2T3UL0BYoruE9ksevOsQE8LZFKnuF0zbhoC/Dk+CX
OKsTeAobkqZM9NrtBGtm139tDqpF5MX/6i2J0plNZKh1tdclD5OGMB6czOUejVYXPJ1qfO2E9voF
x3Wv3/ZJ54GROB9PerkowLWDzhrLYJPbHGaA+fl7KJaK1AL/o0edRuL8wYKPVshuaB9fuBlZorxO
g9fCYKJJO3dOYdd4RMJdcv+yHpHqjWBdgfy5+DZ8OBZSZmMdbgofn9IzXw1uXl+1Ho7+D8SfKJmN
zvn5m4eZ+AykegpccfOrhA3YgPF/5nGmAtgRZ6z9GuDJdDcyW3Jhy+Eq8BDczh8OUAF7MZ8BVmvH
xdNhtM/gyqa2pZ8e6R/8ZmZD7OxK+58Ds63pSxvOdHa7dIv8G24tTsPt5wKGqBkZr2i3qDT6pE0w
2YYtuz7yrzuGpbjBPHVFEKpNw4IYgzM2ARW1oSdIxFyDtYINtFP3C8C+zL4UoI7w9xZvqRVVnQei
PxM79VEFZUl35V0PAxXSDEkJl2aUKzZKAqHZ/+BwjzhPhWf9wnFNYtKZ5kzJrmms5Hkb0+lNf/Mo
etU341l1X2mpD64jK5ISbK4HQyXpYXemwyGWcPzIVjyLrHqCYD8NoCAp5fo69hquspsytcrCa6TZ
35bUZ6PI8y8gFn9vEUuPio0qCPj+Q0SXvL5ktn1/Lxo0tgaJoueZ8G5YCQyuWF83RIUWG60lhr+y
PyEbPvlsErO/LokZm7KJym5Gf1mEB4JEoUgYaID0fK1Hl4FRGfoMqFvT23Frv/9z9gtTw1DU/8zn
hZcSHJVeUQRsRZZhOQAQzl1C3WIxTY+DAXljwkgxQm/rV6U00WO7VfO7vcBitfuEhGmDKSJZ/qvL
fsqWGddZ3G2Aitru6Tw4qKtedZSijrV1g0kBHjLxZTUJmTA+of5mI/zn/rZC4lU/5Y2DTJ3gcDZH
wXVLjfgdG9HhX6yXXo8z4cPAfc2od6Htvep30u9WQlrym5/4OE/15LRtEtMB3wZ6fBQxIqQjCP10
Qr9XCHwx/azi6emdaHTkVOCxsfjUOMdgBA79W2QmHtKZdJELFQou/qLK7RJWvyyx68PE0Fy+cZAY
mJ9czMV7UPTgapzZ9fVgqWfkQsYuQa3+dhpOmmM/x7DIUfBZsRde7S1rDbGVzYnBywRzvLXW0mHx
OYf3xHenLOfP6jCxZ+Uw5kG+OZjDsTs3bXlF2L28SYHs3qbg8uVS8aRMrena6c3TBNxQGPkLnN4q
8s6haRofbA2aq9q2fyXBZeS3u+G38sRSJ+HOt+JgP021l4BQ4O94VMgWU9R75VXqnLVa3MlHHvrl
bv4WxBlL4mchtQ1+nwpvb0FzRWRo9BfBuj3qEuPrQ1zxu4FCLEcS2sFOaqd85DGgCFYsaDrHeiN5
EAPS675rblElJbilxleULJaYFREr+mkxYaeJ0fR9gVfR0GuBiLzAbt3hZdtlm141Aq1P5tXv6zsi
8RBGwRtAzbaKOd44qW2nBcV4LWs3uf2VdrHhQfO1a2mxpJ6Sd1MEcCT8lMt4WCTqm3BmqqzZyAFS
EyiixCb3f5ir8otYseuOwc0/QUb484TRlx5fdLAoO+pbiAhnm8FC3jEoVxwQEqP9CcAoRl9VbufG
VYds/o3BsKeUg7jX6vVDhWaDTHtt0lf7LJLSsP0wKofYhA81UsuuN0bPolBMz8UIT8pQOnkBOY9r
h5h5HA6/+eHsGkp1EP3Nx5DkJ/w8h4C/VQcICu4EXKEJsPlmlh1e5aWf3OH8y9tJJb37DR3yXPaw
VlX+1/DyZaWkrsuEybJrDS5g0IyjviRcSDhQPNJsH4tjyeyTKt/OCuPKGC3gUIfgXH0jPapJShqv
CFTsv/9WWijspaad/aLejiul9SD/pfvvGmuWTw4KKuj52FN3axMUQQmIbQNQV2wlI3G6bbVCS+sH
raA8+E4wQvj36uggxS6viw9EWRgG5floBy0BK+Nmn2gY9vS2ZZoXPX7uaNFMgqOb5+xfOKAahwsq
r90WBz+1jtMGkHd8PafgQo+Tc5CQya3L1jIrYfrehOFtYWzckltqN7z2GNmF5Df8HIiL4zAbKLkD
O40oh5U6oK85qV4jfGY4jeFY1caHMXVWE6mekCBX1fXC06Z3FcwfSAo8SLGatCXfWBizIV4pi0U5
aTtmuZFBdFwhNwbpS3tKfAxFNp3gJrEDZhHRb1t9avWYBQWK1Vlx7aw99OJa2xe63xEfEoHbVNTV
GNrpsYVfakAprEvauKuRaJYxZvAPO6gx1X4zVmKVc77DclrLGGmhkYAuzNonVUPKwZPCHihTZO13
Nm3qtean2KhRUILn3YFAIsI+gBY3DvZZlFryLK6YSFQYa/lybCcx6sb7gDcEzNJRyWWeUyR1+rA8
WSEykocDde+fTBis77NmbBPka0BWlIQg4MJCrB22e26QbRyL4QChf4EJoX5v8HFzVxPUhDwrvX6D
nvr1driqHXuqL45S7ZAGCX+hR3aom1jKpW/3WZKGcCtzDzcSCe/wKMGbILwNtk4DeHTIoRwA9ztp
FM2H9EK9DFi65MdLJI5Sr9xE9e6MZaHOPMF4DoVmwqGOUf15RmKNJodfz1SXaR+1+ZID0oAPcM1w
kxO+YtV1+YhzTnQ1IFgAB1aCRIopsDJAlYB98DBR1FWP+if0MNwHaqqc/fVECezaV4bEDfm/Dmd8
uY0LO3PGlIQWn1tQhkgMrG8lcgmFbgxRe7Z1Bsykm8StBkPHZVb+q7KdK5OQ2HflJKTh00S8EVKm
1mDL3CQUf84JJzasDj2bxOtrCaeKZWEzoUpO5+2C39xo1N/usaqZF7nG8UGi5yRtR5CQIojaYwF1
dwMJF+ht4I4b1m/cKG8y4iw5HzMBytv0i1yNmlKu7DVvwnRiIlEiRUJQKBtA8TSZzn4xdn/lfe6t
Qp48mCPQ5GQ7bZyiiUQ6fD96mDmskJmCLVFu6mRMdL1AAvJgb01lwr4UA5m44Gdm7KbiDV/nt47E
YfnoBYS4dtmsiyGcoiQ+DAATwKtV3c3HSipyLy+OPtmTtGanEtRDdY6A2CT1zWuEdSdr2xwxYc2m
1oL+RcdeMy5qxfoXeH4z28pa0enHpwAd1ULC7ycLemK8ikOilFz7l14EsXgI3WnHq7TihdWoAeaK
aPfJPN9RgLOXBmHKPZrry5c/XuTCqoJn95c3/izthul75aZzh1gh2kVnhtZsTCjIgBzzIvLuhIOz
XVFF9cqJ3DUEb/7AeYVctq98gQ72z0cPh82e8RjHrUEd4zSkbB/eDopeUVfbmBbIA3gPx7ec07YM
eVQKCheWjtgE9gBNld0yfe8SDnfzSYiHXWHEWVNcVqBjh7iCUcmRibk3Lbuz1yWRcvvVukkLFhz3
7IlwNbJky0kdO9UDxarZ1wOifCxS0yKDD5xMXMJPGMFohDyFxAVOlesD9m1b6IivnfsR1QR+ZHB5
YuBRiafsZyaBygQuxhgc4vx1K6fW9rPkAnNXIW5R/157rKDpqtwCrwKnenl+KIPuEqLCIxLQ0TGF
EIXoi6Ttd7WeWM0PqvoqsAsGtfRp/IQQgDctci9EjCZJe3rfsAbIz6Zoq+gWZKZklZBzn1xByRTe
CyQnu+q8AXOUbknaEewZVinScT11AjZxnPkCfUQrfptSRWWT/55eRp4MBsUybZEFpvHjwZTWJf0k
lFI3WGW0V5rbJu2QlZvEpUh3sf7XGPvHRw5biOW1OWCq/QgQKWcr5DRD9J0D47PQ3s5xxqzwLV4G
miO1y0Kp+GRT4/cYV9YJeZLj32QOP97yhT+owThxhsUfWzV+qCWM119Fa8Hb1DSqGllu85ff8+g8
9TgpGvy/sFXYTs8NSAsXVb3FCCyzzIabq5qNZfRMIhWX6YmgTJewd4ZMv/bob1qY2B0oO5sNLlh6
OMC/3xEFgAwtGDK7mCEBReZJbuqU4yCG0SMIfTsh7kqRnsZhIGL0J135TbqdTaTkAeZ6L3EjToDS
egnvEMMn3XgawLLbiwCKRVr4qNf7ughubvHZdhje3VADc6Eimk9hP07POJtG2B/0hoRtDDDhD9l0
7VfYHO4T/7pm3U2IGokyWCLNwOSn8uFOcqSaCLZZaErpyC4OZWpYbyrUsCeYV+TmH5AaPBh0K63E
NyUxj5Yt9S3SGGi3oGBoCIQG7aEsUMOj1hbO/0dH0AekqxJdYmTDBn5F21erlLvzuluY0hpfpatZ
qy02Xxua8tglEj8xTOkEeCGAUDQ2/M+bh6Mv6dBKr1Ika55+bXkorDmnNLUOV8XLngxNUkoi/Dnv
VirIB/xq96cn8nVdrWR/qeOWOYGGFYRxMiTciicZk6PpbbwuYZsSQXRXXtjR3OKmHs6cLQlwwtzV
urTmgf/dYx9Z+/yQ/DJuEbBC0qXij+IixsZFLUM1oX869uHrPJ6ws3PQ5chqrqp89Y5/DI4bbvO0
25J5SOXHqZDP13VRt7wEeAX79Vgne+1xlyt0XcK1PYNEaPYcLvqKdLkTrXH+4duyBFATWl7WSCXr
5eP7Iw2SCbAXKPGARpQCMWzyMa+jC8WWUGfqzC354Suhnbxg5q1879hZ+ickRUBR3n0rqwYsM203
/i1C8at+GQdwHF862FyESRnDH+U4BNuTyRlHIjdIGty+oJh5mImk3tx3BXExtV0Rf0ygKS3jSJpM
RnP/8VKhSSUHZ8n8/+B2nFfsTPtvVLpz1H9hRP7xF/wsKII9J9cZSQ007WiTqUNHQgqX+EjDpMp5
igIiFC/7g2giF7WcCgMbxsPwszej8GeyUmHe6wGYoCsY4d0T2bGSJ71EF+srVdrhTxaplksXgLP1
ruPKDWTlItxfD8GQ67JYdeJbsm3nBZmLjpCFHyqe11307kKCEI0eXRjVhetq1JZk+k74AxKOmDNv
sfTr2H4lNZXWTW1bujP3MBTbVmEMInO+qUDYICQm9lNPgN+sH/b4PmnVCFapYEZuHsgBNuoY9GL7
FVwKmY0i5Al2pX3R5UHRF92W0KteLbY1GYApY/TeDD7M+JpJzXxdfpvqmCHsnc9LalliKgHFcg5K
RdNASiqBEdIVhcgSw7GFzwXRWrVfE6y+Pzv2T+cyR1IC2kdnPnANtYAP0dvCo0crEilWkImkhPSC
5sDlCfbxB0+d/zdiyuiZ/S5jHjMDy2NnWkuL81MblORWxw/sZY6ami+vne8xiKsBYyycNqMqPP56
Hsu4x+FIRTWbJs4XOwrJanXOoRmxjmHb2lSo8nxQyPsCcK82sM5oLW+l6pCk/97n6DSoansI1qCg
f8v2oYbqXjtP9ybOOmIBrztVAlr9KfF5Yb9UARrMle/Bu0jrlha1/Zl/1z9cb4HCdtL3yLK6DpIv
eIxoabRc6E3Nku+5piavS13aDp9CZ/JKUsc0GtIoyHwrYQjkjrh969EvIuFHJdGkztKbMcX7hh22
4AULXnhBesi0hug3pkUnXEQslI83qoNUJWrtKc5GSbQoVlQtWo6Glsp6cRFcBGGSJZF6WTSfOSmx
iGmD7e0/h6y9itIZuQ9hSE8BLzeSfQ13yTNQ12ZVuXDrg6Vz5RwcUA+Lc+C1a3oa1iIAcsyODXwF
aN+7Qh6SQ0oE//R2x8q9hOK39btiGf7o/tn36Y9e064ljvIwzgjtw5T8krWyCc4aGlKwZCm88Shg
sEgm3Dqth1GTJqunGkvtooOy0y1l/sVv8IUi1hhoTr5Yg+sCuQN9mYLA/76BLwuQzuulYCTziTK0
gbL344c7E6q3DrBg/EiyX3eiX92VUhFc/Ce66VFldOmN3iC4K4zbckl3JLIMR+Bf4HTQ9Gxqizdm
o9UPwVLbFQ0wEKh9oUOKe/Tg/T+9i13o1FbNAA27QsEAhctpRWZVCLeI3ihc5iJEqsEBNl/zDG/h
84I7GQn8450nUmT1uBmk4mIpokwnLeF/iEE553YvEDr2Hulhli1JZjzmm0Zs64+1G0HyU1ElsqD8
oBcAZuh31KGqdiPwVrBDOQFrdTQHqrFrpAyVtkGLTnd3jQWopAYyhZdODgUuNOfDglmgFU0yvjcv
ElbrEMaUkyAyE8U2Nyb5LZ0NDyb+bEenZQI+U4039RYYXKPZ7NwM/FaZbETFXGzHAX01T9zgZ3Cj
PxR9K6rfogw6fSDOi1JyrHZQ58tMmawM8tgOb/yIAO31mhc3YnSrYeJ6iVhVNMdRpTSgw0wY+O9g
EQX7el9xTCyDp7iZuD9qsg3XnC54VksW7lsB7m/tzNB4pNi7pgOgpE2g9kMUVXHIgsOp0RCsl+l0
pEK0Tku37TUIYx/7JaXYytLn7CMI0toEFLlPTPT6xgGDrdSZRzBmADb7/XNEe3ugobjJm6qhmXoz
vhZn1JLshK1WiPw+H/75REbziFidqGcRbmOvFN9uUoE3O8qLhgkk6qbQDa/vVc/3m/puFzxUfiTV
OB/JLIJ8KsQSlTis++HlZnn7UL2uGf+CLoYPDqczlZCtRdAxKuXUW9JTJmE7HZ9uRnZHoaSTTIi6
QEF4aHuM3yDQrhXLLD0DMEnMXhoI93xcsuFGmqiqwMzqd0+KiHTCjlhLUGSuAZZFXw6rEvrYk1bO
0h1MiMuFQAyQPv4zsiZADFcnC1WwMRqXT9GLp8QXKVHX4G/CxbWG50TGGvaMDRphty2CCLywG1wY
LYZ4iQ9Nr2wSuqYUhxE/BSD24j2uINPFHMK/hBzPdDWOdsHWgp35z8CBlEDXZ+sTYBuh9fx97qsk
1lZe6UaRFVWrjVnOUI7xQy3nmTAhNidZryDF/nTnlarCzYRUBcdxvtTnHMD+ASgi7GbTfj7DvJn+
rW/fZisVIADly2GRJ+Njd3YJWFUwdBepyO/K+2y8y9F+vfrmQ6U8AJz/KY9A5Wcoz3jImbQzntm9
DvztR9GvdcOlUtkJDdzzoB3yt/6VCf/L3fFyVkJEouNNRggoGA2OBq4NQtiYC1NfAIOILm+q8/n9
LQ9XTbkjog2PH4VD1cfTrutUsZAG+CIHfTcguEFd3GbIjT+e+cEC8aPWhscwGDsKXLbUIYE0IHjR
JNG7HE/PKzlTuovZgVkQr4Tezoa0DZZ5ycy5GnfiNIQ+blBFm9aeCnV3eNgphPtVGQgWD7emjhDA
seLd6XWrQFj5OJFFUUWJo6lwLWSTlcQChoXisWI7CTGUvtvewZMbfeZMkhs0N1NaCkFTbyoJLvvS
oi038neKekgjBkQ2sCg/DBskikMeTvAuRHwsV7EgVlUdhjmR/qdVcon8Gi//MnJTlkKEaMffAYec
4v0UueOfJfZnMDnSt481diCYGjfF1SCWJ8t4njMUw9txhv4+Vx1xnLeS9Kn5S2GQriQFmkvS2A/4
1kalTO/XhEeo8ABMsvJLElrdYXlBsHkwhmfoDoSkcUvLj9ucETAgBShrahtEyFPPlaY8UwCc3AdA
DAmr6xgVchr9fqa6bbZXMe5ZTrjqzhGyNBJPfzz8lspkMTfeYaMxYfM85BfX3YbEA4Sl1FSWSHXw
/03VY0F9CA9QUxhAemKMv65L9qSlw57Db+qxNqgOXgxFs5E2joDDcMZVljkP8Zhk26SFYbaUQYsg
yXFKBQGvZf+1VO1FVdlnIW6Zr0QPKIYsToCNMst/0T+bzPTpo2YyFtgn8ufxHzS0GX+QlQTE/64F
+fBan3rHFNxbAEk4eAozdernRcUxjYIfuWmRV/xnYHA4+fXcU9yAGaw03IVo4ZJGCYD6G2ASfhov
o0QOiijSMMhyA65xt6bqDR9FPXEEiJgnAX+kfbOf+rESf9h8qgk2oY/kLWaMKzQ71snFxOlfyFit
behLZ2VtkgIkXpRlgQvSz2v9xE9tsyPK3c9QnFt8DQXe0V5dn8JdO9Gfd116KMaB5GuH/N96uZIJ
6dCTh8Kps6K9DEjamTz6F9YqOKInRGlD6TFdh3LOK0vx8LcXBk3pS3ZAevRpzXtf6aJEFWxfFKmY
BI1y5Xg9ygcNqD15zAAPI2Fmeia9RCIF/biClNh1Vd8AoTMYg0s7vec/yq+XBSZ382Efxi+S0tw3
q8KhrqGhkhhbpKPvpPn608ZUH1X4deksMCu4bdt24NfWLxx5w+IPMPFUtcVz9SZwWqB6Keas5KM2
pO8lIVTaNSCrxaESJ7qcibymLEXaooCcGwKfLewuJZv43EzDKfzT58jHmdh90+eXHboqcR3K4yKA
6HTVkmMS5ATWFdApNEOnvtSv5B0AfS4QvuA5yXBHVfXblFw40NzQp9bD0Yv5Ku8pU7i5j2rLCeTI
6U4lHZw14907IkRu+p7FBABX6R0/QGPwbfrVFZT0bCBUndftdPxE4ESNQFKVgrwLJsD7p11I38N0
W8XGIvNeBEetGjxopFG8jmxjg1T7zS+p9KJ85ebpF4TL4RoGCY3yQwW35ZQv508PiM9DIuB0rKeG
40RM8ktijFMDXdkSUEOpRHuZl/RQDZksEznMX6wNfXglNUbjnCVceYtttuB4dCQ1qAVwNNxrf/JO
9qdoCBESUVT0Nq3LWwme5cju61tk1Jztmo/FRuygtGPNrGwZBc21aiMib2TMnCgIqTG6wF7pdbdR
i7tbG3ZBzEkCydZeAoX6lAFUymwFaPe/JqXQHCWD2beAFc0hC3A/8+upqsprVhepjCHUq5FKs7r6
obKukgJxLQrr5eEpFfmUJkvbkMrN0PRIJTBVyIlCj8cPV+C0RCRKD9Nzh4zaaCojW1H4HatwO2sa
beTfYbHUkiC3ONULJ9DoNYgKsIHXPkjZABvLDiEmzZk/84E2zac0XZzu4pIaCgQgfy85qZ0vXzJ3
9oEhOboiyw7gLURTIHeaS2uwFlvlWaD6bm3fmJz7anuld/hsZrqU1zeK6j81qTYCZQO+egwyNbUn
5V2yXogypafkWLnPTlvMpdscokL6P4x+6+gnimE7pWyx6gLSa0MDxLVV2+324VOIuuboFZbk1Bjq
yoQryjJN3jG3qnieN4M4nJmUYHuqGy7YYIk+picIiZi3dCFW3pD9cpQq9dfpv5UwuvaabJwRmJHB
kcuw1ozm+UsTikn2aBx54n1ADL+7WWBpsWSSOU5WcweysATeb3yen4tUYC4dhKHYxNUEqUQY6YQ3
b3x5kysvP1+fkcxuKlIafeV0rgthpaHgXnJDtWuEzOwN98ywDQ5OGfdqJi8FSPNdtFd0DuphfVDh
BZ0wpnwDjGcmXIlj2MzRD1Yu+t61heoWgv5cbb8ZmqSgvFV5oG8EkZRYiaJM4GoSFMbE/ctPkRWw
t/Y8ULbjKpC1j7JygNhkGqk6b6GSfRznKUsCBFnqQjD6j3n1DrVA1gK0kTZcdYCEgWehZdsw7JKj
nIYgH4XNGh05UuMkuC5bg8cuFTSO95Y9qjLFLoNejKwsIO6C+Plfr9dAhBhvmnoZQRGtQMUV18Eu
j9sA0P4mGj4GAfHZZ2sgGFAVB5Q9kBlVlcKEMdXYRxBKIdxSj602mkFqZNYLB2tlxwaXdXaMU2+Y
A7svHGMzEMnYthhyFFoSQR4APCyUHHpwJ7VNhVJt9FwBcloGfjrJ/4m07jgMKvBLMhs83jrPHo+a
Ef2dREg93fn3KPkfLl60BgJ2YtvjrtZBXeBTYklq+xXxI7KasIKV/pMqgcAjD3/Htc96mIvRBVwK
BIB/TNX4zJbBiLIa9+uIr/Qz4+rd9wGqMxkNGJHF8UhvQc2Vip42ylbBVDsfxThdBJFmh+GBZSym
os3QJOwwM9MqIOJsAcVIROv9AkQZnHVSkfjc8Q8Hu8CDTRYQx7DBeE2YzXqiGyapdXnH9Q8olt8N
qJXi0pLw9FwuvyvIApFUSOs4O9OyXuXI9uWM3WGSAIHFxWX+9RbaeAJhVbkdAiEBNSYFLyLcbx7f
5uTY8ErlQk3EsVb2mvmFgORIuEFqDP+AAIFmaTShqvHaEtbUIl+Aqsnd4khqZWzYFPgwB5pqFmEg
qhmxVsa2Mp3pEaewmwgT/M/nFMWz7VCkwLfmLbA+/U1JjRbnSt0XOX874KiDQE0RV5twQSwiaA9l
dRCtSKer6RhfB/H/hVzkSu4caOaAqE9rxJYl9Rwq59UP4KOuRGy5Cq+6z3Gb1GfhLl2nHgrln37k
Y/Wbz8PIq8noJ64nk4Q3w3mDVgMTq4szGB8Cx35/uYrvkPx/TtopNyIN4irGqaOFXglrQlWjIYfi
gPjrhKdRp2LybSi30k+XBY6Mw7+gm/N7x8I4TVpRqV0Y5QTTZb3vgykjlcoWuuQzkMOjzVoPBob6
/Fgk9yTwPI57hYFPUFyLOTKzFIDHgMYng6hk7fbBb5LOjRDXpp/hHwRcp+fQMAgVcCw0HjDvuX0F
iss4RBqSSAlCtWPpHy17qK+u9ptqzPwD0zue5ORH1FSpUG2bjBlWIuj/0wG3milHa8/Pw095CauT
D3xuCANCmIwzoESUTKrk3ajQcrn5hFsfOQlcgpJr5WFq5T5VJihSz0obfi+D8/9jlVFSAreblrQb
b5hkRA/MxH2Ob8QyuMqGTwoZSJYZ1u+0IU8gIXo4C5DxvdgsUitT6XEb55fLTBYWjSrpNWKQ9IN1
/Lf5kTvAXBB37YtfFXxYjNrAjrfK52/QW95V+SiTx0JU0ENEcIci+BtITwpqEVjSlQe+ai5wIoXJ
HgDMD7Y+2EeigoKrsBkYOdzAomfFFrufIjTDZ19hEwPQrWr7wB8HiSjSHsykcRZOSDq1ltZ+kyYl
G50TxQ8bbot8YN4tnPHlDp0JWxiv0NiUVpPMwAmAtXqNAS5g6Z9kxYcUUUljm3I5NKHMPTqS4mU+
/iwU4cvzGEp7rwIsX7XCkWUJMw0TRwgeT2puzmbu01/z+nPI3rCn5cxGr9xd1ZroUfxhH/noOQoS
DApY1zoLj4VAA+4QBnXAAMjTBItVJ5ejunp1nTfC3Vjf1yNI25KI66ZkpenJpXjjCWqxQg1Yu+bW
+aT7i5Z0/Y5t6nottxQOPMg1b9Q9ztxZVxSclo41TxknvmTAEePE1R6T2etk3zSiHMR6uSZ/kyh7
d8VIKqIEjp4/hak+CJO69v6YePzat2eZ0PyedcnJ7YUggPGqRAlsJu3N9uHxvKXOlc7jMcWg+R22
CPPVxx9pOL8bYHTp7qRl5B3ugSeMhLlhtvEP7en3FlAYee9OiD/6X4jFMMeFlRPDvnXn7DARzEEj
ESKANjdl6icHZDRNzHGpybqiw+ETwkZ2wv+drp8Zy87MBA33IX7weuVNFmkhFz17mdrbl2JVI50p
FTcXK2kGdoQcBGzMUddAXDf4P5dN0S9JRl0Xtp00quZLVo80MNB9AHJ481xcubA4hq/gswVsSfMS
2F83nal/s039U9YurPXNWC9LxiskNuraRqeF8aO5YOw72eLFNfJpo45LuDCT3x5DqV5dLjUHnkG6
AfXvGbkIiuSL+gsD9zSltwHXv9POZpbEOSMzrXc6wur9txD+KcUpwdGlovjp17n6oXRPCaBWaf7H
zJxxzhvEXE/BLx1SmCuc0SPPyobnecrjxyUZd/ibsv0Ipt1DljkNH+l31NiMDhQ5f006xE2YAMvN
kgIo/oy28jj3K5Vmd/CfiUo1xdPgptjy+tgG3Bk2dwlIQlH8a9BHfjZb7BchRz92rtqh1BQJOp3n
Q3nn2UmYzfXKgZt6vw8x0yQJJTJFbNmVV3rvaFv2REHi7VanmVYuCXcyhPCjdKEcsLyX5LI1NUKt
vWYMjhBe8l4CJBg8VrE5CZD+J0mVHT+MJU62FIyCaDrYGnagRSRkMuWhaw9dGMAs/SQGiaFDAMP5
CCIay/RYQEjAx0+0RhaJUc3k2YZGo/qyyzIXr8plSApgOsD0HGuuQgCjQBj+Xx4H8B5oVYUSlVnw
328x3X6IXFvZ6jBt1sduD1UuHKJzgaiJ+9uZ4rcuiGs1rUcQSEqNPMAsW+CN7QiFArcCnIgrbJZ8
UQkYbb9suwXpAqyrCJ/mTZKd8cmjgm2qKN/yZFEG0liuKNXv6n0pkbFa6elSUDNZe2xw3HTGgOTo
QL2jKfdleC2MGSWHQ9ifflxOtyaglUzM0pENZuliQhMIwiP7RU7IUWJThNQCYsUOKk4HRZWTbi6h
0Ltbo/+MbmdTolyrxxPIWW773zURJKkUnXXl0Uh/5uI1kiKXyDHHWyil1xHBM7Yoe3KWm1PUB4dZ
/Pa35opgKfSNYUEIb0zDnBGZJqzIeKXAeQlA6X549oeONHEBuqcTEmf19as8RPBwmZSD64CYIEoY
H9KFk//k8Um/4uMo2ZWJ9nYU+yoM+8p5sKwALp4HZ7yG+8aeSIxKJMBcEgOHxcAr8+n7lOk2drUy
WZNaWfCDefPd1Uh0qno1BEHY/V/oZnZ8MvEvx9KQteieb8uTQXQvoP8z9x+J6S9fAd8ynKatA6J8
YH510Zmquc4mruwik+83f/VMttZwriPsv0XkaFfwY50iHh1InJQYe8pUww/324GAptwq5jsXJrUu
/xeMByuELq4hWe8fq9+fsnKTczzA0l/b+bUwCqoYBRJq3zvNWdSIN0efZv/2+pJAapK0xburz7iC
E5znqlZkQGecdIBCO8IK64nwtWVWMb4PasGEIBlpWoYcgOuEB+IefJ1+ib8t3Dn1AXlgBJ16M6Qu
pPcFsLYqCeR9gKU8ajmyWUSekNL5zE2C0hSXpB7xhssD7gkcmv/xU6zhfZwB+raHknMjQsosnpg/
Ea8fArBSpjas+g1biQwWjrZ4Qe5cHPLhHSyWH+tw5nNvookyUqxFFPFi/CRl33/yd648x8PYPXtX
Tu+x1AlIqZuhhTEVR6OqTezYi24EolDm6aapMFLjxQ2wK57h5V9DIEa3YbzUCAXNhfQgFPGB39Yr
7EAN2Y7ehCVHj4nmy6Dwe1S6i18zVsAYhP/PwAbLKUSeUhb0Ch7gXEKuIQQo3KWeHMZx1yDSKnUA
4S8XlZLJ6f5Wf+FmKYxhrAKJNYDOyyISKKOjeSRz6oD7YQGE/pPI64N243Qjey1FuL1KXaN43GTV
1t2jyWJxlhtzFKDSQxHmKrp3tsscOkCRcbI95JGBz9yRG5oSO2BOaVMV4yFSoi0ow2WVh6/7KIwM
qNwMtkKfxMK3Evq3pAxPNaOGdZzW+MLs5JF1E2Q2UF+8EeMgTy4wZxyXRLlGRR9FaJyd5seEi0Gz
hxPwJoE61ekuRulApDbb5YjL/dUJHbvTocj1GFLeJdVfPST7mgEO54nmwY4UQF/S4KRwCWaB6BQc
ajjCL/diO1uk3SDOESzFG4lUPu2eXJ+hKpIvCCh7bHooizwueTqJguAOYcIy0ylmC74ZVnAEpGm/
m58URn1eEpvasowcG33WuVjZ4gpHfFJ+rPpBHO9l6A4OayI72RfF6NzqDB7wFD8kq+Bn9HNRmG9C
Ki1mmzFI1gUaW5cVEH+Loem4EY//ibX1yNn58SJWaVVGrjYVPeW+Wc6hNHZSGXA2Bp9SaZh5Ep+c
BLX3HcCK13WX2f2u5lHgZyJF6MfbOKc6rRveOVheFyCfWfsDhjT/L2zUbjTZHiqu+kPBoAqB1Mja
ya+gRMfnTeXoqOwnHi6K/FvXg08DM9fFDQ1RfdXuX/EMSxf+81R8XfPI/fh9QjVZjr5iqJF1BXYo
jfdcpO0dW4KQRC1s4j5xLjx4tE+SijC8/ZaifyDQ43YOxv5KApCW94ik0I+OlzHGrTrYIsGsYmpM
FpUR94BYdgnSNuoSsmYjrjPHCmQcUSpsRoPXCNksrorFG7hZNvbBtHpxYUVJnJX1zb24NvVMtvVM
X3HOoDu/sWR6rTJeq+cNJlTTZ4zcGBuJZUD+aVQoxVlhw5O3lIbddO1hss/eqFp9ee6goM2j7Sue
gMIMYySEAkLbqOKnP6g/PCgCctocqZ0pMxVz9Wa/U22mWwk12bXTmV0athVcAB6pSPFBHHpPlWFt
W7KwuZy8ALzNUxGsk00nPTiXNuqY2icdanmEUOCA0rfDW+fDzdg4ERa6eQ9jZ8200D9AUwOU7ycJ
FEzQsvCrZ0TtkjiVxPLkxSqrrwC/3Dc59Yu+a4D+pXCx4h1VFjXYZ8V8vwjAQIIHhMHOyod1qCI+
h9OfllVPX1BCAUiGO4sWh2RQftTaSCU2Gx+fI9SQwcrZXRcSqKVKb4X6O3+XoCgegIKZfWzdz+sV
xuL2BwkWyn0+wkbKY66wvy3Ts1VIbJ2SJhhR0ro0PIQ+lA8lbOEUC4MBdxbJKx8zdQw4Mogmf1Z6
J28d5BVEUznnB1jYufSoy/sofaLZ0xBSbg84TpFH3hWxCdwcf231DKYEbjv/WWYlCKGE6RJ6Cbfl
dlqEac9hI6zcHIc/eeWL4WroRhjEIpS00cZtyREuN8Q7QO4bWLno0BzR1A2y0QVXbi19IcHn6SCf
IlYLicjL16V2oqGzWRy6NhS4o3M1JMannuJVwtHxuaZ5ocD/jWPmEAChYQpEbXmmSo1jP8tfeb91
hGexGLEr6B1MiLarLinHV7U27TbGXpnGlcCzViRBioaHsj7r5RZ/NozJQuwTdn6pQsjhwyMJ4TcF
/0u9MiAvIqUeeYMKiz7IuePcszacg3l2zZzFvk2+vYSd/1V7BQ401WmK9UFlGWVnoC7lcbQxapZ9
hwtPRUosI+yHW3ThE/5p6usCthf7E83I7sfxR2POgtFdz7/9aLVr2jQpAHO1OLxwviK1eR39VgvL
nyN/Wz9YqGlDcvIy3Eq/XF29ivjGdOEHXYvZkKW2e3sxOfp/BxFCriBkhtNfU5UiLDqV1e58t9lV
tmKjoS8Xkpt4ZWRxwDI2XTZLICd7qR0y4IOGtsmfZeY3mpmtc3Pfg/dNi5uYbL8uOqLxLCY+uzjM
SshU+00dsCCcgqz6JkZO/S+uhsUA/ztK4KVa0GWiyVD9+qpt3snHGFLtlpA0bYl2kpaL/urNnwjo
fhgK2Woi058FUN2wVcTytSKywzYqjcsEQ0iCPsqj4oQqjiYxc0t7XFZ9TswvgUB/rma7WvCCnS6P
++bGtidGvfXXN0GxWXYmPW6oXG7Z8pbozWLSnC4iRGssze6q+IpNWG5rnpDO90yq/eMi52SnycRv
6OJd2D0flP3ymp1cLCe1zhiRe/zEb6DIDYVPf3n3HWPk5NqibM9xuz0MaYw7JvJ0n0wUTkrURxFQ
sdtAJDZHgXXbWUraxraxln3gI3AzvtDibQijDBhwh2psxNiSzUwufupM9pBonlGj7ldAMQTz1/3r
AxwsuApln6N1Le97XWjaTN4HyPo1Kvwa/F2yf8mO7yqqxJfAKstFLaDt9x0T/iJzUQckrUaLQ3qA
xD92IIVLNrk3wonNqV15ViIdv0haqSg8AZ92RRtM+7IsJOG1SJvHBj19Z/vqxdZUVmAZPm0Vth43
q+AT3WA4k4R5Wz6L002TYtbq2PAuPIpPYWN2KpaQxcjb2cgOLc2sB/+wMrIKYJmuAMaL87WwtDQw
Yevh7QGMSQA2A+sgSL1LULQDOeIi280nen5XFDjMQFtVG1969BT4LxNV6eUYUo7kSrSpicQ37pWj
tA/C8+kw50v0Qy2zTk/YHOFgYjjylZLOrCWFlWqvh/o0vAUmKNhYIRynyhEzBrQHRBajsxCdfstS
n2ZWOdk29Wkv/F/f8zHP+yFt1ZpXUH5X4bnnlwYTEEsropjta9dIIXFuXQuTSL5pCIDG9SLNUbBj
4r0y7rtdsPvY+b1cJoEx0qUE4V9CxSvZwWbF8jTH16jkBPjAGy8AolN5FcQ/wWxXRbf5qOZnUmFt
ITa4ibXADDbrjyDaXrDfrqd71ZntudoXGbEJ+2jdJYJr6n9X+c3pLWsl2duXd+hkt6y2lj6h7K6H
loE2bRdxbyKnjZh2CqXdhAgTrI1UvdAxMGJCobrEROJF7qgYLTsV85cvPQ8Yh+SjEeVaDQ7Wgikf
1WzWs7RsAzVbqMXY2hh3P5OjUzVeqv5wzndBbUifUjVhXo4J+GS3XYEJBM7NYLHE9CaJZcreb8KT
dyZF0Zlyz7TTEzJ/C6YmFgkPnJEz2J8Dmof5qo12nQZdVfhiwWIEL6YwizZ7dCwU9cDohVDQpQCd
olQb7kbXVZn4aVLJgD77m1OhfX8dqNTE55kjh49LEicThXjKdj+Xu6unTYR5XrfkyG4pPXHCFZXm
7XuRQADjVqqUWKHfrOPL1lF9svaYVM6qLdX9fRerRfugaD9q2l/Tb7kVsLSjfk3tdSVxHOm8JOME
H5KSApJxB5WJ4cwL752GhLcPaF3D4z5at7uMDOJxC3SggW/V/P1Usxi/lGC8Ve0dj08dUAqdYR3J
wJ4eKio872vF4uR+U9zeCmvkqkPjmyoRkt1Y+cEAT4WQILF4HKV7cZMe4j7AjXxF1JvCxSs//Pgl
BR9gCdsN58yOdD9898UvRDBE1a1riZBG1PCcXrqls5NRWyyKrqAoHKHNhlJn17MCjDcAFi/BrGTO
Q2s8yniLEPmYZ6smUXJCldpbW+PhLsfsy3hkwGKQ1FKYDjJdBSBM0D3Kf1otb19eEPUfaaNg1Ztw
HGvbl6Utf7A4s7buewvQ4llCs0DWdaMzpZHi8c7wxXvBgt/nwg6c8lwi6rKkMqerMobCCuNj1vEg
IcsJI912do/O8dtwk65doOgfKayRjgcyOZeHKxMU6hRCbMRC0oPZKqujg0hQboM2k62sHBZtKtx5
AEg9uwigzxZuJp+1cs15tmcLRt2Cmmw/mdhTLY2zTcWvbqJnvxPgMTjvLFpiGngwrhvZDJazSp/S
X03AK2SpND36y5ISZ6EV0oJ1Da73fSGBAj8Tm8gaxEfamSfhRiEEOmj7vOtxJHYiy7tVsirEBI7V
dA4K6hxzHKyVdkql1JViiBfLDXyY5Jj6lT0u6AXaia4BWPjuR3zVg9jPbjcfabOWBPMpGDz4bwc0
3CpHg7IVS4U9+qA7fS/zMy+zkd1+kQwz09fTZtVkxE7LNA06H2LO5xTVj62maGI1LeWwn+oZf9GT
qfjnU2PM4jxBC78vJ3HuQDT8nZrErR+QjwFd9BLH8EoKU4+uSWnwhKpQ1ZnUHLxLsJneecFsuKpy
qdd3gbBFQo8AgEWsGhct4KIcv8qLPvF8nEdCrmRnrW//ufqy2V7nnXZUShEW+zS4Rmvug+Crpa4+
xtbFgCOw3F7Bk8bDSxLFdNrm3VidJe2U1LWZK/ttYVF/Jq5/xaOQ5VJGq1ftepnd4WxeViqnxc7M
kUCIoBTd4tGzMMLw/XCWIpt5ILw4FGVGrflJ1Hswgms9c32fFLdQ/5d7QSryy8TVnry622BHnVNG
6yTJAiBSuK2VMA6mluNTHsAbvIIN2SsH7KUfD/GEq0FiOc81gLHI7ozXaRFjnVzRPnjsQdXDCRKL
WiR++Kgn/oix2+Kev1HD90qxZ3SxnqP/u1QeZxpKSr/TlOSFXQti110wArdWA95/BQ2hrSMC/irF
MKO6/pwQR1b9IaN8juN+lpDh6+kOvekyHzyvU12T6L8LAgQwTZrIO8kfrN+MCSdgrBkdTDbjDS+F
FTqQz48D/sSCWjCPs4yqNEWmrTLIr7q7hfQCAA/nLklATb3B3uY90HYrOCdFRbacYao0fBquV6oV
js2i7pf40+0JZs+UygCSqdE881dQD7ZUETAurEHQJH05KXmZoUlDv1YW45FKatFOtWGHMxoSU2eI
+fuLOxK/aqMBs/0mCyEHneZFDfjQ13HVAOQVD8660zZQZLjjVKbShS/Lpc/Lt+cSNxtvhqNpqn3N
FVSqBU7SG+WVLT7n1pCr4k9iPaeQlMs6fpXpHYTUnAmiT7Iyt1B1IoG7MME0nnmFZxh2/yUNS8wW
+eLBP6p9y2J7znHOsCYpJJgVGREoVRmkIjli5nQKa1mE0QSc7TvI5UJnXujzAyt/gLy1VNgJ4kyH
BjHXGWG+iKArm5/qtLzWZOmM149lWG6snepaTPUm0RW6mEJ84ZOEwicuyiXKGkmnOYqzEoqvAq1T
aB9a9SUUvqjlX+lNFfSvFg5vetuyiFI33g/jyyLKBAFhMYimsxovCJn15eFY2YVelRunZUxP/SBi
7ZtdlhvSjUQ888xs6Q+dP6pX8juZRWv39mQLuwm+TGq6YmrBVHhZU98AMxSOVr+qxAiXnpy5ufVt
bE1zWZ/EOppV0ok4z69qcjzIpt5qgcWhn8hPUB0GhtERhRuFXYn6eKX8i0BBUyhorceTxoOT5cFA
t3zDz4mF4XaHphWg40CXQci73JgVrp3Kp0NN/hKkZ2FSHqYruHhQjbIa5iX9RO3B/v0hewzG4U+B
DaWAMsde+ViIZDfTjQIBN3biM2RAs6b2A/WRd82KoRBayRDg/oSwLp35bzqhz6SeZCiLDci4u87L
5uaoqxfG5PHPLrXy7crJS3NdRlLYAzzaIR219LQRJZ8y42BauHr3M/9IH222TFgkfsTkVfW1doXF
brt4AQ3gZoLe4/aZ9cIxrrq/pQY1II75zy27eI7+Hv17abU/UmKl7CKhpqh6IbCXG1DQd7a0MaEM
WDtc7g/N6j58lp/v6nILXSJn08XUKPQVr8gfRu+pyXOM75oSe+zCs1QXPuhobDP2MvtwPoldeQCK
86+dMhApCwaQrRhbc4D7vhWlMp7k1AaE5olbaQEIIbmW5wTCUIp8EUU+2Ng1ZL9U5wa52XRfGnUZ
bkNrKt7gDBUdJGcflr3PV1QP6PeXis6pkm4nkuEu5lZfBnbkFHF+TnYjJuZ/dDdZxN5S0YXcEgEM
qfcOC4m+I1PhMcXoUCbrsluyO7/e2I3sdqNEArs5fVTwvzeuPMRfiMlCfakN/hjZcB2onFeXoZEL
szCX5cpKqJ2WVAoLZYDd1oyBUtN2fqJnxfNFHX37DJWVv1RjFHCLuK021xfdRpShOL+76jXSAG7D
jyCjHYFuJxu4mxD8HRm+Fq9ETaWd7BE0hKTEuODlCsxBZL4/67y/dQnjN4ia+8cpZt98aqd44I4q
fIFoTSHG1VRsw3ay7YZWbUqH4v/4COXkpVcnExoz8IvzLIpHQTqsch1Bk6EgWz2PgWJt2qpYCIyK
I+ra/912kPOMvKmPwTI14ABZMDvVeBU/buLX1PqGb+zp5mPeDPLETRitowmKq4CdYyhCkEq8nDiB
+U/Jf9gSI+7kuJxA6ADFX+HOEn1FqSO+bel2XC6aAVnvxkkdr4SQMGkKIZkEGEUhdJYNtVuIJ90o
yPOa3hOaFjAMFgiW1dtCBUkFFcPXwJ8kubXJ1a17lv+8dcy33mlS0hqIVs5/R3tu3cHB4cQimJi5
KTVG+erCOFtd0rG5wm5g9V6Jm9gdAqGA8iZrRpt+pF5jC+dxgoqaG1uYmFloZA4GYrJsH00Xbifo
ren36hfP84sIYSAKux2PacV7LEYnCpCxctBlGpo+TX3eIwEyjrq2Vhp0FjCTtfRtNKjrRoRgU9/V
LVUlaQ7GMZ+rs3u5pvPLYl1WPrf6xWbyzK0LWvxJCIK8GbkkL9pqwDy4CHzxmuIP9nw9M8wlc847
JwPo50MuaPY4c2WjljlI0F2YiIdj8dUKJFEdPNphoPE8oSyT53Y6mLoTY4fDLDVDak/shVeAa1Qn
T/7CqO1zsZt6sKJFnWUfnONdQpJMKKwiWT5DknFXHsO8ej/3pfTJrB2U7tqnkXlaEd6i06upDTNl
qcwLKyxaSpt/cFJ09JEGzkjoD2CNrWzOWAF7pJ2ilyRWZ+5UdnSy67Z2P9RW4gdHOsFz3oEpP6L8
XVb/mXufrH9hDyg4BgKI24syrD8S4M4nJkdpr2zT9JTSU5NZQhKqhWWmsc+krG5TiPdTCjqSLeBP
pEH7kmkJXVv5q3Db09jOHR6eG+yFLIHCKRovre8afYTzW4o1HNuAt5mv02SHukeHzbizT+OEeiFn
DuvwQ6xajoqTUYguEj1qRPJ8pOZesZ/8gfHAw/NokEqcfHPPwzLo2tT6vaE+9Xf++hxhpWezBJTC
amAZjPPuJJnoExjCX2lkrCZYFSMcYea2zXN8HkdF80O1hkqKStAv3weR8qxiBFvWSeqr1T5krHrq
e0VtzO/d0CfCHba4usNyljLclMKIMiGSfw2RRnjpNsuqo0+kwdQd+TfXbhr5wvqLYsU4X0ytpop7
5prJ1X0ejc9mU8trNp3xIXbs7JpExXiir1+hhYSGqKePDK7+RPb1r4VM4/FFAL4kgaS8AQJPmJjL
qynE7OuM+JsxKgktQD+CQQQLTFu5ZmTTEmxmVh8d0d69gsUHzZ2AZ32ghg+gzuH7QzMDzRjIfh7u
cVnH6kE1QZKJ4TVBBcEl9p66/4Qfp6GME1a8TLRY/FIeuLaCxV/v1CLBUcFaCpwpiWPPzD3lVxyB
b6EjE8fgOZVqRU2xKhYZE5Fo0edCKj5LKET/Wl0gSqBDBTJDOInFNIm+TFJv/6mfrxxr50sCEGTX
uIf/kJfOh1d7QvQSLUltrXZZuImW/O3h5xgu1wNzMDhkAHvhbiYzS3ApOZB5HJJavusgzRvX0+EK
AeBy1UIeqF6+t2ZYWXgEU9KAyWQbVvpxNb4Ig7OO/pDua/LY6xarWD8elsQm/VtzLhpXhUwKq0Ib
WktzOmElUHbhwPi0TyIGgjNHK1Wkiy7FaG0tCPgVUqw5tgXqdFN2FsHGO8GOk++je9Ucfgs2GPjc
DOjD4FY8Xos88LSke8fYeIW9oBVU5WswtzNEec9/Icg+BFSCrU4/WQMFdoJAtOgD3bvPKrj42caz
Z93DMLi5dRj1rokovuE83ovoSEjfZPi2tpEjhQGxk0uhWwuLX1boKckyHiH+xg7+Bvsr9peQxrDQ
iyMrebhHjq3IA5ZhztQHpM3MLkQUD3JW8OSUP9+MEdVQOy2a1zejH1UN8qrAHDGbLshbzvT6zyhH
yGP0puoq/HIX2mfcmnDTxTaZlvbwAcjxNx8SFUQxFTB4/GoBiuPDEJKZNIK+uODs6hfUSJR0JQIM
XTJW4q/bsmslgzGugCCcm8B35ZPEgXBiUzSiqNhqmhDRftUvKwPrNVuq+wlcFAeszC/9mRxljUcO
3JE8cl8MCARyi1IZWxOuO+sA25mpvEqZWceetH6TNuFXDxPn06vKQTGFS0wvDvGebur3BZcXajCT
//aMS4++fb0UCt4WbZQPwqSrrBewB7EsKbvObkq1KRJBpn3fVcbtMum2tpHbN3IpkXx/fbqT7lhu
s7In1qK6PZxmu4cqWcIpvlRv35v/oY9eT13eZWbibaYnQtD+wRBP+KjQDdyM+19z/PTzhP1UCEDU
z3E4/Q+jycfb9Sc6vUqmVWt3WbdNXOjTkQHProNdbVEKnYJSy2wSxijQ3R9QKVOy59gxzh58UE8v
8TKbpnM7w8Sz6wvR7l3RwgAz5b95sgI1dSfBcR5EAml+PTibmMJShEX686+ElL6ervRI0xL2tTPV
xTeoG8W6sY/s/5Mnl3ypp9Iv6uTV2pzZi/Na007tckBglwpn6Hv/mXhQd7e2JKY/wyv9x7BiuSd1
JoKpPsNb41LWVtOnqj9E20LPGcPYKNIARk59JJyMOiLrLAMZlYu/OobV6nbB+b88owlSuJYCcKD5
4tckvcEFYO5a0Lho/cYL2zVNfNDeWqLZOGUOEoV5JPokh0GFuepn8OIsqtXbs0d7cnlX9P3IJelj
hy9XRWE7B3egPXOkAVsZKk4UMlfSdxV+m6nG/85DzevNHHN7HgBOYj5r9Ykf/fQH65b5SeCuFWWJ
g/I805Z9sV9mOrtBK6Iz8LeEb9utZ2BssDfof2v1VmHA8/LsUGz2o+BARn/z3ioIAdAp+7X8QieV
JG3fmf7Ze5oI+EyhUIptmnqpZHVUk5IVzIolVrwKGhawml2bDf5Xdjd5KOIvkoTaWGUlMUOgacs2
tz600EYb+i7sy7TfzauOeTovBGcnl45YSXK/pw1jduUT3gVfnBb2FMX57hkOodquk4O8d/fC+9xu
JwH4ncWOQLUbknCr+RD6OQgTRjeASEDrF12eP1b/huBO0WQRD1MI53xkYiu0qf6fKMlkpcnr3pZh
rL9N7I4UiQ+jBr+JbLEiBvfPH0tsFPyzHKaSkIUyWwYgK8TrWsRPTtVQJpGtTNOlnu3MBwBrBDrd
tIjKVfJEAjM/CL0r5I2gbS/xUBboQ2qCy7E6FS4gDXX89eQxQfIECZ7Vd3tCSf5HZvygQg0doEGf
Dts6NEHrcvRfgF3XtpeW3z1F3y1OjfnHMsv8GP2FtqR4ACwIWw6jHnHASBgnGmZ27o00WAILnClZ
GUolM3LubFRJkKgQApVxv3P8fMrWG0XdbrWtjyRmGu8j7lRtn/hzcu1eXbPwqH0EhtRw99i0DDPN
j2gRsXKN2n08+0EbcxNofc8n1hK5UAOf0MXyOBnMSDGFANoY8x3lueeADU3+epVWlkH6S7eUCMrC
w7Cw38OyfoYml9SFOC9pfPI/PUzOO9gI0ST6TZZEtIW8WGgm8WHOhREvOWOmbvDziyCFlXPOYohG
CS7ebf0g39xSqCE8Cuahmasu/AV2ZeJyH7V9tQyZoh0ZiZrXZoDAo9jHVd0eAQq79axv/tQKyP9k
WuuaF1YvgKCJafCqFBQ7SPGgEIL9hBuqw+n5Qt1v45pQqx/sW7/Tuh2jxxVqg7klfprbdbOD2ZEt
eusLbvEt/SDjKgYSHhQK2wgAXLDm+0G04fPviLlBOlBSVavEqzm3vzBERLqvVNuiGTACDEsvNhla
x7xmyP7sfPOIV0VF8DouMU8iuKHlrikgO/8V2MGjTrFDmzeIzdKpJkl74hCnBnmiN6tAEJBzZdLe
olKNnmAIdql1daDdjBYHI6LEwCvJeZ//rVMnEc0m2s2BsSNFSeut1IuI8t1kCSolizfM8fm4AT0+
zyB8iEm8Jh8T/s7ULtY95cwPUoiYLlWl5x1jEUDMX2ENDTskvEkYllw/qa3XenpVkl1O4AzOoVNr
bmXvfluPXexnKDZVTQMFDFqyCGFCUmJnMyfNfCChcXDjrjXUugXnHlrjaOnFWjzu/AqPTVmazg5W
WLUzIRHwnJz16XtXjsqiKZBQ50L8es3sCgoUmxGK/lquYzf7GQOZMK2fCro+yemfnGfdL08NAp26
PVTfbGy0+M7hP3CpW5DSiP0GbUTtGiB51svExfVypyF9VJ9sV2xrTh1LuyWY4xKY53p8xenjoPYD
GI0choarW7u1kFFFZhhZNmng44MVyvuVuDbRq9Iqch0E4GmDWQd3v2H7h8wKj7Ee7a2zq/PZbnCr
IjO9jefJVxXT8VdVoXGLlMkL86ILqefbuKMUd1Y5X9+E6qOnJqYRqDxexxIZmPUieRzKxcmG4HY7
lZ6EGP8CbG/E1JGHW5tpjFatyaaUvtYzxIyJ3t/wjr5Wpj4+Xbx57Ko+jT2x8esWsog2wCzjEc5K
H4tmEcKeRu0cWEbDkfKMKQMDV+6EaimT3mSB/D+TNa1Davlas5sab3wvwqviS8RZNULfS0tdYRhI
mZsLD3ePRTlgL9+2dHuQTlnxYaX8zkqZv3ceaJ11wUMdyaDeBi4l7s5K9UDMMAhnj02Sn4d/5Dvo
T3bsqKxP+ljoD3dBaFnymAfTKa3/VzJFDxz1KfqYLgLimYEIjNCzFlLihI8U40p0nzpocxEXpuB7
MshP2RWUuz3IKeWpxyvBlLxe8BH6o5s4hA1J2xJ8PQ8AaqBwV8J53fxR546dG+2dy7f77hkSq68n
+00Bz8UCPnQTJzAW3dnz+eWXBmyjfJ60VAZox1Y4o1E/mD+fsrnxsYRH0roL6OHeJBz8RPzTjdmx
K/wrabjGKJILpMeHZsFfevVuG7uqeDrHCmDRErTRMehELvOopd73xFgjwm+zEDgxeK8/2WGd2GZe
fSRHFr39Sd9h3oAd3LiWtlRUsanZ54PV2RSfWcdh8cpvo5EXPFsvwrJ88ErRljU5EcMK/LL7UAQL
Qy1RmesGzlgRhMwM0qrfTcr+v3poyPvvdyE43aYGMIt8HSUQRCHiSAz9dw8Udv6XCU6Uu0131k9t
l/SAEtZ5kE7Bk2m6z86QNp2sDyNSsh/uyEKgz8BrVnZAv8rsgMNW2+nvqmjSHI0Ze0iut6hwjnPS
qJhyLWxTqC8fZTp7KgQgE0wuz3r9SUo1+aDvF1OcgkBiuLjJ0gzF2iKVNmB8H5+vjcS/KC5QJANV
ww9lWshPeWQPr6NfXWR/WnXOGo8wpD7BC9SuOkTK885XvAtusMLnd4twrxp8nAOuF8ZK0/5vlNWC
GcTCGlhMJRW0tv5cdVEH6bOA2/ySRmDCuI0YYOMKDkdi99evh7KGaIEu+0Y+gvnhu4nlZEwkOpZa
YP/1Sdlul/0u0lz/q8GvuGYr54nazRdBOJTM5lVp1Uzw0NFvG/p5fIy8QKn5JYzI0iEVvQGsAVWG
VHS9cvX9z7aSkgcen06cHXZT/IGnUa2/kS3Cr8AAhZq56Dk7MyT9+U/YBV8EMh/zxvoeBHm5ov1W
YwgjUphLpytoGIct6Ol3wCietpdEZh9CUIeRiacF3zz0oO308Dq1eQWoCyEl3RbRvkrEw8Tbk0Aq
ffd+GpCohED6BMwQOGOVVHtlSRuhooAvM6JA8uf+ONLFW5Vd/Bz3ZHB4U/9QiQbca+EsttjihNzj
LiB400SyoJ4L5J5i8bvrmE2rnK6v5NvVMYE3XdiwzjFRS7ytIgggnuc177fZrJUE5jg2M85pMCMA
aVQInFuk7nfXDWSQElTKNughA7dxGKqF7S/txyW4gwPZMC34ut+T7RUe38VZ/eQTmHnVO7mh7f+a
M7qnlq4NQILClC6oal7IUtwHLkSLciaEdZgtK1aeL4dPwyqQZpSUKYJFnXJ0We7cMr/H3pfiF4qu
+MWxkzUUOBPyVW9n+UHvA/NjwxSI2PwUfXLTi306XzrV7tmNPtkJV9Dq/JV34j57EluYgOdjCTsR
xPiNznoVOgmwWnPkrhze2vqGf3PEse1lSn3ItkK31VfeDzPihwXrLakp5IpcwJL1XPCKO2sma4SD
nXGTwmTBkPKUt2R2XNNCHk9k/ZMQYoR3Yv0i/u0HTZCWDSlXFv1Vz73uugrQcYOyi74ZyX1ConJX
mGbT4gfBx5ybXlJK+cDXJ/HZwPsri3iWIOGAi7Tpug0J8QF3cH5aMrLnDTriR0ET8QjiqhkRJ0im
tsilwAVlujhv2M6uPEDrca9T6IZkK/zOoqjiHb4dCCrTLHvsN7+BDARQlRWT7IkbbGbg/n0r5a+8
k/fZ7uN2reFmEoUneV/j7BL9g6m1hKNZYbn92CVqd5PuwyiSOlfFaaINy2pqqbe5G8Nw7h3za9qz
yratKK60G3QctYfr4UOESzakolfrkeSFOafBm8QUxavqdN7fVLZoer17oM5FU5hmvpuYjepCS+Oa
q8MPsz0T80Px7r37tEUtCJoNFiULu2zBoVSZZtyqi0+sv8Z5HclkyrAFefrjvnd1tzaDbT2++Gc0
9ZL/3grXC1cgEiSqGoZ5ysFsa5u2dKm98r/EpOXs4Nl0lJRir64MCj3+7pSUr61cNnFysuhU9sd+
hckKOUJXffAQtjp4Dw3Lgxabt2L8qUFdXwZ9Wm22IN+5I/7fxgOQpFElR6X3/17b/E7uRrWimr1S
vV6Xkn1T6c8auhc0hIusAPT3YpTa/jqtnBdmVAT8VwVBnVECXpfWbH2rpzkJTxq1LfcU7Ards3z4
OYSoCihna6KXEcclifahlyX6/4iRJSsVJbOacf6zIWLLCQ9jV8tPh8DITeeWfz1XkNRwxEYe10kg
lA89fuZ3ptmcQPVZU1vtNRgkzRIcXEBtG1Tyd7cHUPtbgBADFItuyST3C2dXyP2BBwIKfv5pWm/R
aEfNEtjXSPrvhl8ll+1leVWWqeN5Lfm1Mu9phM+2N17ZgvyJuRQdxfmI6Tu4j7VYz0FCPzSMPx+4
KY1f+Yn3gHVM1cP60aC3nNWC39L5gKj+J2T50xBtyJJAS+SWV2geeX2uP1xX88t8J8QGA4wZX+YL
yyktCgLFlIsGk13A0iIDFxK9eo+3Du9Wg2rN935/v4f1ZvyRDUOUeLCbLeovOZNWqAfdmHRPDy0A
yzKmQbNWHE0S9alN1LuflqYl9aRzDPQAFaC++Nvk5cg7hERxw1w34GafjL3IPu7Jld1b9Ms7xLys
cnVxxK3MrVBmySQrHNwFYzz71IyPrSOkv3Dl4BZrLYWqrdygNaVFczRa/3dUKQmOxbX1S+R9UNvy
oIW8gnJaYmtFtp4g+vMoOEgRDt1Hsx9ZH7eWLrJTGPh+7vaaGORXEqVKhBUX6ac51MYEDdd/Y7I1
8Z4a2uDGQGuBko6O5JFpa7C2h8cOPAC9QmlvUbScV5BujPmEMHC/8ZBgbygAOR3qbECu2/Kq2kN7
JsVXUl7wSe8iaHG82uogsDnru7ZtdIhOMIr8fnAv3K/6QK0ZAZuK891EEGrbZzVLZPJccD4FzQFE
jTr7Btb44XYKE1j8UeeDSmrYRZZw11dp/7vqnjBiFEvDsiNtxNkezKm/BXYePt2EPKSI+O6yltca
54tjCvv7Q6Qf/UFL0akf6gDAQ+AuQJTC4wczR5/Smb1zciy5HUue7b8RvstL5pZrSyci8XD6yDPP
ZBwnTI5SOCs0gm6fY0xPXkDVr+tsu0CjUtvOCb1/bYU+64eW1OYjjoiHGOnaB4In58qbX6ZZAuaw
5CF/VHEoUP2QI/h5p9o26oxT39tzit4O6fH2DEFlLA2V3rCUrQCI75vKM9dviX0CHn9yucqJygZI
5eNfibyX7TrcmNnAeDeK5V5wArTbV1LDeWIRM0WyGvkv/AbgXCMLwUg46a6ZTDd06W9GNjpJdn6q
Fx/NHHQNFn0c0j3GCBk6MVzd/rmzc7FJ9Trh0ye7hEYzbc39zvKE/ZFz7OmegEGyJvK0aRfOYL1a
JInyK6vOqcU292eKjwtOmV5vm97fb/LQeL4C3TI3Vv3N7Tvfe1YXAIJ31McwKHeOvsJt1GWmO0QT
4QpJMtNndJBHpC8WZD2OykPXuOGjQ7c7WfJoHW0YG8o4E3WAJJiFkg11lzR0jeC3KfZIQllFElW1
AduL92ognZZ38CZZ1BW/XpPoIXzcoABTc5XzzYRWmHaEWnZbv2UDQhG2kbduiwRHExZPQ1haK+Cj
4AclZZB1752l7ANSddpPACmsWm1kaSN+RyF00nfVgFqc978djrGWrgMMkI8DIxogOegP2W0DCF8U
dK5DGKUBzkRUhwM1G92x2I7TWW0u3I5WzW+QCgiqxa3bnNPwTtSSVFGCyfjdCJGIGK90ase7YJVp
oxATnTCEy09ITddsiXugzAJNDE94WOB0wkVZ1dJMZr9KeZpcUPhiuuYjPNIePVThZJS/0oyyIavb
j7EOiclhlfb2ffdl9BfnCQT1CfTGNbD4oW68oiNYyljw1MR2hRFkbjetwD8ODYNaOuXYDPPx2Q69
bnJFeblC//2lPWfcVCHqx3aM+8vDWrpGR9D4yhsWJTdm3GsUBPAGIOt2Z3j229FNB1Ppni9Kxnjg
nwC8bIBAer1FA0d2XqYJiygn08BeLkFCcZ4z+/qIifkbIxr/PCa8/zP+MiBl/QcjohC0ODcR8W2A
zeLtyLuZVSOpF4juViBQzJLeHxnWP1lKXUGhQtJ9QMclkisejiHNm8/Q/ew6ykjlN9fb30YnSOun
5srtqwFXDrRmZD31mJTTsEikrTTpvQ0eNDFTDcVpmzp9zCUVBD7Hn8Wn3xTcKRS1KbBL/Mpt+W57
ejGdm+pSsZg+d68dH3CZTjq23z4xiW0UXmjGXcuDIKwbRr1PLWjK+o5pLMEPYNeGt2hgguwTEuUW
Nk5l5/ITLkkoFY2nCwFpGIze080YNiu8fp4CWSuSo+4AjxO2ViuiOSpsBurlmhgN6DPOToUo0mik
iOKv4LxpxmF7hQBcwCSJ/M2ASufSh0OnjbtulGFoVp7ZaO7uGfLxvgSJmGW8plh4jVmBJXnjHVaB
gRTG75fGgWiyitI5St1gtlob9PEK/VIWUjlM/VJRitgbI2ui1nGvK3SvMuW4Sda67Cr1lcOSAHYC
5LMWCw6JEDq5mh9VcU8JCQpWPSqP2kXWW2oSI52NAVywCZih2saEERjGFeouD3Gl7L4tczrv+Fi9
lRQyzoXTtozVgKtxOjkvpL34BOYyHZt4zEwTsDTExWG8+AeSwOZuGMNptSJjrb1mLhByX3IZMNb4
VtnLar4E1sY4UmGq/TgTfYJAU3UUdT9198uPyfdAUS1wfixjpgt4R2PBLQDNzJ40u0dKI1NPZLUt
pf04IT+HqJmCGdsji7WoFiLwpoqpZca7fHoPaIn1aVbrlboEO6n0mrmcs/dNnz5CQ19R5CNk3iDZ
fsTRRpFf5iV0gOjoPhj/n81ZoE3LFNFhGR8IaaAeWtOyx5nIPJ00L1hlU1aaRuyEDagNsU7CZVDC
FrdH+lCZSrB0d5lqhagJcvLKpbwgOKiw3wQTC7vnk59XkDuW0g5mLfpwBUHO6KbxtKpQ82ErR02A
lZYcGc9+Q7Av+Fpf7boRsaT61p42A4sCpS7SgiafuqhEWKfS7LC6gYvWA6wkIFvBVwNmiV3Xr9Xe
RYco5aRuE0KQGAdWekgSZQl+r9qm/4BtqshOH9/be27eIBAcLU3knhyBebSGg/a17Ef4GdI1ALdb
xICCfxRmDLeNIstLsr+7uxdwwDwUiHoadaB0OHEBI9Xy6Y8cPzsfeZ8QqZUI8BmtzOb39iHkEVvt
X8BisjA0RzU58M+7C44FAQCNbBgEhdd+GN+5xmERgvNAGKYc5qOabLmwoq3BpBm1bgnjtpsa8Lio
MJsbj2Rm5PBkIvncowz2M4WAA9K+VIn56wSnEY3KtoZtembiKLQxFgSXJF/N2BT3CVkWZEU8TMVf
TOgDrP/rky7q5/wv8CvdQrh5VjRHZL5HRIVymqeeZaQrI/vMkv1FMY/GnU4CsvB1wVaYOFQ7lJD0
OTROLAwswRcVLypM1lMM5zRe3dKQtRHf2xMgg69ym+6U2av3uIxS0giAJi1NGFHTIqWGBOq24cvY
EArp4ccyFpr7wy0jaP4mqoOSMkUtdt5GX9FXPRjBu0Dsv/O1s107uFs835lJWcfb/m+Uk8cKIcdL
pFq5I2ks1ZeTy/zlpLTzim3TUZE9ziTCG7YHqFKxA4GDibiHxFBPNiUx47NxwSWP/jZ/MzQk/CaF
5fizZwoeFhWdPp6iFiK5/vCxlmGlKREwJwYT9W3TS0V6K7pb/OMjKK+bPkbPsHndB9m2Kv3I3fGp
CH3WhnwkJyArgsLweV3hB5U39Y9F5/m0mxLbs1pve9UelQPEWp+udULwYd1JzpaVL2sfp6959oZT
eKBKYBf+9wY8jJgvcWtwJKMuYvrA24hwnoynXcc/kUSxlFskDoSxhgX39pTiEgRCyMJAg0BWWlk6
kqIl5qK65AFjYYckIdjTo6fje76pZgCpw/SKcPVu54T67RvcCyAnOdRTihXzcGHL+lmdZRvyOEZv
4FHUOtfDb+XAyK7V+NL5dn7AqKEr2wo0GnFNgLlWjNVIeTE+1V2sadIsRwL4WW8j+HusIVbr5JFL
Kmd+djLGz8ryZ9WWtIVTn4IdD2PmFyMjde7ucsypkC9fWqiUI+fMZ7z0mg2LJRDRE0v+J4gzdL/d
uaW95msdCHtpFI3TkBgjwBqDW3Wp1YcBI9uKz3yultcsjOGwYObKZGGiUKA7Aeny+w5sCB3PstgX
6lZhxckF7+PWisXnypokZ9JJsEQkhf5fGtbZ1kFDz0G6vZQJEKvfNnYQrUNVQEt+Lh/Twiogowe1
C+T+B0NNUL0EZKm3XCxA/YVUBGnuWN0INjY48O7QvAOe5QVhPPLUNhqKljG7B8X0fNrwnOD5yxpA
FqZDnKXTP6hdQ05gwMdUTcR0dcn2rA6wOyHZJAnG9xsaMq6mN4zheUDosoS1za5BIjgSb85tzTBY
Rs4x3GVHWeNL7QPmvZbDSO1D3h96moBTkyhwSQ9kGgAT+ogqowHO117A8DhjKfoEfaoorTasj4bu
J9SuE1PUv46p85TVCF0KaRQ1IAQeMtxSSGXSU/wsBc6E7MibUeYlYYjWCExIYFqyS+wBbDDwRVxr
iLhhDeeSIlng9jFSqC0LHb3rNIfWDVK05eEf2SOMQe8VdXpJpsjIvrDUvkIeMy47Lb5SGFlBt695
o0hjLNpk3QyGkqsM9oaex+nfUs/+XBmiy/iLygj3hPSx+RU2d/aNCUOc3D9dBavJzwvbyMZ+NYUx
zx8h3raU7rCst0WfEO12EBeWCDzdzXhfMPYJH+T2IUEETp0f7qlak+vyQKt1oPb/muxqCPG29Akh
IqSQLVpsSPuH1yzdvAes+t5k2ZAOf++56iLgsODwvmWWhkc6lM8LwgUN2O5P8aEllCjLwr2eK+FJ
16PLwp9QDBnhGbEWXk22K9lcUIJ0+TkA55gs5qkRu2ci/Byzdf7YLXlxWKIHzTR7TqH9f7+nHHB7
4YJvoqbYLDIogrMaIQFhbKZfSyAyZxUVy85dohRHxn5bA7nIIkT0IiNNKk8IyPfkVCOUxr4adINd
enDfIC2p7+Y19UiJg9Dmfc3sS2yfaFPTx0EM+EAVP9cJkRk2bBE8X0sF0XX/6YegadEbiIKu9dU8
0LGfGeFYEhHhNwcuzSn8w5hS/hxG1OlY5L0D5I7GlWySDbFmjgat+0feyqHtuIdbkoZR319ErkXJ
6PG24x0TwXmqwGsT3ui2YDb3ZfNAe74gYmS4BQ2iATOTYo4w54hXeLlbEuh9gMjPdwhh2KP5XAmx
HndEb2+yeSWkOoHmwURf4O7F80YAw20/hZm4SHxGB4kSiC/v4+uDkhZU+tcsoA0PwDSc1+gbzR/a
KtxWPIolZ/VTlKrdlgpH1AR2m5AseCz7x0RQROxh4bUlkoIFmxRA82wsF7DWMHcaKzaxDwdz9kGO
bs1nckomcsH1ae27lrRqk6hfNKe8jXN2X97BGo9dwyghApAMPdwxXcDaiwe39iuyyBllfsRYgmyI
mpxwTOTqAGwrH2NdlQg2Si9qUcixbH9vxUUNChgXPkEqpU4e7V4LhwM7cTfOafozYIQnlvySBj51
6F1J9+2pf+yGwMle/wydrk0OzPwzP9KhjC8kaWOBR9WWVI+XiiZGGhMJRy+clIpGaemDLo71gk1f
iAJRVx8QSb97gfCuGC7vSWxRklDpG2X75YGb7gT9OsPZHTzRqBKIEIwzfnDY1aq9TPDL5o4dRuPJ
OqL40NSsWPIUqm9wY0aBy2bmV3MqUIdmyQ+6a5r6dBhYm3vyx8ZO0BknxnmNb88HXzjBq903UDAo
uvkus3Vk5TsfVkdwCtUMxdiMiVrpgXA3CfmJVKzI2y+beFa1ybmMi2UWS64Ylvr0BTnDF4/J8uDw
JJc8kpVT/nk0JMc5L6r+tPdSKVkruSsIu8QycaAZdAyLK4vFPhtLnCJaaOHCHf3SN/pOJR3gg+Dd
KGZyiw+rCzCBByemnEgYwSl5xS93/WSye8LgMb9EAvE/nGK9HF6oGTAXPt80m8hWP0B8uXJJAG8j
0tLErKN8axYwq7rsK/fjdq32dCLrXYIuPUe2QjFInpmGwFXb8tEMB/y4cgHykJ9WwV61bw31g42E
/QFff0EKV8H5F9bZMKdtbwf0/5ksFWjDe5OYuBKx1B4gC4mHrjxxrnq3/VAh6rMCMTsD2sevQHb+
wlyvOVNWHVPCTNCeNP/N2gcY8QrK2AEgcS4ETdVWosXxcxLWqrgU6eA+hdpT/VnUdcQYjnKgGHkV
RolQB+tvKaOQB1y7RDhoLP7jx0dMNGp0ROX3Mjqw1ViYAFugqrzb7pzzkPV1L2wrDTEQrbn1RUni
hCouVQvXtGgkoGO+bfxdDA+PRtaKUsg/u+lV+31DjVa7oObpCIaDcdKDE2JryH9DK+U0bmC+T5fi
CwRbVs/REYw81hJTph8epswXzKZRdZXurjhlsnA0eG0BQs0sq4Fm2Fuqb8G/dGdqDpvr2cTDzDo/
M/GoC7LEcw2JgmLasnw6OKarAxoT9J5BdZQEuj+fVfqkz9os/sBcYD+Wtxkf2bQqQ1GJYzUbIQ83
A5DtAH/6UhTZjHomVkv2fFrvcD8kVEU2n7PiuVhTkIhsmcjz+/YcLWtU8uMojQb7QtyBYZAdOOiA
0y3rTVaoFBNcc5op/sBsJvDMyaqnlj5ptWAgubN9PyaTioubq3+edUYpBdSGK4ZYVlVxdrovUYnX
RYh6GH29SFw5DS/EVaIeRk2deUSwOlmoM6EI1MPbJk8UTB28CtS8KSD0DVXTVNQ8PlMhYBjtUSLA
KQddeDXhHBYklYHiUv4kznqPYMh9H3CSlROotcYIcPIvgAXDKNJgA7nsOSR0cPq6ucgi9V5oOwsR
PAAcbT9zTWs5vQcp0AurIBgCsMbqw4jiQ9bE8dEZu9rfs8UJS8CTccBpjAz7Kpakzc2FKhHIN5zS
+5oRiTUu6ggQr9bkkWCoX2Y4cCTPWVmdIrEAkD/42TcqPmABDFmWxDWJHQkQ548jofrFCM9V/44n
gd8b/EYiZhA8eyPVUmIlJwW9ICPc4w4kVXUUwgsVSJQ2ElzGc9ju5GtJLHpgMrO1OfmqJNL6UNOs
sgUhI7XXjWhQvkZoAjhgjxRHvOUp5LL+6Z92niH9FfKKOAzd4LGbB+EJhx9lAMvUWlGruomx/ARL
kd/jEJS6yjZ73nL3lGVaa0YcvVPxkp5aMNKkDY6X90LUfeHuUQevuVmRk8pxvpxxi226PLy/sIIY
4GPw3jEiXu6o8YUSdpu8hk8AvzGpMBAO49pKnkNeAIH5ehLsd8BkbtRbVLSZc4piGMjcfuWiArqG
QIoR9f59sRxZvehC5SVnls+u5++v5XpWZ+H8UnlI91rDzjGNyYwoFc6n3vnPYUu766nrdEQQGnkA
iY4hNMt/Uzyb40wLBO5cVRX0LiCFfM2c7td61ELTeBQ3n92LOZPvLkqMAL3c8hU5hiBdKeYo2RaN
p/BeAk4X1BEhIBr+xdvBJ/GUf3f95LSoq0LzkmIOOdb0Vvsh2nbxb5rDL5uNfT/quPoO+IAfujWo
qx0C6tooYjOJBpDdxCJ9AxUk/MCpZNYHoE+bZLk0lWdru27LITMduEMDS78YhkSfOGQblowo+QNY
LK3XgZRGod5Dla4v9QiG1zcUediC+Hz5qQRNd7VQudGfs8/AwfJvNsyt6yCKwugCxaT9tFcikLJH
2JHa704+GAcr9C6v9MnBnFgEluOYpgkUXMbaABzyibasYNMdx2SjrHe9UuMHmES1UR6ACbeqU8fo
QwW0eSSGkGMwYqllqhUULATbNsYKk5ffB4lRNa/u/c1W4r1+QyEXlbiJfj/n9RN4EQBWMAqvmnXa
4LqvmNLvGHRb312ah0IKmD1SocLhUcGujc9u/8LDA0dDaFObC+In4ODgTDNzeNAcHwZyQ0rCNdvV
b4QmJobvsJrbkPJuW+J68yXIEB53M76I1clDeQXy9pC5+qJXit4St1t3LExqkJMHS/JENtkgBOOF
0DIMOqshl/9tl5zDHifPiiR6WE7cKzsQ72H5eS5eX7qbUWLJ+nZf2QxPNtyi0CGwPJQCyUXBbhcR
P5xYDsxdW7S6CjBB2wKwWjgA/Gcj3Gv3LJyZYMl3oP3pj7Jg5CfaShK0Psfzr7gtEW3j1y0Zlr1c
rJZrdKmNt4bpxqDG9RC0EVEZN9tWQiUeMCJmZlqgpb5ibvyX8Zuqhy9iBy0CI2SvhIH/HXhRDcIj
vDQHXliZ+UYgliZI3K9wmmMM+VpRil0twL+5OEEHhKhOqMFgEoO+6LM2vTdRmM0I64WHnSc7tLM7
4CReLWFqdrw9eusJYNPDNQHK1nTDbxNsSq7h1Mrw7p6FwDFCUwO6i6nJ7/GWJdnq2Hx9CzieGTje
1IumgpdwN30jMG9hyPZVApasIstNILq+D+TBkPUwo7dlfhwHRFzL604fopsCtNTvQocknfUuWYCW
68Ty8C57mzhDVTr1+Z5bBiEXNSvbc4HJlj4PGc1Q0WaDrJB0T5lx4In2Z66nhZEc3mKaxifMN67m
h1U5ugssqpIcgtdsaYL+sYOmbHRJhSWP6/9u0VAzmLL695R8Wq68c1owUIWdtILylBp21GqMMv+h
vRlZyO/yh7v/kw43JHGU8FxkM5LqdVmEcB8CR5cCfP0GfcSnhAaUFKe4bS+4hpEITunqpLZ8pSrv
SgTiOcJyRkaVWy9auqCZLwr+tgVe6h/rAEo4tlXDQ/yjVar0UQulIFoaPV+EAs97M4unN6egZ7/8
AZbhMgShhkMYQmNC9RZQyATHbi1zfv0s68FUh6GvqsnLzOQvWgW0Cme3YX2N83K2sth+qi+FoHfM
2p88cL0SQly6XPrXpP+HUwSqkCy+StF8qHdZTbWe4aunufk7J9MdpHIT9TUcgNVcq36/7LKzGKS4
A9sD6a9Ix7GbUf7+m7+wKAJdvZhQhUJgdlJZhs9aX3h0mfsv2MWqx4bgryby2pVctqh/rj6ZT6zi
71ESZbSQswvUSAZfirvBLH5gvX5dN5Vp+3CttGa8a2HxyHaHH/GQ/11+7dxusnxzLBaio0USlaGJ
S6H/CvnJzEIPpkE+IXnzTN/8FhkxSIu+hkZlFXOd7HFZKjHZJGQwZzs/0hZH/lSWwgGwyALZddKC
0zMTCMhPPOTWyS5hJp5F8uIbWp+1Omi0/LoDHZ/jNDcy/ryMYbiehnRKhjlSM8bfLVKwaYdRF8+t
s1c0zFzFShjpgZf1bj+kw/wFzbUm4PGepbL3DHDXYgEvs7koNxekcGMNfviJH3J/t+62yjkC/yDm
rK/sW1g6D6Lwf6Q+FCdfOPgisD9W6l5a5YBvRfikRnYFVwFDJxTcCcyaFrpaJ+qN57pEnfJzeCjB
IbUE7QKNtWe0GQcSv14PhY0FoScGkdp0GCijm+SQB0V3O6q2c8lb63LRRAt4ZC+IHG2oWHso90fN
c0IePZ+b6ljKPVgesOmMNScFjRWrl6z/AZPPCNgcpwv/4XLLyGQmS9WGU91p3q+iQOUt77n3ZnCI
VpplUYaOdSk7FxZU05QZdv//i+IFRu6Quu3Gho6xdiE/UPjnXWJKg3Z0IZgDUYIkzavRgG9Wm7OZ
Pm4l8TVw32/rdRGgH4uNOEX2l0r9SVNCtMXUdmqd2L0t/lzBW0pgS+vdGtuSDy1hFXScAl3yrDA1
VBEXERB9qwJCvlO5ZNGufxu+pJT40QVxBsHwfnTf2nTk6ODnRnMOo3DVyaNTuA8UewopCePxYnx8
9/naZ4FPNcplCveQ3zkWwq2X+eydP+Ir4rbTZqq8Hdny9tO4x4LdYGk6aBoDK8DkXe0w6Wb/H8Ei
O6Jo/FwcM/m9TBl8rxDxZL2Do9a8oBXm7ZhBTsCle5hqJk8FI268QzFV3MOILle4W35SPthDVWbM
LdT2SRL4te3l2q1KihTQW/TvFCqC7qJUoA6aaozKmvyYqAQJlZIa8bCGIVcAhNDiLvrFNWdG0Ir7
v9Sl/kt/gYxAWX4pyrWJwnbguB60KimZzQ+FBNAe5sYVVz0oURd84WC6g7jGi5LEnRnx8/+wYyrM
cFqf3gVSQZEm7QM23mEkSb39tPy8M0KoZIrCQ6BhaESWUk/7ha+MHLFyNsKCV7UicUkxcgnWnsvw
l8CGS/YnEFq+BJRSZVkIzt0iUTqPmyb7KhO05DJ7QphuXVK7o9RVttoxsp0KpqPBr+sjo98Mper9
MRo7g3tICWO1UU4tK2ioDnwzsOCPsoEoF+XfeyddNOQd5sLOAzPwlgJFbkVCJUF+wzCm9Nk2qw3A
BN5+iT+sMZut/FZqb28HXLfxXCUkW4nOZmtNI2qv3A44zt6z76AHojsSQni+HltSUThq0vIUEBpd
oNkp9IGcEk5t1uB/jostnue2k1orUpAUCfxkm9FS9+Joi8bxneeWZW4TiNiHZOnNPjbdJ1Wm+iJy
bN28FjHeW2ibH7eYbTIQAXEqdcewHY2lMsYoJOi8YRLxD2Ey5jgwHpulczmChU7XJ2tMq+xtqyF8
waaq1p736yzzKPLnav5aYiVWGARXiNts4JhS+NeUlTif+DI6fnxIb7nD/7UFBnLHJAOSQG6XNB7j
Qpx1wYa5U/UTYvjWN1jR54xqyKCdeJX+8l8gzagXpx3r/ll5CGONinWkzU6LXhomHoCBriJQaUkT
7ee5KxUub9yUbghrbKPc2MLCuSw1sPUgpq63FlwnRFbnDJYQQ8KSk6xVISt1kw9FLvKdTmx8maJV
aGxjuMwyw50b2VhGtB6O6/gq6aIHlrXerU8DNzZaV/zUGraaFi6PN0surCBUDp8heikNoHIjPj1E
u9LjsgFXBPYpsQ7NUM9d3LR2cvyv0pqsaeIL2OVb/3aFkY8PlaCaqGhFZIHwNvei8inFwkYrEq7/
nTHWH45+kbyGqhmdcxY4HxNcKZzVSiJnBMhNTDttvL4xRR4G1dqJWbGZkE1DUdDJ5jj0mNw7t/ig
VjJ46WTh+oMlO0XjVOIY201NNLQ7AFAn1eBOIHTIQK3tohQl2hsjDXHQNb4ASQmZDOVwq0fSTSh3
/M0PsRqRIq2vN49CzOnXedW924NIJm9WRQUlVUcN/HfpEjk38BsJdShDq0TyNYEowxop4ogEjNtj
Q7fPg7GRDvQ2lI1H7LrUr3A5r0RQWp9kQIUncEaOjf6QAv1EORXLMSijK+AH4LO+NZfR70IH4L2l
Elco2pwESdqHTskd9jyDipmzN8eNotXfuTaOH2j5XJDeLzVqQRJBt96fWHDuUQZGADMboXTbpH3k
dfIn2c9SsOQy1WGaKafTBHYaWr2WJuIIjzEEPwF1JrPSPUoAIX4XK/ohflmsYnc7ko1QAuoWxVhN
Rmgsx0w6gJ3X2SWHHNp9vISAiDX28+OuQEWgPtDg+oZpYo34uneaiMy4xMyvM0FJm+Ac0AIIA8kB
Tkr9mc/sLsYwgudYDD0AO7OnMr58xHzJRe1WRvylZpvwfGPKnLK/22UGCL3nHZNDza4mqvfe4sej
iIXn0s6wS8F90CDkvBcbJXG9rWzp6AmKsIiRd3Xgei+wYXbbo1GHX7dHZAUzx/bbJMtzgbvUUe9f
hyBxAZqrE5rtuEDstIzkhwqNeM4PRNPugxrJt3jXz74Ic6s1pZU6yUqEKWZHC+usNX2qNcKZBdVG
n6lJszuH4sP+OmayPvA6LtkG7ibj3USHxB69pYTpuNtH3pA6T80GX8BMmBDZdP1YUbNJ7dNgTkA2
uYDTHrxzV3/ze1R0nyn+mrbrxtnB0ysbsO4VzQFcwnMcc8/tYNfk/6bpaMfwmnXW7XUD2CclfuBh
Gf1LJdkn6c3JPJS/P5YenpopzJ5RY3CiOUoE/NaA21j9gDOoXuBVbdxPLp6JAjZKg6tyxuWtV3B/
V7RwkLAGm+xd9YB9DbjRy1xyXZ2+R27yEZMXR9XBN1WA4Y6Ev5wyFBYFF7OcXKA9MYHRiZpEn6J4
t4p8+ffvQKnBp+CuthZANkkuPuYTEPsgrJop6lp5c64fudV0GtGbiqiMoV3B4BoMc5ZmAn5Nsrg3
x9KvhQn2SNYFqlw/VlG0H9QzFgl/GQeZnpg1cKWvV8cY00ocpYVmnLC++m9tI4pbT+Ru9xNPNVYC
uS0OSy8NpZA4Pyb/6YCwZJp8ocnun9PwVNsfNLFU8uexGgRvjFehONWlSPfEXMZ082d+uztDRRlz
5y+7K+r1MORsxSfEZJa7hdl+d0bp3qt1oD55yTb13ihwUOhQDZJ059gxeNET3vW/Z/ICEasZTkm2
RgAA5RWIj09/9jwijOzAAmU/okGlfqZAXh7upmvav2JzpQjxlzE77sS9ByfeEgr0qJ4L9R9srFzG
8TaPKz0gH15Z1YG/76TC0nsvj4nFwN5VZmE0NdZpCuSO9vaHyXoK+Sv3oAmSusVCt0YdPXOxEqnN
G3pzv6KOTKYdxwQgd6Vn89QQUZ3nFex3/sz29z2TAlZGPUCJI095mcWmF9TpFMmJfyoJViWeiM5P
Yt3FYsPFg7F5uhiB+G35OsGF+PZ5jxWE7p2EN582yKOt98froGOj38S2FP+8Z2KmiSJ/0Cwo6eeu
E6PhOyYy+HDWMdUQSKQTsz+967B49yncPumUIBDsfARH6cOjAW0uMb5Iu2jG50Xu895Jm7NdJCDh
2do9pv4ri+72ls6H0Lw76J7czNXcATscY/abVzeDwPeBjlF8tTJ02O2gvgEa5rOs6VcCw5vf1W1k
rvlUcmsyGnDL/Hw4I3XuVCxYlkrn8zIhi7S38SLPa9VQ3BiwBJxK0c2JnfpzDE2YWSwKosptVslI
GNyxz6KYXVx1x/ti6+GlT1opsibz3ra4XaNvUTseIPDy8P0GZzvkvFTDy0FH/LfDMmmpEFAeUus0
a4Pp5pU/2CqnDXmUDK33o6FsdR5g2v5xpDsGiOvB7EboMYlEdOi4pYalnGdxA+bDbLXT/luM3KtW
tH/HX6/kBfusvUj7eZG0b7ffwO44fnXRC608DVdMwLQz+5r0EMj0SXGd06/mKX+wugt2clX3waKE
YzJPjokxlAau7cYeScAnOumyGaPIdrY83q0QLkGivlhBKM4DSq40OBoLAKiofW7lgJwK5nCzNcPq
Di/Q+8I/uD4nDAxvSkKr4AHRiWY0Gob+mbGFcIip3f1m6Su+VMjwgBymQB2jLMEwh5nipMd0Ug1b
xbaTURpsIzqmtv+cdO5Zs8B+AS5vP+uOVfp9oihAIPdr1KebIoiQMz0cILno6ieKyRy2cR9odqhw
riAC9iPoGJipV8ecX9UGTNtIIGRXNRecyMs6T1sY4G6qJCJPXwkjI9NrUEr1OMu5tN3FZGQOcnXW
KRqXw4mZLV6VpEv05cVflnye36EDPF6dBoEnpFJfNOBAlBDbgPok495UpkgISU4ZiII6HluswpON
RXktfzAyRXWX8GaJJ8GONCX7r8TmWs0ntp66A+LcvqkdL+l/7lcEMdI/4s9zooSeKR6tfbXeWk1/
HKkn9JInDSx2x4nYBFYNOkl7TmsDpMDefdyTp57Whlqs3LiN7VlbcXOuMD9qxudpcdVcFILU49QP
QGkFeHdkZztKsOMt8RPPo3Z5l7Qpn9soSbuGFP5/RBfL3hsJ+YV102h0LS3R9fjSmg/qv0FVq0ww
4LSWy3MHe52IJ8WqHC2miJCVwLg0MYQVVg8Uck7QlwfLyp0ox5AVKcgRFTrlyWcY7f+NKIMNHmY8
yGe3CJHas0LZSQD0As7iKC3XKAh/glY4pw1xy5nUU9ThIDLWtHH/0HmgKi5NFCHzPudIOmn7gbxY
7OJrCyShX8M3Ut1WQDJwGlsHf1Nmte3marudZOhsV8XViXZvMc427J/MnhCmQs3A6GRC7eBJ9oFY
Ve3t1TrKSJj8n3rBgs5nv09c1gosMkLl0kL5R5WKvbWVjvuVNuadK1DuJ0y8O0ZxaUcGhHgaz0O1
FOgYfV6ZgXZVKgnKMlja75QCjrEPFyM1SXR3/CZmQ5Nor0pqJEdThOTQYTtpTnvyJPW1vB3AIDoi
Zk3WAclEVeitZ0BR8QoCqSDSNrtmd4RKFr9iYTlgA3dIynbY9DMzYp7k6I4AysT4FxOBpV1Wvbgm
yxtQFxGFhaqldpIDplOoiX3yqh8kwJp/dpBxGqcSChvEwcq8ox+8Rah5jmgGG3mSpxzKgK1d3o2v
OUVgvNdwavhH0cls8xRhKt/fKCV321Ubyi2luWxvsITcLoO1z5H8wxGHwvxpL1eyM3hFa2n90XeT
zxjOfQ4VnkfbzqHtx5L1hBlNlOJ+Nnz9CmqpppZ+LYtH0Ax/4SDBdyxkFB+aK+dNOIcwAxqWbUD7
wLtPiN2rGrV98qORzPMy5aC5FB7r4nyys7dJa3rdZ4sMg2X2HHf5tMXVME67Wz6KWviWsUwA3six
Nw8db/SOM8Z8bjThSPlq84MseSrMlXqs30fhw+QpONF1LrzgBkA30lUczZqwO9U8XFeYechJMlIQ
z1xYP3MOplLJBpRWWttEq9xMtGAuRdON3eNr5dTN7Sr/TNR+r6Q/nIIzNSDysQS5ABp6JmKxN0gj
YdCxXEvENWu+nxv4s0n9Kv2FUMTFn+4KhMTpigKSOF+oIzvxPQRSPRJEbOgTIuHqpmXVeJGKVBb7
zapF/fldTCj9HuBnLc3NRoN4UWb6UwogSjPIDkhm2QZnQdG1ID6bdru3ufSIBXdMfrUpfrSxL4SK
jJsHcN/daQ7fIqogQfBUiuDWRKrjJPwD85e1ZgV0AsUIwb08/PriWcFViuiXlqJw+TRbxvRaQRsq
nNbI//qpUg1F6Jl2RG3JAZFtZowWcoNGYrPdrOgWeMdNzt/X1DeHu+hVxhCKGCz74dbI3UUS9tf8
tpaPUigdltMXVUhFqbpxhoFyfAxkGqd+qWPjcUSjt9+L0FMURTQEsvcZWkfRno3Vu0iS1HSX8CRD
W+4F/LGsWaZl7PsmMVCc7GbhAurYtHGkIVOfFrE1vEH3aSDnjgIP+OKJPb1KU5BTEvCU/ictQJ8C
2odN+VnKoaLmJ9pCSEIobIPFfJULVcFQgLeLu9N4eAIDAAXGQk0gBYlENbovBk74+WhtXCr8D2EA
tO/KRo29oKX6Uwk6GUUvb4kTVvu+8NtA2zkP8YfVAt/QXdWTuf3+lIL9fl4oGJP6pYsPzkpPPwM9
R/OTVPqUT98h43ZNHVvUotfubKtm0tJH2h22729KYA+dd7PoPC8QzSLtnKuAyB6Maz72iflTUxLN
+spdCkf1bkt7GJIBC25Sg4A5929DA4MzJatqiFDWgBAqZIDmBxq4Cmt83sC3sM99G5By9ieHCXaw
MgLHKg7RCyXSx2z/ygi/7N3ffu7RWoiTkU3agd2/wcTZILl/0ljyK459zQToe1exOwyshTGIga7B
3GFEXP6cCSMav8bi9/OsXSOWrUXUtAt2PKr0Yjxo+V/2J2njHVhs1yBH7lYAnC0QuDWhhBSFOaUS
Joy4uNp3DfRRV394skLEvFH4IErHCn4aySMJdk/IyZzouvmRKJsR///n8TtB2Oz29LwVkNAReHkc
/GH2G3C+PXgVSIVDWPTmeBx6JNHWBjBkoJ63TmUcUzbRZVWabagLfUu/oS2+Oiz+wNumPXyWSIUx
UxqhZVwzmSrb/FGCiK+pD915KlGMQ87EaPljWdaUvGqqDgd11MfsIV03oFbsr72sf5xZk0fu3rMu
TbfC8llpn4WBsbViGRP0kFZQ0wbExRu37xMOq0lg6IRubcvKdiWxUqFkH8/xpo3kCHXAm6kSTb2c
5gE/4O7XtzoB8FhJiF8eQfcE4DguN3gz3vyUWZUuXr9QrCQvHkMXshvSanzSBpL6IjaoazDh0gGV
52Z8WNeUgUfqOFpiw/iAsISFufvbIiocrLceKvizRm9/zEZoF4vHOtuCK6ovLXTRX7cM0LOZzI/w
8btL4soGMOomB4D+vEHSmxdMGj/MF+V/AIrutUBfuL/mSg2TVt676RqqLe/kwXbwKp9oQfg1Bonl
33cgJcD7P04bR50M81LHQhAl4imLIlLyujRXw/oXO3UrXjw7+kuMRoPFZP1ROibox1/YyLFTngIY
5THagTm7BaG54oE1qLI9ejpH6niJ1CzZnZY+1SVYOsRyOt0VPpCR2jFNfcIatPhQOkZHajpqLGU9
B4PA9NECpsCMgg3H9pqAVSUIiSLZvkeI+wOLcKCgZRlQF3qR/XgQuCdYiM8TI6XH2QNOcCRBZiZr
sedLz9wKAQrlNN382SwmYpYK0YGdtCvtyAo+7erkE2xjasQNOSjRkcmtRHi9IbQ2WWOHjSzpYDXz
vrZ9r//TFpiaL6JRvjbDKIVyYBK2s+hI4cI22smEPL0A3EvaozFLY6yHbLBEn8bPhDctGZEtSlhU
mhDBjxbr/+ZQURUS38xk9DF4vNUNpWgLVvAQZI1GcWYFk/euiaaRcf8tnz44zf4TGsjzHL48gASX
rKZX2yS50O4PvVp4pR0/fFU3D7kzX+pXyTDd4fqM8sAx6Pc7O31Exf3AmZX4Cqf/bNImqeEC2dbu
PCmPF42f4Lmth1z14VapgfMnA0z1E9XHemkmOi9J5Vc5d9/fftF1XLNy955wJ9DUvPTSd+O/gqT3
8aWtxUKy57ygBFCnROSktgfMBbPT1JKBIKoD1r5kVX9jKaoiLi6wHk7SrfhLlnwK22dcUZMH4NQg
i5L1gKIGo8A6a9OdhVd5yJ/VHPdOLRrTprX+xcFJ8P4HZKNoyH8oV1/IrlEW1BIM/LXudLWWgJuc
f9UibOG3y5C6gnwpdS4gNTre5373m8eQHgXgj7weWPjjn00/a6vhHiZ8iu9YYXURJC+whN19dIQA
8j4qmrB5RszW/YvZBOv2akvljJrIT7hgITXHhb05cW1Tj4aQyjz0SaOzLFps+69wD6Md/CCf+iXI
5F+9/fhwXv+9+vuXWLzJ/JRtBjcCvJELg39KqhsQuzX+nI42+lc5BLSUm/jpwda8vhmN5jgkxoJc
bbWZZpDxwrls60yU7m4PfakcP2KiHCxf1jaT2xM6tkmjy9IMcdzUDj/x6sP1zxRqmICUDIUjmAkl
t+KZ4dt9mi2NfW8y5DkKkOzpAi/GCLz1iCFjwMyqOuay7kVCsrHIpADQ/Fn6XiYEnOmbfBTQvzpK
rudTxtaFGy7/GMxKgHAexYriOePRsL1AM23+G17kv4/JMstOtcoY5YsiyeHc/rlh1+mJQq7q0Xvb
xwytO1+7ybpnMo+bFz3n/orp++zW76a2rmiTDrvoC6YPCkDMpB9eoL7FI/PgHoRtA6vNaieg3iRn
mLKHEtLlrhe750YWM+vImN/JrGCZVKQgclKd1ASXxw85vetgYcYMUhJz4GnN+Vf7z4Z2p7q2Mc2y
tRaP3Qxj4ZFzn2piCQG20fQ3kabDiU27zwYsBX3ewyAU5XNQ3y5lrCYIDP+Y6l1F1pU3q7mlMcG0
EEoC+pePMe3qitzpnjjhSMje6gV3zM2+77pHQj7s1P9fpuuP1ilSsQMyQEsnSoYBx+XhvxQ2ku01
/7ju1nVOprxMGCs8Nmpz1zvBx/E/Vlq6QSf3aGfg9EEQH114QSDqqAlQW0xvV9nViIGuJ54l2q9/
eKFpTDQoa9Sj6npZ2FlHyJoRC7gtKhfKCgMlx5aCE94j+KtEfiCnbu8DVCbqjrRdKm8a57Q4I1OC
or0ObGHZuuIC2baj+JCul0hhv4SnJqe2LCDy8Wf4iWNTG8qPg10D8qhI7zV693P+m6Pv6mNR5Hvg
SD6DzhkrHR6znq5gh65ouufdhNSzP27Lgd6fNo5iJjEDTf2LWoNjTZkQMdiSzS8sOPffSivUsBB5
eNXfeTnkbLrTrCLyqQb0bq/3MHUl+u0mWxVQYr3Rdjc9LW6Y+V6po7bKOrqcygOtQEKp7bWhLK+s
P/9u6NiY3zqB1zoY6t15IrYq6Da3tbYmd66T/YwVnCWHcuv08gWUsdCd+J9TIzVFl8WgkA7/Q7tl
22GPrNe7OtMvn3FqYU1GHzmbKJgFwGMKLLwnYFQ/QJJ30zMpBR8+3of6Fkvj11F+z+TdFER9RCtH
0z0inxolut5iPXECPkmVVE3uv9RE0CDoyPbMfVNFtHFln7i7tUltOhwkGNnUX4hwOoX1RuTlI1rj
qpvYLELS5glCoH0nUdXqgGpV9Peunr4XLBo/lw6NpVdM4TfsOVodAmOrqgjgMGptKKAr0KgwJMbK
n4ZQpLYeoRPKK9GWONrq1ijJOD3BpcEyRJ1MwgtOGyNRBCREewvcSg+zG39N3Sa56ZES8hE+alMQ
+kLHN1ecj801ubp80JcR9hvSlMd0x6IHzXrWo5YdFrWtKryQmTa3mzsROzRlIw+Nbvhc5OPbQ4CX
oWGGk1fpSjGoYDvEb008WNuDsPP+PCMUjzOj59XKfsctLgR8uw3X47wp969iQQGMBn+7PpRzqrol
06iBtg45RQ8q2RwuQI4O4oBfce1iAWH4t4V5f0wtjeffJ0HP9cJMiPMA66NWMQo3lt0Y8/vVuXrJ
KLzRL6uSRIH+vEvo9a6zOfunUlws49QHYujSa5fc06qmPMs3YpFBROt03GCe2KqNIQDa/SS6E8h/
1edd0m54hzyMqSMjezry6FBMc6MJRKuPf+UcapTo+sXb9va2xC/WmdMtUr53vhB8pNwECy1+N1ai
FDLxsNLkSqNILPhUtXHLZyI6tLyn6KvSP7H9l0BraUxSSFtupcDYdi1wUGCjvdHFVqDdRbx4m3Ui
JkNmzq6wQXLXWbnwWdm9e08lINMTF9BoxWy7P5/YlfsYdfxKd8FzDP0Ykm13fbLqEgDMiNzA7Pvx
gMhued7w/p6MogUd17fA522wAwzj8PfYFBCF4kiSOxVv7dvcXxvadhubwTQHHXf0BHAg94W+Npr+
msNYLNWHIYaWW1muekXutnUoZGVHXg5Ow3cYzgePfPJdPp76Zd6LqGYArk82j/iv1r92VI/7t3Ju
1n8bYIdevjAQ0YgCCW9znHstJlBqbJPzBVKgY8DvMDdPN4T0A5tXH3gw0yd3UIub668ledwyNai3
RxJpMwFOyhqdf/G2PMDiIZvxaSNjIzPbxTjMMS3lh8DRCSTQnMNl/9hSicqz05nsZ//GRnhBqMGz
VyWDHapbO3Q/q2THfx5AWv+kqyCcmKvasBZ/i32p9BEHT3LVQJn8JL0Uxx3nf3iyvPN1gQXRKppV
T0pmDkktd8nvrxFtKVSQUf+hQRg5G+8fqlSbyHxiNWNyNknPXrfGcLOY9a8HaupU29J5H2THrZAr
En86OmDi8eQ3EJDw/ey3aF2E3XOgyNPqjGcx38tjAfF/iHZwwpXvxIlzUoZC/symKHef7EsNsrF4
KJhYsQMR4cdVz7KSHyK6TgBqN/hs1PBbUu3b6NSKX3R+LaBSuubqXUtiGNo6g59BmK9e3VuC0Vqi
PQTW1QdTPFbyTXXZsllbAVUfwzguHu+NPbX5cm3nPZmVw3jDP/Jbok2cW3lYFlwOgYvT6CyI8E8Q
3E8n2aIg+JWwev6+8HL3HbcOCxOe5Fb6iC0MgRpFGqrvRTlYzgnFJsd0MF0ZMnVIwJxLamxyqlFl
ZXUK26wxxb7zIxOSProFcuctI+Okdc0HYixtqY0pmdUH7UnPVTaZXe7eh85nkTXkkEpCC5P7Fpxd
ngv2qfkI3kbX2W1PfHO2kaCrzWoBHaZu7JhNBYEdMJAI+eHyf0r8ofdG57Ufzb5fo76ewKBv57uG
19OwCcZ0aOOFLH+EptXkoFx4HK+jsE4z/lmQvRQ5ILPxX52FMWgzBroqsgrOt73EJ7OVWaXBNf2s
gnvjKAgg0A7zdgc6PTGAoM9PzUzpGrOytcusOp0ObMpO12rOoYIq9f9QSTUioleC4qYzXj30chXo
IuGuDwKNYGO/nsnopUbSp/2IwxclVi2zQygOorYeHaV/vhGEavzvonZicAFHG41EC8jE13Q2rBs0
vp9PMl8OHa4dOs17n4GfB0iBXvpo9ZwcstNFGWBLUN/Z8XIYToiVeDmd3RA1JMJj/dIAqTx/5gm1
pdyIhCDcRh0GLjMHoArtbiIKukhaB5Ks7cbnshufeFkyfcEzdqpivcMoTKDEd8kU+YMvNudPrKYk
z62lV29brV563TxmT98FoM1gKhZTwe/TIk3zuBmlnx0ZMKLnuScHC7gcShUSn9j9XfsKj2i2n0Vu
VibfiAqC/FAPiy159MJi3Qu0Tqeb57JVFq7hQz9lVSWDNX0qzp9LATZFDa+if5zKRkjHu3XZRodE
uPpre4JCYv7Zh3P+87wp85pUmsXqeZTNcT4qLmvoYE0Eald6SyZwmjbf1FbYNtLWBPcR4BpgsdS2
xMxY+USTp0irwaI6Nt5+DBpbPbl4UNchsdArV4+pOThZZgLbEknMi22TPYWMS5D8vHXtOup7ikB8
Px0Wpgy5dHJVsJ4FiXsTrmWRmRMrXUuToOGemW2tHo4HoQ+K9qjKopdPG4H58dRfsdYHvR5szpvp
H41tw1N82uo0FmJwin4SG5abDPq7WDwrjjwdoNBPLTs7Ni5qA+NkhYePTPGrsqzYLq+i5UjQqBmI
A30xr0qnpxUxqw3D8AQcvYjOICT+9PvegY/8FBLIxucISU/BcTznBirDGKaRG7gDq/cXVVa9HfWW
EBDAmnRw+fNddgUPtAhklkvly4awih4HCAUCCpzFRnPMx7HHmJCfnE053+tm5RKjAkiVpP3StBar
8ZlVfvhB5oACuZvmvfGnlstkFxTgvi9b5DDd65GhkU/pBtDFOaVN5NgF3vMiYydZpnFq2R81PSpr
Ln4eJZ+DU4Wx9qVcKnPGkQz1cdhjjBPA8apeClvij/KS5Cab6Ql4cPqLTIT25QT+GEo5VWwJ6ODe
6sZhMltVYNdkImzHniYugiPTPeBTRwuuRFeqdfqepx6JZjONwIvopp2//Kj9V5I+hRJhSGY6HolZ
6SH+6JbZi1jdF/JKRUpbqYXDwQlgCmg7sYMHaJpasF8jrLE7k9PbFe0nCOF8BpYsLjTAFnLRGCAa
CIK0ArDpZyFcQPuRb58TRvLJ6XDZjVZdpbirrP850szoptJ5lb4MMqOuaIiRF+hoSXvlkl9Omx1d
Q6EHksAv4e+tznoNpjszW5ObAsStFa/6azzpNJFsHbE4us6OBcQ4dlSPH+IUL9VLHRJArLxY9nR8
KkjofnsAMIlEfscsBTGdKYyU0/xv3iZ+RhL+1hN8xxiqJw0qZDnlcHBPLllcivbLA9oUxz0GHEGL
h2vf7WyL4og2ZMtHKw3OHoWcnwVp/OZ4e7NSf9byrpiaKLH9ghdhiHdALJun7DeO5Je+vwdUVdl2
RQJkTqy8C9uyOb33OzG5JPY8IJl4oswzMVAMb3WqqyQmIPTe9zfmxIwRih4/0FJizu8LMOEjo1Km
2yt6KaFtNulyEUGf5zriJjBJOSM6RfaOMgbfd4h9IYTDTu2gIbpwssVoE1HUGbY2H5TRIuzA9rnZ
I4bGrxZEJ6DKVTWBwWWO7ZVc8LbBCEdOInsp3pbceSqGEJxKiRW9DvlfQewBJ8XwNhN8SZS5N/W/
g14qT/CCdzMT7ir5SZt2TtCFq9GoJZIaz4X1YcfA8ZHMgarW/0IUmJf5A3xtz4XeeAYrtH7LKy94
9rYVCgx0QLSG/BHh3noLkeM7FWamiOBivY0Es0KbZiKjal+bv61IICdF8NX3WwrePA2liki/Ve8N
V7nLn92Y/jXP1RRSq/F9tkwKDJ7Sow69/ffDddmR2igj634+zeRf0lMcGxQa/xKfxj+JR2EdbXqS
CgiQKrUp7ndUlaCvcZS9yT/uZ2/EsWtCHscEoP+7EpHUE9Q0tLZuzsXYUJrXPtsmVFHpVDsCviyp
q3ug67/HRpoEaF5F0zjW5UjV8DLx9ZBkRkdeyX07X/0xWELjNY0Yf1A7ttYZgkycnKc1Iu8jz2PB
cGfVjriwVlUY5IgzBBmjm/Fxx2RXlizNR6NSS/0kChkmvbmswhCkrbZXTdqWOm8p7bdX4IoHa7K4
CswfyQjV4rstrrGbyg6+HcQiaOh1ov1cxBjMrOFmPbztgAsHX3JK7051aNYxCviidXXM450fzHu8
PvbT+1HsJ7VjRIgCRC3Ht7kP0OE/0NsRC0dLXLd9Q0mAJ283mA8DNdud9u1RPvhu9HYBhGMNYeXD
9GbylvYsF11WNoa82mBesxJeXURuXTRanfXXvGZJ7nHVtKkEwBtTNxCgr8IHUUbvj+3nze7aL2mk
c1rBET7wT/wxDo4zMiDlQ/+3eyZQXPazIpPUKioI4/rRx6P5+k53LPWW6wbaurKXZae6aOLgTpQT
vlhcbgcuOq2wTKw8WpeSFs41VJMBKS/oYk5ui9YcSsajhQ+wHAptPoEC+claroMBx7D/MP7qTxlF
aUyrEeRUu+lXUBK5nzVaMLIuSst42A4xzup7GeQ0sE5GBd3JPSAjFzc0lK6LXRTE6iveDa0aMu2v
sY+/XN2k+g4Xy/DM2su+qQapoWwEBPN5Ta/COhLj/sz/QskpuRKwGFwRUe2Alv49L0LXHGMz+7T7
zJVnNy0ontmdxZ2NHSH29uOQmElzTVod7iWBzYXk3qc9lXsMk61tfLcDO2LAMB3qw7G1XpPhfMss
cZ2UBkp9dJgadD1RcP4ZFdJ7Ydm+BVERGF1yj7407D9Iz+SqSyUgYU++EaYsq95zQ9g5/awQICve
Cc/2LSEpeVv5HlXVRC6fViDAN0yNGPA+0KDXFMoDr8vYRUUQDkO9Y/tt3KlUtTQXUdDAFClmpAL6
9Yl/dlFx+uovKJUK6n39E91Mtiy0rYc+NFdHEoVVeALVJjihmV3SEh8ePknhSRbuMOWpXGD22D4n
VkU/nW3i4Bp6dLWtIUOFpDc6avNRe6sqJ3/AaAh52k1usOzhCk3tm9t6vO378PG9xLiIC7N2VzXB
Nz6U/cBWaGnqBJH/9D9ga8lxO3CzBgvB4usdk2tPJn+aFgMAeov39K+VWVgLhwODwcev5hhw4zHH
yISbsf3sBK6JTT4iUmTfArezwIvvP4FYGtz1LU0wWjValOVk4A0v9Fji/ihjj5EisiAZHa9s1arQ
+YxmlGs3TsWq5MgasQCd4LLaXdZ5M80+haDQf5FFlfM4qFK9swj+Knto/ps7yXJ4cJ0z9aiYTluG
U2Z1tWm4p8EwJr+VgchmwdQDFkYrZzYSpA6+YryYzo7m+Nbv6n4dH7IRJD8+jqyhaqp8ua3iZbuQ
oZsUPA+hbQ700I1ucCEsfVubktUdNM55SCd/T5mNY7dL6oJbrNg1c6RFetuH4+mLrfTNjl+xVSsj
GsvxIatdCAg3dVYQdtbm4qMiGtYIl8CPEtbDbu6AzOgGwniaX9B1OJEhf53wPyN3+oHWq+dayjeZ
TZ1ix36RI/bdj/HuR6FvrbT9u4zgTt4VmbUPk+Avywf5mz+Eb2zL82e6dqffoGtfFIG3x1rolSce
4DI0EaNWzRs9W8fxWiZT8V5/Kj3g24tsDCZBoLVyuUT7ErUtJ6U9Mm5hf7+35DpGYiFXp5pu9KMH
5EWqaIFPfgxe8QBo0ApQWppIHTbAQOpaBLwXptVoHZ8PWt9BoKu6eQTu0EIv/6x0W1M0Ai2JKkOP
cadcxc7icOBO8TH8RW42oTBQ8dst67aJreUT/XOO+7fB98GGsCQ/a1E8RZJXO/dyIrWHASgI3CkY
PiS/DvtAxbklcvFyLh+Cy7N4HRDZrH4kHJ3wFVpj2mJOnvxfv06Lbg50au9SWKGZGG6CGZq0F4X0
wX/lwh2Ocwp9Qz2iFoSc7pTHWoXOQJoJ0XRlZKPaLykuzbVjlDn/d08AfH0HYVf44IoQ07896Ag9
8baX1DXxbcYfHMptazk1sVZ8WaTFefrRmJ2JP0UYZPG+YlymJuSk3MO8jpY0/a5rLpFlhkAXiRNG
IJB5b3Z5Y1t/F8w9pwWWtyuNpRJfShO0CsVgcbT7A6Kkby0zlV0+kYrBMC5tBUjkYKFj7o6PAFfb
ZvUceVJY8CiU3gsgVXP7WFLLQd9AeS2mXRzzg6yREqBHijRS2e7lfiqxHwiQyZsXZPDj3IUOLkiM
n3D51iaJxXWg9KYNkxUETl3DhNBylJiCSKiWgX04yBoTB8Sj6uogmGzyWJfP8ymWhYCb58A4OULS
bbVojmOJw8oSel1SIWRXFqf/41qoZ/E2bmtVTxZHijDh4R/WEkJQrMARa0XwzMXpDwSrOH3jdy4r
rdXxBWaZI77y62LvPK9sZd3SwrzDdYEllZYqLKam9l7D7PPRY3xkyUKas8D1dcs7Akjid0/NaxLw
fRCFsgzXhNitpPDycRkQrgj7xwfujjhm5kegVbNFtwkk4fP15ZXNemRXdVXDmvUskNVSYh7N8axn
KpHLO+ik04P8mN48wp7so5fPqckRTUNXbyHcD0FXEAHgOaV5upgmXsMdz/Kjb1dAHYc9nqYG1uvQ
U8Wj/Gr4vSFqP50lYjd39X/H8d7nNM3Q7O2KXbHq+I7JR4xYfJ4wX5tZgG0potRJ/9K8RENaT3w2
exPrMj40XUq+Zn8/D3QEXJb/EA6733rBUANNWYR1+bYHSl9Ik9gEkbhrb2sJJCYAnPPHvL9QS3oz
M3HTDS/p/9SKavLZT+0egmjPa4emc3FCzwlCjK67bJX6mrU92+Wk8rkJr0kLqGbTULTa8c8dg1Ew
v5KvdBSy60VByBcgGjBstzvAJyLqZEFb7yp0VjMqzOcfpiuW6b9JhpmP7S39s5FDQL2Z8J2vhad9
QIrcq1JOxn8FEAL67eLpgCfwNIzgtuQUc7PGvosOI4YbnnTjXkd1pYT1FBXhdyFbnIkqCJAVaL2S
QlNBBl+S6foCI9OnyyFZIAglc7ZZuNPQWehIwNaiLgK58TcT85P+IoEHOemFSVj7jilUM/bxUMn/
p5IjZxzMk0SaEfGxsw/t5CYN6QQeinvrnOxzvfgMdFRUSl1+Ukr5C6Mb2bjhzXbM7vIBCqO6kbDB
e0KHVuQ/YJTQCrsm6Yul0NNE+KpRCBBGztT9M1A067kZIq1rufDiT2hYd9NqjvHvqIWgRHjwrBe/
8tTouPHdi5UQaFlwSmXmkaXqVWuV6EjlMGfu2mACkDIFZpgvJH7LEMhKXGiCkriafa3d43yzfC/J
4AvVDmx9yDcL1hGb4b8X7QY1NZbtG7ji1k2kOUEXFujoDnFYsb7x7u1S7mqgQLFWv0xus2XXvDg6
jCrYxw7D6XhoXQZ2CyCbnSOFpK93D/G1L78GLR+AlVLMI8BI6RkkAg5bywgjzZn41wo3Nldel0mD
SFpgkLyw4vWXbHDlnuQqOYf5q1PBNMaQNtir2yGKSzjOH6oB6Mfkl4at2vFtBqjx34EKsKaS35B6
KfBgf9cEiERbaSO1ba4DwxFpMg0uv+Xdqh3K/K0PkGg2CpkxL7LKglzJPSjKfVqkObfk3S48dGx1
hp8qOlnZW0tEY8pWGde5Z7AKwzuC46YLwGLeqcDUoJwbOl2Mh8tAP03xWsjYwlZrGVX5qA/2Ss0j
BmjsSdK92riN1P3fsIJUw7AXQFrJmvasN9Wvkxlb1LUiSOV+NtdIi2sCk6Oe/P5VhMNmHBW72adl
E/7J+2Za/3myiN80sE19ih2VK+T6fY9gr+VJVuJhqM4/XXz6SQbfHmEKk8Y2A4RfYm1OdCBGSUor
DKyRaLvhHXwFVs8Yd1sU4gqFVOzNZ2/b6lOGbtJZXnpL//XCCWiMEvzaL2c/LCGbGI6iW28KdiN3
F5EW28v2ydZ++09J+KUJYpmKSoOzZXdfE8RnnD7JKAa2T8N5vX56X5V3C6P3L8EloTnsA/VaNUrB
5P3sgrEhCA2NJuBxjm3IdKehJiRl1nJ3tmv+rMDDq1n/B0QaVBR+nlzc3e2zwveByuRwbbaGj9Hg
LJsUkX0Ix910bsyhVbkc18qXmhw0uOVhJR0datXptlv90/zX2hGcJfzSYyPRK6sEn5peG/j9LZ4W
4j+Tu5lCn5NFd5iLt6ttNjQkQo1it3HSHw6ufi1pHKqfxt4+N34BdQugaH5BSYtgzWPdAYZUhnSc
oiX8LkraNjOHTt9K0S7AxPwxE+p/XTkHh2xKQUOdTcnsgbG/HCI5Q6yfAM5fvexHqQDQLvIdC5xT
TA0ud3HfPYr0uCvwsgYhCHmo/rRC3C9t6NJ4+MunwX7jbC/XKE1jvOuZpcOr5HU2jwUS/qTPfoM8
G5EPmxgX5SQO9Mg4swkeJzWGYlyLTI6ZoI7feaUJ7USJfyFRycIiaD9EBWF9Ex/aQGsknQ5+jQwM
4n62gyPbznOYaJ7yxhMadTk/iKRkoaNySj/TKhH+UW8NvT18wss9Q3rZw+yg7314PwtgM3TdGa8a
HT7lZKbqMpiJ3MuUGgtpXnN0yWECgwQ+oNQyepVlfNMXTzsyN6CVZSUruIia6qjpbDVsn0O/rbeP
OMTeDgj7Vidg6fH1MVZIJU94S11IAsZC1b5i1nt8W9M1NViT/4jb82kXiTDdA6t1NZjo+eTRsrUD
7o1RYjuoXtZQXm2E1skiTqmNcGewv/RrI/sEN6C13xCQg0so5FhAV0oZ7RFzMCF5ymm5kqKL2rtA
qnFd22VtA0dHFdIsn78KEX29c2B3aMJCj9lPuf2Hj70dk1g4S/HO7hRdKgU3mSN5zCV/BK1k+jxb
o/nqkiZOp2bHQTl4dqD1hWBaKtjEPtBojy5wiwZRdGSOXuLb8VRrRMoLOgaO4uc4dqUn0KKBjwBZ
K8ApzcD9A4X0hYw+jJRQCe+gMYYK6lkzlOtEbnCGHAEpks2BmFSUIhXBxD9LqJufi5Z8Vh6nVfnk
JWzdYZu4qI2feQhEbqpne3Rhx1KYRsEOZVWyZdygUOIBIEnjf6aqKFLDM/O8Jk/tkVXlBIsQGRr6
VmdcQCE21oVQsyg+k/8b7NhNg+mCaA2WYEDUIyHJ6iz4gLm7s+d0QxG3sXPmyT4lCXcT7TGz2Csr
gci3ogfMavKrnj7oxqn3UHOBKlBbp9EXatqhANvteWkBOt7gv6pKMHISnZWAYjTBfroPV43ULU8p
ubmzdqvhgX/0rfC+4nZ+4/i2ltw2sKXH+UOO64xxy7HNR+A9AQ6F2FhNg4Z+2ck0ShYScgGjdO6N
XO+wV5/7imLALCoeQUb44BE0w8XrxiLYCbNFhE0FZEn3yJjFy6BVWxxcxeTKh/sVWWZXn+QzMAbF
TLpVxy/dxp6N5VTMxY518fBYNOr87gcf/tCF9xdmdl2MC/X2QFozY9q7ZGUAW6L9ftenxhkGzujV
3TauqO4XTo37BunqXL31LogwQF7Y4gXlEXfvEKUFISNHngRQjGnaEw1Q2dCcFcXSD/dZjbI7GoNd
VWTrlwgLMmcTnbP2Pw2YOhOWfwspHk5qsaU91bcJuaOLE//U5I5RoRAEj33OXnCf0iyeUifZfMoW
uP0+uEatscGi4WP4wWui9xoT950+ZuV4hdqsu/hc++9PvWG+LjBU8JOtVW5Lj8SktEEQC4KzYHre
gXEUOQ8V05cwQtDqeANR5/bOT4C/4GflM0qhBn6Ezty2VO6y3I+/KzRmp90SRXIEifHIoz7hyYXa
kZvn0LpaYscZogX3+2pgdWyMmpEox0YI1qX8nwddDriEtR/UlCuBjnZHeJRgcyyQDYrAXbSdTgMq
L60xWcX8pLd56dhqBB6qqChVgxxANoXYkKPvqpLHKJvh01fdIp0otsuKrR0SM+qMOtm9K+okqqgA
lHxlcoqme/JCPm8DPp8YsEQmayYyC0ec/TnuSXuQN/mdx1wp6eAprbYhc/Q33GbVEZrGBuvNzPa6
B1G938ZBjQFiDtafsWmsePrlhHjOma9arRRu+733rUoZvNKIkcahJYPej+HJd3vRWhdCsqEoxfGK
41CPjdn4fraxfANvcL32lXuteU5zHqL/OthuMcLpJwb+Axp2DpnD0aY+NY9vhgxO3pr2ONDIjNz3
eoX6a9eTA/HWL+7ya4rtZUUJYokX8fPlpefpjrKAbZWy814NZlYUE4opAutBVW3JArkzZp3TjYf7
AYccmxn4Ngr56z2pwKPf5PaWil7KdpH6Q8QG12zZ1pJDsvxnfLBpVU0e8EaKg6A5nbxmyYetuCRF
QX6Zn/EpoB0KyhNPTzbtKqXqS/+/fef+72vUzP1NxqGvfO1BuVcBzFoinGCebOCV4Vxlqq6/vWJn
XDof7hlHyvmZOYeFIHZWQQuJzvH5qo8oNhCP1/zHbO1hYmlgUJntR+1eC8cPeybJjYXrkfxVnEej
Cc3UN7t3bHEENH9kMG3pa+657Q15CKwLb+mR7wUsXilRJCs9FIxuZe7/VxbcLEOHOSymYZHPB6kA
NNr6Ki7nCrUDb4x40dXyXZ7i+6ztReL68/jmOzET0dhwRQVpX+riazQMM6hhJ/JwFu3q6eaCQXOG
PDuaNLw2Z6aJ5rsPCyJ6+5YScLSy7Ta2vQV0vHSjdA2BbRZLI7lWhx2Zgma4Y1a/UQzLl+wAv2aC
hcwVEZY+9ibH2XmbIg5Oeo75yzc9d1i537lLcBpkir1uC+MVxhryPXrHSyaMzF2MK4mOz3Be4mUt
nBFQhak8aEZRBc3aI/5L7jsTv8BU68+yRlgTjQ4s3ic5MxHqggWQAIIIIYkiPKVNz/GVNp5Bei/Y
7Q61/kB+dtQ/51jWungrvMmo1G6KWDcWUGsDHp/4AdMEwLUpYaALIaQ1IVb1AQhXlhWNLQ+zM+6U
kc+Y1d1PSBAuCpbAQGyOpuLN915kBKJ+s73++hQSHgF/E5keBqCZJkkojRxOpHxBCOzhDG9+KEYC
8f+fkTzZG4AsIksmnBGdWCz06BGhMBpqR3SIXmLbq4dl5ixqorHNYIbyTnFpZDrJJaJOre33srcg
0DSrDZJIn46dNGO9nPpOL/lgrj0Wf5kw8VlNCe6GHyjzNrUrCGy3AaX1MFQMg9v2lj/UfaGSs9UN
y6G2EKj2Drq2G1rWEQztTFOrqPne34klTqDbdq6+gSbRXpyUVHDaBwmfZnMIqlMPQ/c9PEIOC6KF
6iaP4e0A04uuqqiAoCNQar3acc/2mGjvA5yIbkvUawCufeYeV8FEk5M1ceDezAAK8UuQaQcjtWb5
vH8F/FpXZnANPgFhzsDtHK8TfaabvxqcTcgA8KpK6IHucWbup6IcVT9n5hi8cz0hATrWftuROT6l
T7SODm6Ae5PLlbrqm8rbdJQYN65x56q4AZFD4JvHmkuCGylY7G7bN/ThuCs+sVzSjcX0QH8DDfnI
ANd43yv61Ic+9Wh4RT3kWUFuOSERi8szyynNHBcSYOKs68sc0ZVzfEWQcuiVMHXuVbt1j39xxO1w
pxyJy85yiDGSS2d4oK2pnrB8kbSDyjSFlPb6PbbVPP0n9NdRLjbuPQGzO8mGf998J5UbG3MkfLJh
PvWhaIJTkcpqXAAX/WZsSwiIBVjvlhcK0DLdqJeYRIaDLkyTVePmkNpboIVeDq1AWgX/Pk7RO5NH
tycN19ZOU5bAUSa+8TrHmtkcueGEBkdrrZQRlCjZAiTINsCGPG9sWAhM4b5WlpXiOVu8Q/OoK5Uo
EIwSHXLB7qsYngF216p0GCKqM+BB/c16QgbKkIqo5d5PNsD6QKtrpnCGTDjALSb32rGx2XgtA4lN
8OZ8jLLdYlln/uvCOO8rDixCVs0MDGKOMGDeEQvlgXp/6jrB7gqsFuHNBIx4Oktu0FraNVLyK4Y8
Szp6PL3LG0MRe/QgBprVsd7OHtx+cCIkBM5DG90QDkJQAXFPy59z+BdN1yqFWAzDPrzwgBpPvaci
7/wJ7hUti6XT1rfqiFdY70p7h+i5AQSbGyDgOfPFvwMULY1X45ryCxieE3U0oRLruqwe+tKJFJG0
NrXjrnQnkQJA2ZXKsutxSTw5MmZh3ErQH3eoSaU4IApSiqsIGSnxho7VsMHonTYzO75dnvh6ONtA
9ge2BuM1KATvGcxPECzMQJst/79PqhMi62PO7LQmO1IS9I/TG/R9OuiC3vofsEKBbqrjjbaSG1y+
FB0ryqqbYeMh1kdt9Ql5HQWUaHxGmmKBSTSHda3+sXCIIfptqltxb6+BqeaWv8/c4EPO1km2EjJc
/lIUosVlrCYu9sqFE6qxt6t+wtsQSb3ITa2yLGQULO207niHinV5yqFbg4miyzXgYNZyiEX1LpL8
BGRXy3suHsAnc0rwjpALeGorDhB0Zp6ocl8bcPbJD+LT5wrug+5Gl6Q5P7HPWROpTf8Q7VbC+19q
pkACwC9xRc2Ot/Bc8idNNnDs2ZPwgvn6Zbq714Hqv+YDF6T1v+cUt3BzWJUXWTkNBQUcSqNGr7RF
+5aE4L8RlB8CsOCH6xDMK/jTkzA0nKyTY6lqqNMcHJkNRi9Ibf2RXaEcMIb2z+RHAP4zODqo1v8Q
o3NgSc5fQp2kDeWROCI2KGrcdjG3UGyr+SwE7ETNE78qSRn7JLsInFSjIwQi7bsmDbRYG8IUYm4O
CvmOVC3g/C7p4RAKsd48BWm5UbdPp3hyZoTY4+s/Tvf4CA24b805Q+6Mvc1sKHsINP67JseGQVCj
RTxKcg8ArwaD//LZFzrj2vsqyW9HEc5L3DGuE1KYuk/tRR29hPWuZju9XdJd58ESQ4ckYCcL6EWx
xIWVm+lLqWvHMgu0FKwxSjZnp6S4w9DglseCkxKrbLpWFfGB8KgdJj3z/GLvXYHPR8TcihaP9wAG
6K+3uuK1k+5tO9WqRpUumbl7CVZGh7/69CaYLfKGs4g458QIA//ccaPfxp19vJfyCHuSyTo6TPgs
gxmqziwMrVUtVbhKaSyXVSN7blbTIRBjVXQJaurIDJehmZ2ngVxUlvQ4nv5LFyZNun9G6pPvxE62
+q57IT17imGPoBZsdtN8uLtkX+3nbI4FWp5UpUQdKHf2yjAPOig/fBIieX8SMWFFimwd9ys89xkr
eEEGTkLcp4z4M2YQQKI9M1BTl84EnF8mB2tidKqhPwt0N5YaRGzoIV6PkQt2YzLz10Z/NHgKFXCQ
F9Q2dFT5vvEJ0fI8LbaMmgqCEdTltFuXYVbd+Klk+n/slxGLISkWXD2jrU9JeL35iNknIwTg7Fek
ifxewWUP0ydt4nugZ3w89h8o+rRO6BOdVX8a7SsSMiXgxNgXeRRbkSLSVBwPHTxMtNbDg8i+Xq4t
JGUNqL1cp6sJFMu959xXF7kUAXbXg5r6dgFGNQHRaeAIHYRcboUxiCAgaR3T6tKDZcfPJupYv1sF
RdMCrIrK5IFcb0JzlJEMNeiLg2rP+1nWWMbASnfb7lPo0GwiQYCBQOCW9tWLcTkcRQReWG1lxrKW
qozS5LvZ1CxzWmHM6uTqEm+NMK5zR2WAd7BPjOv2JpD90HjCsGA0e2xw5QWEubVKiQJM+6IMWG6K
06GhL6dFhQFovr5lwRA42fjAGIomtcoDzOkinFxJIE/7pVHEK4ZgazKPav9Rdsun/xt7qeMyIUJC
LJeWoXS23yMwVez9gMmIFDe8oS80rnptwuL8Dr2UGQJ2nvOHOkbEFYTX2xSVfdr0RlsXvT66arQY
1tsmwJ24TbPJ0PYivJkidSB8YSX1s2sU92jINkyxUMDt7OzUHtDsfRKJGzcSdYhWsMXOvjoBOCnd
LnOrBphM+/JIdF4HJlHZHIeXdvexGyuToJcDVSkPph46PJExayMzjbGD49Vx6Ipqr+Ne1tJxxA1B
81YdcXIoRDV2/1VWmXZsEGz0fg9zxpVe31rV+mC43ggqIgKIAZHiCeZ7Lzgz0IG8P6n84s/zjfuq
438d0/rNLYNDp3VHUFSMVtF2tAhF4VMUTzeXpRTRV/ep0dQvZOUdCe4HoVBta1rBKkjl92tf4Xfc
xhbJA2vd92G1ZCXQZK7EUODmTg+upAbSY8SQFEAmw3Pw6GB0ZiF3+tNeWn0nEHGT0xgOrdijIPBx
SCGmzOXcxBHhKwRWtBV9mdjYFycJGU0yZDxuzZWJHAJfTAJkNu0d4eGvJqV1TDEbK5OhiB7bghuj
qu/tULpos16Orkk/8oziL+qrKR82nRQezoYQjBYncjKdO9Y5ve0VtU22NQPl0zs+v2hZfYoopG1R
FvKh8cPq6ULV3mP/SHAQIub0/UqyA6wZZ2IWoZNTJ+ZVAlaFKdf7KXvnLfDjsTnxFOAKA8hsTlbe
SthXvcXuT8jqaxgGcqahoKNJsc5IuxTj1zUGOPdLb4nFSScFYnGbNdebvJKDeY2vPq8y/LBTIRE0
qNKniA4MFi0SIAl8Z28aOFVI1FV/Cz0Ek2MFnsW+ff92wYZTywVxB/qe5l+TQjB5nt2HRWbUrkL+
ZxCnJOTDKEUmfDwCzKgmkkDfpCyGNtnrk5SNPdDOLWspzWiGpQRfQQ1g4Q4x3D/I9eUeMo3wF4AZ
MwtO/dY+X/rKNBy3p3FKvb0WGJijL1XNT2qaEDuKrKScneGWhIosUVekUPl/XqbxhwGbK6hrxLHV
oRGgw2HiA58CNpObx02KtwmEz4F8FoHl3E04vW6nyd2WQfl2ZOTtCaAysEiYZiKyGNNjY5Uhb2wa
XSt5Esb387QqtkrDWhRKDiAqmbFI3McwLiLWZIleLCxzAZk7KvUm8zzStfpiWPXLgckOypPJJPse
a2b5xg+ZzJ5JBfRp66G9DVmMTH5o0LolzS/o2KZ7aAzVoYT9Vo3cNNYIDW1ekMtsgQHdbO6xts76
i5Fpkw8viFMdx2JJ+1Z0Q2WZzXp526Z1kvX4/Q4TNlMiUbsrSi3UUSHfApkb8Jij6QNFwyQWrhJ3
zldj2edPVxV2KbGQobRARfgI7dk/mcFIXAI3goEncPiKNlPT4rNK7LUu1+NjHMk+oP7JUdpB9G/o
TIk22YezkJirj+8SzcbWBtLiLJFRGM0E462SOCA5GBF0No6rtyfFnhLVPQq50FhfWTGCGP3Ml201
b8PzcPtIGv3ET6EtHqtFt2ZZz/1QtowHvzy2mH7uB96JfyBJevjlD0SOvKIdEgYQkm3i3gpttnsU
wG7z8k1fY5oQRBKUNk2K0O5x3jFVuasMz0VkdppDFgrpTUPXeD6rP1ePVCUwtVjNoK1D2AZHIl1N
KObA1fEteGDW47pzkMaF4Hlu8jkx6lqMDCWdXGbeswErWgaQ4bqZaYNQqYU4M5LKxtcr1bR9zlsF
17q1a2yWOaWJlz60xXfesRLwWfPlQR1QEl1RWSxApiRazXWIRzPdRzH9PGP7WJ89wAJnZjLUiOv5
fRgx9+vJx/m5SmmbtYOJ4T7TlTrQyGX34HFo2sEn+0TnF6/iuCX6NypS4CA4sU7GvHGu6PkykPOi
bU8qeQd8/8/hroFTrkQasCdUYWyft/b3zfPx4FnkUHtLl3sZTrmbpyArxcio3jELLZYcElBMqG4V
cvmNl+940Ps+yZ/7ZEjHLhZkaqpHJjrPwvqUzoLExYISitIIKfadDbNITode3sPSSQxlWnnZ6j0M
AAb6O8GzuXPQ7BuoJ2ja2T9RYc6N7CNUt06+rtt6WtnaVwzqCuaBb2avbev0N/vEhvIjYfsdM9NS
o8naJHtZpf3BbDlU6YSNdD+HM8Ow9Lk1nZ7VUg3A4a0xzzPJty/K0RCXMQgPalCUfzFU0rg9sBgp
KZGMBISdqZLOn2Nn0FF3F7zjh7y2vw2VRM9TVBD1PKh9bR00lk/5lVCZJeTOvAiKoepm4gRgtGxR
CU3LK30ipo4mAaF6wpL+MiTJC7+qeg6a9Hm/O130Agy/iMYd03c/wFjiD1OsCLQ3QhyqHNulvGOK
+YPAKum3d1Av5eEALSLCpTqKs6O1Ld4m8WL5TYcriiyqvd6DCk9XrhRhbVT5sHgkB1MURA9I9em6
0XIS7wLwfhR1N0xRsl+QSyxHZLnt7OieqRf2ChD/RBOQBnKoxSLnsQkofU/RSrWPvy0zcGU//w//
XSK9SRiJ5VmsBC9tzGrHPCll0MBNiivyudFLw4JRZeF1nlmONtzJuEUUAmS6lz/5/N/60cQ3sjiW
FKM78b6hWQC81QadrK86b/hkHt+zzMSTXTHXQCvmaHaCXPGbhT4a4yeYpipf38KEClONa33zPMXI
q8CrR9f6tlO64FVmzTHuaJles9mYb5BetcieN7GRkWRSeI335nyiXIum/G21B3LoRqvter2onwcT
1RzTqPnuib7hBzJacvI05suLajVEHEdKaEHC59iYYeWdFE8EfmDxV9kbc5BO5G8Ttig/8SlTCCUB
D1+xOMGuHgr89WhD/HamXCQfaGxw922V5+cFjsPHJYIjkWKbL8EfxzDsA2WdLPcfzObteGEIP/vI
bZIjXQgqCm9a6E5pgIJfys/CumGh6h3HvtFeJ8Y7xx5rP8dkqUN2WbQVnJ0V2KNXoI1IXDwEQcQH
ASvFVN5yTEmhLv4tXl422DPiL41S0ugO0SKhwRJweBNRvYljEhmbrGgpmlBWFcyQTbQzWjCfLkKI
YIwTafR+N2gNIXNMSgIR6uGsotXPvi/I9m5q/YBzS93gpNCr1V1I2OF8x7t0fenDXQEUR3+4/UpB
lF9rzANkYXrLptqy4Lh6jgTQxxcbWt87EjmvfFFTyH4LRZ1WXzACBgmHWf4VFd3wODiTBTg57+gg
2Cj8fUdvwTVC/s+pqlnpipWtJov1NBkpeDmDTaRxbA2PrEMDswACdbagMP1B+BH/7HF29Tw70tfI
PQ+MGnO3hssJmYiLaKczxZNL1DY1anY/t+l59dwS16rasWc2mo752zAama75k3F3srXuT2wB7yIP
mI3LZ6pAi8zQsiEZKNhM7bkarSSNZ72wyKy/h0H3XUFC8ZnfUoKhQrmBI2eXsrVAC/aF5XWpekkW
zvxXyMutQ9N4a6fsv0fgzT3uK4MNfgUEUO8wylXbsUhwQFKGl37TjRve/D1djxuoNUFrmT0qlR5u
ih2HwWVgQL0BQLabmAsj/eE+2uFQNXQm1yiAuNpiz9YqJq/8W9uIOgtg/nzvFSvUQP+W4TxROOAv
iDDkK0RNxk3tonIerhrjGJv9yy58dSUzvLsmavNs+57sf3+I56quZjttI33zIvSSzLLc4BbOle5f
togKE7uM/h94BEaBimf2T3EfZ7gjtEzetUE3yJmI9AVXqIguTDspwTCq9WJExy374ADRHQNwqIAq
ZE0HaGzHyAcDM13HrrjhID4KzwYSgLcEp0QwM78Fy/6uh7tQe8SI1rQMkzT9W9kjrBky+ktN8MFV
Dwlo8C5svZOilcaZULSVi/WqPQf+mqbnlgMWqoqGA8Y+echeUWmvL88PW/xwkkBJVjoMoVm5HIiu
E+Yc/PUcsybbR48gTA9Rey5tmtzhH63yMoy6boRNvDFh291r8F72PNCKtBSJmzuVIILpLOCOoFPO
75Jrb22xVZFmJmdVXtq03I5qKKIwU0CHtTLW4CwoF29Gda4PBgexIYjKUqMmdjbdUcoRdTFhXoJg
JvDkF/A7JnyW7uYWqb8UM+zjAxmEbyDXBRcbhdtK8ejTbC+UUUQSdPmuaGaIqtezI75qrRGd2c7T
RBSSf3r1WL6/9IlKngJ4ZIxrV/qF+XP7hRybNyvHUbiLEth5ZHWLA5sp5Vm7zHB2jTAiaOF27d+T
Irf7qqZ/nJ55704/JxByq+JcA4YjQ+0mALffpwsR4M74kx/Zf7XXfvNhFSNRp3sO7evB677cz+QF
98D+j4PV/0AncCsOGBHk7Bob+Z2jsGEO24kfnLFEXpZ5raCre3yyc5//RdeLxCvLewjLMJMevQk3
Bqbgixx5V9L2t23VgozggnKIlCUL5mPqI2P+YWmdiwO+hvxvd7DieyaiMou3PElp/T18FKQABWce
Xd9Ao7Z0ssUz0Wp+YZaMEznaiZMMYSKgGNQfruBFo8spnV+Gnocv9lDVsuD4Q6NqzHW/t4GpqM1Z
Wt15FPlJJpf/RS+MyZ8f14HZhpsYzlzrUa0ddzfjoxtxiqG19syBr8o0CdawuGP1iVGyG9WyP1mO
hjEGtTSk9pSrHsJamfOJXrR7dixYBHmqOQuWsUOeM+n/XsyaeUFm/+hIWd17cUq71Lw+UHi/QP8X
0zVrvCUPd6vOP9TJhvcXT5n3hhDHYembpgrsQ2kb68OUed1HeVPgvza+QJNSSNkWkplwvxR/y9K4
xGD7OvHO6Q2vVQL7oZiqilGOmylFHSCIUrPUk2hKQeiPbx+fW333PcDqjEylx5/yjmhdBlwgml4o
w8OjN9J7Nv5feMhtBkZTSaO4Epd2L2Co0qjGqJLsUgzSL8VOlYaL8BBmKdEr0eCfcyr1vDTwVQPz
rN/CL97edl615kBXKFx240ligv/FbJVVt+6tAMvNNnEXdb0PxsTT3TGFZ9vo1WJ1QAlEBUsfJu0T
HqbsV+q7MGDadkIv6iNKz0wr2LqSsGmjdbKb61rQC+qe5o8gxLYK/gglaHTI0uxGD4J1xAaVX0Fl
xNd9pRp2ctj9fqDUKgF939upqC9Bm1LCP/rxvia+99qcPaXg3N4AhgerAfg0fdIyIqKkFkfLzcbF
jGyF9ItPBAJ0Vf/54In9EglRuXOtanPsVlkedtUqyuXcHRV1CGOxyTrEgeXcWesnwseaOamJZ4uX
WE9+SC/eAQGlkgRjJQvcY2lxCBorF2JtlNyeoQSBm9qgecI+IWqxXDUST6kitF+7Ply+BdcSKHSR
LMEXQUXjvc+ukrtaao4KqZJsmDH6jlnqUwWMyGG4rdU/2HdrGSFBJJP8F76PxY//vvk10B79jo72
iW6HQjiUgrMvgGDbBv3VUOtajmI5m4BUreibeMm7COO6ZNNmmAzujmcH2wcGE88taM++9zf6ToXG
/aXbKn3Q4dopNk35okEm5yWxW3C6WDPdDpezr69z8v2MJt7SbVlvQsyrZXlVzZkRgpmJ8Nj60OuY
e7LlWJ5ajoM6d8MfO7YvBvezyhaNyvn2OuAXI0SznhRVMuFDNAl7qKaOinlirWZeO3eN1L27mo0X
RPE6ceMxrA4B3LQWUmgeHUpZf6WfyEd+/+CmEpIvaOPN/vsRbpdMCjQhB1Kzp0i//92OGCUil5Fv
RrgflUNPjvy/TkakmC7RtpWOdD8GxBU+UeWEDb4eRraA1ukOMH0i96nZSC/ECEGwur4Kq92bfPVM
3HghaL3mxRhKj7yvINb20Lfn5dQ8bJS5PxY/j0bs386uzy8M2J4CpLrJ0ZDdcWGAUL8JrLUbrUBK
lpkloxSxSc5e0Ax179Zdb5fHwmgCgP4K7iWmYFjofqfqN90A6ZLEibEnywuwcwZ02Vvzs+MIt1Th
YZEtyLt8UKmuR5qoM9mBtvxZB0RZXiapEC3yA9GDp7Jj4FkOZWerGHh3BnhwcvyGIatkpY7nFtRa
GCBiB351ay1PqIN6EZAOOrewK58U3E9ippeEscMFrAfgaUbbkTOSBr4HJXO4z9lVnG7VKIHKBqJy
l8rFYS4lB03cGvOjbgjbhcbNLkE00EkWn41XuSjKJjmHQ2cOZLS92Lx9ZTf1c5sBMvarXxasJa9E
cULN08qlRFyq39AY3MrF4mOnzwVEyl9pwPeTUAg1d4b8uMERWNLKpXPDZ3hi4AcEsiWfkz1CYo6q
cWikD0NToxZ5LTuPB4fA9av/4173KSAth+1EFsfyErvwToQ0LPcHpVV3elG8ziXl9Q2qhiiza87+
ZSyJeRwI/ra4sjrcXlmwcc7G7SnKVOzkqpQAVGQxUOA30qTmknpuffDcGoPp9yxp5gM5revGckzK
LQS+jAdUSMNChhW2UXUKIPfxbc6HwGhTgwZHquAbxB0uP0DQ1VHyPKszyYMFms3qA0q+IQ7Pf8Q4
BIF/JoNP8GRHjCz5By2VdWCnpk1Kq0v5o0lGX08vBJ+xbSbn83ndWMUWZh2inNNmU6WokYLu+GqQ
0GbsAmSeoVCMhwJKukLYHXqU5Lh7+UuI1KPde2XAYyjCIOsN4S2ex+A4LUa4xKq+cPs3TTzrq7Ct
uBTSWNu+GVYVEH0tMipPUBLcuKREWRoxXZzUwMD6LKOJ3YmVyS/7PuOykjNePvOrZ5nJhvFpGlHG
LjlJIp/NcwpCdo+OObQ29cBKCsD1gEs5MfAWkjIoNatJYzhlK5r/c15ywfY5YQihLG17CBpc1Lvd
gLUNl+k/kwh9T2iGlpX9tF0A5AoBMAzNVhohMzzzO4yH2ZSi+TwNiXwQ8BGPv17KqDco94LSYZH/
wDaxCA76e/I8gQrw9leGKKdBbU1QP+kvIGnSYd4sSJjOD5PUXj+/QVOpSlthS5+3DDAxGbJlb8nt
x+GPfs4a90XfFP98Suju+nnmFc2m2pi+2BDtRnWhJgO5pOC8i+ltxC7YkeAQHdXCUifQzmI2jOcN
kEyu40YqoOBl8OP3lYf4pZWFuhKgvfj6YHZFQqyNU6//zWTakZcMjGDiFd/I4RtOMVI33FNIZf6B
AlQYTukSXoLUu3VSkveCxan9yz38TJp+ImdN4Uw0eKjhfymmhwIqXbADleflrBpqkB2YvVVlYJmZ
bZoofDU4cuACWw/lVJcGVnXQQ6PsG45a/PXPS7lL/OahjrQtE5DVb+aFODjnRrljOlKUY4mCfBfp
Sk5BFfy7x1xZ40ECG4Pc/JShaJOJiJ6iqSxKMP9DOIeWX3aS4OZMGfnAWJF3RAz8tluWoKOuN+nQ
rpV34PDqUeceGFQZ9dVsplhxhLeWrt5n0YG+vcysJAC/H/zwU8cH5scDQtJgse96bUGnzePjQeQc
RfeK7qD08cfFcPd8rO+RtiYaAv4CmzXZ6Kebqz1NZk58JrmeSPMt6CJbpQ8JfO98VxtyqXra/jRC
DQSGTN0Ex+sH2qXyenQEwIRznYrr9Z9aGJEIEe5uvAH3ufzZP2/OPJChzzjUoApf1ZwF8ZprLccV
WE5Hjkl7OM50CUVAyloHryiQSb2sP3GwhnoXxETAlrU9DtBiHHmjRaiogsRTTq6RV626gUZZzaxM
kZru2iI1bxqb1QiBElyiOs7ei9TwQ/6GK8+ZeUnZkHfgNNc8eRNoFz1MV1SpD1lwER+VLkrW5amR
hxI0YOi9AJc7NmSzw7H4UYuRBrLBSP4dQ52Nf+sfKTgYUJgPaJApD/dLLYYV7XBuuQdenX+yxGXD
Xs61SvIXUU0CKP09Y0YR9f+2/7EwWzfe8qyYdcl/hax2lc2ZwBdGfTIFEz1b1937369PD38RA6Li
pZ8VuXnq+M4iHVUrf4BxaK/vXq13LxUCOZ4X1FXmqM6A563OLuVS0Q8ynwrkwi4UppDbqunAByU0
L0hKgb94d5BU3NwPJb8MV6bTY1fDQmNT6EUHFWcH8Toc77liHBhdKXVPlsctceK4h1D1e8p98LvL
wyUgNHq960PLjuMGBGjW2TGRIvcL2Hq0DQHbTIg8+BA0XGn/gdGp7OOySXBmOPA2iHVkMgFQsbXS
KY3jWnwXTb5/MWVExspP9bAtU/MoUJ2Ns5scH9NwFP5EnIyfbXmRVhh3u7Cnk2bclgc0uw/uuFWc
38+ddUDlJZHtBVO7EhFY6eHPfzO3SeHtRbm8ACFliWGQ8aLt84TuDNBhCwV9iSOTNewv4ukLu0Zl
aMyp6WbntOPHJYdKuLJ3muMh//vWda5I1+Ufiumj22KP9amqq3FWTNjQ79tz8OFqYT/No/4cWu54
BDhIQ0z7OFjj9LWNOPWWQe5mYEZk2dWt0mkYMa8VV5sD6z/Gv+cfYUPaaftrbx7Km2DmVadfTFjc
T+++2H36szIpGlUqE5UMYFNCe9ULt+jPNDl17v2vpJrvkUSbWKRldjGPWXwibd+/BPdBME1Ur3tR
Zqkn6UtXmetwXHVIHbd9IoiiJbr13eS5MjCE7lrpJ0yMkLrGSRfbTimTz86sT9v4KUEppM8Kvdjm
AvYfJnoUnQ5dbaddirZ7CkPYkpvdH7fSPjQxxagSEbobA++nYh30tXCqRkAwEmlhGaKh77Ny+EO3
bgcpRSaBd4t6Gbtp9bVkDsivcrVQH0//yU7JepAA8rrYgBuLak2BzYniofYe4U9sSAHS6P/5VbCc
bsb6PbItAWuRdNQvIHbYE27pscLtqJoTtp9SXRGoIt5wbNrT5vUTWQ9ZirNH6O3pkM0a2W3pI9Ng
kzGeoK04hu9ZHStNp/C1ufo+r5qAjaWkgVr/CFbw28bGTcYyIorrj+d/D+VYQ6ifu/cHX/eqgEAd
7ec4GGesQLczehNJnZuKGXzYihuLFQujkj/fsbdYZe3iDESJiEg1irhJiZfIeqrNpbJEBwDLJYWd
qybf+v2iGTHTVjieCSdLHuBtZZrP2p7x6iDew7jPfxxlDtTZority+Pp+4hlffni8OPtl+aZ7Hqt
I+87clT4Dprnn6W6jUgOlpDS8RzYD3EldzYOnJRsAVwAX9IpMw0iyv6XDmXU7ARgZyQUBwmdJqFt
W/PRYj9wC1e/xKPuU5lHtAdKU3WVbOdCA14e+Ct0NvsfqNCCzM02SVWAH6+oKZjMzYJLEfc4vuwQ
eDyehYJ5VeEDnT+RVHpDtkdAezkeKt//FAFSQMLVM4rLYfxJRs392Jzz3Yt5O2w0am0q6gI2oDsM
roTTkjIuM41vedOhhahQhZKZOwUq63drOXsyJm82RzA1vapE6wixAirnt/jJhneM1TiyDqkmBXLK
Ia3VQ1Y7BybSN/C3yf1m32qMHUJelxKFwGBqhqobkbzPLJEy1NrNFoskYcdcFRSwg7sYXbGif9k6
fGed6wU6KdqtPvU7Rhx9xEtO8keesW47qcQh+zO7tTO/wpvoRwLEscL3/JZfcRuBql+kI/Kk+OSv
rDkgi3WL9wqzwkCRVg2hCYTB+6mfzgHjKy6yaCOZg4g2eYzLfdM30zNFUpxTzisXl9WBMmBs5KiE
p1nsxhi3C/7+WYaQwqv3ja7U01FyEbrPOCuAn24wXk4LJ3tkuX2TQ2mYex0u2QlZhEiOVbilUCuA
tXdSDXbvwsTI34fe95khl6zzHFQ/zZxIIVU/aPz+Q9+Hzmmj2jcL7P1rYnGn08KAYz4gMJxxZyvT
NY65VwDyd33klYkHfE4mmcRQikKg0EMdYOLQWh8MhooTeleFmKoxy1GX6x9VdisCzoXbX26q+Cyl
HLbRjeeJoIOLcYUNHbVqbsYzEnZnrQ0fiiYK8Gxz6TRv3Hg90n/VWx+C0noKAVNRZSOUyUBhyrFg
CBmdBKi9kWYd+0iObfy24Zi0aj5ovfbZZEhGdCdEDQd/jt1VFN8+qBvp/vN699O8+eslrLWATHfT
H3eDhy+e7dSCYKTAaF/fl5kw+DeBc0+EVhuDAflxYJZCTnoEIFzMvIVt8ySRrPH1ICRn/YgDxmai
NmmrQfNVhfbOGfprm2cVrq8gn99as986JzuYA8khUERsqlAu1+n6zTgtTOSOmeNdD2egOidcipAm
O/0t8MnJkwGSWH5mc1pIlv/1wwrvAJKdf8ctNBO55Q1+cBJONlV6WoHtVDAC9gkqrjX+FAimuIdK
ZsgenwJamFpZEv+skOT2D35D5BGpLFL/tYu1D8t9ZZEszFAPqQKG4gS9RgKLbVP+tgP1v6dIFWQv
3t9qId9eyIYXWXWSSWd6LZH22bKzZJMXIJWwi8sRyRPl1p6yysWE7A7XWOwEolKYZv35skHiaVDC
EDmzlGZc2ByOnPLojt+CFinPEzpMFXxao2VnvE69KnJidwHTRjKbqq7eDdgJP8dJ5wIOtPtqQjmL
FdEHWIwGMon952+14VZA+k9fTNdmWGbAQODtyVRRL0guTuH1ulce0oybIo8eyPFUqczPgJEgee1Y
fxg/fK08AwdQ1S31CKiZd4Sgf9PoZyjqb5w/jSin4/e6K9SiY9icPYMFWw7TF0t7rnbwX/D+W+NR
tyMOvzltY64yMsP/ICN0XuMDdeHzsBQI25/0CkLZ294wAqnyZXRX9p5suoukQJ+PGGGPDwuB2HXM
kwbwOzWl26JCBxa/G0RDDBMWf1ds375hQK2es9WTmcP5TZD6UPg7Mv83ac+HdgoVlZFY9T0at3CP
fJyuRPfJCrHKc/MZ+s5ZB5nbWT0C3GgMkPVlC4MCMY0LZ/blgV9Ge++fDt/71IytCGVxJdlRCZD4
/uF5FHZQwiuWhvjkQ3SNXdfaYsUrJ21aRUGn6gnCc60eJ/EZv3+5nwkMZCeEYl3mo0yByOjyJt5k
FwFkZuQWu0uy7xswCPF4WT7k3HuH6vLfVtcynEUihjXBPJwy9kFDyB/VWmcHH2qNzmDB1wZwyhH2
yBNJFCMxRU+TtemHRMl8ixMuXHJurG6ygenz8lrSCiHF2kqoMnL4hIA0buDyl1YGRwyx/O25pGHD
XtaFk593q3Ft7VJ4pEHN9uceua3gwMNE/NIjPyrDboq3rwgiVD2/IlErgoq+SxxYEBXhEJcumB1U
joyIs8AWZkW+PrK50lq9tTBOF1eFA8d3oZi5dHivPufWIqF8/Pbf1B2UEQCsXPJXfE31BUkrBwjS
CXbpxpJxRt9VWaec8qz5VIBxd+K5oDRHht+HMsR/5e1LXET0QjjiEbdze7v5F6JZ6AKiWxNEPWuq
9TEM8RJMNOMqVPJOAOR+GqZ+zvoIqCeZ7QymD1M2ZZM6Bv4Pgf9nuVETZGu7FIUOW5qLmF0mNc8S
1RLCrMvYaMT+tnRc67ZdSYoqHScbRy3NlvoQdH23PuQW2A6fwqIwfe44YD4NSfKdpBHAuosNa1Vo
SlNCJn63zfvpS9pTF5ddi7nRrYxjwWD7rMG+63HaIE/lRmp4U2QOeQilXU1bqpSjQXnzHayTZMo9
QVgI/DcJSNjIHvQPd4aV/VCgkL7oF8mQlqnbeQMe6jf97AXAUGOJG6NmVrkhGzm5eY+TYsjGwPrs
7eVKT22hHFGcXLFrMlgauV5BNPeMA+U8h5/8TplJVFs0fSYa2exv6R3Hb19TOnMGMeQUe+hQ5vBM
fj3p+CQTyUpl/Y+FOc3tUZhexGiqPrUG168EvlJG9fMTp52G4lRxF9Bpn9cah56camaMT3rgcvy3
Tat/J89i+/MZQHsf3HCo37gJ3oBrHZxIYsMAJIgLVUVwZ3XsvJlfxXcioxjfzTIG7BjyteLzFgRt
BaAxEoS7fIYzxkj4EeNyP29EnczbqPpZ2RbF+Yx5rjNJkY8b5AEKleJL4J42Qb242SMSrOxU3muy
8vfWkxiPRoFPxN2cjIBJXPjUInZK0q2sYbBwPpm7H7VDHq+/+NnG6nSlwoWTyxnHJYe7zsOIFV61
0gPVct4XVgVhCnKXn9G1q6mhnwL10eg0BwuJekXVkkVbsIPS3NAKZaQGcUjLbU8IxuJ+g+7w4StQ
zo4TaNZksGeT9CXmAQK+maR6NsmUpAvEft/+ZApfEnMj7DKFrty7czC8LfCMrL8hLN43fX5Lof4h
WuHl9gj/Eil3K0pxxgJ7okYlflS1vpASI2/d/1lpyN+fhSD1h9orn7SYhqSnpn++vtxzxQ1B+gg1
FPNB38xL8wfZWIOYY32H1RrbAWWk+1Yvf07VVTSRM/xSuQRylU2yDqDRcLvjMJLANsyiftt54XtO
B1gbT0sdVnSD9elWWhVm7J3kbdYwNl7NOz25H0Gc8K0eO2lFBhIeTYfmkkL3MeVfABUyu7q6vLEv
YYOnYreaijU6jEeiZssfb7QTlg/2Mw0idOK140tdF7nU/enXwCjzEg+XdqAl3i62xdHrkTh48LgQ
Kll/aFzKFNdUV2FmbgaDZ8uGsHqfCVORUaS8M25DrMnTx/iehGywscyQOIiQwc2pTD9niMSsrfLB
ULLSS3iGXr/tIEohIAA+U7LZPKOcEyzECTXdLfZ/JyF0YFwmJYV0Ayufd7eBqC9OdOwWgno1Hj9O
PMQLskL3J1iTvi4oP3mq8r6h65sh4x5nghOZoiZTMN7m3TveTaPw+K0c4UlJGeiYW/V2fp8RAM51
8/tgcyVtZLg44F1Up1iU9PVMBAMGwk3qHgXrYxBeTq0HccasPGL5SrWHVIa2TQkBOkOWg1DsZeMR
hPNUdgLPRp25VRdMeSAjWK7mZv7nQ0gzNuH3Qu2ivbBW9u+rKXkl4FlHX+whH3qYAVcVeqpoNBOA
vZc9B90WQdv6F40g9sNDbfaxOtKHuUgxM1ta9+53dUsOOpeKeMliExcvyNrdK8xtKiNd/nRe7tsZ
oBBaba185dV0gBu+n2Fu33fZvHc43rE5C+uehMdXf5lni1ujA4jJiYHzto5Rj74alZeW4es6t4HS
jAaAsooUqF/IGdUPZEkpUOx7mzKcOwk+J3f4DByV8BpNGlsaHvPqfYZu0+v4jRhtpO9KA5MtS5xe
/UPznhpinQ8peyTjc4Vb4PdFib1Z3Tn2pX1OLTJvTmG9VNDPh9Ie7+rWX0osfpOl9JRVeCzNnAc0
mdshyX3YaX9+rLGc+q3G63dV1zCwjSw8xDWA1ZIkgqgHDgpFPgxrnUvMw8gJv8Yc0PrLL1ZLXQw1
k6Q/6wYRFwCLskL1hzneqxf4GmZzI59u7ZyaxZwgyttT+1xromrJCPLJg7n9pSWaGEJyQtglTGoG
blAmZf7bm7SM0IJ9h4FGrpFoHDYWQtEra06zT1cOBStGfoAwG1LPfTLe/GUXEcy8Pvp759d2lVog
IkNLSMGV7vIf2gSjHmZsJP807hB7hK30cWgLKDQlV5cmaDmNYbbS6M20yH/sbsVG/bj44HHgeA90
P9D42hGikT1IRleT2fqKi9Q94JS+Kyu68x6q0ghERVQZNUJVFuRO0lQ1B9c3kDW92vgeish+6bue
Trteiqh1Tfc3nFCBq417fb/GmsWMNrOxfQ4HJ/3SfRXaW1EUM/I3U8dmTaiwSpsqgGTvPMd8xMW6
d6+CSMuy9GPKqKbB0rOxhwVuZdX/N3y2crmhSq84XrJe6sj+KPUQO8LiWaf0+8bY2vNZb34n6vFo
J/fC5M3ZKiQwgDbkpOJJSyWmuO+ZsAawXA89jcCtHt154KBVGLUBJpPA46l7LnrqQWji0BtbgzZ0
3keYoGSJptOvp2U8x4BujyLl9wHF6vwviSrLkk5rsOFXJfR9d6R0Uk56IKaZmxYg1ASDg70TiBN/
iagvE4z9txjmZ+tS9eK4MxdVQcVcs06ghoGiw8O8zCUHE3JEFJ1vy4zpEEaO3/zhcp0U6aDiWL1+
DRsEPebVPsDU+enKEGMeb3ylJrBcA8E+qk2gUuTolqo0oHb3lrfz2DDIDMj0frREsnZ8x6R7jEr+
7pANY0/+qRXKAEI+lmEzSXipzDL45A549QvyMLxb6RGd5y2c7yXqrH6saHKs3FkoAqAxWVjdc+xJ
mituTcnjU8+StUZt3RMctvypxHCAU3ZhFZoVhojs6dp2pb5XbAgaMhgXfGTgoPlTB5S1Hbj0/N6C
JiRnhQfgRftbZKfvyi17EIGrRe3UEZWSENAqORiw42UPaW7t6mn56Hd+ZEiZ5uadTGyWG6YZokFm
XcP4rwK8yChlS7HPmIDvW52ZT2ACXWx85LZRrGJUmJRph45UWxL+fDPpXv8x0cS5q26hn326+0vu
GngKP5brHPpWxE9uKAZ3aYi6Pvq/Kz42ClSm0KLpqHG403RAXfCPZW6sbx1w/vApmQcbxc5tO79Q
RhjTyDgh31Q1pj9raH/8k1gTR4vMu4v0UKfZ2GhGfr34c5oOph2pNvSFMccznVLnvJdIwE9v7NMV
JeuyguKv/h2177o483vwNGQUBYzbPgG/OvV7vrFdS22m8REwjeNf67r6p+dUS03KMIKEpmCf99cN
OjnJM6ti8lQaydUCzg1QKOI6Lz/8FK5Fr18w+cY+1lNtr547SFBgjhYKYHwATNS08s59XMK4+irZ
VkDqzKTMQzZUFsznuJFpo1c30+4YhYCFwBWkh3utqdMXi+HZBIlgKIm1h4YN+aIY8TFrcW5XHX5y
996HEPBYB0TAyN1+ggVh1Y8vvqQLkWwivfbtaxfMSDnvOIt9ZB00jluc1rlDzHB89CRNRBQG9Mfp
lPO3iJBhKg3HDybRSkP3TQGQQWkTioCa7QbjpIdaNsSusnSVOUcP5WKKxupDc76SeFwNZnuiPcHY
DwBBU9B5pBgsbm5ojcN2BiQ30NkB891K6xxe/Ikltj6jCN93O9BTZOxQiiW6nI873q3XkazvucqP
7WYtD2P2bEbgtCriHrG9XZJ1yjsTAt1zyEbxMES7qHoUdIPhK71Z4OC+MkK6yMO7UKNyws6jHx1r
qBo8t684d9nMU2czt/45Rq6DjLugkT0q3yDujMQ2My5FIz3iWt2djKyRZBQlJ98vYAJz/ns3SYwc
0iZ6Gt/6oIjFr8rZ9JsrDXyKiT8joIeRNeKInVzl0qEldOYsX5nIkePaBIE0KtesGow0vRoN2C9b
bP02o4+2FxZiA1V5c1ZrKwTPrH1Hz4B6Vzte0qQthxwGepEhEenoGXQnhQyvzheHFFYq8JkIk7CD
96uSLFmoeyUjF1UP12HL77Ox7sZtQGDgVKMiXUOIocXO95aLvnmkSc5P2+ob45PVDg3klAu2DuS5
Cg5T6v2xVVnTG7g+qTyHsg6NwsPs2aUaN1RhaO78heYrfliIYRjvG36VV0XcKH40fsDs8xohvaVX
W6IccDFN7LWSW8Z7B9wyckFVpnWjtRzdtrbgIUNq/Hgdp0CrEULwVhZf9rImOxS83BzlgPUEZxVT
1PORhQS45eG9Lm2DLApAHNM+iTVrc/mQ5NLiPRVdDd7EGt0sci19ENZQKmD52LoOHhJ/5HlN4YNj
m2Fr+0cxT1WUo9pRvq/t2uUjAxh2UP+XHm5m+NAlefoT5zpayR7YHRYG1feVlVbABMBWzFzZAP8k
azTcGQzMWysk/Xojr5SNbiEF7Px2aI552A7GltaCUMYo4wzfUZD4buKBgb614mZ3VnGRvGpgrQG1
xoIbXWQZctkejhjhiSVNvoBPOgWQs2wqrLanAGLeE+h231cmjGUdXn2qeMOirM9y2F1hypxIlzSX
j3uvNAfT1oALVknzBEEG8Z7Ys4I39LIVOz/fs9oUImfs5Jdfkjt0iZFFepy1rMPX1y6OG1voESqu
xro8RP2TnYUpPWLoAodgd8yTktgFzqSO/xUWQ4rVzD/Gdkme/9FaVPU/7dKibSUI810n6QJLgawh
k1bxWELGah9rY1dPRrpGgNPNTFAu30/o7ivRGwwpEZqscC9RLZTq7KtOdKP8gE4A8zljhDsmvLGz
oBFuibbQjGA+nN+nPwNrUhfflIble4AK3gIJk2Es2A1rkcVkmkRma+UU/z+WaeTeGCeKp1+3I1k9
vqAbbdJ/aGOU5oOUNJ45P3BLoC4cBurKxi2HGZZZV6mIiMMkzRI8zjKx4ULlh30reY5t+pVzqWUg
0SHjSB0eWgYc4EW27lqdDgK7vnkgUsG41rD4i26FXXpByPDY+AQSQrSXviOoif+XLxavULEz4gDn
x5d+znUPfxMvc1PDNP+ngEJZqe3tdeEOIXi3z/ZoT8dcFZxKeoPZbZGm4VvckObFyTkF3OjHqxxC
MPBIbBI5FVm/FMJC2WbWLrRxlW5Oqf7NS10YB1BTgp3+sgHaE0Pecl7PMoKGvweKLnRGpWY6rpAK
xzhAcWb3UUinNqlgawyh0KyIOR05A3uk2ClwMqe//ElNGCEmNy6VbZw92LqYs1dLQfvH4yeB9xlc
+mZQbCtzcOwYiGCVXX2tR+sqy/a3iSNxl3wD3I8Tdz5XIcBixhH6JKsgRHU4oXP+FSqb/hrzO+Ax
VrbHArhyIMImp4KGWXTqWd6exOFQj5TvE9SbkAN2/GBn9g6kEAuQXK14Y4VbeqnLd/yh581xXPSG
6KZxPNG9NpcnfXOnTcgKG7qSzryPALSgAxjJ/qWRUcMrAITD1RZXnyLzIUohwPnUwE6Lb9k6bJij
6JyuNmx3CU/uoKIvYlysZ1K9De04jCeufJHlbkC/RyGx7/gnJK4FNJeMGkocY+/6utY5ijLvxKoD
x47YQJVQb31H2givkOVTzYmE6FcaUs5moGmoGRalSf3mOLP9xSPPbry1NkUX/k0UkJOUgSraRQIi
KJuA/rMpHzAvFypJOoSYHvInxIU96b7z1bPT5z5ahpV0wzIPYtphgY5pmmiz6zQPMJviJ8VL0Y45
yf18drqpsGNnsGFtMdK8i9tkkeHgXjPTQKafChNF1N6a1vx2nqevcQFo4Y5nGUBh6+25/fuuC427
uFeBC3FeoelHvlb4Pm66qvXk++5UjUs5y7X1ntcC7vE5aqG80b5FwnpmdSUnv8Pvf6QZZRLuYnEl
nQJk9jZyJpdiWoB6XL7wduMbI/st4g0v4hOfnhS+r0t7O+3NPk0lxu8pLuGdjlA9Bhi/8As2Sy9K
x6zPZqCPWDTampAXN0jqE3eGzZpuMLDdwV/MS2on0kDLXB/WozGeywgyuNfwK15IEE+equbz5U2N
q1CGU7kHsYPyCPF96LNT/ysdYAQ0pm3ljAkKN7WITXZTwDsww1RSp2e+LOi789Z/ApuVqAoOgacm
typEtmWuTQ86B5qnUvt+XdPp+IN6+PnAoVtGG1hpLu+IMCaMfanbThDfxjL0ui98fil4lolDUIlr
fWIUL/MosafCQkAzrRJDeR5vsHce1pftlcI/rovM519thRGCSqBPfcDkGo6Q6vVY3rkhThq+GG7s
fKBeTrBOONOBP8n3Ivrjcc4PuHJ+x+A34tQe4qS0AQIK3oAf4qtMaC19RICYl7jPjQ0nSk2Url2n
4DZJpQXoxc8c/+Zu0WZl8Xtp3jjEVTQUiHjm4wmgBx5qVks4wsYXFJgfMeLJi1CAu5SfZzbfjqu0
l1OBImvFnHZ662vX9k9iDmwU955GP5yI+JGq4/4SP5+/YsVlYnBARh9RfcE27h4tedqXrHYVXukI
+7s7TnykDSZ7a9VljVFMlRdHV9/OTOnNYq/u9bXHYnNGrj2u3MfgIk1UOKr/fYaVsF1Kgcz9qK5w
peBCdqVa/N4IZ51QyI08SnY3ItNdktS49hPiRE/34Y1Bq7MkHdTxPFx2WXxx8BqH+7QJjMkKam/u
e2aaaL2FA9KLZLaU31gnsdO5wqvcDOZiRLUeMNe1B1HAGk1TwaKTgwYi6ZZDOOuYETDkGogDxj5F
3Ia9weeqW89laslOXek1BMDsiqYlFFqIelPRlWuL1zDjZmK963uuZT54fMCwrp/KrsMUJSJPcqAw
Ng4yuVO2NTDrNa2eZTAeVRY9foHbcQ3BrN8gYJ1cQZHQXpZ4CAEKvpe0HPD30gBCdS8riwFvpdrt
MHS58GTezuNe0xaCJZGmv5NsvfE3d3ORQ54S7AJCtVz3QWDhfvDf4+9Q5AjPLxggC/1+Xx6jA4F4
flLDMaaqB8e335RE07Lvv3WN/NzprPpKPkxVUk7tgWK9loN1FWNT7WDJpn3EvzeDhxwc+ulzNkHx
M6Lw+tTMX6JnwuKpzGIWjHtFNRdjsiq+CoHU6yWHb2DkpJHI5JyIyUCpkoLyYwC5TEZKQj79ZEOY
EapzMmYs8hP4xzxUlAaNAkF0iDVqESylmytOTYEGpz5K48TkZ8hfl2d6mDmsJv1krm98UNESM6hi
Q/wpEfGcslQvBBWbKSrjMfq64SCdHR5So7yDmxxiyuPasClg3qzk69ECUFlcVBSqoQp57Is9qr/d
jBbTWN1XGNAncGwahFLds+GxzYBg4Eg9KSGwjSDvVSVJJ5nODwGhbnly/SwiE5+bn07QWlJLkAoO
ASQQzS7O/vk9FJcp8+HAe6nFQl1j+MuvbSkXkFTHqwDPi+KYpNnUa8OQM/A7qJMZ85aQIltsdGFv
91i41UyHaGdGRt23xiqH+JXxsKldIOAAkHMRMjglTr3+3TCFRumHqNmijTgWJb2JNOmIEWXPETc5
fBS5XULIjm4hIb9QTorsuBqjy1nDONWdfE/NZXFbjfBbK3wU/N2k0u/7cs6TCDkQ54b779ixge5i
GsOkx9tUNMzX7hYHw+RGvSRIn18gZOAoJepC3Oi/PxkPgx6qHyuVSb0SdBv3Osg7MMArH+DHKujb
u0DC/9PO03WgFf3wBwV6QWpxnVR5SlWDRO03ZBPulbHjPbrl92KjjhLdPr+LeODChOl8MoJs4JSb
vPnt1Ojx2ddvpeULI49u/E1mndM2n/hRgGJ0tW3NpCkPyJbmu6gfmHx6netFcuFcmdqT9ZumJhiJ
O33ZYKAEFl1j6Ra7GyrOnO7k5rGA1dE63hm0Wfqbx1tp7vcF5CX+VyqNAB2iG/W0kUw1PRGie/KO
Vi/ALo0WONgbCEMN3cHh2nEushUQMZT8pD3fFBDfCJFnI6JtsXeEwo0qlFacSvDvjQzqTDX+KwIc
A2bLCu3WhqFUicB9WQjvM83BitHxYQjEp2W1GXIUUiic5OPRxHxjG8f4itvXy1FhQaU7FZbNfyrq
LvqOOr+ABPXRzmNzeUO6Y8/HR7c4qEBy+BKy9NBWDN82UJNKxgBKtw45i+QqVUcU9LoOwdroNJal
vSmHs4uDCIOrBvurvzTrDeLLJzsrU3vcZKxZf8k2J5XzU0uVhug1Htu+DIApuTeML9i2Rl3odj6l
OLM3JnCflt0rBAooqFq2aQ78JPSRBjFzyz1idihrzN5qdacb1fP/G8ji4NS2ZzvN4p9ZPP8F2QBM
2fQGTaPFBKskqDK/BAqfe9OqJKJs3WRPqLa4DK/eDk8D0FS/9VqJxlZ2w3ChU7hwiIxdTm8WDMwn
1mZ5Gmb+aIwSVkKq5dyqGM68OlA47SrGiyMMP3S4Vn4ZscYGVrHuzw7K8kIRKYsgjsb9SCjQW3D9
QP16zaAr+PQW16HyAk6SoUgv7hEIqpMOKm7RpykIlIVDTW94mGpbvl7XwkDPRh7jVBvtnqW/D+CK
1NYVad7jP1vMg7Od9JciNU5zHl2CNDwbXPxTZQBSP+nPjOSgoX+AhRdemXZ6vWKPTb2/83cvhb6h
j4Iw2nhhV2goakq84kfPZFRYDUBzt8pcDZKNqABUz93N9O8wRUe8gFE9c+szzu0x/6LzVQCLr6qH
JKtELHAzmzcpOkRHGL3u8A3WUEjjetM7zJFVw2xlB7/m0ePF9cwz5cE4wO8DAj6+9sgjAaflxyGc
DXzZvvpH0sczb4XyHMnM4uAfXeXxcIScO2RTCnhOnq0CNdAKFAN5YhbN5u3tbhem/6PN44SdTsNT
WafEeRTcfO5OCAgoB4UHxXA2DibC5cU5xTbcMtdH0QGoZDeyXsWn6KyQEeK7XwtqjZ30XcmdknsC
C0lKbgMevWm34OCX/w1FHodSnS+W9qqf7tmGcSBAvAK+KNH4XSRono7RPD4rCtdeznGMWAClf2dR
87HGIbKFlu6dJP7hNbuTOgt5o8Ls14ERSDQMuU4U4nNcTZFqQfu9Co2lbWFAdRxPDxS58A357A6C
083e/yZJWKiqpOqlNX2CkIuly/OxKdm33ukXyvg/A5B3VhljElpaHW+n8wtv27DKU4kwGn7wqpbI
N8H9+HLbz1PJEm1vputPN9uKCUACvEnCwDJRrtCeq08eJE/eAznJXHTK7/pBqr4HI4vpXqcpkqK3
GGldYEZG3IsgUK53xlg9noKqw0tMVY4lxCcoSK9U8x6PG4y2pI6vnyWPhjueSzaije6DCUKaFlyt
NVEz21VQ4kv1beRgSp0aqcoXZbMiMTGOSc9BjdPJxxctI+ZJJnVcxIgHq/XUh4ZwaBukIjIwTBty
8SJ3ace6m3nXNbFKlE4/3I/WpjnfcZrRf4IUkIChWHX9+nSnmFZ+1YoN382jswKGOXFxKroT0n9Z
tqoBgAZTxjlodsgwCGvuUvdmQoQQ6n7qo9uVwJ+15fwcgOiowjDDEDM04M2L0pwmiNgxGIhkgF+j
FmGq9Zaw0kzbq5IAF8WaC0kXlnAjU5jEGuzHR+q1Q3YGICWZUuPEtwWhPaSS48ROBgLQKLydiTQP
TnJzBZy/G6s9nWVAawZ4nWIvvwwxrwU8edgbygnFlE35YzSiG5tXZ+Wltw8R50pd1/8AHMIOqR8o
q/9lRgJgU9SuCTU4CRTXEmqOIQD1oJSeXsAwXkU5P1axQQqgDubi6DXtAzl10ElYIbtSy9G0HT27
sb/mMJooEAdpwOu1QlkHHC2BgUC3boTh528dZot4XZmM2VjdNdVb4leJ2sxHhkNL6K5qJmepRaMN
WCcISmaeZ42Ps6k5YIqaODcflCFErl7qrd/jDE/o432ylu3IQmYkDm7if6n25ifDVGhbwwIAqEu5
LQ0oaYTQ/I2ay8RIXS7z2CAs1aTM24iXxsV/hmHgh03qGIdxooty3+bvipZmw7368ST/3d9N33sW
dLCIj24tt7gVNM5m8Gq3O5QgLwOtpUshW8ofcwefBvyDDugMdZMVBuuuLjj2o8otRpfw6AK5PEqY
oapmpAnFH5ey50fdr+ULRDIrkdU/x8XHAox/cgsApUAUPEExq3bweNd4AGcaPNSmhlZE6xbakw6U
iA2T+qbyNgfRfzPUCcgoP0rIJpTiKHNljNApede1q1DFHmbipYZ7/3j6P85tVbRGEUI1FRXJldMX
tX2//+u2PYJ9mXkV2D78DQHjtTk/op3FHE4nGr2EFGOBQeR+Miwro0de+mxDjU32tW/rP/vnQyLH
q+r2ue7iXH5nm6IOw7LL+GdWRv8LN40syDPsywGsGl4qLjFnrvgA38byXUeYoO0ELhpg8mEyh/MM
Ejjyr6B3j4fr8VlzzEvghShXBGEphwnhMJt6WU079ZS6vIRr4ElxZv+qrBw+bpl1VVHqsG1e8eSv
b7BVLOqqbNru+uJZHhJX5/LzCexZfuHQkZ92v4O7sn1L9Jrc0rZP/S1XxlgXuCCF+Ukr1GKIKoZ1
0HrpmODONS+UJCC8I4X+NiymY9hiUewOnP4zo/Lmq2vr7WrpgAG8TQoQ+hF5bceAH1ZoFzQYlfbI
qB5KjjrxLKkrOke/TcMVjoOSyEuikb+fKjMrSj683WQn/B+TZ1sm5ZfKGCcbVYVyPdxzJGv4WoLW
MS1vgqR6TDsE4guNUo3zXr1EVfwYRGJZ5mW19pWc+1BYTUk+jQ1/K9+mDlvxmVXB3/mHX7FoFukZ
UTkxTKMsAP3CZ8QYpRM10IYbrsADXwbu6szr1UG4TGte7pM33U3dG2DzxQ97y7ODPK6jdXiQbGg1
63PHWlbiTwA51Y4IS20WDLT+SAcgKsXR+Bft5neXXAQljsddu/MPHu1XHgufaIwLDErvQX/9N+RJ
sjxhYJECkohDjK6LSCuFuicK27igqaxW+lDvGc2QVRCZUg3uu/DPY/IHZsC33Xt5vMdIeufJZBRY
h3PDERCeqyzv1rEBREd2rdk7ms/G9xAY3W7H5U4x3wnZzfRb2bbsx2F9GGe70tFTZN2R6nmAemnO
z2VWwY1OkPpyVEqI41yMbxO53C3s9HleOvQfuM6RGsSt0XYsBNSXpUjjO2OfOldtbesVq6/Ya7/I
VqeGiYVovulqx401Scm0UgEzvXgsVJitjzCL7FNao9ZcU3wtl+LXk/t4funkNUlORtrXrhAPTyhM
xPT/55HAqs2A0X+jjtA/WSvP4R79Vk9+m4V6a3r7835rDqQo6gP7nT/3UfZSW+Nur6LOohQuzPJO
iiqQDle6S8Gg7W7DvQxgWoUfqfuhSIkgTVmafF+c7rGJdQOl7LSf8woCrt0yEIvsHWFrKMyCV+ZV
fB6tCjwl/3E0L6Oj4lf+kzD54D846UXv+UiLzNS5GJXsAWnqmqkbQ04ENX9Ufd5VzjWVA1YqlqdY
17ufEft2cauBx70XzbPl6JOZ7ha27NURjcJpXXDrtC4CJsP1UYcbZ2BKn+VdtFBrcLUHet4bFN2/
aQ1swjz2CviDrRRWfkkz84XggAHXtPp5kUpCZ6foUuw5H+fj9IlFPn1o8KvH4ZPXPkaob9G99fMY
GWKWOdyih3fqyh9WYiiwG55Jp1udXrNIgrzRfbK3iiyavswLKY2qkND2NjUh9nx/JaFD1CSURxHL
x2zljiWebeEUmhnOlqvwUVyebejba5dzdxIoYxKvgN3wi2BwJn0BIp1SDOAaA1VDkUq8jYPPLyyE
n8VQKHNDVpnUvxFGoTnqOnbChCCip0D8QtEWZI1AryqTnEb85ZfqUD1afWrrNylZvgCey+7rQ8dt
/JiHTk39O1pCHwBZdCMEQ+fumzEnW6jLEUGbJtAHZUPiBbqlfcPsgow3Yc9NxYaRV55CEJ1Ya5QB
8GlZ9q+mtiPdN73itaPR2z4Um5q2yCwQyyEEoBFRWFhvPBxRp6f1W+YvWM0sCr2uUBzo+i1lnXTU
kAlfCfIBnGJOSXR7LS6fYuluVyUW2KAEKKEFa9XS3OAky80UQhw2l6u1ZvytRebX9IajC2quqljc
Dgjh3gFn0s+L2VET5J2bb4PeI7Fdf7+8JVLAQy0UTeWB+VhbS5/QZVikzpCKYMGsxFrRplS1sVSL
hQ56mlgXRU17SQtFEnHN9uPMfa9h/AMrZILyxei+k0qdLFjejT83MUCHrPvT/QsrbDC6SmbppCva
E1xi+3vRDFOQl1WrE6zt7IH9ak70Qjk2g9Q8ZIrsOkH+2pwQLOhkH+qPVkTgXX4IqoNExbr63Tk2
xzl5VM1E6X/nKW8HCYEmdWFF7/UdYC1UeSjF2+oYrd34aczaQ9xF9WPAGCHWNIFLXTJrl5jx+g8V
9JIAKywPt0NTOVds+LQwZiMfCZGnahY4l56dLXB+TGxWATHx7I/yqw5a+wyQn5QawWpsKi0gWvf3
j0TkJYQ5HPtOqFfmlDofDyVaSOVz+1gPTPEhtVBzAB7nl5zv3e0TDLnBH1IWCf9LqitjMo60MNgC
4OUnyOfoCxNtL/TvzXao3cIN2/1pnkkgqbwG8nRia6oiKCw+mLXeQNiwkdres2kS5MED/oLzOkcn
0byiLNtiZWl2zmccRzU2nJtV+j+JKHO/Bq02O0l1W+oDA4h+XY8AoeyYcHVcnAnTh/Fx5bbRiUpn
9MaV1C2n8i7JVu3ebSACqWEpiWSNxdSKdugdb4ZhvZBMPFAhQC7YnYu/jAC6YOr1U0JKG4eTyTUL
lyI0RenMDF4/vgnFQqBJC/B9MdJB4UOUjfu/Fgem0EsmkFOB5f8Y7VD26B3btjEjTqVikbf8Xr5c
0RYcTqLZ67H35BKdjbb965Q5U/0xxpO0TNoLa2KVWbPajBlewA3uyQGuFIA+NG+cos5dgebqgJLZ
ZQaKmTmabPhomJYpv8EnpCXtYm2oVisap6pXk5D8JikKaF4D/wa3o8EtFeQI6yrpmhRdVHvf6d2u
M7F/zmrlg31BDWdj80K+dNEjlnbFEnUB6AakQSWg7k9yFV6DUtlgi6XAuUHi6NB5bez7Fv11PM9w
eqbVYgOwBCP0cnbQSwyFefoQW/mop5fIOE0jZmcThJ7Y8QeNBa0TUU8xeHieKHHC6//NgdB+cNf9
YgIu3LJRd/fcCZuI5YpJa0CZ27mF0CaCbxu6GSI2rRlFLO41R3/ZSaPeBNO3y4Mbk5rCOi0BycnK
1PwxG2cQFqIC8RxIKCs1dLpyFhQoPlq+18lCk4HCpfF/sI8B06Euul6LpP1EQ6VWmqjQ/FgwFGke
l82u91Ki1ty6Xks03qHVBiXiYR7xEZprOYIfwC0DuefM24/zLdz6J4W4DrxI23oPvivnvXuy6Aqu
rrLOa3I35mVBI5FkalFcuEovT/XEepq9PSA7UPQ6hxROSq9NUbyhIuGHdiMiEH10xwxnvILcuTh+
gTLYwrhLpGN90RurfOhTXQ5Cq0ccarDKD6G9OK4bK+b8R0oa/6qkNW3OQ8rSB9QbUb/nefDeynE0
vKylWTLvY5v1ksJqyKAOCuWyeqrgFyMeMAu8TnnqDO9S2Mrx3SY2XEjiw++OgmndvVUv4yREsx57
Cbv6HGjpQ/M9S1Nqp4pI7KON7vyqZ28D4PV08ck9C4kC2Nxg8wC4W6bkzaRGxcTL2t3fzs8HsXTU
Yf9CeIgaCmESupu/pQzxIDGHvSeuyt0v7XU0/QLBRrWPJaVqZLzKxL2PPdLvUPOBecsgZbNIk/Qn
w9WGhG+6KJnFa/eUbSo5cvBNp4XBKCHY0XtYcXnGec6blPpEi6WkaVR6FT8BKaBKmP7MHHeis5tt
puoAEK4NZ89JDoXAkW9fd/6vZXnBwsbFbzuNtwsxezCgB2zXMxDAnGVOSwpZoDomAsmouwvj/hCN
igtydoFEobDv7y68scVN5rTAvTjIEqqYz8LKZKahgtlBxJ3XwcD1v3D82rpjn6J9KhmYelQP9mVv
DJFRBOhGRgUuTMUpn9/Fm0Xb3MfxFfaYk09wvhAxkWywq4X19Ogy1TCtfNJ7ZLuWPyNJy0LN8GYw
hLGN6renyYzb472EO0a/NHF/32US1FCNhE4vCPMypjx494Vr0c/qDHG5CCE90cY0ICBtTdDFPQWa
dltNMRFI/3nx9lInjUkFydQS5Tz7XqWR6ip8d1Md5WVcLeoIkjN6DQ4cfD7hxUZ+DyxWu+vrURQd
nyqNMJPiXL8HfptrZEhvkgWA4BShRqBpHz3kb9yQF8e5DSSM0MY3rDse/X5XU+8RXz2atkjsXHOQ
FzJ0o9Uvu2KzOhWyzXt/+boa63Urpy6dLLyhDR4FB5AynxGW9ImxnTswRqFPADxMlokFQOX97YqI
LlMdt4I2YQ4byBhwLDczhzpV26E8302ZuUVcethShY3Vi+MY4lo63yKnKG+Hps6fdDnN23RbCVDp
tTMDRGSPFgg5wKW/Y5DUtoj0dzdKm7HcH0+luAqh0Z2O2vl/DdJe+1LR0Wpz2Wg7g4wB13S8ODCP
1mecHE5IiKjqHykrOi3Lzc6WSOrGbtdIymTC1OUtP//3b0/NHJ1KxzmSI9zwGhd3JS30eVYa+jfC
C//ReA02CoOH1mougBc4kj5pYoNRDBeogJNCjVljRnsWJgbN7Gbt4/RP1W0/uuYN59lhAz3UlxXu
qM+5obmh51Hl+TzaApl6YP3IJc+0WSJzFoxPRjwq0E7XhfZ0vrZovpH1YrNpRpmkWR8Hn6WWutMp
rD9XlL3gUVCJkFqWzeIjcnOJKiXgrKYtCApPpz+PfVHoyM2Bsgbw+W+RxqMA2UP84dCW7gw9eXdL
J+QLrJAdGknPG7WEXfL2L0uPCxAEq8w8bt+IYvvb85VghIIFElsbdFre9C9yMCGEn+MTq8Bj2M6W
wxT5HGdhx+6AjCNpNYALHQDboNMuwe64GxlNR9+TAgVqbemm3KFVQoj76v7GX+Wv/lXllxaUPn5N
OivPZT4pO+IqU0+/A7xrBnRwY9Ti82xmkoHxR0zbuZAfBeoCoMxC+v8MM8+XNVllI9mrurk6C7PQ
ns8qL1fzcadCzrGjBY0giN6KtRRd7/Gn256h7DEsOl28ccA6eosePJkUALZ/N5kiHpMlt8kPKciU
lU5821qjydmF29IIx585vYmgL3Nfw30At3Q4Fah3bXr0y1qPbgq9cqmiH4tq4W6ZohxbY74tRv1E
ES6mygNAGF1g6OF104uNYPcY+dbDjayBwXrUCLnspw7QQK330s+17/YxqqEn9HRjbb+30RgnJYNr
86s4/SyHc8AYUOmmmnEq6AO3BS46MkH2K4OXXtm+QR7TgUpad9m6R2pjHcCla7v2krGU/ADcRCQN
pESZBPt2YZxY6PDhlp3CGfQvPsDeGiGD3zaNdk6pWQR1j3OurY0bUYJcuHnnTZWGU22vNq3sToU0
kpeTOM4vsUZfITp5I0BnatfFTU6FkjsShuH+JsCspl1NROuC0iWlkE8zhnHzdO11sk5JD3kJwV+e
ZDfmtaBpm45wQ/ICZ6peOPEvq5YL+zMLfRI19ibUz6owQo8fG0xMn3/x/2QafYZL5FOn7VxTt/Y0
dSUucfFTpshGzoGI5rlt6K8BxveXopzqqjn4Z3mZRAcYmdDgCq0QpplPP6q4QpV3jJbaVO1YawTY
NvxSqcoE6vLv/7eONWvx/9H1wcz+No41LolEcJnKR47EqDujKrfFSYewEZ6+hFQUZWT1WtzfAzfP
jQnfhbLHEHSIDyczHjYKPXT+MruIKXMud5CPlLTsFVQPjBgfJlIunzjTW3ZdbOYShEtISkUYz2Sb
dLF9ctWTVYDzI5gts6ixVaFxN2yDZKkVWOg/4lnBiNhWdqV/AfhVfdLj9QfquVsWde9Q6LIIe6Tm
j3Zozn68y37OiOwoeUEqoD07D4plKePIQTDyhSucmhijBs8V0ItkO4QlcXEpHu7NvXbw5VtOeKEX
G6310GmMVsCeTMOSb9rnPt3prlv3nwrynm2ijDQ7huvQa9MuKMwEkhnOp1qohTYkfzVHNEjurcZq
ini994scgzNNSTtVU4eHKznoXjSXBflooGQ49Mz39flQBCaUAG1qudBz9IxK0MIkmCsIbAMY0V8s
H48CItOPBqbLrh5TEkVvMTfh3dJxEiBW3whdlL2DdXBQ27liIlA641tkuA06TkN89jO+8HJM/guX
3ERNIw3B+JJGL/PijGPJ8mtU7FaQ2f0qsoEgirgnQ3L3tavyjemOVzbLIuhfcau8rvcoUc4pb93z
L30b2cnFm0okxfIUVkvDZ2LLvrD14amR6Mw895UhkTHfXHRDYJ2ervvda1W83Clto8p45n/nLKc+
b12vbDYj4bXsluE4E8ONfiXEnHrozxuhtiTToIG4DZ0F896q1/aPw0CcqT0f5KZppC+vxtIL0p8l
MmexQAc738iVjGJXVBMmYpL+4l3glMGers/iXMgZPt7keqgHQikFjowprSCF1ibabc/LpFln6qH/
mkzwnBGoDbaGEqzVVs+I4N0mvMvr5nXCzle85/B01ijn5mgbbNT5avHNDh3w0JSx6efnlZIz6a73
re3nRWEPpaYqJUHNApg6DXxWe+CH0FEA6EtemoS0M0pY98p0xthRKx4BrPNvoAx1qv5cb5YJC3f5
JYYvRYRzaCgigqnsBMu2YcdwHsSjB9aO32hdyUC5evWt66ek5fyxg8QtP8wD315qkJM4xGT49NrP
drxs95o9qQJu0wSh2WccwxUygOiEcHhdx504zkhkohPxuSCi+fGsVds3SpyKExLFSUHM8o7rrw3A
HXAakF5ytTgZ/hr+6bR0kFUMLA+gllTS9G/F0+1Cq31TmRyYsoSxiDPy8mwnAjDosLCZTYOn/Mcq
TYqttvAWLBdh6+xZwhcV5GKEnP9tYo9vF8Zd2L1b4Mdauc0eQ+TVggfgm8mwqGmpFwxN7X0bcFSe
pjxqwTnNg3RDR4A6lODW3DErofmj925xnQKQq5LSK9PMRpVmloUFnW4vla8uFtGoNK4RU3F3acox
zj63mFkRRvLW8ECgVN8N22W1H2Hi7NaG5AIh6hp2pyZsXa9za6riGi3NCGqlLsoPEX8f4Ztjg89c
2HYtyJyZ5dN0k85P6A2FuZW+dZoBlhTu+YVMQxzMJN7rEsHxNmKkj0xzLtPoANcnSvXYUYOObuK9
rnHIpWV+IRUp1qB1sFr6Yjng4F5OtfU1oeyxVqVt6cgmUanfg98mBkkGnPwAt2h2NnhW5Qij0nmv
L6NJjURAbJNZmVpiaQPmoYTdv6Wgbc2VquSmYJwbmmghu8W/z44pKvtfT1nagz+HNzNTu/uutQVV
MRrRWrus9fyaK+X/6FWuVwhvqKPW8j08eKcgyygd5pNf6ceSSeaCK9+gUe39lqbOb2JrC7sdCNq7
cRrBlP3svBJaZFBRQGnM3hWuIVMdoxFmCZ6BgV4YmhktXI3EIboBvcGvTXoPcFgHWgOQ+DOmkZBu
qnkmqQHJoGZP4uYufoOXgcY5IAXSYPCz22j/tZNV48TGEDHq//uJRQCUNJd0TMqiubBN95L/h1Mx
HnXPAaQ4jOFiA7f9Lkh2vP4aEpdb03HfPYQD7M+V+TDB8/ES8FQQ8aFog+YfS3friSv9LGM5F3ES
QqKZMufnwd4w6VOjqCsUpDBFeeajMA35xKjwgEmdCo/ECxuWhtevZ4Tg9NPbYheJQjJ0EHlnB0J/
9B1pwj6FmFQynK0i9ylcd83baQCfnxnCb7qW35rNfWLBfl1M3KH4N9W1+MDzdmsYn1Ox3AqZ2G4Y
pOgGxuRRe5OgWioJzb1IOfFdvPtAP6FPGucKWVig1SP3JojkFNJ77WbhXa1G1rkhdRYwW+i1Sd/5
l8TxtLHdM04E08jTU2STOo+39z2VPdK38w5OfwTjsBamW72WU1jcgtsaBsTRSB+nRvYUs5BoRMoc
ljpQIKhKSQgGj3jQcx5BfERQU2BmUF5/bzLuBKOmLyXh4vmQ76uQ2nFv4xa9rtblQ7zv4vVHCxCQ
K/BVZKC5r2eclSpl1prpA2OVfFioHZkWNOdU9haCEZpajIBq9ZA/gtEuZ3+jVmlAw6DCfKr1+Elx
Gm1mFWXBFBHKcCDsSMh26yzw6KDTkwI8vFk6cje+PcxKKmHzhepBeay0tu6VZY7oJN8J/5eCnTn6
E0rsT6IoT+XfA/eQfxwpJi/YUJP/xoRU8kW683cEBdSw6ijjvFePQuj+84bQUzcofJNab5doJPcR
daLUySop4Z+zWj5+fpyAYH7VnOmMDF4VHYIdhDsUwcqoLkMmi5ncawXmT7z6+XPNd9ncq+vIARou
pq6G6ZQo6kbT1jFQoJHGmYudrKGfZskkd9P6YEWNasVSfw4MPnyePA827vJWJtAEJRvaE/XRUHGi
MWjD2Jr7HFLbrTILXiQKtC+gkAEzBb+eoIz7J2m0b8Cgp4HHp3iUqcmDovU7cpsbrUEDz2R3/afx
yzypBmV4rSQ5bwUhI7bKWz6qqHTu2YtYXNKOef0taVg+DUhuh5m9nwwS6Ejga3SAw+9K3Q02Nw0S
RcKXNcL29ZqhsvWcofMIPPi3XE1MsFW28BR/5F6VhbFbNM+bD7x4lO5KHW3aLExElk8t9dAoUmzK
+7ztUFhQZM62KB3YL9r1rDfmEwMLXjDKpqsUOCJjZWmK48/5T136zcANnXkwgM+XuamNUxhU6CBv
EyYk8BcvEVQZ+YX4NdnccI5yXmIG0HBJF19aWfr1uecGuA11Hhun/0I6I572T9WVaLY9t/uDlaPg
Myf7hwqsU1/YPM3IpMKTOmZvFOUuZLiSqwbH8MH01AJqrHyHssZQ6XzpqTC08TCuASPPF1PCnJju
mvvRYq2gnoNuaTCt3C0gGUYF/j4xhx+TMwu41+5d/YreeusCi7a2i6CiOA9QSie/iE58xlxByqsa
9wwp0Z9kkHijXE3r/z73PfNFbJHvlnx56VQYtkfb6ORs0hTAvKtKtgimMa0PzEVJcGR2DRKrmF3M
0ELnPViuHdsDWv/+t2WY7uUKrGc+IGLRnp/bFv9IRn29ClUuJJMAKmmvIpQYPWTMzLrp0lkCgqNF
qufKV/x0gh/0Hysc+9djoqHgYbxaBByVelxzhX1PaLxswRNyEClMr61he23Hk2pH9knuJEOMBT7/
HkWlVxUdAfF7W0ChdwVwzV3ymTUy0dleO7jNcqYq2O5+ELRnAtIEQzMAi8CHdjcXqsPkQGfrsFFz
/xM+rqt6wVhOrdILBsDraBYnmS6Ov4jpW72xOAOq9xKVPZ08zczVujdixX/eMPagJVSsaMyHFnA8
6Z/MWkS5LPG//u9jj9r2c+YyuUMiYivh37N6JFHuFIfvO+l4m417rfFulqK1zgV/HzeUoHwdlr5P
snDhjPBNdBFOdvZtlaUtokd8DdajzagtSasaAf44PvcLhV/foAZNmSc858nf/YsgiO9mqzbrBZMd
pNi5i0A2InAmmsX0X6Tw/U5UzfCb85/tLX3LOa3RBcKWuYm07tK5bkMFYe0UQpgM/AplyHRXau2C
v1noOrISw4W0tvu56qGL44O/S8hO/RT6IB7Dm7ukHRYKMaN5RrKx35P4Kqr7pVyFAXZ92YyyDTJ2
H1Lr4zQhuAys8ewQzinHKU0jKZVcygjkfPWOl6j3Q9CYy/Nu2uc7in4u0OfehENi6BHuGGuhllvM
h01RKmYptsmpLGluuDMBH3gpn4OcwRa57j0/py2eDmySbLlT0Ii+fU4FNJvc0JHR2sBTJ053jHM7
jNpm4tpyeu76YR9XUjdW9GgVuY8mOQbJBupv6wT+EHe2tO2KHLnoOiHaS8gmDCXA9I9aGkodBmqX
wqmYZo54V5nnjDeciFx67Muq6fHjqIpuSyG/oJyeOQnOG0U/OiXcJeSQyicjRfX3nNZtrqiCpHCG
IGBubu3ijf/8WMJHglnltHf70Lt0+HYFFJ0v8oMLtHWifxe6D2DylsEqIjZ60bcKrnjK65B4ftI7
p8plqkQcSfKqkXZEJUhLJ8Tarv12assuPiUJt9q/dgw12k3tsphePjSEIo8YZ4ucIBDkLk0YuUtu
+K9qPRv1VBdY2y0wkGd0FOf6gQ+Kzdg19Vdtxl60ft1YeLNeFnLzpMuwnSBJzhkCv+bG+mUjghWR
zyhBwgw4RWjCtOyLOSej88b7fsr/qLewW4Q/K+eewdne58C6Vly6Z5lQDER9XfCi/0LUG0DKMqj0
ZoeQwAxVK6u9K73pBDo3JN8Hw1jQwuwXYuUAuOj//So60llyeUNs4sHRhRAsoEJyy5Vh24HuCEM4
esdV99jcU0TQkHcZ5aLpJ835EMP2/36QFtvt9C2oj4gXc/BeCNYWAJz7oZxxjc6BCCj2bnE4SWAG
ZjRIsigomgkQFHVGboBhhCky2zU/zWxY0DbzLKJgNHfUw75TKCP9VOUPqFSGPOWwtYzq4YitAqFb
rRAfudHPbUBLyE0DthJH0oKFhUv4jRu07zksqpT+F0ejNZLBmjkxF3X3khN+0n4oqjwkstet1yGG
OWz7KBwv+FRKWUrPozOBd93Ut4LgtQKaZWRGAlpQ/7DeSFI+kSRwk51dMR2SAZ2KdMIJGIEZS35D
DafLnv/JIcImhJssrGhsuzANq29O+9zUuKveawqkygj4FfGCfuphN/lbBH/tbDCtlnFK7m+Y/vwZ
71a64jlpcd8Nw9DzBuyWTMkRO+nBJxq8HMfx6XOrZBX27NellCr3GMgTgoPg3jb5soN/UZKJpYHN
nAiywzbBEqBcb4gBlMxgVW6x3znEXFhEc6OkhzwJIoU8zdn134t+jWSbhY2gnztsJBtb2xf6Fzi/
qACDwpAX4VtuFmeWSCJKrBvvIZQCi31zbtAdbbUCgl1oA5QB4gP3DkXN6tR96xHakt0X/EuVc9RC
1DmiC+DbluZce4OOiWVG1IO13yN8MLayyfXVgNPosuXZgHlQunj8P+0g2YbHvYyRxHpYhSJ624u6
qnEETzOWWcbJjaWCFy2Y3o8lqgORGDALE4UWkTVWIpbEnaK3ZIxzhOKWp0elHoC8fWDW9vzfSxZ8
4hM80sYlkJG5gl/lwBUmQ3yUn9LvuX0RNIVhbeY+jr24x6G3jm8Momri6x+E9FwhzmBQvs95uGnP
JHWt7G4+BWez9U+P/fHS6JaQEoN9clUt3bEJJrSP5FCJLDmjnz4r9BZCi4NfcPIB6kttrcyL0YxP
uNE34IKIGjsPBmBxLRhZkQjESu412epH+aihdGD//YNvIllebldenQ93mZSUkvqQ3agi1kSy7a80
WXDohuTONA/K5EA1SxVMMzGXiZRFgkSqUWvbg/Clog78JmwzXRha3zQTnMBlX3y0NeKccR1XreC1
HbLZp1aQaDbaiSorxMOJ1Z6nveKwXj3T7a4lJ+DVjKGMTRccs+6B1xzwXFv1LjErcHg35Ix/t6G7
gG73iXDNYSHEMoKfae7xN28yDcCrsayStuHaXEMCFQ1WdnUIN7GE6jxHwUJVUtKuWcWz7qg7zeeI
zC9NIBbe/jR3cpTqEpQ5fwyhfO2dFolUyfNxN4858pL3TZtTgRqaxYXd3o8C4FFJp8Q9MviiL699
Ga2+MohSiq9TxrRtvhHOzUYEwiIKqsSlzFBB6Tb85a+LPTQcqu95Dwc9NNbFOohqvaOQi9DZMioV
R12ADzv6OKJfgZikjzoJc59HsE88Nz8SFoDXQrJ8XsKs0ldOJMHtOnuYpV1PTbFZQmPhDWk+E6rt
ygNwdT6mes9EJ2JFNJuKcBeYUUBPUZfO1CQDnU6bhu6YyObKFJXTBnLj/PkssikxR5vtXnrq+/A1
1B0+QZBWoJUxMlMRyM93T1QFR1t4p4UzR+gwoldiKyxywaz5Ndpb/NYfnDwq1ZvNidxF+h9lql1k
J7vyYup5i6UcmVlcROWx30WO0nRtzXQPlf5/tocKYdv8+ApEwbwgdDA5X1p4zAc9vz/hmsKPlRJ+
f+oOAOKfMeBRlU0webVouc0rQ6DZK4KAmphEqYyYU6C8IiEyzmezR66vvfjG5AnQKEhJXsAm3VT2
uuCZlbH5kIyOgIliSdojEj2U7xzXcVwBP7x4P3cQYJCpmaMU65pGbiBZIHIy6p2iV9NEeEYWBkjj
Hm1/K0JVI1V7EiFulSOo2XBhZvJKctJ+rus6eWtTrFdxXA8XbM65uRJGWQgXVIt/aBCb8kVlMFDC
LSij+iMVT+ujV9hXhiI7YPRAatMY7HmO3N//+ITUfiTZHSmNjU9wTIudM2kQRTvmGS/G2pGxhx6K
B2cFjcRtGFqaWfRPfmBw4WuPeKwBNkRCqqSBL60GUlKDKINXoXbJvV9yS4oh4zRpfBu8AQgMyCZW
DikSpaLVCQJ7lgqECwgWTp9Z8levdrUoBd9kJtXEcDZmDK4WtfmzKAkbb6o1T/Wc2QkF/k0mGDQQ
Ru6ys+a4I4CsiI4chQYYh5IpLoZ9vijAQPJ8I3q2cAaG9sa0YpLVREt8JK/4793SrDRuPfwTVRCM
XlR6v9ikThxGvsKtHzDrIbbV7f6qm6hEHUwnFaEQLYWIrRU9LHG1WaGRb+Ib8AlNLluFFvvBA/Na
u/XfQjxnDo2JODIVi4avsXQkDz+DPRygTstOkRMdgO6KI3wkh/NEGlla7rHfrCZF6vokjQtv7fXy
7R3i7AhvPYNZExaHhmQ6KY4dQuoPkydfr+XTzxbJ2JSZmsx7rSk2PwBzG8GrSjHw+n+qiOSLAVjD
P3ZqM4rOZq3HsgBI07G5BJlUe7clziSFEYnOxqEYvobYzAM8fuP79d6egJgqRT0L4C5fjhUjxVG7
7q6Xmpwfd3tS7+lWxNsyQ0V5pbZi5cqjkMyG8I9MgEBgpviTb6LQ/VPx0gf3U7jtDGaqGFOQUBJA
2ZoPx+4t9D8b62R4c9qvy6UT+WDbZNHgiIa6Y/xvh4bTZ90K7zTv0XFxijv9ITvbQVOX3swjIG16
RplwhqUjUY+GYSWhUCJuygytueQzqfHAM5PxIwMEpAHzZ3sdnni0jJaWcDgFLcJPimYh5yLNoiol
Sx2Gjh5omcy68JjlBfHaE5H8/mXcBs9Ml6ftpnQp29GnYHS+XLmQggCSY7awjEJScTKHJskiR+x1
5oLzlLvYRhkpz4Cdp4VH7MWQxoDBhBK8QMhXG7lRbr5OKLergcQ+s6OAB4Zf1AlQACFqzTkNH4Xc
tZqeghZV67WD/tO6LCdfm1IvlhhuOe6t/WZXnl17mYL5cDd9ZyZ8hOQgFicW6iLQBtcH428YBEQT
95vr2r0nQ8AC78/5b4sD7W6ahtwvAtNSih0PDY+9M5vLaXwPsH7JVHWtqvUqnXHkhawonRulsrFs
fi3alXsxp2hyce7c3egAZi9JLum2KOQozyr/A3OjuFrjn+7YkOVDLRruu0geStqoNbRuo4V7xniT
dcwTGeShbAIocUhMBEQCA5EWpB+Hglk9dkkFv1yG0PAo2dX7k150MHlQ0uWG1dMlWMP7WnWLCM58
MK/DeEAxMqzOafSLkjEAK69vECiccHLSii7JfsZ15/UxVNYWxb1S9PROnlSQ+oLheL+sVAVMXPqz
L2WrU1d/Ycirq1Bxoz6LgXg3Sg927usM4//oKvEIjXoNYq8XoREAJFIF/V/n/bZuAOR2hmD4rltS
Jbh4it4oRixrsGVXBj/3cEu+BzORKA0kXkYnZs8pYW9NLRyz3byh+nj1o4yNGssUuIJlmKcP0aZP
hguRU55XRjSMtvKbil9IXHZZPcWaWv+d2t6IAx3OzDsm/7DrNelOfBJEa4K32wtvPqOWJZdSBub8
I7SUIxVa/blMSpSs7kSk8heRwueeV/UzD2NllqxYcOxr1tuxlOB1PKOPJ3MUo7XaGPZVa27Moe8P
hbZ7g9j9YP7VmnD9DmrGCgHDbzVI8EA+8ZTjp2OIrcn0gbavMqQ5brHgQEZg5IZn+tqzBrDLNOcV
EHwLCGbuBfsfZYKEw4Uw8oIaE1q8F6uZLKlAqPUpb43rzdm5LZDE5/8am4s/LOuA5ArnONGsGbsk
3tGZEtDlrJE8xkSMvLOrRW4VTiofodJRyp/oGgtgYEuPdpoEvacYf0jSW/u/aUgcguFyQXAF9XBa
EA9TnA8OGmnV6jEoRCMKXtGFlG86o23rivShvz+p/+jQaidY1+Oo3CGuvUevbmk0JbeNVfqReb81
IFBaaXfA2wQkdqfBhlG9oaIw3AIRexF+G6ntM4Yns416+OQaLjAdx1BHK9s5ZPG0l39Nej92MjEF
B3Kk0BdF5WR0CTxgujzvlG6AwBockHt/K4YXomvy0aBBEAOI1sMrz6jJR2bou/iRHzalJawlDUpG
T+K2K0i2KEbfqIotuBoh8R6huhafKyfBarQ2A+3sJPtZKH5n6/J/+Oy+u+YsOAe32sX19p/jdkpO
XqNKPJ0mxwZhSTyWj8qBcQTGCn5jLRga40/RZJQdvswuAz+FRHfpXC9BuvrpSn8wJ9S2XwEBzB9V
y8wMy3A16c90LycfeKYK4H93hUl3iqY8k0+/YQLWBhLKiYt+T+KMzR4AkE1WghGQw/xbC/VysESi
ePJwkk6hyGcOYLQ+QP8PYD3s5dZk7pARI0FRC2xC5rn8PCo0tsi9HxrjZFPp/CZsR20p3XznKwXo
cy3+nooxukoP0x17iKUfPS8fyLka6fX/klcuC9Eo2kZeJdxCaCVZScSy/7OMjwnXcsiYDRmICs8Y
DCM9p+Nldd/z9uBl5pKSLrqstEj9KqTtrOntJUBrFrXKeto826OetTzBjcNBYos0zga32MIY9cst
byWqePeSw33KgiwMh/YJINVRpKlunR1zOEsloUTrQoU0EulMZd4Vtg4fR3p/svNxGwEOiszDEkmQ
aW7yQOMg+homo19toQPrFtYsObAokkM8FBVxUlarXdiDA+DiQ7r80Qll3KvgbGY8VX9UbuA0vSAC
n/Ujd4vGkNhoPa430ZhrMgbJs8oHXRDxAPDpHaB99WRNDJUXBUu8O0suzpRYOkv+luEfET1qOICf
3JSEk/Ol85Cotq/qYEm8ZMoEQcyhH6KjwAplD4lXNx2kqNKR8MMc8NzjQ66mL/kjq5lGmKSYYqPT
z4M3EGLIevsgk+joGh1S3azUpu/Qrrkfsec+n9j/KCiink3UKOpiXALd+40wguB5QrvebF1pbb4r
g456cF1G/nbmCWD3zQWITBahmvqvnE/WX/lzDDZzU5AZaVzPKaDzu87rqg0Ru36vPvGTyt2kFo1g
IwQE3SeztpeW1Ggb6SVNknSMsuf/qTyZ7Bl+xk69kjYVyrxNJHFuYav5fzVFp2t2e7YXRYbe0IaC
etBcbc0U7olcjb+yyA/DJ/G4Ou4k8qOyDTRg536sr6s+OIn2GR6L8FDDEpcTwWbKiLzq1BxNzU+o
cwk91rYEpSC2GAfyEhdB4bEslxtJJQv09wwrABDvuN33LfUvvZgj59RKvLh3N7h8qKoGk0o3mOkC
fSshLvK0zcpZNpsy2wqc5+3hbVyOJU5lX6MSNPKrC/ELxmRX/qsQPseKGdqeDUh++dhqqZyKMX0B
tfpw85qFdXcpokvXP1VQoqnE7/Ae1uwpSvDBWYZfGs4GWBHYopi/d/ElR+aGVxuZUVrmVOXcUypc
vNveAQr8b8gIj2axOg5VdGYS9A9f1Y8FZiFQobCp/MqhU4LVjx+q9lZ120AFl/eLeesajoC2GavH
yTR9BXBvqjlVLq2oNLAxOj/0DmcJRybPCXnC+728eLeg1WbDujSJfpNcNzGNPVhN17sIJLH23VvW
EFEzm+i3GmOnKEA2AfelrLT11CPF82UWv6ycUn/PSqX1JlW10MxnA6RAMWt5bISW91WeNZcsfLea
fPSoUMcBXyDd6IalxhzS6+HH29FdaUx06EEg8ls28xXP1TG0PAtGuX6wRZWao/b22izcVmeZqaZx
wVCUOYoeeyheZy/uaWWlktWKnW6RqgvVW90cRbYjnjEj6H0mQ3baM1BNDRr//rRY90OK8ZYCvh1b
xbhgjz7T9vEYs8XciIFozqrwFwxZb99f3KXQAt/LUIdO81CKVXCNlxec2B0EtzrdnKi+54hY4TaA
P9YDIGoP5XRK1GR+u2TGVvPlH4Tr8sGmRmkvj4kQeKibw1lgr9GEK9+dvr0DuFQhISzx4Jf3xnFV
1wIoFhrb8a9Fy5H9thMfS+YOZM/41Y+cAcBcPO5aQkt1Li8FtLLfvQR41Cuuu7fgZ9nmh1jnzwec
wQXkl/uDqYOMVMq1zB6sNIlJGAlq/bINNOJgPlA1Yr1ASyL/q+a9H7TyGZg4gofSf31qcANR0J48
52C67g8CKY9sGz3y2dT+YnBihqeeehqI2xc1oZP9w6XncQzmao2NTEb5t2dngvt3nrhbpfklQiGv
Y//zZkPCu1kolAjXO9nBBu/BbboJCaasAeKOEDe5B7E2pxNPcMBsoS/1QJJ+ri/Wss7HhD+4wLXe
P8nstqgo2HBTiDUF0UiIa9rljfT5FPjB6skrG3Zcm13z19OFYnw5NzKB/0Ys1CcbDgw3UZTv6Um2
pUl5ycae/6YoNfhSO47i5LnX7Y/nW3BAGFEKpQKreNPZoCf962zR+/kBBjsgUU0o9HaxnC6omhNn
yfDZvPBG4kI4qug2O7ZBQphZ7BvsCPvIPqCIliVOh1UIZuql0q5dRALqVE5Q7iogzp2gtJSjfLUX
+DY2pKeQsAtrqvJWOLpcCBro5aqD1sv3TJ6qJI8UeGIKfgIkzcF1/LQ/pQsF+wPHH2kdneuJ5ZDY
0uuKodpmV0TB4A1f0+A+angHkFJ6PjW8mrE+/zyJm5AdK3ByRb4NPJbBKhX7X5kJ0YrRd4af9QuG
Sl0ZWFfA9yru0f6O4R0gqlzY5dA897HG0xb+PicxvGLRwX5VUN2fepec2RCaKNUelpl/Gz6O9sGt
dVYzaWZ5DNqRh/XBQfNcRvlHWGQgHbyrsC8YQ1uAMgzpujPWfXdaU13ZrYb+zEMkSyAMTX0c+s/f
L3KySXq5mWrOGM+R5bdtLG6jxSVi1l5dox2RyXoBpNSJuUC1Z2PX+602Ds4n+zrxNaKSD1dBOL6Z
sUF4p0teSGm/GAFZKo76dX/U0FtcAybETMGBb1nCaJPSyZWarmokbcUDTcs+EkLmvC6wFOjj7BQ0
MyW1qik1K1sSee1fVqXxbyFxlDVY2H4oWmxWyoTeSwIdADIfzMPZTS4In95gvhSunetRL9kqtv7o
EseotlEXChCjvBDBjEMGWsVqVpsfkuTMC9DI+lQym34XBq2VaJb6bV8orSUhP2hHJyIhdRnk5aoL
jPkxjx+ZPShSfqNve/BCdmNOs33f+u1b0s0OHBa4gPmxUknwxpTo7zHlYKT3YMekO+EU400+8YOI
rGzV86PvaKCwM1Qn1FFnUWxm6cC2p9YGF0qQX8c/EnJjwnoBU55/ZrqL1F6xVrlx7P/A8xdDYFWQ
TJnd9gItqbSr/ZZzBl8hCDW8a29c7i7d5XriZaIS/UMw75a9grxidkPDs/eqvynHIK/cxx0O1/FE
84/koqNF5aPbIVHzK49Go7xOCqvOK0aKZhQ5RdDneeqtuUJNnsaLQMOL2PFrMcjj5J+g9aFlvM42
Kxb5uI45Jkd6XkhSw0keFXeGV014UmOLsf9hEL9kbL1nRHfCdu8jzP2Fz2mVqAqBLYj7RahMhEJ2
3JdxWErW2H6Pb3CoST8ZtXzb1X4mr1czCsBSI989ZWXpnWtcrhFpoevhHQSzqN4ssK6ynYZuwF65
HPGsSj8pmiDrvURohAyY/rrZe1DDVPuoIKjOa37FWBeP6qOqLsAI2/XwOn9hXhNTEyYpbVy/9CXn
fJlUpIG9EwL26cN7X80Lb3fXySyRkrS20ekdRiXyPVN4rRVNRQx3c1JI3R9HSpeo+qu1FvWw4Dis
QGFJypIYZC1ESzbrI5a1xRR0ROS78ekdLoKgoPzMSvly86U4HqzkxAJY1yAJbqj+kMU/KC3xd+iV
oC5W3/AGyrIxqiJ6UYuOUOinLPQTFd88PpaVZZTLks07IaeXYIKiKvFBNlGo81cbmgqdgJw1NSFG
hL7fLouHmTISOtsbtgsF2qZFD98K1lL8Ybh84dVaDntgVdsB0LQaI4Uls7d//sroEk09wtY2dv6g
n1ir056CsHoGOnchcEGnUJ1NSGtrj8ddLv7jTqwEXOxUbL+aTlvGrjqixYOmNbS0uWFN9pgNjP4g
ptfRWwQEu29K1whvZ0owXvGsRYob0mlZCBPCakWGpObkM2HiIWlYIS2lY+RMuN6KEFX4vjKyO2W9
gyLXMQNL/ySTVf50nJZgYUj6iQ8oqtWE1ALuvAQm1Etr8iFmGZ2QHFwQuAPbFfK3Iw+/fXI71ry9
ApST6E4kMnfgtJyG9vRO3+mzJ4vshM3y/RnO9/iv5W4EGtKUrEzfASZJreRHWqSL2qmJpbFW+afs
gs3bYl65hZ0pghGP/lIrNrof+o6S3GN8ovuWgCmIV5gU4ZytvXQ/ynrNjGLwtQHdt77fG/UAlJpD
LbtpGaOFtO0MuDQkjt9VQNonLHb8vKVKCMbSv3g5WW5AuRrJqBTTLZt1hM8oaEx5Zpzp/gIK7UCG
iUau/8inDpz//hJ5Ns33PaycrqdR3NdShUKsmBqOSG5gk/jSLfaFX1OIAIztnE2huk5nsT4D2d5K
Va0XoIncHKZ6VC+SQ9CamHkkM74Ksmo0LNgzkwVNwjw6hLcpUiH6Hv0RkUd8fPQF+i6VU87I+HUR
sc1f66aglMddS3n0ANqIHWmem+dIzMBByDraMCtnFdEXa6I0+QI/V9ArnN08l4mzQgBefGd6Kg/v
UtMDnh5W2bFE2zzjWa31q9pr99fbeN+MciR7l+8B2c72Ht1La1uftRRvbTh/aOVK2YuK4I3X609p
OnP2Wyi1jDgFeabVlHPqzsea7OnomQJtE1dOS0CNhMaGJdFiQ68E7IsCn56WjfPFWud6/lZRPaxP
xI7O8G+Q7LrgtMvjHN9yHBeQFa1SsohwW/DZTILPbixmJWPgFE0dTt0T4RMCT4NPQW8kxDzkoK4D
Ac0Gm8p/TlAfDMSDh6JQkmjEXJci5PAR3aAXUSauTucsGyfoRakHgB83AVvHyDdrhF+MW1rPsF5d
luhBi1UcLBF7SiQiVBpaQMOGGbXB4CvyyabxSNBxVrqzEBoEOZs+D8yW9JXgdMfD0Gyd1S/DfdPi
i4CTldlrbDr9s2t3iyI+bwFYodDQUjs65Ua2Ui2nwpmiK9XMQMkM/UY9dCw5kAFAPZv6SadeNvLb
niOMtI7Ii9BUTru2sxSC3bVT3YEjkIf2plKPWgw4KIVT5UwuhYnB7GxHExvtkPu4Oa6WhQWkToZi
u9nK+2vW8dcVvnNz73ogC218Z/0t+q0lCyrStXmuiO3ryUpCBoVHecFSZdgJlzO+COoz8jL9Qj4C
obZDbYuPCXcq5UZZ16EMqphKDrCt5qFcuYxya0/OZgI5Ng4TD45FHcjPtVasq21ZYWko7OpnFclw
pDA84wWU/bbQ5K7GDafVS/Q/FW79izXud2VzyFHheml/uVIfmNABgxocSLyAzegpfFrdHcsRCN0K
ZaB0ctgwtc+4fiopMY+tj70hHB2aMLh2TsUZZajqYxbl0hLAjdU3VjvzmRxfo3dAdTlHFGjAo5Ns
ioA5jk8KNhZOiP2wVXx3mGW/+oGKO8OBGVny6YN84xay/RhXU/EGyEQ6KwAeGB8PCQJVeYnwnsm3
WkITmFnm3X4bpaYtCPQ471J/Tm8P0V9QeE9HjQxtHN3tBfb5GXa2eoFvcCZL36xS4EuWKvS8EmRt
fHZWakFiKdh3mmPwaUL6jpBY/jbI7Jf/+kjjwWQNrgN/SskMUMvJQtJRXkKq0/8+ekE72Hwq2mNZ
RqoMlTnST85VTP6nAjKftZIiis+X/yFN03J8jy2Lq5yNmhQRgOjXPRb4O0DcRTiDRZ4xo09cPkNS
Xs3EIBVPM9ueRZ6I890lFEDxJI+Ls0rwEXcZB0Q9EOXiuMiwm26J5sZeaMwJbF6bS+YkOj6C2Pnv
SThd5W8JzzHregyYJa10p0J/Y6cGcInCl1shH/T+Wbe2r8s/Wl7l4qau4IAofgaShiTL0kGfr5d6
kSHnv7rKOQJ6lGuCclN95xfhsj/OsRQbCk73nAVJ+J+0KxYyh61j6reBcc3LO3EQOV7o1jjc63iu
fwRTg0W0o7uGRhe6Z8QBb9UtIRaZhB966w2+LD2i+GZuiCMsAyJ+NK0BZifk+3OyyfcVDEClzFNI
bmNA3/vznFLZQBJ0b7UZCRyQ7wPaDOQVuyevDVWp1N4nufyTj6EY16A3rNPnlq8KctGTE7mxyHnx
4qirW2PO2U82AnOP9lWY7TeIzWo5emn7BHxcjbIoifjR9Ioyr6csSjg/0VBcbG0Ym35j019896vs
oEz7M9KagQb6Wb+wm0oGkmMQo70EzCIqtMH8zK7LYcTZSDw41Se5RCEfDnGceh7V8RdX5jsE+ghV
YlB1ySVpGSIEwA1ydrNesIac2iN6A3ffxXkMuqr1yWnXY8te0PaTN3O1YeSdQw/O+TLtyoFTD3E/
DG95tHgLSVN981Pc1OmaWwtgEpy40KLRRlAUFQsfKk9E127t5cMZVHhxpPp639KR3+wPyh2kV9g6
k3MbXFznyeHZtnbk6bBtgkKf5CHhyHFkj57Ak1gSXAzKTw36HKw7463FEtnCoOWE44qQ6TxoVmwT
Hdu5XBrzNEJmEksoGfgaeBiAk/ORmPFNRD6ZpVWVctn2JuWdCw46AolKjkhmUBeoOkWWi9vxKwDd
VgPBRNFeHXUc65I2su2tDbmII7BlShPoATz1ZUazK+OopqT3dP6k3Rf5Dm1iZgVKBkejzE+S46gB
nFM80WUuXoTBAffjys91BMdEDzl35WZ6rYKm9pHbtgMS4wLsCY9rGx5TEFZSRSexN5R2VzEDfpSS
g5rCGh3dQztFJvNTFHz1ODOHA0vFkXhC6i0vfgap/2g7+jAHA7y+7yw85PtkGDIeKXa3S0Byv7aG
DpPgwU012Vra9gKyVRX0K6AGMWJWFfRUXj1eECrsxfLpskAm3eTlvsyfm8UN0IIaJ9/mOj6FCg4i
4OjIw3c0t4s1axZUIeWL3tkgshUIQjNyMLC5fPIyd5SPmC3ioXvU49woBwojS5M5ANn+51rQGKoh
wA44OdMjw1JPnJog8aGRzYxvpm1dJ3yKF+Ae6BNddjO0hAB54NwRKJrUOTQ9GtaueFwIjA02z1mj
IEaoeXbSerbIFD7LWzYizS5vrC3zmWhfXoD5t7rW+LfbVqgJDXd1OKS16uqwW/LYK9Kjb7SclykI
uZ5kr8cJkJ0OQI2gKtWw+Vi9ChnjbA+mk8zuv+RtWmYP/5FaCTBd4VVu8/rSJ+SlNUR+nK2nTDOD
pmym/RMIwTbSuOrdinV71L+f78D6spovy0d2Dumg8knfu4VJT/yy8ZsbLQO6EldWRkFUZtNKCBTR
AlsLCuyDrn1wL6pALisKSgrf2oVAIAg2Hf9YMGxp7kX8vb8yQuqcRkMbxp0Xw7eCxr6Bwufhaym2
KR60hLijfEJ+oIX5Pj/aGuqCiITVlZt3yQGh74FE/5387CtVONjXIxl2kTXjwA/pYYRxdOzV0422
oZMUUCL8+PuWu2HCa2wwA/EZE3WLwwTv6SPxfXuO7u35ZUAaDJTnwBD34o8psX2oiGf+HhAnwBXM
C3uSBfYPZxrFbl14vlImLuxjHgBIHyoFmmZQr5eO/7TY18rQh8gD/N4UIz3sZ2ciRVFIRdgCylzL
ARDdk3VSt1BjvEj9LBIE/9IMFLQ6wuXQFL9ilVv5DqTQOBEnXs+zSQZiVLqYRa+1koRZn6h31ZsQ
Bzk9c5VyWSe6JxENVOtULL+nbi2Ddc5uoj0CKzufFRsaO7Wc9pNhNlDuAqtPflLgzYvK3zjE40IB
ipyr1jUaOt5Mr83j6PIfqOuFBvzNxas3+m/s4meNGwgJdK+8hEnkHdMg3gqdpN7zQ3iBhEweL1sN
ghoiHWQ90t3bSgPhKonaSnBH7CgD3TjE4TNxeSeWrh/lleNmIwlRShS8oTBJkoWKs4GfdluLpPhY
DQSxL4OWEesQ8RMj2ZQAGsAMQxAhggn7f9glVXNyLot9Gy+D3YQYsd1wcNf0hSwoozXsMhsXRO04
q/2ZjQEjMOIJpMOpUy7tkbbNRf/6/2i+WU9YMEvj9VzoaNmyrt1d/Hjfuoi1Tsr3JYlIzr4wK2w4
1UzxPynvk2wN6b2gh3WPsluAl/SvqjRO7yk0UWIhE6RzKvfEhvqXjNYPt9aPU/n1lBucf1j/vT8Y
1cvKdJ0Ip8eMCMX5nv7Z69Bm6uiAbdKR5SFbFCYuKY3JO3l7SSXkx+gEMyLlzAsPZoOIiwvrHgOo
Q68WZ4nwZbVMGWJtob9R+IBNDbbbW7QErs2nU5Q2v63Fb6VDxT1qtGX/HsTUl9StG8mcLR0oFDgC
ynDm8FZPuyywc8NUIceeBhELOLqH8TlVGpGzGRkpbp8p/ab9RSrm5dVYcfeZWx8o9UKnlG6YoMea
Hn93PWi7M+T9pE/XOnC/QWkxQMJ3IUB2ZuFwFh3Rhx6+1QOg/B+HEZ+wnVeLPRVj9mjpVHmeXjhe
uKw5PoCrWk3PCPBvaEL6OVqZsrJLbCKs8Q4fLWajhm33nyDj2OAtaIcrhUfUbQaR+xhuPgTOK4z9
BSJu+GMQo2vy5NdCBFG+gN3pjylsZ3vAaMNv4CAjdKnRnTsSMa2CKqUvi+gZo7Hcbwzr2rKw5ZON
EMvOoKif6Hq8A4TZLFZdit5KsXzfyDU0bO4R9ZtW/qi19P77XB2DZKYAqO/IjezPaVB1AU0EGq26
JzO0ZU8q9l77kiWfXsBsM+hvJ8mqMesdQArr6zaLRiHAxnAYpHgosGMcUP2cZHCIB92UPd8FwgNt
sDuaDupdbWF5Yu3GSmXmXJAwcX18JhWrnWaIdAIVVRIGuvFCe4fkp811jY83AfqI6+96kxSTHFr+
aeTAVlVLlHc/b+C9GlXUvDJ1ve4+9uqM4Ydb7rYzmFLo7WmGQbvvt7gJzadlJ3ouXJKY6Pw1aLm3
wjln+H2yn5DiFhMawQ+4lMkyqZeOMnE8ortxasA1zyef1FSge+2O8Q8EW5Sq8JqstpXRp619eR3v
LYsZHDrjLyn7j8jbzfcbEhT2J6G+TTJWdx8qobHi8V9FnA2LK2ICXYUOaoJgIQCjwXAFfspJq62+
ZodAaystAU1BcFbeJr0Pyar8uclF4wyhyfISrxIye2bWUZReJ7BB8bYptPd0GJQjp83BsNId79fo
MTEZBsYHK2xmQLF0JA6OrRFtAS8JOlrv+cqpiOIL/L0RBcRVKFIu7iW9krZf4oVqtqtc/hSkLxBo
scExazgWFuTk1nj4ekHJwTDANsTICRSTUc5ozoHfGlB1D3rfrhUGgQQdf/9Ad4EoZVMR5xorygj1
ZSoitvZw6DsbzsHoOo9k+5zFcq3MXjhH/e1h2ZA/NOMhD4j9kN4JQcn/gmHyEESDtXE58lu9LxCi
pMcaUmRpfbdV7nphWq8YbyZJTs2Woin5Nh80cmubnlzRqHjvWi+bScmbtXdJnTaJpYGNuvks/AA2
RZHTNv4P/fOoSALhddZJlNGDfhPxCeFam8OvIgOO1Z8My+LOyKXsI+AjYDnPHM3yLNshgVn8q0Fo
wQ3DryQFxzphH0C8J41Umifms92m4fv2M4TX9w48npd/+xQvNFNrlbim1KFUBLTWPeeU+PjDqj8F
DoyjUgpDfIQ8CU7H5m8UG/5jfvTH4I5/zPJPGldfp/HdD2NCMX/X5+ICN2DxDhJ/jWze1Kzavg1C
MMnooR9pKrhnJS4qh8JNczW8SWaxTII0nmifjrXWm7RZ7jBF1126yRhCUkVHfkYHZEjW0SKpMUdt
irIYArnvGLztDCXjvLVlaaeKyquh5s9sOh+XmRcHU06cpDWJ/Jwme/i94HbrgvmqJBZcSr+YeWX+
LqnBV0a6sk52AsTgWiLN2qvKr4Rdc5DidMoLRbMphJhlyp+hxK0e8Q0rOvRCz5eGVV1SAo1fz2r1
E1iI8jCL1CnTAq4DuOF6TRRlQceemG4fIp4STKU68qrEaHe41ZeOb9MYrHCsoWWMUSeHpTuLsY2/
+glSlIV5Mk3sppS1evzT1RvQLglPXP025Gwfi1uDQdO3+bm1LEc6TYeo21GoIgvMWvH3gj8wd/fr
If9O9DJTBsHx/s9fRPgh4wL13HYYJg4ZiI7eR47ujBwnTNACeKHRxtlQKN47d4Gz3QRv38NK7tuN
lurFCGxtV0Rgco4TYAiPP9CGuUvF11LRWKSAQmIrG5nuJ/l85018tUPxW2w2rNoyHQRSWPPp860o
bXLWjddhDygO7hZjw//FRXfsvI4LEuHeQ6x9FUAqoFnp37XeOIMLZ0o3tvl3dhVldKr+X/0zaqa7
oQIflgO1KgsRTNQTlyJ52WtK8RtGZjoB9Kq7+9U0HA+M9RvVj83jHdhKn7ehFiOyIV18ewBgl5hu
nF95BtHSsZLrdI4POWmVPD029Kurgz+sUCIoYdUp3aB6R2Txe77L20lFxg9QCzG+OylwohZUsYh0
ivy4H78yWTewWKrRIII2Pm5XmE4mQyu4/HqYWwmsNP40He3xoBqainJTmW4+pK3GBkqxHKMesxO6
4E55054Gvf79owurQqCjYBYy1Stt9cqZF7pk7wRXoPeJ3mFHpdWMMFvApySDa2pDAp4Z8CmNqHvn
XmVu19Sw1PcUOHowNa867dNik36bnHoDuq5zbHYcsVTs2jfMKqGB025KUsXccRLO/y8fuyWG8I8b
zp0qyyWLrkTDAa11pJIo+c2ebA5S73dsAC9KkSlIAnhwMONokY8WJzA5/udreV7RduDapxX54GSW
jgcJej+xiSQbQTfvsuaKqMRQsi+KnrSBukwP0Z+AtN0A8ikMNIEYOFeCrXySiX+QHIza8TT7xoqa
5AH0Bw0AewKapGcAi0z5ImJk/GwLhiSviUSoH1B4HgFe2TheQVfELxiHbycORYh81tCb9mEVAkqD
QqW0w/gysKOu7P3tXV/D/PSQShnOsRSmd/nER8vD4WYWcSAMlNGsu+x1X7h7HyPcNdnVPWV9CETQ
ItX4197q9pkjFQuA5UDGNzDBRJjpCx2fr2RzhiW/P11lTK90zhJ41XZTO67Wd0jh5JMjMsNyshaa
jFP2yMdwTV7AsoCThDZEn/saZxyqZj4VsPkTXe3SMz3MmAXjV+Gi6DoVGg8OQmzD+z5a4ehQxB4G
6Fa07Ui+SB3YR058PiRguea4HDWF43LMp9fkuRrVLK8MU43TYlY3pLhEzC+npWMcf3axAUJyLU6g
361OTUpeT6zWj3WbfIIuN+11JqSRg6rFKnPnMvxwTlcd5NAIQNsvOliWiZZmpguUKmPuXfa35SoM
ovn1RXSrZqKgv+N2l/36ps6HhyfgimXpyVKVqKGbtTFNXD3Euacoj/x3Zg5lq+rYMTBCSUyxNexE
fRxVy1ZdMfnYw/p5bYbEU6zr8GTeYVdxIBNg9KdMViP2DY/7fUbEochk4ID56855nNgeMa3HlSMm
Lz/KMb0Kwhu1v8xRiBnzu10yRhqByb/+V3b9MK5mhETlXbS9C6LPIdPliP0CoVoMFAaDKOa0kpLy
06fmL9Z00NtHhVj2NWNBr6KsF/OxS18kJgpS/kZlv3JAjNkMht9NHaIW/PiDYLD5gPGuwuR79uVf
u0Yyd51LCMW+dgA9YYWOZvFDgBfR0EfOtYEHriwN5DyuIGk3dEA9foADQeAA6ukD3d0T3TUk1wIq
WxnSuF1HisrVuUt/bFsV6MbEqs9S1o0laKyvFJdh7JtQ9a5DIjI6i3O3hGuDlHIJ8A0M7ggNrAnI
Fr7X0kqL29c7iDjnm3ZcEcFt4uzgCpfPkOUcCJMD/230CRIDV/Pj8kFjC21SPdnKe/deEb2kzdZU
srclCiMDQrXgSU78Ys4yrHwVWlYHCaetCPegokAPDoxQ3uBDyqpyU4ubgpTkNcOqRgzAS1rsLumb
DsDyy98srPanYCtKOW1V41aooxQqpbulv7tUBREyw84ew3ZvkG4DejU0JbvKZGZ5Y8JyJPizBbgb
ZtYYrSM5pcjt1MUC4XpVHEq5U8UGKP4ZVv4mddS5Isd4cpWy7VsPvTpixa7qf5WuTMHt3YBX17Sz
6EJ1y/4RH3U9gbYPDKgQnl2pT0M0w1Un23TT1GGQyQK4bmrwSIR8WQnnqskiUx7r5Ht7Fb7imqjk
vZ3tjjoUrKLRHYPvbdeSrsyc4PWEi20r2UtIGqynieUVrUnaBGeDtS9dga7aeJsWYCCogpQGwko2
9TWOdIMs1gs6fBLuM/69w8HQvzpdTdQOKERbao99Aai8gcqGryO1MwgPXeJ9Gb5aYfE5wt895VNo
bpogLlnOjk4rJmE42ptejJeVXtWBu3ZoI3gdCtfDkLlmBBIFXEtgXnHi79gthmdkDRmr+mOKv6UU
gjxSW3Lp5zLj/vNytw+4aaj+RrE9S6bSJWC8uMor5st5uOP5/6j3dD1H+mnrUMZHXgIFZOkytmlB
1ANfpg5469GMhLxcQKuDh5VF7GWVeOpNFQCqs7SjluHf7yWc5123cdlYMv6qAHQU6bCiyaCq7YWy
paC+sO1sHoD7Ls1kDyLEolCoJWdQEPJ58Cj0QbcUROwi0J+NJjqVH1Ygm99bMrvGY6xTmnVaJR/T
TjQUCxJAIZkozPGLrCIvmLLDTOyS7VlnI/MeJfok2JSM9SvGwVsellHRybd9FowbOuKDVdN+rqn9
t89IJ6dd7Nvf/4uq2zW9EaxLWeQ3tHXEJdM7jO8Y+hbD9kVnpEbNi5vGaoeIp6Vt0p26Cmv1oc8x
Gn6XVpyHC8DzjTZB6S99ldWVO/xhuYx8SEQlsDgqRbk73o+VqOYZOwouV/GtgAapBxG39TQPr0/V
eWOmp6JgQQl2rRsy9A3smQh42LrvuweTVmuneKR9f45cZLzN0MbhSH8hx+aMfxr8Uu2YR2RjNZo7
IIGIXW5/D8MjHnVmaVSsECxPaFDOq1/MT/DhsltDr6pEqWlppkzvm4AXEvPkNC1FKlUv7MW3WWTx
URxWuwx0vjlVCeGXnB5Ob/fNGbQ6jKx+egNKeIEdiREhRpPbFJP63CT8n/iJK40tXSh0zZnIo9Q3
T2RdkqKrI8K91IwszHFpSViFmCLee+KicdrrW5jyFEo1OoWjI1YRQPqd22zFF3cJtuSu6oZegot2
dH9aiASG3WOfnvzAiMjY9BrUeKeyG0wdH3UR33FUnCe+r8ARo3O70DA7eq/N60eHdXXdgoDnbWWJ
uEq/RQuSW1i1mzleNNxIiYf+HJjxwhLImS0tT5EXDdnrzk813FRhtYzcm/n7Zf8sfq0q/qviooRz
Zc5tLzMtNZlZDAGavVyI7AruCpWa911T8ktJwZvEC+LFYuaDEnjis6KbFLRHwXNGT7lnsevoqfcR
NJ7Qs+S94dli/kG74TUpSJFVHMSOHky9/uzCI+RAAZlQh+iFoUwU60qF+RFmbc9YjffW8dk1e4t0
rXbJM3vEfBS9FdA0MMUXmRpcgJkPKuiAay602XgsKNd7tWIKUSnCwsHUhM4UHDx6wBsDRVdMkN49
YI23l2qx2fJO3oJtcMOTRQXX1onxGqWPlB0MRwTtgnvUQWkuzA0RNNS6uFUAizxcaZNq2UHL581/
Qc4ivLvHdaxmcCpFSQeqDRS8hwNHnGtrXS8wFGvWfo9D9dI1pBBVEsta0HU4y9U4RKaR32RYQWDm
ePCWANVPDGGJf04XOPPg/CoWzl/pX/F771QjTPipV1RhmvgXQ+kLS/GySFkxBXzOSNiCt+BG8fbM
vSEm1JSShJuTIV2d/2WpNKiPdCUrQp8zNP0ceWCPPue5xlXPenOgi3QZECMojPyZgVR3t5K/FmmS
LZvrz2fMnl4YZemmABuweQUH9f6Wbp/X8jrMAeQuXFgfYSkwV9xLorlgT3oJ0a7J7t7XqZW+xvmJ
UV6sbLVDEsz+1yZ3Rp7dgcsHyle+LXblw4sttS9+s8ADQ1hZOIAtM5lduWN414pxVOuOpg7kRJdK
FEWcTFYLTQSal1dbIhcMSvOw4Y4Q3k6JjCqa4g6W8fxkuZeoxd08lwNmW0JXppoj7w3rUSnKhM7B
ZWp63SPjTaYu2AQpJkjNdoEZ1tS6xMotuqB0yEVVjjk0qGa6H4zjMiJaYn4LEz4l8Na2IVbctRzT
n3tKTVFgjChB9XF7z2N4YyJCiV5/qAbO9kRG4fmEMn2O/SQu8MfLZwZVqQpa3/B/wCz+Y8XFW4tj
HiuGMpSjUMtx1kSm/g8qZ/WOa3VvrCpVnIWAbSknx89QZ+NGUJwIcfjNnqs8ws+cu+uhWH1BL4hV
spUCG6AxIGwacKuQqiHD3zG+HgigZRtuExmfJ/DX+UhHmgEHoR81MyipekYB3LbhuEVT7WlFFkwH
OPbtJTxMhXU3hHt0bGIkukM9e4xHwh12BqocswwzUC8Y+Pvqxhl1eW7F8NRRL2mBWrFB88qBhoZy
D/ttPQ+vEGU1RPrycy0aTMTZ52MWUxuxmxSWXzyz7mYtcM8b4ZkZqN8jqkBrYdUfS2TQts/EUlAU
iaVEjomWHRY85bRVSoxfcW4lO/ZxQHIVCPBX6Bo3JcALYhaUhRHsPax4NKC2Gd/dOtitPywIRNdw
Dgp3Y/cA7HvhQiWq3rgucAtdomBcJRF7Wf4W9pnpMveVnr/AAQp0E9EpUu8rTsaREgcnLIaSF9rW
+wyGx74w5cfOeakQLLMiPKyyBfbTpCgd+xcc0LAfzdKpUqUogC+WwhSP37zw3ezUa28TTFfm72HL
mytvk1ZcdYpB4ruz0bAEUFxG3QYtesrZD6ZsPyv4mpU6FCYlsIzh0jlNK991lXH651I543TbGSrJ
QjdZIEUnuN/W0GRCl+33a6y8l8UesH5nKETRW9SMO27SEPB0Gf+ISQyI9j6CuMOq8JvT8vsL52Zo
B05KZQSjN6HPqtGaYYrYgTF0dsJ85bSK0GWuQhyBpnvifF26KJ87MnWlWS0JEex5bRqEWB/MOadx
vM9NzSNGQvMxD6jGTvsHvUNrOV7+UGD84ejFHuyX5qwmo6LkNPRBO1BXuEnHhMUWnCh0QxqwA4ie
mBRehnTGuvonQ1WV8GxZQzFs++bPA2AHlRrlt2pmMow7boPgqQ/FVBDZZftpm6TRKR8r0PV062gd
o8oRBqMXxiqoqSZFavcRH/laENNeTm+W7TWhIyl5rOjfpmcFNS+ADCVn1FRXM/UOr6q4Hqx+TUUK
SbE0AeDRiQamzFgUxrJ/zwcZnRNZi+p0/HAVdZKelojkiPbLLaoXi0TpHoSxuWetp4dLytHmY/mU
rYs5wyd7jI9h6Vb7m1PIgZnyGefpbeJ5if6j+PVAOKGDMQJEfSEVflbeXaFtILSY1esDSOzq2ECy
f2qnH0J9HxSjiwfRmGzeWn30Hc+QE++uTX5yT6eHBQhBspjm/EVubgGiZiJXtYJX+RY77iQ2VaqH
DpzTkneVyY75PoX0PVTq4bDdYhVgTvMZZrKboYAUrfXu4zV+XvvhnsOyQtehn23OFyODs9nIDaTG
IaDfNC2bCgRL+mvwX3K7YXAN/nYfxfosCGTAPw8jJeJ8mpW4XCrb37XMNtQR5/xrrHBNxTnTbhaV
FaDnflufpOid2ihhmiWLN4Syw4zgnJS5dNQhO+VR7X2QvRHWe6vGhfNiqdXaofsOIf4sETbsSX25
ckHiOOZwH8S1kWcchzyw58SHiHBZaZbEDcB21Y9UO0EMhtKy2oFlQYzA7yaly50bEaJnqOfj5VAp
bq/ox34tSA0wIoQ0hTsGNNCOdzhPLYFVw9AhmMuJXiSUONuhHLCqORMzFfkskyFPA7g6mjZ1ZBGb
EXtOCgskujMYsqd8p5dmoqGadMzQukSn7nYzguURslGMenHyazo+m83BlhGtxHAiOip3BY8xdcWb
WRoo4SPq1XGhRf+jAHmcP9tTdPL+YhQB4yM/Fw7sjBes+ahexBw9N7bE3aeX8H2UEVgtkNfj7V0l
OXpi+eZh+Ne35mRgOtXFXPylUntwa6mEgasG8c5slfj/NUJ6a97pNNTAoRKpLpn6UJGx3kbywzgi
riRxJcTvZgmJQwGCN9mOkF54WKqelybCa5xJNAd8qGu6Sf9C7FOlcApTNfcwaB7KIBEvl1Mjx450
MSxCsAl/HhZRcj3P/I/s0urJwLaZcF1hPTxYL//CrY3BWi4rPhy5MqTBvS9PZIUMMaKX/XUzQvhM
gNBSpTDljk1uCAgSIS9vFi0IlRwr+gIjz+XtXWwnN5z3Gz/EGubpBGWtEMq7dhVN/JjUtEc6JdfG
dxnnzwiBO/DH4KqbqciND0O3r2F9iByP/f848TpIOry0qyGKrr6bzj5ruh6oV3sW5XkiTBnnqjcl
VuL1SiXdLNNff6p4A5KbkUyWAFNawdlRB5MT+qIWR3VsxyyfFisLd44nXcGzN0xlvOktuZPEhT59
vlqMQCi2pL2yA1w6ryBnllvJXlnP74vLf3A6Vix3mcw7qMMKZ+j4RWi81oF6+6LOp2km6tF0Jhah
2DcQMVW+dYMbfIysjeiFA183prW/5s7UO1D1LAvZ9cP+POqfhgaBPTFJFjpQOcycU1T7WcLc/k26
ZwVEK5S8UXcpw/E1y6/4Vu6zxgCWKJdPOS0eQsNhWC85wQQf2hUeITzl7mtCnGP/QPipswFj3gw2
imqIRPd08E6T0icTvrO7wItfKQO+jtceaepWt9x1N5r49rm6lfuW+9ZSdDfbHu/24ovxNJyX1rf8
1xG9xSkHUAer/DTyFJuk8A59yNMyaRfFjus7H9UhqY65pgzjcE60oP21+yhNUVzaSJhUJqC8nsd7
1nFDmfTlkrJwzijFGKFIrD31tNcCmvziIgpfzAhq9cJiysnuMkit7Uw3Uo+xbbqrvNL0McnvoDOT
uGTMUGXNV1TC8/qabkQHSh+yLQ7H2YEZZMz4nR65Dvu3vAOv8JEPHel/6GCAWxVPPC+3DbnG78TT
jfFBIRrpf13PS1NkuZLcbpUjN9GqX2e6DK5Jh4xwArk2zZAybitoEpXzycCn10/LjqjgW6wR8Srq
SU3iGSQltJOCwPwFJXd4G5n/mcjQaZLeZjj9252lrTmh2dEg/rns+sSOLGPOEK4UxWie5P/u614z
YUgios3s5uaVtQ/KHWGTn/aFbmHLxMPGBjz2wWgjn7bNbvVqC+VwXgIVuLwaavWifyVFVbjYxNL2
lh/EC3CNyKswEtlbRwtDk297+rt9uZXssiXI9gZDGz7iy/72tMGctL0HxE4/6bkV9l4YmlKUo/lR
1+L6flCyeNjeu+j/nCg6OgfD/3Wul5bzTtYOLtaVhsbmQwn95fbNviZCislNXFdxMLyROC4v/6Cm
rOBu7LM7+cOCfdwrQOTQ4sLrgyTCZ1I0J7ZbaiQgQC9fJq1aOplhDkzzQn6cG8RoABvH3k9kbFP6
u4dE74pOsHkkcjYIgbk46nRNZtvrPkmA3ZVV220vyHmZK8VakY2QKPafolxpklOjItwEDxes9EN6
I/HB+QWfftocn7+oaFExm+QrvtvgQx7/r5QoQqsl06Wzlp6BkBxAriqwGowhJCCukTGY3+MTf/pH
N+sJ3g2RGQmybl7i9z+hz/rEOKoE01u4qdDqOZyXOcCU3EzA/VQzbVSxkx71tdVpbVcqNFDne4ec
YbbBLeNvvzsw5f8CGTtI/IlJ2P+/qV51zhURjFC5ZiAO5vpBiJQ1hGPbnq0C+q31C0e7wRNvLJyC
g99Xa6bUsxA47yjhZ1aw/SFqWpzhBAtPys4Q02igMzVa7zzV51YGmcqsTuBAMtfZ/KIsst4L25vC
OaXe4yeiPQ9ICJltXflDFVpF4Be3bonqOUmlLi3SXc8fR2jGGpRJn+hZsk6LmYhLgTGRvCWCIP/D
t83Yls84Wb+58BZ9huxwZX2jYOxVMHvea6OUg9xo9ooU/yiIoa6CLYb/u3TqUzZvv4VyrXb6L2uM
rgWAwyhaXqdJyRzCLfCXG1bbZR0VV5aKCUYZLTTV0oeJlYRTyDBlBsTCKU7G7a9QjsGX/MzeKVUp
2UkUWeU59Lp3dWZVv1QxVZ8PuCBxZNdlKawnHiPS+al6g/jlnN9CBHbcbUay4Tr0qfMypNFUWe4H
JdfiVacbibWIAg6ORTFkSlEduoRGXzGlFjSUsNKUP4CX1RF6jUkxknvclwUGM/pjggPWMSHQRUtb
8urIwvB+RxxZbv9xPsV0ZFvPTkH2K6aJ9CVvjFRf1jnQ87c2q65ImZrVLvPuN18ceOtz2uO6P5LQ
XmrL7/0j5yRBQ31TNLaLPiWC9bT7CZtjLhCMy1NNwBHmmbzVgoOoKij75RTSJfdqLASLuYYsAjdN
Jpi8eciumoQ+A0cLtZ/pRxdPBqiWPivYreUOJOBhNeGEhctJ+NSLpsaeWy8WfG/EL+38SN6xSu1U
ub3/i7My2kNKFMBHr7boNiud+dKtLq3Wx+zbvLIJlLnGd7HaefrtMR9uQ1a5WkZCkKvhP7fksqHW
iE6A2MuTszG91MIBhPjEYp8zkJ37ek26FVIO0hNWkjr7vuBGHzL/iF5ZY6WkZw+20aqGfmDVktJJ
KncAU/OpsyGLPIGFDg0CBYICimnebN5xItne03Z3LNvO9ABjK6nUmBuv0bx95/HtMQpFF0lCUXA4
duHmtbU37oZQfmBz1AIMpm80Rog3ssiQ5RsJR7wJ0wVWcEsISFZWFdpne9/J8JS09p+GzjQ0+Xfz
+N0yHQrzoZCzAZSRjYrqKS7CQ0//9lpWqBX2OQXEw8U9k0QuQ8LXOoFLVhPIpfHdDLoFEg3hkjQD
U6T1GnIr/EPJEz8VyPKk34DSYi/gnMKmUJeMJyyGVib8a9PwQ+0S3YUE/Fzs7A3hIVqQuYgwFHs9
2ktiKtNWPfrE0tJLPGrRcmnfUHPu0ZVBydwzMky/SK/03hd3yu5ePVZiUj7mHVAJFmOCfDXbrWYp
40jszYvF6k7VffX+V3iyp9pu//tJgV8JUKx45TIMlD0gOSU0aQRUnOu2F6loem6Fr6OMVssMgsrs
zitNd8PmzhqYH1PoINXjVuxel0NiDejYVaWFIxmSCxhJtHHmKyrS4p94vjO05Zdcd7DYq5oyuQ1P
cqk14ujUt3F5yXQkcIXQeg2d1PisvVCAU9Ih/HyqRXhZk/SKxSMH6drPojMKRUH6wLqzlr2UUbPm
tvZE3CSiI8ECClZQR3QabEfAjTSX6QOskejqmn1S+4JjS9EVYb+XDjHQ7JAFvNCJqc8x2yAXCmdk
UgizkABsj5IQ5eIJ4tdj5/QG/CODOMBYKuhbXx9Sr0H8smLOWwQBJS2xSYBq9w+PM9maq00xLVp1
u/0WNyw8YX3pDLrGU1HM4mUhxROMTOFkpqacKxJkFV2kkM7B+t8ZUKiEldVwM4eK830yzH3kmKur
kiYHo4FpAnrminzPSdzSysv2hYUH5OlwRyDeZuQauUG5wubvhnhiB/Brug6nS3QFL67DgkT/umsc
HuQnI5aC/yzD5Tv5m7ysKw0ihxCc5LfR894CElIS8BDQh2YRHVQK6uI6kBhacvutW0hXTw00G04U
vYoY61nX/sGpChfkmC/bRcwTV8nwo92f/XmSFDdba5x7R/wbMqtIyXvCRF2CcwgY8SM0ixaZUNl7
KC9aPGWr/WAn0LjxPh1QjAED9w1QKLGUEJ1IndBhmt/fG6TnX0/t4HqPhLCJluvNPvFZT+nV/1Uh
VUQvg51Nksg2KK/n3a8RMLmyicHwTzCOyIpE5WqimHTbxSdiADQc5V15BYLw0H2nb2JVcD78zRnE
KadqK2BfqFJzgc66U4O5RXWZDgjRSjm0kWaaef6S9Kdog4otE47oOcDqrwLI3a30CY/t/5xSe+HM
6bzGwZSlOvfCxXeNrKzlnpmBMFf4bp9NXxyrzb3dAFyavpk7mpxBPVgQVc/V3JFDRRgrj6x/kwro
dzUP9ELJSP2GOAY4PODT83qgBbBnrzNg8IkXQyDgubaJiDOferANz3CiXI/FJ3jokPChjzyddtsr
+fkR3ka6mVG9LnHfimR4YcqrdL94LnGVZbmD2ViVrAOUYMYedmRuU6sMk3E/f/2hEPSxSLF08YdP
2qHV/7/DU+P4Se8rVCkxsD77kIUcJMZ8sh2AOpByIrChLlpVa9Dy4YQIa1EDn/Cr5lrHNDsiEDHA
97CawUkYLmoXUb4gIU/jruWZw0ECYUN7gi9SDe/FHhoDm3roN9C2iwmz77J3GH4UY/cIVFRGKBSr
8SOSUWIRy1i65j6EwhvqJRolMDoOXvpc5dSEs0Z3/HJIW3Slx4TRHIe1uxIO4jg/6+hwy7SXXoOq
/D7xazXBbT34sKJja9fwA82yMLAWQD46KN9oLngp9EeRhJF/H6mEr+5Qpucw/UQcghv766c5qRfl
y0ntXgtEp7+iGZhsxwrGxfI+bBSEa81284ZCNNpWj+8OfKuCKqAZZPk6ziVsKhJwVPPfPNRUNOH3
lwAb0stSoV0AKV0pIJykjAnfpq6E4O+AgqgmPaUZQcjQ1r/O0n3psfwspdOh6CsHj7iyWoxqsGgi
FmHVSOE1KypTyVNSW0Mwgct4d0tXXy92Rr/OQyqpjXScMEpYSXkeGfq7lqj4tSf99Qvrqlg8bIdQ
rzrFCUtd2LcannbjajLYISJFDjhJBJD3WDolLOsvlmQEbyoTJpuXETPwuORAEH+qQYiuxeyu0ldl
RZRK8d4xEN7ZNQMaPnvXZT9NGjiiiiL6wN3BfTFsah4iG+H5Z6p+OxXyA1A7elyyt7V1qCTSSYuz
3l/qHwanj+0TueYMD7aO3M6P4kUdX6UPJL4KsU6rtgkBhZjmki+ATSLIPph6oXz9V5CsTfzUBpWm
oecQFRMHdKTBXSZXnKfOEFY5NDC2jMNAXDo9o4ygh2lh0P1Nphcyz4f08juf2/RJsEFGIDsxlIEE
L/sJHRG99jX2I0yBqlaA0Hdtf8hWDm/g34UNkDyMCcsPVOT9akVqSl9mbwIBQrL6B6xI+qp5dsYx
LHHo7dr501mT8BDrB/jTE3XpUg18hyQjGBMYBzZyaMdmkYgHlTJ+Mm85aqcNmqVCPCILrZeQwLYh
2gE2rY41Lg6EcSEnsBAJ7i67nBlZ7LOSYevlEoELYF2WbRJOT78AaGm8MrlluXu9pi3xmXI6q06v
2lIS0rnehnn4YYPCujoHvNmSQIQs25j+kEknOniTW3qHqJ6Otq3rvZJzVKotrWXIKt70TyVf1KYa
RwwAR/10QbpeOTq++iJMiSEBVCE9kSs2P1rPmE5sKU9rd140kSwhD6QmUXmag6Dw1CMJQDc2+kyM
ExdFv9ww70C2MNgWBO6Xcj2r47KVQ7oIZ0MdFyyLCXJ5RJkQ2MA2p4lKr08UF4pzBv2Q2OUeoGXV
Q5qWyMd4fwrd6kwGg/iz1aav3ESiYp+JihPmZrknKJ/wNhFezR/xRFsmC1w5a09px7pRzXC8eDgs
STUERGzKPn21kwex4zq891zQGaaU5oRebxb9oQuBNPv5ZYKRjJ8Gu0d2TB04xiroj75lX+XBawA1
k+Uu7rphFvfzFkpKYKfOk6A4E4jFdzFMzw9ll3AzzbFF6S9CHOYHnqaZbGfA0DVomG2u7IuzjU//
tbjDEmnFHadWcfWEeWVT0SKmYdC1Qb+qet9GlIR48ZAF2cCY8ZKwTF0oRg8Gp/LVb0Jaor8Xsfuu
BFAnPESmEuL3MS1dT4uCXlPmUxBU07DFALhjeNahr9gIV1SOs4+yotkqcVq5nziOR0CpxGoXX4aG
AV5RJ0LTB0jqWaVok/kU/Ex0edGXZfbyNvnbJcgQdzSlgDmGwBZiUftbtT/PKvh952gopf2FSl1y
QFeT4xayPRr9BzDf3gPORFAb/5WGlZ5YqCCUVE2eVdswy4eiZVJw8m0E8o3bUvS1EJU1fSONlObL
y3d6q209S50fSUhVPIqpsr0JNRdiiDk0Au6dXmNPI4kc2fDRdHViW0dFGoPdaKYQe2g3wiJqAzJD
qngkdfv9ek6EzW3/00SKAJAoD37DE5EWSsfRnx6AyMyhMd48F1QNDP/xu8d1jWGLkjzVgMTLNACA
5AUhyfwqykEmGvIjhso2LWlrImXKr46RqHaEayDLOzoVuZlV3nbgBpS042gjHFd/DdR/aksbu616
oYx4swAf01U/DELRj6Yt/B8Zg4dzpYzaKav8mLTtD5QUwy5Yh00y9z9EGP3tUkbrD/6rKScZPtUq
j02H1C4ifuOW4XWFQI93j6sw9VXnb5Ke1VZT6iGgG1dUmCzOZwLJuaNQJilCKVk83tq2eylA0b5u
4FN52Htp7IJK1XDuavWv57F0GSuuEOY5hkIlvCjvVEWLGPiDKccAS2LngVtkStLxBs5sazayq9I/
aHJLVOs1eBtKhov27JJhPYCvIux+pLMRtmunWbXxxM4YGKvxL63pbkmbj8CuliXoh1/p3wpf+4GG
WuTGqCjFXcGdLqaxCUB/9Ue9u6n/smGR1OadHeubJyNcsmqkWrlV62xAfbSnAr86mB8ovHr/kLMp
1m0FPdSrCnciYjrcdylqsAT+sg8wX05g45JDjFOlWjegGRJyowEEqO42pJYsafpqQQCtMf/O0L5S
cK5//nI72/aCFUQvZu+q3y4MqJJKFBuZ2ndLSt65ManMhza5ha9xsUzpX4wIAiMXbc0goDu4rew8
DzEJlqMKf/ZLxaHvovrIOYJnRv+SdttQnHLkrB02iOjAV6h27BMALDbt8NGcsXBcxFbCfcRSvJLr
2WGUpp8CmzLE3mdG9xOYsSjzgpAIO4ki277Yuu6wD3A8/rOSQO32NwwkgSehviQqFbbFflTLN1CP
+jWSLL1xUl4jPUlZwvpAAJg9HAwNqhdWlYQ2gZ1SW1YmcfzY4FEppZa+TwSe4dwPdKq+8sKnzESV
ovnGfRg/PhFbHQdYhDCuLRLTdRR4wWlySZLo9qvpf/Yjtw4lkBo+Hlw1PJ3e9pvK1DzcmYXsnMlp
yLE++ohLK0Qa6i7V8phYw2KrQQCN0kVjNewZLhcmptdJz7jL8aPRnsvgo7gKwMvCzY+USJNBNtyN
MyLWTNfsVfGuYnAk15Ct+KrKVOZw9MM6xRvuSH0cjsaWdy13GDU6ZWlvLNw4hzh4Mxh2hpXkDk4x
DLXz6+JNBl6lx9R1j+QD+LLuWxwiQQlBOobvynTjADTU4E28JSa+lCmMd2dvuZWi2VcKy4A+ANxX
tsg6TjYW9QG3W4VV1ayM1eS65XCJO95Yni6iF3NSnufCpTQDtuCFZ1I5rBensXbO4gjZjy/7DXAp
u7tEtS0B7gcHSLX9GazYJjSZ0LhX1eftmESU3F/IdRIc4jeigFhpMAxd1RJwaVdsKrok2PJmr2QV
vBt/pufTElQLn6ynepXon5wmT1kOQNKlugj+wCk6Ifu6qtpKoAUjQ2+99/80UrXrjzUcC7kDi5tS
IlczsgX0pjaDDa4iUHIyml+18KrqIpciux2O9o9mbOqVKhAnVPwgaCAaWEVnmYv3V3gsN6xYsZlW
IORTR13DydmfHkyLpmiQ1i9CdZpWyUbcyTyt4gX+sJK4qxdnXH5+lPuAQZvg0Bieyc3eGqqgovIT
j3FaqsAIrjBbck7sd/gB5tyfvEDOji9NXF4v+3fqYL8K8VtXMw9gFi12a8AcOu6Dvt8ugVqneZ95
PJVqKjDjHFhLfwphEH6TCWS7Go0Lp2AASBd2TIK6H8QCdwhh9wf+UP+5BaESyImqq9wXxMEb3/X+
BVJDWyPEd2ED1v1oSSU6G3/Ar1ewRWH2Ecenh8vhvfL3f+gRyHnekLvydXEx+X3jk0odidoffxnE
5LZ8hZX5ntFX7LzEF13zksU9K/yUBpEzVeHy31RoxKZ4LjmhJNAKM8gGWVv3jFGlwXlJxQANIXrh
UOdhNI7cgAxnANSBxW3bDKF/zxoe3t1u95zbtEXmUwPAeSqbaNcOqj1cws/3/RV1uj5geR0DHBr/
9+AP2t4EV+szVtHhpAOFSq3C3Q6mO+arbejLKn2Yp+72mDvqU3eSQm6th09jR943tqXtViri05Ga
LdLzqAvceapDDN5arvjLNcRDTYdopQlB2fy3ChV6CihnY4aX1bToP+1LC6QKpEjGjY4OCXWsxmV9
s+jWRiUzdjwEn/tb4tCjvbtS9nqGAE0pKqI9b5VyvzYv/+Ysqc5xjFlEAfwkl3t6eOstY7R2irvs
Ob4dWu6fXbTaTCXNapo1vJae8J1RzaezJCNdcn9qCI4NFB4lxq4uOl7C5/Nn+T6vwY6Ador3seYr
m09EzONL2YZhGEFYVJwnJs+KvCqXGrmJdCRYO4YMpUVZqQxl25iOV1EndRqMzPK5PzBDnU5HbPlk
VcGjR8bmu4TVQ2phdYwVwrE6UwzuxUszVqOaTUmbwSdB3W58nUHCZ8YMeEvvj3dzv7aBjt1wWhz+
a4xMDT7L6F70pk3losluHSWbpqLljVY4W6vhzt4jhs6kWBQ5I1eDUt2/HDPrTinlnQI1jqcdLxWq
BNkSnpRlb1MykIPzReepJdZbke7cGO7XPz451sX4C8PN7ErK4Yyhkw0mDtjURp428UYoOZldqUwF
4xosol57BABVIqQZfZp4BFXL+D6f967sqG5LlHJspeuQSc60PB985BGVCsD5yimfhZTh6nC8s9Pr
al/X4wOdHie16+UfzDesXzlkFXb/C3u6ozkR5skASIe/fD0pNRr8ZfVtUfRfIvdqgDTnNG8OCREn
C3pIx4DB1sg2BZtkvhorDzSOiDSaOLo6Hk2s+4UIyGhK+8yZRzQe1mm9P+u1D2ifsVLaH/aA4Ig9
aomYxyTj5DTvOWRX/QgGQq5afrqn+txAWO3izrqxppZlrMua14Rdr4dDpYbbDhvJYwnWNyR1+0CX
q6vyMVW8d+jk8dSR8vlYnqj7ZSN486HczPUr4VaG7d4TqpMtZ6tUZCe2CsZlQdcaaCH2W6NMCqn2
KNC5Lzcse68WteSNiUyKYIUr/A8mx0nO6CCTZG3neD7TPZEttUpmzkT+LnKx9/Lx8kpyhZwSp2KV
nNUhct5eCYxRKkelbW5rwQVghwn6c1ucR0ON6l6aRq/PpnZ5mBUAHlkEYk7iaexqSq1512zkvIkO
tWco04+NjGVAoAG20v1/oDSM/JPveImQlRfDUhoW730AwqsnGRKeimCrMC7IG7b7hPsina4xx9uj
MYzdfs55pmAEbo7owLkLEy5Anb+1u6z8eqUaXkhJqSfjcywMJQMdzZgWYMedapTIvZJED3wm7CyT
WkGM1SMOZeFSJb+5365zQ87wcdqzIWqxBdKfXogCPQXGLpCuioz9UFRT+ATrEeLf48a9SpZVBNUU
oY8K2KH9Hmww6cC3GV58bz6D2kZX39uy9Imm0qJcQdJIgpmMIiZ1KpawXjPa6Bqpxv4228EZbRDa
0mxGLRjeGDItWOQLosgPq3QxZobV4hY+uXLrDL2qZOkDuBlw6j6BYoXrj6j2tzBOrEVKNukC7Gjn
ygwKCUreaNgE6Hhdl68K/IREO9Y0R2exTGFJ8CtT2zc5+1izRVrFuOpuUx4MzTR++RD1hxZaQj6A
nQABbueB7ZgmS0mAvX4tYPneuT0kcvGADD01IQVbqLZNC9/aE/wO7JoIkOgt3nW6Q44VreBsk88M
VneI0j0/qwCIp8wtsVfMuvCS37xegmAF9LFGtf2RzcMTdQlD+CxgeJxdTF2tSgb87SoBiDLeXWgj
wVRvXKpup2C6LZAhUfroo2n09d+ECrlThdtWm6Bcugp3GSa8CJyDIel8A/toFSOCJhwpIPsP4k2j
b3I1pmVufy/3YWsJTlf2W1uKN8RqZF4ccEaaw783jYjQyC47WunWH+HWf2GKlwVZt7zXGue0d9Zl
nwIfO+F2D5JShtja9SDHC9yLWs3NWF46aPXweUxMO6pfv50SNSI2Yvjmlh82Kyyx3bfvVoo+SkXY
HabaBGhon790m04d7MS6nMY1oCy/OkTGix2aMaQVH/tb0HCZH6Yxu9TN9QaUalwnoHmxZafbFGgz
pieEliG6dWpfjIYVTmMN7l9iXyZo9NEeYZ6q57zjeFCi5u2jTqIZ+9fnDqKnAubIn0+HEn8lxANo
ntjCjyapODQGosBYgNJvhza4OgLRkYL3gWiuU5CsEdOzUCdKK34HdR7OaP26tBEzBwmV3quPXdK9
D4uhae00HAxjGT1zq8sJqtUsTm7OsjYTuXLXW9gDp75krt7qxAPenps3yXr9jKlBzq7FPc02+G2V
atqxJQuJNdZifpRLltmTlebOIYpkEWho8lv69K+qL5CUzC41l7e+Kj5Dh7Hlqdjeb7NeCi5Ep74/
+N3QYs3oB0iDxAhkkwo/pkmkWc94jFXyaV20OEzS4d11MbDpcAPwlO5QFYadENfEsMcyEmrf6W9I
RQbtIm0jXjXOdiC0DX9TO7XTVL5j6QOItfLW6xRDTmYiVnxJlUYpbFy77SJItrXmMDpT7ukSElYq
7qkcM9BgSCBAOz33lDH5/hSYKRlWUXXzunjkMfG5tI2NWJlcbjtZWFPPRPZ0jcXb76P3u63D3RL7
cO5uKGEdUntdNs+4bUgvlmqLaNrXJZdOBwFygnjXdt3aeQoexMQwv9h94oLzNNwD7cFqO7SI/VxH
uzF3keoDNrN2pvlfbwhJzCQzqEav2ZzKjzm3SwWwt4n+2tEWY30KEWYYoFE7F6bXEPGatHKKuL+g
7KSuxflUNcdkVAmTOnMIjngXiYQQOfC/+bpnhMWISslp76JrFNLci53dsPe1GUm2do7o5IZwmw5V
RxkrQOgKoYAoFRKlL/qY3N7gXSw8c0blAX+aqkeV/oonfclkY2EOQ7I9Dpusl7xo+wAO+eMVJ624
ouGFHNrg9UEcIp1wxFFdzewTYGpJKgSnyty8Rg4TMs2OJ1K1pzicDXns3ZrMgQEIyB7gNu/FPdKX
iw4BppryvoKcdF+ixyF8FmW5nkJyJkXxWmIEJpHINavLDRBIdp1NcjuJiJVw5b5RqKvK6B/pxr11
oiETD6wqFRoqScXlrWeInTpwkKR4u+HrAaWO3MYARfScdlQ7YsHFTXJ/eehmDPqTtXABWX+TNaDX
LRsgF09HofRkoBT2pm7nsMa/36IK2sv9ECIZ85HCGPTBceCUOv6R5Wy0WosUwldQvRQj49zTUszV
nNNK5wcdcVcS3Kaq0KoO6OghaGhIiHWdnOtASyjxoNIEtjXcPA7xODjzxRfZnZ3MbFml0mjR0a3d
q2zJ3EV4x+2OCzperqdHMFxegbkfqvOmFG7O1nFOauVwkekGrUqc4dzN+0icHlxB7QfsKJRkRAXk
AfTUeXheJZq3kMhNQwpjN6mFe8qux5LqZSGZHpcvWjXExCXyupMTAH/DzSiPfu49meyP+680eV0w
RMIJBx98s8lBbs1oQr9D1VX0HrpUdZR43UiPL8SY4QI/ohNd1jZ05BjIDx0loNaP/T/kTqaiJ3+Y
diE9PoQDypUgiwE4VsggtEmWLMalteRDOp0m8poJbsDCdmwG1bMhWMdw/GU/HLIWRK2sKvtbi2HP
7nJ0gQl4OH/n422pkyicdo7HiqKzPEocysnoNBbzMOE3AtXr3Q+uhq+4IPWUqHlwqWTlQfb+Nzbf
bQg2GBFqBygJ4tRb5NN4FHFzf2cgqGnuTdWUQNi4Dr9+Ic7oJp/oopb/t+Dz+QznNeBunOaBDY17
rWpdJ+wlIk4rBmqjO+wumT52CcbbLVAJBXcmAm0x6+N3BE3BfEIusoZ8X2skXD4cIHvv7gsH5dr1
REOrN5t8dRdJ1i4bfT9akCA+QTBMURTs0cwgOxxubJ8a2FqbTpwnbSHZz8FYha/rGu3q5OEGEOzL
8EzP7PQcVKvGJcMBiZQrBeDz9eoyuh5t/UNtN2LqPvbGKwrHi29rWsLv8ZtADeclOrZXoyTGesMg
vZIxcQvJO+6jDMJRVsqiQHBTqEsI6+DNYVtbo47qCjBU7otLKk2gqrst2NWa18qH9V27uirXoy3u
PuYgZ9Oh6Vkk6w6mZSaIFyBmjaaZz1siyFnrYmPdBEoHb4+oGKEgmphCCLHXnjy1iZr3fN+4gBGh
Uk6/CiMVRCu0FG4YbtrhA8LqIAJuYwTbQIcd9faX5j2TZ9u6uWZUYoDZO25JG87eSYFJuAT9xykj
99xoe3jv6Yn3gu0bnS/Zd8l/LJpzK7q2w/hu4FHdPmcHC2yY+2KnjtUOet6PxgBciRtams6HPQmX
dutk12vPlS4WXV4UnGvcs0Sou9t2UjlvVMZqL3IAuC2Ma+Sqp9RnH0PqEMFebT3dgPXEza16VjA6
F4cZ+w6Y4Hl+0sEQRnhhWjVDdB6cxAiohKpDiAY3v9m0ZHV1+UM6ZjrKrCbRJVKWwrrsjNasNLvJ
sw0uA7AE3n1VbL3yLNomjLiM6dG3rPS1EHKlzmCAAgBUuZ4nmFavImkVkt8f95+9OoTmHg0QbEC1
kvoFAaD8qYB9h8FXvJko0h2/M7T+gE0S97/fNRo7T+Pn5/rUmE2GzZSMks/WegToX9Yc+0WiXXGk
xo2C5fCwMCjpp0YqQ+EhKOphrmMu26WOKL29JrLadq3dQuQHRgKPXlmS0CBtRu6vS7k19GbrD0OY
d5ClMtv5Lf0MdvCsPf9nxEyXcLJvdDiVvoV+evOE4cDVgEBkX39Nn99F8bmTWCXCgKOr2fnSD+fB
NdOkM71G/qjjxleRIp81vbCmVZz7HjY2RPdNZtxzLlvCmuubnI2NABRd347EcixmnLyUCf0vqsVx
WIbe31S1WiuG8fMWIqsMB5SjJz1WmC0G+NcUqcLB+xvxfayP+h+ANkds/E7Ulk6bGTHDBnNYdTF+
NgQVC4UARZy1sC0CEQaEJWL9Ce/mlOyIO4RY0agxK1cAwURjSwGfNMbL1gIq90fqYE2hf8KKbTWb
m9z6quvu63sCPAOisaFcSgqjL8Lh+PAS2bgt7KT8czjhqlBfhuxQdOqxpAFXSdB9bnrEpDBwrsrs
r+MF9atz304sD6EUXf6OVVTTL2VVYTlJz1nA8I54IRJeNeo6twtt0+NuDa0oQQw1HRQrt7fQB+53
3onubDN25OctgbHNefSiINd+7dYgpz0uW2dFobANBN9YW+NfHb31aWMnQWnCOLlexmthyURdvG5t
SXYy8wA0dZBMmpZvBK2H+CL/fmcL1IStyzuaHpDr737gD/tVxivMssd/fpZrFwI+75vBZZB2yDlZ
pPiNKn641BXmx8CJ+rJyPn9T1lPYOvLY2c1nx5B7HcIxliDkoNbCOy6povuI6EGcbljEis6wWNRn
J8WO6dDLZ/pSlm9twyG5NPBfq2trDOTX4chcmJWFKxFr/FXW6mvEQ/rf38UF4ofuWH4NRZjw8iKI
32qqvJCql+SQTXLS1XKo/NeZb7Dgmz3Y7q/N2Lgrs23qqV+LvrNNlN8TGMj0r8argLT+37qCGXc2
9RzaJLUp8qJDWQHBLCd5K6+gK5AAD9OmXfeyV2OI66Fu9N+RkT9DP/avK5ozUhYr1AP52QgDjp4M
fG4xIEa8nSfD5xD55EARY13/QOXgqSpuqPGTm8tMXbO/GcST6fpPIWB8J/PG7lqnc0570MmiTIDq
ckCBPfUtu3S9GoPYwXqhaEUz8HjiuxbMufraNGMANFMlPz9CHMRa9X8yRajMrrQRHs3HYGmRFS1X
Ym65aiQjRsjMFHu8CtyLkc0frQWYFsmtcGULEuIuu+OvlTehNclwC5zsr+VXZu8vrtItTy+iQCY7
iV8DQzfRGcxrQDY26t9pTUuwmR+glvI12Fi9QWN4e+fpd1EGuKL9/D1nUScq9FB1v8DzZIJch5U3
SudKRgtjakMQ4RgwuqdF5n6B4z0muPtSreESEJGF8HZVISQYiiUoVjbtekXCHYlpYmVUhtvt6sPz
r91g47RwCkqjz8z9nJyuXeZ28sDKlPuKzy2vrm3Yv0/BwoUuBo1UfHoEKesObz3WRSa8X9t/Kkmn
8B9ON3rKQpS0Z41PHyaV2DZe/qb3bQrUy4lioJOLLVwhp0bs3CYW7RD0+GrTZx/WESldhRMdIuAj
z3dcJCvJYRizejQnwcwSIOlXYqoM1CaQdLZBxx19qJg9JLoA/4n/+qVsNSkSkj2HsWSE20plBOcA
Sq4Twf/22ZzTN1xHTliaH2GF3RhCkKgEcVabejd6lbl2n6CXFXyI9K26Ju5w8GjiIs8SGf0CVGY7
NyMOnLpp49rfx5QnNZ5DDCQStuRUjsv3HkH4+LSBjvZH/Qk2l4YoO3TnoFHONrNhvp5bsfy4j4bR
qK1zlrvd2nOAgR0CG//3Xy+Xd3S3/ryPJL9QyH9BXdYBfzZycYmUCAXko3BiDknHi9HQsFXTLp99
YxzF1TKHyAZG8pR0jJYzbxUyFiwaSkSeYLRy29e7+6WAObtE9ZVTv58nRa9H8J6BDAdnbzHcQ+7m
j0jtttZwOEJwWCqv6cS6w8k77fNMWu3Z6Ce/EVJ669XTOTqADJOnD8cb0MmDFxpNJY2W73IdCx7J
TEgJhgC5pt0lH8NxUsbD5rYm5DyI29vtsUepJnwN4tIko0ZQhrQQjE0gep9gI1J5zL0o9hhagzPh
BWVh1LM6pAYtEttZgwrhyeT8u09kbWn37gGg7l9EMot6MdE4AUSOPcbcK6xhm0vD+ZuLI2edYiSz
7h4uPLvLf7Jc1I+fwhP1OMwtAeidRhUWNSqIkP0W5bqnSkT+s4MvWpXSGEuiBJDsvWdRwrwtRdWN
mcIPe+6rGT6gFowsc2vKXhnXOtwcOKtXEPouz1HfKznjaTzhNKRGilI62KeAv45Inu6xmFk+Y1so
4e8IIesUZ5mdR1qYbjVy8nujlFh7RLxlkVxQngf1BVS9ND9+1qtMLRt1w6DHrV7N82hu0Z6pqd7V
5yLjxCCaRgIELAQK4rM57A+ufaXfgfy1de5o/Am1E0wpCprcPaEXk2ZfBLss9hLh97rK63KioQAQ
lVttH0W/Q8HVdg+hcOvI4Cgp8vbcmxcvuyl83Q3N7uzpQ9ZeLdpfaGyNho82g+AKmOQfOOs017t3
HG/IyBVksFmew4w4KpNHS5AsaJTO9QIK7EA0xD5O43il0MZ86AxCPop3ItJRLvSZQp3MNiM1Yw9p
JdvKWMBNj04z65lIFONmoI3Nj7W7FNtDLE/QpjHZ/7FBH7s6XayDVfET2deyEBCV9pLm0BRpygru
F+ruGnsd3UhvZTY/co1sPIjh21xUWxhnTXZK8Anapw9eDO/eUx88wVmzn8ABZnJWBrNI7VyeBqeo
jv/ntPgCPxEdrfiT4yUfxlO3w1+JD+aXUwigXtgl+GvxKSVgy3r12RWveM5mFmTAZ9tOkT/jKq6N
yGSctMiWWsqwf/U51kSZjr17f4zrWq0PZbyNRvktKdt/3ez+bfAyLLbEMlnIhWqYFutHCZqtOpSI
pjOWDAashTUiLbUZM5bVP5OW2XLiBg6EuDyj3VcDlf8BcyYHhV7n80uAkxwe5IEh5vuztu0w6F1a
erHZUw6A9AnupSKEZDrn0d6WwxRGl6/7z6Mzb3kfdRNG0v+3L0SKcQK3U+TmtuAHqDftLhCmtZ2D
UFBN4b7yIccmYBj7HmuN65Rt0xRnIJ77PoBvC28vSOkZG0m8xljAAU5E9bZUPuMPDT7M8TAdRmeB
7XgGrTBScVzfLBXnC3r83D0OXDwJuiClPcsGV1Odu3pIFBmiD7z0jlCRCrmsnUvBFLJfRE3E6DWc
d+W75Szv+pElY9k52/02MAWtOh0R7HNEeZFo17IEr77NSihsOUSW72C1/2Nv5DHYfUp2yz2Tg3dj
U3lsTNTbBygCafcnvzZYCRfxSuhePR22NbflrlhANJmo1WIeOIr4NPsFUgyiu6fW4HeFEwuy6FON
h9SULY3VFpa6t73MXfYr53AS0/+8uILpO/SvollPUDf1Xeg+KacJ/9B1K4+oRDH3oHZ/SmhLpg8j
fvZrnlrn1oZvleBCiI54TZ7s7Gh4jJMkpsbFJwv/gkXNeNBhEvFl1w/hLFvXHx9dVa++p82RFwkj
oQPzWquu9FEYyEC+CqoQQNcQjP9ks25aGXbkQ81WmV3ZKPGQVpNh/g3gWpZTe5Ba/UXWR2nSmtqz
5tyYcbdDgftQP3Q0Bebii/XtIJHK98zLJgCY8fpFp5JPVCbp3sTRdKjFZHxUw2AU0s6VHI7uYcBA
gh75mFRO0ANlHZTAktnqPMSGpclgPbTujzlexaIajtfdAHm5/z8C2diTMYQXiiiEC1M6ZrNsTbwh
N6ZyXdSlQkHXmC+9woO5y4Oqeg5yb9iWh2wpEOLSt0lbkVZ2ka+OQLyCPNIDHYMhoBl0OnsSilOq
vFzCLquYG1+5BprMyP+3igfyF5HovyBJkSvFzyKRBTeYPfSFMhcUNTb//OCMhGnx+m/rPKvHZFYQ
BoWN+mhOiKa2T6fmKcVeVLdO6JhDCATX27RAWJLmNOSlQdRhvLnRFionOugsM1Iwf39f/547bOvi
tIy/gNMWsQeD2Vflnaf3Z4DopX5N8fV+n4Lzsr2uWOFG11MP7Qs+VyB59uy7qPleoA/dt5ne/0wG
Y7eXlcemfa8O4vxsclpfJfq1uF7AfFW83hLYY5usER8lj6U3M/rZrdnGy02UVC1+TWIqbRpyc2Bx
Ekfj2oClIoZP5MQwoadA12QnhHE3Rzz0/cmFpb321QoMd0UjnVisLAGiS+ybOq9DHHBFPvqfZINX
L7G3HmofNU2WYOZnFxsxwFU3b5m+jWUtWOk8J/a1EeQZoHaYJ0HNSRHDrKOrBskLIbYS0De5Dl6s
ulsAaUU9+zNFCNqNJVJ6ijBWrDE4Lysl4UPLmV7bRGFs0PYSKJVVKt/rKwIGb+w4tCTpg0Te3lLX
xCv0vnm6Jn1lUO5RwUZZIrBZT14P2Kme36vqcif+PY7Q4nuP5ZXwfPDc+ITAOP6mPttsz/EFhmJq
cQpmkONtUWDyxhBA1aCnLWmcr9MPaWfrJCFdrmg6VIXLppSH1K86TLjy+TmdIgFFuN+FK6TATX5H
eRvCZOkWc1NJ8/EqWmvoorX9rFiJwzYQ4DG+mats6z5fKUeOTvCSqzCfCghEUndp/UjkuRU30nHS
9tg/vlUiaw2XV+IWtqtJ4R4IsODlhQ36WYk01OHIsZ/YP0Z9ZzfHEIGulOqT4DgZQ8Mnl9r48jtD
b5ok1xKdyRXfibqmAbVVMESncGKWeK+Ag4kJjaile35PiE/2PVdgi34bP77PXQ6WaZ+OqhoVuMwc
ofDnoy9MLYAc795Sm6UWW/o+xgzWpUIr6B89YkAIF4NNuVLJCPxhB6ntgKXsXAXrB9l0T8sLfv8M
zoCAkhdJNiw65KQfxw/i8NxmrEeNMwU0B33et7gZETHfV/4lN0xUTn0HLoWG79H86TQbhfc0NZbM
pbc64hyQ4BMNivKTSgW+x6uUQy+DFZKmQ8Xoaeu+9WQa0n+1SRyI1iboD1IDz7OPRRa5FVy4OQ/N
SRw99WzKn0sctZ+9JBS7swYR7J8y9t+JcZLKvnTKD3oVym9IIKSZkiVg+0mBAt1uhH7n1wcio1N0
m99dr+bgG331UYYBgamvR6APs4ClWD8sUgFkD4P2qw9b56DP1K1ar/MyHILj+YMUb81nOiKo5MRu
mIHSWXC9LuzWngCzw5++xiGvrqM56pvFtXcR2BPNVfxtXOKPjsp/JxqeIxbXJUoVPpuTN3bQA+nZ
5gD8eCjRClzfKobz5vabqjTSYUK6MfgM2GFKmh4zSoMo15NVFI//Zr9qhsQ5i2SgbZ9SWlcQLQGY
IBU6Dg6w2S+NOBxVIKVMEnKmZE/l8ZP+ETdrJCzuBHn/53aqnUW37vlIX7TgyAeDMG20z5WutvjS
JbMUfZUX55+V41rv9bW4ONPKc5oQvaZbWG1EfbITCvkPlCuojOAUsJVeqjEOziKmx6cC0YcTE9j2
9pmI0tWDcuZ3bVNnvvZfJ3qAlgGZhpsay+zhU0fylSdhXfp2hiwq7CYi7vZXmJks8o1yLMueR2s4
64QJ6etmQAaXi+xNAtF+XWQ4jLbcQIzBHYmdrKvoSxIbLUDUMwC4ynkAGk1I6FnDXlUBcb3Ev5RJ
Ps5z+MmKI9HdVILahJyjB2Sbzxp9HBEpLvFwObNRcy10vEpKn+ihO8KAnhUuNmzgv2DO/G4C30eS
BXW+ckZlqvmiGc/MX/MIXZYgRoLIz2GBpTZjW/W+rK4EbiVpVO4EODSZRFVdFS30d0M5olaNng4q
JEtkK18AWDXBXBKk4JZMa3mj1M4uuyaO/BlbeJ8RAOwCeHnFDs9V5u8s/bgJAjjKmPJeVW/z6th3
j+P+koF76/YSt1KBWuIiMNpAqmoXVw6mtM9fwHMIBOPQO+Z8FAJRuy53iJJqoMphTGcd1igSqo5E
2x+PoMldYEMEPRtLRZB9R0+n5G4g98ZMSkiYjfNbXXDTDRKavcduTP32UcyujZ0H0FG6m9PCZhNH
NrAwjOdz4Dozf18G/DFL8X8PCtydo2xUfyNcY9YmnuggHm0wi+jP8ZVapSwFqLECuyfgmyy8zKyL
OZbJNDxMI0xD4y0CXIGuThcsSQUycnT5ttTqvOrVUyNu27oWpvf5Xako+uSxNH+tqErCF+1+pB9x
8euqhRVt12Rj9LE0BY+PeOh1bazMeZx6JqZzQ8CQK4IE1io+TmxT5MSe6TkWi27IAcAq1yXE9TR1
WchkwaoL1N5/3EM6dHYC1J/zc8bn/OFiAhh1nhBBTqgmGBbPQeQKO0jlQ2EY9II5B8k1IWk3dvGV
lwRmXw4XsV8rM9LtD5r8pkHNKybFTJDi+SjlnOQWk8rap4ecZJHhnmy2bnCbXfWV95g8chgn1Dto
XSkU3AET35UU4JGOnvUWNJHGmXBygT2OTXlsBxGNlHnxAhqkhcO8SxSYrRX/Cz9HIKwivp3U1M7v
aTo0fBTOsL2EwiUtHBHPLfVNdEVWG32VEBD+OIFcJoUaRX0PzHttdiDgs2y4IU4RT1e/Zr4vYVbA
SG8IknRNWDSoGbu3AxToqchudgmFTmEpTGT3C2cYXEsP+Kd22pu2iSpjq7bAXhRxNJpJUUJ5KwO2
Q33zGjcah+AmW8ALDJ77mRv3Eyf9i2WnZ9yu6ZWFWhL3IQxn+70PzXrWd2dZAvE0j+ZEYAn8mU4l
RJyNVF/6/364Jz/RF7auDUX45Uu/eRlUIwQLaMiwcBf018eHtpLaezMchjPjhthqGXIdYk+wdmLC
VUwRIdvqVf/Oblc5tjr+2oUflU3zSflYn3aBHyRR23wJ+TJfHCa7yuadPyZ47Toel0Rpklwa0xkq
FJR8R+oKnHcwLafltOdHSJ7G6l4F286YLInibiblTh5YjhofGHCC0ir3dEQ+9EBzmdmC4l1hGVZ5
+rKgn/fBmYNaN3oJn4A5lRest86pmew00xIGLLMeah8FboWEsVPtI2y8/oe4SIpjNz+1z98LFIxo
0RsQAKakOA6zktfgb89U7Dkx3njZsFsI2ELNbjFZsjSTakl90ovbddOSOlo8pZ7tzD0bk7sju+GK
K2ysC6qDazeC0NgWgi8xS5fADIVJnkdBRpOc6hp9mOsP5p42KUoy4gnkwic3bvm+uub2VftG4kuS
OUW4ruuJ0cHmWhVxlO/ONW222tOLjIoxqqfq018X89rFmojc8c1gNOOYy5WhYtXiBhTwYAT0hUOw
8sAfApiAN8+FQYebBas6MhH17gm2u+74ShkGUdXLBA1o/RayzLFBnMsVTUX/nQp2yODTFTTS0hUu
tmqOi1WjcZP/uZTf6Y/lF+ghaBRSwo5FCVPcI663iqk/vPAtD8TsjNKdm8aJ8zK6YwwjmJcayyyC
0DMfL1mqswFVTCCXShQmtqa+frnFwUvxfvJuoS8jLxqriL7magfTMHf4GW7kCTJYn0xd5MM7r92V
r5o3YWvuoIYNq7xVCYyKnyqPuAJJZk2Fw+x0I3u2acAgZjSnR378dl1dpec0q33aZalBdNl9FP/4
0aSsdz0Idf1JWAHqj3sIlNNHLPOSUq6Mwp155/SvszfS8ZSeVD6xWrZdOYl4q+dUMm6MfsXRoRqk
cfZdJoYgxsXEjAHo+P5Tt4WpCgr5gjtZ2FNGwLYlBR2bTH+paQuRwZYwF+pPPM6XPnaf1obLLpXX
BKjfG6tQRqSMoN/4LZAG59J25WAjC1k6JPQHwN554WAWrjm46i5vjazFM3xO6fCmx6UinPpoFj3Q
l3mxgyCutAwXo+Pvl4KOwpMzdPFMGljFcRMK34b4IdF92YHdj1JfhsRjIE9dnznsYr6Sizxuujiw
rdkoNIOVWif9RrsLTlJlieQEc4iERh6OLRlHLGJzNahbChQVBPl+IWwQp5LT+K5cuuYfYdLieuur
B9klURe31Yx5yOliiDNXYXWb6SfsisAa8NlIvroqVnz34pE+enXWQ/FxuIUj3v1PivzyZhnelXOz
W6i4hsmES0tB/ctJVljB5r75vPW6wQg8MEubg9dZY85aYEJ16qCVTQ6njG6bhBXS/sdIMaVla+mX
rgFZWhpOMO0voUTCO2/3DUqchvgGpPC0seXThydrce2y3PbcHAwwpfT0+Hjn6EYZ6EexotgnOxcp
9ZBX60p30Pd0LXbLFokxs5VXNKYLSRMB3w78ZI3nCZxX3Cn+jGv/DI+KzuSwVCm6+EJAywhvXCVf
jm2WHr7jzsW8YkXCp5ZwSQ+W3wyMvvy92s640Vj1C6fB+Dg+jMqcuy/gu/KeVH32o5O6oe0rPaS+
m6wwJd3XGwKXUZfMQonoMWTChFTPGP2XC6cvb8aqRBxVaTJLdfJzjgN6IP7Od8AYw+unnlPM4XCn
+Uq0NppwQp5N3q0mOni6t8Fpvj24PrSKhWsdBQxulGYaVr2y8oO5gYZq6eRc2a3iF7aIe7cbQorv
MeOPW4roXscihKsb/kosRfwjApXJEJCT1mPTp7w7aMVmVO5JbI2Cui+pND6jgGp2+FDzhp9/Ftm8
qNSTnNmF2agDkVyWkL6qWqahsiHpelqGpMwIh6nDp6nAxWDXrsUgBGdK0wv/6ILre6gRnCdqXuMS
cDWWBiK2cldtEJ2rfuv7WOe5XNfhSBDsSjx7XNbHmlm5G3NC1RWeNJXtEKy7KJdDvMpEomILeXxy
b9z1fT1tObpxSO4mYH1SFZlEZTrj3hxdHa3VEPqwWHzD0btUbbLpczjPPGHBMdII34Qu8nskS149
TFr49YRSTJHBztRyuedf5OBCOVE77GnITbHT+xf1YPRDFWqSfUjkBi5gm433X4VDBBgc8jAAPu+h
pZXb72DrHmjYdW8II+QD2VlMaqm+FdHwjYFrK1LIkD4MH62FPvFjDIQFvvhnkKAvzv01ZoYmv6a4
XbueyKKsVFdrSYCW/qWgtiGsZ2fF2OJY2kwdx7M4sLxTVSQFFbN9MX2WCSGZifDeTY1lIO8Rhl/F
rikkaDb1w9LqbOtDZ9dvrMLfMb8SSjRFS0PnSm8lAM4XITL+mJgPffjx0uGzxVGj+8OEAuMLL8A2
x1+ipuEcIrM8zG4QbE4XoFrniW337+PjxZKyiflQbFxF6LGJ23AD+SjVUTE9UrjpPoapxjhxipRm
pILLrUdtgSz8hBQ1ID19z7KRzd0xFVsQiVNvg9Ui4MgsNCZpxJcSMsafP3U3z7Ghbliiv8i3ytTw
ol6sK4qbbfM8b1BMGsfI8mD8OV7UWdKiYZ5osyH5DPyiClRaWMMTnBAvkYMWEWbzc3HaeQIz7xNQ
7MqwFNFTj/AWF1qhEzVzB/hBQrSFgCvG61oJW7oFnp4R4PF27W+KZFpYx9k7STA56AXR4V83E96V
F9YZA5+hpGfyEidQFMIBKflGbnC58EX/+qGA8jUpbhhtJ+JUYppcof6GMhVx3cH7oJyMaM/5DRea
0cDsU5pqtm0SWAbXbCemDFNMwERqG4/wH1ir3yY97vPjee49HZT1vGk8jl5ZBKITZH1Mop01/DeT
93S3GIAxo0Xslu/bZ3COD+tuwWyVFaWZlbETjmk1U2osItDTLcyJZ796O7T29ilYtIpxQO6deS9q
liEKPIALmjzDwZKP/17ZuRdcmEaPnlSasHTe1RAA0IJwof51Rl09k8AqOOeGoyOMa/1EGB7rVnaO
utzI3xBm1yfC4crE120aTQ9ySPKkV/qd5KLANS67M0cHmK3pupXh9RmXKF98+ec5R8OSw1fQGWIs
ogaYHINDscMgGRv+YT/085IvG3mfTvdylwj88xdpX8JXsPXpVhTmSglXVHFCHhSM42s409a6Uk/1
45AyxXESkr4v2jnW6UcIYIU7nef9a0MTa4L6nECsCa+XcMsiWynmSohmz8kW8k+m0qMd43FN3UrB
bLl+pNFWOelU5Ghc9iUKQVLiLP88HiCniCsBGwY/FL4hPkSfG8jrcZ7bCqGc44Ye1JIpqANzU8Os
9Xh+eUDFigF5yBvpgEvvATs+L1OH9vh2OFiXAd+NXfsY/ExfreSEefYkJNTtngflfbo5/Ruh+cO+
rAB+6FCIKl/zCR00hNxiL8TNK1EzC8ntO664tWnjLNoz2SM7VDrA2AlICiQALzRIpx/npmcIsnKG
6en0pQsnYXqq9PulKwmJJnF17fDS0r3wU119i8Bg1HR9g37oDIXB/agfkc7B0tdE4Rwc6E1tx/jm
KJgUGhVvJpB2Hc/etdIdsYvk4PjU5wfqwu1gOgy7wYMbgo+buhK2RcRfjQih3AbfFIPO24HDT2CE
3UjUxnovGVbW7ob0ma8FJTPNPMvxPbGsERRT0GUB5F3JizmNV4VXG0ENQC7RGYzzC4ZxpxT9/423
Z42lpq4hT39F1RWqBPhYCQEk6/c+I3RamJ83DGE9J4B5TFKNWRtHgn1SuBwxhpqUVYz4lKn67cKF
XjkFtd6zTRE5XllbDJzZ5h6dSL9lE0wAz/5CJso3fG9p4W1KeIr+DngivbZsbAjPWnOp58QhCcnp
t+HjCAqBiLmgSNvzHDo8DRJdYCYVB9fqqmojZ8exFU2EdgPErXrmOM3hxEl2tWtzmTJq42CcTS5c
eTPANrxwKFNO+rejEmTS1sYBg6DvKrwCa5sEnxXDSdHkJ6XTQxdb0OVme06Py/d1NvLunKf3DY1T
aHv/szidE5Lx+0I1pwg+fq7S61F9RE6F85Qz0PBVCeqe8UfDZTVp8+fPd5d30VSZBwAF8AZDMsn8
i4a+0FPw37/JQan2CgkmkUZietXAskwJxyqS/rZfGiJH4cWdx9Epzu2WUX7744MqeiBXbotBBvv0
cGfJodyful0gIXpBe223T7YCwaaKZhAuWMN7+PTUXOcx5lAfAmjpwyP98kr6IwTkp8buk6JBsct2
JjIVlkUE0ejCap3Dh2ShuXbKJLsCJfecQ2tNeD0990OlFSnLQMc58IXQi6Ats4bjVkB4U1t5PaII
cYSGvLq/KoH9MP2ao3f4NhgmY1WIWWc2cLv9kQED6+L/qKf9dA7uGanhlmBoboh84prScNIbLPI4
Mzr7qnsKc5nZNayZGfLoRUDCtF+3rD18Rgow/qFaBk/VAgi7wzu9CXE8lT0u65ylj2XzMY50YX2k
e8LzozprYjeMRl9+Fxf/lXHo6fA+FdEMzaMQ7PFZi1sDOkfcbzhUOGS7yoFXgn0CEUjPYRraB3sx
FyJI2I2lwgrnIUvfZiT/eNq7ah+uookVju56+iy/ZPwAGjftah6GAd5vBDg+PoOmPAdHgm4gnxYx
lVbowQSgvDkI8IeW/RT2U6KIKsf07Z3fQx+EPXfxf2lGca+o6kU7LqFI2BYlO4OAYao+8umMZCFW
cjDVVFn9hUn/Ai4zrc57Daq8mjzhuwEgxI+5nKAp7pNB0B2EbdrGpZ+prxDZUALm2Pxi7+eyhuj3
XsQ+Ieaa9QTjzioV4EUSAmyBvUxRE/xPqr+5i+yki4qWV7zYxjEkSP0xBxL64dh5QJbgWZ7ipJFN
H84Vp5UAL4VKkLobNAj5xmt4pfmRjFMQWhuGH/rJx/WxOjfTFvQuE2tpXZb+UdWoFL9HIsLzOMZz
tsqageX4iemHFWmmHQZhWFxJzzV2BuMVdLpZGBsf941mv84kkWhjqV0KwFEYM9MRN3EvvWdKHOf6
wkzoSdulgAvD2sEEO8pppJe+04yiUK4Uy35ku7g09ZLaqpVgFlp/nN68aN0mXxUAlYqvE8x7tXVW
4aphVUNu1hBiUKAGv5IJxywF6uO/WSRVFXrvhViQlRrpoo+yyhvparA67WpRs5otYt8jypsJKKI4
0MH4tDqSE7FLZnOiogjJlavh70FGzG+FSgAHysARXGNdkvbutouLbsg7yE3TScxsvO1vV8dtufHh
LvjpdVCeVFZHSJyQaugdCPrDeW1ZcMlg+MDLTTVJ+rYxJjs9AabZrBKSLMkal2t8ZsIlIxyCffDD
UePqpwu4RM1PNpJMwGKze/QCitA5kCL1PUkSK7ShAicwIGRpIqD+CE68NUWy34oHGq32iXVoLMSO
VKVDxuxQN5uloW+0f/3k1iWUvvt8T6+CJLImENzI5bBWsm0HMl7Jmw5u75oNq+pNMyKblA8gPEG0
qwlUn3He8LlXF4MDHc4YcR0xBBw09ZgGlRK2q+8l1lRYeHAX0hHEmf3CJQBThIWPfzS8Ua6U+WnG
lIvViiy281For3R+XUWl5QxFNvpLKV/SPib83HMFBgHfVsOQoBwQjV9zJmSaYXhU2K3aKIQnKecd
A0f2lJt5qFgUlOZ+Wl/NU062vhHbeIx43fAZmeosTgxnRA+CJhgtnO4G1D47/8XcfppNBeGHGw4x
NPEEEwLoY9TeNcOqtMrTh70OD18THIjSTuYkNmRJGfKxtbhvwMTYcjSKxrGqaYwumVKHKmd8te+f
p5pdPjVRwCJYKcrHzVnTFWQvEmYY06sdulC+zix4E6IHw2NFAdfNPTfBniAEcFgqgYECO2hV5VmM
W1VrVcpt+slaZbClyozE1EMgQiU9QpQBs2tec7SMX829/w4nYU8UlXUpNyGKt94iTkVg8/wmlrh0
CrXTtYBrNDN0cxKsDA9IBjgo24k9n+LgshHNjjDiVe6mhffu1Bwkh5RQXhuaFC8a5DF8UcuqXPOb
kAsvnYM/+zRje8iRGfAso69PSB7dF8BRb/MKLBHEDHpo76RjWsFKSzey6LqHb4KMW/OgWIsqHF/v
L3lWnRCPcC3nv67Pczk8FU0CgYQ5nbJVTOcmeT3dkEx5e3BFY4CyVHgheQQmV3gHEDOat9N3dTyO
2ZIOB0pZvYfzMPiMB9iV7LmyRaJZVoimL9rpzH/cXd5O8/joiuaYzE+YYmQqLoeMPWaaTFuyyBo/
o9DXzHKK1uUIuRMk7FzlbM7HGxTMX45AvTmyTSsWmuRl7Zxlo7AHlv+RhkwFJGD4wy31wpt8FltC
xW/tQNJ4IuTPcGVWbwMrvQ9TjeT7Cqux9IIOoDT56znLbCzq6G9vfYzjovyvV8OYWpRFbw7cLQuu
p4mj4sXEqqIb4G8IHi6B4aRlL3Dqt3TcIJVRTNOZOAj7/ye1Lqu86w1J9yNTp5uS52BnN5J9GiHS
BlscqeyEezZhlszbBxGwud3HwTT6O2uCt7GztSRJTYMZpi4wPE+hkPoVisWqxZx+9MAZNs456QxI
1GXWX0FvgJ+RfBpcXgV+F5dKeytJWqfDXXkPJhjq/EdKVT1SVosqCVs+MZCrmnklIsFA12sxFhTH
mV88dJsv2IYe/KuKj8s1QnGTK8W8isn20XOIBX5lI5wfyXghEbku6Wyz+qrPw3YNWNwLMUg9fXt1
DmLqjEk+tpgZpg55RnYPL7tCTmyImQc2tO7m7HM36gpdD6f+ZDU1wpy+mY4fub3gdQy+F40zdrGa
8gdKYGEaqPOw4bBGWNgJOhqBzrQfpe+qrXJRJJ/iqcfH6Sp2WsMLlsQqrNcGHk08n7dWVbPtrrJn
pnONLtOtyvfZIiP4AFeeuooUaIG1I0piFyV9veJYqouCfL6tCdiGkFyzzivD/PlmOFYikoGTaasZ
sIroXRAgixaDX4wnokEaoZguHQp3SjNSh0BK08wE7ZKBBL/NC3p2KrVwW9cALnhwUQpYNTLxgkGO
lCvoDE44MJs1m7gmqpdIfCM3Yq57ONTYYuVpJsgOM9soU26Sx7Zp9gQizpI1tAwQPiXk2AIJNUCO
/W40Qz3FZUhLYEAzsSQ7eFQakWboMBEbwIAgtDbwpdy+vUVllJnH0XgfUesXH2A4j3dUJwByb43N
bA5e0LBHPodbpXOBy7UFLRy7tQ/iLAjqSHplm8BWk88WfYwtPhGaJGHaA3lzxGnEia9fFBsp0ZqH
mrIJ83NtwYUtjzTgVWJb2IHijfW8za1duMV6Pd+GA4yxYlHt+gQpKPnWi2ofljQUqfXoGBAQLbFU
TN1+KpcdHS0xj1V7Fd8LaoAaP/TLmxgKJ+8JFpTM0wroNeKEszez7b+knupICAfHyf11BZdGoEgK
AQrAZ3wfYKf31wXJhJoN9xPM+2eLLRlXaeoEaHRDNV3IpWfEzzLXCrovz2WUgVCQvwprVd4OF66v
PzOoeBmbTujefFy8mPYRrvXlPRJqWIvzwVVNeX2mTcE/B0lFmm/kXtyKaRnrfrpbxWqMvBdUyMTk
ZHIHakfPGO0qaArrZOTrOzIr5n5vd+1CIRcAd7TBhpdNc2Y/ZWNObPkr1LJHvRoTNRi46d0VN4ei
3KzC2t9c8hegQ9QtUszGxg/OoR/CffX/kNPwPqSSQD/cyMNCprpM+wYV7L2hSQUCBbvlkS8qUxIF
GyrdV7bQWCmFiyqr/VZNmagoYLJL0a0qrO8nR+bArbNPobsm6IiZ3lc/mfrcdzEx2b801DigAnhG
IfsZlzyer2LID6gGZJ+33vZSusEBH8Fkoh9oTBoi1CpOd1kh4Ml96vOEFzG80nit4WOJixEftUe9
YPrQodbPX7OVZXHpWvd6VWqr5y76k1aIQSRIJY3UMsEQ/YISahq3EK5oJzEgl//G2k7xkGYPtdcx
jANxZL++VYryfyxyr6D0eYFvrM6hElDhKjgBFWjPSyVJlxFETedTgJvOwr/W2J5IEqKzpNttz6T4
GSCVb90D8ghXYBhgE+VKuzlzvlIky2WPouwTy6rTv2ESxgFmLdqSmHqqlw6/Cj7Uozi/qgM4KZGt
HNep5KeTNw6kGm94vfApTPK3UUrFmXuAiKfF5b8P4unLc+AvDc1/4ZlACo4XzhiQGT/R2TqZf3Ny
7tljIyRHwc0DwM2/wNBe7J983XXaMIZTqJTkYyT1/2QeNwET5jCEKOFmmFfcvlMJfjToHuHilI7b
X3d4ZbUVCAQd9aVTztXxwaHX8J6cKxu+oK2vk1bsljKBS/pZwbzKqvJPkwgzHfhdZsz2yUT3xQwF
GCC5tQ2GNooSe0r1bAjjej19OCTfE8ssmYA3MtHM8mDtBbetzQFZ4PFlGMhItGLSwykolI5hDxsa
BJ8cVprF//IapJU2D6MykwQLywTm1dL+Oxvk98EVsCN+1HN7jxBUZQXA5fpqL44mRquDMkO7tRrO
pdVQptds2tSZbgcY4aja6drer8nkgUggwHvJzokldm9lFnGGrp3pcyB+UYr3UDAz4pP0DhH/AYJ8
Bybn8vYiU9CToHtXTpH0x8D4VEJk2PSI1HRL1hybtwi6YfTbzxHyHlmRIyklU8OJ1nHWbsBvlupU
QLwC5ACwII0t97cklw+SHvvUgVZkBxhf3d5Pa8sE5NQKEul6rrgoZYQhSCMqxmysACc6GWR+b43O
v8ZD74D5ECmXLVwZcxHoy3fseCpZHz7100mUgqDh910zKtvVgnsO9vJ1cWMT85Tyu7fNYBJqs1Fo
bJdIFwVCaiR37/MDc5TLkqh+FLNTXYTPTr6v0l/dijazUG6dnhyuihCTgMoy+xKFlzUDDz5avFF9
ns77D52fowCZYx+Yg8EgPMIqC58AB9+5tT5KMzSrL7Dxs/11dDf383t/cZB92YyG0eJ6csHO9EQn
awsqUEMKXkyuGMtoPEDlaEa8AnRbF33FeepoAMEhGwsOfd4+4wRLzehj5JhU+pUXj7Y7StOmfkfE
wQNvoxIuQ84yHQX6CeLZN2CYcDzGA3z4BZUGzV5HFJPxvRE9O6pall5mUyqIYer+kr5VdD+zP4A1
8MrIOC7uqJGRRSzmnGaZSW51eWzudufSX6+Zoj4IoqVMq814x3Em/VgGXYHfjvmXO41tdHe8r4eu
I191+ECbbsNvWRJzpJcktqQiD3J3fKMZgJjBuTq17n8XUYpFY3Jl98LG3MbOQj+hpf8b97VceV9U
5rrTRgMHbx0CHGUqeUHIPGsIufhKo9dsymWAZir9d3hCwI/A2DipC81sgKaZNijDif/uLb1jrdlq
ihC70hnInrTITR5W5VTILc6v5kRJiRWeqQ5nsRF9+tdtwmmaESEm8dYpgkf7NizLZHyCdzo+Ov04
s87+oj6qyAZ7WPBILrBmqRSORFZKnzzS6KV9q2fB4F9euoPPqyMl2MgBRf+zeHU0Kkkl7pSjEsxi
ZsqyvWifehBzGpXiwb+TY0NEX8lgVITmRPW4sp8z6OqWfiWIt0uiBcCOO3R1WWYDS0KaffeVt6SW
xfWEgJewur41jJOmVaANS+ldy7kwCwoPTR9RXWOtET9nEoA28jugIdCFFNy0F14rwU74DOp97Eqh
4GNRp0C1Ju1hhmTgxkEbY1ZA+Ls6dxK5qTAgdbKd/CeP0Wkq6BYM28SfmjPOn4ZFI6U9XLvLhJo0
D/lgMOYRSR4YM9YnITsRFZBruMz1tNgOERutjpT0jQQpvqJHzx794phV4ty2kMqZ1ajJKmmC3/iu
ANIkDgVeZPsY/cv6UoOkTgspRjatKHdjIZN1Tmpz0TEihfpQuDnLdfsQ3hINd3J0aP2NPQgJD9AE
rVJHoRDAicq7Mp2gLCHv55HhGAJYdAatcqyohAXGhJI2CaY3yAnFY0YZvsg7I0iszEaUvzeD1eIU
YI/+E1J7I8HUixGMj48g76F/UaEl390Zyc6uicMcphZOg3vBSvh2ru09kg+4EEmSK9nuOtptOYIU
0OGoZudLHm7g3gyZBCkrro3Ce1cF7CQ1AOgGtMQKE3iA4DOI0IFM3pJ06+MMy4/rSPgjzI+8tf9E
jte+AgPPqkrdv1jit0xDHpedThZqbhVmJ3vxI718K/Xbfops9f5+JEbyaDwk4cCHrtXV4ujEjnOl
k9ZY2PxcK2Shyxu2/JRKs+z86cXlH5jALXkl6lIl9bnw+SPSe63nvx9+GTQ8O5tak6+a0MpNUr99
mLYTNzAlf3OYAEUN9CZRowGGruQxDs7U2tgdyRNSqSAT2T9D5AGdT5qTwa1TxNP6P7fset0aesox
hQ9SfSCmVcpPmgT+XeF/JbWCgQbhqUEBonPsyqrBzaaLjiVXPx0vPhaA6LiEGixJuvHjDa5NTPoz
fdNHS1mHkPMt7e+hG87OZtHok4gwnHjxZgZQV/ovbRMB48yIgQW6fNoMWL5ygsEv75l5MXPsDoqA
BZL3f8qzrZ2sLjhsM8qypqlbC2cgZHReS0KqLmCume8fB+srztampgGEbQuYCsZLkLflKx/83L1l
p3M0uP9deYzRd55pq37C+ydxaY0wg0GMBkjHkWRYCK5+6eoUdu12/zeDHpALYEW9IDyx+zdL2BJq
obNOWlYqM8p/qdSgB25CBV0z9LOpDjftc1+kgmSi/IGJq89ojH7lv57mAr5r68Z4L2cs2aM7pnbs
srJosOrybCYQ65n2Zh7GW7+irPf2USyX4kpIQ8dla9OYGEiZ7NhLSjrQArdxezUro8CUOCPi7Lb2
uScudU3zsTeFcLZcDnF5klq864YievI1sFnAQN9OufDdAGiZCU9vLI866vlIazef47XyCwXB8H7s
WEGHZX4mpHmk6WxRGs2aBrmFJQLySVZUmi/Eb9Ut/k2FgBVjzr7pgOXQrVbPLKfVBxDzdQUEwFMR
0UcEPGw8rbGgsO9X61xH/UEUXpXJ3ltYHRyuNv6xEKiYcnf0Efi5Tyeh77Y+JHJpHd4T24blZw++
vvFnLizdcO4rr6MQdA4PaTWNnddd7Rrn8MtEyJHid2Z/QWUxT3LBjHsL3XE5MQNu+PXkPZZ7CEE2
WWQ95LGGtVc6GMxf2A/q5GuSXR6GfS7QIWfCWeF+C89pMBPpOTuae+ZtwmyqeJUOWeC6o81xAN6t
2nhlDXb/kSWHG9eAcp3Y0gmrA9YyNT8tporVjeBRGWmZ62zYajtUPDKO/NMOzATuB/zUbVZjxu1i
rIqSx4jeS1c2erDyUqfxiNGy57jL1sS3GNPLcBJHaZ3yrY5LHAl59JEHS9v/aOCwXVu1gZqr1dYw
dgdNPFgkAduM0k24FoWdpgyaDrkh8tev8iVnXqPLfAJoe0ufO2M5KAjYrphizL1uN7EML4qmVCgB
a1sPbqCSuajmRRv6ASgwduYPxUSJYkxLiWAcXFWBDrHspu3hHO/uKLRUYM4N0ZqHS5ie4Eh4yRBP
0gbwgsEhXiD/516YJIEhI5N9Op0TPrlRmSTyNdkDLzNqhTHXu/nYUOhYed9uL2hQNjG0Gz6tJ4ih
jJJ+YUlJXLPVgKqMgqXV0kk26tlVx+DxVJAYW8Buxfb5CcHEjK6rcHc0dVjjDe99Fqr1wTlV+v5k
5jAGWGWjigkbEUop3BE9O50n02uRaEoquB19h60YjKzJR4kZ++dKJS2AlLIv6uJ+YR1q7tXPc6CM
90r4xFDKdf6j2/2KAl1ma959XKcUCVrlXLyT3XlDOmUkmcfXo/PgzHlyw3xD17WLOQKIm5mwN/wh
26jcanwJh6WHkYHme0dvV1opSP7F1sGxCyyy8DSKt+ZSImnhbO62pCLmzk6WDyqaYBEDunO8tlt8
o040m0VKW2lVqLf1p/M8j03t/Nd1YiSrEjq5ApjIWimBMvIqNJhUUxptcx0tAKOh5sS/qOFKYTaZ
sIDbR1HBWOw1jVzoyviPt+IyPpLuB100hswmyID795AX57hZvSUi1bpfzjxEwjukp7dCteZrrdR6
P2k3pJiExsC4EqOVlzCIM1ROonSgrUnSJAxmaW+ho+cITqFf1YN/RzUi2oSH3nDyi4pRqNiLe5VM
ZrMYDMkUpYI8juyTzdoa1FsGNAx9Qubd71ww6QosVjHTMy7+3ajw4eSDhQqqtch46j8NL3NFm8v8
JJtDzGM/tZ/8dSDsk+ihpQkncYd2Kxn2itu41M5gtOveIXegvz6JIuQ9mWB7E5P7tPZFgv+3mvNf
KB/kh75PFGW9/dYYVj3Xg5R+T6hjZpIQ04x0/y7eJnuKvn3vX7wJBLAKH3yZmpvZOACPM5Bg/Qlf
2EZqiuOkQwck4f0o2x2GjsoEXfxtLuwVttBU+aX0SnBXcgnpKlWfuEHIryiujmUbLrbjlz61NC+n
1RTgaJoBX0xucwakiLYVYx/J0D7nx47muKiZsgB1aC6JNOcUAjJcOmimGHdHK0h8+pqRsXryYR8L
eAJeuei3O2/AquhLzjNxklFoYxba23m3COe2TDk7BqWK7LDM9h6kQpSxYSc0Xaru+uS997zhRllO
RKPlLLcwgyBq36Qz5+GsSxzMfj7fBfcUpU2jcx68egn5ak2VkUYUJLUlVq2nLl9AJHiRoOIcqii3
w7AfEe4BtQAgxQvvQBeQ0EYwmeoa1r4njjxVd2tcS8sX+nT5tkQME2oJv5RH7Cex1U2aVDiioekZ
Q/1c3nfvi8q39p+xNwcZfAbrD9jY71Zf07csekGbz1t1CH/SV77kL8O9pJYTCyf8Zf8WhrCT1QgA
1esZXMEkhhf2YLy7pEC/WCeBA8/C/BHi+cz2w+5F8rTRxQR6h8mMh40e99yUhyvICANXPdbWNMpA
dJ12rhGFvZRFfwAxHbvDmJfFT3vTfxl/w/kV7CueBltOAb9t2jPhj56mUMbReAU3fAH4g2U8dJ0/
Nqo2wTqt5rMlI16BKRjNVOtz+6PEcCc0fkt4rdaqVI2pyJgxLNuJ/j5o9YHrXBbuDEjwNru0ks/v
zOokq8EPNaNTHLwUOJ8LcF5wWuIM880zATVVxs4f/nHC/TerH1iOUH2kjNTkdV8Az8coWVYMxOF/
Okqzh9qTiLNBGe+Jia5A/i+QN88VsSxpdBaNKAyJ3TbptVHlOZvUpwU7+Z3c2O9c8hdHKfwza7DY
/W2weL7NxovoDflGi4v+yYvLt2Ffs5So8LbvZcNnGJ2nY5s1ikK1CtCv1F9QzxGufuvPKnDd5eVO
61yAvvwLO6jxg0sbTOLijAveLgAKQX93GenTlDU4rtVKaMue4I/K5sHZ5fsQAMafOjrMrTzwcHiT
MW2KZx99r7xrraWdc3H5adml3jBakSftGlvTsFeiHwXLnXXKNuwrw0O3zwipxrC5IYyayyAoT8LW
F8tI6AMnnhYpxBA9pwUB0XGnFyzC3H9xm4g9JAVp7rEou5JwTDJGG92oltNlsqQGB8zpxbgcO75I
L/igo9wba4y3EszJNuN5y/dvclU5n+yqv05ommwP/eLwU8829+VdGTNuui+PXmVOEvUcellSgwvJ
BOLuanQFPyYhMXXC9AvWRTHBRVmqDTHzJHcwN0ge6dEiFw+dN16bQ3/iApEJgrE2Qupp2yCnCIhS
cJ78c9fYcPwouo/42HO8/1YoBKiMbp9/qd4L1cXFypzG3oVIVyEzTRtsM7trbBVHuMj5oRAeiZRk
4sksIrprGyvSz2+9TZILfhYVAAi8Yhtd9lkyaAP9x3wI7RaQ3ebyNgnQgXciphk+CuNHnzdPwCOW
bbA4b7CKD1ArcqTm16kNunr0reMj5TeusSShiv5JWaN/CoFB2oD9i1MoOpBMlG0INRn9JnvVGeBK
eq3UF/6/FySbXZS9Y5zyPaKBgMLYu/KphP8Ngni9dv9MJeW46U27IXKujjFMSMCs6Q3915tTvfNn
Gdzm2hzdDdagJA5fHrNq2OWWNTLOxI8vNKfvlr8WobxY6JoCthvuky4Cptt8agS9MNf/EVAzTVWT
RmXSg//B3qEHsVpqCK5noARnwwmhcYCjnfhRce8Uza+Dw5htu15zJ78La2KUgloW95FPMcgQ3Zcn
0RYua5mQ+6TpISFrgHkfjf91Ts0URoXxpXluYKx41TZrKbAed+fMRdW2/y+5Pfi1qNKkthyWs6uZ
9Yk2RSBmXt1+Qv6gC0Ixh2kfXJqe0cjNXZCugQZLo4TL1ElAQNh4697lfpaqgrjEC6a3/xugsmnb
eGklL36kv4NxjpHpxlROEBqGjZ7JmSrEj5zdvRRDwG1awiO4Ct/D3Uh5akljhsSZFt0fWEpd4ks9
2hTc4oD0/UCz4L0a20WFvm/m+sJpVm569EgWhpkP5yfI5IDNpTDMDZlPGZwe1ZNpOxRCcRAAc4w0
kRHjCv9S58C9aiNFxS6Hj2RfkgEmrGywBYExUN6ObVfyj4URdu8ahqSTIkuyTx3lyr2Q6WbxUtI5
W/yk99QreLqxCQWNcrBeCl6qI9ie4mfkZkgk1o5QexY2yTxLgWvDPZ8RUW8UsiRcTo0NtUroQQyT
LabRkw7OwcAtqben7m8eAdP5YnnlWrFyLIGBsmnX6SorzjYIrbNe3Bdz3+FPe3Rwr2F6hPgT5KHz
wMkZISFMS2ivXmePfDLvd8y6sc+lwRmiB78cSlLekleX5hwsW2WP38/Lh1QBuUWWMPp894MuVSWn
2zxgj+p9gmD79ZZgB66+tII0YG182NBuAWtkXfnJBc13QDJg4DyLN200d7VE1bg8nYwHMnupe0O7
WAUspBlO+iXppqnzZH4DLJ4MlOvPb71QVlBxxwhfn8wrGo2EKE0EfjKoXcQ8jBOz2d+qGfghEjL5
hkJ6BRNTQHujJmH6s8S+vBIaAng9fuimMQdHm7t6McbCCpUFt3CzjWsKoQQI/QvWjgOLML0FXzQ9
E37zFt9qI/JfzOyeEkPlPSrakej+yXc95qa+Q5AGkWpNG8VeIO7OmsuCkKN8ddEbk6FIaEnIO24a
HpIRlgmpOYtt+HtHamv27yNERpl4FxDfPnCeQi6+fFC0S6tIJe+K4NjwyrUcxVStxUfDeM2A/p4w
zM+BpssPfOJpN9hOxvWZhfbShdMo9A8ZRP1q9MGNP6qqZHQwl4bKNDZ20Vaf6NbVHyW/7oBePawu
fATvDiRrlbLWcVBCPKeK9AU6Zx6bfCYkeAPEitCfRQBGagBEWE3GQhD5fjMDV2H75L8+3gNO7hoD
oxvuuwKM395uQLdHaKv9Zxky+iN4PAth38rLgaz1bUo/iXoam4gMoOJtM1LY6i7d2l7xf7rwpQHa
N9X9MoFlhbxT72Fdl/MKPGTEImHNrff9SAmXXpZEFmjWF3fxkgcHICDkRIwyD4SmUZXPi8kI7LEt
QrVaA9BI81Q30x8/Mi4ZZtSvWr9dGzpSsHb3GXEdSbRQrwGS8GdLsw4avX2ugWGNDiw06Z+lLW/0
pbmFzfznOV9xg82MWfIWj0zxokNX9JOcv6QstkkWTC23x+iRF+7lD5IMoi+DILonkdlANb7XM0El
gtCsQJFR+jQymLteIcBEEpw8/l7DD8ne6mjwbwHt+LoVCtXERciRohTBEDBTITQQLzLAv3nJcxqs
OOJKCnOTttMnRuxCCsY3gCJUT3PldRR8VQYInQNee6kiftvTLzBIcR21W1OL42ZcBT1b+VrmjoE8
Y8/lDUfJbWrsEZ9pxKIygisbNeS5A7FwlhgAO/4koiIPe0tIiS10UT2tewftDVk/QyBP8/LS2BBa
nMv9zC8UcrpoH+ciqz1kuMYJ4gCa/fmGE8Fo9Yf/9HFuaY3N1SpBqXMIbo+WxFVHh2a1dZg19MDO
HLo9CiEa0xROe9TvssFsCkiXgJXGQfOhd/MhbtHYjIfYcDTnMH8kg3qwXWiqayJWjwv8avbuAIZB
sEFsCKMz7gJEGA2Jc4lhLTswmOnkjyTo0HEZiEnNbqEyyGXNGuHm6q2Brdrp0YtUhr31CdyAgSOW
K7RHN5Q6gSDNmEvHf7Dvfv2Jef3zJt2Lx7W2zTyDnQkO7bOWXeQpxqzL05YaoL03cWaMH9FjWAF2
T6MpVRA7FmIsp533p7c9bWR5jM6aCI0RhORTyA8xHQYUQPKxJwisuApqsvxZbM7ACaPxfoXgOWUS
IVr4SlgK9eviwc9fuD/TWWZXJE8Ey34roshPMScSCuNw2/5aBbxrclaYGnSTaIqyxpsMVYXlbyBZ
FHJX1x0TjFigvQcTI1DmRITexFOSCN1LFGJFcgBuDrSJcw23iNKZ/50WKJdkZuGdmYSDGR1To8dc
RmByo/7sMKcDUNzKGudcuCfBhmEmaxQSXFQB1x7BzqR6jfxOfbm5xsustOxoPfcO0J85h5/xfxZl
6+NZ+wjfs6/awdqz3PCgNQl1VM/SWho9epTeWXC7+ePApjUTnty4R7JqqHqRMMVEx216adfV8c8Y
+m+Q4HUmO7D2HljQnDHeQnxYyP/LBAS/ppO2cQ5ZYMn6zIw7vKyWn5HSsBF0ntwS+ZjQMqtZiJZP
jSl6D8Si90C1E4p1JdpnjykDQtpwc9x5NJu/Id9y6YHFGjPjY/7N3V163YrGS1U2FOawkweQBGfa
P7YtrJF7n/E+R08bDYH+nho5gXO+A03w8J5CV+awPFBbcH4edmgIO0Sea/4bb+qqOdbA7KDBq+j1
mY5WSes4XizVhNFwUdxZtpDHFz6k0wfuqjiBYdCljwb4veQkd/jkSS0xTwA/r697FMrNt67GtxUd
NvHJS7/uTApAgrn8S5XSqBTcB5O2LZsfS2x5EysR6DIjQmL4lY0jjTeOdpeBmHbixGXAd6Ul1MfC
n5wkLKqNVQAwJpWuJ+65oS6C4kwL6DTtVtKHDT67gEq932jWXJ7WoOx+nsJRhBI7eO6VAGOTtyBq
jXKk8ZNOQYGEVKvfxsZVEJmgydIzr7Y1pcXOHPYlcqsuKrlOP/LrglHdv8zG+VDfP9wCFrL4tYCz
hMI4gsqXCZ5Fvxgo4+HYwKaI2oCMnSEN6/DW5b8rk/uXXubXUD/3vUF07CM7V6vo3azFYHzIDwAo
uKT9KK2pCRIVRdW1XcTxu0781NsVcfFCJ6vJhKE49oH0XcaixmvvY7d/j/18ZDT3Qd9kR9RDtbVn
efzvAQiibDDIBp6JblCG7iUFumOw5KvR0Qz+YbnIBAHFVJhvi/1ZIh3Pyn60PI7eUsuCxSQRKFta
sjdlEROPa5p7AzvnEbYkJmX6mdEbJ32u3b1qrhUpqXWoWl/zGCy8z+V9feBb+YwkUqbnipyteYqM
xjhvdunddWKGAe8OMhuBLi+PBFUsqlDr1r9OTjmDWf/J96kqVDxe0EOu4v0ZPCXTmISmBbsFL+JG
IXmGvU2zsWLXrShhL/S14AQxNX+SlvHZZWaJ2iErgKAnm82Ir1AQd3LEEicBMHKKRumySqRFC08z
0Ud2X5Ywzc0Na63DduUp5Jeu0xU3HUfzrRcSRsv6b0UDtlzTl+cp0IIJt6M7OhL0X54exD4GrJwi
bgPMdRp95xgEiF45U/321v3txVeJJm5aVKVddF+TGD38TeWKOw7JL0nLAOwRa6r5+lTmMUgWXtiW
8sPJAZNA4n8T+v+4G3dk3vIuKbA7PTgmqk/wR8TxasdyGEVPYEnFtR2DyFTLOPcYzoqZzw5+TfY0
ouQOysFNVX7XBz3CEGkGOtya+0u+GhDeMTnPd34xlmzAOl3o+s7hjD11wsZvO6f7cHqlI7HsrsTb
2HCR6+gANajuX81Rfx+W2NxWeHTArbSbGgJB2063rkEQfFKyxJfPmb/guClnLzjuy84SwUpopJGL
Cynt4KD6Nj1zSLoTpfARzfkBiVsuiNnP04Vo9M1NbV2zPgmQr+D3m+zaDQ+5F3WU27w2PGFr3i2A
i7Q+/r6xLhSs+LAXE2VoZhviRGc0pXrHsEhSyovbv55syE6pMpm2nxO4H5gAyG0au7Z0j90V7sHl
U/lo9qOKm/D0rzXy4SWJthKt4tgGoid8+4dOi94YOFw9IkweeWZ4ebO702j9g6GXD/WVvcI+JrP6
c5w8jRTdkjrVKO5FxJNCcHIw3ORnyD4bv/tEErBHwQuvfWRNdXqTB/3dO4kWyEjREzCd8vB+8bXj
Dc87MvlV/eav3kJzVqaata6fqLmV86qHNSTR+pmAyi85j3S4VeyTSWIvDaPNGFuWGaUx4JhCcgC0
7HzRxaMdpVZlPnIGdxiXcZ2lzx2Vtt7FWojxpI9C6nWZ17ovI5z6f/nEtsrcUOd2jVhM6HRiv8I1
o52WMMcA3dEVYsq6CnP5XAGUkEuDIft0q6W2xWy5DHyiL3k4ExlmUswBRY2wEK572uOoo4p8nalW
TBW59BQ2lwrlRwTObC8BygoaHwAFaipS4ABqcSJpAowxd8c6t1ffZGToDzAPtVj4O838tI35SWxC
UFJN7eMhysHcci+Yp6OLKijZ+gVcFjE2nvox1ZhA+o1V3+dSBKtjrWpXQRMmmrIIJHfV4+f3YIMx
oR0cQfKBCWns1KJP4LakVxcaPzo2wAOQ+8hrsS0r8bXmLchyjIfsAD2upCep9I/BjS8F8lBfhAcg
dnN+X3rRk7VOASP3XrPkQyoznzt9MXmIHgPVgGT0QI7ayORfomPed+nLfTEUrbC4vKYMbkwGKUpO
QuBSVMeLIuCMSPDwWs2kDylDGVIrV0W1wGRlQ2dSbl6ZjT2K11B7uiteZAyl+HBtZzrI95+92EWq
BYeX9d74o9/q6Xlz8FzQBN9A8LDCWcliByXa1okOiMGNYiGmF82eg0urjT500F6nuD2M2omPY4Nr
WpRUkvpxxfHpz8AvIzXImkyh9TLUUcdBqV/gy6SDj2sueDBM4QHsybSZkI7ES9vEdSMratZrX+6U
1CIt8wInAJDgAmtDN1YWnPLcRGatVU5qywWdhyFwhXU+lF56XLn2Urh6vrK8Wxe95wnaVv+Jm9aP
+Y1Yf85BiCJOop2qEY6o6z5YTxJ+heMWclLeJcpe1GB98DyXJ8r6vuGSJB8KV4V5Fias4IgJZ6bM
AvMJOjlqqSQflpuXKB1wp6SMPKJitOUUt7r1ui4OLnQo0EJqZ47/EMtpOlTEdzR7T8eY3kIZ0FGv
69OEfC7ikedrU/0V1KmYnoNUz9FLnUAfwW2wiiH9NPnj+A5C3cC9DFfQ47gReTy84MZLpEHRc/f4
AWUa/Cx9YdcTX1Hz0G1GaLCMIagVSgTXxLckmHrIO4hJEiDKm1CJDQxd/4Pq05i+KjF3ssGWXyK2
Zr0DaszveUOJTlI+8q38iK4r5wR/GNrqP8dsDYmzX641x3mKmj73R9r8G/tGNViAO8G7Sag0skZP
43Dj20HHjV02xQ5J3N8a96wrvH446syBUFGtuRnqmEKyLKHrDRjG2gL32Lbk5W++KQB1kqVcMLL/
3Bh5a/lgKF7zlN5sVsJxsEUE8v/kCgVvY+e3Jf9FnKu2IKbL7QD8Wbx5aNy/LrWikSDrbNqlV1dS
Ss4hP7I5osSq6U3MtiKt90vQUuh6KLXn5ZciHOgR+hryM5h/oU4aKH372xVEJATYGtPimxosAXPc
+ZFh3Aw/A/jpoTCUbIFdmFEqqhSO4EF9+n6IfLTvTvmRmRsUNXOwlMgLm1y96DnzRMTmVPym2QZi
Vy/XnCKnR+06xwXVXXqMWuEaDUmrp5sW6AQtVd5Z9EKD9U7cz5QxdmtCkeBgN6KadeGNIh8yuPjU
Tg0Uz5kSIDh6ejzObcHTTHsmEJsmeJc4hUexHCrcJBqM7muqnc3OZ2bFT/Ydd5SfTbAY8gV+hCdX
a90rEkHtGGftq+mg1wtNo0foM0y1CCaigs2FfVdZMvM1rfWxdHsSDE8300XOks6YLmNF3amh5pn6
AWA/VyVGpFR75ksEf8S4Nvqt7egQWnlBRh5QHT12SrT35UrNOtzANDng1WvF1KccXPOViap/T30Q
F+9/ICTJfNxFOuHAgDwiS98IG6CIriVSXYqG2YMLj/gNzzyt/hGBUlYklMqtoRjiPQTu35eZi4FM
dt/c47PAnL5l/rEW8CdfGglS+UTHl70rjXoBw4YiKkP5wOm1Tv0yWvTxXCev6PA81wRKc+aWIsKV
NIHumJ95BehU5vGYWzf2nz2iebbYWJFdFrMOkc+xOOpL3IQHhxzEjs+SvLCXopIMobpWM8f+Eryf
cDtE8EtzP2qwN+vYvIRq2Hr+FVhg1LuXziwWrp6voWgdeyeHi3W6MdN+1q1Z7bFtYD4VHwveksFb
8Dx1fbY/dDsLrlVIW31uNVTqhZt3O2BM0DwjGDEmkLuY8PgfKhe7IsMj25v3CQW7SplTUNU11BVy
hkogx7GjkyReAd50/3RzXk+vP5gaF3Q2EijSjFaCcu8Db+9C7rsSLPx2cytUqjApJIPikvku3Vwi
MmKH5dODq6vx3s/8EcX+QB0SgaZclrNfVndjSeZddRNXASk+Pj/J0Kuv8qO2iJG8uVMzt/PH5WH7
TglA7SJ4jcyEi5tY90wQHO35t7qfFjaJfbWtrGfoHGy+OxMh4YSPv5sA7t7TWp7gVlA1yDHc/EmO
9w57QOtEbxkGb8Wr8Gewx6VA+CfrhikSU42RHREo1BYFvfPgBicGuXpqIZBkiJvIo3a5eckbHH4L
ccSaFYuPUcyrKQwVpvw78MLt2ZKtfE1qyIKkt3RUBWfkvKb6GQ2K6na2hJ4Kz+2+Id1W7+7dCboB
NLSlSngU1ULYGQBmpQaOUNqXhChdGEauillS05FhqXAW6+iENyC+oR0p3lgnPxDJpgo5VW5VZWNa
1gzyUJw73CvFtyzJbksitO+VnHFi3TFYW66O+LDqlolJ4F1QtylahdMNRx1bOpgGmzJlvH9u8GAY
+uUXv7XMzlrOEaJ2wkqDwFyfxfnr6vrtN4opwASRXLwrBI13XiC/0Qv4KFCDouiGzcKDq+/TbRok
2t6cCFbed87VknlPuHCScEXjdnJO1siivJZZUU1WLyyYmMzdRSfnW5s07GqXS/+E5PBr3GmC6w57
28xNFNsOmhbfndw04h1tkKGWXJkfEWD0l5wKz1rGt2n1C/DOJ7Gh/RlM50ZJl3WnK0WMm8yr7r1+
HAwB19b/oeussMEQUU/cD3nvKzEN7/CQOBfAM55Lj8eZZwDKluYrN0bxEdWtGMurOHMC+oF+Qhe5
ERQu8MElMZOgYwQLLEqpzlHUweuQ5CilTODfD67so1MJkzWp4KtMxZynHnixxKwbgzGdm85m1+xv
FO4bgaDGLFHUrmnHv17up3ODc/4W2HgaGzQdHHUXekdhnvpxu/kMiCYjaGSmwLJ9tz4VHEqhMMz2
Bwm1Ta3ddUAR9NCmn8bpbC8utVx1GXGoi/aj3er//n8LWSvTFiae+ssjVdJe9aI24idejk5xtv3H
m9dboG1NSSasuS7kgPuSsn+uN7qOPIx6hxy6Qx6YwiLxljWnemyOf1gaIE6fPF4OHK4I6J2jX5gW
gBX3WG3MKvoD+mYDprgeGfoughCAbmJe7lXhkHGdCwumQyC8tTMfbfWoMAuP+PhId0jcMjnHod3M
6evj7QoAC9EjS1jYDngY9IUkxbmD2lFZ/Z2iTIjtGiXhHnAQ5RRz1JHHvvapOrsDsgEodpO0PkaM
WBA+ctcVneyGVQTU+3OdxT70Rxtqx0f/kr+18d0kvX8nSzC+T5pfeGZx31l3PPN+9VMXUIjjEonr
37rQ9cXmGAzgSTL9fM+OM3QE9t+Ic7pukWVDSN+wZDZENUQoFRA40QH1Tx5oAnBD1XLsFBrJl4ss
GXEBgJ5AkUxh5oOeMV86U2YPcQPApohe9va4rwu20mU20Kx2dwNxOE6YB6bk+Wb52pRbH6gPvkOd
pOONIIrdxltVsN6JN5raNZd6MWI6xdp+EqxaAVZi0ixJgzNtaHQNkYm/fQ9WHUvDeBSy3IGTca97
0/z3Aqz/OCb6udD1eIz7+LUsHNJGAmnRA3rGmmpzMrAASdB1iHDrTwn8ATyOCyzmPX1PM8nOPtsx
aWKcbpCFAEJ2cUy/G2/1iOgF7scIZyq+PAZxiwBpCt9sLiHgrsVvdomvui0cP7F5t+zrexRp22Sq
W1gMV1B3X4bSEe6OCpzOznU9/Tf2hhacu/flGn0TxDGME5wXpnG9TN7+sxveXzXcnmS0Pomo+3Ip
+jC54nZuGP4P8Fn9oM5zfd6ltM1v0ZqEzfg8yMG/cSzY9CuyaOm7L4/nbEel4JAepuzoiFnNrD2w
eleOKhGIhxsC6doim6l49CwUyHeTPeVeE2wp3n9KHSphUKvbHI+Nw2llu6pgJ/gUz9HfqIpeKY3A
IQYEY90zVUdZlfM522pgx2yq+PqaPUBiKwfS7OltVGyC/CY/sB3GQ1nIuZiDJyb3jZJzvgYaIDxk
CbyjvzTRlTuiNMZiuF8Bmhr59PG2lG6QDM9+Y2CJjdjl3oNqy21ZunszCVpE03cgmi2k0zTGqXx7
2s+yKqCjCOY+NiIVMDkh3bAulLuibXzOOu9NuQDv/Ak1aFvSxV/W1VikS5UE+6+0pKNAtlLaCT9w
0addt0CJ7OPu9ktRQE8MVnFRibdejYKCvOkK6soflqoHkK2WukOPFdt2030TjeR8A4FcD3tNJ6v0
l9xE8ZL1Z38r5cT/apg2lVmlwuYCAvdmOhzPv+QjSOxkWRHwu9812n52Q4eHbJu5ogxX4UOyBAdz
Nk9ZdGZMfQChCi/XtEU9VJFocldr8mdVUKjwQLmParasl1GhkAV3KBHD/ht3kFy9+QZzMLrG/kTE
eF0istNmoi85zbWaR4Dnzwcf2Hn/rzkpVXXr+YWes2CTep04bz4whV/8HTFK5sGXFHfcZGPZX7pv
DdziWOLcroC4IM1OePtQwCldZNDKMvHglpPSnLjrUu046ZzWuViVQEw6XvdoabIAjtd7sKDxR1aw
0NbIEE1T/vLAAL27TAWamG9oH7qU8mF+xVKWnfbE+LFY9RUZ/uvIipWMJpVUDlHWqqWzFRt9hSa4
VH/vjzD1KtJ0Lrc+jljQ7MqqIcQgoiwY0qx1jDf2m4hDsgwa505fLU5SqVRLesI0PQcalHhwiFYV
GopKgce0D/NN+hyWa1t80NzbDOibvwkJQ9WDghzvRhLFAr7C3MkLgPGIsGgYCx6heedXA2tS2RkT
qWg7FN3Ul79eOwF3gBD+KYkHNQuFkLUnoP0QLkChE+zjXq87p8kiTyY+GA005IBBkJQEvELEUAlW
IAU3Ix37H6Xd7H8W4IoaRk47xiGKf/TftC/pkvNanJmb5124uAl1wxT0I0uvpMFWxPnZ1Bw7YT3S
jCf6VTmKJ3o32gKyFASUERdh7uWygivjTyoTqNbyAf1YezY0jFPm1B6oE5Kti3iGDEnAiUfF+UUL
PYN8H7KNAZEhVxFPxh8H/Wm8dPf88wCShM0eJq1FoexPUZBg5Rr4MQ8fic3npQ8M5vTDCCEyRWcS
EvGBnwsaHPY05lpaX8i00qfiTNa5M7HYm/TLqJBU+hsN8beMGQ+x9foa7obkiGS0wbjFwv9YV579
jJ9uauNapI2CSRtbpYoF4atnweblZ34nW+NhKUEBAnRqCrFebGgT/CMHWc3Deipj6lU3N+6g+qLo
RQUEIrWmwySh0vjs1DZu2V7YG7Bd3EKGNw9A80Xbf9xqmWFD0UGKfve1G7VHbJyAKeQGlr4Rjmgr
AE9e/0tvPxvoCFKCSRvwz+yCURVwrgQvVxcUGeVEx9XPaqrsrxg+CD4f7Aj4LUsdzZNcrblPFMmK
fgrxWP7jhbFO4BiBIbRhMMPEFQujiDMc4gCNa0hAtIZEAUeeHHxnv3TLDRL6SJjTPNVnCVM0fTnd
5l/4L5mgPteyuE4MjdEqDcw+bO2JRP7FLUeEFIVCST0garBVZgcucrqYDSN36OdsFmrhBZJs3rea
aW72oL1GOOmbgVaiQEZi+mj1jhQDqtrp9khS4Cg548thp10JBDHxENHFJw0yb7hx8/XoC665HEiA
g/cYN9/yaQWwnpPltbAW5RBtX+stbM8ul8JXqI7A9QSijBCkMZvhKxMrBzVT1GpZKYgNuGNQ6AbB
b03r6zWDABuQmAEinpL0IkKKYKcJNI1j6bjFuoxQFAlrC/XmUuxrNxI/ulMGBDhtvuEUgsfWju+K
rEkLDyAvcnpYYNTfY/2chOAbKibgj2jUGjkraxY5MQDzQPlYpxYMVjlgd0au/f0DiOhpc45alFN9
lzY61iHQxhC16jKq1gfB1m82PuHrRn0/IhVy9u7dRaCz9eeaGDvxEKFnPxnV+6Di6FVzpz8rdZJ3
PGji9tqnsmvhtgl3NK6UzG39a+CM1iWzshlkA8QMVWOwKC9TgUeFrioE2sJH1toZkE7NqxS1T8JC
G25cT1iJxK5xqYgG+4tJh4kRLxLUIPMqAmkcXNB9Dd1hUP67spxjSdoRmhCt02GDoCdRXWNsnvup
B1SWvBABo4l9YQI1Ljc9GOiV2hv7VuvI1WWMLxb6WB4Txmvi45EJ0BGwNP2Gwkc3Ei4zYDduN+cq
Yehu567HFvFgkQL3jJbJoTmGMsttkaBWUk9zFPo+pCahDJoNISWo31G1c7O3kCcRyJzdsmwivvuo
Yyer4BiF2WtWpCo4jl62SlIMdGIFLchc+V3vqLWopbe+Qsgz6AFdo5AVutqHH+YzvOkVXWNaKflj
F5Kyj6i18o7l/MKhiJpXRZzs3G1y0IyoumK4B45FpP6G48poIrh/v9VHgCZ+8Yii8gXvJlVYOSER
lRYY/vHCLvR8Wcm5gf5oMyKemROSqEBYu68RgzrOD0bIMRFNOjKLG3bxKgjNELbqVkmSxXW44HDR
2eFVK5HSpWfvFrZk/wp7bPMPmx92DiG9iY2e33U+zDU+xycytIhgwuw/ZdLzMFdfDkE+KRE6mVPN
ReRK0UVNRslEnMSUYd9glnDwHmh1kS0g8NhKLrjEQzJSVY7Tff7lFe6DYfc1PIpoFDKHoHI3RvGI
wOM+c+ONIwneCaftg71n6RXXiW3W6qW2nPfYvo05yK2xlTMEHW++PidMXsfM9fG1mEuAZZPB5Q0S
YdWrERUR5AHAjrRbJ7M0WBqk4KkGOYGtCfRFcDLSb+SFVi54gr/0W9ds7MkeDpMFrUuDU6Wkt644
Q3Pt8b/Xl7LoPI4AcGpF13HHj/V0kK23K5cMQIM04M9VooTXjKOOtzCi3jw0d28A1JJhAyXJfGTw
e1hLhhjWtyqQOU4ouUto3Skrv3hg60LDftiacpBduHuJrK1VXfHOL+4YOTBMe8d7rt5qBOjMtgpX
afpF5Rx/N/fLDBYxs9mryxi1aD9h2+800XvrcDYZgC0K+FkjQE5YJ6nc8/wOpgKApGKNmkdCYaI5
ED789C2gIoqS+3FY2WCIq4bvTnpcdmZ82KJLUygvpvbzftzoXifCnqhqvnHxqPXxfXV0sfz4ZbXu
IOHPAq+s4nrOUO2Mj4LoHBFmSY0hNHRrETkWYx/K+v+0iKMZuCCoTKk9BP2sF7Ozynt0ZdXMvb4g
R6gcqwWNG/iJwy5seYkwwBJoPVMBkmlAYD4ZNjpyBsQGytySCu52biC4U2OwqfR+H4UeMjdi6x+X
GP85RRNdrlDC5tP8OMQBFc7/KE/npVeWUXgGNX6FT/QqWkYECr2fzqqeKNmLWe6IABoQpEmh1DFB
SbUZB8Kx024a9jE16G3jQ+p24aJKxhT3KsQFLLDFjgeihpKOuT7bNdwUphYcMZfGrUiuOGVbtEg2
U7IBZAe4FxaMKHxcqeBIEdfzAQEZ4PKgV+/PzackdlSAGYpp1GPKzeXpAN3UKdu1uRteG/3lOVXn
BnP0RrNTg4AJu+GkseDFlMPHk2ifK6CafjFVsLGJFD2yYDmWeTbsUAHR8mg9C/GyWdha/u4y51ib
9Bq3MB1cYlWgQ4ICIUtAS7+XThhJTFuuGnZWhd3PGGpCVA0oGpIwTcSoVVmteXwLf/yJ01rvaGIR
TLljBIJKX0KRzUE6F894DLKiNstZr00/640aOsKMOtZ1EcjHlysbxS51WhKS4P2m5TuyCYp8hXjv
dgBkGcFOMAEyAFg2ASA7G+gczIyr6yWgjEZppvKRgzn8YFzHqdqNRveB8CdhKMYPVllF4MYKLsmU
f0lQJ0Y0qMxPNTJlNb/Ds+nQLK9hJgrqq9RAr/09iSMDsZpwEUqO3GxDOuyJmsPHERdioqDSxezR
qvehMO0gV0ampjP2LBps4ZS85Aw18J3BgnHOX25C8NC3lZp4sBmK1u8bujgrWx+aQ5RjNCDBq7xX
U803L3354mPsolW4CIuBFI4ZQF+NA/JpYzcp3WGvNozwWHvL7lE1MRHP+DrNi8dCfc6qXjQuHgYM
gBboKSUvqov0WF9Hn6dAg47uoCYZMEeVPFjzf7YQ3u+0t6begWMmx/BrVL8Zb2PBEaXWZ544hrOC
tdcvNiN5D9mE03A/gocF1/HtFMAJ0gow3f1UVsOnC9z7DfuXYzN4FMqPh8DVwGOpIKHiobYXD8C9
GK8jsfrSr321F0NX6wD2GJHetZNxlZLUFAa1XACsTYYPT+vDdno4vzUFdhEER5AJ2qaOM12mGFni
PAoQ47xbjQMxkXF6YbN16x9Cgkp40Lco4V0v96vde8mzn7slVCCoGoxsgzRUlMJPOuqlGtEGdIBU
t6/W7UH0j5VtlTG64Exn4n5KXfcFHFp7yaMzQTYqxjWkrQ3bvHIorT3QcA6GpSYvxtxbjQ2sVyjF
IwVSRTuSHsQpXw38tgpQUUCU400Y10Y5ofycX/w9HxUQkSBvuRrLWcueUjJxftYtc25i/PPQfHtY
qcjNYcV/hmQ2u4NE6C97zxR7I33O27Rj2rup3h51ggw7K10E6/+wseYmfBqxQEJLpeim8D2vW7D0
C59fQZugPNGq6CO5Z6FoY4hYMFVmNoV81ScUaNsL+7xoyISxsSZc2aGnW+GkfwnT6WyjnJ4QTM7D
3T9L8Wx2Irx57BZqempKv8TTpvqWogaGNL7xLkZC9be0NNKYO08orx9KkDXW4YbUEl7+C0obK2dg
oWdiJTKoB/o1WWswyXPMStnoZJYwI68Knqm+QQYBUZPNV8Yv+a0OHSCQ53lGwO6pigHHYus53+bM
2fX6xcGG8cJ0+meAOsbIEfloXH8xi6tWKIkbUhwy6XY6+P2eGdwQg0x+gYndF8nCLVDoBuojuXRi
KF08jkcaFsveSP27E09jYMZ1l6QzKBZ0HWXMWQ7fyDLz00nidUOsES4dtpQGgaW6D47gIjSm0Eqs
zr4vvbZVRUmOqWI9abkRhvePGe0e5zYYLQuXxeER7InrFWwuLraxKVJLRyfre/JNezvLEP6wIpOW
0l3/5Jv2pZo4kjSjOhsIeGFjY2b9KqRrtceyscJWXABgQsvTL4WsebR0t1lM2d1uVmNz7gJh/e21
k067KCfK4J9CWJ41mLff3q94WdfV/MPtt/BQYcrmoRLE9CimUV06n8FJ42bnJfRE7diBHv8/DNq5
ULslCI1ubLxn0uWO/+oDfb9X+1AqKXrFKkai/aAyExr/cGKwlYXCg5s+r8iVQMEA/jWf7hZqCbYX
XTmxNCaja3t8Np2V9mvdjx6gGdVZeLB+zbPEf1ickP+NJyKY3UC0+wk7yX/PwPlHknX5PF+UZIij
Eun9WBH3zV+L+NhXmfDRKMm00+HAhZFHlkhdbFhr17SCLKr0Kx0MFn/4NpkKRPRwDJXK0UxNijua
QWw0rGWIZ3El70wcZVceq3HXBjH3SkaJsGHHtS/WzlH6QTaHjvow+xQdMjRW8/cOmlt1LtrB486h
Vnq/gdiHrP/kaTRsYVXWQluY/PD51emSl892lkT2JrlNqRLGNGiEzKEMwvn5FHLxq658s4X2KtUx
pV7VofrgzIcMagGSi6kx5psM3JaTe+AWtul/ToEyMIyRIv0e6OKbOjy6fhsrz1BlAHmipvg2jokJ
3Ih0v7gKzXQZqAurlUhwpDoroSU1qxNGiTf/g7VC4NT+7uwrNuuB5EZudHFZC+9R9wLwfmywvGhc
g4maT8xIjVMO2VoY7mZ8G3wREoYDKJU0kjFMXW8mjDUGOr8cIbf/NWAEY4CyD0aQiWsk0+7LOxzN
g8MjNmoIflqYWz/KqAvCMEXyl0XNcnCJ93JF64+XMRsujFQhTT+Rl3s3l5u8HeHkXPElrf+X0xab
vPxOB2iyaN7MwUyUh3KMtPSfVg1jtT/zGQA691ZnJzn/XYkxh6JkQcQb4HTCb+03L+yYrUdqppAg
MbSus96XGiCRUjfhDy5JI+1gKpFj6MSTxByWDQpLV3g0ZVO7iUYuGnVggCUB6RdOHj88izO1Dq26
K0KTEFnlyBsbYsM/vY3RYK+AVm+CbuthfDHWK4g3g/RglrE2HkwkXOqkfHZf+nLZn2KyzVDVT1yq
h83V/d95YRSCPuV6QUXpOC3I7FFpMbEJb/5ns8YWlYbKTf8YJNL/m4NU7oCZCvuexpEhOsHVmULr
4Jc4qhSDLjkHzwN1MEHxtL55y9AmLgTnKQeOSAG7X+tXgNs7F4lGHb3Tzk88weT2lEY0U815RlAn
2evVjVu4m049jr8LvvKXPx+RVeROn+OWnAYXl0lCHB8xTqOil8fSB8bFaIKGuc4rn9/4ErLkdwYA
mZIPH3yHxVpt1ObnOuBf3NY42pFHGtip9A2I4wCpnxUX2+uYHmrtZkW0+gHmHxMB+3QwwJpSEDVg
ImMIRsRUfHH1bVpc/6ffJjZfMIRlWHO2ZxgOZ0S/xo+nIcd+j9yxzFwGFroKqt8jcBf0qYNGxKgP
KGxy5/hYHLpCGoxdOqE+j/tLDn1hczfeRWiMEJ6Q7sDkTO0F/h40++qwAzWIs8uCpp4TLX7H74a9
TiMK9TLcVMUzUzGivNgBqWDxIYZ809hhfIIyqF8ACNoURvre+9BCSk8MiMYfiVTHKej36sG8D63U
XbbI3g8KRUldjmzhNYjC2L413xL89ut/NvGMpx9bZxMV7+Xqsz7fnpCEFB7bxuSuH33zWXGWPX66
hLeFh9SVHfNcykpHncbykM4ojs/GILcp3p7YCDS5S6He45aBl1UUfWDbo1rXi0NSqEqjWy8EUEEB
1vDRk4qiCI5qsq04AXFSmq2azcYg8HXdycdmEH4Y4AYQG/N5PIbzv1lR04aE+60jQlgzR7nGzQQn
KG5LTEnTHRGU8bqTarzhWh98gPL/M/3gMLbYhQ4cULtszmqZSfquOKvbobN1XQZT1EbQ+V9ryBC6
TD/+oSz6w0kGEXa3dltUYP34a/AH6DB+/5ApbhoDX+/Yh8olGcGu+cZUHuN/vdmUBI6AUMcCoJ6F
UvRoJeoPVQAU60PfQ+frMAIiRQMDx0DjoMD17h0X3dr9pNz/mNVs/dhYOpHuNRYvrd6wi6OIDJBZ
Z3hTiXhUkbev+Pc0fq/R4VUDUATWP3QS8QdpBFRylCJeSjvwLLwccJOdVtRmOFV9EuU8c6zFWZH6
VxACFFHXrFKf15KOi6J2reGHaCNr1sXpvKZ5IfYmkQoX3Bw7nB9Jptv0ht3IVBY/rGczvz5hv6Se
W9uef90UQ6jZKFZh2NoBI+1F98BAxI/zazEN4tYBcZBBXfgZFy/hw5SoIVbsGK3fUZehTHN3+WaT
muURI2F/PUEx9rdTOph/ZStPqiyyTmvuEk9VTeO3pMxPV2y5CooqaXL7iKdIrcYlyGntycgK6bJj
8/ppzwvx7Ia9bBiq25r8N7MWs7dvkJzvK7TSWUuKT8QcMo5mMIrSy4qRNw1I3kiZ8AVic86WPyL8
4ryUdQfX62xiA03IR6LN/wPrGkigemS4dFrlynugzlMORT+fd1NBHhRy2WaTkCwlnVj4WDdVWN7l
mSTULVUgY6xV1e8iOb9YUMhLJf2MlGML/jb4RJmZIKwV17SlxBs90d7/ngRsV1RUBKFCE0z7zsCo
ohf/l77ccSOf8FZT8CpYM6x+lJ9eUG+5QioGc42OLS41z/QltaDDQFy4xr7zvco2/P+PvGZfaZ2m
L6CV2W+8oJvmw2Az8CBwNkjYENjYQpj/JR1qOr0YU4ubgWMVcfuHAf7vz1dRhni4K60n+96rmivE
ADIkWlGM0Jh05QfUcS/vfWFRGote8qa4LY8w3ilEF3wEUo04TvaoMe8r2j9xMtefxnc4wRSzfo1A
vfiQiIGQ+83g6+GaPm4WaMHwGsG28EjvuHFEtC0VD2vPSSdnYr3ObwS3LjJPDseLJAkfEk7sVDoG
5BYCIB+yASL3dyiMWSayir/9PX5txCzLqYYmVwT3GFPqzI2veKIzcYWxtJCjIXvHEU8/JF9CqVG3
qb3VQSV4UO7yK38Fr9940zSZgfPqUjYAqQoLGWZZ59EKthrsiZxOqUwqef+QFHa/ZaYrgOjJSqRZ
iKGEwHbZLgaOnqvdc9uicrxH43BGvnE0O2s0ZEhGuB/iXCKeea81iOMn3H2oHnNIHl/pF6ELBmCr
whdFEEPhQxVgrbzOBZQwgYRVeKmLlb3BmaAztyAOcvRnjPE2zrfdMtIaHqX0CJfRLRrhnvjVGxsA
ZrkQ3n45EA84sSl6on3L/kwTFjBFlMSJG9bF7UHWDDpqaah4dV3Tm6C8dG67m0PApKa5r70+c+qw
Mm0k1C03UFud2ZWETptjfd+cqgN2N9u8B+ByrKPnKw+nd0N97f3IUBLqzBbIle2zQvU9q1qRc7V2
wulVKY3+lIPSV5rta6x9QCNAMcxMtj1oMnRBW2NBVhtimVMvbbJDiASMWf745W4ZXap5QaqUBOXD
gqkknaj1HF5VMMqtzgc3KvkGe5vEZV2QJHGftkch1pVQ47Vi6yipUECj0bpf9DTUTG3yukICLQRT
l0StxITkapIOC9RCl0jvx2gYt116Krij5SvIBZy+WMpudtOfKRai4I1pEeWjyT5nh4+rj2NuLwUC
e7qdLr6NlW0HdT+lCZ9Q29M+ukDjah+uvsB7GO6SdC9j1f8DjdMC+qI4XASAK2GgCgeadCQy7rz7
GwTOlXR+QM6JHqAnkgj64qscuQlRRMBazwMqdfP5J8YwmDZMhKsuiOyHtD2yYFnl1qAgXy4mHoTd
c8k6jfePoAV2pjm8eUT6ZkemZCXEeCQhe+roV/e6KCqamyoGbLZtYwRPJvB7jSlGdFAaFWAlXxcB
mdve4vOuS57E+dQbX5NEvcX02FpN0LIyTk86wZt9+7DMYKOXJN1fUO29pqfs/Yj2iAwNU3PM4Hx8
nOtlm5+tncW+KEEhq50owqEpDpLkdsn1l8g1X6EtVo+1YRVWRLHf+vLX6M6d77Sw/6qIM/6M59eL
k7Ey3ISE1N0PtWsDD/sOeLnvGckGWL9tLauGjcJsEGEqJa6fQb9+i1QupFZ9uw7PTWUab6GWBO1l
4nBnGyIfMfkebw09ioPqgoKIHGpr2y6cK318B+BvzcspvU3+bGKmk6qX/i2S3QXBLxHoMbDzJVVI
gaz0ilyZrK/Vi9UW0dhk0BbYhAlBFQRvDq+gAF6IZflE+73vhJpwvOSMt0dJdZZdFkVIrTOlT6mo
L6x2KejchXhWai4Drp0Td9qxUg1k86s7zm6mEgq0P0KzFUf5LEkvr6A7w5ldxwNdZQg2AnCCn3mr
4GGjSoczyuvoli1iGm3mg+GiONeOd3yla8wBPtTfRGBoKCxwcLPS07hmROZ8bS+xQQwE2pYVea8R
paUVcIK85Xx5cB1M5fMizis3l3U1P7yU+H8i39oU8dM49XoNHeG905gEov1eNqi5Gar4mDpkLGUC
LSg7YtvrR9ja/H+804z2uRdlduYBR64QFtFI/bDnE/lO7RfLywYsTNrwE/SiW0Mm+ASyXRuLmbg+
VQuvpqs1yA87BmIwks0m1U7Qdbeg8teiHYC5QJQFl5TCq3CoBbmC37QawSReTSiLROPAjDE4C/Mm
J07hHtwywQ++WOAq4DS+q9mrhDmIRfaFZ69Lv8Tw3kM7UJbyu+Lx4hzjZfHUCwI3rqe172UDSdaH
oI5Qhs9Q08VJNFAUO4IWj6agEcWyemnU8+m2ZXAZTHaQyhQMiaezV4wrdvQexIMbZPlmYSCtZ1xH
nIPcGh80ZhETSDWYjltHwjPMchAZ0IgerXSvPdy6yLW+scqVuQ6hTHgLfEeSkL9xv58CaQ2yMfRf
31U0OxRF6QnyVjB7YsKBOBHClmdvPQh+53RJUkz7jvsMgGb0TMsk7mQuS+Jull4MzD5ra159XZYo
3K0YUlh/tLgxJdY4aB7gzDU4Uz/Qb9z3nXzvGD268jRjveTySEzLJuPUYfebrDmjYpn97bZj3eKr
Vx/dGHnBLi4tvDUYc+EdrCtb+Qltt22Ao3b1GpsdfBozSNE4IRcx0r30ucsZ+5yXZ1ZjQIXwdFJF
c9Ln8ZQhae4g/nfxU8xfBkjKtWg+FbOEM1SU6GzXsAzhm98i8f6e/ufa7mOvcSMj0CjudK54zRFZ
aMSinMP/iFnl/U600yM6W5zyEDade+6DqsOgT5ayI0y6wRM7t0fwi1IKZNu83eZooDMH+BUcDxQ9
XSv7v7faaO6pLombLIkDVsSZSYCraih+bAZuRLYTJg5U6x64RTpiWXh7LVkiX1eGJnJTd+073FMt
q9RuMXKLnracmFHHqKDJikesDMxErRNv4XG9ZPtvbgHYC9Rthgy7aorOw3T1ND8Ig0hUY3/HUN1t
L25zkozluDh9fF3W2mpszuIIx8ojUqKNaEckgPWCDcYh3e+AQSeEIR+DXtns73+IMjk2r1gy61lL
5O8wUskzmghmQEd8KSIC8vjMeLksvycXWSDVDEwiJ/4l/68+hYQ2i21WxvXHU+z0fD3B6TtJ9hAb
hp7jOc5ZLjmJ/ONA8B/SeMZd5pHCXqUMagt6JrXSUwXf3UO5MZ7RijhRYBsklQW9tKNEOIYl61o6
Xg9ZcwdwUI0FdhwW2TUEkEA7239A0MsaU1m74Le1lEAsSHUdQO+kMEsnxEi+49iwSyWba+5rz3At
YLt6u69PfHk2OAhDwEAeB7isANj7tz56Wt8JtCl9IdTiJdG/HKoqqF9utPLw5/8sd1t9dhZ9uVlr
ERLPHUgc+DulGh7cMuc7fVOT/3irgx+SQhACEx49QFz6VkLANBUim7R2A/f8vY2YYLhPI+GPWRfn
xODkmorS5tmYVONlIMvAXUL1Y28SkmoCnS4Tcg6XgLj/IR5NY12nlLi5goCyUkVPhwUF+ZRWH1Oi
KKI2O5qQF3JGetX31XG1t/+E3lBvSW7YIyBg4qZCtvxnPQVHR//D2UsUMILVo1MfpnrV6fRYIvYa
pSsSu1XHCudJx5nxIwxfgwYroMNGeRwD6g04dyoKwDcv6ZlvOmXVo9XW9z6T2YmovJ9V5mXY1yMv
ME4whwqNyM7BxItUKBAJGS+8Ky6K2rOrfDTuZbRXGtEURuICEhePwt+NUYCAe96apdlq1gJJZWzB
ULvSkNCZzOvT9bkmNRPfrPx03t4p8+tDvYUHgPGLWFcx6vlUHx1jRqGt04djFPPeEXyNxNV7ObfM
L3UV9J6BZk7/frn2RI6RAQ6Tfa4m1BPexFdXRwocfnIkN4S46pBEPAncWAUQM32/jG4Z4oy87AQb
z/MV/AcDlAn86XYKuduoOaVmTPBKYwQKaPkJ/cB6J0FSBGuhcO5nLMBrkUm8WZr+2cwTvZIM361v
gzhLOs8pg0ezhUhP0uFTKNON83Mwmh6kIQkf8JOKQEwCiwpOoUihsNlmSBeDPFA2pFojlG7wb2wr
WqhhfE5CYB4CoU6iaciNhUOLox5Y8mudj1p2vjxpkiN7X6iIX6s9pDn/e3ptzCAsQdZr1DvLYok4
IgunVu5K2idJ8YzObvxdi23nUJ1bKKSgkfYBaoTpaAdebwA+M9qFpTcZPlbcUrFRFKNSjw7aUUYk
02CEuWKt1lx4z+MLVlJywxDGuKb6j4teUEDzyZpglYBLvjaTlnAh1R+OcI9xqXMCAxrRIKgdADWb
Oy+uoW305GzAa9vfGjYLrN6nTbw+Id60UhYowixDNEim4GqXlS69X7g8Bznhipj0NkqoT5MkFE0S
ykJUDhrDGCWAeeHcXtP8IoWabNXKfkUYEsS5e/04k7lBb2Tsi/3NIYLuH1itKdNnKAK6IExTIHyi
FAw9Pa/u5Uua2rg0EIFGdh4HmNoL56F+N2sf9mGD8HfjCXvQ3SYMTMdmpukzhu333tIKTYyEhhE3
vVALmdX3oMHSZfB01CkbHXhut1YVHlFXMfjxbv7R4wFyRX69xclr8ZukvZPswlEW5Uzky1a1/t16
VJZ3DcdSeU40g62SU8PY8GCifodVlBP9foRJBuTcndy7h4ST6Dbq1tqUoSj4WajDzbS/XMERwctS
MY0vTfe9R+6H1dNWOAQA/ngBevfpAYsvSy027Q3HCF7TnGQXwkJEitbgSAkI9IefJ0IZx2ilFy3+
qmn1Pv56D1kuNvNcda0T+j6cPaxNdUuNhFMvii/Te8ff3QKe2vPF7IP0H57B40llvkemZgfss8eu
9UCVqIFy8EKwzi2TENVcYjFXeJ5bIbg7vX3TL6Qo9iDOE8iYtmOonsO4nZbITCDXlCwvYbALOWrd
YI+29m1rgndeVSQyCGQnN0z5iDd1h2Q0Qt/ZRGwEAK0SURmGvuGKGqMgG1kiIP5XgJKiRtfWSrQK
qgDRKcH9xqd7MO7/MS0ufdbSBmUkf3+Qe624y9O6oqmKTWGEtCBECpB+PO+rjULidNhoegvVXfiG
yLSeMCeNyMTZS0IaPMrg4y3OsLXVqYVL3NCyrr/BOnCglwu2/MhwAtyCb70dPeiqFqtVUa365uAt
q/SdTJ0HfpVBYm9pNEFUElQlBV6RpjGoa4OSpijuYBWgbCSwEI63rML4XhXFiaYU9f5ka2t8gNq7
Diwq+RPXsS0CLp4n6OBb3rDsxCrYbMKDV4OMVxeiDug+riIVa+nb1LsPPCcupvDlO6F8Tx39FfuI
AULaMJM1XuAfWkTGQCk+Vux4tHcsQNIrb8EKO/k3w1TOWtRvJV/h09d56JA3L3vqM5hr3CvuYHe3
zfObqMmh+G80a95AQcGASwExGoqEtE/ZH6WpsXGkLmle0yZBhdSQxgmP1PYDYLrb7wYo3kRoVb6u
yDf0B7FVQDuhYwSI+QqyCrpSEih4a27PjrpGWIq32HJ+Hd/HPCVCro3YFxHeJJZXJ2brmgS/Egls
YJqApQzgAKW8YdVeQ5V3t2UdQHrsJrvkIuM7uH/rsZT1TycnDbWc3k8Crf7j2Te4vQvz+nzVaMae
MoUP1mgLw+6Pe+X+KSeCJdSzcnSJhEo42rnmKr4Vj1m8xJrzzAOuBrjH5PNAcwSCd9pSoZJQTeLf
63PZe5PoVcYbtq9rQTiUGZgZHa+9toFQTYDUTZff9/+97XTf6teGXgjsnRwxhv7wIPyZ3lfwOEWX
sPqkzMd2Onq/ka6X+XBntd0XhvcyXx4FwvC+9wjaIXa2xOjHEADoRUN+EZPV+FKqpyC2vSWapn7B
21/KQYCEu6duNnJSlbRuQfxOfOMeWDi1zdFO6vZU3uazL421hdYHpGs5sZSYKqP/zwNP1FWBh8HS
LJyL3Hi5AbGxM33bxLVfbtYlLW2U2nZ7IXM5SfyfaM/VLHSyS11Q8/KbmXSpSOJ1bN9NojldNgUH
6mZC2zhfUZGD+Yn8IQ8jEay8iwfaAn4cIFDf15oT4uVRY2TZDQnb75PZm8tIVLcjajxNa9ywCIaS
C+EZeZ15mqngyTCJbUh9TOYiPahnSx3G8/GwktF+2bFYkePvdolngi9h55wJxJBwzJ6AZH7IzMPb
KqO/Mt6BI4ZGkRwSycJAYbpIyVX2ZWIY4dpJAef6oMcLwl110UeGM2MrA+RBWlPSo6RmqyV/dURC
DcZDJ5dtBr9iCKHLLh7TIQ8c8gU0Lvw0NV+ysMiByOFclzMTQN8HxJ6yJF395mi7RhCobmVSK/yg
lVj2MwQlCkpB1WdxtKPqZl+WGJxWNfr4aryDRusKUr+D0lZajDZRUUre+mcP/cKeL1UwedJf4Or0
QF6uhhGuyd9k0qcUoU7M/shXs4HcxzIgRHWnBUb5Xl73Lh8jnJ1jHWzZOJ3dHVep/mz9GraQoJc9
tkTqicmYrRyOna0e9wAgzL2Mza1B3nKrfVcV4wCF5u6CTMT0zqUGtLzxUCQ6PcMhHOP0NdUhXKo7
gvPjcu0u5ET62ZPyP6YqPnRPTGFVHxD6osRHXPXyRYRoL4xxPHcCY9Az28jXQyMgGfIop3H0wIS9
IFNoaPoH4HcWWv9OyHbvaTFQ4TTOmcU2ZxFyhLF+N6+LjJsGf0X2QyDIFYHEZu3PmU+bVllemOWj
yF/uuhTZIIpy3CDCbNjgRDPF+FPb81k++fLwYB4ESDL9aRRh8RIkbb5hWtIWEtgmesWJ1I+lh82T
UE+5mRIhYfJVLjGhOgVBluqAnAwWS/iezpDVVOPxxjUsE0mxbScQvT0TNJtPUhMG5mXXVW/VEm1N
DjLKcX/hlzOLkHY86eZonGoCqpWsVYLZsyr3ouXXFpNUXaa7hiUY+DsQ/p09cf/cfTbdT0GIu6vr
NfqTsADmc1/dp87GXQBL+3qUPOngKX8Wp+GyQ818VyWh4G30UIXzSWDX3p1bgPEvKfy7mNrtYKIh
O1tP8Zbn5jtfgHt/ucMmfSxLJ0tS1v1z0kFiyRrCYwsYUMrWWz8R6vTslutvhbJDYrHgw1K/INZg
O3nlVC9flq+CkYFuOghAQyE31L8OkQ00vAwFVfT1v5o5+g5K7Vh+me2Xc4GaZgiGKUa5u1/yQJ+8
C9juTW2mf0a8xt9JpCY5sWAZtqmtUl+8MVMfwj0YeQ4vm2933yXgUDU5OsAj3EuFmRVNSaeBVbRu
60/D9YavZTQy3ZmXgMuOFLMu9AeTn7toQKhflH4xU01ADBAZo6dqD3wnd8iRl0GJTQyS+FRafGVi
QdajP52R29yHisfSAtI6ZARVYNTIAtGRrSbWhLb+XWwwmEUNnSMe2QUi/NLUEMKsQ1/n7saCQvtu
1J8HN5RS/1vTjPGduBip+C9Kz9oi+XwpiIYDeGggFBhnpCPpl9AQxlEU4hThrqEsJH4Wk2UtjFKs
7SUCCOHrzHKcW1CW9KS7nouI3uSpryb5HyJ0I+7rhNUHANlDoYnv1rPguTQEEjeRzX7tU+qlrL8s
WVWC3jRSdQogF7vaBgDH6A5a6UHtkVulG7Hw+q8RhDqlPjlC+PMG5sp3J1qcz4WQZFwIYEZwG0qc
uLk7BF0DJrsK2U1lnFjK9z3EkOaYnKKEtFcVQkHKuGgKWQAuEKKTGys/ueCtW4WrDHlM77/IMnvx
mL0/6xVod+LVexFqbJ8jQa7Cd+CIqTYDi+UEDc2wMng9ND2+pfwOGe8AjWczd2oKqZU72q5dyiRO
XkK2ta+Ja0ZNchqFAfoPQzf62Ut/94P7VIkNlB0/LDrxeS4NABa5WGyjpS8H5+mnhnSpg0HBYFL9
H3zr+ynIlqwiH8+cYLFgVyfEyY66wE/AjeG1uNENoDgLPphZvmm0DYwne2e+XEwFMV+vvhcR9x6K
CcmDuh5XGvfZqzYGteCHAA65s7CEelOBXPqJrw4PLGNWazYqQdbkFR8Ph04CdrhmnVN/QEFQwz5d
Dn1LvrmL8KypcMmNZ4giYPmyxhvuhSDhN16Ei7RGVgiodPTGOtIRi9LFNbNMFTRMjZW8DF3P3gdp
CRFAhyiHpUrZsEPHF72heIT2zYaMvU+drmLlF9L/eMwz7Q7NiTPU+ebeo4RhNjRVxAWUODRsbb5s
A4SZQ5aGvsUcRqsQgbOVl7F2MPPJU9th+2WuwXCf1jYWgtBDSniDiEJ9Hy70UzP+KQd/Ro3p0+fJ
rJL9gOcVb45DbNIiioY/oCy/MxvfaiHhOzgHPqLSf0HrOZ5fbHLTSIEpFibb7FOaDSfdUvjAJTGy
lu9wQtHam5XZuiGPLwiEtDtpicLRJN8xcyrWFmAL175pE3j815CHcD6ZwdZcyYuImPMBUKMcMuU1
wHyCSRoAtobZDfATlIa6inwuOqmkxE6YpFDGpzr8sFLYtluLHtH8BKcIX5m/J0MmA6kUk6mXmGxh
2a3DtNNeulz9NS2UCN6VJctyoqic1tQhBcsfpEaVfKQgQXFO35d2MC3KQ2Ft2O1YzYbrt0pMt4sC
McjgeqfY7/BVNGMdt/aK8HQkYbaR6kzBFFEUSKtoWPrs11g3ODn6fUyvYY8SWQLtlDB3xapm58tp
md2vk//jQhZXZcKfZuHcPf9DCWeCHn3dNYZ6PQjpAmihjjbc7Oc0E2ePMg/sKUNEClAAckNebuoS
ZJW0JYyzgBsE61hAwk88PC3fsrj/l7aKzk+1CXsiZ0PG0OjJzu6ocA7XJ/txnW89H0srD+jj1w3N
5AFQTFqxwHF2ZeUud/0qebNrhOXGGwb99Nebu2gmiHLqO6aFjIer927UVLd3bri7y+2EwRJOjK5E
rbDLHKqP2pzZ7pmltScoS0keooZPL7xhBM2qXEheIjdLv0mSGfAuRYrqxC+oZYOoxJOCrBLx5PCZ
HvEBnKJEjmptDG3KwKoNs9SbG3AvZ3X61bjNrKavIzn2mbgIJl8ipTRuleqbxJtwdazKaDCrSBw4
23HR6NYujzJNrHg4EJC4CG+69j4kT32uJZ4jnAUlBE3rbdhNP/rRI5cle9Osp/MuYKAut1NWCPqL
NM644a2P458CfbYaKmeNLplOYpMttqsatahfoIHpz8VCwknlTpNLSxqVx9+qWFkJawK+Fi/3oK5W
DAS/0gBW8KcGVmVq4WYRtF2VHdhUuNk6oSTexCS+vWZxpoMiLGrv+ycpDEButjPrkTY0+ftQC8lh
tppOOIKOrm2ZLg2Aj0bkny8WBeysLrzaimE+csazE1QYP177rKcKL40hgd3tT3faytz//fNaJHwM
FYo0dLxWPjHyTH70ZJQVFK9enuZw7+JCuk9Atex45cM1gNrx/dhaaYiiUAxCMTNaA6Dl6ctA36Gw
7dc/GAgKB/l/pqKwXrKw9nppfRKOZUxZbMcdvZgoDyzxaZTffzdz8YBb8Xwf3cPYe72NB6xRepxx
1xfrGi3I2Jpo1snecWVwJqA5ILNbFsGKobZyAvUQ3075Dfd9dZVAvbXUbspWvobtt2zmPiOJWuy0
4moHz76122/ucE6nOm+cUaKJL+xKVQjrJYM1LFP7uMGwvzHCpqR2X0a03ks/xuYzmvphI6mOhG9W
eUYJUlqS6BJM99n/NpCwmrXvk7dw87ySiejLhXSKYAvbT2G2KSowc3Kp1Mu+IpCD42GCKeCXJkgp
q9/qDJOnlgu+8R1lII5hXQvbDeOi9zJnlbKF6T6I2rMhZchkLR18k+53szjxvH3XegtQYGL/p3fN
DVtdo2QB3CvHtTqFwf5PQwzM4nMSUex9XHG2cKUKS94NmAV+vRP8fQZO9jLY3N2HfwjtTu6SRLTn
2Irzo/BJsL50fnIojsY1Qjpdlze6Wp5iCrvHKF/H9qMsm8EKCkA00Ai/8lTM9powOJNtcHKqQ4up
IoSAxNlmzzLfSzh0iK0zt0PV6d18WnU7wIUvOg8ex7y3kO7ASpDuJ6QNnmkzQT0al1wzLfZck+50
YCN7q751tKeTj2/asJ1lkf1puq1xZTQzXBlTdEwaYnzAMyOUZ5cjzorOfgNm4X/LB9t2oSxtyQ4u
JeMrIh96ro7JOz7wnozS8+sdrMOgB/DAB7kOFJGVDBqOoCCgWL05xjn9v5MfyxsWs4siGKnB59PC
HC2dr9X74WOKdhESpkemMH/WGCmumDGTRCOfBtWR0Yoq9X2XnlqaC51Plk/Gq8Cn/zh/8RauugV+
1QX9fQJENiH0qQ/y6LtTbEj3bV3dQgNbSKsKHF241ENJeNRM5jtxmfvyXRR3M3a4dJkp1cYkIw0o
GQROdqUM1Fk/znBZI7fzeyfPodeAwTm8cCxwVajazgDpSRiLHfUKVzUoG0hYzYlP5dlCzNRy1HDc
1CZAJCa+UF8EJDW9FwRQW3L2YKKJUwjwfVLEa4WNHgHreL9KMxVHR6wtjrl+aQUJTp8Z6FC2AVQ/
vjFfVZwThwP/bjFvL5AhaHRnYv+A2Gb2UOO/XiANSrxcufeDru6907YPe/XBcud7EasVWDIPRXrN
MSZaaqN9sYl1TzvmhvK4yW0Eki8INDU0eUtTefX82lGCT8aqcWS8ulwUJzwR5I6xeqFXjnoTkIob
WfnBL8rI98nT3kZsCS0T7TOqeCZIOScdhDRYKmFefrVQAUlrOuJRPuI7Zr1Zv55J9YIKFpeVUNuG
t/fPTG8WY+k+G37vIk/NQZ2hwMDvETxXLrc/+yhZ1MJAwAcuGkkWMDj/l/rO8TGzpO63QrFAHV4j
iizq3blYM200OIjSlKZA4dsUZ7Ktvy1l7Zzi2lj5ah6MBrinlYXZInFqXimrKOH2ffEkEH8z2toa
9N/sm2q3fwCjYstmZgzYcCAswLnZquTH45wfgGvx2Y7+m6ZSVSq7MVi1l3dVMrsfL8vNcYnv3HX1
Rohnk//cGrlHXImoiI+O7MFQhymKt4b4veU7vEjLbSpJu8RXDhbeIt8NW3RrZIHB3emg1OzNEC40
heGb7ozKJdZxBTbaNRjyetqk6yTZmTjWFCVMSBHENSlhRtNBksgUXMvzAMiD27W52Ycqcv570gJq
+XZlKZ1ksxX4dgSJOVXDsFSe86xYMTXgihS4XzI07lycrrQ56nYiutPejGBjNjitwT9wo71olObJ
Dl/dVaA2t4Y0HGxd0NACRBtfNcufe5IPgAz0ZteJBqLyx9+V/R6Fxg8yFF33ejV3BKBk1FtBEXM5
r2JkuYRldLyTJI/+ZLGYeu+oG3Ihpd0Qa9ozzQ/TVxVa78Jed20Pkx1UJ8k5BoekeCehjf/A/dBk
F5deZO3nCDrkfqyjDk+lspVn5xVk8WoRVzkBfQPGdjcpE+R08kaaMFCohF1g510gvhDCYfc+T9cv
dpWsV5U2q2xu9J5HMjZB4W7oegk+ViQO5sJI/o1ttQk1ut7V+0cnqXk7iaEtDvfoSY2y2DV7bPHi
QiDopgzx/xpTq9/VIJaVI3sErMvA23HlMgBGUntFjhtw1LxL0ykc44VLQyjfCeNBPk0t6S9lFDPn
UEBC5PcN7NBDCs9K1GY+eiHLyuDLC5fPLy+jRF+1PgZ182EEfQhpSOKkTXziijzOdjxJCC35VmRD
AcfQ1HkEEoN/jtWS6UuSxcB2D8vquz54yUF1+pWuVdxmWB8jQhqGzo1PJtJUkkslu7W+Ybz+tLaR
pk6W/46+jSlzlouTlL54ZqA5LIvrKW7gh/bmjAezXGQEGTTnPtpC4Fa6JCpElKWvwZAOCliC2FnL
7RVGZuf8LdF8pOn7qc8LcILu9FUqPg/3ZCZsmgtVyxbBbovI8I07usMZ65WjKx4H67FwDvZpl0K4
mm0NWngUx5THzg14j2p3mIcxToLgxyADBz1moR7VTHAPulNddlLw7S+oekvnvGOs39Oxf3uOv/ct
F5awA6PH0b9FueAonvhG+Vh9epngPdGCpfprvLkg5E8rwWh07alN1zVJiVW49oZx2sca8y+kODBe
f+CkC+ROIh+n5zYbgD+7AHlFv3CWrUdUe/q6dzJNHQ+6QjhdQRP4NWSai7CvRe5NNg0oXAB4pcby
AfvjMWy61Iwgey+ei3qRPQuKjVK65QZfhobIofNgmU2yXTpj3mvm5IWwP3DeCyHztmORqu7KZjYA
m5xhzsvkH0lDf9d3lVo1BYDnjQBe9V7kHJ/IPvmP0EpX1yFf7u3nPObDUeOfuP4UzrW2zfrOHSh7
y2Z/VwkfY5qQgVEALTVLTzGt++oW+5gz9/djNXhCRV7NzT7r2QNgu0L992OQKL+4BVANnpmMMVgW
ONMWX/Ys2auexqcT2BlLekhnaSB9oFtqNmW1JCT3yAuuVRvGzKnyKFyZcg+phthUv2NPVLrxuSwi
/NuxNJOAtG+Awx6jlgF9Eg0gyl04F1j4srSw/1cLgmNFXD2CU9u3rnEkjPNzyoU2Oiq1nWdK3Iua
mhv9SJKxgWW5ELP2S/eGe2ukqEVhaU034PluJYBZPyOLzWw9DrskApPythhR97yRs8406TLhFeua
JGal1f7MTTUe8kZf9LzTSgrxQQjiEsCoHpEOzS2RLmF35adhuOTZOeo3LKCo5RE4WMTatb7LUwb7
ONjAaWRduXm+pk9Ou/wrKLPjIJncETripbNt39RjVrzbCrqYplB0F3+8na6Iqz/cUSRn2ZrAVssh
c9UsbWeZBz8jtOyqf5WNRzi3C0xTxVacZ43VTJndHEfBd5tq8GjFlkpI1oyRu/+1e6mVuKjCcGCb
aGYw2lTJ5qK0N54w4X2CiJr0lUwbZcDlcwOHqR1ivSYtdrTev9Xv9j6sJN6+av0erRj7+M9hVTa1
bP8y+eXaXTop9NvYM+8KtJuZLNbfgDn6Y2H1oxO6Rp89wBbBJoJVWC2nHI6IbxiStJFYgdX8CVK1
ivfDGwTKbbOxndPoCG1bK8lwTIdn2ms22cGJYXJ1zwO8u69KT7Wy1e5t5sk66ZlkPkZMx0hftKhm
c3B5z/hzFfNN0jdt9XkWJfXgpIGSph265jCw24BBmI0pdtt9Cb1l/jcDYYe0mxXnlaufX+OLTkJ8
U9k3pSz7fBh80f37GxyE52mbkw0tSBm8hccT5+9NWET/RyNZXQYADB6kk9eEdGWidPdB21N7nvJe
z9bS+IBSVFHhhu8cU64lb0gmRPs2b/tSsKP6ZbIYLB0FGiLu7GhCJtKPx7SqLBNz+BErWTycYM9J
fYv9SnYefceqiWCss/98oxWh3WbW+ikhmo/+vE3TWYxWodl3YMx0JF9f22LnspDeB3z6nGuDI6Ry
uC12vmR2whI8zkxiZmGYtT7pj9LGPt4jRpElgep158DMLT8ltdmjp3lrJxioRevdUwe1jakO5BuR
r11arQTa9/M4VT+Zvk8E8rd4p4YbbRU7FM8L9P/QJdvmeWW0Av3PfydkKD1YGtKYuCkyruWjcn0E
5FVUw+Zfj6MLdkYsaaLtXpwX7UIQwbwHrmoCwZBSi2GEARzqM3OkjUBvzdxosGVHCz2RLvEJJxt6
59i6YwyVm5obmhqT9rwN6Eo8BUVV6jDu8q7JLyn9JH4wEjeLolBGko8DVKkE79XdwXunRf5/JU2h
CHB3KGvPVMDhEe+GHUo+WwzF7Noe/bbVSEpp5e2KN5QMovAjPBqTQmbAisKj4thsYc4kwIpTg+lS
LG0ahczfWpuYF4BpXqzqjvBy3h7SP8R9ebpNQOJcLU4h8stP3jqxcbHVN+/rKHeB3nsj7fwgtrUt
VvP6TgfHTE4UZgLGFQJAgYVl9Gfg8Xu8K4/HjHT10/9h4UewkeIflXzvc4AEt9/eqy2v7moR/tWT
IIU+BCFGaXNXjqmTfkXP7wiw8hv0AjemOK18GsD0F+LCVFKAYziRAXfgavmFan+2M+sIEcUHaKA5
dPcYqELcOfrU44PIe/jxVMvDRIPHSyUkVCEqhwVvJb8Hf3o2y0K0QS0xDokwCkdLpW7CD8EuoWKy
uvwVWILuIb+BWXBvtJSulX/BKf+LkG/o8adSzfm20c8kCEmGMZkRV/02Wq5jqNRnr/ZlIPPagL1J
OKnsJu6WTxa4gafQ1A8XpcEZTYBzWGeJhD6TO4gL2J+aF8N3yozkK0ByrbAxx7zMR6QxbWbkGQH8
7+KqoKsAaQWZJZyHO/IFmH0vrJinRMB9h/kBw71YidJsEzbTUkWiGzgx9D2BJv8J017y3S5G8wvh
gVyQaleikf7pUbJ5GYJMVsEU4/GY0c5pU4VZ7xPCkF0NmSBm6VhMz/YF9vtIfh9Ts0fanRAaDlk6
ek8Qoh/4SxkZLG4H7dT4ZFv8T6/YzBtpE4sGvlvonC1WkElbVHkc5heXd2VaXCHbLRa/qJWk6XVu
/og35ECeaRdWg7towA9AlrVhYitI0fdRH5MEMSgJGWDk8/fCU5BSCDX4W5ZIGtXYJR+83mPAxRH9
ql4FMVr00ju4Ee1/jzfBRvk1xIo+BobGEBNKHSkhoTNmNaTnM7GtESNKcZqEEau3V+n46j5Sp/BP
Jd5j4/7AgHvd9pZX+ge2qzcqJIeEmEpgNje1EUK+jB/qF3WyoRMN8u3/9Hbz6bC6paVxXu3Zf0xH
XZeZAQszPhN8PhiTJQV6WrZnEP9jtLqqm6UCJUlyhNBD+JhDIeWbDGFhgu4tyvc1YDtRx+/7FNLe
jSTvKV63xPrQeOCnNqF4zc/2lvuVzdjolM/UGQgx901cjjJHxjiTVsg+CZ5gSsXhk+3MTzKJlSME
bnZ+3EGqIJWCNFRWBD87WowK24aPDNAT64khJOEEErnX6HY0ULumzxtNErcz7OKaAt33+GfYI11O
MrP1E9gpRJBXYDa5M+bChvVS4rvHDokIpjpWOqGlAiNMdJXSpsiihB3ePeF0Je2TuxdOmQzA8wHy
yJuFokPFPdE7GewEAekaoD6xRmt07NejsMHOj2jr8i15NzT2Ri/IJxfy00IUYa0hvAlydyHbduj0
TgqSB4kAG4LbVz1LPp9ks2op4Hei346jz61kMo/Z/fyClZC1jOrHnkTpinqwI6IBTbD/fw412Lme
VuwGChxFWZVvskoRpJOmZYNy/omBNncBY3JKeAosmwmiVb1qd7g02ZLCMaLcj1ghtOtwdrwis+qr
3oA21x7kOqr6NFV2Z80UtrUNuTAyCJG/4rxsqws5OisHBQLtzMR4SAEzZ/WYszS3YmoRnSt0UPKL
41aaBwJI57XwrvMD3uGnllVpL9aH57sdOfQEfoslylp28uxqkpO9TNcVGwbv17SIz02dqZz4gnih
iCh1cqeOrUtcbmEEnKL4o863KgpkOaIiKOvAqTaYhB/331pogLKah8saI+DKtCz1SjNmM1uqaa+1
MYddt7W+xO1m0blnECO6wMDSG4dH9BRJdDpIMjJCgoVo12Aa7PfzQw0Iyw9TykLP3SRry9dbe4Cw
iy4olXjKFHC7SywmWG0mPNqoYOVgn4kqjQhbbOnzjkgxR/5rpWSmKRGzCmOaZr+Em+FjQ3ZsyykV
v9o1VRh3BJwQOABgRGylm7iefz30FyHiklIvBFOrihin1MfNcvfhWR4/QktZEIL2ZQn3v7bb0inv
BBHTYWH3lnM7vpVGhEnskIl85xyTZr2LdO0D31BekA/I3e3PB5OnsuHk35K3uNvYiE6zp8TgFqgl
AkZOB9GJUZ01hTY8iDUtIPXYtdZssDAJlhl6EOGdHSxh7dczQQcKUQZjdudI8zSDpBG0h+qGAHgL
S9QufS253kqsESAa1TlIzFgg8cQuFyTxykZPthddPbILxcth7SKM+0Gi/gT6r3iXI2cH6ivaKAwn
VR06rD+ErKStpDqjcEPi7D1pTCkNPpgDSZHOkRD9mFmHIAsSeEY4pIlXKDtkYXa3DIYp7oq+8z0p
VNzaCzuqbQba0YfD+hraCiHeAvLl+wojnSiO5Ejng+/0M/Glj0nvUzXA4mPgLZMCZu5n8yY5xCKu
l7tfOW52DfnlnJ5d3ZwRmcUyo3jBOjp9y2iVeNRQYsdEWPXJ7mzoB7TXqlp2QUsh2W1IH8TA9PeI
++IOslUJM42FXBZIog9YNiWF7sJBJ3sWdISHfhaYFMjBhnfgVu48IEjl7HYaUu8XhwkHclHKKwZU
rJ1bMMJcmCYgmqyofRHqXKqQe5daVmTH73ib5EXXH/JUke5Wp51x5VTz9GWMx6DBpvvbrtVYL+29
lnOX3Ik4qLLObjd27+N1WtWnFfn/6yTl+3NZiQ6UtxpxWKt9bghHiJCAzYjozaYviapU0sCA6kaU
f+hSXjtk5EZpJW2U7hX3eViwBZMMPpaoJqp5CbXqiZQhYoLEkq+aX1ntQY8Ds+dh/dZPDKIMfbeZ
DFLWpvGimS/lCIIh5e9k5AjzbkBES4fuSvjmgpfKTjCsZGbNZmSwSsvESUaMsykvq51FSZ8jvE9a
0CE3GpzqjzRdpEJxzlsVUXwlcXrh7rcyHwJJKHxZQ8vCyKoeNiqkoFM0cbbmgAXHek+RDHp8SK5H
0mqmjO+NOhevJFCdU86hV0SJSIE8dsiIYqaoRuYDaJBlyvdHRYio84gjlRaHNjTOa5QOrGxSQt8t
31XuI4RibvHyWxPe5ekfALli6flF13C/OO3yqfvBVy1ZLhdAWtTFRoX9XjHkMRuBNr/2qgc8QA8o
e3C2j0o9u0EPrCp0MzMzo7bswJoVjhhbGL1eWuUlx5taBlnOkMoHdOS/y8lViAJrP58QmFzOIkr5
VYaCvJOnDb18uvBj08nztTjY+syu7uj5eD7d/UsyDVjiPtFrf/o10erEviVp6dzDsL9B5l91eeHY
5WRTQaE5WwRTymeZiKoj7fKJMdY65ZRagCmzJ73E2SwFbISaRXxsYmRg07BvF/RfY9e4j0lQ+KyB
vnvFPZnGwjwqdooU/HoJCnIRGlPumKREJQ0Hoo30xVHbakFV2XBYWxAQlsFBlOVoJ119q/mvl4xe
suVfHFmn3uZxTn8VL7+VbJN2/FcruZdUApMP5Gi9Jxie+e8DxgwJ7FzUFyTw5cNGACvx7NHAo9zd
fV3PoxmMBjrhkjq/OjA+UvrCQYwvABLY5EfXgmLiINy0ykZGyMQDzB9s55Lbdzi9iI5TPpKniBGR
bXJGEHdUjsAGpIDX6blD3ntT8R2E6bR2ouNxry8aHcFiXBGuYvFqRpjsbvUrr/vXmt3YBbVv9AHv
xF+1y0y5Xb7spm3LgJz538MQ7XLfIbPnQDgZieVNniF7+UwSuCy1UzIkVuFZf2UKeJZptKwiHaor
6/9YbtUVX82S5A+cfjZPqi3HRa90qH39cQg5ytKXVk960oGw6hSaAWemFV4H6gXayqgU9QMIA06q
8Vk6hWjENhwVTkZaVe3/tHtgzfFomcGwu1GYcNoRpKfm57Zqf4gkm4dUa+4NzTOSy6oL/tAkmTUd
t7eb8in2zYBYd5qSDsHyOKKSjMfqtvY1ze2CHtIqClkYfRZOsAKXatxrgEVKz44af1y7tCvXGP1Q
Lj4dVohFR3/KTpPZ7yafoSyQDpnC6y6V8XrffVvW5qnu3npuvt4Wl5OHalYmT/lRTAydqe9tTVWK
jN2a9PoMnibfjvfbh1lkg3kMwlXlcPS7/BN9jLBfWSKDi/OV9KpUGicvgVbmkvOkKfJkq2A9VldF
uBO6Mjt2HlU+ZQTqpEA9Bl+oCAGHQ92c+VEe8QUAQGEfumK1VieAVRk1k6ASL4ZeWGCwNWR4h9Lp
4Z8Dex7RRTpaqzGv+8guc5+P1z131mJtYlM/kb28HlppFmiQUdZv1B22K4zhMXLRJVHKbHWJ0EiP
UjQhhac+TEPrIRHrgvMHa734SktDIiM7CjjHdi0CXPF6JJdj3oQamiDWqoXXqpKeoQBRDzH8lXgT
GdA+IAKj2nRC6VyRN0n4p6vO8Hv0KHGlHy/3xNgPZ5gAKoBzdnaO6hJ4dk3kRiBu3X+QUDfU4U+G
y3QfLq2v4st15MG/AjEq119mZxQ4sR4Z9ghxj3oLNpRXqGqhp7Jv7jMlxGcdwKqjEiIBZN4H/qwz
42JdwxjJ/15M4zuIRffZa0S48eB6Ujy1/fBBwqnmevMOM4bMTKqvwgVgXQcfmbASUGSUG8df0QX6
uE8AB43AsLgccljlONqlpPWHCUHyErubv8xA0CFM/awfXNQCRLZb57GMjzGE/WI85slnZewqclPT
xagFCTfgBUOHwWZgHIzLcwt+PW/GUlVxtLQKQi6q7TKEu+7AZjcKNEh6JwRck5nW0IRSGY/CazFU
HB6gxxQUegMXnhTXokdBAg63hQ5XEbsYFu6KsJfNlNvCwhM4eBeVlz0pASsFaynjI75z/qG1chjW
XOGdnvJh4o9Cppub66LsORa1aMQtv4qTzK8aH6+2M4a+IKD73eGm3cgw1QD8l5U0EAcbTgKAEzMl
WnN8KMZGwJT65axuTMJZ0u4rjkzP6Joh88IqVdHnzuRoeELlDgQI8/5J/DS1Wmq0w1GqdsuPYDgC
8cm86R8OFWRy92BBM1ZenMhvrSRZpvk5/qRzOIhFIvbyvowNl8U00ZCXyrX+K+usa9fIn7zw1EUy
6ind8xig5k9t6WjuSqncc45c4qTaLN6/68+9PXlVCE5TVcqi+yTizSQJfh7N9OuhzxnMNc2lEV1x
p6nQ802zVQXgxsGBB5DNI3NJenRxq8T2oYAYwBTIToRAq10w/Ac3d3hBYO8aMzTf8oVCg4KG+hLW
sAqFjQnlJvTHFI5K5Y8xAKFUjG7H+0p8mpwMiLmlMg9BhXbD4vugAir13sWwiMwoSm70lChqe27I
XvdgVt8AelKIq9TEawi74PN7drtAUYgAHkPvJESvPw7fsp06AIeAsS3G4Q49y7WwSf65YPrVYrxN
F4g2b/Y5RF+BEXjpG3D4n8HD8syJX1kVy++bG/Owr5UhAcvqr+1aZyUUhh93NnXJ0dWvYGZAzxgc
ZEyLVKxganPe99Y7dvExHtkaVRc1BsuXb5qWFQ1DboXULJ0BUSYdgUIEHT0hlACcv2c9855yssQL
Qfdo/fJp1mcbSCaIQJWYzdK7V7gDkoLkyB7bzq+2/IQk2Y9LwTHxbfzDj7OhtFnlMN6aTLd0p/QR
Q8MkF4WDMJu3DmxwGykif9OAzgKVCbpVPZPpKFZZbhO5d3jBEvpm80z31EJWS/A9B3nhuluKZP7c
fka5vNLPlJNdSLq1seiXCE9pglXkjipmqxVSR5AckJ+HW/ec1mLyQVhqLVrLk1p6dfH6MVK/eR7h
mTnOTENZE26A0GXxez22vXj3o/Au7g2PCP9OKEUtFAI4PTAPWsep8CCs6Fen50SgE7T1+5CCVmix
o4C5+S1oZqs3ET98kRgnMPnRCJVBqmsLkHf8Sj18+VvXvrWIRzi0s6N+PuK37MSs0LZI1g7dkdLN
HNiZchBf7e2dbScdd3CPbBMUzx+UjdRjP33b70Ym22HmRG4fxfevZDngc4sNDp+Q4FjeACFIUWdA
0LhoeDnB3tdln3roZ6zkzQVzM6r4Xj2RMYAm6OP/PEPtl45+amS54F75oBpB00JH3dsMetCghkNG
g77F5SBNZRlff8+vQPUaguJWH2IrLvqvdlrMWE3/kRibj34NJnsgIKGSjACzDpphQDBcTSp/UAfx
UwBp7FOYvxE5Ip3Ja3ocZiQb22aykDmB5I74iVWaPm1EPuTn6F3FH43ibWpo08LCaAvEpTO355s3
+zqxaldOGBGGTIscrc58bvOvacHrfIJo4hD7K4ZccByNrK+Pr/f4TYxXNLsvBCdmuoLOeXrAxrU4
Ajrwjm3/Sl2u1zSZc+h3N4wEQngN+IMczRKpoVPIVw8eZq9GofMxjEIA4pO4gmlh75rllJa9uaFD
PRLxnXTwuvEYf4e5ZCPrl405HmOU+a0OMFx/aekO7t3h6VygmaLV7Fk/IyaxR/R6oM2dL+QZz/dj
Bmt6/NWZxKwV4g9TbYRRzFePUREv0dhwDQ2XqKemihegr5Eu6SnWfXrDTiPiiRifLhspHgqAAIJk
IVlUAcvyEVjrnSSB/kGsAYw4abqVMNcRofA+coHb/DoNW9fhfD9ddW3B48/gJpDEvbuPSGpPmvYD
kpJzi8pp9kDy9KIf/flwDAsZSmyKaLzn0m3t/MtFZUeIZ3qK/4uiPjTN81qLeLqKtnlD0wXn0DRw
nQMrRQM61SXKN/ZjB8GOLSGUSVuL4Jou6Po7gfpiifv3PcaXQryLfjWMGkCBm3GzPMAMlgDZ2m4v
/9LRKlT40cVkyOrk8dL4YuB7o/c40Z/CgHrAVbzCUrF7jcswyyXdRFI/JOSjdBXjZ6dXwE2tudfq
a43dV+AF0qufNHF5YCVIvfuBOQ7SjvfzfMqXiEYc7jFQuh7b/7uQzxXvNPY8vnumHqOVsBgX4vX0
JDdgTFi+l17HoP1bGISMSjv8MwVRy7vtRuW/poM/12ncCOfYNLVXJ/H5Ez6bnDwl86HTxNbyDB1S
L8rrlPAcGeoGIXsOsTD/okYztBBLad7DvyFhCPU2PFc/qjgHbr5pUb4tSdU4KYAP1ayqLabgwuHA
UwyiFUTkO5czhIz/orPI2SCIF80gOa5BtyiSs4UvWnSkPG0DM/n/bmo+GlSpDg3HdkK4pUagHXzQ
FJBTwyp0MI75aMzATdS/wDuxxGX8pX7XEFLSufl0rRwbM59yRPaHV4GbNzfxy+j47NDHasCupEVr
gxj0iHh5QAMCZER1aD9FqEVc0C5xsuyH9j+9aEpysDl8FozUB6hcxmR27lWkSWmlzVl1MH5+B69c
0fQPHbDD4OJ39UUfMOmhZrUn7ElXZ1srdebztg8oTpblmTequ4A4zqdz4YF4oHrgqm+LKQratq5D
L+hoSEE1nxpt6rbuH8/HVmbLb/oWaLlvwR2Svti76yT/rj+1HmfLyGI5XnbFrhCzYm6Hv5Eb2SeE
u8l0iYC5SiAlRoXR/wCwal35KU67EQv6fLJ8aZdWjJvseheMjIgPsoDsfMm1OFWOQxvqJfg8QYTw
/gcnxIjw4oWQPkZwMC8r35HONrXLl4R+g0DipKcvU8O/c4v9PZG6Z/kSqF7N6nmwI6DU56esA3Pv
fH6U6GTjPYLmciw0hIYUiffxx1V0iOhPwJk+Nr1YB6HAMX7sMnU+RKHYrnN8zHHFXq4Idd9FO6hM
Zd7GwOwA2+KZgQsWDYojEWhCK5f15amNdzju5YLwkSXCxW5JZtK7+DpZj7VqCU981OJrRjJNhon2
iC4oAiAKWwqtsyM9WnERjIzrszGuq+BKl7fuDdrFI6Gc4/5ajjRlyNNcEf2K/Z0BgXj8mt/e70EJ
EoPe8TNxoxzuL/DreS5EBzMGqhidZ2lud5MHgmU9GO4WX6hHO3ESVoxaXXpgmlC777uF48tSA40b
Uxy28vmap34n7+CLRm4WhfWRxup4hIMcYGkKsWXXA9+VUqmrslCK3hh5DjiXZFoBFPBXEbIhc769
6CXcSXyw4vkJPlnE9SKt8AtGjGI+y/UqOhnnFHh45PCBpENPEU6AiB6SxbxkAj1LDyveRYKbLu9l
LTZSVctYs9A4B6BmvvbGNBZZtkwLrTYrzNEERZL9tLB7Spx2ALxsrEgLvMV2DQVM2NnSEI9CdPPb
qDub/X0+czRdD3vnJhWsGH2u60A8igXWQ86eLFi4GsJp+xG6rwj16Un0U3RT4xeX0Dl4PW5JHUZl
q4EojF+SwrCsRW2JOigIykwT9cQaR6Y8PDKonLs51vqz91HOy98mMJYWHgrgeAEckHtXovRjOoc/
iEG+qh3dGzfKKQgCGjl+BQCXgBZ7tXsEXxc96EozF4/lzmurbCTpr3/+vIOETpwXSQg1Szbhq1z2
3zUDzqJWm8RD8dVaLtN/pWA/duaGrMfuel8fUd8gfQucG9q2wm8otAWFRfPisLkXMxsODNm2xPLS
OIFkTjD1emxdxA5Ay460R2wnXHIQZi+LQ9CI5Ekjbkv0XqjIIeVx84PkDN7i8CfEJltaGGfN6QDr
KLJTuthrandZ2OXd0l2lGKbQnaWZfr8k99MLEzmCDfWWWBppZ+y660jWE33+hhAk+ZwE1arAeCTT
fyYlKlRYQV/6WXkBeJ557TYUBy7W38m8XfJiH8/k9qmcx2JiJMezy6RiYmTX08rPUwkWrTetDB/v
Rfepjt1kz9Ja9iA/Q3S4Nd3oeXYHi5uQfvTPjlSggYOTTJS8xnwtjTXASsdkc0fE3U3PufrILOMh
5HWaKAUWBbw5qqA9DRRtchXlyhgrqgbzkSRoHKQA+s22tyKsj6dNGgvmWms9PFL6P8zTkEtuz9LI
pIyZGZfQ69dH1TLtPbhTirdyGw3aOezCGAMtS0/1JjwPhzxCfM10kXPHCaTRuVUAfAxuzJEWjr4M
SSFLfA94XhdtRWrXY+Mf5xZa9ckG/ZeIvmNG9/dbwRQIZxctdPJDXrG1UPuH7JPnGbW/2/1HARfZ
6Kk9HJtNljLWMJws/jBpiYjpz9Ed7UqlbAZr3Hprk1RoqfpuCUcvhHZCQFO2+s4xxyXXMLrB0qIc
K0MsXljbS7dbQW+HaFfsjxhPZV3zepFyC8Uk2Ui3Py9SxoGt/Ftrasg6w4cQdWUjNFCoHvn+Ho1l
DU7lKTL5GrrSgB8htYGI6MiiA2DBgz976LCwj76OUxCYyMAbkr1+bquHlimkroa4A+7AY39q/cgt
rqJA2SAZeACoy0Feh6Wyls9vdtRmQlwpzCfn/dZhfGoAqdgGz3zFRMhrdQCiiDCGppsLeaxzHeip
BgpoMw9jKGH4C17nFT6TJvtZkqbyrO4XZ+DTLHtqanev56DvSgrMWxiJTzl5rXNkN9VGz/ewxqt3
bXsQfm4AusSk1QBPR7pOYYpr/B8R4xNufM78DGPYIdRgyauSQr1IatNndnfSuk3Y0VRNj6QwtTV8
F4XOP5EXvZC0/HrNBqB0gL6KrxHRTDHICp2zgPSiJD/Fvq23nx600BtW60g+WO6YqCxq8ID6CHRl
Nzr0lLKWxxXhhAEwN2sXVS3/5SXS3e2L93tlIpW38pu7UGqjAauWHC60I953Iarz2tWRdERyyAHr
ZutgR5n0GtOImMeA7CtOZ6SP/hOFKpoYygkA9pr/VD2tUW3wgYSs27a9tpD1/qjvryYbMP3DdgtE
dZy7ITRKVETX7hwihoWu1O0EI73NKbV427FMWuXJunQZ4Xq7x7kpV+Eoh/1QyUcGDWYHGXYN3OvY
vgNigexPXGApMdn9u49Zw/yQlD2a5vNyE7Mf303hm2Ug/Yi/vzi4QPDaSKFq85KgJUQOcjQmWrpE
Oafx4XcWgjz9kIScCDlUwucxHMgNrzcCF2FrnYXbvQdy2UpzcLESgxOEL+8sRbrlunpar6JBGUgj
NDchVPXrVsvKVHjCVGkyFZ6Wdb2tirxgS5wPAdX9PetacvnQ19eowrN7Vy13j4SWM9XX5IpROGxc
wgOJpuwXN7EeYsR6YFEdCiahmr2jGaEGh1EjmQ0dMJ2gc+VDw8aJqF6PbFgdqxyYkrp8MIzdJ3YH
4BPvyn3VbrMDDkJu8icjIwszxLA57ETEd6nLp67L5zVZDfk3ZtYbv80Vp7eaxMofOAL0RIJdVC/u
ey95n9JkHnmR0IX5Ymt+AuRhcRZOx+7kRSex1H9vtW9+2jwgKdtwnT/fhJ+AtPhTf8Z+1kOVH/Sq
wbQmInVmuO8qFcKVPZkXIswin/6uHrUc2bLG4tdeft8ROAC7aV9shLM6UitdI0A1kH3hzXkUrCoa
K0LRMMEofC4CD+AlWGvaRS8exjnBL/X9UWN+j9cDq8xd5QmAn7SJMBu3PUVlmb5VMhXSJZhUbAyU
jTR5O44Bc1RfoiIbkGp8j1DoYLW1S2cZ7xlDAnWiv0p1WJcGmasTZXSiU5wawjX7slj88EAzN08u
dTiTZn5tMd35UaA3GWljnV4AYERZhWyHJjIA7S16L+S61B/mfOmTjaOr0ws60LBNMFcaY8JfABgA
k/jUfmQKVwtpiHyGN7Ue2N3Id2jnwF/ngMl01HEq3cZW9TBdWZ+QNf7brMYf5dWP5Tq1IL3okjhm
aNrTzfbZtxMiZ0O1HYX0C0QJmz/nr16uCAc3Z9IsNljKehZNrAzIwZS7lPqfkrJrm3+nhSCswIbk
XQqq5epHQH5qjd93GazUBLA9Z6VSdQb/qESeh99HdaD8GegOqkDr8i4Ya3KlB6gxsgIA7cfBqyw0
+3cRxtHXfhtItNTY6TY8WhGs5P3HdyrmVCsjP/TIZ7XnTLZA+ubcqOW5s8oxyWg83S05SPZZjXOp
pUgD5kTzy3uxsndhV3hGngBo3y9pZL3wbhncjipPRNIAudCKvdZUOTPI8ocy+XLpFCgKy5L0HafN
SF+TInDCPfJVJYL8LknOd3cFgObI6RDXkN209BJltMkrVD5j2isduRic6ijTRyWABGCjFt3B7RBJ
6e9j9ki1w56kNuHuaTWSSLyVO+Fz3Z+cze9UT5safMHBn7EtTVn6oVB799yHU12LrV8Dla8nyeZP
tnIEEzCuc6OqfkPa7uQ0fqatOX8Ee66TQHW+5JTsx6AeiMIcqhXccs8Or0E9xyUsqzvVmeS4b8eE
Z46VzOrg86QCMxA9asc3XY3MuE5RtxlUw3K2flRxT7auxxGVxI5A9bboSChYGNNfqD8dUm2LenCn
sNXSLQoCAcU4Jg8mDuHiXc/NLXAfNnP1TsMiPGDSH2RWkqqqgekh/UKXTYJsvyXmSD1apjcoDukV
H0QQICj24+i9ae31n1XPkCWUuC/OjcphliGc9zp2ydsSgjQxbMZ4J/YRA+oB6jhZpBVdefdNAQEC
XwNU/aonxkAD+GpChW70TzZNsK7fQZ5JpU93IIDDE4izN9yLPjKLjPrVEiMz55nke8hfE4yZgOeu
2YjAkuHOwz78Eohw2ke6U70okoCCgCQKdR/b65DsDaTvsOoIw8cp6ZsFsRVrI7Vy4/c8L50kOjI2
l+HpIMubCUsP+Bruned3f02ijEoCnEYixWSmaCZJtNAwLpJEB+HwuJPa6nytHpQQX58JZSvX7EPz
NZFibF9rdb77EF3rQPQuCGiYqOPSfib++IfbiAfHV8hioSOeHcIcA9bCh1FcNYIZqdOZdeFDTuSi
veUsmk+ogQwQIpLw+ik3NnhIadH8U+lPV0obQ323EeD1LDJSKNThOrjhcfQqRhvLmEtmSmX99xSR
CXIEW9LpKtza0T5VPJxSB7WHJk/hJlFjtNA6jlNRJ1veSHj8HhggD8TWWNztxR2T+DujbP2g8ANC
uVL0eN4si8dIUC4cgpwR6cw+xsfyXb4rBzNoEW7RNnWUK/aykhHpQxgIEDqVFH5AClcK0wX1JgGy
jfqaWkEt3mNNvn9CWs0sPLlBoz9cspy8nAvQNdOdSEpMSmc3XL8+FEkd3CZET8VVc7bO3F5nwYiO
GCerB/j945F0ge9XRrnG17BhSS0XlgVEuvGyZSil3pfTFjyto+ysfS6gElp9dPhlckQPSaFHoJ2p
56KNY/MasetW58zVhB7rJ9WoK7tqKRTC6WEDSBFzmgVRW2vRyW18QRdJ7QsBsJbYx8jW42gtAriF
Ego2W1cO3eO7lBlLGoqEsi89zmyKZHlY6kdGMovL93fuZP1NPFXHia+GikH//510c+knydbnEZTm
W8fB9CJslvlNmHGGMwhUqK2xrHR+wz+jr7Hpq4BVUqb055NyNNIX7L1c5IZESstOhk+R6yR0nso7
E5sDeTQjwyjBg4MS5lh+CimiF8+IuZiECIOGTaCdY6kb4tC+k9nQW3K46AFF3RzuED0cZfyBw+Tj
lGXf5rISzCcXyI7C8oTvzXSeEqKwLMOBGD3Z0vgPfClsubFDYYbTGhUjNQpHk6CsHETMXmayWd2O
XiqV9HyFZmfulS5fLDpoF5yBW7i0TJQn/I66L/J5v9KoIlIzJ79rnVYJsdh8/Lbi0o9tD3Dhlcm+
s5M0GU+JWp2jCOGcWgK+DkTJoKzzj2rQo0X5zwuQwC7Jtd9K80/wwPHrNy4BKHiy18JjBhwCzX9Y
7uA7Gfkx7RR0GJkgOePqMdXBZJbZPPfT4OyfWDBodbt/KdVQuHzn9tmAgcsP2YFf5YW8eMwnzVL0
oSJqDtlmudYBZUQlWPccTTbXdLHasVDHPwkQud12rkXUkkvNJpX8+92shPaTLXroQAtADmHt5+xo
cdq2tvvhpf647+LoWIDxwot7JUvdqcNCDbDqY/s7ORXqH0KD1/lILxKgjv40TTlyr+widQ4nMy3r
m/p9RHQ+rpocJazldw/yZuBJEALiTQILwRBfSG/tS0Uys3VEJNPBOoYlujMycWYcQRi4u8G0tUij
c4jq4lRat2rnNPZ/4iRgjDGaIP0viWR4qVdqbh0b1Zc4b63eSPYQqs47TDHszNkZOyS80DWnSGBQ
cZlmXKUk+TlL0Lp7IgFf93MLixo5eJMJk3x62qVewFcxtlU5mMDl5vNSHOLP9S7vRNlDB3ogUvsL
RrtdWfAsk4uwatDD+gA0Za98kFdgb03YbHRPQZ3KBixuiDvpZKmMBFE3kDpUCa57yZy9gqHHRtsd
HFqcbXPbpZxx7r2VMRlMo9ibhlYmT65I5LX9brplnumaW8HFxdcyP4CkOGoEwNw2zLSgFhYd66wh
hW42iWtWEAVu7B/2LH00PI8LOdNLVeophT+xJhNnpY1K7p9Lbwgffpo3Hj8YOivR9CPI1UbLft7n
nVKp06QkofS4EvaNvdBTT6L0vbUSlHIQnEYxBMDRRvhPl2avy2J1xO3Qm4TFE+fZ30B0bcLVaCQN
n3RnNnNEJcreNG2Z5mx1oaOigFuSg8t1Swgb8nW2Nun9TDV1ir6fsTg9lMof50lZtYAJKWIqD9/h
IARizrXqMoIDngCSFig49Zmz6hAAwx3iAm2yliio/6saz6RRZee6o9elicFX48I3Fz1rdWdvrKnS
pGvfLZw0OMZmW4LX+c2yG5oIj+GS+kknpyrFUJxBxk89oTHkU6ylnM38jnCYd2MTugpUBuuWb8Dw
tkIrpwdVbDPvC8WERWEMluy8prfuyDsZZBpd9AFETKSf3Fzt4T+07dwC97U3w7zu9icjKrEJSBGt
yM1ZSlMQKoUxKt4gEEzfzb5GUoGUh28SfCIGjmZuYUQW+dXxCLzW6sWIb2my13gi1cFSWuw3lWPJ
nMVC2zH979BgJbayHD/S3DlOtpxWP+SLyt8VX8hdLZFca/pFJ1l+WRpQkCb7xF2gBl/qL4hTIl4g
cIsxBnps4q2pzW4KbjVFvy1SCi/lu6ZNqU5qUEkiXQ0AK3DcSGORx56Y/MzxsgyLD10cxilhXqUO
1ivTHJDkbsKvmODaKE5xOwBoOVgrW10a40QhdXkeHhdpcaqZG8RbMmrlefqqFZTd17p2VMBlvBcv
sxDpT+7PQgZ8IARBj8KswXmxXZIQfBvseyjeVgAZx9jjrs4LfYKvDh3QzQpnZblW/seN98H0e+Kf
ID7EFxExkQyZ6X6gWC4U4DVPDR9t8TWm6tUEFQ6PSF6XuQTvn9qtTXMRI5nkt4G+WvuQ6m6OYfLD
k1JMZjCChLCqPO1aQwmkSSPo2yXTGqpEsfkGsel7YlWSRPvYWPjLl5q42hYz0K31RQnbtzXY0YJR
s91AUYX3rMJ7ATkDz/U3q10yYWO4hIQTBondnIlNkPBrJUSdvCPP0iOzWqIXCIxWvsErlqIOqg7T
Ulhuono/yVyhjv3qHabDIRM4ei1GtMoMcOskO0GU/YQTZge+Uh399aYYFuZwu7zMyxit6GlXPs0V
qG/s1W81KQ3rJXKipngsHxXuDQU3cJHFU8XgnII7kQp++6RK8GgoCWqzO26GQ6vGqhTccOjp12j6
AULRfC1cro1kYc4O7n0tNDq3qZcXG1ScBfcVE9abo8hzvF9JKNn/E2dAaeag01cFFbhu6rORt9By
7p2GHOoY+3/HeSqi2P6sygQ51xt82CP6I+5cBob7HDK9kEk0RlAGTv7EpnRfNdMSACFXoSsC7P5P
FbORahb3MRm9wAaaUl4PhnkBLcvicW0Hq/DuNtLWC9xYJQ8sSfIacD9VJf9RNcCa6fBQ06LUE2HC
ww6DMyPe8/JRjOQUolsVMygkRWtUvqfc3E00aYjZ5t0/jWh+gnNyqtmFFEQ+8L4AgiXRe6vWiw+1
fKYsAk38LOo8RmEiaBVGTpsqOsF5Y6BHhW8Q0KgUAIz2Gw/6N6l+wrDHUkYmcuI/WH9FfcJwDlUq
bnNiRYtJYegBmNdv5dvotFoH7bGJ641E6WUejAmegh0WBDWEHlOTqIe1TpIcbU+k4zOE0tBEHt/T
aUqBvQX/hDwyWLEaXq3LRMp0aBNluEDojyKO11TPlUY5f2LzsJA97GHUpXAYpoIihPMgYvDD43DQ
Ei5ld9mhhIHNfh9TEXi6oWApc+oCTVes9VlKJvblmXFNb0s1TRlEskthkSZ5gtdP6ia7/+5VE89C
GwxiQaVNeDMIQIwqR9UJwp3zsHfTfXwzEwZHEHsfQoMYYdxxGIn0UEh74PYwjQPUwYLE6/1r4I+z
R3OwzL0QqqLSoGxahv1snc1pcwZTJpTwTBYc2CWvz+vNP5Y6gyVt9xpyN1ZsTH1SGQkdmpTzKSwQ
xwynChq8YFscuygn51CUZPgUE/sKLAVXXKnhUUkqAsV1owVzMbWS00+IoFeVWFKXP49HngOwN/Jy
9U4xWeFZBbdpClOjEwjRZUtUkSUxkVSohytgyECk5mPidXwhvPX921gkICVLwpbsvRn116ohK+Fv
C2oxnByt0XQbWzow84dS5T2xBtrIl2xUyOJKhq++fe7r1fMqK2xe4859i2vjcsR0TbA1TcDZixDl
xt7WmSKr9kkqEkiTToI7stBlKs309GFNlxwAhjio2rnOJPLUkLezoUla7fkY/ZW2j7yMu3MvVEnt
l2LnmU3ESzQrd4psCwHMMK3ZYMRZCfUNTRgTAqLvXzhQJkhJVeOMe7S/37J6kYFZ/HRceXZ0reY+
3vaBrFOfmSGZvvO1nGVMFQfYw1Utk9As95bgqLxgxJhU8ktEOoqixwBxSmGeUrbWD4LZ895tMS1w
xMCgXVKJJHo3c59CQfL0M4yQs6PlvEVef/9+27ka062O6w9I48imF9w6jPIHsR879DvLozqIk/J0
6QEDVLZkXbv5oJBS3AidEY3Hv0CVUswC/lJeX3yC99aIzLulYZ4dCr9VgDEAfbHn99FprYQ0plGp
EDkIVuYjbCrmo23CzrJK3aX208eU+5ksWXCkupcTKX0mZG0AjsyZfgp3qP8BI8IUrsm8Ak8HfFpV
oORl1p7EucgQ79uFh3kX4WK2J5wHhTmTELorKktJiHFCjwc+esE+t7VK/sudIBjykCOMNwSPPb+8
8JekaoP3zv+FgWpgC3s8tMhTn6sQyTsIvD5vFnqUGXgXT0Km+ofgPvaG2sNlFqQqrnsPIYlxms8x
r8wP2F7xbu/BeIIkFV0AqZbS4GCc6/sa4QqMb/miYRN3KAurLqAoHKoep/Ez20jdlwVsYBJg4vhe
h/GQNOEMWMP3yJXD+fxI92zjVshuPJ6UrzZ32upD+x5e71aHOOo6QFImMFMQWCW6RrALlR74K5vC
YpriXtbdaElMp4ZCS5QoDi3XGkWVqosdDYU7fc3OhT0ysoIiSOeEBRBWvyU+qQOV0qmyv84/mGJz
xnfaulYA9serpGGrYCip8/iqiX1fT8MQfv7gvSuKB8Sq0NcfxboE6ZqwmqHSK75Q1oM5aAnZ610t
PkYcyGhPvdw07EZtUBbmc9e30bECHWfDA72vjhaWPD1/eztIp0R3EhzKg0RPk9Jf8u4hgPoYf6Bz
SgMsMxqyCk2wvX7Wzm1JVSO1SZXpvTELyzreEdY1kb/9/Hec1IjmPHao4wS3Hy/hmBXTNbe+VKqF
rw70Yr+vVFjD8SBnEiTSiuIbthU7FZ+3iZJvA4AFTVtzyypoweJxAfu+saTHz4nT4LSyzmuSENH8
x03dbLvsupS2wDfGoP91silSSsUEUPjERqv6cSFHybUPPETVLum+lcxRjBgJmkrzhlirvB0maXq+
aza+gckLznwl3Iqq0d4aQETuU4iEVLI7Fv002WDF7eWwRKkCrc2LUToaXa81ln21GufGXYJjTrDH
er3VJ2goKpW1CwEIpD/dz1zWKERi4EXOe25Z21h8EtLiaReX2iLZL2IUjhrtw0dhUkVasHgn+VMn
7vjS+irhwLDt4529X4XDmGXfxEyVQL5kuqq7twvcXmahT+ycracwh00reMj/K06AjdnvJeS1Jslu
lQUvsoSImywDOlXrR+A4j90Sx4vnBHGv6IpbvTePETjNnSjlkgGHeKoy/7wcypLWOyHRDK6v3auX
zc40SXREpP2gMEJ1EITluPxzLcOuxHikOsAZykl2QdrdoCZHcVG/7j92MXE3DZubBc0pmV5g68Nj
sHBh61oTO8ipxseApJOwRkNzS4XEcUiZdPE+/0jPHLLmiyHXeaDzUvkvflaHuy5IZ0380HyksxZs
TSdaO1UD06b91iyHf07IzOzMg2OTaBs/a2JtExdtYRQIGXbu/YeqQFPhaZfBihzEZ9seWkkQ2yBW
4Lm3P316sKks8Uqe8/POeCEYmfVklbVJ24byCx34lcke+FpJnQnOLCRXngw4QBTUGcgnxl9OJnwT
ag39UReM7Njcn/JoNr+/iZp07tydTl9/s42lrTPCi5kV9N2rnMfbgDwJ4Wp07Y6AnEAHXkcl3VY/
mVbgCxGK6L+PYcTBJAJ9CcHORv4b9iwtVVMSvJipB6F3y6m3SHRBc9ZIYWDTD86oX91bDWVxT3eX
DlWD1r/joUGbUE5PxVvhiA7/J3n4rLbjg6/mC9IYrYKuFU+Qi2LIXncFVND4+6mxGm5t+qVON4mB
2hQuC25NHzPsauzzVcU2sDf04m6KUiGB3HpWjw0rx6jVSHYGkbHuy/9AKLY85C/Sxp08WARcxNtV
lcdYS6EwvFBKcQdMHm1MfoWYfu11eIJrNGhBmznuEbPFdOqyMXXmNvdmKpw1j8vwsQp/cG4Zc2o7
7sTWkM2MbqZzvfzHFkZFP0BB/7qnctz3ktpailH5jjJvNgJPRsRA4uHrLQmUnkc1V2an6g4fv6SO
AoEm588Hwl6pk5RCxHEImyTy6ZmdeZaWqxWii0z8faeYOKjq4Ro/xTpn3V2EVPdKBZtlukur/NDh
i4FmvSMbOCsLc86zC230IVqFJIYEgNkrtnkMovAMeX6eq8s+dozYgnW0NCBAgX7T5UnWTVYMAdD9
cQdxTXJx4GYM6DQLdZOmP5OnInOCscEbWVQq60w11GTFrNoUk7iB46SbcexcPCUM1xc9slBlMjH0
czuIxxJ1KDq1X/mgsNrDpuyMEkgCVWIIR5RjBXRsB8Lqbitvs66T6YwffjpWiSGQQBCGO1LTidR2
NJ99mPAVrSDbrvAf8cwvkyRwP97U8BtC9Dz3M6AL4fxSS094xUd5lUdrS8LAlFOK0jXPBAORTkN+
c+SKH6ZPQE0Ju6G82SOptYLMf/D5ImzEpLuCigPsl/SVDiJVEV0/mEzubgJ9JNOTpXCBce8P7Ksb
Lcaie+gep4pyKMynhifDeUSvJQTPXMk48+Dizqv5DTi+6/IJAVyeV89Ve79e0+y9P+OFM4bImgJJ
Ra/0QCL0FA84A0UFGHXyfkWixPz8MNK5rXkjFeaJYX7H6wyCH1RR9ANRG3fKzoRQNQB2h0S2fNvj
saNTXw605pMeFk/TdGSfbx6K5zjhdkAH1ibmeExUTLa5GxI2hRStUbtYeHwBug75W+9hrjt5wO50
U3CRUctnB/5/SZ5cS9hjSJd8YQ1eRif7CnSIIMQBxDLp7rgHwHKEZ9aauXif5T0vGe6T2jnqpSNp
0p7Ow2rN8+RDh0w+0oEh5JdPkkK3HCcKmu9mlQkUdJWYQP5sEJKcyb0FJKLH91GiyqZqRa7dTcIW
bZyzng274faNXwKEdQGTxVVnUIoBMIBJYe5fh+Ay87KyRDupJeny8lYL01XQtN7vIhDFYuKfzNDr
qwJxzzuFLTFaecqndLVDW6wsHa5EqRgtpIJqvPFtOPqU7einEFEF9TBEK+c45tF8IMFnKKC/lDOb
jRBCz8zYn7+Y8jyLRFN5YAI/13zpkomH0ljpZbUjlNC8o4jN3VCj5rmIaDE/WNXqw3wcMRI8ouUQ
/SE0b0+3fiE2LqHhsooG8G4P1CQfZxnA5U5uItsFa5uwhEw/NIABhdQsnwf26JuMQWpfGsdDXKsA
KB+jAPD/+t6l6yvEax9P+wKaY47mutqBf3J23PC94OWi+W8FaCRmYV+r8uMJ2hxNtO8R0bRy8Ub1
/DHrUcp7gO9DzNQBVqUOY8w1cjrY/PcAHRJCoWaIdfc9G56HH/9M72Am4uGQZuAx2WBuEqdRc1tc
HLEExHN7VodM0TyC9QfIdXDfNAoQlbKs/XehtXu2Ri9BBXThjaSTc14GdXBVC6sxXDmcth8SnQfr
8H2/dJlamwUnIsJu3GzKU9sbxpvSqPCKFBIF5ekgVnKTeKUSAtlee1XAI7lZUwgypghKHlHK54Or
KAmTg1QPrnsTBwYT69xPL4nnN2s7Ihlvr36QgwMvcExJkKYCvp/wh00wBWDTUxJpVQIIwlD+QbOa
SV/9TjufHVGdhw2+PM1/cdUjgwtTNA1QVtnNZUP2PsPNJk82rBNLewurGbg7DspeKhedJ6G1ZIjH
2KH2LZyFAV98VDWXfGRTC77pyipHINMlj+zkDErWAw1WxUVKrNwV8k/4ukl4VZu0OohQ++I/3mn0
o9ss7LW/l2SsG4ePsMmGGs4ZUHix+rZBUaAeI2UeqZ6nOgIUpUelKXdSiHRdIrlepye3AU67JuhX
SW2IRqQSl5Y68/J8LThcryX251EOz/XG+m85bCei8R3rD1UmQgBr2Emy+2ilWG6GmYlb3yPCCnnU
XpL6DC5P3UzbZE8hFQRaTmLnGex1MzPGGKoY5SrKaLm/2MD9l+7yscKOQ9zx5PCioR8TXOYyiQYp
RW3V8o7vYfMw0VkbmatdQ97wEMvzJoCZ0KYKWsRgFhF8Qag+mV6x/3G7yZbj1veMpBLFchDhyU8a
zUzl22ui3a2BMQFdeg041z4KzLXL5N2ierI8eLyY6IzPkTLSXQ3LCc40895LVjhLxAunwAwpODZo
Y9DeLZmKeZQT/Asb+5k2Yv0LOaDPCPaA5QaS8UR/WTKFGw6ARTHfL8oYEXXqHmE78TLRDF50o4kG
SN8dLotgloUwW5xJ5711TCzjhlrBGGauFZq7NQes6ovkoDbI5BdOHZo1GasY38l/vEqv6mDOKhtl
PoZG4CtgqWgn3PeQxImwvZPwrDw2ixOmxRBJKNGbAxAzQO8sbmxNhwU0NEgUfWmWSQxx0JX2dUNQ
OvWXiG6jswVKKa5yK9ikGkKXN3pETsHSbSoroDytFlbkj0pT58GPFs2QpJgZ3bWrqlruxgAUDpj8
Vs49rQnRwn9E/Gz/KbpEbXXaEj+MK58WnqcRt6CrbtLoTHl+wh1QBribm5n+7LIWB5HrjHBNKfTa
nFw9jDxqAXfl2TDKb8Mtq2JOcKbjvBZK5c3vy3zLhb95nmB7lpjeBKCkxkcG5p6sbiE1c3Serms7
d+n/fmGcb6RVrkudu87lGBF5lBzGfCKUTd6ps2frEzwZOl0LWq7nyBm/ie2WwW1N/FDCE5WKBq3K
bXHwTxz7hgPIEfJXNTibVEse80ipB2+Bc/p0CJa2ts0TPyN/WJ6nI80EZ+m9ATyVIhlqCT4MVsy8
MQeBIi1RsAkF4LEnG3yVeQI0/k6CKy173v8os9WIFVNCk7aUwF3tY64fUrY3Iw0C6c3jT7vcDXvs
zRA7CeQ+RncuvrEm9gj5chsxVhfx6HgWbLn6/euVtyVQwLa5xpq4DE3Mg0V1qiBkM6v5IURhrj4m
7tOHYxY1v/kbvDh4+R2CouS4TPQQ6ZFEvePBpqT/XfmsreDOVrcg5Ip3H4NUHB7HS4wpfCk0VgE+
9Z9QrojTte0F5O+JviysqE/JCXmamJZ5uuoUjR3zbR41SQOHT5VVqZc1XiQ59RgS5PRFNSIGuFr1
pnrCJklfcfreRQY8rGV3YJEPFCIxmdgbUs8/gXHEQ18ezDPgVTxBXefDrYYJwieoSDniAkeZP/F/
T9W7D+c24jtfxiZSJ070yl79KaXQYEH7Pytti+W5sY9enS3fzY2onr0/+7Ym1D0r8LL+LsUUhYKR
Y8zB6Br8laZ+9d37c2WhVzeZpdvPJtwFzXstGokD74TZPME1I9/9xIGRyTH+zXMTdsuBWs/MFOro
4zJ4fAwYxuo19CFmtneoRg7JRyaVAw5jvcPhrI75PkznyczosfExeEpxdPjwe+xclebbviFmPBcg
v1y9+ecmZ6mb5pP03CUt80x++wpj2NkcM8cbkTiF5GsNFeK6afg9VsW4LhPa8odto6yYV7hpgWL7
AgCaO7kKABIDW6mBL9e1p8z9uhp1d/8PGkIjCGAyEpvnyz2WMNFS/f+wBZzSiP8t1gpGwNnQZllS
e+011W6g3iWwhHB9kbsz/Iq5QbOpJZUyXV63uM+mbJbMUflCRNV7eQsmp/7/J2us7ACtn0Lq6sJn
q4w1kQQY2X5Mu+W0A98WYAh8xil83iabTQM1LQPuOnmMMsBVr+wVUtgQA4OoooE+AvjpVgrbwkCM
rZ18pSNGoB0wjDyyB3bEXgVwxNvn+KY0Rglg+JtufbV9jUpVuKDgW0SRfOFOBa1uSNGgG0+ET6K1
6tcPKnuLU/QpwK5bsM0cOkhX5DMtlTATmpUCqL6Of5huNExOBGVNdfpDdY4Ug8mOh9K71MdqhvkB
pYOQPmzIAwdZW5drrptmV6pO5qq8ACDXjujcvfH0VKLeKybV7O0pDyrZad92XGzGSUlkCCXsRU/r
OGbXHCOxIrOtxI6BV0zYPSu2R5xayB1agc0ZStgX2QMbOzbJ2UsIbL99iPd+Gh86mFFHJbGYJx4R
5HjaEjNLttxt7nDzuLn80GCQRdpOY4lQVjuPBE/ARHzR5VuBaN1MKXz3CT/c+Xr4zikm1T5iiCuP
vrt1aLi/khO3tMlZ2/93HFa31A99p/0wD0+9u6z++WCSQWXnAxBortt0fO7B+7R31/977uk5j49T
gNXu4UwydYIkR/kIBYU6cLEewAioSs0rh18PuWBaiWsbMS2OiVm0RO+iiLZ/6gVy/d76IvAP6iCd
x9KwMvl8drXP9kRW3meAQfxOfXQgYABx5/RN1/daXcbS/wTbR4bmCAKZMHnDL9TwakTXKXmHJ3iJ
bUB8AVGxGAO7HbF8vzeDth38JWwOcymn4VJ3io8++gZ7Zron6jwwqc1axHL/qngad/Mg0UGPa4CA
sW49OxG9sO8lAZWPi+zKvEK8Ebu+Joueq9uIHaDZVJcV0QadwhnBxQ24OsEkDQezbWb507YSpsVS
rCBo5ku1ePlEuTRwregxo0Z9sRCymJJGel7mUq3NW21kFOhs4+/C2d9iSAtcllJuGFkI5bRNTVj/
UNMjfYA688af5cnxDzxFp3evZLqtM7mXFlRmLx5nnbrhyRBuW7k+aw/iSRJQp7lYPBLX7ghnkbuP
1VLX11MN4osglEoP/5ZSwK6Hc7uVRjA0mxZyQHNDEytvhdk3hsrfPlep8XS30wvkRo98TGexF9pp
R0qj1qfLGaphuxXtFYT/zbqnX3OEuP1QRwUh8Tkcu3qwru/20KpWZoxvPmJPucV8FZEZXzbtj+FE
BxCdPQwqutBmUdkSpaKlHzqd/Xj9IIWef1qmHSHEFIehI8qMvoS8jt0uTApDHPX4OidUo7gaqbe5
sfsWgPuoUsrGTHY8nu3g66XmKfM9/eulTrUfJvIe2fLLiQAKmr6on+I8tOqteyDI7Rmo7Lvrl+YK
bhJ4kSoYk0JqbqAL2zDsTkJW954TrvmnBlUqzlUBh3e2D/cb1XUdgta2jeaLLpLUPv4IL3LKzZ9F
C55f6QcRmu2ONIl3bzVcqdCRgXBq8Q9bf02UYZT+hygodRGOx9DljMgDlWoyGKM1D5jpcxsT2gwU
6W8Y7PIndUIdGoRWQZYeFPRYHbVn75+jELC1SWyT70CK+vr0p5Hkwo2diFdD+Gdv7L7PAtnLfE95
Q6Ay+GTTNgpMO2mL6ZtxL8uukRPE9UP2LwlhDZwflNoGQtmlVYg0ElWqZJlu0Z8LxBa9Li1eIG5Q
trZE9lWRMNXy58a1lRh/fzq8h9KR1ylCiMKqaLdOHiWudcqNN3K/go6zxrs8sUfpAMna9gEUYVLd
zj57Mt1jR+YLC2hxS5r0HcK+Ik4YHU8TNzwLX5dFS1dMF4gSWYhj6s/4yaeT6L5JgLxdAk3vfCCE
oFBT8FbYpcgGG360y9YWhDHA2+Q5i4ReU+2/SZRnBjEpgbvSPL0TWLMgP8toXR4aPHwJeh9DR9kg
iREdNhGAlGJnsaUeW1B/j5HiLN69ReZXsFDO2jy55OIE+2juLRT/P0fRGrjzXEdgf/04tg+2+4ht
9NI4Hd9qiNJ6tTI2arkJGnvIp5xpbHF40cpdFrAAjeOXBpcaFEVJAIqoQDkcHEsIg7cClM7rntN7
Dp16BNqWmz5tqxXDwrBQLOVzifpf7C+6yFj8czQK2HwifUQQSeRRHjrnxtS2+sZP16kkGgW47T8V
Vk+z0sGbhnPmyifZYIWSvXVuCCMTZUAfWRYcEZrB9Df3Lu3O36MfnHRt1cQk+x18zbP/9CpXvjcP
HIZRR3cV0RfesY4fEzhRXh+AlrDypsztCjzC7wPEQbfnjWS/V0rGYQiCcypgfj/CJsbfLzT65BDl
nATDUnC2lCAatmMJ8fJw+S3rCelyOzjV3ljbON+UiK2RHNBW/uIQfrzpM5iuC1RokdtLjXEO0yqk
y2zuRjJhhlsklfN4afL9rCXdHwINLgofMZrHqCf6FfMNABJkF19Ys/CsnZR8pADuo9aCBeNfsHtD
psHkHuer7acyUDa78yU4fJYtZR0f9Y5c5fAf4MGDwS+PAWPoAXHvbdMYZxktfgJlHUS37SPto3Je
nQK4TD28xkNyMYKhQLpOFwYOBKB+ORmtwId8jrSXNHWV8yFKkWxurh+fMu1ODD5+v9BTrdyG1KBD
XfT58St2haEiV1ktvtWycEn47Lx+gTUYXUMQj46uwNGhhRlyfw+K+IRBwV92Rn8xVaKsApYGGUz4
93Ng6YjMmlSHqU0trsrqiG4kv0aBXyPiHkI1om2C2T1wso/j3+gcZ0T4k/xhd5fbC4kM0SuBfyxm
5CmyVwrvM8kuKiaKpFlA3xLIyzZydBvyHLkKBKRIG87Hiuj9nPWlpDxpQbKoInr7pSkML4lEQfZD
qn4dBSlOLPtCIqnNfLEzAjJCGcb8csCvmUFapD16n30Je4X321rMBnQpQXbVcFCQnHzX4JSrn6Iy
4QxYbdytCmFCCTGWNy2USE8q8YOm3uJ1pN43xBH3x6oL/nOyew+uQu0B7dZiCOHNqlbbt1KWuE0A
w/EU8C4sZf5EmjYzHhb1SEXZK7CDANm2S2KNKH63EB+G8YV33zCREoNdkvf09xBobtdPT7Fq75Uj
l5qd5Z4D/8csifV3N/mJvbSc0tkokLz7EyTC1DGPWhq9FM+2z865bBD5VzuxkzPQIyjm3ONFCk0x
iKeEOAe6DsevK2/dvMTgKFWz+K4BT/j461T9vmHSbusuR9TqCIi7INC/4R6fJqAt0e8M2nK/5Cfi
Y82cqaC0totVHicJ4l9oljFdFc3WzJzbxV4WmT24mqrOKpDB4NevlILRgsaAPe6pqSYHiSAHMp5U
URHoN3CIxGuOC0BnOWgEnsUvpwFrhDWjnLcgZdQWQ5vZBnLI5GYHyeWKyhJtjVxuwo3W6fYvmhQ+
Q16ZdP+fnUBfMnZLRtfNt0aM51xzUObN7VdyRaqZdN0yyaGq+TS4rHQJI9kqRsWUHguGS4VPeUd8
SE+gFYXB3BglqhKjo9y+uCYtHHs8dJNgzz90Jg6IPrfP+kGIvwT5Pfx9uD9yPri8kYMhqusFT2+K
oU79hI3mr1q1DCbBF9IYA3YbwklwTfTiWENQY1R+jYW8mjIIHSq0rdx/ODVb4BcFs5eBi4Eu6kko
NVhAzndBE4pt2M4iT4FFVY7IPNqaSkuLph3DRPH4hIQNJoAnn0Lijut3dHPKdtantW4lC0GMdFHi
ot6z+ZJEE9w1UK1CdT0Gi6bfzlPnfvKfplZ2bzo8gB3x7VnJX5daKiCRq+/28VjPSHanE0k+nFDv
LoJ4oYtXvUFgDBVeZFzu8sOpH8TciMr+i/BugEUMmhqjP1ISItbQnNokuiHpGROmmOnK14aOHykC
ljTh0/VMVPje/4/P3PonC17dakp/JOFcfKZtdJ5cZKFY+xbdzNmTTVb7EjopC/U443FoFlQQHvQB
7Cl9VXGCwT3gYeW2+x9f5jrErXTPHK1DTutcRbBQjXwK1b6fg/BE3BnqB2vV0AKhGTdjmvwF+R2y
x5cwL8aQYLUxE1PWQXdllnuDJ+23zVqCiZF4rHNDl7CPpUCdVtdPVEGuwDqPDuWwZ4jkk8roXUdV
cwuEneko04P+laLYPm2sQPGE6gcCVR+ididvsLeBiIqSGjIhzx59aqvtniB7s/RFtH2cWJi7jb2k
zd+Lc1PutKSulr8rdT4spz7wKy/2PRjynAI5ctV9oft9P8huWJHIYbk5Xht0xC9KYjZG/EXxeNNU
i2XtDWoAacDoE1ux7WO8PpGZaW2eCeb4gBGZij6TPr/UzLS7pr/76fgXMSNDypH3jED/f8HInIGf
q43PJDRgutUZ0lcK5YAM7nwNAQ9ke4WjetjeFqNrTCkkqlqC3LU0A0mBTTYzOkzSgPLJWpDEzkoC
G2zN07VOkkJi3Nde3g+ru+vBFgtVoDZNj/P1+3QAIfM3yibsapmqw3makCFa7L4uyVvcscn3BolI
LgWGJF8NPYI+lu4SoLKwuGmCifnb20lVzxHDe21slP+T+NleTvWsVa/VrLmEV9+BJn9SO+yjUYS4
JMb8ElAeRZs4T37OQJTBeJET5Qlr6k/kJ3wa2eMUW3O63lAZToRicNMdn8y0Uku3q01vmi3V4sP5
xnO19OOel2oOGNItAd/lqrQhg8ujo5eAlnrrzKXZ/yIxukCtzC/extYDBpR4Vbay+6Mv55Nqvp7O
+Ih0E5npLOBOtQtVBdehwxZYlUAHN/48OcnbrGAEb8FBkH18uX/Vns9tXvBzDIW7GGe8F9ghkZfi
29uKfuLjz1F2iiblED2SxmU5rxPFvWOG5/CacvJ1HOUzPrgwJh0m7OC9t+xsrw1S1Ckmwca+/yeG
V6zrsoglCL37qFfGGJT648xsMK/VXlBBT1ZPe9gVohay/imlqLpn3nMhiHyzI4d1n4JyNX/wWgIJ
eobW4ALk9Fp6nQ8D8BYp2NIGs7gNzciu6XSIuQHx3iIcO6wEiEA4ZIoNquJ7ugCHaN+jPcy1QWtf
Bab0LbJRFD+MGGsNlXb3DKVD7WPYL0N6MlCBOjcPVUKxV4nteML5FdB5FVlD5pucv1fpGBE2SSq2
rS5DxBOzL6tyXURIbxzRDcsVCy9E4WCex9/I8LkE0XTA9n/ePhytvg1Ns3EoVXoG5iaMKLfVowaM
reIB2qXvxjUeE6vSI4a36jznDWbZkyCeMo+FFYsEegkgGG1EcoJy1Gw7+qtgN8QL23+CKdBfdncv
yuqG4Bp0AICyozqvwJecw5eUEAgp6ruZ8iBjO7r1KdyP0vITTpnu/dSchglKKo15FWZCK5AtX+OL
Jorbugu+Knajf1ooLDwXIiNZCnUpykWZN7vox9QZ0KgTBKw467MFU+uyyeBeSip8UBtm8Pv5MR+V
ClnhwMoUEWB6MkBP2BGm3hcAUTACpnZUHaI1D6+HmNu13S7c4JYYAjt5muxqYEJG8d0qW7pnXWQe
skL3IGhcK60bu/srUKWZUlPT0ccbAAs8x+Hw+qe1v1XNPuhLhD9q823ZqhR7w2SIpXQLn/GUlFDA
IFawrDeBw7I03V0DuJ9o8Cdgj9SToWtpPWNrdmVgCk2SqaDPwO3Q18ZEuErs0Vu2+YiFhhrocDae
CUd5Db6veBsJfF/3dMtkEurFpseaiO1mC6dq/jgM8vn5iaxbuXPrOnYWbl93kqgOynJ7LIBt2QuA
b1e3zS8DxfPMAX6WOPV1MScs9CcmAxkX2wQl9Lks2kTZ9uJoi0PVoHc+Rk+umvlfDgX/emkPjBZE
YuoalFMzZVlKBawEajqiJt6aDZjY/08vIW8/yBNOJUuMp99BjLbNiqxG8zoDEnBU/Eo/DVgRYys7
L8N159bXewZlMKDW6J4tcUx67/eJDY43WWSEmz3qqGPf7bk/gseajSDgazt9hjy42yE2eliJ9Vwg
DA5YilFHRGyru8J3HnJXS2WnD50NAxZ7LZor+pciV8TDoGex3cWgmwKpRnKmHObJ+zHVRwHIp8XF
rXARKeGPPN7s39DgTsKJErqE4iWiRfZ9S+VI1Iva5KDPvLGhmfyZuQMqsHVPfJ0vHOvcPGDb/bF4
HZJXKeHMFQmPfMg7V0698qYU5VZL0Xp79x6qRWMWqV9gsw9clkbLcyu564idz09GeMtg91PPvYJM
99/W1+Ren9qBJTIctb6DB21UdOY4h/vTatRZsYIC+Q3d7ll17eN+UT3flW7chat1thWb0YmNywHt
e8NyPM6r9jxpuvOx6Kw3zpvhEJ2+r3OB8yvurJ6+//5vHsKeWb5396v0p17W8VpyoW6e/tXuJo3f
zMzVb8g6pSY9+8JYkRhE9MVgHDjSOG5tDOqU+J2Z7nzWtFafSickZlMZGrbs02J+tw//ProEULBo
TzZyJAHevM73EW3JxD+KhnSQIc5bE/8W5m7m+KuGL2TThxKjuAqsLWqNFU2p8/MdPv8RYjm6P1mF
vxyJr+C4phRSetUWhYEy3lTKvBzvFzvX/eS0nZ9fKplxslnR/syY40eXSBdNMNE73xE90IcjPe8O
OM/CUh4LaS7WOJzzYHcfT5QWNJ6w/2ClCTp/nZNXulALYC00HsnFUYM9ej2DgRtu/Oc5zesshoUl
IASkhPJvum1/TvSQbxLiX7a+eNLitkmNmmzQD8r+fuE+Ix1NCaNHKn7SM4FFfBcD7TzWgFDOewje
42g4ozlxEQVXjNOQ2vCGS7ykRVMgokHmmNF3IRVaeD20KsBeKN7Wdo6ydB0tiWmvQKzB1NKMIxEw
WbZs/wIluokNQzhT5phajIcDZNejwNszQSnXS+9LSiXJ6RVxi8lcjeaN+1H+GA71+8CyLUBIvwxR
S2HLhwqu8xMT6d3QLnVY65GZdlfi2rNNBHwrzMSeyhr2HHBymOY92ILCT7rGGhqfVCsjkhcQz0E3
3E2zX9eX+9j586dFMAZa54j0eBaONienkiWJzJ0OjW942SXB+DV3QGEHR+9HaeSN/GupfYAz10yf
O6t7G8KUSXtPiNo81NTTQ7EGduoJzVN+4xlFOkQSqtw17BmnZGDkl32kw+pGnYWZd1jhp1yUNup2
AAfSbW0ll2pjzLBgWPGrEyN8wRKEommiw7GDpWBKQjaeSKh8sBW+Ltb7BRlRqx901YLMODuRWoX8
D9GKr6fq9E1iFaB4wudO2Hv2TqOM6NCtCRFZhHHJvMgpSw9/JLxgGTYB1gusU6PdEWBvyXXFsiuk
XioilAI2ID62JSrnAy0YoQ1oO80/ofZxh9UE5HIq/lQk0K8pemybEi3CJxfJu+RwquB8EZ7x0pQb
HXr5ZKoRZV7+lRP3cVVMA2ya1xAtP9kdei0ORh0BxKlMtfz+gi7oZiWPK05s+5ak8ZL5PQ+PtNJf
hy59eYoKz8oyRDre2ktJcGRsJF757z6hiAqdDZDxvslO/Bsz0KAH7CKCRWgKASIWURtmuVCNM3NM
SOhsa46ScUaAhyzCPgMvEvVggqPX7q0P/XZSWbmAdHggfY7lbfNNQzpIoyPONe0f/x0MKdot6Wxe
CPCcGd7gKC7NLIv3Opekob41mK0YtB1dNYwZ5t7N6syCgcCTXdlz3wYWhBr1BI7jWwlWcRflWhj4
zrClWa/kVeAhlZ5w8jLiXT3ktoINenwbGMwMKtxjDDU+W2HfyLqrHG8KdYoo+ZGFgnrQ4Bn/W3Wv
uRwTZ24wDYR6R0RPzYMg6+KKfn5JQgNN1UK66xnX9xc2sQyoHcuUGwpuGQ4Xigin5ui/lOowWOLb
SGVs8m3V1wdu+hXnvHbbx3eisXf5RmVSkgZsLq1ReAZFhHDp3w46fwPZmrNqIwG/9ysc7AheWA5B
l5DxEfg/9idLCibFPWTkJ8MjsQrABR7bBnQ1q5yS0mX6zHdt11bDQWzm+r7gfES9cwFHKcXWfhvs
h1oAdFfVkSFHfeRTYGIvYsmf2qSKjzPeZ94X3oedTyTxlWJaeIN8WP5OhpUD0nVeBN0ujQch1qY/
J3t0p8Y2kDvxEH/YP8wBMYi86KBoaNsbiU0o0GejYia5dwMum5qISd5wh1rUKrP7N0wIJH/mxflo
bVRCy3mS5+PIYZ9hfX42eDnTeLAAuKNOxIjEfkDV0yQJgBq5Hdq/V3I9HDrhoWA9KFgmSOfJANZa
qNhlgS0d7OSeRycsoUEUPd5DB/oS4kVbj1BMBWZDizBP3KZStaL5iOzB4XooyeUWiydIXo2/K+VB
Um235g2xQMj/M284iUOpQhmH1P88ubssw4CO8Ww0QUXUNSfvDlilbwTnueEbGKE50i9WtWFkOvP/
miLXwnb3YOKdPMX6Up056x4wtHlynUcceddkEHpl+G9dfmeB7znqiNkamnIpVQyRV4jY0ZqLyukl
I0Icfw8PD38gGQCxVAXUAOMD2lKfcA8/xERFI0CaGyE02vgVx9tHmKlIen3ep3ZHgHSSgOWZkPfq
U2G0H1f8JcA9MvcV4F8kzEganx3UWibgN/KHhl/eewX8RcntZ709OCR2XQEFiLDR0vK6eU9XilxU
OSmjcAoL7Cc2OW53Ydwh0jrrXlLKcbBzP5U7+hdMEAzsG/89pSyg4RTR0XQ3hYERpk4kQ5k1/T38
UbKYH25z6INQfuyu+D34+EeV5j5hivOFBgEaY/mifQkLKTF2t240w/Ulc5nNdCHu/lKutsF2JmHb
TifafVGB2GtEuzeCvUIjUPq+uiiCgM0OFi+mk3pfS7vbTmMh51miQ2fgUUs59KvBSdP3cIDVn8dj
ZCySPNU1IesbVYHcvCJQ1JD4fM2pC9HzDcG8hp1db6MfNQ86WFkLx7mIdOnv/fBfB4byRnz3z+Mu
M+EB10tHStHgA9dCIqXEgtmc83iuW1bA8Y8RKy0z3+6QdXFR3woBFl6NWdSOnCu8pm0WJTQmUrIv
T1o3FohcLhYumPWvYEubFhDZHiqPnUhwijPhmBYtX5xldjKmqCvTIVR0oPUeWaDX0hybX2y0CadN
MDpweSTQdUYze2cNcjbMcPhdgp1+DzIEoc6AJOkY+ThAMPD4CkcW1neEJylg4pMeGhn/OZebQFOy
0pUSbDGgBNPnFZFpoIPi6sB+b8lbViI/FBGWe+O70V/koCl9kfk7ahuBE3Ezo4PPk+Jh9Ib3CPJr
E9dEF5bvkysTWkpUCwXUKPKku0dO1SB86rDtVGZaH6G9hCBD7JoSx+Anb1ce22pOkTwGj8fc3Q10
xW+oC8GXlF/l45cxTOrgs9fHirRutPTgFFQp56dr2uOsHZQoWkpBJ2y+yJk5mEufNXe59g4op6ie
4hQFzAd20lg1uJt8DiFZUUdkEv6gmwkP4RUM5w6MVSLxKkxlgUD8Wvhg41bfBGpJUDpckQQUm4cr
fnKugqmTgvP82lci9YYk67shGgGoW2N6nVB7I23EoR3yfDjfl3RFVxSxiXu0iC9SLzYQytl83ECc
EyxYbGG91JK/LpPmERyeKW8s/O1Wj74GhTUHqdiPZYy1rP+5vPBd4vF24V9nTO6y4RBTBzxyE5mR
h9JfpwQnKKS7yEp78U0m+W2IWU47QyVZgtuVR4cvbEyjrZP2BVOpJP5DwdXqLZxuZz3jx2SbWCqQ
XQzWZLgBqo7WlOcXVx8e67972JPdRd9pp7eXfdD4FBcQ1PiVwfenWs0d162dbGkGW16RscbX9Pbv
6itwqr7QhslqaAy9VCPly1hs4kJkyIgu0wT4ukd7xNbII+L6JXxD95sCFFlVF3csJOmhO9lo1lI9
8G9Xd9jZIFbz075DgBHkX6Jn2Xhm76rwLkDvsDbedt+720FwDIodfdk4FtW9/y6+tHt4oaH1Zkdr
rYd3xRQ6beXXSdaDUatcMNMX2P6yktIffo1rywLzNkbI575BT09yuA6PbHoMKZGqgT1v+3nBw/2W
o0gj7uBI9xWX+xo6fxDTBxtQ1o4BdMGA+VnuUr8EacbcTojV4k0mk7fi1oaU+EauFg1NwqRCpp4h
toyjNsHsYHwBt4iuWsiT89YDYVlaNjeAP5LvmYTfeRX3fIe2PpdUrHUFlwy3/kP3S361TYkVfERn
prymYu1/xoLowsPYu4qTYYG9lchcM+3gr7Z2693rwtrBZg0n+C5lRyOVw+O+HfKjMpMyEg+m2ISy
y1qG4IvhUiYRI97iFP0qEgg+jVuZuCxK17XM1Ye4WojKwWmgO6udzBzbghi9mFcUa5JGTy9QTvYi
DOp7lftTy8p7aILlHdqTsZxFQCb/ZOyJDghmuDT6i9lEJiwtMeg2kMN8xyglTvNexzW6kwRl1l7F
2wJGon8SVd8nKAlg2cFlf6NuFxbtFRWOoLmLTxZRj99uBl+BkV08WC+qnzv5YHWu4ol1JsJkYRna
B9ftKUnB+HsTxGPNUtANUdxoKTfSMacwmzvONwW7C3+0AcTf83mB5ivUMxxc5PGMgXqC4RJ4+jjc
S6FSPindmhpINlRInyDbX6lZcOtMet/g50xMh02sRriSMl2PsjdiKDAtrhXe8ngoM/SJWe1dDlkt
b6DjdQHWqnNEr/f1I2dPQfAR9IAAxlY35NRPlx+gYJY08ZqS4nW4l++UNHVerzXVgStmzOlsAiKG
iqFkUrJcZDLaDHAbqDzAwxMLxh+rHeFA7E6b03+5lGkpSOvbM0BokMRh6KtkYaHy5aanCiqQUdrd
ipEZdvA+vgZKpPAt+lCKhciMqStQnNb75Yclj0ewNuvgbmsmMUSFlTdgukaD2FoPuAQ/yNjJvlgv
8keg3N4mFpQcpG7Dgxfz0UzvnJMzrC75VIbAYH5CUrtHdVl5aKQgT5mwemVkHEhEySOm7S/+Lgd0
LVxUztg3tNqCqSNIq6aZusiQJ48isKCxzslgae4RrZeFvfJP/5FPE4vcC2Bf6GIcV8M+bD/9BL+p
EPN0oGyuwnwFbqN4M6ZKBDt5xx8O1e1VyztauHwnCDxUQDdr4Bz8Gqu5yjZAE3AO8fM9XHtg4saW
6MhbN7AquacdqSdt2AR1RiQiDxnpETIlFG4zAXhfz6Yv+l9vGNX6e/GarvsHHn4cfYOiz3XDsZQk
lUmL/3or4/nvSQtYj3ZUn0roLKDl2EifgY4DxmMoATMTL9FRTJHQvINb2ZJB9eKjvQIw4HVa5Ok1
dxbQ3o8Jr4NnorN6iT57pFsaUKN91wp31Y3Xg5ZfVEeoUxiF3hWslDJc558B+7E8bgGd3zubNhwd
TI1LWTPcSTbgKwAJScV2jAkiPfzDrL5DncHdndEu316mtx/BvfEPDgBcJPWO+1iG+eKuWUmxbwOc
7fL0X8hoFO45wJPl1FvL3DGazMsI67rTXAIcgqQuTWaX5CFpu56Zp8QPZpxuEUmOhicNICVc2bpo
V/K+uvCaLa8/hzConplXGQfhyLoUGgq+koBXgfnkONduUon7Ra504WrPsSaTu/U4ZgH+j+VN4Bf/
VmAYO4WhVpajflbnGITaYQdU+N9GLL+2EP3yCy1Roqv9Kiczn9tFWe4g+5EU8UMzQHUvyUXfFdOv
A3I4RKB/B54KSqmZlEJAbUyW1ECS5E3IzVzK70ofR/QAC3QOPTljWdNhwhZawNl4LOgYikqHL171
Ypa5NjskaZjlYJZwesZY7DFiuvqUYrLrbY3AQWjZu89m5aMEdjIpNoAXgYDG7CoozxCOgpHOtgt5
dD2DZPVDQnMmuhpxCyvlBUBBjWkrDQIHa4/O+MI6KmR0Pe1Cuzg3iWWuLfDLIzjpJj8hMyfKGUH+
HYkF3cFIRG3kbAzek0ubsJLl6tqlnqsLuzdyIK4K86MHDf7YFKGUwbod5/7ClXqB0n9B9lfDWWvi
7pmVH6o89QkrTPq7b6tXs/JnMHIZIMbZzPu9C6sxqiS37+nRJ38yQ/HxlFFpnDAGI6dKrOve0qnu
SKGTR8+PTy1ytH5gtRB1kd72LVkE5HMd/+r/OW4RkF6P0hBFbpj/4U4KCAUe0m0LAKuADUUkFRq6
GmsQoqZ2yr0g9E0xNXZsTTOcnFuIqKUjn22wI3+Mj/9ecjbwFLHobs2yZgFvP/dKKKj9N2dB6Gqr
B0TEk80d1GkJbdcaiFB6VBcV7hWdvZ+FsNJY+YRO06BWolEC6EaiL8zXirWzWmsX6eDPFVhUkaR0
nK0ResY3htwJ/yF2DTesIufXU7gbB+6c8LEcSAaXm6cHuN2AcIkpni0WuBMGG0Fc39bEqs0j/Z1v
dK3aS6GWHzjlC7whyXmaNwmSvcuOd+NIx5daXK18LFbHQmo0NwFFKzFHo8qyqTiaPq1ApxM9HeN2
TxCR6zSPMLLJM0nLtLzHJqAaqkYE3wFV6bXQCGzj7nd0qrDUFh5MgOPVMA7PFvEwlDz5bd2TNqaq
EM2rJwAAcN5QTjkQEM6h4kt/3TpsefDCsZGSXzsSNcBQryMCvLKTMqZLhEaB+gBRICpSU8cM9Tqv
kMWw7r0xNyL+Lmb2Al5ZVjrUtA3UCuU34yyBJqIC3r0ZUGGVPJ28fFudwBWpMDwR6ObvPjVbFzuR
hKjuvy7zVe15B1Ir0mahqmqyljG+93RccUCuWKU3voBngJHsqElXjiE4l1bvpqrMNSpAOpb5UG85
SZRQgMVR9V4Eduo8/dvHd8Oy8Vyk5AX4hdQijTruJ7PToWiiRsFan6/v4rwpG7MtnA7baTFFZB4V
ZaTdNudyiFP3t+c9csieRBtv19h7cSkmd7yjp6RSCowfa/gYiJ/iiow+BLyYgQcDgOHc/hOyDB+0
xQiO1VmwRt82npm+7Ay5v3KUaUpUVjkjivEWyPcjw6B+N3Os8DnkoAzaHrrLvXoladAwKeB6wHj2
2DWYu0LOricIgnG17uY6Zq7b+N7vreJsH9F4WlZxnojhCMuz3g6haakbOnUB1Li2BKvIcM229uNx
UXURQTW7BMUYRmckOH5pKWUhQJXzS9G+pjYLDRyX1XjhTuikA36mKQ+tAc3qN+NhkJieHOyZu5EX
NSO7dMvoGJ4akzEE72tdGkpSW6rUo5Kcuu3IT5mnvTskmEHKklUE/Q7krO1mnxlGzEazw8ElEk4W
7P27293SuUQsmmhfFBUn+Z7eQ6VOHD+lzkB77EazbmC2cbizuc0TW0m5qyeitWyEBN2RTB1BeNW6
mKtCH08mhIYDCoVkwlzs35nP8P3SR4xG4Y5bftLyoxSn3jBcXefbtySKDuqzk2XJtsfYqqN6bX93
DW3pM9e4p7/7tP9bpSdubsvcgIkjiLg3b6iDxvG3BhLUH3FRpVN3pXvCsypFujNpEHUVZ/ic5R7x
qwK2hhHq6D6QhySJxQtF6oc19smoPAr5y0RAyyjXqYtts7cB6N7lmuK1k9FN5egWDxayKwaKP3I0
dZZer+bnKFQsFVS+qZlc+trqt/F1ODzP5LH+39FZLB9FfzPjZ+AWZg9aGlH0d2WngmrM56s6VZDV
qqahdFFuVDtJVsj0vv7yvCDsxBdorB25cuX6c7iJ8zXq0k6Xt9OZ7guliY0hS8GCXAeEn6PzVmUY
jzWjcIpgN7d4PvgTKsB4BD+bGBX/esKCY9AabR+YnsyQF9E5usxvzGQ9tgNfJ5HXY1o7sNJ2xVfi
HsMZXeV7QG6mkGWGjhbwFaHsz4sl+1A2CBu7i8nL216qAul7eHhigzmody4KkUXENQk6ILexZ9gY
IxV+tGmZQtvjr0SezchhKAmt40f1E1oXhtgMXI0LnFPToHEbK6Wvez4qQzjzEaOt/bft0wJ2ih+N
DV7MV0NUXleRqLCbgcXdtgp7IOcl+g+VqVN+Qi4C+zLHn1kVHUUWWXjA6AQlJxHHn0LgpfWtjRts
oOz6kyPkgvuVSY7sfvB956BSbtISSQwl8jhDLNUK/fs/rXn3K89tyW8rQ6OXjGkOujGqZyWwrMgp
c9kh/GTCxhb+wPHH7CEiQfutwGknkwD5Euj7JBhxg1jq5bzcgV+ERj3vzlOadMgY1XiIKWbg1Dvo
n5jHndRJipwk75ma6T4DMf3sxKZer7QF7JpRnsfmPqGuSVYr/IcI3PFXSyObggU3zYCkkjY30k99
PFXlX7MPMBYqqO5qeHqYW2inoXZbGKLcnSIRFtoKA93P/xsNDdrLYQXBEuGP37scDve7TD/VgDsc
I03pGQVww45BF8N8tkck01igUFisszgcerCjcJJax6xn2N+halo0mSuMT+VeGfaQbus67rQqwbEX
i8WMEMNNb48BbDAxLbw0lix3Zf5ZFOnoND/7QIUX2Fo5qm534cmWlRF4l6319f9xgDee2QCdl53O
b+WlSl9c2BHu/pxd9QK4f7/GL54sv291Zi8k9Pl2vcpd3prZ27UbsBA4dCMlw3JGrdLD0w6/Jdxf
xE1sAb4+eGsTyHK+San84ZBV0/fFy8/5xR0qW3PhCa7EQ72hWyAITzBroXnUpJAtNAf+5pSIGjiW
4HUr6mrwyRo6S2CYHJnaKx1EPSQWLWeH7xoxnGew0herl+3blFSsXAS+tZqvyHP0t2JDTzjUQdA8
FKZeMNpkG7SLL5iD1Y/QcssbtrE4/7VKtyfmJywRCwp8u57yQ5Z2uTPqigQvO2DhiQ9C0pb20OaW
cN3s+laYopVmyelFLMA8Gzc61o2KrvdXfpaRYcle8E1N+SsGyFkLzSBy7nkdJv0RuivFUIpiKioh
VEvQAnqXG7h9RFJcbLN7rEAZwpDM2rYgvVWCajUe0fM8LU0DeN5a3kDYWX0hW7VerchiQh0X42de
TxZ0DA7Qe4K8D2JvJYdJEVPhr9fl0JE4ND6Ex/WI6hvQvL9A0DpKvgkmZikTaXF0MBR8xbCU2mkN
bcXQvgC97G68HJJsDZkWhE4j31Z756xrnhqHbxt91w4PsDvMU/QP0IspXNjeg1s9Qe9nZYpMHwfv
vVSexvfFL4IhnaIha9qLUuPP5Pdtcme20W+Fe1p2SyAJCxXYOyZExJZGXvfh7E8e/eYqqR+fKmbY
Xbi052l72Z5cp4apO63zu6CdRzihVLZ00C1bqlphqDFmwKtitGBpTx/BGz3ZFWas0cXWtQftVQgR
HmJxuBHj4HvDAAkGYjthUzifJEKY2fM2azpQlJbACWf+jtT1R4PzbQ+qgnXtfDKKDC0TiR25dC0+
HcJt6nkV59NMeMkEpW/PxSS6i7T/Vq3l/cHs0CmDwsVjbv/1dTib2if7c+tSApsppeU2GBGtlN8r
/RCyK3Xtp+EnmXVcGHt3HjwawUg5E0FLA+JZoRlt1x+uxlYgtf9JXT/y0DgOJmvsvWsDUsODcwpd
jpxwNWvoiU84nhjlXQTJOmwEQ7I7QbfgG3qkNs1CrjaU4lk4fzfjV28yLsd9xgQr4vsAhzv3QjWk
kfm9U/B2wovHDloj9TBwRpiTz7yXFgdRBy1QP/hqEkVXXl4DJ0lsRWchOiFf07XU3RjM0Oh3oDei
O+PP5iu+RGuwu9zXdFv28i+gw0RHHtH3h8K6CwTVyGGnvWeRjjv82WOX+qwnkkDZaLW7LMzdV76g
31szpObtGZOzaiVW5IUV5ztjuLcvbk+Hq/ze4v3hKdIQt7U0WtyGBpP7fAtGq4DeUmB9BrHpMrUL
rFGgSGLQLZJYF7/eZB9b0FozOtHOnOrDaT1Ry+BnbelR7kE71Elg3jJ69Es5A9j+QWo2V/GDxqQs
hXczl9TbqbxZ1dVIPx4Se5PqbrYrDhiI2y7yymebuqrrWK782oQAPlORnHhNda0FzHhVNTzfGkCB
fYElX0Fa2HKerYceP6V7UkbnoSkgtJfFy8UYMwWyWq/BMrpmDDyUmefrmNPsAPH0t4XZEYflKFSk
BYLcNsfET8gJhsmtkS9aQs0w9dA1ndjZBbNjyQKXfrCG1sX+Aft9Ys3KMY5kuWh4WxEmZmp2DxSy
ovLQPSZtgsXTwCjUIwgetBwlkNCnMdvOoGC6oP2VZyzIgMqO9CSG8TS84j2tYo351ukG84vWur6P
q8H/4tCLur7tmnsZGl6CDh1gLba6tr1vH71+IE4ubbpsQWb3KT5SQBKmY8KKnyLhirEz3DsDYMTg
lAuN5UhPZBarWpF31XfTpSV9GId/UJbQSZVHt23fD+iQHBa6fSBVeXPCOFqXgrvc5hObbZuCXLlk
Iet2M9wRHbf8zvgraLS8mgY1bElvP9jMf1Q+768xUyA7pI9iOv9CwRg8Zar8tsSEVNLki63Cn4IS
EAtFBrSpNP29pAl3eHxfH9mLKr/3Eg4rER99Jm0lTvId5m06/xYESkVHloHHnIY67ypgnyQ2i6+b
+Xl8Hfsl8IKDcaB04Il+c8X06bu2ggrVTQU6z6FCjmZef+pP17qgbqa3DX0tPDcujJDGLRsASj6K
Ew0XZHjJhMWQO4NlK43zJS7Nzm+9sw8j2fmtD3JzuXnMBVDhyAzdeq2rQv1K4XOlv2eovr/NRoBX
Ljhwv1GlFlIkDNKFACoae4Bab9jAev8vnnRqoKecRWc87KF63Wk+RFfBY5V/fbd47aecVEP6lqz6
R/CINrzANv/uRD1+ajZ/b55OUBf+MbopHb+4ZlKI8qsSVms7tc8L2Gzyt3JvJ89FJfYUAY1ix9hM
l0NK413E8DTgnx59VYFCsOGt6RNbgUfR1FAq2FSRNoRqGOsy0U7xVcYwAXKRdfCjHiGatgdylemS
k1y9rfClgH/k2LBTVmI0+ICMj86wrdRJv4M3m+BuTzbUK0bRUNe9ROie0o/8EvnjnQNp5+iAnf2s
yLtUcIPqwdJ7I7j3CNjWEgusGmlPEQy9jpXdaOajbt3HP19YZgwCBCqQRIVL9AyEyqThMPDSVxOq
dr7dXeWQ2xHdiFe+vcoPldD/qzBfnV/U8O2nZ7fhIPlpd0UkJRhueU8vazEX1llTchfJ/jYeSY/A
QCnVU+JpcnNbJa6SJvvhPNVvMBDFKDdrEB4aypwOi0z6nm/beQUqORBO0MnCyp0oJM6lerypdiCY
D5vkQZZRrgHYSRQMWrPYEBoF5NVBh5eliOz7eoZLDooRYisnplPNnFzQwTFTZ0oBOt30zM+0SQLQ
5cRZ0btYC1+H46lo9NN5fk0lgN29092j1hD053Z6qm7Idsv2kJfHkaHHnFSW1bwNSQk6CF6LOs6w
9nwbkbah3++fUOkoDAw9bHy56kweS1bIlWG4dIBypSJ2Ek6mYCcQZdFQRgLNIimLUsFsV7ePWhAG
dxjaJiiPkfy5oylzAwoARaK86QI2u/S3KiDjZ4YYffMFms0u/G9lb3n4KO1M/PXaJHzlUoYpHzWu
ony+q9ICTKKmDLjbrop9+9NExJjo51mNQBuOUeTAnlaqp4jL1FgbZreaB2zy9nnsTjUlAVcdQpiN
TSrPqRGx+hkkpZk9f7o5G9RxfUSbIFL/FvPMElWOXxpELcutZxoheYlLk07btjMjRZlRl3NfLnFQ
NHFVu9M1vYUkAJyTARsOLxpEKqlUlNgFEUY+PTbZyz1IJBTGDfK636v+DkyKdwkyKhDwjvdTh7KA
GdLXh0Lgc1d/H9aMxtw3Kt38iBxyK9sJeQvf4IiC36UWLqiubzIaGwrrYtmcqmoE46APi9VZ063/
KegIrzmbRucxcDdr7cbYU7IdvTh6a3TeOu8vhHlo7oTwhNWcKNlweDPy++ikmkUupMJb1lx0jXgG
IVwTYzDuIWe0BTuz9G9qQjyDSSW0kUFbklD1nOFeXMCG+yEUx+oOliczOZo7XCFvk/KbNFlhNKMr
Uea5iHiutTtH7NzUW5presG/cO6BsOLPBSWFd8yaPt6d4UWLjTtMc7CycfHrAU/s0VLdo4AWG4sE
lggfrQrsinnOizcQJQeYuvzhCupxxP030OGVN2nkCeXOSE3y6T1HShY2UCD/wgSgcT2MRsD3xOzS
1snoEWWK4XWR2Dmpszfspjo1xoELhtOv5x0PlyrooJIACWdudufc68eH2HXcL/A74R7v3a5ecs+2
4KuV/Ho8kh0v57uVYCBINwTQp7/z2rhxsozQXDvgHkAdl4Wmk41otz/HklVHEuMBPuvQWMuCuzLt
a5IOCe5v0vD3VOU/vfzvgkPqllMZt68bFd7AJSoxsehN1XbJMhcADUFDceCDBjzTLoWtqCwyKhGv
RqqPX1VdOV4fxJtb8nPXMly6PTxNd+stdxi/Uc54/VvfpwscRdZxZQTyew2YXvj90CUEV0oc59CJ
KwVEUC+VPiP+HhbsaD0lj3Suuwb2WTOpZTHLUDfUd36bVa1Yy53hwrWS7JShDecFMBRpIZrY3g1r
cEX+ZpXGBDuF1zqdQ/AM6WKW6lgdKFzCwjWIe553GlRSeEx7S7/eynWCG0i929u+gZA4Kiotun/L
DbZdgKGqCwty8s3mZeUQkYkhYWa4uyzVjK/ZTgiVPi6IH+O2DD/LjhPcgmUHROnNt2Di/dul7qIi
4CZtaMosKXzg4+76qZzFLgMk7owDptmaN7bV4d0UFDjlOvoSJQ53ycUWMWNjZEhz0bAdNQ3+zDAQ
Br9a/oOnKE4PGhlBOnnytMCYViG0sCTItmxdnF+X79BocFdg9t1QUz0SeWg1eT1zj+5D0sF6n+LU
RWovnvvMqmA/ed1iFnxeJub33QTgCE9CXnuV4KM3JTS4j4b51eMRR+Pf2DAUXVdk6EShEqyhI07N
MJ3SGpDPkYBzbmESY53PP4/G2jq9GlPvflBexWOuiEmx2wYQwEbZ1ujhQ3PjuAWFg/Wa5ZN2v7x7
gaDG88Yww6iZElymc6t1o+JyMFBKZZXMlEXrrf6qgEhmK4yS5S42EfwP3SEXdFZ857LNF9fWa4tD
cfl0waNcddOHCq+fB9vIRPVu8iFQWnGwMVCYSIdMmXQWFBx9k5FvVcfaFm3G+viVyMz7hryqVgzG
V6CGkxw9pM4DYStIkr9oPrO9mnjSEHzcioQ3R9XsyzGrenBzq8m49fLvSUv79HARLT0rZeGRk6Ka
a8ZVpXkQRcTY4w8RIx/DDV2gGUWsQJzB6ncKtHXJ/G2PO4G2059H+AjVr75mZDIe3afShELCZOV7
qIZib6mHLV2pxEoTH5dE0Z1f1YvSPNE65Lz/QuQxVpJoRYU4EMFJTlBA7dO1yLL9FnBX5gHJNEt2
rgb2fPRwpIxORWNvlvTjdwQZdHVX8pUweMX6RjC1GhHHQZzJFZDArulp156/mamQDLrpOGZvP+dA
rkoo+h8zDHV5V3TUlVQQVYsomCpbM03R/9pftVpR+0G6MyTSfWv8vBfcXSjt/439BXHk7Me/Z0ew
KwZ3RM12wEv8D8svfm/P0Sv6fU5A/XfMSDqIZl4WoVxAWj+6kR5UuYsK7Lh/9GUhp95sZRQnHdzA
dGmzmLm9BECGhwzUB9QPqgIz8zZNOCPrG+fjtq0Bm7nyd1CLZg3c/3ixplZu9TjbCK7lT2pTu0EQ
PqZCPyK75L/TUL2AWSYzXAwtOu6IoJV//zUEpGZmEbRSp4ui2M7BBoVPB6jh5Xz2GMbnZ9iCRrnx
lOT4tIFAauNeZRMjnsAF5QpK1ATrYi3iPdSUcMPYeWNa333k3eTOadn8288WEw2vYwI+OoksONJK
CYf8rqv3PG0WQxXM14/oZ8BkL7jH+pCKGuJlXeFjFsOSfiK4mIZCN7Bwc9qKYvPlzcPfahmVt8sT
7CKPmbFbtxAznM3q5KJaERqabMd+cvbWKSIKKOkgFNzt5KejYJAl+Nf2d+7FlOAwgLEfwHstMGI5
qmOaTZmcMv/4gmZdxFxUPygmc9DADqNzaSXvdnaWKW1Dl/QCG4483P7+UoXKRL7zRc6W/A7u7+b5
wm0lr3MQFHFYJBgOnk1SbEwziMhOEprPXUsOFGYpPRzHi7vP8gnOCeMLAI6YheKT6uqcJr59kkO8
QcLVFR09EYPNCRvHuPSbqvQT2XYZL3nshNO8OQCMnRQ35wxh4eC80i+8w5pemeWLPgOxEGl1GHrJ
lq4JgR6NIBDmY1MJPDNlsja38Y3jB5V4Jp+Z51eqbMH+oRZSqmCDvwt7qR29SRiLyCDBCwWkUNPi
4XxdAPDm+jm3S4pTOBd2KuFoYtzi7jotzatyaanUFGKFjdnBdOnH6RoBV5Ymd8QiY3gz9EhC3qx8
ly5V0g2OENMNrIBI/IR5qFnpiEUd1yLPhWxqJwFxbQTqzwUJZKi+d9dg1WZIFM4MVFfHfpNy8h87
z+QlKdf8olu2trZ+wO3mBqYNdLbluoPok2QfyrMnS7KMUiIRgQQ/6eXKnFMBIhtXMnCRnnKXlOb5
6wEZlWaXcXyqfxF0hnD0wNTdXgfJg5WxD8h8yEkWA6ldW3jtHSgEJZ1tCK1fNnzCxndeYuw6QYMG
EoW+X8D27v1e320PDB0hAXaYhGIgCTlD3ESKZMB4z9VP6VTfTd610OCoLNsJ0cTi61h7t2yUobD9
ueDIKjRxg0wCKirtiTIW0wc/mGaQdd3RKXWMggwOaM1wN9+5FPb2jFpvhDfwYZQHlLhkczJK+j3F
+W66TgjKarJaTPLNYe13EPzZ2UL3rQwMKbsSgBkxBLrYLbJePlRokowNBd+ZP1lfvecyHBM328di
lrZgGuNxw3HP7/oZ61py6tTYbCnXkhXgbAiina5DzaHcE0N4sE4Nj+RdEJ/i+iGsC/h9pibAJHRL
IdHIm7wOkp0RKBeTti7Ytl0ajODZ2/OmEarBdOEVA1CgPOVO4slb6GrmOQIVHrLthrGIoWqWoNCw
9/xIaM4eQ6at+MYL3NJyjyIsmZ7o+LDxQNOfMXXnFSLhb62/0JPcE+o/bk0jwUxAxews5V8ynnj0
TE8TG5jHDGGb8zjJHFa7sez0vn+KY1uPMJWJc2Mi+WPyTX8ne+YT/Fp9m/oaWwCMtfb7rqauQe1b
QpcyIR0DsOKHFDGHuKdsVYYwkEa+WMbFygron+UxmD+ktKEdxkDHIrfsRljpldOrW5GFqgiKj2s0
xDEkaQIg7SUQIEYsFnCmOHWU4Zj18mPQ3PJzG+HCey3ksS/o3ZONlvHIY3IYSsW6WFFR4Lzctl4s
q9CnQlkYal7/4h1Sf7tge8USoD3Mpv5W7fHeWJmzEOMeF42DrGBOCf/NVmKZ0VfXEI/exhRrDwDn
IYyGdesIEgN4Tr2B7vBkEGC+CBE8FVX2e3gH91k2D9r9YeoOcLtagfnJ34qYjtAHEPxwSx+UnGn3
ZMu2hM7tdu82H6N+LvcPxEkAS+DQTuOgRlLRciybaLYpjDM8ISZkmQ7H13cqsukgvf6VFxmEagXt
L7hRDKBLTGrtpVRPERGu74tTl+kGJXiPDRNetGXXhI9OgxERyVFtydTPUJ2WmgNHI4ZIZw018bv4
qiME7Psu/EfcUVpvEeYQOdHQbvzc8zbCSWGgi5AV1z3iZZ3+lxNKl/nsqx/iuSBk39kxztQd9Dg0
roGGApKo+qAXbqRZvqGEW8BeV9l0mnUU66oayRqaJP+KaitaF7Bt22BenXyACNNgT8A3FDRrzt9Y
3C0Sh7xof4DlUhZZp6VjtWtBbmqjVHwzOjTJxUvsCjxn33VuSplGsMsD0JPFPNOiM80eIePYUBhf
J8PE1QCCLeDMCqgebBl3KsvoReJdWV4EqpHNM3chO2z/0N1pBGoRL6DqXCHmHVhahYdNoOW8gT6v
Xu3M9CF/wSaw4EycgC1MkcZs/0RjHsO9gR8jHjcz9XF3vdx6U6V8gPTLikgaGd70XeoOul3qn3AL
ojRcnbXUruxI/dxiXHSG0vqCv8ZXrWQVNRbC2riaFi1ruhO06qvAPAe5Zp9WkKSuqB5oFRR8f6LF
SbXRRUok2vVT5Yxrc3rzg4P2DlxH3qLghe6L91xHROAPwGgywwyYBM4ph9mXXuH5qy9IEZjUIBC1
siA+1udY7n+aZrKw4gqpqVQl28wYKL78m+bGlPxIUlSjBcFYgnHOYRT9pTjtoG4Rtj+GNcgUSMW2
ssjXQ+6fZDevo1nqzPrVeGxBnZ51Ozxy3RfoFGrP6tMQPq1pOmHPHQLkIFoSbIo1PxE0AAEnEFs7
S+9iYpN69JOk/cV/6yF8KE4DWt95ZcuTL6bqjlvD9nxRKB7rhJ12E71oWwqz4VLo1H3XevB7YN6n
9rVXxzba6ok85wUBrJtxDY2A7Pn7Fg07R1fbYKkoYnQzK1LxAg8XWQCNhgg19hzV2Dle84szfhpv
YkipmJwbH9igOHzdDITBtzAzQDegOYIyceyI61StQCxkIlBgql8Wa1/YxKiwTVu72T1mnKTSChrw
WYMXy4mBapYYHyyhPrqQOhgQST0cI0qUV+9vmd5sVI3V4bskVuTsMf3vQd2FdA9FdTkC2Y4QHX9V
JJpWAtldWbTcubgerHyFtWddcneTW2u3Tq5OOK7P4AsJjDQJKeSyRc7nyX6ip9ctSi59JSMhYXsA
3NHVZ4ESOduRMhoXJNHCplymmxe2WA2gwSzMdmJ7PX9k9k1NtOECoRUq1BtcmpCbL64DZX+gG9tw
LOYCYFaBbTDtD6AZrFHESnRPfXm57Pi/NzwZ6cX9+Fq/yKnuEOTOMDy9fDfxA3Oo1ppWgiN2c36P
mUKsS0W6vNnBjkrgpdSj13MaM3ZiwBnpsAb+hAQk0ZKy4dCOJCm4FZ0M10mZ9QvzRjeaiDSn9KbR
OHmItDbz22xM2heUNySh8/Ld4fYBsYViLGnEie5AkeDLk+HNF6e11Z/dDwMz4kMJlRNSNl1xn/sE
Mc18ea3fSu6UBasDB3TqTsjQbSAxnSxFULFcQfLf9dZZfW/Pni4DDdiv7DEFPyXfbCT8iLhVB1Wb
iowK9EGZIn5BtQiiW/MdEqGJZEfcjS0jGH/yDn5IKFf8bVA8sen2ATk7IfhhPHIQTtc+Erf24uq6
lBP7FMLF2DYekAF4UiFG/mGnONcnABZaG9GFXy++5osW7YFXPJU9QnwV/lEKhWgF4dsLYfPKNhWq
LiwQABTJDGFK0a1ZifdN+yxE1d3c+bFmmvtYQ4vZ9KFihzC8L6JBKIzmd2KhAESVemdwDQ/d+Zxf
8fSgObvIRYg5flo3rg2C8wVDC2v7Sa5Pcl197M891la6BQ8l79IudvWP/zoLfWl7U5VLQmlL6Yk/
4ICKRc1kZWvBEOdCWT5Y66+RacULD+g1AVMLzQ5qrKxy3FtWrckm5j+liGJrsva4cXtg7vHo8Wlu
3T2bUCE9becI9FWzCh/thgEmXEDrnwydi+Es+aIR+/oN/I/NQCJ+hz5wlnl21MnnJTEXRcQLuO0x
S8DvUsn7s8SA0NDpFnilibY0xMErtCWHX22r/4cjIeQMdjTVysSdWhtuoGG2VIgy59RYMGtCmC9e
4pnDNZf8cnKS9bP0pwdkaEuu4eJTqcovWf/StqkggHd1lteW3L3jnNThRwPkFVurbf0qyvYSpPbK
AbaMACmHFVRu6lxJYXsVQUUys4IDwcraqGj9J01a+LkZey6Nn2MERO7oqlyvN2h1IRq+qyRKjC7b
NxoizxEqmuXLT5wylAbccAA9bHZvbQ5rLKd5JdllHghII+6H13iWU1z7V5moPdLZybCyxhrDzlTu
gwAaWc1RQ+urEQOIRU+htQQO7Oiv9m9Y4322UP2ItC6oSQeodsyjId4iU0tzXNThvQz4awJ2+Zpf
mbT0vGShURq4DV+vVs7VgitAeBSM0tpSxYRjXIbexpA+k1xleavtRaTQDbeo0x5lQIQ9u7uU1YXP
q83J0UGFSjML38/h7N99ROK3qBaRbCNMubjmlcvTCsn00O/x4LkcO1hUD4P6tHsPvPiZSdMp6tlS
tsD40sj+zR4QWIMuHzusykkWZbuYWX3JtEABgeUQZJLdNFrW3YI/1hIG4o9aBuSccXNFD8FZofDW
g5kim5aCsHmKxTCuGzGn/gGKwlpf/6Efdkv3CIl4HwSJbeHLEOKYKIBE6WJX0+UFzHtjt5qUdZLD
69TQHwf1+5A/uhAXj8bMb00ZR4lxilfZxmohDkRRqp25S3f1iNQDA4/q/NIAVRJgJdM1XNn/rMcK
pxFdMQD6wHeN8hYefkTw7jASCEvvzIwSlHh5uw7Ie8hiieADaj4gWqmZ3B4JcyGqxVUSgdUxZ4pj
Cl/T5pFoFZ9fZOKjoSNxt45kQQvEMYxu8mQf9OIM2z/0nG4W+n0AzJ3qwjRxxN7MtYNQzlEAhVEE
CNzW4tadOPXFsVbGItWCP1CYuwSVXkUtgL5+EIemLooRphgfG+PUbHGFZEdDbueJ5u8y1l421RZG
7uqjna5WbWztb/IKWlF8VectUczEThmrCyiY5nfRgYFcvRBcUaxAr3P7UuFPYuYc68mB1g3EX77j
2I2EBVYv2wVzdvKjRmv8IhVEPz8ONRijKzWLrz++aIfVdvtWVXiqo8tXDNJUMtZPIrTK1yE1QPW3
gr3EDm6bR1/tpDTA+m0iTEdqdtB4xjy5937SGk9QAc5AV1BESIId8OV3smzNB/Lf5OFhPHVzmT8/
0uwNCtigTUEre1V4lFMdsLTiM67+sNMGa0yvF5TBRnIV9rj9Go2lSHiv+BJegG6kb+srY06eJ+nj
bS3f4Us97DM5ADINqQ5Pho5mr6lUvjTQNT5W+RZHg9C6iImeonwxHuyV9IYKXqgz1YESZPlTAaSn
EHSF/YzQLx/xNKIEy6KGkir4Dpoq/VlEOJJpe7UOXNZ5SYI369GfrB/ZQnpvhqufJAFyoI37npGP
wTpiif51ABGOz9r+njaNivw32wUne/x0bferVQ6+sXymbz+MOTewwfLSPKJfslyWm/k1iQZbc8sT
Ud0HBe3xMMfTQE5oVNgXgzyb2S5bzUK9uIufCup/8voND57NOz3+YeCkM8bCQvQdDggvcIHGdGPL
DR6my8bfkPyunDyyaFWWVk/l68H6ZP7iqhy803vFk1ugS3We5+aUJhLbt6Y9HSoHjpde6uwdP6dM
J4+rwyy8uI9WwjugXd/RBLkVR7870O6B/nZ4REzrKcTbSyNeISHcnZuURi5rvZwiOLLpGtwz8nIM
Yg1ZigE2JsVckI/1mpsquLG6stnUf9AH8oYAAkmXiMz1YZjIaNCd5+UqrbDzalZ+VbD4ryKumpU6
Vi3gChO+H5TzIQgFVykfr4Ohv5cD6EF3MSeMJKyJZvsZe46GfTr+taH6WT0CrSHtwb0o/fTcXPyn
8NqU2bh7CuRLBpJBxxc+R76WFYwTkFEZXbFVjBLQkmVcF9UcUxRekF0YOMHh+WagfDIuZ3gT+orP
hpXPtGhkes3vCR8z9YQpafziFOo+SIBQzNuMyaIFi7JvClihugmIR0cLfgLznYXpicIuvfAyhJQO
BeW79HGyf/sydWWvYgBbsIWwuvJGJBifGJXRrXATbQ97TVDixkDUh2EihCDV8voa4u+i7IjwcCiU
seCD5UXysDCO+iLhhYngMdOtG8W7OsUrtCdwmHNv7eDOW45Zr84BCtcunrUmO6QrI9ZV81+9KYIZ
W1V68td4AxdvK3C+EqQN1duI7cyXgovoNWrpbdhk1irC0pm82HuxFZ0d2wnY4p+G1ELxbQwx9JY6
0iAjME74gAUv6nbXP5A09XfHyBXKoBK/zob1N2QqTtw1ABgJIY0MM2I8MmmChzwNBYjv8BPHv0y9
EqhsvDgTAHg0Lfu7AG5fRLv8rF4NxwQ+t8i01MkZAisRssZl1ep+y9cKvvatxkqoS+bPf7EAqfmR
P+DMTOV8jI/9yP/5/VUl5AB0c65r7klR8y5z96iHHS60xNZvh2v5QAUlxKioqKBJ1each+QLKauX
WV4pMJj9CfQesvwSbxtQaMozu9WPzQt051dECIAtcX2/MHnYYhwjrXuEJnij/c+WuTDCRBueOM9p
5oY3JkqEsxIKr7pQ8E6sDgevhqXy08/K9oaVedLMnaWmh0LFDB77RCJjP1fo2cI2JfpYcYxIyeht
CkU1PMGSGK2wUuPesVbZUpN+bl0jAxVaPPpq7CYIgqoMIyedGdSrwNFJIzDlDeBjQcwNf+8n35QY
FAwsn9UcECbGHxElMxfgRMOyJ8q3iOyIqin8aLUPOChqv6UkrVl26J1FsxYctyrkqvQ1Kgeo5coT
C4M6zHTKoZo2l85ar6dq9gIfkS+JFloANCQzLqBJuM1FVSK1ebmwCQQ9hDPsKEsZx7f6eysatjYH
NaDtkSZYBf56avQOx+laoK60/BkN0eT+W2+d8a7QTOsenE2XC5ZrDSs46Ixno3Ppyf1mvD7g+gJU
FbyJ+6FQMC+2sjKghpIXZPKrrEmLyzO3Eo/9bPWEdzM+fZSgU0hQgGtwG2jsq1+udceNbnao/nWA
6NjinTrNe6m7WYXlDoLuWND6oUAlvymSs8OflCzbHnU4+l77MSq00mMkmgFzwFdleMzmPWLC+XpH
6ckTDvb20//othcMJSIqSFWH3fvLDur4siXl4CV9lJ+2IcHx+OgjBk4f3IfaHP+DlTQDDl9k+4Fx
lDIkQ4wcRiVzQPtdF1EUmAzheZr2kKBRXhRdJk6WPSEe+8RURe8Rtsqlxv6lhiDFbkS+tt+rN4Zm
R3IwHPNMVqhikx6XDqC9h/438he+KNFC9JKX/cr1BX24XR7Z/Ms02zk6WvGvv/4Lx362TzXW12YF
K+iBeD+hHGZdje4atnh6U6zRdyXxiMXnmRXkHp7Od2nXCcqy+KVun6WdfjCMDIn1Wrik1cpgLLyy
vwoCWKmbzLPs2/pW2Pb/FM376N1GzKuBQLwBynl5w/KbC5qtt+pLgFHheUpxVn9Nbex0PhZEAd7u
Ev20EOI3oSEFk2wYiBSw2cS95tMNvq/1YgGMxs8QVotHNj0a6OONv7mW1jHS/JfBgUQo7tGsvr55
Yn1zXDLTnLv2/imJVbX68yteVfLU8wJM78nXpBaam+kmLK/qozUipSiuOA7nSAqZ35UtY21LUlkj
N1M/XtF9PlT2p/Sm6wz9akhasJ4AwHH2G5aS8RQCPQgkPMaPb24S8L9BIWe4GuZrZEOANWFfF8Zw
hL1gWgehVTZDjouv7242R3WrCs//4ate7o+9lTO+KS8YrboqOt9OF/LGuKx8pfsQh3oTlHlXwAXM
cASwHIjEDjOwFYbvdjqRFebhK2mwuNoHtDwPegxDqpu4lu86LyAyp1PaR86iUL7Lyp25ssc2cAbN
/40gjfezfOiPgUDFWkcJcNGYxk5Lv96ViwTu7u4jaDBK6OW/BMiStALotI0EGjex4CBH/AUUzTr9
MSLB7hVMOjOpIsWaJZTt+XJj/pMKoqXURd0YOA078rDK++mffUmBn2BQfxQJJvmt4LC6SiHCLI13
ynJRAaBMlLDRwjU5+nZlDwM7gt5DeLb79Rl8XXlV9DIuNHXak/em8zQtwNwBNlTWx9P55FJI7SjD
rSqWop0wPq4Hjx9jpXLSqtPna/lskSVjuZEKN1IBQhKS9mHQVqpf555BQvAQfuhfDnqGOzCuxHNm
RAEtK1SngdnKxfdrtg9XYsekJOQiOHKC7r/OjQ+bifxjAM5/C6XnrwIJaNgeEodlMmUpgQ863rdB
QmhZjsW6CC3zeiS+uyE1HFyftJKIR4v+kJ7lTG1Y2N1DD1JbuxtH9PlO6O3DW38DjRuJQabR+jpD
yNmw5J7qeB+1vipWfewdBKmeDy9H1NzCOmlWz+jqu5NGNwgXuL/pH8yhibrGxLixnf5ZefFC3bAS
EHeU8vxUqY1kbOfDcKVHR5wzh2+0l5uRGdCJNLHXbA+dzdQ6XyPemW0cjIRfnUFCkNaCbcAGn1bV
h0Pz5+Lp69c3w5RiHhBYT63v2kSjPmNMF0+DN56TE0zUdJ65Ax6kLacLgpjK1FFbO5sQNSEo1ULD
RyYxEfa3WhhJnyq3kg8z4Miy4TLuST8iXiaODj17W97k7SZ7zk7vVVk1x4ogS6yw0F3vsEaZUYQB
MF6mH6ZiD8XLY/MllE9OYHvfzH4/GyIvhcYWZnCWzQUZMN6F3gBbHBBsxAGrHR663LqYnpyKhnz0
vO1HtNIBK1DGf7zHfFDC192AR2B8wRWUK6QjEVAnhzbjxu+UkAG3ncYwAILvZvOzV3GXQcF6Tnye
uwX7C0M5K0yP8zHt3XnKteU9ZESRI7Y9hsm7P3juuwwnUE3poc8i0/5smYLVf1390BBcBaX2StV6
5qxfspR6O9O26IgJIFocT/aBz6wQUiOBJIPcLRsxHe4cKRpPru/FpK649DGV60eScREI6BhsczsH
7SPhu0mfmZq8GwN1Q+1mg5u83+BmDVSK1oeWQfYilxahww9KAxaET5xt0wZaRkrIvnZ0FurI9qNe
u7DAmp66KIuzBLH8eyzOrp1lIWaeF8EVl3aHncqBj/MlBxDyFHd3Na45JkMoTdUieowu4UwLWz+q
m1F+uHkWVRnj/KdsFddjznww5Nty4zrqMF6yqqJH+V7NKJVkbeNVaOXPZmZEz4bSXcFtG0XMUjRV
ntOJ8Dx79buVAZLC+L86Dlr+rBZ70Whr2AwKVYF+pmH0ShoG8syB5IgbRfu0brqfTd9vBAcHhpDy
8AMYtF/ScSfrUV75k36USbHqGh+edloIbBEsf/KZWGMmyc77OnFm3azCkTC1mCsFN9TQqXk5MLRS
z4oRDiPPT1VCSb6BHfiWKQzEv9NIO5IKsnxCm9ik5jOobZMcOr/3b/YcomcL2VYOh/2e9QhCqS9/
mf2bsV/nPuTMBGE+lhaABBIfj5zCihY+8BJal8KmU2kvHlkaeWzWcjVst5sIpQ3nx2zd+ZPm02sw
Ouzrw215ECESLhCxfCjUuGmRCJwkR5cbUiR6VJ5z1Mmm2FWY5H7dv6VS8S6h3zd80MIYwBG69sHq
d4LbnxGl7BqPNprf8N/JecqOqsyA27dbsvpAzMyj+tEkPxyVyC580hAJH90SqsuoPgXSXf8NCuFF
uGAxtu89KEAr6CrlHCnhQDGxfP2wwxdv+rQzwsnoC+NAKlGYfLT8qcW7CcFkwCI8vSlMi4CV5Dby
78GRpSvYxfhNYsZgKwEm87nJ7Z0WC1f0houHyVayxNnabY8V3tVx25LhYdl1roD60INxPp5h8QSf
AWWlSUQHKsKztjfXjmy+xGpSgOvkiOS4cfTYR7F6dzpelyoYNbIl11G3Rgnk5kW1R5BfpRzAkzXB
cCh1ey2V3F3P/tjSezYNi4NTmnP2VKMTS9PZv4DVZslRuR3hNEcCOHBfuCGO02qonAdCJbo2xxCJ
zGTqYD2O6oFHaCOBqDguLB6psOfPKK0Rli9ZqiuvvbXjSVDhX2eEIAXX8CQPEcaTFBFgeVLIcduC
CKK6Ls4dy1seD7c79riR8Fg0TG4sHu38UTHj/Hxag70LO9VrwLdtzCzUZ81u+EYJX6AfLUeZkafs
Odv3Ba+0IfM39ZtjjYFWhQWEhBSzrbWDCaNtqJOLxEMZI5bSg97uVyna4HFxJJG1jH12KUx6DNJj
xj7mDcNnbENKES+S31K6U0gQ97iYPcGe9IuS3U647K8hF4P0lATGaVCJF5vHaxGgc4OkyJzCCn1Y
BWbzrICrB9RRIb6lxQhJavLeMQ8rQNZ+VLbxn2ReYwXV51SL3AFVr3+vMA83PaP4X/3D/8CMcIp1
x8t41+lnPzgvqoR/gXwnDK+LyZ8ehaIeJaAjULKFlxE+eK7yiEZbhuONweQhZM6Gr0zk9WbJZCmN
LWwFfs7OqBS/UAalxIJvsS5XrTh+ueLQc5G+8NUyBWAFbKvL4kUpym3/qI2rSonXK0S6wCNXo3bY
7/aSIWL0E+eRzDTS6PUFrVhpU1C5cq3YQPdSxv+mQGfu4Xc3jKNrFTDYSxwvjen94cImXCt3mUeL
pJXSiWDRUi8XqBi3eCkRZ8oq3qanbj0wB85KZMpgaGN1ijiiGtbE1PlaxH4RoYKU+09XAiEBvzo5
wrwArYEOqpgjE3o5bz799IwR1e3O/fLoMLu+pm622urpuxJnOxNTSZrthh58rfX0jd1DWq/NSmkX
pdR/A4Eo5M/ZCL6XAEtbo9Cjd7hSQtfAmViAck2Jx8sp30T+Rq/e8QTzDrxiQaZN9jqUGa2MJZ9o
OuZ0MmjAkQxQL6lGmYHm/1gxt6MnO39BodC7CTxjLYeHg9xN9efiD9ZpTyTuy0w5OZVU3r+jc/pk
hBnvUaWKP7tiT1PX7LVZSz7+hmjK0W93SSwWNr3ctWiDOVf8dSKNCqbd3/lB24vPgcbDIM/AVyN6
0fW03nHCyBYSSQ+l/xYDHZ2xkirvWhynVT5NL+bqjvtbWHS6DJ0Okg9Kn+2Gq7KYCDNBGR+LObGc
8PzLX0bTaPzJ5EQXU0T83CC3RsSyjMTqiIgDzVVmZJKxupn8qGTTTSM+ug1EIxy/uvI4DtnEXMtZ
r45r6XPlwBOoAIgLCLygYo4uj9xJUYL1vv3iTPvjgH4CwtHbVcmr1r0IUIzMWcUTlQ3DdQXVXSly
6SOJDlOVZkoerM2Z69j7rZ+33pD/hrPsbfsOh39MJ1aWsvju6cP9+BYsGvEaJab3zgStftWGXWnF
/gAtYryjK6RYWBamFUwoDTawFbQwrjvz6+lNx6QLKR2qQzinHrSSgAnmsWHQVmF12BDqQp/sSVKI
sC+pb8WeECGCZZVc/TXAFXAKQCA6KwKNtC8mCdA0/UZUoT8l7MYrUyH7pb9Prn1NQ6gisZuGCzLp
DyvuxdrLe9dchoDbIdSN9Pc4PDEvMXu2eqopA8/hHjJvOl6P5iY+RQYxk35cMDzCCYQTjle1If0D
9s/wzBUjZO1rP5cCuQriaSFLJcSbKg3Os4E2Dtb7MjdxFOoeaHnh5IFISMOWRrqBFkl2Q5sdsvSF
X8OmaEwUAWCRmiA4gCFZHpemRK4d1aa84yXj+xAOjHZE44i1DBBnYuS2DkXaKNrw7nM4OTFZXhF7
Lu7+KE5/v3NT1jAESqyOA6S79c7ihInNQU0w4DIgey9ATzUv/EYS16PvVqMSIIUwTtQ3ZVIPxEYp
Fb/tgNzCU8gCBbuSiPnU8W7fV43cPvp+5vS68RC3miIFIilQA0RUG38fZbGtfogxYWAsmrtxQ3e2
5DsQlEWK2T1FP5KLIhcIQ4+w2SiXZZY+0q/NYaVvlreWkxT14IDJgHZTWrSouOED7t5VgXQTSwVM
LS0tj8pf1TnqDVFOwZPTTl0Z0BI+lu5xczdlmwZBf4IiqtUP7h9ME6CaYLMg0xhGRQ2fmVtv46QH
oR++SsRkz0a/H5iiy4VO7IRTfRwyJk2hnH3RFc+ySjyU9I8Cvjgx5QLQi0DTqn+VXKtPAIY25uo9
sLzXU0Utj1zOiwBLFjnN18FWIN7bwMx6i9wD8F6S+CxpBdYZ+fJaf7CC2uFWx9qiFW1zISTd20HF
uWU0D+BwSueXFUlpirSCuawUliSTdwhWxeCzn4mPVv1R8FBXsgQv96po+INB8Ga5jnfT0dvZjHAF
zGQsHTqlViaS8JSzr/d4vDvul4OFaYqAhQ5cJL5TGGITjOmpC8eBWdeiQynwndNytM7/4iXX56Xh
+Lyxs97fR/XhoPfB1d3S+n1+G7KaWKfnMUBrX7sYJsXj5gPRFFfiqb7zDgAeLP00H60K62gIXGAM
I4/xq4Iit4wqEvvK/JrmaGYOme1OS3Gd13EbZLAPa4MQKZ4ugProYEPzayp4L3jT1n3pPAtED0oS
EdAD3jeovXsqjArAaSD4MKhPTXxpWLK0lFemlh37h68JFQQ0EAO88EgG9EeaRxavW+gwuu3sqHjt
YzZuN6niyp4u9np0yMNieWqlRXp6kukCwAO8ADxleGHH57C9BhCMR8Mjl8bi9dtrlghcMQFFL0gu
qrH3SOq0tAVPwkzernB8kHoIfTk7n+e+ntvSpzaNMhzQ/JHRZgqdPk7pMMWidW3CjcIbYPl0RVkN
rSHQvpYQ6HLnVKal9Br+oWWeq3HD5Z3Fy3LYVfjEXeFldgxhRC90mrcRC/nhy2oFBSR19N3j6pkt
UXBbp6/QnPwZin4vCeRAFuWKj5FxgqGd7esBxkW094KsSFh3QgLzrKBpOkQb7rpyxEkskR8qveK7
jlX7HjlWmv9ySGdjqEsTHZfBHQfJf/xEES50Y2IkjJYBjgCjLnhfQb3uIqi4YdK4E5j7Lwku33op
aXt2END6jRCRKu7YyctlrDRBlu3m3TpAbrOomo4TSkdS8QUCvuHaXtyQXOImrounlAcUF89FLo21
EN2cOx+kTW1nJ+odFuokI1KlHj2hDwZXBIZM023BTPdBsOe7dzuLlnPci50N2fzyoxHhOSIgKqNz
KL5+8vmST2VMtwbvqhfjYP0ZnGyQdDjH7AjXQBTjqCI/aYDZAAu5jhaccAgY5Fo0Uy5H2Lufjuzg
8g5zwp8Y91g/4ew0qNGEJ0vOiPkqPWVTk6zxmyIYQX3DN8oiyq9fM02aO1fbTwkm6pRM5ZCW1Uqw
VhXj0ja428VnNoOp+Grrj+22KELFdTh6rG4ARSqHhmgjfGcH5xBJYmAm+mfeu197PPxTxzcOCX05
NEpLp1XHYA0oS+pbGD7s+uXnysmirym4B0T2mQmhmqm+qqKJh5fGl+V+CJfecbZGghBrYHqXtckL
cLKlDfRuQzkC7EXfZ6IkJB/2vtGzg8/Y4m1dpZ0RUEmUt5ysHXVcyvt/VE2ABJaQHctGcbzH6vAu
dsEbIK0b2oBmVmaVftaQ0aByWpxvBRbSSzyjR+xxMGPfEobUnIuVU2t1XW8HXZR6wiU257BBeTTr
JlBzu5x/IcbX+OF+Ig8TliKklUD4zZvTjCzJuWpSs5JpEKO+vRuidsc1gEhofAjlXkYa7miMT7eT
6pCHd9wHiubo+kighYiGsgZYUYCeC6qM1wzWrP6wB9d2UWFgmemqvMRBbADhoalOwFVuGcXwTEld
whfGBVkeoDAlrIwgF58nUv/RwXipMzb0YwDTyCiXAsojQH2/Xxn8M1K9DYb508ucjE1xblqM/tu8
7w3dBE4xmWaa0YKJ6Hwh2zi7KaRyWCsDaNPf/hwM4IZKm7rfEW4qzVH7UxRrbm16rkmSiLGYDWPv
L2KWhK6KsBteQVOx5LGxY8BlKl2dAdiDRHxHo096ipyqcGVVmunJ72qoZ0h1GeBlGcNWk/M0YC1K
i+DaQmZXiffG4QjOWT447h1DL+myCEJmqqvbxm9x0lFzLjGm8DlslMwB2O6gOHP6/evyxFMy4QIM
Ywpm9QZbsVyhwvAFAwfbnkgW/oOkVJ03TZq3BW1slX2jmfYiXSSfgI4nC2Glgiir2c4DL8XblMgH
BFeTufq8k6lHBXS7LKMsvaWno6j0EY/y7YueWlBSMKxwxWKU3UZvUMEg1+JbJ3ptEP0DXexEYNvm
SN2qv+LrahjmX4HLDCEIHMRWFvJt/PBwfYKeKX1fvv9IuaQ9sTb/8gWOlgt/IWOTt+l6SpnHfjUq
6okfi6Pp2Q52ZpZvEH+I6wA7CIXl2qqbIHIgY7HFjbLGywpO3oFI4aZRh8HC+F7WDpoj4TMIoLuM
OmkKCEOkbNYF8FSHMmlsxcpOshT2zxdwswQI454M/Av/NeOiiq9AlIQhaI8Cmd7QS6QXOL/9U9DI
NUsy0G41Ukt1HWlZ7xfl5rWEkW120OHuGlG44xyptkFW0Qx6qX4iko6QNm4+Wush021Z/yoBZfWx
WKWI6iw4d4FXEohELPfsOzesqPQHC3HAFSE+ORkbBnsqgIkWyPRF3MRn2rmJWFDL9k2fUYPcGUa7
hvvPPAAqVY6YYrkVi4qLL5x1Sy1FRLjQ/2KoXI55nj3CLq6TZI7kA4sdl6cihaAwLxOXjdXabnl0
depx1i695r10rc1sBF3D5XhZcQkb53X0xjCopEGsII0bHt/spZvt3lQ+eawEZLM7mHcaOvuRfF9L
KcZJ0A6DAEh/h16SipTjfplsF0PefIpLkz4IssiuBcmSQ8MMCmSXAACv5VhyVnaDpDJJ3qz6ZsKo
hLZTdXY0NrJHiGs3Nowkw/D0Wz/HTQP8WXUWOR7a/OzhfCu3ZWzeVeI0iye8ePVzEA2TT/CD0oIk
sTY/F22hJxzJFe7RhPFmYk77DaSXTozxCgZXNs9hMfHwrITel33Hwd6qYxODnRKLvmuCkCUfCMR4
pnoUvIEQFPAtuTOZtE7iOrnI59nzzk+IHOnrd9h9mQOQz+5Fz5lf58Hs2uYOZ9cyWmteuwcQH5Ge
MK8tYKzfcgsnSK1D6mNpVb4Z3g5OEuF4cCZibWbdJjBFbVED9quYM5zmsiroaZSz/nrhsqdlEbbD
qIN9yHZ+XUKFcFw4Az1Qc62+Vm30vftKmD1sKRrILkey4oQCLK4PGJWjbbXSLv0vnPWYlQEchfvh
E/6BU/dNrW6FJmfl9ciCbiqpl6nwJUDoGoEtW2kjzylOrswp9Oj+kXRLbvrXXn8EijPBRtHGn2HN
Ufm7B4iksH7prHRHYVHJ3lISt47yE9Wi6uCY/ljy4uFcMlE6ItGv6/fNYec/SJenm5yCHudnL0bB
AgM9ueYg1MLsEOLQf9yyAYb18lMg/RPwvOrSfG9CT/3qerbJSe8bKiDY2HxRF1QDY7uEJtqaBxAU
DaGU7sc69EKLEGnXChBwvGq1V/8Vi2OHGC94HkyvHdBwXH9VjtOC/zi5XAEb/TuCY1+UuMnBEBHT
3/BsWlKG3HJI4Kb7tCW0k1nwVAlpl3wm+kyY0u4H6zAz2+conJgcmWm1WAexARy5q9MNKSCMg2jl
IvXOejd5kckO5fGu3HnWXq0+fIcc1oBbNd1OhckRp2M0e2MkiC/VO1phppB+Y5HXQnJenr9yJ6Xl
B5WoK6RTpuYe6i6fNB5aSaAJ1QrYVVhbe558GCfk7OCLAtcgj36h+pUUZGjH6HS/biWLVfCk+dAd
wSMocwnZilABzQyrftZ3ORmXGZQsRDCFNQx8vVWbKTMGLH+Od2Ihsrl/YG9PDxqHY6wqlepsn0Xy
vyPjmD3lcnUHFA8yIIW6qO1S8tmW/GrOJVXNiswKd7XvnuqmvAyazUKLAFB8DJKKzeE0KaIP8k/I
kK7Ymhy3MLqt3Zn88Il7zcAddK/vH3AukbfXtf+UY/po3rCoK+LZOicmp4s+4MtENKbh+WWS+M8l
ib2DWryoAMYQcjaq+7XyAYqgGzTD2taLZ6ZO41uN75mArBPLQXMWkCI8agjL1tLSae5OcBzjsex2
1In/1WzG6JG9K8ZGY3NW3QKiNrCuYpjJ3iY0AR1YtsbJvst/PbHcArbQqL5WSqfKOjPUX7x0dLkU
XVNUtey+CdrxlPTRvWUj/ax7vIZSTpO3K5BwGxcxANeQZa4GnECclbtJDFI/rjJflx92vpmZEtAn
x7tcITurGiLwi9BOIkxpR9dpvn3ybZjZcR11J18WLfaec1WltfNIsfl6beCu9bvqhWRvr/sdhJen
CskA6oDorxiUhFzmZbSNe4iDA6lZXFeq+lDZFZzuwIaPUb0T3xnc1oI7f8t886xRnVG2+aZy/h4W
HuYXsSSlCdu3bTk68C+Bl2RJ4YxXnpUvN5YgmbOyAV9ESuYm2lBe+nasLMzgUyKjMBB+ppNN7YCT
HXhkPsCTomItPdau9Q+pzh/dg3lwQwmy6vMcvYW0tALfsLbE7Fh6KmkxuDMorLrXppFg3s59y8it
kkCc+O2PeYxGWZOQR7P0qefWmuVO4qb3N+f75kJsklybCJSXB/N7CauhXJi9qt7+LMRyVTL0BnFi
pKXyG7AsvSdTugn40osfi0HX2NF363Yp6OUrfmlFIJ6iR72SIPL/QftJ7TDvg7hhdVVp/EHD1Jht
DPjrJn8XsPG24RYhyK6Z4iGEL58JcKh0iz72afdCzwkbcWtfAIppVfDyws6gDuL5UBk+vPECihv0
MaBjyD/rVmtdxex8DGwsYM7lmIlEF3VtA/Wbxorqk6+QtZT0NPJb16+AAtjS2pnSDgaQ6LXrZocP
anQqt1Yq9Y5/dP70F3D/k0RO6i201uJ06dlknDk5SXvaZtH9GHfYH7xDIc7DFcpwNVrh3XJNpkNK
lG4CdFEG33HeyccgYq1xlBaZMmRd65tOHU36m3FxsceYgGX0Kj4UJUAvx+Dx8TlU3xNTNyOYsi++
/mOxMnanl5V79STabVqlock7uKQNt/kFLiPo9XrM/3ieFCotdL8rQsFlcT4VQ2qdKCYMD6wwleGy
i+FM4GI8fG4AgdFyl2To7UbPu9Zw7pnypQZDl41yS0oRelZgccCXQ2an3kZUv5qcZS+bYKSwvORb
yo0jm938ERtdn0nG4nKlK90PpSlSbXiUXpnE7/zRDJ/fGzZMWUJQYnCgsLfGLbYlY+KbnYzp/gJD
iGShw44GgZVdBB3NBqOY+o1dVXmBBjWIkLvuOsL012Sn8GjbRw7aVk3SroPXBN8sutXuCRFSUCY7
YlXqPCw/uQ+146zfgjkGzBIWJCmNvk+z+zSQWJSCKaqcDdplirYUncLx4lb2TrUfOqiYC9l6eLm3
yKZ8jccUWCSQOcjelP4gf2ycBsSjhOU1EGwdeZ48FJ5p3urYiCS0poX1DzOwT3AJMWqpPFo1eCo1
R9n38gVIiJfQePdnmF6FM/+7Azg3lYYoCTsy78BW9niHb7VxaXIepUu4hT/pmm/o88VDIrKf8oab
PwwxAmTAz8edQMhbQI+9kUwZ8ZnoVfK7jT2gfEQl2Ro9zSJSm8fHp07t+E4SAPTrFSrUNNbUz6/c
uCYNIUnFfDhklrDZNHKpebiBz9imnKYVInEIpenlA2IykO1cxvWC6/pAvtuD5shAA2l4o8KJTglD
dbDfrzLQixWe9btaCV0DP1qOl2BZAYfDUE8dzIxIB1UP6A+n0JyEasoo0Z7oIbbKRHH2SKvULRzU
+Cj6Ig0MDaNmO7HGPZ2LBMSXM7hGpCYaO6WQkCFGpn7xgUXnpn98WHusKZgEEIOijHvaWPR7DEOr
YbNPPygti0MWqQ6L1Lyn4FT+lG+T2KvJFFoTjjMIssGhrZGV6e9QENzsZy0Hs6K+EEKoy0pf5UEL
SB6sdvIGP1qe0EhjFhThmcq4pr+s+svN0LRJzD0vu97bujI7Lz18HcWNWLzwQmAPjCX8GNLBBINA
plZBSx7QjFIAJVw6Zs4m4QwD87rsGdc7iLILjUzP90oj8Eh2mM6uE5szzzLxpJ38V2NvcT6Dcc+7
PYA0HZTd517fW55C/W3w2LG8Xt3sYBI0RIIJ2KUXgShFWbm7CQSALkuFAP/zyUABJkytm1lzFjlo
ruPm3ZZbxZNkAegkG8nKL0yE8PPgfvUYIgx7k+Ry3+L3qXSHf/JdvGEwT94DadQtnhID0jAxneLr
6ZOixDUxIpSs7KFZQWcOAk5+jqBsm/EGZ+uqqYoMpK3qe0SiVVUbP6YCuugL9EUtRa8CWKa91wWs
GQJDzyXXNoliB3qiX2+0lqHDgeAL2vVZa8dyO/hsTF/ezTwuQA6XFetU4Hunc+LugL2BZhKj6W3n
4HPE6Cl10XbVQczpD31f2PaGXt56S5tluwkuNlXAckMDDNG6dDjaCiJlycwgbcIfstJhi8yI9WwI
+IvTp3G2R2ywwjxwV7SBZpL+47L/7WSVjro5n5/bvMZPBO5pnj+/8uaoqB0qSLvzb/feU8nXqyFp
w6bJWXF1tgIKnHpN452b9Haj8omV1DLXiT0qGpTGo1xFUndw7VOzmYesfLknpFD8wUrOf9Yfh+ju
OrBygWvvSVx4VKtfRxrO6Wwuwhi8oHsvv7wfPI3PrgRwKvw7dTCEMOj4GJT/rprUILWqdsyjSjGX
JkSs/VCCujE6p4dIuTaQFigAZE3l29UaA/ivOFGpRyO9IhSVUi+sZMxIH3D5TdniyNBo3GfM4JuV
eXtY1O1JbhWOkMzCjPbb0KiOH6+fhjls4jIXagPjU7SZg8hKstOHIaJSE/HTd2OQBh6gslzJOgv9
M4cxXqbw32VP3NlqCYrai7gAoocvxxe9cEGf3/7RyZwa9Jb01nelPwIvhy3qCgl7IImbWpTHvNZC
TnZhKF+LA99cCrtwrJErEZKDKHdOvar2+UACadlbu3BE2LeHJ4mQGGtgSNVHPJa82LuCsS3yQ3Ur
pEdl+lS26jItRD9oDzeQQiQpcrKyXYoILdco5NsEH+xoOPD7GzolKSU19lrGn2sr7n0AxAKRherv
UpfpUpnTeqJ8d/KVYBiq2eZYqwQCNs9dCKMyaXig0+ZXKg4mEPfEMJG/ntHk0leZOwIKZ9VYE6NG
eGTXlhFkGSBglaRp/gNdUImUSFt4pIV6R19roBJdXEUuEfWo2yJ1sAvPDdGCb6OGZP0e0ljeWnqG
j9S2q35bM8eSx96M1XDTYX7KVshQQzDPvkje9ymRl1wEwSR8z5rdPGa+N5dOL6IHUHwXAKAOiIEh
M4yY5X/2/PaGSJWRPdtWE+312Eujh6EwPkRTR6sDNejoFIsJrXeIdE/i1SsfRLVGb5EvMIpcGf2Z
SjJNHVilBapF//xfNT56aIu0OjhDSXqyZgdKsPa4vysuuFHPZG5vb7P8T67DklJPPCcyCg1Q7yPG
ghe82kchThBrHXe+8plEmPBH1xFEAgy+TB9Cproalx45XU91BdshDFQWPbzffYeJRxz1A/OEGiPv
XeYPVrC8eOrXbl4ZNhBRbrb/D821nzPhn+WDvWgWagEr5pJ3TduVjIFg7dfbZ668RcfX8WetuRsv
B0s95+soLCpGO6cqvL23APhZ0wOZaRWnfpkdlfC3KS2rrMuqPy6De18ekfe0064POxF06ma9eVoz
xdPDhnNc8e1YC7zI4ptiUcbpPwfmc+DzuF/g7r45//zG+sVLNnXCGB2osSElybktAj8NZU4ETtAr
g24cY18dwcOIqCdGHhUZ3HOPSQLmBbw9HPj6G1G+iGe1kmVVdyRL8blTlLmXTBIwsjGE0aLF+HD7
8FiW0Yp3ysxZnx/FwFnhaxG/PqIkyE+yLS3HWGzaAWnkvKXUVSrt4u88pwOW1fmc/diyOztnQPW9
AqGP7pq4zxtRWM8FrGWJ5rXxghZzk4TRxsi2MAJzF5lrJReb04PHkuz8xaz7jYRWFjqT2RIqDQAK
ChyGIkvKK/sAGo6F1HyrQ6JLg0Kmc30EWVDtJuAKsWBWgNbjaAxS72gD59ThqS/CwGqAdwaXMO1d
Uoct8eeICTm3DZ5bIhsXk0Qto8wExAsKiOMBheCc1/tmXnak2UM31TSbcm++llir4ArnnU5OCJn5
ogBkLenzHZo77Gjy8bAW+9suQRQMYF5zIp4zah1orMt1VO5/y242uPY6/wb5NhWWRor5TOWxV5vf
+xn2h6TYE/gyz8S5gFz0PCsuICNF/X/aZg2CWNw2p9c9GHGfjZq2ts8z8glIgGO04lwGAfEEoKc1
9DPrKi8SOy32OQU/h4AxoIHGQh9AmAQNsLcaU/T/9UPwYQzRyHvSoX6ei6HPkMp1JHY08LIUg//e
O3lmnmuo2nxBlL54JKMaIRNby9l17IOZWbh7zrajcvMINYZC2sJ0diGAlylfsIPDbU+VsUc+bCuu
UEnCZMjHi7K8be+0fxws3Vka+/KhSIE5RxN3SBzUzsvFmu4POhI32YRLW8OcWHBEodRd2F4oD2Vc
05xicU3SSIeeC5Iv+ofrZ1iIl3Pc3XS5+KOReaBdEKZV2pFUWI1bgfLQ0vvCSI1B+ZGZszScJyKy
3F2rL5bbmjYx4JOp++azjsRrDRZGUYvIK3KkZxmaBfKyYas43J6VzAFYkFgzbri9A7VQs7f1te7G
TDHOj5v19+/p7rlBw/rooHV/RGvgh8cBMXm0GiIcJ3xRns4GW0WIZnHCv4chKDnAT/o1bm65gspk
ll5Ar/Y0HjJ1ywp7VBQ0UwRsdtchcFoDb1LGya8Vur/HO2mChCRqm77Siafff8hftCyrgSrjHPgp
RMwtIU1Or4Rlob2BTYsVpNNzzADUEEkUzr9xIkobCf3PveQBgzqKm+xJB5UghYLsfiVgXnqwO6sC
2LBJyc/xQWmrneyIoRfIspDYcpJ93Zy0ax8Oj6wN4fCB3l/mmxhq1iaKjc/4GP/cpAz5+GCHU7VU
h/cN34nwuCjeKtzMcIGRnYfaX/2t5lFq2NkeGdTWgyeA6GFMxNn2RyLRbO4EwoV35tmfDNiyeaQD
gjAcbO2ZjlTwJ0x2MN5I6yAxIvkIik/kR05cmhkzoPmGmFBZTGJPUoWlTPNc5/BnCOjdvKwQZZeR
2pz5luR7DgUL6jR34a5CRIefLNFbnGt3WJRj+WV3YGjiiT/vzaEKXH5iDKNe/avTHXd1rl+CUzvZ
DQIx2Tll3RK41iAS7Lxv4bTyuDAF2n5/GHw4c+v+ZP0qcKWYqm2RBixT6jouscZJQPI2KEw2XqGy
zvjfwk+NhwNXYWYw8fRQ2uMwHHPr1YvgNiGrN7qchG4LveyZ/FRZ66072HG78ZjCBIhr1VAclYM/
odqYIt0lFdYtVr4U1zKyyicn1CdIbB5b35mU9q/JfWVyh/QfqtGSG/gJYOrmEAZwB6saJihHNLbC
5KyHppytAaWVA+FSPANjDC1tHOrT09JIX456TfrPL9TfiTDcynO7KXXt40QxrDjcJqHnDvCqDe8S
2O8MaaESV2WeZHIWEMdxXnLgUt4WCYobkMRQLtHrSr2D610mE8gWQZ8qY55gqNigJC8dE3qBkgo9
aNbOIARrFRTxd7imuzvHzrrqWWSvMNjxvJ7NY3w8P6FhrCyENMRKnqLVYE8hP0v6xYF9/VbJwgPf
K2Uy/4zAX8vg8XXj+x/rCwBpq517Ly5EjkmNqorVcIDqnOI3GTu0Z4kWsMC9AB9/jACCeTenR71c
7JmJGE9thqNBye1IvsQRwR9cHLBNMiQQsNaxI7g9LXl1mERHJ/tR5/gGAAhPPH7EgUEEsCFZzakR
t0g+vDshf544rFxrzLtGg+tKhOeblc9vpkCxzCvaW43GRPdQLW0FI7IhbkDPI3FXSioHjn8QF4Ka
/2aVqR77nuGljWVyZVzEUeqaHN42ULojOraHDrYd0l96f/WtTPcDfAV7AZxRU996i7ygOQIgwEm9
5xGTSxx1JTd4lNrQkqIWQCJg4PYuDVP+SX0wyMjzGbMUFSWXRaXi1reNEh0/H9mTCou32w4bSZcs
5jYhYGC9TDvCCxiDWBiqzQwSo4I88mUAlpQXKdQ4GE2cAFSUFNo+KL/7e2q+Ig2Xuyomn4FrRiZ6
41k2W7lZSyQVQeH90Fq4YGXzUmvPyhhp7KEiiO/2/AM7vRnjHCStu8xMMbJeBvrxVFLyDldeHl+D
DDo5bJri1oymCYVl6oEVzIuagtS/BY6wpwz9IMv0bzKOfGw5M0dRhH9cPqdCwS3yDVrqKWD0mTBO
fSklF9o3qnzKrQq5R96rJI87CcLbiqA3bu/z37gHiQ3TvLQh4r5XUhG5a0UWOV1dpVXeAGApHC2J
eh/WakAHEWaWSEWYyFSxzlsIFsQ5z4qJFSm54S0zqq3n33eJgJFiD5997/+9kyjRtir1v3/MaV5r
f5jOj4yLcx/LEm+kSRgK9UT5k3zYDJg2/B9DL/1mg6xmZe9S1tI8gyRoy6S21c6BXCa1clWKmzT3
b4vpST+wgcKXNIQ/uEep6FQhejbOdXro6uNqwB69yGjfcnlZe5Qd4bXAuGwgwxggHZtK1dSSA+HP
znMfyXO9K9GwXTzfCbJ5NJ9OMek84scv0mDUyQsxu5kU9YpVe9dR4AVOdn1g2xQ28G5FTTfeC6Bk
ChpofJWx9utNXEiZi2Waj7K6gW5UlpAQEdfeQ7vRhxAkSmh53hEu250FAKt94ogEXHofhNa7llKo
MRxTneEEb6a97SSzpGPC7QheZpvadIrhm03f/URSCZKqGCQZPqAFValddyNAp2Zb7D47yVXb08/p
nDhyge3tG5r52m+Y7BdIaB7p+SBZnAuIFLbLTF8PKjyvFPl6VVs9dBGh5QET49yc4sIPP5Bpzlkq
bsPLoXOWbEm0EZPr0lX1rAmt+eAyNATvuU6QIBY8UB+bKL9qzcLyj2fnvBgnMMnLT63A7Ze+EY4Y
FMh5/9f24lIJQEWxGyOcxD18+gwNGDCwzq1DKKKYfDbnU3zJ5I96Lk/aR9HvRuo8ygTjeQWXeclS
dl8Dje2pfK8noRitliL9Iu8MurN6MR/D5Fjq0eTfAnw0T9ERO1fhRMrb4zBa+vBlG1fWso5I5QxP
WN3rf6spjiW9soRBMngzYH2AsqrFEcw3QUPHmfE9oCcF5fNd+Iy61FiRP3Lu8xGqytWnL+YUoced
xv7jAaPjW60kLu9y7ZPeTqo82MfXFQST9dQV7oXNic+w5bAMlnm5icJdqfyYN9iQrYp2t4p7/tll
vSGcdTxeAQFtDY5oAbuEnj9tIlOZufIEeXc1xNnbyAOkrITk0q7oJV0niusxdLDXq4cNQe3GsHHQ
neVqGUpueD3s+Py5Y4J9/Oej3JSR5AyYh2NkyUfzHK+SvDyolhlJroeQUIUJ4EoAb6XlcaZ+5/qb
AayKFziYZ+vzVHMRys4F0YbbyATwYUSDSb+EvF962FbAfQ3lujmlTmHram/XF61Ywg+HeiYWoBz6
FuPuVhIoHlFWeSdkyAOFEfVB5CRlxTZBMYRyrN3Myv3DGOg2eYYqAC4I/LAe6SamsZo8OOjs1CQM
datD1bbBA1AU/otJyseaG6wq1XLXe9U1cyNudc9Aqu4gL52YPHOcO2AiRa+I9p3T0pggY1LngpeB
2naYQ5QwXp1BaWYZhSF2pRrWFK6qEVb2RcD8WFInGyB/j/CiCw4VyUh/HndEwzZcSFjO2gq5ZgNU
rw46lofs6i1Pcdfnpe+M0r9BCOst2RJEBo8TZ6X5WXCYEGHoxUpJhf8YLvPFGl18APMelSn6q1F7
CEwZM4RAUGSW5l4/3WWI8MvbOSkoGWj+G55TvwvVIZhzlgzcdIBFdIEt5jiQRGlb5tMe9ZJK6sF+
lCmf0Eqcik0YOQFYlaELeu3Slj9A3PlkP0eJECkQzuoYxkTMK+Nd7uDz7R5jEACjiyCYh16kkYxD
CQatEO3nGbQuwm6SpcvKExwpATomdeNocymcYKQ5EZ58w3w0hriuGd8KhITd2pRYxHMd+JRNsWiL
Z9WAwD+S0tWfE/cQ8TklZuzOIY7nw7/MKPiBlQ+C8iIKIrDl/B+D+VhcC7/aN2Rt2uT07z/WZ22V
ik0lNighwiDo/oZ3qVx+84GNmnmgwbt8wdFY7WiJVLeWo/0rOuhlJ5zSz1SSLPp0egk/zGFlFRgd
IqtDW2om+I6v4osob1enVE4hSgZL/+qvakF9qink/wJT1qhgdN1qkPaHkTf+fvcgFM1TR5lCgL7b
X9jBkgc+2RvacpaeUFIVPPPm8w8VeCKUw5tUId8mCAMrjRrBlS/vwoUc0em6TvJZqeEVllTui759
EABCeJxAx/1sUgbAR+ROFwiHMk0WCMhqV1+3pPYLFSgAjX6JsfHp17gSp+YGlIcnvH8ONFtSRzWE
0aHckqjXNagWE+wTpa1HRWRHQ2eThwMAipKaFMwfbdiNv1zSVsWIF3cIJE+vAxm/5fhqQ8GzbPyU
Z3kUWFlMsRqoR0GMT6AYopoXW4sDlNbQK4+2wqniCYr3NQYtPYbuupznxS3g6KurExhlwMAVB4Cz
/x2wWP+GzR7h/wjmR6Scq/DjU0f/5dEDAzBtQOpovApYW50DRd7rtewM2PJK1Bv8ps9oLA9+/qe3
jJikzsLOlvTOlTTa+z691g7Y1q1YMzH6Iy17DbnVbadE9HNG0C6rt6lvHvwLE1jhNYpxFLhtPvTS
GKNX7fIHEhsordE3ec+ZMccC8DENzeJruw66V6VrX0e6zflNqGgg9S5P2FTy6T5fQKfKgD1842xR
s5Tda60EMctIgNmawD8ITEateqipsNIk2Sf9PxlxfLKS44Up8OXX1iDsgO7Wrxgn4fwPy/Cp+k34
4hdJs8wKSOlLGPCIhrW/yKoO+D0rjzINWKu/QPj8KqDcCISbIl4ReskCmUkCU43KaTfJGmTylLV0
Y8Nq+YRdEr+6nNNgyc1x4PSKwssQg+YVdc6LprMaVm+GyYcuvpnG7f1rwoGqVHaTGhfTdrlwDK4h
P0OSlM2iPp5jzjVl6Y8Ss3EjaeAsUvBniglwzTSTu0PKrC91NZddiKwPnTSjDTrEeNnN+vljzYVS
aUTLscH7OYj0c/lX8oB1jgpbu9QYD8APiNSKgwd6ZbeM0mo6Q6i25d30eraq4LT9cGFDeBDHc5QL
GNjG0FceC4wl51URW/gzEka20cNoJJ7pr+PYBdgEo8Xf5QnBqzMzJbDdKqLEOw5/ONkIL084B8wA
pEkXqEbyvDy+baKkfMaIorrOwEFK+7/9sJuPNu8X5Kuu012s/iBsfty/CdMgHS6zrc31WZ/GzBpZ
nDxNDoZ+sbPmGeY6pZvUIAPKmZYYJ+JFUVwk2UqmhpCKq2MzLXYcJ/qe8+TyaV67wtho0Y9aXIXW
BKhWYe83w+kC1+mK/UhwuMnV4CQ87bwpprmnKMYbuY30bYR4RswHUl7/rAtZe7+nwkYd0GJYXwbB
/2nqPlzQhu0QQNrDIT9elPugEFZ2ctS5LW3M75XCt8mygod6G4KldjVlk63AUHw2vIohlDDnyFPV
EpEclzlmFt5YDOwFB1c2B3Pgnj0A0KnOB+xKnLyfx/LLewf6BTNbn6MXf0j8EIXEiGrVUrIdlLKJ
aIbpcW3czjXsTGqH/6SBvz0tLgE5sEwWtApMftNmfC4jWfobt8cX3hnm+E1HJZlb/lYY0xqIvTgW
NeCsjwNji37qoa1aS2yBJXHiXo3kRP76a2WOkBzjANa1lKs97M3Ery8AYtA33uP4J6Ci89BK73GA
2LZFOBfqx9lPhL3eaRpoqxc73yLgpgIGU/ECz1F5zibuzeb3vkUPnRgb3ETeUGesTrI5/4ycIa2s
N3lLr00QNfo3z/W6R83gk+DqMFI67me9MNadxf5Q92DCE9nHiOOS5RNmtovH7JHFXSEIftklVYbD
F1bhdN/9lpJrTgADKgF1Ev472ikT5bgXJgADAkORqq7+Jg8nxaoYsFUyQ3AcVpNdSmlzfAwF+pzL
NebJVE4nWGR6jMFw1HQyZ8NqPGl4jxwGnZdzyuAnnkl8yxOcERyGbn/+Il70OutVbJsNMcvVAP0o
UXuZAX/eGLlzxIQzNDsXEPlQc6Qs8kSfatkTiOxe20p8+tddSNAK9dGdrqLTdoDuJPFsAOnSfUI9
ZPqr6aIkIWK6oaA7xhJBk91qvfcKmmcWFq8Wg+pCv5/S4ZTKVSpk1TJfuOIWmDJISGuYnt9Buqr6
yTvoR5o97JXqVQXElZkL4Q8C9ibD8Ol5WsmNkOIYec0qm07WrXshfV/k+zlenSY6cobnjGe+TDeZ
/24xV6bdV3VX260QBpw/CDt6aqFwdMHpUooQTqbvPzsYeUfnoc6IrqvviSmf22lLVKzOjGb4BKN8
dJBVABVIwnMZGKePgEleKtDTIgbNuJJXvLN8W+DZP4d3Gejeoll6fRiUbYqDqqxOgVt45IRG5/Ks
wXMzA6KsnFSs01EOahhyh3qAZE1yZYQS7GnIchTehlO+sC7P7CdYmDeACS65l4t6tJQ1B9ptitFb
h9oIS7fzB3/ksw+PuKZVb8NYl1Jc9vPCjCSDisCcDiLjhdDiG9LRlD77WpOARtQu3B7WPo4qgy/M
HvHxIGvZYdsPJGU0iDQamZhBNGxhZWVEfCfZKBLV4+rhzxPAxuDX28SES3PlbaXYSBt1B/XMqx73
3LrBvruzCn/lZNYWzjot9cwErXr4ufHyElkZOxfpxp1OPLXP/NzvwWQ3HB+TXl9iKojawiMoWYS8
XGx3R+cdRH6BiD/nvgZiL0PZU4WwCL3+uUkyGYo/ueaAjgBr6UcxJtYfdKBcizARmBG7lleBF+Zz
4eqDXcm5rmwcCsUiANmhtDBuCseE0Y9TBrP90viug0KvtX35YVjGIE4t6kFQhg9gfhgWXs1hhkDD
e7iIJsIzI//Rc8lvbOMz922Yr7/p9P+AVePbUzJMn4U9Y7QnKTfUkrQUomnWowwtMGwccvsOUYLJ
QDV+pEdxeH57HDtqgYhrhUBfl3ECy1AcTCmvVwkvQimwr5zmOvuodOzTul1l0eVa1mo72WE510/q
R+3LSBCtDZtuyM+YKrlUIYXPk+omoRdMAThhG/JjZm+c6wF/ItZPKSUj+sz18i8nxkMN1JJ4Alvb
hJayg4SxpnmTTAft6Ys5ZgcAysLzc6LLUT2rcDbiQAZVRPXtJQDXN1QHVjkN8v0V8hb0rfYMicxJ
TBJx+cRY0eiGYQeD1nwrU+NN91Xl2a7jQL66rdcNP3F8uFDIVv7V4RSgLCUQXTOD42W+ksZESoFf
YUWAIeWhSbfpD7VjmNrpr5Moy02Hx1i/zbGwkw3x2KmDXq1VlVCYtxBSrRDZ7ScZG5CbISOws7hh
xxeoYj972B7ZmIhvOoO/8piU1xfPpeV9Ch/1XATs/qRAyW4BURuyzf0zX1fpuzqo3JIYez6TA5KA
KrUkda5U8MKQCTmgxVhV3Dghduf/mRMz517Vy1HBkBeCQ8upBXPRkDL96dwaj3zbw9gGczhP+M/q
mgFwnDmCEiqOxta789WaYYeWorXnDCa/7Z8ERsCtLB0MFzXsDYed01feAuhVGv/AzHCfVC0UWGAm
BNxLpHSxmOlaRYO1UerKRlx4ESq1xymJuZo2lO4yvx+grSmvvOIcWbnIMiHMvHfSPbSd04dNfWGg
fxWfY9C/VorQ3rd0P58nLFG7ExZh0W+LyLpwBDcs4peJ/cLVDytnd6eel6n5AC2X4IpbX7Ke6Lww
799q/3IEQTHdxIsGERJ8ZGbzrL5PTc9slqxJGeg78VQtsrgeecJDucmAqxuIOhVwQMcZU3vR1Gf+
SGHp+nXrwcwq9PbFRL7q1ZNqpshuQOG+1bzF5q6xJlYlyRBKXY7pXQdbxcWcfqV+gs8Pfdtj6pap
4oc7AqZpFJDFkbYVv+nspbMRk1DSBFtWBf2nIoEa3CLsz5QSdgFmTcWuTRpaZ8mOoo292yZtXkOl
du+KJ7rAIail8BeJGMXvVgT1dHB7C9ZmudpRMXU0I9PVzXM83nCJDiVybog5STp6rXJ3CV2rJyYA
gleIEQrL/GDXfZy+nLMj9K1eMnoda/n94L5EB34N7HQqf5XEls10a76M5zuBsDJYsn3EUEg5Cb30
sP95xVEnA+GAn5stFMrR5ISy/CaQERkaoklpZiFEkmp+sssKGq2bIg0elYHvnKtzOjWdnxvrQiyw
ysf+lyuf/M/HWAZwBoI+gS/hqzdg9V8/WHEqtRGGdyzBaUjhq1kOfX8P7Q90a+SNevNMg+p3gDN5
EJ8WNv7JU1JK4ZrmIO3Bd+CNdjdk2Iz+fwL8bigHKtsK+Q96m7Z7Y36wmFJc4VigR5JvfghVDAz7
aGLDwJy5S99tuWSjJOCYum1r/HPtwKHeAjKIbfl1S/WrR+2hy9cTucXazSVBMGlcCg3634FA6+aU
7AFMUlCu+e4cf5XQG79hixQf67J6+BkqM9K0S25BLXrFB/RuvywIZBIOh+wIxjtofs96pz7fXBkD
MJrA5IECH5KogWiNcx4uN10zd2R+Yli/zFBqxO/VvjirsR+METc60sq0zWmXHBfHs1CrHgaI+4gy
/J+ZZKuONPNDaRz1+vOo5Wkke1WYZebrvDOhacqIv1lC+RckgDAn9QstI+RRNIGAb+RWl0mL4xCk
/Qp7lbe9vQg7qN2gEUUREUNAnzfiUryeFHA6J6llhTC+k8V1rgwPZ/6MXgxbMg6i1z1M+7WJ6ocS
ZBmyOx+o5F77ST2grsV1ktBCw+BR7BYc5cqlNMegmjA5S1HTLLj02b2y1Oq3HzaPbshACqwXT4WH
Dk8jADcLfJHx2PTxwadSkUwOKIdTAMiWL7jrYN/rcFK6URanIeAUddE6jXWWFK6zwQgoGMNcTk2c
qqrQPaYivVHXIIQiZtf6RXJaz8OJx1wrv3VrLudtzbOXfW8eKHBqB8Io9P3KerA09urtManumOO+
Mva8XM+LsGJwwmvdvxtW3GRGNgVsFc+alDAwjEP/iEMSj6wa2W5B3Rfir4tM+HfELQXZw9bJ8BKS
CJza04XMJPajZTvA8VrmdXsNcBf88JWcCAtKPSM4fCPUXaxKK5wZoNgnoYB5BvBAKsDh+cXJrFnz
Kpq2701as7W9tgwKbCSOjq2Ok64TofhOZxICDeMpIATTtzneXm7AX/+X5SbAKFCQYfb4RB19NTOL
nnzSeAGFkW4Hk45kHTziiekNw8I1bOdzx4Q5Oa2gWiAwKZ6+suhmNc9Bl7uF6SuuU8MmnQf1lP1R
FghL+V+wrquzxFTquP4jxfMUhpgDsI2eczJsr567OG4LKD7P9iLhDI6mO4yjQo5uvQwvnWR/Z+ic
5+MX9Mn4Q4RVTkLaiC2/jwCW1cD9Qi+90cAjQWiqSOYpcoPQUa/7/WjoA6KycH2e3P2/VXZJ7geg
mEVCOCTUsWQK+ajImWqQIAAPqih/G2Fv7Tx/AfqpV8ZlfAjQpAcHpSyClAKY6wg4oTox5nFY9wiD
9cM7NKAN+RYH8WZTBE2Uu+gSWr57Ez89tTjHeGOZpbRNA1aWGPlJTg791XD2ponnVpLHBDCkamGW
XG/AYt6dyCjODkflmKfqshnfsQpgN00vtHctlwC9jiq5iBF2j1gUFcdd8tB+qk3h/lS1abiarftz
q5bV0upInUpbtAk9CYwAC8a1qrFOq/XiXWa1u77BL/c4/ukY32t8g8awbLKGwp5Szhq+IwtfOkYp
cDOj87BFoKr5nM6WlJIPPKMCOpl7vRcgl3g6AcLuwkzn07bYsIST04jGI4zxQ/3jAiuNx2P2tT0Q
kobKloOc1pwibL6XNaRR5gLG7DSenbWwLpPN0TOOf8KjYMSkfxVrGnHx4HiAkxyZY9inKiKwDOe+
R48oYu3N4/KDv1I1BENYM3GmojL+rbWp6cR1glMe9U09AbPC8zY2OVegokqggTEreNfECCvco+r2
F+agPjgiGR/sO1vIXud/uzYGrvWsrXfR+Krg1oMbH6Dz7yI77ctjxwbz296FCWxy5i2iFC5raTBQ
aKvHmHCQmTgbE2d9VpvzAeKnvJd91n6C8/RnOLwhVZauhsflGY5k+3UUJ4QpIPbua1fX6KZguTX5
Ef3ghYG+nBoVXz/rolgS/nfEWKu7ZZNLZlXg7sQoq0CQhhYR8MPQpX695NjPKtJnOf4/jg1oiZA2
wmzd9+JC6cOhAiD8TI6uBgoazKZFxKJwzHPn0z/uB2VkPv6mCQKyLg6pfCdk/buV51j+uuRdb5Ip
aCOiXfAthpndOhtDXEYGiQHJv5GNUCkfjEUpuLBvM1Qy1ZpN+jyHUm0LIiuF4YT7kN43SVt4ArTb
JPJm8AR4IP1WX6BwSxpvJdnfVM2orQiJv6rPjuSpa3kQI11Bhuj4e8heigTMyx38SBfVrfC5TGOo
mgwJ68MI8vHiAYBlwP5uBrJutq3ixEWo0bHhK+NPyuQsU8x2oHAddZ6BgrKTbOEAtMNyUj/uHe7N
pTEZqSAJk/DWyufNKb9XYWv/f3Q06fLETvh2No+7bG9NaUO+04DLDUXCZ7FGZIPeWYorKZ7rFx2l
70Xo8Y9R6yu46Bnskj9R8Ql2tsBc/rAFmlp+HuOsyhJR3HuHvLFCae81jXGqSY8tictOW/g8kag2
woZ3hZWNmECn9zx3Lt2JH3lmpMH57N4Q2a/i+tOLzBNooUy3MXF24Ie4u3JPBI0cDtuOM5bWAAxL
jVv8d5cVAdRY7FgAzl356VCFNdCWFIEDLsG64OUtSRuSiKz3zC51FazC0Rg3MgdQYm4w1pn8tyqa
jtG8XRvMJU49fBeW8EF8irUkitnvQtrECfNv8qBOR3hUPHWwWHh5pkgYf+JtHOCXUzhsqTK6ko4B
ybmOt1jWuboIPWxR8OPoo9s9Akpg7BImc6kEY1E1Q6IXfAuctyHchVhc4C7XJlklK+Dz+EhE1pvQ
IX8VhtDqL+muGTskgojol07bpU3xc3TA1eQr3/ZmXHV23eJWCCB7c1NmvTPi+RR92bTxw1BfSJ7V
gKS8eeTr7c9ceZSHQSArAJpiD1WW7qPgkWRNBuO9H67bO/tRPIzqI+jMD278MSWE5DaIDDp9PJ0V
RAevLK+FZoA89Fz76oUZlFGOifq+gDUWLdN777+/458bigniD5OX7u32Hn5TMCi6Ll9VzCVYzo6N
b5XRYVq6mWpky86Q/7WT6G6aEcFGBsCBh0mnExiO0jngFA0UmtRXIyTysk2XAoDb81FZoAIeQWq7
V42jaBsNOKrqFas28JwHsF5tp4bXTRpLGcWbpFvmYKar88BhwDpzbVjO4RCrzivHcTLXKheeZ3dK
5//KtcCHxadTBrtKhxY3oXGHZ3cZiAyLF1fBtBjuEHU/MC/yvdsFsMLYF329+cos37+Q8OXoHlba
lj9TYbIQEbprQNfWs7VrXdW1FkksA0qVr0SejwWRKLIu1TywiRKnScY9ifH/ZW4IZZZIjXtbrgNQ
c62vJyEURFiVnO15aXMq1lKb8kQ49usU03r0lDusbgFNngKcvjbmbI+77SkHYnmoF2j6aW7FiEHe
rp4FxensIr+ZM3Vf7keogEgbqsO3cdMMi+jJzcrWaZ5Ox/KzDVHP/pnKZFvBOFGlSD04KBRLC/mA
L+Hdhrfo0i5qU06MUECCfZ3Nc3J9NdoLz+XnZybjl+DVzAdbWcRGNhN+eBHVGFF7PjuPm8gkdY31
dhhrDha8RxK7qU/xDKvMsZY2FyCEibth6LVAFmzuCgZzlIN3Juen0uYrkBzHZJS0UQ+tcUW5wXKq
O7iBkA1+jVdnj05M/Jjm6U4Lk1e3GL4gLkMAQB3JGhZJHOVCUwjM2Cv8Paho8e84HaU7xWZ1KHJy
t0DTf6yukcW7yTtaZjcw5bHBHQ69UIOCjx4mvQCQvGCbLOasjM+X4Vp54iHh6eYItV4562wjvNvQ
tpe/z9lGFKWXZ5b8jpxSgGJKF6PgQBVpEMWSQFucOTkiwQWOfbVbpIZLgoS5CBevl8XJpe4aVYnn
kcn3gF/S7bAVCCyVOo/Lg0UhMjmVzksnXCeqJ43xAC1neRE8P8yhvTYyMDrAyS+017ci010BHTMi
aaOc67FhcvpfVclgL1eEcIA1k6Oa3y6o8ly8JFc/2+KbNp/LNXtWLEMwBRIVAtQ5loG8HbnEQ2VY
8oRCFByhMRukNX5x8pT7AMJsllTBdKS8LOX7T4ZO0BsWJlKryPxFsY+x5JqHIyxLevRvGy8hAIpl
GNVEo8z67TYpdFMXRdBnkHpt500MC/K/hiDtm+lSHyq78GvA5mNA1h1w3SavXHTnLn33lY6Byfta
o4TSV3lgpvRFEJUkOukMB4iHzdNC8bCsN4kgC+Jb0TccTn80iVsl63FNoVvNgxr/9M66zRJ+IWi+
KeSb0O2t4dP0dmMbf9i2bZgIVc+Zw5+yY9rEm3nJU5AQgpz0SGK/9MGg8jeDL8ZoobbBsIyY9qYS
+Iz/q1fU5jriGBxc7Nn7buMfi61DG3Lx8IvPRUUeUOQ4CNtjEbqdziCsJ+19fymQn3EK5n0erFf4
eZ0eRkN5U4TlL+qmfeMNhh2rNv5fpRsOy94BkK4di8RuSAWs0nK2Y6Aqd8IeABT+Ri5TBHl5LgDI
zfb3LYE0fAgl4FA/ZYeS/IRX2NJujC2ZC5MdQ7T4fD4ZoQ0kRpSbORMNgF+xRzTr7DhMA0T+k9zq
Vl+GGZpyGADN7kGO3yDwtIq1i6lOx8SvfDYpiWWWnA7uYSNJigp/JA8INXmip5ub041w50FtpxA2
Q3gfN/4oyBoAN/XVQs0nmXzMIm8dwx8fE/TJEzB12mbh3gOUT9Vb+S6QZhuYMeVKHrxT2hxm2HpT
WBP8dDU1wXteBqf6Ndu94DlyL3pxFQjGzNaopA30/mBBNPtgt8bMlWG83JnO1f49CfNvn0zb+EGa
jAd3aWZRzmHEiNPzLGuP2wbRX3vKWb52Wj6zbbaYxHMnCrmx3pvQruw5UIUL87vtRP0xuyikiXBV
kjK2HCUM0fKRROXusUAfQIKtoGBLyrfgy0SJUN5Ll7GSQIGQEX2bXRHV8128a9U7glhGQJyZWz5z
YdDQJTW05jGGP8RvBuyW0K5axLMPZUTMn35dLIp1LpWTr/82gUR08A759iFgAqqviGQKjkBDmnE/
SB9rtV8RzG7hVonbr4EtsPyOmXLNwvIXsIg0sMB9oQOdDW3BIMovhskoqcv1pQrWa/41ay3vuvji
AcyOj4B9d4hMRFxElFU2rrVoi82eluLM52p+lJhLDERF6tHiMNQH4FrB1yC7q4YSHgXTMquHENLO
t9T8zHhSPK6GWLMRnMdROxfi1pvA8oBST/0n96c2TUOemko4OSAGwrhlwgJXhbjbm9h9UWFIvr/s
mqvQjR+hOG4gHMEaQ8LeiOZDnhLMqPc59POyidN671Om6rrIIm/tKko8YBfUhtWDD2fztYiMXM48
SPDR6zEIYNqnb0d4h8elblEFHvP+eYAEN94BFIHMlcY1cUgx1Fp6nedIMhY/Eflxs+G+i447qEvD
Q28A3Krn+RgBgpvryZ61zfHUFU5uIHVx+dNvNjtpTf/q9cFwumomMGW8Fdpd6+W7QnXiBVimY0CS
YW3WqKTNzZ2ZmFXzehRHejHB375rXrk4UBje/nnrCwVYm/U9+AkESrBzfFExEZSZBSo4BpRCLI+4
TrNptMLAlAw/cheG3x36spXIRLPJVFbFpWFGCSrwcSGuCmrQ6vvVudeaTq9s3Es1FdwWljWT256G
QDTau/7m090PWHZDLdr6MaePXwbCA85fl4V0C72SV1MxvoVVnDPMxohu1TFEZBdxl5vGVe8/OCQx
tnB65s4mMqEwU31n3gIWuaMUqsw94TZeMHV/+IiTjccxL3TUtC2mhmHZeu7ng4rSbUbGIQOEBCoV
uEugjYbbmHsWoyZMakqHi3FJnFFIYtoo4qKEUWmQ/0oVkoW0cH0o29lvgw2BjN1uQhgZPgF32Vo3
5doHSBVQPT9BtggoC8nTEf/QCTDbgxZnq50ORzl5usw3QNS0A0a2kCmhZEn+icOXovdSa25G9V5/
e0qV2L1ZbXfOlKCGai4wprZyD+GBwtH1FdqMWE8Y+wDE2Sz9O2n86/iMzsEus9OYB1uHBdCpDnPF
yNJzZODT6JszN0Mp+TRHxzd+8w4rHGX05sNd5c3XC3AoZ9H65tPcYgMb6om8JzzguOfUtbof2FqK
8MfQEqck5sTSyjOdc9J5f08lmcsfSG0ovj4j0XJrHBu5cCaK4Yt0cGNWVAbn9IHfEv/C+B4/bdT9
zOJ8VgwXFFb+0NoFb/pwF7nS5gouNSXRPiCBiOx47jCOYmvpGJDdjCHa+M/6tB1W9jI7oHk7FIE2
k7h0PM9VaYSqH+YVDF3n/a7eXNTcd7WBoEfF9ulUj0o2hDUUWYbSaThiHDxajm6M3dVx8zGp2w74
n1to2nxGGuV02I0kbeIMAJvYMmZOrR+691HdJpT3aOXFN66uR7N1ZWJxKFGou0jkgyO9XfmknkWt
lseqo6sBE3vb9KDp/9p7VhXU3ZahqoqM3yxnSpOgoRtnm2+5vLAa1zutoNCHCtMUQ69vsSc+5M6J
PbyxkL0cmfFafJ2tWYJ0DOvw5MwMhR8eGTIQT15rfKXkZXn8DDv5TkEHa7DSx5BmXTRPeugnUbZv
wMfVg5JAiUsSHajRzQXt/VTvBdrU109x1L1iOf9YZN4oww/CfDL46A4oF1UfGsmqI6ATaSuBYyn2
Gkf8iV8cuOeyEf4DA0EdDM8zA/wDx/9R881o/pr8FU+F4hm0ctuVL9yYb9KPRglqwfEQkJD0z6QJ
JQQDiRCYQB4FCkj/5XSGSa2Cesel9wSrh0EsZqsDqZJGxgE6fs1N09QorbPqz1gegAsytiIuVsLx
Gm/KC3FrmVmAf4E+MYhx9vLzsZRuVlxjFhd4EnD8BQ/4B5OMbyvLPoFpQ/amZ57VcQbkLu/GcYT4
lZb8RAfNd+cof6peK52oh1cb1W+hoWFdQgPkFlhlLbxzkbvOMSQPlLVRzCOQiVzxWefDm2KSqXQw
mGl80VhiLtsOnn8WP7db6Ce0OMn744zDKgHYmOCBRh+dRJHFX97W9Pil7XStZT91CcdWgZTFexSU
nHS7VxLnpLlrmBMxBuEIuihuqg4Sr+Wni/An5ngIpSM6dXH5ac4MUFfawleMPDKjSY5nMzZZWNWc
riU/7mw7acBPZDm/gQIlbkyKfTc4wNoUpK+sNjrgdeAG2QYhdvEKrItixVf2z5eg2duEZiBAjzko
tA6xWQt/3iNk7xV147BNR2he6TRL+BhYU4WupOzaIA3ICXKzoBWdvybozMfcZCSlfTj9VgtrgrBY
CV+8IjvC8FCWdGOR7DNM2qXa7CWMtlwev+3bpTimRgAf9MqpAfjManPvELmwZEhY9cPdyEH45a62
QTXBDpjLCKKQn/EArxrdVGQNdK2cUSZ8/D1LIzBwvY2gnxoOPuAOAIkoQZGuQoe5Eo/CgvG7UuD+
VD6UAf9g9gUYtVl/10WWh5kjKfc9V4dxYlFXkapFYjA/nOPcX6t6fRDTkyjTIQ1qVyNaBlkNJOwv
pvR2Rb45YhPmePtJckR7hPZ7FX0idixaZLjAGJZW/rfi+H4x7wLul+CEK/iQkbSmPBxfNjf895Pm
74AyvcEiwf7TnufK1MIqjNlqeo+8ci3/dVKBOi0r9fTAp1OencviVZ7E7ZNZYp0sQ2w4sFMYsdC3
4P3N1QjNMxf8nnNDnQMTo5uuposIcVjvgMMp8Ac6XayEmur1MKP/RuSN1Nw2yEfFH/KrX4OB8t7Y
XsDrnKV5kt0pFdPViIMukZLTzBY9RwnRSG43hToBWAO5A2VKNL208w3Th1c4WWrpwYu3QMNpN+zq
dpdXUC6d9DNzo4Wo5GuZ6JqOsrmZUj8/nXf+5RP69D8ibpMzYeh8/4gIVvwwh2WJNn0u6UEEKOdv
57lqLmaLmolRkKsgaxfP7V+yll6D0tHhp+h5EZavCrXBnbFzrO9e+wev+qnElAbE3O2dXgVrrMQ5
b4Fj9Fyef3VMbxSZn0dlgK0QAEjsW+49YVbJ5ng9Tr/QncNuYDnYUxSg259rWCBlETfL9myJQ6p5
WmCMepSH7mad2ges72cvo7dMHDSi9A1AY5LEir9t7MzXQj+W2+WuqTn3mqx0E8z/l6waXE32Fs36
mzzOTtqRYp1TdokXpPjelM9PY1w8mXep0HWIOV7COtHgH012YdPYdNbRPCmIrNSZzdEpDG+lv8jA
lcbbbeytSwGB3yDD60ZKghxd4NoiUsp+lUEbt9esPh16Bq4XHEexabwtpgUDN7ZZxkE1knOCzFNF
uUFIgrTVJS04X2OEWN0YnTtXYu+HBKR8QAe0lZlJNhFniD80OpCbe52FRnJJEoCsB208a6lq4CJl
yKGpYu7xPoSm/9a2sAfEnX1YI2NSjY3XZQe9PUz5k9FnV+qq/zr8qZAt6I2cGJdBrzwZtXQsrW7G
6cqczMVIyoIPdAmBmAFzG5WHYdRorTSQAeqFtJTtfWczSO174M+SevuKIfH2XlZmYS0v5Xv1R6V6
/dP5eLP9cMRQEdyz2ZgNg8P2/4RmHCcpnnkEKb6fz34yxjH6PDuKkkXR4neivjCFro+QExsmjqW5
TbgvP5TsWWFr4v1oqJgpA47qCI3+Dx7Pzsdglc/tAfj2BgYa8BfoSMEsvAYijST4gLEOhoL6ezop
hYX9+oTEMd51fdfe6BT+705f8BAXAhYqUMuP/8biTvt6RUdjey9vxWymC94r2RMz03+b366XloWX
JnUpgjoZWEs1BsZwsRLyI8RtZMaBr6p2XaUlYdhL6HbMT5kfDI57L2uwagX9Ygx6iztkxCFrUvP2
CM59WqZS/3U3CuhMSQjb9ca9mMJmzlSAqz7lpdaw9b/Qg+vq8QLXOGE/nqO72VbPP3RSA4YDfG2a
H7d/D4JRHzYLAdW0e1RRmwNpXkNtY0Qf8yq4SEfBt70gzWaJ6WDMpON/ku9OLWlnOJOto24EEcFZ
5ZODLagRqIQjBCDZmZtuVF2k//JZ3vgvhXYYSRAcN/M2YRbU1vWuY0mztUtqIwuNYiLuM6eHWA+3
qZ6DrmSrKujkf4vIxV7PLsVWgPyFKyPzxiUFIlMIU5Ri3p7XTB9Ucu4+R/+hYVd0IBafM+SJEajf
w8MNMyxHYzftNDrv8LlChTER6r0E/PjcYrQsIRHQ56+RIdMKMUQ1xALIkqlW/JLRGabXfbSMz19F
x3r/vtv4H2REG+TAt9Kidz0I5map6bpAwSq+edKD4UoFDbDpncim69ZHh+3C0ZmilzoVwXEuCLY5
bM3u+WqZ+Xzaa46i/qMUPuhB7CKO0J+LsH64sL4C+E4xGSEKkQmjAw5D+DUZZ6T5w19Jj/pSxQBB
zC1VLDzYJ5uQCP9UiTPOoEspRrNPsHffiS7qEiFXDNpLVXUsU2tqBOCRmv3kvw6WwasGwBLSXM+F
+f9HRLIsEVY/spqxF27BpWGwRz8iTZ6/4ZbroPGPrIci7kuGIcNAU5WflYZumbjIiaB9Hr5w9Yiu
SBCoASigDHQOrBGEIIxtFpQSuKgPkSfDplqwOeDsi4v3zPsUfc2dopJ3/mFtkHY2i1IOG3VqxdRH
8bojDd2I8EXUiYcBU5rnhjjE27VmBrMXoaNi7MniQ84Fy6qQO5DXVLHrNYYr4IVYkxkPsrZZ5X5d
YEuKw0tfczvr3uwzxogP04ltwLOMUE8xVlhLtVE8+oaPl4DkSOTppllcYgL0TQD+XjyoN8BfV0ay
0zi8SU8V0n9pqo2c0eWWrXSlLMJ3zVDoAcUCyrNIoGaFizbtW6Et2TSz4vGdErqhUlkopBzAVbcP
5YLH5nTBfvseF/27vMRoMhdr0L72mgQVTWKv3MJgQw8jcKiM8p8OpuZaY3edV0XSYp9Wq/gUazkz
qyQpUXBu3Nir1p18qJzNRz6ZRITSCATBtclDncM+JQ8Gpw7kPbAzTS53h1H0TZqFWCw5pjYOMlJV
cp3tV0pLP7vyUMJ+AyMqnlZf76OB1FgZmeGy5xcWeORYowiVQ5wRhfq0r1FPu6KQnSYrxmU0D1RO
qsxcfEoBwEZxwTp5eR7ElH7E+wFJOUjTZvJcHzsF3qbSYAOVvFLXtWyyFv/YdGJzuCNU0R+U+JW+
p5MFuzmp8Xwi8OdgeepU/kmJuhF9HQrvTzzeAQog53vkjV1pFBRYoaZ836yF2bPBLqb1SW38fFK0
9KRIAONgy76e7HgATWBxAIB5c+Gh+KcZUnnnPN14jUaYtJ6AInPIrJ4hZ/YUU/UbtD390u7zZja3
TgiiC8IICwAU1AutDuXkudrNNm9topVOjGDuzyfy/jECHSIM1g0ubFxC56trj9n9X93xMrdtmQf9
yhfxLmQ6Pw/JdsCAR4OFfgSocjM7Z5ZpXgO3fQ/cfVT2lumizUN3PVT6mVqxwxR6c6lVtGdfKLWc
EWMNXRXD3M1lDwwS/dcD5qFjQ/5QhvOr1JxMtbcPxSpGn0qkeucBVGnj57Mv/XidZOl+UfB14NX4
TUiyi4y2I9YwdTpmMFSPS3ZlGr2ojlC5uT7Ruk4UFJoDR4qNac7WIKhBtL7b1TN2O3CjumwnLC2y
0fWyqshdAagkUeRhmstNQwGH6TLnL/cyqOVwt+uL2AgTA3DwHwig4L7rKZa+Y5Jny5ZY4Et0Uozs
ebrtOHWILK2pm61zWYoqBfcMnSogdF886p2bMd7vTPdFQOypqrb/cU51Q22lZXJEoP+9+LgEPYyf
5EFOpIbF5L9wFwN7cTvXcj/O8OT73FXXprG0etaG49Vy5+qz1ea3mPJg8neXlSngkfufj0EER/Oj
eSeMWXSVmBfhqX1nc7MF8uU1W8YDwW14W/zfxAxFyUkngqaoseuuljyuoOY0YEnbrOEBdZPwGBzv
p+ZPmIWkArpdrfFGdIeTxHWF42oorYhx4Zk9i1FTRUT3W3TaLlac6JsWoyEFjXFhyOaPPpTuqVY1
4+UAwqUIq6NYF93kPPPTPNRyqtC4whT9i07TsKdVNWxhy7M/AELzCvcktWYSpFekS9cRQ1N4TgSe
Dy2Uuxf1auvn+mWy2CH8GisWheVeZre9gurCEUqkuH6EKQqqtpOsJ6N14UMUvzRP2Iwc6ckGXSla
z8gMceAIa+u4Qk60ZdJhPElb0z/8gvdeRxsNas5NSi3LowQK+nkTn4zseFmUIoiedoQL2EfHObId
99466aL3L2EgNWnbiTh2KVhnPxh64YqeojT0S1lfbdh/3CdmLpaxvaHTXzdZvoUurXgYa2/d3cdC
7rvkT2t3jg5FQFy/GEqMBy+sGjGUwQEvymT5WArAhNQBhosjKxWpXJ6E83BXfF8BRuYbRS9RM3zQ
e28d26/XRtMNuUVCA7rKNzvvxi7cnnOttFR4xjkS/AcrVOIaprXLHCNETiF0BePSqf3dEFCi/XJI
esF463hHkib2vnlGa1lUfwQrjFnpauQj2Dx1IEBEa3g3unB3tO5X3a4V0pZCxG1iuNUmm2z/QeKK
8IpJ/kcdBoBrBEaDdMJe2/bozk6nqbK63M7EHq3TNd4ZevoDfrl7vqsKsK8r1dfXSzQb2PibBcM+
AfHI1c5jhz0Lov8QMCwGcwLGI8F4jAtV6dPbEtem/o8hirms6Qu3J3GbDxMQDDEqQzS5SstL1FC9
FW0qFBLbC6/AYt71Ao+E8CpzX4umvJfqt1OqhM2Lrs6A1ftw8OkG/EbnxtvLirrWD01qqNmskjHR
jyRH+nuZD84XbkD5bfmQBGSxkk1eZ8OFr+qBwqcBu4RbDxS/E3tbsUrG/y9f/c0oD9SRTAfiCZj/
7BfwyVnAgclO/7aVCbegrzmGuqKoj+B1nAbP+OW2fuFu7TGgQ533OBRmNOiuYtKijL3JqDLscvXD
nIQrakz4jR+RYWjBSyIfFGPX8C3G4/FvFse9n/0ExUInZbdEcy+PUmviiLFoGD9T9ie6fi2ZWmse
+nb8vRxU+AmzhCqQ8RtWyiXc1CtBVi4c5+vZu2LJ+iMtxJxNuqmGGwvG+wAlKkx4SG0/uedJ+/EC
SdxETCSN0regnEAD2DHjHowddVEySd7ctDTXIe56cl1JXROYsm8hB2lT3ZFvAABnzJJTuZepdKCd
o0ha/SIkXrBKaVAEw6RdQSmaEmowkveUn3MFObEpV8FSs+Z0XdVh7mVPCWDUpgOmItvJ48vr/UPm
moLpXLVLuZ0dXln3lrVNkv897uP94i5zxjrt/prltpOd36UKMeUXbNv567NNPw2sYbYOnuXVH6VU
QhmVn0xfFEECbU+tGQoZs1pgQbWb+9qTVONG6SGF9MxXIZdZh1eE7QnQ3MYGSg1i7syG+6h7NrQ9
wlXlk23Rbr7Kd0pATfSHfFT+NfcwCU5iEOBAv9BnqEclUu7MWNtqMUJvJCuJ8ii+DCpolIYmKdcO
Bz2U8Jb5fnGVFgg4lKByZPGjr5d7R008C+MhBzjpGsDZGfmlkVjBwpMi8POv0RpE3MhesX2DlUG3
vJLQudPWGfQE8/c33W90VbBcZE1mjZ5WBoRCUL4hOBThedsUTQ6amIF4qOA/eHASAJXT1N0rheVu
/YoIgV1xnVg/0WlJgu7ubFGXQy58256+edpAe4wOKUkTvkum/gd/mmLXAXBRKW8cdbETfi+JIJIb
gDfY8OoAnSqPSICuvY9oSNQ+j9gkKYRGEYbFPExXs/3Vj5JeQMqz+cDgYWDNju2Odhw3tV+US7oG
VyTBlfeW4uW2YC14/gy/P/+vmsQKUN2XZisFKDCyccefxlJpcFvSUwoJ8v8rfqkKPzxB7Zdy5r+9
pfEU23py9FNs+eD8SKqb9mh1+bn45B1BkIIUCfk3+f2cBkvdmWmfBxrTmw8+VZ5hevPuyuakizx4
qZWOOCVOKVyfwIHgekDevWV629IFR6lBfwXQ/zCwdw2Zt0gVrNfko5jv3ssCgpe4LfadI1UiezwB
PVLqlMDytmvwx5IRTWrPBypShbQ8nRbliyP102lSyH5Cg7numdbIbS21lsuaEPWAc2k7+dovRtYg
UK6EHHpMeLfTuS9ZFzMjG5pu6uYe/uS+Zo5gLo8RGnDXNMQxydnhHeczvRTOzHNBZWiAirari0+D
lcfc5TzfjbDYa5F4nG6RBE9kCPVgA3Wcbbpy7JUDK+t5oRZlfekpp4G/RzUg4QTAo+qZxUoNym6f
+PSV63CdubkfEjB/H6Rv9ZYJ8nJ9vQjqcRzXz5vhqRGu6zRZj7sPccefE2QV19SjJ9Hc0/2+1H/c
9Ojr8LbVVWHe7c8gzCmDBhk7YEPCFoDiS5CrblOxX6yElOhOc+V4XYa1ZFq1mWHfvfN/qN6TklvG
2LrW+6cfsxpXSFI6M94Jtwe4wsaUEbK6d4pSfieaWvCBdkKFslCt2TgmP0oUuyeADOu5oyvdtmwd
0sGM/i2BcuzKajVTs9SxMBIkpfUTG49Q8J/4ZlB+kB2hwst5dxY891Ck5dfoYbbu38yt8FBwmIJr
u4TGUgU6ZscTYbalCbwnn288iezuWOJCMceeZ29rkbalKXtLPrnpIDsARw2fzyyNJgAU0wePoo+U
+G1s8zW1j6skcu8ouiquczEasDQqoMV7JZQ/tAfbPyKqIt0oFUilaWMtjHCaGT1wM3qTBWaN3+qS
H/C2BfGEUjUVaUgRLjAjIHSLDyUe0AEwlkHNFask90Y8Z0iiTEECY+CGEjoV4CmsTGO/iwflxL/7
YGAEHBm4+zFKFwAzR1OPsO578aF3qBb4zl0LwAvpjXzGOD3xP2zgCUdEBaFBz65ZJdI37H3uGQp5
FXkohTjDIVSxDEGKa4pRv3DYdhh0BEQ+DT5wWtDdK+IGF8QEGm6Vy0v4y+nse8Dts/a/M83BV/3f
eYGx067jmjU1B0Kt67E0Hqtxn6sOcPnpDeuI9XS5Vc4dhEpENL/ephUJQzpxU/oHlCgmEhrkWWb7
RPr568pBOmw5IpdOVCfYpb44BKRZ6A1tc1OKCpbIXfhSZ5gLYJvRLdeWxiFX9QoR9/woCHrme3qg
3Lf/3WZoqsFeOZrwD/usWGoUqSrFrv21Qh85ysTJqFuivJPilziA88dhcz4LfgJb0kPepqjI7YFA
ZDj9JX+vSGrm4F3vLGrInshjU9cL2EpyQ5/GnU3NlB/K/RYWIE+BiiZ+gmlkGy/DoXKwvbhWiBfK
+k02DEEbxMl4UkpzsRESngwMS0TMi2j3Gu4dL+76v/qHrNU5AaLo1fEBKt75aywx4il911i8CyWO
a3OXIfM6iLW12c2M8SbgLqBdPz2KCVakOQC9saXyFXq5dfhC0LAloEk/dX+48tN3Mf783L36xoM6
7J9UCyZWVcnVsTYPdVOIM4VjhdZGqv1/wo08juIZToA+UDYdcaiaxIbC3tQnEt1hzLBl8y12F4k+
zVA0MqN7kpWMmKHAkYH8s3pVpidzeStGY4t3LKm5nbBosvwuCWz1Phfk6ZPE1mYe4b9rSaX67yXI
Lg5o7Ta1Vsufy3ax8NFMJuCcBUn1Aca7KbMFbck9rzDd4na3X4B/MbJl8AVDpAIMa1qHUY0OdjBz
IoiY79g2t/vsNgia/4KTYDYqObpr0DqI1GSgAc46aodT1KwplTE378FVCswuoXjkRf+OBnWHRMDm
q4yM4bhObsZZrTsFIZ3sxdLVM6kUocVp5AF9GY7rNlDz19Fq18OdeyB+ZnZJyoI3oicdiAJ0FDx3
/dd3CTNnu4iYo3DzuQD7sa5/NnHiy1/VYneLqz/+SYOqHG5TCtYCQe0h+coE+ir05MQKQlq+ibGB
Kj87dWFyXTa6AExm28Q+1lq9U3gsTHAFD9GdHHrjBVSm7nphvBk+9X19Q7WCyOArRIXuAc1I/e0I
hAsZln336qkMynHsHhnRMNAdMUfE7XQH9MR7C2Uaz+3j8VGR0kqJP+7O2WlloWk635Od8Ow4dni9
G7KOuHnZoWAfAfum/MsrhWwsr/kB9fwx90Qjglt5om6jgOYwBADD/5UF4HWAjDoeHc2s8h21OiSV
BS3ZRsg5lGXbdw/1x+9qaREVqrhwQf6yIKBd2xegGtokbvHeYyB5JdKHUaNIxNq7LXWS1TYwEumj
Z2sAMEWzhN5NomRZ4RT5jymevGMrc+Hw+fVhCbZQyN+LkZrjTlyOEo7JXfPnzmhlWzpC3YvCB8OX
e4i10MCUEk+FN865iX60KgyD5SJHYMfGSz+b6jeNAw+w2Eo5uKmHlSD3zMMGYFrIhmXo46YjYft7
PbI8PUfjMvBw7t1RlWgjxBd4peRum/mXPgEDzoYleTd1UmStx067xUP3kpn0NkAz2zw/gVn6Txnd
gz3oH0KUVQaxCozRMsDg5IX+fbbZs4u04dFKrqLLc/LUGPUuAlMkpT6xpsVJ3C2H4KhL6fUda/eT
mfhBzqwdIfn5A8w18wIrFbADrakO9p2GVJk4a3p/jQHxJ3dqylDkOt3+K9gbWNC17LFQL4U0GK+7
Wtkp2IeCJWgsph5NgwzNoT1abAWEB4Ej8gKkz3VowYF6pp2SWxckQPiwYHh39pnMLblRGWera5XU
itV2aUd8Bf90LIib7F9nVHPpnRJ5b8LIGyCkZwF7+h04yvDC1xQv9hSprBx4IdSkzuaU3iBDndMl
kvNqmlwoeSknMsSxH9G0Zajs//kON7kdho5P4bd+m9LEMLsyj1lYvKhQO5qMY9OBgd7IpeQkG3rt
syqSQBeMpfQJqdXsXL+lQReJZR4vrq2gkF5+WIR1ZFlFLNd8cJE6H5zhl+146GB7a4f/7mwl0k2V
O7swneDXqPKv5Mtd5XE+4mVUygXmvt/MVu6hYg3/K8uyP2Tdt7SkLTj4M5LKoiltDJv3Pfe77uYq
l1nwBoTMEvu06MoAR6wzCuETzEUhBZaJ95uJg8sX79oRK1LZAIthK52hHKemPebkWbqVNjl1uK9k
TauW8WYXI3Aq7YVH3HBYbKatoTPxts2WkOlbWniLZd4G2klF1uCC0HGM1OKHmLK9Lsoh4A/PD6i+
9BGG3EQ2bL7wEJpd8BkUVv1cQ0NzYn7BT0P5jlr8l6PqbpIBcTA/1/L2v8NsAEWYryn/+6GU/JnY
ZpzZRhnKwEZVy/HBbfQs+3SXcrWQ5V67FhddzMD3fq7Rz921bRFXN8grL+a1raW1ylMy9hns2UNN
ywGewlcE2OWp6jZhuD23JqBsxF4d6j1215+Qsd9ljQXoZ9KH3oKMLQxWY82iAa7JqOHDKyLBUKXq
uosj//hNo3V78DuyrEpY2tfyOEr2Wy0W3+3Y+f/p0HCkR4yZ3BhMADQ+4v9onvQqKPlKVhggYsXJ
Rr6X4h3QcE9TgibsARy/cUu/Q5ByzTtq8v1TrmtjCWBbD4fOFJXDDDNn8H9DgX4a8Ya0G4N/pBy5
x+6RCgYsX1MbQXdLnlxUMBBuSGoN0Ik6s76YDKGZSUREPkZ34K/Ezd+N4UJkN1uXpzIc6KJiIC4a
ElUucG/+t4fx5k9ZaMTgpsNq1dLBFfhRkMTNsTLDdL1/JtI34Ia+MWP40resDSsNEC8Cssj0i39Q
mg1nCEj9bEwqTLyDDrkKBHPliuh82YkalGd3tAGNH06HCDtkPkw8pN/VDWys4y5WyHoPxqOJ5WiU
2b8a5gMLR72DZj2QXpOPXzF8dqyQCy5b7cjh6yew7x1ynw7OTf3JUy/Hi06oD84DXzUT0tV/GPrp
uqyzn+eHr8YqVSWfkEb9EDoAjD+3suuN1AIV3IkSsEHWEm9xuOY3fN0Kcdx99mZIlbF9Egu9nbBR
VVXKkCuLG0jmPbzBf945CCtTXcVPHa3NJAFp610UXZaBz/nvDp9w7N+6hqGSeoDDxxJESL94FREk
QuXzn755uNcG6lrala7Rqtt/RoRpS9EdNL7QManM0+lluNx4TRUBw7H+0aiFFBi6kaBOoBgoJzgx
Dz3oc16iCkAGWxuz8VkIP0FornqCNlhzCchTA0NkCIt4BcNa4vV7wnqJLWRjHx3LJyWMBwjkIh4E
yuWDuwBxqlH8ioBT2AVtd0DWnmP8CSPg+2RSg+MQqPBqEwI/VVcSIEI6vAEnQ7hVFw90Jw7qQyux
gFicqZQXXrRPaN1qEhCCJtHxFP0KjEj/NEsnlxri57zDa+kSLnYWRam9niM+oqVZJCoROV/P09HB
B+0vrVfH9vF6yb7xqmZ0VR23IOzjXYyRbXBCE6skjTSKSHzGJ1EXI1cNHL2JpNo+r9jyQx6XcpIP
TV26b1d+LTaohpn3abcJuIFG23EZm7hoZprlxEIZsDIfBM9qUa4gsjRs0RTK22muPUlT7oTtL4Nw
px52NtUq3mPRmfzeDZgGknI7TD/3vV/3FNqI/CyCuva21dAQwGKjgXeL46eEBsRXMmnlc1h4sPan
GwisxWJr7sEYZvmXdgvO/UlGe2AXDX0LTZmZyiCwxVbku80Uf++8zLRNsTQtiew29gEqnKZIQ3wG
FOyBxhvHQPyXKpPlDUUh5FSxE44C7Yq9GXcDGqQDCzBZpbz9QuJ84poD4TTHM9r3sW6JNUAIqE97
m/fV7wLVyW1OeyeSfJzwsjY4OYzepuA7vUkvVnSnHpvvKJgvCmbY4g4h4MwoPdby/ftCt3JeHFuH
GYCDHtSb8Pgh0M04cg6ovSLq0FMbG/KcGb8/Xs3vTQby9ChDN+NPhq9s/ex3PB2k+UoxAnQ3jU/0
Vlu+IIAUf7JCFhiy5U999914J3nQlSTMzdiz2D4mu+j8RmBuxjMMl1kHqY69QLyzM/F/0cbpQZmr
g6XJEmQRC6JzMQ58RSF+RNhXH5aX5aoTtOQUwEIS44LGv1F1PUYeAD+v2/wKYpd0gF88w611cEC+
JEA+AV/HgeqOGE24ijQosjgZSOQU1XO3E0njzTSaA23NW6T0kgj8A5RRFdtU/St0qd/KY+4gI3dQ
2ubmGw3MiHxcmZK7QckwPnZF+QQ9G5g3vAQlLO/l5PAF6qYqJB+37dnKQr/nnYqDHTHLInDIdjcz
p2DdvDk2TqK/gq+0nd7EhoCtNxH4HpHV9nW8HSfj4Bf7tXDPa6KAIkLGDLnhS8/nRu8jSTSIa0Z1
6/+AtwlllXXty6Dz7OGB1JilpV7kT1KmDh85VKUlKQAZVtgi4LegnUDurLHlAHjTIaEBbPGpAsqA
VUxVuzssY9oIw5ADqLgb9/Iv1GrV4VtE0WpHiNpD1DT9P19arLHqBYUSP+DMvoSRxab5ZQugHCbr
R3tkxjMIU8ZZXJCjFsMgs0esUiN3LKL/Xd8AG5HHNd2muSxvKuJykRrhztRwqHp4XDQyvCI5WSbX
cXhXfo+D0V5oqgmXY1lt42uXkOjh+UgiP7aLXXfu4q8Ex81jKeX0md6ID03mZ8YLoLY3suFA9Vmg
2D/lFZmEkT6i1tPLWJNBgq7wIZ1sZpbz6GCjZwbu3H29Z+hvoXOSJ6yydugnxw2teUlmg9GAv4LK
L7mP9V/YgxGPTZf3WnUJxtOgXjWENdT7gKIzxQZuTTVyE1L1OBGzFrA+gBsW2DL0MOJ5/BfT9hZX
VXiEEOg5eHrs0TMBs7mVu0LHjqgfbz5Cw82OMkPfeSHC9mU9X1v8cWjzxoWanRBVXc9l6VmPvIVl
FfiWNNbm+VrIsbb0TqWJZMYR1uA2QzR4RVcRJuNK2U4B8nSCxBbl4Hb9+xr9emN5ghc2eRPHIgbb
C4ONdSAbuz4jZ/wur0FOtyw0T0snALOeh/eT0B4jscrzzAM9XHXOCyQ6SRMSNsG/Q+X2txaTEMqA
87rzCLrLUMjzMkq41VxI+xLZVr23YJsHDl2JZ/g5t/iUgZXEAOuobWClUNxZvPdsQfSW1xaH/fsw
k7sAvw688mX9fLdmowNKbXSdG8d56SfzMdDMzITRONhq8NpYvu7P1IB6y186xUi17TcPbl0Kw+hS
UC/+967y1lwglaXkb4IPgqvk0hjeZAZHLFjQgbDDSUm7w+HwfogDEovtpD0K/uHeKDER0/Pa/jf1
NMzoVGsyGKdlCgS9Fslp0X/5Bv4yncdjWPXm8Ynh3/gdy0KE3pa0urxpsgKTR5r9OEp6QrMYwe3T
96UjbIRA1IEf7epE01ani9YCb6rAgu0zfKRu2kUZ592CufKDJppl7nv40j2Oy1OsvR8ac9d+72Wj
hKb8W0eEktxBk2X3S6bRVF2JHZ0J7Aqw83K5M3KhUmcW7u1XQDZc/YvX5oiVrycoly7mGBY1fsUy
DSbiUKkp4npC7MGZnnYHmudgiEPfJkkg7EacsSNC8JWH/cJH704KYzFq3dYADInEu3W+UeLGBV/0
Uf8Za+lsh40uYfYyWio9t0kc+9GRt0ZObVz+xcRhyz1IcCce3QT+lTSYg/hj8CJVURyTUykVYI6a
O9hRVt2nz4QGTBjEUC33axsb9pr1FmRxg/kgHNlPqoX0w2/4rLvaTSKraRAQ93JLSFGAUtC+yIYT
FjHdetCFtf/sxgii2LTMB3d9vmT+0ioI1sVQYwNvYXwjtZ17s3+yITAKQ2srRgGaMZJmyW9BVcce
tINZDtMVjgqqKUTVMFLc8CFZKG36q84bdRX1rZdM4EtYRqnfqvNVOSEM2OjF0f8ZZWzwLq3trENB
Xn83j7GQRZHU8mGQcH3G3ASQiP8NfsihEd6sX96wnUP7Llt0spFWkEwPjXHU7KM4xBV3Ge2lu/3F
L1aCUBWPx2k7+vIzAB3kgKnNKbMBxWPJJYNzWyiVKIAxZbrateESlqOpJX+u/jVVfyAjH5e4rKfb
Kc2kr3ar38007+BQHtEM0g1iQzUmkEm5A2p7PvsRM1i3agqPIpKmtbwjt0w6yu8uiYL/FDuHH9y8
5FyW/xkQS2Y6jpWwOga+H7nq6s0WzoL+MFDj0fBPna8uSndPzFZbMQfxK04Lb+dIXrvMPptTbepI
egvF0G2IzQwm4gVeJyx60giuIqeEkbhRkyYUpPeSp5+iAUvwNcUTp0VdCdy9YjmPRqK/mDHgbUFZ
icJq6d7pIcFc/V4jgh6u6uOuHCwNJljUwFI2DkcJCT/iitBQEljKidDtqxQWfKrmeHqjeqqiYIyq
r0x6SsN65nxcBK5qZLyVQxh+J20htnII+xil2xvd4YHS7HIhgdtB2aHTcgrMRYJtPKc8TBeOCpkX
ggzmcs6f5O1oaITLv74dFi8aogq16l0CUy+96CytkBQ4u1Mm3E5Mk+j09AjsWkcUBIBohcPR1bBm
wP7dAeEUHNMp8Il1iPScqMFZ/zyyuCHacDRvrKEcCeFmZGPLSkTMMCzB9fCCCy8RGQyscxo1VcgR
WZVSvJg2cP1+LL68Av8H+LE/aXbO+2wvWJaAPk77Jy+1Z6QRQ74UZLduqerJAk6ntHPYW4sFR2sK
nLzZRyz6KCNIyj/CuXg33KQFwldUKz0xyJptJZx6qkBnFwYxLWeOBDaJJOIv+j+dkcQLqKyWEma0
/15TmLl/32UkWLGdVmAcErW0FlUb7kUGcc4+445IvCz64bc/4Xoi/ywuY26Lhpd/d2UB2Z/jwT9T
eKVqW2ZkibwUrWEHOnkJobA1xjR1I9wDji/9k3Zhqiw2V/phIk9BfXfZcc0jIxysZaoL7R5FOViJ
1pFrAuF6Sx+cd7NU4do4xpVdO7QDzwJkDjgFaTx5OzNTQa1G5AEakvSybcP0m8V9OYrE9Q14h6Cw
2f8MlOJ9CG7IoQGp+pmH0w7j59+cTmjWz19u7ug5t6ySaa6Jwn6+P+yF7Dyio9T8tKBJmUZcHLrd
xHck4iOyiTuUHiqEFE7DGGb6UECR9NdEwXpDYcW2a8KY6S27HvwSADCmebt1Gz8XRB8njRsuI33s
g+ZNMWTaxRI8szOFwoJd9nxrULjtuArvBP0Q67aj5H+WOirsWb2HwXdzZBgkxaiBDXV4BfCAgs93
3wAlu7ONIousJMFRQOpW1b/DPLUR8r88C/gEoRmfGTPNyeZg3c8JuZKqVCtLz1Y9u+3L74Cr2jpl
OlC1VGvC5GAY/U75HMV1DCIaXXjCwujpoyJgf8HP88Qh8KHkqHkxjDQZv7tUySlCkRMFhAjr5nz6
fZzV019yZSIbrhXvygt7aLLyompF428/jbF7fzb+XRPSNkGTnIA3YDYK1tiN4m+GW1N/8GXZ2s5a
A52fCq8fRzS0irXBHiEC0904JM3KnLT8Dn4MOXNcSWqoVsKTJwWQGPsECaWO8odmOkcxb7tIGAqy
QRcbmsRBC0TDXSCVYOPHVIznwUXQmnhOA6c6zoz5JtnM6cH4FqRajtJKTiYBkybOa1cd+DAN3rGK
LGW3ToUmSc5q+UuAzp9j1eS0vhf4jIksXJAOd/PjeLRSFIm61hW+k467W39B6r1M6t74nuOrXDtT
Q/ts01o7twaNWNbbEpNEHedttAe6nSOR+sT+I7CUDYy9gBFap7BdlXeTDDoiwbwq+QicppkOFpA+
DzApXv8M+7W/bsHm3wsndcOMsAV/20CrGnVLE4jqkeIjiaCKhS4c0RndSzOVaQQI7yZfrVTZyDRV
GHl4meQpiOYCHvTeuCHa6hb9OAdJFr5fEXMkUabwJn8qp573j6Kt9dB/KbtjEAi2nZnQsimknczL
ephjzmJTS6e+HF8CSATol4D1T1oJjz7znASEmu2lSAPQeU7YDhVlXdAkCZazuoTdWdVoILOnsmn5
1JjnmLbMpR9TY04iiRbmLwDELoH7zjHAaIuYJDxqRnWduI18T3s8R7EeYYMkXFyP7cbOkX1e4X8u
xeqqGw5AuJQYDhuU7Ej/+NqasZ3Knt/3Xqb3UrEhl10SGyZET2Ac8UFZ+YZ/W7XeyWkqyVZxacCC
YxfxiO2d+9nU4qROFM+5iXztFxNxvpAVY2FhOxWIIhQMbbusm14Vc04f75da3OqmF5LWgaBS0V0u
l2Nm0JLkGZbLlI8XBEapCJczwyC6yhKy+Eu4EqteCPgi4k/xG8RhOzvIC0LqilU26ph5/HW6WibB
nOafnsQnm6zQhIkEEQRcm41VzwCYNkHQrw4G5ixTIQEZ1hyk+zz9RmJyToRjQSbNJi9OWDNeNN5E
uGAZqj4P0gZxyKonRY9OcdADNB4+o7Lx1q3c0AiYN0SoSGX4UiX52s4bXmMcceT7oKiGyB5+CNAO
rD+gFmwkJjimY+xgMILz2tMx+3NkS3VnGSShOQP7FrSqf5IWzuIl6gWVmPWsUsISK96u6r5I2+dn
v4w6wXDBPuDWGlyJPw8tT8ctGbLOUXBTdgIC9CK1p8iPbi3eYwEFJsWCSGcRaaGgTs0Wtp8jo5A6
UgjolbwJh9IAcyiJAxjBOgnI6/4L2PoTIzrWP11QSl6+3wG7V8E9ioHzgAbfxhY8sI1dLPnJJuPf
b3fmp43CrbB9YM9ZiE+V6FP+2LzVikzn7rG/fVi3/EWSqN4RHpSN+VEJM7El9pjYUATNstqiy6Oq
qTTQdpr/FB3cX+zV3f2vYS2JnmOs+wpk9PTkXfHFbPUn5nLbqVC0fChYw02VyXQjwRmP0XAmkVCn
tn+T/BEeAPrsGQa6u2sW/8/Pi02LeEUcUaFm6MEMQ8P3OZuXJHHiBmg5H7aPj2vMV5FUegPzvOjv
Zkm8bZmwPcNpy3yZLof/IYxGnCcfhht2eTfnxFFxdEMbLEg9iNqRwhts8yCtX5NnIIesFMOWyIxH
YrJPLeWqyiiE75qCgdqSjCtnL/OEi6uuXPn4QdhDnctYMbbVRLqb5+KiDz2wJytHezFfk45QM8nC
/O1jG9z/FactcjEmgpXJwUvvD0wNscCDVYxWMothcqdZTFHVd78DMaLlvpaGzmhi2Sfr1imjlxK+
C0qUXE2EXURK0+tWTHpKoak+RBUkcDF9MGyOzC1Ie9n7snFdHer/yEDo0nZRvqyebXPyGM/T3Qbl
9tHk9yBiuNIPs8frcrPdSpqNGAlNuGAKkVU3lc0b/poo3u1GWULqyHKEIhp4mbNjHXQb7tCi852k
PSR9iHcWtiBLPY7EkRPNht9dMw239nVbLWW5iDIkp9dUEmc7l5f6F2kiFiX826QCRblNUmCaJNGE
HfXtbs/AbJ0K29whFqz7COpCGv7dkUFT6yKtfgKFvfH0yfycmDj80TXPif7Bq30McMKnUawdiljU
iNIRBmgWASXAdSrryqMGI34ZZ9OH+xTJCHQKIUKdM0gzH0TbuSmGraBqDgrrbN4nrnrGsBegtZFv
VNymtzZlrWwR+bg2R/UD5gAv+k9iTcsmYlZK7uyiEeoAwB82NKIs873jnvqzifoZr9xj4jkEdwTb
RPfRcF3BeSfb8Wp7oLB4vtKKXvmUZgqGacnQRimetHIjnRbRWOaNw/PvtjuKtvBpySl5d9XOIrcZ
LRZNtjau3fieHX0uDp9UZmUjdpdK9YBu2wZdXK2cg+yOLQqSl64EKGqJ009y/kZOsOtSkPS3jGCm
2WUQLSDMny+QTs3zy09mov11IYl8N9eNHPpW/DU7YdseF9GxfbQj1p0iskW3sYY0/UQm9dVNywgu
cl7jAAYuUsTMVTXQderA9I5sUXzVVckPvIG+nFYwkFsDNpMyJ79j197zpXbRTtV/Wr88dWkWkNB9
ko2cRDmDURHs/hI/RN/63FF8WYvrL9Ud4MrBVL5lfA0sV1FOlI6tjPMiXPutClpfmORbiwWB/PWG
lYJt+IVq9A97x5BdesffOHqFKdWEPKtCdBVb0Kid91WGJVOMdFshm0+PcAFkxebLELRmcFc72gDn
qxaXhqJdBOSH3Nr1hky48frJlcpkd5q5hpWWW/TKME3sjlSuAHkhdFM0H4b7b04unQuJXAkBa94K
b2VmkHNWh1XqyuMjPzka2eZlrEEVnnKnt1kpIOH4GQNpalyj50LyFkeIgPAfCTEkVLvRPO/pvZPd
1/Om2iqishGjngPrrQqsBOoAl/Lj5yJ9uX83/Q3Z5iBTAv4JXmw3Pi/O/AecN+JtncwHL5D/1igj
zcEtojqR25cYvIfBV4o0h+cTtnFmzWUIaeOMtW37GnO5f/YSe0UvkJ6x6jEI4+x1PzdSGxkx5N8Y
mzep4OvmAbdWXUfmnI9NyxEbaGPzWHdBX/SzmgairyB69o1HPGZ8x4KtrEK9VLBxn/awEw9HzwY1
SRSO/jN0IPzipUaAh3R1PhY36sR0LkxP1qexxvTPnym2ePjBjatV6orOQ24GiLO0AFRYo/VlmbwP
RtfyHE64+E9qrsxWfdzvf51+t5bUwEOtXVZ9Bz3YUHwt6W46C2H/oRz2TfubMdFmzi4pLwQ4nWbe
6qr7CbmwyYi5Zg1vz45ye28Fr6jm4E7R1w09LUzah5MC5WzwsBpS6UrMpUVJZL11fsdasMtIe9Vg
gGotmHdh6OohoxMG4EU70BdmYmbpYbpurYtqfD3H4oBAoIJKiHbZs59Jb8HJBZsmmUoIOH8mZ/14
+HkHaT6jJ8rnCuorRJkFbbttcSIVdjp66qZAVQ0EGkpqBSkYDEiIo3NuLWTPD2Dggo6lQVCW28EH
JS23ofsE1vsWAnWllhfg0jTawZEBC7MFT00Oxt1X2RMOhJ4A2AN7bqAqjf4YwfmBu5GZTKWBly2v
llJ857nOi8JZWcBXumKZtgD6KI8peIykSKHvZRFIFJBquqRcAujhQuS/GHLmaWti3WrQ+rRbDGCI
RxBR5bxppCjTcYhYPuUe6nQ8AYX0bOTSaSoF3g8PJwmW2LVRemYs6W97yYt0t3nVGStgBN3LjbmK
pw6X594wcGJr3rMc+82eu2fE99kDWo7yJW4LJo8TvYJPf7J4xNm/yYChdPYWErjY3pJv/HHZlpfL
yn/oMdygDeP/q4Y13wr7SEDNY8VJ+PsWuAWsoO6fvU06AM4ea9YDfGGqZS2xUIaULsCR0v24cFoJ
Yy24EqfTTFmuOeCW8+03KCMfu9tzNRFTsiYa5TlQQXyyylYHnzQKDPgUk+WTGYNkpHzGnqyRTN5y
wG0ctnEq5dfWyQUunpcmeAyerynhKip2Kuuyyj96cidevcnw/PRSB4Y66U+t/UxXJ4xKi31wofWj
5whvoewJsCV5omYw8w6Xp8gYnHvoaWtEKi+L/ieoxylkW44zR41dXnNoe+/XiFhXvaVqeuSsVt7F
uj6Gn+MwofD/R4LZrcAi69CHIS3REDOb7Rp8vWha1yZ1PaqC1nowbGpS9gfadIbfvSlvA9tEoAVY
r31zPG5T4TUf59osCXc3m+x8m3PSsCbiqjCx87zJHEVaWWZB4ThvirKxntYyun5yxuUwH2negxkr
ZORjGV6H8eSmxGYJyYbw3UHSYpDkwJ0SuUv74Y1zZ7OchAhjqM1kxFrlwH/DUdftytlOL3WsgQVI
XBN45T9hT0ud2kbukJRFZylqA/2u2EzZ9XX7nJ3mex3l2/j/6vSjSnxnO1C9OBEdZBikw6rY/92M
knrT2dpoXK1BqzM9tRtjm2BMykTsaQzAon0dulslnO3r+exIsIRgztgOuBH/PilkNrO3vmzg5JiA
PE0FlnUAQ2ltoW0Mw9gaUfnESj9ut//Nyh4tIvZ8lteTBohV94YM+0UV/gyAsQEay/9HTXovw63k
/vtNgTsIExU4qvkGwt+DSJqMi8JqZEG/wKyNV9ZHgGgVdwq85fYbUfia2uCWzBZJokWF9bzg5V/D
KwdtKQhQBGfIEm5bLin0/4vbpn9rIKlUligoolJj5enD7RV2XHkBO4zew8R8XcbrLpfYYdT4IndR
ege70EeG1Euc21Ozb+XJ7sZe/XXHZAbwy0kFD97A1Osv8KuT64yzlG+iVBcyLALxrTGDMEDKfiHa
YthM67bZniuTjZZ3K3zM8ObdXR+LzdRrr6OUtKZ63nmum66IaHQVM8LCZIkNAB6GGimg+8uLhcw/
E7dGl9BIJLMxxYrhdp3yVLqut2mkhEw5Hwl5aKUiQnqoTvOi6/gn3VDjnZM6EZ+2rDEZFGEdn9Y0
VSxBsmxu0nCOiSeTdU4CqksaxwGSHSFHsnsevWDPzq99rsyLZAwQ5nwSsCixlEJky0dl/i0sBoiy
HPcFzINHemaMhmNpFmfcMDTYqXeRSY7T1LqxNFscPNXqGrbrcXJwtHN84Any3Y7smCl+ldMuTock
0Ae9Fga5UDJ4OwLaznh/unYEm55/TloNLQElJIhfIZq25RCUhdEgedncO6SKdx8lgXhQirwFeQcf
flrGByA01zqskEY2NtK9qxuov4L7/mYIR4Lc4V7AwfRDsw2jj9L0eG/pX+yMPz4lPp9lymSr0SFU
7KAmg0njhV58Ex8bXEkQ8N9yd6pgXkGLuOOZJz4wDyhjot4NvR9khLusIF4kIxZGGeE4q6zDL3Db
aCFcu98V3fNwIfvHkKn8eNGZBgzkv0CRK70LYPLjMqbU5zeEmOpB+AfSz00g+cqRq2ugHmyqLNpw
Nrgex3U+44NjJWSPaui0nMuozchI+dPmGRq1jq65dId6CAyNkLD5uO/Ieh577EgyoDf0ZZv125+S
YK4atu17Aac6DmhlHMK3NfHkrz6xDtaDm9antTiCa9XCm7UQVqI9gzii9E/tKNBgjkXTcAPS/GEj
4yHA8UjRKCf+etBA1vkRa5aGbOVTiRpceOPoznpUGaWOIypCPixyoN3EG89mtBv3kG1l5xwBTscB
ncxu3e8kwJHl4R03ABL0ZBufRh7qGBsHT3HO8t1ZVx4CMNpiSPBWnw71K/QksC4TRw0G1ZvBLWNB
AG4RUfeXhPf/Ctb8KA4/HoCNePTvFoo+vLQpFlPOQBqndcVXyuolHiV2+HNeiOMyMZwvwanYzvZR
1KvjXlXRc040GPnU20pOLkjAKVOZiSkVPQHsWNFLgSTfjFcpdPCQ8BuzXDPq+r+GMPaCX56rsGwD
n4rnGpON7oeX8P84BDgG7+JPvoaqXWwp0BN2NedK6eQLZjfPibgn+nDtPcppBZegUQh7mYAvqse7
Pku/Z+qrhDlYDAeUOMW05sMQ7nS7aj5NOgmxKhsYvzCZ/Y6pAWE42unSm2kAWYcPPNHJleJAsNcj
GdGzZ7Jlq7cV2MuxT75ngRo8L+0SfvysYSr7RCzgbmxKIUvFfwdJK+rrPWBXUSm7IBpRNMNjXFRu
0nS9Yhbwk3oog7kJn976RkS7hS3rdUb0CYtsEKBWCl2XcRdtN6VNYQS7k4cn69+hHn0CB5RYiSp+
BqaCt4MmehaI9IOk99RHskx4x3d973KLXE426a4L8eHkGMUhmwwzrrkwfVkcpF7hoko5Uxt1R/Dj
EEc/ak7FOu8dQsMamqEJ0soPO9fY+Z39GvQww6vd0CMaEr/RCeO8Zo+5n6VjVcydZAgVtoz54n5J
usN+r9s1sRasRwZRkW5A0/RJpRyoHqHRW63ui09GBmAIeue9kwkAm+S+r4i8oHa0RpB+zuqnLWPT
6eOM+kNaGeTAYAkq+CTR1/T0wPAXVC0943ESpUWVmCpq64qIMY/hmHPM6rwwOEdfo8nxCISoULUS
SniziwjDxLI04mDTmsJ3T5KwnCMbs2H5EJLwXMgYmNbM9c3ouNg//bmztI5Qb1gU4ylloahHKtfv
D7sQi+MvCma4Oe0pkosM37cpgjHxjZtVNoOwys2kHJGQ0p9ejRGa3kHmH7f9uWCxjpHKWnJoRojo
BDSbH7WS3GRNSZCXKqmhBI+6pg5hGp36WP0JdwigGCJquqiwHr1l744C/PfMZAswNz6Es7ON8w+V
gWlG7h8A9ClvnHLY3btbVAy02ZbuLZnx1bo+nhF4SC2Pq4pcAufasaJB28MyPLtGpAzspYZybsaE
dOPb0CPPSTh1o47dyBNzArlx/eE6NwIRZUCsR7cEZJuPPGP5iussovN2b0XDixP+C+L0QzFy9z9G
aUtpHKWVfPFvNJH9f4xs8Vx3wTIH5oIZvQJI/ITOSxejnBjCfhgESUXCVJ7HJqTaki49T+bfbIgs
wu7BIrSYcznoORQ6KGxh/II8Ko+lnRKjKv28kJRN1Uh1sT2NsKeLNhEzOXtjmiXBEGaGF0orLw6Y
QRuA0S5Y14ncpAjZp72IQmFfkLzBB1pzcSfeZz9u+N+kU5wQi3hZH5Gh2bAcCtRyo4MbAh+bdn43
q4NsQ6U0rCbvTo229HdAb7KJrVmkGLpVXnVZws+Gw9oSws40yj1SInZ4s1SDA/5gS0+9eb5/3KQk
+RYkD7kTYNLRS1wIDcb2YSQKugy/jXbu/DMrMPgUI6ifKFKMgubUpw9F1Tja57RriFo9ZoA600Ao
1Sj0yVqd1P4toqh5a+L5LOsH4ZIAALvkKh0omIdlGtFe1+rD7Sm2hn7WkJXPZJFKT74Yu5lt37U4
OnyWITxdD5liHro8FIs4NgTQjuUakMrN63HZP2yly7t3cq5KzJ0Eyh7pQVwpo4jCnD649uL0sXAX
AwKNOgy/nJdwDgNwVdcE0DKFVKT0F4GuSrx4lHNcxyK+DYSpFahNi5bOlIbwAVnpz2l5z7WgOJKw
jgIGkcDSUvCqsdQEEceQvGOk1OWKmIKup9ChX49NqyutzWYzwK9P9TWHJOUoPvGWuEXt9GBJDvWI
rFOYsVE1Kic6y/cK5CUkYPhAb37hTQhg2R8igKatZ29UCnwWpqOVV/NN+U4iddyGAL/Dw6tfMFN/
0pZkOKMvreEa+88zrfTi0nCp2TBpszbGCM0HldB4I5pXWF+wEmustKiMqs6dMIvCJjVXL6W1L8Cp
fn6XTb/+vOCSM3Fn+c2w9Rl8EDDdfrayG9u/IPfUAYtALO7NV+53ExuCeS4WgAlVDgapOPr5dAnO
kvuetDfcWr8Aah/8x+EqT9edeX1vB2Uf30/Fy7Et5Kctuw+5V8VGXgEVUS/1pJsD1Zt5HwfuKTX2
NhloIxEDKvR7RnkikBMhn4nAgBzP8Evkqj6qxqhv67sx3oQZk4xODMuJRRrz+PuXx00lQ14FHIik
hWvYhqVKUjs1uGFGpPoC5k3Lupj9oGHSIeGdKw+aqKVVlfAd8GU2RzeUW3sM8vq30awlA3MbtAMq
cULdWzJqBYV5xTydLmpwPl+4Jmcv2BSRftdyWRodXEojtamuCBcgIFg1LqmV91TZwokR6pDF72CL
jOmaSGuz708jyyEEZk+7cxpvCynJv7BOP0QtIq1IhjxiMRpGbf9twP8Sb1TVxV2NkNfgdudHudBP
3yuo4AcbdV+Ma3maXi6R556y9crPKnX9XZ3IRTgrVR/MxMtH9nOajUfWaKRbswCS601tUhhPewQS
l9P0ssAL3oAJmHdVdcEnbQVNdlXaIe6cqW5gyICbgDNbClXVX3IjAdSYYqjQn842fw3vKME3gNaX
o2mJVb8ZORLdMxAioDv2MoDHo+yG3L5qsq08tBFcH9LlxpaD/SbxNwhEoq4DAw7lyZSDOyQBiU7p
uJeBULNdE2JGdW50SI8OByMnENZ1V6D59R78h19lTE1zO2i30ONacW3JFg1jxOBw+njyeYXTiFSd
zudSk+9OpXvxBP3iqifThyRDA0QY0P583FjGRFgub2yB/GOp8cA87xYZ3RQay9cP7drSCX06ZNM1
SKtNBR2J3b+IBzJhec92kwBK1w9VbMJJyclNCSYEmyTCg/662nT/X3vAHnD8ptz0+k/qKXpehFoo
ipyWcFDQo0xE6YyiGq0MPSxIQqPM1ZbYpSjY6FK0VQcWX64k+M4Axp0Dp2zDLqWkeTwWVZiqCtAU
X1D/cwDgZrRdzsg3YqINvuBeKh1QQlUPFPbfEtXyyYAFY/Xr5MIlI/44SyWR1OR7PMWapLbxDvax
1nsnHamruBNLg+KzOV6pzvEUMkQPVwBiwxl06+/6Elfn+rFSjAIwU1If+xFYVb5Tijc4bP0nHVK3
VwexYjKuyxxX0+yYo3M6lyzSOCEULYrTSw/idnSnxBjbJBFhMWwkUgf89FfihA4e4yu3881MryvO
UHc30iwnqWcqLbu/RGPu5ssQyOkaqNJxEtNlFiawl2BB7DU4Xe8OtmlNn+lqVP+8JskDzUT8Jsqj
Uk7irmYJrsymBcqB2uQRKboE87RAw6aHhLyJPkJoBFE2gVvQbN2iDZ1jLK2+uj+B4E36x4l6YLGj
8mxRbYufTSMJMFqLQhjyuwAacpZpDcLd05tA5G73DNvjGZPGy2N/+VtZAbL4IIrHcaFXUMNscSXQ
1uU5w41B/tDLusfHvrRX/aiM1FnweAEPuBNNH8n64kBcorpM0jt/d9yLxH4HlrfRaJgloeYd5yfD
HrRUHfiq39eL5xBvvMszmGYtr460hYGBlV/ER1jHPP9vYmmXLxFquz0vtxq/Icwd5burDkqTBdP6
nru7pQinCtNr2u9LfyXVQOMCWpBjGDIM+xBVkQapTAu+GyEr8G/mWFjsCHTiQeGzy9IBSd6v4PYW
bnvjUw2sXJL/QE11pCs7WhWtr/o5b9jzKTfa+zwdTRA9rLplFpjKypj/ltEpLSxkle+0vEQvSv/3
woNAZVrw9yfZnrrHcqg/ChqxTyOL11EHRkNoXiiBowEjacmAbnhdtVp7n8Kog0bf3imwzctvJYG0
UyQ/3FjcJMk6hRSw/WYC+Oxci1+U3Cjq5J3jsMe/eOl/QeeZGWYe0Doo2tfCYWjEwkMDp9xnP7D1
2viySOM70xQJV5UfJrrgOjPhpT5Z8SrdF+kw0OkpO4m+74DO9yKIGEqRdGALqYjek1ubS5eaYtPW
sskBm7xjoc38w7wBDwfX+AdQhk//FkbJjGMtWUrHIu+BGU9ewT7dh3AcxLs5NcfFj/sJ5an2lKl6
65T9xIn6kglSkIooRCLPZ/WGj8Vc2vCsNGTrtYoibWqHyLLZ6HxlnnBNWdHga6eKmfebvje15Rz2
zyMQzkiEL4HHdF7oijuq7Ni+I+6NamW2B69gg28bbjrhPKBhBmBik2cRidszmXewXJRIwpxwTqth
3TBOAdbsQtZR/k85hvP+ktoV4zn2/Voxtkd5N9QF7Q2I2IQdVaZ9UcCwPVU66Na6ST1QROVZUUG5
Wh5OnktmWiV2XCq8z8hGCWfbptjEQ/FRItzJIeVuPrKdWrTZLe20bf4sQZ2kGpMznGR8ZIpWdEAc
QQNe52RIHdyxtBOLFnSGUOojMF6+N+Z2Pcei27aaEKW0kvuPEl6scuOTBuXu9z6WJ/CegTAzBJVt
VM00lmInVE8QR/0EyjQVoVuyUTASDkPLXOza+A8XBUsclbG0Tbd96f3yRnyrHvVX+asOriG4tdA6
y6WtP4Le6qCBvM+jbNtINpELhGDTqxydh7JW9kyJz/DsmEnIAmkyAp59M0uplLo8e1R1knKPtEXq
Yv6gVf9sfbrvDbaWG3943JGU6QamQx72Rr+gKHpYPVmFWRqXfWeyieFe4E03+wDCWcLC24xSVCTa
BnWYp8wBuFmtCk1bmV5Y57riAiLJpvO/8J48LDbX+9QubfpPeyPfC1HpVey4+y28Rcf5QN3fBJbs
GJ0A58ykpUet4CtX5ynSIjJNAEu5VIdDVIA119AoWyI1F7yaSf6+UwW2P9TC1yYqdhrVReGbPt1v
wbZzmzMiZhXuLeVq6p/p5zx4kxo8piNAifzmVZSJ8T3j0xW1V9RAZoe3T4V2m0v1s/sxfw5IwUgC
XXtDwW5BrU3QHIHaq2SZK7tjdi7kHvmxfkddzbvfAarkOdD5VNuRc8l57C0CeIdjG7r9kWK+FPFk
I8aJXmiNe3qThlhCJLKgWaIuP6wpWQL/PgYXnn4x9g/3PP/yY2A+Rsva8Ityre23oHjTgHva8GG6
c0S4a0NIm0wiEmgZjPGE0iHRIjO/N/EYBcc//7XRM2K+t+YxC63P6aXfSI6s2XvSmbEj1rVev8JL
pyCcm36Zp1ITW9C/wwSJzZJ8wT44vr6s8pO50rgKTeE/cQamOLLp2odZtoBi49OCD8FmE29beEKA
hGfboExUeelrL39B9WqunaBm2yDmuMj1MsrMijfbFXQBMZpk2vqIjhHuCyT8XMP4iVSanWv97f86
lV4V5rOIHyyZUSM0C38CdgirBQeg8EWTSYsQXtxedhRgiDrqtIq3U86GrVy2jooRNrE8wL8ifP2G
3mm5EI8EqwTKuIp4tPxBRdUG0UXU1JupuhNvpeoMTIm9qQM+KcOvISRGF8bxPJNbGJb8AYdH5r6q
MByzc3o2IElU5J6CWkI9Brjyi+dyciXdWis05MHxmld33l+/i8RzY5VZhntDr4clGfJTIJgADLgE
25zDZYcTNsCcGlsgBBfLMgxul0IOurAR26ZRleNfv0pPJrUXPexnUQaFn9+hpKVwLKgtKFjn/ErU
bhRkOaN+XFiVg2w7DhJeHxXp0wjAoDd4Pm+NsjtI5GMhPVOstWcjsalUQ9GrD2wRBlR5T9O3kxfz
dyocPyOiYHyi8zI7rfCXjNjpUgaByJ7em0bW8uozsb2BcYsdN8Y0IqQBT20AnC2KLL+JjBj19cMu
abUauY0W4huFcw0gxTShq08+urCbDaQLelr2J4bk7N/VEj8AG/abnp9Fiyd6f0fMm/SWpHn7Vs+G
HSXpyK5uznFjiqQ8Tlav5pFT9bgmGom/Sf1/GDb5AFhCCppbN1wFQ6cvWLq71LuPlLMkyViKXkyl
MthSNKVJFdmYAPMnBmIKSP56HOaxl4Bk3Jp+/Q7f3n6dWO3SgF87HTFuplEJ9fN9rYxQroRFiBZu
+ULZtUafZeG/b4hYkLXdq7UZB/1zMS4sQK5evLAeBvZ5KPlhrqGw7FhgHYCX1bDobLXHoX7Un1hd
L2Jo+pB45M0Y/1/bbRMvnbkW8HQ6uzGLa5o04kvPH0KorbiEBE9xd2b8gjwyc5LBi2uzE8cRP3Oq
4AeiXHv0Lc2y3BPnNHUOj2RW6oP3MTK+tZio3BmlZrX5b89ueWRFcNHUkYIzHfK2C2wATqLUt0H0
qSsyWOG+dAKFgkWlqlATkvHXUKl7HzfOP3bwGmniDy8hiHofNO+kAUynN2BlVU232xXO2THLBKsH
I5Yqddv7vcSJDe/ls8Y9zbijersMjMiAXGWcgMu9MFjo3BpOEBxvVss5/6wWQIW8ldSNAWvU5/QL
rTD1wgn2ji+YK2qzTNLPXlXQ1UYwIYj70I/aGP2mX5Ye9FJeX4qT4kg4+GH9tyPDZPVdAMwyCqsY
vFGh+a/CDBM1JQ32N+SguK9CgEiUqP0hSRO6gTV4qVp+rbW7ugx2pA5WQlD2GGh82vyPhKDIt9VH
7GiV9rQrwkl9d0Gzh6jTMpiMPQ8ox/f44HbRkncOZ4KGXRs8TAU/sJAmc2qiD0PW7huiFP7PNcI3
6FfA1UsCPfpXSKqLSpCdi0XQ5bj6UK0YTpcrpadur591xW8H65JkODJn8HwYzz5QvDmDxGTfr6oD
dM1gjAU9NboF1Uq1d6L2AZREpgEaWPcQZUGBjhbDxCKmP3D4qSPZy7KG9A0ssgkcOE4gsolkTkaR
Oq87mhRlWLV4AN6PGkercuiCs7ljj5DazSicKelwoxfnlRYxOwyaMs62xMaDTClX38TwjR8U6Pqc
d2fmjhe/nOy4pPX7KfxL/LbyWicR8an2RfrFOt2HrA7LklhbldRRrdZrddq6/GzEta/ylVX88zMQ
0bhwDeCpav8dD2LeFbNVLHK/sqQtoVyb7Z/6yRQyO1hh05u4xkgw4X36m4PNwou40ysCcTuJFLsa
XxocDLU6FAZJYx6kuEL3ZIlr9EmLfxeqB/C02UevNNZt2NrlA5xmBwIX9xnlNWu1YTTkUo4wokbV
C6upCfynDq07qgl8hgzpgFVBbuqxecqpfyR3FypC9DiVtbbldE82ZwYxBygRoAWLagkb+Df+aTsS
3VKIvfbz6/R+8U7l+bsveljaYYO3nO0UmKiRglGHRuWoNNQn7t3eVZ3zLhcwDaLgIDdmNptwDLwN
crbWONCq/1jE36UdZvkxq2almvJAks+c30mi8bWIZEJPsUPZiEtdUz3XbkK55MvgjAIY3WL68yD6
1hYfuSzBXRXLmJ5vyg9wiZZsy8bv5QYNO7wHdvB3Pi1Jr/ObaORjOrzGrnOpsKXgUg7mgjDLYj4q
ZlNC+KVw90jaUZE0I1dm4XMH4eJxErd023XxdZDH57v6Epsny3XD42Mln7T2YjXMYi8OTuvPl5Bd
EHP8nyMOmHSXj0XoV46xfgmtN9oRZkvgVVhkX+hFgX1Q2FhzwBjhoeXHoKyktdlFLZ7a1VszVJmx
4AXYkaPN6FvRazMTqSo6uncZxFAwcyKRnFJG8jrubIWrKVFggbmC68xtBXZ6nF3pQY+rI3Az8Wd2
jhqeiQN/ssQlbl+z+39Agylb0/47f7pcean24ykODPszKIi1yXUiAJ7zARqXbPgaSgCxzIXdU7YI
Fgqt6flDCmxLtsdP8OvkOVGlpRSn7FfIRu2sgVBusOKsCVTqoTc8HHfBpgoZ2f0v5F3rw25QOKXY
e4yrBCdPr07CiDbFLPByAV/SAYln2NwitxPp78j1otE0fPY942zmUYNXHKk5QG6Q5H1KsocxelLX
O7JGeuzu/rfU/icaS3c7P86I7hdQc8PopuXgS+JvZy4QtUWpKkNKDqYsDsYSwR8xP7WPUxky2MiD
J+AbxsDku+YQZBu2GWI+1D0Eg78Uv6fWcKwl6rAwBOvu1R3VlxbivOk636QT6SxwdHvBHCYgt2gC
A68TwLyRPHVTBNjm6Z0DjZsKUCtkH4Vt9Cx5WI7rNhkOjYpmgwfvLpDDc5qlNUONjsKJX6cPwsk8
PmC4TcGLZRRImQMqBjWqVWGLAUv2yFOmWWbU2i6+xoqzaWIrDGAc3gS8Oiiy0ByHjc8+7CU1QgYX
fZfbzu2dwvIWkp+7OO1C+ddrNVzpmcv5hZWHiiQW2TqnorSMHS0NuU1zWPjxukRDCKJr3FRcrmwv
5GMCacYNFlVdMN/0lIRPlXLVRAzQH+mN0DMiMAgjcEQQt4u7/VBP974kKxMofMtYm0D0TtWMxJRu
v94up49anKfA6128hxeD+Q9+3eYuz0SNkRKB5EMk9VK5/s4C5KrC1t+bjBPr9yBUqfWeChTrppGN
mEzJtF8CDmtKFv/E+chbEzNg59Oq3iZlsP8NIZOzbClYnv1SxI/8y/k5YfiWEp6MeMIaRC9nL/mY
3tfQtXgYXoRgUgLmev6sHS735IpFcOWXUzeu48YBu8obUqMXMD2Ll71TPP1819fRwM6psdjvMq5W
LxqeRmdOTYXuoi9Rd5mPGGWsYpEjvG/P4cPpwAcd/OR98Q9Cte0Q1H/XrFQpXR40m5hhLnnaKlK9
F3lf1TdzBe1uA1w38DeYG5MPp6t0g0y4MWSAeQm2ty15Zj8Oy7+2Jvqj52t/lTOrg3NUQpvJ5u+I
uewpbThF/bYDCjfOvt2YSy0ERTdbQ1fFpZL8Y3CN6tH4Osp453ahHE0dTqvNwEdCpetAQDXGgZdq
Xbw5BGBR/Bh06vP+JKnJHsZuI0ngavduHMWeC1zJ7wPteN7hE2oRva5EJdxMHUNOvLTaO996TEtY
nzDrhnW8mKuug1qCd8L8NfLTXAbgV+GFJddP8k1vIPogOqtcA56nrEyFhQcIs8nJvIk9ml5m29ZS
MBszWQOwu1nE7N7dS303yy7mEZ8yOK/MD4JnlIbX7qohAv2bga/OcslSJmjCqoNzbiMewqRF8pgS
0le3anvA9nl/XQuZ9xwzPRTuumNRtexbw6tXfT31k21WW72tYjGuX2xj7338WIGipWUL1gqT4Xbi
TjoBNZHocpB5cGjgQvUV8EJM2iq6UTpEEmWQ6XMYd5bIyw2mlC2aBdOapZNqZHkIlboWkgzHnmyW
4XtRpYYZZ5RnhKqdp/u6cuP+8277uSIWZ2zEXQJzpr8RBLZPg4dUILd+BPa1T8YsB4gBOrzjZ5IC
CAbnaLplqIkEB54PTX0qlEpgKHvL1hsrBq4L9StpZZDh85dewP7ToovdA12OxRwmuY3qlSVxaGoJ
I5N//AU9yUlbV2kzK0dhnoDD+1OlYsgN9qV2rndPBuu2SUYJPvy5AVZAMZ9qi0MZEL6WOz6AAv4b
YqtvsIzzFZyEYck7FMTHV6R1AvGaNcyt0XyxRrspkwDMswe5TZCSFewHbp3Pz7641N173EHxKLdH
Pr2JChWGpK2h1v9ocQZEGC1HEXLtXD0dlmVyoLPbL66+2Q7Rifp6rx0DM4ZWrjIR16EDt2GJ4B10
7iA3eEcGCgGM7tsEbEOPE67/SAhrEJBVYjJtqGomXwMN9FiltwXq7UA4FkyIfdSx4j7qtM5C080S
mOkGR6egVO2rS/M/XtQh01CxxapncZeP3as6IFcVBSFjmHmqE4MA1248lUyjc5eGOhAcmqhMy6R9
/gQh/jWKXninbibrgF/3/auMbGiYla/xIOIExpAzuD7Y7foiS5sfXpRvCC6kW4J11uLg4Nv0Y2+G
V0+Br04hN8L3JA94CJX4lOWplwYCp2mf2IYH/I6zpaHoYK0TodguDTosCwKzGdCErJcI3ExQ4svk
Vqkw22RzElO4HEAAkhqAy+3mmnv6aBjqHs+IKtd5j31hE+gJ2Hkxcrv3sPPaQYguegHe3DLpetx1
29vN06mCN5n1a+t3Km2C34nk/RRMV6B5HqvSqnM4O2tRiXzDRFIhV/qh6bJ3cg44BE1aOHruAW8f
4hlq5ysfdk7D9UML8VXIZSwT1ouKEYlaxGkHMhJ/BnWvK37PEqMZyM7Fa+LxRmsxOtnmFqPOBu6I
I5JOTwQAGWCdDgX05uh24LDu2210rSVOqO3iUgVPdQPHgm8iq764i9gJfExTz7B7kJhYEPPccVgY
5lj/6TH/osEqKlkVA7y0VsgWa2Z98W5vF0AOPHJbjV9ouXnM7si0kmuSEpCEOcpF+qtiI/2g9+NS
c87GaT82wnXvBRsn+jo0HSU1CTijv6c5VO4eKy1dTlHJpKN+PNX4NgtPTLlTVfgJ5h2kBvkAXdoT
FlAqvCJYmJ5PNfXfxIzC8ZHiYLId0C4WpUZ5vH6Z9ykjj8SUNwMXqpGMvELsjB640SZeeXKnZF5M
4RiXmsr9jtC7WBzEOaO/Hz9Fx03cZKsek7EEqYColNUaEJL64iIhi/5fdJ1AC576xfyks6n0x/Wd
21CRuqpr0Y9zKN+X94x3fQddL8yjoNXpz/vMzB6yrGzydyHbOulmKoiAJIIFbGdKDTMCK3s5wZPw
k6N2iRIn7X4x0y6t8WPzlsWse2fQPqPYUr//ImWzlkAddZ0ZrAssEYKYICvSBlEdpuzCyUjXSSt5
bYPax8Km9Wk53nyg+H4bh6FTHbgx7/UsLtAB/Xopi/lxdJaxYS8c7Y85XCOl6AikTPxsaZXvX50Y
CSEt1Kjm3kK5xMtdWv37Lbhb1b5IQVb19D3WK7kkWP0iUvdE//dpXsGNUWL7td4lqLUrbDDEMK0P
XYdwdGjcljOyKVDZq7roNm0NGC8oQAyWVIvf5y8vOMCDiRDMMgzzTj6C1ifsNHFCdprw9ocAoyP0
24B9jrVjOYzkVUYQE9f4CRMi0k0CKXRHUschQu88d9J3Suj9lXHVIk0TIh2iLLbzL7+h3hnNHy2z
VqvM3fZtIPwEbpdQ15AA7E1VZRWQkH37+851fgT4PRlK+542pfxK/O1X0++zS/9YA7VHMucNtJIA
X6xr+o8Wba0KQ2ooWjflt8i3nBdTJK46o/8tfQWj1uTarShKeJPciKN1OUdLh8pJX7yKI7TR0yIn
BbZdGfqlijP4Y0AneXmjdFBkiz7Fm4R1WfTKH4oIWDjHhADFfJ2C+lb4RIfEUPPfNj13bMjjHuG5
j0/y17Nkm19Wa5MW/dOnyCZR+qGEcZOjef1WNTQLoLYafQsg2K7jiMYlZ3IhtFcekOL/cFiSnb/3
LHT2KfHZitcankY9pwGIlL4wvZJCfl9G8fQXdcJX0KA0JUJ+Rx+JtUCsoKbyRLX27nFufw0g7wBo
DIr01TWFjPx8HTVFfrDcaYLM6YlMJMaeRenjCNNu1VRjMwPw0O2pN8+TNLsCLAAagVMEBDsQuA4+
/8AlYAoGwLJymmOzSFUXwYC5Uc1anXe/wpeEsR/RJ2XykJntt7NEsy5p693G5Cdgzy+ZEPX2jwpI
KgvqU3/eVgpEeaw/EMO1r5a40UWiW/ubXgFkgVCGX64h/dxDlEVVUqIoUupzyXfsx1IuPnWN4CIX
tJCfY4ZFSU+aNdabT7dTWviTewjoIcmMJNTCqmGpQbetKtpYlN5mjqBTrqucVAYKGLoe+LK57Zer
l9Zrm4Ix75C+n+cJRkKAU74OYoz6wEkpfuCOyzVGQ/vgyKbXoo2z+Zuq12wQZM+aF+kZca2CrxjI
81ytUdFkU0fJpjYsADPEBze265+s6BIm6QwDv46cQZ6E65ZHxINQauDzcrZRTHwwuGDXyjX/CgpK
tLrSv5u+O8xprfQdSNLIhShMW8cEsP7lFoJIFv859L/8uIl7Y9vJGxoKQ+7HzDwZrB8btF4kPdaM
aQ==
`protect end_protected

