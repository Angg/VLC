

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
aEqvcre4Lyvq+Tt5PXDTwx71ktTXYMy4x/0E4dKe9BgxVOReq4m528LoaLIP6GW+fVGwy018LBOH
jm1+bivxEA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
QYrPCp2aMIlbBfuPNfY2dUNw4w+QKreq1bwTmXohDVK/xUEdLBItloqXSCGC7+jUg/Qb5I85f/Ah
KtJEJyCziwj6IUpMayW9odpLYrmaGSusKTx06OZfHHMO82exXNzudcAn72ELL03w+v3J7Rw16Yaz
qLJy0R/MjFA4OGOwuMs=


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
WY4Zr5cvsgwcIO/1W7ZGRcuOPxuu6EPbRD5e9/HsVO16X368aWkQR33DvIRaKE6mu6z2j0ahwjZs
reKraTCWpXPIX3kHEOQ4G+U8/pfBNAeLu+gHRaqilAs+vw9yv9whz81+ixVCKNNcRWQOTvo30pDu
skLTcm2m/QQjNLEpHtQ=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
m6613vAd4+Ikpmzvgk61cQ3LztOi3BEUS+a/u62stTAr62ac1zeSm3L/nrHzan4UzFg0iiv0fkQI
HlLvWFQnraEvQEyI3HNvXjW3i1zg2bQV+yu1q5XCIXhmGlzOkz2w70qM5ze4T5v98BsjMp4dYmMx
A5f4dpYgpZiFnTGLeMS7ck0fB2IZjiquePTdi7jgm/IG+qLBUBUT8dNiDp8GCdQcgG4HweV/m/jI
vG3z9EfAXam/6EPH8epbQzdWAIlMPFNElVQWIXYwEK7n7IkwPHcKKy8h8TIQQBgfI3+K1o6wVERE
QWtvGEQ9KskjsTu85uDfcWnHbHjSbT9CjOWhQQ==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
akC0NqgvB/U73AVdpjoyhrtNQqSO1F1f7/iM28U3ok7yrD2+mcT2y/A9xisbQ06qgSdVkeeZQ/fM
UEmZFdpeZP65dH8ladxkyOXEBZxMn5HBR6Cc/cxzHpMOCwyqreDrscOV//dRgt/fMDUdAzVx9xAF
S3wPRW/FXBzvZQSBlmnr30bFT/LL4Cj8vJGIP0+tX4O1SFvZ4wHGKlU5KqTKs8dVxLyBzSJGBQVb
pymfPPn1F6nJ0s221XFfFykuFYfHfCrSyu+wvMs87eFK5xuSJUkyXUmL+AeodntlACtqvxNeG53J
I6QuD4FQzVWl4npAqVztFXpihv43QWWvfcc+3g==


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
SbRxC27qGffCE5dqvP2lAKXlQLXs2E8yapa9AwWyA+r636Hw6fp2hwwnmJLYUQJzK+qMT7z/eV8Y
OxzIIxbpnjsdHYaEBRYqwROlVe6YwnZ7L6xK5KKxX53MhhFuBHhAxWp9i8Abwj6PqlCffSngelnZ
dnsX8SbNI4PN4MqYSBwgphTtKUTWu1vfLq7rTdNhmsL/7y528gK8mIQQ5SkILrzE8DHO+vA0WuoB
gDK05L8J22kNnh053JxW/y8ZxHFerifahlKocYNdeEgc4mj1EWLlwOKC3M4lBgZJ7fZnJl1veWSN
xU8ddBWIU09TNJJQCC3Tzn/0bh/v6jX6rkbLQw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13264)
`protect data_block
sZoMNwAAAAD30Kly/X8AAOmJzkJRrrIB4/6hjDndlnJUnnQz0acTCCg/4hKYTyvWzgf5W81nUTxx
EgRQyLVCV/V9RIqj6r46zwqkrXcGCrDYW+37vaUJDMdm3L2JbWqunwfC8sUZWhYKZsowJPc/9UxR
hTb2QkCMK3rCkPAZ3uo+FfEnw+qnNyJOt5eJMgupw4+o8wsxk2VSVLJTwt85U//eCI5NfLCzH/8M
Hm5LiIHL3dydfQADiwjIW9p1V21YKdgJ8ZqvruKcr9MskMZ0nRrso3X9DmS6Ppg3ECg3vKDw1IXT
rofzKiS0H/xSa4LpGMGiKgz38lvIMMr3wS8IpqW7F373yttWUJPIj9OmQ++qrApC5YbbfAziOOrw
vE3r/TFgr12Bqb+9iywNGyL5W7Iq47Ypp45GDkxrhpdEXhWRMpqBOAPEz9tnrGtWIJzkdV2Oi/jg
qNHfkoHGtP+9DRUeByfuZ+L2YI9zvfsagOldejofYfUMl6o6rHzxQMO1+HWzWVs3sJopvhp8Uyy/
EMk+XOMpkozVOzSfdNs4KiGZa0cnvn0foszU9tndivNoRKJLWMpvjCZO4/z/bP9KbOuKa02FzTDB
IbmGJ//8y1GHRY06ypQUXz/oSIInE7cIT4Fs4vrrJ7Y9FUrUfHNTzz2as5jjEsV9bIeBJOcFoVp6
ePG7ZlTOQB7Ds8PSecx0JaF87Qn14qbOxS76CyoffBGplFBTVa3s6pG+K53lOWB/pXuo5ix0b3Ss
B+ZLS0rLGJtDywA4lKjuBcL4roJyd2YpGp5OHDfkqYGh07VkBh7GuIOAUvPIySWECutx68iowfsf
ANYXUrLrOvYFcx+PdaXUvMgIZ4ewoX5okRt13L8Vye5l6umK7GDtLRnUt98AK2B5UgdZ/AduUrfO
NB8whPIh/aum1zN3hGWg1MXUp6uveA5lSKu6SrqAqdy3rlyhwUixG2po4fOfSzKNqFQ5BHDkJkXs
gVT1ZBvTNCg79tcec9h2L52ap7q2DLebcQ5a8lsSHlRI7Q7s6vDAQ980YFzoDZenfVy6nyT8ObH5
z3a4rjUI4UtcI6ieBbuuIFRTZR2EKXkHxcLgT3gOXdy3V8hL+1qLe5oCJ/YQoc+EfXJQ9yoCMmH4
yAVjD+MA2cThiGEeRC6b4cjvWPCpp+f3HkQeGKX6Cenj/LlwtVkdHNzDV8e/9U3/3zFqcGskCIz5
sr39JOuTBWFBiqu1nlJitDQFF8Ffc9+4xpiXZ/4CzEw4keEsCNzhrFPWMQhfizqT3q9PChgWJ1GC
WdIKjUg/MDdHZoIi+r4YlPMP8UUgy0nGMHCBEtPGVLuCj7GPAx1KNWtqE1NWfQM8srFAxDD5zmpV
RPwfQuvTziAOpNbn7dj9b2E7fUF/qcLYtaD/N5TaRGuHua/jqfafAPaUQ35t0OVBxz7Ur8mwFtg/
jQDUZneazxCTinEdv2wHCqcOrWCgHMwUv8VzwDUtK9liBP/7gG4Zme74GSLgNFHuLbdeJn4iEtM7
ddhOtYs80DrsZDGfdM0DLo6t1aLspHh4aKTT75fHvu86qAyJQAV9BBlbBwT2k+V973lx9KKUim0i
CmmJjgbxAFN+7RJaWkvQo0e/1RjxyeSA83nqqA55/Ln109TLQlbIQpjTniyHf/2acseqS0gKQ0u/
zm6T6hc5+XMHUgFaN7la2BOWcuVQmZDnErbvV352KSN5fEgMlZHLdmJwqcKSl5kqCOdpVV/3rWEf
616BxLwNjObXhcm7xwrz6tcV2FfuuY1rXnPrvDfNW+H7IO+1HaPBIZdURBA3BRFDvt2HdeEVtZ8S
HioR4nSajywD/kWal4W6K9mzdLh5mi4+tULuZoiAZNO7pBzdQec0YBxJ2yyT6GJkXso5ouLJjdxc
MDsDTOnvfJxVEqcj27ZVyVmanqVnsiJt8wDKAu+vxyezRYacQB9SI2JobJOKrW57A2dYo+kkgyke
qb8sPRckIKNIIuTg1vk1XM5qBRurbw4cAppwGynsg0QUhISTVGBe5PSBqpF8N/5Uf4b2zt/L+xT5
I+frGmWwljCpYMdPbHJ+FKAIU5J30tu8PJW8sbFZYJCjlLIQl2xKko4RBgzUVPzonWpRFSHkijN8
H1ZUrmrPfKnGDy91L2P0FmATeU0Xj76RgTjQtMW/N4g2h7laNe5LjwO2EkX/iXsnoU2wunTqCBDt
VG7NzWK1Smmb9euNgacgJ8F2Fs8E8RKiTjenmaPbcvqRvfuESzzBFQ3suWKCWRRfGlnz8CeWeN/v
ga0aKGo7UNRKA5LKvSAn9+feLHHmPPGIeb4XYpSXHje+0YyvpL82wE2LVpfgf3N4MMlcc8mBGpnm
kCsr6IpOAQH7g3JFyQPPF1uUgm9/NWP6XwTUNsqOExMqsPApHNnF0yql1JVIfr2o8vZMu1j0goSD
fdKgI93w2EgRH+4R/iRPyN/s6lRmz3EdTxjBIIuA9FP2IaUct0Ehuf1nVTtGtQ02efXdK0lZ2m3p
sgwulrhnAlsH+bN1d8Jg6oh72ScFk8L2Ukria7fXdaBtgrItWHtXGUrKW8aHAYgXgJjXxUzS8Ay3
U1eXKwB44ecloWgLNWS0pmhB7bYxRx+n2Y/TaAQJKfF91yFtUwyEJQlqP3wAoepZIHBUeXrKSePb
xi5iyEc9lOBHJzQePAqlA8P0jxo03ZF03K1ugBSeufFhfVvSFMmPuFSuZ1T4ku8Kx893W8pXD1SJ
yIqstsWunLu9igOV8c7WFnzUNB4ulGXC5VURE6Clva3bG+9K1gh80ItN4bSoQG62IRPAzyoaTwzS
gosU8E7BSkYhdOAYRW8bSYz0mly2elVopoaBsNrjm4VwsS9Y69jZO39r1mgb8nUYVkdW7mVvtqn1
revbbshrLVrbiTCuwzjIZpyFeFfjt7UAhl+XET5DHeR2YbY1ECQY86gy67pkXBZoElXrI4ZMneW8
YUDxGvLPCrjUWYC5syz/DXgcFx5zsf+sXVWWvIBAXnzaPBSkkveXIfekdQgjTv1EuFDMd/Lu3XVd
WLWMPeNeytFEqxT73j1zmBC23sCpXOY7hrqRWuyAVGL99AF2t+SgrHqOkvWodP4Ayz+daolj94bC
hizUj1T3Bj5C1tgtKcX2WZvmpbSXhV0Hn+KGlBVBV91C67DkGrIlzhgykBsT39W2KDVRaaffiye/
DM1VapdmURmgltrztH4BDXBTCYYHeRuF3/a6Kln19CzLLFZcfqweUHV3R/b9TzXl95Ox+guoH6c8
w8fkPCEREJoV8/9t+VuBizFXSD9Esx7Knsvq8hADfjvpQ1WLcnjdpCQ0kC4w+1+NAF9XwhR8W7dq
GE3sxPnDZVLaF6wSC7OjyL0OUeEDrkolYQN+LruKaCnsRI/SNfQpzN0LYnGI0gUm44JXkNETAYy4
NOX8RH6iAPyLcHxmYK+wImAxfVKpeHu5dRGwepSdQVUgE4Vc5kX/goEHa4Kkx03cGIB3yhETxr0j
ePGMrLUEXib3oYHCQwpZ80QEif8GHfQI8cOx7D/vH92Rxn0hWbHhMNG/MDCCwpAoErlFk4tRjmFO
jV3Lmnt36u33gcdwKgTV4oiiR1skojHx5xz3O/H73WlqWAf92Mux2stXLhq3iefbDfhtkNMchaC0
zc6MMR//tYgfHMvY4SAN6NnvaBHUVPhxn3hwFNGOVD/lK4ecoy9hw3mmOO8xqvbJQaHyYLgitDjk
LgtK0pg+Af2BiswuQ2Ph9u6gFWPcNNSmen1NYWbhB3DxXkW0u1rTdgDFZHn5IwAtueW+8H3QnWVp
8TdK+kgfH/2OfQwMQGr9pFVoeLUmE0vU9+eBwYCsfTcLV3fdsAd3fFIaRNgMJuzpGbM6r0WmJ2l0
cLoQOe+ZxbOkZqitGKpxxZwseX36fCXHo3WU/3rsH3EAmU+ddnnBFaqWxeG24zIr68zgdBE8duPw
scBzzHran/26ot5n0iWdujLWFjGIhdwrB/QcGPICsqJlPwX2gFdnx03AfEW85U/yr7JW7SrIuuNO
kAYHqSskoBLYkq0oaoSsBWANf7hGX+LCTWEKXZ3zCWSVPUPU/lAMT7vyoImGhEea0QfhM5GkQ97l
Y5O2QcYSGGCAwZmL8F4jCZbMSZWOKTuj5c666nHzHRp2J4vThCqv6amHeX2zr17n5wo5DRcZZ4dW
X4cXC4B/khk7gT1T8O44yXHcK0EQoF3NWDhxo3X7+BNavS/LEyU12/3Ce6kePE6wJyROzCvbp+4G
btIq2ThA++v+pYY56cEeaKxtIc7N7SvbnzlxEl1bzJbPKRtJat0xM4CN84ejdv7p9MxZ6XkvyDUy
6hOU0hvV7JQczs8Wn/OLZOgNlZPjGfOloYkx3mCX7WCN8sSjNn2Z44zTbzCQP3rIMeQK0p6ahPa8
dAUFCEmW/v8AbrfWHRSU2ea5ZimB7+rSOUjgcXzedhFW5Lq/RSD7nTZXP9BqrVlhtlXDyR1a+ZN5
xiS3vCPwXkZco6AMTd1guBnLPpVuLOgDcX0Up2BcFb35f5WNS/J3t6MOrIdvAo9L/tvKaiP+hvOT
yBPyriypaE9YYXSl7zv9vwYoKaHSHqBGAoTH+zFuAzbFfnZs0oxY71eelFBVZVehtgcUVmOmsVY2
IIfMTZG6MLfNOqUs5CoJ5ZTG9tia++bBUAmbPIQTo6nvQAvv+ubtFHQBf7fa+qhUrsySqcxt1IWI
wr5nx9qm6MTIwsHnnG+f/J0C9cnpjCdrPDTLZLYX2YRyTbwi5WrE7O4dK/Ky8ycsUZ7D3BfWHeXq
TJm08Ke4O8vS9+IcL7CdzIEP749vMU5JRCDSu8OrikKqSZzcTS9grA3tiljouWR8Y80AZCk805cX
EWysC+3uTWLVJpprapfEslGXGGRgKqLJ1Yt9kQlbBx0ljIVBcYIVGZ2g0U0/KxbUHjwvD9E0lQzn
L4/huzFjwQmxLcG6JKRyaDXjhdDblLdUoTKXAEoPcX4g3O0IwJlHs914MQlTgZuy97Cg0audAVcM
8Yf/3dJccWl94jrDMR/scpGV0w1OtI11hFt7jm/uJJUSdvBPOTvpAUZHbUlmBECdaJtToFMEAHF1
G2sbcuCK1PsOkBE0PORTT5QpRswJ936oyheunFgIL+QgCybUjjzfcqQ1QX3leZxisSY4OVDSkZOB
F6nzNiYswcSxMH0yiMG80bj0JPWEpxEOxpSfUxJwOSVJmrQGqZJe5hwyVW9786gEv1XZLIAV+R4H
YhGzP/JVVtIv2v5meOz+zxbgQlkxJzGs9BGzjxMV954MtKPrwa7p112Wel9jPCXaKiga9iZJIaFl
08LqRCeq0Fx+RdolLKZiJPXB0Xow17B30AScrKg65/W914jBlNWVVeMwLiQxJBgOfnpc8IU96Qlo
82SNpptO7YG3LLmuBiHRvQmMFWTL9OkyQ+s6Wk/zaeR/M4WA4r0alhpcBx+7PM8LZG4+JshOG+Nf
LQfTBONER3xXz/RsbWBT3HwvR10es4NnfwL5me79zQlnRtwfZ7sYI8FkrTj91pEfyEp8B3DH2Kmh
Ox0Zog/w8972p/UmkLUH/8Y4PK0sp6w68pA85Q69ejb3Jt3x8aSb/VOUQICai3sbxCdaTsU9gJsS
Qimpj66eH6r9taMyD+9C2p6RLltJlJ5BFhCLd9UnsnmdJG55xmVOA04rGtB5RHvw3GYaYiSY88+K
Tl1xBTse0k3n8K4cJz9eTOwEVn+EpvvJhV1WxokNWpUB9SeD2T4/guIUYNMISAeSfBFFQSfC8NTj
bApJ43Q2Xa0jrTJQWi+al6wr4AB6HwQ9cYHlFWo6QBzn1zNkIjBVM2czP7SL5c3Flmu1m2rOzBFB
74M8F0qv7T6J4dPihBiSqKDWhggvLkhKezqoFV03rAk+bpzY3CSY0VgNwZbcj7MKID2PdFhVa57G
YsC2vlAFSu8DehzH55Z0gw4D03o5YrG7YGdYCxSvdmZc3wUwKOi5Ph8nKMkbpgGgqgeaSKtspTlw
sud9c6vJsos9HpNWS0qWChWfQtf1+YYe0xV3cFBeoVQnVVuXiZGok1FlJ9M1GxX8qT8YFhKKQlUr
PogNGACSxjxrn/SpJnIpRouMJNA8xxplm59QLQRDfxFWJrzcqQnHg8wmizP7TpzkuPEs4uC20Hs+
R28w/E4TrKKtkREPInBmcjzFW8UQbfiCHPWodJMoJJempBZKdv7GLpYLhycS05yPYiDU25sgdVkO
f1IN8Nx1ABCR79N5M1oS0KcxjwPixoC0288n4lUdJ/Gz1RIyqen6m8LEKaIQ/FpoVyd9nIVowKIf
u85EBEpOKZkolPyFy6dYFX1BcsmuO9Up87j6s5aQUKq7ByihAvGTpwfj5R7srbibH7MbOyVmhu/R
GkCE+YcOuZvehhsUmjY87qtOrNfnl7OLabinA/5WAo7IXqOgsKfWxuHkI8BBNG7AnDt4qE5Vdw5g
65UnWrZ2e1Jmx60GYMPrirbsqY/HjZFqIpiZOEicjP+7AysArEcKvP8XEfsalexi5zqwF1H+A+e/
I2oFzXysbLAHD30khzSbWxt32Mg7hse4xj9vIXrBmn3qzTlQVdBGgF0dTDGWyi9REpIk9iZBymsb
MMf3kNJYob80iKXnQmPHTh0FRmTJeL/ySuZKnOrDxSleswbLNzikZvXlPU+gzvUiIlBYMbJb9Rm5
wCmgNLAsBfVj5sBQrU7NnYjQWabeB5Z/rk7n5c/QylzDWNMMKsE50LZKbe68d+g74jVLSR5t5Olu
tCo/Y0kmQjlW0PBIWGzxsWACGzsVc6utDWA0hISUaTKKxwxpqNYsdN3RUlvrHknpEXaHkEtmIEHn
YJj1Y655VeLSUBAlmpuBUKYLaNH9ZjKm1S/4rkSveoVwlsyt2qKCGPayXYl/hG/s8uqJssPYjbFa
V7TDjtEmvgxjk33uvNIBqzi9+2cH1A6cQ9m/h2LsJnoNU6BHZ15fHDqCXrvUHfHgE7Uxz10mCYPd
+5lEEC3iuFO0daUjDNSdLxb8OAiLlG7QU5K59Wq5TeC90LmLp78W/5975u5ETsMSAtBYgUBvdi/+
QQcu3pEcvq/VLPMa4vjGx/h2Ntxcq51lRyGqNnb0JiFR8EPMCjHjZ0MQemlx6AkgTvly2IoYz1RV
pIksv8iXtrOU2qSDqPEB95eDn1O4gmAmjl2YjFPm4rM/mQFtwDuz7tiy+BUFkVgKHCJlTGmB2W12
QqkG2OGeRBQ5xZGj065IN0/8o/AEMD3ZtzwJXdeGpyT5OnGCCaqonUpfM0ESkIgmFYVe2TWDjF6C
7L3lCtcvpizBOKfy9BDyphB4k1F+NxiGOriMeDMocMolNqG6YXriBkPldIapLGzQMLQtdlzLYJxo
s/KABzzYVmnvCbh3t9ekQtGK4UiYOKj5cpVYFMdAt0j58LbHKSjQ3tTkzEWh4/fKizL0Dg+U5MVr
AlKWsWzcnMYvqlaz2o/qG4V+0SgLXJVAmdpR/tdlc0kJfNF5HZgC2yXVkZeB36keNGmvjKF65hjL
umlBNwwyLWai5FSBYrXpfj1j+0haw4PMEaatBytN5kZhhnCAl4Eoj8X3/l4hKV4+3qYXAJWfgGXg
L4U1Fn6+oQtu9hAhceSugQcbVlJvuQ7jUFqbkyt6E3aaKktNX9Orq0dHOthc3b1zdGUw9YekvD48
WJZvAn4LN8CeL0gU/lWuo7GwfZjyL0RlRmtWCHP+y4x9rEq+y3m//4PKfe5/1Vx+mtPoBFh6aIgJ
6kBr0B5iMWktT3fGRshpMBshXm1m3TdiVj6pppAUGg7//C4K5ogwLrOg7cdG40fGsHNtnTVOe33i
qjEaGzfDvc6kM4XTOkqVvLhzboyelzP9W3dEsWXDx5gp/ZJeant23VkijcqMQl3qFjmljypH4xsy
4NipiuULdE24LtgFFmHJJHN1UTmGcHtWhwA5hUPxinwS+q99zxJ4TbONTVcX2tliPoJSISqqmosi
3s83MQbKtihnTCsHPk6TZmV5AaW2QOqc7JQNYENRAszmWksdM1Fmda3wGFEe8Wdd6dS6qxjryBpL
2nE1uAala+zVa2sX+xMVS67nKp14BTQyFTRhnhGOIswcyhEGzrsIteoy6/zm6/0kQdS2b30Lrrku
Qv+3wKJLfVdarYeU0fdHxiyWiVyHLo2GiGSQmFkzQha1vkzAWjC/s3DFo0H9QW7WQu/n/jP/4+3x
5R/LibXTjaP7HlkCKc4va7rQSMAOuHK+m+V7uoYkPyfJGNgxuqzAbdpWIVDfDuQlRP1uYSzMMdZE
CKYYAjm51vEwIcxXyzwv1XfF/XUR/WT20m32E4eAbJrg1x39Wf8LEPjrE3U6N3EvTu04+/q9leHf
vVKmRqE9ZupWiLV0kWOSf0Q0DpfsRjK32HMcm4KBiEelmHuj4aIhbF/JdrWF+AlPs1x7lfxIDJCj
d+qksiIdhg7tX659ultG5Mla3l3cGNTH6m4grd4TeFKS0hIxmxTZSgmj9oEk4HaQ5T+Vup1LB4vN
1N0aSxZebJLWhgNjtFgclOvOYN/q1j11ndZlYgt45khX1JK5BKbooFjdEuOCcCBsQAByVSxoERa3
lAbjN1pD781PbS9OeMmrPwXsEhPeNlQ1M4c4LEJJUF9z0VUjpyFjlLlKmVjM8DBgKrC8ESXaGpud
I3QV3+F6TdUWPoSvW2MZUmzCnGc7TbJRdqmtN4htrwIFoG9L4kOcL7Jk/bbdKi1lOQT1LAO/8faK
F500mECbNkuB0N+heI/hMxLfV9LJUiW9zgBxYBIyk5lgW09lxENRgu2T8Pf5zMgu1ZFMDinp0x+4
2ljp2B1NQ9Vw6Ttgj3NmK5k3n6DSt9I16Er+rC1aHPwjhO0YIL2Q+gkGxU5g3XkVVh6Ur3Tzvr47
rm1K2wmzYbcezqphhVOBN6GLxFBdn5ig2Qjgb8Nymx9P5t4uHcektXDV9c70Mdqk63VyQm5Vdr7p
KMl6fTWMgNONdhtWJvgL7duaLx+f0EYxIPZPzJGnr36TxkXgejP2pZG4MhGvyGvpcSuSf3EaPz5g
3K0uehfpAqkj7xooO1B3b5IKkzeRI1IP8KlaDC0Jua0/rKoo3J21XQhO0MucmZ+nFtGmf6lA87Yz
GQ6QGsMcXNpvzwJ0szD2DkjBUnhAXf9R/AJ2/0NlDUaa3IpIdx8U64Iy9u+RRo6Ywl/6zOtEFoOL
h0qR0O18ZERA20FytNMxKMGlApPGzqTILZy45SmE3X00o4kzcfPSFExmO5JPWYj1xFDOEFvQIvJ1
bKp8yRnfPetQWxQNK0X9mgOSedEmLQmsrHbI7am89WyfPUlTLwCgy+70gWrVeOjVDJGWXcfzmAPS
0FaMnZqpDCOHNtpR9cT0Fr3O4TLdzJm5O0Vx5thqqkYivcOIzOb0dOgUZN+mbSYCJsff3spzz0Nj
ZefVC8dzqmynIRq3xE/7Ia3gAOHc31gkII575ifX5jC++8qgPLMedKJl7NuqVyD3R+bWbtflQo+6
K2P1GuoipRxYSZMpz4Kup/4pwFLxaNOQ2Q6YWefYY6EIEWF3UfdlE9SsfUJDme8BXb8FjcqLlJrj
dbOITKrYuj5BmNL/4mVd/vRODA7ocjuX47BFmMMFaLNpNDeNByIGf5fX9ZWb8IoEb56KXSRqCEMp
oOHGH97arnGAaOnLVmE7FSTY9gvU9X9RhG2Y8J1OkMt8V1aw2mqZj/4W/kxVmZuqa7XA2Sj6+DIj
j4oLnKj/85AlOj9r3C57efvPE419RT1qHtgsMKl9+HO++Ufw3/17dhqSvneptJMgFH0aGykCovMF
ao/dfrL7dk79+5WP7/h/XGCVhXtl015usrAevEjoaTfJuf8ejNwgJHw4nbgMDfbdi+9we1vPGYgW
ILfcBU4O8NwE2mpDq2FP+vAxZXh5+JdOkVAr+KgtGkdmuPTtwQBgmjFKm6vC0lb8GvVHLLGwsGWt
Owr9Uh6kzzM11+7+eOzF7NOrNcuGQJI8+zR6fe50ZzSfycQONYFpdL4j3pAfgryaXQV3QTtGaS9f
TQZkV1/d0e9Bgv9de/SPaZrAugDnrwqb/hK3FLb2rCO5YgBVQak71PMfLeoVNDAOAZstOsIa/jf9
38nfeJMbFS9tClrMzyw9YVmZWxVYpTgeaPR2o3MO6EN0If+A1EWXEwtpJAaZbL4JzuJ7B0rtzV6r
Qz0xiFZfwShhmoMsr6y+jtJn06ygfZmtvSSW/7nMcXE3xuiCwsdZZz0g3EmCl74f5PR+/8/yWl6r
1OtavOZYvRVwDL0Cy0AqdVzr4f6ezViwmt/kLLMuAs9F0oFvDv1VhRvNsk50yb2Cjb7MxgtJEp8x
fqYHNFNuTLw5UwpNNXRcLjpHFcTY9nxbR3C95TgYdjmmnMaqdEmTnU8EDzPfYu/3PNDlRN6VYa6J
P0CT1JFBeyoqRcNKFZNBp0bFAwCXXpoPy7MrJgzO1XWokWhmWSgzAPIxpAI20W+/NgSvrRp0N8pp
Ro8E4svVMVZWDyJJp4M2Pxr2obFpnvYCEwkZLaLK/80DXpqQJ1CfG15N9w4yqYwcoEwAPCTvoUCy
SgVIHgbCrO1FG+vcurfkOTXZnPoTfJvY93e1mPG+oViPf+RAEt77l2CmgX/RRSS0MXlSMcDCVPUp
yleUGihSTjzsbdExOXXkzlkTGI7aoLFgcaA9ZaPoEI/2lvqEHr1TVIt4Hn62IYLx/HQyGvsiq1My
T3VfbRK01VBDNK0GrSOnrHnKn7el1EIEwmq0uNnUMM9EI5hf2QfqMBlFScV7FD9KXuIsC/FVB1IU
v5MnAvXmFZT7IelE5hLK9wLNbrAXs/Wfn8qQIaBGBBMvlUAft9pYuPRFxhAd7BP88aOHMswdAEI/
EOXhTNRGx8TOv4qpH1df6/E9L4miwZsLzgaOlf8myB1DcuohYigNDBM5aJ6WJQULth+YEhDugzGB
5FEsdKtUsIP1fjcOoSQyvUYB6EIw5JkdMj7aS7JQbhT6Iv3slsKgFQoZXlM41j8YMCm3P8965RTX
jjP1xvBEpcPG/PQN12WZ9kh/E2neajryiDqjp4s7nJvX4Ni3ZZossvnMh8CrVoFbfJ6C30pj1Nq9
7p6hRjGtMbp3YiyiniP0UhKVk6fOj+lP7XIzusMmVRmavI2E5bwep98cvz/2I9Vcn0MqZsPoPosi
coqfuqFcr5CkPUxVArtcwIcmTWoFuYAdUUdyh4YiAMwn/Vx9Rjscub7p287yaEgtRELX17HETk3H
kEdEKcY9FCCpdlRWU5xgtgHxUgtdKLO//3vpcA29v/z66QeAuTTJnWYcg53HNchaY2GqBRn/k2dN
jhKY/NiLeoAepyAu5YxCYQP8gTTUEgD7bY39Ek/YMuWIQHk6Wk6S+geD1airgDo1rBU2/6WTLPUj
wYE1mO+h2CEjf2F3hlZUZqYW0jIx7IGGDlN6ETTxdVu4HorAcVJzc8irXjsaTCWL4l3dTlPWXzKx
siPKLvU1hx4Kge6XhnmukeAEvPotH8au4BRC5QNK8lgZfd4bd31S5AtIYv2cJOQVVzA8AHpkoPQg
5dHEe248iB+3ZLYRF7hFdTMlREYXlk+xgyZgLLo+TzpDO6USRU1eZP513riaehaOpELS1H01oBR/
idqjmlP7w5JlVpoCtlX2Dy1UzPGD8HNok0glz8B6BD0fPoSXipkMTnkXIxU9OLNUMQPoWyIeJ2dE
d/RRe5Bn+MvHwzlDBA0EQzzDs/i0whtcgjJXB0jjyXZtRd8QoQFdfdgsOZ3RLAYCUgCw95LbNTfd
O2UVpVrHlRT5l2ZY9tBKprY6BoKeGOf1arAyID+lGkqL6K/bukgo8hHcMbix3r797j2hOG8qLLxN
e/NCaUJn8+POMAmC+ljy297Hl8Uv9my118GD5eY/+I8n1OC+L/tNdx8eLWbBtHwqtTzmXtwCZeSB
/3rgzhgGb6NIO5IYk1PBwUQFOtbbFvl++/PfZANqkGIlQv0XAzliSGeDzZAXVpYvOIHEwevJJ3M7
mgbYRyHKPvTCmOJaHUxdk4k4wNhQDCjP8HzLCa1RQ4nd8d6ocZtyhkhgVwJVDDW/2U5BLCshIjaX
G61yE2MYOyYYCmjie2A8kNrFRlAcSP6mlnfxqQ3m96C1awbu+uP0obhshNdkuldO0sTRwUd2tAgQ
Zr9qMyHI5Y+6YT9qyRsFAgM5XWUHH9RqLsiK1H+XvEF3Ufq3sff1ok79fGKcWPW8EuIlSMNJry2B
XoJPQa0Nvt0QcpqtUAsqRY9DdHsaMgr7vBsFo3LLwNM/ovdDksLHaZ/kpy4HgYELv/UqXye79XMV
x6+6yttlPVsBwhdRGIv31RVSv15/H71rOkLWJEf+bQuPvp9ywAdRI155NZ6NNn9wxmB2X4a10uJx
jnmMhiWsfkSD6yYuwMlh+tpIfJdYezs+a/K/QbhMvXkaaib3c+qEQaiU+smOvhAl/Et08/FlA+cW
+5eWuPh16MKk9wXwf6xwDANFcwVyBcRs6q9DjTjMaQYt7SXWX+noDXde/KGpApOGtGOqDg14+EI1
KsHL8qCRSd0Lst/i3qIeh8t6kecka0Drgk3HQluGeCWpuYQxDfTlHx3Xcw9p4g9XdkNCv+Pq5X5G
fyaI607eTL0CIcMVH07igGm10m/bLiYe+7ehvHQl8zt4URcNXbF3qJMmEltAcS/XZUb5Bcyq/1vp
9pH3WyTBIDcjfdbpht0ENSNTXF4p18Chhw4GsLdpkVSO/dpR5IbSt2mzwBwsUdVdgZM2Ia6Ma+1U
YGZ7NW4K4vHhZG7p4EH7x6ZLj561PbxCmaGLOiAUAzAAA+8k60Go8rAa/L0bvgPNkkqjFvgg1EnB
wrm72N609meSJCrtV0Jh37ua1AnUPXwpqze3uo6U5TtvUY/6nvf5kcG63NXIc+zF7IWELq53E6ZI
NnCITVIqKT0Rj5TtmImuUBgQ90i+cIR+Gf+U8w93XUOx8kp3Ip9OYq5R7UjAgau0odsykA0dtTbU
AWrin4MW2STiKbX/w4e5DxrmtcEqK4JBM+qMl7przzFlaeP8YceRwXYikE3v+jm5xeZPo0WhC8ZE
BSGQOGNwyiwpE52isGPggBiAAnyiB8DJy3DsT1yRFu6m7sz9YaOVcHLCF8Ko9xDAWDdV8aoCETxI
X7sMELmwBEtytejMMJbuwNROT6jEF9lXw3cM0xOYYzAb3Iz99YGANaa2WssilRB8vLawqes13nWT
cB5shCx+ZxVTt6nVo5bGTfO+1C88HM5fvjV6MAiRGhR9+wdZEwE0kM8TTHktsxBoyc5iFzMKFcwv
vsXkqwIhzR+qrBk88/kMA2UcikYXQNycRYL0zkJ8P9GbtY3Ugejo88iwfvmVbx6jrnZ/cL8aaUwv
67sIU3qE8KhzEZAf2rzxNLP7RFj135+JB85e4F5HDwi717z3Yj3rmxwufJgG9ezV71CzqD76FZty
r+EIMtvsR37PjJOszyNcEhsDQt3eNzheg3K+B27gmxOlBjtPER2uTgB0s8iyHvnLT/gdHxqugwSX
ww+hhnJYGJj9+rGlIZRpTJqY2VOGOqPN4yL5e46+uspiwasbdi22Z9XsIMCYFkIfGcQVGsEf9tK+
gcsNlFaeUyjGrl0xP9ckSkZXhn+8jh8o0Q2q9iXG2/upgpSPZetoebG6qnS4PFcGAIRcbDvTIiJO
0xJ6CNIoHKb0ktUE/BUvLJNUUqy8hEu0BYm1QfiwUTDrOnHYyYPPve3V0DKRFQRe1jJ67bBG7b6U
Yb/gr1Nqcm1IIQoejT0raF2RH3jxcoCNyzR4S1xS8xVITBICDECn8POuLTaloH4pBRMvQetqYS6u
2hl+zWNSY3/fXWdmWP8B1V32E+EMukQD+OtOwmKGC65ISDdF1hoGDKMbzAcjmSULLEau9d324s3u
M2MPoT9GFT0+sW0pfuNbZJRboDVru2u9tzcEHo4bUp2v3tPX8RWuhQDE4NYeY8SARlE336+VurbL
lXobInMWehXlg+giD05Kn/B04T6smtjgAPVrmD2IEPm+eng4t5hyIa3LCtjXqr3FjZOCOjbRF/4h
OwqXkdaRmBzMmi/RorB3lR8Sk5mNjbUgAEmNOXLGDQC1BCfS4gSB4yYlNVJIcdQGv8ys5sQT30nB
0GrFJ4f2hyR155WapDnBAYVaGsMvkG8s/LY1vO6DgqMAiAySc6YFqW4Lurr3cq/tNnOCpuedtZCb
cyXZykM30XDDcjMUO87w7lP1Gl1C5Z39CJ/ZLx2jQ1FYz9iWemP6MrK5oTqKWVzawQSCCcnTXBGF
gc3vYY0nLYO178bYB6bas5x1CKvWXNA32yzyAUfFQjOVlAifmnFv6Xme65bBbM5WqktPHYFcKaTs
bj4Gth0V0lDMx1n2AI5yJmOn6agVb3AaNAH7qQlPuBrtSdG24GmEGq2+DxMW5bh2KaABHohgU4sZ
XGxrvzVUdsU03RGg9Dz+groeZ/y1mQOJBy3sAIoCpj5/7oGrE+ZwXehz6e3mb8Vr/Cx8WiLNHYrQ
kKuz+jv8oRqQRGn5O27KtfD5wrk4tKSqg0r7uRVrVGkXIEC+rUw3bhQEkhirUgIANKZN20k1g13x
PlURM+U0YOncXtHYM4ppGZZh61r/T5Hx/OuR06c4OoN6f/XE8ePEjGt23toV/ltnkcGEEf4DlezR
cXs45PeMtBhWCnqYDO+IEjnqcqhEgNY8lzDGPCx1OMtWe5gzEAbKGPRhQlAkNboaZq55trNxPODQ
FVDfDz5tvGupJHJC+LYoj0rEErE0QNdf+xrcEOHzOIndKttBq5Bkx8/bh0wYO33Q2nb+mVsJKkYB
m3YIdw73rfP2xaBNlH2f0VNpt2Mc0pepRNYpWPu48+g/F9fVwOq+IpcMMFo16ZofilsoKrq+yDWw
BSJQV0AEVa3UMxtldS+ZwBeUblU+bDJRvdugB1B3iap7L1dBdx3SDRH/PX+pjmD1rAzSVPwM4Em0
miMeTappyytDU8ebonmoTmYDOPyDaWpNRNK5iAvrXQHgvrI0fhxPf7+4CN3CkHxA9c2BCqDGf/jF
uHcTq4nj1HDdqS/XmQCrkZF8dbLp/3OJWPlQDAfU8w6+zAAtCzqlxyMXR08q0JlbSzlbCaaklYuw
ZAnfxg1uVML1twcSIZd/cykkhPUrun7wyCYpYymFSzJx6d1EnD1iK30HpO5Rt/zEyTL9C8ZXAhB9
fKmEh1pI8lCahhn9K52R3NTgpWhbmSEGVHpxoSWmhVBJLsfrqXSaskosCN1gcWVZ4ZOMoKTOIAd9
nVGrN/xLm6X86r61XFJIouXsxm4BBsu23gJEso4g+nZ0ChaLtrwojhogWr73KQMCX/e7S1CfeUpQ
+pXcq8XJ7IOP9Lk+ZR/BJJKIfti8o0pRcNqrfI2P6qh/Ga9q5xMiwBxtofeyHFVABfI8ALZ0letQ
y5RsYyumX/AXdsDQjsy5SH3k9v3vaL9nR9v2J7BJJewG/YD1thMlFq3i0YXMDlB9fCo94UBlNAIl
OB6wz/xlDTCaH+oACJ8AwmSOZ7dHRjsBvOzmKsOLa8em6XnNwRuEaslyCPnWQn8wChNkxRmsOk+K
366ZlztcpgrbTUJrXaRX8lpYt7rM/A7dSH8Iz9N/XRNRfVwub1/N4gl5sfB3ki/lc5EXROJoExbW
/dw/LAVk4qfO7JZW0RFRdqb8OJMc+6wWrm3BPUctOu9gnBDJ1yL40jMJ1Odts4v1CqWYABp1AWqm
MFlpXs2BviCYaxQAWJiikRWrPPAAU9fZJTD77vayE52Lj+OChDuAPSRblhKUuLDiT2BkntRkH3ZM
Aylcej17NGnX+C8yvnKUYL+Wq2KhJQR28lBcExyMhq2iB8v1kaqkckOpdTZFkszkYVdfLx6KUdsj
lcffJ+K6t8vhHEltJo4BnAoWGI2HHBSKIbbP4+sK2IoWmGtQ+7NdrhgqJ5ZsdUKcCijaWh/yLhJj
1D5kknadBU0hYyzuQytrJHuYaakJuJYZsjLQenhi4XURNkflvMdBdM/NH63C6E+hCt3xLw3Nsj/X
BMS/mG2DZrqkgy8HO/OR6cbOJZEihWOXgvWWCmV3pr2veTU+8kK8tHnbynyoF+OJGSo20Cxu6V94
wiy4JwrQA+G8b4FB0Tuij9i0dMR+tU3EqDi4mypdRI1dOVSiiuvt6OMds3vPQOJG2ZR0MQr3AeDb
0DyOkxkWar6j1bfmCkO9vtX6OmpBqHr7VSdXF2AeKjPPdNLuVsXInO96ndCUNQlb6u1I0vPIt0Li
e2Zd34MaJG6RJDVZdRviVR9ZjyOvmqP0NH6YYn+zhhE9DMjmaNvqvptr6OrARyld3XS7IOJbmit+
c2Sg6vrJDbRNL3vhtgRmZUOFOlu+Pp7k0o2ayfqz6+E0k3x4AyqWGWTRYCnyp4YMTRlL768WrEhg
qnIBMkDbQJzNi67585DbFTNhwulUyZTgXNwe1Yw5wPN7IPNj8eUHoTI2pOhAvAzkKboIPGS7Gniq
ZFc4ORCOHTj2qRVPs/CoVfT0xIqs2T+sJ2/PYSbQToNM2diygKx9TcCqJVTJijIMEOutA66MzEKA
6jy9S5Eh9aXWnGdB3as7lkoMJLpCGfRXG2gHslLWFgdy1G7YbGp/dzTqYy4RN3DzwCoMLIlS47B7
kC1/eWx5Ob78Aks0/prSRx/gZ9XlHdkUAXADVcrDW1aZ7f1IfTFpp7fS1h5JpYNMgjV0mTWEfcCd
JsOAzWZ5ZQQY4jrUFBJp0+931nH2QDTECZ7QYFH0iUE/LuYBsri2NjWP73J5cztuyuzhKU1ozGBb
4tfMjEeqf1LcM0sR8MbcmfVu5Mf6NXpE5lyWhG08DW2drNnEgLIDB5MCS/Ll5rnHqUEYPtFMSKPi
iUDKGxGq6KcPTwA4MXRfT6tDvWUdtPW+BE4Y88qlgKreMLY1x27eg9ntyqeb4KqXE0Yxqsm+LXJB
Fq2wR1KfD5TXE7kSD+dvgLyIEQl8zXRf29ULX1PCo25xuPMaRAbD84qJJMquFGKHkF3g6xqMvkuB
0kfibTENJWNyZwFVw2KuHoRaCVb+C2fx7BGe63jk6svWUtD85ANiwrQ7Wqh1X3HM+J7FdexoJPoj
ygHwpoyxxdu0kGBaG19oRYvC+WfSFBKrB9nBybARDunl7SwhIm6Cgu0uodAdyo/YWeOQvD/BcbQ9
QCKUFwIiuHPSBQoRIEUB8iRJRP0Ij6kwjdXV2H/I+aLc9yg3DTZxiNQRHNsseoBqdo2eQX1MCMCo
Wa8xaODYOOWdmMUyR6tBHRN+9CNffrRa0bKkUnWm7UR5OniZCVujjOHtWt2mQLYKJKcLmZ/cNCSw
VBLxe0l1Z21h4zb1Hyo1iscmd2StjDoMwpVGOmozlQZFpK/Pu/mvVdadG4ZLDtwN0RZBGZAmPyAA
uio+CMHMEH+xL4oe2XqNA8Xp3cAOl6SBFRKsAyXH5uUNfzu98mXQmg2UcBmN5o2yW7FpG6wwqoZg
vtcRJeqxNdHLQDd82Dd074sxqBIDSdNowynrS7Ml1e1jJNCZzaAkZbqKTDZQU+JhR6xeTEsh7Sgx
v6IJhbEMCPkdtC/mhj8dRZUf4D7A93TgC/X25k6atH1kJBPZBPAKpdxBDYm37nOhlERfR4mk6U3O
oW+p7Nh0dPQY0QaK6oXqDGc9p4rOW1iGgcJz7WDOT/Y1tG/U4SWA2g==
`protect end_protected

