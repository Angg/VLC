

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
aEqvcre4Lyvq+Tt5PXDTwx71ktTXYMy4x/0E4dKe9BgxVOReq4m528LoaLIP6GW+fVGwy018LBOH
jm1+bivxEA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
QYrPCp2aMIlbBfuPNfY2dUNw4w+QKreq1bwTmXohDVK/xUEdLBItloqXSCGC7+jUg/Qb5I85f/Ah
KtJEJyCziwj6IUpMayW9odpLYrmaGSusKTx06OZfHHMO82exXNzudcAn72ELL03w+v3J7Rw16Yaz
qLJy0R/MjFA4OGOwuMs=


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
WY4Zr5cvsgwcIO/1W7ZGRcuOPxuu6EPbRD5e9/HsVO16X368aWkQR33DvIRaKE6mu6z2j0ahwjZs
reKraTCWpXPIX3kHEOQ4G+U8/pfBNAeLu+gHRaqilAs+vw9yv9whz81+ixVCKNNcRWQOTvo30pDu
skLTcm2m/QQjNLEpHtQ=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
m6613vAd4+Ikpmzvgk61cQ3LztOi3BEUS+a/u62stTAr62ac1zeSm3L/nrHzan4UzFg0iiv0fkQI
HlLvWFQnraEvQEyI3HNvXjW3i1zg2bQV+yu1q5XCIXhmGlzOkz2w70qM5ze4T5v98BsjMp4dYmMx
A5f4dpYgpZiFnTGLeMS7ck0fB2IZjiquePTdi7jgm/IG+qLBUBUT8dNiDp8GCdQcgG4HweV/m/jI
vG3z9EfAXam/6EPH8epbQzdWAIlMPFNElVQWIXYwEK7n7IkwPHcKKy8h8TIQQBgfI3+K1o6wVERE
QWtvGEQ9KskjsTu85uDfcWnHbHjSbT9CjOWhQQ==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
akC0NqgvB/U73AVdpjoyhrtNQqSO1F1f7/iM28U3ok7yrD2+mcT2y/A9xisbQ06qgSdVkeeZQ/fM
UEmZFdpeZP65dH8ladxkyOXEBZxMn5HBR6Cc/cxzHpMOCwyqreDrscOV//dRgt/fMDUdAzVx9xAF
S3wPRW/FXBzvZQSBlmnr30bFT/LL4Cj8vJGIP0+tX4O1SFvZ4wHGKlU5KqTKs8dVxLyBzSJGBQVb
pymfPPn1F6nJ0s221XFfFykuFYfHfCrSyu+wvMs87eFK5xuSJUkyXUmL+AeodntlACtqvxNeG53J
I6QuD4FQzVWl4npAqVztFXpihv43QWWvfcc+3g==


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
SbRxC27qGffCE5dqvP2lAKXlQLXs2E8yapa9AwWyA+r636Hw6fp2hwwnmJLYUQJzK+qMT7z/eV8Y
OxzIIxbpnjsdHYaEBRYqwROlVe6YwnZ7L6xK5KKxX53MhhFuBHhAxWp9i8Abwj6PqlCffSngelnZ
dnsX8SbNI4PN4MqYSBwgphTtKUTWu1vfLq7rTdNhmsL/7y528gK8mIQQ5SkILrzE8DHO+vA0WuoB
gDK05L8J22kNnh053JxW/y8ZxHFerifahlKocYNdeEgc4mj1EWLlwOKC3M4lBgZJ7fZnJl1veWSN
xU8ddBWIU09TNJJQCC3Tzn/0bh/v6jX6rkbLQw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1022992)
`protect data_block
M6qBIftDNP8lBYmZxRpA+6XBpNpJ4dtHLmeHvWdBo1X/FYuIZggi+pYkIHudsOLI2+w50e4/CLCP
MFyGzo3tOiHvb1Dz2GlHNRF9kQU77KwcHo2cWuXBw7KbHuKEhv/dNoox/CORQy6JwXaTl4AMeW3Z
ZsbfFigDSxJZsVQxgJeKfejtpMLMOPsS6MZbej0jSOllv9sVE5PocYInjiLVaia0969LsDfRS84q
oU0LWi53WYpf+Plq4BmrJ3iGuz7HMW8w9zwBcXT0ySwdob4yy9vsuTBIU6O4TgdDMwGygg0CpV7f
eEM+hqebXUurp0+O3nrtyQUi0NU4zs1KZ5C6d4FZfyJGuB6xW6uC23gaLl5pysKFZCjmRCUgzM7T
SVzclyhc1b9bCWfAAYdCOZ8mxseP0Vc0c1oSsjW4HS1PhDKyScC1c9Vii3mXs5mcLaKhzYTywo2A
VSQ8DD7Z+ZpQOK+Gpa2vOqRGNlMCoD23ttIfZfvk8w6AvQhgUGIsWcDLgTWXYmmqaNyWAgLNoKcS
Z/9v5oZ+9Qs51vGEVAM2Jr1bW6KRP9+2RWb6KwEpZpgOintP+MOpxlOgoPC83mnXGEJxJBo60/ql
aKXn38igFbp/qD7/f5hsx+W7y1M8Ku9qpD8ufbUPb8nqtXKbiqHI2UF074n5b0JPiHUy3q37NkTB
EI83vhCO/cLq5ByxLAhDvu8Nk9h5vmpnCC+MkOwlOrZNm7NoRIBNsq1GkdV2Fo8PSqOTh4Y2bA9Q
FvT7uWfTJ04Vhxu7wRitikboujBZmg6IdZeG4K0eT5bB6b67Po5altQ45kwGvmVKKkxm15dsnY7+
FT2jOK/9EsDeL0yiI4JWZws+3/hkwralL5HjMWziDVG8xxJ0lv/rlGKGJ7kgVJ+Y9dqhcmowa3jU
Ilr7OrI5KikcvHCze1hfkBokKTvF+ZBc63SAOhlq9pUCcwbLk4K6B0yjycxqN28+pvrBU7CCYdAu
rQA0VDqtRjuYezxJLDCiCqq8o6ofR+jcGwQYgzUBBDU+kTdM1H75ZvI/yxlG5oK1ySBGj3kQj0+i
ahFaSQiTcl/P937dnxlA0AkFE0+DCsPbL8P4oTOn61gL8hCoAfLndLO3EsiDrBf+EyjEd3jJAnID
Wxov9r6sfRujhrMCDAQSBxAQs00CSvwlcefphLvd36Ce3FeBgUaxzZDVz+PXjz4fLE27SNjnyS3K
/kjsSLczOF9m0fQ0mR/y/ajSegPJyerfTxGOZAXavQ/xtUz8BYtZwum1urON40C4EFBZQHiYtVoW
OT0+097xPLL+DLcb4rD8bIg3//J278A9FRjAQqdpsP0PDb1CcFeOnZsI1tGTySBoUm4y6KzD2iNi
1Q4wKnozDFxxImPRelNerPChKyW2K7GqPoOlPIgWOO4Y4Cq1wTj4j+lOVMHbqfyAhq2YhejbCCqV
QlCJrk/MS7bVfCBOHUx8A00BaPLWAZaDHstZLoCYKXPOp0geT3Mjsahm9DfkVsnI9e2CiZkDwx7P
7Gu83VBhHs4KNcUvyNUq76BPpEc7+Epmfda/UA6eetv5IaT7nYgUhF6JDguEngeCDl7qxZnvEUJK
1jiLk90uezfj81Lhb61Bem0SaWekTzrEFZZnxt8cJ1xFvZJwnoynM2YF5WdZ3kKRKYCFZBxPpet8
agTprYXXGsMo9FNFHDqmVpY3Xk6zeH7UY1cVtM5ZacvOUO7gekvzHFFaslsaExeKCI63NTnlwQLc
KPOamRq2udhBc0/RWwnffnXpVF9pH/JESMcAuWffnRxWIJ7VqLB7b+l51n8qgE7M7c37MjKDmZWq
LnU3UPtHWys98DHBQdqNB1DZx45ABRjj+SynzyI4umJ06mxtmCtR0sV3gaduSGyYm0bPpodAusm4
XcTXRc/ZV32rTefl6CpIKOROP0shzr8Gw4Z1FjHVi06xTVJS8xhk5IVHGn0d3PpcoMm8Jli2XYfe
Pd2YS6SOENFNgjdl6b71EtrWKt8C4VwKL1MMNsybomYtDdRjVpa8ohdt6afIyu/DcT7KB6BBssQi
rJNA9oRZRHjnPOz3k7m8nbI7SHoP7HEc9rrHyymdmpG+Vk6qqcCNXmXVQg3OscR8WEweAoC0eJ8q
9IiF3q7tm3AHYi9MHelrzOxBMFRWENtvIDt45iICHXiajKtaHyXu92f0DLvT4hI6stv5VeTGLY1M
uIrjKpsCe0DkTnzBwKI9A+d/xsf/V42PVKTuvn4qtQsolaRr7hSKCLLnGVNZrcByrBJ22ITdfb6E
E5Jg67TNaV9MPSsWSBhW6Ff2S6JdWEi38ZDLpUKoEE/WruLyp/yBoO7xhP5e1RSHVfXMLyoSdfc6
wJR2iomxSR7QsnfXC1Aog4XEEAuViU6JsjztvUBEo2EDNqSuho0jZ4+ZJSaGXJk1KZ+qdI/cUY9s
whz8E6uFpYvEXeH7K9kmjljsZTju+t/e5RyIRPLHqCgrlbErxZmnTHSzmMDMlZ1LXfdoA4iVfCZY
3swUkcn3DbhUJdsXgutWMuNXP/0AWf5kPzwluLE0ic1leO2F0j4Gr1VHJJhSsgEQcOc3rqSj50Zo
AFsY5hgtiZq26u1pxEZHOL9LlDRAdI5nwSnVw56dTyl7Lp9s6DXnBKo5TlT5gljrJylKvfJh+xCs
mHu61/PATUeteQDeMK/AEHVaH2cVEUyojigYgaJfZ29NfZK9xJhJX+6/3dbzU770Z//TiOA9urFu
uiIIU+9EOEcn1nGDSM1DwDOqQRWcbClM9upYoIkDHQ/Pgfu5GiR8HOrwd3MiUdzzpba36w30YypS
8mYFIs4Nkci808V+IHDtSnv1GqcCmMi7v+5jqEK8O53lY70HFgQgV+ZJ6T2xrW8LZFPsNrE3GKfi
/yGBxwRg39TB4YRGXopTVici8GIr1k3KeRQKKBAvfcXvsH/uxF2ikLPj6xxc/FyQEIgnkVQw/Lfs
Bni18jpbmy1tje32bhzAU8hjAoRU+qoX2Ibhdn5xwvWA+Q1CK5XmLrY6CJFG6/uz7+EPWMLQ4I71
kJyjNZgwzStSsCjyjRCG/L4wY1lTMZM8/dRtmg2AwWgc8lTpiZq15ad43dr1umvG9/XQSRq89y1C
J/PCNlJP0uXVH3NT7u1PDvF3IuLlnQKqBu1St2K2Et8Imx5dyUwTmM3wVEyzN9V5+1PpjTjPLnhL
AJ5K5NSkNTeb1jQYAz/dBWCHR8kycCs5xr0LUK9G+v5QoQa5vjksgHaXxQd7asnEUWbSJRH6aWfN
cdIQ/ngR5gAbFWHdOgDUmusYy6Rut3QZ2Js0O87GGyDyXf7vvlBy8UiNjWh2rJeHkEm56XiWci17
YXpW6cnBYx5Hl2eJlTtgUOTz8S+nSqjTmI+oq0YFDRyO2EZdoxwV1Wu7h4agmIOinoYvzWzkfZHs
ZvEXE19RxO1w1Mz0OsaFCBXrV2BwaFWYzPQgREksz4rzWzrGyLE0vfB1blpXZL0mr4m/EQ6/H8oa
Yc7OG0z0HX1i1gaqWn3Nv87zGmsbIoEk/kG43Uyh5z8Xnmow6KSc7jWOmaqIjYFZ9sSzZchpHHku
ONhW7AfpsdJoj7RUluri35i6ZLC9ea8fNLmIZ33EpVsYJ9Jdey7IEYAfdJqS2lY3E3vIEMrmgy5R
Lti5tO5v4S1dUQtLPoHcp1GQx/1O9HMLxbdk3aQ8cfMwtCjhCkdgJa4o32V0fB6J/waHUzag+AkY
JnP3jlUmad0mFDM0mHiShXKwnS2K84eLV6q2wrZzxvKCoZLR+gyml9M4OdByUlrmvThsUlQVAVRW
NWdhiIQewMIGJ0YT4s35ETb9aKpG1PYtpjuLbTZ9x7TXRj4HouK4kjgQ2ZTVq3J1ikvHfmQYbwJt
G0mxk8JiD4a1ZwYd5a4yHwf9rsKB0dqq/lpeKMbal9kONYFqt72ig2YJB/kBNVgPdRei3TWfDsSB
vqJUJX8xWAKupOisT1+f1NJDKfsm88J3SvShpJ7PA4oswfNZcmwVIAJB+hRM2z1viPZBFf2PQslb
e1lkUIpKQJSY1i8/n1fpSlZQVcALJvyUyoYGaDUW+OdICOGVecjZwuA12AwPOhrwciib17M5fMu2
rhL15cM8qwl+fO3dDunZ99/jvmfM7JeDDKOaBK3G7zb4zKjb2XmKfs12WZqqHm6XoEuf1OdiZdVL
GYsYLcjfv3VRWfxtf6SfQhpMfpo+tUrs3m6TccvYXPYT6bIHsELrdyce0llhmMlWbz8PLi03YgB1
yzHaifi86cWmFEQUBd7Ax8qwokw7S+S5bpivT2pVwNOe90K3vhvGeDFBf9DBchmcvlus/n5t+fMZ
+9f7Q+OvV5diXn3lmrrJCdpAVeJSmpno56HHtoYtmurs8nZZpthuN1XjdKdq2GI3pewHFcmH/0lo
5ZnWlRK6XZVhNaLVkw3JBd2ibmoDYdW9EAM0u4wF3mAKf24b/f4+HRP9d2qm7UayguwQtUyd7Lgs
Kg4byXK3r6Le2ZIOLrTQ3c53TaPe7hzOXHkAeNm7ddK0Q8qBesa7WTK2W9sKU0aLQ9Dp/5Np89W1
KyMfDuOaqO/Sa3/aqlOBoiM6NoQrBtwtYwBJ4M6WdUyEyTyjUSM8FkH0gXu8rSZE5SRjrL5BBghx
FeoRjIRtRvE6sslcuQkuwUCrF5e1OhkcqfqiUlps4OOfH6p63RUu7wXLhl9PraKI7dNOs7C9gy9y
kjwQVqUXjb3eHsobZHA9JqjGWObKi5J/ets5dTT3q9Y+32a+iBk2oBF1XnoWgfqOcGcD2fUrwGWp
mXecK45hwUaXgb6nIMnXryHjVnvZfsrEAeFB6iVrLD5Fe9gGPtzO712Tf+v5eu/vI/Gbj4bkXlll
vcUCDDI2+aurTq2C/NPRWvl2Sx4nlv+gQYT/lWBHD+eoGyER2chdtOFahCwkaGJSQsxrq9wtkCGD
cX6zycA6nAUwv5Ev0p5574719jbcPcJ9oiQV3/KLTpcDGj9nXO/qdOtyOGMI/w6N6dujiM7poU4B
bKvdrC+UBEk04BxiJBM973H+MrJV517ToRgLsRhEaCAePqHl02Tv0fdS5EC2zDBYya2fu42Qm/An
EQfwBbvT7fUpZ5reWMuV7XsKNYNeP0Zi1hsZclE8uuiIiR796Rb/AxIYElUxKl502b8mbyiWvZOL
y6C5Hw/+v87L/2MLAyLTnJyDpTJw9a267E8DFt0Yov/VJplfK9xiLG/8QOqi3Q4uv/b0aKcl6njz
3VzErB8HlMh+6AXk7kQMmJMI3WyQ4AJEvKBevP7BoJwNlPhVhJedLSFtBK+TA7qQa0G0zf3lHbA0
rR0taTritgCgobN4wwoH8nk0TYfwi59ey1Sr0hsQKCA3CLOauY4r5NjOOCtdib3rRUmOeP/85Pvg
GsVPCyEhauAb7agQ6dr8yG5IS13gXR+DkvbhNVKj2f3nw/PgGoX5A9SgOWuowgl2H0vcmq1ACal1
A6hxRMCX0cZh1cvrYtrKpisPRrDysQIk76gLveyr6+b8GGCDZMw2iaY1hMBrC4S/0pC2PisWBPeM
5F8CJmGTnXztP/ndxtaUN37KuirfNQlCrsBC+EBwCmPwLXAENJVEQ8gWS5NoCEPtHz+N1VD59kc6
5+XrJGH1Y0Ti7YhhkzOmS5/S9dmEqP3BPgdR77qKIZT938DuTyEqVZY2KH7alaNajq5yWDp2BLm6
4rJnXcaujzm49ZnmrBj0DYiwy52IWWmYfQkwQaTt8+gob9eanzZi8dATxgKBarg0Vy3qR5TF+jfu
uoNIxSC6OudJqqiSEMLvGzg+j98UBW2VYPmqI0+C5xxuzaNMKjcuIE38c26WwBhUyMDKtAAfQhg2
DnNfsrC8hLPhIvPBGtOMw+TpJO4+Jb10L5blsCOPebFgK966kQ9kcY3SVY/lc6eOjmzZX7E9RH02
aHXbATPvoURxyrd7S8gctcNiHSSTuVn6xk+CwkrKojFrxF76OOkIi2xqlEv7KufGUxHJ5E7dYBPe
3o0uqWSBrKdKcg3Qk3Lu8QHjQjPJVYl5UHCH3ovFuuc7cy2vfPwbFZQiusvTzFCvL0c9bT+XMFd5
1iqcSxWQUiULk1GtSLnFKJ4Rm/aCFBtvFhN2rR/E6jVcFcQqK1zCBCp4YLM5eNRu1StPAP+YrtjY
iTHq+JhciLoADBpoJg3ptn47Fwfm6mM/L+OPWfz7hokHFXVCMgkLe1JxvqQDl0hGXn3odCTuKvrW
XYRYmYBFaenIGZWD4Pfgh4eET9xMMjaq1QaXwRuIDvhX392m1drS45OagFRLED/cuZXqLNibnhjb
ivceJ7rBNDx7eKZM7XS4l2cL4DEFxnck6QT9ERHd70Pdvy0ybP+jlFDDy/0LV5F0L96jySbVzknZ
hSuaF/gWDtl71L/iMbVIkHZdqV4omLWnlL5LbCd88lZdZMxIoFubgOGkzcugXpkFOwgJLAFjJImT
RLMEtwYpeGtFg41jQmBHCTcSg08+2d3TVGLVRhjTXfwb/OvqyQ+B9rlnQK2hJaABl4BOSYnsxykI
DT8AFXDGnYv7vvmGr1CLjIDqoLFc1zJte2/+5iAFahfhxx1fBF2glwCunULqROhmQFAwvbku4AZi
+VaM6cJF+Qpk2RJ1C7XesFtJA/joVryl/Hszxggvw/YAK3OvwD7JtMJNnUzv4k597I1PqqaptJyb
HqkXZrPhzRX96jU6Fr0UIEsb92z7/SUe0juMAC61EQgArJO2lpWrv/4KmOQtkGAHDshyfCOesaNU
trzSc4wvb35dg8tTNQnYTv6AClKfKZ8ko7ZRCx1s6YQg4Z5wWsyfjMzMnt8LV/PjnAwcpd+a8aG0
+weCsxZmt9pU7A2/QbMeMQxPmov2oAzIUgo4PRaPsVdt5yH0+McWMX5U8FNRWXdUwzcJPL8i0OQO
8DJ25BNeGtPYaa9ItZHCLtC/0FEVhUa+WpQW9M6jcsv+mPcWr2AxTs1YmwkbHqCzK64ViFQPnBjs
RUGPgvFE+HKhQu0fyZkn4g9fBJqx+vsogljlARCCYz7qwt1dVxX1TwZk1pqdUMCalSf9V1UMoKG/
CBGYXqDzOR4FacfP4/Hk3cLzMaTdKeY3IjbkMQL2NpmBXpVT38b7zp25OS/M529/yphBKPS2UW8y
MqoIXhM01KQbGyLN7KMPk79a68VNP2fvmJN6gwW+ib6ISj1O44T20mx7ZOhs+HwHjambfuEFwe5T
pOSuy7Y0ptlu9wtXQkWW/kgFaVYvbAHobYEqSdWd5g0pg4HMhsP6jziSfvOsGn4+DEg25yOQTACr
V3/7ZsEnlpiN0/HoOH/Q4gKW0P5bca3AAqbL+gFMb5hQRgDnTpHmlU+ouzfuqC4r4U1i0rQJgwZS
zK/+cA5QD86TkQGz0vwGV8LEsQ4mBtdh+FkuSWUI2ApvMc5aGz4uzWwT2mF9c66zptyRN1UoagEs
hhX7NjnJIhDd5budDl3CH7Sp5SN5cCQKtdicoWeqhv1y9Y01BYPdLjS8nJoFFtz9FgnQavlxKGO6
G+P5XsBv9HWezFgC9ouUGEETQJIfOyVJvEzvS3at41Q+3NuRociNT1dUaYB2oCi4/iszHBxe017Q
H6lhi8FilzP4TRD2P4Nkyx8wuPF33DtNGY+rvyi4UYkc8/fGtiEG06tvAAhqPhQ5e4VLfsBHVw1y
adsVTSixbotdJDBMadD2RhTzZFcwlojf9xrhUsk/4t9PNntwHuDe7DtmhCgpybJSChVkGs+BPfcV
N7Z7LLqOz1rYQCLi90HKTbPF4H98WFvvjvR6fgfKmq9x1SvbfL0voV0um99BDf5A/FElg9LxRrVx
Xkb1eSyVyb/EWob9lmSLSZ2HYSMT3/2VHPZ0UJcSVxWsr2qI8iOC1WSHtFioygDlU3m7CsMbP5xb
BDBxV7K3ZJCiWA+I6raqT9cPwwDiM+6Xk9RAQBMxA3m/5KKR/2baQHZOdmkY3deWw0vhD6lQmWCP
VlkfEpPyEinw2jDKKsAt2DNiJlhnrHpPT/X/mmLEELB+U0SqLGIdqPOTKI8mIJwLuFU3DT5LJAb4
DFmQx5VaLTv9DDdV8HDcfzzTBUFEXLfQ/acNBFm2HzYcu2yi/yBUwgm99CVCEF3EHffckppF+7G4
ryVaUZ4XZeuYzWJgLNJdwDm6qAz/C17N/fgZq8EaAkGkjJf7PphZx8P9/Hu4I+dBJaNp2nprxnD6
/zImRaeoInprr3zaVUQ2EoGk9kl9uoMrTC3p1SUzHim1DLCxHsoUqRs3P1IFUn0T0tNHfyUiNO+z
h7ejfos0Y6Ko1NGqahHgn+3cFmlJzJBHDcQ13hWStkSh3VjVdMyTc/5yoXDcfxo2/R82VJvv4GEw
WW+uHflh/FKvV1l6Ui7WlbX5NxkgSWmEBu3prEgugkG9Wy1yKOeSSSCqh9WTTUN6eynJg2oxKeu8
CB1yKWh8IewfZhcPhLBSfavbE8uKVV6Y1ME3iC3H6iIVf2wEuXWQc5JzvWBBted/T43IZx2zeQ68
t1y05qXEhgwUULyp/iapxcdD5a2WW6nNqURJU5UmCpwDbrNqSNqD6sJAaAeD14lW+DYx7f0MNJxF
1RUKRBJU5wcp7ou90rpc1nvJ4ebuSzGLCi7SsIQudEK/zZSp2+enFWBr05Ury+dZloFSj6v17Ijc
ePkJouNWWWccafhWQKLbsVC3Cr3fH//J/rjwV8kFTDA6usF1kJRIWX9NRY6ukdecHQJUS8PrmswP
kOIbVUxWElNmT6L8LP0V08ZvtR+NmBG4BJcG8ddhb3RBgjDqyBfvkgXAiAKpw3TStPSgMKZnUQLQ
ELOAE+/BeWdxyO3ki8dUd5ja3+eThC5M98fjY3ieSZogx5EX7hFJxlv2gob4hFDEB8S5vVRqIxI/
dkFpwVgiOLxYFIVnOwv4toXCMTaz3IIIGo5xedJW05u5MP8sJIuSsQo/ZEs7hZQGnXRWoSFElIYx
ns3L39SZfWRBEVts+GcP45D+jOMRoScIru4ME6SuyaTzMIUNO6HsWQE3emrp8xrtxi8AFTaErhrc
tjHLNZFrtjmyN1Tbt0zLNPPieKd//gyK7mflHFS585jVqujP0Wz0+p1xr4D+dTFikjdEdVM95Aq0
EcMEuA5ww3VNIJA18LP2XO/GsmjXH7HcaM9SB09lhQki+bn/0EXXFUgZl+lRX+c3z00qHX8PeOWP
1UjcBVcuyBHF+CiD4VMCeR/44Cggmaikrmferi5xCcEQp4Vpz41+fUsTcWtD5nQ7eUDqXhsdCATc
oDH18cPu80RgLWdAoGHGGO1leIhQYqGD8jM1JMtZW+VN54FKxZ0JT8NnYSvGXNgxFVjyf/662GCM
w5PZNxuD758bFim2+W7fU1GjXCUmIL9iDVBxiQ+sSgUqbyCEHfjDnGpHi+q1zVL+jmICOlVW4ID7
gbn94swJ0x/RCX7snO+foEQOFo/B/pbDe2IJSieu+zZdKBJEnttLe+dsN/la1zws8kfkC6Wo+OSA
xGILJ5dTS71h5jSMqrbbl4D5vQxDUqrQMqwqu4OIIW+jbOMUX3tRH4NJFa5eH/NVAjYCimOvHPjR
bfZUKDeEZUkndrx0AGSuMjrwaDIpdrux3hzfbIM2hwZZ+Ab3VpmOHhCqDiWWIXlR12bigThDVSHo
WXVHLLXS20mhVaQGEhR/CTCN16oHN1CiJxQ71vxvLtbRExSF4s8FkhcdpX1QceCtkv1k502xi/7g
HdAxAsUSekmHWMQCPmP+0XCEj+7Y+xLqE+5ixdPm2A/FHGN+NYBUu/RzcX8MTS8cehYRC07RigTt
pOIjWIBjZsG3xP1/h+MyEzTMNdwdndCjB8VzFV3GcCOCqi+fLYYXjCI/b5lPsKrdDlCVjh+WAyGD
wAtfUxq3obvS+O1hGNOA5uwwcDQt54zKxsi4xvNEnWvxQzdgyhppsFaAx9bLA4BeYRosfogRguIf
T7cwcO/ASgw8E4n4cdcbrCqE6x5MZOc5NU2ASr9b7RtF4ZnDkYIp79OoXdHJwEBcVlQK7oenCZIk
8LT/L6mwMNeO+W3Zu7GC5YYGaLjLDRrdeyVhHuKGo9RdpA5+AwwA8erdTnGcWMB5rv9nuauuHIms
wHJHTlv/VcIClOXde/0eFIGe0kvP0bT0HghdqS0EpStdbdSWkbmw3T8CbMlHS8pRMKMJYUMEjklH
GEuzXROaIejuX8nIJUSgEBCOGxFV7uhh7ga0cmaf+2my5MKY7pHSN9HNnhvb7yWLjY+Tbo4nNLuX
Yjmq2kE3k8uNObFIbrMOYenhzbkyCsRMzdM2r6J5AFVMFkPPvgWh2Rvmi75Ld2H8/QsOjDtEnE9L
k5hgp/uU/dIatxEBWgO4aH5Y5FKMiWgApKg2K9O0SLAtTT/3ZfvsKXCZa9sq5rF7G/FUWlOMhWJx
AOgx/16GOE/J3tI3jVyOuo1VOIDp/CwEbVPIvcQKiPnU+YTZDOA5C3KkjmyUofZ//b8dFUjGhQHc
t4CPrqPcY21nbDWAH94c2DxowWoZsG6cO+SwiGjJDLxwgJzgFDtT58wsc5CnZ64RQjaWm6RxrCVT
ny9ZLXeTZhS1cNWO5ktTHYKwug/Tvl7kQJpJRAlpYjPIoGmNV2xzXcd8TPRvoQ3qpqkgew9OTYmM
OhWJjYXm77KQeTXhDhyCWnYaXLyMECvfeAdyShY6pA8yT9TJBpnXXfRfbqG5mOafEnDG12x5YmQK
gjhVHZYniAm7V8Vg9F0SGVV/PYCmik+eDkSZ4dURN4j+rPqWLsWA1rB9qK02W5+Fvqynbl5MY5El
t0908mcnrIRtGw4w1qShWdH9nlLoP5VEY/snPuw+V7vEMpOYGMEWmK/vRJyV0cBHDoKGJstAhjOy
47xCWOMBCCMiSK0bb5UWbaB8VFsdXAQH+Oel3vvXRxUTNd+KZswYkADShxS1RSSUXmHsOYQLqnFn
unahfM6xpAEAxlgjU6z5cSvBdBD6Nf0jHcaNEWxKa44y2aagWIJ2XYUPlTtcWqm2SL0md76UEVAq
ZTYUPbCnMk0wcY7FnzcIxbqwwRVB0C4NfKHVWAUiW4NGEfDbDLcjv4Tg64sn4kZ3HhsI90AL5QyG
6ENAPMa5OZ7rHtPBBpguo9yGOnUPH3r+BG4opq1jFZSBwBNxwq7tmzVw7AXqoGP+SkOE/DS3F2dn
EgZwtOxopp9KiLzyfWSOxzpYw0kFZP1RaGfrHV7vFwWF0NvO20qOrc1ByNAUpUlGw0tSGUyOvq9S
z9sY0CUXp/WfAXu3N09nxoYGWScutLkMnm0GiF6wloS66ST1mVBofoK4H26XgersA+gsJPKEa1SE
9ayH/dnKle2k4sMxm1vdwja+JYw9y+yTQwGk+bi0kltDebYjFKlyCz3QFKMDrPMQ5isvVgFbvJnH
ccsVFINb23F1iV7MCH4QSpVE1pk15TNSe8SoqHebgWI2Mxc+ruXXC5Set/SAvfnQgosFS7s7EK/F
4ZpomcooDMkT+3osPrnItc7RjzyYmFnCgTWzqslB6y7+QUCb1kVrIHTEnGNqgE47WZjFQzSh15ei
NqJRvJH61GRpAQVu8Wxup58y7iHu7XuVp2jCW43LtvfQ6MJiHjCFs4dIOF1oYII73sJBKKCVApJD
iT+vpvW+FMgmJjchqzl13ZK4Kh6UM6X7vg73v4BQwU0nyH9IjGQi3qU3UL9WosGm1kDGfNrYzsqf
Db5LlYNKOIT+i5cdyZxc1W5tSqrxgegjzsCBuYidtOZ/Uut7a7nhJ+754ONrrRaFy4FMetWRRKhR
iMK1uen+kunybklPb05kDgWSTCaQkiAEMwRbnc7UB+lBaGEGRV/DMKY0JSqlGa3Q3TZYmvTbSuCs
H90yI+U0VNlxYDRzMpx895alvLX0CSne4xlJHs1LvgGyECYCm+oYgxjTngF4WEKvVlv9iU4R85oU
rSl6rBfSXD530sP8pARxu6sHXZeqogUxcYIgOegvMb0sx64G4T0pFbAzWrWYgm2TLnCBFb7MWvQt
60aJLq1msY9tzx0Jx6GTUD1Rk6QOKFHoshdLDePPV4mrOjj1By1kVWiJSv+jsPAXNX9YHwSDaud1
5RXLxPExRd82MwpfIBRjUPBDZjn79GpJgSljd65VvjD3kTCtnMMVmbG3M68T43pSvA83pZFeiOIK
S0c53WInfxupXl64f87j2n3s7TbDS5b6mpm+fN549O4RpS+YnE2JlQmix+oPJGfoBsGaZjJJ1ToO
eJ40T1XzKLaWSey86iI00yj2Iw/HE0D1SbSHa5yJyK5DRrErgOYFqHav8EUiAPRimx8aLWAVpeVp
rhDEhuP2Tz7BtEQ6cAZWjANZ/MClOjd1niXE6XTKfZot8qE+cO4otVx6ljFCOqegYf374pIgrdP/
6u7m4/AvT5ZuOPoYbupV2rdEkfCalOSm5xjwtb5PqVX5tc8/+2316RWwyQ4GFhpGllOJgT5VhTov
m0Mr5lhP2uN1+FnMjTCU1/irx6iBgttiEiWTcqyWfQAK+qWJDSrKoA3Q+DqOj6gly8m3n1wfIZig
IDCLGp7HGlgq7B1yfuDJj8wofB9ZOzgsi4HZKErn9sFXbtmofi5FwcGNxfwQkU3KvdzdSNTYsgeU
+lSYPo1vAoYFnxsi/xZk//oTxYORUJx1oA8PqSznjcSk6x68owdM/HxpBhUyLdJoDk0i6eFoT29A
HcaB8OWSjv2FeISmDJQ72+9/oM6sqP6+MYNzSyvuGL4CmQKfyoyVtLkYGGZPecf3AqvUgMME+QkM
XpLZOBgaulD0hPqgOhMd/QkxWLNXT7vkoDIPzGZKY+LN8VhRZ9GrGujsEwHuFM4bMomGkHDAlyQk
SEsIVguYVqqAo776/uV403l/AihILXznWn4hOkJ8uxN54G/6XJKaOKRBciU5Z5vwnTq9T3EesLIZ
UPG35+vNd0DimjiX9gfEOSYCKrk5cVe5q6LnS4bX4r1wldxu7knSM8f13QqiufeU8tdOhI9qrMfp
UOBPP24XkQSC+t2DVSHKGD/P57NM6DXS1VpcMGOZiYvMlXQTqv5ZXOV281p4cIC4cmQiFWijQdI8
YEOT4DpRaVRFwJByZDhVQIESaSCjtz+Czw/NOY3Of3mMnwppLp3GBfJaeF+66kK5fVlx352wV2c8
xqHmrdyJCj0if4S6I7cOwnEZpBT5c+GjokgGWyxrPnazIEXeXymDjXD9xkFtS+/UhrFSZULCaid/
IJq7iFB8HGcEJz6BSZxicydgkkOy8/auseMfrTYPiLUyRYSqbAnX/NSx6idJjYKkVdGfhtcrJ6i5
csqfDpNcbMwcBe71RoBS2Qjy4EkzxH/yC+XlVr4o6sEOjg4s2Ja3ki2QmPAQuhm3i/JwHnEUw1ni
e5po66rh/TUOZ7HBsBcRfn1OWOEBWYtWob9NUycm/SwtOsqmiO6RB2EULWYuA9hefjLT6MzdoVAI
1GIRaoMuJw4T889qhiGLmf3qSocpG3ZJZwSoSlHjVTxysboGsViwHdLa1kz//9P4vARlikwmww3Q
NwHDCpf6rVUnF114WNokhzMqByzbYgPJ7qs0c5cquiCeLDrRO9ogsXkGYjYSwGGsKh0pw7DmDxtD
3TKmoxMJbSIaU0PU1Zvd6Vu20hxoDU5+bv9/pXWWEHTOWnZWO5HZegC9/XONrSCZNsZDBh5bK57R
S+VUsDetQ59x5HDmYByBDtYehnwYyr/PFkbVMYNSNDRudfCfPyQoo0Pqbt1LyRSlkxT+m51IXDuD
wOsQ+pxhnsw6+rTlZ291XTGU0v2fKvw8n8gxirZwduMkNwvMSLrhVmORZdb8BYx+tSMjLGk3hEXu
HzHRfLdTIBU4GukNljkjFndDGP+8EdyZPvRdov4FobrisWp/+cZBBSLbWadZ93r6XWwd3d6KvpqS
cwvuYlwelLrG4PUW7irNlOIWMRfH0VW8aZGMvGLq85vvDyRQSt8MFzUHUTLN2ydyqL3HoZScjxzK
9nosipD3Qbr887R/OPCLBHKGLQLu+Z8pz9WVGD7BABhlaXK5m+KvLijo/rV7h5vGGYAA/boq6iTN
NjH9zCa0bekGDo+cYTE9DnsNEgLMvJoCfqHjrVp8IyNRA9dd/JseTK3LgXqcBLSSXPIpNgK/XXVt
MfhP9yIzyCSUN3xkEygRnfGi7lJh0rNEVpr7vknBwvfh62buDPv6ChOGf25GFtE6AuvI6vdjlxUS
cUo8TQCYC3yGXLuev3A4FcpOJCCNwfLfXK0ATI2irc7HYDGNtq46zm4++jOoyH4K6bBbXg7AALm0
q3x90xSBor0i2D4NO2YFnuD+AOQHVfXQg2+qNXz3T3MMO337y258FlezQ8nQEKL0sJbY+b8J5s/F
/W2IPAGNfAjL+8yFZIWsrRu60L+pJk1J13dFmmV22SFD+6HJiBbzj5FQP2Pzdu9r4fpL3e1RD5yz
uwDZbJnrdha6Hil/mfNOK6Q1RfXWRzg1U17nxK6/gaL30sLuG8N+1T1bogmHeGCNJ3iqXtuKAyvT
Q/PLcTtqkfhv/uDwq8t5r2+bSYydmin+M8xyfqYoaf4cFGk0fkfdsmg/RuYUvADM666KKuqSW+eR
HYDp300eDfQUX58+kvMjSviRZdH+UVWml2IWMaRV46bjl7JrjOxeSA3FL11xu8IHEhTtKYTqeafY
yrxvn4apwFsgAhvqtmvBD5fplwSDhkST2kiLFF0SMr1huOe3EI+OgOCO/hfFVbVks5WQ4gBC+kOc
gvh5sSXN+mU9BFAOfDWLG7uKddDEiMyLaUYfX/aS3NISX8JGG5xXIEr68wVtHDuxUbFnXQsE5xBn
dQC458b/BBJ4ddwXoQiMGGzpn+2QPNq2V0icGNS/w86YpzyDdVKyXpUPE+I8EbZq5UiHqVNXBKvE
GNZAvSYKY2bzNEitdOtuFKluU6oCzcqo4A9JEEnqKJXT9igUpic4OPy0zS0+3rhyZJQnMdCgQguJ
5xKxieNlziZQY7PafCOmz7wRzk32UuZ5cleKn/O7htaYQtsbEhcosHJd8GpjjKzQkaTcQ0TBsXPq
a8vNNOb41BCLLa1//rpvcVoRsz3/+2jJ7MvEB7Pi3aq/EvZb16djefm93hmcG11HPlco79n0lPKE
8pk2J3FrocVX7Hyt7HrhPCXtojXSNTd6CVpIxl+dsG7ITnkGUjeAFMZqzIcMsh72AleL/3QI3KRn
91MkKKhwQMNN67oRZrMS+OenpqDjcTy0Y7rLkVcTPaMeMEUwarywPWKAtODiuTC7bAA10FJ4EV/e
raH0ZHDlIM0yn4dnpLbQeV+WSbTmhyv1monSNXBXeK1Kwrl7TR/HLqFGd6PAYbIP/QrV/ZQ2xCEs
fiXbexLJ0zc33L+MfUVbEr9QbDqwlvObEVQgfS+hCW8X60IYL1knZpoNwfGo/+nLeNWZDdlBgczO
3leEb737l7n/As9L4g8IBIaiYZ2eodDmZ/tHwG2X3ws9SPat4fGDI1//huAAAmicaVgZTgf2/WWg
7vKgOm4kpWnUxH4bHVd0GCT+pc2W58OHG1Z4hA05H26+zNA8voFIUgqIhb7rIQhODKr1VFpg2ktD
RVH14UVBwP55tjyfkN9yastMlemEicQ6xIOVXvUu9S+5JlaLes+jOeDkg7BafR2MlBbbzl1ryvck
KYPcUz/Ls/B3PRxmDIR9w3zpmNa5nFVabo07nh4rkKJv//p5YTpJiIoteEelAvhlCAYi1Dt5AXFc
J4JVEc6K2zbiiycd9fF7pyPzNgwWSlbf1/wG7hvYFuSzVVkSPRcmU7MJbEwKSzk24vbwvSt9EQa1
7zpA0bzQr3OlSbdtzGyLd7en7O4mTC3V/nCnetOdcwFCQ6/pQkGLCIz1xGqigXMy1SJmTQQ4OyP0
jDfm9f2J0pKfr/BLAKp8RMWU9Q4+mmr71V05i87AGSn/VswFv6QIgzhlp184SKpMgijTE2O82pZn
1NLBfYIcsMbwWn/OwQUCNWNZsB57AWSr6QThqbzcWIOHQ7/Wkxnsc8eNDlh3mhqfVnu7ek1OgE6w
As8IdYxoD4pjWCPikSITeeHSfdgy/dqbUaHPWYlJCjBdEW3AyD5YABa9Q2wKoxV8XhESxt0BjkuT
Jj6hOJ4W+3+o0eHU7vZymQ5VFpeWysTzi6bp21yrVecyQtxn3LRdbwzeZdWWZpLlYG8RccmYZToY
zjs3qARMeJgtf04JLhN88GCyERh9zzwZPKyDugNF4sal19Y2dfT9iUBelYwY1dtsFZBQDJTg62/t
d1NwK6jp7rM35JPN9qo5wGc6TxdzGKY7JMaO4ef6QVyg/UXb2fKycUXe/aoeZQ7tuas+jjh9m86w
l+nMMhEUEBEInfGqCsDC60NXDiwF/L+c0irxW3LmK2w8K1zRhlo6tl8oSQTkM7QuvuaNiQn+kPzF
ywcthMbCWUYwelwK/BOuZi2VcJF/HFFqXOssaz0X5ZhRmaxqgwfHSGOUlgEdgra3m2puiV1MJkF6
HcTI1rnXkMsHML93hieq6+athH4H43u6JLzRgG/ZsVaRcOMP8lq435JMJmBLyhX0VdL5qmc7QvXi
G96z/MVmA++UZS6mPN6gI5QgfHOxYzu3xOgr8gv/jOFZS4J8PlMbOsfOXYtBFz/vn623+X0IvZSr
GoXFzr55CVcgFJYfcg40ZmLLYydqlN4Dg3u29XSWNu9oWLCkicEpT8/pQ7/cqKXJfaMERgO8fbLP
T/z3Mxxehj4YXopScDsid89TBKdLjdadaAYrE502K4tGBeamTJllgATxuHF+7fDzkwbhwNfqsGz/
zIZiseo0AwugUHF+GUk1Ei9/NxFpvOIET+9z2sAQJ1JJ58l95EKgABuayskplucsvT44pQnEqJvn
pgSWdsTlJ8TIC9e6QXvgyZM3wvSE+7Vm6N7lmz42w8tovwfpKnMuqhnlQb8sKKdpvxxjYQiJSZDu
A9++5oo1ig8/sHpghLKtwDGOE2rJ2riHCR5LpZMjjnTbMAobYgJbZN21PrCFAc/lE32rooxaAfos
Lr9+AgiNxtcqX+rLjWj2alAKjLksCBtx1c9IiJfNrKoLxZOYl98sNY0Ps0ztVJQ+Ln62Ibv46LC+
Pb55BY3Za6EYmZY5WfIr7inPSDG/BKx40NiVQLuJZNWkKJcrANR2g8XbeZTIcd0+nxyDp3hXEnVS
EQ+nZFKmTDtmyBP5QumCDqDTEOBae4rM036kyF8t7ronoJs4CYUpnMS9vTNd2TUQv1lqdRytPGIE
qbsYj3+AEoT9+CdQIU/0ZK9X8D68eCJS9eaUQE+k1B1KqsL9iFuE8UdcMFU5wc9rtYG6oe4AzdiB
dzi2T2pxjQtHT0Jzg80EnKQWHO7OcGh8/moTeD/WozOaZcvoAZLYA5SRPwCEz8WSU28v3MnLjya1
L02XV06HJ5zWxlLaaVD/NkQhMsQrEcys3GtZE14rOsyt5BRYgWTWz54XTl167AzwK3zUDZZ/3ooq
7lbVFLE6Quy2jz5WgoiBRRSQ2thVHoUocoia6gXgkAmx8ukBZZOLlDMU6TKSPv+5trbFKs+SbQCr
XhTXLEQbRn/cz1Ho86vQig1gBY6OyX0APc1SXi6wPMGRdzdt7BBN0k6i566/YAmMNEWHfd56CX0O
FkaYbEDHG89kS6VKG339TcusnwO3lebmE2cc/zc85SC4NMBGf3BCWg2940EE7RqQrmeuKUW+Bc+o
r4NsmwFnNlWrv7EjQ1ZOvQ/WJACPxecoXwnrY4D70PaGSuHptcMU1aL7HisL4RCmh2tVAoXGPOOq
FZk9tCq0vd6jyrE/LbQxIcb4NBlW2oJzPGGoIVAmNW7Go2mdlzd/LUOoRL5bxTdDEbAYELwzWcjy
MisLn3mcVCGc9kOnHKSUPlTNeST4cEohlNKb/G7WdWHMKxJ7HugFc7akV2Abmw2VGV5hWtJtLimS
0FW1E6TGsuUn6HJzj/kDTsK0lSjMMf5ddG5blADWhm+YWIhv+oKw5DsCeox8WH6t04SEYKoYhP0X
OMtOnNK8oXtCE684R4yZEWVwKNJD6xMolEtrkMN4KMJhhiOI0bja2nBGS2nJ5ZvFyeU+TTefCRPs
e/hPUxOUKAIhHa+JP46hwHG8MFn/9b4T8aTEMC8cXEgGViN8QM4JbjvgsyRNGaaS+hXfmONJIN1r
hSYrCvdqR2caDatpqtaTpi6d3OYNqygFTAC9EegA6m1lqbcbGixfRei+hgZoZTmtkU7NE8Nwb4Pb
rpskgDx2+hg95cOowlD83fAX83s0RIpCqs+FsbGD+/c9c/NdCBtlG4SczANFiufb7gFGKP8atmy8
t5lMOBIo3wL5bylbbYpxukiOFc6kKTpCqtZPhMnwvucb7tJ2RdDOBIXn6Wq7nkErELE49f3FKtwH
mW04aE9wC7TgAamIdRJ+ASejsNnIaP6wDMBlb0cBXym3iyzzWGH7Q6ctDaMWLVnZsjgNusehE5Zf
cW54KbN6yJV8Gdyngqn/Uag6IayWCpj/uk68WPxbDIxracp2G4j86W/wI6yFOdI9QOR2zxyEOoF7
GonrvLV620uuRS3kIwtAIBu5/KUNGQp9K3e+kp23mRbBIiNIzqz+AewyIQSvzSRMaYfKFscL/tSh
+/2HjOdCXwUsqQl6rMGU+ahStPT1vR9W2ATyOJvZ6XhS1bRgFtvMRdTj2UH8pTjoPT/4+wRk0TUC
lqn17M9MfDut6gEIU3ziFjmPlBjIpKOLWZaFujj+cUWmQSzXJeoE3bdzRIRALPUEUD9gIYFZHxAm
1yqr6mqoAusRSxjhw+fSpc4j95eee1suL6DO/2+MyvgQKFrEt14eKM2viI7/reluC2AAhNv01jfP
830QMqaP4DFCi1F9PV9bXnlO4RF9DWOmjUyHUF1s3e+HOWzr0/KLb+vm+phaaDJVhP33owym2iqG
meyy+xIcPW/E2+NTr3R5mpZQbR+a287CyBomreAIQi90dpIf9yzwTxG9Yhft5tgexUS51pyD36Ma
PVkeURxbUaARABpVQZaCApPhtwlR+y2NNe9Z7POU3emwG94yV5HH5shcru8uy7j5K6rleNxx56yv
TlyGOo22lxXuNUcGIlPY7nfY1LbpFC/uHfBzhVwRMNW+OTo3fINoUwIT/Miz6k9HUcivodomCbG2
re7eU61thfdyuTOCejfZLT2D5vQ0FsjCc+GBl8JkYvJG6BTj1AaBHExB+KuCyWpr/3iEAuQOesgw
OOV7b43DprHpLCREiwZuy053qtxVM9vWavqaO0yvCVp6FtoDJvUamSrXaFMwmEKXeAnq5c7nuYhz
FDQ4ZeYC+m3WlOh4IQdbCP4s80XZiP0BWlhpznNrydTRE4LmVvKL905JfPcC7uJTYuQY2ooeJTX3
Z7BQ7qtgxTajFh9RtQST0C95hrM3XDnK6vTq94r+zDKaluzTO1QCjkCcMyO9a2Tr0U+btJEA4Tzm
qJXG+fufOlPXHyHSVue5IhqtkOxMZzfVNO8TRQDRP+ECrCnZAcoHTAmCaVhuwHNRCO7pETm3ywSq
vdtdzB5DSzQeajnOQbjo/cQ9MV7gjzqEW3IOUCW8Pb4HXlNUjBYdISNeiGk0H7vBvfvIitwOFzFC
A1TjvijJuuLT/qukaO77uqnojjBk8j1tP2bmvSodQw7rMgAlDhFmBqKjKVPNzyMiw1sdnQfsAafy
KUeyRKunUS9AmGa44vf3Oi3oj+QSUe+7M1uFCEeKSGkVOqfynFxeOlz4X3vwpstkoYDreAzvEprk
az5NHrLk+ubxkefRtVTI9c436+OZcnd4+CNFMzKj7vBq2iFeMCuEeFtXNAtqF/cqFOAyTmrt1Px+
zZA8zNXO79UkiZSgzacnM/t66cDWlTB3FId4xKRa4ytkSoKdzEOd1DcBO8jtXfZDjf42DXslzKg+
1mhe4AHY0SHaBiR7DkqQ5EJjpYK7IdJwlW1cbNlr6My2tuJKSVoek/a6Zxo1ngOmrfUv5zrpufpB
wieTtfExx54c0eMRDD4o6vNgAjabnbuPJLHcC7roz56+E/OQqt/jsJnAVNogzaF6rg/sCX0rg4KU
7W1xgGKaulP7Dqe8CB1u5MnLvbBRU3Vk5py7GMAs/Yc+BDNWxoH0dYrSklF41Ez7D3luTtvuFsrP
P2U3Z+Yr74dzrqZsFDMUCgftr9Uy7PCuc6+F5Ia5E1bjnaNXFZkYJWwXcrIdmXMVD2zLS4gNOJyd
D13ok8YaJGPUH4BOdcAshFdKzS9yev879C2MwM4aMivyCDmU5BY+DhOXpPxllbjR4XH+nsW2rhd1
Zz2eGmudVvCtK0sRmCk2T5LagNFOgV1FUg0CIjCojAtIvdwR4KlyjpzCAxPkQDegX0vSbp8POJS1
FN43BEA/PEabYiaN3ZFckfOEhDZV5aDvy32Luj/wtBEKh5I9zUDmyJQWrzrZ2uER8IbPdtj2TYYZ
ZOSiRTSSNhQ/F5QvTBTN6pU9b/bGolafsCvLjC1C1qPgYQ9ZBOEOaY7NXQaFe1X8zSKBVOcwDD/o
UlT7gNTXouK9/W/oH6AW9qInoPA1lCB2IhfbeMu1K9ZBROz7fKQ7JMUtftzZDiQDZk8aGXkQMC3Q
2RrtcLhOioNOU0BtxcKSG1N9sXBfi+kAzfLzOfJD6hGgzltVhsT/WCSOUU6ye5FLCj1sav9UKDRt
0b/tWcCaaabpbb5P8khiInHbv731H9mx5p/PsnZ2ExuSWOoQOrU+Q/rvlj64JkKdP8K7Ig6tcPkU
dgLCuUGlZUVrnxY6BUpvJ9bcB+3/VzqeWcd482xOurispXCq1jTqsgXSuW+oV9smbIlU5UQoe7tV
G+Zz1J17m/8bCsO948RchzpYtcrb6ih7Ip4Cvro81gQneLGbCTiMY8LPpFq1Focgavfz2qYK0tOm
669IVRU1Co0Ic8WAewR405I8iqsO4jup/kXUOo425atrtXIH2nLIQy2jEWFIEUsH6HzDlbmhmIrl
EjVu50ENws8XHX3f1No2RWS9m0j7k1gmxYnTd4OpVsT6DvaJ58/O7ojAc/oqpjRRDZ+/At8hBih6
ascfhcW/WW7JQbQFQzODBxMouzsasfq2PLAMkcJoMnAK3E1jOmMMVdNgtMNYPtSQnVEu17jkBDlp
DwyFtChzDM/urcH5Xw8j5y2ojunSvuWYoK+wFW3qnmYnN12xhtjdpvJV0RWIeX9e9EgySt5H47MD
rw7jnAkNwe4+1FOrQtzOoyFcyWhvMvfPFpxVdXHTGQCxpKcveE2a6NIm/fyEuJm4L3DcAljjlZkP
ySHCR+9jwMmHl8o5+epjurTMMzQh3XNrkwm+Zwz3lXMncyD6wQvj5pCITiq0b0sUUfJ2ODRnO7QR
LBhIV0juZMZnToJgJqw+KGz1N4aio0FeXdxoxT8UhMw0SHxGmWAaqi/Zh+rPxpddnvEHnpyhuC7Q
sC18Dh8FybuPTCm+a8Xj1taKjM+EHGMuUDQYxophUZ3T32CrsHa11aHisoR5tkFRZO1doESdJlrz
vbUvK1XGwM7MhPV1FpUdbbOrilooiVsh1Rq+sbAT9Ga5+NwxIwemeTP2lRBZdMfOLGLuIaRyOEJm
A/9utbKDqeeoChk4ukAv+s1p8q7GETFtslTeeCAdjBXQX4kGc5bUZixGAgIqqkXJ0pa5HtK1G9Y+
qxe/ABYAJ4HLMW6RwI9wQGJ0dJ1ZhygKQPGWI7zejiksMe18uCBL5/PnBm6v+F1poabPI9sK808O
WfuO7XAJcVKv0zAW/Sf+U/Y5PuXYD8196j3pluMrZm7pgeyyEHd3TTHZEeqv+jc69yO4qjkYLkkJ
jnMi6H+UYb4v22lC8qRw1izaDVB+23EeJQhZFrQ/yDegQQV9N3IatW7WdYNO3fTrv0LwebMpPatS
HLYIcHXBVG0WXhzpvk3YXeuIRlAd2D3J1Fy+2Y9AoqJA7BI/26zL4bdUSUdOjOjxmuqlcIfxqZEM
16zTZoZd3tiTqvt2VG+bYaMx+iR3/KGsDrVgev1cECamE7NVPYmOnU8S3GPouHeCAJlYh9JANg8B
8Ifzw7BwSbguEDq9Y+2p0gN2QLyl6STNIGvfKjADvWr/dyrpW6x7kiOgyc3ChlY4Dn+JLATEWNsx
+ZzYDPS67SUYtMHHPOv/kPUwcXwQdI8sWI1ktM2O9vhsf6XoAMdtSzeER0bAb7FOd7uLPvQV+Juz
UZMr4eAD5q8KwCWZph6Wusp31qS6YIWc9tU2Sjuv5ZohCtGoRfKJT2uZ4mwdrde4y31L4i41A0DA
wodlhF3eGUTkBhqM4bMRsBrcC1sxR5yZqMNHufKZ4ev1fYm+bAmOsbAo61E7fIzqT39uhLh429NR
z/wZ9RkQhBI3DxFnZI1lVgibuADqNaPLJLifsG1GqtSQL0ZFiTJ4rU2gU+kj2Dn9GkOioCq9MoAG
8rHn1NO6YCqyS934nCdcuyJNAiz6uoX1H/WC4rpUpg829e196sOjXSBja3j92auh5u74O8ykhRXT
N0lDwlLaw+NyjNqRlxesAhgEW0yQkclwEPA1hZ7cW9hnQhuLQimiDt8Zpl+Cx9IWdbORCuTi0n4T
TYGFRgK3zw95adGTmkkvJYAvG6FI01GywddqQr56JCLKbSk5XeIDHEniZltCJwyNSK46M6cJTEgy
Tx0uVcvf/ys0THKq1kuL5PcQAXb8cbMuZ7ldltXWpuPkgSCi7WHNSVu9+tcF7VkiWS4Iz17gE8md
yFRF09px6xIjQlANeaUK8EN9MzUDxySVJBuY97AZOVsmNy9ltocpw6RHutB4SO2xIc/qSoK6kUzi
1GleBqwkoxTqIPsi1GHQSjS0W2qD6fr+O5NxabsqjIsRnruGS70doCAyQl5YYUMc6gpQtXncV/IR
qybXNdklf4bTVnfX1OUM57vWngeh7DNQc1vqRgPMFZ5wp6WbxP3ZAt0LbBE9fpW4S690QT8wTMbV
Cn0ifxU08VQsg0BuIFPjiR1xnKuxtwwguyifJqmvkYlY257xIccA5VnlevLZHzLD1gQ2rAb++ihU
m1ZLvSwJVZGefKh5p7dFvtljuvQmQgg0pUW07e5ykVCLdkU4qF7a7VA1QpkDx0edEZHxxZGzIfRL
jAcuGRhaGNiqv+WcLPM+ShhT18bNgqcS7T3it+j0ZC/G3Y2jFA77HjIiQm8/28V6NYLxtBOZqYgh
nExoXBEtckiN4arZIMMCstG29oyEGO0RQy1Z4iJNKH1/th0nhl3yX7+TTACIyHt2wQGxrufUMt66
22enobsXgeKJ5F6CZHuKAcjk6JRbosOPJ7F6b+nLF0HLpl1/xw1/JWkW4tW6zADJFcu1QKPlIxAR
z8UuPxzeJcpmMjp+fiswl8mjuROnJLx/0ltYN1Yt0DZiQmd6MN6gNG05qImKsyWDYKgjPJ8Oz8FR
voOJRDbvM2+uSIfz0LJqLbTbfv0+my5E33OXeWdS1/LZe9BnZfxhhTCfR6eXq8o7Iz5GhopFZZdU
lOAZcY1wx/xDwhN5XqnrqcfNOOCTLyLWhhdkHBVi2r+cvnu6OP0DmzcxEBrVVQjGxC/X8n1LSLMS
rSD/jX7Vs3p0sXets7Hq+Fq3NXvvNvvtoTy5Z0Yfrlpk2EciF64TuaWKFYsteVmNX5f2beGmbDaa
Yg34azxtQF9DMjgQTRpnPk+6Yp+uEaA/ymkSOGg8puQCGj27DSN/MiMHBTv2B3yRDB3ex2kr7T4v
9mhIjPMrlN2+ItevT4TVV2hEhUf0Owelu5D+XT2NiWiPToKAKJXEUOv1drMIVkDui/jmrdlmf2hk
eV+1pOi3GgOQtP8g9TGM7D6BAuDlabp6mD117XQ9egOvW/+QKxxT21RToY4mdSNxw7XFoT6kadq3
poxE4eLWxu5UFqw2hOe22vcH684MpD58GqP4i8g+EjTUK5lYqMRErMtG9oiADrWN+t8jSdaJD4k2
ifd+3zZzalbjZOAJWQliGMYXHEscPLGWioPyyhKFzqUAeITggxdRgiKRiHsPyFOjSWlK/Z9vTZXj
OGliFpl3nx7oc8Bqus/EGCzy6WwnptkN7OnZP1hTwZuBYwjFknJXNk5jxMWav47TeMd3oE2iDhEW
vm3qgbVsD/OIxqZCRPHMgbGRWRgp4WMOcqo5gLwLich/OML37WJhUUSOFEy2iFPSowLXuWilsRiO
GQSlqYhFlsLxLTfqPXiH7kH2yX94HqYNbdLOGdzFKFkKaUyQ/ypyPFOvhA51tDDcw1MvK4lbZFhg
gGZatMexBXUbrThvhi3WUynOal4lT0DrSHA/zSkgMq+u2bmYri5THtHk4WLO+VggbEDQ1gblBlZi
ziXvq+WYXQw8PiC3eFStZbAQwQTVgjGdf6Ddq/4BepCLCbb7n9K3CVqGYXPYvKquaMKut8uSpB3j
bStvDvlpFKIk6VeWsRoS7PGL6rt+vi/852OegjJ9A1tnJZLQpWg2U5Zx7e2lSwtWoOTtfpYoWERJ
dWpP0HsXslSldMCAszElAIaNt8ShymeOyhfuqA3xXSGBfWid2RYUyGbiB2PDlxrbWAhKYI7bCGvF
X/nJxuegfVc7ahVft8yEIMZyrAZTLhIRxQb8pGHJI1RRSTj609ocq+UayhyqI+7UpEcu0/cSBney
wT3FdImdg9H3tyOj8eGRIiBvlkvZ2RO0sIbz9x0xZtco49h3CuSVLMwXWUXZxuqlR2VLSp4VEAWS
HXZWAvPCbERyCKhVsUrD6d4E0Vh2Cw7eRwVBNYUgNP8+iZbgErXpkueUE82J67vX+g6ijfLTQx07
X07RPdhOXUnste0PakkRcCv0uS2a4eT8bcc8i43GUiR/ort7CQ8Wurms0kJ5WThrB0czLy8DzfOH
jfQ7nKKc74E5SyEiTMeFqkhOPUOw2E9S3/OtkQwHdoxn3BdVVhS+3gG3EF9DgcF9aYSZNXQopxrG
UEm+4rCM5zRNy2T8MwSu7cOeGfX3xRvg34+RROnApbDNyirRkUXqw+7j1JPtYbwgHxDbBSIuzOCq
7ZBexPOz/IgSu7astP7hlBlq+8kGRNMuKjAFyS05Xs8IKH1dsEYv3ObFfnlA8ikQ6zSKYkYwY/ha
+ehK4S8YQMQM/x1rtxuK2erhLLYqhMRT4ghUlyLtvFrlKXHaM7QUma70TuXIwmsIFeerc7QXjRxZ
pJYAM4GEGb+NeGhy1VtINSN6aSkB+2j0i2wyEB1tIz3I8Jclbc+zsCtX3dcNpCyiSmm3qZvDAdhb
PZbGWTuf2/ZHmvz7eWhKNCq2pnLQJxnM0yVHpbxaFKVa2hSeqWfh+QDNfkYYa2JiE8nGo0JN7+Jc
XU3bPCu9z7jJxwEZZb6P5BXCJ6kkRo48PLj8ne9CaIberC3b1dZCBOlYhuA5Z8UKBt7u8X4+7OOg
2mpkZe1bks1e5EPsT3Fz+eXGNCmZ6lfPSgWMYYx4m9MQZFeOc/V9rooaAjbESuJSCbBvZ0Ffnyw9
s7X0EC2LLnF9Y7Kdq4RQHFGnZf7Xryb5DhOEmG6RRaJuYGiOdseg2MZOJWp1rovXRg01qwFMGN+w
2XKVYdWLeGwOfnlPvQZTK3nhtyHfzLSqyVqK70LvHa7/nQJAYdaeJNogsGaJIy5X+M3/NcWWMFjX
msWc9wZZzEcyZcWH6/GGXIUTU+KGxlE+x1jMKyi6Oz37YpbsFaj5xwicicjQMPUu71rWsdZqMFvo
+jf7DxBSeNl5/mDu29hpWKbMOIO9OqUX3X9ydcwgxIAKEihGuOEdQDVcRg39Clq6vUOWi42fr5eq
Gl0uPnCYTGi8elX+qppCJ9ivxT1TjxNqJdbEDN772ydCQHBwx2HgW3yQUc2Z5mUKJXkQSAtpj6tU
oBR34yADsyGFAI4kT6rvcI6S66bsI/KEsSm8QnatnhzvY5I5e7XVnkeQLCih6/XTrdE6NObiSx2u
8awMuEg98kYlPS5P1zYUVsiLnF/U+4z9Cgy6T2PqN7wjz9GGIuX2Q+aeDFIveSF6rcFj4GL6GbxQ
pwQ3iX/RzJRZEw0HQLj99Oa6/8Vt3TIGmw2f2r2O+lV45RYBndVk4KuDTyBOcI4BRU7xKmmIrijG
ZnECcRGjCMGAomR/frRJkdRfw+q/oEylhpxkXB9ueAcAMa9Lx3Pkez/seFojZDQl/STHQhhhTjC0
lErPuRvqfOtaIkdiU9/52QTtltHtcsOwrYDP9IDHlCqTVTMwGHB2R992dVp5fE45v0I+ZyhgE2Iw
dbBNGEiOtgrcQYmGYJLvklaxZcRWLZ7obOfGIwDtQ2+OYMXXFwd8a0VxolYZ/lHTbO56oEt9998P
fjuU7ZKaZqLjH1GnV/M0HT1C1t6MG9Bk8pJ7Ce+baUmAnquOJv+54BcDh3qCL1hzCZXDhWX3TFQA
FDcBZUD4PeYBb6+4YwKO+XGZJremk4UcT2tvZ9qinKk9LcF5X9GWrS7jIEQFjn5grV+joNn5Vofz
U7REurUTUgoDLxsKLpagYxwLAd8nYoCb3RpgtjQnYtxWEb2FdtsAEPIVOslDTEy20iNbHW5VU+3x
EjCZPi4xNymCrJQbDZf8pnApu5a5oz7SLLIuZyeVaGnZMxnE46aaphsAhgGpN57AF5OtBzI1xp8V
xdwGr2CTxgCORqnfa4PF0CJXUrU1uZKhT5YhhrX5xskKGT0vfHGIjclG6nUwyUlbV8baKuuYOOaw
BxhqLEN/SzxPBoYIduWJ8DQFyQMH1EDmNIInJQQpOP9bO//U/RKIpTdn5I7yOxz8HNenNxVCkEPk
l0un//2tMLDjDzsMgzT6D4VEw6ArKlcILFxhOIjJ6WZlMg0WxZ8DlgNDqyG00APcmwpMkdso3Isx
x8KFEO0e6H/uJyZxfliDUYGFxibgUZotqHKg1A+sEy8jfcKM05Xs8Wr41rR2n5c8PdKpITkh+WEk
qRVsjVPzVKAthYuFS5XzKL/FXj/v5HERlZsrWY+Exp9KyYUsgerx+G1MZEmg7ShIOumdGJ8KcUvH
NkKlhsIp3WEiboR8T2CbEY8zwDbU6W5M1kHDaImCRT3sFHfPZOuB94KO+X/njM/D+ZyfzYz3XvS/
x1tojOIDgG2CmO4IkfpY9vKPjj6XM/4LwDaLT5kJzCIPSuc80uzs7W951Asi6UBDfQQv8U1WlmbV
7VeZ/sX1aFxNDg/Sjuh4fu6rdkVYGeLTLnaTuaN44v4tHel5Nn+DtqdVy7Sl0H+oFB8D4EB/YtBu
DvIDLpf4TiefaraOSOY82UUzMaU6WcSnYm1c3Y5nEqY7UzMytY3dz7UVppc7up8HjA9+RQpyy0/J
hljPzcYDllMzJyRSqPaKDGgo9mH+myOBXL+maLuGlKTdVYJz649qBRKB1VKEEF38LO6Iy/ji/tza
oJy1j88Yfj+sYsdYYxljB4ankuEWx26jcpLjsyDQNMetDuccGrL2p0qPTv0/gF3NKiZNqRcVdPBi
1088qdEQvXSiCRL4NYk91u9CM+qjnwS1ohpcltVzMp75i75nMB0TX/y8OjpoTImN+/ZIh4KxSSHy
Dv0FTBenMogDOYut3gpFOQQB6DzhYwb00d4moOEHyfaXKTTSN/AIWEiTY8EtNT4/SyBpwIi6aq02
yJen6h2p6ghf7fV7+EH7IIRcH9oPIWRSSZMloKJjuRoowTrz2t3RZkFwxaqel4ZyE/9Dg8veK+7r
yoIV8oKtOhaEj/8pBK6V69MXdIsK1g8U5APWEsmUNDv8+tqSg2W9jWAB2ltq1VwfBmPFPVZXUtkC
sGPB8fyl40J9CLMQtd/LGJ6l+yEs/r8QXHJERzi9KSTgusD4eJ85gSKgcTGbqr1pfbf+w3XbeZcS
6NsP54CdZDrk4XHzONIc03CqdvNvj/koobv58VP7LqP2ReVO391pvom0oimVFakw1dyz0ewk/b5N
bGkkIVIrHXu7lKg6yGGtdA4Y6y9yb0zicwvY3im/uBejQMVSm9bHfVqJtvrcdMoCgiPeFpYlaPX2
BM87rqh00ce6J0JKt7hnEil5fGlHxZ4gCrc+MZZPxsmLJev7ZWi4UjhTmKKUfOuARs/QGIeA++hY
DkjVqeKlJuT6WAdT47+wtmiMZ0H3+ZlZrVvM8AOP8+Hts5qJiqEyDDw+dqOSSIjVQLeu83/2PSXV
nRw1mCOChY8oLhH9E2nF/mEY5/1Ym+MPnOwfgHy+Wz4SAkLCw3+UdRfFaVEXqpn7KDI9hxzV2DTU
eODI4nMFr4KQwjLwdL0LWWSMoezdUH+46J4ANAAL4y/YUjVWclI/SzST/HpXvf0NDbsC1wGqraJP
pgDsm2neH8BsdeX6VGGxHu/tFxyfKLi7GHC+sBsttM73RodS3Q1XmZWwwoMagOm5AEhRL9i3122b
mshsN9WJFIx7aSrXZQnUooRRUU4j9QcnzAMlA9ozRUymjO2yNcsJaTPXLJev4N4uc8H6vsEEqZ6m
xGvYu8JtkJmcdOx7SdSczyW4mT/DoLNyItJurOW4DGNys55IjyiAlyk/tt7HHbyG4N5GtluqXOsO
fvqXsILpI99eEwym43O6z1fz6oYitDnGqyaQxC64BuhJn7OzL4xxmqSpex+Ph1CKSs6mxOlFtX/d
6g27h6QgCUXZMmxlRtQiseFh0BZNuoUK2lWNCVtqu8/oiEz+MXLrLGSCGF2DNiAWJp0golyMb+de
6NrtybPYz6s72VrJ6ylB5u7q/deFWiV/i0NqWKi5xEWvFbLJWrI/8qtvcmLuFjcYcmy8Me6owAsv
AqQXgytzq7b2z18If+EgDatloSh+XiPlPjWHbVb5ej7d5DJrmhoC8KpbCDDw6zaLBezBKsHe4OW7
5Y4D1z88pRUg8PfTOp6g8hViwWyWvAGroqCMr0DzUJgABwO/PC5F9ELE9U4lwaEqeJdjFzlyjWr5
1hwb+LbA2QRXnQsEPKVZhqdJRfq/uRYJtLC9QitJ4IjIMlXNjBSR21zqknB5+9NlqHIVMEcQt1gw
qI+SbZvTZqPe9jJwbMaz6mXjrXm006nNSMHr7/l/GvYZUeQUQqeuupAAmQzrAo11N+FuctL5IRal
0n/hTbW0LNO+PP50OlbGmvsgGsF2xP4ekg7nBfDB+XXEuUWQYZb0YaRlcS99F3bHJ6pNOePWVbGN
SMcMYLnCbpThAyize41NPMfsbEXxj0rVjvyEqUAvCX7Y8/S96a+e7QxUvP4sxHJwi7DIOa559LDc
diJz/GUbLNrFAlk3tsG5TQMxmrbp6pYnRznY9jzp+vXM/eNvqGCRgdu+/Ot0HrV/VxqotNFaFWcm
3yCtYPvqw6XyVn1n1yX93y+4lR2rYWBwzbwUnLMI/9n2ve+RBubcqBcB0C5XWdAhoKfsSV3hKQmN
R0dMj1QYvAaUH0ZSfU78xhSrl/xda2mYrk3UgYX/ft1qZmEGFD0xnlt/7/adL8j8fWo1WBaOJMCt
ED6QRuR4CRMhNLxe+qmFy6vD1EOcDM6jy8/mTTIqyFqAKxynu8g+38KMSSc/GstooWgNZ95hRKpS
wxGnEFUiNiILQREySKenNAO/VfufimSNo4+FxexbHEDC34eCX3hKg9zEgiZOlyImtjMmqtfxHyeL
5SlscHBLWtmPuHyYvlDcEYRxOrbT7+zuBHBgd0aMtxIhENuYCdRQ+xMw4pR5NdtBcItw03hsgRAR
uhNSnamFZEE6ifO7p1ccg9RpsZ5xo8I9JMme0C7OZHnnu0X2c9cjTafmzN1rSotvjjxrAENPQiEH
PndsgL8OYMyVzUeEWiyeq3bzcjVUfxVh+GqgbT+Fiq7R9aBW0L8kfKaMRGL+ehetp3UYG8iDHu6C
imHsrfR+tyQSOcmpqXowNhmSSxvewkPmiiihZM0RV6qiVHcD5Iz/UV0dF8xsvawZY+wrethffblm
1Sh7eN6yERVTtAEFm7W1qFh1QCZDl2ILmrpTM9iARzpAh7CuIR05BAgsICh0+SPr57xPFjusAVOA
c9WA06gzC8xcmyH7T9krWjSfJe6kUJ6VNUy3XTl4IgDe5TCoHbyNPIsiKn9wLAgL56AiqJ9c7Eyy
5EXOpbLwg6QZ8hvbBbyK5Nev0olZrOcPVD+fExBixcgY3Dx6kFWIv46jKLSaJJZ/hgDKci0Djmp5
VFYNn9ltM/uLifnVGBukbuN8sH9gS6fymEV54tkgUPaC4ScJJ7CnX8eu9/1N+iiLXeqhFuVPe4D3
WREJln2WHi3uIr57u86wGh/pAegB9zowJxqer4PS7+5UVZxXOlq0fXcbUvRN+cJygk9L5NqwMhBL
v7mkaU8c1Ec+lyW59Aiss8+Ho0jnVRhIiWx3xe+xgIHmOB7gvKgXj5eCLhRz3shm62GwyR+QlsRA
IWJbf/9tj14a4R39FsoFi4W+sFkOcrO009NDZNFd5jdVEGl3BWUXAxI2TtdMnh7Z6GYqb8DhiqM1
iJZaP0w9F+XUl7a8iQMxRkcO2UT70POGTD7NEZ302Tn+vPkevQ+YGhmOJoTHMAp5i+4bytjld8ND
paw0jHrWg5ohF/FUa+7YFArZrqsWQ3zT0wwmDRg/9AXhN6w590q9Z5dcv+NPP/xu283DrnZAMzv9
w0AxQug6MJmvv1hM21xN0UaB2XR1ZgWomdIBmkHVmitmwT9GVkeUIQ4wHPOuzkIy9kYiL6gcv7yj
MpjIvJnjbqYGQK6hXhpLhguALiB7XoXcexC2e2iUCrNQgd+6ZnNP47UR9ghzTvEriaTzSKGygbaG
j/A8H7xa60TkAzyozsuNRT6kLYMr/J/47Xh8XjwUG1MZActDlb4HL3w33JTnJa2uf7SWdMjMLgbh
fhbzaCNU83C9U0pb2/YTIOVgl13DDTFEpNocKlG7Sq1GzjZ7BQ9tQm71c5XQpXCc6H+bHxD6v6wd
/hNH7lTPvSs0cEsrxRmL4432jpyJh9uEnkJTUcIhrn13JtJD3Eiofh3SqOaNH2NtNKSYe6EHuRQr
AtE+iYSi+y9HreCy5BRGtpgxY26Kz7QHNwbf93+PsZoKWpd3EShSTYsqBwT/SYijCchtuhlxcRVd
v3A9/LZeA7HKEnzAqnzp+r7mdfBgKhR16pqG3upwu0vSZfBdytyuYVSDxxm2bchRTNw0NQURJt6L
K/Wklfo5XYfsuz2x82vKK6WARRkZDNrhndCJhB87Y4Yzc9IuiPINrlIBObqGuec+vDSfM+Rh9X0b
ax1j5YnrH/mh6bNu5gIz2HdvEaVw1xFSFIOMa1FwPh4Sru/KUC5+xnHg6gYIMESY/Q81/Ag4QBHf
3+88kAd/Q6Aw5ZNrwkg7qgTxQHFQvzM8+UFmfRpAAUwZpH/Njhz1Ss3PJwD0Z9CqL7MBt1dINSPZ
bs8zS8V+eU81g6qmUJRgU9/bhNV8659CK4VBZdvkRh91fKObxvvIWZ6CYm3hrRY0v6Mo9GBg2Uef
yv11SakBNldWoiamS9czwTzBCSIKqEfMzlaCTsduu2UQXJFJv+w1yPzSuhkV0llA3KWPDqsbHGVR
Iv482ImRqNselt/yP4YS12UAW7ajaOchRQj2Gu25MfcQU/RiMrYS+T+ZivqD4u7RUEGVEN1b956f
y6wREPGoFgdzmNHV+9o/BmHlAQdXyfJKCDuAkfkhb47uQyBHWDJLlsBxSxiw549HRvFEJaUp9gRh
TIQtVBH+Va12sn3M+OCU/7BqwIx944CSpxR5cBFB7IvYBeJcoB9r8LVXkPnoYLF8IynMMnyCb23v
dkuWltRuy1zFUae3fx4e54Tz9ZHPsCOFFU5KfhV0l9Nh84PTnwn/Rd/n5HBTXNjPcMfIXzwBhljK
nMcs4dxbOg/HFvfV6IMY6yIds9blVMFPZodAYbkC0ggiFmg5srjk8poWkRSs4xJ6A/7VZ2AwYfC/
CUYwR8PAUZb7fXvjtBCcjgM9nZ6F5ZWyXELuv5Y+W4WpZfWLRgloW+vvC9ah3eJfxr1Yw7+c9Q9H
3AAivT4VOwTd8VmEii9iusRPntyaHbZBGO+k1QUVKITgsWcCXHnQ3+fLC19PD28PKUQcm+E1zAGN
rvYaD86X+9m/7EQqVrjz9QTGbNIMkizBZQlejYkN72M1hChQNgFx1M2r4nmEWQdY+OccxZBWAPZF
2RRHtSsuy2cluAgzi04P9WsYfx5MAfIJYJyr5+QYqem0VlMHv9alcjSYa0sx4vaRFhtMcPPhzVTR
yI8HIaGdjpXp5pnDmos8sNuI+Khic0bxG7dzVzupUsurdmUnSAJuxbX0giWlWID4qI2oG+kGpeTE
9HY9QwZewsreZi0uFCwE2pxKbT5qjRzqwvCPjsavj0cj3pyA2EPB07YDxH/RRBND0U/TrDaRV2xW
fHhMH/DLJ/YnE25xWOqyNErZhe7Ub5AbMEEvmRl1+4uXyzP81VSF+wyyw/exb8dINwnPTtoM5wxL
xMEoAcqLBTTTjwJguUGRZQLnZuIRfdRBNlMbhlsC0rky2idyrm/IfKRcy4nFUe2xcBEfBRqYzhNE
AMxZMr5ZWecxzQ+gF0JjvcsQuW5yYc9KUd9XK7k2aKmfJDxlfwDpvvLd8f9DcP2gxf/iUACAKsrp
3yhppOTxXjgKi9CRLp9saZ5D4Q6TuGyKhG+mhics9mtp7k5VSWWQM7X04JeKQ0oU41J6mGuqlZfk
4yJ+MxQseN2qWWIMl1XsRi/OCG13wvLhYEny/KdOFv/55vBTsv7Z93ay4XIPiejJeGQlegDy8Kz1
K6OY4qgVOLHQ1cJRB3cke2RIsQI65sMrPNmvLL//MvOBOWzI4WIvBOBVhDEGgvq9O35TxAMxR4st
aBXNVGfiIB/h50N0svz3Cbr8ek+ibAC5AYIcokCWboqWlW9OZvpfXaJL2yVhUzGUl53VOZ92v895
BOjXT6HtoNpOt5tHGeK1VtcPDbBCYNBFy/n4pMFcGaYkblLlCY/N+J6aFzxYwBInOfbzsrRapkXl
YIfquLs/IAWI04gtSAdWzTHHU9QbTAjx9ikQKooxjht5o7mpvK49SzBT3t2xPLOF8ia+yTET0DjZ
NZY7g9CRegRbjjdeSO2yHdFtCKzjgshw37rV2TeXKxEae8A5feLWeL2is9+GdKlDuD1vwOY/Ogoc
zls9L5TGDWyL5PQXH65amvCVIb1OhALHbEkn69s6m0HCYIqm4XFQ8RkKfMO3wxb8AQ7f5rEGvNje
24F6k7txBxZ4AoUBGNJ34Ufye1ijitrExs7Qe0twvLTl9Yhrv1znz91+r+M9rHYk8bc1n8if0dsp
XM81NN5M0Da54gDlr4zPDbMfH2Ax0xkUw/K3aiRZKQU25IhL6K4mzKWJLH6VfWCHYTRglLIm9K4L
3vTs5LdTEoeHnXeRFyiVaU929xQ8wZiTZxgzOwIOKjSi+1WcdlfJd0i/XrYZXNdwOfupj65PFSDg
DG61MFubn1ebVRYCz01TRnqj17hnlRffQOD2l0I3Yio6m1TiMFdlVdqDhr/zxZXXE6OffNm2LYrG
gxcclCshs4gqDmSM6ethUJXJzJ3nq3rgAjyrDyXLf4P6axlQ1ZDMNwo6YeXYpjJ41+oAoKADGFam
FerY4YjxEcTAz0/Lo7gwwIfre016tDPInGqlKR7QZrQ/K267d+DuIbcHhjQP6V5/e3NUHD0Mp/kL
/5XSL9zUkTr0q7OmAaJkAa8W76QTn26LEFTfMrG8ozZOGStCv/GRJYsIW6PFDObNmTdgWu0dZVMF
Im/aphFpuyXoj2pjTRtirJ1BKr2x7QUTvQXQ3nDhXALs7uywvUzH2VYP2VAvQen8UYrhEDCGR/pS
UmLFAw+DGw2aC2RcN8mtdS6DaQixG/idS2BeZZtkcB05rigXOXYRjHhcRgLok6IA39geNqYPQ7wp
BdI8RU7ae7Mecrml+bGC+ANSLJ7caiCMcJ5MQJOHxluNg6NnAb+5q6L48TwgMhgsfNYwA4iXr+iF
bKhMqm9cbE1FcLccrwK/LV9z/qBiULJekcDo2eDZJJjDpNPT67XQH3OVozJNyjrwidIFnguQDVN1
atvw1nNq3woqVobRIkW/HbqIZ9pcj7UHRHf4fus+e5RfyZqNbR7np+pJC7GpR2zfv3Ipf0iTRWXs
iDcso7lGsObdWv6WHhsfPo9wnd3OMAjfNTKCuW+vIENkpo+yMMBkvzjI5pREMpEwTVjwp5vpqpos
nhwYWIKPXK1adqnTuUbcSjJk0n/qDnamCjHPGKAw86hYlfDQQpV6Kj0tyI+SUIFv30kCf/w+esIC
8/npGsox570reSUy7dJYA0TT6+aYQ0PAh0MwSz5BwCwRMYmmiBzJ1RhBu1/BS6v0NAGFHvWcR+Sq
eGxrtRGcD96blu2AvzE6qlpNc7c+MXbSVRKzm3ZApD4V6X7Ig0Jm9nxoGyc3t4tWke6JDpjd2nRg
MyNQDBDxGsBobO+yN0c5Wgx/cqw3jUmYxQaG5XYcwdXu0GJdP4Mnm0xcUzZ+jGgnlJPqxVfNrqNB
PBNoLD+xPT/FV1xt3v6xCwnvPJWJBhdJIaNEH8EwoXpoCtM2LFci80/UK22PV6xq66ON143z+HoP
mlFLnrUUscHMD4prgNqM5LkCpQcgv0rTxObzQMRS/9UAnd3JVRxc4YxkEFHLt6I2XgsJJvA3SN9P
xEbBA3hMSprUcaymmtvKy4NdMAFlMNZDdt0Vutms84z4oCS8Ki0osMlJ8Lu/WQUdkQwZqcpIGbpq
rV2aLs5nNm9qXv9Dve0qbWJUnVvn8l8hwknf+9cGpgnl2SeHplUDaXjj2WpjCAauYEGgKfWfhwuX
e0F0bxYlsz+xIaFeRzWNVsnGKzmkhMS3ReAnz9Ck87xMviMkdjgZqIm/pbWIngVv/Oqtlqsp4jfR
+w7g+YH/QO48F9M/GZy1PqHbZGqZ8Fqo7YRRrIIkaEO04Ha+VwzuG4ysS+P9HwJnR9Q6S/xoa92T
7p1LGEloO9TSDO9+h+Kqimw/Nam+6vcrFGN5cYV9wXI6kRXz93bstubwUFnMI7aK4W06h/GLwmvM
iirjti8VgGZry2IE+b2SkQ2uoc+hGXcjJRSU4FuH7FKEKU47JNyox3I9qnP17befzfti9euNg6Sc
bISTOwpSo5RJak0Axn1G2CY9vuqdjnow/TOxJDcdGg9CxK8oLvDeeQhkH+rMEq860arwaCFd6HFX
iAeZW3pdEDmxJT1f2d6qTXJuvJrOy6EcyifREDkOKs6es4NjNJT8vqyChyazLUPVo9fNHWK29J2V
EFdzVzKQu1nVaXaIx4GjAINcPr11JQefEbJNNqUfLYEzQY5+U16LiClIrEYpJ2l/lqlJqYo9T42V
WI/U3z0CaXei/fG1EdJcFmzbqsuSHGog5GFZz6XVjgCZxrTU9pv2lGB5i5t6KQILeADkavRDZHO7
xRv+KbD6nMsMkAyHzmJqYPI+WP2Mqg2AoP3s6l+mrYDYap+cZrQqtxCmPYznYUqt9xpoDw2MI17q
o8AvYWY6MXyqpkEWc6IFPveFwSqIvSzDqBsyw8yxAyQJmMwXfMB1nB3C65KEaJScfauwKGVly+nx
WLUcX4kGFCW5mc1bxDkluXHPAp+QUuxdsTQcsyP2Xc37LXZuFnKjCKKAkoe+gUS4ZmYbbQVUs8Qk
aHaqGhPWvFDBIyn/f7Pk8ST/Zv/GfTj+qa0ioRjX+VRPG47565BE2uhsj5jUC6meZb79Gcc2MInN
Zyw6d3CkQPxe31TS9RCn/X8mTANWseKzwDcJvClPbVct0MqdyA15dFHZvw1F2iUbhu6ggoXr37vi
EiWTP1EssyAcKE3XXHHwB5Z79c6IZL2C71i09FNBNfTBD+l8mxA9KX7xLBGduqYExiQckKtxK0G7
iGYtP95BtSu2z/HiEk+66qoU+gSLsQWSuoY+tpTPA5VlewTFiYDRghDCeBxtatko/7Ky/DpNoupD
s5C0+ERhiVAVkvJ9cHTVPAjAfXUo69kRATU1JyNq/YzhuCfGA+z9G4Dl0edyvk1fWlAkbHOA6w6R
Ulue69VTurJRalwv4dQE7GW898hMj4uVXU+NLawE+1hAlmvyexVknew1ny1jPrR4f6UaZHx7f24E
CuMYlK3zMEbNLzOU11hwDkZ7BY5i7bibXIQaCABonc3/1T+EM3zeVb6KPeEnl9Cvjf4w69isVcsi
oST16mC8M6XiHBFgB7MyhqW3BgR7VmL37AzlCrVU1x2ZVXfZI3sWGMf8ckTJ1PYQ7SNyezg1N0Co
MarvPr46v+b1XeTJCDIcOeVHAh1uzPRaLAklZmCChVvSnpArnCUBI6GjZuWhoyzRs5a0A3ePIztd
0pjimqQIjS1rNk5G1ZPlq3kZO91EJ9+/sZ8jfkqKP/9ZJ6nC3qthbcAfg9OIF/Y7J8NPBui3KNcn
mUkgsHXkSAGUDttlqKE9PmrgXNpaNcIM5yQqZLZsDemjCw546gjz9JlHFzMNqZIuDvKirgm1jOJL
gfOdzx+RByf5iG2lI1GU2Jae1rKAvIllkfcripg9U8Q5o+Hw8zsKghEsnltSOMLdkOnyPjM4sXh9
MEDZqiqysXPI9ONiLe/r+2+WqfNai3wjmtJrODfBAGyYTwZsEKSggYFBhvSd0RSqL6RUxO+XEAa9
YR2XjDtyKyfKuteG0cXjsFQoRQOa1Vmlu3wy+5jZCXg5kd/9AV6dtnHtZicJrh3I1nnChoNxQWX4
oqQ2RdGDDBx8VAYRGiRyQoAn8fshIbBcHZFBqi1TQtcAIPX/Tyh7iKfhYxCSCLXtmMuCjftoZQVh
Z56HvOICYQh509+V87ke4twpbo2AUIMlO8duQObWHTbI0t1WGu2wVLebyLAjSBs+35GnCHJxn4uJ
1H50flOHVRVcGvQA0Eob6i1TJn2vH5ErPLx1K8OHw8V10fT3jKzKIvnBIIrLaTrNY3l42y1a7qW0
DKfRBPff5MKutQj2xAmh8qcyH1zA8K9y20MJelhRZuBGvkZNgr+O8YnUjZ3GwUijssc2Vww1vHW8
wMOHNzGql1STWZLscgf/ZRAC57XECVO3YyWDpYJzkYTY07TN4rzAytwIG0Bg1KlvvmXRXfpetGis
g7OmXfqOpAanCFY9Wxl9iRp0RmoZ6L/uMg5pReB8nhmv1B1xlrWugRQgGxDDkm3sFlaV/NXNGPNW
Oiz7C0T7vOvlRXOjTEMXupjc4wM15QLqd8OyUS+VGBHtmjs3C0xkmqsEzjeqQMCRolIaC9xYR7om
ERIGldsfO0hwgA803DpDkAKsRIe921lLScx1TIv6gj3Ain6Vj/f/ZdNI/apOjDHfGXxxWmfza8aA
ui7EYkcXlJyFvRKHPaET9HOxKDDm+tt+PrZy35l9nCdvKLGm9VaulU4LTIuKX3v4M1X0I+ob8SPp
bLQTj2N9cGEPYMKpnhM6k5st1ambqD9s/Ml0sIAC9KAcuMaT5R+eZBRhMgt+bvB6hOh1jA7wXYxg
DY1d6zc0aK07FqeAroKzlm2nLlIJHXPe3nIrVfByTMGwecTc+5BVNVCmW45kZhbfkTgAAurDXx5L
gIQerbd5Y/EZco0PBztVE8SK9QA4CjO/TqXwDjXXJyS8pavNwNCo6JcTndthixoz1q23T7zS9jbP
73ZRI/zfPZBbiHAx+HkjuXZRG8k1Xvy15MJZR7YOCEGFYf/kDyMKARVKZcHLyb1EH72GlqCr+i8u
nWxIKL1zKxdRozT/0eNVKaYDSc9Lz6cDf/+evLiLOP4ZLlmDQvQAPj5efqaNeAS3hFx/01J7xWCk
VeaXs1/MH/m0rKKichOjzxZWTu9qrZuyzeJre4hjWcC751rRZ9KH4FFmiNMBmhR9Ofbs6wBmLmTm
hOVWK9cqWaQv0qL7RxTbxoOuKWjPBhR3a89BelpIy29jLRM4txFqXqKKgmo1xaNyrkesgXzr8pEx
RManBSeIAMUfj9HItSz0JfpDgwEkYoFa34QFE5orj4YJP+J91HDEuITmSInyHR7vLqDKWLFEtDdU
KYmfTaT2UhbG5tqB0QCBHyjH6IK2P9LvJz7/J7105SWJHnmh5GL7TIMP1J6K90yM7VSlPP5scFLo
AphOoEcydZbKtM41poM7v7Lap/sGgLWxpYzs9AVW34gXSPBP11sI9P5Z7blGqmIVqXx6HFsUfo92
igeBJkQkm2rVZ73NEkSC2Pc9YUZmEQ2IVBjbU5ZW5yE3nMysWadzSCDUOMCHSzNcBzkAn+nVrNOA
Zi3KfySeAQbHJYhuk9GgLdQEpw3Q28zLFIgYp/19NHn9IY/O4nNm4HJ/X4ApM+QfONJrRPjT3iIJ
Da2IrD2jW4p4kJ6HHs8DzGX/0dngnKaA+C68v8Q0q/ysLAsfuLCGoknrYKQeb660zoRCtQSIp8MN
VioaHtvxbLoTUqQdax6gW5C8GrJMedOuaq5eh1x5MnYcAsdZi37oy4MLWuSLoeSAbCIzs3IJXJHq
DAsfybYTvmorgut6mvtE+ELSqLuEmu2X6BdIVyqbiRpUKQcJViKOnCEoEH/6xgBF5MkbikKe9qqq
/BaQom0MCrYlVhCbgQJQjtbu0WDjlO48Luu80rpx/DbeBVGKUPNq8/am4UpovCxb213qqB/hTf3o
sHrKJijXXOHizBP3a0yo3LG36zS1pd9Z2Q+1zmduJH8GQ5/z09lze2EsYzVuJDsBp/xaN0/U1Y5u
C4x2nnKlYypdZZ8ehjx8bFSvWd+v8MosAm9kMm+VPi9Mt0XDQu0B3ZgMonRt15XIjMJm9ERLf5bQ
VX9vdYlGD1PwwjR+0MtR1z+9HuagHyaM4U7EQ9pesdPmtslZTqHjblvLh0mmIgajlxK1LY6EaU0c
ZI6ashSELdzFXrZVZMNjSyqtFiYfAMTsO9m4sIs54ArdJta6o1/D3suiqyy0g2GjJeOsabrc/MKh
xppTTgmiF5w36T/qZhqgmcwS7otpAYtPlYCkma/plRo2GciI/pXBlXyjK2kbcAUCz87IQFNsaWPa
Oxw0AUCwPFXNdlMf3zfkRhMalzEioMIBPGqwzXFgPVRR7IkqrKtMqM/rgd+rH3LPY5aXDJ+ZoDAk
JBDXatiF7LhVjqfWMQ4pGwdDw8nX48QYUJ+tf/1rtyU77boa1SKivGj8lo5oxzd2U8dTmCdG3Sej
mayshzqyBp/X+JfzpoxHvid3uRzS/gLaryLCgNT0hnFW6ZtdCHs4q33diqJhv8zL5v5L9uzT07qO
751QlVtTaktkqGqDk3QIPhzyEZLZHmqiVklBhgszg1VxcZnaewMWpl536zgCn8BpiNpwxVXd8b9q
fIqhhPDzXXhJ5355eAe8wL62Tk3ABsIK3yqpa2Gz99PQO7S2umgFXxIxpRcewdcoGzbVXc2hQrNy
t2lYJclSi54//n3PJV5Hh8pM34sJYhLtMYky0hAgTebl4yXuk3hxoOrvb2RePhyP05fuVmGgOkuC
S9Z37FtXrnMvNiMRS1eZaFL4Eg9Sp0NRk7k7jr8DgqUy/VBOdkgauR5bcHEkuhvlylF9/3ZPrlEX
IcLVTQaYg2phTwRLgDTCuRjuLrrBAdiAWEJWvqQm32Vm6AKYPxd4oo9Uz2Ysj3KNQW71nmYsUhvJ
HiC9PYnuMk920a903HgT68Ipsy1PsynSzpuvuUgEqnX549cvi/ZBrBaHRKgZ2z2skWNGDKZHla1A
OAQBRzo7Z7viHWYLur9gQZQPdpJVZRdw0rf6kxDdiRKywC+8LwIWkFTQgHm7DgRFFIa2vl/OkweS
ynYH90QCKELzzRM7d5CTy2gIJKvEFkm4vIMIK9DvCTFJewr7+I1JN3RFKqvn71LJxDH83kUBH3/l
DLYGdHWpDgE1LjOrYOl3ZWVuL6PknIG/VCLElV2QktQziYZvUe0Ay9I54rXL4pCgls1nm5E8Gfel
SC8m1UvC9PeZCgmAz9WW1YfObwbNeqZ1VDeNexZF41bHF8guluiHqjApMDv6qBEIqLozHiKgbRjc
JXpcaRmT5QHhjOJHddUyhuZZ/Gn/gaF3lN1SzVZHcLAe2VE5WSz2VugEDKbJLApcaY95CEqAaCgB
iQF2xoqCuYWj0Ispa/XIVEoqgUmvRQ+l21rT/uJUwYGDAPWQwlH6kZMWt4pf2245dS1kMPIkRbhy
GdDrVNzdjDRH1Bksv6IcEq5eQqB4zN06iVahjjk9xpk8KFonZpvcWGoVqyi/gl2pdwMs/kL3gPj8
f0D92gJO7XOibIV/E1T/bgYLDweLsy6Ypf3eC7hHW8n1VbCdEVVYki4w4+N7SnfR0Y0NO+sdiceJ
sJxj9bzCb2t4/gkayuwqmlg4EC/nT3ZCQmS9TV0770Ouad+KjHoqq0d+zzuHxig2t33bOo/ElYhV
7q8SeRhJ2CUjeFKCYtnf61icrSvrOoOSFeeJL/sFIHhn5z6qvT8Hg6Gc6rirgryw8iysUYAE/RSq
Gk73EwPqI1Fw7d8mTIAtvFmLlG0MhmZh90Rsi4yaYHM/g5AkNXyi7316CJexjFJjq7ZiY35ggjTg
2DXe6tva9GnVq9BW3CMCKkNMnhzTpDSn0SREkszySLoGpToyQPWV+9x7A/8BQ3XOVErMBsEzyaEm
a7Y1A/bkAwqxlsnE2NBv1UzL/jKvVphmc+0iQ5XuVRV1xk57SDS3FOpv0mq79VatbFqoXEONB+v8
c5/TUtwQA1yclzLn9CPtKgzcFBvFMNKCjQx50VJzMCgXhQ0ZAVXAs3ECqw4l4elDHWU/SslV+FKa
ckANFBHglxRAA2sH85V4A4hXNWT5C8UXcOkD3q0urGNJrbNsVIn0LtTe5Pto3SckHmYPXwR0nZVD
dfkaw74qLNuqMoQ7FgTAvTUw3xN5w84K12HP+U6byoec1kfYxvND9IyHTA2CVnyN01xFWZ5hTVnx
LNbCx/k9n1es7Se6Wa8LH1SANIhd5ulu0ovV01FUEQ2MbMqD8oFvIQZ2IpSz65ge6WBAnqkDVboM
cP1Qt8mDU1VoqsNXxEHHdn52Fy/JwjZTGVRCBZEgX2LmeOr+ctQ4sgrZXbRVR4+s7uu6Y33x9rQG
ll+q/KbbExTsoj7LlD3pseVbxbbJqGVPnxy6frYeFZZSxqYTdaHA+pujn3jbs90KhYrbhlg5jinz
308IXHxYPjdz4i4PXVcVPLdkraKj8Hza5xGNPbGu7Ix+/w5nPtyD2zKOtvkC2Ghs8+hu3+Kp8NVg
ch1wjUFJRXMhpshwwYdzlF5I/9wgNh6IOxAzPXnSu4WBUjajLmMKLEwplcgQxQ81Ez2+TbZxqRi6
szAK7sPwjvUe7BeJGGYZq0eruB/0EU1rL98j34AWrHh6IjZmirdpiODxTqv26EFYKe2E9AsUgMFI
NXVPSc2fau+NBmsfFRL6LeXDLDAg2gaClPPAjV/BVf9Tectb9X3JxiA052Oz8W4Z2+O8+HpBxoqp
mV4I6sQOMdzDZXTaUf+yhinlHzvfBy2asTzHw9PCNfmv6y5gKswjf328YP8LlilBpHNK9wJkkPRO
mGZxc+JLBKgOnm9hHLKU8DihcP/7arcLUcRtZBYD+MvZnp3vKQO1p+i3/XYJE7vgtsWfsvBlFw4n
+OYhDU3Gh6UvzSD3mFCjUFfnH7VK6I0S6DGMecY/IJ62FTrgF9Mhe0ES0yxNfdJtoS9Vv7hFFvV8
VnV6rCZ4nAb5xHQhMGtCfR44WT3jk16KvPNGhoESfCxCFYVYiOWqt2FPnMW8F4iZMm6jC3HejdS5
TyleENOVQVsz8BF/iMyiFRKku+Ca3CHG+5U2nmVkq2EEni8A4WshcwEFbugIXeLtU779xnqkwhL5
1IlqqbgHkVPe86lCAHqxzgQdKacz0iIJEJgweRPEem5z3ceUCwxq162Cnz0rqAZjl8MZWlIDYnUI
y0bP8xKYGrUXpzQE8syCLe8AFmtNwTWiSTNecPMEnJc5PcG6usAIV3auLBL7lgw3PR9itRVDKZqG
e1Zss6hz7xDgozCK2zRVWp6S0dHlUiZ3qQgjhfq40611B4yNmWv4LxrPYtfOhwmIwDFl127VHPn1
BVk/L20VbDtbgUHGCGDnjCB5vGDBEsztFL7rvoTO4RoZm3okrK7RjdGm/U7fQ6fdlOl91wEOFJ+6
p82qxY6vDgh0xU6I22L7a9BSA9MeoILOz5hS3TQl+gPhVPk7vyuR3lljTmwnHOUYZQuBsXtm4vTd
nipA6yKyYtrQXwqZcNrkv4nhiUXf0ZRPPJUPwM07AI5W9QLuZOlKyAMGfyPHf1DpzQX1GtbUMa9N
eYoIa89teMe/Q1lHI7oyeqf08SS7MV+QCguvbsn2BBFIycWTkBZsSBECzqUZdJpdWBu0A2vGXqX3
sn7got7bSnxcMlXX7pQqoYSn0bp8KncJaaxneNmKKVbshMS1DRuOT/hvO+vgJAsPPboZKAC0j6H1
JZY7RFRU2aSeWq89aMjTgam7us2g/uM48oEm+H0u9UeVqhuZHSgjAlyJYEMIohg+ATrENi5kGp6d
KwGmbxm6jOnf74ObhTvTW8c0mWuGYKiF/IuASnT6SVj1H6Y5kyyele9VLK5wfrZtSu1za4L6AmsT
xB2BCGp+pU+SsILWxN1DyYEe4/jeVBSe8dnmT8RrFxdpvgIDFLyhxpJKIp9L0zvlT7bXpQbjwCD0
BzGSwTDdB4sAPE+z0H9EzjdTSTV/hrl6Oe6NMQ3JWp6FWR/tJfx626QGr+BXfKnicpdyaxiNBEVV
e2JROUw4OisE3uPPD+CpgBr4Lk+FGY43C+wW5UtbpFWeZIZpNhVxNR3d88IlzCVQzZjKHlHZLzIz
VLY8sA3gND1j8sxnt/yqeieCIQEhhaz57JnO+OGirteuUS81M3boR5aAGu8EyPjcvDUCa1kso4BX
GZptxkslIx9s9p5x5s7xNjACswvdfJg6zA8bl/bgKeKEwN3n7j85B2FBYx7vja4G0d2JjorjXqcf
zChXPBz5Z8rlCaQPDL15IJp2RZ5dUXVnuuoS6HwX82K4WR6tmyHdlTGdtQa1nAQ9ci3ohYTrc2+j
VdeY/1FocSSyKD008oC0vo0UOMBAwKaJ+2BZF9omnQHlYWN9YzJuaNmmAHW81Ys2iToizHHNl9bN
mg3GQOmb3/IWbM0umil06sZ1oGyK60IZ3R9shqsMM8kJT0w1wpQOAMGNk0U1wLXpOA0rtava4hL9
gu1CzyEK6ABXKo/daMagRvNYBErVceR487Ya6Aykq7EbuBhbGyJ+xXMOL4ad7QVb0jrXfo6ta/T1
f3mQAbFL/sS6zNNFwpsxSltr6xmt7Bm9CQNe3m9wh3/mADcl6RF70Bh5z4E+4O9D0Zv/7BU8EcSk
p3BHuwEXSjphtCGM4a9+TW6KgoskVM1D0AcSVmjkjLyq9rYykU4O33kKy9QOys5EEzFGSrT6SEDU
OPcxeYc3T7XDxzt8/hsQl92ycGcBfIA1Hc3qFvOHy5Lu2tt0GZIatDIBAo8tr/Ex7rSqDfCqp7P/
HYO2qI3neo0l9FfBev96lOtSoUDxpF8dX0FF+bbHXsMRoeR5kaOCPvCNJy0HY1LtzJEtHoK5Zdj6
o5kdTUgssWRtZLD/RJitGWccVYcoxMjV+28Wqtc+uXqxi1Innm7J5Cag4pSkw0JCd1Rg/3AbFNnE
SYdeWELx/Lzqjp3+t+t+jfEtXz5BTUGrhfzOTC0Z7YRbApLowTzf1CuRbaBZFH3Sf7h5TD/tQAaE
KWpddNqxspXwav8vfrMvbxSuSS/WoHRrhO7sXtrpHXz7wcRHU234iUsNku2HDhrXfM3w50oel+Az
PrVrtzdbwQBaAjcGeCVXY46Ywl/nLSi7SV9bJvX+kHHQRte+eSVsR7fQ0jk6popFm7IDW4H7u3JO
9PRHE+/fEFLbCsxF8kFYMgSFfGA8bIkCxja/9EBHq0XWfBwIJrg6/DjZ4UlG4LO7DLsVpzfQ8gLP
Md/mrkAmZIL+ACLyMunFUg3KJdEeTrP7OAaaHHQ4Kr8bxamNAfPsT+iE6o/o9bW3mBkBI6EkYdkA
yX4730G6326NItQkqE2oAsqa9Vb5C5VjWRW+zv0oKdRdUTxRnJ3plD1QzPPrwUY9W9QSR6gfctNT
9WMCdeFADfykiQIb8xYwDP6C2lXTkHFnkqtw2SRkJFrU3djnHpxjZoRHE/zfC/25Tss2H1qagp+d
Z0TnX8WxzceBkTOxK5bFl0kWxfljjc+CPd77RyNV6bhl32B9IDpt0/G2dX1/zYCao+o1WUnSRSgA
sSAlGwCxVKDN90VVTuIbg0VpReqolU7jK5jUzQX95c3pSvhd2liqJzsfWVHH2TGXTQPkczwrELwc
sEyMPLJAsQWx1NFko63uaw+chD/yXyeY3XdDWZ0FA7cLCkUgWqCpMRwx80X2ldq0fOLz19ViPScG
loqcNOfvBvO74fXeKYQfzsDSgUsb9ZOziKfrTSPqrpy5xxBpUQAh70kYHMPNcpGvfiIxY+4nVifc
5AI2X50zOk0EH1h0Y+IC/Q4HpnnHeaTvD4kks7pQxn3BlYI3pfWa3HHAikYgj1gVR4NvVvoBywWx
L3Lm9TwPRSGG1RHB9FKRjYFugOfhv2H4dOBqxCflXyc3+EMu+fRqQMsJ9v95iyFnjbgchNLa+ZCY
QLH80VSkWlNbRf7sdKYqX8744aa9bfaeh/3ljMwCt1oGnKfPwYJh+OSBYdRrQaKKzmB1dTcw6arW
MjahKhxuJNuTSFPu7ym4fx62MsBaYeJk0xPtgsVx9SCd4xtoPMS2NyrqZE7pOsHIDt6v4JAaq2yV
H6VScQyibTCi5PFGwZAx3sPFMYdoy/ZuProIrHOlz04cd4bwSWeSkAUJbpsmPK4HQR6ZEYSo/APx
uGwH4JXcNOlQDfgKvMyQvO3460NmjxdR146xChK/35LtbpIr9ojSG80EX9ptgN/Ou05uUFVNYEJy
cZXzaIsB9JT/lVXfBBLvZjNQpW2MgDlI5UAs1U1htkUpni7ACf3JO6WK1P/tbigM+HSnonSjCB3k
P1qnv8F240Hv5uDJCr9c7a+6ezGLm6YgCzNmHSrp1PTFjwFGp0pNmBImTPJ+yuF0Qk698cz6pU/B
lHImSbYfDqmBoKNDJUTjDUFRXl1F10VgS1WHsIi909FkNwpb65y8RMtvXqr0wz/h69DbvnG7O0rC
m5vNkC9TG1kHZB3U4z9JbNQw7Lf60c4sRqrBD9C+4y2RzDsf2rZRkTu9+q3eamoMLVxxY75xjdXX
GPsG03aNQr1s8pUls9kElrwL0JTzUkDjuua/CQ8MuGjRKjRtPkOrSdkW1V9AD/4uatAvrdY6PPlk
4wZqE+Dyo6tlmH3Ry5GWXaL5AAwhunSdouPJ3AvUVtv/3chihibU/dJcZf79kynOCBs7PU97NyQj
3f6AbV93OCHOdZwuhHtKdmAfvWwMI1nXjwSmY2gwV+ywr+eBoDg1Re2morM7ec4srPMdXuYNONID
NBbH/Ojph0HmSICX8NyJ82Qc+MxQLY3nyKB/sDAdzH0yNerA0tvD0B7JU7h3j4MWdsH5TKU5pJ2f
/8hplGOSuvcoIpGxXsCvwz5cKwpuQldnFB+yD4Q4Y+kU78HEESkVnP6cVFWAksVrXAeb8KNId3Mv
kF9EtSmtZ2h/HlxOlcAhdEgx9WfB8pgxxMIspCne3tfps6d5Ro0tGBUSLfn/8Cot7IzWsgH4oEvq
ggSAPuw4tfLNczV1OjlFvUrXEeSznHULLHS6P3NqQfn75JanprM4NsLoN3Lc+4WcWig+Itqu53WC
j1JSqbjFcadVIVCxyVzRrYtR/MbURJlA/6ZuEErUyeDMkx3j+h8RQp9f47shqHpmmGAG1ed9koow
3CxiM26CJceJBkpjH/cX67oCSEuTtDa52kjUEDyXsKSInpQwezUsu0e1Xl3xmiXGwqmPwiyyfoyi
CKwvY3FxRYyg+5ikGxVmgPK6FqeDaIC3+pTsJC+zEKVp5a5Ly/M6jcX05GPZ3gqrxehlIUIVKDHS
ruXPzwTMbZ45Iy7lAyo3RRfihUENdkn/fKoGNxIi2pONRY2TTLqiBPRiANMJiEncmlM7MrBaHgon
2eR9Vr4xV/GRQvPbiJ7b+ND1mi/QPictQZ6iupIWCE5/oWdn73b/jPx2M/Ixy+dF19fjdEMRo3Uj
eNZYrZjwqh/tKFkbGjwAxhho8DSEnDTLEc929uLVxdizQrb6bt7OJKe59ActuvX9tv1b+xB5s04Y
+F7smUvrrLW691mrNK14cVgB36Fq6+nOnBp1V+RB+tSbXzKVx4etl6uajsGEnQbdU4gJXDHEs6GW
a4smyhMkQaLilHy47D8OlYdHkcO1kTd6FVYf6aP0LOCpovTXY/h6NbTc+t5CMvutJvQ9xujXIxWs
OvM933goIl5ZZJDWpzqPdOHXLmFKhC9sX9q/QS0+Qaht1TBpOQnq4o5lU20EkikwTmrHtA2RThMv
7sjgadMH5qXMNBJBEjcEhzE7v0ciCPqB65yj50PZh43jYm1WdFTNIhbpdBTK75j9jCCLIb1y9gZJ
bl907gc+JZkcvfXokXGqDhcJOnvCiyn4eIUqKZfN51hT55XlpST/EyfFP4zsjUlrWoLO67qlXPaf
eje2qOYuGKxZMZLIGDwLGkRjZW81aJtBV+Q18umdu623CeCh9fOfrSLckq3LkFsz8Cte3y1wIb18
Xqi4YLNy2hn1gt/dnRSYkcE4ZAlp01JmN7E2WnsnxN5XbQ4va1Dmoe4Q8GEXNehji1zzdKqaxXSG
diSfzQh01T2NN1bgVbZij5pQcA08pUITauBNhban7rJhxUl1xbNhySYjvaSpnYthhkC3fIGas2MT
78WSs7Os1jKfb4B3CpkrvR6eAYDQ3R/RMU80XMJ/CH2pl4i4gV0pM9XNRmKh/j8u+onMwV5xQlzq
WzmxeUDb4i/yP2ZZQqK7w+g34YNUgQ3wJOjBGM3vg8nbo4Ipgawz3DefccBHmyXi1bStrhmDpu4/
QNWp2Es2h20LcqECHLEbQwlYxZXC4FPjvYMUCCSNNd4LH/MZYc0F9Y2nxHFHldAaLUcgJv+qPzYB
TJZEIwmslKKSVhlSU7gJQRWQbh/QMHzWlgpOHGxWLybvAcz18AxBQtAVvjFMq9MNUhzKUYTM7/4o
w+mczanCOWiM68kVG8luRgXoBrjfjWQl8ff+pnJ2XpVWDmKeMFbKcDkd1YBIHlvfsJ4EV+x0+WfD
2XCBkENCMJUL/Y08V0tc2C0gKVLsLzsC+cC1TdhBgAKKAVkTDge/XWPKMXcwBqygtvGIVCS1uBCX
Z5eqdzT/bMp3jm9UQJYj0EihE5hE1lzQ9WfC6WiU37kxCjOe99oXNE+41X6qc//UpXW8FvRUeQ3G
OflISzP8ETGtdx8Yzn8eIqahUEIYXWKt8UsL/foIZJFWYcOBVRVmJ0/f/g9EwsuDPEKQgUsh8WiJ
8sBCYkIKTBDb5UKllMfvB9mSjXMBKZG62SSwSi6Lj8Rbk2enciEjXZvX6w2TRvr0yR9Vj0QC36ki
J3ZnoTy5bHXOsN2y9jnOmX2r/X+7o0ERPbS0tleNE/2ouXaAi1W1WSdrlPvGQE/aM4eqtlUZMWA+
vCTTB1emR0+UgVp5eBmTFQoT3BnkwwjH7eC0lzM4sPtkXENHb7AD2eQySnl+Tywtl92izINFjKJi
zxLYV1iSEYrthpzjusqVsKbvjgKtErZY6oNzZMseael19HOpIu5M5TK3FpGhVaOl84NDuzvpw3Ki
91onjKJ7YC6C8nXqS/5EDSa7WS0BOt+py6/AmqS85iuMr8Vfsk6GmOGScwzu0hNnoYTg28CHfI4V
rnkqooBaySd5n+j1dihfO1CmETq3DIw3NF+gHb/q/D/Y5NPgWv/88z8Gq+1k1uW0bIATtKf/N5T4
m9xKl3T7RiRzI5JXm4kj2dwJFGfH0aOetg4EiaL7y4Bi2p0l8PmOAscU2f/1bS/q99RlMXVHrr7c
+LbubkYJ69hjYfOu8Jyb46NFyQJ636B5A53LJTnRBnZjiCiqzqUB8tqLxhXlxVBHGJDMUjRB3afU
ysBrWMzCl7NXih7JEfSyeYbz2BXUdn/NkDY4vzM1YXZcS4HcmKUUOqGvl+wXXBM+hHMbb4DxJeaQ
6xpza56A+UxIOwzq0T6TeW1Ayw0LI1aqY75AkRaPXETLbpUuqDt/L+igYb9utBtqMu0J5bhgbBFH
Tf8tMkXwDfGfVsISQ76mBcMzfPAnqQZFIbiDQmu+0kiQtNPHCV2LAF+zChikqWwcgL7meutzWkbp
hjOqGzzrcgmFCeJ2OeFnCmaWXeSQaQzYpTaTy4ZHkRfAib2x+7Hbpb/bW8hBVJbhOC1pVPjWoJBV
qIj6vq46MlojrlhJlFSa20ske7WWP7ycaheirzJJORq6Hl6SqqwvdibCCRdgyDTK5IdBsy01qvzT
SNFBhRRInWHIFB+8LU18Fp6drhYcqHNgiWd4YjxqoN0mwJ6e1WztH/fGInjgj7leneCpXsV14zPl
1F9A9mg7GHOYg6R0YrlVHnYBxuu9siUbv2AxCGAqNuSzWGVukimqru4U0qw3YwZPKWfJGvJODl9R
LHXeGkU8C4ZAKiy219D8yH8Ss9f3aDnfonkWZEtkM6POpEzNLmmyEJ04SI86+CL08X4Z0kCxnxqN
yx6WhepteQGiQqxRansc7FgNuLWzfBqB3ezQE3GjV+ySHKQzH71EhFdgvoRZ+ytw70pQZkPlFel6
BwEGhTu2VDaMvLfZdOS3zKWAKTP5z15V7gGHs6L+IZltO/1brE0vqp/S9CadH0z+SDI78wm26S6p
QDLLpnqcQWzQP2Ce6tpyVH/h4zgQBXnur9CtvIEmvYCq3B4Ve86qh3qXQJF+l1YzfGDCF0weC2oc
eyK8KR/knftAenPMkc6ERJo/kk/2fnNpFCbfgET9i3oPOKoZ/CyQdGFAsjNRZVjjn4bOsmSfUgZ1
wXeQyKE3u9QfdffeCAxBC7Ns67i3gwPIsNNaQ1Kfllz/w9VvJHv1nlJho1C9Tpq18uaPulp2nRJv
D2mB5wn8c0iph3PLEVH7cEWUfCG1Wpk/0geY92o25TX+8g6nBNEV7k3Ip7Zci6ZWPDd8/Ku5brl6
paewby0HHnzXxvXdhjApBSLK1EH3i4fJ1otSSxiZO/RKHCbnTUTeMkXsRNmzcE9UkQHEbaQH+wkm
lQsW5J/PHroxUzSy0YoHraz/I2DwGNcKtr7jn7n+OcWSrimtMek0zcdsMFFArdIHNLXlRUMbMZ7Q
eGJq7C4ByuxKS8tAj/6a5OTam9VfTRrN5OVcHd7JaSGY9ozQR3eVbOrSm0ZB3Vr7FbU7WrY2l4uP
8BgcGnpQoyKAEqdL92CzYL9aXzOpoCsfhxO869NiCfy4cpotHRAAoLAn1sFWFQ3UxRurt4Kz6d9N
K9Q2fNpths44nFK1ksamqOpiPq238lPNjVXaptLMDrRPJoDwPLViqxhF4LxJ0UFdKzBfnMOjVmMb
o7BlftGou6s2rCQkmHAkmeSCPW6Yfw1hjdZ/1Yl7TgrilIyX0lG4g8ao7MzcfhghFyKidu37GCi3
1aEw6G3tvOLFExnIH3ZBEug7jZvxrxwPVRn+v4emQtOHRGqb0AZP0bCRNCeZpxGG7rIdLOqaeuRb
oX6JDTpItag4Y8MZMuFNZc7aLuwTM8wVUfdqRrX+6YcwnaccQnuMiZ4vsl6hptMEvwAq8USeGk7F
/VvmmrPBHlDi77g8DeuvkTLuCp8ATb3owUKz41UWzmyVucIVxet7B101Ha8Z44ec5AyvGeIGjHV7
ktndlPtqI5u4VUJBze4b5X6tV2b/G3gRaiKqIdE7UbbsS5WZLwoIpIeXNtYyrw1NUEundqZu12jr
zg21SLBrbcmeOjGhytQo6IfLMZljpzyZpeAr4TwGP1EcKrZQKkZ3XA1f5onhw68Jqixm8WhlUhU5
ik5EPPCvrFd4dl+wjWWzdF9Z2ieqaey/kIXaDzn0wILtgzNGRWJ9Jq8KIpmHyQefnjssbFzbWx2+
JVbZ3R1nD8E5DdK0Jv+VqK82ExiY2B0gI+8UBBgZ3maXupLXEfxFSbFLlysBKCybV30h/UBn08Q7
RPLufY6j1HETSCEmFOe07qmpCyMLgZQKi2El8Ttix7lgvV9tJwKTs+GTx6xCjU0BGtueo+SPaPLY
+lntLxTHg00TQeIfAKQGblME4ZhEKAKG8+0nMFTB7sJfUcwEBRosNsdKVZtuALrNoM6OGiFKspNb
nFDmdUdNbZZTdfEU+t3aQvTT6QwvZk6wPzKSmaf6Rq9/kztmHh/FwUrGYfyPEX7Jh+MBGvIwKmoh
BpTHMidOQfT8/3O7ABx5hID5mLqHcV41ZM+FjC8Z6CFkqUMZsYimygO19qrduYVN62xv+PFNlPr4
ZAPHq51ByCXhdZbWdAfY7B+W6Z9gMzA8HuTnLCA78SPrgAuPthjYoWbhE4qdZpU0BwIEssxPaP/D
ohobtWIPmKg/Wl/nfd28kD2p+L2Vlkr5XK1iLMMvecxZun1MvVgO0zh0nQzfNK1IZcFyT4vHZccZ
AaSTTZRARtsBRtyE01dqdv9Tefwd5dSb0NFTCDq7eAxAAMpXoKg1dBa2MH8HxMr4GlN2/OlUnWLG
yjE1bLu+D20z0O9GrRtpS5HOxwtTleLdnOpnSTx+kUkz8H07LsFSV9l5WVBznmdvUtPeO3EA85I4
qHEJX76Y+p9Y9lkLr5ObdzZLZsll0+8iyF9sa9d/D6Va8YwgUv7pz4RZw22RQv6qnKQK0+fZR0BZ
2NDpSIcZNj0NsFBVhteTIYj4j4sWOtV0t1Ft/lEiy99japs8Q5uENmtilhmIV8RQqVSdLb2RsogH
2Zqslp7+1PP9ePt9e+sv0NykUOz1mjl+vtYsjzvM031dEQVtZyRVrsD3EUAEvkPCUAgMwTiy9F42
I1IqHBo9khzxH+bMu0SwEXDXSkyQHiCOLwDB9uE96zetM7eY1L1w4yJsZz9zH8pSX6fcW0LuouIF
rIuIQkrY2TEKf8HfFm30AVUBNLBe+cMYXwha9SHn60nWYA6nXUhtPmIFj16zLm49tMXiPpZ4AwWB
lTLKomi6ZMdntITFIEsJ61Nzj5bXDGtDGdeN1GWIQMElVrRQMZXbHEMEocFDheajxKLEoYoiPub6
uFzYlBvp8H9u092hYmvfWDqIG7qHy4pH02Kp/jWzjPiEKJWzPx4FgW9dJRhkY6XnKvOYGchOQUPH
ueLX5OC0oXFWEfOBaEXKtZxHX2PxbixmRdoeEVS/JvajIU1AC2zr2DweP+TN2+SWNKC2hkWyZrJs
jb7WU314RFzMFqAN11ZBuixCpaal957rauvsWaqhqHyVF+QbT8kgCk54akwNrVIAA0pHa8kQ+7J2
pgMzidDKfxXU1D/mdVgLU4UEQDvz2aOZ255fIrpkDcccOuiCqCfOnXxcEsgB0OfKETv76jvcE9LD
+fbaaZ7afUA+yJS6W6Mmc+CGBth1voJ2Qfwf2wyBmvhjjxZsxSTbQ8qnxeVm2qM+vQwePpjPzis8
4fXmQLIXqye4TguulcR6RRpsDdveL6Dbv0kSJkc7+egHvgCneoIuGX+SZwg+LiKf2cHBjwe5ohZK
QVmWlZwhocysTEbmDAu+JLTgfLIY3ZnCdIGqauHqwltePzHuFG5xuwrkXVPg7rbMFzkPRIE7ntWv
buymU+7m3x+Pu1M+41mb2g1JfH7KMg1ZFA3wRYz1HETilwzathNtjkQIqveZh4EhxK7k1ldANYh7
kKkGptvivQPxffMaOdf7bhagTn2Jo8hBfvqVgNwbTvuYtWTk9XFuQB/lV1NI4f5ZUNh+XChHabMK
1Jbf63JdBal/fvWt6f94UfWOc2fR9Jsf3vWmNQMA66+mF8mIA/D4nT7A8O0LKDxB6yUFkAO8Y6t1
bjENOkHaYS9ZMtq97bD89xIhJvuC50IeaIXPdMyaGdg8rOEYfiFE+7lZ1VO3VHfKNjPI7xvy2Swk
GEOqdyHN8Tl5FAeolnO1qtvmPo2M5r37MUb1guLCo6t2KpgIvAb5a3bfTOqyvDoQFFHTXo8NEUsl
omJdO3wX+vMvsd4IDxI1MNXoDKO3qQXiOw1dOhRNMkDq9iNyH3fQpEy0AQHaANh+FjuMHBo7NP0b
2ASt1OoLOzdy5hf3zBTZRPu01cQOuovKGKSPoJDSDaFU1C4NgtVyIt0AiD4oJ6T5L+sDNay6vag9
0wuLbn0AHhqrOb7037wZ3VWgvHDsh9Hmg3ok+/qXcPqLiUthJw95HFJ7aTx4hY8nACl4AkuOfttR
Zde5sNZQ4bE1cCuwq78mL84ff5craJaouACqzAo6T/b2JP0RAwjT9Rv7hB28YS+XrVHlwcpEBrj+
FPaimn93pk6R13hiU4IUlnCEz7+WoDvPLgONturMQRsEsOhO1Mr0mDLyry+0Rw0/WNcJA9BRTCKw
pc+igqGxyjxlDUHdM2+aKjq/sBEIGdlkasJesDpTkQBht2aJZ6YPkp6XF54zoQsvCp3WOUKYcJzu
pSA/FuZhffnI+eHdn33vrZHhS/qPjea/2pM1Rpw4CSF61Pkf+Q5wY9qj/t2nzoXrgiBKWkebQIHD
DB7iu+UMoqW6tFo7lEIlf6XwXxVa7uv9bgPkp7TXtigL7grrmorlMSWAdLllH1XfMPnIZ4EmoxEf
oPQjNNlpClfvqwnlahPdvSRdqI6XQ5SXv73nzrYEy7y0wA4xgLltVAdbYgcTaqMACyo5iVb0/Jhr
nP2KEIhVrrDdE013SuFAPE+/bGrH8uxzTCEiNs7iU7lpbSNIG3zMbrklv831x2lPR8UBj5Gsfs6E
pBnaqiKks22kXEusdQeMzQyCGM1+v0vDB7IPiLmvrRx9JEPYa6W3LnhW55Hw+qhOotecEJPG2BoX
u5+pkqgSrhroGhGDAZ8ZU3/FnUZt2ECFZ/8bln5Fdzpf9oMvv1JUXuQOP+WzHaPV8EU5jsP014ek
cJH/LI7/wT+wVvUfw0MOxATTJVmWcR/JLj2N+2TKq4oXRBdwSuD+Bh30nLwdFTS7HzqAI8hqEzZz
QhscqQwBFhsE9/U85k5UwoSz5AJQ4rjKnonfN05B5a/HkqVMdiqFCGkjgBxvZLZrlzxM58kJT43/
GHgHTEmTr+EXCMfIWQUnWzOekTgdLBc9zc/dzwWY3wJP2PrM0fCTKKBIFXsimG22hcXqjpLAyqsE
rCFIwb7jjo92cK1/mEN6/yy98fNwPcqACWk5lDFwCjd4ib4MJNX2+SufhO9BmDlJ0KD1hd9Agf5n
cO8zy8q8WDRUzOt7hHXDlLmu+EZAaBhYbuRPymTxpQa2IpcKGuK5Rne5yljfz5xiKTu2QyI59+0l
CVhwhGOk1/B3Vt+i9hmEv7nURp27gnX+Ohx8WdOV3z44+D+Zeb06+NyfjA8sY0OSg07HEBU/9iXQ
2V/hXKo6UFKFyXnZbF+DPxeJxind4lTgAe/R36Kok33Wpnc/jnod28RE7uU9UWIKLXuYDPUijlrv
8pDho891l2U4TUjcEFG2jiMz2JkVAiUld4EmL+p6OPqcBMGAKmTN+oyRDn7+LBoTiujBfo0ILLRD
y/dWLhG7ft+uIzKD3Gf3MaFgq/rozjsaEGwD0LPpocQdfs5plfxVxpaES4le380ZBubgzU3o4hzt
BkLvtyi30sGuHpKy5iiBDX+pRkwzMtKyi5SGSW1wbf30I4yE54tTT160q5uCmSpY/NNhHLoVQ2/B
DQJ+h0MYdiozZBHUpXtTkjcK7P6UsLIRPfh7JNpJs373aisI19Gtu81hywGx3pLIuDJjmRZ32SXK
cLU+1S4363NcC6G4B+9KrkPK2U1xBAHo1sHkqlKOO02YvdeBzNeeraN04Aqiy2evYIgA5QZ4iYO1
1EGNStMLb1AZWx8eSOIUwRlx8UizJDSB21+Acm7y2V+6TCYz7D7YZjYgXAgY5lyOrkS4Xvo8B8cI
/ncTtYMiAOCUO1Co8R/s3vGgraHWgS0xKAUwDrq+iJdM+1wNsQhN0t4YhWZq3MnskgkI+jZmVdjW
QMnST1vgheVPyy71Uds6+OT+3y53R/SIv+e+L9TJ/+J15jHNrRbIJXfp4umsbwCZIljJnf+S+Sa4
2RN5/yLjOM6XED4Oow1SUcZjVz6MHHkD2t60weq2CeocUI43e2OHFye28WWCetPws9LdZHXSPvEU
SfDYbLId49hZfKrm935UP55iV9tjg8BaIrgOq0QekEszXjmdYhWagIis165yXp2TuaRkHV3p/M9e
BMYUoZaTOCtxG0cIxJLg9gOGakU7B+7jKJAYKr2pjAbc6kt+3SAFc3OI365qGhU/yneybplKvd6M
68Sd81khZXtgp7sjTFvm0FiW7CB5vjuK0iULHUyvSByjjJUuQE3SmCZ/ju8Yin0T0gDm4aSoaKKD
NhJqv+bxSqUaNp+FB4wucVgQzOZzU4LiDLa4gkU9gFKQrn5B95QqyNn8crPZtqAizvK6Ttz99OUG
keVq5b5GMy374LMRHzw9R5nqQh+Z6TcGhi8vXulJtAomkyO7OZTtSKPz+GvE7cxjiPn9Qqr+5uec
RM3vUj3vZI71NvAEd2OIGD0Qlknp3D9ybI6jHdPqdsWTK+A0y39WroIOEzM3oCz3TrD5FTxk1gE/
kkgvKGyX0c8f9quc1zQx7pfiCTDyxz3Foc9zNjWEuBFCGwCEaFgMSN3yIFOeOROFA1/tivdDMHLp
q4RU+iifOroX1g7+VYqkIgAlcKzVNsaLK/Plu6fWwwhAgta4F2Rr+mHCYEVAb2Z0+JPDWjnJU3AJ
lD/2jVBn9PCYhe51jJLyn50o7CprDbuYxPghkxzPv9Xblt51TbX4jFVv919nqnKmhIla0/moMnkw
70AVkegsfGyWfce3zlSRbFXRqRzR+Nbsn91QP25m3bsCFAQ+wPtYbh64qoxmme5/Qle85SVLUB7D
b8hGbfXGtqGzm/RTuLuhlncJJTFYZ4gaR1+/E695KGDzY4+otx+XXhw2l6gDnw2p6lV6nq8d8dyV
PZm7QeUp+pjSWCQOglTvV/V0Ij4YTeF9nvhKARcolKt/POzFCn1jKs6WCLX9yCj5BFhYTs0zpVI9
p2x8uv+GtjaglL8L5VkuHDlFz318YUGrdVA53S4YBsdkrA+220spRLUyOSdEdxleDvJSvCtjB0g0
tolQA3uyu5kEwtXkCBgO5tEqIcyfwT8NgcvsQPhsysywFcOl6MOeAsScd9OBldu0uWlRqDjofTi/
Dg2Fvn60MlrQodZy02V1CzrYdKKhG1ZnO+P2dP3FcCqR1nKxOxPDAB/DwGMcyZ9g16fIYQrFbfLy
oCf9KusaFSmDAxDbUIVxSLFWoOK029zw0Ng2ayXaTiT/cM1+ljmAskdnx7JEgVKnUus/4sHpRvdd
GEJ0/PMGX6ZkfCwVeNLC0qUkrEBFGcScl/Z/d4TnsWpARkbqLt2QNYOaeS5lwPCVOiqiGiju6BXc
6Cr0fbVl+pfZ+Ammic8UV+St92kCL1fOaULR1SHzdwk9EmAj41wJrkuRiH3t+arnbD0t//RQeOVY
UUsV6DoQb6IAzKFYsiEHNMo4rrHM5kNhlS2leuuAJgTrKKisMZpmyq2RIj2dvc6hkKipvv+Qiabo
nnIXqxal9rhUW8f+N7mpjdElmIPT/4I9aI8XynBG9e1/Jb/k/KECnu8T3PWHHeiti50EG7tbZMZ0
UHgYDpTH09w6ttGmOMkT6KLEoj9kTlBGQrKiiLPj9u90zK07ancaNnCs8ZCD4F3zWvietxu/7/P+
XukAGq+x5QiIXh6yU3jedEOV+aMifbj21/czmoLq+EQDXBXPSJSH+R6iC8g9M8jvwsELpL6VwVNh
dmEXrfYvPf/PY+wwqZLMBKoq82hv6Z6fR19JsMoaTHF1k5wZ4Ov5cmAvamooRyoSOewTsOdUSWYI
mMgooe58VyoqVr93m9i2K+Bk2GGQu0deFZ5r94QVUScPgamKidBe8vm5PUxWddi7BonNzq45ZtxT
HDSjZymrmvLsLxwpXQ3eDpTGNOVFyrvr2Px8iigobAXXZL4qb8EWozTsjIL1WN3YwcQM+mUTjfu1
5OID/4PTYBZfyYO3sJilB4fYtol1R043+uCMnEFy6lC3eUo0+SurTwr6UK8hUmcuJMWvPKIZqBrv
fbETPqqyEZRgvTSlvHS2dNlAQbD3SW/PoreUSurkhDGu3EdjDL0cq1q5k2Sa/pqFXuWKCpMVgH77
xwktdhB4ij4ZhFEgLa5jspsCcRSnNDE2KOhLdLtKVo/xc+37f2ZLIEDXixkgKbM1plnqzalFj6tX
KUp8dqKsNExKt/KpiWrDT+6Mxj9elG7L+B+VruidBgzsJMEH4saMAsuXtMlmC4BtkDDcN2A4wL9q
CpwacG38fZaVCJPIjsvEw+HKKJ95Pna7f69KZGhC+WXChlLSd5IXjHdi3gZFEcyXWdxa3ZalOVtX
4Bbzn/OsBkU3DHP8L7Q9E/33dDHuFi27TAr5vb8CX06rJG6NpruYe9p+B22sfMQIlOOD+uxFjLPF
QM3e38Df/4BLUThZzt6IAJ/XqbR+8gEnyPgljP5PGYuoIoiBDmRSI3T0PF0gtF4EdF+kKtTwL/Wo
26ADjEAZyo8vHrKrGmuUjXyY2wcXJ2mpVSk/0MN7EmehU/LuD08Y8j+9xJhaiOL8jbhH8ov7gKb+
/+6yyoG2qmLjBluWWw8xcBbskwF2L6kOen1VDa3yImAAEl5iawu8TTayk+d1lzHPkZSzOv4f6joB
TpmUCHeB5mSor2HQ6eMK1zGKPgFSf/PdApEN9MAffpOKZnzgFPcL91v/NN0E241/mc2UqoX6aYjc
VAD8Idl68rqHUhGRdB7YFSi/G0QsSJjezhZcUVd0ddjDefPtEWk20nYUdsLNhhQLD/y7oVT3CyCz
Jmup9NFpzy3cCG3WKz7q/a00eFEBp0/ld45AT818b/gezzjCtKrXFBxVyOyd+gAoQFpNU4KptAS8
Fmk3Nk7YwySoIsPznpfVXNEdS9YdpRm+jMcPIUzRj/pOqiMK9KG7r1ixm/B5e3s0Yzosv3F6vNul
0crmEuH6aRjVxtuK7p/1fU/Faqknk4m7XWv6IioabCHuSv7SghVVrV3z2jSjiwCtqp1PpUYRSQ2J
PcRNik7inE6rAVuVRUEysqjlRp2iFt/CpVHzDuHhTPPR3e+H/VowSXAfIPAjzYLb0iT537DEGvia
+XFDRXblSltx5AWuGh3C9R1gKAW7z+Ae0aVqgfTL+Ad4JPkfbAGMUepZqu6QRlQWZIbUKF9+wRcG
cvUmBE1pOiosU7BPVwRE0f9MIrg/c0YTHjLiB4ZH5RycZv30yhz7CvGvMlYcgK+foug3Idg/OugS
ALqsddQ2XuKwsE+cIvxnjZxglTq+vBl49lrrpt/5Ng/khPMDE4Jlv3CCpRryb/TBmkJdPSNRT0Id
/v6v7aeD9GibgIh3qLt8Nucz8uf3mGfY0qYDGPFjyq8PgCGf2JXLKhG6F621fu2SxKFXNtLYn6Xr
HqpjTRZSmVCXzL3843GryDzldKqOkLUgq7HkIoTcZCY6cD6Zh5RDHXnIEQKs05MXC5Oxo4oHYxR9
B9ZlOR+AC9rh4jZfFzYW7XhUbVBvEqKqOiLJy/kVKviqhihpJkabfc/HV4QkrL7w7O0p4N2R74Pg
T34mHsunJFzMUweEq9MUVMFs0t46jbs3NyzOXhsEATh994VRmdUPL+XiiiasZ2TTAlcfjHPMQ+ws
XRkmzt9Tu0fXoZUMP5qsbq/maSdHKi55PhQ0vRuZCXesjlixGBt7tJgzhbIvj6CNw78wbCfwgjSG
vU/7xYtfmzsePsTsx1WHzBmKAGCeAx8hidtcEMiSu3kz8loZaJWyBkVsWk7Ok6ONKW3B4evUEBC5
dFleO4Fe/5FMSo9e+yKBPdRcfYnADAd38yZNAoUggYyVUYn9ZmoiRB8Dl1geJwXwe1zS6Ph5g4wk
4V9OhjVvHAM5rmAnMy644oDLv6atAfUE3qAAE85fxhm+OGTcnlC6RkQRALI0rpemLoRvlDXTkflq
+V2oE2HLiU8H7D8xpKq9x43n25BrYJ+0spOf/4EGz7eGFuXzD1LpN1iHWWr6Qr6NQp91g3mLFFTJ
23ZhmsIbq/s5uVm4bT6b/5rH6DWjiCK9kR59lrUDqAsPAD+fXVg2Ih/qKIYERaD27of9TT9JXBT2
hbbVWjBQ9bPpYTVvlF6RVldqyZruz+EGNxHATcyAnXLuwjLNkRms7PGqmJenddZUzSu9uOKuCVNj
29D7w/IXBEX4PyyNJRG5z7OTfUFjKzx+FSy2sjWfh3X/c7cH53YLg0I4ZV2Oj/ZFRrNvjvSWkbb2
nf12Ke0p/WCAVpCvqi+kqADbqtjuOJbt3801cXglkXpXA9KwsRRj+bHNYuBI7G51o/LR7puHbCkS
qk+9znIDZ50R5ehC0e/XBjCnLu3/TtPrAI6O43Z6M53XO7dHMr93/Smf/HVWFdenGD2BjfTwskW5
SgYepO2wja7QPMC4nOnMynewYe+fAoXGBD/uCHtycLP7UeVPiXjVdKuSvtcI0vTZ7YwjpDqx5TZs
zoyN7QZB8yGYL25K1YEf9aPgIlq2n5jXr//LNQRTHg2Pne56efgr2W5mbXNtNzz54k5/0MQJphLQ
crOvvcmXGhQUCvw6OYRy8o6ETKgb7q4+pko/EPIGaj0YNgQgZWGu4zE8ch9Lp0vl5urzZQSLHgNw
rk7Pvy5d5KsNNs2qLL7KLdQE7KqnDn5JKKfhsLRid/MHy/KRntBmwnx3KYScg48UPVylFTbeMBNG
8JRNF9rU3wytZLVhKbJJJkKYTbCz6ZRn8cV6qsFmpw/kTrH/g+wwrsFtS6Z+N+oyQlQkicRY4aRZ
GyuKVYo8j+a1NI+cQfLdyMf3tvBOixzcNY2CzEFPO6IIpXT1pmp8NiRX5/IklwYRKsZ1HcL0Vmdf
tttP6gl54LPqIKiTbNos/pUgOJjqANMh1AfICo+Rx/kBfLDDQZ+JGYKbfZeS3JzCRoXxPVj0Rqx/
WodbI1uoT42GXZciOCGrfeb4o1eNSm8/FboxtmRPMxcF4p3q6EYrs+yidH1tVm7HbkebEb60wp8h
rp/+8L1gE3+nR+SmDVNpSvQphK9u7IQoohtuZhTKuyNYSg1A2/eeiqF6YvRc4PcPu2YHYU5+Rwfp
dx/4ec572U9YdliJtg25Sl74iEGagZpWkqNC9yEF4KZ4VKyPmlyMp7EVoXh5yMNIa4GP5FW8vfm+
u7h3YGedM8ripaYdABt+T+F4zor++Wxyk+OfmYmggHnkQ4sZlgfhIj8gil6j3oD39Q5eV4A+6dUj
2svVS3mCinyS5Su0MMSSdysB75mtKhb6Uujnsa5ti9LqNw6IYN43I+jUlUKeeY5Sk0jEchjwfbVA
m7Dp5RvFXIqLf0urO2StoQypvqpsSD0L6Ro/sWfJoQY7LNsX09sx1NodFFCFf4TEMJqNRTTVbnWS
pKAGUWZhWC9cYDfZBY/Ng+e55kiIyPq+e3gsdRNAEIeRQytm2by1xqMb8D41GABkk9l93JD0ujgu
IDjLMLlbblSPEJ4YGucgZJDPndr+yNN4xpKBArRL4zhZpD+zKpJOt4I+1SUOYc3jGWfAZW8xUveX
krVKH9x9VnYhXwEN9Mhb9hue8LCzKilb7+3JsKIX9imuO2K8sAyRbvglAoSppeBIkbG89+roiIiP
SWNhFdhIZ0nA0fqsxZ8pTBRVfTpH032ItCxhXRwtAmYq9nA0NEKkFXfGZ78upVu2mSbR8SRwP9sl
vJblAoINgViWuzECbYhu76kfpr+SbR+ECd9qHisMfQHfXeK13Dbdm9vQEMuNf4OMRnY2qU8Fqitn
F50D7sxVpaV+In7Jfm5WbXUnl+GjTmvjtkTYtCf5ise7lLNYydHuZTBkipoqoseLSKt0UpxwXBIL
vw23FejFkQp4bHgdDSDFK19QZAjzRaEK794pLzQIJl55A6RdySsqh5CHeUU4mgwdVr110H0hl4/B
jMdj4ixpN/Jhn4G1uiWdP2f1bPf+uqYL5v+GGLM/7azzNw+reT6gwXH1n4uFVs1siq0073dl7lgI
9IMgiimSUe6FpRSDEeMpgew54X1lrALpWZzuSp5/0qJ/tMPtFqeXbHxw/Gvi0C4Z+i6De4vmviCV
fmD7uk73+rr5IKDZU1lCUt5ovtc7iRcymuj0YIgfjI8LpNxCi898HzgU2lk+nDXai8g9GIc1P/kA
Z8D0rDW5ubZsvxfS0xH9Lk20WSCIeAQxdAAcrDTacR0pIoXWAJRTzc1/+O/xvT5HCCBayptrD530
+nmOzOApMV4QLX3nY8ne0rm0PxuepCaCJe9nzyf98Fs9Fi2opQJYiLRMElhrOTpyJwbJKM93Kjo8
eIJRI1sjJjMOiYhGFFHLJC/6pqrU3mwc+kzuHqvk+sVV3tiH+Tzs5EP7xe+a++3t/2kYffekojJ7
PgeJaxe52Soy2lqDbNtbDAXBhlzoaIbljTAOYpGcdeF5S2rT3dHyNqURc/H91m7un+k2Yvw9cRpj
+UIzL3elQCtket1snYJS77CseEyFcbblT0oGiQexGbFbGigjuXINF8h46BIzFSHt40en9Do49E/t
j+7GLFOL+WXsfeKuPEqRiqot8hux1KxgcibWDDC1OE0APojZs6n8rROvp1hhEwAVKHGmdH7O6A96
SMcfwgUqCIIu0mwMzESTlxop4VnbM5ebap/JKpU1cNOKzxOQVyI1ahfTxBkmO4lYgzZYZt025swn
FqLhHh7Lwu6yTKMfsp1XIMCahHRAaac5a0wgz1CbON9KnSROGELnfN9pAvvvspJRQwgnyeVoXmrk
lbTBaT8reoL4sou8E2YTZm49uVbWUEJ0PVS2gJrF1camNi6HrsrRJXUUxDe/JdOFydr5SdQlvJLP
6uyg+pmKjeKlwf/bZvPR2ZyWaJ6Hl+4z33IVLhZaW3tWunAJK4VcFREMefqIB1wieE42kbmqNkuY
gY/FhYetU+0oK0F5uzODnrGuzVOAIjC93wpXw9hU+GN8KyLhNWSwtt8DQstMb7jDhzyJlWmLIGxl
Wl2m931EanPIVadY0PY8UphrwgQZVQrxrc/sQzZpuSFCwmu/Qv9Vg3PXs5UsJzNdjTeUek065UMX
anU5j8lOOs8UPalYuGxKeD+SGxQ4eC2IwGeL5pDIyqNuW3fRSXFFo3S0LjdpRB5mQQZzTYo+wfaS
shgYHOPNA94AOhY5yQH0dRINv1Nq/DAF85ai7ZfQbi8RWxH8R6YqsgcfLAYTP6532O/FrxGqpswH
aVL0U45ut/AsG12mfuDZfQq4L2tr5ZtZLEZKxDNsCTAk+kT1Gz7/KxyR2htyy9WYo8RVFoKEk/gw
iZ4viivdc4A7Q4AV/T0WPzX638WBhYDxOoRTP70T2bPS6jAFeeR4NyaDAxDI7RVOueqk+gigcTxs
fJXzy17BnssppkVoznn+ub0v0xLPdNDBNr2ztR7iOY3+XSFz/Aaq0U/BrKcy9LD1us7XlxH3oSfx
t9kaaHZWH2v5rBANujQL4DEmW+ocIGBWg/jj6Bjwnle6/rG+so+e100Qap9FjJqhit2HMctz/Sok
waHxDu+52AehdE33s1qz0hzk9PRPgWSxDjJ0ZlXQ9FRuy2Et7JADFcQ4dtWAKAbFzvo35gQGT8oz
oxx3FUf0FCRdJOYvQe/Zb5YJ14WCr06TjA1WALCDffbs4kogQARNah0z6D3l/OKXeLP2xhiTl+f+
NbBEqFiONpG9ye49+49rjh+dhC9C9CRE05+Kl5dw/0ljtbbHxkSqCyPrDatjC46P3qn7w7iUkSNd
cX05Ju6RCxvnJRW2Rm80JGpd+dhlPkLne9Sur5J12ou8H7sfGkSFOvzKsnF0u86UAq4YVmKPA2+d
NJsbOuWseJneo8tsLnTqFKxriA+YlMEvJtP8lOb2fyu8FOxgUSvCrRsFVCKynq3EUbDmG1npMnhY
oawBtPa77p0lMIeTC3+1NLg0p24/JZTnZwnYBhUAW2dZSaNbMMeKlzMmlamMmkCzvViGPFw+vY5d
iytjxEMM5ByLbzRt/+vz8dgkIf8A4axPdQ28OM/Vaog3rpNwUI+uc//Orr3OFIMmK4NgHt97HkI4
XV4kXMxG2BDAt6DQ2PHkLAuUsS8g6nGqguzVR8dJNpSiOCn/GqFnF/JuYIFI2bTfSn8UBk4zl3xE
rbM+dpSSYO+1gnlmNpCzskO+bHSMoi8VA/7Cn+XQXjX2ptomOz0M0o0hWXQ8KI65ykABvtREh31O
keumMYY5A4N0CKTMEZmI81HdFYmesTuiIlxGblh5tJV/Q8+3nXfUA6CVQsJ9t36qGL7EmABbtFKM
n0wA0XipBtOn9HsGy92F9qyODjX9QZn9SGEBtWGHFaC9Nx1be711sxobyIaXUEtn9Z346rX5tTg+
2vHAjun2zLBh70TgjwBMRZuIVHLgtoY5siNmswVv7Cgpa1zPbtGeuhe1nraqS/xu9HxT/vAhcYSE
UsB7jGkMDstz+R9+dI36I7YpHj1xd/GRie68QAaToiHlKBRvcvUxe72SGQiSrSTmJ9ehgGVBhEYV
ILQLi2r99fYl/jEHrQxhveFPM9jG1Bj5KHGwcQTDcTHDC1CYw9mPg/jWDh34fz/UwN0b08OeX/t+
Weovg0vuOojYGwrWoqsF0sjQG5pAnd6lYxncD3FtS78O3M6vbclMhFoeIBoU7KaHm5q5IYtuxha0
JHSKIxa9i2OeFjXB3OnO+JZZbAFGXC9vWhJM03xM0vr6P9tJTMr2z6ydMgPC7J9ifOQ2SZ0KIREQ
fDuqkQv1LUJjcJuV23ucw/X0TXT8fangPxhP5LZYOHo0Phw8h9TfyeQXw2afagBVQRYTefRjB4L9
Jp5q3ERoz1RujPXPCN99DHPD8Hp3S48VvdB7izmxY0PH59z+4vHNgHcmmZg+53ETip71goCa4Lbp
Ot+U/ne6mzCA0TM5ipeZSspJ7Zf4DiCMK2OcANPDXUSvpLQHk1+r2xmrVJ28ZgL399G8yweC8a9T
i5mcnThbK+h74bHXrXwFLFHCtwcwsyE5tVeNkzmtKrAtfdzAsrbEeI85FC/GG5J4bBl1Su60ripE
eUmCG+v4cRGEJTFI1k/XPH+L2Jo6JHFi7YF6bsdRpNO6mb+VFfBPaBiRYCHLp4rXPsKCc8B11eJT
yRUXIEtNe7ACECWvmTF6N6CX58L85mxtpe07cTlfQVmP2D9Gkdsa5BM6kOlpOLMiJabvIgPQJNNc
ml4H5c8UHncQTq+8Ef576V8Di9wOa611s0Gn7PQcP7VvR4w8VVZZ3DBg5SSMzk2KJjIkDDYdBfXo
v+jtVohqPQxkQUGBIVxw2FsORDPOS75DDX3tJ1xOasm2Htyq7mfmhKaL69u9kVPVgOukfrJiy3tT
Umup8VOuBRG7s3UjF7pYvH8Hh0sZbFwX7+BLm8L510CIHcnfNmgs/qJCdyX6870RYen5ke6wrFPY
fybuEXa3XO1H4VXI57fHJjsXnx4NAN11UQiLRKf5RcjgHWqUrK9xnWCrgZrqSxsEQpKu2IwhIfRU
RGICsDaQkLvLFSSZCamSsxqSiySHqwQsaXyo9+Wd5tv/rQSlg0Ak+hSxWD0knOCcK136HMCVHl01
BJ1cTiO+Z4UwC/HggGxCBT5rmt1S3Xdzklea0I1WlcYY5jpVHI38bpTv/tNjJesdslzIOYHP0vTo
zAoj9ZJnke+AvbJrwUp8HzWwJOIRLWZQSUjqEFk+Zo0bnvSOX2ZLWqSbW4W6TFBO13qT1kZ/BZmZ
TAv2bJORfYC55x0Pw3xUrG9+chIVtuiCYVnqtDf8b/7WfJeeZ45HK/tIVlYoUQ0YBRxBemQWIgXT
gsnUhQLkxRCi/g7jLixx5pMiudsYPLedqwYiu5FJpHPZ1KY+aUNkIQsfk/AFNNAcaCRiZYVY3cYJ
0KKM+QNWISm2sIZmy9YT3lC3cXoCiJuxuCem4st1vhDJQTVJ7Hg8yskqcyo81HHHFiB/+oImBI1E
wC6VMlbJjGqoLeiuvowFE6u28XCiTUT7IVpvm/GGml1EVxGRbv3y6P/KfIgLNyyvYQmel9+l2C54
77W0VqgU5V8vmnSPg8RvLPLcssEix0EOnYzRjPm/kKyC7SwneFp36aoh4BOnRO7i6p/AwWnFmVkB
K7uvNoOcKV6A58KaKHbCh/ntnSnTriAlVVpMA/9qM21wAKWZiS8n4yCR1arT4fx4gO2PUQ+dNgrx
UY9H4s0rxZNj5HWxoINFTNUjs7vAUDY4DQgWf8uJ/29u3qi5+IqZrTKR5UGjwnZiK87S8ivUYm3R
/aRGfQ72y97W9K4xnHnr1o+QUgodPMAzUyPYTagPTAW6KyLyILV3A1XupyoKMM+ofsiQRfOMGCkT
GePHQjZ1lFZLiGap2H/ict/U8HEYdqDQlIAfWp8jmQSFDcR2QeV/xKo2QFoAXps4g0Zhr4C47Hjy
RIAdxjSHGwQHqJYUVYdmdv4Qx0ulEpQANA5x78E/NhyUBPBrBVp5c12rnU/c6yeBg+0jmwSOLBxj
hc0iUI+qTIXWLnu/SKlv7Si6nAh8XetXUZdZE0O54/+gULQnnwKj0LG1zhdVt3qiB70Cx+lgnaqo
uAFw6uTxwKbi+ecgvfvqeJw0YYRjx/5m7nv/QRKmEV0wzFhkIdiRcRM4o8xpnkx5hJGnBeYXaGh3
Ssvc89haER5nqK5jDwpB/jEZkPD5Pt+BaXGjHnyaar+VjsElTiiUJI6chpmz7z2igVf2HUhpk8gQ
qHNVljATyv6NKrRFgI/VDFe15g8bYBK9HUrZzjtuACKkQzEVnwfwHgIDt/4UQC27vOJu9MhDOWmH
X/OCYXFjIT5Jq5pz5aVh8+K1SUP9SDW8+lDX9c7q6RjR+ZeTgE/mAQHmaCww/2GQCB3Iy/UdZQmO
xybfkM1mEYkwDxIXeSLjaTBQVpffLtcHyJUeUf9keS+PrrHBDUxDOwJL3dvkRS60xBhzj83hg5tI
2dCzYkh20hShU6FkL5Lc2/uWIN7+v571DUjrem/iNLkOb3eRB4slFR9MgUHphZ1R2o6sikt7cBfP
c0rjp0u5A7nabT9Z5hZxHmZWSt8gLualU6m+bK48xd7d8oZdb1e2V1HVe3P8iYxJQhjJYAjBsY7v
miJ99mL+XD2LvqruR1DA+2uVyGGQZER3CH8t5pE9DexqkUnRnlO3gF5t/AhbmnIGaA9FcRwMjmgR
B+faMyflGtAqxw6Ykk9z7WF9vw11tFy/y9ZNl6iiihhnoT2cid82D7I1/Apeg4PUYgooyXI2hFFG
BIRtJPcxoFw1wV9CMsj5GD+GBqtIHoIu5m5WhWTC+A6jN7zRM1Kwt60obkVj+Omzhyb1S0FwXpvO
HmhfdxeOxmWjAIkI9AkCPgVJ0t13CaQcfQ4zFYuh3xea1a2k9WrBXpH8BzVH9ROJ4XMGy6uMr+qB
FSxVrs/0Pi/rIzhO+dxxkT/ffHhMK8CpcJBoUD2ohLG5Nojq+w0gYZ761uBzOYb3neU+sODsW2lD
tgjGGh8ZMzqNuwinF1JmGaSxjKu6onz1gL4RlZD6MNBQZPb2q3Thm0MhvtDOCSOrTZ0KVk/jXCmS
qv6C4YSg5H8md02zXZEQLDZClW7FQGIT7BuIkONZyqB5KXWYWCZUNsVQt13pjSk+ODYfhRUXw7M6
CxfC344at+7/wL7EysZqrg4kWFsF1Q7s7MAF3+CoZcPcyEcNV6mYs/3HPkdOkvO0cMTCo/bRw+ub
Xu5IhURYHa1yzZWpLros7jTuiMSVR/mmFHMTVAOFojNtwqmqwMTxga0j1wcwo3TVoEtfeuiZxY3u
5H3zfNpSdtWJTLOHm2dGR/KtTh5ixCCLC1rLsNV1ZqGgCbOIlrehD1OiW1phMd4nOmq+iirGRRI0
jN6RtfyyXn9XOgJgNxGKWieBBV9ZSRr6vc5dQFaMbV6DJwhPWOPU9m5TmNmc1dNf2d5r7Zu3zg4E
vST7NOZBAXLC2CQaKY1XU9grIgcg28shwOobNwNsSSEo5IBRu9v8GlGJ/8YmwHHJvcGKe2xdh/SE
4wg/GQSLS7i2JbEXyZcQ8u+3hlaIFgpl4xRIv0Wbjp/UiRWo5IMvtpzjajt6I73Q3binRu6Ez8YX
r+fKqy6YgPM4Z5LlArBtRVlXWzRJz4PCOsysK3x6+QldRq6XG30nRIe5kq83WoalqV3B4GukXt2s
ZhHF4li+/QV08en4PKBqYkf/lY7m18ngMgov4ukq9XyQ28pT/+8CDYO3QFEPcr50Oo3qbrf53cQN
a5RS2SewLd7E4vfKGwixDrIiGnhQAy+HqXhsaRiPAiKIQ+CIfUfh0J9SJblZFg9qtf2u+x+tp1uj
sYJzDGnCEtuJrnPu0uTLhJB/7pqJe490Y3UXV2Z3WH5BhRnirkN0+6yMLUNHnaTdLqnihEBRihXv
rkm9jRRJiWZ/Fn/Y4jk9yKytHac2p3lEMZQYaHqU3ABOYtQe/FKcalYZKnOaLN9crloQeOEzYD/w
BIB6QKHJr0pcAR69Cx2dJwmxIUgAERlnxsnuPzml7uWFATczYLnWBct6ZabbSf8zdmntnApl4Jh7
cvue2NsFsuPVBzdPyb299shjrEKmEvMRXfTNxr1cofdJeOl718T2kBtKHA3BX6/rFEMnDPKKcM4W
POkm/ym8tZNllkbpImDRZI3+qHWnH3En+ThOHqhbirBk9i8z7TP764MATwbsc/O3rVLnN6CRsXo1
gLiG/o9IO+bJylLRYf80x8RWviopV+tZCboUhXjnUn1dJrbN3Xmfo5jCd9YnT8BGsiqxmGzgqPuo
gRPJrUlFbRhEQtJNm5tbG0r6/JSlZZ1jotGrwYKln0tqFqoKI53M8RIHevtrMHfIFOi82+PlacrB
k0rLOGXT3QhiQaoBy5BiLYlmw7c8l0W4Ve5nzE10YsnJFcIbEjpQMW6mx5qaNpVSDiHaMFE4lIXN
WWVUAe/GI7ZAeSU+rJEtmh7BcI7nnpF4UuXWFAGnzBT1NZ5hjKpsnXAU7mitquNTj9u99ywnhXz6
4Bt3RCMa1fOpNl0xVx8X2qU+qgwaZLMxyGCGJZ/rR4GYoRw5RBWryB3BeNbo6LQIc3+QL9g4yad/
hORFy0YB9AoqPS6D5rAm6BZUQGzmIFxfvgrOJMAy19M+wSGwkQ6gQCvR56U+qGFz9zg3yRaesXJE
/0IAMeWgv6+J17F6DJDROHeKWByb1kmGkwhuItiFiWlA4XRtETctK5FIKUTE+YfHV+i47w67HyB1
CUdU5TIEQNYCE3Or1jpiJcBX44/bcYox5Y3OZksGJAonKOxCcpLD0NOMdzIBQKc//QnCE5mygTWQ
B/VkKz29sTHVRUliqqt3Pe+lKLrEQW4zo12dVrHeocQ3tnFuVeownWCbN9/6pceM8xljkv7K6iYU
xgqVUUGX8yoTJKM6xVW/tvYDRNjg0d3ViILEjUJukCThb+qiKs5te6VuzU4ua0BkQzWevHZdMnpq
RngaDhUHnEquVjLxXs8TW6278YekjkRbJRcgPoqucalYQgwzxkSRnXrlYs7N45R8jKpTUJ0iBTpS
CIYK3SjR1cP5AYYcD2iwNdau/NoQckEvOWLAQ98j6qR0Uf3d7hBiXNLSVBQmxgGygSedXIYnNDHr
r4rGifJKz+2nTXowTwMWX7gFTDIqUU4a1WbDHcTwH0FKcTkGhSiJU7VP+8UW77bilG6Etbliw20O
faD8zhD+f3nPTZFlsqqrQpH7NcFh7fVx/UUCLjc06dxXx9UB7FAlOCm27ZukH9KLtIoNVV50fcWr
4IMW6/0G4Wff9y/UPKsrvnqFpOOAMxnpkTQ6hKJ4lRhoeJzJkPEwe7TL/5+/sOCEGebysGX/0V89
Dd2jdcwz3r/KE7WSUP8Pp11DU2jXCbBJvFSghGbAeGKgGgAzSHN9QlsvI9drjzT+UemLwIgmJFGA
yO150eG9H7yr56YuRrLvaJHu8k3r+CBQapKukDRHOeSZTbzKXn0NBpY1m6B+MyM02RiIeFXxU/Ht
+/CUJvAS7PllXE7/hhtdhIlX4G3cBWRNXbPWTbLVo3ZfHqtKQsBWOLjU0uN+/j7nmbtQ+BqqSTk5
lVFFq7aal6TY05qOir0gi19dZcrnzyQqHnzMfq1XJjlA9ZrNwZ4uTmhMmlOSnJuzo4nMugd0JpBr
LNRAoIfQ3cETCl0HhN/k6QSCVetawhB0pe7CKw0RMpQBmHG6vQ+VqnAXhJhLvguvfbSorXzA/zIO
SP2UYUMA/GrLgknqVTmEDCNmCWCYehYlkDP/89gN9OFqn7Md0bQpDlKyTVdgA8H0Xk0sAvPMGXDR
FzeizJBAq19Rtkqp0mVERwWUvFUP3At9m+ca1S5lA1jX9oPsyKOPU7WqXPD84lgLCREge+CCIG+i
fgItOReqIGuHSbe8PdeeKICtuy8Ylm3XlLmsOUddB+c+Q0PTPFO3N7Bksl9JOerQWjrYSlVwUJ2q
EMcAgU+tAbkbNAyxoxxmHo+RmTCUibfqoE9cKefFk1/d78skNsI7KCNLpMlSUpM5DRUvReBpFPvO
m1TvoSWPee41uoPQnYdA4lvhzOqPsCpT8pDhlJyR2Yuc6Eg5+2nTyY5kJIEiRGs1XAs3edZWd3zt
mqcQQ0XqU9cCq8I4OG78Wl7NecyhTg68ALLGqw2Es1UXTZI6pBNqf6PTjNvpyH1zesnSnQ+SHTVx
wl7nAcdVXgN0NbgOHvq5J+m83iBEZvG5XVyBaRia2ZQaBZjlwoa82pBw8KpnvA7/PbuJCaYybPlD
L2CD7BkFC1xl4eqqEpmbJDE6yXe+SZ+yR+TsWL81iEVPYGQ2flEeOUVBaP835Cuvo2HS16EbY7qG
eiSa5nbrCl3w6KYzO0Lx4vJPjNULk6rhi8QFaawrwKS//Mu+9gTPCtoTwRPN5hbYRMAqq9yuXyhL
DEoDz5kF84pzdmkgxOx2H/I/VUPbj8v1aI5zVUQ9PV0d96iMvIIGgewUAf8U3oFLPGQoVCjGfZq1
s7hS9n/8qzmv1Bn0cWLGRwaXmLvORI0K6N62ALEiQs5p2lcow8lh5XU2ponsWxNZo9nuv8yNIxAf
mxhrLngROm1QPp4oqRnWDvZlVMjlK1AxZcTUhc3aEeh+TH26Ovu7vQ2ElYKolOZxBtP5g0cumTGy
P++8UnXBFtk1IagOO3Qd6s417I3T1Enw7TC/TARfgqF+ICArI4739BM8Ts2Dhqm7Xt6+LAg/w6Ng
BwO3oabMkqwNTFGMiv0DTbhtU+rRE2eggqyPXoLB/ksN10vhXinmfm4QOVOxfwKK/AKrXaLVhvRZ
lNu+j/UVwIIBbZM68MZbyVk05cfAAnzgr+fHagVV3Txpp80ISotMHI/yiKgg3GbmP43Nb/GC+QwS
QBE54sOY6zU62bNXSijKhgossYh3rl/pSEnzrq8+t/pUYx+uvVhUUecCUg0jcj0TuTaHw//jOp9T
o1SM4WO9myv5RwKd2aRTraxJMFPAdA96JpSz3zGAaXcnnSXIzOcaXytwt44elA7dJRrBUfGSXb6/
u/6ZmhJAezXzqHFr3P+SPbhxJxuZ0fyNvrgAab9nIyPMpeLmTbv/sMWurtsJQn41+pHsyhn+t0no
y9pMVK3pEEXMjMzD+8g8QJ9Av67MmI/k4yBk/lkVeOFGXya1axbLcj12Uk22O6CbRjP8ipbED4B+
/2d/GfkIDKWYICgTHnZBUHCLcR9KN1vs0krtgHpKPUKyH0IC/2fTJpipkmcoGNaQV5Yt+WaLXUAp
IABCBkGO9RLOuPkl8UjQpWB/Yav+O0f58Uw/Tcx3LaftyzdxBvGF6sTlqGUFQfXmK19sjStQHScQ
zNzQLDx4zPTRGHI9t0kh24L4RQN8ePxcyUKeZJ93ZensknYHlBQjW8O07WnhT/XBokfMfI22q8ap
x3i9nA38yvqofLt0CxuWDRdUsDFrgEtGLHTcVEk9aS+4nS4Nz/n4M8d2n2s55HyxBOJunuIlxlct
SE6eYopmRJFUsHfMGoiRzoaU1wwrfF1+4D+d2I6X1/otNjXqKWJzeIpU9Omchqsu4d2Gw41unDT/
hdgsTeCaNIFCUJzMOb9gJevUsE8hE/HA4y4IZEmHwsEhwmo+GJrWWb7OCN/7JfPpQ2ELg9J8s9M5
uWi/GC0NEqyfCJ0i2p0u07EOPlib5eC9la9gp7YdiiSLiqqQByYtxpYSj978rEUl7kFYAV7wnPfu
9I1PpZJoydZneioNkSQlweEXNoOcOtzQ8ZYMXwTX3JCOnJU9BgDimFHl1GLK4vMfsSvAUpEHAoBO
9dC2hOqeS+f6MdO/mASn8YxTcuL0ebgit1kN+YpwgfUjGxo9EtORIDMfAyybMkF6V3fElJaK7lCI
hb21QK3rT8gPbZBqqH6enpuyUAumFQ5wxpOXzLQVhBbJMefobB1AOhkiQqKD3zNm/xCNG1/+9Gke
DCe25oPHr+s2RB2yU9XnSMcEqcjymQkdJsMH32VRYpoG+sCYhhjUERkOx5AzcXEZufmFYOmwt/dE
XM4se0TQfg+AYR9KmthFBNaZXZwyEuQ/kyvk22Yjxs8WZ+5FBOZ5A4jtpsyDVJ7WtWWOgIr5INq9
vczi2wxrJDmvlkEW6gJPSWwlODi9MxEqy3VvMrMEY6R0r/3vCfnLpiYg/X4Af8wwwYF+ds67HJnV
VBldrJ/cuW2dWnxtZEV/ywFjmp0G5is0iFxUV93vJ9L5mEoUR4KEvyitU+2CbiHmO/9QtEc+MhcH
LWYWnXOG9AJzd9ftb4pIuVmEiuig86HCWh3vDRLBqdmDzcHbHA5/aWr2n2OYD/LBVHpTQx8OiAnZ
lWEF2syujJLgicZBv5k4d2YO+Vff80vX/MlSMjLwtc5hHs2w8gTVyvJvoy26XsCBgHsJ/62J2rbz
WqsMIM7scT5MKmmBQpTcgKr9a1jtRZZHC1MkmcyTSc5fN6MSHAI/fXusl31pVWnciKWvArf4ERG4
Sf1XaSkUKGtXav7Z5PxfDX3ubS7hvLjmG9xSM/kBMxJHaQev1hzPhxtu4SOlMDoIrO+KgGjO5ENh
Bbm3ucGmLZM2WNLq1rX8ZeTmVXZeMEqqF2jgSTJToIvS+ZZ0GjOScKR8qVyyDVKkuZDPTF5slJ4P
8lLkJc/lrlKRzdBjCR+MVRlUKIeO49Cj0V3bLgoifLmIDGun1zF/JvfzTv2sNQ6L4cGr4Bhbyt27
PlYfdtBvzhGp9c3YyReuuvEXD1VTOnYS+SdWGpPX3+cjWjgGtP+MoHDQ7qxstY7begTvUCvIGTKJ
mmeEyGll7oWaIctzc2OOh56knG5jV3kIMYBRN85UviZ1XesgPb6fDFb7rYKJu763WjNmfydhT4q8
Kelc2un2wj7BjLczkhj97mVDicJ6kcIeFpdczXwwib8f7CoeOQ3k2CXUohn2REIYKKnVCFvqxmIY
+RaIXKw7dDoBfLdnCyi2Xlgmp0UZFQfWoqZPcn9i1J4d7ti5SN9UeJWpeOugbM8ef0UEn+tifNcw
PQ69XZM7hXcd5vzonAz2+MRhtXMy+jEkIXCQb5QJoOQC68jQVvQuMLePHELrsB+MqGwzLNTetQPz
SDIbXlmgc1M51CDcPnYEPPcmpO/YWkRnKcIOZ2dWA82uKOXA58gPTSKgu/R5Sp87ta4wjfmD2gGc
eF5e8PTddQfQW13ybnBFTcnA0Zox6qLW9snAZ+V0TzWrVrwCux54Ov9x0O/ZC6S1XXYlDmEKBQm5
QZRg2xeWFHtS9lVpBHx/lFmIbkNbnMO8SmfUQp0vnKY72S1rW0G6izOsPo/+YZHcIFyxY+2Dr/0R
izFnDGHWfnWXjnYCJZTJzQUDpD91aJAbpCVScygkE92xbc4yrq4gcBJ+/GSYhTpQ6S1Iy+J66B+x
wMIOFMVwWXObwy2FeX4xs1xtTYJ7RtMkANv9kYbb0+5idYZ0czl161SahMiyxo99J5xBgX2RUj1N
XQDLm4DQfH5b8oKKHQ2Fip3a0X1RtQq2Q4DsEnLxv0+ID83dkKU58eROZ7wC1IeBEK8k27MlON8T
1u/tt3jJBY6Ri/tFo2kwd0WYFgSRJYpkmA/2PlHLA70Gvo8JuKkARnNEXe3hWO3xR+G4S0aOTj3e
gnXkGhzwq++pPNhr7eG7Y1NI79TYiMe9cIQVICMUG/0pgA2cc6v/byIdpIBhfjUAaGx+0qbvGsSJ
sxiblv03mW8BgGFAN2vLDpAsi/by9c04J/K7/M9t0kWATwLET6ihVKh195zg1uH6ZPg8tQXHCZlc
7CZEcPogpFLdaUCEGH9Kh+54txgZqU+eUJ8+bi6Fpefr0MOytLzyRYGB1CGaip6YKOwkuy/UQfKU
u5qM6V2w5v0VzCXAsiwkLmrIWRzmUfGa8q6bIVHVHhP9XhsSQdyre5TSNX2uYvMEfkIkdIdwoM1Z
1wDzaZ1ekFOUKqWqPiwCdPdDwUOQzyRC0sB5LBq0Di/9NZhwcLcI9YQkoKBhNSoizGNDNZSRF083
XxjNIqzsYz5f/4YNco7X3aMWYToHp1LOjh9U+rBbSUBExRt1/aKGKlWJGNbbbIvQbZA2Wyora3Io
YkWwaRtA6yPOGIkSGOROpSn7iY3zeZUCzqvto1E4wVZLaU6eMyVbZe8Uq9ZV6h6M1pJvDN1Kjwng
GgOBFYGkf2tpKZGbPOZQoPTn0Kl/IZRKNEhHi6gki61Pi2HSygVEEZ9YMzhWOTDVBuCoYa79sQLv
HHK3SEQSSILX+KREYcq1+a1okaBfmg67roQjrLEA5DTSSY2U/rkY3z8gTkXCrQ+F0oQgQyLfNZBl
H8iqyw4yMb+DRrE/0KaCwl9D5RTknRoydnx+8K3xAKgHdZSWDf2+9VCGkj5Bm2eQFrWuNjofRSwF
WMrE3Hx1KEILO6AfupnDF/JkR9hR/xhyMzQa2sUUguxz77LewjmmAbq3dXI+bvclmiBBajPUo5oy
q/fii5Gfb9NkmUrygAB/3bN4RtS5y0KUkc58zqNzmOcHkWnx6hSP8epg/CuxkE0bczVCIapynmMp
2gIJRHIIV15vb2H0tGWv/S9b85KzrS8zyAe57uKCFo8v1Lx59C8FaDoKTgEU7bJ/7u0hkCj61cpL
kaDt3vD756wNPWbsr0TnGu6eKksssFlKCNepqHgFd4CWHHz5T5OawWoW6fw1yz0V8iMybzpdVhW6
E2KDyygAjCv90HJcz6cSAym03qw7kg/FkMEcpmQ0BUBgXO3zjvioI0lopp6yXOdYBvkJyTc7MsI3
E4XMCWoCz8MJEoxd6izI4PMuqEmsdm/TnJS9knKxS3mgg+9Zr4+0uWI/H4YmFaz4NxWNhTw0bbg1
Pbu4fgPPsPA3gYRW9LE3f7NbfjrgZ2KwwiW/KmN0XumOzqVnmoaKXag0IubQHWDy0UlpsolrHvXp
d2LxSLropJR+xEPzVidfTrglhKwZL9k1+x1qh1Vs519td437kwLYCtUPYnTJFlnixsa6u7a7C4CM
R9ydZvEUthQusC/OQAPVSTC+/dHolirVZU6qtT22zE1yXz5O1aaZTDXLIettdTSy3cevtBrU5WXg
gdec2LebflENxmzxZx/7kHsJE35bD+rrhn4/qKJepHilWxZ4uNZeVoil9oGtetjWnd5K4mPj3MM8
OtLnUwCPELqZCT+xzQe3MG98eK1tSPtqW2p+9VP7y+ytP5FtDQsjgJ6n31Xe3q8lQATZgkiE286v
h3Jg/2HaqCnBise1Z76/IMqOqnEGFE74/J+rS+Yx6/pwNLHkFhYu6YoRs9qdug2hwrkbFFh+WbVk
7NyDSOkQ7/krVoQXTSe5pLUhNIj15FRNS7lrbnGCIArkAIkkdkRUylbyqegZaic+9mehRycmWv0m
CqiyuYMICSV/gHlYMlzany7/6c2TH12FYEZA1aYqywcJrKhxzV1sSfQ/k3g9MxyTgY9FKbu1fGln
Tvxta3ZCY6AAxbUm81wMYmbOllm9XNwIKNfvM2WuXZyOHvY7dFkN+gwWPuAqIi197o+PofrsMw/x
J1Be4yU9QlQ0d4ZehFAFLk1Wm6wlc+UweL+7bHrZ6ErdUvrPBO43A6dL0QF8yoZhT9Y2j6OcJlj5
mq1EaWXia3TnmhgKDFp8CwgyVIgErPrynMP+etZvJrUuymrIP1mrJ22epfrZTfrUt6PfjsQ2F5sU
dL0KyXdYdAY2DD501EoUCobyqpvXxL7WTu9j5JzOhOKEjt4A4C/No6F7BkU69+uZuzUXFfcZ4Dc5
TuqC9AP6+RirlQrDxT0jZc6ZEMfh4LJP/jdyD0WI4Ax9/PtmMB51XdgxF+NCppq18JLWSn3uomgC
HIYhSPz1jqK5ZgY1hYaoG4s4CPCTcRB+KCALBG0VNvyLw6H+RbidxIiDMlxY/Vqev3YHS0CLnClB
DdM0sifnyb1BQoOENju1GPdvmzWKaTTdqYipPejwOQ/YlDASWdzTuTveHAB7+5KelipReNhWs3wC
EJcFZCwjpPJ734/gqIKSt0ugrcuCNXnYO+BFnYv+zwBQ/cIRSRlrK3NQKmuyJAfaxMWrMEo+HJAe
CMhJk5KIjkBCraKWJODco3xkdMtqI17IUpnycl/jxGQLPqFN7rhRN1vMxm/F6TaOCyJSugL9DHhZ
cuQud+24lduN0LeLwbv7BHPgUKCSG5F2t/IhMtXIlUb+T3/wmwAz6xGG2A+LnzfrX6FlkQBWv3RV
8Nj2Lmmo14tWUBZ2yvROBEbyxWszi+bZUzSdURVQadUguHKn5DA1hafqOXKmCOEbOtMlQiDDfgNh
XyIC1fMeGchiNgVn8QL58y3Cj9YYt6MAm6/yFIAJnHGnjFPSKWjoHewtQzm5uG8Vs2xh7PiiYOs9
8iIexSa08sGnHAkzVWu+BYz08aFbhTffB/63Syfh1P5GePYw/rtVByHtS5t6njTroBdzXc6hvMcY
4e5jK4MpzKvE//8wKq20rTUb/pWCCJecW86KJT2YUOp0Bwe0bZCcc5I2mbJ1WirGFtuixZ1EWqlM
N0Ova6y+7iUWUtODAd85sOGUyKLbi1kL+WUhlVXd9+fmhKN1mXqgE2zNvxZSqwm5F6imKb24mN7H
KsMz2UGk3E0W/286qIEpFQbJKD0ctgSa71pNE/rZ81jbA88cp85XgsFoJfY4VDdSIrc95XpcQnTo
b/kkbAqFe10nsvY5B/pOIKB4ZwzPOMHa7J+6POfvzPFKkwarxdv3Dh0YbFVH0EglM80y+MwKFZAf
gkH/G4IGsRSmzApYnyKnaohf75FEq/JBB2vLaQdS5TSTzpSjmV3maZ9uhhpSDG1aTU2tVJ/NVoiT
RiNeDJ6kJ1P+YH6vhsAnOoUn/YBjzFA9ntLNGxMbsZE4CeIBv4v/I9GTLRtax8x6hDXcpyUfmSY8
DkM/19Ikxdt03BKH0OM0qtYInriq7gbtsh2TpkjtExAO1ttK07tTczXwDZGFq1riZJ/Dls46PoDP
bAdAMkwSL0eIZGLS7VkIScTwPvgKVj5wcBUh2jdzZQF/zt8nEpKgtyfHhcQIiGkCDHZmgXbkXdO9
/f6aL/nUVWr1jCLFhZ92poI9UgtdTktUti62erzsg33ytFaWCEvRD8uEMVbXBoCBrfVrapEMZSzm
aP5n4dIBnokCipHTxjmQzF3MrdDekKckEL37s+rWOq5v8K1F9FkpstTNSz7h2TAIvjFO11xJ92gz
qQ+B4VGcF7DAy9vvgO/GqKwWhxuNNQ6iNyxs23cfD3s3Kf822gX+aXumiEwv254a4L94kAcmojNU
VpaYWFI+kB0062N+/jHoSipzp+jGqHDV4RCdDdnLWGpxmpdFjvWVZG1+OIojvybEzT7EJGzb7Tds
IRTNW4hgZG8Cazlmd/H70XtKgq9RoqeGeqvFeEqWXPzI4OZibHifiCiDPLMhV6tYz7w99IIFKRFN
JlM6q03v4cdTCCF9i9I+uGCqoHYOQ6fZf3z3tcLaJk+SOKIt2cNtFNTShKd+7irJotFHckt7VrP1
D2oVHVLAIEHRKxgeSuUhquMwVkYNQBHOUmoKRqr0NKH7z2GPQvMpmkzFCEPR9DWBEijtg5sKQ4N5
gN1gP+IGFi2tZLuj3cQr+hinkR7ut4uqUCJoVM/wadjJsB1Yqy7QImTNXc9J2PGWme24jhYlcyY9
7m890JESpvlIEv6NKA/2d6OCXU0O8172xNKaT2Pe++R9Rp92/iw2EoxhwzMRRTF4yBUUUmcm4ySk
S9bcEOCJow2WzQi2lXsGSB5Lp1Nb/Tgn/Pjke+I2FecJ+yamDIxfgolwdGOVE7/QtgDO3n9bHRUO
noRpGEAYyUNMmQRChfI33Zud0hko6QYnxcdrt/XFRrH6xZX5UZQ5Xiv/pJ4RS36Ao+BwVIIBFEjl
H/S6Z3bvORnaAavaMv1gl3eRyjkLmQdLGEUL6H0/Ybcqh6kaY8YZgD7nHeMPEMo26mcilIbcU2Wj
eAoZWUvJkCVQVwlwf9k4CV4C5VFfObbLLfu2vp8piGNxu0k4f1nagCdhB7VydeiY4UmQ6xLW95IJ
SHGDX90fkJEqngamkBCLsb7rQV8aZpj0vrwkv79bO6tQs7PEkq3n1N3+3pqvgybEGtIs2WF9WydY
uzH/SndV6R3qHmkD/uqlEn4bWDufspcL5K8NYCEb93/B8RC8OBEU7pL/7LqgFlukFlgRuPCsaBKR
bLX62VGWN7Lez832Y5Tmak2CVUgRVwUIpJKiZKbLYZkD+4CKlpOUo1DZo34SDrTV3pVxvs5/vbLk
04jhgBGVF1z4dv9dapkOqqRVW2xO7vp/OdXT13sjvvKgbuo7ytlWQQK39Go2PeXckxbeTdMfuTFC
hNk3Aw9lsP9rz95N8zl3PQ0IoQGm2sbxBRNfb6PTmBw3PrE6NFAdrHiuhbGPFUT84e11WJEAnTQk
VgKmQDTG08I0lE0HLnVx6ImNflysI196RMMXRjSj5n3zWZ2pUIDvppKiGND+0EkApH+t13Lg8Rm3
stlVvxQQwrBqpdWfExdzVcGpVL+lplYA8ycftNW89MSwjX2rHbK4EUKH5dqLxzXIXp3g3v7ttJnV
xWGrMgjig0ctPqgtgtQL5WavH7tBBOwv8i2IeI0CfNKe7t76YiIjbBAsRTCuLIrJ0q3yVFADgM35
oiMS908EKYFatcBE2mIaAwQwkOwg6UzTlLpQ/932hyJXSVBr4hJ6pW21yfQGAl5bSCf9B1u8NhGe
1C+NLIjbacliLrHFQb09BkyLYfOZOVjWwBJ/3jWT1fl3GpbDNMqYKTqYLVHaopf/PhgGHdyDUqZp
YBddoJiOAjDXF0Q4kS21yuqb/YgcijDx33S1XAKZGZFUhA/qoRjSXa1A7ol2R8RKZSZcKUyQ1Qbb
pLc89Ahj0oxjbK8OnL+KKvdp2iR5IIJYdyF9aPlywPqRFtQ04dg0bwhw4BExZi1BFDUsHlf6vYg9
HvgYhdyhCPTcoaM5ZB231AOc3GKCr+dDITmAL8BHPmiou7EDmcXTt3ZbwcdW7GI476tqpIyw283F
zbt4twq2yI7TBRAslbTWVXpPrUu0/O+K0CiN+5m87Syuv3Tnjwki+tH6PI5vuqUOb69PE7WA8EN9
BPsRxiPTZn0DV9EFi0vGlIVN6yohdVyYo5VUiF170SIVRddKe5a6KphVxmiMaqkqOcvNhklZ43P9
1N47wxuV4AI5/t1j4VAUyQclLi/cL782AaX4exahTMCsbgM9rw9HFqUgRrP9AUKJCrxGoBYEl5Az
wdd1OG7XxHAl1zc48VAFfjK6yHiVnU2Ie1Y9DXcx4jNU8i+ph3lD7k1J4exPur3Dq43Z3DGB/lju
Eis28lrXKbuj3b2TaNXvL1sAo9J1JQHSbVITcGhp6UMCqEO2OWcEMNuAqnp3JEHeF068f0vZi8eX
Em8y9nsAcO57jvSzBmSlgwGvxHGlqqBXwmceN9bLvQi9YubGXbkuP4pjugptXO7FmygS4Yc6+jAS
krpweeAV4ROA/KeEhjVpOrvseVc/m5a+e9FGglkcRTRrjKtEECFcZhUzwOsyeiPK+ZdA6o5j/Mvf
WmdFizHIzIOxSrmygaoOwLQTZ6KAst6OBlFin7pNQ5f1kHbCNmUvRq6zgi9GbU8uM0uz3yTLhK/D
DU6nuxOzl1QQ+MZL0OmjezxpIiwRu1qSMmY6rQ5UNp3u6tMcULXaQ8GvygF2zI/iDacweNfabBGe
LMWLttYhAaIifhBqLCXmZDqCV42UvF3aWmURtXsRB+u3XkZsfvtiJgiJCpf9ih2iF9hjHMBTTdh4
L/ygw5Gh8NhtGEERuDV3wmk8qc2cD4dUSt73uqz4q8lWp4hB/dRPGaRleis62b16j//bssblXogd
cF5ofVPesUp54nlEwUEZBdtmvlx1Mg0Kq/O53IJihCvCiAsKV1kOY/wpyWc7YblDYThur4A7cDzC
YgZbF7EJ1zp1ib2PrIERl/c+JA4QdgtPn2BNqlsTZxmOEKJActMWOI2rjzGv5x+LPO8w8N/+wXfb
yQEPr2r2iyXU0ojeFm/Rn9KmbFwzu6p1TU1x8B0qI05SrD28lzHgWm2dw8xideaZYLprh/TZEtSO
j/8+Cqw4+jhxaDJB7irHGycTZxVObt/rxX+Y43B6chMIOeZlASwlX3rpo4ZHLqM7kXfVriOmaaZ2
jQxCIYRKWbqB2xqHJCxR0t791gbSwqoHiUUgLHTjYcLOb5T20/0tGAtRM+CvMoFIT8CdMLAdb4Zt
rGjxtsCFn7sB77vCHfu5dLcjzzunbCxltp8Mlr0P3U/fy0yxpCiaiu7/9blvEetNCup40gOWndXc
rJtGR7lCNl9QIpAXYKq0wcXaXSPel2RNegdfBUnmj/+MgvQtPbevQNisN/qXdlyAfvAL6grrRAWL
eVNDwpxFAm8j+zE6nN2cClxMEaR9xP+P9wXPpCwY6TvXgqeeyAEtwjtq6XDECs3r+k/wtsP1jKn4
iiLvRWRKE70AcJrem07SV99ES4g345sF3jK5MX5MGiTRV3+Y60xg6bm8PMUh7K6d4/rWRVPT4O1v
4rp4qoSsq9I5SKodlXyHGl3K/xaa9FiqvJ9kk88TEOlJKpTTBuzhggf8rKYVH2vJWYFggNYdC0fr
H2fE3ggnsP1040yG5qCqyCzxHdibNfEXv+J9lpwX7dnNlMfxsVTFWwfTuVrRuv7TYkS22hsGBFqw
Ba+netH92fG4uAyFhBeP8KwQjxXFtXePDH3XGBiXgdpU4LZJzW/ukj4wy5/ZG+IakbZt7aUNhRD0
0GODbxfhU462gbIcX+Om7fsuRarGTryYISUDVt5+/EfISwRo8wpgMRKzv8If740I6sZLEKhIRG2g
LxjZRV70xh15kpKdnPLlse/+aBMHXzbNIFKTpfXTBqQcQLduoPKB3SdrC3gqMGCR02Ae6clmpsMD
LXHmQNn88PjE5njgnVN8yBG4fpFUU9F3QJZeywV2/Ab3DzHv1vg8uK3n/dWeb6h3NajyXKUZeEOX
qugogDXqS/9hwrX4H9s5BkPTbYG6GZanZQyYQtNz8R60hc8aY4SKiLcDogU98RSSYGqO6hoF66Fw
uqKJxsL7TSw5jgyXdSaB7OPkN9wUxDvwCR22IAJtVPz2WDXbyXoWGIQHBMUDPiCJWXZ93Evl/zL9
AKSyXbPnOsBCRLNrfSKn4rAJk/z9LIRmm8Po4jv/seDet+5bJbVV45F9scDTzBreqhiFtI6BLWuJ
Fhf4Jsn74mIQsbSzP+w8SCb65Nlso1wnTz+uH3xY+w+9+Hz0HNUhekcsijecNfdLfX6DqT5FSX2C
2gclTWErLOIs4LQ2YMHySky/QTpAZMmgxtrOPqojoDSi6R17+TZW/WIZmK8DgjWdEswh4lX0/d5S
XLTOSz88Lruqwnqf9cxlb4cFOcpgo4CMkat5lDLBAa7zYCEymxYnLSQBXOQQAFK/asUFyySjuuPF
llVHhMGSXrETW71nNl9eZrU8wrcXOFjEK3SJ2+0ZMIyQtF5Xn1ylOAJzY3jbGTaxiMpTh+dcfcUo
RG2YjMzWwQ3h/PBr7u3K5K7vFpS0OFH9KYMEa/HWeZaT5hTBE1t/6EcOicy3Efm7nSTWnfNyuYLA
jpGOS9qEwlevAy01bIK7ds0NhIda0Bcr6GhU4ToeICq+hJKE98cpGy7y4gyPQHiS9EPyOw/F+2AF
PGm/+kF+taMCHjGS9uEUZExe2I+SV0V8XrgSzt0EbfdUrgoo5DYAPWTDaeYy9AJcXynmYiA8WajT
tKPYu2MKTCbqy95bGXLhu0QKKiVfIZ6pk3vvK7Li3fKvUbsq/8YHIYPlnTiWJswxsPru12SS5agg
fUR+b2+YC2nGMHjtf5XrEDRZ07N8qZoO5w4fNLK0EWuapZxAS28KpMeHRy30XvwsGHYeH+dEikuB
wf1B1VXNjKmka5pACitS5dtTL1fQwBXnOXFhXDd6rSkGuWBsQKB98Dj4zZVntoL5wpw6wRdePDr8
1MHXyK9L1G2nh/m6mKlLUqD0IWMezqSbUmVnmAORfhM/bIfu7ioSnZlO3qYl5OIm4FUbp59jBHvt
nU5uRyPboocDdklzRvRVSb8VnUk8trW1q3bB36wzlr6G0gQIF8YbPhxK0ynD3KZ9fVUZvV4RxQHj
g+bFiao2SYc0EX7krfDr7v1msZ/3t0hR8Nk3kUrRlpIybwP2GcWiJCBFdLr3k++/GixoFcgzPDJu
y7A1JVSdNT5SLCUdMHhEWWE/3cU6fUHLsu9l+YxlmcwYq6AOkTdStX0xUPLO1v/gtWmkNYJL/VM6
XkSAfISNiGsg9ZhOGUYfwUbdSYz2ZQHnNiI5xgrxKbUV9Kkk8RjOK+O8aftfeR9wU+RkzED/fUmp
x+OfHHtqAONot7Zs6sEyp7R2J+CkvCq9NsHc3mfjQipOWSZxA3b56ICNDn1buEEaZwGJjTDomXS6
WgAtq7Q64LugdELBNDKCj3e0XoWmGLZwhG7lZPgdA/i6MRK51WaogNspkJ//Rbbd/8oujPX37JMh
pvibnny0VXhetEq2wG8U3uW2+4o/enoskw1PsUA9rCphu/28JIJ/STsQcmzGzR8C7djPdz9CyeNm
F3HN4rxYUFuX4esyuwQnYx/7J0iSuIEh1j1cNOJkGxooW9mTAKloEnAxeX2ue+caExYVkozebWp2
w7NscKffKVmsWvApciK+Oyt2MgQzIj8yJuDZd5YzbK6p0wsC/DxW4nJ9fepmPuh9dIAk+xIiRD2D
xeBQrjT7zETirQKDbRVEw0etf9+yvcplwJThweMn29enNbYv0pdt3LT7sAjfWen9U57vNlSymLwF
mD/x7ho77Wz6nNuNohlGxTHzW6sEGPb44ECDhjuVkQ+gDJ4CT9wPYu+6OEZp3Z3HPOG1bwNmdM9q
RUEcyOEQQ2leXuAADGbRPknhKB9Mttw+ked3W+eMAnmx5UKsPSbWXHN192FYV8lXvmGnsHHTnikb
2obuHryfPBZV4vs5RCeqaUpmsGkAlb6Mz6JRqC1lg+lSpRKVe+y47OhzKhWvIHLB531AIsbqomgx
+4C+bFRmybZUJSxzluVr1+VDHsGgPns2PeX8rzD6U1Ooi8zHgzSgxEbToElpfroKrcJ/IsG88Xi1
brIgO6hi6V6EvcqICn3uvf/TIIKStlD8KTNdBHXJoMRyWPX6ec5MHN5mL7QPd1cIzvKRgqDeL4RF
jByh3t3D5/jtTqa0v2twoHU5qiSgE8cnJKc6ggsWw7wvNHGfAy82ruUjn8sLtGbG7HWaoGEEVDYo
8JpEYClpoLJCFFM8tP1s00i32YAI7QqozvvbVOsajungdcCFPByTwNPU7EPApe0qkM2P9vYlQVbd
MCvaOw+J7A5wgmLxhry/JojHCqnLJvPqBO+Hec1shvj7zfl9NOagmUaNUU/sPrdTgx+txOCOP00h
4QaKA2M480QnnxiLA3B2dUd/nMd1RelAyS8g2tLySslS4PDfYi4Xr5pTlT9Hz1hiHRc9JaDHQs+l
6qTsF2EaKiq8OZ+sWTmmbMccYlLXE2aSUcUq4Dfwt/aYGk8vVItGNUBqmOmPLXTf9Z3pkgF9gNdE
n0qUttR09HIPzDuX8V6lXdW35H4HFKl4pTUl5VxDLhgtDiAsTBmxqaWobj0LKCYBUxqQykMspZZ6
m2NEOPRmT5JO4MvgiYbYEn8R2tgjlDRihvIYmr0C6tffqw2YgyPlL6oKeo12qms4kLMM5exsv/ic
ydQ+UjXqV/YDiXAawTM/lq9CBovq4AACoPeGB/R1kMpSxzMswGDKn78Lm5QhbTLXE4TLVcttfQ6H
YUB1QrTKhAgV4hP54EreEAai8G8kBFrOxwTHM/k9fBjVpiw8Qt6BfCXNvPLGhj7df/VOQkIrFYX6
KaJxXbWawpW+/2KLXrttXMSFGfMrIFLMz4nLSv4MDhcE2+YitE0u5fXqnOnU/LZKEpDjwTrmPRh4
kSqQib36unYdOa5UolUXLFC2Fw3lVKgzVE2O7+vy7ujb/K9xJ8SFs4rIIlVQn1Njpvkr7h49K9GH
hT1Fp41IN8yevCUR5J2zNMbKIR8STE45pBnhkqsc23xmOBgy/fy5ydcb5axFPqKRoHfTgSBz2ayN
YEWwVb6ApvlcRlBGP3RsEmtrSvL+2DdDRnPgH53f9tKSHFrikSjQIryg5WtwMqX06sJWIuB885Uj
hhHXJY400N/IVM3MS73sZ2ht8k6txXbkW5+L3+ae6sZhTEgPhcRKiC3Bvyt9KtOHIr/P+SNWNYAN
ZWk51Zwug3DN7NmymKzMtMGv885PxpOVEN3le8WUHJnNNByPIR2zgtR03orGjDcrkhEK4iCqMhzV
qrH1BEQ8yOAuYxTekYvPXv1vd3aLKROPJqqcxIwUODqdRI4gc2WbIumTtxjP4fX8U9bHzlRhpbtQ
cHBcVHaURGxexOIxx53ipo5ERScRU6wn1IF94V65IpfjrDMHg4rXF1/W5g6t280dDSZP/RMI5iXd
jt37/ar6+l7Nnukbpl4YtC8dSQUS80iFpaU/0JYsizoQkYeXdW1ltvZBRKstzqgOGBn5Cc8HZaY5
jEm+GGDLV+2VKs7cg3Q4cTQyc43RSjDxj9rHIh/zrwHuWrvUcKTIDOr7JymqXNs1TcHnTdy76EK5
QLbRJIpZKL9pciO8WIMwYclknTYciCi0w+JLEoysfPViq3YLwwUvN7UKDq5UvU/87Nks5TMlN4t/
OgnR3XmnCQj+EL3ha9kPEsDsfScQyv/LnH7twnv/E9buwGeTgKMDVMpCcm5wA4w6erdVUbLR0fnV
tt6rY9HSBqSNE8pY1Qu33Nkro/xX7BL1Ej5AbVBOR0E9dJuNI6lAChS27gnrhc8SkbhK4OH1KKsz
ZSb+Fg4HbImgjlM7LNXml4sVEmpC3m3SdFwsFv0Lh1DbdKmo8a6uaeHO1qd05zzgNpo6REWNMd63
fVJ706t5sM41NSyAHxvSw3a6n9dMorxq/XXDtx4MvBbtypVC+/ErggBFv8JEij+cDFQylaoj9cjR
nKwbqIpFMe98o7tWaPeNMNgxN/756m+nJGsT66iCjHwAdJqLTAOzxrzEO3ukgw3k300oNsAXUQ5k
AuIm30N83e/qih6CrUMYF+VOONgP+INZyLNaISH0dLqFRDRfLkJWqPr5l5t4T/KHr4b8DA0PwJd5
ZZ2ROWEuUKf2mz0ZZv2TRLHLgv1hgB8ItDBL/BR1mW8LyCBr4uWXhyvZcKb9/67LJTl4RDUhVkN6
wkSJokcdXdZv6VLnTBrGF2vfKo5me36Lg84mFd3Sm2f8gxdAUxaugpBD3jK/RbR1r4MftTE8TbYL
Q1zjMUVgHcupya+zAC4y0jjFu9+2IUUvTrCeVSAJiP8CQngLgAruKIrssc7StRM/Csf8vTIUgoIW
eVPF+gwTG+nPzgXOPWWfYpMX0zUGVfAUsdT4bOPW/YCmd8Jg1BeOMPkfq6nZxRWLyMG2ESRkv9IU
DchAmlq7Ud7VVNHiLJUle8L9TLRsyNi2hEET6N5TLMmLGbeToY06zgIg8PMe5nhBfn0vB712Y9Jq
nKkXiU8oyMIFKHVGxZSwY/vgHS/1M6o9D49KjBubSsP4CfofeygOAgQmqDflGzd21r0Ga9txnJYh
1BD2FLgXtR6seycOe5cevK2mc+PXXm2DJnkxsWkgcJzozf+PwOETsQMY4pgrWaCnWuSxoaHx6/Zz
yQcgEoRE0UmMv/hlQnlrFQvfiVQTdUMsN15a35yuFINYoG4ETx0PdSoRXCOi5imtsBfdg9ky5m2T
9KaBMcz+hV6AL/w4lXe09PPbWaBrrediljzSKwCcdV/edkSL3MyJZBhHknl+YwxUBqAqdwBmT6sH
mHehjQeOWUL0DqbSW45oiYWj37Wqs3Yo3eDXPkbRtGYdyTFsarl/pZDTGeQwZAkqJh+pYpn46Fhu
0szGSIQWebbwATbS4xarJsdSfObieUMA10TFRrQeUxt0m8wJdH5e0Kzwtjslbp95+GY+2bAxKhpk
U9TIyygCzwQ1W1wNgggF0q5lY9v9XkSFslU3j/gzu+8k78eKlEDSOn6S8Vs2awuS2lDZcZURqDj5
eS/B5LYRkQSSDDWCpBdoKfmkhlj+ZRmNJzS0V9JAOsQZp8GMl9OdK0ikZ7tLntOjBsEIOsC4+0rm
DtXdFyfIWuk2TWBeqzSlYZcVihxi6HQ1F/9Zwc2/ZTZFraXWT3Qh3Gkjyf9mJqEjU71NPGgYA5bH
vuJ3r+mLFiHdoe02YeIXjN36McZLyCWwLupbp66kZdPb0p+ObtIx1WQPgvVEjJE4yP7NaaGFGijg
IdcXSKLfRi08r9sqOD144DdyzeFphx/o13SXXlPjrGtINpgc7p7YIPh0iOBgy/zM/LP3tMoD1NDU
VersWWwyLj9K+9mdbcCSywPLZniO6C+LJlaWwgh4rcraorN0SmvoxXHhQz84cl+l8sVc/ofLKoBm
/lVBxt90sF36Sr3efK/5r56pUrO9g16GoeoOOAC4SAGQD/1UAyXhNwB6omAOiZBpk6X/wfWuCdCh
Wcy/V7rvFDQhAmSw35Rx7q8UGt/boT3r4kSDprAXsQjKp+ysXFLX2IaCQetUQHuu+NpdNtrBMWdT
HEMVW3xW7nctG2tb7ZIGFRvLLN+5HvTa4viVGWbj8ndt0gKZWXxEKGJm5cgfNxvL4EKZtXKyETep
aikIE5DVrKyHvXEhQIv1ORUFIQtY5EleOSGqzZzI8QdBj6xjfDEp5vg24fqrl75bnG79MoVL1RnR
RFCk+qNH9EDzPFxcF+7T2ntbFGeYVCwOVu7i/hizT0pjWey2+dRTl9JAlz171/NqR9fM7M6z6TDy
jsMzEFyQUHbydDkv8MdVE56ISWbeuQpdC+GtueWsrrFX8eNKPxqWZVKLNjT9N9mW3wpgFW8moSmK
VebEuAQLgIPDmVw62IYCeMk7oEZXO0PEQ7gU8t4zal6qiLJaUMi7o56EmHSINGyxBHKkkKXeL2V5
oYuR0nQrWEzwdZY5RS5KPBEK8ypnT9A/VQ6lEJ4alFcR2W7upuw1y/VFx+hh6j69jSeQbGO+cXuI
0sqL07IH+91V1AKth7n7zXRGiC/r55BAM5r9GS6HJm0gOUFJnuerY/+6MUh/6dAcvGKJpah4IM4t
X0OhpOb0QEnqfawPfAiRJpDKILAqdVtd84lJ7nBWXOXigjMnTygT4vJ8DIDLqTZsKXghKu5OFCbO
dqBWvTU1rj9p7RKUKBDoxfUuYhikXuzDOB5dgyRCSO8HFpxGskRo4gEcLcYf8qaSd8uJZ/1BP17F
hnJRpiAIzQYbFj3MWFJAD0wgtUxw+ZW/mvrFwvte98zbazud01fa6oU0hgXIgZMAqdN5+JBg65sm
3zccevE20Aaw9henocYplvnYWYWjS00dCtFdBksj0pDTFL1RNmAXfaqqLLskVSfVA9LLK05XYBQZ
5FkVkNYNpSvgS87cBg6bSOdoCs73mxCERiUw4qFH7c5jdi/nZQ+crAii7HFuYAdzZx6DUftH8Bow
pvDItgCU1hT8F/4SwMv2tRsGsA9HWPVvmLBvyxiwCZZEBqOxSDXah8RZxKMXHZUmbwxW5d2IHVNk
OnwaEMyOU0wUoGTiB5Q0O8zSfGluyXiB0jf66SJPaTlbvGPf23WabFLDKdVNdFKq55imtSvVSybL
trbWTUbMKsrKSm9HVE0N4FcuWn6/XafhqRuOekuRR0TlIUr4c0M1RrmXIDF7WmybPJW2em6sQEun
zKXkoU7z+u/zjyI2dNP95vRvEZauC40nGd4DI+6lEpkttJoVG9ZPgB/UFfMDP3tTcY2PD3Y/sweH
qsN75vYB+Xjsz/mA71B5GerSogc6ClkPjWoElUqtoG8oWnb+dnWoS2UdtZ+5bEi3zIhPQILl49mv
B/dS+BeW6KFgGq058Gn6nfNrVaQ8jLxcUJ5xb3dSWTS3KGCgf1VOxUeUraM3ZvMPZ9by0aQY3dnD
lc6kUDO5yEknXhMlnvQsW5fpreKdpBz7+8zrt3ixyaRujVYq5u1jtXBwKpw1arAajI89Q8h4u1Vk
0Uc61Wb4vF086Qu2nSgn6yVBIQDQBjSl7gB3zfcOEFuFBt0q6RHtcCuuSibxCYI4Zp1uLwGL7l8i
0R84rZMoVRnuqXzdtpmiXiGMhGMEpCwq6BjMOgr9OYFEb+W1WdMOY/TDNsOmu0kV5MwEryinPJ1X
dGeg1Ed5HLI4/mkh3QTUEy2/vNEL98Q2IJx7upZ8zXuJwPIOoQqgKfCtab4OB03KHvt5JBuRMrbU
61BWxJP9TrHmDz5gw2UfVM4bjAq6snrpZUh3e/EHeUShnir8VABBa2SKfYCZP9msVqZN85bzN8ju
j1NcJFBrDUxc9ZkPfCRxVw2St2uOC3YfunefqqFLRcMnZdWkMr2teUZOyNIDYAE8Hi7wcmN2SIAx
K6AYC2WvjKbsmwx4/AgQjwANcQfjD52/PKBEbGzUgYWENMqo185m54SQ4/iSL9rL7gSN2Si4sfIt
1WcLHKX1FwPnZIhyKR+CD4Kpa3wvKb8J8pwJbhP/GzmtBhx30E+usta6rEHXlhZT5JjNFLRAMS7F
s0alx4n1NRYEnUTBY5c6wfUPzU1albv3zsmeta1w0Xuz+pDad0SSYdmdb66bOj/lf3WRH5n7xK2Z
xcIlZOkMAjKs7/usa3IGlKyO5u2AgMTSqW2cr9CtKwUVN018XPw/vjLqUtaWGYYIBUQz+mn1QqNc
1H/uGPsLvPd+HQwODmXd5tNWkHdqXFA1sIsyTjb6ZzqVEr42Ph7yl85yaRSd8WsHxg6wqUYEc9IQ
hRzm+oOTvOcm17JN1ALHn5JIsRIJWyuWS61pLt4nAMqud2TpUYFV3NBe3xl8qM0kLVeO8E1Kncz/
kmUBkbRYXcXDj45ngdw51tSWee7NOVjzU+qy36ch2q45cDSvEtduBVZGgRdZkdoIk937/OGA9ZE2
hfQ4tl0dGKOk4eg5eOcxhweJtD0BIsMSt0rwdd0GTpL6p/qG/XsmJ7bvj+EmN1nzXvIsJQNNr1xM
TcGC50viXHjiLqL+qaLGl2o4I/4MfdR1aWkAVlfb3TENqaJrseidncy7f09f2Z9z9Hr1UPGaaKHC
GN4sMJXFA05JFvjG8AA8OXfpIQHdwDi1QoWq8yzDnL+HRzJpRQti7PR88YPNMNbyd+sEVFLI2ZuB
EMWUKl57Ebia2MGStx+2yjGEjxWWRwf+fCFPLOIf9qcwVpVB/6AJ+4otljtB/ltDgtl6lejKfdTG
wZu8EDlqfsS3gCdrhoBZOi7mxsnSDnXbwXUNqnBw3yEHfFq/lTqvjHNgEMlk6fv4YGt52ayY3TOy
m+ezEMwcfXfKnbXeQy6bAFD2xhSZF0o5nzYJT5DPifdtByEmtY05ukqNblX69hogY1ZrJKx03LxB
h0BUGMW3psfBUmDUw9RWC7FJlD0svjCPjwbV4eiwU/9UnRM0W4LDH/GUVbflSzkQePT8NOjXNhp6
ZDsLhRFq8c74Arg0iRxUxqvbsznFzSwVOc1mQdmDIoI0Nr/oD2HBC7rKD6i4ZIdGq0YNMlG7pf99
AeT2TIXMIKb8wwUbA7FUUrK8D+UbtwQ5Nfm+J9u8Nr802Im51UX3l5/NOFvDK9/9eLZqvPTBqPLy
vwRngufyV+CNxWvwRkjRMg5UI6gW/sykOhoBn1aRRH4q7B4F2WJhPL8rQMxqIt43ZWylxQJqOum4
HBBtXhI9megPAgaVQDuykuNDdm6I+kgyxiEl8UL9iuWiGXUf2JodwUbYdFEcJ/Huk2XrVFQz38ET
wf53zQFbi3vuA/vwimMfae6fiXn2U6svjV6ypKQFCC/BHGfMb/8Me8GNXHFqw1QZ88/yuuwZlH1J
QfPl1IZbZhd3J6RI/mcvOwepA9Bwj7dye59/kqYmH/N63hwrVryUv78HTC07AdcCUNQd9ykstvjH
3GafekpLpyAKdjJGSgI6jwnFOULjd4ZIZPhBLc6j37Q1sBBP9x0aP0/fZtZELZ3QXVm7F58KdHcH
ci3dv6YnSb+2Xso0Eg5OGdxaIjbq4Ak295+RJrFOZXY9ECrKTKoLVvXYrLOmLlnW2/meHqTYiKfI
r4wAkdr0cMZOXXXupZh+n1Jphr1JcfvKrAJWpPswTgXjv3UEJacj0cZhJ7Sp8GyZOeAZTuL3Y56X
ulzUKufK6+k5hWZEaXq33Ren4g535PXJj2bve1bITqTdm0HqL6DBCOoHNtplzNWL9lyv4PiQE/xE
QB9QZNSA9tjDPywPCR1HyDuT6k40hQl0zjy+IeB7JOf+xTm4/34F7qXZQJSryp3baCzSkl5gyvUU
XuA4hZQCE4WpC3vwiMqVLpLyQ3H/PcG+YOR4q4TUZ9FlPjUL12hI6wunfEMzzAgzGv+SNS5PXsE1
Ns4aYMKCijPHOWLI8teldqHc/OnfjEK+sP/1HAcTP46D3su0CEnvQxmU8ZN6f4z3ahEzFasrK3dG
JuE/ZGYieU9auCsyVqwEUR70jO0Rs8UTsuSiZBnFcq8XU+nxzbVxlW1bu1er4pEDQY2FGJDbkHWO
s6bEUh4HFQ4ZxhSXSLgCXEUTZkmTt+L5gri96T7aEU/+NsT0miUAT1gppUeMIskIXmgAqWOZqbE+
QwTVxKIPuzB2/qzC3nIpBZ+bvA2z0mH7ItR58pXTyRiZTfKlXStN+GjDs8WYd+F6EX6uxjAQqBCM
7TbOgR1Vdleb3/oqA9lCmkPd6la+anVIbJVIx7wdR5/DWphnLCoCwD11KE0opvzqgMVlhwtvu4zC
stQDHgu6ZaoKyOpYbWzLiJAOG4KevNOEtUA9Dgv8wb/OWSzdy5FjQfJwDUdd9C78PGcG9JWySTHh
dy2arAjPLeV/ZIsy1NA5E9loEp3cX8te48QytMrOcCK9j00UbVbVfTfqIy8lxLY0Ee0L9hP8OZRZ
uaefHceN130AHYSy/8XthMxK9AhsXlmKDzHCK+launzZltdE1tGedscho3Q1eTBrn+fSXoZyP8kY
FvZhNo+En2QXfPgG76/tbEp5IpVOYLkBvCHFF6Eh+bRniH9nvHfIbKWO8HA1vY5K1jM2+OWw/ZmH
aIeALctg//VfWUuRbbQKd6MydwGPqkQl6EhIULGtc1pJngncyTFJTP0XLby4PP4P0wJQeORnOVEZ
+QEnGCnOoRWVa6+sHqux4em+MwJW33CcyBgsF9msKui9zTKEHGf/Ryd7mtsUotTCabdw/E/NLbuQ
fBewm9uMAFvfDsGCoziMNySKUxA+cqitJe3d62jItdX9ZKs2/bInzj2KeUsl0ZHFKPTL6oihxaBn
SQwkciVkxfAsfkbHm96UN8FH/VPWKI6LfOdmhlQLW9xSehP8eMtcWqTIS/Kg+Yi5glfetWgY9mPH
6R1W3wHT2nyYr4Uj7tsd63k3OVdEnQnC7/2FIxhFK/5tZ+13IMtjjhAvYN9IW1MA4hsLggkyM8fH
A4MEwBgLI+2ng2fKcyiPlE4cXWsTPV6AsZyyJdjB6Z43KNY3MEdMDs+qWNwfmeZCkj1I42ivRx8n
z1yFe6JHE3dUCa6z08jA1RBJUusJg8e0y86k/cTYsZJIWkx3D7qpJmQC7YxIcw1lBGc2lbBMNfLy
kjio9xcvpr/wMiXdQ0sWg/XW56H+Gi48BBAANIKC+7vPhS89bkhU5ULZ5nSaOqlc44fxBau2L/TX
vNlV8uaKPnZ+WYH48oT0M73788kFiWWZMvXPbh6C8hatcE24nB9pgY+t6YvCoWbMMtpsbpWbueXN
CpJOcWYh2cTzu6BwZY0Oky2ePrH0QN34r1h/0wHApsb88aPRLRQxsKkqvacVMJAHR7RKRP6sDkHq
U5K+Nx0URK8t80t7dDoHD9nHL0P5QLm4SrChjlxQfkQhUuOG3WMpyeI6Qgqt1skKAi6KReiur018
2I64GVMTwdWcBB9xXocG5TaNrbBaaGc2EU6ffjOD1bQvIO8rfTjyDPmsZKXR6bnap5dvfnhgv5Ll
ie/H2juUShxQLSutLpDEl0D61I5dGtoi/dsLkupu/WeBmJ4Dd8WkM8F4kadCL/eT0P+pFyT3khLr
QEMGNaXWzV7XSZi6CbT1I+WGVKTG6eyCVbsRBxJ7q3+jEZ/ZWjmlIJvK1C1l9kyGc/qv7w2C09Tf
vg8UbrWgx6qbfg2M45Hgg+fCFJTq1nYbHsmnZHx7y3+0p90AMXJ7+Tha/OWnveQMqZFXrt/8CBjU
tg10Mnp6aiakZd2BPGvh6160o/JUWojUbWL6dGhhlU3sjMKrwJwT284bL41QFT4Fx8CE6MdwPvoB
poSWm8/3ojFJNCCkcXwEaTpq1zORoBvmjZtvItqFqez1D3B6G7bbrjurGkBQ4JXkrHgJYNJawHbB
zweh4i+5BUrJcT911w9uAShM30PBc8pBwZSzdk/9r2cc7+Tjgo6CM4oTIOcUA6NBRLsib5uos71I
SQpkPAIeeYzeDu1zyKeO/JYPD1i4MrqXoGSj/HcQSXKJMPrzXFJidEE96/Ln1usr3lbQhA3dE1TY
bBoOhoBA0L3RZhKdQmpHxKhETxMj8W7ymZYjWtP+pqDYqagoyhgFO49hnOBK8HkQshe3w1K6OgtV
LiwgIvaOarZfUiyGNj8E5kiIe0W1unDbpb4yYcuI5daCR2ucNxyIE0irOHCyYiEpehClRcJ9rxtI
X0GfukE9g55NJqxAEKvT0BZUtud8IlvcbcvR7/3OopFefLuOy1c7TDyXDZIPYxiw9CZIwLKaBKpC
MLRJzLIHXg6UGW9otn2N3o/FZeGcqa2Ya7pzyF5RbyhQhNUh2wOCGSZi119FOIULwjuLquiv4J20
A44m7kyg012MoNu7aP9e/M3CMmU78FJBYoyiKDCBcCfE42/QTTYkxrIwhgLvL9nD+N/ymvGtsSHg
LtvkKBSsl2CDS0D+CJ9XQAaGb0kmxujzLS/q9/ISWi6/d+gRhIKs0SMug3rfmAGu5A3BGzc4pE5E
QBIEeTmj1lGEgIQIblrrGd7XqmTSeiQhtdHz8/3NvOqE5yr6vSB6do4V19IZapcohJpdinzsNWO0
qaaaEb8RjE7E8FavZ1Q+JVjdOj6tdJj/KZNnoVymUQzSyjHdOag+btwNcAbxqWouvmKL1/jRfT5V
B9sPZCm/miZI0SKGeRx1UVwMXalshqjkdizhbkNc4xlhQtuCB+nRhK7I6tvVlVNd+pTzS7DQvXum
4avqFhJPrYLg/KjbCPzxzxz1Mbwt3EfpxHzQZldgg3OBC+LRcqUgJrXFyucBM/xJGZAM4pjD34Xu
Ut9dxQs2Ps1RonjUTIxLTPX8ViA1feWk5AuJIyvV88GSUkF41nmQ68Oui6pKRem7MoWjKvmVDg+f
cP+zz/ddMnHp2BB3Lj+UbJ+JUXxnEOAwgZDsgH50x0AA4VLrCOjVESikQLvAMYk2h88jWw1m+s68
7ebRXB3sU6ib2GOyLGfW87eWqPgWkTkhq3oVvWBUPlDcezy2LYKKgzY//pts+KUtJl6PjjJ7l8E2
iTie/px1lkR+PogXK1nfO3S8pPhHN0VI/XfYMQCyKL9GmiDRteQWi1h1QOLNIkR746C5sWFUZOSQ
ktD7b0G5k7USWmctGp0eEvYUQ2tr6U+0NC0/3AniCCS0vIEIW/is+nscz97Cli4Adfij+SSIsAzU
UyPBIB4ygJi3rPLODoI1z042IZTBCkoZPA2yknjDfjszZnJNk9JzG5/TGZoMh7upYXuTS16fl7EX
BoebjWXwbqSYhyhdQ+P5tZ6i2RDm+Q5F3+jZNAaGgdYNR2s6ZX4JJXo2amPXCj7R0sRcU3lXEkMa
wj1X1hc7krBs6kxcAbbJfN6ykIdjgLyBPT4x2OC4GfKJ/5fIo/Kep8PvUwJLsnfULkSa6O8zeHOu
90pqtg7s+d54gFttCLJedTXqOVu3A4IZJDtMYoTBZEgRBGwad657SARB+LWIrVw5NM4Ws6yQAvHc
TqGsU88eaLKJVmN/5+chzgZNdSai5vLSS2+3t8+hBGE/BOkCOb7xtKRNfHoWikMZdL1AJtJAaJ+i
SP70s7qn+Z1jB+L4mJIDhbcPG8pRr6pb3oXQ5LClKl/EFn5oOssyftE768NxY6bWgAogJKeBorZC
AE9ljziaNyoHI2KHoBr92uOgWLx+VKwvyhFfEY+K83zERM5NuUqVP843GkKv7DO4nVfaoIY5oaks
PtfBlSVr8VBigvZOgo4sKLdgOK7QdixsZdndHug+NwUSrRpgDTKvREoKqb1f7dDnhJ+QOnUgj0Of
8/obVBvpEBs3TQYT8Ttr3B5dkuobT/W1C9TRA5QmoFaH6lsh2/31RTlqQkUSWNCEWy6tm4VbcD4d
yH3bwMHhkpGcriSDSo3yPYcF8wswS7AOgzDtAvLDJ23pxMLDLJr/c/4yd4+mb4JYYFpee0lkUY19
t0/7hNMI/kDfa/KDYyIAH6FbIoGz+0WPp+ZgekxSPmh4nuH8AqltGjypJM1waCwqBY7w0pMFL1HD
9cxWggCo6Vf8Jt6jk8649QbS/xZJfioIu34IW5dwUZPew+6+s2R81M9Ont9/KszqZvW0BUZ0VRE4
kPqItfYML+CR8NXORSAP08UNXxOVWN5/d01HezjKk7CDSzuNdT+mqM3qE0i/RneaN0ONVQWbKSFH
goolefGDKU8oESKwDWiENAtiK+Bv8glqjDMHnxmgEHFMdJsAtO72jlLUrYwj/NP35H6QrGWWE8si
svOyvUq3UFKxtetdoit/YysC+UKqafXrNO3hmD05ZVz4NsJaI6CU8z0rSs15u8Ki2rrfBM8BFfGe
gVxVgpN8Mj1rh1dPDvv0MVTcnUblfoCVrUCohRHbKQ5CqCXrCnyNrQkz4X3K9iyklS13GnaeiRWn
aGq/yDnPJEDmNP6P5Ib0mwdJ0mVMjXcKqxkez4iCAIORZw7e6jrlZjCt0qqBuLc+xnbxaMRGkOWN
DJRBO7P1LMF7KDASKMj+8NSdMSep+WRG9iarTZs+/CGpBdHrDI0N/ORcvGvu/8Or+a3mCAWMPVdn
hqXeT4NJGZGnqC9oMEouJ0qaHvlc2QWln+hTijpYv1fRXiAVr45TZG9M9jzRdegvuXMWguIG86+y
ZZ063JGLlFZG1mL5KuZcdrirFGOjwe+QLXRnH1JGHpfmN9vriT2lxbvVbbB66Gn9UVwfaaxcQP1d
sjnzamQfxX913zd/f32nULtsAe/yNFp2jSWGeKJKjCJuApahbCFJoJ2wj0ubMGuEAWUYUthhge/q
V+dJn3YjxC/iWc08Yo2HzaRFti8rQx2+o1UpO+llqcx+riF7rpikCGy0Yi6v6v/B5inAFpIAxSFp
NU22HQFSGINlXaIdY54HJedQoSGa+PGyHHeNZ77fugnPVbL56SrctgE8RC8PJZBMR5nkRnTpnp6o
DISHuNV64QEEElw9RweXAn4qcU6okGKv4Tz73lr82RAA80ijhCLDkKtgRoJ1jztHbb5f9nLqzoqQ
2L7kkGpsI9osQcLh1z4M3im2vTHtgTaV2775V0aA+rcHlaXERh5jh/4Otrj99U4B98+VvE0XyLeZ
XFB8MBlEPB43blW5PxeGYuKcMp0foSqG1b20sH0wsUulyCUzT6DqDF1M+d9A4L3KWD3axCLnoz+G
E42niShpd2NvIHT+gPU3fPVnkw2WpwPnagHNZv/FOfiS4roZpyaMcaXi5WyNmRA3J8B7ficzVNYp
nWWB21R5bIQRgUyaalP3RmY4xEVyKsIxUJbMY4TXR3rhhf6TXzb2oFbRMQ3WX5c0gM08h8eO/6Nv
IMt/YuBXKjj0gQl0WOl2FtMveBWmuvdA1QdLvBwCda5gs6xTz5r7OSq93HKvjc01wG8tExdS95uW
Uut7YwHy70snKg8PXz7NkTt6r7zxTNAikY6h2GythNdWkn+uewMtAhdruLZcTWuOWUn/4C5Ip9J/
twaCByDdzxQyuNreZPEhfdzPQTsZH8fhS4fHtuwmLAZhtWd3kDnhh5lfvNtPO03nXYsj11DqsF+c
uPsND1vv0gPnWfFdVMvDK0ianV2BBLqFCuE1oR6W4H/DAioPrWNnl12gSQho9Q555/wZ+7eBuw15
EgjrJGuTVCn8k3y86YToaQSiIpNpg2a+sx5hMlJACE4RVMm/Cz4vd1dyyJbOZ0HgdOxlpX3uBbWx
BbVCjfRyPry0PbrqvVbQD+Nn2QWcUJOadWG80Na5gJZS0Fc/b/GszU6ZZrYMNsd7Kx03OyHuFxlb
j96hYe2bbqGsokJ/s16yn2EbgftI11/4IGjodcugsRU0BQocGckEyz2EuXIzY5KmH/2E1DL6reqX
vfS6uy5f4PtI8DXxsNC+wMhAUMq4l4DdOXzQvSTuU/f1Tb3QFGE0pNJ/OYHoQmdxJH2YTiwmj63d
9O1vCe8GWG3WqtUG/hB5oBRAiiQYbtrIoQVeb9AleuXrGJX090x6EMMbK4wkp1LABhePCs7LTgGn
bYlE0rGxN58zGmLHcyR8DslNtoztiukzyMi2dR4okOL+xt1cF4iv0SwDjfhem7GJA+suzIspFGd7
ImmmPqP5uPgk8JMOmYy5GrqeLi402RPiRuqMbA8RiRCOsT7WwGr04RAZKeu2/6azt2VQsn/1qr1d
vO1dAwK9aL2S3KQ4E5II+i6afO5Nsf0aJ7mCi4wIITtpcATmve389pfM8ST8PEmUVQAeW7KfP5CG
lRobXVQyO4n8n8qmnKNMfyfFaqSfPXIL1JXgsOgyqtLZOP6Lo+SbsMT9chyjWR7crDhO2RoTGNKC
MEiybjCOzFklVZC1CoBeMaq4OXSgnQmPPwn9k0P4Kq9O58rBH5G35ljVhWDQsie1wsueOs21zKFq
Wu51dUDroeqWtvVMwf7mXK4jZIlOXe3XVd89R1YFJuPZ1UV0oncBtK56WxhWsrOH57kYnwCb6scf
INp41si/qaLpg1CfLlNWp3kpKeDRtPbnS6pt4DiJzr7wNQt6xJQQiyYfrIX/38LVQG6S3z3EMeK/
K/4VhgrBrm3whuWHnMVuebIMWL9eGgWmk4qfguwKaoJQEbtZO0/iuEJ1WOi7nPx/IjLZ/rxF6mlQ
c0hWNcWtu5Zu2RPPCuhywBhiAyPa8RLR9K14Qq8OA6MbXv/H2cizSpilWBFZ5KozHvaPsT1j4TMG
wSbH8nJ/ESRmKc2vm1rvRce9Fn5YBxg+PVIkqCYogs1HwtMpIwFeoUQJukbLbJqMBs5C1J+u3Gw8
sgRebRFcxEqgcjtq+4yjHa5YWuz0ZyVl8xUyPylNZLOVEMbH6Vzwkm8UnVKA7Yc7uvK3QPGqZ9tm
gu27Qh7mT/wFnw0ZUYSUoy+WogfoEeP+KYsp23eCYJy8M80QBgh1rIfX4Qrj6SrNVDkmhlZ2ECG3
yBpqh7N9wikSMJ3H4itplxaflGB2tNXuGdvLyjsiEx+f5XbtCdoI6CJ1yhFCmE4PZ4e1hXOqB/3I
2wugKICIML9waeIorkipnnODlF+Q0zxjWQixNejblU8W4d0etUDxcOVlJeBVwKsLTSeXRYNOG1S9
GMfPPRRZsL/NNWn8/VqBZq84OP2I3lfZYoV5OQd9FCEOLTZhqiOlN2io9AgnUDvCFeJod4NiH9/8
QAwbqu3yopit72P2/kIOasiaZJFzPBExCtLDX3yqLFFTxuMqlqaG2rTPxW/+VRTI3OYmn+2pbyvU
hgFkAtQcIo8wdRNCTtZljjVvU+Dkj8p9RwSFy/2rCj4gHQHh8khK124fZZp4QRWnV+Du0+K1WNZd
+i90sHz8A5BbjhAfKN81M5o3MLOmRo/4xjsdH2Ujie/pC0aQkDE5UbvrCA+RSn5BvhcJzIx313B2
LYMl0J/HvdlkQwvLThTiGaPemnpmxgklmOnzmI9Hf1KXh6i9S9tkGcZARIPKGUvxVOEJma91a+MV
ZXJrk4HYOUbYUJPeTD7tEp33Lv3QuNji9CKx1EoeIy2fiqAnViZtqyrvdLeglRpTLDFxx43e2ige
ajAs5YjnaOnnTZ3j9418JzTgHGfe9863l1x+1AE1BNErOPkF8Hh4HDHMH3iS2t9Z/KERKjd+n+m7
LL8KFSX3EcWKbWILt0URLuIFzvWb56nCQOC9S3v6nv4TpTtyq0PsIqMzOIE3bSqB7h6RvMoiBEZb
jm9TXIcRBjBoETgHUMa70OdwDOU66EKOV7O2LDJPBVug/YcHdz6r/CbGAYiYaplRBkLHV1pMmlGd
UkKnY6YWyR6h3EQJdZxTifE9VG0AtLR1GQuiiphwmzDg76UEKitF+MEeoLvzo/faBpD5oo/ou2GF
8x75baFkAkqn7/Qc5VEfPmlBLFPRPbB7HuDrQP84MsJk+IkJaMZH2rHe+Ohg3Zy6jl9izmDZlSda
pT3bVIPqiahcCP+JpegUwXoh4MFw6217t1sy4DXUF07AYv8ZtFX6TuBT4zTeX5mSV8jiFW0Zo+LE
i5SOyxCme9qN/nk2gMGB9HwrajkiAo21+8jIYTQMduAEbdYwPvim0KRgG5XSEdgLO3mNCHKykSFo
lsPwB8puzZAGIoEWKtwX0Vddub9iq0KCz/1OKhnOSxMwyMmHvIFrICFmY3QuOwVuXV0G/gQ2FSV2
6OtV5YvDf5xAAVvMsTJcbSoj/3YNK4KcM4FWE1SlUyfC4vzLfBhVczJaT4XIB3GN/QXyZPFW/mFI
PPb8aijRSMZ1aGpdvYGBaWgWKjrwxZtzdPxKbszMKsNbZZqpQ75uBC3ntsSIO1lEsOT8u9satXMf
8dO3yx+3x/t6TQY7FhYI7MVXdivbPKz9HXGpdD4Qq/m9ynBX41vfxuMPpEo4cZTYKKZd0vGFotJd
eXPxRF4I0jpDm4vPTEooEoEKExT3npOtDJYrYPBo+5q/gMTxnrHUM8Yo1xrNzkUDTzxdV9eWiN8F
/QIXAmaoGUEMPxORn7Ah6nSyTiCCXbOftqjVxzJprG2XyZH5ZiP3s6HIAfsHzq74h8TRIJjtiIS0
LFgB1T/sq88CHcHg+q8OGXJMA0O7t+THPOWnh4qrjxfl9tMC1+VlUEsZqtqTN5/2cGPMRH0bN69Q
r04RQK2afvUN8RoQIPlEZKNtIGsoebipzBIf9jJjRw4slxa68tSqY9FpODP7Yazn/bk8Mol5Uxmm
tFH7rFQDkM2Bx41vO9FmirC3y7ot2PaNgcn8BvBdb1w2eRCFsvgFIRnMc23V/47rIB2Gs+o1bjpx
+DNqF4nCaZ0ddBOjbPB8LFtPcayQM4EUu7YwRudOa5nctH6zCdRao+xMzoRYoynbaUmG6uDkYCR7
0gTzenxXv/tgXYZ50faA7XWATmJgsy7BLSzuC9tziTV0lMYtw45m+H6ziwHIjwKpZG3yhX4Vn92r
QPSvdset/TZWE9/mzO4h+4VWYEyFrUqFhqtg5NOhuf3UZSv/Vshpru4WUx9cQg/9BkU9MO8q8WlB
YXhjW79FV8fAJM1YdD9NGtb7nEFZJJesgjlRQtuiZYAZj9gNHXnWjX5NMTsiKUgP9pLeQ+Kmi3Re
mN6WkHKjg5YaibAaJuKG2L1U25xJ4nYzUcZboXdSt73lL6R7h9rKtRfNe3QWmExJzJJi6OLhamo2
APW7LpIiLj03p2CBzfAqUIEPIf0eRzoi16X4k0e+6r/0mF+ShLy7VCTP9wV0BdVHDcxgn4n4rbu4
+lqPZ5J7rUFGNxC251qWrLjz10HsWCWeX1lcNlV4HZOeU3k0Po9T4fmeR5OaUbqzkeN/rs0f1JRx
n7o4b0AfJZewpQXPjrJatjwehpIhi5jFgGhDhAS97xzSd8IBHDYRyB4MG9O0+EJsxXKDS9IKUwgp
fvM3dnELTjZeZ3tB95uRJu/NSoYyfXBjUjN1oJ3jARSjQ2nAaV5kLmgnzEW6jFocQZupa26+fZhs
1WS6kKrRikRy0bqzy6IP1Jsg9EQcIeCtcJzVcVb/p1FAsgAHtiEqs1xtM9drnA2lDbws2vtdUTcF
5AQVpVgYTdP+TqmHRZqx8Q9nCfJqhB97oj33Cn4xFABi4enjjI/l8kZ9VhoJDNwbXaxBPcekC0zV
pyf0QC6ndOs6tO7gpWQVRtEUTiWguGxlBe1v+i1rx7hN4ROkfJDNwK0QcRVmjnd3cSfTZs4sMBnt
QY6hoJK3sq0639fGviCYsmXQZaH3GrMWIcQHBnRe5L0tkpAGvOHeQ2zseFobmvweiFPGWZ5D8IjU
dYV8EJkToGmS2D93cxqi1WdmFG3RUkGhJ8PF/UvvGG5fIqoJRuBPMJkWTfIPxlUsifPst8Kzi4Nm
DjLnPqn9H01BZxaGD4Z9BjzPe+ci43iZggaB89Bj2UWh/19QVfaM1sIfpfZ+Jf6d97TwvVsCl4WI
XT+yuz7FHzSneagyz3qrd0xjCJqRlTtx35SDvrIdnpebJoLP4nD4bK0/E5aPMtzxY87gS1YhvvHY
+YNbA9CFGhCq337Dq95dzwADYOivzJeSGePUNkasaxkNpMdA1JFaG9yDkKdvOi0XVz2x5sQTXRhO
hSHyzXz6eyynz8UsGhH/Fix4Ve4mMaNJg8nHEaMQJUCrVfYjc+qMt+yk/an/nsorYHj5VTVfIrSN
H1Q6cq9AiKxi5c6KwWiDtNLBzY2FXECEgU4LAKTQuSvfPeeFY/LYSejXXTUJ1KQBGTxgg+5QngMR
GCoCuitAD9uXsS1vs8oMHfufkJ1jA9z3unbvYbf9uawpX9B+EtaCO1Pzf6M6rFqZgusMIEIXLWdw
okvKB0ikZtrKjBxD354VjIeN1e6hUyBLaS2a3YG4kgGrmkzDZWVN+APJBoTjXwyxoTXy4hlZ0ctC
n2bLQKAam+ItxsAcZMsLJc5VIjpDVcbjAlEK4NUUSSPbZqwhLWHozACqXjJqktiefHHCH9O1Bv7V
dUB8w0T/b0QXq/vuwhVs2CH0uwxOvCPlgVptDyqns5wvNZpPkAZBTSsvKlJ0yt0k22asedrz7aEt
v1hrXTiicAWCoCqcic1L5tZk1ltjyqChcEju4k2QTDUl65v79xopgoIwu0ee3iDltHqn3CPzvs3l
UcC39O3uEMmkTpberwf8kWOBoYKKcnGpndRcvchc1ofG8gHPMVA8HC18hCN4Qq35j4quLOptul+R
GVTPpgrJPrrQnTq7hKwtuCSNEpF6WXtYDuMGKbNpMeVDqr1xUx9n7FahvQit5cCeVxCeBa+joCoS
MiVX6TAK87Av3udBSuwP2gLoGRKsYPCg3eATu1hlTHPYAaIC3iN50a0a2+L+q4Cdl64Hyysx0SX7
3Skn9x5/26Bwc9M7d8AZ+5yIAqEKGP+3tfFURiGWq4iE+YYWlcNM3d7IWiGcFA15YrGRYfO7UsFs
XS6b6b8Af1OzadllEMjB80BWTt0MGxR1VjOhiBfa8oxMRvUz+d4IdlLRjXAIJckZZ3DiFT+4Eswx
shHzMrATjFBpg5VZoqehG4kUskoyobgVMt9ns5ztOuDnM00510C8mMmVb28Icq0lB+UbUbWIw3aj
PUlNARoLZ9DydDqT36xRf76ZD1f1VOEx2NiubI6+ePfd93Xcoz+W8xTQg3ccvwbZXnZS6vZLdXQC
x1k5dM37w8ZWtYsfVmVovzhKgXNxYp6K4ivprTUumrjBays8Tf3R/Dd3fnTv9IkSuTqwupME/9R4
hGRuJZFBXHVnpGa0nW+a9lCAwiqbQf6msS0fAmJv0FBZ2zLjeliASudUys+WCdsaA2/3tcVP7gpx
Dj6LIEZcloFqvIdkw6q1StVPCRz8F3LBQTtMtCZPlksuaaomr5SWYZIHRRCLKZk+Mm9Wr3I//JWS
if+iK3If08OyKZmna/s4rQANGbrCZ93X0vlm+F3Z9ERogwJn8tDsNWgTLRY6kwLoG919iDfS/tWT
q9qJYWPToZxFE7kZqGXcwOI8WAL1bhroJ5fiiNVoefnKrM2pQ0rDmM4vXiQIr7QlQes0BQAvnSYw
QWxAtHpD3fATyrwQP7pZ6IforP15AZMajcME1Fw/FdWyeCdYQ3K3Rfwa5IxDK7ksdhIyec8lupfq
IIhF8OufE+ij6zQjY8pZS1Lb2RsCJu8Za3Qfk9w3Lvlb/ShrjW8sviJmvEvtHPdMWB+o9P31urgL
GCogDAS5Q+5eNF4XH7cfd/VmWQ1FY5kN4IDtXFHWUdcay3/76h/44aQbFQx1V4EtCuHW7WRoXkPO
EaJPIRm5soUsLcQFejnoSLJf1yVWazaShH52dKXFXVyq0Vj9uPmb1n8je1JLZQaKe9lIPfogZouN
FzoJ9TY2fpQOsUKCHewPHEIEUd3nBcwhVjtLgxKARFAoeKL0OMtzInC+EBu0eBAbnoG9FyUupL5p
vpOG8RTZWvWjvELuRNd+yfhtGiuqaOt/5RHaYV66O8H+MfH7VDuXC4KIYfbycrAhI7sN74Ofqcf0
lCGgv45MQZjgEiMi0+/jKKtf/WPibA1VE4sDvT7Tg5D6/lGC2xCWDLcQYMk06MPFucx/k6ANb0AO
eHIn4ffKer5AY6e5fek+RjJySB7dyU4/ZmQGlv7FsgapuecypDrPCMOMrivlOsY9H0Lu2EiiTpC1
kFoqugpLFRkb8FAV9ixaNhOSvvvOMzJTKx/yMZwOl+OlB2+xVH2Q/n2TmIHl3Z2YZowW7CqOOqap
A3D0IahtDkrhTHR1HsWQVFJmDCvgF3mFRjZPA0NWc2VoRm9lTWjQIsG2Bq/xanjLfshLoXNNp6c0
m4MQoZcofYokI3AbeFFnXLzVx+J6DNK+kxxb1nPp+xyjXkjjkvtI4xmd3ZtOIZbHHPfxyvMgbeV0
JoMXSAOSvKNhghBxy8zGgL978Oe0H/51REtieFfbn+ZvrqNk3hOsZBt1Mvh2tOgiGOPC4ENQ7o8I
PZdZpUQLmCh1Ghjt6QgDa2az2vTTWOw+874gGxuSLiH1H6QMu43HmBaikFsEmAZCqqOxW6wAW6cS
WkrXLly/8fShEz1zlQaTjqaWEtl/7lB3dZfscgomIiMxW/V2Ry41K4qTihr1Glfi1S5jB2J4/cen
NKRQ3Q8TLhH1g/67X4XZGVgPzXA/i7Syhg5chvFVC/8tjriR7UFhWHWFEPUVngLQLikE2DGB09Xh
qtFCw7ezDpUDtcC08I5kO0SSBjN8SXikI4RW+FQWsu5q4Ol9UG59MttKRqlOYG7ud15KItDMnFAy
JXCSbo+R+liLNtsvZ6Jw3a4IFa3bEXQqXCT7CguDlNrAeS/XSZhqqyoDckOzWldFVMTfu/gn+RQm
len4zrRkiEEscJXPIEQRKyS2KMvrhYQYeoKmS5vpEdZ9+0/0DGRAbRTBMT9La4t9kyhSicIGHPV8
zYshylHqKr0q5sU/WWiLHjCRd+5HN2wd9DfRYY7dAt3ZqtgMnNlkYHr/dfbu36U+dY6/gNGWZ9vP
If41hmljzu+sQHP/MQY0WWRIP7u3flzypQUz7w7+DjAi70a3FFOCIcImHCas/YvMgByd4zmlgwe2
LCtSdhl0Tg5po9qZBNcxU7AC8f1gxaVccSskCHygFQSz4Uf3VBBqilTpItPVz3n2d9eYYFXU4sDC
Thsnvfk41sE3WIThYebjaDOOApoKVBpRC3bgcUuhWLPPm8M6xybMl4oPOs6qH5FlLK6xw4rYa5WQ
wJO0aWOFaKT44oMXRjR9TpcQiR+9AcEIZyTmuv11hTGGTnNvQbh2/w40pBzHHkhUTQXlGxMhtmax
CZ/8C9ZmwhoLJl5la2aUnX+2raW/dpAXYM7qmvC+pZ0U2+c7TdlEQDZuy3JyuIRJNj2+J/d8lyHJ
0J9Rls6F/SIyhPObvhnKYewRMBG5pTPlyDZ402BZJ43UzV1I5s707AnI30lFEv1sdMX5CJuJHFcg
+SFrlXDP/SezkTdw5CIWdDt5pub3/m+ciH6bNnnL9c8Ubxh14EKWcmJPYBnSfrj1TcyqXqQSqJC6
gKD/wqDEqs+PupymIoRX2R8WMrVEEwLU9VDOPjo4pwDU7phMN2y4dYnh0+fc8KCEwzzlqTt+5cze
olV4HDTn/DW2zmaDYw8TCEIDDiWC/jFKExGlj378L2berhhiz1g2GmsFDn5+1TzvAuTBT99IEwn6
obzeDPtHKpjyxlsh2sl2m6UZun0AqFl9JnqHnAWwZlFwGHPw9ucL4EGAEPNLys4vUheRPAWiQQoC
GbbFxoURe+gafJqpptnbu1xdbs116a4k3LS5v+e3z/zG2cp5Qh2InC0TrlCZkjQaYTM+K/xFAmlX
2pENLSaX5vvP15c+TuwL9nQ6DAwhp9DnnRCBy8iEmiGd1cFJC9pVH+J3P/PMEBsyULpcgc3IODRi
jQn2hZSurkhoq89ozMcVUcaz5R92MBZGOC9XIxQfvZKC9EklLsagdjC3Ks5XDPBwapfMbjpYmdmW
M5WUR3doKnl0rr6GDLkZUF2b4N41XWsMhaQ2/w3g4nbKcPBSDDPBJCFa9jkR1MgrlgCZ08H41rpk
xsFBNXdHMoDWPIYqJmBskjk/PEGSobdpGm6rSKTYWNkZLPOnIjaNYuyJeBaI6pMdRLymbLu9ISwX
J5aDZ1VpwJE3+GIaHJW9++xiEUjIpFvqioVw66t+Yg7Soj3dLThBxgBSRHlBL+646G59kToshnAx
d1QhXy9bSGeTl28cqVByxrT6ziTtMBQZI/62oW9EVbnXubcmPckDtIHm/d3WJz/fNHN9XtitYAcs
Sol448RvXFO2TvVvq+Vm6Vp9S/T6dT5SLob0rYMiWPBrZ2/ZiHhsRCV9Es4puRhW64pqnVdcGTyA
Zl/Ly5dB9wLAczY2VOyP5JONGrrWkEt4sIt8H6D79SkQK/kkMLnRfXC57OjTRLVveRJzRJ57cLa6
MJECVidrA2XLSNJdIaH7EqQTBfrUe4aPbRgmeA7Q99buaAigEjG7RHyrewQ/+5rC7lc8gQK5F7aK
98AkNyK6+TXerehuyaByWnLu85LQuAIXWnAd0kMKvPU+KmN8oTSJU2h6dTnwEhpjS8aFKGTydDXr
XFD8wbu+/kztEtP4xkHhDeGSZ2GSLQKleJV8qDf98T4EXrJJNVXKeU8a/SiSDxVXk/pINioZ8O2K
JEepthkTUo2nx3dtqb92bEgcxsIoFUh/5O2lHVm6FW6IkT3i6D30EyHRKRcpUv2WSMl7HQL4LY4I
geo47iEeVYc8BSQc54tFEF1l0E5TWScHXHQFFrkCyFjQOKz8VptSTW5BLaliD/M0DjL1cMF37cN9
FcPZl0XESqD+OiO+r1riJrJDLgakrrmrAocPwg/brVrs8myvlohKmplC4ISSW47CGW+OTByFqoKR
Xv8iVac6ACDcqbHnDcgsJ/r2JQwadKT1MaeALtjDSzN42lrA/SEtUgOtTRsPehowsAgVL9coxEkb
Kv9SVHXJ3IMWVe81KqULr+U0aNqR1am8aL8ttZOsR3ebMZSem9CEWKmzowESjDsJ9pnLWIQxISb+
O2tdQRgiHDrwe1OA87yUZJbEzAYhJMM1ndhxjdfexvfxjS3fuz3kXWtpFiggrLXuit3IaVAsJ0Co
93T4cWNvzk7kxQnkI7zNLYrAScIXBqYGEQ3j2InRbfJllnpgMGCMgwLPBU/1dweBit6TC4v8lSNW
JKuVjaNrLtcn5tUycxIx6b8rKyE4Kzd4qhkDMkcT0QW8bxxWbUF1Nh5L/l1NcAB728TZGawxUkDN
MMQcukJqKKVusQAi7JaBmA0oCqrEFqUNGu/6TaovI+Am4aa3cKbK+8J4uMFl2pUxNpJMcgmsVaIg
NKH99yL4UfD1fiVJGuC5Z899LazZDgciWKau83mqBVFkIxv+NcBsNqfMiAZ5f1W+eD0Gk+SUzMDV
dE4aLFphmR3GgKSJPpzU6HAtZiKR6KBrlMYAbOt8JYbFnxDESVByzQjdY51WiZKQfcM2F92uTO6t
rH1EZZKwPjW9L1wfb3fxaw35HDTNYPCkJIJQgnagReJltPRSFT8Nbt6F5lS8yyvbTUuSZQs8C7b1
IoTYQ6Xqj4YCNvPDjHelJn1Qygk42kmm9waZRTyNTZekM82LMoGSR6MOtLnc8N1UN8WD9XfBc749
B1cYLlwgQDnTvjXltc+Mqh0om3L/QZKmwojGjFBvdbhUt4ovikYObXSRasUI8TJpMz9IlgFtIiTn
aZuh/nHCsT1PJQmHfecHOZO3zEs8ZIeYTJHEPKv/7URllu07vLjW/8mKHkL9MsDLjh4AXx3T2R6b
ZRj5ppcHSBPz7OioVWHA94mASlndLqoQiGgSeRQVqs1v1f4E3eCa71tKCrDoLS5RbBoiyQs2/5Ta
dJ6yLWtup2i6J0FU6Ct4rgchfsvcuIMb/z9v4x7m54JfkEgIMK85r11gPAMaRmM+LdWV5ZDvzIlF
eZmSEHoL/ho3PgB4jlB5ijX+YA9mAxcVBhL3dfKQchPvFildDY9Y2pww/VLZBnEoEaVAImrkUm6u
KmcFhvaMQPhlHDOEZGIEllqbxyXmn3opjrfyKcIRr3CoSxCbdqSaaic0ZFd55YZfvzZWkgaHy6KP
wPs3b/dYdMD7KgOWjutMbUESrUmwMtijPf4JGIyzACKQB0+dH75l07HmKOijjWDAorxIc3ts5RVv
QcM/YdSEjBuWtr4XNFuxwF+6w7wW7xSjdBwgbmd91HCR1TEE6HvqvpQuIDyLon7+Tf4xb/Ld0SBz
5QN3/F4RQRlm3BXrx+4KAjLApTHW2TI2+QbWke8jkB2W9Jb1nOgPmdu51ntvQLwtgD4YN057lRcy
ZQN/jtYPdJ6gMUbZvyBATq6OKWeGiMkeopKujh0X/F37UzVe2bErpOXN1GdfYxk5IQaNACxx6Roa
dSzC+/wzO14uBxfiR5SnypxCdIJOVFH1qnvONVP0fGQo8/VMT3wwSqX2PEZAT20nQjnHEUNSxCH/
a99XYagG7ZoPBFzZ1ARpw4dv7Mh1E/TGZKVLOoCGgsVZ7nH4Fp3nL6v4M80RgOvqk/SByuDsKB5p
ShyqMs5+SkXQRP3YI3p+4ceo0VXfAkR5kVsbt5I2MM/UJ83rASGiAT30RQCshbG9OHkOFUPaDMWl
hrq9RmYdjXmw2GEqbPE8Y7sEMaVmqKtTlUlO9+SLgUpldamZqoJt+IsjCZfxkdSbG7JxrcTk3vXd
kYgDzqEQs25OgICHvRIC90cG6ETle9F5/x2QvGD2Yegos9NWLKzVVtpQ7Vtg6DEKwcxJKbMJ7JSg
8gfWSCUX8no38VekYaIiXMYQQ/JyUxcRgR2dZFX8zIYMEAlRaPikMN9ESHe2XOFgj2F+B+wKtB1H
9nTOl217Rorl43AIrcaultF5vQ/dOhaOAMcEOsKUcyOxCDkMsu+hOAqmERnSGmeaEJ/4hfnr6osG
5z+ZuS2RcEsripnmIp6rFENHE5lCx5D3zAteWT3ajsAqFm2nkEDhhtsSngkafxm+VeFqQhn2RrCY
A+UM3l4/zL3/RC9xvqS/lnWDeq6A0NbqSzCoR6LrMhQf6QUIEw3doXcJ3FBChbvOJyADbjrtmBT+
+wCZn3FA7uTdfz8PnSeL15l5BL04Z2dyPAoQVLlNGlUZujFQml4KL7M/FTmuuPnkPCMYvM+b4nwq
xvXDeAgjSg5ON8qP4tnqKd5aRnMR59WorbeUFgo8Bi7tdA/TR82ixrBoaYnTRQH9qrYaPrVLB2Ly
sIyNGcPMZNsYMwh0LL9RQCyV8oe7sJMIFUkYycjmYzY3Tm+EZ1EC+vrEmQbbbaWDZE3u3hNLlk72
YJVAVWDpRp6fARLbkcmP0iOSRuEw6oK8TJ47BxJO/I3WpecgQy03NnXhmIa9D7xI8QQEdplYPgoK
oVWoPWuoJAGDl093d+OObmP6oHNjsUKXcenovFJs+3c0+41qMsQV0uuQ8Ag3bKTnaiQogMe+Z79+
gxTP75RA37+U4U/ZNP+VtMg2C6gwxcgtqYZG4pluSorHkKGVxgRF4y+zf05UH/ApwGpgGM5vtrnk
L7P7KDnAHxB73c3SUFU/0C5McBsGa930zjuOrLL3dpEtu9VX3t0xXknsIjegYv1/fmUumXQwbnMq
iwk864VdICGfntZVVuGraJikL4hpAwkoU1b3k21Yx4ZvHfL4a/Mi3oGs7sJwrfcCgFAemsVM25rt
MyMft0xBIlBs0iE0CWXtsX+XoMR5p3YU1zt7o4SgwxJwrB1mOfmcl5mLsM2YZ+pcwaBJm7F/KZyF
EOXo1ZsDpA7/1vKZgQyjOMcYmDlKy4nBBjKRFv9mAun1MKW/WKsbx4+5Rz54TMq1qLCYqpvhqMFq
YbhECiDaG8PuUoIfKXmr9vGD53wIPhIAUuVXdO8sjP6QNOz6vYR6yr/ER6vCJCOUSNPxcZt/U6NQ
uLIJ/G/EjhnVu1y3DzSp9YIlcEmDoSD11+3plqccaWh7CR39I9rcJAQxzMm10Te4yYX/SGtDts4C
eVPHZtBn3cZrvLtEOKDBF5ZBB4Y/CgLGX1gNM5IpZWQvdbsfTp9OTs03nMz4khPMrO1ynAwMn24M
drq5OP0QjmZfduY6WifqxVznfLGeYnefz7ySpCB4zWpWVEtdlkXATEmnmjPgwdLoD4bF7zBzzu9R
yxSGZUGPloAFjSdSOQ8kxXGh2VF7K6Gtx3SgRIJ7Z2ipCGBDSaiRbIG5RbMivBWeG6aqiMK3y5MP
TlImUmRihk/oeHdIsZkEJ3hpT1YibZcCCeYRyskZM6ZVE8rw86v5JfJcuptfYgysNGYfi1aMA6Xi
03x1YdfByXy62NtFXD4fAYPfYUioylYv4bHSvi0kFxvGGJi/FyHtH7zhyMULpeLqbpLgRFDok0s4
zXA12AO+tthS899lkUd1LgtFm/+ShhRJ7np9BPVQlNmgSw1ciVCq4l6DhYQJ8LAh9rTqXiKP3ptp
qijlYM5zFlPd1DqiGXdxt4vVzkn7k49AOnHVF4bGF5p7YLuWImiAUPcBm2HjilbFSb96GVzvdcFa
kJ2GlHNW430HiRv3E3pUF4kkYmbRY/hjGUika4I2TfCk0l09rw6mJ0vO0CpWQPfQOEkcMyEGGeoZ
OiBOGsF8eWslxOaxrbtNkoFyQW7J4H8IToRylOPY4Gq58WN2qIu68xCQkLm/Xmr9M2BSRdw3Mc8Q
4Yey2qsnCgOUgF5W6xeYHCdGX5J/Wz+jT4zgpH1GLRPKiGpPbJPRmMtH0O+dxTorDeBPK8sIm0Hq
D00hFGdGS66gWoV3vRH4KfrGl09H4u0e4Rudk1hQ2GFeabZ5DkD1kK1kdxexnGoChJhjsIMKV5nB
GWHeIz7I5uAWCeMgv5QsaeCcGYGJSqsJo3Lw/6ntgMOmLClPAEijOnvMsqBR3ZrVvRVPY+m2XlwE
8i9inopOqsVOOYZiwuPc+VULAfRZpdcXncSD60K9iLVaGcvdwPJos5V3M0GfKu0PLE9b5pVLnlgg
dC89Mhuarr/DHuD+banFFa9e9Vndj2Pr1a7si3nw4GPeQTg2vKRpgKY84u2AaND+Yb3t04J6m25X
QZf2Txn/V3QolNx4c7z05QkOX3/MwtcJcReUGP8qBKygwsb9Q0YcHHH2maEaoxIeukDuX5f1JoUQ
7dHpMmM0Ae977YAMsHOZm2CPWpL1oSmOcXnBGT/sktPcrOsDPHf3pZ5pyOz2IfIXrM2vFaX68MO6
LV+AsbClU7PdqnnPWTU4L9hrxMHsnwCf0oPBkrXOFVSbYqxbQ+KfC6/XXQoIr085D9bDrfiqYK/1
zkJFwAXObWr1jWBkn0sn3OacJLy3JuTgKq0amiRR5uJm3LAuVZ5fieStn6AEMjH0Yw8hXAVCrcP7
ikibUk3W9LTdxr73Usv6yybwPJsYpFGSZlLl/qblVZyScd+Gj7kvDZutXE+/GHCCKU1ZgJ9LMGyE
A05SViXOau4adbftTOUNK6jMY56Fy15LsS7vFxNxfDLg40U74nY3uEYPWTZn34bbjXQiBaUattVy
EG3UVYZ2wwAHnFejqcs87u5XktSXZBzp1pnfeVYKZdrY8WQjamwwDFqMH+PeftTpOyW8240WSCFR
7j0ESZnw9zBD/dIyZ7oaQcKNxAVVhpcw8UFTgbvwgpDyZUGp1Bf6wyXCtwkAXzDuByf1S+rGH5gk
Zvzwgmc3VyYMTo/BJyezhAL02ViyNWGArTl+myO9k8EKrTUUv1qR46EX2je7mxjB5Bdx1GuFeY/O
dG7vHhqISEphXj7b4NJ1JbarWP1scCx2umLYljM+GbdtYwRZnsRmtsJgeOzcSah84psbTBVEjQyT
z+3QOoeQe6fH0Vu6I8Js8LxYZAJUrfBcS3cBydJMKtCJSuEBko9XGLQkeAXePxaa39ND4gjtCGZi
nGCv2Hs7JitpjxtDZfH1bM65//NR/JM8mfY/frzt4ZC6mqbR+QZXS42JyV7/qCqp56/XoS/SIX05
OVB72Jg11ogJJQZUBZUthld16rUcLW2m1wVpuikRuWW526AMv7P65MiubUsiq+fEH3U+4sv5RUNw
SSKzltWnnE/N7gTVy6MvIOpugoneNTvuLCM03U0jYQxXxTHis79QgRWBknc5ycl/x7Qtnulzm39z
xgO73YS6uDLgn8n8IjLXxrpE8nd6GPB/rLKzBxKavoDz9VWaRmt7LcNgACZHDFrU5RbJffiKo+AR
jK3poNRnLgy4drqLA6hOkEHlRN9tav64aND2iUyiXfGbUc3WiyYiPn6q6plaFAOZZWAM8R3oTLmI
Wf23whzu/xfIb4e9Hv2LG179kfCRJne4I7MtyA8eCjbyS1YS4wTTZjAPHRp8X1xiCe9yHszTq04l
tCKwa8mnWnkB8Mb4pEQLyaMcXfB+0qkly9ps1cKGv+1N32OqlVRoHQ6wN8BfO0qrZjIzFdmnb/X1
Spo0tQ7SZyw/BRAz7IMrFh0U/xuVBoP9A+N9jicIvbaA9EeoLXogeK8YLvkxrCze4zvr8lWw8dYo
hqmoIxrwMHnoVGhy7VPQ4S3EMEFHyjb1v5nmjUDtjMypXjtFm9pRgTPtnp07GrZqPWwVxBePR+Mb
Tn8OnSugWzv0bbulmQLJEVzdNbcr/tNWjpMTINSL49qmkMWxa+67n6D0nXUAS44Ey/91iLl6dDIR
zYsXEJkTDr/wBlWD1ImOn39vhj10BDk1ixrgKRQAKxieWzU1/4emK5HNZvT7apTGkDYyjj8jZ04V
vOEoB12TUQD/iWo0qe/Gsz5zQDDR2JVHr/o40LxEyEc9HqlKH1pJM3Xd4u2w8pr6w/gbMheFx4OZ
rcbWUk2+ZzevgcOQuAnSw8+Qcsm9PxW3XwNGnmipbwY1roO+0GYNWyyWgwbDI56wHUlFUqlqqQrB
l3zrnuIHiNsahEEfkgecJnJY6urhqt4+A6fAVX+n0VVE4IAOEoDVl/TiE/mrvz6uCb0rdX+URxer
XFXIY3VWXRrU+QOJcSrKxjPwmWum+faKlIXHA1Kbcgrkj/9T4CEBKszaUS+pdGJOoBi2PXwMc/fD
TGG2VNpLbu/WveyrPb0PbhaD4/XVCnMdbH5cj/YIsKe/fp65HXZz2H4c9XVqQOes1gLLpsUi59fj
ikPUYn6Mfkz9PaG4Csi9H5Gutffod3GF/BYFQsYCRY/XvFvYoDsjoJZTwteUhP2GSlwMF4uarSiQ
qab35BbfcFfCynsPIMceONQW3nsBfIiPt0NyUgVJY0hP4Yre/mYbl6QUgSQZujvf5l3mkI35omor
1G3XZT9EVEMO2wJI+yRcA5LG+F1l+e+lW2khnx9gOCdLE2cm/yVw3rWMAY7zIAg9xVs6bMoXTY1h
2EHblt2juC/Cwuhhf+VsfyE9kaUsKGntWKGKhY0LMf8UgDwhOxtyQM62xTBok8gRD8rEF0YOvaOt
43fjhDRqVy0qD7GplvwC1RxZTKAGctAePjmtp71Rm83iTwvtEgGO5pebNqFEOZVd1Y55xNzoQk46
6ktdNZKJFNOY3rPmkdLAwXpYLLUpgVPQIGEprW2Gmz04f+vAoGZAxtpRyxiCNfNXAAW5lklXeKjD
eQJO3+0Fb3OdSPZdsu7U8Fe9WxNrDv2/hB8hdGBZjYez3AHemyHrlZ011JPxoGQCn9k3MZ/X4JJe
2IsEThA8fhfx0uJI9yYXVbRhmc9I5XsCqwX8Bwm+GVshGh/QF6Qf1gOeWLs6esRlyzFag0I0tENE
lGJllGCjAjC2sHpx7H76673VSiDb/v/AddTSVss1cPcvFcrluFJMVc65kQlKY/XT49xYZ0vHU+Q4
vEfB7kQJh5ZBGqFBZ8Hd+Uni9zDPyuevvI82KLtVSodXrhJ2QWU8+Q4ewT75ZkYbx7ZaJBUoT0xy
6T/yd0qG58gbtonNHMQ5FjPE2FIF61QLU99JLhTNeiwOMV6oGLgznxFlOCnioNX3npoRCd8ewYtd
GV6ktFNddCaa40fQjA0M6wZOP4wo5u7oYfpFmUvr+1wRKATk0GSSy+qN/+XIMmbrD5zuLVa5cc/C
QzvSnb9CfsHCLZOb36B4SqCMARB9v2GL/X1wqN+ayHNG2jdxsiC/b7NSBKzTaOJ3Ah/e5vFW09/V
8XF9sO2ez5yIcKs6g3ADTsbAnqIgyjswyn7Ccf/PSSoAy5MV71BtSXBrMy0OAr1d5oKF3sXSNu1n
nqiy5AUpO3yI177bMgxfbNG4WGV+MzeZMGPn/HXfHyFW/3JyTlh6zY4tom8tBITqmmJputze0JU+
zmtWS2qWC40SN6jByswX+4cCAnHCxgbqogd23x6l3rtQR3cZeGZV6JJrCb5M4ZsruusESUcdlrZ7
Ku9QLEQzp0Kn/vn07yiW5J2UArEKxWP07Z9DmixjhLwo6G8NJaZlCNfZaXpTypJP0lqgW7HDvRAK
PtUb/U17djmkTwDPYjIVYT447QiWjYYxQq8VxrLWahdR2dIphMIVP8e6ojXT7YT4kpLn0njp9bnt
Ez/c3RsBdl+Rl/OqaE3ZUdV0jQancnDMWJKmotOFVG1u2fF8JCCLJpCiB/FIqDpPF6EgUyBdXIxT
RId968dzIJdr+UYEc/c86rG2F0XKAiCabaZW6xWj2GvlN2i1DrK6JQf8gSVIUWjkyorjaaMiX219
pNjobbNLRThMMSmhtBXDyjeVP/34InOyxt2fAtoU4Z3fUUOeCQ+QVznXHQbtnmU8BG/wpnzFTaGX
1wfhQ0OxHXQVBLoGAPYQwkGpUJd89UnrdmJLUAXx0ufPKQOziliSF92mFJIl0sE5nZ3BI+sVy7i5
zyPzch5bzYm0SVWHZvigWp5XtwUXrN0MO/1A85YN4ctb4WShQXiowUR3IxOKQ+/tvY2Rde7BS01e
au9Hlvl3abAk2861ZyaMHyYfAcfabSx1uKwDyxoS7UXQttvjhVMe8GoFzIFhzsQM0B3Rp/eVXGgO
iyT/iuqI2Igb/YR4ZLnEFIbBwMVhfYtRiQL2GZOL8GcJ2xWcV64uQkl5p24Fh4IZvYS0lxzy5Zet
Rgjmovw1/cPNWBBv1widmBaZRXorimK8oEjG1sdIQjwwSW6m/S7mEi9hH09W/ydb9G8lYOPZbYdx
8LBkIuFkmCo+odiWor+a/qWgIHFkGaGl3uGdXQ5uE5CuCIz92x7TgRrmYSPqRccd/1+6Gw00WcZh
2dj3jwmaRdBQITMn6/7JiZrmgwd4FwbAi41NFh2Ah+kA4yKFeSvPCha4j9BO6jyAK5bbvKWz9WFY
6lk0SYgb0PMRF26RLffhlgC6BDbkUYmtKgVveU2hP5Z477nINyOXk7ERFme16qN0OnB69E5QGJHG
D31U8pdt5Pif8tlK1NJcTLCJBIoQLeUeVy/Y+3mUYyaRU4/VfcWUOQIer+/V45F5Ye4iw31ZIy+C
2zczqqF6PzRtjWHvB+00+ViN3b75of2J2UYS3oOzjlryROVUpdKYRZLIhzJc8JT3WD8d/PjY7vkx
wFXONS70Y/SPNsXyJGi7kTP2aYn71GsS2KmIzGkRzvjdAiD+4JA138RXauZXiqfHhSW4eUelFWtF
2vTM3sfxWfpAdfhXS/iOwbUFjHjkix29tfHHYd9IY6aFbqiM+v0OTzTSTDnn5lrexyl/BC9/A4p5
efcjhfoMyfJuqAyuF6Sc488n8jg/YV0dndf2XLqkwuxEB1wNcqTiDh0WEIVQHSiZxNPRLL3rLQsa
VweQuDfCFlVs6wAagKvaobYkjO6JPXC/ADuKVyBVkt/bL43Vjpficq4yEJPX91xtPmg5rnLGGlq1
BU9WhWzpfTov3vx5ytJDMOnMtEHGiGfXFs3iuvpwPbjo44y8m19LTyu78r0rYKxNINms04XoeUpA
wCeDAR/uDUWgRTYNA0LJkNrfjyyGrXqSkZAyGGTuSmSuFrCU5493aXUG+YpwgK4T62URN55aOESv
mUl3VN3oCCqSDHTcLGywFsJtf5/32I5Cz65AgeqNX7+Q/a1V+cldN6wDAxhEJzUe8ff6aee7ME1F
4K5mABAThRwj/iFhW9umiSrdoUCIfHwvtQ9II3h82SRBv9mAcgLrE6UryBy9o1i/pJ44pGmZgY51
Phvm2/mSTV/rxs0f1V2uoYtlEdN17LbMuAIKbnBkja7YO5ywobI+rRKU+vmMrrL4dLVN/K9KsEos
ID5aDGdkN9A5WCnvx3HfEO6gplWc6+98qkmlsvgk9PP+bSWUXBLkShKlIcBM6XzMplkgeYiXE26+
/LZnkMWcJ82Ub0NGxjvPr5I9uBrLezyr7d9dF+is34bVMOo7aZcSsoKFoEUHpYyaBBl6HgZ/h3jm
OlnyE/KoYclaIPN8NHNUwEvZeQ+1NTdoLjZiMIc2b1st2/sk0Q3irwUXLo35YBzaZyvJa66bYijJ
5KevjVXmh1RXxcftQVb+EAh4wtALzQrLWkTR3tD6syaNvrV2N7QoC4zhZKL3JVps6Z0jzfQyONvI
r+Lks38Hb0414K+9pWed6vGoWFkaxyP58g2FecUbnUU0JDRRFJ+MXYo9xd86DtWGajQv0V3EREA4
qtOZXDhPuxa92FWrcXafMBetnEvy33K40IbTfj2oOe2M+lt4AGkNh7eVufTesqBxLvATr4sPU0Kt
YxfTsO0k7ijUp3F3/JOOoNh/nwTCEUTHWgIQ8lBLQzpcCHLgtXTaapZLUdZ7c9YKI1BBQXP2OdgD
H5C0bM9NCNqEZv3PQDzbm2ADMgTMXMI2d4hpfyNRt83NI+23wJjbehg5Is6kpiJn56ZCgKYryW3E
ipfw3wzwXNdPni0VwuBXy51b8KBLkP1bOoWmctMXnryuSSuE4MT0Sr/StQIY9/eCcrpyjN1EKnnS
RJ3aKC9sTFPd3iCmNptbRCJfKsAMa4QYyoruIQlElMVDDOMYKXAvNxp2s7ye6kBr4sQAkw1NyZAO
rwcVWSLEObwGAX5msdLpeIFIic37e5Dr6TcMm+VoxL7/+K06CbmPBfXNjW1C5hHdvp7B+L7N8ksE
Aq018vwBO3ibPxJ73773aEEBszxcGnHYiJjFJcLnjWUCQEdjGeaB6HdBHItC71ZcAlCCvimZpSY+
Vsgi8VGO+j//DG0mB3ls2Mtrt1iD4x5X7AlrLRoDLw7d0jtnBWTj7VAIPfyXOuURuIuu3e8f0F28
mcfMQnpzG8gRcBqm79xEFHf0Mo9SOtWW/VuPxQy0w8N2LM1IHgwhMMMz8FyBfaGY0CFfQk+m4A3p
gtB1BZmbU845whnDys0DBX5/tHQM5WDuN1leTnmbb9d5vz6wvwrLfejfZaYU1Akw3OcC9+y87M5W
vfmzHhMHXSklsue/JG59TF8LEJpXlLCZ5so7zBKohGrrTpM5BuI2BZs9XTFSRAIbhGJJ9HCP+JwG
RwBppvg+dJRjaoY7KA579bCLS8DKGoFHjgqc/mSbJgwqVflWu5sY4k5wvnzh68OSbZISupUsNIGM
jdvlxviCF1TsN+gTmWHDHwFlYSrQnJRZTYBTCHs9Y2cTI6w3ap0nz5M8rqNgROXMMG4/bwoOEA4L
kSyla515T3CazpgYCMChxuPB2uvZVtP8L3AjbJEcHxeQi2jsMNXjQuDaXjvMrApxY9WprzQOK6s3
501eCqhHJGK4ZREiETrOqn2DxUp0S0Ikx4UhqPUq2hi+ElqRaauSn6MijDswM6fWCJKxWKqlxbKE
to16RKPDnKUXy5SEXP7O9tcumx0mz7QKteKe18WD0xwyCekgyYFt/da36u0LizwcTJz4IpctIuf2
V4VQksK6dJkp/EX+jVqsUnoSxfr3k8gwT0q1Kaz6PCStF2Nolc61LEN73HKe5s8Wcl/DcEsXMpQY
030EaWlD5d87GvHTOPaP55/LZdXT/mfhZJ+GnIc2YIg6Csg9hQBlewKhamyTI0dwgaoK8eCHWStl
wHBaU5tsGo7B1KVlTpHmgpvyEVeh0ZgtbFdiwFJhKuH6ghw2/T33rdOuOZHmqyrbqnqN3R1gWlfC
lNIz8eTw1EJEalRZulzdSIx0nzxMxIHQB1KItzdomIB5cv8bByYf6DXvEpObC3zNDQVHpFqtXhjN
Fi7qbKlUz8LOMGtgateFE2/OjWrAj7lh83EEZsxs91XgWy/63kBiyN4eEPJdoRsQIJrg4H5ODJxu
v6HY8kGTbqIscwBZoQz4xNeb3p0mR3LDFtyEObS6NssgnrxsBGXAd3hFGVnPXYRctm9dXYnTv+yG
Y5AC3FmYG3kyBmL41xUxbp0U62Jyd6dVcUvYp9QGrRbfOkhU+x1R1j5JgshD3w1w6VsJRsrpW+ln
PA0LtVUlFgLwnw1KhEPmjxivknYnaXG3KqmNzsJY8ry+tiPtDoZcoFrnSjKg7KB6NXiKELZbveJt
pE24pNTpMuOA70XB1/LmAjonIGZC5QlO/07WbOoJjoDMhOE1vqJ/VQOMzf3bZBh6LtDIbO2J5ebX
kx3FlPo6hJbLrQCpYNrUpayUxmnvW4s6DpaP9gPr/1j3aBE16YdgnxaJMM0jLkoqhApO2aFfLe3T
dZJjVGr2uvidtjdtJZlHqluuk5QXAoa8QJocIAZmNt8VHZbmEDpdvsby4f8hL2WRxj46sPtvEx+c
4Le4IYFFeWECSQwyHm15+ZrHP3PhN2A0gKMx4l66/IbR1eB4E3vCIa/037VkIsMZtkvN9i8oN6qu
5A6mr+ebISbVipQ04Uk4S9edIF7WI52gVkmBkaxeVEsk5pzLgnTc8rTyGxQkeefL1fzmjFLrqA4x
qFwyu7na3GXnum460DwCYilBpX/fIqvCFWTVrT9iDZ6SaUaWMHP6ySqYe5dI/4bZRo+LU2PJ4KYQ
aVhesdfkgrtVOjmlFIhEdKmMZOh7xI084GfJHzgwVAUGNq0ReOEB/G6EI0NfS4Ymq4JQxeGMxn7c
ORAjUvglEv3xId8Dfz/45mZApMtdoRpdkAr4i/HOC9xbeByRXAGddVBnqwTIUA11rUTbvkPPCUhv
wHoLY4cqdUMLG8VWH2FwFgQgVSrw1R3iKchnenZupKflE5Y/Icz6SpycKda8i2d4uSnIT6oKDQ4M
+7iaZYCTrGxjMUN2D9FsWFveYpsAlIlOAjNnOq0bEAO1WLKqUtEg2/kkGg4hvaYtDINJkmmLQGXg
BwN4bjU/JBWXO9t0ilsjeV/zA0ZMcmJXo5tfJQr+5KiWK2GFmLhZX0zM8G3SWx+VNddptd+qTq4k
NLYU9GI4F1S2H+vjNxxaPLVubr6+EmWThZa2cLgF/VexBbENyYJs8denopuWuImElXYHj/pbCvVk
z+waFrcQs1oTL5mEWXD/ak2DM8KHorn6HJvd2tSR75tq4YsnJjvPfKO6R1aGK/fh2glUTdWc2Nnm
yr2a1natts6JTpSCq7bdDsM9QB0H6nlOqA1Mh7XAjzLkKmaINBoMFgbnKQdFoowN8FIN8dU4wnZ+
LlIadZULp/u4EbjhkZf8CatMW3QYSYACukhU2T8XiZNk74Ohb7ulyq2mskYLBjlwR9zykmcfvYvt
VJBi9tzB7AFuEQbwvQ8QdExjjrqpfR6XGs1eY+saHUADdeHh4RjADuiu6LNCmST1XyitirtY2Y7t
Z3tphHN2PsgoHfRQei/zjw+bzTLRc+hLiFP+tfwvd0kTy9f/d5VoieD0PKzqbPjqxwqgLz7H5WSD
Kjb4P4f5Es3OFk1/+KDcamTeiOl2HCMi3n3AqYLKAOuPdupqFh+B+xkKqdUb8r1X5Zd7xAnGngKX
bqGdx8ZlYfMZWb3ev7++fKiDn+RvVYUa06OCm16XlFKQjTHLRdjl0Lsd8GANpOt2jYAtJj/O8eDK
6OFIQKUQ35WSwSwybOFcm6uCdOnAinrhOQCjeqYkCsAkGUuKki2+Pk+VBQYn1GHm+KErPD034Vom
dHwbz9SAKjlnLcpQzNVFT9pFekW5CT7CKVXXgFjTcRKoEaccHUWdfx8n6lg2/NUn0vzqtPpaMGqD
TNUpSabGq+gNJCu8zT/Ql0RLxBsikP2y5vE2COU4nXd6KAvjwZ0N4f/5hDV/gzu8osCEhCqiJrhD
DlowoVpqk1NiNMUIN15aZ1bmKo0QcCqQ7mqrXJ7y08epD9LsRjO3WaPM/0VTcfobOMbIzzGcr52M
0FkTRY5WRV5YeocGTlIvQEp7SnyGPnTYJaGlRIG019fQYCHLmstdWKD+TfdFNAGiKHl64yz6w+Gi
ZztwYnip5L8iaPTArRc4P/Ccvi6KI744aI0ykm7feA/O3YgE8G7afU56qqRheU151krlDIsAk63P
YpIttWgYUjK1lPpcJwJYoveWnvH+nO9bBQ/c9u5kvwMQLDcVN0EM7E9DwvucMbUs5vOKY+TPRUz3
OaD8zhC+624P3twNQnsak06ySyy/K7nj4cNrG52qD24mMQ1wYEbUVQ816MjswgNxyNoLjAUH37s2
+6Oev0C0KLga0fAEeb0jQ3qFm2MCXHFT/6T1+jEce5ZsUrxxrmwb/aD5IFY8RN6Li+rZQj1o8bNl
eEx5odft+jV5mf3DndIcXbtDGgGxHdsncqGtC9OPl2yy0zjkDK7JgruVdWhbpfzYVuR01JXqbg58
m+SM5QoEMhK/It4aCwfj4W/7V8FqwIMfhM8VM6z0hwSHlj5WKmHv7aAnCvAKRq8xl6JT/aCkVQnx
L3H9R1f2xdlyZ12qboxyEovBVM0U7lQivYnydcZsSziviIGkF+FAXiqRiObbfBXXTT51mvtmuFzt
vpHF9B338IHkWWQVPE/A7VohWN63lreyj8YDL/SLchNKE9+ioT6KyIzLdv6hFS8menl6nxYJkM7Q
oBF+g/m+wUk11DM/aL1td56W8hstIVllTkblXYnKdhlzZmuQ5f1ZHt9YCcAo1N+jkAG8nG4rRRBF
MtsTiaKNRqZnlmDTkQsdY1s7Q/FCqxJhNgs7MR9qgtNh9hkOhl5t5brnUQUZJszafQlzxiocg8Go
Slv7EUbpaBGYazjqwECDYdc1pDq3VPVqxS5j1EdbG2lvCU9aL/WXcrVGARbeBbCZwxKXudKqk+Vx
puDZl1T7mXQQZFW86FJn2IKmfRU/chTMa5u9laDFsY3xnoR77MtyNIazPdOUBsn0WdhMW4GJz7DO
TT8QD9dwhMxzxFV6Tgt6/deurfhiQ0zkSHDux1s4B4xNjsmtv/GAE59AoJoCYUvRc8M9azyZ71ct
947SPzzEbcyzcivJ/czT6QAgjknp4GDxveqfIFz7lvJOYbG/XF5Y+H0gBfXbXrCv8RxUuTmrz3B5
4SXiQ6GrPCoyvYY6N1h4xQ/cnurcyP+g+dNTtZTuIQuZaVCzU7GJ84lR4zqEZYfPM9FYcS7ypshQ
E67cLRHgLdHCaICD5FGR7x8Cm2USL/0rAScPrnBm/jPKo+HlklwbWZvs5x0JMt+xRu0E+bJeLnIp
s7ZSa3FhvRgJuYzjKdwwCpsNg1c2KtE0PLUZOOuYE1fY/d8sEk+0fdTcIRT6jU1DutmA4ZsC7+YI
b0EEWHjLvv+ELCMtrVl9dsJGoLANGr8ljRBWsOA9E36ou6VXFH7/PTj+BHgG4guh33pewefsLBoS
sDipU106FNhguwTE+ucUuncBWdTWYWtkjIYwXh/rO060tDfRCGhnCix4pPU7Y99v4Fge9jjvlccn
+W8Qu0ZCpz+cZ7h947khn2iKHwQmparuYU9SdUQT/hUu2COtNehS9lv4p8aMy6aVWEgfNUn7Ffhr
GqTl+OiYCipHXdLALsYAmXN6rm/tsDvpknjDgEtxtCH8o9odVG33vyBvyTqkoYrC13ERcgZWnlU0
BEHV0tFOoYpwFB0xmHUXLFmliT1hte0g00zmCb1yUx565f77XP0Zxpcm/qYoRMwJjSYIIj50sIBn
TSKvTB9lexWVaE5UgKxomO9juCvoqaQkiOz8JBun0fKXhO+8qMLEnzJymE2n0Tqp8OO+PsfhXnaR
x1neb6YwhVcpnl60CgSko3Ehz7ALjEeaH/qhr/meGkV7vU0WB3yc5Oth4G5nw/GT9a95qomYetME
UcAmXOe3CxH3EBRaLyq2+WtNXVoEMfTgqNBLQWUd6PT/YjIYtdzSg7X+aC5Io3SwEK0+letRUAoJ
9gMGVGHkkDx2uW5vaA8AXluuW5K9mGWXrKLIsFcDFyiqI1nBlJeZJHewbNZmJIDdhzXBUpWvUQ1h
DY5Lxd/snwS80llepYTFhXRCmajvwl/UBd4FG9eeDHDsqEvOFLRj7tR1w97DyG7QOFDe1PtbyfkW
N6Jm6MbPrZUgxasIOh7CNahED3bDeoxYz6krPhRuba33DH6M2SvnawB96Jq1btcVeeScByagQuDN
jidnHZyu06YcE/MwKFtA8Dr/TKEyQfOraqpGOuwEUQoUpcQEX5n7md0UsdKBWyxtP+7TcSdW/51l
hgkl2Mj9GDiNcPFoqVOxq2VxUBS4iGfZKjaHauEVQgs4+jZwPfO1VPDsznvW4ZZjU5f1yAFXR5Vs
cO6H9NTdIedSxXsD04dJ3wZph6q8Pjw1y0waMTGd4DI3adSVBhbmrxLdj03mggHAanq3jXNpo5Ia
VBMV4EwcjTDKnMKMjvnSi5eWcFITSWxMd+QlfwEiJmW68X39Hw/u1LuWGy6Rl45Q6FZa8AYiw/D8
jfloW2I2Y84NfwkXtVhXXlss+aX8uDSVRQkC6WhS0Y6wS0TKA+vmaLGOhKGtu1bhoc8zea51FsuH
cj1XebkJqAuqD8OwsuQ68Po9MEsFTRbfyIk3RBF1JJR+MQcc9qYOelAdrWME+zpdCBHw1KjAhN9g
EEiry56DqM9N2mQfJRBXGvTIuHNmGjHYRc/bVPBrI8T7MHtoSoTakckKc4lU0S9SduPdG5dyi2NQ
pt57aDkU2T+A5ZXp2l+JfI6s9hicQ0DApIrAfVsWur6RmzacUQWlDlQDrRi6g0tNZfMOnzDpu1uY
05aRD1aPYPelv4PNq/jBfSIsA/mgkr3vQ8DT6e5VfRGFUbQ59lEBp46H3Sw8HQG5fUUmC0NHtaEd
yZ1XbKkWhEvWP80QTVgekUUscYLz9DP+PwExvwavUzXttZlwl7MIqF5HNFf/FPdAwKPsH9OCZzId
2p1tlya4ueK97fgZc2iwIrPBT+dxfqXJb6dCkpO5s2KhpQQsHrHPeH3JlLo8MEjcdzOMItxJYPcH
u7Fi+VpfXuzxsKi8lpY8zOAIMbWq0zCebLlB3M3aGn6wpP4+G/3LCQzMXmaf0YspDMrPhnxWhu2Y
xhIYMd8hlUx2z09ffR21hJbKF/B8PZKPIZsNwdPlnkejykf0GPiU3RZc31uWIqKrLQlk+mZ301op
y8oTY9kY58qWfAWSn44SyT9u9cPRMcyrvKoHNLcnD8GI9kQt2pPpTTOs2vbh21aX7dmw/59h1Aeq
dDvVbk1RoR1k40YKCUMGHCznjVElkPSNE7JusgmgvPnk8/rMskEOACWcuo3ilnffMYyos5jAr9I/
ZjH0xRgbNk0r/AaIG4leoBfJUxP2jvhxQBzi43Rf/h36+kw1FTtP+rUV4CR/29GxzQAYfLx4DqoV
3ijJo3+3NT4ewLoftyVPMP9MYnp882q3U3jQtVMlJcDbHI6DDRh/PPRnoOdCB4vUIKIfFZWtV6ns
9KTuW+1kcsHzI/Qp/z+r728fiUBt/SPVT0z8ODSZcoDQPZH134gghXkzaTNhXzSsqZQr/Nt/CZcc
LMV15N+ASgEUKRlbRIUK9ICJZ04aa5icdKBNgqpM99q5QqjDNtwr70pEK7ZQLu4tPcQe3TP0Blqj
dbtzs4+oCcMx+8WoFIA1VEAuYMubrbep0SM3qGNh9qHX24PzJwfMDpa8mtRzGtoMJvTxeRH7Zofl
E6FKziWSLb2YATQoaK1IEJP9MyW+wPAPCb7d8720vlhO5RFAld8aQrZPVekahg9U8sJD/7oKzMfc
+xeUSAwRkW+tKOFP90kWjSzKetvBzQXscGmUYV7B7JvOYShV6w7tUK90LZLSYy3i21gc4S55LzVr
17GwYKEsiUTHiAnPJw1KISgS88Lt5JezQLfb+FmxF14puasKCBg9tL4sUKYy8NDindWjxptuSsPd
RbRsCDGXYoL4GUW9ncEmQ/kSPs/g+lESlURsUIwIcepws8RVrZ4LsTv77OV6m8WW7utPG+My5Y0o
etmfyVx46e2Rt0nwpv2qDoVvmy4KrZ9VIrrVRjiOCnnvB+WAJoElDlDJxJO66hxVRLAxQi5hLXDp
k9iwZzaTHb2nZkm+0BXp72LEv8blvtvAU44KEJQGX5WsBaiHVnZ61VWnH3BtnRCq/qvHE+G624o6
S7OrWbkpiBC1vusAFwJ06V/8U9wjx3OnZVTSeJxu5EGlWdt/4m4kafhvlw+MFYzspZMKUU9LedMX
wp3wlc4dgv3BqoUervgn0NmQ9bBGJMdj2E9Qg4Bbh8hnE3Uw/GOyT4j7XL4tKAMX/Z9TSWcwi6XA
UMOr/I3HchRq+2Fs5N63tS/snT8JE+eYBJwIl/nEtr6vdaOtAcl7WxuApgraDRpdU8cRDD5NubKt
5is4oGQn37VpQbIPoOO473QQywciOD6SCTxqZ4gN0jv1rKbbzAjSCHcZo3CvXnyhykXD7Dj7Ptzn
xCFIR8gnox/sgdy+ZU69XngGnmk+HnwEDT8tQCZMom73ja3BGxNjb4POa3P6VeYo6f61ELNF2knz
j+fYms1SsAIIjJ/wdAil80i5+IAVWx2VyWbsYYMYtCVZHv6GGWLVejU6P8ADFlvxtRSczpuD270u
mMsAIvcs8SAlrjt8gzk8YsGMB3uEqdIRBfN3XJwmfml9hJ9FLveZCAgZclXQL4wfjeREhVW57lEv
/b4RQrtLmX+UL3R/jYGywpNJui4HW7X55/yel96hAPe1ZQ6Agj1Ub5AL/CITiyAdu3ZG70M4liu2
FApIDCiPyfou8G6p3dZwmeBBtnlY+hY4nOWj8ETxnEZQfWKsB1vP9jK/Z0DFNwxDKXQWQnoY70NT
um693eNcAWZYV1lw0jfzytRpl0Iky3VD6PbltOop3ZNCcGUvC365evbNcN1yPmgMbm+vzxOVxcQv
Spudpm+A1X3ZyFP2pLLgU6tltkQRJeJQqMsF6X1D7jRZdBNBYUEdrRkW7YgODLFFAEfmesOae0vU
DHLz68LLl70iSsxJIJwx40K7bPQMEo/+JfduciM5wSw15n+GDPq5UnasEzhqIzOfHFRCfaerL1lX
LZOnvf70UNYEpFWt15/nsfnPRApGITD+XF1G6931QfsI4vzuP/vQd8FZ/Nr0MzCeiCwug2W7Geqq
j54IqD23R3IMXCITLlz1DcLrf7a37K8YwtMDkI2MFe+gmaJGfmMia48KcN4a4zwDCQ65IXIqsCL1
XpjhYV1QroqJ6csS/IBT4ZID0CRujPT2VWtv3XU0TrslIn0+brFH69Lbr8jSBzvyZMv1V0mgNJ45
GCErMnXLpJGt8Uj2SKLYuuZMib8pU31PHtjWMkVGrOqosposusZRt10GsKW4N+A3kifRx8fwnizo
WLUx2VOTk9Gr/5aLzprZ+jKP2iRqP+NHmKlMqL4yTFSKY4jsOTZVG9I/CmUTlB/3RnK5xIYVziPH
EHNqSrN/SsKm7oZ1j4IAWiq0lmY9gnRGkDGGOPBrOd7lj/fWJS3YuLSnNHDyNQVyB/RtaCFa5hTk
AvJLnY+W3a828Cs5qeE5dMaHiMunpDT5KO086HU2+DflOqbbhg7wNHt805gL8lE0yY00s/1eB5PC
kCskWySgxEgM+VziSt1vKQn9VzliuavKUY0/it6oryie8QoJCmXz6ZXQ9iEinQG+iKRQky/coiYa
M2OHkJbGRmh4aExyNKsWVmztmzrAVwV9fQ+dXI7hhX9QOul3qcfKmakS8Qz4mJ3Jh2lwRrGYGFbB
Kgl+zafggXblMV+BuAMgK+8zI4wisXEUYqF2Uc9bd0c4vAtykvSsxuK87JvhuuhlOYbR2M0rZUJO
Zv2+/bOOex7v2QT5xlkOuWMYNhexft00yFXRwin8XNRG24nfpykqJHFuH24w59D+f5xXpXnq92ds
HpwETS/U03O8zSWV6eeupaoH+7LC2yW4NZl5Ifco1dAhQd2ODQm7VW5HzIXQeL8GFkaJk7clVCxn
EyYcK+T4xGpe15I/4GdLtSMn5ZtaxXKfPrHDkzXMlNtaKZMQxKW8InUQkro/c98wcLNcTImfacjp
NoTJIbiAsYadjdmHytWFVnMGjJkkMzZyIHek5DgKmCn+wwd8J4UzY2uRdpJhv+jhn2PdgdGg5Ck6
21szbiLdAFqe3NjepFGfAhiaOBcFIgeZBk+AYpXILP7iA5yNLVfSJfcxxHrY8ydupZFLLVgaKE82
00ebNdIcn8vAkDrwk2nDF263h/KhERU8Di0Bo862xYXmeg1ZghrUc2rXIW79wtaTrvcWtN7unPpo
uEePkEeiE9pp9OTK5c4gZHANcRP8YcDBeevGU1s2dRbDpfsybiHDQLuJlqc69QTpSzcrdBb2L5fY
hs7yJ+C1zoYpwP2UDk1ft4C1Ku/04kQhOOoexFTyXhUBkmGLdl5aL6Mcokxu1QmubplpzDNnv+Ja
a2nOEHEsPETGi9RoSi3BNWdDino5cgOtg6MtPjfGxMya3ottdlXDpizQrO6PRiN9d5i6Nt46/c60
U97w7a1hS7bC1cRYkI5evx2+7HKnryeLpYFm4fn/6+w64wrOylAFbDM0gBVcpWIH+4pZZdunbZK0
I1qR5vMHjWO5tnt87Imp9pvg8GfSGeBRkw+MZ+vtOML0FTfcsf3Uhr50tY3dwUikoTO56Sqb+kiQ
oDVy5C004KPpymrxSeFOXLimxWpAaVDDBYxYiLex/jdx4JFs8sIPYq2l8guK0v1d1e4vxvMl01la
NcRiyaRdtUNodUlyEpQ01MFPKjIqyftqHHcinLoOP/kPCRkO349iRSwN34q+SnLbz6+IkFGpNIw0
oV9PWlxTxP90aWAfoCzvu31fhHbHwY1LPF+DIi4h8um+sGd/iKqqctYGalhczExdqdKEzWum0mSW
zvwOBqQfdWtlBYRQ/ln7PM7Eb/gg/6ykH3VD90OCO5q2N4vhE3PhgHQhMYitneUvxJbd00rofz8x
rJFwVcSradYTKMfvBUp21cBF4EYrZjtdN4F0ay0hMOGHzxFTAF2N4fpshRu1LehjwGLF3SXEGRbG
GkLrfaF6OtzxddBPBrITQ63qpjh1gXz/rt9i10GYyGcY+hTFlT2d+xy6r0zJF0Bal+irUYSyEAui
MRRerrMTIbDHdnCtUZEZmJLR6H4+iNRioQyLZClM4jo2291W4uCgOkyr5iz+aotuzZBdiZJXCTe2
TfVomxCWkLij3bnYMlD98TuzzWrhV9eDnoSyWD3M2ZmurEmJCoxaqEEZDQHcRO/qpESWLieb0c5+
a+sPmXs+tLDvufdmWv9eCOiOCSzQIpesEwmyKUkMgIE5vYKPU4PhfaagzicvdrzP4ADuBjf9O6BV
mK7FPw/A3jxBr2A7zFpF4UKjT3gQA05RifIK28jJEq/nfKvAVNf8Z8WFUCXK+P5x1hUI90GLBSsu
alzubbMMMUruAMe9mbWlPPidirkBVCS80EkUho3IrzfXpo0hV1onDextCnSNkA0LgrZS8I0jJc4m
EybrmZsIu3nnUvKr9wFO7UY9NjQLAr8bwfk9M7g7N0sWbMLlYOaTCI7wgg7BpastflzP/Nz0anwt
IEm6mw8IUmwKQepf1256HcclwkelUnCj8/iKWVEHP3AxxUPCiwsI3cEjZ31WOy2hmpWBESjURDLH
wMOEv0aHwkNy12kEB6pe733vAlW94/kZ7NnMWSYRexBieHkU2Cj80A+3ENV76VEpgFwXcJOJ5y+n
l9qvvUNuyJECElzRneP/MYXdIonYT2EfST/HA7QMRzA8gGYTQniWiURA6cwRUwovsWzAQEs/SNIB
YYSTAU7VHBAB04wmpwm7QuC4uNVTkelXzGduigisqAl5SdywjWXKD4XER0IEGiIkvj7SnbsGQnAm
GV6XCpmHx9UBX1TlCUgqN8J2PqHCEWkzubHEGL4DBhMr1NqUJhKsvtx6l/dS47fsuEMt2Lgoqk1i
YJsQZ7KJBSagtrHaAPmnSRNnV7jiSgxrooGojRpw1la9yZtx8l5woOOOYtU5LU2s5AOouuxOT2yh
wMBNytOZMGcYWTsyvrzEoGByyX0qk3QyBI4xKfKPi4hXfY6odF2AyLjGyHUax09fCvqX7qcX5SB8
O/+bSmYebCq5DR/JWYc1SwlK5UiMQlDeLuntCBWCuSCbmbTNIZI3dp8Hxiq79Vm5rI88b/W4DufK
y8/VTs0YEe3/7JMCuQejW3xjW2aDVSPc0NMRg5bUlQsSMRc+pYpULbtm7Y2R8t9LmZyCrHoP89LI
HRi6BSA//BkaFUkQ3/HPpzWwDDAaG8QbeHJK/zu+Xd0eeCWwckaddbCK3jj3C7vGvbvSoJ6pukYm
U7HPSBQh1MnNAcv9w29kKn4T5ZojG0k7kiPdrPZ+C9TejV//Jol0jMXP7LfkzXMxlX1/ZrPiSNcy
KYIqBKQo7CvqkK4XgCBZ9VT4atA/JM7u+/YLfXrE0lLzZ6/gbmtFOuI6aFmuM+JT3EpTNr/90Zda
FxrMgq2hf+XuFbOKqrN1wkYVBrxdqFMPpT/ik2JQg9KfKJmtWb9Se0JAK/MJWPCDLY2DvYPotEkw
ejVUMhvckMgQ7RJ73WEJTHpg04i3eJ3lTmaYYH60lJh4aYIvg0Op09QZycfgduLvlNqmCTzRSNqY
4XW76+o1sT11owzE4tK8q++/GG6tBj8ah1VFdBqHJO1n5YywWPXqXYER+UMHDW9vYuEC//Yg1xFi
MYXCNhi1csgwrCpqgst8pQYpmrHSynhj2tN46He6qN4TrfPCPmY6MTSIaflTpzNV3eLTbcnSQqTJ
dJJluA9wh6ObAafcGS7+nsVAJgIIEAwOJISWWQBV75fTIkY6CgG6JfbLOonMSYwJHpGPVmNNex2M
xDsKjFibfFEdE3pd1oBsiSlGBsJhfud223PUH6RYBRX5PZPxWnfh91hbhChSXE3RHHjWZwsZ+mFc
qd+O9mYqvys3vNOZ7DLWbgXkMaNKOlsLOEpLlO4U0Gljyk3D7i0xKov0aom67kPEC5AdOoyvRi+K
aCWyJE0+gXiZc05sPA7LmgVpMkd883DFcGOdfLQU04xBzez/WVeY+GjVJCbkSs78vvNCDnL5uErB
bp4WZ1XNtE/BQQnJcMBCLpPYZFw90jomT6Gcf1XPMyScYGmnYrmcB7EiXGNg9mEY3ljRwGfduZq4
+mOVedz1NN5SAX20EBP5+fNwBCtHcIqBnh4al+KAFz5Hze7lGMOP5VjWHpEIWFzLAJl2vwoYcR1Z
BYQc3/APX5+NVCevIUHnkcPhSfyvAMJvwmoC9NPM/MIa3rZc2uzsRsFuko8pPwsv+1PWjzaHYPLm
rljFu5v83svcb70WkAmRNZuc7DY/tJatp+EvkBRFx4dxrbX8eZ9z69CTvBz+N2SPwujEacKtC/hC
Ga1m9y6zKXC3PqbgJU5sleeruYHkN2rPPIiKlPovyr7tJW64SmZFrZ7BC9JMK6ebtHHXk3VHaWAn
XRMlRTkDKSVdrgMXJoFw1V7AEzdvLMJqE6vyCKpGKMp3NiJyv4911JCrJRyUr6uOmPbmHCekkbfs
+ss1jfeAJM5tN1uDcO5w2JPSPumhXXgAmMuuh9OjEOW6gCjj5yyHHYRNdM36xeP95dxFOQWmVLWi
Tuxe04YscQ8rdEtnui/r+LEcK0EVSYQ5YVcWL38VevPHE0hX63iWvnThK7FDFVB4kfW5XkrYvH+u
OYAcv5KswZqMovliFcvi2KbdaWD7oAiFNW45umBO2H48rYirCXwzkbJuqk27OXi0wWUe1NOhPdvs
ZXmvPsPVhbZ2JzK6mWd9N6Jt0JYCzzCUyXPCskqrf5cc2GXr1DuLJszlRpNmelanEq3IASQFrmzc
3z+yBBsv2uD85CotnjnYHj7LjFuOtTTepQ/DYmfPV4bjhE75g5C42AwaAlrM36Z7LBY/6B0GrwTJ
eZB0UXkqgUOU5s9KThHFc+r7NLsvSW4ekYIPdHwF0vmwC7KlSFsLQY6mwQvt4ApCkhSmasaKPk3S
lMSKBUfjVCLwYCBbiEaMAyfbtVygwcuMn7a8gVCb9cWeg3mv8h2LSTg2yFYmAazNxGPB0hXsVH0L
HEN6BdhDRgZKKf22QAzIOfDz2A1rVwiOvTtFGJFNUkCLQ0QQAc/30JPD6IW8auW3bbwRx91hFvlq
XaOQOxrnEvR8gqETDUle97SWUuC1YhhtRm6xWeWQdtcAMcwf1E8ZtanIHOT/3QJZSlF8iRPvuZZK
Y0uxxUchoizvrmBWnC0J5dl3s58qoi7C5mtQv8Q0T1sDFkKz38ySLk6QdIEryrlkqHOW4ox5+NP7
Gk/HFDQvR6kQo9cPG1IfJHitYjyZMyihQ86wMSDz4IcP7h6p7ruPzLV+xh6BP3jNsItozSnQJUi0
Q0mNSXVGNJig53c1Vak5OXmEBZ17/hwkMoGx6P5Uav6K38najkJV0jPoOobMDpPira60IiOUW92r
CKbOxB+DJ7SoFnCmSAaOJO23acQFJK+2qa+raFxjuaHOt5VHnG19iO+ilbroqED5F4iWgCZ1zDG1
CDBogkQpfVvLQGNQZsX0jQAJB8MvXjK6Gsa2pPSSDxK/Deeu0+nBPN1C0Ncs4QlKrZM1+Nt3FwGN
JB+n454xMBDmPBiZ/CWGz+tvfNVwgrA/czfJRO6lOqTGOqvlMkMBzf59tmkkeb2+X8giMZl8mDRj
/+BC1W1yJkZ+eQKTU/y3b0PNhMgiy//R7Ti7PqzPSTA545tc4q9EMwq02bZOm0A1dkupq4xunPz0
piqaNYQUSP51jkHjamHTAh8zTYP8ZwPn8nXBi1i5rKvmtTJQGntYNggEWqQU7W2yQOxoErwgx3ue
qR6Wx49m/gBwkwgcvE3cDMONnkadPOZoMIPnW5q07A6q91ecye2xJt5Mc+SwAAWDDycnMYn2RdrW
gFBSm5h2wIo+tInuAo0/QMCfvSs/sEJNUgBj1khLa8mbQ8o55jlK8+RJ9JhaLKrlTf6IQVAE0f6q
L8zYJ19LgiKCyJPzsfAWuXhlMVsIMa7zpWvbWBanljmjX1m8YPk85Jswi6sI9Mog0DWZ4xJQUjfc
cPa3ODuWJJsykxu5GY2z3V1ob6CY6Z42nN/dLtfhHfw16sPGteT9gzHtkvoi33a5F6F0dP4yaSSa
DEEvHKIDJYme/7aKCFPsJUitk8KYwac2spFah8c8quXh/3HUxX/6yDH9RaP154M3fa3c87AJekhN
M0ZdcwU4UfNcK5u6Lgb8x4Du23bMqHWjJJfhhOe0Hz1Y/Qgy9EIiv4zJeKbK6Ymq3BDcFRjKaakZ
6lt9cmpngHE+ngYij203GDADkeP6BtLHZlPTQwtOr88IVEnizGXUhJVPgOuZMu2al2RbNMCMUIwa
XRyplDZox8AnTmOG8F56xhPkiEZuZIbJBaNZJ6b0ufej+LQaoA7nlexGw0lX1IgXNJ3dTmWgNJnC
tFb7eYQArmPJLDE3KsZYeuljg3/C7vhQMOJ9eiDWFvjiafwhXxAdTGqJvnC+bwZ8z0uI7B19IMdi
iWeplBqJSyUpNS0cfkjH+U9mHQyOTBamjgQ8a2TqdKvhqizT5clJM62HbBAiBR2B4NZ0xm0aDfL2
sx6g9lVw95FrZSNBKi5jntSIxAnX3uOEaJByRbWXNcLXNKDhNTecscp0EaqBsjV8NNe4liNWMxhU
oDXP8XYA+tOjzbdXMmFmc0rlKxIYGyRzAZk8pN8sxVnyAGo7EqMpVNp7UhV7FPQHkX7OSyfdo63/
hhqrUZ4eHsBtaIJpWrzQ2rj90Rt0K2btJ/s15PMwq5DEeyS4U/1HCylIu+unDPwpS0oO0stVRfmI
Jwj49rztM/Mp8s6MDE5QDyO8Lt4P+x2+PUlUixWuxNHo7Ws5Td6r969srrq4wXuSGOjjMszbI/Cx
ZiPVTyvMuaDIc7Vk3C9+ccZjivbLRb2fNIDTaO/4KY3DRDHtpGVSxuHwEjhaW0G5LXmB2I2zo+F0
v5dqJTvj7z6fyiUfUO0+LJHW9Cec39KZ4ESivbmADOT3x6mQEy3OtotnWKYMZ3a+ih4eQKN6LgvG
VRHpVlTXZoaTToNmwysC0kXxPYGzSGIB2CKXIie5GydfSfDc2HzhNp5075rd4rPNWPaP5NIZ3ylC
uQJcxGdqIJHAExFNvQTPm49VmDLV1KT4SaZhEeO5GA0xFj3FsLZUPtKlVGAi7gPJDWhreO2lWBmP
0oLi9fBOaE1LhAdNgqogHIY9kxBrV/rUR4Uvy5bkhGjtzh+YnUN2uiuJ6Wk0C+WJcPCojTtlF7S3
6eF8L+TJasCNlldnkYXD7qBbTge2PuO1+VHgft+IY3XE516loZk3M7gVVJW+L8fW7qCRrmFn50o2
Tv+zle9TooeIUYbsHXYKlwlEnq9Rx05iyNmCSjwciKss3GQ70i3qLygu6WKKN94u+olJMyotCnba
684LMoe3qwlimNcrip5P8YfRcJu+yf5Q+KRhFhTaHSU1+X6Cnj5/aY+GCQBPDm9VBLQbQoEwEwY3
QvXhZLIwgAo34ZTK6nr69OEi0j4UcA9fPfthKE7vxyQAigarFRwbjZw+iNXfejij7FYAov2/sRFz
Ukk6MqPHcw49jjUCZZa04KkpOhlrkvhcVQTzipIdehGJEDrJfwKMd4tcvzuZxkM7X83E7Ql3l7fC
leOJilg4IKQzYoHk9efhIhZjiOxKvtE1WaH1Cuh3wrRoXxZ49OQBj6emntKH5DNBNFRGguY9kWNi
T/8tT6MDM/DC1rQ+e8R28bsKAiyCKeeWlzh51ALqgWHUVtN6ZwE5wwFhHhAyqgxadM9iYzOJ7GiL
hH2MrJeXkT+v3fuO4ty8VJGpJgZS8QMmIQfUQJHHTcrDAmdvYu+zoSqNnsa8knjHkVPyeSFUt0Vi
HVgYYvaD4Je2deWvCMw6T/qEyKBRdy+WbzOibP+j6dvMqiCIi3oe6Is3u3JUou7Ybn21MA28u7RK
XNUlyOSTbZR4ZV0TJNMXYTxcPpEMwf+Oq28bDsMPDcSeJJoMvSKcAXBcFkrVS+6CabGSp0cv+C/Q
xWyNWVq099+ApbthM3e5R2Eizl464QK38kE0NV4C+zYHMg7vn92VqInixYBbbirC6vR3LEqlHnlB
mej+zp/YF3N++5i0z9aeDNE21j1Aq1Rq3N641SbGo5XwcbSM25vI1GRNpurL5BmjwrfWoSZCV1Ne
fnwClS5TGcC9s2RnU5aYhexCYu9zcW/v6uSZqCZGNfq4c1LoknIVv8/wirHy17m7Nr+QjDFgKA0b
wxHpO+zP0syBKKLoE2Er9KMXOA1KGfGpevBrDmYQPkmOBMoqCztYcI4b8w7nGHBWBnbpxEy99uVB
TbGgPgRpIsVMKRpEmG39ErCBGjHhX5pV1oggYj8hdfcNk4kf0P9iEToy0m1MV4FBJ7tUX6T8Wjop
2Of/+WuZN3xPoYOqgdYQA3rhW0C5rPEVcN5AaCVPxKA5IedX4gF06RAHpMT+4oSno/erY652Ui/y
96n4ZT9eAaIz+5XxyXG3d5bnC7GXbWLUtmPY3BYu+r1LuupcNyIw7UTvc3rJ/XtMhtA5qob5WuIO
buSfqruXGqD+kx6K8qufFubhnqc47srUKeJZB/HtqdFhYVvvIdQTdLWUN4d2ULqCoNXyimow4uMp
fJOBj1iVmIQVD89uv20mUu60dFzMYtrY41m3qo81Qfq/T14yRZgWTCYruiOsanN35kx+lyrjWMgo
XhVTkSC9O5XF4nNZn3m/h3QnnRMmjJ6jepI6+OAXdRyGlqD9EajE36ROXhYVEX725Qoj95U8I6S3
x4FK9wDVJ33BVtcLPZGxg/iCRj9bzD3yFxd3+eTYs4JvcIZbUxzFBYznYB06Dcx/sZiIOM7KQwK+
ufR/pqpvl/ca39CpmoQoGnpqHYTlVZYw0QZGBGPjyR6EMHbAix7xCooJFz/hz5M6rEFX641EbMpm
kfxhR5AMBRVorXpj3T2mNkNlkuG7H984S2lD6j+WW1H4z878hiiZGE6i++I61F7ZorQi5tXzaczo
i0XCf+TDNKBzD6ZD542qVCABsPup1TVLo23OnCZ3oSLqgu2+QNqAmdJZV88Iakrt6nWjtbsjJkxO
ZUyKeCSlYOtE7OH7Z9U31THNr3YNwWCEyzvmnrjky77f4bI0dIc6vr/gluWD1huHUIspQ+T7QFcZ
KsAW4OsajDxO5Z0IVRvwzKRjs8OnmOU2ZETI+WJVaFl3qQVIWYbbjJLE7Qs8M89W1KQweEBh1HM8
Q/CMp6gt9FA/Ry0qsWPU1en9LUfymEzGJjj8f0SX8eKMhlaecarljBQ36HIQ8qNKVGvTCuGb4iS5
Rgedm/TRExwsVA4OmSPyHfI0yuk9XUDguemAMhpq0Z/m7OLnbdQhfmN/RwPc0X0dc9qNGZF23nGo
6c4M8XhOx1mh84tIhp0ijSL/i4XLs8fXo5PnIUX9U2y80tOpj80ViQmpD6b9dcXFiWRYYyblMtvO
1iBiYOK+TkNx0MO8xsMjWgWUMmqeaguMJmGosAi6LRNRB8nyrZvtknhqQAvp5dgy6YAato9IHwbG
UIWyhAMCm+RpTbkWIoA+p+L75HciU84Q+bUr4vBhMoQLMxGeD4fvds3xOcP9AdruEKjTdB2EDyfb
rmhD4Q1W2yNMhnbWdC9OGVl3WUNN0iJVcidnHB9JAyTLX7ZJd6E3TWuGz7OaYbnYXvrB+J8mnWu6
HaBk69mJrnKXjiXkIwxHGGwX/8auWakooeYt4e3OFYAd1SJYGQ0BrIBfrAiMy2Hw9XtvE46TTOMf
HbRHcUcUvtUKPIMu4xwyoY+D6v6x0bhLmnvSoAcZmmnrJt3N3Mu4/toBNrl0S3HOwt8og1aRR6vl
a246NGFNJdZ+oi6b3VDawPATEC1s6YJuew0Q2lAeN96MjosWDl0P7VzrWB1zpKu/hfKOqpqAZlw2
Hey8OdiSllRAsBTttfG4tYUm31PTODEUlKTWjRX2YwjoPyEsXJE4waXg0MZcvr0Z+Dq1K+/59ZDd
koDjK0/b0RF26dlbS2gFw7Yvi0EZNQEkEeiaBy7APKPcV1dC4j3g6UeJsnXcfQKOMYmHrGxdnQMo
PLDDgrjRSj8wkWhqUf1loXECze0xtqArHKZ3PhmzY6P4JVgndtgE7mBwxJJirZW/u2HKWIbn/T8H
gvgNwxURbhZH8Lqaj3hMi7zIENA8O4milg90LxuMcYSif/2XPz8BQgTalMBC+qXKa/UJUeyGFE9U
yKBxnRIydG8/LvCRR+oVHCyQP9X6Z/BCkg6bG2cresokcfLrDhx1oFsz1qDr4OhbrjnTv4ktMETq
6nmg6iDVbi5fYXhgkyg2y9ZfNrcOJ0yZ21xPLA0J2eg8mZ+nKsoh1uA99zkcWdhqg3q138deKzdj
i3vfUFz7Q+SoDnWWMtIGPO7lMONHNCHoQc4hQboJAHa1QyP1E7Uv9BMl4YSaddPk8petXO4CVb9X
Ls7HX2048qWAq5HTpD+U+JIL/VkaCq3Mk78A66PG8eIumQwMvbCMR1M+yqwNYYMmRVwPdQDpoEcU
NdjI26YwR63bUv7MYU5/6JTsb0Swhoy7qTpd5wKwWJMSevLkbtlcRNNLS0MRN4NNtiVtaBlYpyEQ
XHgWRCqf1ujQewfLf8J7K9lxdag3vjJk9KyVXJ7LE5lEmPsws8LxxSVUL1SpqlQSg/7zq6+N8nnz
UgEXbu6XKD49jItCkPMuxTTGREB34TDzRtOGattBOO5D5AGfS3l5wtupIowtPa7QiOUvkbE35gr3
cnfGhswfNXtkWaGG+40RPSODA4lXwHJoCTLVbvvi0+QIiNRHheMolGV8RyUcgtRBrbt0sqpkxnPL
JZhGnsM75tlNpQhlRNFREW2QtDTDNV14R/mR5KO8r2dSrmhoq6JL/QgoF/2b5ZevVWBDW/2jHNq+
LtODXYeQaXZDr1ybogbDtAgRgIJASq3H+eTBqMNhbpR/iff/szRxQVkM2Evqdadw/OZBiAdTIJTA
dw56f5Oc7415Sh0FuAy2YvhWsKtPqVZgjCBoMCrqKXpBhUXBM5IKlNDoQA7S1HWUahwM1VwA5iPA
xI1Jk8kLBovxP71GIzHksXP2j5JRU3xk/I7BzytstcHAAJCkYkDoYw4wpCRTKyJcI/4dnhO20ABC
Ors+xrx9PEEgq1kBWHTFpsmFQbIUSavH6Ty65a+Df8sZ2K/qFnT2daNqGM6R6b7TI8cwIJXO1dj4
NvGclGPMgW1NoNufaD/XuqH2DVszYusNr1k7uk7PbYnBDn+LM0UV50P3XSiZ7tJgZO8dMaPyEfnQ
VG02QyM9dEcZRkBedDYmD/4VIoZDRm7JVTgoyOJRZzs5RMYO72UBhlYKjhX5nzBoCV6WsrMEFooo
QTt80fKKxRrQVuWdUO5t2uN39L68Go9gJFWPcVGYwVdTNyiRm8iVMc8TtPSzTZQHNb5nEsvgCL4J
5EKPrh7TNo0jqkvXIAd+E5EJfsGwrlnWhJo/6n43de/dNIpIzW2sfeZKLdlft/oCQUBg7AzGLOoW
a93umn1LdH/b/E68zcGwyyMW+6uyMJOO1k1tErDmHB8CC8XLnXJNjhwr6lGqYQc0/FXV2UD10JFe
S9XCFF0ZYR+ZbHLEkzndcD6DDAA53BA1wvvFIv7gPHsn90lv9Vrh65dP31O+f3t1co0fqAIsS8Kw
EzYA5ssrUIYCcbVAYh8jzhBeWEwLKsONKi/gaEO2keHOFq3efg3oYXUK1/ZpckPn20zKGH+V77A2
xc0D7NTsmHKdnRRz0YI+Iuxs+4K5MLJWFjwoN7CLF8yAFSZMKYGLmd4uCyZgOr4psXklm3j0bn55
WibxavbD1okJjY7LodTpzjC2f1HKHeVDjGiJGGlA7/HEOsBK9BoPqnxVhsvr0AJX0yTmJY/5nQYJ
/uaPUsDuftrAL9Zbg9Q13Jb3YG+UKzo4lRit/qu8mXCQdI1U7WVmStF6rnSWIgpz026/MW7GBCsj
U8ZMPyXGId3UfvRbJIkfS0b4TbBX0Wwg3jlKK+qvCtiedzHLBdsPlEnjW2KS39LCRsAqQJtcw+lG
0tZhbn9a5C+0uvS77yXXpTPiDTXugu2DBiCHhQXM00P+incFO4y9pIvmg9CsjVeU69y/8C17kcFa
RVJNWeUISxqI9/Xh4kPS+IU0q6Wo7d22KEO8fvS67pCKPKPXoCnk+oVsn66lN3AUD8j9SklRqYth
eoht2EhjF/QBV64evLZCdtFTeMvcxgglfjo5hsCGpONXOufj5RqM9ECWR2cFuqsLVOj8TvonW7rC
ByLnhRqLHlBwgvRffF0e60+BNlvAX1kvwiO+nE+Odc/3ejSbc/OlbaO+qMaFXgapIeu7YsI1K9Vq
bP+/h5A57YkuphTy13gJpDn0t5iNfoEAo9rdNk1Jaj2Ko3hLA7HvFRpzHvZdtfKKZMPT8p+bqUJM
75KI/zzPTOZ8K9UJeZgi3KsCeTcu4zQY4qQubuPR2v/QN6cbR1B5eLvWdda9NAOGqW41jcAfMG33
CXABghT6BptS0+BQozrDar15YnjK31UfwDXfUaFqIRIaWeocr2UxdoCfTgSygW+2NhQrcFfnLjRj
X+Pqun3vwNypzugHlPZWimd1e1XORHR+ZIcW8avhN5a99PbPCvIbsfdHJxjlF95mW0BIxAKUw4g3
EO281mVSyQkG63FZbwEkgUbx70wXFhyHVsuzMqqqAjRFuH7ctDOGUxTKR4z/IsPmutKwayyc7xmx
9DFkUya8Q133AxuFG1Lw/7LDcttbd7FgXFqPpcikCOB+uW2NOWY9+cazcKGde5GfC/qBoNQKhPUU
r5HE7Qd8PfFfyGYmSoJYU7S2lXC/B59spv+fx8bpafeKWUeyyp7Lm705WfGVN25TT/guVP0eK+Gv
ds+xOhqEHudhn+k9K1kx9KAaU33nM9Lh2XwbEj+/OP1ZlzlEfNH6C3zdoKpGvbNtgKG2ndy2Legw
RaxDgqvGRxwARPJI1SOUTHNC5nyFpWRYUBXipjw7s6STNq+lbZoyNkSBKsrBF3HEhN/ePTR7jayl
6jzKO7Oimye61msURkEP+anQeeT2XSK5at8vy/rv3uOCPuHxUKchGrmRy8mzzzN8PMGjt4LVx0y0
eCuV5Sw7q27RkJMRPN9LCSszM7M8vhc3tRhTWVqdvRIO2qPRLvmqvU9yvUH0AZqg8EzB2/6VDwgl
RhAG/flYo+QVEjfSTE7DPMm/aRm/Jro3iQqj7MpGEAJIgeBLnwZwvafkCgbplujsBofPrLDbdvO6
9NBJZ++HB4L0tApND2sMecm8gYdIvocsBuMxREXYJqiWzHOZnO1Lj7h5xIWqjz6MBIeLwu0EoIjy
0uRZ4yk3MqJfzqzGtRqLPJOaaacFWBWWRBLfrDssV2wAhZ248L5Krqcjg5VgSsw+LfSudiDLcD/D
GvQtKqnJlUMhgNrblGNVo3boyu7oI8wrQzbX/PBE3KF8VUg53aZTfAesEe8jg+qXkiEvtFlf2USt
KJpwhF/s8c9fHQbcsDhSZ2ifa3JxvJday5Vg1slyFyIQqQr6tLzc7Io4wUHtG6GmZuR0C47OKsG4
tW1usQdJFYQk/SIVx2WaQVAOmVzmXTs+foNDFoODmaZnT/sTUTEQWkte6fnzWCbEZ9z/K9lFI8Vs
ao6hoaDzEgEfw+8bSDYH3XOWabrCPFsIhiUvwUitekuTYw8faZc+8zfeMi5cBGYmUxs3jG2etuiQ
rYJrv4oK+fqOwEY+SUyy6DVUQ7CDCRYMSH5bnZyjkBsypZuhMzr8PyGtZNFRusOQ4vhtq+yy8w0K
LkdTlMBaQuLPle6+H8ubGjlzHfgb1dmoL8ZRxXPYpFIlwSYJcyO3x/nYaoKpsrre5ORx+3yrgePH
DsoNn1CbyCrBZ+cnXJVXaV8hBVI2e4LaAQQsAcg668bI3KkUbackLl/tUVVlqCwdehSfH/cRny4+
5gYHRRHRncnmrzYIT28K9rdcIu6J//xAlKaEQ8yffqCLQdGLpAjj6OG5C5DuszQbhNKzQU+5+stZ
czgrkGrmG8uQW4viM2YOaOjwRyhynrkIozf/j7QsnISCguILlsSKTiSdMaqjYgKIfNnIYgxxzmuJ
0eXwgaOjJHCsJcU818lT2uL+5DJMaf8Ct/oVPv6WrVl/po5kq1T3IkwLjXGHc/CmmLw6CpVoHA+N
EuR9P1nggFG5Vlt1KKNBHUIFWza1qWA54gS9nBFKSry9WwVc7ZfpQXTBFX7J9wBPCwuwd+jw97mx
soAEDNazLmGJwY47FAeZzU+wfVSwQkUqRfTCU6K8mEUi8MxOilwccXjYDs49395IvuvEe5eKclT1
B1kVORfOCgGAzxSkQTuhngw6bKirnvy/02x5sde4vmWt2pEcIDNiZnNZos1uB67brfGZWEvyb6zz
1ajwPFSYseFyUyAbDzKO4a5vO6xJguOnWVqpwVMUwUZuDgXSu6IAM/jxcpSL7EeoildpW3uWWpXR
mfLdpNQtwaoPEfQGo28TcS3nzCJ1DfTgLU8pEUYJUxXZNpoVs/5CL2mdKxwy8ZD8jv01pBvDYHfx
dXn4j3R3GyLbgLUjVDluho5XcdKVYVHwquUR7HwQA3wJEvflRvG5hULtijIAXJ37PMPNDOo2nXBH
UvXVb2H2FZffBK1Ces0xzmLrVkXNiZ1SoRgrwkdgSVx17CBwi4nv4dQYxM/ReKiILZ/fu92re5iC
k6+BS34G6FVK/YqsbVM0iqqTANzu2X0WFtfnzG0b6utxMDZUfOjjz5N0zub+ucP53gX32W96TlZ8
s+TjJE5Raddevw2v+8gZYzHhW95eCWOu6FFA4GefX5PSHflT6hyjlqk/j9Nq074piSzbdAHPkRyU
1G1/doh9ho7xJNxDPi5UdDxMVz2L1R7lJMPNqUvDpFTtlv8IYgLdmMQXVf8AL5MxUaKtcK7fGh5V
HEf/pD/0EQcGpndct4pT0Xmkj6NI8PJdWyD1ay3/SmlrkL4Xu1MVK8moSPAj6J+3M2xbb8GaHrHA
RcE8eeCvUJE/oTxO20cAG2rZx+Psg5pjYQbc/LEwi4Jzu//4OE9mTOBluELteS5g4CdFpqgvXskP
XkVf4A7AKhACz1ZEenwMhatyesQyAQAVlt7U98H0AxLw8o74eMeoi+9XwgKE+VZ8pzQDJmn4JSjY
Owl747X272IbeG93OlOQG2VHO2CYYWn6ETvo5mptlgAZhZgArLxUUCB9QQPrrU1CV7kejWKOTQTh
su/pIDd6DRRzLlgaRVmYznlT79VLLJi5ZNDvckUu/byPoWhFCRPza9U00CCNsPBD4EQBXxFChB+C
QVhuj2ni5ZCQzeV3fg1YYF7cLQv61mRkDvwWWQFNd3OtMbjSr+xK/bXe+oe+RUmpna6lDdod9O/T
BS86BPD7c2cb9rb9VKvQkkkWJTSL8chrLiMeFacRW2GM5edAVJN+2rBPMZMrwV0aJrZM0lzGx6iW
+U3S3S1hbc6AqlffutDDbN16GmIxwpLNU3NKgkD/iMi34U7mw5SRpV25qAx9x54Ldj6gw9HZs8Ix
PQ42RNgIALZcNAqTk039Um78SNLEV/iP4bJ5Q4SODP63LQeXYG50J5EjBNcSsq0Qtp6s4e8FUziW
aWfuOU+kFjJVqKa5Z6mFm/F8iGrxryk9noDQ6CWVYPe2cPnmoVQvRSlwNIprbf5AdkuvxeMj4V7u
uCzPKi9O/k1ae1meY3qpFK+iLho5S05U8C2PubqSzijuij1TBKdIQRV0GkO5b1lLImRLUTZERUH7
z01uY9cR8A3QzPU9o9nr+ReWGqWbo6CwFoxCP3mfQacH5SbwtX5OXXKBJgbv3ujj04uCis3Js9kg
WPcboeDJoWl5oufD6VDZrmhfT9jbqbJxdxON8LE/1P73jK2/B+HHp2bANTLRcqu9RQJwOmb4WbAu
tmeL28NsOEKfjStJMPrnucizVXNB7XuBHq84hlYgkrbPqLW9jVEkCkrsAlq2I5ZsbX5M8hqEQ74X
4vuhnzm8Eu8SOFl/Bu2VkbhZajCsuPwJXOI6rrujZUVudRqroiZYVgDXk4PxzbNkQ4nonj32wLfr
rlbI3xaR8AbpNZC6b4U7m34PIBvGoQ/irRwu2R0wOo7zFxcVfSODjQnE6yK+Fc7F62HdDUKLwzcf
0LWkjsKRZ4CsIBGVQ0yLJh1YoFnhNXBk8BlNucEKZELBG3Td1eITqN8KF4M02leQb1+QMyo8RTlw
KLcxcHutBt9axmwEgXoPGZi2XB6M0KAYXXKGvRh5HOPzwob+g2N+WpP0UEWzkCO0TzqhuCcNQScN
Los7tPY5KueD7iqbNCDVgoZrfafuN51WyAuWScY0pGYhN9zPeyVhWpmSjx4TWD4rzA6KDM/UE4JK
8/0BIrPW01XpKSJTp1VG9OdD8Q3uj886/SrRmiOSNQqDIY/DcC8yyLQi02XAhcU+jbk5DCTC62zo
dUb+rujYwPSZ63rUMy6qFtrwLlHdhLjm7LxGJzmA1DpybAlWikp6bfzGDkObZ+imbbT7GaRIJgMN
iOrCvl81Gj3N3eYq9NEF4IvIkO/3mK5GXm7kQQmCx95OqCydw3ReQte1HNEhvaRAzNZXuuqvI43o
DkimULqIjSLPmIMFVgxDdOOhroGLi5r2W4u6htAgPkITIO7ttV2KAAGFnjDU3ezfznjHPXfcAibZ
nBA4q7WfRPrkYAiH87EcoZOjegc+XpPcqv5FK683vgWfYsCV2BixuwUwb2vg4izznwJ1n/DClYpt
kctR3x18SR6oFGGFnTHrW/2C3bk6sRlFjbMj5/pd3Ef6159YWBkiUaYg+WZ28/h1aTuMq5pfU744
5nwERJsK/ITv6msb981v70P58Nr/DSLRDRc9q84dtjlTqqwx/HvQoyBRJK4/s7wfe8x/Qcq47c8A
qGGqHuHXDYI4SvsAcR6vBDlv+aFsKiHV5dvnlmZ1b/9YGgpk3QIS4xDcPCOqhOj0HBByPyqnfWjp
KKE0GhK7nYKBNkybFSZ8mgeLqSmIJ9ICgvpLJEcnFsL0p1MiGR4OKBakbHbmDLPtzKZiSjGxTbVD
LViXn8FwUCykwZsE3iuWFU2A50iccx4vkBuegXMj30darS6qAddn9UrD66gy6LO597o0zwPh2MW2
RPu17Hul/o9AO+VhiPLtNFcvURmeO5qeYwKdU48flI3eLM8u2ucBexZ+wxZEmfl4wMrJiMxAeiT4
7rexY4YUJu8VIMadoRYv410BvBwUUd6yARV6i02ygBQKbl3bJn8rsBOF2+v+rLPk5lAIUUkBnaq7
4zRdqJ7tAG06CyLG7qbQSinMyPHTtr+54/YtNobLh91Li20XAOGfg4bvsv3R2hWawN66FwSLQS6O
hVHHRzfGeZMG+K0QzaETiDAYBPGqK+RKn+0HHVYRe4ymZZb993GjJp7hKGIrial6nyVVEwUgbhBt
dd5rY39qWSRDXYEdorJy+eesXXeJe1BRHaRFt5zN1UpsyR/bqoR6T0nrCTx8jpIUvyWJxMzZtbi+
FfiBCe4LD57UkzHLS1A9oKUMIzKQiORfutCaZHVR00qVIGK8oUnGxC2StsmF8mjuw9i6KTWASahe
FFn4cLG20kRo/8MmPB4l9iDoJkHjDBqmWnMJo6RNMJQYRDvAza8DMZ5J7tS/qNqWmocP792SY86g
AlZAr/xxVCeDv4XBEt2LxbTXeOvGNyePouczgEQPM/4CgqFcn7VInu00hwuIwwKQW+LdD7cEowmc
I6hRbsH1Xr2SKbVtgnRxg/iR7K3asW5m43CEGwsTG8xiAMM3zLMqHWzPamepw4tXxlmZVP7XVF4l
EBHIYoBCeqMQ/ENrxTTl3ma9cX8eBK/hcjr1HI+btPkKPxePyKXU9cMdDx0MXeaBFYlKfcztVu3e
jZOCkMse3eoccLshkl9EeTwB6kKduwaaUCRW9i7sX453XoIG8mX4fpO82a2qGEvECridBzHvhB85
xjG/zScynMzpXOSjnrhqq7FgewDNu8N3d+GfBCcS8LO/VfgM+8ODsEpFbx8cfeSZqGaY5rDgZKSh
xGQ2Y6LK5HMZt20HwdjJE8UDUvJEAhtTk15bx35kKNbIacXYZt4AJLrNmhpPL9tuqbua6Ui1FndL
jfPM/DzeV6V2QoXASSYWlDEnF0YHPFalSL+oblTSWOv3jiZ1m2aHb9mh/byYrqrCoEBgLktIAxPy
WtQtINlZ6Ydk6IGKSzLe9Oyc9hQA8X+s91p3Pr8GOzTuO6uXEHR0++lPQIj/ZVxBLp97DixZVrKh
typkizRvJsLYMKjUtmcZTudECaMrpC06aV1ZcTjrqrdQrlDArzH772Z6QBlC7lHPyvXNNbIvJ5oL
431CxF1RmJWfOGpTloxeVjrMchwLA141wL46FFDzuNeASPi6neVGxVWiwEdJ2z4bE/diz5Gs3s42
Jw1gXPNwgTvB57O9nSbt6OCtaQtTGF68nGleKbTGrHa4lanMMQheU2aDTKqBpxQlT/q9CmkRvWEB
KFcIxZXFKF0DrJKDKXrkAdqH7tM5AhTJ5yft1y82j5HjXDbkKzm/lkmXN34XXYm8emP65ju12XiH
LMVpEAD1NM4ZNdZe5dGoOLek8vg4xHDzLwhRzwKiaGLo0txR8T8WNMru2uHc/HY5F7N9mQq9w1+f
nrx+TbIBO59/BlYSBMMNGHCRtAJKtUruIBx+zaURi3RWxJwvHBrEMp557E2iCkEO/QxZhD2KAx4T
4ifpIxJd/Ysx9GbKqTvqIkLiXGi5n4rpm1SDNY5o5cmOIsEeKrgUhgWJ/NHZeofd6X08KT7AW+Z3
XTL3+dfLcMYW8sKqugbmHfb9VPqI1XAdCMF8GdW+eUowRTJByuee+yeh4w5Am7etJLSDIaWzV3re
flHrsW0aZJCsnt5Yf5+iIV18jrgf6NKexFlww1DmyLeZoymhp8biteZgN7nEJGlQVMftWdY4/JwZ
djz2dKRfdM+Cjc4ibtGRDUFp0y+tiWAjhG+nwAw93WEE/3jLda9dxUbFvTxkrwpedseLabkd6Kd3
AxcEev6poCKMOjuO1td42tSBr2x4W85k+c23N/CLmwkxtfPDJPek+t32QpsvUY4EpBmmuPLlH0hY
2ZatxpPmsHKWoJg91btolzlFqN/UZ8UVMGrcyqy1c0pGWmv6sr+Swr2EA6WIrNStK4lNt9GLU3x5
fJKxQYn97wj6+Jt/aBh4TDOapyX68xP7mal21b2dge4zwcfP9oj6ZVQbeTv1hAgMhd+TledYR0GX
6ZCz0nmMudVZT3hvxk3Dlv6casHuHHPyl0172rlHLjrTQHRmstjXYd4ClfuA4ebiOBF7SZmDBWqX
3ID3RkSz9706wAucSrMchqWzzzApLAzgzht13aJmgALjKrE0wz3y9HsqalwyH4CDyKhYl8EefxIM
hPDgMWxkNl0AknZohhuZZjisJWpnugVJhkIVeiF8wqgcao527H/Z14mg9mBZMu8gZP1+HODJ3i5W
zVY0Gq2C3Xg+U5gmktRzjFce+e8xa0030dQ2ySzHuIMjeubMWNunevBNl+OlScZUPe83ACTvuWWu
d3QBVJGTI4A2lDtL1J9SSbRvrup4n6FsN6/vvaDnB8K2JX/llVZcDtCP96wA1MbrwLjaejNTrY57
8MKSm/kFPUOpLBo3zNiAU6eV5YAnoh+V2NsBsgNEYxQbp/sadixLnyVIFZ7hCZSiF+/NDrgtcR8V
2hHCwjUBoDohFLMc5NMOGr1sK1t9atuOL8kD6ugnon+2x+niPp1T7+0tLMMJlBUndj40MchmKUbp
JV1xdMZxrWe/a1uhblNm11ZGf5+CXSZ8W2+OKy+M+EPXNztUe+NtlKnSNR8y/u253TfbaNRIfdGB
vxCTuq1LPY4+bjHN7pTLgj/75DabYZ0Yd4BDTJqpuqHA9ksOKj2D2gIUjBf3PrgOQJQGxQjOLHhB
KxDNhhybBJaylgXlJVoIpIegCRgqJsoUBWZBKrtAoxpW0UgzwOJIfxLbaJglnKYNPwB08M8Tqzl9
v6wTTQ+hIzetHIdSIK2EbFWDUiqD+G29IcysY1c04cZ6MkFXNiWmFcj41wFunHHn5rTsVmRRJJDf
sC9ivnem+0MEk6UadLsh+JuhA9jeH6+SbLCED9ErNL3pHvqU3f/CiaMgwi26W80CsgdHc2gTZZlh
2HC3NuNNOeLJpxgwsegaM4BwVtBhK+YPp5/3638sajX2LJVkMrFo5PKpLVg26xdpPFMc3NAtLzqV
RqNnCiNFmtEMLYvM/xLCnAWMtrpT21vCupg4XNPMDxuFX/gWe9Q5sWjTFtTR5nwRpWjbouDTueOm
MYHcpq3+oggsC5AXkwu3KuquJyngyevLF04IsgITSbTmdW2hpeBIlO8mqxReLaGDfah+lFBWmOLD
+6NMeL8v5TgYow02g3pwnv3ZvK2FWBKOwGROegT0VbrqM1u6ARjeUz66uuhQLN1Yl+NK/D2qFSXd
eDW2HJSJBURD529qrj3e0nHxeCI3+gxNvw5DC+6c580jgBZ+VvzNc1pSbOhRgn9AXJhwpY64appK
ugKLgu5ZFCzMRWVrMMMhpxLP4j0cSq2zpKKzFqGXNQ4mNoW3k/qz9oXTZISux3G467vmpfEWR/2s
9+wkNVbq0jnGRyBgZFmZZfHCWHxBYbb+5VgyDzv9P5emiX6nhEwf8IQ9KO4p+DT+WSJJDlqNXdVs
4wvgZ8Bcn0zZfjFyR06Ib+EUMAkPIEPqtLrEyk6AyI8fLQhXLsic2vAIRNuj7gqRnx9rqdjtdE/X
admk5vc/MUmoGCHeceKPuGHOgEQs+rP6ewNQX144dgYPbxHPCc4JVDe2Emnzc/EeUTn1zuxsSZHs
olKk/eOGnbFaDOGq6iiPLrMmTcnDx7G5H/A8Cf3389nIGekR0qsUzi+LZJ7Y7QZc/21FSOAorIpi
pfDwp+/L5wvTjFgwSzdGxPPRy/m4RrKjxiZbQVOFg4dJzzL0st8NLui1lIaigsdv2MxAYsSJ9AQ5
TEoBAvPnsWq/bv6eP4djdCFGE+rUy+qSdGdQYjzSfYq98y1FyKG94byoQfXLviY23k9v5BxsxLrd
/ZlOEUNR5YN1+Dnvyn+f1x6MMBZx5TApCxxV00nICSbbS03XFxVXnxoYyXC8Y4hkPb0JLbEKWvhj
m8rG7q+H5M/6pDET05gSbEsXgWyMWXorTK0FjmYxVXyCD7I6pYs+bBmG2r5M98BMGqOg3teXGou9
Ky3gQtqojMwlqRFqT0zI5SoO+GX6P8Cd1/BaoOVv52XXB2YSoZKxYhNqucSRg9LFRyXhsuXyhi+P
q2qJVsIz2XrTxVcmwEutewTx5gjmM4VglCbQNh7hzdd35tXRJrl/ZPOSz0lkWNJueUjH8DNTd6u5
giiBlkuf5Lp93BbVcm1BOBSVfFIBHn1tijw695WUIse1X8G8hnr0skVrjTbtIXieQyyZMk6ufZ2a
emlSTX0KmoRmA0XAC/hyaHNnxxHHUbqL9Ma423VJJ4fLViFruEsAkoXULEol4iW/mE6mIMIL/2zr
Ftps0tL/3qlcJpOtvMfU/iFqnq3ApTryoY2h7fTMgzZSyyomPcKi6KP/06f4vXE3HMPWte2Z81pl
IU715eIsYdOJK0Pt6Arm+D3eDytWs+fDsTR6nJS60ivlOjiNnOijtvvjCLlNrOtl6OpLnWmHeunG
x1A5HpOs86A/eTr1+BgdF2O/eyTyfUh693dYMdGJPhDThv8m9OGdK6AjM0geRsL+csV7M17ZFORZ
oeNEaW3hLWYYvcj06VsHjAUrCQ6TXBieS/pxpypsjBXv7DsL8HWosIP3xEge2vC0kZxqBUVxffsD
nCuHd/CSHW93H4pYrUxiLitjVkLVsA5T0snkOoFn4kcNPGLzZ1BsyI3Qq2tTmwuQqDgydSgbiLmt
ojZhPlxSL8RnZ3EZoAI1yRH8MKdv7VWY/rLlcTAdO5j0gABYdrEsVl+MTRqWokh4n87vKWn1IEZc
yOl+x2tfBI9Y3e4p2JiopVbqBJn7UUW3KCdNq81Mur1M7y3l/g/P02szyL3hXOZA580Xi+7ySpDC
9L5nPDRGyVhRr9vxVnC9WwiLkvMD3uk2/HEOsKildtGwloFJHtJrQf7FhXnNyfrhWGTI1mUzuyes
XGZXtzRWk2GVdOQcJ57h4ARWiT63ou/MtQUQ9iBlzJDDtb7hKBJ4OJybASCulnX0f+pVp80A2X1N
56SQKl8tEfRhDIPNwJmfcSL3Gie7HmpHxiBSW51bpf2JGMWr3fIwk/aq2nD0ffnx2eZPNomTqZOX
pT6jsigzpQBVSl1srEQq0C4YcWfxTsQTUCFSQxGnN8HAI9M15VxORISlnDCgyxERrPMZv/DAXO9f
euix0W36xasW7hHH/46z2NUDCYk5CM+UVuvanXCFpi1jymXAdTpDADC8mgJAkYODY+SViySYBvJ8
fYLKiTcpAGE6WqnsWtyuq5ZnmMLPXwig00YbSZnjL6zcmNU06Io5zj7+if5NPPRy7nQ5dq0Autj5
SpAJnV3lV2iw06fKc9f+squ87RkzU2HW50K3Z92WbtqXuulB11Pli+LCGTc/UBhXe4PNgDblq7X5
5SibJN3pAJN84JHyMYM6FuLW7ApmCoOZOqO37L9OgJjYr9L1R+sGaKd2YP1U9U3EHlC2IzAiQnfm
TjKav6d9cBbHiTKHKmAcI+D1KEkVp10ipyslCVIq177ohYbfF/1A/uVPOjMGBFZtxXp8PrMSNF9A
2n150SKQRw3EJWQcMjItEncSJAbFd9Qs1bHCSw2gIid5Vw82CRwnLn599yRibgPn+f+W2zsEzciO
aq6xiIoiKspejkvzZQli24yi67oyrQ5MtBIrfhD8FzdN1ZXTACjaFtD9aOKvm9lzyc68KY+5gmXN
T5Kj/wdmMTBLYObtpyFdVef7YuWWfTKnhIJDYgcm06GoHdUMftlkvDWcJsjPy+Q+T4RxoM6kdpd5
z5hNL2LMUxrBaBEYdnYx8YhMKee0gilO8KggQ1OOR7peeyucegZpeOwgzAd055m3u9hP6INfDvdf
gBC7MyVPBHylfx8wtIfBcMkmkoihoXLQ9X4zedI06EFoiG5il5H8S+tozrJ5tSDSqtuQOaa4s1a0
MKosCKu7sEuO9QwStNmBzhaZ6Z9DI8T3AIf7JDz0cfyUYMFGnCSp44lI5ycw9Cp5D2up0UPGzvQJ
nvPTSnjHTndiXQyp97C84jNZRoLpgFL7FKvKh4rXcct6fsjHDeLH7H1PL51kvQ42hEkaqAdKQDYz
4YctIZq9g5/gyI4F9V/DPCymZojfEpeiKXNPmiHJ42Kro8hQwZ3u9yLccFRCixE0wxjpXKkNYDnn
Fwbw/vfTj/rV23OFMLq8ls1I/tQO3njQ9EZV5MpO16bE+2IOogbD86t9Plbft5w8W2og6sEunAOG
njaqTvFuD70JD4xHcAqOUfIqDnjNYC/bVQyoeWcR4QG22pbUOrCRoXMcKdQjTZjISebMJ4THztmC
p7llfi4QzfmwLZdcybDgCXWi+8ZdfpJ4vGo6GHI7uiJjnf5FwXj2kP+8ejdQe5JHb0vJyObw6CAE
z6L3qEp/CBj4lp4dDET8Fi+zn+FSOMrHfVkwNcWtuigz1Q1gFHGjHWz3RyTRPQs7c1BnHQhPNgGt
fUWua3CNeSSX3YyNS11Dsdl1Dv+udydii6wZ1lba9LnvJx4jps/AUGlS9IzusaJDe41suAr3HeLx
75gzwtBt0NJ7rvMI/SwEoP4jcioXKyOhjdNTdsURIapd7Y58IKBp6hLpXZYbLSBytLGo73pFwUps
wH+MIsOV0FFyYnGvJXnXXAKjgoJGFGM9S636akrdtkSDGaBHIb7KP5E4tzaCJEoAIkPtV2opCdG/
TIsCFnZeL6Kpi48fj2z8VhlHmOrth+4i+MsRgujKCN9MKAN0AqGiSt5beeNQMM4jHkmF4Iz70Qn3
Lc+ie5EOqiqReSQwHjYfI+pj0a+XhyUIoVJXAkaW4VEJAAzDI4GrSyh2z38PBn2kMn/qYa/iOU33
HMYg0qfvytYrS3HGRY95okpoRy+n3qxkjGnqq9bN658Qfpexm5zl+MR1lL3/4r4rG/ezZ0jWiFho
fE08Dq8PvRNSj7MrSsHpDdjD2CZ408wwZPpALlVOXghIMMjVcP5qv1U+LF37FBzoo6wnfJTRtGeX
G4X7Cs2JtN3Y5eYjbYKLloceiKlxtwtLdYGd2wUH6BtNQkkUhoX0qH8cuSZCiAZ2DiuGc+hvMPV6
r9hHaCbIAAIbRsiqk3ZiLLmHakdvOmHG437PR7doY3Qloo3JIEme3+bunCQ5Ihx5O5+1O+rPRQK1
JaIWntN5VPPbWel31JIf/4SfXG3YefHYZCVS/D5/CoguYQLmbbCJEATl+dnCYh3xy6iVecHQnWVK
8LSZCLbtlBPxIoL/mFIv9gB9yd3TggnKwDF9xotszV3Rw48HG6ly7x6DKu9Bo/b4j6Pmf5L+fybu
4aTcuwJqKsFYfdZc91psZDsPDH1p1RDF9gk2ZSfvfctZFuYEulNaIz3mgwXHi9O36PHFUpRknlQc
eOCThuQ1KEjLQzEiILKmO087X9//vJ9SC1D6eAjBHqKWiwq33/99mFnEl2NCVgS85/HglfSleEHO
8wlMcMhEcclUI4yTU+dpz+1o2caHeBKk4ugab5VxrpllhWx3UZ9O7Eg28DyVXNp6GZH0gAWvfb45
qlD2agbsEh8hHusHCxWzS3H6JtWml4qBhwJY20W+Dijdb8KQ+bDKwwA34DTiEXNR58j/ujjj9faw
DoIjvvfzUpVNm+fJbR+qDmKhCseN6X1ogNBZuMOzeuALvfAoGvKkFiTyLbt69D6KC7/oXA02ht+N
N5hapU4eLY20lySiN6g78dmad+nh0qrenAivFsC/mSWmVsAxIhyKta6l6k32PSFmIYb9Zz+xo3sm
dVSNPAeFkS1A1waO2rFDUH6Wwh3iJS3mS0qeQc3728EhYzd56WNxs3xac55vnJaxwaBix9i/0+Hm
Wv+rDywl5WYs6x3QUzhHPYM9CZMJA9RO/cDxTcZI/xJGVo4tcDaI6wK7mdZFQSvQu6FWs4VWZNJO
+dbGHjySOz2gYU+O7+3fJpMeHLfas0zzOz3hzFZdjFR6j+htk7zY5s62g5rz9jk3LvC/oOWxZcjw
kdR3u33LDZm3AzCi/zBAiff9V87bozFVpmpPFYeLC15+zEzTJWLZTSLsxUxD8OIpAtPxhaYDcGCm
Hll6rfJlV9qKFeQf4DvW4lJMyrnTdo74G2ZTIC5SWuBjexMtpHLayHbhJRWBeJ2R4Txn3lLHAT4N
iefVbBznLFFmZ59xlcYoll+apP8KcytR39+4S/+/8gCEh//B3w6tb3VBhWWBeft21a4SXFsutUOo
2de1PsuO0AywQ8kVzoHo+e1saYmYtdQ3mokyjLYDM4a/LhjxahGskj/M4BQjxqHa/C4LE1+27VYa
nUTou1KfWYbWPnRAxy+VWLOxRTdTlmqBfWESO0c51ufJ/VC5rQs3U1leeBB4bCSvSOXQuK2xHWRG
r7D1ZY4tk4pT4EIVyAUHlVZUvNSz8Qc2XeVohX6l94Sda3kCfZKPnKRlhX0DtdQ/dLHg7CFf0YRc
3YK2ukaStu9aWaT28wSIZLTxKDo6XC7hlUTbJyTBz1gQBZRJEw5M3zHlSrcqS6nJKb9LtcW4HbI/
4ign/X9toRzJq9uYU5lwnISALnGq52VudHqcHX4G2gLC/fJs+I5RqSf0G5EKRhEXgFIkBc9+uOBy
dtamW03KKGxXvnZhAnSPfUEi8bWkajx3ysEmvh+mv8BVY4dEU5KuD1lN0j801JP60OZ63WZMGVU8
Zd1f0rgykeWtWOeqWffdYJ1TfyHavI2Pw8ylzNTNbPl35emiHQ95JhxLp3N7DPlhH9VrKfwcSpy4
rmMJ1UqOLSPi21jR8yMso5zVwoQRnQjT4HD+hLiD8p9U7ZVgrQJaA80VzPH9DXL0pbFiuYQ1VM/n
na++b7+ABR4tTUXaPW4IFhoj6VETOAWcMHG00xBoBCwIybu9s/OAJeiziGJ//7dfUqRfj7VUXDlR
dYi6cPkrHhnXAfEWPRho8Dj3f3lwtOb1VwXUnLXv1YYsKR6H7VTddeheIe18bmCrZzOF7dfNB94j
M6utqzRYZ8aMv90rKUIA563s3eX9td6qWIZh+0ZYy4yi6TY/UJhLNsUBxxIM2ldIC9xIIMsvWm7e
6p2WGBUyqdJalTVDYybl4KP1k8lRSg1FhQSCusmQl3KmjA//YN1M3C2vhzcN+xCmGYSwWWCktwb4
7JVgkYV8Aoe9vqCbvByy6vIhgqFOo2MXYLhiF473vfZT+YfQ58enjjrbn5GGzVcMirAUyVNmrKvf
hqzsaPR38v/9fU3ZZHJCMz3a9ofezSwPkAEWn8TTfChYH+iieHim+YAwOHo3Y33h3mXsNZAklndn
8m5wrFqw3neQVUUhIO57N78wzluEFzCu9ta1TdXg8k0bGCEIusKoqqhBMheu32OmIoYCng35KX07
0Sl+UAdJyiXB7TkOpXkmgdWJhTl3QRDzFwFkA2DLgpUriuRj0YFiHP9h52jRg7NuI/GQu4liKHmP
1j2prw1KGXGMhA8QbBjvAZtj9Rmv402gJMLS91aUXiDwNm+UEfLQU56gG5lEC952tPmKhZTyz9wC
qtNH72Q8ZqasuXK9qDkso7NGGKM9WTh2NuJzO7ldH3s7KBC/PbwZVr2YACHENGssw3lncXr/alu5
wWgm8XkhXazDvKRIT0gzRFVj2L0NsEQCG+H+8tUHFerM26fHoTnEhizl+I891MR7NuUZCh+v3Um5
XFInm5p5Vfg2td82g3oKZywG56W/BTsKgnzg0OXDGETclTJUbZk/ixPhkZSzeuBvISNwkqnQuDU+
dFZyIUlOdcU1Dzamn3YolE0wdyrQ78JWc0XxHtuCMe6eQ46QEkO6jJbDAJ1/jzm2qAcaDSUs3CCc
vH5dNk6Eqr7z1nByGHRKDmygyBkokHBzLYOgPZQF9bYeR35nkr/fDy082vRLinlZ9tT1jV5LVQGT
uK4676EIQW/2d/mTOeQNBIJLi5LDSMjAKkps/R6LhUZGYiJsT/CZ0PBWgJPhlxyx7NjDTn8Md/6Q
1C20VWszklALBFPKTSC73EqLK5irfMuhv2avQV9j6MFsfgD9uSDK5h9b3L5uLit0C9NmIJ45MpOB
kdhrOQ+4IZzU9qEOqC2XcGpq5aAJBqEoTzlXRi2ZDkOBFy+TyZ+YVnGTTTTHju0i3MUHWO40fz0T
E1cvj5C9J0AO9R383GuVp+39uvWmVZ8WFjcUahPzCTx4BTMTd+MT8F2u+sMd5tc7LExcWe9YeQnT
Em/F17zuremU3nbn2JiC3WJrurXB80jsdcNpRSFSVMQ+Ql7irNwxMtYPwNB5fEZlzut7UVSiHNR3
X4YmXm8EGMuDCoEbqpm0UrCdDLH+//UWTI7ZvrijTfelwiJUAgNsShQE2qqCUcJh8l8hebyHpBQd
cEbfkolMSQ/Z5GzCbeKgOdsOEb3QRSSBriejCzxynFGXYd82H2iXMTKAEf4YTzU02/T2uQFbF6us
mSLT3edeaFAfW+X2Z8n4zfdSII38tQfeTGgV19lHrcMuHMduqZcFiW6T9pq9hPhCMBT9uHlsd1DM
+ss+QIAW53E35A/6fISWcaSkWvQtH6O/SoFRiDT+keJXRPQ/JxDaQQcmwianrVaP6xZD0Be9Hoy5
USZLIuOycBgZA/fcUc7G0OBa5KyikbonuZbVXJSm0gjnKFPAyzH1M61d+v5SdBpeCDvgPxkw1Cq2
cGwVGcJBT3r7jyjgyfr/hIN3bU5FSWHAtVEoY1x6CxaWKMWQ6yVYd8W9shQ0uqrj9XG/7njvTd6i
uFr7bYgRkItuDnb+bis+W65W5ugeq6AdYlIPzkkBkZ7je4FOULl5Llyv8eo4J13DeuMFBry2AP+3
NjDPQdkzsJpWpGNpBfvp5CheNtDZwMrKelcITudvciHB4GTUklL4SwWfc7CVZzUx31n9hX5x2i7Y
bnXTA5TfojwsdopzS8jV57CtKuXOeBxK7WMjEXp9HAcQVDm/rU+oDID/uGSAb2NPLmbDiphuTAsC
7jznvLP0VmaetANhVhtfGOWjypriTivpcyk6MZtgaLztt9rSNJJF4gkdaRt7IQlieS27wPxjw/aX
uyO0BQ9ORjFK4nlfznvO7Fo+6KoJb1D1zL5I/ZWaOWxIIGvdWweq+MHtb/HqIfYp0q57R69wkVrj
wlV+eFArY38Srwp7js8+YZGG7FZIYjQ0zDKqzqgeUZW4T6952j6ptmA/3+HxJeE9oV7qXKuYn9lc
BACBN5StcXYncFteYVTr+5eWN/gSTWeNkN1T5u9cuSqZt5UjsFj1Kb0y1mvReMkuxIZiqfFvtS4F
NSdd1cX641hMTcvmeCnxST24BxvKe5fQm3IbDyTUwlaCKFd5HODBb6HKKpxrwOvSol4ynbSrBWbM
I7wu/uqo2rhy23LWwK23qnscLM0qQeeESXdRpVc6B48eYC71l0OixXSH3mSqfaawOSi5QBGkvdDs
Bj1YaLsrU5n2EysVXg80m4iNmT8AinztjgIuhec22NeJ2ERNZkcwMAAyT6tDdQV1sEzaqZLG9J3+
2+OoM3aTD8L/VC41tJeJa6nhZkfGM27fyjKZckRj2+ZMZU5DslTzT8Jmcttmh8rAMhdXJAFSSSF7
TP5oSeW+GXRHVQhZItXzhOI8p4VzjY10JtIiHAenPnNFsNzlKiwKHRMNCy9F4ICGcwJ3KlTx3zm8
j0F2JbJ5hCWCSDZTIsRGz1wXeQmTzWzQl2CvD137dMUpzUOb+kIuVURqtp3HFcKBfQndHANvf8Nt
CGXaWqHXyFCjemGLsbXko9bqDTVNMqL0M706d/36CzLdLw9iU89Vube+AhnMjWUAAYHNzcdE2GE0
tB97BF/71rFa9mZM+lnv/kuFzarmMqqTztXoZUy6ZmGrb7iQqIDONtDx7Ax/HounYbYAW3t+M6fT
BdNZ3yTDaRO9Tqhae4pfEyKRAhOtI7GgzBuK4qCXRnR/mICxOF3cKkhcMtAwtwbbE2EaMP/ZMcM3
7Wx7dRwRC3Hgh0KO2HG0z+dVkU4/PA+Xc0vxMKXT9xz+wSNq3xKqxcCBGDJpxP6eWUSlKZRkQeRt
FyQ+RzGnTN+u/Or7eojMM34UUGfPMrVDobAHWzRcEYUPvVUfdBqXiEcjcLem5TupknDhg0WlkXZR
ar211HI9ilPNtcxhE9o3NdJE210zXFusm8+Xv5lIZC4vvN4x5w/AAzoCL6cnnFI+Hzr1+hjPpfRq
6PUZ00PBoNhKjV/3WnhFOaqxFet1XGhW5UpQA6pQzWAXrWni6OepzpxpdLeaaiQFh08i4oBkP5KN
V4WWslk5YKJO+Im2kcClIyfCXtliIgSP8YzFSgq7aiDq060P4no3x5na0AZTiGWEYY3MPLOtxySO
3wriw/KSYWelEYdWPDKJcSJP22GgrxAjEqbaJsljZS7sp9v9iybkecxugsgsIehSQ1d3zyRLeXmy
q4OMb8HtMBq7MNpQla1O3oS5B+Aq2FM0E1reypBLLxda03oAlBy3vRQsdu1g71UNT6LfNUQDShUS
a03JyeT7Hy8PAlraIaVkeYMiFWh3JfiZF0iAg6I82+zI4jgCbJ67+t2jt0BOoMo+nZXfSu1kZIh2
AZeMPTk9v+cguEEUAgHzQYJgu1mGl21mQJslI8QBQdHFHSFvniClowdKJ4PPTkzx6z0UkPYe+Ssz
iofGfqtysg8OxpwIEUJKzuAcedJdCpcf552UA+5rUmBFLCkgeww/QIwNWI961X+mZ7dv6aM372qa
FjAmOne72uxUfVb2BpG5KENYi/0SBwNPgb6skpfbt4sBt+l/nCdC/FGYpTt9r057dUy5SAQrMyNn
f57IXALwNLkiJ1LW/X30ptLpEBwUdbrhh+lEpv06rlmjJF8N+ZiGtOtUxsyD0F2QToVCzgrCugAA
AbX84Q+wmXEcn637YwWRPJPnqNpbtuOnKF7KpgbDW5lyG5oaY6FVA5AYuVAu/M5LbPc0K4ilRwiZ
fkfE8INOhN8xjSUgsbhFKy7xxBJYhD8ty0HRhk3Pf+06RE7u2EoRI+XAZqP6IX4O//v9mk/m34z6
aZ/7csE/kBLQ+7WyUGY3Rd0jGxbxE3k6aTdTaK5nyygjDjf2Pj4XGTyq4gOaWgibxa5YGdEpQ5mY
74tPB1vUWKG+gROnSdx8bLV9BitWp0gMCVVAevpJETF5YOihw4/P1oCME8bVLtEqKKyHQZD+lH/u
7ta+SjeOHxMupJyZJTS99v2chCmDO1BaVfXKBj20rK+AEYsuuGhBuhOw61kGxSe6HoDffEPcjIM/
/FyO0vaUuVOc4RD39EuAJl1zSvIC1ivDSiZyhW0AKG/1bR1t7H5wqyhSJjLxTN093Wp5iy5nFVjb
MwPxMTLrnSfVFQyKrBNGMr7dn7J3CQMTukQTyxogkmOWMGVod/36xxuW51d8aW6sgSm5kkyQpeoT
n6RG3fp/z0TpkyhhznJhSvMlWtYCOqkemt1B3fmXJFDa2IgLyJXHtOp2PdetPam+6AFHaiAr2/Fn
npCe8pHTNhY2CqYWXQitRMx99jhjJSjrEsnAHvsYjcdxE1y/M/I1e3cxenkmDpzq4IQGUvftokYc
VC3R/X1JkKI7Y/A4d0PHqla1LXSb6wmQxAT93T/DbtoT/78wmlm/L0sroX3Yu8U+n+V6ZNSSzSlT
CI8FUFVY7QijRnflvAtTMtW55ND2o5/KhGlaszWGU0thVFTtwvC+WX0V/69d0r0hOwSBofta7fb7
FG4ufoo3hpmYA52cescDubKE075ADjPmgZwRke7hzC+ClrmzIksw8BQ6p+jrm3QDIV7+pSzs1nX3
PKJPpDDWQ4B3Yb7eUedQYdvLk0ICVgn3qdkAVohlwh8e6OMT72eSpwl9OTQU17+HNyKtdKztTPMK
0pgv4+4no2rqT3zFdljJt828xv6YwURtUG8E/MsK/gf4I47t1+QxQ2Q6ISdAKhAYWwPsN0Tsipax
6PgddySeMee/wmmx3flccj03HAIpGE1+0lwnJFrQYW8rNq0XON0z4B56r6uxiuLF26PIuOwokU+j
/TJ+5Rvn6j/HUv0VZrcU+qGDqF9t0/JS4HHe3hUuVog0542LyqZigX7zQnqENNahOjm34ACq2HVo
x5dGXW5wm07NYP8SQBYKvaZe3T+aBoK/VsnoKHaWHRijdcQ+nqJeeZGA9KaM1gE+eqY1Lm5qryXu
+lFctVH7QatOlWVdi8lXpL76ZYEso4L9HW+WxzTsAprzUbIrLSsySDBJ5cAhnA06NgYcww7ahyTl
nQlGL+ee48pV2DEr37qly1E7w4Z1RHtubMpr/+Qhm5GR20D3MrM/7wNsIprOIXrbY1Ozil/V0WbD
AszTZApmr/gYfuOUJGkv5bFEmGAqqaDJXmwon8VJAkq8oGIEVexWeJG4KTkqcTxztDa9aozTDe8T
3BxEDtWoEW2kk1+LrOiT+AaTWTF5QFQLWduklxqg8R/JFoJ8K0TJ4ukiyEz5nEw6x7YEuOuhJwkH
nVgkFEIG3svjylBZW05ptmk8ev/wuop/0igSJzS8Govdf1sOXD6IIcIFB8R03MoYiBb+/cTedGwl
Dtdvfk1ovVd7sBvnIk72Dt/D/Liz3rBQYcxMI8b2eFMAabFfI5WAMk8wFTeuaKkqk98PfVmVJkoX
D8IwEBl6gW+1HKN3tGUhuKM/OwNsBjXwIOM1rUU/uREmpSVFIW+IkBWjs7ZC64BITtSKCmycMYPL
8hRVQg5UmHPZ6Xn7t5MDKjR9xWR5hySlpIMAvv+aYqFWqQEf18J+rKy/focU+pAP7g7y/tzXsA/f
YNvfRoYbixg95jY9xdvGXhBe6wa/tIZoYVUcVhIQePEwrbW0qLTFc0Rn3BDH14JTJpwoLCDIOX+M
mVDSwaqaOkBkewEffviyeZ/njvr9X8sBlij9L1cdoP319EQdpZdNuFdedN3NkYshfOHtRL9sYFCU
I/Rz+++O9AEu93UftHP1K2dUl0E4SQG8ejoqjF67zQInT4ZVGMnIGoi3LO3518c7dgfYTCggNmuU
v7qptBIPn+BtnSM0wqqosaKatpSsEfqxx1x7XNtgWBkVDnIe7MvGyfJ/9v5rZstqs+DorH5UPo29
dY6e0w6Bzb8s5NBPtM77qUicuVgNnRKs4AlkG+jCyTcE0P6vTnGWnZKsJW5LiqRd9QalW584z+4j
yj5f1loitb5cxErsZpGrTgc9+dMEYkUkTLy16ymmLkMHkMKAhadL4qP00VuCvNiLoWV45CGgVD3K
D9Owz6g9o7EV0e58LkwgflRHcEnj9Ow81RlHg/UTQjdecu8JWKkmiu5+ViCCzmfxwshtZBj0MYb9
gDiUYi+5aNJVggL1aDj40gCen81W/6jKQUBVC381zydEgO5gxvYtg3q9DP1srUuXLS4c9cZjwvsO
BF0h4CRtxlEmBMldi6L0we4kxVy2AgNYyMmJ06J1VY1zdac/Rovfac2a6/M2KcIT6zMgP2A0QC7q
2f+p2f6LnxU2jv3ehor6/gQDeO1V6meCjI+2tAAInGAqDuvpy0ns22p2pdvfAAG8Ye3J3oUzsUEx
VttqdwroKKk3lHw8CcepP7tUrxAmws0xUuSZ2w1Ue7IdBiGl43SuJuiqJjuRYt6+vOpRDV1uTvGo
FXiik4EUw+TXwCmPbpdQE9fWV2cqW/Fv3Q3RPs8AOh5bNBbtep108wkFq8AIIAIk+eugtYEXE1YR
7xgdVttLJbHHPZ13oArz8z8+JmlL9KOmcIoA2OgBm2r0Pk31387/S0KfDfTJL8uLcYxMPNJeNRX+
8JXvVmqhX7HQasPhZ3NjTBuIcsmxVeW+3zWciJmrYt9WqTcZ1dlGr5wGTYKQoLEgvGZCCC4zvK7W
h2As9E+79fieuDMEA/LOmP7c4o7se9reVJb4C94LVldu4xUhzF/7wp5lnRwyK7SThdfT3NXJWMAl
1S26dpzjSUheGWDdMmf6pcuiTI4ZPGz5/siI9nR2vkqDCZDD+//JsN96bOmp4I4jfQgMQWh7arKG
oThhDWqhpBYTeZSaUEm7QQ7X675YgF+jKITnhgBN2Ln1nEPBRnElYHHs7H7d6AaS4TQvrTCM+dRW
LrI/O/df0y312zeGbuVj/LojA06f8IRaPdfPHqOp6lrqJevfai/4zofwmUQnDGHGLSqJLEkymiFG
ua+CpftJL1Fiv480cU0gQ1u0bJ1EtDNWe6Pl0flv8kLl7CIPawPK+WBmAEfPtcdgI7XJXkEfCHNi
2r/kkQxhb316XHN109xh4T+MW0o1qPx1HiOlPxsgJLm09Ck2mJSiLXU7KAD+u/LsT4WmhfDx1n4U
54itSwv7EwbTBOnAxR/JOfZ7r/U0EqFu7Oc81T0Tj95AfxTkHQD1R3CxaTee/3z/yRHcXBObWcnV
A2xKp6aIw4NUba+/ZJgE0DsD2syDy8cQqKlyRJ/aKdh0TuuAT/42E6+viAzrHp12409bLcBIk9am
C/wWvmTG+uYBgpZGX3wJ+Ry74gN3HQoHyvRG13V6phSZAF34UtpteZUv48o/0/Q1u9218i6jJoRC
DeXVzUlZ6/HUyMXBH8Z1QdRCd9oltxp0TC9qH9ZAxGSkeWfL1XWaaZyJU+KK2byKnmRboUEtveaN
X7+UqvUymCwZ9WhUUDuTtXk08MI6qHsRoaBjbkEk6dINu7VfDjdUTpJ6yTNzpckZhfVUW9QbSJQi
MWY0MLprAjb36cIIiWxq52MWYMnMVY7KnVMo++oIo+Im9ETWgWyLflIX9DndVgXf6S/k3CVCX4kt
nlO006E7skdlnYTLZV0xWjrmyGFkC9IljDfIkIASwlNx5kA6G27aBp4X4p0w5tZgoPJaOo8ULD6y
ombS55M4Peyw2Y/GhIx7BLfx8B4FS2PAK3I4oAGtz+4VDV+n1aNLoE66TGbeI6Amo7yKV4XFWbmj
3qogEuLW2NhZouciJiqWW2HPhOMSKnPvWTPr0s+VnbgByT7EhpaaJJaxiXIvWIF15kNTlcaO9fD+
MHzQ7hhuHPR0/3TcmSBbQTNbbo+rjzWfqI8ir5f4FlSNwYnKuAJcE8RsRWHVVhdYWvfbvh+XZlga
as2dNbX33IA9qmaQAHc5e3G5EAM+ut8+xKhAzVsasfbECBTnNUx7UKyZJg0MVXGz23ijvopfQ4DG
+oLDFIu1BDI2i0Xr3oya9M641aeJ4vXPB5W7PhZia9uw2kQBslkOzU/f9aDNq8Va7lqPmubB5YrQ
Vj12nEkggGeeCsX7AflPFAPJiHA8F/bwXN8Rl5OQCbBQRfS/fqYIqQby+Qce8VSjUVCu3aoWUtTL
MyJtPqkXTxwTDj+NKz92j29JcqX7fciTMvu4YdoV0Wgjtfh1qk8I/KNtaQRCSUwn5WolUmomjhFf
ahFi0x+o6Nc5gFBfiJoXfg4GMhZLobCLI8hXOYx9Tydz3V60AbN1812d96j5Ti92RDp2pIqxwqY7
R0nzzsj56cBqzHZT8Aff4t/cxcmMIv8qjTz69oVv6m7U8UIXo5v0pvhx0aA4XcjWVUrrHfHKREKQ
vIMwCY/ZQaqSfmb90Q3nuUcvvIk7L6a7mPKzkVtnTnL1gNb+x9IkMT43WDJlkStGxzdPBBxnUOfM
422MMnvAlQxhJDwHtcqts9HlHJtuFhuoq2caCuex3PwheHLGVT8eEws+8Q5k9t+XNtysK+CDnchc
3CmDqt3UYU9T/t2BHduGQbikd5Rm2aXiBIwc7b4JFzNSxVwTAr+8yEvvZDBGYyzaSqFAUw2c0KDd
9NSozWXnjEbpaIwET3D97BKYx8gR6M9naV0Zlwd9+BDu/pSC4BrY5WTzHrjNUybvBlP6Ma0KtYou
oABZJ4Jl58njxe/68N3iU+ujBRqan4C4fBPdKn2z5ZJeCv8M546SDTNODlk8UAqQDOkocQppzIUV
hIoKX1xYtLCft2KCgIFCvDZJvScvGn4UDijIA6qa5Ff9hDMtf3LPwsS5DunUUNeAzhYqU2dnflCh
FEALrgnFVS+HbeR1LtXXy25RITZ5olqzA02i8MDxWycb5hO0aeMLaTTgjnMgVs02qzgWk9NI6Een
sTC83QvkAPMGPkModwPVbsAIAK7laXYZFef8oEkEGR2pjIlrYwVVk514M5O8+5hymiJSh76INe7z
9NuhRFLoffx2uWDzK8OMmarH4ho5DtRS9Dod5Jl0SLNPATWzXfHeuNzr3c1LdjON8ismJziOpxtm
NNgn15r9tV+RwsvrVI6xnGUZxfg2Fkl83kZqA+CqV1OnM6qKUUNhRRapIdg7JqiqQIO3fquLASEg
0idxgZJW2nfFSLFt6jO+2dp+R/EBnntwyrBtWhSJpKqR4DVcXAwheL6bRbPINHU1dhHkZYwPBRHL
/SXS6nS4kfEv0q5r7LNOK6GGfTNGW4kR9KE3PaPBQ9Fr4s/cr3xn4ODE/98xYzhlAWRdvoEdicaN
E5I3qh6eVnm/hb64Zs7FtuWEcCRbjH68Cc0k5FQySlTflfrHVBBvqgNuXtO3/JTrmtZJhnCEPnS9
luBVcX8+F6rEgtXuH+NEmk/O0jivMGLUCXKHlw1rA3QemD6NsuBBAIKSEHSMA1586k3u3x4N5apL
RdKapXAbTuDdy+5uyAuQweGyj8a4+3XrdGv8b2Wkx3cXOwe+mMwLBsZgTWwIETPLw+rcmRjTwypo
cYrU0lOftXG0nypBZk8yh4NgDkfmhBA7fYMJdohdWon5M/WDJe7vaglwWvPKuOZGpytmrdHPtmKp
1AHNLBZCmm3G95udl0pEqRGsOWZ3oDgFLgnySGVVZezdgMAJZMMmyjuci3e4BJYj4wcGxwahZ1U8
DF5G5Mx1/abL5+sL8zApTRJabcOQuqCB5/PgL3WY/I1kR2FsCNSWEfYGuuwwnVrYm6Oj1wJRgOqa
RpsH3MBVx6uwbdG6tFGdZr5aQCmRAyeSEFB0F9zDV9eREnU0djMPEkK//ZLW2aEq6/F5QBn08X84
+GOgSMv7GbnLjMVYGDsxo4in3GzSy7fHngqBzxJiRukF37/yu2zux9E6HzMnYiU8Sd23yBbb1E0E
U+Efgjx98ZpEXe85XpRtdebuiZ4mtBG87qzzPD24YjwrplvTXuSLr4TtWC46tiK391FZOfyrC6gK
Y7XkGPvRzaLu3UfemcqY44SHqgbi6j+bzWBVSad5fZzoX4Y/LgM7vk9F8XPBYc86ZzWDMmu0bHgK
99iippeFZ+VHGufj6DrkD+VBpC4IjadRJvY4zbOXPIHdzcRA/tlYua72j37JddVR3MFtl+iMYsHZ
BgHVB1yqo1AGIGUDCCilzsZ9vB/TaCA8O8KKYXQzF2Ol8fkKyDFQ4FN9nfSrqeK93W3hoEWveZqB
to142aVwygRBtT4ZwNtbhaVr8HaeTX0X35fyWLm7nyMLBBm/tNEM0B0d/te9+29UGonfJqaLvUws
IphGqmbXrzUuW4wVlLyyjKgOhqFjjslO3DE6ak5sfX4CyLd3w4HG5KG9WJFZTf2I5wFWQ0Hmz/ei
Mtuwt1GWqNqiPuC+CmQR/urWseNVCAH8+q33kTVoTkVHHtNwvTqKhnhmTn0xJiFGmvDq98/y5S7v
lwdrDC1yMvkDaqpXSauYEDl+5XGIz4ITbIC6cLDcHoclNtc2NNBebjyaMqMRGWtWTyy0DfJT5dbV
eJU7JpxXLf0Jt9Nr4xwKazHLj/ktgPjE+NrSory4T6/wwJto12XmEmS7UPKsaVpPRFhisT8Nk1VZ
A0QOYiC8rMB3GnZdWx4UX0UHtyzDKYJF5RncGY5n5C0imcDYzMYGIt2pS0M5h5gD+A6Ac3nQyfa8
o/tcmtk3D0RSFVZjkk0203FjCldQoQNkC3cW0n2jCR+RXwGmi5m9w7cVEqzcffE753Z0+fxliPOM
J5UauU5d3s0tYOvxGbu8OzMbGMFE36mKHoFt9bATxFLmYbf7O+CCCNJGIZbSBd2zu8C8PzZAnaqv
DkoRXFACk5r9TUzdH0TnBr3ah56oOfolxrAqmEpjE3eWRIyQu+NKFxKOZ2Trx8EydQrwHDYfO+F5
K1DUtZc1QdNZhGtOtVoDNPk72WIyw2eY/0m1nFgteunf1fxHV6zdc3y8t4zVOkV6BKuopvtcmUBq
MZbKs2J9x7I0iEMqBGKOJrdAJmQFewa6wffYxuAWBlRrGbadSgW83ZI3b5yfvdiLC2KP7XMI6Zio
1nEcyhOjKs/iohOfa9bCpGtYVftmKFOWV2mHhROQhEs1X2phDMpIieVobhhXpAoLOtfcf6tblCQq
wVPQS4wvKiZDiROStgRg9aqreJ64tx9lCmf84lhfWT5xP38nZ8W8+uFEqK65K4eFCCx1SG/ZBL3f
A4Lwxo5FJMHIvYhsAWzMrcO17K6pw64iQhcv3UneSZMt70zDdo/JKNX1kAZ8lx+CSF+x7jzIwQwN
XSrYi7jhVQTSVCBy0ei4YRvDptvVq4a6t2R58HaErRhL24fihn+j0ZBbbJwFdmqRYfG00GKnm9XZ
kbbKqFO0niYdZMjqrMuf/9Ma1V2MdSL3Fbzw53fOzATQ4M5TqFDXknpD62qfYP2yVVdJQZ8iGEJS
YTf5mcO/NSv7TKJeiR+cI5L6Q/pXI7wiWKIfri2bVAgWMh9HyqcYzPdu82ZUxlUJRdoXIbNtEqd7
MGmj6ESxQZ96+/3YP7hpabtgzIw+wdUUCPF6ELbjJopVgwkStBjvm18kk1frTCd7yid0QNnnXnDt
zibHu87ceB8xt/B9S5GcUAXDqaO4042R8mHL3J9lOO49xCaMeCrY+7tz/3vZrfBBlme1fcxXTCCI
VAiBBoc8naTWr7cK7yOZ2GSvqg0ufXHX0zglOHYhHVpoGThhs1EMXkU9EWUdYF75WeKWG17+mAUt
eiI3gQAMCGgdrN5O51eNcltmoJUV1cmu1ogzv8iF4CgWDcFnosUKihf1WrhayVfNGyj0pWPtoiGN
iQJZFptZpV3Jpjmo5kWNJcYqnG2OAO1zk34j9y9i2zVdvQ3rNjE09B/96u44LS9xNnf5aYl/vGCB
HZfUFcE/66BbUUN+q349Sq+hZhYj7iDTV4cOu/08BvzuQz7vHzS2WEUC2I3A6Eoonqr/WNXUWHqF
vTckGaNvh0folfz6+sTjNM5cPHDEWvLaPb8pCzUcUOFuJfwXWtkegEdlFG4QfArCG4LisATZ0U1L
XtA64F7ANdRaqTrrxfu6Ov41i+8+e05gBNehPvs7XYN4Ma2J7qVsIlTRzujA0dX0KQ5RELa9n0cW
OAStmXaFKOogcdWQ72uBNgGKFF1uiR3ADUukHR8hJvJ/Q8OOx4tSjQfz7xbsxeRKLGfV+4/hV3e/
RitjjCaCwOqeIvk285CRSJdRxlTI0gRwQ+ICGfdKLNhupKpflruXQMt4pLdkVD0HfDsnpzngOYgi
d/KcH2xamZXyQKp8lnziTYgdtkfa3O8IUGgOJfqqErF/jbEjBoBepjAxBkuyQsUYdkwjiCY+1nTf
FJGt5zP3aZaLlwGnyfvnypxYfdDedzYPrsqY1vTK1hyFkYJWyZ/SCRGivto2siFP9pZdSYyZC0Qi
yyr4v9u7HQ44wEjSRgaMf6RRBuMrdONLp7mRPjLk9qGgR+U5le34VoA8AmiSTjBuEEBIvrsMj7fR
8n5qw83oNP8g34XoRZoPGpZxDafym13H0S8qq/3bGfpB6GZL9VZRqdKBhRO1MW1rY2C0GzerOce5
yF4JQXY6Ptg2gC0kBREr71g5W83qS9F8qcOYSbt86xlcHoQVHX+xyvamxkcZm21EU7sXiS454lzH
ZpluwgvWlswP8h5ixgO8Pxghq5vVgMfB7MUGTA+dfLSjraWX67xNptdyPMOxQ/l6k91ubQDYWL6M
aobWUGDmBdfAZRTkdgfAfJuRLwTt+2SLEpWrzwjGUCpSY2u9nWTlPEjXvfUxIiH/hAjuiizNfFMK
o4sGFNF20CMRPZOw4cAa7GRggox61aRlVu6jxvnbmhmClT2rNpt5ddGV8BZPHisf68weWIP8Oki9
Vie0hkV5KUE7b5VlcYsXCBWJHkILePQ172MaNOMRW08NThk//tnFK9HeNOhXtv37TwB09ZxzELxM
GP8mDL0zjmo0+1+utyWSgaV8qjaNajqMbqWdZ2E/nGa62k3uMJrYDbO/JXZ2ucxaF+gQ4P2/dL+e
B361BkCNdENWL+1hrFRTEj80/1C2C+Y3WmUuwcwxT1AkuunoZpHtN5FIIrO+JyVOOgLqDypznr/8
rheEftVq7qF21NEqQ+AnwkQ94QIZgqeXBvSI+L7Jl98Oajt9xozshl36UzBOg+88WdeAjX7G6kYJ
5dkpsaWkGHHhDT8/t/GvvHlnQK1m1Pffh9cIYO6cHf+pB4LxoLKhi17WnpzrRXY8sKY9GUIfsAA+
jKgWOxtYSVDgCLc8HkWFNKrlaxNS86reZO0iNFusHZ39jUq7I0z6W9TY59A3rLir1zZ26lDUGGRs
yE7DCzd4KP5ABJaYloq7YLlmx6oRjlsAX+lnmNpTm/DFQ0qIHdevuZ4PGJyszxsnN8Haa6vLuY++
sdQbgezLQKaqbLKN00EEEc1ZLsrHbgy5CqMaMh8TwmUXS1ZUoHz+nphFhFh9EGB5TiTas2BQuw9F
N/YoOLuoK5mcpGgH0P/zReAWRzBQLeSt68l5zLkWlZQFhO2uSs8B4+jfgi5n0X87IwyygZ1f639q
6h/3KW+fRSLMjf1qCeTdh9BA5MLmrsd6tSGdYYFqm4XGMUFESoy0ohjbBzDto1vI7nS+A43iaxTX
DwL90kP64q7XBHmoadvRb6rdfq1WgjgZEN3CnQJvhjO2xkKOnxhcm3aCImJlOn2tIji7h37ppY2Q
rS68Bd3ChTKW9IYr2qSy4/dMvnVLr93ncENdixSDxhEXAAWvraQjMLaQy8dx+sNrSuT6NIaI8eN0
EXJtjeo0A01ARke6Bi2Rwu8ri5JLWdZNH5e0UDfc+fiytGHjCH5lJAo/3tnnkcQMcWXsVJKQRrwd
g4/y08isV/JpArDWZa31tZEhRfeGJ+JG/MOj/Tt0EQEjTjaJPfQk/wXMvnOEJpq9ogISZosh8ElS
A9FHaS79v4veY7SPKEQ1pkTWRupPVFZpq3mkBK0VMHDZBLG3nwM7szNAXpNQQPxxV3MC+54o4M0y
bBYiR7JUn7rANrmNSbtvyWxxGGcZ1Arwqj8UUPZhSoFGNER9HKEVaWajcr0q/lFlnjl5FhUt/Ytq
73crQE9AWeSyz+idNFNUv7xzudQgrheRiw10R6mPxN2a3aUB7pBKv/+PCjqyVaSCokJPLtLaF2by
bYjKUJ2G4+xHIvlrE6SyROPvtLs+ky1ugPz/d/hs1Z4BRxQ21nWZfehyZEQG0Z5U9QUPH5hAq37K
lfo6PUaL2yWERtFCYZ4ixmtIC2cK4kYxI0oQmDGkgp/tD0fyIHUXilzLac+DrTxPbfGJeynh97IR
AIhWxxa/HyKKvrlPHd0vnp00YdlNMPbp32DcEs2ZdKWICBH4U2iohvEKRt8fOLvQZRBF1DC14ATd
WZSfVWlQlDlrQQ8Qdvdwu/vhCSZe3MduI7+EDvx2lDBGAe6iSUgSnabUS62MRNHw1sO0mwIRDdDb
2XY/vv/UhhPXyctrHlp0weBHhihBiOp0jlW7u/JnTlxlowIjxQUuGm0Tn6nhsAzbkiI7GUTYcl41
HAwDUPus30pFnoGVdwSJaQQ+nfkQIxxca1hNhmkV5Rtx927vt4eMzbQHlkKhRy3DVAxBr4KxtJqX
0d9keU3WOQqu74wYjiLFY3lCTrb1++FuXGH/64rgA+GPnK8yH7o6Saq0JGaH1nBAG2pneCr70Wxu
ZpHMdIXFY96I2BCuDb461jtEbbVpYFUIaw4ksX9oZ+iaSdKBL+vqgctZq23tJJj3KVdjxBoblYKj
Rg1nJpKTfHQOBED9qfTgq+oRYY6KV7LmsO7nIbo97HLx5VQEHufOFONJYcSz+9BpgdCFxWlz8e3X
Deq5B8OUe66gIsmVrLxig37mhukZ6+Ef55+qewGpUINpdq5CXmVu5a4t30905hOjcEl5UDERBkbe
Xz01vy5Iwem9eafATzHdoUdv0d52uQPUQsMpAlt3AJT2IcChS6Dd3mVuKDhp8RaMofEx4vN9CsD9
WbG4YZSVJQN/3UhdDbCSCH0o+5gZDFvZ4ssUVzFmnaU6jhvg1nlAg+MU9uu4wWyYi+yuY+Gp9QQA
PfDNXmy9LXUWTh44F9E1eVhsVKvl1+f8/ubuKByG7o3g6YSVXNWnt9RBvnMSsM1xhXS+Xjb68VNT
VniZozPM/A13ZjSYLp8JJBPl8yP9oEfh67ezvOpNFxXNRyKieSY6nTIJrhbmTXBXGxd282WFTMnm
8ib1/jlf/tPP3fxp3GQ6u6lqRAh8yXTwTAwrI2/8aqjAexUGIejefxRG9Qq+XM+nNYQAvxjwTxfl
FdlHVeZBg7NzDUhuCDs3ZZrsQXVjPh03TIprC38z85dPov37p6D7fjuQY3lYmVnYJrI/7j37q7AK
kzPFPCrxvZKo2K2hXbsrjVRdf7IU99wowZ1+vY2A852WUtVF89andBGXwM3MFr20syIYkcDQbA/r
Sz6CbIq96flqEqPsnF1Irna+IF2+bvG4bFUYD7mxzHmBPSh6bvk6OnDKkUwstQx+hbrwQBUKCG3t
FCJfp3DYnEykfIlZQQ+OS72IDLnoHTxKibXcscajpS1lO5+14f2Q6QA6ikixBUu7t6TRFV3D91ky
t52YJcY0xqG9VcW5tbwVf/sNQFf+mgRyl3ZDJbKpG3JhmGbZFJLMov0e6AdjyrtyRfMW+GMfjSF5
1ngQfV6VmGXcdRyOsiEithj7v0O8RNXRLnMbfpQPMocezChs+vXXSUHZNNLQFUHKaf31TPp+XZOD
k5CCm//7LSygL14djhFgmDBADTWEV5VrPwF76WXZhs66HwdkwdzVJ255z+r8R56nnoOV+5a5K44y
fF5LBVFZ2BallbyFQIFvXpQbcjuzZMYDipspml2m+MnAk0OrvVZNIDFqj6WA9SlUx1c5PEc0qVtg
bnXsa3eHPBuyiIDCGgl/w8pBB+D90Ysf3y01eY3Z8CCUnCYRXKG0WtzFwOJBk38CVe/Fb8pzdg9k
8f0EBINqoLeB7MPRwTgmKs8/nKQxJpTIj8TXUvmueQOqbb1RtSyK6Gob2StNqxW0rhB7Oy4Sakn2
jNZRIGw7TOL4Nkro/fEFXN7+aGuqqyNVJsEALqm6BsToUNEQBETB+b5kUYWvFrOYSATvcG7kvKQK
RJifGuNE0Xu1mRzYiy+nwvrnq243vMbGjvN8ujpTRuH5hywvXbSCsORkj4+iYZcYj0m2eUJAW55B
Le7II1nKj/PbF1qoyiyJJzlhQ1VlkYSgmhz7M6is4sY5h2ZYL97Xy99N8gmCQyD7Hr/YlAjsgKsw
b0MO6p5xmv8WeKd/1XPH8e6I0U2NdKAzOsO/CVYuenSe2E5J2GNFoIUVeRX8AUNZ/xBOu19gdajK
LrpnqWhGwgQSvEaDWsDnMne/kihZW/pEm3wEIqSAwGEXDN7s4xWM9f9tBiBxFrALRUmP2jqsV6r6
UGkOoHPWQhBS2hqe0lsGiKeYcKWe5sHNjZ8TgQoBYnR7LtVT3fTqJREyvSDfhLPVy2Si97qaMVEN
ex1I8qJkWLRROt3LT6dl7akapZI6lQ/KP73KZBY6J1lRNSatugZJhux9ONy8qkx4aopBM/ghRCri
H6/jJJ6mM/Hi4t4Ewol5f/BotWlYQkJEre42c289JNvdOKsnafG2rPYIES5hlsrfoG2NpIPgqlZk
EQGxewRooMFs9mgTodUtDkcS+oqKzF3I5UB1SeiJpLASSA/H/CdLSTkB14YT8Xxn+EKmWmqq8fAU
c+LEtX5gudiFyqCBzdeNwy/n+yjGEB+En1adUBJeeDjDtI2fynSDfflDa+qweAROoNVdjW5Q3VUD
Nim4gDwL/HNkgVpLj37g2v50VE9Rgu3zSriBQxVZt5+gxxEjM5CFlWB2uHEqp1RCKXPgLGoTwZPS
RidiybA0U/GNNeh/Pzhm45RDqv8QXh7rzw9/9m12fqdSL955UwG0ul8/1TURKV33RQlykfGfNjT7
6L4oBzLyW1X9HpFmuQc2kYQ4YurEs3HxV2Z3x2xhlJiUS8Vzqi/Ge9cTOFsNfrZdAo6R+Lj0QNO+
S5t9XeLi5xdpfFBfVyRti/LoPH6AKyNetxFLw0SijuKtUX8WzboR7Vyw5ZJ+iO27ldTe5q+iKf0q
yIjfdnyi1N6QZHXDiNLKlgsNy31cA+BdNR2uXjrx7Gd7S7Xb/28Qeo6oGwHyWDlUrGyol/2BJ7AN
hLpEruBAxlRfuvbAEw1VY15DOoBGPGVihSVWZuG8tTXGr+tIF7Fzb7HErR9IcYrwu117e9DY/8Sv
54vilJwjvGNh+SA7Vl4wD0X5CynhlSPVasXWOup1pEF6QkCtwoRvcrBMRLyoWAb/dMX3luR3K/CR
EJBIQMz2MZWXotnjPkmZRBREf2r9p5Dp4DiGzk0hBP1aLD7ZJz0YjXX+FuyYg1KRkWBndx/xUIrf
Ln3tRXm1uc9a1vb8dG+bX9lvaNiSAQ9Y7c4Fj9VN8NI4DEtIc2OTU8pgApDkw/T4ox9HXqAx49cw
DLqM4xf0DjVmXf7WQudN1E3F3wdC/nO/7v9YTSQxiewIjUp1MzTirV2rZy4LC9YMa6a+gq5TBqPO
EFFdb3qLScdSlVIGHTuLE9QN5Xwb0wKZtTSH/h5hUzOUFxxRK1kQfHZSZn+nYrOgehFQhmHSRrxt
jsYQ0xh1PrsospvP4umAjCyW2pD+0zBxxPwjbpiWjEAyKJYcNygpBlrhucPVd4nbtI9EmO9PfIyi
t7BjP0PZr2HFKos6J6YpxP6GnHyme3+n9npXunJ6cpO9DCddWIxP+/WKpvqMSMibWFBxSE2K33C/
GU59QTbD4hqQbhF9FNehn+JAy/QWYO+DtY+EjtyPVRjBcorfXxDiOsqD8ZA75QwJzLwc/sDnoxLF
vmhoIXXQFs3fd1x0rO211m0t0vKPixQ9OzIFEynUDyVvyt5Qj9aBnQg2Wm4UTNGAaQ5srtVXysLW
Yb0eZTSE1IrhZ2vMWNgkIH6yKI3XQ0+yZBaT8qZIFURSgPEJ+Cm9PFUfiedKLdCCVOUmEQaBDeZ3
Px0j/nfuhkpMfkLkWXqKJI75pZTbTk2xN9+5jK/jvGfB7fQMgHpB6Ns+rqVr9C6kQXDiesIGtnWa
gAP8GH38LA7cEd+BCMZcmZcFgR6NNXtJS6jwzmmQdX7mxQug7NNT/dYFRZNDoaAGDlmXpfXQqi0K
fcFQ4YV9CL3vPE5QTq2/QxyKzkpdMbhPEtrU8qJRy4QxlrCL5HJz8Er6RixC2zkN0UqV+0hVE1da
5xdXfpoH5bykYGefm1KTFgOpErmsox/JiU+MargybUIkxfNFKcJOkjxJEFcrjBzed07+XiFhIj86
ChpJ5CvdZQfQlpb6U1a/aW91waVPWRf/GRyJTGmHEwgr2TsQn/kX8djLGw8d+PDAL0hX4y1/sIUS
Os9ottTAa9QdZozZKOHPqj3Xl+yMzYvHa7adCqCQ94d7s6yfBp1+k//1fg4PYoLUx8+d/MdWlIvu
T87tBNVBoJ5aljffRAq1qh44JGT2KVZPMnD+OrYbgX/NhTeSfvUKxzsnBv6ydeYps7qr79uRsnbM
+iA9PuEUl7Ti3pUk+L6zJrqqyHASB/FLh68DrZnqVKcSZ3RoQOWShMCT9VInCyYuGFXTAKQc0YuN
VKe0KB6xaVG6YOxDe7QvqKWZF8W8l5KjL8X633jhjAH6yuiAfgFfXAP9VmkuBuBXtuJygd41wqpw
hZeNUxEdWUPW9nbEst4E4SQV3/4qPm5TKOIa8KgsP9xtw51UuKTIkxxGfouSJs5lZslW9urvz3Vu
GtPFTFNuk9daIT0m99atCd/bwFMZUMYPkzOudUwGjwU6nsc5fproWKl7ddPzJipTtF0w+BDLOOjU
qCaWTybIK8OpDclacHZXE+acQqVb4EN0WB+C0UapG9EO9msoJLvLjB4C4DI5U0YMulrmfYGYGj5k
POkGHnFW6BjI1y+2FZOuIybYopeJ5DyuuSKzmYntkSXdMMf9SbIdTq3qbnmKIAsWj4/Sg3RJXZmq
jhFJLF/k2iXARsc5Cz6QQSP23x5EFATKk6hul9m8HtzNhWGTf1YdPRqqb6JhSn3Feyds+JUCyg+z
leEY4KDvGp6CCZV9QrCkY4ryaPOONqBcmMkyBkSBC0LQNdjF1zOvgXx36e/ZK0nYyEbTaB6LGhFA
Ea2pX4cTEwXRaNOLEESgUUqqAo/8knmPrPbbBA+jUxVfENezBzZELo6EaCyxZoFqcopKzoRzo62c
2IQkx9PYFJ8RfwAN5TQspoSoa9x1b5Lp8PIjEZBFA92FugSv5/4VuraSUHSm+FmIhsFJ1uBqUogQ
KAyMSEXSqrXCi5QAFif4HXtVytvVG58iUPX81bAQ3gkiJYtXsM0E0cwuGtTwT+PabWjSbCUdr9P9
JzFweikRxkCOXBn+32FXeTN++lSL17U/Cj0dHZKW+0ae0+THRNfk1qDIeorzitEDxSsp1iLw9znu
RFJCc5X36pw619h3VTh3teIizoiY/JDFpcXaCcUymfXpqR2iFJXb5BrefbuDzF62CSSlNv7Z4goJ
RT38nEV8TkqlHYHTElGjacUouUkxJNEltTgJgZz5TpGwPAXD5OXxMiMLeRjBxL4ZnuQKyVm6oIvl
jxmOlOaB+Z3sr/lAo776XZ4GKmR0TGTiNI+rxbfgMGgIhwVPwdT3J+9l8p6XTotqkElY7m4B+NIX
c1wo1SGRD3pZCHuODxjBy9dDG2eSPFt+ms/5WVcLsOOxmMxjAqznWM5YB8PviAJV4QSs1cqnfVqG
NoTlc8CBWHfPiNykMBavRtUztXMPJ23XynTOOh+BoJ9t9fDGiSv+LfasYFMrSxg2Bj4k6k/blsiK
dM5vHRuv0C3VAH90hsD5US1fl0K2YQGjDaUQMjbJckUpftIyHMRXZ/QIO4i6YbOdiw+xCDDJlOol
Tlj60J6+uv4CjmKckkL9ZV0lMNB4LB/XiEBz6Iv7xSd042+lU8TsjjANVG109qavJc4Mk0bQ5gAE
u/JJwN2NOhQckXLu2qE8otrwZdOovPRNuB8+atbNCyvO+vdlAC/nGO+cyHh0aCAIwh/dZVubiUKl
z5I91pDyQ7GXJV51Jr6Nubh7BQvNt3TrIuJ57TevgvF1ne+XTNe7b8TB8rhAIHTIU+n+56PJekqC
D6R1b+RtwTPfv5i19omNjyI65kX2N+jSr4zKP45gxb5erfEub5eiHLUvVKy0AbWiZWcpsuNTQ0IG
EM1HYiYl5O74IrmvVayQgzLVIUJiFflsrucBYXOZRtNdxirszsv4z9E6We8OTDng9RJVrWl62m4c
aU2LuxBv4gM09dzSfbNzO+aKypPY+M/kvYEArbS9kZZjvV/o7OFtel+54ATN7KeS+fE5/JDtApXd
xOLLQbidJ6ks5+opf5x4xOm+vV/bBvu3VIJziYJa7YFQpDge8gQhz6/LJV0bib4Vzn+OV5tIwRsA
uFrpYbsj8H9cIkW5pkt1htdctZ+D5PY1X464qmsfII8qyWpDHNhBOBkR7l/yN7PJ08YBq56qvs6W
lGEf3iSRiJQcigwQe+HDyFPftdQFEVhmPC29BzHcOw8ALbw9t1CCMbWNuAIppL8Ls5+tPhEAEGhq
9nROefpk7WKwd2bPGHK4SiOeoaMvdZkYJRKhFPSOr+RQ2IvvZPkCnGCVGSz+tloTxJ7d8dLs8ZsI
BUE0qfL1Bvh+SjlbrxMsrpfQG//Qp7KVTanL6jR9yi2IdhPyAvRqzc/BFWuKPvdebbP4neGE1gTX
Sat6sKHPoSR6FMwVaryxOXH6ClpeIPvB51YkNEpLK/GBS7etRLit5gM/w8AXgD+la2+430oumHIN
H68dFcBBJr/HCNcFJT1/KilI+HSJSXcwDg9UrFKZ8pOmuApduyQM0df4PFTZTg55HsH/4IwIPb3U
debWb17br+YgL9GH0u72acKfj/BiHDKCmEkfN5uWv76ERgw1P8EKh1TfUq1YkLasI1fSTZXoQ3QC
py/lYWFfHEn4FqjGX4GH6mKzbZ8njiQ9Jm/WUt3F/33tfPj697GG6sfATSYAAL7F6NvrxAN8u1TZ
hXfjHN6S+iZRxU1nmtjd20XZY52r5D1JRwvvcQylc/cbuknPjR3+QZ2L9vOLnhhd5XD3nNGc5gnY
emMo7YLYdf+sp34rECGB381Q6tiBbQIn6IqFL6Oo2iv1jgv1fc3lblQ5KcSOXsem1SgNKG+SGy6g
sK+WaHVOsamkKLg9dSFlKMRZ5UL5bYR+F4StLBsWe2fXTuVYJfDf7SN4onhe2bjRNCoOdcUdPCZc
UTsctVZgb3GFjCEsj2n1/NSwFSKk2pdCfTck0cau0l5eaH/H3rg6KU5dSejsd8hYmmE62ZVOD0nI
FEUtc9ZD12E3iUhY955hcS0F/e9dZf8Qv/4BAdpouSKGNghQhtIcuIBkVbtq12iTAv9Et7icgsWj
GYg02ndKnRdyMQ6yA40M2Gl75pS71FSzAPreqBqtz1rZ4F+YwUrKL2AkoL/YtfUzbI5yQPRXBTgY
Vz33wVCi3df4ImueCK3nR9vjzqhqYU+Q0XH7eQ8dqeoqp4VUxXOHQbAfu308DQxkMGI0Sclhqwvo
nRfsPvZTC/PhPAi+A0zoz0Zg2+wry6GGWcMb9tuY1i9eIj1vkIPZUGLhgUKCFNmUJ3YY/SFtGYBK
Ogt2iwK48GQXlZ38UaK5z2zIucmfvGv6smyU6TDsin9T8/MuDksi8INL7UW9z/pIdg8koBJMXC4m
bCHwpdrlrf0hkxEIfxwDsrB6fFJkyG5pDEqpUcKgVOiSBMVCub3IIuSgxtZD/fixgazk0GrtPbgN
EWjuOQ9cWG6F7ym+/LHAuhDMfoX44TxZb7V2MDO0+/P/CPRiid5pVcaLRyCq8cnttXIvd4WW/iJN
B/yDMhihuSZzWUEOyRuf10XZo6IizVhc4IdOlPYx1XOofLBy7NJHEmQdyGQYT/Y7hTPhGYVOVjxp
blSxj5ocX6s5WsJ1adSH4Kxy2i2SMdZb+w+jwmHGjE4tM8c+vrEhiEo4saJWKPWWGBTNKg7fSGpv
1k9Y8Rcqr6B/yxWlcVwfepNkLKbqIE29L1e3MzpYxrigxrgySQPfbMACRBUlV/2ql7C2xP1xW4wC
0lo3mGFVOiIBrttIthwa6Kk9V6dXEHyw8xL0/8IHX55aaieoDDSFWmo/d7n4qCUkS4UqyxeScjlS
fu0rmYlBvNwId2f1i+yRrANwusgEF4iValh/vjHSnu2HeIdZlUupQ6oY9MHmrKosKyBn8lYrphbK
EsBrQ9En/mXiG0nwCZc80yKiDHz2tAXfs1PiasBGOTw8ix2HyRKLZSjAvq992bOAWz/T1tutkEDW
vuf/1IOPY+NkYNMR1s/VyeXrTIJiJ2X7hQkQ9hlNqK3+4GxuPODC/ZwHxsJdMNRMxjdbJ2o8Nvda
/uyEMZ3kxBISKTQcqPmgwf6dEyNL4gdeCGg4Yqj1CM8qmgeGigx39kW4SSvk4ZpZ+KMSloFMCTzP
7X+qX2OG1F8+w7moECGHWcnq2PcqPsdoKRke2p+AX956Soo9V5EfYXo9jf1coNbFHga7yf5Q58rh
PRHHfLKok7K5pTN5V9cR9hDBNHG7tCodS4Lki6q1lOW9mN/Ilb9PIrhCnbnXMe2Az9+YfHjiMC/o
8j9wzhNY2IHp3E9gpHD7p2tr70zfcA+a/ePUWtrXlEj1zT3gUhxRAHdOd44qsUG95jbiLXhCa98I
jk0YH0pKyWwO7z7vRJeEda18HAWrVeTEvZ2JOC39kWVec1S8wRQ+khB1TbiwYFJ8KUYR6awam3pr
Dgh7imB0IjhKKQrwX38N0HKJxPuijdsD+xhX0e7gPqNZUVMXkmjTY/UQwac1eE6nHB2RdBWzggn4
hS9oF24odsnGEOh1uOb6b4SOY6659f5Oiiuiky9cu5zmHq9uM9JIB51B4k8Qu4v3jMkqbkuYoMft
CMr+LuTzRcSAxFNVHwjyhJJoK6UbfIhaeAr4qvLPiTdWDjej/xNtPBT5s8XcZGdiYoPQT3Ify4wr
BZgKXGKPtgfXSlBlLUgmwYqIHklR1rKUQblryk50f+ZNbbF1EV3+Nj7obJX/yjl/N4YhWW++VBfW
zHKUqEqkgRiQEqET3H+EddzJQJ9LYPqQI6NsZLTul7V2ya7iPPDq1lVb2zDb0+fNeeEcEw9Z0S8X
4EWLkS79bZyRKIodpniQ4UlqZJJ0Se5bmoGyLKYqjwCWKfipP56Ipn3YN0Supim/mXt+26g6LhRn
5q1iBavZqtKAX7RjBrKmsUrcXKnbRDTzmwigTcF78TjLeh+buuKedKdNe8v4VyKKWhzALSG6SvJS
cWcMlbqco6ZhVhtk0kPWzY5+mPT8Azr97RAuUI61twwJIdAR4AFHTp66CrY0lTBB4I6nUhedwinB
HJdSxZ1AW9l14YsJZYoVQgBgdBiLIHrHZz8UqzlBSAKeOFixyo23ZhuCTQf9TV+vKLT6mMvxj3RF
kM/FQ992XTOUWBnUxL+EygcDlucpqlaPFzB2ivJnIDQMZy3SQXgvvl55KMEylf7rAdxC/eOmQPuu
dSNWzrfXE0kfXi7/yBY08sEEPN6M6T0nbBQqjZP8jWWEnc//oZS8X3gAAxZWA5+p0zMX2KNkg86v
PIyUPJszpXWwacrpcOApZwq3vfO4VeLtgwiTPzWjAyq8pNOfNl7Mw/3ldr4nmPuzAQ8QA+gMQCMW
aTYndbaCx6SEOs+8uoLvPMAA1+LEgUywnbSewVUgeU/6b1x7i5L99PnCED6qk0Om8i1OCnhQ3Nm5
U6Q/MgLLlZcuB1oxmjdn8QnNzoIWFe/8iUVpCaoj9DWvLWoYUZlEwgyF2YgIbfpyRQkr51nZgj8/
EXDJAjH7jAXOkFco7GseCQnCgXmilfEvHapGixCZsBMRfErEdBRzOwF1ZDmStczHaqSMKKB8JCuO
LHuXSmpUg3tVJ1smkQ93Fwcx8aOSI0zjM3q8OolE5BCWHcNpwNxp+t8DkgmO0UaBIcCvb+N9nhyQ
uZm7aTcQrmrGoTHymOtsO2m3MER3+vf+XoxksZnsCu0XqyVBex8uFpEyCBh5S+RYmlJjlsme86dD
vnVm1zYlqenkGOrHGqTCRxGyJ1/KVpOfyVNOf/cN2y+KLUCFEwbtl6Vt9nNpmR8UBAr+ASoi6oMH
pL1N8OBgBE3+J3SgrenwKAnu9JtrEbW427+Q8Fjyn2dp8HmP9zLefODszHqpfGBpjl+Z1xJPYJNX
1XOm8m44qNfsne8Jd1SvUCv9/ASTqgLLnSEq+0lHhbT55s5YtVbQ4jW/HxYgpiQ8oTA0utt+9kTx
BUGZRqvWTRmHh5BxuiHwPnximDUiztM0FTduuTh0A7xRzbmhHqniiaxGmM4GOfL2xE3WFWVdzywr
WVCCNZ+9u1gzi19Xj9rmluXiwtxIDCJLPJOu9knQJu5bY2UR2ak1b7t3XC4K01miOm+28N677ZKc
zZRBxWGCpAkkRe2VsXFoDAmyLEdgwE1hV/mRd9JG2BLRxj3EUAywRciM+RrxLLWx828z0dinjux7
0P7TCPRCtk91BZDmfI1JoIR3xv5+/s3rpT7sBwpiBLqDtH5BzwkyYSvFxCDpoJ2hpRpRErM2kKIT
F0CqlcEwRG93u29hSZkF9nco25xdAMLno6gV2FMJRo1e1s0a1M4dC1hfXOMsSiNdrPoDI8OlQFqb
x0wqnQbKACRc53UNSAm+ap8UIVDdAVn2S+y3mKJgqPeukrEoiCyEc8qtQ+2znZK7NyiiXkKbI1rc
cIDTMI/ziugl+CexZA4oIhaSPPGr90x4m081ltsX9vrg/l02C8jG/v8HkQ2YKwpnLH/6gxCF9u+Q
cdzGDw+Eic1GYhKpt2Jlnc4UJAdlygs8Xh7LASCtFXx++5btioeiEEOavv4RmU0EnKJU3YaaxLJP
2qyy495uOpQEJxXRtE/Bihf9xzjJFSxNjuPtuMhXE2stCqyBedFwHz2g2kD9ff6ZhAXdZH7sRph5
CxFnMfd6b3dpah6QGXhTsLHu7uFko+PfBFYwe+iLj61AmU2Q+IrHq8X+r6HvSly1CEHVAY5dOdij
oz1Ouw1YnRpkDgLKlFccz0eqtcrm4JxLqh2jIGfI8L0pSNphZiMGMoHPvyFVdLoMK3qN0YF5yLRq
OqwGv+eXiS2sovB2u8YzffExOvZOGKMD6YbvS8sdfcTTxvUQvr+9nMokIWkfr23XXCsLJPiySX7j
aL6Fv+JpP1pUmBi1PdwoqWhyH92zjtGP/tctPKLxxoRRCCorzN9h/xYcvBwz9G0fe/LXfOeB9Ank
x9EERq8ZyshNU1wFaFBOMh/hegIx6UE42WT4KhKpZaXmhlX8PJf9jO7z6rehZFSt2Pd+Mgg/joNj
F/qvGINa4SIzh/PrHIGKUhJxnTS4SG22YhcOGbsCSmkqb/DFKL4d0yhkw7gSRXFj58Ms/7vaoseB
4VDCp8/ozoQI8C/ZVL80AG1IVpUqsj2TYd5g9Z71ANhGJtDymYqXi7s+V2GfkyMBCkqod3XPXqoN
zpFyRx51KiN3HKjb1eSyVy1ZKSCAzRm1VY6i7qfwopUU3oSzc9TWD2Vp/CJCQoVK/L83tuYd2gy+
fMRDuPzoggUTGzAIIl5H4VXUvDTJeEdh4g1cL/qV28Qs7tgOdpnb9EysWQodTZwIwLCYVfAaKw5A
OPADa0r+bYtMMPZfeDmsFnP53dT+la5nSZhc8NIS6WPkGW8/KV2+J+QJhCWHXxj5rlHKwpMKeNwp
6m+My5htPswj/CkBrhtNDDnECk5vKhjWC8OCX9kO90Cokup192BtdQdAuL7jmZTDVs5kTG90NiRV
STxVt5cDyXmU9ky6iKa+RP2RYCOz2TCdDIxZa2yhTA/uqNDaaaKEghZ3wJ5GHn+uoFvDAgiowqP7
Br2mu3ltpKnWnodg2iPh0GA1yDRK+YQG7MuQ3L631UMsNwVcTE9LfK0zCmq9g8V1mMNPc9V54ZKW
wpWbYZFDhDWW0QJFgu0SvlcG1Exv6m54XjBcyIAJ46xJ1y9TD3Bx1k/xeA1Fn8mCRxWLbMNphiCM
amyIYRV8TBwMRLMI3Hk4enS/zv7iRWKWR3sAZDwRSRZuWxl4ABTrVVQSQbm+SC98WpxoCY37oeJG
Q7Ne7d+/WYEP3tT+3Y7P7qy6eJaaLSBXN5tsNDUkSGKqGkMAn7gglbr8kNeSm61ucWG75tsZ2I9x
OcRiAWoSnZAWn5elXofopdjCOBS1yZWjH6rTDvvNQb5JlqN/q6V3S/DbAFgycFWEfkkdIpIOnetX
O+x8HubH4HfGnVirpPYPi9JnNln5fHnqa4FEfODKz/K2wTCX9RvWEHGEbzDyUUHruEbdePYNG3Te
Fr925Vk1fvByv6iZZyPhrrXFJR5skSPNHpN9Bz6L2R1u08a7iFyfdSt0zvWZSeJvz5ER/R1WFq92
cdFU2SgT2pPjt0GRFEEIXB0Rh1+3siuoG9oL8DSnfs1pYOvA8DRk7gDcVPZqDNm1cNHNLDvchv7a
gKhFOeMsi60mMJdr3QN3JcFVc7H0vTgDUPYqD+XJeVpSTDuXbk6hCqHBL35kCaqmweq60FoGbaOL
mVLHQMbdevs/X4iaS0oFiCZxT7dKrELGtnI5JjPVOKejjfYPPJz2Zk2ct7NUHmKMhb4ycbMCODtV
o9h3Idb+QUe1G8+FRVIgt65k26EkrPnEo/Pep0NQ5yKWA4WDxM3Z8JrPKIH7XM+XrtbLz0CKXT9i
ff6LsvRnfMtPy/+c6Pno9xcRwzM36YeCTRVmFHs8HCPxPQKLP9Xw7ibx/QqGPvntjBcKlUXgglcW
mQtkGTPrp8LmNY+BG8gJoSw/ak26vzsCxxNtILJcysBirNTAE3e58UCgMHnu2mkkmsnt2goAI22s
ALIxHKRC2Ntn2eX+1GqEHTl3bD12q8c4RbFDCJouZRJD6Up19hHwLwWPQ9I052KWeKexosu6U4pU
13Pkxwfp2zPslFy6PrzRYrc3CF/Slb0VAN4qqErzAdGKZjWDtZs94xhH0lcrg6Hfb1XlnZGTbmMk
Gvg+Gjxt7blgSq70ekTAfl0VKnCHXgSuoYptBIivzCI5qVhrAl5sAaEsH5DGYr+vvtInBc4bGKhA
iLOtefp/bdxENsEJjnPTvl6mKxbrniPXTQJ28GdV320PCEEyXUzaAfXwYJsMJ8Xi83F6sPFLK+mr
cQ4/a6DXfBQr4Xxf3BFvBgmMPSchkMHFNJzAAUBezv4F8KXbHjv8AYVmgdkFBF3ZgiZL4ylLraZL
SwV6gZHW9wAojrYql16316z55ZQ049SylhsVeVMzeTbxvzP1QWYUHPkwYt8K16CM+MtcoKIkP6O3
vM2vwfqOu0R8pPx5+6va9K5VakeJ8jZx6MeiuHT9mV7kqyQAO451uUJtyXmVXI2jYGK5XLa0Z5/A
BvzOhBm7EsnpSsbsANX7nKT8HVBBwmmQwIWc/6W6uWzSZOfbGSh14AU7wWH7UPPZ6r1qGDU599hr
shOQDQcw4xxOf2K6rq254fkXaPcA5WgZobs5OtEGqgqlz5rceWprBwccTCLdAQJIKl94FnqKikwn
jAkqjDY4ZO6a7fKbqSGO6XioFl+TdYJhyhcnGYDK3gNfimEuG6MM73sRcbFMK6VXgNqOtZ2sE9oo
uvPsJK/+3NCehV/CT5WsD7YioVRrguSSXqf62QFB0xxcSu19PEnD2fbQkMhDC6f3H8hdrKOxoSj3
73xVv/55PKYH2llp05zoR5/S0I8MzJQxq2FvjkUfwxxddKOxE1I32GOqtgC1PcQ5DBtD5tjipBC1
KJGF8zVOTYP671HyzJ6h3VbrPGKjdTus3HyC5QhNGDBNOk1LDA9UiBb4lUk4LPuJnNkSvAJGpKQL
3bvgRrCIZODIYD0h+LcsnuWL9R16LaxOBsgqtjzszEzVJWMZrsuTrQMwBiMf2tdK89g3eH5K6QJO
wsUG6YoYTgv7bwjdvd+K8Eq6nplzU5vKKme+BPloDI/17TxRvXJW4NQBZdLlNl4lMXc4ZMD/D0tm
4n2qd9A0Dmx0sM0Q/lLfsDX8cY+h73+0mMLuCV7i/6zOR9HgQpJJIRcFzoJnRYHhNBSdQ/zQJSsW
3Fs3Nw2yplmBFRvJqsBu6SvchAMTJ0jVhjBQdWoD7Q49KHElR4Ar5urSSW9DvKvhPReW+va27JTL
RQD0H4MuLBBJ8PkUwFo5HkLRdKGHa/suzqm1ECsUI6QOIcj1NurAKcmzpiFV+kEqTasfcgnnXCfi
JBMUimzslWAgstGLQYvLKYPCW7ywew2lf8+8MNpLvkAI6X7sX8syWMjfJWKs1rYeDd1mrlsVFTLt
uuRu2zH47f///c5RsZBXfreQv5NxztP5/CgDjUq+NZPpbOliFWrXvjojFG56YAbjSIMchib6pYpg
+B/I5aRN5AaWpNlSIkg+edGl0zxXIVdxSbBjWDIjxEe8qN8sz9SphcXorTHNqVjSkbyEixK5FfBL
nEOpOaM20HSe34zv7bJmyWyC9d6lHdpVKoeQ6XP0+LwAAXRSy8mtRDJBPmoR9IrNM+PeZr6pasUS
eKgKSapkk+RwYaWykxJElmpbcoUDnjRFgh3hHR2xvBuIeN52elh1NyLALsY4kBc6WgAly7RXIMJ7
qd9NpB7ynqEQn59WsZRDet+h2Z5wlkRVRWkheFrRUOR2VZkFjJOMrEHqgKjTIS6uBpYZsoxBDhKY
VOlNnICGESRLsGfdYKqGS5km0lp73+Vm0amM6sw5f77X4RklHkl6cz6UB0KNtj1uQaZigpdpBELG
L+spGatpgkqR/gtCbD0vPT8X4+g+xkZqMNwW/AGjzUwVeRTacbdIQ2gV+TawfJ3hmeQlh9yABBN1
tSfZ2cpcljXA22HK1StS/6VirOAbIUdsK3u/okCUHrakrgc9Nv8PXVqHU8VOKLxK4mgJRGijSFOE
1W2k/SkiKiZYTgeB6T6f21r/OR3z9wsiaIqjn9oCpUAJRQx4u92vq/rxXbzPJ/DQYKyZ6GMEbML6
gbZ8aO8PzgGMkEiwzzrGOKLnWPWr03SDtoap+fDEDLRbhKKrxfaLXDxecDTJ7qClPETb7i7ifICk
19i+v1JOLoLqEyzA2273K4x/QgBjJNrJiW4YbhwIFErXV9V2MMGRZATQ0EHow57zH6tZE1TJqhg/
hh2gcSogDYG25rPJOsjwqzy08Yqk+Vq75nhGfWc77/PCuIGQIFg0G5uuDs/Wokrd3NebHF8I6XlI
JIo6OGx1To01ejHzCSzfEWP16Fm8on5fWhDAyCbIBjjYpVKoa9ZUdQdkHAkWw3dOubFPenygHPT7
FUDoQKKXB7MRxJJPAmurKiR7B/EqES1x1C3gJ6fCgCbtawvr5AAvnURuWsUdafz3pcmd6hzBGhyH
KtQhYXaj19yNk3fTFnH15HgjvQ8/iNKQ3gbJ1BjWc4eKt5cs0lDyuik0+IHu6i0OjXBU4ihD0P7C
jaH5gDLwG/EloVgYYby4OtOrLpCCqiAKTXpyUNIri507lXDmoC3spaES4gHsadb1uLBuC1DNLsmQ
uMCenktnuSV1zr4JRSpjGkTcoFgZwOc01RpTRB0iyHUrcsnKQGgoM9+w42yoV8cvZL+4h7+A8ena
q1fOU4wFJx9iI6xNrTJ+FNG6yG1cuYjDKW0hLZUeRolt+rd6sbXdOrOkfskm8I+2JWbY/lJXt8tH
Gfrm/9KIvaApXpKSQ3U25zog+XgzqDOWUcWI9CD7vfLUvqWiinKKhMS2lhK08f5a+xWLZseoWRzb
gOiHXiGdWKFtJ5/oKR11J7bFCLkgDt5Bo7S3xE6d/Bx+WygQaqCAZ7Mswxj09NXvvLiUVJAgBy38
XC3SlApW70ZSM4bPEe1uLzqlaZNHx63iflb0doIiOejf3ohYTdt6iBgmEBm3AMmcieOcNz6AbqXH
9+vEtlWNJWlBY4liEcsanfKJ4VLTmqPI0aGcrIzqx2ZGUr/JItaxOGaiEMv94TbZa6IvnF7I7NG0
RHDU82UAJroG52I3mkazohhzJBkmvTLyhp5pat+eGMuEK0qGFXf4+dklAS0kMxS1y4ugjeVZAiGr
me3mG+BHYeMsU4RA1V2pLN1W3uh9wwbejidgjapUY1PWYI4XquT/M/mvku6KRH5Scbq8sXmBrHXw
+l/jNule0Ubecfey7B8F+c1/rHiceN8LYFoLkRLgUzNtuu4eKoJ2XW85N+fonHe/anlqY8QJ8uTh
hizvHP1CNkCbEYV7Y5JcApSNfsM3YKYfeC3bElMza7YcVxqSUZ14EQcqjY2yTJZbwJtqKneYEGyL
7C8JjFog4yQsU6+nlWXubl0P7FCU3X3Dz/NNikcZeCwoHFFPifzvX8nXSLcRT6IhC5Ua4HQsDnK4
WjFOWyq2HqkPKsPlooRNiHmyC3uMwA+fd3CAZ5gpormp+WWDh+pbL5NVBWOvADlBJxmNvcYQ7qWE
1ODSXpxRnoT1OcoeqlWE441SKh+swVAahI1rHziQsYwVNH8hJNlZ9H/l10o2x/TeqTJBRlQ6RFqg
4Um19LJarKMlhFGp35jTETWvp9xN6ffrEkI0teL4wktmALEqCtbh0G9yUAm/myBkuDWj9SoGg0GX
IJ9BQezjD/xntT5m7JPBbYpHwHao+RkIZQLEU/AgYwy83+uXLW9ote47RZj3BqDWOS3EGTN3cEtQ
TwvP7rdtScG84PnQkvKvmmVAaRxNRN8j91fKlUfWEnaftHqldTODQ4FIkzy/rvoGofweAzv3IL5Q
1QqbZWPQIC9HCJYaENldEKXBJETIsVfEYGhs5+a/7OtqUqUqz9zSElIqfxuVdg0QP0sXlNc+oJEy
DisZV8giXtAyywoueda75D4thSiAQeEaSCuSAnTkS7Kx2/ZU6MITxRDbwYZ6TLtISuHkKd/EB1Ck
D5EtSToMaBEBktMPRWcOKpYVzDAa8Bf4V+Ecy4PZ8nJSoBjOLcc7ss9yprCd2Tig5LD+KJOjsyHi
lLc1N4VpOq7CsUToGQXYD5b8/f0eJxTWyrT3hdO/28og19q1AWfk9PD0sK0/AW8DDkLO8qdDi4GO
JYMWAFmkYfcfjmf+n9O8OtIJKgXg/ZVcbizIHLIl6fBKL/w9gtUBa/rnYKeVxJKOVbU7Te5qcT5C
DFtyxl9dUgNnR7V4tmby9MRYb62QOca+/6jqEawqjT3s+Idf+hkc+jX30oCCZS9LwIgC+6xnouMr
p+JPPgmG2C12gVONnxo+BlMYCYTtBUJ00Ym28TKcK8L5IpieVfaQiy2KDdizNrwgvqLge1Ar1G+Y
d29Whsx1IDVHlieF9NJRLLG6T2jqXtsiXio7x0qffSkgw8aoUCMpfafbVhBSnbmY3t8t0XybHrPJ
vK9f0QRfdC2GFP2kSLzvb618SIdNPmZwtacmvY6qJxxRmlexOO0L2TEke+YkI+xMmJ7Vu8EGYgHg
QjzDOevbqaLXKz9Tuf0ms9XOiJdHED6Xl3vcb71foUKTPrnnwDI/7147tFXgw7EEnXKLNDz2EM9m
jBUhrzOZGfN/iDAki5rhzMX3h67XsBKxnHg9nm2ANmB7ChTk3G9KPX7lYAgan37RKh8X6I49WoBb
CQIv4hUqrDXRRQrTUJMCo0iy8OH+xflvk7b9CGuroewinDAoePyNvMogPM2CwWrpRShBkt1r3UWc
DvAMWJs3VWlwM1/AjWzgbBwoJSDjlIkqqfxQW6V591NMRUI2ZTsQ4zhQR0kxIbRcqZkMHhgCXIwQ
zmtivvEHA+8wZQHdk041iz6zJb9nAooIXPsDrkQxivOyoa8Taj2lMSfu9Yhh11lfzTGytsh/UQ30
0+SRpk+mJDYuIFdf7klgOxeYO27NPcTtGQlqZsxqbchOlRQ7p6M3PElpkUd4OlbuRkM8AbVykm/J
sKq0LM9YjSvOkBJQAOHN6gDCvt86bW5dD6XfaL92LgUPjvxTjUltrAy5sjFHiJ24PLIV7yyxwETa
WHDrf7jpDA/+ThGh+KScttLrV8k/nMlPH0gORsTWz2dRiKdu6e7NR7tWGWXCANx9jV8gvSqwqmYN
W5fGpXvFBwk1B5Tk4K7VjIgXwvj0OUT/ofy6PV8GJbThLiHb5OAosPi2Lal2yDwzOpAMN+uCpU1v
azeMkMvbS9UAUvqBiHmmmRlHt7ZoY10EqGcxY70oKRFqjEJd+YdEoSiivFnE3eaT0nXxplAyx9mB
S01DGes/fTMCILguzIq9zhycfTPRK99b7zjt8DUc26huE2fprVtE4EUE0pHzpA+bOJ1m1FsBvhS1
oFB9LWJtqubP1iBsL8ZpC9u7beTqoR+DsG1mbSrOu6a+xYT+y50ffXlEEqoGaaiHwV7/0HxdRZek
QTVZE3mC11+SQrYpgSs7kamMLdLYskvObvNw+as5S0TBdvFqqePe5lav/Noozbq5D4jq6Ap5e+7d
FVKNx4Eh1kGMpe1UvCyIFCdepzKMEONx/4J8BBnx4yKGX+2s34FJtFJYbsWzNzRUMkaqs9/F8fDB
q5EKbwposLYpWY2fjkDNvDhjFCBgULrP1J9Gd7SUdlurB7JqDXAj7Nwx77XOthm3oN4GpMuUBpBq
s+U8+s/YjxqRDjTXcBCQZb07iW2pxpwU9aKpwUQEyUn+kMyy8NO1KMtcEtSAt/sTRTav481Ihp+P
k3gHZxgSJh9HxRoogqUS1rkPHjEg+ti0S3Mv+HuzepT/rVpeBMLDgUZCejjQtsRTtgw6NR/pTsic
5DB5emp9GYXKvGhDPK9q2GRzoma4dnA20ZnrTDXWEQ01ZMhtCPld8nG52VcZvBQ2B0KEniHok1Ty
zz3Sxf87oAMdjdog5A+uPtip3mlJZtIQar3rf7fGg48YiH0mM+XlROJR60PCtkeamZAnMiXv3ZXD
LJknl+u+73BYB/1M5rh+icIl7cTp1HaOssRTap32AohsaGtMD9b4r7CDMZw4xfXydy48xfQfe9iO
fDMQJvbOaEBacWaBbRY4ZvR3A/dQQSxNAiq3/vCbKYP05EF0DpHpM8CeJ6xzXrorPuzxZgth/H/L
WRRjwRZN7Ozn7/YUv0+J1x6kJWIBmCnGB+eQC+s1wfNXwIQyPuig/AsU8N2BL7df4IFniXfWkIMS
f7gys83tCcDC/7ZpdeVnC0s98u/EJw4yjzKDjXJ7+stUGrW796/D2YUkCABnBxcrvSENr15UdyCr
gF5Trx5PRg/quot8Av5gQ5vFL9ff1M86fEqN5BuJOY3aASQnxNE0cNVp9W2tF4yyZnLvQASHlzZp
pgsk/wnWn24nBxmbE8aYhC0BwV7oDWuwUszrCm0L7XE7jMFqWDxGHZH3pmb1RLQj5LvplaNQZHPG
HoQqX2SvnH3Q9nHEBw1YK6BgLP+7sKuMoW1Q8PXhF4bGVkdWKOuLbeWH8qmnb5WPPy5cxEUEz7RL
IaQ+xh6xMQhtFBiPxFkhv7KmLqwJPlSFJN4yWaOl3HZHgOI9uAGMSJL4ahTey3TadMw/IP92/72u
wYr1Q8JVPSyCgoSvcpG9KKm/Lc8J70l8P4Wu3iDfNGlkShlwzvpfDM5wevuwU4NJw9LAB13FO1js
pYBZMv6LJcESbkZ72IywdPtKsxIDNBcGj21V2p6dR4N42SpiqzTODsKkxINLzxVnZHEigP4uI7zx
mRq4KLcbODk5sL3nOvdLLFxObnLVfa/J/1X/EgjoA3nxKMoHAgfwsnQvti3N5gzn6Nq8JDuHu7VB
OC2j7YrjUam1AUCE4U3ZUKZr1oqJgLH0k3oYTVNGK+nTw+1FHpNsqg+7Vp2pv8B+tcb9aim8CStF
ODOKYCfuzNKSVWtlS9/JS4d2uS7vVVufOjr1mRRFK0V4Wy1Lor5gN2lnjj6FdAk5Uqn5r4fQRSgC
voLZukGh5BkoFVhdgwYzu4J55vKCCt85C7Ue9mDimCGMviy/zOod4QSXSIaTkkRPFpfwFo/2ZjDo
ThkaQsYkWDGS2GMqbPZfSLGh1jGDR+XWYX+JiYVlN4BzF6vdInuU4BH5ZxZG6lOlVpqlhfDRfm+b
9wOx6Uko12neKMFMFLUcvKwVefc3E5PLfvJxmq0Lf+myev1a/FuXeWY+QOCGIHBwWdI9z42/eLy1
ifLB77ifJJsmbfz1sBUdLBwPkD4a617cHoz9SucVMNxfSIeDnT0LwLuAQhhpEJPAnXAUx+J7TY0T
olyubY9QPH9MOkN4ioRJ7/ZDnyMAg85Dbov7z2CLKN1HmOelYBuk5d7aQOKjI+7Tbqfka+9/rY4G
nHdh9B37IvrdRGx6TEVmGdif5ifdB+8TFDuYo62ptPVhR3kIwU49zEp6XM29y/ub4/pupDdT6Gjs
b2lx7R5J1Tu6CdV0aexABSN0gtMWltq1BC3xdNIf2vFS8UnHCWAamFGSerIjYV+3UxqRuKiPXryJ
v0L9yKI81gXRb8Q+J8Df762bot4dKGUanjOCZ1By4M0zWRcO3MbONikgIFmpKCUY7K50d7OOFcC5
3JYtdyhgJKClXQNUwiIl7Ti3cOGREp7M/6tTsie5ai3PacNanltAqau2tm8XaWs5UObA7nXv4eCu
MPhAuaE1GHOlsTsnrtidsz8da779R+wkf/EfglvkrW6JmuHtpXiATrN72fz4a4yOd6ZpHynum8Am
+yEoGy/Tywjwp+nJL8i0jWb4QZ83WmV946EFkdg9yuaEPMqtMcEI5duTEonJpIsvlqcLd+YdYs5U
fkgSD+4fC5aKL5x3dPxIb/OWWriFxSyKydiBxAtXLo2/dSKOTL+Be4O8dMGogmr9aMW9AJnttl+m
3++X2T0CQRTC8wQIkNBQXJU8pfOksQSCz1znul4ctuDco0739EEG0Gqv4DkyAKtNS0QWzysmSsZu
tBLffUrn1ptetBCUdV6i2KInnoCw3sTxapsxncK4zOKNMrBltz5vSyufGB9954uERrTQTOeKzzEw
nyOKTahZWaruJT2aUxAKd54B3z1BYGCss2ySNhSfIKuXUfoC/2Nt6PEZGmxY4JswLdSs2+JlwBej
rmpNJH3gi4/3xcbDpZ/omja8yZbMVakzptfH3gKLPof0wrJTPQiAOv+em41ZiuAwKCXy3rmPQ1ov
zbTPMo07a3MYKSDgso/lT1Cc1Iq5OAWe4sgB45m9qB4dYNVt/Oyp8mf5zOIiDS+MRTSTV1wtQvoz
DxqNxIz1CNm098mnUpkAvDuHxlx4/w5voUtgB4uskm17EGSOxi3z1xicflhuxEcacfOehnlIGSeA
aWO2Sxi5fZ7ICnFLaOpm9pQvNfzqkIkwFR1KjuaCp3bBWhDpkIgl3S3a03N8gtU0u8pE65hZA9pe
rXU4Qhu5fTvTHDnKtcCnC5oZ2j7vyLIDGrZM9H27qDPJiuzB/YjMqMwUb4klsOs0+e4cqL982VSh
H6Dhd4J9zCSTA87p1g/geRIpiXRoQeDHYAhI8JPLrEGqAzZUSndAzkWEVAd2Rx236GxbLUi3E9ZE
KE/5sLCGSZFPOeeyk8mmxVr+OKUDFqbSxNly7hd66XC4Bm/+qQ0x7nDSXYvlfurWq+xfoKfAYtR6
Rqs11r6boQqoAajx213kPxSIK9mgTvIk+pKo13vL0SM+A+kOD2k16w1SJjKgp+XgMPn3BAuDL0/r
vvz1tn0vaDIyjaHy9vIFnTogLm4brii0PGL2KX+5F1OuMCI4iV5s3x/WbE3bhYPhh3NMDWagyD2M
6xhDcok46f3+XVODhyvmMXJtlpnqmGNWnjulwXTCGFwDA7HJKJHxqshi1qFpfTT+TJMZMX4y8gc4
ntv96H09owyFxsMHXBn9T/DfFGxjoVkX9IqTLwjYmvB58wqPrdZvGjsbU6mW7NaTUvjk5wqWZuke
qGE6JjXXWsWBBg0DIth+h6F4WC2nmvRHdRnEdr7XGay6jW8GTZroOvgc0nj9w9xUGMAYXpPgbXlF
A/2C5+zDyCL29LZXwKZD3rp09P9pXm+GjKZWCe/+6nEWXQJovNF5iqzp7E583r8FNRbK/j1K9sW+
nQTHznHx1K32c2kTe8qXSx96MoU8x+n7VQsqhx/Zo9TEUOXdn3eHhXaDu071du26fpqATSytrVKP
Sg173Gfz4+oO2pcwU07jGPJsfyTyIyV3f+4bL5zL1V4v2xf7O5URlNxZcJkzJp4uxuxXcAlaDi4g
hl/4ufNR5TGEY3V2zbpozrQkqMMuOZ0t4YrQ8EWXc4dwqn1dDJtoHTn/rMILsUE04XtvFawgXAip
SXZfK0xpzD/nZ+aUzINQUDL8gegw/lDWJuDjo/Xgg9z0lg/MQDndQEReZ2inLdyt6NIvb6IUwV7I
ZxlEKuTlSBAe788NryNAX5EPckozU9cOfXywpKEPgIkRg/lC3WWwdC+8Zgi+z3UKtIfRMXcAitYQ
UP5DQ2wEyL00WHvjXfXfVnrz42EIJiwijZwLx5m1bZCNuA5YiEJoj/85FfWmvqy7HS1jlNXX5jqU
e9NiO3tCEHIJUqzu47yWT9tb8qFPI8XcxPFXaOESSzCKdMSKtN92veeagE3D4+nJy3+8IRztva9c
2esaxedBqs2x3k+aiSjGfbC/MeO7pLuLPeafqnJC07B+jlIT/22xbN9GOjxi2SvpcCIK1AW+VjkI
wbmTZdYk5AGfBaglobODtElxiADI0c0KZOhnQsmYJq4CXU20A8S1fsk4udL9KBmSqeU0sga4yxrF
o8D7NIkccx9eEVQzI24QbQaX2SHdXYgI1ZUfHwvXHxwJ6Bfk5/gzMbfGRMQMl12pmlOCtlzH7umI
EDHaV3K4BBy5UU0tdKIgor5x+HGzD/rPMkJGIRbDRkGyifqZe7xyk3RfaUrWfgXVMc1TWdPSTElX
6ANVQyFtmEF8mW25K2L0vAWqh1r/JRpbRxXdzQmf41Q7OMTqlidOUhfFRQBRllTZqoIO7JOtLLqm
QG9teeeT1mJuDdO1vA8Kwq5Gxs27J7xKHSvrhrhhFAHd40TSseG/rO0NkQqT12OUNBiWg0304mIO
s+EopUP8CgrWDoFYWujoWUWeIChSGv++zSs+rbjEs4YeqidevXxRlV0PGA2ZOc+sfOzsxFtK/Jss
kUTe3CzBAreSaaJqU+I8BG6qaN7WRr0NHnhZeKyd9tdQwF2Vitnu4J/nNY8shGIuhruaQzKTXi/4
H1LE3V8lT5QF9IKTQ9n+B2dvwWpNkPJIGx1FtJx3rQK8IjRAbvU5JfLgwjn6Ps9GtOh4WeWXG5t6
6KdhPLuZBGqdCP3z7aNMHq0CI9nT/7kDS8jRI009y3gHNPDdSi0CdUB0YxnY/QNjYfaXS31wr8lg
LiEvSTcF62rda001cJiXFhIgUEExK8asUawvMl6o545kKoGx/eLa/bzlGjQEag6Q/xg4EG41VMhu
p4yTWSeLBfyugLePzfFHjtDvri9cSH6PKc+RcUjh5SprXcd/gRgey3HpJyMWLTI2/94l13KtZFtU
a+UkOOaCQexHW5AIf8DNTnmk/1AOxudNGCJHWKlKdR0+HZKJio3CO1Nuhh2rIWVXsNvppmLtXX4B
AFzD2VudPS52pQ/NotExp2EiWObEfqL9/V6m1voeBhp6/1RkXcn9kxZfUB3EMOJQz8L/nNSHKpkG
TIz9YWi4RgfVU9mW1oAQF4q3s8udqwSYDxpPOIGd7kLGBN5PcXBeneR1jBvmQESUwCOsqSRJ9tSF
S2zZNHPl7RTIWai8ZXQUEE33jOkNkj1U7B/eHM75dDFzDUgi3DgqLEqqpnWqY6XrqIY9rJz7CUJa
ngWTEgV+xC8/Kl2YMuvLl6gsg7gay/l1arOwAx7CBAgaZSDJNgXcpv6sKGyDrqs2l+DMVipCu56K
QP+avnvZxMomT15LNKLI56pR9FCjlu+3Yqwbfpgm+dUozHdemAC4Givfh5Qx92T9xYAvkU7tZN/L
Tsgo39Mw7dS2Ok/LIu6Ac4Hf1ek7Z8U1Opcpm3C83E2UmzuwkQcDK6q3/cVX+vdv4IGPiKF7GT4x
oHpfqlQ0ahNGLueoPvTyjglOGelqz/OvvKqa3EgBCJ9+WKjGSNJpDn6aebT2r5axPiG0w8Jzaoqz
p1QRGV1vwTgQk/n+u/BeItwgFy2mAXRWoA1+wE+gV/pd+yXNIb8tWNKfOdRjzys9lpxaUJN1toZX
Dt7mJ4ZQHd4LIJygsI6YPbA6g5652oRCyzUaZeB1PI01ivFvXkX7YbQ7jp3MVwsISUYv2MtfyEma
N48rkaHgsHgxAZS2yoEK/Wa0z05FfPJaLg4B54D5MJ9ArUADiltM30MeZCpHlVvOyFatIkB2o6IU
hsEy/vGFuqcaNeaHs/6bxfIPelE0wftUm512/5xwvMz3K+3Dcx+4L+3127lQXrEYUUcMcIIY8uYR
pEbUBsLsMllPJRfFJfavUgVjGROfELclgBnunAoxyOjWOl3AkjfzKogg5UYEVAeCd1otZbMYC1K8
QHUdp8ieUI6flqTW4Rjf+b7R4Oak4QUsAJmRvOKMxAhN7aCPe1+yNVk1u+nrdea8/RZtb7qa4bKs
OlzIOY3rQ/Rp/ec2sm0+l+m/XPG2malI0wx+gVNESUD6hCLFJ61BlYdddJ7NnCcoO894+5gF2p7o
uUSH3iG0vhSvwU5cIFiw7ZLG0v5HyIdRwPVK+7EYFFtxQD7yooUe+sQ8AzkUtUpBUZTn2/N9HmlE
dByBMSc32HKqETKRbE0vKmXK0pParjKFrGfxq+p64Lujqsu7wAPBE6QvSJysXXjSzQhS3e2hf1Ao
QI0tndC6gULqCLl6t+1qWFIPW9iVJd1OlLjXy8XuNGOpY/AU+SxUWBaS5EhYel7Rr/vnNyxlhYta
wlcL0PkMzZI26ToKu5xBIglyZts3/l/SbzsUjVGTleIahTQjJaVJYXOt142R/XoN6ldObredY3DN
NmpKV+QBRxQleCJtHkvukunsA2bv2SnxX7H1vrDCGXQKyH9A7na1nXm8Wsnt1KKn+XSNsYwMFo+h
aL+0l+CtAsZBh4M+kvxpxh1AjXsxRu+V1Jbza/jByCy8lzFCw/QhZxxlDbWyTntl+eFK2BwW7MZZ
csrft2wVa/c7yeaiG6IePRgTkI0arIsKKEs9S3crv7Bh9qyUEAm3JrgiSPyT3kfnIw+yTQV/Y4am
adTsom/AAT+XCm3zqLsSWi9OE93k0eXkxMVW4YBPoGHr/Xy6SGU1Za9+jZhV7wtwV22I/kHCyT6K
qwbcqhzbt+Gbg/Jaowm2M9zMwvf9QSEET37o5e7XnrlUIkk4dEDyncglEzQ7CJr9MOgxjbMPMC22
tXPfplnJy5/J1hR2iwBygXJVhsKvcG0/lbEuTUk6QS+Zdi726m6GxsGtZuVB8NA7n2Jn82925BCF
SaYTmjff8Sc7yspnSFHEe+RmuQVAWWnrmZDwZeH4bDCD/e9QBg1o9t8JFxluQTgrM84pZMho5o1R
lga3omOJbYM8EKxGMhMsU/YaK9LLG0i7oMWa5D5/IoGENoaCH5UrByxeRaLQ06daBkDdpc4h0+yh
LXAwnSLpgh0ghI26OouP98STdIKmfQe0BLw6HiTBehg0ALExoIN8DR/5S2mTeZ6Vjmsgs5JhD3Ab
dMWEfEpcXRy3+jNReRwdGZzdEaHI2COsHbltouMMwhNRqANN2TQ3Hacx6/jTRIgVzbjmXlHeZvZl
lmcJfMn9lbdKARsSX3Wa0QdXZdqvscHjLujbqJgQVJ1udi9W+ZNUVw7o47DEO3U1OKf33Vf1lUfJ
yWooNfZhmHWTOe2W3crfnXHqJ2NB2d/xvG2m6sNmTgjOLb/3tV/SoQDMnvDmBipPcZYb1nPs/cOF
TptAX0A4PrqPDav3/tvPEYNNf3EW7lhLwkZST8ApMfkDARXygObN8nFA3JPjWEvA2bO0xIn8sb1T
/cZz/NcM7veptNzzYzORcYnzxHPDb0/h11inhrVhPqdjbSwmTyKCyADWcIDl7Dw2j42J8aZo0MRm
xLXBb1k5vuYxGqhAhtNyIbxBrh2V29lF2nLQg1OQM3fdjPHakFWcgzBBghutwGEiASQ0SJv56+1H
oymkakPWrhnPcZW9tgpDK5NDPLQUi69CAo8x3LX8TpSom7IB1E6J7za42g+cSznvKiITyRmlJRf0
nd75m+ablU5A5Vewyz8pDrm9z4A+jaKQHKC5C5qtCFXXVXipL1cdakSOiLKZJuvQTqXEqRAX0hBq
olm9ye18JR2+3F2WdWlE6/OfY95+WvViTVMwn8XlhZTxiEMFvOm2T/FxUU8ART3X9u/b3hiG40l8
h+oUSm+5CayQdZvWhNIUxTNRgSwO3IV/WVKsvQf96cojjvi6LeQ1yZyqXPF/VnqE1JaE2HJ61z5M
B9N92BGCcCfaRaxmrBBAtxO2YRB3IRdEeFEmmbyV+BlW4JjhplnlaVO2jnEIPuoXSp2+kbToq6J4
siKmxpXEdVc9yqS+sCP8Vxiyi5rkPqmleMN1Oj92herMxIH6O7HkXL5mzYt47SsI5j7BMEg5yI3q
bvLN76op5biCQrMKzEXWjgH8tnRcs8RcD5DgplKANydueCgt5oqN0lDQGh8Ukt9MNsMmVruxnOgI
Fyr5LmE4SVsh8scJiS9+KinCYBUEX+8ueVKWUmpibIQdSlnKZRyWMgMVmoF7BeeROft41eHzNwX5
RxSBFBXlo6zYUdtQr3MMLW9fTUsY8TGao6BaxIdqou0lIhX9U7pmnwtXeI6oEQvZSiPFOOA8mILF
Z4KmlXlAPjVDZR+Ke/OzKK1yTD8+f4i7tN8Aifg1mmWptxPME+ue1vfTlVuQoeKDMI7mQpwdM5EA
Bfrefr+YTJTIJTS/sLMC53Xb3VvcRavleZVWF+sO7XqubTwNr0xRWK79w2w2LYKrZxQ6Bu52rO8e
GkN/TJtsDjlRwFjn9f5X697Vnkddq+bSpFqYD/IJYedyYP4Tn+jvi+MmyaZOXjzRFygDL2r18GYG
nv/l+P5nB7aQmAHp+Ly9KoX8udytezfUHqp3n7QatPic205pCsnSAN4JSjAMDxxxvdUVUs2/3h+s
dPX+PHaeVacFjZs1fFEDcs6GeConu9ITCROQl2MbkUQE/6Hja9o6HbApiRC1Mr28iu1VomN04b8b
M4indazHhzZV3B0/SpJUeKgvVzs5ufGg9qOXx1E/DjgTlvhXPZ0yxDfOhhXIZuqIuGbKIwnTTNx5
VJwJto3TGbpzqpxUoGos9SGGBORubtrbPpJ9o79EXyQqSR+67WlKVo2zaoi3TmmYjJzHvCJaKlRy
WW4HyW2+JcjOmvbMBVOmk7A5+5J9eYxnkUkhdcfJu35MR9fp1oZa05ZGjIJq2a905SpB+VK9RZCB
TKRH3ieaNwDl1d5Ac/V4N9d7y2Di9y+39524V+CjRIVmmvdxvyrrpFY7275mdFpmpBaG1TPzaiqd
YlB+gHJumoZfYo2Yi5XTJJrrccBQREmJJIZpRUeAXZueTRR4A0TAbIZlgrkB+3R4GyBshqMEv+sb
1Mnh4P9vEvLtvNqBvmGqBTntKK5nzc+7Zf7IknJjFjzgd7NTuVnSIE3PlEa3lbkOXe2+9+e+dMzM
qKXM1eYFDOdACrUFXjpYnXxkskf6A/THpcf+QEkyXvFsBSaQqbo8zWKjwomOeFrNjOJbz/y2Lndb
YG/poRD8SoqSltTDYIXeGawOX8TJ/M1RTBo5NSRCBKojJN2gWVruvMi3k3e5ogbWIALjcPZo0fnn
6jSG4VeQds1fYIy9D+pXr/JslhcNWjZpEk5ZrxQgmtZCTuAibIK4qmmpqLC5ASXoamxF7PfK79LU
ui4h2um/0+nx7derWm1c5/I6TsaOF9imzedL8ATtHwH9AgD3rXH+ekQFxzCLTkHL1/cjf8qKfsPs
kHXHnFLWkklgmr41l/AbJIBZfM1tvWnc5vAJQIqSYnRWY/5kA+1A8SM4IY1ewpQaP1SBJJXQsV0J
5KvUBulVsP3wDdPVcLq7T+E6eB8Dc63aOJ1W5UdWrn3CElSjCRluFkXiGmPoGDzcylfuiRfDbiNq
zitbYxxOncZOvuzyf/KjuSI4X+wptJ8MdqqKe34jglglgLh13UEQ8m+PfWzHMuEp/xOuVdVWebiP
sB9m8OrlEpkX/qqpmRUSHUDV+nwb9Tx0LcuKS5uWnol3qf8cVbSDYPbQjfBb5l4F/w+aWfgKm22q
gmaK/jW/Wamx54zfHdBh83ysIIkOxJiWagusfInZhMT5GprvtWiupoEo64SjQJrvJOGkrRB8w2Lb
KKEgy8JMMsiY4u7TxDm88l8pHKjoYT2k9QGhP2mQWdqdHRxHZeLzJN/+SEJXcOn3qMiY170qAR+O
UkyFd+J0hm4nnNVdDky9iW4q9AF+wrNgaqX5l51QdgJzGU04YawZI9Gm+GnoMyk/V4lsosUC/e4n
v3DcitFGCWBPmpv/WkiUwv7GPPjwOmwjF1k4aEnrnoZngdXDKG8qY0GCd+w2TPeiR3de7kmEQK/k
7dgu1nWBRUE2rT7bPk+T4nZ50lBEfb89uy5grA5J4OvDttjYEZJnW9UfDXuOQ0B5S6yCFy6Ldjej
yMSl9JUFve9MGjm/Ce4B9cXUYNJ1Zb5SkXp+j2HEIOsku4QNhouiZfwHieF4fR7oCVdt5VI3UiZO
jjaSB/myYxwIkAixGgjpUkOur44qcWgYvhU3hiqL7v1ISasihKR8+clbtU/pweXJLkcM3dOFit7n
c5/mm3YXPKTuJt533ujOCbQ/ymXhRnySp0FDoxh84kcTUxz5pw/Gr3q6uvuYQnRHGd5fQWGxyK4v
P2ba7YitB21+nFd8BdQCoOP3SJPSZxOsIz9U1uTm4Cwx7J+v5FOPMAv1X6cRo763mGueFK1IfET0
4XVTahN/GBnQlB2hNwJOCc7bNDL3pjUmvqTVt07/vShRmIk6c7lTtLlQ09GczpUh+iOZSSdaJwVE
Tg0C7mJJaQQ1G3kndloBaBkOWkNwBdZPb097nJY9ceusUrSmR7idyL+3G+YokNdPBznVPkJoXEJv
GX0wdVJL1hjPbtwWmIU2pFJ7YzpvO5P1pV51Yqo/4kMtwaTTEn0jfYamKOnqbBhDrxWbVtgdV7B2
P4IZpAxBIpJh8ctu9hVUU9b8PXhjTtaBKqFBbzkVqAlttGFG+zgt1GjEQpZvaI2JKPVNcBCgvKkq
B8DuhdPTUaMKwugMEVtPh1nbv/YIM7OScRarv3rFI3VdgXoH2lOYejp0GXBvPmx/do9c24KB8mcu
Ew4p9q6BI6eCz/wd82BU96P/PEFhMLiC58CNQufabIG09lUOzMUWfn3QPMk75hdL7fSINfUflHsn
cz7Y2/YDEHZt4K51tvwIo6tAzO38CUPNFi7bp/jlHN7JkJcsV7b4kWAos37IWSN8HCByXvvQRfru
FPTDBI2qlaV73eW02xdn+SabeG9R+3jrmwAHGEcEuATK7bEKECCFPKKd6qLbMWtHO+Sj9JolfGTb
Oou5ygib0GTOusa01Jeg6y8UvH5m9Lg5hWuENt4JLoxDMPa+gcF4pAKpu9Xsd0vdB0Kb/SSfVTpJ
u3jgMYnzRNq2WDzAPydu3uzdx/nPmM9grZozvdHYGB5kwqCfYPXXV/zpvaTs1CnTrdXQjVtYfOoE
JNNOxaS2JMmOu5eKU6W1M9Aosq08VzjyI/x316M8lWMR0yjnjSt/ws4mr678/dMEKasMvYhOGdrA
4tpvNDR7TmlatVn8k4taORQ9kXEJG/SBOcBpYgg5q9Jji1vS+hwfr17mywXCpiANpi2BRTwinZPy
2rHgG2ZjVws71TJ/PeaxPY/r4jbqoawyNUjr1zdjkX/0Gbhwlf4zTecbhy90fVpj1Xx5uThfCC94
6sp1FUeV/WpfW+/sNxRiopYmCIA/ULFTXC3Df4haaMD95DJSYgqjUxLuUnBDXV/q+Q1srj+aW7eJ
59U0i+ge4q/qdXRoDrYgYZlwMGjugMlAxYwMn7mMbQLeg8wQiEwho1tGF1VzBgZqnUiD2pMtsQC6
tpQ0OpoMh0AjNto+tBlvVCvZKGqX7br6+7IqUBPj2fOB9X23qHz9zXm0NEp1LESquPpUsVEw5nGO
XYk27cVgOZpdCMeaQdkubFf9nKO3Tm/59gJpj2l8SiEfRKowniP95Ni6ZnvOPSe57pwNNoXJLEY+
vdJKn94+e9xZhL2hgA+9aM/FdNAs82ggrc8FdZpePXtR4XjqYugAbHpMi+3WnjwgFR1q2QdCiWll
/vLqg8pSR0QtKYQ3uGA3e71TO7FJI20nucL8kRrCrVCiRISJlDujQbJpB+CNYg+mJ/9ys0YuJnSp
KMTzomHf7a6Onbc4ZaALd4nTCE08cOfpkzYUvacYC3M6FsJ+aOI6E/qh4PJbLW5wZOikH1qhNVgG
Rz5I5XdODkO/jrsiV8EGqai4rKf/+IXj3ZxjlKyA4slnsUBUuyVbP1XDa72ZoyunJvnlyfRX/Gq9
pgzi5Uo0ZY/IWZPKHtTe4LQBUh6uaLXLpsus9BUK9KK+UIaenHi+WTuBvTYjK6vX2Os/eKtcyqbc
CwyXjH0HhF2vdBar//7HgZUz49etLRklm2LvBSSRRLmRogaW78TT4ko1NWEKlp2zkpMH40zvrQdE
0tNijeqFg5rTmAb5rsMkiy75YodpPFbKtI+NtADxJfaNHj5VjLJAizQjStzMvFONed+qveUnaBDk
15u/5t1vu5SZAPr6w9pyhvdhagw5KIN9C21oOjY0LRXK26MX+vjTvsoogwVEM7IQBP5mVKHRwgKm
Dex33n/S1CW4euLvkjDttMhCHWuvncO/Aux1hD7q6WdZxuw+op2bukdRWi1tx5Z9jgsTyEsALOcL
8NkJEiOQdSd99CIpqglICkcVd0nHmvYmfbOO7diW5zkC/GxQr6mG+Zy08MCLcT3w2bpiSUBMVXp6
tfdPGNYs3QOsZmg+Bs1ScZ3Vou6VHkeC+RuD9ABsSkM/H2gosTG6getFqcDx3/Uwd299GK+Hmcwv
72ZvjV7ipVwMXKU251v9USm+H6gsk6OAD1rcxYDwuYVYu41AWQ5mq55YHNTOl26I8mdDB+Lxgrwi
njItbkl7Cc5DZkISLCnlo3lC9BVOsBmkY1L2ivZvxeZLlSWTsyajsNwR0KDn7vkOpOJs38Me5UDi
qPSQA09P5I/8ZL/KlGWVCUMWRGttRLxx8W0y0l0lV+TzRGkoadsFiUOi053nA9mRUpf7QdQxSQ9a
vSZUu0eW/KQxR+1zvQJqml4P8BrJ5bCkBQqZiSnCyzJIf/v8lZO9so4KF/kxPc2Rlw8Pj5JzYMeU
5OKbPQifSk80Y9GvXZlmJNLOW+n1WPC4I+fbYbHrPMQ9u6ikVnNL4iGhKJKjGXaq1JnukUn5glFT
0gVzOixbvWbM6LK7nBoiOXd/nkGpPWk5A20rO9Jq3iYK/yLrxvyVLfp4W2UlU6nSM7tkfNDIEcM4
ujaOzIHIaLYlV0uymMJnJoM4V8DZIx9PdipDMRT/HS5G1JfuHQJpGQkuIXUzQNazHCRBUxsUblMP
oT95+cEQkUb9pNgsMshKmxicjdoP5SRkmnFo71RPs49XheNaoxVmHa6T1NfxANSCTjge4kLeWKOr
TvyRrX/OheSZ5k0Ad0s3VR9BlntVJ1tvpidRDI5qDL+EI2cjOSX8o88YldOYsATehuCRsDauw5a0
6VvfAMBX/UXuQnLxLcrb2f8pl8TkGGb/BvZM0e/eDQQiAwYXfaEuwQPZ1FApUf5a3hFdMv99TXto
0aeBCf6vnmpU+7H0cj+KGscel2iuz8X/EZ1aWZs6SpvuLfJ5g+wy1AbHvjkw9d/a96xKr+f1Pngc
mW477uDxWwMD29wyXcuEyqObOjacrN3Lx/Tt3powcjmcv8Lh399/Q3nG9jFMY0IUdKvdArbrF5Wn
i6+c4yizJHoFm0gDAdEG/oC5tOyEKKMVNIw6CFBKWTYEdKmCeNCzFRISRVQ9rX3U7td82f4C6XVb
0xrjS5hYZemCoB5lAaJd/e7h4ON2facv1vxjIyaYle4LGYXpGRHKCtSLwZQjRDKot/mFx4FAb0k0
LvXEfwBLDt2EJCu3QvJJiD+78vpRtqQbgw0OjcQxG43KTKyTgpFdYiudcQYApG2BwR+DCXgVUEKZ
6b7mo7G9gS3zWzoQIlxvo0hxpaMjJx/0tqYeuJQW2N9FHkmuaqBXvTQEJnYfJsIvv82kRJi5sHbw
ZCmRYsGoQa5JLD/o03QKmQrfmRHwlQ9uGciiiDMUH/NDxrgaKtmrpdOb/T+6erzKNEx+rA66jZzZ
WdlKfkj2Vr4g3bXKNmXuo9jW5dqDUf8XH8JiMd0t8gwF+I5SYmYVHj8KZNKQUi/XuQZZ8ZeSpIjJ
3jhkGV2TmaJ/p+LyO/UB2HJCC97JxIfk3Z7HrU61toEyMp3ofjECOaI5HK7H0vyf6L4HDomtvtM0
ojwL8A6MsdWCucCDXfj4t/0UHjPQDa4QQIQwSI3BCJ2E73T+b5aEJA+f/Lg2J8B6JNi5YkSgcK5O
TVGK6T++DxkMzGZdTOu31VgpIlpF+f81gzBCVxTVPpFIgzHdlcsqmYcwkxegngIpAMT7csrYI3f5
K61t3dJGfoIl2SXEq4V8Rx2LTPkOAX744ie/ERzGQt+rUxaoDTmqY0p7XO+MDV0vuYoze5OXAVqQ
9weHSBDAuoX+oXSkH0wM7PNJMm2AQBJ7wOWGQSr/hV00pL+xizwcmhsxOVL9QoI+bMTFQLbXvkje
j9U+zg0XlJ72tgXIGvAuvzWGQ6sKKBF8pc381P3Cg7lDkUpI0ODFu/JT5prfJCHGSud3h7Ppdegh
96eNkhZVZdLygpscZ5o+axgGhQik5UQL2ejDQKrtIZvEjQZ6ll9ckgCDL+Mmjir8TeEG4HhKz96x
3VLFfjlwCOmLkr+XgIM+jUXpSMhJhEEoTeoSoJNd/x1Vpmpjgd1I/7VOSMTjRKHIHDv9go38ghPQ
oRdiCm5SsregGrIHKvzYWDc/Sf9OdUWT3wmOK2YGEEefZPAandbVTikbhh98nEFua5xVHNMhGQWz
XIOxpJhcKowC+HGYRryayMKpAd6Fn76IJ9YoEAOkQ6ODNnIb0dPIc+ME4D+s0N2z7hD2xEjgLydP
u8TDM3oboflaZZaiki1YU00dkDMr+GH0hGHQt+6xQXj0Bgn2uFIfPCTS3NEw81vllZwi2imM8WGX
8wR/VbrKWm8OVrxm9HIh+0Lsb0RUnydUwl+pajiwmUR1c5OIGYejQnh1OM7yEkjiuxyIT6sfUHGY
tiDeDSy6TR7wEvubcVjipVT0cjPQTHdpYmeHMjtAlg+iZk8lN0k1UcZuSUO9OaW9v7bdHhCAbJ84
qE+PyYhnDudJ83/8YgEGhbWfN+rh7y6agmfmvgZtaPZ6WVykv5Y5Q/k9Kxk9bNLKQEQAJbiBhPsn
yk5OCaSGHBukxUSVYENL5KMFaGsfnTmskMWSMDD0nvVvee6feJ3MY72RT7OsAU1Q0Rpp2w1y94x5
nfDvNZcWPstGaEHySCturFjEKXrrWJ5KYVnK33K6gHMSA1PPsmSrVOAiDmhCqWBwTXBjwZ3zfE6b
IYIkn9N5fGFA01L32AS3pNRiQpYBB56YCSL1C6mH1ZGrWaUY1ytNLlZVhsF0A7P3YCQ1zM9BU9Hl
vv4975GLY4vIR6MhozWCJXOo1tDEh0JnWsh/JRcVLbbPkXpfqDw+Q5MiWAVY7ixsNeWtVoGOJcgg
gS8VtaDfiApJjdWpLKRDfBqIB8jv3kQ93T0xYunuPmmfGp6yyBYgmPc8GCXwm+36ifIBCNlsjud+
xfGkLSIMPsoXte8C+vg6EOs/82W02lQ6flxiO2RbWVZxK7/IcYbVU54QkQBAfCgpwfOrLyMecIT9
sxkJf9smQgXVeiYR5Yha0ZKyxBMranGgqHteDyLYENOpbjlYKhlJgd+m4NZhj1ppi7GotHgXs/gb
s8JFgcihsD0iAsqG1Ys5ZCxvbsg9EtSpw61OWGOhWQjmDzK3Z33HvqarStSMZyUu1wyziV6qNRwi
5SRsANtaFAd+V3hvIvKkdVZAb6k30Sh/pX+kiZrMNR9EYqf8uKZ+WoHpuAPk+4HNXmM6D39/Y/Mm
Jp7LNcAmRXkzLr7iwKcjqXdwCI5/MBjBMVIjtwAD5A7VJiX8iUMBX8FdPf8u1Cwd0LJ1cb9uut5x
e07me/+7psLqqUb9GE2kMqzolknhvEHVP+z26aWVLeANkXW7wG5ksLzt8p6WaIv0RiL3k4WpHf3S
vApUjs+Whu4ZvjJqTjNj26VCkg9/eUPwqJtEg2x4gWMW4GM+nol6COGu+7jSpMaO02nDSK34zJXX
KHlqIBVK8p4RMPntVHzullQZzyYRfUFnLLbqFYRpx/GGkfFixRZXf1kyJn3T9IJMpJ8nUIocI/Q6
6lYgAam9fqre+j8qh6qB3zVNtubNQRzy4fL0OrT+UgpDi1dKiY7HeIUtHzAYZLBZ0094fmBhsoek
D3P0L4Bg/swUFluOrueSqnQgX2xwStyYKkPpX/VSWZvONRZ/A6VNtlhDpbd++XVu2p/GZOuIkpZw
dZLIVSFWbTX/AdeeJmJYQzMvEUZjXO3vnYEbS8s103VLPb6Ad+69gZm3icRv4jyHbezPh76vZ176
WoYKT5xkZiODle3zu1q7TyDklsvzCqMn8BPz7pCgnF7v6sNm86q5LcnbFvOeN9DGEiukzL9GCfR5
/rPmbu0ioUqfzsMePaOdA3KJrAr7DqLXgjqLNaWfDLwLFt5l7iV/kdvcLy2g+K14q6mmIZ9GblUx
Hi1vTcW1x+Y7Q0xYHYLOFWChbozoQPlTJW2keNR3nvGqdamuy3q8VyR1m3Mx4OsR11tv1qvHxTFq
3bBZK9zCB0vdACryaFXzV2fT784hUjzTMoDds9W3G/pIjNM6IXhGW2l/g3/7S4gDeEQu3IUe2VPL
Ej0YbC1pRXzfNBfx3bV91jiwSyNd1vevKMOK9Pq8DM4QpRQVZ8GrnqVCtpvZirOolzg4aFy7VjZN
lqvFyLGXK/jlVQ87uDOIpezdO3UJVdh/ZJpm/OFb/vShUcKVsHX3n3g+23eqKyrbQMqUC6J2CHXl
BGx7N+AiIk8uLie/UCeK8hQrHKkJKpyHjKOnFdO1zzwDpngLhNrGiIP3ubJZUxArcLIaghPzG6Tn
z3cXhHXLUOjYWOQdkvvoOqiT0voSujmIxFyJ/FmXA9MfzdVwxsu13f0Sw3PxPNMTZc5ugsJVPNvB
rJYMQ/0yYE2uVQ+hQ5Htvf5IZzy4pRdta8IkoMxaRrReoKvHoUhxnDZQmtvbK03fupkoiAqzGl2c
/ZwgAQgQkmKKIPy7KH2j2zCssaoIJ/i8F6iz1d9q9hlX0142n2T0mj0iiRgA2homlT4b9+DPDEBG
ZJb3r99RxJR9vQraHeJzc7INBxWN8mTPAM9UhRPsHTdzjjCbWiV2Z41mdcONJL0QvhDkrTbJTNZ2
4cCUonfNB03WWuStH3bm69i6ImHtMGTOKIEyxauu0qVf7F7sQ2R7pJKeT96KDLsXC9zkJzfSNlAT
J6JAyq/Xv4NBkxG9VZiE/r3jfAQionjll27sc1Jb1stPRbab3fz86omviY/ktocyk+hOKeny/GIq
4BvkKa4ksmOTu6H7wlaOcyEbbsbiVSFaZ++tTApDZyqbcloFJX0mz+3m/pI1Fht5VcvY/sqHu5Ef
KAbByVm2jlVWJZtfdK8FRQl4fnvfUTeDBVqbJ1iF9+nFzidPL+lC7mcwj93FavhNxOMs4+DADrPx
7O7jlyh8xaN5stZChURClCwCkwp0eViO7AVDiCQsM/b4qTx9+xB6PeeDI/BAEvTPg7dCI+ajCak3
3nIpcOjB33JcGTFbTNYYzexDEGcwNlimrO5hpnJvQYCVrltDaLNCDoVIQ6dokLvtuOwCrk4O4tx1
papuKeljFQuEmEfc1CEG/QvscqnUY0ZQOL/CSL1G7C0FYuz35xOCucvZZBH/hAjjY5L4J4cBLIoh
GK1GQ+lmObHNfTVteX94z6F5fHYScZDiIAnEEDpLO9AjLEUacQtZxXHxJwQZnQU4Y+vBpEHLuLeb
NIVlBGDpFsIGgMIW5ubz+SHwBIdXkKbxh0oHuFzbC7oEtGFayCF0lSXTcESPig0T0upb9WfMgzbX
v3HWPZ/qydmeoG60vHePj5R6Opnqhs08EoK2gL39a2MA10u+qhn91HqJxP/wAsxCW0+VnL2wXfwm
lEwHquWLm5dp9Wo6A0f5zJZXcYiizADTUanNd+D4Dn7NXc/lB1oVItQEqfbUEv6YjLJowGhmuVmi
x9D46Gqd4aWxPNXwQmleRIRS0gYCtqEV0ON/+7+c3B8xhkizyQRPo+oXDTzEQjemKoc4g4t4OiQq
raxVA2vusNTIy0S9rrl1tSHWjR6A1ugYRdPwUCvwjOWF3OPLeWGsAx6jQQ11jx51HA8wVffyqRZa
a8NKZVa03fsO1baGfChZf38NZ3LUcigiCi+/Qi5yNh6Va8QsMqW5thWGB0DQ7eHLR+OvGGYTK7GK
/6O2aErArCt3nPUyXZ7qCR6D11djmy8mzig61NwCv1cvDEcxV2GZ9fhItmchgx2kNYMKBg7mLC8E
yPpuKqXOB3GDnTIUYP8dWVLoeb+OANUxtdZMnnJR93gu+YfZqcZN9rqPMevntgv9F8t4EZcoCB5B
GUvXicIjfvM7uU4pcKQdiIZZkYrnioNX82sorGPgja1opcgJagKmHtTdh7EdDI4sX2EtCCKjT1/b
exn9ydwoRKf9xsMJU/+ArDTdm770JxdmS7e0rntH2MfOgrb5cS5+srKBxoWnkzdBFe9hI36WLDbD
5FxmaAElajjBbsSrA4nCsZoDwu1sET+ttBhXmoB13eDkmVPr7/fNyxnPH57pG/AvSS2hBQtnpWb9
RCcoOAEbOPFfLUD/muIVT1Iui1uCfH+XbSJj/eI0LDdwjMuL141VEUFyXyvjedRRnB2Km49IWnkg
KpBNcyoDHqqzDK5QVbU4CxO6vygadh0YbO21Bqluyzeq4t2LxkXoHu3OQpDMyd/6cYtugdn1IUfc
yY1tZHeEdt5kRXeuJASOBrGHl9ZvPzFK68GEZ4LJDfwzVS3dcZmie8fq8GMam11KF587/z5dkCp+
72TI99QRLDJfMgCEQ+oBmLVVu6v/PGVuB/c/daW526FXNrdkFNM+o8NqrNMyw5GEJnMxo6s2v0qu
+79bz3oq/Xl3gefFo9yCEeeeP6l7Y7XE50YW0MsyExq6/UGft0hGJuMrZuUpXwvOYFPjfGWk8FZc
QsUXtdhuM2M+h7Ava0eHqpqcXjicjD1mJHtWCKqOJ7i+0tYDbHeFOrSFmeNRZIhWlhxoE4cuGJ/J
VnrSTi18wFqlCxiUicSFx8gewkL8DCkvuOihyocKrrRAGWoF4W6hfK6qZfdVlOI7+IoG1IEnN+5y
sd0dPiWQPgu2a/74s4f9JLXAyO8sLOBcv95S3WYars7Gcb+UWj9FlnZyvDzFMSat2IoYvCGtf0k8
QFpp34yAvAG2eny66P1RIetbWgp5rbwfwwc3d6+Y1DknOTJqGHrGYU23YEGLSAPD8l3PXxdomyjy
whYLKUxF+zHpKD5BQamKyYwQ6QggmBlxkXaUpcDRRGdGbLd29bVGnmtNx25WtGUu4WBJvjtKbpUq
KShU9kYmg84Lqe7yt3Q7v0IhcGoZnpeEUmHBNEAMPHhjE6BclfNpwyMvWr8QtVYkXAmijTI0dcjI
X/wQyiILwe6MIABQzYEdZJ/xulO+CmdPO+PXnXuDK7DUfTwAXHOpNxZ+2faqB2XCyKJmNJVkNs9K
6Hy7XHUIQ1URLo2a0rhbXaHiFk10QSQesTiwD5B3Ja9L9OvWSB6vh9aeANiEWqesvxZNCpJfIU3j
ii9X6aq3/hgqjTel9m8AXg4v8NeEBlnT5cBHwdhGTSBf59CB59uiamjyPZ++mZaMXnjC0Y+d3pYE
TS+P3T1Hi+c/D00VxkQDlsat2U1+6wUThYOtqgsn0O/HFVOMvvdsFdP9ArmJj0sVF05Oslvjtyhj
+QkJ3I8bhPA8KZTQASVyJQlzcvhUXm6yF8/4QH6/nLU7ixgJf2hJm7Ia07gcL28mfJdLB24F104M
7tn003mgyRRsKfG6/ubUhL3e7Sz3qm831TcJnBsYGb2Caq4T0H2rwg3E26wPcyFprPHxERhOGHdp
wHb9UPaBd4fhnDKIIGJM466nSfrF5WRAeUBFiL+XFUkfWh3utXi2kHbOTj6JUIaWO/AUjZ3AUqHP
G4DgSDyGDQ3ADvvDpIN5+Dxapm0VQ5cuhxD1MgiQUdRfbZZJz3Hwx8OQfhabRG42Qta+mXDWQ3mS
lLf7g1fEAM33x1mfdM9Vp4sPYfEQV/BC1yrprBxHI1JGPaO30/pwnGE1rrsHSrprkLb0IMX3gguw
NFpCIGrMmNjozqq55sBrAua5YD9PIAFICb6hggOxTibVz7dV8jGBKPiEYzZzRHm59Blw3CwN8Uus
RSeYHg9rfRc4HR6ddT0SoE/FnGzWZwDCPmunqJ9rUhVW4zMZkUmeqo4U1FExMo3/yK9joMGqOobK
tEAqth31jtg5DRxHEea+FzbwtFs/dKweO2eVFt42v4uw7gD+G7Wme9MxihnCgjAJTKBvv1n2cgwN
wLgWmsQ8vwJDRqKU7YlSDvLtlvXPyCibUoHQdQRBj5LSnhEdKlS8em65uFpsxJeEuHb34/gjDwKJ
zAClUxRFrQoq2F3eWxZQGOIYjox90vo5FiK5k1w4tb0Qk8xLaB9Jl4YTiGrecsNcjiUvkGXoFI0u
p+XxQhmGKJXeELEyREehut5mOZgR69FTu+O6OmQkDa2swQCvySwqen9/3+h0e9WFMlH+xeKnD2Zx
GXkk35328vDK9U7IARNJtMWlCor7gb6E9XNert+dWXBPWU73CQ9j2Kul/mfVALiA3C8iWepoB+tt
f66Nmr+BVM+iW130bQYdUlhgFT1gZFfv9G3ao+UKcgIbvJUItB0Trj0Y+nBXyxv690xySir+B0p+
Vj6uXXJovrl4swcLP3E3o2BMRhT/YI7r/DpDTtn6oWSQ8myWVi/eIPhVfJhU9MXQdtuKtXrY8U24
TfIlZRspcs5298IOcFContGIfAuES2PanmHGHzmXm3jyRndQdY+GQZC0YyLH8Y/c3E3af7EZgxyg
OKgdfUGfZniyA/57T0w2CTLrA37UpPRdH9hamAcpRV71p9QTOPHvb2BGlJrTBAB4rhR97dBbgxDL
Ttc7t+X6ftuDM8X9lUhgD8ceH1X71QCU+49OXtdsLv/fpo66NOuBW9zjSxhOT2onG2na8IteI4dD
U9RDfmRtB/uQTTxdRGfN2nhPTuQYcjjSmx5zr8VKcz+pfTDxZbOhK1NcuPlzcdirElnXlUL1LKeA
wrCrKmOjrKBXQUH1rssetNF3d5gkUYxMLfVx3ADkjSAm8o5eWY5GyHBRZtBeBEfufBYxrNfrzTFc
6J5N+JEC3As4nLZO4wmVFIowBnL8lanr7Ct5LTp0OTnjzNcwn8BkoORnMUakOnMee5BO8gwv2pLZ
jD2ugAN94J4fHE+vV6qoig8Dhlceqjo5ZizJNCaxaZVqbu7Fdp8ySxQpPSbEH/OPMmMkV4Nhm6vd
3FKTmVMVEwleboAUCBgrfeM9tmGR+3qTobhOzKYmCeTH/ISFP/uBUeF5Ts53DDNszAiUCLtw6DKl
1HfgwEQeIGlGR/Ba3HcalOzvvt3z/J0y4D/MQYNPelSxG15zvRE/13sQBLdgJGI72FjfPIMLj9zk
ecVntRkeg2DgPpIaRh/PStUw/hMrk+Bd5ht5cuHwkIlBnHSLBsVM4ZiGcHXb6OPAFxprbg9qLQX7
HvP3JYiauBgnk/eBJOLQG3F+1qRNwERtvGR4gVVw0kVqIbMf2vVH5+C4wBp1JUg0k5DFJ56PFFQa
FCiVtSu32j2ZkFxfk8tyc2tL0jRi5xtRIAXujsrSGgor+fihmAmeRBvL+8nXXMRdZmJRs5iTyowI
nrGrM+6RZNsRnMnPpRMVtqCObCNSg3hgYIk1Nbr0roxiKoQAYeGZXbcd58HXwbph9L7iSRMRYysQ
xmp2hDovPQFWS7lzURDMOhtt4kyYVRHlZL8lDsdMCt4BCpWCJfM+MmawZEUssCtQstQk5EBxHWGy
rjQMnlSJSj9oGhvgGYT22Wz6HV7/oCAlYz+EdnUu3OAT+leHVdpwV/f7n1NFAEaTnvMpOk/lYwNB
0yEdV48VhhcB71iD3TDbE0ZKWVgBk9Wp5tv0ODkXs+7z4a6mH8TcLZVsM/v7ppw3gUY00p7qTNhD
P37TR1Is4rKbFJzvQd0jWnEUOuZUfLTXkawsOpa5ZqKXcClPvstGt6Cxx8u0o9vTBcQMoHbBTSzn
P5dedu86j1U0koYliibO5ox1MbdhfuK+zfYD4beO99AouKCeU5LClC4gcYaASoG98M4y0tQw60Y3
Kia8fgZre7pujZNBO8hu5Oz1ODgr+6uFJ35+c1FG82IlDMuOeKtkLg3+Cux2BG8r5txCIRbdoCmc
oWXlnOem3IgDRfYSwQjxNtz+P0+soyBfNaTpfosEZoaQFieVVxV5+OoQB2SyIkK/GRpSwOQcTsfm
pN8dkw283gv+jCXdfxniL8HOud1iWNpilicUUx6H3e6Czk7qqIQDtM52q7eUZtIp2haTF7HXZyHc
h0hFpU89C1DcEwOn+tSmBE7MI7P+cahEveIvMoXqaypcGDuKt2goFoneuup9vucGzulI2B9vZNB+
DTHZkxVZwXpTyO4pWjjMJkRthPnCJ2Fi86RtBr8ADIpNkr0TNw2Q88NYKAGKiyk3gtxfeXw6uiWF
oUPeLOW6/+4XZ5vZM68jEfVMqkp7Owzpeg9AULNLe0ODRnsHUb8mZ+uRQEA7QeBeKfk6hVIeOVKt
33ujmeaVxguJMkbXdSa1R4mE0klXZZUmmnS/W1Ufs/4rYeBjIzecJuu7Eu/mO9naiXYXOxiIACSe
fbIo8QYy7z5wH0+nYam8JgV6IhCPO+Idpq7+lMrxebU5RVd7jxYhSmcYi3jDr5gNxJ4gK31OSATg
DsVLBTIrxesecMGYQUy+dVenwyqf25vsSX1yNqpSPBwHaAFPEXaDo4PAB9YwOPg4xS9QNp2ePpbw
4s5IGQe/ApENscipA1NmEfX5728rvl/l79nzT3kzw22mXHBnXXsOLmlZsYvaTV0eM2tlbby5sYg0
jhf6xmSC0boMCeqDVlyJukFGx/yzYYZGFR61u31Sk+d+Fq4Bq7YETD31LE560Yj3zyPfOGUnPSJa
zwTUH4ZdqBDxA5gKhMrZuL8AT8pyIBysLAYbGMQ/c579DPDPHe3scKvYzSC1aBqh2c9q1TUEzBhB
EjuyoSPH5R2Zf2c9PuAqqdxAX9VDeHgDSg7sVcuhWVumBE6yI6GfyBaIDcsU2PP8voaAvSYXcJ7x
A2wHiFmO5Y79w0w4TFqCsBJZ18xe2TS1sZp+xhh5SAPAmStJJxCxOI87Am9G/b+LnZo1ELozhSm2
0vHwG6MCjWfs+/eMfX6yoRIqFfi6sGBQG0Bp1yBjkAbKVrgDIF0fc/HyqJ530IEsjRr9844lUgGL
goV7zCVGZNrASXC5XpOoVHnIlrOf+GGL+dh5qrcyE6SHr9KMAEmV+ZjDIGhn7UT//Z9Oi8gLLm8A
lzTf+5cK7gsmXnKCOdDIaERlP7M6A/OuNTLqFe5PdJZHJukbJNnoqVVHZbgR8MzEAnM1Sd31M3D5
Id1szRwWXIVCcaaUAFTiIyZwbUurQfelZOKq8+8J0vkCFOKIbEe7Td8FiWmJvOSn18zdLUWOird7
YR7GRc9N9EapMutCToqNdLKDR2EtM3hRsadBb4Yu3OLCdQFuS6DWcCN+xksp8GxcSefUoBERC8lP
x1LIo4wU6MY+7rFaZwhFg5pFPGUsIsUt1Zz/Zb2cJOH3xUXOAPUBpATfj/tyOir8x68uSvREcPfQ
uY0XjC931BLwjtMPflrkie/civhKidqkjrokd6rMF0rA8oeHqk6jfgqZUHskzKLKnC67sgO/D6Bg
cOa8m0xFO899xCGEEQGrsvQ1sNN4gn9lsSWRf11j93Ry7DlbtUQGX10nUYzliamwyx53NcMIh4qT
xCsiIr3LG+lCq6TEdu0Z9GFXfh3mq7027Q7gkPrhf+C4JvezeA/kA0eA/3T9bRzzXW9b93gCHjTe
PuBgTabemesmpW5RU0MxbNeGkrbJjn/AvpJm9VnHmFfti1tncecR1er6MuKWGBw+W/8QsIPA7b13
C8eu/CBMGGKACL9xLZFlUh50d3cdMAmWu2ieY6Q3vgo7xcwf4jDnMiv3OUe5bjo53gCOFRe3qzy5
Dpdyj9qpDNTbNLrrEYLg4QH84yBmfCCqt36i0mdv4n71kjJZrb9QZ5Fin0F40xTX8S17z6vNqG0v
rHkVv4TPNrJonpADcfGNDcJ/A7VFfufrQxd6RjlPwIuwoxpSGdZ7m72T6IhVXURINTEW6slZ3vWf
Qq8p5HtYBCB02iQwMyz7/34VE8tl/n9SUU1txB+BQp7hRqMEAn9Nqjh+FFnQtD2hTxEx4LVMfcka
z1kJ0I5bCoBX7k2elh34tb7tBHIXdBgOXQDFdivBLWFX8LBOZ7sgAMypEzcliDfmT4MocbQP38oI
EIMzNVOthvHb/xNUV+VdjRCoRLcwMcgQ20Bplemfkzgvq+P/cyEniiodkakg3yXM28y2llUK999y
7tguZ21uR5mUMAfHOm3wmWQSKOEGKvyu3jS6zTBmth5j6CSUhFLkiYkRSAHkge7pukReohx34EXl
aDy5GFKiC9uKzyUIGKgJApOVn1QSR4r+/dYxofIHz7s42Gg/oaWjYomzlFm12M66zLEwM8gG+6r9
9tA0aUUjxjzlIXhBlZfRDZGrQpWqia57QcS3Y8cjjz2KrfQPWZWJ1bR3CIM6UYL7N3z5+laODrbP
6hzMCI93TWpVXL/qjBEYp84Q+286yxNG6xDvJAz3SlNtE7UnZJCFE1L3x/mNp9F/RrPPz5a+QXVS
Pe63JN2V4v9P1hI4t9XVtzz3eri5kdD2uj0BiWy3eyRoLuPS9EcJhahTQHNkD3O8qzx7BzflZQWd
Qg0y7VCLhlDjCdhgcDCJCvVdyeeUXQa2+uV50e6vxA3JTeb7F4U7YICwNoz0uKY4XWwqL2KJdXg2
T0SVmPQFtiPyu7MC3L48DYAnTtcZVM3cihkns47rv7O2E3XG52g5VTytM5I1u0h6NmhflGUepmiB
gzhnYTsXr9mRimyktcvVK/cQ1G6n8pTcS1l1I+StV5UcRwhJh8UAYs42dFNY5joqzjXhLzNIeSgJ
z2vt+dkLUTp6GvDTLUOy8yKdKmFeuafAC9Q01rz29/KtPDryoaLK6y9QdP6ofX8jYWSVV+8OCn6o
3p92vl+uQ1YETFzemF+hfXvadfCIiWsW/azkHVAN2JnljhPwd6IGMQk9SkHKlx3UzIpFT6QVsTqM
iP2zkyavw9/GfHaOM4XKyoC3wrY/V/AGvR7bCzXdkz+HZ6lfrSbRujpJllQyMgrM8/8FlLwEj16V
6k26oa4pfHqGOEtvBD9wn1V8Ug0VlDJrv8kYF3YLpBqU9UhjNg36Ll2Yo67uFYiMJnm+N8lOiKgm
hEoLwlZNRlw/n0zekhJ5v6IfISf8pFYL+pyU62MC998rwnILoAlRRwCcgo5FLwBsbZLGBLxp22au
ywN0R8ex4crW11sSpyAjcujA/+NvNVkoUF8vodLZHE51hpAmS9y6Bbs1ZcNrQ4VIR49mecze1j2/
W1DXRqNp8HiYSV9xm2D3h5aK395XjHNh4LmuUGorPWPPyfvnlCeb5EnGBlAMCnfAPGDQkFz7hDsf
3SjMzOYQlHJHZn4OgwxUdh5PHgDfrn1pLrFBE/5liiT1iynIjKMDfyaGWqNqsEiLHnAqE9syvjFL
6YGJR0V5JV3zNxKWVI00b/lFTpWwSlOfVVjQTCrxdKMNq5Op8tvvkAroZHnhQZZIt9CoS2wzEUOQ
eooEV0oxm+geXxCSL2MXshOX3xUPCd+cgfBZkh0OzcZdaYj/q2pf/kmL3uKrebCYT4pH5ZUTTC/F
yNI8AGpc5ijkuZTSNQ95MSazXjy2KoCXLsBYi6tjT+n0rlvpWXWhiBN17nlIqEdearFbRdmSb/Zy
I992V13o2iP4y8U4GYprzmkSoOAjtgO1XsJ8rOTY+lZ/44Ht3Po+2rtNtycsYJdSix6kLGzfDQNA
J108pjJusnPa2JRMpEB5bu+16M9Lm8XfLYFs2YyAA5icUq+j0JLCsRKFImqki2q+z3pQqEM4KgR8
UUKJAM6h5O0NKcztN1qYvvPUbycelnbYstOF2xnCnvu+Bo8mz0by4TJnFfmgbX8T1yBBdZcKcaUE
5cawk7rVO+qf2AAbxqxfrZ/T5ViG/AW2gbMZWW3N/sNlhnFGefds91EJ2LSOhmbET9FK4S/1ATl4
dn01PDypTNIUdKS8ummR+ess9ip64zKwxttgcT/9zSiW56jtaxhkJv7760E7qG9nMpBQEdPKX68S
it3fXm8rnX9meA9xiBRhaOIwbauIajMtqgpUy3frMssW2m70wCJgbprqeUhlO2BRYMwVExubrt9H
nb+tfNgC+mrH+MzqM2jTknU2cz5G830BPRyaZPvuL+lOtkR3hl+PeOeDob3pzBR46FmNCxruxbPp
LNgjKaJnyPX3BWRI8Pahr7gmyPlTYQKVBYiziR1MQG1wtOtmxOWtsg9AOkz0bUYNHzLzcE3d1MF0
hr4N0IHv+LwPIv9He9k5klUasKFgVOmlz/mqg1tpev+FQ38g0GtCaXddPex3t80cIBLmi1qRhsv5
vr7zkBBnmjO1YCc+ogmFH+W3cp7d34QqjKOCBmEb3sasKiv7rFRQIOKVmJf+REPyL0I+TychgaKZ
UrkLF7uQGcXRlILDg11Tygsr1VDSnljfp4EfDLimVnCmTc+AS+lz+Wsw2gXHha/FR9n1MOqP/aqw
8OoD/EGtJl+Kv1VTYNRH26iZhKTkMKdwVrdykYIwwEsoBseMmB7SaZ9bg3vKASealqBV9epPMbdh
g9ciCgBGl0p509G3yKLdOuqEUFEX3I5L4IHEf7CThoesAe9ZOWlhg2vbuBMBwgqwttYS3xvWs9zf
v8Xu3E396XM3xLykWeWnduwEJp2LXSu2Mm0UyWeONmESKEYontNf3PzxY99ARJ5eLdc3VP81s1Qu
8LcEU9STJ6NiE4rI+xvlXzmYuHyATDTMPySotbtfX3uvvk47nCcW4PLtQeLYHhj1gs+MKh3jkz57
WEIk9WRhPpbNRlHJv1n7tg8xPhpJejF3RQGe4/lRvdGxqrtlsLpNWpRtEhmM5UAHE4MhD4R68hNg
cwjFr7MhzaLLpYK8CdaF830IxUVZ3T+qtYIhhN+d5AqUNuaqukKq07Zdb+cM9i03/YCQd10AnXgx
ZNdnRNAuuFBa/yMkRUYeOzVTBZ76r5kjyHhSCWy5LJZvxyCDFJDV+MKlE1ebFHY3q7X9BjBvtejK
gv/z9aa62EVdiLtErv8SvlpDfBqWOxCQOJUMr61jGy3kbAwepAjl1tb9eKxYK7pC14sEB9YD7WjB
YW2KR2HM0eosPuOWMtfJ4uo4luDsZB3p6yLUNhlgcTEuL8FZMyZwDzlg2DJ4S43GMwJ2wcLJds+c
REDzdmh0Qqluf9m+PP/AbtqYT/5qQ1mCg7hXs3X9Usc+NKw8kQBoRComZC2lspQIVifWzMpAdLwa
vCzJ15E2bE3QWtbkyHMc6H6HaHsnZzrAtR8jOL3go+bQoXz4T1njPhAwisrI59DfxcobTQJBG/we
hS/NLH5SV+DTyVCunzKIvXrwLKygiSdGi5Fa1PWLaZlvzmosMylZVHfQcf8Cb5ZSzDdppErSWhES
1LGfmEXGg443APbfT1W+IlFILiAhWU4ZJ8i9hQtEGFXcy2/YKUEy3JQHFWywbqMfwwd6aZ+Zw/WS
JBBmztcWmsk8MrdjU8s18SYVrRxK+yjQN3bCjdOfA6m9xjxY497IVXJTZZ9a4pqlMcn0LyGKFAdY
czWRII4N/njTyA442dEgWlW55oT3T3vxfyy0AtdIq8QGZQS4q61QgWGb0rGAKMc/rsftfGBh6qEV
9wWrFrtASzbY7OAOcjpOqyd90OroxwXun5xDqWWLQvxCPx/0g3+8fjDP9goT4nU4CLEpnFp4F+mo
CEzG6i62OaiEsd62JrAqMW5pqfUyY+TeZFGObf9eWz+wQG9+yLNf7/J/rcLz5T/X10Asdw+3hRwr
s0pVzFIIGjpf5wAzVEHNaLjhp7UtJ8tWktxjWzMmSXeXBO4Ofd8mcFfE6dwh7msCwxQBChBxp5n9
oGVIGiIjuNmUN7mJgE2VDOX4vOgfAYBtlirr99qvtzLoVcSzsWDaR5IDaf2u5GmytwLs88D7GS8t
H4wRg3zgegkGP3G4hAgDXduF6bQyvChbvaTajdFCjlwFaHlbpGoQurCsiPjEm+GnHzH9eugFQnRm
CI13fdbBzYsHrT2kSovSDEgEJ6A3qvtjcT/tk9nTZpAS80B0FwOw/myrbr8gY0KJ0hTzipezg520
QA6GvATJMFeQmTytC7+xcMugw8jM+r1cHnSvK1xusoWiTHrwriuyQKW1wK/Y69bnrzR7QmO8x4ce
939JFZzdnRrX7cHj2Vz450Ov2T2T1YZZKLDmNfPOhm6uKhLQrjYfK1XpxlhuGJhnRhvPqEl/o8jy
qjwS7I7MOiA6wmX3UjRE4ItolMdPA/fBspiEzPbbr/x4F9ptlu3hxHulDY91bphe5UxZOeSJORvW
h3dA/P2Ce3VRVLg4qtZPlzXXSncoWCWLUIIfx3Q6GuHKAcpy5R7ifx8Q3K9eVbVBjjkN0sb96PoW
EicD89c0nenOVi0/jjfiD0eyc/RuaJgbW+XaLykJTtRF73Gqy4W5o1l/NRvCh6DjwSn9fSKXYy69
QXBSemqB/RFXHwul814qvyb29jixCW26QJDDaDQD8w98Uz9racyQLbUngM+ETknlYTCgMDHhojnR
8wu3hS7pN2CQRXQrHnKRZAXRnXSLJnQuee/z7U16aLVLoRfItTPq1e9d3iPwrh5N3JYsiswix7pU
brgaOf+vaVt8BQHZGtBQ8PDOT2hRaJ2F+v3ibvA8dENUeCww91VNPbkld65vI3+THD0DJ0H7sApQ
ko0i+LJGhbApQWIbzJ+AGHxOD3XlMZYjZqAPMlhWu3MVJXjCOh2qpKdvSX3OHz7e+2gjXyDcnset
g3E3LRqWOnVZ+6tqQrAN2yWB+5VdnvWZbb0uIKIfoHQQesfX5UUgnoYcGoare6/bFnKx2lUoP9CY
zYriVAMDZbVIlGnKZ/7dJVoIYGgcMVozIZdiwElbHxiXWOzJnZT94p23gIi1887zMuzTjv69wgDd
SCgaoHom7SUuEXNeHEoxNIElQx8eeUwtSRgbLqmoKSbd954qRLg2RAN26SdC3fe8W1xLQCWS0T5M
cnXs1dD7FpdI63YK9ybd6e/wwEQJA9QtF+P+4hcTRZ0fG2rDKtCXxNaTi1keFc+lLU+NkYqTvKpi
9eabJ0DkRE7+AxNV4wb7CpkvhruNvH+EUcvnzP8OJ6LwV9YinjHyqZ/A79NnH16DvZfoNto2XAjM
4DmlUSk81hkDpvf7xRSMBJ2owickFckwar1rDjEB8YSnYz4aBf/p7DK+7Ydc5Nl28fVpJbJaXMQ3
dIBgxWOsvYMV+aUdrGi4A7mZJl7m7RkaqbKiISPIjJIketeOSPR6fYRWo7cv6ZOKks6FXZpJt65s
R8HrpMzkjxSOCB3OStGE5R0JGOMdV7j2otYL8J4Ya5tabu1Oa4IaWf+j/jR0lFcum8sCH/FbNOJV
X3HQSfrw9S9Td0VwL+X6WE/v1Ltff8Gmk96Y+Ifhp3gJMQqx1TClH8WqGCLXw2FTGYKK/Gg0cPgP
cGDQq4+70Pszfb2bY6oujCtopN5E8hnT79GkqSaDZORrQN4BF/LoG5AuBk0Yg1ktYAZ8B+lsHT88
g7pU3CCTvXPl6u9GslDcoNSgV4GhQ1uDA1nH8D/luT4LMxLjqYM3xrxoS9cUCol/3Ww9kyuEhqnL
BrK7Y6hpoB5Vs5l7EBUpJ6wpFo3brLSDUn2BpxfC6Kv7xqWI4thTOh/T6TR0Mfk7nSVlLNDnadx+
8IrBRyjUQKaTPHbxgOb9+4ImLXs7uT9o9SSH+gDGd21B1xs8uS0UGuS+NZMsqpXsVqu6h1PhF2Lz
ar7VY+fuYvg4+r0DBa8ytG3P1JVLcA5r0AZTd2Z9IKYGI9siirjMK6QXH0Zywk3TKQCDtx1L1f7J
ozB77JE1rFs0eh7B0fWxCy9jNIvo7kZGgQdghWntuazwNCStghPtp1tEr2oqJnbjMuzm6jLj/qHF
W4vaLJMMf4mJye2lH7IpyhrSSz6dVEA5rO1d77aPD9li1m9SQ0B+mbQ82DS3EP2t4iFHOBlI9hAx
HbsSPdW1SpHt3Ei1umdT3EKRSlRnqU9XopnpozXlquPGg6pmhw5PvJqX1ecz2Kxabh/VkkmYhiit
ApQ3dMHvrMy+IeubcTJblJBPHKUOaltRsH5wh4mlzxArnhUgJkGQzYbAzKPMLfW+6LBoDLMPwAT9
aLO+1dxVsEZN9d7GNDDtwV7VTTEp+Gh7jyLea3u+DbbdAFuaCpnaDi+YTBMlK8r7bLtYSu8nQ/cQ
+xtSmaJsKES1uCTU/XjyX0fRCd5dwR8SAGstwg4Pb412flQ3WxfuoaOXrHgW2ZBAXsQZf3eEt+H1
TV/H8RvnjOoEBCeQsz8wOoMH0b81HOx9Kk4l8A6R5dpLoyQ1ew2tHZOkDYSxlT9cFLIQSYgVvp5n
4eOcatn82d36dRnzLEAAVNl/O+sLO589Us9oeXGuy1UbvTJQ+3ZFIJVD42zm4r73Hjox/p15oe3B
pU61Ze46bnmabulUAo4oBjShGUBvgPGdCfgALw9am1smxTkQC1Vu47f5K7LQ5T8uv+jpZmBnWim5
Q7DyD6PvxHwWCqtO+600/XMo7lxyGL57m84aTg/oXTIpSEfmW4kUHcDNQLIKeVpHy4q6HHtG6Dr+
GMF6Vwq6lT+tKebWy8rJVl0/MZ/5e/pGjbth7yVKPfBKRf+IFgd9XA3uo6ocmfUwBgm8hV9wTSUk
ElDUSDjjSnfvToQR0Meq24F/APGqu8BRZz3jxsKX10GKfhkYB2dZcerO2G2IXY7v4Q2Ux1nUSmNa
W/geoss+DR/KBGNJBN11ge4Tp7VQ7M4NP7VsXSUSpdu+CijT1syq/Wu4IbJZ7LDbG+s5KvzkQLdH
UhUy9+tWXMcB7Oa2qibiNhJW2Hyc4M5TptL7aTU9xS3KqDgAfXb7paY9eFx3G4Hm21h4j7eyV4sJ
QzS3V1vu+K88XO+mDQOvd6dZTz5PGNZcuiDjky+57mcUUyi8SoZRNAg3NLz+D5yJRnYJiaF4kwTq
UVwg8k4f3fUDHvcjFiiPFbWpb7nMbtOsUYd4mu8jKr+YftKP25pQIH+MxNdjZNi8gyNb3Q2ihlJh
lgQEGvNXMO3y79ZAYZ2xPeG+LZ/2WZuqeX51j+gSj4lbQyfiErDGupUIlpjmwaFBxGgqQaZAC67v
fZfWaGbSdOOCu3ZTnEmSIXfflaBu6DGGlanAgtCKHq5tw0q22lYZ1g7kTJXqNLNGbv6cJd4uTrYc
GSSGTBapyz5zkPNWEuGZYvCBaGAsDtR8+pvdwjgeLY6rFpcGbanyqeRUzg+cNc+OuR61C6Cc+dS+
89ex3bgWrbjisClpgjVkWTkaKxNSmqsfwzlJ9Okzw4myU5BIgbvarsqXyy6FsTswFVil7XattXas
wskG68LvcCF1EglzTFnEGqFa54l4iKoNt/Q9PhPCCTiEPqmoSRN5vkdxv88JNpYQL7G89K6KEChL
E1k0xuAGLdPfjAaqHcW8AbLt3Dh4QJPXD299ng9VNRNoeCULDmeqroUWj/dBFCXMrztgrzAu+oBQ
WnsW2dwSQw+w8nZHE6aaDMTQdoVEOQU6kFWJiERuarVUPgqEMbC82lXrSApjiqwrZmnXyy9vaStN
Dazd7vIMrfPYDLKjt4BkAwe7cqovkc0zm6SlrS07IR2mGMaW/GZeikeeqazWO6YMNUAdmg9zZPsZ
6xIDYzG3vus34Hg5CT4AXeq0XMUmC6DWTDNgVFeJKCNBLlC3mrqZJiL1NPY+y/3azoVweM7rRR1f
p9Rpud5O+7/tohKndbkysW2PQl/11DIUchZ2I/lXgKTBGLFkSUDWitkOGQgljxB9rggFICs8CDfx
1K2/tFpgeBZzUWlLxnM5+R5fc9TK6LHy/NJP6IvBAXQEEQi2y/gFmILlpjAGHIH4VcM6lSagLaO+
1LUnxZjVFw5YHBmAQnyXmbW4YnMIFTgxhyliVlFojzhchCQ5i7byi/Bm+kAs4VVoE/hXsl7WbxgW
bobuQMUCA6i3N94OVq3xR0SyuDKL/pemRULw6WdwOL5RHd02pcXNrBSecAO7AVh9zhYqSgYZnQCW
iUcFwSERC9cw/XfeUzgSD34qrJa/uXg6sQ7jq1Yo7LAjl+E+imviTgh22/mFgu3vS7tWEvn+jMCI
TYVeSFjZ+SgcRJvWh0UoTzRzCpGyR3/CM3a+yQUCkj2BEuhLU3b9etOZDWji1nCHN2/ocnaU9T8E
y9lnpep2NvyAk8eB9vF2deM4yB8gvI94u62YMNWUmoX5mtU5XrsL1d/djwtYPKIrhPEOQgG6NpIB
qgy3jiswEDObo2kRNDsPlIxY+H4btymEybJlZcnAmZ9+QTkOGqo2g8jIa2QUA3YxoFht2MeI69HB
kD4hUe5lvdbkxa+vh/dxrpHEoy1bGe4HG9Yv/Fsy6x/cRjkCLHoIehb4z1PigH4fHRdGUPKvreKd
nqoBy9w1HLPV0p3lqnXUseAeranBrysZRy8k5jBQgNi7bBUXXiFKXvNxcP+q6qalp7ncXMVMJgu3
F2iopP/0XHCeP3ItfUUwL2uavQO1KV7ZzK12HR4vRnisQEq6aC5Jaq5pMrDIob8s5Yopvec6+0Ta
a57Qx2LOF9kgY9/Ggf+wYGtaBELuActrA/Qk5U7IZ71ArLqV51CVSmwCAx0LUCIRjQ+2enDhSHAe
Ap6opCOqOsHydMagJailbAbxbmh+pb6qvpqC/GR7nxQp8fJjEEYqEV8GUO9EHLtSERcP45VZG+Y8
Rg6ttRob/s636mMgbj0eiDPpkIbEG+EpKa6eztJrSD5oeDCqQQE69yuUxMQYLeD4c9ozz+MdhHrK
slj6dHIt3yu4OC+Tk23YKy8IWHcdiBy2Ou3JfRsvxy2bRLT2rg58J4al+iurKZM0z1A4ZnhjGcIM
nPNgCRXFo5/AbPDg01LdsPDArfOw32wCiaTy1csNCq1v3PsRzK9+brDK2kifa9sF4lbrZ8+x2WEa
ywkqIJo/qZYiQ2OIXMtvgBD+Zj++qs5uHnSYzHdiF+UdZq3q0BPO1HIjXibYksdnTrKUrJ1GfodI
hhwYLMITOmF+w/pLva3Fdr1A1Bs0EW5I8k0wWckWUYlbn3h0oCrlYwvYircejXBJ2G5bVkfXXXLj
oSJt3VvwiPMGY4TEN3f5Ar0wvtp5GCZW3+ToCJueMkEmC6VEJrUs1nBEeYFCLbY2lW64bKUyGRuf
KQxTmoKcqUf7boLS6yh2oyi6JaWA/9EDEQ5pUY7w9dY1aacV8+G2xnH29Xgo2IOhQVYHOmsvVXVm
y3XfXKen725NqrHajQtA54/m6FpP0IdVHSEjS4VjMAGML0L3kKLJbHyThjQx3BertzdqgaIkTnuA
cf/L0sLix4o+owkqoQFYXRuquf+JHGWA2UkSyqUk4VZsy9TVaGPWtVd0ERoHS+P1AVSp0mV+bKty
XWPQWI2fbcPbEZ/KMTHvsLIrzIqAgmrN7BPAj6MUwzdIaYdRgr8b2npzcgbJQuRJ79KBxjyE1cYM
BWAzLRcl2U6bZo+5DI3JLP+LRv0oDWwBI5BjIYUW4t8BOfsYo0thnwUbIDNIoopBNCKF9NESs9cr
eKUN9WOUe8QjfXWl2RGRQqi9ThZh3/sukQHiveWEEc9ZjiTPvSn1S3bOFZ/n771Qd5OE4rsq4Cvy
Ha7+nlJTIpMbBQR1QplJQIks801YKovk63wnS/c4WMMMHChjyqsJMeUA0/gltftLCUYFlQY1zDDn
fsVggn+nuJ9ABvJ993muVgJkrQzJ3cbp2wRk5F1B/nmvXa6h8yPaiYgZldHVjS1E0mWzalmNiYqV
nr4uugwTTUXwx9fi5DNr8y2K+bmeasn5barbP/+jayFpSmS7pvimYhWZeqSfjnAq32GcaZUgV2ch
hfBgL5OaVLw/xVuC5dKLwSK2H1qj5mRzqYOeGmwIMobiAbZS/jpxVGQiT1QOC/4UWURX0Fo5g0Gi
6uQ23gZyMs5w5VFFmcMprKD3lQRWKXBuVEtWvl3rioKHcDLcPnwilJPgyqpU0+PSAV0UG4eyT2BZ
jjTVuZnI/csNEutGaX3UU0lnJ7vS2a5uaVj0jh69WnA0deKPiNQ0BOugrV8+ck+gm2VYHuurAgAH
2IoH2Be7FEMmNWEk3NG2mwuSx5DR2/MS3ygbaUpcvN0jnaVZsukwiaMeM4xHXIGyMV8t5TyRhpR2
3BlAtt34N8M44e527qs83Pw3DCT7idI7gd8hK/JBrAvx71BW0BKSEWkn05/Phl9RMsDNyzbMt8TF
rYo5H6KqK5SUExa02+7C+bFp9RCm+GY65xPzOOD3Aru03mzie86gfFT306FEFmjLGlqaPHAzlc3m
vqu7KuzFphDtP/gBj+FUJPJGag/isrQlT0wzTLG7bjHynf6H5KEXv3GpY2z1Yn5F8trSo8WSVF69
2q5SECwPZb20mGPYRaFOTgpgVFh/EKEKYHo5QeuAejssr5+BgUgRXdyPdJ0sSMtP6OEeGWWZElv0
GHMjJHMtsAOXkm3+39N1Yd1pV7+gBGWNX6Rnb42zzQuxTwbvgXiazeBpbZVoJfLc77XsG98AtyP2
KuMwbPtz0/aIA+JjhImdxsfuO0r4TaFZIuvnBC7ayNfhbvxSyYGTUy200//Y51Ac5Faj42QKijIQ
PStxeTb1JByPYLLs5P7b9vxhQGmWkiMPv5//xJR0rwZB/RILzvDeOnJ3aRIuHBjijvyAuS5EFU4k
TiVunNDR7oakDeBLZ3N6lV7WeXjXqazegsuOIHhrZ8NNvAKMQuRWFu1PWoCjaoBBCvm28L2zHIFN
hVrlAtC04coFrs9RdRtVLlSPxEGsiFyIWDIgTrSfYiPwYKC3wovjYQ+zmYTxECwy+0nAwCZpX8fl
oVA2KD0327qMcB9Ptccj86DDa3nX/w/xKmg2U7EhvUAnWweGCAASPKXjD2GBhdHrczbsPvBn4N5r
4JEJBUeC5l63mZzTER5q5vSSEjo76Dlbib06D/Es5lKHwazO2v+4/TEyuWmzTFw5h6b5ip7G1trE
iy8Jxbugyay2j9rVcXlhlfOIyU5SrNx4rV/Wf8VRRyXvLcbDBGt3U7lDqI7sHdOkXcEffaNxcH1f
pAoH/1qbFkEXg+wjoZHjbO1z+2vKBfTiV7IpOAdrwhO/sroMRWz+7YUO636QfhqgDbcLIBXmrONS
qeh9TsV+ONvZLoZwl4uXS/Dx1RsAxW6Q7kSp9My63OzH7K32vu7d6VmXe5hXUnp4PogFjx2s/0Jw
m96ZXLAHpwY2MDpeAh1hviGnQJJzSPEXu+X7E4FhotE2JSIa4zoOjGAnpIcItkQ8p8N3XSo4iTcn
StT6DbLBSH8qndVgxLABwTdXOdrYI4Ngs2AIhp3zevo9BNKRD1yhcfZD3Fm0BaYOlB2odhsjnExx
bvU5FJFynQlSQLit4qhTFmrF+RYhDQxbu3/jVtWtVdXkxUP0cTVNPaAmG1fqbC1V/2mZ0RFwohb/
b1c9JLU4AWQWkQk08dUcUaV37q+RWnxzw9cT2ZOEJqlU35756pPxSB4Ca9C7oybQtH54qBkEIRSp
ObyCiy3QY+fOYA7pKx2Lqk66S4WfqiPhInFgNQD0raIdfbqGzW6tniT10h3H8tt2Dh2r8u+J/5wa
vSRGgY92RafHsimP+r+C445wn/FNYtxg+Fbmm6XpovKiLVkMcuDTEC6r63AAp1zt8zJjXd08V8TH
FpTDAoFrWPQYoPcMltBxi+lbeZqhjwQTMNE4fY6wXY27yMKzqFUuzmEZCN8HV6YSCL0bSyvPCLZr
4xLm3qaspqZEVXdD9iBAmiei/STrRAPQVGJ2Zdv57rpTsqxEpAA0zx/3Hxt5STxkuk4uyoKrmcOE
4vH2yVdpym1+S7V02+4s/rCDsgmb5Tmtfr9qd8v9bSuSXw0lWgXcZN3EvuSC1SXAFmtWAL8cfCDS
7Vf8BYare8A92Zo2Dp+FNVisagZbmWvs0xDap8VkuVhhLzK1CvdXf3OKzqDg0EEJaJ1TDZOVpBgX
fHdq0K3T9gQndmvqH4rNSGiuuTpZmqalzQl9zZVDADFXeCXKGikif2XD4mYntwF0SEL1n+U1NqEr
OegTYzOVUYfbveLCpellFu1eGTChR2Kxlnun49yKUqlc8r/3zhJ4sxCSDjSQb3+aXa5yiXIkyNaO
f40ej/Q/iAJXWhD7smnk5HpnRAY1+DxCG3xmB5tdpKFAVmohCwqv8A7vG9qU7P6CSF9ziNVDHAx5
BpT+EECJnhljMt5jF6op/g6lA+CC/J/dRiisQMxA1WdlCGeWTzqcm+7/vF/+YYXPdPzCiP5Koehd
OkZdaKfVWwlw7ZxxbLqfSMpNyMZJttI0CctY5ijwF/sIvr1389FGFraPMvwWz6mrFPxLNLDrrW84
Ryt0Lp/UyW459zxnMkthPpYS90t++Wf6ATjgdAFjgDv1K9RvLDNsi9ew+JnrvmI+fBfkKLzSCSHN
bHEdFbmb0oggfuuBAcAHM20PMWXcGAaY43FdW5xOX+xlSq4F8HRsThOXLSIJUPBU3gZOals/hLGX
4gvkRY6dgMEZBVo7/ayHt82sIvu7fBCVCn6/jCAEoUB/P5bMHtSrNel4cmDDT5X38MfP0amcBYJG
RnLQ5x0gyckhNKDDElbywYQ0j8mzFtKGigxh9g55Edqn2cyzobJ7ExKyZDxmTrBDFMHn1NFyYZuW
1YJymKyG4w/k+Owv72AKzNX1YyAXS/61vhF/WPFLwTNjV4SzwJus9eJrMORwRQ6ezUjhEN/ILZyq
asAU0uBY4dZ5eK/wbyGp0TLfM85avouXWRq2ySn8kraOTmPZHd3zv8aufMmGm+puYSRbWmIy0kvB
4dfUo5NnxxyuRYUdDoMJbnaGeAqrjzHYnHcoynEuoyMiUOYusrRDdtANXASNY5cdjvSHJOlQSEGh
mCDXaSc37DSszGgo/mUWfeqFT9g6CniHjbDAR65sZNVwUFROxfdsezD/ILQ2lQXo24ggPNWeAMd4
GoP020UYJ4l0PA1rlptm3gtm312eGBnia381tTE67DnsEM4DOmmIRfvsF8JCr/wpOcLxvxbXxhgF
JoQ9pzpTat7ERhTLX/UjDbLyzcaCVKHx2BzkZbJUuxiDvwvBoHFvgt75LlyYxqpIrRFsNYX7gSXJ
f7L9XMR2KDDLnu69tEnG345/n024rgZY5IBqENvNkRZ7I9CvCrHMOlKoASDWcSPYoGChRvKsPUgU
exv+Ncrw+c4LfDxYjBbZyVP89CMrmLki9Ote/4YFMd3U2RntRL3PKrhxED0B4LgYKvsDx+JWBfSY
irsOv+909rSMO59+Hry24sy3gR2YVQhbsWwTKYqjm6VI2NKIwSkY4SDSY4wdDQUFFDJqiw5sgKiQ
u4gh7ePG9w4edMMXo1JBrtpZzJvN3KfWQqSsN9vR2VDp54DxS7YkIjKaKxx7QRlo9l9jO9fpwy1X
iiKQU1RvYfU5cduqj9Ti4sDy+s6D3vKV1vSp3Fg4DS9wXaF9yq5b1ohxBDCQscsvRCl2Bhr9w/6A
KYin6Y02jgCbrHYGWVF9cQsb+JvB+uWZxcaEuxjkFgZYTg3xPofFZQN+P3Yq3mUvyoB+83O5XYLw
CBYKAmBj1nbmf8xrcwR4dk1dvd+lBfZgAgvek1xsj5jzZF6FwOIbUUw/fIZcMCb36krcSv8Age0G
6+Nj+ol651kjB6Bz3MebZ/PviKXTK26OGJVBv07O9mxj2o1nH+BfrL1T9xdF7hWs+E33guM8Y80c
8nwT38LRoO/Nm6ZX8DXge7TEARjwJJKAoXJJLc5armGreU2LeymiJDprOZsllZJDKu6bVVdzskby
husppNbD8BCM6+qcp/qEt+pM/cqg+FYRPBkevTgfhE6oz+smHODFp4WwOyeSZiPJXTxIdSgj92cc
0DUEbUocGDhSOAArkhtuKIJIenf4i36ykVWuoJe8zigewitqf/pgX5mVQ4haOZ3jrYhw/7ZOdZEi
dw7oHP8ozvmbrWYIb+wuenmdI/bZFNvH0VpATxrktz2IdM7YUo1uGYlnVuuuCk4NXIDt4MkWKAiT
6x9J60fpR4ggb8sGB58pAOcTWa2Y6UmKsg7X1mtBt+xWct/zsJmr6JjdjEhVscskt4Pc1x50r7Jl
khDEpiWgN/aftEC1CnHH+wxwj34aSuN1YI3UchyUYYTn0n5Z+bCp86yV9Wpr0rzPq99VCuDz7TvW
QWInpGc668/YpcZ8lES991kRujXNgb5hM+jZoZHMdxbS4honnrXYO2c6d3IGZC5Zq7wkhdQI0mxd
mFNxen/STTAbq6XPl6/MONG4i908gVTDNrSKScixnChkJ6VXgOUr6NqPYkTS9hTs+tnAd+3bvSI+
EFkR/WMCXcu2/8LXT5QW1xF6yJip9olBraPK00EBuQe+kYxd9ryvzgIBYgZ9hY8a3Bp9kNBDf2ey
sNHsxQFSzqsLBOIg3mOFSii8nbeUfxbVYWMPdZLbaUR9x4u9Us1J3M3ghywxHa4ojZdUMHPiUAkr
qha4ZeG+uqI3riEQFjxhQ1+R0GDjj0m1Cwqvpf5VpwM4RZqkLBXPD5rhz2kIY1YdrRzWT6ArRSDe
U4gbmuWfs6X7YkAMzomCawJL5SONeJze38SucjOHenNZVVagblZBqWCmSabz3LaQQx/o1BKQCx4j
s5URvVjNa7sQcsU23GBc/M5SoX2gBPFROSju7YmcO4r0cYZK/APbu/91ZGp2PG8HKxg+oXYWm+As
eUh4CCQmHrTH1cViW6Nq9lqIOj6xlaB33xhjfBomS5mOHjLuD2+Kh4krD8ZSKVRg+c8aRIUbsmdA
OS/PlQDFwWONP/JThHY6tgRkbYwgYr5EVGZjYV/sTdFK0cuuNKVE8uyTv5QKZe6fUB9W90wRM4ZI
VvkSTCxw81k6H32sZ/H51oLTiZmIWsX3JjDFFh0gQRgu+G7kz3OGJuvhqEn6qIh+EIgRjcA23FrP
dYhKs+ERrle2bKa9vIQYXNrO692SwM+PkeTdZahUI2LjAaVbOyD4Ol+JKNHJB/Wyg/4lxxQlxiX6
ilTmg4ljMZfyA/e0gntc1fQHs5owsEhwr3jA7x0SzVC94OqSJs0z3Eja6l+HFkdAPBCsCORcM1Cu
2cyDJqWR9bXoe+1sysLRykeg0yOnzNHdftTXY6lct66nw9VOviFhBVNtFy+hFJknmR8XgfBMFf/y
n8HufuaPOWEhiW+x47oDibR8xyEhpEpEb5xXBVMZqEzCjToQ9wC/DTuaFfr/0MTSbC9jgKOQM88b
6Jw/BJ10f6pnBZTx295gDpNAs1s/UGmO7OXjBLwbQ96QLRSLuUXD9UOQ+qj9YhwL0L2tsyBxJ4vk
Cyjcf+1k8vYTWXItmfusMNw7yG8skKE0jMhdj2Wxqd/uFdqFZrCin4gtVDrDa5HWxCkNb2T4Ts+r
iMIUzLzoZuB2GXjLVGy/xKDZldRRzzit5kuvMX4mrGuxKpuCL/da7A+ap4g5TvkIVBMGy80aeSHH
jG6GlNyjCge+9/jwXAVyxtTdV/Dee5aQ49nDw1+1n16yE4l4R8SRa+2scM8+yIH1GdTDZ9cXtV7t
DBGF28dmc66fb97pAsltLM7THeTPlPfcAHCoZwhGyorC21PYwtX1/Q9p8wPGZ3oX/YLaSJO3SQvb
KCrtxtt3ITrnFaOPBRSQbcu4TFG+WUH7YpgXYwhghsO0wp2oqElh68dD3RypZPRJUqpoff8WbGTp
ZtX5+lc/tl60AEAcQ9Mn1UMa75pe+rwmo+TKyvnZprEk5+fikJ+WCPM6RgtFzaOYany/S/cgt4zM
bkCBed/UHjdUtJ3TInZ9CwLMghCDkbliUGR6F8bYlO3FywpY9rJXZ5ZejuxXjm1pyxb9CM5mRRpf
t5ipLCqpnIyI0Kuqa77EGUr0HNuIjXYCrflCOpJTW1uM54ON9ASOdDxlWHigOOKZvuRUIn9udePF
0MBihA6cL4SxasaWAnFqVH/o4nn5ZVzjDA2qXKdiGWUWaEkE2t7kADuWl+FKkcNWVHWMkRUjUtk7
pKfCOs++n2zKcAqB/etxVyZZofJf6YXgOgkOoH8DtKFWqqYH4SWTTLKVMWpK3dTA5pJ8VVP0IVEo
VUPa2jb8XyfSZYMdLZeYpKalQhxt/el0C6UtgovmtXeuEeQH0Px9Ox+eMLTK+CrskrKG4GpZdhYc
5UKz28YRJYJJtoKKvdxkBtUdxLC++7d86JU8qPeVbX9pmUL2wdIcXMsZTKPun3FerlUeNG8GpIDi
+aIXeozGTYR7jH+ImovYXbC0fS5N8zsEkv1siPQ8AHIGKS//C7aS3NQT6Wwp5DzPA0aNt/sMWp3F
V+P8HBGpkr+H8TZfEEDSby4jEmK4dE6AzvVE0raCzv57DG5tHrAhsPLzt9mKr/cgQAdyqjS62FXH
ImDbIWxXvGLH7mH1wpqIUIMhp6Hajv6OIFfZW251TVTUOpalPZetftISKpbFM2Fkb762JiOItRcy
gMChlHTt+KoE+AN9HyyrprWN27UelfaCgJwj/9C0cKChhG//EBfQ2R4d2jBFAGv1Hv3EUPBhhMYR
G0dr8Xxy9aaO/2/cAii5o8N+L7umG+1RJY3Gcr/j8xFj52Sg/eQGOaIZ3imSawmJaU6sx0Yzey0D
7tes63ZvrufB7Hms1DdKAqZ1IIuMOEKEeNkaKKoRiQO40uI/hrfmV1e01OhSXr3rFE9Ky+X+17AN
E3YsMS6kDmZAYXJZXztI1L3j19PULGI8nhx6lv+kF+7IJ73Jay1gzC4QbSQmyvKK1wsKE98v+XLW
6kEgrKYog+DxtqHSaszUlFK+sy3wwrBaCeAT5Z6gVs0Y+YWT+tOegEdOK0otmjYdiUGWgnnCxn/2
nw7lbE+h6sZiElVrhgMQoRU5Bzi+8NtVnQELF8Ov6HXrtBSflGWXk+3sx1d6FYhoK/xdvFA5/gfO
Hu0faI2H+g/yRrQIlgrwUg+CN7UjC3z91u6lRDcqARwtrCQIWJ3BM2d8IR6vAQosnXo80dM7S5AC
LqIgNHkhxiGiVNLKTukKeGzzx/DsyjD4evGsjm3kXsRJXbu26bwI5vDu2VA2AmESR6VdRnUxameM
haZ+s1es6XkoKBD8eGDJG3TRmY0RLme1I4l2hTtuMRgQI6ALPmmI/nXKukWU+SA5ijH0CUPkEoh9
v8rQN6SmZpwblHD0MYtUB6z0rga8nr68oa947gIpuGvWl+S9UVic0jlObx+xnfcB8sTWutYV9q3o
b3f4h7+PejYodla20ltFS0Kv38BlMfR323rOI8wCT1LIOihFRLY/tNa29bZpV7rcTIBzQnqEA8Ob
Y6OmuM/pL1B/O2Z6xOpTDQKN2q3dByc3G3kww/vH0kZJGCxcWD6x/OKkoJVF0gSLUZgw0Peb6XYB
u7T6v5LUkWbQpkcHI2DHe8M2amd8kWoU44jTl3H1Mb/2W9ZAxm+jUywUNHlzSYajjogznGnvpw1q
npeiO8TNYNYMpdOu4Iqbr7BZBmg2z5HA55YnqcbOIGoHuC0cDL9PLfafjS1DEbECSbY6kgT9cSPE
BOQ7XkN+QCx3qzVQq//mjrkVH9ynr/EbTNPEC9WbI6OT8h9/PlI8iYQ2FMwQ+1PSIu/k1wfpn+vv
+3a6UhhKjxvBd1JdDCWxj/zfVCW5ny4UqkIkauTYo7qlAOh2WOS+Su/OXeyWbQsjgpMlnYG4UHhW
bCXx4T/e0oxS+Ohd0/AwlP9cwY00z1Hi2mA8k5qewokr5paKpl5ChgKCB4zfDf9042dqxCALfLSe
kpqzdjHn8Tf9T4Fssl4nYwr8t/cCZdUR6VW7ubWUnnoQUn/zi4NJDJZjlJxYzdUkXQRsCgGvmPgd
WwuUzu8oMEqYQEwGekYD1mbiwRAskhGATqJKiuCr2EKvnyz75gYl4U1BJ1DgDlE1XMaZuisXNEc9
kD01BZHHbAod029uTbhBd/aWnpYRXKAxBBwT3On3w3WdCGWLGLRkN/5ZUBzHIN3SXdIPrpH6WuEX
QgwfkJOnDWd7UxQvK9Kuw9V7lcQX0X9ZrEQGOBJiOgykp1f9fOLATRUFMqAsPAIdWl14E5mdBFH/
JGpF9nbJ2N3jbDOYcgXpoE4WqPAjBi4SKjRU9n3KxRoF1bvgG3zcVC2dWv7xJXLcREvbLPJvSTiX
IBzEPpQo89L7LpqzEfxS2YuDODhsVLcasNhGIal7V+W6IBawlYjD2V5MVcMEFMwEFoz3XOQaI0x3
KSdMBHqnkJ9EnwyF4y86cMFzANZVrhaDkC5G8ncesnqNGokbDyBmoSeZ5avXvmroyz1jiOZkxyUC
nkFP0imOg2RbttNkk/lbFys/wM0yZJAV5/i36Ypf7jeXlu/07DUyHQRilxJxRlzxFYMrQ92DBgNd
uTxoxSmOGGh96w3Jpgur2xxyYVdPFwGEQ8maEzHgAO3s73gJcOiVQk/MFxQ7RLsERYz5VvSXbyHZ
lbSVFbneIh8DXjSYdtecq1GbobdO9Q9rWVWs5QdCnjlUFgcILS6sAbUl47JBtmO79MqcxWmV1VI3
ICu0YHPXbsCrC18MDvJuYJBvOnM/69hOuDfft35rdKeP3UDf3TrvheM12h08oXVLif4KlsOQjSVi
lgF/3OsRriRmIDN9orFv1SJpF4PtITg5f6erZPVkpMlNd2SKR9s25S69dS5ZZ8sExMDP+WScOi4H
+tvm1WsogEX5+ZbCo+tYgu90jHhEreTDBoWzXNqUum6WjfLOTp8QXfhKZ4d0syS3OJkmy1NWVqwN
LoEwInnehx45vTzEOj/RV5aQJ8IIIm6tHzGvKSuBwODd4ChqCEKa7/qELI7dW/fi1mIXNL13Qn97
KAcfeG11Vxexsv882j++BgnyQfPRJyo4hKFjRLLFNcyruS8k1PUqODgHwwa6u5DkT/zWHoE30Ss8
jMFKvUrVgI8Bqz+Y7TzG9XEijUPl5FLOpsfa7W69mD42jSfNnFMv10ktLnxEGG55afmEserqrYdH
SqPGogl5m+hfs9BsyVj9nBnqG9boFxATOYd1MQr1HOupOVVNRtkC+6akmKnb+yhf9M0qmi4mUIZa
GN7EAly5wkyUElkIgj/cA7mAQuftyquTMLbDm3oT0pldeLTyNmVRnrVKlXsI23qkIxYXqz1sRI72
qZjCFYYE6rxh31CuDKBy0VlLgs8bvwcsJBfsJlgGQ48DbQmVmRW9TNcCxAZid3JoyhBWmRNC76l8
RIr2McKd1NfL4l+oL1Cxz65tsSEKDtUtPWXK6mBBO/zxscWqY4pvVwvsqPBsHs57oKtfcD22QEXt
VufcjOwICLa/DuSS/BML2SiluUdKdoA94HVOSBHCnqXbF893CHChU0qYDghlOwQ2bRKR3oK+5Kd2
7xMiAMFZeo4SASFVQkkx/xUADVEoqasmIfuB2xp656U5kyPsmUN1z4fT0R8bT4dq3RPQi60ALnVu
KmMw1n9aS+XRDW8+4UdAkU76R+Wy2am4wJsZqZUFePtigje12LS0aX30AEAQvWAleLyilbhNVQ9N
s0R1+1eqm8JxfYMVUBQUdDKHOvejFgWeBX88KMV92I/T0Zv8h/fXH0QHmtsANSc73uTn8+dAmcNw
+OnOKKcEsZeavihsz0oQncO2oAXNndGUpS4/um5BX5xoc+IsXwS+mNt/lKNr7yT37ApM9DCfvdn7
4VcBzRdrMlfLksne3sJ6b7ERRCv25b61KZPUbu+fLFi6P8MUcMxyW9JP8Zajm0H+QYZMCRrh3UsZ
PzL0fgm8HvhJmIPEUmbKscdKxU27SoRmll3pE0/jc+Hq9Y1Qu5QdxDDz89qecp4pClismy0jrmJ7
BXwgz0AVdXrI/vngwQFdtwaoH8TQSTN1dDukvR8UdYoc5BemAWKyKaLAd+HdlTIIerfPMSNqHnNU
ysGAvF6Fj+j5zJ5Da+xDy9D5Sk6+bh3nwP9MAYZF09XijMDDVYq1PuZ3V6iAUoYTOKPBwPVurCK9
DQfdl90r1rO2wsjMOadVwsmoGRfEn32JNfj2+e2RxB4cYyNn5kuM/4y7n7VeqNjANUm8E/MkPMEh
IJdPucB8o10bclERw8hTtWNZ+yX/GqBzDRPlnqreljAAR0oE4lMyyvf4qcFzBbQB65cnDbdX3CQh
Uw1spmpQsFFnwK7FFnq+EifUrid0F0YNx1jr6mzA8rTGOVcY505coCSDCPuIrjgdhwUlz6GN1o/K
cWplpI+pBLxgx/K4h970qToTFDQxusQi1hDfJah8W8j6xnOziF15V39vdYYzFToi2Mu4rvBC/s5B
he7FqZ338IxxAHpB1iTV2xgXDiEfB+tJXMg9xkNuUzwgEq0g1V1pELTEhJ6yy7x9NLnm3tBbiZyM
EC9o8BYtgms9CTfaIC9WEqfP5EtQ4dvhPzWoznoSKdipLL1Rl4eBQo2URwWQX9b85oXATW3E3TAJ
8r4TS3+Xk2W0e/UJZACIlr4YxPOuHCXMd9cbh9MynBHBVYZ00jm1vhnHSERCKA6QlM0mRABvej01
vko/MVc131+reGpH3SPwGv4l+CfcWJ99LwBlBweyElLSaD8d3Tl0pdyQe3c3Ul1jKVgHzsfFuCBo
G7nXQqnPqiJ4/Pyw+VJxTT4HvCLyIUEnOyIpI8y1JFdK21oeupqQqbjnLRRiFZ1tBZbYX9oagaqB
fFoMup9/veLzd/qgsyn2QFVc1tMeNm/YwjsLa/yr2wU7E6sHx7uxvdfPV41R3Iajc/ASXk6qiycP
lqSN+YXbmRuF4qlh/oGMp0Ha+kaUYBT2w6HgWatZ2qnQu0P2jDh73n0vDggnuANoOexvVHFqB5S7
9tX45ZXIVwUZuQ+Jcy0ixdOT8130911GwEulfcZpIANpvHA1jZp7fyP/1ryaVIZQQJQJXZEaH0Px
Cx1dUnsra4JkOcLjftB85sq1Vzej8RhVcog5QmOfFiziIKTqzvwitxVse9YX9JxEfSW7naZzm9Vl
kqY3ZNJTFcGHx3qV/Fr5IKTnEmq7sjcbvGxS57loTXDdEc5y5OSFisqNfZNqbfXnH2he+u81jbPN
Mx8UOwg40R7RJDLgLFLBkFGccOeNSqBlWq+j6btTu/UpnDfYhz5pdY6ETFW94bvsp4roCQD4d4eQ
DFlkjWB6vn+eHHg/iFQc5qeF8CfgW9cHnVzlzs/Dd2zlcim6JOBhFhDz0jpzDcTBISyhVShNM7+o
uXhkRB8n0ZSd7qB7sc4A0eg26s2ssA+mUW4BLte8txKIZvd/n3YUambjeR6xEMzCJBPyOtm/7+0P
CkPiqxyrmYjE3MxIqsYDXGl8bRJUO7wJcSCCUGJZPkKg7a4snNT31I9pfcmcfQHNdgVGcPGrH94d
0dbkqsJWKyBvTTSPD6WXMoDQaOjqxrheD5Bi/tvP01fKrxxU5wGxI8W7X9CojCac2ZPQqVTfsAEH
YSgabWSOSK28WuTul4aHhP6vaFEwot9ZEeF8rgiDWiqqi4GLxlDiWOnB7+X2DdVXl06oZDaBtBkY
zvNOjQ7SPPnKOpfnUHQq4Q/FZm7KCREoW+pFE0kM71uPIDqynJDXAN5BlKON9vKdhEagTEOGWu6G
ErNjLMT9Bs7gMiSSaak63kgR3+1zeeW6d6sEVo/WSV5b+YGQ4Z8CVHbnNRNAf7uMzuNFeC+aPEdR
RsK9FlXYOBuANBS5/pxr1QWectnhODEaY1Xppntz4LTNnTvPh9UR+RVdb9y6a4f3yZTcaHS6vvE/
UiRSv/Tfh792+HqV76CJ3jP0p9TyqUH7Wrd/7MKGYGmJzeqph4qmYmq6mPLdjgejxZ/VckN/AZYi
MM7e3wN9GRr8rYu5kX0o4osQ66NEzwcFfj891gOAHIM4fk0qMcla42GW3luID+pxCL06jvHWfqVU
np5dEnkrCkprRc+G1ekBVKl3DP0T+YhOJqNbAGrMRe3cScB9KGm/w3CSkteZuTlRC2ZT1Y+dofR2
H2UX9WXcRCUzNnuM5yM2hjx0ts1fpRNB7ZD82d7ajG29TQr7fTMhAdf/a0vBEZllnJEgWCeLzQin
qhZPuPRP6V/xeeY3MvL0SNKuuzv0QoVROqq+gNXtsb/iWSFV6kJvsEcDaZpPNmEGlO3Z9d4MDD4e
XX2+/4aS2rLPVdDsedvaPdVE9a6kFST4zAcGS+Bq2gc08w3cJoyWksBYZ0dQCZN/QbPOz00FZzVV
UkLjZBIxbX6WiapFR2qj7cJVa3hnHJeOn/FM4VBoA1ug6nSXcUASctgspJV2POKpQNURjDPSB/E1
ZnUEFKpdV5uuMWyfKDl4XbQnAdGl2rf+wyuPFxtRx4279KYRfuKno6aXTGekuJ2y5ypEoQZ3Tu7v
YnSS737Jqgp2WKpMIVR8mcmDkLKyDhTP4xOidOFL5dwwvgJjlohXSFvN3diT4pCcGdHAf4O0ju2F
xwQAd1ECv7cUW4RVI5MenECBUrpgM1qxbwUpnw11i1hyDNU910KKpHR9bhanVUMTNKjaIipIIUFE
zJ0pzMWkw53evHImowZroDVcIL3DRhsa3SE0VvjKhV+DXwcXKmzPwsKeQznDBoisJlNvbNJ5pxSh
qZMUdD/QBLNlFlqMdzU9HDJS3Hh/rDw4meu3f4gr0CKUTLYO1dqP9VUtCWYY2H8gs5Umo7tCx41F
wHaiunTcdohm6JsXdQJRpfYAflf5+gDNsx/ebrQDIr/XfhFaJASOwbUQNFk16ro7GJE2B4n13+Gu
+1LAEiYnBWnA4KnxCBxCfqI8OP6YRC+/5pGEW2akyAJ10Ltoxu81qrXjj/8PnOvlpDDrI0xjpfYV
y4csDW8IUHfKbxX7sFgNtTdgMTgKYfxh9MqV4wxfs2iDCxv+CN/UC376PfXx4NFQxJ0Di+CLZSjz
4qhwCAwRUFfN9yfLaksQXflXE0i0HgbMDxcsu1YWejZLXiFQH7+6dkVtUl5gak5Z1dp/PnvbATmK
xjc1bzf6A16X8e+jbVS6UpqTpSVOri3lIm3S7F4LRuXnyJJ0PDGzuooknaCTekbzdyXWNRPnsP/k
tbbj8K5QGa+fJ3QM86fcnjLBvuphfE6QFTMOYUpCz0fon3KVtZH9bDDl//ek7NnpXDjSEcdj9/GM
xHVTep8chD7t411QNi5mQImEcgY2YJI5NTKNay5dKnm5V+Kt6tCHURrTAlaGdX/+8FhMFN7O7PHM
8u8dFfvVs2zamqUECy4YS2buDG66kBApTTSkrM482pVoBCOKJgm39fVqPWHe9GD30weKbbomZFxx
Gl+ws0yIgv2d5AfrlBF2QZuQd6Ru/JYBSG3WPQ/5FCltayhKyQZ2E03CLXDlNzD2DTbTkCUGURtb
+YQM384QBzoPwuzmk19AAlcf+NwtEWn7n9L5KHdZ4+r8qgkla8DuEjWS37fuwgpxHxNaiQrMUSEp
V4ngXC+VRJ+9+g36BIn0QIQYEdbaMlnhRL4oxbt/BSL7eK88xxUlb3aictFppVHpjIiRSDLwBvkp
CrTqDcKUVkNUnY57y4wzvT2pnqksFUOhj8jpK6ewECL38muDQxGsDwqQmClncwA2GShdQ0iioHKs
EXu1OlcQOeH88FS4g+RLJyozWqLRImmuMnuAqlR5JK/fymAC+d2wq5wCl/7oUrr5kHRC+SiG3Pw6
OzsApn5Kni5xMcc9AgQZriGpg55BvmK+b8bGEavQqwIV0pQteL/+yxrIBYdwKwijfIxFZ24lT7Vi
7SqB0JQkNhVTIjRCmqVhNw8xfno6Fda0oJQS97hfiadjjtyvujriydTEap3axoxK7Y6JQHfg7KJG
VxZJnbT2DPtc5UNpV1tUTddT85XACnbpvgD8XS5EqjiAgRTvj5aSIvYJBMQ0GcO2yzZH0IGrNe+F
OkKgZufzAIAEBdKs7rGlUXdAkokc5g1cB3muYKDJJSEmvkuXmB1y4k9mEpGlGfwpfQUaOBl8c98f
FPjbVJOv0YsgOOzuTV54nEyDBIfgVdsvg2BCv8JVz+vzVGiLw9HS/8grCjDtjpuUz2X+x7mE7lcf
rQz2qgCqUDj1Oremlghl008IQhXRQEds/zNhBCSZhNgvOlI7depx4W08NhTGWMDbwxypuwNGb5/X
uxEvhC/YeZcmVr9IFe8WtrGQ2Ie/NiSzUsyJb+8Ki8QekCOaIwwcnt2ddry7gGNWK8WqJNUJb6Fw
ATgE0S0X4dQlhyrahy8STUPoAXNr7WmLn3U1iJhmEvnR8CFY2obAIAIZ+vT55ciqYbIDMwj6EqC0
EUy+DhXu9YOKFDKO9Mx7yAuQ/7NBPqAKep2bEE7IhFcAbJzgyhTc95QdBpVRAOjmTo2sflFb02nA
Jv/pwWfFENvirB2iq+ZfpPbfm0ltSQ0fS4bSplAkdcQTIiCM24ea0TPzjgVjb6hdxip53sVnBuNc
8g44GP6RDT9396v2NZTQs5Yin77oIc63hsUwwtV3jbLRQnmv4lxvfZWR9De9lU/ach2qPLJBqDM7
ppmAneEe/MlUvbR7NMZ8mJUBgyDfy5/csePmK++eTN+rIxjrloHIrIv8wIeqNbZxO31/zkrvY4DA
lNjdBuhE2ZBETeSLk5PxmUIGdb8sw8rkjO9cbBL9HP2S6Ls6QFtOF4iI6YktsSGDwqs3TG5aIIdz
ywlUk6vDo+MvudA71bB68gLAbE9Un2GhVvGDqQ5MuwLGrirWtyKCOthauC9bZaSjLjOJKQoMBN2Q
RfhqNT6DoDalYT6odSiBVUlS3hmWaDRzQt9H3Pud4EHMnyOLSUJGIZnlILJip/kFl5T8BRwhfrjL
pfMcmM7nT2idbH9ty4xcHRVFd/XpcPQt3k+1REVrtM06bU73qRYExVUd2QehiR/8xDG0n6vOt0XT
Ty9xiUDIEOGUvQ1s/MdWSmAq3vtgqhFFp2CO49eeOcZuQUtIJWbjEy6yKevafK5W/AJ9ltqcQ8In
XH8C6AJgEsQK8DwEW6p3xMfNxtYe62+ny1KGkP+64Wp/jWFJryKyfsstppM2WaI8QYvj9QiTSuFS
WinyqvGZFU3UPgNKw0C6FIDZHtklFFZXqjS3GtD3ueO1mEwj08M740pOiB8XFosr6hlz38eLcNjt
0naGIo+5s2MpvTk7c4kNFEdmdplECUjjTrp2Y1ZyTSbY99mt5Jhaa1GO3aO6ZU5K0ssq6mytfwWd
H4s2bCuRJ57u1qKTh2VUhofppAi8Tx61j+eXFGMTwKA7P5wf87QIkHRB1aTiJZjOx5h1mlrX6NJn
AfL1pWz9Vwxz+iBwfZrdaA/WWrw3sDOr9sOpbjnf7L7uTdahrOqAn+9aPX8G7jYIlxvCVS0cMNNx
bHLz0oubE5MNsa9ppQY/JgYXS65tyhZSoriNLGRWq18cNWtJ6qfgXyiIyn8+DeHlMQo90RgBTJ0i
xyq2uZVpC29ahnwQ+9lsiKioaLgY7VLbQGFEB3h6XEHDzAM6G2ywubhXlZCwRoBzGimgFxEQJSUB
di7QlbqtxUPtmEB64s/lW9eNmlZQHLlY9bJ7W8zkpKRQwOGc8FcxFdwTvgjnZKmPWhfyi1OumtKU
rjv/MEfAL68KlIyze7K9aOe1T9YU9gE4uT/8t7MttPwPaFcQo0qtqD/Iqc77uuw/3FdhbsvOyOzS
L+UtBDpp5U7Ov2uwFQgQP0bEnBFnI7Tpeme9FtLX8vQFOwWY7kz88WuIOaoFw9kiHTRaCQSgi06k
KP8LtggtDFBVpzY6ABUWz0WsccoITrLwc3ZXE6cVuEl0fouImAqX3lxA38fh2jOYCE+/gzKpA1Sf
hyMqUstrQ3KNTcv8YJNIblWahRSLoLhtGmxPtBsGd3lA6sUcPeeciZSMBFTABSwrhmoHnIpXaV20
ITxlJ+evus3PJzI9k2T9zB5gTsH26HOjoYCOdjgpjuQWRs+wWoX6yGZ9gpNTMSj8X2LoCPWBYTqx
S1tBPOxDTOVTL06LCndWWmnwhsYRZUL+ygc4RUI2t2W34jmpIA92j28v6hZ2RRU474D3Ge5qd9r5
LYAK5n1sNsrgimcckFdVapJQq5DxFgsitRlQkkRyxgn9h8GT4j9FYNweuOf/ayA5W+O68Mn8vvnA
OV3048Ng+4pvc8x+U4fuaL86lzjIco+uWduLpA434O0iKRnx+B2bOVttznYNygq5391zVX25PpTk
z8uZz/0XXmhaiwmA45UErs2uzL0nPBe9K4iBudvn9i7lwC2RyZ+MUOEj9SHGngrGgTDPlXj/y2rr
6/zR+0xLAxthiFjxIeAwQibWM95+gVuwFiCTL3r0DwX3f/tQVm8Bc7mey/NIOolVrJ9BkZjrfnkB
jHVUdoVmypaD5rpKfIt3NvmiaOrrapjHwIkwxfpsIYmfz6j+ugS/2AOlw1DpxsbtgnBhGR6wnWOP
Q60nPOX5mwoS8fwbEwhRTh5/9d46erYK4DBdO8VSaaDyOSxdO2qhLGR0yasY6vJJoxnBLRDANQPl
kKAvx/zN4a8FFDNU4kPDoC3GBycxCTKTbvGOH2GJIe+DonsDSpwPYThYoUvnbxIun5pfwfu7bvhD
wt6rBDesl0svYBeb2KhY4138hBEln9mwshdzZqMdq4MD5/Pd7nDPduZWNv63Y/rZ8smZsEUp0R5z
W5ErLg6mU4cVVrIj3L+8FHIYkPwQ5LqNcKOfeFIyCZYICyeLrPvIsFNjl5dENs66XDLOTXy74EFm
U22pFAK+2aptdRanjcwDhBnVA3gzIQjnpce2i1xV/Nq9I5OJ3ocP0tq5DJog8b5MJfWYUS8aUt4E
hBVL39+OHbyMIxEHjuu/miO3T/Lxo9XENOtxy7g+n3lOKZ4R4jPulSFjyxq/SvJtnZv0ScQDNhMu
fndcvqfB3cMb1PgjHHNOzotBSA/PjmGMBP10JhJVFWYJnagjLkQLDLDtLsigW6QHtCGK8Lr5vmxQ
0OseEj5ZSTBoeTzlmIroj7x9cEddeqOAMtyabbbyr5cpRsJW4ce/ftDzgkXHAJZVQgSc3ne/tNbs
LYLqChcdtm9V0EXLPW3IaUokYdl2UGJthy1QLevEirQnRij5QMK7F0ZtVrNBYuL3VBrC6YObNxOr
w2GZbHJoAMoptJiJ8iF3abtqVwVsoznqa1Ut7/yUH1dJb7q02UodlXYPV3Wc4zRvW0CWF3vlEK8j
ZF9gk2fp8xh4VGdqt/IR1zaV4G/y8a+ppooTxu1WLHDgZN4VWCSaIAHP8tBXR0nHmTCZJ2zfCc6C
vj9FAoFcopiPXd+VmIVA6X9X/nKXKm3v20s+phgRzsBZH/i553PHNAcOffq5BM4pm5hMaz5bGDI8
AVqPJBRY/fn+roAC9nKbELr+tEfyoKrLPzBI7H8ufzgy/PrlX8om5hSza1awHwo5mQeDfnWZh9hD
WI62vmhgzeTFGlPZX5h20HrK5/YUXzxgEdr3KmgncCxv9TUsmxOZTgErvz0omwWSnZQggnSYAUwD
Ickwe5oselWAszRQh3rrHtdjcUpuumf7kJm5UU9Rok0V+BNOpnwpLmhxWAxt1D3Ci3lV77u4DhTS
iv6425eosL4Jmjwrfowb36ilnR2rRy4oSqXH5lvWpfKUgVIXxFdngUs4pLRUqwxf6xcwj+49G5bK
WBA8KnGlDUj6Z+n75psKwJUlGCrrWScEl/M8KagdOjhMxbmB2nYTuRazvaxYfE9Wx4/Ycmu2k90w
l/NqtoIMj3cvUGmn0LIv4LfS3Cpw3qZRpLNL134Dmvux7I+/Ktuym1g4BWCkCq6WuJ4AwhJkSqYV
JU0VaqL15naX7ly0khU3x8x3n/xuSBj2Go3mrPOh2ogVU6a0YquojH0VC8UPJ/Eu5k293ksLUJBv
9oXlrQtSlZ5YgnkCwiqas7UOSDbdqAkNI0WE/zy/A2UxY+ky1AMd6taWgOrrYr2focc0SFnw0x20
0flOYyA15lx4wmvTlg59who+sL0njG0XJY/wbmuDufOl2hcn/Pr7O1z0fuU76DyxGTBOJDsYFd+n
ggzH+g+zEqppO0ki7Y2mmO8inJ086cMSSxZKfd6ZxfY18sGTXm3Up3lx3P/hn4dly8ADNDPhIrXt
Ly9dA8Mp0mQPLqYDJfpAMUtchnrj9UaxMmHO+QUXuMXnnlpZPcF3JjU1oad3+yctEJ8gs4pvbhL3
UZ1ttrbcbLKMqO1kYs9NDJ7g3o3oZRHzhcw54HRlgTj8E+XNgSZfWrrf7zN883QfDIY77W1rORYT
GvgBteEjMK/wW8zv9SpBVwkP+Ko4eLQKeoBeN38I3Szr+89NzMjolVGbadHsqi0CVI2/uMy7dn8R
mbRv8hq3a5elNJaYDIQNvNanh1injbgQndnmuoGsbIJvJTFAQKRG/EMaHk4dsG0w/UfI1ZzY/myJ
j0YdA84bfYXNUS6fXo8pJYSgUCQivaF1sG2dXGE58EniMaYHgWrASaEzaQX9YVokGDVrk4Ms+5H8
fCItiQiyMeUKDvDER6YkNs5HKtK9mW8rckYl359VdYumcs+kYnH5RlHCFwUp9zX9tjJiqKYH1urP
lRPj8TeINBuDfx6T/L0pDOwnD994fi2kQHB4mcMOhTHCilDHoLISGyv2bnwnk/idspjcmLFRFuZ/
FWV2thqyHOMGy2qISvKu32itAoTYQO4JXjo0J35p3AmTi5A20YiKhLGcIoMJEhcFQ9Ys3y6rc6r2
8iNC6METTUWpa2hq8TezeBvWlfvkbS8FovsBeTMqfnHsrZLpL+AAHLarT9tll1OAIwQxtXsrpH/c
h7XhbFNAeeznVVxMSYKnh3GQuxf51+djwji5+F5N/CLmrdx150lzmHhY49yMbC0k+biduTppo4fH
nleZXUqqPXlNNp3vIXe68LpTDGsbdvNhkZXpCafF1WzFFvYWptOBlPV2rNeJBMfeov3MkUTl6MaB
QzhBkjijYQDVZpw7znBs0wIDmlvd4Ah33fJJ3ADr+BQOuVOPYENCp1vgqBAWCEdcCpFgw10AQM8Q
NEoI/S1+xhEMZJyBIqhsmKcm76udvvQyz9GbaWKRI5DwAZoeeW9VWP2yauY2SHj1b6Y3ls6K6XsK
47das1HHIg57nYImC/rBqSxm45O+tW/UJIy6C5gx1dYYuq7dMxSNCIjQbKfmvp5lFo7SBqnvqNhP
1+CryGrPHFbL/UGOoYkLUNvZjWla7YtCvj2996ndhSP0TTya9Pr1OtxkFn3QN32rr5xJQGMoi3aC
uyLkqEcSWqfV4HB6yu18/IEUsctckm+kRHL/V6qX6iSW/azSeVtqKBmA8dHWXma/2K4oUERHiuJh
Xewb5gtDWAj/Rsn7UB95+JyCg5ZHenzj0HwwAlR2zlK6tdEcMB/5Fu0RagKDUzZ6LLiEqbUwEE/n
YE6lLbfEIEfWWWPtU2yj3eonIYWYkwsSYZnqXeC8jAymoD/XwlQqcNFldZQLE7eGqVEz/I2z30no
lVdt6yPlbXJn2QjbXK02HB1w8ZYd2XpQDGSsSoZwtjpIBHgU54g6RR56QQddM1mWX6HwrsMycimI
89NwrJRGUo+p6HC1t3Sr57eA5IdqR8lR5sXGZOb2ilLXuFBPDskEtz9X9km1HjAM3lvY/MaVcC31
Ca5/V+mi+1ft3kO6NjM5fP9giO03DaRDgRIBLBPIgQZNYDnp5JTo0YNwWlSTR9HtXDZHj8r1fBSA
u4PEGctNNbQuFeXfG8AMhWoLavlydVzBUyMoWjvJWdI5dXZe5sdUbT1dbZwo6o1hMLP2jiVxEEpk
PfCOAwiCwFaCpJaxN/y/jupVvj8xLDzrGWPEvdAohfMl/L7PkaFpgOoF8nOY8w5779FJyODPLFdU
Umew/v6bHE15OFC56r3ol2GR9jWu52pVOD0OkucRkIxiNe3w+prwbEoXqp2K8p4V6b2brKqM1McK
qrShFnx93w97N50K+NiZgdhXeasYVwqQDCTx+79jGaTwvVhuHsnERpmHbbeHIDhZ6Stq852VaCFp
MyT8p3aj4Vk8LN3lpV1A2azj+VNJ2JDHc4Le5/4n+5bO/R2ME7l1ZlehNDyHcVNMr+PXAuO0m4/i
xMih38zTeln3a16yGGszNkqR6+6LZLIO3lgO4QlG18IInhNnxEPK2K5R7XbzoAvt4WHD4trmNI3m
khwoX7Oa3LhBJN2cFc08bsgXr8ECOeIrIbP6Hs5sjZVg50tuNXzRdLZ0P3QPr69dNS/kAmzhubGR
5KpbsPRAhaLILvMqMLC7swBT78V5+7iFgNwNvl/9II88V5NeLRQgLQ/L9hrxHb1FqUUB0dHKmOu7
Nyxnr5TythX/3sOwwwaxcPjks2CpdBPvsP/1WRBWMx7y1yckaMFDdvXu54fNxgNAb+/gmLS58/Az
KurCFn5vL78GvNesNlrP7UylGb/XuffW1cOl9eYgCltDORfXDNSFEZGLBoqPaL4qy7XpxV+HhiYe
XOH2nv75pFujspGnR4Q82LN9vS0TScuvOXeh8gcA+mpfTOsaBDlXwluVKU6Ljw8H49oMc2L2o2Cj
kwfECW3VayrDqkEZuMrMl42JSgbj39TBmHcmeQvogNKC0xsHDIv9/1Rl+cMMVcbZv6B8LiZmbrih
8ixTPR9HBo2VfpJJMfxeyr7xoqESpdpNTDOzmkO5UKn03j8jHz58RqBNWLSSFDPW0ecqBc9AFgcZ
hlnZcWY1JS1uZ7LgPC+DSCSokso5grw/J/qdxgEaRfKNoEmidN1xrGiQlyRuwPEIHYCv7TLEE5kp
j8PU1EshSwTwXFrGoCwhQ76Ak35N6sO2EwVAAnh3ePBLAOqi4T3qqMRbzQMbkUtx4iVneEj9KLCo
lNoU2ffN1Ww27wxgtDs/greePBDnHeVxi07kPzSxmqpvzeshkzTZHsO5WzzudeXa64DAodITK7t7
TUO5QHyHCYn2Fm0kgX5oMQb2Z2MRN6su1qT3kekElF5xaeV0+iFfwy4B6jRG3XfMOas4UfT/FrSH
cSSmL5B0pUORORhcVjOB6M53XIRIoL4oSGtld74Q42ipGMogvlXWH9N7KEPWehwbqI5z6YNykEOX
rXHMifTMC7biy7+ntVVXiG8ZT+WOm+uZFmyTk1M0SR8tvinrsN0SJFERVM4oII/D3asd+UcdiFDw
STnQ0prXvSoktHPnH9rmQJ2k9RGx8NpjxqF3ojZaH8GFHFUAYhgy1LiORntHhs5tHU/BtseBaNit
+y8X7hoqTBHzYEj1asi0wcaufuZQg8aaK54BccPdOn/VzWAqTxzF6+QkC4PvR5vveWatKcExC2q0
Y8Bv/XoMHilUexz/SwnbGCVhoABYIznuoOplthVkRp2eY2NyjoeN8P7OBXG33oT0f120yBWfnhJ7
myZowyvWXcXFdB1NYHNJdw0vWvlO/yJRt5jTtJWvdVHrkq/46vp8ykL6mddoVEa1O6z0DApg2yfK
5cXRLKDiPpY9nFrOXdwBY2le2KTn4tU356Bu/bANXryXiDlGmtg/O5d+/k0Xm+wPVwFueHc7IfJ7
SdeU3JOY5cqEn7QKP8Hn/fwZsPnZhpHiA5ne3DxNeOTiY0x1V/PMysrzjkQSkrXhTn23DlH3D68V
ySEBOTcz3XHapwaiJEgRnJjSR4/+8jMtaMd8ki2JDPrhq0KPjYAzYmaw1c7J7SPfUQOIct3PR3GB
PrZP+bxzJ5aIFA0H5N41MKhJnCqtoa/cVkJ48gcSaTBtMO3QRkjZtbZMIs1pq91rHnDKWarANu9e
+rF6iPyrfJF2XF48E7k60r22LWO/1nYqv6Xk/bWhRfuKEthuHEqbqzZVTYOKoLl6+D4UnFIi1Q/5
6tw8AMg/pLkaBiuHa9wkLEzMcf1yNhFVPin9LHMZF1I4iSOEpCo6kpzNtCG+CTApKTAFLSrny/Cj
Flc2jIDuOdzoGHtCWma3NtckpqyNr+Z/Qt0KJ9aimp2jcEMelVKu6PM7Jc+wyu7gY7KOSbDikco5
g1/F2b2LKxFvaATycxvn2xh7ojISK6W4tVHviIkJIU6Pl8bfZHmM00ljyIJXSZR6Xj9oYcm0lJcN
oRM4c6iaAsg7eoPmpgURPhUVA9T5pl4tqNLiLIsmKnM1Qq2F/kox9Dq5f6lr9gcR9b1Sfs4v3GFe
+POHFktVZz3kFEdU2iZsHSq8uqu/Kl64OgVUYA53FPDRcyt2+lPEPC960ND6XqfWDn/bcwTmDd6Y
XPTiNjFLVZj3PBZ26K3nBBCw+ov8SxmiasVtfCLTQsYV5mb5VWDJoyiu2Md5UgF8wId6j5kJ4Yl0
E4YlY6rAGZ8x7+vRKgnILuvt0ToQ6txkx5gKKUa/ypLF9UF7MzegAAISkuZFbOOvwJejZnsun0iP
qOZI4xlofhOoqToOA6MyBBHYkSaC9mqJApAC0LQj36Y/4pUXVo2ijgkWnmlYJB1T8QhUK2bvkJeb
7NoyRsPgtK2Z1UEaq/Mf+OkAM+G+MaILBigU0H9ZellZEqcNnhNgeY/D5RKYtB8pqwH3gJn2FMww
qXaR7n6HYtL8dJwo/e6n89mO242Ez4oMfUjgREJJidCqKgWuxMGlOlsJEH+O5b3resoU+ZMFN8u7
oB8R4SLzmbrJSgcavjNkPUMFCR8K0OBSmcJ2IsK2puYcnfzaCetJ+ZEPOKq5Kf08+NKzkf78qrjX
wpeGlOMxjqENjj6PMo/RHOd34WQQ2pFPEAKIcj4LP6LkO/xiqCwp5Es2pW3EGzNaG6PJ81tDb0mK
KTS2wXGfWxHEFYgpCMM/KD6YrC/yNNlzuyVvi3C7BDSlHrUfFgr+7K6Ts15I57m31o9K7sOsfRda
Q1V3XJyjbQTDEH4hK08oYF89UHHMy1ew8UwSPdxnhqgucKqkKvHFYg0qDtIIS6LoMvOOPMmrT7pL
f9FUa4LX5y7EqJcIgDnoURbdH4aEbb5dgvELbjFIZEa7yhNvjt1nAniclKJ0jgg3tcbbnVA+jXEW
4neInyOjTyYHjK3HL/D6bJa3386qZD3C0C9RSU7osv0rLvzl0Ii/nzuMqwbFrfPm980HLDAC/aIU
2OQ0iJWzdzv/fkGw2azkDfAkHzZRTM5uHhqghCCdOk1jlESD8XQFff0xv1jK62l8rJyAzRvlDkEg
2XyfZtAQvMcuWUXjsSOrfkcJ+rBaIj6x/57Gv7O16CsxeHre/t3VUXgY8LdHKXGM7PfTu7ysNFU7
3NJwRzgGTYUt2ojs2QXdumgCTzMoJl7KvClmKjzI5HwXW4c9NlqnYbcBA3FUdAknA31r3pIpo5YE
vdmAV3rvQrVQzkSYM7Zd8YnDO+U1o+v3B+fiE1OEFsPRsFS7mlGtAwaSiCqGT93YUME1ux79UGK+
90+XupPMwWT/1N21eAnffdpbMCZqF4kgpqJIKc5XPYlNQKsjKpxkpQibRwsZeiBHegrWOF2yw7rq
kZFUnOO7z9pVUA11Fn1GhRrnvtyR6wN6FhClbXjhzkaZ+dmVqtG25e/BEIWsNaHdxKQdDkigxcsS
r8GggC7s+vith1kxb6STFzfJbd7DNf8AIiaBJp6FQMmK5sihQWnNi2nQnAQePm+jPZ6rENOSKLXq
foMZ3QEBodbv8wJ38x5PXMoqGciHYPSVkH//XWnsuNcbs0vf5hEnJ/nJkY3VgeMDJ4tflxEs/uC0
9XVCcA3VxyadZH7Sh7RPv6Y/LLBlgaoVdZbmtsplYaXtqpOkcr/MGimUZCFZGilpuFcPLd1xip4N
osVnf8FHDjD0Lyx9fjvNzjkiAGCyPA5Wp01WDCZ71Jz2Md1iMnkUhDgSfnbPsb5J0m5TYPZWHw5/
GTwQggy8c2K3ruhEXbIHRpZ6lI6JE7k8IuRGIPuIhx8Ltv1DJ0N3nZMMPViOcdfImmBzNOA7W5v4
W8+4DNnzqFRaaZb8XH0/EtVdoTvHCC0joQaVm9b/OeRiI1+xJ0+bTSLXr2/NySV6Yj+p51KCVrq2
14smqfFj4WIiMLNFVpPG8v0qLr327PxeFR6U3gBcgO/kC4tP7tuXhWuFpPiMeUBSYc4E/W2kf8gS
epNSpD1srWyJknIaPvLgIa+Lb3Kmo1q0XgXCWkQNUEt5fm6xmAzahy9pNptMNEKKYihQ59KT9+vm
JTS4fb85qwiKq4JY5/k2/7ZZkMfZ7mWvoIOlxq1IZlIhhIqnvIcD3E5GbYe56iVHT9RqlWIhovQJ
QFYx256SulnkKNGNVuxSLsAcFbKY/55WyT4tppWLweMaiAMqeVLQZ+bI+BIAwOKMPyW3Zpqhqc7X
cLx+CbgsSf0GUXqUY9Gq7Cg/VpLAhZd+Z2I3EPFWJA4FbowdMoKbGRxLmxKyINptYRWDXk19H3vK
NuBnXKH5w0b7FX8jsCrvmVOcnIA7rv69bZhBA1PcTBqil8t1MfD76qKXrvyaP98ifnxEjFbbQWOc
BJcEVdkTxwNKLv9wWT3vEJvcyLgn7XTL6Z7w1V5uJjUVPVuzXmewbbhj2oor0XCG4K0PQKExuyMW
OoRBpcgTIWa2+t4yMjBI/WTIPw41WXKQyJY6iX2w5KHECtJSprLc5argdJ8qCvgIeZLIB9PvP1lD
zhffmBh7osAZHMrhqMZsZdLKdm1klTaM1Hov75+ZSd3w+88cjHTJq7ZaqBMQ8/iIrtjRe0i1Uvw7
RCQoKMDpH1dajKJmXPd69CcGJClBgK1S4funSrM7vA8CHgel5mkLQY8HY2AW6VRxlMxAZz0PqW20
Kqaz+M16MP22wixu5XFvrx8gA6jRigSuBu8gEdei5b5xtMLIxtrXEx7OwJXq1OSyBpoIrWYKg9LS
cqt5H8187hZ7W2MT8L6JBnToCq7QazPoFju+RnOCeDSAi2nNR57KOywxJm/ig0q7+ZPLD5Wj4hZE
AIYkDloTi29+bafFEBeCtsLq34Ypy1kvElvysGaft6jkxoYlFQRcrtt8hABj3AM1SDJKpCL3ZbqZ
6yy/X60hTBXWmsp9iABoIijP5AaD0IWK6xkZnvXEkbQHEt+rxoH6fgFyM6OIRNYofVgvYKUe9MjS
/XXKHnw5sNU9Qe/GRnJQiTUfAFw2aoX73qjsneZ3buxFOULK0UJHeIE91Iad3ocJmLWhMl1Zvlz7
tL65uQgsMrppa4oJdYCkk2VDjZoy7Oii4leodp8u6Ol4QlDZGQy8fk1Y4Mdn1rJGlNuKv+SQKiuf
LGsGU7gMHJAGYSeVCVDs8tTQe1+fUtu3Iq78ic2+zeUWFM53KFSJGfdvHigaVLWjnAiwJaDXxTvb
GDwE+VTsqPON3hNEVGWe5Pr4wHtakIjfdDIB/51blzh9ZHJDK1aNS3m5vlGsL/FQ6ryPfQg1zgyW
1DdJQRkksEYFOYIfW5zuComRzqnuwCB8HaGk+1+rtN0Mnvd6PSE9lNKH+TZQL0siWCOz25205490
J6JUlOJtw3619Zbb4rXTHkpDnQWNe4zAQeQ+/CHlAQUS3iDgghGwRmOveyD8tjVwBukXj2sdqLco
WMqg7N8R6HG0heYYvFc+tGQvC8V6OisWlRrhqVwUyGvwZ+SraJm3TzHWrkcMSoYF5ASg8OQhMlGZ
G9Xq39j4O12dDHYT6B27LW9JVsK9MpUEgzqiWWgttYYMt82CRli6JIfBUTf3iGibw6ScHYY1PyBK
nQsbdI/Dn93wQ7YJhPVieODzQpW9WJDx9KOunETJBC2dMqbFa60vKiq4LuPioKM4/TAHsP5BDIwp
vZ/DEbEeFqQ+7aeZ5Rds1k3fekfqDrASHspiVV7O70IccMGo1rxmtxLwFxm94ZOOv5WWdkoCvInj
02RabUvm2QJyiuZVwN9oZlI3sndePXUP57sdNT9dI9DgmH4idnbmRcnBqontQiZbl8Qr5+Ja5cXY
vgRmYJ6lXgW0fF2nQuuuQ0nNffRIrHMFT6+12KNxift4aAeUSDnkJBNra4kVKn76DZ4PVntZehEU
a8cWQDv+Lh8bbpKAXkz4VPLuh4ZTF8JEifRJptim0ZB+1Vqutgz0cYhN6ExTFx2oyGKKYNeB95MP
7bv8ro34v6nj81vZH0GzcTjjNKr1LRlv38BXYpCA6O5RHUOSmpdLpfAwqpNytkAHNSo0bISE73lF
tqdwY3SC95l99rLW0aAsPsVbpuh/maUX2qPc9WgHcTvJTAv6VnRQ8iArP9lg9RKs7S5KF+1JUG4i
e+FlDAGryLMkumxDnBjmWTLbJehiO6OveTymbHUWU6rx+6dZcbp6Lmz1DolFrh60Uk+G+/atHKCI
XB7yb9B1SEn8+cQJonkrc/gTsUkwbGfbeMF17E4Vr4xNk17HRgsTxmPbNbs49amP87rDBRjpPEp4
gg8x+Odh7jy9oaRlOeqjaUQaJTyIULLLWxlYrQW7PJJXB5drNB+6UlA4cbZOjqqmyWUEhhSgt7J9
3xT7xhx7W993tL7lhBV0VXPBFp2/Q6Welz9CEEXhlXfzZsPD9bzN5hrohAHB1H13CpmJRi7mgrmE
MuiCxZ/k+sDW7O7I+3ZVsJ0EIhuuwCzAeHE/D3vcEBtfgBzJPsGL5zwqEG86wCCeMXBeQAIpGBqp
CZaSMBi5N04lp7RT45GqD4iac+SsCcfXhERuYWpLcU0x2Aq+gJWJ8/6pWVYvJt5u8DC6OeBjg9VK
/IOJ4kmFGN/SXnUagjOT27IkohPYdQ00SEuFjC1RlkufP9ssttkot14NivqqRzzItVznXekYT7wq
o8y/ihEJUz+NjSeRHxXdOBy2Gukc2MXcslBpjPQhqWTzUWMILg7/D4eqfjQFZb3n6DjzlC3L3K/Q
ioTQPjcIa32f1yVECd4wZeusc1pQdZf6s/pzY6jJu9SjC+pAFZvRPl6ULh9XCVlsf14tZ10Ws7Bi
RexeffgqghI917xWttnYImf0zHSEICcQ8FMGwZCWZre9Hb/994Yw1jcPIPS9247Z0kdn846HNulr
W86wLVJRtIYUJ6UBN7Mamo/Y9rUiW2DQ2L2nvr9km3NIJoBHTJUfLGxGP+eU76pN9yegJes3wV4j
y7qKgeQNUAUfHXDA9KYv92gNak74AoD6HiPnK6b4/ocFegFkLXDoh0M0ThdviKiLStbhoR79qtKq
85DEsNFsk+nHUBvMiHxPTgR9q8McGX31T4cGqHkVVVHj6FppeaC5yDEY0O8CPzIErxSpPAs3SOaT
XkYPcNO6d7z2tyk3RHqWplOVRFA7ACt2F+pkrIGc0EK0+StrQO9W2NS9u6eb+nK0q8eBBozKpbLE
dmfFaydde4zjohKt/7tOECfSohC+kZebfK9rmhWt/7mIMnVm6Ij0Cuq6Sso3Ggrkm/55gfr5T8bP
eznGHhaDL+gFVmOrDJ0jj9uwyKH1B7taNX7VyHOWT9fg3hz/3NouB8Gs+Pou//8kYqupAU/bZQTM
PPX0PvWQKLK/KRDKIh5F/qcbdHkzZxAg+KIuJDH5QZmnZOM3WBF2qnVZzbR8x23kUIVa36ENfsk4
QgGw01Mi2Kps/GkZAbRJYCdJf9KuV3O60TlpdzgsRGjShpcaQ3Fl2ypR84dTcCNdD2VJlBP0XIY2
x50ZbgyWEXQE1ClNiWpVHrjRRFAt7ne1PALhjUIshqNRsziUk6h5Rv/pGO2ELaxETu4gs/nKJqEm
sYSAYmJLSR1cVeaVwU9H4uBLCwuFzsmh6NePVP2xqArJfsFD2RFUD1mwDSAZ743s9ba8PhjFWORy
YdwNCdOsHjmWZAmzeaOaKbDvKfHbzFqGNFNbLicIX8XhwfwPZI15kSDvKV/qM0XPYSYYe3iE0mPR
GjxEoqZHMJYMNYIKVuAQId/e4YVrWmDPeywhWFnT6HLeEcFN1e+RX3j+QkH4fgnMyLJv7nGvH00b
N5SvTl1VN7DGPx8CnhYB4rSyjhM5SKdFhH5bQr7o5O4mYWjLbinMR5IE/tnGGBNFD/BbWwsZnAdW
VWqv053nXogVH186sv5im7KDje1RXqxaXgKRw5sUUMKnPXgTJZWUekjRVb3BYw+C5XzodlOMRmXJ
SAYs/NQoEdCT21q4JfsLjPqufnU80s7HHgIuo4aaDtXLBN0wyHsmLUYLtNHUZEtG66FIS1YgTwiM
mSdGdgruXwx29VjyCb3RBiHlhhw06gzYuAPZoi5z+o78DCBqGCCSy2lDL7OMCWQhAhZi7lfojo20
dawNJot5V9B+L/2Vx4OtqrjIbjmIz4Tn3Je76IYYFoEK5QaR/Lv6PqcRg7MPbRgZgP/p6NgAb1gK
dwOItTGlpnMUCair3tBz0C2A8EutjL0hMNbn+n4Dv5jPTK9oP43LWwvhYYKTcUGiLdeuMh7L//Dl
omjK7WTg4WeuSX2nv5gBSisVAnXbKRD0VpSHY45QDFNAacjM71VPxWt+ByZVxtAVBdXNluwz7mI2
Bt2XKRDCLX5a96uvpQedFcpgAacLPegkSta/o30Ff/AyD+I8QBsFXxlKru47CRXcO/YIG25CZ8Vx
ZRGO1+4uAuWmH9tJLkjdxZLh6TGzFbaQ+yz+Bw1hzb55wMMGLXXXbSHKzDopt/dzWLmzmAgJ3HHk
sgrPthPD82qrlzRVSDIu4GEWLYb+7+yIjQR6fSKtR2PPxkxFm6XWeiWHqBxxLF77Zl0BFjMFhnA7
+Tpfjj0T/oJr8YFfv4RFeStgy7z6eF2yNXUUxRQ+jQe5uF/Lslcu3QDmrj6nBnzyR4MuqMmH2XCQ
2Y4SVxJYhf7syK0Nd/cHkr1bNoCNGhsw3Ztwkmj2zVvKvTEEkUCB8MivXH+i3zHi8b/mKNEUg93k
NyT9q55O4CiXzQkKEOgw8imawbfAxkRECs4rO9K5e7kIK38jAkx9QsxahI0Z1Af6Ts4yAb27rZ1t
roYu10a9d6H9dNY7MwoVx7mfGSJPqXtR4CBs5y4KpdhpPz4KJxXaWHbtYXeuzyErELP/bzR3xiv+
HbbLBDvOKYa3bU21H02wcJbAMmj9qDquz8Gj618dbp2ocGr16fnKZBTcLR9IV4F4bfYQJKNDQZ4h
fHa0JzC4Qi6bv+MMs1SkqzIKofUZf3qrVNijRU864Efzjw6BwU59LjSbdqTVzzjZ3pX0nLqAVrha
nD38hMCXZjp8WFl3tHbPsw9T+fWltC3wvhJjyQjWs5cgNGGhHsDhSZuXVRXN2MRrRek96Lbr2Y5o
HjZfkblsv6rqHagiAyRPwpN0uiNr1d1gBIBAjGOWfTeLkOGts8QOfsVSBfas5jrKMhzTfocMzhmc
WeG81WpdU0KLE1LerOfzJOZXhLZtaFuogT3NuUl6yqxKxorB/xoZeLb14ufLs6rObi9npYK1+JfF
kHIfIRdLUeyeTzMGu2HblyIqlzVwg6M6/7AH//YPrut24m3is2rYiaHmISpR8l1Z8iAzjWDNuyyU
Mvn4o5JNMlwtk6QbjGfUxnnulVVtuyi3ngf6vsCeyyqqAze9o6S1qNa0Z775G1BsHyLeHlBPKPUy
f1/qikMQ2LjfixReyW5xWKHojLcAlRKGL5Kc1+w6c2W6v1pySd/x9xT8uiQ2O8G98Zci2DHdZuMy
4BV3ZhgJiyDbbWB0cbmK8IR56nkAHFXeyJw3ivSd2fLkdQeKFodw5iKzHk9CMv0Kku4WgGTwGY0S
W7k2cTCyWSu3rVLtFREyZor5w/laU7Y5wQVNlm9EaGK4eM4EefvoflRU+DWmjxK8o59//fD4uYWk
KWNCowBgMrEhr08rVOYzDgkNkjYkYu6LV8YwTB4G3amWsk2NFrHmSOvSp1GxDxk1Db4YSF4D7jdA
xm7vNLsA8ojEH5jq0RZ9TpEJ+k8OqyY/v13eUcubJ9RYA/1xWcbtqS4p9uDXAEwf0QehNOzmw1X9
qWJul0QgFDO9WxXylDwxFvP2dGJOQPymyZpXV9/8UOcqdaxX7i1OsvsmgLk7Vaj+sLcSUjRncivQ
VFaWcuAueHk9y76bI0bkigca6dPpD1Z3qPpDhy9emsZXvqXBB052b10C4efJWN5xCQzeAgM27IR2
9pfdVAB02+mkJL8S6eAg/0q5uMEAtDNACXmudlvopgDH8hhTrAkiKPi7G6lrRIWa/EfL26/+EHs1
ynDewibmOcZoy2YPQdOZNXjFlGRNTT0qQMao5HETz8daoJBdRYG51bEdoTv9yo7cvMqsoTA81j8J
XMQdvvfqKeT/ySQlGaDQoc+Qp9sovw+WrprvSQLRMi7LJDlpL2mBmz3eGuJbn197XmvPSm5dZcXh
++1P47Yq5EFtJK+Z4nTPuJCI6rYqTCD+CNY2XQUHEFpfbFo55mqYHtEcA0O/mJ8HnZ9s7MQl1Vi2
LeWEBYkponpETAOc7O4RropUask/sIsqJYMvYXrFL7rIVVCu1ORiV8sTppJFe193gjkHYjemLpif
3Y/EklzTanE+A4Wo3SAy9JgPFmRWlZ3GA/8XbCS27qvz3unrN0f55e/80TMv3CqtCTVVZjnsIzTL
pcK6AZ6SFu8+V5FZP+FM1TAl+deaoE2bfKMwA9YfsirX9Qgu+rXEqAYNo8IgHedbXFILTD3W29p2
BUcbGRukYnp7g7fwrv/GuwQlvY2d3FNSsIH//ShhbRgPa4GrtRIy3gcsWPg2Pk0oX7TzxvxECGhS
dJ8XVoXLHKeN5+DviIzk+CFKqifPjw7AgVgf2Z7OmPe/J0IYwfgp9PxW8H9IlxxTZQMac7B/ljOH
Sc/TJbPUsd42pmh1/HSRYKqGNvDWj7JqEeOvfGODWKSzNa1IFjCprsntfNEPdZxa+C14d8K3uKIM
CDS81FoHlmafBxSEyO5ulpq9npVvHq5wMJFVmwiI9uuxwFJ49TEW7kqsfgTWeWOw0nfmWN54HUrJ
k4xnhVyDRUewAXiYDCMAtOSKKo+jdXulDqwSNUTg6W3EGWUq5HUtrB95EyHuuykJmGXJDNK+469I
GfH4osodFVO5yRcigT5GxFy7cIwyyh0B3uM2b5CS8OUmKKWljtzAL1gMPMtCn1A3ZvbxZzuKBuLd
667wY7MZ+ZPJaMctwdVCIa4RzWYDL0Df342xePW7Wh3zoqK3akhypGvoz4+eFyAsAnIO1HbPaOt7
t+V9Qa0QL/82npVl/BQ0ZVlt2+BfwupK3+LF3J/JDxi99XJ2ZU4y5mtcyAeL2DGHdBGoCIiMUMh6
+R7guMJbCZw9H/wNIT8MhafkFgMhE7mrid97CvCyo7yGf5X9Pgaci3KXod+KXlts+hNbmzp+MoB8
1esaGvHVxkUvIJRbkLCXgjyyWx976iAywIOrQq/2LY1st4FN70p2lHlf6ZT4SEhnKkSCtIYYmta2
9mwY8D7NJHc6eLWi01bjqZ9hTVkz88lfEs9jUCc0XLZbNZt9cn4LwmIQ3BISDBM+xe0/E6Ax7rF+
k3Uy9DpPtB15njBXEiRpQkue+M4HyFaTqf+9mcfikLysgJVu0+B3TsQHFs6pN7VXywJj6zFWufeo
BuXJZcURZ5WpcbIkhAKTsrGVlnLdWxiH5Gd3UggW6MBEUu9LSzqIsKhcPDvWvtwXXWVpJRRbRxqR
o/IDd5tFVGMajTZESfEpEW73ngVImaL/kmJTSRB6ejCTpI3byAUNCuztDTyLPK1fNq+Bzzd956d2
yay47d1xRgspGwSkWzhWG/hiToODWMDNnw4GlNiXN0X1uuS+gU7ota/A29R6BHHNVMlDHCIHNYuV
5aAs5TUSgK1gevDDo7jW7BmnDjayNJzEAMq3gUjr3iypADUM38mP1mdNZVUv4TuKhjTs6CKpRWZ2
rPLxd8mzDGMm80dCE5tj4QXGUy8R/Y85ugJR1IpCSMzHDMnSzSQ7Kgmel1pzip03F+NZSJfF8FBE
WA7/gzzPI50cvuXXDazgdFve7CJ1EWxF30iMMAHf6o+M0CgRt7TDJu0cuq3Cvl92hXahcvRixSiJ
QIt+SR2YS3rYYVF7s3LRFKmrApetOEiI5Eu5aqidzIdLp7XZqbUkMW/hEGNTaGVEH2dFwuNtZV70
JtCkMtQyV0aFkgYuT3GVmpIqMKNYbF+brf/gc04Ch9F2+pVa51EKkoxOEoqWgAvsJ3Tyi0v9mPwM
7kC0nK6cmaKlb3Rw7igEgy2bsOeu/t696Olc6zp5G1lIZgVE0YbUl6EfI/8U/6OGWleEIjdQYyCQ
FTdlXfvT3VFR7XQZ7YSO+J21dE43xgoCrsVsUAb5YydBF9CK6en7BRyRJF3/T4v4nATzPnNdqvXt
YkEOiPY40uwL5cBhO0hD/DhZhDOLty9Wrip+4AUDkfgkiLUEREbORS80vM768QRkxEFPfQxKJnC/
9csGnD4XeKa8FSeb73bsY01l9lX+oxReHwKrf0kXNgAZlfk0nhLk/LfPAa10pQV5xrQMTHMSDXg7
MiGTdnB0rRLiKmw+8b3jt+FuwtWaehfZJcrYgvyxWPeCgDxgsMxRAiB9nc3Hj0O+30iB4+SM93U1
sun5x6MMKUOtGrZfGT5YXM/SRy+7g/EKUZRsuqQ7yJtIhwLfk0BH6jp8mkD5+XE6aArayzIcvsXq
oTMwxcJdzTcxlnWSvxyOBLpW+uKohF+5Qmrkt29tFYGSOSRve5LrV6raggh1r8pBx7Jx/CBzIbLn
CT89y9K8Tnz/X2l1Uww86j0QAwyVybZDm+R58hPh3y4t57dmzhaSASJVAV0pQRAnJAa9+/BIFrus
AaLdcOlWNrrkJvcjsHpQSJRRjmT0uKH8vtQVqnuFPAWlXQhpdGK0PoSJdGHKqunKHF6ZSbAT76Ci
pu1H8Y48BulD1iw4xRKP7oQNZA/5fPxNtjJEu4wByRjY8CSNUjUzlYv0a8T4H0Ik8woqOeFb910g
eFE9UOXUAE25I72+HexIFQUSVs2PvP+BqriqVcFYcSkjsUtZpYCYkftms0U2tC27qDK7OD43LPls
tIO0hdt5Vf+ZP9DcBJQhJPl0F905vEi9Bmej15iGd596HE8EhAf0pw9e/fx69NFxEC6uV5D/BfIL
Vddxjoz6QmnKtm/MXRPRSMeOoBf7wpaBz1gb0dAUH9n+gNNL0IPeKrEwHrZH86Lg2W1RND0rMI0x
r3Cg0hOIxOW0O3UyCkjojR64/j8SVA/jrn12Ot1oURJu5LbOMbSLA9c2eOmGyYo908ICDmz+DIkh
CIOGVBXD4XWWaPap7cLUHUbYVfBiiMTuaFzdVC5Uu5IOSljgewCyTTdXxD1/aMSCklAU69/ajJrj
M5+tGo9ROV6glQyZWe0loRC3F6zQFDWryoZOPCoLwNGzHkujEl3nkRuN7Y0IJUhF2iXro3MFuoTq
8nDmhp4/DN55swrJa8q7an/HziWbJp9HT5UmQNOAG7segC5qoigFuNjy0KieVFpXxf6ItkPEcmfQ
66yNZhV0nTjR7Gc24hK6XAmbuq/aAlC4XwqecYTU8fGcjQ90Orz0Q9677x9jeE9VicE2HsRccypZ
Vg57vMFqR2GplsahGy8keMHnOdR0vcFgFIOcNoia225lS4cQj5bMeXXE03LUJyg0EHzn0XKb3u18
XRIBe7gE1SAS6shLsGcPcpoqD3VtRtW4PXDrkY+I394nhvXjr6fUO7Sd4IIRmfpp8w6AgKXJGSCA
SyQfRczm/hTx6IJZ71RpWlZbcOspREVnESa6RxNqPKvpnjZ7q0Cm7aJjeGNgm806OfvN6XV/0UYA
XVYIjUnQxfyqJK5MgGuBlenItxOCyXUfS8Ew/IvrLT2qgApq2RBj1+w6PmDEF5QUaB/3002333VM
Vptg71paRCuf7mloBh7vQvkHWFcGoPMpT8B2bzSEcCTrQgCi0/kcTzJWOj9TyMyaUFX7NhTJG3OL
d5reWVMyI4ni+SWs8q7FB8Sx30OvNQ9E9AHPYeZN34ghqp9ZVUKHdisqGHJ+8STP/LIBFu84KEMv
V2Fhsnd7f2xFo19oNxn7vXD/vsHkHS3aViouraNQMzwxh7CxdNCDXlXo7suN/2v4G1ChxXcnUFZW
Xpu1wP6gHW6HtHGkN5ZDraV4fjtw31PzoLCptjRpOm/PgHPQL+cDkcgKY+olUr2zL4lPFZJDM7NT
3r6hQ7EoLaMAUKbsTtQs57u0vNTcmqLEcqVG+vr+EEkUGRWvpqujRwe/qRMElJZ7/bo9D0bbHPvl
FmBnD8aG/1q5+kFNCDKb7leOjiKt4kWEOmXYola1XRR23k1/TJQ0DJzzo6a4Kiw0GLWG2bA1gF4H
2AK8lRM9n/dAhnc6wt2g1RFieelDjm9vR2kbUPqF9N8I4zUr6+IYdxxo7f+ZZSaj2f9OGuuL4wVv
vWNzsmFprpkqInlU/LHxKePfxtEPLYNjD1O7UX/Be4idGtUy9u1ZUR/Pox10evREgegt5klEJ4cH
XYWlHJjMd2ULgINPINHxywZTTmfqUnk310tcn0FlUPiNdS6xy0xBoW69bmhJwYNHuLuE9mHHFXw4
oYKmet/wxYifydnb4+Z/c5B+/5okDNkZTzOdaeUlscVku9dYRkCI4KjjJaumhS5oniLN5ZpuLecB
a9IRVhb+8MnaeXICIEbsOChWBmfbe91ao8HmiN26qs8kcfdU9UwE7BFBIakXiJ/lf5CaPOIFm0bO
HAg5IPibNV9uEjpPLZu0Uj9KHxk7r9Civ4OK7m7+Yy1ivwggs1XQuTGdma2j+ouHDwItYkHeL1dA
sNlRzQn6hQBTfNaJ6k4dYFxKeUQRuRMREkxV5gV0QeT9h8XVMginI2r/ijkdd6wRjy4t/i67pntn
PJUdwvfImC3d2JvmoEsK9/d6i/xHa/NU+aXqrdedKdBbekrhxLUfsOUGsIbyeDhmDqiECiFnt+va
69j7jmx7voVN4PoDm9CJi1u63lceeD59SwMakA8otFzkKf4qx/ubJ5CEvnUQdYg5iGH7iFmoI8Hx
VSqoGnBGRaoS6PjnCVBcEZintDAprW1q5PaXhOG2UpkMHqgbkkmGg08uNS+JCs7Fv5y7Z/DMCljg
hHI0hNfvCVa3iBnfobom1MN8wI9FBzadeNhhCSLx1alV6YVYc4qrrny07mmX1sgmbrM+pRygofDo
0y09fosiMPh6eCOrXzx4Hl6kbhcoGo3pttBPGOkdVMF+hy9rP9WTqvIZ0jfmAI3JYstgeW4Anaqu
2S1pSIkpmb9gH3ZcUZFUzxJHNlZPQAWn0Nq78FOiE026cMVasDje5enL+FGcZPA9KxSqIl40c3VE
hw4J9F8qdp69GN9cbo15m49d4E1Wdl1ucJx1881H7NaLSxYE3wzO9pl2C2jPYc0oP3K+AAhySd94
WAhIvGIpq8F9JiXvNGHHuUsBeUV66yKa6qTIL8b5kz7lXrXWMPHO+qI+fOoBv6W6omWtjE5O+PzX
jU3IPkpATZBdAdQH9DOa6+QozXa3hHjtlX2gQ5+nhzy5lNocsxIULdKUoraMGz2aK5KCQWd39OsB
61pSaNAbYU7F6kX4kioUPTox+7xMTT+AcsJDLrrRGSDPPhCA+cIjxR0pOgXcVAOox73b/pzs7DYx
3NRMRkRE91mpNO42mk3i/VjbMfMVArjxjeMBJKT6pu7zT7eqWv9pJYATQjwSweUIj5j0Cgm0jv4G
Z4joDE7eD6jadUYH5YTuHvuOOZSW481A40CZ1HTIQvle6D5jL3LfOV7Z9rEhJDxntajjIkD/cKdP
7lL8UabF5BMxFe33Y6iQAFs6fYBzQfAS31fjJyzUkAGBnlhpfHec1gmNbujrG8ugIOQCeOFZ8kDR
GOnCRMhTLpnx+PjRmYb+10Z8c4WbzUH1QkYGjp5YKcwT994blJJbezG8TSIqCmNyNEZRPR09brKL
CHgZ9FpDMSdDr8gp3WxQP2a/tkwbV4BXpW0wdXkCdgXECE/KBwykqekWybzT3wu7V0PzIsljMoMS
t0QeSjAFhkap8fNC1dhmWk8Bi/lOKs8nJjSUUZNFO7kHlXnhW9LswDy+grj6B5Iz7wlDJGGIrBeL
pfUYsI+S7in2tdqKFVarG1lnMi9xNTuOeumren9LLPPoD9b/3ld9ubQlEsjrEfO7ZJqXCdVI1dfr
22agA2UAQcu10GbO93Zkx29jTVJtWidAI1KKFMAh1htIanhgjGtc+h3wivOmr8bI9vAL1hdDMXYR
67BBHh5XCRs0yzq/lEN+9WwwCLl/egXjqqM2Mqc8kAFqGfoR5LbZQZtMOPCZEWbyhkHAfDGBHO0Z
FuYunwYRyBv/dGF9n7itlwuK8NhkYwh6NA4fjPHASmAjoyY5HbBZxz4OgeO3g66XbCOHmhmkfpVl
uwAJhjXSmVVaq9b2Zmsbebmxa25PIIaNeClriCoiCgdZil186hFcxek9W0Z2YjQVpoH55dWw7zG5
f2js4dAOUjtiuh1uJiFqgqS8go5lgXrSFWYpNtIldvMgMpzfJCc+b9J5REOJYvnyfaJpvE9oOLz6
t8xC6AK24v9UTjsw8dELP7xKAgd0UYNTtQKDQS36SbF7r5GIVjDa9wK1Ua1TiTR+8NINNfDgLI/A
LCGC3bKD4Ka6iST8yyyzrg6S7jBAq3aHpTil0IQJLpKTwMZ6La3+hvgOvkM3d0MvJZvYecV8CGOH
3XpUFsRUyUxdXcMo+KmIduuGgQncLuvhBipaSTswMW0hu6ZiOH9y+J2n956NlL12VPq18kALeWsV
Ql7OwvuwLFTZqqPCkZD5DRou3GSksvd0U00o1lxrBC+K1UC8fdG7oTWml9CLUVAMTOFVwLqryWgH
J8Efc90u9wXKHRScKaOgeUQm8BgLRSdKXSJQFhe9Bth+i3KWt9lIbbcmupo7Pp/HcTRLIYspoiwu
W9yAhlz79dsUZo0+pnQ9guZSOZ/tGpV2HCeRKUm8BZQ6jlfPuGMwd/iLYLQ12PBWPJpD+iA0C7WU
g8tww624mNzEHaeB2l3jvc7ctf1I0ANQEQMaO2yJt/tkz1XTfj24hFgTGBgPl4AqIr21RhBiES0p
gJD9URJEMfpGsls7cqVfbi6a1OkLfjG7r0yXVVLQD59EmTSDtXdL7N1gRn7C8bn/6lGfc4gD5+eU
Y4MUNEIOh/YvKY79oUOaopj936fQmeySvHcUoc8OiyzzUyD/nb2p7WKaaoW01DcZlP+KtOeznSOd
rwJBenMJU0S6+dCn3DToGi7d7/DzTZryWDQgDroA5k5pbfOvfhpsUfRl7zCM9ayExmJMuza3ta4o
VmpaBmmganFupVZqRB3Rakko4TDd2a3dv2IbE3XcHmIzH0TKy828gy9zvGw6EYNg04dueE2iG0wM
4WWq7qOulqb0o+7GxdskiFVknnpfJyzjSXkfCtpYp5PZZLQpjjqBpWdHdmGVxwwpBE5ZSR5Ez3xe
uRCMj7abo283N92dzDw3dVTwSkrK6K+YIKZXmkbfcGflWNUI8mvpxd+wpX9pXu7uONSpSXyePEN0
LIevyrXWA+tD9YNpbJq2H2o+yVFpHFRQ4OAtc6Dkf15u8S5kHiriR+PmQ4pG14EMLWAYCvlP22V0
kFCbn/8lDekoHrvfbmVnZPB+psV2WEi+WcnE8MlH98ySWp3dLy5q0PkdjZuUqv5gShiLFrYoeSdB
TqfswS4N3jUJpTg2IpkJTztZ6gtGV/+vKjSD/gf5QnXdXAUyjm4a5IaOocYZNr6WcIMIR1OslR0n
TLjPL0hv/+r9XHt+GHz8zSPwpm4IOVQaS0ZaY+H16rTo3vBxm65+RsRvZzffrA0Tp8i+sK+JeuVn
GMB2PEYS4OCyohmm3QYXM+CMxm7LRjTFUcvJgf3JlIuAYpjo9AL0xP0LnWAC8y7Au6gbRXw2kWsx
hH2Vb4amM7JSOpy5Z29+6YrpL7ZLnn7/uXRvX895nRKBg0IT0K4BcrCP+LOnntcWpgXNln6rW+HU
yqzopTcjiYE6CuLj6HHBscT81368guzEYuv5Tlk1vom/4XsWbUvnguFBQWG3sv9k1//bIdmPiUMh
uVUt2idnBRPvDSUTBNHXpNho99sIZKM9SUZyUDP5tft/ACyDMaxDykd1a528EqD9oXD3o3M8ViUe
3OJpv91zTSKU6YbvUpFLX0UWuUE9vtsCw4LT4dF8/l8VPrvszxkuOPe1VTmWVrYLR5GwwKrBgH8W
CYlLourK6WXQd0sin20PMzJ70o4l2nK5wK73DE/mFbyMr0Pnjc4VKnJNxw/cyEsV1fBENzSycg5c
uHmet3Jb+zGovd8d2JZZmy0LjqMvzYRrKG64FDr+Cf3A8qY8UKQXgKMoarW73dR+A5AyoYRF8fBc
KcNcVdubwYRWRzPhFc9jFjhoKmIkhZ7SBTaYcFnJw8/fCkhHiAMSFfk5p+rTYxX7azlPmNgffenQ
1Z/ebWalzLATMj0aoFUYnw2PXNGI6Kxvoh9LMSr8/thUcaignz8QukLN+O+769VkAFAEi4ELalMb
kKvE56NZgZ+erZQ8VH6k4SaFBah87J2J4xFbYob5Kjarc/grtFlxh3a2pr5YWCKe4w97nxofTN8N
vsZuJaWOOuVlSVDDah1bzyHrFiTJ7CE3/73Aia7lC2CZy6dUJyWFOlTtK/AeHku0HGMHRMHA9Ums
xvfDZN/IuyZvdYXKkKRtRQV5XVswEkXD7bNUlYV0u4qIgZtuxUlQS4Ec/zBKXl8diwyJsRr7QyYE
jGsBp4Rh/3O9zMZJc9fiLA9L4ET4PQjJYw9leh7lPv3WEoHJjxPC41PYkaXJYnRd+aNpywFo/6I7
cVla7/yXPhL6PIBcN1cXLSz3hpq06udMeA4ALuNUwFdcQKX97/jDq+Dn9cTahUL5CmLsdyvlRUQ6
K3+T+rKP7UkC0NCg7Tm/cEW69KLQEvsOC7wKoDiXMykc1hrp19TbXlWIGsIgufGnlY/PvIbHc57m
wJA8vbZNZahN/VdySEVebx97NuormFmBhti7ccDfXOsBvPzBS9PhUchEImt5q/QbX8A9M4OLNuH5
a9dTs011Vzm7jadSAJ68lom4W2u2cXHEEGwtXVMJ80aAe4zbhgK4NPxB0ynJweEkIceLw9jwlfJY
ml+b3hnVZ7CI4AvfaXBF5pNCjxW3gNGcPuRF+ZB30qHVP2tEGU+msw2V4IBgjUhZ40tOJel2kdhD
07mH0so44YJcmPv1QxYKzIP7z+PXUdtO1LkXNmiydVN5TGHHI2hfarPHGTJzx24GndlpRVcR5/2s
Nv33a699KYdDDEKPGlPbQFMjdOgmzkH8hbqfbk8NuYn46hSdIJtZzX+fDXqGtAl4P5+GfkMVFmfq
wYVIZ2jiiQ0INpwN9xSkXhrPkK0GouDT0sm/wzLhGPu2MRVyl1B9G0YsuKIlfXhfNFUbaibBtjss
pQ8IkQQTR3gGYAoG5gZpXOv9D1zFx8bAG7+WFE7CEWNCw2T58We80rN3OTd35oT58M9VJ41wVBvx
tD23uYeRWPE3GpiXW3A/bM3UbuwLlUlJyc2KoatqhZX0XV1z2dl2y/e/s7x+z5cPWiW6q1xcp6g0
aiUyDB+xC3UBT2WzSas0/zYkI3xkeaPX5wWcthXTH5VuFZL6vrL/k0vFTQbUJENmlmS78y8LIFtA
ZpMb0Cthyd/FCtHtpQ+cekWDBhv7zpXdO7qfaD+Fq2wjDEfs9oByw7Wjc4AvuaF+AACgZJhvWK86
U4yI1+XFz/TeYANCbtVgnUTT4wDAFkFVKtUupL8uD/rM0NR0oyOBRYJ2seUro2ZpqbOmX0mAN/Dp
2ZpALY1tkMwQ1K3z0f8a7DrMATSYwAFRTz7LRPmwqH9K0ykmmZbHPnTe/uD11JYG11SKBwPKINSs
3uuOR8YUAX3PHOyFgtOpe7b1COGKz40MUu1nDkafhpeu5XsKMF/J5bsE0wZxcaQkdsRL6y7Sakvc
Niri4B8g+n+6tfsypPHYTfpnx2bmDSt/x3tCcnQMNdaaLOMxwbe8gUjI2og9UYOK3z92N5x+QjXy
rk7g/94iSEMFBTZO4uPK0og3ThBgSbG6lT2KqsHEzedf248uKLuoucd5VXOSmVA7+3CH2ihLwNVb
TRSIivT6z9sHQzBVvibbOqFWq+xJIHdq8EjiGXxk4xufc/L9RxXBnC+R9imADKiv1ulD7E2yW1G+
bB10s1CueITi+kqUl+ZaAMtrPWIOOUn2PQJq2/ySdZjRA5sjr5zId+lLkjhXfFMdrqa+KY5LSRLw
G6sQBM8wRqM5qFd5dFvzPRGRcDiWLVA9fKsHX7bQQwFx0cruJatgTEArOIMzBz67AhLghiPJWoML
FGWhEGDG/QVQxTruSj9XtRpNBBe81G7T9Lf3kfWNc0wxZRSG/UatIAKHYTvx8Vpgk3ITPapyHhqu
dmR6GVowofFwd+IGIUl+RkGA/AIGOhbMN3QRISe+VIRn2a7B4PQGZyu0hZYJyXyZNV1rrqDt3cIh
CAK+N4mPsY+S2V1R++GRLNR+VA+apnXanSoEFduC06JgsUW2/+zbpRmKrgF2ctp77QQeqPDSkUW3
UT1I/JRt19YL/jFdymxc+szpUMOfOwtOErOtc7YUqzkliVl7cn1hg9UulGkpmSBcZYk6iM3v0ivJ
N351ctsZctXKrh+DtIcpalo7vvrzGypNPTd8ktFuewMgMbBJlCutlj7Q/uaHkNSi72Tz2z2hiPnh
ZNFmFmfhxZ0dCellfLNR/OW8A+2YeaEhPbrXyH+UU0QXlWC9QtVYhAnHWg8Yn8YKjqO7EaJzKxRe
nrawccmmpzfOfDVZnHp5JKGROf9kJunZ7pS/uE/5k+CPokvLIPimhpArP8fVpNgvRRq7/PX6EwpA
Nc8WDsr764ARyuZTj6Z31q6d+vjKiCp4YJGFkXVSSvDWoweYef+Ti+UV+Y4q/TFGxAgx+tKhQw6P
765QATD1BFqrQKuPQwPopS7XNsTYNubfaMl76HzXuGB7Ahgs6HqNEi1no/Ckiiq3Ut67wU7wnx8F
H+lZgShovuNrKfSGpnRlpryB1PWlSjsdVl8+TTbQEf09/B4XdgBH6zCO7kUQU6LGkl2yhzU834Z1
URdWyFtaQRPVsKSb3MGdJPBB6VJ9zr7AR67evbIQkN5N/pjCeN97Vfz/c+OLrYWioelGYp4uxo+x
W5NrSmlsw4wqsqAqfWEkVlTlerhky2TQwkZYqEiXWeRdRiCectwt0TB+FuySyl8I+sAQj295gwTb
kHx2xuFIdcieH0hHMoPPnitQ/sHRcO4FvrexdBsaeSwdR0MaZhpwb69bDkbdCcaVNnoHfAwJ9DRz
dFubuGnNQUIcjufxZAkeI6Q3fKe+hjPhlxYZ0jDNnBk7PCTgFVGeaq75+RjZ9MblMN+O3Pze+HAM
+p6ipmZGaaTMuhl2y1ZLvhpkSvK0mYv2HOoH/2Xs5QeJ0ROwxYPmJuk/FSbH853TAbO0ut9ZZtWx
aFqXjirlRpGvr627hgZ0jaOw4Ag2fg90VJN/c50KMyhZTztQOEw/u0qabzcp6tMHWiXYl1dsL8RJ
lkjIa8zZ9MkG8O66LCTlB9f0sY1AgK5IDsW4vlXSkPwRVGlBMGCjSNYuztduAckz4Hu82oY+6uhp
aYG+QLVxPRkNPzc7slp+kEErt8i/QvJJtieAxygcLOExJesI/lBZZhtNAPgVW+OPjXXC7CwkaDp+
GAj7+iaJYmDTQvzADNLXhsGq4iEygGkccsY2w7nyPJMpSWH4gXPrDiReCNSvatlDkPRuglvOq4AP
AxqF9SzXfRYxtaA4sWJvIZAOgpuZT6grVVwwKCTtOClr83G1c/3GwsQVbyFML09yY08loO3KjpeW
K66WKCHHBRUeRDOjb42V8oPxyitYZJ3i3frp3MU58ldvpJcjuLSD7wD3hjlMc9gwEr1sLn2p8Sj4
BFGn7d7ae5MCm1asRWMRJLgpyFciByf7wW77e1GkjaiTa5L4EXUul78AMCWS517ABBYsvSXkBVtd
wiOvTbJgVFJUgG5GjTMwVtwnnrr7vEFD68JCoXPegtREKm23YoI40bQz36eaq8jdjQHoU+MN5pB9
+/JyvVr6Juzcz+k5QNaoDzgdrQCkiQE24hlz0/+HqsXjY2WJW5ZNUf09DbqvI52gjdjtLC0+inNS
27K9b9YmVad+c35FO+3n9zai6Jf/hnKHB863zoJGeRvPgHeke2FI6wVsHtGVJbyO0zEOSOGYsz9S
rmiW4mYIFUA8xc/3RIgUQTG6JIk46m09Q1FWoBERqZw0FaDEsf7blWNiylqtTWyraBUw20OR/428
1+KkGJXbuWgnTlZtE7Vi5UiIfn50VbjNM/bT/cptiiD5QHIuFyoZTA+Yb1/6KUkGKr8Vlsi8xqCd
P+ERe9hphlfKMgL/0Vc6V1S3hFHJceP992imkLxiLmadRCu5Gs2mor4Gj4J2+TpOSlFOOh6i2/Pn
iouGtx0V8YkfXUpJWZ7+tDMsDodLyFkhFA+W6RuPngdgtaSoPOPWtm148mlMlG4dciJa/GFRfbe1
e77tm7Uq9CohcxblGMM+CpAM2tHFZFvHiVClJQBgyjyyuaA0kuC/ZaOpg6fpfxQS2r6Oh3eaFm6G
IZaYFv4UEwKopS+7UyrHAbnxKU59OOofRxmesaTG6oKsGxecmrTMWuWYlKXMURakIV7bdbNAWnTM
C0Po4SJJAD6F/UPSWaTZCHVJYhZW3EKNpv2s1E+2gZ2qXDfUUv2CTFHoah7skYJ/9kAw/d6EAcuI
VO7Axied6UzC0/dCe3vFRX+jbxaWLQbUsVPwovoyHNE1g7gLohV/T5JWD3Pxwy6tihGoRkj5To3x
Fp5NS+UBGODOk47SntIGscmPtyd5rgxzlhnnNIPbpuXNZW/LFWK2DdaOF6SxT/Ukn2H4sPJYrFQT
kNPFRFLY077jsgdNxFb1dslO0vYaFeq0l2djLaQDgVCZ36huL/jHMLSfbTMPU1aWMG5m5Ghr5aEW
4JO6QSY7vh75xQyh31sNENuWb8agEIoLIX4YdKnfth4WSSwmlDJtd85LSMyd10KFhPR0lbjT3ov+
rTDNtupBnFo+d2lRVkH+PPPB2cGYA8f2LViVg2II/MUF5iww6L1fLDZJ876CYCKpITNbv0x04WH3
BWSsHGzz6Wy88SLCJAVkcpHzs7Sa/SGuFXFPctwQcSA8Xlyh0fp39M+jHMAZwE34X/2BQZkPJbRm
VjixR6++yutS58KQ2BGJunUXAPM8Yv62XeIwtaRUCwL3gujzuzh23bQs3CICPM2+Z2Q6BtHjOEFx
rhBgSKAPsW32LbnvQIf05OpM3ZyREZL8wjvYa58NjZ8REPZXS12Q/OCNYDpSm3w64+ZUZOj1LWrM
qpP+rQriZ+BkMrAbaBDiWUNnSIJTxKc2pzZo2+XD0GhhfbL9dQ1gw8ntZ5EFrFy0XMu5I/14CPBN
3EO0DPNQnQdPMjxoizsHV2mhQx26o9PHeSNLhDaME/vReyhFVeBOk2sdhhd2czt2Nzm5VTxziIg+
as9nr6JtJCu7nKgmnERAC/nfusvaFqrg2XNcdQRRRMa4eibgUYfSCENMfMPTkd776I2A2MnzhFQt
jfJSpRJ1kldl01Lerw1YfReEhLgt+XXSXtZNn2+9Sm7lBnOtQvtngvcABuXQUUHCMVfHqBA2uPa5
wA3NR27dM3Hh39N4wI7inyjq06y230RbpZWDzr0V+Rnbcg3qRJA+FszprPHcfLWcHHt4wiCeed2m
OumqlqL5pTenS3TIi+ZD0Dft/kDrRJhnAeW1fK3i8qzn0HGYWKACtUtmqJB+dMKjzOHfvJVu8m8r
0kjw6uSKT4F5Im7wZq4z9WrKlgn46ZWdK1YTU/iLs8Jl7Ws5QIiE14MiPVeDnDPR9t3eoOltGkio
UrbwebjoYhoIerijaVt76Ho9J0t2o/OHgzxayhxjxyTllTysg+NQ1TqItvxJjSP4kfP8VeUYJnXb
He79fNo92xdqBMxluaaRQvcWaeU99F2gyYkYSdlWvjm79hxgP+d+w+GoiONhTbZZQY4as+S3Z/nr
IZRQiidkK5oH170XeyxLfnVaYgz6vjHVzgxPRAY1Z3pIRPc5OPNdtmjg58sh80g1KpT7f2yFjmme
KzbGgJH4opX3PEImQaqx3thpLvDCcRk2amHeiW854pXdSwbacI6RCuiLLD+SjQeIHLmCNIQyccUr
sBTCqOlslDs/GWhPOGPr1R++HXvtulh4jKRs0JWXUoPumUUGfOz7RGf9HdK7+RYViXRXKGJIucTr
JCfO8IprHKcbMRMaRIP4ZLGmG4SLG2YT3mOjo4p9UWvtPo2ayGe6ehpZwJx52+wjI6OYs/ED0/Sv
DD0Bz/UoHpSPYQL1IrS26NgRxh+KstTHTl9sm6BrUzEZNjipjkYOdGkBjLVxqEkcPhpRJ9DH1DBD
8ozNr/faBWksXwb8h/BfG9nIFN2aCXuPmuhUtbf4IeckBALVqoWxNB6PPWYvgqh8vH2m4YnTHYOJ
aSCzUkFbFY/BoPV22fhTdq7xn8q35XiqL/qePdhoauG90tcTiKOG/a4QjAlJWm0xmfr+pdGyEts3
d8vLQrJmQbZeuDlkeFG8MEqFVtPnQDzT1bzM6LuXeuUkkVsL9KoAYikywpfWtS15mk4PqukySVZv
Qm2hS0rKEvc4Ybg9ObEFdkHGrtnPqqvvngS6aLZB+QnzPjKEOpoEM2TmmORhQnU7ym1pdswRdL/7
eu6o2aaFXpqECzpkXO6Ucac+b1DIX30qW9GUXRl3MJl85uZtJaRzNabEQnidiDdnbq/2SAgzrkhF
zpFr5Yi1B6NI2pIU4/PfR+1QhBp8l2FfzT/ZkQiKQV21fJ0wJ1Fr2QKFS+e8kmp3O8ZoSc1F3QkJ
MRm5wdyX4eSKcVV4j9R5rv1xumWq+AXSoKN6u0qOVcmdv5ZKjsQqujjPTKsjdJ+ivKmbNTqQYt9X
xJwDLfHLDCbAzf5s6OAwx8L/QwvJwTgh/lc61jEZjcVQARuQgEqGH/goRgCnsQp+YNjmbTvlF74O
vU0MOciKuB6f8yN0HNEJ4AD6DH9vOhXdVVnDoseiquO6HvDONhI1czaa1B2wT/s21FsE/4HBfBIT
C9/KzDNjZWc1+cTE/lTITCBq4slX0fKgOornR0XSw6TpxCqGsxLiMfrgSRJvlAJMHFhtAqs33En6
A4jMJuOWs/07ROsFwXRn+bqKQH2aeIt2mmE3/n6LLjNLXhVUS7iPXpAJBibWhknomXKeBXZdhtPE
wafOvsmzFDw39o6v4DpA3pgutX7GijaJbo90CFNf3E8ByqZGieFjbS1hpAx4P0wxyjteI1AOmkwC
kcUedKdl0AO2394/2iTXgfTtsjkR4NRz+NgGiDHDpsYieATFEIv8kMF0y55+z0erlovVgrmvdfxM
I47vWYhtOPX7DdVRMHvO4F5BcSjW9iw5AJYKbBHxR09Z3mt7Y0uweYBA8s3QNYQ7iXZzF0KjQbKJ
a/Zd2HQ/OMagFIhb/68od06m500KXcDZTrmMsPHDwRZb2aSWzUtfX/GobL3z/d+N4ah53xIDyGOo
HuWLhtZu7td9QKXY6z0WfxDjM/dRnyHw2AdrOWwJBg4x7k78ueH9vphYGMtzuPwYRhFGcWtnz0sT
jlazXSoEUGg5hmI0Ei3oeQmDf30qP3CkgLSWB+H2mP3PWiaRiAzXLDA641NfKGZZvcKD4NJj7fkP
Iw9/jsmmeCWU1MdgS45+LT7QXkqCOAEfWK47mRaV4IKCyfaUmbS8+KCYjANmH5fTN0a8BgDbcpOo
zlk8uPhgiwN3NiFL5AVJghtRbEsMmjYreTzlvCe11vfoqyAC/B/VCZVPtZUhjlCcoWeweGS23+uM
VWzIdEXX7R+vKicoOv6oE/QcpIMO2LKHBYSlzNQjnxKBZs7tV5wlq4pUnEFbayRKWpAX3VSrh4XE
b1kcEdJAIIq+t7C7XlF0bZT6LV/AT1yN8vUeqTinggQQzKtl/2EXgOEepXP/XatX3U2bjHyORrMh
xzmuozxJlopk1iQuXxRqK1LpSm6+w8JnaKLTFiXyT9tVDnSq8gZcww1OcgE4x2BHZSJa1J473Yao
DBPP2JZcSHDJW1H51zuXPNhcvVwLM9CxEzzANV+iRbtNS1fLUafrsawJUH98Cls0ChF7n3E8IlUn
sCRBrPm9J6xx3OT/c0CzMyuUig1Kz9FTkWTeNfAXmI2OQVyJ4+Xm+IVqjk1DLgq+JNlLbelElcKG
HS0qKYTtRSDcLMSxIqckd/v8xUU8vKc6Zjvtd5FwKPGsI/TtKutDIJKse7TsiHHxTdSyDnFi2Y32
PYha3Gq+qB3tAbW5x8vKbg9Dd6qZCbxqDxSIdKDA4C0cCC9dMmvx29qeaHP4ZnSVcnP5KGvVSFxg
/E46vVbbuecrJWUgQtdLQFj9lipXlw4TfA8rx03WylA1TaigRV33An5VMcAdyDX60EOwE+jKBxEc
qnskTAukNH8Cgl9sQHIjs7Dw8NK7gInpjetaT2QpjL/inu/JqvloH/6tA6d5y1kGd89yGdOfdPza
mQaD6mlkyi/uaG1lhOxUS5qGOG++9bDI44Z8Ye9/K7A4ZcKFaPGoOqu4mSS7S968ImPR8TxLvCIr
jc6PbnjPpe509LP/CS/2PyT+RNgL4G9Ybr+kBwaRWe/Kslw27TYvoUa7LxOlQIodWYaRDfGanJ7u
VA4HuPwwHZaV5elj+aDPk/SULfyQCkd39bCypMEaJ33v9flfWFy00v3KPd+JLcTrepESd3niGMcA
YqbC0zKkpRDy8VY5V1qADLXbh6XSNW+wK8yFNQoPOzz7YC06HJVdnEEf1bWXoZMV70zlKbuBORh1
RtHt2V/oyA4+SD3QFRuLA0sMVoCaL+GBUfvQix/GAO4rEKyf/j9BN3GJMCc53lxWhoLIXzwxzwtg
u1G6AXHizWIIq8LtfImAMp6s6aIKteCcbKIi2AKEXZGwLtcLgpOOuT0/4ypR8Wok/dGTdHHaeeRf
TSRIC/vKaVT5MzjFZlFX9gqxTlCiCASLrQIOfRDVOdCjeeLyGxLm6yTXKVD2FI946du0rOPxEKFM
rV2lKKfNl4pbHHnREPLfrmXWosZX/9N/0k0ckeqfdryS+E+HKIWqNtHA+p081McSXRuRxByvdE3X
4u96wydCuIoFvVuoJ4w4PpOnFiUx2Jlt/U2lRE1ZlQLs0lxpSi+eUN4roB/wNZdsxUuLOk/xKy74
+nMUQty7vohdm2gUiKAmeWYcXejnw47EwEpzw5JeycuiH5V5+zjASoRAhvI4aGc6XYjir+DaE6F6
9KSnuBp7yOYDv54oEc6vKNuhCBo+F9UG1zuw2ZRHrTjESH/JyoCwY5KCzarKnpZhuZx/QbhShFsU
5vC9Ka4is6oI+hL7cJRv0lBhbiX44qjOeWGF88xzLH7ZZoOnlfCzZ+whEDabchG9JtJOAxXPMIEH
Xe657b/bpmJVXoMVP43t+Bb1hKq10S8ugRbh69Ydd9rx0Tg2J9UkBTxEmTwS/dUkMIUTdj/Pnoht
N8thSIoHkGgOMbUZTs73toMrUdhBVFesxW/oLLzo7+E9J+v8a2hE3PuGMe24Ip47KAzzmwSpAchF
BPlH0UVHKkaBqlg6KfOntL1twLtUg41LHda+SGXMXCSmxoFqFLtw2f3sg/qzqPifjOJ0td7oxkpC
f6JkN2/PbPfK8QqdUBkgzXlKzCsGmkMWNRgU4+754ksGpobd0L65cZ145FP2REJPJRdwfmatLnuH
jvJJKi5T4I+whodLYD5fDL7/ISBmWeAgXsMB7yVfSgIMROCDU6uySsv6QOrVGMNCb7cD3G0Jl7qL
ox+F/d57nvCGlSe/9R81TmeHRLzBvn6B7OwxhVCDoXnCvtDP7j8I1d0mpEI9yBTb3ut9msagY189
hGJkyt/RirvFD897oVEAECipp5izNuZC75kBZx4sjNmnya7igTAMS/GcTsPDVZdLJhvJoGuEpQ72
RqBMwLPlXPMIYUMwMxZaeezh4DEp5ZUZmpmJKm26TIbUcy1Q8xlCaxZEj+F6UJUhUJJV3QQHCqV1
sRYxCe8pi2i5Gq8+pVxgx5I17IaaYLKiLKBHOCfZvVtHQC20//MOgdYh7UkuYmv0R56YRWfLLefx
UzBoUBpOS9mzvXF19BRw09v6Fc5tJd/szrY952e0mAvFUbU01ZO7kV1czN1cN5ciB8P/zB/SAJJG
EBbyWimx2HAMokiMjGw8xbA6ldDwvNC0inYLf4Mc+4CtDYxTSyGn2CYnumED3dQHNmx6AVfZq68t
gYIBzVfw6xupPZ4J1e2np2MBIyfiFD75Zyd6PCWYMj5EoId8cjSrunrxn0tqj6ENHJp9bdcZswwX
RqQq9f2wIQeJo9or8u11ZB3+eqH6sDpSBnti9t5LEeRpKV9sHUjlPtLr4EUnRo8UG2kolYXrDH44
yz/OV5CQx+ikxw2wJIE3I0+tSgLPJka3SyBionQlEtKEz7nu9OiQPPT1qS3fIJgvpwrmKu0fylT6
xcY9CL0KVySr2IGPQSjtTtjRMAmufiu3y8W219RrxcNvd8hv9FsJCd6whEpmnUohYJlxDoDV3Wms
zrZmGpKitmmyYoFC3vO5lUMuxDk6Wr5gjXmW95rHhLjTY6Qa/bvlqvr/SSUPQhJEem+WSTvJtJrb
seAWTozjfuQ9RYwCaDjP9dpfl6m+G4v5AcFq+oYHTzPxnqGijak0lNWz/wShbGdakK3wWd457k9Q
EIIZ10+zY6z7CtJhjaHCafSS0G0SJ0mYCxZpk877ayCsY84ARuqnK+4eklJm8rmQ3OjX5eW/dLsv
xb11xYOzGbc12Ga7aO0ohdbR9bGsjzr9yXttp6sERqQqd7INtBfD+8keEJ8ZgIueY0NhjKtjzbmY
b31Y23qClk/aRGu1OVz9BQEcVhgsFeRhBPwgsAFq2HCqG9ZiwL1MYBQcuV9E0AO/oxj7ccf/RrRF
tGfIoWK7MGpDaMwMv51ThtEwdHWo7p1IGay5yqhi6sHldpSbR+Pj7bUftYURcBcRVTj3wqwR9MQo
jbHbHL0NR3gZYMXIhkalxFNeJuvqescgcVGZfeiYjyrDS9v9WcKeNWJZnt7aWbaR19/HWJDlgAP4
/o2jFU8rQT6mmfVnZ+vDEaWI/rD+lgVcZoNKalIglCd/dqktvfkXrczAoCv96BC0v4FNhXDn9Dms
R6SOkLbxlffCmRvnfJJnDyKQ/TEIGCchjGhZKHEDpCpVxKHXu7KLqzXTIiIg0VC4Pc3ZabKaeLuT
gho3AG9xGiuzO920T6stN7mYjE0luGsSWsroP2jAWY5SVsPlLqgjLK1i+gBsWqOxwZ1XDrw68e6K
IFw6fAdSQ/lwszfaPbNMmWIbyGKB3MNN/VX85mkAGgyQm0FhfxI38AtPoIahNp1IhMxTKH+j0LfC
b7CJkB/sqJFWoebJZ6dMtg3dRhznn5aXUOAe+F+Ig+JDZaIrbw0qf5xn/Aph8/71oLoQJTHyaCBU
8X8Xyvs1936hSCjza14g9NISkBMH9yJdErqRAldw3t4fIIN/O/jvtkM2pAoEvORoHIOX8X1vKvKx
gGMhcemgcmePGgclfxGwWtnn66iejgnu9faWjNsIAEgynWw7F1BdpM8DLlXOCHPRVi/JL9+eSv4F
Ozjp3ItNaPBpGqgmcmykFjCRjTLaX4mPAvKsbYPFXL344EStXSnRess9JgQ3kqJXJLEv+IUmeTWX
boSl87LTmcj7awhAJaQu8fvBG0X0ak0jz0+KFxpJ1W+IpQlkNrE8ybwtqautCgGKPJa6lAVJNmZv
OJwvTnt75rTprvjtOOo32fUMkgD15+yM7W9eQNJjs+4wZMxp7m4cWiUnXNOVGJinNCfOkO9mz7QQ
HQB/zwozphOkrU9cgHkK8Hcx30vSbMGZ8mz23bHET/G18RW12VxPRdKTnkTYRwQqGFwSkRKnnpgk
1C6d3SuBczX1VtZxGF+e4/zCzx289msHxbPxMRVPzGuj6nXcR3yu3yUaFAVokpOBu2ur/ZMOU1OK
G9m6W+MQGPSLTpsJtFd/HArT0szMc6pS87pfQ5QFMBMxe7APl4j7eUOLDpDjOgdvi+XuJlt1co52
dr3oT48HEpvwq0+gScSAX/qR6qt9pwU/uJN7RdBGr8WgQJRtXUf9GqJUVgKEI7SSc30oqEEX3Utb
RJit6ZvPPpDtILh5wcypSlwaGgR9C2FQnGOew6gu3HZtxcIkxSA0b+2MTHouOL1dbLrvXzicb8b0
5QDu3s0qhfJlAAaiYViI94CVlYc+sQud2ECkP/Nn5srfkqzRCiHx3M6lSiCPRwC7T63es8keu4e5
eXxH1Eu8RqZTSgb6oIXgK3Ic/fR0g7oXnlY2CRty+0bcWhA6q4wBP8Yh6z39FQE82I9/r6UNymqG
G8Skio2ZxbHrOPZFmTBRvbVVPnX1l1yHPo7A7lJsGj526Ud7tSqaUPP0YQjnLeCMlQNpbAH0ftaC
rpF/W2fKjsnshxzMJmc/D/Lrnqrbdi7bOjLs7yyb980P6HCHgC4UpYvE1ESTiTXRouZblSQNgUsQ
Mgxp2JKEYwCUZBqXFDKKhHi8vhDJYb+CZ5OFSpikgWrnODU5L+i6M68xr2GAFm8ysXXUaSn+P/BI
xF3uamZTMgGt7Ts84qT5lnp93G9zdagZ3pwEjrBBgHXmflsKyzioG2lOQZCQXuXUeFW2mfuXzAHq
nEQvyp/LC9LsUQ3uBrhWQKJZOjcglkiRAbYBdPTxjslcI6ZoIyH2ekfhS0sBexncpxQzy+s4Ew68
7Q2uDCw1WiHzXKwKW0lgBBeACzH1YaaDCj96aWgAeNaKtDJQcOL1Fk41goBo+YgSdCo93ijOEmUp
BJ97NzLTux/EJ+5LsG7xDcsrqvJW25G3Trdgaem6mBM0Q1RLtYQE+WJSqPcxSuSBlkwzDuDnK4Ru
z46hTvwunkCeUKVpj+J1esjcyliD5aBBHIMInmRLdX54+awZyHEDhxW2cbnMqIsAkG89+42AS83N
LZFwWYt8pensXIvUg95MAeLUVRbNAoKlpFigM7a/4KSricFpbIN3UA9UKi4E4QuIZsr49/Be/6Zi
+JcHMUugpw81tVIqeTd5v/IzotAtPED25lpOgXJ54hdjzR8sfUwzaa/pDyTY3xz61++i2MtuaWxX
2U9opxYqjV6UeQ+JHgRFYC5Ts5SU9fYv0hYP14koZtRunsT92W4R3c1K3ZHZXhIzrh2RjcOVf3gf
N4HS8y5SO3praPeQ4h5A2I0WSpFkRk0Z6K+e9Te4YwcYECH5YLLV13yTpOYYEemgP5oR/K50e5/W
rQx607HOUlPzCSbC6wv8W9O+hrZEucOYniy1YAZEl+kJrJdPwc8N5v+A1HflCIUuG7SBGZgsPpHk
ilMEFXbPAxyf5rSTi2KANoUcaavz5AT6zfoBa8J0msaMLMqYammtHN2UCuJyG/+NgVsdCoXUvvpW
I4yCJAxh3+sdiPTdtx4ipeKOpAQir1xPJQl7WsPu5HeZ3kCiNxdpkGSoXvE9S8NM96yDLhG88vIo
/4m/xfwbR1lhoYow0/fH/PMJtA2Au7h+G2q0mM4gIlSKS/LDE788ZA0zcYOzQGCs6tznYa39lioS
06OzdjlSWZrhpu5ENYsIjEajyji5uDpFr18hXJWHKVwSHajzsJ5Iq0lpR2Wt0FFCkh7ugx7/rvPV
oHE2pWa/7/mO6EIblMaXGNm33GsZFbsGs8S0/zaEAdMXxImAgAo/J/gdiUODjkyISwMsz7CYpA07
ZRMyY52T7+XqUNYiZb/4b9PdQbNYXRuQYzl73IXrVEZ6143sct0gVxzxWirp17Dgsp+JHy4nk/Ga
9e2qUu40i7eVaO/r5x2d1awd9NcYbcp2xQyZEIaaq72CTn6MnU7IggTps4toPx57KHgck1oop5rk
NReiWomE1X8AVc9FluheUmqk58RwU6lR3DkOOHAG35l4BFnu12vs35IfrMk5C9lczYifgZ6W32FP
ZG4C1KK2DmU4N+OQi4qP45TjCKQwoKx23+i4flZo32vJmPu1yyvZvGwgQCcb39wO3TtqO5h4WOny
VPo+U0lUqhGEfxpBzZFZMislZxzEhPCYfgCUmncLuwoMvwZ0i5zjM5N0INP/dc7bFKm3Ty/4FSXN
NGoVsEHgkVzUE9vfJsZasAAMYoJd/vCGRUZAWPOwU+hyVeEzgCxVNjnwUE64+LfLxjiA8tJt0udU
2WCYLlXTAHT2mjWecOx5pXHCF23MBSg1SCh6/enKhMvqwFBiZ/pvLXHTmf0FrT4nDE2jUdxw3D0w
ptpMz4hL7fFx92dodfNNv2WIpudm3OZ180zxwhqPsImHHlMQexszqeYnvJiymwGOJkOTHXVJymId
IIaOmxSGRBTdJsRH7dUi18oYfzXoEnmuAclJrZozxU5Mxxmo+MAuuNQIrK0+f/dOw+Uu8SajBdET
H9LcrsuZI3nG27lMXLxZrsMu3QlTlpClrTtMUMaSWddKTF2a3sSRwYn2d2XrAxxkpIYTTj0GSXCq
0SxLwFm/wxqHH/y3reCI60FrZdQQCpS5DOxuRNVsNzp7auKYyM936+jIYN5+4Co+G/DHKyuwd2nW
YDpHSe3fXNbr8U0erfDlGg4snMYJ/hp+M54MVtF8h/aOmx8WAvnfFitdlTajo+PXiWRNLFvh7cWU
wVv+e9jrgDwgIiHGp3pvE+9GGy2Fbn9RYa2+1nzuFcuNZvmJYBAWJC9oUz3qQs4EJEmlup3O1nKo
Wv503ugUtwb+q1B5e3Tx+3xXWPJnrRZxamvadtywtuvbkCuZgfLdkl1NaEBHvHncGXlD4Nne4yqi
A1UhyJ1uliGz/iI3ZVXoCZvbjX+hqvVajf05i/9EfFWIf9yVVVgg7frwjdKnM5WwSkQCgeiOIrD3
Pp+yN5OJZEnUt0IprfAO8qN6Hn2F4cX20VtcHfcpaI8bWtbRbb4iy3ssjDeiNEqi81tAHOQd7xpd
dJm/YZ/IU52pCFVl/5xYrU4XEES9oPxjj8Dpbnl0X3BAIwKVlAZBSueWI5zvVty/m1gKqVy3kSKZ
7ZsTcUz4dgVQByAjTqPpP06NHwQybbVmOs8bsgYOMEFtU1ruMqFOKX9Y9HnTzeqWtq9X/qgJcYBz
d08f5hlypyxNjWQebRCnBRMpfCDJhVXdZ+XiPdt7KsNjomqNAcDBoc6M4VaobPpjB1O8oT5ubrtH
9p7WS3WjmNCncBj5MsuIk2KWMcR3d4ncKHNMkV9fFiLwBBufViVPY0bKKNC7L4BhS6RpZgcW40hQ
QOEspLzf+FVIvajQjTqP8d+q/cavG1ThlTIRfEUgP4eI84lujXuSSMV2aGDn6wnKSP9YABc2mBgC
XpC09hv4j+O+jGFQ9ex10Zg5MpA6KrKfvGuEsgJSa+quNzZeIuxRisSESBN4JBxuK3FjqcvB91lm
2YyOA09wG5bmyn4y1E8/p52S6dVH2c5xaO36zZa2icvJADQlgkqY+657AfHGBouCUDUHkrU/UXvV
vfOPiVjl48D1s7Y4R9ZilVyQaJEpzMJduQEhLYkyfP0iDrrkRAzQn18phHqutJsuG4zOTuGtVwLR
2KakpKmwvvteENUd8Mpi1qOgFtO+gRmxZXHS96yrc4MZ0DeUNbsj4tGnaFJFsTmshbw1EFE9cZmO
1Y8+Swmp5A4nrs1qGdgcUKaILy/2TIVGqES+tcQ8rjv25UU2MTHNVkTJh+tVrC4nKiUBgw/v33cq
blKupkoNnvwbqMyJIDOZm2NTMay5QX/0LoxoUVuNjp5g3LBaACeU/9rB+xf+/IUVeTfj0L2FLM3A
MrTuI0ycGOgoIDfwV0hiTSg3TqKzEVP5jBS35D3s6m6sdQvnen0QO1J4+Ld+SVrsk6ddtiii8YT8
Vt8zgpeXxG5K2/YhorsZEzYHKrHNYkTljS/DRQReDIc+qadoTQNqIJsBhYVcIYSb6TOjj5KcXRmj
7jNxIlAtxhizUxkGTkKc1u5oSmhsaL9dvjgfsnNMoF3A14NH2ORixp+UpCzrDxAWFxw5CE/8SxnM
GLSCm1Gd6WQOY1g1xZjrwoL6baGHwRpDNe3bc8qiIrxSuggXANp0FM5V6qXMG85lnJNlfYBczyjJ
DxPLwqlWznmk8BBl2gSqTxamXaHhei5NxCu3i8w8tIda4kEbn01MgoJO0aRozCk5TmQFtVjzawyP
YmFAr+QXzhg/tiPjNSBS3O0SGU0R6HYSlKKlZRDZaBf0oHOryevHfEbGNFFUS0xwTBcscZ4MHAgf
0DiHz3mtceAcRLpt3jSGBI56FgiRDm4c5dCAY7u+sSpgUOgDRvoJWDEOXYeBf6PKMWWUzYhkYQU+
+WFTRPUsu9B5ogGrjH13KdMNspDLflkB27cfj8xxE2dgPUrJUPp/hiamhos9QA67MlqDTTKw/qw7
83GWR4G2HepCewErIs7i2OwPAJTyQgMULjGiL+kjee6aN77dYz+gQuGh7PKEhQHP6iMI+eUiCz7P
LpdZ5h6/KYEKk/NpqzDCV6WDzq0WqCTyLf7lfwmnWVPBqFChFcfbAc6CeEBa/4Tdl7lt6SAAL9yq
+1VtQeM3weYS31Dj7AVUtpuqwrK2Sc97+HUo0oih+240gh1QPOM1vgMTihVDkf4LdnCwDPwt7bf4
PNrmj8Vre6TIRqH4g9oZMDApFVXReAuBDpx/X2MWxenU/ctnjADPliDGARo4VnA6XSSSlEdktYa2
OHTQc2mIH7pZ5ks/pl9JMjUCIzBwK6j15aAiXdJ2dMajDrVOsznIM5WAnhJgflkykUvpxfqQV1Ra
y/xhlEUcScJ71nCL/ynAttJMICw7DhtYCAr8Lb/Eqan9Ns9Hclt8CX8vqz39/ViXP8pXoyZriSGD
qEK934tMWTpWjvflVRhHr4tXB4wocvofjCK9sA+xVpzRRiYIfgHxvlaPu7481zh1sGW09puVEHJv
xsxfz3+ld1AVXB84YuAWV7yu/CVYGG9W4z0elf+XKYUjRjaNGyvDOj/DX+WbEdg7wL1VOCaiKj2h
OPPMwyKgmJQ9OKlwaO8nakBmvdqyEGGqePC2GLBXZ9xItIdgQiHr4A8fk7Y35oTy2n0SoR5/OaJ+
eLFw6u6TQTPpnCt+GI8jNpXejlq/oYf7JeG2lehta00ARSuRaetMGT7s+1wwN9YbJC4Byl+l6W8y
74OVVx4O+brnH7xk4RidYtEl4w41uUCxKUQga3HEh4Y/NP0nrJawSYFdNI2ctO2BDCaHegb4vqCK
85rDxsnXxZGOysarFcA0A/GJKkLnpaZkkUviP2Ew/f69ahwUEv4c1CskzcXYFc4crzKwJ4XrqlL6
gtafdr5P9ZJJbQ4D6UF5f5SIxHV8UuOjcRI3fpf4Q4ouKh65T+RK0j6efd6SX5ycK4s0vc46qnJB
PT9gFf5PsiMaJ7xlh5BcoV5ExMuqPtUWZaMs7Wm/o/9T8cwwfNNSPK1jO9TbAA5FC0RQwDWBGs6e
yVGhyeJ2ZhnowKKp1ZfiIvB5yfmTgP05uCEG7k3R1u91ocXFoDnFqMzoYLDDarwbYTrmVIUFQd24
TB7iFRtrGjE4LxaJdTrLJ0MOFtgWSf4HXojugVA6RKCjMbDX5KkhkAV2BreGrBfEArEq/E6mkXhZ
B5DK62dX2AnVxvuI3ZEo50Q98E2Ti1hFmNYyGNGtBNpH5Y9QPEOYVGxtakXDwK6rzzXWqAFi6H8b
mquhUvYwVgOVKilOgTQ0mf0hYMWzleNEbk6vgsztUt7zSxNeT4olRNN0sL2HLEeDZwOi93jYWgJb
UQMbfT1Hy+T4+DO3qSaBVJU65zdb/ySPT4NQib4b4/fMqXYmKRRs0JriknNjEu35XWdeoiFanfLZ
l9JqzTr92UxXXDN73BhoHRamBY090luYvtbzlfkOwsKOMGPSG0HWR/4hSJgXHsIgbU3VTm7EvpwL
YjuYnKo8efB6I+JCwpZfz8tWEltQYUS7ekI+BbpdmKtHTgRRf4TouFOhzvMUBsR2KmAml7k8US8Z
D9VdhQB8MMo06aWNXJ3ZntkNR3OLCYlvbYwwwHX5xV8Y5k4GkDE2eIjhZ0SPnxwhHkZc7jfvhmyT
Hqbk7Au8I4D/lqmllwr7h1H1YXPmTYwxLOHOCIzia9P0P8vQRBYPY/Csk0R8RQL9pZylWOQKw3+6
euJJVS2HBm/P6v03GO3weBSt2572Txl6nvJ+OJFhFnSJOdN401AjA7EK5sKYO5f0rg2tOs+I5C9R
r6jUVyt7dK/JfARKHLmRWFLV6kJx9Rgyj+fOcRMttEML2EXi9HhKJqWBKxDM+eyzBbgIjKGNxlVI
GVtDguQ3Yle4qf4P1S70T2gc8WXZGDZ9o4HUtULpSVaNrRsJfFaiLy9XXBIJrJKePOMn83NWFFfr
kAJa/RaReePPk2tlfkh0pl0YB7jpP39uBXb+dCgG4rZub+ZoRamwTMroPiRNdOR9qBZ2pEcic8Z/
JCxWHOBmdvWYrFpXLJ4v+PF3a6AB9XwcOV6I6IeW1wT2iBViidjj9sW3L/OIeqDVgnRrxuoAbT+l
o1U64JnsoNGGO2Hl9kCutKGG44HQthapfhNXorUhUvzzyfX421Tjg3LevXkyjLe2a2O9pHBIDd0p
CzqvUlwI/rX8kpKDmSWFHxFTzG2LcTVapIGou9AllKFoPm9l95JBqKymLieLHTHAyIbMQpHc9sAM
mm19y0fTArOC3K9wLLhOMhpOYkFgAdsiC4gVC4mSZ8KyAPZuhi+8xtKLMiEV/t9OeLzzc7sGbwvd
EN2RKF9bGrz1GmHP9BVfXRX4eSALzXB8SuSXmzAejFFYoWQp6GKCK6u1bcsnqd4kfMsz507eJNru
Q/RTsgNJNhOtROv9YDOF3Ym9c20D3veeI0sNB9KGzn3KzpL5aausxy/AG22LMBNEyRVBlnuEDOtg
TvD+ypg0ug8Hk8V8j4VHPCJl5t/cVKyVnZmEX4/OVDPPhfOlUoETLXWH6VHjsgdjp3FAbUOopn/Z
U7hImULiv5vgIAnzeIarPoWtpqFf0wYL+BUt8Zs0OANj/M50S8ObA1egLaqm/n6yBoLBKJGd6ywu
74iovu63OO+EQrQyuvnXnJhDqzJc4IfQFRXWC1hRRakv0ifHu7MJkICw989ml1qy9Zhk+wpu2aad
EgzOOiHmCNMoMTrnrTqc1UOOyv6WIqKmUyLFvMLDOoLnC5WAwWk2vbEZ1odbGVBNWPstMbf+bzZ1
XOpRIhZmLRICfBQRPKM+MwwdkLdss53EAAMGYX0Z4v/QDM88PaIP2iwaxvkhIkCAgqUSuHb7/sN1
p4cBUe74MqqlnX+qu+4wk1brgl8QBetsV4NHGcFSgwtSmIP2omlpAj1DPaxyFRKryxv4k8InsvX0
ass7QyC8iKWKdQQS2bBxvHGCTO5MmvvhYlWtDd9/7Rf+aFy9fzIUgSVzk0WMGWIgQ77padOUpBfB
RAHHq1mV4oW8SI391uq9FDaOyS7aLRvJ4khUvWOqV08Epzl7vFOnis0haMTGSyWlTbqLsTAshpV3
WyzubuY0U8ckqp8b9yGu1azF9ok1f5d+8eI0pXq1HRdPPBAMtiuTFuC92kEUbvHFAuklXYogoKJz
NdUm53QgMmG9GU9eiqm5S1OS4zGy3rLSAK5qVARt5K8A742TieZakj6zHH+t+Rh6MjBkxkvWJcW7
k9n2LW8ECrryLybC0XtCjCLaemxwUbFxAgQMGUN1YEjA+VKl8T0z+HPNc0LfJ765loCyAX76Y1bn
dr17x4fCLe+77ly24FBDhtjSjQYVDWEyfUOVDRXipPA4BN1jKJ+OHSueXrDoYH9aQUFJgN0dwYSo
ciorn+5ndjdtUWq18zPg21dL8mY11LMx8so/rRLW2Un/HX/AaquxoMci6tHiKC8P3kIFQ/a7x23u
dvFGK4xnU2Ho0tI870zWiD0wPSStqr3/L8K1Kp/liRQyD9eR13lXwkt8TgoMqRZSdBJp5jFSLlab
98xdbRoDyv2udUhvKCxho2gE3qUVNr0o0ENtpbm/pBr9yHyuTbMLVLAbL45sV1cXwDpi8TvJtlk/
+Ku1h01cmz+1q75EywO3sgyhYR/lKje/6nQK9vy7XVTgzlbq8t78l3M+SZ/oGNlMN7tW+dkswmcg
JDtmLSz7EjDDMheqTxGDSMF78Z5zoPsdiZu+w1pCFSZwuBm5JMo3ZIjWDIYstRclcjxr+9nuiM1c
YImiQqhN3filV9xTEom2mCcOXFGhCIvTXie6/NVjqW7rbqM6KySvRLwPdTxVIce3xggwpDm+HRBO
cBt281Wj0++LAa+XVb8Lr4usWtfixq5kVwfzVpkbLyWGP0s1GytgDz92jzF+ncmSZ/BNrLcKeLnU
nnJbA9Ixga7BIlD4bZE6iau+4NmpHLfL4vBrxAM/H5Uhnnc3pH+wocs+Ep4hV+MKOe1zCASQdbyJ
moVR59tPTo8vDJvJ3WQKscyn7XjLs7kDympqyQqKYhEmFJIjafN9Hgf0G5RjkGsuMcRsqS8n3ull
yf6Cy9R8kdkgjyn59fZWm3IFnhjH+UCSzZTndQLYD7kgO7CCkvEntV8IxlcPCV7nEi4k/GQ2/KoF
H19KUT+7f0fRIAH/d3rWfiAWZ/bjsHPjMO41078yXvvEI25UnNrXRRwVft2qbJYSIKmv2lWi5Lj0
a9RAw5QzufDMoOuCBH5chSMZtMh2h7whqzFmbgLqu7O3aH46J/dxEgu3+MLXwHnep7dQwxQvWl5i
mMEddNNmNO4cHVQoVJA/iS9B7Zdw7qui7wFMfJbkdYh1ASoLm1L8HlrU6QPDzA1USfBaY/1XEAlx
Eofb+GrKuBkwZe8CaUwou9sYmSiLPlDfPseFilzKhMifb530yINWWl54nuPZ4kSzWdUv05fAal60
auQnmowwTm/iM5VObR39bpMCEh2i3vn6FQkzVHRXSJD9xlegzSkoekFPNlWGlPffI4Qg1xrW3w0Q
dJMawMzhnPbup+KuiRa173oB7lcVN830Kr7t6sthgPBex9sdLY+RM9lVnyGJDRd/hbgE6yqVdmJP
fT+g+/tvlDT6in0rDUnFdPc8Jq2dAjFFKVZB9qW8La8GIlR9CPVm8V/dXykt9At9yGfIrOc2YmFZ
ZLULhC1+qQ1yA+uFQ00nlCfoNn5wSGXyXbpaf5Xk+mHrkxd8kTJHg2nCGc49bRIfYggS0A64fhDp
r4JL3xEHVl27kO52KJEN2yc1yyOHMSmgUBSMepPdEC53JgmhztKa138UMLlN3ldl/yWjOaMqJZ3z
l1n6Gvht3i9UUDeIF5LKGPZtiUY9qlCG1jNw0I3bP//H188nBLPIbkzoUIlYjK2IgK0Bfzl5UgBU
G1Z+t5J+JLuskvQL1XdTWGXvcc1/6/tnMAwhnxN6rISOX16r2hu3KTTT4zvUFeGo9L72qkZgU1go
wmos8ZuDDTSemyvOuC0BEvL9bhtGNrVDWXI9yf2D3EP4L5hHaFYbEvnOm9EhcEY3+Nzy94Wc2qVk
Zp84BJ9/vzudB1WUAnjb+8Ua+pRczTbqKKZCMhyWY9aEK4csCudAiQvxCT76N1APtRzNflY9Jdn7
Rt+hgoAkVb0xR4Oa3VuzKY0Xg80hcFIUT8jSoday0LgreooLoJ6SSjBNfFk/hVnSiefsjt0JOC+N
4i+Z+9Q59MsT8wy3fSQ+NOKxglo2BcCFvDo+hyp63uy1XqOIYfBofCeUwi/AeIN8ylbBs0bYFW8W
n9XsOaYi3q4o8Yv8c4ftOClC56kpq63feoNZMg9CoWweu5OPWyiDNOm4Shyd/2wcPjxOgYGxrwM4
23bjjsJEEWbmifcla/T8mzoK0+Ek3XRRWfydw8HUQ6PagS9SVfVByV1VqXPNpDKYEf9TgQ4s7gWU
giXQorugWmPH7fa4auTibtgiQI3LhXTxaGtvCxDBxlZOZxzq8rMkfRhr3iz+a+7OYnb2QDy4A3s7
qwrrtxexS/eXmj3srIer21SLwLq9cihvPHNd/fb1AhED3OVk4njcxIkrVlQ+VDxng6646IOtW7aV
ey+KdxnDmKfWVY2Flfst5ZkCk4p9S9gpeYKkkvyT2Np1IwjUCbW/4kqLYxMU9zu5ULC/gNn+EWD4
2DqLPZTqAEj7JYK/e5TWz3JeJDPdaLn3Z83KHbtWPgqdr24KLuT2Q6L0LDOYzMsHZPJr3tnepFZW
1GU/3/dlbFgz6YItousagQPj7YMo5NbYcsr3xspw+cxSqrADsN0IuIRZTuoMcIsKW8/PRBpdiPuC
I/aIdEhuA6hOp558u3qs5qNuF0rUbD5o9rY+8dy2dtKADfmouxXWuDwJrvLVW95M6B+TVmg0pPdC
kd27QsQfsA3iwlyBjaibnI/glgoUvTt7Kl36O4QF5kLoqFeUgqD3KWagj0MbK83h2JCZp5F0V/av
F+6NEAcrWfvOjrbEqmVHxypegsaghoEj494MONJ+dlqfnT+79Ov3w8rPYBwtiIyhdLWEnkl7p8AG
8Aij3Xkve0qf7J9MHjq/+15huy7N1Ht2cest6Bm2FafEJJiZyriNzjc8DBQEv1DOX02KFQijHs7E
OMbKoIcz6lwjc2nWs0NupuYbUqrjnaThfGOxImeD+p/8+Zz/VyUMUkjWwNAIWBEBV8RWpabMEC0d
58HJhjvvCw/GrrPGMIOkXj09+g+/LL69y79882kvFIwK2hJUKvb27iSS/OzAFx4le/7IeRWmw80F
7aQZO27fzC9CWT+wgFhHBBik1JYFffFuj9eH9mHweaDTY8DfG3YFi8ltXqXNa/KKrs9ZI9rHuvFP
AV/zMaXhqeYrLbpLeTX9inFgvQ5eF8kHpAcGHan5nLpaRHf0V5BkAv0Dp/VazsCSeD3uV463BJ27
OUorSO8+x5fffKrUgkx7wog+yu89gvEjre8cWoKQp9MY5+JHl7L7zRFQg99abRxm3kDzlJXC8WPJ
F5MZ2IAa3smP/KrGGe9v8PO2YQSXCj1sJsb75kdC7Vkpyd7cxjfTu/cSqopUpRj2U09UX0pWGE86
fb8U0niUfW7KZBaLVsUPK5ALw1Jxnfl4i/ybIZnu24sTN/oR+7L5NGkvgcFsm8oHYgGcdLOuVdno
GJE/O9Vos52rZdgkn/fx2c78O4n700uIPCAL3Dlkua1CjsY4+1KCYwBYOWZgfEHcsbwdG9MVUsxi
z29SuQPl1bxxYrh7RbbtFu6sBlU/Vkb5TDiQIpy5rqBBEuqyE7rsrp1Qn1amhJs8KY7+HCv3t8+/
/AGzq7YVgtlZcj4NnCyJ0CzQ/7tSRZqyKDGpd7VQ/IY4nvSibFs+M1i/4hZTXbUtamH+SO6Rfks2
Okw1s1TSCNCTLO2aUoI6LsfESMBVJfjzKdxDCNoRzmJOGGVe8P3LybjA3tQ2pQ+9UsbxgqFXJ58j
e3KZ4QJ9qAatJ4IBCFDt2vv/Es8PhhdmzMoi6KjxjP9Bfl0j/K2FCddojz+TRqzHZNvfo41TspFG
+xKSTOI7gOKyKlnXXitfk0KgdPr5s/JlmSquPKJzf5WFVK961yni6ak/TqC/nJYuNZM+W+8Z9iPj
UrICPB/PE1c8M65XiFyGhDkzSNncYkcDj+mi/m7/nlXg+i9ZR9M44oA6GhtQisrFWp1IwMPeKsXm
zbOYYBzZCBI0aNh3Yg1SUZ2SsO3ff7jU9k1Pd8S8VXNGWvI5NNRYrkDYTe0ekSiVtiTI6CK0e0oY
B4GaPJEz8gZcEVGQL548sxunPAT6F3NwcofG41vZ51WibTZKfVqoD5DVYM63uajbvYYzorijX7U+
p6/zQPq+W9O5fRywr6cHGz6jTlnT+N4cDdfAF0FwkhgIoy9QjWjz7eEQEr3xY1sbvD/a2g9kdxYE
QtxTLJ1iZkgDGSDDzqGu/moC9xbMiRK6zUXe4zPWUOyHQbbTlTmEtDlHUYE888nbX5/M0/8U2wsC
Dv6RU0PhZ9drgiBZwQhkbFWuxl8V3PG8HORZSFs51TkVXvCa4p9je2jChMlM/H+QoNJ6t1iihI+S
PKJaczm2wTQzNC+k56Drsb4HfeD1kiyu3Nyp0Hiel6gv7lXSs9yhXYQWHDiPgkGBA0gkRi1jvMch
SRRrR+KseD+wqq0uCusE0GP1QgIKxFGQi5Dh6hS24f0h1mLQ6ECOa6hNd2BjC33uCSuJkg3IjM93
hT2JqizDGlo+6FAqj7Azo1ccEa35aL6M20/76JZDzMiHfauoHJc5aqF7h9doPe2g3ZGiPSUGE9nR
sayFbnb+MeDErd/DsVNNdK6nF8cUefJdu4u7LyNM+VomPBrVn63eMlkCUOuOVuFkW5KMOlci96IT
erVN8MhvrCiUEQvk7nuqEIPZFL40ZCzKmcwhhZaWyMKAV6zKmAwlFhhRHtGrwv+4K3vdCqeebQdk
bXfIitYHrnYTuZ4oJoF9ZLAyQRLRTuSVrwFNjU/gicpJArQUVT44ZVjCctupCe0lThkFCgNSeAlM
fyBc5Uq1a5L954PLS9/j1qmhGmPy3E7FUg6OprnHHzfEJUi35xxDExX7T0IIbbQAvF6V8kpKrWrR
7ihQ1lIBTkacqdgYO72VRwxQpAp7YAWzocXqvaXCJa310x6Col1MoU9y/q3PAu3Cdlvur2ouU0IW
Gp82wamhiUuBSBBdbCyudLSfKoBEbmDrdrDxJS48SLlfYzLltdKxSGTh3nZhvtLzrdGfxgiWsR8P
i5HlKyCBw++87CAhuPREPI489VyoQ3N/yfgBdS5AkbAM6KS1yj+GESUx89T+awJGhWRrQi99V0Nz
LyORPJBqKvJFxG0nuFGZH+GGfPHnpdusB2nzSKFQlnTg9qIw8htcsQp7uXyFzSxwirzjP5+agPEC
hccuQw1wRrHLu4eHKhE5hHohous45MPpH9NyFUA4fBliVZBrp/NHJtU6v85gqkl/ObFB3PSNCWRx
9UqYOx5MqlyHKYxPsPfJuuH0ajLahQY1EiNrbQhAKhAzgJr+Cq5nPxJF3cQn64z5eQtzMYYIGI/r
h03cNJVTqVLZVWe11Ixr0UsorKssz4qNX4xD837Ow0VyxLKvAfo19NVfuVOY/Od6AY1qyL+Qmjdj
ElUXET0tv7tDtK8KKDDD7NRCalZnCMhgFspYJI0o+sPT+n4jckSyaq3k3bEHHT5l1MeWJHxIjo0x
Xheqw460Q2sOP2u9Lwi1qYs6N6zLos03QC8VwHAPQnNiQIiWdhLx+faRjwHbm+fCMWcRka0ykM75
gjxKrai+N0DfOAfxNzxL+Var77x0CpFx3ZZHcd7jx3ESkTcvbRRRlZRmtEI+klTs2Y8pdQoLt7e/
Ceq0BVDKl8gFnPTZkX7bQ7iKTdueG/EGsgMKmbC7wSHteuxuY1TR2rXwYG+fT9BV9yt9P6qOq3dJ
tUquOxz2UD9YmwJ/rxBBop4DmD0ybbuB9YM0BaXjQqSouXnn0Hld2PoxaiwPZK/zx44V9xFK/GsA
UUH7k8cfl2szPvUGFSSpE+vezfS17QozoW2t4h1EOUQDNgNyGWr1gH5jukY9xDBCFxoIy9ST1+wm
s4Cyye30qnSYLRZbbWXhDWrdjSiRKOfQ+D7idAjyvpW1Fwpxb2VsOK0PZf/HQJRYwqSa5H3xNWOl
lEqxA0arYMjCN05t3RjwzszeM1H2jz92GU/M5aaPJrnXcOLmOOQuWreXe1LrwZ9nzZ30HC940IMG
RChyRd7HgWH5K0X43YyX7bBbddfN0/vMgtjbutJJ5BXTWdTjm3B36G7/PTGGpMusNsfT0XK10b6H
jg9LSIc5jAScwUCVQ5mBa1iV67KwYXY3TOjk/2ghmeVzxE3NAQe0F6na24rPjRHe9fhhZryGxOcm
D29ghgInQZRYeaKE7jqpgSVuicrTEda8UM36hfcJTQ1u9TSX5aS1w+j4uQ7dJoLFEKu248+4VUYJ
nW9H1OpHvP/J0G8OAm80lpWaKftYC6+txqcBbpOAqpOxAVoqZcxMc12P88zdGuyjEnWg+FjSZxvz
24U9/bxQtlPJ0Pxn23eLFYsSp49iwHYvUhR+BD6/6KUHCXGauZg5DNoXR7t1gghg2XAhG+rb1+Ug
3EjEOzB/SrDsOAQSv/Pmr8N+yXfUUOcu0lXQwSxsMjLsu7zeCZbxqXJDbb8P3xn3lLObbSKmkb0Y
jpuMO/cM9FqZ8BNXU6VOpvs3DUl+uWbRxsFqPIS8UYgKxxQNaTvC6bDGvL6/V9hSL73lRlcd/lfs
vzGaKRG9lsNiGPyx15I7AhjSAuYUHmFwfMRMpaUAPPnpjwTIfG4eicLFOiYXlse104EJRJVR4Jqu
2SMJ2z8Vpq1y05VZ8RRO5ZImbxBtqrGTUzLb9XjbfpIblLpPDmO3M76Edq/l9BCmut1Nw9JWjEdV
FsC/UhksD2ULUUKCLMtyhEaJUYT7l5myE1UgHsKud+L0DRkKmAu5O4LF+3E8NQ8juj5xpTXhdixC
+8CbWf1vL07B47fmYzwrTQtFV65gvfI7zx+A94oKKr/9ANpKBoMuvau1FZM+KbYemyq5zgauRkSt
gp8yBI7TMjtKWroPnEicdsNApwxssSMhZlfnuA+8XGMKgF1IeE8+IvPQmcYUlQsCyDdmxrFC/kPF
wRVskjBF5uqx2vEHZeQQkMiYoaCM7fK5QaW2NUcd3X2lK+unvm+w5bL2+MrZGYW9LEVT5S6XX8l4
u5f2RSyBnDtMr/N96AO32U5MLXdeXxVFkzsjPdQCwMPiOJWP4Q5Q+Iu83yOqrHYuaDPmuP/lzLde
Zwj5oMetG3L+8EHIviK5RHH8tWCa4Mk0vMrf6ZCSjy/1WRTKfKfi9/Acnjwtayj0SJ3CzC5jnJlv
5uaL06tfRJP5CNScXihObDYrFjDQsdvwWcgXBBb2uABiiIJnJX5WcFYHKmmtV0ZyM+Rb3q7vmPRC
R5VtkeG4b/GlkNlD4aLHc7Aj36KEBCAYwyEzXF4jcuQ5MAzI5mkmT/3Wm5p7vkT2jq35gZTWaJta
+cpEf55eS+2pax/In1OMy6N6pGtlVOpE4azAMMFEkWBjlfHPxNK5er2MaLfIVyj/UmehT6eqCAI4
KAGoe+4yk9HriBpe6Nwc7bcnzf9ifp8X9M+79l/JmnV6Mvws4o19vET1vrEh0rQmrvOkw2VQFH99
s4AJsyDAKcAyJKcREeLqP6yWK1QlZ9brYomBDmPaMDywwl3JiUEzbsWaWZsuZ9f74MAI4MKoovOb
rcDdQQ86sqMyhpNLwPtUQ5ZtGre4CvVu0fclMmiWetUJV5hxm6qDUCB+E+qljQ3C3vWhJrFXIYUi
LDtwpImO7DJojdNQHF71ImrMAgYvxRA9+UFhlkPxUAuvhrypUIJtksasKFnrzWvVC5lyODr8N/zG
M/I5C7eCOjFqvbiLwH/sBHaExfYa33DbUC0ey3erKsPR5bklKYVV6wcy7vhaunFdBE5UDOm5CNnR
kc9dy+sKqtccB6jgel6IRbNI/tBkPOH1DOIQbtKWOF40zD7l0m9WDXdPLyHsD8cutwDtTOW8hqFR
ycgRAv4QwhHjhXAjoE9sGDSwfawS2U0DPa5qQXk1ORuU5s8L6KWipx2JNSIjDbfXZQ/2rpQwdjR3
sq48KtuEY9HQZe8LZzKykfNeujkCRYcfkrrFDGu+Ry7VvDu5KWvneBBgHaqJZY9ecvphUVicG0H2
6h01k6DVFD7+ggs+qoTJkAxkdXTGg5eyyUy9+BodI4Z8C2peZ1i/OMdICaNkGFBWEKTkZrS1HlNI
+dt3/zXNQVgcnU6Puy7cHkgJ1OpvZgbCo/0hpbH+ShEzF1J1Zo3U9Jlsg7PH4sJCICVhC7JjNs0h
ns4+d1+VvzkO5oL//kgbAE0bM4Fd0WN/M0RE2/UhGgSDSc45GVoGo/B5oeBZQty99IVWmI1G5cOS
jCQj1v1hrCqAu8YlzSDf2AO8xE3rKrRPZA1apz2gGe+8y1rIV7A1YLW1FuJpyUZp7VBIdtjNDZNF
pGuBG03Y1SUqNrGqoqYEjHLZdrgPPewdKBf61RyhxYstH85zhiqM60iYRnnW4gv4V+YvFJqsO/Qk
3S0F/mMW18fyggnzhtSnQhhquOpJWQhp4GivXDleb1CT7P35SJmRh5hCtoPSSWVH1pnlbnTqJnzt
vZrOg65RTVHsYKIOUpblrqFBQeG2bZUXa3FARvGjoAlbrmQmspjr25SrXEFOUk8J8PVKuLm1FrPE
jJzxvOhYr7zaPBSbJueulq8yqO3SAXHBQkbyaQrKmuQO7JBDTHqHGZ1zq9yLVwAfeT8PlqazxqMO
146tDxkBQciQjAZU9j/sBww6ePb7G34SKcvsspoSe0i5VQG4SchUvgfH+qKMaWSs8pm49lM3/OYG
ULRowBTm9BEn/zAh8NlXkpfr1QY7eZwenRP5b9/ABsv8UVuKnCaBf9aj5B2HJzp5ZTkTs7y8Bxdi
UbZ4b3sXuj/kDO7kMmfnvvwit1BPjALht/ys/KUnH1Ssq6hIWwhxfMVr8Ss/XJYRptD1qnPn2QP5
vzT1UThE795vjm8Oyzd7T/ApK6FgLhUCR3lQpPCFsi8PPw9qSSgbDd8akspEETWzQMRc8Jugh8Fh
wqnMtX43giZGBmNsuHSlBKqrYGXwLZo/7D9VX1c/egGvZkxAq9IzVsYgFYyHctx52S92fzz9ymrL
sV/GZ8uybc10cz2VuJCfcTuF4flIsK2xHQoxgIxJ2zeLaQNlDz7J2KHUiWvtiLmXQjhZKi4R4hTm
0qsgaYlNgyZOTAsBYC7lqjIq3gxKZ/MrHS5c7cTkG1YMzuOASKv4/9OMPIEsIGvSpyb680Y9hLga
kzugevy2FyAxUYgjerrOlVhfj6NiLGnpA2Qpp12oWqmHqeGkpYqsWcAlQ69mtuczTyqVcb31R0aP
I3Rl+iRMlM2emiUqh4lSm9ZembgDMcdCj2HcHGvIWqaGYgrlFV1wObOl/blPwpFXKObU2kYcU0L1
3MwDtF5Bb8wHB+ZsUAxXZx1oVx9mLl+MkEulzG5JEnhIAajaBsN6YG5rcwCYJbKvXW2c+oq88KVy
phrBMTr6/IlVavZr3TLy8W/RJaNSS6r2pbkEEQPW+X2sNGhZbHs3gGCnFMzNl/l06QXbFgaf6yKY
0tn6FC222+Z2og41dGuF4AWFrgpOHWYVOQ71Z8mv4W2u72Ve60Y84gExKtjUhdO/RiVuRk2LG2qX
NxJAqtRpaMIkEaxXzoiKNw/JaULzKCeMuyQnFiqA70A4WVp1UrOHFz7BCcEPnh4fF748aOhUt74h
xzdJSKGjXlv/UWNQUtCcZsuNg1B2TRLcFh37hu2sGTPKlcJ8gM/qrXJHqc6T1PmRTgcXBU140BaH
AIi9MAl8nQYZrUPUac/MY8G7WYkm59wrOL8ybg3TdY4aYpfAon4wVsp13bfLW721L7ff38ed+hr+
s7N7ItmcSzm/f47ss+LlDaBnAWj+nwFpoq9JEpRojd2xUuhbVRUMWx16oPl2yUIR1v47xfEssR9X
32uh/amEjNFS9/t2sebKdsJTgSWMaWKtmYR6RJWlPeqkSBRMebO12mdSrlprevx9r9qkWn2KEekf
C76gpqAis0hAhgGq1Z1hisu7elCC1WIcd7cSOvh0lV4Bi4H1D5/hGOFZs5ivByJiu055f0QDPr1i
9li9JdfzKIjma0yG0MGfEdHbQJC/VFhkAou7c9EWkzo7FiO7hbKpuoymJ5R1CkkZ1Mlwtl/h4T4g
huXPMP0DWWTv+CjuUpBhhpdrC7LgVldaMvyrtBYuRBWnQtieUJZt0HnV8pKI8Cuku/U0LXfwiWwV
AZhu65u13A5BPe1ojW52ltG8jkPokUsUdLOAE8CH3x8rX2Uxnadzu8mpy/yc/WCUp49YPN2Zm0GU
phUjJdzJDxaJBoXd7VRMrGE7/M0M0zCAZjZTnABUs6D0ZaMAJt/o5kS6cUBYzuKnguUVCZQuR7sh
Va929r/HdEhNTbhcCkbPu8fu+00vnafxSV4u+WqUaND5dB3wn0JMxg3jnjJ35NE88IrSqkJKZi8q
i/TSM/FfMLiK/Ch8yKLBROcF/DzVWEBXLauOfCl2w7UGIOa4wc5lL4kC7aR5lEOzyIN8dWzZAtmG
3GOQoLVI+QRWjkGUQW+F7O1AIKXVgR3X/LUlzGv6zxWhRWuPd14PXlb+TCpXJFg38GaydeTp2zvA
os58mKK3a0MIWkiwp9xvD0FePPcFssASGaTTCkoYLxfm0bGZbDTeEz5Qkn6zId7saJL2fOwjsF6P
b52U8S4QlIC6NROm3pRibiphVTOT9Sa1EkqXwr56n/BX1B36TUjKlL3o8wAE/Qu+q18XnNSXinQq
WX4dFfEn1wHsPva5KS1hhg/6aSVLWrbP3Wsc3Cxo3TXPR+lcOooewcxbZhw7ky4mZ/f0lFUzZ/ju
um34yCzic9q3boQ/Jlq4J+uUwbxiGiwi12N6JK8X0GnbTII9IsN14E1vGlr8V4x0usvZ870dZTAr
fRmnfZVhsJv/yMwY1m4BjdjUA00CU4LOl9cBhNZTVYz1KDKpSD+9r7HoooakAIrVbwp6bNGaDNhc
pDoek5udpJPjljZn4f93VPSTNS/W7GwVoH22cXdKhdGqqbjqT9Gadi321anmcBnvzG2LWyoIYPrt
+Lan26+oq0T2E12HXOLNJNSW9ZfdRqHZ40hkjZxfnIzOegXGOTvpGha2KDlM0Fa04FCi4Z324R68
N0XxZHMwl66hB9OpSnL8xCe3TXg6G+spqWvEt8GAjDrCSKBD7zhFZa8XV5Jl++sJF+9cISOfJvXq
yonisF1eKvQqF2k9gPHDPj0aP9OD1WvjrXrlLlsxlM2HZw82xA1W0KjackWX2EgumypSGS5rhuVG
FtwjbV/CkzM3fjkQ4gzlZ+vcujz8rA5E3rr5St+4fiSQ7EW9bfznuaORNUKEKCJF3Kc/UvjxtGPU
OCVc5n7gGSyqTxMKRNmre7MyqobSZVvKThjmQez9IT4+YNH9WmpO2O1pUBeSeyQLU+7FJatw5lin
h3BAxXK7JHd6TUgOk1S2TCcJ4uKbEDYgNHrWrZxgqVbQkP8K5YOSGf97tNnn5c0w/kigyVeqiHOp
hQF1dz5wu266eIei3BcTNLmeKfiYBCai+aCSaw7gUmCO+1sHlqF14amzF1kcsx2XGb2OFfzshygf
geRo0syeJUGA3cG+Tuw00JNY/HpOUlfxrNG8tDiEmzLNsw/XTpAT/UG+5Ws7IklSs7GN3oOKqJqu
cgVuVWhjNeoo4OKxkZd4fR9yTTKsTnc1ChmW6cpGJc4TeQNTYeZONScnW/TM9ja44JGszPlM1E5p
+FF9SemXbQg64urz95QQijNfHVgNnXvevE+dExbNNnxgUHKmXKjennV22Bzhhp98cikYKeqvGOLQ
weNEHEEi77cJdj2AACNfMdvUlbw6Vqy2KiI3kRcg/fTSxu3QdXZDRyMbYMz0QWGj9NHkYL67N+G3
QcFN+TiOfWCeqgR1Jk1qFIZ0K76h1Sy7shhIJ0HqRBdmR1rzyWlO/JUlRNNAGl/loMALsobX4QrA
aygXwxpK7kVpx/BqGeHNij5Vrg30AKN3g1BbVSMFAwU9mn9Y+pxSzxgooZZg9P5JUR6z7HxCkqjk
jQkTzEcv2fYanimcxxC0C9A2MRkEapNDk5t2YLvkXLnajKCe2dtLjIhLNjIaFMNum3mthIwlgfve
Xcl8+ZImuRUK2YMjjbPdmvxbBJw0k5WfyYBiTyWf3rWUic3f/EYYDVgUZjGtCsgtLi78UeumETTB
y6TAHwOOZZgheQTUOHr7O8mcA6e+7pT4CvGF2q4+vablrD9zgW6zMeTI0x/WvO5nkY2ScNFTKIff
R52RFv6jdcMqwnYaIVV+jz1iRj+EQBqR2N3RQYASkK4QaIFw962G0Hvk8D8kXn8+u6JlLhkkz9Nt
QaIocjoSbj3fNFtGHfHykscdJBH8xBhGAfEFTxgn0W43IsjQ3K8PN371Hi4W33kM9qjNaDrkghVR
sYqNcB9YI61v4fpxMkT4204VmY7iNd6Fnf1SzS2rlHehdcWyYMui8qhmCAZtediwxyNKgNq9iIJ2
st3ODM+5HXPgWuApOJOH66WGRABpAKsC1mQ1fCIt2ZyvUEZ4Db07b+M8806ZjBlb+Rky9LKlZ1Tv
NZBnZRymhgXYqVbtcV0L3eRJ2QMiTFarwH5LGZBp1VoEiTaIINlydtkRgndFTY74nt7z5zl/6xte
QkT/IKGgtMQAVNRw2L2k9EXiJlPBw4L89dqp7I4So6dqcyp6kMMXK0Q/3rpXtAS0nx+u9AoKZ45V
tBT3fted2YXu/7xbkl7iXmf1v5ctykMmvzqCGTyKaOItkCAEnazsPcclMAWYwch6isnfo02WMP5v
Uls3xNcxH3/zCoLl/eDGDMZHYi7dsXyLFGgJOr5EKrWWVwJ2Uvhc52/BBIrQKVCs8kGTJ09dx5Np
JQRiLX3A6N+1GLfikscCA2GG3TSoD6TE9xxYVHYxgGtYI4oeywZpn4rBKtsvu2FglY2GQig7kZM9
bFGE6zTY0FVcc27IVegI5+vtPNjUcMCklbdMTNVUbQr4U4LnGfRyOZh9bP3UCZ04gL/2MROaQ9fk
oE5o6GsABm3YRg9OdJ0yG4yOcNFMmMQZBvFS9N++V6LgFZES1VfcQpnkbXNLuCHp4BYQIwZRYCgy
CkQYIt6r0Xg5taddZLSeubBfPIaRDmVX5TVi+7WJoKFcnMYn2ZCCNspEfrRLm3rNjw6gHqoW1hRP
xAdYrPXPpPam8LG1hENTP0gg7VrRIxqFuAWMg2QSZ+yk63va7nAvCM6zS+vFjbsK8tkkl5ZOPZOf
6DB/GKLGAkJPtT+F4/2JaqWcqamhOMtKJLSkrKSU6yoVHFVwMhoZC5hSypCdUyUAW4L19W/nh/vZ
Mh3hcoYCL9qqr8KJ1e1aOqDU+Ea8fcF8mVQHWNnknO47KIE0J+2B4J9gzkFOVS0WAkyOHrqOxP9w
JpiQRLUiwAdi/mHCz0UBzqShaAL1NgOX8pIe1X//aQDx1KeNWXcPiOG381MRghKkMIv9dAGcx0EV
3qeZ7HZnD4aYsFn8Tldsz90qyE8da0pHwnEFaxK6Ev1kJmtsjke9ATl2uSSEuKXZplwGvJJda1Jw
JVE10GH6NoY2VqRqNFkEgK4Rr0A1APpY9/dFuE/h8wraGiPl+IIgDIqB76UyrhCyhiv/abqdHV87
pI2/iKt25cpns4hWHunoUVXvBAlRi84NPcHQCibNhgVwm4IZbz+2ROcZyBykNYPaM/dWfylIi+D+
vVsTpEsS7OgUwyOUifVeFZeqC3dVQ3L/rlBUJgtxSACR5vne2yKwjh8fVVGFCBMN+7spjvZW16as
T5DjeXzMeqg7hVN6uIs7kyMUbhtugb4MyL5ojQ2u2DHEWJoVAZHSxV9yzKfHlUZkX2Z3PVXI26pm
EWUGQrECq+e1l+yYRmTx1ruQLb0fZpqzlQ3DkE0MEs956UV3Loq6ab6QkIlOhjjkX/mwLDNpI1OP
Qk/yKLn+OIYNU4iVGm5kk1WFkNXcZbCwdJRvy1mF9+jfPLF4Wa6HHZhzlSGhGuXAyQsAxsTNzViq
BJ/xgc28oQjRsrwftBcpKky8CNN5tMtnqeIuQQQ1NJjrt0UuJ5f79gUSiaiIRp2E6VnRJdzAH52c
xOrzQvmUInZ/JoWWAMFwVsN7Vn/dqQXYtpmOr8Ua8Dk1VPB6cwc2YIYVF/c3p+ZaJgDkoA1NFcGY
+Afw5Vn7dBzvWBxQLzYj1kSMfaiNZPKopgZxPjC4KK59+84Dd/JYUOicwqeOEn1VgQIwFxw1nFw0
sys1yKYDqVW0vWZGK3zRouYZ2eRBY6RaP8x+QH1e1jZalP5G+Wt6Nh5/sJAId59UK/7tp23SZflj
pLYQh+5+ZToNLp77NZz5I8zVPx75n1l6fn7AwPSDepFaTV3r+WzDKYLCL/vydR/hOWueBN5XnGne
BD5UDTQRH6p75vS0OpBSOliPbdtW8GqXPmhw6mIAH4nq1M1sAyC/7HRWwwMD+DjvuvU2TCNQk/SK
L3um7owp3s378NZSUuO3eN8xkXk+0j6kRlUlvBUG0XQqfa7+8C3LeVWHou1M1eSsSrHd8PJOXU+A
EZ/8Q7eVAcp+1hS0o9YC6yiJ1vA278aoZcZ2Qg7LfShGcTLkWDc+p4Vaf/R62Ll8OBMyonozqkaG
7bb8QnsblMVvzKKU+GHh9hPS2L/XPiqIlNqHLSpCqwxEz16GF7Rk9zBr8IU3IrLYUO3at3jrJPR+
0wHhDAE+Z1qOAfbGfQeQc7KZitOgP0eg5zQw86Ggq62dOeweSPy0rqAVyg6AlQ9UDLJ2+vwgKewk
/U8XkPZm4v6Oc0+UrW9C2vy84NnhSSOnf/KAX+jq6snZoFURM6lzU+gmbI+bI7NS10nD6qmM9g2v
Wmd4AmIAZUs8Er2JzcGZKD3A7Johuo1AWUmIeK6V/1Lyw+iXE5PI3lYYM4xqvGvYoj9rSZnffecQ
aRaoFerfLGkV6GTdmcIOu9tg+am6MHYg9R+WiaVOOBiLZavhc4uO3jHokuGppZSOD5gAUSYeoOZi
B4OEFSylXWI5y4FjEEqm3NEslWQwg6dt/LKa0SXZmmGqxgIrXfm00v5KE/x4P6YIHY9F/yaZ94yX
DwtLAKXMVhUOTAw/90yiChBCtLLOlfoXUUS7238c6w2GI4C9R36nl/MEQzQL5/YwvR/39nnL2z88
LgyRNR211wIhv96Lxk7C7WPVIXjBHRgEbvYQDtHVq+/r4y5iBcKL3cEc1F/+bQrq61WMsdYOBVgJ
+/AGzBLwwtz2/TMXW+Vw1K/wdeTAl8g9BVOGOAT8a+T4kf6piv6eiYcbK/WUIQiauf332cXBv+rn
eZzd+7FWV7fuf2tDYgRl6j8zrK6hfKXnMTB2pRqsCthGGda0AHEDpZNbxE0/9sK3KctgtdNHyunx
qNQGjCcPd0CZbQM/EmidmIdTElTgsw14eHp0dFpknTNpWMJh3EdZDaoVXldjNkw7TutphHi41Wjq
cwQ8aha/gSCAIL/JW+yCcPoydg14HfY9y0z2dJTGa9broipr/kxkQAto+01eUp+SeiGa2CYGDWiW
acSS/lKnogbZjHzVqYXYpjgCQMVtiIP4EF/u9y3bkNyUfowDzHcUmOvw4nIr4JesE+imRR8cEm0v
qR85vihF+VPU0T051YGcumqTCzOXSji8OattVRLhLpBGHHa17F7pcpXHZyFYINn2+u1JOrWETgRs
F2uFUebFBWOXnkSPLtW6nq/IYQB4cLNmXv6VeXQiMvVD7BVKYxKgME9rGeBZnYUfKnpsiSsVRhsy
KFZF89rYMcNIFiGgkFyEnZSJNupt8mveyozjY4O+6Yj+upIdLreHpbgoRI7CaoA7kMqPx0umURFW
Rak6MikBKkvoF/gqe9ws+uiz/BFdo3owjr7tGr4pP+j+sIAl16IXlRUOz7TAn1MaRIMkU3ZBhvPw
lcgwJImWOh1Gu15Dtd9IfyqXjm14uAYhywUP+d3qd6/i7X4RmBTC1dArVrtFMcPbwyNSRRBiyMXR
t4Hz28R0MvBQjsCXbAIYgp4/EZYeEAtJn2lpnBBGRGBQrfZLuwysk5ped+G0e3KiW/n0n27FmnDK
Wpy5goJLx999Msv4xkeWTZUZbSLLBtjt89snhy/Cwq0txp6Wru5cEQZNVp4LY5RbLEMvOo8PQUNs
x9XYp5UNp2H4i9c6ew26nEu8vmrdK/tOjJkhvkjmoRNOEiPnc3saMSf7UxIGTPs5OUPDBjbN+6Oc
M7NVtm/lV2sQ2Aj5vM2aRwLR+JGvXDds2rbDCw3zwdO9sTSSmpHXViOX/dpJnMnOksDKxMe9DGDZ
r+uG1E6ETOih4T2CqnLHYledamOzslq5Ag2dj6Td+VAeUHOHcNscHid456iIWjWLB6W4kOpMWqP3
ldI8hn7fZxhY4v3wxQ7MJi+otZeAPjHBK7iAFtY5OFI0qcejGS/ZFLgMfYcFuFFIjAgqnSxCjmNc
S2DMVQMuZB2hPO76oPr1TyHQbUOeekqJ50ykDHFN+X+QlQp6ium77+7dXIgpvHWAPgvcoZxpjV4L
c2LCCfXQm5XbTT3Ki85P05PJFHhAFmJAA4FTChfT4fq4r2rwJjuwyEOZgrQFlA7MYGfSjI5YO/3k
z50keRlyUiBYNpzf/gvfnEPo+fx07l87QB3R/QAH9HB+g6CabHlYJTCtxhGPjRaHrQn+aVonWJ5e
DCwRmfT18Tp1mtzCPIdG8R/xhu66XxKEj4adOLT476/8wb/daxhik+QFDr+7C4PBQ+JgfORIS7kk
M2SeUNyRshiSO+Dkh6EmwWqv/IBV2cqjFJfcd887cZQ5mpR0qVpi4WHW/JkZZifWfI14S1gJhXIV
4MdZvhQwbxVeHNarixx+6EXCCQ1Sclfa54rs/imPQ2jGqGBSfqv7BYB9Mqo/+sGQKuFnTJMQSd2W
6HU/SOCR5JR88isLf8p6TMoV1sm23qtalR0pEppPBXiGqQ1zUdW13aolP7kPLpbZjYv6+/44gKq6
Mv9lXCuRgVlUUXDgilpbl/3gL3qOy0q7mFSr1EfBjmQomrDo2Zn2kJP8opmD+mDj/vzyFFBVu2d0
2aEmPaegjiTyA4vF19MjwgtDlFEmy6pwtL7VKzaut5jJVGFz92AY1E7WYcKUzWQoj8svCFSfxfHx
ML9ogt3tKCPwi7BsRQRaD75jmOr2AEuj0QdhL50MAgKrbqh5pKq/wtOzKgLWbPSrhDMYWwEsvHs9
PPyYgLpLaY7RKMpY+tl9mA2IXnxae0K4qR9RxOsKYmLOACEuxWKOS6CtjcsU4uoCEWzEkxK5Bx8T
Qa84Vy0uIzClI+ZbeVOUoJetYMnzLxZKHgPaImFlC/FFK57p+hVXz06T2E9qTiWs9vFcRNddfLDy
dTD1qw3UfafdmfEP3cIocjn+ceA5eU+kvGuzpJXpOYlknSswbXJy8SGEIBP6jZ5f0z+u7Sk3Xf8U
oaeehadpemXWtp9mwYBF8vWmydaZ3PZJxqee4U09XeCSEwkQBEj97kX/Il3qWMMGhcbVmtSO7K2Q
Ca2S6xXJogm4Wb5flgWc0NPSI4i+h6slQx4UWXeijHT/r83BcwEaMDi2RkTWHnNO5Ept0y98TE66
2Kw8+FcIZwU8pJy+VaYCTeWGVCTJ3PVYojIcunOZxuTww4mICIPJygvYJE0PURt4yBaO1vOkmnfb
GAqu8FfC9s+3ElWkNsCwKnYo1qQLLcy4La1peqEXaQvUqLrWN9bPtBkKJ3h0Q9YsD5+Wr919c1iN
XzJPjowYas8y8Wdw4yBcKnJm8eZRBfWmF63wg/b3AZtCbDp/1NUc3Mg6j4jJzEx5qu6KPddfcRx8
w+d3ffyk/A7dge7vf9/biUWqXrqN3Jvwa9yR8uhbUvOyd4qhHehK1hev0GM/NUF/28UZvyx7grPA
6jxp1R9/i8s7Vb6TBVZVEFTTbDgc4f7Ny2q7WS0t54rowvHLRO3FP/CH+FD5BGj0R7bO0VRaGtWU
6WV/cnmYMQzn/ylfJsIA88qUVGVBKyxBDtcuHgCk+lEgAK4kKSv4vlr+ATYP5GfyfDROL2bFbTQa
5bbxdGhKDPYdLGkWK7ahQY6UTC5adUVVUugFCYti5rqfz7iYfae5FA8A5+LdMSdFdVi8o5rgtn9Z
LppHJqCqoQKtIm1DlbOOXpdTB/ekqcP7m3N0bZih5QkSREzzj6pyHcS16uriQf8U+uEXLuI9NPFz
s25YzGkg6n3dUbmZ9LNnc5Hs8LXu3hoyfPvgudQCD20yqrRzqQe1bX2Oz3quIWxAeqaYC9C2YWEY
9tVhHK2thGR2hOdSsrG5lPi26s5b+sJ6GCe64PIIGv8W8A8sTx+HNJHUWao+DcRtUrtLF6xa3/+V
ove7EzpBJz51wB49n/CmlWd4VYgWUfSvXy4kyUqFWAOy8Ac0IFnM7qU+NwN3cWQ4eRdU85zstmp0
qLArhpIAbDXkP96+aqa4rwjMuU8HWLbYyJx25GzgWHbWKh9DAw/mU165mOraIa2l3W8eQmHpBZgU
v6fVsGz42PraEPNc6dkkBt9AaCiRJmNYmfwSgs3KqEXIu8BYPBw4mW2ulPwzupyYh7Kk6atY1f5/
nflceoJb/VIUJMaSGR1EbkfdchWOMn18C2+ntyc8ve95SA73mbN7ZBaDv6MUnLMkwUvF2gyUEXLT
IuFKI4lj38F1ysPPimdzGF2VN2MX0xi723tZLD0cPs9Q+Ljqe7H0PYK2iZdm9NgWGIiNeP9Vkrit
dVDo8dBmsdjgfo35oJ7RJ4uRDoOlGsSyHmVfPlg688xYx2mW1QaKvuddwh6Ps8bW7sVxXfLpu7oT
7nhxQYRDpV5KV0DC+KxG89hUeQz+LIs6Rme2GP0qnWstL1uI9U8GXMmAUz5UGBQo7vxW5v0pLCtp
lR1t5teFeAn+b7ADtYiw+GM9krEeh52fSPcmuzeFcqe2E1gtHkvSbOpdOM/ZzSut+YnDkwboPr/4
ZQlgnQahG/TJC455fJ0R0TjQ4bUerzH6c2pkErrJlARswwyQEugmn2xVjTZP/D1RRN6fYaXL2WFq
NUEpkfoXJA20dCGldunGSv3RsHn2DgeeEKImMKJJZH6GdvheyixaSV3Nhp8ns4mZhkvtk5/EN4U4
Adv7KrSKbpk+wwc+kC5Q7U/hUf99C54aOZ8G1H2lfHqQfzfltO6+OvD+J06floPlqe2xFusCxTn2
kZ2CW/YmERAousyZdQN3ZQFzcCSD3xZMJJFsO6POafOBXaTordAjifA/cKfIypiD5z00bPZZSQUE
6wyl4einU7+I7NAWqwvc64QDmZHLYxqjnP4czb6pTpdYkInmW1mFA8b6VD3jH5th51oK2Yt5QGwS
pq88BjkW6fx1XtfmW4ZWVQLCq3KvfQIqC9fMn7cYSfWqKTNv0fbgT+O0Qa8kzg7tbupIL9ePrMhU
jlKZvyIVgbBTcWxx7pAt2G0fzudSD+Nve09ZwP77SfdKHsRtbMwZbGyWRf666R8anHCHY4xx5MHf
zgJOEQ03mi/YqeBfIfRWhXGqFTzLlSph4MDiYAzlYIO1qojJlpZWKvcWXQAyKbZwTT9YIjiqk4CT
UgEVXng8lyjVNj2uerHaLB4O76SDin1ZBu7JocQvj4aN6Wk9Dtw/HXwxrKLpz2KtdWtMP6fsBFwx
cNPMLtHWjkbMSaDynRDGgbARpGq5GcGwL7ooaRGdAhK6L7ZSyONVn6umolmfI4ILAfV85GkteJ5/
E96/01CBMg0nqmvjfUbi35gnbJNlF1w4KRxZCSSBeZGgdWKneX7OohPUvPuGwTILMSjvimgaH4xB
c+duSN1MOqHh43qsY89tGMD8BGuswaCiVz61Vkd9CZd1Pl12Y6FCY3KDnAX1jTV0s4fJllIf/01f
CfvdmmkC2N9yNrJ/i2euTmI/UXcd1Eh3UVmG/370nKGMGfUOWfcxXY778sHH55CLzQ+GD6uBdiE8
2J5PSWVte2WDn5MydoQXHtKmq5SKbddAgrf0DhXKrzrvL0298fw/L1sWOSN62TaiE+ABZ1yOBUZ9
eqkfIE9Ao+NpD47RQKDBiPl0UBUF9lFOrrOd3LbOnhSYtfIuukY8hUXxi9+0bO01vWYJ9gDtXknf
TNyV8BV5uB6KhR6CoAhW9VmfF6znz1IC4qklwmrf9kyOu/fuSnMFiJ3T5JL7Ct2Ji3gYy1kiXGyM
xC7Ivqc+EXeve9c9Q5tdOinPKLlxgPdosS5oPhPIxIWNCYuaYcVpe/cBqFJLHMvVzIOgFAuW91tY
BS91ckJuD8eV6nNMtrCkq/V+Fw7ViwuVhkflsadpVflBCa5rHRt2Llh+dUOqYJ9bWdfr85RISGJ0
YCLOhCPxbK6YD4t4j2RWIvT95xLxP0WkEgMAEwc7kL3nbwg8H62de9efedGr0n1e3FN/c/mmwY1F
Z7UkOGOcnwYLsg4AWgppeYbun+lAJnbSO0XiUzGYPQERc75c/3G1/G1avyX4+Z5GCtr5dqar4kRC
dZLof7u6Rr4u+Ms1+vQKqpBwQHfJTmdnqpGvIs9eYn5O5QotIhq6Gr2kjsK4jSd8OFkff/Q9rftU
INcViyMyH1fsRa34VJ3M6izige14KXA7nQmG1dvQ0F9YKie8BieTJk04PlBrsQ0my1wpzPtcgSGC
C8yl50IhzkM3o19q0z3kpAoKcBVvywxODM94YCIDUiMEqFEg0Pn9hB47rtN8dpFxqDiQtyGM1+et
t7yTqNK0/UHpbNw4DvZi5GoDYU1bESTspW0+LWNgNJeWWBeeWZXPpIVSUPK7H8++n+43c4WlH004
ZK9wy37kgIcc8SD/qOf/bsAkzjCssa/WJ3G3jTcuG3xZtLZ/99yrSHbJzjb6DPQGABW7Ags+x49B
sG2KPPapl5lKgWC1d8qa6KcHSmvniczG3VwcGsH/moEsVWJLNnzPXx5HCDLnOa+yJxCfCFfHLYrh
PIEleKL/te/bmzxJm0hDPwH8RdLp0687ezajtchccrG4nBKeDZUEE2AXrc4qTg0F9cirhxiXR+MQ
OwsHJUwRnur6eUZYZeLChS/Tvjx/epZzb+F2TySl0dGcaY5+wko+iB+MbwElIadHBJ9yZBoqQPOu
IBbKQRIZdM51RwoFoRPFk8vSe237HTtNhJnN7SA1xfpBgRXe6PXkCuxUVGXjOuzFtZSMV2LfjtS0
Iobmc0r5TNQaaZGfU17Vt/HMuUTWRecVGivoafzKVLi9F4e1tglMQqirwGUrB8czhKNkU4GU992x
SCArxh40TzdJEm3grM+INaG6YfFoo1hp0Qvyj9zSdeVL9BoopAb39xQZD4/EBowhLuTOs3rGvWOb
s/CLqteDJd8PWlnSDQyToaa3G5r9TdMRntc5S4FL8V7nFGi9yQKoOxmC8CDe3EwZiHoq8EPXtwVQ
p51DMwiKGmFw+2TQJsBSMkgMa2cCGeZXLImwadGM64D3tM6PZ2zWOZ+3MdePygjlwG7UkpkqHXXD
w61pwHB9ZQcShnLkJ8NuV2gQHDwNrov0YGARJ+C8JUB4xJxH6AynQd+VZ3zvF2iJ37eYZbKGfY5h
vsDIGhwbGB/DxrSgihLXg6A4bQDT4ZzgX4wcv/rwNOblrl6beeeB+msg42TZMtkSjqmXezwCUfs5
NQ7ZG6MjhU4SfzWBXdDrBLOP3Z+XJUezSLNb3fqE6tNRGsFP6rXMGhWWmAG1Lvpb7JaRySu99Twf
4Hnfw0ar24gY9rSi5oeZ3i4GlzE8WUSToJoaSakCidou0joq2WWSeqsyFdTqqYl1W2agsCo9buxp
3jPJPKYrU/jVQxZmOUySHiCh91uR6VNtq/hWMPH92G9OGDk43us5CPSPSfeXuu0D/2ry1Sxji2yM
bHxRo3TeWwHdJ4hEE80vG8n3WhBlRba83RVjoPbmjPCkj75Fys/CYPsD1+F66mkllOqP/HSIq+Qa
1DGyg9W0B/rKtTFufKMA6rW1wwtRKuUFMhSBtxW7iYodyAF/Ccb3xjY3vwMMd/Q4A3fT9wzz/r0e
mNlkzmuIvWS/x7NK9PAG6Bz3MnHs4Fftk8hqknlW2BzXJLaIQ2I4khteOCNvLgzqKmQg23Q9LmX4
gvFEBg24+QJdB37rZyIXhDwUE/z9E1+BpSz/W6x4PA3nmcIG6mb/XZtks3ceSG/Lhf88472n7d+G
G0/4CTq/Ch31XAqTtYdo71fev132vZeXEZW7Rp3dtQiRsIi2YqoejDc8S0/b3rkeo2QMwFPVRqDG
ah1Ddfe1jKaupPUkogHcfAusN7lTECq2ruhk/8Af6jNYCKhYvJqWwbjJaFjA9vQ6na+QnpU7HTEj
9gp5UsES8ImrqR+xJjqLJeQ/CZ3OkIJIsUuRvgyHukBSbem6xWKc9rAkS0LZSyvxQe97sf4I3TfS
tc+ly+EaoKztwVB1NM8Fa2q7XHiTLpbUzbwRujNSPF8gwZVYZD4yRF99Bl02D1FykehEBiLJ2yTC
TZVkw1Vikq3C5E8ghsp3fCD6+SSeXZdagafqR+6nWXf3giaH4x2SZLh8FxOxC+QVYVfePwVopDmD
g/zCrXGtDaZAsp8XfVAVPA9M12to7ITaAQ8PzO23XmSuufCSua16dLMOWu1+bunCmyy8MJbjZEo3
EhcJrG60/qhVRcC+Q5xXhbGDqZo7JBe47BdUFj5oSrDPKclzvdGF2uMAsS1SddB9SeYMU0V0CLr8
gcCrieCL3BOFLo3k0Yg8zFnyAkPyKgt7o1KIxuWtNE33XrPJZgea+8LFsn4v18D2JIazJ7sNfEyV
b+8C88Fcz6vwU/8c940n5Dc5iquqFoHxWFUgSxznw9WKIivMHwi1W8uDQIMzK3p6mRJ/uZQvZS24
HWnEJSwH2AndaH207oJ6BKJq9n0AkB53hYI1c36MbIB4Gp1M1BeM38uNmzjf/bmlaqcuzMfdnWNh
8ElfODnfB5YlrGJ7sMvKDH9Kgvax0CXG5mQnR9B+G2CHui4GuYe4RBu6XB9ipt6LbaepoYOlNNiz
Sa7jNjEW1HJ/9RzRPQcDEbF6OlldONBbjumDX+Z0kHM97ZK10+bEP1K3/5LeY2XJAXAghugTHhcU
qkfVq5CAV85xNpRuC93xM6cCORh5BrlkwYxs/7mDVw38eJftfCD2AWmi+vuUeEfpaQAjzrkdf3/I
4CYJlRnEl2DFWCpcwc5M1RhvXKEhUCF9G8N+5L/i5a4hXz3+RiKHYo5mQa9J4cYPvTmXNeY8e9Gw
szPVzAQztHYTQoLplWGYxy5YcOd3+njc2yF4J+ukCGgyI09xkc2yBqLfoYRk6JDFItd2NHi+aIBD
rlsb5zQZm6Dir9H0355kk+eO9xerRYpWtzKvBmfeNGf3qVQgH2l9iKxZMjYyY5dHhIiiojf2TGPk
82mc9VGgTR9BXhyFSctFSysONQZ6gD8hjWE+Eis716gLVKQ3bw+klxKDeDlzTPOEvJxkAUxMQ6/0
RaFw8RHzrua4S5dbAKh4BwQGxJ6Rn605K9lqOBzVNjI0/uKWomHT43yjNBDm8ZSQWPJIgfJcYvLE
KxErLudmp3xZMB4MMLlmBsCdvIahnCjedjhK89fCALzVLTCu4trUYtR0qA6iB0OsKUD8Aigj6xCZ
p05KhJl6HeNZeTCatw3ws6I21o/U7WlKF9xnYKS/Cr7nppf4lYorRoqXjSIpFYEMVz4M60wdnKJv
tmnSFCVsEixRQqbmcLSiHRgD7UT+ISPEVgrUANdfyOMIEFVLGyEpaYFL83YJwQV8YQosn5UBhgbn
qo4PpaxhDGFBWTwF8qdHm6V9jBI6Xc7hmNAB+Mzkjl4chgja17FguXeRwBjyxtci+Si933fu8IPO
YDmfvKsPob2sEZ7WUr0mwmP2Ttf1+JiUj4HpCLaFUNS4xzxCGph09tXs234Nz+8MTpn9zsYNENtJ
7LyxiDCtBXfTEkPd6d4sBZy480iAHRdmEnBZt679uecess6hs9Mnf2EHK/E/VOcbvEumr3LJh6qx
ZPHPw75EPJJLFOOImI7UzI+QLnrK9HUhveMwwfzX70xheNmsPp+1TQXKanHqPydBVU0pjMXBIG0l
hv0zrhYZ841ta34A7/CFHJnPLHl7298F2Oe2Wzzn2pSTtoM2u2N8xuGg/cdjzAOX+qDgIcorS/py
cvborzRuDIFkyR05xZLuMT3bDTRVDaIpzkAmym8kiJkQ1hz24ldqaR7mRqurl60IQOF2dZyeriXe
NKyDoYJgC2zeZpYwtyMhWU09IoCl2llByq2CeGxehCvhua73TzeP9xqX32jjxbIm6Br1Rwjt9NJc
oJe7qPgFgV96PXwl5bbriOGjNPqqdlfOLnqOB6wIudDfa2a3QEaPRLdVsY59FJSzesYfvnyecd5A
lvH8efvFJtm1WxkxCR86/Sxeo9miF6PmwYurKAR2UbXNsuRnozd3DS9W7V6Vsog97RFIxhb0L8TO
/M7qLRjlRP6APy6O7RqE3ChMz5JdJX0ZRFQ3KyTFsFG33f2gbNvx1C5lsswTLM6LkhBDBRVW5sXQ
wvWheGPMDRvy4ifUo8G0mlm98vpJvF2DUhXYqTP2FjczKzH1dM5UF3TxeG16+cX4o+oFo/ttxHjK
qlcHEenDOtqhNf7hQkVwdIk7MbVhYqyNiSCwruqvrkfh/iGxlpgnnA8pPFDd/9JcwkLlKexUlskX
okpOEhirhwVmbOZFmEHzOomO9zwn7yGpZqA5QBPgDw60F+Sm4lxgrJWlOzrHtTgNb4/pDe6T3HpM
KDQialr0oOGn+GalqsEJP52goy8BGuonIsXJ0/eNVNNugPfwgf+H0BuAaB9UHAGcRksHLVfOA3A9
Dsys71tpZuXfKOp+bWtq3QRfdKok0ouhde+sj/yuMIaIaX+bgQ8SJAga8aZE06/phFu0kH7rpB4k
to8aVpF8LiuZSbgVeYwnWQcGsqm47OVnMgSXutC4Kry9DmadrEQQnAzejdTE6VQFEH2AbhMdgUlX
2iGiu1RPdjRMAd3yrj3DegOzA19/oI1ptPsKcPuwOpSA1baqD0M3rROE+55hzs2sipVmMXub2kT8
vshrFalfkwEI1pQfo9iHRkjDjBpGG4t7W1xfnzAX49VfiTTkZ4E0oqKLUPPweebruwVqjf6uonQQ
fyxfE35GHqTHoYM+xyL3pz76t93tFRR+hny1rzV7VcO6YGXB5IyrWCYGiIl72rLeKLBbX3mNS5KA
PXJb2z8zo7oNtz9G1bgyGt4ob/M2rW/yJcy2KaITuIEFKpPc4gUHXi1uJnp764qOUeT62tuR47RL
be3anhbo554nyGPp28kJFbZ18IopwiYM4LW5DBnv+UyrccrJG1+2lkvuv8do2ew+d4KR0n62MJLy
7L2Rr9NlcjFk8+qZwvK0v4mYeSXuVx8GUYZIbP3GaCg8mXGclGN23YKgAWQRj1oT2gPs27gcTK8k
uN+BDrl/5/LsaPszZ8vui1EOIVOrfnxzzNI5kt/zVT1R5hrE8xXu3YKEtUj01b4omyk2Z+dhRvKJ
QaHTnRFn19hKHGn71xQcpWGr+okYpqnaJ42m+2lv/jQD8YN5FciG1iq5fb+yXzUuYKVz/rAR/1Fp
VU/rL8gwAaDVNT5JGrdtCEW6ei3Zb2d5ySam7sw3TBghg9Cprjza6/JCaFOjeR0OJkuaYH6k6WQV
AxveoF3FnBG2Ngu/IsPAKeR9LD7cHu1WUyaOWSvLqUJQaq6AkjRDJYJjSKNSWkBUwIGLyNRXOy/+
1s0rHkRfxwaWjFtpvaBXFsGGisCL1rIriyp70nyqWoC7T80HXr5KU8D+3/ivobKDSH+qRfLkNlrZ
ZtDLePNiTKeYpGRGmqiwtTGzvHVYcXOLGxLgjp0nnfWBjOMdoES7x2aa41ashnbJeSevg18nJ9XO
kMbkA8rPP2Ol0lfAqHFSjvPKa/+S5NO6ZPzaTVh8kA7EOLZzTR2qu1WlpeChJSkE/HtgzcsM3Rzh
X8GDFVuxxyXhXVx4hGmE4G5mDuT6yoG98goAXE8ODzwr3tyG/f0++95fNW7pZCSutXbtyykaOuBT
7UflZWKnnW5bcBQirhArUyU855643ZMpqV3Fu9ibikmmS7Q3sp1BDioecAuhzcoJYMtLnj/yM8yA
5nf3yVIlyZlkE+O39voKOagB8osciy6vGA4MX0luKu4jQQrg7ztlpz67drfGXAgUTEDStrcMCRjb
X8mJ+fannFShbJlqL1ckmAZKOIHG/K5DRsQ9PXCaNm5KEodOoMbFjA8XrRAoZ/kQIfeZtq+LQgQM
TDdWFEkV+kQqZqeCMb7V4pLZuK7hIkgGprrs6rq5JcGFfbErpVuC1jFpHGaMZDRR+Eaf7Ckp9cVg
7SVDebvi1vTvhQKJuopvWcBWHFEYklh0OBfabjw0T/k3/W6+x/JmKRnuOZcS2yeRlX34tfp9moJz
sclLQ5X0PCmfTQTiN7TulDQVFQjutkcQEZR7GJ41HwBcVPI7a2S7SEGsH+rnTHt2i10Tb4qfrQZA
L/mT4nfajb/Hnmmxu/WL4MVRNA0y1dPpu7/nrr382tl3vdC7mQtHYI9fUIcXhHytxtfvchFydfWJ
mEUDxNiQuM5uxM3DymaULOzDgt/3cXTZkEYEPS9QPK2ykDMIi4B9cWfab/O1tJq8THte0TEyMC/a
AAhBJO2QJawCvP+c/DYsGvdlsBnzaCFH3GZ0pr93M7qrS6GqsnWmxOWW6J4zrwbYVIbVfNg84251
SlVxWUdcox/3YDENL2AN07+bnxVLpwDL6J6F2RopzHb3Av15Acw4r17yKkVmoHuJpVRtKn9UboQ0
auOXN2BOf9DBZcWZgmvzcOajHpLUiny7fYXAbTgjJze2dK8FIXU1me5H242EXyygPdh435+ic5Mi
1z5/C3zs5Xrav+LXLoQ2qXNs7HoZWH9/aYu9+V4FtY9oDw39kef8dPz6EiOPsnJs7UJ2jdKZMs0E
aJny1xI0lZsq6Ox8Tvp784rtznuYTOuZdlCT0b/+Sbgi8+hCWf/XEZzM04rIcjyz0ML6FcL4ZW/V
QlsC/zjfdiWBfB9V4bAZdL/C3paSGqvvIZ6u1+swvlT7usdWq2MQ/mTW4cV55pCLL1FTLzaoEWbi
CVFaoErIaXDzYERZF9V2gKWaY1axtoyGFQtgsJ2+krT4z0O2hoIZY44kijHN+6WxMQdfGOhbN/4C
3AUbYSUKbOfK1mOwMtERhWqPkkw2OFYQ+fNg/rzkRLpa+v4kji05Eqznx39qTY/KP5bfp/paf6ld
e6uu/m5ZWOIoFE+jt7n7sEuy36V/qzJ8cl8NMUgIN5ToIzebfMi9Z4HKCiaUjWDRC4tkRTrBCsZ8
4WO525OxqbVCu/HGOrW0VpJIJluZrDfAho9fAOS6pR2nvYB9c67RdYvIoMBT/DZw15s+dI4RCQQr
bFO/KHIETImnXtIEcpcIhp52xku7rbjCcUjTSHOm2up54uj2VCFnYbld+na4h7kspXJ0UpdOdlho
MAHJAKSOSW78M/agMAwPHZs9FG7+TRHNxLYY1eMehFZftm9RQUN3/6nPpceK9DOLrt8CsHGjCKyR
XeUPD/E9zOQ3hs5/ald/M5rCx8WE9siCtgnJy0xps04XEAO6moopaQGmJy4oDFOGY2M06JrZa7rn
4CirDURav39FgSjrUFMxA73x0XAhMPP8zHEKXCBnoRB0Ic9xZILTc6FUBrJpH2B1rqLeBoSfYYYN
pVWa3ZoBK98zm5yunbCWaONBAah2K6S3Xppzbe6EX7BS8FjQUjatlHZo+mTe5A3b5UIjUrXwNl+F
uo4uo95vySqbUtXvPj6yNl081Ou2kFzftduVOCUAot46eXKTrDerVi8oaAhHc6FYCNQhLvbK1D6x
bt7NrVrH5i1mawjjq8kGHgLJbWXJ7j62wn0KOvsCFcPjPV/stb07vGLFMEY0k0YvjUqyqrnpjhu1
AG+S09QV1n98rAT/M2gEtOUAV3DhXY+w58efxhqBmZFm0TdcG9HyD9NV3PbZtTKMTC160Y3u5vw5
rR5e9hPdf4Ir8BHPWUop2a4ufapCjhDpKIycQd74t5k96fDp4+mCjXmS3WDqGpq9Zl/0f8Xv1Aar
ejqlqaXD7erZ3k9BtuR1I0vd373ra4t8WR5ziaVikF5onY1O1aFeuIkIH0wopzyFQyShSssXgFLk
Z+iloBWd5ChNQM5Anz0J+A5ukCsuS7F8l/+XywUOoBuPmb/6kJWbMin1GvMgodH1tn8SMhFhGDIu
Jzu0kKSINlp4JlNDTfY/uKN/CDthvZPAWRZ00LkDPv1Usr2byc6dbwNeq6R3YIz70HHN0Q4nMcuR
GBQRxllgMaZpaG21d+DLyLLY7GcZgbrAwVlaoZn09hy55NKQeJ00CJ1htjv0zOlXe3UdnWsihg7A
B1gxLT5ehZ1HMGW7fgOpAn8oF0ZfHutvtd3Dp7s6OGtVwFTIWGKKkgEGNoizBp/zqxlJB9DireQL
hR+sNnYx9qntuj0KE/i9rmw9yqw8rknWKfe4Docz2l6uhNkzB4wuwAksCFPXsRFp0pTiO7IQFWle
Fa0d0+UGh7Oq/vTmlEkkatnxqnw9eHWUhg7TQYTpGj85GuPhYLP3nqczH+t9FWVTmOybIGBN3G6K
l5H7+lTexE4Z/xbn+pC3DmvEFpQa/+baAxz530szD9XyhBeGWyZ7Bcpg5Pw/UYRyryGXKwDMk0o7
mxCs2rhiZQ+6HRSXag2cXFGnmb7Rp8SN967CKQKjJHS0RiRi6HbVAwbQRxT4Bdngy2QkdWpvqiMy
aP1w0WywbeAoXZqTTimD8+YB3zcHm+bkRt1zys3ZpidnY+7y/zl81HNf9Q908FsJuXojtPeYPOCx
U3OAv/ssWQJYBgH25FC8/3XKy/ACNTCJ1bikcS/HvPK9b2yyfBipf1i1/K7vIXY7OzDpbFhj5b+i
V4ZAF+RtB+4i7X3ZT9je+8US84mrM8W0LxmEYDcORD2ffD0B5xQ+0z2IAr3mfjGCRbP6ACSdnDAQ
4xeCuSF8T/KDqFvh+DNidTWtNDIwv9O1btVqqR/0gJ0CoOOQUMpuRHO0XqI8W+9m5tZ2jM+HjsTL
I0itCp2So3SqHRGX4iT/KXyqTPLP9RMObtryw2ItOhjknuiYek7RjSUjulDIuLyMrm6NLuDObvF1
SzPuW4EzFtMSdozGgaDjm69sUkAhneLrjd+9qVrgQ+QhMZtQl1mga6YZ6D2nsxqAfsE0Qxq5jInI
djINDTxllsvmvZ1ibXeoUTwrNsNndiA3wHdhQCCC7bEDQQDJbvJGtbTBP4OVyCU+sKPrAHip240l
e4XS60BEtKcydH0yMhzdIKX81+H7frOTG5JqZTeRLZrbRkHjvJo47AamSdn8eG0sZUxyNgkYZ72n
cDuvzxJj7zwNoW+nQChInio4Qm3yDDmGl+QkoWnlGO5LyHQqfpjwfpVoG83MhMdumV1a2NCNvbI7
4tM26YkaLhDQqMGmSSuec9AhPI10f31+ayeeL9gWKgrP1fSZnw0YrSqWhoLDuUUfPSGf1ki31hVe
7eHS+GwcoIw+9COhRR0giEuMVCcZPc9CSaqO0YHUGV6ftiYC2uSFX1uwbey9x7oAbVNWUVssl6Ym
BH0DszKWdr0idnsxmBCUR1ab/t36sDOOv7JQas6QRZJjUYjG73FfeXKkJnuaFK4sV30e5cyRNvMv
BcOaeHSP7Qhf5g6DzdZnbxkBPvEKTcVT55JavTIjijv88pBA7WFsdU7c6BnZQZziuq+JNAm1QPlY
FWK+G7lMmBeWL7stdLjl5ramrRjCEqFAPmOmgMKnIMjBjHmyKALEE6KPHxTBijfbGaqBZq4FQSGo
BhMasglrQxkX/qGNHclPxiOj/GgIg3KeXo0aOEhGrMXJ3kKExAU0wJpFMNhx0zCmq7OIljGtSMcb
KrC6+coLZ3BRXMpYf806URVNAHMAjljKos++w6DmdNzTLWVXqBZHL+oCD6cjSV0kZL3DE/v/a57+
EwCHrmztgxOjWrI1X8W/FWixU/AdLJ5U29bUkdMs1vz4HQLQxPY7IpTYEKSgrGoZq0HfHzasXdDk
YMsC6y5k8jgT/8q4647kZTA6QSA2JO9IiX6fbsnm22mYYAg7htOZF0yUys/9bUu8OtDBnPvtfKSS
uNi6lEAC/PAahRU/KiQjo4k1fJ37LbW9FHALJiM9PNGfL+9ESj3gwoo5HK9glm16BC0OxKeMnDCA
pUReCWrJpkNvYptBxrYP4VU3hcA2W7k3/YI/l62RrjpSQou/+K+dKNbLlN5Fpkm/eDon/4Gqtx0D
qaZ9XxsyZsoST3rJ2dTv+7K10wdLn8jFZp1pzGQRoIWbYFvtrsPgZymAi43kscR4Daf87/dRhMSO
d+Q4F/35h2gw0qjs4DzAoLHvh4S9GYe1Y2jeZFm62jGCbWObuCCvG9sJTc0CVEKt3xtwG9MobsrV
SfaBnUtbpq5Ii6UcGfSQhCyqjBVr5t1dtskXmoODFbSvemxJPzw5hi4WuH3b1uRG9N13oqZUlp7h
fs0ewJvk0dfCBPyt9w54R7WKeBg9lSpe3jXcXxyWlZv8LwpOE2u6e98ReRAKBAG7RJ0/5M7xAmB+
eGSLnnv5NUFXMWJKigaWcHbovmg4gfIpSrdwTfb//O4x0ZS22XADiq69MEvtGh66u/7J1ciuHKwB
e5uuAjriTRVabNHv965BKo6DoDwHggwt4H3ziz1mQkcxgBhrEgE6dyETKmBfXXUL+N2zxDunE8lB
BbieNoEddPvi/bTJHDxzNI3AUOv7BVH7eXkcmaH468W0k/GWEzzrB5IZlMeHpScTw13iMYgn0ZtB
gNMiY876ZRLvXZWVMSbrqP+EScDS56miSJy1nYnPyuF5BXcQjq0rkKKrG3eWBd9/y3ZRPu0DE3Nk
E29nNWhZ3kqbw/Llg4YMH0ITHX2eZR0+OvPhU01FSi2GAaI7m2AKVsXvmU2y/oI/BCa4R5U5sJ3t
Xnx3Hu/l7AlOodp14iwbWghLjNkCyytz81UO5DXx3ByKnUGuQUoOUeTdDWlSATDaDHGqxNlxYPIt
47coWUTM5ZzPOM3Zzr81wQz7gdrqYgRQjtPNrYtbeBkO01WJ0cuaM10iUrNbmHgI8i8uu55Xu2OD
SQ/Lah5+6J2wp9X/lIP4n+ge7Tli0buB+ZtWSpceFPbPqueNLNftHSwwOLCi1Nw1/MH1uAjcM90W
Bc4T+mZUt2KBKG0XgN09FKkn1OI7b7+hiVqXWvIqI6A3lfSuq38XEeegZK7LrUeyfHOpLEKiXKat
QElK+uq0dEPYlk71riQmEVI/56OVYCksdvx1VnpmtvGuv3jeEL5OHfKMsp2oe6+dUClipheU1pa6
t5CMv9QWBd0CBN/H8tL8ryZ1p6n5gLZH3xEqZ6dymIRGhNI0UP9H8sqHah7r7VRC2Ru99FI2Yao2
Bur1fObYVCdFzNzFIQ46MeIrkoUW0FXQACIwM2YqMWhmUvCaeHNuGdNBSl7cMZ/qoFXAsfwf6XLB
DL7LFo2idPsrbWGDAPZaOEOnqDkVh9Ad5C/dZGi+8oWNvlpgn7YyE74+p+GlwM037tlkfhGLfoAU
3kAxJLgGJ7ebVxRJyxnBZTtF/NYtIazDgR16pFAEvYCk0wz/KpBZbT1z6CO3qPSUU2ijFWw3E8Go
ht5ZV79TGz+wHNH3yyCogBtEJZYfYWnlShl/T582HLR7zN/jHoWz530Wca2XOagFb2p/Zo+/m15b
bP1banxEu3w9QyKrNMZypDguoQo1B11wWCJXcFtRyUxdU4bd8t3F8iH3OIgI+nxw1a5u0LoRoFyK
B6CHH5EVY39LCsb2w7VdWFcX/P1qPgIL41aZ9ydJrDQPRl5TGceeRWx4Ovv/nPxrg7S2AM8aUJfs
8QUYq7wPa9qHIXfamkfDhk0BjZOYQZ5gE/nikxp9wTObL2N7sDJNiNTHHAE29hGyO/yvH5qSQbEZ
S87BulDGaIhzDUf275FS+z+wW5YLxPIQQYM+RdgMWxiJGgYtQcUURZASPzc0M6FuYQjym7qk+vgc
dTYKeURFcKNlbpO1Hb1jLUuY+9/Ca4poeW2AKNkXZP5LW7/8FGLpIGhwrb+zd6YluQ3tSGlliy7V
NAAH92LTeZ4AAAaDlMwfhbWSJWgfdK0B3ZegRQ/tyxTA77wo5lDHpn91zqU1wtdYfYjVdUTQWOIU
KwRqaSkFTYfqbq7IVyb4dtACE2W9oqyD+ddBgp/ODr4u8Y9MvcnmuIbrXWyyel8ZpW4fB5kSPJpr
AA2bhAgk+++lXTeOteKJLufhWIbpk4rc2qx01PS98Aqrooq8IQp82IFPmF+XGnAUQhveJhVWwyt0
rMpoJgfE1uepLod6WhCwmbSmZ2Am7kQkdwPC6GE8qSGWqDchGCxwaQ6QGmX8u3bLae88GtWmHGwZ
vyctN11bb4Y54nDKmSiNb99elSfSnQuxKGceYxpxPuhIbGOuBcKNrsSqPdu9OxcwC9Aw9mQO+p8r
eA/RP3WHxGeD5faSNTaUJz5qneNFDSy+QYpwf+MuFbmwygOUM693Jvj2SWJADiPLUSxfi+ChJs6C
eE5HgwO6Xx+JPkkNRkkoflGNGM2rIw7ovsiuy+6UkW5/dr/f+A3uYTZZ+bGFm8QzXh5oolBgSPL7
+/uMwbkAGng7x3EdIHIR5d4dgg/GobMtwnFzZ7KkpHCpv/erDPKU1RsnapZxqH5jtovrP2Ws6LRD
9gDZu2B1EzGv8uT+Dtp6a43c0FjT+ztyug9ZtuW7wmEwMYTDi50YW/xeK3mN4N5Z+U4wr2nHyaPK
zhKckbwlmqrsW+yL+Rw1V1jJVtMOjjfUAvu30KvRQx/dM7uvqPJPWvALLtQo2hfISJUFIdmoahf0
7RKYmqkobGrLFoLxsq62TE+xx2pcdVO0RnY6Oh6vsJrc5660WJMZa/PfFy5Kc8hCnOpvkXh6n60f
lmBhfWYPjlSy97IFmGR7JRx4dqq2hyvvjwONAPbbJEAfJqLu4qSRE13Y16WmSnf1H8e0QN6hV0lR
a7xiktpLmkSy4Mz7q/X0ROdrt8U59jOa0xQ7ZPQhkqD1Y9Zkq8x9N8hSCQcCXvbI54+GgOWTYL62
EPs5LmXAs8VH7L4iohG0efaC2rugoLDr7UxS6kNWKYVTfqGNqyVLGqaRe98IIiVBqaa7DbGBPSqv
qMocOw5tCafh3k3rRR3dkq6Jy8fkowzGBbnco6nmMw6NlIoGTjlsz2JcVe9nfgs8tHtIn9SWxhoD
8GehjywTbfVvChufXQ9LBBUPvLtMyBdAUXPXU3dJS8MsaKxJRaOEpsousEUFldl+fIK3k/fCfI/D
8cDU2Sc0eqlzfT7/bfHFDisGGihsBLrymfzYm+Gro0XbGJpw1UTsYEGJX8xbvqQlTJj70csZ7kxb
+a5RntIVVuLbDyUCHhVWZzzKtet8r/g/bin4L4HUVg9EQITjxUpjbKbbfyaBiRKmZQ3r60oxJ3hk
Fdg+t+BsyxPmE4IVBJLhVylNfB6RFCnxsWAELWbGACEg1DQW87CKRH7w+gUksa8ToEOzmSgiaL1a
QtZC4NWuBg5ts9zcQncm91pjd8JtDcjgj9chq+0hGk37u04FuI3m61YlxzuoYDJmTo2CqWZSo/U8
68Uzo0zyQLfv6EaMTij/7DrYQGCvfQhJmvDJt6oVTHfg9PX9HTsCHv8ao4mtADZ15KH6xH/UP97x
Jkpst6u1eKhWq1mcaCxAX7YyV2fLEmUCUn8gnwjX3KyWFOqz6aKDr7w0fbg56y6p/JWnK7/taGz0
qz4zTdV0bIjEOqm6WMU9UK/cJB3sULC5cFCFDsYGpk/wxC7HJgq1WsaDXl0QoWPsMPZA5mUFFd3D
rvliFkGbmef6B//R4Ryw2RZDFquagkL9QTyhiZLoBIyIMcknSdzB5Y1UOUFDC9gVB84F/b7O2bmK
lfpZkcOT9Cu0tOBWKXQDN72Ef9GEXV8XU14bZq/OBCveUiAOahTKJvU12az2Zlb2LxRjZzkDtiNO
GzilGyjIl+a3IFO58Mr8PIMeh34ROvaLgRhSi1znRDK4+74qYvPqSc8f0Z1ucWWJwpGb/eopc1Pu
RybFFpkz/ja+RJLDE79O4/CHzRCAobLBeuAxg6qA0igk6u+inaA83l6KHBOG1zqUH+iNjtqmK9Hs
6Eo8qrl7WRAc0SUJr6lLY8wsNIvjJMhxmRgHii6vEFcm/CGeqKlLNYXQS/f29rpE8BnihfcIos5f
YgNY6iyt1j0BHJ2V38NSJkjciI9FrhX/Ih7j4ArIzcbqxUEUl8HcwVHLo7ryA6xEygODR75Yn/1g
o15yOxdbRP39mypZZJQSYJVxMXPDqrjMJqwq1DcSipvdg/JNBaQYQu0vxS7JurOmKWnEsZsePTpD
MBVA9hAvukNzZmZl7+B4BPI/ovImoe6Cw9OklPGM0HEhLtNlYc3PC7pzH4/A84N+oPPFV5AfJWb0
iYDo/KI+lQp1QXn3fWglJ3tG9LxsK3uOR7gudapjvvnMCgib/r3p3anGvnWudf24KePwuvfP83If
3UDdjittuPyF+BYv74M+2TctveHyCaNCp0UyBTc5rYqp25uFj8t0qNpSXcKWuhHfE0hqn/2DSs4Z
ZCEzjSJd2/K7uhTC0HSlDo+7ZNYFbrW7TBDRIZiv9pcIGxLrr/zeAdcGnQOpgE3BUSYDwXjLObt6
KxCJnpKfEL81TpwflZoAtxWk82i3ORHuETFcgzmRL2KSQphuT8XCobh6Bs177pfHgZomAeRoXsrZ
LSdWGEuknT5kWYqMHWedV8Kr40Ixr+33gC8XXkMe267p9DAa51M6cztPm4S3x0r8yJga6ShBy51S
f3/d84cZmc3ZvWJ37BH0iC0adOywaCAPsov5/j/+ILPUapFcDfuxZyrq6VpWLTgSe7Nz3AEP3CRK
YFgyR8xnYRoLbzrCrh1YXgu1rzpYRXS1DqGtci5GmRL6N8USyOLW9k5B0Ii25r2JKeQCZHdbISGn
O2Tp4JJDubAD6Kj3paEbbmFHmCzmZ7whrX47vfp2LD2lMZSleX/7EoKlcg1m4tdyrqHLyrRhcE6y
XnnJdFpBsib5uOxM3m9m//QvrT/hBsXVt0dZUJqi5UUUSAwCqRcGIN497JtgHIgQI0T/+/I8mzgo
J3za1MRHEfNkk4mykbT+5HqqQ0IxGRauZ+8VP1mnekM9se6lYHzLe3kXMpTpM1VaLp3h+jPHtbQ7
PjRaF/UIB+0T4lQT/n60zs+sG5WBcW7Ph6a/AlSfGiVZuedXJnc1JIQEyJrOs4u9GbIj7G9Jhtsg
UBnVq9DcbZKiqxpNQS970gAyl7Ukw5jzGNyF1g8cfOwYuZpVq5Hr8dalKztDFp7gKvNIRDu5NDGq
O3MWihBDgqALZxhMr9m2CJYvrKc8J/OqrXtiDX2TqqYFEebtP6Z9IHsqyAg8XwKmcavwo2++dfoM
/VclezLo0gUNifPVw+LAxqNTDz6KnWhKds+haU3p16gCvxhW8IpCeTYgxqTR6S7ybnp3sSUhcqX6
+is8loH3iNdKBoY5XiZNGibrGrHA2sTua+I2RkR8VJAV98nk9gtJUFTtPYvQeZ5t8A/a+qR3tbQ+
jqZP6iRlLLpwu2vS2trUo9GuAxUnlSEB9XY7aq9+DetvRyWoR8yYixFUMQfOCDHPPkvn4AIBEg5G
PRhWSacdae4/1K1HAHcF6XEtTSKfoD8PiNJrSu0ZrzlRBSQFWatInxxsxJYbOgaOr8QzzjZhbOlG
UimPQNqVbFPX/5IS3dG5CoN0wPiZC58KWTEFS8/gQSIBhJ8Yt5EEyR4BoILBxlNi4Agg885pl6Qw
Gp+ohQpUsKnBwMf6RC/dZLYNpRaytC53QkNoLxsHXRVn10kPBRyOP6IJgafHB4t6Chjmqstws4eq
WPUSYnBgbIpar9MoQ046Zvqa6hlMizfHSBTYh3XgYuRptjlvfa0eUHACNvhQT96WtHk9RyFKLm7n
0PfbjatUQ2UPscUrX9lfXDUVB1/beuu1ZtYncAHualqOnrs0MN7XqAYEtW/g7ZBhwcRorTgkSuBP
ouPb67ObvRFqOlq/f/mbLLrkX3KTPV/qcO4APo2/AiKW7ylcMeUmSOx2LFbrNQL0+wfULx+Rkf/p
o7B/SrXUbmKP7Qp41skUsO6PM20CWDCM02u/3mMT6kh2gxF6KOMtsVuES72tH34rj7jSFD2jDWxx
E87VMYtrbrYZxhcN4h0UUsgS12HTNWAcS/+AZ8KsYrIil75WHLtGnuglhzXgbo7gyXYgxQvUg/E8
d16vTv7KcH4yzNc7TgJrSYNTZ2/bCwNAoM171P7eHYFy29VdTcTDDYgvy79qVueE7rl2Bqcv1aKR
mgEVlmnqLSSA8KYMK6DIH9uwWGAjBWsVD1B4HzEYz7CXdR5q6uyOe2/px9KlPCDz2wgF++9C0IH9
cHDtNWxdzRzYkQtt/ZLNBLQ2kRrbhoo3aXz9IwE0oSVycp/lTLhhMBQpviSdMsYjwetXWTXXe5ud
1V+91rTvC8NTQkxNZO1uqIXNrsNpsQvHE1GjAUHiL6PENoc6H/Y8q2Bao5JEkFL3hLbwQe8SPCZv
Ns3AElIXvEDw3EBiJ98+epjZC3JR5PagixXmPsxo8D02xza6H0eMtMqV1RcEIP5sh5wJPNqTfKaV
4LjSAg7KHqyxC5PuppQBQCeyyDqpIn/Dq75MgUHEKK49uKNhVhybrmGNU9upVeaqxmKaIrXZ/ly/
xjkyoSuyzJJlkQrUrOyuAgGdXaWGAiC/3YfJYFE2z8mF1wGHNl0Tkz7K8nO40G5Q2pEbFiiTzKI6
5Zbe5T+jBphKwttTZkNJwz2aKL2MQxlalef8HaYz8TncBxGx2D7uuKZVgZp7a53yu50Gp4DXs1dL
/K7zyFB4ymbJfKV/rjlHssPQ2QF/f2Rc8N4qUY2NAZDEWv3tMgGiFfQsS7zaAH4gtfTrdlX2/rct
jTLIAqt1he3u2naA+Z588qr27vB72zWOvVy3bNXQiAcwSVXS3ICMuYg0zMgZmMiOcPlo3fgLHwLc
EMJipRAZYICR0wk8sr5crDOZEAfY+IDbpw/uUdDNDc5/jpfBBaqu74X2g0GL5/sMivcKZ/M88bP7
YVtlnFPQEfs+nzpIIBZYf0/YvYdR8JC1Q4F/VqDI+xDHv8B5Lma823AG/W7G9o0adfQpoP2i3RUU
rlDp5Wb5V1aCdW6vh6at5bw3p4bKGrsGHSTxATcsiGN7vMuek/jDUEDtZnZM+dSWKI+2YOM5BltW
vMvdr3ocaoMQ8M2OtuLS51fGAg2/NrS/9TaVlwijr74SiDVQVjykfv1YTTLz3bLKqT7+1YxDRszo
fkK2LTvvPpOaRl6QqrSfARcvHzEoiGvyRK7ptvp0aoOvNZVQPynhtO56W2Xhusz9UhS09Q42hcmh
KPlqgX8TTXwaD2yaSDdHDTtOibY1e9rDG80UppzVmfNIeY88ySjFWQYRBwyjAcfp6wgab4XdTaXb
9Cg4XyEBeqQJK6ZzV35xJbHNFirg51eYum16lszI4HYEWDFvD2LSu3AdCKi2USXxhkGpABiBA60g
mgrziWizKLlkFTJqEnUaDsY1MzhLKI5M3e62am+VoMaPZlfeMK5zc+ixVPeYslgr3uzW6ijZu6Rj
ELsNfdxhsvNvgqCM7YcOjSWETg6XSRKkaZgQJyXEH1KrXIJdUWSjarJ/4hJG2KBV6SLtZP0egbQg
kWPS0aAOURv9p5+ZvCx9Y5JjW6BzxcdZTX7qQAUGDWuznDyZIUJsNo3YbF8mHD/+FAvejTJ8sA3e
BbzKagjzsu8mzRgij6PVaw7UFE/yet4XCVfOkz2JZS2AnbiWAbia64qM3Dfh0S+bneLcvvchAbbd
luRzf+cjKyPv4WemF4QLn+jEaMStptz+a4iSRbjhYdmDIsCcilBRCOMPfb3aOyyb4cWDvkyjVQD+
zrC12jsiZ4XC1/5BPOp2AmM+p17cnsfQFheAkuSkvepIT4SNKSL00mOY4lXg090NRP5Ic05GAGq7
lSXbFAnU6SkkO9pd1Uq+/vmniIOgHrvi3L2XhljYPCa/tgotPpeesXC/9Cb+x5ABxsZ1O3JWuFJg
VhHocvXk5lN+0Qilnv89y05IG+P3RcdyT11XYsCyz3HXNs/rQieN+O5jHPn3dwZjjVDAmvG2e0UC
eXIiLiCFEA9xsn/iKkexglsB+OlSD3X3KPqI3B1RVS8rDvtaD3WLJwKqB9K6fKuadMZYaknNLPSE
l0If3EXm+C/a4L5FBQFsBzZ51A2T3BsPMG1piBzMS9y/n1I8zdj1aK/CtiXAX0YE9NtnxxCsUDrc
vkyjc1pjPVpskasNmcEfUks6CsHOvBt8w8pdEFKtzTvMePF6f0hjtPZsUJkz7cLVZuhk/tstV0Hi
RaCITLXRtdCIvQIWlllXqQQYlsqwPh5cmHoACcdP6DL4v5tD4MAasJqjWtka9HXT0syxu+KoIzeM
XTG4dAx863QlmbsxvqGFXxeMLBRNhDQlYkAHQUIEPLOJzoy2HZFdQWQEAo7LhyzHlafnQdWmNlow
pWvtPNVDLDwgmEYSZ9lJFhjbwy75ZFU/0oy1mk41N8T9uR6M0dvdO5kza5Q8F50nolPOgjx02VMJ
xDoufQLKlKbnEw/fDEbBo3YzgstyjiDSS1/IasyWaCr3516BFwhw4zzfgTVq6V09xeoDjaGZWb3u
FRcoZN1ohddAyktai1c1y5fOsV1EgvoTrEHOilA53jkXdSPSL62oZkP2k2chz32/EopdMliwCgdh
JE/X4zOl0bXE26E4NQFvI5w8wcrX/H7UErV0NuGj5uZOGNprfRk14OU9KDf8lIl9jX0zH3J6icIK
CaglwAmjvO091FtqsJ85pkjWbQdARg8puVZkT9D4pkh4YfnMenxhdjftTu/mfSzZ2WTsQ92h43gO
mhKnB8dSxQZyauDholzjM3fM9d9TB1W32foITLYrruFzscQ19tEGAwmlSmIqa65kLLZThQAni0O/
2cM0To4ptIbeQKNk+ym9RH89dyImSJAFoR31aojSUcymtljeYhpZa1vLkSDLHtge5HOEjD3aF9jP
HPqoStXfDrOswdakn9IRE0p4wKgMhI8xrYhr12EtTJsjpz41F+5S1InZreeU5BG9Xq+Z8mBeLdR7
Otd2Hp4tuPfrnBOqdWgmSWu2WnlDxZPMlZCvAsQBRFbCTrVsMqtjITUSGpILU1u9n//up3wTTGoP
tdhavyI1AObcec8hgVPyQfOfkPGovXv2yf/+d5Cj5tIJTlydbNjMRiVsNkUbE/gu7W2duef/oKUI
yRgZ397M3J6r7tox2PVNOxdbfA4fRH2VmuGkvIAlHjtxYa9vYaJDzRnwWEOxsAk7mI7HefFOLv0D
zAqxv6DE7wPO408qq2bMyyxs0SQB+F5TfjjljxPTPM8q603NYvVXG38A8MXdW9TDkdMGSP9sgiQL
4NR5BfzFnpe/h/gJa4WD4BOr30YB1SAAwm1EYfpFqT5BONVGyQcikTBKh7QqTELOupKQo4TLyzmp
TFWRlixHo7G2MespMSbq6dNYaK3bNVMEToeqWRP49RdmmfEMIHxIcVMKKTmt21xdStbudtMyo8/H
lc1+I11SFCc3tlrRzxP97sTbUzaYPHTVyXvewDgPbyNUrk2dVxuiv4PK683lXWpLWp4OIH4fIQ+H
2OZEnD1hVMPoy2gZ7vO1zrfd0OhJSTxjTkicCl4FoLVGdjN8x50gvc0Z0MtI98MHlnDKSzyj0tOK
nxsZH+v2TapVyEeVgsXz/Srp2F1ukWc39IOTlpUsKsu7dg2qtss6uUcRW8Krtm9ZSTxsmEpnXjfs
b54ZbjZIjk/Z4hRYG2Jpmy7Km6FD40EBbyYp4pVviPDejHzCTuhIqIgsWjZlFKBYUtzo1Tj4aQoI
bjpbNrAqfjwpfhWiJT8B85cWXDJicJYfzShNqnzY2/dZrdJzegySwOLclTjn6sfy42X0j2dZ1oa9
OKGSXbc8clOE4tb3a0lygUvAopaJqOAzq4vBHyMjkIDRS2Gq1hkHi7BKaL5I8gZYah2jAFjRGsAs
jes/KNlXpFMRVi7eo8V7Hg3ELMyJ8g7M40Hyok6A9ATXibsPa+tU/VFRtxnyzFwnJU+xFsLbjVQg
NvAXJy4CaeekW/OoaMErKMbCZYJ3e4swZYgTQtu6ZiqVvU5xxn4LQCQq16YWFIVSKAz4lu9e5uGW
vpdSDr7NHcmKCQom/iwJ+zSed4p3n4zgkosNwLwQ+Acjj6dxixXQtqmSLon3UubKynC+/it5W0iz
FZpKKu8wH35XEnSKnwL2X0h9TKh9vOtm/ohjE1pMMXH5h5YegC9Cl9W14Yg2Zf6T9GHJT8rQKUPe
bjUUDxtr3djA6cJFD5HSHiWzmsggi51C1i8x/yR/elJE+deQTStVtt1yL9HMEv+WzRNn99ARIH2o
HJXoo+oC/EykxSh3iM7KM0A9UUgXnnsIPcmckUoySIC9o98CTgqhJTxa6qo64c0CeNrW034BwyEE
xmTd6ThtSkRGcXNtM2DqxQAuNc7heooZF5MXT5V8VuyOUGVPnwh7ntSBl9iLTstyGlRX35b1WrHG
SSYX3apdvl9Ir1xslmfqRRnqIY2cbCgLx7/k6Zab7eziFTR3IjUBqNdlA6iK3mLFeFS6nwlIe9lO
6p/MJD4rcjzaByn2UFW+ndOy8g2Av4fDCQ/M31n3NIIrrQCh6Le3PII+Stb+VWLfoBPVmLgQNj2f
yfXuY1RClifW5lw4QGqpacHPwZl5mOhguKOOsZBTQg8m0wRbJtmKUQ8OLhs/uZuUAV1PAuCRVRpR
kcywyaAdds3lGZIU5uKe0YE/eKqMsKo+U7tEyg4MifAMQMuxrpQzr9Xv3CptMOJs4iiE9nFqI7v9
uO53GY2M27+CixW1LoekTtgNJYispHhICuyBofqLA3Hi1jYP3UfmN5Lur+kSiFZSFDq4sNd1cr6Z
kVhUo0bUN1S+82owei3pTTnNHcyxa4hnUQbFjOH+9jfynQU3Dgels8Z7/EZY4M3pIZqaY6C37KSy
yKNJlmltWC2GS5YgChP7LWsD2qkAeVg0HE9oPPdHa2rRe29pQAWYXTnqt/XiAawHSL1fe+ARtqBu
6y6xhucDb+jOYkpKSsUTJ8MeZlU+P3KwncTFnuPRnTh1Qdf1r9Ggvwcqy8sT9y+VvOzkrGKslJDN
Enx/jMEYPzFb8p6chZn6o8UitF9AdrY5f4c4n/9/uy+3qYa+++rhRDHVNh5LGvt+wQnEu1m5cg4e
HN713fXZZq1vZq6w7WTnfbDG/SX6IPTB+AofOMdYAxp1fpBVed/Vn9NHAVVWy+91pozUIaLkyhvV
c1g4UaEsJuBa635wP2gNu+/1Q6ewIPhFGy0KQIFCnyHvXi6S7ZUvjKqdZ/PBqdjFCFdf2pIMwHMj
UPGCiuIXLJPD1nWqu/JqBN5WyjivbWTVMt7kOEhpMuTDzsLys78MmAdW2dqejrRj2ZrEbNa9hOPB
7aWRLkGUs7rbSUPOGD1ZDhU+1ArZna1HtSqkzhBEq3I0hfYuFYD2S5mHCAbz9BCae2XXrKBKyWSg
3BX4ibixZXCAumfH0ZUlO4Ht6HAtpL1Zo6K1B766hIkOuj6IqjPCVpBieO7I+WB1CFm2BylCoG24
6eaWaze06XEO9ThGyqSAKo7L7KfdtPTo3dSrFyc4ftlJebXOfpNM5uiLeyPbuVsVRQNYr99bdlFQ
3U8TgMAHSiTt0cFF/qf438qnO4dDrUWcdXyyUc9cM6az5IVZJ1doc24kfFuboyushxYylYOjZWgU
HDI55AYh0JzzlPq4HRA/+dIBduOmLFJ+wNgm+VAOsv78IWGJn3FGmwMCsjAPc3g6Vsut49uPAhax
Wm2jgIrY832ePmPZVzw3wJvaApsKM6qG4ttUSfrs6VjDHOkuByrQoyymC+JN5Q00U6qUNSu8lqne
Ii3CJj0g2SP4eCFyP/TRXzAVOawBNdLCnFIWTwTNIKT8XtuY9qfyQMHSvl4dskUddNV2tUID/sU7
jPkqn0wUWc7vYB7MbudGzr8nJXMYKRmRar21Je4oToLsUVo22reEqtOt7Rw/vno12QL0pUWu9mZn
cVXnFVTsma++trWT0qL8Levc7Bq2Rr5Ovfrh3th0MGSmykT7AsVeh/6AUm6i3XfEh5AxUpeJEYbq
TwJMNyTgSPBnr8Lw1r3SWqVDcUuwJYEZMpktujuZP7yLV5bKuQbvL7NUW2UnAZ9XXofhpbit3B9I
LdU+lorfSR+j6D4GKKph6RvsDVY7b5s0UrzN5CgLWCCn/5Eb4SnxILiyPeshKiPSrrAQtMvbH0mq
ILWEkhzrA1kDrJSHGCHWm3N3chEppVYKr1kOw9NlKUYJVClutMwTPMVpjDFI1ZUYg7LoGRObYgU/
EcxYsB8lS4gq3KAAmVPO8IlpOs7BCzFgxA87Y9vbNpkNWZDIawxCvdi5k9MfPOjmroZ7r/+0Ptpf
x3B/rg/aPJz4xteS+hq4G/QvaAtGfC9C3LIbdZUEg1UkBY2K00uGt0PpQJPGOv38HfR/mWLmMvBu
Lha79AaeTM6xxqcTwRlvheQAPDnnxyEvCOFCuxySV+eikrGI5GgazJEEBezt+wEMTKdZuoxGIrzV
EryNuKzVJ721QgM3EFGUIULMTHp7sZpX0MrM+0+r5JHzTefJgUX1GKZXHk/519OXvsI0R6qojX7M
eGFbPH81llqZsSSgBa2ZhZOJDA6LZd14bIOHB/yT2QJVzoW9JjwSz+xGNcVCHr8zQKYfD1AiuhrB
N9Nyo+udJmWsLvg7317Pab8EgowEErALQoNr3sSOe1xfFTTFIxb8uKCMQ33EBGxkZrZ31QxEDpLD
eXOwAzbKikA6SJH6SBRLe/lO3oKSh1Q4nQka1BKhcYClkPXa8L1qg3xjKJYC4hSt7iJcq93LqLl1
dSgWcpUe2UYYuH6ourWad2+BNczAwdqOnbhYSr4Z/ffXlZXTQiYWWQx/FT0PkPaemCSrs8jCpOYj
4aRUsJhWz1uxpsGPwrRWMR89pKSCKp9BGTE6wjTc/uOIJr0t0035fNPSHFOEcu5cUJC2EvOlOdjp
r2iHaosbvi6CrBO+tUw3Ajzj7pGsb/F/wj6bujj47NuRYp9w5xEvIXPpsfP13z/Bh1zF6U6o9Qw8
Lu79S4LKb4AbR27D9swcGr8G9TiNuW5c3qz9Uo6qpsfyd75j2cNEFAEMv6WBlvWdIBzCstmxHqIN
lKkp9PEz8KCndLdcD5Wr6jumL4QzTfa4vfrQ0G/RFh9M1DTaW3Zp3X/Q8/Rn7DR/1yx1S7eggG4P
m+0nFKAV36KhKZkH+Kc1OcN95kbadWRV9DcZ7sJfLusaUXzXWOQTTXIRsup2G4dezFDmzdEklW+D
Ji0Ut/exEbrPTzwBVN+4FNhEtqIv+UQH0swz1KHc9GSTU3M7g3tZHkyskT+9SOal6pCOQpgqApUZ
0vmqD5zIcCY636zBSMLe3+0fTDU0sISR9EA2LUkWfQkUG3Z1ShutVSPqKYc5q4RcjEWmdjfqTI1w
At7Llf1qK2S/RnTpm0tgNZafhZFUCvpX3ocGeku9eujE+JRab3PclHoovb8i/59HSto92snm7uM1
eNd8GBtOWz3CL6/PmuIgebLpsa9FB/63l6tGyZsUNvruHFNAVTn8xbx2USm4MiP2i0LwQcmylpJU
dGGnoGAJhwLOXpbYHYe1YxG/CbH7VWIr4G9d8sb3524jscje5AjnjwSTV7naGxYTED9G549riEzw
lCCENVRNYBSfxrMy9Ivk6R3vweZXDKG1ewb8YV20LzGJ+TYPiC84itKnkvx5hVigPN4HPvefAcWn
M3ax5eRbHrn/idi6ZKmsFgR0O4hArw48AAlo4jWtcksPTbkMSz0eZxV0A92u2vHVp22QdZsk+nlt
WGBu1LD0T/biGYeynWr1wyqdd204Z1kcLCyUP/qO5g3yxq51NCrWLJB481fCtYwx5cufZXWAuRzk
PaJ54OsF2aFhNelGQbH00L+4K7xtFNj4tUg6U2AwfNpoNrKzKbxj7CeVP73mMKNxrqtWUNMcoMio
tYa9mv6/9g/bqGGlcnJptZMjTmZ9DbyMmWLonJ99XxLu2LyZ3RLAkEOE/vj/g3KU1yhCW4v7lmkz
0CEOhNuGg0UX0jcbP+YTjT5MIgZBAwrAB6ybXMEHnzbZWVXuAKKy9l/JadjwMSooX0kUMW5HADEf
uj+EkwBe/d/8abg154N1MolzVtolaRvBTVg4N5tAmxmGo6vwNzfDw54bc1O9GgIDlQr1KYH+kzi7
Fm29bmONXXCwlRfx0ETgEFdkflid3lsC3if/e0Vhr6bUIycqVMaJF6ryiwnu0jaHZCNhZ0nnKAUe
N9VtaxsrYeBovUMdpbSifwB5ysZ/7KA7VisTG6v5wYUczSPdrRTdR+o5XXNItfHmuU+hJuYf+Pe+
Yx/jCicAh/Bty8X4y8DhGhxFfNqCAtXwp4o38gzhZ1xoyCT70M/5ilAJ1FYycd12R90LbhEhUU1w
XNmUaHKmAlCcDdRQZ9RxlU66vikTDD1uKv8pQbzsy9nSqKUQRt0lsk8EHMVKJ/IDxuaPfX3r6Qh+
EnQ6CpXqSpixjpf6uWCVA2180lftmk+O2HMx79+gfRzV3gTyXskXBo0ceBg0YD+o5aBTZY3Zmj9u
Y/bogmE69oVxj76D+EX1VDs8Xush5bzS3yAcDCz+hHTFwe4dHJ8PB0uv96ewKYb8lDxsLPINOQWg
+2Fa9Zk88rpGy2oEdQ1jAC7c2XpbAKE7w+oDW47QChHGPqIoN4dzLlodI/OsK29I7JltUOHVzjS2
wB9GtdjhfUfnjk0oSHFKffQvoPd7JmHoNcatnZ1cxuEznRH+FEf88LP+COmSJNQCNqc667KIjVv9
rH34zBCXIajVBxE72iVd0VrNR/y46mB4xA3zHEciXNQuh5GJYqEh7rS/TPQZM7Vwdm3nGjJGtpvp
sGT9bYiJbUq5eEuUDV6Kz6qiXzg9mewznG59kKb3a+3GsebCxPt026FzVK12w8BkSm7aXO9QK7IS
eIUxRVWJQ5XwCTcDrXGp3Iohun8mOl6ucdIr9Eovs5yw491pKZ4SLdp7ytv8Ce7zl+/kEixxpAV/
b2/qoMY0R1KJBSpaEFw3NLNY0BQPLjQAtucoU56xuE4f4gCQ6JZwXHIEtRc1N8yYteYxMXiWo4jR
ztiN4qR5QB+4dlI9PATnui6yyjJ0blxNbsFzWQNCzf6ZRL2RAyrsE8YZKJDjts5DHWbFOJhNXr1p
6YNp714V7VgZ7yo1g+Rf/NUN75wN8o32ITZ6i4g8H7cUbw+8AvQoLZaxgBDd4WryRnXHqbwY1ex6
/+vbtrh6dK4emu4vvT/9T0rlz3RKjn87qQh/C04arnIAc88/GHUBPl/VdxE5miCts4UrGUVUgmSm
mYMWabeGDTAXWvMTbrKki4ga/AHaxz4KFz5S5c8zvd8O/glhuxkoYkBVrxqsWlwHdy/zqMHIkSjJ
aaVe0aCeq9D10lI45ABhqvxVCHtHrpVNq2hl2gc0hYmbQmqEtNBe6rD6X8iyEVjuESVIfUgM7zld
9VVs3up0KRMLdwAiQz1P1gwqXOdjgvj6d7pSp8bZuUMQ5jqoM1oKST3fUep+aKefizxCQaf5D85n
IfLTin6BZirAlZThdXbfagWumBQ6ETGyOcwxr+xTvF90+qyC0a9eaEnsl+AfVxgp4snSve+2Hqek
jviZmUFxtiyuvjadsc+tcPxVZp4zMKDljndxsWnEyD6scP7XJOOrIZOfFlOnZdYmX2VLoONzGShj
kMpuPbL61nkwL8K2TIixV3seMYQJxU5mx0U//QsWFiheBU/0jQ8IjwkE4pGBQZgyiMwjHAsWGDUo
Ncv0py3dVgORKWC866URRwtWnd7Cl8+VXCv1c8JH9N2We+VgFiiFREjjquWwuwMQBAWgJkSDFn3O
Zazr62tpIYSVa1n6kcqRN1q5vtUTui1YWu90IvTyblvbxpqjHw3o1GuURQGHhqHCazcq2d204BBi
RzAFWbHLGeCI57ib1qdhGU6X6kpl+CgAZefLvWdS/PRSIUvEK5Qg0MFahUuYiAqxdUMfCzUSbYXe
6BlSBVFFYt665+QwBcq41QykE+Bya2g9eSwjkc/ewed6s8LCNz3nqrGEgVOINUpn+4UVGL2ucF5J
Pzu+buviIx3WpdRMa4Qu+uROKIZv5JqyXFn2FjJUDCRZYEUheYgGXUUMmOZn5R6BAWAdzYK7IaUx
kPnZvr1FdAXGfe+6xiRI05y7wioN59KSuuSbf6SXuuNGdIaA8d83gWKvi3i1mrOi1tqy8SKBkBkd
si7COAy44mgDWpzPxP659FgpYhZ8FZEvCjk836X8gnBMWWnYNZB9F04ZaS4QhrktsfywuUW5BYJb
UoppQAnzCkpBcV+Flqd0YY4ejyvEgbYqoY9Tjx0jQk5YHkw99qpc/3YaHBfuZb+dMSn5krorksEp
l0Ior0l4AhfMfITCwVAxLeHdm/4cgA3RUqAlM0DJdWNd8kfojmtsUV6r299t9LVOJWbZZEFDYK5+
M3lUgnJ3UPE+oHfjStqYMmuU6EE+fxGkyx2vQc9sUoi21pXxz7bQiQB9fVQHaUC2ryvyUVnX4UrU
TvuIuHkMUZm0b2Jif72APaTi0IKP96t7SGJintPlo837piq93kj3OBfuFHBqe+qDLCCWrUTljc94
qmPeehh1phnB7K0Plg6uMiWmDcjL25aESCp6oe8anB9uhN9lJfopmM94PxdWJzpOD6MgTZyb8VRE
AjRTuZNLyQZhDcZr+h8vAgNs83vlOHUxC81ZNK+QKuIvUMl1+l9zuRz1O191CZEFJdUViKlIPSp5
KAnvz8NIBPMpmYFnHMuUO9YkAX4WVapUx+SBGgKiMkclit/wa2HAxli9HI4QNCMV00jDajHz+5Yi
NwlGOhrcZXsVWIV2uINuASb6HZr7eRyDFT2NLWQpTFeV3kUrnXVp4knsMTGHOz9M/jlqm7KUAd8z
/HEgA8h70MEpAKuss2Qx+57suv7KK7+iRz02W+R5kzJHPjx0GCCQrFpKAjjyCWIZLReA2gdto8cm
dL/AMK+9xhmzAbGSXg79zndUn/bCyixseWLQ7GqU+aIeN+MFR8Fg24re2aSdqdnMwPOsuwSd/RK1
2ApfthqRur50kWIig62kBIkjTFoW0qHsv317FCRpchfGF7bN8h8blM6EGKn8jN3UmwyZJ9TJnExl
DLqDQBMoEsZTeQ/IC+Kg7IWmZE/O83g6tOTJx/To4agDcPJgCXpW7wcP7ECm4CKsESBhVnNzOJp5
H4ehIY0bo10sDtr/8ItrmdSZqfAnzQuhK4YfwSgYnkineqYoMwqptF3ylB6qBxsz8VekB7JXDh+r
Bffbx6CLOk/jXXezEB9bNGocQZ0ehh8dXF6O6Y0ClYsp78vHk9m/YUYGhbP4VL0U61Wkq+D1KklW
QeqQVCRGW9LvGWj7yDGNuBotCGyIA6HvvVwLGGnUq2wok0Mf/xA/pjzgsIf3ttWLyxufDqAJaJH8
JiqCiMUUFOKKsP0U7elfR3lCqaCNJHPiPozEfFcy7QLjhVDwlAT3ud+R9bnS+mVxb9lQy6cXARIq
sQ/jDR/d8RDB6FYKgZtSS3U+6AqR0m3tVQnTZDvSGSbBMaY4MEyB/lF+pdCxoFyOSpq6PN8fEpyw
PS0gdpIpXCYdwUf/2h4CLpcBm/QrIG+Us7r6oKt8CZ9CXFsICdz75gu8GeHGWBRHT/etqtl1W0/s
SZ0xhDb1x9WXu5YspEN5heJLVw68FRaK+ykc4n4RfPjlJKV8JyXe7oiAZu5XgUKTx9e5Fk/hdoGd
4GYOZXQup06RIkb/bYdEyRgccTUSTgR23wnjIfVQyZXPbiCzFwXftnJGYV+SXE4P/6IHOUcK8KUb
5qiF9XOiAFoihI0AnWSTcglx7iFmz8rlWgI3BkdsqOdkBhKcFLEEFeQXDt/XtBO8MuaC869GgiCM
RcTFZIFQOt3r5f1qqJek8KRzlQSMltqbF4nawR1lBrhJpTUdXDxw9Nl6bL6Dk2fmjabjLJfvFiT5
W1yd6knb8vTwyp3ueMjLqTyFHH3oanG1Z2i5uvZ0+FcyXl5iWkfhptJPPAvIdlUR9QmLSNqrkUBS
EzE5gPWfPW1+Cz6imSf2MQmz/7ak3n5tTPxggv76gWhk+UeyuPmvnB8OBcw5KHw/dnvrEP/KJADL
bs4LZ6GLmtdMy+zGVzn4W9+wss+iEroDeG9D+vnCMSykBZhD6YMt12ypi0YApnrtzKj90U1JSLVs
AZNkGbrpqbX293y90RzQ8Cpo5ZXjm89QyPU4zc7RjfkizxaF0rYW6ObvaglUM0FEZdFfbdl/XbP7
uTMSi/zRQdNWsKnG0vXbMaRh3yHut1EHmpKCi1MPwfFvb8tqIo0BL7b8UG2IOeHugxsS/MU86HWd
cdxpBj2Q1UYpV1er66ka+YK8oG3Xwaup6Exvo+WPhQskr5MDHGkL8FZu08GjPWYcIZ4/YOsdkL7M
GYWL0tihmQgdZkLOKkGfaQptWvXMIveRRl9Vnr9Eh/1gt16CkU3aSB8N5HAxWZ5FS+arRgML8wla
BgYyKPOKnzXzW42spDCfJ5fJyfvwv7u4Cctj/JemGSMyjsDj4nXM4dhNC9BVo2jHB/TOwnH2UJ+3
L1Y0AxdVWlqIsHMyR+IXoX7bbRsOUfYXefwy/dUMuor+WrkyzI/pEGHzlFcAvceAvWKOPa9ORnwk
yBhLScpNJPkFLtt8H8HGe8SqE3T2mGulc0BUlw1JbJgQ7PqNGz+t4yReoLGcAytF7nAWZvJihy0p
H8leAb129J725HvZzSpfAgaATvQPRcenwcBkojJCWuSwqawv0c3OPJnBzpVe9ytBKYxpcMUlW1WI
EI1bcBiP5B+jaJtEnroaAEJNFT1MsBm+Iuejug16VcPciph+q2aQql9v05wQnKy1SOuBKFNECtbI
Z485u/Uued22R6DfaXI4KkT8xnw38tRIqahLqixw5AKlWUe6MT6BPhiAiYHw1o1dUNSRcTMRgLtk
4BgtWgIeVbu36GThcghYr/huWxFjiYDmw093yOUSyhumBqvT58IM1Hwh/Cdt/HtPEySK3iDS7GHO
wSYh4kBIwGNqXTP5NDgrTDmU7gOpAC3WtfHWwhfWrdI/Q3UvG2NhdpzF4I+8uqVyg1qU/ewA73DL
QBR6TasIU4X8t01pRuzpAjsJ7ZWZEThXn11T9LeBN4b6IRvyX1nH95kki1ixABipP+I1fqcKTQO+
rtHhy2Xn+vHObN+ARcfKQqxBhK1+x03K8/5t651XPIB1DBGKrKg44tlmkqoiE/DZBc5gtbBPsBGH
KpowY+gCrHvLFkj5yEMrtM45DEbG+UWMnCOkh68cFJWn19eZL5n6FpoJZhlWFipmaEGhokb3UOa6
oLFQD1cbjHbfefnIYGLHyq11QSCLl/VL3lQpsHXYLRWMufx45OQbF6tQiUtaNprDagFIYcELGXXX
5Wz4nycLg/Br85803wMRRAD+4uDQEK6Iry41kwLAr2QAWnPkfEIfj1Q15/Zna6YPibtsmYBcQiVx
h+UcmA6rSIPxwMA+bI6X/PJ0zR+n3Y8yTOLeJGh9Xvlpv6PIV2ythD4fOeDlX73OkaZUhKHdKFRm
KC/YjWLiEs8X0WAN32IHtJH6APztdF+2UMIdqyqaI3mewRelJP4krpzcJbgyPJGBfYaDm3IGL/4H
dgJwX1DRjdfw+ibSpRVE/HeqZZI5HrXABnulE5cM0fiVpKbyxIlWJwRaWV5/LqOX9rRVAVrNpWND
P17PbrYgCEm3YQZoLv6uWhF7PpXNj/+v6rvSWOHLT2L3U4yP727R/GPWqUwCTzmHkiS0SQYyJcNE
AjzP4sP8LCflXimYGRD3S+T9oB6JNrI+cdPKQPEVGNZsGW/WkOyyvpxbL4NY/ybTRry7Jjo5DuwU
TuaAxQVuRPQVBR+2SVf+1rRpWKrviNbP/gGymokmlKn3a8S0v61UezjfUrBuTAoaBgMM5gknSFeI
1TxbUXIHKc6kC2S4nyloSJ+iKm4a80KodSeVaKfdoUDrtV4ZQ2H0sWM6nJIjHGT0cZWIb77SBBp5
FP5QD6ePEN7Q0JtiDfu9OKNKuo6zc1OYiV90rjEXGpj6W0u4EiX/6wKPbmk6JwgSHYfNgzmVQ4pa
TWPMqNfzVnNGv+soECBacdblNQ+2mqthkrbZx3dFnBao+EEGRYBCVFXQWQt5Q+p128uJ5SBJO3+4
l34WSWrV83/tu9+kk1huOxiqSqIL9yZQJUKbsG5g4I7NwIrC0D9sPImRC/U9kbOywueCplEZzy6K
45fwyYVUgGHZsHmjVB6bKK0Jxmbb2hJOiqz3MqtdTm3XiBcANTPrMA1GkSkRYfhVfZ99JiLUDuba
e/yCTdZTJwv/O9FBR3777EMZs72WWx1Pt/8gY9lTif1wIwkysyXJkXLHnwUk6D8u7Z49vlpgl4wI
cxsGsj9MuJFz83gcx4KWbQyRJYi8IgLXC0qEKs0At99z7XYo69InPWUsSkFuVaEXLTeNH3GnnOlK
SNLqGYwFEYQWobOw70vxyLjVmhK3pvxkHb/5YyD+Bnq3+oI6P5oJDvQYOZaWnC2WEKBKR4MiZ1dS
XfcETHN4jmA2ebVw2XKd5Azid15HmxK2llVcJOXLZmwBd+iHp4eqklLLWPIu9ycoy/7nQTuR8Hds
fLG01a8MY9fSrWryviOqmaOo86Tp4BUGR5jbsnfH0fIt7ObyY/SXg37IIaiRtWT/2+AWIzYrACfT
e3WVzLoxgO2i2+Co+DysDuCys1iYChEw2CYfGab7FiN3Et6Gfa5NyUaUeeWygM0TgU25/q/8DmDi
Y1/Jcxzc253MCqcmueuCyYSmN/p8S6nMGIAMcXJZ+9lUpjKZQqBuU886kX+0ZGkTJLYJcoTXdulc
KGvk+W3LauWXI1dz2l3WFatr1ZkkFYb672tlk6hunjLqf1/xYuBt4yFPeHesSt2XfNEkuyWCP2UH
tk3FAPrQ8yvA1ER0NCODRk+g2oKC2MwwSEpw4LTCki+cEHHbSjqv3nR3GJ76aXu0rVcXDguZSUC3
NkS8l3yjBLKgvbljRZ3aJhYKibBk8W0NaJHGuSDC7uwZYwqIqzoz3TvOXc9vnu9ddbkgXfkpwkPS
MqAg/uVGjQ/KKHPFpq6vkKjPc09yIuuT3EBoBsrClpPp7TXu8T7sjxQy4806S8eCYriC8zOZJZfa
6vFnI2FHkPIzYV7h1NCzHhZwGmwBWr7FRhdIt1P3oUnpPO7NeJ/d8KR/CDZt7SjLYLwm8xEaWaIM
elzko4Jnca+SV2tCU/sQy/eyLW6baiw+wbAZKIut4P5UTblftG7VQWouhngMy7ayiA8/cQl5oNEt
wWW+u/eXld99YNJTiZDEqB64aI0KmN43AYCSPe63oyxZTQvA8VoOcZA8aT91NV9JgULN6JmmYopw
lXJk0pSqIPKDg/pBFpu5tWPN0m+6046UkXPSbwftQGDTn7Pe/XL1OCvl/0VsHJczoCCL6d3viXLP
D2yfH3SrjF0MwPDOE0+x9S3tzrawLDMNrh/8Zg1qoSHDDZLUfytYhr+qiNgXunf7A8x/lvdkbA2R
HFqNg14dSEeiNBme5etgvdMduG17leKPK5ohZEuuBZfCHcgN88WMXwQ+bYicEoNqw7PC28XvOmAf
l0ZFPaoX/yWJBgWDb3GCEIN4d6pvq1gQThKvRR8mVTZgl+T66sOBoJWzJ7yGFEJOiUA+8N/P7FwO
cpgqy0EVPIGQi0qUaDqVCx7xsqGj7DiPliqEpnd46nGSE0U1OeqdVP56NxEWLa8ChBDTeNNzXCoQ
tEuiYJWwePn/217puXWaq4p4Z8ME1lIWU+Yu98bM3ZZfTu9egWkMdqbQ7ITIv6fD1LY3uk0jhMcZ
FtWkxJdjC0iMdvRcTH0tIOUBIBwTtMFal0jNialf1lCQHUhDcQQWMVM/KBmtDUHbFgIJIlfSwJKd
BPix9uUM/7QEyWW3jVDByMV3uOvpCkPjPkcI6egoN/qs8QGcDLCb787jvHJI3GtUoBmeFWj9HiOT
HyGAVQlaCNvc27qjWPEnOizyzWl7DA+zi8L01G0HX8TI5slDHAaWuojsahP9gc5xjKXn9/Wv0NGu
KSSBh35PaFtQfA/bTUBpNNNi/exv0ZbCM1ti71g5Q5IuyeauJg8iUslMfcBXbzD+vc/9NAqOeY53
MmmTivsWThZP8QafUQ+LKrbq1BDCSWaxcOjgwb9a4Icd8DxuAZmN2hrVKWOR5hwMRlS0c6hvAupP
UwS+bZm3vGOWCkzouweAkPLUVfVOryGRLOQz1G03yxG9tGNL3nii/tibp7frd9C8llHzt6+3IPOu
q5O9W8O0u+CC9h2FyuJUZLv9D9e6NLDXHpuDppcISZqIf5Qov34Va8yWXNKQtHCn5dfSMdK6IDF6
nwX7cGzq8uzPMkdUYxmNR1wsdZZ7+PORPuogsNFfYkoyIbh8zayIHIhSOyO1Q3JCnXl6eGFGZWUN
aqNnSM281Qvr2tUKNAE1Ne/DUH6tFKqm9R6W0kScWZbAznuEoLPtMg2Oe8Yl+vagrH+JP8kfSKIi
fhDvK2DXK2XxRochvxf9g3C+OldW0iBdp/eV70AQx7+8lbTxGGtieqvtIoOA4IvO+OPNF4VLgMhm
kr0BJ+4fTVBJm0GQYNqP9LMPh6qrXjpP9FLITM6HQL9W2Na75nTQRS1YSJJX2aXxcH8oZD6aZfGu
XBnuobzmC3AEDBsFtN0mUNizyAmZ4qrhzNvKGJjlk59YZ83RFDjUP/IPgZiDQmDngecQbonbHuBy
8YIa0bCLqwaGEuRDt48zxEEL7BecSD8r7f9NNt/WV2LwFJfvhlaHfUXiF8v4b1mYk1I8D0YjQJRI
1t0fi6KelcYEJ4D3PI8NZn49qPmkDFBAPmH6/qeiTOfaV8Mm+ZPoQ4Xhd9JIJ1T+iW1d1XCZ0ivZ
feTRc34bo1HV2Ket36dFBWO+T60KeIwtyVMWobtfoqGpUXVqJHuQPJrRSpgckeifbkTR/6QdlHeB
MiBNkEEu/xJ2ANfILuHV6MQaq/+4Bg4ZwBXaw1gdWYppnqVNoUcCUsbMRvM0Se8ZeOZjGsPOVYfI
XSAdU2d2mWj51mDCuZ2bCoBz9Z/xWLGl20RSwjcWhhkzyhICIKun7UdBkQOYcFIZEdZn5B+s2/m0
5S8nYcWhLOsxlV+pEEk4B5zVkmfe1cd8AMMKIJFZI3h64t3Pz4AFLoNFyz5RuRjAdkXrT7SeTDb+
6JxtO7lInFMPl4tW3/SZ+pRuH116oLIj1Mntr9BAWxGOfigajRi5yB6G7fqtJkVQ7f6FKbViI2U/
lXKinVoaijGwEdGCNc5SsZbl/lOxpHxzXbriZItaoeS7ZdyF7V9cr/OxoO4tfOhOvoZsEkVVABM1
Lck7roKJ5TTYtLZq8Llw5ap174ZIU+3z20McpuvyygF0JYCBTxPACtTGSZS+SYphqUDXZswAzWoJ
YC93bG7O5buEteyhLResvLB9As5etSZib2CNJxHoc/OIOdHpo7UvqCEkeFK6AP0sAoBRQZ1FJRCj
ILBqbOCXZZ8T6uzBF18R56VBMkyMEiWGqepB8M7bBpS4AJBk7AYYcC9ZBuk77Bj1UXObgSh1mSTf
P61m4nSnt36rxoE36C0TX05oTPjaWqe19Ej9as7gMN9uE22/xX9E5e/0BcUAUd3STvAgwUcuz0vt
WxGgZ0+3gU0OGGbEuQmPZVmKoCHsfw8szAACCUEVfK5qc/HQsM74OhvkpZ9RVqnfhPpgGxoOzd8U
ZW80BpS4fgy5u0qyWVfqf/NgVa2F1NBCpf208o5LbQQS5dxqODS8/u/OlobWu40i+tPRNfjzJweX
whnrEPNhRiUgQhJGh/V3hgmXYMKZJUtXqynLMbDiYdLTzYA7gwvdQxhDyBKRFF+TVYi5LridI7l+
6R8XvQT36rJt0lyNyXo4ELB6rCR1vuDK254ATsN99Ta5M9TyXJKMOphYf0KaEOt2Tfz7eE0s6ImN
QB5rjr4ii7QfQcxfE6AID2XJVlVIw2rBX6Id+fTX734LcG+D4ULgGCw8z/V1uPMJXSerM8Z2fCqb
J/ptv0oiEzW0x6uu/6PGahu29jgsxu9X771AY4LvJISkfG7PAgW2gxcSQvjr/T4eImXqhnDK9a1m
V23THGMu8torbCeaJ5WSVxJcy8x7YH/AfciNsyX6f+lTyfqmrTF+V8yoqXb+Msmss1cH8XRuFR9B
blf1na4Ny7JukTEaBFIuHgri4mi5zDjepqm/XGW3hBw8zP1CTHU0kJte3MH0b9FwPRDq2tXLZdhT
5VaR4Aj9hEmOZRBbHNryqggwWrTtxfOXB9c7pVCLbwcQjhyxe67J8mkKo+heQOukC632ERc5VZxE
WMiX5l6FKKEmVtUAGYDjbzwYehhvuawXl4+Jy0t0BjDa4ySTrsRkGGF+sl12p5uj7KnttIfjNjU3
uWQFQIzYcn8qS4J/geLOyOK6I/whUTfWBStjLE72CH+BTpsFmEtfn/Fru+IuYAb0OCv+pxRWqSx+
ADzzKA39XA5hkjVJbcyyftGTsn9erGUKyfau9O3caxBA8lkJzMxP+FmL+jRojQqXi+0ZZX7z+WwO
bz0nPCqCkbjNZ0Gngx12vqmobFAu6j8HHJn9+VvrpER8nNXj1RwHmTBWBKitAISiHBSvTgfMuH10
3sQGLz92jcNBFtgyLA7lPHf0ZOn3wnbMeM4V4riPpLkRU3eWZu7xzYH1rMhwB+hLFcBmQs4knZyp
xv/4QnvjCSND6JT7jBWbAetH19RCdiAMvmgHeZGnojQj/pZzmcGa8z/lRABIG9WuJMzuwHuinbRd
dhCF7nMh32/nyNbXWssqefrOIsePAFEAfrq6uFTOzr5CyrMMpqn6nSi0fHyxafwQb9Va+ISkURe6
RWf6NfOWeZvm5E+9dfs6l7FFKLp/JOnlT/FrH2VhpXs3EwnoWwBkiN1odW600n309kLHmRB5QIS0
5CUVeKYvsZipZoY8MuJRPEROcxnCwA+FXeMZIlHADwit9e16PITeOVzaspRAUpu57Ahw1d+COkBq
mgo4B8XnVRHrgSxcRYu+nacqAmz2mXbJ1wg9O3GoJWEXIOL5Owbin4Yh+Y11In4DREU/S3pPrZmq
8ZgV9l8Alx5sIWXsb4oPGE33ld/2xEXu0fx9gju1wiZcNVhoWARm469D6hLL+7DbfbRKf6dzlAzP
XqwrT799h2SyQFOdpJoxHzarKmgmqXGss3RBkze2LN9Wrb7zvbLoLdnNkYZBXPYfJd4qqQTW5/9U
fku+/7ejHOG2/jYxjJv4i5tG40qV5Ergl1b5O610k8Brt0/mZuCki/MPEYBsGyyCS2e4lAiWwcGF
JVZ7pWCfrQafvRI8vzjg7c//NzC4M7BaBtOvMle70tPu6wHXx2nJkzepHkqCq9b+Z2HLx1XfFmYt
fB07z/Pt8/RDsAu9O+qwYUheMvHj7bZeCdDq+sn3qDcIrw3iumVocPzyzWZqZyAo4a31G/BtlCQU
KC5MSk1Dhgq+SF+fZTAFDmFFDe56lhEI/ayX53zH/RiMQLvZtwnACPgiMhl0cXDQ6hPgbmsQBMN3
85EImlL9MVMveFD8JzWYImEhKGeV2nj26P+qBaYpK40zpgDQqN/emyz8W6ZZNLXW+gY/81ffSdMM
9zW4ZmjzzQ1Y6e4oadtUNI+UIsydaB5ecbx9Fs6L+PPhIpBl/8mdFYo+8p4zioFkA/XBnqSONK+q
ihbJb2IHJLkEO0dLuNuoM1kd4Q6ix8iEa3p++Ku076biHRlrdMFSrThAyctirxoSNI7Rai/5If5v
9uc2oeIrNYVrpFMLkybrrcWIQ7YgelT10EjQixsndeg4FKCsmxxaghJ8rfhCgv3rOC/BWwNFI1Pl
XVl5oSPUK34r+0YQBKOG4fdmmatGTaQjZOe5tudGmn9py0idmkiiRIy0PBh1GyfgFo4DmGaeUj1W
rR32uLleD/y2x5sbysLGqkzMoT2busAo74iS/g8614DFEwyDs0RaobBoz7qhsvEQtCkRkF7BnExF
wykCl+0RSU+/OAlKannwvjqWoJyk4eEB/4S5DAT4x0S+QAP3yQOIlqgwtlHWkGXBmPMEZ/7D2AOt
ekjT0np+olvd+N2CGyM7BaHgIklug8cqLQyejIsuP0jpVtcbo5WewCaVNcLvggn/eIpV+WTAAiNS
ILfn2G4raNLeco+nIce64XOvVrLYLfS5GGT+7cq+1vcyG+Un/xkDELVM4PmOZ1f+jZM8L12fFhqM
sY+J8Rf93UdboYhMcJ6ova+TRDcnsY70WPzLObth2U/HUmSy/yhNW+iPUmScaABj31ldgY83uXH/
F2A+ICBMP8jDF5hTacr+HkMx8zt1VRnqzNt3FfbbAmLDQ3Wrd1O8XnNgX9rXx0offoltKZbliJ6g
Tydgmbh9jth8fOpRZhuBQ72v4ukDvchNQFqFnsSLipwH8bv1JKjXTHYMqUxbE3VncXp8k5kL9R43
g4U2ESw6tWVr5mZaGkRUTi/OkaGvBqTnhotb1OlvppEw0P/457u+J8a3rF3B9QdhXbk0yK6OZ89/
PimIQ28/7LrHRoTxm/WP3H94B0H0Nq6Ru2nr1lun+jmYP4DUE7FrXl6cSNf56mIHWsOV2diICTMp
8asksrhVbdzeVdGFY7YQez92POljJPjhkeRzlLwqBOib5LTcaL5tTIC9q3N3JtPo0+hLoWY/edb/
rb+XZ0lTDnJHf3AxjSc1BmAbUot6YBgL0sVIBXFOXRXE5bxx8NLC2Q/+WFPlzpLOT7Q/EP4qZ5y1
dnU0V7x4ugUlXarC7uJR8BBSQxqIjaDXvEODHOBrMYo7VhYmfb4AkG7gZuX+rD+mxlmvPk63eZwu
55BAGNEFVHagZ7S4hEq6CECUYNw5KfQC6avNfXu1Jky5roXwiS6DvhrmPB4Zk0jOwroAwFyjSY/7
ecauOsqWL7P7SwMC1XDym0qCwPm7QAsA5tAyI/qjy3HgTAoKLg8k8n2VfOrA/+ORpPo7jTAFl0/4
v9/mwzALJwFzK7rl4UToxW1udF03+GQ9UKGGAsCihtUyTTuErwm6MGy36zGrZQqzo/ADrCceIbyC
b407FVWE1orFJMaKNqRDAwchm5ZBHfSPEVvaF1UJmBv+64rTvvc04RY3Ec5iyYhPX2fh5y/nyl/u
dU/UDjFp7WcitfrlYEKO1rLKuqIsp13UAB2AHJ69Plyoz6Rxlp/eEVHHoIJGyTZsOxOQWMOnX02g
YVGebGYMD+VqTy6lJZKKAOFi+fOhE5f8vXmu/da3a10l53VdHrypvgCEBGLZOFFAc62t16zHdduJ
KPTsIXLXc2JR390zQy48mopYUUu0OPaaOgtdqBT+9DDxDkhKM5voy/eoOZZs5OXtY9pCJ2w5ZWn2
jXfhakcdL6E0l+PPHJmrgNtdV8f6XtKBDtaz1u33v51ReziHupn9d4d4EfqTggIqg0m28jEi8I16
1/dfwzTIQfYVSMh54LfsP2hRvl4U9PA8jBk1+AGmFtn39weRHARQaHOHaeeqpyhvVm3P7KdJMZrJ
5CYk1npeZoemOovKIt1eBx71ODeXxsmf3tHnIfF+DOoPiEOKvVdc2zWxZzZJtliqtwTr/5hb/1w9
fn0BdqES6rDCNYze33WV91XDy1n1k9THYu8A1Kp+ATj8EM0CEWWuy/9zoYyk2qHcOgYuZ8up5+p3
jDvBYEBIcoNpJ9WS2dpcNK62adTbJg4aCYOP/jg/RuahuHlRBLwERJ3OYwP/N9ijhUZM/K2pD+e2
iVqio3TfRo3oCce868NYiVC1d1S81EpbNOS9/3BwjfInSi7cKPPxGA8UVeHO+pGmD10FrLSUdpte
lhAD7aHP9kCem7d4dUqmb44fZ2vr3g7mFf+8+uqukAfD7IxYHsBU30SVJ+BBLG9xanH4cbNAWZz6
XHWrd4yleWS/jOVwIJMGkXDE1NUnrH91dNqhwWYH66OPUfAxr0qhgXma+9ES7vPSr0kQgXvtRYA/
5W1viJmupdUBXHheJJ1OikjqiQyK5PnlRKKSpVJSXXWOuxPdIFyWA8R2ykqOGHATX9mpKgHTfhKN
NFLzvO5Thk7fEF8ekBqzW7ns2hT1LwhIymqJwiup3VmI8lrwZm/3zm5tFFE1PYpRYdxuqpoawItv
E7bxwzaRCyaMwVW6zhnay3SgkSkorSlbF1i1AH8+fbRaO/q54oz50LvkrftUdb+SvpFUMq0PFFuX
gzH7DV/jZzHLLFaTiF4YSuxQT8Kyl0EP2CSutEyIToPhVQVBffPoQHXSoRP+QnfyEb10p4DIv5FZ
T81LS021K/P46/VO4UuUgapgC97Hn0vWSI+XyDyDN+PZEMk2e014uN7AXStL4aDRGGVYjxLONuwd
yiNYlZ1JBVQpQ7XM8MztxS9jjek9pUH9xlW+1siY/A8XLgJL/OCG0g7NrqiLINstJsi7oYaRmBWC
Cs5QPi6Lk69m/i1Rqgl/FXdGgb29MukZ7L0cfJBj0AWzTmPMeFPQdsd0s2pZV4o1eOA0C+a8/La9
LlzvVI5STjur2C8QEWVJasuZ4XQwyWIghlu1Xj3XIj7aXeshus6PqND954KdFHSoM6B3BCJUSbYW
ASdt1T2TGtFsCDn3FHfk9xJuHzMRbKMJXU/RHVMnoE+ZGiD/JpdiyyHtI8twswzUDJIo9QrbZeiB
as4XWLmQkaPNEMYVcWLTrqhvq3AvgExyaZtJBLaHXxapFVEnIqrjmmDu/MdS1I8vzY8ad3RPs60m
fe7/wwaQr6vrqv8IIy9TcivGoYXtkqkt5fJA+0NuS1KUKng/MHq/ReDEuPqG06KJMmtc7Y3Hg/WJ
m7Ll/d2xNsqYuYJf40zeLo32E2TMGA/vTwOfleNDiuaYfSSCs65ilsgDDJ9B8h3VXWHrOqyFJhj5
raUx94tJlD/xO8dtQGOwYc5tymgBGY5O5EZacHTIA+VtGk920S8pGUNpqCWma7Ii0cxwnjeauSCs
X2Cub4jkShoPWltMogfj+UnJldXRME/FqoEBf8RbB1mTCAoJeTmdoMQKXnH9LtLwYq8+ZobXQh8t
2cGOGRdFX12b3bexHs4HkBJcOVGg5yjVgFe9LJdFYzO8YSceMlZAiToo/16L2M47QZbNXQvC7cMj
nlAByYjuV+dmmkEXKL+W4oBMydjnnJsF653YwWVUmBqaVAXQnQF8V760uJcasJjReEaM0HhN2R51
+7ZHe8VE7uZqsZGucyVMnKj8pxfWlPumt5Lv5PGWtR1dxCpyR9BOmaJ9GA4MqtVsnHA8stoMmZaM
wD5ppo6SwnMJ2UqMOJLeAfQjJH8mnhBUlvlJHL3dJuTAT/WYL28RKeO2XdAe4DS+SD9kSO8URk8w
4R6xTrcWfUkvm4HXqdR55rawqDPXkgjgF1fp9uskeDGwCsPTXB3g+zcpdKiUmh/kOO4mEXk0C/0R
NA0T7VJGjigB0tXk5ma8LJF5w6eOZykEJIGf3K5R9qq82J2T23mHmqON+liluBoN99TTf3dAYtyb
jN0f37JQIUHk9oyhp+QGs0EA2drovSZzXQLs6KKHa0gm3FhH5rM2HdX7lCOLbk8XnwKpwvIETzpK
BOMh/B+d7xQY2SfsFtp+wTTPJ2KTJuQeuxcOovpLHTtqCoknb5Sz5nmquGqtbKEpqmhz2hjZapZJ
aEO2tUe7/fLh2ciMufynp8hNF5iIxojNSt9CSZE0InHmscpZweKhTRF0iVHlY1ALU6rGeLp4UEwo
BEU6TBseOQq4OA25P7XtWZD1qdtwte+cro5vN+SldezL7DJYAYEygxpurXVn7wkyNG4iyC/ebgWa
5Pi6v2smkD824vgPszYyiNkqWdFyHEHJKvNpQk6OVEZaamfb5pPilx/pMIaY2Y80QjWDYZjr1XEY
buEoZSfpSpO39ao0VJyu7+b7M7FfJc/G2eybxo1j2N1sXb0yQ72jFt+TVolfzS/Xl49CcUF8NPNe
SWG5+zAJ+aFGh+RNszkYDJYVKcXfF9jhn9SXH/zY2Xno53NRrMYR3iNSGM/tkBIjNp8aNa7tpr6f
+bNx5/2warVOilq+2E5PLu1N8KIGAHXcwqiBDZR7Dxuonq9zjZkJGfmbzdqgAMBrmAL2ATPuuknw
AQWp7Mg6wui8qGjk0fqT9SiUnlwAsNHe444IQsGUG95kWYpILEVd5uFoPT/GWbY4aCOxdNgYq0w9
wvAYfbz4E0yb6Sq5bXIDohDEykjE11IeJ5PDJ2lZbO0wUDnyClVo/os98rTe5wyWLs137cRcXuVW
s+gbltJd2PRRg5/OufuggRae9M7QcxkLvVz3I0yiC/xblVLoe0PG3aeg0W/MK9cQSJtkjAb2qzj1
ybzDJ6p0dQVPe+bZ3NMHahf8z79NEiT/D3K/5gsWWYUyVkIAXbLDl6FGnBg5tMY1c/2UHZc+8BZs
GKhqAJFW3fnfQHcdTcW+XQ8FKLVC2VJ+BF9NZ5ZKcR0dij6oQX6fQhLyLbH9u89ImAJI3OYxWIa2
ATUrQ6PIZZL1fe6Du0cG642BL3fIaN4o5dp2xdLRaY4VtF4J8OjWlvmaawARh/sOzDB9MCPSTNMl
aXMCl75QXxdFQAKjYI9nOnd82KIt6rNTerxVzDcQCtSWpgein9os0Mhzp7Ro5zRGasB0/jrWy2x0
6MSpfpW8TUmwOKX5JJCThM5EUD0SRKpVM6CHWQc77TACLLw2U2yN53eT3FSQiAwysoJ1zLvuZwgr
guvR04eLCBT0Zjgvjfx8fV2GyhOn8hf14F8Ts6Jh3p2XijmWAHaIzJwEw4r8yyXDkcR0mHj4euaK
OiBVFHB/u5Ag0SKrxQACZhPbUA05l5WXUZ1nB2cdoLSlI/mQo1ZbWNnU2/KAJViUBZHC+Fs8vmMx
aPrW2+mCKRUlUxrutR58m/cOaFKQVlj2VnHYPDK2iQi2gN2NLAOlVWVWTS+prTQOQhW8rulsBwvO
8YAaV1SEXUdICVGyrDrxtEM2BWrcfQdxl6ZqLyv0YTTTAL+7b97kxspJLeI6Lv9dg2VyDkW1z+XF
mnIbaA7hmHWozcileuTSYZvI0dE7jE/Mxvzm2nNJ5UNLo04S2lYC0eRX3Jdxd87qpiTgPWnBp17R
yIunQGkMGjESU3mczPdEmBV1Bw5MP+I04Q7Ka5qeOAcwrifF3AwfrKkSvKcOJ24NsCPdmzJwHajH
FnNkbIYk85mjMWBmdzmOMQT4/h1RgCSdukR2ZGLtdtb4qWrDiyhS7CVZLyR3At5HWp7xvYPsV3zx
Zwa2ZIAvpXsWobxuZac9UtXQPpVYY1amvqVvkvZA8mM5i/oUFt7FA7xyWfEAgNHgLjcsd4Kh9xTR
9Ffsw2wmMkBKBOzHURUjSYbmBi1XDJKyyUetbsbtdWmSRFHdu9SmW1WlcAoTJD8jN3AiZhXIAXA5
yCetho1qkLaDLrYWurbh0f4FS+0eaXwvprQbmQkF1Pq7yeqne2y946ekJhkZEo3wT2ymWqi8hHJQ
ZJVQYj/GkMYQZY1a77cm2KceOfJCQHNX8JO8HvQi5C/TdJxSkx1z/651GqcE2GBg5ILOCWNdAxOH
M6Uvr3nKXGK6fzY/x01GvOCy7AigXiHrr8mTP8Wdl0LYv7RDBcLbkJG2lpGOBLLPuqSFjv67AIrg
zuqGrx+CC3ZlcJN6R2I2nAYYFyDE/iKlkkddAZKROewCDoAxwcDXoDG7neL1tNchZGY9+Jsz38RG
iYCofGmURnnvkHpLNDqPsC3Z4cdHRBI9na8iwvU2hyh/G98BPwBFlz64AgLFSj96cqfPQVj5g8Oa
FL9w5cmMQ7MDrt6ST8tHrLRMKDWpR5/9hWTRpySqO9mae0arS6bidYgBYrVNWydRzhrhttJEmNvv
smXUpfplTwC8E90uqEg9OLcQ0tGrb2lEH8UE1t8AwzfOtnk7iTsRpShjrDBNfElG1oEjqzbMLJVL
i7lr9NrqeWFn0leKHylNJxu1PZh3Ov4cLcpIu9gvgydrkNJunZmosBQxdop09mc347rbS5x3S6yn
9adzE+GvB5hOZ30gQ9z4G12CaJ78SBxx/iVEW56PYk2OANbfqdEFrktdMopayO6+Z1MEOAB7J4sg
hGftzgn0SAjT8ufjAOwHy7BlCGMfSoiVGWMrO+psJ9y2wRC+1HBHgXBEE47k98/Wst8LmJPLvo01
0YlqvZ/C09uGaBL5C/R4WIgwWBualqMF9eSKmW5DeB9lrsqUBH8wJ+AxZgmV+prcikWilJNo6aTZ
NJKruW1E0Onm7jzuwe/l0T8/ufJnKQyZ/DmpS1zlaiELmc8/Ng2pXhR7p0GqfkC4SElR7cOPpDmU
kh4qD8TcLxe/fHOlSTVyXvPxTLmZswCa6HGP8qQk+GvZMrGfF1ROS0t1EoEmFhMF/6GYlybugN0B
8gltTQtkgWVetnKS+8Z5CNBe5XghSvAKlDUNyr+/O5y/rJpU1W3C5jDmGmYEMGxOAthACI6eS/VB
GgIycDKiznro6EhRBOm0SeCw/zGBBPu3xXs44ui1Mnti0HZex4HSuiNvpje89nV5aTcDXCn8vROZ
f+gLsK+lOt4yDlJQc4oRTF8lGciseob+QnMQKayGiNt3RXvzqpNhL9z13wa4x0ksCowTgS1gYkzs
sHFdp/cZ6A1YnNqDtjrrhwuJgG86PSrPxW8oZhH0Vbml9cXJw/X1EybNX16tyTZcJ2SgFaaIJLlj
T7Lm0x+Ax26SOtIpfntlLvljujlSWY4Nr1Vy9rku2tCUFcGHM9r84tMaGG5D9C7nBqIoB5IzKivo
DooIHVzQjogKpr0+dOQd8eoitILim35tZZkbmCzXT0LXDdfq64WWfnHYmLjH3M+gS46WmDyEWBul
sPbE8uV0L16Ct+lpC8TpK+h/s+HnXs8hFpl3env0i11tsvQR7gnjJtFe2qcYGnLqMyHkkGWdqgbA
2rPoGTD63NiPD4ntuzvkWqz/Hh2FmfHT4d7FaNUNusTUd+q86veCaT7fL/GW61zDN9L/VgNoe3hT
slc9acouqsmEfWtG0D3vBISD+3/0NaJnVOPBMA9DXJ/8R/nwJ4Ax9x6ovlecYC86WTlFvTSsHSp6
5fSL9ZnHHmUbqj8xMq77pGWYelxvgFHWO2RsJs2Kwe3woPPlbFdBo+F3VtILv5HOSj+lIY5/um38
clMFiEJ+6Utt6bXA/SjFJ4HQAz0Mm9LfhVtJm5cbM9c1ACugrqhI92ym9et5Kl24UfB2JJe4YutR
eJgkYxzX7gxFiD0GWhs3skSCP3nBalPds7VaMyG/A7boXC+SAeSvDxrhkVZNJgs1lv5Whj1JvrfD
QfORs2uPDfBGbNUIV4ghwjxzr/FheZohi90fdR4q29R5gNp3/PdozAXXNWz9B9wVE5j7hSoe+uyn
75FLB+/NL0f5IfWVie47cZToBwjxUijpZY71tgCgkGH8wdVtmauQ+zCy2IBPapsi2puMCo1ae6lE
0uoM7q/hAuzx1mhakjhvvsFc3ud25Y1hnnK3gCvPPMtQ2cV3GlQ9ZZvV8H1qtembeNdUv7Ze0JPH
uZNerDARo+SOZGyYpe6IJs7J9WFV4UZzLhkrU92mbZNPNJAdoQcrlicoR3330nJa9prEZZAtZDTP
dIWz95Q4A6R4VWMn8Vc2N2S6pxNG/ru1AZEyrJdUPPKJg3+Yu7TOQGpjbGWw4GujtA0UAenqZ4mE
/BTZDmD2pRn+Mwh2OZ7gc1maE4ocrqfjHa/GNmdnfgk120SgC6GeDVpKZRxZ7/U7TgeGqyC2KevG
SwmWUnjN1tqF9oRt6n8DrIxUKJAmbDOipzL/mZ4FdV/bvyHdzXAmbwFQBrOrnVsXL+MKKAI/1Xv2
gKatAFBxUvfZJeYJaNQ4zlIMmYKUNWsiNatXB4V5IQ4/Dk6esD9Rxa5ggodP8jAH4yutssRaW2Ki
kdP1z+CbJyG4K7ol0ogRYpFT/8evu/wxYR4DSZ/0jbDAKUBWU7qPZQ07UCkha/zMyl4s4AtUVfZv
HiLelfqyp5AviLZdqc9PmqN9r2gqc9fTWgXlE7Hf4d3toAM1x+/Ted1N8/dXjZhSxrcLnqjW8edd
YWdQeQucnA8IjQRS1lRPvehqiIgAVluapw2WLWpX2GYTepP0QI6zsXwXVymzk3saV18kB0wFafVu
GKd3ZEds6f3fZWev0abUzRREoNWdntMrzycM1FNStPRB8pDf031NbQEN5hbI3UZuXU0BLL8LzEPj
53kXHuLAe9QOGDoy2mOAZYAqAq9j6F3z/l/sCD4+iyjNqx/LTaN29X2Z2+LgMGnIm45L3OfTPNTL
ZkHcPJMDes9LW3V9F7Na/Fp/5OlOhedz7OAouUBJEkf3SILsjKZ5v8Qd7IIrBA9dDg6oC5vQk9yJ
FlVR7Pb1oRryG5s+YgvqZVPOiG46jlrxExrgyOFZBKFrjJX2kdhYIBX7RgGrxh3nYCx732iJ8ExT
w17oO3gGDrO1+a2lqigyIAm2+erfqZ5ZBf76IPiCrGmTibN6Ql1ZQS49iNI5WttPmCdB87G2PqZq
/NQ4e1QTGH+ghjpWVZWfSHPuUtPzjAlc92tvz7AyubS+eg1RmvwWUsD//e/Z2we7RB6BqVusFfqo
MrfLO9aPoAE3z4GRNvx5iz6Ap8YKLImRUogIIpsn7CuybI+Q1gM9hAtR6L+7GhXFpU8yFduPvcmR
PH3PmHUKDmVpqZekutINnj0CFDDuLFW3PTAVFnPYk4f0N4MVq0IqEiHkdemA8txIYUVCyECQZ2sH
xD9CsoYXkKC5EzTgjgcFwRYg+EWemG80o4iu9NsH/gtziNhqF0EDILjr6am2mnsugnMaAuF9qa38
J6jsgLrAlhMT0rWlsJs8kqRNy/gNCnXL9i64W6BbZbLrXR3TIyLUEOY/5CHGjfZO4HZ9+Szf+l/H
HtO4+kr1wANV85Hp42dySG7lwCwgvpnSzFGTzqT9eS/un6L+14CcLdi/aTeX/dx/wR7Sfcs75zRN
w55a82Fe3UD+icxakhJ2dcofcXrtIojEwGFZaX1QrG12VprRnyuBeleoaj0ar2Vh6mUePS04UWUV
vtLWDT4wof48XYpW3Bl6qoBHBnHOV6jm6RKuV7RhiBgHqkLX04U8rYd2UVpg/DwU86Cz1z6mGfaZ
DaaQ7nm1+BB63GulKygre9XLdgK1GTrT4v5/pi9u4YVy63TiqKZMJRXoZPxQAcXd35+2c/2tzLyC
VfkLn2FYgc9B5KOKoWS+FsLxEqgy2EuSFnGnmne14WOXOrHx85TQUoLsiB2ETvmnANyKbmvmAERJ
Eo6zXd3vf6O+OFdE8RFL90DcL7RuO3GO/lleOXL8hoxDGhtEu0Lasc2uFTwrUXa3vn600GFwrtkI
WOZbvVvOFa/9q7PaA22AGAKKddrQd55l6v0w2+Vf0nz+SbTfzZYBpxtLdYOPE6xJOSY1rz6xgno3
BhoxAFaOrqW+i0gq7gdktudTMQFAT2v2RJu9CA9dpVQd024ELVFv2txS1zZd26E9O+cMCCbD/WSh
fSRkccyAEJiwDsI28Zk4/Z6G+/NBxaywhSEJZd+3j/Gp41JKMeGON55x9ylsyfJCYZEYU8b15MBs
hiqAmdAQ16pXMgxXxXwEFOB1H/Pr0npcst7+mzDe4uFm3CUGaBt0Qac5j/If5KlPNxVUq/p47tuV
e8501cfbb/U5lXGxM7EvJrNUTTmQnCmH0m6OB0kbNYwGYfaaigr1fE/EA8+TjhkS3eD6eqMyrHin
MZWBBD4S74DWj493NyyVOAbbyuzW9IR4OMsqONKmnhQdXsVu/20HELxHW9o9sAGd2OB1HS/VtM/l
j8wOtTAgAqlt6Yzo7NizBDblA0CxbaRcJl5RQOpUkUqhfgeOU8hQrB1Qj1tfpG+dstjRpz4Te5rV
bvjstoXkWJYcAc//Fk3DPcwkXjBpnTsT/94jpKnS0Y+JWNEWIlOJR3lh17tikegXZwBuyXdW+1Yv
bfygF4zxF4XzJhZ74R+9qRmo+Gh40WVmulIDU697EoqBws2RSLbAbjCnT3rexMaT2oislS4CBWs7
fXGK/r4LEUNudaA+ON0urfNEbgnP2rdIlEbs0zz2zP5rk/A7ptVgf4tSM3HScktvGpG9tt77bPTk
cBL8PbjLRWDlBhuUeNyiZbLJSElNvqmjaKZ/yO8BTqPRCOQHZJYp4uZKXNloudHaOCwmwjCN9+6n
EmyA427gDlUXtCotMv4xY++U2DimHHpXKX7iaykDvkaZ+RyKAQW9PU2G/akdMjbGEYkQ78cVyIYG
rj+LwSaDVIBKWYwICzumbzJBAa0qSduRhjSdyiaUEeHhueckG2t0i9WtwNk/FpXmQ937yiWF/BpU
y0cEhWwtm3ffrT7RiDUoQbzHRS+fQd/gXcA/di1pPDR1ShRfkewGPnJa7JcLEj2gpvcwEU7v5WhQ
E6FUQXAGmd1+6lb1jVJ8ky7oBoeVMCoIoI3V1DcfmnOAWTzvYl3qYLUH2ClP1mhGPdlf8MlL6ohE
0BWKYTd+0JrU/MaZ+8QGLQhaLTU4yAHaZ2LHstASZl/vSIP1Hn1etnEASeoTKbF3VcQk0OnqE93a
fbQd1dr5CEabHvKBNNK4lijmPCVlTc46nZVN/XP2YDNzQJeiQzkaa37QNEcXYIS4djBECBTGD3MO
vWbdn39JeX5rkfVULbqJ6l0OemPyyMExz9zIq/WpgCrDtPtBexo0BllK2N6nfA9PWHyIvwirQbM7
QJXyb9gmi2fRN6xcciEdtOX6V0Emuqpgc4EgTGYiOBkRDy93PAKtKoiYSeEhQIaKIZExb6RuJ1Gn
gjAEz2gwyvPsLZuqaOk1AqpQpOvwzrSd4NAmkP/3ggCG5kXrybpnwCyJG6/5pVrLhZWt7xVnP187
CwzM0GV9/ABNk5sOcaXoe4Fon2jhWH5BNuxbfqlgnoU+5unPDK24D0i/cWThFmUmCgPZP0xeeD1S
6Gci3kkM6deoU1+VK/d/qbDud3lS3gZlI2xw6GfYLbwAg3qNJSwVWJeHdCDJGG986Sided3kowEf
Mk6T9sWgPErZJDaiVxRjHUpLRigRuiBoZDcwO08hPNxpFi7D0QaGQYL2neHih1vNF1ckvf+mtwUq
VxvzDATgqpLc5rrvu4J3bSJKDqLkN0uacLhbQLwZmSHTXEF7lUfpaWrWSJ/Na+mXSVmQFfKFcBNC
UlXGoAUAG0mtuJLtvf7mihVSQ9q4Oqnfctxit1wkJnJEgrhnoT1iVTxcbAlHPihaslctM+19HVBg
5f6+4aFzl9CztmT2rvkHev/yp8ecBrGW80cH5P4mn8wi5HjjdnZNEFJyIh7mdAfnDF+KD3Fx1Lii
iU6IcqW34w1Cu67qCWJ8vxGuJ5JZCJwmNpqxeS4dds0QyYy+XC+wDGirQKYUVT2Q85uOMKUemp27
s/bvJnuHs+htYTLC4PPt8zUazPfXrqHm2kaXvhod4rW1Fs7RBwstVgwMdUct4JDijV7wlmiODni4
SCdOmMOVXI2Ba3lcO5ebH5g7sPB1j48g5HX4E7AZj6fLsOqzf5oPFOO+KS9MXDorYk06fDoK6JE1
rNBt5i6LCT+Z+balrBk7mV7m/Ld6X5Yh6pdIFGu/V0sq3541k4GqMyI0ks63C1RzS67mGB421UlZ
i8jqCVIa+wKrLVB2maPd2CB5AZdqyFfiYOc+d4elWd9CFx8gXlrvpcVayMipMmzs882ySb94dBnM
aegVn8OppsojaUu/AHLTka5HHddh7gI2AMniZ/wYnj5sl9djxQBBgwvaMhC4V1b74HSr030JwDll
m8Kh2Xn0HS55c7BK5tVAlJ/yheWGRmH1P5juE/+AjF5WROROzvrxXTsujm79GmvkvNdWNXFrpu43
ntaJsfmxIotNMCYEA80tATe+hdNgvzqVwLnp8Qx5Ru1f/jXlMZJ5ouXmRDQfdpa8jzMFeSNgD8oh
jhlEufPv91rH7H6B4eRoNyirYFNwliP3+yDni61/owFemTjszJP7aEKMnqRft8ExcokuICXAVGw8
0gr2wwKThswv+XutontMf22H0KsS619Z+/6d2w0Rcs6QhI1qnMTDLyjRldOSKW4AC2yCgaGHKfYM
yhNCtUHrUpGY0rlg264cnQ+Noc8se/NzpCOHThE5wyP1quBOqFMzXAIIWIL2LpFge+oGKbKfvw88
XsprHrlWeRyJIbcCaU49T/hbZmOHgw0LTwwKDowwFhdhFAQURyhfOKUKAICk/5NPpV8TlOtdq1yg
Gv/zEI0CZHRUIgEhDlLDoqPHqhiIT5CJjhw8ZlxHMXn8zk5dyKsLpi8X6+5mcImut2OTH1o92h7J
AOefkhyY4wAYjVv96nSB425rsTa99MUwePxi5FXw34uTaa29bEECsOwnyaomiqulIyaykS6zEhZx
v1qd9ZltBLXscRQu3b8Q3R+iCcCpaihpodZJZcvHYrjJRAj7Xly3LYOyT9Dbp7fTwVQoxJIf8xYg
Q3MSJz+cZAAvZU/Tx58f4DGNeD2fK5ZthI5K5+I09Kqf828Glz1dChX5NrEn7tWK0yJduNGiYaZm
oC/sz4dUcSSlqPjAZReR3PPBRHP9meEKp9XhYkslnwjdB2fiSr0LYy60LkOQT+9hePHBez2y1i85
M/OaMQ2MLgnLWuqWXLsfWd2vXv9K5T6VIuvVIwguqjMN4ucN280Tux7uD9FD6t7rZXiDl6o65cUP
PI69m23yamawbaJDOZAupwAaZ7sT8HMkY1VRuPrDwG0f4NvE4rP5VVeziazUQ0eyxVsH1VRt+pER
DeapIAx5S/QgM6g1E6ldXbmVevNKIHQHQ66YWp2oZXbEBldjEXObSR7cUi4rm0xkpV34jI4cvazY
WKJopoLaO5jZaRDeBXhUpVst1UbVvaBiUqilEV1+3ABjEhkEbnpvYW6/jR5OT2QCKczghOcu56KG
f0QXIKnorhgzplEoR4jIMnoI6lfDRaRs70lF8kIHGapg2d8LOLX76m37bAtO/wTMwXKWNlxtct4Y
2IFW6hYA8SGUKfQ4XIYxCLN7nnNELqKRyRhX9ZwLEI0R9Eb2pMz7XGCiwVwug67D3YtuyV3/jVVA
WyNr7xaXBBmeHyONE7/rOQq9tAfz6VdCBXGZarhFuScWsAMrn3/WdXeFs6OWr/1R2XTWXq7tN9VF
705d4HdSB4LmhF/fSFxDw6q+P5llYugAKbPrFagSfuCsC5GGI1EGDRIu7+HaQV5upV8puH1ZNvkQ
dPGTyy/24WEJD8dmFFebUuvrTdPykqc/IyZ8XChfRkhiUKQdJ3G4O5S6z0hVwnVkdMyxbot3PdA/
DHV8oPAriKol6qbAToBgBI0q7NqgwgIrSFRJRk7UjsN2HelFbrDQniGInulyxyqriwuBcOmoX9hI
LVua9JKz+qEVTgDrjv5489n8RPCKwCJd7xQ+pSwtJZoxghscV+JRM0yPbdHuDWO7OGYz58wrOTYy
+ceWMi2r7nLhCH3pPZVW9PQGrNq/OxmAxBTMosov4eUFNolHBdi+0yB3ohT2eRrMGsvlCni5C5al
Kjwj+LRY+TLGZtj/+IHfcR+KpjWyXSug/eRavzL9nyAgM5oZcdoBi+KoK5DnmJrGdIrqr6IbDLtc
K7E/UX39d28I/xtz8nNak+km0vl+gwwKWhA7CvG+dfdgACvX6DqnmjfERmdd0Fd4Zy9HizVWy9nB
AvFtu5rk81XNp8TIDNH1Ux7ntdYk9ByhRzoFQNZJVcdfHj9+S26B7oirENr9bdzKNDZ9Rtww1D/0
hC3Fmo77gS2YKLUXRXgyarto+KGeg8rZhU2ZdCOsKNNK5Hh0Ox51GODtBTCjhDOZIoM7QBJc7yw8
e8M/Q3XpG8LMZ4IiPyTu9iyPfwjtNpFW6P5FU5Kbes1nUVGBDZ6BHK9YZuetRTOFf177ZHoHQaxS
Iec5l6C0v4tr0OvJkU930rJ+VbTuf0edsmEReBOgxp1D7lG4MNpPPsaWuPxzUYjHntRJJpn5/o0M
GFUpjfLOvVxwUfmql8lm1t061GQh9XFmvtQolx5wCsrQis2lFMKU1naFVyEdhy4cvXpgqiPpVGLS
kZeeM6IrKAtDchUMAJb17ihmXva1epgKu1sw9BxUkOnFQJDEc09pSwEt6KUfOkYaBTpNEUpdzOhb
8bEPEmCMLeQMgCXNybN/h/s7opd17REj/JQXpUo2K6JVhIsxlNwTscit2keXfZxX368fLDkJ+IK4
c0l7KkblJ3MxNyhqAL29Mv1uwXGWHVqge7IGyQbZIxVBdx6cpk5s/6Pe01vieuslxtF0lzj6evPW
pRbZ8KEM6MOsVMUav9NIKmIDeuGey5QAESVJneJ0alvvPMlCnjzOwrapNghr2SPp1l+ltbWAhTme
lrfLYoCmdHfacLbL/35T4XGHouYISmhXnh3INpIMy4L65Tn0m76pmuF2cWmjyIu4I1D754nz5tpW
gyJNd7l5JvYtzS/znvyeiMIUXG6OkAG4Ze5EaLjrFa+PrHUuoAAJZjYbzcTxGXhJ4nU88ZwcVMID
Y7taGxGOxOO1MsmNBNf9eTa3GexM5UXXuFLK35MXWDegKbbk6/jamorwJnuu9aNt7u+DFbB6jo7W
lS7cvxWhVzBuR4QdjTYENa/U07m2DesGsqA1DeKVl0aKFtkgcMJYXYgHBFkraGLBCrR+2nkSURUy
SXUcgWaSa14l0C46Sb4IpZRsdQXLFwJb02Hvuwf2MSA7zW/LUmcmPE1ng+h+4qv6dJvGVlLnyl4S
Cmj5pQWVrff0wQsEFojVI4gVbiUeIhcmfQHwTB8gdDe/HEiTYLwVtVL5T7NSRcGDIsYGE8IIOmo6
pVoBthPtv36p1WGolNN18RTQ5iu8TVOug39pqTOGzXXtoyuGY0nmBw/X/SF2HveoP/UqCeiEwXHU
tuO9zlhCiOpEAM4WorUMy18PJPfi67+J8wc/2l/bYRiZRo07Ji3Mn4oKcFp2sB4BCUHRStZbxRUh
kjn0f+XJMUkqd7Z8/izH2f2m0reY7U9L7tvzRXfzALob7iBurxOkD86AqdrDjCqMTKn6fRZNZBhs
rgcLhAk866Us8KndSn5L2nuptZa1Bk+Wa+6GXoWqv76BbNusuXDf+2x1FH9n0NVv6X/FigUKQ0xi
I5vfAKkTRxCF3ysmHXu0PKyJD2+pDhDCiOD5sJ6Pvfy6870S2qO/Np8sjxF7tnmFn5ggkJzIiolE
9u1u2LYzIKAQAwIJ6Dk9Fmp+e1Qux/HsD5NgcycMYJRtu1o8ObUTTqgHxP4EXnkRrR3Y200HcpbS
mbrfFzaBT+9HOQEFp9al8wmJ2p21Dpcdw9NM4kqIp6UqkQ2GCd+l9HBfB5c93UGKJtml71ITw6J3
gzokkQpsjn/AjkzkEwkyaF02ZvVKY9DSxcqK2XM4nWwBL3KdlwGcR2KdGRCfu4B/5fwzEdJuLEbj
vAV0g8ggxZ+Y9F4JnfhnQSs0OG1Wmazgq4puRb2y0V7JCJx7aT3AILVR7VmFfQpX0R0EhppJ8gQK
0IguLdqv5LrQZaFo6CbnlYaemNUZs3wY3AaYXhpZoh0JNkqgYv2tlPSIjp1qPhsYBPqkTcmpwTTs
+Am3dI1wv09tKBFqBZCAMK3kVAePyJifHiDqLU/r5glvvt8dj9rEpnSnQqui1qgYNNhftpd/Bu3E
W0PV/Wm+1mw3jracMamaBKADyWsyf+vQbigNOdx90OxrqLmkTqNMWkRaHuJ1aB7iFrvYghgmpMGA
t7TvJGBcrD2reyISou8+oF7xdB91+MR/3PBUrCoLOxLD+Zz9NtyqRgQdd8wjIFa1OgUaAM47qjW5
/XaXNh77+qZrvqQ4kRkB4ok6wtFrgYG4NX0JrpAW8I9u7ZtoGyTD0Qwe9k6yu5fRbkBhcHSQ9Aao
3FniAJe7cGIVfFrR5Gnf2PceAXd4aRYdCRb3+Vn4L0H4gHwjwSb3MVVzn3YkGZhbhQqApu5Hi+6Z
mgMBcWfhzRd9u2iuqvxYY3P1ZFGkrG3a9Vk7rgX0SsbxoMlsgfNRd5i0Jlo++ZvF0QVIkhYlrYid
NroLfOJzOkX7zsOByVpIRyGPMHWe2Ys23fMY2AdVRlID3ebABXpdoNFHgYdhYYfoJEu9bJiIrNeU
5Uomv+0ws4xHwCKWK3B3WVF4eG1w7HouElJtd0XQXlnQEzAWJnjXfxU2G+r6tMZXee4piWYAtDU8
iHiAgTPQChJVRAW7olrQ2LBFdUxAiZFnGyXNqtVXMMtsfyFaF6m3lVRT6vMn77MN1dkjfMSVsQaV
nI8/ETL+Y4QFl1lIkjYjU9Hc0f+1UsYq+t2usSYDbNOU4NsAYTpaVu3jG1HZ6jPlvOeN6MW/kS/4
7YB+bgPbhnRmbyII1OrhLdQBmCB5QeadIVF6KSfZDCDdatE2q89oS/JKqLKRFbWUeIKgxkv35mIy
On3RZGISTrt1e9abqDXvQFTvC5FWmFlI2DX8/0WnkmH5tK3FKqR23mcmXXh/PlsNoeaEadB4od/H
OViLqWnJLydbnlxfliLOyWi/XTVhaSlkKDrmFmznivHB9Pnlv2e3K/g8TO5a9rYue4yIPqERHDfk
+9sst6DNnW9RHdyCyaX6Q1VGd3AsI2cQ0GaUNUUxeyn+UERJcHvDaWvPbQt4xIIKx/7qADVC9o2S
cXGmrSCJnSbPpCksM6BediSb6xizf8oimB6B6W1XSBo8Njax5lGJnzC7K5odg5Ve4Cv85Z0AOb3d
go9FBJH4MQRWoXAxY0W64Snxop8N6PCh5jJZSjX8y6Y/uoNza4rkOR8WAoWVIJm2CKf/m4jv5iuY
s30wdBfI6r283KWiESMzY6A63OnDZoaQi8V1eFi+DK8QnBv8RmeY99Ds5lT2xaC1yzBRgUezKPWc
K+NRcrpmsJgvngMF9YrA3qt5QEnHJFGayrzYFJjuRtr+ldaoxON1pm1avmLtEqaRYgN89ihAbcTt
3HuXjmQClpBSpnKCzqGkza9F9J1IV7ZY0OJL5Y70ZKtk/ANP9qvIQ/fAJyOxY+CleIGuh9neWM1Q
2CcBG1mFNkzeiuEuVlSmp+lQBELMJDqEiC9VNkHgCSYcKftYIfHL71ZL0k2wWGe5mjUWYigqhi0R
4hDNDZAvwPB+K+m4skNWj2tQr7NOkPzqxzP7zs8pshmy+qCEVbMXi28V2gipp0iyL0qqgjpyr3Fy
Z+fDxYYflPjFP0in3CWNwtm/L/F8/SjSOqplGGwrTwqAkxizVMs1yB833qb2n+hrS0m5pcSdDKJQ
O3+0c/r8p9E9OlQCpIyVPtd5qPEcTnIOFL8xOG+92IMBPMRUdfstgntpayCZBYoXs360UfmI+m/p
AwDjz38hTIXoHmc3hl2VqVe8ifOmaiQECltaDs/kvUtm5FTY78hoJSUNeWSB1HSlHvmP3JSjc+s8
e6TKlMjRpvC2AcV/OTq+1aUAHXYr0yAbd2U/vhpndO06JCN5zAGyGQdNtGFkHmPZJhOZxxeuDntj
WVAZEwEATgQa1c49d8CpjBlvQlH4pTvkr4MumcbSqFgjEYyfZ7vjWftsa1WPwP6TKi59SseIBgmK
+pyzzU+IRkit6C3zZoBPO5V/iBtl0EkgqRyGlGdBy7b0PUVbtWOmtM1u1FQ+aPeUrK2dNrqh2pZO
/kCxjXMoMR/hmKz6UM3J96iReaDVff/Gcmxl6FXglCBf89COJpEiRH4Otx60fhkaHmVF+ZMPkGsg
Z+2GfNQ6JN+U+OpERK88enDpbogyQ51ZgTwvalyy5z9DDBhvPwx3QBqKRsvZCRkkFzqlMj4BFC3b
6cPtqgXIZ9L/Rgdks5cuNm4Zj/ytOAQcAwY64K4fb08xDsy84FfrinvooTUE78VxysT6KjrDvc9y
9Z6yviQsLoRY99edB0zVZCPFcKFpWJKoHxfrX1l2oZMK6CrY8ra0HnbXi1bYDFneUOarjKGosGHF
M0kbcU/Dw7Q3DYTmL5lMKX86xYDgFhx6avYvaob+idObLdMO40K2QREZkm3p87wqrCyxOzV7LRAU
0N7ce26q3vifC0+Avneocrf4vsM/1OLMgzyC0EFxILVz498lVHze2cf4NkWFxhsZj5/Kd1Ms7Xbk
qFBhRs0TtJjPyGLTN3vfXGfhQvj2RYqzxdDcB+sUkhfaJvSbkywLTf8bzj/lkkmt4ae9k7vbZkEr
Rh33O/8le0I1xPqkC7jYzmYy9pF9gDyBe9RvaKV9wLQIKbOMkoNZVDAq1ZRp/SlpcpWlhvww3MAM
j0YyWBEJ947A79tziAYuHtUUn5ia1pR2hGIj6U9GBRWHhOQd/jahN8GHeBpldWoOLlNC5zOsrJii
BfoS0BS6mZq+qqsLOOg4psWFwXO/RDQCPwwaLaWW/68PybiyPRc0op7iDaWgvbXyA8HKD38iZ1Jz
hwVA0DiqHn7IipcWyZcXRDUtJYP95nMR8KWx5+/HwLhiEcTZz7uA7Ds9ZtceGRsWNbpuio3MlWdi
Krsn6JJmfqsUWhp9AexgP6kMmePj69GYngIUlS46vAlau8wAlItqxN86X6ouOvA4o30Ecft1WpQc
72Ua3kwnk7H2ZiGypbDq4zdOZVzn1CvrM/0gvtb6CSuAGjyLnuZew431F22cunaaiWPxVzCr4rGe
tTW4LahC6U9TalL1g1fxCeN5CoJjjRJ9FdD+jqKMMXQmzgnczB+8d/tXSjo47971n826V5acK1zW
EP8TZJBfFXHwO7UuzSQKYCXgfeqcXW9sPLgtHiTSiFumQVBWJQzZftM20ILycm85Fj8AZFx+PTkb
I/dpzj8SHyg2Cz2u8lN5b9mBJ03FVII4DzZGBk7EVrhH7zbnhCGoFnxfXAztIBKtEa3BNe29Y24X
HJkZyBhDLtJLTIzDN8NbzoN8LBGxd4n2oWwNplP1gQ4t/Vdczzu609jP2uzeyphRB//j9Z7ZHSKg
lhk3NnRulV/qLRhaq1EZ/RyAnLU+8h1XOJgt6lg0wWH+fslhKwg6CN3Mf8lz6CXoithL/JBtF+am
+ENmI8/xVYg4H11Hgm6h5hQ04zJyi87U2bNJwZzEHwRiJknQECp4wZcm0hOdnaaw58tTkR2LyImc
Wvfpp7aHoo7ah2wFnr9BinYcX3G4KhjuaAa9mHemDOlwEtA5InLtMo5aG39rJeE0MI1l70Q0qyMF
NuerQh1eLPOlS3c0GFXX0tUyVdGueK9ImAzYR5JZ6QlbMbgsU1+Oh/0jfJYWxPyAZH8twrPMFn3E
p5kr01eHkTEV0NScgCaUTKdKtwYAlroPJ700xPJ0XgLv5oWKfnjkk4d4LHiIMrIXxIecL8Au4kzT
9npc8nGMkqerilJQc5ypPpwx2ocaoJBxJoIq38VSE2+3QmA/HwnWRWBfMhpu4j084kl6uTyNIeKG
zgcAXYNbOKem+i8TvdT1Ak2zuJks4BE4V6+dM4RIaRpzlIfwJ36MbiS4AhPaf2UCC3gcZQz5vEHG
Gvm3YKlGTLKpIZbaZwr+Gcyihe8yLMVU0CCUmwoxFPEt3oqmjiL/nrs/ZLy62jQwFJVKaOT7FHkj
57a5P+ioiFCeDU22h+hSBjpVCgqwQK3eY2Q9W/+8DFDqgmdhvBMcd3+X56UIZVfS6us2k85Clkz/
+EO8h/uYKm2t+3EF8GzZUOoPYeJk0h/CTWxPsHpE+fj05zzJwWNcomMp252xFhdRNI+WC4PB87f1
UFiyWZplWBcqAN2FPyd2ObkmiuR5eMPRKU84LMrokiI8Q7GvK/MyMkRdPrWRoudXgdjcJs2rmOrS
n7pZW2xmj2MlWPxULM3rzibknPG7WeL69xNykSLqdpGmUhMRwqnplBUaZO2f0c4wDUeGhAbYnL+T
UbkNTDaSRN2LTs8iiPoL/VGH9+arY/LBcj2L93+Cs3cOypi8tsk7eAvTWgUHmx8l0ITv6Mi0k8eW
nnVqvmqDHdCkjfPhIcrAeqQ6fjTsKiRhkFKNunBIBSrHtZjUEFlW6zmBBrqR8fZNNbKDo4CucU7S
1kWZsYDhq7xvIiOrrri6erxSIr7T1HPABJRdu3wUnSJ4sViOpzvfxYu93+NxvaLjNpzLJlWU0EOC
2Xn4qsV8I0ihvpjPphFZvBlzNFToeBJRH45R2YD9/yyoLBk4ButQLZzDnWKFUjW6Bw5QqM/C4qbC
n//2kYcRuu0qTuq3U1GRPhozZqAzHuAHmxpUZHgC4SbMRsuNpj+1j9RtmRuBKF3sCSuiGRMI4Djt
+sm9ZnLhpk/41Z5ov4XMr8egEsDuOd2E80zsvx/nUR6fIt6/cC9UWVmbnljjJc/DKU8JrCZ4gha7
0R7zUOBBaZe/tv7B3ZfaW07Cl7v4zE/1es5cDxHh2kqi0+uSKoYCeXLkQjL4ZxowOe+d37Thi7zE
OHb38iR5N2PAsLXwe9kLfHTTUGWBlMBtLuOVXk5tMJzvJaaZ7ze3qRY1E8I0MGDVpYQiuUAvEo71
2VhowFKo8XC/hCthfca3uZdj1x9hX0VQCR9OP8zqQWtkQR1sAG3J34EKl4Cq03N+s2UU4LoILImt
aqqliqKtMXaHYMsZ++lOTcrCYvD5ljE1kWloDG66yQ/hnaxJhB2QrQy+MRlLZqmDV8LUv+uLCH2h
vNeBBRvVUvGdtEmA4yKWQxJmaIjkrbr1pC/T4dIxd50iIhDELT2PK+1ab9ArRL9Mc8eQ5rxIdSPI
+fIRAtkQoX2z6YWDr56e6ac3La6AeyTxemaGs3DyRpUIzjTOk+n3z1kcf2J2dWFM9nWoJRp2A0xQ
N8LPPOWehX6/EodUu0PgD27Gug+CttXsYFwNIdT3YVBFTsWcVVcn+Xpzz6CTyIeWLSATgXUVWfLW
l1w0HyFNUG8MRAAyW07N4Vt3o+Qu5XQ0j2YM6gYH/Zq4zVWWuP2juErhhFGVw+D6/X8mm2fiFwQS
LGseEdZlruym9GVX/I7Xgs2Rc56vAghHF+tCDxepWuXtW7tswNB/CVTzvb4XoNBoPHzZi4qD2GSr
imWCp5VV6t4oNbxBj9p4BK8BvzCVmNlWGGqUW8K5KvWwIVSMreHs0dP3UsTl2m1D+Ds82AcOyik3
zwfHo/W43guz2hMQ8aENTaTYzvHHRVRAxq7+yzeAmg/JhKUHYyDxuioVvd6lNFp+9F/HZuTBqxUY
5DdEsZMPD09NlW61raz6POaP1I9G7EpCdw0wBudOQA28XdO4evXrdQvGB/1qBEf8LY9l+eMOObLg
4+ZIJ6vkQCWnbjB3epczOQ/WUnRq7g14j6MN0ZkkfbVoOCpwCfKLTQo6EGDK1icbXogX9C6Iifil
b5YpOKU6UQiRDUbyPGAp5lMzA58ghUFNAbJZbmOrXxZe79tltcsG+WCWZhXFU927KYxbMaq+ZbUx
ClLrMaAQN2QDsupoqUsZjc0pGMfNHXlHIF3xex459YFtQN3GJ3HAttxgXGKXnVM15/NqlsFkWJLd
2fIMNqa9rnMOPvA3wGFQF72hq9wPIXqZzTxAvCTPS50zUlCZm63W+X9FhBlSnFMAw/BYWBLXUV9x
NEQFZx9iSKaT+dswFvnm70awwyBkz3orYK5qXJX37VdHQbKY2uW+yXl00ULbicid3DojvZAAeia9
1eljfV1DKNRCRvsxveAB5myHReeqwnPpLNo4KrpPROirVsWtROiT/fPjuGUAhrTon/Pg5jGGZ5yu
rFw2yZNb+ZO1Zx6wUQVaRRRcEjqSvIYwBKNLgMOyVzKCNRX8LtvIYntuTa8SPEwhfKfgXeMhipD4
YKs4h4qT+NLugW/PTC+aV9npbNdEgUkGLe3oRryLJN8Zot7TM7TqMZaMnH8Rr6d4ul+mV67qroEV
jc4riO0nmynILT3JXD/qirtikKs8EZyVziOlYeqnotTHhaUfd0a7/IDZQkPEsYpZfXvJHG8EzRwk
dHXUqpDEg6rYMmibC1XdsAz5GjYQjkqQQMXDLEV71h/h0QT+XDvX5uLxxaSIpU3Lzc0l0JAACej6
v3IALnDxYPFJnUY2Bj3yZ5ycaRUpQr7j/Z3Az8QQ4cV7915zRNYjBwaWDya7y3ZKildlZV3ZMgLb
Z2YKNnRmRtygR6K01HT4lZr3nMujagFFDx7dNIxDZtfm1cMc8Vw3g2yhgYGNWEH9P7FJsyrwfJfh
wNSh9CubNhIelsBTSq69SQ5ix5yuYw7IQufi9a6yB9uY8Z/NND8XbJs1VQXoq5B6yDnUPP75i4dl
WzNEEOgCTXsT4DdecCC7CxNwOmwRCPd8fMHUJSrntTTV+Kj2EfEniaYcuIiNQeQ/sJa0yVlrSyxi
YoIb0l0lP5L7FLitpWC8mZiSsPf/H2SF3Q3ASoKH3lBUhiOyeyXO61QJrTRKFJjEyLQP15u1U2Cf
2NcAom7/gfQXSUQppFSMfMtxvzuaFkgrttBo/+PNgxaBkDF4rc9i6/+Nzdc1KjHmPmZN41NxlHL2
/MMHlsox0cG/PmbJrSYAaRrlfHBfoIk9UsXEYhngQU9j4j51MSiP7Ul1A+4c/DY1Q25nGnbvt+IG
vkhKsFobFDHKb9tMzpG5Y1ptYoY6Zd9VrYvJj0eE2fTS7C+OBYfgOC4GAswwWrEkIKP0rFVXT4Vz
/eMC+Y/ysSAsHjra3DIJOE7qg+A+atqnG0saxu+bu9Rnvbf7pIF37W+CXyekyX4C90YTRRU32rW+
ev2UH2HZwKUWWx9unIWUjBpwY0FJkF71LsnS4ZItn4R2NddPpDVbl6ioUo/uPkwyHq1WcqX/XDwv
wPrHiLyp7dFTGbKGvYDbN3k0BK7/lH7/VOFmAUCYrbhR35x37mZs+TJtgIv6GRWVxPvHrum7q7/z
O//AQcBxOzC4rJ2XYrUvlfzZgeGQ6PwEyRwM4IBMybSFtAsw7A8/1VHyKI0kd1ebtM3snKawDZb4
3qnaePMZqGrvGWETjk3wOoBuNrtGEjjlXsRGLhY4fIb2ycQb1rPUwI5S3rEclcXCsgdFPy4wET5h
9at0kU7ZvKuZmhbd4B+CMbllBLtvnSwuyJJYVr+PcB1FcrqUZa+SMPWm/Y8+0YZZeC3/s3WvZ4dW
acOT0/AYTdXnqb0q5tM0FcZuCPDH1bpIAg1CuM0HSO1fOBkuYz7gD789XeDHo2B3N6WCPDP9V2jh
Akz64tDDDbhRqJBeTFnS5iAs/qPJFml+KkAY+66kO6FioDx3RedVUcswe8DFobIP9LcgPe80f4HN
ZFevGrX/T40okF4bOR/gQMHd4i3znxPM86uVLPGewz9cxkgnCkERK2nYk2PxwGx3/0NP6/vqhnlq
0ZslRNZNmT+2ghQG9fmPHq9msOAaHQ0IjOSEgob/rKQjNtNgFUJmHBzRvuQ25A/GuZ9aYqhz4/7p
GtieBRYOQEiRkRmDmJvzN4wFjBhsdT3txa0ZER1wlrKv7hJgurjLlqGoUza+nb31S2c4I9508MVc
Rlh6muIvInPrnf7oyoMOmRiFuReugKXsQ0veeW8IpRbG6sCTViUV0gljEyD/qmm15Ircn91yGCws
4y+Xo6EYqgrUv3F+d6XOEGOTLptWG1qrCVbspqZ+/ZzRh34cxlO6MFeoMD0CrSGQk0a/pAHfj9Fb
3Z3JFAR3cm2D4sKoUfVC5+PevrtmNk+uu1qucaS4PF8D6VDF4voyyg2/8FgnDRd6q0lPe9OLfWZC
jyCpPvWKqi83bGi8ZsvPi//ZIVQ9DPiuq9bsCxo+4B93hlAEtsguOpVE3mLsKJ4UnybGxNJqZG+a
nEzCuJhYHpJUN1cbFVl3lo+14GFwDyqEnRXozwsU57lrFoJjqUNo1ZIq0ppoP6hdMcOgLasck02u
1XNkH4YWM7emd6MU/q3KhuhW5phIhrDt3vH7fSJuTyECiL7I3C42yPUAqsxcmcvDA3IIZ1k+uYpv
qb7xKJkW19ps6nrq7klBHCPLDrm/aQAs2K5G+j39VJRmLaq9rpZzLjbiVXhZX9ncoG3/qNRBzw4F
ksdHUwMy7+jJ7DIks8N9I/m/0wsyWdxF34UWZWn9RnSWoV/zMyCmb+2u1bir4S5B23T09OiblJGu
z3Xg86tGP8ngklaxckh0C4M7uYEIBQ+4jqKAiAkY48fA891jPrAyA+WfVoekFcea/ylCjWO7lrIx
rzlFy2MDZSnyUHWi7rrQyOfhzSoIzZz0Og2wlAsGoQ4W6WQk7+49idFeZAjUEbVV+0WIOuYtMd0u
KMYynnggsgEKUALI2seetzfmG3cXgGK+LfIR3g3+l/k/d1fOSNOqpNNipKgL0Kayjk6o4eyOZl3H
2cC4rz8mBiKK6xTV1EMznqDKeDBAYYshUFxoDIcZn3k87x1QpFef6FnbyDePOICnFASPBiFggwlH
t3777+SBOGPgZc7ljq+lXYoq2OBxE6qYIneZo7hH4RXM/LXS2/BV7tEC6CjJ/fGJm29mWTXNSrqi
A6mNWpLyytzNA1e/GxI3exnch1Ysa285oZ9vD7IQlWLJskTBWwLB7LSpCr92Yd7wQ54lV91Ggvaw
+wQd3AwUr4PChoW0Y9IPc/yYUd0iCYvqjAIdLavugGowLFDQUl7r+H8vkNCtFNGQZKYW6GhYUCur
0XyJCLzj2YAP5L21trIXuWt083bG2bz8PwHVsXhXwOrZVwkkeql1zRr+w5FI8X8yF1q5QpgcEzPD
PfXd2ixZsPAxldG4UUMnOL47KFr7kOa7c8tpLwLZuY+eCCt1bY5xq/B9JUvU7fazdIGPO9rYhJqT
fFEn9ciMYn/FpyF/5ERbw6NhBqiOeAGny/vxDkMliKCCfz3qkNM/BC1wtbxYxWU2L+kHzmF2VQyI
d0yyZbWIfU+PZkE9ShvAiLtRjV+peAr7dRuN1UEM0x5hAAY5t1jBSFssP1zttL4X12tl33pATdBu
LAoInqbeEDHn0HeROuCW0OTp5Qh2Z04fjNN+fWmlSQ0kRuO+svTv0xJe75SWaXZQdThG5ffr1TIl
Oy5odaN4OjHhsluNsZafzZ6MTTJkcnKDylFDEleOnE+L0uUWgF2ulnBMbYtU67jPsAQms2H+Bw2M
6KZIes55xNC0I4ovLd+3xp3nl4pFII0pvaOsEh3QfwygGHIbKxX/6BDbOr70omktm5b3sM5RztQi
3VZBPA7bgCI6raMCDenW5f5N1q+wlZhtG7KX0SMDngrmotKG/Ew9FEthcWWWuZSb/7PnJE25u6k3
0JXgBd/r1RtGVK1rB+PqZJAVbJVP/yZphQhoIQyIugkyOI56JpHka0XBj4wsNQoARx2NVfOi+G1F
5/go6XbBTWfPiqPmqbFJhlQS7/wePNfFXMzhzXk9tZH1KrRCkgi4xWKNc1H89us+SgNOZxlWKxh1
zhRQvUzP/qzLbNK5Shgdo0f9cDQQGSpAoweR7LqG4lNfCqSq/i3CLjz6mTVYfw+smFx4TXSkT+WU
q2AMNYHfsSh5riOUxZ/mpoXAOoQxuUtbvn3kKCWLAhCfnfC8402PnWipgG/kLhXWCgJ5GeXX1NVG
SYE8u3Vzp0iidL1ekYHIe4BpmtSpvedkb8u+sJWOhkda7pUkwu+FjQuUbdsoZ9ZFEAR1Q1Y+IrSC
PTOFzapmRLiE/Em5qlSs4dAQtz2FGwuovGbCPKWExWM81BJy2pHNwVirjzKNYDbeRtbahBajgnOi
Mbll+7eQTdnBoKdJJnk7q/IDBOEaWZTw1C7pjmETqRRYvQu/YNgwpHZWJ7+MOarIyy8YrO9Ko/gn
6Odd70fW9YkwU55WBoN1GL/Dk7VT/62t9T1ZL3bzff3f4n8RJfECr4j9a0pGT7YXzQln5rpptw8f
QLN1NibVgtOm264A3VdS7foZnl8JN2ivcCvh+aVcirN5L/rBQb0uHp1HoWh+J7rob62IzdbvzqGh
C9B2cY8KhaibV2SnDyLPMDJzj480GDNP2Xppf5X1pUj5XIm8klQBuwGt9RdnWOTF0D/Wt6pHsJC+
vesllqD+snOBXy8YoI15dOZB4EYWU2oLAfXgAuomAZabzZNSjvR63za9GHRIys33MtFmdyVDvyto
BaYyOrhNsFBZpXyJ09mg9c5H9EztQLVW/LfXqs8NS4fnT/olvp3pv5xm/O4n5AD4r7ZGrzi6bYCF
o0fruxZFs2SwmJ7boyrOzYujafYAMWp67aJpbdqPYo+RNYs5KZwmKfSIfevHnKVFsvCDo44CQnK9
W11SkOIaj+iqZoX3R5YbYf07qWIEf9mXYbZcNuUnTD8PKkrGqgUxJPmR6P1+MuDX/GRvvTdsbeoy
Mpm5UIyowjpDvPyXANWzI4aA/M8Kk9lHEDs7jRLUUAtqIj5bKWqasGrLPMDi2+xC/NfKgIKji6p2
SFcgXbbyvMDcvPbhytAD3DFSMWd5qy352I4+QKY7CReuB1EqSKdkPUVqLkkBUZ8+H8CHonoRGiIk
IrMZTLqUTUinuDoDiQDylPx2nEUgggL68D1sKHSJWYbmv6pNfJAX90LqDD+iCzyPo07fQ4JLpWaq
goT6JvQp3MIuyEMecox7XzVreT9khYOFIpdu1VtEM2T77RZhRDSTJg+1i9k2hX9UY3Zx0Fp7MnU7
5ChzwL951LNSqZMEXEnsxDeXOqObyiBDdVF3IQbwIEPUAGt4mJ3SxbVbPWMrhZ6sifa2rjUAoNmc
36GBaeW2TrxLNtcts6ycshNpE8RnNNqMlLEbEouzcs2i1YqPROqwdkCcM0oo8/X4I1VW/QOAcLp5
IbdHHE6H2JJ9V0fpu5RCPfqf7RimnxiQ98Ib8U2aADLy435b7b1FsxLF49ihCpyiYydjIxVvHmoX
hR8qy9pCou2HegUaQHcVE07vJ3miV51AEXpoar4dPDmHMKmvdrMJ1x5YzWCf0VdHeCZ8jvTrXVoh
bBOVG0UZfKt5fNanP4OMsbn2S8+2yszNk8w0IMZtpKqJ78b1DPoTPbETxqCexEI3FKIjfuV9Asnl
uFPLUAPx7yna5qdy/wwrmDtjRwjjGMBD18FZtM+NIgUNZNghV8iFoQGgH9psyRj/sVNh8hbEm0Vq
YM0esNxKnbjXTExl2rzfUQfXjTJA/Gv0G5MPl5DSmeI/9d7/zdBlsJ59F13pHXhItNVaxHkzk4LK
shvb8XUXanaUYBhaMa1LBaqqfqdMwBkUeFwIENtSNtc7DWJmuGg/nl3sdSQLFPN1lp5f1IUGCgP+
eUc8Ci4Ve/9MmP2ZaKy2L8MS4hnGbvvJNFywOP5bh/TR1lyq+3kNs7ExDJt6fix/1V/Gbs3dK3TS
V4DDdi1V6ZoVa1WV+9LDdv/PprKwTVJxg6n41O4GF73+zRAh7Oum65KYcD05Mn/a1KklK2pEJ+fk
i0Q2bFl8tDF4oMXqhKtpNvPgJoB5sEfVeLIqwQrlkxYXK+F+aPYHhblZGNk8kLOkEHOeyAXkzXi1
/TtuPNAVq140AH4+5r+bsyrIx8C8YQGwl/ORYvvWhoQ1wGTrzyPbbRl/TheRW18Z6jzHejD+ClOq
/WyGbgadP8en9ODovX93tyH17EToEcIlNSp6DhODK1RLQ6gLKaudASZS9qD+i9hy8GzGc8xoRNOO
8LE5U/9/HQWP1wFBgnr9bxO4UuYESlDIiJZyV+7T1ne49Qj5bhrPqx01WOzWWwcLorKSl9v45qgt
zBu7vXBXRxF0kphcdTSPLGDWwpYq5Ta0nRy4IklwmEzpne8KG+OyKubz96J7/rkDi4YLS3VcWwLC
RKxy44rIAu30M5gFywX+FyCfn+zj6NlCijnUUm4o87IsLBWFyhArDd+2+CJvIpJ+NCaECXvf5jHL
sJJK9Gm/mlvvGMKPfNBennO66josr9BK5/+5pgfrqfTAUAuk+MpGwLTp5e3Exwarv+IESRjHvjhj
PK6lPxger0WmpEsg7JKB2U7Hd38bdvdTDGc1gRgh1sT9ac5j7wiuShSdFMWVdc+yBy6bN4Ne0Txj
XO/pfooz+qpcCW1+KLKwtRCJnE5WbBk64L0W6tzSuPIHBNTdUwlbcEAzGq7Og6idz5qkMmzcEYOC
gvRpvV4prhUiwfqobBRqo9M6AJKmnhgYcdOPuJqPGro0PG9rlTvZPqBGu33WK9MPyIOyZg6J8N4Z
d1ydTNvgFTO9szXlMkLz1u0FnkVBcEEBb+R7u2rFyE8pvshJL/dpLfelJVHt0vFr4x4ngQd4R9vZ
3I8Q+xUo8CDXmAkPNby5aW1hNLo+cf0MgMSNxfDn5FRGJ82ZO//ucLRKoQazHpvqzhdmqcX7yofw
8iXlWODfGusnqlgzU6sCTBonct+zUObhlB0e4abbnRqWL1j9ww14BMJSYFYzAI9jzvWlnRdh8yvo
khXvLYz5Lkd/v0ZMB+OLQrycQlxRpMKwSFJatKvD0oNDq0Met8ZN5QwHT7BwjjbBE+3q4H1D44Ns
+PikF5DjVUUPlxxN/wC+xEPM6VjwuFxjRNUw96MtttsIK5H7TcbiagsgZKaQpwRdDlH1nah59VZi
zrebHcBJUuQId+t4d3/QB8Q8DX/MfKnECCG+KBJrM3IRAHWIeeDOJY0zcpLURhpkhysjS+X1yAQl
8Efh/f/203SLv1j+HxHfx5lBNHiuNgWmbKt5HDGbj1B4cs4rFr/EQ6XzRGcvLwhqQAY4OkDOD97b
R55wNamb6TrFsJ/gKhIxw/UXdCOKLgcmf+vO8kPLtMraO5YoZc4yTTgKYqYu+5trEpfnpsPSL3+Q
1ohflbBdhZ6e2AYuTnqNH1myueG3CGagAzaYFZDP7sOJNJen0lJm5qvci2fuZRnrovO2cYqxAmvn
bQbfAi8/ooafO0EVMsp9ZG3Nfee5cYA2s8olAZvX/fSAA6/vpmwcYLNQGuoPKy2tlAEoxFYnxih/
FEfU/OoeScMapNKEqG2Jz/Iq1qHIm1SoS7ytVUnhnR+dPP+8RalIC8ZzCVA7x08VNJTOijPneMsy
tfElbEdqhmkVS0MPSz7jQeZvpB0nh2p3mmYHDmuzFDH6d8rz7gVTq4XRURKtIWXTCaNu1tddBkal
syWoZz5yyhTDyY+iwOt/qxazYIzr6Z1SIpbwy8yrsn/swgG1FmSxVxk3lf2k5wP4OQxnp4wMRRBN
PDPhlUuHkvB4qywPXu+PktHnkhzzmGK9EyJ8oTDhyzFVmHUEbuNVowWQ3z0G99Sa1C3GyWgjl5/V
joh6o7lQlQTPh/kXat9TnRJfvj9U3zqcDw7mWio6jkIvhLvWMn1qVVrXVvtw6MNHNVKN+/xGFsSl
dJKR0RILe+ijQct34kBYBkYMzolHK5vynpqN9Rl/3Ud3iTVakKeeCudu82bqe2hlpy54cCiN0HDS
O/8qLrgFwklSOAML29mxR3mqDkvCoD47MrMZ++Ewzpzzyh1LJGZG9ixNzmVOaR2T/sZMe0w5CEru
pPWkUdsbvhbHdqIq2vvLmXbfTsxhaCIjepMUU+Wzhf+MKAcA1cFltHnbQUQOUuUTrlVkLP6/9war
wR19am8ePbRGtC2MQQXYej8DyIq1UhgbzcTqWfgjk7tJglZoX/dYt+luU1TgqI/I7L/sQfTpCDPo
8Fx+1emOJxvbSfj+KHHJSnXhjxQ3GL4l7B2mI+uDCmsCqnJXZnfh1vZAHaBp03JXIlrfmlqFoLMS
BI39O5BGhSyGNCoXzBXym77QgM/90CiZekQpTa0xLIohaTuVlpwNB2wOIZFPWw6ZNnJqj9xkljC4
aZuKRn5YvKHP/lZQqb/QBQdi01M3lpEbVOxhX2bWfyiOTn1Lqb0pbbb2LjB9m3cumty/erEQ7yJ3
euqCsuNmdwUfVRZL7klImvoc6A19sQhBdxoxijOORvcbbUtBHVbFhVjkbMIRWVk9Rih58bLtQIsD
aTW+YMqKIX0DICU+llKlW4x12w5g8YBVfGmWLHtSMvPEq6q1ifXEa77bIH0RF1Tk+CAgrWU48pFF
EovfgMA2iO1cuDbQ2tsfxhDEJtD3rb7p//Ebs6T7pOXeliy802X4G1lFqtOdtp+cJE7XREo6TQr/
g2mKbFIltx36kmO59mvlhxvnQdE5V7NkP2o5SCwzPrsvJ9smd5P5KeZLciSRaDYP4yhPCzC+evKx
HEUv33YAO87W9Ol8r8OJMHlj9d/4OoSA/BZgndDjvswm1SGoDXmhck3LOVQlgk91GMmY/dtrrFT8
PFizmIO40b+JBf+qAZVB0bDoFfbjGrwx7LP/8054u1J08F8DDJAQdqAOxtYCqoaKFAI3vfj+F3Vw
wa3HZjfgfJdEV8Z1ikU7sf1B5nEGiJ3CBxWRn9N5k2UDmRRDd1m5L4YpDo3lfsjoob8YSlRi0x1n
63IFCfbUvBPy8U64/JylYlSOaoL7RG/D93vZboZCQcCs6HtdLy3BT4OHPeY9cwP0TvMC7fvqGuW1
Y5B511ZbOEqOu0xTrxGVm5STgBMoM7JRBgnIYsVEHpWGokhyBQ8S3lCWXXb60C2B9r7/nwX8LsOs
TyYCaHbKVz4cqEglQk6Shzzdq+8Q26gB0JC21lMWMOQmodn5dj3KlW2heBKEE84qw5DHfd+4l6Jd
TDhVXjta+TTUtM3iGVeti5EzHk7h8pQi4e3QG+2r+6QwkWLMYYHA2Zj05AjIEPiWYF+j6BxmOReO
3Mhl/VmcG0vKayjLRBXAoqnD13yC/+cbYmYFXm8HC8/Ib9EKircOyXcGDnnlDxFUBbroNS+72JhG
SxtSLQcfXJULQdtl9LqG2Yz0cnzHjmLGuVK3W18YAOFJEc6XY05wip9stexGtqV8+ytOrgCmomDl
XjJH8Ew/ajFH9OByBwowAnNknhL6Ec3oPnxFOUfZ55QGnv1XmbmQdAHLSrho5VEcdmcVH1vaTi3c
T04dSbAD0p4cxQYx6HQHUDsFo9BOnKAqXTwf6C3D6wwtLgzftVIsOHFrJTZS6q3ueFg7YVqORZqe
dYZRPZqmEHVop2jvq+k9SRzXlLIV6jDbffsrjRlpYsFRUDW00wS4BUI98C8vDEDLYc6MMPYNe5qN
m5Urr3xhzbnhThFindzPdEMUj6lNofbf30k9n+cuNHd/VARcURRl14MN18UAcfYgL5hHCqXUhh6n
Q0r2HGDCYt7WchZCbG2OInNMEKzbbT1xnI6e34XSxrgiGd31z9wXBj6d15qLYjEWwvHqBDqrzDdj
LTRLlbhp0lQIVcRS6BsN5vNuSwwhRiqltXYwFyd9wlREsct2eGt202ssgjOQ+0ngtGJpEvur52Ob
akaFNloL9um6tJ4tXv8Ub5DFQCa2FEsJLaG3YURVd9ydrGOsOprTx6IoeICjvHJMh5DLk1oJ9e3V
Ajki65ITa9qDzeGrX+d7lnAZnO6A1AWI8Q3rIuvU3HnSQ8DEvXSM42MCTHejVhBQqAuUyJ6hRvL1
T3EFYkiDg5AAW/GmX2c53bKdTWKNoHy3+dBx+9IlPpD4tKhSxcDjiN3BYewbYFiLWVR1JEIwzRAH
rjwk7x5Mp4wdMv3c/SnAhRVcSl1nAGx/iNKBZGABxutPNDpkBg3cfoDnWov3Rsj3PJJqh+oj4QVv
az5IAMGsnwgHkBEYJrA3ozKFULDn0X5tJvotb8FAJOBXjoVz7d1FkUe79SEZWsi7e2fEMwkpr3AS
C9sLAkXuK5wnUyqjyXtQmWN7Jgoy4yVU0dIwIqAja3h7Oj+MLutFSXDh6WBr74uEFeeY3JHHQNmc
OXpwfBeqlx8WYHE/iZK/NzvkfWnVVIG5lh8XyYQkHDYwsWbok1FFbZ8XUMuo8NnKWQ1LnCWxjGk4
atpMmxIEr7vmPX8wLNMh1FlGMX1fdKBwwQoeZIMzceMSY0VmhmByivQaIyAxkW8G6OCNLim7LRjG
0ifdC+k8XXfBaNeVv22Fe2Djf7ocyfXBfGl7C0E5yz7mZ7M7pMkDZ+XAUeoUS1q7V1a+EC+9mBnA
Jsg2KRgwMzGMIqya2RZseO08bncy4vkGlUbGE7X6zMylSvB0ta6U+dCcQsj260NpHL5TG6WO/Oic
Nzui8DsGFBz3/GoR8KMkmLpssX5aR5d2cNBsVpJz2JLgimQ9AR6xu9b4sG+g4hYO1yK5TaqDQbap
xo7fyqydmPHgi+806rFnp+7kp8/pQYt/0wnlrNs1Zx4/hV0Xaiosgv8eKX9yLN3CXp8AHD5adYlu
bNpgVKobmUJhacyqj/HtTMedFo8XixbbPf5ods/7k8VQuA28E30gXPiwS04i8rEceNRqvxTAFXrQ
HkbDB8aTWEcuALlJfhJSdqZOHPzfJI1Kqdp5PGqbgG2T+UdCyY4RpmbQiCH6phzitR7K6yjZUxS6
dY7GRWcfN9kX2y9IFRtyqg6b/G8Su/kwN6nycrIFzHU8hcB0OX2Ef2x0oWTHbrWnoWqf44JoYKhI
glxjfItKsaVh/e41wKhs2PEP+AUUdU6K6vqHht/nARNM3LdwoYg5KlowBFz+c6/ftAB6jCUbkxCc
KzCKh9pwBDbqITNmIOa/QmdiANWBkgEkl2FESmOZZiwOWseLZC68Gs4j5esYEr5r4u9PAWRbfgpw
o+hR3dyZuCyfIcBwogBYTtChaRm3NL44Tg2L1t+Ai4/F35q3DTJvJNTWsypIr5QRIfte+UsCieRe
27kt4v9B/VlT1FdYkqt62fxIzlXzLmOHRi+gRVXnAUVPQ5yy5nUhV2kqEyd3lxgFrfgC8cKqOoiX
976ZUycziRREu7tNRxwV6OPWOHWk6Fw7SGy6TUIdtldIhwZjLaf5PG+tZpSlf0KwEItAMGJ6vj/l
AlwOv3yCP0VJXMeWvXqj7vZR99xnR7P91pRJdm4M1so2CUqEsj9aIheTfu3el5XwUiNufV4E2bP7
zobSNN8AqIMruNKcCFqlvH+bLiITKOGfKh4A1bwOuZHixBDHtgQXu4Lm5l16fsJfQmXkOoB05e2T
+a4jTOM6WjzshY1KJpoeXN1sv9EC0U/T5TnOivzM9DYeMyVfG7ztawsTzinLFWv32MBR8KM/f/vv
qLPmsByRfxTor8c5CqMPQDr3/YxBLQsa3I1/pOIfPEmvv4pl9uII19DzSsmyDinegYGMSb2aqm1/
L0C0EoZllMcQIkbzFCbfs3T2erM3X4D0CNBRYyXo5M0g5Hmmqr6F7G0H1DRtvtyMUFg711SPF66N
ea7ynnWlxDvUP4QO8v8cGQCDyC9tOmTW9FRcdkXH9u/JQsvGviMsPY9oO0hCrcW3zIITiX6VbsW+
dolYgdBibQ/K5kKQP8Q/KHKLUiVPlI0MrbubkV51ixLo7LiNZtrTj+QQVx3hHPHXqOKp7dt8HHHu
ZjIlbV4YtYvN1shAeLf7iBYiTe1sLuuk3PlwqDJbH4dRQ0Ikjbh8KmG8GYBuduAJGArBHUwhzYjv
CAqH5NyVS24AbeqK6kMThNbW9bjtn4yQdeKpdZaMpOdRj+nIiVQaOOtm3TNf7EBfAgw23xAoCDf9
j7OgG62pyFdTJTc0L51ZW2jukbMDfAHxYrK9eiZNUaNWC16pBxNwoPQGS77swkEZ+LssRyRTQtwL
sCddxyEq8r9L+rxezospje+tdwuTLJ1cVIkhUu5ummJqW7FEwEOSOt9u8kHlb1LRibeK8aLlDM5s
wYwZsMDLtdV2ted/JQl8BxbqKGtGfZu9B+8RD5DSYkRayAMLCCo9AkBJOZ/+fjf89HzcUwEzZm6D
F8Rh431v6g+IQxZGUiBifdbcb4Pzrume0kswJ+SJGnbtp9+DRfGNkrEgXuScrzrAKWd+l1e2nhpT
jU+oUEVqM8f8vXBruoe89czZcvD9qGcaowtxQxw7WIfX+CYhlDg4wqfSxk5W51npIKLzOyd/2HOi
DlDwSrTaEFZUQZC/DZN6z34QUgszCi9eBJOCSkuCFjyJjGExTPnTSt+/IWjvGrKVkjR7KNZzThuI
jdNkSYSYSqjs9tvCGbpQXCzzJzGHa8rxeE/Tmmtkj0oHzbzykhBGmernVhuy1Dj/1t1gIQdGULr1
MHm7eRAsbx8Te2jCJ6UI6Po9DxToYXlvTUyL/r01v5WfM3fTvs3Y4p8s9t9+krxM/+P9txpCYS+a
EF7cB2rAPrPl/XKvXbDQ+U/2C4/jLpS85Qh+K79NzLW1UUS0TFc7YjrP1FZvR+5lgSNc69Q7Cyji
zRFezu2yxly85jE5RZmVVYpy/BDTu53kBxG/DYhdvBht8EvWmjZgersGcvTr6hDHq4htYGF7RBp/
Y3GxZInIAXpvhWJ8qRiNO12Bp/w+2CzWdokAXqSwxmKH37nhy/OvmOqXVBG3UuhCJau10WLFwjMQ
WQs2H1+SUPBX4l1OYU7iyQx0h6H6k6N2E3xCYUV44LRabixjfP5jCatoKOFfUCFiqKN27QeNBdsW
w6DZx/lPZiIDjfbJN19g1xI5BcpUq3zEXPZOo3jJ+FdW5Ie2oK0qoJX6ks9LI8PUUh2H9Twfwrbq
HR1onYVraOwy7NurX4rr0hT5d1cvWfSVy4WVRd9UJzggIj0y9ob7DwSFdTrJC8FlaLJ5j4XYVvOp
Nb1Noq5bnHY8izDppJ3gwgR7XFzh4puO2GRvIN8Ca29X9jtWeRa96pdVHaUiMKAvKRgnMCOuYwx+
Ksuea0FIcmGU9wy7a4TZulS/qFXbSXQU3EvSqeQihELPwLNUIe26JsYG7hvrDDeUe45n9V9iKY2w
1rJRbJgJspvIBYVGxSEXI3y7+qn9faTigRHoVC0z0eafvqmoOV72ft+KQJxdI59ogpwY+j4uS60Z
vBnQ6N9AMPMXenRPR3ktWaOTgesODan+YD7wggVQ1HxwEhuJVMwuTaDTYNFCwzSJCCkWo6qzHQLV
w0OeNfxMu6p7M6mYI4yIBEzaGf31wbXpegS8mtptJnB7Beaqn7pRzQIMKLmw9iPfj2T3DdnYNm4w
3qR1XAsNqyb4+zZdw1zn6rlxzCIkasDUYCX6ivulDOWz9vWqSnvlurWxoo1HbbWYrjTMFk2INtCj
+PO1MV/9rfYgzglBoiOZBqSCxc4Nwk1Xzx2o2ITqkr8SxeY9HEkAtsfCGBiTxX1UAgX2QqOOMyWQ
eacUSiWlk66sCE5Uedc+gGMl4N/68oLaH9AaoThKwVfz/YCNVuhduwlc39gFFO8FLyJvGfBoxC8D
4BWK+qXlwREk3zchr/rjYInS391G4ciPCAY1TZoG/mx737zzWU1URWnhlo3+TYuOEVkIB28xo5ot
x+NTQdGW1VJCkJ2bFkS++gNgGsjF5oCgfehBS3KWL7HX0ezzSxWQrgc1XW/6e+sfduP17ivl2ZG2
fDY2FJrZWIuAvymsNuzG07Ohp9/WTLG7H8JrcwtBhr4lA8tnE2IjcvotPkSj9ZsbXf6xVXTbo9ey
BC4KWYhPszMe21MEg+HsyWNAsaCN3nqhLePp2zYhi9LrIUKLImRbVTkr1XSI9a8G/pWyjHoYzLPO
IyXZRfzqlc4g+AoCMqQUXYdxAe2mY9qzj21Rkuj//EBRLud46doEiT0BY5Sjcx0c6DDEfJm7l/Dh
cImZlkFeVzr9VHYgDoN0FVZFbPYzyGIiGFd1FdEYMLSos9+6vrdz+jBS8C/HrnnNtGPqJbeQpl+k
fLs/ilb5yl2d2rrafxcZBnUo+GlJGYO0cliNcaqlBmWpqQY6HS4BF3tcjEGVf532cneDS24S7gj/
uVwu8DY0B+8ujybUFDZSbPeqBlAJwyFHTujZe315t3WrxWRMGaIOKHsbdQyb2x8WXiVLMDoMJb+1
YTHlsQjTXqfG9uUw+StYRlbmxOBZKq3Yr/rdFFnB1yrVtXblmiy4jI5DQm9x9D2odNn0z9v/fJa8
zJB7qzmMoFFlJk3utDaXNu6qeUDt81CHAC1I5Noo2hehXg+OxwBY5S5r+r1xQva8oWprWJgfn787
qjHczoaIuNRJDl5y+JFQeC1Z8spSHsmU5N16KbKBWrYP1LKmA3TR5wdQ5bX+Bl5bcmjlFQm3bq/J
/mEYNDFMqqbhJjSRMdDCT1e+vrCiYBmfnYmai6m71N9oQigBRGdneuyzk98bFsW3vUES7RmmjIkG
+DrKi/NUdh+bymzPn12fAI9yoTHbhrhQ0zxnb94hvrwB0tgJyjzvSWhuY0P7f68jm9FPQadaUxKg
RYyede/pn5/MDip9W5RZRiFGIXG3br/sDEiCW3m4X3HS/eFVAuR7lBfpj2S0vmX9OLzT4e0ZvU9f
4XbgKHP9PR7dtY8QljO5i++YTMYrHr9hKrWP6LhiTA/WDaghRfIP6BgxYzm1WFCqHEAGfkCdc0Wc
6zwqlHHek0Ln3iDLQ+NGU5tLKj2c9kM1DOenv3H1sVCO6rSybblgT/emhsrSgE8+H69Z1lWGjIsi
qEz2Wr+o1+6OExMjh/sTPvaevShvmFgmaFKDnOYS9TaD4pavPMTNMZZ+Zmvvf1DopJmJKJH79b+2
j+V1a8UFDvEvicwuzgq1Wp7Kcz92/y9Zww+jSOLx2VdWu8cFqUWZh95A4eIcPG3orAlL5H1Eev5l
RhY9GBC2onkHw7eCFDdjMVQj05f0YgVG7i8KzwBeznH2dfUiT20BFHWb7HABJ0b6cHtlVpeR++pI
iEFBWc+MdiKi5+Ju1ovomysxhdpNK0QS44HPiCsK5zm8JGmoKd7quf3ptl/w855QH0x3fLkWEbMa
3l80gOa2kpZ9iG+4aFRgpyJrqfU7hhR2Dx6XZZYfB2BUN/ckPq/46Xya+rNTRm1Rm2X07f03rkBo
KMEusWwYyE1kGbCzZOaEMDESBaRHCdXyYcNmKvThRfAqYPWrG3JMzqFEqrHmIpbTlqW0r6qTUcdu
UZJFLqN5/PZbReV7KbGVe+n1AQl+GA8fcOgEwyDthJcPJXx0OQz+qpZBn0eJOlQDUDfuz5mSANyT
oJy7LUINtDaYtyDjbm+5Je1/GHM6HlTrlagNBg8hYriOxMW1HtS7W+MeDQCU/HxblD+wowb8kW2U
fhhAq0tk+GJX82vs+4hjjg+o941rf30qWeS632CNXbHGIGUVfu81dtfPP2pdFqJX8B3uzT8ncvGD
0l25WxoUQ2dyLwTZRST82pn8snRxHzvhyQGg+0ArxwhZ6cerMdRv2p20U6+Wd6pMaQbTTQXsJ8OC
6JQlkBI4Qegx78hncMdnCCmy7E0WlNMN9K0yiO+PZyFmKMdeziNETcKoZ08sDCCVoLKM5ojbrd8O
TMSfX3lpsDuOLTI32fzbn60hqbbMRxLRQScGYmvLY8XiP+owmGSkj88ZhfZcEkih2hGMStg7lVTb
0tcuiJYDiNfDNWPJBL157oErOr3gBQN5GNuq3zv0S7+YJhoGouHNAC/+/1IjYgWNfmEm7GuU21LT
uBa91TgaM2VS5iemz0Cjuxb2acK3hRkZWgw4EwALF0jXY2F0xI9CbpxUumLe3LIAD8l9k4Ax2qPM
7BAy2xoLAdEDJc0obW5NVSz1UQeq8Td34sjLqVuigwkI0avZBWlXT4me70g3Tg2YT/wzwA2aaB5E
RThY2HhGbQ38Z3hKqjwQ8RdewOt9wGiQqU1RaO8rgXPbSNOxyHWY8Cm5TffIK0yRYzWO3EwximxB
j4zMfHC69GOAo+rwKMOIhf242wkYkOVn8+xtA3hGTFPqwGsi/kzjnnNMXDVjbCykAX05lilD/w1i
fXGUVwO7IQptCEp5jVFFuNlr9W7p9hXqIZ5Kio1rNKNqOZpOvWjhUoodvhYFMqY489J8wdC7O6Wg
MX9hvj+UFznkW5X2seSbYQcValNfdHhN31PmXFZCwBSPTkOPzPH8mhmYo38Gub/ZY/Ps7b/03H8Z
eDAO3F+CXQ/cxvSw45Jb6dTI3BYUEM5/+tdB3xtShXV+Aqn78ddNdxK7+RguTwZhtlSUHK5zBKtd
sZNnPS3xsfwb0VRyuU/yCu5Ddj6JxvGQD61DrMTDOnnObpZQKTR7Qu6WxogF+fiXFPEvjNo04knA
D3JYR+UXtYXuLRLs0iwDkaFY42nDxRhOmC8vnE55RmmtBebyzS51wSBhCv65HC6CbxrxV/UkVi+M
uoTAG+5gF0xaS4uEgDS4BISKfkihee1nW5wd558Bj5MerMFcen75Pc52sh4dV3z6tWZEhyKxQEVd
RhOIObYQXEm8me+JYuI0aKjrzdSIE0auU27bbR++cvOfdhYvbyEGGTd5SYBp7ApqFZQre/ari2VE
7/adbhpWLuzHbsuZWHX9qVi9Ombs7/uGx0b7RD1LN4h+zTJClJA/JalmK/BY6jO1540bSIav3ng0
eBU3ZehN2H7DO6eXF2RwBeRC5Q3Otm0KP846wKuB8ylW8j+ZIc9TlPQ2hfI2CuCzJOipd8MJT/lO
j4V91R/Xcia4ltwZ5oHAObGR6UWOZNeYSHJy1mtsyXq5LwddwECWrOSFJ6ferpxw6EemlNOWA+Jx
jwrPPV58qcJV4oRe6xreiqm41Ya/iZCYy5ChIefhmNzCa5rkSvZenxzpDc4o7Gb9ffGY07QW5fIL
DGg1DY4iJ7XY8JlfjQMOtAGaLKFTpqUazNEYgx4iHfmKvtmkDQbVe2pALVDtDHY6Hgnw/ccEt+eV
k5fPzvi2Lo+d7nq0Em1s3KmqJvVHabeOFVatHU5sfHLjjrivQXBuFVppg2Y9csUyZvqE8lqX0Ba0
4JxOvMk87ODHL30SDoEQiulj8IkCtmFGrv4UB8NSjjBKAwLOcF5Ut57NahhXJNZKOOcy0pXganFT
oZ8/Qoo5Ess/lGvFAyxtd65UPzsuMQITtm4lpH1g13bEkPeCvL7MXAdhkKdBZwxNLcI5Q+9VcMqv
iuBGYL3/vGy5K4bdMeFmFOwdGXOdEizHyT0ejoZMAOTkuwpKSNxVI4W5qZ5w9L42z5agnF0uQznY
jUH8lIyHI5B/8LemkWoqO0SwOSBoqi+z1ThC+6XHyIMhMWV1fYHfRF8Q14DlnkDc9JGzug725YGQ
NqLKc/+l9NVV7U6WqE1N7VU9ib80uaB12IqckWMfM7NzJuIUs/rvc4P6uedDNT1VQ7pvRAaMfFUm
JCfwMy6h8O/Hn5v4tj5eFJTZeK34jHJ5erRcSpnBh9EOSiHGpy8GqEfp0cgGVkrRvOANmegalK+/
imi9iJYsx1sjqoolKDOCe+uB8dIIV/GWnMiZYNiAEkQaBqYlgMfeAFDaP8z+GYlGhXRwkXbpZKtc
gZ1Xo1+yfS9v+Bb8SZk431bIdAxP7LjYTuNH4XZEokC3EogycUcS523GGdYutzqR1IPEaHLmERDX
c28bWyDn0CAQs003s6ZgVt9ZKGAzpozdj6macgjizU8Pz55rXHQLGfCq8gsdGqIyOhzXaWclaWgs
qro1U+tna9mLpTfVAEICR6ITromoa+HqR3DI6sCkdzTRY/REXVErSCYxdcZ/vluNPZtV1dnF8YQG
uibaMNVs6nA51E9jdaaOMdwtqSj8roUg09aTWqblxyBUyeauSjs3mKGL4j/dq44UX5XgVHTwMq+M
texo92VA7Aj4cpQRcdUcLNR9uI5bGq9XwlxYd+zKasHkcJ+8fV3Yvvd77Ym7riq5x2RGyLgnPl+X
xpqk770WZnFvXem3ltC1as4DaD4vDo8obNP1fxR6YmX6qMcePNh1/kWUzmPXY1Lvoj/7dOUtzt13
xm++KNyk874UIT6BQqlA91QB5O7GY2P+KRvIRMKos/s/0+5zW7Kmza1THkOzlfiznuxZvaWhliMN
vBzFEL1EK2kUiHyx9ebaX/qsP0kQBVKYOM59WR1M8/O2zuJWR4+U/WcUJWvfwkK/kUUMliDruqtP
LPFfsGxdT0YCEF0lUdbDEH2yyQ5qCdD7uQsXmRVVSRAyWqRH61xfPOqkS4/wIeeFYXear9ArdGTF
TRD9t2kVXbCt+Bd9zghwSzIqDwtcVRnujnywMlDm/g6fr7cGm9feHtkjpaa7cxO2REFxu1wbWgn4
M7Be3PS/qH0KguLAZOlZ5r4PFL+Cy25Hem3emlr6s1GuFf6AFsxNhCfA+wVoGlnhPIAtcqClO2o3
yrhD8s/vJkyuQvgbDUWWjArLxPrc6+pBsdHk4QLZ2FEMs+YTcq1m6SnZpSvbQuiHTrYjVhepblJT
ibfUVis8uqWl/GpGmEB6mxCDbV+El60dOM38pO95/gbCAGj5I9q6NKXUKjMFDc667x5WUpgalNcO
eLJKIW4vJFmcYKVsvlAZiiH0Ou4c3JVJ+bPbV7nhfy6tWNjQN/di4dj6P4VO1i1XEfdqKIbkSc25
X9MTA+tQzvVJ8Q1WvDppc1Ovr8kiD/X6Q++LeuCuDMOI+qJ7lWExMWhhxctipVtW4yXUs8HYyMM3
fjwRS+eke0QCh8sqZ3W9HEfYcGlB9gl7xdqqgav8fF943iuWJgcTlhFMHWlcpz4Hp1UlKdcqD69C
I24mdFa1aRMZNzqDcTPKpi4Z/sx3ZGjtrT7mJxDb7ZaFDCoOWK/Cs8q5CqrnZUrjAGtcOVzUFkbQ
ysJaxpaamkTNYYZg8loLyf+DljngIe41B2dzDJ8b+KvrWEI50uSpENSbxSCW7VQJo9j5dPYDtvT9
infR0WthmS05JDss6/i6Cu3RALCjbGCQcDVrNQ+89vVsoHj3ABsR3CiBNabf8KcFLRSAGU7EJM8j
DP2W6NPkWMPc7qR5fZmvl725Uhp5jFCdFh1YGpeX8h4uf9Z9xeErLTqLxRsdgpFDolo7Ds9qxTdL
CxKOZL0OoN2DkjRZl5Q22lO9SkKPlgaWE8cYpEv32nOgmBlyHjfxcsiRrrm+KZSJIBcx4DZpgeQT
lnYJ4cKMkgltwxiqyCSmBLea6BS0D/vZMKGLS1aGzu/NJQol3hHt5Al/w6JlXixa7Hg7MZPq9N9E
CXsZt6klySYtAWu8tfXj8lCjDSEv7advZhTm6ZfAic6xQUtQkFwHlBpNTXOWg5m5yTwG/GsdvUSW
TLwZ3ziH+iAb8zo+kDFVAM9w5LlHJhvXdmiXBjbj36bE3Vys0ZuvQg48GU/WPOtfJS9G4/WBKHBO
xdEAzbkb28PmoWpKDeFgdrffc0h6JwWoy2eLw7SfWnQIODwUboItQWmCIPNeuHPAMwM2+FQnJLjo
TerCJl79w43tpbEXons4Q+kau+lbajxMti99h1stQLiyzxOmhAknFhqMyiCg0raDJBlx1MMRSeeW
ModZD7jZNc2NTNb0+53Ziwm1ZTmpYt5uLEtlPgYJB2byMNotLZxivR3FhdORuXP3L3xvAPoK+TKO
LkWqniyDIlCleeabwdWm3kkNPjYPXkpzPnwcuQarCKBVg9Ow+nvRNCcEPNhx0X7NB04kq+REcKBk
X1/IWFTvFx5R7TPODrZT+n8Q8H/A0bPWxymX3GRDuV6lVWAb4r0m/z52LfU7OruBHDJ204TXyjPE
FTivNGadSWQPUu01Rcv0otFGWdmTIRHLXDyy80hkvS8mgQqo0tjBTeew8vzATjIa2avwcEk0sceW
+Teblu1Ny5O6D1Z5xCQeZ42mqx8sbWlNM5tSPwVYjWnbJ/HK4Misjgs0696jgmVOsx0yQZrskfzr
wLgL99fbPpEWhf9Hhi22Vfnq3tOtcqHctr0u9wettGYrxKi8BGXNhBGMK05g/Mrd+kjFJ4sBliv2
ZXQ+XULOBnZN6kyeXDXO404JSXo9z9V1pkmyWS3+w0pt9IhAvM3LT1G8pr8IE6EzxoF0s98YD4AW
l48I9GIWOHXcUsFPcbJ+a3MKwunj1h091KnYSv2NGguFYK3CMKGYbEXwuOEmE4PbqEg0KTgRt6Wg
lV/raO5AVszh0yzvB9TPqE4tycWn9v2asQcED9FYB4Y+rjCZWDpvweWLCi/gKwcMmoUFzqD+Bqbw
rfhlYgrXM0C+RH6HO4vnaDJakgj7SR2oFtCF0pnw6e7DazdpGH2bnJGfEcz90U6ZVUdLCEHBSbdU
lSKnFW0gRW3zmLjGHGinkW5auAZKo54cN+GUVOhjbvL4xGXchkAJQcsv5CJmJjiDKNnCP+Mj4ccw
RQgA/aI8y7nT0LWiZyuAzH5xCQjDeHk+r/UKyGy7C9E+gc92CKMjVTd3Xo6nujqrcJqa90qawNxm
BuJXwWUGsS6J2vIAd5OFDquprktVO0EEa1RwUYdkQZ58QUcgXeT7nla+iuMd9N749VdinpK34dJf
rQc2yJiZHp549pgYOnLEjd5VY4zJAMTFLMrbz/GWiFpDaMxcu4rLsOGvq/jTPgZoNr4aR5WFHDyI
4JR7hYkMtzhr/l9N32nhkPAfj0BWfCh2crAjxnrik7c89Dh69ivfqzd3J7DowkVIQnE1wdIYbWU7
pPGf2a8+QHbezsuXPJmi7ExqW0wcRYuBOOWirh6C+5+hlCwUYdCpdS/9CpwKvKZnzylEFcIMd39K
2zuppCVVOGLa8XEF7xSKM8188SK6ycZfK7FtojxjAl7NASh0/qMTz1QPIn8bibXQF8Wk0bYUnD1m
VPRdE/Sr3KunMcwy9DF4esQ7p6gXZUg8KmDSgONa0ZYH1aYl1YWTUy/L3jtIlSbtO508x+0DDkxc
YDd9D4s4VcWKUKjKE92T9YPekgWvdZh8Ni5flH4P061nogkEfWFmOTrEgx+WMZ9UPIcXnH2ITNi0
n6sgeU/FgcbmCjkBD89nzKtI5bMdHpK21iU2TU2ApvRcMmlMutbRGTvNsC6IUL2E9pAUEnRzrCG8
RXroUtu/TXyeVuahOS3tfhobhojgCnWn7GHG4X8eDV5pLyjQvv6pIEY/IoDEzXqvue04Y8V+PBJ9
cc97I3KuTxfLrWB2mWQXH2VFPNXCb2KWcJJNT/K4blAE7FeEtVqqWLdFjm+8ynr6gpAqmJ88YyF2
RpOTCnU87sj9i9Rd1N9Vy5Hki8nPjuH9V+hjDHMaJhOtrFMU7CyeBoh024Ish6ZrbaKAuHMBqFpx
rTc1OnO90alKp27Qijqdt0Y0y9FbqX1dLOPWMAcil9ToOXKfoHPqRBNRw+0+L/PKfPTPYgHGnkEI
nHTZXis3suXjZ9gOVfG6NNUaEXNcTRmCWWUEJDNcEG0oTLRXh5PLLL+rCPOU+LKb61/gsgSgJ0HG
9H2aBLbeerozEsKCo7so6G4Qb850ro3wmjWDFmz0zOQNR8AZraIn2P3eRFeXMJsrsvrAX/CO4W59
iIBYa4+KhBWvavD1haDTGrvFYhuAKFv8thCIxDNN1goEfQcVwgqU1bw1piaFEAUDux+8b5cnrpEV
SA5h41wF3M1YPOek1T6pqno9WZQpdW539fRL++4qk5d56iJIQOzWXfnkQyr/aXH9+GmKLZVDhApH
V6Li0bdjW4SP5eXCE6F3dQn07GhcdcejgFsRZcj0b87bEz2XY67nkD5EKZQ0SlD10WLLc98jx2qL
widRaJFBvl6YQoLdmuEd+puIybkuB6AP/AnqtPxxIyZJkwkINkj8/RP4in6/eyLBpHpeE/fR0uWu
ACfA/JnVxl7lUMsXz2+Li4YIdSLGfpcumAg3QwsKWmJ/XlfVYDCX+GNIhZMugejyz9K5dtd0HvN1
1Biem2aJ3iLuzaZWZGhQ3/TOA8D+snGGcJhWbAdJyKMQ9dgwOYg23HMKa5V9uM2Uu/0bLhEb+w83
OUSra+2qQNqr3rMfCF7cgZSC2ZjUc9qCSUhb5/pDsXbiTerccoGopdhhG3myZagMECktPL2/eaMt
hXijeV3ZzSuwyFScliLnz+wQSC0s4fq7E7Z+pnvogZyk2X92dNT1GlRw5RalhEatfWcr+FlkvNGf
zyVRbBOsYb0Q/nD07Xqfv1uqyBAmaSyjNsIjKg+lggl1kxJKHtAzLvV6aGQkhP4Xvu3BglNM4h9b
vvqzFuFVquK5axhO7j7TYbO2tbUJ51Uft10H3ll4NYz5IRUYYMp7HsZFtlDlVDICkUZckMmS0zZB
FcIog39jIO6jn4zqZGqIxZpFA1E8dHl8LJ1pDaP/3sLxsU4c8026SqQLNEh+wGRl56T2p+bhXTV7
XpctanMqx7FefzSPnw0lZgNjnQ3FtcM8OMBLLeQ01YcTMjZ74zX2WF05n+crwUo3tmR+5of1qsnF
E40ojPhg2vi+IC7hiNyCQO+Fm+dIq9ohe7aYaRqzEx7S8A0bmWosndTfJTqzpt0ehJ01l/VY2KpB
WZwI0aqWqc4wpiUWGHCeWv5EklLvfxFiJL1vuKTnduOXdqBHRWAwuau7C5iFgwuxmMgCGwPy0tfq
6tZ0axZCtOtt6VnaQS7Ra8IH1sFdcCHDGvoayKN1ZrkgEsUCEjsumxw6FY16bieGO37Nlzn6x+4x
Cu63c1dYIslipXWwGINc2oTK3au/P912EMamlEu3enRIRffR8g6Gze7s9z6Rm6W8gCTNbCO0iEI5
y/0svk4VavxOD9ZGrMTlr8ug5FcfLis4OErR84fcbJC8Qlq9OqUCbjl7/vvChQYmtNchACWdclMU
mOeyjewOjKdTENxs+sa2Osmd9GCAKmQYvHZW+PLzYNtq8/qS88q9nY/bRjwygL5RIQmPVnvGOoYl
lqNH8lVBUouvylngiPtgNhs/otW7VArnR2Ty2QRlQ0gUq8Kqsm4zt/2rveXOp+Xuh3or3lY/ISj/
Vtu8zrPDhOZPJODopvAD665pWUuFPqeTWPuG5vxzpyXsrhYMfgdBbBjg4tlde1/jn7+kQmJRt34u
bvyWMgtpFvxhgzx0u05MeNQNx2h+9oyWzKc4Aag04fV7ERVzUMY4GnMZL3dErUIDpgEEYlTfL4QP
0GS+KUa8w4WibUNoPpJH32GzRyUeZ7PTejNfnvThQoqFy6NsmMlPunkg9keh/CJt0xb8VlUXWpxK
7EYR25Ex+7apGVqBeqVxbQXbXvljE+vnHoT+f+mDsyZsp3uLWMb4o6NeyvmVNPWQWA3oSW5prBEj
6dQSKwMhSQ1Pn4KNOJcW3/yM9Meqfu+PveQ5Xz4CE+/yRTvBFBmnJxSHJWx0ww8v8kByMRlILXPe
BxRBsPZ85rS0+3QDU0RGG1+djyHvw/3mxGZwvQ4lJkkNIFYEWLqNNMwT3Lqy9YBS4NwSBTOUsAuw
Ly6Iac1RRnePY/j7LbmKs6U/bdBM00lHORJZBQrZoojZeuRpe0MoL60Rc3ngM2Yyt96qTRPZ3xfN
TftpCs1FVHXS+o7JOWN8ScDsVsXbZz3Wdgr6x5VS2UofccpOg1IfVTIdytNqNW+S31o3jwGQNB+N
2afsZblfDb722zBipDak34/2tzLZF1uc7tW4fScybU+QU+HEilki6HBK36+oh/O6C9AmMnGyPhpE
xUkOkB5yGNhUmflT4QyqCEnwGGcOgUxho2N/Yxtmi6tiq92Dk1CCCDLV7uETrZP1SRc2SpnuQ5aS
mK2IqHmkBw01xMKHuCnobxJ5lVouWqb3U5R1K5tXip0Kr85snUxtT5PSCyzG2DwcWcuHILAVBtJS
/ZCrEcZmlbEtNoi0UkT+PibSxgs8N4Gxnr90u2IK8kxSnGFM5MzR63lSVyZ+QqWwQOPa7ZwmhNYR
P3gU9jZnURkIoMJCshJF+4jiX67TbQMTvu4qHs3rpdDdcRaKAxsM01v6BtKnz+Bb4GWXIhslkoIg
2x5vtIQyUBQNlDHQCjdX6vPXziJdCUpk9cdwnkT83nlLxaQwgWFE6eRk6EbfR6rPurOhfp8FGkLz
oOt54MyPqPkCZwFuPs9L6KwwZQvLfgeMa1nJmZsIRmsFfj6kGV75BatigRps6JrxrVmywtwADpxJ
fAb8hWOVg+Luf+bKrqRgdijSuW0tCqUOnIKoVEDa0fVNrD1L8ONJdl9xZmBZc1ECYSS6MRESkdJR
gKbXLRi1CUSdoZQaSYYjW0uAAoywOtEt3wvLq60OMkvaPBC7fzjF8aJ/jN+0v74vEVfISWCxLjl0
jYPL8v4gAybJY+i6K1ARH7mJcGnBdvEbADgeIE78Q2B7T53vZK3oNr40nQpec9iT+XNFMiRLDuOc
M7ZseCXfPH0aRKB6losHskM8SFP44KuM7v0rdPCm5IvxF0yQZeK8pTe0ZQ5zzngDPBHB4WmnMbcI
oKwgkC2tlV+5bfsW8to55Mp1u9yB0yLSvRJeYvS9CBa/hgyC1352aNqmMrYQ/cijsDXMj/pFro8H
Zr7pT5h0Ct3toJicBEXGZlN6dR+hoClwfMNqBPgC5UQkRTOSZOAnQOtfYFoMzI/6crcXNjUvcyTW
PTSeNvAVbWDtWlAS9VlaSUoMdEE0NogMrE/qMkNIMZ5FOUCiU+w+ePMbpAuCq1n5D2o+5WbnESHt
AHNXm/TDyXgks74zBgXGNvJZRQSeZUC9b1MV8FmSRRWR5YK6UzYRBiUvVdfvnXcoHff9tJXc9rFT
LL0ZBhmCorJt8vTW+B7VJTtBB9lEE47kjq6dsA91GRbAmm+HZYDuMruIId2hKXXdMwbzbyaRbzaE
BalKWcGH3K7fk5PsU44oTj/fUFQhUpWPQzbrtgsCqrXMOWn7wE/2UYwMEdHkjtbwFFmIpgU6apXa
dVC9uk0Lo5n7R+s46m7WmHWEgCebhIl47EfCLiRWjm3PEOE6roxHmHFhPOHuDP1DJCPdOPkbKyIM
EsJma/mpcdFvMwdrhRzNqzXKELob8pefhlp7z0qhpIP7GJJdaBXgQwagBPHM2CjIfWtpDy7KRRI1
UwXHf4JBaJpC89ad2nTF+vsoC2bgo5uK0n0qcCB5Uret2UG25qXukcCasPIGNbyeegCZuUqm9he/
rE9db75M1eMnv6IMq1B0+O+Je8cqAk7V0zstDaZZ09kDKsVa3v7/r0CtHzCR9xmQSYZz9p95Y0CB
xzLhkc2zBp48JM2R/zniHcbIu7cDA+sbRKJHU/BoSPRoGbAqZ27eJ1qmGVgP0BnZNqsApdJRz4Dg
Mah324cGzIhzrtkCXOsXmUk0NAN5mc46kGZz6Iug14AFLLWrYf09ksXh4hm+S17Bk8xFXnytamdC
yXY3saXs3MIJze0mMVRAPIFP8Y5Et9dH8hM5Kz4rbHV4YZHSpmtIPU1do0013X3yJnL4uq5VaF+B
5nII/L55ODfEjuJjTdPysfXIDYb6MmXZUswm4DMvsw5d3ujxLokyoG17XRdIC+5C4wCboOQenrIC
+uNBNohf7nFbE4ODAIUWH4kIN4AGWeHYPtpmuACUrYKtnfr5ZnNGWML1DWhGrcgvuvjkGhQQl6Iu
gj5073qsKrsoyYmrK2BTVqkYsxc+YEJRfC7pebffCuRW/OH1QQjew7xXqu0wf0iyjxL212fGgZGV
RQD+5DBkLBPlsb1Cp3PS24o2ymkU48HyDArPICimW+VQI8r1cFrCuLrTu36nO8D3yAgvw0VmwFp2
BBaR8VtPaf9UQHQfZNFfwt3wAGhnLDTR0Hew20Q1VqXAzb5hRHw5+m9Zd/UrprmY7w4mGnzZxCpU
By8WhyYUIrn422Y2bwJzusaMqsa26lczQvN3atINzDIL7dO/zMD489YZWRHox/t2hItvupBEc95U
c9Om/EbWKaxPEOgMqSzam+Iz0/HybccG5+Wuev1J92aFP3LYCUeZoWKe8WsJQVwRciO+ulXZ4hLB
61LB6qU0WohkoDIDDJkZYVBTCvL7aR7GB6oMLF8H/aaPHB1L2jplsEvUYAPHllpd4w1A2mRo1hRS
JZP1qKm7glSnjXvIvpRcH2RGj4oAvCmrsH7k1slzxavaQ/kOW7eSJgezRv0rSQZ7y3N7FxvWrVKU
6p7mvINqxx1SA9993X7aupRWpUgBqVlyOTcp2gHM4OX/lWpQ7cdOUzkMeiWY3kEN+xckwUdITzhW
zsiHgjmID7inNWWWwZ+8C8bRQ0Xfehdcr047Ba4t8ag+viA8AZaMtNAa09eNzgEz+vkPcWg4JxBI
EOihD8NK5pQoSC11ToJBi/6V7odGMANjyV1gz2uaAK3khOxZSpGYPoHt9w0JD2JluqYwYcCD7SWB
ZSulgpR1vj+05Eszy26MZAMG2CwbqJ2bOfrmDaIWkqietUGLb2oyd4sNcVj1TkCHAYSvPWL6aUWR
9e+SuAVATax2TlmS/NONhz+pU9NyYdM8KF5YPOP5J1kb60mCUcneTMERA4e8E6chnkoUb9Rcg3Zf
TM5ov5DhRLmVaywQ6MVuRuWgkzeHBBcsP6KJEdzGgo61faEvWRYxiwmxzpI69pZqlqX0mzlm3sph
IZ0CJ4gwDedQg+u2rjSVpYcpiz7h+BOSI4+ZPIXbFRBkPpeTd1tNSmbHtogwcc6hoqs8MajWXW8r
gqkuG0hGwuV46A+CX42OBejzHzzc5ML7NjsxrIgzeuCi6/KDMibyeE2T9fhtlS8uHbdK6356yLJV
92m9Q9Eo/sgVnT1VvqU3bTZNe8pCOQnf1XmXiLl4MGS2G9xiGDtFswG3AEjgHIHwiSQW5M/KxsyE
k7h5ruitikbryomq9plX0eqXkH4MJKREa5gV3X3JN72c9w8rTceAjTAxDwtUpEQEL8jUh8Y2JlG4
qjcXY+NgR2Ongz3gPAKJ2N5CJ+N5hAf+9hj/fpTodZavG1m3trvy5bScWHmcbwdhytUxmhlsiise
0jpbp8q9dve2Upu+YLh0y8HuahECCQ0ZB7oPIgHMTl3CjIDdDCSWUEwlAXXYPfsi/P5ccNsWi+BW
ldJI0bKBSuFzhtntlrxPC2kAcLPWXdwLv1r61bf97BRBhwgbmwIAsuN0BEUSIsaBkBHZ41OKB4iD
0ef5mbpxcPKh5Y5ikb7BrBI5HSJBK4CODV5ylfDUMzrLHALJrfy/ZmoSQlB44jrXUA9g3EwSd/uz
lXS5L5W+WJA3n5BGmpt0esqeDNC2iIcRDNMjEoWeGo7W9HeCsido5BQqvcN6vMpyDjNiWplCovgc
z9u9JbqRCI+609sqf1lepXZJjor65LRONBqWmD1A6f0zV6lNRfIgqBrLtJl/xHfM55zm4WbkcTg4
DWbZjxW08HF0OT43A3TpiFV6byQ2dyekuDXtd/r78e4ov6IFjKSMlZS+aZPRAXAKCoQyssVFH0Q9
WMnT7jSjm3I4B1DNhxzqMlGP/Vaw2aGArua1Yvj169q+eBPgSg8kV8Y4ZaorWsoT2++i6ZJzIj4z
izPcm1ysqx2Dh7KUchKCU1h/D1YSXdKd7htJu4ddKIIOlqE6NunRmU8bK3R5sm9KWVvXbUAjGuAl
PKty6LSb8+6bXURyTpit63y8tQ9rgkK57i1Y01SEhsY+5/06UPvzX0Ytiqyz5FAGTwuHjkiGQ+5I
5P3pWbFnijwWwuEEtBi5+JBxOfufnDP3C8AdqYu9Qvna+CwX3EC1rC6DME2itKQn4mJDLTei6OK+
R9AJAiMbZRuYmdC6af7XWTEGI4f1mKlA9E6hIwCoJDIHhp+yrL4vWy+6S/uCJ1zdBj/E8auWT/lN
OeafPTHDxUJn8HodIw8SJ3Y/JxvpUae/KqJBxtmB6tk8Qd5KEcOjabpZFYmpc+mG1TiK6TDj52gp
rHh9vksbCp1joXNpjfmfCRHAiq+XwT3t4w08ArUXrsRIQZN0u82+SGgYrzY2th+QNjwBG8AGEaqs
7iZZmuvmTM2Ik6mvEkol5yYJ8PpB1wz29s2DwbjLwzpB7bRmnbiNw6SbaQ/i3tDw58Z7DvxBodJ2
K3T5gj0gH8uWjcEZkCG8DC5EJ7V+/Rs497wdULVmfwTpAyZFVk2YHMLQ+Dwx5wg6baB1AHIakMw6
2Y0xjpL9ZLoyxdhuWkl0lVD0KxRIw/op1VauvzQBJjQalz+D1Dgczd6wPDe2XUEhZKhxaeVq0+jF
EPbu6tSLaIDIhD+Mi5/IyCTy0aigui9VxKdhDREtvZMq4sYsB0RIjn0txeXhIDTDt3DAsUjtFi/Z
i4QXH2jQLcyoKt/VNtXhvpdo9pOvwRkQw8kKLb42E8xZvxv/K2/gD7EZkvUBNgktAEjjyr5IkR5S
b7lXU//SA63oLZdpry2mcUgyirhP7s2Ai5y5a+MajmdNPCaynnIZ7DIWr/UgGxfAjrHdbZrzGRcE
M5vQkPpCpT4m7YU9DeFdh7151jI8FYVYFKOu4GFjam0WIkYztABmgFmKPsR08I8nttl5oR3659Ab
Asd6SbWP8F+Ql2C5/49d8cAqkUK0p0QNIi0KR8XAAtEu2mmDUCRcNaFED07EHaTmXklzyqcc020H
08wYiYSBDZB9gghFNzUCA7A3NlPJMALW3HRbxxf6/kJi+KGzL0adXVotZChPYe77LTHZ1o/wJ23x
QEUvbJFsxQdzx7afTIjvUUdy8qyjMRYXWzV0P0ToPamTT2QHaqLPJ0VIbA5Wok97ox3b0/aMFF2K
owdULv7dRlA+5cGG2IUezkyjX/e2g75dhz9vAYVHn4Nt24+GmY3pD7N7Ut/ApE42Q2ZWFXhN1yxM
Dwt0QExxi65lple/pTD9QgGy5RfjhIJw799wa6XY7zrVHxRGfOd0hU6V2k4f4EVnQNnuPqy5x7Yb
hhw7HZADzZEWiDxL7QNZ2TQMSlY9xzEDGEd6l2l623IIUMUgf5ST7AtOKwjzNeDgZ4AgqpgVQGzo
uUV5jJKlotsVEKxjTRo+SFIHQQAQNVBgA5d9rqqOrus+rhZWX2PcNSlj+leBfU+eULvxTlCI/g67
CAKr6ey/JYN4qJ/V1sjPI1a2Ci61z1s+iH6tRcxCdEEuQiOpfYOql2ynRjau1bw2+KgkgevtduuJ
J6xP2zJT+BS3TPbGIYvJRVHtpImQDOgyldOrb+UJvWNcU7NuaQFQaiVM3eHeYkV4epRstUTtGloF
o3/JYm5OWE8khUYLLm1YmBB9cfxGLqaMME0+l5EltDyhdBqv6SyuoN6Us57FE99P9uOiEpdzIkNf
qUkc1jgOAz4/ZPNuMOTGhy3AD7J4PTg9hD2uun+mnRTaxZYLUyD9Rv3tFXm3NC2SM2tcgaIqLMul
sBsm4dT2R4/ta4SoQMNV39fQWwEf4cs5yVJ5aLDcqWJ0kikSBAJJARjcsoRAyehryAdZ/9QvbQbh
p4wj67JMaNcl9OpRZ64CcoRPEKZY/PmAHg22YOjh3MR0d4QJ25VU4TmAcsDzi4ImHnOx8shajTsA
3a/hfp0/XUx0lz0cvrgTQmiPEjDY8u94gpn2PwyzAABZP7rShyFcjODwhmpHPgnsvL71Bh4al+XO
EXTkpllAdnrAAJgzWCaqRPbJB780xQrPkgkMcCn0X7LttXBQA5TS7hrrR5rmp4sOH5i86ID7ZwxH
ydh0ScDdkNUBIKhZeUzhY9BJxN6C8kCTW3G3+F2LFIn/uVsaxJOTjwiQjlYllyRfJT+zVa6Ira60
09oAkTtHwKgpTViMd/C5XJDrg4n4Gdzj+m4EEwej3QTXOcfDrQ2E5+ZeQ7Q4IHk4aG3COoxU8Gew
xJS3ccLrohUDjo1bLRO4Awf1MUJ2WVtUH7WfWe49OSR1kRirrrpdXiUJpBwkdmCAMujsjBiG8kUj
14eWae4novNyim7KlQzsLUtVEqeypf0bCibK+ClcYM33qoH230eQJGnQ7oQNJisXZHmYUuceA0Jr
iWESsUiNNdjq6KTpHBvjg1YSXQq6CpzTaJVSVrrYKkIkBYrFnDhjz3my9B5rZYfRU3PK0Xaw6D/5
5PCk/s+/6vJvudcwE41lEGeRDZ4nDUslHgsxu1JX1NPp5d0HTTDOuAxEadNoup3RTCJtPDdOXT3b
fT0lmd7H73CvPnYe9iMkVCU5dxpcZCT7SKPKDhKGQI2oX/EZP+0K91bEOLjeODMgRkM4m8X+1OlV
HfidmXny3mgS76y6TGtZfoIuSe/nlSIbfM8eRWRkzAIjS0sh60KbpdRL8kuyCt2XgeVwRzwqmw5q
UdmISjaJ2hXNjObg5u82uHqb+a2ZjU5psDvM+G8lj/AmORYirNrZ8NY1jc0H6Nz51BrRRoTj9jkV
UMJfuQzAqY20gruP1cqcfTOrp00lOXZeLgDtiM2oobiBtPm+/dpWlPx1/qjzZKDqgeD4AtyjOyaa
rvYZn7EnL8/DjUTFBeTnICZcwYNgMwiESBQmXXl+fLApeyBDcjZGThCQ+7vriIkKmVznScopUwZw
qXIGzHn+Tnd6xaZsnOSY18e6k9oa04MhXomF9zPJrzzUHZBfItDU2nWfv21qchbZVyoutuEI8woJ
plraGAxR+YMHfzBnbgPOx3fM9qSKK4zRX7XC5IGvvhVqvb4NUJhS8/gWKtPf5i2aYXSHmUVCHC6Z
7F/nU64mqi5dd5+KSvVfhFgD3IGNME0f7ldCecCfSsClJjuY1MrrD0MuPHocNHuXBBEM6XABR1XL
ZfclD0b7QEIZPnVMHfLSv6ZhfJiMGjHjtWfYTTXVoUcceGYmmCq4iCbo9h7RGLYiS9yP8CJaqY0M
YzjmwrIylueL0SKb34HOXQ9ctoT5VKMC0/H4cVY+lbz+Uf8xXUgAPpQnKsu+Y39hi23WP1Ga3iMi
mspZhyL8LjrSVlSAhrNA8YluTCVCc/NNTlapwQVxV7QrUrsVFWQ4+95YtQFE8lEZxcS2seFKboui
Az3zLBbLsnKIRPvDn0vT810npv7qSpWVg9VUaMouCio2fABtrMzj4OFRbny+c41y/UGtnDKLqGuM
8A2/t8W37xJZs0LDbD6GHT8h1xoWFrc8BWUvfaxG3O08J+QIM1aM1ofzxTe78q1ttPFgND97d6Oh
dHnsnbdDxWdrTw/KnxDwhciiGsDAJIAlplSIOC8TVIWHmvsZWyT+XUm/A0WJIsYMwVpsKx4FTIE9
v2vVYR9Z3JTYKtrASl2zt/KtbRMVgJPocp82t71+Qo86rHEcBvfzVbt8+wkRDcF4H3cHQBNZ5Lxp
IpLFvVkTujpRYkDQmbP9YTpBtPuBZtVogtSwDFljbSJR8KE9YIRXmb8OtdOSEt9whx9WjnYYdWpx
lQQ6S18+yLNOSO0siimXd2bLhPz7ut5rvMuBgJWrWo9TkSLElOJgVhmiykwTuFkXKh6oxSVTp0gr
VrNZ/YYfC3jow42DdKsIePXBfR/f53ZpngBcVOXrZ2MDMzXbtI9a/0czOIrrsKgiwqu1KJG9u+Yu
jRgKELZs62yWwTfFyDXFuaSw3GBtULS0+Fey+OQ8R12cTEbe9BTbSt/3fS/pbPlGP3XEkNndzXFb
rr8UtSp/CNjol3A7rDGn3N4L0QtAmef/4jivgeuTONZAKaxjfrxkx1RAwqsDhpqtdQHNi/R7NZPq
WlsXbMCn3RuTQ12as6U35mSj9frJX23tGp2zSGiZn9fzKGWQF7LCbJwC3mP1UaDqZgMG/Txxs4wd
FmUwWEDnb2YM0sw8W7WvYy1jwnn80PyB18VOTSHnPbiEXFI5POzKQu45mNMC6vE3jmAG0x/M3pzo
xhsCLEvuXNtjsy8ETND15pClZn7St71/FK9n7Ma5zJf9gj13TZg0+vajMcU0sX0wQ2wxVTw1FIax
lvtK79BKw+0sRourMOGnzedlusZfWsatjHqV1Z0lT+kJ793f7K67JBXI9kUhfC6ABBOXbz0koGhr
YMcARg/4UesYMj7EnXerC5WNoRoPfk8g7v6yzRgCDBISfqjg3ncQ8ZGtzSHeG21MiLkQMjaXMCEr
9xAjjzc/4mCpmM+uSz2XNztSOBXmDEVb7w315SKHImq5xaJAcRAwnsS4hcgpuvuSWx6ujJPNKitW
BBi88TVCqk5hOcKGE8/XOyZ3xbNgy5ZpAcHV8VVI+4zmhH64/YJ10mItiWHkbwY2n/Y11uX545zz
qBY8ylLqzxW2jvr4LohqFyYZmWbnVPBM17l+Z75Y/9SlxGCJPjksa0jah2ZBwgu1pPcgsefGmImC
B0TaaIEX++rBLoPCk0yednZ0+cVFt6MujG2ayhpUPlSv4bPJx0fuy0N2ekqb5o++fKoG5HMBxGi+
xGAJTM4C4xaK+7eZie18gflu88OtPlW6KyhOi6D7Sa16AaJJZ0xha7fk3puheRwuWa+TwCvmwkal
ofJVxupSAtjArEgoPKpvXuNAKIrJRmSTWIx0yLemtg18NRaK1s8JK/kne7JjX55NbAiHaAqQjP2S
u5k/ytJlHVxkuFB1riAbgEECF3ZrAImHB//5dm/QH5gKsUETYKbtEiizn7xLWEdyRKiZquqc23+s
uHWJwEd2qyxvNdUDnS9LdrpUhtC0Vquj2okZYzufUnvsMtsHmzx04y+TGxRg3D6t6b+Imdoih4c+
inQa3yJWk7A1kTtoBjOl0KZEW/IEqh50MmO7+Bf9bbgaFB88P6ekGsIPIBYNLu7qv0L6Fhkzzpba
D1rU0Q0F5os4QXSBvyFG2xqDh9nDSEiVUswJU+yB9rU9G++ugbPmO3IWKweJNlB7PvUAeo53fxhL
aTztToENNO7wv/KSj7POui5FV1YsVkre6KZrQI2Qt7eZ1vCGhXa2kw7uSypMSKksecrNYOwctKkI
IlTlUU5HpU/2PuUSiFBf3BrMTGWUn0W5I0H5QWS/b6f5yKUtF60RmGj0kO6lAHT61IrX8RB3MujU
vmUj71qOXR+usW+Dri4JB699D80dXxdtOjZ8rFPNJv8w5kJTSAWSbzx2RKhEx6BAJ7a1qyVlovNe
RPh++uAVB+JNWp6k3vsp1R7K3UvSOkI+4ndGihp2qz+7STCR/kREdlpxYAT4rqeNUnjOBSQmESQR
lZbkAsmRht5btTuC7EJb+NCx3MW9HEwPBFaiJyT8VEXfBNInBeiB06QjtUhQsursBw7HGdvywQ5w
eV5LYizKvNpGGIMU7nh+5Bw1jPawWwn35O2T8CBkxwH3izkSPPJ4TG4v8z6/z816/PUu5g8IjygN
ugSAmyRMv57VQccX6T5uJmAUtn+Mp7BzOW5rWS676edVsan4Fquq7WE6Rv0lnpgXtXhGEgUiRxCU
EWMk7SzJh5+r7I0PS/Bot4cyzqC5z87Y2y0TisUiy4hgjdwvoBeIVRLr53ZNvV1jkteUU3ZMCUom
yD0bSTULBXSUt2FqFGzWtUMIOtUU6/o8tZId2S/9MHCzVwRUk9Bbdkr5Sy9ka/DpRZOWGFmRdveC
lrcz0ZDGxqPTHmzQvfeCxsd3F7WUyut3U6I/0fQFXqzM3IQYi3TM/jzwaoF/sF3yje27GlMb0fIL
KOBJAEBLzWeVbDTJwhOWFC7vrF3toN3i469KS1ukN9cQLfaKH7PSK9iFmrs5L8OCVCpiSg213isC
MRy+oEPiO/B7WrLHEfIG2JjyipKBqKfV/PqI5fog8uEmBiMYaRPVjuV78diEWtMt9uj2YCfTp/K9
db3p9bcmcXcS5NpsuqB7E5RBg2mIxibYWMm5Cge5/uBcaiettQNgQxfVdjWqzmPZE8CSJme0EDld
pNo5psrU8ZEkw+9Dw6ZBaJgIJx8beGuxIYeqwBaWT5AdG5STAuLSd6JMIw4qabITVnB3BE6nT7ba
MsV7hXBDRmbw7dCx2/HlIyy9DpgSK3CE7fXPExZ6JW84BHgae/SkcMQz86wRs5C1xn9WRebyUz8/
RqrRylMnN/Tvvg3K3LL446mxoQWAJY1Y/oa45p8GqRkrqYML1vncYt4geb5sBeFKRX1ez8fZJ9m4
ZUP0RDxAZ/TuHB8aNwR4YL/kYsdx2d3bh9oc84FB28g95/PEYMqiIqSvDNat4AvRlI92JcQNEKqV
USLFxUTlGmM8kQS97SHQnxOWX4lv1fDBBaeik/POKDuNNuyBRjcZ5sLRZlTOS/Dif4SfxurSNzeg
AxawSprTrJD1t4saHUB1ClD0BxX4SLbhb11qj/DcXc0+SoDUoZdogrKozbS3ob8fWH+MQodXpunZ
uzDVwNR7jIfL9E+KgcSr9FfcEwzYtJHgCI4r3o8ZTLTZ6zZu2EhgTG/IXMaBK4zI/7E9bwRlB3DB
lK34vOH7InGAxcfCMGRQoPBUb5gzZN9Ieg2GCfzfOaiJIUCdbRd2xPwVGNkDqe7u/KIR4z11stT0
2KepBsl8cSXZ9P5ZvoJ4zEWo2+fLccD1LEqbmLIKaZ/lktN4cVR4RtSq1Hv1CXE1o1XtGkCjJXot
kifvvumJi5yECZdlyAK7QL7rS7Rfr3HaBqOpdcvLsIRdBpy2z64FY5z4rVEOyCfvYrUVxzvRwt2V
idS9pfALXp0Y+V0kmMLqH7reRc03N2trKmg+AUIwcV6JU5CK8dyJLi6v5SrK3eNSt0nBpKAbEmBe
BIR7rDusVmC5g599GgB2T0JGxW4LDJjI6greY8gZLWzE31ZRbgnr5XtPtHkJV5LhPvYR7BelN16j
tUBFW7pZtR/4XnA8Suzmw/7Xp6CW+OoGtRLqhm9aAhEOF9/0u8xilt3aV1oldfQ9uvuG6y1C0oBN
BqTsXM22YjekdM4dln//58RfzzLUUlBcelWETx0lvDjMLZmTxD+I9WihLzro8zBeqzdwtC6GCdv4
LSUfN7FU5qNWHNACDbicYzvZSKwxpNrUjb59frdccRW03DE3aEK4vjcG9Djqmm04deeJokxTY8VI
F/GhdQlwIfnOS98/Je2qaqAJ+fuji7qcby5DPTFm+OK27qw3D7hnb6dlJfh9PJX18MNqmy1Rp1wN
zBAJuoO4LwWEZdZzy3uz0o9NK4ISUK7XvtBeOIW1L1kqhAz/2gEb8xWGYEFP2xJZxI+hucZLcRCo
RzerrM67qGuM8SrOPNGS/vv8o/AvyVwUJf4qry9su4cG3dcmQCjuIjZaUHzLmpR3Z4LXzWN0NbvU
bdtct8AMxH0ux8pu0yK+Tgd1EUl/KXb1wxORvn9SgGwL26/+swyqJf404brNgIyzd25Y1BEvc5va
cnZiAme+XB1M1lSkeII59LHmA6Eyg1pLO/85NtRXv3hTbKyDbdScwAb2BpzK4vpUEXeKuCKY83s/
DBSfgjjeigYrsQB25QCXKflem51+YDAbB+zqSdBu8YSHhzOdRUaaH0X/CpPseQknjEFVnmR+axEP
YZCMxKYc219hNfLS2AcH1jVTdH8zrfx8ss28xWIBMYsvT8LqOpl9SPxojsjt3PKpT8RNpcmmGkAM
CTOFTWHBAdKCAEfWKH0Hl0JqJSe8OPxuTPhPoEl9mFKA+dqCTns/W934qOOSBzfYcDrnrIYKrG9K
erYxOXE6Np8mlDOBMoyiSpX2s1ZwL8CX43Pt663ANbbQBczJeMohTzJ6DZdvCNpOE6oR6Aa9LEaC
3iXrRvuweWJ+FhFerm/mxvFFtB+pbw02W4qXenh5nXT9myWu2mNJG+tuLGDWtCBkJbc1hwKrXNMv
wZbb21ONhuIrZb/tI976ssA1wF0MW+ld0BGYMIV8A4digD1beU9yz5hkrg5mYx7QqV8q5YBz1jCQ
ywraowLPINb0AvjsnqY7RXU5nGHr9qY7gfq3A5N4KMIO/nre47GH6MgPlz6HPtp8AgTLeNT4e/To
mRYH/76QF6+mVbUJjoT3OUnjWusWF+o+V/KdZWRqBhCOwQMfEblcxwNMPvHdYJLrn1t2oORTxLxS
peBeVldzx04IlzIworrkQi/wFobwp0pUbeGwRB2ZDxfy9c0vyhRNIZeeXvIlmlsi9fvUwyOjoFCV
qKjBxRHN9kdL6G2dWAHF+K99k2lGbuU2aBkcSAI2EE2jQ/lzKYu54HWu74pwW3pWZhbdDzmScMfZ
PucsqXoyqnsiqwCFiBxqwzdFSXuuEBZzM72QSmSg5lfjptrVzDsCH0CxR66XpXpujq7Suyw3RwlQ
3Hzvtnzm6PLQED5inbSjcpb6fx/LHwXqdYJnkUNur3f774P0UXxuKH9U+Uz3i2WpAnZe164koESV
MIRcyyIcLwCMcU8i/yHLnG8laiyWST1RBPnRoF9TXoqKeE0JEyJwKqM0uBQ3BiMVVm+6mgHm7obw
iF3eu3eJDv5oRNbB3pAXjX+V4eYR8n4m1zsr+y3/0dKGGdsC9oD/YwvwpDP4gAoPilrOpSFd00IS
iCkXzUTQdjI7TSSUkXRh9ndc1sFW5bnhxoRFiiVccagEdHzBxET3XOBRrm+s8Nr0V0/bJYNmylU0
mcQTx7+fFxaNw5FL5ulpLhJ58Kp9YMXHH0iJTo92WTKWWbLm9Pdur3zicwxd4wc0pAljv9K45hWP
9eH5axG3oxxwGCQmU/Y4Jev9EuExvTQOlq1+rt46/9XjX4Ww3txp0Gsbzl6OjfVjhaOnvJgq++SA
ELHiAYqd8O1+7TMo2ULeq91u0YIv7BqpwANnudA4n0B/yAuA26JoQcToIxXvpj+Rz3SuyB2VWGWl
VeBy+MoHZ9wfq3A2R9MldaQGRXPCcoE/P2D0oi5pl2GUANo6hIwUivnsDkJoDDsSaAgaWVF4evgA
7gcn31TrBEzVpTDKqbmSDl7jhO6YF/VxJLV7owW47Gqv2fPSnvhrrbTA3BSxBzg8vFIRmG9qwJhn
lX9A/LHRBrxuyBPohU0Cuib2hmV8ej6mow2Ownfc4ZhVXazSk5JNQ5oaJfm8mPPlUMqyh72rLS2P
au7MZNPR7jUZPivGwahYqeXadOe93JYmScffoyzUxWCLZvDfypMNcn+VuAUeljeO2kOFo076tyC3
5Xy85lN7D2chK9TFi63tPshl21YiYw7RDZH1m5oErbXdJhQbbX5NnSGWwRJt8sXqRst0e5j8x9NC
Zw0EXzjgnQsfHYco/zf9dbhs69GbKhMZ9fF4wM8qjzDhWdfw74J2DihPOEapYiztizAo1tHK/+fU
1eCksgWVpu9qmuet5bveGKMGFH3Q+eloFbbHfBBO7Dd5/Fq24MDbExGyQ3ml9pxDYIdJ4Mm40Iz5
C48AqeykTghKJcxWN2zfwvA247yUxbQzsA8EoSf7fdD3cAIFfhg7qfoaDGMpYvgXVgonxc9pRIWZ
hZPYBMXGjiSDKe79Fk1rd6j0BiCRjhR+9al4ns7CJSj6VQTZxv1V5DcLR+ChPlwOVLzJMFe/r7FH
x3Gdfpau/muw98+UlC1ZVzlPcF6rqF6Q7PuImhzs86mKErOX43Xu7sqm28ca7yjsnmG7L9xL926w
HEhodJySLUvi6wWL5sS+BhUCjU1/+05B5okNdc5ffooR5GiAjRwV78Un/WJyBo+8P6/86cvDvKqS
LWDLjW2bX1d9nblveG3zKtNrj2WxinF2Bp+fLbLoKWbLnv7ucj2LsjOqela6iYLtd8bg4B4WQGVx
41tQmfbmdi330MdKhbEC7RjCP/6MXjTt1LUSLtKEWUTQoM84OJ6HQwdm7khhLF4JIsghNW8LR6ok
u29qGQdKPxNjmb2CGXvjJRUbfjHtvM9lgapmSqXU2kvCLwfHDduofIX5VU/Zp0whrdZ18xDFvCqd
+O6Fb00xZh0ox3EUSDVy/aWbQjhchex5R88nX416ZyIgXZc86IE9R/BJLpnzsz57vVBPEP3GZoDn
sTeox3H9r/7+nue/Wkl7BTT7jHeg4FE9d232dccD37bClt4092+1r5LzniOL4YiaMhgqR9dYyh+2
Z1TsK3SzU+S7BfPV7DDJFr+StsTKy4DzZSNcD3TQmooOVt7Tgy9xAFUoM99VSBCPRhCfqa8JkE98
RKJS4eOxmSs+wZhD5r2K+hUa8vNvA0tqzunKlJvC50mceGfHCIfiRDm1r3655MwJ5Pldf1JWBEIq
0I0+kfQNQjxy+2BWKT+uAvHGO/4hkZrKeOEnA2VtgOTwdROAhpm5rsaQlGPvQMB8drDAGs36Uxbe
guM+HZ63HI5RszA0H1VVsPHJa3z5buhme6Mm24oHk7KbErYv9O6HE2nJmgHNQe076j7AFrMSygtp
F5iQd4KUueIKc36Peuw+5HSJ+BfjDIy54gRnaR2sTRZrUKvTAzR4qnXCd6a9qXeDPcjM5ScDxseW
VPMod/1JW/CfM6YBuiqaVekcT5tCUeIEeVIF0WL7rX8jO9E72kM4N2kHILVZGCopkmf+8JWqrrIi
cslGaxtS91gVQZ4fOow/5iC9TihDFClxiWyf8zfHPbXp5imIwh00+4XAtzSXulpGdbjRVLa+wvS7
pT73LBP3iiEU1EKG3Zq6F2pXr9QLADPSwvl76KeRJuDj5QjovlLtZcNLE6fdtGSXvBtvn/NH3zAe
FK0sksHlEkvjwMCOe2Z71AXoIK7s4Dmbm68NIs7eRWjzw6Lgpz5CJU4fvm9SrK3NyIGA6r1Vhl/2
Xsrq0MlxlISITsv0OxlszOc9mFmw5+i3CF2YlC8an4QuhDXJRrK2G1veG8q2Wpl0jilk90gFffn8
l9amvpMGczIr6DlawA0w+kwhAUTbdXDTpqNjyJS3FNEwaqNAQYl59le6enHt3ZDemI+Wk0gJt5rE
/JzCIvmjtovyQ4g95O1WjefDlhtMCpnF5ZrDH47AEooHWnjRq38eqTVpR8YbO2MnPhn0gQHp5Grc
LnfQpdlRzGS7tC9M9+dh7N2vKU1UEHgZAYdzdOR5EOzwBuq25ObnlBEz/uLvJ0hev4UGcv4zgNO7
S2TFp5rF7zK+1z2GG807BCTRgDQr+9MM0WPSTLInh0J0yTgN0Vi5c2D9f9sqTi+6cShrRwFu+91n
W1NEfqhGchV+XsjOWU1XQJuw1O6oNjmYH1j3YQyv0EtAd7BeDoDCFSUDAtU/J/O/6Mz02Hy9o39x
MN/wEsP1vizXat5mVjkhFIQVsX1XGoE733fUhG6sTOcvyOdwLgMocdUnMMeeYQ8U0XdeNfrYTtR4
/5SoG3otplW6zVy3FGnA9H3tIGbPW+gIDaZEHYy2jcPu2mTmXPC2a7nb60tJ0J0grx0IDM79Bbpq
mGQeLfETvfyY1mZm8L8HlUdk6xpOELRRfAd05W8r/HphO8MTrDIaTp7V1mOVrDcT9KXqpl4lb/Zn
zyarBqCn5mxHWOKsuQagk2IlQR6aNbNlWT7MR1CydZHCJTu9NaSQ/QO/h0OHDRdYQ7UD0IWVSMPu
f8JLJBie2vOKHL6saSunPLYUu2OHWoPc2HHwbI+rikGMSv+j9Sbbxwr7yDWroR7TBoo5OtWiTuD9
k9viKuA0H97fV/UD8kFnuv0CizzRG0I7k8Wldn1iAHaSKDAoot+uBb1gZrkcOxCrNplghgrJQsdS
Ws/OTyVNf7bMWVZu+K7YZz0CSjsYniguue1qDq2POC+xMjb5IHW6pENS4K3TZg50RujtArwfA8kK
WKtZFJPThVCHSKr2rsCNm1+JFWDDVzMEbWQwy6GBItCV2ZZGUERVzUMHuTAuKZ1Dmsne9BADvvYX
rv6FMB/7WLOJ4ySFVnydXJwps5zaV1boYvhc9yu4Lnh6PV+VSnl+tqprMXc5cZyWy1ywOdOviCQ9
IDgm4dhjM8lN4LqZDqaXvYTC5qbr9eOAbjFCEnHMTa9n9KWw24A+12u+Vm24j6zfD56ZvIyWcHz0
wzzCjpfDtQvsFLw3s4vZleVuIMv+BvnlJvsyhjHkFAhqCDBixucGVRwJkYgYcuVdzhJHb+xAfqrx
DAmnDz67r2Oxw8NeXeNIHXQdaUTvziU8S/Yjn3ucq7OBYDgYYNQwp7zWdsN1jvQAVfSFPVem0zvB
xZQV4x2Z6yihl4j/7Q33ujNQtdgAxR++QYZ8Q3GscftIiuZY/DZlnBjTylkV6+cUPig50fE/M7bx
SAEn9oEZcPodPk/j4Y+C1hBKcK3zcKWybjOSHitfIFlvpYTocgEaU5JXEibEFq0TFgxUiwG84PiH
4SOIO1Ix252Zi54TnwKd9uLe6OO9C5OxxmBFbl+BxscmAgG+L+bC56kN/rrla0kpMGSJrCXm6KdN
qRDo8/o81xXQUT9rS1GKVcRxIE3tQlbBlovu/CVED3oiwjRYuDlvFwj7MXk3AJtzDCM6e51EGxI/
kTKXoZ+uM5xtPejnelQvl8ceDmCya1Nw11+xn9aeQpvquTD6AdWEqmOKaneT49vOd5f/GH/FXD6y
mkC6nbC4GLZK/dI266EKP5tsBg1lE7coKF8JPrN/bGJ+ZYVqNm5MLMrGh36iizqmRiVHYgmQUqR0
iKARIysteoq9j4QHmKAHWGDRanM5lgfnwG8VDWiflrR233OZSoJNTJOUYpA3MeYb0df5oVzX8ruH
f3CiTRIjtN03/qPqBSgkvAWDL6Gp1Zv3GeH6wUzNByrKxL7xv03X6JtCRYnQJ0BtPxeJq/jVYJ10
mFo6QaeXC/pELki1Sxb0vAHTclMnCAPB735qOQFei6s25fffCB61yVBkryRngWtMKySSFkE2UIzC
AlVBkPt9+zRzvjUkixpcQbkUbvflyt8ARrQJbONBW3AP1qHT5aB1zoz9TxajTA4xj0GSb/aYrAt8
lY0QhoagrPd/i7K0DMBuhDklxb6bSyAZ6wwrFTItgOiV0Bx+slEt10xgoLGY0+yrJoWnhzFVrJ4U
ZkUjti4YaLDW/iCkZiHhM8/Ii6MyXZyzuObbp+NfUv2TagLUv0kG3BnKA/wAkjUUHObIXLSOeHMK
UeuSzgkQTlqmYuJyyZ6Wnsd/Xg/psnF/SgNiE9KfxSFgAeXczhf3BDZAXjfEcBPp972CUwdUtEgK
0gfj0zcFEllGloSK8uiHupaAWgk3iE9SiKFi3zbv9inZ8J1AwtxRLlJtEdazG5viHF2OU4j5JgMl
IZ+wRk0JWHoy/yZz4hxos4p9Jhol5NEyZhrS7ERWuyBREqltTVuKNoA1KZnWV4S1JdAfXA1pryat
l1sLUH8Tl2EmkF3GIGFLVTd91/FovQEM80nWAVMHsuZ0ikSSludhQ9bnz5AU2stfrOsm6YmFktao
Jrvd31pG3UDXrUgd8FQ8AqP/aN3uAEF/Wr2seJpODKjsU4AR+0FW47P/zzXH+L84I0bSj0SG8MyB
qPsht+9IubRew44Bn7LQumUe+DHbhB+fVmsorg63KR8f/0NhYgEr+wNsgShpB7qQ2jPUvYcXchkF
kEsNUg5zfc+dJ+wl5XmKkN5izgT3jTQzS5mlJBylJ/ljPwZ4e/6e2JOBcNcUqWq2wyMV1t63Vbwy
v7Fbb0cCxER4LqhEAFSzAM3kf9ZOfJIGvEqUjyhur+/eqs2dPNmndCZ1U3g8RO1GLAX+hsBO5vL/
xr7vBk9EWGY2z1LXQgJuBTzn3h9Vj5GAigkH0uHmOP/JQRNEqZrugpZeWWh5fibqRvrUA/IyJQid
jarF0a1QDhpoqdGA1SG+rfHGUYFY8OcvmxqowzB6IRmqdEx+QnUUd9vz2ARwXF+U3YHdsLJBC/xr
itqk0LwCAZwR7scrdnndk0lNvY6xub+DSZcOxDDmJzmsQh4O26pLIC1k2Pu54aVsyjvFDhR7q9Qx
qhWBjBB+DUD2cA5DzjqBVs44LPSePI8TdqMgfPyv4j8+jw+zpPmAzOw5LpXHTFo6+y1iRqsKa4YT
+HKlNeMeao+f8oPLWKMhGTJlXF9JGqJmqJ+eZod0j86N4FzJgYkJyAAQpbQpVHewsM8wF6FqDhE4
zOD685/11YHuq+XtBTvhsKifx5nuAzd+V/G2IIeiyLto4+K0aIwmi2C1WYnURYQc5Q0KRttgPS/6
r2uTSbA5V4Jt9592El3U106PCNdP/QK25FFhHwkOSOh2k01uN2JecLpp2o14Ld3OSfkvQiOWqvtY
AWxv9fYyiNUPCNMIEUd5d2MJHPKqk322QA2n8mpQEmjX/b5/hkJURT0pPZoWBarOGSr5uLZjCwfZ
0zraFARqjQQTTahBzKzE8rKhfXUQDGq6qKUoUk/FYSgLIg2xtJNX7LAYsLL1Z6ddu0u6klODOl/A
NqXdRGeeVj3u1yUATqHnwSxUKW4rR3nM8VOykcpWdT+uXH3lJDyBtvkbGvElZipeK4wM2Zact3AP
fG3BD5GvixKDfn3n0x/3ChBT9BEABQkGMDr99EIygJYlNBAs98XduUCI48cFDoT8Cg97E50Y1Fak
AM+xy7TPI5Dv3NoTuiqsHcVn4RHkXdj2NsnU7W5wd1CdiR0RaMVirs0SqysXteJMdAJXnCuiwLfm
My5X9TL5lcHPCSZQmD36pk/cG0B4dvaFAMw9ha+lZyZTrkJDiU2HMXj9sQnsig2/tZ3KR4CXtyrO
ZZY11DK36GAk6HMGeXOTBFy3qX0AxJXI+7G+sTLppBhCFL14RurCa5lPL2SqM5Itm6VbvWEoJAXl
p4PxNb4qGFpnzC0PZx321ML1X4NDEumOu0ovWvBZ99EzZy4sfYo/cDy6JagdILROMzx3JS1jIbC3
S1KMLDvUjALgkPzI/gOPXNJBYAH7vWyf1z1DIAz0rQN5trLRzPoeDsg8yECJK8VMSEK5KG8lECEy
RPfd+OqkNrVT97MKzA78dL9o9UuHQ6oWzknmQkgUsYrTxVgoaR9AGQgrsYLT+9qdqmdDtRSo1aQd
xwJQvfY2Ky+ELR+Aax9d1ByWWvORBz4LqgGDquxHo9be4fUQuFeAigSmHtMx0sqbCMMxOYmU3kev
tXs6vwCW6s3LV+SYOdkXF7Qaw5ThXc01vVzYseOGIelvo8dCRBQmrDSUC71Ls2bxdXZerwEjI3lW
Nb4h3ThY5ESo2tu/sLr2wLOn8Ffnur8e0oKT0xh2RXFoI8yhaVnjI3Ir9O3hglj+19dP4RibjWz6
lzmhUvSoPDeII1T3LT+p2UBLztveZlls4zHBevSJCooQCvAxQiL8WkDh/Von0uN6fojn+kL9XcKQ
4Op5AFGn5op+zhFym6TkwAT1KSt7c8pe6+wBEP0nY2fqcPn8lBxvezKX4xaDiUBbgX3FJU3+DlWQ
BupoUz6nHx74dlmB84zRs2SRSTSIt/Mnui2Q/x1KKIMnLzxecEY2Do0CnHHS2ggevTVywCeeXSJR
jyc3EfJe6oAM3L4d6h5+prirIisKjq80B7MWuYi9z86Pk/0W3+voVGbmG3p9HJ3X8K1uVhbxvH+J
N5cgiD+Jb9KBctyyD69NVj1rKn5Vm0eslNo86WrbM1TnLMjujNK/6Yt3iNXW+pPQZoWzz+JjaJFA
XV+V0zsFozSlfXXrOuBo1XMaskTbIJxYPcI5ln209yt7LxLW4/81yp6NSTis9LZcQBLWHsilrM9/
11k4nKcg8neB6ItihrenQ5dbjNcC6QL54rAaLx6tuZAHLZjrfxwgtrwLxDCzzXm6K3lDixjfkOPk
bl/xMnHQLGLhp6nwMJ/RaoxeGzilsfRJH3MxE3pCylRHNMrMdMNY/LjzoxWVXw3ip2tp3Uxhorun
Crfmq2jy/CB8pKLdQSeZg4gW8F7L9gvOekvIiphCahoJIqo2o7XbeoU1Bs4lyR030vIS6nMPCUtu
8G6mwoYxz7ZXWC1NyAY6ciZCVfmdKoQyqgsE8pUE2MfV33kc2zhFCQf4lx/aS//eb/+AXpwLFe9z
wCv+eW19FtU0cEnvJC3yflPbt4gZIEloogIT6l2R1aZIBhT1k5NAr3z15DKNdaS8V/j+foa48Sll
n5/+clNogyKkvVmrmy05kzq7Z6bAvAEYVlULTTjon7Yr1RJgbJQerTA6tsdmHjIG2rMGIWzgcxYs
2vM3EuPXuzOiht9B0yxX/4UOcdMQSpDVt7x7lPrLu4Aba6O89jOQQrmfErrvnZye0aopVxtuaNOn
TpH3BM6zb2HvkW8efGcdbR+2jQNUKpy5ymy/ac/KKtvDmWb/hP7FStO+6tP285GKqM+dO/ix94Fq
xNxTU/2jmp07rp76F82O5pCTDf1evJ4S+aVAKWQ+tHHWjDJYEb6d1+X3fz6uvO76DROPJaQ9JpD/
DQPHzkFdS9tKe4FzSNqcA2K0lMHfBCwjnCGOvZiZDTfijYsRu27eDeoPhWdOx+a9c1bEheZ69EtL
5ytY3EaQAHC5Ui7MXylc/DvNmOWUjkgN1V+U7Tz5P2wJtZrrw2BTAqSRB0EURPPjRF8Yj3+DjPD1
TOD3MhQFvHome7YyES/HpdfdPJaGovbRtUUGgwmvDiWzeKx1U42G+xQl2P4fzseBtsFnLYIcGght
/FU2+FivJ8xYNLAmyDjmkRjrxykfM4W2Ew8UDdDLPl9IKtVFef0Iu7a/KPoWHnOURRPckiBjovFI
uR1IPX/MCD4Y8EtS2wmO3yT5HZrugV7I3GsP6/xD5Xe6q6FUJWqKLLhSy5iUF9J0rd7peGt0+Qtf
EUm0wyftPuoq0Z1DPjlTisVNJsSZy2Jnnt4/IKIpG+XMs41jzLa5ZHmcYCwpihxBS3Fp+ltklvtK
xKAxx6KHAtM443kv7YmjUllWfkfh7E3oXzDQVw31SNACvXePehEJ48Y1iSjHYvHFkjYita58vN+e
bOoszZXJvtt82z1TKXthbPCDFC30kBhxCqsWyUuDyQzix/DNOkNtI1AdPaXR6R0l4wkROIbKV+lO
mFv+7PmhrRpScj+NNz3yYYwRL80He9iPKIkuL5oae1yEmY7ygO2IaG8GcCdfhtc9/WJCfNIs9SZ0
M5m2Et0Bio/sInObvfavvJC5ehasTrZd3ou3j4Meethbx6wo5c8IeixKm71MpB5x3S/5NX/JSCo0
9QN7cZAbLtWAnGdduCgDdLy9nGoevWCZTmLjXKiRnpdl5tSVrUJhxX9WWn67rPxXW9XXFlHTzJug
N1ahC7cWoc7ikqeoyA0oelWuBhQCneC6Y9kuAK/39boszHECfH8cM0bA9vZM1UAyT9rcJ4InQMo0
cWvpDQ5/UX7EGtyQGTaI1DGP34vsbIw3fIHmLxVd2VSePRYNss/gsCubD7Dj0yZD3KCnS7VKWWp8
/PCu7Rw7iw5CGi0ExYZ/2YIGuAp6Nprl/FrZt9qJUJgTpbFQJiMfnskhhLaOFqHFXDcCydR25CBy
KO4sZmIXHWoUpgUDP5CE+bqwB6NnmTFLIATv0LkOkZLbLBXt371Jdcjw8a8QEYCUAJ4XF5DPS5Qg
pmOZRatPXJBG1ePorotPunWmf/NIuqlIJ0iJceDfceIR5UO5dn105qOd6GE9uXeRgtgXLyqpRzNg
z8nJHifqAFv5nfcG6dbcqik6Be0hhcIqx5k7Xchoco3lqBaLB9G+L1bK/OpLqrW+S/e9jeWxkVvd
BH6FAgtpArtbmxTG+Yi9YKeUNNSkyp6iGPUaBaxZo+ncarAYgXE9qms9drPGIwtsVAeZuR9addCU
zASLc1bzbYWU9zJFYzFzBTVoArLUCele8B31Nk5M1B5ttG/kmMeFSYv6v5igLR+3C+mQELuutAb1
ndLdhtpU1Afr5BCGargE9KKqnDy8dQPSmNsUHNVC9OWKsz17+i3SCuY8E9lQqeJM+9j0D7pW+t26
f1FkrOTz0auJAXJwq2ItKIWRxtylTzsNWw6g7/LN5RyT+/1MFo0vWWbm53AjsWUMMGc4k7BLhsNg
2yW2g75ZN8lbSQMURY+ApEFT3A77keeQ1FIw7xM5dyHjQoxihNGOyV974i/8j4tPnuvBueMsPtKz
QzefnPkWb3XSI5bG5O7C9fcZaq4sb7Q9DT53rYIIcsiRjGCwHYp3MWG6lxOTDjBA6CDfLLjxH3+M
aCx+65I10wPTSu04A2Cu25vp5CFE9K9s6agFqXAibkPYldCABiWKtAYEON81rzj3d8EUAetcZNxN
ye/YrJOsQffbXNobm/BgyVwhDST7ELjP3OMSF8voPxxK8oqpRuGS+6bvV0YdSRlTALFHEChjeLXG
mdNWtX5zgwkGJX3kdZcIYY1hbuVhA/q9i5xj4ibjinCqd+lGfPdMYmlU+VaTqk6AlNuf3V3kyioF
pc5GN0NSc3MDuh7XAhlYVFQE1PbKRjHzhVk8pphiC9P7Ic8eK79f3aBCI1YUczGC3dbflds3PL0E
ENBlGiL656OPWf58AHHDAmGVTDJ1mxJkBdmx5ueBp3oAQ0Crl8abt1X5LL+RENNsyE9wisBJZqS1
DC3d3y42SMomHWCAyD8eUoYLIhHox8Fdo0UQ0PBvyFmqplt+357fdezFnVCmEv+SWl67gm6FjwHQ
Tmvm1QBDUBwN7S3fE+hu4wAgUhNWMIg3hlAuLbtkh+4qm+sOQbE3uWBR2YL30Ny/zcuT3V2hvX0N
3me6ykpMrhuYdFSnAD5D+EFrrx7UHCV+eB/GVrVgo0/y6MOVg6z72B1Ak1BzBLEYqkp+I6FNEXwI
nrJYscXzauR5PUsxkgBaKmwzB7QaSxCR+PiPxLy/xUNbPvjw9v2D4oAqA65S7dDCiqjvbcBxcbyO
8SRYMBSrax8FT1FFqCDbqif2flcn1SpSFuFPhnw5e9GHlicB9I/LIGXeG7Ols/YvJ2jIAeIAKjiN
DbpYSUfNuYParb2FONx1vYJmsz9g0lKBUfVhqKS3/+LXiPEvwG+GbpK9F02AYC7y6ArpwfPnbwQq
/6RhmFvrS/7BtHTr7cXSlPGaNZnB0IYfybj2QA0OkZ7+P/4YEGQguaHsodJXsfogdN6Sbrzx5xjJ
bPiT7BE94KXGH9b5ybxLhYHgOnU+cEdi5EGhdiD5PGbVAtDVF0HjEoUCCk4MNa1EDbD3Jd7YaDIv
rNKRr9GFmbS0yoHNsdCzTdK1q5C0tGftZoho7m7Lrmstkvj9QyI2NN+zFk6xG/pTudBHRIuyN/ct
sOtW7AbXXISW+Ra3TYtKAgqG+bgXrVYiuf3KnLka58m0WT4So3EVsclYL3DoH9nNWZplyiOW9UJC
0Jw28CbBA7/xCqO30wcTrAhzfI0M4yhBmmOSGaywJkAWbPtEXlMWpRXrIrl2OdT5/oQI8eWaVYcO
kIzMUQnMMSEgsU1x3zL0HtUY6CQo1ixZWxqA59peHsmRgjPlH6XvKawGL6krdNbjOIwCNr4ZcExl
r7L2VKz4F09MqMvoHad33gBeJR+YKrP8jfkM7OybK5t+FACRLHgb/gOheK9UzaQwrZAOXThhuJzu
/YMkI8bspyvnruIG/Q1eMh6FczjCCznvkehhOPkHWh9ck+lchU7OUup4q6olr2u2uez7vVXSirGv
zjPbj0XLAKd9JW20h4Gd7Q5gMcE8xMEYADt84iDhVJQTwsdiCHgTtEMn0QIbvjXJOgla7EL8u79C
Hj3E6wIYOkvIMc8o4+mL/YM6J2EkFfssHV+1bfKv/4VHi7BJMs7U+sMaZDOFZC8kY8thGYW2SZH0
Fu3FwahhU6ETwvr2xZOOX88if9c9qVZMSeRaoPzn/nGumR4Ytkcu0RneyG8DoTehhMhg2jm8LNFS
Rx+6XG4g7j16zO5lwkBiLfgSlXqnF3UdF0LkCzglBJ+srSwDSSLr4neAb/03oHX4U96zo4Hn71WG
f/xcYxNYr0INXJGlHYbLAxLPsIxb/QsEed/sIBaMjC4u+14F3W4NuZY511bPAFak8B5TbHi62jE6
8tknJ6mUxkZt959kT69UZds5PnTl+hvQLnVlMV2QC5gkfqK/wgZbNomgupRavo2LzKEQCspPLMcW
v5XD1cYyg1FYW9zXpw63m1bP3bCEOYHlwuP6JERo5+5YN404sS7uhG7tZ1XGE2220IL+OFFKWX2S
yGzTOJ5zNpuMdPonNsNBOxCgOoQjZC5I301L+0hQ2Isnot8PwOZvxZKWc0VkSdGVIyBjDpnxf8XY
0rTvWp5/me09ARU2bSjp5Kw0+18Vn11H1YgZt/4rNvS8hXw/Qg/SeDRrkr9hC7eBvsTzYdE+Cu5n
oCqb9uYF2oDybSxelYQm0fElDZ/WgR08T/TVMAXKI3JGjYH6f1UFh7JSbjUWAJiO/mUKWUJqygl8
PSaDaAQIxxghqGRoWNUPljQKgrEHWZgbIfJF5Jz/fiqFt04tM6OBvHOJlrgnRlMdacUW0hWX7Bmm
1kYNF7uGAtWw3UdICGa/q2r1YgGQ2lj9glw2iM4r1rG/yMeTF5Z8TYw/7TynpRm/HcsWE8b4WvkT
qG6unXJumHpjzgqqVBDmi4pYWS9Trm/2lxPZ9lvaIY9U6jU69OT8EkFEtcq10GrwF4cvcHZy6Zig
zCtocO+v7RR7Grixq4fchVhjhUK9AZCuTp/jc61KTAgnXeXrRtHtSViei5x69w8GHF7DxyLidDwV
mzZNLE1pDJMfd2L2fBIEgpCHte2Edeu1DVDG4WhWSM9xR5/prB2jAka1X5F+fuQqBHBwRKh7/Hzy
B392jyfQXfjajw2igGmvEtjF5RNi9JukMmqatzNqLJZNFEKo7k4f6585pXNP4uyIzw32qWHLE2mt
HJ0m7gSLQ8tpiSMeBRlyGvrdNH7cj40k/qOsRmHdv5iV0nXh53tzsmMi0lFYqz2myFUfR1CJG1Dx
i94aUN/SOs1KmXmBlLxacjeyPendv6N/EQnFV59adguFQk+2zoYeYulqsSHFKMYc3Whyvi3CqIk0
toX0DnLdlcgTVEzQA5lwKDzHAhVtKtK+7zCfN2dcgMdKdX0Kgg8+Z0538QYy8aF3XC0ZrwE9JvYt
KcNTTtbdn/rtOpdTzEiOKsA1JBf1gyMUno8X8UZYUr0JJN8STND/zR7t/EjCO6DIuTf7SvKcKdwd
czRVljfGyfNu8gT2EjYgtAhx/Ba4ZNCfNhNgC+xkwdCdIC0ue/QJfwJBOSbDhLMigLxIh5JUCRVg
X3y1gW5JHHMx1ApZu5QNuTTVhkGHOmz4+di2zOho+ab1jC/MxnpQHCMMw8R6VkPLWu5/jMJcNeJ7
6Xv9WBz9szdhaJ+rR90sDCytpQy3XPfZseix3xlQH/bTlKiKAVEEK+2ERXDspOUNB92E2sc/Hsaf
4E/PC0pBbYoy5P/S5i/1CXgo5hqso3MphebSWIGNeibLaropEDvfwch+3KSdBqCv4944KzMtgEAR
QIyc0H9YE75X0xLFRKKVy7ia1KZTe1vKgSjDLjLdjV0mlRV/SF/kKOFh7ASurO0ZUsKg2D3Ao7Uh
3hMGAA8Iv8cIao7PIaYfcKBMN4ELSOnHXd0Il+zrC3zLET+HMo7Ns3hnz+Z11Hyi4APHP6O4rFGL
jENUJbPNbvraZBxUVygQwXY6GA+Kn2xwEgfMMXZ1sLcRDlVkgh3iLvIt2ECRY8SoGF8kyxlupUxw
dDkPE7EVkxQdbSD6pFxGtMtKKs/e1LihQ+rzQbZHFOX5fn0+FDDp0AUinavTjnmzR7MPePm8otaZ
6vqhihXwmbwSx/eNQkG26yxKBMOMPnR8GH3PwJmFOKijfWZvlWlU7wkwG1KzJ7PNP16iNlfqfkcT
VAT44seKz2nEtEUZg2xQGzCeBf0308Lg/Qqp5/1xCv7ERWuzf/zvApUePfZoiUZPLjk1ZJJpbm5E
cLxmAs6/ja6bpwr2DyiKagkFT9P+yvUC6l+gKTSY34Nl3MzLWTT0s+ynUIbhXQWbPFYcRZo9PFWp
pcXwhZ9Jh1rp5Z7HCcZ3KSPdpsYTUXHGd+oXZL6ZtYa7ofd5fZbHgrj9emQT4HJMlGxUC8Tfal2f
Lp6hAPpXXyqE3solGN5Oo230Tww+vkwJJBqnEYCTozY2E9V3aKSRdiBsxxbgG8YBJQ4En+TBtibs
90+wrnL1V/4fDc/CKX8TCe6je0IP7UEupMa8crRMDibo+hJyG3B4WFQ/zGEk4VaAMKpe2F6/UIj6
EZbFfGV9LqC92LLF8G1qjBFJhd83moiv9B7jUesxx4K/gwJfiuN4NiSdMksEFyMEyQr/Y7yv5bf4
N+pGzUcFGrL08+Zem6E6bbEBsNWRtLHW/BC0P0CbVvXDlgpAtEpniwMEXlONo+A1z0zGTxwiynYP
huecRCx4ArhsvGHOIDNlFryQrVjy+xDzVyKHKaW2VqLH39oOa1i0Jzh64K6f6PDR2nZ5740YJbI4
gwv64XROza8BClUrXbJHGCtrx9UiretMZ9c6S1fZjSebPwiZqBs2xOEm4LDpaBUuRTVdInfw2+eU
BZhRZ4FvOtUFykKFa1/QS9zEDtPZTFJrPRj6SCmDVA1HHE0/YX7hq6Uj9Vd8EnlndftOM+ZG/M2S
bbTdbnKmZjdLm3JZWumR7VGsMbo2xLkZdEIH10WCjznWlm+bIoeckxJRDQJeBopfglsWfNXB8onE
m9uIoKi/qYHXT7mADAzNohzqOSq8kZ1MwFfexwSLnCCY68u+UJJg+xuiz+bh2oRMr0Z2i+EINs6B
RdRgN0XI2pVEKaWI0NZD2kRtb8PXK4AeNmS/jJ4DuLIyM7hKnNWuM/lnwBIS896FIcvE3Psz97xm
pDtEVLV1Yz3b1YyEvmbRboWTdc3ktg2aMtfwbwg5dfeOZmEdMK1iTnZxFGVQsUl1evCElxq9oPxQ
MX6UDIJnQpUtkHDWxtw20O18DxksFAD62Ugp8VJkSZlL0nE/wCt7pM1NAOXUBjp8ZUp2iIpO2wIu
epZsBSd8w879CfjfW884SMZ1Ix9sdzdmExbu439WSwq10d/RJolCaNc0SyPyVdG803MBSN+6oMnh
DQYcFIxk50PSvZpXqB8Fpb0VkFTiVJGg7beSEtjs5YS95FdrefRsaLuja8Ox5MJg9LsYbw164qyU
AhpnkfNVHcAxFL/65PwzaZYhPtWmpUV30QZv9kTCDudby+golancd2s9qXUNr+3ZzeZrYRiM8oku
V2s3oRHseT1UmtRVPwhCpk3JqskGDfLZnz2zT0zpvpohTIou7V9oZZdzY5rUoEzlGF3fSJAYscoX
TAGahghp1zzyQ+495r/yWbFfdYL4RyXdcgN9ax7/GFR3JZJ1tMKyCk5vlMnCCMeE2igUn8RJEo1W
Pb0W3RFMLHWxE0cnxAsXvXMMLaJcAime7wuxUHAw+7TnI7DgRTLsHwK/Of96EddCccmg/ok6eK+5
+pzsHjrE7Xy7IIbgtViOz3ZeCPnUp84w1dF9oR3SDz0oBwaX4VLEXtPOpNALMGJry12XvU/HSvyR
Ot1Os+fTVGA4teLsRcyCW/41EiSRfAZ0wv3Q3LLEQCuM0LS83EzJA4Q+jGuqvD26LAToebi3AQaN
KNMhlf2NOojf9cgIEOBtR20V4cH34SXt6pefPfaHrsKqECXfT4247sbg05e7uQHYXz6siEu0iCP1
8cv92gJlFqmOyDTgT7uRdrpTk+Lpp6dLKRItpFGVUDRSoRiB45VG9Cf2jIAPyV1xrZ4B2q55KTD4
ByWX9BRka7zA0UobCj1SLUBCbCvQhbI4ZZcyV7Jl/WoKxbrkT7i6maEx/grBGmurb9Qx9FWDGcug
6/TJPOWuidIxVFuEuKc4naKxejncera1XRiJS/4HjdNCkTHnJFvtJeV2Z3FtXyJ66mI16JCR4PS5
3jNfDJEuXpDhvodqJhnc1Iy+75uh7+eOwHHjJDL0qoRR1Ab3MinNGoCunSGfjtQzrxJQdF/rIZ6p
kfOb+Ar0/J7Gt+dKTwnP+VTbZKTmLZ/BWVUY6OQVt2AEzupNZq/sI/EI52k6qE3yddbyqEcaCnki
HQFjhcUba3SfNjIbFGBiegXpXdvjZ5rnleaE5iq78vvS1POUVFplpU5DJdTguubJ5DNL5GQZoqxL
B+v6lXv4wLQHGgRQSAGb/NO1ebwWN/QC9yRBwXF5rWu2xtuD6JaoMtWSMfm9BDnDq/aQOLbwMW2e
gZpkZ360NoDZKy1s5HdMD9UXJTLWD0ib7sQM2Btsz89V1isARWaRNr+f3n+SQVVfLjoESmEPdq69
glizyI2UjZYWG5xt5xtjFSd6x6eqHf6k4MOnPxdPQYzEtfQ/i4/TbyP0p1P/KctBAp0cfXYk48IY
2FRq6ZJhG2aEhCtXBiPF9NVRAQoio1ZP2/UrQcFGL2eLwua0MNqaYIoEg0WEysk6+ZkPQ18sPkg1
UErHCKXJ/HeLgpXXUnd8tqo7IONT6r5KRciVPQv5kwSG0EIE6szDxOLrHMEqXv84FiL+qwnhEHoV
wWN4BdS3HYGngkQKP+zLzp8T2aUb+BqW2nvEMQ92VazsP8YftDNIr1+0HNwivkuCOIntzkrKv4JX
pnwiQGMZlgSJrpi+9C9G0XAtKPpg9TkUdDg28ERUseScUHzW5X/LCJFSMku3tEhHBOP8mPc3HbWJ
oy/39K/NLNS6ed+UM29JeARoToNwa6SNmlPmg6pzoNCjO0uSw8PAFdyDlXIHAPk2nMPSljcjWkVz
8DzX2kt5Rhvy/QPqQn60JlKfT89MSxl9kDPEVljEXTbfMKLXugiZa9WEs8SJMTKnBrEr1LA4GVKq
RSEYTSE54DE0jYfgE1G+2/ycGcIFCNd79wR/Xmq05RjOD/E45N7SdofQWZIR1BSQ2d+ldCGP0q3/
F8Lt9TYd63zesIus2owpH8WtrGO9puP7flZ/N8WNemY1suHZpMryTc4pTJvgWepW8RHXQTaGZvCT
1hLj91xuepD+jn1WaAiR/KLH0y99U4faY4DzDkvN1/y5M2LcWqs3YpBp6VyzVkoLuDbVzHKCcUwJ
jvs8IKHlev/6gxCHOQfiKQZqlIyqxskkZ9FTWlqF21dzy7/4nAM3hYkEx7glrdanEU7ILQ0LQ69M
mGodJuHdEbpQFoRxiCMTDeP1QbnpeQq/2BTF3FisVx05BQn6vFB2odjKLG4INANJjY0/fnB9oIpS
S5hu1S5jdRrQWL9NE96pl7D00P38dhKB0iqb8CkvfqynmoqyGM0hI67M0aFVDhpEP+DMB99dm5xu
GyAXQVgTqLNcoyGgoR96sfVaEZHYK7Kt85wKizVuVM64ImXVKPyiuOB6Q+f8CrWjRCSKKNzzP6Vv
kUo+XuvGOVzcqikbWAZ0aPieZljz7Vh/cR4/iduc6dDYROXSDjExwvu+WtKfb4nKNJ2Bw163a2eD
YV0Wg5tyX2xEiX8wEHHNKjR+bStmaHeSbH4oJ+AaRLquRscibmxpjVcl6og5+CLkIc+Cdw2fQRMp
Z9ZBpTWveorcTbzFklje6eFz61G6J4OSLL1zvdlIDuKbB8UA1UmAB28Dh0b14LeD9beud6WjaYmY
3x8DcGamLVCfpgmnGVi/9IeU1dsO8vHTIfbhPqt3CltYC65WRFy1O2zIaU5XLO1Jh6ArECl0b4B0
19BWNzkvjYXQRyLnmlHFdTwRCOQKbvHykL3YXKfvXrHJBH3/2E3knWrqQ8Tv+eERcQnXXgie5tLJ
djksiKMCMZjNxeIV1WG7Gv+ZDwSa8eReZ1rWi8iS4qejwEYLm8iB+V4oJiuiL8vo3vwUgVDWdLaz
r/vYrxv2EI6Qbsi4lqRN1auJdVeKGy/8JM/SgJqkAARi+WqO9jSlMQHY0SV9nEYRwlxlenjnSCPl
bil3ikYZfdzWELXF8BJ0ZC1eD+pwM3QSOzEJm4FQDWXyYRn8dPWXjU97/jtze/8er++W7VqL6Vzi
mLd98LWUA+g7mXA4bwh1K4o7Ko7HHQn8MDbopc1vT0C70Lf2Z8os+0uFyhC0enh+/mQjAB1xOYN+
9s7Hzt8KMhZu/pr8puhyw/qP158USwZrSZaWe0aY68j0slRmW24IaohjBaG6mBeqgf5H4XJHlvfG
RiYw66hhYWPzCh5ZpuDy1fWEHvbckbs/ufzqmEgZKHJzha+jg3lwWc+YtF499L2Yz02EBoa5WvhX
Gd6yq3WVdrjCI8bKLcsEnSdISd9A4XQRT7Q3WyncAEvBGNGq4/XIywE0NsUVPhbtug5kdXh9TSo1
PLzfGd4YRseNGwWmy6hjFbPxVzOOm04zgNHuGiePypqi6VYYT/zp2IXLg5g8NEJMmFz2tXUuuZHP
AU8BwDuryv4qrsUi7LtUWIsK8+C4nYVLUcx5rzH/c36eziyZ4j45yIEF5KDdnCOgDNMwi4fMXtqp
he0zTxRX5HKxFefOp/vYnBV8MaKUhKapUmnL2jbZzyrPQaOz4tczhlEjiqE5cykacCYYLVjRJhyT
Qzf8+BYPtS34csyTNg5iUYBYVwjt3YUQ3TqHreHQaY9IPYbr1PwsD1uK74A/NfhbnKt/vXetL8x6
HkomP2FR2gbqbWfGomnEEXt0lwbhirltqF3lAAxMStVvmh3IHSDvOdQWmOJ3h+nSJZUKduwnrY3q
7gJ7ql3gAFiDCLkVfdhVzgBoRMSMkDQ5TaaUFzbTwzbSVFqFw+1VdW+ASl7YG/Kd4ffYG8/QgVCD
04U1OYW+wQxVpnDmofXo8NV7RqCleUezjzPJDMiRgrhFycufnV/55Vbg91tQt9nwwqah3QOMf/uf
ucP2H1edUJ4W11L4tyGG66sw+8wRHYtzV6bFO9RcfxpHsWHMaBMa8oQluiOGOvtrvrfOBZ9hHOjN
LXrNZxLcMheljw8W7nsSc4MSM2vaHQBPM475VM8SGNRafi2oBw7/3pqwZTcGKwykbPw4NKF67f1f
NKXp/kzF/eMHiA+C72CKuOelco/20QCduLb/aOIlTVhHC16xX1V9DFpf2k2y3d97VP+qNaqT+0Oi
2EN83F30quJSjGWXx5WUG3QpgLwjobbRWoqHOVkYE/B2F4u9jk+tWCv1k5XB4VEL651OK1hTNnjB
O5poaYMzWew66W3DQQ3fPsYH1yXmGvIcI4BROBxm1PEX9wUdEW1aGXdNnwwiOv0O2D1Xe+X9jUfE
y/CLGJ40HYcpW4ML0Vg50Saaaqq/xyuSBTRG839nxVbncHr4LJ2jxU9ZZRXXDrCOLt/AJFA43WyT
M5KSuz5EijUy/Qum9kwp7P0cAelhZquyQeHNZvl1ts1Xj8nz+BGiKkgVCxfJAW7QL1Y934GuLS4i
a0EzaJnuuS+aKhkGfMZc2J+vrjgETRsR9Y/sE3d5QBD3tMQ/GEj8mlyo0erS2i/JYhxZ/QvUQIHd
2yAaIN1aP2uifKccWEcv2HiOqmSDl/Gj0Bn3yeLAu9rfM1yA6TsrDjxTjnZW8TlZuOBMq/sBOSqn
dwCRPKv2AWTlGJFHOgIS2WxNgaNw/gurH9p4R4PRN6PtjS+X1hxnGpAKBZ5k1UmffVPT4EHBV1PG
mhjMJgp+QoR73X/R11PW0mqRNe1f+nmRsBy+QaR/s6/jgF5rIcu9UfANAsIjPKBGSm6iOzdRMCsN
a2AT5Bo+73tU+acdSiqdshPl1wlJK91kE3uP8uF/9+WOjnr3maOfGZTZAL7eGxx1bsfiYAeCDfSi
Y58JBwgxhTASZyf5vZEfvuNoTtFoG0Xj7kHJxtMfdCEFN3KLfD90masYWLPsNUHPmaLBWXkpUsAM
GRVKo+gVQLtlLLiy+jE4j0guaDeZaNdZE+CXh0+yCP4YQ79hOQEyU05j8s2gvJVNdsloLGTIfQpE
N0E3zhGpg+8LD83gfMPeADscPfCX8n7W0Zam/w/hzrN5wzAwVhLI+/xJoEgJ2WXM6wRMlF7/RPcB
J64vhPicy9cqy0drz2aOEMbwpxPlphurH4HLV3iy5Cj2y2hZ6SYqA5Pp+iuP4unKQfdhFoZxVzE7
T9uiYYPH440uOPc80ueE0LFTvPCfoacrJ9qUaw12RX4moIiBhXPatI32oLmp2QhGB8mH70rClnxS
zB+gekXsHIgLufjew42HWH1cZy+GLYXxy5cuxacno7T0Bz5fms44lSohAibZEjXuws4QL54LAmmU
oMqbZTDRffF8+r334ZMjbD4OJGjS5aRfg838Z+3TEDs3EsTQFDQX/qQ2VAaoYVKA75TRclSlPcrG
q22zfEOM+wqTjgLfHceRmU3gc+7mGq5mP8npcVsRFLlw2P4GZsyv4C3ejgVEq83mfafciK6vcLci
gllrLha5Z/Tlqc7DOXLsPBcdiCGoV2GkIcFTCyLFNny+JIvN3MRNpCDdiAvcSmJEYc2dk6Tqp9sR
dmmZAXmmpKfJHHIbuI619UjAw3Cn378Kgaf7UT3XdwlFksvPuR3mleTk1bYrOf7LJ1VHAVn2bpYq
B8Y8FGENMz9BIDl9VG/Y0y9OWwja94Wxvr1wH4HwoVMVlRW+jfU/CzaVSAVPE4LNMMIUrnpoqViH
Bb+i6SseZAiJzJSLiXI7wMnDb6bcoFTI1buUBFObUtcwSzR+R/gKnVEKUMaoN7k58Mi0VQCeYK70
iVSQyNziE8HvF/dW6DRyqBUh/9pY7LAlb8/14YshvME7Z9YPUis3HjfxxPEt9q0lA04IWMApI1mx
QXx2eHnsxK48+UMMfOItSh+tGccqBZx9S+1xT63snofmnY1nQjPKGcqewS7ntTxnVOShTSvNvVjU
1ohWE70ENRCROkyIgPPoJe7ypy82pKs0izq+JkD8WZLHLH/6U/PehusLAuC2CRxftdcETeJJ5Pc7
XK6/MVLPPQ0fB0VYePBUYwNEYlxHzFreZJYDdlFxIkAi/TXqywRGV9IiP5KZjswZOuNsRXjAMAxO
jqTxcXgerU8B4SsZpQYxg5N37SbRaCBXFhvFKiJtwGkei8yU57+uxHCTdfCniSRC7+iRy5o5r5Qt
GwIz+fVS5PN9WRgTSVTDfr2OYSbTgm/qNfyJn45FPKZklU6xCtlie+KgS89SHZXokUDAVRH5ZyeK
OSVqzmK6T02hssiat1ip0m8c6iqdHPkDXhWoTs26nUMLD1lGWEke1GvDa7KwpBp+OAAx3OSutOLu
FoTCAsEFvQAUBbKmeKMFF7NNof9lq/O2LUO1KhKDEbj1dmcu8PiWQDPBJ63CAeNnQKoaza6+WcKG
mZ7Qcd2m1sWKV9Qjf/FMXAf0bc7onNX09Vtc+/d5IlszKVdqHKqA5WzxmMCBbpC77F1GZT6XGLDS
o+okpXKaYfiqiMdNhFhfvUbCq2dzNr6Mw3y8OIA2yz+gY8oZGcPD8se3/OEPtOrDa2WjLyzVV3PM
v+GbMB5G+Ex64N1nfgI0Y7AyCyWYzJzWco/FuetLSauugLQY1s9DutOYYL56GQXj1SZfF6lrdgMJ
vmkHhtnvEGzO30je1jUt8ryivQxKxNV92YhnBp643nC5EpYrAMDhWQgnbjDF1YQoIdzU8vO+j+8d
dYJrNTm0tF5etV3YOCZ/XxQAbW6X9f6hLIiKaWtPomOOR7HMantL5m9fpS3Lz5vx0/VyK6MjQ0tu
5YAZGii8pzMF5Osnw1c8N4B2eho5d6xEAlhGn6ukeIsxqbIMmi+J7xxOx2qRJ55Zkjw/O1yZ03b6
pQCOOVcyHc7kfEAJ7Jf+/VVvr9X9wNuIx6zuEYdMlXZrD3U/05q4kN6PXjTSRjQEC2cqwkQnmrBX
gA6LZ/Y0uHpkUrcART0zO7CPL3CQNKl4s1OvX4p3r1KKPguH4WbJeUK57cDuA6p3YDtrVO9Vv1Sk
i8OhStDMk6qSFNqGB6TZBiL4nKGRHVJ2WTd7W9WeJHxMb0dQH9Oi6qfxb4pJiOt6xkUm6Fd8H7ed
OD0UmRfrx9tOdXEBGMD+jd/AVtiUZ4cgo/fNfwfyGzMHzPC2otivo8iNcYMl4CNpwSXhyiKVf/n2
X6m2SZY8QGYbb+vJLrgwopm3Qn2XigpZM68SFHikP2cg5KGMlCSrYT5lbO9PyOiAMNe5+F3p2wwT
W/zYMQvv4rs4Y0hRdB6Gy948OPdSJOHVVsyBYtIAE8gAxlAEf6gwEgYrdsR2fa6W94fvwRqnMZwG
H2/Vso211OoDo4O1OLHRgzJvPO+chLSB9IPzL0LdKLOIve5lI46OX4FIMZexmu6VMxPLY0dCv9aV
oRFQlBGK5Uo6Qwr9ekve5cicZ/36ZvQZrH5e2mbebUdHUaHom+Qg0O4riZ8GTC9qGhzaXm2IsQdx
4PNdbbe+wApPwN1tHN/zV20TampkEkqd9fIFpFTx70KIRwlkqqrgvUl6ATAZfZWBFTkzwD+PHNAM
4zFuoEa6vonALqJEiCAzAthuVP7fsZtNVOYSfEtIU5AMKjmTrrTlY6EzShScu2P0e4KYi1Vv/dCS
9KL1omHFruEoycpnmli0BqIAlh+tyBd/xblbdxlcdmZGVSXOlJcVGFL8vzhl88JuLPz03xwYA7yF
6AWIraScDDUjiFZpyuCz+Qg97fr/OTnJDvIXuIYS3cdcQBBuS46+orXoCCQLlUmpgp9xft2gEhUH
kEquGMQekpcOFLfzWwGbyEjhwXK39WVu+/lJtmj5z1MSN7ZIaw0B29TeKilng84zzH9pwCH8k7c6
YQ5PugFW88+YyX/Wwc66Z/UH2ipzcNJrJHQz26qCFCHo2+sr70UKQU6m62OglK30WBnhNjDHJd68
g8xXyHyQaLwQIsKHHvE/Zruqui9sJidwIWZmvsM48zjwGvU/VLWtjxMQIJhlqRK6uSbV9wVm44BW
njIBshUlxBQGFqcIeI+cdGM7iPVSJDnPWNufGBW3qwCKmb7ifAdFBIbmq0JgvqsC6SwvxVkJ2lLw
aQUUtclTDj+99ZoVIrzdLhxWYzDTq3YBeZg0SXZAjkP/ocPBmeXC2JubaQwORZ4ytpUPIt69hnCG
o9Rhzpdd0IRBokaLFYuLRRBPlcJh4UtHL8BSs7wYKR4YPBRszOzPjQCB4bY1M3IwCalq4SBNtvz0
/l6MyBN16zFZv3+kmG/hcUO4utlDrc84LSOxoVDyWlW3ukrHYsYYAL+kLahTuJmQe/bcin6u1J3F
nvgLUYakxvR71av+3ikdNkG4YzpKhfBkbJvDfgk8CFqmxrco72uR93Zo+8q6AlcppeOX2ZDm2m+H
fFdVYnGzbd5y7zh2+R9RqXjyUwhktcqncvby1bRbXI+y2jnlm6OkTowo2gBlc+1QGbK+zCPdSs2B
IJs2LnChxy0VkMeiSx29Hf3bUz5+OvFwuxfmJuWZGAb9EwHHtrdryRN01u1S3kcFuw089yzaABop
uPVsermJ6mC5cmESq/Dt26dRHZiOeApMGArOZsBca/a2tHwLlAhLJYHKckxdSzeKx/7sIyOMhv1b
K+BkT2T4jIwWMB2WywItxOyJeD+OLjv/o8dcFpa13KDtLNGRu0jMc0Vf+kWqlf/yt4NgnL2+bHP/
A1HTWwQCSwS9m9VOvVp0LYGdcsXLoyKGfXxhtFUHWta+n4Tz6om18TgR2EAIYaHNw/j2XyY2/Bc9
CLDIADfpQFZu+QdsEoyeqhOA/MEsaOAoq2qnoAVdjGou+VGeMAbpOZI20Qdg/q6V3IqzwWfXSaL1
uHSckdEjbV4usdHSA4jwZ1unhy39bO1msAf44HRKP1uqcc59j4tUGCm3/vWA3bmK+FbTBaakktq9
zUbL834nTmeMMxPZAAuWiEpYDaYP9xlz98dvnBpC/Sb8jFu0E6zTzwfZMuWMh5sWEu0llBiz5xTd
o2rn4UV4cgXcCxGkloFnQ8jLFW5U00DtkOJeFbSqJSpP+JQ++e6r2A0KT0Pe7tNgyRQ9T64Sdcy6
XZeFej+WSz356lIjNP7nzSw33lx5/21WSTr4sXyiP2y9V0ZJZ2qvk/4/7f2SXfWjP3SOG3+BtHUm
RQn3khRi5H9sJ/OdWvqGXtkSZaBah5G/KDLMIuCEOO7AYakc32ctS7BJrOUGmb54wAL/BZRtNKlN
MrrF13Ca+ZS6p+tl+7fCKW0pQdjQvMU70cR8OmjuU6h4pa8IpYKACKT42QagXG90K75l/09mIpzU
qQj7Vi3c6ZpTMppxbF+vV3+VbZXyNNjYE9Z+rgwcRFpINkjqlV7PYl/TbKKueIviAdewO7wqA/sB
tSmnYaRbNbFBsnD8iptray0ze8IGeAkquIZ+6KBhLiSu4yiNcVJ0kf63RcfgXvOOvYcFtgbfzxKR
HQJyDT0GOiF3Dr4BK0E1i2ugwohjVu8/edWYCx13JhNH1MzTMpyomUyslLojYHXHimMmWR+qTwcp
NYK/dkQrhF3CC+/g/aCIkUFNVE6ZqBXLhaXm7RMXQpkEFcC6YA6x3VsqnmeDJ1sydNH/FtdUZkyq
LQ4EP0OToy3NIeZlCm67xRw21XOTx0P08ReXIYFRKZDqKwQVaigvty/2liFnje17BigABx3bWX9s
vDkqOdd5/6O59yjlKUoMa8oTdUtG0/+mw7AGBKQNRGbm6HjC/MHcSzdkvU5FP2/q5b8DNN86Yzps
t8FQ726pPVUr2E7oo116zZsslmEfeBl9mpbR6St0wAFx7ML8IX22DYaGWNpCeuqdXQQLQoWzZlCA
4mwvKsM+km6Tk3oaGuuxHHqtx2XXPyl8Wv0oCWDQJdz/PjfZffRXehvrb8uvwyt6P1I+qA4J7L2i
cEPcdqSytix6FQqp7hio3c1HMcc5p4EvhvKq4idYVjMAaxd2k4aimvrDqFG2MOyB4Hu05jw8rJKm
igsfaBw75yxjIJg1RCXrqTcyvX+BOiHghQ68S6lN+v/DQ9EUHdbwxmSeKzxVuf7+k5RVDWL4n4Rx
a4ufHOBJkPiu2zI6lKlnsk6xNZF3ISRoZ3XxCt2feN4KClVkLOcUbDf/djisW8iXDnBZRHFgAd6A
za3MVdCoDyPB8LmWBj4gLg1MIAUcz9nSLDVlZSSDRYa/SrT6UIOk5eFQyZzdFs1dEGA5tfjlKjxK
W6UgDNv0uEF+afinZ+RResW++iuXJKtj+7atBMAZmPe3HvzS6rLg2rFa9e7/9SboLt0CH2SVdIU4
YjJmvjmyHYhHnXeIk1dGqSVcs0zA7l6w76znlezN1DFZWpISIuZbhd4WbUxjo2v3QRiTj82rdylc
xdOA/c8gWCYMn6g11yPU4Ovb4WeIpSq/ubRiWjLCYAlG2YgZNYl8HY/mzXvj4IU7+PXCQkO32fmP
MET8WJfJVu9Sx9CiXXfuyyiorrOKFYMaTFx/1g2tHDwn9XKekrHcFm8Ntb+hF9SFBfn/6WR3UgZz
kHZKdOJDWhqZDSpnn2IKd1wQmajJmiitmwBwKp7nKMuVsmyxDP+DBLLE5t6TLMMPkyUMhOaugzDC
YSGI/ivC/8Bjurin4bIR479ICKU3EXR01O5lVufInF/1L/gbshy/URCuTrTtCj62IQ8UBqwfwjiM
6eNPROyte/BJQvPZ2f+DMZsG35BAapeETgz5OuHJlR2Q46DMCWrYki5EJvMaT1VairPN9E+gY5ls
ci1JSvZ/nivrJmHhQOiFgB8I8ECYmogQWkTkKIy4FHaTYvz4EL9nfwkU0jarBsP5E5bcge/2OUCn
N86cx6ekimvXhBTIUzZE273EgacAVJF/A6lJHiCT0ic7z7En1sulzLDv680F6Bmjz4pe8IWbZb1x
PnIQD8AUcEpKKHrbmVXR7o+43PUiA//Qkow24GI+qAr9W+8yXWIDKtMpcqNrD9LF9O972fntEUVw
VXyG0gEFJ10K6dWHxkIACxtp+l8Q25QHAKaH00Dj4eSNxP8XYZyuh0E3lMleMpa40YLKTc4lbloM
A6zT2c6yHOtOSTAAUYTF4CObTcdOLrNpITVCBnFb5o3EwEPcY9WEDo9950vSNrnQ3i6y2AQ6MRS/
iAV44g7o8ZPf8EtbTLR+E6BWGIPmzxvgPqbZHRG+L+WPnMh1I6997IEx7CzhteEaeD82FvEB/Dt0
iBw4ykyNh0ygDLrnqpaZMaK+yCm8Hi/QHOGhh3zovC0N8OQUNRgDnLheWelCkNF4k0V3twv2K5xx
6TZ6SCsQIfw1K37HtBxShAsE2UjLFm1kAgXK6x8K11/eqykAWL3pD2xq0hsLVLFkD323TvrbK9PR
MBhP2MpNkLZCCX4oQRSO70PLa1Z7VhLk4zuoxizMMzeNmNEUBKOL/2TrJf6ltRLx/eMvQTvz5afZ
6fbzCa77PW9k//5nFWF2d2nDCg2RMmciCbhAnalETIzxllgiwGMVqw/KofsHPvBYZZZI9tTMsqOx
uOfMhOkq/SQHfGSmf2erS6dz+TwMbyrzma0oWlrWMn9SI/vkZ76ThU1jkOgfKQO6MBR6KNbYhUXR
FFysuwb2vO0c4mEcY977nWjwH9DtbmEI3r3M3v2Rqd3Ra7jFQ2iUHIzkav5rDEsWR8aCdmtMBGlb
3eyhiGVpAh1JbPUlKgOyg/DLkpmEWlFmkl/CGlhkxDCfbbzIlMAp/Pv6DTSmVDql7dk4IujZK/Ir
4T3h5oEGkf1v/yhJxg92UAnOaQo0I3PCx2uADCsex2imu/a8eyZoTZzNBYoP462Y3WfzvGtqNnB/
M5yFU0nwEr1HRFNHk8iJus9iAUTNX40oEF1rB9O3I232BQWAvcQ1tiFqvLL0hUBQWw+iTc/Sigpe
V3x0sGgw49DFCjnA9ada+cf7KyVgu2dSk9jALnLYisgNKvHy8QUYfUZPVdXJ8ChXvT7CNK0HJ7VJ
6qXmJOfZLLCzd5q/j5rGKoDS/pbwJyCoEoLoPN0u+Z9y07aJwwKeGDZqLprzndPOMH8/4/QZ3l8b
gUbSo8v2SfBQnLldPK3yVsIGHHikGrrm/Wbgs3MW/qj5z+EO+VcQocawkF7tRBaCTDX1mywf/YYv
pPrf8dxnR6TKtGwlRkej+nYJJeM56mSRiKVlCUEF7LKuu2HV4ustWdCml+dZ0CoK9d+bkUTeueF6
XvMDwKpr1NTfDIt5ecHxLNIFYoRl8FYQbSCmvBmDigaRAq4m2ZwtyCMhI8dxoe4oi50OnwMgC2we
7x2T5kjHTObB1Mutr0WNrSQcvOSHrod3WiLxxN+uOymzRdZGf8KMIkBTC5awlZm9YImC+2RT/7BB
nVILvHrzNi3ts1sK4wxA1fAKPVaxtubAOI7Uw8Jt1ePFVfI8SamJZ3qGTZnXIhrXWSzsJpS1x5NN
eAB/M3F1dl2ERW3pHGK7t2cCokxHNhC43CdlzvSDTNUpc2zJFyBXdVhddRtGFXe+6fGS9ShPjbHs
D19CSnPVkhBKw2K55yro7GgWYrMlL3qsPBL9+Tf3p4VcCmmrUvRy7MRkpSl1scgWOCOYOv3qIrRc
JbkI6xUt1/xba13cdiXiX0dJXlPl8xZK9/22cgnX1kuueALJ4PW9zgwZkOCGm32Wyrkpbmx7oRN7
3qmILFmf3g5xunwzK4RiRatgStLtdm273nkuXMq6QJGXscgipXqRSmGQLozKy+RM6OsP2J1zBRVz
Q5vbUIHjwkpztQIS3twRUTIYvNz531zIV7TLQts29yzJbqVdraAbjGHWaMvilv5FTEi11HYWYvQA
yVVqf0zM+FD+HbovzJwNTs5ZlxjEcCccsAmKg/h41BRdXi/i89NhlJpVnLCUrw5Zz9yomIZ6LB7Y
HC3Pqhomgx3Bp7TfSbCIZrvOpT/2vcsQf2Hci/q7zdViFGsXatv4zOSxwtLc6H2ljAPZPM4aVKSw
bR9NVrcGbBB4TwcZPPkfQHZxQi+2csae/Q2t36WIlOj9C9+bXYO/qDERiB30y+FTv74VPGG6ePnR
zl6D5VUI3dwqYedJn6H73nMsZzUseyaugSl3HkPJVIGvFYzoRRYazfsPilLpg0rU+CdKJ+gWb6rK
h9O4EiT15j/3ZNbu6VRfArvimSGmmC+3goXS4DyakvRYHlS7wWGYB3yom6Fanrsq6Gwha+jnZsRw
NPa2zVxsWkxUCOlcPrOxz/MmjJJhLTe/ljj4J/pxAKKHEtHtzgjbALphS7z83slA9fECOQKJy7h2
xOXNx8u8yoYOGSZ1h/1uxIaG2aX/1PgM4fnv89RNYy0UhqqZ5j3k/ZbVVHvSH3SsRFojubJmZ3wb
cVNFZS0eoFJHvW4b4pqG+aDt1isJq2kwZallVdm8qbXPL1wmKEMAnKp83pdaJstDedihYOAhBph0
pqSbMPyHfd/1a0sUB5VFjp9d+TmLBGxysP2wP8Zs2W8uoM9XzgVKJzXyN1/iUbnITolRLakPNQVN
a5wlPPd9AThZQcJCK/g1I41wh/+kikDiIeom/q8K8Npvj1G6b+52qE493sZzb+fhCMwaYEH31rcr
6YW9G9UPGSYgLl6nd56cbkeyUhteOJiOaCUxBg0EwgL48hwKS+iIZo48shjoboypvk4I1JHoplz/
CbAuxy9G/Nb15nA1GNd0Qtoeiiq2bISAE4mKqbATXAa0qcYIXHcFMIOP+JAuUga6BsndsKuSuj9f
BMHsTKQIBMGsDN0qe4Dr9YvoHcZzrA/l2U6V9cWoMcLAfD9B5lwhQ28MSf4ghcYWVfd6WEzlzu4t
5b2XckUg8rtW9y8caSrKBqVdIB4oYYZM69NIRhCq3mZySXrDRetPQMoLY5li9sVPDi3AJI6f89vf
QjTOynNX8d7qQs2bd/WEODMu1hee85x4G2mkxecgQIedEBp7AogPdDRgrqb8LJpnLWoveCglXHxL
a1+jlZKvp/SJVjw1e2tHMoftB/BIx+qDcrQJqzWqOLGJORBA6X6MMnFChMkmwIYFA8FbdFHh9szw
7CvdryCK/eDy1nfq9yILYPzEisLbHvjqVag4IDmCc/vkCl2YdgUAeDkqr9SQrhWPZCy3UtMpA8wB
tmPNoMeTEhj5eagB/0O9N+HphU3wRM3FN7R0VL983xaNySYHazhiIO/3x8eaPDy8Qi6hM6dH9IEi
vF4QFEHT2Qw/HpAM5Ru+E8QUQ6wOKKPwfMRSEdlWJa2qVvl+g0tC1l9Q4nIbblLyjubboRMb3aKS
ha9+NOtBjOXhMMKe1aNozx/ynQBfpj3rXa0jMmkBBEF3iIqyZ1/qnN+y1iKdDuzRVJ+SbA0tD9bv
pg+Nmpzr1Wi6KKxFdrCI4WqggmL9W2fbGAkq8gMbjTitmIEZr3dZKo9h5Wkm3RF7+oIiQCgOl2kL
ghmXarXSC6288MK9CImiH//W8vEhT3NqJJ0kwbPuzCMkho3SVe+SmZeI8y4QtmLyi02e+GiuthvU
oW5+zaPDLr11HVJJpejnCJHKosPG5eFhMYDMJFPOGVcod3JhCQWf0NdmyWNtJBo/HAtrtjtsYYh/
WxE1BdiSwuwwDxWTbCCl3NsUmPBOdRtpIWh0HUzm0o1rmAL6ujlmvot/ZpTHmuPrX10EUO3a+nx0
9B0bLGo7B8vNHhjaAaowLUGYUMlWoH/wjNqAVi342EjdtZjDUUdzengbViKuro/KuW1X2CzcW38X
Z7A/YMTpkt8CKJiyOhfFXgDnYFQUrWkTrqgd57C7sQDUY+5UPTE1xM5yHyvGye68Ggj1aGvQ4Vrj
yfJYgrub5CARUyuXH2puufGrhRY3zf3Eyz1ftRVSweKWU3ej9ydoU5Og2MozYoYRQRTQzX5IuEIT
LAF7fzmXmZcyHaJ0Z6nicyoOzR7S3m/mtpoTB6j3LjC2dW8W3fIhgEUbCuzdPvHNu3ExzYjB0CkQ
k6uRz6bsoNFLTE7XylmJvRv0nPAEJFghQXDVe2ie0IOCm073Kr12JPkJqET7Oy9RJRBYFJ5mRt6U
iMRqUZXR8fqH4hXjuemxZO4lT5Ar7fHyj2dbR+8mkwr2v99rtYkm3buCoGp9PfEsavLgxny/1kzc
ntFPk5h0IoR4GQ7AixOXD8RXicKh8v/MFINWRcoZPc4DLts9yWkqQk+4aNc4GYO0/kxjdW83gZbQ
NGoZO9CQF+InfikafwfTuOPqMlTSQbbd4BHFsQyTPczXLZ7x76GgpK37C8eclBCE9dccFHgI8qFO
cYPWwXJEnu2jmR4A+Wp4TffWObJsXJcaalm67v5jzj7AkgDUI0jNCkHEEB2HDFfQQUfRwiz6IzhH
wnCFpj7cO2+WGkUp26rBvDLb74B5sn6wnfIucr5AciM6X1GOXBNQUcDzWhtpZxYoxZRaqfDvFAdH
lov614gN5fmUHw81AbUdOwn45O4FI8J3mMiQMOt9tFS/s4mKqUUXAuJfUugGCFJsmjs20Xt0/UDW
7Ds/wTJjkpmAPGvZ76cS7KtjA3oIa2gvIVyuOeibPwdCuv7mmPwC1HOPaWEGFjPSkoU+nnrKktge
h6fnnBPyD4f5Nk3f1E0mkE4N1LbMuOVuU9r0NZEaE1PAet1cBwkpCodlTX5VP7kiYQaT4rnIohNv
SDW11m89WYCzsMPY21ZAAoOTXJFH27CvVX3qwLbo1sq8DNCK4734B9o/3U2Armh4hrujSrgtCzbx
qdqpYGVQvYZqY2iLlcqfuitpatLkKcAH/FpiozqA1j6d7852FL074wAqyZRagj5ewK9rfqbe25LN
9OQ20EAOcEEfU/iD/Y83I0QSKNrA8J3eTVfSjoX5QkxWvutcxeEnO5Gz0zlwTl4x1Gh2wMmcc4Me
Ih7kL243td0PBgIUp8tqholOzV3hBcAKmIJJ1x5BImHdI8I5yvokvhdWm1PNGpRctgWmfsOChZ76
BOWT9w4s4GIsUqJNWEydT9aX2y+kTeGQjAQJWnQMEeUu+Sjais5lg5f6JfyoLm3a3ilxjKTzpk4V
x/OtHcKzIZtSC5F4+ccIIVunAjDmZENqFj/5syYPtKoiYdbvobMg4d0TVk6NQOSN92i0btebn6uk
yVgcFbNs61+ZGcUr53Z+o1KSCtbxpOg23ERDe4wuibD5Ide5h9Jk7dCnNoHHqpCTc0OX2uFwojg1
nJGva+xQEpctEgQnPpTZmm+Xo0U5KTNu0taOKMU/OxHmZNJ6Qvd4/lQROIAzXiVxUvwTpF/XGIV9
50rx7c39cigA9Xl03unSSqYLBE/ErEeRZFVjAUhEXqXwCH5aOA64nl0KL4z9/uMFaRQTdPdLrl5m
wNRiWFwf/E62crshNdpMdKgxlcvEu9IwUuOizc/sTFmz1BOU8gC+HxxszlG/o8CNDMtKRufSgk3n
KobdyFrKJ/rZ7GUkhuJMi0S2cQ+ZBJxEXZ2Yj5jHnCPENla9QxcgxPJDmQhAwdN5gjic6dwV5nit
n6NnKoT+95wvBwN/y0A4VL/KbVgfJUW6oOiscnAcT2fInkCFGIGvVX8nZiArUn9ooO2ot9CTIOiS
gwuSv3ISLyiwUcMQulW8voneWmeFuxZ25CDol3NRwwI5/gitZrCv91Hifrt+3cASsbi96nSvzGqW
3O1aFVch7bliQUbGjD+AfIG/sJ7tlK+x7agR39qPHAnI2T+SDN9CZ+KSXmCMVV19GatO4wA4VCAi
b2JrHZp48V/hm+umqrSFa5Ef/RLBPZc6Vhlly8Rc0Z7XR5SqQQZPPwa1xELSLp9Nhc2zZqoQfqXR
7ZxRJk2oAuJMB9ws7q75IYpIwOnCcAm7p1angUGwlfEM2UhQEJ++pD4xTZDYZV/Tn7CT1wP8X2d6
Dn/6H1/Iki+FqGSKHAGAzDGMwSB7MwoaRq+D6hOB0D1S7QQK4qmlMR7XyNOS1vpkohxIz7C9zQLF
vGywjTNpjkKlayrbjFl/jDGFB3XjpLuYE8gSlhqVoMCkCRTjoTmzMTjEKYILV1UkiyClrR0SzdXb
UzsNObNMrIOoZwHRnqxXW5B35Cqj5SM4gObPnAYC9NAfzGNuSenoGYjU6dZ9Zo6rYYYRB7K/gUHm
5T296QUGQeSeorCdqPmf9uxMoQTjze/RgM/OW4M7eVzNIuAitcYz48aaaKSpc6Jcfai4MMpyWYjw
gi1K7hpt/ZFmc78KLF7L9+VCqY41ANM5ZYd3nqdhlPkA7P2xm9BatWI9V9VSE/wRKWCYebPEXJs6
oE8sqtIw1iGbdnfOPIP6HBYoz1X+/mddaKK62YTISgTcRVeb4H/VzUsAwOnPEEn141icgdNJk2sj
5SIdtO6scFZ3a+VHcyn25ejT1+QZmKFOs8Dc3DhJDQl2IFNzNLXRlOe5r61l5r864VzjMcAfVAkr
qsV5xrDNDpG66gAlxe0RmLRNLaIoARyjUDCoYzB1x10AsIposlwmZm4LOhftwKlJHEcgpTZFS8fp
d2zKEttkqRQL49MndH/4Si1MZQYqQkL+5Ubs5vZLp9HZk9CFLoyYzGx6MVyf/D6z/FZdBjoTEZQb
Ca2Mi1pQ9U/ov/VOtbKO6MHCHWCNjQJftq6zp1MsbCEDtby95mZtdzkj1L5gv3g9LhWQMhg6C8+R
XBq+7P8tP6fRkVyMVBju+H23Pl3hMU8mxC3AGfCq9jaU0lwvw1K5CMonr2W2AHdhZxPS+H8u3Rj4
BWu7UftwLY64qRMSFSr3S6AWupW7sWOpYT8R/af9HMB7Ue4CK6kt9IwwcgD5H4CNNm+fZWZkX4G9
QQjwZWWIHiGQTeFYJHSWtW5yC2NqiuEtH1nSSsssezHYcm906dZm9igD80mJl+cRaQIqIV6ZKwbZ
gl6PCKv1Gm4BnTNug0YUlHEjidoL7byyaRyRl9vA+nRtB09fVIv+5uxQK0GTws56tHiFz30g2Qlo
gYSyDqC+8zEXZXtPtWJ/aNhx0573ths1LwQzXBuWamMpxfeg/UKtSM0qYwn0tMp1pG6Az7wHogY/
88BWveWAkucc4wtoS3fxK3pG9/UZIBIJdPhoTw1TH5HbAu83naO+VMTO8E74BREVczMpLqGK0Shg
eRhokVi7Xo/xkJC+NE+tn9rqCamVQd6MeHR5CyPHuZxFFiO8Gi1pkYcd9yXehcOVkiphKWQy7gpr
03dsBGbraZd8M9igP5vynfZhlQYeXxUrU7hG5585LPFN4yddSnHoCIDL0zDBEkqG37ArUgIQj3gZ
EvZq8i6DDycTFjUR9HsYPw+VG2WwL6xnGyfIPeH7I/1WN6qbdN4KpYvsb2EpX1weIOWSBI8f/Lr6
xO6L2RZwo8MfOkTCfPeEia2akqclpZGIkbNS30OHBXdIp+TtSijIe3XrtnnaN/ZiO3x7PSenRdfu
7mq8wFOHe0lDakbIs92dzlSALH6bIXzIonKFvMlAlHYdQF9+ngH+nxCE2oDrZvtIC+S9tlASlie+
TcKfcLqZcsLdwW8DsziIXCh9eEBtJ6Opfk7KMddonnGH51B9Pf3PPYdFNq/yKSsslqDGf29MsdHs
xPGxX+6EqzY1HagA/K1GHmEp9NSucdzQCU+2udpVQSF1J1bdMZvthPTf/ezVLd7T5LF43NaTd3R2
PvpAWhuMmzp2qZ+EUHFldsXHFb8ToiSHWWqYerQvYOKFwWu6tJEHL7B3/ZqP1B/3y13zpO4J+PTm
ts514WXC6yC6ruPd15O/oOwN+YVoy9Kj3OcDHYEr8axFupAy1UwisqFCdG0ewZhmkITBnXxroqKA
x4fgyAMWw6m4gFeCy5nTHyFPjPDd3F3pBvoovorPoHYPomv7VFQg7981Fr5SMRBEuyHwuSytWJFT
CPQ9CH7OBAZPLys8XSgwpTVOjWyVJ4fvMLEDbk/PjndBUT63Hxp+ECkWb81TzQa2qUR14hnlC9fa
iu35B5pfEprvG96ZilEDvneiRaYEIdd5xRomYp60rX/g5+uy9REyADkIR+KjNiuEna0R5NnX7wyz
rbOqvRzjWY1l3U8UIMBr6kHRDI5lkBKaKL9uWeMyVlDVuSZmkrxib/OQulLXWxhq2/X+2NqTWmfL
oQZ5/IA+/7F2bzz1gUEJt3UcdQvsSoXYuh2jWqgBzUp8Ily54SLBrD0G0kX0yNK5FN3cITnaNEO8
4zyFtveWLYs3A28PB3VM2cbMpCKij/CbVsjJn3WLg944ccP765ejuc/EN4NtPTidZDhk9rTePEab
oWGl95D7jcnJ5hW1rU++XCNvyzArcUVBCmcXZbnyC7H8zOp+HosTMKDn0oiIZN8xM31eZ057HZuz
OqYH5+L6Ni2cPWVIAm8YW+qVN3Cs64PzcpK4lwAKW6ruugz7POTOrnx6zHOeiLhoRTImQjRQM1bN
m0fwQgD/1fn1kaHG8kPqhhjgyzMXAyvnJMRblHv3KNZbm55psprhT2UEfHyWq3UJgOPs6Xm8Mjgk
o/825/hXJF2pWPPdhgj6+vdtDCzLj6n2dCgF4oXEUjrvCxFI+aY5A9SetKVucGG//UkArHp3hf1N
ifdGFUGQRK8qoYNRJIaBiN+3wlsF0MgvXHnSRHifcm2XChKq1bk1OvVcKHOb1bIa1l6uhqNFXX2j
+dbosJohux3ChQv8dJWlrNyUJPV/ujhsJIIduRfjfbHxB34AtYbDwHo4JKJO0KCeT0AIdbbaTwHc
7rDdZBD5vsX5osNLv3tM9dtnH45TeMz1bXG8O58yg6pWE0XRjChdvx/aIJmqSqOcPwiEJH4HOXus
2JFCp4ex5pOWdZSGB9z/FZVxpmgLfyzD9Nsz1WIvXtPgCUaKfEW8laIWjbZdfmhwwFMBOqYI3tmB
vKEY99Oh+bS7c/1Zv2hlVl2pF5klA0lAfUegsyAHBm3NgSxvJCqVqglEJBc6ZhhAu+zUilEvDfHH
6pOD7wOnjyDfJ5Ese+al+WSfOPgxYGENhH2/4Bwwyhnl4niFWqpRTT03KWWbREDBO4a6RpLITgC7
JL7gNJT8pMR5UzbJ1LaWzNF5NLtyHltAr9UmJ53F5dBKt0+X2HfKj5BdCjFEt5eCzDYkNlfSMTld
rrVasCZ+8kbzg8sZoh6lCz1yzzNeiMDqrQr1UKnB5rfoO1hV/KTO0R1p59pdaIOcPxdIIU8kM9p1
WdZ1X8R/1/bQWQhAOn1xM2vs6kkvaT7X2ZGfLOJ1YVFPO8iKeaPx7EZKnum74//tNwT6xukjrod8
1BWAALvi4ndk6WxZmB25jpIkELU4/1erCDdSCFgiEqFrBmHdh7WfXuYdvygqoWFqNFxLz4GbfHoq
wrdcJ8mqjb1gL6v5AyOtnrFUoL6eN2KmLmox16wB1wJOusCYdS3X5ca9iYq53+sjrEqjXu/EYcFk
/waXSNvR1u1iAWJ8sI2lN/aLsM29WOmLOITBjpexiOr00l8T6YruZmW4YggnJt4hDHoy3GIupFb6
B8DznamhLiPQRmLXr0jYIJmK5X1K1uM52a6HrDrY/x4C7OTaoIpWvB3iiaxABDawqIMH/SjAhfa2
j+IF1UsVyDapfB5JevFudIzKvk9zaFdXMzP21p3rSqYtQATwd/0smFZXkLzABJ1lgohQIu8aeD6f
NTZeC2zumZcn93/GLNXa3vtqtke+Udk4e0mU6L5gaPjbZxhqPRzv4iNaKEqSqIWIY4ViYZRzk8y0
U6v/MnBA45BDwVn/qtzZUIi8HxKn+4G3/XlhZNHmgAwbIxLPlNOllEm5RIEvxjn3Px0IJlnZjTJ6
CEM1m/mbDm6jp5n+uGHoQi7emi4vhZAL1gJTH9SRRfkw7kYcD93tn5T4URbKYK4frEQXbRN90cIW
KBJjj9qRE6Gk9imGEuQCgg9QzPpJiPl/+rDqrl7U7mRo/dK/uOcrTa62ZOjOq8WOQDzIyBhkZzap
2z3VlpAiFe8uPQvwpDqywUG0uakf+JVhxvU+vq7xOOJyNhRSEjxh0LmhhWu1uwZ9Ae64djufLBEl
LMKmz6TbH5Bv7l7vjrVl01AMbH+NK7iZ4OAQbYwom73ZcraHbdZPl4xPAESnLY/xjWXeutwmgrEI
UTbYzKFV/HFb6uWVFlUo/8yX24Xni8kbz64R/Shx1mRYGi3YO0RGp9jGWFrtl9+IzPHBtY2Oz4P0
3/r2KKQjh2bymfVOGa9rSDUuC8CzFR8+X57UdOYAnTu3Oaf5Ia+j1lbRcHmP6bcp5ITyniKzwXCv
fOOrf2+RmbPqGLebXysBteAQhngcsajsVlImFMs+41Nt56drBjgdmlr6GuWbFUnonO16608atS/V
C5dWJ2lotCCUQZ/PIBTxyjGuqlUSslAIRS2QAwdCT0oRg5m62TAmIZS3AbPb4DgIUlJppFZTUF4i
Xe8Ah4hJ0zUE1MDffSwUbuwDc5q4PuAE/Cb2M00hU/7TUG3+cfkbbZIaoWFUOsJhgfk7ptlo2Imj
x4wRuC1aUj5Fe/f/vYug8FQpthHXMW1n4lIBJSR461fynEdkChXyJaEKivpbNqM35tMXpTpMnmcW
h76HiibxE/1p/h6n6gxvkFBqjTasCKTRb6gXsHLQ+mi/IY9J0Z5zXE75pUhLYtkwIlOqGbTcpoPR
E9ywnkdnHwD7uYmdSEfwCL6eRGyeSyB2M1pnv9GUcF9lzKlVJqQ6kJmpz8FjGhtZZwCfj2CsrE0W
At8e8zpG0s7KbUfr43QH8vqichztOzBWxQ1l81exd/WJAnvhbKmjApxFG73TkO9bCziiE6RNW/8f
HvopL3qUtwplK8eZ/GtmKiqpye/N+PUSTGbve8gXHVGL3j/DSLhXbqppCNOKRljEl9XDRkw5SFPr
PYB9iLOllkTznGAzYArTWpC1LG1sg9HXUAu5+1S54sHHbkE1wkgTtNdBCpdSeUBNegR5VCCqS5Zd
69LcGuAn0NobkSq4o/stwohb3J+zWSjvlMenqr0inqCQgbwEu+C9hOgY3ZSxtqmAYitJycxlJBDr
CHi+/M2MH66XzPlW2OnZtIVQDMBhqC86HeyzKLzlxow+YoKUzlXI64qqLH6eexXzdscX9FjqblkG
mboyoXYIpk1Nmc5WTVh6qEgMpiOMO7QktZ+ZqJIN03Za8XayXfQNOBQeakQ6ubsk6EzoojKiqGuX
guDmFUeQdC1K1qH8POShSU5bnfbVhEXIYERRUNTAcSMvCqL99Y2B52/JgMKG2D0roPEEUfn8t0TZ
NavTp62EYfYA6zBiktM8LPM5DzrqimaL6BCJMhzGqUoiS9AiknI7diha8Zq4nXDj+CqKTOVj1PrC
JsTsn+3oIdryMT66oceeUHvwCmjriOPaBart2K4nQMqVcR1rlOp2RhzxDMEmrz1ISiQDDxL3tPmi
YxSISzMmY0tuZGmgCTXhl8A5DvJMN91VbKTF7UnMvXy/vHz+UT52KXAC+9lCxUtI3sE0UO2T2y+o
lNs3t4estF9VaMQsS9qbyZvyW41dAviusFrFwgXp/S/aUKa4Tfqherq6r95FZx5c2ODeCDIOrMUD
Ggu1eXpo7Unt+yTf5j1yZ4aUoJZfsI/u1T3xuK/hv3LwAvTvjfBRJcPLnbdo9mPKf05GjLELx/nj
jLhmveAR3k3uiwuhrS4XHnrAQCVFYkNh17DJlC+LS6Qe24kT1Pnc7MwAArUNxZAwnV7z6aqW0kex
Hq1Oh4e7cRM9xiSGT0aMBSIEtFJETBAlruHcGkXuh0eI3szcv0/SSr/5M+9ZEPH0Uy74RiMZ2uO3
hmTctK4n1ni6Rwz9PYF7QAHD70UUBcVc8VItnN19tT8e9zyNA/fmWSReSkZ6NwVV2mQew4xcaeJZ
rkoTeZv3S7LTRHrJ+xURcIQ4Ku3KUrBBoUTbTvb/T4bjvfRS6qnlPvOU3nEkkWUhBG+tItNh3AAy
7jMLeTv/GJUq+owqhcaFbXn7HikCTYlE77Y1QQucISJQond6SZ0VyLFUFEeFl51PNAXofFlMKxJD
nICn4oie8X01LgVzufiymlDpU9g855lJ7Izdc4HYt1ryh6y+uWp3CqLCcvDcD9Tzbx/QUa31TWhW
Bk8czs3nOCBqyZxzMyLOi78YJbsrQAkuIxykWmIvurs7wPtXgOGqRPAiPiD0rw/DH5dYLS8IyheX
Ux2aVbxlfQqw4buN2fIiylAJnvZwA0p3pIi+hOC8/LPWybPkuqQ5XOcufDTEDz4h99blSAy70YYX
A7rF0Vwh8x5HdfbjjZkuMcFYwai5L5rkdwx66QrCMJ3jvqinPg7OF6w3VUgnGCNmPhIMVjgS+YMP
otgy0qhikm6CR79+oYthl31uLnmc3Mbgm6T7rkG7V6QGCv9y1NHo3jgi1StMh3BecfsejQBTgKSf
GhavOtUH1Qx3qLLdU/FqHxSLjkW0/p3sXAuPP+6H2maL3mdbf1rGhg1pEZelIyvorKpYMZbJEfLG
Asu2ZucmVcf5bT7yN3YfbDCzo0N2bFYFbQzvzfTcflSJCmrzfkPvOdnzUa6eOgqoNiRVoGRUoeN1
oorQyaVxq9U8V7855nnE7O+aOt2I0MmqTo4x5nRN/zQ8kvnYiGjSbQXCxUCOOTt9YIL0q8db/Smz
qsmRdrq0DL33nyoov016Pr/H9Spy63zi2xXW12Outp/cnZnLYXWQZH9uac0+SFKt1eEY0mb/DbTt
RzMaDQNwIBsqro7hYrhJRTvoG+EWJhojhA0/2xRB2szQb6Z8BoJitKAi5Qi4T6JH0Ek9w4386IDV
kbkqiKpWBhewTyKDUvgvqDsrGsdIlD16UX/ieG73dHfQH9/KFjNgk7e/XgzjQeC2qBnCE8pCtD5O
5eRuM9ZpJ18/6bQuJyRfW0gf+ecZ7FIKXL8p6jrDY4WT+jscGl4A2VBdcw+eyQIubxObcob4lzdi
RlbNuJ9uZKN0KX6Fs8uIsN0Wh4njyG1VsyvoYBRCIgbsimHQ5+WjEjceHXlGTiegXxvrT3ZxQ7gH
DVbaS6tRmO3Ee7BaIUdfvtf/n8R3uK5QeYtC2Jgf5xFAJxpn0GYgCNYIFQXjEv6jJad3T11Dwk4w
48E5iZhqJkS5LqdddrxPRc6v85z36aLvnbSAVJBFFYriNc9oades+OSiKgUNQmHjJkK1RWVGMBWW
18uzDhlis+M9Hw9+GJ92o+0/Bf2IM4biELNDhEFUF2VT3UFpRWphU675BvRymqAWlh6ryR2q/uxW
P6rdelMeZNIORry4WSV4wqNSZsSmiKfYEUJ9Q75HvP1QntjmikrVUO1Z5TCbEDKevBQULNiWeBws
n17dUuw67AhqDFTfHqdG5Y9Uox20kilB6hx91VaE4sZH//OMtnhGhEYC0y9oeJ0paFQY5MxUBG8c
JGrq21BAp1J4ku8f0q4uk5yB86t6aqSC9ja8CMQlC2TvXi3u1VHhVNcbyp3T//7wBhkRu+rPkucd
v+cS13/sqJDRCqQQGwDj/0WRWk/PE6q8sRJpmyKBjsTCq10wfgsfAvS5mlinYj7V0HHAoSdyQIPz
s8U9vcIGlQcCcKz6uOA2UbrWKjD/grMkvPZjFgUjbbICT6RmMRbUDcG1uNc7PKpe8hCWlACkY3Is
K1+eCaewklQCQtmCwJyvR/+bqnm7QxUXNYz05fSBVFscgty8yAYldL7YmfzCo3kpK+b1uYIu2FFU
Bz6ogmyYRYRVmKhkFJoMwLoeM5WTG2TH0c7dop74CbKpxLDTjOAn7Vg1RtMwfhNOqtD0mfoHpuZU
7Lo8V+ZEgVRULgpSmYNyNNFxDhbLredJ3PL8hplqg4eNmNMwoJSmDffLziXeeqoLl0YuNLI/iXwi
htKkeEIpyAYwwwcadH1MuTKTkPnqnEBJaIGAVCk8xNz0OajW6jR1urKYAMzXK6IFWP+YqdLrsttk
0i6+wDsKcgiAxJCkKPEir+sA/pe5FLnBJn/B2XgCh0w1LcRBgjkJClq2KT22sJqd5+CjwDQLRWTP
7X/cmwtW16Z+aMJmGkCLgckfiCwiVrLGNQBX05z9ZAn/BuMzMd3GAdNkQaH7FZNw3MjFm8sAbVBj
fwln0LjZ11eKq89Tb7ykrHl649h1s/RrOo/wFI+aBS6qwIIT9XINXc7QbIxCgkf+8BVVUFZ37Y8Q
0rBNwyrtUWAaw9fXgiPyYr39eoo0ziPOxqCc8YsnaT+q/BATXLxHSbO/ElHoGsnBgkY6uLrsi+Xr
1NoyzKBvc+Tur/nQ+QCoy5rZ3VOMfaP/M+lZoyHH48mmNntIZdGfL6dHXIPWsJFPMZ54EzKpSp/G
j45H1RQl41p8uUVXUynrxt1IPrvo01Y6fV59yxD09pADTGxgeU0thmXcFbQFg/ah4QFxf8ASh75o
YCVailnEcYnCJOJGkgloD82fginKfQ5EeXR3RpotjfhuLs6CuKCzjBisYCqlVJ/sVliqM+UKrxdd
5a8n7b/4ZaGOXXFVTCFsV/vQ+mC2EX7zpBhQO3Xwe+CbQrIps6a6joKJ0hmb8LM1StsvX8saGzPZ
4XA1zhhjzskCLJRdcSIrDZ2RS9UZbaGzaNis0BALTK1gPJGiOxLWRprGXy6UDgSZIIpDAUUoJj9x
DTuPOHJ0wxIfCClELwoTuyC/uETqbmvCs70G53YxwUp+yYnm3khRC5+NtyprlB8bP1zS1oVgcCBS
XoE+b5P8DfC3c87fou9Ovf84QVTbkDMUGRwGY2ffk3KCE+/IpW6BMKwVJ+Kj3KKLCqvqMVybT90m
4Lvmu6ndDb9tRuXlxt7kVRizUEzaO3nVF9lh0ycnGhHAbc358OdvUFlXQdz9t1MFd3Ft19wHCktx
Fe8kwP6P9xblAq/aSox5K8eFBD2mBDVSwVkmw8jLgEyKu5zIDksskhJrvdAs+5svZiEt4z6pG+7t
ZSOPnR36UFG6K/Jnih6dTfzgsKtaBQe1DqQfLaElX0R4OEJXPGICA1AhXQEjXLIil8KSy15p+ltA
20Bgck5YjRciOAANw720948m6rJMSmzANK595VRAzgG6Z2oE+ScG5JwQqL7bedoa62aXJ9r6tMUh
ZSQfzfVFY1oeNtuLpBKgzhaudNa9rmKpwbGxEhfclAL1NRwhnVv8JVusSRfpSIBvCcGddAmRYSgV
lUvI6bnOUd4kAimo/QmPZqYO7pHMc7tDcT7fZAeG5o+kSalk1qxU/ETifw8yGD023qoFTA54u4bj
dDhtRgx0L3AeSery5myhV6XJFVKvg+p+SH2g+QkM8v2paISoVjRdnfZrl7bhAzIiezOQbNwXaKD5
Id7YuT/K/Vp4hOF6YC13xIpFP0+IavoFdtCtnjjJ8FI/pMvY69xFeHZjwVE5jeixqUB3rpnmLoUC
7cnraHf+pDp9OkKvNHTWVgFnig0mdV2WqAQC4P3mEsLv292LvMB065Ve4Z3bn+4SO1kweZGmwj6a
W60tGfGI8qlUsX6sA2vu5L/OWCNAzCFXDQKEnAroobqFVQEpUMGKan32N0kiM8je3e6pKlKWVJmL
v0cQkS7veLyPGRke7PoOENK/sT/og4dwmPwVz1rnNj+R5JafuzfRXNTiFKUBVGjzakuxEJVOIF5A
rjn26Ll/K6684EO8zDXHo6Rdp1FFrIVDuXAJkOkt3jXj7kgbcgyB31YOwUDSVCFaD8DMtAI9mHnG
TjEM63PD05j5HIgK0pw9VpX6fUGGNTOb1rAhLNcKHtoXjtHy53si84u6tKeLptSoMEPRMsKbqENk
0J7diFREGEtzFzJ4lWq8npYqyeODKJApeMv33Bsua82GYCLV+CzIaGbkU0uHvcQHaZgBhWYCRZda
G+EgVGHPiLGz3iAgeFB3G5uCap5bNooTc6WazKzjovP9BDiW60ov2DimYIjMi/is/34j6U5nwXCB
JJLTDsNDECCBtd/hKPYCFEHmljpHNcjP0SreNTz+TxUVUQeNME2GW76yeFPhLHSnQhhwmxVzODIy
t8IyWmayxaKIejlneSLTvaY34tytvbHjtYDxlxgEeA23MqdUSzIu/Slc52d8kbGCc8/dBiH/iK9F
d29Cy3LbjKaWYRBaxOj5KEO88ZR/YEs7lJL8r2rI7Jp/q461vsw8jN6+nV5EsRzlts+1/tsc2Vrz
IArbm1fGtUymvBpKb6s0ug+XDf2sN4vZyNH9WU4JGkWNPE7nHOlrJPUr0tWUv+t7H77GeyUJK9RH
Ggl6uxgt2CoEskFVD960jgC2HGoYJfDHRmAn2cSYeNZUsUdaYWU8CtAo0KECbVcuZjEXJ+pW2L6E
xGkFbheBMuv85P9NnDgAj1K5Odr9qPTXs0oeLS8JTHLO5+s7whPA6P7g3Q/ZYInbNgAsk/ScKuhJ
V8ZcQchnU11RVaPDLAR1aCaqWkfkRa0yDozQDmLiD+Q0foD94ymHy67ZuXvRGU4I2Ntkkcuqw0oW
6rYNOJSSpTqWD6jIeeNDz89aM+QMNhdu+njImR4OtFw8a8ckekhiajokmhYuC6G2i7XJX8O2WNpt
qvC09cOf4J3ovDpp1KvLtNtMu31AE50jodOW8w0JNWpRrinU14BLZVtTpnZrrPAuR19elzSQbAcK
OhQw6yHc9/0VbECfPA//BWoZuOXat0y5Vh6xgl5RGRXGszQ3WMQwOlY/W/DmRf9HlKyYco/ajQ+1
XhGhLF1+alGcB7yduINIHXL00MFbO9ijqdc1YRMlTizjt4tmYxwSm1KjKDi8caIKgbP41p8vKlF3
H0hxeY8O71wSPLOrdsyh9rTVQf3SzItrIpTPOsoFF3D4QnQImIXsOtu9DptIhCDafttMY8U3OTvE
u20d/7c4PiuUW7dpOXRJj6i6TZH8z6lN0gVcusp4Phmb/+7xFjyZc7ZR6Xzd7KX2TrDf/9L8L8sS
Ig+w8TJ2kbJIgPPYPgJFwNCyCQD70WHtTe/HaL9HWBWz5HBGHdccViVDWdK2b8SHFELWHf+BZO23
27g1N7HeeV2mTopAl3f08psQTJT6TtpLLvZ0FvONfqsQ3RYt+TNJBYcioWUdiMYeHf1YOi4mJxAD
cLcJ0/7npX/lhOFvniouabli8wuc/QcZpZTYc6tn3iCSA+ZBnWqj4xcMHvN6JC2Ct1Fi4TWLr6Fp
qyZuDWL76KzNAoJWFpBjzXYZjwlLa2nPMER1H0br7MvM1m2LCHnK8oRIcEXT6rjqT8aqckhha5S3
Ys3A5P4fo4Ap7jn+G3MRB/7JzhcpsJdS5Hqp+ERrRqFyKBlAwHWKSb+UQrk3jAs6jrzYrf1O6weJ
Si9Aezhg1qQv4KKzCOk7FW3NjRnmjHDEa7wcq910sLgc+u1tIAOCllvmLqoT7TV2mG5GhDpxWRMR
4rkD67MOuIX1RgwqEKA1aeQiIi/fmczI6Ytn09TvxveoKIVgT7soMBqiG9m/ezO7TiCV+zETWnOI
2WPD8xj+KOCLS3EcfZCKOyy8WuIB5D6dJB13STfw5Lj46cIRVEr2Xr6NokS5tPE72mBD/GMYQFMO
Czg4CWwbPFW2CAcYdItEqzBGjTFZMoRUZfhJVXe/UuFTbp0AS3p86YeSxlMrtD7GoB0Evs1NYj6f
asly19ebFJ19aSqorH4ywN04A5TAm5OAXYW9H/YpchZy08npbM42Iz8EAEbji0XE7Zl4W5M5+XvA
oLEqGVOltvrOeciGpPWH7HWQu72gKffa0HCq/WSqyyEA4ZWUBEHqPd+5EWLTw0RrHgl68/9YNRYU
UgLy8s1jB/CCWThvQYyih+rb2qy7mCm15vtF0JVaAA1SHE1Axj77+Yi1oV/10fH1kLbTn2/Bs7om
G5hDpZSgcuEm1L8EDsQlXVi9hnxd/FKB9n71EnbjFZNGNbvL3QFFvm59Hx4VA5f64d/NjMm2qyr7
B4PrrIgcaQoW6s4x1ldZ2M046l01QREdRHiTOZ4bcluhi+rcmvuqwGEr+HAEcjyoqjjwnST7KBoR
HUlurYVVoa652dQeaaXWDf9n9xaSz8MO/M2EKRjVDiAxGJ7D8uYBDhvU1Wvamyru+df7EDZ1QAFN
qn9TWofeqSZ3shT2T24VUte5MdBJAQSJ1D8GR8rwD2A6HQuMAvAZIaKA/45k376BjmLrYAdFuDs1
QaxA0xQ/8mNCOMnKwmF2AbCrUw2rl2ZRfm1WePaF13+mh2KeR78evfTpCDZz5h7PqKPAPDNftQYG
TqDZJqOfo7PG1JCea0NXB1JEAXXh0d1k7yCBV0P46j02yw/VUUXPeANkBnzgBq8ic6jiQkAgn2XL
Lw73tabR1fOSefBNYayXaWoLrFM2vCGJbkEMlcOQ4cYcAisAXshtKzr5rLQF+3S71cL0wAV9r0nM
5U0YTMxa0of22wBra+6Y4n/XgYSsxPnSWleK77683yskKVT08JwflW9t+lJVXr4v9W3xE4PwALIj
Mhu5xeihPYYrfQDfiC0v2Iq7hsHQu3EyZlvJx3jYzpEtmz+DxkwXSfWHcytSC8vVdTnK6Yeao8KH
C1tEdtPPNc03lLMTzJVVilVb8nidq0GMwbl/KSIeg4OmvnT0JnmDoYkfbefVBJbRJDVWDW71brOg
1YIewCViMRuWDsjW8ImbOMzJ7H2xgYGtaXZ2Y/aZeq4xiCYwhn8wSZZ56uQzs0JUfrVj2QK6RsQk
ojkB6ehJuPX/sVbPEun4IBMQCtZJ0R6ghdqTtSnKBSqY/LwXjApnDKnn4yZDL22luocPe7oT1yE0
V1hOE0Sf42/JVZitMSclx8QAz8tvSV12FoCWCaSiNuK5P8ycAb6hdr5fke5i9sI4bADpG9Yxte+1
Q4UqCyulzJt+PkO3GqV2oKE9iBMF15gVmZpbmMPsUVDn5tGJ4rVpLKDpm9RkLGClF7ZsShZiGkEN
aLb76WAia4GqwO0ocy/mcfIzqlIUAlXRhDxnHUatj01AdfNwNk30WL/Un9bY71TULFUQFhtFch6l
65VcJR2mWbBNNyP1atm9r03Wqxh1yXAb+nl2RFvAoDuFGxnr2J3k5f0y+iLIXOBJh8h0Y7fR1dtS
NG4sca8j4QlEtsoMxGJToWHLxPOmgiSKD9TgAQEn3+KM5w/7K4YUFIVN0cf9pp1OAD9Y1Ih9/trY
jzqUcDraRBaT7kBPI5Wn7Mn77Q1pQbIcy0nl5rtPLJbDisykOvd0HSRpG0XekYhMy4eEVmB7OrBU
hSTrSLBhY4TlJJE5t32I95QN1P4+cgYB4ECSk9pT61I2wte0EByurQGdth0Osw3wi/3iAAWOBNdS
1RCID+XH0MGhOI2RRkgmydS5Et+ikMxI8MNgb4IbR76pjR6+nchEPJHl0CCztjQVeQ9fUi216mEM
DFYmuEDDvjle7NvcMFcooqv+KMNttFRFlhd+mOXEjMJJ4dRYTx3a4qMHJpg3nCwDhsOsPz+z/eOV
3/jyZ9eaw0vdmCLirj6EBfR6HL8m0p9/lP3IUS+g0hVzvCnJgptZCj4KsKR/UE4LZfbJ7hShMsMP
9/Xb6TZOFBncSkR3VRknXy1HqQ+9secrtkEXSftY356l8qltIA14yQp6eNWyM/ahGCeJMQwzDuYD
+uRo+5mc1gr1z7xezaiDpu3g5twI1VLXlYSLKNQuzfc78JmS03MsptK/Xoci7WnVOjbQrzY1iGoF
kf0eB+QbXiQEt3rMRieQ7rtbie//YgA09cBk+gstiyDAE7npyffJW2s+zx3B9dpVbzB82fwolEdT
i5ykbhJ9HvyOc8cd5JJIaAZqZEcncY/QFb202u/pDteuBV+Vdrlp+/8TKPl9ZB3YI8JcJZFf32DC
YL3Qosqv1U6EAabglfuoIPjSBbNP5jAWBqHH9ynk2DhhAUqQ4Fe9c9gjH/tVntWvA3FqZh0jCEjQ
8o+vL6AUDkY/KkKN8CQDSu7MXMUz2l9lKbpQv3kaL51ErU2/XJ8fPj8dpYZgLwPHyweaNL9afya/
mkAZWUrbGJEp52hSJwnDcYkynA8YNBIsihjo2nIrnQ3N4fMy6xYm7jkGbc+sm7chmZScyQ/ZzpDH
r/ZbtEyo+52TGZGn/SZxpii6hcV+vOQ6p6xb/E4qSeQloJYHBeCP3YOeyx9OcH5uWgSubeFRwxPs
k8QRV45BIvVX+ea1AklFXMvk/rXQ0LFm0bNYXptAgzTKEbJLDGPMpKbd3W5TnG1gz45a5CJxk6Ca
un8KZdLAvKIDYU2aWKIHVbfdDm2EO8DrhXqR4jUf1KyL/LC1f09whDrLEacHWoXUNlI8F+E99D/r
NkbEQom5Gx9s0mPkQv305P+hDQKMKtK2eYPeL95w6ZLziw9/NtSAYXr7yoXj1Fv4VPQ6h1QHwZoa
A+W/JN7Yl0IktuOK5ueG60G+mB8Oh34ZknyCKu/YkJkUt2ImzuJ2bx0cfzwsgTYOzaVljCBFPFNU
0iTVlCSmkFWEnveSZNVqVdsiOdNO24ZWhFX5ZqouHxxWkd3IuG3NSCNE+r+aMCOaOppNyi9sEnWU
ofRHcO/HIct1YgjfSoqphC0vnwmS8kdgBkomkIfDfWgWktTsw2IsiGVBodqtiztYecpTw06ifyjI
U1dvQqP/6rUsTKA6vyGOvqu/M8WUQzp0DuyxGsckjRIRrgZEdIJGvBD8yzW278XlKGmIOJ0sB/4d
0QFSm40CCiSFzLsRo5OcDWzj8/FdC6kKhJLx/DHS+M7b8mxSpF9O2ivA+YZaXJRE/pz8OJHRkyxF
M7U4NhLKglhGPxkORxY3A5jsbeY6dQhGk+gP0AkV2osmtJf5pRKDaVnx0F+/mhE7YerrYdnhJUlW
TKB+i8O1/Mxk+TIqT3B0uSELszgqt6iTleCX9H0KTEqeehwgsIyV2nJsI3j+XGxSYsywo7qnC6L1
vGEzHubDn33rJSqaQlu2btnHiokG1c/mIkKwVgGQwP2n59bzTSS3DvezC+AkSY86A5guHYOtruJq
OwFogBtQ9Ntu3IbRw8NH4mac8wSfBX2LLP9RcXWIuSbTFiPhYMahTkMXrzYvjkkKeLS0yyLpRKFx
CUZhD5osRjyBcWjrP4n2NWiw96AKwNc7rqs63VVkZU7msrMIKGZHHGd0kuT/YOIZ8AkkqCU/Snw1
UMkLTG8arkvoPvtQZ+f1LiPQFALIN2Rh669FWXlxMr6z+9cTqVjwnqG2qLzoipEb7HGS5IaMOiLQ
splOHQHZ32p03lWoy/7bO/JLfzZ+9k+GWvw6iYKL7mQE8MMrKvLHQIUj4sr2exnC9PbqEJR3dPVd
EbCAQOo6oy5umzn9gSn5B4g8V7FN3Ej1grzA9TYiWG9EgpoosHTuVjCzq8MXAfLcXv4CDHjnErTm
mPTgjjqRlqZFmSSMYrnYLx3n4pf3yyjRY+QSXtX926qw97shdn5abK+VKVZhgQZR/VmoeFGJ0vWi
S+rwfwf1O5ihEs3dPO/e5tfO63kTyMlCVVKgu9IQPiXQg7xDKAWry7h8ovl4qZOGoCIbt/Too+Fd
qSPmjQfr1OmlhPLsGARmu1qzOr0P8WJjN0bbJ/yH2b6BLwH0tXtp4S0O2RB0wfQbhyyJecGq+O/W
wchHMmmVJTrZwmXFzHv10olzhK7PFqUzHwnpVdMIzPG42/qDVCQKQ03IA2U/VNqrXOW42dWF8ziA
knxnjGL+/xNdaPZrkDCPmc4eEksE1Axy8rYeyJD6uyBAQ/TObj+2lTKn+J+pifempabuonk3kzs+
C2o21e/+BFuY2W1fPE8Tk1OLe8Dpdq3LbSCDHkSarIc6LzSaccqbf2xPzVJ1WGoI0zmMHu4zCUDo
H4fvKxz+wxS/DM4Nc6yCvAnQqpQOR6cdnUhdl3CEd5gNoXX/Ow0jc4JL1kUr9fWu5BgNpOGgKIaT
A1wBGnRpUJzVWzN1W/vkUg7Ul+S2ajWQyYll2RRM677iYWuiG5OXa4JvctnNvuFa0eDF5i56hJc7
uW2npblFPls/GBx+xYjI/BU1qv1b1PIaENacXZieP8sMSqCIwfWol5jO4aW0BhFi1/wvd6FCHCML
j6gGY05BF6QBnfs33PQnZx8kMG1ooxF3uoUkOsEVVwSGkVz81hbr3aJrMFuvToU/4drYyjCq4MSA
nZYwIfzUW8irFY2/V267cSnEava5Ezn44+56A19oAkerE0755/1Pc4tHIw2no92of6MEdQcSxGGC
oTNwWey0gpPpL9sg2OsFEMkVSFQULl/3DvkjBUcQiHfVG20ZDLSb6qgWH0yskPoYA3ZfoCei+Cde
k8q97HeSUk9V1fIWm2qrpPgcDRnpHOcPMc0ILcG0l2BKMMaYn+IqB65b/Fr99nlRjxFE1y2PtW1N
YDH9rgIjVBj+Fi7T8UdUs3ypKgua3S4fvf51HmAJihXvooIbVZVfJVtJ1NaVEpNm+TsHAsXjFDNw
1J7qDJ4QGBVWsIE4HwLFglFLegPXRyZXXITorLGnect8eODATJyg+FasAj4T4A1/sQKcOp7S8AKn
GMBWmOPsz2c9y/+vZIXkd7D9x1zKBui4xqY+NtZTbZ7bJyocHPjjZDdk03f7+ncKjU3aUJhRvr4q
RGCx6LSziJuueAD0ppHr4/+mW0UFMCA3QtZZcHRhf39z2sgw0rBptIbu/Dmd8W+ey68417BRLc2l
33TYxEUVI6t4xXm76GFl72MONTlqcpZ30JUd6yK3JtPte2GpRpanFQ3EuC+4WTSiU9a/CVgqwng+
xe4DfWfShijWH7IvlecKhDT2fbJdWQwiJWphVMIvyqJ7+liaar+Dt0KaN6PuAzAytqUDW9nmzrnT
z9MkeJOqUAl6qrqvu4KNmYahkhxC6jmzLismm442vH12kdDhUnZq0CmMMyzotvGkhelyIGhDzcv/
TxfgYQwFaGrFNEb7y1BfXitpuj08S7iAQTbhSVvM/4W0UXMckqb/Xh51QYoNDAqIDE+ns13sOF/7
OFYuUuDV4w7rvTmQ4UwpTlSxZgrq6LRVzot9KEpIO14CmyKaI+DERQw4nM8EphEfkGFx8nnQL67l
x+l/PDcWpjnsnHTC1qppgrkItN248QPzzlvdhN5m09BcKD2dTYRe+1w/c6IPPOOztRb3WF43vU2x
gHZ4o3PEs0LDHEXWT/05CdZa+6zCkMm1gDRXZ48QzNHTwRhVlctF7Z43neDZIrOXoBedZBP7lsII
ncSvO19cny30HPaZjfIBk94Px6xNQD1RR1NxRltS9W97lng0OxSj4Hdtd5lLzWu+cwxqJuCxofmI
VrNmpC+GJ9litiC7exlFb57sg+FDddabsH2MXk0b+G8CnFCZl9WgKIKPb7XQUNvVKhosC5NnqjOQ
JmJL/eJSq+wMYpIyiZFcFxmVBCS4OMogG9DSkPa55kidHN8eQnYBKI6kr7tslZjKZ5TedtXf3s1d
rb585x9PoSoYTKyGIw05cNLZIOyNUAdAdoenTu34RcauAj/t4oCn3ouybzByVlAtxz77PYOcRRZl
YfybfwSSsq9Edsdw6Cwq7/gRLK79NbVti/OYVgYbYRs8cTVPoxLAZdP2Mq4HGfFtGEMWqwFRmJgM
u/QkV/tTKhamzFiNKDC1CcIPAeZG63nyUMhsDbSYMSl4ppvm1sdkbL3EPZmUrvF2Smaw7GmdTps6
cj8dbj4t6e68gl5NN7yRohJ8kTdLilebDh3I6n4Uv/2fgZZVEeL3/94FFUOjULQNrFzXF2qq7ABD
PEAdgVhc6/PL7cK7Vjdo4zx+l+GJFcJn81xZYGddat0Zt3Kv8EtLh3KZfWbFOXJT/QgsyRF11xXX
WGom4kbj9kaMpHx51eO4uiBZpmGpI8IAEjdOTuRchw65H2V0OncE0ZWc5TqLpag2UXSb+TU7LEAJ
rsaP+QnD+1FPP0ld970riNnQkF2vwHYvdmGtoVKwR8jK8wksKRc/yVJq9qX35jDIgUZHNCEYk0WC
pUnP0QNBabHAiFQsU+NjHBxx8sl0bAsJQKL92MY70UaQ7X6UnmJU+hMjjORovBHkfvYKX/0wpOYp
EKBFDrpRWcBeroaJXGarRqqHp51f9QS/R/DwqJo4wQorKwm8+AqkhcYoviA6+eI9H3aV71gGE2NR
pOCwU9PfIt0zyRSf0FsJqhu1h+mxq/GAP9cazj/fnFMVvt5NheANw6WKEKidWw5ex17fj5kBp9wC
ulraCH0l3EwhNDUb1zRwYW9VGC/qSv+qn2J8LZAOeIRjEkHUvbR3BHAQuZpU3ZU58TSxxrjApnYl
GwYt1v+u8R2lYiTSx8T0zzCR51ebEJhD7UrJnhi9+C3nSUy6IxxDsAagap6LsNBNS0r9sqzy2fCG
pHqrztAdSiZJhTLUj6k7gpy1e1M2HpOTrNSpQtJqh3O0uN/bPqTrNRZ438tpNe3Jz2bAjxXh2N2p
ptr3V0GLi6EPcs0fhFqxrSPzEofeIe6dkqhH/DuFZs5ki5SfchcN3iHX85UnfkzBOCVMVIjXF/gE
NA224WLXBpBSKP9qIKa3p2GWVDeBXVUMysLXGF3iHDZB1lKyDSPBy6AUV24hA3M4SOWjE+oIn5N1
HPToBLmhEJhTLJfVweCJGxGoylDtxKFMoKbA6fYCjG3PegHX925JXMLb2D268ToHP/C7rqLpOF5w
xx5y4ixF3OSwu+tPLa4sS7Zf1iU4TgwoFK4kmp3gQFt0x59b5p1JxlJQHs9uRqIM2aYHQCMqg9/0
c5l7qQ34J0QcFhbaf5XTaHMdXUw7RhZV9wuZ4iUJzU4CtZDDbBaV2hMn7gjt/ByRYy9EbjGytrT/
6MltMs0M+JOyZb//kW8wRI/C61C5FSoqeg/ugsUR+RS3SDUbU45CbgBhvpy022nO0Xk04LwRzwqc
kdrqlJgpZhCOvPfsPdLeo+XQ6FgMe9qouwQVOGOvnhYQTm0QWzNcLwVlWkHZA2ls/v+wfmlUD5p4
jKV/XrUMsG3bNXJuepUGlsJXEPsNqdSLXeKlBtHVPc6jrybxfDfI9pW9bBqp0quJ72V3EaJ7EcEj
isbqCa/rCM/wqRv1F+lnrOJkwj3WnDMbyFEc1jtNZMLlgqpkLNo3IjWdLZVK0G26hB0zuLCDm0II
IRMyZ/BRm3fsEPlwMaIW4SksHFsXA+F8/u/niTITAfozFrJbUQVCX66+lgx/qdoXpOGX7p5yO5W7
3ZRfDakb8fJb11bzu2ObHPxqOzqN9PMquRciUW/feTU/8JTNa/nAWdA1OZA7EwSlWZRHWi7jDOI5
u3Pr2EOnyW+0gJPy5i3h3GEeKV/LOWh3ZlYV2w979vix/SyMm8gHxJS60s0itzNZypfuiQFxbJYi
8Jwwdvke/WCa1zNu/uN2WXLmTLjdXtA3/L4S2rUcUvN71UobKOletPLoowi4h/3WzSI+/Ifs5kii
DONRi4qrTo0Upp5MP4JakkfoRm4xX2el14GM4zPTKQ7b9c9SNnB7tQ8gpy2BGMvSQAfGFNkgsMv4
4ghMFd8YXwAnIvcyKF4+egzvNrQgCNG24YnsHcK6jx89052kv65OehithRXex1FbLBkZP/vh9MHd
dTDbhPDyX4FNdVDxGTQk4z6ihW7lH3CETNKKwudEdiQhpNnwFI7lHpDFea27fDCXY7FsuI6jY5MW
6GT18iNdwz7FJValcURQ6A8BIn7IecfS7vFw0NnaNW4UPPpaK64llxiNarWd6On2RgyDntbJ1l1t
8drvzlWsFonXRuteGwPZYtC/ZdjujC1jqp5gXhlcwUbGspqa9nlZaFd33YiJK+bLA1fKlWQ4NbQN
651NQZID8G7Vg0s+4GNMUFOc+lfzBx9q3vMjpO3gjx0uwwp0HhVjOdTDY4MEq4DTeIgYDmQuQWSu
oovHrUuqMPffQ60viOrE5IxpYk/Fh6w/LUI1tSEyLWXU0F+f2hDTNsykDA2n97lZsIRTYzg2lJPU
MEz4HoOzdtIHLE6PWH+mGplYpnlS+Mib85Wmb0sY1KbhynNEukrHhJ/Gorj0WGB3M7GEa+H2fdIZ
RkByyjRTvDJe5cHSJ/rdBFX2C2dIEGYF+lw6nz5ponshHE+hBoiqlcEg5DgBv3mrOFpVvARvwN6b
LEEWNsUZG1zOUVaJID/Vnaz4egVEihJEfBMxYJ2p311VNqdMY9kJfNJvA3Yh5+f0sHTroEZM6QQh
sXyWg4yFNHsZy/5i1U9gyNtb7VV65QQj3BLlODKy3LvgQMIn9/uV93Y67kqY4Z4dqw3jr9EwE4jS
BR3+s1QtTG48nwdQay4JNsDJyfNDK7NgTXrsA/b1ZZeLqPLnbxbWRDIdFWierBWstsS+SMMlnc7O
/to0mnS9VpS47dyYuMew2MFIJ27TbXofFDbjAmhArxVfwt6FyzO309qLo8C0V+MVVlRmtSx6Q36o
r37vOp5kUTz/Gg164p6r/Z648DcRmYktTCxxrQ8Pk18MrfAdj6yJC7ytXrqDSpKgkK3E2N+28A98
z+1w7xFMLHdPSDdIyn8uDBLQVz9SEPw3qBgwnxiuw1KDl6/wBSL4OEeUSiv5l5Q3shlcY85thpvT
P/SL12+ikxiuT5ZlZk1x9Ce7sMSk6iGDNmULO/rN4qv7yon3NuTdr3oZ1/kLvOA0bIykIEA+fIYa
WItcx6lSwaiA2Pr6d2VOtF4lEBZirPEasjKEr2lDV5VJP19XFXQUcgNcgK2n9qPsGQKv0/Elog7t
mZJk7Jq2rjuVZc5N7qVlAsj5FHk1VogKt/03wLhlHNnoQ5uavx9dxr1Psx2w4/2cFZLxlivA/JeE
oF/h4xZj0fqdiAbLraK1A/I0a9CqkL5m99IjfF/qhQVzJ671tpVBPxrK6m2h7SttlfngjS04QOMa
pxkIYOOmAtNOK+ez8sYDnPfhEUSzdvIxGSAF+qW1HHZIRIQantqq2mlSnz7uQXt0gDh/yzIiwWjw
ddttPmajDnfpTL8oBCco2uGGFDE1fVnPxraGjbpoBv958lTyhDIJXJMO3R9wa2ClugthI0rgSWYj
OckpHnVDsrRJZWlMwVdeFeRc7at4dPziay9l49EvZIL+6J/HdJVLfY1LTyI6sLxpZdmsNmwJ9Nnu
i26X1k7VCq7Ii4eLB14n4yGzttqAbJG/TO3FuUudjy5aT4s/K9FujJi0EW5/3RO3SlON0gQi0iST
TZjyZJ82IZts6D6C7eV9qsPhFbA3tgLAQyklvElS676tIUFlhGyVkfp1gy6uRXvNj71s8jlQMVKF
SFM9qZmXsjwFQw8BBzGBkWnctla00HF5zRop/4Z7/05BS8A4bo1dK0MqwB0RfWhQ2UHkFNywTEN/
/v7+RVC2oHd0Pq9V6NSPxSU8TWesVqCvcoXyLGQKJByFJvlZHlgYfvdmPGUUzYiNlb4zLqReOKg4
uSUJJ1nZgFz+AcoG6iRPzqIxnt8wFwstXoMovE0IKwUICrkXu8RwYeYgEs7hDL7J2ZxVT+teiOqP
iSIPR6feR+0vQa4B1msy7I8H/SaPa6n6iWrYTgx8KvYkPmKunaO0EAXSa2eDcshwWpH2qj7vBDnU
6z9uUKbrsmzEsuIcbEgrbdyTIdtnOlxpj6b+8qli6JtxlDx9qQoAIsdt+QKc6Iq1P/VaGP5wmlmf
/nmNQLQSq66eTW+cZ3zDqw2NGCJDkOuqg8AuGB6fcnYfumaDB4170PrQ+2K4mo9r6dqMGFKe36Gx
RW1qtG4a38KoI0mAHdsHaNDtv+1RHA8QxCzEl4dtKGcL9NY1bB4Vhw9UWQre7pExXJF+w+Bj/gF/
l0tApZt+LLPfPBPINQQRk9HGgtfL272Q0+u7WsPPVA9MJrLhfEGmsMnGKKSdjXMOH7+cYIPba9Ok
D3Z3KpO2VL5+fhByTQHl+QXfJaoPjDgJJuMgvOuWiTkM41wJ5V86ZDP+N+oL+rKfWVrpzg0I2SYm
zSiO69HMBSUk14QqlnXAVVYLjLBvh3zgX0Pv6DrJ5X5Ubdf6T20Nydx4W98kd8VBSTLbEOHtSt+p
I4MC96/ZrQZtxuwZjRi0Tg47+3RgcnZZvVQs+fZf7EAgb90xV41N17aIa0l5+OVxT6D0aGwzVClB
GUhzPUPXGOJ5HmwtySHrDAAMmnYmZShBv/l25/3nb6jn+it5/1ENTkD5PMaC2YulkqDOXmnlm5HS
CB6kXNYYycE2dqW/jyskz3eGKRd+tQeHzx0GAqgOEfd3QOcx/sTpD3jh63cSuEtD5ROFvIUFVWQh
MuYbvLhWizzi+3s8M3rHQsF5lq2fQLh9HyT4DOZDXoMjqJeQrBzsiQOL2puxUjHm7vdyE6pKnpYE
5woWC0jrOLNDE/pPFqf/G+YaXJkQAEJL4J4jzM+krrDPNWTKQpkU8T8nYAOpFOfKOB2OA6eHrb46
BUKADEtBkmwdctT4tteTNRqbhXvQX/7DwBniS36lkr0M+M69hQeTq90gT68Lni0Ur70JJqqIwG7v
6ETmYxI9iSWVDKvNU/JNI5H5wbDI0VF5MkSzG8KQyGmbTXENWgW5Ey5vSEmGpm9SldTiCj2wOzJV
2NfzLhJDm76Up/yEpnrAfCmulm5zBnXOMQpj7b5Se0XFHvl/b85x8amdyS5WShf8Y5XdYZj/KKuy
BhqW+B4tQjnaGc15WO/yO27lruNqgOLeykRygJvVDWEriW5eqC9f6T+zf6djYJO8IBoL+V7xL+Fn
qYPAitvIkx3BAUrBAAshVXi6b34KAIRF8VQxJLpdgq0zG7X0TYG0ufsjdfUl5mSto1xXv3awj/wJ
BwIiD9yw0xdd6EkjXSRqLmiGpllUMHkSkHCZlwcF1W9PovPx5znV8lfAbdmDZDQFTDmx4Rh+GlSv
pswPffHYCMJ7iT41OzoPtUzlwcgSMFYgdOrUCN6RxVX3hcuiNwU+ySzJz8oAo9MYvHhSQ6VUfOfW
Db5a6aKxPYtkOnRKRqZN5My0fvFkcsekgRFZJDvE+Vs17BQZRKeUXnDC87w91cgPatZrAPdvQtAf
0TcTKN1v0OpzIi+sNXoFk+HFrKEo8wrVoLgzn5on7GTR12EJxgSI28Sd+oXcILsarwFMSQBaOsyG
48QkUGab/q0ANh0E3LtzfLvxT7jTNypCTA5tLCEzNujcLr7syzknFmmrex6TRTEcATq/F9Z7I+p4
Rpm7C3puDj22cja6pSW92qN3q4OkkiZ9RamNjkMhzD76qsbPQp53/USF82n/jhzvrQylW+oYg41+
N4trx5c0H6hL+PJJAlSPnwa1/vjAgkaicWBeimIRhrgPO1nHKhnwoDM7oO4lbIlY9WfERKaAl4T3
RwI7AZoL1tJx9aK4dcdknv4JOiJvv2QUosh3A7K8xKWveZ7G/1VChLMFqIk57+D5WEwxG1sIGVJS
ax6FCWhY2tE9GJRh7b6zF8Br99HpmabZqbF/I9Bs+pmUZmvNrSdSB1bPOPEcI7EN7Qy7RXGYiC+y
QE7WOMGBDoFbGB023XQo9NQQOajYQVAnnV3p9xzeQ5OLjyy6RUR7afSpLrLy8yawaNjM+d8k8iqp
srA5e4dCJiq4OCdJ/43PPK5+vuOJGm3gttYN4QHV9UbnaqWi3LBB6h29sY9UtlJJnE3uXOoNMRri
4TMF1edp675KNk7kA3o/Xb3XkRX8nFc0i2QcgmuOzYfFXO3xv5mPuXOHt5eguUZJY5QEIbtYn4IB
s+18JW4+IpZOGli5g5z7Q/F8lDU7bhKoregQdnr3VZ8hnHI3OV7OtvQ+V5FzYfjXyiccWoN5u/M7
WiD+A1g5SvF9CMiQW28eXNa5znfz4uUsIHX7r/wgJy4QLXlE+GAxQpoVx8mbbNxHf0F5MN09/Qv/
EBSjAHg4G/czf2piLrLV0QZumG/PxwDCFkkCiu4bFPZP8h84dt/cB2MzaAN/lLMWyC87tlXWwulZ
KXreLSRxmnPWRUsVxPwEJDUVW6RCCr5C1NvCIMHiKdUnDMqu7apQ4eIPDl2SJgUs/x6fed4ePIum
i1glENhEaWy3DwuQMZvv7UHw5ukUPjKkhsm61JaMurQ8uf+HmXFmBJDuSupOT6tkSC/OyBaRMda4
qKmL6U+NSKF2TKkVrDB3HRr44vpy3D5+2nsA/3BVZJ8ZVSEKpcIBH0YbWKTcLmA786KcQfljLgff
Sh8Sv4wmZF70wpzDzaxNVnnS95cKldvKZpfPbAMVNNdx8B99ucgqqg4oIduqzONjYSL1dxbZl15u
MIbmBBIben43WkrimhO5rXN32euoEqc0f4NOgQfOqD3CVA2k3rLLilfFJpLq/PzSQftzJx2jQxcu
QdC3QCFbi1gF1HO3naUA5tD6lpWYpRul07crFsKQ1VgcggJnGQi7tAd+vY4A9+eKrfp4YtCdQziF
10xMrDaHc9B83IvLKugpcOlrLPoy2A9u3f+PWhmMDM5ti9m3xxbcJmLv+f19QNazB+7rpnGXsHI4
/zXa/f0lnBKN7JfrexjXMFIN9Eh2vg8fEY8Arw+sa+ncUw49AjEMLTrMCbyZFuf7TyUc+kROTMyQ
SKKgccE6eDLD6uMSO87/pMignD0nJ55gaUITF4Euln+qEMeC/wRYeWr4eVr1Q49oUUIFI+12SUEO
oeqFv22WEpXnpGWgMev0oqGN8SPPR8uWWAENiPbt8xzWxRyFJAj2GNeX/d4wq15/o+5QH0x5Jpfi
SmDHZWQWlAuKMJFi+xFkuthxuiYA8ayjGMbnm9lflzr/vrCP1WUc6SXuLhgRdMVrH9qdq9sHd48X
j/R+oG2ywFsNmNAeNGMPW4DQH7JEOfYrECpIIk77HgtgBZ+5QY/ZhtlC1nz4vqEgIqxkOn+uPgsZ
NUTshr0oJUpwcDqVwW/FiXbu9hU6qBROZQFFIkA5BIPOvJA/USM/R0SILEg9AroWBj9IHkMOYi5/
SkjPQwR/K6fpD/3b6KA5bxPuX2TsyJGlYbMo0TVVbLRLE0ONTlCDmonGhZUqSd+pbgLjQy3/uaCL
zb8qsB94xeAs1g6lpdfbkOCS2ml6l4ZrJDVS7zktfoFxMOV+4o0MqdjNw4atg5fPHKRPmBzbzQIF
fzh8jPvqH0Y2jYvMYLyIwk8PT0rlTuARljO91apbTY2eyMqgHi7sFP8LYqWo/w7l+IQRkNlZtgxI
R0dMwrT+4X4qGZx2KS8TyDYPv84Cg0LzNbeOyEVpNRcqQWhWPnxSBSVX0tNswx2QOL/Fq5nyaB/h
f7qF8LiJ5Wct3IqRlZPqex+P4qCobuPfDwzbPiyXDO7xiGndHifwpa0m0N0ZPijJq/c7MPLvy4aP
QCcD89v6C10xjyl25lVMGcjw9BnfBLWj+tvQb//NCrvwNtGplGipUZVMm3kFSYDxqLaY+ABVWB6w
UXB7EezTKvTR5evulV/PQMxJM8CrWSn5loMsz9C292cem/YY0ngMYW3bEOELXeFO6jIzg1MMbmR+
vm9ALIY+EcqeGz6QO8/J1Se9ZmIHXnF55/2/cdQgyd0hCcBo8KhQHaTRgv0PES3h5I3f+hVfdt01
UuOIXReuXiosn3hBAZDTzm2UE7Pbokh4RdUNIf2gPzBRh/Ypc0pZ4/PCBNXLidt1QetvQ2FH5Qqn
wNiKuJu2oTLGhJOuqk5OP07kd542gioxyUrnhNn/QXHQMf46nk9jdcVQrXQKDWeEOcN2cEdLjt+1
s23hgtr62nDaxsUO4IeAetr9Om3SGCNQoIOWmASaQ9jEYMlWq11kDX0hYiFhLrvZQRxTnsMN8Dud
l3vXRkcryy2VCeU4Iqq/sfpsEKQG5nczEuY0E+HXe8q/FxKhtNe8STGIHcrlrxTM7ADXFZgMcV10
REJ4HoxRhlm8ObDWP6ZU5w+ea0E0U/QhWxZLC2RbaPyzgOSZdDjs58OimluIGLuYH1oCDXudE+U3
9pR/wa8HT0NRlZmHzERyqMRBKVpPnqwNO8OlU3tyHx0kkVJFvhZAHJtxEMM26MSP5Og6GAQd7hvj
F59B6psDLDCJEjEf6MqC2lLgpwOm8MWjYVJqTTRIg78+5DOWqtyFnf+d6tAIl4HpFG+EU/dVYe09
xmSeR35Yrpn7gT8yqUEWBczhozPDhPoX+fvSBNay9zCvAK2diXIju8ACR1qNFQanhqSzCmtOTlpn
2R1ENWKmpUFYC1AcrY2BwbzkGUxq4Em8ojk4ipeLtQeDRUATrsD8ymcjT8KrTmdlzhvTs4XDzLwK
u/2TqioyOKz/Wa5sFUVxBLrNKiCv5Cc6IwoCmUC1LEcSZDuUvVb3pGmik1h0SKCiOEuEC6eNcaVJ
FzaPuIcAP0CXwp+0eNejSzMclADHd4PfTsjk0/pVY4YHRDnCqMB7uH3gBuNMAwh846lWULw2RM38
pUIWoVN9EEwAgiC2Th77J8ecADMWP7XNnERPlv64YTzac91OAEPWhYA8kzssnjLDja5ZlwHWyKh3
w4XK0NnUSWcrcrVgMAm2NJTLnPHmGXDG+wWuct+1ppR0aHApHf2zAVr7KuCQ31g+4IDwdPvZ2EAJ
pVC+Ktv/eJB2AVcI/L8jsyfYydKuuWQwfyUDUREIL2iRyOQJ3Gejg4q2a9ZvZkngkkdANcbp1AhT
GN1bZ7L2aHuiC5CKGaz2hT0rBVvRaa29uPxRESci0HrLnCffTd/ZsivlyWFBo5+IiH/6kRSq7Vvt
q4GrSWUDyoPs1r2aHczss61EFPhTcP/8ebWKwrDUyFXjZpgHVKsFmhEZgz+3lMyRaPbRANpig+d4
oK9dTzfYw+uQkqL/JNGMyS9WNfm+1/SZBrRodZDtqxZoX9LEWtBNCl+fKSAdiT/qDdfkPh9vOqx0
HRR5SY9s+CZvkdYcsugevRZVf/0Q5rEvldiyW5djLIzskoTDYkCLe4ZxVKlALA1bHGk8agmqNbQJ
88GQCKMn4vv4R+wOg3/sJ07A+8z4sFcuz3OzgCSNbbji5Hy3b/69CQZ7x5El5ni2x1AraES8dDQj
yOwLDtj9xNB5+68NCAtXOTFEE86Cv3WN5myafqqk9PJJ4uSETftoYNjOZBbGb0oRiPi8YwQ+H7XT
DhZI07tN6ZH5DToS1CkCByxXaWWqs/QFXKBN8Y/QCe8nnJZ4WNWRT8EhNsHrTmHWJ+lrx1qOwxYL
4ISLZPbNIfcrk0rBhxKT00wjBHfTMlRy+7EL9CCt2l496D2jcm8c1mXDXfx0x/FX7/gVjpRrbavR
f4DGVSt5dr58cbxCo3rt1Y92dlzre8fvVizwHvVcjVG8u9t+JzmJv3nkHG9kymxcE3xLHuXzIsgJ
WGi/l1ZW+EWZE5vLfcmQp5BcBlI4DG5/V4/QjmlX4oWEetP/wcTW8gPXSSW77ndz2opp53lDc9es
/sdDFJBJtiVhWyxPThdDzwszeL354Bt6MTPzVm92p3l8Iz1n1VjtMtQOJl4O88gXXEBRteWpwPnk
OFRabsD45pTdv6ZfjXSARll6SMZNIWU/M2qXgRiWePATJT6QcuX2gb0Rt6RCCLOtYKLrjbRoBtNS
HulWuSfxaALuNGf1WGTwIAN3So4W7gaT2Y9EWqX0M2lmkHto/9/CDPEgmnxyhGF0vhPLqjYEBh8L
glzNgfRdijx9YOILop0XExog2nWmrHWDXFK1qRuLjWc5XzSAZ9LeILDqj94e+rwN8LwGyqdqqxWy
p4NWXY/RiJPsaoO27HHvyvpiTTW/X/bTUu+1zJdhJzHmMsY/A/ojnAYIkAWnp639N/aQeBpaUl05
hNSF19YlgyoptaqLkOy/So+3YEQxTwbBh8hJwcjndvNpb29JfMtGy07neSwUM/ZUjw4Qas60nUGK
eSxRg/XBfOqJfrG9QFXIylYI6dYbbUl/vmDxyBeIJOqqKj/KS280ZMq0XdX4WNnKwQl4/U2fKZVQ
hxULF6SzS753XFTSZeRvJ3BeZNBScPQONKehhTngurNHDcuU1YEDYgmrHLXlG3WcT6s/G7h1f+lQ
1WHUqtkSO8kwVDRRftkZPoGFQcLXY+34JeMV2znWhTJkv1jw8axZuQwW9VOAWW+5Ui80nNxs5H9f
Sthxe/TySVxzArDKxf9Et2bvarlGHLdVh//VBm8dslwGHza/wU3VoMRVotazC3NUF2RQTCSAX8br
0wTi+BRmXiM9WDe+eisqGD9w6urYJKQQeo4cW8Ad+eOOLgYWUhE11VFmugpe1g/0XQR3bwlNnnzU
LFOYN/ifSvny1/qOmimwL+8KN1hMgiiPnK+PcBxDVqYFjmIxqYZEOC7/EeXCf5OnSE9vHDGs4xmh
2VmMEFkGj2VaXd09lyBEuMa6rB0vQdT40xZyklZilPVHXo7mEQCM2xRkbekQF2HiAGzRbnYZ20V9
WgynGlrnvcfH874CeisQqCqcqlhon31fWnNJPalmQriLD2nDbISydP2YM9R2Z5ymBWlySWA+r+hL
xHI60Qoj0IGls333Rfohe2Ti6vxWtgMnATDI7x7JK4VXG/cdt+VE2c4loNWk4HciL6vRCTurAx8/
PguwwqH8pI06fIYUf1uJfeUUMUzeDH5iC4/0j6ffBKRjCV0S3NeGAkFmm/cRg8DpQ1z3TmpyU3xC
7jwkii5L8tf2bMUJjRYzGFELFKSppioxH9P/4X+XhCABo5gHmsw0EE7FXIzi6a4TuafZOiuQBN7j
vjmIMhC9Itirb2UZpa5IwVVsOkqLpZelZPU9/A1B+LmQVbVQbjYzZ88LYu5pZ4UmRo7Mals9p49E
8mBcTpzMlWKgvYvR6/XHmlouOi/JiP5/v1o7DNFsL/phEHx4BmdoBAeKGcApwlRfT5hA9EE/2OXb
CBi+xuyTz4mgatirw/rR5WXBt8LQxOH4i38RIqKLgUgUXs6Sj0SLShqPYk7MeuEoS/3tbcvMOCmd
FlehDaqARXCGXn+VcQ/T2/y0c5IoQ+Az2ex5dArIViaF0b8TQwiULDaQS6d0hFSttZxCIp66+jWD
QKgFUshDWUv0qJ9iHyxTE8+SYhhA57jZ/Nep8YYDGhTSrE2kzepTYlFy6HnOUpKK2aFnUhSC6dzE
4TtgeYjDo/bFiuDgExkYVHnUrV/bt4dURdbXW3AvudFNP0hOUwdWiFi7xDdOai1YL8NzWY4037Ij
6Q4iuGr9FQHlKwja7y5eEbRtZ01Kv5vdCjub/Sq1PkAzEMPEWTVjcx2J9CKEEM4c/NMN6rRKWW5W
TXcEfgbaucWBo3eSQW6yBWJaJ4wiFCJEilhZsFtVQvc5ySfodjNzk60QkKHjMF0YrA7u1jv6ybEx
BItS5/BJgGqv32t7xAzeKJowwVg2QNIJ3UECyCByOZVO+s5aKXQ85VGiToRjpF4/tYyLlKIl+RiM
Eq701SYmtCvt10qA5UgQQv5UiX3LVBHfjuh5ZBw4h4yCPLlHuMj0CBJ2/eoA6gTCJ1fkQ0z0pt8D
wh13hUHHjsQlaS9olrpYge5kZUUdHHMa8Wohj4p0PvOXjLbJrDX6YTeGelyf4URJWnhKsVuhBCX4
MKDNpgFc+1u42g5SrNO5wksCHr7ka/2VUAA80f+rjj2qys8l3gsOAi3M1ljSoHP9PODFXCdpKcCb
L0Gcp+GTg9cwOy5f5z4mNyVDRigkTIGuZaDkLP2xoM8MYGGSaduUa34z2eRmZ4F/ZyT9EOaKL8xV
K1P2RRqNwLGjOVgkwPxC7KgFT/jE59maQBDjUGPlrjo/3Ur4/57iTErF8MX56UDX4P63bE/EBc8j
TEuRs+XCbwIqxZMoO+CDbMX4OiURfIxav+MeLtUtSsV9iMZW7O+x2buQU5F4Uaclhtr9wRXJbKyv
NiiSisD6jlts79sXNoRXlXomBpx+yddZNuFaztvX2TAvgISZ76x/yzN4XxA5O+4IoDW47a28HzDH
TuYhTN4Ef6186CDw+PWeaQ+iVJznhcnfkzFZHfH76QlCHcSg8L+1DzcM3J14j9bqGC14OTUi3kfP
yGE6BMVXE6SSM/zJmTCp0OE34SqciAcGfOntMYOE6fUB9jkWEn/+QG9Kxmqn9Z+bd4lrcaDw3uzP
bvXZRD1Bxer3j6LXNQo/t7gGtVkuYTgu8zVDR5ZwFL1/8zE1/r06y+gdA8Gz+cbbujpLaJ/TIEuh
EOVVXM+ZhAYOXA8vYUe5OGqhmheHVTLPDp4mmavI8fhveK6PxcDyla9rUWLpbtfRLmPo5/45Bwk3
7ug6npkjk4+oBEupuHH2pPKvvNay7QTih5yBlatF90IwGEb0iia+Qpy5dg3WddeRbBvi0m+F8Qmk
zBKWS7jW1LyICxvHpCIIs0gxzJA3+HlvLvcZUorK4pbB4+NXt9WSe/q+09XJ0n78s8fsQ5VAdxOp
SzRBJgIbZi52G+vbLUqFZmIE+PLsosUd5o6JYr2kdGYVVLuNe4DLg8O+sTuX9ErpfRxsAERhQ7Df
ayPrpGlm+qnkJLJJczbGZ2j6+ZV/3PPoRpHC0tMFpLj35zdtoEIW/o/KUH0A5+gBWBWMgj0kvFi3
VX6JCRlOA9FGRUn0HME8UTJCWvOs9ZL+iN3lUhpseM57RTN+LHb+6HPG+TdU+VHNEr05ZGkyX03c
exyeacM0Zh/BUFS7/mwW0bwQpZXkwHX66oIbRh2Uv5VtFQnvm85Ccaj+wLEZRErgPWt+58WCuIMv
n2VkyW9KcRK29MSRx/yz6BczF2qHg9sH9EoWfrwYiwp19bL+fMiPkhW/AIbMB9m8cKQgbQVSiUcw
hYAnycnHxOeaZ8VyEH70JF1rgMyMMhLxXIvYvPsTELARzIpKot/8q6061NJSqnZ1OrRs+OB8NthW
DcLVS6Zmu/IfSsrCWzb2o0/k9NUJil0R05k1XYwGhm08X1JMRkjbS1TebCFQ4ImbphJ5/EdcAnPi
QfxL5bom6dDrXH3YRle1CYeyAqI4VD3peH/jK9FQGY1w20B9J5JKI3uXCS5w0NrId+zMPMyhyK3D
dtAO/3jnfjrxav2P8vzjvaebjbvKwfGVecEHguDghsXKOXSHSZsq+sJzSFfK7424bh4DAI3kdKw7
aZIsvF/jX92jHFR9nYwY+RfAiYN/rMLnA2Y55OB+n7f062AjIIHYaVfIO2PIXM6E6Ws5VtTBVWpx
KySHwkd/qp0bfaMJ0wJlrVG8ghTtZ2evdIzvzxbirdIHyph1HI708qfQTjoLIOABQV2SxOi53TzP
x7AUHAMpJ75juegcPPjjJW/D/oTD0H0Y5qatshjhvBK7hWb6mtbxDhKjxkcKxqBhGR8/S6Hm29RW
x3IURAs4l3XFaBW/VmMmFXR9/U4S35CoSkpkxNTZRirWYBkFWHOC546MlX4ZZxCC4k4CMqczWFpR
wsp6fvEBISzsWmxsjUeWKilnYc4qqUch7FcOSTDwIihhrQyTa0ViRMU2ZwSJsLxsZfLDswNIE1Yf
SSf2LEmfzModTWheKu0rB4qr1cI8oqvpwbSouhs8UPBLZS4wCcGnTBGWssjKWJAKMxWME+g9ffnq
QPBpAw/jB9kY6GG8h2u+2sXGOjzhM5n/xOg2gyEfYHrccGFEMHuflYHybcybmbvoNoXvrfGO633S
8i9rGAlut7Nh4KHucmnh6N8w9NC3zm40u0kUIY7XGnUe5O7tGdfICkggXwIgPrDr3L3uwa11yK04
pEkiiWJyJXhMJlEONe1Ds8ZwvUManoW/eMyJcV1JPhKV+Uu2OiR8uoiC0c8D8+eiqL3O9uv5HxqG
0N69B5X2hgp7DbK8V9t26cPgaGkjHA8m11w0cMd5BLgYox7JPVZXfpODxXkVWoT5J0l9jmHT7F8l
wmLMbUQD8/HhDyoRVh01A/Yx4vb3z/aNpEQOw4b6TemFGr4ZGiWcxvisk3qYuI9t3bbRNHQ02FQ4
nJZQwNm9EnfULR6RNhgYwqPj573/Jtl9IELYQP2/xjb7CxU8BQ1gVkbppFKgqyQpq/prLqY4v3F2
/C/+WTzva+y0UZgnfGEO7t8Ds8jVSnrSE0w2/bEJFkPrsxa5jMBLsVj6Hug9YBJ7Nz9UzYPxQZFb
ZnIHCZV3LqWKY67qukMaKUG9Pk1LsgddIdBzC8E9qJa/p0b8kq4ztXkHWV2fZNysmQKxSWcOWqNY
NQg5q4h7PcvQmCvk3yL03Snh3yxd4R7OfSLEUqxbdRZca3fx8wl568XEAo1C/UCySs/7A/Iof3qs
RczYgqS8C+dZFYenGKzXjs7hWF0wlEo3EODwCoO3MesS0Uzzb6sb1d0BWLP8wZaJoaIAHuKBDGdZ
2E1oQRLfnpK9og0FONO/2iLBhJjdCUeAfwm5xXh4uqqvWrV5m+gmTFD8jPvnfc9WO229wJ6SGwBT
DK/x4hz0zW7Hsa4aYRQKFd0UBxNPTTq+09PpNMv8kYwG739K299ttyKWb2MctpL/tb9Zn/cf3EW8
NRhp6rtYBcxyBwroALc3UxVm5jljlNSdmRRhSl8SZhOqqY1J0+q3rAKQLfp31/BZTiGxA0kASQNA
a8M+LTBjmJsrXLYqpiE8MVfhBLLXXFZ5LW8XRzOzE5El3iGZeLpvOMC9GezYzzoyqHPylxqBBrMq
u+ctvwvbpaxq7mhTHUdggIDXMR10Y7cBQQupj1NK7VMLksO0k+PMAX1LGJjgaoNXLPzDRgcuI/Yr
LrLeOL6tBO8om3ioc3v178J8Z05CmHWZ05rXzRpn9ovdEfUvDBaUImzdic8iLg++ArNZes7a2iov
virS0BT5kNibbRGbCw2ZN+neCQGSU0G7WjmjJLeDlTw6uW6wR0h3twbc/aRq3OCnHe5PR0kO6ITi
0gqrw27Fuo7RRfRzh5dgpdePyazsusm5tyYZKqEFRR23M9VlA48jhNrJSDERjD3M2P+Jinl61c0L
dEnHAM2rUb6E1wzsPv3ucBEAV5Op7y5Fbb9d3Y9cGwScF7AZtsCIWfyW1lp+jQvcel2umlQ/JTor
uPVG50qZlLXxFT1kX3qXnrFWRBJAs18ahEwBQwAalOlPT+jjnVr2zbmK1yR3cX4p4L23vN//VgS6
dCR58sFhOedD/nvMmizZr050xNghQsvdTjWGxqbJ0kHdpNS8VqPoaSBs5GC6+SKTryfcRYso8WLp
sLTG3M6QZrP2BQ8vN7ccDNL7e7RbZwxP4ERtAxTAfDX32kWUtjnQCCgfxURT/6pXDeGZ9pesxoKx
QM5iaqR/FpoXC77onyMHccyQTxGzwulMXOdOeKgoAKWSpENNIOKKvcFDAwZKvEG+E4bSN+3aIa+Y
UH3i0cR1/blPOsZ20o/X7/MB9cxF7oFWMDXddzdfyvDtoqnBIH1hec6vc6Zqlh3+VjIvy/imCko0
qdCD7BGNpqpSZNmuNMEBjWvsOI4pEOrDOxEW6tkgUCmmDdJi342rAgT1Hr6AlbZewIx30ww3eiDt
Cg8o9RwsDmfaX00YIUky84MJbfm6RqGhCR6fcJdDTq/coOcgTI9sZWxhYgUBslh2IBtfJZKR6CYI
2y0AOG9aFDgeFTwh1FqO4HTpJ+7rFEIh+7TWh9kX2CRaXkxH1r6rJY7PmF+m0/P7fUy+7uAEAGa3
IvVzrm80/L2jn7hDkmxzEARS2QoxK61NImq8exq2tvHi2W1d4bn8Xz1SeLqhOFa7mhzu8PO4Ycp/
XU+7Ew4yW4i5KMbf8JV8fugBjy825Zb/DND5uMW0y/R4lzrMc+2V56AColSpmihTjJxEXBfJ/vij
HdsW85oVwjSFy8t4drQYRZwL0uRpVwbhrJeujQmlOFG96609uk5gzW3TYpwPCeaGSmIFJOFwVkMB
oaMUC2cyyTvCupwUHSBOgiqN736WYCqhPYkTgQ7EJczQtxEbip8it7/oabnU6lCvjLeNQVRx1cGJ
G/FvwRDTAsXBGztm7MSwYvHcvVCgk4l9FZfrN1+9p6ReMQcc/hcWoAp3Cx0DtMEhk3WVNON8iPzt
F6TRr+COWTyvlMsboyiVummezxqg2+l959wXTlz8wFTqpp+GeJM+OfBZCeXewSUb5wyrAbYYEBah
xYwPXXZPa7GlBdtLPl6bM+/bzhYf0Bct0MvVJNWeW1zwRaJV+KCHhBp/QOUJfEAtYbhtFRuxwBct
6L/MmEUCgKIUaB+H+UndeZCXzLmaQ6PzHALSH4ZvhLfmP03bgtevJ0OK2NRrqeKnB/26J+72+wXs
8579XnQR4iaiAzcsrgSKcF00FYuLDH92zXM12sYsz6qkj9U5pccM2YJ03p/R3iJTnWOpUNHk65aV
xk5nqUuMpxHHb85IgHhWjBzjCJEqnCOi6/FEzyQN6CJvLTpwWqd0pJBVR9tJmql4u6hOXJ+APCYO
FLZrkhHRS0gLXj4vczdPgAIuE9KffvnK5/Slx5VQOlibKgpeeGYe7AO4pMw3BZNkXibSgxXjt8CD
1ByGadz85CCq2YjMYR0W/Ouu4z+943o8BgIWLlVTT2mDzvXJjaIWwSjvK6m0P9HnMmw0kyuoZ2ff
2lublfLF0fqRAsEifB8g6vwZ33VLWrxTdk5exxRNbL7DDfqTiaHYGD/epg7H4oY3ZwDYq0EcuDUE
t2dDhJ0RgFMhzKpCg+XWKTtkQlwIotlPUNXSVCys2dxTY67yx0HMuQU2AA0hPx6KU0EWhIp/mtsd
5/SJjfS2zxRWrtexh5Q5EiNAG5DwQzvRoi40iPSPTBdRReACEp4FB/2JqV0n0hGILf/BlRoUFTvZ
AZll/auBgbik7uVmdjiribewX1gYxEKcT08uco/q4IdrYtC1nvVSCXxM+UUbPJFd6tTAuML3SpX8
U9K5ZybJvuGjKVGRKArxVZM3BygG1ly/nGa3cOTlkpyEnMJSM3XM2dDAv7LW/Tn56Y41Ic/nhRGn
lu3/zEkzFnBY1IURZmI/A6O98ASG0mdc8Zb5Mxc8I7RB6uYO7+Hvjp5pd9vH9ovx9IkqniAwz+6W
6JEIWTiDzIomia4s7nf1cYp5HNj8R3sc1rUtAjvB9Bv4zUerHdsF47ci8m13b0Cum8nTDC/WKmsk
8xgbYrXqxU6YbP5Bnv9YvspLFQUvzLFjhRy8CMNW019qPpTzLmpSKiKCUufGvFnUwPpE6kWCwy3L
sXkVPi0kaHQiEl2XwEzDTi8R644BOwN9bK3kl6J4UuzwtgR3357rMACXPi80fYmyYftjaL0q5ajY
+W3x40KyaTzfOpfOOLZYXNh6HyAq8lhc9veYUU4ShzTlOsZz9oztjy+zAgmv3O2aEAKVpEiWd3+4
TTVEA4mAp3qj/tjmFAr1O4C1CYJm/EuP+bVMYIkvc1YCc78Cax6IgoQ3qFkIbFOQfM2rJeDTgKul
sROkSKmSxd1Jm5hYDUPkqJOJSXTGVNGr84mMvQ6NiyT5iAURjf/IxSfJ+HcFWy1gv1bHBbjhsAI8
LaSU7pNgUCKlDB6Py7ffnACUXTN/VwgYfH1L4AcJ3EhRoUDexIlk3OZuhAi76/rtABDdU3WF9Drd
mrNBe6/psTgUf/scpgrfyvzqMehLiLfIi+wBYPBe5Shq8BL8RFShVnXtKzww7/vXyfAU6Zxpmiao
TyhlwV10PioBiicF5dy/x/P8ayhqsy6ErFXLgYR+NJ3j045wZEqVFtvvDsueNxNyw8lVzg4TYfcv
kwdqycRUPnsLIQfEasQqZmk66xviwsAv1zZbZ9f5TlKFTmqMG0B0g5CqyEAl9eLN7hzLDmWTiUeh
BgggpMJ3MLfXVxLBZyJDuvGFgJoo3l2dFQcGvkCRGf5KvXCuUlRj8ikfASZOxR1P6vt5MLy4EFYo
C9UOpVnTUbiDCc4UPB5L5ticip3wEBJ2q4QZWm/Q+zZSzsl/cM1qSOIHrmQenZzVmvW+UuliU7Ak
i08jiwthEUq11Zv1ayjGyEAcelf1Uhtp+4dAsPY8P4x5Q49KOFc/tWELdhR8zeVLwnbo+vvFFvSO
QfJRdNjVoIAT/Xf65y8Jq2tnE8v1ukQ8VSe+s/Ha/B20ei0ZGLJoVpa4DLjUNAlLBTe+Jg8Cz5Yj
AMA++a17famXobYg5JhF7rA/i1ZDrD0b0krTTeVJJpm8w9sG3fmP3yw62t/Bz3NqGAVQHp8Ts/jc
XaTMm8dhVv7hPLEVSm9yR8FbKpL/NS/W8pIAH6+fR2kQyYiROyoeFdhahiPJAC7XOmsuKV1H/9SC
r28Xjn+rYeNzM/pWlTrWmWpzhVvsKRbNrqzi9fgzcAsl+2qn06o/vye6gXjUNZ3PZPYpPhhI3Vd3
g5Nc7480FSz/RmvQtyhYLdvdEidSn2tbUrgmmrGkQWJ2nFvz+EFBDbx3csxgBzDZAK8j/zg1RNmh
sS9ISYDGc1J8Dz2E+5ZusV06uVD5y3wtkwviqgVJnsql2PVqxdEO7xQUapzR8eltTmhv22u2Gque
cCQ4n7gp1cVnnGV05Pnq3XKecAuxoKLslDEJxdCfMSHFqi69UC8igq+5oazAATff9qgQx/WZhRY3
W7bEKs5VLMBZtX/Il7jJz0UMKncjMJSrhb3bN19sB5NXFdqCO+/TPL1kB0Mafjw23B6azX4qJNUP
bwuiM7xvfCLGBa+Do7vH1pB0GiZbtZG7QxPRWAOKueTL7AaBfMsnL3zak9ipVhh5aKiq1v2AGfjy
A75bsLNaBJCN6kM2w5FHsCmYRV9b3EHHJdDZ9OWCMAbMATnfeIh7qQUGv9RfgMIS0rRBoxwNc6aF
M4b/+SEdKElAgIJnkMY1+uIRpnbVDKkermqPjRGpqRutCkJLKEEXO7IaXGoH1DEZgOu1sw0e+QkZ
W7LAtjYXWKf7KoGyzfn9kY+mSg59N5HpxV+oGf90kxzoQpN1iTRtPvu0gRhYeqNNAoub2lIY9aGN
Y0bQ9366Qw2bkrJidCooyUZGbtrxx0EUcDZL40umt2VTyYAXb20D32/HyyCZTgZ9uSuOPta2uW5p
HvXcUUFF19O8kpAOYXiNKxvddpNZVyTpfkXEI45xlBhPk212lq5Xw76PdW6nUvZ7Uh20IDKwQAdK
UlOZzo9mJJqiB1K9B2g38l8RZKJ9LSmIW5rc1tvpbbFvIcVa8tS22KL9btMJX0UBqBq6B9xDqswo
+jfExbsVDYFAtmtRhIXGoTvt9Pm8I2i5VYN/qVWQPDMxY1VruShMoE80Cu4sJcb2OprpDQcs1kK4
lC/IMcMt08khXWc9cQUyAz73+DcaV7DW7jLWtajhmMuwqQ/59qwBbLXN9hUYW06xbdoVi+REE/6m
d9XNj5kS2ee4JclPB4MEPbuVOHVlItY5RTFy5IcQDzkiB59AL7iOWiFyR+U6lCo1qYi25XuTsrOj
wLr4sWhk0saeQ4uKT7oe5BIkd7xXWthmpeAZy+mJSW4mz4V2d1cWZCnVoASGgOBFdYiOXD8asnHY
qhSQoX4jFiAcHl8OmzzgU9MzmDCD6lBvwhqOrfXHXu6KmxNX4gjwwMsPgZGZDv74MG+Bqux2bkv6
H2uBTwZi9/nZIWwVS5E7uZ4C3kd0Yxpke6Y8xVnj6uYBWxPl3wE40S4J6RzqwmRaIlKQX/6BLfKR
g4LW5HkLJLmA//m8qfzu0hEr8R7ete06zEVagr93xhXmqfWjleSh+yEDxwIjjfcOzbokacYNVdZx
qdVOlHKjnht32KPPo3ZRju7QgOvxQOtj2xYf2iEazU6PVtGS9Szen/wHLyGuBE2BV4QuAbs15sqa
VG5uhDesDuNZQSR4X0GA2caJEAjS+ueW57mdc+GJQRlZPpL741XrwB3lXrgBsnkUr7zspypjdVtr
gXMDxZR1TqN2ymyg4Q5A47sFqACNCH1a+WT8aPHA4PmNm5qa5FPgW2xa58vYDqukiAVPg2W3I5Ka
IKxn/HuVH2ywhNuPe+JMgS50Ggq4SKH/xyCWAPgelmdtvKoRhu6LH95OxM9/U6mw4E3NfQhhp4iV
fXMGdxZNSRiMF0UC82JV2O5dpW2NQi19hOk/rH0+5LI0VQY1MIo9mvN3IEKVIuj2tOtnxIL7iVtO
Hd2sfcYDQp8N7ISHtq1FLlMCDQuv8Q/ejcAMe0+cu4jxK7p0RIo+OHXKtzosID5KyPd+iQSMXz/6
0ILdmPuLidT7xai6N07W6/m1jYWYx+zD2csQCNY0+3ChZ/EZmJTk9MIPAUoXEsqbg0vVPgWpMEEb
mdUmESnjUr0qWVSNGxziwR2umde3qowO4hOb+eELf/3RqL/AJ8+vMwUh9HaCkEFo8FVCrliRA+Up
AtZ9sVrwPo24N8H7ZiDkv3jKMvvHpgf2wY5H5pHqGmy7hB302lSvUSgqlqRMtYqxlH2Cfj8YPmm3
lDHtfZTfZVZivCBqCKvl9+c5VRCu3S/agCkmms5wafcn1zfwHUP8CoCafv3gma7uASFqi/pulsyi
9CX9bUU0L1RydvdLnzlqQ7xLDR2DYkm28bkLE4MRYoIuaPYxU2j1mF/FZFm1fq0fwjK6bdzkz39p
ilwAFZteDKvKF+isCJVQ9iYQSspIBPCPPCaFTTg9zUedRpyPanRuHV8sRRXgx61ERRvwOtrRrvCG
ATWFKOduQbRoIBtqik4ITzkNYxBqt2xP2L4rJBJb7Llr+R3Wm0yoUdvNMNK4GUc6qC2mNdogiEGp
qweGqJeNxgloTwF/D2J4+QNMgbJpvk8hap1q8bjlKMkndeeIZHHQndPR2Wi2786hoiE20Q4C1XHD
WBPHnRqAvUoF1cXoUkN23xihNYz6Y7WTBON8wsIc/Pmj5AmnKplLjai8Q+PMzPBKMhiHm1qi0/yC
oJBnbU9o42NerYNLxT1j4QNF+CBwpqbE5mhEIAp8kV3SPf3QYbRe2B0rLPuDItCIdQ/gMFvzdZmO
F7R7j25F1gbA4+s8Lv69zuMQpWOmlEx5QKipfqCsVmzFW4LceJpnWgVVXGWzl75a7AF5qHrfZYox
s0sDYkUBXKxMjIXMiOO6ZhCDYjAAGyxG8/pJJg/bIPh3AHxnOnXM756Sv2ZAXMyZqhAEbID2PJPM
Vj/nwCoP6YnhJfvjavwATWvQ69O/6oNix8NFTeu9hvM0hCwY2Bek5hb7teey4/dL+EOD/LIh/03S
NgRFUzkCxrMAFXEBkxMMjXCDfKP3ZnpMJonPkn6PnCyAhwmVwYK833aTa2nWnvksDKrCcswm1ZR+
GAbp2rO3tvAZlFM4dtNOmDfwT6cT0/6OwKnHsngCH80wNk2BwtUP1JU9vhL1kCfDFl7Tg12zSj4x
JEYzuk+tPpVuNZUYlhkWoqq5FGcEpRO/SVE2lIysQNTYPf5OV3xbKiSuCK7izGhHFNr84xvv6Dtz
39fQ7EbI/y8MLSYlrnZgNaRzV7IIuq7eEQa8ylKVGpD27NOA9lgweUW3idDrdtW+UnJDF//KrDcz
CgCWeq9ZHs9E30lwqYyKv6UtE2pkHgow8H1LwNI8X/QbmB3Rj1I5QPxStJOuWMnCwO3SR8h7GnMp
qTDyV8Yp403TsnPBYn/waS6hkDqYjATaaKP6lHyerJFdhQrHblsL2k97LEWRjaKOuAOjSbtRwSFi
zdaXix2dereNl6VmgbwukjHb264QeRHbSkUXzg43JPI8ztnTMNj+lR5YfGW+rYxmeuBcby/gCG+l
9PkscAWKdHtm8JaKM1z49c3TVwRSVH5dNyACAMR9aN85pk/Da5xHY1tkR5NkaU6I2iN9hntmqocJ
WDbx8WotFv95UvDqq9PGjUhwcrRtoR7+gZnNbmqCTctckw03g+PjelBiEosu8tH38Fo07YMQGzGe
cdPNQd2bRfx76uiK/R0fEuaRlqH7/d7fbG4flQiYesxyLBYF5oSbrkKSyo983S0OrpSGc9RkeNj/
gC0SBJ5Q8AZA0yY3SpGFB7sV5NrnQ3qVy3KYmyBKivTIyQz8gtg2YogD35nkQ1680euTeqt069rk
6BjtdtFM22EeSHcrtj89kfxbZawZNxIZCQMf27kHnvhnMiB245bzwIknJxW6oyov1wlh1n3YQXt9
eciDOXWNtkWZk7Feuh6ZI4oBcmi0csXRp7/LJcdPRAvM9iIZ8AVgjP7vGvveEZD90paZeQ6LPVj5
wsC2o8rLrDACcbc6OzVcoLhNNQW92u7FSW4KIbrdgYzGTjK1pJg1WjsC9Oa1KjpcVb/ALASWUFFO
EF9hNHZMKdafYuTy94ApdUWmLyUzVyjrP/6UqwDeNxNw6uq21dcSkaKlL8mMxUa02DjO9DW0uzCS
XMV0CyHoUfgYU3oTSrcFb7gFO0yWWbS9C1TATW3QVlTfkuMNlOEtLqUhZpm6YJcv/Ph9dHXO8AOu
pfzXzY89RL9U1rh8zESMp1v4MLAyZNyTW8t7UXPEC3cyaSIKVT1H+ATK9Xn3VXt4gsebypWduyYa
qvz58TIKMNCRyegnu6tFQfyNvOk1JAAsN8Qv3K9/vC79gIh9BEWmsNH+FXyUbP/eVmLDcz8ZyLT3
ZGEj4ETgtwIkVCZyYbtyRjVG+7PW8XOuhktpoNwfekcclAtifcvzy5jW9RNmfMKymKS1QVTeXdoI
X9G6wJfACuD6UfbCumsuGzVAvLo6lhfW5oNIAHYgqu9pjRsZOk7Uou7oUY0VGd1OxK1UOkPCEdPV
rNbiJd4KZpZ1Spehy1wLhpX4FgF+5lze0PDyZ/zl3YF5lsmpOHzb8Vc/ugr7TjSdjpgfZwKMSgdL
3epOMyKycCz48Baf/FHYI+Z5NXXWXkE1KycKMngQXuzfB65+HMCyNh56BCoCw9Hnzl9eu4Ih7qNW
n/CA5g0P4PATC0n6pZSF0G+IgoOqazF9F83IGB18Vn7zbzxNyMdq2Hc6uk5yB7L6V5Pnd590mNVC
tz7TW0+lj5PH/dYr+hKIConr0LcSBp+P5YucDEii5vXnBSs8gLF7wGyQeYCVYTI773WrRU3WaEfP
0pj2IpTXS6uLODVXqMOeiVkwExAEsogVFvNKX3C/maWrXY8QNdVueL44Oq7VaZepEr6XHXBVhu7K
sltCyJOiZPH7YYJtz1k8Dxxa9QMsLfoqZzBfEMF/gLo8vsVFgD3N26i/mA4eN0eCeMmNjSujKBIV
LdPb9+4GKxTuhg9wWoXY5L8XGQAvOvEhq7l8zjJpHq9xJ3McIjGuOsWxiKlIzEGOcJfB5J95FxoX
FdPgRjtGM4EUZynOmJhuiwvpUbBK0/y2sKmHjeh7UDCOYu1Q1P08UOV9HAnD8eSJsQkoHz6Jb2nL
lFi8VbA+BOETA+4aTK5D5Svr0jj17vLxC/XcfnS9enbEicwEzGKna7eI8E4mz8USYZwe4ZwFVdVS
NMMsQuTH1FSiBFrlR2ve2KMhcPpJM9QNX0gle3aI9yzZJU2S2Ecjy31v908Q3r4xPjLbFMVPaE5Q
dqQhmesEisO4Fjs0/EKW0lMCEuc4keF5XDrxJX5XuVl+YZKuZSDxNzPy+N4BFVMRCJsv15Vjka3O
P/qLkEqz/BJ8r7GYUuGB+tb8rWGwgL/0J4RfrUM6AQu66p6tW/V2nhzGwQjV90uXmsGCoZE1TLnM
xKY2JYIpGioEzQ5rPhnUidA4dcfJt1znLIfVCAPNbprBTAnDlnn7vWnxJxTZCAXZUcc3z0wZ9E2o
et5DeN18gGEd8pSkvIqVRQeZB0/Pe3+9/vZ2DotLWXwupefvKF9Vi9w26bKQEy3khFI43UdBrrnJ
Qn5Ky/0/vzo5LIlvYc8QNWGwRCS8lTPuTzp7q4zkGvFZpnOh61RqDaZtTAy3RWsaRKFR4YRtUO0E
d8+zKE6BiOXSd6fHLIk9W1v5u5c2eNSW23NM+Zs7wPn9pheMtgT+2Sc266oAfP1cvP1gNFAiwRix
NFUFSqCCYPRT1ylQq1KXYdktENcYTa1GXNdMpaRfl6Ysmc8rIWmqOz4mShXOelrdPkfVxonjCFom
H+d1MaBXnPrUwNJU1Ipy10QNmhY8UOiJxMteOc+NQ3dQoeTZ1dztQExouZzpBjKonhS/ixx8UOOg
Iynv390a5+hooj/XxtFMWXw+k6jBmOSFKmPSSjPqoEl9jYzg4zueJJBlyAkXRS8zKZJAACiGLLT8
y1sesBYi1ynKWHhYIJz/Ft8EZYpiMPHshCxNq3wtsGTlh+0Dn1LSN1ncZcg6ORRcV+r74ONVMU5W
wursexQ1A0GZM6/P0I1xygR3pTgmW7n1xwhZVIZJ2ceCMJFdfPakFXTPAnwfxD5lae6oO/WgWKy3
8EgDbSRnJrHDfwJ+gDa9G+6rpwNUoN56rPjSBO44kYg0vYKX24v8WBeWHfkqnuXiG4aSfOLOvFUy
8pKr9ILs1bP76Pyc1/vVAHrbAtrvsmdVE+AHp7p0a9DoMUfGbBx7ba/qKM0vFp1Ass5t2V4Xik0h
YAfgETPbN6du68RQvtOt/EJXYVkAzuAs1v5PWNJ63VTviiDg8+59m4TA/AsGVaX0yGbBAnWwSusL
s74pEgAWwDAsCfpJqFlzNgRkX9R+VRDqPkbBq7jxO5C/+olSwwtTl10rTxXzD+hoAfzIKjDgkyw6
7GRG+n5d6Hv5XiLUHYgrC3GbPneAji00mfcfu+3+HWznzkx5jvr2P2rKgG8a3vn+sO0lTjZe2AoX
/Lupet11G9tb8+ngirv/tQg6Lvx9cCpI5IcfJSUvrEY8uA3ga/zwlzv4Rungdek5XXPRMydyoiF6
tRBhbYla2iketP4DZdesjijiY/EupYv7GiwDg4unrXU1oQRvHxxwMzxcWvx3ArnitAXBmQ9DQE5q
zjn8esFcUb7ns0WvwMqjr5cPxS7asmLunKs32PVseGc126LFcwRxsTu/7BH2Vk8m7X6PBLahrOiH
5PnSJNfNbp49y7dqbj5RYljJidaYDpk25KpKuTyoT3cE9yTGpbYVHc6sVIbTDHTnPWPbm627S0ZF
0ccWmINC2WMBiIv+EFpUYyqSPxvy3HTvuPeBePOt6A653xBYpvkegbdUlbbDbCK2KEIMglgncrtq
tXHX3I+MltD+kDiYQnOrfwb2BLmCF398KkMpFS9bXQL27AzFovOHX7Q5hBmr5+wzaOaQDoJqrpp0
yftaFKvxU1106mHBlF/fJmhGweYgUscCblJBhJQHb7QwUK2IAk/x2mf/oaUYjFc/pZpedluLeg4g
L/Kh5I4lmEGlI2wIWhp4xmyFTJkqpk8MqpieMvNQZ+wYZw5gcI1M3s6Zr26slCfRcIWUfLtjLroT
maFkzLXLbUGYlQ14NDDKvI3IJmcgTBOGiThrjenJ7LlNK2w1dze+JicIDsGo9K43h1dNokvvL9o/
0HZ41zY76bRhrNDpeLNDijevbZJM46HdO2QhcBjns2eO5cLiPg3cS9jxZbtZRa/OSh8uaU5O6Uuj
an2MgTzzhkDTIFRA46JPPLaeendJjh8Jq8BSk6grwBTRxXTtd0fQWdEAlk8RWSSvCANCUA6JzYND
9kjJA5xOlPDQE6cjgFBsw+CsrfgHdpyDqA1m7XgznBa5mk7x1b2rkeJyLzyrOLMfWbDIIRZvokGH
6NtBFFWNMa8gEC73m1Oa6fudEuy/M3Anki+5Sjv4NjYoq1cPNVLgARxOiujr5K8KC8+cB6A2DNLX
AgwL0oxnoBKclMHrIYAs9T3kAv/VWUp8681cjamfbr0xRzelyI1zlsH3l5mzTt/wL/93AlBKdyy/
uSGgKzlbrCDeyyta7LqiDvBgNE8F+gtev29RcZPIcNjcNAdzKpuAOtciVghuJTYnYdB54I/zSuLx
fic9MpwgMZWLT1RVfgS9HFyR8rXIn+ATt1lQMyE8fP6Rz1ycb4ZHI8zeyoXQOGTDvFUIZwH60+ga
FUqzprurPh5JCFETlAq/nyOh93JS88VI8295KBWGInuFVsV4XyC0HktfqxrFy2AYNjCGUtZat4we
oULjXCZ/AJLkOzfaRIdPObpiWsY2QzVGXiGQ7P5Dmw8EowXeYrkjNrPinDt2KR1N6PTOUA+gprLO
ISh9O991YIJnW3ln8W4SqZwAGnQ9Rgl3WLhN9G1j3dSNt3GCIicsAQ5SdBmSmQGGKF/sxLXibu1W
qlCDrWGrATll/3Gyz0MnXqun7X4T2qc7/Hu93FBvlVNXT9q0QMSbAM2xr4gSSxg3jn5D2fHyh2Yq
F2IqkpRHEbH49ItP8hUmFJoIz1Die0qMvqgUiZBP702ePvtZ/rS6Bm1XBRwi41DQbeg3SP3AYehc
TPLJlOLVHom1i8veL1Bl3ey+W0v0eVJTIRGs6/bfr5IKeuFRUxjQCxNR6Zy9IvHfZjaHugWFUCy6
x8SfiQG4PpmnFStdyMYN+lsf2XWY+LU9q3ytKuNDnWhtphSoWGtLGHKKHaqph0/4WomZU2Pplf6t
/aiTN4I40DbswnaF/Qjn7E5L23GIIUTnoIN5WlwD0FfnkaK8Peg/rkp7wXpdTm0kHUAqlXKwvNba
6ikXmYdDoZvLATsSQbIv/E7y6K2wSTGj1pgPAGr4zMzksojcudEsl+ckJPsIWJwj9a9fSEcWLaPQ
wfciKuWCjGVFU+Fmrnx/VQ9N8WGSbSQ+siK9knxXtCsaK6PK/GR1Pgsv9XPQc2lsUoxuvCOHbHZH
yVfzvED9PBDWLrE7NSvGsQ07RgoqSKbYbJdKWCq4ZNcOsso/hvMiqu/7H9A6U8caSzcy9VfMWJsv
J1nBr4PBMDcsBegBtjcUWRDXL4Li+z3YG5DhgeCI8teSGyCGiXefwD8njXkEMJfcA70EHpMvi6cN
blFcPLx7ZpYyPMUQr+Mo/wOt74iNiEM2kzM/7P+uAMBQryBgTGHu0Q+udrj+P9ZY16hh/Ae2GR0W
/uu9Dh00TPMQ3EmHZJBw6+pgi1aeXriLVeaNEcmFt5UhcmyrIP0oOEiQagv14tpyBM24/cquJuNN
bweqZImZA+GWFTk4gcnKZNlbuCeDOHboR8k17LZsXLn8sD1GlSHscUs3nirbrKu+aYJZwaXnNMcm
pFGXlSbfhz7MfFVarIrkeE42bM8AlbZlzdQLJTU7GWdydpPB3udtF2w3l0BzwUT6DKgFvWpcYW5P
EmeVwac/+N6Zx8rgl1J1O0OB6vSwXYtS/DhOOog8uFiehKb7/ApvxzxEP7U/CB+btdrGM6pgfeTb
+Krl1NRnG/veJUzoHXaC6msgIgbDwA6pdX1sbfDia6aTlTDKir/1qNLSqltN9wHkO8slf6o4LqGL
brPHEDVcad0hhYLtfGd8wAOJrFDRlkgkCaTJ4xNnXoBT6jT6SIrJIz0cYaSL1byhEdcMJYNXi6rU
65Y/vxKmnDiL7oLZvTwPlTumkTqapEUFaeAe1qT7R+KKbymz3e/f4vxR5VdjycaLwadVO8v/bIT6
43ZhobSu1l9ltBd14q1VuTvsbUO/oGdKCaIGJuuweLd2UrH1uPseeSgHtCub/95u3qbdSYYF+QZN
xyE4Uvo5qnZBKjg98YGKCSUQifmvRYJZ6+DaOhRsyNmmqwAEEbNiOKuzbcZ8jKCFtJluUHV6+xDP
4ZYF+X9og+pDFCAlJe1PujDJcsHVQSeKFda2yYIfaHLWvAeNemZE/BQCqeOhKF3XtbZ/ct1i+qlB
uM7I8yefNBkjqtxZ1I1s3QdiywkLSmZglElX2CIGAweEv3mcPO1bXWktroDu47u7V0o1ELnSnPSP
pa13B/s2MoAWrGs6sKQWrSaNFf7uGvwZuGLzlCPVVomjWBMot/zOMBZhKuxcL8dM5+w/HMcP7QTW
jN/eizAkeYazyyGad/kw0DM7SCIItUSB7stVli0Dy83in1omTKvKW5QEOJAGSSY83/+C0/uwh6Tf
5p9/chjnUOci4RWoOkI/PfahnmLHiO128pW+iWK6N9rxv1ypuKP6Lo3fRCNu2g+wsya7/BqwumXJ
0h4ybDpYNmbnjbl0FTXrDitOwp/sKsiGMdTRpDenLARdm6SRDKPxE/V+lcITyviWTPmeCem8Tqa7
J7RHG23gc6369Pde7V6OPjc2PyatEFDfMEa2nTmFSaqov5w26NzMNCc5aMDyRif4Z0xhQMg0DGTd
t9HBnjur74QMdhC7L/EDZVb7R3tJrixdQCHnohCPsbdO9ebzOcET+NzdsCvLA7cybsaCcLT5Guqm
n7Wj5J+kARkCXWiXptxVYwiXT1Sj4iX+ozK61YAupT12FOLFPpb22v2COuQhntY5eeGdNNXljFTX
CojrKIEJE77QXL1wT8pQwmZ6j2G9OftA6gDvvMVEYwTVguhNL3AsCEsw88KrDF5enu8fqC/EseZC
vuFmXZdnJynIjnAByzYRAmgjkdkvvAkZxifp4n/TYIX6h1ZkAUdVk2+AyplKZfYpTUTFw4IFa9oA
8f8HCwdIwfBVY8r7W7/Dn3Szd/RAH4hMgcPock/QMjyoekZGeVpyeVE6ug1kr4X1408WPkvjZ1Sm
+wyiMZTlsGFYvI0Dgm0ZioQQ0X+U3IgtKiCabWOLx9KocV395DpQtILvrDR35RHgI+GvB5Cfc5It
HfylXwAZ2DuA0CVdgkdOmKS9SOqrIg1MnMY0gljdEL21FUs90n7Rka7tci5zz7YqNOAoNBlz0M5s
peY0w1JVWqg+gxSd2Ya+GLPVyn/MPsGEXJiSjGsLYCeGbfr0y4eOMzcg7iVn0igVewSRhqrGUZSY
06cYlmU2itCLNftiyRAa5czKqTS8HMxCIaiOR61AM26vA/i18CHLQ1HRa7N27liwt7HossRRyPwa
lykLp83DIZlmJP0ZCVmhkRQcyEMwkQP8LDyVYnt6DhHP11Qh+wWDHLhJmdCPILQv/bmylUUMpYhm
n554eflaSTXM/p+L8ejF96peACkZ2/d19FhSKTa9OasM0aMieCV7E07tdsO+kMfQE0k7qNZMgmCu
JNUOJ3Ex+3OieWGEwsttzizhHaqjeuUf5CfvI3BsDN8snKb7AcZpyV8BEVxPS7ina65a7sNH1oEu
WyWRVIEZhA+5QQU6plLKTjyVXwMjtF1gCxdZlE1VtafoBzv1+qbUleYTjDYvSjX7ErKrthMDT1Gu
lLlqqFLouZQEyee1f+dOzDjDN1lDPyZowPSCAw+tXzi0lujtrwjhD8Dw8+aR1IqOvWMA2/69AWi1
4uSAZVAIH64cFR5iWLNCkuUkBF2w/0zb1SCr+KuUCo2VXZ+d4aCqMpnzTt56gPmienV/pk5ORvsl
E/GfiM8of04ASQTaSGED2zvmVTnTNgxzH7JnanpxkGu0LM7loVssbzEtTW1AK8nAJbHFLHNVH/vj
7fgV0cFu5dm5bQ3/CYW7b+WzCKrwq7MW0dlL6xfKM/w+zTnksfYljTPC0a51W6L7rFk6UJj46qsj
G+3UMwRbcIHhFeKLFrOJAqwgr0t5r7sEEg3lLFIP+oFt0lX7X0seBU7X9EFbVpGRVjTe0zIkfgKJ
relqvhpnJ63FHBDcJzHnZWgrE6dh0VeRxz0TIuERZxEZWY0LMVxJhobAGWQoedQbVDK5SXX/s/l8
X+0FGR6ZhPMXSblPwbp1edgoFatlNhcAOaugM3rRb8++fqRS5J3wmxqrpTrq+PsvpLr27c5wAXZZ
Aqckzb7XmBnKCCqh5vecqvjbtcwWbZLJJVysjzENPGzmAyXWAtjyn1ZKSnm6RoWxeo38BrPazHtm
69Znu6NEizAWHN2xFdPJMxxV5CWL7AESxS+YIb7/wNpjxo1zOs/xIsJ3T7MNtW87uVxazIgrHVLd
paYYaqHNQxpJck5ytiyKF1WxWtUD9zQpzTYhCCB1l89AXJZ+4f8vLO+GTJjcXNxKq2XpjSFjCWjc
M+NS4blLfQWRadUFeMc3BLqI5C/plOVekO8ZqvH6QiaBeKZItc/7FVVXOJ7G20B1E2rY/oHMr9j4
mUNrNcGdFFnckr/sne3CbUXqnX+A8ZH596AKqF5T31VFzmVZuub3gZvi1kAF+hQIRVdmi9LSOBS1
Hkc1BgHmASgUnoCa76H49fF+QwMANVGFk6O0YYlDNT4YyWSq5cUi/E5TiIxRnM9a51pO053ppisN
X3dZ/HYLUk+de6w2JJTZdyOAWw5aQCh7f2MWpW1lnCZB3Fn3DSBCZBTLk96lVw7unCIAJeeLD/1P
Vm84qFcPyXQ6XqhoRmpgFoFVsJbB263YqB5+tF2hS7/lDI1UL2K2E3mfwsQpDYnE+ytfjUmicCrq
f0haXY9HMbGCUCR4ur7MFQotL+WA9J8cnmSd/q+cL4dsGMyMHCA5LwLdctjt8yTjQA+wPV6FPV41
DpJj9FqKDBCj/jSuJm7kRx6HWXrCCF5w0dnJHMf5SJSFeGiwkayZvZ8WpW0cpPpkorE038uzCpMq
7A6kYxWbVkYR+97NWqufzY0Zx8Jf1ctx/0UfSlyE2VdOD8d6nxWXDQQRBWA0fJDpDGkJekAcwuE0
1fHgG2Rn85AF5/292GSqfyVVJvJRYVZfqi+JS+9DPVwwFMgTWqubzT/0L3v7afduUOZiBJGInS6C
sQLOcVDWV6TWEaOEFWRvF2DzionJDRTblVbaxoqzhnHrnbQHGDHRczCCyxFpEeKvu4Fwoo2dwHx3
ARq9P9wAJmLKPgkxD7jTOBqRQdwadXMRAgOAPyDqlEwJZh7MLGyKHxGSf9m7fnPkiApdAvOXTb0R
8nt4PImpNwq0qpz2scMpp7Nntvl8cn0KqMPSMOLR3bdtrigJ1oMjX6ekP02bDrgQcHAHG29eAfKi
A1W3O/Xi8SJm3j72OPZrza+YUoXTiXv80goGJeicZuEqoY7OuxP60/LDD2f1LafJDxyw4Qh1XEj+
oDsaB0UNRV6LdZGq2tPDHPCpy/UPkfEDev+08zEqKn8dolZcS+Tjg1aEPYQIK1Y434buyrTUMcb0
mPkjwWMIISVprGejhBbA6ZhRBuvfrvh5Cc0tfFadqJDqfuN+ynZebb0hoFrJFF9yEjvjhZ3WKq+p
kUfL9pEfjzFtFzD7A2ULVoVlLPalNXD8aYkARSqDsLZjsmAndPB25JNe21fFRjR6uZNHOCX+58Wt
KuL4OX/i4IjdG2rYGjyqlZ9oN42mI4Wo66NFI+oKTl9cu6uTCe72duk0wjTh+TGONdtQ5WvYG9Af
OIMff6FlPcMHGvg8v9HwUbuPnoU1V/Sf0yxbLmFS1KaSV5bWaws2nEvmhJgf9sSdJ0cnc7jUHRJg
A5qtA9C7Q1cswWwDPKzkZNVTlf2ojLm2+++JdteQzuYZ7EUcmGCDy13nNvB3RtjfayLrTyQoP5HU
qcp09FroIAlCCnY6P9BXdXSO/eMtbRezFBvTcGLajF9YPrt5vLR4A01frDPOnzaTK4ys4sleZdwy
1ry56J4D90x+bw5MtLlZXRdlvnB2FzpydV9ZUedzEi7IwNxp6I7Pvm/5cellnS3s7GAlt9vvmDUV
lZH0mggmhDEjHzE3kue2yC6CFrXsEpxmbNh2y1Niz/O7Yj6gkpAkRCGTLoiuvAnqrxHz22SCGMWv
Wk5wyKP0fU6K2rFr1Ig9eyWx/8Gd8Y2jA0QFLireQMvH9jfEzNMUM8esPiz5EvGgH5BgDaYYe/lU
Nai8rnSYIezXSN/Md7+hVdzBgHaBVsYr+Ptg0af1WBcxaD2XZ8MuhPjRbbqUhkiqayhePPJCv90Z
aGq9gaylW4kLOq6SKQcuJW0LRuIdPTq2nOXz34uHxBQ1rkzRPD6Z5e5M0NMXrt/WK/JX3mHtSe9Y
AhaoG47RSNTVvB9XBrHE9r0Z4ckwNmWseQhKILk6ZZUNkn+bjZ9GgO0BGuaVGRIDRJOAacUWZFxG
k9a7Hfdt9tvKCQdN2ID0nEQbLo+nfGHkZwJ0NO2kxcQq/xN/q5nD8TpyRDm6gJS04QB/z4wE91Ig
enNJc/xi85GypTCc6ipyKn6FgvhVJQ2JO3MDAh3VXNgTDAnrxp1yNIUxc3V8k8NcxEP5qZ3cbc+G
Cc6Go1C/3dYM3yCHW9ECCVX7K+ZZZCRQkRMackoazjFp7JDBirAndWS4KaOItPp3Rjl5vV1DFT/M
3XWKJN54TBSXPJK+c7Lg8hpLdn7jYLKF/9XCH3K1qO3ruUUGWsC+vHJsSCbfjhM3bgdrFNlCjs81
tgu+TMdFI7DLA8GbD49WU1L4RhWGIedVyz2VKprY98Qtob7Vt0VLd3hVwAqwe0Mph6iOIt93b0Pz
v4QyP3v1ZCkmgJ5tX5KLgV9Nc9XHnt4dcgx6mQBlbgcQeO4xX2rVu8Y2THMiIa795nBC6u2d66S/
Paej61gaJHijfmb8717ePaDmTRw2MNQsvEPPndedzyIHWpB0O/iN8pJLUj5YVPAXj60HCEOe4RZa
fABD5f8+OwRzFej4cDdIwTVPka/lqF8IOqrkJodh/PcFxwMiaF0OVMUIRl28/L2qoD+Rei8CJx3T
K3y8dEjSnOI/Jt70Iuyph2+qC/QpG+n1SWPjRjb5J9kuUFGA78ZayYztFYn2BUa0APypAF8L+sbU
qbE7jTCEnW1pokOuTOyuUyveNSlAN/yblJ366b2C1vJfvxyg1YMAvgXY48k/ZT6ssC3Yt/2zB7Rn
SddTgK4dwT4jmG0gKeVvXeF1rShF6/dgcgXDHuFJOqfs3OAqZIL9wVpA7ToM+xI9TGOlfpbEBT4+
IkUqFwAv3jWHYjrps3gPwRK+26n9I3ik+vqCy531PeZANTjxOL283XAvuen2OTY3dkmZZjMTN+yH
04TAOc3Kl1sYtsLjdGIzyGmXEFp9f5oRFnyZS5CIN//SNGn/uwRjvUP2tx5DqEojHg92unWNx6ca
HejKgZyki+KtBil9NINBe2mb5UFObXcn9WK/IT1QpIRbPZ4vtoEiLjKgMfAmjuLd6lBZRVSfQ7/5
4UILTNbS0S70PFHxOg80cyXnlxQT9K1nKGnudgWepyyEONvjac/6PYTHffzVE4gfa1rwWYjYLRIP
l1xl177C7JUeVXR8Ku390tSjlZi4JObFwwVBq1RaPfO/MyH877xROEXSMuHF6N05MbemjWTsDM2O
OChkHbOubkAmq6im6KXP/Lc0d4MVjUJxdENMbiz4IPjYRuNVSVAWmee4xKmgRaGjx2hN9Uz5ls2u
0zVZroWSODabcCVuU/dLWuEORUZE4zFWeCmnfNyE7E3M8sXKN7g61IjnBtyY1zssZvWZ5S6ykyha
Kn6E4e4UwRPYOoynpo9lZdOS3Y4hrDVDgLryKlFJGrD9WLKmoJuZZDCQXvgLbg0DopvWblBeorut
rCfYQFnTxtp6b2o75mED9zJpxFg2FbIyBvqaD4x1dzjBB15OoDif9/va8SgPMeIfmrbjOWoKZRIW
NqqMymSGpaHxJjXyDxT+jl8m9g7CdZ5IWia6narQYs5UgFXT1+glLEZzpMVi3kV3+G+JDXnv7la7
Ast2SwLOAQLhig/fv3cO2ybf2QQY/8YVzwVMdT6jhgIV33w9sewn4Xp8k5I9h6V15RLRJQH4dYNx
gqGiLlk1oxqIOM7op3Kd7YIRUeSTlVr8kGQRke+7n+5hFnjBG00N8ulzhJ+0FKl2nDZEUzYS8r6H
9fskNIZepqJky8VIBo9IBldzQsH/MTJOPUl2lC70us2iLOBGa6qKQLeC7MN1lSy57uql2i91Y4ei
BW61AgiO9G4vl3LJkY029cM+oH7T/58jUJ6R1rhB87k+KRfn9CRuQAWY9f6D3aGX94mrH+8YrbXs
HJa7OTOBfWmXBdiTKx9rPVt0GglZmRzopr1FZdlcuiluSExJ6a5cQxvCT5ISqT7iZqGA4gWb23fx
s0zqnLJsmHnQWFLgNyJCJX/70bF7yTz3cdt0kPpIQ2LkOLhzbRdjlJ+ghdc9Axuvv86zpf51cDQX
ub+Aks2uw5ij9i8fTarGD0fweyhDs8PhzsRnvDydx5Vvv84KmGlbQaTpMJAmeKuUKZjrA+fqU1Am
ibRx2hnSqyrDr+HhXr/KrfrMzYQZ/avaCW0GsU/pDSIJVhv60tbucbSjfA0+i51koPFTm2bv5ls+
KlynBKu4+ZfQbGLjFZ+Nnb1k9KOypT6cMiQuZu0NJGq0nWHxwB+5UXq3keMiCbPC6Wh7jHuLLqyi
wtScRQhOGYoC0rxw7hZ/FQNoDzgH2GUi8pukHiltItRwplCd1CxK81dkUUInccpGYy0ufgJ9jH96
nBq0aT0BZh9T/2WEGYX1awY83tS2/aanOwQ1RnFw8eNSThFQGy29lGkp98EkGxWWishu+cmxPIHX
GBLNeBFT39jbUD2iGpk3eJYB3afZka6zTHPrxHHwWiuXlbLlDC0yTlgajRb5U2JitGegTsQW/P7x
KoRQNwv0vSDPuXAqfE4ndtxDRabeWlPYuUvxKUR31EBzueSkc7F+h3c1B+UzvXqo1rwoJDNVAOcV
Y6icGiDzUPALGSuSI6JZHRUpkZFFbi7/aejaNI1AKnCPrvnTttY0rNi4lzDIX9Wvn1xswSb8OVVZ
WW8+O4CoN8KBuVonGS9QCjDtvyGdHfJ0mN+fpBoMoMe6XX40K6gbsE77xq3Rmk1RCh39XwjmVNUX
U/AIxjF96oelze2KaacN0rtDOYoXVemsc390ZJoe3UhI5rmwYZNHMsabX93ylRA1oxEsl3xeUhRb
vXpbNBuR30hao81efEo64hNlDDqW0yail0oYVPMyQdAoRcuA0UfCrOJ8K44pBnC9gWKwyKMSrCXY
648ZRZ9RrvWRn9PTg5GOSV30oCl+7An/cdXz4Le2bvuIapF673lzao+A/PDzIph+KPhRUoDKKW8V
sek76SvG25z7v07BjvtxmvfntIbLuc56N14fBryghwoTJhq/EeGmUo7k0O90eZ0psZboRzlBPjec
xpbc+7SbUaIHEqOaUb7HU1CemouqHf+IQ+++K+vUG3safRhUF3tZ6CQnmqwMNR+5ylKYo0rkXs28
Tcz9WKsOSHjk7TQg2nGtCK8fhcEIHRgAfgQpsJNKPUNQ9tuEK9x+4+3nt9Ea/YzOMkCC+18LSSC0
yMKtQIMxfcbJAwwIsAdzvKUw8hqy7pMU8JYOmby9oeHMEdZ8Wq/HC0LgmlDifu8PIpF8YAXnBL5N
HDxpFx0YYB8RROpDe/+3ppk8cmwL5nxeToJMN2Yp4BNpFV4vCdQvxGOaAWBSeGvY6gzMkxPMcSaO
HXYyy1L0VYUWvCS8QgRtsfl2ndKjIYUF++gnnDjwPO4g56QQbiF31joTJDIxMAi3ZRhYhcHegxE/
uUTEGb6Ny0xwzxDpESb3WM/bEvkxv5nbtNtY2aPD9iQurptRrtIwJEVPwmZUqzzR2l9yaju/WuaO
BuNnL7MQfTL1yr8exlX3p9xvD3wj4zOXFYoQ/zUshoMkoS8rHdqVSgve1+TuC5dsFz+fMguaX1YY
j3LBpKUBhF5WTl7nL3iF1jKtSMhHeX60GGMJVFhx41g6zLiY8V93hN6gDBQ0uOqQvnpXJSAruyHJ
BBYsweSQnQBlZt1fG8ylY7QJIdKaoO8uRnSHAoZQ4unizMQp6VfQVX2bHOWkN/Chkf5NNUiO8fti
/1+tulaa5WoJHl08jfxkCwWmuCJIVszp3wUYvQJx3l6qvgUY1Nq4Y0TwOar2gaoMGvdk4QZC4jZT
QG0QIjQ1wwR2fZHsYR3VHcQLYhUgCY+7DW1XsqfDwXoLmJlMl3ffrajI/7oQE3JZ3ZXtn5Jpnowf
FKSIZtvxqfiVGhgN6CIZegvWgfoJ3QMY+NVvLtPhnA1t12aC0aF8U7hVB5uwkK7pJmpjwz/OTkHP
sG4722pEGjENf+FPYOL5C4tJxfHXShUpKKq+wFnkOcegw2zmeclIDPjmaTNET5nTUCK5NT4nipqD
Kz2hjOct/Ggp8qftqv4BUz6ILlaykT0nyETrmmVjBMexS/Yrc5JTEumanxOSk346ZWVFwPhRa4Ka
Nxy1JIOGWLCjwEIbZaR63mMhf5QVkvOtu+FHSlEfL0i7Tm6GgOh6AqYD1+dQ382xSNLLwHIjKx4p
rhnbkP2PUvbE1GSC6sfwUzmGNVaRjVMXBlnlrsXYpzCb7KFbMRwv9NcErMY1ueUChgJ6S/JeaQi8
+vl+TCgiWkEIIvL2XMPjYmpqO9SP/ynqTq9d7ZOtOmmHkizRNKrKLvjGHEfryAEK7MOh82vS9J5t
EKGRgDjTo8e4zlUzIIWcHdjYkmdNaXWXg2tjiuhqosNQcjCskwCeN7yVTN2qSKmajUCFfY+y+o5b
9fDH3GoiqbRenSdKo1JMGYuTQXYaL+aFgUh7/jIqcTFejKFRRxpQqYISfRJTmFdhe3ZEVgnx0AnB
WJ5k9k1PSwKIvtb/oi6pHxa44UZ7Hi0uq94ST57qYRrBjZ9FZWmXNQUaKKE/6LrfRDragzXTX+g0
+lOdsqEXtyZz0FfRYAVe08+5w6Ede6BGxIp1eluKnUuwPtgpJg0+jwD74LNfeEN511PgYjxlVcK5
7knNg60u/Euo4gM7RcI7vSGB7ar8E8ybbh+yPQlq5GGp2KBYHkYiFiFtgSevZkRCTkcQqvJdy1OV
YhwqcbkX6Xkve22cmw0OpJfoRUgUd5BqaQD5HLGCubWkCLAJHAmeb48skZt1mID+SrdF5gPXyc5C
ldS7e6U5FZg6k/S9jtJBxjm0cIt6rbz0rjQGtOIPMLz9HjEtysc96ctlIhAf7peMdUziDgTuz1SA
VUOSjXlbeHj8lO9UbD/ZrjM1OH40lZffy1H4euSmDs5AE48cUdAf39FxX7uD/ZEIyTa17QTLk0Tf
lbkmLh4hqCl5SALA0iYEQuZw8dqu/BtZmZ/mBMZ2+9II4WR114LVSYw1KBTsyZEf9RcBeBbE/SiO
zQC1l/TV9sqRDD/7tW/K68ac+c0krj4SofQXt5DEMA2ZFb8CAE83vcosT2OL4ST5O/Ul3dFLs67M
6bJTRN/YzMdSIPmSaIf21OkH2TTFwPxtYbSG6eEBq0bfeb7C/K/mz3Wvp1+HqA9JWfY7AQ8nLt/J
po3VbAn0FU1OaGBgcTcqFQM4Gbp+kM6GrodtTdyts8SeO6jmmXeABTk6Ga8A6Yfb5aNfay4DuRni
B/gDB9u100HCys+5VhCMj2uqYDPiSt6TABDPbzeadD2wfVry0PpMMYo7uGpVFZC08YOXzIM/a1ph
w38npWkJjPJMkppnzG+vczE8EK8iTATmnO8JZMgaa2ABZe5v0PYuX5k8ULAKzawS4pKXqqOKlBa3
J6Ih2EZL8LvMDCm/BiQPM35K0mw514bhzZ7wdb21MF7rTOh9YKurN8TbNvZnosU9q7SkF6+SEcFM
EMLxREWn7FNrTNqvcyXCvbvzC5jw3DjrCENHkdf4Fp72YnsxkblFEa2vQynOHQwt7e/7ySeYPoWw
3rsl5NDvhpY7ox4FJDJ4keV/EhMRJ+Qk72bGwuHg9PvtLHDu9jiC/98G0e0bfR0yt8XiT9PmUVzi
j7GTL3mve509kDl+70c43t7bByE0bHeduW7m2oyVbfruE06Sft8UgQ4pU7IveLXE1pPTjpNWTe7F
l2YKVj85ahOIDoFzQ3FJhLB42exoPhLY/xB9uhKPu2PqMDP0w4voa7wuqzPudFokfLhQd7ICs8MD
2EIz0tt/h/tgrG3gdXmdQ6mwetcIjU+YobSUxtODpXuFggSDK403+eYRzVpchUdGK0LFa27o9Wtl
oh4L07HOXiTOQkgA22ToBQGeApZUN5nvySMR68Pm7CPdqp0OuWJoR6jk85BATe961kfQDeE1NecN
K1Gsv/MZnsq7kZnsZ/mw2AlbjE/iRJtk8F7RgyPfFTYRfu4POB3OQY6ooct9EIH1cNrZKcFIkJnT
sEyN8oXQqdsO1UjyYImOpaL+RJItND1QmDnzPeTXU1wCCd5HZPMa59c0sDQnkCQtCbJoBGylza/a
wMCE27bhJsnwJ9Oh2L3p9zObf/76a44vyhWsRcHk/ePweUsGC/2BeXyDDBPsFmq/f/8CcX7XMfET
rMMebTwCr4zcoZVKhghm1IR/0gdBoHglOmqOu9GnMM7tQTx0tnH30n5dE7ICJ67lsTOxtWkcyRvZ
sao1vMvauu6hrnJzxAYpWSGFW8EnY/OaMGa4wkU9QJ1fFFbjTEwJJ7ojt8Sq5byvHRlrAscffgmk
qVQ8Q3FDuuTKt/uQsMYukTjWOwOlvDzJTUHTdd8CklcyYjnrWzc8pzcxAOY/qiaA6+TrhpoHYan3
jnDdP6tbfUVbEM4v4oD4I9okqcIfqSFuiqt7wdEgq7/GyiKKzeo6Jzb3SqhyE6MvwFjmjHqWyozW
Km7BXsRBE8fnmdKztK75sjZvUYj/wR41zJP+XkeeEPaueG0NjZBFohZMo8u4FVRtsQEQD1PZf9P3
s+DikZOO7wzPwRVsWHTR5pTwl/ZG9BLSQXcHV1QKx77gAqJgh06MVpbsjUxlKypoAvaOyUqxGfTt
6gvGgqBK5MqL6nM8GjskLuHxe46JkHa9Ur8zP4tRZCggk8Dqypjyy1748c1mIDoJhRXXOvC6+Vf5
myr2pnMXRML/UZnsTPpZhFKrKNw0Jp/jZXhEL+MDHbL+GJkFCxQX1ODyQBQpbFv3GYyWFayNPqM+
FkxmcU5lgOvBiqvXH4K4gF3K5iQVEYLllp8szZicuu26iILBW+EibrkoRQu3exr+kGDZjIoMOQQ1
pPKJspt63jiIicyJQ6TJy9h4oWBfSVvKFQEUUz3ak+rMNBGHWgqq5Qnn3qIFptretwW+y/0I/thO
7Pb6jcP27dt+oVYlBwCFcosa8ZUACDmZezbmB3Qtu0SZjZsh0usiDab6sWAP6BqoVkwggH/r6fKl
w4kcvIPuCL8bw6VE6FHMIDRDRpL1+T1cjKxGiaklNa3aWq3ZiIJWSBQPqHhOhEAQe/TMN/5hcqFN
13dqe55mudd/ISDr1h6yOX76D32nsWYVYHYFpb/pp1TnViP/a366QHA5IPiZ+6bkdmF5mgTpcXM+
9MkOBPdjrs4d7xll2BBzMNN/6XSkRHmIIN8idySbwE6GYCkgZPj1eif44Q4llygGzPI6rImf6ZdF
Fh1ngOSfx2rsXs2fXoDOXDbtBadm7rDQOrmRqvryEXPvdmv/QbCIwLIL6YJR19yl1uvJ2wX2mfgZ
h9FWlfF7O+XEHclFzo9UcXmrBoBjy1esQh5likM/putb8d7sJsZ/eKgpj8k6Mg8dmm+7QbXd+20d
AwBA1Otbd4Um+wdDGMmd5FJPWC2xmefMapGd+upEX6N4qp000stKm/BTuWll6LMxTPZSXOThfLbf
jNl2rTZKFzZM02PP0oKsVeylQUw0vwPmuc+JCsU4APRHIqS/GU2PDu8dYUemKmb8AGCzQoUGkVKx
smtl/6iT9C0P8cOdWHt1WwUmpD8HY0w0tTdsxsxbGZA6XlZqK5KHX7COFW+XAvlPqgvi0qfTydsp
he85Ud4RRjgO04V6kgYvEFhktR3N5D1WxFkuX87rRZVw92lHTP5OoR6Zh52yPifzxCQ554q/cQU0
OyWtBAsZlZdBJVleQdlKyqMQZ9e4LpCtDnC5J4W+Wy0M7w0gPBPPgP2b9Hyd7p3b2Df2aQwf2Kw2
YMEDk0veGr9+gPs96S6W4cfBqfp7fQ2dl5byNQftomI7ZWU1NTjm5Oaf1hJdrKHduL6Sdr9gEkkx
WCxjpGTCqnK/aWcUOnr5GGVpJ6w5tuSy8UzNda7eIHpb8cg9jPVfwxFW4uVEVWL5cvS3ARcTYUTj
9HUANBMDg4ml6cwYXyCT9MhunwM+Pc39GMK8BY57PGDHpIvJ4u++lH0kw/77WRHZ8icLKPvNt24P
EWI1x7JlOX4EIgmQMKP6mMTsNSOOu3ml0lDhKn6/DEo3O9An7Qixdjr2ywWOthfQDS1ghVWavmu+
CQ/68lGU5nXuMDlouw7MR2DIYHutFsGYWP/uXOw4sbihaR8f5TKMFIh8scuWSYjPgUY2WqYT7oXh
gpNEY4k0OvuTZzpHDb9GowQF/WVvt9NxTAMGN5HVHz2VUcsv27os2Kd5aV5sW7f8/p+czjSl8D10
jSQnG3nq2yhLGCYzXAsEVIDOxyTOjkmLwY7AClmioPWLDt0hTl5CnTkKEE5zDEyJYoLc9lkFvgR6
Y4E79y4yLEtw6kmLk196wOxu1XcPnemyJBusXsh78doLkTmXZweX716K5imFv560yL1FDSrDHsRv
x1HQE+DjHN0gZy3uIfrYgO6liO1p7eH0sRKW9bTlRUYY3q9e6n2GYpT4fgYRhnarqV0ka99Y1ZHz
ZNCSK1CbJeZtf78CjB4HTJ7ht5+7TdnVvLM3jaeKqLLbWTTkXzxdajz5T4CryK5MeP6sdSdZDjCW
qESGZeJVuQMFo1of9wNYXrCslHA97UAI5JOWr1hQNfoIZyUj+Zp/NrRyFEMHSd6S8qavxpzBfriI
0i74w+EyxRWwzoLyVH2lXp2Z5RJoHkW4blA6DyejASyL8e7Sodpsvl4CoRrNsJsTIFP+zXffiYpX
X8p4IbhEe4Erk4YKfTABKnxxt0zGbfg3HU5K70uxMlrEvqMiJUv32x+ELZ2Jv24R/raFgstSa7f1
bx9/VYjnryn2Cb2ZwaHWjCZna3vz7ndWrBU/k/YNk/xI/146n8NiWbswFOFBAUQxhFMuXvQKHlSj
z2mfq6UIQu+68quOiz5gPz2PiG0cudfOplAJ/78r9CfDft8dRUfzZDaXNi07Il1tDrf+O4yBaXiN
x6WG3xVAegubNmokQF80D/BYITPNsdMcxWVGporJKYhUCVmsOJqtcmIl516Sna9ZJD51DMQFVX35
J2rJgcr4B/O5olS9y82V1uDnDPQKahhjTvbo1To5jzBUHe6fm4PpgTi1qsEP9zBAoHfvDx0z2f06
7p/wZvt9bwQoB+EfSWvZkBIz5Sx8OGZMG9G8iGtZ5SWj+DhsHNjEIBZA8qJKeFilxnbNv0cAB1F3
QdbpeONvOht3jovaYLKaab/iKprAx+tgf1lOZmTScxl2d4wVlioJSA3NVewrT3A+21KQA9M7RVyx
FarpnOPcuo5OoiMp57db2al4J1USC5l+TSiUQPrtGNmQtHUB45TBG6mwMJ4cgsA4haIRbfBAfFep
FRZpRUEKTzZifJRhePstEVxSOk5ycjLbw3iyVO+XadxwrO2gO9QBfRaN0fSUy5wJwSL6FUpgTx+v
VI2YhJ45PaTAif0LGF0CkI6ZBiGXjwoqRzih3L3eyspwg9TnibavZUAmX6LbNtDVKMY5cynuG5pE
tbZ5iQzirqRzPrv0YZ8hwMAua10cUCPGuSfTiZ3BqtvA4pphfMhrHU0eSk5+ETH/huyd5XTSBccU
0hG/Q9NW4lZ1/y6zUemvxXv2IJPl/+n9SaAF2IVBlwZ7vH5VWLvBYLgtYfXSwXc4YdgVFFNbKBgq
UWxd/elae4oWCcfjaGxdA2ovxUCTKH/p+ETIfHiMy/lDerD3p2X3NOTeZl3d1LXJi8PJZMOZhreE
oMJF8rYrc5Ukps8v4/qDfUHH9h6T/+RNMHvUNwct20FWUy+AxaQ4v6LwYDXE3ytKSXLt2+6Fe7cj
EvHgqUW95wmhYqrXyB8sbO2Z4d3wSy92a6p1kmfbn0KSyCltIrLJwolhBy2CSzwsvLvaEA5Y+2l5
y7KJ+EVyHyjvc29BnHDCdAL4F763OizAlq5PyI+hFNIqAoT5wEYOil+oVNO6lg5oL4b5uW/nEvi6
d+QQqcLvKV9KkLIM69C3cTb5V1uNJJDc/ng9k6R7Yri3OaV7l+nuLE58HkbtF6FhIO7iJKSp2Zt8
ir2yYrOmKJCDl+aCgyKsytrAOIg35K0f6xEbfwoF/YR6/vllwVZeX8yIywAtLT/RaEM7YhzCn0pl
9PsUtO1REc8CMAUerHA8rwgPc/bE3kXjgaiWk80nzfr8YiSK1qemNTV2urmqtYnyXaTAiB7HZvm3
Ds35NrBtkUGGsIi7TbYG1O3q5U6dRFIR50sVD6AS9txSN5Q1xR09LwNl+PGOE89AtxM4RwY4K6oX
yEJO+mVjTmNGZWXU0b1qw8Q/pqCdVU6Jx9LZAAfhswsm6GOaU0+Iu6JovueKlxNg7AW3Z2PXs7H1
WJ2P9yvQEfFfu6UDngxjRVBYXvLm4gz7w3IuA6ZY2vyX28m2AnAqyKFu2ylfeuOC5/KydyKjUlsy
NFeKVukby9HRncpwMCArDxED6Ldo8KpfGehhU7LNvG9h2SmgClHfZVWkJES0VqtWYGaA6DdEAbD7
y4tN45eSJlsXzRHxVDNN8FKYGlI2zNLxcWOCFTe2wqnFGVqSpLiW+ZIaCW5kiLaB3uNnvKaiuy6j
mLgkaOsTVigJuG6iedaNkiO/dDcBJ3zH3PAzbmQr0XyjdKBMAKDTFjx1xJcmSyF3fxz+1O4N7itm
3mDmcKAd8h+kdFy4HiIAH+ioV3GnmUPTpKtlDdfkA4x6bKqkyuv5ZKbHQBFWuD4AiUc0LqZ4Qwgp
HWraL0+05Q+rzRUazXvgijQoeeMxaot+BVdDn77Zxa4fx3UZbm8bRjOUS2SXj/pjvS3L5xliEAHN
yaBZ+rVVqIOq9dEi7pMfOj/2dj61RGIemhJDsC7dioMF9Ggl+J3QBeqLFf+TG7wOKAvkFndIbjYZ
hoZ+oFg/QDu+fZnBLGfX5Qb/cwxH2kA5kLyMOursKomsHMnlPXDl1vxjV/mDeCzJsUODhvOfgiGh
3Wl3Tql1SZzwRseMsId84CUAqh+g5d7CGo2gOlyOAmQ4nexqdk/Jlukgh61gxp88d67g3Fudb3sS
a70c4Y28cxg49aOgq3Rv91lXFJBRTXXzciIdQhf0r6p1lFkH+edjMcNFLGgsE/rdLoHtkDN4+42D
L+EVV/D7RiOnqoHT1UVnTSkOt/s3t/FMl8ZT4wJhQsuLa4uefmZBas2Q4d4E4CEUGJ4uwioViDuZ
uGBB2uRMCP/4b+IFB4lK/faAxLNGzTHaoqQnTfrfpLXPn7xJCUeC2RkZkpqGJ92Y4mXTXF29T8KJ
x7Tb6urwjSa0R/Fh97mKgpL/uDl2GbK6y32R40x4GP2kNmHGpqRbrbE8EskJFW7TcHqre0D7sVbz
zKFVkFepQZeYuyY7oAnNIgcTX160t/WMqEQk5dPTJIq9Ri4LXTNN06FjkAfNQabg7EJWF5P+HcCK
luslih7qifspxgQKeNRW+87EWqaqJKp2Jsw5eKaGnu9ZTu2bIrkLpvO5KMsDGuxheWmH1jrvmebZ
YjKmL+zwEoZZXtgVMzm60uyefFt8j7xQp13VY6Qk7PFyIi8KTTJAxE9p76hyl/7WFexptXlZQgNu
q/P7ioZ/etnzYRe23DNyHMtJFEy5hEs6CbrpVgHzvXQTPaosEnLVwiGildi1c9MXH4v0axkuf+lk
P0nJDfcCqeeczey1PhZNy02k1CwilwwdrvW9GabhVwuEyObj5An++ebRI8vEAHvzVy4gvVhbQeT1
oSArtXHpccDRVvnM3PW635qcRGXj0Z7UqGBI1EJN84/qGDKFT8cG19A2LsKbv8dNEPTnxXn2kHCa
HunXkk6nmwL0VUJfZicNjktWGEJH6p34V9N/kE4vXG8SkB0Rx0sOXduQEkfUKP5q0togDXpPj8zk
dAz+tHasSCZv2UXmioMVSSsQZe4BAKL6XW2k259mYCL7vIqhuRsOMC60osPBZmpWZFto4pNU0bYs
Ktyf9gXw0Yj6oAJLu79MvmSBHSxZjx6Sbttp/ZzUEPYEBqt7QQ/crVm8pz5v4dBP0B8CUIzdxViB
QkFtPpeKqB/pk/h/rRZ37O0vePCv7YnDgHUYT2cp/Z2LT8SH3onBiQQN70XNS0xUijD7OlAllcJH
KBp2lCgmwuU+93guOOtQ6EiASbEnXKXb8JcPsX65yz20SiwE9FwJKoOXria5HTYh4sv/pN5XI2PH
7gvGecPEVLFafHNbr776kEAKvKal1inmC0pPxZVfBF9xp8amXd84O0Jh6ZRoqlO1aDCdSr3cDFXD
8NvlbmgiIkWb9q/paY0X/8h0QMY45Kthfgr9yp+ywjpk3T2iWO3XF7vsLjvPPxEPqQ0PI0BM0zzo
8kvqm/6kOe263XeBX8DoS5zLT5yTaNjDiYL7pE+LI5s5+RVIyYw3mx8rTr309HQJ9H7CdsJznXgr
oV9RDD0JCrGBG8sk9cWbtbdXWMOIJmWoqNb22tpIx52wxFxy2xVLYmF/j3tAJOChFlUBpUIlCa9R
fX57Ti2ZjfPjNm83jPuWusndVo8QedI+zhXZF9iud8oJpryX8CPVijFxr6+Aicx4I/LlZFkeag0r
RpQKJCLfw4yUbqnZjMe6/C8bruui23sGB4spyXLhIZvOPV2dbRZsIWWAf3o30O+DBxe215+FiUOp
GIzeOu/yhaPZWAbcsjszV7zQ3J9Hp7h7uNorhfXzYkSjhN/+v71wGFTBqpLx8Jqv2SP5g8LQMC48
cFnnDUVFd386LUEVEJj0S2ZN9wO462wReeTP1SlXnUTn2fBaMHXO0q4rqmYhs4AhvQFJHG5xyagq
x2cjqtFLJLksxopC9oNSbkg6B8wQXRGAfiUNlXLcHox4QVM0CahIT14KNzDC27AlZ2Z4unZ3cQ1c
XM1VajqvYdhkH4y9wG+k2jUX71EhDNekqvp+4jG/1TX2igiq9xXy6GBt6Dk9hJtVgXCpnNtAR1ZB
W5ooBB6B/ITULMbyI6T+ef4goTQmsH7OBJ0bvmjOYeX+jMGKK+dd26Ig2s0CwYH+CABosJ6njozF
SXrx35wybrrzkW3r0Lgs0fybbaEtFR/+T+IRQoiStuaI164MGQwd5DV2AEbICITA153FBiiQgv56
Ry96HRKgd8F4HnC8t1Ghir5Nti4brhvEIR0uVJOp/RtFMoy9eplTLRoq1RwP719hk7VUOTE+Xs05
NjaUUjsdREgQ0q2LsSfEG5yw0PVGIKxyGbDkc+kJjdYw6GIJwlcEJvXr9SKYbVHr2E+B/ZUfu0Sz
Bj+r09WC8MY1SveC16/JW9+JOekz/xRVrfT1PwTibo8aYdSUoktv0wJrH9S5tOQoKsmqq3G9HVqW
KkTIwNL70pILew2f8J/OTHO3oaiiFpV1OFaaX0mb7gxMgMcI09xq26IJNNEAaDvytm7nKJk8N6NH
eAkk7uVPxO1xdoQHwauhIBgckTQ5M33VKRcxSZwPGuEI24g9Fm1LZxma+bqrZj56hIJNGSJ+0Wto
PejephjJDGfYxYQdfefrpnafzXgfL9TaJWBaIY7t65wtlo1Sj4dcQtiPvfN4fcMktYnapL+OGr7x
3MRD7bI+X1gEfBKIy+5ZBumqnZ/r/LABMBcHYHMsFw0E9Q1abvfowbMDXfI1m8PIJAI93dYZO9MA
VSdIDBt4ks2Aa3qZMotdbg155W6xzJOGO4ndjDetZJ6L/ov+lM3f4nlT8cSB1hW7dxiotIfh+vW8
9WX6sxDiw6FXl32dp3J2rKVgs+lrBT/50pHy8T3bMDGhLMdv6ONphXtWvmeo3sR2hWeoHezrMHQl
ptI2GMv7rHuLqV/+v2kt0XVv7ZSGRUrVdBSmdRSn4/Bu6TBlXE8oQI1BYuiMwhOcDvQwaNaGckEF
XIAIgcmsw36cR8/Qau5COQdBjZaP94Ltfmoato19TC17qVx/86nad47ga9jEcRYyXK0kKEDaeYdt
JsKLgGwNmls+T7m3dvboni2pDygD8Jai5aGOEfJ8poTKWABHIzRSlQOcAjOTrz6Q7l7Zawb6Wy9U
kaSiPJMdmkO2ayMHUTU/qB31Q2DGoMSSn5JipGwinWIRqADgPRRqfafAUpGXS2VmIYCO40++0exw
SktqD7GPW68i2PP5JKOGAT3glfJ7pTuTaoDc5pHIXM8mF8Q9IuG5il3yVJ2/9ZNWkOsXFMFXLCnU
lUD5pOz0n7oLr93+lwNnb1ieT/p94ZxyWPAteYtKGP4pYPAS04JwvxnKn3R1EyqRC2d/EjRf1oP1
YLvah4lVAz3BDUn05F0Gm1L5afHa7mmg66J1EuMBx6xl2CEALpK1e9W+Pu5rzV09qomUUYl2NmNo
WFlLacrN+zVSLCCJaYCOzL6GBj9GRIzVPr4KgZiMQDgx0PitKva/sjla1U4RLVQNubCX5cQfJ6T8
DKTyLZPkNpVyRknQkdqS3z6SVHUkVtHXw97I0xTIlzOdK6uFh/IZecnzHJJnw+Xh78XSX+bJCRpA
akSTT9ecHZYFFxsK6yimg0wlVDcOQMU1Tq12ryExOq5y+qO1F9s0YVoBeutFzQh/G4lZsKD8BxI4
u402+MsyqYvAMP5zXS+nCezknh24Y/QKdc+y7/83hN6mJO2gArntP1B5efzRG7j3g2d1eG07RIK7
UrcoKBfj3HE+xZgzYUQ9l7IrHLdFN6UHJJe7f460KMe+duCC/4xfjK6pOqAd3hC8KoGr7oVGsu/X
HzR5tDEyqhj7WjHvwvRFwH6eRRpigO/0pPXUQp8AkPLdwm5GzYUkOCtooC1kItrsWmvhvAShgEnf
8WM5LeIRjSMNxtcDw0b1iLqe4/jfMy5xohcuoleJqI45um8ArWV2K8Hpe9pz4iO/4WJ1jvWGv4he
Dx1WqPuMVZgUO9cy/R1ClHltT/eiiE6I1Xhp0z/5DD/psiAeO/33YpKDXOSinS6iCICbjbMdLprU
oH+3oyCCPghlCfhO7axcQ1m0rfad4BEBVWasVckbFdf4u4bKE58vOJLTTRkorGwZNWx19fxJQy00
kSmrChTm7EhnEzoXiwAtpygvP2BYpk4y1MmYIiSw4I6JoYFbGQSGa5NIswoNvHzMQ+F0pNSxV12s
CICFF0m9SzkedAalIEnYQEph9wmDlTYONAhI40ebmOpNni6IOWJDp754KegB5fwSteBn+ITOJRVX
SMaFeb/0+Hhp0Hw7I3qlE9UMOeXMtYvm5ttbkL9/4ofbyavf29QgVHCEwUXTBMCyIFTe2dEuyDWB
J4arPOW59zIMgkQffb8IFpa6QLAQicCz3TPtqknUtdDlB0jS1Ts2U8CABmmGXrhLiPV/hMqOOJVw
UrrM8KqnGQF9My6o49OE1d1L+OpLVlZhS//4kQpOMhL8b6gorAZlOvQac+4xDWRJ3fv5th+0Ncr+
+Ghs94ZM5mqOmJL333sDKH0CSYicYSiabIedzlAp1VS8rOdVXdL4gzSWcpI40UVJVp1QFJD1nrb6
F1AmY1KGbja2Trd3+0O0VbWzjBxSemjKzyG6qtXfPm01tqc5yPGyVlE1JwZRcgojlTaz65quWPlo
IJs42S+c+l4Ims1fGr6r9KVNrH3Kcu7SXaMC3CxVAfn8IsdMJqczs3qqsgNfhcAc3plmhjVflgkJ
52FDQ+DdS9gKHcJcZ720eysKdMzZdI4Kmrl7RMtT0KKp9rb7rNhUn15ML6vqy9bR1rtg4YnjaK8s
uVIfxHESmYHcWaqPBbP1KXK+kMdmioyzeGg5o94irDOeHVYr8RQjhIDBTuOgdrS6ywUp6AsKBcjz
JrU1UWhpinG8nnSjn9PF3vltvjjF2gidJ1sTYF9dmm6tiPdBXzB0E0jqpPr0WdmFyIR0LF2KU6tT
T/KaW+psZ6pyFKI8H16kG81vT2Z9JwWVMhueZZKBZrzR63O9BjYEW05OIfPOXJcxEUjCLSSJt1XT
OA6Fjr2Nv/fQ/yxJ2TQNob9XuSWxXGw216E5hwLfyqyjaKcY9MRuVw+QcyrcvpryzRaJsMVPR9QX
Fom6kpt5cXhl2/mIRO98mpdQdPkFNuzNCWxNUVdj+9ZfGLSBgIqxUJuK5O1kd/69yNNFWsiVDC9y
tZS2u5C1lzy32TMLKL3Efn0K4DDTU9ukT7WMho/6aZgs+FXZoQfqt8NAo+5derD2G/WydYe5sxjt
I5nc4bHW4nuwTbdlx8hnnuSiyE8Zrks3uQOo6SgecGATY22NRWkWhBJTr5Bbjx4WaTHYR/9wUZbz
FWyqp/zCpamUgWuNCG/wa5iv1gC3KRLCWG3CAC3LOpjJC6Yw2H7E/TG5Sjpv2YgccrhzIWmtElCf
BKctfLNbF1aDdggvbu2JXXwPVqRf8lejuY2c3/vkzY3cBChyIiyBXl1SudUMgRQpSXWY9vKF/n+F
4W90qbJdyxPLKMjKuNmC71IMxl3qtixHdixIYeitPxKuoLncSGVqrV7D/gnuxjnkuoaiBTTkPSvL
QDRuM6mhgmmeFebo/ZBOz0VB0N2sbuxsltCJPH9jCrFaXLVNdXy2rUmmdwSub6vrbqqxwmyIjIux
iGh44lCyRZEF9MT4cVBuy5lVYivecNvuqZQcgpwZTnysi3knXM9Y+K2G5+u4avKLXg7+Kn/gF8T9
RRzv059L2l+SeWCv2aB8YVdiy8M8LvAB4KKsolXyFUgvCYs0ESvtei9eAnHae8nONkSwCdShXhVM
7T94nigHaMLEodsZPBXKHHQoph7+ygTnmZusS5y7jGAR7P2jPLs3Ey7RdRT6bedrSSGoNCILmpLm
Ki0sFVhKA+DYLa+Uljld0P62DkYynJIqXfguVfjqhxKq5CACQB6KYEjNgUwGopMDpnsO+2dDGPmd
s5qS4OHRn/CB8kSHvxXQt8zRHOa6HXkU6nkNahKDAeviDw1T9dccfhljlG8k4wmk8qpK0e/3wApH
I/b3cQIG29GkO3ROVy0KV94R1Zc/Wu/f3jqnKD5frpFJs/ZqbFK2f9GDIdvOdiGd9x/vWgZy9Wvk
HjiHZJuHkmdqYWlUg6HR8UEUnL1vT0J5rNmvhC6qAEcF7LL/YC2rHNQ4okIWnPFYwjBYUplagk2D
SRskJZ71gfRO7HHGdWR9po5g1TvXGdcyYKVxwJhzKIFcqsyMb6B0iBTvs42oJS9VEEL4YvAoL1M3
yeY3S1blwZYzP3BOcPryQoFtlim/ZQHq4Ul+a5pk5LWSsCE4dv7/iDY+fQ+WUqXj0zkBQubaE0q/
9eLYsSGaQBn0GdOjGo99JXNz1XT9Dcb1ik1m8+udz/9qa85HeTpYvE0dUCLtgy1HGEjXLqfTpuTe
p7QZ/JneEz+EdOOWdETe0SkJunRZBu9t5nFGPp3bT9YE4s3hYgzv6ehW+BMp0pVeEkbxqd9W5uoF
fKiQLavAHAmr7h/HiFwcioaahsRzwCi3KSL+9gfb9hyQsXvuZGiobJ+htr2fpEprtcXP7tx3zJPh
PLy6/lLi+TgY3MWDMmpwJBruc5t/L8EjGHa5mcq5gCH/64u03+vUHW4UjbyZoau5QWgwvMirFPSr
3Xmz8tA2fR+rDa3OSc9kZRpOwTND2GkFzAJUYwkaRVOROlKFvcli8mxDf688TwkkUy8MptfCpWYm
daxSeg2kSZQCG5cn1hC0EHH15cqwfqY91E6OHJhumppo23le2jFJbYhlV13p4TQ7QE3sp+260MxB
pU6lFECSiIB4xVBWqN4quEck0LIXzHrxiqebMOwqczFPFm6nLu7j4A4774Rp8d2ByLLmw99U7dE4
DcWTOTb2iQnF278N7QZ0SvnFK1R73XiwaiI/NLG07XAOe6kao1EknDh7wv3vzb9T1swqO1GW/ahu
uh9vVRph7ITfzIqZ/e6E0o9unV1iRUUdTvh32bOHQ5MRSxb70jdVJX9tllAKr1EniEidVMxV2Pjb
GxW5nDdMVnkvTqfTU94DqlYKMDDdFbIwrJx8HOdQ7v0DgD4KTIkmJZuIcyI7unb5Pc3OJqZvF0BZ
uCF3/IGwsSDtMdH1rj6i3U1i2iQISeG1neY24tnSRCKP6cVjgGWq1GIWGQ2bXmlDZ1brNNA3924t
5lY/OteqHosjOMbRLRTtI0EinaXayiDQMWGYWqs9C9DPLKTiee0f+gr76E4r8HmS+JCn83M8E6F3
CjyjkdlrS1rUlG5Gk9/o+Nz0u8hlNX4x8fhbWj8F1CMnutIsn5gJqpWuPaNjXZB72RojfNgDMGyt
HrRtd3E7cp+NySfhLAnjmd2tQ1+jqYA0U/yprIqtm5Chs4NOAnIubEa1BeHSu7RIgqwshBNxOZoO
kztmuhmr/jGc8HPpnUqisRAy81EnbUiXhL65Hsu1+8Rk/2P8JqKx3IxefYUI0LxCg/p/vDdKnYYw
PDQdAuJadT7RpZPoS5+0SKre/AJ8/t3kiATTkfSeQS/bjd+DAxMb3eFK0JnAWl4fZhsL4Oc4PgML
mGr6B9gXL1woiHE9Ya5dkKTkmu3XpSRDeEJpkihz32nx5+RRr2RjJqu0+9I30XqpB09z7/k0yVD8
vemtFglKVEhVGwzxsRwPh8Jk+4iR6FbzhXut23QVHaRDZHeDZORstd2M3HJv4W2VuvMwP8YE1LH7
O2ixig9hD8qiyx0AOk74XSrzGhNKbhf3/Oe5m52ZxRANZUMNG7Hw/F5PJdYoNLsUZOAoqBZYXm8f
wdKXJGhku9MbSTJlaEgIMuYFHyLDT81gzeW4JPi2oAgfuIFt3nF1NN/JXagoJqyuAPgoCAtYU/bK
zmV1D5ZkCchhe6LYjF5S4fbhPxqel3gAbIiFM0O5pjq5Vif0BSRCS1sGko9TObdAAnT3HgqWHn8N
aaEJgx/kyzRypahY0kY0+0TRfH9fRLuD7jueoLulUKGwkR6a8oaxWc+j6ranvQAjTu1P6HfJDWFr
fR8hMH4/05bxsL9bwOpZHtpAK8YY8Ef6PC478hc1Pa6E5O35gg27PJwc5xodLTzrl5SesaYmauTD
M+vZA2OhrJSeErZAZE/wuYe6WJ0TP/2zwD3QAc3qOM+NhS1kfNprieCQGxG0Pz4ZovdtQZkbCrz+
uujm5WBR7gvdIVv/6tm6MYxw7uwSy6fLt/tn7w76LbonQwJchcOE6WJrATOpKMHQTTnTTMbgJe0W
vqOV7YtTtRiF2+nxl/b4tkitUsKrXGC37WfgWELMkQEI2QudAPSuRPIVYsno2EGc+iZPzpQ7p7XB
INjBFXBf8cwBBh8WuujPV8fqndBgsObY52fHYq2XeHqNsKCoLVCK9Ha0+wMaSehbQkjw7ZuhFMet
OGW+LLC2VWKBjgsafIr5Ky9LIsbGvWkbyWG3LdSuZkTfrZ699jl+BFUxJFgPN2ji5pNsLtaJiTpP
lK9HaGt0oGrZZaRyCrK0SPGQkXQ4oyBV8wh4sOkbBOA2koKKaub13+JAOLSHOsGWmaTlwhG1GXh8
gM+peuqBaNiZvvnf4gVRFGIx/DNVGdxzReSaanGShupWOlQDEtR4FD7RBA5ee0E/9x4NP3tuRxKA
8VSul0u+NxFW/TI6D0A/MR1d8OcUaIrgPrDQuxPboVmTgDriyjxZgzw0foBFhtzaSz/aaKDaK7oV
NWl59cSAsb3E0kbVaQ28D/80VFrp0PQDnzKktcegkiazBhdEIhcfr9s5kpRZ+4oVXi0iRYMpBydF
LklM7i8zIlB9ErcWbgjHaV6aL2ymGxlp6lU8tja4REaxutc5TajTMG8RgliOr2soKsu+1k8KfEmc
RALWf0flnmiDuhNoz4rnQyYcb5QAsQ4Tzg8CeKLNmyLx4xgTg4fqVZObRWpV48jWgZnbAtdC1Q+0
Fe3dxasNj8YeAuP2RirRnMHO2oBomlFOwmTJ009M4C9C6dK/mT2dm66PFAdtQ/sTJ65JDFQic4tl
OQ85/0RyZhCoEoGDRyFAsVH+smEAlCqoAKMHhrT7AVJQNnIkhTyBY/569pZcz0WINmZK+sf+4GS1
4Cx2KJ8t8dyXaI5IwjvVQx7haNa5XdnujmQELzU0OUGGeHJXNBFyLhX9ye8hz40p/VCekSKCbYma
yJWSNKFX2ixMrd+aDXlkNvoFko9+htz6fddOQFUEHuIG/aT211sqvO17a8oK5zJ/IiiH8KAVVY/4
YNLewODgPaHHaxZAAFeXRi3J6Y3PyjsIiQ7JxObMfmpQAx0j1GXx3yVpeSjJ4z9UL249+xhLhQBm
VEpMiZb2VfydtqMC+zEU+WwaagEfdI2BmXLs2u+NVKSRAmSEheg/epnTJrq7R89pHHclGMOXB9pw
B/FgJoJ5hc+Q0JR14V3h396r2QQTQqvDGmjtcHITh4TCz7K3HbmOgDGJDjlRfzG9Xs0XOszzYOMB
72TDvbICh0PIUFuvQ/c/+ybjbrM6Fn+16RagUBkKHygySbpYijNHXmRdcw1fB2NOmANlv4mHl+u/
I7O7EFYpKlEfJghUG/0wns+qVNi3/0CTZRiLRfT/A/S8FiDtJygEo4YUcNO6TNK2kPTSO+Rqq0s3
yW7+hV3Ck6XVqYjKoj/znOgvMSy51b5Vy5dWBIHYGOtj+DV64sEzEBfPOc4fiOd/OGjeAC6ILj2V
6ciJogTVA1zzex2dniCTNmgc5lK4BC8syMdR3q5VdEJHGbXIl8kivLIl0vLl+p8XmxWoCoHqp/ge
HVSSmcNAAbdN0PJmiE5LQpVaa7tI0ZTwiLLrtkEFYjQ4G9e4lX5xOry3aVB+jaK70NxFNWofJ6V0
Dp5gGSianDEUCEzRd74vomA2ky6mC3lESXs13uofWDiWUkuE62pBMQw0kquMRrmHlnalQAYzUOxg
afkK1P+m94d8xc07Ikkv8VZho5effjeycdPZTfW0ut4nIv0mOX4vedYBQts45g3NEqiouLFxJx3z
ge3ASb+ljcESdWKmfAIH1xfiJH+1HTsabwMc7U2B0XopFvfABnqpOpbghvHEspWwLrX1sT6MWx1S
KnyTGSB4L1hOb+pK3JYhRTQCCkUuv+pFeCGlD6fFwakfp+z6RiX8XlXYcDk7ET4r/Q8YLcsM72lp
HfY/N76sDU1guGdbWg+LhqoqWe/NkiRbzDIrbxyNyNexf8B/k76dQVVXmPOe68s017v+1jWNumwb
SErGgmlvemIkXf1XuiGXOnULW/L5DV0ihVHAWUjv63ltHNcTRpEqmlH36c19Qj8fi6NcPFv/snqo
unAonPcazx/kFYJvIJiv75ofwpfQE4dtkAJRQj1CmFVrrEmfSIDuLfATLDUR2ofUnOCRPiVMKsDZ
rHXXAmySVNYWLNAvEeVS9/BnxxRQoDDXO0R1XbN28KdgcfWEV0oEgiQd2wDlHgp5M0/KzhSNSFeu
pgCzGV9LYC5GdtDQqkYXrhEvKkTrSP80HSziGz4PyHWHXzgtm7BN1F2/7NLjVTrY4rF0sNlb6iUz
cJM36xjxtSZCk5YDg4KgcrB8H1lOUEMIVS36z64jBUeoClsufc4r2qcAYhVW3NUtGJmAQE6vGW2N
Zd2FjsfLoL2gTmpY00D3+LHDTCR32S7MS7tA7QMHCOe7GmEZTe9YIm7s6XjZHa/Ddn5k+dIO3zWU
4Gx6eEzHCEzbhz5XDZlvu298x00MOHIZBftTwCGesLIJ7Oh1RlH76dFW8eLAEWw8OWuLfl4LH6s7
zpyM5vxiHGjYOdrCL76upxdFeQx3u662p9qaAcIhecz5pWJ9hE69t4bN/gq3jceLMbpuux6tn3ju
Zf+9Hc/xyjywq3ahhlStdNix4pWDjjXGWkZGb0EYHmpGfRwZ6f3i3EzildaRNSiJPnmzS9OSK1sV
gbeX07wHrBZM/uPIGSGuZsGgwlEUquJnpBECz/RwKFNFWh+SPfJ2YXpF+ANNwq/OPAhQ8tD9JB06
kW/WTUYZtEPZOk58fLXbwAI62EzoVXyhsmbML6NIsebbWNra36IBOQkr2yjOjDi1EgchvVY3u+fa
QQt8yeo7pLm9Cr3IAT7on06I1l4uUxL00kqja9/gFGOpEvRaZKIbPAGefcFUqhdAsZNpwvPi2b9u
63RgM23loAcZUmwLaTBbY36TsV3KawUJzJtDW4xMjZIjvlcoT4vN9Ru/YKQ1pNnHvolacdFjAwzu
0KMTPbeHbfzoiezqyMqIxqQhJTpkp2x7TQ5sxK9c7gA96ARuajQ9PN2rH9HMspsW6t1Wcb3cjijF
IIaY6KSqmOq0Ofz1GYaeUJKedM/Bm9l27SCosmtbFgNqvhrlpI4eF9iPwVzgg1x3FqXQH287IANa
IQNg9npCr+FshyIhxeDXDIs3lC4jF2z0aAm0HJMSYFMyyA18V6IY/HRQur3AFzC1ORsdQF5aEOf/
v7tb0O5/zhmXlEBLVOiq2u6/7xfFFzOD+Uz6ZF8reBWXlnfyOPwZ6TpUX/o00o13TGG6Owzsw8nm
PiteaiIRgO16X2FEEueQpewmW7JS7EnpcVMBoqvO53zMw8KPZApjW2I5SSvCkIVERA5Z0PgoNZj7
AutHl31puynJzRmmck9TLBp86CfNB8beq66A2QvqKOwgIbuBZO4Sd8TsxAPAGS+Ol6D0Npioi7vf
Wplzt0fP3IEfvm7DApcciNalEHQhKGvV08FbnHPV5rDUTn0hb90ZOmvTAUwpg/93bHaX9749lnIg
WV8Zv5/g9ftoBY3bTS3pxzhjzy4EY6sO0OF8ia06/n065BPfu117ZyfyZaHIZQ7/K8N0YmQ+FY86
hJBNyyPH1TQEjuchTrU3cdQ6C3+JzXLFo5PRBNSDesK8Kg1QI9yTrmH/omT+gUZBmTCssEX4pRij
WWiuYkVZu5B1rhWIKXaoTdUFK4B5F2wkG1pmLa46BvN8B0/TfU5N0NKJeNalZNqLaKfoK6AYWsZa
sIGKNy2jYWa9WBl6O8VaRm2inPwAeCmrL0T9Tafzjkkt2Vg1Lbkq9Z0Vx/tcdzZ3b87lie78QWDb
E8pvenkhCjGBAmKu5qLaizDXb6d8AzEEhWFBKPcuVaVNzixfXS4oG09ftdWyoE783wdiB8T7RWEh
QeNWTB0GpeQ8niJUHMbY/lbT3t00k9h5EdGf/tE3VAekT0+1hue67y+KsMjT3vaSjvATYj9qQfLG
Palayj8BS5jtiz+W5qVuGjiIrnM/B2uTapY52sLbfnIaCIEoTEEadMcBSVkJyVwQXsqESV2unXiz
7Qfk9Msfs7M0jV6y7YYVTiyMuUQwEFcDrLIru8Yaw7fCtgil7zDn8qZo5At7e2RnIbPKv2IMnL13
K6thuV1T56fTvhPp6Ji3UDLzivD0/C5wvhi87aMAKxdl0e3OlZ/ZGu/cBXIV3wMOk4M/aCh7Xh7l
G0jcRL7K+UCWas1ienax5Rqs8tdtzeWCB9CZzK4M3zHBqzX8egBuxEY9AyzTSdWcvN5zhZSmPeZy
DzO/nNMaXQwDE25fY5fOiKvdG8336MShQpdqkF8uJhxOkk4x493+p3XzzODJeysoM38sRm+cVcpD
jMr6GVuJReQ3HlzMU+t7vPiJLdyStV+gVZvpYmYG2VKMOkwASiH7c7nus0cgPpp5yJ41qaqDKXDz
WTAxj48AF2w4Id6sdu8xvZLP9XOV4WrS1id8Xdy48MZW6UMO2U6kceFIhu2/RNN2cyeFwoSykP57
xHoq5S6owHvhx3CwdGJi/WUB/ji8SuvCLyQ6itNvfJrSaCqelC1zTrTgQS7P/DbrZN7NIWHw/hCD
W+ToeFFtcWXCl5uVMKLpIQ3tQeVNmt8cbg6ojgFhS9gE0JEcFbM6YF55r3bHgb+czICCSmpWqRQM
ixqY/s5ZLp9RekvrKrDQmaSdpToy3jI3l8dYQtamgBEqfilLnwiuoNLaUVUMQBdY0/U4mBohbOlM
VhAsth4ZE1DNCVusiyxCPPGvlttlZQGKQrHAeHRi8vRXvzukhRyXm9RgO8lek3ajzvqSOhPHFHcx
jgIQCAyDQ1z5bwKr9s2dZjZyMxBU1scsreB2A8XqwWB/0Wdmb92K6L0bG9sIyKM6H/pSJiNi0qL2
vdZFtrWfU1ql1S3b4ZliuIjL3pl7xuxzMGxinh9ch1KH1e6GZJKAZ8oaN+seyD2eyVHymdstx02s
P/81yfoxJxwdSKv1VnKL5wk/Xj+zJqrI7U+BrJyCx4SkRG+LPLYGdtkOszTs4/zv1bK+JuOPW1iK
LNbj/G4hEOMRU/Oi8BfSdnVxj1BslgosZPoQdmhc3MlqwgoXXiBdHE/jhKV9TK70L6/7UIHqLZsb
TeNV7CWm+mimKBFHP9QFqSdpHEqUh9V/0BDEz6puppfP/oJAarSPU6g1jGfEgqU07aWqQOOXLDZ5
cGV3LB9NyQBfWYN8mSpdNgVsdPWZyrnRNWdYlbQQbRYlUQGJARU0VSnToUCif55ka8nx3UyMG4FM
2PfNqDA7+e9rzfLsospjWcjPIzxpBVfMEIA4KR3/9Sxq7g1FPptykwBaXTlri16CY55Thl8VgUOE
ZHT2He5BxoDu27kSogdz3K2YrhfHxTlO5BMJwq1PNxo9FrTHjDHW41s2lyQEPuc1B/Pbl9pVZYU5
3DHl0UP3ZxKq+3sAsYTYqacCFK2rNWosN9izAN/kyseEo+1jSesOm4DTjROs96L0ubZZgdOfgICH
c9W1QULON2DuQjwdJ9/i4S3qCKw3czPnhEZcF4gJgSt9F0ImsfoNw/HOFFe1bUYZSkGBMdBKsnR6
x2j/CTZ+NuzcWYtabJtbpqu8gVDoTzPfNwaT1wvS6+bAXfcOJfETw4aj65oRtucSeYvm6uXOUckw
J5+hw/phiXEvo/394SDujpi5b21Og9fuq6rZcR89fl27IvuP6gDdGuS2Z3psXcNjJWxpAKNlqNv1
xky/oOLd9EJVy42DIT4q72uHWbpb1YS0qLKzoshzw/JGRkVWkD7sKZmEGjb44ZkFyM8SqXs9+Yvb
vrtROHkH8M7Ky13PeP8VgPXUsJu3RxAVEnw46PdbLNuW4jLqp8qzZfGQb51zLKfvE+xxckgt1Swn
H5N0FmLr37lZGHczW4yX0kC90Dqw42QtqlH7/mAHgHobjHuX+HcOC2KvPHMpVSKuW0/xardk5mLr
a6TQ3KWSdMJZVXtMv8KIF0v0QX2ntoR+CTG/98/tI9fhN84AmMO2yprRa8nF/aQPjk8Pe6ijmT8T
X+rlDza1reL1cvJgArr0cOHI2Nz6i2HzvWaluc+hqceSb/VcZIu30AQjDXRPfyqMgGf33CQOJfLM
GHeyL49KlGZUeU1a2xYfR2CbFJpql7ec99aMCEtH7Ay/H6iSz1Id/X6ktiDFcfmt+0legz4bE98U
25hkzxS4zfQEtpnCGYh080Nrw/fFW3cTBU9H7+S9vYKq42fMnBNbM5SCNkl3sw+zXUk9JyJW8TCv
lpY79fkBj4Y+SDpsXGMQPOap6r7LOOHELhUpx9ECaWYlZwE4vqjTXHTWV3ei+gnWvpm3wSKNCsF5
qLQDj9ETvEJ1lIfBD5Ufnyp/P9VIGZTllJnZXncIeY1kewQrb7LwjL/YpIlUnEHzeDrb3P5W9f6E
58acaQ3X596dE3Kavf7QMELdrUpxEs78vysV0f0phdRf9aw5cZAHIRxdxq1DkPlOOxzmClNvvJah
iDA5AajUdNSm50JnT/7p96ev3hPBfaNQcZkQizMQvi5/O/kgeuVlQdjYEL6P248Q+vU3tiHc7U3I
f0wRtBvUf+My267uxw7rxCm2D4Xuzwm+jBzyKSQvl60Mw9WIZc+Iyj0tzjif8/vqy52qja2mcSWK
MP5RkI/oWa1EoDmNYLbZqg9+gzMETGXb7zAePZXblGH61QYARVesMTdMNx4jhQ2oH3qzjiSxrHtH
u6jHTAvSB6sYiS5tMVlkfQEgMXAU1pH4N7hRUTGWac5EIl1tI4eZK5CJLnAXF9I3fpgoXw0VXDG9
wbxtGt5OApbVLWybSE/VqZoOmdkavpzRWQtEg3VMhc+ePLG7Hsmx+ozASup/rBqniX2oSfD256kK
9U/1Aa5a5b1wpEtpj6fFc9ixY6N5+2uZWcJ858yIpavSBPf97yW7/HOwFq5za8oXAfUhDiz0OBtd
0/AzC1RomT61yelKqGTbp8NBNUq2F3Eo6yBx3a6wh5yquz4qVjDxNEebgexiLx+B0oWmsxGTwd5H
f8RsOCJOrk8xVzlWnPqhZoqOjTzbekfzlPjWVQWDBUIaO10IBG+oqL3PcOXqOszuQyObNAg9cwUg
Ri0hpMGqTbdZi4mJ2zSIEmUzgv0pfkdZUTid9ESEN7hx8awBn72t+jw60hP7Fyt1b/XRBihlVsat
6uBVcYmWWJWuFTlae1eRFCHXc1vkrB9+IMqtNlZlAHJCjw0GWrdNWNETk9ke6CmW96s0MyYPQO2g
xPE7mS2aUvuOzoAv8MrOuKyZXJq9LH6nuDTLmNpV6wiP8HHScsCplSHmwwPfLlKd9Lg4806/LLKt
lHPoVi2djh4hd7OFV4RWayv/iOKj+VPaIi7f/yhQArXGlmqDgmLsVhJEUb3YpcJoQyRwUHwZ84ij
8qeSfX//SXSynEU5D3d+r1JdhdskWPPIEdUiINU99RQB1eHc3YvAf9/CfkEzWuiL7IsYwrABBEX9
6OhBmC2PnVOCHfGzuEQbKQZLtA9+NaYTvXFBDsGwbrYdI0azOO5uvz0FUgAKmKcyfd9FsXl9GpSy
yx726fMpsWj1W4nynQlCWPo2IyBgpDnSJGkLjvMFZJTQCPMl1CvUmQvzTVUFAeRqRd2JCgPr0j9D
RHdknqYmaYtXoEiFtVFg5vSAW2cusDccJqa3U6iNMosdbf2kxPv9MPkswyxxZ3XZakgtFNzyI9Xd
ZZkdHSRYN2ipbU+6G6/jluxGSXnTbhKnmLRncIj9CF/iBpGRvsq3eIZTL3BCUxBYiGEA0mAQ9e1s
zF5UZNTfM0AY/dha9kfD4e5jvM0SD2myo3KCaFDZ93i4HsK7yOrQH/u2PKxUouplGfbc6Qo/S36R
YWJf3VZPSeeRxM/ludeMYOH9H7tw68H0MA0ZxuKKJrrdPJYlHtLJH1OMRketVwLKhej+x1Z5xKvK
vrAflaPJc0+WFMRIGwX40RRl5Fjuj+etUuomUe2TMYKkozqU3Ukf4IM3rNuCdHQM73iAskEFOc7f
aCEYgMq35BTnSXIVpeFW6GEZYVaay7cmBMJT21JETQanHkRQ2dqSrehtCl3OZ0E6Ow8nsPcIudx7
BywmJyMOXQ1H2aS2FHSRSVdpVby0MRFSvDALFQcxY0vWcU54rSUXPprNQW7tZrTaN4zHxO4eRn/q
GXha+vctfYFT5gmEC2g9GmyIVRcXdrMHqCpHI1zrAr9aHFTLrMGMxUS4F9o+bfIoc4xBpNaxb0Ge
jUxWe7gQZ6GaPtb7m8xTX9wRD9cgEjHHBG0KwTwla/Fqz67ZDIyO+kuMJT7Q4SXjHunA3T+Irtes
80hxIIjcmpsKCLnbCIOJOWS0ONR5cKsYrNZkk1einO2gd/suH5JnFpvzI6uLN18SYv47CLymtHAk
Cs5CkvWuhwgJEUUyp+tpnq8tYXCvrcDGIw0CnuVVFJUcik0wB6cQua9KCVI1BP8ViC149ba6w7Ha
1MYC/UMFj5hsGG+DMGuYN4S7XyxnXlo8AHUhV0CITeObvM1Axs5kyHSTuHg58O8ibEHkYLi9sl6I
Cb01PCK2juNuhEc3XB3m/kPsn3oprHVMJ9ph9H04H6eMjk8+BOpsEvZbnFCB8kYJdbVLlWnAjNVg
aS35WtONQD9CU4NuaC+Yn6LOu7D38sZX0IeOX2VP+ywzOcGI6yNfdZWH3GFmpY8Js/gTkTN1x4SZ
xSLbF0Re4YD6Z1RPIo7Ge3LjVxFT00G9WODe+qZ5EMoEHV4x/Y4pZajEQdaKgYkywrEAky0gYy5w
kLynuJ/eyqdNmSBNk2UtIPhKonnf3KeDZH0U2er6TbjTM+mhkpzU5qnoxL5RAfDlRv1jci8zaISW
3fiq3PXL86Xwi5uv6ZxdL5oqUhhuYMx6dSuUrKsIMn8/qThxTlOkhxocjWbCHblUtCylIK8aOf87
SL6ZgmMbcSQvyNmJwKxJj/+DhIy7M049AssxTree/LbQ8j7NIP/VamsZsjhSwyN01x6tW5LW8s1C
cWvZPlQTqQ7Zu3u/H/+4qXS0qLFww4zDVNEIhnCQUsFqCu23A02ZTpiVfM+4vquuGNqe2XZLEfa1
RNTripAI6u48HcdnYEdu9l4u8h1xOStp+cSkfHRScQr2nzQzQRzC0gAZ3JPM+hcjUmRK+DwzkqUu
CXQjHBezvB51Q8DgO/PJqZG7XlK5+uQ78D62JKH9ST0EWK7CnkSC+TDD7WPqVpg8IQfqg8hUoZ96
zBD+FfuRR0hNeuU/QUSzMpX2L58qocrcHc1JrkNEGeuLdDePS8UBMaAklc/2p30SQq15aMHKASaj
h7Kwfubo1Ul4uPtfDPoNyablNHTiExCM0/yMxp5TWiH4TcQctYnu61NruCkDkA+/Hnn5BzsFePeX
WJwmFi5bPBTMl9Lwy065T0As5tifay2aDnUSZUnj97LSmUxdEiDrySIWZ5Ucrto8bN0b984smYbp
v2rfF0FgPBXTpXN0VE1xfDgXihvcGTmA4TTPUlfLVW06Ut88djo1edBOv5yNOZblH3l/Pln4BG02
dwmu9l29knNNVlwZYaDqGEH7lGgdsJV2X9uLAIBDsta+IbujTf6odW+Ph0unGdreb84OKVjmRjUB
SUQ9y02wvnk0qspzblnnOpW36E572f4zf8xCi9SgwOi3zrM0rTNFlAM731HqKir8OYxTQ+4rVgXh
ehx3BV/XHUAsoTjE98tWlSvi5SLFyrJAurNZefVgYsjRQiMpnB33LmuR6IVdJJylLx7q22ueENBS
X5kIUAo256TAfELzp3V1GSvIJ+qv9ZdXLCAtOHd2KBLWAIQj8iBH7alWdvH7/i5lTEtN76hz1SWu
PpMYtPLIBj+zMbb2/ab2pifIfchpoekq48KCyL27MMkoa9UFAsrK3NVRx3ob4TwATrB/zttPtBbs
c75Ro/c61yAfAcKxwwARZbpCQhKLudKk5N4Rr1yXO3UZIUdePKDJD/u/e7F/IHyCn/NbVQwlu4Wn
nIivIBmCIgnQBvb2flDzy308x+xNHvuI0H7EZvVtaZvYOV9hjLsLuhEYBwtdjoQIf43A3a/FN4tF
9BA7QEZQsKkRIuTKB8B6Sdv9TU0djYIKsWuqtJ2aWfBhI36AfWGUuUzQ3wzi/xLjcE9vXP1xkwg7
I87V7o9gzU+BmZS9U6l2/CJ5JJuVWbDPRIvTX1c6WAqPWXyVPebh7fNlqiZvwu0IGK+ZXF2YzV7Y
4mv1SwQp3PdTArEU+BE42X3TQBjE52qS3OeT4MWBsAILegJjJTclRA7hAITWVjKNY5iW+GjDtb5F
oxuTiUkJQfaR7AZ2D0dNjeiIRH/ZT7Cd9Ti53raJxN2m8u7sWDopGTHAIV7v1c+uSRV/7yA5emxB
Yjg5jTb2hK0DfBrduL+7PI/8MEFi9h2k9i3iV+nIedEZsLS6h0bhIKYZxrM17yaXhP7yBxInRMDX
9RqiV6MwHtUveWFXlfD6bo96nrw76tZnTFCgZR+ZHr1E5Xzj0y/QTe9AoQprwv+0yWAF9B9DH3lM
c27eh4cHQOik7a8hp2I0uBf4h/VH5In8fZ3ya3pcPfMC+S+rfBCDMeRDsurAG9y4nXnb5Qxp+oo0
GNM+aezkNoVnsmwPxE3yecHXjrUSgvi55RdbTlZx+ktjLQ+TrXsgAVaS6W99u8l0IbaIXqzQQSzq
SwLv/gC3sEX0H4F3CfO+8/evSZfxq0XTt/WTB8esun4be0JeJy7xBiNh4My8CBlrTDd8k1UXbMVT
6AQh6AuvYfLGfu5wehU8UyMVrA4iOkwOZvA/wm2MvGNSgpUIE8YwNG0eH9y3z0MQUxPrWU9QAA98
dexXrdz+ZI2rTzrKACNUV/Js/2HA2SIFZgT5qsMyL5+jq5/iwDQvDLcwFxMVZYcZoEQthJvhFv4y
TmK5KWVYhc8LPl/1Sbug+1Ot51x9pXMNDw82hpWECnAmF+mQ15OYnLW8lSUsJ8q+bh4BHpzl/KFr
4k6KboRJVFWwAHaXnbCQDce4/DlinGO9gsx36Ev+wlybUjmzI7jzMAkhUk4KVoAksRrj7uco3aIQ
CaALQvuSxLJosIgtk4elkjeYSxQArS3Ai8zqjuej62nJgz6zxXUMTrZbKBkwAFkE1qwKvkGF66wq
pm+gm3Fa1UF8oygw9UbPaAiYpMUMbqmZO1TJ9fREhHRt7+yh8+1bGnXUbi7gYbj4eiUj+0+viZyF
j95WnKBk7edix5EthCsLg0slt3pWUdPVILBbWviv8ituSfmYbqCZ+I1nsAoy2EUZfMvQhprzbEXo
qt6EaPgLmZrbE2qeuRzzAim2PaZoOkIYDJHgGL4hKEsqPKG4fvFS9zemDpewMAV8GSuh8Kbq/8/J
sr7H0Kw+YanRSucJzYb+uPDrC7RS2eQOv7WZqZVSa95vLRxLFPrOQzqn11LHKfoKWQL4dF/Vrjxw
0il6qDyn9HMA+rQUaAv8TvxypAiIOINvP6ezNY7zLWLcQau1Wm1OCO9OxvRg0P9Ry9BBi6NgSAt5
qrOKePf+dn8v2CcIRLzXNS/eprxeE7nVdboLMm6ZU5iWe2b2heaY4CfstmIVWVnZDPusZImjyKW5
OmbujWWbStDpA6XHcmnnvPF+Z9UWEDwUKSfHeLuTmWwOpg0uUc/b6iR+6Y5T0FVBkI9BIRxoRBtB
bOHXov6AfYA/XVeD09sUpQWQp9I0jrKJDB+T+C0PdHcgl83SQKDfqfy6HXl593AI34KSRJa0tnjc
eI7sJv+eGmNAzvaeDpQRL4iyO79V04lsCbLyo9lMdRtF6eTZxhw6iwPEu8RZYyHuhzruZ7Dbwbh2
S1y8JMISfuCps8svoqkFNQQ/6eG6P7DOzI7VDkgHGPIrq8HO6CPOhAqBpKA2IuGxXljSZiLLaZ9h
JVNzFDT38ONXkhW0dupWyeyOkz4qBjn6D1kbLRaqP74tJXoFoc/i0RKa3T+nPbbIV3NeR9UuqkDJ
lY+Hg/j+amsVMY2uuMyD1cS35MRXD5CsYo2aVRgk7RRFgegsbH6aVEgjTkana6EVaMNf1WFX6yx9
GBkmNtFqfMS+jgWcomRdb/dtLGL6u+PaCqIjxMR2bAN3gT4f/A+SZrH5gDvoXW7o0ZUwh07v2dZ5
D1YnmonANrzi4k5rAh7Lkh/IJkasia16lbeMDIL4nEw/2ZJdEf1byJmzCc2EQ6HaFslgGfuPXMi+
RuEWDkxSPsutw7dDZGTrkWYtQszLgQ5v2Mm2c2rrlx/oneFid0DU+lZKtm7Gk0KgH/Uw888ld7oB
z+dWc2Ca8URXFyoP/ew/z3L+HBvgwP8X0b0pHRr2Xt07gFwPMyxg0D/wyqpDPVG75AWk5C2W8z6w
aJ04p4i9SPW0xvIK+Krb4H9+A9kcElA8k490Cp0g+jwdSzOcMbf/hN2bdAxozz8xC1r2qUQOwoQh
+BLTQh1U+TDnKYXRz8HCg15shC21PQb98XGGNFHdsC8L3e4KLNa9ymkl7z/rSRLErQTF1d4w2y+2
IKZv/cgYLTMvyzraTwKPvH3bPJPIv05zyXAFhPmtM1ShRuqGr2XvxooFeQsBRqO3vUq2lFISMXJ0
bHgBKfacEawozcHaQi5+yQtUPlePtnviAbWBIY+GGdIxLk8+hdsKeQmEgghPRNYmPEml3Az8pA4M
EDyxoOUTCM1L1c7U5lh70tGsyH29Yd0TMCpDZOKfFPkLdX0veF0OxkWOL+AlxsmMZIqq7sZNQQLp
HwP3/0JAzMj/IIGi+Yq5T3kkIQGBUVInjB2ue7PDeQUvrYlghE3GFyIWqKS5E+ky84NdVhydjBDT
Z6ZCyxJE7OnA+bA83jX9lVs91ik8Rhr623C/Yxe+tM3OC6bEuW4NsAwJWr1QauxNqRYinaO4vRjD
x5Xjh1yDthoWBYR0PUl46SF3d/VsnZ/X22OgSlMuVCya+eS0uHBNxx6QhGyoQew5shwwcyM9kzXG
L3rnpe/sSnGLbFRf2T/wQl+WNQd7PiyXwfwPQSJQeflL6YFgYVM9Q4mt9zqwIqgNTYHmBA9bFwxR
UScI6a8kSMr6uio84oD2ujunYvqE7vtRwxntkAftf4llk2uwAsrlwBoParA3iYeDqTIcSSBKTjgr
qB4Fa51ZHWAJtDHM4rXu9a7DseogyxE4R8F5rbBZ/FZmAfRItLqMcx5cnWpAKtprFIs+bBxkR88P
Hg3vwshHgied7sTmVecpYYM918lE+RLioe3Kx6ufbV6XylheZZKfPOMkrvhkQDcI5SqSvnY5QZqs
NFuzI6FVSCfqwieDQVWW4E5VZma8/q8Q8pL1mJp/NokdnF6M+6YlffFzzUx3Ht22jeLeAAJF7H5Z
/aATMkpUL8aA4h8zAgD2OJqtAYheLvShqd3Mws+FwH+4t7Yfv/XpfiXY35toR41rO1Ca/CUofj1U
/0JjTBZOUxtrj5dbzPpF/Tc3aJ0NHQNxSN4g8F3zkz3L20qtwLBMgEDu+69OSZ3FY86Kjg078kzT
/u06iZjX4x4um84MfGfszZpgx9u1B2R7U/henHiIPdIvXv5q932OGoLa3FVf/wrfL7LQn8jfj4zf
3MvRl8w//6sjzM+It5QjYH2gPYPyIUh0gIgDp4C9UKJuYHTeFcyhx3YXm+VL3mRQ670Yq6kTHDXq
hYW2RLc1ID0hspJmU3m6Cgj42AJR5z5R5g6EaIILBzpq8oWvwIKFFFdwVIvxZncklgx0LHbzU1xm
OgGQcwDvqCbJOlnn9+5lYWTtI/sSEWV07LCEs5UjqfED5s2oAkgjyotMGLyc1+5boRvgOssItc5I
ejqY27HN2xCu7j1wo3YNg6tW2dWtsRADZkt19hfM2ZupQCFvDSpxCtL/kbmRzKeLY788b9nu3Gzt
17zPej41oliEVXZfzVyHDjPWUg/qX8IsWhyy0DAOkfULutx3hiUrBA3aJT4o3b45950G4b6CcKua
3gpAWKEVlbai1VfitbZ/jxYXfLZuGwjy+lcDukCMr1dYnsMJG1L0xFd6jon1a6VKvISP/0sGcDib
Q/7Guqwo7nuSjR4n9+GO0d0r/tUDO9TtCZ5+NYYhe/1lg1WlR+rk1otoNIOUKwiSoj+r+UHBIbJ8
fSo7wQjsYmNyE4NvrQt1oqT+9bmDr07Q6YB1oZMRsje3eJk2sZ1mNABlTNv3kW1tT9vXf6PEf+Lj
S24Hq4iNQGq3Vnyt5reNO9X/2lm/hfpr8MVPgHm8usUz76VzdXO45pkes3XCM7s9oX5WOacYZw/J
ulGzgDShdcIcwlUCzHQmxAwovLB7WgODChT9PpvtzyWqAgkU03IZkkd7Rfc5cgwDmBX8Grg27SPf
zhzkNs1Jf848JVYobu1haiOUz6207rKX2nxr1vz1PgXqAM62tIeSwEvHE38KsjKLlcpN+AiuKFXE
CbHZPl5rfwDpRrzQlZaILWHc83X856dBtXIRNlGlgD0+hBQ7npBz5Za2LmMVw7Y5pkkV5C0nqn2P
YwzrkgR13wIC1oLGu0zQGgpti9S7zC4ESNw/2TKxcKER58M5qTQX4ROCIHP3G7uOAGDgoIYslSjo
426cYSAKHXRzZX263O/Q6iD2fCNPhIOpGa7K39++/MAsl7SN3IqKuNxuhr4ejVj2s+1ldi2vIYbN
sk0GDcnZNk6u7V/Gm6sutrTgcau0QrRH7T2MDKtltBBasF+sWkaPdcMzfts8MXkXDXpc8FglKh6s
E7KkstP4OuHEym36+WX06aag5W0caoggpGtdmnjYuqB9AVLr4tKdY5lYjb3QTlArtuwiVt9Foimy
gB4WAuu72t1u6IqyCa2K6UYknN+sCBkbcSC6ny4QducBxh0NG2y6b3IuL/5JjB4ac8Kc6vjg8AO3
Q+N8m56EOMQhCVXrtZmKpEKiLvvSYYUu6firQe5F9iYha4dxqwnDA6ZUVZaslYHwLUBnmzJC4meF
rfZb6cT4KOvkGjnO/9yIUPIczqcAqUWdTS7LZkgyuZMqQ9tFlpjx/A0tn0ieq6dzzT0bC5zBvwle
JVpyQBMJaveTxem0TU9CVwD6ysDKK/axRVGjVW0DPjrwAttVfbmNnuldTsfGXzjiP1XVSOQakyaX
QA0dvzb0zNka+SeIVFmP+fOtb6cQHPo8TFAt6BRkEjtKahGJFIaABtUZcpUEfaZxzMikpbbQEari
anxRQHnvB+81DzE+N/CN6Edh13YjSUk2UuBEPb4tsr5nUb7u45X2rrA1D1oNWlta0+uFeJ+Thkzo
0yCI8cejKgz/BRhOktgn5zd3chucrndZ2CId1R74SlDVGho68osB+IcZvGJsODoZlJF8tO4L9gOS
sw+7FzE1Vj4nLJqLVRViPtzSTGf0A4HiKZGPSxFBUYepxePHEhKa+VZ1Oa09tqEx0cISZSl9vfhG
c+sr7k3FgpbIJihrMRutTnMytId07ErReQfQlZ6VEzCzOLQMa7FEZU8sbkHt0pQOYDVooP0sYrdV
1QpXnxQ/BKTdCW0Ljdhbja7YC+1TKn9CJosuuCGqOr7/Tu4McEH9pIAX3IawwjXr4hl6FOi5pY0J
M8OkPDmvbjBT1fB3onWtOIuFyGLIDLWHMbZpdoK+SJRZ/zYt+hm/Gr027V3hIvrRGBdlJaloqrvh
oj6QdJ1ALYqw0AEsf0JcGqeVW5+Z9f3jAZ857axieSGxZQErcrXNg/1S8pdvgOou0b/3HpEM4N2r
hvp+jz3wDJZxJ3s7rjPr5ZTMUypqLdE+9IPeIWXG460WZiKIcLq4wIrP4HexSLDVZe5XyLbM/lqU
xTQU60Ksd9P1XqsphbXslBtSnxwlNFSLZYTMp2xIR4A2aXWpPRAEx+WtfYUQ6X+l7HuCrv6U2G2X
otcpKE9uNFUnQvZL+wrFkMXp3z05TaU5ITBXIinZartqrpdkylxIY1a2n2vL0LJgLDX1xwqPJTUC
nGh5YLCPn3Kc0FrkUHkKHnj1hPhcPBrWHOfDchyW8ciM3EWHNIM9Mjtd1Tp0b8BPTa046WN3iEeR
f/W9Do2iFxn3jRGlEbOL6eT6/Gj4E4m8/uqzlUOLSp2yut05CAgofLbJmGIw1sEW4oQK5M5Myf3x
Yl/GAY35lZ+w6qARRmacjwb15CGfVV4hZErJUCTsCvvmqV1wXSIHFtmJD7cdDriW47aUUd/9wA5d
UsUZJ/aSUwzTgyEFf/yLd0rrBLVni0QFzGSeI1B/ilDXPD+J/W6fHut5odQy4xwmEZzMS8wM0o8k
dxKHkV+0MVqJF/+c1xEAt1jCLx9KNu78jJWThcyvqk9gdbxzi73ORMvBA5dsmX30K1MQtdLNHX/Z
rIjul924Dcp+rzxooegQVR/Q7DEnYyhMifwRR7h34My4a/DQow1Rhe9ZT6nZuWiKuZfjk1+P+C8i
NoOg78H3X+j9ZsVQ2AxbRaKcBymkm2wOW3hq2s53Oa88GUOSf1QHKwo7rXTImOX7ZDJ1jxxiTjio
xGWlnm/hNJpIER5Pk7dteavQD2VWIDcRkzcJP1VITB3HC0+hGDWhzpiVySJzdwwST7lpfCSttms5
ORQaUCJjodFR/nG4HQ3h2ErcUMw3JP3HDx/KdMbMMkUb0tucRXAqJzzlhBFB+VSy5zaP+xHL0co5
eTe0Xn1DOJijsABNTslIIeq0LVGXCtybd/Ju6S7TcJgJiI5pOq/2H9Mvqbi8ajxBxGRX6W0MncXe
H3qNs4vC+D69GGBSVfv8ef0QMmYbPUpktEg5/KISLxrEHdPC+q4Qj0QG8TUY+fLWwjDnkBnVTMmu
YNaEm3k25CQTvc4U+GWY/7CyXnaDIDBLvQoDKhytic0wx1+MNkhH/wHrp0Jv+B876zyjdVYeYBdz
EoBWpBtaJC9pXwj1JeWUC5pzbOsXzs2cNEmBBSFkuJYbelUpHDC4EM3P/iTMOLc1DnGMjx93RDrp
GTrEpKtVBBqglZuwy3312dVcBA0s+WPf+onvgsKB9bqXHPBfDv+3D11mkuKkGBKLY5YdnQXzhZ3j
CAZo0yFjxHGu395OxUh/OUaxm7qfqA1IPq1YlD1mC0tVWI5mERuMSwiKvgWZ166UZgsd/EZvBNKw
lq4mE9PsOuyoK+SYR2W03lxR7ZZGfDWF6IRvZe1hkmrIsIgRzuSTeYx2HGX3UsyYb1YEwDzHLqJL
MA1D2LuR9lXT50ugx7A+Ot2jr1ZOoLcIU97Wx8VhQFe3zDzgqKilmdD5OMEgABcIaz6cTMVKsrov
MZVSJkpl3qGQwuuqj8+ieaHbk8lAOG0XpsKEsjgn7rir2peC1eJHe1mF8zSvWlewaxyST0SzPh+A
7kK3jnpALx2170ANVRhnOY68bAUAylbmSAAKxMKkp/0bZop+8Wzp3D+ZkxDLob+nXftjIOGufH2+
Xylu8WsWyFrPZfJoV0WbOiEr+pgD5ut5BUiSoL2ciVZjZtXWFGa0INqaJHiDnNebUnBRNE3JmBkh
dK4vp+wHVZuK2BHxvo3zD2hkXLoSg+mtiv3HJgbb0EG8fQe8saHq1YYpxWl6hqjESFbCpod0H/y+
Bu9Evrhw0S9JJdcIrDpsdeSjqG2aRVUTbSxJ6UXxefBTf2vRG8/ayBTsyOBR8dEAsWPtC/SKAXY2
j7Mx9mKuMbLjK2xhpRE+fm4wFFZ4yQaloWKdwSt9w1O/Y4ZYoi3c/eJ1t8m+f2YFRcnkYmuqKgiv
PFseN3qXRp6LOpaiq6sx8l2b0MDXPGaf/vjr2oFTserw9qB+I/BuRmLzru2yqrx0hbOzoiuBKTej
T378jTnOr9pqrtjPJ5q6y4i4Oh/ZuSOzj4UHF6biUMpls70J9y30ad1x3KswIfwiK4Z0sRKOhYim
vLgKiZ29n6ajYbDTZpYEM0au2cwG6S65KczXx8uU1TmI1NMU69Q6Zqi/LmkZu2oRyxY4U/BCdRrj
Ot0sM3iKlM6A01sZkDe8ish5krBdVxPWyehlu5sIffBaAklsYRt/F1P0wMb7ZjpfPqo6OoRFwS2t
06DzrQzg4jSzE10yvD9fh8HC9J12lRzXbrTtXslKboeMvHa8E/y5WDaD+pE4kkbt+WE5tfKJ+0jU
70vYkI43Q89h2jta2UkQNVmZoChB2uj1BEdiaz8XiCl6PB1+Bkxj8JD6YLw1Grf6PWGI9KjhU92A
dE3iu1cYLXxVn+CXMOdkV4bVBLOjUEt8TWUW6Inw9X5O7ldTkghjwl4amEIFtWah3x2YumZ4qYna
IJQCPiJY1g+9Y2bTC8P7mKScNzZjuzO/xdN/iFeJjRiaw5vvGdXlE+hZ3jGiV4c32ZVIu8OMfJc9
6IV5qtH3cU5BfQGsdwmMjsG76empWyI7gHcOja+F8QLyqCd+5HhcUrkrY6qxss8u+qgzQzct94tn
zTC6InIvgSWjo0REYJdyCh2qEYoQXuxGkUpyXbP5Q1aa6KL89pDVWWJXGZ8T8B6tgRVOam5hzuzB
nvh2aSv9+R7sMnsyqVEl6+A1aOnA1/Ff2P6GdLjEFPwK/Y7poBpmJUHA19Bgx2QA/dhs9Xse4RLx
ghSBmwwoDPVo7ZweH58qDyfcZ78bGDA/eBAYx2r7kz7FNw+zytfhKHWKcNL/XqFo8O+U5p5ir033
qs7DruQtuOYqJH/oIi1CuWAkhqDfU0njry+IKchIK56UwI/bnWM3nYl1on7kkLO9Khfe9kUzVYFZ
ZtglYm402EYBEYnUTbbElWwrbTI7FxbQZXyRFob5fvk7mFw9yIninEoVQMmlLjmwUbYMZjZAEz+S
R9gWuNuFonijS9S5gz6pU6ti/4sHIG2NkME0dhTAp498cwqcfD55pzU2kmUMBaMPPPL4OhclMvac
KbwENM+acn3GM9dvHrWQg92ES45ZNlzBElXraS1TzlOakdWQjlPm2IgOVBGI9f0n0d7P4O8+BSsJ
ToKYd0t0L01kMqVxuK5xdy5m+SvOpDbdPLNgkagRzUUCK1nruWzE/FNo8ybxLh+WERmF+uSMCd0E
XAX2vXMqGGLZP2LMcnGsAEH/CrKVA2769fJkzOGn+z15TzMNc0km4enuwGDWB5OSLjbp2yUHKzb/
FUepPPhZQnM32W+ek4ciJpAqd9jigMFtSo93gpWlIvecRKC6CP73NrZHdI0d0sCs0Vm/9Nfu5nGB
szjXGIX/Bp1z/zMRg37syywXinTPuTobZmzVIXeZabxphl/FqnymuA0Kqx6rMmZ8PM9oEjxg0KVU
N+uklhzkTyROUdeH0J4BgefuMDcS17mSVyCI+OD5a3++s2R8V7MDuH+ppJAAmyeHnk7QrIhRFTVX
Jdga2FvQIX8hBDToQ7jby5ubtm3kDsi9f9Dh1IPl+RLi4PfWFgLr8t/4gErAHG3ZvgFSsB5vyJ/y
LDwcfHBY4b5J4hLxVbRY5MVgD1hLfabvvKxPGOXvJUtY39ngNImx1wcLT6ql/1DNQinsHFjC96fR
HSScxvf8mJbYjxUGXNmf1lZSGNvoD5/LSat4KDujo/w/x98mX3Ex5+im+N0uVa69g80B3O62+ldm
VZF6ybfYaqti1O+foslri2cB7+WbkDPPXluadXxu5reUk5Pj1D9jqd1/T9c84YJCLMUWWG6AmYma
VRnIjfGtxOas951gDa4qX5dp1amg32kfk+hXm9IQ7icXgH26BixWmXGOm0wB1HwvPKKJyDuL1XP8
FuZlSmne+nqeykQdWZblAvhTb0QZWLl0W5bBzNivFMwIWJgSPdI5lI8JrVzF21XxBIn5QP5SEv7y
MeMvruGkGvuVV+v9gCHXTesoZr9GYZ7q67tTOsW6AizX5x5RFHGIQL3YXZOTYuPxbg+9Vj8K5MSG
NcLxPJMx6bVaIcEf0Ho27QL6ltz5IxIaE4urOGT3EUeJWFzllx1wWyLhMekMDMhDE0/r32FIgt3v
4EGb3c6FTPMRRnfwjTJiWo59CRD0zh8h23oa+iQzw2KFRp/E2VMRtJSDAIlHFho5x3fXPC/2gKIM
M7PYbpf/tXyJze1oqCwFOBFJj09NmhulCRIlILO9F4ugIQn+oac1aHlPnTqtzhRdPYgrFpl974wX
mE3PFizo+bPQJWExK3Ga5xArog1qII5mFxXPC1ZaYwXSPY9diMf3vcXnQIbocO4bmzyLcsbK+Wg0
3Fc6FxR5Y4sX5Du94u4Mqwz7vpCYPWT/0mpG+B9nsyM6N7mOCDMA79a5CyFKsSH/0nGsbSbgXOem
IbuOsOJT7iFl3Oke0o89eiaMSM2jS8hxOPSpE4vZDaN8gukwQSY1tGo67amJ9C3EUpdt7+eOhcEz
Z2L0WLW5t9bjQ4bA80IEY3q3foKlLbmp9CBDf5HeyFtmjG07T7GC8HzXnrE063oqzKO2PYV3gWqK
G4e1UTef7hm40PQl4zBqY27ZJAeFhG8dg9n9HWK2NSbfVGoeAS9jyc678zRAA44W7MFvjnu0dYH1
/fFalhIR2CZ23a3w97EfROMPS8UkYcu9gJj9B/3/ZGdC0DEvENUGuGNNbg6overUV8H0XXAghGRw
fva6avBZtG5QDBJtjRU/mDDUtwJiX4HOysFYwNGxd7mWo111OI9L3ZHtVuqUGtkYs4UNmh1y1cdh
DLI0ChZGMDOqQnvKx96lKCkmPznhQl63JU5Su58Qt5tQ4c3JUx28rSbVlNfy2ZA8D/R2U/GKLwoc
fQEor4V1RQ/5XwFLh2eEiucKCij/cFlmSAf5BlEkmhJ9VoxkdQcJ0qYZHZbRxESe5rRwxDMocb2e
kuXKQ997BVIc8snEaPVa7cCNDusmWvUwfit+rQrxh4d3xtsIwh84o1kz+ClPtnmcpOp5C8fxg4VJ
enGxZf1Mie0x54TmS18gZvIFBzrZ2K0IdEhC0U54UM9EL+sJqROsiLMADGF71w7SWI+8MaPbx+R+
6MTvhgRm+LfS8wCdseLg17t28+8Vena60NFXfkA4+o5mMonKJBseY+zmSBQP81BTDjRolrJY7XEr
CuBdULDh/HwsOjKQr2biP+RvPYyrioXdK3cvEyAjEmd5klY/gt5hKs2c1tHZT41Pm6KxsHwxM6YA
LDD1mbTqJ/beEEYZHyrqg3aiF9iS86DGqi+S8IhB2pDuJr0EXidEttDGD1MthKGq+6ydhMH1TsAU
UMZ0uCrUPhH5eQEFzty/S/fpfh6xfR09FzWAN96kE70kqf7HJKH0ViPxuYS0z6v4OvKBYqXri+KK
CrhWvqTmXDo8Wzw6MNsQh5nqgxqg5y+ZZiNqnrOVbsYYReCUfCF73YkaOxWApsWZ3+hfX6nyC4UP
gA1mb84Ud3jIepejlV+ivZJ5JZd69D3g7zStXxLyzUqtH7vBC+MkWTh3rL6KSqcr7Z9Rr/nADnFW
Gis2GMTrP6DKOx4pnXkD11akX8fIM1F11+J4WIWbTkr8P+SpGWONr5ZTegr59lj37KAq7lmfKDjw
DeLU0BDzLf2vmsL/IkGa08fxQDSmfKBqupN8DXyNK/0EyF8ZnnSUYak0g/7Zji+vQuTHIGz53iLZ
2UKHbJpdhbVG8J1VqdFkrEuMcLqLpgj/vg2SJSBokh6Rxb6+LcRAn41RYkWU71hL/e1xpcnx2CGZ
5LDQ2zXs9lXTz5egulRZnf7jNbral5gb6d1cooYnEZtHbTYTWSZmPr7QgmODdjys51D8M7zxjejq
zxcRdahgFIb3/ay/ze4e561AHrC2PAl2DvauZz1S4xpmk52wWHeL+Y0OxUjIQe1DnkDY7N7mUBJc
ixJ9xw0qB3uay98g/miquuzaadAbcmEiz98gmCJDprjSShFLan+Qik/ir7a5HHgx9N9JV5V7lnRd
vv+Ik6GDXkcLZ7XnLfKL00ezajzVM6HxahSVf8ZeOwdobFEpoywWWsNT3r18lBrZhqQ/uPZ+JJ5N
C7W5q6xPNuhdSFZoD1/T1bn/efhQ0vyIb95/XVH55tVLUiLy6lu/Hwc6sFpB3ElgR4Cl9jByxx+M
9/08fgk1SIM53SnBkD2UPqgmV/Oc1ft7D34BkBGXv4paP3Bcmv4BHOaH4/Ap+u22Kd/3CzwriKIy
TGIer735fQ3v5h5vUosSM0W1mYE7ciX1Og13Pwaciq+6+IafpOhJAs7bi00U4C1SOtIlwpc6rNuD
VCw7+oKokDXmZr6NId3/HThMwC/TF/Ft8NvexkOQkvudHgtrExK2nhl5kC9ZEZ5grBqZxUQ6zM9T
0ML21hOsMkC8K4D+orOMg8jwhEMjQkTcz+nLuOwjVhoji6+GjU4NY2X5TCVaVB0izPKb2W1mVL83
Ko/rC1wYhpdvaagrHKgCfwOW8A7c9M5NHHX6VMg1a+0ihphdVLER3t1IDuZdaZ2yrxCT1RfOXOuD
iVOGz1BZklc0UJytJMv0Loziz4Eq+iabMOPdSg8xPWUgjDxDO260qIujoUOkI3mK7VBI1LK/Ek57
1kxmMBplabCxgQnuYLgEQYJbz51is+FiFd1AgsnQPdyEOrsh/LbbKd5oKXYRSXZdxPj5k65grfPp
AApqWC+U1Ln6lv28bZHqDLcgjZBZy5JMJKV6wcGDFBCMkILI3m9W4DNwGoOarLJNtyVTUbH1RuBX
bfQbR4JHcw3FKDYv5MI/T69fdKTalnFkf0zEMEgHp8PqXUPui72Hj0aNdmLcfA79BrsxqBr9D39N
hq8FT4T0mU5s7K2To0zcyGW4irE2uzTexoJhmIWwQ0KiIIV0zptkWhDJGPUWrFifW1Vb3AoBZjxq
51EcanOVZ9yRtNZ5+DVJUq/4fhKjN2k+VySKwG8P4r79zst1fySKlmsd8riXhWePU4pc4/IMm2HB
uYTVqLLRMv8+YVc2W+jymtbetyFm75H0kYs/J21eQvAno+NB9l5wsI/U+gTBMAT8+OIXMapu3L0L
++hxgKIqgcGRi6TvzvBNa1vYUbu11cSkqLx23Bf3cZJyXaRdFPsrZLIvb84ftXCGnNr+yb+GxPMa
8Vxnul4LS0kN4kI0uukqKRL5fyVdNxwx6ePHjQcsyUBKEnRfun9gLmDrhWaleZLSuYSC/u8Sp+KB
EybfHvk6ktmkvL0lLkXNse0gLCdSWk31wRyTPF09oPaSYKJbuvf3Ljvlud0CZ4acejP/ddMiWvBz
7CcUFwZ8beuJpp+YhvZPpLv22E+qBkhpJ/scKCICIEh29zLlQ7/r6W7Wrb6pNgHbWJOz0AaJo9qP
9E2L56URCzzxEZZQSl7hwQZfkNT+DpI88RriuHWlsYSr3YFXCpYzRw2MTBYRsywSpLUxNl0aJVh4
0FM94M7TrSXK+DWtxgqOdG2qdh23+N06Yf2ZnzlsuLatyRn/5nK2X0B1LeyktYYy8qZT6JcxKhps
C8UX279TUVf3LDJjDACio1XRsMaOC4W5eKQs+qWEgqvI6t+kze3sYo/wix841Ae5K5FgwoZ3HuLr
m4G8FjyD4mEVt2D9VGh6/hY0ycA4wje8fb3oOEtLRaQn6lheJPnTB9mYBXDJaqoKDeZob3r2ralW
5CFbtDBgDeJU83bqVx15HnAnRs/cAFufusqUoA28Z7+rB3qS7Bi/5YCEe+uHprsSTbpOdUA+g+BO
X974YqtJppKtlD0hT/g9lC/V/4IkxFifKcBXueuTXenud5yg04d8hvnZQQM27MFIfb3EahnvQ9dO
0Nw73vuCU0WMTt6y8KeN4VzJuGQslfbdeErLmian6gEspQR64UrMfKvfDQK4S3woXYs53DxGhg+5
btOMOZYsrPOv3J0Ofs27HXi6isXXnestkT/7Q29VOeMRJ/pjmN8yU1GSuucLFpxB+RxQXtxYMibO
wlm2lbhJ3QwXzqFUU0UHjVoYRJn0zBCl+lvV37y2R1r1xdGIpWTElzrjc49Xu1U8lZax1+acYEaU
NIJrpw78aAXjndiJkmHGoCMtvUG7AIK2cY8tiZmwJOBBv4prCM7AR8ZA9Yb9fFrICATLXk1j3PIx
Ryofg84yv9Hxyu28s8j+R3mThIQbIbkhYyRoDUNF7azIFhcCyczek1ZWfnd6SDbFnZeOwCTMPerr
cP9YbtHGEwAtWlRFJjt2CDVmRwF46fQTBhXf4ufzfGYeoG6K40lGhkqu4SSedePBgZ7C0CtvPrJj
y89y4Fn52l7AOaKU+UMRaG4PxGbuzkaupV9CPvyhWG6MmMC4fsOdu6C7RHIceNK5tn2YlLb3f3Jv
qzwkbTjxw5rTvJkUd6KVmp0Ld6gZ1xHBNbaOks0E3DEO1W1IHtB1dw5uYHvv1KmnMba/PU69mkQB
gSg8dxqRMlExRHQliKIHgJCNtyBrUNEGjdiy2TGtvkOOOtCbVIMGca6lDWmqZE51WkF97AeTuRm4
XVX9BBnYP3KC5szkC+Yc8+LePE3fVXmynCuOoCgzlINdCqv2BQsb5ZXIJsbiUeJ48L72BPL6B8B2
DLL2cK9OPnGR1fwfW9OF//ZrsO7TjCh/hbtGsQbGFPKwLaHShCb4/p3vheIVO24fnoHiwqOC5ZBF
1iMnGjIWZmm6S9I2WHi106Neeqvpj5o/RZruQQkjRdQbuMQ/Mej1rVUsw7vI26j6OQ8p22RC+diw
1XDQfEM4T2ZhLfskufgPGnj25p4NwLtWT/GOTgyxGQf7pGvFKiGa4rvE665IrCkgci/u5cv6WVhQ
YbOI0bx8gN3+kSKFQfnm+9pSKHTkaTIYcc2B3NIFXjwtGfy4sAYQ0FQceeDT9Bf0MwwDcknP+dvU
mVw5lm+mko4RvtxDT5nhOn7ab14Wi4dzGBV23jwckN5ZGVq6yAJ2EEAc5QFnS/yze450RwEcL+5E
8XVhnWanasDYrkb2D5UOQQQsaXRlP9PbdSARs7LXCXVXZg7HYXByqvTpGL0gOeFJxk4VUOwX81Af
3+LfzPy98utS+lvKpBbwaWkXmMCaINA8cYeTSqDYZ3QVuu6iF87eUR03eLVxYPDB1J5dBIIoOeqQ
ap/kkerJMUozylS+aicPLkGe2gK6IMXsn4jw22fY8I8dJDU1vUQGRSvtpIPLNKDfGxGXeuQ7Gx5v
zYx7cCi3+PfqGIv+UDzlTVQji1SZEOt+put7/LeNl3pHzkwXqR/nMmGXHPeRsPY+SZSiUOEq6X83
lXUgAPNtTzfyQkMYVZiK2g6j1MScDoWoonVrTcj3TxZKXPZLb6yc7VOZoGjTV3XRvJWHvwQwHrln
+f3Korf7aEuBLz8dMd8Ff4QFOpAVCK+Xl35MZacdJUMxqDVEJtle7xH7Fllsujhm7b7zIB8+Mz61
aKlGDYiwtLABH1nbPuFSyBy+GwXEzNrXUW9ejvquXJ7p+QYeH4huenT1asqL9m48eASOlJHrUwPT
EIC1z+3tV1Yb99UMHd/5A1KTlWzCJS2qVDkG7NUMRJXG8b+WIeYGjwPPzY4hSfbOrUJEvWC9AxyE
4JlWq2ez/1TcKiohMgpwHfmM0GQjve7gc8v9q7nLiZshrSSfBWwJtMAlGzSeSEVXVvJrgei/D9bM
g03lrDKrDqlugcGf3fFXAwi7l6AK3wCPsyqkWRR6yfq06RAFqPkMvReqJzIlSm+tAs+12xiHtPB4
1BD6lBplxKDXUW9UB6ga3AwFNdN5WjQ2y5KY3VjvNfFrRoRpYyYiQhg0Wcrnoh3RidJyI54z/hOh
GbSKoJQkKrRJdJKvpE4frYrB5PLGMF7h0k56aQN4zKqdo8h4OQthFcJbq9qbawKPZNrlzLou+2Ai
WyoVKTSDRZdxcyXd/wnvWXiZAWvBqNcOSgxi0tpLalrFWlO/fvzjb6SVhRggaAZ4ylAgRxRHbHd1
t4CDjV+v8iqHN6FLQwNJcaGkTj6Bn18XsRRIMEQ5XvwrGp7nPueMnNiHZOlHJu0wH9ZYML0oStNT
WzP36nhcI/eLd+X0hw3bNjzkG0md29qRZXN3Ij8PIHpwhRBp5nSr+bHRqdNYSVToYmxdgsxyX0WO
0yTiMpKomXS65Jx/FHTvZP9f8cP0FHo+XZrDyK0YrWmqcokbNGjVYMmpv9ccTr+9uO4BMaJb5ii4
/4IO8B2Eui/kOAcSCrZvEPQZxROhkRWFosqFAuPWT47RrwQuHTxF6SsY45ZeYfPIbumTSk9n8B2z
0Uf8VsEQw7aS6w6OT7eTRi8cSOBpAKEJKgWt25/JW1vr9svEms6mMdYZUndWVwOJosPTHfQW4mdl
D6MLfCaWdMb+dahr0sySGaOMxewq4Kr6hUNc0iZliaYcWNu0jEqxrk+ONiJclWnaWVvHQ++/OF8O
kb1XeYxS2xFOxsGArI5qIVVecZ9pgyLqHcHZbV7P4IWAyzIYsd6SqnFM3qcCPG+AumUjaoXLUHUR
yBmEsZqE6llzWhYaZ7HsNBEpXWvbTFwgJ8gTITNLCCH1FLtCU1ruidLKKuKL1wRgBNfJwmUEG3Kc
usLZ7Jw5jF4sCdhuPwumwny1yH/w4qiI1Lkly0VtuyICQkYuwBHYuRwXe22NroRnE3kRKBinioLD
+tf4sWtxo0qzYSHFhI5RGQfI1I1ESIo+kzlpO3koucy9/Ma4vSk7zfJAwE5YmSjhc1W9Yalo/EjQ
TBLHHq9rspkd/aYKNJXVNi9UofaUfkwGejZm0USsRRrsaKz3mOWSQdz02UQKE+FntKigAf6KSLuN
+GkxU6uFDFmv4FW8OoQR75pnBR5BMEGEgt1CUb3NY8IRnCkn3k6yL0akYEgttB611V2txEP3D5h+
XFWORs719DZyovS7cw3NXJfvEhM9hBjFqOE3I+8TPx6ahX2LEfW9HMkrU45VO3s35mMrUKBSBHJb
Ag66WiGvWsywanoReoJo0l+Hbz8akwi8xGvTrG3ykSe/npkWfJrteYL4f73W40/kQrmbpu9TpEaD
CWCflTF0bx1mG8hN5oh85G5jaygwqBg0LkleRL0txNRlxdF8VRyg+pebk0LzjWQwG7tPmPBUdOYq
x3eEc8kR4UUKYWYjNLvfZGQsPH4QcSH7zI7DLNNfrasgBHfpzmBhrfUTNqiww+Qfve64hzBki/R/
k7rT9z3kKWdq4TcbI1sUd9GOK4HMyQKqXw4zA2DMUBA3D1VE1NKyzQKjHr9yuf+lXecguSa5jDu0
kYkwNGv8jD/KQvSngNMAxyhqVImt6pUeMYTHghkDvUmaMjw3oTzyMaPcbx2EOiZNiHfye9n7kpWK
XHB/lYl9LmqDH8irI1MQcPuua0rbBzK9wSb8GoQOnF6gPIea+bypANYB9j9eVnhj8mDX5f3sZcih
fdP2CffF1Ejy9CSXhTIUfC3izGbKTr/rkIQIil85bYA7GqZlHnrgfrmY9jVP+IAHARCQEg5a4P/7
YaY60elN9qCo832KXc7gw0ITS4PppiL+t7f36BbmGDBI/Q9kNsnA8SGI7nJFat9jOrwE5x3zJw7B
A8DAG01gEkSqLB0iaEc7C5Is+dj0GD2Z7O8wSSccOKP+4LzofJg4FWAdsFpLfk3sG5ms6NkvuEk2
oHpyKLDqeLBLF6qRXXO3fTQbcYckuRfqpqcy2c8y8htVX6+/TTkBiaaHs+AxZt1pyoLe7MMO2jbj
RLv77HAUWL8DsD/Ei2BHXUnWrKOdw9mqi5QKP9TRD3bXEYm9Pam38c0qrLz8DVg/8ySVmttWaJK9
IfJhqZPaJp5XojK6pAJqFmDKxE7sQFYqT213ZI2cWBPjxE+Uu0SlZu53vOop3GCNOjATbbL93YRq
SVwhW406YGCGFhlUgMGPMW+c+52MOPaV4QtWjrcF5hZ4mRMOIm3fKRJqNklxQypYff3YnbjI3yfI
WTRCON1DWLd1vzQRSFXiaaiuPvXyRWeNXrJKzjrpQG3wzSMUQo9sSlfhSeEF0QBU392G5FEJe8SN
f+YlwgIg59uvQIlw/8bKgRl1PEBBMTRoEjmaBJ91DHivL32bCPeNfKtg+CF3ND3t6s+7bK0jwGCz
1S2zQwhekvPAg35GSO8lRwebBJm0NIy113YEOcHEmNANushk6R2aci0vOo/2P6Z3QWu/T7jwot0w
IS1LDCceDgCm7LEjfB77ECdhkfLB+1XjlB4N7CzyxYZE5AFJeOaaBmz4SAnFcKHsDmsf1LtXC4w+
r6wh3BIiPz2FsWyC5ZsUquDdvn9FmLycRs7PNTJO82xfogxn0UHj3dOeWOMQoek52BO5bPhIou1m
uJ4KaTJz8KZrtBU7fMPxi48+ewd2yjsvwFmO/prZz2qevRvagYfBJOcqstLOZ82lOe37JeBWPV1i
IRrIo7MTSVsDUtQ3TyUEbTu12m0pr0Qhkp1cWCMR6DhxGO9rl05U+xw+J1Ue0IX/vquzvCOpdpd6
dh0lFjm7RS5pDWSaK7tGjjD2zzwy0+sIdQqI9/DFdj6dT4+euac5W/tqU8b6W0HfLphecPakpYmb
E/fateCuAIKEzUt7WWHHYSfpOdECQFxxP7gERS/1gPkdtLZglQ49fgHIWUe2juYt4izANzT2lk0L
y2OAxztsbGB/hRDGVVhMTv0HmtlC3flfDfEOxSaVLIKXkIsAwdWCoHOpVfO9F6sGIwVj2v1objHv
T0cdrHpx2x49yskpiZktgICIJwErajMx2qsOPk1hWV8IgH8EduZ07HwWlNbP3fqAaB9tw7qVuIwO
e6H0Ci2JTxQAl1H2NdCY6gKZRcl/JfenDxA/yY9AgbrPm7zeM7ZfrlDsbAZ0sHgLWqU3UPJNgv4q
7MwL8tA0s55Ci1SpVmNP/v6XWuf1U8gqGipbYOoSNg1PsNti0vLzzdDBriQnGHDw9VMBsFKX9MHi
uNlsMsJ+I1DfFupqG9P437oxbIPhJ1vslxDGSrquDZriHxjYafrH5i3MqsDb8SfjPsDXLewihg5M
kgAmVVjWvlcp6ZmWVYtXaNa47KP31G6qrbtmz4z02jNOPNC90pkbprB4YUb7ocQifJ/mqH6TsKkf
WVRSzg9C0b+2uRXu8mKsEeNP9pINAi9k3+IwOEIYCKFUftz/LuSpZTL/9UxPnvcTE2C8+LU2OQOy
2/uZix7zrGQznV0dk2MxahmHFvhikKPC02tIZs44hpp8ejiVnT6XSEtyRAljwQmvC6VbE/5wljD6
X6DuJ+0Ry8SKVQawwXx5+zLajup+yR/NADWLKkP6DKcH+wVzLQB4gvdZSVxg8FkM0pvZ8ma0bV4a
g6tSPXFXOc8mF+iNrdZdWh9ftI68Ny1HHN4ZIGl/d2JjT1oIci3yziNL7Cpkw+DGRnWANLodmnis
7wFrNceUou+KEHCUQwL7z2b2tzMfkeHxktJBXaDcBRl6ANTdEJExVRQoCweF0swrrc5LJpdDxDI8
BsRBZyP/GAJUC7orv/HexgmAs035mqPj+Pr4O8okQem5bgP3zzA1cosLjfFTm32FMN794IO89nqB
o/aLotZLSjWyoLryHSdmXKdz0rYA3JKxWM02MY2eUlK5h2mzkZaNDrpmX32poyIdm/WhTr+yADa4
u72rT5QXid4EplPsAprMjc7z91nxjNHNsjc2LGucRrw2KazShJAQHuPI3qgmDo9mXxDXrggnOkjH
mSdb03NjdqlLd65cB7hk6fqKWhbGTzw1kQ6PiDFPLvEpgKpq6wAEYPzT5BYNYaKhD8dJ0t29qjnb
IUd3e0/69nVPwAG8PJWKSxUXOoTJI18BRJU2dVEosgb0XBqf3QXYMUJkIwVYG93ml5Ee1C8KX1jS
u/4Z7DpiBy38DNqyP69TEMaewSPnShC3pJ0Zl/gWv+DiY8k1OY9KoRytObgwhXYVaoosZq4XqHCy
NkgL2eNKhAqj4GZqCMNHKN3Qc1taU1v70R9o/16R4OQ9lqtijt3q+PD8/EFZNlTW6gAaP/BOIMt5
0kXINVu4KD4N22UdT2SGD6WZFjeVqH/ga35fbPH3sVRC8x4KI/fGQrAPPVurj06aAGHSYEAT6Aj7
vicTimdVn3o/1W3d4RW3kzXckKfqsDhHgPes0I7JxEU5eJ2Pk5in9lXzUPat7LNdBy9+Mz7mQqAE
pGrp4uI2S399HlsUfDqJZJan6FLZzgwZDzsvJYlFwLggWDJpnCTMOnm1aX+Jde457JS9OzsDFjWG
2Ivc8PvvB4JecHxv7zjpg7aEWG+gnVif6nDC5eUv7TOcIsoMdO7W86xD2OiCd9P5IuZn+qTLtgHc
mzP1ppRWORPXRyDuZmpIdOu2bV/NsDwzVtFtSQgLD7FYCUjvHmaew70GRd5dC+DaSmpSwmaColEn
DbkNQpby9h2sSXbQ/KwOaefkeOQ3sYeRQmhgIxT2Ebgr9dfqda/VGubhknsz/zwQxInLoRmvXiG4
p569GPZLkD4GSen1uv2RGyjfMQas2m9jiAcE1DtoOO6+LkBHEAGbQZGs819j3g8+wiRLdHaHP4TE
mvGVJpu6fFDSy65hE69HrQZTdfYT74PXbpmwonssFEXcXUuFGKruhRzICzmbsvLKdtLCS/LvxlK7
4B9lrgcZo7sulQzc07WEdBqzumxpHyF+gzBt0QvjCeei52jCYkEqyDxdPbS1R4AVg6fHEXqxV3tC
Gi5lhDwr/F3Xz760YUFPSUDn5ATNtzsmGM8fM7HuX2ESqXWw9c/KTZ/vqbmGgXLs1hdXEfEyNIOk
tUeVqYtPMStm/UfwKkTO/AYuy8QDeAFiLSg/wL2hhQ6AR4fOToLrdLVmPIqQ40ZzhsfgfBuE/OOE
ziFKlxthwoM+cHVrqVl3DmKFeA+hxM2bwsdeTzH0KvGZpAg1b+B929McrZOLkuTVWMqtCuwjEECb
S5Ckfj/bLfmpSvrnVFJIpfKWaPrALK1v14OLB+KyFmzJu6GEAhah1jRKe27H7uuWUc6dUBaA2KyG
88ndNk7lYloKQNbQfLcG1lDyvVEgAc9MKzODUklbtxHab6HsuL2yKBGF6HwkHeSG8+xEZexT2Zkl
bFtxWhlLBqbW2sI0bLUWDA6FXRm4QIEACQZHHcVjmTKG93liRDJEBzKnKkF/qsAexg5bgWa0YRrq
F1z/HZV8Q4D9TZVktZ9/2r8hcff55Jwvzt/UzMr2VvkVxcu3NXNikFpRY502imHXQTxZfLzoxTNB
uoDiXBSON8Utb2amEhbYR8SGcX2LIk4JiwiVGK5B8/cShqPphjS6F+Yx5Yvgy11XhmKTJVVPcdbJ
6Kfp1Svh/YBjQLDoTbb8e7vQQhTuyhp5Ibc0ZG0/6Ps1p4l/ReD9dTJtrfkR5B/feUOOs9WP6b28
WioFpFwZDjWvLq7ZQ/3qU9OdybBDz2dBdJtD9Iamh0pPeXJtj7GXWpD20yINd8pb5d0FqHMsRW70
Nrm0wLFySGy8v+7GoNI47ZDX7vA1LRAWEFZyJB8Nag7i0kk86+JMkc/Aum8X8wnltTRucswcoa3w
YOZdSGp2uVsmRdYXII3RFxwVbsWi0MbaSuj0GT2vt3KvIOX4W1DqcinkGbHHNsocGedlq839H0sS
QXbZqBoZxEeO6TvpiyS4FPjQO0wdnXn7y3iNnASUMu1TmZM60zduE32tnXygADs5J4mysMmaiYe2
yAHbaiCPDy67O0ieyH/X2PADfzATIH4snG+2pLFZnnjS6KKu8x/pwlLIYK06WMOG9HtLwTcn/gjZ
l9O25bs4jDeR0Kc+h0/4i0ECGYwWrfDeq0BVEfb7O6iRk8+Yb5yZ8t8dVdWPsyW/fk94eCKjxC3+
/J/lc5nsreV862zLVFVc+4FGxKRNiNgX+CJOAR7+7wTiLq1GSKUp9nBknkRpneXmRSjMWAGLxhhx
UQOuTtUX2SH6gP263HdhfiNpA61YfWxQ+qTrW8NR8fKVjcEPGDDO1GA+mcAfyPtoMOeNHJLommja
pwKXHNk0eU9qG6RXsBEDPRYgEnXFVeP2p4P9onmAx7hWOObCHurl7ypadJ8sw0+tR90pg86BW/8m
ovux5442bWNKVhJdO5pYgGnXOlykZDIgYoj2F6eXlWaFx26AQYN/aI/nHcH6gXTo0fEgucntlcU3
XM7lwy8uSUC45qa/xKgsQqAxkaHyCC+PRiW5sQ7vpfJwTD1YsQckcP3qlj0nm95ZIoxHMZMo1fS5
kczmVt9DvNlO3EubEbAUDEdV98edDcHM530KwSbH+ZRtJWM02figtKNlGFWnCuKQpgDw0lxTa2T/
y0R3l5nPzIAi4zZ6B5UhGa8Dnd8Fx+xCi9/dI0Lo3zrDezv5xVxCMz1xp20f2fbgmppp5weZ3uaE
lSfdaJsUdjr79+rjc3dPANrXcyf4Xcz7mvOqTBULr2phejyZc5sH3w0H/yN96jxQZvpkgyboQ+Wm
2lTxcwPcQADI+6vgBXAxLCczqNZPDI63Frpk+mlTO847ELPOfkEFpGtLuIhf3tvpVUqDOyEGHvgE
ZFCJu5SPPzf19CZyTiPjDoArqYSEGfFB4r2lBrhSkkxEPYl02dntpPgU9YgAFI/ftTlZcv+9QQCJ
cgiTipsv9CKjjaR6SNdCEgl5MHks469DzevnJRFqbrsve6xbsPVfQeWUB8/tzbKLp7eAIMAI7gV9
chgF5kqPVzoRHctWJHXBG82w+oPhAw5uOF4Ynfmv3Der+1ghR4kVlVukR8nztBtdmYk6gaBSTQUp
gHCCHuYS4u1BWZEaEWBPfrPDm7XXLAIUmzF6MQOqLzoPIIR0GZknzfPOoSifY7DscXhx10kHGVy7
sYnfmNlkcPhMvS5uhKvUQFnPdebqqucQXD76kFGk7ZKVbRSZhbvr121QgyiJBHOYd3v5yj0MQXwF
VkvxwMTuj+9Drfqz3FJypzrHINC00dwsJioO+7m4ysrWwL/pW2uUdFrQ0l6q06PR8yB+8oA2tqFH
90hUvm6usFxPCZHAEFOXHxLtK6Yq6ZRZH9yxzI0pFgI37Yal9zY/DJEPWLtqA7pTzzbw8+GQn8mx
kI6xSNC8X0l8K8CFjL/4Ld3emJZrzuBsRVfWS9awk43+BXEWbODuIJuYCQ6k9orRtlHDg6TkxCdk
la8YsH0ImHROZAZ5LnWetFI+kI95sb9B+tHoBs5UYYdwcqADyI7P1LnpMsCSx3ODV4xB93tQk77/
bV1g1SjE1CI26x6yV59NHFfZEsraXdekRIxtiMfOrP3cwDk8Yd3RQ7incM4aNqybfabMxUhbWtE1
oXhpyQenD+nUfBWQpdAuCKfolIFsBKyEETkIwW+MSe3st5feRT+iyi4vH9bvDHmBpOM1aIKF69d8
x9V1v+pDANaQ1vs/qH7WBmAWM6KsiDySNHe/2ntZwXWF5PorkXDghEMEtwZ6mPCEFZBiL5IcPZ2G
1VVo8WfhZUPChuO0IN+dJdw4At89dqox1ojeJ59+6fJB+zxU4nZoJWEs6H3IHaWurLwqmkazDaKc
68R2qqxYn1DQf4tR1PSoFzcr30ygP9OZvzY6TKAcVAhKNxeicmzYeirkz6TzWfsoh7DiWtd18NrX
DpaEYxgLX8mIsLO/D5Z14NQ7bRNPIiTvgOlXY+wFy7K5CvyxXlOEgjD73NBax82xRxLZRh54c1H1
TNcJdvhfbhTdkFkjMIEFAkmGcE19KXW4G0MWa6HZthNgobqjmAJIzaittL3QjOGLbFuuzXwIVbyG
jvvKk+DGHNasudp8dE+L/pT7pqcGbEPj4tDo+DPrh1aECxRL1/WdmR0q/sJTY/gklzmGzeZpJV/Z
wZX/vM+Pzau8uxE97eOTkeO1gOY+604yD2H4hQwMmfQvTLNxZzJQhmJFpi6cSHGIMZ8AYxv9VDOW
yzzoCRQ5FLmmPMQq1Za7T+e5Cx+Pati791bW65McNPGEPtyIKDokdBh7T8h3nYF1vpj+YRd5JRQV
Ps8QPgTDTxqve1bZNFbWeUspyRMeIOW2O88O5TczvWZf8cxKl9bOAg/7q3XyADbiE5iT8WBrsu8x
Sg/0xWePUF6RNL4NmyivbSyfk6FWbFeZlzYpiOtH9kWfKl0sgsI0AKjJbyxzwuXekcywvYrRKcfA
IF9ej5snOcUFmOblnrP2ZD0dcTGb+5MAyYaKgVJGdehKyKEHIqZEJ4Ag6ZL0/qH5GqgIvigbPPSq
04jdHBauOiJGJID3uKebetXgV0Qui3fWlGr3L0yo/sBEJQ8gyJoUhzJEmeVSBy4akmrsIXnyKUtn
jv60Jj6hoDAve7RVEDvd8o8vSJ8cgPtPcvuw0oEgrsLzZX2hvmUjTQYVqAjsz4Zr8hFjO3C3YpgD
BBxAESn09xd9DK7r4JxdiZ1dEVO3goKa4/KjA0yHSjcElrDzvB29DW9PBN084y0ELwYKFqJvhA3Q
VbmylZZLB7pfMEX0WW1Y+8GH5lD1EQWtWK2ZIt/6yZbP306MjaZVtjNJEuSG6AmZlRMRHyzIiUWu
b11IP+uvzfsKmTaD1z3YesfWdk2ZfU+2wSTFLwAk9Kf3wFCUHRFXaL1R75MNm4oVb6eV4z49usPN
k2rDm4UXMOVMOH4dCrQhDFmNWIlgwwKWghE2qeb9Rs0NyHVqJr+9yPL+gDwNVFgisPW8xcjwypZZ
AH+IryIOOIvR6ZdtczDnLFNt/YnhrXRcGfKeUmcAoES3/+9G9FNrLzFiSKLEbNwUHnvE4yv3IuNN
iN1mPRQhmKSobesSbUgIGYu6tDrQoFOscy0/BO8GbzV4PuWRnSyhc4MG9T84y4IPUlnV8J5oNkaB
9QI72gdj07GKM6NgrZQ3SSSzfYNOjfIppyT0S/rc0fl4+aD68mSwtXRZ0CT0jQ3ZbpCwUU1jK/3o
l91EYSPG/jXYUSKV++q+3ZVLTXW0n9RIyYnL5Rzkii3gudiyIOtJxLr+gVKcm6u4f6ltMpCzikQn
lYthpiT6J6EO5KQgJX5lfxLy+yhM4SRBGJCESYKrEfchqbY1G7vap9U2cTfb8cZHeEouJLoCEsUc
A5jIubSLO+mm8RkkzL3QyVMRvPp/NZ+WS/C+2i1exuEns5fOzV3TaWiC/AgaFmZiIUeItNszq1Eh
E/PBOR4BN64iTGESEcC6d6wEx0NoSDTfdj/BwJvWP0ottnHhh5xFy29EgBpF5sy7f6xPOAyzifWo
BLuWbiXFwuaU0UYXsce5gl2T8QKf1bwGy5XfFLUc52z4tWRdFMdcO3qJ7TmwMjOE6wscZxbJ36fT
Dt60RJbMiCyiHV0KotT0ay8ZW4dJWWIAlfazizSX31B+JUD6fqTxKuMpS+b/50TnkNYqoR0c+olq
G3E1YnMDUMnYujAYGaIyybM+EgRERelusaY/EGiA/sSA10SDXSrJ1Ko0tf347hi1A+L4nYJR35Y2
BrcgwtFMVnr488gR3k9iYnIQaH+F1+wa18DQl55GHV0a5xmjRUocVLc9MhnOY+1tbdSjD72AWH1P
8wYB26Rf0j2oeBPDfqcWJyuCWU4MKykmN4lbTeu9l1wLY4C8Cvc5U5SZ7CY8wUXzQh8KkxqgXefC
XCTOCrtgw80O9JGIx1CsUzh8TY5X/2YJc7QOVbZIbSBXmtv8pCW/4zl1fMZpVG46bnYgDPp7x1/T
Cyyi5eVALx3hCj0SLmtdBn1YByPr6pVv8iBP4VIQONtFOQ8rd5svSDSA8SRl5j12UcZaurfj2Pu0
z9JLJvvNVMV3IURh8MTTCNANrIjN+YRFukh1dZ8tfccTAaybBuDz3z3xt0ZUxseql64BdTMJPTlt
E5KmqgbY1cR4BXNeDjOJB1Jb8CJeJpmKDN0uPm2rdPVmTzVXuuozIgjrMklpiThG+S2PgLQ0m7Je
8zmesEX3jY02zaXT/cDqaq8LESwN1JnYFTuPTVtTfHpsuoQLgfaKsEp49P+YImG9xoaPnQwMww3P
FElYLGSyGmXlEpQwoA3U251PPXqvluK61mF0J6XXPUBH+0rMFK9vQvOtHQHTLzHOYHyKdXB5psX0
eB/rWVqOd4iXda/WRRiQMKVOSLBIry24ppIyYhLa+JD15FIfMm11EOFDMlTZt/zWl4rIU409wSXc
KbVDWA+5fbXTiWG2kwlQ361rfVJ6gnTLXGQbzJV8nyU/M8lFhibsgoFubYt0hN51mavhrrXUr4Zk
Nc7TyUVTyV+i0k7jWK7KWWSkF8S21i+fbQLOLyrPEhI71+IEEgM66FOX5Iu3WfX5glwZ5bdfWHKx
G9s9oLg2yM35GIah2v2JZWkeQdMr26nzvhTieYIRXGUgRxgqcyhR3opLrvcFmrNX1QtQiP9VfJWR
3TrNcnm9etayUAGLbW68nxkOirTbeb/DJZapw06+LdF4LkoLAdKiLCRjsr3Yq3CYYDnZ53unwGmT
KxC3Tx9l3jKsH96M+MxW5MBbeYwV+gorhnGBSS+2ZbfSbPA0GHJY3Q0otfg7bunNr2DkTTIhnKnJ
1FgnVRxwtDV+algBHts2KwBfekHwlS2bJRp9v2KXd7D9a1OPxI0TObSuHoGYox3px0GitHnaFKaX
YlOzmaoGVGYv/gd6VtEVK1va8omqY7Z8pDynzl1pHNWxbLdwIn12HIdPPwZZ09oK7OM8DKC41xi8
MTOy50rduAvinHDcHzQKGtvpeKR2sbWxCf6NDUNKAlRxJ+EEPEYVHsL9ZSfYlq5ygRDydVa+MQZR
pz2KLadX27T20BdJVBZJukYDzrrsufnjJ/pWLweQHw7EUuNa456m5/5FHfp6nKnU1Vni4X7+rrX/
Mo3xJQjbGwqOAsRZxxLf/gX9N5Fq4IvgXTjsLklTizC7jHJpj/7LNVy2A3ZQmlmQnlz+yz/0EgOo
09Lpi/JolhMXWBpW/bdkuMqjaAMQ7gmNuUbf6HU9uaxwJfEdWpRDD3OAYrrkkfY9UyHpM1x/s9CY
g/fA2KA4ILcqZ2s4+COG9ghOgUvGZzXP70ZFkxIM/WgtF2U17Ob7U4G77tWoRpwycv4Ntrh2La3c
JMSUY1viWBUVLySLzl2q9b4IJyKgHzC/UADTx6ELBxhWcEV9ULeDIkGDR0M5kjhv5pnA+SqozN7t
ylm9h8w2ES4HbkpnnZpXMg/tghuwodGNC1LvOv/rZbiBhWxaoD4mvjVfvVoqzroX2tYY5Iv1L3mM
mWH3qLDWMggZKrhZ3PXzysjYWHzH9xaAP9q5clqe8tfD1sR1fxAIidwpmYqDdx1vCw4NheQ9VL5u
JKmjOxWM1SR1BN2INN2Rx+lsOHWDNNGxmcg6S9u2iR+ZXNFEQAKD9ccA/vDs1oQJb/ITAqnxrguf
jdUDW7XAk06hjxs1MMkoy5iYKoRmiLwBHiQbu3kW5gefVNYQItqu0ZaJ4uNEJMlol61B3kUOtX1V
V1mvRUeB+UNfRTvNRF3hFvysiJ80aNhdpED7IgfR/QI+EWXl6xq5V6Rk874IGIMQ+WnrxopDBArV
SpYiqfRJWI03EsAa0HRKG4cKYz5VQoy8ZsUUqm8OFAZ82OafjAp2lcYn06Do/M96jSTdHTug0S+p
9vBTQv7hn/hp88SimJgUFTxuIhxQS8i0cbU4oaMAFkA3RgMZySfAFhBeRF4JuSBMCaehfl9cBNCH
0S+jH6/6DuIlK4EZwCG3kCiCn9zJ6x/v2Y/5SV9xMIrQZx+akH/MjYrEYyZmTGhRJ//2me66acw3
4KozoRE+EVH7bLHEtd0+lzygkv///r2A2ROerIf7q9yAnHIB1k1mRAulc/Aw/LteCk7bpR0bqIW3
O9RRR2lQzmWOZtDvPuy4FV4RxbmV/X1IS3f78OOCuaQ8ldbEcQ6KR42QcyODecBWYrDXX8A4vU1P
TFV66m83BJnPNlEcwxsEiNpEdajbrb3LPE9e7j8CszLHdIbwgSUpdG3XyVLGrB5oqJY6VeEGmd12
GrfB1fFGolTzDzdosnqCVI9AWaQDgN58sJEeIG+wGS0XPEqNrKNRyWTIkWH9pMceAVgnhAWDcUHS
tjNC07IKU0y7VnsIzbxiwA0Q69cp5efUAdOPNcAoVxMSqP7wvd9DEcda/hJg0sQvwDYf2bufVQfw
r9SCqkSQbzPhB7osewW5uTz5DWXNFREDXrIXsIQ2LUTu6re+U2jo7D+MJbwsI9osUX/ZEUPERIxt
4KbmiXR0SNcp/Aqgw/SlmOPHtJdMNAkwP3a2fv7sDZQGii1jBmh2RvxsedU3rGKP0g5LFENipRzl
3RK56mtIGOhCkRk3FgRQkmFd/p/JyIa2O6QDWvaY4d2LBozsGG3+e93fPH0jV7+gIuPi7rMxaTRm
FylZcmXPjg2Eqa36Ho8WS6pqnKFNSH2wqV05fKEAvmwDq4hJFRAPoJAEMqKu/dWKssATwXLy28to
AO2joQ3oh5uM7KS0jWqg/yoz1/ewyQUvoogRLbnAf5EO22M6UIFrznx0up/s7/VBzaUfsOOOeNeE
6kOScOnAodRFEGjO4maaXz1gdePIKX6g5aHtDFt90hOQ5HLsm0KF4TjzYOzv6rsmyJ3A6MK1+6Hd
6TwUIJbM50KTKlTYKYEwisuiKItrpthYLQ7x9vk65X6i27sCQBhQ//xc4D8JXBh6USx9G06pMP1y
XRJ1M6njHlf5krmZ53w8FWlmVNPjn5HmBMhfzqwH0+60FdVkaJNW8YI0Yy+BUVrdcV1vfLhZppge
YDdhWJKtMTTkLlJ+JED6MU7pNDb6ayzmUM6mCLLOlouVFhU63HXwr0MwMSDpP+JyFGHl4Se0SwLY
Fb1nB7vsbgrY8inNUSTpKLQZwWXWeRMW0g7c+vK8Lllm4WNGFqp3v4xUcHd92AXN1DP2H5dv1v5x
54TXxxyUQ2jegpQMg9NU7R+j2+5YLzLOoBi4Bb0ldHTcdslPrbGcnmmbC2VOEZPGPmQdVqlBBb0v
PD7JN3OdTY5Pn0Ly0q/MSfj9LbNJr5giteFrNmnRDiBy0wFwYhtMV8NS0JJOH6zgLfmAwwTGikot
yAszuRG+g3eL+qaMy8MX+EYpg0rNNOX6bVHJgbFhPBiis/kG/Dcoi5I/yueA36MERtz2RRU33Ik1
CBJMg85TgrKQwuPyGpPmA67qo/fkERDF/blEyw55T5KTPMO8VOC18fiFwr4/Ow/xl5ApUVWQp7ix
vlI4k2Ry6yb1Hmmz4wgHSmKdlPN+TlSCVKrRI/OVSa+2ALmcxjeQS980HLXWsQoQeEuFCJUa5tN9
iFhR+lDb2SqgwFbJhkp7Cred8nReji/vpUtfG1Hm7xtcDGrAfbvXfa6+RB+I8iIuXzGyup688R0v
n+ylazlwpWPVJ5wOmL9LYLUDhM1phh4pkQuPYseknI5A8buLlOX6CSPv/l6CAEzO2CQ2T3isykdX
titOcFWtrFvp4s+h3kS4DwbK9u61UOoxJ+zBWX9R8mzDmCWOnyAT71Qf0BslMBmhp+MFo1MV0mL+
lUMOkynrs1HUKqCDUAeX6dQCWn4+CL2l/9HFrKtz681u9yHz8Y172XpmHCZ4v7/Ms2T9r1Fsf9PO
vSHHabXFgyDj9HLfui3LLTuDAW/ufGEI48cvvwKLORtg1Jshc4Iz0QDoAsMVWrKWnX8JI4RXaw0D
xnOa6kgIk8LfyLcC8M/xdkKQUQ2cOBMSe4bN9YzQ4793YFJrYL8G/oVsDn6Nyx9EjjomGNp+3cFA
0Njzlwni6bqCVp8ZWwWiYU81+lHOnbRUnx492MPhnwxsmMe33zXDwi2X8pNU8iphQClduW9BeShX
3Azo8OxPwmP+qEIv9nZWRVGM1+b9+YwvrHvFe6QRKbjS2fn5IbUIzX1G8wR1oIFNUXLbFsrBVN2I
nbpeqSvrW+hYHaUFZdVh6FG6rO+2NIuySOELu4gk/4PXTD+SP9JyZZi7URlG0OkKtc9aMT+/SfZe
3hWhsxbXlL+EELgwUBvxJOMuE9DSAeiVwreMxEL4fZzQu7zJfTJV8u5Kt4PO/xRmLVA/wmgvoyMp
bCzPkPP6Q0mgcIARSQ1NeSEET1pUTujxeJK/E+Qlz4UtjyEbeXNYK1g+RD63dEZ4YD6v04tBRluy
8VmzIr1sfY0xeDxqHnp0u3VD/ffX3L5JFC8jOYzHzUwU1r01hCP4WhnTmUoWioFu2Z5ZbpqiXzTT
iQ2bDQJwn07kONvOimqE8TATU5oHEBVwKRXOG+1bKEt0JvTgjzqICZRDfIof/U3autBk/CRaPrYD
rEuWtuS1UeY+I2HLWGyZM4P5rmONyxhOghsogkM1RCngLnaJi5VG20rKYzRJHS44mJQ+qfnI90/y
TJnVoPQJ785kNgcsqdnbM3FzsGHoi1DkJ3WmscTqWXXEbGF67/JmOXgeJk/58mxUsb2VU0ha1qjO
sdwOMoRAvAaFwHV2VMq0Z0+GKcZZFFj+fl+aBbHwqcdfD+EMezUyBzEQgsxhIpKjZn8pwMxONPcP
4Y9sUcLYTBgV/1JXeA14RpWTgNuMAwna//c9cIbgZ7s7VtfyCl4R26uw+KYtJkExVataFgAavuxC
xGMsEFDShf9gBoDZ1mNAdfKBddbfouFU8YL6yblDVU/KBGixndNXMAyavytDgyaZvCys6VIkr0kb
N6FWEBmrDxqBiiDQHlF3FkDsajjF1HA06D2BmzPnvuIupvAzQ3rtnVW+thbriTZbNze3dbF05+2m
+H7tAEOM/LJu+vpzO1KN6VlZHlmNtOeAcq5kbrwrX8uqICoGoueZRBrJfG9YIjVWsLJuXePB4DmJ
T+GbO3o2M76jrF7PifNNT1/sMC+CmIhWc7mY+Rmr8EmUjviZ6pLwjlqUQl8WUL6KOCFfaTFg9hWq
WdICSWRoWCOGEsvUeXpUYrbWmpQzRKVQeve1UXueTrvu7zJFwxQluv84BWnX6Z52HsOL+Oo6QBPZ
as784j4Fv1rQlngaTXkhyu9Zsw9OLsaRh6Id1N+w2vXXA59raRMxvrDsIgCAbwe+psfZrK9Qx0/t
mEjr3/BLPpJRYx/MUzVIy2EkVgbp97M/+MUdu3p4z6BvsmEgs9Ivkzvzjl1cui45qpn+n6txFINv
VAGu+l72yjEOZxp5d87vJqhmGIRcHc43JsllDk+UPdZTRgbf0IOU57mf3TsUCKOe7r1R9enGZvkK
QscQlwiOJ+5zuodHCrcihz5Qcv2OtsQdw8SEHfnRdgE8ltCWg5DT/UDdAebFrlH3diYvLQkC2Upe
q7FBjaqwmU/5KVM9VWVA0GRscy32ThL+QWt6mkxPmNhsRhhCxJjbNLfWX6xG/HqpvY0v4ykzTeBa
5ps16uqQQzskqggAzBgt3tB0jCZz8516mGwqIFlobSKQexmhxaFfPyA6pPMwKxsfLS+oVq0ZP6dU
ve4uAjdH9zq9gO1ds0ziEFTjqzsvyxne2gv7KigFzcAyZQD0Xyc3N0uxHwEK6Wa7P88L89eqMmFO
Z0SkfO2NnqV3yCgeIWQIF2eFjn+7vTPM6GTA7DPVZEzTjY4rrXmqyTrwPAKn/eX8upUr0c2Ga14M
lo7cTC62Ow61IHPfXAnidsi7aAGmxsJbNvzxWQqFrGJs7e3cgosWBcJYoETwKsf4JF2h528xe2XI
zW3qRIrkDetenbje9acTY9HD5Kr/IAZwwa/5/qlIAuEv47U/9x8LU3GqtfLexxAR7N77VfO/NIyV
0/BdlUmC/JNbt4QSJEbxD+9rjfjDpPT7pagnaidduMdd4znZnnAoC3q80eFz5rZ+zaRqVrnHl2HY
9x/u0xgYt9PuVVKD9YS/IJ8YtU7gOX7ZR/FCqdfgZPWBGgkquzOgbKsbkHTxePzyRwXZ46BbVrKx
IWLKTnpWyTtNKSyR6L0Pv/i3ADCUZgf3k3dysasmwzuwHGPB0bzrlYmAS/UM+sEKpEy//0ZB38b2
S8d9NkdoDWKJgojKxiZZ3nHDacZno13drTH7nzJLiBLvmnAOH7O1rsGBrVXiGdxSk/Y08Mu0FoOu
5agAs43jA3LQ1vXMZ4/88vlDF4ZKF2hYzzNal/T/Y/CJsf0u54Q2+omfrtZpZZVH3aR8X2L/ZzMf
9B/rpsVRhext1N0IoN0kFLy2ysI+iwvSbejLZ9TwH0F7TAhV6p59PMuTrl74F6PCQ/tssJ8buZeM
gE/aqSDRitgT33LmYPSwjbuEIuqKChZJ+xldB7IQntuQYAstCwIAqqfEoiEo8Tnr8t+tSQs8eoaG
a2XOpC2oRuxMowmyCWJ7ND4xS7BRjO7eQlLh3tixwKFNNBwNHvzkwb9w+ItE4dhLXsYPK3x293FU
1GEl+aqPCg0dUupkRIPQVWPenyQhCqB5J8SPGWqnAkqhkaboiP6XFsYN4U91tAXGFLLCbXsvXNsw
eeWyaKIDcopmGxXzjcW5MkqjN01H5LPM99AU8vtaHVcRRd8+akU8QHJXzVfNLjq6b9PJoxBABEQC
QSPQiSMN8O7XS52bthu4ijRWYBMKViaDRharnYs7HVw6ggdkyy+ZrXSowvfoj+SQxY2KFDBPvv79
wtfvPXviSf70WrrFeBIjoCuPWbqdJt2THo2PmgNmVyW1b+op2A/SnaX7LJ3lL+dGruxLXuTcRuOo
XrOM6YnSkJESrtPnmBRWHpxVOzUUw3L97Rc7j4LIiR24Rg2+Nw+VLuwj8XhnIumP4EAgkmRjd835
tX+ylyWkCRl/w+s6KCnTfQEhvMD/7R8uNm/cNckbZy/NKvtWTHO6HvnDLe9A4A6i2HqsD7QLptOj
7rAxR8LvBTcvfvJMEwn7KoKGMI6Fl+1SfkkuYu4cAaRzDpf93CgxmXeCr1sSQvfjSO6rB4m5/AR+
t2Fy4pzbBx8BE02OjxDnZlwVP6mfwKlpjQafw7GH62Gbm/RAAj38WPR4LRQgjOTwRD2KndYQDf/s
OIegJgTmsWQ+u4gjdVLzbRPYSEaykcM9MaHqtV+7526LvIJd+w+jvf5zVhoykUNVVXYVKEglS3Dc
oDz9EuOxX3X6gQiRk1/DK0T535FNcL7nsBAEuvCbtS5PRXSLxpk2ecIlnmT9QBFUhKFvfjjwMIXK
lw5uu4wyc9q8qb6648YRCsZObX1E3OIpmHQDxamqiXsxYlWRyt8C1fyDDtNcrSoAnc3f2/rX2XNv
8XErkbZttdKJ8lGigohfYv1GEr7edRzO79dlW+UWnGlKks1ZfniL08IRvkxJ79xeeH7LIOccGZi0
rLoYa+QY/UT5e36bZEG5nvDHa0AsaGYvBzBfp3BYNe+MhclI38BqimxMVG9SP2mdw77JC9+tm8QE
1tO24om9hT99AhUWBl8mWiVStR52RYpxHqYzVOBoTaYTm/iLbncODI9TiZvwvgeNc5aR+vH28BrO
caKEQ/dnfpITU+hxQKCEmrfh4Jn9yl2jdYWGf9dtRWZZzIcYP7Raq1cbySpH1NUTLJY0zmeXORBc
m6H9S8+9odIhFUJbQkDa7Tkg7oTAfYbBRMLXB1THm1RL4/reMidAfV4aIuqyLVfwm9qhJqYlSp1j
c7bQp2+tbVRcnuD/0JRM1fUfsdW0HOG2vEgTUe5Soj5q54wJOggHgMLtCup4nt+zk+MyLMPLoD1o
aUYCkQOvDwk/nXJfiFeF9HwLIRj00ijaYjKV2APTsLmn8Zd4Lb9WlUoZL8e+GQI7gBciqQRMtHGd
AEyl/6GMUgtFgu3jbmW+NCNOYjAriYq0gs55eJCgTbDDxnjOvm83KCDb7V76DuOm/wqQEsnmBTnw
D26xAb+j53qiidkzpYMQ9GH1XPTCAvVRYlC41Tk7s4+/Gq6bkW/AeifkQGd96M8oTjAK2rwIrAVZ
fWvUzvr9WEfxaskJsR+FjSpPadLNXtXXPSf3iLNvlzgrqB0z7xYaaDkmSA0oOoBRUgv7LaMH8TZ9
y7ntizntidYdsrAD0Ni5ffULUA0m5YPqRlpoJXR56To2e3lk1XeNyvvDBS1XkPVeGgN1327u9IIk
uh7RCNA+j1cokrm9CqxpIT1q1L1SFRmY5SiJfH7qgVZghoBmtmgaApMmNUlNTbMrT1s9LOdL8IoF
Nz2gMLN2wF3N1sSL4B3fClnY1wovRhUaamO6Rgkl1JgPwFS5K3MLXP/0cEIy9zvDnI+rRB1HDDgu
gQJAuu37luldU5ca71ZqrBFN6gd11QhA0m4OEMVIHTIsRv5UWbwLZQ4+nh+UIUBq+G6QQWoykJRP
1ABk5uvKyTL8IaH2gDKCU3WKIwjP+gIeCXcUx5PXNaejS3kGMA+2C5TUW1raDrjWHgJU6M0bGk+Y
vjQuRrCiHf224PNOy2GJDpN40yQvX4R3HIAdkC0C2PUd1cLmB6OTBLB4iJLCfrQ9+3HAOTeN+iRP
wQUsSoRZrWFdbPgU6iPhpduPdm8wErehjj0P3Wpgw5/hI0mOnvQrsqPTSB+a0Y5WCB98AD/u4Yzp
ezgFGOG7BTxUJg1JxEkkwv3NwXc7LpULZQ/psADRjWXv3pfP1PMQ5+K+EHJltbT3y0zb4j6LV8yz
ecugmlZzTj2AfKVIfotse6oVQbpwLMtqXXqM6f0uokQGpkfvNK+1WrHbc/ooCyZN8Mxfzg2Xer3c
37a6kXS0G71nhOMKdGf/FcLdQu9wkwEwSALgKWSh/FOi2NHDKRd2jbJpMUwSa5k/J78Aa8dU4EHP
TLhCoSZTsgNbNy5dHQyz9JQRdV1mJIdr8j+IINxgpKQN1NR0xJDlQD/OOzqAbcAiqZXdGuq1ODdQ
HkXHgdITZtnFdtpFH7OgkAwwf0h/Pc4/+6SKJ9HfXq/SYQW8XWywFqyy0ep85ev7JqDJnrte/thI
3T770o3GPVDgqxF9qtHn0jVDqcbJeZVRQ8LTpTwFk3vpXHbsRmkBLeeR8aAiiMhluNb+Cmh4qs9m
LSPBPYKt6fc4VaUuufc9s33uSUS6e214+eNbYQg2YoTlBZ0tv10YDoj7hZsKihM4w9+6tHIZ9fQV
7kAOIg+stLSErHc8WBf2atShUTqKezYjP1NSsRVXcAP86b7GSfqICKfsmvDVvZALLclcm7nSRABc
HfpwmgZ0e+nuudLG3M2G6bFmlrI/BZjsVjxfX2iexRTvlgu5SWprzKcYve+jblt+8PLd/l3XHsSP
SKTJfsjFnEuNb7qMx+WLrAuN7LqyEU97fp9sfRmmeu3DAdBskpXaNtMuliB8DKJAVD1SW8ITwmIl
PdMFIsY6OfWRpK9HVuCbeHp8NUyuBtELF453doM66GlNvG5kBGqxXMwvAdvTjlFnlwaHsvjU8Mj8
juid/s0lIzC6q/HnT4rSnj3nLVK4tXBanCgb0GsrFpKzSyo6HLRD4HfIwZJJP4B6dTRgL/Ri7c4E
cWkVaozdsTk4XoESZz8P/7nnCqSQb7D49whKt1Ik/vXxGRmprXTT/hIR28P6NZLA1CApY5GG2DiV
Sc+6dVveUV1tW2mLK9JaxlyGL/r7AGtK1XtS/Ub8OtQGbBXlVnB27oaQJM6ErXIUA1lkckjq8Jhb
YL1szJtfWDFKgx3fh13sCS2SV1Jq9jb+cbSHdVr9xvTL431sJApz3AJzzHL9DFGC3U4MunFSEDbe
PHY9DfPTIVve9cImX5dVRRg3QTD2J47XUReOcCD4Dup6Hz2ORDuSn1XjxWYFtrtHifdCLfKsjGh6
wtAYUDSEuBRISn+imyWqSEMtNwTVRqXILxfHtUwTUGquGZNzC7E3/9ukcksiOZR2kXa2Rek9Cjn6
II8+cLZkHrcJHB5ihiqGm9tG4kaOBI6LxbHpnty49RcwDwB8bQRCs3m1WMuXo52wLCUi+wyPOeUX
Q6vrAMVjWK9d/fetUc/712olK19orHqX+wyfPiBsJ95k3+4Ma+PhUpq7Hsx16UYx+CNuso4PibCF
LKP8rasFr5zMK46AdcXvM7mFN24rCWtrWZF6WQ1qEEUYzqGGCnyrLFl/yONBoorxSLlTXNXA/Amq
60EtgKerv4mIONGqs+I2sqfnf/IGS+CzesnZN6CHGQcaUmMcmsSUhNBZwkFJjiCEk+Cy+JPNiBFq
q0ZkxD+/0g/6vAhjA6dA7UJXrIKUe02L7aN1SAr1MDFPcq3pXyBnyEJoqZkTG6lyRM1NHTfGqWb9
1nM0b7PbeAhRsa6dinSsJ04bTU+Hg6J2USGAHQkAaoiD3gfixOvUO3xgdDra9uwOzYdukykUH/hl
7JTb04nrMIZ/liRccCXxoUu0JcQIDJS4WwZA4SqbJmjEK20FKiWExXQ37R2MlllljtbHAa/fmkkH
3PDoZJ8HZ4fZouvURtLiLqPo1sjvXvytwHoCCwKeJu8XATfegwSrWpyiZZVJV2t7v/H837hEV6/B
kgjkcfUHLLITLme9N5sv+h2oynNI8C5UAZLWAICEBASG28LKnAE+2f4b5RnRrYVVx/AklUNITBBx
iqQj+hGs5XMZ918GJrYocCtngGDqYAps57Jpzjn+dzJvBpcxrnQ/A6Z3hI/zHztqXsokcnuh+jZ/
5RQcddKK6igO1RunUjlGBEHxjrjMblJi4mRLlKMjzo8Y9XjUJe23ioKXb5gJ7tujxH1VPj8uUclX
aoIpUO4s9ZYrnx9PBEGVY0gWnbylKndjQTRL7mQPlz43f13dd0Kap7n+gUsCPmU+4ZOiPTdFBjsA
DLSSpmGoLISJR7FvE/hF/VJLjfJI0noVfkDkols5in8Z2x3qR1/05v96ffOzKhxDm8h6no3LmE7H
7IvfQPv+Ysud4MJ1wL1/jkTy4gf7+swjC/wtREpN6sUivh1hjFMO/u2cqZYB59MQlowIp92kpvvN
8MUbeJc2sjlg3j9H/foJVX6dMYg4suniJ3yW1u+bgU+Aybf7WSkgvCUJQjF+PoWJqffvuLGWIF3q
Q6H275STFC2Nxr1zTpmermEBoQotmBkii9QnukFC7XDEjojfDhACzkjpKRkQNtOTSQMDSRxa/L0O
gyx8eM+fUVkbEGcuQG023IH//o4NvlWFmIYdoPiaEyohshPC1PsZ9rdNKBAipEDBZc8M3LLXOpBr
/OrUedyc7mjF2XCvSirDkmzN2Y47MWo9A+pvW2//LGZA8Vl8tQlV+nN/VElHsVFjXiJzYHVgxpUW
HShgLEYMHWU6uhFeCK30WgWkV7/O9gjxlop/CinvPCGOHclbxaU1/NTBuFM3aSdWKVE+/imk7aOU
CJqkc92qzKZl2W28hOJr3X+e9LKEwNBEgOCSPiPwzDAPnNW3Bh37J4GOqTqZ1/8UyQ512YTrmqiI
D62ONru8SIfQtPgdfRMGeCMwkD4SNwW04W5YWFTi1DzlgqwOecWQla4aOTEVbLdoNqU9/2QHi2yS
nd6zsLsOxy/HJYJS+SCWjKkzMbU9yVYgafaBhtnJMaH0hjYCn/wG5txK5XHM4eo27PU3Wji1fXGa
XbbV0vC4CJgQjEgPN56dT9BLn8IrO6p0cj8Wv8dgCaoRmPIUYpfDJ+kOD+b+NfZE9wE95kuP2Drh
FHdHWctO/7MjnVXpfj8u7UR7/jC+JRzD+rnTX87De6pNrKv5zH364fzpItZE1zswg1RLWTMYUZgS
s4Qa4QNNiwqr4+tNfUfIyvFP3gZnbxxUO6+aPrN4lzEG7dl/XjIgY0Z6mQu6kvzFm/hgljMCXfrx
zswp9TYM2y3cFlTZR0+ALJeRkqKWKT2eSkhlEC5AIytNsaiGwybPF1Aag92DxdpJIJtFJbbgqWpl
I+slqgAEGEirarjkauchUVPxv86jhdx2Z1Gyb8G+u5Sv+cee+ukEXauhWjnOy2buahsOUxXTnK9f
BOHmc7IAsVtI2d1MDOyygRrhM81hNnNDOG/nmxUZqmMbz6+vjsrmUOIeRjuZlNroYZcXOVsgQ7qN
VU8/O9Dzfqv9Zy9OGJwHyJ0wnegrIdVZFTk/M9rpw8ZXUgLl0n9d0Aplh5e1MYhuNZ6G1nE2b3bp
6BqoUvTKgWkiVMWqeMKyWjDk2V85oqUlDurjFJs0lZl2P0EIEAuHybRrqZvQTAbGCw5HxvoO2rec
xkUf5eCP65WLGSV3l5FslOeM7boKAkQf5k9YTA5obnTU0vXCNPkNDyZpZvUiq5yeAef4vgEW0eqe
PbFYJ6tJlRm0d38V+gFNYHGYZ9bOgrj0atXhB0rVB8SzpouN+pLU8WyGpxZMjo7oku9kN+6stxEy
FVfRalTMFK3kjaGbdq5rXtDslL5RojkLgfgHIdp0mp6xcIV3xoUvK5ywYJVniwGRMQEfYHWqjqRe
HOobTk8VYG8Oh4iFF7RQcG3tMgMvkrrPMhm/lIKGrriewFgfyR7vyIYSTAC7vUWeZqymi4niIWxe
Qz9vJhgfIgSC5k5BMypPU5A2pJ8uYbFkzzLI3Z4WNEWX4bh9Ev0E4UiX3+qX8GrQw7AEGSNbaMAq
I+1emHFmNvmcuKKrFfbnDQ2bVJfyvhpawXG/YZP8cvNZq7oaT/O6PWc3Vgx3JZXRsgIjpGOfghGB
JzZpTvUzekFKHn7FiPrSOLhH9s20/Vj9T97H7PqWAh68uad5Cq8p9WmXAW+Jp6HoWYwMBcTIwItn
iWHk5RFvJyhFm9Rwo2MS9Vwhl/eTwMOVbmCf9iM+bq5Qqk/n3kRK+LuiQTS4CDH91EC9UvLEsNz0
eJ84wniycC4sdnUVEQ4/E7QYzKK1TXComJwCdrTV1eywaJtk846ljJVmPaU0gN+KDJYPkpB9Dd8v
QQjrr+x2S8nGjZ3dvvWmDhUrd7MT7M5DcgXYDOKGvNmkn5EqEfP8bYpm69DJWZYbExFSMJk5wo8F
xLq15lytIURwiWC5XZBa6mP4hubjFCjseWgocGJSPoYn3/RltI7/zyS99LuH2a2NCBXI1gCehDop
5h0wPKnR2UXq/xAnxzDvzk/UoGoaAId4N4ofCiAquhn4/L/D5Jdfc+BCaxX1Vv0HqlppHoddc8Bi
TO+GAJ5I4Oqcet/moB5CkTETv61j8wConWzIsX2vbrLbz6WAzsPIceFjZoYMrAy4gmZC7s7TRuL5
rlfxj8RYBDXMoDYXo6ANI7H1gFGiYUk1i/4h2uvggLt49S5QqCEUOllWln8pIsl2jRn7VJFgrWkr
iE5stDrr95pHlgyrMYHjCYhM7P+ztG6Q1FYE9YQNkhy6DVaBD6FYu7C2hJZpt3Ny0sBodyQVgcbH
OfWQEsHPLcUIs/r6VypmRRhWEFXz+RAqI6HGB7lh46k749TrIgZuM3rp8dsgmZzdVTJyvkh8Prh5
uAKTtQRQxMQ6FihwCT6aNfF/BNejyqZkus9JQFTutW7mxMGNcuaU3XC3NOBs/V1QO6HPWwcR4FRH
WMmckBVSdm4HQOM9gG/MprExiqqx0cJyvWBZWIuJAi/eeRgMt9hKuIk3ibHLEVd7hn2jIWvYpLsS
5V5rd4wliT0vYWESIexnisnj3/coIiJhp3GIKpIZNAZHc80GDC/gezHbgkvaexuqdaTDkKaqAhpY
qEWa26qaR3u+vkbd1Tu8afOHSMczfMsNN5R/zFCVoUdcY1ESA5FmeyVkGkSczK3XTdvy/uUrMZh9
Ppb/BRR2tYZ2wtphCH61spbQy3EmiFyAu5wwlElYyxEYWcGYlH7I8iEm6/N9/7+Cp5jrGQ4JT6mm
XwfKBQok1SadiNwi7Z9xMtVgin8VsEIV+WPjSeEsirZW6aZdVf2aUMFH8boL1AxP5MOLgnl93hEX
HBqgCcghMYgojb/RaJRJiXUv0dBj+5NEAJwDbfHgtqc+MsBG+twiaJF1Is8/POO6Y6WpdxpdS9Bz
zsnhGPuqOxQ4SQz2Mw8SDdeP/zjLLlDrhKxEJk8NbFB8CBlrkJlN4YZP1XoAeBW24/ILBN/AQQBj
Am6+ShUupvQEtIhygXlh9UCSnxnfTNgw4DeEf40d+yF+w1VPS+rdrD2ZBoZEdofFd8QzUqRoHSvo
YMG23bFDTh0ngbOcoq/8O8iu6gRemHVDutrwZGEGy0AaRoyjVfXDICHAJX0oOW6zRyY87H1JGHv3
/S3BtSZEfa0Q3gCXW7tNgBKuEj+R9zUvORWiVSM489VcIkj8f41IsI5vFVuHewXpgF98LfOVCPQc
7jqtTnmOGutfLSCwjuDAzBmmeXZnEd1XnpB1cffUusDyUFe9NHyhsZ3ugpQsqPgOdQ2pQ7PndWBQ
3kGr3xzMivstcAP/fwREB9o1/0kSQ3lYIvkeW+7wtic+hc0xA9oIjG6HH46J1BoG8VTH7834Kwu2
NRvWT+vBfgToKJv01HQsvCfMq2E6e6bvw6czAqho3D6oF+/eR6P9APYnP2890BOb2LTn/O2AL6Cp
VndqJ9ZT9SrysdFSo/InlTnPZ5WcEYtyuj4nSzbvtKuOAf25CX3sOEXyTuEbiL17zCoYLiNpIcoq
lhm1WdDA7aExoksg5b4Gd5JFp/ShRjUheWGAl20h9Dj04imvV3U7dsY/GuePMbiN7WPr5dtbpxOC
ihAzshf17IttX0ZEwuIkqwEQmJSVcKVmg75hI9jxumM8ooM6I5rD6YVuoMz+9VwktftReuYVKQBo
U0/flWYJ033oikqSI372RkEq6+eP2sJ0A6vHNWeM2q2hWfniiO0p3AA8Ueo4fOw4Nz1QqBdj2pQo
jlS/3nMdMrHMmA4l1YEL18opXfS5BYywuLZ5fmdKU5EUcj5pVL4PjjNz/+4otdsH9zn3i/NTRFHG
tkw+TqiPWJQn3KhbSUPHosLfo3rmhMCXOGXPGHQy2lSuNfTkHCkReK2jdN2f8fW407RJzhwbMzEo
W5zHUYrHVLk3RT6WBI5HOeyht9rGJlKwAK3y2R9lM6nDpki5HHIYAKxru71vBwu7s791xrkY41CN
ULgEEDANJuUhfEQNbKgs+cHy01yruvZFFR/pVlNM7thxwK19K/ck69RY9kE0ohTQTlWrAB+mUdsQ
+kT/vKQnBe9/IwtH6P2Rk60kHZpAphvTOA2XkY9aX2aSXN/exp0SBgpNEUfludnSlaiB3LHNF7Na
lNnb8tCGd2mChJPf4E47L1fiXPdCJxNCZ0FgY0tw0P/bQ7qeqskvOiLnHmTYRU+MQNUM3T06vgGj
QEOkTICEW2tjFshcSUa/SYH6/yCvhPrHCUuWCKpZwW6TTrtNLlCpld0zTrby7C8JkL9Fo9a2Lb5v
ae7Ah0q+4HKyBBXQHtu+G+nLQT5/4CeUZQvqWir0dl/JP82xwhRnwGcfm/O/lFAKXxF2tXN8/hNL
7/nwFyZyQl7OV6BGanQQlWVTQIT2pXXt6uPfVWQhLDpibwQf0MhBQ2dTZF+G0pVYvQ82FqDxLRqX
CvrRkFcGNVS7lY7fdsCQsLzWCeGJWD3sBBwYyk2epdAqAntb1RFHAN/AzL9vPFG1kguwPUu/Pgv+
h5HSLOOUzIOEfuZL9Jhd3ynIXhMfrMPNYac6Gcm6DKq8jhdnPjb0tnKoXxQeie98EjAjNWTz9quV
2P1Z9Gs8R3rMEUsur8gLhiTUOpiyTAYSrPQYmCKVb8ZHStGNOsg/ayiYVIzTKtN+uBr3JHFeyPW0
a2DT9proxluspAzruJaj8irIjji0Wsmu3lztJ0gJQFdlhcCfgFnjTTzqZ/981mMAR/w3YiTwgmq9
a9vwGhVTmr1kgbxRSMLcKEA+HxaIobwuaAqC95mRku11CfOH0+YGbht4zr9yGM9dHHrvOrRQBZ02
77owYSfBt2Ns0dH6Cm9clscYQSqpkbWncOv8vv9hDwgx1fVeO7VlJigHbmXRX3V/DdMyiGYRqGHB
iMXjeCYAja3OpOv79kpU+ypocIp+QNI0W+W09sJJNVisv3yr0I4dDZX6ILDweBKjnSFM/oYoyKyJ
b7WxRpTeTclvvPqAYz/BSToVTDuOKdynJu63OQL5Ldmt20YE+CpsQFk2Q8AkEuFsqYnqnifAzoD7
eFY1SZ87+4sph8DTY7hGEfSRGdVtovmkgYUWPLHe8Vyw4drOR2GDYZjN/1om3VINGrIfm1RtmR13
BojXFuiOzL4b8DvyA/Q3wXqDUXtH4ZAfDYODQaS3cw+NkNn/juFBVWGwFrH7arnlUGEjdEfDPT1D
zt7SgmfXWKUSc+9InU/Zpf5Myref6oP931BrqYhrlCwX7kx2LQwLJMOtjtr9Ol9kSrl8/NU4fqzR
TYDJjRu+Nh/ZcLlg7G+njAvImEehdsMWdU7obx8v31nuoGE0RNj2FQ6bpQos9y6qXS83RkWrCbRS
oDEm23vYX6XfEZ3OfZUeH0FM1KUGndWS3IQysg4KbFSvyJHdiYOamwj4/8y7qdcM6o5f3Hi4Fx/k
wngMwIdpY943sIT/A/n47Q8q/KthJRCgYQkNc/QXlLIeVlONlsjZSBrZ3/+R5I4UR+AfqSazD8EL
1ha6ymXNEec8vtQFfMzaXcnIiqsW6FULPMiFVGJFGlET+kbYqM7ur0M75D/q/aHiKnFj0QbjQp4L
Y5QioRVjzbxXmvJtrMGmiU6Oj1PGFTSaLgCnQx2VhVufcxQH0Ecg37byqT2H/OSe1/Hh5UN3eJlF
Gsdxsymoey+b83nAov4MXuwd3vznJXJaDZ6K0ZX/VX5BEqYFciMoQ1noXVIxaXqK49w1Xn+/vXI8
53FmuQRECjAKsjyaoJ+ffxnDC+j0nGc8ix582iNWV+vsK8hrTfX8ZltpFTGyTHM0hVRdVwe5qXFE
Cr9ajK9nBtWM2TgFeKwqEaTdA5u1DfSE15DZeG+riN41sWFe/jinLT+bQFuxxiHCXOEY2CcNDwWQ
4CahJoNGTYyjHhXRiIDLymaUNp1L8TeH6+rGCFm2dn64u8vVT7+WiUkilw9p40grb+7PwwOkKI/H
YJGcTIt7jks9NUWHVKDxcu8qxNjLCvp8oevRbDYDPfH62CguqI6ofnlARaeGO+w1tJz6Ae31b/TU
0DMijV1ejOrqcdUB5oINdcuZ9FCDo+G4FTMDBsThTCapq66//xrRoyPcCctVGZ1jR7e956zgF1UJ
nZbmuT2gXzZv2+D0D8bAu+Njh7mRmyrUiaxyHzmaUjDHIMKQTq3W4fCtJU9B6HKcb6vqoOOFpUeY
hQ5j+l/88+1bQHW6dltU9QffRip04E16qAq+3d637m0ElfdzBlaGP8aKwII7JoiSCn60/vWqHBmb
iEXajdpi1V7hddiHuidUgERDwitAqUXW4POMeZzok7GE9vxQwDtXtJU/M8M+/fWWdtdOp0Nh2jyT
x16yLme9UfFzofoLkXCMVEKUmpCep3vp5t32RX76H2tmQIcbVb8wsrXBkN6GdQ2lWizkmDk9LuZe
D83xNd3JTcgG567J7nFCzsfWdtr7NVGKA9jpYHm4d549Rf5UK4W0a1S/4vGM7FZDuDT7BnjivNCw
BUgVB3xwjGkyhAyhs3KnoD4wN/XJsa4iEzt/UOhwjC5L/37zkZGp7QMMMNlZeZtAB0TXDw+1rlFx
PMPmRiffhmIWBTMsFnMXVgNBi13LfBaO0inbb/lSdxOiNlciaQxWUMXeJbMnJURdPrRRQsTOOHc8
9V+//rjBe7UYDMEt8uOG7qZs37JZmLD5TvASF364G5iMoCJtGiwRiTiWZCfBtZbg8bMeuGjjq+Cm
5FYqiD18A5tqELnsICzSfY1F76N0Ra9J4z5wd2sA3mPSsbKtFedE871qYK4yeF7uuXNhxAfnA0qY
k8lcOvt5wbbhbu8TN9ago/KhpYkwsOTkI+Dv32U7VONkzzUGWL8jVk0A4ClhhcFHxrUn87RADcWs
pUpYIktXwN1C58E1gb9///zgQf/+0HYWGKZCMAMy9WCi3d4xJGcZCc8ZN/sTSA9QLtUpdiTsOmlR
404Ru0gzHbV2uj4IX+7wMHCXH+cexMYLK9zOgLTnSdtwOBvnv88wQ4ZrAJlmQ7n5I1Tyr8E7xgu2
ZTy/goy0lNjBssK4ClrVsQVCmlvpPI+e3BJbOroqrzXmyV0P8SQZgEQtPAGME6UrkqdXsC7bp20F
Xtebp9EliGvikY2mJ+6zlPeRt8TdLGNLfC1iMgVfAe0Wyqb53PAVjnwz1JB0cDcZgG2Hvc/xzMp0
GydwwaC2ODQqO10K99/NrrZJzdKjMORTAEJiwMoqHAozzWw0sc5pIbp1Usxyxyb2yH7hxykQmN0F
04I3OAV9HAGPqoaMt5dMPGlD9AVd0Sq97EgMqa0UceTej9Ei3eE4+Te0yakLM5oSgPyqI66TuizE
6oB/NX6CxV0EHZglVl+WUZzmaURRxEp/zxyJ2wjJIENAu7HAKSuV0ksGXEIiUR69mjDcf4fd8NcI
S2u7GLXF5XVFh6M7OfNfMD1k4/nAQJO9biH4pEy1FiMS9Lqk7mkvfUwC5O19k5JsF/lmmQHG1mes
kjHJBCpuSuDm8wCkQD+kqqCXqnU2eRXleoyWL97nzgkB6lfYONmwttRdnch2bt0iSbBJHqNXylZx
JobEXht67YxXmCaNgw58HNTJnyWrXjU932k25coJmCl9RZ+FyoY5FagSsmLahglpUViGtgPZUeIy
TzdmaBsQbo/lHriJ3CzeNPEr3A/xaVFp6nnVDc+w4jpH5Ybz4ER2D0RdrZYtTDNoQj8DNE5YjiLY
oVhPserLzkyxauh6IBIrMLjqcPSmnIxusHNI/O7mtHV/uiqGYVldTiC+JgyKc3CyJkSYrVA0iBw2
GyEG4JS2Xg7PyQkZrM7VkGLPjQE6rA2FTvX+SGwuU0kMo3JjRoo7raVPsj+ZZr9q2xJv2M/ZMlhM
eIF2hRn8ngHU8pdLR5ZYZTzyRHFGpCSayTGEmy6yawCSDQ2IMnAyVawIQO84fx2vJKAIqIvG+Bvk
dvg2UDMs3LsXqcmeAjedwXd5ZtVlnnmQMjolYDMrzimqN/2X4pjd/td/gK2pk8Z15xm/Z0SLBMh0
Lpt3C96vPt2UaLNsbNNzXx04kfyLU93lKd9+Y9LXLSG16RLIJUOqfT9hsgJRG43ChJqdA70jNCOh
9DdykBcUUDhoaYivTSxvtxrC6jQEsxAAXev6z8er/sO+c3SiZ9+pgh9yrP0fDL4EhznivRxKLspd
s8+Q2TopxS14TcvFJQSvgYkSSVE+bmKbKxih8Es+7lKPClvmiE3vOS5MeYCJJ/ycOqLMYbv1ovb+
cpp34kHEBAFCtT7L9G9DsRIa9sL40BquMkOunsfe/oIdsHBl8ptLysSqpVUISj1psTRSgRcvuFNL
zpuQ1zz63a1wPGVvIdZ+2DGZptaGCs9NQDcUQFoB5+DcBInijVk4qcF5pNrIN0rQimnw1sPpP9Wc
QVNjTYvQDsYUuiNFdeDB/V3xmIEtUClnVQW98uFj9SrrbCgXfqSyUYS4kLfr0bqN2O4CJzAj2KG1
aABWa/gouHkibCbJdkGj/nTnLQX2GHfFWr8VIHAdw2zGZLtpgrqe+X6dGS14MhKCAIbJ+g+GJMjb
l5mdfgyAAbVOvVP/wtl4fDCfKl3pb7LWsRuYhIYqFv48NB5lGwmMtm7V8a/Yine/EgVw4UDmZNPn
kaBJT8MGkVpu8I46JcbXak1wVzw2PmYGw29UuIQoNOTzUz+tYVH86VREJy/6ekphey5zKfXieIjz
KBU3fBt3941W07uQOujEgo0Afv7/qs/JfI0ZrmrIbHGa/ZEFBze6QMnJfz3pUbTpPRY69i4x5Nj+
cGHq3KQzsz7ADf9J0eQoNC5oXowv+4IyDaMMhE0tBPCK6n9GDnIoiGBGjlOGfhVKGd2pvfp1v1WP
WBe16aQIwBR36pW1taOpkUtHkfgz1JczYSqOR95r16gxnh6RPNhCbEoQzNPLuUPHv0LV+9f055VE
l8HN8kM1q/ZYubnqYFl6nJdzQP7IG3Y4Go71kt6ielsVEZY8y2FBgKs53+LYUA5K61+vKpmx1Rvj
kvI963+tg6d7mDDXY7yM6UMhtvirCUbMeC/i5+bgPke4G/8QicN463eDCgAgh5XRB3uTYLHOBYei
i3Q+D4B41X4kfiQeR94NhBEws44tIiV7zFGB+gBtTJJkYM7w0xajxgc9Mi0fi6yUSCS54HTgNmmi
1SaEdZn/MT+UtZhrdEL4S5zxNeBKUWeuYaFcG3Zk34yoUqOigckWJYcbQv1aYrV8MMKNDHZZo9+n
gz/t1vQTrhm+CD1++rBZ3EefvFvMmaFe1kHqq9QKakmvoiM4AeBTyFdnX86OuvdA8+bakITBgNEA
Hwp+0xtSK4etK/fGSDHQPyqyRoNd4BmdDF0v/6lVH7sn6dN/skjMwu4wA+h99/oxcSrnHBCyYu9m
IoaLqyrC8QdwPTZauox1AbvD2WAv6OhTcEZUGJ1csC8S2LOZvmZSxs/wYFuRtdQSm2xEg+3FiqOq
+rbPNkmU0W1cbKm0vVAJZsS2uT/TGL4eF7pe5rv3zB6UoyY+JtOp/r3CW/d/Wlw9Jg2X2rkZPYQd
xNhjeMhU1PvpPS+hXb4qfBGkiXW6d4j4QZ4mcT1vw9S8fk1nq6smbkoT+jxL2mpj2zm0apCmcLVT
2gU79+h3dGm8oAJyFLWINOUWZFFu40G8GEwIb2jHUpkkf9uKtOpal9R9jyojstPRqOpp+336tPPE
+ec8Gmd1UYCJK9lvMGJghyEe9vJeDpKpWP70lp+JIPNBmxKV6BFRVkoqj/Iq3rhNuMjz+UYZre1m
bHgdfo9hxjksIGlZDw8Gl2/mbY3mEquZjiEqlYWfEHj6KN4mvjm7COXSDuYCS9eRBwhmrFPliSZ6
SU/QNT8JPZ1a00NcBu4L0fowz6+jCDIezR67uFMpkbUiGbdZRX3X7gvvf3jE2Ct1A2A5GkrrA+AK
ppvsUuatr6clkeeAMUjg2FgkH4rIeC1kHxHTypZjQ3gSPDStkPSQKIkrORsTuRggLfKAimLdVHOM
n/MSoIGeQuJ/zc5GmchWvRFyVbvxpup3kIPFGAvTueKOxTPFEX/D/RstjE6iATl4ECGzSj/rNyP1
zOhs3SlHtHbwuVYbCbU8JWVcINrSt0WWKg+qCuT7bxSaRzRjfsUjn0y4DMZiw6e3SJjWqtt+bcG7
3o/tFaAUs6FKbij9JbRiXLod+NtsmuGjer35DlL/zYVd7CWYtwpG9tFRW8Oh6rTzZeDxEIjWprFL
3WrJWwOf5umZogWK+fRmcdghyyKpzlIV6utpePLY0Lk4Z8lBL93rWpcp87/Ibnw49NET0qLtsGYi
idlOx39KMH4T5Q6OXwy4Zb8m7RSJyf8CV3smHmgNWb4+LLcVJt5IGcSXKpBvxlcLPmCi7BW8JuLJ
NC5gcCdij4+FhX+yQrEYQpkiBlc1UUhUMszgeMQv40gYcQ9LF8EUf65xiiniRtN5+5CN059sGg6i
f6s8wt1s801RtKV50WDZx0YL3zv4PXQnl0eEEA0VUVfc76CMF13TpD/c9D3N+oKPr7WfW+qWa2N6
/dYJ3r+GNzI96vl9TbQWMK7Fij784UGLxBH7NkjWrEODUwtZVI05b8WON4jymXywZePLHRoFsb5v
m+LLLOJ6sWLfyjEHCi5z7QFcVWczhNvhvpM58Fbn7kaKpuA+41VO1lGMWa3k+e0wXO5049pAtvOc
7nwCSj2DS8CnzESsDVDRNMYHPz8g7ZZnpf8KXZVDUB2dr+wrNh7i6n7GXoNe5N+ajbbZeDf6NvZn
deL1tCqferO0ZFV5fNhh2s+IRKPmJna6Sfv0o53LJEqhtQa5xLp9E0RW5Zhfj/fBiJe4nJtwoiUN
5IP/oMkJubwJw7BqWbDvbWvaosTLuUEA2roEqmQhWL00gexokmwCZVPnCAxNMzd70nEyOl66yhQa
1Sm2KCpXiRUFXCm41WLDIY9ES/rzCs5SBpv/HRlCAh0+DjM4epcnR1j3jpIbb+PBAfx63cAM+9nn
yZjzalypsTs15oQ7YdBN3b29F4Wj03nqj7c+8yLV3dB4nerraFbjYgKjQtS7seRyfjDxMdYTGAuF
+E8qWe8+/DM3izdlfy2yfzRxfm6S+EnJ9L4tcrtq2D9n3Y6NoxF4BQK8V7TEQaB5YXzXzcUPq7Iy
m/Q3d1840k/AGYv3TMJ2irbCDCeG9HXRmC7s4Gk4IUxDrxauZm6AmtgNEHEJHJv/QT1kzBBHHXyt
ZbeOOpX7cszQEkUV1OTo3bA/b/3XTW4y2pTatDxDw9/CaWxS3AvaXj75GhFoCLFc0WzEUvYaqAjK
YbLBgc3AdC6cwcqE5eAZzeqFT+ukKz6EkauU92v3YkmdapqBRL13pAV92tsxlQHgVjYFLgZ6ndvf
UF2UMqoOhcKK2u/DCom6IboPg5b2VLVs6EthvdXEpklsIGicnGQL1y2/WU+oNdJ2ftUBxucfkMNR
eq6XCEfZDbh3gg14steXeQi8GKEcc5SgK8UaPfOAeiY/e2OC4f0WoC7u9p1AdEl4VCX1G3QYRdxm
0uhCMXvM8hmbFRf5TEw7+sB330YTouPUdEftW2DReW+J8HWEkni/Kh/PA/vD5n/8Js5ZI8zLjk4/
AUuLKjPZkXa88Da5L9HleSa807Nqwm8B3ctv/T//QQmHIJkM/66KlqICtLrnkseAZR/gu7ET/xFP
a6Hywgcuv3nnpfvuXB6FYWj3Qoahle9mvg9qlOOAAtVzPoT+TdYmunRDbrAd3Ohe8Fp989WZT1d8
pLV63XlDr9M2RRMXIONE/xLo2L4EIznCL8zrsBs9Qh9V0GzW1Du33bc7Hwrm3EJPQZ82KhvhJpqw
wHfN26qtf1DHiZmN2bJKqYe0YXqS3VFWIML9G8r9nh1u2rFalBHnLIx6xDcXFdR8R2D173pEr0lN
ziswh+gJHyKwxJSsNeCS3UxkWBkSAXSeF1s2l16GVvlZri0uK5lWBvFTyCX0mUnb8ojoYKfsoYAT
WHYePpuheBtya0KyGPpxFH/RDE/yw/eJx3Q/eHoIdU9tuGZE+mXXmzZzPXUcfirpk5Dj826/c+yP
ZKoD6TcHfftGtkPx7nEmmh9ZOVVHpzUru7o6Qwc3nh91w4hgUhQ64zUbGLx0KvPw+0971FftVnNG
DaXE7uMcH4d/R8n1Q5q9dtUzf+vxkZdcCtsRZjXx8pjh/HrAmT8/65a4jtI96yv/jPJH5klTaelz
fUjrHSnSyvFNB9PJVfA4RkqO6/2yXct9/QPParOtVxsbiQLraRKOVEU0OVqD2M+ckngZQ2WsEQxn
fN7nWs04r8OfnyI0aNlOsLzm8/0/calpU5zUVC/8rG2BeaCnAgjzC7KnqwFNxfUmJCbx/nVKDRxE
/8IkQVmBGcqlvXVjfL4js2S9yE2fXcp6+U7LkealyNVSwQyjinXQmXWjgTMMRWlMO+oEWhys3Xs6
xC1iWDCWNW6bf3dWoyGsCSIZXyvG1b/InyxAxfy7ZJu4q/ODQhSCf7tNba2EbmDNhcLSwEuA7/IP
Q7YNXfvF/6xbWZFzD6f+M8eKU7X8HL3frRxaodWbZWeq0AUs+hypGD7drfDTCVSNt77wEt4UJkE8
kqMipvZ2UqruP7YfnlyWPMGHBdoRn0EJ7H2jaI9C4By1QGtoZFHL/UvusspKodRVVz9wv0xdOhsH
wIou5MM0cwZOTci6mVw1PoXC5y1/tNUSgJCVsHRkj0w3DYmHIJK5FdNTq2ZmUjo97Mvjds8uP70/
nQs9uOtyJy4DgNZeD+MbjmzpwC+aIfBjTSvLAWQZ90Wuj18HDvyVN1Ff3KEa8HeU6+7WrZhrF+T7
bEl2YB3b/hocfu1w4+sQKNi7sIqRiGn5NR5xyu5chw6/0qZ3+9pyA3P9Aj8GSvUKVsxQa0tbU+dz
qaRBIowt78LNDTqWor4cJ9YECQe2QYYwOQT4LhwOLLIpb2xAI7KGvCyGdTpdAJGPQsGvVmVeLisy
yCCDNWPl/oK5mJ9rPVWoBQ4f3AdLADUXEWFUDbXGSpBZwURLd5B+sDOgtkQ0DqYF6ljgVJNfswzw
c1lZjmVo3CtDYJpQoSkVy5ts1EcOXphr3CNQEIoFOlz6imDFLOKrySM0UmYWAfN6M36gZ0Fs7sRC
WFNrA1dwMuhK+WopuzjRPCpn1T62tySRRc+2KWGaFFcA5M80trWS7eAF33ndsR6UJdh7EJNUQP9i
P2/9Lyfj8HF7HCcL+WNF7OaGG1qWclETvRog+eMS7eeyac4oLXqjwHrTSEoVi0D9D/Eq3b+8YPyU
K3sGwDp+HwDsFKKbXRIBr77WUVwloSwHfe2hhlo8xB76hAvHWL4kclFyY4rJnCfP0WRjAxLHEoJu
Gm7orCJccmEHrLQ+DABsHwpoe8jN7bMhNCsC3gicKQnSIOgutYXy6ffpCW837zicFoOkzMm30rCZ
O01NFNIe8ziYmMSDlbitDK7bjIFWCmTx1YiwJwCaS57V95uP6lxB4E7l7b1ErG0FRoP8YUCcPBOu
/7HouwdnSwqwRsiW1js+U3FfLbkCKbkXsb8qqDRglGR1PVe/6RBbP24jOQoc9vLcTNpx+6CvePHW
ZEkYzI2bbxxwuSpMuLjQCGRC8xAngyjvxajDZnUEnFqMPIvIbsDNZ+gTf6zBKg15wH8i2fv67ZLS
6bGD83XOfh59XGbVh0gxlNsNwU+PfkrYcpYLcEnf53ZI1NtX2E0ECW8FnSxnOADefPLM0DAUa7HG
sOwWwov2+4twwJWH6bhH5o9Wi0kl5dCTKu/pzMOPJgPsJYxsKEcEw3O+6VhEV94deYRMzTN7EvCN
xNi7KXOxaMnSmCftBeWVZ+dK9ZKgvt7ukaDZUMyYPoC2jJJmCuqIDQVQ43/Or97hu/DLvThWWefr
Dilox0Zr4thvyluR8NHm3zCAWqkmeVSrcvoaIK74jboBD/WIK3tj6Eh9oziU3UN5EsiJ0lzYY/N+
DSjqjimt7Fl2qzm7/oUqYaZbKGYdXzo3rTECuWCxfKS4j3oH98foeToDnqXnZuc+CCqdmmK4pV+L
sVXgtGUkvHszdRa7Wz64aF9/UW/yfW5+2fZIoDonb9ggeknN9CW/CIuHJaQ+Pnne0ePs7D2iTd1W
VEmoJJD52qcDMMgV/b3MtT7K020t0/JUzWwUZIWbTCi0NfIm5+6l1KWuqOmZGGigAa9ZCz7bWkxf
FumZUAUT1+oWVQzlSlOgltJkA6x1LzFExg6pBI96LKYvq3TTJbl+IC6RqemFaDtdioRJZcBKo3ln
pK7DQplQAY+uIOYI9P83vjTu0oR3JGDhNGkSN3iCHsHoTHAbK7phh0/pGikgGBLRg0oi74qROJzG
zjurmL4lzK14ywU5xgQ4hQPtPgEH5sS5FqenTxkdRcWjT/03mbFlE3ax7ZeN4ky85UOCHCUYJeoQ
Hxql2Cmd9XSIPGMd0oAcDMfbMF2KRq+3IsfTTfoeVu89QikIj7X26Xj1RxZLdk4BSg0Z1qLjlkeK
cnBKExwKqxu8zq5BWdPTqltnzaoANyytkDcNUb4mhXhXnCTjemqLXhLfLOnxKp7gjlZysNhRWciP
0mUWyIcutwvXzcYBlPPa+Sj+TtsoRfa90uSwOVVJVvAKmUzyEx4l883Vbhkm8SKF53QGEneqolOX
cHuWTsS3bBaBMz7IUH9EMDJ1sX2TJL7FnOM4VRVbtbzimTL6MHvO0bc/dQWEiW0e8sPHQojv9uli
4IAtBz4z8r+aHsCfkWE6bg35PBVKq7zMK80MTdM97Zz+OKR9kLO8bfXpanYlvX3JcCm0A8sR86mO
ILgVs2ZQ1Pb5IXERGwiPyh/9mU//XT+xtLlEP8sgHlPBfZh6W8yWv2wFNLimcs5YVZ8zW+uOT2Q8
t8tUAtLjeruDdD5BXJC7Ws7MWP4hX9u+l7Fy6R9lFNr8EURW1xqcq0DB8wapnRV23v7KwFpfDDNQ
YrIvD7MGDB2qMUJ5jspIkz7ubR173vmjulLRFh+H16EfGIO3KO2wPezcMm33LjhFWzeZk8dZvHZv
RTnvCj0RbmJ0mbWb7quroIaAHtQ+28VyxLsAITwiVQySYkhadKAy/c/pkak4T9+yqc02gZwyY67l
yXISr8P1QpbP1yonf1ORoAtLX+7dCG0XtS0hbqPiSs3bD35HM9GnEF4mpl1ySYQA+4OFzcnF28Ug
L3yOvGfYH0erWiDz3wbCcE2vqnR1BqzXv922SuKKNtejnGRNHVMjF1vWocVYxcC2gSadlCcTueRb
O580ixewIEwUeRjb4KiXBujds1SPVVSlwj5Lp1D9QG/hpnpajsYvGg2L90ppszarML4Tf4ltB/n3
w6LodDpmo8p2YF84nx61HQHFNPTk0Ivmz8gzfo9zulDSzx/w2lz5NFChkes1VOPBuBh1+EGxvRJa
6W2r99eafeBIvWSzjFOwHXTjuYcbXUz04i8S9BExx011RmgHLYpn7P++C9kCItjhucFdZENv9z5C
3QZkGtIyZJ5WwsnejG2GSQO7G99sNtvp8eMqOXaRLnPSufKgPaf4fxmTTq4Cgt0c60fjvLGveXbg
kPN44Juq82liyJo/1TaU4ODL2z5uEBaH8l+//7Xk68l1INoM4yaOsOUptMFKdGucHiQxxPvubx9z
9FEb97DMoU1TlIG3WPm4RfjgmlOdLYLWLxQEAxIcKa7i8k/IC0OXfEpIC4Qe9i7RJvRtMgOzEsPj
YLsPjwy49mze5n8rUza+btANloh1sCXVjyRi0P70h4Zrk54+JK+3rVYFmtxP8DxKVqK39YQ7e3p5
Qynvt4MGlyzNU6POG1xERdfd7DiC+pdXl4i8HJNqLNhAKvjbIqR6oPXCJ5dhiYhbAWNIz134yVR3
LwTxPXITu3SsGwRcqsNQUihs0BmN/iV1Z17knDo62f/eyWcC2gusDEpylLeMyMqu/eUxhd04T9Fe
2ZPZfraGVOvyppivg4V1nRG46uyMDoc09tmZbBJ0JjYUKkY3+QnE0lf4bjks21Ig6e9yqQKkcn5t
9Mg5ep0/X1czLqjnam/o3Od+uIXWD2OcpMyxHklksYoEw8SzBEiyj4vhP05QeqCadq0iLuIWemFk
sHJPVMEV3/YZfdOnMvStip0QRLJmchPmqWAduJPgYAfxMHGV/5sXs/Mr3osr2GeAaycxVY4zvQ8K
6DzpDxV9M4SItSBWga0KbC/CEvsFqXCexDXEYuph7BZLxKVEVpb/7O5OksnSQgQ4WHOq+0Fm54L/
2/BgB5WwqjFA813crdLizdn2yFBoQ2bR7adB2NRcexYFv64cHcv4RMDTpe3vxKOdMX+3xh4Jtgkx
ywx355RzUTsFN63k0ODtMsIHFVYX2jQ1WEo+yD6o6+0vZ59x4xVe1nF1VwWYDUr0tT+G5d7KC/QW
yO+heJNbPLj61807bHzYHlp1jxp3+vAXRbJx/DjhaLjz0zzgRJHyXY97ZEfkJlh4OA504rWCRHT9
j7MhWUsm5ewEcfbW18JGHzqlNO9vX1iJAI5PBq0+C027fxFQrnhgVRdk3o2UrjfeD8F9hR0na6/R
mSiSeMiJJNgAM/EnhZYkhrBe2jQ5jZoizphL7weveBoj87bL3KcXwX/t/hsB3jH5JnAa52QiSfA9
3Uv5IkT6GYgEVnFrzSqGEFXa1LyBexIAbswZKHp4dRbBzGda6j2cD9Yt7ixA8hUSeaMjXbvUjlS0
S6Aq2621M2A7gj2++XPqU5DyRcPlVLGQe2e6+2hOLjspbujQKFHB+3H6MwZHKE/dpkwxX40E98qO
AfdLeZ2kdCPc0hc9P+gScy8CFbTGRqL0YmlD5GKiku8Hu9nI1K8B+zmQ7U1BcSmU5SVZFoyerPMb
uvnpk8sv0G8vxhZRqCG0zQYYRW1IFIYFWhCNGemeL5HASN+dhazxcFpeCO4j2T30ZHiyxQpQWvE2
WgGl/AT++FRDbd55L2pRs6W39i2oxYPFmz+4fuutwYAajhEH8JnWA0bCcwzZZzMzFPhXQOCXtBqa
8EQgGg1l3xp6011H/aTYqQDSy+pxe0FW71Bwv0TG6XVJwBYe7llKqnjTBC3S1I/Tq5vqxWB0XzzW
7cIFE8zvBvL0DqDyTjDyt4WtvRaHdK16OsCuCsN/C53ibjtkRvFTdZeJ3zGjZ5afU37bJw/s6EOt
GKpdK6rS0Tn5edNNIZ7+16ToKWQLmRd2JcIToNpo1aVBEsrJyAI5ajKso11SEdBer/n2wK6SZKoW
NTskmh3eouJNibj1b3GpCL7ohmOKqmICP9Pje/TofgMt8TNDjBDcY87ijpKJWOjh2udnWzPSgsk1
M+l72ou/QvTlILxXoJNQAkQi99fRWQ/dodK51hVTry+As+OuS9eEdOr9nDD+G4g/F37KtHyps1ar
NpefrfseDC1q33j9ADhzy205P9PW3TsedS6zOSMmQvJTBEuvB5ZcNRoZqV4TBKXK4r9dqZCpTavV
1JeJRFuicU3VlckFYPBOPt+5grdFNmqWRDhfDyF+xv0jDQ45ndwBndYR+HHWlMnZnHpMmpLgCQnx
Vm7u46KOE4P3zD/J/z34/3kNDtnpe9vaSRLLDmhhp+xi1firXoYs9JpaJvz2Q4q5l8r4ewBF1gW+
VZTceCxslLYDH2LZzcFxAHgWMiak5A20TUd2oRKySHmhTQcn4jbYFQf/ILGRuLiEFehuggTIQMTj
8KbpzY4dG/rH4VhJXUKF9vN5hvh1qTH+ufAXP4EuEF5wKKW7g3fzIy8MrGOaCARNqiNP5QYjowZp
1Owlu7zxW3c1Rg37OdD38BYaiMpC6Hf8UQL4/a8ZNktca4aT6+W/DWtWgzT9MPfHRNKVSRwiIgcJ
2aOEkgQOOCX9qrqUXrbWZxTKy2Utsyi6a8BYcbYq2fCQNqDDCDoQVKkDOOFnN9DzQr7PzcnTzd8I
wWa/Luf2R+h7LTcrzllLaVnazqxXW5Sno1QwVqfMUpKepLSw11wMPIfKuEnsCZb0WQrsLhWgj8df
BA1Fu0Ujfh8zCd7vTLCDd102sX2CRJePTj2qNAdHzUn+TC/R6BiaUupw+of6D6kyPJG7701rh2mD
QOcDM917yEnRzQ6RDkboswyZ2JGhxCO8smKPWViBHE9kxUntCduYTvD+LiReH3ujlr50pJVOYHG0
uWV4XcCgNudFis+hLmxSL/jsLdx5gsI8poLwVicanrzMJDa+Nhp2hXENpWFp2zJy/eRQNNQytwOv
zmXdQwfGtI/Hd5kALLJwMrDrh1y4z7L6rY05eWaYNYGWh76jM8TLQKYP0Ce5scpk+i9Xh4R9jz3Z
USVAkUQtMTP/8a87tXlisdAtd/9vlCHzucBmSuQWo9olgrHnkunM/JR8PHTYUbXGSklDouqOvsSA
fL1hEjPgb0/qMPVpWT//R++a1uYXOS047LuoRMFQ0nBvBworXFd1Y5IB1IUm8odHxAfaqT/pPR4a
dAoAcPGHtCMTJD5nqo5Dwt+CMMMVhHZOjjo54Lmll9Yi72n9eHM72APCIdo/CLoVYioa3ZD+K5Xe
1hkcr2BsJxqS7MAK+65eu4mq1JV6iudpLtsUmi40wPqz1quOl0vvufPD70YYMqqfILPheDgePIx+
03UV0VGZyBGYDwAlBabtkkBmHHPwhfKQOmdq11gLtOpUhd2gCBRWYgL9CKn37qW162GqggcXdYnO
Xz9yv9rApASPqhiCduulWXg8piCFRBhLV5AlWlMQzF+6EPQluutEfbN7LKpGQjYAPF2Zuoo587GT
HsXaQxzBbprSYyu1w/gBaci/iKiL/YLeJRLNJV1rs4AfBuaIHDhkclr/PaG95SwvztuWyTBuxeP0
kPxCHZpaSVB9500YjOYZw2x270uWsmMauUKLnY9IwwnqrIvvx3mIEGjy38FHItr5ZxqqWCqQsLTc
xw7fxrJHguqXahtLxgXiMAEXCXf987W5zkrgUBpYvf4NKgdHIlmVnG5foQPaIGHr8TY5sA3nnJSw
yOn0NiBrAR0u4+qbm5oBKOEwnMLhDW1Yn6hIFfVmkgH309ITGiRRYd/hj4oLRYkBChEdjw4SJsxE
XXPRG8pXiJ46uNIACNS6GvghfAhqIz/DhLmLrlGdSvNdmuDIwbnwMjSNGofWfDEY4p8vH3tpeW2Y
cEuSf+Nubhc/1Tg5DUvAyqCDma3mbq+w8YU615m/y18mu8IDH7g9CNbWZJPFToHo6sCes7qRPrGx
a5Q7R0nr2N3aOAye8KeS8hoaxgQpfjqdi0nzkgOklg4aHRAGX5dsvBVd9HQ2p92yvFrsHZMtkCSv
sDSBwA8pN5qmvsJnn57g/OrHMhH1ufHRCjve2JfPPBm+A5T9mLlWa80DIgGjVpr0J5Z7L3pFkdQe
VN99EngCW6f6EqFDgoeht9+T29+OExGxiYY/MY3KyR6MVG4nB5dF9gk4eJU4Z/8xQ38wdx22nbHy
AIW3JavXS+WfjJ5NJGtAFxmRF7aUnPwor6vUvcIjzOr42PxRheFfhS/hnoqH6n04jfSKV3W3nC6Y
a9DlO983bq+uoOAC/rTEqIHF+IgBfBw650FR0zvYpNL+k2r1VXN6kkUudHEeXiMDTf58/dGD0ewv
pXMZWH9mcK3ZbFJ2Z3sNoghGwBd4YYGEuveKytsYMmczSOT7xlJUUP8jLew/kWLr0vxsVP3oP0D5
Bcq6ehXrkgH7C6blVg8kCYvQdCjSivfGSf+pf5aP4oiNPr5CebVXOPUU6sporh3nstOetgsuo3DJ
RmQ00B/CcR7wVVzJF/yYsBulBvh+9s0Ztm4aJ+FKRLPGFtyo6C0GkHX4b3IwKr/PNeHpWO63wHiY
W71ZVv4pHmGkIob1TXMsZbZGMs491Ezqm7JjxXMse/0BPeWJiCwX8/Mgnm+S7EiBd1NYEd4Vh9I7
61ELO09hJ8kz8FcXP/AIRsWSwOmzccKaQG+ZDOgJM9NuY70amv2gVv44VS8i/RxomATMF66awZbL
5Z9Hn+yvT34C+3sIjZMJ5zCBTUF2nfy6MKluPQ9YF1vdsJta11yp9kUFvOnYYzGSmJzdYP5FetB2
CmLR344hRN10qd5ov0iDmdilEcnEd0aPOIjMJ7mBzyzQJ6R4DuJFXtzKjAIrHFxoP2hZZq1fUsT2
L58TZz7INXnwm1bQUWGnnu/KIdifdPqkzH7xx2Mr+qwFU7baKkeHXEhXeWs4C+Zvimyz2PW0d4nY
gHPgY9uxGBS9JqzeSMY1CDhh/15YGZaDN4MbsxaXW1OHuZ/IBWlNpMD9KdtwON7N7apYxQ23ZVO4
JVg0qi7pVEBEn3Aum4YVzyuSVpqAySLd2bknQ1wwGgoCnGXOo1TEUnpjGXcM3InCSfzgPS7fn2Rt
bffuGawnjYV6ku5+IDWVtdv7CfTJWax8kiOm+ULsvhgWd1TEOp93HOirfEpXJRh2w4OtEFAnKalw
sKeA1yT4ZNj8Yr1OhZGbXUMx83+OPPpvTWXLh05OK15EP9Pozt6RIoo8NK6ILlnF2JI6hvaVQQnG
kE3kyhuOZOUZLbciRYJFykhHezb4y6pkkpWZ7qKdQOZHKwBkJlKMWmnZEJyNM3NFmjEyEYsn+byE
TuK8AmupgWP+HcGngeA43ULLB2qF+Ij50/vId1NmkoFwxi89wAssEcc9FPVhXshhso+YEwRz6Hb1
fTfk/svvzpz14uzzazEDW18NRVdrkJxdzKPACoSoOY90X67gK+E0Nu2mVGFGfr7+YPs1fqBpFu9B
MTFSbBMbDYq0IkYM94ifFqVur3es+WKrMze4Lb5+iMvVfp2OhwL42ZXzgmMKrDZknolCeJY2Derw
aaYrOH2Gf2Xsi1RL+xOsA/ZeoD2xh9wsHWXbZ/+TkZjOEmQTHSnX1mfCeyCszpZEsGXrx8hxhJr7
2yt6z6V6RtCcmZWx35ueL/MCV3vTvRNmKVn5+i6Ocv9FJjGCGrB5bWw7yPfHFI6cHKOQukVHteZq
/eEhsP2so59k/IL0ZRVSWeeBhpLpmACwzzDZmXivxUUW5EqvuIK/kMNkPJdRhjXVtPlBMN3L83qu
Hbdxf5z6qW2ptM+26ZD+AaKuuxBOmJkB8jEfR4qk8VDQn0QIlJ90mgibJslezsys0cgnafEWKXGG
kyYReDGZpiDgZAddHtGzA8WbRp2yH6amfFnPSG5oGfI/ZUxovj4BXHIb4df83s2teix+9F72+cDw
lJkp3huH0bjM7tdQpttph4i74I4J7kX4TeymY+ga1cBP/zOV2fOkaeyXPeMuwf9hwN+LmmsE/mhA
iD8ZigyOoVPkMQ3WXKFKTfk8kkscMq4pGUqAEqdCHAMwFUadHVLdrKL6hdKCGAxXQxh4Br25kSRD
HelvNdyj06mwJfRWOdcipLIlHtc4A5hQ8GfzHsoAv4pskvvk6fIhza5cuBAYpaCiFQTXwD39zVN0
36p8JfwiMzrJf3pvRZZ2yQMgtYY3iVKghb/yocb5Q7ogCS6Q8Cc2VOnlcIWPZQt/W4JbIMkN/69m
ugrI635Ymryw8RgeJ76vWM9LG+YW+7o91b7US2/yKtZ7qpuF3ml4VnRk9Xk9pVGSah0diKvzG/P3
6rXhJJyqO+xS9reOdyQeBLLUFDxTPF3vBhJoJdZ1W14mIQ+1YatTT0K9MIQaweagqroUsDVxzmEg
eAoGgF4d4L+BKF3Vs/enaq7Dc7grarun11ieXuEUB5HjwXMglyhPRGBxDeNXD6UbJ8O94uYQO5fa
5/O50F9ijY6hyW7sGrDmiwJUPUEkD8FdWPejlQ88/zDwLyXhsHYZuQwB8epO3pgSNpoDubWlzaV/
AwS5TuXRdLO6f6IvazCF/Y17l33dRV11yF7nD5T/8zslVJ+g99QAfVj+ZDjuqyPRrtA0+N+M/VGp
5ghQEa+pmVVRqNm7kiMuvaPB2y+Q6erhxr9zkbV1z/4KNY45sslEp9IhCiTunG69c3VbNhJ66/N7
v/RPZpEhYRZDotXq0zObhHPr7SSXZktWIw+tbP1/lDFvZiRLUe4qPLdF8U+BEvWG4hABxv5j74ry
b+Oz0tX4uwxT6y1E0FyXpQGJ+nGBUoCZUV7tunvzEZwViw8q2LfA4VH5OIfZrXqTNmxKHlgQs7Wu
bP8pn1BkeBhYwirsmjini3kQ6KPljr0dJoL9nCPwHcjL2n9WJDdw4nuAbFo93kIWMrRwuIklOjkO
/0aqkK7WKgNGTclpYqnR7gFSIKIDxhI3u3AamyXXguY4RpzI/7KlZizrX8nN2tnS7XEj7ixdju+t
5Eg3yO7F2FUv3/BbaO8JHQJSMVn1mjOVpGH2ax85NyM2hzC10nccXxLAUoDnhkkHfPDjhz4t76kp
35DVGkZtxSlTrulf7P+cPf4Og6tmaLkTe8X/P+CVCSWmy3RQMc9D4wuA0RkdE1cFN9mm2X/7rO2v
Q+EdPQRS7B4IlE5FBtDAwdHCIupi1U/0Mcv7kTeTcbgn3ycK8e0YwcoB8zegVnq1zXpoQ2FVEiqg
UTBWfKsTsOoqc9TfVVWnDewsLz7C2fgygZxLxqwVEdseYfRdpz+ey6SIUMU3dsfd2pULP9t6P/bc
xcn1cQZqKgRg+Qtp/2ybOh/B7o8maEtMLE2MoWP3l/oFORv08A9UpwOowGezx9sIOINBE5w8Yl67
q9rpqMgXsoBxImfi2CIxG1fOrasJVnf6OQmJgUl0PhKpwk4KoK5X1f8b/WPfKB8Jg68hEnuLY4LG
Fmvc1RfOxRX/b3meAAhwL21mdCRgZsWXVE6BGCmFlV11jwY8XSInG7Z+xLaUAtMnhAyjm3zNMqkT
b8kFuryvelP+MDCCaefHGa/dSnLRUa8nPo+JodDir7oHMeBGxCUFERyxZL9lc+PP1v2Rf1oaOm6i
tLYuyPXzPtDZ0Fcdwu/HZotJNMkm1ECjeONREWzKA0VCYo6bFo+/6a3NZOPQ13qP5CDL1sxtmxE+
VyXUxzRU2ucVuSazma0u1dFUCO1h/B5ly31W3wY9+Z/oPdf3iE1KwozZ3zO1G7sBY7CIUW3cJqtU
/wbod6511FFQnZxuG55E2fGtuI++2ga/3DFE/k3gPvbRZbFvjo39TDxivTGc/oVyyuHJ99Ugiaol
Y+mIqWAsMiUC/YW71a4SJjlpdmsDDMKTAlCfWOFBA+PXu2NvDGYehxXDmXT7d6jR30nVDZ2noHFX
Oj9j7M5+flTHJsUfVkKI3L+CwWpjLhPCYrK6bNH2UoARUWZ9bADHJhmRjMu2ho/tpXFMHR/Br95Y
KLvGbyHGf3duoTrzDnfUKcrLO4WRvmiiKE6tmbOgQc0W6Humc5mzpku4g0kv8DvLGv29lqjoh3zW
cE6h4VDJdzo3bNmrIzZWY0RVO1QTQS55tMwNHnMXgXaCmXJcrfQ2XmlfQlpKIxxVNSRSlq2dhJ/t
cOfYrPEjv5bhlHsacXgxXo/U7r72/prucqFgFdohxLVQwCnGecZHWtzJwKO51HiHwjbbqtqjAfh0
oCHPZt4ySDEQsSby0SOpNDlwQpM2Jg/VOZfyXGaaKIcsEOT9J+BlfzsOYn3TMOwKGVMC4H/PJKw9
BQwACD6fwOQr34ap3JNJD/RVEHlgeL66j0wqGrU2ql4wkRpppUr38kR+74TKuyVnNhIcsXQ7COo+
Okevt0esP477lKdFvm37i7CTMUYsUDNsF6GoOU6CcGe38JBLZ2JNjpeEodj6IBM8AhXTKIDz8NoD
ojJiyBP3T48vD9N5HejKGFgn+rl2skC2+DELroysxd3XzE1AedFWDKCXqkuttxOhLJWq0gt3/VMa
C31T5+8dix0t5sn9kl6wzBxHaH6C+465z6wsFBfMJBqgtMxOMPEH6g044j8BjbMXOxsEW4axxmXf
nROAw8spE/hWIExxB4I/m/tPBPjvvgPMfNYOLgyrDjGlYi5xfwrTOHGJVD5Q9+irK8qMC1gftf9E
el6RKKDSsd/p1qHzWsHiAkxiqrzAKy0g9Vfg+SimImqvno9Wtqras4rVfg08YyusmtFMxdcOdxPf
7DgH19fAne2CGUieE5Bchc/NR4kvrPY+UUbpIAuAP+IwinewzIw5YnjPZAtvup1ug3IxyNB8FmlA
/SaSgEUPhTImjaf+f4apaG7VdcfPr4ruVXQUGJBRIVSnE+GVzqVVDi3fhi6LleMx1haKewgx++V9
xbuOL/0gQHtHMwNW9ijH5xKlpXm5JyA+qYD/7puc7+nDX2MAchnf5hV4zDhg+X6VIBmXRNiBd6GA
eXxc9pHhdvrkuGiRSSzLDizBvxlGKbrMALLZL3qdCnSwummAKCUWw5iKfsLeBl261vSdc1oRZY9J
75cVVR9PQ3RrvQ+OeGdqZoWoWXZod9hrCt3DsoYKtzZRwKbH0KSCmPYxJnP7SxWSctCOXtMGqymC
PlTJInK/qyKn0RWSfrNzi/9IrUKUOeXy/cqaIXa/6A7jLSLnc8BXilPMy2XKN3nSsiiwSc3e3SLx
j+N6s6YnoCeC5pLsrRM81QHmu7m8CcNbH0qFOHZXTqOtQ6A13CeLdgfXZ1DsXUcq05yfUA+R+EEx
wG/vLORVzCDADEd4FOwpCvDYl3bKCI8UwgYFRgIECHlT0YQvIvGi02SBFoaukF8xnLP0iBq3XpSd
zZU75P8sqkQxBDLjxAXILJk2lElAOdBk1bszncxOJJClo5hcFMcNvcGzUNMFaFS8I2B09qewtc6V
Wv/0izf9OJec5d/NMdCBg1H7KcoIul+i2J5Q6s3pY24NSyvyhP1bb/N6a1kfIpoOsH5dfMr+YPkV
cEre6+9Ta56nyN4d0ya4pp0cjuHcY7NvvUD/AZXFEksysLWbOo49wbfyrbN+TJPkE2dgr7ot7NNc
o+yXzsqxZmvAvadWOiIdOzUOfvIZMY/GqcNBvzXRwmuvbrizNO6OHZogXRV3NF/3PHu8TfQQgzl7
1jkrx7AurfFdu70KtKQOFHXkNMvw++lVqQQq2+oplvkvGEiyYSZO1SFzZyhu+tcvsGDjwe0aZ4GC
fVQGzTc+2lJc6Mc6zE9cEk+mBfd18rKSkEVymXjApJuSBzkzpsx4vpSTX4+nF6hFFJl67q3vjC3d
iHvdvnwh7qqEoHxxi4thocIuhAgSkEAzrIVBMA8nVu6F7ZCyEQDyLJPbgoUqvilO0wwi9KVeFhXb
0tIl1AR9UguR1qHvheYdKN9uABy+ZAIotnwsBnCFzhM2GejuTZMmPpCLK89AYVi29xEdS45rwxfP
RC7hLQzvcVmJTCumk0ShFVP27DHMJEmYEPOVL13X+k39Q/LxJbvxQ2JBubxOB2rdQHXyqHHFGD+k
JQbkhCD2yKZuI57C0NpT6rbIky9Se2sJessSDBB60+S0tZG+OCfmY1qkfzX5G3L0eGt7i35obA8O
cGD199SeS7mM7QhThQjw+Pleo9diuihD8BqIaBs+b2IYY5/jxeNGHyLVWbShsdzAwNKQpaXgI5OR
HnQUGRFgl/bcDDVLgIfZQoJw7WdHqCZ5y/1ajOGzKlcBfw/aatZiBem5NEr5RraiuowgURJYJuVc
M+RZp/FRAetpedHbqYWagLcFtK2iRQFT2ePTzUrJoP6GV8I3bg+iwLFbJU5342U1FGPqsXm2RpN2
GJRZmasKmIVimQ9GwtnCTDcSxyi3coJtHiDMFOYygeWvOEyqbPInlBgh9L9fAjE2J0XmiKmhCe6N
g1/Rz6vWl/a/0qB8y4t2+dl0Yf1gcDKbYcRID4JnTHVxM01rCjVmV7Um5qH7/bxnGCdHlPNq5+/h
/FPVMu+GmFuUhdMPqKWNc/bhq2DWU1OVssLkngBLlQpTo72nDxQI1uknS+4OBjIsF00rBqY4keHr
Vgc0+Lb5WoWvvTxBlk8KeiDq606YtlnxAcNz0iZnKgSdNUnLSUNoNBdwJGBq3gFff8p4YGt28MF+
fMUZYz+xGXnrjjuOmO02zgLG/YrIHY8UViW6L8tHbEKEum5G6QmYRDxfQWYPe6PBgL3tFI0gYog+
EvaRS7QsQZKRfaJTkOj6BOuQOJQbRxxhgE+Z8mRSHQyzpTqNBzRvf7OApp57vtlNRGDjl2srjZdx
aYboZkaeI1qssLgc81rGq6os+W/2wf1e+ufltdj+Fzg7xprnqhgov7XFdV6EmeBmwUc4kBEn880E
Wakw8ewE/wXONTJGPeyMAs74ENMO8B0wykEsrNAkxX8OiccZfymRk929o6V1o6dxusgljwOa3dOw
dho+ixsdjycdGs2HSx9c11jq8y51nE/XbfXOU7NwBCz9xPmUlEU/Rd4eD35t0QdXAV63Gi9Oo0w5
BEwFWwI+/tMKnb9xWpneS0hTk4+l7uRDC61v2PPUpl3K73GoScrnXLsLjxBx8VMNCZJWR0P44hUw
CX92iTu6hEVzBQVW6+sh9tJNZIEpcTsn1O/0W7Pi2+bTNWc5UbkUhFJiRzRObg+OvbmWF3vbpmAA
UevQJZfLckC5hgdmA+9jUl7FV5vw0Z9/70Ko9XijTMNrTrICEhEKhaootHgHBavWIhYevSSGJnlu
Xfqk1b/+hLeKkll3nM6cprLQegSyWx0Rwkg5i2943bn/EYcU9I6Je0wdPRDZKKU0y6lwHGXI2bXh
tEF0jLmluhdIArFrZGK5Q96F0k4FqqjP0XkqOEizbzR9bQgOXST+0dRATOrS5jJjZlKFow7VJjSQ
qw/ssirySIOPQJx1L7OUn7ycjViV/gPfNyZfSXmVJppENc/GlhQIDq3viZhmH6jekYOaT/H8YO0R
F6xz06JgyyMyA2EGH+5BwCRBexLJzHRqPoYEiOlx5kkpI0NIaDd/EGczaiBmqiLn4QYYTtis1dEH
yOAnvglzvE75/+itQDbAqM6pQbvFJm4MZ6kRMPAWORz9ma1IjpQXTaeGqxh4F5Em0kQPQPj6MNlP
5kxYTA95SFkbxbNLbTuq3AjVI++BF5UJqljUtU+D1lVxxTuiSOyXPngQsyVZCVSOM8PfMvTQpLfH
+AcVeC/98jqo/SVQ/vujxnOJZ8/wd3X4LWsQ8MzfFxasrWKXwqDHSNk9P6zT9rk3RNWnboWNXEL3
0jTEHbJ48JemqPbi9+GWgzJ1XdQ6/I/DqYMJTfTQjQ2HEWTEIR9gSeZE/kP+q5dTgM0UhtxFuqZs
lPwoEw7btCKQ8vr8wXMj1QLnxMjTE8hqiJk5h3FHR5tcMrgEE6+jfeO9QGNU1s8VuDDdi5XNCcQZ
yBIdUmXT9J44nwZtkFmJ8BjENs24riJvSxEkPozebg6KlScluuBgAO3e5q4HUcxbV2Ait8Q0M73g
YIvZHvnQbSYXSOx5SbLTnpcEoIIZ9lnj4LMf1K5PZ4wADgXtpw1ulZBV9jb3A0TRM+ZBkMQ40Q93
OA1/oXUkSfWVmgQPuuStqVZuSc/kqbsJEFi9i4tPtQOdlKxyMDp001bfz3J3RQIYGvPPS61+HWIF
itp3tf4YeD8X8sqA7dXRn19xQzj7/jDcyCRHAIyk8zj/MReBlA71Y2vMnm0+T1338+ZZ3KkXmznZ
EEH9Q2BG4MDFgepQySzDARBbONNHPWZjG9aGLwfwJd9rKEZtGWTE/4ei8dmSTQ+wiMeWjUmzGGLR
wzsZX0mvSAjRHRpIHrG1hHBEBpsWmVG+ILzHs9AR1dohT5o/fKxwTpGXrDX9E9Q8s15BgVgFwMdL
h3EYh+7Fgp4iOPyCif5HnZRcBa3Y27eEC8dQtpZCN00ObtHqbcyv82khvZnxNNB8gwQB75EAEheu
XMBw0YcyAJqt4eqCQSHn6G98z2MEBoyXfdjTKXfR31kVcBoZrnsh/n6FQGvQB8w7NsfzaweoblIV
FUlEx/0JALIC12tYGQkWW17oFWNzJkmqUwGxTi5vAEVn/nPEgLK990qeIThPht6yEEZ62wFdv20q
gZ9tlUVHQhR4+gWlfXqa56FBoVEGCMuFiQaIcW5Bzk/SQj0hWahVrQidymQMyEoO3bZ1uCASWZ1+
8xTxgBTs8qgJP9DtXAmKn+mYbBScLoF+i9MzAhFqq7egvIKXAIJVpqkmqVXH7qF1H+3qEyuilL+M
BABd8ZLZ2rnj/z7818HOATYfbYKRmr+oT+f44xefEhKVN2xMRog4D7kJZ94BEMJ2ppq6ysRF65St
8hOnATm0fjMxEvut6If2UZMLI1D36mJmls1BzhOxuwW8mSVKgMElL+rnJeZEQOHlAJSUiBR7Vf4R
iLn56mxTde0LjKPR6GPPihqC+wMLxHlu2+MLNrGbiABcRaILY+n73q92D6yLvgD4tWgt3xHMqg6H
e2il+JzR/7gfc1wdgpieGHdZZ+MXoN1A2mKej2VLtPOvhdV2E9tglaZO9Niyss9gIfQk4v5aoi6Z
QygR/0lIpFBikQ8SyxGyXSSaLVfl5knY5T01fJROXg6oj61AmFUsTqydPnddolKPTB/9Ae1mqs02
sejgtZTHOba0xpTtLPRVlJA3rlYHr36yqtpJhwTYRASSbqx3Sl5De13lafHHj6JELN5jYO5YYFaR
lJ+6+uk9AQPwxCINIMxcdXvOCatGSRxeaqeVKR41Xz7Pt6XRQrVcpQhK/nBI7wq/Bzoy6MnOvIk8
HJ26D1cmORi7KqHzSW4TG6X0e7vzV8gmVycd6VHE8WgaexIebarDlIRzSnAcUi/QqqJo8xYZs8zv
tqtwoMwSdbO5dYHVAngV2EvQ0G/cpxxIJyYvAOgW8NmP+s0W/aPBVPi/DMXOGpxba+miqDRhn80q
0McXAfMspwH9KX9qnYhPiyeufZgYZzTWQRjt9yi6Xyun2BweuAX4zo9qjnvz2udVBHFlnu07z+Ja
WK3Jov7AZd8f58/V0BLJTBOpVkqx9tZeKvnSW4OQZLGGQKCjgHrdH7X+1KakN1dUTMEugd7NsncX
2T10fJNZvdUneLyluxaMb8J6zGX1P8vIS8rAiOvBmkGjut6JfMnM5d8Kg8oXI4Pvp+KhSOecFn/2
nFZwhw7TA1+TjbhWznSnnbTVbi6M2PAtPmzF92DJ8F0pky+sFyMc4qob3O5X58zy9SfOeCmR4GQE
zfhyY/Bq3Nn8FuzNBqfrUwKO9zArS7cs/EYzkt/9/lxbeGUt/COWp/J6PJ8eZ9eaIK+anNlgXozA
/63B6RT67SmT0MrqucSHYT8DA7zgbXqvK3w1LXIz42U/tEca+BzqPY1/xnXOF/EmT2nH1ueFs6vJ
bCTCnwkUU9yrvjQ8FJQftozEQLPixVkn+evABsTbtPj8yWMMSi9h/WrzB/6wIR6gLB3pU0054B31
+g5/gQZLbR30XLwYMbJp9kH8+c+z7hJZ1AjWZpfJ9c0WivHrmtYyq+9hLw8UrTIC6pbBwC6Gqkb1
SXzF8l8lRuPnMOBZkP9KrdAUPk7VtOICTcdTZdK36P6b1b0yxlhhdUka+MzGMiGFY0BiIcpOKYIg
bgfmIJ3CPJHrV7Xi1wd5b49/YdoU60ztTTkp0TJRgD4xFks4pztxmnvFv92J0yHK6SLdFiYH839s
0InhNGOekxJa0jg1vMH7cQX7q68zUZId2oHZPUY6SLLWIs6Zl+EzlZ7KrRGnQG/PQfWM/xvDNnDM
QkyudPTICNNLvnST6VYO4TYn4J7EbGP2flkFjsawxbVF686yH6IT50Qzydds/3XuGoUuiHY8eRCk
WNBa7uZGMmEJyO5fURUnOKoPUQ7Kc1fDtcYt7F1nNYamhpVjXpS0OkDID+C738KFpp/XS68qhall
prw/taRjqA1iyH7Ggqm79ZOddILnWY7jwJ8WOjWy9RuBeotXvWrNVoi22lmxH6nNh2Bs7o4f6UXC
EsT2JzusmkEDK6XYTupfzytkFASS1D7IJaV0rXdwRwFRPPSK6wjzDu7wr12JA20i2D9Cseii+yvY
BpIcCnZ87uCnzm7Ed+KaR2F1MaIzC2xRx8q/GYnHreLumS46v0AvGW64WzNtevZv94XQJeOBNRCY
17dZ+/U/mjngsjpHEo7msCZy/MKWR5YkR3z69byN5hwvCjTV5ip/diP1T3uAdwgpLbqRwYzf4kpx
Kz2JKTAwOfRODB3s6+8qFec6E9eBvETp3QyjWIZ0HePgWQjz23dohBH+aS4z6OVQ3ZLnsPGQVEpK
ldUFooMlVmyWwS6AxVfK0dXa0mrbPXQrW1iQm/w86qSbqP87k4NOERvIaEw9UMgSGkroMLCXg/lm
swgl0P4YJWRXyxIxWtFopRwcOZZydxEJrhbuur/Ra5CZQtRXIxgTCM26ssH4Kku27cHOJkEufgWB
t4KiiyVZei1CeALsJoqB/JaYV8eAGGrx1Mmr8vza2snCCUFVSaKynkFGxpHeOo91jy8JKq1d3TZH
seH/C8sNoXXIObX24j1c2E1FgLyGR+l3L3enMmrRYd97dIHjACe6n3aYLrZvN8Mp0x4WwL6s/Q3z
h04uuRcIHw6A4zYSKOeXBLqGMieHXCBDLQ4WTZ4xkVjhzGG+Jm2Xf/4KxWqIObqKG7isjwzvz0Kn
+Kamt+wdlEEJHqM0BJnD5tLmwv+YiA3P2MJ4DCpfuMtdKi/S/pfW0XlVFAm+7sOBSKVuX/YoXuw/
DWOpL1LlPxDKo1yawIZkoW8lFA81yLLcMWOEkKvGGT9g0GaGvQ028BciW7yjvlLHJsXZ5MkNzUQZ
j4cWMs3eCdBE2PgRW9dM3NL1EGFZ1qcZ/nBkNNsY7jCPNRdnqngbHVTGrjw3OwlaKuUy3gNI+VOd
awVV0bCBYSGY00ZDmKJy40YNXthP6wrV2D5/trgq8iji7BNzryP2cRxz2Prse58tqcYUSSdgXcDt
DMr2oqzJfvxlC1OQqiDdvze6D8re+gfGezHJzMLAiH/auTZ/YyTRDTORBicVqLthMhONPosyL0TX
aBs2LAEQWG9N72XqAl/O//bjIOql2fVrETqZC1wWDlJ/bWXP46op5BYn1jMnrePKF5G69FknO6Ns
Ep7WBD+TAcW1XNA6EImPZhKyMvzoShmXfh1fqrStN6F9eWBUzoCtexhie9kMjXHdgcJ2oPrECZ6N
TbQYqS6xLgWLxb4tM+3SaJZwlYSmCGEwBXXQIxTbLYYkn1Nm6Pt7oS/q8kaoYIqgRezjqAM05w5d
5bI6Ifls51hjHu3n80yjfFMEWh9yLVHpUNpKL4qhyURceJQhjZ6XSxH8gYoKe3R2OdlDM4g3NnOM
f7kfGei4xXqbEHVLgFnxM2TBOE208lFTb3Y3x+ZK/Td3bO6NN6MW2yG2kyoY1y5iyVTBvbZz/fc4
ESMai/jn1BVXjR9mr3zJnlIOOmnmcniC1qjlaQtf2TYFS79+z43lDmK9BZn/rpwZPjKarSeak8Il
57K96Sl7EkPv8Ne1Uw4ZJDhxi5Xh2OIP7VwxO4zlXTmCDQ5R9dX6p6TedqVVIu2HonzqJQvAnfak
JB+qNfG1q/u+fU+O1YPLUHS8G/waUhPWs5rQUWHe1KetpBl4h+z+TZTjfVdTjdWyyrdCwJxKBGEQ
8DMuGF2up1vdJZ1XPElPN7Me9VgpPdsoSR6roPKjWiAHPDTMimdgoyzpHJ3c4Zs9AiJZ2xNMEJs2
dClrQ0yg+lW+eP/ExMoBsxcMFPEFi0A5Vzyq+FQ3jGgL5tIShthutj9R+6TzBNZSPlXPk/q5vK1R
H0tGUvR4CvAVeM8C5cNlgJq+TDM4U83d5B22SJmXz3/Rfn/LuJiDee6MZjqV6LjWU1IG0L3GOvBJ
ZRIxrMUo/FVoGks5jIX/35ULqEi9svWftHdrzWRASJ4k8DRq1jDp0MRArWtxh0nxgF+t+X3+nmrI
WwxmhEuvKGZGNAWF/3aNgywpdzKavFKhWdHrDuwlXBAtoBUqDY+wBjqyHv80DpwUZ8MJc6gAc1WV
oI5/RDCozIluK6b4xvd1BUQM95YLPFoZmtYbdySY7YI0OFUoTci2bGiVPZYLfsADGlgyK1BZAy8s
DHOvhUo3cv+BDkSa+W+jE2Z8MtB7PLXtWQ+846n5SbHtMWhyHedBUtf1VmXVJu1lsGwyRPZy+nUV
lr1I20BGov9pjdZZuXJfyrp24OTk9ZMM6RpZWxMzQmlONmxrP3FfkT7RBkbHpdSYoae6L23BFDrK
yX1dlqpOoSbfCJhTLroE5WwgJFzdICuFy5oa9Uiw4KmJrvtBAGMJibr3LJzKixkCldxqzoakWU+j
Mr9jeK8aq/QYYcldDGnry+YKz6YC4BqGhqSMpQGM9+cQOnn+zWDdEBxCvoieR6v/mEBkUad8m1d/
5mFQ9V27MgPNSst3tGPW7I5V26iiFkQBWBTjsTolzFiTDU21WJ3BHA9PMvtA/1fhtiqkGGm0ltFP
Sp6UP8qN7vfQnTW23edu7kpm0wlu541LDsU+q8a+YolbAF55ecsSYWhVK5onxuBc7caZNWqMvU2A
oEaj/7l3SznRil6je1Xn2KJUd8uezACGXUAKcc5i7J9pSR2NYFsUorQF3SN5fEr581Ru5iQUtSsF
a85nwBjEuiEICrsBd60F/HC/MitBYrnMCDyiUn2xB5gpe66vaNujFPHkFlP9Ah7Xv7n83dMqhB/r
eNpj4MVMlCVbTUdvQGJhKK+xTGAsCPWOWl3B24p09v4nxQ1P8lyFSBFhoJN+tfuDrfNLoZTDUHRt
gnvtI8mVDFg/CivhRY/ar+hFP5+qBCQme3FYVSTi/IC7BvvBgnDgNOTCAmuOE7D72k2UcmlKQ06n
wO++V4KUukA/edF4lpscWoJu4BsidP+IFFBGCU6qSCl+MmMYGNBAep69PkOTMkdrTeE4CXgG7eGw
iOfjgJ12AlaHBJjyfO2QPBqgABrSJedI2Zbmzgz9eSMUCS+BZIyoQKsfxd4pb7b+zrjXfGRUrOkZ
Vg7hckAAhDLj36ur06XlCzUUFbtAEER5Gv9315GIuMmuc6EKiPLuM5E/BxEldVuuebyb4bKoTBEw
r4RLcogQtFQH14+a6SZSQHCFdPQ3WGdiZoETvot3ujhcqaqukVE3OIgKertH/KWAL1722FlNP00T
Lx6BvINn0KdjOfv4yA+3E6ev3oC6Ot+Ug/CUtSzwpWf6hAqVxVLqMKncwuRTd54iqP7knR6HvBLM
mkqr2X0tSLF1RTHpEIAmQtxrtEtrjlgQ6vJLLpsPoMfSvlNQwrtpPUuPm+CMPZBG/2Yfej8dZmDv
LUUCD9xn5f2b7BNFuZWEdFDdr7hNDeuWE1uR7jKl+N1wKz0J8NdEnq0SK3DSAX+T0viaXrQMkjWI
iCXB7c3Pu5uXyz6AL22RS2uCxoNTWV4XpcP6cyqFIwmbk/bRTgH+bbc9SnG5WClBaYn0JoqVAJVp
ooWNQa8bYuiZMy9ZUWC+afBx3owckaBK1tAWaO5xi19k0obNAbvn/460NzrlLZaeJImsCwEZGoQ8
+h68KW7r58L+5nbAyjLlXzhpQSUUi/FZpNSVYQdGENBiSpcWYf3ONNpvx33KVIta+Vj/Lz0lJ0fJ
V4Sxau81O3L9Evt+46owYloDkI1tBIDQ27bYTjW4E39vL21Q63G5p5PelTBqCc1xZlDC5DXY1OWo
KzqBUMEyezLdRLMQ/i+nuu2/w6Q/LUdHJ+G8UNxD9tDfT4GnXACtnLtbdaKSQAww52UobpTh/umq
zAhufRnuCWoevk98cwOiPrprwt08Uhd41batotWMmdGNL5cgDK8Nm07pCpjvARaGWyf/JEJwTIDC
fqRQ23/QY55Ezo3xEjiilTVmtd0gRMyWRgixI9+DvO30FCASic91I3oKnAMe3Feg+4wl+98khAlf
q8aUco/9QiAYvUO205SyP30qT/JsLYhuzB39CUnlgncgb72BVk3Paf+gMrO6IyXp+Yqsnlys9OEZ
YEyBCNyks32vT85PEMhuk96lLbOIiEsGXHJK7XW+gQu2uXw+G1BqZbAar+z7MoBFQjsy4hbVOrZl
7bnsi8JGYPmsJlTvYu61EtXZH2LYXY03OXwBg7XWh2qjXZHyk2fnpDP0HEZHVP2VoahAwlQBfkmi
xPjGLdlBKYHKJ6TMfJGqp2FalN05MAPn+LmfqJjIbHG6rZjAVJ4OhnJxvR/FAKH1BwlpI1VUArxv
Q9Dq41EY6H3V8lTlNq0uyl8gE3M7FbKSybBKShp5GvI4Rlm3W3IbnYzNR3E1F4SfLx+gvJLIln1E
B54loGheYUftrl96gLOboGDmCo2OkbKPDGDF9lSUxuQO84eQdiEUfBUewXAVMoFEUYoShe+evwuZ
/5EDWnAfjTRzJ/lKkEpn9P9NLnUYgC7FTwHcSn2/EAg0tIjJ8J/HGU2Uc06qqXThQvXRZHrZ/wwk
qyVNamMKxDUyKWCHATS0+i3a1UgNytKQNtySzk6HrtAUN5VP9u7ULRy06l9Jis0OHRXndbQgrfiE
2ckt1z99MqKvWtAlp9kjU1WAKEX/DblUbDLzjW7xOfe3sAfGqpG/pdKNLc2U2cofiLJOc3Ni10HS
VqK0m0ihTqo9kzWHgm5hVuRQR5+iXETZBGSxM4KEC6C50hFMwCSty1L3Rwof5YhlWivLrj0aEW9L
n4jLlgvWCGLhNlrG4c/UQaBD6yixLQklgmm48krDFpPOlsQAQDHN5tbIbqiumN8N5Z95taq7s2US
NKxJUJeg0yEhdOvHra6AK11bc/YKSCnSMRnZTkzALjttp2EeugDyVqjde1xrVFrAkIE9AtNyU7CC
fqdGfPa1x4G+WFWI94g7FID4fvy0G/Vm5fElCuAwN6mZ4earoZ+jgeFOENdOfAxHSQz2cNt6OFN8
lmZim8CMnF3c+l2lhY/dbmRXKoKQmidrXO7tDeP6xJHb4hNxw+v106wLDa069Mjdd7GsHhUzucMG
AO1U1B3WsOiRNUarkq22tpFsgwRxo1zF2GDvJmu2n0o7F3aCtnK1X9V2Yw19aNXhimcggE0eN1uY
nFUJ9qxMAytwz2Rymh8pM5EWLAGeJ9zRXBXdBBgRFwSb6d9HGPCxqCPTtpViWXkE+EGqnwJhiz4y
LQh88iaQLToCU6+hpizYUzcRlPVofRNL1Ubrzkihcr1Q6GeWhxgbI+Y8702qSiIi9wBkbADcFcUe
YXRUQBeOJhYuNZO8eNRMQAxAySxU0s2gm5XuA3XpqqAEEsyma+H8JYGdNUCDXfNaEEMEjfHTCkMr
N21XUuwIYEYK41OeUlvpf9aJIkntasgNNgF0Z3nj4Zx2FjPl2wDQ3W9GO3pyDpMGw/C0tJmsANqq
2uzL6/SyZAiqvZCkBO/7n3Ud3Kl6nuUcsmYE6Fcn8AeLjlGidW0d52L6NYgBtoJgA/XGWRcMVIEj
AqzgdPLZJrkQNLqqYqpv3bUfXunrOAsfEg/jT9U2qt+WK52tuaCYXd5pYT9FILie095NXledvDE5
xHJH03nuapJnW9SVyzcrBXUYRci4+uHEAXgSd1X/uUmbZPFEwCUhF8MeRDP1AvWVujdgDJHsHBsi
hNgY4BpEpzk2vka008yONRHT+Q83kTRFeWMsIyAWVvaK8YeRso9frZjiq95SsSIbD/T8r4l9S7Nn
XJu4eO2t4O6NEl5AX3CwpM8cH7QdGX/Xhh3BXHJPo0nj6Pg1vqlCa5QdyhJf1KuRJIXF8yJcvGt7
0qeOtXCOFc672dPVpBNKthlo4agGz+9QnzcFLE4rTSu3DQyKm6SkK9I06582W/kkk7TOuL8b6fSq
zGgu1msDzNTf7yrgHwsYYqcvFt5B3qBgXIYiwlpDO791pxJWtu5rPQd++rK26GRmMPVZP2kk7hC3
HDsgmBtBem1hugvhDPd2vpd+QN70dER0y7REKdmhJEuTeoQPERUog/ehaWP05UitOsqxBjEKsAW1
VLfIuStFBOnAsnES3itmGVM1K+p3mYv/a+3BJRT5Jl0/BM6naFPsw1baDD5dMs+Rq0xxr15Z1Dsi
osy8tziXcWvQ0ZA9geAyEcyYmA7QM6Sj/8Okf9+VzIyOVLvM2u02G45dxJ1i1w6NtqlYOZnURuoI
ZpL2F/5dyg7kZiQlhtFWf06jvHg9uV3hvRqkhv0GW10GrPK/uyNmWouDgq4yOLDi1LohAcTCKZ8w
hhy8A2WqQOdMri6GGHAvuvtMhZIAJDfV0gjtqhAG4gc9bY2VIinr3wxKee2V+IRShoBGzEDrpD2q
TlDVRlhU0S5Sl8zu5JWtpfhUfZ80s1PEOwPoK4DETOEO7Uo9dEEr8m+Wd2OjmhEsqdgfmX4S7dSz
02ulnDGtpYZcVt/CwlFpTOqTZUxdN6UteQo4HfR+geiD7EilB2gIAjGtY01Lg5XwiLuwVx12i8nm
wBsT1rv1RLW30zTCbmeWBzSsB0573/g3IxLXfCg6FeIkyRmRhJh53OFvzU4tEZdb+5maKzgDY6Bp
8vb12Zhg/a1rIUPgftRIPHQNHrbIvwbRbAQdvVjGs43gNvwHvPXJ11UB/JbPDtiWCtRTvuoVmMom
CdSWyP4tEdFsfwhTlt3JCQvc6x7nWRoGuX/cCwhh08/D59zn/MuWlUMVDvvnKHinl6iZskcGmmk6
DLfjaK8pWQhr8TSn/FJvA9I3FY4TQbO66B62cwJzKef4lvXoQo06mGdvjZK7cFE++GaINOTw/zTa
t+EjGk4MD5v8gXcf93cnhAzMpWTwxuXAJbLB4CralAZ31lcN7rwzORJw+k6CeuNs/ZkkeTlqM/a5
b2ivzVG+tOxmNC3AX75mNiDB+RY1+ZnDuyT2al9a8fMPqcdqsZsu0UnEYcqx0DZfWjJ5FWaOgItP
GNEXc4q6yhksCpyf9Q6Ohe5xE3xDq4VzbwViMguxKirm5u+alo4tR6A4TBGJXPnlJ7oNGVx+pLzR
beN+mLBp4BcC6kAcazNwqFXnEjaNQy4hZkZtsVls25iWrpcqdHIrBsf9QXZguwggiqB2Q2EWN6Il
G6shLOX4u8NeDqPopBLutX5W9w4w0YE9Et4GE/LDwZatS+0UT3D7la5Y5VGRGPXudCZwe40kt4Y+
ZCY+IzdxHssn7tTv3DHfDBakbsmPuUlB7CRcGjqe0ClvF6X4zG/5EaeVp6qFuyIpzHzidV9QzFTw
Afnedf8B/Sa7XD47fON6CsV4qOw/gs4RF0/5NJ4OogOztqsEqsSHJqGf/v2z1DHjZyZRXnj0Z48x
GyIB71rGpPQ7tw8FcYNuT0rbB5Mjpu0+H05gPIddS9Id1DdlkPSm6mlw8z0oBs7s7YjY6J4tP8eO
1yPyfwLPhwy1BbUZ8HLN3n2L+R+acDZzphlVgxfpjkaA6BGq+RWjcilw0Dm/ZjbKc9u/R18pXGvz
bOAUhqcf0JldGDO36N/7e8W5ejGcUMN2I4C3z1m6h4PhDB2dyxB/ncIyyl+52dfcG8hW8ACIHUjI
5tMG8hZ0gq+2T/LIluDjB2MTMZUPZFMY0oW/gUhufvFLXW8PLBeqtq/AhEZjiLrlg8Zhc1SqlYMJ
a9F+ikFs8U21IrJJQMbKDyTXX9CWzrHEaiH/4tL71ac8Ak72aU30dLIGnKvlajNxj2n8ZIhUeG0e
vSXsIi/oyZYW6eujhw/hXaA9+RQAUZ9hu85FLTBXTi4r3bmjK0qkcKZbL8MrbDfH2cUUgsgus2PV
2/P/PtUgXVUUJI55TxosK6U23ledKZxmHSV1ewMFI7EoRmAo7FCeAbtrmaEDiRkhPWQ2nVMyFWBX
8JJRVN+SjW0Xo3TB9DtcHj26r2vod8bLwA3/GlqPhIuQGZFHSRFg41ks4TNoSURdmlTggmwW7Fsm
O1clOwS1POdoYMpExyx+MiidfRDajFarhrYVkmGYCW51lwRibu+JyWBRF/v6eGoBdyk01P+ClaNF
1jM0LIpp0ZqihPCmM2oTVGGp7rnFJwg+u8iShEyIUrXddAsAFhNk6WLDnu8xZMHqlsDeBWbMAL9H
OlEZgpIErOHVlHifm+OpCTFRKvFrIVgjVnQYvqVFiUK4kbFj1BDQNeZovrzW3pmLNBDlU5x+YLD8
8pGuDaseke8MY62NPYj0lY1PV6W+twKif/fbLQMo3j8RMw2c91gcwLcUmpd4vRl7aT0ug7BX7JFc
+kvp6L7Vyw9iYgyVa1Ck1XenJtGYvx0o/yzFz95E7rEQiyeg4DycYUn3F3yNV4AQ98CiAmO7x9P/
0eoREhSVnV2KtpzvpARHBL8G5VSMWz8tXyHGMsckU89YseXDi9anawppvY9gTmk+QzZzdmk/kXoE
qgYQnaIQ9weK6/DvMq3cj5qu8l9Saaokjco02OuH5GyBxo+FchuxcUvfwwZpLT0otJbWHG/11cFo
LzDDnTtfQeovNrZN2SW7iNB29lwmr9K/LKUbjMELoVdK2hDUIPfQhtzEwhxJ4z4aNpqC91Zg/P+q
/Wi2a3Qk/FNAqiMPxnM91uHy2TYCg9EOPN0fLWibXkh11nW58QJ3sV8Kyy8wYOm3mxNA7fI2KQvQ
DqwRw216KyauJlq+zDQPAXHZijmoNvKOF4rDFxwwC/s6kDrh/YQX+QMY8Sj/hVMH07N40hLwrBXd
ncSScB85BwaOomSvNZxbCYqjx2w6lWNTPC3tTjDu+DNOTdKuYhVyDfeUIt8AneDAgSQsfaqxM3Lp
8SLnedRkotfvzFYq3CeufokROECMp0fktgbbDYL5qxE3U43QBjc6QuMCzrtcUf32Htmkvo4kleyY
DJjt0s8mQ3pZ0P59qeukltFUxIroMehUH+ezQYQ5U0oN/t6s/TTp8uaGxWgQqM01uVo60j2CU9iw
MwwEP+1+gNkuoD3kJhJGJPsAEN9j2OGz0mC157zhpt0tMugkMUjj2pACoZVvc321PL7SdsnJ6uEv
hrN579zbTOFwDIDSj8DhnNLdWhKMq79LQh6GGlLHX0S5OF4gp02G2sEzxb7w2UNhoivg2IPa/K/V
2E9PUjFZV9HqHv5aCyZKBHQSmlIlH683vGfvDQWThZ8JGGvx5Ut8bR0uUII5to9IiJ7q85EmtqrJ
5ok4l65N9sAocOLGKFL0mFhdKL7gDWHbox3mQarZChpdBECz61GGNvEDv85Amzvy01ylbm+XETA3
VyuAziSh1dMBcG+x/6b8qGJX8gjdRqdUuv0zp1CFYOfmrkOpPT/JJi0Vmz5z0H5MZB+mDMwzxW7+
A6T3E4e9kx/x4iLIugWnuR9fYOM7zMzM4WUwgVchdEh73kMbOgZq0EdYq+juuiQz3vrQgMF8fDY0
MH+fumxnvt4OoUWTcRkpXM2kRrEC1qkePV5AiphffMcKAhQLkFGxED5LVQsd2/NugMVvNtmR+0zQ
x/O1TdWGBHkmb+7rShymSFsEJzg7Nj8WBN/Y8gqvOCAayLFmjGQ+duduZgHKgdZHejXmEN04iokC
3B6iAA341cEfKslHLItR/DBnSGDYtICCNJ1VNCmYQAycde1qLCf2pa94VPpVoi54IJ7u/NauEJL2
zxKZVCFyxHvfTYlxhGhVpIrgs3Do0ftKg8LdZC/Ecovlqt5rel8F4PxXEY/YNc6/TaqJb50X4KIt
7vpbldBIVLltLTUFjMg4Pmye1XfOJtY3ehRNr80N56bdygb4kZTyWBCmTa4qfQAVdk2+UUrkwDcf
W5eZDDoWF7zivnVcXNvrjBqhqIuEQWKFLkzgvHU6x9vmbQ53JXxldy0EvOuF65WmaNj8HwV35I9w
D98oHY8HReuXXG44HznkROj+qvhoo/Uai6afQJ06gLW5jK9g6ByYKoWd6hDH5maeTqdjzbFk/TId
sxGyj6fCcEu1sym7zHYI6302wTAlaYlo2tjOdKlnbJThZs/vN5Nlt9YaQICCdaMcUrdjw2dkpIZ6
fZrkjS6i5swQ8g3fEK+LT9IVdfvRaXI3zFbL1iIEaSF32Ypl+hh1To9e1QwPLM/BhhAirkIJPnSD
LGokuKxLOgGCWet73BOGhhq3CdGW9/FCPkuptMGLHJxjfAQjwLfwL1LRLzU4rQhWhPT4lB19zt6H
JQBmlQDs+sI+f8x3W9U0GV8XJeuDxpPsYoQXy/dfpXY0nWhN6mJtRg97ve7psw6YGXf7FZ38nG25
ODGQYhZ34v43MJyi/Fo28Qflz0vvvIpVKYs9Vq8C2c7Lr30rFYuYEdeJSQoPEbv/ntlUci4cGEps
1gpuGf+Nj30Yfpw99wEwF3qo4VhiESFNimnPzwE1XSS+C9+2JQA2QJw/ZaZ4zOowjOjqP5HufH6e
U5rbeNnMUsJZRPi8HgQfHY4hk9jWZsVd/O+pDkqgwFvvOFM8a7+WHnd4/AyQIqpFEPGKrb99Cj1a
+x0Iy5qaF1e592Nc4qaHOSk37983SDF/Zt4Wbpcv6xEa1Qxl4fRsQX8JsQ3HgEdOWFZlpfIbKYM5
MI8NVSw/4G7lY6BA2anmcIpCN+kCVLgOa6qs/avpjO1Uk4oS0vCtmzHBmGNODyfx/YsbKOzfrtXz
pxuoXH1YE/GBKHGupmEqa6KeuQIsVwKWQe14H1ibZdAM+j5GD1tjU+hyQzmwZuRy2HGfxzEE3JtN
AOTV9KZWdKQEe0VIkSCf63WTtm3EIQE5puqTvnK3wk+WvRphNSxxgPT8kJpgXoJhqNwMOCh9LDet
oRFzAAjG9Ohqr/PQ4/J+yu2AfO6tHu7sWpzeEhisRuzQYoqD9kExNDGQH6Rw160MPOlmh3cIOjNz
fVa5zq5whWsyiDgoNFYQ85HMLDJcn8OCSKYtL5lLQTv7cDNSFqd0Xx7Qjc/H/kL5Bc+NOZeB4xxT
co9xrx8R/6936/DSnsAl1Aq38b9p5rGmkrIdSDcUWJ1SDY020PO9Dg68NSccLBJF5XiGvlSSfeyc
Myhpo24QIz8OQYbFfkAecqzFvskgd/ekEYqsiP0ysNwi4SESgTmBMr5XBiLsG7LV4EHfjmY9EFr3
r5044OvtCz5RWShC6u7KG9cCZPWaMLyTnxVmhRoLdv2rDXUUa5hdNRMAjfzikbqEqm6ZUa6UG0So
RY27YizXiEylysWzTPOKx74O9RTBU1YFcWysvJVJXC6+bgN8DT3wqWwL9ZtmEIOPcWQh/YYR6Aqy
vAgRz6iL0qkrtLSyKcOj3UqwxT3c9Y9gclYTJ+mhC8/XyJX+ToeYYxFugKPZpPIPazm/v0pvpNqK
q6Zo19+dFIRrbZdDqOgg15pr2IbaLT6MaTWXPX5oZKCFJvLFYyuzZua3aVOmQmbzmRcn5PoPO0rc
c5f8NvEy/EGji/1zqkMZZd++ChbfeWel/AahyLGY+b6g2evhRTyXdCG30uxrkuMUE/O9vJF+Ze+B
KqrS5T5iv85j3MNyXOtFrqag98lgavwDRooZiosaQ5dJpmEOhCHjWFqHCrtb0S3VDoaf2H6I7UjW
jRxBOtg5zG6tq1ovsTCO5iO3YH2c3NDiBtnTgpdAMm/340XeyfmtzmaXtCP8jHhl5hZgKRKqfmzd
CHa24zEh+L03oZP06mBPIGY7dciD64gzVDtbdHUjcvMXohKzQYkCY5SjgOoxAhL4+bj/E36QlihM
7r7zgZksn1R3hmDKfp4u6+yWC+FHNFwNgP1phtD96fEVtpezH3IvCieOwlXKXA/TTOxNAc4b77BG
OlANtghr8qxvc14f38nKs6/1KstOn+yM7tjYTyLBlZC3111UCyt8I9dYv1S0Fru+724/oigKKiOe
HUy7V9CUe7nxHrsRD/xD8ce4TAzoTIiOw4QALTUcbZ2x03H2JQG9c1x7kASbc2KEeyJFpwWRO6xa
KEd7HKSG+bJhzd13NF6Xbl/BuI61QFs8lAoU8wvRIe8QYyi1KU2M2Osjmb/kp6w5Mwp+Z26qp4n1
wIQXmRyGhxgusAGsSh9AxYxeV33EoUyr/hXRPG5OAcoBOvXeVZPD+sYXO+KKWT4Irg0sJIhLLI6l
5N5S31apETq0/fKf7ogAVBsRotTSrlTwThChDHCxv2E1X3boxjoa56WcwJtEk9SDQmI/ti3tv+JB
NJGaw51Gi+Bx5I6C3mEKBjXXqVpFVEfyK+XeLRJ1mo5kO6CnOenTdMTIYF3M73Ntt1nsjipU4bxr
ZRe/6HJl1j+u+0W+JGBwym+qyFOQvLyJjW2M/AxqSDX8MsosZuhTxIKnPVXTGkRd6ZsLwaPmEufz
93aOrjN7Cju4gaRYSBf89nqxkEb0SQJsdzetFJdPrVKvIHRazKr5aOKbTZ5XubJKp5uNZ+SPXGrH
fRiuVyiary6rwaWs4pCLDvrz9KYdcd+5PpxD86jyoebP93ppXo24tsz2XqobLRnXgXA6Y3GmTA7/
mKchIvJ43fImi4Fj3iUTBLOyWFnyt/dnd/Bp7DoJlB7jLlvENaIKwj+kWsSh8JgPN5sKRoytPOw8
zJsG1SLkj9jyQs+qaaiY14hjda17Uns5BmoSX/eCTPZP+zPUxzDa8bWiU1WUIW7z2cPnhpxkedse
mnOLz5TJkjDc87uvIIQK2Uc44U/lCuQObtHogSzVobqC1GaUo+PwVeVby+tW4LnnhpAJpc+fdM0l
4rf6DA6FhzABXwsXBiyQJbkn2NtzkU06qJ2pnS+9bp4Hc28JBPQFhZdp5mIRTeVVtkL6FMNdPRi4
kYQ+LM1tqccbapzzl1qqk/iKOLzFiIz3k3Ou4g4dJSCln4+WYF9jOrO7tWfNjpELYV5pbq8J0KmD
pl+THgR7S0rH93pxSGfCWRGE2Y2pkICko2d8R/BuS8GnNQ8u0270M96gSADTUxaxG1XkL5JRzEqz
wJ5sYHazd7+lGR9VEVukNxczedgxxJBx0pmJxQSuTUoD1fRGXRPIWxZq2WgfRT9L2c3IIqr9nDPx
VA21Amd/I/ysHidTuGhGUrK9rCYx662TDa6k8XhJ9JY8ldhDCGZPit4BBY6FIhjjw+7yLSX02AcK
jW6oXE3aWWSVdWpmBmvWAoNfCUimam7XQd5lMoQdyh41xkQf9BQye/gFMOFuP8c6Ph1v99BvfQ3R
Rsjz1OauG3fZE6F14ScTfljlMAbON2l2jQhNOeSi0SdJS0Scz9umLPQqz9HK7d+NitP/CUDMrIAx
13VdhGUeVro01iH0noN5i4MfBeGCDdwlbE40G7U3mtIdsDUw6wjvkFcSU5aHQHaELk3UDkhfswkh
nYOYR7HdFAppda2vEjvoXEA2hLgrOc1Jcyw6vgjY1gGd93wM+0J8SD1ZCj0b8HPEZUW/FRt/q6Rc
meDp6UD44De0tO/mdFg6hj3NIm/bOHN2+R54OHlxQhoS2Fi8i0r5SAbWW8sApQWHLLMKOMKFKy0P
hXptGeC3wF33Lz+cVfk5KXeuTz6FLzu1SVGz+wbMarqPjb4CoPNoS05VWhQk+1yw66Cn5CL3wiZ3
Qaoo+pZZuUwwOVPdc8/ErETW/E0cWxjwWCbahcUuVL5+noxkGnYZiXnyqpJuJJYd8uVxwAUtYDQ1
SgIPSw8/2jpwkOf1EqGO0zF0XaWc8eJDm1XeoRO5F8aETeJxy+356xRaSOpSF5pfg4W5Q9lb+fNk
OeLgUtoLcmKXODhReWA1byG2Q0CvaqkeNx7au5Pm2SNBAeHtWH8O/T1IcAMmsB479EntGT8pA/9V
r+N3ZnwH/ZMqqMxbI+xicsgVL+OHnYcXr8XfCIJtUapIZDjndMTBYfAkneYqWF6TmeRVNPC5Uno1
6/vfxr93bX8yUHE9RFGMTZJLJR/vnFKrDj0wmmG+IsEQ7R6okJG1zjQusOKCpFVITSu9fYVFQ+p2
HOGCl65iT9gyMPIqlGv9L6Gv6XzL0z4OYn2vCSiL9GgE1OcThHB8OsZkTIfW41r15Vm2OKmy/iQs
lQHBKsHT6C7LkcEN4PRwZhY/9ytm8rWwwMIlQ4LZN0lj6ugJikQhe59028mX6zgXNraxE+cGZP/v
nDLIqktqAoXiwOJtteFHvyEH4xS9zOqAfPrIMYwXzrZ/9/oo/94kf8sFRHazmz1piNZBo5BF8SKs
lcz748sYivs0IeW5x14Xpyrmq4RRYbDzRul4YC4OT6B8GZMUit5hf+fD4jjI9lyHQW4LcMSV82gY
09vPV3pQIByS0YShEY/Ke9YThopLwmsLHxrI67mZ+FIl61yDX1NPDJ/1g2AqZ4DKRwRHRveP5KsN
jUnHBXpVJjoZ3Bs3an4BTYP1PtgMDlTIzYaSC8zllS28zjM8W7QcTHynoHa+vKUOKUaZAAUfyujW
nzm4XwpYwxef5idWiBva2AMXGdIb0SlpGIKpQB8tQfgLRvfSXy2ER5QApC0YDHDuY5icQ/k+xhwr
MXZILPKtJVShQPA5MiS0X3AZIYNsJv0MXpt/6NRPmzxwD0tTXL3w0OTIFMVXC8Uj4dq3zK6o//Vr
NPLXW5It8GjwDi9FL9qx4Tj9Cpz6Wr1DvslLw/pB/aL3ASreWTSQl5Wlu+T0LVJcDQEfEMeJ2Cs7
R7OcUbgs+lLXX/jKTDOz0TtYiJ5OPVtzI0kMq9UDB0NLDUIBvLlFSCGBRB8DdUeQPARRBhMjWsgv
rPK7t67PhW2On4wxHH+DE0AoypSDi0EgH4sjJppV0j6j8kB2k4Eizv/gLkajqGjFolt3fLuYT/Ox
ejZUtFJXrhPe/Np5UN/aqui0aCqZdlmUOn9aCV1jksPbEjbOvjDrHwtVCgEkxkTEH1U5NV+13Mxm
hnB4FE4WhRHtHXiq+Ts4GXTCYKSDpJWOGUGssv1ITcRgblF9QVDQy7Bw7RxwjgFb8G/w1aC2D5XK
VYOdXb/NwNPBcQMzOEjwX7cxUdZfrXLnxB9EVfu13VW4yslYy6fFziUWKYD5pVYjn9sRrdA/+nb/
LyU/AiMh0e/qJ8elcvVtd+vrFXqgGAO05IfD8Obh6YaNO3xjl/Viv+f3EuCB86ApqF7vMc/PEwOF
QjEDFaiUxrSsE/EEbpw9mqSYhztsLuP+JccSZ2yCPR+XEd8+bvnqnAh93/6148IHhlJP4SUgfw3p
+Da0IBZenrr/ZXyaj11+fs//w1j7LI0zIqnlMsy8vkUc+OBw7xSBTitRjbotAjJLkkp5z3rm0LH1
reY19OdD0kDRM8eCxF9jc2ZeBUSo0nY1LAqlyJRUg1F/+lUHzD7dpsWU/HWrbjuEbSyGuTYjCVbR
VZXGn0RuGgTCL0zOZYjCzWnKQ4xokLBkuo5BkCnwGaXMOp6xsM2CvLwt1ioPPE1FgNc514BUWRQb
SkHIzv+iu9Zbhby0yxlzq7Ogv1UmjKVy1OijLnfmpklZv5xeEMxEInE8xCcEtPUwHZjzj7+0t8l4
bIMtJDH0XBiCJArc5Lo2vEupOl0WC30ZIt+Hq4gNLPLjOBkWNf9nWAGVgDPX9wtYaehRfo8Fp5HH
IRZHsMKbA4BHgToSUFjSr69acdX++XoIRsJlM05VyXx0igKO/gxvuLwVIMTS1Ai4KAt/nfwHDa1R
RSJWBCKN8A6U+iWzEl2ypFalbXHxPnnqxqgJVZTJlHY795Gj5QgMek6jtH0cE2TWwu8y0L3umLCD
jQ8cfdpLzVbAZ3mWV4JiIdAqz+lyq8wAh0EoFNzfDJV2G0G76G6iOO6rBJGigZI8ryGMUHN3eK2N
OaEf4vz9SRHr0Mufwgu5DJPZNLqM92Iasy0Wf1rSBFtxOk5LOnOBnI2+OLxRq4JvPJKsibR4CDU4
33i/IoLkqc5l9Vba2dAgh0moZOqR7KQR4/oJNLbV5ZmmN4BYTvyOU2CU251WPW2fqX6Py+Os+TnE
tZufndOpqKgoia5eTrNEpii7EgIrc7sSCAv7vaH06sulF+0ocAVwBAeHkV/ceHhL6AdMKnjcSOr0
dWwmaP07qwrayZqf1JQxvZM/QXEqHLBCPoLX4+pi8FHzkdUKALDuhR3v2/r0QJmqA8FcTL9xLWK0
LkzOB708MJFTK7pyXLxCQndzC8F3/6pcW2722orOwLmV7/Dc3O5OQ23L7PwBn265lDOpWc1J3Iez
0K/sK6gNLqmPjdZEp4aDLqF4o11R8MyeuZBXylmjrwtyDHN53QS4iw40//po6bCC+4/0zZAgPqfx
AMmUHfyLP7NGjtgaSXq5VO3mxvbVeU+/eTkQvvn0nJdtCeDpsGC58kYTRxkp3OTKdXSsSa8IPkK+
gDg6su9hCrvyWJgUsERWMaCz6u36hAiYaayUJnoSUWIN7IwK+Mcm56ODzxFtzspRwryND4xJ39aW
1uHBqC7Ac9cmPvuhbqkQyDqcn/MQJ/rgiqtRvXRYekKUMX+bATxTPNU/uCyoDuTiTj7Fi3jGF2Ri
8alYUdpLeFjQbzFQBeunPP/NjZxSbl73l3JsCJCGPDbK44a/V/Xnbk6bt+Af+9cZyg4L3OebG3l/
fiII1ssJTf4igbpvMmzO4F2IHuaNzg5C7ig1V8Bx/dsA9KKxzxY8iZt5f5DGafFsses1GtOSbhIL
DUERQUEH2pXP9mmep3/zR62oNHT20+X/bNre0FEA8dHvcurf3XNSaQZrr+qC9qT96/bnc+Ed3Npr
TZzZ8qWYqgXz4fvu/1y5Lgyn8aBFnpSzvsBoZnAhcbj+wMZDwGvoYaj41dXLwebx3y7RDo/Qk4XV
R/vTjJIz+EHAc6+oxP72gc0WUgl37TW4MW3Ziiq6S5Y7h0cB5JGSJtrqfQPfGyMLfT1qhnuve71W
IfChSn68Z9OMUI1dgH7orjRsfzmIeArIzjgp/qbTAgfHbTnClsK6YD9SGfULaAF25igzjIbI8hoM
uN+41+xFIYbSf3RjB2/fOGKPAprNpujgj03+KoYD7SvHxvnzf6lZGFdzVxcePYGFoEgWWg74nzUw
af89cmLviLEi5IKlW/1qflxaBRXPzkuslUfDxyCfAAeGVTLdeeHqg0QgptUz+sOQK2mfCny18Kii
ROWn0LVqwdS/L9QspM/vwHHXI0lreG9BQL1lgCxwehUMBPIc6zpEYL2G0Q7oEp8mHUVeOO8o5IPo
3RLWjJzcCpR4GvzQWHRdq4QO7h0Nn6XjX1etzccj3QdfxLhmn+J5NC0dqW+0agEsiwlD3d/vj7rK
RRS0wYYj43IZaLMFiULaxdxgwaTejCiyIFsrKqdltCY/EaupsFNeLlEGgX88HF6h/uow/CMMTSif
0SX9Pexo9XtcbutyHt9o2h4LugZt+s/7ZsH3LYYcWHWgbQwUDp2FUEGHOz/r3EU7nvT1SYjnUap8
XRqJfsT8KF2cmNHuIMJAhRkiuhsWVXdCxFmpZKlF7/totioyL400zcHhs9xIVwrF+pRfeMnh0704
MI2TMNuh4Kap/ncC3w817xCwovTmPaQ6zgWX0pzuWjwgUXwJBIxUoaPaG+GYJqF3C25FPbVq/iBb
YfSZoawzIyacWmnA4/j6czMvr7CQ8CW7FkZZV8u8NcqjsywnGAKPDxXIH9+LcOTdbmzvqJfm3LiN
TwC8EtsKRRmbqW7qtq4Mhnlgb671hoBvSsrjuJnOtY8Ogwkui7p+rNoeI390YZWzj4BGQG/oDidW
zjLLJQPeHqHvvRYj7RDqNNv2GG/5FLO0XbNPaupzHh2EtjUW4xkpWITFcwx65ni0xEp046nnSwHX
csh4fgmOv3e1QduEOd+HZSIJjG4IUoZNauj7Cece3J2JIjp2BQx/pz//9dNqxZbXQ9zZUx88QWSC
af5yK0+pGB+t8Xrm1CADnXW7uqjfBx3cbifxUySipV7Lbo1RNJEiZOU5vp3VQzEnh73WMl42xzCp
72+cg7OSYeAb1kHowZ1iScAuHbzFpvuwdb6DMssG6gforwpdPin1qJ9jQE0hPxwzN50nzxJLBAck
N6f3Mu7IXYl1/gfKkwmL0G7rb17Z3TgHzO4aS3n2LDdqBjEdyJRUuvJF6WhnKbxnlTseT/rEJziU
d67LTku6o0PBYIvtT5SrIwd0H8Oou02By7y6EnEmZgBVaqGWaVXJsBNfUFgUSNBR+NpRoVhZ5uq3
UQgizCcpV3bRrt9qLAqXM3SKJeV7nbEsPciBzAtFs3N3tePlZUGmxWjRos94AqPtU+Hcx/wHTR4H
Rol3568/5iRGsIwQkDyVMVulWVVZxWDJNy/jZQdip0DIZJmAOSuilqMJIdXKpCYPGTH4tmapWmii
qLWWtqZdIpPYr/ScFvS2MdtFSuJRiehsS2eWgMTw6auBCHjcYhGOvw+zLDXTnMRGwRue7kgEsrHd
I5sRTQ85NBpFJn/F75FB6WgbR+3ndwyljhpElbtoaYp9NSy57vGRcMh0jCpJxVdrZfVVHFG0qW5W
zioftF45+X/p2ZRC589yWbz8ii+NR4A4R4nlmbgcynVptR6KRIxt1Yliaj/HcNWMt6EKU1YAsnlq
TjWsINe1k9WVyJN/bIVO2cPYJfKsmpS9sX3+By91p0GiRJsj9iqU5gsuMJmMh2hJm69Pi08bJ6Mo
Q/MMJp6ymobRSb4G6r+SMqu2gB8/esU7Iw2EJj4ya7iNcwFxHyg7hcOQ5oMqJqWx+LxTX+Mn/GBm
+1JgOVWCaNcoGARq37hI4EYrwcHFZ7NVTJqQ8ZkmSV31EMSLJvMTLLDFbJBDuBGl6i3EtylJ/N7Q
ZAUBO1Hh4FKPs9O+onsWBgocWlOdAPCKKKVAjbsc6k4mBYsQ7V6kEds+nuXrmlQg7FjEkanHVwFu
/HENx9qBC4GYcIA7v1Z/O6Y+X9npulJXTKZLpjq+oyU1qC+3ZfXDQyPTmj+jnkezr+ZMmpszEuOn
fcvhBcoRM7qGvaZ+YsKNb9IDV7t9R6w6f+1KFzM0ZO0C/prvPeiHI/ukKKitZ+xV6gJH0jbeZLfF
xpNH8lfUqOV1l0BC/IHp5uA0Ptv+jBPe66lreV/MSQwnArW5Kvodyw77j6nH12UnarusPhF6VNYL
wWs6OvEyBUtKd15JPuU1vm0zQ05q2VU/m6S9n60qBmDqcAotWo2+gFWxh0qnkQqgryPnehNuAyfc
yqBM3U38N3OXanUh+fPgI7wepb2vK2fc2BcM0jVc77XsIc1XIx0lNb2Er5OhoOJ9RhO584GPX2rY
Dhcw7R6EnASgLdxs/fVi0WeVcCCcx3wezjsgWreWewmoT/RCCXGSd0ukIWkGHpMJJfuXZwPOkBxT
llsvCKr2sLjPMb2uJm7Q2nqQgWrVHfCSx0W0r2t/WXFTJZm7Np7NRzfxMlsyUyRa2883u6pTZONX
MK0ijgCHCtn6LzSiSvGj5UG225dGke70y04pCZ1DHLISf7vAO2b9FXzJUedMLZCSFO/gyPdazcgw
MZ9c7ewJvTZXKFk+/lK56tmM5diRu0fvjlltFqldyMkQeXzKR2YwxqXB9pAKAR8TY2HWBGgx+lSS
uZcpM2sj2Sfbjuwk2Wq2hwR9xDvQnzxQOjaL9BxYzucPpnK3whTGPwUImUigiwDIWYFk20ebD3ex
S//riKgOQw1Oizbu5vOXIJLqkT28p72Kvms4DdYes5ch0SyXDKWcqTe/l8qntx4YVk21uSrpnW9z
bSaJmWsqRQyEVTkzD+btWsuoevMgfU8LezYP4xFn6nAoQBMeNg/xyPmKwmeoAl5RtZh35RrGDkdF
nR9SNkH8u1Ml1mL+rkUIPmguTcGIp7JKceQDi4KHp4TE3UnXnZblmIUJ4ScMqZU6B8I3f7gIULyF
zm19x2RL5EViBwt8atO5LEioZCEvycpUdevtdPHay/zQ31kNSBkGb4hgi3JVkvd4wVc/f0z7cdQN
JETn6KnD9m+usCU9pqSBFJwdR8WltFimtJ1Cv7KbuCV//UqjUPesPs+fH5nbge2yz3U2RsabGkjs
n1in9CithFXuDyG7xv/OuGre/XzKGq8IRkgsD3vIJP/NPjHmYEItZnvbBIfmyWfB/wKvMdhqA1BX
C0gLGMIag9YAMdkhGGGD9STv7/7sMpaOz+K+PWXQ4oS8/21G7907EVR2bnqjrEbbAoHSFs7TNezA
wKV3bcGB9XzMx4uArhnje7rlZncKl6aA5QWR2r9hOuXSiZGZ1ijwn3NlVitge4hlxGTPgBTN8XiK
1lSaZoSa1HivN3vqwlL3FueOevErVjAb9XKwMVLnZAn12K7yLVGUbW48X3xE1yvp26/Yl/i2VcFt
klFkmpBVg+qgFUBD2g1R4IQzqLvioOcAo1vK0qp2du+AYQAQv7P2ykad3ofeoGJzEYtFegDTFb4i
kuydli0RpEGLNq6QEB9vJQvGsM87lVGeP2UI+QHm0AgRK9mQtUs7gYZMb8S2wEe5W88j4qQZvV8l
ZkKu+Cn4xtvKhuihlDqyDXBvYPndno4HI/gyvMgZ3SqrTXEUW0MI5FBRCI+Y4SJ6av1tQ8UYGXkb
lSY+rqPLcoyNnqiTQR1tzvYmalaFfXI2pHqzRaNcSIoouyG3bhJ8Hx4scx1zp5rpxqD56zYBJAqY
5/zg4FwE+tz/zGlxF86uuLVMk6+DLr6JTO+9djXq5HEfkDLSK9+4gPAhuNGHg4VxB0wU/ZeiPPtp
cw848VJw5jSZ8NgkaLlvWyPx/AKrSEHPAHDX4MCYnTyrWXQH9BkA77tz2Y8s1ZEqJ0bq38PFvgKJ
ZQ2yUI7OzE020NQOzvnKEaZDem+TgGKING6nBfE66wGlB0+14xBEQidTY4SNKnd6t3yCtGn1MlZr
cVCOtsk1ZZPeSmoPzXDDRWw0HbVcBQO6p/tBaJAGg5GQzgD5rdTLWdLQcjDYkD2luus/sv1bPE9P
mPQmdulRENnko17TWdHxAB9H9IBVZwhvZJ7JJT82Wqgr7XgH3GiLKA7G8ookL19H9Jo/ISdQYeZt
I4QK1XraHrdrcx2GjWTh1SX9RMOc1Rb27sTyHZZ/BsGkaVl14+HECqkvwfqMebJE96sWYKzFoMko
4dCCEGME5kfk4UW3A6jjlM6mhOk7L6krphUMjGpcbpoVL1I/+TeSXneLAlfsrA4Y0NEs85b9FHrZ
SHaX/RkzSLnJMYRM9OrwGPQEEf/RIxj45XzNaa00Wl9DmS9g5ZG47zzIaSyF8TuX/Px8y6Sftt/p
ERUQXeMc5YiomsHF/RJJej8MuCu76Uyl/xEaTlV3Li4P+2RDa7Kd6bikzI/q/KlhA0X0a80wmz6S
HnYTrJ3I0xkzyrAd2OyFso6x8YuJfWMSZ0KL2MKT5NFjUdVV2zpI6+WrT+9UMsSD2XK9sEoKzFYg
wkZOYpwRf1bgtmSqfwtAU/GzSXaod8GrGC4bAobFMSHKa2t62NtqoPRS4DxBNZiin/iLRxFNvKo8
H3CUUS9TLd25YidmV3VgUGJabi8CHM1T0tFlr7wYHnhQb+/AT5Ki9SvOhzdAgQyxS9IuuLXdi9yU
2L7sClIbCTivOG7UmJ71Q4w0qxuIVg9KpCjOvUknarZao6Nd5in0SN/D6VnaKlJ2mSi1TV7Zbgju
doSlsmpUpJe1pnkewc10onbcDF6z41v1olevKHMSarmxDmDlHhwKKL9vQRzMZa0HSkcuThyj1NXY
b8dLyvhT69Xo+htNU9rDa/4l6w0FafnycCqEniLq8LFPPsnLqd8mujqVhpQDoEYn1/DOcwpb66ek
4SCFuM88aT5cye59l0eAAVqfkF+tH9FToeXeDhYrTvzA21W7JQyp+FoWEaxiqCdOfskfjB2zLyOs
+XeEeZ+0XKl0y+aV1XPU8JVnHRMhM1jEcI01I0j7BhQSfKaH0fgZk0yWGTQf++eDStEBY6of6JO7
wmG7DVN3Tppqz4W6kUyHvy0T8aqZc/A80zcOWnNCo03Pz2xtSO8GfnringAnZQsakLcjeg8A+cRL
DxTiGrXDctsX9l/HZlZyc1KnsfvLeX4wqG2dDMapEG+uP8wX07HrPizW1LqVSidI40oK8s7734Zm
lyQhMc9A3VWnLzH5Jw5uuWufld1MbjZ1JGIZSO+dJd70f3Ny61VGs7DoQV0mjOMAfrwvz9T91637
MtS3amAdlPC1IsaLTaSjzl1tJbDG/ZNxGPglewamOM0yUDphtJwvJGd0WIcZBQDRnnW5iDSXi3bI
Jf6XSRFcka5MLc3hUdFR36OQW7wbCyZFCMv2ZE+8LsWcedsO1IRz3KLbJpKEIhqjnvrg0yIEG/Ow
ebuRqnuI/osJCyGSC3Tu7v1B/YC5l2xym7jllW39aVn0lBCJdqE9CeKde4CNym3v+qRp2mJZ59UP
epEt5pP6pesRST2yVEtd7QwS0XMKxYl8Xhxjrl58mlXJZ9WOdrtncOEdAMrADm8kGICcEBrMbRlD
aAlF5acaWOt4eKDJHOqKGIbYeR+RF3DW3xMYbnHju+3NXNZHBOanP6sRQuGUtX/3aBHm5P0pB1ff
COFJWuUYv6+vcFm1nCzDVjtrG1esB0l8JeIQpHxyyhLVN2C0H2Of8hrnqn8LcmAzNnqY1iYunWnQ
FczwWbirZaMmXOgKZTN3FTYTB1s/ppZfKVN8fr4BxWTghTAM5D2CUH0T88yV7IdqHiHfHUTWDP11
nrXsrGmZ+B1XFR88jIvlNjFefk26ZacMUuD2WlV3XwfBhemCqc3WHQkUTxwm1vShXY6btifYPCpB
HbY+wckbZDAu7pAFqNXuT5k4sRxL9S17AuBdnWx0cJPU8a+RdYsqmIpOvcIrkLM9218pSCQn9akS
Zax1pQwh+G3kluzQFZFI4CPWL+5LgR6um1+/shQHUwsIMsf/2lj8HasnZ5u4AOTD4rpj0tsGDzuK
VPkKdsg5th7W1TJaxIK/vP9yFSISDF6+gjCXzo5Mb2P5oa2yTNm0V+m1KDWix1KwWjMLUUMpP9is
TOIaSh9JYByb4uqWbUaVEtMIUm9olobeDpZ/7JMvEjlnKNh5lsx+yireEJHdpOAt3ws8/AKjefL+
35kbzexWd5JTl1jX77HvhcXDc/Ko1cGICWMi8/lgfHq9t0o3btSBpGk0pxU7YkeVi64vLoX7Zds6
QIquZq9NeNAHbH6De56ERh8MFACE1/3LEQPEyrVEQ0+vxCCCGsbHm3ZOWi9wwzjNkHO9Lbz5BWZi
hcD1XIUZ3J7fWue9E3hSL6DSqQHb2X69Ud+lxxlvNI29V+IE1YqlMfEMKpK3lT0/X2S8sbLYLKrE
QSgbLUKF6plHRsavXMVSH82wnXVkZ7VEoLIi/hwwmSyMrti5XMy5q2unDOopNYu8XFRU37NyDGgH
vS5+ivnthsgE+HxndGoPzDIuD5s5P+MIpo1cS6lm5nQL6mx7MoBRFsOPbUxLlxaBpu0i6LoK7IBI
yKcB4lOdwQE+3Ovq1UHtq0zKWzb9N9gJ2qEZEKADc8iMvFqanMR+9F5C+v1qt89UxAgTA8AnZGba
bhwVYgzyCQItTzjQfwiCUn2sGVJ/p5I2Axd4HK0MFCNlH3ohxzd/z0Wu3e6qwBdAL9nbbr55OjkN
VNJtHT/juL8C+yTkms1ovrhs4cenq+wkyhehNocYHFT1cnm0kbGQ3aQyA7wukJl3RaT1HI5UCxxR
d/CKVJEI9KJZCW5lvDCypojbBJtniQ9yoiTZ6Gvoxgw1n768W7CPK5As1tKYgsp8yDfjkBhkAtyr
T2k0M4Ezwa/ixdia9GIWRwuGFxsSzPBrITjCr6Lk4tTsymv5nIh4qqfG6otMXvXXc+RNY53FI0g4
SVomXbXt4SmEVI8PDfefpoiLUpS+/xhvMV3JUaxjBvUmvV5zZc3JHuoHn0eZVHpOpmgos9vf6tVd
zIdA7aoNnRlLPR14mDjB2A1n/0pMmySlzybLUNH/TojmVYLLKTwqt8L10Qnir4V2V6InC9mMlU5N
aJYS26b/Lja2MCH/1W1CUidsDEzeSpqJOxXLTJTyaDDH+AhNrmlkCpsn8y5XOmPv/xDueSkf68+p
qbTmfHPJ5z1oxPNDgFjkdQGm9+dUevD4n1V6kdGKibhc0xRCi+X2yHTx32IpCooQMjTyP4v48aKf
Xsk0tsYhnydI7kEjvH+c+vR15Uh5rxSMPP0lX8jS31dkbSYOo661FQ7Rekw2G88f4DKxEZUAVfRL
rsFY92ebo6u9yhqHK8ilM+5mu7BeAgsW8dJ/I+6BoVyKSBLkWxj4Czrauz1R9ALalSW6dg9I8+uY
MSFgAqB5ArpIBbGWJAkfTU5Xa8E9AKjJuAMnBsURcV06szAX0XguFMoSDl0LST3ZQtNae6y63Tq/
kvbjKNcFu+Ko2TmL3BGhAd0KZSymURMWa6mbZ5jHx0bD/PEORGw9FQcwoYKkMmuh2c1ZwiFdVrxj
44RMuGMyL/B7zS3BfJ6BUAkprWR4KTFzW520gsInUI7kclFrhStBP+RlD1Gxv8VcZmIywGpSmsog
BkpVr7r3DB+7tNcG9witC3V8Px4ueeH31tiEarh2aacXgPhhXqw42l8GHnhVBcUEy466DOXmOp17
gXC4oWvK0YiD9rSwomSKWATzX3hobsrvhdeTn588ofdFIZDATEwLolCj1x53xWf9SlWNt0wDMpAK
u3I8mVMfyLgnSGiZGiQOhRYLPW4309SdFi8uxh2KKMWuY7QpKGMjLbrTdycLoEzoyyVBDFU4XV4J
qjsusENGgbvpCQq+Atqvgf9QUN1IQScQRJmwjFNUfjZyy7pdrtuwv0L/F+Yyatcl2wYCFJBJSz41
PHc77fiLQsoql92fEcAHp/Ei2ErjqCK8N92S8g+9KP0m7UThq7UGGfeTVtYvlRCRrVUFkFRx0I2S
QMABJ5La8Qg3cGEva48IMp18V/bOVoVHJxiC9wAhZOl+Efn11Zja6aLy3jfaxfWZWlNk7Sl6KpOU
hzqkfVND1jzUWNJse50kleFI0dYsJxG8rOhvIO40scyrGTMVf0iiay/hl+jlaasiWjIjjWvVBbJJ
0FBiyKQcrIuA7AkwA4JYKygSTmArY/aJOe/NUhNMpYC6gz3hiB+sI4XRvxHBFet6q792sDPIimJI
92NFcmTU8xJJZx9S5l/5Jvqs6m9WvAkz0fZ6xghFQMOy8y4fIRLYcRE81wHT5gGApph2vDplrBo3
3C2dgz2tvHMPBAE4UfQ+WenwPuOpArbJ6UzJkMpwP33tlEooMlDJVtCNdUQ8Mv2B9uAtZsSKQDL6
jwN7pI867vn1aB+AdxaKdTb9LStNm1rrV3ApwkmImVshON5QhuPvDbl+fws6IalwUxD/8Kl/v/se
og5xy8UW1+j/tPxnbPSmlTaOQpzGBIPclR0h/UO8er8rA0oGBNIiqHG5vfUIOf1s1dqIfRO0mkJZ
vl1vK7VkmjUnUsjEgNxlAhzlQXT/NQviIPXIJ4FdAJ8xRmWu/0M5/4kw8zWRb1tSYmCoqX0Oxwq3
R8GA1oPdiBtUY5dajWKQG2lIgi6ARDBeJDzbdc1Uenw8rOqLJQekHfbDRaVO6SvpyrPVFuuZB7Y4
LiqyY30S1wwQFaXjKdIDyxNwhawICF2LJGQLdyFvMm7bg0aL9SfPQqPxDpRojYHJ9m7MYkfQO3HY
EI+fVabJz6Qo5z8sYGMxM+y7P9T+3shEJbOaZO6voa+mVQt87cPzGt/z7z3EqGL6ZUikoRrN43yY
tMeYExdDRYPpt+8OOa3WO1OKvvrrLSYddLD1VEzvO72x72XR09Ml+bRCuZyzoKfrDkKzrCZPPDPn
qzD2gA5b7DxuL9mEMomW5r4XCNPUsHLyroHQ6JE/2WC71aAckS0Db9yavYgORISrv0Fy9iJH4BkN
mEdBwZ0mUJdAmzHnBPrmLDypt5i7IN+FJum3ukMutHKubnl0/9GHU9EmCuynYFoxNwFTDsZ5vL05
ezbyW2nlDFQ+iTf8PVMAukFvc7zG3NLxKnplkqd7gMdTk7fSwKYxvH4bq5iQ4uddZaB/ZHsgv/jV
w9jx02TWM/cPJutrs+IsfgW3cDIDZTkXvGFnxjgw59UVw6Gp2+6uxNyL29ja8ESwCpkcChiCpzKm
BKlTVJypB9TQIvJoHBkQU/LpyHuJ9llH8ai1pdOk5wx0SYYxHFQxcskfPATgWFWMLy9sn2wtav+J
O1LnxevX82KLrO2tCmklL+eJyizAJyetrSyckZjHUku2LKSpbTP98Ed/KuduhuLdOtpo+fRXeWZG
NXEFZjzG/TyEnjxguTPiH+eHJ3C0mijTHNT+dto28o1j56iCf2kOwj4C+WK35UAUtsbMF7ybTkio
FB3bto9Oj0bMHml7HE9GPazQIqiSGPtBKCxN8z8gJcdQqSAdGbwFYOOIIPuISf5Rp/NA5BMJE06d
CiPLfYkCkvxlNWxHxMIwxAB3cHzbs27CKgzldDuaegpOUunx7TkaYPt+kGIy79lfeqtB+oeJ0LV4
owB9kJ4MmxBBwM51a98amDJjVBaz9VyNhkmZr/um8wdkhyCPi/Ra8zQ9g9deAzbh/4ge+4Fqfo1z
DyzaWydxktw3rGympMvvgozY4iiT3PFX+OaDuh8sHBaXQaV+SWh589jJ9gU9QBNI2WLYil2eopzf
ieKozw3Mt8kpf96a8/C8cJhe+1mqvXwg0fT/cjHFLwW9dnITeKCU8ug600n34XG8HO7YxD2xg0JF
SycBuo5YMz4L8wg55y52Z2CQ1Ow6Asl6saSYAayS89lZJiyEFuMKMNirg3sjmgdfxQ07CkpjJh7B
AVV8G5euCvGCkp9elU+hCq8CfspjNZbOMvpe1zTUYV50TMmFcvJu7mdR5ujI9x3OV70Yz7Qf0kih
deb9+ukUQDWkL4PPiHTM8yFW0CJSbSuWuA9cPz4abGZaiDsIDHj4jZT7OPg8LHfV3bhOAPkjCPaY
2OJMhqLrheSyAEhbX8mnDAFsP7wHsDQ+i5QbK1K2pAzCEQVO2uYSmbV79ijPVjxZ5AqcUB4dNsC4
G9bxxaZtglNaUQFDAliGCTqeVjLadGBcHWqnKM9TH38WFqVcoqkGLWpvk51p6l9iG+glBCV9Itpt
Z+YVWNnoVpRzCltgFEEyeFIX0zmHo+pVRLggsuPF3tkYLer9t0wgYiAty6Dr4EAj0EXY0J+OaWH9
5kfc3atORMJp50TdB+4YLxt+HRnyylFld/n+1F9tGk6uk2H+14mZkljaip4xrvZCLkVA0fOx/RcB
QD+GaInBc7+zTABDM/OzEw4Y29oaVQUdFztQDN1KI/wiNKuldvtM4fyBl28squlhDcZQLW/Kkd8O
iV3zm5pzwHb8EBgDX619jA8IoM7UM2qyEZL78O/ED38jijhJa/htM4J7GvOePGGvRZPRcKIE14gb
B5EGjp5KGfXtKUJ6DI3Qj/6WZosfcnqBsxgzPqhwaysElWz7TBrOXl5klrG/uzHLD86+Fcslxqtf
fxV0VQsSPhYyE9C5m6X8RUMIfeUC0gsUBMrvYJyWDV8NZgxEc3HTf7MikP1Rl/h733ErrHoRNBmK
2s7L2uwPcUi3c5k2TuBEGzPPLElD3r4knX9o1W0KXf4BemZFe8GQvjtQTnib4hTJt6V2FwLztDdP
/l0ALvj5tOIkyxoV8l0a1o0oLICmImpQT8m2cVIc0yO39esHHP3QLWVq4nRKv7G5KLay2Wi/visI
uLFIT2xRs88pgM1QPCuuD0/TPyI4QFVqU77qiaqJj84ulNM+1NtICxS/YVrHsT44R0bL/kdV8YQN
9OIVQa3tOThgknsEhed2Axyx0WfvJ6JVPifk8i1mV2Afbc6ROMF1IYYJiTxkoo+lJwOSMJky5d7A
zon+xFCT3UzDKwSanFFzL2kZ+w2rkNh5aW64AOyxU9cw2LuCnUyXeumymzrW/wu/24hrKDBMkutU
2WJXPpHjs5zjTnZnDh+fTOTbhiN2L+IrvJu/8mAK4LEmJoupSfrmhywNj/YbpLNQ1wjtxU39Gsu7
64skjc9lDa2zriMkbFZbC3zKM6o7dh9xzMkayBw+iNLoIPEOvZTdNd1dUYwZq3KgZC6eld1XEBsq
3CZ8HqM2tyikkwD51YY/G9jMx1UE66TnJovvOYRpPc0wCMmrcX42ULFa4kkwC7/ttiT+VxN86q0n
RQKn3MUF2lQRTui1nv7aw6HJIqWgZdl1wm3GeXTjup1I9y3D0G8dB/smq3QTmYTaS3zcbppiahSp
Tw8gLksSZkCU7fNFNqq++EYiFAw0S//rkRGrkxCfX4+JtFGGixHyK9fvGYu+KRFP2Yq1r60lHjON
7Pi2pt2uM66daGBIwCH1DlP9lispXpjuoi+XpfVzlXGNKz4eO7V4z6id4g1NcnufS4Bvojzga8kr
cuUTkl3TGA4MrTOS7suJ5CDmVZw3xvgIcK+SBGQp/6HcQR+W4qSYJ4UdjH+v+MlnpYCfWF6zlSBG
B4lv8EwFguonr/R8RUbUKPr3NNa7CKaEou7e+qCjEuZaa+L1Rj337yKduXSpHkEcb5DhARq9+6Lj
syCcmsdl3pyONbnfgM/z1itzrjB84G486W1218Sl0jBSgoWPCkVNG50Qa6v9H2qdhvaL1Wixynp/
bsqxK0rAf3DJ3YCGWOY511xyEoGNz02FsgF/GJMbwQ9qw9PDeDftygGyAeaGxQgL5A/SoBhgFsQ3
z3wYQ2rWmxuCzL+kfi1a6TYe9CmL0JfaiFroxozfPad6ncDscS7TkIPp3KyGqSE2PdnYbBsMdk7Y
M5whOv4YyMTIYeNtkXzHyBw/Ng5ZyLFsWsuAiTzkBSHy1nRmY5fDa9dhdew7dxP5Q4zYhbd7sOhh
PX4jZFw5UFVpSruJ6i3e+2V6yuGNcP4F2BEtQwPsFkLtRYGsp1UDq+xrzfo2vNE0V2ShwzckAmRR
pJKvZ+c2uoIWRnHgS4V/tVMI98Jovr07daJQ9cFTOK+bwoivlhtmyaT5ugkrTwfSO2ZktfyzyNJu
BXMDll54ogLASETBFEF60bx1q/wy8UpVKMV8Of37Eb2evYzyTLiM5RG2PMzkGqmMsYMoFEh7SiOS
EQ04lIrTfMnO7X90rBJI59okzw6q0JOpOSRcoQ1vqgdLLveUiYUfwYo8z4S6I7PrSCav5xwE8yk5
smXnwrCJqzpOAjxSku0ciGjEtnq39HHOLubbrdbHENvUGIZ3Ofp6jc10yiBA4Zrt30wicSXgTk3S
M4Neo5R34QyJm3dB6YRX6RvzcXlk+Pr/Ut74AZThI0nvMoSARsMrNzdniGqkvODur2i3mwkn69ki
gPACuDeW01r/NE9jkBHWd2mBB4BTsf4vqpRm67q9iAlV6WsT8ucjBA7ePqXCHSlViALgtQXzGOtz
hHNsOfpVOwZ55hM7VRbrYDMTytuqvAcjrMfeghdt7M4ePnkxZaO6noGBphj5RYLjOB+lk9LZe42m
2S4+HuL+lcutghTp1uFnkBmnemWir6M1ATjYkH1Pm4YqCEw0dxp26JSafI3Mzt5V8oxWzoPC/N8n
DD4qgvfSWLnFyUUMGya6BhuzlqJN2GstYXgmEayGUaejoEhYGgakDYTYzukXFMIjNHKcm3ar1ZiL
BKHkMF6fGFZhXvbRi5IssZ/5U1PWXIoG9HN55Dssf0x+G2ObMtAiyMnEV0usPGDnk5iV7VcAn3d+
21su6UfGq6NYIyc7Di4FmATDqq0JtXbb0bo+xbfsJ+Umeg4Y6GTVKFYJysbz2N6MiVsNyb6C3ktS
HnCSZVvZd+0uS3emMrTy6U+gpvvJGXxOKljjmveuVAYDaecuDiIV//3yCY0MlpJIQ0SfPcEF075J
9p4ZFDY1dQ1D3znaG1GY2X/ZT5bXxM94T+thsPePnrjE/Jx2PWpqndOH9575eopvdQejbrBDO46Z
dHEQuyvAA5yLwXYuQCtPKUSEUBESlKtxXoF5bPjzmhu9qgqVDMe6ZmBL2UmGNd9BaJD+poe/62ZC
7+P/wQTVLOtrdfqvqtF5JYnbPQubt+5oJd5W2LV0KVcQc5heRTIdDytURtD/Sc2HDHi6t67vY5k+
kkc3OyZecSuBcNC0B2m4HJFwjnriaIjAT74xmODnTzQmPkCXpRwqOGfh6Txh0GYFugv/y2xEJcID
bYc1lNpgob/6A4ZiFxwUfnP4lPjEBd65BCO5u1f3sMNpLAu1XioQMZmfqlLtFAm1rwc2yx+BrPl6
U3gx7/osesIpH7ZIgdekDeh0u7rdhJYcJjnaB97clW7K5OVjof5ep+0EGTaIaD/c7llbzOQ2Nj4l
iT5GwbV713Ot12kejfKZHvGI1neU+jIuIQ4s+nLDQDnx0IyPCF6uns3DrP4cT7Qw/amn/KjHDdiw
Y4W+GB0NpYJiH9qIZ8lThsuC6CXt7J2JSeH70qe7mir9TwtCCgHvH22VDUPzYni0331hz41mv66Q
DhbKUJgdEWHy+T5sYMESWp8/3jICVU+Uldq3BqISQ9pB6IMvdZmi9CqzNoi+32RYZcVMsVRBZ4QY
m3tNQ9rB7f7//6gBREB+vK8ppgX+ZOCjW0hhl2Eg7fRP5V2/59ZfZC8s17Kbjf2VE6SEEUM85ORa
Ac2K7iGo2AL4AxNQtuw4AMCmRogZ5wAnBcxQq5QTSySmtT/YwyTS7bxprbmIwj5ivgda2UiMLY9H
2Sl2cIluENmC7uXcFT+r2qYkNZ9Sxu/X/nKwo6enKdFWKsoiNMN5ZAUkd8Du6pGaoKBiisxKan57
udh2MFDn19ssdXX+kDkI91XJgCOzBFcjP16JzWPKf1+3tILx7dPxudwxEpCiHa5uOOo75xMefYCq
KGaoXuSpQbe0zbl6bT51iOx5VdFBdq1ZWDeHwU6WSruCPqiCuAihzvRaEmmIsqa965kZSUKrEcgb
b/nWvy/hy5dQZQFo9oME+yTDVIAFA7Up7MOloIfRhl5bsuCTP1Czb3S0B0gZDzW0mhRibipeBeWi
1U5TCoQIC9HzJI1pLXGR7Qa3AztdOwo2xT+iC1+7PStHFB0Ri6cH2W4dvCDYA5YgnreDgOMkFywK
0/AqeL+WXUizumGWRBBnbUXuaSxaTeu8Aj2GKBGqAIRhbbbmx7AO01jq3jw3rIv6yOgG0mOJWrBg
g7uTC7mucmZ9KAveT99IfAsWCpLshPVwKx4vSpkEgsDiaMIic5GxLyMtaaI27LhjK30mta4LaJuy
bAqmMSkKA4g5iwG52bUTVQ1MabVARdK/vh/lk+dPfTqoCy08EVHdh/C0IwiWvh/dz8O/ek1jDDNe
wvZ3PcHg3Bvtl/VoXCdPaLErGrAdGJfoLBMbuTwlvHQn6NdIfd8eh1dGdvfDDYUVnOGpg5hSB3o0
kkmWQeYoiJYH6zQEZiZabBeLUI4lmadJP3bbGlqHXOaDiAmu29ZK7SYe8yY9Hxtup590bj82C+27
DSNXwaqt6ouqldEtaGVzOotvszDSWhOxEGROo03tz6u0Jdj3orxFhpZukHx3G5SHI3uU/CalFt6q
UEvVWTobfMubCiK4hH90AJeWKxENn3TlQg+jtsXTt7tj5qVYk2jmP+ryeOvJS6viACgmcavq0dO+
DBFL/VU5g2OF4zyBeib2uryReA2yMMNqjMSQvXS+a0F0zEH/qHb2zt5zlaLTpDbBrKEFbaHEAcX4
fl2MW58Pjp35VtuVJ9fLtzLvJ8Ak2eO4lrg0dw/c5H6mt8cR3Q8554+P2aSKFxNpsSqrhTtCmN+C
GAQfAOVD1iDPMX9yOjcbzNJ0fS7tj/6eS/g1nma09offG8KqVUgM4XYFBn3VCUfe9CW1tMIkj5mW
lrlt7QwVLVUU8iwNn0VoeEAHC3R0KMN8KQSI5gfQX0OVKPiYHu3+WzJkUbxwklIQSGtVQ90ZSHJr
6bFsMX83NAX7ZIHY/ef8qR7xCrmHIJyLGAQ7SXjZB9B674RKwY4cAdCGVfrfaiFvfAbKEShwUGbt
A5CdTiSyvqTbyKhXhQvfjl0rIXUY4yMxbgXvwH/dfuzPnWjEF6f3+u+hJ6N3Pi47OVGTBXKEDxAR
Rx8S92zFWFX3V+suUhNFb2s6cpAb0jRq8r5IIGymTGgvXDLLjGwyTz7DpXu/ZgMkYcio6IoE+5B9
h0aODOktG2BInERegGj1mI3o8qGWqtBwyZQe6sywdizySlaUOcwlMxnUpPDApnYqG6VnIc+k0KoY
UJ+XPWnXag2CJTGxj43ecUga2mmNawzjBxKkAGrz8brd+eeFwoMOO6myPSSpBHdKdjTR6cO7mjpa
TiuYeY+NEeJ0AP08fwGeMqrbw4X+tgHtwLvqR/d8o1OY7aLGo4fc6pz5Lv65thclMadXC8hggqoN
bmn/Rc7HLo0OPqFnpi6Dj1HTUCh5uzH7wiH6rO4LX5RXqSH0XeYjf2uRBoL7+M2jqH14kiAQkZJv
6jiN6z/MViHBZlJEiqx5iXzLWU0Elm/jphS6iIwS+HXZq3jv7KnnvmOfn/oXTPlAurAklmBxvLEy
qdyabm3J4jfmiaikslGCPINwsL34QgOQrFB3a7yb1HdbN6AIldRrIlarydwg74/0B9zvfKemHTew
ICXU6CMMgEcsPrLQgbRHAjZvmBgg5GIXaIvlxoRdsc8hwuK8XSS+TwhW9HhyKvnr2VA4I4Alj9o5
z2nysbInwFtY2LkS/ENhkJa+1WL8sB4SAuZVjk16xRX+4+JpISg4s48Q/PBWqLji6bP/C34Yzwia
V5kbxolhRjGAtd62oohjNOiwWMj/W2L5WZSCxFBXAFjXPrpXEBGVVndwOcBT9FibwdwoPQhdIqOd
gBc3NNGR+XLWSzpSV1oOmjDkDOXkejKvd2sXcexjBleloUn5g3zK9bw0+OaYQ2dC/m4YgvHarfmQ
0mGfewVL9yDtxC4++GIQzEGyMOT9LiL37osaeoqlGMLJiRTIpQYxPlRdLI2RO6Jql0HXrntB1ALg
vtqlsnlOwDxAqVwppSNjh1T8VedBwBg3BZjY0vnlif8VjfBJRXQI18vtNJYxqvgZ/jIg6OgPJRYs
3lhWkBMhKOseC6VxvgSgDJh2O4gOHRYnfKcBQqbUVEGAaH64mFpqmVdXOz56OKFkwbS+IC0S4WO9
ZmJmkFzvs2ziNgN4nIxJAn38/CyXQc+9o1g2dmMh35MaJ+NCmmbemVZBlQBhovv0DI2xn6+/RR0R
giq5BKjCO6ttJK9PSqZtJQnj575JxyYbSO6Npvgs701P6b0Em7DiMe6kmojeXcKx0m00oO5Ec5xS
x1y/i71fEBGpLqNz2nIYWRWvKkgFY910hhArt83M/iE5IQ7PO06sJedToVDkQO6gNEd19kW9W9it
6UC6s5xv3Uu37CS0V2TKgnrhJy+0HDTexLS2WPZKefQ/QyoNN2r8+PT3OeaWBpjMmXNVQE+Y+skB
umOac2Zt5YEHB8AQkLJnhNzZJ+dM9tbLyLo10nCkjL5fkL66xGuLQm+iX987FSWPgH9AbvQkGFb0
na0wsf8gBsu94yOhzS9unnDrS6Q+m3OGwVTvJA3nkS0DeLhwEmsZGyiUXQZ+cCRjO8oKcqGVAOti
L/5fZY0vu5iAI7hOjXFMWbfaoSbx2Riwk/lSqHVO9QSrr7rtXxEzvWtLMoAhfj1b52zx57dU9SXL
A9a6gtCIfOsJW4/+nlDDC3NOPnxsquHyQD3Fzrb1LXOp+lo+ghNWrZ9OqcXlsY5sOlRSM1iHYc5o
wFYC5qw+b7F+Q3ntzq1YEZxfyn2YGdkz82wgE24F/JTdonMa+0hY1YrVohFBvgte92ByPFMOOvW5
MFqQqgCauaNHc/dHtB/f4VzyPwWEPDiF9GAO+3v+8sBhCFq61zLqg+xvBo0pUq9VoQ3i6iZOWDER
w4djxmfWI7APbHpfUfq8Mvv/vbAB5k61AMZQtIkYaxYfSfdYkUgKA7oWiib+w39ISE+vwwyW57WO
XJuAi7EPPOZaxEKHFmdP46tX7ZepB/Q+thV8CbaEcGCcBfLAaDglIHmUx7sevMX+N8hN4+LDQ7SK
+T9zPqZvascK5pkIW/KAdMrFhy4So+4oYF9IFcXlfMYbrcmeIEaXHyXuo1C7ydVEcN04lFOg0Tij
87yskv/O2eClY4oGXAIfI+C/4Patqc/3wpo9Dul3nozxn6NAkvQ0zfo5aHubGp0HqumMiQghw8cU
v2ls/+dZuCIASdiTx6HB0QTVSVZ/ibFOunBt8L6P00uJFVgP8HQOh2iRON8v4sKk69icSwQecpKj
iEVtbuByCQr8OwTn3iAvSQysebHx3PBse5gguEu9k7NJmqBWw+EWx6j7VQF3d0T78xvErJTuIYeZ
HrzQZprQ4ffw1G+kJfWiYn3SxHRXlO6RtbZKVT8pts+20m/6+zmYURaEb0sLbCz0a8PUcFjT4V1n
DTerwuOi2CstY9RY77hUHkg8QX3czjmfXTnMfgYZRYh5BajwXNprv5ZhH1F0Ruy73l7+G1R4yMsb
EpTgYxRH98rKSqpo3zH00pFYlxexsThlthW2B11bTOrit4PprEITLBVZ46krUmGg3gqTy4ZLpdcg
gw6Jt7LQBJlBS2D1Kn6vTs7zXltE9kncUSgtjOoCxyMfK7IdyL35FDS3dFUa1GsUYX6LDcAP2qHk
6+gZQLt71HkzLigVFLaLjPTp2z83aZos1dHnJLmlzhxYFlcIASVDQcvVNm6gVbXFrGOLeYg7z1Kk
U9hZwHdqBVOJ6ioaKpdXstzRo2RKlOKsPbTIVuzHEa7iuTv7mvZcUN7hRp/MlpsUUL7jKG2jAZ4t
3xCVgGTQ31jwxymUgtKes0wVKKh+tETJfJb1OoZNdHKVSrd5TOt60grWF4syjg4RvYVi858Um+sL
Ubz4ikVpqQwQs3Qqq/hMrSgsUMWflBfMA2G74u+rOt4ArOxXCcGAm/f+yYODboMuQyrI6ue/BX9H
NgvwStYNiY+n5UEjCzVvsmRzA2rEmpa8XFvxTDX8/pLsdiqzp0+vBtBpoEU39bt3K9nksg2XxKx4
BH6BlSrANRnPFzGhCzEUbUQvWjSYVJ+Xaxr2x2oXBWvosM0zacDYk/6ZkfUrYh8FP0M3fUpxz32O
TEgAKVNHSCG9ejtVgbEL1kQF4O8UemT3GgrZWBjN5jqHu1MFP19iIm8a3gEnVAPHDoNdqqXRHSA+
SD+8eKDaJYoiBBQ0CJWkvrZ+PCS64QK0EMoJp9UerlBb5gFoNoYycHEp8WlIdg1i+5rfm0MlCMEk
q66mKvh8etkUvNCA75rbaVWqD3rZpRltpzSNPczgXemNW4QFz2lCJaieexTXKgcdXGPkAq4wu6mX
+EnbDZJg2f6fAMsBq4jpehUWMlkATo9SOno53ZZE5g/dpIPFllrl2VDT1ZfMGHORnZE2AlQj0p6a
B/kWI++3yZyN84O/UIu8CrDlyJOs8jlIZ8eB0AUZPO8LWP7N7TPptodmdV9yl2EVHUCfKhjA9mde
4bHVqjK1d1gaWKa+7kxX9GNHkK53HrXO1SaaKPuJyd5wn5fwB8n6GlhdisuhPS8WnKc6pAGxkDSL
epFRTBUMQdrJPuZ/quPo5Rt8Cxv7QhjxemuKeSYCD6fllBZ/4dxF0q7yw5QFqMYatsmBoK9qPkm+
yqoB/VkYTG51430+eWOerhr8NN4MCrwFDLUv91rJjn5DFUWn8FKHR6XFctWPCsscACkCWuZUXkdd
Zrc4R3qw8g7nWAmOclRqR2LBVR4o5N0/D9p4ix61AP9T0ZK26/+ueXk4BBxodxzDjHLJM+2N5xL0
sOYKbCXZDuexBt6Wl/9f0cKhop8eSoIDca/3Q2z9jrfp4Iwhq5XkMTYhcR4DG8vivmczbP0NzYfa
WW774FiNxUoSSmI+bzTWXXmp1ZEtiYikL+bp0x3/1v6KEIONZ2pFwB51G7MJVJ0z99w2SDCto6Ew
Y/UngIobiBncZTDPH3uZ2jd8Feschy6ViuRzDdAU6IIIla9FEa9t1U3MpYTI/qV8Tk888ZE1um71
xBOJMd29aBcOAhz78e63ZU+BAycRos08vh7O2NVx/XR7fUPRhjdAk/w0hmFPJjvoIKOI0rSB7QMc
vTInlsZcknuqByv9JM8+OMUsPve4Hnhcp0Gor0ffh+2xc/2Mfu6OVw6h3fRfea43MjUmb9Illtxp
/54nEi5Pn1DRYgMj+nEWzexBtxLFJV0PVmwQxCdpcqXo0EfPwclHG6FVYdCl4Xr7Jrdh0zELg+ni
ZctMzR2hLjEXsP7qfPEEYBlzfsSY0h6gRybUDwEGhNU2p6K5AulAJEsFvhtge8jfR5GlT3Os3S2w
N0BQYiVN8z3n3b0ATYIPCEaNNGgXWiDFWOa7L8/MsxJUJYFSq+zL2KNNboTXblU5ymuAwl6dLPml
TuEWLXkRdefbvR2+le+BBTlemSnNNxsTCxSv5z2wE2uo3J0LPdD1Z4SHfcvE2qulF0ACct5SwDId
bVX23W4oUOY14YJoBk4wWdreVkJyXDVGjHeGiX+QzVs4o/fKlCwWj2xCK0elKDDbt7Br+iIrMOO0
hPC57xzCIrkM8xw/EH55pq62NS7UySzDrZ+nfVvjmctZowFAHrAxfWM5ax9MawGBLpfpUblbzCqk
8WvBGVPdm3mMKceA7TDooPnpzJGx5RwRq12p9eBZCkAjm9XpQ3oZ0E5/z2Kj4/Oz1Dnqd0yNb/eu
j8XrYzxqCyzkkEtmqp/EazT15h6SfCgV39RDsY7/OyrGAaXUMV+qrCVY5kZSNdCQR2OyqZvFOlBe
VyYodfAjiaSPwzOQpACnKSVqBXLpJiNqbzSBiH5O9XGmYCDCqJTzcxX3UHMg01VHf4/EEOvsh0rv
Apv/cEh2CqSuqIsZj3Sm5+kbKz+wwer12rxszfC8pa9+BKnTvH1KK1p31dA9fsYvHikitqWicnCn
ZdZTxmNlZt7fBmg1n8YbxadWQhAHqgjydl7/WLQHlbEp0sGq25zh5tC3ucmnW/KJ1RDf69k7A1aX
UDNxCqUCZ5D/mbhpyV0fXKfnlbg/4u7i2CVoQwVcAofiVH3muOsh6GHNJhvoIYATo66rh9X/fJsr
PCpzqeKrDbb/QrocCoEmMkBwRNbXLCG/6m4vwTJMYq9Dnxj71ARvf32wbq78PGrUhYwuvMPoAulr
Awzovsw35TygBbnkYDv+zfxEx+yX2tjgZpwgO3TS7pIsaZF+ctk3RakikWpSObhi7OjL1oSNW3op
4hpzEwWNn16vRFrPGiWvJ+PzFqMIqQcRFTOYszVeZL7ZkS7hJbFMoProxdUD7LEB1v2XM3x4svF/
wpo7NJMl+3zsDYjXpO/HOE+PtedmvianbhcON60ui0kbqsZPts8Un+Rl6Ft3HDlFIFXjqPtZLVeQ
5JStK4fLohMkaUW0dsFyGMLsfTA5tARapTsU5uacigst4EzCsIyoUaGXgzWp61hrK/U8cXrnucww
LqrtMi9VjSRmeOIyZo03NpTbXrOrTtKXDrWQk7sd2CKlbYMrjjsCtRcbEtRZDGRCiv8f2PRrEgeO
XxU85gsVXKPMq5hn/hbESo9hmRhWhffz7A22/yCeedRCkIl8prIgzxgbZj557B2zrhMaQZobvOw5
XzV7uq4jRwoOpZWmuWIwyIMqZg9wRBS2zHZs1wF6cob4gU1AEYjGeAFuUOwNX6FOx9HJhdXvceKH
gH8w+tnBnAq9YWX8Tn0XrbOjdn5kqLUt0jjbp75e3s5JpBHPrhZ0dYwO3NyVpBUX9LKVhtVcETb0
6Cnpq2Od2Zduy9YE73LPZTn43r8l4DMx6zpIImzxSm50l4qak+TscfVt5o+7FO8XjGLWBpDjxkGx
mGACNzWvJoAeCmi3znPgkY03AZvJzayQ/S7Y1oN4vAP6m3g19iyxChf9AMmDUB0+nM673e5MoWFT
5lpqoST245YSZ/ZeiIWzdoh/Hr5aiaURX+odaFk4tLE7IRGKu8FUsuLHWL9UMaBF0FvIuvA6WQpd
BcmzgU5qHS0woyWrwjG1pJXrlYmw84ui7MGI34zVk9XqvTUtOM71DC9mrJd2Jt4gNCCwe+yIfhZt
SXQJDkZ8F2+b5Q9XgPJt8crSQoHyyC9455zCCeWJ4Sy+RpHwkMui8xq6eVty7ro83Hn5/KdVDn49
Dx4y48K2SVgi9EuT/Ip7NSD7K+a7snjXC2/WQCBsddwMQMPqyF+ZIzYddr8/W/+RwVYUHgG6C1Q0
9wskLqLvwqAcC3Pt+n+XpZQvpEpE3ksIB5rTNs7uDK3bBaMJEecmsCNccYp+84UGc9SD8UMFvvHq
e7uVw0fUX3rnvbIg3M69I+qi34HSHJI9HMjrMwAwDsC/1LkFT3in2z3IvDyU8M1MwDON3FTxNSJe
5fK60Zl8ceArgQt0TMR99ol/BAeg+mk2ie1c4dGJlVQPL+WA3g4M2jHYdhBt2ZNVH+Lm0jy3QDCV
eJmwsGwiYqCWL+ckiuE7ir1nxVuKnmSGGMVDuHLCOg03d14fw9MF0Ftd7CK7gxHiKd9Zmas3Hvz8
BitK4LHufaDetVk3a2aBeDwA3oF44fVv56Gi2/+1ZtUqzGXYjPYx5E7LicL3RFVQsSlBQ/sd25Qd
Fig5mBZnyUGfM0S70HzJD/JeeNK3kah+KJAWXtg/PCSOaeBDD8oAU9AWIfQVmANbBUMIvEPho/fQ
v5tku3V6B3MX2gZXl+L4f9nhp4CMyQTZz9eYS0RhYWJn6X0Lbr2FYRiJncqcw7rlzno/1ASWt1Bl
iWWwIgw4iweEHm3Xkg2AasLpp4D3Uf5ySJjc3POSU6my2+GtYdASCiqOAqiEt1tqBEnhGOtOLxED
lDeqoBBhTcks2JN3Sh668Ff0+3zO9RD+gsj8QzzuzTp9TZ8MkNfe4d8Lk0C7PFgo8JLxpNSChMnN
FVcHJT1w/JGcLm6VW9zxN2bh5UAEQTiXQRBRP+VNP4AOETbD5idOZtPrg9/+5U32PO5SOIPVdXd8
+fMqtHlunCpU6BbIBl8UuQ+5KI45C/t37pocbT+Fj32IBmBXYSbTEkWksQeKCjf0XyVSjExt9uZk
lbUrgY54k17+H7KgZcgkTyIRGDSpZl+ho3pDNxc+692NgnxphCKYezoy2IARMaOX4HKFkoh4s3fs
4P5SGr5GYiLGvV1xLIdJ5/1nzaqzxKinHrnYoM2PJfnuZHMK98iQVu/fWkefMCooFZO2op1TfBvx
WucrW1QgZZfFC7xSLzt5TyRsWVWYcc7RS5NMQj2pv4ov7zRUbFgvHCZ3BjBrxFWSEGcmpC99eZYc
2OAHbfxb+yB3lkKNMuXK8wkA7DedDwRHqR3lISPdmXVCxVJYeqm3qNZyBnRujmsEL+EfjBgAyBQp
DCkRTB5yfniZWiqfX4AK4AUYqc5o/vXajklK3c+dSx0YceUdPw2GJtHDO9iiyQLsOuxURYp2HsN3
T5o91Sp/ggFOD/b7P91b8V5WiWFQcBXIYN/vyCTCB3BDSm0U5PdbWRSnkT9FzoPMZHRvDM978AKR
RQRgMVs/TGcA/rM5vUBK8zlWXpMmDTTKn+lArjF1izKSBh8K3Z8fQ2XM+uWHfggiatWt1YRuvLIb
0khxerico8OiyoF3qco0jkzD9LBkaCy2IXA83/zTGnpJHUwwNQIeiCgNAyIUuT6kanmXH8Nes0YE
4QZhsRxhecpZg+codkwqYbFKy7Y/O+sTOlI8U57fv3bxRCrYrQc0lkNfMyrkXgh4Vx5vRKM+iA/g
G7QXfqHc3UygETOpUfY66ktTONQn6mS6lnzN536dCVOftWHUxPQqf3THg3dlVK6EkXBOa8t0zOnj
Hl8c1CylcS88GONvoAhJWKNcmCzYElH1ZU54CFDUgWe693dHag8+f9AYX7nmGjV9dgLlRywKMm6H
EL1D1Izp1ks+ty0c4f7W6XFZKP49agoHnKTqQVnJ578m8iAhoiVAJv2MlOgLRgYIZms3JjBcY/zb
FSXLaCzo2OVUobPjPshymOVzQdDOaVlsIBp/ndWcL3t7Jet/vzBLvu0BlDzGvF2rspC72eCSzQ59
kaoG1TjeJNnjiFguBjXB3WzNwHW2kr4maYWHJKoG3tr9N+Rj1cE1AamI1vD+Nzy8CsCHq607r3Xq
w92/OSsBoLJ9TMKK4VLRvp5O2yZfjUnbcIVxkRSGK/hJT1W40H6mfQ0ntrsXEQvpgPZIcdMSPso4
clCsaMgJf7p7DJMWT84jD5VzenAJaZxScx7KkM0HpqtZIoHLRxchlpZZ6oU0t32gFRrhtu8bvFxa
GjLA9NdLcXV2umJHnjOXVe9/cZ0YFWRORfT3HZyv2epz0X0ssbdvV+WG/MMMXTjLhANE7KBsVIbX
M9U9hJOGvZfVYbt1pcTliNlyuZo3SuL5kkMgI41R653EWflDvk1dh5YMBEY7bq9ccoOEa+QQ75Bq
5FU3j82OB+UvjxzVTgNb6uJdY5CABAVC5h+rpL/vrExyfHOgT5yzoZaMW25L5OSL43mG6uHP/qcQ
o/6PQyzumrt22BJG7c+mWXnIHuiUXJsxEJamOZ87BS4WSJVDo6HMcwJNCIhxVuPfLhUS2ssrupyi
bVt44oZ3gbPRg9kDxEEnUI5bBlzFr1OulMj8pTJqhDEVkO9H2W4UM5pODplopakVv/IrbYtEAOcH
x1+uKscL/Y/BiZnykVFtLseZiL/b5K3c5ZIAI0w/TgmkTfCSVrr17pSQEGGCpZdcmHVcbV0/nKtJ
fjci1rATgPBqJKFrVu26Sr2aw8vLkuTT9fBuC90dP4zoqUEwyV7rEPTf4mzqLG0oKAPVsd1Upla2
hmCcM0EB9Qx3kepqNEyjCjPgpdoJAHRGEQezMonMKWmB0bYQogtzlH0uqO2codVkVIbNprM922Di
Xt6R6/dukYDomQk9hz7v9yLlixlode4UR/FlqOmBE6jiU/LBbnDl8zBsBWnJn8i5ox4XmPjh2SLu
lZlNoEA2nzlmUHlIJv0dRFtSZrhtOuKidboLLTQTlGtsR27ZP6Fr1wQaicT9nqlELJANUlFB7ES4
ktFkM7p5nt1lIwpYnQl2Q63xWr9zo+vGGLWCOzMi8itkQNE3AT76R8RpqFoI80DTO02+00kyra4w
8B4+6Aq/zWsZyPKe8dIcyP1xSWCy/mo4W15XkpOx9JobhXhz8dLty09IfWetE7PizN5lwWCASAae
0tK6z4gL8Ce8K6Hg3beXkXLnWGqmxYNg8g4TAXQEOmlyiu+Sd0bcNZ4ivhaJb+ik8vMvSpi0CYmC
n2pg8ByPGUJy746u35ctNk47brpySP4tNzelcoavbdwsa0/NKp6AZvgAzcLF2ZgcScHz6HqYsDlw
yy1OuWk2aipjlOoH1vXBll5u4SR75xS5/kmwUUFL57yFwCtU7NJZJts4IX3IEQJV/GG1aLjvyLs2
5CWZxqpOgylcc8IdOv5s1s1uMKPJ9VSZg5NROGOfOeVQOruZ8DxBNDCABj/ku0/MPGVIRJjYNFuR
I6Icgfcfa7Whj4ej6CFD/zAJSmNGALu3Pqbj3f4Tosh02i2WcTZDxHgDmrGw/cIPIZmZXGXTTeqU
Q83mXLd8I8yDZnY6FyEYZx7zzfqKovmYjULOcK09EgJyo+0rQg1TLqgYuuvQ/ZFMix5VydVEzBSE
5jvGcRgXL+oP4atAtlxi0t/RP1/fN7LFq47tWvhS9+JDb8Z9FtLjbNyWydgf2yntPF7IZqmKeV/a
wMBmqlqiRo0Ww0B2W/ifhRIqnKtpp4awahsnXPFFAFzq0V1FojA8dEDFiOAdvjGcakY8TAnErvPt
NNc5g863UZPOuavZyjmwLxp7bsJ1zm7P2sAT2Z9/UTFAog5YiuvUgN4EO3qCUoz3aIxj55E0pNvU
SYPsZPE+tB9IWfmyUkwORUmEe8qwqx2d7cZ/tO741FuKgidD13VH3Gs22aqEusoT6gkx6XxdUHjU
CQT6l44Rkz9H/8JforOI/9YI6WLoVKSnTJZuITYBzTFJ2i5tMCeIIPCxZ3YsmzlPwM+p0I22j58t
WpMv93mYkB08htcbtnLJNEa6Tub1zAttOj56XGJI/xAc5M0X8w5Wo5BPrfNBFtd7nZKrdtYN9b3w
+Puf5YQ90T+4lclDMiKotlY6n6ZV3Bh5LKGSikLhaeZqKhal60vi7mxA5UB5eaBUB0QmkiEfR8jf
1ao7tEFyRNXa4+nSHxTk0C7tIa5B1S4I9gs9H6OXbZ9Lglc8b11rBXOfIvatnkqmXQYgfvchN6pj
Jkg6k7Onm4QHMObXECzHIWibZFLR3W3t8zwd0ueXdUH7yVv2zuDrSdjFAcxUTvE5cAwnobysTF51
eWYmabUfYk+8cqL/iucVHJJ48mjLkwDJ0jqK3Z8N9V1LCawHtFrF9/kidJRYFZiRRM6Lpe8BG3Rf
KTahcwykBvQsvqqvrAV0a0b83nfvvwCUJraGQYCuG24BsdlDt8wmSoIzrQSBCOkisbzUqWV9IFs0
5cy0PkmGYDhyP48wd93a105j1dUKiejzHLQZez25Bnc9zmgiAunh+ACKDOGzDgYTMAmyyXlRN+ep
JxFw9E2EmUyWvUhWR0DQJN9PWAc0Qh3GJfslW352+jkeFKtYqz2Tx5InoQ0ycXPDVZk836xXM+P9
cXeSQUwtJzHXCUdNXrpR3fgIJDl8YzeK+GftleuyDcE5G8+/lfuyThds/2Yh2vZJvle39ZH8MH5S
gWM8uUEWo/c87E6/RkDRy7mwP1ruHUUA4SrXJ/nzAzctTznJajxGwPl+2an2Q8i+fdabWnx9Asru
OvAX2GFAY3wccST1+Tqbu76HhphTTl723B1blliBNRy3dsXGdvollPj2WRaAfr5Q3mtxq+UUuJHF
S+ku4FWyiTn3uj+UgdCSXzyudY4UmEbJ+SYb7R25tVufZHrmom3KvYnLLZGSoGb+DTN5XtAKww2H
tzxKdFtBEln0QFduaYy4JqfOu2hKYOTloF1mJYmW7ma7F3znuGNQxxaW4pLNwCQsc6WiJrCzDTyt
f/jqQVr6F5RbwmLgpRgsoNH4wzm1gnOnsGOBYkpmdJbLP0L3nNUIvEulETZwBl0rJn2gf+BZNHp1
7gijgvtBenS4Ecjxy7gZoeGhQ/SCaHIv+YcIdYQi0/cJ5vF2nlb/3nbF0BgUAiwRHbP1KLSyAg/i
UvOjBSLCX3y5v6JRusQiaWQ0JtLRPBTLlMytMlf9/3t37RNB/7rdk1yxvlqNxT0/509txLCLU34E
rXaJO0/X0r5x5fPrQlcBmfPP3b8PazSWAdfUZV/4oXEzvY/3t7+GB5JdAbHEXV46RCTrpNOUEBeu
dH6dM5tKEosW6h7jxovwyk3JjyaxRs1VehJKE4GPQ62CyGQgECtunT9n2r3SehzcC7foFlNRhvDf
Wga0TPmWBQeta9wsPUTD8+3erwGcY3YjHjbWpIvNL4v5DaP7t8XJVVAMN8itf7+xUmYAHYU5zeRN
X5hYKVb4dKGL7F0kKRrMOzCeIvreSzINUZScf7oTkH3Y/BKTVhyBS4CDLruxqr7zZN1vW5BTlbHT
65FG6upqa97/mTWyfcqyZMCXZK8wdjLUINfo2UHAR8kJ3eDsQQH6AcN7bz5wK1AYWS0/vLitCDt5
8+PDF/ki1IjDACuu65EmF2RXf2haTPjvWaA+xI9eD5Qt8u02BVNujdF6/lyMZTTFY7LpXQpB0ALf
A44oTrorWqHdWSbgb0J69nxzM0+dfxCTc8BW1R9LxSjCrWttKjjJI6lXoXguqLqg2kYHxAlJR6V+
sYtz1mtaU2YrYaRnhj6HQ8n4jOQegqO8rhw0MTMW4ceT7Rb6mbvlhvHX+1DQ29sKjIrWR0yEHOc2
0B1TqOku0eRuMez8Ff4tI4EagsWfhFBObSRnVJdqVjy4iLS2p7LjzE8BH30WWE/wDv5JRIMr5spG
gBjKMX3l3W7n9e8FguNN0I8WM88tFAj5urNlY29uR1/ujoMvzTJQNXfiwgrjxD91wqu1KPD9sbua
djEkInw0smfEr9ELpwVfHFf/00P/kYlxA5Kyy9CJAV8jedMqjdqOaFc7TVNk3tFbO2dnFLpxRygT
RYDplQwrQYgO9t7QENl49Vx/F4x/k9eb+hGARhUWtZA/hfhteNdNQ1EiDoSdtJWW13f2Ggy8vy1e
kxKSlTpnTQoPPO3THxLDdlWQEzcqMxwimNFEZWUkP+rlce/mZHlUKUCjPD+MhDrdZ883nRUHHunt
mev7Rf4z/EtKQDDHdJRkFyBWo9V30r2W9jBQcmkkronKOpLXYK/m1WjymkmCBey0+7ggTGgW4F2M
MJOEtKMoxyGJP56zva3sRja7qS2Hq1pzuZAPAmwewqTzbU7gWq4HP9HaM9dXvMD2svOHPgrVvnB7
Fm1uI5RjHXZB/Is54Lnatt/uA+2uQ90/qrFopEzoKJqGA5x+qeM7lepg0wFEQOX1EXuhvVRW94iP
iSa89edbkRNokk/caUfOtk8Cf7N+zDB9cnF1WbtcJ5rACuHp4tDduCrs78aa6nuC3epVQsmRNDr+
OQ9JTYHR9pTLoy9TZGjucV7XGbZ4BuBlfJDwj9Hkcni7MYvArhPHOhJTVqNsujXuhlzyoJfiNafX
ClIjfagE18aQh2x6UeEhM75G1sWft+qWGIl3IHwN2AnY5AdpZU5xjD/lC6pPCgl2mIn+xCWjmAY6
Zf56yaUs4bNw+9yJnRdCClCp4QlcUuZXK1Z5nGt7MCVZyQI7VqvaM0sCCPvPEy+wBhqzBlWhmSGC
qRUMFlet+FCzqC5Dcq2LTR2UDdHku8WcoJgrDyC7TAF0l+4+9/+3j2aZ5kEkhGXhjMO2va3XIusG
s1U317imRqlOyRCh9eQdjYBLjpm5bv1b0SZ5YWL+Emv1iaAuOkRxiX9qmtfLTJL6IVCLPtkJ11Uf
E2wkXbxO2XYEIfUzKTID9UBWKVNOAL/Fqj+64cjEOh4jd8+Hd+GfpMpWgjA2igNgW+cgVWa/7DYW
rMNSabgfQE50Ni5MV8qmM2D+afWpiRCAudpRdwiLz8Ai7PprtwpJQygvX2o6hJtipUVucB7l9QFt
8qIV4qLa15L4Sv5Nf7OmXX/+y0lLD+Tp362lGlfAZZAoWr/ogjEYSXe7clrSUelu2qZIAFQTumS0
qKmkZYAeuYoAFbFnQhS+hHmGRiJ/wlXHg0uY8BnbtwPcvzBPm11lqPrzYHWpVF7Tk17uhPKIEeN0
qcaFO2htlHg1+RqYLrPfJ21hhvJt1judWqQ5xBW5rzrm1HmRS7lhAeh7k6tuToa9B8PJVG4YTdwU
QjcAPFsaqdgUOSs1QXErDKkqlI/101V4mSucgmQJqltbd6wKzcXrEjo/Th+/UlkaBjb05TvzCdNA
PeDNEUzGlYx75vqWWU/wKIkb0hA9orqsQpNICN8WLhvzr+kurX0kJPQpqA9PZx/S4jYR1jRvyrFx
lhfP/9K0O2ZMu8GoX5s505LSGCre9yqFlu6LUdyzjEu+zSNPiRTJ9GIR2A829XUFmHp+HwtAgPHg
CFxsazSSqJmmqKuz65PmG2P0vdPTSn1iXEr5DtEmoHxq5bDLnPg5GGglQhK0Hfu3KcY6ANZGOtV6
ikfOlHMk0d9UQmAXWkdNemMuETUak/CkCIipMbn2C3kIf1ItUaxDu14wEOICJv9yHykkoB6j66x0
Qdsw0PeenxXAWjt4+mY/65IAd34jBLqoufwENKc/6YXG9Vnh25L+PP0TuAL0yNmZoq5VlVjYRUhk
wB2AVIfqZGn+YQ63WfF8nbtZT89PguTdkisiX0bLSFplgNO8XpUmjUdX2kAiX8yoPpqP92rYz+pO
tUUt+6NBNd2f9cttdSvt2Kbdro3CrF5CnRavP2w0n/wNScC41CgHu7h3vPPZaDrTCnI91AjcuvsD
Yi6BByOB5oNR7Z4RB4jMM1YyZe92/dhZqP18xTywzc+JY7aAojffjqSXpVnXDFrVNLq7JYIjcklr
pvchPue94YojPHI3OHxRGg3pOPCT5QSxKY1SNFye2cWKy5Lg9/qB4PysANtxuLk1FW78d5Nogafj
E4vSErO5Vp3gkJedyPo1HhEjGc+oNcKOArb/+z5if7yfyt+jnikfTwbMPaqOxAbm0ZzopkyS7h+S
fXG7gd9RG9XKtdag8LJMlmQz8NXHPizD2Q3Y+YYDB2uMtMFWrhqHGPr6MZfhzAEOGewq+SwcBR40
+bH2Tpsm1ep7nKkSMN5pV//AqcKBzmOklnBdlm9u0Hkcu45YJ99jGlIFrH/pNrxkh18xtQQpXv+X
8/rT03hu6IXhnLKdlPjWGy7B4ovTZP6ULRIDkZ0ITJqKtdvrsUuSiUPhNvdE7idVK68veop1LagY
HWD0G7xMM40U+lvjeJemVRtsr27ebnBQYFnjdfYvx+vfYEUW+bPM6SmtQa460ZrZ0imFQwBKVGUb
wzEKdA1GchLYWCqplQvd3l89iw3+Sc7rT1koFaG/au09M9TPEioBbRIrK5SQa9Iaqt/F2i8dXijg
XD+7BaVND0xzZ11k0J5YFJVaskp+9aP8Kn6e1D5z73sIS3OGxQfGvhyBj17sABL149wWPJFltkPN
OR9e5mLdH2stDtrtB0/+Ro8tfRVVlNct6d5uXIQBW/c1HP4Flnihj6EroWJ8DvHx5lasSXEwoDcy
mMkXe6FoyS2Gf7yJ8Bk9qWyQTnDQcyBPGA2yu15xi3VQHjdzzohy+G0D5g7RjeCNtLvKp2aSivlh
1bVqKLHnMTm6tJFMFAZsUW0B/Dz4G/nU+jAzqzKsZG0xxT2kEi+q5UqXcI0obL3TaleXC+4KzDDB
GpkGjU3Ed4rY1STZE78hrgA+5yG+IDngj66IWiDR1EAlRAHEGJ4ci16caQ4183Gk6Pz6xbLvDvWE
hhb+wF5mv82rzmJEZC1EWmVjwv+kLQzWKxh0HFB/bW3umg08pn5I2fx6pZaybfHAHF2mLJM3C0Am
BnX2GCyBdjq5Zq+Vgyh/j+jHmr4vZ4oOFcEbHbzv/nbj10KafM8BM/X4Vu2ME/s0StR+WIEOpK7B
vKwdrb889Nj7tRS4/hJ1WbsWtKfzlFlGan+w0rhooA5iswGDugRWlbYcwC0IORWmf4bGh2CQugqg
a0u4WMQW+hpgJOftISL/lEGtdE2Ns72d7XcpPf6jVQHojNwnSmSATYyGL66Dx40F9W0we8Jqxhpl
384OwmBhtrW5EoHeQFSj4VWYL3QED0NvGah8Vgfg/ZUxUnshPwsAvYwa997dwI6cMH1xZebOTGW0
S6I/O98TejaMA+PcbmfrFRt5LtAiFGQ7SMlEaWPqU7DEdJjqrgBuwWG4acwYajPOOlvj9sJvVGfj
xylu6x//tIsvUm+gOvp0mB5/kb/oIeUIK7pxGuMxY1LNglCDEv82v7xjxC5rd1t6rd+NclhUIenN
oH3a+oQs8qWGN9ugB11W8a5SY5T8AZxLEZphZ+0AH9XH6mfIAn9+SDpCghGa0KUVXYOQXuf9fqTC
fnCbelBYyILmepFitkrCYUT622y/7sH3K5LvJHSeU4uxOAOKp+wREfgH7fITCx7Okl9PUy1wx4Hw
mHLMbXSD2qdHgR/F3Sh50gcexmqTIH2VFHQ9v4xXfSYGt+n2xRxCv9TATFpmmDRA4YKiDZkyXC3A
2KA5wiz5t3V9lPSrH6IHaar7ZhpJ0Fp10JlP3n6mEJjvuss+UBJEc5rhKM6MAb6Bl23E/WsUijl3
R6NaUNNpi5JGsYsDXCSv936xAr6uQrIp6A7htn+xIlvtdz0LBc+ThtheYnKiMiWU+jUP8WT3vT9+
AwmWNThEi+clhXPj6V2YUJnUrrm77dY0Iu9v+aGnYq5MM/O2UQiRfEtFIQhyrdpXc1QALtSSLHF8
o/T9RjhDwSinAwWrKS6maxZjf0DrKEzMt8vS15woQQcbd0WJIO7DAZyCUrlsh4DHrXFx0v5VsYHC
FZNBf9Cc+/pzhs/OYsgAIcpBc7xCNt7nOhmoGQ7JkUlOVQnsiEPvofu1csrdo3e32DA7qI9+Z3Ta
PlN7HlsVlcdy5YuXDEF5q4h/OUhikPbQybtXpNVLIaCJQCTnh65xdz4REFgCYGI9FcAM8lGHO5Tu
TeCggebNxBo638JytF9IU4fLGAPt+RDoCdn2HS3gEAeOI/Y3PHI7DRVsbzpV7K4Mmv+kN0Egrc4p
2WVA8cWEUMR0DgSo8TA8ZKKJIQN/UAAAIhHtvw491hiIUcGPhiL4yXeIr2urBly3rn5g3Ty2IZkA
JfwC/M6PZthP0NWp+SswhJEbqFSvD/aJknhfShDBR2T4vHORcXSeoqCyn1f2aDGa61senTJASFd8
FAQA85KMWqnNwc7a3EP4cmLF8OFpSrfNuJsoeRYUC3Hl9QgrKn3urqV789+tsMqgfFittBXgzR9w
Q1RSYvp+QHtzR0Hcvv3zBad8wrzbjJobcDwiY4Mm81Ykwptzz2hBb2yhpI9JXiy6nMsoAZMoG/cy
XgjgvZ0U546hVX2/0SaltDxid3Bmu4oqHE2RpsgMNVmZ3pd842nKjYQ0fx/KXhnpdkDhTNCHnpj1
ox4dZtQQl/gwzfY3p5NACj/1DHDgFm3bzkxCXoon4ESkjWMVTnUuqLNlF0VyxqmucDMaj75Vin56
I2X4+7vybrX5s+qzhgUu8+ikw5myw0xPo6lYmdNtcerpGDpxsKpKu5Uik3TitnMhwXrVG25w+NCb
w3PpSI2KuyE5LXmacZVvWsAJBq3F6qKq1B4hj3Md/o8GjRXB6Sz4mgwfSHRn0Bv0FlI1NpzCyx7d
DSvwOLQzstrGSv2argSLxCHIr+5MO4fSS8oscnFrDawyd8lIFl4W1g/BLN67ZJdEdfGxmcRknRc0
6CuLLMk818T8BosdH31kyu6FpRKSHh+397cO38zNeCzkM9N9Rb7jlhf5JfyN5bqYa65M55JNCQIm
4CSjEahcyBO7qnG8VFpUJz7cqQITQF5AYOUZl0xaq78esVJNp9Or8spdiDHEy4N0ecXASou9vGeH
51C0SrG/pn+cHOMsIxDd3q0i1LrKchmqqiXcl/rFdQBn5OrzdBLbHZ8xHDbW50w+oWlSJB00W5C7
vOqzz5h3W8BRfmJUcD65Wyt38IHd/9Q4x3DXzPNACAVmJnJh/rWrAoS5HSolUFBhtOiPaFzq0CoO
/u8QiTdbd0QJl5nc2Y0QMhEiMAyY0AbQUi7Dwylm+ilMI1xK1TKCP71tregovftFKzzx6yXuSHNk
sHtB/OxwD4o0SXfdjivclDCDF+T+JMc3uSvB1ujD4x2YJe+U+wBfrL/SG2Ax4oJBYTWGg6e9Zz0p
fjIIZfB5lnrCJFfNkaOOUkhEUUqE5MH/XHNbgR6GNY9UYfUCdkCvfrpROfrw2xljeeEc+3jJIO5Z
8b+sOzcMMDQdx2uSP9Qda9/FAeF90w3F2+UYJVE1ymhXi+QeBxVnQ7qXGDsfVEJKbATYcy3pOOLx
Q32BvLIAv5Ghbh+2iWc1MNpiwk3P10zEXSxuN6xRwkbhKIC/n87CUxXeGbXG5nL7XYes9vUIUVvH
94I8XR/wvx1UWxbfTDB5ILz00mMpgO7hGunc7JA/eCXeSjXeuck/vuv/VlboeKBJV/DvDMyV0oeN
n2aKSJiEBuxw5IHAkKdWbCTy0BuSfHX+/22FWU7q5ygcch+f6v2ZB+IQnYPOGpZPWqFXvERs88Np
j+06jQg/RkSmB9d3koKlwo6+rLShFbozpdzPjm9xYBhkxe3qQ7mUrEbfdctO8MBJtlClH/nZrZkF
6XOQ1VyuBeS4ut5ShOm3Nh3CB1gHK/4gEDu45u3kKaVrJozPoWHqAG2n/5nPiIQqrcz3ZJ3Zc3/2
brleeW+M8BLpfTH6zUvmnMUkd1mBnJ63pxIT7kxD4por8Yh6j2f8fb5JDfQFMroe4Gi5qrNuUlzw
zHkq4YIVqkIRCPyn0KZsdFj/xNSwq1CrCrYt/W7xqd61nPaZF16YL86GWj6XXYM2Vo5vMQnpNKG7
/YErtLwi++rqE2Nb6VVkHtGa1I+YwjPV488jHpQVs5iecyyiQFV04Lrts/wDOgiLIHTSbDCPCWRU
4sbFsjKq8vDId4JeNjUSOdB4rARVG1kq3xzewx9gbRFNmuFOhC95REOjzQXYbp87200+a5rqH1I7
yqh3sL2Vd9XWLlteUJ4HE5zuVznIantOoNeg7FXm7hBaOmyy0Oru8uaTHI/1WgG5niB7EAo9LpjD
5OpeP5PnGQwhjMEv4vLyI5fBYDy/VhKx9vXINY/5KEoUdcgybt/7QTqeN5EJTjUy+13v5WAbhepN
w6DkAK2mlqi1L2Cq/e8lScmO0OyPiK+w0U5VpsRKHFo8x8aS9EhEn4Tea+5n2LvuyLhzqnqemisF
ad1wkmDAZ9x16cRLqATmgNrcP/oJnzZebo7SOFblrxYWH9JBYPJecT+JXlOLi8oHtXVRACkTTji2
1A2cg078vKDl+gPsM2rAQSSHC8FXd8Kmm1Z2sP7FWZeUoUfx76egrb5DkIlICWVtqHLVDqOcxzd2
TFq3d7PYP01W17JjFMlFSXS6dpWpSfCdEi1BbGkdDkZDug89SXVWRAh7gJrYKzMkFKAVvVJgf2cL
PczyhRBUkUcsYL+s/VUVMTxGVXMu+lUmNafvzexSNtLZRXGKyxkCRhWQxDVVJi5hBo/w3rVomV+T
j4XkbP8t/jsoGEadlKobJVmt0q9xqAWd6vQbMgP4o/YLd5PQHSWvPB/jBluUIJ4tiTG+boF0sbc9
Z60F18QFuWeAklJBIB8+N5+bAnLnQM6arLBYSLCDecECAB/oOkhY4cUTuy5FbWp0DtKQHNCLwvnV
rhAIedONuCv4hyCXzkv8x/01ORBAqB/21gU7HxwBmw5PbvbcegaVBmnLdX9AiYzl4vnGg92WIYLt
UMVPOM5nE2UKSlIdUeMdMAufdz6tiPd5b5CJrIWcvPdX9/eZc0L1rv3ckKxp+7L0hAWGFgFOS9RN
REvsm1mfc/JY2UMPxXIt+C1FjN5QGvvlqUOoSuo7NtZoG67eYTNvnbNxjMvJt/ufVFGNlcqHYfeD
QHNeyHafQRkaIYiTBSVvBnzqu8kQNUXwf4GabB6l6DiOAqfROSGJPwTckmRyyumw4Ay40GmDUNeR
xvLVK+6h1qr0z6GKPraNKB9MUXiA9dTNWzbr3zB4S5mIL4JnyvLe9P16zk2NFtcBghbqKf6+m+IY
FwBQmlK21kZR7X99zN5nTX/HvRRBHErLg0xTwEvwzdOdecpR/HDCH8S7NNQPKlv8cuqtxp85JqlW
HXs8U9RyVzrwGEYT7UR61uTnHDIo9uk4GfIMnuaY1icej/K0o/3aarKTNzd7xPL04+8SC142Zp0U
YbenSB0AQKi+E7vuVnIHO6gLsqPhjEfm8cXwK2vG60liADsZW5xxONwWabUyaR1wggBltKg1aweA
e3LTYhc8xVr2ifat4h5hAXWb8/3AH+6/E4Oi8G8vOAam51GPD7kvwYHFuwvN8HA8MWeLPT9BqLIA
l8jTrvywXSpzYfKgrrzR3H0KkK+lfU+0vD4F9hM9P+oiV5BOOIYAALm7W41A7fTfCty8LMAIFTA/
HNdIrZaqHGT3qOxMtiKb9PLi8QfUtpVDx1K3pSROPybD1aqgtfnIntG9l5fuUzGkA9yWz+8dLMfc
Z7NN29CP353rt8EkJ3eb8oQG4znkW4az461+IuUa1UyuxY9PITvKTTGo6atrVKFWrssGuyQokj9/
cD6Z2vPrS6/X2yOgpYJDPhwMopeBa6ofl37sW066AuzW15n/0/TSd1m4YPbYGEw3RHCHWh3cBUqT
xXDOYKt9gGthpsH2kbSIFBd6/qPfan+oKLTyHFkupRkLWp1AFw17nExIjWxUqwkbGd+stcs4c8Rq
y+d3YKktYYuOas51KolECQv+7HBsK6zEGvoCjgKOSeUKr+Z/98HoEo57sTiNYs+ZCp8vFrSXTxxj
4ytJPkhMUnhWIn5u3nRfen363uf0EzxMXjtTDyZoBMZkbWhnRs615p/0CJ+AWUo8tjW+Dkj2RMbC
bWPHBZmmDa/54M9+y/CrAKW8P5rKSUTF1DvWmcXQg1jkwJb+6kQC3hWzgjU6txOXE5AoCc6FsYFH
WcxMca3wOs+OkD6TQuAUhq2wMxYyNZfUKthdeIJbRGw2PAH5iy2I+RiUXrvJwCRii8ajdCuVott8
qtbnB7xNlkNeRPHD7UpBaY6LXWyd2pSunpZce5pDAAJ9No6QMZZvre6CQcRwPslFcNxVq7RtEhN1
nrlyUEab68XWFShdnsPCiVixeDX0A61/sGiLacaOMVGTN9Ey5bceCDKUphICHqIJrWi48PigUv69
IFMf2dgLj2bEpPSjIRAvNP3u7uYmYf3qDLu6ef9QvnNbF4SdCOP1MB7CymdMhigJqQZqBcl8JGp2
QrC5uMjqUlCc7YjCLbJq6pz2Rk+UYyHkw52aoUhSeMa5pnpxJFWaiD3ZFFbwQT8n3FKjTIHvfqSB
ECtd2Vg2bN70K+WUvNaPW7eto7sqmABP780RWs38x+TAGunQoeRJRvI6KOPYOix2z1/NkExYW7KB
yROhgFwzu+buWe0ZlmtuZtwvsAcLhPg6jJnzkAF2UpR8ODeaSIlsbip98ZWVVqV4q6Q96MyhcRKN
c/MJt9dGJabgFOmepMT+S+dgxNjwvRIC9GP8KbWulS1VD4qeM3GVrp1VC+lDNjePpz7tz2nwryUY
9VwIHElp1KYFxLxofpgO22rFN2/x+xtGnbCFu2IdZWBqKvVdn/lGMw3JeAJSyQgxu1iUg7VWWYC1
J9r90Xzd/hogCpXOxR+DjKA0d/5FMfTYNltVQKcFbVPDSU2ks0kaccndbvDbv/a4IuF7uVyIrvKw
SFN2gGB7SRFXwd2HnxFaG3ZsjcBA/SwawvL0FUQ55HhnUuIxsZW5xdFv14Yp5EfpWvSsUMaOAmmu
5fyUD9fgWmnFGIuBSxnOKz4CRchNfsW8dE/wcSrqu86bkZ5JUhytQUTDZSdMfYfBtvzf0YNovBD5
LKBws0nnsVe5RrA2+4WJePrpieVgdLCUCD59tSoe/nZj9SAk/fy1zohXQaDhuy2AeGaBTATHnH72
98b9oHAgd5LJmpG3/vB43EmpjxHYAee5pZc/Qsory2EOe/hLpCN3p+02lX8QmW43/cOZFqojVHaS
Q8YNhlUzjZKroUgsoDi9Y0HfHNz9ZZ8sD8kH6+Mfnf5VzS3sp85M20OGZda6knkcaiXb9bOmmqsi
u9C+/gmx3USXNnZ1aRFztfAr1EDJ7WWIbwQm33iwQ9sqggzREgUCcOs6/gPTrKMH8N7xTcd0fCtO
nReb9ZPfKTr5RfNxV+VRg3m1Ho8qZtaIwq3EPHYfyuW9PH8qouQk1VT4THeoQv3M810O+xcMRANu
zEZdnIyMTBEIpuQXb7IMp2/8Y0zFv7ARa4Mknl8jjhlfc2J1Cd/womitgmBPT8NiW2XkjtTSy3tO
zh1yrXzQiAPZ8tMhel5txyRnwdzMTqSCj6JreBrklnx87hn8qBRAv4MhMShEh1Ar9gK1UtKRivgt
Rij2ISErHsKzK3fqtFRpf29udjvteVVPlqIoDfA1BnhDWtDHATLiGlwI9b3tPlm1Dj1548YRsBGc
+OIjZs1xFwZ6ZKFhuR12VFON+akHVEBWyK1UMan7IVZ3Fho5e+lCk5jDNkjRLagQMOSQQk+FpqGz
hWYhxjsAZ6wS9EPiui/4cHTdCTQO7ITGNmGfE/xdf7a/qf9UGZHUKPxCPUevR23JScz3ydxHGKg8
KWi9/J9yVOs1eG5XUTYlgMpyjXBtsts7p7g+QiPUZQnd/me5f5hksRAT3GXs2F9pGRGGLEgyauEP
4tLrjbFuh3zMQIF1eWnx9WP6jJuFWGMgeRoYjwn9y6W5G7DQ2DDGEpAwsjCSsVQnAP5F2BbURIkW
IpbA/p2L+wJDTpKvEfOFYybvhhHfHwfDWsNKgrde2hw2W3CMHId7tKJhx+rsjGr2VXe3UXJXNfmw
T/p5SY7T3b+GUAG75WZVr1A125apf1/xseNdXERmCdhc6sEqZygqPRjF2fLbJuu9YCkFb0FzhgBe
QlvBiS/ewwgIWGf8B09jUeIQKg/YFa93NzuCbSVJgL7xHtqlRb/fXYrjFK+B+CYR4+PkGUrVMQtZ
eFp/0LcWlrtwQtrJOTgFxBrAUcbcAmKFyqdv1YddJK0Sk/edp0aaiCMzCLea9lcW+irfzl3xUt/7
X6rhVWgEp/HwpNJ9VGMeEY0FzggYhUQ20bQhYQ2a5U/AJjFyZdzvztRCm74XR7sG5V/PzYLSY9g7
UBO8eg4xE+UxcSv0GhGW+kgatQuSu0tRkqH04z5CCq4UQZf09KIaXEOMXq+vecFd1pnIUERLIcGg
7XAHl2qVL9R08UGpEI4yZQjd9MgsiwT3j6ECNMhzbbvR+51DS5A6e0mPjgCp7ePmysz2+qYY+uKP
yVVcu/8nmDub6eJ51pxCskjvF6CZ8gajIPVVu5Mo+ZcRPl9HB9Sgnuyg/vTB5DoAzLzX+D2jbFWR
g0LAQwsMnA4L9BuEzy4cP/Ikhe4j0mPLca8ZiL6mCaPqMnW/uHlN5GkK+rIurFZ1yCYWxdaobVP5
rC9aqZW2iVXZCezFKeIp+dfW5oKwW4nwQTLlExDJCKSEtptnoRfbEdR6bjAYfnyxLD0qhglT4NM3
zQYiMnVT1Ujz5jeSBLz3JzqDGodvZ/km350in0SuATkAJMu0scpFCsvaOSZ0VTl7NS1fBISQqzCH
2nH2WqjBsS/0xczRIciZvtcmiPJUyLRP+YLuZi/li821phR80jknLvGthp+1w4Is8VvtWYoADd22
+v9G5rNY+or696hQdJxW/9xqpRXUojxOo3csWVKhtLiZFT5+sHGIztt0u61IhSg5nQ+hE77tOl6t
8yIYe8PKFp4FQxPJSZmIJwBo5CnEbsK3zGF88w18weV2h6XU+OvQnRRbwaQFlAhnviQQtm8nk55j
pMjs1a6g4IlVG46f6JuPb4mD1jGBBTLMYwRXOizw2hJycw7y512IPFQ5bIDvr85s3oVX27Ce1Zl5
PF/A56G9rrSqKxT5x/QKs3G7tnXPChSa5eWLCE6m6ohlfjjjBX+AE+ci2GRID4b1H1c6IWU8DnTm
/4hfh+2PJJt/HLDbYSpigB2ZRrwjLApwjSQsjo6ejZpOHGlLmfYr5VpMSnsRxfVrxtPbxGYzdbao
JWdnzNe10qTbPN2rkEM0qypKRpEScwSTFL2JrSXkMcSaY2EVDtzPlds3UWz6QkrV/oRUqbjbi/Oa
6PGJPOKQ7Nn3yI4u6Ot54hCeOTCakYu/CWpgn5m2AvcSwL+Cv7fIUhreBSvcjImJjQPlIJ+p/9eb
X+gGVuq9ZglpHrSj1wJ6cIgqfZLvIZM97ox3bbJMxza7OUxIgDC/dR8I5ogDc/BBK1bBckTCx0vM
jN9sBpAc1kpaL+NGS89OpLK9cPG7a+LrYPnr9v9YHC+CPahO4WhwgbA2rvDLfiIn6fG8+gv9hwsd
KaAaaVUX4tLKx6YzOhLL5wsP9d3GTKzmTRwhQbScshxGCHrCUEOjFWCUOLEGbeRcqVAhbQC6OV1U
zvE9uzQDi5vgzMZ2S0SS3J026lLwMdYcE9Oz8DEiI3mUTktQt7y96FI7vu7pd6fSkCVXYyAMZdCm
pe2u+7IFcIT0Kiyw2++CTzi5Jt3Fn48v39RdEwOQSX59+KN1NtNSRcO6twuagQ7vp4Z14oBLDLqD
oLmrpmTC6P4XDgHQOUikKt/EqilYyDiq3pUC7ilXxioIH9WamRDzaokzApxOHD1JLnctCrHnc0au
xesfHXYvxbocs8inJtMCtMgv7MGkGYktsoZCg1vWcLQ4I0r801QN/jx9Ohic5j1kugmMfEx9LgaR
YoBboCVcywVVeGlzT1NljV9ojhuXbs4XTyOPzMAFzWbXn2fYmiLCFQeV3MKHcD9G2No3+9UHCko3
L3GsXxWylUkvw1c0Earfph04TXg0pJKK/AZYmddbY/zjvrCILWwz62sj+UGP45xIJD6YXfTfrvbx
0Or0lEBOQXRr8G6Lpl5MbJ6t5rf7nZX4Qh4eLQ4eoh8PCal7cx4RPBqNtX0WFD81GMMIvm79qJX1
SlX0230n+/5y4sIpXwLyZbN1dg/MQducwfTlcOrdQkTTUY/keUlF+ZhbpTWeIx0U5t5aiZG9P1bP
fVqNSw87bLrTh9AKzYm+3dsh1nnrvp+9ChaVOJ+a5rQyA2kE37ytPE6/IFvHkgc6onMM7z8vdcKv
TcySNXrRiSjK6/CpGMMRjhI9K61b8pg/PxV10xro2kyKB7+AzTDnzt0VoWBtB3QzO0ur20/P+cuJ
eyjOsR8zD2vxTmaZnO3XL42v97z/Yo58O3s2TCqNzPuwGr/qZmlkhgXgcXaGCuR9ap1PnQWiFNvg
a/Q/YbrcRkGOPa46qRAkN6aibSEpwUcHmjGLfCawfpFBTthcZSGNROQViudc8e6rm9PBmpcyiwxi
2ODVSqdoKAtJ4dR5jWVOEfcIj2BCcwz87NAmx1XjmciPYOL0juze2J3UDZif9fAXRdbWBnUyCSfW
G8JC3X++Jjf+AteX41PXj56SOGzRw56kxy0G6FQZrdX2v8iq1H8V5+PU3TAB/CBmdYUte5ULk6oz
VlBDdi7D4RuDvd3b4y744+6YooxDGewChk3jDliOe+X2ckE69qycRDjElRdCLUs8ek5YVTVnqCvR
wRVV+Mnqmz5RWGfBhtmF3jkYNpFOrLyIb7/6FhDQytxw9nQPJmEDqEW3gg9++Nk0MTzsJo4b7/JP
+O4tlfWHNUWItW5p2OIQRTPywCIIlNsZ8DnzikDi3jhdE6T6/Lc/KtNgFkGWVW83ssykKSG4HIpe
DrSVSmoawhgMNw+gsDtFW8I0E1yUTu7ziEMe+BvceVFip7iR641/wgrHgkJvgPZPTxlb3ByMf3P9
0YoGT68S0rXNjxueqjcPiP2xMaa2jfabhRzBd66c2Novyi7LEGrGMv9oEw26wy4B4BUmHwrK5gIc
Vnys4lcENxvsxpYWknAmXn0XkbLFp80rQL4nw0QGX1zfCVz4CYfX30exytAwFhDq4G8xQpYfkeZF
xBPhyJyIJUqlKLHPlaAGLNOqT+CBHPWq9YhnAEkmEnozh0GlPCJWrGBLKbfd8z/UrYdaWLzl2BkP
8Oco9kRB5wQYmwTqM4g4tEsz67g0CY2DLsGG+szH/CtS3Vd3iHtKOhvG9nf9ea3GCBVgvPLQ31QQ
GsIhi7HmEgFGQ3LvxzCVzGwxOLpo2sY5W8AfSw8mau6IDV+WyqRF1kYLfdGiJMWyZhmhAM8wsjvC
YVcdVeP4YjlBR7JMByGSQ8+2ibwrxwqBX8s1Emf+s730FRig0y04HoH3ZvE0EYVDBqDRxo5sM0Jj
FoyBQP2+O/WGog9OXpxshzq9zNvC5VGlaEEtkKYYbgRhiYf+d93yChVnF8SG+VEafKf9HioMv9pD
1NXQYlL0s3xzU1lcFb1THKswr8HNhT7O/ryfsmM3EOXlloZC/QKUY9RE0bxJfVNOlObmK280rBXP
WyKxwMSmtF7ec4QJsHPAmHl19YPIarwFzfVee8EvWW61xzFZ18GB3ZDq4DieDdGxlp6YspNyo8Yo
UL/HQ4gtKyiZB/8f8b4MYcfwFYIq+RCAo5yEllAtL3VE9butaP+6UsNIVFxRZrtO3n1ilaRFF+gt
JmjegvYHNnCzu7oeqfDC67e6I0DeLv37KLDIKsozMOpe7r+vxm/tNWuIO3h8vSJVmaHsQd9sj1xv
tp3f+tx8bEWz0imSAsmCKld0jOf6nP5BbeonkivV2R6qbsJ8wtdCeENbwFlxR2mcb84hodsGo742
/4RZYdpTO02jHXzxc4TUYsXZhid0AL5IolLjjK49z2m50yXRsWgNHEv2N+fnHb92hngLinvOBXPw
p6R/O/Rip/YquG6OK023guscPLvDNZcUPM2saVi2ZXjbGAlvWZWcCs2Udf5enlQPdbENcOI34HnD
FICCe2eynMZsPljd+gwM7cSzatgm83jJtLPUNId3CgaGsjlW8OsjMvV1H6YrZai13cGZ5XoCTxNv
8yzWLEDZ8LLrvmL4SL7kdgnhDoPRXq++f3ALudIXeN2gnqPBquN2Zm52iPSUZUzo6tncP6bboqI6
smBTbkqvNQKQssZ8Fdu4zirOcakyuHJAcYvh7cujD+Zvt20WhMOcj5HEnm5n3vwySNalmYWAUdFR
p/kb/CjZTS2m5A+pg28qixpUGdPsSk93BRSlkXSj+y1f/NcM+9QNEJ0gPAP0AZ1f9hgLnWOC+r5t
t2ibstWczauxASpDlaZKmZ0UyKgIPljKl3HX7x+GygHH/v9P6QYyIocruU+vMPe4peAU8OZN7lSv
670Zhx1LyrROk8tjv+ySWka13qaNL0E2PtKFRFqb+CXBFNkmxpGCID5bviIA6EHd2XLXsFBOYzic
DVOanWDa41PsjDc7MnoeF8vW4NbeEt69IAQKUS6kEa/XOs4OXLsDkDQQ5IPk6ow4D8M07rMLcXFc
Jm0W27mJGDZ+oF0i/wITXAEWhyDgTAmQO+Ej1rSdr3qljYiCxp6sILAzOC58KJdpviXI4N/vi8IZ
9tJPX4WieMtoCMsXRg8kO4MFKemcsrxpuudOlaqS3wQ9UY6mvtMes0WID836L6hjzbCv20aI8XpY
/fdlYcIVwvNYkpH78cXgGxFpEauF1NQ8/HBfTH91sM7t6FnH0XwPk4fNse2+dXVTTjqXwYC4Ynmi
eAW1Ghs0SwZsvNBv2AVX7y1yDmdBfD0FOztsf6wIC7Frg20D9FbHd8k/KJoa8Sd7hCUc933Fs/Xv
Brr5kdb7RH6Gz1u94xgMEBYJggpTw7fCZkqbWUzZ9Kvf8bbTjmbsNP4zJ5Gv9OXxZiMDOotQISO3
hJwWPY7xBpNPEJIIACufEH61av/lCjCL25aXLmS3gtIxODqgGcTlnXBpxlCH/0I39T8aIHMWgAOf
1Jz9PohUcVXIIuK1FMC4Lm1ATq9VIuURo6DJw0xAZejPWjOVtceVFOjgbF3O8JXB3RR+F/7r4DuM
RovG3w1NxYdPoyFClV3tAvqE4ezMZJPaXgmnwr3cHJ1E36WSZE+gmtO6rkJP+U+LARbaOKsP7RYV
LFXG2H3J/78P4OIzasJYMBijoBD64mktITFvJ2izCW1q3NKbZw6m7bctNZtrjv9RdMPvgrye0Ndi
TsBf3yt2lIJn/S8+t/abaON1WVXkN9exImV4MVWTKLlRbs9RKaKaUxzpMSd4SlTIuSQql/DHuAJg
b9kr8Ju/myDQlHKm/1mv6nO57ErROaKZkrEle4y9GJyBE3vxF3Hz4axS3HuVB8ayuMCJxGqW27hq
J6ugAGrpN1lgru0d9GcI+t6G5Tqz0+AB7rV1qNZZNycNNQIiWvy02S6RXmdsmiQu073AFo74m3JH
10600yAcWSc+0HKCKx/8XZebDp56irfaacwo+0NGEBaFpAbs/YLR26wIpUkPeqnOsWVTStKcUDTO
0ZMGzYdi5KV2OTAMa3fYKNcoBzD2jFvbdg2KrzsLquB582qF1F1TnFkv2QkuWhUdAQBgxwzfbAWo
RD1eBcHCitpzepl0IVpuo6EEZoGlgHZnuZrTa3Zo+5OdTJAIXHbucp3WZNS4Vktb7pULpVtXIkCv
6PPgOtxYG1O68mo6XDySYOKY49WuuuCg0nww0KEBPw62VWTH6cM1faT1yzHMJqbUDBf8BQglhvor
Yl95btzHXZF7tQaMHvqPribCk+1pxPie1aR9YX93Bh60HwgCeVYUawGd15TNl8GUPNmDl/L8Vc08
57Aia3Oarm+i7XOZCOzU12neuKMlK7lY4J7ArM2NEk+yaTs4PUPwSP8tvrdrKHd8+xGqMp87JEWK
vEFBoO0V/9t6Ei8sdBeARf79JL9GA+UNBokGXy+11c3iV2C5I8lvuMO6GXk1xpTPcxYcWAWbdbOh
GHzAg8LY4iMq4yYKL/2MUaMET/1ik9K+AaqhWW6KXZdCEkNVAriKVuHFiwOj69m5urKDZbU3I90i
CLoJH7hZXbQzBCUJ9wQgbBFnKqYRyae5w17+47AZwSipuR4YJipG7D93H5KZQYfp/Wu70F83hmLe
Luz32MrcmqYFkGqj/BpmRR1NN3nFZU5TY/5vSkp2HlG5oB5lTlHtP/t+AGg2yN9wpe3G6+M7y6fy
P2F2fYevxsfpCSwbkTykRic8m62v82FuxXuKhBqes2H/T8D6iq5VDfnzQYsVJWvNh7z/LmoZG3it
5BWhfC7gvimEIMNaidcl5K/sTipRhoPleogfRg0SmoezDLLHrE1npqmZCPGA8/G/ALi9JLYnrR6S
xUQiD7Apg/IrlwjsLnakTkPnrVjWAMi9JA4Ht2y5uXbd/ETtcgvbXv47WG7MJ8Q4NpVH2rdBnP0Y
tZbpCZRUujazkx7FPLo40LRnL705/c7Yv1ep0xtCG7zPyCDD5GPZ6Yd4L8godElHcaT/bHQ1SiE6
dJVyh8PsEVPjxsz1x2HoXtwBFh44q+4ZD1wFJtpArperCuvTQkUcECrGDF6QrElvIZJr57Gx0cf0
gvvbA+fxAknJu3Th+/jRfWQtF3Mn/NzLlrjs6VlaBOubf0srWNVpH+1HPI3dXgFrNfEjtqX/ibWi
oq7cEBeGcuhdyFYHIOE/Fa65BWDrcJutl4hDLBzw0V4nAssq8TFe9j+dWHnZG2P610iyHR6MZYe9
RJ+IGLzM8l/dxws5wSL2KP6fUsHmmBkQWklHOU1aBxTFH+jQRP24wyxHO1DfvGrGLwNtaZwu01Ol
16E+7j9hjUTeLT4hR1RL6AE62iC1RbzUw3ifeN0tcMCrOWzXATFunzi6uu7xkUOkQ47AJNVmSi3x
MVyXxP3mDcot5wvmXq2qzoHbkQJ4ulC/5Cn638bkmGA7OQarBRrEJIcoQxS+rlGZl7rRvzydujSy
Y1YzmbN2bhwBdkM7zmpCyUf1hgV6RaoWKeE2fU5M3uTqFwNxNa1SldbMWHUzcqEiFjJ8ScpbfWTP
P4WXtJVAiY1LBQzu0pX0ctXc7EsI05wCYXePl4WDGlSmFncweGEO8NFTreTD/TDTU4BOys0lqk56
XD5g3UYB2aiRuS7BcPZiYXiBfqMRbaIS/Hrv9fwovhQWsq76Qyq0KvtcwPCPpiwSp14PEVwkYs2S
pmL2W20XTbfUFXwmfXFqJmMpJs5ZMU2e5m10Cc+j6NKv9eY5XZzU1B4VQbggvgplf2RjgKujhSR0
nt0HgsCNLBSmOQ9+8YnML3IISjZAWERX95+eJSmOGM3vqAr/VFBoa6PX3NQDNzD568N+kQC/Kbhp
QOJAzzUhPTdYXkdcgTvaXUx4oINrydE6i5yCOevvctx/qzZVAspGR2aA5zPepojnW1uRR/CDkKP2
8ZVaWpNYryM12gacfi3y9EyDG8+m1IlT8nbHdDeUVSVViau/3wnUe4bG+v8gcvIOijEBqKfTnM/p
hbWDSSKzslWVmEtBQPRhwHrbbCezrk7RF139RpammOPqyIU2eHvIBOpcQ43VKC4rjcs6AwIICOyB
3k4XlCOMFKQYPfSJOCySfqCHrcindE3QzLGnqT+WJO2axX57h/RthdwUinFVpqqgFIV+/yT4DeEd
WQ+6345v5SbUYf/zTLAgzRvI1jivW4g/ZsEj4t32anHBJJJPnce9y3cv33aeNyIgHCYq5sOUhTn5
BLkXj5WvbsRDkZvKnPX219KQFifk46ZRizxJc2IuXQZJvm99eqFAYqI13+PK+If+jjvAl9sDkxKl
yn6mZSrT7EWRTA02vpZ9PtrL16sbHp/kED/FBk16dLbNb7IhoeuGg9VNm9k2K3o0GX8SQ/8JB4Bq
oXtWKckz02EM37UnsluprigZgsnnPi94Uzq8qEKdUn96ChcQcTV5kJVi1XcSrcvLa+lzqA4TpDtg
Uydygdpttb8lKaVKevhXS5IPhw64Q5fwynmowqJev/fSR9mxYHP2tj+RlpyrQnEtpVv6/dv7rLfc
kjP+cMvlmka+li+hjaV/TX8FVl3atlc5YAkGNRXCrTQhqsYNMqeYNTnmCUj4g7zLIbN6uYuVZwG4
XbwFlbTCvqKgPVXmHo2bHB8nwRSAVe8xkrJywZe7hdg77B2CbPVpTcpL0g4v7BTm7uE/c7+bY3wO
FLG1rvUVKhFzYAVHvOKTTGBpVO2GP219aXTEg5sT8FGf3/coHs6bUTvFR/6iGJvXc/54lgb/jmKh
XhDkyQhotgjEJ4f3VYAFwhQLTw3+BOe9cEW/XhrMzH90o8i6c6Umtv2PdQrDAMQwFvTAaLdrKYmd
TLgftTezSekvXHJCenxWsW5s9tAaGVqSPYXUmTHwFmcNJMrQ55v0gMmnVw6AcRJcZGmmPFZEuBng
gba9WIpYEsfupT3JwNV/B+slJJixIimR/C40WxTkMjQEo/pwtZU5z98cjuslBjBHoZpk8g0Yc2o3
twujnB1H0FE0U8WmRwpeQOtgFTs5d4VKkCbHGBA60CUzOHOIrq4hHzICwxazB6bygHXzOwuncchZ
lfwcAkD2O9rXoOwyw5KrGIoaoVZIeQoNSU+t9Zi9yvXQPj0JTxx3ijrH46ep8VX8Yavjy+TMK+wn
kLBt1n175xpmhMK8qUSCKltVdAXi6NZl1mazyLKAX+6qZ7EG500pLSecnJIWzdKKaTJROF84qFE9
MMeonpqGd418VYAF1A62o07iVQlliitSUzAjcwKiS8dUuiGAyhZ8Cf0p/nt18crgxlMs/lyBJt0V
W0dqh3MHA1cxf+CMtPmi4oELkmrm81sX2NKQJp9W7/69He4EiHh6PgKgvM9OW13iEuLts6VhVmYo
L5FBe0EDuaT4Q/4NnpJMZcgQaLSwuxXTCSmk2hIjMT03iRkDof8xwn+crJAxNYQB5WPsDb5QXHAl
LDYXk9O8AIr9lzxAJNazdNI7gQc0PKvHGOt/JrtQ4bVZMaktHuLlqM9mps/4/D5Zzu9roUtl+304
4AYU3tqbPCQJzR9DUr5kjvw35HkqtOQy+Eg5+Hsl8BPyasmjk27jcEmXJUNfb6RwRfTrCSXzIQSe
B9lgpV+abM4h88Pgjv0aR187W7Y1wL7kWn7seXqV/ZGbRFYtFqI9voszA4KP2MoWi48Rl6Gzrz+H
7gIIQpBfqXyjgckD/h5tE+3kw8qCkNxzGOaWOXsKfcA4BDnsaawab+5RbMTz690+iYtSi6KoxDQK
+k+iAeP5Y58LtYma41GJ+zs6EWj2tB9s6haZWCqLIaB/NVDm14N8GgBVg22s8unlTfl/8qdS4pPc
E/2QfOYy5WP7D7ezOG2EpBaT4tesbTVJ/dc5g3RO01pB/CcjZ7oazo0yvZhtLYE7UOeBws9oC0ya
okiB4HKUtjnRGEoLUvdTl+/c4PdN1lRrYLlWj0iNEkkQ6Vup5bDfYyzv4OV2rjd2oWOGBBOCDR/K
EmLxZfTzCHrcwTH7VB3KULaF8WIuKDjRm1cmn8yl0MOFdipi/6RDoww4DT4uVJHRXCnl429/W6VT
Q+dwCDO6cjdeeAzJNkevGVKu+tv6ZLo/+OSgvP9MltGqVuiwDxqdH+Fi9vTqC+QTZTpTUtnx3poI
B5ItqoRQYzvcpzipMvCt/b+W224rj+KyXwP80J/j+KKvnMTP47NfQi0DvW02+agFgGa1Wj3VY5w4
zbAj0vaCZGd2vb8gW91RgIvzQFHBPEkidU+dj2ux5w94EmQle1hOQkW5Ts3op6pjq2x6yaSz9vxR
HOVWWlP0ZXYADRG9CoA+fC6NBy0NJEeOtnmhQerzOhUv0fFH53RitiUp2gE+j2rtwNVQKsj18F3n
g+sQb718XhSm6HKtFAgV8fodn/AR94ZiggpVZcSs41tVDISRAmWv9Q5ax6eQPX6dRAkcBXnnCxeL
nAVA3WzloeeNOZa24kcrUNnzTvI1XwgVM4gXLVYvV+cb80CA3oky5uQDgQEgbDCF/RrmWILgXyfC
JstGFCKvHVrdsdZmZYOE4N8ksXX3e/SZwtY6apm+SV0670c/6sQkDOzM7Rliz7/ZE4UPwaVZU3nG
adeNvsUUVHzKuOc6NzhLQrTWylykdyEq0VAaBHU+FRWyoKgdWQdN1BFZKQKspzGvWVhJ9rStEac6
WKSvb/MVXqO90cmt5z8iAhMVSxyOlVE2kEtPUXPHVuhwdUa3yuSkXc9AGmCuHBX7dHMzZjeekXYL
j4cDRHAenfEy4lSwXu7i6qI0h7GkzNLvxEcWRs6+9AOlJniwio4HRcbE8mk0isqm82aUsQ4Wkh+r
3Ykj4uxA8B0kdo8Qi2TCUtgWkIue6PWZrO3B23TuOhJXsIDhzRs/H5UHFQI0oVZ+VMZXJ6f3hD8N
+fPvjHa1Y6G3bt8t9wi7LFQukEBTN6iRRSBc9X6mrPEw+BEpSYfRaeTEmkJy44zX32n3oGhRuifz
frcMr2NV49BPGTIjEGWYp2fiMgEXMbp75ldXPcPbY9zqa4Xs8mtMby2bGijJU+Gzkp2tkwb358Sk
Budj5NeNThZ4hWaiyr3gI3WigMNzPvsOa9+Ug+cbHQuoh7rMCmOXpEKi7oFVLk1Fx5ytizZKxSu7
EI4dxq5girxQxAZiZD6P4eaN+Xmvoq0OkhVLQJYu02tzDZ481wfsHyy9tmAmLu2+Rt8SnQZL3dqh
AcbVxD3PB71yKvAW/fg71stpzsZ+uf6Cc3An8mvJWOCdhraReeVrKcXp58HTbe6enC41GMbAMOPM
BDtzJMUdQx4VfsmXu1GJ8vAAiiALxAVDHs/8thgoyBNa/G49tlLu1G6HrynYZJhzhTklhp2dH85q
Lb4gEXS8obdb7f5hFcm4Sobclpbi/yalq0gmVZP1g1/IguSsNtbwksMtR2Y3MmbKpg9C9sBLIKDi
Q+5Z6+zDdfkbM8HgnRSbD/QvpMpPJ3kMgRPjHLFlVZaV9VMFf8FjFBGIlO1poxrftWgh0Nw2YSuo
575PIaldp7O5frUw0Yvorqt/9IUI6A7F6v+LYf4E8uPAMIz8kCWr2jK/9LZlifcwzGi4e5/QtPo1
/U+XfVgcjO0iIkQwZMrjjNj1kbkljiDFJJRzKQ+qMIiVsc8bnKIJKBT2vBy7ZhPXL+B43IDPMe/U
DWB/n81lzpwJlLMaFbNHSMPWZ4tZ63DtAtoLut5liXb4X6AnmGkoqkijkSvOMV85yfwRoInqdIRk
8Mh65IrUf6jI5nYcDa4hlpuUvZYw8zzkCyhC8R8bKPHUu8IX2Zsnv5BxBnTe/ajSB1yvBthCTh65
7jjotzIpp+2j3b1UHYjd3c30UvpHpXUk40SetrPFESMvR7CZmPnkfVUT3UELPzcHzuImop4+NqUl
/dNA/DlNDku3MDUy6jyiOSse+/lzcDTYcorUrVpoJhsvv4eB9j4FDTsRM3Ivdlasc3G958/DnSYg
NDT0HyYKhf+fuLv/9jMatIyP4GUEn0yxx2BlZkPnlfQ/7LvRAYq/bq/dKufSbyzs8F93A3tnHMF4
wfC39aKmp9bkBVg+JR6acEcTm1ZeTKLdofcO0+AiCCQSeHgpeuAYJqh0V9pcfXZlKpjmWkyUWthy
bTJAXPQXv4GYZrEcKxx4nL64viofeRtCPj0WBrjT8SUNOo0hnN+3avB9NhkzSU3wOql0DcqCGuWI
Vpb12VIbdZ86Tlx8xzrpYqrrQKKdDhYXqJl9ER3zu/arHEDTnrKVJxfX5axOUp/BeA+T1/ULCf2C
0wNKts5jTEEWV7qPokT2WtZ1YLZ2nciXkiekfUO4DKa3UfOpGd4p/gZWHjgKr9oLx9pID8V1sXy4
/W6K772YGk4mg+LnCdGOEwfn3QeY20JRLn91bxQq/0oHYgSrGa3KuqeLbIfPuFASJAceeoTqLXd+
yXdtgvbAcWv/SAlqZ+O08zyY6617Po2ch/ItrGIzISU62d+3NYy1eSgM9t41O8KdBXLjIw2W6UPJ
ussv2ug2uNF7ONP/P1gjk4uZ/xD+vHoRLex7l8PSN8A2hnIJjpmAVCDSNOpjFBabdeBk+hpeIdQO
n/cZxdASCwkW9WDdsCBKs4nWMFuOqDG+O+Roct0NBVmuoelzOFp39y0qqBM4Y7nF1oLQcO52Ludi
ccKE05yxOzeI3pIA5eOWXL/fYOAhjMx8rSzuSoDhnWueOT/ArzwfdvQgLIW+WeqwYD4ixh0TkASy
Fw6JrH+rbcsR7S7XQdyhTyB3oSAMmpqbOsycyY7txVBvfzyjFZobNCaowPiCNbZp22NyUpHIQlf0
3Y6YKH8JAke7rFbDCEDvsOSb7CBwXAp/pSxarwXa3avKuY/nbeoOclI2eQPNaPWok0o+FxDDmbXt
QuBPj1FVKujVfeW1FnUSwhMwzgvtYWjs8ViSSQZZb/92wy6coAkdQ4KCywCAZ9ZflqPhzbsaUgv8
gKQ/i4q1hwfATRzMqllvq1zNkFO1AKZK/4ZLw/tHK1YW64Kwhbg7nprmV96ANJxhmokGf3B9zA7w
O4UQroqmxh8JzqfvAEnif3XQrqatIcX4BiDTasDCkgi2T1jpcHPxS8r72+A3T0T85p3s+kulUp67
kW8gMjASneXX42QH4rk79fCyBMfz9gszvkTMzxafESVc/UbCMnXOHb8YjC9EPy0+ntLW39KquyhI
wkaK6nhyTE1EPaDn9oBPUiRBj5V6kJEBCCfnQ919FSP3XI1r1jnvJKs0T/IWm37RSkwg3ERvcgTf
sMdWtEJeptGpgYmbYRwvKjE4JnJHEDERAfV4v5tUTrC4n73qmCyCxhn/KP3pROH08ucA0cShiKPj
mepaXdeYkBP6RDjLvAqQCSYBkp4e+TXhhDBxH3+Ww8XGhXjhPkRGlgyuAlf/db75zMI4WbVk2yeJ
Xkqmn5NBlTe1LgJxUZGTEV49L6RQx8JZrdU3pPKZifjRvBHcfkL9hY6jYybbcrr3EV9G6tVeRehS
LNDoKHbnKZ8nuU2F3/yLmXrCLlvsx9ZJA3K4Bm5XbXe80YiCQOETKojkUzvQU7BgUHiqW04BMrmd
AKFCtr6cR/jJqmX5GBtyhotNsfV/7kEVlWWgdeVKWw5V9liNoWh6MUFErAgChZvZE08HS+ulYyBK
vq1FIgJfx0JjELZO909KOelqdjo/bqt08YUxYyBc94R+NsuoqlfAboyH/rEMLOg72NSuxIwycsm/
4cUd1txvljavVhpUph4hKXcmKYpvGk6Sw9AjSZESbr3R4DoSjWB7gwsKED6M4FXTEh7DCHW54S31
L/zfsOoLFXRl+WwPD3B73MHXGSbBVLl21IYUgdtUmS3iBOlyM4T73grK7FyV826BO0BUhv0NDAZg
0vNMjNaXVgahjlMgB4kerjyDzlkrIiLKy6c97uNizQp/DH4gDHBYr2X6gwrqzI5cIFNlpWVgt5Z5
cHNLeqo7gC19vMqYtxanjjFo3yQ1SLDisjU4+eX+C5tj8p5gXAXi8u/HmHfGdVExy7z6ju9ZolGV
soBrG11Fy8vZWvWRTXUD+ivGqyAGpDadYGvKiVoQuE17nC/X+4YCPXa/An9ls0i0zcr8pVxB96oW
fUmLotyD2r0OrOzcqNhpvE80qWMYGA0SNEO+hLvNsBN6Py+TlYyGTFVMh+P8xbcI3dNpVbTMxMgT
HYfgkKapXECpDDPQRQYJFYgvkrtQ2Wtk94/0O4oF6XxXb7Lj6sXyHRqUWOzrHP4TmSnbgjiAVZ6F
rXjF7BCdHEp65LvMutVGODJHAhj+xBOCgXo2ShxZDSCIeIRSB5BHGeWi5ZN7xAuejvhs5lc8T8BJ
VEfzDKGXooAvaCLV7KRTsGZR7YDeKeDEnd93o2Vzo0oiZmYJg2KxI60uKBuUnODqmmXZWVtjUKfj
CNoIOvciXLpAwDACFCDnm4cUeZp4RpgoUkRJ21P9bWoqraX6V2YdCDK7HXlYb8H4jnkPUKRd/Lrp
V7N1Z20I2TvRWg26VFvmZEN1TF96CPCtOb8QXGzPCIDMECKSe3YrRkwflgc4IHEyGnFSDnvlHOVY
2n3L4CwJ6ro/QmMtdf6m3Yy5GjemC8cE9Cf9oUHq+cljuYwsAtOwlkXjPcM0ko5hBad9Pc0u9uzf
HB6+jCLLNsBs+bfcS6cb0KtbcIAV3B1u3xl7zeBhU0shoLb8wMoRQcCUYucvy5V8xtTzEL/NsPDr
gVrKiQwHCuZQ7/auaSj6Lb86Rl/J9UgDEPFIPalwXo1WuWtR/1pDcsOfjL36fT7dakw9wBxkaZrm
3uOf2O9xS+Fgd7NWQ6nD/MKcEmbxl5+kEj8ArBVXypfZ1MjOYNzZT1cRB+CM/MCOGXsQp6RhY0cz
Nu8k3xmc9TH7+swqJ5Mz2drVnTrJLJDLp3XAgncr8H1crf+rb+20XDQ05X1DFKYM/U3LvzHxfzNh
HMl/+km1FrHx8onBseVjT5JcMyLSc4KEafb7fywCUOMj2UtIVoXCBqcvc6MQqQ5V6du2TnVHEDDO
PgoPqD7N7JYXQ+96vBl9TDj1j47e1xEc6nwDEPfikleifNEyy8/MFxfKQeFLCN3PptjsJLbeGDA5
LXsqQPVWAV2vJsquUWZOSd1zPz71Vwqbe0B6cn2FUVIp/8RLOEDjXczoRjGfpN48fcbaCYIoEfby
u4UA7ZnOR+R5a3eeHOzo1jDWEb9Z3ahOLa6C6rgq2HSXEZG/vZ/VTGatYDw+6TQ+ZhGKTiQ86ZXk
qc6jcuWwbEkNO94kGl0/OMk+192p5PHTWHkuZhUimIuZdyj8dLrnXsiVTxnZYmgJjB8E6dD2DVrE
r+VtiNo5R81mCWmKWh1W31x1P2/lJeByt8rWGILZyOiHxRhOcB/Fs5dKVpJIs9fCFcuhefIfkSZJ
j8mk9buXuqkBz4BgFlIR/nK6hhdT7KpSh40BLfYADQ8iyYRNfwjanLL9JzOH73gfekjChMV0yI6K
5uFC0Ta5A7sQUvxhOs1dQJYx1KW28sEzsDHmTBAncNR8yGMuM7avxuR3LClwWAd6bPb0BRu2wA0q
crW/6EwitrlY/zj0AAEBzqumVu1y8CaWRuvDXttLB/lt3vN9TvYJyyOiVCn0oIPYgtT8kTHrbLTo
bGavgZoTFoJ1Fmm1u8DHfTKxnCaeQt7UjSSyo9tBKhufaN1UQ/SARR3hARviK+rzS7cP+d+CbS4J
lcslby8X/QJeHUboaZb8nCBBapNsKPyvAoVBY3/oNXu05cE8q74NYbjrSzh6ar6jyedwwYYbbM2v
VHKibasPtiELlvPzQToAIeYoIw1lvYKXkmUCvBvJtvC+K5vw11JqQbrFefJIfLjTeBsDjSM5+9Tu
kD5Hy5z2OmKGAzo/md0Y2wBO6jFfdC3eEHG7X2MJj7BhYF0y1m4d6mR4Zye839ivSXqwDBa7/zas
jni/laiaEQHUKzMM6tBZ/dGdULo+PzvYevzin18X8rWH37rBLBemeJb1BCpMyubed+stuNxoyaGt
O8UwlEyiaY7LTuYWipk6mw7x0CJ3gv8SfePP8QHhTAekixyxKQnLHrEivH1xjXYCHWg0kN2SMa8l
AMWk4R/wzuMO4WkLFz/sQt2ZVFMHTPDstAnf4Y23WEOFyLfungzlTqFAfmR9pBDHTMDWyUgb9KT8
WdZTz2iqzMsdPDotzO3vlZntwHDeAiEKxKp9D3fOUDGbKFWnCiH7609D7rlkjS/CldZqIi6I5a8G
ZYujcatPd5keU1MsI/jBxTvl1NiYsmKTDLHILm5PomIpdrJF3JKrzOAB9IIsJ80K0mwKWo90XELY
FxwEnnULc/nSzJKdTUIgmUNanVC2kKCn+65Shq/2vlLboimts88PWSUwRuSzbOujgeOEGvKNk/OB
X73L6daSs3D/TFXRt9pRpy5tZC324uZwKHjWNbNxbcakqMukboxHakm11x5P+in8mtoWBOo3Ty+i
7Purs3qpv7522ifjQFXNuysVdMnCHgPwge9FkXkSAZ/Vb8DbLmejf6WIoUbjfYxMPJ/U/CTZMRlU
QvYc8UQV+JHXxr76Ab0fRd0abgoM68HEdomoKEEr4/uyb6j7ZRbhw/JgZMpuNWzvO2YjF4W//hMi
jpNWJpHqVjFuOQJ36UjBl9U8lMXOyGjwhcdR4fU+90JBlw9oMK/WziA0O3iQg8X8R4vtiWMsfvHz
8Sd8DNcqelaZUsA/1gLJoXNHI0LlPlHJF5LdjGeSrVpzx6hVs8d/RnZHymy3prxIP8x0CMwa5qF2
RdFBcULZmdXro1Qq/LVZgxu1Lh5ftzP0XJQYgUrb1RPCX7ZKt5lKPjgtACo8m9gn7pCBkDrktLuJ
p8yVW4Xm7LJEXyKB3UNH3SJ7HyXtH+xQnuTlD/sKmjamV6eVOV1eDMYEdrLzM7WkI6qhsG0YrDuZ
XktaMYm4amGU7rIHXdeDMkPA8T7pIVQFPpc5X4BGt6AKZ7hHXy8eC2dF4pkzVRdOJPXUPVHb1myc
qNlh3T2xTyWJbpzdEaSUcVQluYfIU/JunZpXblxYDNjhGvL7e70nmemFo48p8ISqWu71B/P7n7sv
FWz70FFM9LNSuKodccNXzHimRwuQtpOoQ5Ek+AhLnTbxa+9VTCtDJd7+rXe/sxF8ZuUFKj5yP54/
6LMKBB83tQBd5rlZrYvmdOlnXjudo2GX0g7E0PSVD0jTilOOONDk3MVuc62gyZ1SUBMcEMcBVWLk
z2hlRHF3tf8DkZYx9qcuSwoU8OBCDFFju1VbACEZuoWlVX92lUsJPj/FW9iEvGMsGHKIdTb2T4Yk
l9ywaXtsPkmIbTm/flUfV017eWO9BWQUTH4bHVR0ClElxA4Z4CJ/0ae4Ty5eSpI6JQHl7mJOm1EZ
32brlouaW6khzTm0LjVSbaU6aUq1jH48yksKzWTbiifQAasxqStXDNTT1DLFzRYHxQIKfAbkggyp
KVcLx8Q8eXyNOaos4xsxQ4jMOPOwaaK9h59LW6qguxD7Rhay0v6145No5LEvaJHxmZB0qe3+66Tj
cgVzCafeqJafAA0R2138/fZq/3AVatEEZwaSzcHTM5UF7n+jO83aLXNaYCIrzaAe+gP0DbDwdGr/
9g3PIb0Mt96gYiMnrL12/JDXmncFdHAD5q4rxoRtwIiCth/AWoc9zYGnbAuA7reoJ7PkaBubcDlN
Pgct5wm2pFQzhOwB+UeOkN7z3T4R2hxDeYXnhkBTuHd5Z5p8HqK7LF1GhJlRs1oZggGsstZzvDOS
Sd2ZzJTVooI6HJtug72KJ7Q2iPgFLLRPbxNSpX7oWMCiwHqHy8wlW+l9De41Ifyqd65qVs3Co5VK
F1PgRaXQ+gT3UvVzfSgDYeOjCt4pHcNV8Sdqk/gcVy7wtkcbSb/LzRr/ukaAfeEU5Yb/il+TBSVi
bc/wlbdotny1r7G/EUeJdT0IwGckVuODWq+0YjYMRJBsqhjwJs5V0Huxevasu6UtGNHhNfaNGOhP
4/yDv4n194mbpyvRzsKIDvDldkU5XeCEg9MDIXbHJJuHoKuvpGbDz3dSGG54pHJxhzQA5GvFnxoj
wp5oWeGlJnfU+gBmwKlYh6VBdxJ4y7e5+P+xnVeP2xTdiKlEyL/s/6dCUU1rtEidlQl0uKlNBBLB
uTI62vWEntrimRixuSEqtk7tDFt6iVu1HJ1IXoyDQgc+TJ9RK9sSXDaU3jzFUid1ngdXITQb88Mb
nVRHQ5Gb2ta1nkZVGEeERLANz5hQzN+SgS85DYp5F3qULe3byBa401/e20RzDKiyIRKhwbqvTAIr
Eg4AzMcSL3Gtf2HVKRtzSfck+icWMpr0sAZO5iYam5hS243xAN+OQaQbjsDI4U6OFoYZnx3OoHZt
xVmIBQCvCHC66dFqUj80lnPi5seh5nr41AYF07JEsHKgfga1I8ICpPsc/ONwUcTcdaELk49k79HJ
fEzugwwJBMmsFnPkV5p5IZXGtmmq3/Q8VqYSbXNcPHTmcPaOoLEzeKaTZogU98/0OV1ATT3qCRd2
K2XRkH2XNSj4ph4z+ETsovL5MPTP7+DabDt5elX1eASafz1pajHY+7YG4IlMSRC4bEzbB6AdWdDg
tw2GxcUqIyIapLP32n5ZSGG7GrCt58OX4R5dUgoXTittDPfd//2Lb/Ur4KrNZiPD01hWm20x8o4Q
67288vfe4Ey7Oqe86ns/bIhFIV41LVKc5XkjL1ljyqUtKwg6YdTPRbtRnGrb0A76fYCjsyQxIvES
pQol785n61mHeeo9dGS0SvR5JtaWqDmvTlrflXaJtAOSBAhwvf/29ENuhivZR0gUJ+1vZ38W8+2j
buq3y9ODG43XZydah1TDvMmQeflwRcnqLfRyG5IhEp3wksQJjf4UON3ooznlqC/pOLFaeKCNo6yE
ekzYma4NMTn3x0HII4S4utAHHw+51BlOviV8hjrOXKDF60r1+o5d7YC4gIb4z87O3WXoLTB9dKPp
yCIxI0W+kpNpfuZBhvMRb3YaeJy20OFav1YpB5r4awuo6B3BO/abg9JNJkWcbIH4PRG/qjNQRjZM
du8GHjW7xCR4h5anXEKQiMsFauT75dkjEI705oB1KZZkJGLfCEn5Po34EnWHPOyKO1DmzZYuysO1
Ii+5eJnaUVI428K7E0BDTxjqX9tja0CuDx6K2OtE+SDy0hVJdbU24wNEYu6XBrZSvf4q0/Mmli4o
z+5mLsncDI+Zb/R1/CPZ2jm4c92+d/ADdjMYF85FwsLpJ58MonHPRlCSB5BiRnVtMtieoj5fXLdz
L0fK4S5ymXxqhMk3To2oyYQUEf4FaN79v750VJ03fAC9g6d3k+kSrW3975d3YtLYyN42QNniyVRs
/+eSgHNp6jj4JZlibn58Dbh/LqMOEirEGY6EpSWCMYDOzBqblyjxaygqvqYBwTv+GDw7zuI9rWmb
T62owHypaysvZ02LoMPqyaKsvbV+jjeW2DhevdD/IXtxZrcrr3OD3edhoMUAz5R9lS7PJdmwoABv
oC1PD0S7cEvIegUmX/1z7JjpmbzHCBFzmaK7jX0L5prZ3do1A5fGtx3rhu99nbTWiePJMIbSqzKL
eXtR9iX7u2wdm8DGvH+2iWsFI/pV5Bz7rLlHRk8jxeXkq6wjKf4gx6MRDgDFPFlqbllBYP/BanBr
nKyaD4oZrYTcvfWxVC6my+S+/imOGzJwIGJz2Jmyw4uHHDGj6+u7D+z5nPorZnIvUNJdzM0liDvK
p5ymvkyYotIPIJp2gU+vD8RVI60s3IZx2pjuk4aaxu6N6PrsBViDLcPAaF5ydHKiTW26X13IjrCZ
1hUVRQeb3TJJJDZPat3EZz8A0FNAsxgOZUaLUR08ptImK7Cr85WMUkKkX/8WbUcMrKTNCqhxGxHF
pD8jAMiMaJag+s/ksAOxNIVNsetUbU0eJcUyVksUmp4JnbA4xVwzXyXD1KZzIO1GVpEUtLT1gnnv
q0RWPGFWQy2JrXsN2bjHsSRZN/fokIdP4jzZHtaoFvGlyXvZb8vds7iRV+zPW5T223Hf/oznYwKM
xHz2y7NJxUjAKmpd0H2XdRf75JhZGAJnXyyYLa88P6GoDe9BVSAXLQ79uCAIVRhbFyOKlJGpnQYn
+RR18l/GT8fZwf8KZMuvdVBOf2eq1pPLzuiJWkz6oQh6bJhxLQkGDKqQb7dhIiI610pqtzdJvIuP
2WM3UVry2nxgwWDdD6pTm9+ZttXanSwa3qn34nHjA0TxQl4P7PtqjsHo4cmiEh3hC7MkNov5q+OB
6GQBU6TEqlqclkB8EfDy/jAYTWCZ3UPl1Qpghq1sWShrDMG+5Uf2XKuR8bMiz6m5AFN7ulsRe3PD
zq5LK5exuYrFEiyOxt1zyjeo6LHzFscBsHyph6IxPUB+nN184Ud5+UvY31clDzZb1VIf9hgNMSRj
1pqfcIB2zjPOW92S0wSqSagDiqtBKdsEqN88NJyXgFoFNWNSELvCeAEHygIlJmB9sI0SEOwd86CJ
Sv0uKqZjLRtYadNcDWSY6gehDW8vkTjunlHcnbMxRQsaJjO8MqhoNde3c8EsQX/W2otOduhM07zs
SKkQkkQzeoNVcHCLlrYR2PZ3fALopK9dv+IcFiKn0K4pUk2lB0Wqt685QUTl/JxjyFSw06T+35rv
WgWFFLT+7P7L17lxGyTgFtUkiwDErm1oZYzoYAWewRhEM7VkMRmYGe+dMZf/Ixg6pKoNkW75d9st
VlLKD9zCux4dzOrAaX7WwWY0NXsSr1rxeXjwOmS0QeDZJwbd3Glqdp4MtNTJ7XmkV5VYKqT37RfU
jy3QMYrcRRFyU5OBOC27N82xIacE8xmmK2yfxz2bH9P5/LFPmdTG9edLucSoAX+Y3C5cGZiuXkvj
1V95xuJCTAwxF5VJVgCVUgsFQof7RJ9XajoymlnEFIaqmMLdnwnqwf63qnw1fHOP1wJq4jX3I5D3
DAP30DKUP/CAuvvFRglDWfXS42mA8W6luv1rDDi2U8ccfq0okSRNjUHb91rfoOodCwK21mpO/DZN
VDo/qEUUydW6BAuJTcSI8ETPU46njjWRJl1PlLy+IucFdpsLeaELfTwTFnViVJkIpwXZolXuTIWr
b7/G5sHLB8mbQMow4mZoFa2z4n5p2gI1kpyOKFLanm8yt7nZbHY7eDbG1f4oB/CxeLBAT29GiJ1X
uBDlRMIMRJhYYEqgbLE6DwPatSlC6LlLT/d7SXbiUruVBiYtYg9jvkaC+gg/jgtO+fiZSjhJh28I
GXM8WPqJNl4Kh/EQLo/eCyMNccilCMA9dnv2OF1zMcGwlPUKYYmNeIeMz82fUQEjoHP/MhvMmjdw
VZogr6pvsFQrowLeo4zifuUoSsTvXCeLB8mu4GfBjgD604Fw8EYnw7SgBKb3kjy9ewHBtlEYHnQ4
Xdh+HJcOjTj3yVqOtt/OaCJKo65QQ8unwa+v5snqqhaPg+Wh58ZxdGjHU1xxehfdg9svWPsnX6Wb
7CC88GI3UMg05o/5zetEzudkSYmEYiVCKEqqzG0/4n1xJ+zuR6kJXLBisSBjJE82PAq0+2ocPpab
yfPRKMZRsSWOBT6xe0h8Ne9HG7YrsNDWQ0kwTzKeo/cLVnfJhTYrzq50AShT1JYpet+3zdfjVAvj
97DRUkbbAlQLYEz7xrPmySinsB0OcZTYbYTC6QTtHmMIjftg1VozE4KNXoQd1WuhiHrm19zP02eb
xEL6+wnb1J2LBGEQCPAu7P4n+Z6ZuplbyKak1d2ea0xoxseHzKTo9cb3vPh5fZSqK+f84Jdb3R1L
6OQry/9ynHrqfuRaBtkysFhEjkeISzLemtTtShNFn4XL35cKgwFyuN7AcTlQ28KvR6DtASAwWZse
RPHrir/kPVPX+MhnF3Q2/JvypQ+t7y2L9Tfig/V4Z1aXw7Q2sZzj/c1srHA406pqLsFQByMsZgRq
ELyKjtvlTxJ/1QOk9PhQBIp/4edLmgPeR2oGzB39xDu+my57OzbnRin4psk/Gtp63QEal+eZFoZM
JPxtlnOGIF+qmlVTg18UlUrjKr/kfOJoQ1YG5hZfsfUHNTxzwyNfBBJt9Tmr24R6Ky6Odmlj0dOh
ULsksVf1PcnYWClGxC4fXA7lr/ygjBvxBFW4miIP9YWo9ekndEfbG9CcSJ1LzXFsdcLmo727DWFM
3c4TBYJyZfE4nPDokgX1l9ZhHzLUfeeCAdGQNbtPL+9ei8idN0Nq3stFJuN6oAOSbs5fh2fzf2+T
mLaTK6bM7n8/CsBVNrFoUbAIEzVCjhR7eFWntNFz32RoFC3+EUEMx+y0h42oNjqkWIM9bcOYlVf2
MszALFOlkBuWEVbuVRfMGG4ItzXDQAFxxS+IZy+CYxZzsmtAV1SA3IiXXh0igJAO1KQZtZlyEgrn
bZg7LEMjNuS75XQpP6v6412zDdEwPt5A1L4mbXKYqNNru2oEHj2DxOoSBNQQKdOhgDZu6da1B/98
PhoObN+n351ZMBmAP1GXTmzf7RgRzHWRRuiPuhiZqdrcMQYgNNffHqF7mC1aktl8PxaVr98X+RJY
fOJq2lMjP4Cb8IBhIgI0Dt1k2dCIxGLFECOMMmdRCX2WBLMonZs69LqgQ0o/6FjErWCr4cEGqnt9
vkGFhpYSktIx1oZY3x3W1dZ/QPHwq0Zo3Nity17Ry/364bhepH3rkK0Aa9m6UTg6CcrqU3iDEYgO
O77cljWZy40ZLB91ii7jyV4y/2scpcvrAUoD3Ml8rjWHWArs+Ab/gdnwFDaX+hR8QR96BZBSUZX6
lfvUbHayYnC0kwaRL8lOSVfSw3U+qMy32JUh9O6J3YL9odTj4OHcAKGuPXTUmO9BcO9CLzqKRfom
djn4ZgOm3wSlz6LdBw1I6yOmU1QaU7Hq5SYx/cyTded39RyVdrGB4OvFUOxEUwI2mhetuG1sI3vc
dW4Zt8yIuiBbUW9vh8Tu+dgw7Y7lrf2JmWnMENVrwMC8WGZfolSTGTFQj2gisfgtC73l/fofTaUh
1unUi9o/ReM3E89Jw9QtyHBGWcQ7GKmCcEJP3TjhwJFxxL9i8vtyCD4GPsbfXcKUNG8kqu8ax4G1
xIwi6k7HkSuT7G6h1l03HCiyBtfn3+dXs1fZ00JDN59sxGyWKxnFSk9swzPBMyR3milro3Mo9BK3
7hHMGLHj136kALottbEy9mLhaKMqRULpuepgqOrPJHV4oeWB40oYUeTB8GeX7WFFJR3vr98yj5vI
mVZQepFTKGEO3HgXPGHn35Ve+bX3NWsVkfT9y4Q53DuIsrsKz5un8khmeT3MaIQ+HSnAqlRsZBT7
WYmf6Ufotfu9POuWIdSfzgy5dOoiqBiT5glI/lIqU5AqbU3fauhCc5TwB750bCJ2+bO19FLqHtxE
P7R4oAs8foCszDpLs5zs7QjNWC2BBToDmBbY8xREErGwcJ34pxUMvSG0v80xuJqiznIUh+V6yop+
5nibitTsEWiMRcZcbOFV2TcfO5/Tu8nso0HJB5/AYEUlrc4eEOAqtrbPA+8qagBv6buBOtnUqHme
wtEOzHRGik4r0UdbL6CcPEk7L4tkkB3zc+t2JTocFD3exhOe7ZzqpDuD1AbRwZ55p3MetLLRCyI4
F+Gm7IXen/Cg5xz00+jGBFyRGLCGFFhGePdSaUhde9dhNCTU2KHdNwR3FZAFA6u/tcd1QK0/8/IG
8kLNbidSLjENTtefFViQKF6JdhkFG6UR59BkP2Uap9r7dgZg9qNbBQZAZgahVQmZBLU9fq0Lw/tL
8iOkD5EmFLg7I2xCjCMb/mmQ2Y+Cu62pvqvVtRCLYzfzVvV8YsLUqwt8uXk+KqMspzGGC/Mw9vW1
rCJIyNSxWgoL3hSs/W0ofzIRs3CZIoCdkZSfzzWd+SCKEuKTVvtgMLbyFHYzUAzIjZZ43giu13Gk
AXj72D4uDknYr2ZojAZBBsYSCRE99GfkIOE0Yyn+vbPQS6bbSzfkiF3zAZetV4VyVPa/ESc8iYz2
GnXgaFyO2rCYae6gz1sSgwcWo32dEOxkZtuCqgagTxCkHYfHsOJD3M4MFacFmJMUv3NLb0+MGCX8
RLeb7lTnX1HUkuSfPJsdvtazWlnMjYYgFROAQ1fLTkv8mpS+Ny8xrSsYUymrXGATWpRTS0qlWeAB
XkkB47EXGrHrQ4fhNjmjOqrRnqQnMnawgvMWyq8D1QPJXKGk3JcUn3pEGyCyeMB/qIEa7/gIxtzs
GB9zVOgLUYh9nQhp1Z2mvDzoE0/uPCvFYefBWxNJpNT9XHO92D3MMhfc9I8fkeg/m17nQReMIWWH
/KVs5BjvXLUv9szZcGqFE6vTzXNrBapU7KMv2eHK6+zLABOp+LkABafup+kS1imoBjoNI/HKKJmC
KYw7pW5dZ2FWAkoUkW3sSP0HAkea6A1aOERJ6punj6R0WSQvpdbPhrc1ZT/Kej8lrPyg+TnQhhNF
DLdQyPRJXb6HFen5yoJIHtR1TPd9mm+M4dsMODxF+scdK8+EhmTVurNqxbldaTr5E5uDEMNpuzj6
y0f+nbSmjm3cY6cGAcM/m43fYuCBjiGj3jO/kwRfg91BHF/t3LFFMmryyXm11hpo2mwHDZ7sUeQ0
k+bVoiL1alvdzCfUnNzH1l2wd7u8KdtUuwZtEX7Mzl6WbGOURBO4EYHhOIIiPOAqCcDH1iogDvM3
qmQZKSPfLc4iD7hVBKONsN6r3UdrNEa6UlUF2k+osXpNjFES1L1ME7gmnM1D7iG9Yp9Ne3BSu+G2
op4NMlDyzHWOnoas4Efu5Gc5i/oLjrGUj757jTqIQSAoB7NnCxPqdfXNvLe3mOz2+kFaEHAl1/Ys
+Wiut1KQ6D6XPTq0Ruj85FFYBfTuqBE2vKFFRmbz8kCgORaIxVK6nwGvx0EBLF89nL64mof2FVvu
JXLobjhnyOrlvcxlGEaSzpZLdUcSRRiavJQfLSeM7nz3WNHBxXSDlTAYsgYMxPSvmGoMDh4WYPXe
75Vd0cCw+4oukfkVBk99UR4Umfbz31KC4zN+z1ILkJWFqKSlqdFnpMXry1b7X2S/9Ei6TZEXgGUs
jah2MeE/v7Ot8Pu4oVKFaUzQoBPjq1T+JOK5V3ZwlPBS8Yk8tTsd0rucKkb9WjUCJp9lHKthPSho
d4ZabG1yiL+37uQ3/RouCdKcPss/MyaL8s+hh4bcaOKh8mSMdKQi18o/jIX2z4kgaBCUwdoHdchk
jFm9W3PlMU1Xa73/34HFMTvsSys4wmCGMYeSUp5ZrJg1o4T7Sf2GP2XrXrmNjvrnJNgk7K1Y0Fsw
7sJXMts5HmgJ3k+WQjJr+UnV3lF/VThYi637A6YMCQ5zTHUyRLwNgqw3tMkoRQRt2BMEs4gNEtlX
cJSJ391cZWdmW/AYnsgcn5DSOBveA/L8fAgpJYeVKfkkiKgi5irqTJVo0Mz9UYJlA7Xz1tfTpWnO
JbYHn8/HR2hgwkPeb6VHq2mf8B2uj/a9r6bHp0uL6F4hkLG0CpXxfLlNFe+xGxggolnrRzBh0Os8
YA8EcrVNlx8LKlC8DT6KQmyClEhCSXI/3CGWV1RZVrEXaAzGaWmqBqA7QjnBDya632cRLFz4nv6Q
bQiJBWCyESPZxkvWzlb8z79nfABuEatf5Eqkpt9pTC1k8ssO+I1of5UHn6txLtxgGkrw2qAcRmG+
qVqwXJ9KIrSmCWXwmGPCb0oPzQmE3+eX9qkiUBdMqfbUmlSNaOhlSwyrreUtXlmz5POGVvXHsQlw
CADH2F0rans1Kko9/CND1a80Wnnf89u5ADfQzpbuU41mTVHdBff3QhSdQLJ/heWvdpgDJ0tKbrjN
KwSETnN70LlqVXFhpkXn3lrYl16VPPuq13VlGxUUcrYarD4D4rjAVEMAwn80YSmSj4jYHmYCqIAC
88NdDdMpAkCf3le6E1hNJKIgyglGP4WOfCGWu3z6hKs+3L4tPE+JiQ73QgMdYy89zMEzVh6d0HAV
CxeEyC9s2TluEFCSLdscJxDhfuh3IxgD+5VDOJIpo+juHAjwCYwicMmCkAtOtVY+9WaVgHO5fwhR
EXByGVeo7B1lT6guT9n+J0Dhkz6YZNAdcvFWPN8qoSuGuwJ4aUEL9PMZYOBZEAT98ZLYW0xdC6I4
/B55kc/n6J5LVwPnCUQBycNru2iJe05xkfeH1emuVPQ7UoTtShJ3duF00qDqVMUCUsnsNC7LGKBg
0vGEGnUavy9qHgWBKGXtqq7vFFxEBmkyv2TqilJ7JMZvg+JRaAw6WpCpDjawL0y32WfSCYGdpIvQ
uvGzWd+T1MWZedYikK0rGyrn1E0A3N4UPqXNz5WRq3pObP1l45oSNk+w8C8Iy4h016JV514pbraY
sOuUAUjygEg5h4I6ihru9gB3jQVNIRjZeD8HruZOaVXbnnr582ENUgpAxBiRv4JWJsMw2fHNrDwK
uobQ3k0uyFqZulTYxD5KB8W9BnrIjZJZMKprnCHXaeFTg7WzDA5T87IAeNIAkZUsXthgCAQxowlN
s8OAqmD7HngXkZp8tRfFLt/3nhTOGQtwWLVzTwyyNk8i9u6D4f2Z728ZJUzWROeRg8lborrJCR79
w90S+52nQseTteBiZObGonAoirJL9fgVcGRtF7xtLSsH+wat8k2LvttrfES/fyqra5JLEqmzXXVB
MZOsHj5IRN8Umd6GRXU2OB7Qxmn4Sd3VekXL1mrLYj+qpPSi/u3OJasN3/jrcSr1SIIdjEEYoB4E
1wNguiNDpjKHsJWkm8pkIyAZpkh/XDG/3HHfaAeRaSUFD96OIzT2U6LQA3+rO5nJUEF7cwWnQXYa
6iPoR4SDdtu1MbLbzZcwG2tMyEWgRgENS4cVKFgE5y9+zgKonAIK1/3QmTAKqs/ztmu+PTmYAfmm
3qvdoOA2tpeJ/6yRENrajg8BLKw2v39jmIr1ZWET+0ARUK8+HN4VvzblJuyQMzQNL3E19MYif622
XIEMrTNg7ye/f8AZiV223zKA9LpnuGkKQDCpyZutcRGco8uJMEnHZcoFF9dUn5LiglTF1Q83Tust
EescbqFnNSX7NyE9xT5N6h8SZhJZQHx2wWjQyM3Gmo/Y2y4gqCt0A+CWgwc+8WRaNRA1kOblGt4h
1MHBsMoVtoNYyr/AYob1vhRz+RYUhJdrbRuzysPiMERFxVVzXlJs5Z9Gy4KXF+TmSGT6A/jfwUSo
B5R7PcKfgBVu5w8hfmuD6iQ45lHAZSuYmK7FOZzs49av61QPovxXrA2NGyC5no6v9Ce3UZLe887u
Ep2JW60VkTxVd9Dqg3KblY04JGrDSsVWsjL3WXKaWSLIoqdEr5nATsMqqoj3aTOc7Zx61+XdMhC6
3PmN91sh7L2Qi2wpaMshX0lBKf8aUcUOx4WIDDYQQIUj76/C4Jo+KWzRfGkFMWduOwWR+JFrK6Bj
aZFqSENki25j6GbKjAa7g9I57avGoLqtUSdAG6UBisd4F2Gp2Hz96ifhproFdjSqbuMtvHdtSbc+
qVoKibeA/WLB/DwdvtHLsxwJkSvfTtK6ikHlAIOYKRZxE5cyuX2qK5xk0QgeWybVd63Wfzj+wpBE
nw7h/x0A4sT/bH0bdkMn07HQoSxKW6TBd4E2BCzGG709bFL8lZU/CsCWHrOdJq09DbTw79ngX2FY
5yN8imsvOpAb8YqoLJWW9y96cSahX/2nadvx829twCdVoRxNcXqME7rdKNmYVkQKxNyZ1Z6PVyka
QaHnEw80923HyrA26i/eeRmhmo7Pj+HsovHbHzIAtfG2RV/75oImtVSuwXpts810hvMnE3XkkkLI
G0+/aEAROzg2MOyRcLd3tY9QKiNjy7t84FVzTkrm/eVQ2HRCykB/04jjM9dkiP0K27Wspf2tYqZl
Qf7LHMO2CkHPc+z0QENZzOVUXgwFZTW7sYTaKoD/ks6EuVus7t6WjOUnQLFjNVJU4RG21Ga4QeFq
3hcHrI9pGyQ0nP9tqpu7ytnxKyx0h+CFYl438gmZLwBrfYzjFEfwG6UaKNkik3iFEUzEhsmGrGWE
83J9tftA2SnEmgTu43iQt1m/cDz/HdyFDegaaWFcGhQFHtwC+gxCo0fdLNhcgc+1CODt66UNKiqg
8iqiZ1LhnJrn8n29ZoMQsYiZJ8xrFWTQ7j5D0dSUGQpF9eDQOQkzkeRA23nymB6i6PXmAn/xZBaP
ZBlzIU2jxkSXNTfIg4+oef7sxRutk4D7zsIcaM+xvSawbjr7vQ8NGb+G15CZxWa4pmKUtNms5Nd8
hVlto0iQkLiA/fJJT1ZIh4zEgBBwiUUw8iPbQaAds/J8AlXHsjkEvVZMSkiEDo5PSjprf3KjweDl
4Og0vwuuyNIWREn613zbJUjQ4QH6hl1SFWjM0ZVTlEW5ULMG9lZ7mVpMC1TZ8AodJ+Yd2o3GQHBD
qWUCGtvu201mWUGzXQlzxwnVaFLtLbTy1g8ZjOGDcV1/KgiyDcdZe7zfe0uuxPR1kI5duKz0+u3R
AZcknNLhYVhy/IIKwFUNv7MIwPJO+DRXXts5y62L3dflIM/mVz4g1KrKGIXaTtWgqWMRezf0xh8d
DijpSq/hsj8eIFaL9jwq3cnz+1xiABwpC3JbiUDD1O0bXtETULo7BuByxTGE8iRwSeZutvbIHuiR
b/y67Iu9HP66dKyM5wXONGiZkZvbLiBiB8kTCV5XRRm/uKA2KyDhdBdGPe6TiEbkgwMXbqhRXORW
h9GmK3ka0r7UqrxZR5ixIBZsxzCyRaJ5ux73WnliwiIrrP6JrVDiB0hPbAqcr1H5glVJVh28ech4
YPfymZrCsM9xQ+3xK4+za9PYFP6rSXxsuoowE/yXZIi7tlL2rHa+yJP9niSeACtmI5tRcbAEk8hb
howmBRDjr9Zb0oOtLazT3ZUhqx4dg7FCc3HzdRU5mKLHksNlZcZxLpzi6p0fYD+3W8orvldY/a+p
l5djsI8gdEIEhiCS3DRRYeRSgplDxnLDRLwp+J8rnkgjqa3LXPo0ytjMVL0Kh6cUXsNQ84KyexWk
zXxhkOY6H7cTfUXAjjjFLlsEVpHIh5Cvlrg36PHGyOELgQ0ljy3ufJ/Xc6Xpsgx+LsJ+aA4/BlAC
j626Z/kN98ezgfUfhOv1A/vTDGUmDRIrxyy+Zn8zBzxWkvmKVhrwL+2/4Q9pXD9bkFzMo8aKhDjk
vdwYHN4Aruzs3l1qgWOp42Jywp5dlwgbnh0h1D6tnpUYS1slhE+c4wZLlEa6/OzU3fHKKPERRsbi
K6Dkk95kPiD1vU75ik4rb+VuhunGI+Gawo9+HJg8HI6J8SkrQpsDxahNhlqayh19F+i979thK1fN
fIFYlZ872TtAb9fJgi4bWKjCeDAdwsNJEAJOVU4renjdj2gHsnwLupUhx1nSZgpIBE8NG1V3wrZt
knEfXdRWdKS2R60U/ffnjVggRR/TQ42uiCOZiHYJKkTjBgz+MYwk/dpWtPcJ2xA5f2P9ICvO37VN
rhQHPePXR9HnSSIWbILN5WAHtqiQb7pnOMtekW+B/jdUEP9+UVMOUuTXM5BiNUv02jYS4boakF8j
r+hnZFsJ1YBXc5XW6iNtcDGS5uk8odfjipGx49WSNYGNE0ps1Aml77ZFuQytxWHhnZj1clS2v+sA
nTC3VPIaKPaAZXjjRM9ueVnYY3Vee9EqtB+A3tWTmyt+GO+mK/SZ0FBlpPhLPfUnOZ57X3YaWLjh
Y95isuIPzH9TF2G3owopHZc17qObogelCC7uFQFUREBlc3+yoECM9tI++ADdkA5s6wKaqKvNliq0
GrTxgT7TnY0Jqcd6pEnNtseNJarsSaPU8QYzzZMVoFytbu0KT5B+CsBYW5u5sEVokPP/5FkJl/6W
/20OYSASifgeS4CGg8G91m0EH4X9Qdot+EU9po/Pri5fvZNl1dcmrftD5sNdIwEy6o2MRQVPvemd
6Kg4ijtfQDcagi8GuQdZYv5bM5f1UYLiCbUhP5W7XfEA00Lpk9zWBWtaCTdRQorHNgcqsWpg8hCf
SafT+8O+yHio0mnOXjQWicyRKPh0LLXSeP/WoA/lRL9kRmilRkSYkOEzkumgy8tvYmFkDAHOpdmK
iGCaEaYughc40neoFZ85dpb6yfEyn2Gyxymi4/kgVgYlZIs+Yaa/Wpo6BR/hkMiRp8l+oRZbkJBO
lllaCl7bVCBwTMMlCohaLZhK0Y9iDg752Av5KFWV3WJ7iLO8oC6OQ6INy12Rj5J5dRJAoQOCYT6B
KDEmFjpvGYlSTXze6F13NyKFMBT5FARdSnXZPyCfL/OiD6EJUY1dLYgIP3FMO3i1SpvUl+wU9XIC
eFDZyAEs9XMDv+JLYp3GYAKdnNMP50ug1VTrvza1r7iwbo+xFTRS7H7fj8zK943qjsIRAkedhlmx
iVdXZPvT14IZA8cSO2iYECAdnKMEOMMsrkLL6ulfzWasBJrE/S9OB0mp4geeDDRFNUiHcAhv/tr3
IoOiYij1tGgM8q0K+8mjwz/m/azTETSg2Rb7znWKJwVzOUdONfi8naZOkJyWTpJvPFWHUwVWijPt
a8VpLCjlFp25xQhuPRNDb4I0/OiI/ZriILwJRNJII5CzljquwWetUCnVtcv5Z8HAtJMGFWMnVh8G
7FlbKx1DDu7jO9Sj/5qjOA0TUxMlU/cbBYhk1KatafVB6xIuqz3Qj7U6SsHEBIk6EHRF6Ai1puNT
e9lYDyxSteKtNpVBrdmquceAFRskmY2mzsR/BV1UHCfrZxM//ZgnSxFSzWR6oe37AXCxFwmrAXif
lsw7MRX460DC5rQWbmzhTsHsOQhhnMOYSGjOOzGOzwMru8Jt0H0Zn7vvWidTmHu48+mB6whNKYPr
+nMX8ohMCY9+F3Ny2u+y1SkZZjqVBMnaGjg5FNXEcpFFVtoYcFZKFPhQ4EheMwEt3zHS9xUr/fm7
U+AqMzqrPw1NvZoqdavbdHyGO9QAF1rHwS1Z1rFhdWdArbBcGsViW+uqoQSO5pvYpxK1YgQh2lRx
XvFbECQYr80uA5sEt/z8Z7NQ7s+fixa2ZbYeLhwrlsZBr6I2ApNujBkrhrqmiS0IbOPxH7++w/8W
ShDctSNvx/XAwc9qWhWxh0q4qizf6NkgSupwJk8ejRrjs2gptpEtFNRugf07g+ypAWl4thaAiM1F
4RPpvprFd5cE1FYoWcEzwPw3NHUai3wpFF9S7WfMqP1uUKRB2BMYSHlO/AM4VdqJiGROH4z7x6sJ
pEFmnv/93G07RR9+/G5YSc1kleV1oWQMiInPdPHz2fddeLaL+kZFL6SZeMS3vFCrWoIrXQlCrviA
8rvBI/SsMahxM0MAaaUU2Z1dOz3kz6e0nPOAZ2niuBJf0mzidNOb/aazQ3lS8sluoOA3We/0GTUy
snkdLOLPTT+g9Gt5es67xRenNxCAeQi8o7OOWt+K3dHo/GbIgZMp0zXLjomw9ck41GAbACD6Lhz+
H46OGIeVn3YEpImwfWxYsrRfPWB+yJt6u6HtCP0bZ1t6/CPN3lTy0vKa3L4nMwUTkeDIzDKCiNpz
PpnFg2IcylFqepPFrAkWVgZUOhhXBvgs4ShXvpAePsvbQgb00OMknYyMFDtgLi6lVWyGHS0IgYOf
fkbAM+43UbSWo24bpM+dFsNbdyp+vHN14Pbf5EDENJ6TnXW7/X95IFeW7DKIvZVMzI5A3EdRuF7F
kTFkk+7CNaTEx6AlxUDYo7/SVsXMib2l7VfCVnLObAk3HQdwxNh5esGsIK5tA0zRfGGl8sBOPlLW
iP16xg7k60c+A7gEa0/YP9U/jWUD5/iL7W24/toC1JDwHvzjGZJFMv+ozdofEQYGaDFIxlHUxa8e
966jengHX7gnL4vpo7MJfps0HNv5ZMtpBEW5OaLauVABH3GMtBoQPK4EMav5EyO4UBuzBcnnINXE
O4D83Ssj7jFF7kvqzzJq8Gd4P5IxvYQeZUJffZ4fE46e1H7TXQ2h+0Mciuwq7lhN96jMZQXHf7Ap
LJat0Ikh1REegO7WqteiJK9OLXveIaXEO9AIys3aqYh3429qjzBXu4A5K4GImS+P+ndpP5ZjbQZA
MYkZYuZpFP81yKhbt1Jibbpy4klQZ6tc3cI+wiUWh9lKpNi3JuGai80QvS7ymcGP6Ku/N5cNSkYd
ES1rflFjvgjnzw9RP9GIvA6o6B0XjYTM1xEi9+WK1JFRCwBCpGyrFRRE7Ks+FX2mhQaamOZ3oh+y
L7/8t+PjR8EWIZFeVnckI5EvoBom+1XxXWn6FnU8kCyNmqvocxehpIaKWT5fw1QX13K+wC30cecD
YuzJMWLE76IXY3WM+CKv+dCW4ftihl8i3Yca7aAzjcugKXRdu3EJjlXxCvFsWKnUK4A3+T5J946o
nGqwE1nIN2DNflnENiVg5YpSBY6KJ2ToXnlHqshPPvuUztkCzRrgYXGy7Qun3sxvipQgekcBaavD
oxTl/Q50lK4zz1eyMPRn3grwH+hnGUz3wMn/53GASYwdK0lhbUH4u4waAjkfgGbQzMavIM0V6aEx
RegjcjyR5oEWx8jriygDREegk80rbOGtzeYaQIdmD34TK+OGZa+WUzZfUuxy2RQifQipkYql4lTg
MLj8bjgooo1k2ncnN0zOgY6+BCdizPzscv6MuwXK5TDSEMed76XTwLmhHhuH8kaA+7Ey+H9IpcLt
95w3PxauYHJf+M9a7mPfWUG9FNm/SZ94X1GaFPxxr4rwB+kAfa4ZTePCguuKd3BXFXugdCiEkWwZ
c3SGSx4tLQ7+XbPOwKuWyJuA576a8UpreNeTRC59r9CGdZoYHIOwj7SeLpG1nxnsT+UovZipXF1z
lLs+g7Xuiu5StBPKn8xWP7WRT4srXJmvYqtIgwtt2711oq1aCU2G9rApzO9p7gGCDf7GxZl9y5S6
S5+QG09GfGCU0oyX4uYczgTQzoFFL5OcwyPKNbKrmWCjn9H/5adhvEiAq0jxRS/oI6z6DN7vMg+N
pHE78O24jBDrrgMC+EN8oQvxvUsRquiViAaxUUsO2JXpFj+KUe/rgXqVjsYsVOQ17irnjGre67zK
OPT0lSmtViKfniynye+DPD1fYxoDZTTdgP2Lfo2TzCiE4edQ06b/mp2SWuUadQ7qLL0RhmnDSYxZ
/aIVg9vSZOcSgyGZ1MFgSaoqpSB+M799jI/yYZk8dpVPujAvoCokyW33y2kqYfV3Whl00mBwYI5n
t8cUjcEh5a23QingHalZ6xnwtzozRd6siHZXVJI9jSO8F73SXgSB7Q1f0861XabcnPnPL4P7opwq
Z7M3s2fv7eZrItPPP9XO+oPDlsnSmanoaWLRlPQmtAi4xucbVc5pcznxFcK+8EQM2TMNRtQ+AMG4
RrbeNizsIQIOUXHAo3mJ98jFW77QYARUYFYgqdA3/N+xJeihHMkBXBrLUBV9/AkUm2bsRA6tM4XD
JYoPC1WA9pEXmz2xJtTuCmkZBc3Lz1EMVH9MCDU3C0A5fk44ub9FKuKtkj5V1jikeD1FC4H+2xnT
Lv6Ek1SnvPQTVTAbNj1EcY7iyyyquow+IWF3pZQKULvgdGMEv3ub0i8kfdUD1HrFc662rD39IrL+
wVVPtMoV2Zp1KJ58TR8g9+UcSBQmnwoOFfkP4u2aIlpqbMEPCE8gosNTpe0Ip2ocbWXmhttnAwXB
/qSV4Xnjt66HvEDYs8hjeLXpE1ZtJRGncjgEzfi1FJfpxk+jPQEuvA72zo8yUrXz8FW4/BE92xsz
Feh5QH+xm7nrpF2z6nMXsyTpjOs9MG0Ehp7vCw3R/uuQqjiLDrYQN8jqSHJT5buk9GfXG4FzJtnK
+117ruoZMYYe8pJ8MgDTSSr3xDulO1wRV+NWx83enVVgzoQW5IDloj9tsKcP8fTAgtG3KbLdRwnf
GB3dkBJ839oFNot87aeIgWoFVGGF1fP+9YvPRlrEjnCMR7eq9xq3rR6nh2wyzX4oT8+xfbX3iWy+
eH37W115NOes3fgtF0tz6be/fTFvp0eWWXZYDtUlvaKK9fSp8PNZg/bAajrEsLRrfBZfBwj8ZUDo
A+cNp1KwQ6g7dcjtd9gk315Pvyb6xYTNlXpczwyf0Q9Fw4h7ZsBnHW3NeGwsU8Jzt/KMAMebRRjG
KS69pvVCVd6iIQ2Z2kX/ID9DRykurE78iVE+gsQGk9XVvtjz6ZDNTLem2d6rejd/6F/2nJDbxkJy
504aIAOprxL2cv8HfoW4q1BKh1P+bqXcnIF6EsxObd7Zb8nSRIrgaTqa+c5lAbp4dlHaIQYdWqir
2xiIDgoF0v3NCPes7mvol0areOoXBclOD5YmbNGDhWcdk9NAivxCnEc0u68xX5xuq1+xMvDG8ZC+
4fjANgExdV3Ti6dBFSwm0q6f01f2LYktPqwXbS7O9IzV2CB4TmNKFpMTqlTwFuQWZfQQcW+1iPPx
5qcKxowcDbImDpzEQX4YxuE4NkZjkTmRj9rWHeHg3ZpvcbXFX98+NviwwLsG3QnyYr9WIG/pOuUr
F/rC8lpFcOUBQ2zc9MyLgYciv4yCQ6qfe/CnmErq8RR4xIMubKQdOOBUm5y0ukHQgL6swNzafly9
V7MFiGLoKoE1ruoZPgx8pPLUOvXW7UYyii98xo4VQLVkBUNA7Y8oh61DheMuFQQf1ICgCUmazMd3
NRekIfnTwgO23A5J3I5asg0tm9yxQl1oeYvFjH3OulzyCFawqSIjUE15a5FpMO6sfAL9meMasAVf
YQxP4qPBScqbPPVj7q02iSiJV7LKMNlpopZtU30Z6v3++8hQGDq2nXLDZ1ytbEKoE42UttfUUT1S
jJdD+pQEEBhGgVkrtncZAbaFJp/crxGRNmTIVFfn61CKn+mrNqPbOrq1W1X3MsYAzIwzZl3k3+Q3
Ofm8wBiCjAb4HsZa0fjqNPJL0d17SP2jc/zrgWRhRtXMQQZLCK7z4vDC//GOMarGK5sZEuWIGitB
Jt7mux5kLtJWX+0Xq14p+mxU34Q9whahA6gKpE042EYqjjAlMOfQ34U6XWj05NSo/SkX/udAAHc9
LqJl7pfCv7y8kDz1LHs9j8A+RWECD6WX2JhjS3cni2d6YfV0khm7C8PxcLW2lRrLHm/VCusC6DGr
HhS7QuqYvRIkbJYVYucndGMwlrk++f/+A7j+cWQuoKtCMN3UC+kB5PFAV95xvKJobqQgUL8uW5gz
2VY1OyEXULZzy3E/N/ZWfO9wzdch7LH/5GlRKydywI2y4y3lyCQNftsuTQjVt8yQGJSa9CBYS4CH
SF1S4rnUwKWpaN1aIAsQzVDjMWN/K8qCeBPCQwk5ARTmrkdPA3GleFrJJYwG4RFqFkLkYzVlB7p9
pQ1QnF/Uwg7sFEXX+/cMKwpOTsqRzX6CN/OFYK5yCtCS1qhNnyj1yF4ZRy6lNgr0MHY/4OY75h9e
ryPEcouIPQd4DmQvdBgr+VaZH2oeznK3vkLpvRd4XOMNxTf1DT6njsYvEWvH10LGlFKW9dvRD/Sd
mBg7A2R9LHz3cR624MQfcD6PY5L9ScV/3J4DpM5V5HKpAj6ml3rdfszazTISKQD+cnjq63P/h9gU
NhSzybaOV8oSrgwl60BD4zv/Si0A60ATIqw4IyXyOLIQfxfGusT7kz+xhQBFGpuyaHlRRALeR5Ii
tutcoocX6Pag0cWy8NsXYrR6HprexbjV9CmjlBt+3ozGEbWParyt/ThYsbtPterORWOBUisTox/3
DqvujgV7qlY5vsdMawmdaJny1WmzeJNLFX9NDUxyJbRrhJPybiNxiIkPBTkOkZLpAaftUnBkK243
sJijc3FpFclYpRc2Xd5/QmkWwRkMCgGBHI5fEJe9i+Ng9pfDEvDVtwrgEDVfSDiVip37cdTeCH3S
BePIA+IRY8yzQ4gQhW4X2rTIV90NG/y6+cJA668tPNzuwdtUqMAmLFHyAxy+kb6gPl8lsmeaOb8D
FMb7/6URyw/DbtWmpQqNpBEsrb3SRrGgs+qYM+UA5DNTabkENGz6bdCyNgCKF0k9Dl1I4Qt4G+dw
GoqMb3GANdsE8Cp3A9M9dTKSAq0xFoILyvhPqR2b7mljVHrN/90giMS3vPx5cdr01AAHhqDUKNeX
++fjgB2L1FpguvZiIk0CuVQtHS7aVhlJwA4Fgzn878IOjel6OAj4AMF+d/oCYrt+cpxTfdUTMM0p
hAym5ygsoVskp/iME2fyo2yJ0Arnox9XW7XYn9yjo60CcHIPvnuarwa0xv3sJUe2Yhqb/Qa0k2jV
cmfc5hYG9B3CUrZ4aNdLxGj8zYT1ZKlH0kHtN0POaZLhL8SonSfnHkEIh16Bir6OUg6w/tMb6b1e
LVkgCNqO7zaDSq0EGJzlRnJzLGYuh/gOh3dGpI5MODA1cn0Q8GPMerQuMZEwMWCiN/MOjsAvJ4s5
1B/TSNyJ0WBh5InqBueB3mE40s7QXLu98F1iNizcnDuLKG0GpUGbToeFudGejVjG6TvOMwbMT2ov
ip8G9uPbW/pb3yp/coa8OkkRGgoQGi8leaOo07RZzqMR8wYNzE5D7VpIjbdlzCZr297grHClCKsM
JWldBBg2+ByIJLiQG9GJ69TlvyMBYVPR4oxMD6MYcxAwzGTUWYtdm935Mbq/Ccv967HpuVJe9JCY
gwOqQsRNTnAvyPxfvpjpY8mINmxUARhWIQ+AjJw/cVGZGh1K5rYIS6RVvsiNqYM0Gqt+VAcOqP6o
+PKJ3yll1mTaGv/WQ5gj6tF37CM58E9CkoBHQ82UPR2bGRaG7MqzrRoRIAodm9rJQTp543C+nwcO
fxpva9LYgH0loNt2Zm1Pgd7kZi8wPZpmHUP2bKJIfTLBS0RtWSWxRN4GK3TKhhADiGd/eslCHaBj
j5NRF0Bw/Zty8rCU+kawoM0um+oiqv0mhgSKRR/hHiIP0UfQVc8NUEY8/d1QHDGZcevx8QY9/bkk
qmti3OuVZ2BC8h5VNK6+oxRfZpb/mD94tDjpdyxbXh5ZZJhU3Njs8tMixu7GARPDUN9R8Y1/cLVj
udzg/r8jUKXyrz/pWWQ4dbXceRSi4em9yTv49DELz5Ugj2UQ8lx8PBr5hjncM7FYlH2rxsLwL7E3
tF8dGFYKD5+z12GMAKwMTeD68Fakd/WcFTeQnpBg7UOUn4W2HPB/SWailc/gDJWJvQfWQQzUp4yk
M/ZPJC/Loc+C3rnXgz0o/GEwa/gYVy+9N/jJWxjnUqQpCNS5TL8+R9kawkguLF8QJWgwl7RXKnsU
6/OV+fTpBGtjyMmw3HuY5ZRFjGUPIHKZFONq3TUd2IhM21dBMZvSZ8WrH/Z2a3PI8HhnobLMOgzX
lCDlHKQHwHgVgvyGqHoAw0HWlXx6IZDSS75bGc6OgDnss/7NUB+tHNWGjrveO0yoxv+h/iAEtF1y
Ob4OA1NzxQ+Xqwpg/40/fAAuZ1yx+WNmUW/1QygvyKHrr0b1eZSpWcJq0zoepijPneCYuYESmsJU
iO65U/VCx1jFxOBCNUl5sj5KpiPH5f+DGcExJKmZJHDuwrcC/lt09YVFVKv/cWfqIJP4vgwTJvV7
nScufPPeIfXndodxk1jb1cyXUkxQKelIWXtfSNW5rOqsaxOgaKBoyBZpyrtRmxp/ve6oATjluf1F
iYfy+s3XLV3+O6Ve5ovSr9B+Qn07Ci4/TBeTsul67rS1J2U633YRdwJDY4MxjJ0wS2fGySgNczve
PJetyo3cvQglT2u809wZ0/9N3xTXJydmDZbNDlmB/jHH4LXDYZGcCWqoWB1eX+ubarfTDmtROYyH
GWa8p9TtU8OTaJ/s+zIZ3v2uiorVzoitEp384rfJc0edt3RyRwb2wuBeCw0X8G4+j5SIZJ5Hlk6I
7AoxEjX+Zyez9LnLJmR9RkYYVWjebzcDHuOUwyEMOcVwBCbZZAu0SI/F+aEKCwlt4qSWl3E7icEW
yqsKsyn71hn6vS+FxDQ3SSVFvXVsXI3CfULjdiLu7Zzf6++OOzedjfu9MGld4C+s+yiH6AeOGZ/L
wGA4J3HV2fFFN5lJHjXHAWSPjnpXdivkOYp8mi8CrQGI6+kU4Pmyhuh75n/RaZqmM2onmjinQzru
6SoOF25lEGtCkKK8ZQArdmhOI9OGkIUwWHZnaXjU5cyX6xUYNThfr8R+VtKIQ+DUhPjQrj44tPpm
t/pVoezu80vCrzX+vIPKtOoqrEabisZuVdRHaAM0RjDwiWE4dtz+iadEelryNd8DRl5rSbTTLBaB
6neIpz66QfhqTR+bLumvjisy15S1mqmRlz7qYWcCLzuhQXydNOSMbk8lQ4EV/YAqg26nOM2BtfCu
BpQyHHEynxMF//+yBtcyVsife59jFm1pFAe+VaEZgZG8u2z9VfHSiKPG4RyM3rDtQ7AVsUdEParY
KKwT7zpVkPTuYW3K2bfOsozgG0jbDqRz/tLMF9Gi2JKeCW7W23L6+63AxcMviV4Wm0xzWX2Gpvga
bSDZyKMbmRvvAHNyMVaC0HKqzgOAdcjTKxmvt0t8jO0gWJOKITOVOJwi6XsmrhumToV6AI9Rs+o+
z2czErdwWg7iB4gFk9Pj1yQArV/cH/DSm2/ikxBDclL5fY/qvPAcr5JyCRwtaWtcKNDpwDktFT3n
37g9pSi5fRI+nwAQuDKyqbDkZ3iLfsxhMQfWyNDKG3ftJRBHGJGPDqBCSlwbsaGzMJIZmGdNHstb
L6iwoxD5mE8ZbK2Agz3QmnSC3qAIyr6AnMkPAaz3+ZlJJwXK9Mpa1g0Il3N65/AwOCr13Q45iSKV
JW4U0zg6q3Lwt9J+VYDhBPkWWbPLGEJFov3TqoDH5ukNEz//3fhOuTw9QKzWVEF58QuoyTAs55Hu
0h4T7NVxQUjWOoAMbbvWsNzhvzCTAiBfy/zsb02C/XNgOTjRkx8k3pi5RNKePbr2618agI7MnFpx
Xocp9HnUa8caVXcma4+fTCiXyMAKVwuo66s2CrI5/K+rae5ZtOijHDOrD69xmTpwRkRwGnoSr6RD
64EaAAkgO6YX5PLDnAZxj0LtJVIP2EY0ckmXcl2o/CC72XVFzHpN8/7cMjxBuVrTf+D9EdzezzvU
XMwZ/UjFDbsa4Z/52d/o9lxmc+g5RqhIvQw9CM1/z15hCVnyBa02zar9Ti9suUff0tPix6dtOn8a
85N+7QxZqbwpSDN0+PC6tslmrOBolMgU3s3SwxcSG+z/5bb/CXYKzmmBkL5tL4DirdI6Ce6EOf31
OEfeMFAINdBEhbVEXlvkyBcRWR9wvKcZmNP5WlnWKP8FgbhitReZElr/dAhwzMPqsxxRWD//P5hI
RzEwHWdNsdcoc7c8/wzJxl5uTpl2Zmg3R8IyJeaWcRYa01kmPJyhGXBisR3uOYqDy8xZSQIHStdv
80goWvXhcwxbCXbhFItM5EsLeiYdUICPmKiWuEobOlXUcXLfxPywf/otV4GO8ANgCHh852sHoBYl
/mD/rCOcq0isP0eeJ8ju34RazrviGsr9EhOW+QN3TIdI93fYo+jlRRY/nkZvcaY2whoM501rPl4k
9j2gkKHplV6WG8PWcR8MTI3jQq34obKpC2/ozVgiF6yXKODEjEnZtsCR+nV9EK9+lQk7pLTtRSFI
iIU7FAeiBwQ8RY2nLohgPSfengWHgxL2QPsBoyKAkdH5dblbCwkOfaefMcfTMz5pTslgcNTeZmfL
9G+c7OA3iSwVFdX62nVi0JQHOcHV6D8mcAqyiUAnWkVa2cKqsdUyJ29+Gzoo6ofaHuq3yECFfbJ1
oY3I1kUrBBqYpF0eWWdyiSkL7PcT5b9PuaSOLsuScFiLlEmO7TGORYo+nr7ECVljM/FR0Bg4oNEH
T4Qy/thTWsF9KgHVQ/nP9E+C4F5kw8lYfqlef3IT1W2kLYUA8yrgHR9t1LJMeUw0/qxbVlBbbGWc
9gc/GcrGBUqC6JExB7PNv3No45B9aNbNAftaGszOI0kNKe0ndF0au09TsIqnUMHw54fucZGMl0sm
JkX/AWwuij4eJdo3crOAZA20vXYVNvqGJBOFyICa2uSRnIg9bEqtcWIBOCMLUviwRb7rdekmynG8
bVcU7XAGHNaLO372dEc3FYeOMLt/byiPQK4FAKjlEDHxPhtmomsbLZq6v/h1cEWkrBXjdNQdk6Wk
OYuuejDeTb85ueRf2B/ua52xO8A74zpAcNp38qAgqila0PKc9tuGqMo9aF/4MYzcAx2EaJuhX5Ze
kEcH6QpqCY8gj/Vti4W44Ie4stYkqeMbSFnnyig+DsNVua4e9yTPFypZ1aUPLZCVVH2Pyw3ev/n+
IE4UKSBwP5aSa9ygOqrJxKjjfZBpmrBIhnQCQ9rjiJy1JY9NYiLp81Z1CyS+g90Q1i1S6fWPPupK
ZZdRTe88EFjc3hRNJ3z94ns+0qf1WnpRjWc1CWfRoCMXqSL10NxLjnLrgUHAagkzlETi4nSC1DVk
0TCTAT3P2sS5M2BJGtqQfht40v+J5PkkVfGA6kQPR/aWrDdOZrfIRq2UWwWA3ZRhwUWvzunTtfZB
2JOPQ2M639xr/6+ta1uaeTvwtzdRA/x7F3V1jHHM5qxHZqxt0/R19SbnD3pvhYzSeEP4U6njymFK
hSJAhbB/7CQBEpcj/XYL5ks8cWp2/nOBWeuZPCSPrK6fij8/sfwj/9zILTKzUAiW4QCC5gNXYqKE
FiLQguPvBtY8UnTZ7+5DDYTZnE8FIncJdSWRsQ5+hLzDLK4xiyDUszSNyHtCNvd7IuN7Pa9t/XSF
13s+g2xVbTajwFzIXmdbukxKR9KjPJ6V0BwjeU3VH8fbyU7l/UUapNlCG/qLJyH/uRkeX7W6KJs4
OLjogTIAof4LRS9WZNdfjpVDpF5l3Ld6mSYR36ClQvIUXs/Pv/vLRRBSR7r7NHMS3hrbxLUjJrMJ
EwCGNRND1dG2Bn7yYaEdTbxqz+j3TCDZl1ct7w1iN93QdqWsjGv5picSaLupY3hZ++pRHGUUMogY
HXHq1WZ7Gt0XuwWwW917dr2Ov4BWxJClZ2n6bx423CcHjfLgTLRnSCbLE0/8kyyR4ySgvPsGnzHz
1S9k8+h1sXBJiv2u0oCqQ2dqfJAn22HyhkTAEN+wDpupaADnAYR9/yHJ9PtyV0mEH91uGOijetbl
fq554qJ+Iu+tMd/wwFN8du7QWPrs6xuWSQ508EZLzMDNJNETOMi8qtNakn6SlESv33NAW9G3a6ct
GCAzQuGTGXz23jOambq7tW4AUqtbL1XSWUYoQGAtuC+gcHpOLspi2/ODMLmqsMCIyY7OA20X7ZG7
u8a0ntMJZ8Q0812epIm0HGpTAF+TXO+c8WjfN6cld23aBwBcIa97trHROciA1/jvbjBlKda7W1K5
HaSrCh5DvNLJybrm4ii1s31LV452EtRT2FkmKbKQQwFd51A+DMhnnNJXoeheWH8JGF59e5vCNN6P
P2A7qHquLXE0U5nFl+Frdve0NP3K5IFJTWsW8rIE50oEp3zfZhu9gDL/pMHJJe+SywmFuHQxTG/5
w3wUEXS81yp9ZiBVDkUbuzNNFNChvxWh5ZWGfTiUVasyB9C/Fqnz6QaNLh+jWFedeRfB/NQl+5W9
VYWHU3YIavgkfnld+kSD/9ccg9nk4ZhYoGO6HXlYSjRiM/ERPQSGZwbVFQEkvTVksetJRn2ePq+D
QqS5l1MU54cEp5J5BfdE/EoT2AxYf24b5FEB03/WnPYl3WtjsLzMBoIoxdKMg9zI07yf7xc0bzdM
r4mlhJfBludmOmftqM8Ov/MbGCVmiubdDk3norhmeOijck3xZMYXeE+KhRFx4hqU4yMsdVZOQ/0x
9Bbhb9fBXgcsKQnM26Ylw5pVa1zH74blFCj9aKcJYQaH+mPUsuBTaIwJH0L5P1MKondChZQu5+QV
7IihQ9yy3sLdia3jkVZOJluzp/f/2ROYv9i4l2Ha6wHgW/AYQ1dY0YM0dE1ttk0iNcUBBTu/Pqt3
Zx/6N0YVo6XaJvboZTH3ZAmJBr3GH/LiXZuOt40mwuKg3WsIRfYjmGCZ6vIxwMCGD/vxVeAnBqzL
X6t275z3fLfxURkPaHd6VtOiBe2bqM7qge3aHz3IcgAUNugCeGkehg09Yu+kKcR+U7zTHVzKxIIW
tSNrHoGdeYwfhlWpPKePKhHlvNbNFhSgiYqkJTbD3lv0Wj3gT/K9KTLxXe38TJL+0Gam81n/8PNN
Jdw/fMqbP3/32PJcjSyJnp9NwV9E+AyKiAkabERdwVaq7Ytl2icupYEuSh/dKfY4TyzPZM64BHNL
8EJOGLr8lmUKq+ROlAyEuqyuyF08yvbwdlVxj5wX6Wy/oRsoCY8Nzrd7H8rEi9/y+0sFUCWDkSFR
owypaYzB4nL1FW0PBsZZ/873MPUV/yX4qQmIJj4gpDXqWyxuPBxsHvstYT81+YcXYbQTP97Rl9xQ
ZBt1sZybC5jTOLCAJGqs5rJlH+rNsykxnVRm1BV2hoe3dvOMmO2fqGNIPvxOr2ybDPVypSzWJbuM
w6ARtrlLdpHK8RMdswij3gxJuAwLLMqx7Z/6sNTuysmc2hjiuZXBqDKlEeBLzqMJ3f3vD5z22KfN
sJn3BbgiOsYd1W3H/kn/G5I9sAKA9Uz02kWt4j6jMBtN0YWrDtMpKJnJqhndi0Zcrhfiyk8HVlxa
VUClgkzJcU/MULgGDHLXsv1J+2TII6Vv0CPdnyaaaf6+3QAO8LBX2zW2UzCaCH6/X68qcV7zo78E
jJ6MTbfTxwCirsXC62UZU5nB7waCs19MU6CuOGCNZ5o0jB/wq3fwbgyosmqYYAZwuwjXsu4EdkT2
aqc9WgOWxJ1Wp0H7NjlXGeiVm0QU4EkjsDRMQuNeFOJ27RbyTyB0A+2sNLjK53aNXSXbyX7DW2rQ
ppJ3KnMg9rckStVu5ihmpIIRKVntknxdF1cPKjs+QntE440VJuND0JYp0nfnF7FtnGeldRzh62bZ
VVDex8UExIs0DHba32bWTfGO+3eKSDnlooBDB3npzjtvAUlftPNOxNhQ1C8fG0j8raHX0jor4iIR
9EiBDj+84lUtEqJ2ITH3bbisdOwqB4EARm6kB4mnKOXSU2Ik4a4ozoO5DFlXI6mazy9V9KQw5fWI
xvw1lLahxsL/FitySgtqKUpz+G5FWlNA+i9gXHQiQS5wh/7HoTcvoyWgMehdKNhbSWrch6zW2t9q
P7p/qyxfH9jwHYe3n//IzMXPz245QiWV0YZvfa/wQbrB7TJs+/6O4g6FJm+PNIIuNzdkp32+NK2i
SC5yTBScGriuxC2P+/QkQ6aQjp4eDAVP56BFCGVlbBYP5HzdK//SItpIy4ifAiblr2nIR3c3rZu6
lj9m6kzJm+DbXzfIoe4xEWL9YkcVSN9M6sdqvt7brrUgmfjvubZ94prNy2/nVA0guPRKxo7XEiN/
LSPPT2hUMRxoGu9SfibKJdcqx1sz3O7oo3asc7Xe7hAjD0TQ3fyP9+INqEGq+Z71d+A8hATErkxf
welCcEvCPi5DqlNF6RKN5/xLh3ls3cmeal6YwauyL1sH6V3AIlRdrlH4lpqlP+F10DJbFlRpJ8ut
1ozC+IZG5SMa0Xmqf/j9etSev01FAtgwUuG0QVpNGTK2oVua8cs/HvlP3QvsqmxrW6dTJLZrH+b+
z6l3DxIB+BsGqKO/YewICSa8WxjsEcI0cyiXvieNPL/ZGmYQ+M2PuCJ5YtnzfpXmG5fJDmRVbbDw
lpFgHaQS4kL+SaMYNl7E6BQdIfPGsYl+tPxupPZzf6ar1B1nW0z4JyVuPEj6tzRd8Cj194JPPPn5
yHEc2ZKxRmn2b1soua9xSzUZpl7XW6NQ3Rz75ZhwYlxPP5OFTfpnDWlEUzfO901gRRFApoY2XLCz
nCpyakvXl7gUgAtH4DgNM2Me+GstrPux641l/4ccSxAV4hOW9hJNtqoD9m/NreSb72xtg8Ig0rpN
HsPBtvvU1WTwM5mFNfLkdZOLtdO1Kj0JbGLRLfqOB6dfAY2cwCeTWCtqoQoOFXTLdVOwy6KtbGDt
1YEoPITv83AMEPjfqqXTEGhAMu/w9pwe74+8xQgWBnOq9izQP2hZCNETEwcehhiZK82US5V0QRCn
FiV3wa6z4sqO4JAgemRIiPtgbm3Y2ZJEkmHen7pUBExQsOJ6at3zrvOytSGFk3tJPk/v++Y+TOQT
ssooYXj797cgXQ/tc9wWAxhsR7ZqggqmxNXiNQvVEmN1tiW5XFDbEf4qFF1M6T4QZeH6T4IcBw1j
54PgT/zW40wp/2WH66oQ5Qj+/VdxU4Pj7WR1W1EQVRNJNHHwydwvmgLco9ILq/0yR4ryJLUsu8Xv
TfWTYSh4qoR3c6YhReqqpthCqlSmSSZQNl7Sr6jyz6RQlqXt87zlI2olr1H4Q+W+u3Y9JwrVa5zd
Hp3ID/wSPxUHXtVF5vLrccGEdOp2SOTpqM28a2y3O6uRuPAIL/b5irqHnfLaxAV89pFRcd4l2zUO
L8OcQWZw+6OMtCdftqbGzAQqwd+aZzPBkix+JIwVp6CCZDp+6kdZcBNegfkgpQijAx1P+P2RFe5I
Yxa3JuC/ua0iSkPLbKVvzGIe5s2eKcF+9x5Fc3v59yxUeNo12dGT31IT1FuPAVnpLbtybnK8H1Tg
6jKnKriCTxjkck7k0c4/GhDfVGMNIxCDwuxdfTH8o+UbTqk8TLYHzIws7Wpb50Cf3eLFZZAcgRhe
U6KwpDCq7vsInIWWI0Wg44BGJ9GxUgYDC99utTMJMgzUPG0RYCQwQ9m/4QhsPp5+s2Vn1uYIkLaQ
5au8gfpbCcp3+NZOAvtfvf/dK+H7FfMCvbx5ww78YKWOc04HApLXhJcxvQ0HCQ+Goanlys5w37r7
CfC/LKBeJiUfKBWksTSBK2Vk9md5yT+Deh4cA/0zY7gga+U5RHK09dBO6C2uIER1inriTXJkwJXP
eluj84sn7GicURosiBYLwKmHmLxLp9pxFsg6lvTVvr16KBj7Na6Expn0mkMaydxdlFb/OryxyqWf
k20M/CFo9Pwc6SOS5crDORiMXbo53MKpCNe2ovOPv/FKI0lHy3nRvSnm4p74sf9xjd8FIA5Zhw/N
WBUBg8aOPOR7e0ujCgNJ50dx0hpzKSFDpycJ5up3s0luT24jlj0zrpXjCNBS3N7SiMmHq0wnkC+E
NA8g/aw5LZaBQ2eWUK8PzFErQW9J2mtgLyLkGpI79IwYazP1vifyGQC15asakHpLx84iYZVyIxDd
vmKN9h6VeF37k/Aa9uWyWbKBm+xba607xNG+3odc8Ow2bNtWiQjOU1Nrm2vuCYYhY8OJ6JKKF47O
IF0T/GmDbRyx6bHc/qg6nxpFaGlxuO57qLhg9EMQ3ubmKn1lCDbQhnv0w+lUWxsMWZY59AUYV0qK
2FGzR3ELme+oxNeajtC1PbkbJ+ffN179YXgt7Nn2fLaots7+Yqrol78mAHDyzsW93dMUW59cL/bX
NDiWtD9odUtI7NCuiVlND14kWE7F87yhE5L5bmN8zJjsjIIKurxXKk8RCRJJ+tvvCYIshbB0xsk0
isjaqpnMLoHe0yafBBmH3JfKStXvR9qdRH+7DPyvaHx1qJtbabZslolbu9szX0krwpz7PFr2d1fD
5EGT8+0m434Ct67xeGsPsvLWFn+KQ46pvfQCSERPL4muCxSGV7bRwg+Ng2jjaJzNe5gAp1bTIxSh
2tlGffEJTkG1rOdFGNA6U4jVAF4EbW3+k/64AOY6ar9JfuH/K40zoyXHdDfsaVlopSiFSEsFyUJc
oVApPVeRbkTnOl1j+REh2hiICUlg16/biVoBxlx1U2uuEzlcc4p4e3O0yQhp82N9evbpFrDEY0/a
SRYwWAETbRx6s9292NPLA6vPKCZFz+1SuEe5jpYM8YJZnyWJDxxOZ64rUMjC66535UCVGCrdY5Ce
Pf0yBJn/IKpvwmn6hbRGN9qnsEwDZtk8zePjow9RkVC8vphNguYwH35rJ38M+PRL2ElE2NZf0Cgz
zmEUUInFMN16E8WO5kD4WBtdT/o0vO1jJdPju3GWNn0VuL3keW2p+wDkiPShybVWt2gCqV+WPhdt
46f2sOu5YQYwZZys6+LDRjegcp9UJ8fxqgH+yKmR4Ju/YSjijdNWJtau3WvsU9WAXVbgaUwxEqpE
m8Wu6xxjTDCX53vGD3b3daSjMgR6m1u48W3v0r1aR5l0oFjAithfDSt/s8ovD0cqsDSsU1Y6WyMc
ZxwZNJ/qoInmnf+K1+r1YZfppYPJQ9pm0yOTDVHwB7fvy6EWPNt39FMBGC1z8bFDsPIs7L0tfiJr
RC9/Q8ntxOl/81ElH77qQrLKhae7eNkN2/tLUyNShYqaxGcNiI0xHEutlTnBZhnrToqQrsrbp8Vr
z0f2rSQEsHxgk70x6rgYmVD3xeoFStYsjk0Bu+RUOXP4Jto3q3vDbVLeUyD/vcaRX/15PWg6EBOY
FM3AYXTjerbrtsj2WBTqLa/Nc4wNd7Qe3ivEg51sB4zw6kk+T0MewG+prZjXrOIpJ+UN0ZLebuVR
+muZlJ+8KCckHPFzounMKPngLSB2u9ivXkHaSrdc5BGdanDVjv69UK6foj7ESFDw59OzOEd2H7Gy
EXtx2/PCH93et1wQLsM2dhQKiPXbg8SN7Ffmi9Z5MUJHMQF0yImNTvhn8QgdsDphjxo2f4eUOhFK
Xyjf1Gq2RyoKf0f/45gDayye8gbCl+bLh31I7iSCGIVxUn3uFcDYJumnrKFDuJu5IIEGt84qCiI3
rRh6JAUTr027jI4LUSh+z7E8JXjooj0noisx/F7hHkXFjvgPDZjnaDqgWsvth/lMvk2LKEz4Ehzx
tmgiJCeOGKhT8xhZa80x6TTuAh42Mwm799e/YBzpocmW3UJ4UfnZj4ypkqH5U31HuvVy6oq17rjF
pOiRnDivuRknwyuoF1DHQlLXwy23WLH2fSg2AB9d7bDQ4i4ae0OeUFe6bZgYR0ldLaBvtVqS6l4X
eHMhSboLbK5FHnEE+rCc+53NLvlm5IFDuYjCNl1wCM43NbIzYoBFJdOgJFjrYbFUoCkTXYcnH1mt
rLqf7KrquI3xCBPnVpP4T0kSPTw1dpAzOxW7bNhBR5wBY9yxTGqYQvuF6Ex0MKzWCGDTfhyjeKP6
JhbhHr8FKS1asZXZYSwRj4PsOE+MOFQuvKsA7/lIB6SZ7dkttz4CgDzvcai1W67aeaAvrhb4w9/k
E2qMZayQaBkNf6Crda0Be/sr2F4iHSFyQ/kidfEAcDlDXIt7ndXNfGBCP19gOc3PFbwaK5CpAFFV
nS0qFuBCwZvq07POdHAl2HIylSXnghOuLJIvqzgRWZJozEu2Nk8hN9NfSBZqZrELWY3FwxenxCZh
qCh2vrPnp3g69Ex0A05JZJmZvb8Kvx9N/jDKUKhzoQluXR4AFa2t9/WGOJD1/uOTzcBGzAUYIBTB
M/K8wVE66JQPW6DGl5lo0wLzwyisfGb2/QU0blwfuCwh/fUbZFgpG/xF3IEGXs9Zmi+44tFk+mfO
XA6oTdSWQh1BEZlTZUqmLO6cUSZVkbJTJotPu7vKl+m5XxP3Ee9ZA1Hmo+/FuSRrU7On8Ggy53bo
RvgUKCp5ySuw3AfowR93jGsuUs2KklAXAsS1PwkDmrUi5MzJcbKHfNonxGV471byEkgNc06Ip6g4
83a+cxKCO9nRAkZoirD80Jesg6cxAHnrg+p6ZO8rPKbkNZHPjgJP1s1M/r33xQzcDAJjptpTaIP4
lkgRt6pOrHj2LMhR9sllInUmSQcvRXjtdgDqMOjUm+LPW7HvsZljB+gobZbyzzVaI6WKEjrsvHZB
7BknYLl4ZQR7+17maRbbaE8xfUz5Hu9Z8Q8WCLVen14lW+XL6luNxdb4Wr4+rt2RtIoTHQMHneY7
puay7RRpPebg0LoutWZc/Nm6WEcc+r8GPVrgyh6CF/PotH5nWbpVcAtgsTZQNohqBuKiXgl/WF5Z
J5qsspQWHRtalV4tWC/0MVLCO3DV7gjwb7Le5w9K2lk8qriAPaor7Q9lkeHx/YSI1nsBme5bHXHB
dlg29PJI1xvsx200B8SaMoEPtQr62Y3vul15stbfFqymgZN/vgJz4U9tFRYfdTvW8yjLtP75CJaU
owyXgBI2wrRVwlzcI8bAQQ3APcqrXPA8aruYVwvkm/jFI/MQZ2BDJ1J5eVoFUiMh/1Stoa9qeGpf
ovZyi/0Cw3OfyLv6W4LGLagWmLWGhE6ugQTPAZnY7kAms7k5/T0yrSktOdJTBjvhsltofiduDuHo
AhTrK0m7Z798vtAXGlv02BhmxeBw37hkdtGg8+bOZR0ZE9fXNIwAIhXMGhkDTWT39898IAq8DTSc
y/BAqxoGMoNMicDXAEfB3ZQjrWnnSpsuwtCMVMxtaJexSSaXoNiZDviNorC+MWHVdaWh/JrqJdOR
vdY9cLd3QhjK+JObIEg7I/WCEIIXnZXeT7sTCGg6epB3wSG+pv08FYLRyXPlh6eODoR0nZpI5bQj
239imdUmrl/umtERXfA2V4DS2Z2ChXGVdVfRC7MdUhhJi8+7EGxotcwQb87ih9MRjCjYSqqGvjtN
d2eoZMwncVCEl5IDvY9La1DLnWzZxBzX9ByjOOOAC9OhDHK7EB/pdLPuLaiA/bsESafkL5DuLwoc
upkjRN4o1Rnfa1NfmQM85bkXl2ln9wphI9IzOwf6NA4I80gSUEBAfoIZiiGbiHkfOcJT5u/WSz0k
6oDtDREuuzkO6+txgxzch3OnaMwhthhnYlF7/FfsrolR9Z4NXsXCQ6C+iGP4eAUCHL8qEYEy/qEV
7ijW1eUvDS36uOZRpV1SpxIviypIUExDP15m7h8BgS/AuiSGruRmOH42myvspp9dRuvQlzMUYhxf
M7p3ymUhYmWjIA0iFziVoloNB1BjYSti9Y910thVBxo6BFLn5g5pblPtlKIM+CqNtbmdRgGfMFyw
G4eqykGzxemrqguji/0n/ff+PE5/48ORQXoby3JXntPvk+l23FadvR3qfsDLN4uW3zVsFun6qrI6
YitFIBIdzWHLdgPNh3poGzqJuOpk64ZNKKA8PQfaXG27O2KgbnWsdksNgfFUizmdt3r4GVjydHJT
BSBc5EP3+RMpO+nBYvVVwLwCJ3rSVePKodmhramYKLKhhseMA83oJ0/jgUVbK9ufw6UBkw+r+JaL
RBk3/O4gabpMsVHFugLAqTnckh2qpncSpQvx/xXMspxEsOhIzpWvW2idilchtMP6/BghszhOO2pb
+xEIfirEcHGJreVNKH0NgeHGwhu0Waaqfwag6Ks822TVB90M0XoFJbl6JuwH1mhx3Q8fXs3gnpQo
M/m+uW2W9MDGTCrHqzevMRJzCoaIpfbquBNj71RztJ5CS2sNtobjyYr/M+/6gE5hm9mwKfkzA7c7
4hqmeluI7nR4Iz55lyZNlOAxSF4UEG9LJKOyiXKVJD3S61W19HYytfLt7O6J950ry+90X+9lWwnt
lgOaJ3F8Dfasd7oOAheLYiL4uaVYgKA5ObHRvVl8N5QhkAtvPITHbIGQaF6GSKNNGrI/kawMjvYt
ot92pzIFEKof4vFXJtGFUiOJ7bLtJYAX8BN/L8ZyX+vs46Mx23zOVmH0ksBvJOCcs6Bg6uKXNjKf
7gq+Y+iOgk3WQZBBFvmtEJcCSzIs06RBZ8ac4haybezV3XKlutIy7NI3iMsPjozoJD6a2SQUniPt
dxZXJ2vrpBq6lXEyoYmswnIo5EMe//q3tbyyVcZVqFY1tIyeXKTbX50ml/IVr59mKg2vwKOV376R
ncf9pNQvXkhAV+f2px7CTDqVtc1w1OGAQ1leSuv8hk6qWlGq2zjlNgS4qgWBPRG4Q4dGSexXAnp4
rDDq0DNN2BFtpEaaCYa5sVl0WhqHUdHgjBjzulbaLEUGJAwBiH8EeALbLMZZs94gmOCEHXporyGZ
nHR195ttaNdFl6/MaqNnbYvmL2Uw8V1o7nk8YNHQNONFDYio0s8VbbcTEgXnKPIxw8zRhnQRJhEc
fe0j7GCAHcCYQVU/xdGj4bLQjWWeJPRK/Bn9aaNdwgw0dtwybvXtwNKwxkj4c8w3fPO3SnBEnpM5
BGftfwarJZL0IY51fZ6j3UT5hh6VV9lY2MvBJafq6YGdgMYbH/okaYBZyRtiytfXckv6Vr7wv52S
+UDuQwX+T8lud3izx4sHL90LLZeGwb5Er96mZfm+rYyb0aeJItCUxgsMBkEHUiRsfh/4N/1O46a9
OthmrVkp11j1VyU3CL9h7fY5AMxIniQ6tvWGYmt6kkghTBd5v8utX2q2c3da+k5oa0sMsvJalgOl
BKu1z1Sof+07L5vNAKe+I+PjCk2j3wIDQ/wlZsCVSTil/BcKKohRossM/0n7KBkVKZi4SvIHwwSg
asOr+V2/ffq1FYhlRwyeEOelkvyrZ5cPuizC7Y1UcwBotepYRXebVPvntV3VGSFNqi0DnhEUhKv8
OcO5FvOIcXytl4Sqnwa8lMQQ1TBjHB65pbcl1auNGdZgJbrW/gDxm6mEzl9yPR8Yoydfqn0QBrrQ
3e+ltcLmu4gPwLn6MBKblL+LXSG8VJl8ZJxHDVu370D8BQmzbS6AUt7M7b5Y74WbDQkgjSkzmWl5
NHJydcd98ycsThWWBpoJIAHM1PfIabAvjHgy5VxWJ8K0df+2zBMGb1h/Mgcvcf1iQPVynsB5kNAG
qmJC1VcwnpJb0oGcDk0go4NmAyapAQDAlcysI4PS9bcfVpoRBfDJoglG8KA0HjiH0xIu3FwZwCac
cze4rIJoCoRiMYOGlqPGjEzRv7fob/A0QE7/M9DUpOvlroPGeOH5SNwZuVkJ8+R0fucf0PRydrfp
TX2ChvpXpYZUzybNu0esmjBj4ApYaAKL3OxwaZr/7z02tDvHaCjzQ2kzBwz2ppFB3/ZfIsP7aPLO
ibWksZFxdUVB078u5KjfyEUI2TWWw1L7hOA4l899Qxzm2Vtfrq9+e+NF1GoowyqW/ZXTEqb8j/MJ
H5NcJLMzO9EVbJYgUJ79l4MyCbGjaTdtc+GpFZfB93KlJqQY0KVZ49UGhne1Q9fIxEDTkleNmEoa
beRY2VMeboaP05ZNUumZmIzIBHOxNIcFT767auaX44crRB7grEWWAef5jqdGHUkhq3+uLT8VkFdg
VkAjaH6t5x1sBxfd42fbcuZnjFYkBkFZQ7tws36OmKICNGPcExfez/r11gnZY7HJMBxq/DeW8rB9
Qa3fxktEiI2G25aLkRlGLVZoCuy9IT/+YTKyZwrSxOyxAQmLg8QkKcinM+cu/uQrveiXa9usyJgr
R8iwQzK4SOxkvgwoYmzraxUoGpauWTWh34w+r3AmjxeeAVAmF/I4jMYlApb/L/eNo23v9PDV4E+u
aEUSI+2v5jT5FdqW00DTGIwUAeryT5QM8ypdSRBjluKP07ErJKHvCNktIwFXOGbi8gnYHGRpqiqI
6zPQ4khr8TvdnyncbmF6zTHF5usPAmlHU0yIJVuloTg+dOAKd0YdHVNULHR7YPiLb9xOms8LRLam
WOSe3koMBOHbQupEC2LYSp8qkazPQp/59k60HZdaq0J07x6ZguD2qLSOlLUojhQHwrcu9imzNjTk
Hx0+go7muXkCU/D3wXOmzZrteuAAgS+krnaV2GEtfTZlpxr/5qs8zxDI9pi6gegyFMB5cCEnZJhU
wBmrTmpf+am0M71zEec7ARXK3l6oK6UvZloOx3zVX4X8IdnIcByedfcdfuh6lEhd8LWVD+B+mfx7
+TUg7XDrJwxbUmpvpwUMAKgOhyILc9leToH2prLX8KsCI6EAFq6xWFv3d2x7n4U4Xp2HLw8W4eLY
tuiPKALYe8mKnaxc7MUDrlNtroLcwvh97+rfoJ4Q8b9atfc6cYsdQPb77LnvLT1jAAcLf1ULbCoK
Agb2HEXvJw73ycfbnK0T3JEQPexOPf2afuyMZxOdBi3sjZRZ+mTyRd271xYhkEgHyRTkeMnJPPcj
LaTwe8qbgV/Gy0sLImKsHPlCkwOx4uwW7burZCmFqEOBvZkQf5jRYw9wQ8reU03nEqTBjwCrFoCW
asa9TmB+wt0ODm5+f0SJkiqNDMbCCAbYq7xrNBaIifuyVIs2U8MnctgtofpUginS8aNLJ8Nms1Px
yYYEvWHAkoqGk3D6rwGp5KwKVyedD/tuAZL5chfMDtZ8SEA65ZsoeG1f9sSFHVKB41gvza1w+Dvu
BOAuWZjeDoQNDWey2TEhKv/hPSmQXAv7HwQdQSEBXHZk/Y9G+DgBH+TxE0UBBbQ4NQ0AyJ+F894w
8rXjMcVMgd2Bs3Z03RU5DaaeEQvYExOMR+HCy7yDmLGO6vSVXb2ayvPzPNkRejvRZsENlAeeAM/a
R/GksX28atyJsg1Fdks4zc5nziuLv7R8Q1f8EE8ijvT1RdA+yfp/QMfKIpR250/dMh67AIJEumOd
lIYnZZzW5mz/ATaJe0MKMBgF4M/8X2gTmovyL9Z/IM9VSpqpHmHoq7ttF9L+IX+vTOn5hNz6RkpM
5NChYHtioLwy14XGGjQk/mjQ/nPGKb1blcHmKuAh29mrN03mVZtgOa9oDddZ/5441qenQ0OEQRWN
Q1suBy+NtK0DDI70IXKbPhP+VlsoPBTAsYvTQABta//8ayvRjrM/gI85hUf+oWJpvKRLYAfjKRDF
FwpvQOTDz1tQ3htOZik4zh7Tu+RQM0kgYmfbFhnQNktIKtS1IDBM3CefB2Iz+RQxvh/BPZI68KgE
AMGjZ/q5N4FOQbZI+WmKfjIFk4hCOuWKo41bi8tQN31Wjcv0/rDXlx7forr/cEB6/PFFgubg8vgB
lOoa4KN+fyqS933ic56eN9gEEilTBMuNSvbY0gQtg/bGQu7xq7W5OjKg1K60i1nHEctpmw0O49hu
05DMW2fRTok+S6wIzMZ7LCJRpIlEtvURylDOMcxpg60VFuKWf4zZ5B1N7gkbzf5YQiQZzjoHeQZh
opJ45f96HTxUJjPIYGbRCT37zVKxZq6llMaHrw2jrdLyI1Q3KY/A7mmTyi3w5nsL2sprMyMUS85B
nOrYPNXmhel9Is5mwncOW21CP5/6WopoW6ZdaHn+QXIs6Ah1L0zXABGfcOMhTlP0AW6/CnOS++OI
k9UzZZscasjVaujm6SdwQbpw/D/NWnF6DMeaMLLEdTUpdf5GS79tLXqiwPcWglkqAFm56jyKd/F2
jige1BivxQ6+jBUTA0h3ixPpCULIhVCbiaHD8/JKUhoWTw2l6mlsz7Xiri3Wp61UhteWAZDF32g7
FCcewSBa/nhpu2LZqKppekJ1N45U4D4JioAvIVdaEzQMgeQISWZ2k8dz6+Ip5d7S0bSFWYzYtdr8
Msk47c2gzkkTZD63Fno7eag7VXwW3zHZ7b76xWxccsq2h5ep/m2WWjc5B+arhltS7uYO5UVbd/3I
AWHxaWXlxuLl74CXQTg7QP+06MXnleQ/iHt3zS19p18fJ3kW+rhUj8Gv2BbbPKR5DPU9lfE84V6A
jthPrVZqtx6HBOo+drI2TiIrx5GDtpnDc8tPI3XMRBwPHn/ofbConiRphpPQWv8lLuzTS397zyqf
Iaq/xGzE8H0jBwStr3mquYThxl0UHko52gVRujJ0N9MTnw7YvXHEOa8PEBw/JPw7XgSZswMHwJIN
U1n1dIXjcdDAsnkATxtFWxXWILhm6lW8qbsiDMbTAInNkVDZ9F28gfVrzQSS/8udh34VW8NltZ90
FR+N4qQyUmeFz8R4XdAzHdGaPJC0yDZx5tQJRrplzdLcTNdskNp/wAPX8bnodrRZlp5HGWe3k0tR
em3s7tqjO65hgIjyTFRAZBkoLGl4B3fiHQyqyWyysFXfFqhvZQ0/jh+gp5A2iEoaGX9a+6Bzacmk
KqYcW6UcV0ISQ9/1cme2ZKihmp/BNg3c/QXgFzlMwpV7lvpaR2RyXFzgXf4S9Q0YRe3eLId9Rjrf
VkSA85T5RUrvrveEo95BUIlFRmr1Wp/wOGa8u9SzoPoUqPaYUcvtyTbjylDnYw/ChkGj//89B8Z/
tDSHYvI0STYPRgwM8L1l/gqd1fuioL3qxJulXTFhHj9pp1EWINl4O1a3i5fl9VvFP6q9HbJi+YLG
MXR+p4qt/7Pemxv2D3q2jpFV7sK2M+ym/wlgIO6Cz+FYGHh8NGoe/lpRIdPqR5sjJhhUyyZi0odA
0arTYRMhwNrICsWtH4G2lZF8l8qY6/Js0AtGcABYC1zZLw3/1Ij4Hh6KHBGwYVIvvE4tUNsohi7L
P+rx0IrDb6UTWwntFhaViZP4KAlQOSYF/Ed40wYppc1ttJiVV0J3AVxvjlwQnkUE2mKEb7ibmnKD
AxzOxn92dFkdutTSVtbBwSJH++xdvErOlnR0j2sIQ7XAFVJsOIx7UAw43xhIvqCAT5+hgPCjr6hU
gMJDiPDwZz1X1sSPDrHwC8Hdw+GKJUuNFuecTBZG4I2va6RfRmp/p04170TvhlvbZGGpOE4e5NV+
vhq7vL1mx83WPeaaAMwWcQ9uFfPb4mf2OZGCd/m1iIZson3CiazY3ivYVfV6W5i3P1w1fYMWvtqC
gjUdY7wRS0PDmhJzOxJ9+cYvnDLbd+7i4NFULZT85f6vuoobre5rmb9okGZ1jEfUtyvqn/olV/eW
NZAsSXGopGcnvqsvFqap3FvYifkqIZZAI6OoSXPb1+T/81ik4DZUqzSI2u7eFfVF42O8jRNT7awL
rgRZpcJia335Xu7IHGNao1ETHdb2RMNk1/pW7Nzz25empNSHsUnxY0XODB1L9GwVuNdNLPPIUIXE
W2JNCWauZSaGRxPxwx5g9HJHBiRiOHNpBeFGiiHP/I15KZLnzEXoE0nqX2D5vWSw9m6k7vcEo+Y2
yiIWa/PdgnUxtIEQSsrU74iHjNDmXhKFeDDwDuITdu/dMhwJaAs9xfQQQl8HAHjRy1G4S1xbyDZM
bLMKssJ11gUf1O1KeuasBx2n87L2HboAxsxAOC/ojNLCHIoxO6CgAtacZ15NxtBTue5pZ76arhmN
u4zmU0QgxyYBbet6B8HYf0T4YoQOLiEf2uEm7m99zjatGLIKoVxPLlX4pt+0QesTuJ8HDxTI0IfB
B4CUcL+JOKhb8AamuBTYisYwkH88JFJtkI3M0eCAdKX3jH57pDIezKXdpzDZg4ariBWu6v5EZK9v
0gdFdiocS9HYsUnZZ51F/vJuG6EoTvYpn/KQV13+Epwgt50rVzr5RKW8gc69UCsLKYbUJtoL6Xx+
u73U7yOlmXkMIJ3zRgJHQ76xgrBHWrrblTgjO8z9H1opyzfNLo9QHEDLDl52crKretqN4c5mKcNi
FUk7pWCyCKoSoTIVROezZRjUng+XbxDLxnjTsltO2ylSZHvj2MAiJBjmACWYcEs9cCFo5Q1fjiYd
kxJXVtLNjdaeIObHcrzl+LREAHI9OXApZCGp5lE4E/dGKjW0YY2YUlYJZe3NkzCK2qrx5l2h18eZ
rDju/ABknQObaVkOsrTT2GAkwOFFBhRMexvjvQ/fiHYHbV3fb1jaj4is3WmOkimAxxn85M2Aq9SC
f4Xe8qeFzIlxye/eeG/L4IDu99W9JLsksLW0rQD0BXb+LMzxIxnQV9pDw4O/rQgJbQtmxUsUw2ST
YskEbg+U26R9gkhXqg3FDe40L9k4m268rmS68glnDQOiu7ZJrKEEUiOgbghnWZ848XNiT4SlTAbB
Rhgp5PBCXsb9yMKChB+TLUix3io/PTHDT62FEDFs6wHSBvdVA0iAQZlAwhFaaE9Druo10bVTTLR2
8bW8VsRtTqCe6IrFLN5Yimmq9oiZrgnwNdAlypH6JLieZdpYZdg2ezP9tJRq8yv/IIBfvWmL5YTN
d+7NxrYgsJbPnF2kuwQUWowOemV5+n7wC2oeAsW3DLSFZZaYX3SMifurEXU77SsK4a1ktst7e997
4c3lgV1AfEsxcnIDbDBEAF1XTYNIfIf3crvT6TIfdaCSaZNCwleh9vgE12uIf9cTMkzNVxLdV9uP
Z02Hq6yIAPz3z9ioGsTNQ9qCFI4AxjJtfpp4xVekZbszuINOqnOqULpuICSdPq4DXyzlRZl/K7KL
6l1KV3FWlib6qomJ3ZNBJQAtbLBVaVw9HrMGx+OUaIQrA35bQJGJlFfMTQfJiCvR1Uf8eIugfvnB
/z+OyGzFvR55oSqRI/DBXQTeLqEuxKdGZXdKMC1f5fRZlRszacU4qsDw/82t2vlqTPvJSmFEYKnk
ByF2zfNheUH4sMbrF7lMMkb90SG+HAFSA5ORll7JM0EqeXDsPsiFBVy7vnwWY4yc5TlgrSIKmRrX
oHqahRzVphPCjg2qejf/uHoNaZcXn6lWna2SySjhmz7KkxUJ3EDl9uZIkyJCvkH3D/Cr9epY/xyg
P8yRdC/zhBPbLpKYoNHGuaEhJvU7jeJBEJbW5iJ/H5XAS1NU06vp2O/1m/yRSK+FEe+4RYh2HGmH
IIIBbEIDaW0r2UVAsXekxQA8f+DAtsPT/SATLg4mnhaXd0IXK1lFWY5dnriI3JYoNvRUb42wmKAv
NTJEaQHWZrkuz2uBH4DDxzf+NHq3MmKoVlhwUYMxc7v7qzsTPqhSYirUKSdPMVusfLFvKxsShTHx
0TEjrIUlVcBdh2hb/o2+T6qcfp+1mEJXZx87LuEniuE25Yu/aHNQ2VhVopPHhYxA9PhMBxxf5sAS
5mVoi++E3jxmSkM+NXndPiT2m35vFpMJttwlMcgCTnP/ZG5RhvrssMW5JvfS8mXfVtpNZOePIsdZ
MiFo4y0FqUUB0MfhjSs27Rtg0cXeUBHJVeFsOrnrV+2MJSvi9F/5xCZ2ELfnfRK3J8dRDi5tIuU5
5C7PybqHKgj0Tq6fJWyx5Gfu+q7nXepk5LzlbFmTDKJF3BGan7kl8gFyYzHS0PkF3BPwuoeEf+8w
cxyIuSAOiyaEHz+Ss/+BVj9hJ/bRlJfOzXqGwqccbxtL68/8io9ga+VS+96wpPSrd9NNgkuatZVH
Fhc9iOHw3wXPybaEzuUDXQ8UqLO6sB0yEktjqwpHwSugd6Y2ZQnQpwOKpXDO51h/Pe3WQTSe3alo
c5gVYOLhrOA2vYNYETsHZHV61jguIZe246IylI/8CGNJKccw06Yu3KSWdVOTv8L1dFshA4h8u9De
8Y9gLRX1BOM2WkqylZg+NRjUp5/BJi4ndUHePfHZ8wmDAColHflkfw/VB3CCWY9f67f9/Ut/n6dB
ED6UAV5k1rTds9VhPbUiMQWiS0UGRwrjsdmji0SDkmxR6xToGclwYfLxKH5q7fC6BLqliINIf6E3
7n+ZVu0krt8K04gHs7lDp5IxYdmcgWDDn6t7ZM5i15hwlnJKHFGU5TF/5EEken2CJu8h9Q96IOIf
hDxx7jDdnRP5TUgSY+FV4OMuqv1Pll55tProXK793RYOL+h8pVq0NLCzWeNLCMNXSTGheGCUX1Vt
e1XRbYR3ccO6XaHzJBhfHvOG4DLWqX4saUKmPDe5v2FNRPPT8FruWUUfMos/XA8fWmulvmpFs4k2
UxgXeuBF6Wp47fm7DUVxk8red84VfSjOaBC5jnpYg53fTJNeWCmgMaKEcnLcf4aPGtiYpI7Ox2bG
PBDsWW+J3WpUWPWyy9jpQrSX65o0k7i81kk/VnOS3hgUr0SwUQfkjqb5nin1D3/s5bvODLKw6+6o
G72EG2ETGqudoNJtnyBFyViNk+gmx3Qkx8ZXt9PQE7XhRP7wZGNH+euQNXi44KGrTnxYf/YDQv8s
A3Z0C+B0Pyrg6o9d8B3Gn0FF5TBNNXe2+WhoytSgjcMiS/UUT+gfrDf0PGpQcJMticbH3TJB3Mou
wzu9bpc53vb2s01TZHDObmpj0+jbLULEM/j3+NOvE/OLt0RYi82k3Pn574Annrr1BmtKwmK6YLYk
GIm8Eo8Kpt9c+oPZH0wyKr237XJ0nzMFc2aVgn/SGJCwRb1CxlqSyhTEEuQUCNyuoVilAORdH7Pw
QdxA5EufDAoUCqyQKiahzyijJsDvMv9EVFhS/XHyWqX80INnkBAakHrytTLzemgQHi51FaiR21Jq
QE1SVfadWl6jowwkWRAKwOfA26hYSPw2a6d3/jxW+frAuWLz7d8X3eJuW6E8uJrKcWy4OS3J71KR
8AJGdcHbB1SzSo7RN2/T3WFmCEm/U5rjKb+IyXHn+YGTUu2S+WjWBM2VJjNt5WV57m0rvD8oYn9T
aiisGQ9LB+qY+ve/UvNpBIv0EnMeVbpP8nmMUAaohV2EGCV/zsl0L7rKPY/b8beNnhJ/XIZIlLvx
gMq0Dk/RcCxkAbVVzxOYhDP3X4l/rCzn8L24qP8egBPumZUXMMzEApL0IXv8XIJjjOgREuoyxibg
2rxgydWWzBXtI12e3N/k30gD27O4GidlDHbJc4JGmok2hOG7OpmQNZvAkyWIZrXQg1SERwNIIiwE
Wu5Pp5BZwKbg/pQrrIX/+9JsovADRbFX/pOYLkzScXgWZumaP4X/BKJIWa9RIyIykkUZnp7OE1ps
W37wghQf93DLXb24+qBe+kZm69ZfDKmf4PslQVmCYZDU4LnDTM1sSXdXiVxWt3mPt4iunEnqQUKD
xpqybIouqZCWej6mySQ7zIJk8wPbOhSCEhwbWCHWBiNkJXL4aKMTtAkG3mxouxI/ZS1BgiK1aWCl
2FPnbzHSi/AZ9vtNfFEf4KBIe50ol4HY622qIKzJnEOgrOwrAtIWPzhRP48nDiU+vPjNnqkSzSrA
CprdVN0sYl6feWMliMNbX+6tdTo7vqTPuGLrgTDuOjUSFd730QUp+rXr+FQ0DMv4BNZk2wcWmLXX
xmNJbVjEzmW6uJFRKh0q/aqEzgjmMxDQz8F8AmcRYk1D3tv++Bfnirr0H8iTpCJJnLcd+5QpSzyj
IO+/EVLFpXeeZgugw+6Q0Vd45KZzc5qlgq1DNrbSEwLQxRsuPDlBMs3qBu3E7QYjXguJLHhKJoC1
Tt3Qy0+bFCI7/8wdJ8GzTQZDlUcP+PoOe9yDHG2+48KFmxOPkZEw56vo5TFdmk2m5VSYTeJYl3WM
LqhxMQxv8rqtLfs3hQrN+51tc3BmuBxsbYgtfq0ACPpV16feqFihIeFT6tK43p9ZvAs0qBqu4jzS
goj5k0SQmv9wfnf4r2ozfC5Xj1buNHpkilrrycuRrTA+3kJDsXQEj8kxJJjXmjt81H+q/akf6xzE
4SBvmGpw06xubiAjg3LVODW6mcgxKYcFnGcZujB04Ou4h9mWUoEpGO8Y044TmwoUMR0C+XwTyWJb
jQPR4uSAC6pPNs8c3nM09bpxJCEKtzc3lymnirdrDbO966u3nFtL1AzymSBT1HPHDEfm1FzJoM8L
YsiQZixnRNYO1FWVQZGhDGztpfQT4uvQhGjUhJ7T6WJusxwpgrRnn7ImodMITPxDo5th8na8M5CQ
wrkL/5bmtWJhgNbVEnHlYrUChyKuwHDqfJKT2A6P1Ee44hEaWm9oIVgGtqZ7AS1J+U/wOGMYpgan
ADAic/+vJDFeDJM5cEBYJDDkz0ea95YNz1vHpYB4ow5iPfa0zR3y2P6G5AhoFczZA22FXCc+OUG+
ZvSYu5+f9RHu6up3t8L92vw4/mSMJf2X7tNCQnSSotbrLdGqelhHIyWV+nRlEV2d6niaY73Q29n2
D7yy2Bsd8d83/Nb59chfeQDWb7hZwmHbDCZaV+sQAdhrQD/L5f1e4YBXoMY1G+4QHRTQxlZPMQZR
1GAfOlyDUBsbipjh3htGvGaBSZbYZXH6n5IB+9oOz9dVhS4XWpsqepmr2mLfBNtfJ3tiKbM5c9xb
CZ3oZckUmP5DBdLHQv1ZqyKOLJdT3mg8njIFYRpkRccl5MOjTnZ5XmlcWVb1x7CFPpb5/I7i8NsL
fJICAF3DfPHVrjeW83L/NjS7dRKCBg23qIu/3J9iOyk5dbixePcGbB2c4SoDeAz49dQggeAnQtFi
k4tj+EuZoA9KbqLV3XDrcFm5EW721uyDrzSxGoX0eUTLCN1oq9ITUtyDp3MPCiPqTFDC1G7ZX9/H
MSjqSRCEs6xnm1bQGErNfBSOS+Ta6p2efom73htP25NkpllL3wVLwc+8XiRgIrG46rglFIlmE2Uv
rCBUNBo6qMMU24/H/aOb60bpPQLvbe6XQZb026Tr6N84fOIB2QlxM3B+eTJrRFDfOF8fqN6zUCmK
7s5ZLdVrY/uLSYHgerdLUxX8u+16KTVM7rlNuiPNxSOU3Al2NekSboeaEWcNAxZb83Ft7uQiqaKx
QrpX+AsKXd1hag0gj9hwBPNPh7neyuAOrLbarfLW5K8Q/aptJE+46b2yGX8vhZaVzkobRYxJG0UV
NI88b0m10N7g9s6GgCiG51W+F6VcdkJB2CMJLTbT3EEJXO3c/aZTM6wJ0f78+iXqWu/OJmAKpWj0
AZObE8Bf93kZrvsdFQPKTf6AMA5tpqB7dlQYGf/K8l5kiOsxalYIfG6QMJ6G0z731l79NNgbefjt
pDp2jnI5OCLC+QniNRrCwwm3SQIwW77EQLCKWn9S3HKCfBPdnQe/5qMW9i3S+BCcsYy1mUf5awUO
WF9jqk1N9yHfAREPU0J+gsKPV7ih665xP+JdG9MXWUavJ47lKOBkE+67tG4GIfu3kSFKHwGNXpyb
B25WAUQjbMSjy6GxWkMWWD4WxAGciMj+WWJLI+BJCEDnZLbcPwRg7oraE/fmULVuqnyOuxvbNCOM
4lJJtrmtDc8WSOsUwzKLTwpUKYvJrZVzBghiD+A/FMxCYHQoauAU0HGsa2SK0N9KNCOnwaQ482/Y
jS9kOue8Asc/PyMKPRd1dsF/7JsbBSXy8gH752/KQI45kxzH7KpEWW2YyrBkNC39UpzwEVk6gLEX
NModI/DwUbGCDeusKSLYIlBbYc9oD35ifVkG64gYJCcV07CBpmGi8+9CH0Aa4L75azPZDvHeMFHI
KONSOd2nmlTqHQNMoZF5EBiwOI2bT2U8bLX5guqnZQrii21O/O2fF0o2oIyuVdbPKF/DH1xW2rRT
Kgnq7FC4oxaDSRVArJ+kDwI0L2ss5+vp7ksUQs0G3Gz51mhWSKkRGDLZinz0tev2AD9ao/X5vuqT
I8AyOQI+hIsq6sBHMkwqGU59bY+7UpiWytSb0snmmuI21BGeWu56zgzDynZ5m/hlp3xxzWwwoH/Y
u9iPnWq6sHVQ8WMMo3zolA3O2TeO0FSBFAiS8RC8d8bVu3yDncSzfYVFCh2J7wo/qHP58ytAwMQ4
S7Dg274s8xohOJinJjRv48Eu5bMGMWblmaWMG1lVmXEyGoXqlIzeUUN1QPbHznD6zD6GDFGczs7J
ZIO+ArwSL+OiCC77FIwYzS5L38/AFg+i2U3PsTNqp21jfX+G6Hz2msPvJM/KXE/Xl8BMoQsVFfP2
+FmOrJq+8N0lwPIX+MTFl5bY9RU4VnTB9vv7rmKKUUvGZQdun8TjQcDw+zcdtMMpjfymPjEm1gWj
dK0M8i5JrAh6Y3EKCFXzSNe0vDF8Gd9L5/htEhc1YjIfOa9m55DIQ+AVQEkBu9gMeRI6pWSnluml
SQq99ISrtb5Wf86UhJ1C5R76YJIS5qJcR+1YBfmS00Z3BBIMlYGQf7u3f+AYFn3AFXDj1lBoaWMS
qXudMPH3Db29resJoAyVpCpRe0dWhZg7tlVm5T0Ick0mrqbHjwTyxbaOr3iRBDkI5uyQgfxu/fn9
4JWdT86UO8fRMglRqDVhamOfOOb6ewQxKt5rWupiFcsVZhNIhxw/jtF1BryiHlYG0sdJ7SyCet2s
59vee8rVqW+CXremmdy+OSy40OMNwCRJTE/UDjuH6f8Kh2RUIjP7QPMm6dDy0ptuUpr4Tl43fu25
P85gJ2IDpd7wZa7H1JhizamWseLarQA4nfnXVTksyDiOc8rVWXEu505zRpESciLhzluJKWHpH91T
v0h5CysHmPXns83sL4K8krVQ90VGcGUFIfPvWk2Nd37G8BsMyBkFi7EE/uZiPJzJsDctHo3wX89T
QnoNVOTT3iKkYnuRqP3q9zbhfueZmwLNeVpopu2uSaC6CI71EYYtTHxwSXXKlBYrGVfJjh5zoHo+
yoT4vx5QhGEoVfta2QJfGD8u3DUTHye8qIzzt77tP4MZYW7zjekCiEkp/zP36k2h+vpJcEJHjdjb
TVsqhUycYi+1sluYLRDvb7vfFttcNCVL4UxizxeLNqeYhyQMZOvi8LNQHsfCRHKAU9Z0ghDue8ev
1yFi6KFatfPNhf24JKpvrGIJX2EWEnTSzE2W1iK0Bu8/YSMKsx+TPI8elmV4x7JB3b6zGJTNbtDp
UrIHGpLn//ebyVxb3XEgyQYNSGfzIGAqlEJYmLz1pgl/U1K7unbiGG6zbcQ3nl5/ef9lIHC0G7eI
oN2MloCf/HfzF0MbR6M8uR4WhPOiJsMXRhuBLJ5zDtUG2lcZepgxvAWavfCszFeumaKwohmLDMWM
RGnYXkKfYZpg80u/mMZ72iCXMljjY434J6veQ345jpVe00hECr3iFGH/IdcoQGs1f53+HJLnFZBE
7pTIDqvKtvuhqaHLyL2yufK6edCRPijDhpjwlj2zxKO3hUc0Q4rfkk8quPhiD9JR46As6rXbPN8i
RRZw2goQ111aXbxBjbwJXGryRNiG1MOWWBx8y5HEczc45JU0FJfoNKM8N9lHNpZUsYQlKH/UfWg/
5J0LQhvoyx+1cHBK1+IbU2A+/vIQAGg1QrFVmGUzvVns/s9aqY2iMMILGiODVcq+DSrcoyzW2Lq3
CpnRDq5NMHd9tUlPzAle3MTrnNq9zjMZaV7rhNkTJJw3RWr+1OSOaSTDC/9jPBLOKnNSFQkOgnlk
TQs4dCjz8LSm5kCzaXR6NJnSjb6ypois7Hilbs+Tq/fOOjsjcsvFTe3C2Ttc4EaervlF+Rj7t4hf
sWKiio/1CZYTvVEj9grmz17ManhXCA/pGYNqSq/hHf6JAzznciLH2LV1OJ6Z9VPPxiPmSdwZ7myf
++L9T87U7ToZhifv69YwIdAHCjYj0vFG0y8n2i4Yzf08Q5WdKUGSFTTMFfGjoPPcMyGsoyf/HA0Y
T8sQhiWLoRRj+jURMcGCAZ++Vib0tzx3zIZh8+b464PMd5r2M0NZRNq9h/pusYR26byPuIEMgTJP
rXsKYkjTdgIETbN9tcwfGaMAAQznKrkeWYpohdarwFrg8B/wbKLWF5vqi2gHZjzC4UvIu3xmKrlF
rQobkTfOB/ovOyzT1DdJO409IzhgtPabtRC80iAPU9d6ubnPFqYXPSTxWFqMSFRcRCR/gw3TDPLy
CSxQTlIPa96m9yHX4dxUxvGmHn8GFb9vFz0U8eKZnl9378jGFWRdwm/9tFdX9Uin/3LyPJRTVgJL
fk6pNY+IfT0NBDrXmX/okSAa3Jgh+SVkrpqzxWo/umSoiBLDTxxUbdTlh5nJS/oyV1UwgtTGcBJN
1YJwRTFaJEOK/H/Zdgm7RZ2EJyuJir+N58gu4i643lKv7w7yejonCJUOMp7zZMH8K/1CnIrBudg3
iP1H6g/bKeWybaUtsd+ZQeQVBSJ202T6W4pm02AXdQ4PrZDfpCBtI1/FgjEMHDTc2zvuxJTGW5/z
vNCLMYGArIAisPHPoAUDR9LfD+Xct/VFk2F1i9wdTmqq5KwJWK45ow7s5axZZUs16A6RrvUDslTC
Qoi2Z1ishWB8ve5GB4+q2ufzGPcYdEgYwUJP77JzU5QaqPiK32IpscSrI3rxTJf4Un87DIcCqrmL
imSG2RfqqeG+6xK2amd6oAZsJXze+sSzXUZXw4Ht7RbaUHMUGw/TplXsaqm1l9nUDF4cvX7E7c/O
pV3O7wI3SnwOnlp041CNodXmgEO3m0d3qmnE8CuMAfjKYr1ysoiSzhEXwxO63XTXwECJrAdAU+av
hbKjhO7086oc4bhv4h0/rGTnWRjcV3cOq5Ud/D1DTougMRoDVpEmJE9Gr+3DqIrIYVkmQn76Fh+i
LsJj4Btyti8UKNvE3UTk99vNgw9lHzLQ+qRESriIiOeeAYwTHClBhIBGQ9WqrF5fxDVPVLmkg1qq
2UjkprhilB/hSwVMI/I6TfXi/b+EjMzZRKDAAG3bjMrSEVDatkdiO0ljadzaxgVi73q5UReOViFf
AFqB9XOOq4w66S/GbmPYZKKRhg2CNk+KAKErhFqbcm+ehOM6mDFwQu0TTiaCbH5Hk6B5ryQSMvZJ
27YxV8YOJtYWGBtVFa6xH2D2+sWV/JC8vfi6uSNtYH5LFuPHxuiZhu6ON1xWnf3NtULEgpr3/6/x
QcTnLFnvXY3YpJASkCzHTYdKFvWGW75PUucGMYQ1J7t0GipuXquS6LDtQPQXrlCSzdBPxyKtaR6P
wP2mvK3pN2ecY6nA/3/rr7Xj8WLYmJkYNQ/iG3ZxMSO+HoOUoEGHwqC0rNu5yeH/hyjdorhKzFf1
gC7lVy9NykAJStUQt63LODe64lkMCj3fAidwf8aau7y7mCyIRcBqwp+db8PtlUF85dplX4O+zF4g
xGnyaNcc9hVm0F1cNakfPr/gkibvzx6UW+kQVs35Teou1Mmy29t/iaJWS5jgtZqs7LAKeaET8Qdu
ugLnX4Xin0LkV0knPPh5oLq5HNheSn4GRNeNWuKZXtfY0vzuRcFrJxQMim9izIXPhEwVMfSGC715
fUUjF5vNjn3EC7JHXepm2+/9PCyD1ARv3yYpJHvJD7OHJNA8GfBHklYuArGPMLPnAEQt/1ReWz4S
BA5YjhmTmomXQ6QUqyjb8fxKIMusFYtoAXVrZR+IjuWzy2eVBkgGMTyPrs65VO30/UMhX6UnP0uG
EGp6iE9vh+zDxzBawYBR6OAyV3hr/znqDMB70E9TR68hFTiD7vJpo3Jw/5C5AvLUwC3lQOTpME0T
a1GhwlDWwzR8c9ANVeM1cz1Slsy8J5995cdTESQkQaOXJa7OeZrnkVs9NjH57Od9sK3lIVEf/XjB
GvIJxhC+ZFnI9Iscne+jA3a0qxR6kQFoN/whjpArVFONqBwk7nuKr2EQnvd17OAg91AhlnoCzlRv
9Y42Vfi5iuWSwueiEOPt4rTRo+u4vQHSrXvLbYwq1pvxP4smnabVhzA/Fd2/DeKSNOip21VdCgKu
EJ919gey7BXo3vpF4TlOIAFGcq5sW8tuLyGwBqiWPQFmvgDyJ7uN23wCaCH1SOcTpfwInNf3t0+V
Q3s+Fp+UfnRbM6LtBSD+MewmwiFHeHymtBzx4U2nkiTTp6F8hl8FprZ1/nvbO1H+STruYIqx45xk
1C0G4jGyqq/Bikllpy+EUZ3cig67/crmzA66EhUu/TNKD9RGzo88Vf6bJWlJSTrMXeEi1vTwHS9/
SS8M10PyL8JOpX7iM1tPxIEw3pZ3w1f7a4ADi+c0UZjUULkHnuEtB8rv99ZeSJDXIhMKrlMhnepZ
foIUWsVtovONWdpdcKgaTwcohliNh4FiZI0IlkAHUMfd3PV38+9P4eWurc8KFyV95ntjU9CiulKG
X7CVqQDHTaeLcG5FaSIVGOl9fEKH06abJUSLDSsqI7eU+vbeWDudgGGvfxuVfauA2M6JFIf+Nnc9
Y5yJGJAROzth5W21M8v6v0nKjHElPR556UaW1DqFjpAnzBC8cYfDx3RZvlPYqMwC4K48r3n2J31k
fdgQV0eBq8DDCDkXT2InFdkzMM/+uWYpjulrtY3TXuM3ZCbOwPRH/E7+eaJOnAmpBXtIOHHE536e
v+6gua0sJYA1bMrxR5nO6iOq9n+UYD1AZ1Hpu5O1bVMiR/b1Ct9VUh0ORNaSUbpp0OufTRsDdgZm
/2jdlKKqRQ5weOxvGF5xUWfllVqrLjgoSG+oxx8iZ7DgA5fKuI6sw7xQi5eHiVnr0C0h4ZTbSTXx
NTnhwiTO7b5MMjRxTfT9noQ7a+ImQeD9kC2kODpBfnzA2cQRJcGgLu4nCuLlsRUIb4ddRH7eoZVN
HYf0dF4YO/KkslAU7ynT7FhUaMrLKoDZzD1rVcpfHaXPrd6o74C4W98Dq/Rlys3rv0J0LUFyO3NY
6BMpLVdPURfzuWNrl2K/WNWl6C6x/N+gb6CocdTXn3SPd3yJksP4VMvi8ZNRNlyBuKMQ/fidGDNr
+cfKPTS9uF1wX/IxM3dSmgit5sgaYpKIjvCKW591ho1rKhcJJc2NnM3tPtFSKlMRPFFqOks5MZWi
lqBl8dOVBHVa4UPS5s7ENXf29u1raGw7dNVaQChv322JgIIU4oKe7GzA7lZyg372U36MkOxHqvIq
pHXHiJ45ivk0S+U2LOyZeJkNeH9m08tb36nMszvDW9CWpIMiPHXdNudACrbQ0+hUONfGcDVc1Mgv
TCTIIaStTju1xZFspnByUu2WOQi8vqv8hv0yazPtEMhqcITi1cDpiPCIWgGTrI3VFGov/iXzna17
UOV7oclRVFLNsP2FHh2pTGni6BbUgeYtQ8f/jXz7jxUeGjIaohGiiyjAEE63Te0P6aByeB3gouCc
pA5FsFcQU68OKDRVMDTufYX4rA4Rmx/rgTUKroEYIo0O6oD70VFPifr4UfsZsp/EJzLDvrcuMhy9
M449LInioqCcHbZgu/wfVDYaROi3jXI5mqx5dDah/8ZCl3Lk4iulxaAXm9Q1OA7GhMpy8ovYmTyd
SmPcH5dZ2t/5qpHGZlyfoaUQIY1VIzuhqAlyfEX415EJRkwL+UoEqAEFZ+UEr3iDWavAUOiIIKJ2
Bs9jOHC+1TGe7lbooiQoG9VbpzXgGutZrIjNGQuZzB8rv+yCw/fP7kjBk3+pozSu9OL6KnYUuArH
Hpvl9EVSAydEPQiwpa6tJmMx/z7aet+5FKmGhkrkmjlFStDyk5ZVx2l4G0fWQukGRMjxMy+RmzpT
mYZoyQpfhwen4DkZcHr/Re9qR5W3ob215o5871JxY0tgGs6SmQ+9FtO5N99g0jFQgReovpd10s9D
msJJ6L3Pvmwcw0IRw7ZifwM/c+43G8f4t910l6U3LxHliXAfMaoQZ89lrQtJFyhILPYgsCwn44M3
6ywKKO0uGml873EZlQCrql4wB6v8UqPHoleC9iBehYvh3OGx24v38E4uyCxNaeg1Q42mu73iF2aH
ul3c+kGOnjBLZS9PeeVMV8ufFiFzOEFEvw2RGIbONGEehxiyy4EfOEpbe7e/FNbH0o/+4HWswkq1
KV85v6mTfG75KQ3K6LhV5AEXuFQNBlQcsUvaR6zIwv2EpRFZ4I51TvOjjO/85NLlAEmV6NKFg3Ew
aPwl7ggmdqvNpUetuc/M0EwG9uZ5TBGMgk95XIzi85OL2GUpEw7q/s5k3r2yzTdn3n/Q2koIFyop
q/H2d8UKliSl21IIsTTvJ2izS7WU/RA9NQ3Ena6DUn4ajsgCTVvwjRgA4XWa2jaF6t1bGvsdj1N+
yNY44Pcnbn1MvYIemM4NBuZF3mdQ91JjQDaS2ASEldrkgNsnPBk2cgpYksPZoVHietiaMab2U8Ij
kI4Ty7MJAJXOGVJkqTA4Hq8C5Zjgoim3MRRQ8rjJhMK9I46fuVyfYy/TYokaI8LJis+jwkBPeQ/i
R4jfwqxS8wcByflfn4gGwrMQ5sF4ZUwL/pmRx/eKGGs6WgKK76O/6U6a3o5PDWbvuTQ8O1peMV+S
3r4/rYmPlBsQbp+YsuY++kSAogPBleYELFFiCdhIWCuPf6XyscFNrXiVLCpVATjMbM5/mCDCKxMC
qHfz4hZDWx0FGp+11g9jdbfJtu7xu94q5nf2fIITwJN3CY1bp8ML9Jcu0x9CXL/JawR+2jnG26pr
FCQQloCg5MK9wbAz/q8AN+QBq2APSK+V6IoqoJ1lkmDK/4XzPyvf10SIv5zBBHsyUQL+/CQsUVMc
3k1nRpxkI/U3rAk39xZMJn7zzuWy3ksEF9RexyYXGhdbLvV86gMpKvvA5POw4rsqJ/x7f5fVTTVf
TgO+Q3kOfhdFdUcJCeojyTefg7oV9mvoiV+qhn3wIDmOYmkEC2VUw04phK8bSFR+ir6QvuTWFdU3
8168xkWwxqeanBQ1Of+jrrO1d1yG1BYRI2g6P4ekMg5Z+omch8KTMkckg72eC45UmCnCkV3UiFTm
Rcj4AnbO8uYGZbFLbgtxkkKYZ3lAqejGcFE2umSsEEDGmgJ8gqr8/CJ1GImmrUjZa+kRRW69LZpZ
Rn1Q9PNhlU5A2fSz/hZR2yzxp2Ye2VHBWw6GFAIo5/7OqeqSxfaPC8WeDvTSh+8LHNdctyNmlJlh
rWFZf3C/UUl/1uIEkHK9YDzDNUYPuDJZ1l/65yerRfzvpLRcXUwPzNje99L2E52BTTebqCVrSJWF
8rip70eghdYMdFUNaebGXJhecibqcj3tyBGT/YVwJChIRaN350g8quw53MZZTSQ4eVaJ6J2TsIet
Jvt5w4XxdGHRIJWX8de+m3hKwEsQTJ5rKDD45vgN9NONnxU3yXzg4kvoQjCqL5UlF7xdJuW5OdT1
eq0mSOOpXwW7EaBGdP8j+tvEUQXYgNPjo9Kq2Vmisuorm8+al05pTWxCAP5YI4sC80u9pzAD/QjF
aHkbTbwvBkvSCA94/1XdI/E+sM5NMGLSu56qOQme6123qv4XwoPEokizZpDVUSSV0s4QLLROzOcX
05tjcYYGlfLAmkXxb7iAyRpEijeewlamUN2SXjje1RgKRs5xKAp+SY8yTH+Psj7N+/Pa6PrnmrhR
CdSY1S4ACaasWRMAXjt9lLK1ZH1Jgz5NPcr+qPkPLrEcSsr/V925uXZbe8hSZeMbiBlRTk9ZWD8j
/W0kTtNYvKY95JJBQ9fHHUUpfKL7ICSe6ISx3SQm0YY2tCecCPLuDbFIcSNuzJ9Gi34nW3nFKapR
eL5CyT8i9tTMjbAQlEVPN3y6sk7/+8HL+S0E2gXIxz9+j6Bf9XzghMaj2EDPZNpPSnYKTBf/QTUe
tXDcIRFW9wzxjhq5nw9V4NgTqXjmtngZz3i7sbxWwv5sD00NiG+W1A7dbEq5FWk8a2b9XhSNSwDN
Yxw1hDc2Md7scURrdpbKMVW/62+hW34myokn5/aiK93pELUnyh1WNvxpZhhnaswmMq5bo+GvEjcC
wUfv5kfOIAuY8KFZjtNC+Sh5XZJk3+39mRzCVbdwGvEnP5+0pb0gbF8Rrin0EcXpbH9iwptmM3PZ
Z+TULyGWGHuggPwr59iFZRurO0Q5EUighLi+Xcc8ENIX9+e5zS3LwPomHtLPZtedUTvvwWjPCPMP
bsrUseuy3bWof4Sur2YH6O8eJmR0Rm0WpxwtKr4aVYaOGOaDXiw0Z21ubGk306s6d4wuA72nQZzE
1Qaq5Fz5ik7HGveQKW//aYBjlqVZmilmq9ZLk1MdEfFzDVrSoFKe7RRIYuWF55VWWWCYNqon28b4
dsImTeTJ5b56slfVvqm52x8rgrs5W9HgqI14oXrBJmCrWJQ+3Z8QLSL7k9vMSKfe/F88wpeCBeJ9
BadDIPEy93WKBI0ErC8i3Pb16btG2cD+z8MA1yZN43skJezjKU+KSQUTKhfnj4Jg0+CRVgmBmepi
hNYZoq7g1flAvsnFUGGwt/kzGL0iHQQKP7bNnlYieh9MRX3WwVNa3X1FwuBFhDLV26ZnpuqgM+c8
b6PetbErwA/ZVXoai62aYOE0pWfz97LYfPBFpH6DR746JK4/ntIYh8VgqIG76Aifg+YgZ/5j3uH+
hTsXV+quy4+QXQLT7ayMS2XtUDSNLQ7HPZItptle1kmHhWNmaSGU69BUbczEP110taEky2bzUvEV
jy6EJexdjMEzEtAYs9fkdRmHLvr4SQGOLuWbnE5JcMXOFAVsE/Zgm2FbaDs1yJE8ZDBnZtfZDDPR
WD4NJ7fKkVt+jEQz/HNweBzbuR2rqXogXwzUlQSzOgzVX8XizPV5c7IW+aq0qyo7GPgglX8NPnPk
zdjx/UmN8eV3D8uSqCmnqR1civFU2Vs3KZevPezTUPho63vI+b2nUyI7vxRUwOwVFSQbUkUDpxfK
ClW0RGND1AklyWle8zKg1mi5n2qQ/3k7Ld3VjOt2mo/hzY9Kvm/3U5jIF/2OHpX9cXuQ5/Zk4ei/
gxOCQwOKkLpYB6KG246AwFLYmLN7KdSVNXnLlWisfNfBNU0TJdz9eQKl/RlYIVmCnRRU7SFoVEfQ
XL345lGKw10pRyHQv/zb3XYJSizUIkMVTAdLLX5HB7JtHBkC8IcNgKh+m/Z+R4oncoU/EukRwiLQ
qSpygJXX1LQYepRmvl1ysbZSl7K+zylO2xorVEg/WZKgG51/bkEUEfKE1oHhp/DyLkD+Cjxny8E4
txzH4A4TwOTKVU1LsqwjVlKzIZxmx7YsjTNrkf5lgicXM9kI08rM9ojp84ARjjfdjuy4uhitvXDJ
PlW77Me73LzIFGkxEhRkRz1V9zH0glETe+KFl4jxAvdlUOFiz3UTbbohiUDPvJL002LN5qJqJXxS
t87JU2D7YiOO4D7/gIaeVoRG/n7OCpnAiLfW59tA9c5GYzrArnzplLI2yCz7fB7FNr1J1mrDYYkq
/Wx4B7XjOxnVdWsoyJ9OKzgmD4dnvQr/FMaOiRSjH81qXcCmbUr6tDAqdt16Y7YlrtNgVi3lEVPC
v9FdNc4PBzxMWo9SaANZQn9FDK7uV///yqoz4Tv/XqyJHNMdbOjOR3U0NIGlVGBkE7VgEcpFLIK2
lmvtQHFOdJDW8+zGhPID/0S1j4SODTMzQsdbhIRVF7jByUkeMgnlKMklA/qfnOul1pUZCTr5poDj
A0xFXrduJsjav1TmDycCfbR2taijnwgdEWwJWEtbiL+hIXTwOs8LapYhIpEgYC3KjnvpL8aRojG4
+d5UxpEeRqDf9TT6bbQsRj4M+sSJ24W1nxGCBfSWtSb+agGxIbm8NmoneCyTkSVgP5uvC0RocFCE
d2190R2Yfq3zuN89i5r99M++6Iaf5VvCvWTqUDLnpJfcc4uWm2F+0xQd2y4HzlJmWusS6UIf8eMk
E39bGTsQG9P8TlLhaaoajnh1zyN9UHcUqoFOCq/VObpeNMi3hSc1GJuQ6N2b2HSY6p03VhgG8Dab
PoFSrEHi4wxvaSxZoENdKnvjzKFFE9W9zKVsF3RUzLbHNKIpRfE92Yt66/f1Vbcqqw+bQl1DkqiV
p68Pn5rlmkdarTq+MFImwUFEyPH5cuNk6RbL1yk8kdUnHd9VCdKyqWiDcJ+rsqfVbVm7zo6izVTq
znlAk6TlJWocHLA08j9OGVKZBDc0ReNpCR2j74ziWRi8BrqhRBIyNMyD3KzKbZyTUzAbIC8fsCpU
4KdyOmJAE0YkF9O9XED+jkIlALBkqNj3RoMnteO7YWTgF33ITA71f/ox4WlQJL/z/P2rLt8e386E
gTB1M5mHKHD4MMU3Z4HTTSxrxryHiLz4x5gmdGyHkza2T8SV1EwrWC3GoCM+yFLk5LhC+KFWrkwl
mzqt+amye4d34lpYw2o686EPkvTiCMbGuCC++D7Af7sn87ETdOx/KB04SfNylwQnb6kDKJz3wCwc
z/neVvYAoocJdhKLH15k6X1KhunyTNGSAdxqkjFDVtYs2XzMwtberlUMERGuA8jHH1l592hd9s44
Vhly3xCqlSdqWEObee5WAtTy5bolRNl2KrdfrWYcDM3s+h1ab0zzWTFAXVb8aZ9uK8bHgfE/8HTQ
EfrwwXO4oRicdplh14jJFMGP6OV1UjG0EsxkS3lx8Oxtt+9GJGIHRgSzUkC6x3SimpVfKFIdw4/E
68qdjvoP0zLcaZjGNUscWAgJ64yCBn0eP/JxDl0+WKSCwETGBoQt9TJUUMyPErohM4CTy1ZNCq+C
aMgwjni+BNVhutr7oL2q0JxModXLuZBkBUmSew71JqJ76QA8iA3ko55OZY3OUXqCBnpeCI+V9ytY
+2LbCuQ8+3fiys5YJPd6NEk3msK4R/sVTzg5N+Ijb3HVOolA8i701ZQTLJSPrVCj5Qckr69N3Smn
TlDqm0Ic4O0/k09c0thrr4RYUAa740wbbbPOkb9SwQmF+tvMEDkxOOn4Uw/tIFUcBvG0+YhqB/2m
fdTik/NIP0zhsgPQpA7SjEWmWcq1pXf/LkyRVRyTHkyhmFxceXPxblgYRECKcQuWQ0JypEVSIuHh
/vgmdtelazEKTzSUmk9j/SEHm+xM4HKMrObMT4ndB1vMEhgeKxSm6SMdyB8eWxpLYQtIzugCw9Sz
xyLjPtkc+BE/sCqs5N/hX1OSShRHgb2bG9mlTI6nL/KSuckSuakmaRpWqQt+0oa37Mh0ehgpxlLL
Vpff8cc2ez3kppglnBfgHzAMwysan+tzGH7LHuhKLdhxPNpeE7wri0YlvMv+tXs2tgZ6fw0sGMEx
ev+VaALf5lPX5+BglDRTQqKTXc5ACQXN28ZL1wdqW9zjV9dSkIrkNqF+hhuoCN33ootoKqsFxx0H
fALK0XtHDVGjv630h9jGNn9kjckxHvRZOChNLsdC/2lWzCtSRhSTkRR++4o0oUoV2lmLE/9Yi0Pp
ni3EuvygiWgW1Mq1WTatnH9tX6NMYNJhRW/mDo5ED4+2B8W+WzEnMiRDdr6xZu8zSK11K7pjTt4b
Rzdvp90sEjvyY8j0oWYdm6JUZrFLoRedNLXheFhCN/YA35nsaKr6kxfK7k2W7sAYYpj46aTHi3H/
XyQ81IzCMkOo4vTsN64jZspnf0wFJhcU8sacftLOIo+NfZcEsH32n/I6bha4X+EQ1AJ5V1DH/Stb
q6TaDeGGEBoySDZsbNJQEerRNuPr4XJns6rhBs/Ar68QcVCY3T3q/V48itBnHn8HbYqXeSi2v15B
4MmiVMo0NRYhfcIBy6RoNeazbGYMJU8h7k/bSmoDOWXfqOtOOOktACTohHIblzE4qplWBCJl9Qb+
Or5l2VrWH7TPLzNY8kmVldGx2n4vQOlc4kR8z1Ct9v8fdyU3wXS0/RFp340o0SYqnHGthwslfcR/
U19DUJ5KWa+panrJK1gIgGI5SVeX/I/q2xMP+eABqqSvtRR8AnnZRQwMI7plqUMpaDoI0uLpVki0
AO3jCxoJbKBXJYVcg0d0/5INuJI1lTKAGHq3XDfchzmCef22wUp+1X3MPFr7h41BEl8bNbssFJcf
F4MyRCsI7YPYPXppPaG03py36cyiJgPpo9mDhqUhjyN+v4uPUV6UcstQQ7V/48XQKavJq1iG1Wex
0l0JMpJuVDTOv23knVA5nX1hS36Yc6X3Xo3C/GEATB3nvK/lIS2Wze/0tEKj2ASN4+o3UWq5l2QA
slDkSsKEIYyceEK8UPExlYMw0qN0qxK3BZ8zGvu2LFR6nJMrkAa7vGBiM3svMkcfMc90Lc4CAW86
sDEk1hiwINlknHtFnA2deYrMODQgrz03oIB5G7btSg1e8oLQucVCG0RevETEdQ0jUHD0i8MYsocw
NHP/aMPY2t3kM9m7v5hapA+MuC8lbckprrjKxsrINjovld/7dhJ3OOGyHc37wX4v+1TmqCmoDbiE
yjD8V7C5eOwPAgBHo16R0xXQCLCskqfM1eoriYrG24xAQY2/l6ccxoc2tsugYhbd6JVn/bMwgSxN
QV88cYiNfG46RtTvjo8tr2UXG5KA8hKm+LlAqTSZYSAW8uikvnMDpPCIzbo2Gq2yax4OIpAUWWZh
//1aYWPaJ1TabX/yEUhghK4YCIfJqVhcp73LF+ibjtVazjxmcJqw6dcAlnrpWEojYGsiLKHSQOrW
3NamFRrat+ybFzSg1Y6G5oOUTxcLi4Nj/R+odC684xCwFIAtzyoO2Tn6KMqnvDNkWI1FwA58/Pt8
lRXIxIfdIdqHT+tA5E/OwkCAJVpiW7swEnF6Ti6cWHqNIHVZA2tbY5ELq1YZuGTmGpbwwx1LTOiK
fBxGyUz58mu6X07af4zvfbV0Ai87yqhpaS0DozZQU/6d5QleuAW1Vf3z+Kzy0g2JoZpEoZ5ez43i
ZCL3/1Y0Z1xVmyTk+no59+OwqTcgpZz7KB1NaIDNolmGH+PGZFOPikMC/t3mjNWuWl750xq2V8Qe
d8AWa0cz0spQFaUPYvRVPpf0/ENRGln8yd6aA/NaE59z/to6XVB7EGdHLg4IgGQ4k3wxApC33+Mf
t+WMz0/iELfBQCjFG4Tk4WMeEGVQ+KgU3ZSl9dq2uTfJbYBgUQ+In57KV1qPbCp3bROt8mVVp98q
rcsVsrSYuwW9IRET3DVk3IaRC8oxehbyLNQqke5H5seWpemgIGlpLZSoua74jSVaWqa9V/FO13vS
fKZ1K1nZQGv7oU+rqtGoK6X36XX28VxduC8/cauJjfo4g24PbJB7JlZNAN3abEuuj8tKCbgTgiJu
G7gN95zKvR8wKlqU+NrfseZYwu0FuE3WtXNyIhXxpm5VFShpsb5i8deFXziijAGOltQuWvQ4xc7G
X6JzcRDsJGqXDFkaJ2gk1Vu76kSIRsQ2ikxKcYjg6wzfnX7kV+2AsebSVidGMk4BubSPJyjdMmzK
jpKxIE4lB7jcW3wWUF6scjkCMXqL59XudcN43fd14vCU2K8oQFw83BED4IwYd6RrBs+AHsiKfqj2
NaarP5oAGO0RjD55r0UyWpSevhSg5DzuAxvZWiI2DWQB7DGRcqSzB+wp0EI05fxALI3tkhYT9srO
OxEHfzpZI4pHyDcycHTKfs1qGs+4bdD2mcOyUuVVMHBkJlKVNhFskfk8GBuxd70leVFlNCjoA1ag
19rV428LCOgEVJd/+CcVWLaWtMhp9AuABWe4prQVlwFdYctxuaFvygc4ASQszW4MKecDSroDHAR2
4MoPxkS6T1viRnbxn01YKWkmmLQxvvKiROi+FODtMqAbRgW9F8tzeC4kLYlpiqenLLSWVnEL5r+l
V93JYg4vetYnUbEt9vlfwlYoPpj2k35cd74mZZwToq5UvwIR7ig8BarLO8IGvGS0vF4AguFrCfI0
BfI3R8WDPaKZFTNpJMxlncfigHk4jxnvDhrbI50D0k5vq/k6Cj6L/G5ckNicjAfCHJyQ/EC1YwCE
KZWLtPxWeidGYT0fj/Sxx3ulTIdkt5TvvQ7w0Hhj+SDbmpE9SFWhJHDMOkytFEJkTwvCjVV9cXQQ
3JunExG6KwzuYe1uNgKRw0vgYjnM5vysTkpT/UIJoF54Kaux4d5FeJGkEnX5Z0Ks4vT0w+oebdCJ
o8gyMNk2t5y/rqEpW+SUd+a1XcfoDeIw/6BY3IuLwpy1Uipfm75YNNO8ToNrbLdzXbjrni9xfipO
DGbqbx5JBaGWwLWc9H9anS+941ZOPKVlgRfwHDTGi58zsxidLF+Sz0NuLo8jCL1MFm5RxqM1S/qs
rvuGuHIpNK19yYIJCdO9uSyzhJ5xqwKnb69jfAV7701Jx2ntG6NMuX77tai49B1ZclnldddFojy3
GEoB84zVsVRxOIZUXTVAcTyzjX7/wQ7zyDuyFq2NHDOnfWxXxsKaOjX9ETfyquqFByXKdzeaF+0n
peVVjdRrLQt6YoNRc5/DW0dVzkGD4TKW+4VxgUF8f0MwdQ8tdO67SnLOphjBit3YYOpDJBk8JSPd
1+MzaJmCEqN/d2msk1ew/JbKjiefPOxus0TjvMLABczF8iq/LAP3Ce/8dKqJDEGZl0LS8mJO4RjP
qd8ebUsepRhGB68reaiD1TIu4rqT63qyGo7zcC+O/krtdX1pfywSLBs9bmdTb02Y7lDgP0rsfpq6
HmKjchrg8l51HutYM5jnfCyNIS+BEGu9l5rNzgz4DesZ1PwgY38LpLoLB52IaEtXh8TMItWIiPPb
4IXencCf8fz7lHoU2EVdKivsH33ZL2Y+F2e+huvSw+ZZIcH+cDYbFst7MF3Mm+yQp0quJrg7orTB
gXDiPzNOX5WTSZGqRb7Z/9rFDNwv+Ar1jkspt/8OfXtw1HBgVV8WI93nTnghxa7D3UIq5eInL4TS
lPcGrFkgxN+ufhxxQXnABoHvtgW2Nf8EfvPHz9AJqyDMBfNoAewVCY6UKTzNH8S3WycqJAYtJnHy
QfsF501P15CiWfGPBv9ayFohC7IctsJ3ug9doDk1nH4kyHoTvGBTs2wDyF+eJ6N2lMIYnxY374Ba
Wv8tc/poAppAK631jzq8GongVJ3Q+G5O05lILUzb1/RpfHpCwYQf6XFDkdXHD1ySA9q1AhSOckNs
i3OsGw8UF6YmlWm+t9DYnIQvMvBG25XYcK1rEP0ehcUWFxXi1SYfzmFTYQ9acLcu2c5zXX7zW8fM
eoUNwtDDX2rJOKcygWrvWECgZ0vq6q1kL67QA88M+eNdW96aNUjlL7wq0q9J2ksTFx32rgEp50QZ
DZAShyjLA6IcHsXPTlpaPnpPOtcMQ0YHDFgMg17NS2JUGPM5dCDJEzfLIH5DU1RIrZACxw+Bt9BP
7IUFDa/eOFKCHjiARGSyms30J372mAAQUo5/kmlDpviQUns5YlRM58fQ2VG16uanz0YupQv7gEql
4inGgMj3GOsk9WP+Ok0qHuYgecQcFIZjmXe5hldwZXWEZG8u67E5BxJARoP2UbKpUwfe7YWNcdDB
b+C/PFRg1WPb6Nj3qQpopZXRLkvgS0iwvsNUf2p+hfGmkFnmgEWww4f/9yylUKANAxxp2LBv1OJd
9dixlPAJYQ1puG1mSJpokzxbaUmLPV1/VBUDZA8Re3fcAYdMKoCIxxI4EAivVLau7qt7fFTBCYlS
EiCs1DSg9C0JiqIemFNP5B1Dsbixm2qYUcws+VcF21y1VCzoMo7Z0kIAgf2cQvm2qEuQq8MBnPph
2oouWe9HOGy5XKHSMtV9NGCGVb+yzvU6rgZsyChxtVuirNHby4V5rKFaGbJgB1JX91OFmDp6PU9T
mH8nBn8uETinMu3YHMEhruXcGh0PWWNQ3Nam/3VsCkQ94YUn44kIuYzENBxHD4elK/rUd1VkKQBi
rxMJuI5+j4LOLceVRBNXPGmN5b5DjDDhsi+GBD8lFavMX82J9fHMUSI7PgRRiyLls/n1uAxeplky
dk9Zq7qXciHhM5XLyfJH2eFd3Ny4SwFhGjLcTDReLydgfIQ2nYqq6crR1c1ST+xjESOfPNstgG4z
4WB96MMJvApiZBz2NqhIAv+/dlV+ZQIYwckcH/+jx19tJ7DBb189DJercpb0zASjS+Fa6NGHmAWO
DgyWALuUe6vKc6YuJONLgQzuY02RFMn9MbY1mQuU8fMvMGukaHSpliY3x26UYl/NTWFP55LVQyat
5hbecT+lH+i+Y05RsXo5lb6bsXQHTs2RCJBnxvw0niydYWGvRU3yoaY+RzqUyPX06xlTeiKY8j/H
/r3rAg+h5C+H/CTd/emBnOsa6NUI3vWo6RGavRZBkPyZFvBiXJl86vee/OJtOMOfiZP/+0I5Yb+P
OdeYhND4nXOKvycPiuOzW9ydUZ2yVd/TI6ehN/WtAFLt6UZVxBcoXc5hVAyySWVjOls9JVeSuIeD
h6QEe+prscmE0P/HQkoJgNj5jr1aB3/W0UfoHGlCgVivAz1WU/D+zTJSnZMxpKahoIlAzVNreV4t
FSUW9msSpcnKOurbO+yNgGgwvmuFS+YUF0R6eH7O6hy4Se9tqueltrZTP3k1BDIbzdjGIDdQpmeI
VuXgodCYUhZ/bi1u986ONvZN3ceJbbKhUJ8dXr7pUhXRvqZ+jOtCsJ7umEaHFLKD9rwxV5JkRj09
ldLRNcFQpxeo4Q2fha5TIAjbHmKLQJLzNBku2ZMQ8ImrEmuF8fz5u5B0wQebx+Kv22dqBFsQfDoe
Mi3oZ7HEbVZkSDRXSDQCGE5kw5Z7Y9HtvCsYdu4kM3DQvQPCkzyAXJNF+keRLIaCWtsOGy7FlBfy
FCcWC5ryQSFweF1FC+innuZKll9Y7OSKDogh7FglAV60y1OCAP86qpIaHf0McR/NpFxqwrJPKY8x
JewBz/qtKDOOT5Sx3Kvl6MHXRBEbnuXU2N5WBW6gAnHOk5R0cyp3NRI/vJ4IvPO5lUT8Z6fr8/mv
Z9xj0PRUvsuwEhzt8J+wTX2jwIgKj5VC2xsIciizO1M5fCVa17/9mwuaqelCmqU3oah5Nu7YvsbD
e3BUg5CZZqyIfEL8IKM3LSltASd/qQ42r0TzWN3VpQBp97rpjWf/lWYZbUqUSj6IWS0Ea3sjhNAe
SQ4FqE5uzA8xYWJ/aoMMfTDUmj6ZSjqarN8Rs3LOXRulTHnftA51uDpIVtjrDO1XlbJiWSByMrJ5
g16jLh1Ko4PCk9AD09Ry3FTxNDP4Vr1VbfLG0fZzMCYk8KN0CbAoLTNphbZtfdjGS2lqCZLX9BXe
PhIgYQb6u6zbcIwF3MbL0h2moAU8bPmLCMuCh5ufQqdh35Dwx1NWJ/6K2P1O4/o16wgKXr+7Y9Gu
BiA9KGCmXKD/LQ5FjkBriBUkhGB267EzBuN9FvLHM+wjfF00bk4EotUFSqYP1LriiA7Sfqnx1XxH
eIItc+fwcLG+6MUB/TBhwC82m5ddUVCOi31zUSP/1K1HXJWUyc/sc1rQ+oA/hArW3hco5RWfrOw9
2aFrSj46GHJICgYVPB3oGuM8NN63WY1YD4ocO3f+KteEh0IR7UcTGEIe4afpEHmSAC0YBfJ2HnGg
vvTwKPXpez9y2V28WvhtAYGfVi0tbG8Io8qBKTN5ZCXGUKZskuPGTei8iEbyxC2Zfwf0tUSceGm1
Is8WA8U3uSdfe+/+cw+xsKQlEfTFOmKDF0+CSprHWsMDuOm3GA5OPidSNV4Hgbm3kg/hkONOHdC5
Ca9Lk75cZvnCIgvepRgvx5qYNBby7waZHOSpseMGETj3fz3lubmw4P1j4GmuFgDth2ggGrfd0B+i
G+8Q5A2tTZJCYbjwzB4NiUu0FfVhGOLdPiIWWd54a9EEU2+CYcRzo+5gWTj++g89uF8hlRC3ec4G
iSJbrNIFutyXvnlYagG4my6QeKNPoYwvrFEkA0+Gm/sinRCi//xxNwZ2Snb//380PeJWjV3edZFl
P93qAW8h1htzAFA+UJdG/MR/VZfPNWdXpGkrrQuYchy+RC3YGCIaa8rodMQW8uq9C1njBfh2h4Lu
j/CeHyt2BOtLusP2wORVm5WupntQpLXc5Fb8BHD3pTTgtbqsapjNeQUOT/wISis0VQ4hgs/tosh6
3icsJjWoIeKwXyHqUwcclRhfQeGUF0s6t9GWq2MqWaqBFA+jAwRXrvmGcRd/j9vHtt68kcPZg2ZI
YhIZUOyIKVTvw1WxiLfIzH3kAE04DeYalKpNVUWkxy9xILfnTxAOf+m2PvDabN5tYCvxNExEnm2S
qfsN7s+IpNTbGnixt8iL8OCPfzL8lHZtz9GsbB6qfMpvJA0BgSk4DCbCSnKEVs10sNuExhaKHaK7
YxXa1sIPsrVP30Q350BxvJMNdI2EwnHA5Q1mZREYEhZKzpthKqvJjHkYCdP2BZGLASlRm621TCQn
/+emDtbwj9NJD+C6fTFKGeyswNra3D2+FVlBOclfATjr73m3TEpiO4xcPXTaXQxn5pKx755Af23T
+5TTnDphrIvxvZiDkjNMp6gIJpg68gB5drE+6dVCPrCwbkfncADPZ5ssWu3BVsaTa7R5MZk1jorW
rko71e1+cPFymQDHhfZqKavSV6DZ3oUY0PpjbcyXX+b/N2vMZ/SVuKz0ULODIEo2b8uBIcrHInIg
92gdy+1UpSqBREGnwhh+VsR+jJZZI3E681tEtNFp26wIl2hQMHWN+2TyppvYBRhQrjKV/qxaAq2z
EjcKOuXd6YpAJoZYIkLtBS1qt2OprMWtwwaZ3kp7M2TCXoYqRzG5s7H13NDqsTyD6flZl23QcMSV
luqyhmelQFbhX3YxOAhHFNc6DgzzoNFVc4Gx38083YMpmI9zLy4vo/VN1ycQufkgSPPshduieMaZ
q/jzYLmzwHKCsLllx4w6IXrGh8W6HS6TwQ9xVUDx8SEISi81nYjq3n4gyASF3qXsLL/DpjtjEi8v
5a3CD6uurupN64RhyPMLfRnmCgSuOkO42jzQnQnB093RTvZSQP34Zw79p3CwNN0NsVQRZlE5YQL1
5tt7mJbJ1YiZKKbwfXzchG41XMq/rQ4u/lh/y8lMa/CQAHLqd+7BnpRyB6/vX00X/CV9R7Z6U1CP
YlZCPzi9Z/4GAYRjfcKP7XCWWPJblk43Nfaffq64cU2J8ONTc5T4uVYtn2XrmGBlKlbrHzffmiJ5
uF+L7lbIs/qx7B5RZF0HpefgW1ArSD57FAYKhF3rLn1jtDc62E3Mj1dGsox7vNZwPTcCrFwFYYVl
RtWhwgVp+n7Wa3xms0cJ1SKfTBvwDylSZ+Ooy5Y65MNWa3woz36oyMlSYVbOAHYvC1PRywOZGDxo
7mltMoXWgVOria4li5RkK5IeOjSsbWvLwmKJOZ4kPHgAvrgkVA6LM+OpBWmbpdSkG43DwYosFJdq
zy6onGDqCKLOCcOGevGgtZ9WUGiPOaEsXwwtQauPKiQO7qGRW4k/f/Z14j9nW8Y6gfPTuO//7rJs
gBZtrCBoKIFVEfzzlce0ybB2qcUCGt7reGMe3fjjloA9utlyAIjKIRwc+/+IdohZHxtwH+d1JJyz
Av7yWRk2O6/cza10hBI2PrlixPLLMJPXTLyqh+fmV7n0Ui+lmRBwJAjhmjzKQ+Lu/dFAtnCc+Gc4
6fp7cYM7SlHxnOqbX4qfx8NAfM+uXQ7cUPVvWOPeozod40UpQufWbt05TbzDSA+K4qkDUIl2z2YT
GIWuenpf0SyplIT8xM1FKS8I/2FbfxtAs18K2rdM8xxKIsfiiNQzYAFHDxWw+Uv6xQ8TAALDtKym
UFZhi4PaHMLCheAtz0cpQwS+h/dU2ZmGUAJMjYJZVPSkG3aj+FhPa0BxGhP49psqJ/yFokW0X7g6
zL6dak0ne13B3yK4/0yyc7fVfNpy52SPgIWtdIU9aFJ8UmwVHfHeCAifxXNBTrHbEWn67Rp+GU4w
KHlBUKmf4EuuZY+HsPd37QpCGjSTsZrM3B5Xx5AZ3Ni1AcCFDxRz+U9g+TDYSOmCtiC86xku83Jv
DxXcV5WZw5ATi+fv6D9AnmvL78ggUij1p0GdlEsx0eeXSudDQQFmRWy5x+jDYSEpkdf7DsX+b91r
iKKRceDDaL5sA+OUAiUcBL7bL3EHSmWavNboPkYE8ynlz+vxRg7hGMpLLYVBqdnZAcgiUzygWhaV
T9ENOr/+OwRxzxk5DArkVyH9zRn99RZae9cO0ot/T8fCrrobRv9tIhl+jeSZikZPGk5ytqoqygJi
kZwGrOC1WUs1S7GX2gVJcAnFEbbW0ukkm3KnU5uVMkgHIOnNd4Oo1jawxFSn8CMhxlwYtZD/cOZf
AdjjsFPlB89d8LEFcclJilsJvh/4CNJ+hG88ZpFbOy4o4ly+V58y0dkc+0qCtxbADeZPlmsfHX/C
KDV5qqUAUHTT0l1215HLvrYwGDpN2qHit3eg0LRt5xCKZpZFmicDLg/PDfgGrnlSU93Afts5qfEv
4oZfhs06mWeu+VPCs7qxHtKx24XewHxpzoDonv8KGp7EzSPGqG3gb1gevrx0EqZ6z7P/FiHq2sqE
rzwAY5fBCTrlUw99qnVHsWvh8T+kfTiPR10aTppGq2CXxOC0PZWhaFevTpy5NpZoZM/fj6naRre+
8VYmlNToIKgb6CS500RPNu6bJR1z3gPSueyteP+0BKINJEqsP3Jld2kJCLwXiVtuP/Fq74HHx9k/
GGH1d2FFlsdlLjwJl5O9pjVyVU6zG+X2PlA8TYWvaWN5IJqTg592B7dgPgEV+N4REc0EIqu+b5pv
JbMLxQalfKJR2PwUfoNV9S3zebQ4WdPvP4GsLgAcIb5XUzIO/OxCQXIn2hRrAmo/NU/vFzG4xB8W
6jI8lwWFnW8ZxyVnlcU6rmnFMZA0caqRrqNCu31lGzsKl9Q4Nd/LWh1+pPBztB38beDrjXLpHAQC
Qrq7sYYV/iJLIcyE2ltRAtDB6ZJNwC4Em8QmksyWs7GfwRk9q3d32ojBApqHxZCR3uvm1UbAGOYZ
3Q95IMnbCCUTudVpCASoG544gam9vrfadtqxj5qU57NRkPM207X0G/rH1A9ETL9zgBncRP0Kt+7Q
krd2rUTngspyxPPSXE1JDI0XMR5H/d88XvX5hPAh1OkZsia7XMu9xJlKShk+TPA+LIZNgTvS/6+L
6Mx4BsxfMc+4SVN+HqlxHfVIUIsxeXQNKn5P+Tch0OjkntfTVj25jCR0ubExrPJ9LqV0umuTJXAK
H9q3j3f7dvemT3++KPg+m91R5zmdu1o5RifgBXcqqlsQ5ZiRp3vlHQw+nFG8WCs4RxyQRAHb9xnL
NlTw5riqKzTRafvodZBetX01LlmofMQ65klGls1yYlMP0OkngnSwdslD7QvEtmc+MHHha1oQHDDo
W4y6bO8qEXLMiMyNECfyzi4IO+KkK+NuqWwEjITjovrAPxxU5/kLau+n49s2spMeVledeCftfdDN
0H9jZqWbt9r5/kcK9QH8otd7F0txMpjUUJ/SyREiz6Mqpnc3De+7SJOh2Rxr/b76BeqUS/O8avJc
qVhDnl0ydOFYyTYUO7TdWCwgIc1YlDoPJJLzqzblbFYKsPtnWDZiwS8yNL9bdAwdIAsHOz5zOs3Y
ikXArpTqDZ6XBGtqfdhYCyiPi14Xo3HYdwN4JcxBp6ZBaHWvd8H+fgcxEdtq1MmOEwE7gcTxj/Cm
cwQ9AnJzILOnY323Xpo2ajBaw2QFiUpBDcdwmqf7gcahbY4xK9KyEmD2DxQUVGOXNAg0eAbWkpfc
nsJ1NJeZN7I3HtJRDbhkEk+Gq5oV0ZmEwMuUcj3UsMbx27+UqY4uLIkCDLHyQhBsiJXxbGxm0M55
iJKLVYZDfXwALN++U7Qnk2HDWC0W+39aQRwJAf3eLgo/XpJsVVc0Fi52+4NQz/4fLDgaXVwYA1fC
y9cKGEf2TF/CJqowGya+E1p6q1n0q1XR0bCyrYGwjLblprat3tD7M2KlTB2EQPXezMxKNwa9/biN
sbVzQ+4RFbx7XX0lFNDL0P+ygOM0lUzjByVB4SWxjPfvGM3HPuwU49LorBk39dIMI8rRT/nnikLR
Ua106SGokdphy9m5sXRv+sxrfU400J78p/Fr4m1thmkFi+j+pjOAVDDgC9/mlWoC2iHQuBbusS/l
xc9N9aJqVt8mmwoSBdH3OOG8DO2/cK+cChecNpwWBcXbieVr/hXklx48gcIt1iKngWvsQXoyykdi
joHN5pLZ2djQvFrmlCr8cjsPOwPBJ5VcwCllPk24/3gBT3ubTbbk3IuNoNJEQoXCD4eTfCsLevv9
M4ucVCioyZKlbuSUOuQrkKgcCQBJMJ5RHBEvU+bRJrJkOoy9kgsuF6gAO594VKVzhTH9QSrbl6Pu
/GKA2ZHL8QuZeVuunrP3WJkYqLJ29bhfz2OUn29UbJJlLDD4gHRLM2erLJmXes3NZlVHl6DZa66q
ieFzuEAPE8EMrky4A5IXdKpOu3Tca2XxZFvVYwkXz54KqEaXLGflTRvhm8kndnR/P7yfFEE+gKau
/f+1ZpRejGP9X0oePfqCGV6PCuUeIndMxq1ziW9X49vFYmIdJ6gNCgIHYu6YJhcqYryGRsaGz4a9
0ajtwSmmb+JBbJzpBy9BENFtmqHbiU/NerKfwdOBa4cFpYmgyRfWnQfvqESVBNeJ4BLAMEFwnzPA
+fc4eew7z0A3T0FIzRzrl2gsH3YS2+kUNt+187hJ9GHklC8TNJtfo5VZvB0QUneOxmaE6FX+Iyor
h7uOvv9XIkvSZc9wUgWqo3zXZvgkh6wWmejHLT+6mfoLcfjjkO/BAq6JDQuTrynimnlBjzLLvpiI
OiHy6muOc+HIRCwu7Pxiv1qWud4+tY1Yx8NVbzVMcGHJNFqfqVgVKQJM0guXPhrIFZaJdfBmMVXo
SCen5TjokF7+Ld9lwaus+1nmPjOiN/0hfySYDcovN2WhuP5jKQ49m1xEogvk0kwjXK8GnD4Mwqxw
W0s3FZKSpXYtdoDRGJi0biGMSlvtSUh+wX5n8x2zoUfnKc+JCNfSaypqe6ffeLO/8zqkD/KbKTsk
ifBj0h0dXkKQd3La0C1+1EpIWdPWytSMDFfr1jNAI/I8te7E688phQB+I/W+Poj6ifxUDa3cKWo7
sehaBbIFEcicOmwc4O941nf/saYFtO0ykGlwp81HSluY8sR8UvrTr7UQr6inq6nscfihGy0x0TcB
CxzQZhq8fUUWxyayTyAUJZiLQXv6JaO1+7umF8olglz0KZaT0hp14QTup3WRfz1ALtKXOIVuW0bT
sVUMWozsu1oQYMyaIvKptKxdVX7+cbyO/QpGLWvCSfHj+v5cbOXifRgaW1i/xtj+dXlN7Uoqlekh
PfaG/lmPRwNSN5GOdZ6Uqbkvt64kwzB7tby3s/IPMrU2wyKzuhj0N9hl/0t7UOaB9yGZejGVcwrP
GQwqEnnoGiHCaqp8jhzf7PmzNiBEWu4zba40IL9PWFsNsX9j/YM6+aBTV7ugX/lGvtMdfl9FR0B9
L/2i1Q6aObufl1dUfp6a57XnxdRq6akWRvSbiIXj47d62YYoI/O/9cBdHBL7D8L3tC1x97zt89F2
NKuGREirjForqBprKWjI51+evEbcHfXD25c2v8Zah94ePlW2DOU8o5Cq5ta5psss3eDZrUQu1nlN
cK8JpAmCnlaxibhR8BEISWiLcDkv1B6l9VTKc7LFel9ucIZqxkmaI0AlgCz+J9YaHG3YsdH2CSwQ
v0906HM4UX4DsjIHQ583vwkiiNuaHKhVFa3hWJe4vHLZ6rpMwCqQUfnXUPHkWDaBvN0MKvPD+ZDW
jYa61s1kiaylrdPfhMw24WhqNe2K1drTvCDoWxY2g6WV5yDZuOahHXcMm1Oqkpd+/iqKNeE46D2C
VUjubtTcJpmHdfTok+SstZZdJojs5yTpx/wLOnXUglb3TLkO1blJ4Vil4Rn/B4f5iZrqh9yJCQVn
90pio5X402lir55tiLsaPm3UFz7Mh9JX0ghsreVnwD3GBvTOlSDKBCS33lQIydnEtX3V5xKaZELT
aV8MTdLN68d3LIOW9Zrb9GhHCjCuwUiZqzADtR/IDwJHMQTqFMcMj89UhtwTx23732QDYyo4Fj24
Knh5si2nJ3/qlbFO3mol1nVLiNG4n8fC0L3/ATz5tB1WMJdrIYwZSFz4X6YRjy+LGcif7F04Ku9m
UrU+C49qVPx2c3hUPF0LZCBxqe4KkIEgF0zosEWNQEUmjCNn2AGwI+aIObC7SYWlVJv0y268ol37
1xRTsjZZLv4llxGF4MEgTfx7zXJz7raOhyG69GxKyWCvMPvD9UKdRSX7pMsOrfr41OBNJ8ak201g
lgNBBaUHd4PeyX9qRgLWkWzPtjF2Ci8lEctSs/0Gwkliy07PltlMmgHITd/H1wemcIHYkwWFRoMc
tRxGynPre9dhJxUlX2EgU7EoZfs+OHXm0H9s0KNWDtwK9OwB1d7xVFTG39RGD4oYrSXr5AFNNI45
vHyYVfi8b1nBaAm2NK5gZ0pXD1+zMFy9/ZF3JG+tR/3rztj58qSVkkR6F5vnAA0vZFoE1gGiwniJ
X5rhmSmHzMhuCKVQ8RF9lme5ooE/NmyYwMVLkBtQYNr0ATpQTn334U3AIdq49N9UsMovY2258I60
b8le/6SeLox029lt8zYAR2HZVUmIZtpcLzDkBEDeui8pDWzAg05pjHLw45c1Sze/24UW6e4klLCr
EiH5GK5AtSU9VC9WFls1pyOLZ/2Oe9YHtKOqdaRyaGl292cUIRXu9dEmb6nQCAOaM2A81qxuIzUN
DTUTLowdURlkHrIxunw1srcdU3UQfqkklxaCrcZKMI8hEf1YED4g8ar+Zhv5OgypKzLivCKMS3sl
Ak9k504jyhCdyz1eRdLg/YvZTn22FFgEIDqDA3YV4MXW/Lu/Dy+S3QGLphNyzHMd+AFU6EXzZdrH
1zpeI2gP6xjrolg9+7wmI1pG+zlAF8+b9gm+KTgdrHBJDOXHld9BgUvZm6lKoZIilYf8/+XQ3vdk
kenrslsP4QUtYYKIfuuYbj19d6RevA20XeqdgPIM8vmOz5b69DAqcsHObLOUyfGntd3CYNJgFdlU
MQ9K+d+WzQRM9vr+YIsaU2sN9CB0EEotprQyEz67Eu+Bx5IH6irqfY1t1Xc17rKhx/gFUhdckMMO
ESYNzV+9C2PvG5txe+Q5PmmBgB0hW3EskrVpBIVvcIqNViytLMMLi3D17ky/0EFEdedQ5WRBCitk
wD4ikLrEADTgAhOnc/1lTPn5i9lOgLLidG2K1S6WwMHKVs2ZSaJkT6NdBpB+bB37jg7ycaNmMIIT
fUFZmh8Iai0iHK1fTfD3JTtb9xdo0/MjDcjVbXI/3ToulZnH44RMjoaCMB4huXSrhyDjTVLNnqK+
70qoQDLQ/A8VOYrEnnwmQKup/uxbtmJ+DHFYnRbcMmoTZ9DT2+lyJhGRot7Xp8Q1U1Lphkc3AI/f
TVK56O6JjUftGMozW1tfGu9LE0AWCKZIqdJr1uH9FZmpBq5l97XF8Fpq2XiNXR/GUYBeM1v3FRnR
fvkJiHLZxlsQrbnitNYe+up0dND4CRNk8DrfZ6v2B9FeglN6qOT1sq7COi9g3FcMeZWs8RYoOU/s
Lz8Gnbunm3LRgWQUzdLexOWYg5Q6Dmfy6nlTNv/nIoYBPqgRbqq0j+OyhjQ1NqVK3lapg4waPDM4
FwpBbqwPDoZt5oNP9iXfdl0XarcSjcrqtYsrpJQWWPYJhg3NhGteS8WBm8M9QA4DEoROc8+XItsM
HZbLp0Y/fMvtA9vAvyh/rvuD9/q0aHtZY4ae/HHFsvIudqs5fWwHXpx7dD3Aq+YhsNDn1nnFgoMa
gq75rY+Db5bdDxI2vLfrBrKT7nFL+kUDuzkUZVE/Ngfkk7l5xyDh/D3WEOeP8cJ8Ua8rF3M7SH7b
284tRK2vNR57FD3jo7kA81IZWrEmuAifBEsy6oDPY1UjNBSh9SMeiRHu+FGdMZJnO9jhlvkVSIBf
vnC0oN5umtwejgyaJfBzAxWPOPEXxZ6GwHQBiH+oHTnNfkWysg2CydodK7tUPHo3ADZT/BBfKtvs
CbuVCFE58Le3ZIaCUGYdCcFkZqfjnwGJ0bjW0V7Li6rcP/41Z6gqbF2w+dbnIYAeLW8bgwxfF0H3
Pray93mEsa7/p2mf4oK9EvzK1PQUe1ZtEwWZNdU7KMAljQbBLi+Og9JCbpFVoo7NtkEV9QCse69h
gF5y+a0ei2XMEKH0OR9bd76vFQtjnsFdTNB4BC+Z81LlloHoOaztJe6UKoOjlpKMmg48yiPvBHMs
hFrXejgM0ur/KdXDsdJTRsD4K+wMb9Cm4vu9ZyiKtRZBeYOUH70R7GzVNQm3pRIZLXPD0cXD5XJi
8gWYDD7pDqVJ8xUmc4Y1pRWKBGfZ14kGP13TzNRn16dn9JTVhurIa1MVs/ZK+0sjXhRB5l6wXTwR
wVkEfOTpq+5athTzo19JY218uP1s8WrtpZM9xZ72skqQRhtMslrViiAfI5Fb37D6gcAkRw+doucU
ggDU2CicwKOzq2+j9GZejCMZ+KSDgClaQ8wzO30T4ubD/Tq2W8358oX5meR8owlJW7olhV/pFV2Z
AIecgn9IHq0l+Lq21wCdDMFvhsz36oRMd2za93IQZ6i2VWYZVBJySRSn9Z99TtpCbjiIjqTyUGua
n4TndQMmU4Nq+Mzt5hn2DcULq9nnVHfxO5vQXtUJOY30oqGucxeSrZxWbOUngzH990dxQWO6H2c4
f0Pn3FzzSZBMsSyxC270k4xg64GAepjjAlWxUuQ07Muji3obcN0WOUIQ4/jJzLqROqusUblayosJ
cZ2Mewk6JnaOgjY1H/Hi5Bvxj/8DDh4vsHG3Pm6yLEwqmpC3pmDkAVDHN7d1GwlgaWrzI9xgRbtL
virH47uB4ZZFfmbLfidXUDjUeyojJj6VL3llfHUS29wIQWKX25U6/SanguGEyyjjVRIfrqhsSOV5
wDSYP1CPLpTVKlMARFJvoQPltR/N8mpAJc1m9hAP/K/XrZspvsh4Fl/HxZm73Rct1KcsvD/NfLLQ
2NcPBYvTriLylH5N5h57xhBeuxzx2Fw804BRUK8kbunboTttlVW9LO+wGfGfh1rPb99rbM5N4LE2
YBwPhKHeoo9SAgVlSyuHVa4UY81Irs5AMsRbYIQAB6hcwN08U9JrCO8EmRdOJVzRJ0Z7eYZ+tBo6
zBm3ytYR8XXvX1WNYwhVAzshfwfbz+IaPrW/AJ20enPgkrrYEhdwcWmhm90t36hsiBOvHUSCNNgJ
KcCb5ZWmKY51unxuul+lajCKJQ2D3OA6OoGkHJiQcd3ggN4EWVUyHp5dn3Idjt0EFAbHFGuTpWZW
+QSPLhYHNhqHW6JwEOn6t/wBMwrrak2yWNx1VHTOcbxrM4IwvEwULaA4z0XrfyGJ/oZ1dSDjNX0T
zb3hW16d4rzyebhqpcfw4OwkeSK0fTyObQHkMPQZUqQyi7xVU1RkETds9gdD3aF8h63PW1nZgb13
/kOF3LioIV+xWi5KA2zUAlm4UC+JiOd1jHkNCUks+s8AyFUK5M/t4zRDKIWNyQARxE2/MBEs6yHE
Pxy9BYv7OWmIpeimGpM3WmaMAgL5WANCzAqcBQVX/UewZVDjhte9CdC9+SIG9wQhquuVFgRZHq7q
crnUc0Hd60cedYfQIK56RlruTab/uiWlIRFPOvyPTD5ZSLVG5+UUTpJpbnaUZKVOZsWUSrGKAadu
HNhvkz7H86oW4vKjSsyfFetcJKPJLgmpqVe72rIJifrBkfHvG/iWzlLtjjmRkh43C0QrlgcZDXQF
WZ7ycqmn+ra79kLWWhQK8+cqcA1SnNvJnFzaveokGOVgZTd7Uohy+qZ1I2FI2jnd55XJ0BpAPXVi
2J75UHyi392HBJZBDaQA2pPsJ+X7kdFAKo/ywQKHQYiw5K1d95M94r3Wr5UrVXBofoaXEWLZaN9D
F/Xl76RnWEUX0vpY22/gmuhiSk97gOwCrpSpGMKd/3kb1cQY7aaW7NyPxsAzqFoGLO1gnTsvC8Km
GYEZPywLZ99m8onv9yRzDkCHFtz7i4XJFmMJlBg/Bx4xDCwYoAUPHp4OtOfRsZtDTODe0PFa+Zv7
194BJty1jncDnvJwoyKjKv7rvi0o2kTw6iKPKDtd0ssDS8K6zhOSuJfJ263hE8qTXvPBi6iJPz2y
Qcr/w4Ymcixj+Nw0OQRFhlHUUeabjdSb7rHWIKHAMLxUxuUxVo8tKvHkQFNAESCnCs347ws4SRsT
4vqdH9Ia03z1uWgvGA0y3WOvctFK1BeXNX8k392r4IXXe/Jx17odcqUxe1s9EeZGKhMqkiLSXC9M
3q7MwQKgAD9BJiM/rwwFaCcL6TFlrWgjqYdIqij8QJHo1jxZFbcFJLxNP04/h3JiHTVrVCQBsGuv
bq8N0l1G41foO3u4/cuzXlQ8LigOVwTa2KKYTWLJ2qaysPYNXc+rLiab0eDS5NQcHVW9cUVEx60N
fOF+6fL98kzMXZcK67dpfWuGbgnshsTPindmZRn4U3WGeF2Nujz310t2wK5MNZDQ0KLXz7neawDg
4ETt3ci+FDnGJ2l6rvTxWxHWGaz9FTdFPNTw+UiAT/rdrUreYNn30cQ+x7lW6s+e+k4CZyMDeLJL
KPhihwiZJjz0iRs3KomwjWruOsWQnoq1UupiacL7mQnCG4YV5o/92+wy5WTodQlPxAbcO+HdcYB4
2cqz2JeYD/0D+PYRMPE0srMHsKMYqvVo4iJ7oE+uGar7WewfZ8m8EMGutDieFULL9Nc3E2zKWlcw
vPTyiOgABx4qf57r25tvX3+NC7LC5dIqu7kK72q30jQn9CzsMHBssJTD6qrV+x9kffdDpmbFnVLm
qiVBfiKEJm43ueVq87USJPkptTTAd60Tq0ECu1lTNV7eQM/tLVDRO7+Fu9t+UkG8qeLbURmIJUSu
hj4XLhBjN2jTSkT9JeLfPKqWxX66444Q1c3h79WhA4OzpKMMSv7Cew0bXZXoFvFCN0zjYP4H3W01
MWZB5TKmcqS0+4nBhZDDhIzElKpgP04RKz4L7h1+45NObRC2rstlU8CDjiFqPCRrNbfHa8m4nOqp
ApNTDmuINSZZpT2Uphqs4NfZ3xAJRSjhuq/M8dEEcQ2hcLSgVRj0s7NEv9CvdQdOzvK98RfX6sqJ
QBq5ZcJg/MM+O3uGJOYoGONeyTjyGuTQpuT8zSVOXHoLALJvspTq2cBdBS9MLeYrIbvdULido0zD
D6Qr1bSDRhis8KmWSjutXcERmT87n1irUd8UjkdWGtt34kvRarETQguhfbxZu2oNgF2ecna/edFx
DutU4GZRCoMjvZJGITeRo+wUQTdmuQd9dMTHbSG35m4LUEWg+qI7cXTZ/l2Kpq+UELqyAMofCI5g
5a+aZXrF97hhXunL+D/aUhpKVDgDQtLZbVWFAEn8fCI+2IVvWUbhuLU3toxfKhPTdaBgwEVu2tZK
kWdW4zFHiQPk8kQHMpfXPspbAoQlAGdfd5/z5kdSTMnHLpu88U9VYy4FXuaTN9vPHVzd1s8shmOS
ZBsknYy2seLOp8bwefZOIzIxxVaUUBZluk/bIVIPmTKBipJ2b9sR5EvqOMREgxIQ1qE7fR6XoKCm
8yHNWnYzd7kx63Wg3UMxMmnFcSxP9/q3/I5CtYzxioMng9rY+gobuQnoRwiJ2wez7PvgYCjacaBF
v0VD3+me481N2OWXfuSKB4Co6cYxlVD+azmvPbLaxik8uzoAyEBg9FJAnatRTjBIoZJJ5nXdQIfI
GkVTUh0xmLP5Xq0MWLk/AU0U3ASsgU6HDnBR0BisdIYSmlgElZpJu5y4BYHVgGigco0T/SZ+nY6i
VQ9qp/IuGjaBDisg7Jl1+W87zD05u665g0GCSPXM/yopmAwkQQB7RxhSr5UvI+z7haGUOn5OQ1pT
eXn0OTIJmuyLUeCA1rWML1hUOqzhUMcIjNRqghBZJ77Vr4YH43iPUvrkQpbHTXD5hcJule1Yp2TB
9Dtr8J5gcAJZ7oxSaf4inGMt/nHZhlR9BSrrxsbQAvidyw0cM4TPITesCDAx7okY2X+UdPAP3A1K
qOOADaTfd2a2rbWWPyupwf6Px88MVmOoeHznfqElQuGK/zEDbCNpXmnwgMZ4B6fbpqy310bGybXs
RYQ4uO6DmR6hVvCMJa+WLKAt8hsiM2AsR9lpL6rd1hHb69PvJKCPyzoM7heZLVhytGvkUyEntDGA
fHdTzU46oUjFQ+RhqzNSL288Iwv1zgRftVEIIHB8CyrMUvyNbOV2Rw7G9TvJRZNgUyVzEe1k0s5W
pdVNSkddTUwV5j2J+e47eN5e05wKXzvvjj3bbYWHhJaCazpSpTcMEKrvaijTDPusvkkPNCS3Hber
WzWm7dvbyFbBsyqbluy6bvUsX7pPWybGh7v9uw4sBdhdFdrTmywH1ayIB2psEtIktTnpkEaE7cXv
7pzMJkLzi7/IvM4K+BLAyBgMoQpvzMrUBm4CYL98XQXEuRrvzYuqrW4pvHuWAu9lVorOQ9YCUKPE
2h2ggDpy1ghBrEUb6DqCxSYkpQPTOTzVAlQZbXMfaSR3iDsqWpM2li6jCme5PP5D4o5HjmzSaF14
lq+NV+afKxshx2/uPdhm5h7vOccelXf8wzuRsO+YTiMwodwmXcNePrfCJgo69kNYpWRVr9vJl7ZK
+CakaaFZxyYjyWFc2aqoKVHsWVf66ISDiIvneGRFtHzEEyOFe9ILGWCd+xevcv2bbpWxiW8309+L
dFT8nwF+UFHtTjRJz3+SkGkmEQng7q2/8wPZkIlgKWqy+7Ft7fTcqcR94TF+lJNEhxeJMG9jRIww
qkkpM/YCftyr0i9gZB0149EV7+l8MEAmGc7xmo5quDrv92rf1Kt4DUJR8lJR9IsgxjXcGTZEBVWt
dtOoSCu8LIBGQ55vg5P1K7aWkQQ8Jz+KWRR8PrNK8U24qGK70mhgVqNfzAGtw7FTqG8IcoL/U3OA
B/E+nKnOWz1fjPAqAJ/dWPXQVfmAxCGv9SKRBQ8OE2WKSbZriwBhJgr7tDiytK5lEvZ1pKordF2b
GayIU74EW8RcIwVBR0YUXaN6bxnBKdxXPNk4Uc/Beeh2f+X8KNwxdbGDI2xzruR4oYu4KRcVuRru
Wh+G+unRkaCtWO7Lk96/EEumBrcFvLvE+1l0zwDXZCiBBkOEpZnHm0FFaJOsGTQwfSC/6hc5oYWc
IEW4am5dXTWDfOuBT3I2QeSM1H0DSwr1ewfK34fqFgzCx991iXkX81m4A/nlQz6rO3NVhlSbmsZl
ngMo2jT723MN51Nj1hq72Lfn+3BDMuZ9ommNeMH+pwJbi0bvQgWSQps8F7LG9Lj9dwT2cbryTL6X
WuXdvVKhf69gAMbnz8C6qCAz4p5BJm3BnoN5T7O/T1l3kR9wusbOYh59tq+S4WjirA5wFwspuzUX
2QOzX5Gf7/uAOwLUhDWdj6NE+8bD7VGsx0y1wk0t1xN4qLzgZA+KX7nHLPwkV8lmY8VWEDfbr1la
lZnuBQngCax9ZT4h/US5Qruv2BnxB3brif3wOy2ecyKbVNXZX0wjsJkxDfFlCXRaO8WXN96CcGTe
nxTPdeAiozC1U1tRUDafp/dnOBKO4GxJSaMTCQq75j3VthCe8w56pcdkyFExa4k491Aqtin8D3VS
Fp84QNbCL8y8D7u+KdG5vhJswhkVvh2/wPSFVdU4eeua9Q9CWRTBnBUpRvuTEBZlNx7xUiM12lK0
hbSWPvCiEvhD+ihqsuuNN47ffiY9Sksska2YRTrezs64kqTP/1mYhNPsUQQgm79rU/42JuQV+pxA
Orm0W0+Gn6bjSHO3eo6Pl0ulxFlzGdaqWf+Cqb0/a8bum3M+BNW6z7KTqlOqbWGDkP2/UbY0lG13
fO/CRsYAml6AMW9l81ZhZcZT8f5E09Lyp8aK4KWQGIuh1GTgTk3OwRX1yBafXHGZ+Zrzq+/VGtK1
h/dL7ekrsFstI7afwLZEB7XpZzUIIGCEED4j0qqTEVbSnBzTKVqfja6syg+4jm0jiwihhY6Dtj8o
qXk3DQX8ZhvbWK9SYF1sd2HsFu5UOVwNqM+Rdzif8RCIyJj0uMYP3QlIHB4y6xE0ftFCyBZqzCXJ
8zVXks1VCVLbMUWdeQOtv3HX90WYuBc+LYE8LiIx0Hj5fvUlT5IafSNBTYC0dTNBXmqk8GqOeWNS
/C2pcbfM0TZDXLEOOO/FnZj26hiBxjztg68gJxuWC2GaYF59om2Rdk6DNatGu5nVF3E60MQx4q1x
wY0gyd3iJFePLIsyV5cbK149LyTUFrU88JzpKaRjcwRi5Bf4jciW4z6XpuhA4wyRucyVwy06Z1qj
DJqYea+aKVGi8UoC7DvCsTUKUGBUInBWrnLErnRqaMO6+JgC6M5yPxsTUHrRfWi3xTEQum8uIsQl
gf3EA6afjzgc2pUq05b1AMoLP3eodRvfJb1VtrYde8WX/wii+rQYFodm3QhEfTL9VJtX0uZR1hvF
4+baZ4PxzzgGEAgPdbaIpFAizn7RDIwUvbpXPdjdshTvHr/06V7paJ9SgWKwZfgXTa0tToi6SzNt
zc9MaGk5Qur1BGriUjeJOw2pnt1hYKDroclkQS6Qz4AtzDbo6pMsKWOMuxDztXuK/UKPYe31wOeC
rPQJcvvSJposPY3j3FTzDvIWSwxDzU5fLLL8VtLIhoD5F2UhK+Eg4q6189cXrH9wEdxoYFDfBGvt
JpUu3cI543Jt+30yzyxNri0+gyxWpPI5zOXG0x1A8ME/TR5dv+OyIO2CbteBOab8xUu+082EIt8t
sCT9soIBXqf/0IHiEel6a8nwMYxESaGMAOEX5emWvxfkMsPw/YncjS/6YVaK4ww4iiD7CQBgTqmg
ReyvGo4Ysuu7PfxhDT+0yvFXJgQSjyQ0HbyqkRxTzj2+DdKTsq8ntpkhHj5nQ8+MbADmaK72g4bb
n/towKdbVajEAxnYZL4LeZTKF4Jn+vhMswlKdXb8AqRmQ+Gcg9ij8CtAGfiIHM4/sF/68HEVDL3B
N8TgmhAfzgCS3GOtqKoWdUhKM6qm8U8CeuC8CfRPqI18qkTD6tUFaFsBzcKVEeSYMgRMDH3i4XXw
tdLwNvSAp/e6k0Gf2DJBzj4cd4d0FrNxbq4/0SqRofwCDgsioPkOGNIjCqd4exAZjfYwSQOxnhpb
c35a1/79K5gWtLdOnsTqulOBDMVcjiBoGbj5pS5thNPcwG31zqoSg5jYB4GVWVaOen5I39JbC4JD
WPhNFJi7YkecMxRtOzxsIsDYS34nhMV/TWofqiBRRs1/iztO6OvkzFmHxIfqYmf3VxVxWsg27u8d
fl5skkdqsLraXpLE/kbAwTEHZKJYs9NNCk3vWmqz/eKxtknkaWbbO9Zsavfvzty+jkvokQ+gSAZp
x3udUwrNNdLZLWQZxhPcPTRVX8MGxNt+H4CA7L/tJSwK987D1nEzpkUC2XuYHYkdvUemJCGYgMsI
FgL9IdK/d22EzqvNSU0TrmO64V+vHcZG3On/BQAoNQ7pDFrYrrpCVJSJmLFbTdv0B9iuA3PvpI8L
mtJHInQTsBzV7pxiykOSrFLn3/OBs6OrjAqLwqV1pjL9Ipttd6OAK/e6hDw3amleuUVqeqp4HqNY
TnH5fu0oQ23udA2pJ//bwRoeg1uXNtGWmlY0qYMqaeIsOczyykx4qZuFoDevc0xLXWlM/t7zMIKe
4pa6meXbKVMETvvWI2HIr0PqvB8h/rvtOddH7YoOryA8hu9zNQwShoAh/4wSW02C5e3Aysb0RGRg
YuanPftxtQ6AFGvKAdx9X0mAjTWtmwuNHhbgBg7eXrdbX/+w9+NiGV3N9rkCLS9gqOFk7FPC4zUs
Q85VXwUJe1wbfVzEgT8cVpbHFf1XOKu0HdRCnrdYLHdvdlzXkv3CKygmWyy7RoASaY1QfUzJisx/
3oFQIncY2YmH9S/yBWXH5u3k7i9osEq+io4DadqgdLW5aXmhBYPElF7LNaK5KsZv+4Q3SG1BvtCa
t2sEm70owK7rXTnCuvWxJo1PQXR3R7v40wJthEI6szoFONxKsGz8wgT/eFMbTq6WDGhDuwsz04id
BEJNA5ExKF21LKigY8J2ObelzSajAbXpMvUrOh5tB3uvNRDRDFLzauVwZCEkF6QICgTNby4Am6MI
ZYihOCBaKXn6vLuVANkFyJcN4EeR1TBD1oI1RJfzuuFJswbpgcCIOLrYwrRARnURIjC5WIjOBUBx
6oep0CZDcaj7pYDmD1p/zxnFHwnKXBAjyiYSC6AoeFyGj9yoCg5Rak37IOPmV5fNQOZUTeiY0lk2
SyUI/kfG3g43JGFMLQyOrboHaEoUp62TBF8Ov0qVF9xh7xsg9f7F/jnn9zAJN3Stb+oKSkguOHFX
9KcLkipy/8w6sui6Ej/6dCpVkHoVgdlJKXUhazVSeBzgCfR1ql6qQ6R8MZgmP6/m5FtDTtopeuQP
Uno795obgG76J/ZaqxbZvKGwLktuVw7hk3zeixu1WB31BDo9GxEWx1LXh8BouDkFouB1IkByaDTC
0b0V95bHXYPfYkODXkhcoaoyNR14Q+VeHG8mnpxm8Hrg3cULEstE7qR5eDDGZAl3ZkSihtRKlrHA
5md5inVUeDHsQBXADbcEwjTAvaDt5FYmlRE2H0oLQCaMAI/ueBbrDUwitlEXwSzfm5u8zG/tQdyL
u6gHjbQz5dIh+db34Me0h4/BDvQ/QmXHQuzBPD0qCvi09T5YGKYPvxeHQe/AYnqIeCNWXCP6s6O7
T1+oH2Oe66akx/nmT1jMuou/+CEDvtIFple36GYWs9rNkyI1vmwP2nrsEZ3C3XJJfTV3NLC4UjeR
dBZJgF6jvfXWDnTpbadUw1xJ53w5VLqo+BCrIHAWzplIiZeLuwuqhTLNq1bMt5oCM3o4WQpurza9
8Gkr60GoJlCHSAIj10UbxGaZ/hqUqMrHiKE4bJ+EGNWnE2ZP1OvJf7XmFUlBTh8X99EKV//IwiCu
wEpYLaVmzJeqTieKIMK5Pzm2Xt7V1ntQv1sToyXBKMPZWkJhDyvco4Bm2Jw7n3SWavbetTqxB5gc
zy0xzJvtUje5pp9EnJ3+DPnSjqwqlD4BtKE6POU1/FnwNFLmZ2+g82+3OwhALGS6mBSNX3nsnlZn
QZ6DNV0nLzjT2bsCTBlvtI/cB19BSphamnXs5AT+dCHwc24uXMSYkerUx891eGqf0WtuClb8+zmK
H9DyLtbxnLsNv2khwPCbuXVhd3bbNgZuJgucMp5SV/urlQWHWz4hRL+i8BMzxJyytqNX13s+ps43
l/bWIoZIMqqCioVuj0V9Y530eSKhXzzek9FunMYyHPNvG15ZiY09EE92h9rBkKDr5Tfb8/Os7MX1
ChUyPqNQ12aP/zJlV0XAVayMHNa1BwPSSDVbHUtOEK1EHxNEy9mGB9Sfo66ljpV1fwqC46HhygYG
dWLH7d7NmxOm7AkSCeDximJtQ0GEoAGlmbULkv1PY4Qgg8cLEBQj1UMipPhv2AZOobzIcJJ29Sd8
5krrPoZFInGQd/51OASvLyD/2RGN+UVkFXnXypSifUG+0SJ+SmLG+iazUuH0xuZR10QamU4w995Q
6R5MB8zQfycbrgE6HJE/TiHY3LlBW6I/8y2xS4InFATtjwqEpe8hl5tHnZMupl2tFeXLf24hS2L5
ZDhX8410ZysGQah6p3A/P3nbRrx6mVmlcQh/PttumeYpBWSFja7PsIESeR0sXADbRUsfJniRnao7
eY9oyg06YlDK/G0m2WDk2tMDzsGt4rqoFRtWm+Z0xaz6SmNaeQX3edX+aFYhXpu0XGm6KL/EIPWY
02zI5WM1GkOcbPmJKMTKK2pYHLNKA2+q+Cpy0eGTdGWmYWGdrjeqqS8VtBpIzEthC9BwNhUtTLDT
bA78gSe3IVzATdF9Yi+xtyG9vtzRgsRVCmrES1F6G6EN54RimP/yMyYBNOBRcQ00z1JxhfZYf1P2
m/gRfsZd2oWGw1g7xMQ/5keowH5FTEo/JhYovp7UPlzijo/dCFy4gU6gOW7n8WuFBrYZXreQhq6v
0929Ve/iDf3otyWVjI3yx+OTeIaYAX6AgIU4EUjInJ3XeMBpKEVhXBgtb+q4vd2IjaVmdKXjCJoA
BgajabgT4uVjLDzbEhInl+A8ZDvyfYlSYaYkgShEhLkEyyuDlA+lXZbZJ6y6vimTkvcmIBLTyJil
htd0zsUlW4lJ+Sp9B5vSofECroivrEuH0eP1EovNMvqoc4UYLk78ph3xBCLLY4ewUig+n4/f/2Uk
cbLr10ML4Y0yqag3dGeojh1ICPeNpkPEj84mftBd+fDB+cNw/6E2seXE0vx8YPHVLsxNeHtN2pLm
xPv7MElt/6ToHg/dIUPuaxhjTMSI+CKB7sNO1W0bcZ8euXIEVXaHhZbT1/aWKvYIZ7zV50G8gniv
XJfGsipNV7ezN2H+RnfeZESDxSQsr//bGvGkkiY5xJCv0ig5nb6JNhITEUpUpXSURAxqc1ir9zlu
8sskCL+lqRf4i2HMqcKqMtTFQoYfmNR+Ufe1Gok8FvwE05n4tNw8wZdVzKeYp8q8oX+2mMc1BrPH
QF8RTsRoA+BrvlQnH3xoUAHk0WAQ6CMOJ8pS4wFIoJs6lRFHx5qi89uY/gJ4CovB+MTrEi9RKUs7
CnxekqinBj7TfTU5Fzd6w1Z+uDghqUfN3xMKZ4lHv2NwyLny93g92qtdFt93S6M36ztwNIF4OZsT
iQmfZ4A5omw69jJdGD+bvVGdxtBnH/Ysl9J3GsAKiARqGh6+tH+1nh6gq5ZbVEJ2ElGPTEkXcPs8
/RauKK1Yq9v137crS9w3KM+n38Jvp9hqY/jfxzqEUUwHsEv+/Qsezjw5BiO/nVStnB7xWArhBrL4
gFkUERtIB3KdZmRaReySo2q+UOXv6MDyulzC/y0ztF1aFZUuZLf0+0HXt5L/IlCB+wdf9M4Sq2qA
5CZpi7M68+3w5QImOh7MW/tHe5enELXpMh4/u9PKjz8fH69fG18YeIZXGvYrKxKaFBHtSkHmuVh9
OZkSIk7s0QtRrp6XLerAEEnQ8sEwHopWAfE3xk4Y9C/OzM7P5icGJfQ/o+i6mlGMIXhLvSMbRWn4
OekH/FtZ6tRBeFOdCeVICABJwjKQVcH03v4x4TnAvCEDvroj/LJ3DLfqOqgs6nhy9MVfKApPbd7n
pquepVmYy5uGqgtX7DDKANV5uwMC3uYPojds1cCSj8vOd1QskZ70uel+dTzojNQdt3hqqexutxZn
rwPfn6D8uewhAICjYpCdexEKmgICFxFugZzzz3fK6ieCea0M5T51CC8jhzL63xUAd1oX/aBN9wh1
mInGdGo1Ptp15ZP4pLp0sQ9y7SsjpWKXZmqJ777cVgpqZKfZ7ptAUHb8DWwNjw33oX3YG610hX+X
sW/9Q9YM2HTnHqZyMG71RHHV7yYPxeYlfDIrF8HfTkNXCcdsyvhG7KjIVtTgzXobjcW+YLJiZkO5
0FA7r368MZOMrOgDvXg9ZQPg8fWGBu1RuoXAsdNArekUqXWk5qW7CX+VncComCbHOxaOMLq1w4wB
o2RiliSr6pf+tZhSCU9MQOOInfhrzD7WX1H2JDi69i3AVlZK0HwDkaZ7j4R6/5b65ahQ1+ldT72n
nBw4VQsbwKxdeZvLOtNbgjRy0uiy6gxKkF7PCdblm7SfNNoUBfyWLUQTlyr3uKyKMFc0f+QxFZ+r
mngE6NOs/jPuU0RpIuCQry+FIk1PUfw4cQYnaRXk5IPwtMHGzcKGnCi/mqZxaXqSiC/gm4A6f/Ml
D1v44RSFNnegQ6whALn2a7sf4Hv3F6UoHAWtW42MaF2O+fYQ+7LTuCmIXo1ICMCkxSVeYxkS36VA
MJvWH1dwxWdKi5kwf6iQe/6jjyi5SinIPwqrok722/EPn7/N1KnMlgInk5nNd7hNm6JtbrBcI3XZ
RCvGlaaR5j3WFJIxq766WwRNMm0qXR+0WfBGmArY+f5MmQNNuen1XsdX19pkMblrtDiBBfre+edj
OsKbSjbPNQa4oKo35Wm2mhn8kZ4oLok0pfcnUsVIr+eUSXIMF979seRHXZ9ObEcmmqe8ZioVBStV
hi19f+rHF4GEZ+YTTkU5ezpDP8rMWD11v82eEgOnn5O0rSLTDLcmze2didzTI81prQvJ8NVVsVZm
ixxQAmYGBON238DO9RbeW7u64MU7Rl6pD1zSAN29RjjLcUcHw83Vn22FD4sgU2EDW3UAsQDBVrFS
8Sr4BFbQqkBVWNxLCyomVGeIwV3qUThKiMblvkN1dPspv2xOHyBiNtNhGqmVcl2F1PNIxXvpM+hy
eXd3+ifnHmN7+4teoBh4z9nM8mWbXCuAJYgT1ARAuHe8/8+TyyyiuwlfXoeKC8sYADk4rOS8/vHH
fJKQF0ksY75KQlpPa9EvQsgIXjuZTj0DlA6nMuka3kEL9ucR5/hA07RhiXLXd9j2al6bINydtjMU
9K8nSDy5R7/cNnxhxxK9fsS0zkS7UM1kzl07OBJ0j3ADev8buZgNGcxr0TXw1jzBJ0GI+J8zyXzf
3bgnILJmF0PcwH1GO1hrFd5rUirZ8tocT2qGzNp/Fe5V7k8+7HyS49xta0vg/PbG8vg2gV2YhqOl
rcpjWqew9niEMWprEcllHdGolRDQfT0oLdyNXlU4h2VMnMy0YRmAFqNxjTRt+91zAlb/6t9rgA5/
v2Gv3qaejB7Fm+IWe05epJGo23/h4M4AiCTvQ1Fp/jUprVg+JrH4etN26/vu1lpB6OfIozDGDiE0
xzPZssybgBq3PLdTdmPDU5dROR/vCCa1nG4r2yMrxSNl0fnF5g2XCar5CuFigTEHu6BVhglKoSip
T5ct/A32LGBqaYuAEnJUb4U+z9cRoGSRP5/wIECgBJb7mrSkPfSFaBUsRTFjnsNBao89U/HcIx4+
Kf70+NB7blbGX3cU7/+mMdc4KXIQ0lhcZ0COJOC3sFki7TvNJqV7/OLP/YfpXEhkSB3D9A+u9dNK
H/MAEuwCN6VZGE20gb1Ik1ltCHY2QlFr0uf8ZdG6qlk9kwke7oLkY8fyEkuD7OwvGKTuF1IwtvTu
YxoDKvQI49IIbhhVsQz1rAkdc8SnpUXiNTLz7ohhvouF+DfxD421znPwRYAZBNJSRCJn9eOMJnwH
kRyaCM+QQJUumuu71kvGOqp5P5U0aqnMx9Fr1kHbUQzplG/BYtoUKhSXd9cyzjvyqL7W9hbnfg8t
HcnlKqIfsEKeDscwxtAel4EQsZB9vosDWcWVeC2TEDY2M4o0ZqFfu+8BcfJCY/vElYBMvFzO+dUw
v+RDDey5CrbwmFD3scfgLY43ujYqV2XSM37ahOC+8BQ80tyUEprogv9NSprvZJHK8VPZfwPnqiZs
Mm9/TzkV4ZTzWDjbg5k7jKOpDg5X+6rMkYMwTc4lhEturlgi8S64R2veEnLjvm4iso5zduk7nfcA
9HdDeB50BA6sGb1+hZzrL9hAlgj6VHNGeGZg/NNFt9Zip4OiUmpIfWiXpx2YB4c0JVDysZ9nm30U
h42CHECC7GZdctUK0WLkOIq36Rye7o2sRPwuM/HBElsEKofcC5mwMSJvchLcR6ZGHM3pwWq3rMSZ
EzyrJlpQybaI7RpYb8rP5U8F5JaNQ1qGWyiFAtTNtNEKxZ0Go6vDInrIIs4E6WgmmwP1d3q952Md
qJkuJW3UIjyuaFE2dV/JrADN2ObqjqQrZLOcnDC2hT4dsKAM2eDKfNl2rUAgKbfzEx4J9uEMmoSS
yOJT5Ap9Jit6hAAmnJ4GXGf/egHafdJaj13iTXoGFgs0Y7NXTmmbinVAtCMJ4Lxygf5zBjsCNehA
RP5mWsqJcR2PKr9tsqsc2imHxax4P17te0LWMzqbINr0FkF3a9fg0NNRuu8GEz75xlzJUsS/arKw
8QbgDynUhZaQn87OPEof2Is7fhbniaTvociljKVXmRx92ACOqAddoMUIcKhRr6UNCqoqBEhlyfeT
HG93IqM7XPTHBbIiI7Rz3AjDiXnQQsK5Ck8XjhRNBDI7TX11dao1w0s3jTc6CpKjh4Pyunz8idux
/G3uAijygWa7QYauIuaV05YwciMf9KZnlB7PP0noQWiIsDDFU93PxOD+DPDz7ExXQYEsgeVgROsz
90SQ2851gmsEftDPika+e9YgJxNFDDH41OC7XGE8OpiFuSvuNlwKklrzZqfm5y8GucJJLgdjjKi5
brsP/CtJjN2y3L3j26lUKfCIxVVrOcTHpycCnV9L8wVEaxdKu5r0mxVdNRYzb3SFg2Jw6qxW11Se
IH53G4AwNa2XNGvGKQEJYBYayhrukI66qUtqkRfc6XhYfkfjKN78r7jKZRFuyzgZ1D87PNMYi1c1
B4llNnrow1zSBtjL/+2eL1lJ6WTrDTz1Hun80K1UzyIKnb0q5ox9mEfrS6OtoAKu9qaBXJCvqACg
8rKUYOrWZOzMU6xDvJllkAdXL38PU337hamM5pIaAwZbbghKEgbw2K3igEuFk13CY4PusigSeb9Z
2H7tDzkUs5VcYwHijt/4KBiNtJ2QvxYwKi7vlfZ450kjNN4DZQqJaLrw5J8Wn5BQPgik0mSm2SNE
lTuFeVOVR/jeWx5I9bTQLMBVSyX2bJYHdywW37FqEOplKnQI4lxktiB8Y8yNt2IrOrho2QNkaX4j
fgfaYpVcH2ddwLMa3NQoBJTjXCZDCRGOU/XKLf4O6FvZSTQcI+YN34W4hQdl8D2VkioEdyrpS4o4
CNhmzqSwjAvGSb0DLeEfi12BW8PcZMviPibXWCcJA9d5xaUNGlKoX1QG49rsF71OsfDd0hC1SjTA
QGxv+xEEeVCbh/y3m5ATkz9bTX4fOq4afEFMwOz4V447GcIHr1ctgRiLobQoNSeK5+3HU65DeoQ7
f5TTDJQPf+TsGa2mZUsOyhaq/FKMNiapmMw6ZhqNXzTHkTnBbUZMrXdXmpmltJxKKGpGW/y1SAnn
Sy6KFr5wHzEQqv1QEvvSqpIbF1F37xocpzSJatcaTUDdPu63gEdeG5J4eg2uAiC3aG5OUQ8dyl4J
Yn2JKcFn1I5K2lvmPPn6XLrq/F+2UbcG1jg4ttxSVFxGdM/U8f8qMUQb0tgaKFBlu1HR+VqqcLDe
sk0/eW747Xmx1CxQPpLSF9nj9L9BP6Em9YZxxGuRqDrcQP+7f09tFVHJw0Mb8VTePdQ8WqPOWjxg
bETI7RouiqGcvP4AH6z/EcKwwI/YsALtF8whvkpwvvSJWIzZQyU0b2DS6iZyu9ZHruNIshzncw+5
U9kdb4OkKkGHH/Y/wy3TrkhHIqCFGXkjOQ+NeGK8ygRyKuxHVg5SLu/LIrsFf+9VMDOULsWIXOZJ
W8v7miuVDuXSy9jd+t4HvjX2SeJe/1z1+9XO6g+alywr+vtoUG7AFoiAvyz2HduXXp97GQ8QdLKH
0YWIW+0n1KfEWUughSe3jbVFzS/CNVMNGtFPigBqMHVZTD9YX5d4Ww25IfgBIHxSWVdkaChhZza/
WfB+k70CCwVGniu1AhUzaTAk1vKbxEEwFQwqTjHXSYXZK7/HMZGwnmPHlKK7Zd2sOMEr8X9VDCNE
2aD7epmwpyFWGlrQDKn3HUfkq6KOKR7cLrIymzrqdKfhRqQd2R2KYKfi8aAvpVAInY8RKafQGo1m
uIPHT/NgHKz+WNCoq1SaDVyyHBmwsxHoX+iu0ASvbqwJD40FuBMUCgyIcc+wYDtbDYHeuIVQPRqE
aSmNHXTo42QdrgVAIFQOK9YmVqJI2LxX+RgZMsaWxgaSKrzWyXs7/oZ31aFRxKxzJZdh1HBVHDta
/IZMP7OBZR5yXaLNV8O/HrMSaJt8yCqHk01Zpm3/bxyvntDtloTs4ozVlnS4MhDIevy8wksi2Phg
WpcViJlytCPhzweFW4L1jkbJmdAmULlrNqNR9LgrbCR1pQtZzisRe6iDRHfa7+74s0bGhdtQ3gFc
8fPgBii5lVCJkePhW9gxPaeqzm4l4ZBmFnLH7z+CjF0yfUzxQzuKr9Kz9R/OF4fAJPoH9dn2WyG3
V/wRhAWlxrS2RTAtzz7l+rMqDxM+z0Hm8h2K6wvFa8Z3n0XFWuUqguR52eL0ZjheGAVGVwtvqcGU
M9SaDc9m+44CoupXKmImws9Lp9VieAWlw//zeUPUdRTQQx/6nOYMhqvoYbOvFO1EWCjbYpe37+o1
kpIBzO334tK95RlkBi1LITujm3pp6N+3k82Awbzun0gek+Wrb0HI3gQGIysw6xXMa9HppXpRZjah
1w7vQbHqjmcDyHUq4AyCIM5AUhpT1i1v467RkbJqwf89XqpM9P6yeWrXohnIna1oPPuKg9OPemtx
Z2cJZ/Vge7DBBHdCVWuJJbzfEYcdZQZKAjnFCs5ThiBDCXUZz8FXLCyg253cJ3gyL6u2ipYXMU4i
9HnT2LEUHTRRRt0dSD/wuL3mkgRhpBnWcPsYWFgXSba10AgZkzaIvk6bbdYzgzY3sqcJ2XgylzOT
o/6CAOUqP62iTNxD+sRXrH0gpabQeVl3Sv33JIMcmDODoUFJ6tue1oDfgWni6ivc9nt3crJV1TQe
eJ7jemqCjC4chGK+Vc9J8t41iUUJquU36HecquOtku16UvSMy0gNRMjbJWW1Y3HxiVCFj5tuAXel
4g3WYdfVnqB+2Z1090GxXrITXe4AnK/Xcy1yxKRGRVS3cTqsBHQucM9d7UZsuvLes+KgpIYOiKuJ
F7OSGpgF+jK97M5vFoWDf0oZ7gJeJD1KlleWYuDosh12/HiI2Jwi3gjk0toIkF2bcIa3zCyUIFsp
PD7IPRgbuCf8nauo/WZ+AFnHKX33yIZOlmpSlKgYgZ8BdazLKpkkE3Zv7Oni2q+I4cfQdvRq0SJK
/LbRTY5HBbzqSfMcvGPKdTVdKntJWuXg5jw1h3wVHi641z2MeJeBIebVF0neFLxiAkjBmyHx8wwo
RJzQwmNyN2OGPMMymrXilpSnEh83qoa1Lm/O1NkL24oaXOmfLjo48dGJ9Y2ijOEhYoQZhh7XjWA3
iPFGkixJCn9WpZriGLgEfjrDyxJg8DaOWDA5pejJm0AeVApmq+eOiIPZJffWNqolI3RzDfAlQQRe
inDSPCTc/5A1TmkU7xUSJi7aHCbfNizdC+XxtflhETv8uEHX3rvML9V0gdkdTsMy1pmEesKVOPD3
SDvSZQFO+94+TdUnEp5rymlM+cxanLafcETgSADEeKpO2ESekdXepRIDwOju0mH/AJaE6ycMGaKw
e5t5rkrfj6fAnb+1huE7jqxgJbLK9W6Qec4wcXZR38oX9c6QFHNMsYRImLJ1BqWdwecjjAcVtxMX
lwl7/mYaN7pgsdSBAVMCFZg3NAwydMF3U9/Hpbc1zVNuX0x34d9l0zrlXefV8++lYULWKcEdAXgx
JyLhXEHBIdzyAiXyy2phkF7Jr5TJdMSp0kwSJfEEMDRdS1YWIorK4qjWjnCUO5S4CwbzrUzFbV/2
l/4cHFTn3B2awp0QXkS3SiDfVhkDsq7gUg9MeNOvZ2kuns7BhEy9OJXW0mR1fjOv0kM7METEySd9
3vn1u/1e9twnbz6Q1UC+Za2jaiWJ9GnPHyY6jaGQQKg5rAURJrIH5iOuH9Ld9NJlT/gW4wdleOs6
xAwZAKz6n5uu3fq50Rne/c/RB4hWsSHxC8WJP2V20UHkc3v/WB42SU6X3+MfA5mrgmIlL6m7MTXS
TyX4YipPd6kE1Tk/BPgVIxeeroTO5Ej61j8zoHRXWHm0WxPuXgSh4aPXh23yG91OmgGXMh94r17L
U+0HgZulsxVqyZSs/RLYVyobmPF6br1Ts4tghf7JvbS3UBO+CW2sL3epH3DN9ODqEBIB9OeGC8lU
5D2CHm3V3uSXI8EwM2N7fxrLJAGO2MXYV23GGQSDrkLith/c2qrMgJdQWHTTclDrC3ncq5eldzAm
O9DW8bnYyEEzzPAyttThclfkli9UEpnR7xluPCXAQSpq8A18tU9cJqxwrkIEIVNFEVGS2OvTbQzq
EnX3v9MuhgON7TZKLIix+3CWvpdRHWugnCDzvCX613n+5/SHMZJwwTvHNjtphqG19bjaiSnquaO/
F8JlPTdLcxNoGrcU+KjCjczWLsUhSOEe6Rw2Husp3hTkqtxnHqcfpUMabH0xB4ZKnVlPj1nfeiCr
au1KMiLaAglqQAO/6ByH58HuCLGW6AG5N5lneDgRjMckkAnAd+w783P5Ix45TC87iAkkL+CUywtv
s2PpRS2Hn6ahbu2rWQBDLPOrrkd4eOAz4x3uAGWWJ6FDYpURbD4F6BkLctxLLvlyms9ByxZoj/PT
UT6uPu+oTAct9hT4xurW8BXqu2U+8gHHW7iKSb3ayFMP4EdmPv/fqEZM+sgZUpR/d+GWHKxzJDQY
kxRXGdAhGh3Dc4VM8QPxPUMnnUjIFQ5L6BltphFVP+dBBxN1dRuKohhLU3kadQwBYaSdKyFIP4lm
7GZwg/xQx64zTIhXZ8jttRqL+xZi74HrMKzS7OtbPKKXbITV6b0/gb/v4CJhZDh8PNaPyCZ0fb7l
QNW8h54GSdyu/rxQrzx4Y2iF40m9TNqBxOSu7uEKjtMyG7ItQKPkifPWKEWfPDlSsDQkX5XUQ3j6
Mn/zptOcZsYtsF808TTNCxkLVXPC2OGhWKGbdahs1cSvqq332IJVMVZ4G4XKV0Lk7OcOMa7eDVU4
QCDcCLd6X9qrgtxXNxGHjva267jK5flQR+76MMabxFxlzolFT3ClQHs6mwsV+uV6LsEyEcQJ8kI+
17fVqROHRc0CMJwa36LUhYO1caREE90TNRNAVXmw/TFWUPeSjhTEWpfC9DrWl4wgMYXNDuhJzgvn
4egAn3TQ517h5JcDfCVVyFytk3kw0yl2GuQk26B+GNYLYGD575Zz+Gd0OO/6AJ7LTOEfVzDhbUj0
Y8np6XtW2MFUt1XCNEOvGIGXldGArlR7zkwOjHqQZ+A6VGoNBBEaLDfCQToF5Dcj1Zug+G6s8A/i
sJcy80sxqsdbnqrffo15eXs1hp+1FDuFj+64jQ4BR3Ru4/npQrX227IIOzNgKi3B2X5VaM4y996V
HNzcZQPi9cxBAJi/+rerOe5essuA0ZEhlTuF06LTcJjMNjQZ1+zb484nVf62+QJ9wKY1jRPknPu+
DsuN33PAyds2FMryavxG4b6ZTQGwNcD9qOOiKz7TjivXgIH3Is++ZIGDGHoB7qhDGObfKPOi+G/8
CVZPwct0PLjAkpZNhQa1YfzLUI78taDMXkyDiizBE+AaJwW8eCpTuZoYRLE0WqdUB1n0zWHR708g
WUkfa36cCJ0NAAuk758cMvI46zNYoYVWo6EcQTGMh+DAUc3Bg9w/iVnLrNwTcVlayl9VxjyZBNYg
paVsjWlnK1yf/oZeoiJXcp+aCL8tnH573JECcsL4BtYk8QFk7KaJCepjdNAf6s1PKN8TCduahVZu
jrbwKVPVHZb7ov8WveFM+SOPg13LM6osGDXach6+hKdaE097v8QpeGtwoqwt4ymU/F80xk/4D0zw
9pJs8VXlSt9WxAOt7H37gGqMfrdnLNsXrZVWdYWFcGFpvO2n7bmP5smd7pHKbc9XwwzZLTfuN7S/
NJqhzMr1gxfYAHwREvdRcRzhjOmi8wWW7+NL87pXMOqW6JvDnSFm0O+LvX5fc838KHwdBQUglxOI
PumZaDfa7tBvC7C6bwlHvwb9LUqd1aVnnlussxfSFAuIIoNks9sFs9cU4P2NuCZ7SX0aIokzCMpz
fqxwtDPundSE1cST7DQ2Ir3bc5IzG21Nv9LBy7k2LcDCdOExabQUNnKAT1uWpER9PrS4tYYT9TN5
ksSB/2pjkxUtdPrRkkMFKe1H4/bv/Txz1xKdWiBlj+at82AhjM/qjnBjXM4cegcqY8PBSaljFvT6
UDN+Gqb+XQgwFHoSAbej3SFwx3uB17UbB63GchQQhXB0eEjFOg9/Z4XJhyAa/Gu74vEN93MFQdd6
nAaM16HydAgAdd2Fnmjx/UJ5NO2m7ll2sDxUzDYeujhJyQ2EoadmtFkUKXouPH1Hq2eq1mZPGyX0
m9w0bxIqp6rPGMD8YabRgJxJKSfyj9ltVoGkq1el/UT9FP02sq+KAbwG8fADy1MrOX7gD2nj5tdP
l9/4Oz3gcgmrxCkFKWcrL+Nmj0JithIfVtmgfnM9nNT8ODBAMbo6L7emctiQo4PEIjJcKMTz2Rnt
oLXFz8nZEM5ReYejImsLOPxpoiwbkn5u5wIjvCxIyKAz4Gnux5xu1tVbPqRWuIVIrpLY7OzQxlAv
8Ie1kKIPgjhDjfMKlmDiHxmah4hJtP8+/zDUoeGzDdCzy5CxKmLKc+sCnaZt8FF8jTyZcPvkaq7H
YGdYoKAnOvsRXMoD9NSpna4vz+9mluVAtFBOeuuWdGkpsvQgZ3S5N+nbH4KvDFklEDP39Hsq2mjN
LqjThh9yF47/xBMboI9tyBpQ2Vx3B5MBeufD5KUXZ4uvp5NZkAFko1i9Q6XS2PI8/Oj3fUS3GQWM
4ldvWD2wqmVaPIkmJ8HTExL7tGZxm9VIR+0UpStz6Qitb4Xonq03Proz3lwtZo237uld3XFoIG9W
NDGpi0Q1H6hEsDhfSNsBpUrfH39FBRgH84FT4E6dZdam8XnndYoTfX+1xJhV2Xw4aUSoO5ezFU1C
I21mLxHXL5dHr4nQ+Tqyi324UG31CK1k+ZxRWprpBlXJdIg3y3LEeBdBUE9QlhjVzL37qbwr+iJU
c8KBCr5v1vjvHXTfauPMMT2sIIWyAfnJvH3zR7f0Ha2yZexh1Q1lKvY3oE7t7nwmHbAmOg2SEK0k
+p6oE55PHiXJtXKllr8QHU6ulWCPcFBwCUcZ7dJ8DTK8dDN6LX/h/4ZOe44ukjfOL8WK4wgjc9ZG
FsCqjzP6iinEx1FsQBN4r7VV0rwXRQWL5CGOeHQIDFr1DOv+Yrs6KewXh7wrGoW8FchwdfjeFKHT
z/lxuWpxhEcJqCTFl/8sWEbcUna6Co6hUcevDYiDZs9VndBxlWMMjFVyfB7R9d9OybHZJlb8qRpu
a9Uhaynuwrl4V6OZBg4D7/riV9/T50wPpM6T/A2JAOvutR0ftB+hQDwEitz5RrdNRA4qY3vkjr7d
0cwbQRWuR9FPEf4K5yLg+Ml7MaI3tKQfV6oDJfDcEz8ekaNC7rTJaLhvAr6k4cZGn6jhZBinr3K5
Y5yLNKVVx1UTCV9NtBav8/6+tFILFtjFfRGUjHvmZg9Qd9hK3Sl+4wGQPZswhSYHIcGWcHYVY5x8
cFSyAHv0PV0g0F+meeF71a2jZoxOAORixtet5UZ9+E3Yhf6Qc+v8I6x0oXlT1NrIhszdGs8KEr8t
mtlTmPUFVq7OM866/saDqNLpr+Y2h6Okuabj4Q4q5uP3I0/QVcm/YNQ0yzgBLIQ+jhh+j52U3jVJ
z6zgcuJngEMLAM6/SQgeNY5HAjS+h+XqldO/NJHap6V3jtTvfaX4EjS8ymZ8As6fFwQfxMo/05yy
W6MB5Mn7ORQh1gGGu9hGW04dp5VUb04pXAGmVAEROWb56B//k3VgHR6z3MYMq/IP+oQC3/wQx7Qf
vCyA043MbPd+rGONh84QXj/SKigm6dNuoviMmExYSi1gSnR1Fabaj6V7q/ptFIcBBHAlSVRf8vtR
Xf8/FYBp3B/SXS+SWRloNzYYmFBjnrdkZ4+WQCOk2uri4iSFzbAZHt1Kxexq0zWoKuz2m2hisVyo
2CoaY0aHDvyJEp55GxCak/00Aovi1jZ4HKszPwbD9LFXpj2wtQk5LTvi81Xn10uD7qnl607FW0Fv
2UVByp63uyaCLoDHT3UsoAfUVNcz26a/36e+/lF+eSTSFxrzfgaQRGlLdh5jN3bn5mOVccBQCZHF
mq6Fw7OBY88lo4R4y7W97ipFL6HF60hmZzYKBNGxYdfjyqm1h6Co8kGQq2hcqTEEpYrZB8g8YXku
2UKmq6YChMZh6Z5Y14PPl24hCDVVt5J+yUBakBoBuT+/heTyLx02JG1y4N7v0ACglFljtwAKroHz
QmrrPrG58CoHNuqRUbw1ktIp0iD4W18HLk9XFOGJov5q+rxgmLXkTUkbTb97otcQWdlYuPS8ArCJ
JmsztXvHSaABtJVB1wKFJtri5OWU4i2PjH5a0cyeUt+ShbF2b1Vzp/b6+/EL60m7iCFelCQZxjIb
VdSjh1+CYUI4WYNZ7527CARAT4TuXcn0GJSOOGtB8wxgsZJONlWPfB29f7wfLJuM2CE1Wahat6Qg
4bKYz4ShZo+8umlL5kQf8SMC8vMq7kmh3sLiYF357P2b5OHHz0HMRC0AlWPJ/HUdoCcjA0rVCtwq
lOOxOYsKcH8eZrUUl0f05FZ6W/wi0PaT7xqDDDjq0wP9In/c3HW0N55DEhIsejVJ/p2FMwrONhAg
RnaKAxKCqGpxrwtfNP+MgrnYbljEZUP3AaRMBOQVqH7WtGAnPU9VuuPZCUNxZs2BS0qHbOFX/Fl8
o3roLCcuqXKb/WbG6qbgjKRZ5tGruZnKV8D5a+zqKgalJ1IuGCEEkie2K2LQy4tU0GC9WzMNeF11
E44OPuc2T+rqPaXY9+3coNVHtMBKRekCoQ6fEH8UBYC6L7O6AEQFvthnD0I4xmfgM58HupsJXA4Y
ln1cMgNZacUhB1UAJuSy42oO2AwKWm+mPb63Dg6kCgK9+zPb0YX5nlxtuTbmHVOtcyQZRIYMME2d
63PF1EYFHg2McHUZmCSTzQbgVHsFKtBVyG1A9Nvt5ZlG1G4wk+oNyeX3U8YAyMEnztu3Izxzq3dh
/hJZyMM/6t6F/0sN7mIzqk5+CVw2FVF04LueLy87JlG1r5w/IgsKye2oSxzmsSlfqhOugF5XErrx
AtfzgwoEP49+mN2Pn5lLT1Bc30YGxWbMPYFjW6K7P5ifbm+pC3rH/azIuRByxtQOl9MOnzxQkJis
8bVCfNr3cfra0WXqXvtEF6we8U1AFtas/V9GboEw0XPjxdaGhZua+XNDoIZqyI2gp9YrUxtLAFjn
9CxPUP/RImOjxtAqBT/80qh4JMtfPj5BVo5Hqq97/0u4t8I70mLE3aU8FdBNsXwjwdv2QuXb+6zx
NXNoJ/jdrOcw8NCNIUfkNRjLueWIIO8GiETZuANVSJeTFCxqn+Nh96wHVvzbiY9w/164eNK3uAPh
A7wPWdzoeWoQ4rjFT7Ncbos4VSt3qy21fMVc8hod1N2BXUrKNh0GIFrEi38nFksPy5BxWZ1sVnpN
9hqiW4+BsM2GlGb9d7uXceLk9lIP9cF3qIB6beQSToMfD9TYpK5z2e3+3XkbmGUJq8OoPnsX4008
jBTAoNYStnr1ZmmkPcLqUrwZpOQ4zAAUQWz8hBTaKHiBpQHM1JhLp5C7ZGVA7OB9LhH3YQjQ2+6P
LiqwugJlg2hBVR6qu6NfLgX8dyb0c/V5ezso3ASAh8xIxh/hcCn7mRnAEi65OZJrveqyMPxYDBtE
p1C1YBN3gPpFL4dDm5hS2LI/K1Xw3kGRcZkggexHYcoiu4CPxSvEFq+jIiXIwxtjq+x48Pi0jXv/
ecrEKdDLko1BWZdA14+XyURed/SEy0Fl4945gj03W15mPaQOojV4M3vQvYtaQJZr0pceyMPF2bPa
5YS4aI0QSEllM11sCI4KxJUiZ8Qj33Rfqd3OU/V9doQEdqNJPv/n2LF0mvr4b+WIs1rP9/N81NqU
A8Hj7/u/ljmnt7kyLDExwOhsEDp7RwI6ihlOX2gbdHROAE+9x0hQXtAxkIHJDh8JlisreYB0B8yt
vsh0zaDZf4Mk71vdfNV7KzvAlHF8e8gTzS/rM4KwauX5+oZBym5IoQki/zl9B04PG8k/dJa6/ATj
G04N9I5kYLwjaw5hiPGep5ej4EFVP3qDxPek3wwDe6BRDVbzjW1dixbNTyw7xE4/FUsPSVvyCUZG
AuAv6VeHzkNH1YGWzl6EhbHLdsMH8fzc/+G0DIJEv20teHc5vgEEhSQToNYeXd/6+HUp7EXpGvnA
bkhf8QRs4reWKbHKvh/k+t/vczmPZMQJaEFTvfjQymBPt74GbAsa7eTlxYfgZNloTNEouJasjAxN
x1QU0rwPdyv4MoW2dQM/5cP3USUiWd8SjTRJNGbFuYbiG5vAeUTWu7NB61OmsHRGm350tUQpqOYe
d12c6zSjd/IhX87TSyLeK8xLb0rGBpW6L/yulfjxr04SZf+ytojKKfr4EMcXpct4HlKO0O6wEyiF
HMId80YljHxq11HMc8ygre27SpYEpUtGFfkCTXAJWlqmeSNWzKxYS3SEoBCAOrazI813tmbsE6Wu
siFRKaqnkciA8DkDvU+85sohmH2KVpN1vTh4exJOrDLRxE/yXulDhuM6RsEw/knUlKXeUHyFii+M
vC8VMFdlJQsvNzkFagbeuBOiqke7k6fjangJ/DdETfxwsuM+Iz6dDaISE6A54+gSW2i/oBIf08Z2
U+zsOuE0XFG08N9ROgOdHkud2dQEojHzIdZpfcB8Au8Y7a6bQp0+FpZ/Ci8GhRk5J5+mo6ue64kS
ZLog0X8KWTTTDrEZXpxpwLEt6XaWkXUmsO2M6QXY7AnAx8oafBj6DntAwHRf7UPLBb+7NGlQOjEM
DiJMwb7Kqm6jd7mDPE4/A2W7Fj19ukiEyQfy6iwirIR7XsO61UBQHDOi8nbSqzsjkWf/6+6SF7uE
Q9lM4TnD5fN6rYpNG51fcB/Q0ZPaHXiJdLw4mw4wyEH63mtB//18ciMcmpRZl2unX5hywMIGL3k6
YBP0OfHcn8LbKIa7FJSkPjEKpL3Ihcv5RALpiw3jhSSExroDJZhngF1Q0F2STyCIeo+OfsbUzhn3
vxKIEY4mqHFar6achmpnIZQFWbJzGnhhtgnOAzPI3B8kgvDeCi8bJIMowxCJ0HelycLw++PxZjgp
EbrQ9jNGL4be2uOeoVZPNk4/UFxOFbIZjthIUBy7wwo9nt8T4aFy0fimGJppSuQrYK4WugFGSko6
mVPxVWZ+pf184K+DdbTp/IvHLZfgiHiZ2npBbox6jtc9hO4hImBTf23ahx85RMniqvVnrYEtVwY/
1QkJ5BzE+F2i4TYg4rbNKUor/XRKw7VUk9vWvMEO69fguFlPh0lNECWbOfT5MG3ejJmtvG1lCV71
knj/W+4kvVGl7gVZca6o7lT4zYvmw4NrjATtFGnP47c4Az8UeAAUfEMRi8X9/yqgtD6nkXxyhdQD
g61y1tHgtKCRcfj7zyuaj/aIISetgOynAOl/me7PsmkmXby1lWe/k69Xpp21pEvjHvv7LYpVhB9t
DT5lPJMK/aN9OgnANZhnh/itycH8XRNoyVca7ay33QJkfjpjGJ/U7ltc8ouXYp5ehxfbugWxfqtO
TyWPFHj3pz3fiYDYOjBw7w1q2k/4XvWkOtVGvLhMifHivfKFDWw3hUhN3rf1dZo60Pge0aiSRyQx
ASCFVXXatLG+VDmosFKGqilY4Q2t2dT1AOVPH/yHgQm6B/GKLMPRG2CZqiyvU///BffntgRN5zR6
9yVsmdgMWu6Ebv0Jw1qXbEHp0JVbQevTfPGKv+P5XNZgLd8Pm9daJt/2OjzLncMuBoPzRyolr9pB
ekRhcoRtIeDrd+ma/wr16TUn9+2gwO7hSP3qwjSnMCo/Ip+GcpSxSB4MZslxjjHUfMSHdcExPEfk
eF6OJ6cWg200Gv+tu7MDleCf8PZY5uaaJ02zEzLrUhKsJjb+e6U/THA+5iF5h8xxFanWylFwTEqP
Hk0XyYEY8jVAaO2nx0XSaF+p6YqLvXbSny2LcAG0BxUk7b0I+7derOphtiKlmiT0IfMFjiQdGSno
xnbo7GPOWIXMwY0PcB+EdGJh0UaJ5AYM39lZ3IsrpNgd8BJxkTdiCXmYspGwrnSOp4YdFPsuaWDQ
p7jdrOSDLFCOyAR3sdc61IDL8Ui3vg0PQ8UjdUOvhYGp/pnMGhkwhwIJtkxpCk9LuNdKmAYvcUZb
fclKvNHkAGgtZ9GyB8Hy/2gn4X7mqle86LOqRcfm8jXYdF50dOcXFz/VyqjNEJkfMz1MIvvGkkez
TD2MrSnoCoqLRZK3CVCwHRXuhmwj46/DS9T7rBVtFXoXbVml0DaMsli+BNt+VNDJqBEyehFJXtR5
9J8lL0WO1OM6BvZo5pTl4jllYXLfQg5wLuMYTk6hSsoo2LdWOT/HLer3xSu1MWhab7xdM4IsO2Jt
7jGVDvzdcGKrWs15FA4clTgpzjMGIUjKdTkLRtbvkDBUYRo7RRWl05ALkQ1t0wX33uQukuB2p8Zg
f7BcU+wI+KZamNbxm3pWkP2kzh5QJ1DqLG8XT3yNslkJSAmj9jngVT0z3BTYPlkxyVGqUpIQpw3g
839/PIL/8fJTNNx8HVmZ8f3ogJcsOeIPACU/Ywm3joGs910ONFTQCXnYbJBPQDVUOkdtv3uins0/
dssgf2ul7yMCsAVHyaXxNUgD4FpsF/FbW+JlOoBkzlqDNk/IT9KLGEZPqzxQvSZqCP36BDuI4GTB
JxRF2sEQh7rb3vmqKW/yn6EA/CCld/Qnnv/gesHHzRDi4tif8blUJrdvyE7XaE8TE1iWti2dtHRc
Nb+QMuyjyecSemn/PAKSBlM3NhGWkY7/mmP8/Gj2SdBIc1yLzUn5o72VJrwlGHHCNpLpa0Kyh3Vm
1oUvgk/GF6H7yPK3Ah6uFYmW0evKH08Q/+yFm558J5w5dx/xqH7/NvUWF3u+xl7y2VfNx8s1r/Gu
RZBMd/m8bCevU8t2ZISlVYSmViLue5n09hjwtWUWc7D5PqLZDyTVzap31EcPp+9V5LG8nezh8Oiy
cIEcqh/q1s034OVXNDCvHdcoeaRv7CohYZSi3jTWYbE4F4M9h5jYubgLyABIrhnc1gx3If6vHdWF
4xHC726uipc/biUhc/+45SKElb2oT9cEIrqg7WZKq3j+4OK61l2rTMwe6PdXif3V8qYVZ31QG6+W
RTqn4AzqXJtHNWnl1LxloWnRldmYnHN5JdDVkgBPpblD9j3f2inR6WUN3kEevATzfVkO5TcNyAJk
+lHoK4tLeLYhQohj6C2VpnYbLguk+ytXvUX1xhBlAvqGYIX1d+Z1uH/TFZZop21hg/tMqeWcS7xs
Lb35g5d6hkOEu1SSUj3YsDov9/XrzWSW3sTfWLd1Xh6Nz2jyuTPGmXBZ0y9p3Q2vrP+d8Aui2ZqY
75jdQYahd+oRx1QrnUuHY0IOcKA9YILYgOFrCnCsW5+ypKPeyu8xGuEfsoF5MCG5+Sa3IQUugd5P
C+B6ck0kiZex+EAmTrMZ9PngAUlcx20TNcGN/7uUajAlkR6B3uVFmqDVo9V8skELc1zuFMH5IrvB
yhaakUQ/y68x+O2nEN3ZXMyY4Jd2+8qvoFhLsJg+HUbJoaH7u7tHEcqsFMHV4fRSwhRyenhy0rs4
ljrrK3zAv/zbevWFUvvj+6to7WQEnSpIdo6OiF9d+yG3NBbwu5m+MI0GlSlvmH0BVKKWQ7xExVM3
V2dyFd+VMYG7qQiseDegvFc+X9ZsO9NopONZefgR8YPSxKJSGW3BqlQajHvHxyFl/b5a4L34SkcQ
FKBLhaoy4rjSATpfAlIaWnEafoAZ0nzMX7wJG4hfAQdGQqIyi5LCMrDJQW9rzex3PK9Ug2a4/L/Q
fqnWYhrARsnfrWwpHMTD24wLBwUKHe2/w5q1gVTRo7+XvVVaYFarSdbDAGT+IcA1zlB8NvRnwUgx
VZ0R12tbIPtf/HXYJznrySWRzlYXmiheflX5zu2KNxrKX8MpsMIHjHXc5AHlKoaDND2cY1dppoBL
xwdsplVJjXwkYHZDcKEAiKt/9S3+BeAEs0PNBoA050eDXzHXsF74HeRw0IlAWqWPu63zky7Wd3Pa
y7HJvDoP7eU36I8bs0YdVmJ65D2DrcSxke5ST/BznNaPOcrjqt+A7gKyh6ZPlCM/divzse056MST
2+NK10kKtxWqw9NNycgZT0MgF7cv57t2PDJNh8TJP+XWt7yyomxDDM+Y0jDHpkVTSksXWE/DwbZ6
4WIviFyUq3igt/W5dvOfWvhfI8Yjj6iT2zUdszzXzrINbJbKrJthAeXzPPoTgb1c4ha/0mtNHTzR
h3w14J4LJI5KTZv00OeLtwu9tIEYsaUwSLzRkvqt6G/zOAdL1aQeslyv5s6cr8bN9qf4NZwg9OSj
OP3xrVL++D+5KYLLk85fdGOsVWxZawYa6mJT2VmIIYCctqBkx7gj7iR+V+e4hlPFFAaXcqfRcBsS
au7w44VCqQW4snhZ1sZjcN7jDVBraJBbym8Vl8qzHtXg4FlJ5jLswZgMY2gGlphfUkscCkp2DwHn
/l/kqxa21ueQFZeB1QXaGLOPIimf+8N8F+igqcqnUt758z/upGjdANhcko9T54trxxGCT8TdEISH
nOEnn4MlURXR0NP5XB3U9VMis+sRFDkgDItEowmB10zYomFL+JQycuxZQoe0ISHufgKA80bzGm/V
Ajbc6DNuAO0vjnbbt7OSmmNX5TSzNsnocLCIM1CWA9gmIuy2hNrFeh8LEiG5HKBd49GcbNW5+Vih
PhyCJdzpGolBiwwZLBXe0zoXo2EUGx5Nlt4AaIXLlO0fK7EAgX83I4hbuJOvcd7ea8Z8nmUVxN73
iYtoylg3MkKBXeKXl2sOOOKfxDRsVS58j03CfufluXc4g0GSdbJp14Z56mmACEnS6iUjgYLUG2qA
TgUvvgl8OW9YTtavQb7lVfPkoKkCvLbKPaARGfidMxhRwfJ+XIxrpUzquoHOZzFYXRGlDlbp3ERO
/sYJFoBKMAYhxpmwu0bmdE49o37XqTI8EO+/VFS8/7NVT3p4KnfSvrk29Oz2QX8e8EXK4HDA0gUi
qw40EKgCzzcDZ1OII0ifgx2+LIk4hRaMCOFmjUxR2S7AmANPhsARZiIkNPK9C+xTb4QTpo/MIJAf
acTbT5yazT3nlb2evDotjmJKoQLzgivQ6/WCo2CU8RdIcDgNpymtc92itrHXbLxHIgVus9ditx/R
24wD8fXhb3oL3LD1t9TtRbhxblGW2MTIZ/kx0v5OWveVcHS5A1Vho8OvjxVr3W/PGKi1Wx1fT51X
k5KTINO83j4YPiPw+5w2miw/itiwEvodQTqhaW+HsQD4S1GrrNQhzeIzWun3yJO5qjG8RupcWbJB
hhsuuCRzd8WB2y1hBYNLKnJuupiy2QEzheue3bQ0cW1D4IQTXRYxSBbzpkbW4hk0j9+DgaPLfcfW
la2qkxSjgTbityMvBugIXxeAzxtpqA3jHODi8LffrjTav4IWPhivIMs7L6aAsycEzQbgNhSiTQ1B
tgwEfkLJWiPmO5Ou4aZSA5aotwVArl6uKhPUEBl1WnyKzdxD3aYml8zIcjTAPlxVnCtBRY0dp3UV
pWpyJtMFSqApjJhaO9bW50beBS186tKwOQl8eYGES5kqAP60CXZCIhFbImVdPXkUgZ1nbGoskKrk
FSVImZ8eJEcxW/4my057Pp09307NP2nrEw2hGsKlpt6FUQBqt3iwUOxnI/G/VkAh6lYiAr+1s8VY
ebz9yVyFNsa+ldBlAL1o5BbX6zR8RPdQwhrNw39Ks2bw4AWBwzhzl4arJKFFaHPB4tse9WVtuK66
JlnvFT37GO3udqI4GX1whdq4xpl2l8dNH8POW4Q85qpCBs6nDM2kXrWsi0Ext8BxmFGc9lnWT/7/
xWfMfVPnsRlbBdRyTVFRDwz4CHde9vBBrZ11zVJEWMGt4rKz+D5D92W+MwJPacgQOE1ciU1nb9OS
Ct83i7/cJHL/NmkVz6+UKvPDQMril9gd+1+LTD5AXwWcCek3oTScgENbHtovRIyMqvJxbOqSN5/h
s7LZiusBSdSXwlgAU2u1dyN1kctGDTU5113XVuxJV/6EN9Xmc2/cOa/OzsQ1H2gQ7diS45RrThAh
V2KM8ZnKx6cgBnB5EintRataMyOiYBdEHQ5sHIPDOnEKqDmJTXGNtACUckgVE/6+uMpM693s5PDm
1KMcUzsfGE28vtAdaZDRAR2JC2oWGmCjcMV3EfZTQVWj6Gwu03CaU++pmdhOn0/3GyFyQh9RM4gG
QitYlmBrYnjgufHqYmrLfoEaaq3IQqnltqRnD784PH7axooDvKj8mGe47fv0hkJ+MTjFGctNd9zL
aZR3DbaQk/gYHrWX0/yUHi5u3yKyVrsMOYauPSJGnenYkcCyR2eYu9OXWSXEwDtK5q3n7a8TY2Ng
uCgl9iDK291/iL6mIa2wPb1RZSGI+AodY7uRLbiVvjzePmelVUnzUyVZLm/hZQrPILOhjUFhYdfo
5pDb0mP4RtYrH6jSTsh8+PggvufW3cWsyGcUaqBHpJSKDTYOIdasrT/4ra60H4odZe1v1Syi+NrG
euxfDt2UQ2orHEQrZUxMTPwa8aNu2a9Jfx/aFC4sIQuIoZStZm13Wip98G87Mi8l1q6ljXBu7yV4
0DCncuveuDHRchYOfvwkYQgRi8PF7pmCImLbPSdD+XahU39pno9YN5Ywj4625S52nfD63R42mnsO
zlzIcwf7x6JrK13+mNkYINiLesF7RgIs6646/TW8ZzR2Ewd3hY0NFfNbvXXgYZx7R8xK4ThNqjrR
t/fxdWTKkbLP9B/PZjT3i8pWta8JcwEXIN3/WSA8or2F5l34LnzAYFwAPOC0lT8FbBizr4a4sfhr
8G2dsGKIloo4aofxk9iYDO7kgh2XhQyVLMeqQaLoYipA6CCcdMsmVM7mLNzMP0pRUc/kym1olqZh
+NEKAJ9HT5FTFLPlgZ0FOa1hwVyju0jC9D9fQSFJIT6Z1MaK3F7rKPt6avvZuT/ZS+uDkI63TlTY
uX4uP46JbNEwoRwOscEN+REVsS4GSUc2gzvKo7Ck+61ASksMJlxxr3THBPycQMhLLJ+RLA1qLk6L
pX0lGZjncRNzMrJstERKM/aAvKT/sw7DhtyeY6TBcyRTA+l9A3ozdn/yfKA12JHwzjV59pndJ8co
wuoNa5zNLAvacETep567d1DWURYOb+bYnGGTt9q8MfiRjFHtBDuyzlPi+6DoMjft1/Gw6WHqJcxm
N8IVlOqg/LIIhx5J4tLLrdiuwgQ+7P+84doU+ML7MB6/YgiF03mfAxEymveoSFbS13TafbQtCTFz
qs4txukkCE4mlvTP03QgYE5PABMC1r5jiQfxgNzk2lVIACSNdu+ZKDNyfJGhVcOm/IjV/R0lOqfZ
t6i0LeRLNKxYAnWryQg+AjFSwFDbDxOrdM6YSrCReO0amLVN+E5AQRtDPm/ELIJ+bE/wpNAF2pra
YVT53SpHdP0fodRugJvZSBTcHUnmWSMYQlay4ZyxpO5vt9pGufymsvzoJuIXgFKE4+hwcUdWbuSD
m9KSUehLIWtThJ7O+qroelqFawlDcGkEwG5aDZcVIOyLKm5ytWjA5gxlVNglsXOjOfahe5zaMR6Y
QWEZ42KZFmfIDe8Rcbus3Tt2RrYHmUtnZApOe7W/lAj/lpw7OruvONnj04TfTLxQ4712kMVKH+4p
6Xd42/hAfMtQHSO5HiG0VLNbfToFbLzayxY7rtFIoo4OoWJFjxD2KMGELwY4u1mGgdFVs/9p7vTz
VePwgWK9MaFB8FxLNaVBE8jQxV1M3hYXtddc3ce+8ZvbpUTnsM8AwdDjRCYGwGWrFc49gpgIKgpA
c0ADecJSQfewVRiJCowneom9i9Yw6DwCWWAFuUSls/a55+uYx4wiUWHn5Mto+NW3zDyucb+ISwo2
5BAVYFwV8oMRUTFYjJIUE3Zo6CjqV+XRjJDf22twLn44quCY2NbwOHN4VTJmzjNnq5GL2SALmVlT
e1HRp1KVahesJnrf1YfF1cLIOIUHQ7KYkHACVW5vg5MlXU1vybMQqtzO7+EuBNGTPcmZIeeNCwC3
werR96wBKd39udQaQ4yvDskaf88QH492uzYQVJZF9Pnu6hpb+UwZXDAaE1ZUhjYvfc06vsMgHIFR
1lodVnUv8fxyjTSQGO8KMXztFbysbnkHJGXd3lJwkDx5uS0Uyx2eqBN6uK3HdmQ871hWXxBaqqDJ
WZiBk9iZvWUiDaBZqabwAM8LfPXDgqygjrhGtCyQ2X7B7aGaC0UZXuAYD/W0Uz6l8atYL8Vb515K
3O3Op92OjK4NH/MkkwBJGnb9ihMljIMwCRCSh1bWaDVi56cdGZg5cHWt+qa/yiSlVup5zEHiHZEo
kZKx9On1YUyrAIToUaQQNzJ9737gED3IJCnpNzgzcTx8PmfJQJ+tKhN4vrbdfoKBP/tvhrwlGZq/
ZkDf0KP8PNdGP6P4VnHRyGGMz5bzvHb2vj4njMeKYJ/8744jdijOkNfp4lQ6NsV+3I5LiK4URapX
aM5LcJI44UY4glHwnSVh87XArOO0EIiZF7eS3+VyNMrgFyerGRE20oTUIcGjKccHEOXaLBDWbzXX
YAlqxcvlgLcJummFISFSp5K53A0dQKzhrv9wKBb1TdcHuV+yWtXnzj98vsqSQdeR8FwHpHTKsLfO
z1jJDApPQq0Kdq31O8G5lUwUbxfMaFr5VgrD7VGrl5ugL18aBBCzobGzECz9QF1jShBEB9X0Rkga
SJvmfbsAI2NQje/lbol8eCavYls+nP+/mMwM3eL8zam3wSYs8zIi1aE3tGvuG+gAPVIHEgxf7g3J
fW05Zhu73ZWx7TDoHwWMgGidg/rFfkE75nHgZEE1ur2gXgYMKHlnVkhcI5YjK+pZ9ecS8uVY5tb7
vzdrkbIz+LMU4YdUAnuntjzEkuy+yFUsQh5imVY+uwqe8UsNa1PJTgcwCwn2nPJJrxy2/z2fSCae
/b62TCcWkJWEOF8IcF+NwHzF5RrX0VHNujvDPcVeZ9JqCrD5gPpNzC81ThQp3D5VfkFIst3xxrKl
gqlZ643u4yktTFwx/FSuqSM/nNxm1WU0QQIv8awTJh3PcUtBXk+VmUbpQKbs6qQt7ICwIpyboqQp
YaZmPOxskQUnj16BXRS6S6I/DnTn7LkkmNJSyi18yWT4X8Nycj+kWymQgtHS7wO2Gz37MfivMGOX
McY78cgwsXs137bAZgkS4xn0TS5dvmfrGpVEOxtcclkF5u+488ifBbr2F+O3r94eIvMOQSjR3t8D
D+qxuXbBMrgpW3ZXM+1TBrWonLL8XBuQgPr97iFDKBwtkDfkTPRU5qNiAcungQQgcG2SkaR63ChD
ZGHZCD+pyDXJHZ3tyL+GtLpKQ/UNznfxFSJbqvadoG5vCTvgB/X+43Yz7b5YNPOfZ0op4nxNBQU7
nlMEnovfTkdO+7NWT8XmlRx6NWtdZ94RfNtcFPqZ0jnBSn+cnfRTKY8awVrwNs4yEvJh+Paj1Wkl
u3g97KyLk8r1A6JlqDHdQ272k/MdR82qDSqz2Xkoho6QzqJbTXpKwtaK0IvejwYlHT3j2kkp0kBP
T5d5d0RhCVKhQ9182S2VxzGxAQjSKiHbZXKZA6YAc9ZUmYZFgADEqKwIXgwWZE6rHwhLVxJfKGFD
x8tGmCQgKboQfzFmi4NOrmuAzYc3RpBHjY+bd8niDk8Xec7+88WBXvPfP+DqlwEtq6WzMC9+pPGX
yHKixDzljkV8KBEQGw5k4iuPZToBaG8hL0P+KdqV5lMpHtUsRDZsE8ADeS3wz/oy9ox58+LIkFG2
rROVn41ZpYQ9vN8hB3GqEZVyussA8ApORDzYL5NGtxzjeXnZ8wElbVHWbuC78lD+zYzpwtpFRUSJ
Apu31guCO1/U4HaBdjXFuowoSqzIGjLfRdHjcfujXyUZ7iLB1EoWNpXabcxP/k56YzBfyJbYxQVB
waunzis4b9OuGHiS4R7qY2GLyACHICuSCrcdg7ShyqSyLbvyN+n1O8TiHNH9ZCutl7nUtgoJibdD
rXn3BmlSOtM0elwGmZ0iwYmK8mKcLvMUC5LW9Rt9L96bsx78hgADsP4jpKWz3eJauFaAF2W+R4qW
rtUr7JJQR9RVMHM/VtcMLpJnfpnZKRUliUz5xnL7M+G5eRXpC6848O8e57suXZex+MzwYYRmBzWj
o6AxxR08KAbcjI679z6/Hk7g97uaISkEjF8f25XPVs9he7LkAXHKOutGsfrGCLidAlIPXGNa/NQ9
/SG83jZp7JxCifcgLC4ewt5JJYfgK9aVDHf2bnkUhpXot+P9WWWs1CGwKMf/7549n805hErIEAhg
Sf9M4ob0B0Qa0pJd7KSWYz/xwgQNtTlIWBr0LYJepPVdEzk73IVcbUVLrCvMccBKKSjUVezTsWl+
pvhzBFAvBNdEkv0kTKQaSliMnIFzXfFcFhu0G89s4cPUvBHVOY2ZmoQFpuH5pi6WcmdEeNaBgY8o
euw1CZmbN6Wy4kj8ovk8j9RAjX7JTF7jVxYuoGOGf9V9RPdKbJYIXU9fILSGVYrUU46PsWdNO4PA
Urkn4G25BGeLfaMUhYpfN8JH3uXDVDaE49s9cXRlKlbuTX036Bnb+gzANxrpCppDpD/5lmz/pSUa
D3EEIc7jjNZ9AB5kp/Y/CNLX3207MwWyHWb/ouQtYQNQaExvlZvue+sR8LuPphogF/xASxq2osg+
RY5czod1kuMnfVmP1DAkeBUu2NxfM1oikaD9h6FbSC1Q6b/LBYqCGg+q/zVNz51Zt9gTsk9Pf12P
YzO859we//3Sh1O/M/L1l2lx7G0jwP4UIaZVmdamik65kl+ulwr5We22FMKDa88w/r4XUD/0gXI6
Vcc8xM0RlSapZrb7lP9pMnlFX/2BGfGfZa7ywXcA7dFb5OtM4aSDqLnb7vwBcweLAt2LDSz+DpKp
KiF/Xdg9QwSnD3U8Gfkdy4Pk8WwSWW7fP8bo5lrwxuw1QoDWz8g/Kja2JYm+fA8AsFKW7TytP6dR
Iei1pEmaxaOj6FDeGFkVzQpW7ekqM5Gqcn4kEVFWuLDXBhzT56r0KB1ZMPesTfRGFp+4XS7ieYxN
kJJW2eLxjquecexSF5BZ6FzVN3lZ2Hpc0UFo1Uuyqpeclrp+IZiZmr4IMX7+eo7BoO6YJBC0bXvz
KWxzW4pZofnuh7V3zo57CWHCAryeeS5rJHQ+at7DTv3EMTRnDrRZRoSneHB5MijUKE0N02AQY8re
NYhkMB9h9ZkEzuu7Mv48QVKMv1fayWBaxerkcqxq1RikxYe0z+tZWCumDa4KNkmVSAyDxRis1NgK
7XEJDzcqgJT/rXHAt4ZD3+ZjgZWlGNdlMqa7d87A7ETCYpB5r02YGTsyax36zSzneUGtCJcdiiXy
UYBRfmSQXegMuGdXCp5XTCNuII+hxbPnxwFEJSp1ivkaff56a8rhHpdpllvrovgu7Og/HmDH9uAL
EsmerZwFyzhM1Mp5RQ+9CErhx5UF/zCmu9D9IUO8Mhg6jCVi04hbnpVVF897jyRYOqCPSxlHBpIR
lybpPo213z5R0qjHB5OjMp86IHMm5Yf6FWcAbm3st1hvCw9Y5IGK4InULSlfB5KthGPMx+BHS4YS
vKp7koXZVuHyL/gC5uIwSXUmUUCL8AVuOoL8HNLK0W18veUmxfE4EUWhZLu/fUwsVwNTdbzTCTyB
DekHDKOoZ7vh5x91lhH6pBX3YbYuUj0zl9KOo1mEk+X+gFv4W8++a+DyhNuUVCmeO926FfSWuuk2
9/fJFI3gPImBunSG2EDjsHl+iulbhPlchWSGJXKh+nsXDZs9krD4t31hVxAg8MfGJJdRaS1tQ42g
s/OUgPtlKTF6WQWSakY82KmGB4qZ0baVvkUTwcMNK6AkcTn7EHsaHvPzt3EPstndaK4RQmdqqOXP
MrAd/TEP4IZIeBa7IEIrbKpOuNIqMstwEKoHCLaynkp6aPnQ9WGJZFTd56d40WG03dsnDhq6h61G
+sQ1WmlzKEvuErj5uI16Vn/PswCOS7RlWDA3BGtOkzWH5nksOmBUZc28w7/Q1oe6DdakpYyeJ7th
2GKg4r2747ArzTeipUFynDgNiEeF11sxoRSiRKXCtDRbDCGjmD33IyV5tWjIh9p2HJkWuj8GzAg6
ZM/XO6xrB9hiapAr/U8Hq3GXOqxRcnZ8+64ObGqzACP8Y3XI5xPBrWMoQFGBvGsZOk/VJD11j6a8
G7hA8TxtWZh7X3OFb+Fg+ehUW7kxFRDoZPCRb93sVYaK4m6Po1Ye0W9u3LMib9E490+GO6wqUxW9
5i3mFn1fve9QxgRGzyBphAy/og686eU8cv+4oLMbJlqRLW+c3GUnipcYAuhrs0p4Oy69qBvaTiGt
E11+Dh61rHcP0uEPVXsTi51dbd2PgWQKoPZulWo2Jk8E2RUvVve5TFGArApZrWyYA4vN5tAx015R
B5BaHzFszBTwLei5cyZYIkQLGVOByNMRXw6GTWAvj2lJdOmGIV15kzcZgUp9dF35P+wgRhTgs1Bq
NdcncvUdoZ/dg4qnHZzT4AxXZb/EhGJQIYVrWVmGMq/EHoBHd0a89/I+BxJdnSr/9FGxOxkcKdSv
ZMYL0VHk+liko5vDYQ2lH1XCQE1gxvoxuuu2V9OarQGxYSQrcdfzKtmSkHosIYuPiZv0m6ZoERee
xkkaJOukinLq9l1EJGUhcQNmlE2dOuVarlvGxQwFndecur+2sRXLaT1lqgYDouvBOtwTtM7CRZpY
g2HaBtZvYZn7Yt92+HDF6PucB0+fnij8q/bWJdFAoy7TP/wPC18drWLLuWL6fxXyMZKx0tnOBfbC
3KtEAhN4U6ngjl/5PCeWTzyNd6EY3xWyMxINPZEPSG1ZPocQhd8YpB19kscmgZExO6tQHBT143p4
M5hPzPnysDof2DelrwXw6sWxEpPbe2igTEWp3hwy5S29IpPPe9qAP35WDClaYmViFHv409XgEBLW
bKKfrC30M/XogBkQLUaUI6bx+sjbjeaVdRN6xUGMSW4wUa9r9Lo3RK5YQ7gjFfppGuRU0cUT9z8z
NR19fPyxlwx6ex/XaQZFePBf/OHfAEbNVkN/5ws5XBgtM7+6kHCVQ1ajI+tJE70/8uGYoknQ8h6m
2N5J6SV6/XhnBg1PsTRT2mxIZvk+AeN1dk71kKnK/DpkYjzg4RjuHengDs4CPKuXlNL2oWzpFNek
8T/XS0itvyVTRQ1+OEpoj3Lc7CifSxPHQBdiEO2sTNIdt3zfTobhuEEdDHyocyxcqsLvVN1a4Nt1
QsNvJBX8ZHPgdemfsrveIHbOB1AN30uNsTNsKzl0aDRw3WrJOeX3uH0/kw+FdzQJfTp/3qyNmT10
aivl8J1hfwSgHu8B6iOegqZCzcXFt3/gBNsgrlOH/O+w79lYDRdKeEMJKzRGGhGA4tSHEip5S7iJ
mTb78vheROkFOSzkUoVBFLSNNTWdDrmztP8zlyKCmZDECqTnqKDhTXEXIeuJwwlJH8cF9/q8AiQw
gEHfM1XaObPxbH/ipQSbWdv0eCX/VhNhrME/PXg8/dv2lujJGxt3WBC+mB46P8BjHWozpPn1ZqUI
ukuLy13TnQCJFLXvN8HIDUDo9uCAHHmJvQcC6LeydQ8rZCXoELjl6mQ76XL097gD/MVeTFwEMhTx
87M1hAVFmIamPrba+UOOrWnNel4bubQD8sNFH4uZA2HtuW26d6EPlhhgmRLfHEtxF/ZbWGwcvRf5
Hv+lM8oDFZuy9Dkx57iKfeGiZXOADGxPCE+SgYjl9UzFL+Re1rGsBGoqjGKBDpX6KUXNc1z5llyx
2KtdUklGaXyJeH6m/BiSv0nUZg/OwvDHbLt3BL/fdX4rqP8auUTL6w/85JXqR4e7orlCsFvtLhOI
6/KMO/QEpwOiI9SU+ylTqKyFoOyDcln8MFLZSHGERr2+rJzlCAFhQWt6at5oQoOg1L9T9gLObPNQ
dQWk6m4NPzWxGLUEFXISQZ+p+wFczAXcHlhHa0y4lAbAnwpjxjCExFs9gJpMia7LvO1ukrJMtDfn
l5t1Jd/OfIBGjEYSysCO5uTdC3F2d4zEv3ur/eCKrNpgTk2muhJ89ublk50TlsdAhb3N0ziXSLk2
vgLfTRGFi9RnuLl8/Wl59syk0vakwhbWa36utKGfE92bJzc9UYQHLqhsmt0D6yqD1geFevV4QHax
f+RUyAiUTQMXxzO2G75nJW3wxwdDXR+/JGlAzIyctVBtEAUB3YmPpT5tQ4cnsttICoMWq6If3ZEA
ePZP9KKGOwFSz7foKZAnXCJ3pUUTY90Li3LyzC9a3hknqSy/yhB9rebin9tRfKYEeqlx7mNZ7Kji
qRJWvTqAQ7pfvvXxVh1ZOOXCn9nvcU/mm0IX5mvU3on4LI7AWlg33Ux7tq2261PtchNqSV92ejp9
7kWxYncgyJUzVKUvn5sxWxdFMUrCXiRsCWzuonO+MwZvwiI0/mGewzCym5NAWuat/iubuWNjHXoY
0r7XgURFmSbNyUfVDbqs9ngxk1CRLDMXnItrB9QXsRMcpxhAnUYX+AO2wBWxJj6RijTzoHIapXks
UZQ/cuFpNFYOj4d/75QrMNF7qDNkIXBKN/7i8bRrWTo2ekU+BwHDXcYkXNsZV9BPCuxIjdxjjp50
HrOSSNs2FaFhgaZVQwSfzRabGX3JZOaVpCc+bOInTM9uON1AJ9Qi1w85rGD+YDp16IZBugliiP2c
WteT8023M/jriXufGIwrbPJhBEhbPzAbcSslgsgQwxnHVadOu8kqHlYqqM0OlFYhim19BP0jQEVS
jbVd35OcsvdMiZKtvUPY0ycmVYPIVmpYx2xn6BiJWQ+IR6MjKvZxiX8PRmWs0gJzrZqSlmdHuT9e
Z7KDeNw2O0ciaG4ktNsUCt7jNhMtk3v0+SPo+twXobNW9llcsuTe+qYGEYxkEm5m2BgKfUT/cZRI
CGsECi8l4HwlFvOmcG4RvMEsKcOjMcJZz/DSbUWHV3x6roTxJRobQncyIP44nXrEmFOHwYfjtW7R
T45WpRGZhjjpjw5lxwVamwenFgjpVWeZCDpCG1RID9IrMckyRRJmHsvgcOURUVSMH7jUA/eBe19s
9OfkjcCHvKI2qW4LJuPtISgmB78mpBmuDsRyfAE9gqcFz7Gx1UrHns2xjpw3aDqw2n4gFsCjrHCW
2j4P9cBRiCeXrSDz5G++8c9787AKTyYgk4gvbt9Bua9I+/aBWiENTYcZKGmbWWg0VHrC+ruzzo5G
0G8tsi3lvLckclIpPBneTiRlYNnkJtfb0fqvdUD8yQQkewAW+0doE/E5VRBkqMXxweqCPwCmyUNP
TCbZESkh8h6qGDwOh/6ulQE6+zy+phHskrRWFiot4jQoAb9ON1NoTgh+vftYVuar/aBhFzcssEb9
iUzuom7LaLjMVHISlswR7YVQT9MagNZKfIMUgcePF5Pgckb3NiFxpvZcXHEWGsx+MQysgGebW1tG
HjyrCl752dFrh5ltWzvel6q+1TNTD8tcRVekPDXa3wBjdBPHCk4WMUa3YFythNfkyYXR3rAL6ids
Wb2vN59liW6ExeHwSZKf/M1NvmdXpsd3UQIST10GQ/+JP/YfT+ksJfQQbwZ6lv/LD7O2/EejFWcC
/jKWj/PVfYPdmyD/VnDcdLuhsXnKL+1cjPUM2uVYx8+ZC/Xal4ZhxlXsMl2dyCGeSnETIEPMYagO
SNPFRuD9oT8PlDxl1LgbKWFmHRwj8iHYngcXP92/YYptxG7khvWOpnewwaG3434cj+6fefIAHn1f
sv+Uf2l6KznSp+8GGSLUSCamZyVyRCbd+pkISDzoXIYYMZSqD+3IIYp1ivBKTe6sqfVPclL9T6iT
DCiK/X/6vfKsDSwhnw8hfO5pZGaj1mP9NysabPR04L3tl5ANiWOswzq1Su9P+YdH/QWfr5RiCG4k
kPuNYNrKHqCTXv3AoLMY65v0zBYZA3/QaTREUp9JUBE0HchCwfFAqGRdpsGHXbKWfPvjQHt6kUaf
GVuFSG48Y6qRCbZ0dD29U0opbLWY1swQK6SfVwy3Yufduk7FYu0ZyuZyx2iDZvfnqmqhuxXATln8
8r9nZSsOD50FPC5uWtGfLgzoZUHyvy+nlsSprOaZ+j9wJaWUxExClSiqZOtiTzkYJaZ3MjMlwpDT
5WSSK/SkV8vXR7NEBMPHfYOSqezCxK/cdhrJDBs83s+8fhuzMwZYnOHENJJzrr8qhQidzIbxHI3j
uzLYPxYyk+mNj1YUMtnmLGaVcyh3VC86Uig14Bj54AxPUKLSrxhDiFdh0t0l61uWSQkbjtki2i7N
FQ7aXzoxFCeV9TdWPSklCtVsrMggwnXgbG6SJKyFXSYIgvLfX2K5mtSEsV046CQFBcACb9ip4VIq
Y/HT8EFUvfLd0d65qsTke2lEgJ+ZU4680dHOFUld/abd/4TMV7gMFVXwnwXL4kaIEebmDEsoTZjH
rd2LuIz5YJCl55rO74cFuaZNMZG4DDRfI83egifjNuFEBD/PV+Lb4V0rqMFCUHckETvrSp4IbNqS
nQz6rTBIbpwsBKzOuVj3AzBEGLw82DbkoOj1A6Hv4D/6Pl0f6PGGgqEQXbU1VaW30Zi+e+109LUp
IXJP33E6HGg7NEhdpxB38ZaYLc+/jzYup9DvS3BA+ZXCj28jjHcUq3l2YXOP8BM8KQS5wQFZ8s7P
QBaOvHSob7O9VoQnyEzmsAzmJ7+j1XlK3rtauLtmhGLJvXypW2Q4xrRTtXW1JB7cPXYFNAY4h4VW
4GoDknMaCvZE4VZr4NSMm5GahXVzpFYR3EcXLqLCtpudraFUyk+DL0y+7SqNYCNDwEBnxFceJto3
A6W4pBgedNGDdUD9ie+yNK69cmAYBhPFrLLkkLVipf3uyLsOs2LEvhQ/zbvEpK81TS8UheBJ5uUC
0pegC6DL9QfEobzEsKwUc1R3BmTAJH2bP3jbhVQZkro4GP2CtKeeXN6RN4LF/ppQuNfbJWriWYtf
JxRcTPGyHxOerkSV/KNvKMTNgdzEhi9egxKsu9/7wfsZkwtuMyE7wv5C0mEjKqAbjuVbR3xRDmeo
nb52lH93xHZfe5HFKRbtNZcMOliV4Rn1tkrBGjKRyesXMCxxJhsth5lZv3xsQatZ46HVkyL22uMc
aKtkPK7tqqT+K44LhOy17gux683DiN2jpGWuV0EWpEeWes4ax04+v24SG1fHHx945uQ0q5bT/Hde
yHSUnoa1cD3afJetBwEZda81l4v978xiw2Y1z+/i52IAGO7YTtpk9k9YFZlxb0evXFJVqyrB3uEz
JMQG395g9TqDjbIFeE8FJu81jLoCQTUQCyjM7nOdBkDdiAcLxENAKHL6MgkxKbxixKqw3rOI2BeI
y71NFoeoP3RHMGimgJU7oSglAHNvqZlS6LoUM2jmeA9mHh9y89HvoTu/MaekEeIDJLcQYaODl34r
h0N0tAHZpj2DyJ1uGbn0R+nzTLreFs8cCB0zrt0Os8H/VkAVzRKypOjoTuim386Dgz444H9AXwlF
44dtq+sdFTauzZShbUebyIpHZNqvuhngQMOBbeZ/PvTzKIexuVyVpwKcckMHq+76j3LQ8/LsyidY
Oe5Deq/aqCo3c9KB+ZjbGWhpjZexdHW7DT5xSuslkTxowMXfqNIO7bNjrj2G3am34ZwFRkw27pSi
7Y6H13dwCugihuPvD0IWgmOK5NrZOJ2F94wzhL6R5+WhsyRRL0mq7vAzjnwlvMqEP++ABJttRO68
yGTdfSUyJs/T/MXtc0iL0u/lAWv9wrt0vGg/fIR9NoE1uqrxer/i626VXqdiX6+fqOs4IONXwAiE
4AgpLyPoGLz3y79COlfboAvcQspyB95QnUEW2kYILMQC+8jbGXvleIttd/jEEvPWHfbqQ6A4bzjn
EFxgnoJYUTCaeRdpggje7D2rFHdXa6bdarYYzyG0j/HEEjB3dY/2XDpK1pphUR6dw6ilii+dhMfo
Jbp8asOwhEx1B8zL9rDKgiAYY+JGMQaXBbba+XU0kvEbNr9oPMaEIOMaDdG7trarQh7Nk/dITcEn
NH/4+alFmWk0iYMEbfC7iFMEdEFXZk5i3EDF1tKr2lsrrpMq3ohDNhUgFn8qg6fMGMxePJiYZxYp
hKMYgEbUO2KvGFyfzrObAGtEE2eaCInI+puS6+PVlSop8nU6fxTiShdnKeauKkZzKeBQCsrsJx14
rMLwsnAPRYhddyT0ho5wXCSTxP9S3pZlZpT+aYGDPqu1uISWJlmQ7mxDpSrt7TSQgtQqSOr2WMHS
04s9NFcaUqadoISKeS9+sNxl9acJPHSxoOZubpeuyWUHubLbrQbojyI8HWNhwgzSaWx7fuZxA9Li
WAVKs/GRuNzHBM2mX5OaiYcDOn/dBAxU4Y5e14iThsH+T9a/9QLbxp8pS+s+VBQstIrpx+MGmjnF
o8pL4/fAR8bZ53dOR0lT2Kz61SZWt2TVUMbkzBRIS6z5yMLeDPrg0InFxN1sWaMeoxVranNhz2IU
UUUwnAB8xs46nmwYWQnS/dzzleAm91ii8DaciSE7eIK8VkSBLoeCApsHqk0IW390f0bXqLAWVhpK
rje4LkE3uWPQ1bEfOoELM1OtJPQx5+sneyYiOnbrPgh4Li2FzYSqYYFyGvQlsC23wmt28bKRWE7r
/mdYqw0gTKdSI+ZVoc7vNovU/AZQRNbgjcQfeCcHbrkFo19w2eDiKoc10inmh6/ffHzOVdyrLgQW
+mViuDZB8X0TYkjoUeKX/YZZ1o9awJh/xWe7YV3qrCntDtfx7EF1SmeijmUfvp7NXloirEzqkgmp
8b09UznFBm/8/VGkemKKphBGn25qGfDbxTD23adOEjpZxXv+caULWqkb3N/cUTJ56w7rALYhoHjQ
wFhIb+nla3J08KjGFFy/MkdonELWdKPOkCFkpc6sJhUgsdIm0azAtETtFTIiUKvV5kgQtmb6eqSX
o+KGUejmdVY5wfiDP18l0w9DaCGWAln0RJbjCU7GE14TwCImtu4XuvpAXibtUY9iLYOrWswKFffL
UcJvFVW+AAdzZ0fUO1Td0JjKvL6/OdmYXIna4Gd7zA15UO0+NnotYGceU+gzSP6IEhq+D5D3YwRD
WS3f9sAlyeXtv6WX8Qb3D0Ylk0fXBusRg61Tt1OU/AYtw742XgxMurYoLlQCgaq8T7IH2dT2Bk8h
0MLsHS0w9/Me8YS6LJutkiN7ItjZaXGos/qaBVu299AJcUvmih8KqZdgAB9dTYIbIQg6urmi4r3u
DsgZIXeZhDzjt95M/4OhVplgGFim6nYzjMAaDu6Xcey7l7c7txgzyIfmFo8hadFCHzzXqGtZykbZ
Bmw8hR7jFsox9Re2cUOFS6ybRyikVaeNqUZRM2XwFadXgyjCimlupqex9ZzHSSvxtfM5XpLGil1y
cEluWDJWzVa4l0ov5o31Eu5WelpiXtYgTOq/oEoRxCdomIzESDYhivqcL69Su6G2psA3q0O3wTPc
ck+qqVK+BHF/AeEmH9FS8Aoz465B1eLTmrdHKn814kp19TH2Br6fyjn3u+S8MekaTUOR/ot4V5wK
pPqKKAZM495PIsgPvNBaePaJjFTbeoqTDDJM8Y5jn4tRhmTQMzP5K73UOkVz7Pd5I3jDtP84mvVL
bWLzU8SeHUWHB96sqFKciJdbFXGGJNlltAEH+I1Y2AGcoHMHR9DWwkXYlefgADE+D0BfGCW8Vroo
E5n6O/gY3SHs4WEmqdQ1qCODo0jt6rvzJf4vnG8S2bUrxX6iaLfMa56xyyeyZURAjg9h9qaJLscS
DGQiNJDPaFAbc1+126AavGwSV0mK0sZnwQboDtm9U9/4QKnd7c6+L68hSny1oMfx0BUqUt+VQY26
WCiI2O2HC4JXJB0lXHCko+mic26/VFaSvi3zMb8vVv4r9FxrLsVaCfnF99s3TT9Yi4j20ocWyKHZ
aXzx63DYtFbOD07QfBNjsBDuIB6kC4RdUfDrldsXjGnSrdXLVfF5KqaUfd3lwdyASmHs0VBDwc5N
T6yDGVaTTkql0w2jh/oivsV3qTYDGcb8tepy4TDK0KTAqa7aEnBobom0FT67cq+fnA7AVwvB51El
ZuoGXpuCAAW7FH8dNszungws2xJxzrUGCh3V3x3kPKWQFv4JUDiBSwVhY7EWyMW0wHQBmK6kTcz/
QbfpljMPq2oY6VKvu5ufylS5ne/l07jfgLQsWBe5UnD2IJH9MgW2twbdjVPiqL2TokfIN08zhY6j
9iGakQUP7g0dqPb6VAmr+cCnk7BIMTvXETrNmGSfbDotp8OlzywX7OQDT38p3JyMzgJtAoKkYTDU
GXRiNXvh/2LNGBvXgqOEt3se9MO1zB0hnJQWZpFbb782s5joN49JUowelhv+6hzeA0xGgHJ+RX+T
MgFEoKgW4YxjK0CqQrafNgn2fSJzbiOttMgjiNB/uJfIX/mJ5JwKhMm42Xe/gDbdTzNpct55yroj
KLlvNLP6VdE+tQ1jfaQfezVWoqk7hPe3GX4PuBNPhjgIz1i7H4YjeY+d3tJBuhu17x7fSOqAXpyj
ugYXB2b2jBqKfddssYa7Uy2R/zFQq5rN+3t/25dutpWCw5+Km8g1GgHrYSJYaYBac6lIWIsZBY2p
lxrV7eWhg+wxTm/4VkkCFYHlWa63xd003MjBaKqjTUZlRml6hszSTbNi8cthzCYwvcIk45oy0IRl
IH9dIX9nJEkN9ZLhGBP9r2HqJPEjbdRDDMVwlv0jnl91aqJN37CxUZKpDTjiB2uR4OYzU2Zw3LS6
HECZ5OUk42Dq4m3AN3ReoRLPjZDMyRfiDPLNz0POxj1eXbwuRdpleAi5dvvr1UgGMpfbCwNx+/bh
wmke6n4j9l3DfmtXUjWNDiJbkme8VLHmcf/IxGvdtgz0NkBYa+GEnCHeeENyOirO8Ye9NvTW5ASH
TB9mQPTb2diiQxuY31nHlbNQ9V5mbzj3RvY1zN27BXM4Mm4/iHTG8r3rsF6nIPKAyZjtPOiJKPC5
9GPvG6PQql41hog+Pwrl/Nlp0YWyjefKMTOeiu1GhiIfA7suFfIxADSI1MHHndaCH/1CXby+vFdK
4/+KA+AqhJk+P9MFJqH1AiX5Bg8aPTGSZnHlX7Ec8dZ+TKrVhpZ+PKlXXWxgJq/nmd23/teSnxpt
o9ymetgKqqm6r5S/jAj44ZXYFnbRbmS/MiBpwyRiqqE5ocX2Go8kUegPAgMZKq+xM1/hYBDTeAk2
iFBIPCYJlHMZKJKznGf6IzC110SbV0mjdNCA/oWbYqw5Ils7thH1AZKder5n/yTSOCwNe5SglovB
c/8Db0KUYIfHIfw/dJPRrvQnb9VUFbhwD5Df3BYz3epg97uTIvAvTckVayiPmHgCIqZXHxFOlqMp
0Enu2xkcvZIpYZMC1wCyN0pVik983eWeXev7n/zGGha/i4wxz38M0wErC8aLnT4xEVhbnaMdQkxe
a/bVAAlGdxgQEbqElydOhLnL0SCQtCgx+uW4Z38r2rgqJrLySYUXL/Bkl/ex/rN0kIHGncjIufPd
Z5V9K8/N6zj0L+ZM8SeQCn/mON6Ata/pJAnxzZsJhOzDM5JTQeVilc0a2XVXoJoi9BoOJj1qG7yf
jHYrFnLjSyO9cz3g67W8njoDCM2CBaZ/9X6jEFncPgIcPQbnjyJCc55PKmLBrUy6ct2TkVfcnuHP
UvAnRV4A3ALmSrQLKfxIEnkZUXUMdmI83uS9UulB9AwJrFSNCPC3jAW7Wk9ZPznQCyEgIQjPMpLE
yCGqf3VOEQg0NHYUUPAMyHRRBXdDD2oovaxUMYPDf+xg9l32VUGiSwPL34vPYk4FU6lsyCHHiQ9U
ytulWugmLE6G7lZGa0UBjKQ77tBdmp4BhOsniZne3WX42ox2jg5mGWLdOlhj3XmfmkzskWsuqUAk
Gtdw1ttozRM/yDLphxavG5dFc78gDJFkP/B+DVx+og/yOAb6cy2AbxAJvhU2iRy+0ylRTR2nk9lX
PLOqod5mb3KxdYX2cnN3FUiu4PsxVbW50ker8Uj9Hj1cJRQkPJFZfO+yMC2kTRmG2/DUmnrUE7Gg
4xYB8wNnNZRgY6KhaLVEJmuJY1BM4Zw2fwaP8T2q0BBOdMdDjKxFbwUXtOKXLUHRIu3/JXxWxdJZ
3+SLDNljOJCN43/Kv8msJYgq65PyRsmexEfOzcs6nYHMQ00TySE6Bm7qg+ou2nJXx8WF/DUZ0ZVn
TJ5QZuqJcedoPY+cdaIM9WsSariIwVXCHmYiOdXZtsXYw3AmKXrgkJvzBBRJju0liXz9p3Yt0YZ6
+9Tjj8cxIHcCptNJyIyCJChP4B5PmGICD5cW2xhacgn7FvKnnnJnQi5J84WL1ZQnfXXtOaIaVOJF
+H/8oloeA5ECV2QRTCfZg4BWLh6cBOCNsrctjozVvAN/BNrEtwbPCO2ThDooO1q995+Xn8gnIVnH
wGMI34pZNvN/uyhaNfUXCrJoRYVunj7evp+xLcIoL3zebCZuQsiV6+r1le6ePaMvEZY8gtehRrTP
9AqoY4dOetMYbQe+vdxkxh6RVQ/Cv6bAzoXeQh7MirvuNRs+b5Nv/Iu9+1snzKrdDRorwhSFuNdI
+zBDkKo0bB4hyTIzt26tKJgc/EYAAn0WKkyn18ctrrkBOtnSx1iv6QalHtd7RvQYgQZQCB8O1QnI
XIAXoX1kGJNIjFB8kgmMihJJb/B4CKmHcKPaObsbxAqUzP2kVIbwQ/5g+qqpTAoUmYUxMB3HwGR0
z9plSEudGUHW3RJsX1IV8pEQwrCavo/LD8TmnwBxz8/mVeY2Gp1ve2bWWt8UThhjM4uvBqpzDt11
hmdHnIJEcryzjaNqdNy+Q/vMN5xtMs6EK9GoMDnVzPYODmuKMTlnE2Yc8Fj5dw14G8T9HgNzHELG
UGbzjvyGTXzipZ7Qk4q5lgviLMhkeqhHI3B65x0rAVqodIr/AMgCEgpTnyB5UQ55sEgSBy3v85TW
7EvsfmAAwfOmTmxp5BDNOIR9Ik6mWSKfMZm2sLG+uiOtq56ny8vKLUp4en/acAuoxhtXC7WKvT5v
GNfSqtYAI8r0ZftOe7Ud8iASW6Ep80piEifrqhj7dvwJ8ES9vFdPKeSy1xNVqFPqWwuXoe2fs91F
QZwG80bVAZjDP8q3nLVEDpLm8P2Q///K3OYevxJxfTWFJWohXYkNIICisuLKe/XztwmKe9NO2l2w
8mf765k45kbeP/a1HUJS5FV55nOlnVs8nKAOyYg9knrcrKoxwb3e3H7ksb8U3MMhq0sxlDO0eK0J
kOY1oGM9tUtRsZlICGaw6v2PJl3HSoBP6gGZ2cat3WoQGA0QWqwyC92JTa1BHFhA9qBMOGuHZ616
9HgYgEyUnJmopim75DDuaHLwhOcmkt79uGcPe4kJExVr3qDLA1H+oZFD7LuiDvC0P+QK1Qyo3sgF
CSXQrw65NTZW/P4lfzjIoodX5LJWfhUt5/TvXKJ3a6LO+DL70HlDUIMcLSISCAs1UpoxB6qEsEdd
ug1RdpM0c4AKYMBIdkBTnqEP55WFIfhVqdFMtHDH4qCp9dPf/8aHIvPJAIIsMiOUe53oMNL7J9t4
HkdmqIQlGp+nfUf2e/ZtoNcGTRLcoX9KYSgqA3JKWeANd7lINI0XHonBo5KqnIapD32Dw9aeQw7z
dPOfXXHchm/9luOVKK9zKS3HTTxoP+wEVf3fyn3MQXPChCknCCz5AnUD1CVwVacxjHZRFU/q+RKW
kk2mSTxCLKFOoJBqzMc0ckCvNphVCLuGaxSLR8lkvxFlxHonDC7j/iy54LOgWou+04vaGpfylDqf
XHU5Ph8PP1A8mtisDw6WraeEEceuFsZrAd/Ye1xMWqUAirC3+SHMUwC5vkKv8MA1Ithhzwga93zJ
3GlwhoQr9Fnh/m9Pbm8mQyECecYxRrwoRqa+h2BMFX1qtM+HtAhsUALYM8G14lfdmjNYw0N3v7jn
dL3Q9bHBucVpVwhP7TvEidiQdz1zf/whT2hRJRxYpERmFXIn2uMOyo4Y9GlQz6aAM+NZwe2ML/OU
NyJcuIYfQxo3GLwgUGQwJzH/Jy+PGtcxMxpGRP09KVe8mXG9M7/sjuJVe7PcI/WrJXxSryMtIrsC
CwEitgRsJtTuKZJNLncwiLJeuyQp8e8DQTXGSFJLQSUeHcPDuyHPW1PEMNwiq4xc2aHKh5PcnG0J
QMk0CxV7DjeG8tF81NVkaIRlYKzAHbIZ4Si9YG6qD40JYStUeR8mvP8Dwras6oQOSWRNzsO/oMYa
fqxfrzX84xPnMTlgINfko75/7hwe0kNyW/+VAyUrUeW2u+T7bk/H/yVcZZvUqUtd8KppZk6TIecc
BX23o5mlaI8H/BVxQmNUxwPrW45s6u7fmHinA2CQG649CGlEmK+CdODf21mMoppHOKEPCYM+g/f2
zACch3Bdv29ufW/K9zDcOxvUNIjp1wApbADG2dn4OQc2HzLYTf7f7PzSHS++zMatIMQgwAnmjUDq
jb+kPF4JMH2TT0HcDv33NDVIayryjLWAbesJ9TWPhcUNMIlvNL67d2T3VixZ/mQzLVw4FropejgJ
l+n7xhY1HChwsJn2iksOvlQ1kUySafv6Hg7SFgDlhHSAEcbxOrZRNjw29l30X8KntMiPmduD527h
4i3VoScjQUKZUQnGvCtahDDxIrFvlI+KjLmd8acscBeNZozPNwpczl0MsluHihfdDdZL6SjLkkod
0EEAYSHrkWqHkjqAM/zKaphnwc7VNgqY+b5J28O8YL3FnKDwszChKBtGg7cJQuDAKQdU4g7lLJDX
kiiWi0+6prJRgm33qezToVaV9sqkhEGVdSf7IkUT4sHAaXc43h0UQUkXSDl+JnWXeW9qmgPW3S+b
/O3Ea6p9X5nXe0+fx+jufsIc2wjHZqblvWxeQiqFHT/caQ1NBygBe+26sKbSNlSy6uMdEZqqoqz2
zKKy6QUXt3BsCFO183wxTCWP//4IulkbhC8g9RPwQa5xSnZJCu7c/9SViinqVmMGU5/haBMFORh5
mQQMogZyPdECrewBI3K7n8u6FBp+rW6Mi96x+zdhfew/TEJ9FLb/gfdN+d/OWLxq/HStbV6VnPeV
fRHkeoSQAyKDvFECHHCSr5mXGtlnRbXXgaDHZJ/sn3n+KS+qP8V69TV74KmAvt2v3sAe8gquKp/w
enoTyErTDOBSsbFBlAr078vHdVcJX1VTSaQy0RHpaQVud3naT9pO3o6kblx45GWAqJMwebimnRTH
/LDDNqB48cxVofEZ1/IM638eRc+rHejMWdarV9USPF4wM8tiAc0ur4LFEW+wBdnMJHoupKsU18iB
huFfbkV2X4dHT+sCPv7S4BUpsPJy7+cyBjimWIj04R8GbOkR1q0B++NlxflWJNiLSf3OaDzfapin
bi7BxtNLfy3cK/KO2LFVoLAMNlodiSCy0eFSNbSEyyX4KUWHCCS/ln6TeD1kU/h2hz1mEvgFMXLp
UmL+rx5qYoLFOXlM0IniWE8nymiMlJ+Z39avoG31D/UJzwz1HtFZOyLMYfqC1K4cwzY2V0tY58xY
79xAUIiafmhkWroh2+GK0Jbv31t2ZFnNqRAKFBYAqbHnfdNzR/V/Fj6mlPpmQyhazm9x5u4atL5Q
PLUWwUXrWabb80gyC3O1+Vrzyf6fRt197Npybc8YMTLjmL2WojEGRypLL4xyXDf2ln1s8SSgxdyw
nCwBdyQSkci7V0lPwKNjFPsRQdfZf3OtaSKLsrYvA8qpUMXuXAs1ctSk54R+HAaXTuBvHNouB+tS
cgTYUnhAN8xObUTSD9lydzmwFIbDA/NEyiUPGsL3jHaHMgVyCo2WBsv0Z1sTQ3HwybnwJItkmiEH
qdjfiTGMMYwwPWfRSajjMKbNWFKT+UYXJXkP/uizq++X5WtREbo/LRnGc2Kjsb1S5JGROjVPFJXH
Atj9x+yWtX3jdlwXlo7KrRyAHJtIfATlLokFXg4+YxjOWGFj9lfKdcZzOSs8P9E1anGnE25OcfCx
tWx2mbvREcFAKY1GlARLKMdXBs3dieIiAyGFNm1kgOxNuqPmlq0m9RakinuI4gRGuL4rUOPs9bzI
EM0cJ57gv1c1BicbOb8WuAonXV3l4hKyyuapyqguXe0uEC3C8nOQLo7wSIm0CkpFa4QuPHBRDwTo
WAfFCCry85hhBkUN0B2R3HJ1w0icjWT0L387QZa5mij8MPfPA6A2h/dRklBzOSS5MVkmgBPNN0jX
0h8VxocVj+s4S5s3D3Xb9X4EPj9jD+XLNicO/E8zyaNWbSEqONc63zTqx7oLl5G6XoflItZ2EDBc
DRpx+n1ZPe5DjzS74BwgAyn/BzG13OEWKNfJRJGzJZKNAb2EI9MztLPLEp6lb5swNuVhhQjRdTwt
wENk03P4PnQyfExWAX49PKQl9buLc4uCSvHwoc6OzqMTjXXO/K2QHRvQz1scxWEgFE6WFrgtQWbi
gLQY+p6VRhENFImPxnOFw3YoL0br6Yk/HDINzg8a4D2sLb24K2973sepJMHNn7wp8emM7zCVOi4K
peUbw88LRGpLIMuCPu9emSl1pci12qmOCH2juZz8KKt7n+ISbCIgaUOusz0ixQUcvKKYlS/BdZzg
ugJe4nUQyXE6RZ2szyTe6eSYil8oUOPz0jQg1xZXIIlBoUPykbS2oR4DfkNDC1gc7hJDchCN0xjI
p5WcP2P3ZpJEziSBvSzaQz6ed5O8tWyMiDlJYm5sB1kxLVywcumBWi82QwIDC5Wm532sOYKTJppT
86fHmRyStgfAkDQ7wXnwhC6qNSE8G0qVI0EX1gvcsGfEYPzMAl//PfNEp6rW3eHw88suQdF7sQMw
X00aFrnNPFTVaTNNI5fyQEkpMEQtJKbTQIcJglSJc9HTOVylun2VIyvkFGuEhEWxVK479aVeJ3ji
5MrliSX6rIhZguybN3/d3RK34IMFvVipKhrRlbzO3kcScRFPtYLVx/M5arTMFG8TlVbFoHKaCOO4
aEXcOOVL3aMJJk79m1EeHGfxlLgF0y8QUYSqnu7pYU2z+bWuAVObvbsKDMV34U3hUn70HbTk4+kS
dn5vBLXpotrUyqSG/w9rHJToQ5hEbJaK7hHML5OQVHyKdKd/swXI5lKiXBix+Ck9SViPVGlZUAH6
DgGaXfgDcYJqylpd6ckCyprQs++INDDIASGapn3EaU8xNpQfiNPNU2ALlDkrUbU6WEuscEkodunr
EjUWQOyuqFs2B9X72mQoWIWpXRk1O4J75IlK4WlVom0n4qt6vGyNEwiq4XqLpTU5d7Ka1lhRNJ0C
eSMkEKx55Qohl6+dXjlmo7O+OScQHvsSZm4WQ2B6fV3VkQZXNsaa1r/0Q5vX6MqPa38Xgp1L5hKo
mMUtYdjSkQMXcb70MNal3F2Mwt3OOV4N1rGcZ57mgk+MGqbs6e51o0Qu4YLPCOI7Wwt23YIgq3+O
P8yGCYWekv2491LHEgk4KctLSTUs0xlbyqSRnyvaWQONjnFBhUUNWZEvHmql/2TNSQrA2sfkCTb+
mC81P2MnGU7Fh8E1AjvrzsR5RbpoD9tJMqdUfY2oXpSJxFZzF+qyRwNGSXd8C08dEdP46CwzSXT3
Fupw+JapSh0Zvbf+Nd4jbyrkBOOTy1CtrOHvP6lvYGy9iAeL6i2Od55zu9mR+Yenfu9+U2J43Nj6
WrG7qMBakbXd6+LzwvFUVPLUevDOzezHS3Rmre8m8VPmVDtn4JsWoTCpeLdUTB1Ya2Ze14eqoHGk
7VTlYuSf1dlM4/PmTLooTur2re0p1C+5QQz068594XPel1r0E6FrL7z5k2RInjubcuOwHOoAE5ZG
hA/sBqWeY4j9EtSvURtnw3mDyerHCs685YyUP4aY7lJ42hy/TeOYZkC+GQvyUzD50d/xrcsSPedL
o0a9J0fmi2WD6ayx++n38ejx/2vedVz3rRR3eO+zOa/ulM5+Xqt/vMNenjBXUd7ykvT96+t4HqZe
ISZPquhEvCeRdNF5U4XYXfrC7UQGzUfZL+dzaBglqZOwdPDUPVZcaqqwWcaS6TB4t/MtrczHQaUH
o8N8C26k2cwl4leUZM6HV68GBd5GTj9AI4rUILHVVibxRWmUXZvSE5Nxr5bQQdaw1Hwr0/BseRqX
RfT0IYD3yrs94YT0h5BGMZBgp2VCXtoTOPRTycn5sLbAzOShEw9oZszPVOOCltmSBmj+lwXYfqjA
cD6rhb016VqaGxhAelHJ4x9URubsTJWbYF/tl2hqUAD96h/Y1KpgizNc+1YUreXuTyy/dZpwZSqX
ehOcDHppQhwRqTUDpyrO9CML01lVSd211myp2HXX/Q/w5W6/6lIRxjBeUIpezQY9+nbF5CnOmrIf
NIzQekX4qqE8zgUhDX6V/trvE6FV+tmEc/ucZutfSTH6xVWR7N0E0mNcnVno2Evmz24/WFiy7Y+B
erHHQQjmvCCQX5NZRyFIvH3N0lBo1aalPQ7Y9tn4RkjTKDo5ilrhqSrIuMJwpufPGl5y/UA02gLR
5pa0vLjPct2xMPQvw2fdlWwFD8OSEnuTa0x6su6A3CwidRWPO/U1ERhRezvwx3+g5IXHJxA2Nupz
lQfd/Zx3uXEEN8uRrRLVwLKvGMATg2GE61qI4rK+BBnwdi/Obt/qp8igA/3cZWk1k47tcAnow8cO
COTSAMhD9444jenntpUxHq6mL9itUVhQfFhUoruNhov2ufzFkv9xpfcvTNxZKM41LcMLNrgE6v0L
+AAQPkv78k7CKXbvx//+45BAKD83x2QztVET50vYlNIhtuNewh7tSJKmFiNuAldwAMxNPkDgXl4z
0QLV5uT5aYyqJzebD/vWaSGV5KCE6BhxncEE0U2+4b4Rmd1dHXipgl5Vmkpk4Sxrnm2hBLOOqTMR
HpJTskWKsq9uWioigHkwKo62hgHd0AvIdKkJei9a/VFNbJlbbjgk6Co2KIxcHMpfaMzGt72lojJJ
VG4z6D9Xjg5Ap1fDYFantg70VBqQ9rMerlTetvLZwDleVoPFuDg0K4xAfqzRG2PzwddxmT8PUcGD
oOwc3UsfEGJ7jlO8auPZaY6LyIMXLWXJ4P9fvsGosv6A61k+2rfCIrXq6WdCPRCJfTbEAB9yerqh
xyaFHzUnz6dIO4EUUPF2r4ID7+F88QRVizvO8SClZ68wvZ1ug2v4XKBrJoKRtFHlkWPSx9VCLBrA
mniHERZlI9Ia9LnnEGdDG0XbeT6DsJMzLIL4ycUD12WiIdzgNiGyoCHr8vWXT2wz48h+c+bPuM6G
B6rUkF0ZVkFROGRKXvwb6/EskCmslu7mOS2Rd48b3TDPZLZRAYVjZqW0d2I1hbnnkH75SxLNQi5R
m8vN64gMo5y7h0SOo4UqqCVOCdKHrRZfjy/VhixCz0X20osPlp+VhKAIiWtZ/xW1RGlm2eYdaykW
qFX4OPg4h2UKNTlrQ0SpTLD16tqc26gKW1hdecOEIiJ/nETQAvUSGwgBtTgJc8Ic8c25ibty5t51
gH5DpSXEz4b7l5xqONmsDj4H84B1QrVLEXMDuyQXDJQvTKXWqzL0x00IRGJ3BxizGsyecAG1mcEw
57T9Y1RnrUG7Mbw9GVE3Cxt3WtiOzUW53Y4Hm6vJ2JzLJ0gEh7lKtnGJ2tY1uFeDp5r8eDTtZegw
uZ3qgyPtKsRN52+m5+g1ILZc4N5+S36U8J2pxn7CQydzlnQwPjgpkl88GuqRBhX8jp0VLZO5Hlo+
pQgxX71+/YyVtaRxu34YCr2iunlJHKjDbgVVhnlPYy70sXbbwu1/+BqPAQgKNCTkGymnuz+1Kp5w
pHL3/553HtsE6Y2r85iZTZkIhXPTeDkyk04FGlJBLO8MddmiNwSV8AhPkR752T5IT19hN34l5Wwa
OnDPFU9mfQkMdRdHwSw4CtL1Kr9RFb5HbxUosD0w+KHX8DMcceSq96Ipa0zhXUPC8vnuno9XvKbf
uZV8sBo5E6+37M5cAMhJbZeM/T+hk/D5d56UReXH10243Th0gAubD1xgZ2QihIKz86A86Xju6oQt
21fz+d7xy0mL82Qc0qI6DqhneuX1SUc/c5SCmRsRMWtl5tijfT52HLxdNTxR/5hHW7W6DCt1ZYm5
S2WGUqb7I+fsl541BrrPZJ2Xx/mQr2XC3hkIcOogJIc3JGnZWA7cSLukdTyUfvSi4uks0li4Zswi
cSo8j/RNXCQ0iO8FAGTbKxlBQZgGAHE9WVwrNCul1h4jEz8zGFlQouprbV6Oi1ESh5jTwRu1konb
QFawRznWVN3Q2uaj1oGQmYuM1NR/C/9TFeJxLp5nd4lSe7b8js77A9rcJA9IHHwzFZ2hTJhSsxiM
Q2FC6sBsOnN6bPqLKmmFF2FgURylPQjxKwOvtSYNIKSU2ncMCJ3K8+uTSI4TSxv8mIVV+OFdlXgd
l3Q4RCGvTN4RaXr1AiEEexq677nWVhAD5BZD0hWJ9r311TKxary2KlG+5ZGGyMALETF+ugo4+Ocp
xvEosjIoG00yiMV2Pk9NFBEbSlyytz03wusiBgW4+pxCV/qK5dUavNvCBqyl1CkIPf83qxvPZI6p
NordB1sU8btodXvnNUh/oGtpivgDqQZuFTyyU5CaUn2EK+lgvn/yrj01ncaDH3JYxyM+qZD1Kz1C
5BcKG4YfIxbXZgcKJRWtmH6qtoJBqVXUODEsgZy6WKNjzMfckdH4PTCnP2PXT9FK+PKWDXtapz+j
XMC6j3sIn26l3ZGJMKhD6vMobA7P1pLEM29Ey7o4KUzWrfYf1aFKkjGZS7FulHEI4c/Qx9JqDRyO
NqBMO4SNFvFZZ7nbFtX6ZHfyUq/tydl2CzzGu57wVhFLplyRQLaNgkdhsNmOd0PFh5wrBgMN0W+A
SciiidsKxiCzrRvNYpu7qRSWQNbeuZRaxk/8LSQ/fmX3x91ah/VqjCYjy8GAAg0ViA29GpvmjBdT
4901BZjvBCEen7V8V1nTtp2Tgab7SO+nHSKv0ixlGAKiIPD7KBpIQlgPH6FJUb3wtboQu2B7Grk/
Y61Vb7GStMUHle3XPY4j/sACkgKxYK6R0Gq+JPf/09p92MVejRvShO7CmAV1vIJa7NFO4SWBrmLQ
Vt3Oz96WJE7Hzwz4X3BlKiTM7gHMawJNi8j7OnCmuc6L0HvjgwLmvpqV0MOZz7MbEoytfP/VcGKD
hMmNN7lVYC/mKFOEy+h/YljaE37rDRuNMQV7HyWnQqQqfxa1MD1y4u61kq1ooWbEK8LsbGDcmEur
lsqCE49GTiucf/3zJT+7yPC8iE3u6Yf9t1sGoZeSgztViwVKPkjbJKKQynztSWXG9Z9vmRSCa2XD
MH1CQ4ZNKjCVs2WiGSr4NgDfIvoJusCl56VxCXKOf2Kf7jGXsrv/+8Sk1fiWWHbuNrfrH2+AcWDA
65O6HGrjLamz88HnJOIdpoW1WbBUL4Im7yqgVIWR6UBpOiz4Mcohp9MaoCyZ1RBRYnC+JGNGeeJL
VjYjERkGnGiQK5VOMMk+iHxq1RRFMCzDN2DxLpvrW2/BLPAm0d2T1nAEGxGKPzBWKg7tEmgaJTwX
HGSwkoZA21HNDmLn7gLXNbzvliq23dRNihvP7fTh/BpVH867kpc7GoeQBrO0n328Wsq4a/i1ZR6V
Ti8bHoSkYcjN5c2WT4jr58OyFauBAzqqq1POs1x2dbXi6ZGB+OUpOkJKChVMhBxBxbbnHacahClP
CqcerLVJZZBEJHZajKqHFnOPjAjO8XBjSXTzfjoM/bwKzyg3LcWIUYQQGOkG3VodoQp7pC5yFeBU
SD80WJPGB/y1wyatH/sPip1cFEYadqtuDS3Tx0/X2GYGCJZ3i+pfeVKhl1Kc9FAtRrCp4//bQxbf
xkIHg2dd7eEfmEcd3zs1HooigVAz7dVZQ18ZL/BE3XFyMBaN34sCjJEVKUYPtw+gqQO4+4YzGRZA
eV5hQTTsndF5iQ5rK9C/9jqpzl1xb7/z+Cu1QqJAqn9fjeTvMmFOIt6B0CIXp2+aYzCx1UvJGtzw
AYtqilYGMedVlQ5Oa0PH+8pIUguQpLBahZ7QBjGMSk9nsJ9rJ5BYxaCY6CN40KPwkFTKe0Q1fOgh
HgY9bTLoCjVKIUg4dLk5Vsey+x8wznos7ijUD24RMvN4Aabmm6gm9R6xAFCu6nISr+lEThrXOnde
4nmbKuIBCBrv/iGDRRhR+cSeiF+SWEhojMKPRmfVc2AXL/srRlDkrFSyH0q9kkTsI5Wpp+q4GxPs
TtPJlYNkZNXuLNMNjFZ70gaEN1umwQIhILyA96l9bSAmmFs6oHgYm+YnFPvdXUFVDb5T97WiAZUf
aw7KaZ2auzpRdKb30E7L9oAXh0M8Z5/Ux0RCIAflWmJ6yDdMiydSvmHDP7kE17Zt/u9ahZ6Np7Z2
p2TIwtga5zbFcUTFFUJbxQKMwjH/w0cmFK7O/51CZH1gMObtvg2TpRMR4NMQ+gunGuv21v2YBqoq
2Qs916RKT9wgYhs4FWB2fWhwkc/aVwPayaIauhx5QNODoKARRLo1uBnjXp5xzL9+dCjwzJ3AqgqS
XHNmMouTy6eeOcxxiR2Q1q0c2xoJnQ+vYIORgNOmkZ7Lj7STVpDz5A612CC3jr4sMr0iS+SajpHY
F8pLRA1tpX94V2FnA0XKdgPweFi1KqoVXnxcexk/4tfSi41rG7qy2wujl6y7mMKy+skBii3l1q7k
MtYPlPlxJmWv/+kVrBif2SR8htAV2nm47rlTHbAKPbTC0bryH72UbV45iPJfygoSI0LU6Bwh38hu
+E2Kq/Fw8vUf1PSXOfZ9JT5GE5+c9uCTRypH1116jO1So/X7inJLkc8k2JuO5BqYGmB+kJA7as+X
bQ9U/KlYcWIHdQ8Y54vwz+1EcTiievWbroc4GlOb1frZyXoEjo6MPm53G61viBRXMKeLsglKT0bs
31YLwOJrVBE9NbxhAz6D6m/US/+c5Dbptq8LtDTWQLMLRtsdVaS8njs/2crilSSix4skBSLXBQTu
xOlcXxSEMOdRHI3kOhvV22QYLEJh3B7+ErBGjYWwZpMB+Upd0NIYugTzf5wnB8v/6+ogtNZ8S2Yo
I+oLqhrWj8jpHct8D0efl+0pa3IDh931T2datYj+h7yX6BxBi6kjQwXP+Ze3DEVUWGfpeNHtPprt
z1KngY2JVba2VNL/wvGzqRqUIz39aDH/QidMFmTYm/xlKSPGoWEtyhy7wBNGGTh2Y+Gj3wbKc3v9
YNhiSXogaTdLCkO5uWgcO+ckNtjpoo5xkNS4ghCKcCucbGeLIJSvtJ3scaTEgk+te9+UJNUwh5tX
nHprgci+T2Vb+Xxk+QbsRCJ3nReDmzmqpx5tF6gqv3aQe7w8rl4L2bAhSS9UExJgURU7URuXGFda
MwuBMLokWIBwqUpDAtpO781Z4jwEORctngvYVaD+h+4aOmywD/p7/+/TqR9mO5aBdIEq6XIdVfWl
d8INMxPcAk1aIFJ1e4GNJrTkSwlcP0LZWV5REDM8KBIHfwM5MVdqzPTzX/OoaoK9TViG8kXH+pjL
f1E5UBotHlPDFj/tc3hBWMv+P96HRF9u0RaKhTNAyMl8K3V0YV1gq4l8Br4+v6DRckxrPRgfMB5C
iFep+dgtmhEGyP7DZ9Xswa2QC/fjnXhf/47t5tUEzZjAoJ5IMuEJW1TE+pycdPeteTEA9k+/H37u
+X6gJmYZT0ZMEHybm1sGtcd+nYUiZdM0qEYFm+DHdtr3vkvnz77pnKGXBkh6kdYNOm+5SjUxf8Py
KkUAuI3WN5yio+OJQuzBjbeF+oQOKByjnSCqMVMYYet9BA2brJxZiFIMbdfYFMF8kMfHPZRcUQtW
EbMNSYwFzikoknYdbPjprkxLd7Mb484OjZj0k26bKu6FIWDARyX947PUJnOLZZLtY51g3csHRmWA
cY7C1tiAG6vQCczl6HHWHUvde+09B1tAXOGchOtIhhq4lZEIgOkAjjh6pWvrhsLSU0NNiCqylNip
crg0EiYbLCWbFlNjTyLKde1yLMtPQdXsQWofYF6x2vwMpLgkEv9w+FaBbgL07QSUSTpK5KEUqWct
K3DSh4Q5hLvtESjy/JdOG0Cauctr1bD0mKYGnWGvHoA9rnyEC5dPLY3DrfL/KLciz3WkMNbfP4Pc
OYFi/Y+LDuZbBLPsoh9QBzCmH0CbLS/gKo9rB++Yi8LmdlubZKxB6y6vrJFS9BGkNgVafWyiXY3+
OD8nkQRHivGZfGbSMU4emWJ0uFn8i7xlU6kCoxa0+cDCH621EG1pEGqBuPix0cH+sfiVX3c+rxSj
Y/vD8pFP00bqNCpXyEw+mvdef7QmfIox7VD+dQB9SRvjQgU+UwWs7pmoku7YkcoaUg3zJlbVmlwG
wn7vAVV/8KAIQMjocFd/Hy/XBzUrK1RKYCxwKePSAQL+6vGyN1nQOzuwQCgW3ujXeIN/e7l+EL5J
V9lFrjKY6SyW7Fm0kvK0NOKOZqtR8qH45m11es506PLyIlH0umNVtJQzSSSbY9IVt8kaD6tVcceC
y3xbaBO+SKFfqhYsJtmoNyMGxwrqyKQSxr+kpYLHG4guUeXH0pPd9hDAgbDYoaCIM5uqdmsjZvEn
iH3Cacri6lWNkmgwXBENcD9n1Knutx4VqwwGyqt2ipS67519ueCacnDl9o7YyRIRxY/f9y+tc11+
IaMohPEC2y6rDPvcVYYf9X+KqXzD23q/OhlEv4qcSTEkSE++vLbtBuDOBxJ4hN3GQjtDqsWrC2UY
xrDvA/Stp251lnT2pEGN/rts6TEPmo9wWcEcmm3dUeFdFam6e1S7wvdhpHzj+hMGUgR0aM0U8jil
u8dq4/Cv/0YDDyz0ghZDHj/VN7RXyIn60Puoayf6bSGz/YPPeS3xCF+j+rCjB+3LJjr3wAfBRM2V
l8wUr41KHMpPPcqO66L8S0tI+PgKpc0+r+3OD6KFQz4RpsN80rue2RiurUKwUPs84Gw77UpNBgU1
UJqaK3OcbIOoJZ79FX5EZwqy+URxFwopxTWkWIV4yyu/kxFqVTTpKtR5wPqHg/91+gUhZJ66Mkpx
ATZbizQWuYz49Q2ymR4J8KzKnKVV+WwvuJlHyxW1B5lAP0XNr7Deq1P+0olJLuadajwqfP3pRFVD
d/MS+T/LC46swnGiNzh/25UST25JM89kSN92rZe2VkiymOdV41tdR275O+SBN2wAAszdyHTHZ12L
Eo5JYM4irxernEVkgHjM7Wq8Pi/U+U/kTWsSd2TG91l7H/Wqjm/vgaZlNXiiFGjueSAhRHflTQTH
d/sgsUw4ZwIkFP4KJ6sFpJ7GOZbiYzYGlukN0xvkdU1MxvV8zcE3D4WzN+AizhgULPaQuRKKcRoz
YFLtrLnz5snL0Se+SU6aH6HYZFKUNWP7PwA/CM30TPlFSUbNc4aRLyyE1b9+OV+UWPD376koX6rJ
qASJ60qxCQZ0nESc0ExDnK9mZpyhLQIejLGgSy2mP6P9flecLXMsXV2R+S4fqQwfn3EDnfg9f4uu
PJfsoJqCh7Kv0CH7pvyKRvm6fEnoSe1O8kPNYbyJWm2xDb9EV0TYZaoJCBNjOzfV0wrS3mnaOSJT
RG+AiZb1YzIXsVGW6KyHXaQAt0EGVgEPlwEGOO3c1UdPi5mahXp96L/4WTD+CAwCccB23HbOOe20
po+3+2cffwJvbBK/0z2pQQyx5omg/VaKUAOVnofelzZkYvgWtwgctRmBJlUS/6kcHlMOgGFau3zC
Qr1y8q+Hbo2jEIvDGrFxx4p7zrROP2ZBVE9BD664RlDa4d4rEuC85FFv6FMo2QJjTGb2E2NTfbVP
s28yo43L5VtLpJ32kvapkYonTz08N3WPrf0YhphPV2Q8oOZXU2xCEUyEsHSDa0WNGc0zv4o9ICPU
ATznGFXDoPI7ojDrgIm3k3hyt15e3Ufacgw6yoMJRMLO8ycuVS7I0u4QJ4lzLrh8FrrRGkLJwR41
SiSybvQ3NadK8w574UDCB7DCEWmEA+WmaFe4A2IilrTvHxnc7ef4BCIuC8yZ1Y4q8G2cUaEk0qx9
FIZuc7GlyZMQ518Uz+kOZud50hrjmTXvMZBHB9ETg2tdneTo+JTlJmhi3vRsnIwNXmfj7OmEr5su
RoAml1BqAYjxL/o5yKzUPX2YntFTuyI7LdNsPv4af/K+t3Ad7yjKfeux3LlrfD2YiH8Q2T0MsVRL
pKZz2z3N72HwnJo7TWNQAjRmeqG9Nk235pzEAJQW+FZinoIRwrzmdZviWDR8vrkeIpNwcdBM4ziT
JaKExIy6GT+9vQaui3XNJPH3Nmi6rGFlF9sf5LSCrc8UcIrNQ2zPzWIE927/DpH224zYR2Fc5v0f
g4ubNlAx/Z2Zp7FZYZ0rTySuEntIGwVTOzU5e6XzNScpRaWVK/lcptRJzICYkkEjES4aq2VVRZdT
0tCYXwVUBz58/y7v6eyNj8rIA8Yc0lXFA9LARZ2txKVZpjEHpLNvvvbKXHQqpSvoCi7lWQ6G6cj+
/SyOumecPCggFDM62cKC1FlFCKM4emR1hpo6LZSb8NYOumzNRf0f39OtrQqdC/QWB5tf7Vdxn1tT
nv+ijvau9OZ+5yXn0ykUUKBYUpJKqIKKQzXmhJJvSPFcr32LV4XNuf3UITu462UtCRN6A4bBiBRL
4aABpokrf5kaTc1JRzHaOtuz5QZvcvJQlA5c9INYHFzWtHxXYdtN9rjY7QQcyfq/IFmCfO94Xqf0
jQbKIUqFMxyJuY31s9xF707qtPEbjKGQuexa9UrmfaH3tdFknO5MccH1fJhFwXGFOuJ29Vkw8YJZ
8M4k2cCyJmxLowQixiDWxVK7OaM7Oehaaw9SmwaCMfNnQo6RV7Ev4tcKZ/EHE2WfFf+9fp6Co03J
kQHvcmzzUl0jaTfSxo40rLQy2XZ5pDpeQQRqp/pr9UzSEOtZX00azLBkT/8QdcsF4Bi6EynIO/zT
MjkoCeVv5jIJEofPyv5TeF0WEzTE4D6ZaEo7xzHOk79tHMMxOvSnHXBGO7rXqXCs2g6SqkNWuLRs
2Acapzm4JTJvc4NdrG07QXbES3oajrWCsRFU99DNCFTiJryRknLthHFTAJJectYDTEEKBh8k8xyP
/vWfrQFDsg7uweLiU2qxdaGk1MyxOC+HrMpWGAbPhG3spSGEhbsA9tGQmh8ySrzqGz6AbD9K0vKm
IJrHXYj2soI9PUhdtL/eiosu5f6EZnDttZDAJVdzB7Vt+GJ7UzvXN9eLtPFE33qwy3ndyWYGTxf8
gXBEsDMp/TVBi2e29DrMbpIKaQIvlWIa3gKQYRuUo9Ty5N+f2t/S5VHIUxytoj2hGW/+I7RDjH8r
o4NwpXqz8ZFuEH7D/jbm+vxSqE8R6bQkuLMja33JzK8mBTndeI16o5/eXNIYmtrHDif+f4FE48SH
tBfhWMipNUvIvswg5/gnHfa5jyfw/VAeN5LlZOKHQlBivsO3DWap5xwsPXBBq1nAVRHnAVJJEqH0
he8fk7rZ9d+v7OdA3Y0WK1HUquS+yl59ElOCzdjHIF/pQY5YpQgi8smdr1Xryfd3CYgRNW/r2j+l
7HG+gjQRFlleLPNVrbryMh7AgyaRoWx0iZKf7X7h47eoY8+zdUprjAmEu+Pprq+b81FA8aEs6PWi
Rh8uM1U+YINFx7mS4XxhK1x1jUDu+3CtQW2KIgnONFarAvzqvNG16FZytrwOYsf+MMDGTT4X/9Gw
Pp6XilXgh105+ywCRNfppi3VcGt67M9olOvZ/WiCLxitmfKl5zNmbN3iccBXq3T4TbBpoubBFK6F
ZCqy3xPxvnBAL6Kq8W6AdR+4dYK3uw+Uj58d29gVbijByRvkzb3+12zf/ceRU67iodes9hOo+ml8
gTS9AxiKikMolijUG8TjUZp3C6Lh3fuYibPVS8dvOkfp9rZtvpj4r4i6kaFQR6VDF4G6QZsM5Mh7
RZEnU9Xd7gpcfpf3R7gDpf8g92Nqhu5N6/xETnmClBhMeQsygmtTZogG+cZBtD5fi3SOKkmo6w+R
4NUSisjj01QkjCWyoLuRnoIP4A2Eif8AaSUfMO+ILCPZ2sRWZJwWbUtZ/twR/ojI09ci3htPPIJc
adp/mlL201H+aUaSjBOHSLde4cYd43hx05mEkmGSg25JKV+DyrDJjRdTxjBaM3ZQZNfQom21g9iL
+aaPk844Bk7ffWMuqtXZxEjKk+jsqxQnkLsH8cuqYqpcv8jedpZooe2Ybd3pusouz5Rrlz+Tf309
RoDvCd/C1E+OQHJl1pbPI0AHgn7KazpKSgmBvG/cPlOTytOGmIvFj3Bgrs22oRRWqQS8/Lp7Q75s
l2uBOvEjMn7XetQoBHGRaAmT0ZpQUUuhykwFzpliUZ5uqramBECK1w31VESnTG0NvypmgnyQmJ4v
Qf1a1G9x5FTthxS3rJ6XQ4pTx+HNc0ZsqE0fp8T8KVW1JAKUkuQnWaxOzABH9YnpITBWmhYb78cr
XkwX6ZvzrPsjzMoiWYSzKuDdkNIA16XTVz7wb9aB1KokH0f27MBjBvgfPx+9Fd3UD+CJUXGgLsed
g2HE+KucMwkTRGLoT5NHtvT2WgL9Iwc3aVsMR3vEe4AuLScZLgebk6dr5B+nsjkexJ+yGRA44WUF
LZTo4KzpUoOIxJvgsqTpTVG3KUkOpHeOU7IxPkaS+pfJTlsU0r2HPgJt2g1jyo4lp4W6msCZUhOt
pTRD9Z6rL0tLoIbmEKnBjH/rMUknDl/g1BRkXsn2a8M54mraT2M8tQYL3MXiCsSQR4cCeni/xe1/
NIeVfcpIaiqZ19vXrBFXduMEaSOdiXQpNYEVm2qDlt4XNy8gWxtVU+voJlvdV0g2MdGd3hWqEmvR
IescHAtoSb/5LSD6hi9NuXP6kE3ue+P9dgt6LSeQTkpzbOb66SbULBuSsggM4QsR98QxYbRosH7n
a8E7piq0Rz81x/ZU5nS/5yaXxbpZLMeNlG6oyARF4d+psaiPFZmL/P3l6xY5+htIrrZWHOgX470K
JLSsy6toL8PBXKm8xQSvol+86LrZhPPypVUfm0tex01GkPCcbGefR3nY2FXqt2QyegWiImQ4rD0r
0GDxTdnT6tirP4tqrzjR6A6ehHUwQCWtIjAybhrfvbwwn1OWa+WfqajLoY5jgZctkkHbKXEPdZCu
e19oo6G9xcNcqsAnAcCL3XNetQjDnABoLXIQJhUeuLiMVXxNIW+ulTHYChggCLDFiw6As2zxvCWw
j4YeSNe4+2QmBJGwnnf+Y3iqSQ4zllUZnYFHkaPfLKRIKObODLwZmBg1qCmwM8dajwKZwipY75+Q
q82ICdzwjgY+dNo+lVOzjsVPcf311uKuNk4woycx0G0IFnXyjm2fDda87Fjw1GAO/uQ/qdFab0xb
Kc/AQNlQ+/LBkSkx2GCGpuCjgQwTDrKO0x+7ZneMFIchHHi9mdZdB2TL0mY5jW/OTV8mU87k/QOM
f81fkEJ+38UaNKLUydhCFpunGGC0vznnM3mswC7GO+x78lAsZLpKAu+exvgiD9SOqlG7/gABhuF+
4EwnecZDDWiKb6kuiICuDsNBcURSDdGljhyU/eXsOZVyQ53NG5lyUkMLu7sPovkbYB+Gm2KzWv2r
0L7MUoJA5LVLlgDFIuMUv3JnvItobI8L64lJrCgYSPCepmU5pNuD/qY85KrxyTD81u16qsEh9W3X
954kZ7iJ0SRgW1yON/ib5QGTueV/WQEsSccqIMxNLbvpUhgiz19oIvll9tOGwul3OlqrRMFVLrJB
n8GAQlIZyJNw71hKz0ZzgY4t61iTa1ocQhm9jO2gzE5A6eoZEfn316WNzpfPmJdC7JUtLCN6M9P0
TBzFtnVWjzYfOL/m01QiwA1mZo7QD6awmOQN3w455DwbKIuF1vxrTRMrBF6faEgO5wdF/hdIL7wh
Dxy0MdSRuGmkr/kyr0mLhcdXFwn67WlfGsJ9Tu8KgGleUSfMsVabN7la7RJrmPlzvnK3e07teVeP
QwEyF+u11IhKClhYY1Q+THXFhs0AZfIQp+Z5q0bk5075JDdxma9Gk6Ost3MajVhb2GPJhsHbZ9NO
v+0OY7lQMu/jeAzexpLzRRJE5p/vQp86e64vaIw5ngl1Dx3k47jO7uee0A19whNZLFEcii5JVLas
uqofkaCCF5CmQJ7CTZLAnCR6+vJ8v7mK7vsloZ8gDw2KBpkZTTgJCRjOcFBj8xE7S0olLf6IRdhD
FyaKW2VIemK8Qzj7tkooD3N33+w1FSx3MF/bJuSa0RiuqMNgaBExrgtQlq6oWCGNiO8DCr84HnI7
Dh0Fx81tiQFlb853vt1BK+e686OWtQc2DnFJNWHHJpJwgaskN+SCB2BJfx9RiTQP/VsnCZf8w4FH
2GeubhZP9Vr45/6K2JC4IiiKyUajMFQyH3nUm6E9wp2RoQ+a/9OP4+Qs/7L7fG2W5IX9XJE33loP
HKv2vqijbL0Yb4/UqVnpvOyTPQGRVkkbQLhhll/zIV/YLuBxmsuU9UbR7D4oMO1WoFIfVtHb2KHX
IAnG7fsjn1VhIcVKyX1ajwabyUQxm1hGkmrVsEplu5qspIDar1zvzcMzvD4jyqWDZFNT6ccShVMa
GZW1O1OsYplwEv7qLKgAGLZnh4k5cQqSd6zY64g7iXzpTbvvkqmZ8e/tm1gHtmx9WXs03zYd4CsG
YHPyl4rw0Rz+lvwbOoGKev7bn9507390RI1eBM+Rd5eCHkXLE6K76E8kmmIWQn70f2eHEUnkK6h8
w2K50zCF528cGC5k6B1I+D6vdrzpz5Yzt/n2n/zSQ+5sBtywQ4NaohsQtBseuFDooijsGL2A6z6t
jLoy5kjATus9ZP920Obdt5xXNsX8oysYWWWoBfIIgsuI/mCKDZUxagRLj70t/ZgrRIxkGIoeW7UK
TxVa1BtQekCVvtcFL1HafoZmRXUSPck2yajD84BW85WhQDUt/43G20KpliqAWKBdbb/wm/MAv+T5
XQLXRumtisrCRX0tCx7/ZxrncJvqzFXcg0elWjR0cBklrGqvgH7ZbAIBBauXBa+d/0klmIinumqm
5xxRX7QOTCdthiLlY0cdczwCveFUFZqrcI2ukdAPjnvAZr/KQ58Jd/b6Va23bRP3P0pv1XvtSeqm
MbUEnloawykK4WwrJHGiYkoJldvo2HWE0EDkwIR9oJTUFI6HCx2m0i99xfh9J/yKQyNQiE/JJZQP
feiNYNJcNxuqlzX4m39Hhi2nnNw0m9wSKmOSk9q/HxJ5UyNGDNa1Gb+NYkdfmoBiPAuvScLdJEP8
ugEw90znwB16aPI7JDEj8IG74FntAy2ONX2SXLzRZp9L0uFVnbfPXoBs2bSlBNuiu6ZSAW6LpOxF
lL/V2kTSwDPJJ2RHw19eYSQzsr+OAMngvAE839oLaIonEsEBow76swGJFK2W0uE7aRinCdtov4PC
4N55GtkF0HZRTOdErYzcCZF6axQXLmfxWOyjP1pQcdWuX/UL+/bYg5n3aLOWmFbzB/UJS3C7swEM
ux2p8sxPsqgKUhuIsZsert8VyZIsP8sUVIHUHyeTvtCJgl4kzZGA/3or/ZGyYUDv6dVynBauW+rz
RxGNMYruw1HlFzl6+vl/Q8ce1+teOsPdbgP1n9drKUw6oo7dAtuI5b4pO97lEGuxDnDR2gj/XJLA
F5qnbCsgNs1WQZ16mg9x4RY5uODOUa0bivjfpo+mkUWUFikdmdvtDx3ugZ/niHjzybWsBb6DKfsQ
puPwz+MwTDFANAtbsHbkMFYaOwUR7+GLAtzsrSyac5ehS3Np8H6XnEqa4QkqpqX3v1QIBJmRo32f
BYFDsZScAHIBoSxOT1ByTr0k1iTkMVw224iB/CpRfV4aeMHSD9wIMC2xAT0GeNcrgf3QiKGT4sST
beJNv4y2n5BMT6sDvVHvkENETum8jCGa7Z5Aj+AcvZ+EYmXezSuByysRGEuzxmbNKvQWWhVk7P9f
qoy0e/KmyluZ3Y9c/G52yUD74Pk1Hj43C7L41qjJ3m/1n5vxOVedULofSsZlEXT/dvcgyzCvCbxf
TPhXj6QGM506wXpLY3P7AHkfAu6j+rVCf80X4DfRkVJZnViP5srlvayi5PaHXtgQHnwSQRS2qzW/
Pk09ZIyVkLqDX4rO/RExvJuSZtgu72MoLCCoDqSpTNoPPVC6RrRS6MIG9S11S5KD6bth0w/0vFUu
EAiX1EiLOJ6FDAXNm6e3aZd9BC0BVrBZLkYZG28VtsWP6NkQ66LqQfiDDyrPyFG2fjdiPsGHcCFB
7urqKCWwY5zz53zmtwHWFUF7eIouZaIClRhHl1iV+WW5ukKiYzneffgINydhNlS93DijjWFgdI6+
hBLBtTVOkh0ztLMzsg/tBZk1Jtt4yeyyoBcMO95R6PsSg3a/7QWvSKIb+oBSH+bSbiXz0nC8rh62
5HGw3CTxg+92eqxYFkmco38c1gfNJbSYRiVf2BJRZFPhtgXzmmEWJxQl2Yi2jw+3KWy2nE8oaKPW
KyL+lsJk3QEDqwxJEfn8hcv2vB5FuelBu7/4zICAcBTKGDLB1Vu+l1BRIhrPSAOHnevDcjriOlsn
jv83SyP6hS7Ucp8V+AuCClwAInLPrakyBx4Iomfx+fTvuQuayp5G919vsQ3zcPHavvTDw5+n27J/
CoDdqB1AnFWoE2o1LiMnL25tAiLfFlEMZk8FtFZiUuWXvIlo8N2bhF7szw+mlATd9VhnPn7oQikK
tiWVnDo+Gbr58tIHsfq9AReKFec7B4zc0E3ME8/VGvSw7bnN9NthikgRSoE6wKALVxokKKtHCHOq
IuOOl19ZFaOz9TLYjhH7UMXo0FLnsPHvAn4HPpSDrBQQKRDpHSxAFI+gaQRUoyVXYGj7wJiNHRdE
Yj7eW30hxnaxK8m0YMsOWZ0zxN/F9NdJcN9SbOOuvtWEawH84DEYP70yH1wsSG0XfdvGGhiqs/Te
ZTRA6ZR+xONwR6nv0SgQyRTtK4SQ10dtiS4Cmd3q2GMja2EvlR/8G5lDS+Pm0HGV8kk+Xd0BmMJP
wDwPdRrIgcw+c3zy+mvIOm+ojiAVbdJNcas5sfNL72T3wcrmewF+JSUe+lt4YfuWonTOUl+KPQzd
8QroPQmVOU+zBZRi0JUvRTU4DqeeMFhufPZflngyRn5ebe/d/n4ngnTelbdAKHYsG5lNQBlrMFNc
KwM1ZWBOUDDYKP4uh3Srb1BN9bB40FZgCRrhNIFBxgAk4QeAp7/JuU9pRIcR9A151vHJuZXk/gl7
fSSjQvOQuUfaTZpolC1naqUOuI2AN0ginpFy/SN5ZHWeYwiGA9BobTc/lIKOhdB+yExFrey9jTaR
nzdkWrP5sGalCcItYyNF5c7mvWP8vyTeEeTo7xBerqixX5lJEl9O8h0F+f1Jac3QFeMMlRc4DNYi
344iVxK8ONSsqo1Rlvi4iF4NWnH8HVJ+0DG2/f0ZNVtQxs5Ed/u0DVQYk/EqLckThn1RZp9ypL8M
UpAByWM8EHDcAj2yXsWpfk9Zc+o6FedWrZa//3OcyxgL6j1yVzjcx7jmADC6/P5i3C9uQqQbYZqb
ry6GMHWHTWZ2uYsRVM45GbNmDXhie58IgePMyYpi77HLJ7iz2RvI6zpFgqzYp2lmqb6URhzmvDWV
HcafiSuSoJ50MbvVyTlsJNWGU/jEbLww89P3U0oTjEUhGBHLjv5yxe13USM+BQbCgUVoSFOu33GY
9l7mEkXvAJ8bEN3TaZ9zHx0eiayAh9RuJuY8d8UimbXgphBRdAP4Zqlo4xE9wsPRV4G2dXEgcKnW
/DlEQx13nZ4KIZWPKZP2E3n7nt4wrYM5yJVzVDS/yBDQYDoXckq0t7cEDGBKnSX/Imybcwh/pnAs
63tCJyNL5eL47DbYrYvEV+HwHDqEp4WSqurcReUCS/JcMtsbZQxdBZGpqbuUt2istALLzZ9S0rzw
aiiSAoVzDob2bmguTR2IL3f5Np9WAonvQdTcobY/SUMhw26G45xuXZcmalIXtcLUkfO0S4h1di2+
SYaiMxKbs04XG8nV9q2zrSQp8XqK9YGR78a3sca3PP6TWaSrdsytB3O1XcihnfKjXEjES43OpcjY
axbLQ2L5ahurIyvebd9yUF95kpS50MSntSIHncsau5fptEaJFzz4fY/QXW+7+6J1dTUSD/QaeNcS
RYJl4Lk3BTFQx1gB3txD13S1juoEZa0nuwxu/QVhNa3VnX+eqpinsREuKbRVqSC+DkJ8Rz79QkHE
u4E6RsShQ43Dxa1rE6PN79biN/wQsgrwA+FQqwwzNTRN0VEkw/edlbKSWHVa7CdEFSB7ZrcQziaQ
zPv6SMINzOhprvQhMuTjhNI6BXcm50WJM+lyqIvrsu4+04h1lOrxXvmjdtXSJve48zkwzfHNea9N
8Kc9iIPHRlc/Nz4yyESawg36RE+gfWY8ms89OsoFad4TNDtf/tFPoqQlXEr23e+dNUwq0tDvNhTl
WPYIVmEC2gNxsP+iRMQoHShOVNa2h8sGQmhe6SLCAaxDqJ5DuTnlZqSiD+z5QuSJp60ETrMc8seI
Ftm0LtCpX8pyyFrobn+zT3CUchUUrZ/XQaSq8Z5s/r/UYwoID/v3gXhmiEGcjUVnhrTs+vhhTaAD
myFb/PhVywIVac4wGa3/q4s0je3SyQCvcgyCb/Oz6IpoNjMpHFd8WDK1QnIpcErTQSdgzXDQ87jm
zfXq7zVPuRsgRZlkFL+8ZvEeGAsd7l8CHRQk3Y+bV6mmi5rqal4pNB74XhRQ462OtIaQgLL5E3py
9WS6ZXS778UzUwzq6+3wQfrttihHEKIKK41ajLTv88TKnvZQNwvlALY8HKD4tfBOcoqC35mTI6QA
lfAP6hzjld5yaeO0VO+MQK7lvNlyTx87V+h+9nbsxP135PGOFhLdkHvaRFAZjITkyUDKV1dJz9eU
Y7zE5MH+XGPrakBClxHN3M5sFpmqOcN6++ye0nZfGTSNGdIZ5IytPA9RGwxg1GeQnNOawIFBjVuM
NvR14K1UPrcBjh4bwe6hknbFUbRO6pQ7+CQQaRjHsIAeAYTUnW4aoJc+rjjZiVIWIdk/7tN6jZQN
ujZ33TMTa7dbzmDw5jg47zCuLJIk/Q2LUXxoGrbWOvGDUeDP82BB4Knn7lWSQHtiwuRvySbKgjhg
GobE+nt4QSUtMwQIxSrxKQEEmcnTS3se/70GChYTstxAsSy1thNNBtD0JCXcNWE1di/XPdSYZkAI
482pqLq0vn/Im4YMeVzpUDZMYTh/gj8HBZi3d4tdLKYoY9rTzFyLMS4sk1zTaeG8AyznlM3fR7r7
CL2yb4G31LuVzC4QMpmibCwDs4NWai4d9vkdKMGyXE/Wo493bTQ6A1MGSyPL0s2kbZMfpg44rYs7
HCS0F0UCmH97RvF6nV+UYSsMBnGyPHkxtY5Bph3ZoWzgiTye+J7Dxkd8jwzcb/M3gSddRZy7muiP
++EN5mi18rVUGqso3XpfvQ7PqmBoYU1gKa040wikwDNfkMXs47lrwjVGienuF8+rBI6JMYFcdQjS
buUAjbVHd0YF1gE4qYDH5h7CVjCw/EEZzMtMSOsBQIZArwckn5Wfd+nomb5dZMMpWvu9u2Q8kZhS
Kyw1FoMyxEzA5mHPjRHPi+M495LnejNwQXpcUy6OiFfksCF19K89ALPY7NPv9moAW0BgJhux+ABf
B4c4xWvyBZgO/yiP0NY3nPZtX2iHtyyWLvRJI9yBDH7ZgSH+/f0RptiJ5HMgf9xH0rkNaYLhB0AJ
NWB+Qyk0tibNB2UaO0hevq6190Veh3T654sn9HpiQX8D2t17x2cSaFRDXj6AyaZhc5z2PNWrEBO0
KlUWpeiPzTG7Nlivj7gsCw/4Nq3y+yixto4CQacFGog7uu+WuDuNyBRZheTKuaDqkU9NesHzrzPi
7kuIX6H9S4UsFObL4X6o9AUtRLHAtbISid61blklDkQvB7gqmRcciUtd+kSgYXG8Eeb+lkf1o2i1
ZWmpMP4OjSmYIbxWldzbCkMYm+fVVDD9vqn5ID3t53Yuf1TVzpX4CbFehqhPyLiGTXy3palEuj/i
WI+uqfTwm++mw4h3xTMMG5B16NlieDDMgfdYwYXrKzHiOhnvetAG7uoofJJRMYbVWmw0o0UU/eUW
ZG5QCslC/6DIzaHxsdj+KROZnb14V7x7s1SrJ7+u41Sz6skxeckBvK+ADQF7kjrlldpurG5nJViB
Nk1pa18P9imAcCsRdp5oBliNVeLfh6HaIzO2blVmAhyQP/2lTD1dni2o+NepBToLpY0yH6gN1m+1
wS2a1+uOwAaAO8ye+XwuTBmTMe+3rMIyDBdVY2gcux1ifSa+wZ5xHlZxXReEwQgcJM3vEwXiW3tm
r32ckVlsmABnc93GR5h1wLWr4v8H0Lil7Ub+OHaMx8xHqesJvmJYHIR5TUbeRflQk91eG3OHnDRK
2AuHijzhYxE25hi1xeC0fZSGVsP11IFfw2RweiAv1RjjSx6DKl0vRsGPXaseLMsFdGffaRaNFlN6
SO6Ptdti5ygeJPk7eD9si8hJAC3YHH/2uk0um1sfD0tHMsAtazyZ15fyZCNBzmhwejuP2m7R5yME
+FueHluXOUKCG5AH2ZkWZHDRzI6uoHnXg0gFh9ysQ8XeXQvu3tcMSZn/DuB4G0mOE/0Bx96MP085
NVNTNNn6cqMncQ0DtyxUOCgQuorNpjMRrjgRCl4aPd+/w0Ee/Nx/PHKMyow1aEDG10dnuEUmQyjF
PQo4GxmQ/EbpfdpWJULLi9TpDDfy93zZLjWoXG2Y/cvQ8ftyPeqMzjsBHvMMUCEMZlkgbVNCWMjF
IyfCKzpu5o0UWyxb/yp/0+WWhPT3Aax0HLLy0Y/HeuBZ/h1t/DKozzkD9RXOkFQABzzZ4Dco0bJ4
194XLdgtIkoErFc8eu6ha5M8sZg3aY+44b6FoAw08jiF8gyeOVScsFzkGY9In2L+mvCHk//bzTrW
y3cOR5Bi5NMIqkwRh5bKzTlw1QoYdAyIAOxBgla88uGnB3AwnEszGUfz3oysvkjW3K88F1gsHiGq
vgfeVLc+tlWGTryhXzttaCPmmWjx+uqYbcFQoDHlCkWZ98b3JLn4OyXPxxFaFHbawjKe854f6ksX
xN/CdlwL1r2wzUS9rnIEctAB8rlZALoBi1NzxH90CaNqG+YD5cxKMlRLsQtl9kpBqHC+E+GudvQ3
mo/hMxZ+JMRDUllx26gpPQo0f8J6XgyZdfP23Xl+P0AcC1ZnI591lmHifVxzPAJSnMGzEzNW5mN4
TK6Dll5NOALj1GJbSqFcaIQc1SioOed5i+5U85w+LSPIM3CnKiY70/mbRxb28A8IAM+lfl3jS3xJ
9Os7qHniqH1yuoZgWBfC+2GZ/WbTY5DTs/G23mSXzS88swRp3by6q6bCIPP8GAy10dtPI+G0Z87Z
aCAng2vpgihQ+XBz1HMTW1dRshd19LGlNP117tKhymeiSdcnbDUaMgqkm53OJRZf0pw30U4i+eH9
O/A+E9LEprqF+NNKPZGh4WDM2LDyggKQL3pmkjASEI6zfrBQwIuxfsxjXJzkcSscc3IIBNDM/SNX
5wPU3w9Mrrz/O7dAQbAfzB8AsQMPtSA/NK4iLj/ljKw3VWvkZiQYPiF+hN6tHHyOXOdjW0XMvytg
uLoFnPxugTO6YswBeTQ8pz9/24JYti82nzOP1KDApX9/79GeiGiO07F6v7caMk9Jj22w8uD5m9Fu
Kyl4zviSAJ4OGn2JUrXTTZ4DmF28bBaPIANtujrhhvMuDOq20/kOQnYb3gGTvwcVhVg/bs17KbqM
o0//SqoxcnJlmMGTVyY9O0r10gKDbIeIuPxeZccxmQwaPcYBisTwd4BqGugK88VCSaszbVGK1FtB
/lBNF+k5JEc1HjG6N2tvo6oe/52oFOIsBMxZggd3hCGBwdLVj9S5dzdjPIhLEsq4LXFfa8fP+dLO
Sldlb+6Dj7hOjRBU2el20M4mXlga0Dh+Yxz1cPeLGKGHmtQXhcgpDnLxRd4kzOc45Har/Uk55UAe
YQ/SuMT0G+yELytyjV6jbSISUXvMWW4/SzXzf+lwV1XUSFuDtUSFggwHk+1pQdyFDLBude+8vUvY
X9n50kACm5pDKIcrH6d7xKxklNxayBAcd4eEqS+qQKRYp4k0o6nzqRZyJPKcUB+YkmmvsNvc6HCR
1bNBmTeV1jFgURcTn3yYLknbOrdrMBzcK1H0rFigOCFUVc/t1kpxSfu2xPbikINrc+LN6q4CbaRF
e1M3EEcpknbeSpA2UVoFfJncVAL3uxiv/LZk5FpCEr/odRd4Uza7wF54QQkbOhKY68cpx1WzTMMU
u+Qty0sJ+UvOn+kGzxS4VRL11xcjOi+FwW+u/J68RDsdzqjJ88BtVL21A9h9v8Gd2nPW9lQrMztv
PxJWaKW5aB5pXSd+6tVqlS/tkNFyVlC61I+uZdFF2+uyHmfdn02pmniqQ6y5abcSmE3rgi+YYByZ
5U89oGb/Do9gENtoUANo0FhOMRITNEG6gNAmVGKEWDT9OFNFGzA60p4dmr1uujAbj+Ug4ckcUHts
nO7c6Bn3DIQb4A1p10DwGXA3MbBohkQa8lXxDeySuD/yYKridWh9dgOGMc7RXLai5f3giUl7VikM
3fziUvz3w/bc63KiopVSpv5BQyLUNsgk4L+NUi7rA1B82H4ZerijQO9UtGweNvra5TBt4TzaLgVK
TjCKgxllulpOKAk0/9myhL0/CWuK/8lD1M/8r6wQlbN650wDAFxGgl1RVafmlBxHkXDsdi6uJI7t
VvSY8kyjk2wTYxbZaPM7HunI8tFOnNVozxLNM5MlacogRSybIv4JSVm//PuNEBM2WHftQ0oO6n5w
tcOGvrpNIyEFOLLPrJexeVTH+ysw21A+hx/hRWYutSDD85Gh9NHRWIwNhOeWhdkWCeOPfpfHIpDy
gM4vO5gv+UXGUUbQVLxL3ROxK9rnUIz9S8IKemJK94bGS9in4Tg9C7kfLIL5OSIPeqWyEC2jmBXG
fyW2xKKAIMS9mQSrFEJLw3owT1Dg0Muss45RHlap7vfg+OhA0WbakL6G90w7fhpQjyTzGeS3BzaO
jeDArSZVWC26GyqsuO7P/j9RsCIQa58TnlbVzF7BfFPsVNLXO22rhA5nl4hBOYfGei4aLwIzNntJ
xh/Fci2NBMgGPPCZ2sO4OURsQcyHiod16l+Or1584q907Z12EFdNTnUCq/AtUnGxPMmABu1iwVNY
MfO3KFHzrP9JqaA18+IzB2o4stGvRYDfQzT8S7Ux4pDsZs61oR50HGNBpPMFX7Cxfo9eBLcvHIcj
Thezmq4jAn1mgbFXUOcEZ0/WL8IUTXcCC+DGScyrc0AZbVQY63pB9VhuTVk5YFIB/byTZHhUmv3m
cXl/mB994qQmuyCLHNPZ2qkL87WorXGdpTW28NBJWgw4FgyU4YH5HDm+YwYNm+KRwoG4ei4pe779
a9aG14ui+c9EVzuyCD0kP4sguHK29pSctvTDlroovCzD9UI6Kz7um4xL6UtZvWEyy1pGIaeUy5pY
NSIY76+RS1/2bE+bAFkLgwfdcI+GBCGVp08njj8BiJSyOqw68s7W48zulmQHTpQFGe9sXXz/zQfF
ZAr6jas+CcpiZXqXa0jgZFoq+nAW/4OSZbCMpmi7G9eh4Bxzm6PUoZqhAU8W1JoReI8RKKRIwlWu
zzRrQfOl4YwMh3b2TZEf6dcYeWrdRaso66F4w18JTrC85U13hcaJ7zGuvnaNUkIpEgr5n+krKimH
OvZ6LR9M1bIRE3qmxt5nhwRnrXe3fI5zOcP+9TAS1pGdyBXXgHpBFMaO1yFL6j/xrOEyvPKDc+oD
lFLb/ht6KDY37GBUCx7eAZHbjRxsuC5i5G19Wp7YkOXk3YqeSgpVIuUCAcojgZqgIWNzjRTyBdFY
nEvp7dD1BgqTPfjngfpuABrMa+CzInEe3Kj9nU09Qbs5NMoaJ0lVKcY8VvBK1udTnFxGaW/WA+oD
U5y+NjwDrVH++KihgUNuZ8tQ/MA4XwXjwS+RsOVAC9PqaFLqSDbS3zmziT5ixdvTzMWNy+BbcYkX
zDTrWY+yRT5zo6LObpC7J5cXMthm0kR8Pva4AG9h2IMRnHj0Pg1Z6yb25qY58r6ph/Z6qZcD1vDr
UFnEbWNBpbaet0/gdnPsJyMuPJnXY667MBLblbzNmA0njkR8uf5xCsuwPpS/nVqNl785s1RlbJCQ
3n6feW6pOPWHinYEziklWtNeP2EupId6dviR1jSmaL4kcGmi9fLbcbsyVQ25mPVMGFQONgGLawrv
CngriZZcJRdJoGx3vmrIZi4JvDJ2Z+q6jLfVo1ulbprXUM5yH4KsXxeTAxq5clOqVFhUj5B4ouPZ
2egnRQN8GewEnRF92ZfDNsKTkjh+E3banw1XlRHqefZTOy4z1U+X47OD730oBPk/h9eokuaxy4Oe
cT0RkszCdNfR04GFsNLiqFhc00mkBxP/aZ2kdFlWlCriFikPKFSYR+xy6Pbjhbmwo9WWxxIWNg71
Sy7UocJ6gMMk5x/DaQqIrYS69SfombN0BGK+30YMfUmGT+a8Y6jAXWzbMEZYQ0OBb221P/x+CLGn
W0f8/9BqZGyjbQgAREadVDqEAG35s+u7LSSyVLq1UMLREilhuH4bwqc4i9LBnfZO4aTr7brdOvly
kxPKxgkIFhqFIK2fC/jG6V6GV4ROe8wjiGqGSF1ZUcvaz61PEl3rkjBeQ7Ikm307tzLxLk8N03ac
i5fSrgp0uZciwhykdwuCanscs5p9d7yWKI/Cnm1HR1BDt1J1Ep4xQpjae2qGLqg6ypntS3Jtgmj5
FA67qM6eBi8kbb8UpRuAPMomofz8PoXZ7Bk6Q53o7tRymqmidX3giLgDHwIHDCoxq8Wn0CdTEF5d
YycZKN1XwpEIe8XUyojYRKcYHI+KxPvbtBGoUCePzu6R5HABLOzEaTexGYYGjBuoX17ue8+ufOne
6M1hZe025yWl4XESOZCdMcOsAgLcLiFZjgm6e3wEwQe/DBJ/0Arv0GTPH0Lkr/5r6YWcttLJ8bC/
tcy9d/68i/rQHZIU+RdzL+6aDPrMSu0bM0QwrwOgImN4po0fdBRRlvxGGfcR1ARqQLRqfF0Qq0Se
gsYA9pYZRx/4hwzhOmMGd4p4ZcKeZWF2e5nsPNv0W+e+Q3BtFMidnPADEj5s9mtL+KLhmcfFqcTp
LmpFTaauRczensXjFqLmszQ48m4O2QBqIWrzLjSU8FyEAp0kzUe6EPx9UZyZp/QYXZgPbodiYoHW
lmx0ZNgG7wGbtD6XJitKEKJXjNkJSoZnjKvNhWLz+DR5e7bwUOexUdkFaslEeN1GmpyLQA78FcUG
Au8GJCYQ2ZjLA1550VjHq6M+Yeb4XjMpqbfcQ0Q7vLjJuS3Z1ymqI6SAt16XP3wd3rbFOnqD2Z3/
yXvH/d5FhnUvQeED4icK3w6dvzbBA2PMBXEGKxMW07rVHyxenpUUMFhGWnDp/FXBCTb0nNn8v15q
VCdbUkqEA3JKa1ojxRw0wylibKOlB0YRotFwm5T/Bwzu1qxVbeVCBcu3WzoIlijoiIgB4jugcQd4
/pSKqGuKPU3/kTVxq1BZf7jjJWEFOkK6XGLgBEavDerCtbQXbHU+TuRJh16jy7gAC6jf+Nm+pKVf
Oz267BlX8Rsjh6/9ppCQ1caKx1duqcUdxFyDn9v7s31ZzJzdcFxS49w8CDQD1aT3bmM9BDFFTPrT
pnoICXS6vwJBKDZOfGPjPBMsh/4tpCQVzsKjuUppyT4VybAXkAnL8VcbOpHX7oGFvhpcLD/uezOO
5+sLB+hrPjvEvg+EHNvqE7H9U6MMOv0lUbko2cOfuSt3gt+8L0QSeYohCASyjQjWeiFdrR2GHTzu
1mLIp46KFZpN9YYtLsYK8E3wUZI9Lyecaa9i91acvcWa0Ex1Ae+CspRQ9hQdlX18hvmvir5v6JOQ
EmeUJ8z/VxPaR7UNe1HlBa9ZmBwgddwaArRXiOd5DWoVyLniwIRlIVEqYs40mdqJbvWOA5rw3fWh
o20JMwu6QYDyetQVYmgdTM3G0qPqCiOZCsJYipza4ErrBGRx8pI5jTF7rqGqXrx87qO5WV2Gxm1e
8Kn+77J+GMYytAjSyiyOk6zSJPsEkcObuSuUm46coAd3tltspS3WLBuvnVoy7WGlg3V70kD33uTc
hnU04VEf3MCmBTcgI6V1txNMiaED3bhRUeZY19XwIUEWv8aCUEaeDN9DAyemQfK0iT8x58Z/Hr6Q
5HYyJqNENtZZtLRA+3diUEUg6fekK5QKaLM+8N/8UzRduyN9LzvZSbBzegD7VYD3p3d9vB89/vyw
Cxnc4RsC2EEHGRRQotGThwH5cWLp427VzepKwDmtUJxNlFEQra48p2c+gsasshy5w/hNJpCPNj+2
qIWPbnsdos0sE2RsFU/eNOvAzLCS5WOMdu0dA4bqo6G8LIU0/aFVgzvQ1+TtGyNteJjp+bx+aawT
8wEiDNTZdWUvyQsuuoazFyCdPUvD8KAEdTQH22qoT3JeqhzYOqW4KsziVCU7CM58KlcWr9GLIgs0
colgl5kR7xjhTMPTxue/hVONP6GgwxF9aewxYxwlEg99+/a2V5LYkkBTYt7PCIsa+r9tthX/W5kL
6iGvhEVbXS+SCQbhSo+0o9u4mH1mRH3ecX/OKbhCn7cKmXrjW+s3JVIKOcMnmmy7CDp4AZP07bV4
uUriPbTtCog9+DIHjqoIYRPwtbtW4IzbZSB3IfPHAVYSJyBfCFLK5VizT5x2p5ZgzjAENYZ5CYnQ
EF4DS2fVexzdpsa9hC4ePKYS7juLL6Y9wVoySEeqAYoibZ/yRn3uRPTnA7c7/eHc/nB8CqOWU3ug
+aW1AZjJ9crucoBxc00F415K0ii7tGip4ZH9w2iwgxLj9fkSyBA44v/J9UHqOraHcS9LXZLWXUZt
25Gts91l02RbD+cXGm2zgQTu/0OJjZ5Trt317XJxl0dYAv6nuWGnok3ncXy64ZcNvOlaEFPj8a8i
Aj+MQjg7nT/yVaoQ0qUK4p1Cf7t3VeE89uTVA+VAGnTd31SIKfB0KwK3ubL6lHDMLFpt/wjpSR+L
nMTzkVrUVB9EL6FbClIuJpHCNJRAOqOCcI6Q7KNGmaut8/0Owk+n4dgyqhsw+08hoI34aejF+Zrb
veQFaHOkFFOnJaA9+tXzd+Vqa9ATdWFTby2bOdwyUpDiGQ8EeIyOxCiB2DWrbY8DWUVr4GEXIfS4
nZITWyaDZExBn8STHfL3TnLYw9G1Uz9BrtRjofaTnZBD/nPRavYdzyz5Si4JMeuESmPGh5oF9q2A
0noRohMYYqQLIBtmlbDOlYcwrDTTHFU3zMT2g4eI57wQ5t4Ffpig3EdTjWBNJtP9ro+gUpu7O0Qn
05Qc4Wc5PGg0atMv/hwmBrWik7cKIQtjY1qywyZwxChJgBtXEpjepczeAAWV3tI6wzWs5uF0izNk
KnkB+5wG1k+ZNZbuUCVT8fs0ibswUfvdV9kCJ/J2Pi4Yh3lTeQ8NvS6whzDzeg5jLmFCtcQvMAlW
ERIwE9+4wJteIHBifJS6IbZ87Krb5p5P5Bzg3YSyT+0v0ZqHzpy8xWTOFX6kkwEfn+DbRgub+Rk/
ReQgGJ6hvWbiyZGzigBiQZ/kAG/+J3zNQTzqSUyk5ufS8hQGTEciQcVM785oeYREMqw0XwQSdulr
UzsWM5BD3LnmHeeNzxevZZA3VJeDU8Dy8Jwdcx8grZUANjFfsSyM2XqeqkL+WVq4Os4VtzpZLQAR
1A1Zu0M3bJtguRwJWG77fZAQYRDlrSGULqqCHpE8qawJgRFW7SfJU8j2piJZk44v3QWyijPblOgY
Sxfx8f+/ASu1+OpPhsEpToC9JcrjjeHZiNO9/7nGaWXnK6Ft2PqLDx7oPacU/v2fL8/U8lLb08o0
pYmDElMFte2UI0QKgl5k1GzvZNilc+jrufsMP4cIlc0x5hfaDtD3mxU7R23APzVYWW+ihzlgGWug
WinyIphaOT+BgRoDwlyE3EliEQbI3RpJUfoh+8kJM+Rdu53zD5WXa2S83w2iz9EVc7dxTmRtXeEs
QU5ygs+NFQjBgisapMZ6Wknr9mvkSn/7SjE0AIJsP13hKNW49Jm7I9hhIuT/Zx8RVQSy9trpLT08
XDYZaI2PuzzI4JHRCTRrCNE8YgJ/Cl2kOCrWHdMCIQAkbSX1GY+MZFK5dpHK8fyQFDvR2WeWbD+u
iBn2qVVl2DuMazO0ey4zKSSDHhXkZgiLcbd1gDocQfh7jIgCbwRihTCEfk15aMNj5deuP9K8fokl
mcFaK2w1o5IZEkSfZEnuTLmgkQJMKS9IfrLxFz/j21Z4iEXOwhCy6PyL8ZFlh2ENzGThQ1LyG8Qr
CcxTourjDCSZzTSxit8VlB740C6AjTbrx+Gt2d7i8tA5+REABhAtDVqf1k1sXbk6QJ8l5oXN99+b
jEs7++svNst1hVYs0yoSbA+pVfLgKQahxSbcZ3A8aPkqmU5HGt9Tzwjatko08st8T6jgtHcLXFTp
+J/QFkcuUlJK/KT+dXYSkpF8ixaAUgj6TWbmjytaMQp1es3GA9sgas/wpZXPIvHV2Z5wGOWmh+xn
8nFq3Xb8nPcWk5fGSk0Lh9xNhp97kkQwxq3Nz+8oy/K7JO69mdSx42pTWp+H37vuatGt9rB/8HIU
pBcjX4fFoWUfr506oBqa6pxfSFBk4Fk+miPyOXoaZJIsOQoCWffNlrLVb4VUB6QajfvBqN9ClG0S
PYmYWjkz+rEjJL1951Mz8DqQ9zpWhYxY3RQliG5f4Mv9pCzs9QPwii0kdEAJ5I3LklyQ8K4xPkMl
pHGmu5Jny9/8I7ZflN5Y1J/2S6Mq8BUtkiRpIHMQvOZa2vCJCETLdLT2iON/NcWO55ARX5Bsr6fF
iBsmTa7ZTGBiQqYK7xM2/cre3LFeb4uLBN8XAUwjSRU7XfVCMQkUY5oYdFITT7Zyqf9bD104ku/g
8fWt9HTNL/PYcSXnbpo/6j+WEZgyr31TIwVqJvQ+tfpYu+i9kE1BRqao/ST4kbjO5PhvpLIhpj82
BuiaeR71zu5veLDaGbQ+6I6028UL1C/LTuWlWihiXW/enEvOYzkLGYpoUvL3TB7g6qtipUjmZcK1
HQl6boZtrq/tPbjd4G31ascnFVYOhQjumRPvnXu3xC8bscKi2MFpsI00QydZRtNNxylR29UYongU
FGBro+uNx8ohZez3gVNaHJlSL6YbjzhAN+JPyZr17hWTv80J8cek6cYAoIkOt4VNdKPnBEa4/TOL
IMsA4udv3H3atYTBbbjrL30Uezzky6P7VLfw7nP8c2RWG+78momFcetrbu4br3Wuyokpx48mAll7
1QcMzHOIiyFwFkUHkX+OcxJY9RyfuUjgW15dWmGYtQRLeUaR0Rj5PQ+2IynfdPAUYvkbtZ77YxI2
74DPTkwddsD+JrC5L52rFgng/a7yd/ZiTzL+twTC0FkP2LlyykUlG+3nPZZhosh8d0fQcoBTIgq5
+frJxxgPINGgbIw5oDpRhi/HmlKL3HS+GjfsBqpr7TjOyYc2MonJSZO8kycaZf4baYTSEn4HSt5B
8lB71Hknti2iyrZYEK85DdhZfpoMkJq1qvbtm1IQZQTDghiWB9tIGtBeOYRP/Wc3nuiQH/pjaFGv
Iwe4j6+aVGAarTRyxW7/xEj6MuLkLWYBFUVwue/R4RkTnv9s/TIwX5AoJaH0hlmqCT/FOFwVaoSS
cPf6/+DqfMMh6XTd7HZOlGoaWOevQk6zbvdhVBRXJoaRORUd+QMWck5M+6riulxjmCqrqN5r37ML
FXzkj26ajkcB+Qpyo7AImKHrF8gbbvfwshrr+ffQ1A61Lfkkfat0XheS/l2Hbr4De+0j6jRSXIw0
/5mCBFyaYFG8N3QEI8PFrxgWmRYAJ6xvAElbi5DDNDquA5xN6nFYAYKNh0oFpgVb9siowTqPtPeD
12a9hmU/5PjHLSbcQ3D4NFMtHSxrSEP97B+4O0qwCEq0SgULd+undyDakPVZ/cgcxfVS/KcKXaa8
590oOu13TGT7azIJ2/Vk8fqQuUxR4acCIUDKNEiwXKbePh1yfpzYzu5VOqOohG/XmXMAazBCGy3T
WofwW3NSSMLuO61V2I4zrzxwubBLF0+hERKBustj4KO1Q5blTlnty/pq7HnLS/nOEC+YgAt7Q+dh
xXQWMJSDIN+exsazKBn16DYpWG0R0cThi7xo6F0a1m+koXvq4pscc1CqCFBgUUyMT4ac4SEDCJ5T
po21pO3NjrpvkQVvGqfSPKWTE32Vb84X6XXAL8Y2YU5t9yTobwbl2B/0IAp01XXrqiyYCmS4Ww1K
yG73u8J7l0FqVMr+wPTl9Paq/kTHi2y3hShCiqg/7iJD3hvtPcW+aUKhihPuw1PwF86QiCTm1BFZ
puiSTXouivQO9btx2H0bmqNWiYlUprJByE7uMlE/dNQIL0s2r8waHdGm8wlqNpcci+/NFTbQI274
qp+aq+ejFRMw0IacLot6zRfsOEQ9UD3HPqQxKCh3ZFYr8eCfm8lGoLPZeaXC7T1JUvClF8uOhFk+
DccHCYQmZb7urFv/n1GB3joYuemX8ObpqUYASyvp6bbLTolk+BVIztRBM61UUCo/dzadXfV+bMAK
CwTl5PIqnkeHJf1iUHHDtiIcznjxXkqvXXZ7eiJjIpZxCl1ecdB5EXragURXOuF75+jdhavfAGMH
7oKxo37jwORCuu2ctgef7h6I8GQVqhDhCinrB+9qx0Et6YQhchJh90jNyvD/q1YwJtYTLvNxnmav
WdgKgBp4yime1rkHJL8CgqfXzKKy9cKA1BdZjv5xBpdYsOJ68GqiHP3H1UxrKqOP0/4myH73XFrw
vix4Yr8W+G8gDQsaTNmys0489Ez+HNPo99DxztZgae1TK4WCzUODfdpTehQvGiCbGKs3Bc2xWVIk
vVvIqGvvZWVuR/u02eJ24X3qlIaVwExBC20TtfCs4nWcS/eVBPfCQs15c9xSJOANM8CQf52TB9Vp
IfZrJp4mkix+j8TE54Rtuj5AJpBT3TxMLM45FNDgU5CR5hmGB3x2ueaqTH7WaxwQ9+i9BnRLNMzY
9oj0XgEhfq9jlid/SwehlksPGWFSIY3q0fEsI6isNv7Sy3xdB9vbbpgZYRhJDPX5SwBLpupVPRc2
v5PT5W6eOU9SACU/VNR/lw0dvKnuCqE9snvYyRd0I6gZ7vvJe9r4rmUt8OM9xx5CIev31+vupmgc
UIKa4YjYTMoropPAr7nEVBn4GUeUMfwzYz7C5ZcEYxohcSFFJnlGnmavdO1ObCZ6+K9+rawHpz6z
GF/G6Du51in9RF8fNNbStt1E84mLBRK9GvrHD+kGSQDnVfXZU3LgfpYHgumW+VdBsAV03ADutYMk
Befzz4j0xuYHvKWuEksqbRz7sBXmb8JxwFhxj72Enf3QZnLb8XbQeE6p/n/DChIE+arqvt2nQe8T
UofPGFxIVuuSStRUQYxgop20POffV2wmC4yQ+N+o4XyH6m6qeDUCrzvp4woJkVBaBr00hqqzDm7f
iDxLB0DTMH4n7vsaZGWtCKHM0PaXfFCWZFDQzHnYSYJVtHeSs5HxO0/pCx7+FkwUwdcQXgfaGJdU
Ve1X6jLYw/luDZxGoGPh5B3izzgMGP8kOl+GWQqbfJ1/KFgqd20suUQZltwgL5TfNeQQUvGz9IVp
K6URmeoVVQhCkcXIeQUaKrHaOw1uOjn5Wn0jhZ9GAIvhLWru/3/EWDlSjd2gxW19+ivIQQfzXTO8
eLcgVNka5djIx5CMgRAYlQuKXZZJqHkWXc8hze+DrcnVwMCQOojhO7ikwV4uslV1YavFRCB9ZUyk
qnJUUfpxAXHkv7wPcPOsgN68QmS1y5vIcYLbb8bX50aD87WBKZQIYq867IkN+eoPpuwO5suiN4gb
kkgZKP5HVMB++54pQqMJyUACEk6oDdyWb+yYOlmzJeMKB/pfLNRgRISjyG0QX5l5QYlhdJ7Klyrw
XwBOduXLtFbSX1q5+TzTYdGOAWNy33r5YsOj6SX4OoJMPrWvoYgu2LrVM5i7+QF/SCshtabr3o40
Hnu8micGXd//zIso4cGvz1rGcY7hJmQyrrx+ydTuDhHUo/08VebkLycSOqWm3QHdU3/wrO/RuaK2
XuG3mGOcWKPUk4me9XuoDXzJYNd/DE+Z2t42eE2rraDBmpDf27sP+N776YdtwssiO21NXT8j0mz3
jiBY6jImuKXztqmzYhPdBJVyiqxj+2zpapateT/ptqfU4shLY7Tk0YpvMl6LMB9SfIppPlYU6P6k
NEDVTS+cy63S4gaWoxo+E3Lr0quJ7sKNE3ypu3T0whQ7dF3382k5tbF4/FcMu6tF2ZaVct6HDstn
jTiyyGd3KCNbt/hkSv+N/1ZQ18iyMzfS2X61WtaKhPUtSTGBy79VmWJnGayMWcR1XZnm+e4n+JCX
ByiSQRY/mcjI7X8XZlp9B6shfoyogZd5LgbyV7Pjyu+iDQHYm0ZI0L3Efg4g6Q26TxQiPNxL4ae/
4VSrmL4EcN5TE3IL6uG91cGZ57aislcbEraRoxkzSZh2i+OIx8tVzlE1lPqsIBcTH8jGTM1bDJXg
mS22CVzTbrm/nHivZqU9ObsQBwYRaOVjF/s6b5BwrEPSQHk+N6adelNXNiq5pxJaMX9yEirDT4V1
ut0D6UuEl9203a2+mC7sBMUMN2FiVC0vCmoSaArTU18D0xHtkLarT7cb3JF9WtZxF8cKP2qnmS/X
dtleKCc6C15MjpLuJ+ya6vMpzHHoiouJwQSiur6e599W+PXBRfBpJTJJLNI2IumK7ACDuA9BUBlj
Ti8XndFcXtDubXzCOc8a600mpXlD+lgDQBUHKhOXntKE+VA5rp+sGhMHB/QilliEcT7cCH/LWcKP
nVIqPyzDWhbxFxSCKaFDlyvLM+GivBzWBk1fVLb3W+eVaKdq8dSaj7sz1t/v2NCL53dcdtXHsSKT
wf042uQfAjwnMPQJaNaEiljb38B8y63PYpEg9WBKs4Jy0LzZ67B8cHeX7yi3ns3x245DZZSMa/Qa
cdtg1EDY2TV8ojpiSUpFj2kYiVXH51KL2qFdXa+BcZKMtAeTPiUKPD6JExaiHghb/QjAvXZCsVLn
W3RzgOqv/QGIIuNyB7Y3jDzemBRDUNKAOIye+1bNRpFEUAEhNb1EsgWFuDL2B0wjsnovDqNc0pmc
eZkQftBWvk0bxeNY6RNfY/rsTNR0urWMyTFv5xXK5YiuZNP4bGJxPk3dOrb7V/bMsKvmk5oGDT5L
5req84lfch4ElEGgLezMIxIyxhhUTxZFBzUtcwVoCMeZghkaFRlQFcl1WMlD3FP0rBqJ6t0fT9NG
JZuoMrvtDDTCEbAfb3RRt/YK9ATQGxcW+OvPb52lzVD4Tdk5ipyIk10X8H8RtyxufQEYKaOusVmd
+PN+DdUH0jdGHl2aAs3mC2CQPx/MD8FmQ2rNvbdBwRQgE9XPg7afxr+X1MFU+/Mf+uHFA/G91TXQ
TDHwA25g4+ADlFacX/irnNjXK0SgZSXtx09TlrbjhtSiAvbjtBOp1LftR5/L7YTnifZnVo3QmNbU
Cu5aW70U9GII4E2WQ2xuUyJbmJMDrUbwboUE6HtKRGgI2sKjqVOMC7ZpAx4pZ6SsP9uJu2sZLzt4
cmjm5fFGojBCC2R53IRYxlMVKNwSuMVltRxIUjhSYBmlwzhVB1Qq1I0GrMSH3Pz0nX3fOnFnoO4K
WM+hzmVa1z+nKAkX61bGaXCHGtQnxxCit5AGP6fBzjHECah8BYjh3B8dzk9gvLaipKm/LXGCTH0k
YVEWbmwvyt4P8iK6SPFzIkY0b7upxCKraOSNJKIRp1X5t+MDAEKHhM9WywfEMP/gEDn7Eg8eTufO
zeJgrM5PLky46zmTme5QoHxGIr89ufYS+2OjwoioK1Fx09p2ua160gkauta7NVA6hUV488dRBMrE
+f0WwKFuvTKotWwxc/Q4re8a3kuXVB30AnYM9ZHYkpIwk8wpyNV6WKiT3rBNL2XgBJlpwNqWIDZN
fiZn245tQg6wX6GJ9y4a54HCdrFL2cT5SZTTMoKUJCjlWrHFlL2hthkrrGIul2Jz2am9CyQRyWUY
5MPNbUc+nQR5QKJwTJU4lqL0DKlgP+ir1iSsmMA+UJTnMxpCgxIWPOE9wSYyXN9lGkJZU+Eo11Mw
7vG1nUScXwluEdBUfi26Y0W3/cKh9fgWRcGd2fnEYP7dm/xqSbFY/v2TYN5RjJWGiBvjE0p7Y4Fy
6xRrTDajX2XLo123VnOlUqKbtrr79KnUvjD1Il6w5Rd7e0qu2jjZHoVf8q7EMTXhI0ILEGdQ56US
UmUdR0sLRRGaqw6aLd4fzIB/gkbrF3Sz/cOMCfYtPlqci+e6Kit1BPE1KLFNyIEswuIUsfsWn5BB
PYSUtWMgUIFWcQCzuQUGjTKqYE58NivFSXdTSH380lj/E87EulFUWBwesZ/r85xNnonZj8X7fcl1
gmvke2d+D3jgdUGdXd7/u86fysqaTlXHmiHl7XXLmPuyaBMY+h2xS0lrDLr+Uv0u6o68LZG72f+p
oZPZ5Pd8KU3V1Vm73vuJ3wn4OCyofHaZdufx04IsVhM6rBxHYUR0IhFehU9Y6Ctx/8l08Mi1QP4S
Loyo/023cNiI1enqLns9H1m0gCxQMfWN6CpeAiA93QKIBOd7bX58oQ3En7kvNk6kAbaIyPFz0U6y
Sx8fgoi6PlG1NTj/4Q0Ft2kg648utDdHQI4sn00jIrZmNlOt5rPpzn9u/2nRNvvGBwS5feoAtCOa
k5yzJWXzU1pbiqnTIgDcfEMaIoXRXXKTB1H7TiRoyTsXDf8ib2hXDHdGajPRCIH9zmxoYATZFOzg
TRVv8btQPn+vqopoN2FCDzQCDczx08SOsvI32jDaZyVWig/jCpA+Xoi7ntAmTctmYYohTMFTguPR
3yQy4yTHkuezJX8U05b2JkRvn4QCNwchg22mQZYN+Vu89yF7fXyP0p5Qr0FCePPKDgBLaTtIAGjT
9tuu7xwrVnTQJXVslOOd9ioY24GldZrn2DO4UUsjNAn9zyhkG+kbVk7/uLpJqiZviUulpHaBOt7r
uEml1EinlNcvHlF075Ux0K/i4KZUHSpL1SnuI+zoytTuEenkxJ4UsOVmpev6sSN0XMUdEbMJ3/L5
bTPClRbnSQJzGku3gg32naL+lysraRm0LTJEBLgJkYpw2A8skAUH0mcwqVZkbJ5GwYp2xQQsaiG+
ER9pREG0SzPVdi18/5dj7mZieelPQG/58vqX81wYbmC5p5mCAs5ksr5BxqwnziQC2ayWLSjlYfPw
dJPxJytrhAXd5T7GW3heIrZGvYLVpMbQDb8tRP4ue68Tfgme2sVAr8qtShQvbW2LtCg+a/8PD50b
iEQrKKzxeieXa9EejBisoKyWcP3OTHR9cQAh7MbO60+tKNPF7t11OCrooOubC0YuzTt7BVcIDT0h
uuB58fGWuwrCossMrUqOxgNGeeLADpkzCCfuCBSmGbRfuSqoM++4Upy9MvRmdDjLj6yRDs0UfK03
0ZAg3AjYabBF70EARcPD+7oeXgh4xGN+dteRDuQWv8lc8CBh9heLcWwmaX31B38ZhG1s6K0z4a6H
2nAiNKNwQ6s0GZJFa5ZRU38xMB63aSSN/vGwW7kLV57FMtEMaU78XPSzCzy6Qk3efdk1P5lHJI9u
yRVqgIN5kzdctuxvhxun12OsT8p6ehyJ+k6w05xhM0JKNss/58bXUFIPGRKR1vHHAwyWijkYmQmf
Mvmad821jXeFJg1AEBj+YwYhC/0mQH04uEkag6xEyFrISXsK9lhIoX7XWCZsRgy/QOsdvt9OcRwi
wJ7UsPC7YDlw450uoK20ohmaMxytsk7jwLkRH2M830BV0li6jDfZYCiQar4UO9N3ZMh6DUL2cgIc
DuFbl4kIzAuwz2QdTXNzzcEMnhJSoB0XEG5aEiPrlWQUQi6n34wjIT4ccQD4icoHZOUMMRl537Zd
D1B7eW807cvllaH5cGfxyvqCjdjBKM+IWaqj5Z9b9CWT06QzIP8XmlGfKGOeuPfu8cK+82ZvfrGk
b26tPLAiJCZJr4HD2596Y4h8RyILvTj9ywC/wiPTQpdUNDUBAfF3nmafRQ1lnVTFIaIYQVL1OT+m
qpp0IAG3048gwNp8Cnq8XlJ0OolMazBexhZZX3sd60mPjM1sMeiwLinJSnat3CNIYHWx3DM4G3ll
wIIQIvdSaGAogpuE1BwLs0HknzpT9uUSwOFvwNI+lFqGtbi+YfRHO3qWGTo0/vqTOfS2A8nHt6Bv
MmS5uX3uIGKL8mTL0mfbZLX/GHojNzV4tcFF0jnWAtIjot7KCKgs85AI1o1RXspDTIij/UHSD3b7
WYo0vunDB0Z03QC3oFUmjJ6ghAzoRSFBr6sMEDhucgo8YUzl4qHUMh19WelT7lZjTQl2parFDsIT
6sEuLiOpsTUmFTt3xPQyqnGzSQ0AS+fDmcXYPj8QyqiN+rgVJ+l0cC31XcfUi+WDImlI2If+23XB
g5ifMR5q//vYz14aizRw3rxhvoDMTsE2WNTzEPYT7nRXZpf+w4O8ac6WX7DTRcUZd9lE+T/5m2Di
1YG5rHTYBJeSHJlavLju+uFXqpToqRrBi5OLP2/vOFqnZ4nmKBiIYWULLPEV+O3zO+8py6VXQfSh
gNBCnCb0BEZTWna416ahznHuQEevlkySb1Uwm7YPZB0H7HblcgPEzthBKjxqGqnhC6+/84AqMx/o
g/Z08xvudkbnA2gp81sJB7iTUSnpON/9LgkDOUElziz2sEx9ZktMGoNqhtsx1sdfzLRRnF/P2+WM
pMKd0LDMlqfb6hNp5Z+luWqeuECD6yww7MK30txb3yWN5ydX1VNRcX5s/cftQQVUKFjCDwGA8ceT
RCzQK9ieGPfYhhxmD6phvSrmQF+4sy9YnV7yRa7ER1pEBWnxPran1tYM5djAqLTZdcNHngSUk8ok
GleV5Ih3W5Hk0jEdQPzm8c1j9QVGa1zQV/m6ldUPJnSzolTpx/Iy5IetD9AVwu8aUbND04Cply0g
DtLTpWpxPssU24JTnGfC4yHObVS/mHfrVIEyQRuaCrNWCVJVPf39BazFkPhsKTCqH0PB7dCR2Cqr
Q4yXJOymurjZZIrWO0AHd2zxIjxzJR31Zs9WIEqgP6kMz8s/0+HJJs6wrX/6TFq7UWhhy5pWTCq1
UZJVQ7ZFzS+5W3kvGUQMTgDZk7RqjsqNuni8ytYgAW6ChLzNQdd2qo2Jrl09pnwhr0vp2c3WCGrA
pcUEbnmMC0Yi/mFTBP5zY2S+9iViuJVopSPvB75ACorwZegAvGBoF/t9X0c0RTB8A4LqQggDXHSn
xGANV2hOfJ1YvrKByV2l7KfDxq8p698jbeTnelXZRTUuGhVLk9nqQFYs4p+a16qc0rVaS5ehdWGY
1cxQB+9yRZOW8lwRyi73g1NbvrN/KUm5o9twOt9FmrbZLF1B3N1oqT+fYm3WlXGG5/YiGWQK9vVR
ymSVViFNMN7WgxfrKB8OLnZ279wqEBAWJOmwIMDssmR2r/LRe0NCT4Bpwk1Tzqpew1ylYaEfzNU0
9rs/BJj+B+4C+Q6NQ6pk0jHnuC5QG4/9VJZevk43aOOdio/rW04YSQ7XOPQrVFuX9XfwHjDl4S9e
FjKpQ6Q/8bapUsrbXztWr+Y2SYmqwcJPbUev9SedSs4h/FYyA20YWPOAuIpbVhc/Q8RWP+Kpis2R
iE9pJPelLl+/G9FH9M81yQIHkSJ78Bzb/Q3EmvbSkR2KntE9DGpatHp/kOtSVQSklo9vcucX3Gxp
X9ADVngkFdIlEnaLr6kqS/8+loQ4+v3iScyVdXHfiQF6KZonTfG+7gamwoNJ1Lsmh/0nV9DtbtgT
TYNFTnWOmMoovqiLerA91ExRWC8YxAc2mNUlo2UEOAiH5k5dbqfRiQVM1id3OIPlHFHj3t6TqF++
AG/9JaLfLQOBEO60ZEKnQ9KTX2SlQTCyKTQZMKykSKBhobaE4cJ7/S1ryZhGIBf3yNJR9eE7TwOS
tyx2DCVZVCCgOYt9bwUcPdQBFDCV3+aA2vfUEyJTzzVH4R1nVcI+4ttMQmAjoH2lfHlKmEEz7XqV
epXu3Fu24A8DYJfhWEdhLYRViYqJD88UpCSQw7gRAVUr2xpIOtowc6hOHeYP6+jtomXVicjJrQHS
8Nmrj6mWA6ia6u0F8Ry0WjldrlF7/fUE0Q9hbMDgY+5UraGEkkhaGQ5M+HDBqOhzkAnUE2Am88tV
7S/Jfqbtzzzt+HnLYvFmoX1Meew6GqcVEEqekUs6jZl1ewYmyMHWQbkrrvXvwuRnHdcMXhl3mP4N
zJDg65KMFyXXZdb7mUuVxi4NyQfrjkEO90+Z5J2Nd14kSTG+3wNkCoYg88xcQ1VYmYlkaEqbMPVv
R5WwKh3MuZ78nph0PPvw+3yuybZSFRvxUbGTqV66tPKtWhBUktRcSjMXZ85eu5xsFHpnYsuN3aDB
t35CLNFRn/yoURMYmSTspOtkFT5pMrnFAsDAr+e0gqZT+nGtIlDSx/VF+gZvojKuvCIyyfhFWxc4
l0IkGexI3/ERFHHJ78SsAEdYTSsDDIzRbLZ4qozay2XaYXbOSuDJUOy8XihK1u9dQ5GJ92Rup6A+
xZme6UXBwmvaqFq9NSukji5pLEB4lOBxBW5mcp5MCeSwZ1fYQZqhsAQgkows+AWh227D5UjK3knw
U6RtHsB0T1rgWwzWhgKFY/p2YkWhXtLKbsyDs6gvNCpMuHTe/ZMa4nhQrP2cZlqSxeuxjh9uwNnb
BlaEcE+VUhbgx4yMZ4fyZnXWIpLQvcWJXIBf/NjiUrb5HrP7dYP40MYQOcgzSX4bBuHlZRt9QDnk
AMN0LrrsacWZeW2OVdCVQigj9UY9V26slgYAbrId2ZUYjxTVk8pTQnbVbBXl4i72zuiNETMhVRI7
xRpQ6TAMSt2b95J7oPgPurJB2gTtNsgN1DgKKQLFim1nbFamCzxG3k/l6cUW81UoOgH8kGsVn8Tr
8hYeKIhDxaaCjLGIIED3WgjwRExtOVYvyZx1JsS6ujUTyKQXo1KQcw3EqQmGUJFUzdO4ZM3vRjRs
YgkFnDsU/iddjTWSBw/spVUv++qJDeOu+0cOxGfls9U3b+XlWX0g8wFrOzJIpAN8k+19zn4SX983
8SePtiAuKv1/jBlGRw3bZ5l8g+J26B2AxaNSlNCr1qIgq1ZqMah8+EKT+8qAQTK/92b9F9pkZ3cV
PtR9nLGyK4M5GG8wztiKrfAJl1UwMkDbAvgHoksXHsMUXnwMuwthrkrznb5mha0XfCMZJIcpvCQz
CQN17WbGX5y5LLh6GO66CUKOpW+W6L81+IOjwJ6LMec2F3ckwtT7fQhbBH5p+3/qkiO5OeSnanfF
bKkJv1IOmGeVOOKZAgiaJCrvWxT0o0NQnZj6PRkV5eDpfeipyuNZNsn/z7okDUUPIwLtrHCBXrKP
c3dxIKxFgVztHR+VURqdZw62GLtaBol0xuIVOPdLLHfjzlKFtgkO6cS1Aj+jhIHR1xxhVwy2HtOs
EnZbECA7xAc3CuO5Tj9FKYr0r4u1k6o/t8Hn0Er9N6dA49iR1+5sALA4XKlWxUGBuAqoHQUXBPdT
4uLSGEJZFjgjTB4UT2qlr5krtZ30zVfwTjm9dkVxuDqMnqjkaEeEumeS81mMRjoPfkuypNUT7/1D
D8sVq7XLxrqWF59zX8egKVtWNC30uZbyb8zVGTrxAfeJXFA3u9OLKyH1rsZi9kkiZU6kR59FitpG
PwZNd0fmxpOutRuj1Hx1U5u0fIHrbHHWvSx27mLSSSQXtq0tkiPkKgi+Wt9GPFRybCPwjCuu6Byl
7LfWId1I9ZPeALzOuTqIP5b6p9mh6TToJo3qQYnWV6SVrVn+jBip2ag53DZaXJaUABZtIFyOGe8b
t9Xa1tEcEyCKHv2xc0BRjoazarm8BGvBx95veWja33TkIAv1BNb8WXvP+6x+nNekSUEYZ10tgNpK
Pw9baehAnPB0ynjJJ0zkFPhuThU+dWWNIHWyOPNFXkLNgQXTWxc/ZtMs6fprehSgUvxg4x3uJKr9
q3BnOciQlXJH8vdMV6bDpPH1mRMRuuNk1jxmlpeYGiqw2hKeG+hSJGSYQbzxwwEMfCSLcQLb9m3J
RXjkiPg4PWD4Gs0ppy/orcJKN+wJk8NDITThB742WfqW9ynpuMyREW23vkFwPLivD4qoGhYzlIPN
13dYrb6JA5d2/HdI72hK7fKbX61KrjTkQ3/RrYG45OQ9S9kS1g4CuwjwRrYi6IJFCOnN12FD4Vdu
Fr8DNZ6dcReVDYKIYA8tCXxNfER4PUf3R6Kq6xl4Je8VQ4PnJe0A1F2XiRplHTB8CVk4okJeDD/e
Bz7w64YlQAiu07KM/splqCgtsF+lmvso1PZts+NuS2mLHvUIrHbFkssL16yc1cLkoiOLdQSsH8el
Mke/xZq9FyraNl+sQgN2vmJyJNAFuj8sTr1vTNGJoow5F3w9Mafu2wB7q2Fk3tr8813ImMd2HlMW
TB9Q0a5g/AjmK3Xemq8o5ApXNmM2rbNaF34acX/+cGBTBQzTzp91c/PKLUUYPc0eRyH68HjaSdMy
tRxAAiGC1NAVo1YGomR2ItMB1X5FR5ApY8e7fTyKO91ekCpMmRgEVmn34E3z16AdGfmI9raDRFWe
JOj4kUZmNAGCgo95tBVKmCKew/e9BI6X6jOSrs+0auxPO2FWpr9ycyH4063TTuhhuceCVScIc8b+
kq6hUmKzjBflk+fyDaFG7alCrgYv5Gc0EYfcF5TTxTNVsddM04sXa8Ktm4spjD7YsGOMURIuN0Wa
qPCAazhea8m7L84Oz5ThMecm3KogZMbU3WemZQ0NHxbkRr+GP+rpkClzpwA5ycWpmok00lK8Hr1E
2XW42BcZwerzcfhRCteGTr4r1ReqnglYkFagBE/9FcEyi1HL2IrdwSOhiNAwMVuvPBv0pMlu6GuW
7tcCRPCidwbsQkt1vaxnl+kr4NIql615N9xPlvDwtdj6UHQzJGWMDu/Zqfo+md6TtqIEHvHaPV92
5x7q7gTnHM1oVWvVljDMbdidvfxurr5q/YRo8wvvB7S/83znjEhgyfCGZabcM8ZaLw5FE4cyk7gW
STmcc2hpN74rQSUaF0yUtlesKheXSFlXVHsiZIqT4HC5lbOu7NC2Pr+vgb0/ucmaPgsWCvxxPjRd
RPvNSpjhvZS6hUSsKAVqY3c7yN6s1I54uYDfC97ma5tKdLvBql79YinDA2wOXS410aePI8oMDnkw
xRbUp/8BZ93hbUBWANtEJINKj1hHXnYAW+r2TcpDwmMMd5UW9WbVuj8mXF49UsXiusQ7dOTW3aPc
eI1DVW/UPvZWPzp2BmE+B0yO3rbGC7Qy0dvn54BfFDmRviP4UtpllZiuxJtP20YstyMP6q6s+swA
W1ZT2qveSQM3sd2Kp+stTeJz7vVcZjN1nqxISPXuGStHtxZgKGLINd/3Ct0vZ+4reR/aRDiEr4Oq
CQWkggxvpAkVroULQfZWY8M6hllWGHbTIZZGwhk4g85gOTPHkOBtBSFbmOYu+1tkfejN5xdfPFaK
EekgGUmjYhlhW7c9SJcOxr6/C0267P36BzMFO5E1ICYr3nM2aV3AnQMSkIOg1dnFd6bUbNLEGbZl
OF9xD101UQKHXwUE3zZEQU4qUtiGwzWz1sUGctU8mqKrKUQMvF1p/YXlkni0T/+fCkuR3wAWDcAN
bcSRgCZGnZjOTFjptYSp0JLUoh/9Sh3aKE2/qHqnjfSPZOh5i9lxTJLHUn7et/nNqoEVGIKXXorI
gSM38hA3jbnAYXBOJAVf+xjVVSl5kaVD+yIfN/r6BeJm1k7Wo2zKbfTtsiecW5wN6WSFLRzAuSZH
QjOG1HuKzmUsnqfuAvQI6iGFXFHUNi6Ozvy21RECIV4Rsty1BtzHPu1k5PYxfxXWcEdbLx/X6NiP
bFax0Iaib+YnQmPj7at4OcIElbO+L6t8A6E/+eL0Rns4WMPx/mGPhJyulXxPTKJ2/q41en+g3x+p
DN+BjWklrJ5d/Cs/8/yB22Stv2eBcSE7KUYJdUE00G1KvcBbnkUOgJ9NDW8ddIayifIloa+T5v2+
dvNmq/D0XEMtS7CGLXWI9vzHH9YykvZYnaYpKQKUE7q6Ko5UVJQTpJHlfezmf7b1UWy/cdFbse5v
6W2DWvnhhwvzuUN5I6mg5uesSrbmJ87Hq3PsMAyaE+rURNx0sC5hml5zKqQfZytcvAHldOAlY/+A
0Jj4HnMvH52OR1mz70mxL+b/i19JHjNRY6AbCkdnkY1FEWZc86wx+hvC2fcce5RhfEMbysX67tMB
g1RoPivk8LeWguQoLEKd1wdIOkEKb0vFvA5hbtwCBMEhyg/BNN20zNMCigH0Lf1WZE9xSxqwk8Dr
LppaynZ3039r1LAL8WlLQD1t3PnoBeRhULFd8D0J/hU+mBlOmC1KxrI79bgcj23dxKnuCAS/yEzP
z7EVh7vK6BB0dShh54YeKeSv03HP4sFcycGjsZXdrSQoOHD5X76+ILAd8bfQVosbK7YBMzoAAqXa
546+zgNalDKH/6KR2oCZoj6B74t02o4shlMmg00TM1Je+DemQo/oxyLXz7WxBftPOlUYqBYeUoVS
poV95Vp5Uo76o4WIJ6pdami6IvMKn+htIPaVduokzhauF42KZ2JHMG4iecKOmqiDOMcEdNT/6vUq
hrNCDU8FTOKGboKqDkElDNlN9/Q3R+mZHU4YQX+31orfMCL7kdGdCU16bmirfHTPNHoDL5SjhriG
a66Vqdbd1SCWQa4PrnWNx4DQeV/ntsmOalGIWToMAcRPypNUvWSRFfbZYcgs2yVYVxo7qt83Qfqi
g1r7xJFXBo3P7urbTRnwS0UgmJlInNKhf4xcP0XsTS/q4IOOo1Wi3ZdYqlm9r25MkSD4ExsSA1ys
mhipenfanebPvxdJfLwKkVCsKR9gQMQdtE3KJux0VCklkHkxvvbcsFs3v0Ka4lc2gQgafcp4hKVd
6xftgKDEnON/aEUO4kZNnwTSxABvsHIhb3gJpsaYX6RvhbgIrsyB4P0uKg9ccKgPmllyHK25dEpN
3wOZbdJ6LHypF8U9aDPbxotAbgOV9oOHbGDarrpGH8Kruiw7V7EaDAq2Rvn99+z0A4Noz1xL/oui
4F7bezj68sXEOM6zcgG8o3RqKUNs1xMsLEBs5OvdwEGLqF21VBi2LEMWKbKR0OvMupCOO+ewiBV3
YYLKnyO5Eo+CK6kztIEnMyZbQhYd8APfWcbEAKOeA2q6BmbKczs9NiRTBaiFIpEjzcxH5e6gu6As
NlH1AyWN4IY3GMeFcEEl42n26ZOM4kN5y3fdUwCpcUYQH0s17KrGf5GT6JWpHRCkbdA6rBKhX14E
eL5sxEs/5Hvw0OUpyCQxcRgMPPKys8dmyh0Xk50hMxf6COi/leZgj38Ux2eHGtfHMak/ZwxQcx29
b8SY8XkOmHp8zGFpncoZjr0II2m3DbK5K9Va1BN/N2DSYmj2zv4tc/zA61uoMYSRTUG17lgpVMkP
hrUneaW6dps0jUR+pmDfO5+mkuQbSZOlCpG8ARN0V3rmuDiYjnUIfFTNK/UbHnbyCVoJoZF3wlR5
MlD8yutM4DH55CTXntiHkGXlDF0XPZ3Cf0eiDBBmmVF0F1jRAWIdXusKxt6ICmrtFTZZ04sLEoJG
TsA6pyXD9v8hS3UVnclXypc/T71lvP1Yt7oJHSp9OKUnaCLhRWyodGJKkydhoRgJ6++vKQdnF27z
iK35Q7vgs6J4bi0GDtXBMwvgzl+P+m8emAbSMxXchnHlezYxz1BdmV09/s+U5ZyyZzhtRahhpihY
5MRywqzjED07G0p/qKWbkA+AOmzh13EPZMUnJg5yJ2vSBjHCXXgqMpgnR0RhmoeZuqLAWcGv7Jrk
CYxaS5wODpbvbGNxwjo/Eyef/vHS70icB9APGttueCG/uCIwztDYVQGk9OMAW7bsDbDsNq08bP1+
/jRzymnd0k67eoPDaHg8yOPfUtHCrGiEOOZmGUcIC62/20PBuz5RGZ6sjdH0fkrG1uT3O3/P3aSK
5+rtUlieRkMaWNTNIe1NTlLGuW1gf3BOFexCHSxTG0ABISR+HRgaVtozjQ+ClVh7gDJE04t/SHGN
b5dHaXF6qqZZxLCbB5JJ2JK6AVbE5SWreRusMUc7TkO7lrivFTjd7vnNip1uF+NPVVBUMuuP0JMz
QYaujEmS/eIWpFB8PplIGxruq75J2vEKU+tOXxm8vJfVOM/v+vULkWExXkWEMug6ojY8Kn7Y1/z/
+45VRoeHP7cOtkIkGaq8nGomZHM8SrirUeq+15AN2julZEQ2513r+utmwYZftRh/doOkdius3SSz
Timffbrd5eqZKxIzScdpVngtKb91eRQ2h91QaZBUMBghE5k0WmQfL4DlWv6yerMxyZuM41Orc/VJ
VJ3XyKNBa9HNA8eadOhvK56qFadCJE5Dd22Gk4gboS8IL1Of/djme+Co1pplRqLxHbHWZBm6bWhL
DumbJtvH++8+eM2dA8p+DfHfQGW1iDKAziquN267+A6EXjXDlEX5noiD9JqWLsndFm/OWBPrtZQf
cIW2MYlgV1hiwsLr8FLE2LHGhUGXB4nGmtB0fc9A3RrjjrB26PlqPMNV7ZsKBBPIXSAAd2b+G800
Ey6n3C2z3JxK8oUD/GU4Z4giKPsBfZ0P7dPMcKK7wsXXg96hypPe6m3CE7XwQR4p6l9/BY6Jz56l
0tXbD6utD1BAYhIZHAyb31nH4tETJtKjn+KU6edugtBlxdN946fRwZUDsD7xhsNur4n/k76XWDdb
taBeu0f0+4YQxBwdjOKBPWcuSax6TSH0XCfBS9YUsZV+Ru0BrHOqyj0LUZ3I67hvvus0rtfBllUJ
i/fV/9cuxTGgANzZ8e0zapnFckLhk7SFSDayVBXqkvPRprCpsDKKwnuy5GYW4EvLDognV7qC0ZlU
cyV1E9bJUXR2o0MZWWSjsFQszCKKVQw4CzjwO/4x2NDg1mYJ0dXW98KQXuQewQxED7sFat9YgsXI
rBedA7zhFJHgWtgXlP1/buMZFiQ8Ol1+IaHgDYgqEieg6z2cT1MMMgkg18HNi8VgrpSOQ6hYsUma
yb5nMJEVNNK2/tGjM3F2WBbXVF1A+TKQbM5qfrchYQ58W6X4o9+i5B34VMbHVw5S7p3uRAQo1FVI
3/bq0QPaYo6kbKQDyN3GE6Cqy5d4WFVQ26zCx50wlS8S5sFZ8V+gB2VATFGzDlFE+nMCVttx48B+
g+071pJ+w0HZy5U2mTvUcIPRd0klHqZzZRaEzZUOzngS0pSNUaTPDHiviSwu/Ed0ssYPx9Y5zyzL
s3gzYvoWzhoRkvvUIi0Y4lQBRfCCjaTV2U7RSAC48nDVAQDlmurX/PZpViALUGgzZ2oHI0kBuEBr
cq1Q3Jfnw/JvJUcCE59BgwDzQ39Q5WE/LuCEaLib/IIFimpVN0cHhnm2YqA5+o+Qotvojr7dWFj+
Dp19jz5Mqp83Poq/JrCqf96DbE4wlF3mUX0n44imoRMBHJI1bFw/U62S9vYvGPbQxmkAbStv6/sV
4KfdGynlyWb5IPgTfA34sLiLe9h+2ZMs0dGYL/VXWWkbc/fpR7npaB9BCT3gmhhnZejL3qm6Yp3n
9qk5ZYog2qG8rEwhWGGsY1sRcMvtMMrpqUg4AbK1egAOHybgw8JCJ4J/He1jfLKIOD78YTN1jsnE
aqOE28I4ER4W4w02U/w4/C3fN98IU6aUFhH2oTf+xmBhnz9NepFW8PDeH1Un+ybNyV+yXH/t0wBu
DVyeGwCGrBevB5tyyVpQhSY/cmPnyjMqhMTNm4F57D3AtAlJbXncvKtWBYWPZAHZ4CiMMeLRDc4o
Qkh794Df+fvEgRqlQv2zUDiqWbkMiOvWHcdiI3i38ecmR119TK57D5LaDgT8qT9ckY3SwVeRb3UH
ItMNaTZ4Y8Q0TzKuHsebsSMja4rZymn8gw1xcjMyKQSJ22dRUgKLAZ1BgPKwuaZwuuV6aqfkhIUE
ZySF4nEzujTy+nbmiMUpFFSkbky1gSD48dx9WHRBcQPiGwHUO+7jfvoDf8S2qJY19lDZ3w75Yexi
T4t3RrWebwX/Vzezznr39XA2WWDy5UDaQwgTqMQVyayfl/fgmpwtal/ufOzb2nTu43wWEAVrbRPr
aFlCqcjGuin1nQ/J1Q21KYuaPikgqBvlJf+4PuCxm30l0eKKzvyBagIxpLTclHSGM7yHT4krhxNb
9voPbAWeAYEcOrynJU9R4l2MPvqONp9JEzi6hJJbp69wJmLYlFjD35+NbCaE7rybbYxZ2I+HGHOZ
PvUyCaz42clg3KKWYwtLzCVGZR7vHLnk5sS14Af2J+K7i6jRTcR85j0VpCTE07maifs7m3OuCUTf
wOb0nu39+cAyjtF8qW0FOP0hQoYTpLg/E+ZNRhWmPaygb3QHR/4TVG39otP8VxqRbLZCB9+WLW0Q
5u4HBmC+FlPOV1sWy3sVHJ7Uvz7fsWHLa5itucWX18jKTbIi84rRpVAie5e30PVRRVtyRwCpOghR
r9CkRtMBbZw4+llRwnunxcnQv7hD0xJWy4cr1MgByodFcW5752BLCOumuUICLdCcmGhKO2pPIFGV
NobJdQF6YQv/w0OTAKt9D2mI0vJtoTb9RANEX3/QsIZPzEtZpdwboLeYRUFqsHkjQ2wODT9RqXNb
iaoZ+IcGr4nahphIR8ZvczOP4PN9pth8toAvrPrwB7P4rlsGwWY1q7sJud3q0HAJjnaEznQhmPkr
+krBbWIQxO39ixldb0LGvyrCSeO24c/fhMaipQhbQHagFpMPskcHXPsHarpTJAPlVToxEjQ9TWgI
26TAfLskOHnJEki06nz+9M0rbm7g1khaUInAzMu9azKlsxV30SUUsWK8E7T0eZImr0luTZijJMf3
QKFBfSstCdwfg5XdKb5AWikeopVHYiq7DH7g8w5EACMQjrjlEh7Tr+YIxAQUE3IyS64UR6t3/9rx
Dq+jM2EPCX4RonvPyALzQ7MCdH1OIhDlfh4xxtoUz93Yen2DeilGxB/79FgHY6vN1uHAVfSlMG17
V+0NbTmAfv2XUyuD33LzQ7LQaVaF7VAI2WarQtDL0XH2BxCkeHsxMCzxQgyncWo+HhVFPBdDvezs
GBj4duNQZULfwTI56VoW+w2CdcyZjMzIphTmt/WET9yn95SUY1FywJnl03yUmJAlp2DX0HyoLhXD
tMH5skbWIPCNbNoqm4GSf7sEUAzwNDfUa20n3zmC3HFjHYVmB23/NBcGpglP188C0liSELgkr4As
fnl8VmPOmklrk+fqGeD9b871V/qi4+jPnVmr/BsIWnA/xjVUXl00JFGMPw6cvXtH+pbJqybaYIB7
CCAq1rmyQ5vJit6c7kmJ931niBXdi5WqApxcawe32ZVHgAyrjTcLGAT4t3MT/QaOGECV11yxj9Gr
abN4zEhsuH347V4s7nI+4JB/H3C16JKinXrayLI58m8G0GQ9xciWHJJOmSWpOTB/xxSgtaKWWXp3
99Qj7bAuEzWuuLtsRKS+mDsnkXIJbxAqgJyPNmIEhKqwsSUCbuCRpPa/+aMtvnxAeVYRyfusBlsA
KzzVAs+LexmSKeWZVNAxq0JydfdMRbWbV/0Oyp0+iZKgw/eeNduWq4blLg1FV50MVKwerRGMUn0m
/1oynVRcnKAMJ0MXvMe2fIhGcB0bampouWl8mNowlK7OGFBJVQyifJpyjqR3NubwYfP0eilVqmqM
eeLRv4T2MGMbeBr6pq/LYlbr5F4qkn80RLnNI6Y+/Q99iDLp3Fsl21zt8s2o2e9YYebsDBJnfExa
fXwMzmrNOqJY6U3ANtVHaq6fvasZJ0DAzWxpQ+E0a5b3DUKygk/qB9Sn1AANuef6Qt4KagECtFEr
yMft6K7jjIjYWr2cQLJFFfFLdPzdoNkGX+n52EEdMYGVuZzw1Lf7GfwqpndzoaVhkq9jmVQZhBji
hBXp9P2XnYk/SJGoGE51YabuajD0/JocD3XAGH68Qnl7hrFdKxf8Af28ZdCnUIljv7P9WljcDBs1
OcgqGFhNEjFPAo7Wu26tUyR8ixKzQ59W5LjKdFIcN8rWwaQXnhrvT+Vb1YM5j3ymDUtahztgdd8v
+ncMnxZqdHUMADtLBZNURfAPhV3fK+02Xo5MCm0Ekt9HEvVyxC+9Juj9BiYSbt4mvqiKQx0JOzJH
XUEA2buz0UROvj6BCY9f3dHbb5lOSllfI1Y7x1UdUNoBTr0twnOaHMGLHjiiJLKEB/ckHOg1JaX0
PvlL5yI9UDZjzQYSazJ8KfaI98eiHC4sqIL91ZBXkh2H+115ZJAljtvX0GmZlJa3r3E0k8qTuwpe
xVi0MX+dmMjYgAptkWO0DVUDw95B/VBUVKDwGVdyAi+cJTp0oN7+bYQ4kogH0V5Sq9aKvU4PovEZ
ppdoH23DT+c0jyorkaN7DtCubcc3mmRLdgdCS7xN0Y+mPMkCRFzN1kyGrPRaIVcyE+mL7px5cDol
VLM/aGojITK9odNdQ9Tu8Lz98DvI1DaVeFaldY+S8j4A6DKnJXmsyZZnQ7IuaNWPETylKyC06bcW
ymmPxzwkHY4sCEHD76o3ZOjtsAelEw4r9K/326oqKg6Xm1jiCyXi0Wh5cZHFXlUHhlcJCLAOMip0
V6gS/GVlpK1a+0SPN2bMeCcqgj7KUPLHigFCmQCj7As4M+OFfkePEPGTBHkZMAaRJSN2l69nP6MO
jssFb9C0rtM54krsxc1zLCWdIintXwCJH33YYHwIPVotj6P4BcRKbN13/EM+gunDK5op8HaFrVEW
qoNFgJfbbp63DsRfbx59OmIQaSFxlwq043bYOzQadQU5UfnfMM3wsumeWAEu7b4CpCGmP5Cjpw8/
oqRWVaBQVTv5j/VB7d9ngnSDt0SkDSIvYIhLZ1q/UiE3lax8cTqmU0DgCdnO97ZofmBD4+8NFQC2
1guKZ/KBCgaKSbJ5696LbOR+aBAgZlHOkrJzDwdatJnyIeRnNcI5+8lWkFkC8eAnpH1taLktLrKW
DSfjEKuPPaKKg5Z3tBkJz4b8WocdfwjniUYeNUl+BhIdEOIdQIK3aN0r4bjXuRBAeU6Vbr9g43Hr
nSoNk2c3tcYVNNGGgpDab8eu+EAasjwAaFhC//7qSbuBOkQcW7weeQovmPMphq8krogOiSbd+45g
AAT/dvvFMnj9OXndxDkNxUrv9N9vJNv2NoKeTkUP5WGn1I+kQRt+WfI7ku1D1JuQkK9O5FB0MeRw
248TxayHtEgsfJsAF6gbCmoWbh6CknnNZbGVCWvF7k5m5d3UAgem5tfok3ziw4QvnpP/MA/JsF04
fWA3oE0IiEB5ZLWCxcLLZaOE0RRnGxjxh2vHNNq2AmpXeEXWcrBswJ9EMw7La7DIr0cLU3MeQO9e
IoWYTIXmOnXyW629rjQRfg5wIOQ8RoaXFZBd3hZyOo5isZHjTi1a6I1wkwCzHan65ZDkbQjYNiM7
eafV4QeCwj4kkHeVka0Oj+beE7uOh+SbAnkviRVShgumQVKJU5lRRoSe2d9m/fbmI2OnRZ0iPHXi
Yv9BRYWtzqcuO5wBOG8ZNXp0GUaq7kYhXOBWmy5JUp6FQ79P7FgnnET9BM5sMjnJanBEWkXVTV1n
p6YesnPyOEM4yVkEHMaNiy1H+0npDdTYxZz8CIrSC9CAlkJxnFj7bV7Zn79oGQKyQSnJe5sczzqW
LD+7U1gYfkSLK69dU8y2KXU0JmHRA8FsiOpWgw4zBV1EBSulYrPVQTgpPjz2hh5RXC+G3ze26wrO
yrLAN4ujtwhSRGHfxnNfHUdPmyXbvjnvzKa3EvRjp4W/bk+Ojqd7Q/331UuzaIl38KAShgUQVB4r
nKA861MrdjwR2/m1+e1cPBe6B1J2lsY1sf8T3gpc0Xzdgq282euKTxmGcKBjSGW4p7wleVv7rRr9
KcpiaNwLB3q21ep1OuxXqVDOxztzgzLesWMka9MkiImtFMkPMgAsSTbigXfO2y7ctBQG0HogNmoh
SCH3dXj3h7xR9lm9IW09HwH+y75h6yv4ofaXu8RbPwYX0hJ6A4VM2wpSwjOfHA+YtKZzwlwyoodR
jQco5zGJlYDIOpHm0XnLkn6L569NlehkrQbJLGVf7J0k3Ue0o3rQubHQXguuMK8JX+U+kV1fWuWm
jBETjA5mAJw3z5AXv6ltvjLAuuHhOYqjQxW7Q7KOl2flBtgYn3z3jV9ZHg0l0ltmx5O+v/UJ9bFU
5Gn80/BOdwYxy+Bs+FojVdqkjAvqxWeXqCfK4c7WewuagGDXIsEaP+xIdOMc7qSkGYEwjStbpMVi
dNAD7vYcp7L6brt5NhThXO0+uETLi/NZwwQIqUxFMar2KbRWQCZ7FTinu/ugqZtiHHaNQ5j0DpQF
9vh1Ph/vaFQapFvevqwkqik+QnT34zAZN8lo05sDIBxF7ED0MeywithhJU2C580w4jL2IDN5eel9
KcTk/L2Ab4zA3wBC9ZpdZqNYlU6ebNSIAzSEXZ0u8XV60pRgdrkFO7iObcn9ulToPLzLwp2iS3Zt
Cww79a8eD/CwoKlye20uNbQK5vTonptZqr9hzpn5BaVLzrdWASXe8Dplmggrb57osYgC7OOpnEnM
QB9S80g1jwcUuSyiY3RFXWGwmyXEdz8dYMq7Hw9fzznow0iXMbjYiAGpmaUnDd4AxnYffwaEZs6J
usqRTmTNz3Z0QWwPGFAcSXYUJAiFXX5OPfKkzvqGfS4THLUA6mft9LpJ40eOGFnjoJqODr9W9Zbs
NuELJr3beRG6lbOqz4dKDsks1IozllJOrHsPvm7txZtrba24F3l3Eaju7dp3Mc2ZgkYbOk8AHoRs
bOm2S5edKHQ6b3mpkKyYaM8IsACX0m+n2+wSdeQKyyFcRpD2Fpd5f9BsbaAutGZMNd98SHzfio3u
LjTvlT63R+NUkzpBksjYosTTP8VkwyJLH69mSp5nH9/QHCa08Dl8hvXLBWYSGEmz4umwQCaHlrkH
1Fylx+JmWMPaM9X+y23vtcN4NKFFTEsCOV7DW2fzisoE/sKOK4nb/9e392o6/ycNDEtjpCJxojyM
C5hT3mgYUa3d6AuZh5N8N1qgcn6wesAg9f60+3WCwsrm3zK75/D9KUDD0OOpFoRzS1Z9YYFxKm1m
R9uuv9Vf3+vAWhzJrJ4e3yTUN2qUxRoTXhwApZIr/2i1fgcW+BoDzld63rl9Nw9FNdDZJ7EG37Mm
ski/DcpXFdZpxCbA1GuIM+QkFoMwYNtjmXR3m5SU0eV2RAGUA3pk71Ol5RXTxjNm+JfZBQsbp1Id
f6HSBXr0NouEf+REiEQCljjxCgCV+L8SzQhQ8n8Slg6jSTc8GU82kqlpJn1MfU/TWnATdwgqG7Or
goDVvn6QzepDrTdbm8pJrMoovF6ZLnjXO9D2saJt17EvXVJfKBBpuxleDlCIFGnZo6z2mdmoQpj4
ljmTnO0TJOGTLbHKNjna6UxSMM9D3kCpIeWaVq4lODjt+zak4IjRsekNP6h+ELBlfE+cMjcJhPiS
205xH94UB3pK4g6CpGvE7yK4GoGuK/Qgf4subXAx3RTk/fzm8wS3r7ZJm0tdFR5DrCbeSw3FX1rp
32t0+HkEXeFuIA2t2j56Ffu3B9uDXiV7KcRdjsBaIkf5ZP3WKmjgZomXSGGTSbUf/RyukRqd3rrs
6EQx5lpdHZAeTBnMhIJ5tpMMrZIxKnhst6rO06kanbXOtPMwVE8KQdVeAlOkH/lwL623u/yRU+ff
LVajXpqEGnwwcoM6U22fU0jIKKpMP0CQVNYiWcnejsnE9r70CCtbu2Zn61vWnMKfaU1zVaT5/V9M
yy6w4PeFkk6pB3vC2h0rBtzuZW5uQyz6kjW4cIRZKV7D16Rxs9LOPdypyGd1uMIsPZDczYYb9iYJ
2woNJbllKAIRYnFMxcLgfHX9je4OWi2PVVzYHJW3JQXnr0kMfX5bSEbvvDCrlILa9Rp7zgqoIyyD
dQYoUT0eE4kICm+1vGGOL1bAYMm6t0UESI98J5qKN8uz1w17FcHyrA6lMIpcZixRp+7846rraQgI
2zMz4PZGsnzvhaLyrQ+AeCQeJkTkESZ4U715238VtfnNqgZzfmqIYDgHngnDYqiKl7uARQOFdxPg
LqLCG3dSav8BSjsY/OQFD/YW8zYirpt8YC0rHeqPG4RraUsssyVAJZ7oVVwtMCHXdsaau9jmRazJ
3ehImpkgMpUoJPf8u653YpTk/2GfJaJvTqIRdS/0CxHEL2KDCn5p+SpH6UNJnYWa4VjlfgC0z0+2
sLcdgkNt3+Nn4dWZF8UoQnk0ncd8lG7XXV03b/czf7Nx4xdt8ZN63k3CmyR8T5IyPJH//Vyp+s8Z
3yGUOrijhDtEDAD/RzXPI9pHaPYx/5/yTIxHOVWlO48mCiK04qfMLbcypVFQPEOIuK4R0kMVbi7V
gcAcv2+GSaJCQJF3Gj4nJyXRn7LobBXRGJidGGsISIMeeJ0iFc2j3DRF1rfXWS8nEoBsD7YBHx2n
abekLg9IQusdQ0tlAEenXpf2C6eUnDQ9tTkTcM9SIEuk+JtgTPV6TsK/rxQCzcWgvcYpEYnW9y6e
f7YezNGG7CzYi6H+cRA0PJf2wNDXh4C8LtXlN9Iv5/eGMNCQuK+/hz2R1EjfKgruyUOD9ucwaH1L
YOpf3c0Um27p+hhivSgLmY7FGSxUxhOrsNSIWHYRXYriAsijl37aEyaOMLZRREcIBDZruVPbTN+5
Gcb/192BAhFMlXfL+KwFIUuuh7iwtxsUORH2K4OUewPs7UP+QAKhcrddrUwFEwyGpKMIfT/zTTIs
WTrthizIeB0WnmUjTfn5RUJxwv0xwJkZbCz0Co0EjTS2J0OfW+QRpwrVPa5oA2vNcScYPLAjTLee
IA7BAPoXWckMfHUbiWDpF+MI60IzDJ+/yoTG/F0pSR5ox1zFhQrc7lr6hoi55s86D/sFjTXpoDeg
hfR4eSBZvPOwHUXgTN4vW5bWK1nUgHUAoqqk4koDBdCYkck4/QcP9IXSEUGs/RzyzfxddlzXHKbx
E/tcq9VvVN3hDNYhzoJ3/1Fr3jP9hMFbGEdt0gSjfhZ2mgjK7PKUPHDWHR9D4YBqcuov25wf8O9S
iAfd4bmHcuDIUGKNYfDt1NQmXmheVma27SKHENg85IZxh76KF/B1cMb9nTT8k0mMcBY9hDlHyErm
U3T2IOY9jm/HkuiCTGhmEUDwig6alWPDHHOaw6vN7C/vCge68+pYAB5bQqooRe4UKVsbphh1hgIS
y9opstBiXs/xABDbEjAvJ4W4xnqiY6e5YsKsQhC2FP5+x9F01Nqm9GR5v6XjnI1s9HSHOg7E8t1k
XwNKfYHSNYq3QorsbhxULAbMQHT8J+j/gA8t7zCO7b+eVn/dnWCPTJt8C2YsS1lvqmRw3PJmxzkQ
UBi+M73Uezr8wfGT0rKGLWbW1Y/hOYzCQRKYrM0RN0739HPN1a1wTBN5a6hXTSmzkuhPzN8yJ42H
WjTgw/Ht3lR6nNdur4dkbgeBikDvZjs6vpQudewNemw/90vMYR1QmY8PmBEtr9zj5Bf9KpBcX5EE
Jv5O8YvAyHWDrQXk7WgHlCoPwKRUql6w2vw81CYGby0Frfzo3XPL6H/SpVuj6BaKLE8SLAZrXkpR
ddCWgbLW9YsJnznaYqRfL2B1NjAYoreXpSvSatRcTAsdb2/V4Jey3PYlT2rbUpMmU9Tbk+Do86jk
XKdsPuKzhPj51Vt9gZ2o03S6khzvO4Tb8+RMlBNxu7KZS3m9bbIhF1JLqu0kKJRMmVLWqQrGM3/m
zborHDn0aMfeC9pSQpHBMkRfnAfapjjdubvlVvXezSextkQQQHa7S32D3lQTDbWmIPXxZdQ1je1k
PEjKKjD32CnggwAlVxAkYbCeg3dY3A1uRiVtld2O/ZipD00sYDbb5K5NXkRP81E/rUMcta8ULBKJ
mRJwes/ZSVGBNjzenTpoBJmP0pmSTLrcIL07Kvjl21WAg7GnpaOX5ByXPGv3QrW+1QEQMyQm6tQX
WdX3cAVPQEKdrJsreRldye8TSvjfXlAQtJCZlo/TPYEnHmM3e6SbOFmPyd1Mk+2BvVY6gIwXLUnB
TcH54XJuijCCgMQPBO1gLSS3IDfwq68oOwezqIxOA7CQ7vbHq4inBq0d2zFBGGkGClXkvEZ0aRHN
Y7y+KlEw60MSCekVSot3WiIOMbTwLcpAp2bKcjUMnMIdEH3umhJxBVSgrvw6hNWTu7is9GifXGpe
bzPtIs8VAcOdfzksGeo3SQ7QB4Ot3E7rzoJXnJQ+kbbHygxqukqRIpaKj68yJKwdZVIkZgbMDn0G
Nule6kRd3uS5DkAzZj+q7NzW+aufzX1jq6MlNaYj5VyKvU87EcLre4u8TcyC+qRFyeQd598dPtYE
RX6K1xy8tvHZHqG/oEmhGOd8Jajp8/Q+U70M/djdyD8Zws0Hzy2YrsTEB+QG78kVxMmV0d7xb0l0
7BTDdR6l8ojpxIDAmBu59KFTl0hubOkO4y1QjziQy+Ef3xg50iPyb4j7CGrC4yLzqP3wHc0fo6Y0
oBjZrnAdBRhDnRRQyUCoeqmeyifiLshyrHCEx93qW803WhGeHrYARnWSOXBvfjWSDIVXmLnipl51
/aS9rbqpbLOODP/t4z5Qp8R6wihB3GBpxtIexXoaYAiU5yjZTz1yRMQfG90dnQzAK6GMSKH1DjGf
SL16djOTgdeU9KrqC6bGZGKzzbmjrzp0ToiMdaf+2pPU4rjcKKGLPb6HZnsNeKw2bsjPpCSatl80
r+4A78VuGoltUaH1jTlTV9OytRhNO7+cAuxI4V0XwuIdfjnecXjhdaviKtDmiMvp+J73NQtd9BYU
r6F08fdGSZYEJ8k4wI+g1fni42SkyTsA2oWRVDmh2DIgNIH2BoI8iZEnSRLopAfZB5quiuovEAYH
3qjv7XwYY+KAHjbqzdEiEH+D177IsCPPGSCDwRNaRb7sO6zieOEAL/ZeKIEux8tABiHEMGrO027k
1i0ptGJd9FoN/z0XCwni+7VHboMupxjPTzwWJHm5vl96M6YEwZWQPZyUqzI/DIN+U4EG+Pr3CSfE
V/Yl0i4/+mPpy2aLcmEC7qmT4gT3E1ZQMkl99d/8XE1/lJlN+dilcDopvaApvvFNkOGL09n2L/QF
uH9zkMhJcAmxGuKqHR8wmjzqarDlhMUZuT6cEc6varWRU3/p0me3lOUen/WKzZzGmkTKdiRg0O+R
p1JUGb/SCRAz0n/qshZk3taB9yL2krlqsgqkPTxZyj+YL3knU86AUGW26m8JhNeapOapURTtfSq8
9Ecc8lDeydM6QQCn6ZnSJ9ZeygF6gXWg5JvVBw74y2Qja0Nr6/O4XckR+CVt7Ili+8+NVWHAZPRI
iC3jfSmSu/maT/h4lR6JYQsMYHpOEJwhbP5ddH75Q++VpqBjIsX42Sj/9G0rLThH9YxStmh+pCO9
HLecwtlbOTDLBBX0JNP7lCN8jnH5KL2MO5QvuTUVEouQIOGtmUxBUA4Fkw1of/eYgSclVHEccTCv
WMu606OKcVHRwUrqTXXqEREsUm55sCRG9IuAL6AiU6J82JAx8Yyyx4MHT8IIpRKI0zSSfV7i7KUr
HM4f5shOWHyfJVYqqgZ7BNWN74iQWQYOeIerYINmXG2jAKPWDx1G+Zx1fHhTrq7xKaBKZm6goBrg
30TQ9JoUFo9hUoafuy8L6SIxvPZ/0FdtXVw3ryVL04Nqz/7361op63ShJ/Us12tqTP+zHaios3uS
6NZYhgLIsiHNEmLQ4+vjjHX0kMYzL3k65kfs8p86BzYmQyiDaBskEHnrq2FQKG7Y6RvZ1ZY/usYc
m7Kns0utrWNC0wNKSYKq1BDkRGr+LYaqpiA4dxI8cZBiAqjBK2I5ttzezJJiT+6rT2aETDHf+W2x
bLhWwd1whvb3cZuzTmHnanAytPZ+t5TlWCiRWHUGS/Cn07Lb/7dhpiSMsBTuIQCOTEPSiaEH6W6F
zDgg0gQ8OFubbV+wlpa6n0qzBIIGI+5SDk1K3QDclqkhheeFcKRQo91rxZoJPC1mOsP/XthLeeiE
tGxseirlyvUTm2qgvEtO2wIJ/KbIb44Ige8VELqDwBU1Zf9ydw/GniJha2AQe3+6bBFCeGzP/dsw
0jKVU7HWqZHiQdMkmZWqDBWAedVy+vCUqyh1ZUTUg+NllZbGsNNM1zcuX7Pyj7IIs9r7ZZ46mf2P
Z+kHmt+IKjxC4MSTWY09D7KDutCTD8fiyi1XZD+vd6UoO1Xec/nvOKw9gpkcWFHMuFpxoRUBaJSm
K80P2CZ2tsCYN9v9IBJHpeVQjCWHdn3p3B3N9diQEtAqon5Q3n3RGUCM2rgco3m9Gb/BVd3lWeyb
g54RpaBr9yEeYtB0Io+Qs138ADLpPBEgODkL1t1OwYwr/ROYXokHo4lKgK55S6VeTLUYiOomi7x6
tB47Jl8a0dozQVLZK4ZfT5wVkhVc+Vyrj4P6FSeVAiFXi/yUoK8znuRGOvgC+m6OTeGhhqg+SMxf
XE54dqJg0RSN2tPBIWLE2OVTf9cQgVsGnNhO2fSWMRkvm6UIU3jUw8xj3t7kwoGKlum1+bCUUK0f
6GWJ3KExYa0s/vKuRIDgoVxBiu3Y+BwoSsWwM9qOyBzh4XtriU3dMoukK4XBWjsyhHUtZqKfEboN
A4KDm219xXCHTICHGRo8fhPc+zSlp5A3WB18vamgi8gPj7UiAIst5GI+pnXH8z8rlQbW3rPgugK+
+Vmv13Q9esc5U2FKRQCtEdkdpLLMqA2yhLpHxmyxJ6AnL3Tr2+Qxlolhj8GVlPWsNPXVopynvsNy
FdZpgQu4IK6IdyFTOd0xrAQZS2k8+7gHlrzHN2/6K6++imEzrruzw3rofQtG4EuZIaELxsJjs3gs
IJuksHapbXcdeNNVblOViKPNASJ0Hysnw3zk7STGxt2aTSLIZzZxq7bGzIlqXnsvIH+xsHJZiBVy
V1WyQRpQ9vGUT0zVkvXHFqHtEOiv/JQEmgukU1Rjsssz0hI/07cY7orkNypzJyQcanz2QpPTmId9
fTLkjpZTsiokHHOKMMe+vkgKztym4tdi28OJhlrxmzM3b5IHokcXZLtq6JHJVxs2MUoOWJo0NeXj
9A+UMT+azhjaZ73rUUN/nbtfAtdrmMFyYLMWwYzH6/nTPMu1zUTENZApP/XfxniqQI44N5akQPL8
LTeC8rnxW3h9tqLUY6zRNot0nwzEGxyzPRU1EwY2zYj9IwLiPr1UPeQ0omlRuaruyv8sinMEtnr4
JdLspFYtwi9kOFFJf66oH20+fJMXc7HZ1w8RwRgibee+GVo3GBTT2ginnNDCzIG2qsExXzMI/OrI
XTRf9L6Hdis9xj0t1KLrf+McYVho3CxIKH39y3hq2Cc0gCBzEWh4vB+B8Hu9rOugmvb85iJpt/33
v/qqowWKrwDH4djL1Hl2PSpkwzwO9bSg5U6/Nsep0oUgI2yOo0RIWsvX49sr27/MMFEHAh05RO7s
0E+shXjv+HYMn+/cfCoBF4nli7K0Yge5W0vkCkd/Ung9Ee5DGMIZc8rlft/6tJe+yvZY7zUiaeSO
6siHtq6aHZJX6Xl4qpAR3IknwojEut9JnOEpEB7hT3jX2VNAfY+AZlEIseIGq62dicN3wqXHvcIt
V04jPJ4HoeM6PKU5nsCYH+VgcDSnNgjBEgSzbL5FFlG138Tq495RRKe2cmVQ01HK3V/3GuKmTXJQ
XZIivFt7aB2OrN7KGkp4VJvQccSHTRkIZLO4un3waS6wic6AzSUD9TGRqSng7h1eS+QfhVvn2G+c
wjeUSbHU5m5pQ3we4G/oxVE5lwQN54r4K0zkd3GO0jXjyGpnlTKtBAMbGZBDqFM6GVWJOvLx3OlH
2BIUVU9p0jCKp1oeKTcN3tbpvJRmwD4aCF25Z1EGN8kHLIPWG3TngL45ZerD6H7r1zAP6kWHKzPs
ewbRscgumaKg2vTv+928S+QtEel7teY0BwV9ix/0fttqrXglssoQFxbYEBRErdtArNL05XwKihQ3
j45IhmTXGBfGrM5NGugJ6rPCbSH5sIf+/UEzw/LBz/tymBF616oQF2RnKinPlLjVhfgp1kuNstKS
kp9QGoYAPkdOphqtaJTqIvH6Thy5h46sXIa4cYO1OeeK4dZrCOktWJjSbcuv+DXJW9B2Yk2fO2sZ
1iPry1KfW1knnNx3CS0xhtJFt+kX7U5XWLMbyZIpc0oW2iUmWRQBJYl/fgYBvBF820LQIHQWTrZO
gmxLC8D9+/kzfzvfTwiRr9zxSndfwluZwXeMR3v+s54HoMMzN//nS0OFz6/nNz1f+QDXsAxPJSeH
cmBFhsZdnkSbdTRf+jozsV/X4Qe2dZnSwnwd81iT4vDhbyDT96FkrzoWgrbgF/jscBIIe6xGjyIb
0LWsW2tY/WkNnSedjQmJYMcGzQOpz5/hV+LOD7pOEI1/TzAZ/VgM1nP9AaGhCTSwm4CBrObw+XX7
uTLYXfwTYSxqiaQlNi5bkKDx+8F5SgoTJX5OJ9Tft6XnDj92iSIcfz/7/0Ql489DsuLDABHcNMKq
U/TxexcEC0pIFy89OoaGqrHiK8+czKMQGhdQTqS4pB/eZBHCOKfwbxVn2Rlh+nZUK0Gy124zqDet
uIpu3McEz25LCi4aMphHfeBFFx288kPl8m5VSIQFaHZ6xNebwwP6YBAZmmk+sfBZEi405KtK99lq
UprgnXL4MCDlfsQA/EDDTcQ/ombgoIWWRdRXagl46VrPk5Q4M+63PNuhiueoqIMg7rXpFfQydwq3
IyB5m08iYvgmpSGIQUY9hXhC3ySqWFNJaAr4rhsskbyF70jfSpXT+gdRR1jphslLi8uO4QIRdCJx
+oNQju7ScuiY3hI0jSXnehL16hBgQI14snflpQK83eGjjFlDM2O3JSaIO/P08ptXL/6fTHvMfrQe
xciuoqE1QoKUvGQEeYhpLATHnG8jOXueCaIru6Q1l/K6Ig2pdCdxRwTqGYOiY9OrcWRG2L2Ip07v
Dg9t936ky6kisNLMijFnC2rWCqpYSZvIIXo2DYnw4HX7qSJpj7LVTa0U6oblJn7+4lUC56lLd1oD
Ov1xo945y6vc63StuKYjI/Ww11H3RY80y5ym05MKLqQ1IcNgfJgE/qhtJ9FztoHip+dBB05cPVbQ
Ap9Se72xNvTeHWnzVG8vf/VTih57VyBSQDru9gKI8gcE3HTs2LNuAIDew7xQorky32EeeIDa6wL0
EtL8kkz7ne9IVWmrOKdmrK/kYGIy3KncVq6ivC6rhMDYuAIrrr7870ZQON3FQCDeOgaOo0/LjRDW
yrogO+CmILy6h1O8eZyrEpM5nQJOYH0ihuKwq11kZn2Wwo2NPcVFEOffpjOrzfQKkjPreSgJXE7I
JjKcrywYWDrRUYLC3REXp1vGycLpcNTVh4R7QbjLjua80ldVbUkkF4Q8ydZjLppKNmoInKnbsKKb
nJ/pYqOBmJQ85Phe4SawZP05TIkMTUjKvet1cXXnY/E9FjBDmDrD/DRKn1cwgMWtA+7cEx0IuHlY
1gKcs33D1As2oy8YrtVkfHFlpLhGR4ZDbQb1mhraahEjC0i/sTi9oWi/zUSBFvs3vpMoQkZ/seFw
RbYxce10vNbTLkg8vFedYzuaHjSfit/gLBAA2k3RwhLZnDytzRXajWiUdAT+xcnb1MQfhSW16Pl+
L23Lc8msG5CTLnnigkXae08mnhFmYEdPoITYgdYjmCiT6wmfRf+fbgmUTfFuU7tb3tkgPsFPfia3
v3T9l+jxplzKP+JgkJ5b3bpe0GWM/x9t5DNm6Rup4PcgntBg5XyHQJ23Z5+4VTCMVY5Sn/KbMp5Y
7E+laiZirOWY4Lb1jI/asUnkmtrzqtOO+xfZZSZmYD20440my2IytNCPXuwTI4t8s8gyBdz6RYsb
G29DmrMpPO+5iOzG4vTj0d1zfJFd9Cbms1orJXGKnv1Kg2P180Wf5ik67AXsXbKXJEdNtjSA9uMw
wR2uEQwPhoSEb6rO/q1i4pQEX5ZcBFcEVqqU41Ui7f3PlL7gUDPEzBFvDo4yTRXRCKz6qhyMaCw4
tTCby+j6hdyzrmjs12CsZTxexyuy0lo93AvKxsY+i+FLmh66KD2/3Wm/czlBG70oXIYtxpBPWt85
no/Uqx8tOve8GGa8DNMX/SNnlaJUZLG4sNyLfLu3r/A45J61tFE7aQsUecBVQDWlwUT8rLJflJxs
w8smqqQwj6+ILvh+ysykrCGR/aHxIkT+1BaV7SfvHxDLuIEWO8qz8JZcaCcGVSdTFeWPTle+SrBd
tSB8trf1q6+19e/EcuCkI58OJ4H0/7NDIXbtwggxBygtERHuje6KYIzUA+WKudorazaF5rp1CiN7
26K9ottAjYqv+26FI+h/cLJXrJaaxueuc0zP6dctWY8kwRTAhGUj5Ln/iQm/yaTSP+k0JAuqF2JP
Ew0xixOpF80VvkZyRCfiqSyRGoNJe2N4cerWcu9QpdRRY8Zw6Q9CleksSJGVF8sT6X6QqWxkz+PK
xi9wUlQEubSf0sP0s49yrNnuU8XDi3XZscsDnEyQ59nr0e+9dxj1TvtAqbHgyyXS4qJFDG+BDjqh
kWrRLnHD5rrskdX2KbhlSEzJvUnMie3pxxXJP826UkM+VX4SrQOkPR8kdBXxbWckBjDoQqHI5Kpy
WvdCB7y+hULVMuU+iO1Eubp0wecL3GI0RkakY+HO5DVPH6ceAyVjGwxjdTSKFVQHn+EmXjXxBu96
6UAP58qKIxCkOXHzr9sZR6CbLLLilJiZZL2u+UJvfggf3eCsaFjRS1LvDJzzjOgH5MsWsqdlMlmN
HGeNB17GuUUBElzUYzpZMNPpWGYSYiXbE13huzqUUcALESgY9/LszGs6t8l/sZaAJk5xJWtJsCVJ
UPIs16IuF82og4RZU8z4JJHgCYLZ3GUxK+cUC+ioPmVUGVLmo2RtMdJfnnWS1x7AdGvsqRDmKHrC
geN3vbEBDuRXyCQXP+R0smZ43vl0oBQ6J+pIBgDE6BG3WTzXNMb5fZMoa1JDtouLmE3OJVeeyQEg
hKcAHpCzmD8yA2qkWdhWrw7gUWbipN+OyH0N9do12b2KAIdnXjkonavIk82xO7X5lNqtxd80nwoa
L2dDr3t+hk+5XB+yqcUeLp2MQOXHjTwRVOpyIpEqv+YEgoJsRy/eD0uNaJnuDiKYq8ng21wT7KuA
SE6rH6tT9GXwBrBEyuCHYzyZri8ktauoeZWnCu4tJ08WKq2eJT+YBE3mkF+KXMwD2PsnH5pIZCd9
Z0Gn2J6DVjRZ/Ud+A8Hf6+dhqFvYxnPeD4ssUdlmr5vK0zfo4AA4hsg6BTn42EeL0oLpDTT6lI8w
1FhFMqqfOSZ20UiF6jJoxdb+wfwAbGKZOH1aXt1Op9Ll7eDpMu5ZD5SoBQbjWFDyG2g9/3ZHM1C8
QOVi3AHxW8yvBl0Mcr4tUoIN3EQZ72z/2mXSJajh1iFWLGDem+0EYRfqpxiYore+AtBfvsDc5zUL
4dZ5D5xW61dBRYHb78ayphp21NW4kice+DoI02gGtHxjeGwqsqiyhX4kAUVcwf6BcOWf1qtcLaEz
w5dYDelV9OmjYCfKGFtN33pK2+PGvc2ngw7B8ZKkG0jbkCLK8/B3fH7XVo5+tuvslyi0yClBUBHt
IXrqnkeY8OeE6mutXn8IVrLnptdwZFWXWyam0S0MDLZlrvhW7gUSr1EfwCVn+fCpezYwjkk0l9aT
XQDYDohoTCE3V4ZFqGHk4SwFOXGDf5F2oGLrgbT8tPIg4hI7iD2P6ItHyI4g6YRZzOwBGQ39rri9
BLxJx21L3YqFzW+RrWuU4X/Tfrsbsgu9nUerlz8Arx2T+fydKlJ3+dnXi7Sc39ILWCKJIaoPjoz3
gj+/4ucxWiNyw1EIt5am5kfoY6FwbT1zFB09dY48KKDJ9Ksuum9Jq54OqLrP3sTx5AOsJvYuxAoN
n2fyUt1P8U7qzMmNbYYhxVDhicDfCV0oWHcshvnL10YglU8oONylvzxdfCnNrYqYiXlcis6j821y
LtOrZM111Ci9bs45f1uJ59+WSJEZo0lhe+7gnBSFOOXcHKl0OxQmjpEtk5AArOdl7rsKXwZEfSMG
flDNfFv5yewslyfMy5UE49B3Bjh/mQA2oY9ofClCcKJO3zgkrfn4ZfrR2+eAdypzchCbAikZ+49J
HPe8Zwt7TYfrejzOioc7xgg9oFhYAnxN6OaZLLA4tTivOkrGC7vfMo5Z0ZafvGitG74xP7/ko19f
1E2FJM9SpkSA0PKh1yxQmA02KGDwY+Kmq9/vMqDrbQOfmU23HEHQ/lNTu7myvmD10HCGEds+DQM2
6FXBj/rv2zOofdNLGOsCTgih3PorC+lfezxc/YZrN6ETO6GAVyjZ5I2KA7udPiPcuEWOOf17D97I
i1vR/k0PySvjXGSTmXoZchOjwH0j8hJyAxIirs3j80rxq7MNNeHoLoK4OhC4RphALLbhuQOuhwwJ
UdDBJBF3orJgoQngA9RDBJr8WCjydxEwduTnmfXwDcRMAtrsakA9sAyQQkl+78Kxiqnw2wdXdW5Z
l81X/ZS34zow0pb1xokzNAafa4XDZQgpmXhEII8QBme2iJ59g86elLWZGs2/tGIog0+OmIwDhoBk
AKtCjrqb/28/wpM88Z4DzGZgJoqAgRJLJjDvmb/+YMGevswitna6mffQpoylyOfcRHdnryInNd0f
6ptyFI+YOulcfjzssLx6gcvktjsaexh7ovjMmlugi2t1P4kcNawAix9FvaBRGvRUo75Rjw1bQ3vM
1N73Ah0wbTE5ifuO3xjWH3XoPM5p84nIHicU7nPZzBRDj9hYE9UxNdLfLZP9vtoqap70DN6haDdN
uQ9qE8HvrDMmKFd1HMsPEWdvtlmWpiLc6jhEKCjN+H/jQMl0gDvxl1vwts9sveE9ZRP/DEHEOMHb
neeY4JmESioOo1RWMwnPEANBKMyN09Zc8Xf8VyeL+4PqoMJeQf1EiCuSyoXUInZ2Pq2oB/qz/V33
/F6gmTv5WCpNUV3RJUqwUz/kU3PbH5HJfwXa4gPUI65czxHibXHP+SWb/9OKPoPJZxcB1+7lAjyl
A9Abq+/mnYML6gp4hwHIk1mrDYtpeKQVdGylj5XZgDSy+Od7OIK6jzM1B/QqmbIbp2/RaDI2BJYD
Ts7y6rnvH5rGpkHX4aecgRH1JWAVLPAQDpWpGZ0lJ97wSH1YvO7S58+WGy5tTzcY/+6zsoueRVny
949mNeUECINBTIi06ykVcjGGpxOs8M97v8Pqi0JW1ao0Hz3Je1U00bzmkzRnQhCRx2kbtQyNMC8B
yBJnXiOnXYGwCTJWin+PjB0i+dkXtZ7TMiMJsmFiq0/t3+EtKzv88QzczAQzVqsM0Dvwn4CYK3ps
CFZ1jn/2TlFMikqOj7s2Gs/uODadLLQmfNXempRtcaYPsgVlRjKlEPJDG8+QH1A65t0b9PSVOsN7
yZzeyhetng8lWRPLh3+aQg4KgofRYw+yvx5Z/AMNxLrXAbEpfTjroTrLJ2YnndjpkGw/xrwjW/xa
gOzYi3IPCDfEarzr1yLNyJR74LRg1T7xsx12ahTovbPgnSohH534gFvZ8V7aA0R7N1ah/K+61DhV
6/ODXCVOeiRmuF17N/oEr3sWbFXoawRolo48Lc4f0TJ4JXtX8XMsTgI8coMJCGhY8wqGw/34JfPX
J1SYkoPjJMhd4Mb0ubeDnyv7/24WH+ZuWRO7y+UzVbJV1K/H63QFaY8n/y/8Ys6N8limv+s7f9Nl
GpuYSkm/qqRB4P3gScb7lNvUKYUH3Uzou17OasuXc9lXenRsW0uqUtdVVrtw6uSm/1JFkbKlIh+0
fSBaXeX3YSZi/Fwx5wOcpWO+ogEWn98gNaqDEWNHLj5bUDi2I1zBYjZQmstFR4spenbh6hIzvL9H
3/FzNWBvB5Frr6rcGZ8kTSzBMMDrV367nrctlU0tMpWv5Qf1GDcyIxMdv/37Rf2NK4nqKOWUIntk
VUIl05SuYMalMBscfxONd7XZPbx01BpwEJ996QxUQ8Ph+pcfvixZ3OdZ9Qnoo87rUd3WxCJBXUWN
5aVE7eonzOVLunyDozTg/WOHiJfI0iD9YzYsR2XRPGzm6PUJ647Xqj5lDzZ9g9Rek2uoRwifhPP4
JweYi+V+ha+84ud8l+iBJN5kRP6S9criN7cM3/Kw8FFc4cOWuMUMIJgi962D+FLZxVoU8vQQKpTv
MqEuCo354ja1XJcjU+ZfiFgnMbYdiNpIfgWFz6WBLSrcvRV+SOMfds+5erIsSplkFRtslYwDQRJt
v+Z2STbjQiNIAWcR4yc6OqrdNy8eNhw6bbxxw8nt+8o/7vQOFVB7jD5zn3Fhitca1AKA2Cme9SE2
UqMPuV5IEFQuMeSBfTM0EjJLcQ9ll7CoBDZV7TZcjCe3fUXb9xWLMLv+FI3hLeNIIIM3AntJfv9v
A0iigA7zmpVusvA4BLItSF2lhiu4O6NOgDPvi4g/vfcL0GcaxOCPItb4eExqBJ/qdV++15F4f7yL
hQCDd0SDnULscwQhGLI7k0mcpr8FOYPvO9rp8nI0g6ZCzZbdfei0ZMeH8A2YaSpoALjRcVHSKhRz
WFNnZy6BfjVwaL17fL9doyXP6OCSgTZ83nOo2cYkN7Ua09MhGHkfbbxRBPK7ArUqXUiMr33K5NsN
7gasULM17OLTxqkRkPBKrK+jC1zF+OTJk0C6bEyUKIMJNmedUMWFDrNpFWzqnZWGRbN+SJwSNIRw
HNisfYwCEG6ReM7J/bUFTmygw4cZRYjw5096HoD6acbW5X5XRwB3jOKxwtwRdStzlORGRW6FRo3z
joToCaOF1H4rxk5UuilJK4HsJyVIo2mRAktmUY2MCA2Db6DGx+/mMCn+I6waTLYblyfDa6iaFpCo
K1d6izyUw+5mpLgc6uCB48cIKdJMEK5FBUwR8Y0Q/geQ8AI2NrzGSiJBkFlD6XJo0g7tkCGvqy0y
5KH52Hjd1PH8AfRTpoA+dBmfzPOv+xkuSOd/uhyPS5aPfjhWeX3zmGeiGLfG4nJH5c1ntlfiEqtn
iCGRrleupliASOQsyTyTjL9exin8lNAtKNLrXxWivxC99HAOvmz5qQzh7y6/eCV0uSs1IdwTySiJ
2D1g2YgLsJA5A8pZylPsK7ovK9mtqHTwbjjDFb5XkqeC9LA4UyyvXwOZH79576qiItWp9tzIq3Wi
kUeWxydwYQEoizED+xxa3gw7bO9skHnKWIBZTIYVsSvs07m9JT3AQxollzhwT2QvB6z3RK+1VjDx
mEc3ZPA+gSaV4AZCsokV/doVHhuLPNmrDAFp/zAq/FF1m1CiOB58xCBysC1ZKd4zeeLP0mZStL1l
XFW5lxD5VaxXzZU1xWfb1PuPhtENi+QwQx7hmcwuiI7JM7Qd4Y20mDRB1xqa+IluFujIWt8ID+zU
1Xrn5mOiiaDDhFE7O4xyi4WJ67KYJgLDBF/+fisfY1RM8m973NIUPpliol9R0B4tC9DKtmmtQO6o
OZA0IAunT1+q8kJ8AXYdMsqiLHpIP7jBAdi1P4l0G/7MncrkxTWmp87PTDRG5XhREwWQYBZCdhx/
16je4aE41AEd+5uGRSpMdxn3iIVnT8xqivmJwE0eAkTylayfBubMbBdoTGCio+ePLn8tBYqLjiEP
10UsfHiyz80t+2r7dBp7NxkQy1LDDiJt8vfllqJdCqyQP3FlyQItvQfP+zzNugxaKTJ+m9Q/XG21
8uSKL15TYztrtjKj4rafsGoIoRWpmkMlKQyZQXzEn86OBHkSfP2pLsZPnm8OsYB2pE9/f2J4OMzK
S4jyupMlMvfGmEAqvpYtLNDYTGS5mrfIMmNewlP/PEEVSQZ4z4yR1IzRGC5F1tFUeAXUxHEYNIeC
jnjrSGC5768/gADusyZpyd7thoESOOMGyFRMV1Qs17BaE6g5D7+hGPlGymfEBkflI2N2NwgtwmSk
EzujZfE1jpC8drZOz51QLNwbOklETO7R9mMB4MDTII7FUQLPWIHojWkF021H/kYrULD02vCNX7c7
OIe6nPMlIFmdpQIF08GN9AtTV+zQeSCE1ShAY7UGxGKBxej7MkqTsQONh9UFvsZRBjlNlFPQGO39
1WgAC5qI2AmKe2xjxSDjEjT8emonj5QBg5+dnS0PeBPIfZOpUa0yjOHZZk+luZT8TmaOnGcv+WXK
drTOCOqXt6xLyomTHnMYKAiXCID2PGrnfOOtjcWlatAPHkbBh0oDss4F5VIXuHhpjgdsoz8eV9UN
2y4TFakAXlXRkzeV1X3Rj3yV9RPlaq0D25RT7Nl/cy0XNmtjbiIHD8KuGgtLOGIfFwZSiV9bv7x5
BwTBiJv9U2pbTwT1iYT4XASPeY3pE1vOqS11qT7grIHoXTSvu/P1w0sGCb4NPxlia7JMQhDk2pPG
3Pa/FhRGlovOMSwI+KOtd1WmlNFL3crhw5gJm8o8UGAhDvn/lrx7aRk6BzxHzIF4e8KwlRtUFXjD
j/DQHVddynQ2dEtAlLewL+mfZb34x5BmMY5M05I1CRkNJwU1LmpJoKVyuxJzn4HhsUtunHBj3jP4
UjzkS/iV8K1ZLvmlyH2+gNOS43SJPeWiaP99ddjHIuIJzTPt+ocUuolq8ZeG8nfo2/Y28BUfoZOc
7FoLOsVrFq9Tyc2OxIRwzUh0YhCB6NNQyp0+IS3qADb1Htv9i9Ael/V1BeWJHEqZTNtK4uXnoJ0O
9SBc54+h8uj0tTcPc2CmCLiXLUte7DgOBaW5HLr3vemoZmc8UiluMbo8txRVdQVgtgyKmph190S8
1ZelX0+pIAtDE+fItsPaFtMP5RaY30RaRC+20S2xV1IeP/QVPUWZaIir+XrIES+Gze5Lwlc5ifX6
V9zL1kWDNgmxe/gQRnk2p2hVHHQGP4imBp4AwxN/1N9lfxhe6Ui7K0+8UVjJ7xlSyRHZwQpgUBJt
zq580ltyokdfSDv82Sx2Kfq+jm29h2/05DJw8LdbTAPQ/DcRSo7uf5eQDAiMeo5nhuzs77JLCtBC
/gcoeZNP8T2biCU3QWaEza2pDbq4mbUb5pCt4BoDQINIVRqsMTVHvQyNyBaXbeli/K68o0JuHycn
Uu/Wp3yDugyDItQxUGy8Q6zuoMj9NURs2Ne8TC3r4Bnf4hk1cuJTSDInVPCsjRBIVJSX7qRSb8UO
KNNQMFKRmyDgFx/4AJ6UX/K1gk1VklXNDWKjl5H1DkEsLC1xPRsdGm8y/Dx+6/6Pzgqd3Xk6T9iP
1Ea0eK/05b0CTx1qvzq1cy/xHNQhtysuyFO1AB/roIIBFkQ98niqwRJtpaSDl3RwT44bTo0Q+/HI
q+IMijNgOi3znUhwfaRyeAYXW5uT9khgytsb/wYBd896T5SnzgJGLH0lPVL4bRCgES/+zhmv1qn8
QVmnAqDBIHNlcm7d6H8Z6MjWnJY5icY/HKAAeEHC24CDoorYaO8ly5D/2BPNi0gbhj1nWMPlwbPH
CmqttGeZQwpDfF5m+pPA7X/f+bseB2pa4e6zVwImX6L402+WAVOJLBydux0wBdzIgPom54FVRaLm
S38k0qIiXr5YBs1M6NDqSQZ2uAfDMOGbtp6o8OBmtMRyMPlKZmCNzjdLUo9XB8DNVLN30eZrFc4H
N9aLDrZA2YjhvilNO7fyqizZ+zK5l6RI0hxzjgOo079laTclhs914qlwum4X9HrwZwJw3Cu6JpY+
USdfenLx7J2AuNNHQ1k5EF6N0sAkSns/Iwdd7MgWBTMU9Ozd2iSTUeDegP4W7bRfASZ/knVEpeKp
fPqggDNMHPqyLrSwOdGpgr6mtaRz7OVUnrhmHy5Fe4k7PcaOj6N7ZcGx6Dw1aaIqAJRw0bVKdJWi
GyaOy6EcehYozQB2F6J/W3TsgPDu4LomYS6OY7NDfDfTctGt4GXOh+I8B1/P5VYrXfxonbreVdJw
FbpSsUNBPlNehAage2QbxasikQmiavYjbztPy/5/ZgBCtHE3KXWc4A+x9o+WqUaZfoPvfUwocP9Y
eI9/tNMK5XXdgDvgCLz7fY/pusLPQUDOLaw9anQrI22c5yp2n7FQ4/orZgLnUrDwQYEzvJGZ46Z0
WS6GpUnp2qtBLiLYCSKsqbG8ZZI6XDjQreVY+4k9313/yKU5xfe1BdmB6lsFRSwO9ELw6mlgd7nS
xGX2W3jO33bYWH86cwEJO+OYMI0hrik9YcqjjIO+z5KNbQCINP5zXBiwxFNc0hCW8VGa/4gY6WOL
WtA+7Y9c2GPM5X6K8fWo7yUM4vxdXXOHSrz5+Px0QMq/Nx/UuxPPLJ6bOlBu/1Uj5wp/m82SispW
MREgpxP3z+v5SWD9kwzizuJqnu9c1hPl8jJ+IQvLMjeYMyGJS0DqgQ/GIL5iYdLN7g0O4HFhXvig
n5HmgfYxTMTVPS8Kf0cjucD5/sTPBmhH5aty4+/bZS8fRwK/ULdE+ktDQGQdz0YbN6ZfMXR0aI7V
l6yumG/w3N0d4bX5yza5NU4DigqKEwB6MlTPGFxInOHke6HRGzhbx7XMkUuwQvIJh/VA9LT5xP10
gMrAtqAQlr19qifA3703ZKOlBiEHgW4ZjBvaMz77UgjAnXSwcfGlHOYkEfaZviMMWdnXywMtCHfW
UAY6tiyA4LBgs/6upKXPDGBpAXNn0nJtn5QoSKOOvCEPyOrzbFGtcqTdqhrlep7FOiJZNER3bqiH
qrpBCQDqZBqef1mMMsm1qJbo0FmrEzT5AJTYwDvMEjr2Ks58EBe3CiAcrWpobCIxNSBl3eSyhWLa
WPYAP7cNKAhvgmj6p+oui+cN7BTmv//8pswjYluBAv5zs8rXIzR/+joG8T5ncujX5gi4PE+aWdE7
xnK7rga/wB5/bqw99GtOrgTi0tX1RMvlAKfdTSb6ZpS6TTX2PSEwKrSCxDtdA8UBZVhkvJSKvnAB
OM/cak/vX7jvONqFjwpvCM8Lkg9F/Wj3s5BgD5CO0bMc5rckBmKqF4AUdZ88doB4rrXGmJNYd8nR
vhLj72xEysFtE4U5GqpvKzlhVu5u+2MNCMXZ3Y+0Y2Z9tW6srXAw+5OwvFlAtd+TNBT1m5aSDA8P
C6Ge5aBoyQPlyd3Y4tFZkQLh4T2MJGBtKNDs7Kg+XMkXQA5tWs71UypHqqI2rRWwcJfqhVr8G+RY
Dl8pysv6Mncc/JfZZ7jB+YsVqwIIJ8Y1RkryNvgsg22FDxsg2tf9qYixZIQWFSdUSNdY2v8p3OvW
XaXonaakzrEx5T/gkLST50ed02kWQlsxtMcaTQ9wZsn+657LgrsAqPlr5fjQTm1B0g3qWw/hEy/x
Cz30+sXmWgQ5fSb05FoN7JSfPOwpOtbO9+aTnLfkpVkJugOHmlswiEdXsX1ECwICmlIH3o5Z7Vaw
VEeqb7KIKiyKRwRMqZ06TzZxjczXwLdcLYEsQpAC2J8GizM3KuLGXhvsVAaxkj8wV9xJ6A+mQ7vE
Mkmtyic4XCddd/PCzfeGyl6T3tgZcE0hpdzq1PjqhGRs8cJWrPl235ghZef24jOSz7Obw1cEeXBa
3b7wCBBczHLZzMuuNhhC7OTHCJrXrFBf9+m4Ub4zkTjpS7yRye0c+G3MvZ84q4uClvis0v6pQm++
mBbttcbVN/eEBzyP0AdTN7wKN9bv/6QV/3ggJEPVWVmVkiM5cDc1VCuST3/WxyQ2dwTn0nCKeCbo
Bcgj3rxS7LzLZi3IPr33GquzZy/g5Q2jIAJ+Sm2DcT4RqxaKhpk0IJZpSkRu/jkJNNjve6/inh1r
DwVVpiA9QurwVI9kWbsNbjWX/RQJ5Pp+kBPdCj20GvjWp8JtFGKJfAqv8YJVpUvoFtnfCz8naP+0
zmTRJiPw21FXO1ygr1DdWuWjvkq8MissNhdDvDYMGzKI5eygjXbGOCnH+9OHu6Ko6g+KeTxMOUu3
gUAfllng7YrbflBNDd2qs0n4J0z97sw1Avz10yMWGQQQqmPO/BURY1beXDyag+n2xrd7b3LPD6aN
EStkgHLafL5QPZilkDihqdc4qEGupL63bBKGHteevCf6sc1hW5IG9ZGzrsYFY6Z3jboxFFGm6tDq
uScnGK4GZYXAgmxe4eeZHcZuWTu/AkmjfOVBbPqvIroWs4YkspTKRHVIPRvyP/50Qu38LBT3BRM2
lq99ZwJSOfpikuveDP2dOOx8PMZz4DY0HBpANhLt2AGcWPlM8/5TyZnXVkG74caev50Pvcrte44J
PxCoDP0F+SPhgr0NZdq1GAB08vZZ9/HDWtSobJunxZAhDR4WzjDuuD1y1jNsIoQdrK3Xs13IODjV
XIJCuegvTSp7V6G9qDcLTSgGhp2dc09rRKS9013KJETocGCPH97zlHbP0rOXWJKVvIV4m83XWHKz
+bXyCUhTIKbGzn8oseA73RnBNv6nNkx28ZCdiKgMA4DErMSde7IHYNTpfw79yS2WlVAXnl+M+oVU
OTSLkFO6k3WQ9DTAbRS7VSXVn20YpmJvk4Qs4fF9fUaunR5TSbPUiNaqGWhKJKHZQieVGMu65A1X
rnmZh3Jixjh+H+ZByBDhr+m5ueBB01tJqg5XBc6Gh6WdtgEcnQOqcM4/0lSBSIvCoKlVF2M/54Ns
NWPIvEbsBhdTq6dWJh2IgTyxHemDsPox3pu9qZb0nZM+/3yG5cSRAFJHUuUtwHOuS93W1H1e5ln/
RAzQ2Fpcm7MX+Phw5KLow9XXiCFSTDlPvqF1rYgFI1IjsKd1MXt0+GAvMpmh5m0SJbziFB5MIbB+
jte0Mp8cv5y5VCQDkKehF7aVeyhm0wWJb7JPwQoXncLJgkbafaoldOJwp9Uz9KoOpj+zm0aEMCmH
bILLCKi4GsM+2TbwGQE1Mbg7sNYQszZWifnJea2S5pnW2yBIn2O/o92fF9kE+zvwi/lba23gwjmE
/ckDj98VBbdpItqCiR72tQ5IEA60rqz0fgJ9YiqXq+WizuTfwaGNlYAmZ666kcjFvsdXzhgyoG9D
5bklXu7XQjr+Ma6xHz3UhyNACd8fgbT9eGA2tcfeu8NA9ZAoOwexmEdwQjslprt4V6pcShiyF5JD
mUvTtwLKwnidHiqURoUFWK74WOTxHnTEXS/ksPLl/vhzI5l/pHOGaUyZo7rJRhluAXixwERlBK1N
94CsiDZz+ZMkwLia10W/S3eEKvRGFhgBPlyDUv/2SZGOV0kb+FgDv2AA6HgHl8d8mHVjlmn7EXC0
QwG6F9o9YYU6k2kELqqzcLIyRpUpODi0ipCWcb3NiCJbLWPr/qw3GGTVYGotoCspHrsMKHIhaCJm
txFosTM1LInR1xc/AIZEdsuTMa8riB4eriyFj4PKTr7Wo1hvQ85JENYrty3NjJpQPe3uHosX3n51
FZY27HjT2RLKPokvqkEu/PX3BSw8yN+LD8lfP5ewJOc2Qkoxx91ZrJkSCG0H9ltIV6z/quxKXPxc
HUGaBN2Vu7z4+7ODlPGrKP4k+dzx/RZrKkEcovsM0PIuQaKre+VascGVx4h7QDe1fRSpr6yq6xIo
OVvmds2hdrOMF1H0RP/PjK27A6KYw2IEA4JaBjiMqu69ycGI35dpt4zr0+fLHouTU0lVs4fejzuc
AWrY6hAkjyoC8QJbiIppt/HpacoztAflbJzygOyQTZ/sL9uLFNvtdRzIwkiTGgN+KKqYZo+IAsnk
qQyxxaROmzdtZFnQxHTxbFLU+bab/y7b/lHHfwVaG9r3Plbs4D5BSMmgS1/aGL8f+QBNaBBS0oRR
m433GgRLTM3OrZseslA9/drtrDgut+a02Rw7yqkzqIFCCbmL8xq7vto4kQaesqwp2YZYnXgw892H
E+DRy+xLLkgz2mgAp+Z95WETZsUz0gTDft8kPKOXDREnIJCTW7GGof6Co6DaukDB33aSANMShPqZ
NRj72rRv6CiadFvAn0O+TvqFGbJpYRq6v824RyXoKG7/f473j8OgWZzGqGf+bSwwQf1wx+PYk/D1
fqdUqszHXemZ3HnOM5bvAAVG25nk9e1jTv7n7yIcHoYr4cdmXkLhJ08Azj7ga1Ghln9qgEv0s21w
Cr4dM1nqvzkTJ0rF5arUOgboJX+PIIMbG96seqrNSVImmyR44Wv2OG0QXxkqGMKTepHUdHQs4xWh
hP1VU5Anc7DhBn24mZj+U+iW2iu4KtaO79M+hRKHTajjUbSXOeIKsg+04ZOgkAzHJuUhnXxZBNzE
/kQgfkng5/0F53CqsqoFflck39/toSfEA1Fz6ciQQ9Q8CCQTqN94c0K2tAXdSo8n5L3NM0zLW6fU
imdsSA07v89FjKoRyOn9wlHRhpsicpuT9ryZbxqAeTbVkov8pIFpHUrcGgjxYmHf8/S4hnySGrEn
1JhaJ7ySWnPbs7i5Wst1uZFFhjJAflyymoIEoe50eMYzVC1DRR+jaWBfod6NqnBpKhzMAxYuFA9F
IOoGi6ph8QPDISyh/NUJmVQEUdHdhGb/PVA+55TnLuLOwDyXJc/8SPdtXfWgGN+7/rrmH8X+EUFt
eBlkwl5RUds+5EsyiTJqb/HkBXna8GxjclFvQctEZEKYfbveQRr3fmEXpCWbErerFpDpsA+VtHQR
ArwBJzq0zEpx2lqkqmTJiPkLR/QOu+D/gupJtsHfq7xau0U+GvxHq4jHRb5xdmbX6MdSi4yF2GeL
hnIIBbhv86vaZcqTik8PpUoqr3zKJZHJ7osT0ntBEt8fAK/6GoyGFphNkNndC7HHtwor0nO6T2/Y
fZUDpZbUo0devJ8y+6rcCE+ohwwnoLN0blJUygcgp4E1zbEb3lWfc87TpKV1bza/pIKHXrNAEDR+
vuef+jgTSb03OUxFssZm49MdCfFb9CINMPisrpZwe55alC29fzZfTVW8cqRuiYz+m2xW+sAB74WX
ykWJK5Vqh/88IT9O+fMASyb3Sk2J/7Xf6kigxgm8mSCy8ZUG+lej1UBDNCETgQcxOzCiFb64wnT5
6iRqxeut+mnejO+iyuQuWtUftYn8+CXTAEybpiCZ9+oNgY3Kh99s93sA+BH/aoj2CQ8+wkBjBAmp
cPbyUjSjmjFJ52a0P7GVq5tpjHsciI5EcqowKz9ILSulVKvUQtdRo+gDpkdagzrDRNoQXzX06iC0
VZmMYL9XzQrZApJ3sWhz4xLrhE0Tw0f0OsiU6gPKffar/KGP5l5TjN3E6LA09qzRPDBa1pGpgV9f
nMQwKCwqUScTQU6TkSJVGaIjN0XJR+MfJKS86aNKzRTxZPWBBDWrQhhEHMkSJbZLJmNdjOFBJvU9
IP2yr095U1QEjv6sfcw5vtPjXGAM0JfxqabnheAW4rEMvIY+Ne6zlgIpJzbrpDmVTdI37NT5CzLw
wiP0v/MAILjiqge1/KctsvQrk3GppNi9R+/roY0qxMdo7O4NuLI3gouy8wghnUkROa7EXajqEMLP
isMBrAOV9zO9dqm79gP2IyR0oyAdxb3DS/ykwhd7BhKxft+sjBK8gAEqiaPeekrGaeloxvQidL1D
rskJJZR40ymXxuFY1Sb+n2X9biZv9fLnLGBAIblknVLnbrtMrnP8UGTm9tV5mjwshvOC2ApdHsSb
vHmNG0W4eZfl0RWjPLGWklCGmMnV9k+ZpYbp1jqW3YcHrIwI65ZFrsD0sDyujaDzv+5ntEfvWd8t
HcBf4AmYhNCRRJ7MbDU4OXbHS/jhWh6W0upF3YY+HzVaMBerNTt3HTO4TBQsQ24OImRUx7tUKJSz
i9mSju1jqDKMHsFQH2JzN9+2Fs1NNXAPmPdpSoB2AVlw7cAPnuk8gGH/czOaj15obd5iTqABXIRB
CfqX4b4TjXAj02Kh+uOl+98DXQcsfCxsQmUdtELI/2IMoSTbWlxUZb7G26dINCe6PtNtVZEG4d00
PYOU2IsT2HHmpYgwpxCAHL37mQ+WrKyWgBFhctC+VQ5itSNltv9I8lChHSxGUj+48DThWxQrbwN7
jbNuRt+dNbPBcicZ31u8dq8b/VmmNGgZ9daTtCC9e2CbbBmbBX3TFvC6hgd2C6Vg0sjLU7zk5IzK
tWBaZ5JswOG/8XL+Nt2Cdn2+CV0ZcPfQyn6Vrs0bY5HconQhAnlpNNtxiNfuwCE4vfSAzBLxrRnm
EcRDq6okBQsZi3RMbKVsFAEBjANC3ToLc79+mzCTzhCMXZi32wOhfJsUMrDYcJ3sTohY6cAIm8EV
sK1mFNLDxhfg2cO6xkolsyxMN61v3+sfD6MEOoL7lPOaiScElAnyyGPwMv8mFF8lqxJDbIqhyvoR
WWMwj4wVkQ9/kG3170WstN63pKCE5k8V+oX1dbzr5jdnBA7yaBDg4KsTlnkyDI+fAllovVyAwPul
SJ3/YziBEcz0TuOJZjM++3864zNSBlrIyyCHdy4HLp18we6AmWtU3YHIiYNztkkbxhNdtnDuZ32I
SacRFOtuheBEWd9txrk216Rg3VYoJ0hGRyVJV5yqYL7HlvijnHaGjPG90AEUu5nkRyjGPJRL2T3H
gAx/dQM/Diuw8/Wa4/HKvsOyM/JbNohNqtvEqvcv1sirb5RDq61nEnzIuSchrgvodILkh/MTamWZ
zWBrwf+b5DW1CSO7lKtvLC7euQxDg1E5V5uc9z+1Dbs9MItxYgAui8c0Vdo9Zo5OaZosIw1xBpkw
1T8/qZEXh1eM8b1pq/LA0XdSAJQRBZmGsb+iq5uxEzXq1/eIFY4ZrCJyyiOE4scFDu0nex+6LAS2
iHlo0WJwidujsLZ3r4PEAjZwXaU5BPZA/wvFNW6qI4btPtjkYGsj5nDgP+jKUcOjTUl89TqaNbbe
9Q0LAqiJQyFBwMHa/5UxIr1eLbVEBbfLdxNDuOWQAkfj/szesMq++6qkqrxsXf81n0uK6Xaqddeu
RcCkZdYE5nhKhgTIrLL7zxTwMO8M6ohDidNIUWRNOg/DdAxd478YXsdhrND+7Xy+BBILiZlNIv7E
hY+HCcX+c4ncw7MdPNm/rZS43u9ZJlScn5YjntNp7hWSSs7cKPPxGr4DZmZoDgtYVYg02Ijq/O2u
lVQ4b7m04hWCgLFZBox9Kof0RQr7JpR9fSpTNteQN4jTh9BF16DADV3hm4MvrKNSMyUsI+peuYBA
kH/NdzHIH92Cfy27BUUQfIYX+PmetsvL5TcRaOyioRcsADDtxXsSwKaEA75SSSrf9RPSQRuMtB59
LHdRPd0mo7+9p6X1fNA59FJJU3Z0wpuMaSUJ5SIGEsVGVVULM2PxMGFKVfte1AM3NZ9Ok+n57zZl
x+ZmbYwbeBQnN1Ofm/4JQMzBhEinFy8kvgJNd6sy8BjLTWUzKXzmB6f1cXBtFyPFk5u/qjkRCjlj
L05DRl6FtvaaNTDuRNoIv8QN8TxzVTmFsXjI4LuGdwSHrGSulfmTxufUqothPcHcbzKH8e1KO1JC
GFME0Ydr/QouQedOy6MbmxRJtmWx4n5N++yYN7tV+TA2KP8MOFSVc1kdOe8PNfm77Al2UHRafk+v
wESXYmd3EzVZK4OiGauUROZ3OKBJg0MdtvR5DljnA8iFN1w7mx6UWRbeK9aydkj+me+0IXG0JlIE
jQuzrtF5NMLx7AtCqmfL81dF82NIQEM75CXp5e1EhoBT9tkfddEVAGg1upm0xgoMEtXXmYtswufI
cndKu2Esh2iifYoPZsCaIA/EVky3x1RQLPVRayg8z3MfrIP09cqYWsazV1dyhmpb9giJGI5suWdz
Mh34jugJ/HdlICs5CpPbP36+HkCq2oY3Q7EKwQOitDDuG+AfxsYOLtkbatKOe9IQ7Jt4rP5EU3Pg
yWdCz9GgweJ0F6ZMjtKQJNjkaNSBsTwf9er/XDO7Nnq8rgTLdUaxjHm9nKksCU8beRgZECSxumMy
HNTUJJvrfT3tbcORqLhC4zg7g2riLbEq8kLbL7ddsK/iOqGRvPlQ02wINrnyNIY63Wk55CUuC5mh
qTUE7McEBIeA7tq9977m/oEDo1PjP0wxmiUdg6VCnxD6+8TW8KQwju54VQzFWVyIoloqnyvbwTRZ
afmNhpVruI0JEmB7ar57JtZ0GBT13fY2DVRhhaAHo42LuXN47FwSmW8XM4jTIzk+nrSWQjAe6yYO
ws+qwxLf10mX3osH1gYo0hgaafiM1Z7mcUnphA9DPIy4b2uATx5Kc8kdHrFbmVH/EMA+Vc0EJeMO
gQ76yuaCpQB7QKNZULgmXQl1+eO5HEgU64yXHLCjAhVQcWAT7Y5KwR3Uwu/Qm5YZeE3G9MmGgK2t
1/ErOiYIZRRvjPGKNkIPMgDfN22VtBliIaXeMQCThW9cTYF8UrdVJhkoTfd2RFouB0BllY2cOI9Z
r8IG2FLbr08C536yDrWK09txFoSTYfFUuefv6yDbQj+bqghSx3H7+ppstMEoZcfYSfXTKz0fAoz8
F8wCZuOFAkFceI2M3CJVg7QPOxuv0Wo7w+7ht37UkyO8ueNra7xvjMJHJ0ejCDS7SNo2wfcgMA9r
O9fvNr/1sYo8+TSLQgvQHtszU7RDCUqRUZlLQvN/P5XvAzEYRuZRGYexOZXvwOSELX+JFZcF3ynE
s+bKaK91uhjmm9GtoSdmPA3Cw08lOhHMC5MzHYJ/nXfpHLmcamrSsInYxgdu+1WJrqcvXezbeSSd
uOGud1L3QpQouSQpWwetkWtK1TpW08gheWSQG11+x53WA33wyuioFuMViZp8aoZhrUzp3NaNrC5f
TgB0uzFyRM/0CRBg8yOd7SbZFfNL+Tb51twO5cu/Vk2u3fLIkl28r4Cg2d46YIO4AY6zFGwFMQTl
Igjg+11IJdk25MGmTOXyQy0P2VO4H988GHdVQMATYzL+360MPgvQQs6syg6lwXyltsV4+dp8RmCX
UryTBVBJkga7QR11Yf5gukeCN96ueCQutFUUyC5T5PpJcuryY73u1NMgO5jl3yHD/toBgEzXAFV1
rkVCHWVturqDF0oRpq8KkNrfN0prm8oDMvyIOG9x53wpDwJWTDfLXQMaOScyZoptpjnM/NGVegYh
b8MuRrIpF2w1YpLSbSCbJXGCymOu/zk6eJvnQjTG/rODJA0yL70L83E0GK1aM/V8m2k9rO3J+Lzl
mQ6Zq8BoY30GkqhKxZD71fDALDE5u58qu67sfUHsMO/HtXBpwED5WrCOJwuyJtSsYHbSc1pAhrC0
ONb8/1guyKkar8cT3Z6aQMtnjZ6WH+Z1i30Jwabq3PQtFCyFV5mUQfv2o0hIkXbE0OehoXGYegl2
4qbFkbYSALboekLxJWJuW2/B7/C4Tw9DI4Dnq2lgypUBJOYRWbOjiO8veTaY8ol3K9YaO5IwQojF
cQunlKjuteocGgSG0sw2fhPdf/5wCeauPSOqXFpz4jINwbOPCTsDESsSepqnjm3rT1Mbh+xSE0zl
F/VSCIxtvvEcu0wzbDAl/Fnw4PG8ob9QTb0SOM41PLzVPYOpYF/asNkoliA8j5C0I7sTDyKgrNMv
6ej3elIn7dkH52XN5mW1DZBBZn+HkjA288lstEeRVhtNlWdZGaq+CjF8echWvMTh0QbgST5Ehe9s
+gTGooYdmX7mRYQCtvRSoPJ/Jyqte6uOjE8zLshDe+Y5EVn2mK8O/q81GBPWFskUNfJAVYyCSHMU
ABATAM/r49jnIpuYdsSYMwG3HGiR2Ic5QwylmyBcSgsr90e4ObgBYSfaE1WZgbcy6qAYrw1bk1XN
TdIOiy3Od1hcUMEO05sX0/CsNyDxSxddFA5rnEx4I+4EdIXhIQTWv/W0FxyFEbxZq+hnkVBU8c2k
RBgpdFQGGu9l4em+cd2Vfu5VfvuWixvmlTlMZJMwS/FxF0VQYACgC8k19o3LIVW28776PAjPxC+9
PkqLqlsAAbN6G7rAGAsnk0AA7AOnTHGWyvctDWHJexKNOwvmz40d/+61StjjzVSeEMzbtCDp0WW0
jQWcnoNK+UoSf/fn8Idwemr/vImd0LEzA+ecDzj/x/kr2FqlleEgUoyRMqlpMblSPUP396orJRC2
hGhdyUPVrUukFfi0S1wsklMZqXcsYck1ox8CRQbr29CapBkYRNSzwqbfVT45D+0244kgDhyOYOUs
Oxca6aO+1dt78cG9HWRWDRFesV/z7vwk1fSEOApQRz5TrZ7QWYqqOLKRGp3iqva8zskORCTFNRym
+JyrlHYjQzwk+gSiKV6qo7nSoSUi2aA0t2HFNfmnTcFFNS1FHwGYTRXNM56vxK+G5gsIRNBtn6oR
olCN/Fb3RsUkRs7DqA7ekNwYT8fF6V3LM8IWASFigbIG03em+tylxZOffvptxxS7ddvCgIpgCNTB
bc4SZv33dUSnijlmUBjvotwW8/cVHJMp+vBlqGr9UT6IDPI/OIUQ1eLemsqN6z13dm0Guca3Dw7M
wRe5o4E+BVXoeIWFH+Bse41xIDbDuW2g+0Rq96eFX7Ni0/FILoJwpAAjsXYKdmUdzmvl/HE+g2JG
qYPk6V6IRrSKeEy0IKLQezia22i28XuvBFfUSjhyCoI5ymLs1W0xc2Kg8FdciTq8yWXYvlyChZRM
V1dJIKPg7uhzXTmSkiZFm367jPRwbjEsJ5w0eJmIhqZsXmKpOwvXxX/lTIT1bUKkWrYvbDmK5GLa
HOOfOGG/85eEDMdAQ4eWqkxhrQAOjBV6ezKGZy6yraSduw4GQU3JDRVI+Q14XfkyXNzKoXpu68EX
lmJ7gqSVihG8DK2ldROjYrFdvEe2BGUVMaqqxP7E3N2fyaIDgcpjK7WCQahAgTOkGTJwpMeCq4qV
mmENkA/LY2UkT5zqvsvxd44Q2hpoBI4OLh57uqiVyBRYLHS09fycEfanxmx6SOpO6AOORRHkhoIZ
BoZAC6+kgajMg69zR+DMdnXDrFlpFjaLbIEWjTD65YmoYX9be48/ZJqyoop7u2+1oncfwQ64uWo9
1VX1r+IRuKLtWkwmC/K2TjmA11looacHK0brciNkMJWC0SGmAQjXcHWI1nNEPGzqp/KAwZ12ocaj
tNRHx9i8/rh20EKhqrBO8sR30xn36aAYvztIHOvXilbS2UF6iR3GPI8lbH2qmNgFCD/iJ/zVaJML
MUYnc9oS6IDmRXw9Gt6gQkhzrCdWeC6HuWY1J/M9Jbg0qaYqTxzwV2csw2kmXDHJgTVAO8lxYYYa
u27sfQ1fuhCuY171dVDMp/Kh6Ni8EXN//naforqQEBS0SOMsZeYxgcoRyO2PpCatrm3GTywOxnWu
fX/jwvTR3rXnbtYy4o43aL0w/cqk8G3ecJO+A7QJYmRilEIXy+ub+I1Ahlq1QX1jAAat/cnQ6QBc
B1f7l3amZ4nBpH/AsgZx6b/elR0RzMScXV3mZ2UzdaRBW5btzUa+zz7vOixnXcS7LvD3hVIvmJpW
uoMqHK3qBkR+V0nBqmNP1TdPPPAKoy0wKMbKvy9ECv7+0EMYw+Rs0lFWTrSlKIYRiF56m4HuGVBN
ZtdwX97JiY6DB7Qh1f7NO0DOO66BsOXP8WiLsX8K+ho1kMXm/NSuKKuJiXdtRI1IqlRw+Jc0dJli
PvvkIDRJ2naOeQgjDe7U5ly5YL7cQc5SRxig9kGZQSDJf9QDhSev3ZYxLXq9yElXIMa6cPHFtuMV
vYBWN9QRo4ro6mZYhmw6SNodevtdGEJz4wakjFIrqTV+sBo3JKFi5Ab73gW8pzAwoPQpRt3W69Et
X0XPmI2iF8Y/uZA4p5i3TQiegYlm85wR3dgWPRna+RpPvscWQMTA67jIDbFRTpK0kFnnmkGiNMe2
QxjcMFolOQ8ggN5fAWSCvt2hspLTJM+caG+EGk5EwJ3m8cnH9/9Mys0acivBsCMVpQDCoZSU61wY
68mqWBJSNtjLdpbibbhfbGWX8vdKzdXL77cvpKIKNmlc4yxeF9p7ftwFM9gXQOIRGSM3RD0ckKQ9
xzNIjxAEYhuZLjdPmkEnWGJWnusGUSVcLCMw7p788muUOn6CrxJujmQdZS1oFJwvd8FbB4nXuJZV
9tWnfI795fw8I4QRjFpGGg9gFEnVt4lGYQH8S8F8qzXf8nrvUJVqKYBbj24tHLFwEPR54Y8m4pAl
nbmnO2dwHvnrW/NbgsnCbsy6ZScmkIkGefU58Yl99gI0Sbwj4OtpXZlMiQAC33QjkUNnlwgaB1dV
xwafHtKJzwJmzSNzIQra70sQJ60QAFbNSJPUDuZoaFvAnB+jz68iVCcKSg0k0Bd1HQ92qnBX+X0X
ZVB5SUIwtr/isoeRhFT7Ht5/E6PqlNoTxjod1cbh1biHrg6wYvkZjWIax04u5T92Y4cq6Mx4nX4z
Z3f9ESJYBytu4SLcLAfn0YFkHgwRE4UxrAAp8PLsFa/Z9hYkq0yN59Y9RBadOxIkDZqUzR2rlfy7
KnFNyA7qxZvbjVQbTl+ZM+AXMRMqzheOHXBHGY4qqAO2try7kUTHH7D70R3ZT4F5mIhlcrPAWi7k
PNSXhIYQx3dQKiqfl4vjLdmbFsW5nTuXrtgy2ld0H9VCtO6S71OMi/HCFM1nuTIEUdhLKen2EQ1Y
zNFV9gXsQgaC56v5auv3SsOZTweYfRaxr7dVMz5GIMrWWxq3AQlNM9/7Re8sIvty2wRr6pgQKu9c
SCUiWxVIyoqlCihxntkkyWH9l02lDM7fYZaaBZMJrlXxZGU/X1i683W06tyuZAo1lqv0f8yJTAfd
tDidyccasZg651LZnhKO84/ygiGoudH5oM+uzvZtfFJm04GeLHuI48aqlj/SYLGPF/aNgnCSZx+N
+ZJQWPv8hPea9iQf6eCBqgLh1k1PBetEIzAQKbmuL919YBKLG+PynJpS71A3xHE599VoPdjlvkNZ
oA0OaK7Br1xXVaWScWIWFUBo04LzI6bfMP/bP68u8ytYScbXFyf3n6rTGTUEJIsLO/IhHi2IluOn
X2jUxcjR7l4kC5+wyigvIvzZMA28gmbUr/jbaShSf8AhHbPO+qU5FTxLfgB7l47bn18cU1Trv1Oe
CF6LjTIz/XBV6VUyA5/0y7re9SYo/efkRAv/ASB15rd805ByJ4jWD4YlyZSij7BQIRw5kZBjVU81
2QyciskT7RWSG0jPhCyWNMKJDAN+wUt1YU1ib/DIvJT+dkRffMekEevaPTXQ6KuXoDGQhsrQKdzj
tw4YXUxxws/PnL0Frf7HZs6fLpCrjmfna12uxHxMD/Wt/OIt5VIb8o5kU44HbLkEf14ktmHRBB/x
lKXZW0AbB5EUPo5OUWLphr3VXa9qlVcpihT8RpD2g/Vdxf1O2LuxdLndyvVI56tAVTMZcCPsSXZO
UGPsLBfcglJGE4uzBCbc6Mj1eXehM4X7ecpaqGVsFSmfQUVNtq2ZIbtnJhnhTi7wlvYJ4QBTKkg9
pUUO8qScabbAEa8tW2w7lTraL6VJsSyXFvHl/vj4D4j5pKB4rAcFuHwu8cvUnuZ6IBgJUbOU2snC
FVGvztonprf8mgO8FuGze+IyXH+VoFy6LAme0JEUa9WqMAyQUe/TGNrIayQlpdLcElXmnKSG7tiX
isGw3/Lz2bVc5hJHamrgjbl7QEnZ0V26+NNDHPkT/VgmGyZi3vkH5/k0x//vKUQyYcToBFE/3yhM
VZ8vEHsOh7N/ZYw0DzFFVUDqK9h+5EAPhxr/kf3TyUTnHZmCjFZV7lFJzqjIXu8MdBLvS0+rZpfi
650phtBzmUhaduRFYfQ2WGwFmFWNlzb+ubvoM9FfzqBBRULIxuFu4uIvkit90/9Wyk+HoX4CTehH
4Te/Ow6JNWAt1ASA1xxpViKEl8TBd8206NJXMe8sJ6rT+Q9q8mx0AOBqHwYqFCIwsGZW0GzoAfBm
HrmMp7AO6lb/9aFowoYtE/hC1pGiILxesYV/pXy9OF/lERUxO4T1MtTdeVpCgAt9SBjdhhJ4t7H1
IGas50Cln4LjFJe9rNWIS06kUXE6nZMsvF9ndcEP4mKw2tBBldhpmrZ8PBLtAalylfV5Dbx8bcDx
mwdngH28yIi5rDk7HPdkG0qSZU5vTPOI2vu1LJAuyKFpLCEYVZqC6q+8DliehvMBN4ohckmFzSov
mZ0nA+CeTeOBROOH8JZ2N8RqXMGMci+lJRGZKhMOovtyQB4O/g3qgwLWw13kOEcjWchQh3nOd+sM
YGKCddVG4gHYuJz8wbrZn+unm7gPtz6IB9rNRxIBkI+gaCk1+RQQ2UqKLhnyiBzQUONrq8yv+E9y
TLtkCSYEKePgMwlO2S2U8QVhnhBH3C7D4+r5BjMqK5KTzP12XWpXjmH68Sua4JNeCXUDLZ5k6K05
aVd6hM742oW2Ed4oi/aBWBEBoLqd+9hblFQ9COvhXn+c4cIDgfDwaUq+q25P6j+H8b07XMeprffV
Bi3C+giNhRZvK8IwIeYqfpvKnqOY4uBvadLNLwyczW5c+W5Iu5S8WDEJjiC0S5mPKJ9Rf6tYQALC
V/7RVkJOc9iQd/IXquYE+kYXJ1Cz27xtjuHJ/OHCf3M1lqg3Kf42iJZMPBJyq/6T4kJRkFCg6TGm
tthiAJnEdOPsZGoPKhB6iAVaDVLTnTm2nCdKfmUa+q+reZQVgyijzXd0FKZsOycOLUCp5WDddD1w
iBH3btNYDKU/RLNqEfdZBocUiOMrCpruQZEBGsD+ohv15oGCywvB9OGFljePukSvS2C+bYbnrlPM
yrdYge83KQzp8N8j/0RjyGfYqP9QTRU9ZrZUIg0uGq1fEVhO/RWPW60CE+07ZmheEAfbK5eRyhWD
XwGPzuMISP1ExC/C1KphP+EurH/NoB3uYLbUo2MthBdiatHZxuui2KGwwxsmK6SY49hW80FdcnaZ
jhBjoQtT+J9iaPSf4NyEFEsiZ1ImkW8g7X1zBqEb1dSc5rRUZg9Jde4Ljk9sDqyYQq9+8Z8M/9lH
q7eDvvk/8NtpIzP2dv+X3HtCAvooIdZLc8Vv/54Q+EQ/0gFsid+Oa9FU2LqzlyUMCZGJHvE+GXiT
ocRwxYAqtlNq2DqoduEY0fUm7WnIYrJKxIIQKf8DmUTngga/4D/8m9xGAJniCwX686cOF+ADTIMC
+QjlCURFOGd/N4kQu/TbV9MefpZRiDqE/w/gvVre2KypNtNGtOL7SIXUqmFkHxONcAj9xHUt+ixt
COcPKVqy66pRleVYhxTPNjtqWO2UzCB9ZDzFU73e4S3F9dyFzJaOu7UXyHqIQbiVSyGhFS/PNZS8
b6B6vR6DgJwbOjTZM2eOSBEWXaraY3FgubX0bMHHLhdH9P244t8SRL8yldiCOBttnCQAWlTck3tj
jJPuR72q87uaIeZiHwlpgHgfYHca3VFU8KGyCQojVIJdPehdiH6VQVN2FGZV94W4fPWMOP06oPVq
6DPwdznI0U1b+4CiCJOkKKT3vEtv2y7eea3asgILXFt0+MPI/XI4XzgLlh6Y2bzlGty3/gQ1GyQ1
zyZisIHKXRSxrguSKhxlr41VDJXTbjbbRkT9kqi+gguSsaC0EB2U8cJ7ViVgYar9UV+5Q+cEToXe
uCFAgw5ZgUyd4P9H9dmxazFpTQcwODKrZCj+FX9xe2IVy7lhhF9yOe0Z52zV6YGZsz0W95RWqShr
b3MUBSkJ5uGZZdRPcA3nt7ND3qiy50kzZn1xE4uqODPxMZq3PWu47WRiD8Jx4zWIboWrkcSw7EVS
y7Z+kwLsrb6NSugV0sLqBMYzK+MATu6o/o4Ze1/cWe6ON6Hx+D8HuWXO0ksO0s3hOZsBJeWsnW1X
/pFkvbISV5yy9kBDTyWp6PqrrwLMFa0TOVq0rSiS+3OOTsuATm+vRPqqi0ZBm3quaf61WJFIk6cL
GD2pbXU8+iMYmQ/Y4fpKEXmEYB+8koT+i74g4FqL5tl9xnjaSguncbBcYEGku5axHOVo9PCCBLsz
zLl3kADB5xpTXc0ilFUUdXQB4ww/jPpzPpeBVQe0iAgeEQcdlFBXA8ClZ7EMFLd+hFcCN8fw3846
MUKCW8flxg0akB5NXQCfFuGP/y+NIs1j6Lxed3Q4AQoEvyPws53z0JHhZcN/VDVhp9YWiX+3hnuq
ElHq98xplnyFNl5gaXIdAV26yC8+QlxsbWb7mZZl0hZtuLpOAj+EIUhxfbAty3M7QgzHRMm3UOJS
W6qTFGVVNeYGP9hnb+YPfMQ9EchZrHC0g2T9YdsBNSQt8uGPLIeoJChHtHkBbxeCyP6nybA6RgwX
5Af9bXLj7oc64m18aPylI0h/y15h23Hmr0WTLqNJ9sZH175jScAEPsmrkjzPFL8tFfgNZ85XI4Rd
/8b68r4Mn2T7SOMb68tOdu32zd8RNkLbsVhzNrdsIdz3LlUXDP618nCClmiFp0KsOU5rcLOULIJK
JoaOK58i983K2+tksFX4MJ8J1t24bh5DJTKZX0sFPzHF29vTpQZSBGPSXxtRIip4OK3itlmkc1Gu
eHb3+Rkb3KJM8QW8MnLgoFWbfzUDDA7G1sH0v36AHqxoUIAKt1UpxXUasAUxWycWeDUoSS04Wo5Z
z8TH9ST/zVA6gtWua/lpjJC33UkIsyPjRBg1hmCx5eB3Hn5xPbu7GTiwhyFl7o4nqMAfIIZGPerx
zUnC4qeV1Zjupyskf2Q1OniMwCXppFCHFZ9V6oaweuE+7LFT1s1pHhaG0mDk5G8MkR5ANR0sXm5V
NFXJyH4gx/xk0/v2z4e5OjNbdxsxHIkbq+d8kMLoUUSfWdJfR0G+r16ME5pU0P4rIprTI0kWnDvF
tp6WJulnnPgszhdDAAhJrLQPbsxY7F1jKaiqSiNGsZum82j2xxxNRRGz9EM5pBX2TiRvdFmOkPLj
b7W9oLlSXpZfiFeNGbW8cmzqZM4SjowxvnUJJDYAXrMUx11nWWhr4QB6UEYaaXbfAFuODOf1Kptn
Yrv9VdLxSupEdrmxyFTxuZAXW6exz+1dx/4bRwjupzyNjIEXab9zD3Kdq3NipsZL8DcGGvvOfwpq
CrjnUCpOdr43y8wrzsCMvWAx2H1vCuDsE5H8x0LWh+fOBFyYwG5JuKMjVME+qRU0YFnXdg11KqB0
JS8QFhfEwf8bco3Ix+tbGUHBALiQmcIaWGaCM7UEEGh8f0O2cp7CEHpGZbeeq68/8uFrbzJO0zhi
QEwjoEjUoDqFboZYftizf3vcwo4WoE+TvV7nGEn5sGQHet4LbNYN070RsWH93plTIbo04UoUbWBM
bG6h3RNCgBW4+yIFC3o2CEe6CvkSOCSzu+VqUYBFfRE008uTOkUNGkMwPIrHL4SUahfDknGXQJ1a
2HFZFzFTrGa2mwsXUxfhYmIibrYnjEwcI4TQV8hPDRPQPLEZAFoFuDhTn/DXYesqV4nq6cANqEcb
i52Oo1199HVl5bYAzlcFiF+QHJTdkeBChs3sfadnJq+kVQF4dB3Qd2i18+wAtwRm5soFs5N6xspq
XGMz4xKG93YhluV5OtSxLLSf6abmYvbWRZtD3Ckjiwy1kVfNzvUbSsUddJtUxhl54zR8o65vG8ff
LDsCL5PZib2N1upVgcYENYr1zCIS5QJpl3R39iy6kTD6Mj/ds8RjwuLmUDbHctcdNVq9NL/2FvZc
V0lzM1gO9RMEyLd7dkURfrWm/mhW+E/30q+7MhGwj53mQme09fST0H6ev4+MiRyUIPE5eDU7PGsg
GNZwPhl88+4Mnn0gozZgj/vSNCp1BHi5C/pjPwZhMNC4ZAsW2JhG0FKMWZXs4QrPOIdgrP+TWDj2
RUjbyaYSXi0S/TXnGewSnrfndyGsKJhvKKLoHy0X3WYKhKZUEFzTgi4BbTwzKiabelAzNj76i9vm
KdTUnO99+pJusKLJwBvs6jZDiDYhQjedJ9+q1n69s9gNTYYsKm5VbtnWn59zs3vxSk0akguqJ2B/
VGS/+HXtVZHfhwR/WbdSivaSu0dm9dHtQwxQ0rrDAel2HbfHhprFFnkJpEkSElNWUqU9hjfg6tJu
MEBjZfsIEGXJ1pII+l7g+bPiyFadlP8VURohtx5gMsaINuEk0KFHaeUDmZ42eqODaxkbtc+rUGVr
b64r6jOhIce1EpBdLXZrZ8/+z7WatLXAYIQNnGIw59JvtBbr4HfVvCOucZpb8g1PWJwJaSPjRbsK
QSsvKBkk/sWubgONvqtQB6zLINN2woiTMPbagljNMqszf1QZ6RNQ/F7HD5qnKY5f7PaN4BbLICZq
Rh9s+nn31pTyMY+YOzqkWjKAFzutoUZpI+s5ubkMKwH9j3aqCKY0KXwTIf9C1+gsa6Q2zwODojs9
y0wE0t+33n0CoPWHffOZkQsDBKJqcXrytGlUmS/I6RgN5N+M31zBMIRk1kyBXOctEKnq+sdFEFdY
dwRetPQmaEBbHtvxE2hWQ0aMRiJzOsfHyf7AKGc4yrMlnjyrA2g+D5QgnG8dseEhMjQsBGH8jSdU
5hb84U36zztS7Rvod+B5TqAiQ6uHuPrI381GfzENhY3YiiRdx0pQdHvSpgzxABzJtwIPJiA1IwLt
RIjp64sDjKTAFhYlbPsCbfplxIdUKAp83K8Tv3R0fC9UVzMNkwo78LObZ1q21vhg1o4sizPPxMn7
XhVoxfs3NfUxO6JvW8EGRY86IbqRmfgYyCBuGMPYjJmpO6MIippXzQJF//WCqt1fDhR7Rgkvvvsa
BYEi3JihrdLgsNXS0nRqdrf2zfv3+RoXO0Ti42X823Ya4CmyUE5fpXnRCzN1MEhfNp8z/Qw9CZ/h
9VaS3jDBw3t38ZYSMvGkqaLmUD3qrGVOmtKq0YmtE+0GrmqhFhvhqO0Y7WedeC2ZmdeEGLtngEeJ
aQkd9mgKzxxqQYG6+Ub7ibNsvawwiKlflkB5bPPR6yeyYO26wSF8Mr4gvahHNsIaa0C+H3c1UiS0
2wGPwPZMqLXAHCFPaUcAJeUQBP3OlCF/woAV0jNaZJY3IQQMRUuCGjmUqZbiDgExuMJyt9EH4Wcy
P1BZMKAAdV7YTJnrBbPNLICp870urO0Oa/ttxS53AnwhcuVlc1QgphAz68EDI9OxrXlKCSTnoOha
mPS87RakhVkoBK85j+FHMifgwZ1/YjxMhRs86+6Ky+E4UbFqcJF+2Kft5iCmpBbtZYXmHasnhRlT
lgWb0Mvanhm3x2Ywju0vyHAZZ6rCe9lJCiEgRjNWJ6BM30DZNkfCs4fZZV3hpicem3WR5vjOnEQ8
A+CNn+wsp1Y5hsjF0GDlNZqqynHHcR47usEtxN7NS/r9U/1Fl3dyugkYMLVGlcJHRpenzp+5Qo3j
W4KXF6zkZ4PoMuqEoe1bP6/Z8qFGNK3zQfPLUnkloSv/xtNgt26k8tkGYwFjDGvRWc6A5+u9UcS5
7HeqiVoT7QbG68tkObp6z42qK2KrCTdAGG74lEP283eybOv2jqmFtcyaxLzNxlKklNm9qn4HwOF9
Tjh3OjJZInQvR5ThFVWEGSa+/DFRg4RhFjNWW6G4KA8qTTWszJlEMvQv6d2JglU4iwJvYT8N/K4q
7e+nRGXGrZkxwiplH7kygZ95lN8TFbQ82ApEpBDt5SI5OoLufWHyPDNNAMoMrQsFqiHsa9ZMepyY
Y6omZx3cRQg+IczSGWDaD+j/CqCu29JP+6B3xdlm60Lk9bnR4h64q/aByb0lcp6tYVlpa3Z64lzl
cbJv18zQwghm6uva1w4ydUT+55SF0DCuO0091pdZWt6NeNb+xFtnpSd27LhIZIIWdlp6NSaw/Wwx
w5ohvYjpY1810gWpB1ygXcZ6yxiZSFLtOnJOB4Y2Kqiizz4fH2aDThBlFznzDa3Qk/2LsfuAM6sV
5FF19G5XTqQ7oUwyzgP8KFuQtQU7tHY6l3qjEJyKYmtOA6jAQOLnMOUCKw/k191dB/vkb6W6hdBX
5a3DnzOStmMurQAylwYikgxBvbODa54qX1rT6ssHcSl4FtyHyCTpkcSmw0SarDKg/GZqmLUqOWFb
E1sZ/8rHY8x6jWB6HgXjfeKocszAhKjaYl11NsqfF3adnxOKgqySKGZYOp1KRXqve3kQGcAlZmaJ
1kSC9pvSGy0hSOjfQ34C3AAzTH1HgAwtn034oRSnMlRLHFLtQQ7PtAylVrCkFTxaauvGPIXF0W4B
4gh/1Jv77CMSHFd+dZTjek/5DDAurwfx0Anzk05tnTIAph85e4m2NT8M7vSXwq+AN0ph6Y/e6iti
veOtBcVfm3mLlvF5ftNhfzKcSrdvumJdwIuWV/0ErYh1C2kvsrIS1FlzrHk96P8vhEthT3KSPjF3
rvlpv+1aVL+CN1JHi7Bd2YCY8MlQ4YCDbbd+qC1nphuJMUWPwSEBH9phAHQxMnWONa2RQsEXtlHi
IXGT0JHJA6rYs7fEUev4LFoLCTIu1pkbMaURKKfhSduipRdmAgfnGv0va7hYLfKnukihwcIxcZkq
FMkGpvHpLU+T59AhIvP1T/pQGwnByNhnJEaSCHwkP3FY7fjiUmqSnUr7w6Yqn8lwjQQeCrZ1RJyi
l6fzmN/w00YuapwCikqgRJKyK3Av6OThBvTJ3ijTaZWI0B5Gh727grjBwktOYTcMiGSXp88//z0c
39aIEyec+Bk10CEC5rSwn7BDw+FHXG/V1oOgGPrYKS/eM/a5UV9kMTqXCCaVTVRVS6h23MKglCXC
CPv8iIMOY49jC5QR7DLpTs8JRHAbHJUNutsMi6MHTi2udgpWoj6C6E88Uhb6Tel2+/cxswQbmQ4J
GP2JpE/1D3P1owBkFa5d/lvYURxPTq2PKSraaxdK7MOMA86FbUlkWUNddjwECflK6yQiCxMrpkgF
ku2BUoY8pjf83SfEzFjwtqO80E3Qo5j6/bvRtoh/7FJ3nqBUMC5KMpGHLmNAAbKqH9slbLrXE3D1
MgocWk9CLgOKkSt1MvpAhOEqiHvEO5u/3GUjJ0r0KO2TIczfIi2FWsQ2DK4JxLdof6k/1M3oj49i
zqwjZxFlk6AxG5u9gvMU/7TG23R+iZm8N/WkA4sRmy3C+Rg8wEB8Yb3UEP42vAXaplobKtJh3lAS
SK7kk0FDmjU6rHHThg/QRGjNQHQSAsO3o9oJbRX8ulepDROj135S6LwtR+evmYGDJscMOjUrQb7v
R0om5h9TTVolfXTYq8nmneWZi/dP/620jrPm3Rvotv+F9L8H/VGcHPtn4kmHI5tnNYS+lnZpL/aa
9aWQsQKN0zbeWe+9F9usr6i/uZeujpwtTfIYnURh8wigKtsB6fkXDkfigUXV4Jn+npTB5wNSGvWV
j5Kfj/ME3WxTfwyWaanpWukL4hALDEplqyszBXSFmmYM0JySvOFwMfRzUbMziJXKsgobj1DCANOK
lWxnH7284nL5noLWmFO4uDQNzqmqfwoXaYCAOY/fNJzCV3FYdSVi+ufsvneXkdfoBo2D3z70emQH
2dugkzuCtOTJzHGpqqznv5XUZ5EuFYuPC4sJJLkGJImsjp3Sa197hQHrs3hpLWPHyPgXQaQZoeBw
72SwQ879r+tBTv3vPjn4CIMs/xlBkrNaHFEh9TWDNeQjgRkA6wLozD8uDuNfKfeY5bBCTwiWHORJ
8hTN4qS0y6JHglVPGyazE0lk/qsVwmm1UIyzDc24AZqnAyizU2/0MPMgeh6EOFwj9ZfyLwKciVb1
TN5AdIri8/p1iZMciQ7YuduwJzv5Y2gjojquF+JGrgsX8Gt5ODkR62QDmGeKRqRKpfy8+M/sMjee
+pAoo3fN70ykllK9HEuXzV6q9o/E7r5LksI+hDsiuAqzcOLIZPE9BhOBiIdcwRK2MDibjl3QaU25
s919yUuq3CiIUp8v+LTg9fFyDdpQ5MdTgSBYgTUjJOfi4+DDOOUmJ/lweqGlbaIW8LdhCxEF7/Kr
DwPV2886OIBY/VHxI7ZQoLDF51hjCmjJG2P9X1N6lNealtMTGe1Zc0xD/oky80R2WVOYAtP4GC77
WVrAHDQnKM2EYcmunb1a04ZzzrULHu8blhU8WJpyRAZBCE+50izBiIy3froMNN+8NWhX5gZoBmgF
zWyJf3E5zH+V/gZ81vJ0bsD1fT2AFXylKEg0glh7UcktohK9rWf+S6EQNqkbOGOhG+MkC1/JHeS/
R7ftvSltIhc3bw2DMqDfAT2KDHYIoUF0RiJrjx+LZH6wEt+WMzODdbt/zhLs5hq/C7ueD24eiQ/W
BQCzSD0JZPnh+wYvabvg64BI/l58TLr5UwAtT95mwX8Cguh8RxII02uuig0bDUBiAhwaZq5pv1uY
oXXLs01mXBIi3b+4KyhoGTBXz6JfQNgOCAT+nyrRjWzYdlrJo/PeUvlN5NqEBXUb8x77LWuSn463
IRIr6jWbWcURk33B3sjq++MnrHGvs7dP1DgyDxKuaFm4lqOCOkEc5lwcfhcWTxN0d7dP9vrzV0hy
DWqvKf6DDIu/42qoyCDlmXa2QlNZexNgX1r+62GQjXEjwPmcmki54KAsXxgwLPCjqg1RbDvLcKGm
ghE4VqEkfayN8iXzGMkgwa4ppJByY8bJb/R2XupV5nVguGOXMW5JiGkttJGKVgUDAUf98yhIgfGf
dV1TNRlAnbjP2tnGzdBUmdjs0vtWiLusAwbhM/yVr6rQAS32N5deGoYfknpuFYFOTgKpFx2Jv2r4
xkpEkpjhPP+ebUdMjcCal+PJSMLqvu+PQjdTAktD6whg27JRGlv/2utCMsmaiYVkag/7KPEyUuN+
IK4lbM9lTFYkxJUe5GHulqEyxc44Nlv+R9AzEtdupLfAVnc7kdGplq+9SDP+aAfUZtoiO0FaQVjt
5+/ahBZS9Zxn5dPjn9XNM7fhVOouxt9sRPkaSI0NC9Enef00Oy/ghTzx9TfeNeLlA9exLE6aGekN
kaHw5OwHRCIGl2OfiSgV5vsEJA5YVRmEZyyVIV78z44nP2upfh63qrV8CXLsKa0UFQuZSgHxopFX
xIXf4HalmweE6eMuahNBTDNjr59f5z0BiggJcsl+2xKUhGm7DkImXz/7cncUPzZzGAqxlupYqB6Q
qaDcdV1DaW07Q1dSYZKyzSVAyMt3yRyXYu7j27WKEnFyqTp86kozmaaTZmozb6ffTjv166gdCCTB
AA1u+OjPKQxFLPsWZPuQ5rF3NbTuQ7iKpFKZ6yfogwuXUUXF4eGZ1ik2OvrDuUItSF+XpCuVmop+
6v9EeEpy46yn6KWnuNRzYBv6tc/UYisvq6vrNjg/plQlBFCQlfEYhHEhquqKcibLzX+GjisBgY5u
Mr0k0I+UROOYslT5jWl4tZhev/oypUxyNszZDOt6xLv2xFZOU2zc+2IByfGRLL7grJXFkk+oAElu
GQhbxTYcKNV1tR0fp/7FfeomOxojfO2uhdmUq8/mYq5l2vdWHuQqZeGk5tcLydL2EzGH6wkeC2Ol
l3lKB2ZsEk6zAlyJgeN5LlUtj7veJ9KPE4YDCZ1bIkCaatRFbF67IuovLG2SZXC0NLMotfaCWSSG
eLM63hlgPhn8hoJTgcVIVSSRxftSC0kEibgk0tZ80XOVifSzHGKir7jwKElIEazL5gi7v+Cu9UDp
7+qjOP5HHXxwX4YgdLgBfcGjBscaiYez6PtZK7MQzY5RNzE3K8b1+4zCKktRXWaAtnUtUNeX7w80
fPZ033/6D5WarRXdXelrMhwcO6wfB4W3okLBn98nH6ahJMphIez3y0bK1p+bc4lmiGic72udRkE4
QI8s1T4KEnhJlgWW7OR3dcdq93eqMbCUb4h4Lf1eKSnM03nRnlaeSmX+SZZSNUXjNn7CcC4vkJVZ
ByKXVZvhhqqPxT5awgYBxfA7R6VYOq+vaYaBZOcYW5AbMHiKPBwTCzAJIkpIqgVVxzmWv/vLJlG6
z7gIO0CC4GbYwxaZqLmMRP7+JaSIjgD/ki2xQPn30xrZs9BZtZvkcBecXHCl+wIQBi/BFfbMmKOK
3uOs4mXKrltUSFMVqau7nHpnqUK90M6nZ8T6R8x79HXGmGVsazhAfc+M2yYuWROP/CzlNlyNwbAA
/dKoofOPOqpY9342W86AOrel/UhjUEaaO8O+KzfbvGFCsSX0XfrraRm8IdNtLp516ZGa1MjwdKjt
vBbPsMOQ1kTmhEnmvSFoNCbaiGb3G05zlun/fkH3JHvMT2X3GreMkY2SouIfzMz2uJ31Mq3HZx7Y
h1f4NOOHDaJ4tUioNvZmxah9A/oRpYRnRbulxbX6mRDS9NKo17HyowRESx88qTkwlQfrkRDDfJuT
y292FXHUOKZxXKM1SPoi2cEjE1Hzf0DIuSS1SZvw3PchKKRI8NPLbMYWulpY/bf4FBHO8zr4C3VB
jR+JZGLWgpcv3e31SJddE3CSTp8SJL5XgeayU1Uu+d8kXzdFxi73T4G2TJl5leRqgWA84xf4ld/Z
U674q63WdwMxC8b60e5wbGDGfN6o5UJ8paJYerHVFAHoEsXu8nBcPioNRog3fK2bMY78GGSu+bBj
F4MKTc4A0bO0bwT/ISHsXlsB5xsFQg7A/oGC9HxiDYoh1NzJaWg8tswKGQeGE+kFj5pDUR+DKqR7
RLVUYTmIjU2PfijJVV/sMh76JVOsZkdYjTnu0k6IxPjIB+wcLFBJ2H3k8tkrU0zi/1Q53Mu7IoJS
aNFOpH5R3+sAbyrBBkIOfW+nXpoaCS0zBaAG1SsczkFvnz5a1LnUD18lZg/7d9MA/NKLVLeMdWFd
Nd82sVA+tmfw1gf5ge91mPUwmm/gMaqaeZwroPesEdaGRNo9KHGEPnHKBC/rqcdFvizVLwaMbkYg
krhxOVlMP/DwcaSjcgYhVGF1ZClMsSeiWmPDTLe1t6t/LAaWXWzaUSotnE6vdkPn5L8VcxQSgRfY
f5cSM9PtG/1y2eD1qJbTzOsfwJKcuclzqbc0STUwiParztanbmZhsMthUyMlwT0DfNn7zzfBea/s
xeUmgxAVg81WGXhS6o88/HfvwGDYSQKHfDSYBhHGJOsZUMBD4UnYCrE2j/xg85OcLGks9CKw5KqL
DSo5qJ58l7VCJzd2sfweoYhQRfH0C7N9DXQOq66+JPg8Ho4LU7xOQ5YgMCf32vRkninsxcu52vUi
XgwzW6pr18Tw5hdMQlYHSK0C+/Bi3LhJ0WtrVKKpWCzHZ6ZkmreXHl4SPPL8xQOtaqdBN7k5jwjt
4SFvDFBLKUbnnAmBOJVMwbX6u/JsKuxHWPgcy25yNsHPx1In2vk4449wLYqxjl1sJqxJtFF/DjTi
EuhdrRX3DYhAKf2McyzsYnlpSPPOyYLACVFgF6dcx8fVe45NnZCEOsfwmar5BjNoyhzc/JKuXR2i
ma9mYuykCHFqjyhs441Z18DUOCeFuyazle8MkBj1U7+mfxeVJyA9WUGv3bPdIxcXyoN4Qi8157VV
9QdycRu1PHaMa4+qonpkJAclyFhP6KrFW4CnDSRa4JukpnrjCoplrbWIvZxuT1l6gUiAOCOA5r8o
PeNKBOVs1cACwQ70+df6h9j3UBRixP6s9jZYPXBvL/V+n0c2NKtouj1dPSYIasYP6PmfGRSnKdoi
1y8Q1pUIQ84Vgmt+dAEdpOQtl2n9BZWxDePkShQewRuOvrI2wJ55IvOJr6aRzxMcPLE/OnMorH5s
UuWITyFYqib3x1SHhxMH6NddVXGklBEERnwGCKL4KlB0RPyC2lQcBeFJF0vMhZATdk5SfcTDaTPA
w834ALaj0oiFkqV8knoDqC4r8hJDsUtZp6SuD9DzXrmCYCYqzsyGkTIKCyZXG2z2HhYv6UXwQXOh
hyFSwLLd0Z1H404yu4ipT/a6nfG9m/oYlkkWh+X6iVxv3U8fAuSubTmUyaxJAsWzpakqubl69ksp
+j3loJ13Uxd9LKQJL6cUkbkehsaT7RI9ddGI2nBmFKITOEgZ7SS6HInsOlQfoeHuRJNTN8fkE1po
ZsiVzGlhIxYcJl4VgETYIJKbr+M5HAakh71woIc7WKlW1/TdSwP7QtwGFo+v2ZkIZsO5mHz8Et4Q
HY6huyZixpwUXY6A1rHg8z2Hc5j27CN39qd01ERI7eyYAFzslZgGMTKCtfiyL9LmIBoXPRrBtseC
ZfPoef3MqjmTsd23/8hfEsPhBS3lBAfqksx5hVq4oC0F26L2zxKN1nRJ4VqD9hTZnAnFM1lrwjFa
JaTOFbt+af/XFnZ+frm16pw2SB6GGZ6jb6nHYFD0hlV6KfLD71ePQ5zeNY9fiMIBKuC3MAsEmuAn
MJ4vBPW49mQAFe+RGf3yOqZo3syneTI3Ztj8GlmqmoAbEwQ9zDVaqkUE8dAwQfuNWNLU56CcFiFu
96md1JwpKd4L2iHn+UR0z3HBS1OxhiYeiDZJQnEdRJElI3UuYvvHq5FrC1g8qkxJMeNrYZFA/ac3
Z5Ht0g14G/6p1MEfLALBPhx7p2WKbY7xiwpBXhEaJ34vF2dJmZsGAWAGz7860mKgRQ5+yorAZN02
TxkLbT4Hi2+Mcpqz9vc73Iz2uHLsrvBMrworYplas4Y0yu+cWmC1hMSNEeJtf9G8lf3CFU1DqUMC
ySKB3kdN0aEfNH0geowbMadQ+aZ0gSL6nO+r+cJ1H3N6KzlH9jap/RoyYFxgzGXwyBNOt1a+m6tG
Y+1Mg9EqbJG/FVJHGwPqjq4l33+7hid40NDqGJCMZ1OSuxOij9uaqs9glZzHInEEsg4U4nZW8dJ1
ZOhpDoELEGtiT+IMgzkWLYwzpj1sV5ayPbEup5zLzcB11juqMMisANiD2vqRPuPrf2vIbleQiRhz
5SuEOt/0rxFRZbazAwpqTbBRbHIYnJlx5qTgX+PHs0BVmeP3VI/uGJPiJkKZOul6j438XtLzVuOv
MZt3gQsw23MaeX4APZ+6EEhKp7qyIvgUNp4Rf40InUsP5NS0qx+nYW4MEsxS+aMcplJ3+PlU2N1i
r0Gcafvlxr7IR9iQm7R9poxmpBNMnS+Xvf89HfxJ5EvksX/PE2jLDJjj7bX1whNeV83WLbB4mGGR
V1XuD0TEgSItyIFBrgsneNL29GN7IsAnRKsJxrjzTN5MeEsU94ye9g2t2tJM86kZg6SFkHbh6AfZ
vo7X79mn/zOSq65d8TNuoizq2bjSHyEdt8nsMOtRYg4v+t6NNCmID5mATOHfNcnx2n3AxSTyhAqx
nRz/n2t6bs+GrS7MLd8sM6J6GzmXdgoJZQv6iIzvg81C4iZqDtFEgjMUMHXUXaStk1In3HTDVS4+
WraY4SYcZDwzHFxSlDUcPX+QQNJSGC4clS9RMcv0p7/6zFFXSPnTnzeQcmExK9/RpKNqAkXCKnoG
MXHCmkObjZBWcawMhp0ma0iBi8hXRHQ0Vy8T/iNmTbnE0+oCGyENvEAJryy+SZEdErlNaIoYKmXh
vQF8O2TqN96mfLxLVY9/E1HA/iNnctzLIwdJtIUJ0s95Nh9OYud5HLlrlle8yStUvbLqB9UTUJcF
CZ1GeiTaQaT7bx9rKiQCGFTOUyUciCuRKVLm7jvDu4Pie4R5ii0fSuE7uVZ0XCRRLjLdBs6HS7/a
tSPejfzngpQXE+d7vGavOhGiJsg4Ymj9ZOe4KJDepwoN4DrsQpZr+Bs+EmtZvp14kyS733AJs71Y
lqp2zm2rmHMRSrgcUvQLZXoYy66B/eqPSJsTO2HIoPUMWTUnJ3TL4hdehsl6+bGzlOTugLDBdVQd
Ti837rK2OvgQAYjeVJTA+DjoaOLrC5+KKBrqFlQ1ndzhBGOWIEj8nTQpCRnx/nRSZqBdRxaJ/XP4
Jha25y795VG80fXj0hq74EVfkalhfDPEhdrlI6zW/0WXMeJN8KNU3bPxoS1Vr8ySnsNf6bV77Sck
QLnOqYyNdIVet79Z8F3s045Ptan/88KJpAJEiTVNqRJ9EfmYtIbe+hqf+2wsR1kUbpES2PgprtJj
N2Oi/ydwOy6S1SGf0lZaUY8b+pT9tMcqEPt/FuTYBUH3B0865wVfJpbAwsRkZAMEbFloXd/XEjqt
ptY0dibQlXygtfZuYZefJkmkjyoIJNY/z3lR+LTEBrnz64WjtDvgFFvPzZfcOjZvBlp2CLtouzX+
kZ7lmYbOtbip4rUM/HV0cwXZFdZHFJBggIUr3jU5w/IuXPQahN5GPNmj8d4/ljomIpjHDRXphqrK
G2ZdmrIp0XL2flVvYFkzQeZrx3ZR8Hhko1NKlh5XgVrRnAL48dNdrvca331RSblCRsr7NZYYWL6E
qfg87rYtX1YrPLXUqXg8acr1kc4mM/iQyPJXVelvivK4jnxFAE7DFucGp/SUMZplQkBiB5SFSL8k
jE85z0HiMJriyEU3+6BS7zZ6j62IPw7sJ3NNkdPGNNz2zJZ2ivzQrzGnLZDqu1pV/1E3krLa74ab
GvUYpKX6UZbgrzjE1+MKXB96oHA5hgq6rroOWUxcPVHNHamYf7gCF33KxMc3HQg7HXoWluqjhDxi
ZuxnJJySfO8CD0xzDarMDsSg0CSaPPA1kPa/bCRGlr/U5qpzfDrDtTm6Mx2sOYFs/t2WlSbgtr5i
Tbpc8XWHYkFeoxgJu9GmCTZ4Btx1cXjSg6xyOc63rhJ9ixPW8qaRgm1iQ1R9bwgO6X1fSnkJDrfs
KI9pxcRtHp0oCaxTrNj+J0Ndd8URRnaWLJotmvoUdHWbRBsVYBt5I7FcFImlPniT/yQGnnPq+OmH
qchGFwhVoKsd11ajNtUOh1TCY0pGHzFvh3bjswJvN8aNTJxrDwV/1fQmwS8f47LAGmUhANf6+9vu
GwU5YE1H/TP8mejy/f9D0yhCFBOYlsGurToGXGuYDpCBkAEsg9ibgDzm0+6CwUgsRfHvaTbHMK+K
AENNYx4Y7G3VJSEA1HSM5wI3rLysbpSgSMYKu1HO3Dzown+eqrg1woky4iSOxdjuWY1svUpxo6u2
nOt9fqM7To+5pUVWVNTh6FhxTAbQtwC29Gjd31rV5z9Rk+Ix80gehK+NhGdBCrkZJLnerJmQdyC8
LWrChKZjX3OhoKNPHX+t+zu4hnqV4hVB7/BvgDmRRrZm/VSVabVl+MWNT/BAN4RNAq++7hnPtQZA
toMK6MpyEo8r81U7UxLf4YqjuSXP3pZg3exkptkrzt3w6P7ozBf8HEFHvBNqFRLD9x3J3FojkWp8
Szt7fuSUrzCAn7gXaN7IT8BbwSLabTKGiMK8N2xvuo7ijZK2r9VXglW2o12yiTkkn/vN2JFZyqw8
3UFDlMkHr055dsFeKqVw8MOLs+h85bYxfPn8FJ2midlrbaNmNQ2IwXsuacuWBQnL4U1DxE2ouDlB
FLJMbQcU3QX5XRRma+FcptWkQLZuSPZ53ehOOSLZapLESTk4pHkevCR8U/g2youNv7qOjMPycZht
TljrWg3WR+3JcLgQbkUjMjGLE9D9/bTIktHu71Z00jxfrP+cp0voIo0ogXC+MIPFJ8c8+nA6t5k+
MROP+NTralGIeXCXtzfWqf/BmuJLo2LRjTfu7m6hpMq338BsAXucxv0l/WkGFoKHWCd6oU0+7/7C
a1/OT3gmLkzLrbJIxYImn79GlJxxh2wy2KAp727bKydhhYzBdBaZHgRuxgqO86Qvw/zeFltTk1Uo
BOJTWa9jU53EwePGv7KDSAMjY9ExaJureF/Yx020xfisR56GjCISnKxmQvMKqV7QoerhTVnpk2J1
sgJESYih5nIPqeMyYwiFkIV5ySDhiHgL1eL3ZjVmNVmCrImhLdz8N2B5kXtVOXLE5mFhRJhSPl58
jSssWiSUtm4heHNRKCOKso+SL7haHuhu8L1tCHqsEgvmeOFIE/AOx5NSstMTRZTBMTn1XUJwnIZW
xKQkt02uzbsRkzwXzcZhimB03y4BSTcsuODzYpysOZNejgcY/EE2oUuENxx60VMV9KMrSdDEcvZw
l4nsC+bsyf7+a1LfcUbx9FpEPHVIy/g6MmCeJjGmxOgK0UlvMW/PhCOdhdahrpZTyK7kuViAOqxK
tWDj3EyGirkadgD16A1VkRhOF038HanVFw72Su53Qh9SnvtNBVXAaWKFWRSu1mdN95pYQodVQzdK
T8lqUAOXC9V+Ww8mCXrvzZfMlOSAn7IEeJviCMhqXyzUeUyepZO9sW7wlvTd8QHC1MqZKAeBQff9
E6HCia4dbKLClkyJZxM+8RrYEFAFfMXxyoegaSmunffGrOEyje4ILb2W70ENsx0fCY0QwgnYLMwW
4X0pGu1DfQ/2castwtAQfHlKKHVnOfnvzbFT+IBa4negCzT38vaHjehma3Uf/QY8twzNKxuO9vHW
TloHooHojqZEb+2sM7vxFblCTnnVX9JmRmcCIWIb096jmo6ablOeuJrsinIYkC5T/Q9xt7pKv/aD
pa9AoaqOVdi9FX6FPw5vUebOjYSFYnrGMzzg9af05wy78RLUTOAPS63ycaxBM6ld3NaX+ZqzNc/x
dF1UwEbytDsdaMfL15gFEBAGiqIHoU8cM2+RcITwXWgtrbL9Fxz4Kk0Jh53nd3A/qaFVp09QQH2K
CHMfbu6aUvwNiDMgXE9bbECaPETyq2LyohmYSIrvldLtmiulsEzyLX6rg2/uwfxzaNWmByr0sLLl
mkbFgLcYqEkOV0TQXQ0P3MQ5uDOWyka/IwM5jhadaZiVKwtTX+WqPPCy7arLb45MckpGzn9bxr8E
q+CUT78kKHvrl5wU1oh7106tV14kcHoyH7wT+Vz3q5yFYQcrjmMWQMGvhAPWv3RL3wi1pK7IFi45
NZIvsHrJF1ULyUB81nBKoBj7OztS72Sr4WNygodYuWk7MstYWOT4SqZyfIFysF33dcqTqWml93te
e/SsrRtZ4sVENL9y9HcKFuYep+SlmSV+bJapPvU8H+0KqG2dwCINErrljl6N3wb9UPiZGfNv+Yoq
NiBknL6FX+dNE9ToSVr6ehw2igX/C9sBNowZ6ya4Ugd8E+qwB+MXt54DMq6pDeQ5PLPxnTfr8Mg4
m1vAL//PFkGWAOryvNGerBlgddmb98mQ/QBVu+gWp0XUV6Nv1lu1jbb0M5h2Yd1gM+dK8FpIwrtT
/QMlYBUgJAdMDvA3S8ntGdXjLmPg4NvIgdZc4uHy8Om4yrjm8FO67kJ6HI8I+slx9VjSK3Rh56Hg
sImlu5TNU/Vss7x1+jzYLX1WKdI562oHKsECvdbHRwC/KE5ZOcct8uLhG+JzWdZPZTmiPWnEQc2L
RQpXdHJNIucjEdUBOhyqBkE0gr0QVHqUc90z7qpzWRptu0boR8i20xALP//C+Klg/t7/sdext+Tl
RRg8mGHiEaEoeAFHhFmw4gbu4yjK5w6DL2xTnl2DOjjTADLovEJh5YZEj2mgcDAr7fQubs+1ihG8
tEcpBrWa1cjN8jgW8Nd1mkm1EICqbVmEqwfsPAYc2XcNMGPKc43QYNnBD/1+gXvFAU4bAh9hlDlJ
OMsNKI9UZXsKQVy7q/xZCCbJX/9b3HCT3mg84lNPGSDPVR3LpnM9aA7uE6pe/5ex6+FvOk3NEOmh
Ggr4kwXnFL+4uJTFr/xwhwiOuG1ZwL/cTm1l2jlekKKZnguOXVnG6m/jHIUn71tL1GAPsbgahhR+
5ovyJnlnhqbEicBX+BY/SElvAmqgzywTnpJ0EImXCpQcJdrEo5IjdTGZtox1WvS6IF/8Xxb3g3hz
YCq8JYrAWPrFj7b14dND7xGYYfnD/Yj625jZZCtBnmc5XIIEj7DN/xRLVgsA+cK4uzZnSLmkmLog
3BXC/VGZrXHfQjWIWibIQHQ99GvoUJQHqLShKfOsTOL1U60iXYvOhIjqoFuafH8ujRX6qJb7dlEB
cN8iuhbKVCui27xgZUz4faO2uPbPWsIw1mqgEi7OfaImnxptDnW9Kj1GcxHQQpp95vO6mOuSMrix
oQ986Flf4s2Hs7pmNMd2wYvTQ4SiiPzUbdSuVOsmkv+nGFDazkFmqtiVeK20TcT7yuEVHUWEWwnA
nVedMRBgmob6IZzINi70EHjOkq/c427ktgjV0gPLBmgg+v7FDvZEM9yzTMTsTyZq7fE0rqMymc/l
zYVDA5do+pQ1zcjTMuChGLOvv4BntZuD+cxvNG6yw3TLo326h29FPhvu3wi3rhFkEKcQ72EGtgFf
9IBDkrrDT0VR551Q/yFiKlKJtwxE3Y4pKg5VTFLzKns7iyQQKQcidbIU9fUdJ0hBvMW9uQs+LCIH
iiXmy7U5M6+5ehzU29NS7X99sSdCZNjnM29BeHpgrVknx1saOR+gmz6jqqldPrTf/hNUlt+Qc8ts
jBCkoX4kO3TTlApib3Gd6YgQIelKGygg5SSZIDzI84B1+c7C228wSd3tWx4Fh0xeBetbh08Y1u/6
KGW1A3B7hSM7EW3F1KRdG776cf7Uwu+7KeaOimIM3nu91hM97kaIRP9o9a47IbOtxuWogWi6FoKX
3nxVpp1ad9P4CXblOzikZc1lzxZBF0e8GzHzgsI9ZiSH7AaWY05577dclm2uBujRXg9dJKMV0267
AVQNL6bvRTAjErBTxEE/hj2gqyKpnerfqeNQcFZX2ATFaCANG11WQaNQjQPNz43I6/Caw4k2UHEo
RNka3kdRCQZB2tN9qdQHv+oeKLsO8u9ft/3nPFlBfCxoUNe82+/ZNRZMkZhUpJ9xWYdRCanoGEww
WAbjNFRAvguxh2njwTIBXo7HkBf55IYVqKgXwYuy4azC2J6RmlwTVgGMkVzZMjk8AjOSihotqnz6
A2isYDQ3S6AoYI5Ez/iqRdPCI4scUXu3N3SeooWsRJKpI5+V2hq2WJF9LEhNs/2bjpZQX2hgxi8P
tW9KmlkrEbxWwU1TZCCdBlx08jynCBbEI6DduvOxY5rnKmxMdmmccjI6RcjzijPDCGx9iDNV+/Ad
St+gRD852fArbZscOPYgw6E3Fwjde8rsGvM43Oi4Ls+7jpziydWZ2WR/h55ToYk44JkbbXtqXALN
urwm08MvWYU8/u58dw5tJ1GPKrAcotHWCuYRgCtYLTGfYSrIeIJ3WECrojsPTj0o4po69f87ef65
ty7baV1IscDvEYoxxJseYbsSbjF+5zy04exp94SC7jxb7tuZnn3gNJOC/ZGs6DB7AoKTp3AG0dcw
+8Q4IrJAD/AvftLlc5OefYay3gScfO1sQJMQ8MtSaeLqGg/PSbjZui2F/QEELluaBAQ3M+Xlvd7U
cYLPxWtgC4TnJSLQZd3PmoAAJmjl6iZHCTAiHQ4RVYZgN1fyAxYK58IavVc++JLyXj2oq58INtVw
oh9+iGIUInj3ov3MpA7TTPxsMEENcr32GcHB3Huzw42aZzL7eH+VvpWgyHw62JAFXISY0OxJQ8yG
fuxZNhIA+LEmWkPq0++ClfnYncVVyCkKTEHA7/Aw5tAJUQsogof8ZY4dfFD4WmOpNJUhG7CzenAu
fHF0ZvsbfdCJYEimCcwVN2IQ9i6/l+w/7GaWAXHjvsenlotejifoLORnQlV0QDrITF7c3/y6nlP1
nFG/wYxY75F1fpxMnxRXW7ajE2DHqhFn0EpSj8e8mS+CI/bsdhJmOK1t9AI8MRxa+cMCb8IB21UV
StUzgvIXll6ds64jCqzYxwQVLodt5uU1ykOFy0ko+SzTFUPYH0QuCtgorp/bU7w2w+D02UtBtZdu
uQQ38SgeDLgpFGQyybLUduJLQu/hUE5qpJICWltYEiC/HM/PYVhbks2dPpF7a7tO09RyLIgs1gGS
g6V3OzeazEoB9s8vDPNuu/8F9UxxLkdH+Qq6hQXf2Vpp38FL9oz2ulVZgzNqWqwlO+SHfMXdm6u9
g3dqW7pf64wY+2v98riWJLgAdpM2lM5YBqiqqRNK09gUFbsLby5cHq+UZu51qIb6vForIxyYJAVM
SuWPa+mu22oJ4n9n79uQNOqOPnkWQtsbF86ZCty+GxWTZWYYN8Zq0tKqvh/Ru4eh89j3uFLhfgEu
neufnsod8LkzBhEbbLZ6OIinNt0WLXdVJmTYwwhy7oR+Fcvui88qNdMV3jahGk+tvJ4KBQ3u1Atn
N0CyR4TmOAglSzewMyMZYhBVnyGRweplj6SlnrDMAeATYIia2Jn5N2ALVC8v954czFQIWAc59A4J
2B3bSSrTYZpB7YCcTBlRxIl+dZ7lDSIcBN2GL4wP7i1BO7hLwoEUG2WbIYxon2KM6sGEsMCo++X2
gWveI8nT2ZvfPoKzjr+lpRq9ojrqkcqgfqjsyGUT0kKWjbBG+DbTotm0+l/bVm68ovL8S/ZUEczq
MfpX5An2dcfCy89WKQCelkn18fvxG9VAn6dyVvtesVxvtlxcoGCOyXOs8UqNrirfBNqsl3lEs5bc
Hp8P5/DGK9Ef6+qDQZw4TZ2q1QLsVbF2Uvp2GEm3I/pzsRo2t/GpgLmnFuAVwRNbr5rrhJD0dZwT
U5PjwR+gjgVTcsyXf1ttPtDHd6yeNIDqJZNsznoo8JpN7UEtoBj+FOcXoEhMQNMIzT5OEx7NJPwt
qA/aoXI/gw0/wPBqjXeHy3q5PObMyHpAigC0mnM2/FM8dxCsDIkw7MW23jI8yrLgOvgOEwf+Sqis
H5hptWnElNXm72gHjY6j1HS5Kap8Oa0vlvLBXX0ekdn9GFsvzAkSfjr/UcD87TOoU/PwDLXwbThh
h0cMeRjMotqjVyqTAXmKxEHdNmuV5rY29lSkXJ3prkeRbFXsG6LLW93LEYMZVK2WLlCDaPWKH3us
FRUY9zzsBFIkmO36UzF9XdE6+50UV/CQrsdtDAyBsipSPGS6BTFY1/bztzoCb/Ej3hU+BlxnonHN
wKvB4PfSCp82061RczRSsz/NcGWnN3BNDWiDIDPzyhKvSS2CrxA+Q43IIiBlfT8xMdsNyEdpN17w
EuUf8vwoJ5DQdTMYbPtMd7RLHV40lLhPpDs1V+rqM6EGSY4iv2QFTkotNts1Sdnoksz4wquXO6f4
fZiUsHn4PSBlAM8koqZ+paoUS9ZjjY36OIZ6QwSj0S2K/GQk5/13P0bVBQfFUOtZVK9FQqhuVQWu
IOLtS+lfx76ozNvMHqxS5ERT7W+M6PWN5gutlXoIp8Qrzsgw4/MRP+BVAdbKM7ziHoIpvzaiZlND
eM54cZD/p7eb13kg8z4bOia+qV71vK/BbyE67xzAghtMv7vHIQqvW6KmKhCsYQbWtJUKhpcbaoq/
Zn6ZvL6vIw9GNJLVi5esOJ6/8g3z0F//xrf8aJpPS/E5MmvYOG3kAA6rpYLEb0aQzL0hcCX/IInc
30wj7dV3Lz63dQZ5sbIhCxLvcu4COungnrfS4q37jVTDMvZaGaIYTP//PX52/z8ZBxehVso+1Wp4
5Adk3RXjsnF1d/G6VgBVqJPCrmKuoSmdizr3xnatEQXrikZg4+F30EfJsnT4RxfgUk1RmsZqGkvg
G+LplKZC4AAguhrV0k44OV4sK7TIqTsogbu0S+xAH8dtdH2vRXeyzqv3sgGieFwy3iPHs8CE71p8
qAh3Hq9R9S1ZPkN4EWmpu2BT3fvODG7L23hf5bWkCOVzYQF5xuoomCUipBelWTLjLGQSwAF0TuRN
IKNePDqnPgUrRommUby6f0gvf8ZHc3ajdqhQNc+HaZlkK/K3EJx8PYbvtBqQehRdPt4LN+wAm9y5
EHXmi3qnUP36d+gde23NsNBD3iQ+Bv6rWtRxbmegfYFpJB99lSlwMqF/vzeeeTvLEoMhwNC005qk
Wvj6gEEhA3ZA2yVjB9wZj21GVwGlTLniIissO7NRwfvvd8kxauXrAVNoKVsaXdPiNp0LsQXKTsYy
AyewnFRZT+FdZjuiM42SxyDMcpZwfVsLZMZMuUKt6nxW1UjPKlPCLu+3CSBM4iKhg+QtMAkI1c6h
7Uwuk/J5TB2r9Hu3w2nvt6uHvz1VwwpuGB8RUiNdsRMdddyTY57f44BMSFUuNpY4JwI+95IT3PXj
dDDXhrO5y6aRfx4BBIA5unoZRvEluffg5b1DHNN70Uqa7yN2XTr9oeB8rrp+VM6UZzLwPaHPyVV/
WcO1Dww/KiXmigqFlmM7D4M+UVaZpPji6r53iwiBC8/xqLwOOhEk/v1gAEU275BmiwA0H/ebEKjd
gbW0erSoI1XVOODFR/0R0qGIluY2H1PUJ2Cc0XtxrsWCQcNne3dNQx5Ryze4ZmxCAWKmQUKdR176
30Tak3iZXpAMK577PCUa33XqobYQKL4kHQDFxM+geSxo3a9w8mrVAioWfVmdFrNXKOieA+VsE4NT
66i0k3wfsWdU2Ff8beNKRDvabKqvUo5Dtd9gEP97bhwuNksXrvCOcnFB165drY4Yhv2LFne/8uT/
FLOgK2nMS5zCJG1ZYBgCroqBCYLTRd03HR5boFbu1fd7swQw88OWXWfNw327tmdY2Grihds5kqmu
i17dREbJgfXZ3MYI+AtZov7RuPTzl3n/vEVdcJT9JTeNCWOIysQ7CBldUksJRahcQLMIp/cFHHXo
HtpDZDOXTmpgcoRsvsaA42NrQNrLn+cMLtpkNlBSDP77JFN31F96ZBelJQ038wFFB7VWRN69nOfo
NGt9fkmUz/su9eOroSYGC952r6pBWa+J+/CrBXnfZYX/KU937mAoxOAgyBR0l3d0Cj581M1klzEK
sMbXaF9OdK4N4Jb90dahsHmAMxho8iVNoqzEI0pyIaOazQ5STUvrZ0I1i5Islq/qaAHSQAokji8O
VgXBj1rKMN0pn66dSD53UbAQPChYaha/B+OHOQGF1q7roeG5pYvqd+h+GI7FeWm+Kn1TtJGZHfdk
Cu9n5T8vUZrUin8haEhY0UdQviRai7H7aVvpv/nSOILgAnntbuypM8RNi8/D56lrPUYRSUjhxZ59
SIwzaFmtK0/tgHLWcqsVGEFoS33qUKkpXlOJBZD6aFBK5Eg1eaOVeVZ2GF6kzwt9G9scLHPU3LyX
D9R0plSCF+Oaj1FoRwGr8Aw7R/8sc8fjOOF7YX3ciPSFRPO8fruG2C8uISj/xuhiRp0kMxPCuxjF
oUip/DqDqpbTy4S9wXmy1rw2o58I9wNtq8TnKydmXUk5i28Y5BQx+wWvniAy0tblMGKZ2CS8LQNy
BmBd8vN/Y7sI4MyCuiLxiF2XlhU0As4Le3VzsUtb80yZNe8DGu2AwvLhfS2Oh4N9bq3PLDAxKmKu
YsHf8IZkzsJiG28wYeVQbftL91eWhcTEdFhF9419QKdRPQLm4yeYWcy1IwRo6Op6hngOLJzl96tz
mJmLT3m5JcuM0yrd63wkNm6dn8zNaHf1KeQDRC2U0jsf4e3p4uX1xlY5AfMUj8XrmdQZOcMUVjfY
lDJiFDm+KWltemtfglKBi+RejQ8vLU8/kad/969xxW15aWQINyjo+uK8s8p97HnD0HZkagyvlqjL
qp+BvLPzPMNF4Wzzne43s3PYwtWQRI2Vgr7KJvsh8y6nry7Rrxq/0itblx103GmR8sr3DsX5pIIx
393LvLEwJEHxXIRUGBqSBuHaqIms7q7MQ2op2T7MV6z68aOSO7/pey4mm6EwpZ/WXNP9+8eBVVEp
a8ElkICKw0PlbCQUnu2/iKpnOFjtwRX9ePiIw/JFoRMYCpg1qAD6YLz7JJoZs2kw5ieRlnuj89Br
EONIDoPlBDUtim1yju6Ev3V81hemhGuxO9usiq+sk2mtIqz/BoytdmSe4zCgWWt/Dt6GKi6u1phX
4dAgdZ54jOkkIplo5WUE88AYKPn+rK6O8lxgB29Lyd181uHXg4eVGfD9dd4foFbBpZimJ8FNAikn
9pRmqEviVgrYZUo9pvAh8HCzMKSA+MvFJpj10HIitONSZ6cdR3tNw24k3B+teC6rRIxoyhjhpIqe
qubpCy8tLBJxSowmTvh0CJLAs1yic5C1xiz++9R6y7l1Aqu+FBhrFVeHXmJTlV3fZsgWa2UW3Dvz
sjN30/LCpmQYO3diT6tzAoXSJBLSNda+j0fVH2iGqFlsuxk8vTT8wRwyjRsvEOnzlmVEJ0Uaq84T
atQ3ExKvoG9HJuNnlSBK5lcK4VnEDUcgxzBIiW+KpMNpiHlZSL20zdiBYVR2Rhc9oHbMFn/0oLvm
/wFFefy3cqeZiL/e47QmsYLpD/7sHJf1gPmFQGBahI4Y55fraHZ/JUqqGARer8EqNT5vAO7eooy9
a3+b+yN9IzHQz1BlaImodOlxzjjXarvwYjGjDBQtOHqUL8NCFwCE6Hey5QR8UwtiNd3LSXEWttWW
2MfnoCeYmE6HjhGhJdTozzoGSDEGs7VI3lBBaZJBvSKweVAQJeqAoD9qHBiDBPkASwJrfRsx01kb
huDI4Ix2ZcbN4f9KGNrL9JPR+09K48KlnCGLQuke1Mo49xSDGs1Q0jjrCT+SeTKUXgEvpntsAnzy
vyCrpZdiZcrJYIkpewTtDvZH7XXk2MOofVoEXQl6JGOQTLLtrKcv5swebV73Z/8lMi2IVubkFkZZ
/3Nzx4oQ4gQzxBQhbRpyfjBiG1RSr2gOn9ibIPaOnvbqlLf822r84wtSIzzlxf1iFtgo0liq5kdX
VD7nYBEOeKluQpPXLQZwM+s0FtSqyaOV76ncXVprMHwwqcagnR2XdB+VU+5d3F9DTm18x3xHw+Y2
ivDAKPOpb6B/pFEniRCqOZQObYXB9SSIlZSxzJzfU5pxsy8NRRq6vpdjbkwhE48ihg0DhTm3409k
tQ4/CPMWUJmtlm0x4xBnlGQ7OcADMdmZQzsScC6lWedt/ulsZM72mn+vA7cmF2x7gS/YmrXHfMTP
meCf2KDxnSKnVg7faZWGMwQPi/OtQK5t5Kja4T8RMt4BDf+NXsQxaANLKhMwl78dMAzpB1vtFinw
11OG/bKrI64ZBhcJsRDaOCFHBW1TK30rVb7nP0y8Bt8zbPDgNsmmKOsNuvnBtRjpDiPxypnB0hFb
xvgsdbAwJ8w0mnC1rP+u6sBVUORa3Z2W33sXe4VD8JZnx9XQNPg9TELOoo4+PZ7knzEoDx4nBCj9
/0DZaNee7nNHAD+V1vT/DUMo6k9EHbWp42bA4R2cp2aSCfBjQOyyfVOnyKDYym7fvRvzxKLQIz0j
OeovefMrZX5d94beLZj4UxAOY9swmubW5I3aPrO5VZaWCkFB+u9Gf668sM5GoV4Z8o9odzpLGlm6
senQvj+FM6Ovn/ssmXY9ycWF5/6Scd9qHcDVf1o8QcVMBMJfY8AcQlTdtH+3jJN88+SDijSGK/ID
17+GuK8lVTN4wUgVoEpMxwC6wYQOsS5mne6gh8K0EhLGRPKnaKoeTYyLnoRA9a/UQHJ8rSBN7tf3
YzP20Q4fLSCPEPME1thwvtyvS9eIHIuu4F/Rqzzr1Vc/pNMLcFysIJ4xYY3r+O3/ntjsl/IuS2uY
SdQgWC8nXdDI/iT+vp3+Z+jr+go9UHCzo5aPoiA+VOk03sbcaqC8EAzhjqN/o5nlJ+HnKcthyB53
Sy2a1eRYbA1GYZ/IvS1C62Qcqev2Us4Av3UXWW2sYn2TKluPvrdvvWed8ywHjmUDsKHiPghihBCr
K6qLb/euW8uRXsR4zz366rxnybqR82/rLHtAnXmZSwS88Oska7xifPVnh31gf/j21XN53MqPaIXV
8sEzSG7xEauodaD26Pq1tZr75WHH8Ok4iALR9M2rUjbRv+tMKA7VTnVcvof7oApgmgs0EUV2CplT
QfEeJe6ZDbjNpQ3bAdRLnexCou8dtCkZ5J8XHpmqMQbDQy9DK04PIUskT35E/hZB6p6Q3N9YARub
PZGG6HV54rehVzdL3u8oVTOpG3uFI1IwguPctPU7LuJOlbmYDRvbWpkmOzwabREJZYHa/G6n0Fgp
dbOlsGObCcWcs5MJClAwYJgBgp620uArsgt1Xr2s8vgiaNyMJyfuOW173syegv7FK/rD/WcvtKHJ
zmHDhi6r/FXCbuzfX304C6s0Z0bK65cHXQ6WaJHkXNU5bISCDzvESvwxsik3mDrr1k/edFZdbiUp
DpbgwRo+4RJ2zR+jBzxoC1fqAJMEDWm3ICWMix0rYmD5qpq2RuWH5J/LdcbOIco0eSZn07usWwGK
E8WJqTT9V35T2074RZLeHn2XWgax9fbiiIoO4nvtbWi4NAjmYaHG+gIK/T1+BQgPrUtpV2K2yEUq
lHhkcTpasy/u1MuTAQsuc7w2C7MMFEuX/oX+YeRhxY66PZ+rHSnmExQbR2gpaZsMoeO0xnILkx6M
gabfwmT4990OrYV2Va7dthrP9d1OXX6t04DwOmNn/82ExVElfM3miU/SozaQ4GR/ar9tgxmv0+T8
1yWVpMksV3ZTjri/XL4EaYKppGT8uyHF5SlJ576T5SmfHz0KuEb7wt+mfPqNBojPrzNPq9JUy0gI
v2zXzxhKRTpM2wdPWGrBImx2+yI//Xg8ZEU15Y4HkM3SU8kXac/vFSBTRj9Sjpc2kV39Nd3wsS7M
tv7HispqxRQD4ElLcsi19T9ohrU1WlP2haSwVXjQ+1LuHi78B5qCY5ZhxCKFd4pdk3mBVYc2vHPV
muqaMNalTWw6P8/73nV4XRwSVF8Gm3h01slVm9d9Vbeu1PruVNywGOwcaQHhqoGv2JVKecDPfH9D
hYYjBn10i9qmW9q3CSCMIC6c8X2lXc+b6JD2HWYbi+vmq81nxMf5E2HuI4eJ6gllx5BoPcpT7qEn
rcgku3yk4FreASmt8xIhgDVICm1ga6bBU75GAv4tc+e9RbpW0MwSgRNVGpEDT7PbUYzbnlVwo4bG
6v5xliGWK2jBFdjdAyPLdcxdg3joILE+PaHon9LOpftmBZBrNEaeDsEr9tjXvPcqYCFCy6gA4pkJ
yNhpY4rfI0Cid+xNl3rhmVi7QgxOS3QLY6tTAKTCV7o641DIBHaXWJEE5MfvbmFHHvubdCudYKBW
x2KwhWak3T++lvor4fpxSROAi5c28p9Meddj7aupddQVyK3Gcp97NVUJ3tpB3u93Io+a26wn0L1r
WY26OgdBji/3G6kPApk4yxTQoJRmFWBZ6bRE6eFwN5Bc7xKNpfKdy+Y+7fr6OLzfgsk2xOcnc9Kc
AOYbB4UdX+sDhYsqpoBlTFdyKI2ti96Xp4jj5r9TEqUxvxRE8z8BY0MGV3Nq/xCJyuf7I7SPEZtr
jwA7XbEpvf+OdDZz77XfR9n0BFoNWJKLolcnRzs8s9HShIwg++qn57WPlw/zaOY6ehD4R6ryIdtE
HruJ5f2p1Pn+Hv0zscRERgONQ7FArqXy70Qn1NtmvBG9uEDxKTorqkpBgnfZ4k7cKNRuaFfU0gW0
pynMKpPqzy5CCEoPse2urakS2Kxsq9STHqb3M6OxUXacPSYMWWAcXE6lrkIDxAEdJsP1LAiVp1Lv
dPWXvGwGqm+su7mck6hqw1O55h6Fg+WLw9lNRhO/YnsXKfR3bWE97k6KV4oQ75KxN6N54qY1yiF+
z4tD6P6p1FuhYtOOP/x82ewQS9fRgVyNPpN2w1nZ+0xG2jjlxTW/rmrGXrBAS6Fu9cJ1qqQRDAPX
cUxIc8G4lE9x9zYcMUJL9wmnn5jeBLyLYV2GribVB2igrVq9XRfnparc+OyHDcD9GCtVfaEorwrS
loyUxrXy4kc0bJxvl5DW4DGgcyOXWCmn78/d2cLa+19cD3rIZrEeMN65dCt02Hl0v04nbsy4Pmc/
vNtTS9C5B9Olb6dOWC5KC57e11nicQftnkEYqKBvVx9H828OZrm/iK8kbxiazYSEk1hG5RyqBQXp
ES3YBVZN+YObjKzhB5IOlN0Im6LK8MCVFOVapUKpgAbLk4LW4+w9ppRGM69YNjk4p6Pfm6r6vMX6
8Ird9rvCw//KndhcVYrHQHXYk+8HjYd2r1fcoGK8UwT5n4HqfoxsPrmIK6whkPDX5HulQsF7pY44
wV2k+4T8qHzl9pG5D2R3MEmdSjvWFR3MftABmzof0rfB7W6mgeHGWmVd9xSilTx3gGud1UkUoFX+
6kQ5FCKK63jQH/Nq4Nz2YyhLLIO3sH0loL5gSd6HG02RflnMfYk+jMBSHi7OCgM2fo10VEHWWDgR
0lEBPcmCdIO21od/s/wesUJ/Zb+CoA3fcNZ7QKfbl3vE0B6jrQwhMKgz9v7ZRyXhVs1+iOPHYKLO
a1ENHfCRSM02Zk2NS8155hETbuSqCzF4JsJNesuGkjPzFz3ERaO60L4zW0jz4qziI/L+bBUXAf+L
kGdCkIW+O5dmwCmXC6IosuPAB3TgMhQrSRIpKCpBD1Uo/naYCq0FVXvMZnns3Xcrp1QcNRUTXGOg
/XDaHuxFueYIaZIIRuJXzp7OKEcM5As6Rx7rBM1AZhhQHsfKqQl0vSBqK55XKcPru2seAKZ4pFEq
pECSuxHv+ngrUQ8y/XnLwn0pDDBUq51nyGIzZD09zmdGkZsHWb+uBZHkMSExZR+SBJ+MQ68x0VKG
+cuN9ZmQnjooE0P9IoJh6SjX7qARrkRrX0f95IUoYUeRxkBSLNUbR73qh78kJjRJr8nwx0awGjTp
t156P2JXA+toEAARiNP8Ic2sT+jfmPFjFyfWRcta1NgCi7QX3yIug8rkGnz0I5z9802wVfKDkvEd
Stb4Ot6z+OglgjSqz6k7GG6YGfAV8Z6jk8uzKlO1JcKZzG0IEcojBcmcuyi5Ek9wYXbjowPQM+ju
v636eN8HLWjY1hi5nC3Efa0n/dD1OGYN9Hf4MJ/03pM1lmygnmLPxii4SLwPIgaJrXd/GiDcPeoV
EH9h6BSAf/CQdST60x8+U6NOFIQw5ko69nZzUA/K0tcu7nTJe7fPFtrknyt6nJgbHszQyM5kf6Ou
cWgye5yvtaCamXj5U/6bSaJGyWf6X9fKcrKCUJ4b1G4S3VpnCRDS5S0/PpXfzAJKrDFubMs0QtPF
wzcrgdSzZpPxDpaZlOScXUYQGDlZiHplki1xVto64+2gZvmQk4ixcCXiBLRcKNJTB+B9aLsbYyxR
U6ZMDdT0UP4G8SMxu13c3mT+HruNrBWIDdAVlC59U7fb5f/zGzcfwPcDVaA1PqhxvW7nbB/DAKxw
2QwiIOYqCyvBl80mnT+/0N0ePCXZgAOJ3ayJ49fgn4qHgDXiIEtzE1vtecJjklUrOcIu1mDI5Vwz
ZjtZXgGwJ4tsmw0Aqr2/ypI3DaFCtiM3FVWFq5yLd8Kt41zgzK1XgHDIa7Pf8R23L9Ck861EU0fU
jTLi8bqxMC4DvwfEw6KGvCPq2YmvEnMbYWqtIQdR2olk/HWMYocQgh+GRPkyOn+0uMyyJwM2KoL3
mHb4lzCT+chwq1wAyMU+l7/jYjrDmXuYMc/jLKG0176Bq9iFXKiOQME9NHdadvSIjpLjUicFd9Us
n1bFwwJ6+vxHgyh9Y5FWlervj5p3jahRbDrpOLmOaGgRSaQGz+kJhe9VR4/uJ0ADv96RacuY4Kf/
/xlcBThE7uWlGZlMp139HyeNJqfqn7YzRSd3Z5+YhMAdQJrU5QGRtmgQvqiVP+4I4tyrY1guDBoP
mJxOR8C9lQo/1wrJ0s941j8/1rgY3sEfwWEi5WtNRnzIRZUn5Z+GgxQ6u5kHnIWHvt6jK/RoMMu+
X2Z0MHmHinxKHzn6bAGA5ngFVp0ItO8Y8BYuTn397L8N5H429IpliR1/0UHIqJvh0Mk1GagD4ho2
Rc2xyvR0cbOzjmkM18WRfotrCB4C/VqjqhM5Tiko+Bezt/JyJd36MvGJbWNkiyQNbo2opfreDw0M
/LzISMaSLLImRgXzv0zp5NQ8tiXW/rpwcsQWcX6vNjojHKintKKGijD1dbpVNVeti7Af5LsF5k7M
bOl0gI2rAFZ3gB+4vKTk0s+Fh7dGE2dL1EVkOIrKcu0RbSGMjvF+lcneWfZAr2tIKeiv3y9T4zbM
0amY7n/OkRgzJs93MzoFjMeww3Ayn75En3qewy9fgcjkGjrbPYTfEX9C6IQux0+5UlGzMfajLDBm
qvgIjUZHzzI7WrhI4lNNNo7s8GlU+kwgswKRBgPScSN2pILosfwWXIkB4ZS7uIRqNhpMnlDkSdHr
r5yEKoSqJHuNDtMl5cXlnoEFMVRoYbrlV6aM1d9V1ARD6h4IXmqti3pOaVBwsJRiFYko8v52rqSt
MdCCqURvF2nPnN5Bt8zHUfhNLTRAQZLO5Rj1ovFs57/20tXPn/0Yev7mlRWMIL4LSemu4q2XLIYI
wvhn8mKPUqujEhV5mlHRTu32cQTHdJCEuZvrjBnP+AZwBt1dRNCow9y3DvPs7UReK1Y0KQ8+lCUP
9JiNS7geVeQa5XFl6YUehVS3r5EgBQiUsHeLSgzcSR8SspR1IaMDoIwvah+jZqaArlGJk7+YlMC3
deMueffqTvGc3cQNM1NErEJTh75aPVVy5jrnir0WXiM7DTNhN7pnbIK04Kr7GqmjkHfRn5y8K4yh
+rAaZP1FTcM1T6iLr0adO+F0TMJGv6oWpax4UQs6YCZHD3pE7m4iJphw5PvpBV9okFG9yf46KHjK
/Bwu83efj9Vxkupmuu3s3WsKoDQKuuPqL2vOs0YRz5/QiGDxTruEsEESzwcft8Qq1BO9K9zb1gfj
8IQLvGaunF02+WLT/oAxA/LkUSQm5eQyN4phS9OSNH/jk9v5WjKiIurQaXSKVlUQYTPua5s0AsyI
HMdm82xIJRP0DSTBUy7HusNcU6uDI6HpURbSieg4ZQY2e8yPvGt/R1NdCT1xhthfF0uE8cURRSE4
nbI1mX5otURedsLtwJ42E4W2PUWwfTOY4KD3I4mNrsY7DHMLnfAn25Lcbh+Kn6XCigQxyQi1L99G
5B+giRv8kBA/wuipfP02yciHuLiJxEyqg4W+izO95hjAUEXRPAOEpMOIF1HE+Ez3pBn1I3vop89H
Nt29+3lJLC4k0lSkyTQaCysoTD52jXFRKwvzVGGgdkq/eWMNDGu20h1tKfoS6hBUb9eebVa0bLEX
K+oR8mx6SIhd4nwF+Z1XirCYKe7kSdlYLAAiTD5+ZrUsofVl7JsFseFNuRPCPhh9fPKz6lxZZgHT
hQjjZtxxtiOod6br6+5R994LQWN6zGAVJSgcnD9QW7LmxO3v0vq0XFC+6BHB1oA2qB32YgCkYYgw
A3hcM7sJxiPgh5qJ52jjy8Q/b27oaQw1jmuyJmZOsIML0j+RkBYC3s6foxEAD3MGeLHnzD08HYj7
ZEBVR/1GZBlVGb3zgVcB5tp9L+84fEzGHW1ovSSIU/blWZubbhbxlvCxIMX9xW5SQr31sOdLN8VH
epiEq4TfMIlQsaYPbvqQTeX4JucQq9KcJYBiRCUMPrEl1qSdgE9oOztzL3N3g0zrCRNXUnY16knW
xbsv6V6ihbiNtrjMnfQLjTDaDIzxoMo+HTZMJbMRI3fIcVM+vtVkvCesHdvXJKZVQ1Cxjb3DrAyS
qp+T7V62qNE3Z2zJbqtU8lUVQ3FL52a8aoKAW1hMZ0LCrIzGhhjtd5aMmabr5k5Roy2nUmB5vsFW
6oWUlErXWRSX+Y6tRItCoSUYZ93HcVw3UOrBvodq3SFZaqo/8sSY7RMaF+Qs3kc+DBF2799/90MR
9SMDKDyMs68gobd8/0J8C7JMXiyqBMoBiYMQC+EeT8h/sycmie+xcY7ehrkCbnZoVOyI+oX68KMY
w6cC088L4V9juxutprKFF8Jpz4WwCLAfUXgidsrOxi2iSpyQ6388FUcCeVkmgr/cQJT/KMWzA0T2
SarGKMzuwz5k0EJGEYU3aLBMmSnhRU/V66CFu4SijM45IcfdPrYD3BwUqhl2XX2NboYzXhjpaWTY
K2q9ZflPxRePewXFQNNAa+vxH8GCsd6N9O3Ib+8vuYJMZZ+3F/dDxWfv+lytmhfqsK3XYhawpjuW
7Ufi7MGmEiuzAdr7peoR97GzJXdnPEOaEjxbcVXg7fGI5/q8rH/caGUOnWtqsTROso2kCTXM1t+H
mq7ve5AyZaaHStD3p8l1YeTIE0YW9KPs/1O0gwV2zAfTvC9VbuJkgPOrSb/+4na0vBAU5S097sTw
G4cCNt/RcrMyzRO6Buv2DeGgZ9iHRZrsthRqiacpoKCCJdRoN1Cg7Q381XKW6bdo90S3dI8vobtL
/O+Gq7coFYTDQ/oXBOgvKJb5ndyvZWvC5By3Nj2cKq4p4aRzQPTnS76kwGwtpMAGtcY/7bJS56ec
nzhM7PCIaUFTYI63a9WtCWp5k4ZreFKbJCADCbhxRp7jldiRHCqpSF16RM2LnwO4aByxkPDT4MZn
Gz1QDCNSVYyqBahbYoRPsoFgSaQFrAMs1IjfcQHZz1/FkdH2WZivu+1egEO9TmWRhsAXBA5Jsv9v
FEu/ACGhEzPu6rj1T3xCHc/ZtZ9LfEdJD+BIuO1dcbvWfeXcgLxy5qpP9EbHUvdRcMiyNM32swcS
VkM/TMAtDHXNMDJBpQOlutFG2CFLsVnTbGIhLakZbe0dPMmO0P4K54dwRkFLMvigoFqUu7T6yPwY
qPEJhFM3Cv94zN7LfAUOpybr2hg2ZrWJBLALrEwPbFxTFfq1PuS005WWe3iHsYMgGdA7TGF9DFhp
h/M/hswyIY6rXnFnl0zcfU54kOcdGp4LASejqzSJjv1kw1a3fR8pR4aqgnsAj7bmVtfAIm4Sz/I/
udPX+pTsO9Dg0xzIKhpvqx5bd1Je8b/oIs2ylUAbafIS1wvUWJdI0cAjbLAj4LgnixBf6Zn9Uz//
0b//PGTut1r1UwKhsGxnNoe5z6RjPTqf0Af61WCoL7CaBdEPo2sZRjpPgiaKH67y/Yz9TjTYnH7H
q0SoG0fTN+hfABEm19ELQDW43W+xyTUDaeGn2hZk5GK8zLmZT6pKfYaq6Ec84JZQByykYExhjIAe
jvcroD3/fPjveLE5LYjbekTyyFP+JtH85rPIF864e0w9iCF/wsHKV6q1ji65eceYozyhJ0Y5uIb5
BeAITie1muo9zrvjL6BNGk2Or8dfIvU9TemwnDBC2ueKO+Vm2A3tVgV9w/5vc4F4DkV2mzbef8yu
GJLCsuohQPf9MYs8qn2rmpfebCzva/Eldng7+Q89NfSjF5Gl59RCSDdBh2E9tCm5cJTjFWqaU2gx
zL5KQO7nlracL+yiRPBrR6LDoUVaYK6Si6VlAnUCeg7lwKcLUhjUcxY/NYCfDHA2gC5TbH8XPqqY
bRjwa9RmGvAB7QVQQbtxHgjtvYfJDA37ZWACeZSapE3pGPPlCk7VjR4LDBgoVRU2jTVAXhz90IDO
gN46RosggHHjy/tDB+ccJaPCgxGvGLADAbY28DbAIbAbLMVvaA7DkA94sC8OUUduKnNgxo/9Px2D
HeUlrU/0g73Mj9gGMaUbMfz54UvDJIMQwTVAg0wGAstk7lNNz3IL2uJDLov9SF1SCK1DqidvdAbg
Uxyv0POwGnw1lDTYI3QXJUHc0C1szKWtOoH28iY31E0OEVuNHMhHc9yidBZMmH5iZ+954SARHviY
RgvuFVq+4LqSsKn0w0N3hvWdzD/aquu5EEflVbjQBbZWvhBEWAOkszyVlVxLO3rU7mJ2rPIi+y/O
6XmAxbDNU1wC7J1i87WzX0sgPwdYNt9BOIgMnWASg/WJ1cE+diAS64Sf2sbnSA5KWkF5hIlR4r5E
wnt+TgnEpGNWgawOrsvoMTBCUYeVHr06uPWAOmlVWMiWGl9sCyS5deSGPdLRL00+JduupNLpvWey
dOjtLBq3YNbnRkfUfByssm4BssZDmovFPY68bviqA3GVGG6uvwrI0gDl452Vr2sq41/nznjesE0a
pR1lnHqVQU6zuCAYY418x3Ik9UpdbjUrKq3JdP0bcMwBHn9WDN2h/b6eFmswIT+Xe/OgbK8hbsfb
fSzHKxOb2eQsnN4YBdpQkVFJ6vK2SmGnu+6hFkeydnX6/eG3TRsajnNDY8/xDIXls4VAeabIuCTA
XMm5CgH3rz/LpW5Hi2nRtCj2yRj1sH0dDNsFE9po3SGqtGtYhFsRaqbI1g2xiE/iX0K71mNKLkkw
aGTfrlvZs9tAuZCPDEH/gpUdafj+G1/RaHOREJePkT3YkC1BSDHOUB6GMzD8i7go5o+agd7nlahG
LQO3px5D1ot67YvSz4V5o/l5IVKE//jRTfl9lpqnIm+uAvsif895IGtIFay+atu5ykpI2//+CTDW
shR2AsrFBaaatiQUYL/FQ2C++tSO8t/adSys7hUD6GeO0esblIUMlgYKQd5BUcRw56EBii6nmj1d
M61prWKqmuPqQOc3Ahel1ignywzaL0tmDXdHj9sJAjeydjOuTN03RAIV6RrUJVGeM7JE0JmULK1Y
MMyt5Dy5cPr2UwtPCXdzODHMjrsJOQ/OIICZhuwfct/cmQXkbGBeBEx04YJA69o74ew6idvnBKKh
xNGg7LdxAgLbelfr/qvWi4NtRg4kF1KLqT9wDTvdZwQtX8Jfgt+RE96MR4ToLpAj2qFePZTwsa5S
276UT0bJqNSjLYG9ZxRm/geVZ2pwnrE6+/Q/CeVxvMt9ZwJweZXDLUeF5qLRgASfi7kBzl2P4DTr
8cUPSe8tA6MbvNTV7crYa6505Tlblr9bjJRivCDi//WvX+sBJapx2RKc76jjbd72lmNAmmeuVyVJ
+nrPUC0ofIrXTXNCfMpFzz42ZRkZsF6nAOW34fYU+D1Oay3H4ONxrSDDKkDMNpUgkI/4y3zO2VaB
ddeYN21bR0OxrwMeuVUkQjDqYtQ+5Jj/PL74TsDUz5Wbi7ry0Eq8uqYEire7FjFHS9FB6clO3wgw
fvB+1r3o6FzEdbYknAPdCngVayNAtrKLKNjrEYQ3oj1QcbwPMuQ6848r1NkGcZsPU6Cwaais6CDn
rof2H1pkWhZwn+ducjlYqBpHsWQTbpIhyRxXFDeHQkAtG8lKVXAMXEyMUUtk3RpGrpK3UTFrueIh
DLXYX1Vgp7ktE4A+9QXppBBiRB89OppqsyXHc1IKLA9tmyLH0bmEKfx4dUBpVuXex3yAOGdgaTK1
gDH3SfHeGE6zngPsxOY0cW73+ggr9kQ9GLk746m5CB0Qcwn5740cYv91BtpbJ7xyLor3EmovPVZB
pJN8JsBvHp3VZNwnLtUFRgDfXrWdqN3EemmDZ2LugYZ4AG+phvZe6blhFVdg2jo8Z8ubapnYuVcd
LT28ziMa1wKwsfHyVRZyIaqXoVvpDLN/IyCSGYW1C/zaBC5JJhI7+6JNPCfTTInBenF3sg8kX7VT
6K2Y61Btz7WCblzFPlmNM2ylYO95QsMs0pwf+PJYZR1eFDJHR5nuMFx+UTOPX9FojD0wPk652Kd+
vDNUfZ0Kk7gDn1L6JqjuYswVF+QDXa8+aK4+nHSFDOMp4xM4LFC6QtrjW2V5lZbBTMd9bfcRocdP
M3x8MBIBvxvdY/ppDvRAtMk7/t/BWrHH7tEF2uslf7kipWprpAvbGMcoV3BLl9qE87n3tKETFLNc
5INfE9xSd19CLLFe9WT81n6NwuoIw+ytBJBQvy8iTdD6vAj+f0FReUSPyYa5L3Chp8Q/aN0TJoKg
TqjgWXat2qXnq6mk86tvl2n8CBTj4vPquXktbsojscuGSLopNZoTI1xi1fdrudkDuIOl1AX8DeN9
NmP9VUobpNWv3jwYcctrX9wUVtahqpcCKg9GC8dJMPkbXK8OkVkH6krO67ehIQpo+b9+gKw20ARb
TyR3MVDIQwq79mKhd4NOAINApEqDbvg7UYyDbSr29YxF3HL24ZLEUENYMqefCRMf4hU3Tjlvv1Ss
+dJewVH6BYhkaLssvDVXLq4YL1SU68cCRY/d3TajGu78wFPMMPt5bopJzP8TqwDtAgkSDloT0k7R
kkJ99fy06JEnGNNGmZwbgBHXOw0+aBSUI5gc6RWaZ8RnyNLbrZpTTvOEdt+hk1rcuiuZkiaruNYu
DoULMouum5ve7oqGfMY/1A+tNj4Qq+39BIaHhwmm0uBnfKvKVKkVpCc1l+Il/y3VuCk7mHZ6XO+V
+3ubr3XaB3yd34YMwgjPuR3gv0PNz+pffoYy2KgeXSr1XeUwD7zWQ5YcfU6qV/3vdCDX10lNgKqP
KI88ukEvxPFIKmrw1obf2kKOycQ/3TBIwJpmGsAUhTPzTir9wNdevBBMV1IZMMITX9IEiqX7FcoI
zmyvnyui9UG/Q1ec9DDk831V3I4GWRS+RDjZ/RfaVo4MYclfeZjZYZ20lYPSizp0h/pjtK6L7JPE
TNcjhgr6eRWF++KvTWH1wSlyx8BDaFFvrJwujjnPryEQMiraMl32ZFLmD2jx4gj02bzfX4Q6M5Ds
k1wSxoxDoS2tUPoN/VwVjeKybrsyUjMzmdtPeKgWTJm+2B+qV4qLfk5N+7YkzsDXdS7dXclcLQ91
VfBEDKHP/iCMTmyVVqaoHyFmJcxyP2sGHCQn46aiaC/Q2gomuQB2tkatz5cHB+CNGHqaSu2MV4mn
XTRYqE53EOvorXgnlj4hzNLWZ9JKIpdYEA1auavT1xSziN3K2UIYN6dkMzieZLQWVY0yXUF/yqxW
7dqomVV1sMiC5JPD706BwKa2OI2bJb6RbwLtApSOx/tCxRl38/dhOU6VzZ++ovudAhl7PkjpFhON
X5j6DLEKS85HtZsaOEydKI6nASpba0BRvrN7nk8tXjtYC0oh20Y1PEQE/cobhYdr7rLP8ZmDN6Nw
RddsP9nKQ7qqQ/doEo+SuJFmT5ZJ+gdp4ckgpXoMGBwsKDPA8sqxLRW88mz2FsqyVkt/zJXyVR9p
cZ8dacDnVDXsOMNxY3QoXcMnZyisoKlEP55Vdw+d7qA4bgCAW5/v6dzgU2/yaQ02SpMz0UUG8qmv
YIKtdbMMPY2DnvwBKvikuEubf3OT06AUOIFqQXy7t451IJYLytNkFRvWr9os5iOjszWnZiTUd13K
GuyYuzN3ZFQxBCmUb3mutmSHzx4eQfOrA8B0JHI169ikuATyDloa4vEbC0tOMzpVdMqyGsijc4oh
UAnAnS1I4uTnNFl04YhmNHvLt+vX9myVq5/rAYvhtuoVrav4ak85HnpgmzrGczGB44nx3op5vJPC
9Drl27JmNIA5DqqPdRoMY6uOlUvWVDblC3flOGmxbOVXA/mQyPCg0KwNBlrbzLpr5wO2AJL6An/J
0bJncvsY+/pC+q4sl491N3p83p6PH5C8iVF0jFM5f0YL4ME7kupmel/WE5Z16MkcUgkGP4Gf7jah
6o7IaUCy0Sw21Cx/flSHNUj0a+F+/AbDO3EiazVWkTxIdr+8Oz01fvSwJYVYCYthPypN0MGcEeJa
n7NptS4tPLh15Naa6/8dK47H3lHWBtNX0eZQjcgSP6WM9qtctue0fiW5xXPF0TQNQKF3LBSvuzJW
w2fFA0bN4bCNdMArusIoDtHPndI0MmrpExgglZoEnJyCP/6Y4MHlVOP8+lV14FpK+AdoH6wYk3Vc
Wi7ecmDU/oH3EEgApLqRKdYY0qrzjGG8xCUmJMiUpFPlZRb7fZtXMUnrEI0jVU4w+8DD+jyZdN0i
EdaLiZXEsM9F2PlCrVTFU8gnovOSW0PrJiNrKENZX2dGqu3s8s4XlYMLV9SzJ49GFfPQaeqras+s
LLCgE1notcBo41QIH+1IKEK0jBkO8LChZ6pEAWiQLP9KTlFtVXe2bZ96Jqth5wqLLwQD1h8kMPgC
RgOYOIReVkIHOsDo3ntJc60oF7v5bs6iuv4TNOksweZR95TKyRl/uAfnQwNPzk6MEO0eAkkNh/cy
urdfhieBTxy29cJfZoz93pLB0t0HmP0HWzzbiHpycVciVF0R+uwQ9h5/pUWVPvhrbdkY/6BXkbTW
elKw5shyXDtkFPScce6lngvMqXxEpaUmC+DqzafCfQxa6Ts77dMhCOpTMlp5k6vZ9Eo7fX+95IWD
9RcU0yLOVtSeXe+s+Tn0nwWFESnULzgCW/cmLNxetZ9+3oK6ZNCbteakE7jvHM59Eci4hN823uOw
d74ALqnEXaJUCnohwtu/1YRuU9oSvpNr+WrICjUDL0ZEqvkTY3rPc3CthNSvsPkif3CNtQHBLYsp
0Q62ToSS9hn84Puajbcja5FVPhcTRVv+Lq5/t/ZmSrTSLb9AWq1kOdCv0GNYIVCnnGuHSXcGn5oT
FSM07dUPkK5uJ7TD21sdm67rMUybmVI+Rsk6NJsebpGMfL31pai2JQEN/oJSNZjejbyJEPvLzwHE
9VPSXIIRZhDG4vJa/EuXS7o3gj89xXYCmrxqtIqVIm9nDbd9/J8pDhKyD6anYZAc5IVonpRILb48
o8WQtu5PDtg3qQCWApU+m0q/jXufiz/zhUT1OIJkQ0YvDSH1t5KeI6UpR5xqvN/nPM8DVYu45pab
gSX2saPSYtM6lKeFJkBgg49WIYPh74lejJg79yTMyWYYmAULbDHBkrONo7BDXTRyP/3cYDb+NUL+
uxNdvcLOz6fdP3izmXfAC6mrXaiJxbHfRPzmrSv7yxzxiTZq8FQmxv8VPk2EJpSOYYGQYrPt5vE7
h7NGIih45RYCcyg9Tfl8Dw96wItfg7/LEH68AAJkUg0vtqBhPZVzW0Y++gmAmxbphVX6zy21lGoQ
xB4P6oov8Y5grY7hhspQNLQk/gX0P3Wkq6psqOhcKV1Ghqbp+cAB75HSZBDopqEzZAbWe9KYp+6l
yWch9U//CC97LixBzNtJ3n6S/c5bo9xrpVpipiSQ37zFogAUyTI25eakWAPP4sGIxQzJe1mOCwR4
fz4sKgt0PjjJjEGYHCyci5c4SJ6J6WuNVHX8nXsbSNVGbLsrssDWazaP8IRRjHvMh6g63tB/4u61
NTTI+pXkox45w21GCV7Sjti8tCJCJGaCOls4+xbgTbTgYv7CRlVWgo7zokAZERiKxCmybajre1jy
V6ITEp+yrbtA0ZImUOYG1QF/Hvn4/UMCFjH7iWhoAyqlYRYGyUJrwaDf0/QXcTB/QVXE6xOvkmow
ka0vRK47YSnSFz41K2S0PAW8OWFndKWs1JIE/pFdx5lS8Tjl3HWzFGcvKVijJ0PealWU8AmmmS0h
rHqoI1yXupUw13Az7GPKi037FNyvCu115uSkFALdagFMHOJeJnQjrW8vqRBHk1ndBPczmWxKtpsR
0BQzg/icFL79Aga9zp9/u/xQjEOpg5qSs72iXuVZBwW+k77EzGn2aTKeHuV2J5z3AK4Pkvm0r2HO
LyGBcSU6g/kh//EAINGGXZWMr6b7nbBqyvpBE0g8ik5ARNxTmPLN6HO+oNC6BAPnSAxlAyrw9l5Y
hokwZrmv0Tww9rW5rkJT5Q5SvyCwgfsUBoe2U848xDJmBiIjrvAFJuvjuUGsmlpqRflBE8k7r0Qu
WPJaq/5437skuukKNDVPhAPjeRE/8J8OybRXgsNeqmkay8ZSxXT3Ktb+J9DCYnWUjjPa0Fu/Pi/m
owacIzpqg699CE3idD1HiQXsdA6tW291OyqZIuIU9/mxXrywsQbyI5lpxAJs69ocFw4X/j5eLsbR
SCtcfvoVJ1PUzyaC/2tByThuLZ9pB1ADi099AsfL9U3KunzIAPhcN3mKAXkDuloOr1SS8CQ+8Sw1
GgIhqHVp58QuMuAx4Gb6Q9NXafW2Bby9Eptl+K7jqeRaM2F679eqMyRRi5/Y3GVyDi0pfzu+FIYD
pwOtcIU2RdkzMIQnJtxZPzSgz/Koh/5NjvdSn6Bu6UkxkHIgawwoskkWSp2EUg6ICG1jLEUUskYg
AZFvflbffvOYoGSBnTwOIrx+zNuUbAZKiNmXuw135JDvnp7NO7achpPrRxho22GPopwiyNPVoEW0
YV3uO1CEhHpJxAe31qBkV8Xwvjj9fYdtfDQOCiZXMs5cdtLxQ3vAqwT4SIHW8wVkH4NcMhrGUEYi
rrO1j4OGrixflTM4koE9WsaeofObevkYwOC8lKH4LgmXTPeuyFxR3G+YoxhwDc6G5D9jxuPJxaHp
wgGGUMxf2kTlfXEp6VpMJu4grq0A4nvD/K2aJmolPn8N+6SCZnDJgLKEFwbUUkaqfObHdgWLWV76
pM08S8gn97YTi+jmvqLMUJSh9e0aBt0gcn1+RuBYZgVU0xNZrN8w3mQkJP0R8/45MV6GAve7vvZ+
+ecfQ1l33zRnstchaJas+pY8Sk8oygX3ajEaqAfQa/5zGi9nu22Yz/1epf9cUdVPMtNUWNwh1Dko
H4K1hKlbhZ5LFQuMHQi3BQF906ot7nKjgVji/bIuE75CLbusAQugqHGb5jROeRzAsnNh3TTzUSmE
NSRVxlWBx/du+AS42OmndyryaFWjlhvckpnuY+yzmgjTBL4YNWbS5iZIFj2//O0uR3CR6jcWiz/N
xWlhm8errnaTo75ZayWk8aLXcbsrspxLDEUMCUdwBVgzk5aHNkxBQYuXK1FX9armT+Or1TCyl4mJ
IGr5zN+Ojv7mhHmp5100+lv3xApdH5DT71I2lPQvwgU5GRgAjAujXkShHWmAc3v9VLoN0+7M4LN/
E/Db5eJMFoCCY83CRiYS/en/pNM7u/US5wySJ9C7xU4BOOSG/5LGRDcKUeTEjRYY00vsI/6N0CLf
H1CLvgm7Xoz6J+sJ6bMHgxtbEVVEsJ1ZqVkjx9PSOsmKD3NHr3JWBkxZNR2mh3iLlJOO7zzRK2Iq
miwY/t3xWsewVDeEld9z5zbrIJP7M07qZI2kl6xajnAf04TFnsThwtqs29hCiC/8oWEzfkHVupwB
uHnAfWnyGRPDrmcq7XKZ3Pa80PO1RePT5pTvJYfERfqWyjZHa5J23htcXXhvHie83mbm7X/xHWT1
nmIySSCZ4AFKUJC5Uxyka5lz9nJYM+pYhC5kooS443DjYvTph59/Li0xzCjkDykKKsds52CodNMp
cy2NfR0JI4N7VqhMmHTNtg1QHIHqxixnL9289uAShROCFzwj00+TbZi/DYYEIGZCi98uvowz5RD8
6MxbLm5UxMlsu8PxXMyd3nI5eoWC1u6l67kYzL/cET4+3LVCudgmbV1PyTYr1snQNLYMqFAQQZaO
WvRDuEld/Yh/hIJubKkdA7qxCV/d2T4LxR/94A/bddthatBVDbR9bKwhoUOmQAx6NDjQtRFgIP4O
cBawm8BdWUAGMKoN8FwT6npPO/ewuRH46YJyCwOeenAThmIWQ5+r2NhuEFiAvgKJ0S+7p3LH9Osz
FV2HrkO5Ox0MN/5AT7MsWki8nQks2P8yNeYRbAH2jz7R8EEEyZDbPBjidZopryhD7FrQnPP7tgeR
rXT1Z+1LmzVN9JcModpoulmuNbKGM2bF//eoroIfAiSP9qwXCksy2kqreJwkWdml5c/Q45vqReIs
1FW5uglHDHvDHHdA1662Afke22aFQ9fMwry18cddF0T1K5AeY9Guiyc2SkotVOMqSyKs0+q0SD7M
6a5XilTf08GR87tDvbQSxoBVCj0IVGS0RwsH4U0LJOxavP97YJy5MS9o5QmjUS8JJG5+TxRss9rZ
ViggCy7MCSeTzKlbPqVgpRa2cdUUti4ZvTgBQrliXFHzpU0J5QGREbWfN6vuaR31SS+lwguDmC3z
5MFVPpYn0kFgGD26YWhZYYvSBrMofhP47MMgN+vptK9p9qSvP7NMhPqkT0qU62AurqC6Etqj5gJE
0llTbb/kVq5U+RDli2lnBFV9ytzhD5FZ6uPKsc5bsHhmQiYOiEoxN+YMcq7GzVv0U7mn+SeC2SY8
bNMddfyvicQFOWnrkP4jHHA/ltFzPKxe9CZ+g4/27FprU+VUld/ZAZWmeCTVma31VEpEf704b9EE
40ILibWM+JtlDl6YJ4ezd9Je4SaWMem5ZKyvieZhEDKr/F2bTNKRjai4vzXBJQC9fU+r38Y4t5wb
aTiG83nvpbd7C8OSjIDLCwq3dstAWYTVFrxXPMYk1OSE2//0UngRK2ktXGesEZBdkum62YmdXY8a
H8niucrxi9xfGRYhM2deWaEFslzli8l1vAwK3QwDoUgg/SzDVBceMy2/owZ5fbHPI3H8aNS2jDZU
dmVyC4P06nbM3FiZOYpC40qqxsZhHq5GspNGNkx7a7hJAqlAHIYCxB4Ie2GUFkFhkCtT0Wstz+3v
OFE9pqFX4U8v/CUOxXzL63jhyZUGGVLHxg/Zg3ufTVVdlj4FoU0OspkXaUC1/IBQrNB6hdRPHOVR
xJplvqTmnclBcrvneQz1jFBEg78rGql02jEuBYQMAUGYc6jax77cg/JQYF0czkrPlsLm2hVlIrjX
g9U2G5HWrQ9A2F8wkmx8Rgs9VhG4DOmthIAvIr3CEx0MOD546ZHnFcq7tEA5pPSZ0tbFewtixnQr
GhGL8P9qfzh86teDhEYJfBXT4zMtvlv8fyE/bCzDw5TaLOUSh9U0Y7UYvP9S6Qxa5pZ5jbWj5yxq
lcqfkb9SrIcj+7m/aL8uygqbiH65LxjMymeMy2EpyCiSurlUpGOuEJ6KOa1fHaVx1gd3+uxo80X5
q7W5cZ4SxdYSJ4hzF+b/tsfG3q0BZiD8cWUg7jCEplzCW0vtNFBfc7PAbzObUbFZ5Ty9CiWxHk8s
zY976tqqK17Qm2uqaNBn/Iji5K7qH/kpqGF2TrDt1IgAtcRnkJV0BF2bvKdVB3IRcVRdQIzMCvV3
MHPSfboZRVWTUNMbZD5Q0pxj+nFdiH6Z9ZopGWayaAxjsdo1tsul5cIsjYYV59GnrtSBl5+ndlXj
cwRG0VBWtnL1brK8rsnxacnRIpO9++cSTFNwp49zXmbvixQf3XHXOCe4lT5EYFuMXC5BkVVg1asF
Nk1xqFwtLO6Zq1JWzEE/Yy9hYRhJk2qKNClwoDOWY//1Nn+bS1csAqKiJXcRU8BVJ6iOB+cFJhFj
+lhhgSy4P/QMsDIlu9/KMy1xXXPXrStnV+fhFzzn2r/EoX9Q8+C9k86jppnz7VEk1IcB66uat5Yl
pwDgs4fjMLCc/2pObOAfo136C91eTsMknyrH/l+bQZZ61xF3iOjvcd0cfermDviJ44B3Q/yRgc89
F3sRfncc9SxYIdLzmbYPfJTORMnLjuLoSgvUzlDkAPtdCO9xl0pPXPMwHsHThgMfBYR18tXuZJPl
ZYftrCdOTK0b1FP5jaA/5ttATQXeCeZuIlhki7xWibEwSiYtK/yImP6abIcwDe4ms4cgbfa3oeVs
7FNWgDmQOoL4z3hGIQSg0cb3tOvTr9uLGHATAzNwmHKQ01bEUE4IDcgUETWqE3cpD66Ph86xRsrA
b++m1sLwieTfcarIVzvE/hcdHXFeQxWDMTBJXEz+lJrqqBZFM0SSUa6hmodxtIL3dSB1BKpvXHf0
j2WMapFbLyrrqC6N8OvebaxtCNToC9ZV5Rsy7YsMU39AEhqqHvLuRkK1QiDBFezqJlIcDRgCezIA
qI6NSvparctzXksZb0uXUoGe16/WfSBA7s7uVEvPo2P6z1FIyKnsSlAJsiixMAUk8WnACF6ceIsm
CY1LS2wnmMzNSCpMIbKsENfKa3Q5rVDZgkoFctiBORzjsPJ6fPN+BgXtxMiS6TvZZiJBccj958CJ
7dGXTnAXClqXeg8ohuSZ1qd3ZfL/SEFaxWJ/p4IIKl8aQ3QfANSBvdRhDkDtLChX4JzruNWFHITV
mPcQSjgm/OaSej9Ur1rLHbqgZlr5boeK5IFqaYXapFS4ZHk7c10i+zPDX6eXetrLbvTvSKbWSguw
3zfGhZGUElIbotp6B0tgeqADADZ3aUXuKauLcGmFTIs9InlB5IdJ6QXbvI9XaVAwvKwy9W/zSReB
zwxIhED/JMl91kJfVxf/S8vsV4GwRjzMcksbAIqS2HmFclp2qQwXIhHpPr+jxcvsXW2nIAn/Sp00
LCtm2BMgBs190aQ/Z9eWOC1gOysnG60igYjipeCFA3gfGL3q8+KVJad0rZSrnk68XVs1bHXq4Y+u
0iKatTyYA4HIHpAbbkv0+YnyWJmNcZzVOjrDRerT9t0dKpaNRqODWVtXoszfFmWmO5XfVfsCNFKm
Sq7DHYOar4LUGCWDiT62CQO6S0o5BtzQGLsXEwb5lFrHnV7oKCuSGTRaltYEBTUi9/0EV6IQkt/E
kd/sYSMWECmE3pBetEsDQnJ4R+RDEKCvcYwDSJIb/rLmdqbT76sMtGY/eOGQ2lzfxNCu4WJyn7Qq
VdLdEuzf2adFYPdEHlkZYnO0OEZMVlMVyuNafQr8eC5zjyuAnP9k301W/TQVwT+AV1fsbMghlc3F
ngykHInvDpUiE7B+vsUDJqNyylM7AAQDJgH4pRXxORRJBDefeDDjcU0gyPqmKg9uMHODCb5SWzRM
HkcJZ4jWNdgKv7d6Euan9X0i4+KVf00a1Y0O7Xz1rpl8U5vi6byIvE/kqxG99NMggzHZklL679FG
sscXiBY2uK4p4Gr0kU0RkWdfXehCWQc8gJvQAbovTJg5sEIdq8kzayqHTwxZoXDvuAcrVDrtC59b
qRpzjdVJMUzSbjd992A3W6lV2v5DXa4zgv6J90JqHo3PdFPye/nZJqmnoJAEqEmH6JG1OSeUoV5T
UJ4Va5TGQ5EiglA2fsDVNHcq6PUFsgKd5ls7TlbunrJybU13TGEErt+c7AHZ0GMRopHQYpotIbNx
FqmXRzxjNzqt1OSG/UkHEc5bc+8bKJYH2A38HLRlM9nIsA7iJ6/QbiVuaN70dSJ7OXFnPnKju8V8
lMNTWJbvdbbpHynnQUxYjsnIFql8jnKsz5bMc9XwbVsrCLtdgTb4mCYr4kXYkHPEc994gGSR9jJ+
iXWQl17bYp8G9Xx35r0JGa5CbWehx2ORswfBv38fL/5HRbsfaKp5ndpxbZI1RRSS2V/KbD68K/ED
CQk3b8YR/VAb4q/7iGsH27GnCenumuue9SzkpWezJYGxHXM2MuAHGH5DDjosK9XxONzDAWi/c2+Z
atnaR7IP6ti8k5CpvcOLRVvRS8w5/CRk93Zbhy9eI7Q6k+4yGjjyoKKFZ28+uwe9uoVIxdQbLZOY
SCVVNCgG7ywkTskwuh9JPrVkvp1+pbIg+D83/WBjftUGW0qlSQuOakuQ0KMFM6B7DD7SveATKzLR
DRtZ78QYYf/NORyAGrVhjZgO4GB97SAYVSTDh9yWwVjfyJH0+SJErEl+z+/WjYj4dL98BrBvcki6
MpYim1YqEebKLicme+pOSbs/Q2upDJ0ROcw0k6WibrQVuPE7IwzmW5W76/rRqEfeV73xu5UTgdir
nGSEJ72LUyjmkTMq+4znn9GcjP7bRYgEQSDXd64FDNwjO6ipABmKH2AsF2Byo0WSloHI3U5ZcyGP
ink1Ad2czBfb8yTZX+/faaA9CUcf1jYJLKCqVrI+gKXPkPQLtrubBZ6uYE+3oFvFmxQHwBbtDf08
EuotMI3ButBJbwhPoY+vObfjZnTplRuhbZksUghWqEo6ljTO5GW4TglrVB5LxhDdUVtDrwkOCRwI
Ax+wlUMF2+8W5WvqSfORzCueqdTT+4ykAe7eij0ecybXAlpUKEdpmVaWI3GF9NwbrykAHT7PmJd7
OxbNKt1ia7HQi1Wri9Or0dCF+MdkpbNmgj5ANn9e8QYy3deAHr4t04mdA05C4roV3yWNhJxGIQ83
/bQza6bXhhC1lBhdDl+UWbjbU5gaFRXx2WHefA8XvmJ6jOSMeCH6836rY5UvuJfnfLVaIp+/SBLG
E37qNLEjXvK2unHZ4dIFts9HMCLxTb4FgZEUEM5+6gF62UaKU6VDpYS9yGiWy0pTh/dS08M766wD
3oPrR9ZidpFp3S5iwOF2RfQaC4udR7N6ftmxBr4LxLakgAnm7nyW1Uog9sNzxf98uqGu2VouCRLS
Gsy3qbqONTLonHWfbw8qF1O6O3LLgmtVXXa0vlSOGAL0m43Sn3/TObfLyub+bZgYD4L2/bH0iP+A
/MOzMMEPrWaA0wKGGF2vlmMjztTAENt2GFTnAZlbSBd8vuG6CMnB5JyYicBWkIR+n/5PUZ40EHjs
JdSwiXL57ZQRCSsei80DvnA6suLLaGRHH1ROsE+hl2V/HObj66WxfcmYcYFl3b0kCxfMxV1WSNyK
WMM7oXDfOUNlFdZ7FqnbEqLnNnUPQ4uxbksdXqO4DtaSPcYDaY/jb7n4W7br5m/VQ0sj5S9Ook3+
QUxYCUFqQlCRFKx2N6OlX3diNnQZLWb0NbqDF1hTkiD+Vxqx1I5PsNq05ckIMJBNI/xB69Zi4MeW
1gt15AqGnAAQWPqf7v/Hr6M/kzIivTF5h+lyvC0Kwj/XLFSzssl8NmnF472nYDtj5VPetH6eqfDj
RTRopge96DWvSPWwaHEgR+s+/1QVhZ2+wgwMvrWJVM08XwX6HEzUeBjuwph4UdGQAjTOUMpgvohd
QowloxVfZf5duIqazQYVkDdDErz9tV3RfMgKv2xX8gxwT4ukMqbnGNefDyef69WZUbulsC96uiQM
CMfJkn9Ku1kca9LuNQDz0TikrdZduYKth6Fh4aIcu6DstqeNH+hhc7j4a36866gVYLrbhISer0RP
N7PqcL/SG0iqeHU1hq/l9Azlb7txGtVswlKOMrv/cDbFsAzHhIDRkTrj0lCASHg/M43ysYtxCxzr
VXOSWszLZk+eUXuS9+nvapTkLJApFgQlxT0E74+bRWcTrs3SA/aSclWyNUKn4F7y0rfjjkCr57Ro
qAYV69sWVFfja99I6Pq5Fs+La10RMU3w8OyF4DQlbxg2TlNurTPMZgZiXnd/f+TBeI/+/xAdFIZI
958e1CSWcQP5fTlnl0o3v8uGVniIO+5XW9Z5m5u7bsN7gseV2+GKj38KCR/qo7MXGd9tA2He/Ad4
q6atNo2eVs5ZxeCQH4k5lwMymwPZrUA8ofSLGdvJXUhk1lSD7ndbLObAFlUTKsxaIqsU8ISIdmGL
cN8M0OUXtSIvbNU0NSx0nY75/JQAEiWk8WoNrog4HTjbFtNE7jYWa02OfpqwrxLamxaDmRhgfTge
upHpTLuX3Ebi+51gmcD/G097mOo9TYn00U5qOY9z5R28BYJGq+GvqaCZUF76qQtaNiCbARzs9sz8
XqEvHz/nsq6yShAeupEi/Ng+9QfK3nLQNNHbAFBw5pQrrPY3e+AD+y5qPUbaIX3GqoCC8lsp4pZr
JPwsRMBgOvGEcysz5lsuzBeYfqbybYcwMSZvZ0zlCQcOHtA0qk8koBClH7UOqo9ptZaebZ2oeSNV
jZU2oxyWGWKhxOmg03K4c/Kl4cBri0jFuVVbv1FUphlR6BtgXFXgdc9ph/ptPZ3/oC6KD3GhYhZc
XKqbViZi5aDSAD7yFbZ/7LAeOwSIKjrwOlkpm+Isu4XLwHXNMbCaQKsuGNo+eFRKWEIQdzjmVSLI
EtfLvMYKTXHFveKtwClODDleovbKCaN5YW6Y3+K41guirSn2zFa+zqkH44GX480K7EKV57fJDivX
tjo7PsivCOANURa+J005FHaiadDNd9KnIZL+f2gBQT/jNGi1z7grxZq9qYgcDyfOQlppxDFVcsCI
qY8YmK0BJYbTUjfKc/swSgvRU3E+dZwoEgJzGBY+Co8H918TNSfzC9oMoIY0ydyEwskZORJJuNHa
v1bRK5YpUhUrToKTDmpfSDUH0vaRyNR09WT+piAbvrlcw1PjZI8uNG4cW3ZuhHZFmRY2O4fWI6zO
pAYq6gs623nXAdU2fD/GYJ/4zTttuTHf+iJpDd52Veg+nTyw9XqwiVKLAAZlr8kdy3OmET2IX1K1
umxTLg5W1eYaJc73rRJTlRBgGgqs1xqtZ/jieCLlB/73RGToiywhhYr8MtRsYMo2i2rwXd0VhDC2
fE7ybfUYCyyr7xoegAsSzBHBqh286lv0vVUtmYzlLFQfMoatwKansiSiF7RSYvDE8DJWrIpjIbHG
Gf7AKSpP4v6BkKh4pGjbpF7/VzIsCUDgZH3KH8fo7Oye8oyvHvQXcoeWXrBuIAfIQi0Whu38v2GX
/1vqLLa6AQlHb6BowKxsN3u5exPNE4IymVcEfol8A5xZobEuZEuCTFZYCixfw6CnYEZx7Mm9pb8y
G61O6Ws8KcevtpbfnWk0ufNH8la893o3qGkYK6y6j2FvSnQVnfokcBHewoMewoq+A6UlGmZ8r7zt
CSyRJe8s+fIPEIfYceAIRla+acQgBL8VZ+kKc9N0dnsZgwxdo1xkF3mA80PD1aHRtHO2Jl3ltszo
B3+04AppFUrzfU7X0glWSDu2LKMTPOQUZcZZtpmYt/VpmKIgLdPIwia1Vq1JRZeTM5nRMc9Jc/fM
HAca1Mw3j6m2lZ7OUbN14u46z0eu6agh+5abx39gT5uExx610Wp9Ipp8AoW0u3Hy686M2OxYo87U
dEzl00jZt5CdHAm50rd0hVZvbRhp8L0jppJCMHbnYh7vz+Bq9Ar9AboS71kUym4kroLoJiLwjqQt
fo2SionjbO/iBp1g/ugFLt1/wgRR2+vcJkjPUolEFaw+BR2qw+4/lTSCEpZ6zDZFj2WlWI/077Lp
2iWpk/eGt64hmBDWW9Gj7QtK/GB/BZlO2hM4lCEqzsnBQ1fYN0D7PtkPRlP9EHaHDuc7KOpoTUjT
yLUQrzU5YdIhzZ0wh4AyVA1Euk1J4KzrNVZeTq6sfAIg/IjHi0I1fjMKf+XB+zvvq6BKG3QxYXhY
VMVOA7LSjyfln4xSTk3ha2092Etd4awSFmAxnEpGNfs9ts+IogJTGsZiXUTVkcsSZqlO1U5uc61i
APO+c9dCaJq+WdFllWP9sDlxjMI+T6OWZKSyhvXOvRvlshSbmRGztBR5swic/iXjgpvFGsPm7MRu
hZqPAGnsiti+/NE6G9+okFMXeyORAQN4nvKWwwaphO79gOeebSBa+iwOwm4EbBqsQS1I/HjN6F2E
3WKYpgE5s+n0ENyD7DAPR30h9Rnn+R+bBnfmDkx5jtyZlvfl9e9cskla99LTLlMq7FXxD9Tgt9a3
4LhSsP7Lgt8EC3JDBsGVJqMiCWjmDX4psbmPXNkU4tXq7x6PR/4BS12yKvQwKpqzKlBWb3qPeqmn
5bOM+cRh6L5U0t8sUjOY9GBtDILHG3ua/7r1/lNeSz1p53SXfc9Bh83cpBSIFT0Nfz0lW21sN05m
DN2Jq09Og7OinqHTV2L50x9zCaR7zAT36L4pGhv/ntBitY8ObjnRR+GM98mRRXbMmkfPmFjmWU+K
zJawOtSTPD2zcG5RCrYOq1eKd7SWkynPql61sUBgEua0cgty5lhpzxVfwtghSXiNFYmgyQTeOrFO
Zg6DJruFRpsowEAlvm6zq2uOx1GEgGd6Tpd3w2vPCWEtK9W9vR6vu5uRQdia5QQ0VWVfXcKWpQEj
EQxEGi1P61i1WXdDiNe8cw7GJGsqqEU0of4X2D5M/AdoNRj3uBSSLOoU46v7gY36xLaqfIdfsdvv
2PMzvJXPONBdHKvOoCpNHJ/jUHPIsaFoKupP7LS2x10JUBvl3dcaGddS5LUFqMAV96C3Fh+vQsdD
h0kPyGeknzY9ncrWZt+UDu1zZr2UMl6ecYAm27kOvcA7eUFUgA9BaBU3CHffIQl038WHbn4Bw2d+
BI6atLIi84QAxMO97IE704Cs9EoLOkK+7nDFl/8iNZznY9H80ZUXjl7tUEUz3SLD+gxoAkLj5SA1
N691KOc7Gsf/hVwS5uSaJGZwD7qWvYoThbiqN6QrAGKHGuxYJIgAPGASzjlOt0oznf9zJq5rPbOj
Arr0on5A81evl647BcBSTP5+SvfDdZnkUqgfyTgv1O31RaHpVYaXXlIv2ajhVB6NBT4Qef/63aKQ
NoSbOsBvcb3tIndtNXUthT43DSrzyTkuYoR89eoxUDQkjbjC/8emporwXiI1IpxkG2cUBvP0unOI
GSnYQHgZj2CkvuTaLAT+zUleLx/dHKWo8l48MfUBt4Xl4QXOlr3RtT6LWuTWzRb5Ysbwuctl6ix9
rfpoW3n+cUwC+rJgIkbESLVwHvtiVP1hebKOMvJAhaMDuU8hsggZkjaqYf2CdMs4dHrUcwfNUkel
MxN2QblTbki9UdtmT3K6EXD7fhtOjwyMC0TUUR9fNQ7pEnApNTWYAa2ZBBtsgDUuG404jah28GAg
9q5/c72XcTzb61aBXfZJITHO5JGQp2Ctau2QK1ykkS239B73URB9Cd9WQ6SMMhK6cf+TR7JWUsW4
FsKOK1rHriVOA5RtE1zQLHCeFF6l+N3m3zHTb1HC33skWY5ReEhAswog/4b44N6ovlsWPrEg1ZiP
k1WM4KL6ASQJCII9BJ7zMmOYio/TreRXRcL6BrEpVivYGAmu7k+Tlr0RNyseWLPA/iJWyWNb8Pev
u+0CvTh9ssRXV1PTNnE+O3guOj9iZqREBVxf+NFQWKgvXq6ONXz2XoWit/IFwi2HFZzd+3eRh/yV
8v3UqY2kGYwrcZewpqiea71E0BedqnrzD/IX2A47njBaiJtbEEJiGj/LO2kw/fzS7bEJRlZXuDpZ
orsY4rntUaQTFnh+BCVXgskpZPOXtpnanKcfcGA9x7gX+sqF6tAQ0XA3qVETaBNsu8HuBeI5QhBV
10bUUXZ2js78A63+kgb7VZXYSkeQR5yOTVeTa2Ud0R0fj4kcY0u3F+I/PnsGdqHQzjFaTRy3cdZG
Am1cUc1GjJBwn84d4nXfoqgY+Fmr7j6rOcNCf3q9vblKcYpg9HxrLI9UpmV/hGyBfVKsG9vT3nxr
Jx3fNCw6DXiLZnLCvNDpldtKnZg0PFuOhB7xlvYBis1nUit4V0A/qec7Oj9vG5+WotvFLLhGVuR0
rio7a9VXiNbxUsuPEPONwLepkNeCFLdqCzz8Ym7wZ/VqBN22uF1hxysZMe99WBvMIhljx9yRuQMM
kn6Gw+ONSv+g9ZOtnu6MZRXhr1AAZvSNH+SkQgUSRVmOxRu8CEVfYHmaA5HENTlOV50Ar/tnOcB8
cKd5Hj7Kvdc8ABOG5IuBQecdQ6ddQrNOOFLpi2K7n3a5XJ2yauDUm70FDfZFTP49+lgLOPVmn2aD
ahVmugerz3/KJXR555XEZ4tnzu/E6ozZVysdTE2wDQ/nYNTERpOhBgCq83YLYgWfavSsGo1bfo9z
bUajnk6M6SvPQHSFH19DvDALobn2bm/UEJaomnPM5aaLf5BPpancikSnJ1i7luTUCi9PHMRq0J6w
fiRTcqFed5VIrZZTFcTgt6jJ1V6FP7jNdWGxjZcquvzhuQYkOhcEPHZBjdL/PF0/8qT6U3TimseO
mB5nnV1GACcqWf2mGYrm3WQzmZBKF4BvAglq0s4NyhyzZZOpMoB88esfCTvg+KeGFgrsraBQ46BH
WJRyUOsPCAuDKSAKai3mlthfV7NPeGJKFVg5fy0zF1mkbMG6SOiaEorLVKc0fvBsOKt2tEIlWUt0
0MG9uwxHsDHHbM0LX1e0zMOaOhWQQqWRnyPH8ZVRKsQwE0pvuxFJ3KkWAm2DZmJ4zHDjE90kgIdm
bf7+cglqginGqLugoK7lZ/deoapsSo/SKp2OQKJWRgChoHU4r5aO5rBTrtCTxtvOyO2HPgg3Dpq3
QPgifh8Jcyp2egfuJo4Q6OLpjH6z40hXIxxKAw/mMnSrEogBpDZ9eHVvoTIrY/UTKrgZCdb9ZQgY
HWGD1WMUdG41GLp+2xDQe+KF0lZ1lA/8hqovH+2/vuyMlsqQ9ewbBax7gpSa0odicyXpPX5J1ItG
7EXm+fSWKbOe9guBlVhkgVKQRopvZXYb74irW1Jg105l4HbOXK1wDsKzNw1aQc85WmqHokJrxz8G
Q+WsKAdBKSrTRc+5ckFyAIzcCLfLEVn2IerroTFnUZfbNvDMGCssq5YZW/wGfHbJCI3RfU9gFtMr
EXo+GseraArmvXPeguNuxSTXorZcVGogN/ZR/8g7OtSu0Z3omHaRiKelAKYfZ+2ISE4rFRBMhBw8
hiO8QfBgp/kxgYIRmiDJE2iONKI+9g8ahHmJS1164ljF1PHmxdK3TyjYCJN2lLnNQeliSx9kxSxc
8GIzQOgN8sLY1QWMhivPK7jMaqOiZW+1NHrlsL7Vv5rrIR92qbQy1+ExnhRANACHvVndGmZvSu3p
zm6LDlBq2TxNtAvGJCkR90IMy0YfCVI2my8MvUZYGXKOQZOL8G7klY8tjOEhn1+GCqnzmXecmQUD
cKDVrRl5judfyO/lIwdhYsfkmBTlUP06tvHdVeqAi9jP11uY9N/O9i6MPeYMaBzyHRBYmDXw2tY1
kAFTyeQVCKLQH03gYeio68/QpPPge9wveQQzJN1FWk064dv02+cwaPyHiEQIu13tLxcCwk/dhqAZ
5tY4px+a3bDIUvFFpnAiCySDojEtqpp90pYqlb14BZ1UUVjW3K7FG4Lk8dEoaWUK5VaiP4d+8jCK
RTlL/ztjXe66TaOiYtDEfF1Xt1RNfVZh3L/d/CKIXSUaL2Pd6JpzyEKoDIniH5JUolzKOk823ixp
YRbuNZMqd/fY75zwhnwRKkvxCFgwQjan9bVba/Z4lwc/XDcTdxAx3khDQZFb2WA3NNezV6mcByn0
o8cryP4nig1PRyeWTBkSX4TbbYL1QXr3z8RlncWSs4h6D3SfuV9Ot6cAv0FlIInSVzaarQ449Uhh
KFOrMFtiAto4pOMIFhBy2Ln9E/HARhbsZ9EtoS1YG8MQIdsubxIRCueIJQOP7avvOda7PYKbmREx
6A5C2BNcdk/s3yOX+fPqTB+W70MbrMoGXnbqGeldihiFoNbidrjpvkUM3ccBTfFDQm7XpNIIq/Bn
HgJN0g2pjJWrBwcoHMv8lvqOPEHvolfTLDpEvhg0az8Xd4or4uRFS/bQNmnfGUVJt5rZmSGUEj8V
eiImqAq5c3UJsjuwrqyN5YNvr1ge62Fdxe0UVfHFIO9i4QUq0171TfMHwjDEqLVMbBf7tQgT13Nh
dj8TEGPXI5rPU3JnPxepeK96hY+Aslk33UGBfskT+E+LzLmWDVJIK5yohhEg93FD6uFlshB71Uow
vWycQrQr7ItwWkBdgqzEww/yNo+IwIE67brSrC6gaPBgmrJzy6Mn7It9AiqpY7Zw4O7vjOn8MORL
ZJGGT0ekwzUCekL+xic22iAPL6zq0meBltQSBNwl8ci9JkcyS5P96XZ+nm7KnzUAG7DKj/KJMh/R
hdP5thgOJjK/GVOlhXRqYolFmw6Cgz7W29c/Zrp3gUn75xycR7qlOl4DgEctCZBBp8gvaLidvJ3R
LWXMsk6hRX3SI5GOIHLYWkqtUKS07aBWgR8R/dovx7TkuXf62BP92AS3UWHYw9gvhT3RIqlZhYXm
X+2q2jsorWW9nTjznabiEnJofbUX95WVuTAF0MzMAXTiAYOepLdnVu2V3LZCJEJg2lYmVommGhLN
iuGXwVvXfoz6frAdq7l3aaRPcJqZgqzFpcSz+FzVUdpN7K7k0rhWqHFn9DC+jONDgu9tZvBKIg3b
eQe6m4UXHEOk7uq/8iaWtk55ZWl2HJpqqsxmuwY0d22sFteef+f/lvzRPhrOqajhyflUudIt/Qa5
0SPqZUo1jRgz8muEI73ZlgBOufdJ/OvqvDHO3n+xzukK8FxaX+U5ZxCZu1kBAKsWE1ARArjtN6c1
Ochlf4kRB3DJ3QOW40ywz+eB6o1Lk9gVDYll/sHi3mrPa1yyjC0qftrnnmJ5B9QPzqnroPuYWoTg
F2DElhmJ4xNXIdq2lG40ka/YQ/mCcPFL3STyfAhrBC7quytB/3+UxWHFB1PrCPO3aXTCYQhCUUFk
YUnhsGXbAiRFRspNCCkax+lBM8niFE0tyOmETBrlJnglChPX67cyeYGk8bUcUBZYrUwy2vYahYGI
+NS7pJnP8v2IBL7m7BrATo1ovuF6ubT69w8dusxWjBfFDWbYTTLLftBGPkjP5pCZYuP3oiwXIXQa
PG4gCk60HKxIF+T5h+4LuSUB6984z1ikFuMKXJ7XL+7kAeSm2yDOObgnZQj6t7sQOC3/zjXO6sWf
Zeb1ig5VYTXsENIQ5Dv1kHQJWxkRE3E4tXPPFjNslVDP1HPSda9LYAEK4RRwUkMjacCQ2cgCMvna
3XHZHcrQPG8R4+AYu3ND1HLAP/QROsz49JMkiMW5NHqpl7iLf+ft6Y2H1yLEOw2ZmvqffwkQXt9s
FABqAMVJAlcg1NkfQEOqLGKgdu1fdjnNJcSaXhFjH6K03IrkAS/jzoGPtly/XbkMXI3pm0jnZ4Cy
2GldQL9W55yHLm+RXWEQJ9M3WNE3D9VLpwfR1egn5ebJvTf6pmGIPEbXDkeiRkDFeqX7nlN8VZLT
QDDcCzXh9iNjwWHekHgcfi1vq6vAKcCftFkK8gAigotaFw0LfJgC5d1efFDPbhblQb12Dl8wPgZD
hriSjM9v2J+VcSoUzZvyHfdGSFU1CuC9e9fIf3ITzZYDC0IxO2ubHex3Ep/YOt0Hjib8CNmkBX5o
HTc8d4PXFhWntvg4o0JD0qLPygbS+EziyNAl41XU0k602+CDYuIeN8XPzlPFi6b8+rQADs9xuI/y
hBHqQPs53g7+nBD4fTZ3+tO0VBwTNlHw26xDN7r7Z7Y4dtMok/r/9leYgywucC3TW6fEbCoxqj+l
3xaeCXctRWfpYTYwN0o0lS+b1N7Oq6qtPUX9LmQMs4UcFy4B9JCPrNjPYauiT5uOg3UMde9V6n+j
JmuD6IgoUBKfF99v7BYja6rDyDflI383MdXg24q7EIAGMHPUdzYPs+knkNYXIAS4/HVdsK1W5AiR
awi0MD1yZKxwjfVhZV4LQKJdYg9jMjbd+5kKeoK7yojWw1gZw+BNv1vngLTeXiBVN7GrVNsUTP3J
QUDM4Nzi5VxGLo8M9aBO53sTv3pef1nk+ksNNfy5QY2xd6ZmB+o/GxckSWxCJS4fv1L7+EFbSbyX
UnGAdeTTd+ljM6s14miOKGR1QVupuzKVt8CMgG2/n+U+a3ekV0D39nwAHdf7hwVqMkOjNtoNE9dD
r9rjxJz7ME5ksTx/6oJnOy8db0lOaKIqXzEKTf6doM7d4WrUwdDfKUj1GOcQsH03xCKLVxE4hk85
B4DUbrwrfCfghfCKSJkdBd+T2Pky6vgEk8LKGDDB53V0xsJ1TMFiE9riL2FIkXhRhWvl59sCm2uh
3eddhGAzAAkOLMpBJ3MsUgq2D2MYWHce8n3jU7H335EbLmUV5Wz/hGjXF7Q5jzmryu1Ok2asGD/j
6bYoG2IoYbW/OHe8ekmw/znWs+isq0+t7MrPETClrpa7f4vNy4fsnyERWp6Hp+uig/+qMbZWLTod
5u5EulSd15ax8HAmFMWm7x5vzxD/HqYCz1fyiiIryxk84nk4Bi+0u+jh/EybO0UfT1cD5EoCialW
lqXAK9G2MjR7Xi1Q3WcXHMWsRsFQZCo9J/QWoAwbqf5rCE0nC7ga4SmUI6IICD+KAZf7oZasYPN2
7x3Fy/ulMhuGH0TtGHeO5im+CBvmIx5BUhksZGzI+39yQgm+X0adly1RWngSg769g5G3OQYbEuo1
HIQIB0AkK3VgJtnybVoQi7/sEWCVWFT6m1YGTexGoASEdUiY8xrsuVN/XTBQNcPnpXnYkfFoe9io
lZrVt6Vf2KHJtK1INzOxzPP7p5JQ0Z4w8oNL1t50Q2HnZT6xsRxax6lO3TcPw9EUBulG7Sc337bs
aSDQQjO/B//5LlxQHLaJAPuYCT0muGmrgjkUlVI7/ZgLvJG6aIXTaheD4u/KZO6GLYPeDSO7GdGy
FoMhq1ulp9x/TcZlx2JQnKry2tR1PCYggHgnhNbyey47TymvJ9qyOkybSdhuDFAAqqy/bMQUz0uM
UHJ0d9SxHl5U1ohNTOa6aGAr4FnlEKARNMdGQwoMWNkiUknbpOMgb+gWrrUZKJk8fq0pXmcm1iR4
ZEy61toKURVKWWmDo+fM99d2e9GNYhEGSgmFsHDLI5UDuv1eoh1VQ5jvRw3LiHl949uwQa1luhPG
/G+4I4QwOIQLd0/4oMLQC4n9uN9XbChpIPwPRD0tohLYxGAaTQOF/jowLvc01gX9x2pj9X+IUqAE
BnnnJufjd13l4FF8FbTp8RUpxTDBeAre8BmtYOPsaLrS1xZEFcJllS1ixx1nHkx9phQYqb2huTcb
q+IAqqluH5GKDOKYARGAODcpi5f/0zivGOIVY1vl1RixIrKn5P3tiGffAL5DwsJ7MPv3m3St12g+
HKPHAwsGbzxq7kJdFReHD93yysYy2GBt2yU73Co5Z0RS6tYYs/xKMnNBE9qyuWYmpeSCCt4RQn32
1sl6aMIVYSQ9m5ZMxfgmcTM6hFsKbHr9Ctww4YsqU8JKmJNMNN2wfYMrl8qoKYlkodU0mg3QY0uC
SGQ/SGxcf8q8udBh8J0G5mTq5eOF2NFcq7gnXNvD3eLZAYjWs70rHy/f+rgG844wu4TxQj+pDO85
Of0zvzI5y+oxTSQ90JzhUoL9tjxffR3aZs/vbcZpy4JXgBsQ3jfAPONKJHm/cEKGNQCvec0GxLmL
+oB/OOxkDXXom0l6CBwxR8TajbMGzK1idefQ6e/w28WrNk0QUuLZdZ9xQ/pU7dK9v7/QojQlvdon
FuS7kFqTlKspwzxHqtA9KHbq7VxuxWOy0T0/KJ6kbrxiNXpyH53PqvHYgAwAfgV/Y4AicMmAyhLd
1FrtHjShnDol1d0HAUxPnzbT9xulwqWZOmLJ/AW1n9mK+yDYJJU4Y8Ao0avT3BzbF1AFDWihHieN
spZIUJesUFfOsifhmDpfISQy0ENOgKhp1iAehyb1rki8n0K+j2Fg6rxxp7fC+KQPYfy4GBcFwh0X
Fcdx5UahzzuoKDjVb4499bOo5Ai18kvGwfhPsjOWZNaMZsRR0CQLLTTusv1sNET6IAhO43EzKKUa
W96N0h3ii2TrYwbmgXvIC3luur/XWK7Rlg99cvhgO3adiUJq2OGdqwuFRQe7+hLdbnm1fBHFYB/v
9IZFcGIhZ8L7Xls8/lTcqiuzcjPGqioq0bCvhZBKvEulKJu6cJBAebFvunuXnV4T/MR0c1UJvtB7
7xwyuL1jDGFEceALnNvxkZWX1NQdk50SreK9v/IIopLV/91YTSvCK72Yldgt3a1TqYRAruMF0eTZ
tihmE99W6ZYK3st19lDLyHoAy9wSJ4i6NlzHctt9ag+Xp/wY/E8RZIDeBbpryA6NF7YVX0OnEYtR
Q+LpYtH87vp8m0UoQPIp7Yff1tDwiSKq6ND2CrVxW5ZuJ43KKZ66bt8aWdIlO0dgnGeAfZfZuRE5
P1ZxRW/FbO+PqV3DKehzV9vBy2yDK9H+0RBLmTDSVMi0GFx33iW8WN5KxZQrSrFcZsraDdBtbbNU
REtjAwu12a9U+KMCPEnOf3C3feA4Gbp6V22cvuLYtRvOSytYjPx+8bbPVAttZ2ejX5z426i2fJNP
a9MBZmqbKzjBxsp4dtCbjNm65kpw/txRiGTxGu2IaBWaV1WCI3Goxv0rvZyEHqESiv61POcS+gdd
jia7B8PUeOUzLbLrqM86HmhDhdOa1cHKJAx6t5OqwOVLX8TThxXpwhB8NWR/++aM5wYzp4TA8bb7
xuxXyYC23xFcGmtFg+l+fXcA8cNVC+5uYSuuFQImcBTvFCKrsaInta/SinIsopyrfsBcs1NS+7nn
zJqB5M0MonrCeyRP6vsVegfwOebX15in8OcrdywMlXw9/5qnQSSwEYYvzVQswrFARMl/HvH7tsIJ
W5i7cm/w9kwJyYHbrcnMkRmfIzEVTQgZ6eI9110Ft/1wo5F5sGzXYQQu+jRUsGnZRkxf3ikb1fDJ
wB9tRYcms3Mqfi1xHqOiz2xk6wGAWCxN2Qy50RzcoBcHX2wxkCo6/fSxK7xerA3k4m4o9p+fP1YH
AS3YI2cNAucKhQhpbkrPMe3LNBitav4mK8hUEYQMUm+pcWD+gDlT9tvjQJRMRq1xgADCXInt4iVl
hGRjl0357S1XSKPu1O0wsH5jf72jYoauPp3kY7hWeWkKlOIlwCdzEXnQ8FAWSw+sai0kUHJ5V3uM
gH9vV0q1QAjx41moLHpBkJSeUYYDbz/993wFjwqFva9cQCigPvO81specFV7lmdRIOnDbJQnVTlf
+RAPeyPm3yze45WW072muFsvl+mwB5Y4cU82rMDbZqG+/B85XHcUJyK3/j925JGsi05pzDbFpBX0
V30rPEGirWzeOhZIE0jYSI1NGpH6DYaXGBYtFRJJyeNfs7NUWhDMHuLJsQOeqF7uQ86aBD2UeFiV
BC+0KJy4rGstZR1mC2HsfSfS+tXgHLuuZRVbrwvBDvh8ytTkIrG1PP1cYB7id55Ru5brJTxcwnsQ
BL9TG3whTHICoMNsSPkuDXJOO8ozfCssnmquwqRaKVIIKpmChtfxCvtPnEuPyr/DubtO+cD6W9Dg
/GBf1429GmKrb5LhoPIOB9ra40JVkTX42xMF/+E6NCG70Fk6qcRqCXl1/ssbwam8UPWkT7ldlZDG
5TmWAzdOIXNkxi7yXkZSFIEXU/2vPpvqvnVT4zqJwek9v2fJmyluU5wUc74jw9nxrQ6o2B7IOdwP
ZvGC8F5OaNEGXSmAaTHPdCZ+Yc2HrpQKzUYfYWUnDpUhbT5ce/vB7RqlPOnM1cyFVEpvks+Lt5nE
JiJuyW58NP1C/mC60cmpM6yiNHxvx8bl4FVdya54CcI+rwc6vtBmynXzxmBsXlWJShADphQcvUgL
eerjBRULQBPjPw1fy23wcgMvSKTZLj/CLRL9yxeoNJLbPyNSrE350IPXP1CG3PYUPGouAAlbJYoZ
D1zXNMHQxWFhlLREJDjJKlmKNGegqQOGDcrDyocEz5ksMxaxiGXHoi/P2DlnMn7Tm/nObhUMxoMd
YJNxGngGt2MVIgHkJx82Z0MEd/heb+WzAM4I7Yw6JT5aHFarqmpKNxdMPZX3NX6GYJ5YrhFGc3zz
ySbI5CzFaECFGDSUhJLe/JoqDKjybfj84G49bnE+AKDGHgSHVQ1W2sU9FnXRn5lLXFhGiKfZB7b4
8lRQY8Dr5H/pK85DeiUVC6nbPTjsxe399VlkFf2SZj9xR0MdbjH7qKRHYZder9GYaCpPYdXG2a8N
/JpgIXOO+/mk8iq42JGsaxe7M3XNpX4RZTv14Y9E54c/b41gZt0wTwnb8C60CimCP6veZLF19BGs
Ne7EOHOEgjst6kBNvksACG/UXPHJjAqRmUtFRESFa5jxBWDQXsuoVbon3c+EW90v8UA2PGXlzdro
RvrNsH6KyNIj/f+dkpFV6cvOugqNjjlW5XxdjNM22Mqm9Yn0Bbb6K6p8bkd9efXFsWVtPPDkuK9z
UMbcqLpVfcK2fNbELn7ZBbmKKPtFkROJNp+kg+8UJdfYRLrg4JusaDBb/h19F3hgBGhQTCIhaG6o
EZPe91W5BZQdm6Hdzpz/6CIqQRGtLYzP1As39ESQAUZR9qCt0rkisK8FmlnqjAP+/BQGffvV7ydG
SStGMgsQfhhpQ88BzALSSNY6u/5HKPVKx78DNIaHuo/6Ty2JYC/9fd6BjdxkvHpjZ1WnmRLmstkq
2xk2zRBlkwxQAJGQ1lyk/oXLM5lnhnOT1RYeaMk1IfSv3xmTc2BfdV0TvRQHRcZLUVIMn6756kuz
NQJWwKBfcIQVKGdby7coM8Joz6XHRCElAuCK33VSjXMOBM4GKsrZ1Q3R8Y1MquQPA4oYV/vvUkp1
XaRvnpW9mQzE8ArrQefl5M/XHci/DsjDKxopDzR7grGBHKKzKOL4+Q9xBaFUngPIJUOmoB7uwtVP
p6W/qxiss6LV2x0pqxErgGYSUjBcFmyM7lVZcrpJSXsXcICtCI5ATIm2xZTo2pYkp/KwpMrT0UGj
bfd1k/+ptVa0WY7OnH4jjkxJxpD3/W+aXwWvcgG2eGZ8K2KucZgqDuDruNlSLJegqmk8VOAF0yMf
zuSLX7LkGlx8DTMZkH8gAYnRkNkyVKItaI18XYHl7ynEeU4G0N62x62R53MZcPgXcKxaETG5d9+v
hyHFfDCkRDFsDDauSwmSUIbCCMpKH5ZEEUyRZojLxqGGb/pzm4yRimMXqyVs6Gr0Z9ogfOVa3OV+
l82q7teiQcibOVlwsiNllVPrBlkRr9y8Mth8ubMoYEj+gyEva4oVfQQE/YyeQ5OqQL3aUrWdr4jY
7k0DvtVzjHa7NApMDa47N0B43Pse+y19Qsm48CHl5jPZAtzPc9AuKrq6Nh+9bp3VOsFM60lQ/+Si
en9+81KUbHMWiFvdB9lOPkC+QfI1PRqr/zl5vbcYvQEl2DBRp9sqv19WakdH4b6FSUjjAUB8TQyP
f7GsLtfBy6+r2bKSnj7MyBGKaa+KUy2InP1QjI5yQLc8duJthOgul+s3lvrJDw0sz0nbw0KUbkpJ
WRrsF+FpheonZQDuqEHHVqlUa6+z63kvR4k/xvXAjP3iXJVRQIN4Iz6hYMAVaEkCW16iNo8z2y0r
MQugSnt+KDUC4+u/Fh+WTs8ztcNjKi1pCm0Sl8+vBaN91/sbLWeqvFm+wUVwYzLin4IX5jNggw7M
ySOHl1kphTF8Rxz5GzdFrmrN10YflBaXSQDxAvnBVZHIs2mF1oFbfwe3RvWlZigp9ER7oBXuE7Sg
IjLNmpzLnAiB6NGdfzzZwLu/D2Z+ITwiTZK2bBLAvPcTe1pPg/y/NiYEIHu6vDvQF1TZz9Qf4civ
vU+idi3MJAHIwAFTr3qa3y6UqUSZauXq0/6TlyD3ZiNc/chZyuOtComo8qNUWqkmwYicPutjZFyQ
IH/c1Wheq1WpK9DO3XMKCQMuM+8T3749VRVQkGMH12ROS0N1d19e+fG36N/IS3MvmLNhif1ZE/t7
gww2IMPvplfGwcNDRVSorpmxXbEBL6Jr6GxPqBQTP5mJ89eZajTMyK4EaNJ3RjW3zWPV7pHENt8b
qLDEt05kQMs4Hr/6Qh4YiMDctEkcl7NRwR1nLnkr7uRHiy2z//NtkrDJFkdJhGMYlVTKuoafrHZN
290u3NgvFfZdron9SrdfKgg7Gr70/09gJJPhhL/+etkb1EYjR8ZjSt38sRrXMtKdQ6p/sayGv9iJ
XjwhDd7vIYXydQC2+aLI8xtfzK9K0neBXY90LY1YhtC5K8qkPAvLVf+RFuo21Vy3+tusamU0/Y+T
W6WUwXSpp3ks3Uoc/GOi7d86iBMpkHfR/81mzMaR+qt1EyhMRQP3pfDyZhWUR8nrNEd24kuoGpDL
Fc53kdMNVwIxMqtQRCaNV8WMypvizOZZlTi6uCZEIutl1Ca0huXeEy2edi3QI49Xr48VeVwff5vQ
MK8OJLBvbB7js6XvZldZ+DAAcwJXz76JgYxnWaJj17i+DL0Ic4BWJWCPFjM6uODNAgcOEptzMugN
y+XbYW/qRjAJ/JYezkBfgSZSbOV824++T2eoG4ekzDRD8bb90EMRbpKsj/qv1+ls5Q9lvYBtN7KX
8lVr8b0eCEWw+jdYR+ZNKSgSSOowvAUIy0GVYQTVg3KnBqmYpXE1nPZo93jDEGjoO5d9hMrck8M0
W8Ryc4cmQ+OK37VwWTAhSfGGSrs925LpWuWECnlM8T6Tl/bviVibFdrYoxWOm33TuflDq8G8tKec
nDFnE0uTXSYEJkoQOlxkc1Z3fZSaoq36CU/QtnKKkqMRoOEemiI0nAPZQ12E5xAKKgLxc7Cp6p2h
KrxPg6jOy5OybFC6jFn+GgAFu62Eli4n9BHMioWBta/9v84PgfSb2vEVnIxjf/1VJOGb6A77NecK
8P5keVHdeYMTmccLkwuiodpuF8RVFaVp9ccg/2r8kRcHzO7z4Rlz+DC4/rnVw8fMyWMm544opofC
uIo8W758sahPjd8IZqN6k/xQwL7PAzcRc4S5eO1EOzDoI8tHnllTaktVbLFPdhrU7DTo6Z94B+fZ
ZCvSnPOFK/Iy3hINQGfthqWEIvomphv6yN5Huu6bsfurpkBi6Pa6i2jxlc//xC6rojT9D5Tp47PF
QX0QBy3UyZ8MwVkvUA7w4tO3Knn9iENsUiau0mqa05RNDHDIBe70R3tj4h4qH91fv9VTCS6P92sq
nDzjAa7nKC0SeMxY+lWV0u+EW44Aas2t+1EBJyVjln2O20HjvSr3Wk6jdZeKY1WZNjqdBGAhy9u4
NRTDEiTKz/obIF/Zpdf6ahBNjaGmILD5ISENOzLYynasbgZ/1OerkYV9mhXcJBX0UEVvqT7guVKO
VmDzqNzaJ4N6SlnVW40n05z4v+TqX+PmTb/8hBEO6gml7v0XLRTE3XTI+mmnWU4iV4x/POBAKYNz
xqdaY3okbqtYX4R6x9NxQQlTPM/0fqw6JZnu+4CnwXY+XCk2cDWOsny+DnY26taFLqCfhipQEcIi
afRBq5zyknRgqNaGW+/LcWz31Hqcw6cLfGv4pCfecKPzNIqF+6wHUV/C6pGBgWh+VO/VC856NHnA
qtxhkLU44u9q4D6QIKR0bg5As4yD/WUy3OmAtgsOmKhQ/2c2CQR3ZYJy4mC3LC8KeJfoRKaSkqDA
lnY1ChetzMQQwQGm+PpQ/WC1cpgY7SEmRUTjA1j16IiiQzmKiAh97k2BzQCQ830Cv6ahFZM0WxJN
H/+aq8BmJ24ZNiPKM5Vbc0MbzoNSIV2CPFyQkoum1OsHreGCE2cbhhDJ6Epg00QHQRAAe6nAaYAx
GQ/aWU9y4ABrOiiv8NZTmV0OggCfZg7hKU4YmLX46drorVPcVOSnInv6NGMcGu8FQzUnB1f5ktc0
Xdaw7bazK4BMdfbu7dtbC5z09ca7dIIDz7bnob1PqYirDPwQSIH0sXAef9K+0jtDrEoFYEFFNbbt
Cwn3hS6hVxzBgD7cpb5VHkE937j3eUzpyEsov2yAIXw4RKoCkuOD/Bju7DgvNKy7DJoDEZx+EY0O
6xB9zgK73m0abBouCdcF8gi7096MDmyckPDIo/bFvNEEBULYF/fl3ndHbQThMs8L3Mu5RZj334ec
3in2ne/IUZryZJ1S+/5N4Hmb3TQZgI1aBK4m34K58jao9H/uQGDN29ugS7oPuQdVPRRnFJhl574m
/xGpqomKnihDR75okJKgWYpQ+h2wMlDXRHkJtkKyFRq/ZuEUC98avvuSsXoRTbnBc8uoLEZZ9Soc
yAFS/Aa1HWG/LdxWshNO49Gfv5QqtIfIln1SFZg/EqRM0LgJDKlrwJbAgYZdOctKkmV9xmH5nlNX
cGv6brAXLcP8dSryspTZtiJOIq641LTOrZ5GMonJWmXEv/v3drRpK+AfFIZVKLqS0DektJv+844I
7fcUEwJGRRgm8No/MWGcLsU0dKh6VfCK7nCiOkUBi4uDVkCAeKh7QW6OqNHOQHVzAUPubb+114o3
lDVmTUzjiwQWoMwNBNeeoHOh9i/CHjOAQhwyE40VZpn2GMYcfdmN8Whd+OVsvZrtI0uG7aWP1rDe
wT8pXi0FcItMlNbMDgkdAxisUHeU7W/seMh6Kmbn3fy3YzA1OtTDPkOUuMYAPmnThp5ny6bISgeY
eIXT9qSNi6T3Du++PZ5PGwnN/XUn5vzJuJ+KaL12xr61AKkA9/EN9YoT4kueDqS6XLpCY0wAaeYL
R+1nnPCV8zOKtVmy1Cv8nU9D6NJJOx5qOHGGmMhFR4RR76pEpn29x961+f2KnoEd+SkgJScO4B6X
KfCVkULNzVeFYrd5vVvPT0SzAOdXcAOL70u6HLmn5YxUQhjIp8eE9y0mbJ97M6QOtTLRGB71ukYF
IhyLixPYh54jWn9CoLUXhPyI/Dj/yW2Gzv5db16MU1zRYC0kimvogSatzH707T8nYxF3DEaMFu0T
b/MNnG14SrCNgaRfjWvPhGbwmE/wMuf22PJgsSroZU7JnlTBAEY+KYLV1PXfE1yq+iZuZ+g/UJ8S
h0sKuFmNARzRnj1lPWtqp4kNJ5leLinZlMFvh9/JJ8gz5V6UbkDzObC4uCd9faoG9Gc+27f6E2U7
lAkSi9oL3XXdT8Jsnd93+NpHhMKPZkzQH5UEOr//z8hFS5BMGoN5KureCuQHwlBDwecCzfnXnSkz
2+fTMEnDxa1Nd8zZijFXY9gllGLmWm9m6ybagwaYwU4LCC6ZMyGYIup/Wxs+qe/DDuv6dX1k60P3
BVUVqi7bDVY6tVuKFiKtTDKLyVQPQIi3CpQirEH/4GNJZVNVPG6wd+Tw9hqCsAynCrGVTvlJN37l
IVeJI0C5yCkGV4xmFdryC8E+D1DDzy2aWXIeyyjydwTCulrEtBmRie6ThA7F4RlCveGlvl3XDOxe
+ldFRl7Gf+VZ4tgA+3SlMKbTXvDGkrP/BsDnZdLG9sMckqDxNoNHVglZHmdDzf0yzNfA/sdNtp2c
f5i/bFCazlQPiQ2Fu+UvABhTLYs86RSCLVFzLlZXL3LLqlwonMFhD5SE1BhL5jR9BOIPJoro39qM
JftzAFAzkjaQtk5orXEJ5x286vPpUsJT2Am0lfmpq6SHyYo9BFX/IPin5xdQntrjgZ4uockcjfEH
Egp4qb3nS3uo1JAfERVwghHkaJtP3fgG2cbYth6y1ftkx+VnQyU02DI2h/PwIfVX43xAy0Ch8euX
FInOJt19+MUxG3EzD2dOQwCAWPrnmi+2RWx7D2XlTAskPd/qn/ztqpRTdIU+1/hIlnJFKB/QF/Vy
BnlVS9WJb15IWW1nFYJo8mpuTr3ZO/8LwzKwdHj0xHonVYAV7/98fdszw584Uzw7pNGpvtR/NsL6
nTaZvJC/WNYmkDxLh1Ko2sxrlduJK/9rw0dP6/ZizJ40bI1nrnFs3ZC1JLtSVnn2JS4wqerIk38A
KneZsW0GPqggVCNbLw/r7iELs72YpYrqpCXwD4mxFsIbi+MBEOe+sx80sK98NT71eoDN0ReqZfo0
qBiYoh6U1KqKq2dEXfHU1RvtBllQjPAr3OLS7uaG+hAGJN5slh62rNkcfn8ojqQWm3XlFH5iBJJg
e97xN5O/28y0jeWPGWrXTdRE+6tlxN3K0XtceW4OYj+Y//G0QL7tIsvvAsn1RUDRuSIDgkYyFL5k
U7yJK2sqHYfl0rZq8I8PszOY7BcjoRdtwRVfRtYMT/QqV/tK0HeMlOtzDMtnzjt1+NmZPl8BVpgO
rFDteX80OTP9D6E/6lBRtNRZXx4FqoP9BZGzjblEK8jJggI1pI7rTlv2/JH75r9ErTKhtM/BolL6
3BqAlbrPj1Q+dxrYYRPOoMSfZvGAraFZd+eG1ZnZFFCTeYxnYOopOL3DM6nJRXouV7pqAjkszjs5
1cvIn0jl874TkMuq03Tu15y4RTZtnGNMM336Xve1ZwYH/YGYgIsjDmswQOA2zAbcqlpHAErvqkBA
642q7IbTQngMHJ3dcwX1EuI92i6Ne1pWN7uDIiLPzMnXQv252bw+jctg45pVIie+G/BsRB8nz5SD
P05Pz+QTYedvkScdoIYZQjY0m8pmeRHvmNDJGCn+wvt2VBSdBn6slN0PLvSlomI8Fi2MfShw+L9s
pLe8+W1AqqJ/hYRI7sKPzwbwa0oachzHdRo/oP8aBonYI+qb/lTnPGkhkaOIuha32IHXPTiBrt/q
vQa+l/F5xAgz5mo4vRJBhKTM06EPGlv8JGws2l3LKoDQCulK+y0cGQb+k7HbNZpoUzyw7voAgZdR
onjtXIVNnsLfJGrcpqD9rsVdfOfsDpzyj2mq0Qmi5dOUtDxkfQWYiGea2ioi/bwrKUQYXY/LOzXW
J1dRLFVS9f67PZyNUHA1mI4gyge1Ldydpp6oW5jNJSVqcIU2/MiRLHrfu+taIXlMGThsc23HEnQL
k0oQgSdmgTDaXHU+RoLdcsP0jnkJ120OPEe/WQnhIq3Db5SIUkmeoLWMoXhjNqYyECvCuSL8EFnM
LnkNuow+q67xqWJoFA0peViOmeLOIsDUMPd8yZ7CpSiQytNubkY9xWWQ+r2gU39XNFpJloorzndQ
tVOLBTN0F2b9I71WWvouiZywF9xvHvQsbJ40422+AE3Xz5lZm4Z3TQBeGLdUNHPcA2imsc0SyP5S
6LXKuVi2q6MoW8GI+FDjfWzmNxERZHqliFqgktfPwa2BLTcIg6DTILGwQWWTD3zZXRMJ8m1saTCP
Ysi3YmX+UnTEE4GuLLLrPm0ScNlAqNg6l4rPxc8acSr20T1CYKUPorKCbJsTsthdHBUWAWYj9dkV
zmFHf1PxYSWx3QCTcO9Bp3wdbTbnzLUig5g8Jy4Puu8Z9jKmvlWCcEG+zBMiUJNtMbDPUbj9aQGF
o6cwC9+omFIQa1ooJfx/wpWHs0W2qcdqA4S9G1fu0mFc4Vc4yw6ZIrd3VirUjJEMOHxNZp7/sBii
eb1JzDCXqK0jLLSmU/T0WrkHxJEtH9UDZsm/sXHkjATVcZAJBkyTf6+fuWh3MCVTza/MPwf8kiDG
InHNkiYn05WLHrPMvDggdvXdB9fFlmKIsgrcFqfCInkJDqN9cB+fvIWsvnw7ueHH6Vv+SHjBFFLC
2dK5AFIDVtR1nhG4btRn2O54RwBUQ/d6L7Jgg1SiNR6a7AEtTBqYFsMLBo+N0xqEHAWOTXWQTx2d
z+2hQdFZWwxyEy1QNnkoud0UkyA4poFByh7jWCEED7tv70gq6J+SQEUBd5juIQj9O+7ncK1PuGrc
itCCVTG2Hod6FDrHAAOOm8ze4/dqtX5Chjuz9szsUNSEWjw0dc8dQyngq/SxlCl1TmOR5ojaktmY
aFHT/Pf5hZ93D1th2Uhu11Go6NF/iGUouc5ByXWuNAyjsfbIWyDJwMMfZilMEhsketPXHIJIA52T
4ruZVZhxnOtmm+Klsf6iw93Sr/lzLcP28U1Qy5qXAd+MnEXlCwPDwmuLjCz/OVs0l3xEhcHzN+fV
xkyLi8jtcaM1wdXINtQ+r8wdnQNm4TJLnoyjX4E0C6PXOtiB7cwHHVu+Zd21bgHD/+H0bz7BGMAu
4j5EfSh0LIxb/oMmZxLBa89do/dTkxB7Bw4UQVJJxg/mzbGe6XkdZ5uofOrrJYLrSVXIKRT/0T0f
OWHKRK14vW4/fGUxnnmV+xnTI5LogBe9CCtvA++5FOh4t6tZ76UHiNq2uCuPXQWe/bob9TNFWUhD
IA+KMElkxzAWrTL1nuE7NE5HwA47hhqZ99GEDVDUYOsRpwz9oril4l1hFbXzqh7Zlln2JFGlG+Na
rYioLlpk9uO2/mTdvGQ31JcopEgX1jPeK+MZ7lkYCqSvrbRpoulkLKDqC2UK2sHgDztHdbcCWJJO
+wzpIf749CJAcKY8c0IpebUG0bK7tvRb15oQZeOWz5+fl5tww57m+IImeFCw4xwGhGw1Vstcb8wR
H4gcchkNLjD6vZSGQIYTR2b0i5n41pn1ifpcFU/HLAIzKpbtTT2kEQGIxWlfuNLdFcXX0KRnsoxL
cTzVPyD3/eN+ewlhhWnyKjvoqkhWjznJY7b0JIvlJpbbl6V/+X9xcT53exfsHzkMqrnjgaQIRY4c
Cu+aTD/g/192fp/GFyDlwGWyXy8YtL/0RFJoJ3k9HU5i4DX6gNMMy1PHLQhVUHJq91DJjVGH5w0S
I1TMhlhZTKFfLZv4lNbhl+8hX+bOqfxbRtsSXUDozgEYRtXjOuz0urbJZhSNaJShiNQpI+CSN41X
DSHoykC1ZCWY7/nqPNXt5IFquhqjMA8l9fCq1xFc/yBa6n9IbKyuwKRHc8pGARGKrFj5fVulfTit
lnT6hixdNtxRYnXQbRM268+9cXvYQ7XzGxPDVrnn+WURyuF6myL+mUU+PEkn/ZVE1zzI2R8ZSreG
pYDXiBWaj+k0wykIsDi6k/7MriVLpVkf0LCbPFrFP5qOvwaWM6CFdiLaXXtLpeVi42cvkJPNKa5c
RlPkHIUrFlOIaDdNviNszuOAYPtu2KWmg8mcbixlaJpHRxOZSn+agemH6dEMWs7Xk4apBSUfV1/F
QnybhnoWQwxJ5HesEmdiFKzOI/pNvW6juFhGUmVstrQxDyWzzpp77LhRNpKPcc/8lO2NX6Jm2AV2
IRTS5uSDTfOnY/NBtIkaZOTyEdjnjTdUVmxUekgi/KIZtBZDCBNEHJkEf6UNR4hofBwAh15hnpJp
hvnWvArXGH7ozwsPAX7M4VuenesM1wvhEA5MXhQii/+wgmhOeecB1kO1zVehJZTZk49hmNdx33EB
15O638/gTObLYzfLqFfKlfTQJFerb3sCd4B6mb7b9dK3maqIcrbOPUFPE1Yk53WQpI2DB0S9B5AB
alix5I3/yCJwZX/J7WPumocieKbm3pvRoyGRKww2CzZCPblAKfIAdwJGeH/7aGy8UgfLiLErRegW
mdsUq1pDS+XOGZOrExZ/bxy/ahYgA48VnWPW0tKd05hNDZ5891PmKe6+TfiEIJrmwl3C8fy+X6aJ
23ItKO0WC/8mT2G489hH0zF0L/XqcE9SjcKaNR31ah7kaCv7j2UfWcEbkGHCNSP7+0nR/qSpbgQT
+5BstV2J3rl2C1sDkZyhZ6MkRgzvyQ/6mueI/uDzUwdtNZpo6KxGvOwQRcFn6QqvxpIzYuVGhedi
0ZfTu0USTvcPCaFdNaN3ZRYjdtUosFrsKYodo6AQ56sN8Otf2On4DIjxN6yo72TpW7PtLMM0cVEN
qyaTtLbbhOQUeTH2vswFr+eT4hHtTqFuBvCykBv1d18sqHInypK6h+ZTPQHZ/QA8YXnOS7U96671
PZ6OHaiXHMBFaGAkz4c7dQbym7ZrLXzvzq9dYcwr1du6SVRPvybLW0e6mR+/Fwa0kYciIKGyCo/l
4dVj9gsPf43719NtuaLWHOTk3ZtECUJjPUOxr7tPI/uyr+z+iiwfmUyLVlVchu58bmqQjg0Ce6ul
JZmqruhMl3k+xX9iFpHh4KrcV3TU3t0K9ZbpT0U1VJsBC7hjY0E0k5DeqRnfWNqythkeIpndUp7b
P1w4ipwcy7g5J6wT4Mwv+REVav586rG5n69kkKtNpNH3cWqxGwOmKSrcpb28ZjpL6KevGt7z4iro
pU7qMWfupetV9NOmrxzYGtB7s8V4XmEng2BLosvhY3A994V2VVIXf6+tSrxjMPLiZV7nVapGhPZz
Nl5PhihbvZbYFHKPM8ilJR7AJjGYWSBoHV5wnu6EoroOFmZ3ds9oJVIY89GUDy7E7rO6P2axZjYN
XhxOwDJIy1Ou0lDj0tfr1UCgk2vwvudD1H6/u35K+1WcGxAeUGWTuQtDjQLXW03xxZIMJ/QC9XBF
32v6S4WaPt3+Jg4K5BhPqg/v8/F96KJtnxbP8zk13w20Z7am+TUL4tEy7KYpwPpHlBzoJ/AeB8X+
QqfxB+k7v1uqiBLkdPGph+6sCB18q0G2eV2x3rHRmPEw18labDiwbfJdHQn2aeh0voLJhLWQVr6y
6G4TqNPmDFzLDgNnxNKZgpkwbObfBQ92jqKAcwRqOwAwE8xK2akaP1pNqPS9hq+d0ExKfDBWit03
oYEmQd8BWZWD/RVx4zNTgnWQIo044EUEX/OMNO+L19/akMfh8MoeuMyZJ6+dfRXjMUUaz5SpaK0J
FBIo/RhvCPgyf58V/U197pa2eOCzXmuSIQe/Ts2K9lSG4sQ2+xcua4SLoBtm1GS+ufTyoed3X5HR
MmGwfDOG+YD/smU/r0rsZKk/24hsjgEGLmIML7o58GDlqcLolIOp1pdmuMd2dYRQ/kWq35OiZyie
M4WGrx57CuEDEBARym8KXoLI6gbOrzbSX0El58RxsqOB7VPCoZzRNSZSYPnsueliBWm/8F5StxQ3
6gxEE+sYJByZE/ttZXIvznrc2pP7FGQU++zHkIqMRvS6vP0yTOHi39dgM0Qb5ftq4iB3GbkRevTb
5u442Hj1jGhRSIljUtjCryZIorI2Y3zlKZ47Aru5Ix5Tr9obDcnYGUWHGGYjXB4m0P4xuA0yg4o8
3WVoYSRM9oSjaRiv6Yy1x2SWnUvMMZ97a0wvm4f9Gv73zM9b/SypjdOIOfYPYuPUvkCrmnhoiLmo
lQ7eJuWWX2Bb0fyT+y1agIK8pevgwTjmK80uHggH+GFXkLAdA08eeFx7tDPk3jYQWlUtbqD65vq/
jieoffoHE5KhBbGxC91inBmZ1rMsVtX7k/XZ/3ua2zQHJ+XGqoakKaPFQ7ZRlPCmZmA5kBh9MqlL
ErsykY1bK3n/TPWW339nlnYTC9FLoE5+31nqOZHkB3ZHR0HDqoW5Yd7/FXzJhTzWEQsksahPHOkp
S2akDpRZVsrxtw22Kj2inhUnpTXdgWGkNtSZIacYzv5kFoChL2MjOlXJ/II4/kraCy8fKOg3YEae
K7Uo1g20S233aNx+NS28tS9+XHl4GxQKECs8HBXiNGrvAplStq+htCFZAWKwlf/I7QGDf5bOntKX
zKDdABn0NMbWVSFONItkjks+CZmcJwii5ibo6tB+M/HEhgfPfsWST9lh1gQ5XmCpA9Upc0RIOc6Y
fTkolLELumkQyKWSJejIm1MxfFOh/Fk5Er+WcAspzHR4CNOVnITmZWj+vCXu4azcaOThqxplz5KI
7O+UxfBvW3Q/X0tDsFERzoRH3RnDb9E/gl1qPe5AL66XeoAfT0Fj8B0GcKOkH6NfhywVWc7iSED7
0zsUIgEh9LX35/0NvjqBavL9VQiXY2NiRyWJSCWL1V762mzyN2i9FDoOjHo0jo/lsW4HFL9AZqiD
GaQ/xmIYyHZVKEJhOFxy7Tm3cYlfzOXWZVVoBZbo6FZxnsmBsXM6g15DiEJr6n3wxyQQYrc4Lbo2
Bat/h0SN12Zf7VVO+TEJYEIVqtuSlxCixkyJx08rRAv5icLvc/d9ejtz6xwgPbvrvDmH5/0R7hDC
vSKskMkzAs5dEY9h1La+xnN8+0bhTw01K3jkTk2r4laDRCoVHh98oQe1Y7Fh/Vawh568y1t9+/IO
9UD0cWeXZHZrKILpsItmFdJ4tsEShnKyvc+xWqSeBKKY7bYA1g6eSR+iKkEK7HVnmpjlSca8Mvis
MPEvMXiQPf3V/w3gJ1AOhMeg0xW00AEMYuzaJGvhPcsG9uPDojU/MBRidwIfc+ZDnANEKlPIbLMk
tCXrWnzsgMRLhGQH9S1rjtJycyOrPbOUvd1SiYKKYY8rHhG9HwEqaDweByDayvdvc7uzFZthaJ4a
tEyxey927Wxx+sLq9b+0Tsjo9f8185cGtTs8LpE3eJ1mz0giixy6gxzQHps7veSJxvsOE6/rXGy4
UPa18Go/ziRy27bvatgA7Zwj/P/mHLXVkp0J5qOSS/IlRyu1S+HkgyyxivRrQRudhoOeF20wf7tS
zKFExZvKRxCcevGpXFnL+bGucaC3EQ/v8nFYUx4/SzNqOKkuAu0y2QJq/6z0oCYWc5SIZ/zpFwU8
SqKSxnng31UPJbAhtDulUjY45p2wFsTpVv8p6cJO8sTtqsFCsYFcj97PIidxM29yRQplg/sgREPP
6hbgWCZaxb3lfs6X2LCNCcIxFVBDOLRtF79V/jAT0plavdirUplrju8B95vkcZnmNKZ7A1RVzajf
Od5VDcK6MDMgq+xjAf2CF7d7/Fj7N9QXPa/r1bTaYchi1xDYfSq5eKoff+rT3yEwD9Fym2gTQeJ8
1bP+1RgtJ9byZZ4y5zE2RnQrWId1+4foRmnUacpox18Jn8hbl5QJ2y1Zi9yUUo5x8yqy/7u7fuB9
VrKv+LueugWS8e5FlcSqY110cy4UJpszlTKsl5s2or3IMBbyx9OSTer+iPckK+0hodadhPmEACmP
ETzCzKNzapbt0Wyju48+i3eXpW6RlzivKkvWIZEv1h6P0c5GRlqW2wnRZ8yB6p6gEd/56HyhREK9
cvLeo1dAZ/7nEx1P3EJheK7HJvynGwwEsSOJoy1XAmu8P/5VDcxKURtOHW29Jvnrw3oqztxzAKMJ
4HtoEBKR/THZKFCrc4E+me1KlCVddfHLo0elvzlH6PXttRcxZWQC+FiIEsn5BO0B6YcZjMFJbGHm
xCb9xtTXBW1T4KLfAP7gbczBcrlJOgQLWnz0RT9L14ZVaWz+swKUXenFxvXwoVG10+HKweiwRJM7
SfPv+VklTqsX0sz5X9Ra4y6AvRnYKmKtm+p/IhUlx97n4AhGC2payhzUNZmN4Yk3Pe5uCw40MgQb
DlIKwwK3iwOm0o5DWV8dLmreN74eavcLIeuWx83uEJIyTRyHgWrwv60I8ijecmga53v1zL3W3bRv
Mwuq01mxAeGpil5+RJayE1c4sirREBuBylX00JPYQvWgh2JB842uoRMfgj/mp/2vDXxyzRYOoWkb
PT2A26N7TRcNpmfi6Vk2xWaPdKopFzdujvvn7iNYSXSUuNfvTKb5WUHK015exr+0ijGvH1y20Gtt
8conjpguxda1VpHYMSz2OX/Ytqaa77Vj/cTIJvomG9X8MtLM+sQNuWJXF6knRSvty1V8+byNN/D2
bzHiK2XGU4TDDYo+altrTo8qbomJjDwfbs+Uj8C/P4eCjmxKljfpXz1GnbVEMBqf7cSBm4WkPlkf
XvJ7SG/lsXS6b5e2mGWTBnZDJnaWiy8gffk8G4HwJ5KaMHdxo6AwSBhXZB8NGxE9a+k1RB0hrfNG
oJL+tCfarhnov2j78yYLIBWgWiPnbdVnIacLgFeENw2wjV3a9CLanNT/PbACryJiF1X2yE9rIccf
+U9TCs7YAZ7WmZzPL8vfv+VFAQum7ur7y298wDLVLDR3m5Zm8tPN+7uNQHaBDtqVF5fK7Zdcky64
CBkDsbh41dPXJKd4TIGAokyyms45fmWNbkIBCYm/gmU2AWvxXKUETAukPSA4HTZMwl/FgkwP/3Ce
cfWtdJvitEy1fxUreCpiJbsF/QdMSK7iBZTXDyuCQBia7lsHsPMhFSqz1CnXLx6tIyLknjkAGSRr
179GJkKNh8l1Wc3il2zFMa0wyI7XwC4140XGJG1rNEIweolsf9pzGYKgjZaVqjxuj64dEyozja/C
lzmXgLpc3viiIspP6DaLzyznFiBt2073TMnDM9HMlIu+LUYmMt9TdxshCOH0cMeNsOgecaHWGvBt
J6/+p69saO/cloclyqK1+QV17AuAA2+d577BMiNS1zrToUNhUGenYmW8qlb1YqqS30ulTermnY3w
UFy1YsyJSTiRtNF1hIIoHpg057tC54nxTZACHfkJuFl7BZgFYRX77Sv3b0g6WF5gi6vpWlfVLq1W
v5lD7ZzqsKC6LUDSnqO8iZ70CoBEzs5AHZrhre3yT91PGwBlsetYfegXthjKesOFVNuaJUHsTVrc
2nSqH44uJU8021gvKEilEw9+sHZpK2+eq9ORmex3e+dP+eHXndwtbbbUI7QuM8gKlAf7nHr+yVSH
Cq1V7D2deXqxbhCxOp2Z5vw3bhOGxzWWNHg1iLLI+Dd62fvhEckHrl7jrM967WdQIrn2HIBF9VYc
Tq376p0/oFu0YLj7f5Q1USUR4wiQYllk0+MNOI7eWoX76zQ69BGcjbp0oEutb1ibFKvLFGXddCvv
fzdfipVgg3MmP8N3Nhon9sfXJSNFIY2+AV/nA7DxE1TznxjgSAxWo/4upHQSTXShiKi99Zv/tZqX
FitJatSUVWGdMc0OiW2Urs5NHaQMoLM6nYe1GKtW1m3ZFJYES1YTJ88/m7jqLIdp+Q6aT/s2nQlb
R81lglr+S5TWBen6ymTou6oWRMDK76W3LETpOl9iejWft6vp1u6+sntd1vsjISbWybB5dvcx8u3Z
YoGLC+F4kHlHS2DGMi288bqG+vT7u8UEEFzf5X1tuTBmA4+JRRCgYoCDoLcZh0NQNBbfyP9stKJn
2wt/fGGD8riFUOqHIxfu/RhEbSDwrPYqwlVKhZixDXCOZ8amKg/G0PmbKQ9d+mVjQsHnvRZzuy4a
gT+AONbn3cL8N/JsbNvKjgHpuQyvim/n0H4LhQmUzgUqaUlEq7GNAEQY79Vj2OYNH5rt8pHZbSqK
4JWmFSJx/CTHeuQ3PkN5oqYY9wn46SqoR94sgo72rNmGCoMp75riWOCN37FsXx9azY3RzNfRVXPS
AZh9fOA/Q0TFvGbmwVVVYdLyp2TEPclosKJ8MpXBOHQ0Sv7Ddqbfd53SB1/wThT7ogWKZCtDwehG
zTQdRkg1tA/ZaxtYKOvmUlUFbAwUagsAVIFJrn7p7rPnbfaZKM3ccMba/3lhe2ovC0eAQmqc0KB0
oep308JmFrZgZ+JRKlD/EH0RkMT4G8a//OaIp8OjK+mpAs9FsO/5+Jlxbb0OFczQy4D2Jj04MzQA
qTDTRrl4Ki/+kq8tWVKIqeD9SWBHs4ACjtrnHMUZWcha6cv3A0oqkN4XNdqYDrlK29bKvsHCJzC6
2zb+seK/h52zOgjt9P9JX81gs5EYJhoEu0yu+DpzI+Fr0vSbR0NQipVgamppsKbsyvsKN/sMHIz/
G3a+q8NVVs8AhB+vzkU/4KUtyC7cFsy2A4SyMzEEPg97p7vvzMxWEz9la+6AUuoDRfrhF2RfUFea
1Ql9zskxyWgakUAUyYgALi16QD6w8S4bm/PO2uHt9gUeCJckl5jl15+XPVkqNGGrz8N6kAMBVKLl
UeclwIXuryTSNZ9le8P3grfnbAB3FUCgqHyqQw133y7v0P1CNPr+QnQHXQNX6s3CEofuoIKJOPEB
+X9vyl3Ts5KPfqL0ZydQNhINEFoC7nv9IIT6dXn8ig9pXv31+hxVDcyjDC4HfS4JD/l/Cane1qiM
FAlD9JrkutYgJkKVFlwNhApTodq/ebqaGKmvn81mjFighkuiac3pJE6XtjzkMgBh10rb2tyiIzbg
6bmVNXKyh3diYyhDar/jWyNms97TDThYIzDD83UrB5wgtRC2u+5/c0yzlSO34w8KJOXj4ckr4V6s
gcxLF2JoaBOW29K3chMmiQtCtf6ularJLFfLavdW+7Cb92Yn1XcEWdFgPMjBNUPLnzBMMOGwvhCg
YIn4PwYDLQZFLUhCQgdqiRyS0+hPwwN4BbedqOZWd85wlUUF8EYdl9GdoKoR7sKYuW+f1tndJTh6
PtqwwI7rp54aU2IHAokatkOQbDf26jA3EeXrmXlKv5PKMpEPcukveq7ICgvupupOUhOp9pt9kLUQ
KhXQFxiRVH1i8pJWhJwW7L9yB5raJ8yaZjC5NryqSbGtlIiirUaatS3VoQ9oisIoNYEyV2GFku9s
BnHg+Rr5XmxVSCVK2ZHemNnjSa5qzAepH7iC3u8EbTMguzpiYNc79zMpCXkHHZ6ExmgwrfZ7oybN
kJS3ptAo1Bu3sWZey0Hi5HSm+mc25x8EzwTEYlNeXU4b+VhqOzmTo8NReLHOiDiyLWsJn1aU4Z5o
Tq3IU0OPfGu0gFm9aIO0SemotGaacv7EoM9ljVrUsDgIdwIM3+nvrdAFuVWPRvTtD0P3u+4ZlRGb
+O3b5FCk4fZySfbVplHbRZq9Hk//uVbUj9IT6acGkuSgt1mx08/svBZ8niTiExxMw/EZNyXCkdZE
ih7jK0175POa7jQ1qLE8k+9mo8xSAtmaRoKdfe7iyUSKO4Lhn4RE4NFWDxTek4/JeL9Wk6IMBsAE
feOV/y3LTyILkdJC7GYypW1JleBukOum9GzRqAowDV35PKSih7u3tO4SB0gLWgK1x9oJujGEgJxW
BFR37z5oZWf/JYo3nCEMwknLDWvpOqkVfrZ51RkwuQauSwvDxLMQ3xtcje8sGdxPwJZ+ltArxQOn
3aOw6CFwdVey2WZC2nBGgh0OJQ/vVgMvGvyBZsG14dp+x2T7gW4AKPvdprua6iEKBoTaoqfdcFTe
jGquBviEhLHMKwTR/6aBA5NZtePVG0KAUVA7/a9dYhRjqCW7FAL0LXP+HfTBMGteV2WOTwUj4GCh
7pmox3+f38k/iWQRFtr86phRNhtCBetjDXNv2NujbNywg3UH7xHdzDMiIJkPhpxSZyhkqVChKJGQ
LiL8FQdZpWJEkwdMsi3+JexETPLY0vZxLHN7hFI9yQiurJnelVkDslryQqS4q9ML3i16rB8BI/nf
eoU0z70CL0Z0cLIyAeOiHn9GNq92d1QEsvwPtvQEcmGuoSvAEDbdYPibRJEksWPLwkmZ0axyqxN/
RpI/9WeZH/9lvtPGdkljlWnf6lkHjvE8wNW8jzsTI7gOR+N+aAvqAHWxUK9LUsgUa1ur+H8KZp6u
igQI5+kHe51ptC21fxPYTgxj2uTUpGluWRYcaWuyhDtNrrvCrc2v7t6RqTG3Ze2U6hYVn4Ae/g+6
JGfCdAQvJp+rht9JrzhsPN5b0QiHEflA/FL2frdm1XEUonVH3BGM8m3rPME2AtWDkmh+F+XAQqRx
8cDcTdod9i32f/Qh7ZpLdpR7kG70vOSgM/YYg9i/a9wGKAaj4mdcnHaaDpaYQC8sVj3TLmHHrK1V
oo9dMdy2tmhiBRWGMD38EVbOXKsHcDaicUpV9TzS4sLwITh5sFojtKUrT2u3l/eeGKjHf3ujuXSo
azx9fyhD8q+VZGwAo+O6NILF568EoyrPrwngbnVVCOz7AT3wFVkK75UvuJMU9WIXh/6MECw2KfQF
hyyS9VTa4k/5CHMtaq1Ob8sWhsF6FfwK2ovP1K+qP/2Nbmbs7qfOUs/DgRRruQiT4jK/14W2HNGs
xK+NoFBbW1wbLetQGqpUC4yLtKmhf5Y35aRBI8UZwsKf2fWk4qLXhfOUBzE00x7N0M5e30GaYxUs
YLYA+Z8FOSEKi3YnoJJcxXwQFC3m9zSBPT6JJfgP915g8J6BhEopWyV2dwbS2EVB0Ex0ZCgi7IJ0
/eXOZuPvO7mGznFaKbOyJLVJMCYiu6oBWWEj1I8ELgnzS/EgWNcM/w9pQCeaLF7dVE/GGqR6PimH
7bymLaKKDOngu54CGLHhNeQkQq0MVN+M0wDtDQ0nIlemV0Egzc/xsMqal5jP7R+CRgiaHdq1EfOl
ffSm6cb1ugMlFGEFRS91paOFOb6JE4sqLxAg1JPIjxO249UCC+YA81kowk6JM1G9oVeXNb2CUbiC
XRBmPsfxU7O0y9DHOwgpgjtc5feDoqjtDJ2OYvDgEPkUX26U2LpyIEVJaJRJMqIdDb/Mc3Zr/CGr
V/m+u2mWSeU4QA+F3gCRas3O5N+92bvflr2fqHE5tswiFC+uVJ0jvC8e+Sz6Q0TIZ6gcIeCKIhBt
OFePJ3UopI01aQxifdYoPmuT3ntFKWZrRz7i3TLNTQ1TcHDTDLIFCVullrVVJoYgH9JUYGxjyMeZ
LuJCkVDKybPIKNzkTkcKBBKZUPNRxb3hTUjLi5SGoxzgmJHSrRRKhosu9QkOK/oD5dcw9XTF7h2Z
TeDlSZMuS6tBCyF+8Nm07tLSfM9FiN0uS4exxnV5Yi8vndLhl+nmrklwdbI5z+JqUBepu1vZzrt9
Zh7T4l+tUY7f8jlI0lhm4PCNLQkiF02NVJ9kb2MuLWBEprV/CCF/HM0g1x/7L//aL5nwkCNMgcTs
jgLkxY/GN/7du2IAY1L3t/Wpdu5eN01umxFWAj6+O7v6kdcqUyp8qF0w1to+iNyT1u0p+QiWRxgF
lBDkjSz9tMPGulPGFCs66gklUP09FY3lLde/qeK59eD73g/khmr8iyqTor4Tgaa79Gn6Nl4Nqsje
60OlmIkWCkxxw+uqn4zklnBlAuiZQTaplT5CZvtctU1fGoMXQegsiKqOW5Pw2qgv8SfUWjwCods4
liUViAslPiZM1QXpXQjmbNoEdbIEuyIUbP3eH7lTeosnVybMoG1sZOJ8a5JIfU51ZJ5EjLpGzZ7Z
J78lrPODp+Hq1ZZfTiYqnLbRrcUvnhJnPVWofHMMFbHMJWhf9QCGviuxcEUulJsp392ibruI5550
cqRM2RUHZiIhdr5JHG+t290PE9fuIz3fuwNKXyPFs+BMBw0NfGcntVB5heWIPVloJqfkQj5BJeRw
DfvfJFq0qzfDVif7kXoPfNSouBLjVrJ0BEJSrfYaA2WTRW9qdqebdOHB4t9MT0FD1NN0QisV/nFS
gEUEbCRXZDgioXRxVrQXBq8qD0gOij4Kxe56Ehqw823ST5zkRk/9VOhEIaMoy8AkLms6xTquO+qO
LF3Cs0SV5UD6H4Vdi2LRsPd2hj31RiI1nQD9H/NsLBNrdpa2Yt5sJqZp4EidLJNHdEwI3XSIGFsp
e5iVSd0ls4HYAQM/qaaqN1tHu4NurIg/8vr7//4lOhgY4YBclMzMO4N6mUsDlDq8BDykDbLgr1sm
uQDbm17Ox1+HHy2ClX0b3tSJLLi7nFTZT2z5KK6ctnqZYFP6wIqxXnPutb0CP8kh0dmNMlqQ48CM
3xY96KMu4Dmz/AwNCFTn4Dk2LOkN70B7BGQw59W5aKUQgSBhdJJfAd8KU/RmX+r+RNA00p4+UpWQ
ORfw1QR2g3RojsgnBVSe//2SDubllbkqLqUP8c0cY32mBYqHgDVVqy9TqY7ibj4cj6tc5qPgva9M
quFKxhaCd5cPnK5ft/0xYdADogThAy8Kc/Q/0e4ETBRGbHT1gv2FeAy0bAAiY8dovu7kEWdD9AO7
WX4SPqnMykl87HbPofeWGTCP3GdgmDdDGrj9iGENxLVgr77UoZCZ/Zf9eH411TaJ1NiQwiBZHMu8
5tR2+ZWoBHXIRGdybFaKc30LXi6YrMrEiwonpUiqZKBQv6+8lYdPLcJgDJJyVWONV8F6wO1vrEdn
8LVEbvhLSWIGO8BUbsDtg/r0/LBvTuyMFOdepNjZWr5d191nNHagTXqmQ36vNKrYy3c3NQaRdOw6
HQx7wf4njIoE7rUPLhgfYeLCGwF2VhCf1QA5GjwfSrgsOm4t6C1wFhGbamv7XzXUsnF8AWGn96Zt
lPBXRdot0UqvR7CleRrVGLkRKlBM/OP8Epla0dmrBDTiuAZsg3nXaKo1KKhOwALx1Hu7JpkkwSEW
GdQHZlHlINUghqBab3ijRp2rUZjm5pKkovnSKFsk8SLd+QyaXUlrILxvYyOtJqlPEQMaw0pGccOx
s3qxkOEcmlZF+V2Oe4UlIXID4QZ5WgWbbdnKRweHUfJk27P6nDMECI5LWQ1hLoJ9ytWfDLcm4MMJ
vClfwM+kFPzkcpMQiF5DcQ/z+ZNXx239C3BMd+sB7Asxr3im7AQ77jbBVuqW/blkC9P5N1/aTvNS
T18gHnXNAk2N7B9J9qLTRAn3xPDcburaG79d9jTC32oDV0VxnhSn0yBLHwKWOW2DgcKOy6Ha4JbE
OuqlbaGGudZ8SXYPGUqYLfwm7EulM8HFFeat5sRlVVRQ3uwiFqij9Hf1HnSs5DQgHtBJuiAadNvl
89jd7ITFdXWX/HoZRe4jXVclmUtuwjMDzH8EoaHLzoYOD0G0Gd8eLNVwWlx7+FUlIfocNoPfZaUd
ZK50FXxxJozRtKdsVg/2xQ4+XUKYAeaqEdZilxLIHKZLCcsvoQVhXR7KNJhclRCBAUNTkaWSnhAd
HSpmB7k9WI0NNs9jiQreqtnKa1IU2OuXnabUIRZTWpRn2J558GVbNALoqHoEhgwAKdTa2JC0pBZm
FeVbK1FY6V0Ed6MkPZz1cdmqUvTLcZf/2i/+RuzS9zj0PavMtzF4M3PIODwp+1SFKDoA4sZG57+A
QIC2bja2/GvFenw3UFQ7j2PFFgPTCRW/z9Esc50DYFY3tAiDE5pegmBU6UJLyij5lxDao1OmBSbV
5PMN8bKYzzQG3D+o1alNi5oH4kki8rxuHwvq9zWL6JLQKx1fIxRngujn3WG4PCZXPaNIpLJySJsJ
GKCpUezlHHwE1G3pdV/niFZibe+1nk0ryISrr6OKbHPhr//szrbB19AfuS39jPHLlCbANGFJUByO
qQgVe+aYgtBGat6VmkBbcFmNtcM62L8OW1u2wXca3iQ+iPMdPYVBddh5Mc9haKnhIm+BVyazX7MP
93pKkA2gxB+WPd0yuA9BrwJOeFFiwA+sSr9fM7RtY0k3bONHezKCH+97zRF6pEj6wQBozpOC7ycL
prHwMOUARXxigUBuMYJwV7CRkRe1zka/h4xdwTeiXReP0y4LGyeOj/oDXatzkqBMVqk7qaQSqiiZ
Ye5y0QT3cxzRATNqmD4uWajWS3SXGW/ygL65/qwgVc66HBgIbU6qXwvGxp5BlSsuVRN4RQo6ogYL
Fj7u3P6fIc5cU8cB0Z47D62NQcXAv6YMpncoL5X1pCHF2Y/1XNdynip80o8bAQL9YTLdkZCAZq0C
nRMyYK4OahHR0NY7527zOgYS4p0me8K0pATdR98iWUXPqYFaKhqlsTfAxsnUnJzf0EtmvmI7HpDP
aP6p6J5F51Q3rmofcqqYN4Tn7gTWlKgKuRhamjVTKcipHgfaiDRs8UIvjvmSr9zlu8ExzAyPhm/1
gSBcHJ21ZebcdbYxCi8V5Qt1uGneEewEs24brtcD1xMbqnxTaJXJdS4/W5N3dcnBzIGL8efbO3Nv
8XXe0k6Lj5Zge32hQ7vI5JayaGFA0prEDLkMoKCItNnTutrlawXCXfuBKKSR+i6oMCOCR6+IAC1O
05W8HVy+hng5ELDBHWRS1mD3hobQXYe5sgGUk0ybvwAl59R+GfJ5rFw26aqsm7mMkCzycFpId8FP
oqGBIdPXB4mCSElIw/WC4yIN8HfpNxrdetPdf8/BRdJ675QwgoEg22xJVHaJsnxim9YHTplyBtDE
UHUpi2c7RLAKEQM7xMhy4evkii3vgOWDESUb2jqK+pLNx89iEaH/7LQRyn1Jv5bYTrMK43zHLf2C
Aw4z9mhGFjT48CnT7u7923Pqf5ku0dSzuYBB986edL3MW2HGDX7y5lX5Ni1WDziGvwRu/Jd1lEST
QTnBRSC9FXF0C8VeVKiJvu/jpizSef79alS9+3ufaNxAcy2gkcVLVHDUa+mK+m0u3mpogEvazfDH
HXsVfBFFzMgHoEGUoi2iZksNmkp2pwTpHyPtuIjJ7sLRVqtTCBpJdED5CGIkWDj/yaZq4q17SKqU
tSEbhT/RQ76lspnS7948db+6mcLtfsNyWlekSJbLprEUdMlV6QRhB7VQoLLOU5cXiavdDx8Le4vY
hAMZaHDHttWJZ+vwmE4qq9ZotWzDeRyO42EME9TFxVvLfq5QfS3FTI3CrkAxCIjbh+ucL5CuNiGx
w6w0eJFyfq4H3j1tM5XKTOGdBFt7XbvyenrtKBXSQUvOxWoCjrvlQw7VrfxTy3FC2IAIEqRq+y6f
h9K1ew/g9iyvIhXY+1cmZSZsoI8VCiffUr3IPLwbH2qN4E/D8QRwGau7wJbFJ+4SIOyJ/IReC8jB
2zTiSzMRka7dqqVapHNHzS0QtVE3jh/1Z2vVPgPYKQOhj8KHoYr4RkKMmQIBE2Cw2KW0AHr1VmlK
bhq4Y4bVD+itZqe3uXR5nc//b4EFmFceYPj5H0Q9Hh+1AjXxw35R0wHU0X++4lgdoz+vwrR8dyyC
pMLef1pZgPKHxPl03h9zHNFs9GIZJQlYjiyccWczOc0HvCZSAvpq1T1W9DIfyrd418NgugSXobmp
NMy3VB7DxGrOABotUKoOMTXnxLmi8gia9Wo0TApxcvQM344BPUtOhLPl9V5aYp4mwJIUIqghPNiT
YPXx5ifA69AI84GVEQ3YwR9WIyvu1LXU3k9AiZkSm38M5YlvfZLiaQ9PPdiWYcrA8tmj8ni6+1F7
iAHt9hF8yN82l+PbmbEIaFcavwGqWI3z1AVaQ8SEk42ETWborkzb4K/DIpGzoFwdEcZIIJRQ7FPt
yZFM9Hl/P1Wsb/xRpEyU7ygfFsrndqbEy6dvyEfVmWRfmPFoVuthApVrrx1Lejcc0A08HIJk/jMa
0dZ6NFJjAUTKM+8vhxXRfMZauZzPGq79qcmCHzo6tNfapCbjZoJUGSL7y9EIKA8DJyV6kQgip2vF
eEF28uA8ApN+uoEqNMb3AER6q2a1SiAKv0luUVA5Bukr1LxT40auPzcNPOXkDTVqyGr9k9C1rCsg
kVKhWhmjaJ76mr8R72IuOq5wr9rlYa0ZABt56W/CM1qWr/PvvYp84JJA+Rlk8re+AaBMqYuiA5da
RrOcomSPxwPTR/5lpoJTeBJRsmS8+x+Oiwy5K3Q/Ml5NjfmbgElOtKdGk44/AS++1X6Kn6pCukZ/
vcHWMhqsCQxm4esMEx10Efs5UOxNzQsSUyjfz5binWVCkI1Cm65TcDWi4etcPAQLYhPdKoAIzZPr
JRuZhMyMXOVM/7ytaNjfsZYqGGNvMZnLHYpPyfrAFSxMfriMpUiIvSBoOksuubUz3Df8boayUreH
Sb/hltEIW0d9V+WhfeRirgLDWBROw1ol9LoVIntocXafqGHwaoVdTtEEM6dXRSc5iCPaOEVHesgI
RPK3y2Zz4ZM26MRasncnOGiaCDMsDi++3jq/PIn8GfLYPd/Qf9eAIxjhWPY7ubXsX+ROJy3Tc+5Z
hEqG3gz1iWXpBjujyFHiJkHFBbmwLppASkPuC4zO+CfIMfuHoHgDOOjH1w7AXiBYVracXaRBAVKu
S2I5uN1Ombv/bN7tbw/RvnG/KjykGaun8ritD6oJTeiGmBqeQ9kMtWuAd1BnGpNGklOyGoZUorQs
rO9/qjiVJM2eDjzCOiiJw7zVi87QHtrOypXbGD+WlntIzLoMrSEi8nX907x0GrsozYIxSJSPlIvF
PeIsh73WU+kcarkL5uICG95/NJGjJLQaiHWK9YHpZ/Q0dlA+mzUCAXWXgJEdm4e/USibk1owc3zX
6G+7ftvbg7Fkz7XSjb3OuE9fOaGcrbHPQU956rkjv4bLieLmG4ygiQ4np7PEWDYhTbYxMIcCH7r8
M1YQ+yGutBOuv6YU0WN9i1kCpn5CdIX6KuRBZ6pY4aEsIlsgSbUC5PVmkMM4uTk6vVDpmMygAipB
Dhz3DHxx+VVGZRGmYN/fRGDwzxF/0lnyrq3E6TrfrEv/B1U1+jfnOkIkoZ5CMk00dzqBvIEK1zN+
pYvrnp2PjUQskNqeFWlyzJXrKC3Lv6iKoHTEd73MCZ0Vv2karKifQz0J+7FFrbvjltgCqL8ft3OT
cHLNxpWVTHIR2uQNTYW75Q+QbpaJ8Zy29/rp6/Mm4F9cB7fgyC3HCjsjmbMgryG+ct69hnZRKGN+
E//kSLO8/NDmdJxQTjLW936+w1Ad1sK+VMzqj72KlJ1kKT1s0LQPVXNJs0qEG2NFHO9K3Jh0IcAy
yzycaz8i/kRr4d8algsfjuAM8Nz8mdxfMbnIfJfRn+ReSs/a9YFJxKXYZ6csQQ6XRXoBYKVT0KhI
KXkn//00yLCk6aP9y2d5aktCQuImsgNultpAFcS32bbN8vCwyM4DDrunhuC3D+d2l1O6gqEm97Q6
t6fmJrI5T/YQEO2PlLPIQX7ZSiOedixOoROLxzVL6hOGxb88xepTo7MminSV48J3dQEW+sPs14Co
q/Hq4XbUR9esCsbWQ5XI4r2znmsssu9fO9zHe9ZahTJ/WphdzvGPn8FaCLIT2BjoQay/Rz9GSbzz
IXtCQh4BBVxxoZTMlwfBmSQ4UKgcLZ8uFAqpAvu4f7oLcMTvB3rpHObvUWblK2WjFa3xNpe+Pk5m
qLUqlcSdiYwXpkKEqFGWfcc1JspuRluY3cP5D61eivkWmP+4HGNfaosSiIxK/HyOzQv6EXaM51Ry
sH8L5wOBBdcHMQYmioejOt2cVOKZRf06GcPJUyGX7uJNfDLRLGUX64s97Az3+7c+B/0eKs8Y8Eit
0B8fiCzvRUGCYeJlIJnPKZA06gbHxvxUeD4gv7RcS2fS8Jd9EtLz7V3+UpGRJvVA6ctLnlqMnMri
2V0td4bO008s6IeDm5yN3oD2+wEMoXIh0tb6lsl5rnySNHLOYYClqTcJcca0pnL6/kHYiT/vEZR6
z0IKRILwTQPNQNU9jNHb18K/WG0Ua4JoQW2ceRYRocfd1vqHrmWL6Lhx88I/Nt0NNkSMexpuf5Ep
zWpO1aIdAVrLqFmcMWzX9wF+jsH2zhk6kvWqE0/ud/nt/5ICF6quKMQdzjRjx9uG10xXsYbbfB/5
TO6063s0Gwg/xQ67Ti55XVSPXM/igZdfOSl27Y7RPY7Bm2KhZudXE9z96mshNxZNeiTBnFnD+kN/
bTDO/wqSxi9Vyy5OnFGi/sZlPVTg/bN+q7+NHjfLUJjBYe2bkSw8JnSlQGEqUdUrPdmuBmvauEqm
ywKWrMzNJhjvuSlYOoWrSVl/4IAxTgVs1E64ld9v8TuIP3LmkKJknocubNbDv14MjfmNABsKlo/3
NEk6s+Hsq8HRaup8o2Et2kr26EdniocKD/jdoql0UiCuDQawNbkT+3Gjp8nZclvt0nF1+/vBj6Ct
cs8G0nlwjscFNkuxyT9ZFXmlorATR+JS8gy8arEA8ArKLIkx8p0oODUIPw1YEM7SxyfCYJ26fQ9B
cgnpSdlORKO4rY0GNKeyArEq7UPZIZ54bvnBtNXVs7kNwjU0ZPMvS1l8WlVEqwIt9F7Zv1LACm3B
aSCpeTAEk1n8VIu52/SpGS0aXGMWhkgZLTvFO4IPxntgpbFBpB6sMkC1wil9gZQe4EY14YWBNRX4
UYZDJDV63ZhDJ9uW9v/8aD5FYbpuoEaHsbCX46Km80VVXsbfmh6aZFtFrACivqLYszV4xurqtLOR
4WH+ZfBOIiZ9znb8Oux3Ft19vxnflQrQXti/oO9lEfXk0/Yd61hvcuQYICaXVjV9JKcbR25aoWee
K9vs9SIo2L87Sg+a0KitZdWPr7BudEQncYuHXONvfH19gI5uO3lltaTVBdLorwPC+XqXE6t1AYZ3
QznnBJC6pPsLw4z7zkW+rWssJCZvfC/EGPB6HeW3q6XX1+jH2Wi8083PhuvGEkgdb9eUyrwaWUAE
Ogj7muhoO2zco9n2N2gF8ZG3PdoUeKdOieQx4Y1+g6Fwu4LN6ulwpXs4tdXKBlXYh2S6M0F6vxOU
gOj9XyFSKpxS3Q8xY4kupc9iJ2fArW402ALhfp6+yMgmvbPgfaCuZKCnMpWSw8I4LSe0oOagfhgs
HRKTnHFVtjeG+cfeKRg5BepQMLSSB0kFJ+roZu8yXlFX12CdssUnPe7he59uNSJalpdLPP+fxGXH
UTm9QExKbXa/YReUXZptWkVR2hd2Rh+rcvPbB8qbGJqSaqc1rhEdodUN7yCcuPTUPC5cqc6xiCKO
dbhfLfS/M9ts41PbEYTYoki2eCvW+v45DN+v80YN5DgxWQuPOn/N7MuGRJ0E+yn/EyfpLZ4NVQdY
cUkgIvaDnyTFku0SaDqkktrigNilG5FJsBUzKvFK3f/aTKc8wqRCcluGpWRQsnFBNHQ+rYIhGv3L
8fODETzWcj4LRpg1xv8wF53RUDUoptLuqKMOpkUCBhV4Bh6mJn+0vMYgAxOk/k92sv+0U8CEjJY4
tQ+UtW0dc13EdQxqGHlrA6TBIh71GvZsolunjSu+RZ/RHoTjrsJwY8KEVUZHPzeElcyDdxh7KHb3
/w/gNwxD0/b5CnhuWGZz/JKC+yU1Elnj0nhfQVMBElwXuPPjn9ByexIHZzv7olbTdGOkMEEqZGfi
rJItcMDCEMw7hVpj5GmpMJBnm3FuPjGFffyycWOV+lP3Tc8qu3VgMOt846PzXwhE3X3qvWMpDIcI
jpsfa/fNXUk6w+BVsWOAKmp7J/W3KpZPc6oLvar9wqnQ/zHZ4oZzz/Q9PntrshYZrnr9P4QjRPIx
ECurI1O6TrIReJXhfK3yrXHt4GfMobZ+0jkPOa9ZyAip9/oXpiquAYrLdtkkBmepVGPrMPdjsOxK
C9CEVgVwuzRky391Vdxl1tUoWXydet+96YqOuDrZsd/SVnWPV/FHXEu+ivUm7XGNOint1GsXy0yV
0ifv/skTEF0u0Nqd9QHdARwyRxooB3+Um56hX+GHJEaDGUkiYDctAT55tPkbJ+ceng2f4dvjX0/s
Suqtpcj931ZXrKV7MFEa59p5UpOhlWFvAAjvmRBYCFIWNWiGwSrSgx3ZaIlN6yDrl+lqEjkj/WFF
NZ/tdeUNYtKNr/t6neHlCHQLF9tnvpcNFAGdP1suDvSrdWRv1c7q/AIOfBrCncvIYRTiSpJv3Y0A
C4863+qIEBEOrZ5qRUGj22WdVeJqETqOTmiyYcWlarPiBdhbMBPAUjgE4ty/GPIk7cV4eN/v3U05
TyB1gtu3NUd+L4WhepZlj9gqWARaR5MERZ4GHBCoCXuA0+o6iwYQbpT5RdXK8OVp2a44kGh/rSAu
bIy7Ei5FC75YIqGwz1gXi//N38Qmy3ve1r9xZMl+CGfLWzXCdaqXfLITK1nvMeNnJyYe4EEmvDeX
t2AWLP+s7K3BPr+3r0TJuYvtC5EQnX/Ntgg0viopL3nfWbfHd1/kCmTlh/FtkYnx7sRZ84Co+IGn
yKdx0CwoT3Ic1GnjC3uhxr1JZt0nNzRVtU376TLLT6zaAyOPN7XJ8GN7tww66SzbhhZc4V0bs6dI
K8dBHP3ljiDE4Kx7bJpcDgtdiftvB2+Zt0vWz7Bm8n/BE9HIKoiR88kEdP763uATEcqptVEAqLSq
GLzapYse0a4qFu6DAiGzSSz+tuhXlUrhiDCGBEf60M3RjW91b9O1QvWJ6wphtWw59oYLcOHaiVub
IJ1Ox0475onOzJPz2zWLVLESWHI/K+nzl/nxg+HIaXFOQWS7zfr0bnokYCBgZ9JRLeNeDaopHf90
WTZu4fBwlNc9tKWxksdzp5mNSaolQjBmvjPTwdtEiK/iR/ETV5sDqi9mERMgcGhhyUIgexkKBvaT
rtrEgAlsxwyda1ThLcF30O2ZpCTsTX2WOu8TyTveKpw659oTaSezVdRc1qYoTC+DIC5r4ImLNjjs
Taeqg45MecFhyz8d7msE2E4Gds6rHuVQDBmXq5Q3518573BHvYVGxATtaTLl353MCGyAfNRGVDa8
4P4xUVN0c95nni4QPwFk5NsCi490U6pJepurV/S4Z7pEMy6z7HGkGriwC9OZYFO4t19GWFTnLnO9
bkST94q0USdtF9FINc8STAb8RBYYdklWxZys2UT/0ykdrAYK0W3BijSBgp+wxKUdMD8SDukxxAPS
qIrLfSmz0ex8wjHIipbt9c5MjQ8UfSKXzAW1S5cxJrZ+/Fz8hw6sQS1lua8THW46CcHIg/AV7kAi
FQopnIpieca9spG6A4ia5GCJb81FrRKXvHu87tjOu89BISBXeojveniF6xr5HRLRNwys5b0MMlky
4sFWXvCAJ7/uUy6eZE/GgkDUUukXRyG72bOlNiWCrKVqR6GCmXn3junsJe7/Ga9+FzRlQHY9PgD8
TmoDHSZzVwLSw+SKdXLRHUZ45fUCOgDLRYt+0xFvehXzORmI68WH4NrkIzEp/bOQyuc9tW2P4akd
is35b0Nrm1DxqG6ZAya5qiVJ+66AlWomK6hRXDcTNkCqpJ7LwinYf959y8lGLJjw5rNTSSzCVvwp
rlVGuw1WGsUlKpO/iB+zw6CotiYDeBgLQc49Y9ly9DbBgS377w2dYVsVqAHKTQdB9G4Mybei5Elc
51WXoLnsnPd7ilUtJyO1smv+vBNczKRCqejUuluJs6ePDgxl7KTbIi9NexeqRcmeksOzQtO9G4AO
O9+aAvX5bxVsS2dnPpAyaCYbkw4XLttj5/Nts7JsraX5ocoYwVFMU1GP052obej0Poa0rg5+uw6G
RcF4VnZ/gqenMIU2eZwgciIkrCZDLCT5MH6kDqtNHqwk60JYE0dG81dLQFT/H4BcZStXfIkuJwel
y46fG2rcRC9n6CMxkKRTQsdohKAC+SMDUkP5V/olbIjVQEWibL/xvC69hzTr7eFyj1MBYhM9scGX
doPkSywn1vNLPehi7SrSWiJoQPbqGd93TvFDxlSONI9xCW3f+fT2FuuX9hiehmgWiyCFN2wzJfXC
F2WRtjOdcKjzDPSa0tA5EsfaOVaFxU8LaBJvxHV9bSqkMFMe4SltipBFUTISFkpaFPNZ9bZb1/Ni
MoQTUWifLKNvujV9OsRPa6ABr/7haQZvD3CHJWR6fSVkxK1c4Q+rRE/QwAP86ogVaWErN1bpiAMr
mMrrK6Fs7GBe8xIpHEQRU2OssXSLFm8jih8eZxkscdo6gdTiDhhcJRzlp6+NXFVloYFP1iCbo1Cd
T6KFQRNk1NPFmU0i1k+v13g3nfCVQfOEJCe6Z74tbsKPuXTU+yd+SXJcVqyW5fAOqjFU21c486V9
ANRcw7DfA2dilfXEaXN6Onpk8Hl3PW54tvRmulYKe7DZX4xcL7WkqsSTqp6DSTYfCNpKiuNI2eMb
GK3UlAs9n1R+LPGS5SF4WAn6O2Waw1bVffcro69NWPChTto4AAtI7QwWnIiySjyCI7IlkndV9tte
6bfSLd5G9oYoOI+KBuf0Il/2rZaTRz6brneCdCSBN8lYD05YM7146c/Gm7ZpQgd/k3Zt3/8sOIOe
YkHZxva7du5JR7pFQN8TlvWaoK5rfKafUyKXerK82Qkx8Yw+5SGC+X5VhRgCcloCuIQJU5zd5+yS
DoWcVS0I7d5UQGIHQsLYk9sBGrkINMxDCNbny0IBArdSItkTVmNG5PWBeze921ItmH/QbDdmtOIq
v5OX4VVEjBoqAfOVWQaMwg16qIb1HANnWGIjvLp4W1cVUBu0J3JgauiEKXPjsaaj89f/IvJwguOZ
Xpnu53dgoprAMVBUFOjnT1TvFAOedmYi/b/h3o/fSZtr8RdYeLXzm4YCImRt894XEpgSY44AVJTZ
x5gjpNRJ9ifqki8G7HyKKXk3KWsVCCmDw9TPvbnzvbMHJx4m1EqFCFWraTjDXoRsX6+6UAb5X3JX
sftKFfOJUkuuQ+iPNLur//smRDzm8ldMht4aSkWLX85NHbcoOWi8kilLFCdN4eC2fvKv4oFJsYoQ
3YPhTIaKnYfWFbVkPCCJtPnbl8gZwDZ5ORBSYnJy6US35vtg2b3duGRNC4t2BjJwNsbW7nrCyHa7
ERFMwxQJprahfTeSHDXosCVH7TmRqIz9YFURXAHDJHGYSHcv8tXn79icl2ABoyCxlOnSHaxTtA9W
YcvMh1yr+yDUzoZg3nU0S0oN/LwqrGnx2+WSXYOm1eUYgGkemPAyRD9FON+hJMaA8qlWbQhHnujP
nPIwviRl3qwHZxW//H9WS5xDsxKsu7eks8b5tC+MU9T5Cm5Y2mG10HtoZXYX7CQzwfc+HsmV12eO
j6PChBD6gZLr1Twe3KaOThCuJoURzcj4owxTLCkLoPIZFk4MojgbraB02ctvtCt5VN8RJ9J5CraU
0nTpJKcKBUqGYhBKsJmUaOcu3YXIrUdyrktpD8XvukbYU3A8T1jWGHzB8cuUBTbpcWyhHh/cWKjO
d8WfNBl2GICJf8yo+KeHXCn5IlDuKCjq4MB5wWSYPp6K1FObNu2MHCSN1uN2pssBnuwPWtbN1TKO
P3yOzw2/x9wQEybNpp9b6m5STheBjz/8jMKAIGh1S6hPf0MZ0cQ3eVttdJNa+agi1QYJ60D0roH1
fd0BhEEVXkAbEUK26jWEx+INE0U+29+YIt7qK5HaNd+0BcY5kPD+j/14PfuEW9kk3WIDEvbDPBNO
kf8Mbb1+TN/A+pDIEKIwLKjiGvuabtTdMo/p+Xod8RzrOd5lZ8GV44fGOet/nMOH7u3Oo57bi0q7
DHBrEAkE5nEJZmZnSyvqfHy/ojZCCGEHzDPieRj7lcp1QSri4lCsZ3MdAzlCuSdJEb9n7n1S4bPF
OXk79y+JHcGTfMhB20CnwmN0lpydRk6RsxtudO2o5riQ3whcyJqiSo2NIUiFMjikMbRC/X8QjI4h
a7nsrD5onLSOUGKke6vhAfbgtT0X6Nt20pYht9j9d2hguv3x0A12IKs7LsEyX86+y1jge6eC3+Av
NaxMSWp5bcKS6c2GqKEa+nebKUiJF6GeEzDNSJRqAk18IAKab01Cmtn6W/zlD2Nc5SRtoQRIK88E
clu/PuLAN2AN06XRUYgq19o7LdLQKkvAX5Y3Qtv9Q1Dn1fLNqac54oiUDwgO3bWHUcOJaTRrj+lx
PpAMppLZLKzj66MJmO3r2i06NwO71wyXF+5P/j2t76MwABtYVk2fX8BW+zSGBPL6x1jqvQP4AXWE
zeOvn2EinaRJM0GEIeGHclqRxGekBojpBx9boHnwBcVswQSOHUZdHytlzCMps+uCWqI9EOgku00P
YMGgY51FVz3t14AOCrhoeBIoyCX6JjpTS/UhPVmFAW1/tXo7NOMYb8hE07a+qkHJJ7SzkHPu9P0u
YqDVJby4i+v+C87vrSwne7nvzdYpA47yvRg02nuab2FisFj1EqbvapAF0tL/Id3yeTitrMzffrFQ
0ghTAvAdP7GiZI+IOwziVOfVxo5avBD5EUtqePIDJU00EuVKMf7svHaK69tHjKT2wL4pmWMPTPd8
z2A20kZF9zqDla9fom6nFbtjTDyXUy1VfsNe3MpIUZAlURS/lEm0Q/xDXBSnYrd+5gJ+h0GrnNkW
RfGmO6cdn5BV8QQFoHGbY7Tnhq8euFLR73jTYSRo4p2dychI+DUKGcAvMczYj0TDhVlkXEjXa6kG
cSNKxkArCRxOq7Y9g6DeIA12wjVz9SEAixIiulybz85sUjx7owm0l+KyxOlfQZ0O+Z++bR+5Iypc
DZ6izx0l3fCOJiDOXxA+HrVNzQ7zZOEUH17va2VsAPAJ5q5tRd/juOwpcWOCeZZF97YhnwNWIdLR
xkpJHf7L2fb7hBOgMqPDBfagLx33Gt1UpL9Pzp3Z9MT+rd97CwPMv2+eQBxuyVFTyf2kCn+WJj+3
o2U/kT6+JBnoQkRj3snDCD7xNHP6GqDP97eA47CfPtGyjTuv+b9PZvBODCHgZuD35g9iNahVQMf7
/y7G3YNS+ofyNmpciyJV/jI0F7wE48q7hyLsCbEbZKp8srCy8VhMNhyFvxwPrMs2REF2zqvL/XK/
wLSZAiNhTiGuu9evNq/sNN9/BRUFTZiS2WSxZwRBcWS3/OU0WRSqXNpwm5y/jzKejH6WZAiaWnE2
EVEZPoaVIRxpB5IPW4wopjHgt0Erhd/Og/QLWG1HdgsD/Jf3HmhumlkCexoe1rgYgkxrEk70afm6
GznkPLGg9fVeiP/rjzlZZVEscxi5M8D4Us51w9TvFte4ZsWr3kOsd1mp3o0PcTAFZI5iCRxCX2q2
Yp+ckF3DQs7EnKDY2FXI6yOCGMnng9vI+ks6Fk0iSw6908PBVwphLVl6pKt9FdzY5kDleGZni9mJ
uEN4hmMbHDXBqj3wnBXYSTYprZHmg0ecCg4pmHIuGJA16MaYQTJm9PXIlYG444ehLzRPXU/HXyRl
xp3HeVB3Xa3VTK614Ypt35O4Yqg7pKo+6ArMv9aeHZb3n2xdhEpCOXIozilEm9VRs5TLFX6T5sR5
ROOYjr2GArLtyRUVaqLuVzbs5l3S/6+/hcaTRvlOFQSTwekqSEn3tebHvwUva/ElTYIDLWhyUNbo
wNXW2wrIl6WWlpocb3jRt1j+TAmjkwWEUNcu21yaevgQKSXgdwpm1NZTMBdfCOHtwVOgdd3N0SAd
DwGtAMGMKOGk/+exuMUKoYrFEsoFu87e2tQFTrFfSrzJbrvndStld4tEpZ1LNM1h1XiaFLOjYQTU
MzTAuRSnEShxT+VVQ0st49pSri/WECH9zxj3u5lNW3ZQsZexb/5FSGHpwZWPd62Sr3vUjiOR9qC0
21XBcHzkBhLyUat5xAjAJy/4cfSo3Ks4FEcs5Q7s0YFSllIh6JkS+152I4/vMbRa24Lg7RjTCC5R
25PAv2V5+IGC+rsOo1DJBHUlPiPUXasqwiky6oZWkqNIhWjQNTxDKDNYnNcJokgjzUD3J/q91h1Z
e4hXq5OLjJRfa6LFhWztyRHWvdMQgj8sCGCmY9nDkbDkQEwgoExQf0MuyJa+iss50xn05P93Iejx
aLiVJlo6J200C7hRIPvvT2ZpPLuiYj4YdyKDt8okKFokVgyg7m/AXIcQ1pJqTaHTNYi9L+tzXi5H
rYuRyjRaM0Tr5+fDzIrOzJ6grZpQbJLZkOPRxn9dAKU9qSCjWsKYICqJuaZYsiiSmfOEGiA0YXYo
EYMOcqr9czVU9sR5yXCVNND6+UKEjFFVx0Gz8o3kT0O/QlP8wBY4c4KDjTKPnpcpNErGFr4WTyGs
hqBdpXmGcBRgWJmSDiPbJRp2hx7tVzwvBUOWoPDxdeIFal2XP82lU2YDg6ahBc91er6tWfZ3chV5
+goyURTdyI4qwS6EItV5WO95Zys6n475wlUUv5gv9R6ZAWJlTXw6jbSS8z8vvm6pYFWi7BDZ0BGh
eTRPfGiuJT1Bnt9yTomMYDNCcwtdrcesVWqKmoXiVymAMnTXUEkMvejdMZ/Oz4HujAO4URBG0hcq
1kBXmRezDCSuboVDaLKTg63eppLWeitEhhJluunL9Zw2AZaFXQuIyZZ9376yD+zfYp7U1eVDuprg
DhS357Mt3S3p7D/uCCxuheCzQH99qGFa0IWlYAqf5ZiiI6eMS6RkT6OxZMex9iDJTfoFKeVP+UeI
riOfbVhzbi5x8TpaTI7j6uvle6cJfjSlKSx0hBAMo7aOUbJaT9yb/7CdssSulBMzT3lbnl9RKavl
0F75l7ZM5NyEmlKCnHMjB6O7F1tPcYkjvm3oPm/Z4AhIOx1fVgEK9gzPdUHk2WhFnjQgAZ9/JQnn
twVoTcI9vqoJwHHfu2wIyQmduFxwgVla0UvoVMD3G3V8BuDeESKijwlzHRPJtCcMAeOZPPRG5ljG
8SuOfHjUuXKxFi/o2c0VJAJGSTrfGmHdqanzCGsEEvKDJxHvu4HETNQeP36yvK6uumawFV52VYft
H68jY3jFzHnsVSSbVjkiZ47IZsVmPz0+dhrKij2l8HveFev45iPoaoDzQGIaZr6qoXalcSMulYk+
aigIm7OatUBb96TdyWcCUe3jiuy9u4MaDYPiF4+S5nlB1DeOmcNJtzDgmb1DuEWH/i9ZSLPbhYm/
oqY/aM6vnHpQozbF5noMDYuZXfURkeZs9IKxmPSJ4oGAo0m06VFnC8r+JeO9xBgojalRBTupzEcV
PSm9oefxRNPxsd46D9QTPuNkxO8NE+6LaOkTGGClycY3fG3OIVCrCUSFY+lvi23IuOm0pfuaKxzB
Zu14h0YJLkQ2XPYHLGlfJ//OrHAB6NqLHP0SR8aOJyV66tv10iLvMjY7KDlovewwQqvb3yjABnMB
5itJBzJaZk1nE5fVo4CyEkra+wcarRNdww/buvafRYcRo9AKx+QrfjgV7HtmZQrJYa01evVmuy6a
DbNhuVJavhyAkT6l19hrYVQNXTQ7vhcK5WmTYctVFrDoHPiP1GEUP/3mp5uE8JacSDMYf6Gsvnnm
PNK1By2vXxiySD9Bt7bcb3nEQ5k9RRPi0j1LqAUrQEi8yQji0K5hL7EXDYCRjCVQIJaYPkUgH6wy
/QfEinYB8jMBBKpbs6rdJckkVYnru1yMA4jmhsB46NHHTEk5iieyqubPGv/RyspZI5SUQ/Zdjvgq
fmIyhcf3De9c1z8RUkyd+vt49MdHVOkk6X1b7jqJ2v+DGFSyrO6VtFZ97v4+QbXlMNVYO0P1Y3TI
5j1jTXL199+c9gnsYKmU9dsPAs/SYhKR017oh4LAfuyI7GbvKZ45QgnmPepp1dR/nd1tF7F5Aa0A
LUavLjXo8qP+0KZPuHMkYr6D3rkfbUDcisESqGkYbtWbVApRBahSyaAOQ3VcXChTthiHrBfnTv5j
dqn2h341eYykuDFUefO3BEMsKLgmoXrBGUadt2rb+RA/Z0cFe4tmduHGxbuMzuVAeYqBorVJgZx6
6pOTV7t/yD6WA3NZPi01I9JK3SShn9hxHBds/d47B8DEDXZC1GXAP/rd+RirVrRLrA67Bu/MlZg2
w7Faws6v3qXBcVkMeK5kLPp1rR81inzIZKD2Nw6vKwFlubGTa4svL5d93VcOyeJvOkqoxRKpFfip
V/vd2mzIqfWUoxbyh5wHxcidjdAOLuWbmN5dhcMKDKSJEbBYmzX4jw6umhvJRZVQFaGIGf4MigmR
U1NzWPyWmUso07L4vraf8I+gIClMcWhEFehoWgJVLd3IR7ayP5+giw+1DIUgBwlQMl6sHjoUvlFC
aS808bVwEl456vnrect2dFGXuwt4aWfaMyWfiAiJMnV9OeawtU2VY2zl9tDXee8Aluj2xBhA85g9
GWeKc5LXrw9Vjs9EayCE7cXcip1og5rEhII30VmoY+tJ0GbRGz9sI217ndEkc1DGoHG8E8CIgZMD
EOoHG9FvQWRb26I0p8Bo6QtvlbwtxplU3TpE7eUOJ5JEcn6pJFdnnwZQcGwF1mhRbZEpur5KsxBe
TaOEvCQlz8iZnxboeKQfdOEmFIrWY/HRCDq1ck9HcAoLnqktzyQ3vRMPfBY/Rj93DyI40CVjHVH+
uK72N0iM1yNhRjsMZjI3WFvuCLzRrAFIRbrIiT2Z50IMXPfgy0HXNLWrzxcUDKvoGh8gy7fOZ2CD
Jxoyt9fWWCMo4BLR/nNJVcS0JxuFulJZ7gmviANQoZcV3Ooe3PPsX3nip38NWmFW38MFQyDZ7pxh
1sApNLyLcaQTN5r2BXrBHC09jnZYA41HozRJZSkUnQmb1br79cpyvaoHOYwlu/htwHxCqAdUhu1o
n7W0r+d0wOge0E0qYXWP4JcgUE+M+s5W+MlDOpzWRmhkiRAr+ghWFEamf+7rqmODZ9MXnypcurz2
JIW0L2dKc8Bgs7hG5IfBCAiBVqQimLgmSVIF89TyfLxWRSVHbGrV8RevK3NCY+FEybN8ThB4/85E
K0pYkN9g9NLAtkhWhu+xI222pWsJukk6ZOtUjCMgj7iCAC6cP7F+mRF24Gl6FZnY9ZB1bOtksKzN
g58Pd4SRUz55ASp21LCtyUBBibjOB7ObjGf3wG3P4d1xWZyjoEFYV5WSrYnzxIurn9ykZl1GBxCN
TBvE1Zs9diiENosgF0XUVeZVC7u4lmn1ROY/HgUCNLE+HOvtok9gneZIS7cMWzsgmy1yotMuujgs
ppJjl9YSPMvlemOsMifKUFPIN1lOmsOFokZwmNB0D8eh0nagZGrYFoHhJvktSf/ftLd/NKIOr0DU
B3q8ggQL+ph7eS9nh/aY3o66XjT71OM9zt7iCXHh+YP8EfQ9eoJegL1Xs2hB0PTYqntRt7Ro/klm
N39vlJ9NjSqogJf6kPuBCUdopzkMDcXRsnHdAVUhqWVh8QddPbQDgd1B2BP6BOoO5/mSA+2Bj04j
WwE3FNyTkEaIfNRcPWTLm1KZeRVy240ixtlJ+CgJGGk7K1ViXiX3YqQ0PvQfWkH3nAIQTp60jUGZ
X/DJB3r1IE1fnC48TTTCorEvv2zJR8e8T3cYIWILpHtNIZdP2eYFYQTijVbLUuehq9sd534PsYfa
Y5ENDDfPrhbqAlDuTIL+yQhVW54ghRBbi2K6g3cVeQvhbGnSX/FgNV3Saxpx7cgoRc2iuVqicWTd
zWicrsXmY41KSCWRKu9TgQJebJ3xw3++hh8CIaqeyEdadvQBefuMJ69pc8PwnVUqaFK/jHZc2aNV
cUUsEKFSaLILoT0kb1XnYpcwOxZ05wJcj7Xw3UJNdeTl80CMIzzltIsQx+eOQgPSvF/Bn/lxob7Y
xLVN9EawtDv+a8O6MqhPtI9OxpHL7rEUXsiqOgBJPoaHsQd+yQ74bk6nXTrqCErLrYqVr2Nasxfq
wuITYm5lLCP93W8Qok9RdjByBbPlTijvcg9aORzkV6bDPFDKyyOoT5NLwHx6jCRvnzEEPU0KmnKr
3WtjlZU3LJpfecgCPjpjj4S0GBMKTvSEcbrO5XiZCP76IlukRb7LWo3qn4OWxQLa5vkFHdouiQB/
adbOLct1JMig5tc0Nj2QUyXKbEjkDKb6UMZnRILRO1/ZIhLFLQA64Yt1bk5wBc8GMdb7JbdGbcUn
jv0HPAmH1sLkah2e+zIfyZLBMadOjyqMY2mVnZ0X0XYXjz9i62mI1lbsSOJfjJDDoQcIR8WZJd99
AVTfHZCN2hYssyFKu3aNPYajD7WsR2+tNVlVtfmwf/wlJ34IaZb+uWiwop/lZgq+QMCzunbEwP7d
4/dkZEJG1iWXDPjt3bX90zw+3B2IKE5ecc+9xrAKDmI1248yZM3q+L7aPFyACTRy4F3F6T7t2nwo
HZ/LfKzuNP8gq+AaOnwJi+qyZ8oNNnOM+RTRWkEPjYcjdaf4B4yjsz5KSDBUFnRcjjsR8Lkf0i6K
SWOVMO4rTnt3kH/T69XlyvgEMOVgmBAxQSPbLF1lzx8nyDglDFLExanShxShtaTDK5dFfE+InmJh
XqPXogFe2Tcf1Se4v1dXvJIfVcXnXzyaYuhja1S32lj8g6i4C0FomiVuPcGdYlHuRCuCY1XVb5FB
EpcS6/z3peuMzf2ZipH1sUKvClrK9AfmEqKlchtXUyU9rVj/hcfET2vOXUYuQY0Gwqrl89n1H2Nu
fcDQwIGo9lh0zwlKZz7AIzZWHXTdshz2vw1wInCPsMtZ5+uMAB1mCAX2fkV8IN9AtrnKAtu12aZ7
9y9cRAN72qFhgAcTZMdCh0zd/AIso9a3VtzIvSZga1NNtPVuMA37CJ23ZC8sApSk3sUZRjPTJkZj
HU3YspQH/ZZK9eSTKiVu9OMjDcXYVEA9qNLv3c6afAe2NZOFWIKXSWE3gM/VrUvOq3cX+ofOJ/sm
yTaGDsyd0QDV6wBuU8Cn0y5kTNkvbLyCtUkCCPN13q4+j0+CQ3Hhh9F5TgZdNceAoShdhDtoFTWf
znuGf+Ei/XjJbv/UrbGao7M/Qpo3oe4MgXFSb7mlP7MG9UYOOhTV+SNcgrXOgltN/SkLIhtlAc+q
KfHDQJE5IKkv04Ok/pcOrLF0DcB0Wta+nT5J9qoRDLBbxZSM5uodePzRj5wNka0DGZ6nN1dGa523
NfNKKGko396YeeT0p0rzXeDjKvfv/N78WhrUZ1iePoTh5DPWpurdcduH2w9BuxVAmX96yWttQcJn
F1ew4Ltj0jmFeYvwrFV+8zmG+a8zHHW1vMkMMTuC9NUHgPOCKjcFKqB5MHNlAZuvMQjHOQoNH/v9
SxysSaaK2ZIKHnBayhsueA2N8pWYs0Lnxj2jDoBAJHAvxAzjjgJDrG22Wu2f1S6D1nrR8SAI+Yfk
XNMmugiGIt1Aih++E2kxRoJDKeSnXrLrsx8MXBcQoSIXi89rMRNgzbLUqMczmYGNwS+/fZa6O1kS
InHuTTqQfzfp8HpWT6DQutC1iM7p0PIlDycCY91fSlodCF7wW+2yr0Onw62+Y+n95VNTsD/2oIGB
U8fogUjQgY9BDPLMkSd05T3OOmaFIT3OBrk4sI4wZC71+8ZG3W2q+UvK110z6k+Y2Zq9phgflH36
pe3+VBG+1oq+hPC48N26mCIDaGnei/SpJD3wTtu66XvPpvYkUt/SBATUzgXEDCm97LnccVpeQnHk
eYdZdpyAkxyy2I7NjwdHIkCe6XD5zX7usi4JqMLM/U7lSdKn54nBAHf1i2Jia8VwRGf+4r/EnEHl
MPTa95yQpujoTCqgphLR3FosuPuZogKzKcJfTcGewEgIbf4nsV3oHwOY9HAdd4TPq1Si7AQ+dF68
FuMKQWcnziiVwzYf1aFgOVAZ+OnZXHe1qtOLbLEodvCv1zvGpFYRQGTug1VxwebRnnJil7vcbdbA
qSLbyw56DkOL3ux77YKeyQSrhe9WfCS4oR4HGS3vjA+OJj1OPpZWa+9OcI95kVKVqGIgV615X656
DCfAUn1+DHuohGWFdKYl7m+DHBsBvLIXoSC0C/9GS8XB1Q5SDQ8Lj4bZwX1JR3w5wDB+d0PAtuGz
AfpomnqDb4/VkWEUVDXHBxe6nn3gG6SoZHjHcz8qAWAl6D/yRCPD7+l57fYZQMLO2KsEm74iwPq4
9NGRkPFnfyOlO82IAytGtWZ09Puxt5gEjCQ6ywG8Q2qUZVb8eAVpPih0TyC1mXRw0b0vrDUwOwtD
BEeTZZhFEYVVwdBY4Lx1cg6Nv3V66BP6V1SZR3+a1diRC2aiosXRIiQlIHWMad4ZAhnSPwCNVFWZ
1mFovsHbYa+wcV4yZXm9KjASRHvfrKUZm63H8y+UsA63yC6eonpXzzkUR27/EKp253jCkfDOqLaI
heDziC5xJBH9t2Wjkkr1S3bTvoP720Gi2wsxK/TrNHqUCYkEZ0psXGDrym5L6Yj+H+7IKOMl4pYW
02V6UI4FpKu7BzwZLJFH+2QalFNgf3w44m/lGcIyf/KmgiOT9pQuPCRlHRKkab0bCAFkh0nfcgh9
qMoVpQNwllcCTL7uVRTMn2hPSFkEhuqH/9YX68/QAYoiD1j4j/jo2vJv0b45x6Bohck8vahnlGIC
OBD/WhSF/gJXd5e+xDne5B5pD9ESAdu8BCjdhQZTH+ILRw1EeBPYqvbWRdQ84L6PbmMy5W5QZiT0
9K0TMkT8pImNqQ3sapTnKOTbd6J9pgexBgSrKcDtDvw436McZs1sgIKBltOuwM7WkQhpmpcSff2E
L9IGsMzD6goZfeMpuPEQIW4HuutnWD7ERh8/Jvoxcwvgd4c5a3f3ejWjKNq3yylQZ047cKPYjyzu
/QZBtfGOnKaG5nJsGEHhJJM3hboOtrPsEXkwmJy+VxIFROnjqyiH6K+fUIM2u/lzC1i5Wd6k8wvW
tV55v7ZUCyr6um7nBqLTwCD11cFUZokfk63ve6nKTZkIRj0rBQYIJhmXPOlzx2Wvu5MdwVq4AJI4
zdLM+juKQqUrW1/XMzHbXoWyVIPytDPQroyzcAK+T26q8bjFkNsnDOP1vbWuVPW5xPtJKwdr1PNB
BrU5cpmDO9HcJfJ20UTHW4n+cr8AwXg4/q36Au0nTF+87w80D7vMks/pqvyeiCmTsAMjkTI9Kl6X
RoEhNTS8HtVVD3eSCT5aiTMgG6owKcPQ8fyvtSMU5UMN3bBXm2Bx9/9+N1EJJeVi2hrsAZ4thErn
6CBdYVZsliBwWw4H4/39plzA2M4zs9T2NTAWmmoyM6XsAOeqBzJ9VMJRp1RqGL24amlbQFjzovrT
jHjOXS49YK3Xe5tL42W/uOp34hp9PdQGZwFo+joRP2PpWdJh1qSbF8/gF6qZliBxC+zDvRw8ymYV
DWsEe3nzVQOXQ3gCxFoyn3F/v80EKONmlr1Tx5OYm1u0lQI623RaLVKuw87bFoTGl/ij9eRVkdhs
MePDUNXCobo8vAbYuMumzRn1J+2ek8PjkxMNglz4REA6ZQGRelEzAyG6iOqa7GEg197/G4W3IV5d
/EXjRXRusmAfCqI8ef8xgmBUI8vSUU6DWExKo1dqMR7juWJTQ0053hfZwwo9Q8QARwWhwL9A/7B+
n6JTTQC2qwmWbGRFmMYAFKtkd/czlgkoiGwJjMYPCVS4xjTFiSQWCWMxrQDfVISyOxreTupE4SK7
v9OdJuSekf9p3pQtbeNVIsrJVCbGyrkyGAYXpS7k/CGIy7dzgiNv7VusCi8vMOUCFd3lQcr1xITw
v4+4xFTVxudY0tlBMFXrZIl6veg53r/r9ZD9NyyZ5ymtp0xVx9gyMePKLPrwXh+zKBLfbvHZOS/+
nZmJcp/o7dOLCebyM9E0YAdsxOk9GRlohRq2tY3kVsSrboAVL28tEzfRicbgHWVZFYzin8iyEsSs
BsP6EcJXFrD0NF2MQ4uOAPfskTCyiFwlB9fT4Oc7jq2haMpRqG1atOcy5lpEdYP0rWflvzGCvMS3
qW5OR7cbwRzIzjDcdM6MwUUMENjZ5DuDPGPkpv0ZUji0+hoV67jqgXKbBR5pXbdyD29gL+ANimIk
jt+q57NBy4c2Bo3czTkXqP2Ua0Y0F++/Vaug3ygSz7tbD9nYI3pxLFPL62ulLUvs4UzWknCS5YeU
J2X4zZ5h6TG4F6qhlCI4iETHAJK8eoKcT6kw/LsVgEJutN1r4JCNSIhIEYgAGLlunF0DhMuPgmPt
zZ27Sl8t6lOVMdIWQe6NSu3JJYvbIjHfPImXV3FHd4jFY/S0NrxBobx/u2UhyJJy6lr76bX8kTNl
Bjrpyu+ge1wX093nLE2J3Wb+fL+0xIWXmHSDMGFwfnpT6jMq8rGyRKkA7Bgk8SJahozOh8bNTfBz
B8j2uVNyAf2dx3O+bUgzOap1ciLpIIsjYOfBBB+fgMT7sKr6ayQBn9xbt5HXcKXQMZG7Z5qAxZ27
lnJ4VMQ5BTEA1qA9+eEvjh5YEfU547ja30NOM8pNy/w7VVtWE5aJukPIYvP4UZIXWUlPdBojH+B4
+Ymp9UdeJySFT4hF/FUHt42CVmhONh7POe6J7MX0w8TxBjXNt2V7EPp9hRBPHLLZEqvuRADp5uSl
ewybsgxT5JBl617eOEOKa9dEThL50gR3zfcuiFyuab3NFQga58pJPSwwrqA2+Uu8yEhxIZ7y9W/n
fnNqdK9Bly6euhZxcWYZNPK3EafEwZwhG9okPTxGHA4DtNJTTf4JJ+VOvKQfWoCJCG2Qb0tP4scO
vdYyxLWxY6ktjt2oO+jOPcIDHrKnKGIltK5Le6LmtIhDyWoW6O0XhZmnQrJTdBcZEPW8A4isIRRA
2E0FI9s04FoZHI6q0BHQUSR2sAii9YOMuwxl2ojAAfWg/XIePPBVXiVmKPvlyEsWCrz7J8mrCNFy
akbf7BLT/pL1IE1UlQCU8/dxk6+ZUL8LmTQL09qFjXCIWnQyCO2e/E+cGlzJp5BYISI2ocFuiWa9
bKtbEd58bKD8THym74mhPS7/Eopg8niBVnbvFoz8hSztCQaqxXa2Z7NOB8d8pHMPuyC1J23KMJiK
7WmeGzUszbGBbfHZo33/fmNuswc298KEZmuo+U7lLpw7DoTbgUr0glgkTkEJYBZfOqV6MbUbWt8/
LwOJ3qwSjWy1G0pemplipYHNHh6mesR4GVANJZ37eaVrJXBd6b1EpvMR41WsB+8dnxDu8x8H4FPV
KwveSiyP2PR9zMuPp6o1TdDngIp0KyXYtoJmeuPVTdUDA4F7//t7NCuV9xzxg8dQqpn2AYMQjIMn
VexsjqS0e/dP9S0b+Choy8xJsWT4uR6AGiG/xaho7SLx9V+Sr/xpz9GdydLYoWEc9kSuqE2Rr0/L
IwEgXOJFg3zt3RroFkmVwxkZGlZh+47VShW7FtealgBOk9efEIq4V6vy9HKzabl9fRmWTKFziRBn
d3n0NxMQtYpi2PcglmthaJnG1KFxBlSlUEFQXj71Ihv1qXhh3A4hyaXNsIHbhTd0Jc8X+uc6o/AL
nlMuchaQTpxnxm4JVney0NBA5Pb95vtPI5FBOH9rsP4DGKQoQXfO4amuwy0aPrYoBTdD/4M8n1CT
xWb7wJh5MeLWzgLJJu3HgFpiruQLcVyHn0EchpBVeCqvUHV7k3j0ivnnm9uwy7gUK/7g8/nLDVBT
1wkpNZ98wPxb+rO48zN98/tHSsN6CFfgWrqnCpLhbZibhh5bC7MJKsnlBxIVLpkcCxiQgrlaQpcV
hoEWqzV45At0XJ1bZUp2q8286ZzNjwn5C/9jO4pWcs8V80zGXgEK3BCOFKJJVltK6z8Jiu8CYnQ9
Jta6v29LQBq77307oeukgtng+rdr7n3KDUD78wDksTBBqAjEtZeGwKiizGF6BUgWVB5BYDadTCU0
5S3NWbXuvOBeaLP5Huc/J40SrxLNt9BnFJdJI1P2HQMaND59afx+dc77QT1kUQhrV8mt8RLJJ4dI
Pxmkvb3CKoGtojAA4PvSlKXeJ8MqZEC1yQCgS/l8Cv/pnjRXlIexBMNWs1l3iNjjiKd4wOgd7/Gb
HF1A1fHNuGbQMdRU8wmwvDuHXio4Cr0UZSDqsVr8b8vn6vHIa/sEd5HHTfDkI5ITAs+ZoVV5yOtQ
kvF/NJKu7qDlhraQFl9YG31ZrxmhoGRHFNHGD4MhGiNEEbhzG6FuACmXmcLwvMd8krpVodgOBwhO
VITRRZ5CPQCI/vNqYaM0jFdgjShX9NAfSoyTH5i6Q8PAXqpvZrlZv2UL9ibYnKED5Qpo2jepIv9j
N63gWE4z7ZglkE2WR/PWBPAVQQKj89OSaD7IFtGGJk8fRoOvQ9C5rwzk5jc1KPNzvJYj7pHtUK2r
umz8eZGba1SsDLh+1UU+tgOpc8LXBLAr3RqDYvq3oK7ME8gWlOq3WpOZlTmihZEj6gTCuYSjLW8O
yil0ZiM/f8TDaDJTYpCGUa5xif3JI/wXGxGlTzgG4c/ZBzpeOQyl2GwQ4Lt5nqmJ3ycqtiaCJ1bj
lXfD10eXB6tIlfc2+yL90HAbQshWfTM6TT/F49nyrkzS/SUHQ00mIT7faMFJqTwmq+iZwI4un7K1
7x5a/w7yIiPwdN+cbOrCEaJC4UIolBe5GFUELkFvQJanl9NFFNmCHbOwl8zaGWvUuIIe9kx+QokL
6qVJfMHqt8NfoT+xrhgm8oWJoyy5QZFW5szX8EcMDOz7WLIOTpX3zH4bZDHrSCYaWCLMU+XgKWPD
bKET+zp5gWDydkS1AP3a+Ub8967/pmj8+TL+v0hn4uxGrKY7jDKcrbWtPf14D9aa5dAinBcb0mxP
H92cVDLoSqCYTt2NNDD6Ib3ppH+IVvFCk1N6FO6nfGxiaJTjYj+dq0+KAEAPC70bz4wSZXrMCsYo
lR6wX2bvjN/f2jjYxZZjBQQWbtbXl4QuDpBZjbYHJm3C9A5y30iWkh6g6KNgatUvdjjtK3BXHV0N
tTRmSZ9/A0Ud6r/UumMancXBquUMw6Z9LfniWJ9k1X8KTk8HS3sWKBPjnaGO30VSg5MQQN9ko/+1
Ssnp4h2WYvUzar/QuwgSZ5tBQx1oNhyOs7LLaC1kjGZLDrMbFUj1mfjqIJuUf2r5GweFaZAdzD1O
uNJ4YG5Yab+7pJJmRnp+/JTQuf8CXxYJTT/8ztUJIaSMIhjkNuQx+fO7qPuZWgM4cUI7NxyrGUow
LlnE7J1KJ0ULcobtIZemoI2EICxkg1ZnBJZaFhUQ8UccGZUT2mY6UrKtry+kEDlXzIjhgyYbll5j
QymkVhWlKVZQdxw+bEI99+0p1utC8WhkpzhIf+MkSteg+xCnDbZVS+3GNJo6JbaqM5ZPIAY9ucds
d/Xk8Dmwibao4PiidoCmxGE234OI5xGERE2yKyc9P8AmCo8F4uAQa108cgP2hicPH3dFJSGMgJEv
5/ega5QTZF84SxYGaSJnEQuN7gCdP2kYXnN9iqt4j+OS83CrfcdhCOrDCDBYtvJIiyoh9+eOKFEw
2DBBHtz+gKQpt5w8v0KnSYql1bjqnL0J+xbOrWIAh1mNj7RdKRCk+QMcuPehR8SHGL0btm/Ttymy
DYPBlrA3cTzsY0K1Mf6tKLP6MJfoqgibpUpiEuNNe/DEgMHZ57/nFu23to4LJnoO2DOGZ+GqHbve
Viwx9FC/cGFTMnYeLj8gEbHn7lCyxUXeAjrCgfoBkGvpe9oS5FK2uuNJ0ZhtM40R3z3/PupGvHqD
To6j2vlNC6XUvfkiQOEhX0iUfBSOgqu5FDDdbCuXkyChE0a0UOuzh2LR7zzp7S40CXiikylI0P/V
g3VuV29Fpyt/o4hb7093w4SEMkoJX/UsoI3rkqeaKLdpEtkvhXRVgQiYyysQWH1HqXovxexrRAwR
ZIjml+A76uCUY1fspgT951WC8TrHK/dVCqgSeRaKtvezfFfE1b+daUdcIff9PMiPueYIwbqsKD6Y
+NC+v2rsOG8WUH0l9avkWOUrlANT6/4LdTRrtgYZey7O9vUthw28lrJZDzzbStPROTU103hbD9Bz
IIdVwJY3g1zTTmzrMHfwMJIiqdom8nDRh063A1tI/dhvK+iGPW+YKD/1iyasj3EGeA982fib4eAe
OFK899vPkh1EPUjs4NA6rXdPvHz0Rrtb+HeF0hxfc37dIYEM4nJ+WuSveS9Czz9BjpFeabg6I1of
P5XDA/QTMh1PFG3AkAKNWb0yk3E85VYFUAC4zo3bCkV2okBH7kXlu6ZoJcI/1KqOdYHuSSYCehS+
nBgX0I5rTcKoPrfxe0pyl9Hz5lCPkn7ZolmIIkMg1KDlAMmreTQc59POxlqmanGFZTKy0e5vWspO
+225S0zUPp5pIOQ288oSXhT8ttwIssc8Am8aMFg6Kn7A01szr/690dymdClLWSYHQSo9TLgayPmz
Zk6Yz8oB5G3Kf/c5uRAhV1mJGtj9zIMwgSS2EGdW7AwMz7QtzAIkasM5CMBjAPMYaxpkz/Ne41YB
pzn397ISA8Snz7lUncpmv7x6cj4s0qP6t0pFuN0zX36LvNzUeuz3JniPNWFZHxUV5uxsy53WICaY
b7KQ44e8O82SrrWMrbVWmg7tWUPi5HFuHwau6s14FgPHY7w2RTMKSrz+7TF3qS7eRe2/SVQFW4cB
4ELwhWKd/4gczyHSvDPJeqG34+BEOIBkHyuzwd3iN+VzcI9jAt6cSQImvuziV/eS+wSXWAglO2hg
rrWNzxQzMzCO9fvl2ZTwzyawVR0/lQqcxBp12N3GCojnGP8kMpaiSdp6OKNOGFu8K03kgQ40RtcG
7wkMW1cLCKNjuA94VjMWnVgXDszs6+hmpoxPK1Q09yOxpMO16gvVrz/jD53yZsm9mf9RyKyI9s00
Cp360j25XoCFBkvRzuxAg17szvpCe2rWI0H4VXu0cgFsI3cQUgoTfXuoh3c4X5KOKgs6050lav31
I8e6sqS4cPUvKuK/7rbEm8KPrNliuwTCLr2VeZM54JeH0kdKNZ9lpWLSJOtXvN/0He26CgeUGXnO
7Zq9IvSfTjdfGH5CCAGXFjEHAlhRKk1rql2M7pnL2OhOy/8ibR/AA2uXuejgeF3lPO6yFwAdHl1n
0b2RjN+JnA4kZ2rgth+ECgAwnI/EKwkYxRJmniJe14YVZZ99X5BShietZTaTxvz/7Tue6IZKXmf8
3tZ6zF7r8pSe7lLVtyr13NXGbz0UMia4G/DCMPJ5F8lUrUMPYZZI+s+je2gvmbb6plfY5+UbZark
FiqYBYKNpYG6Sqe7x+e1kYGWsxZK+EDojC71IutXco5R0zGtZD7p7swcHlpXoQl595ykacqPbVDe
CTKDbHkUwvVAAyaFrbdw/HrRHgiUGcwnNYSUB9qX8Td+QU1eHKx50j0ua/ENTaOsGOKOsbN0rDpA
2d9AEAUCofP2InL7wsPXuAFGf8G9YjipsEJnQ+6mnfFyL5hckFHbU53Ugu+6irmDNH9ofh7fUsb/
iBQ/6jzlZWsJtZREUM3YZWN9tEJY94ALzZed5WkqCPMpjAnWwDW4QmJyvi0WtLBia5sMHc3IDicj
ij7tU+XBj9A48q4oHSwdy7S2QWTkUUgiyl5xCfT88XvyqKM/3NgSYNlo+YI0m9SlDPXlZGI0heg2
x3fXXjcwI5dXZehiHbE/LHXlXcQisJDMsQ+J6SznLtm79InaAHaSrXZYUOwbv36t5dVGGWT1PW/r
cJIu+adNUkOmPgFQdHnbGA8lFYHJ0u2+oU0tM8bJxL8l8rJCGVoOEpkpg9wy2F92tGdcmCfgBeA6
yExbFYX3XT1FKScO/Rggo80ZAL2t3KNMKuI/JeovrzqVkP/5zncnDDufqzHFapYXcO90yvLz2Lqb
rETNPBU13hKjAwe1hjHIgJLedCrPJ2ig22AVqXnNJE5dPqWKX5gwCvzv+SrCnQI1gEOIeuy3cuEP
/lvNUWTLsqlzKf6R0CQhpMvBXsz8Mx1rKAyCdfUv9blj+L++bg7Noh10XrXX5I/Cpu9djL7FJqxB
znJRd5pzkLd7cqii48SVnX2GBPcYsUAEGAiULe0tEuI4T54dJOB7lxDKLKUvNWsA8R+OirOOu1NU
ZT0GlqsDzxCMJXvgeC++MKlVXvDhtZh+OFYMeFxiXKhMwollS1Es0/TfGQgunYths/+g3twOpJV5
y3xaJ5TQRiga/+ZeqwvbBLL1yCCIJDMbl8HOL1hll4APhxjs9r9X8j6oI2Kx0evuAuMILX5wz5bK
aPVIBtZhJT6iEHnFOwgwJoDXnyVtNLYpX7TnYTNO80nfRk9KC5/3rnCXB8Rm1jAoxmIYo9yrhZp8
4cjESHQYkjf6faQBuiKBpqQym935k8vUlr94wFPxLSiJbL8399APem9yauaoFZLKoqXnRoyuTxWc
WIfm99sbXwaXQLjBxDpIrs4en1T8BGiWtzgh/8dBc6yXpKuu9YMzO8iyIUknxajmOk6AZnh4tj7d
/jjnSnMgpQYI+zGfu44T3OeYq2rsEyW0+JWOp25y6JLTscaiP+LzCHOem8jbzFndSWXUMvNq+dFX
IvtNIuYykiBU+Dt5W5IEiT+RlSdOXpFi1TjgAhDzNz3C08EgXoUL2SzsNqXnY7aklNkMN+Qo+6Li
+xEaodJDhnczuKBxgOocEb8Zfy8mXAk6JSUkU4TAhGl80WUYUjzhXxlLIOmSSG2mNtWCva7GN7+v
YVYxvdTcXzLDlIbU7krT65aSGGJ4r0VboOmTE3srqmaeVOoaAURv/mZojdQds8PnhGOlahrAgz25
wqt48a8154dgtvpg1XxlbxPHtgljmmIYysnT8SvfQ7PNuAIY5nqFTTS6MASyVfilVf8fXTMef2jf
g4yeP4UiGFsJNBaMbVjmAoSxmJHGXaZh3NzwmTDBaccroq3/Zxj6/HbHfPq71267DgdBzb65j6Ob
SvutYnyh60SfhP3Bbw6ul5xrV7NBoERCVgbxrMx4ou+oE6sByb0cOFTbJcKCjdYr2MG3QSnXJQGt
D07l2AVmE8h0xiVw+GJGgE949dTrgRR0gnFlGr7wfZt+UGPUFYXJFkkxgX9BI+FPYVFyhuGGG1Er
XkU8t80feVD9IXUOEKMw9zx2lHxsorEEJO4F6l44khSM8jBqlwORXO9KVm/GQrXjoSO+MPCL8zC9
gmWDk3uZLHxYE/rY1Yv/VsjBspqIEmHl/o3I3vWwxiTezRrUQFjKE90J/b4c2QzvNz+3cnFMvTnD
6jngmRz6kiea44NrcQrxgjZZ2+pbZgZONku3HPpj82b9LsX+6IsP3eG2fov+kNNb9tnYMnn1I+Oj
7P3xkmShXl/seSU0F5/5odAq1F86PMY1nKasJ4svgqueR7WXw1xN1w3ngoO6PK+XaoRTm042whsq
Lo2SzvojHhlMo1nMgOqI1EudJEPINsAxCUweCfHURg5l91aT6LGmb5xyB8yoYqbwC1t0X05S8+q6
fKpwhGfr8ap/lPafZYwNm6ASo8N7VEmPt+b5WLig8Se+PpDF+KpRbASWURHZvVSbfCo1LAJtCMAb
DMRtjVBVgY1fUF8UA6ytzBKfeKGbnywJrCCVuYOl8bNANU0Iu5Ho2LXjRDW0ojJBiBJEkBveUes7
Zw6nK7FshLa63xBj/xqcF+J23YaeUSQy+NQ4j46mOmsmC84aFJt83rIko4+TdStUrlxn9UjIKKoX
6Fsd8ZsNrDj7XybFoQOH7Cc6eomYuX7tbj1kpNWbADjzfHA+ps2U97wNzwyt/MYfDf6pa87CYiB/
KFQgfbpkjEHPsqyRDqsD1mtTM09SLBwAfCDwGFuO0iKr+OdaJcucT073QnWOAy90reI2KEj75lOf
ZiBUN5tfOAtdIRGBK8YHgIn1fd6iqns+68E83vQv0vYO6ui9Fj49pWNsPNW4ugRK6elJkODOALGG
d/dT09eDx8EcL7LVic7+d5NMaSIYla3ia8vYTwun27lGjqZIb4uau0Zv1z4jK9j2aBcDZ949gPot
iVg59VK8wcY8KgH+If9KOnCA6UnOIkA0S7pSQmwxdq0dlgg+ddgGgdhJGGilbD7rC9oByycu+KTh
+kW/Wd41spL2l0PdTUQzqAjKFJIHOR1ho7x+VRmzzIi+Ubea5l46RL3GQrMONlQuD92LBIvNEb9C
/egIthsjtdpnxvhhXcnL5B24vmZNG9ML/LoePmy/jTKIt691dYnp1HEhKwMqTbVSSrKPx/l2tQoE
wE0/gIRss6qx0V7BytSJvuTMi6HY3A5wFtsx6NlZNNynqbuaSDB1tSNE0i5+BlIV+PTqrlLg/2P2
itPZA28eGt6YWhZtM8HJdz3Ide83+1QAu3rinOrvBte9jafe08bwkU96DYRpKYsS4JgR6EVVOAkF
r3oiSJWnFbxgNygqxldoZaP6orKu+7sesqIi2VOnRpWLBSLPjP5XfeuAgeiWHzqhq5h4AMGntgbc
gtHCE1U56kz8dWcpWNXcGW/NogPc2NjdRKzbrFooiVi4mtbQeLlIP7cjNHrtA6IQjae+TgzkbrJy
JdepRdczp0ybYwQVGw503Hn+rtRrJxli1uXpu0pGpFR+n54GJcZ0v7rFGlFzXv+/7jeHMULXJn1d
/9FCMuJyEm+yaM+bRHl2TP7QDKW96RVaARux5yPqH5o6K2FzJT4E1n0F99+aHb3u53Xhax7ydf+K
Fn/v/Y2hUlZcVhU6ALdM+b98r+mXt/MOUVhs3dQwltSzYUIkPyUNDcaVjI4EjYqOSvTrFI86mv/J
tbvNyAiXyVBZMseN5qgZxn2WV1fzqVydxq3rU4HocrARuhx7PcaFAPTnMwclxgFGBmVKwQO6Tcvw
Z9ugmK4NtKF0clipa9FBpMtqyxtqB+p5e/dgRhHGOpqNZLwtLjvg4MY6SHvvEjUer798DWoJ2ZLo
TRWRvB0lpESGoMDFeNbOHFpxjnmSAh0RY6R4l3YrmtJRKlcNp5RlPF6hQ4O+Mcsl5l7duEobPr3V
UfRLXMkziQ6BP0xGfq+dD3jRPHhwMFtk8BGDy2vZ6LzU1roWXnuI/WD3sTl5EUksh1Ioz2aQofe3
xZNPHmGtRT+bT05do9sz1bFvbI5ZDLsrqwOuoGEd9DpxxDG09VzAOHu7+b1Yl3oKu7jAOK8uoE75
KyAuWACJEhLV3PXKlyFRSv9CG2whmNqmhhV89C5zDntvXnovnNiJQZf6DQ9J7YMfW5urinV5rj/u
Bnd5Fnc4wzFNUI6Ab74CRSYWunbDCMImSsJ+v66KrF4Xz+KOyl78s7ltqfptyrE3ZAA5IOBxwsnQ
DsXnKiEWFw6TSdSGTNp47UlC1s/XWAxPat2BVoaokoaPsQJiBtKoFa8zllBgsNk9n21890RtR273
HpIArcR2mL1F0tfj+Wh0aRiDvR7E0zd+EQDNIKhM+ka8kj7J3iI+h7WRvgKpblKADvgfkqF2+jVI
wH6ZQZ8Vs9O2WxwxFLhPWI3en3WzmuE53f9ET4ErIJX/sOikwQP9bXRYX+E1NLbI+Hwnd78LGLcJ
tAZsiC273pqDvPD+rkBtB77GmU8vyyp2I5d8NoONFPJoPu+Mekcd5yzplt1nT/v7aLGoRV3tUAfN
y+y0+Mjuse1oZZZOR6VB+gXW46JekNNo9C26dy/HyO7urdK0Tyzpdc9wWqxvCIkuZ7MVyfH5OdSC
1/ikeDf90eJrbzcGitL4KoXeIuRjnmrmdeR+7COX0PG4nz49PdoQYJ9vbd2zKEN4sGplj8B+6Dan
+GwO0Klic7FCIkc/Da9sNyTEuKxU5d+Zt7ro8y4ZTBgdhGDfqhco6FCrVJcOJhIlglE7LnrehD/b
61DeNz4R+3Q+Q3Neb5AFr/UGFjxZ1pT3B56bvXU6/glq/vA4XxGLnnYCLrQpVPwhYgwc9B3wVxgK
4cdilcj//Ap66Fv7o4f1fm4Iii9LafjO7JQ0FSomnm2vMxqTBYsm3pIBHpgG1lFLyxnTVNAEYy8p
y0BtgBpx0UpbBwxvqGFGVq4Ms7PbrS0JhG1S1FgiPHoLULwvdr9M8224SgwREBoU8M/fVTy30yGp
LOY4P1kT3cJSqWCr1Kl7vaVJTeGCku+eJGFQhWAUPkOmB4woEojWUsgNW5WQA7Iu/hLVOcuC0pBc
b7BFYf9BNZTajaY5fTUEzoMPn9XZOPzJ2tXpulKypzUr8ncg4GiCQfTDdlr1srsufDRGn61+tO5b
M/ICUSrmUj0lRt0q8mUKT3LOG7dmoO8SC15A+Qlbz5IZdTiPe9UnvPU9ZXYfm+BgpPIksvaKKjoC
kuOx7vJJQIqMEPV3j3dxkcXW3xBBfqDiLE+65IWZfhVCK2dfoe5CNEMjx96t96FEWaThxwMNBsWG
0kzosMkbalNmpABTqMex2PBpcC//V6H0ci7dpyWNjz+PyVUrVMkbDrthx5346JUIKleYBwf8RmWX
dfaT2i9LfiJ3x1aiNxL5vq3y1qMNQPMeG8ueu8Bk1FRDjifre5qN9PZwFW7TCwT4kJPKliQgYpoC
9CR5gd98vZk3mQ2qZdAmLM1mPa0NX8xKIK5spWjYiQ5CiRU1FwR2AKGZsPLaragngcYf64DiSlrO
VAFsRcVkI87mgkVNUMpvYcySXjNI2cAovMSRmF60aySauofc53lz0O8S5GuoN93Q1fG8+5EsUncV
aomvW3fkjfhf/pxW0uq5wa5WRXychy7n+4QrnkTOwHLNy+2WmIAI7f5ruZUAcRD2NwMbb2AC+iXM
f/1XBgFeU/YYh6Ya1kvI7v2nJroLXxOAtDnGKIJEahn+cz3bZxsxZIYajGhLpo1sOJayjV3RWqHP
dddGQuvHGgErXXwQMczl1I6zvnUwRwgVykydTLHz7weAKpNVL9Tv5pOXPMf7aO/NOo9BPjPT4ILn
AK+LYhuQ88O+eRem0L4HofpOyL0dkFxVoybi+cc6Kccx9K6QQEgFwBWhR1tO7uDH0UnqEVUI8lKF
zdXHdIwliOMKsOM5FphFqkOpLsye6PztWyU9ik7fPPv5nzSPtUxwA4wfBkDk0ofQl0KK82piQL/u
VGRUaVWroebOsjQooowsFj39V8Bnf6L1x2t4wh6nXpPWqQtFXT8aO9hfnkKUsT3vn9oP9h3mjZY/
iJCirRV24wLWcrXf5AMAHxOvAuDJ2j6Ji+k70t3jkEqwIM/rvOZrsEDlMW7IB+I2KrfbaUleqQ1p
GQZ8TcbtEz60kwF9MZtdovDtW9s81+AwpfWaqhD9VnLxPmPeiie39to1Bb4/goiRAQLnPAT11l5L
fAuwZUB8bzPt69zP/dJNTnwbjlw22kLjMiGGngoJ1DDwG6AZ42YzCdJFO74Gi1i+tyjHBwvx9rcG
QF8N7xD8X1fnEbiFh7GWDpIoy5uaIdWkJoFQplZlUyq7u1LW3P+KsAYcMZfBnGtZpeGMzgone370
Xva3RuJdJ+/wFD4I5OnSsnAeiro9DKfNaQsjfoHklK+oI1znli8N0wMtxH+euAZoC0dra2eWa612
b4MFp3RTTDjfKWGk6l//kAhjiHiBcZqtVoC7cuYQaG8SUkFgigzgT0dhhj2Ruz/9pQccI+InbRyT
A+fvMtzcAPubnQhhHQ8J180qK1rJ3tidUXU87a2LVTgQKUG+9JDmxX/qFxrblNGW4eW94AxYGfyL
hXBiAnOGgzinI3Kym1ltETkJMjlUoRQ+/0Tv/kfWOoUX0/rHUnLvdx9cDyk+eblkgLZZ7tRgQs4h
q0Y4DOY86wuxeQkwuMuY77EKe0aU4K/Xd9tcRvJSSAnVuM81GhmWlopFUAf08hmUfNnkLfINMsgR
DqkzGxBDhWgNbpLcIDtOzJ3VIQfN7JWnGptSixUWbpWc5jeobTYVaUokGlXzWWQLHq99zgE5OO6+
fXmGoyG12FoZlYOoeFuaKZ63P0WCsypw67eyWIDV5uhOgmhdhzWoiUEv14b/UJPrxfPhnUo466cx
uR7wyR3jzcUcqaMqxfGlx7uCkqs6RT5+h1y/w6eynqWf3+Kf+tLNyaOAU7irwrjf9diPxtWOsYPX
kIh8IqVxTTWBO98t2suoIx91J9XD1kkgoqbtCHaMn3K1T6WOCQdouwXOWXYIXd0T4a5OEBA9E7DH
OIDslIj7NMYx8qeF3n3hln8iUMf77xgcO2eItWFbVzR8dHFkqIi/hsSqWs8lK/7+gFc3g9dX4CKt
SnZnXRnnuRgRHDjFrFRgQmmfkV4HfY3aXCZXC+uVRYZKEWL0nlyiedmgXV8KiMtk+gpbCKNB5h/S
eA/v2RT0suz2P7fMUMU5dFMtqffvnXg2Y8nVKgCfz0MSdBHslx3cKzpLXkrOO4GDflkQvg6ps6Nf
gNSAhwIg/HturPSQ3rMKprdglkjhUOy0rjEGVTBBhT+Xmrcf0BscOf8QhSKokAGzUS8GfTpbuH2O
xhNHnWsBZQThLkG+Ugh2h0KRqEZ/TrrqV+PN4AiyHWRZJBAKB58mdn9XX4K5+zHzl4qBNAS7jfq7
swTJ13GqkJ8MP9UqQQhN6K/F+FJsQrmbtOG60wAbEUq6BW5wUcc+NwGHUzCcUAHBM6AqNqp0t8+g
ESBFT2Sxd3WvbIJFv3NbTdg5AzReVl7j8zc1lGqWREDJZgh79grlmhoswThWmvSTvtuDaypRx5OZ
3QRxA4ZdCvrdSL2T2i+HfTanNDslFUoWAhxm2hvjJFb03ZRQDBjdTZsz3TCZVGoIwqw9rRmYzbtD
DWom5Ug9Zei1A4o1OQ37SY7ful1RAG9TbjC09+sKh91neQk0VkbdA7kEx2pjsIe8Q7hC6lpy2Okf
xuAZskagP1E9c4xFU0E/A9p4DI7EjeE9K0tFTImKJWX5s5P3dAuPyRrdMMEyLeDhDUpNjHoIAi2M
JH7LkQB+CURIe+a/5gnH10YWd1K4BCNcWaL+A/CBcZYBl0qGrSTw3C9pc1JyhlaGgQODSDaSqEcO
uecr+sZeyOb/x6yc6//819/cMjQ/vta2lIAP1PHRydULbHx+St+hhGTwk2OL2r8JmwLkP1l+T4bO
73e/ZbxGwo7KnjXZH2PfhMHgk7Efe+HSoMSyYfClhGbyjaov3je6mXA5X8ucP9a2z6X5CWC/XqXr
Iqeb1AMCbvXy1K1/LRKBjxhyil0idRcTKOULrRQkBegJyauydIaZS06bymxFgnVFp2gEBE47m5bx
DSNpNoW+g5DwIMVGrcv8mILS9PC9FMgd0lVfp6b3KiNr41/BsUwsou1jNg0xxHY/2L1PTuck+GPm
ifuZUVUyFKcTKDg8rTz7AbZYF68P7ZXPFX2pY1pfinGzhUs2qadireUol/ZQKVzQmzSAcwzkTH1X
GXzFPolbvF93B4R3tgCIsPYxAl818A6N3RB/6XiBHt+VEVL9m3Xzof4BrXpzcL/xg9Ay0Qhev7dG
AnYNeHfBpCq/Ul3XSmyF0siQU0i2TaLN+ASfBWyG3R04uoaESTV3/QX4PDaXAtBVUWr+TMY/HOWx
yAE3GvSUB8sAjeENltPmjKGnaRymz9OFir86ow/GKTMIG2akfWkCt/ikkKYxCLQxlG7SSSeTdTwp
DC27IwrhoGwFYpFIWY19j9n2GxeYqGjFrSfwLEw9z/3vo4m10mpSkL4i0s4k9wF+3GraXDUhpayH
LVV2767N0rTIXSm1GgedqlANoPYl48bBf6fRtMdJT+snlnk7XMcX6tg+fBvIUCqjH2fGkNolIdU8
Z73eMynUQm+GVb3IGvWjr2ZA3JYNRiC50RRfbUNrYwvrGaPkRp6Ydqgb0qq4Ua/pCdeB67KSan/b
MKGBpoUgawsM9gjsPsiMkm+3moVCINXB/hTzcgREvX7RgdSU73nd+6/lvE2Wg4EBMMk9YbGJt5d9
LjyYBGj2Goz8wCS1LZKTCUkvdhSMzTnE7L/Wo5KtuGshmFodHV3gqa/3qT5qnJc/n0OaTHQxNydv
XUaD7eBTEt2UCyPCrAqZzFzl9kHwM/9vRy2jCuGBG8n8lhHq/gByoNfE8eVG3Ab7UuDptvrS+3jF
ydB9ooFIqXtQE0ohREqahczz6S52DPPagLL7CdL5R23SZoeJ7bTvukHOu2PJh45AYWCzFcw2Utr/
qvSJBEm2+Liwc8iI1TkzGWBY/BySUmcig3gLdCq6uEH7RZOs5xmlZBSTo6OM1POwTdMQ4BVlG2Wf
DgcrVjy71jsWneqU5wFR93s2q7UqGzhhMF7X1bXFJZxt3PuYd5uPn9p6roU+PZG5YV+/DstNLn5C
MwWirgsFV1gleakAix91Fd45qtRocjKPHcMSjL/cAVAzILrNrXmHWV8babnHQ+1n1Vpwn2v0a75N
3bjppqn3LsXlHXFGlusARFVbkcEDLMsWw2W2EmhLDnY4myNsy3rII3psrOBp+bdbhXKy4J7RZFxx
qYBGxvu5mT8x3tYaSol1rd5CEtxuHjtNsJ0Vt8H2YS9drR8u1pYvL9qSNu08WU8xfmYFYTj+dCX9
tdWnKLVlswkzcmVOWcv5Rf9eQ/O9VCP9BtmJQ63JDOEJSDTV8oYncdjlng3xvdAoN18K/ab95NQ0
BOfjN8kJUkeyhN6+Tipy4Jxx5hUrr0tp78efYeTw7kxDpZnzHu0uwNxrQxIUxArPGVAvXgr0gofj
xqdLoav1QuI406wtmjnPr7uNW/FcbJhMhq1u+WCv4wBbaIAUhK3o21NrDcmXSr6KUFJS9rU6r2z0
i3vQaolUrC0+PzAWjPwPbBeUEof/nG7FxX3DID06XUtMsPsCoby+iftuqg4gvTVqkSCSCt1F370L
PldG6LxznN1UJaYKeK6wACDs9Pj8IWTwss+G/x5z/CMH4pRekroTNxBDPoYr7a1NqNtxB/guiFpH
COUsoM60SDqAdemCQUzrnlEmtCle6TDjniPTmZhM4pGY4D/lxvCDUvQi0bwofYwxkb00t46KrlEM
IjxlXbBoA/22UAOisXTERp6iOrfgB6sNwYQJZvaL0uTbv5H/fX+9e01qmTJFm3bFngqMWUPvqUPW
XOnOKwGrdAzDmiV4QfGoIdKIOtRu2p+/hakrjS3iNNjSxG93YScFv/rBSsYenRfWvgCo3+o0qZ0y
VM2LyRuhIgcbk+uJjXssL0iZ+GxBokHaNAya47VaBPjiEabziiIeknGjPKfE++QwP46WmOai5BRQ
tcZ0AFlK02/ACMLZ3P8q3weAs5sSTHGtDjKCRuTj+tJBFrvGeeA/WvsEcqULFJNxGNoL942j15qX
uln5BUYBjlGg4dbQ7ebj671qIHUN09lbvOYwzNPW4vBxj66mhfyBEC/estdMagkVAoDv8lCIllda
I1P/EwXekSXCai1/2HkaCR5uPBt99KRqAxmmQQQnoidHZraP5I1EEnAnNTU84cLvVkfDqPpOE4U5
CGSDvlrOT+xEHkYOX/IyravOQIbUajOsc97ttbgxvc7K5Xs3HSuPIw3IyqhsaV2VTHJYCKax4kUn
88n3jNApydp+F6DqGLAYtDJhEcDCL0YPznARXkddXvaLHCahU0OGFesKYuVqi9aCAhnBd2YLmRs2
fNKMZcsgV7DgZYZo0Pu/EHGvr3Cc/7NZMMmbUCpN7TCnjq6nSvh0xw2rbW4Mbij//Yn/9ncKwI8D
1MEH2P6Bn1Mbyo7swrBSFh+rUQ4lObYkslpxzyymrZ09smlPw3UN0iAKb+eSsnU57biYVFiPFH0S
RBX1f0Zhvja+ZVywshk1rccmmTUJzymVzFvMRAxU9009oYhv420PvRaxMW21b+dmCv4dvnSIkLxG
7h7cOwOBZKjaDtSgzq64yE4Z15+2dMeFssdZzrK1g8VIhVRj6NWjWFuNBsat1dx76+ag0BlSJ0Y8
hNG/D3GT0ODrW4cSpYM0rVwjjuTldqyQz9l/a3SabyT4pS4WCC8gpthzaF6WYbcDhdjb29tbVZzD
P6dM/xL0wPVh3Ttmd1SI8LApTvbvpuSQvV7Et5v353Q5HzB6wfYoQl+mnAedwBEb0HrWu7hHAsk3
xS7enQ1U0Jo6iOpU9ylpRi0BWSKLCLWn3VdE7OjFrmALZmHk5J8OofRwQ82ZfsRq3vbGsBQJirh1
Czs4hmdS++AKxJ6w0WSvfGc68Z+w4UfQHx+Pmyhd0XN0wFwrfH8fS1467IaSc4m9I1ZtwP90OYJa
fVd+3eSuj03PNnvsiceZ+OHZFuz2Mj/hGsnvfRigLriVJC6+f43jtQqvgdNcNCXL6YRbLZV2gUlV
BxGWrD2iDvBoR76sS12ntGnV9KkhSeTvYTJWpzDVBfqDaLHtRJ2Xqk46MqLk+QUbD7URE0qBrMqB
c8CEimwvzrhOogNerWjP24BFeJy1x478NBcDH7kTsYiv/AMcI8oKPaQt4sfFe2l6wm8PM5qH4OrE
3SjOOMWcTtIQWmyECuoxJJoq/isdIsN7e1+Ym43VGU3OyYC4Xszxf1zekKmktqSluC0a8von+WFU
iYmk2Fhuul+9RrPe53JT+BlOKIO1d+HmbDQ7WwQtByRV9qA/xyKrODKBxsuQUuaVVhY5+EIfcd36
B4QEvai2HDvb6STnuhupGJmccJiwghnmHNsHQWJi8M6PNI22ZSgym6neDBySZ+GzVWUZEN9KBc7P
ivDXhp1ovaH5AWx0kXAM7NeyRT7auKQlYcMSU8jzS3Z9aHjJtKI3Y9jYZ5YWw99JlydIAAFFokr2
utLI2YmFuKvELmvcaStyfGjbD/vsPv/bmeufuwSLAkz6ambwWjDxPSFrBslp5E+crR3bODaRBa9Y
0OW1lIvRqbwSOx5YDe8yTkhIcl+hK30orvWJyxlH8uusy/4iSiemlqu06i4InbNllNUPozccmLA7
TuzdpcmIX08KvO7Hj8g4UylTjW3ugnAACAmoONp2YJiYetlhCN81DzhbGnFvSdbI7anEQhIZxyvO
y9eyW8jrX3DW7Ybw00d0TX5l2bM7So3mK2H0KM2WfpvMTene0bgAsp5lvVe8gDJ7a+HbOHNiSWs5
E4CXs9CxgWRVkwlyBRmkM80tv9snBGDcBGHQCLyYEv1ZnrKJMEXKDpci0rz3zvYuEAla2TeDgwPk
V+cFilydawd8LDPSo4vYukLnR5pQJ+muqsJ6aOPn95FtRMxNj5xLumRMGh9vD/BDlWO9WXk5LmdQ
cGA9Qjfq4ji4oh3DeYrphWleOu15OsMfysbkgtBbiESm0pzvwMN79q5n+8YkETTNyw3vsOgzjnji
PpTR+/jG8HJca5d3E/JfhxTnaosUIX9xrfMJMjhgj2Jo4YWlpEuDryiYu78AaGiZcbuuOD0X4R3H
l6yV8yM8G2rPdCxkLiCLhILZMQszGi+JjLCeFRO0753wEEy4T0fP1XRnQ1DUse3oM2hWmcRn2Tdl
ihqs12BxGCN63a8XggvmpYeuGV0N2hkdzPpw2r4pMNDiK3xqkrI50XG72B9pq7wbZCsqBs+n/eF2
0owkNMel21bxFj1EGo6G6V4sc/JlumRS5x0voaHgiTtjAONI6sWdPJuA0j8PTN96yksjZTY7DVtz
MQhAvAr0UIr5YUf1AmziOk/6EPXYicGgNC7iKRInZJL2+xTvkiQogx4+ryoudtwjNpgWEALdqz6C
nkEK5+JCF366gp8HkC9kTiMAKm+fwITfC3pcmoGscHbX/QSYKiwfqKXSTP3YZAOihCRXXFFY+47o
yziy599mZVNNAIwEGMIldKs4fRObZM7U9T19XkrjDA0JuBbZgVi21IQka3Rj+MIq8XONfZto2FZI
Brl8JN3tUkFvcwmYcwl1HrhVBETdNZYuM3W3ccuAZMWmpvmiYPZuzpacOkZ7QSG7ReLMPHdQO+s9
agAPcb2PknuXJlUGqFpLa/lvX98Hs1spw498wel8R+Ok2PNMgMstDhD6XdExiN9vOG2hNSgaSE3n
FzuJFucfy6Y3S1+Q7ONg0SKEKEPnmGEh06M4Qetg4XiCQqPq02TIp9+VGgNCdavU66d0vadsSdZX
VyFJukc3VtRx7sVecM8NM4y3zgmafHW8udIqfRSQrSzBOCN8d2UapqyDTd6D8kzmGBX/I+XUVPbR
Vy+ANegunXsc9wxKxpzLeOzWIZfj+eWJgBqTiBdWhodt459TrvwWpi9X3l5gU2Xy+et4PbtfY9KH
tGn3sGpnCc4AYIVqsAPc+Dtp9wfkz25SFXvddsUXeYT++Bzrb4t5Y6/lVxtE+aU6wJkoX2yXqKTb
5gN+H5ntsqRioaZqjUyGLNJAIr6h04L30W5Nd/driDt7dwk4m9MIRwzs/pkVqMH9P+ziPMM5X5l3
aYhx7+XSqAqilZAvjD8FQjRHhVWZsvFR3GO36IOFAKSRdrqS2ORukANzCD3g1MFiidWlq5MdflEx
cEc2ce5LNWEqzkwdTAF/9ym5NYFk+nhtfWstmyE3tzn2wy8r685t5Rpk3tHQGA36Rqf4Eon7GL9y
q2v56zcm9jNjfAv1Vi4bS3COXOjH8Xab4xMHTCLsejAhZxz6sTwMX29blBryvQPzQYbyAQZj10zC
yJu16gjrTBZr+UMv2nDq0OkeM9dL+Vvif5iPU+7lFj2PorjNuFoDj5+CHK4Ey7MbfD1BKHkF4w0D
23kwfZeihGQgc0wyXD0ZA31hXn1AdfEbreVYXVtKgo8ick1aGhWju1EJwxikG1zEQZ0dIuAdCa0S
1UFneeV+lVn/gzJma5s4UZdyxQCK93GbgG47NBGeGQqmHnF6ASLAeJHnUydSAmWVSE1XVq22dQLz
6flNLv97rgNAHDQ0pDKNxxtoYWITYup1XtuDBQLJfC5VEc/geHsxNkq77ah7t5pI/LUh11P+feTy
NirFpfingYVEbhqUoJv0MI/B7BZOLpb5WRThT4lyM/sNyPuQsbUkEflELHDaLlooLWONJZ/A9qxN
bWDm+pMobD9uil7b8L0qXMkJkupE+j2XF4E6KHhANxlQlGeFl68BUHpBvm+Fbog8pfRK1tvVk3Fl
FGeG74v6/DhTJxQ/exzHDQKYsYOqXY+mEnadGIScLVV+HDR/Uoe+NnCakNn4NAip4P6aB9xQ3XLj
m+34oJ2vDWAyoe4oEUDxBl9FJMTP+aVtvuUkdVsgaQmI9hnILEmsx4aA7/m0GC/TpTk9nChq3eoJ
Qd2sRUl/7FXeDxiMKpjeqFk12afL7SpiANIz7xheppFrbcv3AVCq1jdlbc6BYGrd9D7Hq6Vc3Foo
ujyzzPAWtgTNMZ/g4w+N1B9HsXIgNTWm6CFYsq6NZcqC/AS4+hXpK3gnfQ3zNZwQb1SZujic4fSI
qGqYMYZljgkuiJ8RnX5biiLAtTY/jvNWo7VR1NCUwPjAIrZk8OKqjVI0eUg27ovpnEJHXTxdj1+r
Q8KSIfgJJh1iUXmRbjdf/imZpPsM2Y5Oa35tPD5DF56WKRXoY6dgYu4LoFW52Y7HgnwxCAmBqTAa
UwzBwZdCitLG33Xa40Qo3zrnQutQTw4R+rinEWDdhavq6bLmlYA0wM6xi8ZH/SMCD+btrXSkNFOS
Kpj7Q0nKNRb9FK1X+WrQmDmRmkQ79PeO6bA+WY0XroAUzDx8Kh2OQ55ItVnxVMQJLHOzaLO/vqKC
yNsv+F1xWoqoHcrjm/kh3O9UztqUUszbJNrlVcx8lFUCa8g1SgIQGHlBswt1RY+Mc6eeVsO8X7Ww
Z4Jtu/ZGBlMP3KsKkUWNftZ75WoL/m2eW8Y1b+cstGLUskFAJRUo5f0b7OLL/PxI6oJ0sbulIKAe
s27lCzxqt680IkEr5wnOFFzFlz2SbcrMZGT085ETI9pNmg0+NpRpdEBPmFwp3l3YdGkXCUAV2ZOK
5d11Iv5GPGt+k1IQ5e7rVQsfJr90aUybMpg+8m/SPOF6+x6Yl9jJ5ESZdBLVgOk0i9jX7mNqaJRv
BmLT39vwPi37hjuqb9U66l0PCXRBVk8jHuCeV+bRT9PIbAqHI8Q+O+RutlbDGv9QLOuOLhdzaZKc
8q33pDqDcpNRbCd57E5CJSJmrL+l1PySUmd2x3iqlZbVZLfevpG2wESI1b9Twc6l9AADdBo2dNW3
rmCZ/1+mjmUssaEKOKv7QvqSh1Z8rM0hPNcIV++9lrSZd1BlisG+ogYYn1yTP+cwbDgIr5cOzvWJ
zdAvsAa9kIRs+SpUSkLBHNF4gTrJhdN6BN6wF6rNmvzMiGph7pMwnRCFCMkUn27wv9vCOetxpKHl
ByMni5/IAkpwTmx7IZUiJpqhERksIibsnz2f0Dbn6MXmtdNNPeuvKHVJaulaqYrxpwZXu+XHd98M
Aiae/a2M3MaFov2g9Q200bsAmMYKkSTa8TSHMJzWEPQZZWrAri/Q1odOFVbN2h8wEpT0EQIXpDVx
y0IDHZrrvSqJjrOOVcAzbG+bsb2lzmDQnJrN8iTB658VJjK6ZVID/IiIxmyd7PB6G92N0S6V3khf
Hvg+7xPO8D6kvbCDGnEWZb12WDzANCjh/3I4xq8sEE3sQLlNyjdqKrppNdSCjEvf2FvFsccud2Bm
ByhluOWf5BRPJnuS90RRR8TkpLIU92ZzqinrBkHo7bJq8pVn/Pcj/ppvpCyn5HQhGEgJrIVUR9M4
/+wKl6AcN5YEl5yH+d62gfSmO48wf+Ysj9aNT3f7wQaaXRjdxgCVhTtdLKPry6wSwx8dD6PVxpT3
7VuxAWWOh+quQMoBgycOZYo/eukZqtUx4JZmRE6YnxiJkpNnc2wnovNn4mnoeE1VBd+JERBQ4hc0
qSK2i11JWaYrKtsK558E1tsd4IScy4/FwzsBP9cmrIGj90GRJkfPpWAbO1yJrKOGF0EOFB+LcuWN
ZD//o6hCzRzHbRJ7iBMVr+gkp8SP3SiCZqnx3VEBt9/JU2v1ez7guTaaBak0hR78Z8qjtA5EHwEM
GtSN/8VoodCvDefmgHzapNdxtlvFEJj8ST5Yr/PtCfD3xWvqlEjQwFFKtuUcAonieC+3mAGy9wMH
3CCyuDOzrJERyfq5o1wTG2GxiqH7sjb/WD3TBjeV6+4aXnGe1tDUeNa+aZQEUwLdze8cvOabjOAb
ueN8mKSKTRJaMhMx4tZiScECsdV0ytvNTX59gLb6zf+3YzzttWi8f2ld1t0B28B7o5Ewj7pwYl47
U2NQubEhfChGF1MT570qEIQJhv8J2nszx+mqpLA1MAvmzck+HVPynlwmawZY3CjCXGpgk86bDPnQ
rNRDA+3Afb1skXE+9VGX6/UXochol+ITB7TFRLVY79YaIqOwvF2RxkoEHJ7B41JJF7mkGzojctXJ
IhutYIWsaial7SUfN7xoR2/u27w/2Y6ek0t0n7ZWwoKQ3+rAx94Lu9+sHjeBuiOiSd35z7EpoCA6
Kue75tVZEr709SI3UPMJiRHfrWJ67EKgDE+k9U0DiuTnBzaXwxq5fTNXPleoYeJo9e+cdAxPpcOD
11EWz2GZ0JCFjstIP5d5AtvB7qNUCb6cIuZwZtcSnnFFxWnUAuOGPSrZxVwBAXQz2LWxORMgnyCY
4qBYNjAl9kfl0C4zOmZS4NPK9eASTDB3C2uy0ZY+5IXb5PXRzZFZZzbf//FTrQ/RTjQ9Jso3nE0n
EEo+0EOpj+H+S9T+oM/spgAO0S+h8n5Jr1ZO2nZQlj7zWkTvpun+YViiI2bJVdQVCOK6+c7u64/z
rUmLLO1ucGp7HAnkB5DjBBoad9KNdkXuDACTfoQmfi89B3nDKSmVxBwAt8fTaynpc+FVo1uqY31I
uFmLta1Dp9h45erGdF8OQpp/ZQpZj16FjJ9yYu36u8JI39w+xPWxhXdKeXHn8s1ggm+UTDVQzoSm
baoTRBJ+EeXJxzLlVUSvQgCc5ldWhgP5dbWTf7IjDz3kHvNpb9DxtqQw6V8qW7A9dM2R2m+moJx7
51brX0C3w3ARy5wZK40GtYm+UGpE2rgl+OiNhQlUzG+Aftk8ldIr3rtuMnnFBJD4I+WC/Vp7W7Aj
fi+0DBJelZOJH+R2ppzxMifXj4WIciKp5ub0AWsjJIrQR2qqYBK/0QBJC/AMNESPqCuAoaKRROnO
NXRWvXEERZK6yiKRrqCNEm8vmhAZmoWGOsT1ZGGJsslpIcJFXdiUDa2asiINnc6CVfypflavsTE8
bBcr4TRbtyAfbWkr9qssXkzKl5gcwnnE238uKawV3JMsnW0xmKYl4PqW2Vnuj252WOCUIj9xqEPA
rdYmu3a7fmoJpXPTY1Cn9C8BmKcqjSOT1KJqCfTB57ud0Vvqivhk7pTmebofbw3BOHkKhPwTdFRS
/IDhfJrmNZcrzRMXJszcZEkV/EDTztS2aCyPcKgju8soxywWycF8TBI2KNPe+24Jkzk0KcHYEI56
p5P/GYicuMOc7HkRc3dCcOAxXQNI4rsOhhk7wpRVXmIR7y+VuRwuw+1ZbWW4Wqh8zCoQczxHfdoc
roIXba92aa9DxPT6InbvN4FY6HbC94her5zzklvSm1WdKf9L626LfHLQ0OnlbuLfiw3nkoyGdkfj
LxX4CQQ+c4p1z2Olcb/goOcfTKL7vuXCMylg8QmxlpXAAQa0hJathBfsCEJBDaCi5II9s4lqnQ3o
HhmcaQ+oUKiaMOkB5TLqVbrkOULT3pf1yuTD789nC3wwdZXWc6xlWBXlqB5dvxy0ilda2lEvuGMD
0bK2CPMvl8RWEc4OAjWmZ52nZ7VsqS3AgP95Qrv4xX9SUNZR1Kq9GPQUQSbvxqAAnHbY5SCyJMVx
WOc6ZRPMbufgg4e5bKgsRVxz/uQiMJZjp0fCZvTG34l8KPngnBbD1hSnsAQ5zMBm9VbDBFUqGBKL
Yw6tQ9C4NHrpoWClJAiCM7Qhqr1Km6mqIIPYIJyqQ9nXO3ZLcIS/3Ir8+A+UIFU1pU+FSz5jyGX2
Qd/x5+6HjZxD4dWJNpP+VUtxS8Rpsqwgy1E8QcgsgBcuxXAUp0EWVrkkpSbAsyfWLuBzkpOPFJr3
H5UjI9m8NvQT6pOMUoD1KV3SQUQE08KbU3COdYrEPhelcGOlNhMW+5hpPKcAO9xyWC7n5DBiQLGD
5mEi0Eir0eD3APC7Dvt+2RqU0iGHKdcr68GV2UaGB/dPxPPsR2VQACbyg0YAMK63+8WWgOOi5GV/
Zwo0xWnNSo7epDM2MYz254d6Zcwh7xsRzVNfraSGI5y78gZQmi+1ceuj77ws+WwlSG7efRUM7OXP
Ymx01VBvqDnApMzN8TVVf2ypycNjmFcPPH3/K7XCGfYu06wTrxWPuK0Y+vpoMLVZXNH1u3zKg/gY
tklVONASDaztrFoS69nUDdnqeGQojiju0NqhFKDdzjDE+7RT7xAKI0FaKURfFWcyT7lRBlLKAcxZ
JKAw+u/NiwR68IeJGYmGy5skTI6eOmFhDVsL494i1E7Arbdy04+UlO+c/9oLtSYdAy5IhumKkMXn
m3Pkvxz3Rwc+Y+4Aav7OUmaUCsl9S1Bup34ieCz2IS9KG5T74KYlbHEAVnBgLsnyLZBJ1XxhgN04
31aXIqiUdCQrG8IY6MYkdYhZZ3/zkZSrfvb97+y5yf+UAv6eAbnsWC8AYa0eUO5RhrcJ5N7jwvOd
sUN2WUI6MGfFM2yzeH1UIuWOlRzmfx1p6fKh9BtKLohtzPE+KD4xJVR6rNjAvS7SaiF3cX1JFVTF
9aowRoAVwZx/wehW9TvWBb9bidLhnekv00xEGi0554dBLtX4SHjgzyL0LCE/Y6L8Mh8jj45ESgh5
dHKEeAOQkhqCNwpMKgb4rBhLoYoEe43Q3Rc2VtpMLCaX9IODJ8XlLr/fxopI+MMtJoBL3sYfUiOw
smPVyOxvqYqh2iQdqPhOBFpv7DirN8NFGe5n5t3043S/8+NkyRfwVfNpHGMZO8a3x2aaqsvD3osp
5srM6CS30wCd4kQ9KF539LvhIr+dJmg5qUae8J43stfhww6ucTTZ1ANIDSZuoDYu6hg1Gzud2X2T
rvcCQFw56rVgCg+67NYIcnTEVkLqFiXS5SJzsL2nFy2JozP/xUmIX9p8RHDlJVSiFI4FP4syAeDL
EuSCO896kBW7c9YSG2S9ViPj+D5cFY6ORn3oC9zkDpcU6K1FtciRlbLG3E6HO9XLR4WSgvdWNq8G
JwxD03yuHUaCAHyBAgqeM2kWh6JIoLsobkkNo7W9+olJtbznlWeq2MpO5DOaGpmmFnLEFjoDQP+W
gan+0DSet3aCdnqUOt4f2L/ov9BY1wTzbJnuQGi7V65QbOkpiscsEICkpOIUNvDFIaXs+LbR7uE9
Tx8NU+bUF9q0LD6AWzf8DUt2n2bssS6YH3V64aMQ6ASrR4eADUWNeyRcOpXe8Az9xjblwHLF7shl
qSRSTvuldfDwIho2+idLnlKLkhg3RyMxzd6daLIcluOI1I+6ZxPqJcbi9s8kfNRVYxKlSpYmJ2Uv
yyG18VjK16dAZLLqfHqtfugYkcauVGwvBG+nuWolTozqjxP2qOXNTeHs6KKiuSYaAZ0j6hzahN7Z
tVarPYntjdNwE3/X7ZaHuD8wJ6voeDCjdhj1xHlHIeNU3VCMm3JQuqU380SD4dftWROe0lv8IySg
/sOjG/1DkHQfFcWUjNFesppGcNesUunwjCYSlG7XjmFpnOcz+FBAfyqCK1aGOhleZNUMTH3oDbw+
bLcbQdAo0BdZIDZZEVO9b02SL8ULL5oDpIMyAWYonwoUmbwKx12wZOOenqiL0eFzPHVPHO2+1el+
9Ryemx6S1X5ufnBb0P0LImsxO3cbkzp9s9pG7uOda4rBX6+ygw6CT5S/aM+m05QCNvUUFaBx0xuT
iGH9sWOMHTw0XLlSz4fXRj/PQqBMy0TvBVKUKeJQP/T09KslETCLmuGrIz0gYdpyicF8J983j/P0
e7XlY1Rj3yCiYaCS8rxgpkPnmPPHGynGDRv49DC6u7rhmxnTwNzddQVjkSCTLe9vncfBB5PXHTbh
CvAAhwiW1ZrSpL/PxoJ8jXeWLytkroHCZp2OV6c8R9E+UOhsiCCyhzJ/Eqj5wQpiHCuzIsH1wwJL
7OnnQufBKcaEamAaBPThGBUW8CGrxLu1lKYhs+2KV4U3rR2SaQh94UMPX4e5u35x8p/THA+D9d6u
eAeChe44VFgLCXCPYn3Ygzw5FBiOJUP7FQPymi8gGQAzkGmyArb7qLnejejJIqOfIZ9xW8+gCIdn
ZHOchyaDZ3Mr+ykIxuczkcQTMTrwclT2hJD9HvICK69QKwzFbDoix61tADwXS8FqHemXuon5Lm2F
FMWUSkdl3cb9VV+TS1x8bjtOMhRQCoI+Biwupi7hYF4V7k8Mu+Eifq56+Wmo7PciQWZZ1U2GltQj
zqxngPp8jGViYlEZNo7wh6WLbnZEpwnAs6ZBh7SsT2ouNsSLXOq6z9sphO1yK6HpH/HCMwApucPr
2Q7tyS4LUt2sj7T46FQ+c5beXaAHaQvt7fjwDzFAdZdJXPaVqqCBHfukViSHEiBowjbjnMD0LjxV
lhfKxTXD/Kp9PKNrVP8FKYSNAB6IU3XFhwe86F0gKQGYADvD0go9mFNslGZ6M+VUSHonDrDU/f2Z
CiQnWbO5hOQy+I3GqLuADTecTCAVWEXEydF3GgEf/y8Pxl9Zm8dy45fHQQizmTt65Z7P9VGxKfst
4V0wbXdO2c1h8CIiNIKXKVge054fh60fY0v/wZbBk5ciwRCZMDEtVUW0dncHTg//m57pdjoiGphK
bCR9pyo7cSn2wVmyFMmlqdaPAr+u6hZ69Wbd8aRBXEa8ygkVOnLYpJyVDtllloaMKmDtl4SCVtVb
NHOMukSGWuwYwM8AtulraoPm6Y4U9A5atrrr58l89f9cFp02EqRdBDapjiYr4pXyG8g08l3HDLsC
mh568jTxk08ddnvGKN3ASW4KK8i7t37ZxN1gRXEaxFwZH32Jmd1fxeAkRafE9DDI6u1LPPldDb/J
bOHl5pa/lPXz7z9cUc5iWC1wmahXXa0onbqzkNA5Zz2c1WkJL5bC0BjLZXhXvsWezEQM8Yk+0PxP
+o0NlmjxDQlli3jU9vjAS6e6zPhbc4tBkDl4Oxxuv4gNRslJ/IBloMvedvph38o7hbmd9wvc3Xy0
BKph1aTlx/pQ6lKOqVVAdngmtcNn9KCEjDVBDVhG1NMnmzMdD08n9jR0ObK+1gv/kA1mDAfDXdn8
yQ79C89zfrmUd9Tb/1x0CzbB4iAMNXaRazml+rci9zudAkocJLyFCoYA9t3OCtx/Oo8CPTtf7CeT
zDM8jb5lkLhQF1XxpUtF+h9hzJXvZMq6af7rimZXHZeIBHlkRiGjBFCYokHU9FGojkpHICVU2RlJ
kzkRW/vOY/T62be4IzFIwgPHXDx9/z9e0XXUk4S+FX4RaIDUIGbObopHPEL3F7upd2kHRZjexn/N
Ok1Cc3fUO1HwzVtJ0rut49PajI0mamvoLeaVCA8wloqv7I/7rdanyB+JD79df2Du+4g1NAfDqf7d
0NpKwMZObIoCwYrVtfpuSPvHkAVjZwfE1ZxDC1+dcaNqZqhLPihWpWe959ienpWDFt1diOl1uAyo
bC711qSyMMyrnKNCpFu4EUE8b7J0eKiu14tP2Luf3W1uXpisWLUIoKhfbU5Op7OgfyBhn9UdJv2b
SaxUbNm8+eSd6IgPYhrx+nRGSQSLi8HrapORnQfLFYSS2O4NSAzirColT/sUkPw8rCJIwZ0StIsm
VOJtoagatfYrZVhwTTCqIgwSuf1YceOwYC+43xC9Q1EivuQ6yagcTeTB0gllEuMElijnWb4TALCX
idE1c7WBK4yYJ78bn/MSut6jBdAH0M1cWQqVMiiQEGnylKJ8P3071KRbIpWbwQ8qj0S8TzCHPqv/
QN9u13QvV/qCOCoYNpcSUjRV+q6aN02Nhia3yo1XnDueIexfVyXajonOqao+wF7goCs82eiEyCbi
yBbBYKJhcJ1RXHO9kgcBUk1xquBbxOHVLOyFhRwzl5LMfhM8I1Y6lqgg2upIBFqjEv7/4+hqXJB9
G0A2DoyFSKgzZ2D590k5E52CK2wPUCMHa+DAhpynC7cA24WwyFPhzyqOhVe+Kw6Hzhgjq4lxdNyZ
eZbFyPDNVjsJSrtat7ndaF4R83trg7xyM0c2kZ7CpFXG0jABLLvDW+/S+IzQJCPSeqIYZHZKPe2Y
Yjnr48QpBZvzuqNw+9v1Vqdm71b+ESazhWX7KtlCcagsWYgQo8ZvNP5VIga7dC7bbkxb/g2ER4x/
+LVWWXBFpmz3iIMYKTFBoxmyGPNPUqptZoDbwiavN7ZrtuUH6wUslCJdrP7ObVQPn5x/rUznEO1M
n8PDnRGvD6EQui/prBQrBq3WWgmqv6tdgRU6R1rH69Ruvo6n+shcgKFXHoKeCZhP1EsukLqFK/JB
PHU1tc0zZVZpXCFQxX2YLkqHP0ImyAzHIRQqnhPSHMqs1ebk4/UI3VtNuLKiPL4I5PBK0sv4nVMV
BW+XYaxV1T9oM2e0mr3q0cx61mLu4tFUl0ynEEvhTTohPtfFb218JPqkLB2mLBq5uRupmVUxCL4q
I8ZehkT16ehy1pHZCs5SHQQbZWs0PeuX07EoQl0HzMfPeRvEJO9QBPF07fUqzBI9RKm5qi1omdAX
7akUrHashDtFNd0zYVlL6uw2WbGAjiCm02Y+XeHV+9Qa0dWY6rog0nCBXXc2rN8aZ/htCyhk9Ssq
jmMapW/NOXBYPImVjhKUrQTRlxCJL9JurHJcJZulOTlUE7oNvEfMPrwXaAI19cQtuf5a1UpeNqtS
iBoJ4mkbol0UQ86nMx6UlfsH5CIU/o4cL6gQQ8vU8emVM2npiq/UPVP4S0fwswG8ddkO0kr2gHWu
m90JsawlS34CKHQO/M1GVeUvWwKS0wpO2dE00Bz8QsoDrfiSGId78z0IJmWB0a9+kO60QQvOv9uQ
SipcPeb079Ctp/GJW/ZmsfBit7oYEokGtUTcQ6ZLIie2mj4ce5jaqAik2OE/6fxLTSit3mz8yVw8
yX5luzUNIARGj4QMu3hB1nQ2iqK8Kb8apD3yqpGatFDCsx9F3XeFsd6oKR0M+LIXzQ5jzl/B6rfX
hFxcfFy1DH/dBREKdVVTi+ik9ohvAvafG6gl2o0aCLQvAcbmcg/68QHDQapSYhslPulAeMKOmkJH
jcuBbZuyEzQYzR+WhDshICsrspC+VNWlXv4vOF0Q0Mt3Jwqe7mriNW1G5qElL2Gp5Ala1gtJxQCy
RsX9ETYSiWYb781IGU0I1h9I4WbFwo+RZfIDEXZF32oQyxeFOjxdTDrkn1qRpT08QkbKE6K22vBh
tGNWIfT+VqNmr6vaaZHINewTjPiZCPYI5CgjwfQ8XtrHBbgU31NEp3ClgjFb8DLN4ePCL2kRa5GV
9bx0UzElvnyUAEqp87jGPTqDl61XrAE2WVWfYvrkc6p3QX7SaVt4acyapSFRxPAoKDKNFyMiLfhB
HbdWPWKQSACDShrxD+/KZ8peyAYUk6Ihplw5PJnQ5zQ1dp5brL+YIHZ0BLsPnKhYiFIhRLNjTyhU
jEy9UR6fmfjrBlHHF1OotePDp154CPiVgKUryyv0VPjn1jDPyza/een/cl7HVPdf7xgDPhm/pnaL
gLfO/rYT+wpIN+4qz6SYiCiJT9+XIod2NGhrkv5vkKf4zL1YYacEuX7MQWtWyaaUDraSNVRLkagB
a8Jh/SwWPFE1oYCFf33v/W8GpSG2L+2Qao2dVfJoDyQg+bYstC8VSf1gOSih8yUgsvwKlrHq3CTB
had+vT4dkgtvKWa+Rcx0NhC+muZxYbOV75ouYi3bV24jNAtXTMlaj6td9tM7cU1D3wVDEJNpWDl8
M1DzduyFZLT7ueOiOQ3oC7adgUkes8aZnVns9xRTimdr92ntVDFKK22L5TYhza/hVzkHuPieedA9
nQGB8teBxE3PYqCcRucGT/7QMvHDopPEXYLHDllWa1znH4fZnx7g5Oszc+oDyTjKY6hnuvIdeGUC
u9fYeqPncPqsHcxSO730E4BgADsCiVm3zdFJjmCk/s7WZW9JUEZk4p7I5G6MwYdD2vx4UG9Xz/fu
ynKW+AIAhhSDAHr4LDZ7T+iOyv43RGbKrK7q/njyBbaQ8OPFlM3UN+S1eXZKzG5bc54hhIn3Xfts
Wo4zfBTeIow7r+OpJ+/eGRKJItmCkPuF7iTqDlXyuAne+B3y1WKXuIlVRvLfyrVyX54cAaOx4aaj
prUJNTPHK6OC6K4DSLnJiDa9ek0w6qW8Wp1DyXAGctHzJwzCy4xbhUP9+nETd7Sfx/3cwPCRsVBi
yvTquIMYNeBOAl2q/47RMULiIufqRWTcpcRBAZvJYFM+7mIrNAPw9bPaUgeRxT6s9vHYLOunxkXZ
67TmzR2Gnz7e/CDgNQ2sRykFwAyuYEhxYQVVlTqtSSb8oCrOCItnNWD+U52KnHPE26cxbqrLHanB
IMcL9J+bF0+ADY0pzBXdAZsyCB8qRPaGaHDjDwHFSxGkaiYGcSWocx7mLd1Or5joWQ3fEct63dYI
7PaKYx4XFOZcLM45/LUm9Ztwc1qzt1XZtCLqqgI0RLiVwn9sWV4Q2vMtq7iWipzG0qsYov1YbBya
3bDmPiRgT9daiY5HquauG7RD97VHZBuNBRpMFutX2DVsGjBz7nLWMDEOJVb0jSWx8WRUjhzEGtgM
SOnKsVKHEAPK01py22re44i69jiqK0NvUTBNSHfeFZCusCQCtFSypVTmaBuuKGjYiltDHZqI4q2l
bK54YB0nDFUy9rWgdY1H1mWJFoqyGkBEo7iivdfjt8RNeh9xzQyUpCISIsVQsXwFuQzFvYveLNMh
k+LAE9bEpZbRGN/wI9ge7zGzfXZYw7n8XDynDsfyjP50QzDRb9iylFBQzckzJxKHiJI/aDo4jeHA
7ql7N742kBUNXkt9lWtUsrFI/VLquxy6LcN55BesUEVHY+qdw2Rimj9TlwC+2RVoVgBbDnPmU8Rv
Gc9xiLNdJsgOVmmlHB9nOGjFTUSwWXl9H9XuZsS7nd97HvN1HmlWB1ZlCu78jyjllXClaF07ioEq
iU+wscowwJCZf+WOyTrA1dM0bl1N+ErxzjEm6hHMJQo/5N6JMxrgc7IhnQYAEtTK6W7+X8J+CAe6
uQhnmYxQEWNgm2lx0oI/jSh0HeYMsrl7IvWULL/ZGy9iA/RCUO4XiyClqZxDb/bSteMgGJj8S74f
5TAlEAQDfic8VQasQZLjcGuEjSn+4xdZ1s771orh5s4PHZ/lFflKlwidsrMmQiE7IUV1Oz1t+Ne+
vsLePno9JC9HTgSqBHEDadCD20owXtbmql1uOe58NaYRzGCwrou1p1490hr8OGUSSdVYvhbgSTby
goamqnr4C+XdAoxoPPA2+09uUmFMvfkCMPKDcBTnUSR2kWAiB2E+4CpNniU+j1X1jb5xXEjeI8iX
+6TS2va5NyazRECn4Rl+QwK06oxuBj/HGhjrUKDbHkgW9np0lOKekrDt4caAJF9YDl7UkXq81h+4
7gOZBXt9n6rJXYyr+1vcuXqxknuPwbbq4xOdoMLfJxTQGs9v0QmfLaeHq6ahQQGY0LhflVN+rRnl
pRmRjS89G7NvFKuLrSncNk5VJrGjxyDRegrHVrd8VwPVBX4G4KP5fNpK94AySzqwHvyqcKJBXpnt
81GW2lmokwuAHWYp8hqM7XR5mZTTUpBbr+KrgwlwR7x5RkAXUdjzikjmm1n5oeBU9GDL0RdQcfU0
5KXnjLjtYRqQBM1XlT8JUVAMOK6IHnwiogstsaOE0aSWiuRga2WbM7BYwFjm8LM+ciRqh3jiBlW8
wSVVhWrmf8ADFwMWkwWVunoK75Dg94Zvl7BipeV5B1oasy8LlCXbKh14puZOF39wzd90oPQd8Si5
T53zfUVMjjMku+/Jp5m5yBwHlpT1jM6ybTbKh99oUEKVidhw240wTwwNTJ1wzr7CSE/wUdCeZmqX
CB6bPNvf4f9MySJ0BexcM4r2ZVHmiEFcZBgs0F6r+cWAD1+bE6N+KRqIrceEl8iEx5MAJ1AJQiVW
FK30Cu73RIXJUfHcMrpVtctprKTfCjTzGz0j0UP2zrlti6oczB1U6U7OqqUZpo2a4PvUQhY245mj
mLclbCMfL46rn+HZXQJRlNaMjrSXS5Un00WuGa62eI7SZer/GBfNXiFTtY8R6NQPvWt9SJL6XKKE
QomIMfjxOaBl/De+NzyqOhb7VxZISq0hKZUb/fA5U6j8mhzdcJCos2+66nz5AyVZfnfMZ9yPKxsO
hb2bXDjJrAF/MCv3D8KxXAFUAV5NBd1JUJWc6B2iLg0EVHj+aMfJxRnmt23y7kw+VJMDX/ynJFY/
Iiz4hwyPv7R76grv8AU+LIUxx2lJ7GETvm1hQPt5TtGA5qrBWDIP7qKOAQXLrZVNU4I06WSOdnq8
lxNfmgpuXKiDtbdlk15rl0/EtZMgr+9Q2O9CyvlTqNf5+SealZgZ+ZBepUeAOKT3mt95AuXTwnK0
QkkUB6aAXWvVGswxgfu2bbvjdBADxrXCbur3pdGmnc7gHwpPp+3t5JzUOecfsdfCR5yVNa4VrXDP
XhGIlrPgEA3JWbymzNPgtaux4t8BmbeNxHRGnpxLrxGIje43BokHP1jwAEkquRwaWH4B+RDCk9ue
LzV3JW7hy1BuvpF7oJlbfq4gkJJqYr1QCRm56k1Vt1n0vL/UoTgq9CUznfnhW1OkJsoy0aAmwlUT
tVcqdNCllSsLEExGnfVgnJQQiaZX+4TeAIYvuJ/BmfTzGDgJ+pzTM0zqZaq6XZDbIYvpXoq/nMH/
QYt1ek3w0fi0IK7k8uclBqVEHh2VmmeEqkp3+jbK2njE4hKEzyspIpCgsScVnUSLlxhOclLpspGL
zJacbefPRFKKjkvqlShixyOPcZ1Dj8BnYi4CwGq7FBVQmClVjKvd5e4bfWbUpegWyr1w9dRMEPvG
hXHB95ELovgu/QJXY7TpG38N9T3ud7EnqnvHh1f0Gb9TF2Rjb4lWg//zxneXSPdRKEeGCPIQxM2L
AMYuJkhj742eynKBlPtss66jjIGyLWJoc+xwXGYH+cE1z0Vmeu5BO8q4oQKAoRe+iAxE+l40/MDn
WUdC28p6EhfC/aPqPfZW2R9hy9M8+XZlmfoFhjWMJIfiZJmESgyluzYYQRgOGwdD4m4za5jTt1wR
Le96byqT3Vx+3svoSuPrv0DFN3qPbXlOWSFwSTNXtjAKO9xw2nqVll4xXMy+yV+ln95dOUu+Orc7
m6NuZAXOTZgEgQqXAsilTuzoUhPAJy069Jd1U3WqOzPZurcQlnG0Os8puss8OY4Qnq4ZRju03nY2
KFm1rW6/D/2fKSxBlujJ1KHCzziXpPPYaA1We6gMjzk4EeWkXw3e/X7dRKehAJm2nLTBs9eG47t/
jE8EWmsmdqoUpbIug4/EybBoS5WwOjSkoll6lEh/XUJIAQWO2RvaAbdudSHwQkfPdL73oP13bT+9
KSGkQ7ZPIk7xbtm7UPcnpIRmycHQVFCkNom42Au26CuIlEPP4268PMyu/cDYyQwUTD/2fHv/k9GO
7GmmbxnZIokeOpIXGEwSMqcQ6+tqOWNljJ4YpN1jTajrpKphWDd7CVIK9plq9yUY434AXlhSIC28
u95TG6QunNa5OO4/53PjhfUX6Sx3MNTuatH6/6Qnd/h8K+PqaDbaHDFksgn34fdrT2w2u9SuXVnt
44UntUnSLM6ymsxQjut9z51W4xmSbgKoNXvU/WLIBq44EuiOn2FrzjUxPx1Jr9Oht4xhMPJiWVOP
P50GIZK9uYg7z5k6JYL/Plu7N0+ajeH3lx4eA5qrW9TU6qiQekt/umB6xvQ14DGoJzNgTFC7j7VJ
xet9UcmxjOSOP5dO6fY8UC2599KSXLrJi8e3Y4NzjuSPxl0bDiW8pIz1dvFSGkR7ZqgcsMxf6apJ
txN6AqUtNfHAD2oB8MrFvd45lTOepNz8A+r/gREsNLbdXRWecYQ6TwIkFSLXaQ6rnYhvBKYYE4g6
TdzoQ1SA4Eqw/f2g1vGbSL4e4nHsuKAuXuYtGmR3m2bfw5mG4sHWtvdCUCsHQCvLGb1Ohmgjh/o4
wQ/ybaiQ9SzFcmfm7+Me/8ZGbGBwzGG56FxR9wjlXH9NMzmfw2afMzHobzL19BGH83hh95eoUZgk
mrOsv4dYHWUmrGifIEznoI4JheAvP+u23eRYPGS6v3JboiJLInc/M4ly1SY7yKjLNCBeMjbh/q7c
KqrykZ+ZfZnsOKM+cz1RlFL0pZ1QJ1iMz+LeiHdl1rPCQiSOMauGmHjeBvgGgRjSxgWHkFO27tZo
4jK7XbTQHuLVlkg7WOgH+C2SafgVIL4GuGv6SzvGYv/DpgtkVpLg09HCaX1JYE9R1iJB21MKoPQh
n+7oAHnlLkBLrNB+aGrf6oP/cyFVAj0c8+zgObGiH7fH7l5qkEbEIk7defbEhHFj3sAGNHf1G7qf
lykP2OIh6cumVVGgoyso1V3XfhHe3wZwgHcPu1NB7pW8zPCgwpnEK7/jamKB20L5ZGfrmDd9Vg7O
o8f1/8E+yzT03NwbY6P65aDtAqSDldtnmM6/ike26YUpfngQYGe99n1gCunQXgUNU72XGWwLv3Aq
pBiRfWzUNmH/Hl3HwHMg2vjmGrNxF9WS6GF2iYF/apwM7j8HlnTHE2WrxpvSRiRe/valBxrtAWVV
MQY9257vuJyTVhvhfvCH4pXMnj78HhvYcfbsS/U9wMKEYQvR9Qs3mJUZ++7JrhfraIdeSawLwEp4
uXG+tVI9ssTmn7UtuWMKgpTCfvA0ebNRH5qGOe2MWWgmgAWdaF1wlgsb7dhnvk6CIcCOBWdaCusp
QZ8bUueTTWa9BHJdEJYPEUS7bjKzBSdtbnVubCD4g7uu59GwMngVwLGflvdsn2gYb/wtTqIdEzC9
cs5LDHegb1pakddGNVUn4Duk81CfxongTGR7KN0UbFjOpK0KJkPTSxGwaGwzT0CKYvV7VZFBDKUo
qVBpm3KsGHFi6kVdn49SCCwR8Z9UON04b+bgQ0BCBHsfXVD+sYGI2aha+tJEl1fkZ82EiSsW4CKa
Qcx3p6aZgNwLMDsGOuds3+YSqoIudv3ddYJBZKsX6u6BqIDui/O1Nb30ZO69PO5exhn7K4grGJE2
u9KsJHUXrkhpzL1gSoT6A4ghO/d5t0smgDNFjio+Q24KmA0qNYd1aU33jH4BnnuK2bO7ncdfmVqY
8tOKu13l2kOBEgKwp+PupeGmgd3ZH1dl517TnLYdO/7ZiOU3PGojpAlDoa02YG5GJH6aUynZXoyr
zbWBpuQmvVb6F3pXEsqlx2rlzL989FqLg+k35Qw4PEcBk1Hc8slIai9bIUtNihbD4vdSjRzkIpSG
cVAbyvz4DpOV03kCbegmWArwpyu8zNgRUEoUnm2VqmNG2ODzhl5aIWefYaR4o4m7kzyPBScmm5kY
lR5hLxWvCK+CS6ih9/HTX62v0B4j2BKB0lNnZaKXA2eOr8b9OsCjawkX4yYciVEir4FSMU6xeD9c
psWYzEfaYHBqtnj2zYT+48+D8LtlDU3KwVpG2W2EQ6DbvLdhHJWo0n5w07/ydmlP+RxEa2TH5AXJ
i47Gqn60W687X/h5KzQDGzQo5CG+P8S99iHFwh0YKJ3ybpf7dv1vcoUy4mAuj4n1yFgsogPCtmns
aYGrCHqf5syIxdKj+ZZdQr9PubC1zIxVMhTqBMd/E5u41DEm/wrn9lmOn8RSUyna9F10oh992lFh
vNq3XKcK7lHXqVLYW07oZnxvFf7COkw2apsWDTRsi2YI/GNXDLkI6DQhhvZdhcKaBtyAN7Ex/OxL
Fj1GHQZ8VuW+qT3xdI9xrHWybJKgS2YJMRaAfOiT1UJKXCM91k8DWacak27PBifWr5fw4UJEEgZi
T8bCxeAwBNbVbp7Gzk0SqwNhzgaI+N/SaV/FVxk0Ac/Hs5ZA/Wuig5SJyhESV4oxZwHgFAYyzjur
aNn3GQusl6e3qzOrplwW1XW9zV+PTY+3HHwamZUBhm4YSgU6uR5R5J7GCW4PFDuGnbhAxIkeQkzp
8zWWMlZNCPxyy4x24EMNFWUlCOVUUq1s3PcH9+pi78mn4w+/Bb+oyL65KTsvp2D4XNQ9nPNKmjx+
VLcyKVwT9tvMgI/4ux4JgS8SzAxpiakBCz/T8ZKgAWfT3DerE98Y5uJkXOihEv1ZutVmYoKQpY2U
2mSOB/YwHobQgwxwDUoHfbdhNVizvWVPDTbd/2Di94Jo6Opl0+ervb3cqfzr3Hn0rNVLtFEkGk43
0eLKwyROUj746f1VLfG5UqNbgFT/oOLfFoiovbjneULvLyHb3x3po0Xa8JPuoMRW3sXT/XP8WcmL
XGg4mIXKY3HDPZAFfKQ7PFaTseOmDE2P1As4wOtGdn53ffKzlM/JHRYpeklKANOh0WH1t+lKJj7V
Xsr+UVqiB+Pvms7kvDrc5lh/BAQysDhx5o1ApklEADrLX/eygNf0n4ldeqHEGBP0AygiaTVi4k4U
O0FmcHay/PNeg0XhVh+A9cEy1q4nxIgHttVgg+QtBXH2WdNLNJmHjf7t+Y+MWbbhuYEwTcPj6PP3
gNkhr2qxx1tbH+BTU7y9yyexjXQaaKX9KHy1XkaiM+aSsn/4RJjtsr3E8xCRGArzGf5D8A0H6JY2
fEbCi6Q3RhWnnRcqaB6wjBBmUSLPAXu6mq4yN5igxez7Nmzb88SnBRKo+/Bh/Y3/1M/EO148jI8V
Bezu/KVz0irGpo2b0b26hCI7OPjzmPts/CP7ThwfKL9EbfcisyNPbkt4V1xPFe0BqIcHyJm+P4oy
qj2fBxTiubuCzVYi9vFpmxnvHE6FUKboDzaKBFN56iALv++XHdESV3SbxJbZdMSjkdxILH4AN8Bg
qNECN/P7cB7mMFlqmjBUoJ+e2nt6yD04FuEH3tLxmRtWhZQwdX4TQmdZmkxBdKbYv83l72sBD4wz
ssIs3B+1Rwt+8MXUgED5ER/EebEEqWksjtkXxrDpVbEr+1BWBuD/o9+riN77b00IoP+yWGwPdtzI
5mwDuyk7PI0CZThYZL7JUU8AXH3aD+mkZp5tu+I9xaEyvPpte8OSnhsk8+X+WxiYRZN7jLzBBs04
TDTXSThgGFF6MgCXoExteuAWfPhbkHiEvtm3hcYrrFk14pfOhv8//aGrmiwwSDygTySTymukjD8A
GF6Js6n6wleD7plChcm0ShGactmcUV9WY9XdZT33bjLvmem679umRttfIIQMraY18hQvV/JlUzoT
EXY5lMfL/1pb6InKUzr3NMVnWUG5qgk7r9GdSBqdDr0JtK3iTyl/U96P5QUiZIl39K1e1pR1b9u4
tfjHgOBOaxpRPXRj0o0H8ZtEs1HLIEikBmKYUFJqCyhoqzCcy0VeR+JvreMJCHSWUtu027RSRmI1
HtS1+CIvhPM56pvGBll1CWqhHzNmVJHqliLGiD3dHC5A5rQ3j37L7HGdFSNu5WZofp/vbwHwL6PE
IEqgWBJruir/PVGBqh0Cd1lp3ncMy/l1gF49Mu9pBEuEtRwXp8LQLQnZPr+v8uRBqOP/c8RZ3pS2
8fsg8rIal6pHXIgse3eSFRWJndYTdPJ8mnTygbChDQ8dDk/67Vxhn0ml7He19DRnM/rH9nl5UWY1
Yep6rrwn4BnkoBjk5aQ2UiVExlv4KcX6DzKez4a3f4zaIz7i+83EwnJtFwbrpz4LETzpQumQW/9W
DlkaBHg9eH8yDR0ZWDvyA1/LtSDjrV6tUZfPiTgxSNHoaHaXYCDiAjXc1SBMlknKPg54VWBjFKe8
T6zeWoda+CMcE605Ul862V4edh8m+9aQnRfq8OxYlNJB5Q1lCsm8oeOQ+4ECzGu9PwBX2u/UDJ0I
tOUcpUOlwK3+YWUOBQ2nFRphdQLZX2LRbJbo8Jg0gzdj69qT/xYKIx+hcWcHT3HlZCgx1lIRVtnw
V2iSwnJT6rl20vsEHIDaxTEo6YqwO+x93qMR5m5Cpggntv5+R6MlIwGsI8J5JT7kiXk8iI4Pr+Ho
ovhsBLCE44gEeDMjxC57eMbkt7KiZ8xghtrgHiUJnvBVSouRm+8A5Rrfw5PJFGBF8ryi49S191zQ
Q6ojXBDraGgEMYjYzvG1jzQwDOKAYw0We9DFP6UUYw/fqGP6C6H2+qdAVkCcmcgbSdz0KHfeyO2g
rJ2VSNzUoi1pFqu4/pbO+PMo/5YebHW4hXUQpHecQkFyYDKYlrbCvOomqTRe2zO9XY+nnQ3d4T9y
SXNUaScD7GVt3P6XU40MUHHcSQ4jYe8dKSJuGEHvbhhtcfXJrdr3KJ/vmXKvRi6j/g0V5ML0Va5o
mBgOGuAa61DsJoUv+VcP73Xs/D4kxlG9Cr7QnKx/KFZ9sWRH08t4u2oocXrxd71GxQ785innim5n
B42Ym6zWPfu/CeYt95nYEY/IRC1Qeg/xVbcpBKdf4JPDKpSJT0SBfZ7/2dNv9jf/WTzN5OnANhR6
Dh4DT2fAIT1+EoeYDpCWDoTYxHESnf65r+FNRMRXUKTAm4C6biBCgK4Rmv1RKNRskuR/3UA9TWcw
E8hPhBloIwUe5hQt75Bm6smGv2nYqB+nbkbQhp09dxM9jYdtaWY4R+eMab5q1Wzj9c9WhhTXGmL5
eTTK2kDJDnworfQYDq8c2JQ1SLX3UmthQq2/FvDAOemDnlKGcFyiJzzFPEZvHOPuLmdeEw2aIU3z
XDixKCFbX5gqeniEHjympkALZlaNbw+3KjmPZ6ntNB1CkWe4Z5DTCt18DEWpdDJCC4MzNaY2sG/t
N75mT/Cv+XZl0i6DyYsxso5CHtw9gTwdBLypv+EdzBKrOuDU/OJrVwGXrhcLAnVpmFt22kPQ3h0x
I4r2YwBkvN66tuTkYCV/0/Eki1vVbJG9qMIOtrkLYNDIAdH3lwnXMiEmETRgPVakJHpUiid7ZuEs
3dTX0jPEHGDZjxCvnA7zqXWroNPgGLFKXlOk+CsWqWEu/a/8yQ9jB4T9h3EPBlGD3y+QOsECc2JL
v7LBNSK9MwEY93O4RZPRATqD9ickRq13tCSVlotOzbLceqY209o2hqRspcMxckYiyD6ESja069Tg
fo7exxqUX83atRvuNaQwXDpJYQ5zgR5j1JrWhmDoVQjTIwPSA4q1hcOssdmqeALMCfc3BaqNMLYl
xEjcdSfEHBjb6rZ1ZyCvT3tmmOuUQEuh9ZT5FSkdqWIEYKCTZBvpGfbzKyStVXwthtk1CdQ4ZtpW
I+eqaxwXxayEqNc9PZdiGb9dJgI2PPMgjUaCkOYNvbL/ta894aKP7uexdK4cw/DR8x6T8kAcytAY
cSE3eedbDXcaa7xLDYj0pbWsFwZjlLz2KU0zbXlfVvqWbDDsOyuWJ/Rc1yQCooxSYarIbiazMGEp
kMgbUDVdhnaRRYLsILVdiocb47LSywiSpNi+GhKe8PZgjI1fE2WiKXBFldSdDNwM2ICA0nZwwzbV
66g34xS1UX1FAmhwAHLyqEb1JS9XOBJhgDOC4xBkKTtXjFJeO8X6YsnkAkf+8vN55lrg8DfC93GL
9bablOG87eewL+GE4AkgkE7vSPIRpOINLBpIO28g/WDStz+Sk+He7TfMS7xcC2GN6GcQ+3oY4ygw
gpBy/7HATbZilyv/al6lWAJOonjnO9vo+pSvomUb+3JfKw+zcu4tCVZ4dVL4mQU46SOvfoTm+BsZ
D7nB1EiinwCDedhQCuj+ss0KLLOu+RqDKwAWal0Uc2kdyjgYlzBtCSZve0Pi6pUgNSNzr7c+uvR5
kIdMaJmHO6xodPPZkuYcOJzWvP9Y58Oc+ue7NCkg3aiWMFl8lJQvX3zIGGEhvzj/5gY15Mh0wFTl
onhcj/eacHmPGAAZskM/Qd3JOuTGWaGYtVQYvtSHAqrDp8GWULwczQV+TQdlVLyfksC1+vXDqBNE
7vvsb5DOnOwQmtgJhnXcatJD36H+mdPr1mFfz6Ey0Hw/d7cFOhHaApASLUyy0Qk3q14in+5nTMih
nXT6owVodG3Lleq7HL7+7i9oHuj30d3yYShfMJZ9zQAs0zp+E87eEP9dCbUunALTZAbSRbZIukwq
yEuhlU5p08rk0tJI7G9lOrG+XEzH2AWTfPRfNFxxqrz0kBYHKhLc3eB89dzNS56NRjGuSwNsBXcL
Rt0PEvWoXeFJ9JyXaKxBGT+H+ILACrHwpUyB/UqRIWc/LhV/VD95qKm6frTxSn9dK+ZZyyylPjvT
7I5CtlnTc6VXNWRNL8GFuXD/1XSq1rRe6FDEIp42Edyr9Fc00K6YyqZ7iN6y3V11Vl8LFcXDbvPr
aoRUKvtSi/ox+DIT5b2WmTBej120ITslP6yhA8CIPEtvmKNmKlQyh+veoP/mpunGuVgqo0RwAwM3
qOHfkdstNzLK9gMAbIJ9uTQCeJxvZT2/XOeMYqK5QIjF+DLcGgAl9lVfmswb4A3OjAlSSaj1Mf6z
n97v18FjMtJR1xyl6j3AFtYglo+l/da4kKLawGMoMO4qL+3izfpr+xST6KKXW+8OW0YA1AVtOgj9
DJsw5XXL78m4wMxf2LXH+o2n5nxp2lVqIMc75cc4UsBoi4C6Nu1qKBpI2kZicUKm5q8ma6JMukm3
0cEK+93pAJHa1jXmT4K4FcXtHXG67LqIGZx1DeF6fqbGOILjjv4yWBIfy3J/uaJi7UGmnUT9rik/
za+nogjXQhubBQuG0K1UGoflMXtw5Y5ELELirZpeTEwCVUXy/OjjNKFVZCEpLyBsixHvELxwvwNh
kcLimwLV6IBzl82UWVIqHBIs688OhoPRbdbAgDxpDMn1NOVgMz8AWl+70qW2zRSxTxWDuSz1B2iM
CBMWmYXMgeUNw1l0VSjD9SMFwu7TKgsRUOmt7+fKYgViVonsBvkRoOzJyvAH7sxoCUn8qSQC1Jb/
2SBb1vq6O19tsdyAAtBLblJjvLuRPFsikB4u+4EAzJM2bWLdOMCOWiFqQulsTHv9aQEkDz8BNSHC
jERegkp+sx7cNKihS0ym79kyh2UFo9OuJm3kQoohkfWz1AgI0jM4PUDu52TyycN/9SgZ/LurKXSa
YToVzS3EIDmzVPlv9TqZ+TWB6SH0ok2TOqHKZ5y/VfItdwRzsKxcLw+AIf5r7lAHuSjECc2sGOcP
6QfXjmKiwWoLR4FJhRb3socrYr6oen4vfg3L2Uyrgmey8Z8tbdz+mLFQxr8pwf8VpJdGAj9KvHj0
9HvRssrlvbVDeEjivgvYTM/5cTnpoVLcYt+tKCrpeCxw/4b+HoZwrzXoFbSfEFwBr7gu5MO3ryHg
YK8Qgj07xfPygnthdUWTjG66qa8raH7J+Z1tvKI1zCpn6o+IcLTsNlag3zN/dNQFX6Ox0Osvtlp1
k21jpvNeHNB1HOQ486NYv0S8vTWfSTgCLC5N0ekvJY21R0bZ4ZYsndEo8uf8icbwXb9FWG8sOSzV
tL7J8wMkD4tJWNfv/Jkuz0fSYqETUSj8zpo5BijxboJls8+ZjOynnhT8jLsXJCHnBT7MTJQvd1FM
CxcJqm/L9YyS+HkmmMQg2pxvMTBrwnrApQV/6He46VoaSS2se2SGPWAnsxV2ZUdRCwjAUvQLbZY/
mo729cU3N/7a7U7s93N7j1ORQuethIj55bzHrtL2LboeC0+kRkpbbSVBU9YHHGD8SlMMMjH4H2GF
UiyeN8zg8aViUSf6hGN5mjaaHG2VnXqnx00w1l680Sl939D+5SdP5Gh6b6qrt/Ig56mIq0AcsnZS
VtM0/IroxvBj51RNqlCJGjBbZZn/Ev8atU72jlHE/nSHrOSuYImk7WbxGqkIWlS5e5/Be2mvo6pL
0C4rb721lff/rEFOgdsVEMnzajXf84nAtTuQguvAJEeZ7Rmlx6qJ+ewhTpCtL613gSGnanTgg25X
hkC0yQAQvIprBz5W6lLuPfPhecUCTTrImOlUkKtqI9Y8J7P9QlU9jIZPlDn0Yq23eVpzevk5kuCm
mI7RwxsuR+q3ybkIWTvvAKHmR+5uHAkuujp+KapdmSKT/DbXGlFD1lS8nPU8U8VYt6zGWmc2rWWW
YdIa0siqdwcPmy96Y5mQDXJvWcu00qPdJz9eM5JhZgyP/EY5uPrLL8OuLWjPuQxdWlUAssOqks18
Wlu3izCU/gVbO+zCDA4rJp72L1r73yuPHjTqfWvgWUCIZzaOviuqdhMKiK9ftFZFk7bv388nVPZY
BtzXk+XhmA7EXRBfrhTAQeONv4RhkmOWqsakNYNSQJLG6z8bMhjtgIxxBGudLsPr1wGeBGPJ6mX6
k6oLjDbxp70cCNBOViMpzdMoJG4jYVbR0SsK5aiy7Br9/PKVa8WbzwhHRUCFXiGa2MXBYQJ7oAjY
Zg0NzdiMEbQeL7ujJPtym5uD9nnvTq3m2UcmK6x1O9JqXbOx1pCWX5WlWnfGhdRFd6KWZuPqXD6u
UR6bh9aNfUtNVm6uGaHtjahhMPvgIaoqeh551pbxcp9Fzm+zpyZB0PQeus2EWcj6lVfN6Kskc6QE
RPZXmdpir7ebf5Bdt3Dm9wJDb7MABnXms/SFkVPWUQ/u/cvM3r4Ai7agI+Tfc8WI2FTUMTgmlF23
FkYRF1coxOWH27dtsT3QNFHWy8Jwrsg9/4Ha8GAN/Z1Oz8fTbiQhvBXWVZkXZjSCPKoKhrFGYT1A
wl3VxWpddqIxfKNnv5IfhUlqV9blFZyp3t5/XXHJ43KvPEhFEcq0m5D0Yk+13+szrp617tdl7F6Q
V6PkTnN0/dRaeXY54OcCZfRdJ7is+GuNGuFZGXgk/1Dl1RC+kJm2TpaqhcfmejuEm+Dy9oeobzHF
7XygXOzn5Mn87HhL/LS67SMBbD+XELhgjfyySFpz5/Ij/sO88JBjGhZCJlMRIPi3GJSCwnp/l2yX
VFxqoMWqal1ahIHfPZhtuOZEX1T91Lxs4KjIrgsJeF88kly3gTrWf1ryq1J9VXcm7qTS3g9dcUVO
w7cVqDK5hljtnl5uXYb6pNR7E2j6bSD7YN4egdCX0QV0nAVaDOp+WwT+/coRakjXSHR0HRyUxOtw
9kjiByxmGjGmX3T0GkxTwAgrwS5MU2pEaoAk41cfPJFItNPE0x6Z7ZyaDlm43An/riTbRt70pNbP
jvUTIXZrtkx5CWS71aZuQ/8fkievKJdurvnMSW0zQudfbcUbgjdKTRFF49HdX5UOwwXvpElSli33
MAEeVTFfmDpLIGGWwH8wD5zkPPKZfNZxNyE6bz7/ox2nJGJb6ky5IZ5P/UCWHTQ/LkVBSCBe5H3U
KaxB01gc+8jgdegPSC+Xynzsl/6F9vRpMEV5xnb03y2GGGtn6tGArxaFGlnj9a8Dy0oyULAdkkVc
OdlaAD8aseGxb5fcjKRbjmC+mOzSGW8LRsSmq5v+H2UXGii8Zo248vvtxo5+c1RikrwlXuAQCLxa
j8yLlw5oiLeFdSBZzr6PoiWIkNUvXn3WTp97jEar5gjOMVr66fF4VSiTYDdmM7XjwiSBkZE2oGV9
HZ1GE4csr0QTZz1up3u+Go4Ei5HXUZ5O6sf6IuMqblzJh9W1dTqitEZ1uORvZJvGWsewN2uP4Z4Y
BBqGtGbJWd39nlseNIAJLjlkd0z0i3z0iuY4dyeW/WtiZiv8R8OEGoNULIqj/h6CEjIr9xwA7yii
6F2Pkff97m/KhthhrI8Iik8UgRK791lW8cd7JG8J3YYBymSacjUa8RL4W2833ecExQI/qhllVdN+
AtGyNh/7MAZxEQGTmhiib2ZFf3B6OeaMb/MUNrIQ4v3xuZG0sjFmpY7OQ0KtuUw+JAU21r6UC9hj
gdSCG1liabdPxhCZYQSV+vYboUiAY8o7hIL395eBQBii3MJ1o0JFMC/qesIvQArwOyOnV77GIsA7
9gOeKfBRRSi5lByv/ECp6ULYlua6CLWYDl+UeyazTJd4nxdof0IK2Ci7m/vAw8HdxPbrO7ZwR0FL
RtjEgRY5EwgwfOFbHG/hl7VpSnECgpuNa0Y3MpnKJe4QTpQSiWdVm3Y9ZlW7/JATgc+u9/0OsxHf
E6V0THR6Xh0Y6EkPmYgx11EhYZP6dEonziks3dDhMlwttPJrMpaibCCptOYw1kh6wWq1rygySyQo
BVgm9Q+k0B7xwkO0KSzwBYcBTZqKm5azl8uqTWj01ZDDtvK4uCAiC3f4BSQ83ksl82WNzP8GpuSd
70GWlDNBYRskAt3Ygr7ZKik+mK6CbCKbRK4HXIkudWxhj4PWCY3x764nPyAFYDBw/wzW8UH6+ijt
usIoTWmBqGQ6jX6qbAcHzbx3yocZVHtVnL+X6otz9mT7EkJsy/JdcXrChBjj5ulbkU1RlcRTJPG0
BiEXA+SnX+KgCyDY3xVFmYAhPnJAcrN2fq/iPW7POKN4rTRaBQs1xKKOaFtOGEZZbS6rr09v+NH6
6WbCOIbmQ5a28E2WuWyLODnGriIRZwTu4kQ0vC5sEzDLJnFTfScsouPNGi68S5DlrGBQfWzStn/o
wqcbZ2FM9O0Lw5mYnWVaHnelgxtbSkL1E3BSYBwJOHabIyravnBovvICRojHGjp/6Y0ZlhulW2HL
7WIjlgPUOmM0jQAkLt/Qw3ix6tB8mvwVdUblhCdYGIOan8Son4OHUBHV5/iGlzm+EQ6vn6W9t3kq
NWPnPL4iGkO6eAqn6Boeosjpv4sdlRsJxn6SJe2czhO8urDgCnecbLcmPu+LZfFjqidTUyu2Xk8h
6wo8x0GZoliLC1MolPriu4PJkv2Rp7UP/OHLB3/CtAznpxGrCAq5DpN4tL4l3HuQP0vWuqgVmgwt
1mtZEEXG+6iqAtpZE4EtYP5gmbAY1oqVboI2IlImiGNMVfoVXMir64h/9bNpoIqnnguRocj4uizm
yZWK9EmdP6ycgYpx5L3eo/800S9pbav5Of1oC+C5IOoCTsidxBJTO7tJRGy/UH9HxzW/uQxZ0sze
EATmz9xcvDOSterBGB9CsjlMp/Tj8JOZLNWXcHTig2v6t+cOvkOqQX4EhM0ruN6FwIzHPgV4H/ma
uoMExwsNDw4/GPiHKVRQcv5y20Q1CD6TwdoL6VJqWz7CJ0ojAhMuT2cgOfx8KUTi1O+YBkZcMmUM
GVRPr273kt7J1sgGZy7rCX/YrWZgY33AsaFfrmZzt0mdTHQ82kTxOMu8btSC75me17I2Dj2lA1HO
aSCkeItYh8be/bNJCFFyR3rJnVs9/037T6h0r1JCkFUe5T1ChmuGYGUuqhOUWDrJO/AETXNpCD6N
l5R3kePfLec/3WLnqElibZZJzbjdyU7qpAuxXyIfsVvp3i5IFB5UyiQqmh5wAXPOXo8qyjjEbRo0
WcoyWCM+6RdTo1M26L44nq4ni+IXyqpv9X03zqvx4DyYA5anYYNu6+Mpcc2IYkcEKQbhC8SbV3Ym
Rbs+EJMJWgwTCBX6uZHqeogXkJTrLjM7Kn80v0e4TEV7879EdyuqpHxcjSzftbbJvsQ+0rn4BmVH
OZUcNbDonqMTv/lEj9nR+dXANTPzCOTHkQuHTIIDpbcNSf1biDq3WVnwgkPzPZfdJJUZwUUv9EuE
nHS+yENuHNlLaUPadIEH+SLTJZ+L1CG8hzLN6G1jnV5UeZRubvrKDF2hF509GaRZG1i1BVkKt6eW
PJN8o6/rZtxYRwbfGb/yb//rGF/VFO91Ilmz2e9KFR3weq93vADDioQ8YukzOnQeL24GrRjHA3Zi
AoQYTKDnh0HIq0zqroCKHxvtIENBEWxPDWgl8tcNzULRW7OVFuToRTr5WSYlEM6HAP7VTTyqRvLg
YIiy2p04eRouJl2ZtLsnnxITnV0ICpZ45ycdjOb2D09lg8eHqD8Ge0Bn9XAtQPtqpXXn/sKhnbUp
G4bUYpuy47qvA8DWJZHqq+RbsxKpkW1lDNUFP9gBdSws7QAp7zjFseZvnXMkW6W9+WWka3SZw9aG
W8T+khUJZKrJ4sC5wFjPtPNhVnZiAWkZdcG1FZ4UKasDufiLg7UpEn6HKAj112XS+eC9uug6F/7r
S4mpUCFb+6kk+MrUltxF3B15vDO2sfi+vyyUYJyHfB1a4mYO/lNUNvaaCmfGQ70Z3Ex9gy0QcziQ
YaanLDo5oMVxbecuwdY+JplnT41EISV8fnjpfkvL1BRBEwQxxeT9h/vMfT04dJWsir6mBAkrFMzm
6NdpvGCNYBTmZep9piWKyoID7qgZTdzilyLAYljz210u713g+b2K8mE8REZ8Qjxdj4RYQR3IDjFd
3lPXgWoSPaExv43ek70rSm0gf1qUIikas9bFNbc5ssWyvUuqJNas1h2gKCcYPl/CbfyF81pwqjob
ew1dCjSAIP6hd+OXfHEU8SBKDkKg9Tm2FE56GUleuPaeucONZHLhVF0YRmtMsRYbywjcx4b8i2me
DfVDR6Ohd3BORnGyfuikVmgeXj/tQeqjl8KIQqrRrPSv3cF4ZFAzw6PrD7Cdx3Rx+FpkX2E2Dl1l
aJnt+DBCgO+d0qua4AdEQOMsttL5V14iFFhX1yqmcqMAjXMzuNiacUh3VM0J+v/J7xeBwAs0qaSF
znQPKniGR6H2KXQmxvUUvmC89dXpaPV07mom8n6FYX1e9t5/itsbyu2lBFdThIK7DstC8uOIBowl
EEsoTNhzJBYKQ8ErjEJaoiBoNscexMvRN6EQ6y76smzYudhN8HqdcmlisXcVOUbqmzq7ocxIRIC5
MdEBivkcXNUCo2xt/iLMqOUxnCVJz7Vm36GbI2QClYxjLTOVB1p1flFm/R1rr9kPnesGC/08zPJA
dz65m8+bDkMUXEQIqAO6KmXbugxYjTa9m0k6QUbFiNGKqzltrCcDtZpBCtg590yRmvhVQYVOF+V6
L13NkVeYUVyPQwg1nJtYLlNMd+hTZNbpZYjCWd/H73sgywdKEt1l/FyT0NehnUFxVvqLew0UfXA9
lWGh+wVHQztbMnY9Y4N544eVnRJcDQ7mTb63UkRlvYF5stsez/8EkWntHfrolguAebzSee277H9+
egGOgBVJ4wu+/+GJfNEVcHlW0Bgbcj2niSpzqaG+pIJ21de8XKiRIVf9ZGl5lVH+HWjm/DpZ9vw9
4oxxfJbRjPo1JIbiZHi6fa6tcI0mz5URdRNyzH4McdbBSqoerAlN93JhV8lwQzht3llk3UvxY07I
sl4jaIz6Tt+cVhU7/Uza1o0mMXWSpn5KVfqXptfcKLN6Ei1LMGtXRRp4CnTZNorr7bpIJpm61ncl
j5s4Q62QaZT5xlCxgbwqg1Jqxxt/cEdizzA4IfzkjrU99Iu0gHeuaGsaACXLTWlavNydSV0AVvuN
qRdKLXPaD8cjqLbEFwxvUek4qfDnmk0Tq4jUP2ZMxig42OwQQQdzR6kw3FP7pPfNhgXyKNERyBjN
QDOURONNrHyX7ENmm4p8CVDbRBo4DIqsO0XIy88S9l60+zhkGKFAalLtxKPrIvxXiFwIOTdVNPcx
xQDPzduedXiH7EAzpiGfGBz+JVeRQouQS1JT4o05reKj93JN+RSUn0Q2G2OquYyfdleCssxUuR1U
F3EGea1G7kCEC1776ryTtf3MTFG89XNXxWHH3iKOGPSu7LA6SrvEwh1wBEuZqM1/GuRWjdUyGoqp
wu2TSN2Ye0VaGQkNfPere5XRiPHAtwoC+5JTGfdhAWPPb/zROK3bkZNph66VQGwRNBUtppK/6Nnb
wFWf6d6n9+g2UavjbfmL2P3P23mI0hX3Y057/ztUu1UUsoeStb+vlyPhOyFA4QaVzx6TNm1fuEDc
Do9MHZJ4vUkCsOy3z23nWaROnp7P6Bo+SOhUu75elUvwNSRA4xzNyDilYJ2kBWgsU2fKlYqEPfN0
5pynhpduj6c2294QLu7ecm6r/4dW/RRZphRhLadBmbNty8ZMhJGzUgEu+ki8oI6zbL5eJ94iAW6o
6JHNqBIkP/1SlDAwMrzWoi/dRyGm397df92EyMr+xnV6fWVNR6F9vDv/OK/9u+EZcDv0r+ZZwK5m
E3fW/84RDWVjKZ2Ogsqzfc1dQuZK9losRN4mFIU4xIwDIr121H9Sb92lHiC2uAWUrpwM7NQDA2ws
Gn3io7aqlc5G0WFx0XC87ozQS8q2qzZwX+mXloeuBLYnE55W1n4IqQ8x8So6b518myyLjZv1+i2Q
pBVq0HMj8stQ5ttRYldo5zZwv2LK9ZFo0xlvIEeVeyhGa2HMdB7tOyEayfiDdd/FG6vIzgjAa8ig
DsCUU6zI3GFsrGuPBKIzDGVG/B07vIf88IiNAEq4qlDQ66BA00kz/aRsNd64IWgPZLX4D+DZrFdO
OHL0Lk4sssdx5txjqWQrupBGSAraDsksTS9CuNLLNqwQFN6Z3P1RJS4fYlFgPK5Dn7EUMyoa2Bif
MPlrmsUO5R4DQ6XehH41ODDkmuDlSkpdai4SGXpnlE1xd0EGsqiKVjFgfCCmBa1w8ejHiyfNPYz7
bM+QQ0HGE3CPZLY3oseXGBL2WLHJYypic7NPWfj6orMwtI2MBnPKuJSrY13W3Y7EGTsXXbbwJsK+
kXLt68AURUjph/6unejqr8HxHPhmM97RxCGX4zkzP7g/Dpj6zMkhbzMcdq3jk5vehr431JN/5By2
z38M6GWDbL0/BchjdLkn/I8ZsU9vJ3bxxMNxJDSJQDnfEiOQhD83R7z2ZEKu46+DfT7vuBATG9DK
UOBD48Ke8/rweuBG3b7npf+najv+aA7VuE6DTyKGyixALas1JGaZxCEb+kBNYnC8wzHNj9Q0VoXG
7n38bvfI97d2e1G8vd0U/Y2ZWWDKwe8/2evJ3AhJEcyXsiiebgqmx+frDgEBSVCAMcyqnYOEu/QM
Lczgl5bXzNWB79T5ullWZZe4ZDgVfrwEmumHdrpCYivQqw0qpdvp0HmcaalB9OZJ/JVrQKuq+Z51
iyK61/RB+4Y3S6itXuxSGmSAIxWk27dJYa73NyPVgtQzSa7nXYA/GAS4AUADdK1mP0O1/8c7k+dS
yEA82Yf5idENkqB5hKg1hAS2R+Kxn+e405vmw1D7vQA5w5Im3NVmK/ymkivFXO6G3z5/634kW2oh
B9W6ejYHsCkvMYQEwWZfgHKzcLGfpER/PwxDvjpuNiZnTa3D+71Ip22X+Ns/6vDGSNcpHD8jCBN0
ScowwvVvnX8ENedUiWbWfN6NmgebQKLuVGoPOz/wIIKaSVGnVcWikZ7ZOHgsMRTLv7+jzzbwPsbv
B/JNvZxPtZnST4tmAP03FycqQIe/Ph96aAm5JFyVqN+0Tk1wa7iiILxhPgmXZH5FdqogfPi+kXzJ
rm+4i+fshZYWiJkciD3VwauUviLBE/gqFwQRGju9Nm8lwIX4dgHOUH0ll/uV1+dGOsBnJr3vdyun
/Ab6tqIjzHcK26EzlRK9ecqB6T7c6LkWuN6hLPOMHu7k82zoDODpDZ+T9jibe/CNi4JS5POHF7NI
ArnTtO6y6/N87Qt2S8eGS8hn/Y3/8yT4DrLpIsXbFvzyfrAYB2YtP8UGPHALj2ppegthVh1dvrfl
UVf9gcS3Mw/6A+kG+ojPFEwDn6+KZmeY5mMBPH/wtvvE9fKwgspwOI+/5De5+Zo6JqyHWoCCL7IG
8YhRiuA6NyixPXtx0CvrM+vGYZ4kNTHovUydssoEFUaGwew44+D6Jf5BZBY9SfzxVXGVcA+fUJTF
BJc8g51nOeLO+XUs0n6FgSYkln+t62kCGm2po4HNS9ORFFKngSCJ3s/KNqzwj0bMCpvMATLlkBr/
onhRF3MWfEUmK5R62QkGkBo9WWUd3XTfG7jpSE6nlXTFqYLPXgpaGxdSGgv0IvZv156XVHnL80fe
D2HRYiwBRTGIfW4bIN9XbzzpgcSOf/fsrCKdjwHIIR6euuSYSDkJoIzxDVC+Yy3BDDk+J4K2if6c
F16RtUunezcCyybbzRBoYla/l0nTyTQneTez7+uGfnjke7JEfeavy9SBayKaOKd+d8J0eyUrU4+1
PnIJKOamaBD1VVSGyAJ/VJT4P2Pt26HTi6/hCHXwWjTp/zuwH5ZP8rzmohE2HHLPD8PBsD5Tvx9f
BSdUzYunO8pi8vgam5zsLRqaQ3pIHE1Bg9Sojd0ln3z7dss3+6xxvDaXKsOQFG16PcGJvlxYcPvD
v2NJOdv6LP6Q/nmWNHB1gG1Ep1HfQhtEfFbMmUs9FIeUlzMNnzV+rmLdTHZZbogSq08fUeNUTno+
1SL/zno7EIi8TN8QeK0I+fMlIAW2Zxl5zS2uHg4uX3DUSOHxBlh9pZlsKbHgyuCuFv+g/G6uGnoK
pMj6WHikaj5yRzHApWXpo3tcXxe0hqjZMev8/iI8pD+gAXazI51FAkELih61MD+N0OiOtOk8UaKD
4/h44XFJvCDubzgF5XJy6AWhJTlaZSzDixyOlBlgOnwP6ej1StCpunL9ROmOVb++ToaPVG9anOOw
5/UOR5CQTBFbXnMkHbrc45qAP84dpydV9d3cxXTRUDma9GgkguVwujW6fcCEe10MM354VzAsTCHu
Tb6YPF02i8Xy3EuK6DNTFm5NFAE8YrM3buFloyZyhQcEWdwT/3QgdwWwfzd5VfzNw8HMNiseYR0M
NDiDDkG1b2VO84U+NjUkqupoLCHYF2ZXpwVgGCx0he2Mjyj9xbViVUV8yRxqCDAuN2bindt+Cvoi
Apz957Bosmq96sbPU/uj3ACK4pORJfcyxCAgebnV0hoAQ0JT+OQyfuymZb6QfY496acw77dheECK
25siJHbMJX2R45GGi9tHD0g/RwkDcbB4O+2e6/yrNWer1AlzKkvm2NxWRiGHFMP1kDsPcvh6hGbK
jm2/pA0D+OGRT50iEOTM1P0PxCnGmEZUQFiPhc2KqKPdV2LluAgrGdP2YetZbSsqrrmKc8/4HeDT
YNbjQ9DW5MIw7mg+JN7Ms2nwmLzM+4M6xKPH6TmQTJgtdCy54cUZZTlFS8mM+vPHeYsUG+rh+nnu
WblI5fZzFk/n4mGVHPW5ozX7c/eMeAng/Wjq+YAy0iMc7yaKlzPjY41ESUQsoFPawpOj5Ek10ceb
NI8am0UkWl8XQ/fjVyGsSu8U9h62HlKPspwELJZMDWaa8bz6pyuxv3om9hO2VnzaQugLmMBMqSpT
gyTCDDGcUnQRC4ZLqc1dBKucbP5nFjt7neT3jMSTgKOA/zEj1cAFWYPUBG9sfyKz5p4UHEkGHnNg
SUCf6b0SqGnb19FG4hoZAkHvEIXmNKsAYtZKZHspGGJoqvq13fi3X5ce2Guow1HoG3YZdjao2dpa
QdgAmd2+xcH/7xAH+w9Zh9CchvvfpxYWsbgqdgfUIX14qfDs/AeIQh3KJK+DVb/HQ8EPRSNOAfWJ
iSt7mHZf/S1zUIhlcU2Jh8Mf44lGF8tCKAGGNFXIlTJ/aYGsn5STdBvJhOmjiT026HbDNo0SuPKB
L0tKiDGUBgY7xVZZ9roOsfAPwFMcHQFMZjyNodbHMABdVYHNoq0OEQgNuR54RKQGbsLlBpcTXWAv
v/MCJ3taN+ya7pf8AarftQdY0QSkORJd3HDq9cSKZI3NlTHpTJFlExmdPJFIvRIVusuYd/OdvON5
r9o35HZ73rEHnzNJMrYe4EZA/HeuFdpFNPyTlyHGBv/BYopmxmzrtR/AIbJ9pGTBcVx05IwWSBO4
KlZ1aSnuXDJMeA/+Rj5XvpQh9kq3YglHF5Icemil3BznbEeCyrSpey3TKJHimqM/uv4X5lRYFSJW
Iu2SNlXokXwg2ZrtR8UUgEfQhYMg72SoUaUwwRlB7qJNq5jKwVeSci7/pbTZMq7yISg12mQiyQVu
d2iDFgQNQ9jG7jdQgfCl9OjQEWhXoT8JNJ1S08vFcmgO277/BEA5xwELuOjr5rzR26vLP2zGkPVu
bJpz5x8lYbagMvwbngGrXPQyjY9uRt+bsJXIqgNN//TfVHn7YdiAEuD/EZKNmaXj3i61cuJ4bDoe
tv+OY9a0Xff78nUZGGXiNm9KzLScdkjsIsSFyjGZGOFLQOdu5wfpW7ufHLjsMvQkT8G3h7B49044
1di9kStrle+UGQw+8zm3Q/v20DFUkBVMVfNj4fiwPNMWNdnMMlzlirk6nHnKBg/jgbAR9/dJFSz7
kuybssbhqVH4aJBd28VkFT43OQ8sMg4CeXqhhgyDtAToM0O062iX5wJ8TGcdd0SRO2q8A31trCVJ
U1nC/XyHmawvDM/k9UKvgwV2SPi//pyINXY5Q5TUyv9sqtVirV5CpXH994mFc3dqWlxe4fyK0KlJ
NHqVgluGiNcDF9LkJ6h8W+tdzsKLVvTokgy2pv/gQtCaxF+I+0Uv8MGyAWSnFFj7/kDp57P1mnAh
tQsfxcgxnyEchVCHLbeiU7wf1N5YLcz6kTg9BVTR4Kl995PVmH1MdrOKRLmWQaBRAdfLR1+G+hW1
AUWOgTAMoeGb3XY2RDJy+EUyfdZVi6twBthIDawFLyogQoIyEmmbEkF0qmfr5Pf8O3Vf6cOhPE62
lxwrZgqbPfxZE0hkTwJaTSPUE1Wp6hqKg/XrXXdnRhRvg3ccjoqwPEumdhBxsdM+0+Elpic+EeW4
NPvyqiMcIfa5ayVaNygyDMoo3zTCZF4UHQtdr8x2QyElSfFe+vM+QVRnZxYMWJuvL5VDr6tvZshY
5sJ63NXCni1/NCQ4+7rcwktQdF6BRRTZeQjqQHR2ab4RWc1RNQUbItgG+b+IvI3NOwYfxH8aFOno
LOMjJNDFIse0eDdUHhVYIK4wzKwu8xgDliC27SxjzkWwhvsBiSwPbvIKm2/mI+iK9rgHsgH2DEs+
DNAbh28q+p+jeNt++3EOwfz3tOIRSfoUGiOPidz7BGUf0Aw3jg1d2k1F8VxtY2Ns897C8v1gMOae
w1kZKHV+GXQo67q0trOU1usUMgogb+90SFo/9yj+NfbzdaMCBYSLPnBZ/22GEmrt3/SO8GelaMBZ
GDPrvPkBMIklhHTqxDRmaWsOgQzGvxwR7XH5wdHVopLrLB9KosIekzakqnJTm9iOgxp64xc75yzm
wDWWkToMOwa5jgl8fFtRPsYh6sIvTGN2qYbzDPpQnBhLXMBOejegysebuYvJbnzVtvaQhLl73JE8
ROv2LridLmOqDtVMtafqWZfYAFrpnEF2wOoWe1XqzwSxAz3qNGGTKkFA4PmcUQ32tSqgz9cOZPAD
inmK1Ii7ib4Ik4ITNN/4NOqG+I26bv5Iy3YSg0/t68qAsbqmXESB1hyqRr3NGygIY9mDlyAu58dw
AjuPsv5bcgNsL71VmosXPqkgGQgfRIf0J/k8e78rGJBnwO0zmlS2ndwldVJIo6KFx0/9NeyBLFX3
IUZz7H/Rq3XNObZBaggYLVT8hBZ9a9zZ28CtLGgerooZl8aEiOkPr/QELDZP8tPAuX4NMgAcwAq+
cKytrXHfL7dO45g5rkbPDgowp+jvlSPr5eRDDplCKaYOt9FHyw5mQJRMPvvUrlXAjGyyDeXc+5Zp
GcJgeYSojNMVVaVk0KXhJsQz0XgTPS1w+cX6yNO3BP/O630z06nbm6TnFtJczc1icm0nZ9C0yBDM
OplZHwXMoq55Q0XUHrSQ7Gyk+qdwEyVLnV4IoPP9j9snBRMvmYrAYqxESF9ltKinsAe71tGcAxeY
FlGl7heWsy7V/pyNvxuGSkyq4B18aXvx55fKfoyAdekGHHMUEN32JSJscZFdjDl01W+EswBYydjf
EzrzoH6q1NGejUGZG8eolKDJhSVQU2NEgOZGZEsVxlVNU1PttBo/pehtriy++NsFvN+i6SOn7t5R
VeaITOwS6JP6sSylQQ5Jf+/Mu8qaoj/tYIDxIK1TYki72W3kasgS3JPNRR4R2IcsXJgu5gzP171g
fm1TFtUE+G4QUUFnQBRbnY1airl1Y3EmRLc0WFVS8cRjZgrGiNGtGgzEgSp6LmkXhqqcCo7E8mhT
xo0BfdBcf6jcequuy/ipCECUYE73UpCDY8F4n4nkTWlKIdLdB1WKiJeudQ2pWOM8NLQ19LKVaYRi
UOvWxdol/BS9vwaPu0+DWcHSKsj+ielUGf8nWSMR/DM/XLwQEF7e/HUNjCorZntiTIYxW/Y0AIAh
Yw/jCzfwKXWcAG6/OI6b50D1lJ0KsWHc2BIvp9TSr6+01RvR8GDEuddRjFAYPQZ7b1QSlVi9cl2V
98eblgmAHO+c71hkj20OsPl+s1MKVhyKefC97RBqsmB/f+Al5QinDYmuvPlHBSMJdTTQ3T0Q08bR
nFKmj94wE2x88vrmo+ZMc+9rUxcT3c1DxiTPC6HJIhdpCt/PjZAgyxHCb22W5cQmYss8QzpuZrIt
G5laVH0ZSPFmWMznphhw9fUivXvPVPOGqqsQLSBJsLHyUy1u04KhvPtq+H/o5JqdQ/vmfR4G467b
Hdc3U8j8a5k3JZnAfK2+SCYellf4vmOXNBqH61tfGqI7b2ziSJvhoTtxAHH/DSQMpV7q5EtJI3UV
yTScYuZIZo3UlnhnfxJbm5eagSg58j130ZOffbTtI8vGYwYjb1IXflgBNzkuNIPin7jI7IbbzYfW
3k+RaTIscpmpJChtIVHxBJ2mwSw3/d0E1zj7kjHcw0WFymiG5Dj/7/UwHnDFwnMM6+2wxrBewGtV
vgcp1uI9ameaikl4sWQRPvT8GHGh/DvBNr0hGKHQzSz7/fLSWxK6zqXhtyV2q/nFlrRqCVnnSKvc
B+kfIvO7lRbD1npzPGH/Bt+LbRT6z2PtfPWo+vWIIEQzE6X1ZIH0RmJ/0bp3haPCAKRTJzSqLv2g
v5nMR8+/1UdoOlC7ps+aN30mynMFH6cRj0r1r3X4+qWx+vN8R6ALTXnE4z7MsXizc1tkdXxYYPzQ
f0m39EwqVVSSZGO7u77S96ObGLWTRRrbLbG0zKFyyQEVH90guQGLVxQrFnPAvr6O9czdqfTRhsM0
rryHLwPjKllRB4l7aiT/Tw4iA91EWmPNAXDmBoPYX+6pE+Ntj//imJHd4aF0t1me4xS5iX5TTG7y
a++p4kZJ0G8cXfmO5uF4KYf3UVXAYYTQ/39YO5kpPDCYS9aWnbs8Kd+FoohFs4eJ6i8e6w1bX4vA
bxBCVBWB5CO9ZxK9gnt+RrNwNIJRJ2QxNyo0UVglQrxdmRrpiX80qEPj+CorKgexOUsOPWR4G2G2
qsbjjqqtSK/yoF8W+ZvVDb+s5dhRkseonkSgtctaC4a1X3rTahosZpBYe7c4ZpF0irFP9n90QAiS
AW+GRjKvXfoy/FWiO7PQnU20zJb4qS84Z1HjvTHg55ZWKDF4RY5Zcp06zF+5eQCtAk3DHvufvUZ0
VF1KgWVKNEMVGL1/AFWyUx/RP8uE2hHdt9wtYYchd5y6rk01FBZbmd7meb4r4c9uRizJEYDpYuhr
Rrqe4UgEnJl+9ChpmH/zY0mabCFxCLbVllWfMLOZvWO06cFOAgVrVqe1gzcVjRNonTrTEvZUaJr6
kjUab5TmyKcZK6e0DwEacUmcX38EjphmROBHAi1LrlyueqBrlmXlvzyNzP2o78vu97ssWy4nXwZe
lRAxjS0NZHhJU9Hm2PiTdm98t6kfkvZM6EygUjHbupR5MGlIv1idXbh0dbH7jxFfbZhAC9Xo/Tyy
YYA7h4MyMuzvzI5MGciCn+fC+cZ9fl1uHymf/HRGcfcIXsMZu2IAjz7xVm8wQ1ZrB4lJzCwrS7a/
8Zos1H+qqQdYPzWfFG3IkvrowIwQKH1r11Q8/jelwAQDl5TRskc0hUYLXbJW4ADhcbrsF9vAqL80
PWG9lYJjZaG4iDQLMA4KgX4x1cPA74cBXvQZw2TLXVQsB82adeLQuEEc7ruGecRAfhIyhQT3Twpk
z1Eib8jQhZIAX+71E5wgq8XGnTDJxkI/12gzeDhCLyYpl9LjYnLwX6+7ymEnQRTL84GnPmL0HzY0
QCFcxR++PTs41qOs4ZX+oy3C8lyZdIWeoQGGbiEwgVlcDxJCy67e58um09+BeKpsierEi/B/ha2G
GzxT5V10tQzZZuyYy+l47pMnk1g3cZPfjnR9M4I3iWTpMLHP9As02VzJ4qClW3ew1mp9sUpWf+Sn
oBdqDT2gqdF9xTIacs6kPGuG37T/cEKf+4q8BdUsn8nYVABOprUI5E5Ca4E2Nk62R9HEcplkTuuN
jANlb9GDvtua7zvtN77ElJg9lJXHB3mkJdwzN8gGsRAOS5WEAPgY6Y98NL0Ye5HOxOLrDnZ3qIaA
Y+EK9aEvXOluY4jweCLl/HQkULROhVdXy6xg2czs61UVww2pYLA4JQ31ChDoWiTAY9ZJMc4jIW2s
uw8Etfpy2sQYF3GnnSHn9KPwb7jMHSX3IHzPK9PgehjJU67/clt8nKXqpdUk0fhUXgFhZQeU0Td7
gTeY+5pE7MNNRhHT328vi00E23SQMvhZYZZjkhfs/0u01Kg2G2qk6loOYOLEuzoONGBSkaeT1rNz
9z+b27oIGUVjpEhh37uDyF7zAwugvrrp0dun7WKDtymb0OawmUzFJw9FqZgv09r2YwXE7hqZ0tGD
MXJQA67jtx07d4MRbEwlKc7bT43Y7c7L1O2857b1ZLw0Ye98RncqG7ct82B07DQbt8aYYYBpse/l
MrWWtXwBc4WRG/IDw2/+cHZ/cxAXmxvhp/0AJcgMpFXF1In4qILD1+LzhSSl97WCUNbjyrJZrgRT
EU/Ir7v02EGcDQwuGfiwtUHRd3HTTpcGbCO3YE0LtX+fwMbo4u8ZyHmSrPKdEJ82r2sNJo98Mrvn
Adt6hIx2MOuhYZYmxaCvbmjpRUW8gT2Z9b/aTfclIMO0jICvwLB4jukU3LkNEx3I7yyqkHXe1ubP
Ytff9UpSCxqGMsbIl1StdcwrDulf67yxyOp58X/nnW1XCe8mMJ6IpdcDOhBdogvZ9N/4azv+8uv3
tTGAiGUKS387AH6Kczfi5wJPE1KMMgnGGZ3nHIrt27YSr8IaEVVA6JTuF2zRLTEvUDwlXlfcKi1a
ohsbF5Zh9A+h50I0Z0Ufqe8jH+mIn8iLOSlIikCo6AwyNto9ZxLJGZiVFxAlKoxnsDTstXNUBw2Z
STNU/3SUxrD7hbi/IMqJuQC5YZQZaTqkR5838lOODq7H9HRZbhljzLzXl4yLpU/54MqG6COuFnGx
ngM4crwI7FWg82TaDPkxnbqr4gzerhUJSQEjcthn8gK/UeBk7c4HJLIZ0hkenXO9gOzPgzHUJhXS
scvnID1zscPV/ToGsLAP8McPUw1pUvCNEwyPx6vucbw8eCupEqbEnlgl5tEbRwLAl+cf4QA9xsOV
h19HAnVZliFsUwKb7pK94sU4mydi20/60wFJqiiDh4y357a8HrLw1seINtbCO2AYCn6nOjg5d45K
kXL4DYDeqmdhNJRW9VG/c/GpGqUgRORDchW9/XgwBOs+cpjtvegE9RV1QtVkS47ARgwMv31bBITb
UKTG76QMJkWpEJ8w0LehpxF+9FyHReGodS2VCcTjUGL3ylAtxeCbp2/WzujmrMsI58hW16xh8QpZ
ZBjG/0ZWVHboRS0GyGNzRH2m1RS4DGS7hURPNT8Kt4lJWVtAHcm+4shrOEr9up1tN19tQoGXauAG
cvEzdM8sc+CLgvbQpOI9XuVh4DHzLj/pLGdR/l2kG5nfaiMBIb6l0c9lFOABg9GLoYruw2g6rpOL
XIZyhSa4ckuwA/EAbguyvqywpqc80rQei0ynHU20+vLAsK52RzdMCakngpoXK/OcSTZSNx1IGak9
xu8V+9jTxb4a3cn6nidrW+NS14+bf9wLHlbko/d4N8VWbFkLxT2Ao8ciLyhEbDY2yhbwLybrKIeW
X9CLZ6y06wvdez6KynxuRT1T6P/LGDC4TOEeMgM5qyumWyr/NF2GCgkVNKk6+DTr9Vitw/TxBFjM
kVfPFMomRrei1I1PBoFix2RdTx7zPhXWokaGxzKpjwIT+mS69WwjAlh8+rYIWHzNDKz9XYpKjI7l
zVhtBbpT7CYMQvnR4eCS8sQdKpjzpc0G/N2Ioh61toqUJloVj+hV4B1s4XryXFKa8aY4dUfhbje2
ASjCIDdTXRqwBiV8hpseb4a0E8LqQg0gN2N7NTGmmCvgua6Dm6xowLrTTK2aLZ36/t83J+IU90G5
dWQrHVo7cV/oQls4cdfMjQjmJwHU8Aof6Jg6yZO6fHKNUar8RvolLCExv9TfgCU3E2X7MyU9DFu4
ZsJL0DR3FwwSF5USCwLPr4SouMKJni67g25DJNvWIZH3KhgiNc8bOiC1lvg/HnRUZyX4n5NYlUEq
yKv8bMNnve5ARdnmZZwqZpgT01Jd2m2KAjughtGEsv4Hxk7T1qpDDle603tLRHePC90fs9sh7sq8
6m1Hq9VTajoFiBdnNtlinM/ztYJRN65oi0p9uqjJAeVV41yGcWn4kcjBoHtAW2V3K2KvBHBXf/Tb
GWYRiZ9/uiU+cicCPxh+m2XEmeQwT91TGjE7iWfSYhRI3cL8k7adlq165ReWjlG0L/rKSE0bqHUz
SWomNtEXDWAgleNcEVT9ROT9YRVW1Vl0YPhfK+DUIowNqIwuN+mea9xqGp2X+9nF/mdwq83mSJ9e
Q/SIBaOXZIR3ZQN7xOf5gO72wOtlhXAgXVBqvctFpm/6a4h4+kE90miInkVuo/2ZmGWvvaQ4bF/y
Ci3SW7PrFLWuFv3i46GwVilIMCixKCecUYfP63IZ8ZttWa5lUlp39EiiZ3U/U0pycWmUyAs/6cjo
spS5GmYGzsFnprnvY5bCum9lD7MpAc4cm3t12NfQskPQ9U73UPmTI9wXrUXW9AGrZRO/rB6s4g7r
fdWJB+pYYfdE8deA2uSJPGqyb0LIYVfz9rHNKp9Z72nJ6220xU3l+2gdCZIIqaqUq1SoM3pebuI6
NxsZTYFraiyrEbxVIEAIzy5aSZs2vVXMPDWG3mFzdUJUTfxwBTLE9FgI0Dmk3y6Zofez0JwMSwQS
EB86IlHF8VkyNXX67Yg73BfMqOXDrORNpwH26q+GzsFhEq/dRKk1l6syaF3RNUv5lW2019Unx+ed
jPPvlFZgA0rhi0ALY3UnWAeOh+L2FqH6mf4ro9Ej3Y3GWb2aSDZyC4KSY0SIz/iDK8noB0DvUwJD
U/izJVjWd7zht9O3bo1AHF6Mer7XBxvk7L1RfIt0zeMEsd08IklfVw1NpD+EsWpGSQ7sZMIncoJV
WhsWdVLLmhS0NCoJgbrwCiQnzwoaeQYh5FjfUnj4yunszl+zfV5Tfysgzl5KKEPbbHT1bKInBcK7
mpgACI8DelCNyWg1KEsYyI0nWhCLD9BmIwcOKPHpinz1GuAVmcQXec8gy3FSiiUBPK3sVAVxWqll
JcqiIQcp1u0dwc+sNCAzLyk6x0m88amDAaRfJ0xzmhHTY3kw/nU8rFnksVHP32G24fRC0qFKnRn2
cVsaSGHhUJyvCAZIgsShZP3gBy/pkvySRn+OAOgzzxCXf9urVwr9geU0A6mlH7RrOsLBgBVDjwVS
t8bSNK0TDn3gOTSl1e/tKcZp5OuujzYvjDIkocJnUV5YrkclFYpeSVGPalxhHUotekbdHSwM8McT
H+vlL83Qi//ei7MK5LAc1IU5L72DkpxL32Mzf9onhiISzpu+/2MZqmZGh9gjI/MRuedB6JvdZ20S
M1QCFfJP5N8slpPsyiIx7zWaGOm6OMvQuJUIHz9N0c2MvEpKb4Eg1i2IReOQZ6mv5CH+3MKJnUtA
Qsb0hOzKkSJmQeS4PAy0jSLdl0b6Zs0BP7HoxKK/CikHEeBHqbIcRQEQH0fXGsWnYffxOINv6XpD
1zNSL4L+ukTJsth2yxhDjHs+zwAuxDx992iXCiq25DSgflYm7S3L1TQI0rHHjx6NzU0qdRz/3Ipp
GEaijiJOJMjfr4fug6MazKKLj1IJ9c4hzwWG2Q/rtEFMENHK5wZWzI4KJEAzvuJV5F4wC5SvU1uo
bdO8PhstHtyvi1anFhhngyv7We3HwdF+5gfMIuXL7ekFHCnQZ2+L/Xm9+o7ftGwTn/gHmNL9ZglF
jHszMl4P2psCrTHFFX247T7vZYkgxAlqaupVy11tyNRuRwNZboFekuSz9lqTdD9Mrjn6Q8NxFLFj
oh8YRz/+PqOnhNjUhmODsH3ljvyraykKp4SL2QngDzuRhpNM4urCADqHHWYikyOnGB045zYSCvo6
YNmAO3DSKU1i0dH/9a31oNjwgLfL1tEvDSeH6sa8MvwSCIl/JELhDjtMpttTYz5yOn5pI8NrhNlf
nhOCnLmqXrEydemBD2EA3mwb6/DTfdRjdyXEaeczUDzdSjmjgyML1wW6FFl8/E0a+7GPjxmEP74S
UdK3Zr7l1fa4UHgQFkEjayd7RdAG1WkdDjzit4bI+tDG+Hl+fDB1iEDn/QtSFg+d2qfLwFGpt7Qh
XwfdNfwv7+RTHnE0m1p6sjJoBawQTDzSqnrCvE++kUkLUquIBB2aqyYs6OHitGcL3KYGiZzAZvSY
ruo5z6rkfJ0xluWpVBM0Z+9C5NSCzs5bnngRo/bx0wagXMLC7gDOjrP6TzHSxN3N6NJLH8y+RU4v
mLlOELo69fFyuu/yMcp1BKGdmITgfMby1h21kqN0ORrO707hJJZ6OuYNH9bqxEtmyvOsSNcw5hn9
R0G4zTVn54mR0Qnq0cJ6Z5Najs5W08jHC806EfyqVxx8SRjmPtDtUH2TD+QWPC6h5016Cz6D3PSu
3hC8RyBEOLO8yDonNOEw1BSoQzur58taRDTBlBCDtqq06n0bjyQhJ22j8esycFcDNDgobwxOyH37
I2AxjEEHQaQSf4O3gyvwc9Q7P7dFcrraMpgD+ZWwaXks5xZ+KdiVBMVa1xfAr1oVpinP6vMJpmpC
VbF4rjk+sltmu35zNvpJIHMjFWjUM7/nXbXe2a+2LESEm0tlSd4zxHRnBfFqAl662kesw6KE+o10
kzls9hK8tEO6ZuhqgN0oWoe1lZKLPyQWCmvKyemAywmJRgYqtj1lnoKiPo4kDOHeBni2bRILTfoX
6f+SO9NBgpmHAfCCWd7I6lBG9yBdlJmD3BKhJdQ19U7KGuEKGR0bgtuTfzY6EpfZctZjVmljLtlW
Y1FORbYm/RC+4xc9C3bLO/ICQFsQGQ4lmj9O9Xs5VpGTpaZ9yrMRPNgTaujQCtgFPoWZ/kKjY0Cd
HJNFNJjW73SxOO/S81aombGYUOWLcW292D7K7L9YWECh79oCEtcGzFEe/nNhOJurpplTLSVS8tgF
qWdLP35aU12nyfUi736lm7hlOJdmVROO7qWMsBkFmuTaA0jAzVN98NjhgpCerBN5MKDM5OQihTsR
YcTi5FHaixxwAcmiznEsnl1kDe1Y9LMr8uMgJOgqD9T3vrYrUogGaKYtthDTfo4SQf/Y6kpinWyb
R+P7biqIJ4/2SzW8pEhpEl1iUG73BwBRPYdF38SE6EZoQRrOeupMOhbXouowXfT56uGLxu2JJizq
yyVvJCgCgDU5mGJbsksGAQfkPmvosWaMz4byqWJuBN2+lz7Ymi/Tmaredhvz0RrACCKmwUNgRCUe
x48S/VvLeLM8dAqQhzTcbIdkqOIRj1aJ2RTwFIk3LjBBwAMzNKEZ8vFeb3bU8ekfYObwag/t2fSS
RbJkNcootQtBWAGVi+BtG4hiHsbQkl5Dou7N95stnnSVylsBDWeFZwaDD1uk9U8KitDerg6RSTmx
cZHsmWvpxDDr4sgZeLyXCXF6VNn1D9ALsyVdGz/YYN+NwJwKGUbWkvH1/Vsle9y9P3xQTavj1EkW
+iqQ1oUiVThkMYVbPrdRX+x4XPAjufdE4uWFRAghagNx9tLbUbADL9tKc3vVB0vx80+YMKX3Ex3G
hPoFq9qsSBR9f7F0TVFFGgIypP8VOqxPeGZlHeRzJKGuIHqdh2rayyhLT9UCf3Me6H+Kx/hRZ+d/
dERYXAX+NZAaixkKvjlZUizGnJar5f+Bz6Lj6ouFN+UvOcTZLT/kV6EV6SxequgYNZ3xTexlDJG4
uUtbMDKmULdnUbDBYexJNFpaHheD3IKebnu36EhFiSXfFDBt3T2hRwV5ekEzw9AK9Qseed74Sf2A
ANuDvnVZr/FLgIjcUtuTtjWitktPIELlOOOIRWxxQHzBSZtv0h3xXuY60mnunh5zIH4hAO1M/35G
2mLXTFj/tCi88GuCtAjnhRbsnYpJ1ahcRQ+nkBTuBVLv3E+Catpl3GSWmdFuvdJ2o0IB7TEAyQEU
wP6tJIgy7bGqrzpZWjhB88Y5prAZIZ9t/otnPVcHuM9pFLy+o29kL7BJtnRb2N9X4A4+uJp4JewM
436VHOvPuJW6NKJBBla+d6zmbY/h3uLPJmktHiY4xkyPwV2Zk0seu758REKSqsEhknw0Lii/AonH
CTDZGnRv1f8ih6bQ0v6TaNGr7t87Tm5/+txivM8QmVO6PAr+YPubcBc4Rdb2Iwbdx1H+nwFY2PrC
O7rt2aTCPSNOKQhvcU+sjlfqhEJ9e8V3HSgcxdzuZ6MojQzTJu9Efcxt/akyPac1P8Tis2lff6xy
PiKu1vqPEZqSQoVcahrS9z+cbaCSC5V/2u19BhB5RI/eonv0HnqRDxsPOowR452ZQmBxXnsNkfIj
k6Ujy2YHZSEbYykCER6qXU5APLj39LzXW5dowWaH77lSemnWr+JyOvsypEeLdBvbh/BFkg20i2Ti
abcIbGTxfGKbiJO5zp8lmpFsNXbCAb4kLhqIisP23zOZY8fA39DXfBJuiiecTonKBxs/LKsZca6L
zBxv8wz7CcqCczQd/nZ/qqz3yCcXttk1i58HS8vG/IP7+dxaxxv/L0xP4/VSlRmVIhk+K7Sy8+9+
qxRXtQBRN+pUOPuMXipApH+HKJxQPzPfTv4WbQZBknBPalSizqWYfhTYQYaqtcM8L3Br5dzp/Hvf
Jq/DK6qEDevO4Lm39wFvUTPddTd8FqCt4hIz/g0Zgu/N3IFjpxejOeIhpC2TOaJmL5tA6dfGIWR3
DbPJzjmURCtozjpYcOQB4VNtKpdFc3AkZLfTaC5W2Xp66NUedpW7rsPtSGrrVBJKyaX+lxEjLqv9
toh81cWat7rlaHW+9GwKKc1/NVeBzLAIbDRqXCW/1xK4ArlOJusx2TBraQgEJ+8QTSWZNPCzoi56
33uvNGmbYClRfAdNCmfss63vMC4K4l50W13dhl54yS2S+MIxIJiHfuF3JEj/IpVAIYc3ivfdUQNN
CVFs0BpoTK8rNdHNRd4+Haowp5XqbHbMuMgj1p43a6HD4cPEIqyDWbAqxGafWUOSPijRFQSYxPV5
qzPXR0UmdXGAAdQlstd6HjLMnPvTiz9Qh2rmjclcnnl85Z+JQKEtfD8PpcnRuTHnlzp/DtJqpkHU
DTEuHJL0+d+6LtiOcVNWHrMLUMqRkeBG81LYCZ6Tw8tHd/D2uwd0Syxyz3cbb/lq/6ml3cbkBdvJ
8IK19cP8wDCID+mOF1tEvjnXzeXXs1ZXckVlnOy2j+oB8GspEa+s0y9GmUxl2pdiSulLv0YSPQwa
2EG1vn6c4jzAFzpHVK5PbxUjl7Omu3Hon3bFKmVimJpSy9BFI/laYTMGGjokYwVvdtt9+Co5WLl5
fH+VF57elc4WYVGhkZD0F65OgEPMSknm5BRcBRsFtIpnspSJXAxWPVO+RWji1JkEVHKgSoYO27Ro
YY7EUV7WQKNBnKbLw6KJj8D2jKoObIYQQAxxgRK50xhijJ4xmUYA+/V1tdiigHkLONuF5MXyUJRf
KdScynfoXOm9SojzGzW2wk2oufbLSkII4VQg9tlRjR7q7xdsrTGec1wzrj2Wsdjc0a1OrDTUOFUZ
6lZbHCSqU7qXWHQqOnulVI0j1l4UHQxfcBgF1BC7FVDMHL2E+zXztxODLtAg54BUF3txR27pZCtR
tBUs3R8QIQU3J0AvzRIQY4bw67Ft0UjFxYM3v992n0N1rDF1W9nxequYXiMuva46+CfsWtbGSZyb
WgFqk/4W+L3Nr7Rbi7qNli4lqE8sNE+zMvM0lF6HOsK9jbw0B1B+S1OVyxazGzKYivXpfsNXysm7
NvN9KVodc9DAAaqxKFucXNE78VI7DDLXZkHB8Y2kD1oGVhKcdRcceOwEbITJVmwuvuC4mu4xJkZw
8FkckmHtyUq1a6JvCeYzfwbOGZgVkMqRV8VlvAwq1dejEPCC03TP82d3n9sBxx1qbtNMrJC7ZW9r
41+UWF51RlwMjT4OU1dgYZKMHf78F1xYMVcW7pMmyj/HQTH/SUAwJbM8r6zkKSVEQNzZVSge5sUz
imC+UY8oFj/h36BnaukHuNKC0aF9GXjRqQ8qepR+QdGSNDmuDVy5AV36G2gKVfdCnHRo/AMJ6+3H
+F9FLS0vHXfOun9YRew3XQUMCutwNY7Bl1rfPG6nWUgE+MaTvkvTJpeofQ0YKdP/d7HXr4MHcUve
0UoiF9lO+zKq2OJrx7lp1qLEcXoY48LuYOj3/OV8ih7GEd3K37v7pRvy2sv5P7vmfFWnWYZJNQQk
AL6qrio5D0nvBSZh/INNquE9yKR9VFfpmh84UquOdHSJGQ2mTOJR7DJ65cArGdFr5f3/DyceKgg7
MWhSr9QoR8qpsUYUXBwb82Oqosa/YyEoYl5gKLtYn/316beQyWT+ZrDKFx0JoRWHMYxIrmmQd8Iw
cu//o0C5Ook1acwZmV4gi1B24t2qFPC1tH9cJXYbjmGF8AG8/G+cwyEsc9h5veNn5zRbGtR9OIZn
uEF9ygL7lMjfc+XfqWPGZoxw+xwCFlk3AVV1viezwGAHfc0QkYN2lpuO0KMiO/jN8TgPgbHq14ee
ojZpOhcArofg0JmK2ZuR/4Z/k992X1EewwcGR8mNcQuw6UEp0O2kz5rWUd/cB/qxRM9/mr1KQjIT
yMj/N8MWwTC8nBmdCavj2+a70zhEyKS3v+jOqXAOVoqOZ2RCzhr8j74SYLrOdELxpc3yMkqGbuKJ
63g/ppnmZh46uMnGU46gTk4nUXgw6GmuDWp+EOM1Ka7Fso6a4DHhoJWjCiPTUHh3EmwBvvsEN5HK
PHJ5kidVM9/TeCL5xxrcV6wCM2MRE5V9mzSihH9u4MANDThlydAboQZ4r+oRrb9m+3vQA9fsFXQH
CZI2fvP8wFStnRNdfBoahs96PDdbQmG5B2haHSA+dSjGPgL5aM+UEjTOiz2kET1JG+0bghW6AYmB
Ea6ki5iYlD6u2jqusSumMUps5BdkpCqJvyzIYYsHiKXqY+Eoxj3PwsKdGJTY1Bze9J1SYoZKm8R1
cw3dQOSBu+wlU3nwh4uuVce3FjJ9f5XvX/nnSXHgEYJMFtE58vBdnkfECC045k6NNBmr3Ku1gDJj
yttBH/pWwzT0LakE2GeBYR4BPl2t9xXLH6AkiT3sQ7b4jOrI/KB5HtKrRUFnrMnGmd3Mpot1d0XL
p6G+B3DNh/BVYoXq/bK9rQwk8Rht4XwxEmI1d1It8s7SM2x+KnU79CXPmxrlnkrgHppOQsJeltGT
K4GBTuairRtpiSNWLowuYWjDeTyiF3DIkeNnRLA56Wym7MVWsTL4nUB+aUz7P8aztRJRBS1WROkd
rqFoRW0GBwaK7gAr8ifoU4PImyHAzKJ9WzqSkw+E4ejorGRWDGBCB/O2pyYjyYtMXiL2RyTrHjD+
frv3IpMvMMrkjzlINiFr65vwZc+6ETjZFpYQKwWRtVZbgeOrqdLpdQLHGhXTsYAqtj3/HrFF29w1
GFyh9UsoKUIn09YvnouZ7Q0DUGgVTGA3avbOTpsKVmW+vhQnBhUssoI/+Vk1cI8pwjabCctceTB9
/4zzBzf4RhLDm1A4GM1YU3LJQYE+OFqXAvANSOzg3r/KRE4Tmdw9H8HKbvyPvnqv62/e9OWNR7rT
hQUeoK86iCBfv09/FNpurpPi5jruafwC9Mhvo0sxkcl1p8BP4YiIAdPd3k6WCF7beYi5LR099WyG
86PajvM4bGcPJnKTrXVFFV0ny+0TM0t+/Sz+MwkMmyMGoVviWgsMXPjB/asNBpdENRioD93MRXr4
COkBEdPfOUU92oj6c/uhuoLncyzi9hqrhUJ9nPSAll2J4Jsy4DZpdnqafc1NDFFpDfBWyH2sVan5
apqBBX1bI1qL0bI001/z9BuvFbe83NMRuev4KYe9UjjoSkgO3tHXJ6WmkdYToCOSwcTgiFT1M4Cx
CNO4Rb+4BAWRpMRDeE7L9rhvk6i0oGPn5RTiY19HHBTRR0BZfA6uCOACFl7Vl8KQIFWCdB9wPC8o
AM20/q2b73Ul3S9qKxbzqY1FDZ+fwq/UrHlb7Ua4eiEBg8j9G339r3QZrcP2DebRGXu5A+0WDov2
VTf17fEdlm9/aJiXzrHlcSF3iJsCuGHv2UP70fAcVobGqokbrdEla89JNJ3x9+22l9Dmi7Aji8D9
ZopgVA0lsVMh0cNM95Bvwb9+WyHO/XH4wS9hzRXKD9iAIiVPJOXxjT2ZCZURJNpR5sIWTKmXi1us
qO+350afMFJGjWG8kcRFSdh1LoaK8/A2mN7hWFRbxJbN2WqCIiqB9Sr2/6gXGuzCEovYR4oJk68U
A4MlAccXn2YF2jZEEefy3aSnGm1wgdwO6x0tN69FCOJKM1PODcpyNdFFfU5p6ArlptpvZJhRpxOX
Z7bfAJbL9rB4G1BxsQcdWfmNBXAaott9L+EG/1h19Uk6bCTjXFipTXzOi67+d5Q1FiD/gMOo5ppg
yUds6K8XRtvxBr/epW5HB1GElGa5tg+1g+NB+mEeQifrRI2Z8qps1fSFc6I8dwggz1Q5eKddOuU9
1P6S3hTvYPuiORW/jSMDuWCPHQ46XucvSBDhb0TkdoEDccVC95nktUv5Tge6IVb92zU2kPnMn6QL
Pi3FP5JynmvItcQ5Jv+Ll7IQRm8gk1R6yU/gZzzDr/dwJMlIiF+P+2Lzn6+dC4gyeoybsZHY+pIf
hf7DQCqCqVUtY/BfNIAgAXB0rQdZ4mGSo2lB+OrWsHcoUW2MRXnt76ZRzHojCI0YWnLO9W6kOv8E
+84OYnh8JP78FKAvvBQo/u2zxODxpE7lkKuRrvvwauGGfyHhzDkvspnG4YGbLIOjcX2cybPgEYgr
w0Idc628/NPEvwlF0/DyN3ROPxmM8HJwpp5Xi2CI3I2NYp9mu2LsJF6RMDl/5IyG9SF7MZKpwQsn
fRJcQrEmdz96dhy5xS3JcSf9wCtu3P5ehvUgxw8CxcLxhycCX7E8dHf+PMjpQsvfzttYkbzwVzBD
vgP6AwJjUpoQvw1TpLUXa4aXY3G6nfyaLRg3OgTDxZHhRh5Eux2jgiwAibADBQ4ufvSlpHUQtCWf
gSfxE4MPqP7bED3xFJ40zFTjIvhAfYu1PlKviJ3FBsNSwMj4RxNvhPm7ASVWEOPvW2JUilcEhyeN
sWesiBuB/I9yirBUswlawiaOFEffkx4B2AIvr09LjjsttoM6Lo/2V2N6ZJ/lNR9QcDO3lz5Z9Duf
fMe09PN+jj8DdwJs9Ly7a8Wp4D0LWboV1uStjOIuKdWLiWD6Jg8NZ0PuQ7YCYJAb9F8Y+OXY7Hyn
OgIs1VWGPbZBCOtGbz2jc770LbpnfStAFFSa1nTcB6fqJqIuZuY2aNCArEwStmmf1ikILdP3Gzqq
NWrl5Wlg4qRstfaETqDwnGGIADtMlX+bbXNud8tlOb+DT+x7by2X+JonOkGk8jRgbPBK0DKtPqyT
4w+hFeKeI6KdJ9cc1ahp4whNZMb3+mJb7mBW7eGrjVucouvXE25ghfuq5klcHD5ggKxDGm7VzH8Q
JI4zNM/ZJKCM28tNLcTXy9lIs3gIU2QKdSMpDxB1Ug57TWhT/aH3J8e2n3wmdi1BhaChoYvCzDgU
2aJQj/hzMoQelbzaNpL6LmoRrw6rckHwJ88SVddGi45e3NnPVOQVdZ8zi1MyYGjhQXaarK4tHQ8/
MdgS8goDeyz52MaIw9SiYMdVsCcqvT+WvfbycM1l27YFxg6zGEMmKk7nbyhZmwH1lkqFMV7QpL3+
Lcq2SrmC6G2Der/eNw9oWz+haztksZn9hBsuYcORrc6Ul+a8d9/LcBpP2yVSzI7cd0/DjOi1NZpM
vcxKqYF/dJT5s2MLuhyZdewbYtg7UOMLq4c69/UBg+FOfJCmj76OrwRlaB8XVOHMhF8UrkojKyL8
KF2YgqCzFjS+zmkSWVQUXmzkPbfkXFhUA5MR1oBEuEHof2YbacvRnpABD8zdUD0YTio3LrbQEHyc
MtCShELuoouIRPdPWkMHsA+iwpzKGRR53P2ql8vDnGlQGEiteF2x977dg18WMSgvO/cBJDc26gFA
zQe+99klmE6/NOA0wu6J2dWPFV2fiCqW3NotMyYkdBjP2oCyyzMkt6dV4PPgYdWXW4rYIORSmHFu
bBwyx0rMfCsmsPEXfCLzXBnALbJbC/Pp9AzPOgfmOi59F4IUySbUvKowUqfbEbr1avBhDQfLCfPD
N4eiaUhpi+Q/Dikl2bNjtgVEt4cnEy1B/53pUiAzBc6Ue7UId12tbiZ/1jAW/XzJw3oZuOmkqAzW
KC6OuCA7+KRxhg4tpBt9cKCnksASqzCTvS/kir69PJl7pSfnRZocXhQ0uAMegJaSahioSGNGLhoB
WsLib6H+1j8MuB5Zk94FEtLxafS+diRRv/S7vsqbWd5fxv+9wEIoD6h0QQvqseQ/i3l6I1DHKVh5
KLV5JlpS+RWp9rvkTX0PLk+xT3ehNTYPPyP4DuvK/JziV5+IUNxhqRrDYodSrEKY1sXipwEySflB
OuVnvuF8kTglG+ROfZzjRbwlJkNzjGJXyUiHmhFQnWb+q2Hb8OCcOD/9se6ujixCmMl8ZFzgOmwW
h0HTJCbacUkXaDXiM4U6Lgu+7l12tX8jSE2Imv1M3fjLAwr5KtkfHkRIihiUyGzdyCw3dLIir/B/
NrdlnPsPy1nExBTAy51qxOc6g0UGNuN2b9bRiOR3gIJvn45O94VXmZaohOAqVztkPFJHcMKqcgCV
M+PoHqEXaGnJZbtpgQW1OKxfUL7pMOXzh+2yXHVmME+hz8eLf85oLZEmdstTycyV6v7W/AyaEqIn
ch/4znD3UfQ2Phz0RaE9tOUpuKZBLsHg8+xkbqXdmqbBcH7p87Joo2NHBKHnp11MrhfqU5C37g1y
XVLmGVdQ/sn7wLiDRbaksqkTjgRS/E7037jruwvLNnBwzluJDQIV4nGzJ6kWfHtTpFKPzepoyhu5
Pdu8bUAj3/n42s1JhLIu2WHFc+CIlNVKGTrqIulI5dj5kdsMzAluVVOP+1CsxKmWYqhV7ucJMmg8
weLFM/X6y2Zr4OidK/g97JYj+C6YMr+yeJD2IdJqYzY5GiGMypaKYNvxIY8LSQIkZqCO2BekRlsc
us95U2REyXUjYCj6O4oTgYMSRnML7b+jnVq+magR/ZmBG57jAaMX0PmQ2QVzdr6XdnrFUAWwBA0F
I04+LVrDzrLt8JIEiDZeLyBaH8s6DGbHo30bbxInJuzXOEE+O2Q0zwcmXdiu215obNjjhMSsxNOo
62R8kBCnhkZ2gad0cgDGPXVvsXufOa0FjwbqnrvJK09YJm/MHOdFzk48JfcM9Ob4mRpOrQKyhiph
qzlJn/98mib+GyPL7zrussvZNiepvgq3Fp7QqKLVT+uiQ4ypaHyCdoc7SrZaH/6ur0VBSoaqZBLi
WfbSwQ6TzxoaFVoQvYNl52dgtCycUB9nBh+fIlRz8wCr1TxM82couJTpLYTQGi2LwR7vshFLxTYu
iTcEt+6G8ZYLkOA/rzaCIFd/P819Bcs+fl3inS3/aAnMMMxhiOwwquvDR6kC+khefUHkK7XGTEtE
Fey4BN8IgGCyYlDXcKsyA043DAh39wIp9+bm9+oCXI2XoDbhstAz39vNLljwxZY/xNc/E20Lprel
bhy2SAXRNV2x2oG5DVGZNPh2pCY1xFc6LddIl5lpYlTJEuhmaWz1XzD5KIASoYhGagr8XDhSUHOS
x+BcfxXo6XAcK2H+VaYus41++5zYuvIR1Lmm9eF5qdIGFgosD6yo/0+QqFYrvheaDCam6OTaTfOm
nwb7SHUwxq7sfgMixuPelyfj82yOoCmuxzTBIIySKvDA4RvtHJwkRD5pDGo4ROLjYemkXD0tZHzk
3QX76qc6JMUpDPfGXeKgacBOUJ6BGN6ydOCwQZIlTCtKHRCbmCss+VuroDC6bD58upyPnQVu/ADr
UsmKArfdFEeOlAb3SlXPHhYOPEiWmaKxTiyTOoEgeSYau7l1hb0D9ue25bQ3xw7DSpn86SvGNi9l
1urLOXSajEj8UcDD7n78oBUvDsZSwuJd7FNwYxyXDDDtdgXCl1aLBGm4QuRs7RoH1U4crtXlPuU4
LGTm38sIwm4z7VMd9TlLFEc4v7MffbhQBejScv2k/zO+HOfy0SLxtW1Y6WJJ/iddDiqZ5kDa4KTc
P8GnDPG0n5tff9X3vAEhRoIw0Da247iUwrPQSkLIwcdLaHSfAEqpuoV/h0D9r+lv86CONOprPSGA
Ej84tyYDpihLGcK/wYF58hct6c2IMEzup4edQwahTZyZtV743fRb+8/0n08dNlly5DjPK+DgEkH9
aPKZB3sgN/tj/xvcpj2sefB732+KBVpXHHQfKiHbjvEdcaa1AJfLkdQnHp0ipEyLSefJiIKPqDs5
PrNUFLxBOtjCAxerg7MiBDoMnHAVAOUsibLwsXA4VszALCKyspHvp9YEwzCtuNDDh95muliU5ggW
qZYZRWiI2WmXsDuOdnwd6/XazUxWBGUqqvE6ZrmUfwmYJUV29Wb4KCGLjEPlkr3QBzZzoN2ml9PZ
DB4WFGXR3Uc3gZ+zSSYbWzdpsAv3PZkyfbPZNqXQpf3z+nc7casTmLZUbpxgJYd7Bf87fzkjKYo7
FPWOXUrpR1ZxEEf1D6K7cZSrjfoVXTccYCQ6TTAVWKIWmCCGUE5tCfMIkdzkn/Z3GgVH/XJUzpXF
NWm0Ll/blVqEtD2KzB0kOr3b1lrIpVDVJSm/iv3u/QM++aofvEGk6Jc6FnNboF+N2SE9MmocSxFX
O1LJ2bI+2Sx9tGWh8ihs8NA1+xX1jUT+tz4d2Y3qunCqSSaobuIgyTo9s9u2IG1PcMSAPrGrF0t3
5Hm/IPWN8KDsWmrqokB/Nvru+eYaHybMK6WUXhojZcVnlDKyiXKN1Fa4+pfsuDl3Y7IzbgYlCmWP
yyNKUVHFTC+fWVroQUTn6tn7TYWlrwG8OWGcDpoMWZNI7CWF1G1fnDqtzzXIuax16eduVYm/3BB1
8JpTwTd6Hckb/fLjvJrCqcJ4GF477uFCKDjwWXBcihd0q3qGPX/AlzDgcKZ3XlpVwWjFNVopMbPS
2k/IWZHA3cEedmuPTPvyqx5p4PDL13V+EKw0+5IhDW+ojbfBVkP8qcVMalCl1mIujWpPY7RaknmN
r4gOVI9cK4BChtx3f83c7rsOtLSJQ17PKWkDddqqWkVCuqcU+5FA6X0THjiq0nPP92ZzeoqohpPF
839WSdzsZh3i9pbouNFDaxVAO6fa1ODtbL1ItTlg9TSxYIg8FNCLXZymIxGPZrOJHIIPuuMzrZZ/
zthPRBO8OrLu4xbsfj6hpjllJZHprqSfxJEeh+pMCxAGQ3Orx2fAaQVq8BpIiqTWDSwSDeuaARTt
fu3ndh+B8+4Ro0i08e/Ffz5E+/nGBJLuQqCE+RGg+5HxhR2lFnpFmijs32sgDqvGR1KdOypP8E1E
BtJGXBL4k95O8TaakIZfTrN3/Xfu6onIlDkuNZRrG47vaYznu0sfqhFCIOpDfJX0EfgvI00Gg/2f
D6iG+9Jb/NhdH5XgVzx7MExf3wP5VyS0Rol5fuu+9cTGffiMdHRAsXv4meCgbvORaI0jo6I8PHmg
6Di0BjbuFu9bOcV7SIKnySK5MX1r2JdzKLfXC7lsL1Y8T37EWVVcvAhB4EzcIUxCWcbciMf4FiuV
S6aGjUQW9s3mKSo3qjSFDyiR6gL7ZQbg6oEHvclkNP+RnNGu8LBfKRT9en5sPbYmpZv1uJSosaG1
Pygsb5DNkxz3mlmtfMMBjMvHtoAGeR3UXa+V2Mio8yJtWq3Q3yfC/9Pv7ZMD24fxxlgytxF5JqfR
cIA07ATEgAf1OushWig3U85TNFW2Rsmv+CiDm3+MxkQ/cHFTFuKduHAwV3Dvf/xv/GkGbXUHIMW7
RLkuMiiaxXVXf/MitfF2QqvS4Col+Y8nMqk3SCKIYRSR7uJuvgiJ9dsWEubQRIOdrDvkOxAij+Dn
qOUsrstYoxrInOJvD1kWskEbWYkcT5jMVeAy39bIiV0eU53RAfOxoiKYsufUITQiCdPCHB4CvD5i
AytUaCjzpcX9xekpZzg1Q9FQFcaJuMNYGoAy9DwNfM/ZXSyaJQT4CakPVtR2B7s9IADUziU9PkRD
WN5My50FL6N3xWag3LpDl8w7EvEHqq0qk40WBlqIWRjN1yVUpjVKq4X7ukXaGaPigQhtTLfj2K11
+Ho/npFn6oVCcy65UBFdHm18kLEHRP1e3Apdj4cghUT0edGe9sBkCUzhuuAxZXQP+x/r23nyY15C
BYGhCJyiBzbDhg+CpKcKj/GTGizJzcAs8q74DaSslGpxEMi1bLhSgal1abPfjESvFX3ojqMSBz54
5XuljXyGUueIwoZLxVT6b/4Dl562WQsw5Ahrnm7mTfZJfAKOwWqr04OsYFucA0yHb5vp3Ortfidc
Y4G933vLGn+Zm+8YA1sHnbDLiGKxijPjZ2SqXo+/QldSAQjpJcqEItpUNKMcsTy/uF2nMmy+2Xk1
UuVMhp8YQppc+6AdCJK8a7pB/OH5oyDvWeAiRRGR5MiBmxGmqNS9xy3Bd5psoqoxL0d0pHJO0Puw
+7LPCf9dMlXUnEV9le1LseCcYKS4pvxMw7RCBA/8kcwkjRaGxIdnlicGpz83kA61Fb3cuAX78deX
O4/12oevxyDaHyFTiYTZTITMdC1uYwaNBQiRXE7r4zNWM/+BovC/5MyrIwWORpM9FFT7RoFjHDXe
YFy96gAjEBYVKn+ljdaeDGGs5KDyKDjCSP7ZhtoLC6g71brZvilvWCEZ7gJcxNgzZrSLJqbjjm2T
p6J60b423MiWxpFGtF2BCATAFX5WNnmBNTKF1gf1uOyZlBqA+ZWWUmu3+KiTHVikccmSkFVwlgaQ
q1Tk9kMyn0eKjD/cBGx7sts25IJXVtmk4hJuiaHBiUWfR8nHEbbPYDumy4Zdr3rFSTXDO+ercdvV
So3RFijS5SWe9g1uSnr4T0/6CY+bjvXfZfZFi/osGUjRhGSbFMlv6lHZ5OAly4V4RRscSVKRKxWT
nl/CdOQpPNht+mhxSgyMZwwIL08viFNgAB4NWCZ7pVoaF7+BAgVXgtGM03IqOrzU+G0j5QIh8Y7g
nTmUNqRfq/8K1lb3FdrayEcohTQYf/FQ17F6Dh3rUOfVllxEShAa4Otscu2SmZhGQujtIB/FPPv9
XpWXcMH5ajvqZU2MRxIAbfXXW6lp5zh/hOt850R8hOE0d+2QIW0pztD7sZDsWv9mqDaY28xpOmgT
+ZfGW2gZ+j3eJrB4glYV2IMETwVWkoRqiecO3JeW7L31/TqhXLwSoWs7bfX0XObD7RcJHc0otssf
rjzr/ZG0ucYLZB45vLv2gdcrDqkX/51G7UpSVYnrX+19wJaog7WXT37IsS0ctghCmdqmSngzdfTu
Mpgea6eLgTLXRSTwDUA4mGCYHZYoZKAn0i5JPtw93bg0X2T27EWw6xjtSJ+esEvLV/Tw02jO/o7h
vnCyyWez4zTT22nhQDXWxfNB0vQ8nNdAxdQgjWZ9hpAlaP1VcqdnAoe0B+Y6UNa0xdQ0SFlRNiWy
Wj5Mv7K9lvw0BDpXVH5v37uDo0gtk3e6qalsJmOKQJueSpOJjKrI4MWDXCA7xqlzKOenV6Z7wI8S
28g8TmmXlt5piYAiy6k/7Y4IFR6SAVihiCCGfjRJx14FWHaJFe3mMUWYsmMEMjWRKq7cTQIyRbRx
bIq/3ivrDYvSxVYE61MIYT5X8iJAZLHucYvvQV93rD0ThPfxIs1i2tKRd3wly2RuOe4766XawYSu
F1HztKDpl6G7CrKH6IPzSGRIutsFKTMOC/nghklV+eBJYcropNV82kTmf6cFu1HOXZ619avP6yQh
wLDYzUgIIQyZWLYfROkgmyqKEn9zPe/uhuSlGjrf0t5iQpHjaRTIhrh8j45ruvwHG20KsdjtNkAV
oFIGtp2GDNEl0IwDm7wVB74j+18TpDuPe8ebYSH7EG7BTUrA7FYY4z27ycO1a0NzxLjp3wYWwMDL
uAjCXo/yNSxCB7W5AzxinDQ4iGhn9wkOYRY57A4blmkCfPi58NtY1HIKTbS4EDOZyTF0oWkrXIHn
f12UPvdr9mzKpWNe3VGReDQTBKr9LtIaW2i9b/tDgSczh2jd68OVFxqawl68wp2n+rl9tGzGbmI7
2iuhivCxuJduyh1UAmCajLC4XM9yXzlzRzdIh7SsGfQOxroXc3CdPsvFlVqSiUMjhpYdcOCNF4Db
g9eKrdLTD7SFCA4UPml3p+RVe15Nn6kHYijsAJ1vlpCdHYp62u5fRZSfVEuOzdgwsfo9NW10AIXa
DlpthxMold+KfZEWGWdtmzU68RTOt0REmUC6gbd10sm9PJqNcQGEonB3n6cUO6FpWAkuECOn9Gl9
GqIJWPvQrGwI0El4JQ+69Yd+Dn3N/khP1ZzX1PsTstA+Nyc6CSNHqN1UePw46XUy/qDCAgw0jtwP
QyvpuX46or0ljoepKDEGr+UNFEtg2/5uAh7ArTvk0sNVW6cvdY6g/K8ut+ZxXfk9KdWIIB+QbKWG
323Lg3mAKS78r3kx9SAN3iRXljmnx+hFw9OUkZaJNOUI31e5bcGyfjmNCB5l3NFwGryh7Si0893n
RsOo/uw0EIJ+TDOoleD7Aq24rcdoM1ym1YxnQPTOqettS3LT6rOQ8I09FMy+z50BT2YlbcecZ0MP
0s6ckGJy8Q9m0fg6zrSUCYwnWswOp7rycKqJyDres0RgdfGQ9Jz9rWYcBdPZKKK5mWjmDNiuqIiF
R4n3E0vTVE3U/CEeEvJjYLAiVk6c2ud3uVrMwAk/JrVh+nwN0TeabpOJ4DNnc2y2IXZtsTOPP1Id
3+p+pdNK7COXUlOHg9ahZjBJlmd7vr47CSu4+oFww7kWd6OtgRAyAx9+kFbqIj6k4j+9+SKUY4lq
xTpWv89mo11aN8QtrtwLXL8ucldD5LJRKx28YfpZ97BX1PGE/kTjrwgdnv0ACQE2MtSAhHL71rxk
bx+DHyAnn0EjYbEUF9ydGjJLbZQKREymF+F9JMSl3bR60NtGl/mXD+L+YjcXUZrxi+FNZEKXF2OB
gF28bpH4g9CWCiMuJ+NqsZ3yqjfTkIZCy1UDzJXMwXeFL2RwKGthM4Dlb4cClLPK6cmAohT/0wjb
LzB9+6iWXkEAVuZaC702fEbO3ZOidBxmKgL/2S4oh4TlcLmcdG4WA/HdiKWDl7wrT4r+y5EB44GY
DDVMjK38ATJLB/5WyGJvatcM3aJqy/MJLukYSUOO2ZAnezd7KE6m3J5pP15FjA2hwRjDNwmBpV/5
ZJk5unhw4YljbE+i8W7nqj6uF956Gw9glbQsunGBvUqaWosgrcxNqjjxzXKtYGnsszFyb0l4bgAn
wEWWsoQE8cUomFaa1BifK8TDNPff6gl73fyYwau2LmBvpdJAX5VD7EdI4ev2Dk0pW2OxCskfIrLn
INXF26i3GdfHVCXvSQ4J0AoCxy/WJF2o6suXD5pDekKDPc8gHXqM89AInlT8MuKst0yzIHTu4htT
5j8rnQlqOq3elVzqivVRVvbTp4QY0Ol+Rn/wTMXptcnOfmU1HdEjyYSD1f24u1+tAv4thPv6GlXS
Xh/ECwR4uqB1Wi182n/71trjy9sxWE8sXRLJTZTCyluBmi2fAC1kDcE/twBVihZJTL8qFicjMlDs
MKU+QM3qQSCMp44Kkn/Vqpj4uM65l4CSmRhlHeieOoTqDoe5mGyFU4Q7Ao2Zv8WrVfga8pZb89CP
oKiJWy9dHLfW5mrt1HJgrIJsizxJOLV8SG7kPGZffHV+3rZKeJvci+qnwOiP6t3jXBYdpaFshjED
py/h+y4Ke3HwqLXT9L6ayR2Zwr8y0Zt4IU+h0rRYp73auIaC254+mgnTAXO3iVu0DEtcSvjnHMO4
f262qSRyNKp69DLxG0PEAl50201SEVXAXKiFwh9TL8N4FLD1lLMIj2L6s0G8ZRDub4lCi1wsI0RQ
7IEW313zDW4xTTzivsKl0UnwrdnCEyvrDvmmp5zUisCvLC+CeCK0uwxziIfl8aXN43hoevqlbp1Y
k+hfc6JKrewM3X04XlaMUVH6AdPY7b/tKaAdDo2RlLpFlcux7mqCOzfQ7uMZm+pV/r+R554FRXuu
K77CXYdGsAanzaYBANrKFxkEAXlnKlgVQQ8sLv6zJ9jQYMOiWCYdMzOLcdEzeOmUu7mjphTWVcR0
lDIBImc/OSJydGBeGJmakRV3+IbBG9vWmaUu1u2nslqAU9ZkNl8Yz1R4E3w0g0iK1VfwKVr0jm/H
VVkNPOo2CqxDxr+JxHSmorICI3jRbsppI4JlzZp6A4mTAmLWaVVTZe71WwEDdPBha2LB1g/8xshk
Dob0rnlIrf2z4s2ZWU+qL074xvUhoLbeubRoYTyhRGNf6aG5aY0kQcuhtuV8Hl50ZmF8mXt9wLdD
LPAIVb5dHEDbxIt8VGs2ZphDi8XHBkWNSVKTIbjvnEvYHeveNEqpUm15YsDIE0DPYXPyNvQ3inNX
ORkDxCijnDCYGD7+ztINMY+n9BXTECEraJspYwWndYfSLLbRRf0zeXBua7bTh6oQkAaTO2eFJwDi
AZiyyhYaw/sLsIhUq9iYm3ENl7GOytBNG4Xmh9SqrxznwAajOkRxBti2laIUIBQ7v829H7sZQQAr
bFkDOtyB1oBOyH7y1UvIMFeoHrxq0VxbJupFEFt8giWJwxgsVoP9GicDud3Xc1PvXR0DTmWSi8Xi
iNo2PU2LtjxGckPW0FIoJpBAv5WKgKmUx23aO+dSwvGbUBpKf404xPpuO+baRCb+d5rfXyGiZaGX
OBEi/ZMjs3NMqiVBl7wW5SV/kPXHIyz0jZbUipGlP1M4Hn+TFFsbQjt/34DhZMHlOq5VEpPFAmdS
rGCn7GSFx87OGNJ1aMjtv97Nl/jSk2JHvgshyb+g1HoW9Yd3j24zr76rxdvU88JtZbG3nAlyAmoI
na5zRQwrFxPgwQo61Tfszk+Haa3PDamTVvslqcmGa3LAw5ow1Gwlymz0Q1WIDIYjQ69OcEXm6san
GU0+pGTdWqYDdsSaOrHEoqv7dEwDw5l0cAeu8deaiePuQxTt4O+kR7Y9rpATTtggKv03E3Vv2CVi
zEWIowR99n8XFzhxkevje0YQZfnJUBV3ZAnEVzP190UeGU/gEsxIkuuq8rFY5jTs4naSYV8l38Cd
o6ddoWyOY4FSihyzJZIAoYAMKv2VpmhO0Vqix77tYrWB9Fli12AKNnGFCV5xTJHb9pmP7O/6Kx30
gr5ThTKhq4g7ewT68Vfh/E9aSyYknPPd2a3rhh8kbcsdcINMmFxi2zpqSUm8VquJ3mFKo8Pf8/kA
NNjfdnZCWbDMC0msFEcoZ1twq5SUr00+nTJgwdm1gzkEyv4Pb2XoJbzjaujMH2WcPKpB3Q7Dxngi
uJHxpa1YE+S8Mu3Lt+j10wDief59tfNRH0hpfm0SIjSyfMHMMcE4I+h/Eh6zj4kP+hyvp6xxIwaT
FdazBWwqJe+fvkowK7E5zU4cn79VK9XnCHppHVCCa6/OluIpJfOCuY0hdkb7iuB8AWfCiex4+4z6
XiyZC5KXOPV5xDHCkYWTQnY+f5vz3zAjXe9D39ZnTr3VnnXsKoZGeC4tuXtEJa8NqgHZ+rCYWP6u
F/wJGtsPIc9qY865RyOM+yxsFmDiipz3vx7zz3KZLuBjcl1a1Y6EXg5zjZ4GahB0WStTFq/QCzwP
93Plfgr01vgPOLnVivnd3xZORGYNnqi5O5aDBri+6jB/6bDVWOxqeviz+rkY9Sgq+yLAwFx1yE6M
znDY1g6gKGySciGr0+aLW/ZxaS2H3IoUoMzS7Hd9N7NVhSlPpIDPUFlY4lN7ibGZKmbcWVhTfGgj
1v+MuGQt4v4JMQEQx4DZtoRkZjThHkNbG0Epjud9p7+QK1KK8ihhNhS+cYmuLu/RploXn3PYI/9n
L2GcrliPvq6I6DE+zcG0rVwAHgUv63oThKIXNHTFdhwn6in10rLIkHM7jJdL2ZUz4lolIv7Mjnok
jfAOTcGMPcFH5QfgOoKk1Gf+LoDakCFMdBRp7QOk7OpbygEcx+NhhtzivuRThZLsNGzpte+yWzIn
hWFUBHpVPiQUUYhJkptTQWbdyGvhQZ4DytykSZGMVyBJTOjk9gTWgrkL+TfgT2IxooU4Fl2Q04rB
GREcIEJ6Eb3d9GEzyGV4p0Vb52Tq1rqtwvVaqYQDqlc2clQO0Sl73w+W1NlHLavmMS2UF5e2qx8q
ViXKHJDgxHeoKMvawTITEM3zhUyzrRbpiYH8MYhIkaGSWp+4OLR5358K7AGxvvESOiepx7iSbuT+
9ztPVSXW2agpE0x5t7R91n1zWyV/OZkTuKOSrv1LvME2wKfOIMFqXA4qnFiZA6SYRPtLcqyRZK1V
cQ9qZMaDvqOxjhDKsAo0mjL8WQFGGm1s1xrWrKLII1zPLidHvIlpCJbKODtkZkE2AkMxsbWVTysh
roPzBOungjJjm5gVzXO2WyMg/rxFRc7sQxBp6xKm3LFGrmcpW3Tiab4e/RqAVjNKDMmid1qBWoyd
OY+/6wsrqzaYYXEH9H1IA0ZpZNnnU4oeq7NGyAvSmPY51yporhPesKvkcaIU59AFEw1QQwIJuMGd
KGbD8A1R+Zo3+qC4RTsjV2oNz5WqJsylTQ1bGGr18fyH3qWAdEr2zpB+t8MKr0AWfPpBpKLE+QZ+
cwFcZNyjp4+a+aZKQ/tkEqWB7Ar8Ww8HvqgrWeEjU5msiGLf9Lmlmou5PnIqhxi6c79hFwg29xnQ
h0EpOcPSaPFB0Ph0F1teksrrf/bUor4zGxx1iF4o//XX/1cbQdsLA/sReU/zoDlZjS4muSmqyaG+
bneM8YqlorjVehZQMAjRl9ee70U4ljMzUANmzP3dQ2IkrRDkWhp5MwkTeiERFjN4nD1o9vcCETEv
trE0S6zP/Fe94/DlUfJxhddLqCsjHRLE8A8uL+R10wvux4HJG0t4e+keCUacTJrq5EGvKxw8kX2n
oU5Ie73zruHQ/kv4jG1UFPJ7enFSo8KIIZnZ0wEa2l/tij7KL0W0pcQc1w13KhkLl55n9usGTIz0
PPKcIaaK0IEmYgigyKfy/FB8Or7xzC3ZZ768xqXma67WFcJrxo3nG3ZICCsMc/5BrGYLygVI47Sj
FOuJYpV9AHd9xm53HT5l1IJEe4C4mJ8/6keGaKlfXslJ6q/V/Oztp50qAxrrhIaYhk7mOecgE5ta
BEKRvXD5GPBKvbGOKtGic8H1X1ylK9EMeO/MSTAxtz9AYcaMkrS/Zz9JjyDo6ensynQk8ORoxpUO
9+70ehRn75VHIOspGqGEOs8WIyL9X0JYaEEt2k0zGfJu/++JsevjFPtVpJ7UXSk8zN/KYWkegTb1
OAtduBJKXbJctWd1kC5deFwqd1Y9Nz1Swu0mmjAQzX6U7jgBaJ60/w4TrlxKc3wMWHXnnq4kalRW
MGhZu338iZP8VOwM/2Vo7wdHHrf2nriIiYIsQEkYi5Vj5h3Zd1C88qk98OC05D1HY6YzvqMWmeFX
IOsUg4in/mr+dnV+dl8q86KPaXAvKZxYnFBA0B+5XUqaUZrPhEbt9TCfrFH/gSa0j4l5kXPyDtQP
6YxzQg2pnZbclJPlGp2RtN6zen8GViH9eNVOnTCJa11GL/fhi1Pdi6scJp9F1HvjcRSGprQsqRSo
YMJHy/d9g9OGNZTCpzLCpGe1/USfsqNm9DKcdfpOq8zWeoK2lE1/yZ+vAHh80sVCOqh5HJfidya/
VmLdrS5PFvBBQcgr/dlpiKbJXGUW0MnaPMgZX7h/QzJ5VPFKk7oovxv/Yv0QKcc/derSOzaMeg3v
3yVQ9eEw/99jT7+r+R7eMLrNebhHcW3ZCafiKvH7Knz7KHhCQwwDE/NIdZax53d+0YhE3kCXLEdz
AGfovmjfBc3uH47Ef6mrzQiVbgxzxJUv5x9fkNm7ooohuRnHas9fuWFmwa58aB2C1y3WnCTSVWHf
k8px6pxGTCp0PHDdrey8wVlj9zMcN+3fR+wReHpFIGYk6CmucpWDOYtBYxIV1LIRK0xZzPmzQguZ
t/L73S37mRxIjgcWxYNgRrm5wg4XS7k7BafNTfTQUEQ7djK8Jr1HBuKVjqiKy2fSxgi8tKGhK5mc
xsIbg0cBsqdqoFx7FBaMsH00+/s1OP13x3evH4KYvQt0r3VBE7/WszlBTxZrpg64pNwK8YLlOVuH
QhOxXbcRk4lGmbktYEB+0yXcvfVQSLxYui/lx0hsNBFe0liMAeVt5CuVoRWh1rKn2KagBww1gJ9Y
f2vDSXOYQ4tj3WwUX3BfmLbRl6zIG5zKX0q4fcHe1hkx5NQZJJIewx2ytQ7o9MsMx2cqiFgtHenp
APd3CvD2/5ynpzwjiKypjgD+F2S5GKhgY/j7k6vakjVM3WVwV5zem9q1DmdE4dieZkiemzgLhLKQ
AhhrfuFGEBvoHKz+TL4v08eIJ/q1C/y/0zDjg3l3w54cKmwXGL/t80Z0ZSXx2LPB8LcLNQXGKggh
FpXtkrY04QAcK48fdpm3Rct57xvM9833rJlWeueGJS/3e0FqpzgKMk4YTbLcDstrGbk+7wrk+Hhd
FVX13XLulXoVICsUQfZGuPDZRxw6UPgDQFaRP677+p+hpH4XPBDgTzGP2CH3ivyv8SAQoPuFpGft
oY0+Ctdk1vfAeAaxOVNy48TDPxyD86urWixWh3cWh2RCgrC6aMAYZ4jukMFISjvDuZGslEF6zVlm
3EBSYc1x0g3GxNz6oqL+X8TXiVsb4L7HErNiV4FZhdrTwm9FDIvMrd5XZId5uLZz0/Pikzfw9dmC
3dw20U0mDSPKUB7i36MFSMGEDLBVzR7tQo9Dco/r6i6kteRa1MiuRTcnBoBz1TgG3eS/XXuNN/oB
KK+pW+ISRbR6+2kk/g1Z/T4iOUERQ/Ys3Uf5uuQVgtAy4jLHFW5tSIqlVui4Tw1RrE2/iKzApq1X
jsnEjllyINPicSyZluQ2zluO7t5dfTWO2M+VmVFVhAaH+7/93er331m/Ou1jARD4abUCn7GXpN6u
DU33yVFNcR/x1d4LpET6CFjrUYxaSfqZTTc7hrXIMkpauWg8g5jyLdbPHjvyf98GLeOKsrpt7HBC
Rf+XiY8G43klc7aQ+DElfmOz1J7UYAPhyPQioWirhJI8VkYsm+prTmwhzJx52ZtzF6+y+8tw8qrF
88aZ388NJL/6TFNk69AAngi/z0FnHt3p+qIRQ09Dlj+O5Mejy+r+bdEKfvf9XqH3NIJHB0bw6pT6
kJ6uaKdzikpUbGn23UmCAMaP13HpYlspDsMa6IDU3D9BD975WCMdlkly7kBIkqpC4XzmGN+kkCYc
ppNXngVMQ0+q+tc1nj98H/tBRBjSBE1mmgjIIVa6uxuC9L6XNHTwyzTJdsV55yFBlktGisT1G+88
ba5LmWnWE7VoAhV6v7nuN6OwIas87naIRtoQiRhM3yoA9EMVugdpWjOYEEj22cnZK2akPeCjOWui
oyftQ9BETpUfB+bVuRFGbbAZSH1XdN+5vHpgJ/DHbgHTadvQzHsbbJsfSi9F/MF5GmvJayfTH4gR
mJHcDTJAKuIcyT1BTFbheNlOiFOl3MfA3lPs/s5FUO6fibriDllyG2w2DbV5Ma+L7fkmWOtiIaMx
6GbpkHJmqFvavA4FT82k1YNDt2oxL7AOc1gSw2tSEMKLqGq8+MKKtqEHWANkmTMlKry4O/0lMLdk
/QadYuCE1yEWKvbBNAS0/5eGcbAQXpwV8wp/N6TwnTNpyqIck5ut7m/guFheIcUBP0xKNUFSgiCv
rAvArpiUXIGstoW+O5lcETFuOxXe1RDgsVDcXVXNlvK6TfEczQ8nkHx32T0ugAxyzgwHjLKjp0oY
rw/ZxJpNsjCDcl+vLWQDCcjm85dhJPJiBNRqTlG5fXmRDIMDQY468jSfDA55xiEi6HvLuGNhveKT
4L6SxY1NMTBQY0KFLnB8K3QPNVdTSUU1ZDoLSlee7lwh2yBx5ARkQNYXjaTVJw2Izxck6a2BNgzg
eBdzbHYqNBI2m14/Mmq7kZIrZZA5m88y4A+Z2i3rzlZHbSzlunkyojPnUtvv4whpjaTKiFrPwJyP
jiiuCnR+bMU1R/zjOw+m4oM1D88eWwitAC4v1xYq8oZr4VGi5Juttm9BRLDie5k1PlhJ4Twg5KM3
TiZoPekvqby4EvtzDJFbZBsw0TkQzwTmgxSoM82qebJ7Gb8/eLR60IHi/HNqW4qAL4u80q/fXTw6
/XKtv8jgS6nGzkjWuWXL8k3ZejFsyyKXNN5oDpxbt5/q6sd0p93VNlU0aT0Um7UkBGTJrcShbf9f
MGxmkOqy2N5TIV9tgvctL8E3BaoILzCQhZMw2r7ZYOzMK/xkn9hSsA0qIS1wBFdB6TTSwOsqgvl9
XC9Inw2E49hruUANE4KcLdr6ADq+pRadYHo2pmyIwV2jN0jQ3WHWW0WzGKsuSF43jpPeXSclta0R
mS5XrXxzqCcCr7k/BTsmQ8gvchUPSVU4enAw6Ek7gxUCDYnuYc9mlCPjd76/JxVEvueHLIzDFi9N
V/KWXua6SBrUGMlW1dDJejMvVfgC/KXHZpK4E5dEtQ1djUeVWImagJFW9bK1SQa78fwEKNH2jrQ1
HeJctmaDNiN2saEQ+/cQHxZ5ospbX3PquW/70QschDqfnkMyaK0RFMg0MpKhgbRX1WoeB+vwcXXV
Hj4B6RM5VwzQfJsEwRVkPc6rDfBq6VJtBSAdaYzYHWN+VcTlZbBopPrQ5DaQUAOMPBO0Sdk6Mf2s
aRHz8xPBMlX81k1FakSXjMhZ8sjqrNlC6F+83WPtsnbdQPK/ihXJKNrBJ5zAGQoYAhuYR0wofJU3
3AjF75xlIK5bZQ9D94bLioqZqN+IMnf3Y1HAVDZYDkwWN7psuarJJcwTzp9A9+klwr9u96MMMOIX
Izmw0TkXXB0v4/gzdCJMI9BOsdZDSb1EGNUeX27d2ZPtpl9ZfvG6cEqYqyOG8A63I4njMv9me6re
2oZXuJuiI0jHV1rDUDuF61oK/Zrmu4uWNE3ZE1lxi3MOJ0gQ7yfrlSsdMnudnwlOY9RL9kpSwh0L
+xf+PkBVplcjvOQv5TZYX7H9rVtf7B7WYgLlc/NByLckjU4cI9W27U2d8gqMMS7rlLdD8hUY963+
iXAzdqeOkVIXCQtqUOCHlGtrRa4NrbDgEXmbUcMU1O8G5eTO3XxDiK6dxSFY0taK2shA2wUR4QTv
DHZzaOngKBCwG0TpF1rgS+N09i4rZq0dqLNALnUgHDrBY1Z3I7ddWLiVLECWVefjgnhwi0vqhVZv
BJtyyP4/f7AQVpmW3Gr/585T8XZeJCdjTnzzCiU3nXtXTr92/nUcJ2tJJnM7WhX2Kr6WOh/jHydL
dKy9C9AbzbMfnkcLm0rCp5gTAG5jyAADXG80mYHOYClEIIT7iV10LhXCeLO902CGzkciYxh94dSF
YBLXBTwAPUEYRUDKpqUcsZ3CH5WWF5ND6lh7BhdTxV+DzHQ/n6WLMzfOVL5JsJ2umrjw2IaL2tRN
YEENBycaao8AJaP6QZ8LF13zYp6WaT3TH8JaglD4XXTmw5anaMGBBMQ9yjm46YthuFFVSKSdTWvU
6ntehp6guZZCePTarT0fG3JbohI29+a0txQERINqQ2lk3Yt4UzOOrSpIylBsZEaSxCt1tnc+lN0B
zaF6mcILd8ZJN4YaPfvSpkKnHxxbd3d4Us5dlFjcarG5hM1txfcl8Wi5y2yH8shGwIlQOh0pb9XT
0uH5FeR0iwpzZRZMwFUQzjcOUs/4KhZX8bAWNI7i6ghVm7OZ6WIuJZwmfbK+5GrFlWkLJ2rWTQl1
0sucd821PysEjnBo2vmftHPUqVnnHFpUbjIEu4aGcRJzJ3SSCwBOhLDIgeXpRm9sojmb1UmcCv3S
XeoR1TYC9IsFCX2YAqlQdDPELfUzEbv13qjw6xvyNS4/kfL9xZbQGQsmaNTDF8Xu1VMizboF9xDo
1F4a0wmozHsbV9zIoUJkeebWjhLiVg6b7mHrWTknyx712klEJME8rbuyE1U9izh40H5jR5Lx3VU7
SafPBs1kP50a5JqOqr056gc6gb93dHERDOBa877iPkHa/FV2uHfvoBHw3vVtrr38eXfqJfQnl+IP
+cyGJP8Fv8wJ1Eon2r4TciilUXHWTEtNxy3zSr2rA+xBZNA/yAd5gA84DP8NvaEOOU8kglBz6bOm
97pWDq92aXMI1eyZoHUBI7lr3Fqy65FNwkBIOy+c3iTiBJXv3u9WJQuRI2WvP7MxWxecMGqu+JZ8
o7PGYhArUpyeCGS+HTK0Ui9oyIMeSjhyUUjD9CJPqoKDPQmzGbpGK45uURxS6q9QXsQ/yP3NP0RJ
QBhuJghId6iJrL7r5Mo5KM82guohLNNgoKeJ1qx0PdK3x7QZuBv6jE7iVqf+HMiqpKGQfZKNXQRt
JNPt1sbfTktuHww0+OvYu/AfMAa4DN/HImAOJR4M2aZQqmxWBV/gBy5XG+6vVC40cGX/tmcN3xrJ
Qbi53zSgxNwn5FE9VkNBGVwxJnwHh3Xlgul9KnnoTxSDLAE1CQObdMpxX1qNPd9UDbxOLK2rAhNL
WVtVGk+bQcQjj793ZynDmPXbcvE9sVKHHOqas5a6ue3qS0ogif7m2RbDKLWGfvrJ+0ypgraQ9VP5
gpS0/m8c0ROyigz8XQT5wpJ2TN2ZTIkq2WTCfuafFqkG/8nJtiGZinsA3tkceUTTlrJZEZHkHqwG
zV6BEnz/++oCNzLy7OalDjg6H9A6o4pM5a9JA6db5NWyI4Gd5HvL7GsO8+C/PclyDPl826lVI6qZ
9m91t6WN5id/VBU2YZC2VotF1A7QSGN8lLqDthc8469gx8tQXCSd1AdJi3PA8PRyJIv2w7EyCjcP
bVNqkPvrcWk0QPx7X0o5z0650pwDcHELAMf3aePVtc8NRr8RdDj/nouKoTMUchuqSPsGlW+kyrlS
xgH6WrBWdps92BDy/d8Uww2Xk94J8ODkRkM6U49K0+DnsuQ2vJBG5F1IkrQEreghQWq2x37jNPux
McGVyL86HePMnAAJ78oLG4Tp106bqJolc4g4fLmz+0akkiqeL+5SpoZfB130gbx3QEQVr5DlcOx0
DsqDOui/7VtM0j2mO2cf9hgJJoKjAl0SWVvdC/f0DiHlo8v5QDA8i+3cxGpVCql7HR4PeMJb5QMi
vnLEWIfeGFiM5UrZ/cc3+ksXfR8y7bPOyCTkS18joL6nVQj3Wk84vt1jZpNKA5y0mSfPTbw2HsVF
OWoKTfnLVBg4h5UIzr0gaHzpMtQysyu3Y7xm5NZcNXzdgVLTUylQRIDl9peGVLIlesYNOI3hle48
OTD4hckjnnlf+SzRxAw0lECUjMxBATdpoNxNYBC6wE5wJqP+sVUYc0Xf0gRkvcRWXUPXKnGmwvzY
X1+vamKBJIe2POMBpFypqDPVo5LYRa/FhtLxFD1HMGp3J0ar8IL5VhSgUSdnGTlSyk1LLUaSqg5s
KYzAsk64/TY3IFTdkqfpGhDc+w0BvyNTgx6UuVuBHoTtz3CyGxPQx7sVZNDK1DzwfzU37ndR98pJ
k1odqatzswe8ohmnpw+lJhW0NpgoDmtpVswiwYmnh3OzwaBuIxepjjPv0l27cqq4ofNe6F6HGOME
0HHpm7yRXnEB5vAkBM9Ovxw1OSLfbylJkxqmTXUMlY2VjnsEYy3FNakvtUE3EzCvMG2NJ/SMKkrx
vlH9AdaqyTo38OzXcCu1b3BXdoc+9W1zaKyLIMIN7sUzWy6JtGD/jnKFt74DU1MZzjp+vjD0Umug
+xy1GwtHo1mpSagSZC0RhV+oeet3rZ9h18VmOmLKT8ZcR7yQEHUz/kRFUfkbDvzGZimjacsvAWgh
kqKDMRoQVZ+ng2WLmqwOLK64Fr3ay25f7Nil/d01KHziakYMOTkGk6uFT+p/RliPOH2Whz3CvYUF
r55cbEJJQ9xtxAuh8SjZjD2RrWNbm8DvWip/qGKIzLsnQji1imLMer53yGTWa4Up8pZqXlrZVEIY
SwpE1S3NGahZmu87HaPkd0AgVRMIRTvhacM/uXMYnJxYFhS+CNuuoG5KYk3vbSvWun2UCAUuFjNO
68dw6ZkbvC1RbTU7jRf4WHSTqpb3uxnVYTuuVR6Dh4Z6cRcd5n3pjQIFPm0lIz/HIGOVI0+VNq5r
f4u9p8zI/xc9CK4iag8Z2jlcib0DkDk+yygYLY+NeHXsflx0mJLPQwYAt35PzsJx6llVAsQi4z2L
rWngZqkQg8dvfkwq8KS3WehJOWpMf+dKZNGr+c/n2BCHlFRgYkRv1m5chU2OgZ+YP19OHV0YKdWw
XagEccmK8nnxyABmsG1sE/4EF2jk0qXdEDTd16m+eHej5b2mXOKDOKnkl8CuQryjsH3mYZ+Nj8vP
de3OwLjRxDVUbB+U14bv8i809QlczdoUYCcvLLQo7P0wHk6GbTzjCXICexfOp3/2BV9pZN+HFRM7
qpZvL6vhXZ7rMR/jhPB9FDw6/SgMLGIHZrLqiz8vxaoYLNVvdbOPw8qS5YzXZrAUCrYeYG/zsHem
HXZDawpc32uH7vu9bDxQz9s8C0NYp8CJoY3YAKrehnKBQUbiNN1JxiUYnVDBfUgtiYNC+q4LBOXQ
ZAnkuR8zOISwRo7sZYsTPPSfTFAnEtw+bBrtq4HoRGVmpAiNeqpFo4mqfwmQika4C6PtR5U6YCn2
C3ODnopy/nKAmCdEOnivDWQ8iHrHB3Bo2RaH6Jy3CxbubrtlwgmsCEhGdlDq4eZtwOC3aMQIPQD1
khB6yWKlb6qMr6VzJ0RAirQvgNZkzzugqXL6dF4XeNuTYs8LenOATxjZXvwfa4GWjzIgen8GfJ1V
dk7rXsK2jk2qn7OdE9Zbx0ZjZfGrk0iMi8L/v8O2e5oA70RiL1KBRh5vwSLCBQidoRYVlKMCSdCs
956bNIfOELKQAorcZVldQsel7LN9DrGIvl5KFgit3ldMaEoqX00tyWUV6xp82mBTOHLO43toVWZW
kRtysa7K0Rb7M/AHviJfVPHPKAltsZT37ONRszicBXPzUcTmKlHH4Q2h9HWN6Zv0GivU3K5dPWVv
Y1dpnpaMF2UXktAPa9JdMfqipeArG0JcN79Tp7khPd0E6NWcybmcHeAJQgLtHY5ACc9ZDwsh2RQ1
shKwegph+7QE84kMpoiGWsmQoUPLTDIxsJ2zhyk6D5yoMrcBoHKw94vrvemgmlUhsDrReMM6HNn5
xA/6y3bvU3YJ+iJ9Naw9ZDR/ssgsefrhxTBjjfXgyAR1d51RIcTrAdrRfe39MHtITNeDuceUtoQp
rrsKfUmmQjmpMClxaLwqp3kKRUfiw4NEj3DBVawupMIiLy1a75Mmz//JZi/VmlFMam10zVUyYE4W
uEQ724xowWdBcwuU2U3Y5yjUiqQX4eV4QGULGsZZ6K6Qo3Lph6+nPaaVbJvD677V6BZzUequBl+R
Xj+aXNCfhRx0TtAFs+5QnmnY8fXZ4jruSUn8muXP44hXUYCl09mXxe3lf9WmRFom6axxc2ieFrVp
8DgdhxSjzOBp4s8BgKW1ROumrz39WM+R6+rg7sCF61/Vr960f9yIibXX/nIIXsJtHM2gx2z5soC8
f1OjF8CQznPcLsLmnQ52ZNqxHh84jcS2Ecx33Ci3BiCGWGZcaMuFx8ZnaSaRupuNaLwqIOPfCIRK
pRdJxO+cLnwkJNJ383mXaNWvi7vHl9XQpfzNTGB5dfMFTD+6hoVatq8Wk4fnQePglnru/mraHu1C
HuAZp+h2d9SpAcg487xF/VDuYE2EcWeYG2E7agw5lCCtpSWFPDMEiognd5p7JjGe5x8doDanLjNw
QGOxPlxyDwKfL+8EFK2wRdfoVGQQgVxNrAuk16v/2EpEmBF15r6xyM6kbG7+H333VRPrBY2VomaB
3nEVkINststXERe1X4+TVtjJEji3qNv5hUhA+MOZBFE59VIHEylhUqB7EBO6LpRLmfkhbaTSJXLy
2XapfA1POjfaA08IW20VZbCDRAdcle3DRRz8Jeklab0Zayc9Y8HnSj/SbtCx8HWXGQfwHgU4nzcY
JE6VGe7GnVeP2cP+o4PODorVANuOiLCM3Z6r92//JSB6pRlspj4spOgNkIqP0qr4G842NOLMBgXH
edf7Xln/cZPt/aL7XNv31ae8oFwlZfL6Vh8nhSAgA0L7p7Gpcwc6NbFo1NGeYmL3Uz1cy7vNlcNp
BSsB5Hp8k46tpZ8E4WYGKZ259PwZFE88AesIJ0LUwSOX5b9JotvUz8kGSeNNeDurqymzPFz9mZe+
TbJKIkR4EAap2B2rLL2IWAiRXKnP1CA89enVlO2JnfzomlZYGWkBGrtNZOA9B8KF1OIHvQXmZWTr
Wu4/FVeCUhZabmSTASWZxHyia4uZsrHx6bRnmjv4NUfPX3GfesDLRr0nbdKEZHuphoD8AzaXyATG
kzcg+9FJcqtDSYmsbAC1rge+7rYP9eGyNeZrqZPSokZFMa3aYKJOs1I/IdjSdxu/PNPgj1WvJb1M
uSjWNc98zv54dE69imlUPsGiL9WcSEiPvkRClC1kyaR06B5ni4JBJG3cHweo1yVjDQKcizsrPX7R
h8/aFA8aTqC9KpR+UFfnXqYzFUXGclWdamZWpwo9tj7esk2KrHyQxZiGGFkXJ4sWqlw8K9A/YOGM
FT2fztB+PcGv8ZA9PmSAX/5rAXY29ND/JXlcGc07enUWWdiCYcLHV20EThz/0Zt4cWCq2boMLfsP
JOkNAUL9M5tkAj0Frshtj3ECEjdmusVmNbVzFrbpmO2ejh3YRNKC/KvciQa/4vACbJkVzQNb/5lc
VDq01KkL/FHP1luw5CARNBhV74J/WISd3TYSTEEm5o3wRV9/XpekD08QW9A15CCj/eJ4YwG6K7y1
jMBghzFzHHADsZBx9DedataofGJs3g0Yk6oVGu0Rd+QM4EO68kg2MmTyoSHjZ/WB/6gyvPInoVC6
FXowp4sjMXam9ZL6orZP8qD2ACENXBf8uBXB50XVNSaZmC6S03MlfRSR0ughvq0zusDOu0ERt+aU
EpKmji3iwcSvgQgZWwg5K2J/aLE/Y8OVOKosNBzGceOFnQntKlpC5M1xvUVWDbsCOeInWxnxNy2G
LF0N6Jo6bylfJgvnWjHKQ0qcsfjsru+Om9p1txp8k1xb7dLhVFqbYECDsHJNy1mQHuFNJuJzlO7K
vHuebBNk/vMzzYiPJE84yJ4x6UUKq/dGUkB7skrdO/dry6ogpmffUNyv7fSPR0hQxkc8iURa2Fi6
1RfUz0AZ70NJykwou/nazFRM/KQcRFbPPNBSAC71FVUZBk9nCcxqppBSiSQ6sbsVp2/HuGaAn3a/
Ib/gjpyfyfv5OOoyvk4uBIQX271mjiZm2+rvgaO2j+4gsR1y/JbAcmtFkPWXaS/E77zloBUdPXJ7
IJXxAfWo49s6JH7YgUCJyPxT28QIq+b/cUqdAW3hkNQgbDeZu6DNJMZcjMdnPzM3qExLie928DGz
OHMyudYeNb1tBkg1R3cHYnLmdWj71YgGrQWDX4PdGl/hcQfOJv87crcKAtCmedFBhTyrsyO7cK+j
eYLAbmIWfJ29ZXGActa19022/N2BG9MKc9BymOaoTCoLAdUkSMjlThqvXF+Hf7GUt2DnLvH1oKFW
M+wnq/2lIdfojd7YMgKSuTCNRMMqOAYV9xmXstEICRj0InLIC1blvF2uEZkOanPraUA9zMM0mSqr
obRBzUfjNmlMmA4gRNMmc+rNaEVvsKgfIWpN83ZNcYxqwoyLya5I0xbpj7mf/zWlx7Ld1jS8ezn8
88ufOgMxqA7vLahwhIiUdhQhWpeYHy15j5PrOcQt6TTUc1zNz5GOmUS7bOM81+7EVfjbW6fr8P3o
6Jx4mQKigEFOO5p/Ng/2TBzmH48CENW8bQx5Rg9ukOuAYEH5iJDGPTLc7yx9zG5lzyECFV59fOEP
lrQVyUUgFb7AsYdLOToy48j30KgvyvNYuCRSHIjUhoYbR142YKzchrtTUrQ8t74CVeCu/r/pnMpe
f7wlXeC1F+pIpFBSPS8YICp2ZkZrFXwvbr7O0MkLstOSfbSE3e6I5Ut7Id0X+thUBDsRl7y5Jw93
K04SBAAuaby8BIuk4jT47TL87C9QxL2b/NEEGy6Be63fAK2DidexNIsQykM4l/OUHw1S/oFp7dHD
9skwI9fhocSXw+nnuk6VoSYJbfiBlQAcbUFQ/ZdTMi8LtlRZRpRn7iE1QXlHvFCLhdd1kiaPvo5t
GaRr5If6hX4OVJu/Avjh/busICbmFi9d1xPSKrvWX/Oqmz0HItbWuGrUMIZnddRdrV2LbIek5dTc
gAhDHUl6i7F3oiZvbpeTLAYnHChmZd8jQh2ukQnLUxKtKpCFmeKO60BcaxdA7ztKsZghDdeUTnFi
9gzuecYzE/6R0Yqje5TmxQDbP2bsWAyyVu8L50ZM9OICAbuCUo+z4PRGV2/T/qteFcOEfqHsYs7d
8r/wPuZBfSdiQzKokOPmu/6I8yxu9tqh2zXIcqXySJ+qRoTCBDhoBIK5URZbkfVprMDEQVbIPSJs
NFa8WmShYH/E3pwoAVuB3qf9Az+iq0Bdcmye2hzd932+022VPfHJpBvb+co44rvWU+/RwvplHOqZ
AESJt21zuONAFDZsR7lJfogPUbzGXWympubxHxOYr9Q/zQwHGs9NXM+mB/yxLnfpAAh2VA9jBgUn
z9daD/hP94qb3R0CdWx6e2qcCuqoGd/VfBvhebEyMBeQ3NwuLBK+8QmOXFbie88fhM85rnEsGfYJ
ZFXFAznRGZ+1mrF4XHfJYytfApYOd7dM0dLLGDVctbhvjMrq/fTUbO2T8fa1KPUil42LIvs1nYUd
+8rAi+d3vc52tez4WqZ2nPoYOeB2cbRjl2wyLDSpcjygbN89OQ1dBkiPeCyUVGQG6yt3hm3MRdzR
zaA/kQQfohNMkNw6GW9NQwzzJxSGN+qtbtTiosN028NnH+FTA3KLM4jGkOqeS3Se5raxyOkrY3SE
/YhJSC2TqxJMv40AWGpG+nsGTEF2j2gjp7v2mfUKxIH3tIcs02EFI/xM32EvlH51OOWAJvcTtbfy
G5AxNjk7yAHfwxxLW/voWgQVV90t7786Mp8KgYKDiiCBhbfWFQCJYXI5CESljaqSzF2DJecdxjkJ
g5SNRN5mAh9koQVQIAhIlghtO6ggkO9Z1EYDNT6h4oXiN5ljoNlhxV2GH2YnayjA880/NcTsgMkb
awtfgkD1y6O3ci+j5fLnA9AIYaefJBBUb+hjO1VZsI/aBSi103zyzVcxKerv+p1wAC+Z1X1utdgn
TAuWQhkErFxNNAIU+gdmhOcMTBPwueoaacZcyf8lJa0ZbcpR5sa2Fb0W7JgboCLWJaCOusSVyUw5
iQGDCQh++lx4wWyb5szzxEeoopRxl/1qsU55sXQacjkqt+rNBC4A3ijicstXrJ7pgNjsNJkQ4EDx
V8jCe6E/4yJ/AXcbMurUju/myGh/2RDJADMFjwzfQIQQ2Xfihy86EvSX9to8Hb3zfIJV1fHJFDV9
51s9b+QkLddNlyIzcXi0EyIB3kVPrNJB6g+TfkQWV/PEcZhS125xaidk8LgQyzP6h5dw71Wc3r9a
QYtoWDSU38Ef0TPg8OivoNaAwCY8l74qMX2PTiil+XF94aGMB553U7IHkHpj/yMwiGWYwSU72UnO
c7VkjBIdewGa+Fm/CpmULPC1Bp0Qzhvzue1m6XeTWBOgrV+yF5BfvobuodQ9Exh6ATj8EHwLXG5U
p8/GJjlKGRLtEbn0v8dU6I+zS4dzccUUI4t0TtMtcxxluVTI1dRVtgDOs6CdPQKlsyqquKpaWa9s
cH2JjdByDvdEIFUkW0XSdGhJtosy87PW6ITd3rhHvax6TUkOOpQjOGZoLwuQqXey8h1QHg+DDhI1
fQPeUKLq++9VprMelLF/W99SWkrxmcOSSxRybPtfuMfSVNXu3d2i90/nB6YNoBE0x76ppD/IA6Dw
4jH/d1rSyEqcHvLUh2QruWSV9UhzWSKb5eG8e9DVErL647vkcqLg74V6FbtdFQvQGUheIj5RP5ao
GiOVUhjPoamkC2FmrLsfBY+DBSrRjwTS0/hBZ+iZC3WC2M37VJKmTrDLUjgVvXit1P+QY+O2IBDf
iIR+TMi53AJaPFQMJSdsr4T+VpPG7PEOGiA5ShLkhivYgwc5mRIaV4VBernz1xfQwIYjlBjhSinD
Xxq9XbCa3+2/F2OwXU7nBCVmJ8F8tU/k2Rqsp0dDbepl8G4ePTkaquSmdjxu+x9DjKsUDdh93dgb
8thRYmAdZZCz6j2YnbQaqMwou86Adq89r137aWd4cb9gO0n93PA7lj7fMfmt3BaYAlqGq68r/oaE
1CCQ33o4jEHxdjk7GfPWXPEEb52S9d8ayGaOYA+EHq5utLPr8vdWCwmToTOGRZU5H+XfKb+3TyvE
M69+y0eqvFU9B1kAtb6el0JBwynS6IeSAp8NsmLYMy4Q+5HZM4FsFyalZlSteMq8dhN2LG/PoTKU
kyI6jYRC4DOz4SwnPhnGfem397jb2C1ANEmlTYQ3MK8NBD0QOqCvVqMSN/jQ4qGRfdUgqo38rVez
icxAfiFnFrAHXbVi9KhTQCIVsGRARxfA89KMWOtgVDfDQrzCcXuPjHaKjdUr1mbAfC9PD6UJjPLW
52k+7DYoV6E5C+VeDpQpPJHEYffy7ojK3LgZfsf+YlVYPiXM4HNAZ2lZJ0Isitb0+KRXrAS2MbiN
7IFNbgWQcVDls4j6rbE486j6Pe2I3aXFOTlzNgcEZFCQgHEpl4MOlU8yhu286S+aa77R+8PeBu8X
boE2l3OaF/uqhFJtAGEmdtkmwXVZ4jqpd3Dei5UKS73gKPhTppCv7LitC7zlStOimuCFDFTqwzWd
aIMusBvBVs6OZPtLpntoTWcjROxzqyG0bKsj086WGJHO25fCn7c8JWIo85dNXMRWgW32OgXHwvVI
T56RPaqrz7baRZNQu29TARDGvzh5lNcsdeyi9+FQW1oUas1NmIKG7Tdr/PYqJC6qj1bizB4PWGGk
OubYHPQI/+j3DM8GjxwUjlmdvwjRFQSmEmER5ct3YUMOPF/CkSJnK9RbPQ4pSAr7YLfHxDuB6LSh
LB/E5u4/YxoSw6qKCTAabRBOwNST0+JjOaMDiU79dAKHLB8E1DGujDX2hkK9nA1WQPEYiOFfNuFH
lUCGHl+/AW8+MYDBs61qFcXqLvVQZPsos5UD/nJdUyn4TvitfMK9KXFzJiu3qYm8fTfnKsj+rfPl
svPUBi+gZqEaZ/Ur6JqkAPivE8CLrda7Cm78ERGfhOktAqBSa2v8eMbANbgsUeGUW5KjI2T6fT+K
/fbxqal2kjKAlc4pDgFEx58GNVxfduLGp69sOTgM6SEibRPt1hG1ktL0aXnz09sgtFByrmjGazMa
ktqEJ7cWpAQq4IfQHUM5i4B/cZMLGPW99gL4vthDKHcGAaUCjXIP9cRrfAaWS8A1BDIXJaO6yCZh
fugBQtbTW7rlHpCRhFL+jHit6lW2gxdO6VCOXW/YzVuFZdBt7SfZglk9xbukqRvCher3Hsy9nwhO
zZv/RICYf/OVIwHgx98T6eNhB/ETXKyEE5+gxU4QcxZrZo4hRbSpsuZ3dIMqLFl8FneCKZtW4vDc
lBQEhL5lp/yk6CTuiOH5XSpK0MboGGvZAqbm3rchhP3V8L4Ml5JKFcBVBh7WmsfqS0YHn02Zyi3Z
rF0nkHRPlaiF4h6eMxz2N5ilFQthGZdAnhyQJIF1l6azbH97v23R+SXRcNdFGzkora7t1kv6nyaH
QfMkPW/t4Gh0qsPew0kmRCkwSv/RTy7r003s9A9+0PhDKF/N8i2hdFh3oI3GXWsqCJjZSLRlvvKh
caH+MImKI42Fo4/IwLrZtpdwATRrzihDEXkUw7ne2an+Q9V3zKVrOgzIx0iPIvoDPAa/ohc+Z6RI
bY9YjAnnNiPXePjBun/Cycq0tRW0LojavEYNNIK3QqesbSgMHTieD05Pvd+nTTdsUSKnzOj7xp9l
xgtazWLfdCu4z5xN1tgRpPr1mKs0N9uSVmCimM4HscTSjXPye6stU6Xp7DRluZh7VWc4nlfMGFqM
UhpurS6acPsGVsKSiN50pSTGmks830XqMdQQMFxGJNbElGKe7YWa+H+kpzXfmY3roJmRQqyI3rcZ
1i9alCRliQTRTeiiux8jhpXaaaPhui4bAxDiaD/1+OrSvuS2loEdBzbbgqbPg0kLdLUYjaPsZOgc
jaJG0zrRNjF98qSyqXM7PliAQ6JC6pkogQ12RsRhEAB+v1fBqrhI4fEu2DmS592ilrkAoIZ8FhEu
QNwCHyFDTI2Iu0Z0t0NubRFv8oZIf/6wO+V9kOAsEmwWmxffeUzUd/nIf9Snu10cyTF3n3Sw7TrC
gjD7d+SXxz3SHjnH3B4vDBjkky2YLQQmbpfkR+/00pFgQxSrzioIIoqxcC8W8Pg+POsvp3F6Qbp2
ijCObj2txrP+2wRhJ/kHDVan/sOUon9HkporzAbjcB/ITWIhYwHNhMOZff8xLTZpQ2hZ/PPGMbvk
k//3+qmizaLDxvbrM1B5Mc8fjoVZC3NCBUxIFgDBSAXOh4z/aerzRr9x1aGEy0HN9iNbLxB9rPrJ
WDe6RlB+A3s2Pgg9bnbFHUVYHN0epvQmyqAKMalfeDvbQ/MySEXhjotJDT7DaWkkILVB/y9QVVCZ
TPamdwZ7rEiOa+pdTaFoQeBiHVId/KeFIf/WhWxPvy7980bvEnGIvT+JUx71g0SSQeQpcSjnhVfE
bxKiL3zry8Ezt6faM5MMtbJKkA0tnPb1MFI1V44Gb062S41LPhJPzCUQiOHrMSuR6aIm6WEL07UC
RbDxV/tcCelDS3ZkV1FCBETVIggNCHHvUv3R+DyWp1I/0hKWLX4VADaxD5F1NNj/qYne9P5u+1XR
x4sYiylRA7QO9z7LQqbCIMf9UmQYG6Lg05JSo2D4aVNyrZy8ZAsOw+bya/EOzuhYB2lDAU6+2chG
cauVrPT97v81sBtITOQFCfnbTT3qIxYmH+eqAJyhQbL5gu1v/ZSM3R6oSnywzIUJXqnJKEFsQE0D
ioAtsdz9DXqpUaJfXJ6TvZtq2aj2x19DihrNz3fvF28vbUhRtYnHw/9v27qganE+HyBnHqMqOX4F
xkDI9EqOjwAc2aII0oHINLXIQvKnhIkoL4qng1Utno4oypv1oQH5jHlks9XCc9xQlWkYzFkShbxt
g4Zd8nO0zquQdRGfW2dQYZu5yPHzkoUYZRKAjq+kkWzrvLgf/556ZR65QxiiuZjQT/igaC71bnP8
NSVhtBffcSUzLzKgw/0i4sOHAJRC52XygKVWiQ0Kvlv8reavzvy0Xl9AVPkbANA6SKxbt2UfO1X5
+wZTR2FdUywMsvUnt542uqn1SP6gMvVNVZWJiV8AVW6C20sZRa/WIg4kqrXB8ar46c1HRvtXExO9
7YXAQxheBfgUAHSWiTwp/8RQuSusw/x+aldnQzoKKKK1HCNqBLkSYHG94euqcFwodfQsdacZ+YpQ
X8KOp2DltGg+pLjnU0V87oLEAi5A9+BXwjn4X1G/EhwBv6UnEZeP/E0se+xR7etlMqmrRZ31vhYZ
8Z2PPzLOXkYlqHpItoXeh02gLkB+naBxTBWQPGnGGcO+U8thrc84xt4J8/Ez9cCEvc7TGcXQQNpE
iMc2Ga/TWeWc3+Zq36Fa480WfZqvuST2j5uqtqR4lfE6ULdLZXPHBIBZ1qj4Qi564ShllGS6jrxi
epJg4jos65swWnrttfNs8TfxI3jiZTswDjXmMRJV5hAnQpCpxytbt1N7wRU8Kk91q0HVwO8lP2I7
ruagJNLt2tbmJhGi1sb9svP2UrxdDkjbeZSJigiV8d+tm8sZtx6sdOJTRNAjqBfFTCrIPXaNIpHz
8wP0hJABZ5pBIur3XLA73D1wiYc2NXnpvw5z+qD5bqcuZ166F/dCWYgmFWYeBGfEN+PLJYT9eE1M
58y6KV5q2pZEsnaj6+14zi6MoqBBFcCHyAN2Rm2vg3/aGud+6WCjBbkgVuaDU0G85oydh9bgus8v
s6lrjbuUZf/DBG8QcgP4ElOuytUXtlAjVqY9FvlJ/ZN8NhO/Pcjq4/Tv1cyWjPDiGAIn0XILnThK
bEF/FlWYNOMAVbbTU5yimq2GO9se/e3kemKk/aRVhREh+Ds9lUNMVR8nkz+mZIVjQp3g4/SJQLM+
xkAlfcMK+o5deXk+BKPyZ3/w+AFiAzQtOAKnZ/6J4y0rataF3+uKdFQi0Sj+FShuDP1/AP5QZT/Z
EJm3fdMBSbrxsmZDkcEj2A5ATxGXwEean3VuQBtMWI9+xxAaxhGJVlQnb/3hg6smMw2lkMAtHgu/
/MAPus/VrVBcA07SZAe1+2mmVxufXAlCB6KHa3ZmT35tvT6Y8T8Y5utdUbut6WX1DnIjGfdOOKDq
vW6G6GUoUWQeqO1uOFrrsOub7QfhHThcScrVsW/XW4qYVZt5EY48BzswikmEFurjCPHrhqKqbbY/
1TeFgtHKszKywKT6Bj0o5zAIoWM8F8Datlg/GDDnYsH+/jiLXfr64AnYYWKxvVwsfUCLPJHIM9w2
faUrcPeLx5bKpAoIH1bEz63vkRjdB4hClUTHhwDAu5cJw1jNap2QM7L3ln2XjFXufuzbJiTJUa9l
IWbHyX/pe2fOnrahrZvJC3RJYVpkg8yu7Iv1XIfpyaX+7fphSDtyJg7mLD7Won7Nuzes39u+WwEI
R1V0wqGfGpbvRW8ea3EGhBahmNXddpWkuQF34uYcpCB3BZ2PmWxz+U1qhIMRA/BI25Ez3vCX2Q/I
rqZA9i3XYS1G9pkOJbTgSF7wCry0ivaM1uTIAf6IYjglm6gcpyHl47xAELj9API4uT8NQ4BIWorx
BvM2R074ruJlXry+ZnBettXtSJQoAQuym25rX3X67hcmG1ojA8wGiHFIFeELMvVXw6TT00dly9FI
iTd84pgTcJQCDED4k1qmqyo86csFoezFh9M+J0lekoEs3odVMLWNV+q1izXDPX2vCqzUEnM8sok2
I7tFbu7NpmHlgaJMub50VEgiFLq1900tf9bLhn+auWoyqXsooU+84pMvD0rhDHZKNv5Tgr75sHW2
PDXwfmVJbionLMRqsdfhn8e5iOLwp2fURxGmMcDAWkbdn1aNfrcM/MG6azousc+JCQZ2HfImADU3
wRkvg7+UY+yZ+Jouff2MFy//ZJORLHfmWXtglP/ThDauW64r5p2MjVygnm0iIidNa1vh2Reh1yzP
rgy+cdGAfBs2IhantSirF5fIKiQZuywo/KTEl9ax0t6r3miNh7R3C0Df6RtMtv3ErrE4QtqmZg+m
v5/PsJ3W+zQHe4QFH2tMVC4mbwel/MP2q5C5twxoXiJQJIb4YUtFQOpcPblPAXiD4cLUFzJG6ZmQ
8oXCppRK7YrUiaF2ImY/r2AQUQA6pG8RiMKj963/np09K2ecPjKzIsygVyIHR4KxCx0pGghO+1LM
dI2I/mUwjTOhOudAUf/bec3bOH/mt07pgNwbTUdkbTdvSqW8t56Of7wuT01wqA0UiCL1+MWHNR7l
XrIJoSbjuLIiC8ZvQLFCLLMtQNIV7gw78CY2wWMqB0fLfff8qFW10OPHF7qSerXXp41P2hz5T7Ax
Td3GeEQYShMl/+5o2cnrcreDNhgCVZzsOri03yOmTDArG5eVc+IHy12E8bJX+ZTYlJX46eAZeN9x
WIeiSjEqQNPW4fZj4dtQN15qViZsCNRmwM6v5j0GsEnygCBads79oPkHOeCpX0wtBNw4bqu2mfkU
JEMVkASPvD/Qp2DBfrMLi4Seb+2E8tPDvrAlnlrvw6d98GzEKhK7zcc39Qh81m69C25kmxoAV2U1
yzPi5TghdWO7PMhDkZ36vSf91jmxZgQEsU5fJzy28jbrNnMkaR1tLikb5i3nWMy5llQvQc90y9km
YpEni9hItKx5C4BDkbdd31IOwCnkaMq8YQduAQXyYzXq/4TLNp1MyLmCPRr60lcBzx8RjEWhmOFT
nv5u/xqAeHE0JToR6D9XICApdlP9xbUoIwmjM47FrW/xpmwgzl00N/0QGa4EIrNLX9LxiCKxs+ZJ
zo/BB6J55Dj0ds84saos7amCq4gDoh+TtCBdXObJ0FCFWAvmSRgkhetwx82zhCLuWdsc7IVDuk5G
VY5HXH1Dav/KZ6/940FaF1/4pF5z+1ghLsI0PyhKvmVSid4u3++rGbMQMrzsEHAgvFIX5RXL7VUI
YeSnyCAAcXUFrcjJhb/F4DI2bBxjiT7oavTbljhJUKm1JWdUZffo/SQl9KqMwlGBwFIeZtII4+sc
inWhnERlTotl2mJcmaCIe5nZWl0QhmD+UBgXdxQDmvVl/XZpY2gTFFTzWuxsd5x/z6DvTcYZSoga
PaozD69KSeaceg0UjzkF7j9nh2h+iqfZcz6/WSI+146xofa0utBqGn3oY1or2vnQzEbQjqmxzwGF
+FiO/M3ekx9IkCSmJ7U2crjR73hNBbTjg+DfdekZZIzV1TYQGhKOIXVsd5KpDDhrxgfZ9SY2EOaC
qA0cJuQ4KhuPC79vHeOuDeZP3pa+h3S6FD6C9IRlNKPfwQ0AmEUa7tGl9jBJlVwV276QvEPFUalX
xoMGzROBvubj1x15YGbOxnkakL2tbSVwcMWlemKhoL2U5Pk5T/hzVQOX5clVSPKWZMm40P0YpVL7
QHOXMhxvtexzNlSbbz+vlyGbW+Ms3veC8WYAOxBOpmqYhkChK0tFHiRgIrIInvMmKk/CKUTU5TwT
wL/UcQHWmC3zFFZY6t9mLSlJ9Ovdeah03wKB1pG0nF9TXDLfdGtPx0R40oY/l9xQ31q3dAaikS0c
MnresLKvRwrzpcWSvGrZ8W24RasA28KrqxITU7adRPFAbI5RBGFq/wqnxVEaQKyfIkmxY2uh2qwX
kmR6ULhCbSpL/s8x4/pzJJHvMhag9NudxW3PuuDrG5IYO2vFeicA2YlgKe41z9YDh3zR0slhbUa/
mNlgPuYIYbqM3epUDJ0vrd2oNOEzltg//Scb5vD/HycwgasjsMMz51Rrbs5l55p0mJhkmp24zb8B
k/24Am2D4CHypSDlsf7ZQU1wtVkvmUj6hfAufmo+YUXf7oF8kNJMSrq3ERCVI44RicdAZQnrWAOw
tpPhqu+hC2wfJ81DOExfHNdutq8MwZQTtDk6i1HwUqsWUbSCELFwTHbTNbB5EaxZRW04NqKJqU2l
OlLJWhbb4bZXLG1Z+CDa/AyTlfhgQXplyT1taCq05DiAhwPFvNVTG/Od0HaGOkRsSNQvZnPdkrpr
kMsXTdbFqQl7fAAnQ7RHuL5kjdF6iqGWMSXslDVie3IqiTXwXxHozLtQB8eqMR5Dz3TcyfWEOD6K
BVI2dH3WveM3qb09f3BVaLRibDW7K7W2RF3smTGqykwQHLox93ihh2kuTyRoc5Z16NodXoBvJ5FR
JpmWLsrqS4SoAAcrGtcCJtrwux3xGF8oqpZahAfvd3iWYvOVGOivtSIl+y+2n12mK9Qfxf2s3a4/
HC0O/GQ4pIkbHRigIFdo0wqvmfa4PC/GaKjnMM205pFisPF0EwwtYw6SJzJwtTCnESOvIS4SXQ57
eJOzxDI9LKH/+AqoNfRzmJED9bC8xKh31mC/8XAy3zyPDMEcVBKE2/OUDef+nDHHrPrJHus3uKSD
WSW9cz/5Cih0oSGJSxzkV/45odKoXdqAioOImouJz1bJtd55TCdRgax/skG80X2lEb1kGSZDaPsl
ebMQBkOfs1ajHyvBZltI/ahl7zsS2Kvc1vR6YGZu2NzTzzy/I7K5VQBnROrYmLah1nfdEGzGYAJ4
3hUbIrye9bnZkVfsTKlgDCeJMpsjWc01aFHLUFbHP8Wc6hNUUc53naf/bkbXIn5s0vglTTGoUweW
Qje5Dr1X9UH4Tblti0LiOtwtICwkcLl7FI5VjYUMMpO0E+IiF2tebwTRezvFC9l7SlMYDE1qT6P1
QHZ76Cmh7RTFG70EW4h/SSzJmylS/tuEzsEpuXZmjNpCbCwg06TLgB1/6AqzSyVy79FJjiw5cxr/
BzAbvfGruvZuxwYiZL65kiG00s5rRZnNrGr+ylvVauf8mUp4Yq3Y68MLAhNtEjQChPv0FqNZ2fjw
vlfBkqVxPL6V6kP4+raK03MqI87ZdExchJ7wlCq1Jggvve1Kkwu8GUtWPlf+faxiVQj5iwUHXmJ9
fhTjrKl5ywD4xjEnk+8rCLPcUoMTFeDfPP9LxLlt1xRR+3d8R9adHFFSQ802e2/saBYNN0KjB8Pt
dTnH+qKom/ibNCHUVGnYahgCOvQlRew32hEv+50MAAFiy1jtacOQg5TrgEZBRbbGF+IXetjyuL5l
0tofnaF8i4hoEgdQRkX6rB3OdYxLhH535XPzvob75qqDJq9Holjx3PyRaV/iGHkPPyRdx4vj/k52
PkqZvjAleFXCC+DNr76X+5yLIZ3nvtCkjcl1DUoGmGLzZcPWwzCKfUZ8Zi8iigmaojQvdgGnLqmR
zy1iw8jiqyxRrnc+u6HI/NaonJ01DUkSiPMQnXGBo/tSxgbUajhCLsX46Q2MFB0KS3pJq08bL56R
9E3x/y+k9YmGijrxGxGlvS2C0DCTCxOL/Qng4GHLM718UtHHIr7y0RMWCqKXGrc2OLQMuqUv7TCW
ec3M3pVByoOWGrPu+u5xxVIce/z8T2GJYA2/7nJ3k5VzkFIoKT9HXW9i0tRPlolUOmge6R+rUAz1
pSu1PslqRQQ1KiEr+eLFhx9Y3IouSIAPf/XE+WtFzNb/UIOKfc1s2bFfS13omTCy2M3ShBZpo5rB
lGB3we2HCPhg34zQxHVTVCnVGcOiIDJ2VglNolX3ERKG5kWxR9atCOXxdgl4G1jinowo9xjMqJ84
CycN/yF5VFCmkIBAGGVKhAStdB+kWnDsdaQfS+p7O2ryV33Cd4V2/UDZkVi0/p+pFh+cxkmMbio/
a95nZbOg2A5bn/tKrfgLnd9lsorI8G/J+u3F7f2IAb3D9qLmweLfkDN/zEOlDRNS49jdsU74cx6C
4UAbDLDLdtmq3AWkaQr+K1/ve0/I1jghzTgY9N6oxS7e3vjKSXMt440ETlc5DeU82QDtN3dPZXDl
VUPisc+6nlNfO8kVOk7Lterad6Rpz5wD2x6B6e4XfwXIvy1Sk2LggstBX1TK5bRc11+0Rwdmii06
wIqFjS06RP5mP9lGiExzner2Ea5fuXfgwLcKxzzA5cpOBcU8NmadizL/HiokrZwNj9miLfhMZMEk
8p/DmhTJeg7kk6RrWtuqKLCo+Xc2bKG7iUANlY82CyL5mqM5a468j1L4MqRU8a6gUKEokNSiZI4N
+6lLAm9UJx3H1/KqV2AU1kAxMvbZHdFBjwb2EFL882T+GUMDFVkiCdl4YZf0bMgPkVHVlcvrAsu8
B1P97Rfdx/1nOrQirM+uMldQKF62J7uRuv2h43WwVn87yopyGqCbBFFsIEfJB7u+FeN5I+KzbHb/
s+YiQ3R4e/7Zm0cVEsO4FmErBnFV99SsotDOuA+Bc02BRZ+oSsrfBp164iO4NXc5BKYmPAFFCYsW
DIBAJGOEVuXUemH++fsVWiivxM5u8GYt82NJecSQfyiWWaWnXtGeKJUucZmRc/ZP0BlxFtjQQEl/
o9EgQAn6/GupCc9C5kvBmj8w6mNH8hoNqkUl/9zj62DaGoJ6CGqi9bR1CD3uYKKWRpDWgL+TDQPe
KNgfPr/LwMioCofrASsV5k9RVQykSTvQBqrUFuYgF9iOq4LZRAjLa5Douw+XqEPt/DZ9w+lmxVik
+/tTtfBmGDaUNMpVNEy8fmGDh6VSyFfHFodzq5wZMeqvMymB8zNzZUdCXXduVMqgZ4ZOB9NgxcSl
UFrtN8aqjju9Yst27ZuNn4seQGH66wjIe5RYWLwtM4csYjvK0ISpWyYs9Gr7ACOXL3KQxgBQk2ad
2p+m1vZ/aPmY1rVgCCg4R3Q12kvM/Bzwg4kXrBTFHwLiGoO+LM4xQZ2UAVAaLmmsBwRFBEufE+EB
sP9SFE/nFy8TrMPo3iwOdtfsMOqtVlniOrxYVk/SC62cR9AAt0QywOl2yS5BNu+hFrPJkY1S3tGS
SVhWUyN5Mwvz1opxsyqFU/445LXsUHtW9aX1Ta3VHVx15BAHjyUskVbQTUyVV3XskfEmH5bHkWY5
qCeSVjiNvFWgirUsUXE9tR0+iOijDCQFu3GJ8ukFqdRfm8N6fV+qJ6qebfh01h9GdyU1Nl5Jhnqz
xN35S90fQBC3n4qYOoEP4CGLgyiQ6ZMQ71/Ce1NcM/UxDvAYdhNTFmA85jLGJfA/JTzMhBs67v0W
wND64pZZQih+GpQmNgWF5Pnj/cXC3fpVyJXwYs8BoHXTT8fdtTmIVaSGVrq1UGSutQ1SI0/wty6E
Vu4np2ign//bnOsxMGydtPPwK6/rWQPC7U2k3YwLuHbD0L+TV3xCX4jByG5JXKtD6aPOnWmDrNbB
ykXcIMXZ5nvwlMUfpm+X2kn71abq1uztvIUbH5qxzuzdeCaN9RgaafZB0hfwnZylg6EkiWmCuNW7
hKIfSkoD3si/abm1ZPyqgCStO5EOO16JbvKh3H+XtxC5bD+4SX3PKMG/24QS8A1dcO1DW3y8jAth
IpVn6opfSqH5MDefAYgpmAX2FW8fI4/Tz1LyrBgiSJOJXOIs72D/+AuLetv4HKQmxM2i9cZJ/pt/
YKNIkWGML1EiACZzYcWQgs+QR1LHYGIB0fGCRpT6e0RMfkZAmFjvnA+wBWGcnBKzM++GiSLgrj08
mF6jJcquF2RVLBA2XrST0MCTfVV1lRjrevp1JJwEdpJWeZsAYMB+43tBm/DVe6PebozKx7aZfNna
hqCsXZ4D195+69OzzMnaUb6usCmJcfFaOQVU3fwACrI8hopn3X2ln7X3udvcEUm/NT9VMPV1gygZ
qA2kBEAyR83OkQlLEw06lLsVPU4ZBqiAUbavzLkjuP5aXpgDKFK1mNGTAIA94h6NwuxyxuaDQJyB
+3OAMGYUdrFQevCXH6v6EcIj22IgNwj+wVkwiX9k3ACTiDhnaXl3IHO04gI5o0P02Y58i4yZeBLu
+iu6ZwWCXktR2oo6N5bRNnwkxuhx5tcfQa/oL0TEQVrmZ+FXELKkludQHzrMNp4pDnMKIh6VmBd3
D+2lETvPX/c+Vp4HulPiOcmtn+He3Y+FXeJf7PdVaO6Ttwa40qC4yWdJAc/k4BASqBcwK4Jjz9pP
mIuqVhTHfljmYgIxFQmm93ZRMaL1vI+UEn1vULsUPX70gH6iCtZjIih/V2TODv+hwtmLtgrRwCC4
UOqqBk6K1HDUfYfmIpCMKXdbGV97SK9hrqgTTqx+ca8a5E5dE1DOmcRRYmVVa9D6ITKWZptP7ts4
rpy3wOcQB4KPt19sRaaROWKiyn5X/HRknr+c8jeQWRSK5eRgC1NZjFbqhLcEzGrWwPA47wj6DE/K
BHUzhYiHnrN/Bdn/Zu4PndIHAa29khRz8Zp8tb85A40qnJCu5F1UibSWF7nG8vpenuhwOb9Sv/UU
BX2bJ3RkglFVzuJwNk3+WSU69297K3r3pVt8PwGtr7xE3UrOepvC7rnI30Qqow/1B4Tg6eWTuhfz
0EPnFvcJAipDfpzPp7BLkgbH+CZ9xfUwzdUEQNiN7TEebXLikJHipQAbwR+LmUp/ZEPixwHSKGFG
1S/pSk0Qfx1AZS5FIbTKhEI4GwEEkIiYQbYDCaxRaIh6W2iTXNhUR1mipjnb07m9q879fNYAxcc5
rWWED3HofIv8yJdRvDN18fNKPkbmcHI6E0nfW0AOmts5gAx3Q2VHh8Pri9K29RRclwrD1IaIxBlW
2RfcT7J/N9oonu8YGIrNvg32AH8QEbgsVOzCVVnPtsvT0RdDWteDj2cFRnB9U06rEOaCgEgA+SDR
Bge9AHlPsT7eQddLz0WGMwd1JiupS08YxSrz8fluu/3YpGhQKEgRMnj0kCuAr69ZIXTBWqlZxFMx
BQr5YEtDEreAtp2MMvGTQTsf34Hel44xBhIet0kR3NyRi3EdLSCfSku1yRlEECeETm68iZOPJA3U
qQeZhHcjQF6QV9wa3PNmRw18+evMRk9ae6HhaL+I6oleXmmaFodfgVCM3p8daSV/8mgyRUumF13e
qp9qEwtN94L4lUFnhng+19j3ONgQRD5wk13oqu9gLkfkZblU14lj8O0c7usKQ/oyJhcW55TKyQm/
yxqJDHnw2oFewx92pgTE65fpqu/LjhHM4yTpPg+kSbuz4BDwtE9dJ91yhVMRfSHMH6yWzQ3URX4l
Inahvi3ZUfPVyVnkwloakMbaGYiTrx2UnL7czpRZDFTNWd5tv4vm630XBy1h1MH9w2VVFDfMaXHW
xUYtqtEb6dN8nXx8wJgb9T5d4y/Uv2fmFxXMRPONUGcoehO9AUhq8DFdUqc26NwzT8i/HYLnsXIG
nY8WnIoFcQjdcUyoPRnDfaC8LJOEMr+0AayvWGoAyB3tfeoXRdv0HB46uzWdUFXagKPNnPOETYeo
LNZJ+TMP9W4S2V9YJp61MZEI2F84msSR8WuTtw9xaWGJFu0yn9KeC7ar9IcVInjSL/MjT+j0ldHS
7oZlDpmTUW1wy0ObJ+Vm2gAyAaOflcQnPEOWpwmDMEznQSQRJKDs2xOxfLDNZYB6hJK66VFRP6Df
u1j4uxWa1hUpURyOuGWiXiIdl3U/ovd4JxlaWVOPFHTV94TkJMTrt77aQkireNQ81yUWkFlz+iZ0
SuE4Id7hU2dtX7tssjjgP16Ue6wTwmdd11SySRplhAw9rq7G2FD6T4+ZuRWVmpQIewnYLbg/oVLz
h9MUwLi9drn1vCvplMcXA1E/F1HRBXCDFrIzmulFaV5cZrkY5cZS9ui2/H8jU+J+fadRQi9dQxgw
cCFICEJDxjhwF4D5QpFOOMVAVJCPDpV4tMUwsH0nfn9r0lY9jJ/BxGNAzLTlBP+nTVa6bh7QzbfX
4QXP0JpppOji2dozseoWGUXAD80OXYPBiIHjw14otyUQ6ZLCOKenlPNP86x0GOhLjL1YJ8zGmVFo
TqINZH+1Rcl0V9OfYjvP9wqnOhBcgUYSzIcVDktlbAF7LmZmnupGuu8/WheQyRwHBxU3OIQbJI9y
iQIqOohOfu0BEQHO0r6NYfZWx/hYHOdYw+a6JJWkegh2dXHaYrYZGiEEkeJZCFo7SraYe38ryiWL
p/HNhD5H54QaGQSV9dpK7d7zYQIinC0op/sgz6SZKMuOV3OTt33cpHCX4uG1+GTOOGgVNOhFfvUu
KLtc7GBG58mOAW/DyQhxsg5IVr3YxTZ5t13/QjtPnICsAgxOeBWAXptMnHd09awJGN0BYOBY1AJx
m4xQx2FB3avfYdOKk9yyanooew4aLtjuC29MPT5mdJYGMlhRLgFbW/2Lz3P9WR9YGSol2xVW6UcG
vlSxm+kPdMOgdqjW2RAnibriB9xmrloNzDhvr5oFJvmYtjSZVSfhqivqdRM1Sw9nY6B9pzBTAM6I
MvEG3UKaaDNXrTU6fC4cS4NLjERzgkWNwNrSebiM3ybPeuN6Q4s4CQ4aSWeFGk1d7df+cZxBA+xm
IuMKazh6rGhcGH7M53YUhAv09bhdydW7H3NiRvt+Nl3bNQSzr0qqxlYzT/jiRsoEHKuaH3G3vnmM
e1zIGzf22lUQ/kSJJWSX02ad2M3Ib0s+9OxjMO4/bDWTIjKsCOsuPKB5tlOF+aw4gBkg4aInlGFK
LBq3yIg1N3GZGpCLHPgOUiq940JoAUOefXiko4SqxoCh3ry09rs82pqxuYEjno2pkMzgpAFlMF0t
FX6zFw7pMeb/oc6SdyU+R1i20/G+gff2WBLHmUN9jkZmmrkAs/UAG64zcJfuSwmpPTJb/TRqNLrD
yZjkEJTfRri5OR11X5FbqZO+SkYOZUHOev6PjwEtwE0ji5y28cSjBJMn5sHSqeeXi0EhdtKorqmH
TDpUv4+Tbhm7KPb4VAugav/jxvZkI+st4Y+Bfd1TN9aQHFjaSR9kputKxBemi7gwtnZoK6aoLm0z
rh2FjPS62RL+SjkQzH0tV8G/27uXubOJYEwc1MBx1Bu+NoFBGRRU2RcGv8UFdbVkxf/O4a+97k45
GTjpWnjS3xMWFx0Lg6t/1rSWPUaioA+TAF1x4T+vG5hBSK6eEU5Yt2P1UUi7356vlcAtwSu6a50i
CRmwO7unuY+Sg75+BXvreSD/dxQk9PML5r9cfYNew0K6ukoW2hOKAJk2yyyFP5Sv73FQ1EVmVGfi
TnnZkFGX3nhjHGE6MIt1G5RkiXLSqAAokP5yIrcXbFp6l/6mJsCFamxOPKJv+wxuCjyIVaR0g1Yj
WFtROB5YoeEhj6u63LE7BzWwfNqcJN8zPJfCLDfV2FbNTZf0teZAP0nbRBLssxVSe5JCSdFWsoRx
p8SHdUvARBkdNp1wZkqHAOC/hPvaiwCbZGpCzQ5Pz/pD3tFo+MPB9Lwsn3JL689BQG/Ytbp9EddZ
IHGogZFAjq9e3kxTeom4l8k/T/3882AlZwKpurjFrtRqJfo7leauqUQ1Aot04zdizlLXnTrw/M/b
YrmL6ZUP/D+w0jEReAEUcZu7tgbKM77pISixlpg7pZ6EmEeb6sDVPnBjJVRFtF6Lte/4WKwHef0E
F5EOAVD8coW2++/XxOMq1aVW950Z6RZ9SbfCYM39yprtx3FLMYL9wFksevMq/MAP5b6QgVPuzZHv
hnKj4/5l+UlGZ8qVMUW4btPa0dFHgIur9OJHn47tJQgHKixCpCvYqkyq/60kzuTnP0+BVOcFdF0e
aKJNgbJAij4uFPYybiqXvRXrUei0K9YMlAEBcCNgzium7o7tjDDL+gitl6HuEH9hpjSLHkXor70m
Oj2aihiS6WSSBcQVmxF3nXoSFiHIdwpVHIi33s8JSqQlD3wtUd9LluaF2dXVnL+HXVJhVpjjglHY
FxGmH1vPcgUn3bpNsR43KwEqJ5rIqcZbOk+Cesie9qudSnD/HAMZXSw8wXSb3zJmI1pXO9+zPfgD
QiQ27y2tyIXJTAutn+DXU2O7jQ9Kldb4rloV+4kLbUN2O7YdIUMH/8yDBsvL5yEa8C4yLUr2bwP7
jnbFH7Ewu7j7NEQJwiu3Yn7PaAGtaCbw/5IyuodIn6ZxK866q/UqocHhQU9c4u6wlw8uUPbmMyDd
LAf5+FD61/aB4KlTlP9UYc+eeoG7r7Tmf1RYp6+anXkNhtZCy/Yls+d7EnztxHya2k4g7+Oynk6M
QpKN2tKTvW/3PABewVyBDauEVHOOxI15FGntm3TLiuQUyfLZtaymflhncwqh02YNZxrJEb3+IA7I
7BrAA8YZ67GPCDK8WTqlMIwnP/nvQFdbOm9siilDeTfFhbJFnct/YEq3BcDuV+GhnB7Bd6EMvN5P
1BUYagqvS+nCoNvcvbRByUH/ZULGgeQaad7CUmOsKb5Ch07/tFzM4CXJpQnz35P9DbNmVX8SwkjG
nwEaNBuzkzdF7jDGbeY6YUkAxX9FtK2Cix7//lkzy1IvcBOduvwXU/3sEPT0mxlA6FqmhyiOcoFw
6oq7Yrnk4Bcoq9cljmuQ99I/7CXV+Th8QJU3OL4JXHuv+R+tTA4RCX8NUuYBVXA6A7KCMsOUybdg
iPGyFS2Puq6CeRbZCmCkBRDweHcHy/Cpg3OQdN0dIXM7/z6HEQA4UiOytNJC90QSd97I5fEJTc11
aOrqEw8zUVSRY1DQt4YqtkVN+0g8KWbqABaur4Sn4WSZNU1fReaLAqVdrWPw+wb2iriPhxoPNqBR
5sXWihIkM6nsnIG//IV0ibZdwRR6EJTngExrSqo4BreFTEraKQzqoezv52secDd7xYnpjg/bsjAS
cM+ZslBm3VgNTh4v82SQodVHlzm0hI4okb+3VGqlXRy/ALv/j7RiiHk7K9R75LY9d+jK0SO1D6PT
qeAwLEe3aMal5WhMGUM3xpKLvpE+IQUHOBxVviHdTi7/BgT2EVgL1gr8wiChaOjYLsYvDglKW4Hx
XQo5i2emz26ktrOgMB4Ge/2kdOs9pyr8owW7TwUWpJ73lJxuLzs5FwlEbmOYBUKrbS2GeHBrYNEp
1oFbW1iF/+BGEKPv2IhN8wXzSrTXWoBy4fWosFjyxFyflBUq5HGOvzcJytVQza41hVv6Px4SgSjs
aK3uRw+m5UhgPt+04bN58MYzMfqt3vRsDjKlsVfssCJySjUxzqxIEQjCTwfjSV6fcN5+w/lrvxZW
r9wgyjyfNj1GLAZM7ghEodJxbegQEoBUwNAlojI1axnCTCE1hwrc7NVDZHpu8sSnuWX/p/+QhP8S
HU9JE0MaNto51tZD17FJkwx7O9VvlKU5Ydw+fge9yD2SZB8aNIlRFqmwaaystGXqMGSvQ/gxL6xQ
O5KgnDdusi94zvvf80Kb2ckGQsjOpK5QW6cTrYo1vw52r+9qgHcTiRzdGGM8bkGcZlU24J1qkDa6
iuDjJmQo4f7bnmaQ6fOp6ES3NpXPlutpQDB5D59nz1iTAeS/fYjafX6Zzylk00vZF0pkxbBp91Tf
aLLf9GAbBI+R1b/ImUUoL5MuPcncPGySMG5kQC8328HVKsRsB56fHSxG2nFhWSEQ0iaZ3p/6VLhX
DXzFCmCoYZ8hYbYoPMMC/SKbSR0jPhiXTNGSbuo8TOeZ+IA0khZ/DBrZElVXkggQJhOL06U6RLy+
bNa9Ye0EwHz0jX+x3nDXB6+JGbu/VB38VcvsaB9hZkme9tM6/eMbuVBWp8KOxp0iB92SEdQ9bjdX
e8zAHvTYk57riX6+vfj0J84QMrw0Moqfg5m1jHWc3gRK4Li7acRA2k16q7bMb4+mcN4cZ9VorQJZ
cY/gJsOQjX8aCG/E+ZE3STKuaiAo8l2Chiz7RTZyFyKXCYSh1fdFCGACIOYE/Mw9gONFlzE4MDmg
sw0x2qp5Xy4TL4ipooh4l5HQqbQXcO5cSqs1DJpVsqX4Ynw5F29umC650rv8Cj/Dk/zQg2j91/+5
gNAnLKyaV1zIpoj/3mz5NFol+dEN3Ch22jxdppvCKC8E4rdFwkvP15okx1Ff4iPADfFg+mQ5sPIP
5QXzimbj3X4p5NCOHp7/MEE2BBrytnOpXqEW3pFVDnufVdbVz6lGdmRXla6uGQdclufhsn9rS8zE
wbkhwLnySwHGqnWJOFoyhZBHA9pD1DF9LgveB5uTlAT8gf674iuewHFiG3JP1lpHRrLiLvvw2moN
JXAuK6fsedx8E96WiS5x9KN58SAxsWRxjKIijzpGazjsCVwHWNMhVTmHwLgIpkqg+Kaf/6ut1m3W
Pj6+FGp+c6HaEeFyIA3GDdTXAEq24uV/qE5sxlLqZaBfpRl81HOhafIDgGViN1O0IObebLKLUGjA
BfjqeTdxvL0in8Bwu5HQSzOFkBTeWGt9UOwYky9XlnVjRI6la52l8gONdgMnWABSziK0iDN9bwgE
mx2CAfT5lxWsUgduNVMer3wneiMRcQGC6cR1Mv4LjZgCvgCLAPER9qYMTfgCDFYcZ0UxmfxiWmQg
ZPKVLFgMOKtnZpugIckMMeY/p0D2O+UM8fym53iAOXxNEu/nJqy8BQfWxr5cBRNmdY4n8THQkpUv
e9L88kLFy8I0uuvSSSw2Ef5xyOFWtyeXf9Eq8DRXtY6eHvPM8UO8Eobs31gZ2q1Ffzj77/LaSdQo
hYy/G4lNG2nRcLYDsQi8CBiv55MyUsqrQebABphTM8vyOM1ctGZDeBp8NTePW2ysUGIzeUVyIBz5
uzId5lrF43jfjmrE7q8QlEkojlU/zjkq40FZR3DrkTn+RdE+lJPkdawQJctxXUuw5skpfjfTcheZ
Qar3hCUfh1VfOvaJ3vkolBOIFYqMAEStW3AUMl+IwfI98e8ZUlFV05v3nqzRXGq1RB8Wai/tHZ7u
dvtAzTX1AqbENt7CW7NIKanB1swWHyyng0rJcVRaFgdBOTTWV2G7n6ynCcM2GdNfLygRcqyDGFFD
uwmC/Lq2HCu5p8NNxKmRY3OUk8jnFKxBYUMikitprhWQy/4IKvu13qA7YVzS9nDxgecnKV4qkMi9
M1knINnjnWhj1F4EE+llWNSOSybRNaU17W76zgU1DW25Q2QSk8BR730M0AqKbk3y1SzYIxiQYe27
txKsJR0e5i7D9S5krIVoeaS6gfG6aMBulaKCNVpXk3l8TLuHgN0ITn8b4bZZJFy3yu7wJtRs1i/O
XuiiHFovNwIFcTBo4d3KXNh/cIBdRLoC1iq9typQv6iWrrHIh9hwHJSj9BbHJjgUTf95NOsifpNM
w5s7qpfnO9vyRLyMyX5aF7QB/FWn4toGAtXuDggg9nb6cJg7HvgHGQtAYEQRjue3WfoAB30mo+bL
rfGV515rtkIWPL+yyICSknJktzaZ+IWkqlMqIXq+04Hyf9zzgBQe/6lUM60P/Y5xnG9VoR43uQCC
Em/jcAE2V4APcWeUvQh0Znmlh/VV5hL9GKLbTBad40bq2NTXKmVhPgOG5nArHjNQJuzV8AXor2C2
YDICLFeu8j/PpxZmDM6XdClTiJf9bj+4KSziRXiEPNTwrMj9TKpUVWVktnpJaEE6/RZh5Ai0+z4k
rgdW8SMsbJ2X1XUhY4gIySdElWi5gupK6WkEqk37cskWlYvQN2cuzc1hD8OPum070+gO5FBTbkRO
fAskmY1usnj0VYJkhrGHI/Wr7cxHDlJRLr2SmwRcPX6p5no3w7Z7BOXSNfcpnPdMJz/92ja8gx8b
t0xJvwNvjeS0U/KYMc/HZi7oCeZIRoeHIs91H/JPlDOmiOrx4cYRVXv0emRPjVjU5FbO4YV6MGIM
Hqxt8ausSbgWqTILrN+0ADk9bxjCsZ3exyGng+mxwtEnKMa5K37ZdiEJwiHZIFU0fx0UXNaQSgTz
NIR4XXY1P6GTx29Yaufb1vLZH5Ot0sxsLW/+xS2+TSb/JDP1ZXLMKlHO+PsNJFkDlv54m/7j38id
Xtq1BDXAt9KRCtEgpxPIGs3+vRwbbGK76s9v4wEMdMf82R6DKB2mI2KjpHRSyDa8U246lawwWcuo
8cESkH0ed/1Y7Q8VQJlyUCjn7PpP9BcFWo1OxSbYst5TyofXGYNDMbGwv2plYRMeQ0i4x4fa9Hgk
6C8TM9lxxtXa7Xx3tQYaq/LS2cqJ4oIwYBlYzEXjd6HxW2Q+NAJ4ePt7cmJkaHokt+R0dbTqDw8E
qlFMXqk1OF/OEZuQ4cpBC+emlQ4z67Lq/HfMSV+9aJalLS9GGeMBO9FHH+GLD/BgJTlnaYaQP7O6
LIGOPfdRmlKajZliH8u2v3LDm+1HuUYArodMlDwngt12l0od7q5uFgLXlL50iocdATGtuRUNwqUt
BqO9xiGPMpuXAuL+vNihyPXBFQknyz4MRIAz8kKhPW04huGvUfQbJUmtnokYWEY3JpMwiDPrpUKf
nP4YTWdGRpkJvdj+vmT9YXZbnhoMJQlTaA8dW4Wbi9+/ZVml6z2F6EJSYiYIYGdpOnxPyxoVPl0t
Mf1p9xvS255+JoprN8HOsgqn45LPUS+oi70NKmhXn4pAXlhetrd48RB+U8s/SJdiMk5IpmOg45A3
qwdKHd+Wg1Tw9yTC9Hpv+P6zpT/4dcCscC1cNS6qSpd2Nns5PHpX6YSx167rnmqRn+0YtjlEOERq
IcNdkHqS+7jAt8Qo3uXxBHFydlTcr3r6NRk8p77+TVzTIQl7plPM8apG39D9O1I1YYQFXMobtRVC
WZYaSZXkGEYvx7iHQuBITGuxBNFA3HiAgj8cQbsG/dHhILoqItVHT6k32sLIuAwgMubR/xs2K43H
41iWmAPiNzcDZwHL4rxvNq2RpvNjxMcBM5p+5FbxFrj0rqE69GCYmspeGV8o+C70k7Xtefddbqhj
EPwFTlKSwNIBN66ExFbTN2WRRixzWZFqSPUre9tYW6Lr/1EY86ZZ5D7Tjz04YvohJjAjPjE2znzC
85hrG2Z9anZcPrhV5M4X7uONcqS3+Gd8wR/S0n+PvyF1MGwu+R2johPWuHJ/032wEr1um2bfCeQl
0Vdt38PLKH4OOANuizl1Ri7rwQDO2niNeqyDxe0kKy9vwFABrNbs9MHMeugfHgwVNyFUMwH7E8IK
k7R1IkxLMAzZHHkNW0g2hLvuD9YNG/tEiPG2pXRrq558vVIx2mumqvSwtvx8klu9bjSolvsM9fFI
9VE5E7srrOJuTot/iwhXGvQQ/Apd0UdXPlLBsqU86u07SYqiJO6sS2VQJXE6xaFw8t6oBusqPQHU
tTL0kUlzCB7mwv0MR2DXaJcBYI9sIcvzhnkjduCN37MRbQ81g8G4juxDJvU5E50zD3wD/OcEVAvm
QnlI1tP+0ZCtUNRtyCorwBLjF5dYilMsh6+03lCWGX613dgIOQDojuNHeB9vF284a3Hb86LBetn6
FsA5PRGedQ2SJZi2dFd8y7PyiJwllPf5i9WfsURL7vzFPoLV3JQKiZxACqGKSllL7asv+j0zeQ9p
KEMQegXetc+/Em6feVy1WAOg6vpmf9d8payTur6pcUelx+VJ92sxbiqa1xtzvbiKq9OchO/74V9I
2tufKfIxkUkLdGsRUEp+1O8P4CQSyUAq/ErDzlIq/KDCXhh8kekF61k05Tr0GVoGYepFQSSd7Ghp
VO46EJo15sB2JwJJQoXhWUZEiZM3WcDgWg1ssAl1no+z1asN+WGcCCL7xHraOxlGnAiwsFEkbdQx
IdosMbQo0oXV0c0PtvCMFRwuCX1HOWbHA7WJaG8Ge7h61EHdiw/4MWNUi2PO5dG7IRVghD5jEVNv
IXkonlyMBAbD2MRH4GdAf/BvUh/3B/BGPHODt8/3n5otohRIRHg4f8HxQaG1hXMHTviSlahEdR4g
exOsUyPGdA3vMYVgo50gYv7nII2TAcpO/Ydky1FKAQsx4/UUJZQbcC4R4db8AHwYKykS3NScIozU
wUGj0w6BCzzvpy5NnuDwdLDtncvEZM094H02WX8Rk0d6ek+MkrTlHoBJOMQ7DveOpO38720AdpJG
3U8jdvPEA6EsLRrwZTi4LUE2sokrzytWYfvce/pEJrw8hjTks0y6OBZfjyl0SJEByOgTgU9avqr/
J33jhPzDB4TyKQ/S3UvWyt5A2m10B0ZZHHpsGhZpc5GZr3sF6VszjNZIZQ0szPUFxMHWfmffgztL
T+yjMuuxcBU70oehZBg2QPNixL+oHkTtLv9AyLa0y3Jab58RyqXpHDEdytWlsqqWmjftusRImjf2
cmOYl6aPcM0hrgu96ftjlCIYbiteRY4jq8sN7YO9RLo7VkNeT4ijt8mh/Y9FNnncnwCC6EmjBqGv
f+RNU2u8qdSiyqUYOgDUSfDHxIy8ThIbmizwlSAdbpfeUgR8AiBajlRxJMu4sv5/M9JkII77EiOm
b3S3vXiIpDBhLxCVCg9a42Gpuajy18FuMdNlio7yiMASIiL2nsEEq9yLutvKNdCYnHzCB5JNm9sM
DI/WI7yEdviJnOlJDOBk3LpZsiBW1L+JIlaJp/+WbUTZ+YsMRn2b3Wgs89UY20vByXcnLRCzlmZY
ixtYbfrhB3HT7BjBRWh95ONNEHxXNN8ivdu1bNiFQbWKblPt5Zso+3TzloWGabcqdWHLzBZd5MJ9
bx8cdQxfbX/REdVdSVXIRNK57LstGUy3GE4+SRw0uB0in9qfn9Jab6v41xRGw3jERKcMqEK/w1Xd
P2/kVD+zsdkwoqe4EsKtCHtAn6dFROMfEm1iZ5k+/Bq4lkPF5X87xJaWCnlLjxfXHTjF62lJ2lf0
iouTPY9p7NcsHCAhBMj5xbGySAxIFPPk3NQibf/LiIqM1A867Y+V5dkJE+FqbhJzUVbZhkJrDpZX
5qyAzCLM0miajGoMgxRX5Ackp1r/42qVe9RUmyJ5ZtTiYlFpvQ1XRhakB3eZlqrF0ee/53lQmxBf
8kE9xe7bxhByJ/R3A0CvHK8qKKmvtObWi2ndA8vk4rLso+EifMMzsTVG60sm9suC9N8pXnHzzBZz
yy2De2bcqJo8+bue7Df0oQ3wL2+N8lhsZIKV9sEbUVCt2n9uGuvp5PY1+pojDYgxImZ0csVD3zpM
UnkUtiQhx1dH6bXZtTsFT6CdNaiHVfO1cNhvdQ517+fdkl2ssO+u4Uyfv8YoPdbzoCHhTf1NofJS
wOjjpUkHER1/Vh/B7k/+GrDf+cDxHGTzYUUXJHcH7giLac0gnD/raSd/uCZmoQ0sJNirUGhG0CBj
VwjCPj3ALdrX782ieckAS7czffcLYM6vi75BJzl1AIVVobeKT5++vlsN+q3zyQppZrMgf37tWV3s
WQBv85otlTfI51g/NFhSkMmNZWxCB5D+58/LA4zDpdjGGxxEYdfT1hjRuVpyyTxhJe8YsMT4gD4N
KD3x2BOHhvmo4ABxngQc8HjIE0If598ZdD8iiUOhgN6QvQmSThoXjbvKCUwN+XJVELiiPOkzLJ6C
8riz5z2uwZXrTqI/2MBi+2l2f1nGLen9BGjm3hW//ZraxOE4qg5W4Kj5G1WMFzyOJD1QuaOp3//d
Ejq0SBell6R7f1UhsRPT8PAF6qicoo71sRLPUJlkeWeSclvbXv3nALNEhN1IxfJ+fU2EfRWfgRdC
PdU+8UEp96Guy2DMoap2Ni7aM1gTcEzQDdML6bjXGcq5tLenqa51MrgauYop8rxA2E0gIl5EjlSr
bj5hoWXrBMIPhYHy4Kyweco2VqyXTX7bWUKG0htBOn8YL9hgotn9p+QIo8265oZ7wZFniYq4w38S
UsNa82ATj7mf9PMdTPLFUlxxw0UFidFLF2I21/YC/TQMaU6mrm5TFl8ZaZoLzAiDZIAADM/kRVTt
HrnIz7MJAj5G5R7pUlcHllulh7Mb8fNzPjizdO7/1/vlnqKzBrtpZg1GfdYoipI9442D1YS8+a2R
XLqcHH1wvsFVJhKxLIkHrUsgitgyatTUQKQFN5eQTlMyn7jVbFwZ7c6Q0Elnqmu+RCbAag8LU0l6
1DF9m/l0iWFe0sRVxJdx3qYLZcl60wWWsUIIx7fL6xyYw29b0i16uBqsU/B5DX5KtRlth816i0Vo
RuN36lVP6+Msc0UufELSEuVrEGcF+D71mRmvza83MamOJJi5vzStRvkh6vU+BjWc4pSrhr4e4fx3
2t7Sq4ntLIIfm6JHc8SAcEQPzd2QQ9V/JIV0vfghh2iVEY0d8k2OdLh7aBr6md4cfHbFmu2d9VFf
Ly+mzu/Xetojvc3DW1hzhA1TOZBKvRPsEbDN+7YaRJxUZuiEB2fBJ6mPF5pBs6Nq9yM4diloQUuk
6i7wDaJ6SeBLqkof75w5s/U1kFbO90pKkY+xSGb4SqQ6KzNat4daVmSQsncE82yiHG5l9P1Gsz4g
TttEOjh/2ReU0UU4LMmiLo2X8fOtBEma68kGp2QMidm1K3mYreTtJnpZRUT0Iri4cwll5xOpLx5F
95R3pP1QobKdB4D7+W+uYFYM3pLwr4Mpij5Rzsl1gUcbuDkKJwZkn+TPk51BnF52hcGGKkEVyaek
Z+5CpsbNFc5MlQMn20XvGUInuihenKwNU3vO5R3vweVk95hV1Z1Je2XYvRPSzlwMXqjPk3NDtbPe
Qp8jjma6rroQU/x7eWtsmB1x/0rXp+Jg0zRyZhadw//Bx2eA/pRh6Z6aTHbgWrij5/yPyUwz5fF7
ixvY94KlykP3C9oKixQJv9DdoFPx2x+ilyqYxlB6qIZPlFAPPSrs1RUT+eJ5olDm21I4klbXlFPg
FVGvPrVWUCSDEwDCbsa3wLIE+X49cuKcBtbxN1BbMuWUkTjZGVT1rar9puDOe6B7bhxlbphveDF4
/oXjeTi6EysARra6BaNidFR6ydvcTIIpGGCTOmZBnQaO+IE/koqskonsv+nuH0VaBGIW+5qeRANs
dAgMJ7cza2s+mu+Y11PVhc+URzRFIGUfjCBwuDmAZnZOoG2dV3aEx2AYTkf9f2GflpkQb98b5gR0
gqsP4QgYN/VPlZgqIYOhaW3t1fFo9XFCiyYtbxt1S55IE1r3BN2YkCv+b1YwYQLYEEK/kjrdlYCY
w4rlN5fyeRdbxAD2L/ZQ5QnwCo6LvPk2fw+yawY0N7WJ7T27rTg02XaKVs6uRrv+maCegAzq8smb
2+oV10VlNL7UgNcrgvIcXLbfVsfRRTgSv126NGr+WEjmLI3Qzb3QKtan4UMYDtIWeoKao/8TNbSN
t4jtkvrh4HTMw6+WQXTx5mXAu7vkOD8BvSu23Bvkab/CKMZ936JNWWNqUlHqJNbI5tTgDwSkFjo+
jkpA/mkaikJ9K6XoJZbrY8T16DiJeDeInxKXsWYAM+AeJEMiYrN05nuCVHSouoajgCMFaAKomX+V
7VzifyaQoigiYzVZ3dpEmauNNnVDBK5glEg1s43G/wAFNvZAdS7dKoYFGw6WwdA2b5JX+1fr7/iX
vumPrlLYACMoD9xtUv99IdxAtoAHWmY35uWnDE82qQckBjA/Vsi1E9A5pvU+X9oLPMfvhKawtsWC
r6ym6BmggNkl9B2HgLb1K6/tPM7oMxYjymVRn3D2597o+zCAsN3TKmn5K6nEBC5koCKPzxVIe3Ul
43oJTXtr9s3lzKkx8BHOnvPmflvfBVHLHjP4vFLAQmUfp8N5ZECpORQ2gfp7kZVj15aYlBBrPeA0
18WpeDH5H/AmXmo7GRL7lTRvl1Lc7IrL//D1KeIsePuq7Rc1RNREu4b5GycB/TKjxNF5RnMdqnAD
pqWb3Z9xweGeMoiAlMgXlSIKlh+Bc03yLPDR+yKGLAEc6UWE8DNmfAibaZV7PfQbAG50h4huG+Av
N+RrmyzEcgJGDuYGeIVQS53YYtc7Oon4r4u2CSl5tkrzWt7r4QxF4FfBua52vtgTHy+bIOJJi1wk
jUSC2QMSyhs0yNHWq2NIYBCrbRmpefvysfirRWyul8iaFJ23SBE3goYNnPyUVVJShVn56PTRTQQD
brOEtuWHxw689qyh6yfQfGc5wuxgB6J9vwWt7T9ku5IAB8xTdwAVgdZAjFemKepXy3pxUThbEvyE
kL2TnSKENXEEOSWzinmB3VlZWocSp5pCHqdVb4GtlwPFP04gGhy34f0xWuKYWk243t/PLKzv+Fjw
6MayOmd5IYMvwjWpFB6joq07dHbOKcBU+1J7VeYCuop+YoBN7pk3Ek44z9FGxxD8HMGhXsf3/loj
P9CnP4rF6SokHMjF4XeBU8PJaeuavhwh4hOXafUgU73wQBre0EqQ3MKXgxanUVGDMsPXiOndcBbJ
qx3aEcHBQ2wTCbMIGjTjx/KVF6Jvk/x94LjIHXAr7QS0stS8vg/rj4A16/TyrnetYvwBkCKbtLSa
/Nbr9y/TDPsLJcTZJXlwCobG2YU1uDAhHTDkNwv1qSVhkUlWVo9tpEDUUQVWinYorucOTrQDo5H3
LgDnoH5nWJMn58moVq0dr2odJIaoFu8okbj0czh6lr/eOaqx/hGAC1lZmLXnR8nfeZ2qm2WGGIU4
cymD/hnVtkOY1Cri7+jdh+RlwW5VuuqpQg4uz/Q4SaLN2RbmAzcRiARBLOjLDZRp3Q3pq0FghMhy
t0mlvYEDi4W5XH+bL5XrBEvc/FfNx19eqCRpWb6haHmGcHqNCJWN2IYluZk1rqrB5DnEYYltIrm0
JOzAqxPKIZzXfrkOEY8D28b1y9c8a8jvieaY/QOesfq3cCn2CZ5GGXIMq/sL0fYOoCk+I+d48c1W
rUvJCqnJRiiM4I/dmCUl+H7J71ZN2IMFM5Vu5nb3yE23H3Ywco0+8uTEib0yol91ucQ9VFDtbbtU
e9C1RmpjaFjxM4OKbgTcnhJ7J42VYlOrMXzKODeOCu5jGh/IUSZymbgoEmcaw6o8iNI0eHcx9duH
ZDE+8NeYicSK0BxtcQVp5W7xplepICG0ZwNwrxtK6xEclX+zDp1U+5Mz2NxVpEU05n89ymzWdu24
mbmJD5qlzMGe2G9y35cIMQLBByjLBXnjcjjUWYu9PDcd4I2OLHfKi9kWVvTKDezaQF9d5CbhYPQF
HU2Tp8ehMH6zyH+A/oLHMTik69sMPfmyiR2WsOZYPY0fJYxevz8n4ATGaLu1FPGezF738XkU7bta
UXQlh73phXT/gICnEg+fsm2NZlqC6jMqRNO+FZINvolZWCu5++nk19x7PD6rp4yiY1J9SDC09SPZ
UobuY/0DLNMujF9g+tBruUwN8wcaVnnJRdj8eCtjipsxuEJ260ZiTmY7Vum+REAi114NH4r5cF+s
YEEIQN2OC/hB5QpxZnxP9eiNv6ONwyPs4lECobtbhUBm74208sR4s4gR+HYgR6vTIud0ibofGMEv
2Bn9Wi0KtyiDlc5qAkcTkPTf825MHdewIOpPiMoPUwGzPUpW9VbpzmeuS2Eyi9Pp+K5G8nQnsafT
yZrcO1vMApsqgxNkvQB5XsKrn6YvqM+NLqIGrIlgnFAttybuE27QrjUtafwpFvL+JmZUWExG7jvZ
XpIN4m//wruCm1x1fKP0MxbTLFr9QksEtvkqN7U3lSnp/ZqmgGAxbr4shFYmG2BpJ0K78uME1YXU
fM3ReWmZ0LjdZwTYTSQIR9egxvdyNqcEZ3XyvrUbPo3dZ4fXc9xEkj4D6GZSfFfe58mLdwt1LzsW
LBacnqvq7WDdBMFRMl9C9s8n3pgCF+e1T9xYx5K3vOVPx0FXD0BSMcdFGqp+nXkwk2AfgLdad3Pq
Dmoxums6nhrtECCD3SEzyltVXIan9pgUJR7aEel+Wtk5mfBEFXXuGIFop44V7lmFKxtmvc3m9WVU
MgFSp2XL3r5aTd/ftsMNOUB9/2FcXxBTxR1Laf1HrYQXNCOeDHihtgvdDE/p5iKPC21cKv6LCBJK
YC5mXXaiZ+4ZPmpxi1EGyTM0tp7XHzyHI9PxMG43Msm24f0YHWabDz+hOO77ER7Y2/lk3/EbwldL
nx864oCAUmq/g+mDvwC3v0YpGe0Vj85YTjgofffROhMx4TA/mCVZhIMnwKo/oej5oJJFAMMivylz
eWK55u/JfKWZ8WmTp4hyo5OcwlvJOv+3x1QYq0R97DQGGHYbD/yIvOuZGljEXQzjtHuDzexJnzhC
FfUOogHdhIWIXLyscPb4jef0KtVIBb4YSMxRgCWQ1X17GT/vQSHSM5mY1xRmAuNxOZURNO8v+FSV
2+r4QjNbtWy9WaK0w8+To8XM7C3YY14qNgrN+UA7wTZsmygvyBZPf+TshuaGZO5UlqMFFQ7JOJpd
CLhWblwZMkOYRJ2VEj9vhhWWd8tdBerdm7X7qWBShL9gnsk2v+GaqSy1S1BOAGSPC6uIBfFeTXag
98rVK2frgojLH/WYq7Eue5oA0NQuaLcg3vJHn0z8patQV2xBg7oJ1L6xbOgvU90FTRtbMgmvFU58
cF9o4zWftOnRAbZryRVVSVnU5bOa5l/L+nAZfCVPfJW4EgN4YL1f/VJzSZGY2rm24AuxdjZ5wP2o
C09C9ebhKorkj5fU6PX2jsIe77cRdgdL4LpaAlR+b750pbkqj4cehhUcFd11f7GRi83TPPu9smDT
PRVfeeoHuoWFu9TcnqNf0n2t9En36Ahbs7ONd0o3Xb8xDLApffNgQOfEmuAnzX5URgOzDQ5w0uh9
qOAcnfyslMenbwsdGkUgnvOnX/soKPitSRvxFVS2uk013WK6JnY3UP8rWqLdFWEvqmMbvAoxrnxY
vb5SadaNYpuv2A3KW2JjDKhBtcheyxELN60/qb5wq4lKoRaSy9N9DqSZT+Z3wk4kNnWRd4j+0vaJ
cGSWlVgdU1mbs3i/+rQqBTYAIrOTs7JLRLjDAmI98SfwvMjQ3YG9njG2AHqUHGU4Gyfu0whVrBxX
AdVtj1yfFAGHNd4gUzs3H1Ne8F/MLvDVXrvDK5vLOT4+XwQxXgG9LcaVYSkpLeLaRztL6Py95Orc
zzZ1rWEpyb8kwJE6HzRv+l0+FOszmeqr+Zsu8P8oqmjJqxrmqCwPMJ10oV+ciQFn01I6L1YORBkW
FBsrFkdC1BYtJTt1QoppKpf+MThTWoaASPP07Om8wSB+9D0zdX2QB02xD7xD9Kycnq8+/5C4mXvV
57ZgyievRnc3zpH4JfEDeZenFFonBB2Rclw/pGfJzfPBWacJWEYjHh1LADovA/pWx6cpt0Et9uhK
l6DpftXv8vCgYdm/9cP8VxWYUpZFUHcTiImRH8zXgrgFN38fM53NE72T2LDKcW43KAZk1waudl/9
Rttg6qflxIP6htESOA0U5Fx4VT+aAOy2tYY5hhzXSZjBssc0THGu7ZJA+GQaIbhCQu4SX43pjdqN
jNKH64Pn378Bm/iERC2301lGlDEWZDogd6rcDouBETSHDpE5LvRvG//bVF0jw9Qh72SSRpFXqfzg
SITPmtsI9v+uCDpNwwo+HJnmw6RxCqCM0bO2B/oSRtj/D04bwFQh1J3CEvvKRJ9fLnMBnNc8mMVY
RnvDr9gKH8Xqbh8z69kVJBFSg48JD5ft+2BR6ZsNGZA7ViTaxo/K6HDx9b5I1ry8jE6y+q5ASofU
p9D44p8RTrX+ug4Mv3YolJSN9bBYfW6M7QjdvJCC/sBOZWw/X17YqBqf4EzS9D9K17Y1PFz8omPf
2CQZertcCXoQW3OT/cPXTQD88X5ytbuMJTXzfD1tfIWRP/FEYtesLME1VJyBsKLql+etcFIj0WU5
LommYJkOUCc4CCQyTa/ss63JqZ+OixYeOWyrKUBNuVQSjFcmM7q9ChI4Op9G28vatm8Mo+5HNXQz
7QlalS50J/a5QV5IcEvNpTO4umzOK8MBZU2YXYutYM+2h9Srf83xIo5/HljQphaOGNK7FERhZktm
Jo4sCnD9z3jDruMQ6lF4Jg2JYaN/3K2IgtYYboZbnwEP6nkhedpRompOa6KT4KGRis+fJUNG8DPC
AiqlO6TX59LKdV85qHlpRXMD1uRhhhYuUI5KjsPqS00D7VUTUkkSLuRcQ1hcvYPvgT+ipZdeTzQ9
cCcB0VymbZLhJOYCzceFbKZmNudvpKC9A/JmefdOvlJ7VE5a1XjjGg6PwTk0H4ARn2/JcGz3sdG5
XMzmfQwm3LQHuuMTARTjO4kUNisFwLSSd5VwCPd+uh6Y0/TzkPLLqnrSi5qAXq43XeYxtchdgqD4
cVRy/zirHlJrFKUk+Eryz4xdx0KJaew2GZLFtkIywa4xY0ScVcdJaH7NQL77hI/FxEhoQCEchKny
0zB8fDzAcgyhhsHF73CfxDFG/+3HtMQro8Bk+Yz0prcdrlgKP4oyZSgxmBg1Y15U1eV5k5EpeyxG
QIeMBM8Fq2makdCB9oTauCxiowfugxdIMk5d2Lg+cBzEDZPKvTZNUsIxDt1/viT1jM+CX6M7FvRh
yNNa7yOTKyCsYeD2uk+NNpr1urcElYVXjaS0orbO1l7me+Z8w3bjriz/xf6IEpSSEwIXpiQiAK71
6ut6uUlDgkafF+1Z1Y1EKi4rpajt5GXayZD8t9T27c1pXcbdkCLaU6+JdIfQZojtu0l+B3fNeWV5
a/jyc1K65SevyEoOcEIG/GsH8ckJBIki5ZcD2OhGCMqQWGlyFjInm7RT/BaN9b6rjz4XGiKjuj/G
8W6r4y9gXd0dj/BNvFAesxZof9ooJBYS3DKPLJR9AJSoRO9g+EtZbSed+xu6KIrFwpmM2FA8bKDl
wP3HJkqJFS4WeRqOPX04XtHKTY1d22c+WbSdGtKOOwAB4jPt/Xbbv8AWrgqGKkSU76kuOYH4/az2
/VXISMUk3fBQ+qtIMJATW4uWAfdS0RkOQo0L6/T/oQqhFF/62SeCTxqZviibXhpIZOhlv7AIQ2TD
fvkKwE9JfoL0Knduaxm8G2X/XcWUBkBeztc7BmNzOH1O4FcOhhFHpXnTUVWwV16hliq7ehUflUyI
7onbLIA9jYSzNTS7CjhIqqK6B639UJL+KSXLBJ4JIlnnlGXFGKDF/7MogNNYZ5hlUeLfionFTL/b
Homi4OcU9WjsQNYAV4MqEJCZNvhLDEop2vpIP0XJaZFnDnp7MSADIdE+sxl/7drwDiNJ7DLqcA/8
R7yIpYkJjYnvQD2FFzEDPwQvWGIqo5sac9jRkdMObXmvxDoiuksk+MgRyAd4H0Udb5bAwyj2yPEA
rk42kYDSqaHDDHrSpJb62pzytTGjzHYAngOqhoj7iMNOI0iVaO3Une9mT24RjUJS4ZjtvFZUTl3K
iM6LQZK6MxVaizxpnxOQKeJlwR9RAUZWwweLQ3YJirWZB4Uk7X21Vp2sprblewEhgb1EdD9+2mFf
OhPoVtQ42HqcDFWM9oGCsMlw3o0Q37BQYTBmHlYHJ/LC3KR5IEnKKrLDEuJAO+mFW1Ot56PrWICW
S6pyoQCTqbFgmpVOt3UevkGR1GXrAqHf2zo7py4kpVOsq+dyWR8J0PFDHduOdxZFGOb+VENX8yhK
DtdoMeAGA+iE07LkEKbX87HmhkNU2+KTG4xoXCVM9b6dIv5NtkKKLx/AiG20dbbrlHd5iGFTsSjp
9OU9gaNZ7iXUGgB7omJe2+S8Gl9MpOxg7iQU/PJesFtlGL0jnXyqOhQQw877A6Qm2LCALhwhWQR4
6lBesiABlbO8v2O1YQGTXVSSN/Ijov9pgLgA0+2iF8ZfuqzL4JA+qXohobG1L+eqaBI1jn18mK8D
Q4gh9olmqv+bsWqJzUxfYNjJDX66m/6rFEoPWed1tSkS4INk8AH2WLj/ii2l39YFCtXrAUkfacm5
+l/ZP4A9sNWUOZ16ZGcwOkZzzufvkv/8vfPhGxJCY8dQWDAqYqm4vXPntViJiVjWQaAO7EeeqDs1
ouNHGgyY3F1JNjPKnpo5rt7OwyJUpghWcTTFTyf5eQKJc12lhdBxAYOAR03lXiKh+lLX4g8Z7NFu
NtrUeBhy6q73rziywQBSvQA71bohpPjwzsSabPcFVf/cGjnvQYh/AB6VPZQbYZ+G6EjgYZmmWKLS
cseh+Du7qqV7wP9vdkbYxGZWDGs5tXpXOAh2TJvgMXvMLYOGsOgxlWRnzh6Po5+K0i2LEpGro3jg
4L+kmJLZrV6e4ouCj8Aqq6lfbAUHlSDZsvPzvnaZ/KavByQE5+uCYh0murilRZ9idgbpGkZ3jaMY
g9ukyASbZGO1mrZvujCgMKTgY+LlabZwH0NpqwFIxeMqYwCY1qYS4PZx7YaWRSMzhN87g1fEWpFI
kpd56/5/W6rrezQRqMG7NUZbCuoserglvTB2hA8HqG50OHs82kEQASe4MzqipTaKDm6F2Z45Kajo
cuxoW66UIeqAnh+lfpaHN6jNSRYVaMXffWzdAp9Jg2TJ/vDb76Sb8MJ8QCmGvAmrXcTMnEfuGC6w
8nqk9wef4YZz+iLek+dp2WdjGYF3KmzQCXDZDI81OtgjFJ62vU3La0nFAd0kLFpeEr4xbbkpZWvQ
Y34UGZPxpGkALwia1VsgKTdtg9rUcidDmxJOFTskqc29OSl2OVQhABDsvxfsZObl5uGACBQoWn3l
7oHyNHEueCU+LGq+1ITdEz073jz1lUjKIAWfY4gocpyTZaFz9oMdaKTBgd632KyVYxuzuMDrp45M
TeBmQjSGzvYNv/Ja20GiEZ/oA3F6w+dD6VRi4gJJljAwf9bXcJNFv10/B40io0ywwIO6GtZ35PmY
vmFbTY2nYce3hjeqz1tnZvMG1Dk3nl4rMppiOxq3pV42Yb7582GWkLrnMsAl0B95+lN7EtxxOmOC
nz2HuG6oBXQKQPJ+lLoyUrGA5H3BmEMBjWEHSZEDBhsUmx0DQnz+NBUy/1RaOT0WQ368PKukTn8s
vyYIh4QjdjFtljWkBKLUy5N8f9QvAjKx2kwpSD7a/38qHLb3u8su7+ltah2KcEOsBrgr4kdzBvJp
rk7VvuLoJkC/VAZrCvfzRxCPJFyXN186f+JeBdUMZ9rO5NwS68HSwBaFRhSAC+nXcH5Xx/y0EZTZ
CdD1W7NbbOP198fQBlY6d7hVN/AhDN9ia+Iw24NN9ja43VgezSQvOmq8AAXK3sVEp+GiVxdpPysY
1w1eBDdz8+Jxzii3YBCJ4vT7p7fBrpRnbuB2XPyuenVbl2SuLiDLMP/4Rc/pHRHf/OQTvHwfiWRF
0DNJtVlUzpWcm0u+vOXRaE1qZonKMnKzCpPmiPXL/QyvQByGquduQnjcK8DnaQBpk0kv4g5Ys+4W
12F0n6P0HzRTd5Zwshq5piwtBMvy7uItzuBo7POGQSZe12NAM+Lbl9/H6LWib/RniLjOcdBZfuc8
Zh6GWScnANLg3qBLJB8IoFOGY5XHadIwM4Btdn64PfPH0regJXdRihL6EdM4g4LQQsOAUKEHS7fS
gmMHanmBcN5FbOWsVmfaAQUq2EwlWQi8uL/tSyIm+a4wDKoR/GgWXBaS3ulk0B58KvV+meC/xA3X
sUyU+qPOpKadC3ETMumpJbMljAb11R+20hMkotmq20hZyuYbCFG20RqjYVcTOOung6pCpXxsaGDC
6pg98+2VBT0jEjCqNZAMAFp+JJjsX8B2GZ2s6ti68qHMmaPCDkt0VzNQCg17JEn049C7T1vQ1KTl
UVo//qidgvsduQw7lFHLC+cTSWv4X7CcJIfmVkqnp5tz3azAJ+fz4xvcOASiA7ZY2c5F+9pXlg1l
X/MuLCL7DEIqpeevfLLcmf72MLZuAF6gyQALstdu5Kr3tpsXE+J+eviW3Juk7ObryR6EaUHJkK0M
ET86pAySc4Y8lCaUnbafkkx3kfNSRpJWWu9R9QKp24uXsyBFlOwUNZdXhHti8LSBLjRT2jNsOsPl
sDhWvB1DzpXVhvBt9l1rnaySaSYN9vM8qOsmm5Cq3zP3cDraLtNpvl/eRtaSi/1pj472biAq3Hqn
a24Nkrf4IAX9DtSVpVzBOePKGBEvT60nPKvPNrzCC1vOUnx8zXOKzsG0XpRoGNNjpcodeaZ6QXal
rpJ/LnodDqLndcmoAw0kl7n76JMML/GtlY70RAZc2cZhNrrG6AhDaTpsz6VFfu6FREN+/+EdAEhY
2ThMPm5D625lDDmCbe1pkyJLP728LRGISlPNYSxHtKp8GT0MY3seikXKF1LrV1EgWK/LQTmnwSAq
E59vVXAXBu/MfTmWnyij/aXF5yzqslvE7z6aOWB3A7vpR4MCOeWq6DiZIBn8ztVXlYoamcyzVZMG
RDXMOAGif2IkkoTAstp504gYZOzeMjXaQS6ozD5/TdbxuyjhmOniEGNZ/DCWYbo4fjh7cmaLSLy9
qCTyTgbwjup7cety+c9Kpdp+p56OmoxzWSqzEF6/cl84ne0YAmRan5TuHxGQtpx2tDnC2nWLHHbO
oO39LqQoCe5Y6K4GeZEZp2txX9yNtAE6+wgvs76MUZnxZbO+ykyvCS5dtCwvqIGffkE92ug7QYp7
Biqgad5TMik24UEkxmKBeGxwQAg4v4/gOH567n2PklsiOBvR09pMT9EDlib3zWhKcpg7ZWBVQsQX
mhkVg99pF6E3Qs5c19qLvB71BwoGu6EhsZwVVqPFM4D+48zjFwkLBTAQzvIcGTRPukIfKDoRqDT1
JfDArHgYae/uSVMY8aKg3hLRqT50GmqAiR+S9H2KH+XwnxfmX7MQwK9bR2ElTyHfPG+TnwiwN2V2
V3j+2GZIwQ0V08Bh3iqfZ0wn9mZWs4Zk44tNslKsz1IeHkwBNKYSj7HY0avm85dLVpCpnsqby6dl
O4v90wh1BEZ5q/qGduepIV/TKrh4a2Z5YqXF+JceqrrjWuuolZY/lABBBbd+VMV4OyW9ZQhkjKM0
BUh3Zrie+CXL+P/qCXdiub+9QbC0OYxPuYMq84Dv29wYsqi9e4FmZtjuwqC9ALYCIb7JTzPvB/5Y
Q09RQFHlWTuO7f48Rysd84sGFeViUutsvrN6LtB818RZHNeHaK9XTU8qpxeplZpxML4+du1OgXyt
L60xTKBwOWM5631tluOWMWpLCedrSm6CspY2k0tragIGDGvEjwi5xMYKstM195HffUH6Jq4SHtZy
mlkayF9u/9t0gBUF/sZUtr/KKzXMuzV35wDKh7PM1SApARmbm5YLMu4B/240MeXHyOSgx6/qkYRr
ZaBZIpspWMx4mc1yHutfXgDROBIQTgjuJS/2G0JEWl6WY1MHJc8mvVTvLbd5ESnaog5xOxXfNW3Y
hTgFtYaw0k0/DmE/C45Wpdcv4N5IYN/iMhzAuapiGHv19EPMVmvQriKIvhCWyHClpAepSdhezRLS
aMozLVRE+EjhZyhUCAKHMn8NbAb54X8K3yVPIDsDeIFMqTyfsgLyTZcPSDSOUpHplIifJQLlLlBt
88u1AWZi3zPH9L9X9uLe3qUdQnmNZlHZ92aj3aNFVKK36i894cnRpJkxX+p4EWowwBKC/Bg5W29N
BSqlxdzhWkEPmOyiTxBU2+fejkobZNjoSqRSbPE2B8ybMEG3wqPFrz8lArhCCCVYjfus+wFXTWYJ
klC9qaneYheR+ZTFkuEEvgYUXUMtLFcoYyzUpkBiwDpp4GduDm+Wz4mUg33WWkaj0qj28Spm7SGm
1VowSBlFxnfCJXgjWUY8lOqY/hAqUbff/c6XQbGO9OCpejWyad7dLlTh+taMvNVvRScSu6G1mGEv
SR4xod/E7UuzI5TcaUp/le0wL+whhYjkK04nswnTItlM0Hjre26l5fui4IkxhCC1qqDhdJAD0mCO
5Ozu0AcWw4W+F9/E9mqgCmQpTSvz72F208hpi666DOkvyj0SxNcHjFe5g8ETi/b3daxcw356NLgA
+1AN4zD0LvD4OmVR7rzLKU4RRyKUyP38pNd4U2UiRvf2QGrwKOglHpc/eyWVe2k3n8f2dpbnSdhB
AsbmEz2HnCYsbYbYX7Rza60Yx6GvIVY2hMeVLczsBzdQipG5CvS7RAT93oc3VIlcPPQ980GDuMXz
q2pi287w35sypM+6NUoE2HOwWjutenHc35u0Vo/0mLXmaS0jbJWQH0a74Epbpc12tp/LqVvMBCY4
hf/7qN3H7Up4BmzvmZkc6uxGUARGjDOpTEKLz2ywS5WSggI3tAuH6PlYoFzeBotPlieUMMEFoZek
HZGvsoeFeiqEFDqxL5oltruoYK5kGI4HN4+JmUeWJRbhXlyoFEAsusxdAv4v+HAL4BD7CjkraanZ
G7HGrFblBw1AHsQFrzqgfjMAOiVbpjfM74NXTCtk/WorKq8cQUgr+RK89GotCtCVXVtIi+jj+0SS
V0I6C74i52ppdBezFbZUmuOXK3UWV1jR5rMTFwBFUmwrA0emMjKWFA8KfZaMKomI6wzIibG7F1yT
WU3jtClOWDQbvWDiS2BmzZHIOVCFlZunqTgHzg5kD76F+zbO9qPGJmy87IvZnsUkVbG5c0zhiZZX
D8KDX3sse0uaTvD6OuZKe/uT0sNFoG1I4EskLJdhp9f5zeqXCSYfcKHVnRy4rOpluK/LH4VA0DEh
GWpsbsU3a2R5WqpKqkSUFj8nXM/5EkVkvFpTSUA0J89ZNPtdIg4cToeCYkjReW4B1wPcjVAbn0RR
cuKbYyshUCujY69qsq/pTaRwSAg/jalu3xw6tY9cQp/ikFXF+4jAIukIxaolrSEcva7RW6GPin+B
ngjdG0wtcdA1+5Brid8SbQJhaNupelvd5ilEspjr19fnPUjcDqtIPSfZw6WoqVLBhs/mh9lIekOo
q2uZrwlAbaebUipM+yzShpmBkziLCYmCpNk3Szy0goGTmeqXVd+5G/GjiDY6wTQ5sQhfYlgg6t4N
39gfQPpJVctCIYNRB3Q43j0WJk26QuYN4jSNOh1lwa3A29hXO2In0tnZNeFNRCxjgGzkhnNVlQZC
vtsT2cx0K5q/enkUWa/y+mipNfYjK9JCY1YlPz2nl/phUfxTD6UttN1euzIAOOqBa8LR9miUXECB
c82zzZfBWEssyyWI8t8C/XQm/elxgCtPxNfeU/8F5lUtRlmqWPQwf9Jd3P+Cf/gbhf5KXwdlF5Vj
5SELx1SluvHHpeNq3gmw2zI6VXIggLdsu5ylZlsHrO2jPTkz5mthtt9xz8E0mNH4VJjAOv85IwMh
DaRgoyHCS5VRjlgTjLN5nOHKBXm8mz1uDEO2nXb+2KOBc9Mvqn/GcAZh2mlK8Mus15Vsu+YyG4+m
2fyipf3/Tym33nf+Wwo4g0/CR4n04+vt1Wvt9+EH+1BZR/7bFu93PUv+aP+OXMNiExvkJn01s/qs
NzB8ecgd5MRmd4NJFnD4vvthAQFfHIOS/BM4i//gLqHMzoEg1xl3rgiYrCW1qqff4+8ixV1qpnlt
h36l0tW6r/jKvZxiTZcfMNfb4S/f1Fjsnw5TbQqFHdAXchZbxCa43a1ZwM8khWIcgc8Kmod0G5c3
DOs6LEQ/a+tQPTJJ98mSex3NtRAmwdk/eYijziepqeIbT06fuVYFrWjPxdaDWjrtM7UVjMczYpyQ
KwkDM5/bqQGcO+ypoYdfp130RpPCQ6gdhfKPtCwy0iDsmm5ZGpycrGq/5lMSwR42KRsqRrV9B/mn
VwuEIuzPl/CbWmKhtMmo9qppjgDQklWsW+g9XP326jS2EfoZB+otyYgEED8kaEXQu2UUOQb1/mTu
q63U/PCkdtPozzLh+rDY0zIPsc86YDvx7YXTq8ZK1sdiVoK5GoTXcFU8YTMWeWiBp574eiR3PSgL
BSQQJ4wx80x8Z1z3h9qrEYbwcCxeLLrPveNXS/NWPbBQkRfzncprx1YK4sU/VygTJvSZaN3XzkC+
NFmYhk5CjUT6/jYxeQD7kFCUQr2Ijp+akRbQ4IygxaYW9Y5sQD2xXxvEz8HqWCseeePdWmavYTUr
A2Cn7DJjon5NY5pkhSEwKTqPwoGcoF2iCL2YCKRhTqsrQOS2lu/Ekr76hiCqHi2/ZP9ncxyCI+0O
GPfFmhHWpmWBCpDIyDRhrYExDotB/L0nQXzyYnk31oce7+DqSQiEURsMwyU7Mtd65BUXNq9sCnjy
Vx5ggXYZaaCccWICcbBZAVGTCtJivHeCzLj1ZsLhpoOxE6+c1r6Fc8ue2qKkiNotw/VTYqLdCTGp
rMl7KIoPWlYKQpv4nhuxzPXjsHbS7i/pBOIcisuOsdFqZWnPShbi5r3Or9sKlfkzFgYkwdy++NPW
QGP6m9CjMyK3fcGlWs2THw9IR1IqHBo17CWMkYQhhC6TESVOTsRGZgecf1fpb5+CgSjeqHp47XAY
y2DYDzJ6S/bbbqOZBCknWZeIqXObZCnAqc24/9gdtcMN36G01Oom5judLCerwhxpnYV7GYBpAerj
YblIJyZuPEc2tcu25aNtLHt78KWNEEJJ84dkMAMZB+uKhDiqurdWNE2KuabfJGKqvSwnN16sDGa6
1+GrHqcb2xGrCk/qGeI6eovgUtH9BD2EyurXyfTtAsyUjoVWOuCnAsLmz4TTlGNxODElLZWtFIOS
a/359OgFKIAjU5ETFX82oNHkZd26wWPF8UAI8Bd+XWP1MZtXuyvYI1pf0Y05DtW6XQ+RVTw84OpL
2Z5XDk6jtQGVbaGcjnqfnZYpX+Yx52rduk7gBlyt0RGeOGE8hUATJDTNimX1rz61kS2bT2Z8VHrm
YRRgwYr3LOP6LiGxwaKUWwzrsajkiu4RmRwucIkMP629sqJXQN3RzOQlrg+FsaidxWgqGB08VZjx
mLFBhjtlNsavZPa2y3GW4kS8WEEiNXqSTMPx2Zuool9Ecg/lnFSYinmfxPDfbiqNgca56II6dYOX
5IuGCl+I08sXZ7mvKACqJnj6tTbN7VQwIAOiEE8PAbKNXwycz8HVybUDBM75bIKre7ZMZr8Z/JHJ
c1QrT/Q4EK08AzeFIvL64VGi9YPHSq9ZGKxJfJxEvLW4ROyXXPEPxvdLWnRtf2Y5mCvYCOuf+ast
qliMCEDlVKFP60o7DVznWLS+wdMSlAb9qRELoxfqpWNkn3qWa3LxDXPaE2iAYjrwpOp7yRV59gXB
VolvNtBGFkH/iKFanfUzdBWcnkvjPk3ilIdVDNp+g60iT+/qC8+u3yxVVCz0HeAeFe2ZgndPjSdq
1V1lXyjQDAzOhTgGszf/bpz8r5TfEG5q2qi/dAB3aDB1v+GNX5u02BNFAav5TwW6u8DM/UsbRZKB
IaYfX3sj+KAgHdgoCB7C/kfzI3DhPldd9OnAaq16jTK9mk4s7+uuDhal4UC+ZSPUtYJL289kPPuc
X7OFIrJAjJMFMDkKtJcx3Skzo3YFXZ+tsu8M2gxztC7PLgB/g4tJJNkF/pyN5DxIgd+HZ+qhmKwR
sZTla2C/zyw/Iiem8T9u0FXGAqKPbuRKF/xGhIDM1bOgoSworsKbFKT/4GQui3GS1sS38LdgHp1Z
tt5WvAkLoADMVaCqpzpFE+jxQvgCTzQfCK8J16tKBzymozC9mWcI3o0o6vpszDe4T4Vp+tyRqyaP
JTRg7Fj9k+nOZeTYp6S7lHfPcu328544JBEv7cIEecglTvv8wGkRlluWnxbVnmHJoHXrniw2SPlC
K4BHIAWfz8fiTRbDlxK0MMvzgvY8tN6Of0gmAXQ8yEeeZA4UOYIu1Og1FF7RjKuhvNdrYorEWdXK
aURo4BW/JDPl5pjeWxSGmUDCsEUbpwPjn68jeGvbLCswMU9a9IXv9z757iUBz5M+MDCivKuNACgm
i9fsDglzNu854wx9EjgIakgjmSvM0zlWKP0KwEf1aW+J/hl5veKdSIZAbrV3r46j095JF2ksDLC1
8HmfZtNw1uOodpeJvwZADXPHFCoaHskSaHdwWZqC/C5pQN8h5Fhw1rYHVg3uQj3oCbRcJYlyx16y
c0WxPq3GehIpMt0AkPCC1OYdFEsH/tYlXMULzkRIjVs3RypV4UiLhDSKBj+i+3YvK83JsYyW6SHQ
JQ9F2rr5sC59GiUEYq6PqlHFAq5v1qBMjnKpBSBy5EA2QiIo0FvlBHsyjph2QkFuH7RWEvoFel3Q
/fxj7XQWqasftYgiaYJ6bZNXvMCxEiEkJS9N2AetGd5brp0xJZxs+lxeDEq2jLeUbn1ADLbV0wNR
VhGInIjn1Ea+43gCOyVYgS4A+TP9TVUyOEzZYqT+HqlybpJXDOVj2nHjGBiVaE4Q7WbvbCh/FFa9
mfVqTvPt2UBffpEHOUPxr+GspKgmkQO+/xPgfRfpmDCUdA1g8qEHdgAzF6gZxWeBXxHjdSUmUNPt
gE4oT3SZqGhYE03+csH0deLvJbTLRCs5O1ubmelrhTlzIkqqN8M6MYJl8mEdCfyhK4K7deJi1FNb
F7Zn7QeaJID8MnohErrjzjs7YeKiPO8FMQ2VdtfcNaBiethkviXYhZrReKeEgcfhUXvULvrOxbPD
KiYRezUa9nB6pCHaoT1DqxQY4rku6A0hSiJxtavXZ/j9+1SAn2LEaDXrJkXheIaekgHg6yyUfMLY
m/PtL8cZIHSWxNRfzf60gKz/Y8T18GnD8Rmg+Oh1N/WZSxMmK5Kh3rWnEeNaRo6IiBhvPlR0Tryo
2VKa/g/IyhTxglwxprTVlOKyVD3c91Rg6DJ1nJBDOCAEbF15Hre8SBeATQRn7BUoeWd4uqxaQWGS
edURuHtzkVRyAJId+/hKBwMezc70gcByX/4Ls1yApQMBSZtIOpd5S/r2pigZ8SbgYy7RlaX2iFxZ
Ym9fbq9oDQlQzg8tcEqQRvwbz/BoCxoXZwnsoEjtRmeHbcxJ+cjvRSb4XBVdceYEUF7ux8jiNuvI
stB0mg3+H7XiFa0AKsNAkXtlc08ydysL/t7naF89dtNaYlUik10s8pdmN0XECd9GDlcLl98QOi1L
/klY4GZQR7x+P5o8+vMxENGI3cCAfxeXv3kf/SGopXA+jG5B/QiNIcPJ8Zpg3vtRZDiey9YWRsDp
l37u65ip/zEEHuGCvUJ5UVBhmUk6LER7riheRyf+tlqdjSz6Kf/pLvx6MDlWCvKKANDSXUgP2CsB
hucahS7/hFOHpBH1AKvQTLR/60dtfAVPfWtg4i4IueKWI4Km5CISOXQwM9pyUx9keV1upHv8Rpqy
TbGGhi7NAP0BOMPwnri5jswIyAiG9gkGThJQTNPpFU1HTAEGrLoXq3M91CRQogdTjIMtI5poqx+w
wmlbbq9SwaaZh/MFn++9izB8EuPU8uzHgaDW5US6g1/gyTnlT7FUtxxF15CMtrZTsf0pQLKB5Iqw
AJgx4jECqdpNbPGCDrjg39eXfjmo5JbEomnXGFU6gnIjkQ1joPga7Cdv1pT/YXRzGD6txJ7VmOz0
KK28fuGnIQaCiVG42vdvP0QFjowRE66Xnum4OcLws+y+SRDAKmlsu41tBfxMfERm/58MDBVXVPW/
WcAKSOZCEfRf49GXKPm8TaTDFBTs6tuTv2L1ixyyF2pIHsUPKKheO5T7rekG6Xcag3hbdFH2tqac
8d+gNSjpB01Bu28M2m7CHJ4HaCozYwCTrasMwdXgVGmT7icn5D2tQ+YR1IHYdao+Co0MJGdK/5QZ
reNPam2MJCC1dSMDQqCrQIEmklhGqO7hAN283tgbQfcMxpdJqBQwvXekyBGfSypx6MLzJC+3go+v
XKh74F8LjoBAmCfCglcl9GnGtrTYhIOasxxCXCCqGA/lMte3yvAqgZ8HHg2bGdeZYByomiE5IcLi
bJ1A4fUKx6l6js1BMHZml7aogZPyklvHbiWkfwXqhmB7haF7YDkFAgGZzOogpbWuLEMGIbNDkRbj
FcxE7CoezaaDuLFJXQYySKH2Dxr5pNcadV+axhTJ7C8yn3k5/DbFyur6tUqJTrBlWCWlR+tpYudV
3GElJMVH177S5kCpd9cIzM3V+KPJyXNZImLDRdN1wT7mbO4TJeRs0OKxZo+jHyxXglm5vUXdiLGa
hMWHnR9PasS/dI22n2ae/0xTcFsoHUoOppgy3YkMIQ8nfrdKc2WPWzD7kLu9nAfQ6f7vCiFZn/0h
Y2jxY82/soaMK0VYoLfS0EHXRF4Oh6J+GUx1b+KqxKkv1zDYWq16q+EN2tNaxex9XcnIva+iHMFt
1JMI6WCnZCI8d8t6ciC5Q96CdFIwcdpFAOGaduDwhD+6riZqf6mPeVTL7IH70/9jWRk2nqLD4YSE
qdZI7FjnditSQTv439C6Oh/5gANFLzXNdy+GX9EpaWrw4FXCYYGiG2Rgxzj/WM+TkQZuIjq/ar7U
hie2zEUebzoTnmaQDzns+2d4Iq9akMmpeh9JRJ0U2Kmw2TgAcY2gsFLXcuo/WhUwRtQVUUIHVCeD
EdIB8V19AkC7iQvFnKCrCpkJETYSCcxvQ2VhhIE5guGCSdGlZv0y113v1wcRP+62hiNW1Chrc7Dq
4Dn3/QK6RJ1/h6IfQiYtg16raqZL97uRe0Ckk2LEacFr78iht1X7pgKb14odyzXBe2cGpt6LDofg
sqjMQ0f7DfSTbUd2kU311VDPF33s1VKtR2TtaRILMn7WY6PjsHGi4Lqe2BXjHbUw7PwLHyuzBkZ+
Kl1AGLb5b8lYG4K5uaRiP2Ad5akJsy/STE/4oiGPa3R3ore4tFzu8ak+odsgbDCAiqoiYw9nWbnD
QkZFj6lB13rjjXXh67BenWovrPWrPenkw4NSSL9uizyKwsP/HbZc7LXin9pgrMkSGDHkRyq5JIfX
Z4v/D5NMZCWbhzn0tXDCHawRESTegumswplI6QWUr+v1D0eaD7eyhZVpgTQUwUcb14gQoHVAv5/f
gdTPbQWFA6R/jH5z1MEvkWo1EeloXDEsbeFiQBtALYq2MHTnVaBjzJm5Isvm6Qse1Wu89d+o41ky
p/x+nl7xwOxTbP6AqSpz7CM9x8u9396uROK6p35KQDa6DuJGCMCddjxqstLib6uOzj8+2VYIkNxo
sLLHwJD0JyIedwdj3UcdgmRVbyXJEKhJnmdMbSCoCCvZ9k+h7bEUX58l9rC259zinTRfCpaNB617
8X+QrJ8dRhkbs3pJqOJHlFVZjCg8LajDK8p3kAwG1EfiNgaOdqek9UvB+mjIgUPrjHIWOlTZ8ID+
c70+I7fWWki2oDYnBytSig+1CrVekCzMMf+vufyZL6/wMuxf4OF/9MTq4VDcQy9LiuMcdKCY19cg
yG2rWKcapNmLgtsnbLqz0wM+wHBTkAqeXyR1c/nVFMTIzwqWxoyW+bXtcSiYVJdplZp/w7+ZoKIR
vkcQkIAMo2J982eDfntUt+6ZZJ1k/PNRttGG16M8P5CBmYqERD9B0yh7TAJLN4M/O6J5K+wjuMPH
krWbcvxdWiirGaTyI83ungz4u2pWkcQnQ+bARc7+zGAWZJvmoLG2XGDrrhlB1PaTU+Orsywukt0e
ZGGefacVCHdwKsVLBD3Giys/W5E43RZIzTSvyl89OghWPhIKQX6EgMa/asHrSTZJnreHC1SdtrOw
3cQiiILTg1uzVfdXjJDJXHtMQuqhWLW3TVm/3z4NOPMeSM4ZP8J5zmoXDIXgwAcAeX77tm3LGrAl
SMWpgfBS7Co5UxfwFV5P2PKhPucrbf6qfSt9Jftd9HdVoBg67U9aWTDmVTBvN+KgI4dj8knx3qYm
E9VDp3Us6mP+BbxUedv9istcX+ZBVGiF7g+lqGKU9+sUmG9lwy3dfK2//1xyW2FAe+1/RPaUk4wn
JODM9daUpt3qjnQnVKlc01Dr4LmTZFCkbxROon5lhBD7qEdl0m8KxDydvJY8apLaaJBy35yJNJvs
U7P99K9DVNX65SlRglrvDWD38axME1RVelX3VB24CaMB/WWKB1lQ/9vD9pWrXWHBCYHCyySTIXAr
RHOT2ps8LecCQ3+S6IRrxdmBAiFu2MfrcyC0+5hKu490DfrnROKOCdpQgeohFDCqLYmAMChFso79
Hf6rSMEeLSE5JizNQTwvsHjzNs70XEZmRXzA5qip3iFcMf8TigBMm94aGjGsZx4DuqB3cpGkQG5u
xenS1uN5q3Rr0yrIPtfGqg7pGRmfn+sK+/dMolYTteDFefLce3B8A/ImaOPfnIqkDObabI4BWTlp
QZer8feM8Rm6iz+XVCHveQAoJjEGToZAQYK4sCwXrZ7S/ymM8MfUD8AaFlifesffiUTihdMfOz6Y
ikZADmEpMudH9jpXkHYzHG2p7pzYYgAtBEnnia0l1UJ84bZrGdOAZOR3Q3bimQvhh7qLuYHjkF8r
BQsiU8Ep/+YepF19SDdqAefs53YleIjlYUJr+1NtAI/Z4Rrq+flWFiLRqK6rqSBC9pb/oKhp+eXu
7GZxL1lTPSffAZjbaHD1JW1NX1JtgLRgf28vaBeDtf1fo4POF8yDacLncRqacsUcnnOVFKc5GxJM
kMyQKdbQfb0SEB8WftpiDCTGQFnU5sNSZiJGRxmWcPC71pxoLymgSQyPjCKh2w1u5rqNestzzqPp
T5jY+pOlmuTSebqsCWrg4vvHy31hu/nOD27VH3f2nQLxvGH+m16Ye5kO+9Mtwhl7ltHt4ZPe8R47
WkYS3Oyvj4lS0SJCIM6mEjspt7h+4HnC5ePeu63OVYOmJSloF0ysjc19YVZRcouhTBDPmjDJk3Ud
HHmOuPwegJOmdVfVmOZUHEwHbvxG/63Sb2/ArHa2PozOiOQ/WsWmr9ss6c6dgQ2V0F6bc9a8kifm
y094cv72dKLlkanNr1k03zCvfRiEQmuDKwI5dsCipQz4HfjmUEtR7MCB8diAP1BBVHWCKvgNgac7
q9FjBKrico87Penqm6fQo+KNOynw4yvq6PmVJwWpP4UfwItgi722TDRFqNDGeDYXWGTm2voJnZxH
cFVNITTICGTv/8cCtQn8jjUgkEa727xaKcRt6vE7vRU6enm9dU086KjT6nARCy1mQdwFNssImpZG
T17dMLaGyqHYzo2VEOydJk36COZOvtJ4/8HkGKprgcVvl/+HpCE2Bw4nkmPdex2ujifBnbfHOvgD
mviBi6k2LJCUgjaGh1nYEy6qM7J2xT4NXdCLIJVpwY/9Ant2kWPykT9JI7ADAhC3+K4TxgcT9jZ0
YWSFLLtLk+HND6/30HyzInixlWlKIGxGOCepZwgale41LxYJojSEo4SR3DLMaSEyCaQfXO/vaABm
/eNQr5KgJ2wlYm9v+m1tcuYIg8wTPHwtCkuaXMF3Umn8oKIZFRN31vyzSmT0YHrNDR64L0PuBqRW
L0rOOLmQ8yt6NcCVEYd/VLAhyfoWA64X8P25onU/2uwKiSk3vuS0+PgJl6S92ERZaQEwB94kAUfh
Ojg5pFgFzsbf8jl/CSRUekdLqPzPOSPLY7etVkHGmdz0vDc+Tma71nJ6lk0ZbYbizgI9eH0ha0TF
Pssyr5B4p/aA6J2t1d771PAk8LouGjtg90N/bTf3mnRP3PZ89IkvC3CJ6nseXYCscaQCPZ+H38+4
o0+3tlD6mvgOCAcbNzgktt/1WYgzW/Jlgbnwa4QCQIdH7FuukZKAlFz1WHrTT73jpI1GCKs1u3hi
DoyXmjNuwhlpcrnJ/21QPR4RlywvZ7IwbI5/6JHhIjHV+n8K7ag0nLsU+RbqnUOOULk4GclPUxvV
BvCPW6TLC0jr31I6sL/x7wKZkhmLIdnz4u27sGjBfdB5yhTJQUSqwMciK6DN+vd4ROrju46HX2gn
zX3qvMiqiVLpkT9vaPchYeBk5Dc5xbBBqK0wwpgZxa9LNf640TVogQjNfUPtbRH3Gc4kFS9fI5nY
L54OlSjOFdU/l1UZEQGTejskuSVbz27Hs9O7lMPnYHeuT2YjkjgCxlbB0Dqn2pCtbzMvN8J81psI
6z1avyF7zzx+gDqZm1eFyw/7gOwVc0qefsAcnm03FjBHCVb8/69ulV7bKkwoIqBesfYL7ajCsNgm
E43OsWryuXdlGfAWld66BeqyG2h5f2MrR0ijdhoOanZAyx1U+TS0JrslYoMFjZzHdjZqQXGAv3Mp
r+3cPvA3wPYGWbol8UkTdWLBi2Bo/1LFJxH1oMqEcgol7yFXF0/vFUcaR5I7pMACG8/vQchKp54q
rOlOzWLS+KwJ3T62mMfXRs6FY+NgNZAAjW4S1ewVUKUeKIH7t7AThcgZEa73QNAs63cD8RYYia4Z
Bq4MBMgXoral6W772cCnhmtq/pexGnzXt9JycCybg96RqwkrdOxh801wsP5iuN2pFM+OUQYL35jy
oO2Uns/j8WBIURIiO7arWvGKA9dfzeT7WhexRLoQqC231JTWaxwXJTfQ5E0qgcit+vJcDWrES7T+
WyKqSP7rzAnzBe2qXktz7dQQUxv52z/qORKPdcvlRiWvQF9dOCG2JCwdFRcDQ6eR28QLe/dij6TA
VmDDZwKrXbgseaGGbBHsQlhp0K3qcKpsJs4OhZy/awvXs+DKMO1TC+ntz+zqkY3yFI5t8b4EBwVd
yECMGhJVPzCbTqNjktQgsF5iP1g+qhHvghP4lSFO2quwhG6d4wgE2BCNSkEY5zAY1IGmXUTIrdwT
UzqeRAXBUdM5PmzHRyX/4TSBBCuEVdLD75v5ugL5+/fPPJrCHBXmZIp7jqY4ntOxRtqG2yZxppEg
7RTXeQekj2u3H9N1B0xRHPV6mWKE/6JPLOSRjyNnRVdQMoPlWaJKYBuM770P95Sd9qAewW62tFUH
VhXRPl9LEQbnpbDw5wjAIQodpPBNvT3q2H3uaQjvh2i8hrCYhUwUJq9MmXpaTUDrIrfvAifll9q5
VFDN+2dyi8tnqkoGXDRxvPGp4LWhZCNxJL4cFbORNa8XIdfkXEurnY0olgMWCnNu00XdlJMJoWzs
+GEaoaqkp+Aec603EGRp9I2BjUq0PM5ECOT+YoA9dwws139UNPr0MStNAVuIk0ecMSK7X6NQBRRk
AxDD279YzZwW36RgGjSSWUI3+GgPmQqX1/WUPKOj3Dp+cMowyRASMr8YLD2Cfh6axAEWvZbF60Pp
+sBwXiYqePrKufYO1F5ybyWMZfTg4ia8VmAn5/G85FRhq8hEzAc1E58V8cy538FZD7wiMB7LimHw
61OdTRZwNGaCHTxcmcH+RBePJAUl7c9B4DtiyzMFoG0NLYWGKtbCdPsMyT4AB1Pv8RhIWM7sYWqx
RZZ25jMj0T/mbgHtRe+8Pi5zqAqOIPx2g5MBRH7MYYaiKoxVKyhZU6YstmZZnrEwWxZpTAxthb4x
Ejjr+qZFcL7k/1yPQx01HvlNDsuMKSdsdYBWqkL/itXddAEWaQjzl9FT9UJDtwL5DmeKZLbyw0Aa
yI42h7K/vTTW1A/HFjhP58S1xcLq0SMsKSr88pC1CMQu3igCssARb1w3OSRhzI9XLiRF2cnKHgNn
rvpn5Amt4Tx/mZVH46L+rQr/q7TzClPFAzWL5BLukDA/8wyA4u6GO+TD3hqPt1KeqrgVANf12I3S
akO/HkCl6KWAezJhj+yH1xfMCRyHBNIDqZxcQnhy3gAshZhFu9ymeAu6pEEUG6tBH+zFhE+ZAeB9
584V3jcosCnKk+AiqEdfLS9OvUsJbqhTMuCN9YVX5XJ2q4qyOBIpER3inT0pfLFbAbvzANpX3q+L
h8Xo5+aeXAMrtVbeXYgJxbJ978zECeGOLompWXIofFomO11/A3+RBlggfhG/nCNAPtGbRCRbhS3r
I/LGxkzMe3tZflgKTDyi3CeG5eLYMoSFrC2zMiQ8uVOx6CjYvKu3uKhqymruIwE5M/+wOszAaZyi
phWwJAh5GqkGHu5zvVYDvJIAZEp4lD/QDAjwcFKrx7ChgSTOZQey+RYFfzaWaSINaSAmj15iHZ2f
6X9o9aQwZJPH/MO43qDswzmsjXQaVvaqvoXUxMNx4YwpeXE+4H6E3pKFsuOsVbYahrEGh9Zif2S8
cOYovwExTC192TXTAEjuj4GIVG1RNNfGxcHzhVLRXDH9devR5X+LXxGJpLw1XPwBgFL0o50rZOfl
MmMO7iZ5fsi6eLoHtar6n8isC0BX6MuekXgTJgNcbNwUfqj2EgsxRlxjKvOaNwa29CEOUzOz3Nvo
kyHjEIn+HUF5f3H0WUOytIjCG5xOdmfHZEsi8+lzCwKzJQskWxe0Z5QoYM/Jv5BuuSMUNOWhTEeu
KrcMMci6cqKvzev0LOGIjHCoHhy4Dq+zvGZY20g4OvDjCXioBVu9Ea0XxZOru6M5WiXnrRl8Ln2y
LUDr/DkmXOVskF+kY13HRDpoDGyvriTIF6/McG9XxhpZO/jEDlbiLl1O+COWonzqpPZlGbF0p6lV
53TNv8qtRS5FpbMeX/PylkPedyv9SvhcLwp2bRgJCPpgRRlIyazeDKsXK8x5QoAR/xJy14Nm2KdU
f76F9002yC+G1l3wUQ1+CIxRNTRqV5mkwvSG41xGT8E6F0fN/ws0DsFFUrm4v+W8WkG//XRw7mi4
3OxLbzcVkfwiW5EZCppsLVZqY8i+Qbt5R5GJMnwIfWaNzlFamfDbq458SusKMdqbLTrpgs3MQg2r
5/xk2xQohTsUqS5wV4aImD0EUvmthNX+5KRJhctGHMC/b/6snFgjGM116LXjWXrf/k25svsRXBjq
9gUUjjUAB0O2yRf+ilriJ7KlAMdlrOWn1F2ef5UrpTBjC7uEmFInqiMbo9W/x3+Dj7e5stPn4QJL
9rb0aBPr131bd14hPmsWWOwecVd1/G7/KnrWSPQcaLzKG7c98Rq6hDXwzcVaL9bLxZYVMuk6dn/J
4yjzqhzqIfum6AdnpZM1nIeSnIS/EUz7bC2JqjTMXo6FLf3wo4yEfrzIrSw1pl6O01KR5H1QHk+5
FX3z5HS7opnvLAtxMewtAEI/T/7znb7WarrM5D8aHmCPjaq0E88CEXqS105mIjYoMvExShM32VW9
FMSSTOu79tKQp+0ACd51jhyAVHwqP/JjG5mhFHWy1ZoMJGezOEqR8yA2HrMECVbHNtnMRsdCknVn
yf/y/I5G3SB0XJw8GTo6r5kkMUKm8ASheDKKF0sRCuRLehucxzkVQshjTo21iRRf22RE72Zqxda5
wk1rZj+v7PGqDbO9OLnD7w8+HvMjxuVyKZKX7uDDiKZmGCcoWzH/nmYx8tIFl6JRY2E69L6fSxD/
+l6PlqOWJ55NvbhL/QFOJpX83enFlmQOxIL90MqT+0QCIZg4jmYmOCRmm3WuaTYVfxY8EeigOHeI
OFL03LOiLC83nNyhuCEBJ8slJvhRjKJGLuu5u/UmV2pAIYRLJJLNMH+pI7TAf5NgbGg1CrecPxRO
MT0eUrzPAPrMfVUeEw4MpIrWA2rXIEOXyISPT3fAqNtCKcMH+RH6QJl6ncCCCrmWBtCBFw0iiKle
7rWNCPWNFXipGOXHCz7I/FpbwtpVU9sTb1VoAr8c76WaK/6ySc54kch0ZnzvPct2F5F45qUvgDSw
/gMcoMn5U6TBlKABuOJFNoMb2Nw40y0ogZ2uBOkflNIX+yuXbNDnxQejCNICrtG2MxBA4bbtauFD
ss9hDSwe6SR/Gxuo5AQrDqT6G9DSXtEVS/OINo82hMWJNHjxwZR7qUnaESTNQXnHmgzkr9MiXirX
M8K3/XF018ZDVPpxKynCYc39xkYR9K2jVJ6cwBV7/ka0YpSlj6t4/3/MUoBgKFSLk57z8zXvwnxe
9JvqcWheTBsAMEqrpHlpoD6zoLO1udKmtOCOIcuNQEQPikAYtVKgnVGGcW5KRJ4GKAP8wOlE1DhA
qRR7EQVloorrCPohAw8r8UQLhzm9Annapo/Ryia/IC10opUKYRQovVqORmOTPsAp02bgu6hIzCJg
osLcvZ1uAq9GkjQUvj1CP8zir4Bds45WY2gdHUvinwcpHhSQzSIpyQM8LnEV56iS24Dyt4ZRgdAF
8oUnjPMdNLSSf0q+SBpZLkMqyT3SREj91ziWDHJJsx/nz25hvIfIejlT+ftBdLCVn9eN0HFSW6rU
4H9VlXusnx/bLN/wVsnoTGSm7NqDyQBzPGQmtIa+SGYPv4wADpsPPC8OgU8RQwPplIngK/lm05Xl
6ZllQughSgFH9AV5mX+Eh2tKvSbvSy1Oj8VqfrIZIMlxSZ1knrqcS1EEesXVWNu0fxBcT81Zt3w0
Ml7nqGRTnwXNDvk2cHkOpegRoYdjhp1a0LLR9A6PSFhtfd8+t1PuTxD2ef5v7s/H0HCdMtD6LAvh
kLsdwEUMa7N8OEcRy2/a+QcRu0cT13gN2fA6y3EVidb4gA+zfgAVfiV4A8QACHRTotXcL8yN5h1L
rxZhrdpxkH0ALimRNsXyLdxH9LAsXLqnIgMa9pu+n27cnHNhcWiqMYN8WSMbeVjXZpEHAQ8t0YxA
9dvTnIBNqYxKPXJiY3kV1mX3PLIF95KIo27GIV4FGUzvJNnfZHkjOeYCSlfEkXg7sFMO4E1w947J
P8/vDFqpyS0800Sky33YL9jM2tBTQk+0G4NDGABWDAaDjWWoQzIIHxfv8cjB4G6t1A9F5H51Ex5m
obZDsciLa77gt7tUV00A13pRw4VdGDPXFSzSgIq/uVp5+yLH0zCxNaLH/QZP8l5Qxzuq13+7e9z0
vMQXSlrTzDu+ph3EO6fJ6sk5dFdQl7jLS0jGXM7USmn9+hUjazxXrl5R+FiuOSbRwxS13ee4J87z
av2pX0Ij6reIcTH13QjKb1kb///jvaR3Jelqu05Xr83smfRuUDxS77WWkNtxC2UHyNNrIsXfXJyC
Zh3rM/Q+V/n8DdenvssxkzsyKfBnhEPaHNVT14pVbXkQG6ZEFaQUDtEewG2nDe/VRjKXS5rU63Yq
r7/cq2dfPddvjDvKMASYlUu7KvFsma3YsV+7iNIl26oIC/lLSov3cSwb0luy+8Uhpo+vCRLNwp11
colRF/aDiNhS6N3QIvvikO1VBdwiH1/S2YtKkQWeTfSI8p5q++NbrooUCU8wFC+VsdQvqQDlWW41
wzsyAscWQHemSywaAFo5kx1U/YwLLuU9x524+ostuSlFf6QIJl7UBx3ewyUPDf65sXPHgh206zyn
ZM5WIdI/RvXf7jyrjH6IPJJ7L2kZxm/ijcKzdqRMH8by1v+7UYbcBoggdLrGh0ShXD3wYW2KjtB6
KKyY3ArbabR2mYZltq/akScZKUdEnsVRffQrN9hSfQEBg/SlJubkAEDurAaaQcLfl3VNFbAxXqUs
A1L5hOol7TiZNvckFKSUXGapOx08M37vlKdQ7MEreQbfmdoGBeNBz6jrqjp1CzcC4vl7Wbk0UFiZ
FXqYjTHJEXT2bBj6ta0ucGIjlPJ+/uzuS6MZ6sfWJC96POjfrDXRr9YLcW7+twhxBu+ZuKoanQdk
rZihWgkD19KOyh2EA809U/6GMLLHMDb/crYPHih5WHHmvdkXT5QxjlmFmSpO8/9wgzeEeV69Zu+O
N8R154zAgFMrgV6UoX1nNgk8zXPd857hPK3a2r8NinpMc6LK35lWOVZnNo7r1Sz8RrHvp52PTPnq
6MU3jM0kpv2nZaUIzGnIRANFESzClx5pghpeEbIudjbPZnKfSfvdRS2YHdWieCeAiueO0R027N/n
b2ifc/TQv4g7FlYMFiopMG4HDxNePvuxXIl6Wq0rYis8YZAfrWv88IebHhCOXU5pZWZq29bUC1e5
CyiV1s++jU5KFosXkaP/QwSe/MZCudmJnHTM9hRMTeACaunhanqnrvYBJPPJcQ1gYty1LTCHpXYy
wDGhMyj0b+YHYX71t9JXDPO2SJ6u07OMXkNrgiPucjLnOdSVfr1vYC8LPbsjlZGVxgbsA07SQZtw
jCfAKXbcoyZF2R5Hmbz1YbiCE/2XuNAWeP3iA4JOCvMb5RxO6GUkR+WOjUvnTrs8s6BsbNUSs6c6
u270NI8jwyTI2zisp1KFyM3X+ZPu5vhAGqPR6LpvZSnW9eM3Iuh3HLOWWGsCBfRvcrQibPjO31N2
qLOR7Cgs2HVAm50ZVcjLPXL/o1R5JU2wnWbh2r9k5zphZP/VXhLA89PwyOk98iBIrCLuSvPeFtLq
v/eVao5YZF79+eNKlsaYLvnXrOBN+GxsitpN0SaNDctp9SN8GkeqdG0zV4yY6nhmYant0E2GBRaQ
m9qHh4PWkIQXEmNy/QZDA87dnRlBFOk7BatVQflxzJpaSNFJJSWEOOX3Py2dt9mDR9rIfEgofsws
I0cqvcBMxuHXPw2EAiFMPtVZY69naumao8Icovvkl6GtT64G5jGOCt8YEXQ8UTmBcd9mFkF1PsRQ
T3OXlkyrfxRoO1fjrsOGJJprRwNbo8lt41a3f5ELXhGFXduuJmRwS8cin93kPz2IzKjiz/V2AbSA
y0kD6NQybj53ISvSTCISceZrzB7+qnNkmwV2PDgu0emLB9YNV1V2yKvc6eCEU+mlQi3N2ra52mTe
uH5FYfd+MWzT0yZWpvmj7Atps5waHNwS0WLPU/YRjdoxohaFuPevhT5dq14BzMRbtgfYvXGqzYGQ
bBtCrkt2Hd1PTewiCxj+qQIuim2H5NjpLxbG9JQL2BFWJaqPzFXgsYYN5gJdZXTHBPxADmsXkV9z
lFuGzAMA9oUgfIaUkCyecnyys81Iku2BLC3RbOLaLJz8mUPBq5bsVm5xKP/m1xlRnTv8gmOz8o1a
28NbwRu0qPWSYMgLJ3tSuRi7Y7SYyCb9rfCplhnZIwvbuOFoEWUzFg4X5qAoavry4KOeb77oCbrL
dAPjMB4101HX7CsJB8BfpyCNPKdhbW6jh9T0/sDHaGer7v80SkvvpZQGhsu+1rtfctU2N4Z0WD/S
mrsSbojCYQTCsrYfUP1x7Me6NDLKODqRolmDBMQqTx+SLoBofaKnmkVwa+MJs5vVbBf/nIVNfyeZ
KtK6z9TQKOLt+BMKVePUsp/+u6zIZb0QU7Q/e1nwa8eIVF4647qtMktYHxX085LK3VZB4ouXBqw8
dqWQSa58RRwJOYDq8FQD1j+JmRZfc1xesACY16OIaL+OaIUQqenaSngCWu/CwVXgetuh49tFxdMO
n68ewBPp0bD0ZDa91aLexSsTgW2c16B7xZ/lW1J7ie3+ME59LVRhcEYiEqUm/JsoOLNwUqsOHl4K
tEvAe0FAjUxgNxaOvzQQfehyYQm5M67OCFNMBKdkqFDgna+wwy7FekntWndSdKDs3ZXpC2ucRD7y
bOQHEmJPrKW/hiSjZCtWQLdCUHgV4bmuLkQ7aeTYECn1SLWUqaghn/1ffRjN6t0V7J5n5and1LHT
FOY6jTVwWGZD35bOjuv0Z0l8vv2yL7BFtYS8s+euSQ+XBbz7UeIKydYRO3CXzbvk/VQKl2AgeK8y
MBZ/RusFrfzwh79BZWphyAQZrwPNItGu8gnEhb9lFvCBK7+lytTJSFFMC7/Ebn4iG4qL9FFtlpFR
PIRZk4s7W3VetgKX2lNg6TrjDFtRP02Tpa7D7WBQpOIZadVy15/ym2Rpc8wL9sUxd9/IHg7YWHDt
PEUWbL/YMik22RD36wzmvtjXHdnMn8RyAZCJJIzGjfFjrmRd8DLr46xA0LJxnS0zWOLJewmAPcHn
0xvSBrXO+uZNI5VVM1fFXFX5M2k5vAE+cWM20oPG/PAV7YsZqj1QAXc89lOne66pTE4cepSAAali
Lap4TLxjA/k/rUvc86O5Tp5CIRDRIFhK1gAqL9QMA/QG9qoIrxHuIv9mQinZsyGxYSBehqeEunjE
ahUv5jBa/yanonhmjD5XbaTbdlg8rsMiUuRpMyRUzK9mF8T5oR/e88VqdISefv13l1ah6vrI6iq6
dH6hGFbwIsUOv5HYcYxmLCOh7BEE4xC222qA2EtUUeeLFE8whQ93a0SALt14L25FK53oxAW3AlCK
B1rxCK9SquLe7vIfeQdL+pnXurVgx0n3cihqqslj78RV7VBzY/X8qdNr5eb2oRyftIGO8/lIBCrL
WC2jVwZrtgTWiEgZEBexP+tmhhtegRFbbH7joyKBW233JgJpWJtmSph8IDacmMtwsf8yYW6DTnkA
jPxquxgVazdUN+mQS8RsoXb+rErXeWGxH9ineB1rRITFrezUAh4kCoJgoaJrpPbXy7dXkTtfKr46
TZhfPO8iDQZeTv6tFEduCrEi+/2GQpObjCdo4zYHxnK8LWDlFyc0PbJxjZF1Y4vuCuELn35T6zp8
h7+X8wVTxkDn5YqvkqdAWJG8gVknAEnAnrz10y+q1wvdwX8pmIH45DPA49BF6T4/rInPCbX+YobY
8rDpaDxGHv0lhyr38FeKnKGKAM6D04i8OEFSNwktGEBJcgH/P2bYA+F4H1QALPxfhHGzYipwBmo1
ABt7rArHbF1yo6M0YI0NDqP+UYt3K1fsM99E9LcRXh+f1yA2sZq9U3ViMqft+yjVaEOn8W87nfbk
ODSp2+FOe/EI9uB02/qYcFcSKTAO+gV+SSbwNuKMYYW3WCh0CjGOg+FshqdzqjB0rm8VsvUhqcG6
phUXaxj2HBkieNdEj4BlQ51cntwJwHsvkAR7lkiutgbvTyIXWFwYmNwhaG/PbhSbwpMnyk944Wmq
hvhwMrf3dFjI1CTKeQcgeAxrV/yQt1WET8BbrOc5Ofoe2Jyrl7XUaZQX+JDquvPaf0djFiXL32hL
nffj/VlKYVZx1soXNkIvhswvNCfcYjKWesSPH7XIYApRmdyj+OwrTfEhO5tkst42TLcUDCSYNvQi
Uq4WQGuRXJu6nlXvHau3xxt5UxBFARZDzmnVcaaN8zVfGsgxwpYW1hrcFfMDcSlRMledDuqpzrw7
gKkEh9Z7Q12f+HPE3l4eOh0a5RACQyNLMNaAhargcLvMG3sl12xtnuRoosHlxLikyD+ErTYmXIPC
mheQ/q85/z45H41SBRrXDyZw3Gv6/Y1l7lgqkSNkLFhgUwGIxzXlPt+54fFv6dMAHXvw1ve/gD1R
AJ4zTtJcLoLnpCocNokg4k5817WZFWf3Gbwcr9i6JN6Y2OEKLUSo5qEOBnCtn17ef+e9hdQSWFbI
QwD6IaSmrNOK3tW10vfLoJgkGq/5tZysw4zDkMw93gDrKPfAt5rAf61cG+/M1N/tCtdud56i6/iB
rkzxa0mvSazfDsVts86Cz8HlDGKvvKGOBLJYWl8hhW9Dprnpo/Z47/mQx0lrv6LMFfd45482QU5E
qGd1Ifpu+jcibr0QC4BNByUhim0+rp0u6b6WfalNqaV/FoLp9JWt3tuntMWSZ/BCdplRSuYZlN1M
9VJYZ5GKxlqbQlL0PfUGldXF7yzjpDQJmM8OJdXWKR8cAUkaEW7e43pJPAool3ELtjeV3C+ncYr8
uc/FU/YvRs5Flj/19+KLhHbETaCyewlPfqgH8Ucy85KbiYsn3McK3vfGx4vgaY1BxvTfIkh6t4lr
uUf6RVXFlNPhbOU4OvsTASgWNv/0sUl1uBLe/dnkaODreBrocMjZSVI9oo1a04MvkrRkyDIVug+0
I59OtsStFgmzoace7c1KC8Mq4l1Frj3ggbzRdKZ4nMvTOtCBVoSWVHGFdYb9+kg3uSOEbI6WE5XG
Ir/shfwzxH3u2n0nfJ61QG3Kpox+d4a4sfrI9M/WOtgUpCeC5NQEwJsFxV+ZEyG84TUxd0nwB4sr
Q5RclGKyFzZUt7z2h1KFik47YA5bi1mVrtKkIAW4iJl3FCgao3Uxyr410aD17iXl2Oh/YVmT9hxZ
cxeXtNibox4FJwS11bdaF9ktgFoRwaGrgB1GEAME85pQRl/oTbcezZbjqxrxDg0GL8k0wuBKM5UK
SmnDObzeEiEIq+4s6xRNGd3u3200RxUj72ckhZju/B711utDg2SzUustH/UDhsZ+MdFxRBoqOGpE
g4BUkGC58i0dfTexrH5JEQ57YG6XifwB8JqmqsIXo/IDy6GYt5xovl9B650s0vwoEFu3WW2up/1u
zGM0KFX1nnWX2OYltmAT56/aqiVlOMdxZ8rMI+MRzYLvb2bwNevHMf2Fli3P3hpnNubpj/wGp0Du
LjwZxm2E7ULUKslCJFTdAKYTb1Ub+Cygj7FU6jFZXRB39Ag6GE2PdsFoOwNTe0OntJR/LB0T6U8n
1LThTFASd6bpIdGoIX8YATCLLOIs5Mt/oxCUqg2nk0iNluBSnGc8i8WqzW4+7QyjW0zj2XD+i1+l
sc7kvipACnSrgzlbyCkuU4v09uliwfR/ZVhvtm9/kMkLqqt0kM8y8esdN+JpyQC7dQwaodh7+lGy
CVi1ZtUwyihWWG716TJICRf1BeM0vxmVm58YJhI/fabKh4UbwkJkyWt0AwJxiIH6R9DjP/ViocdH
i8YtUdNl4Zqr9CBMzzpxzPL+vuPrPaSx+2wm7YSMuunBzahU5rFVqiUhCy82k0i96RCsmIf8Pzl1
T+au3UBjQAVGXBzGV9fZGudJvPM7Uz49KH5BLL+kVVNcDDoGjBVpT9RfOQu1t0OJptsozC1EQEHr
4mv3wQJgcf9V9itE7hFyOTfNOm/XOnY1nVu93Eo95QdS2yfDxwblDGI5HxRoL6NitVpaN0+ELpGN
aQxwwAg88XF6bzjyFavPBSyw5mNrlIre7QDCrS+BIc8hAQutwkbzeiGX4wGJ/HrJy1UndUr6guvf
JupsYYdV1CbrR8s5Se45lXxA57DSHqJknRtf18Q1jFTppiRJmq5hdVtILcWNKxKHMWNOrIq0u3DB
F2LwsACJveAKoG3h3HzvgCUdpXG/ksTO9JX+kQgRwIUsQRBzJ6fxQsvl6vwu4YYl7KWdKoKDWiTi
8EzcN1zxjClVRbmzAPHe9RfzG3GdZt6djac1zOHDg5NOqMr+ajLGIN8DueQPFhIVlaiZD2bNLi3C
rnPwtuWxVMO3Wzet5Ye0O9vDnUC0B9qS86sKicfYs7Fj+kbzlDd0Vbsx+lAJr+LCUonQFYcmYxk7
/RgO3Q9TukGMI0M55KeVEPLf6urbIHFJ3mWYr4a7/i+z2HzeWbgVkZbJL4IpatwimVzSi7SeTlf7
XS6p2MGN/51eOX106QtFc65GL6OQ3S8BxhHhNw9kloYctGCMIhIkwuDB62e2iwpfWwh8O6rNSpjc
CpIck5D4UY3qFKsQYVyU2pXIXDo0tmvTp78UrqnB/8ElTZxK+3dziKo/Z6ifw12lBDh5dJz5r6CT
RP/oexGbhl5oz4ewgOGpccaFEpEMRizSp2J/b0qHZD4nFU7XrgTwJIQY/LP4OgsWOO7Ul0PziTON
SHby9Z+Q16HH5pS602OphVICLZIrh4i2bQ8ncG26aXHilV+ox4VszzlLxekdPKwwN6vuGqnWtv4a
uY3RuglcrKc78lyajncrwsSFZxwhZgm5LizTBv3V69cXxn8D7/m3rlO7y+DELz31iSmaAjo8ynnX
FSonV8jfvXou9hGRvfVttmXjZb6NRFy/Gb/J/kT3Xls5jfequKLiTjmfz5qVECDekPit6g6iLu/f
CbLEkITwF573BPRPkMqp08pqBI1gIEakaZ8g9CXDhNQl9SpaBvwFmUY8osX21wmXY7uocUFMUVTa
CYjMWXVXT0glNLHEdINxoSmpfWKv5HVUjyNvfR+XEKEdj99pB8yVvyDcA7I/XfCGXgaBT4Jwa5cR
LfWk+rCTqKq2vgEZqh3eShknU1L2R7363YCnaPYnsIva2iYxXPs9nCc3T+rqmt/CA45L7p8/TfHr
GgkfTSmsDN6SCxGsZXQ2KJ/ZjCkCRssOIHIdw2U86ybHzWgaQL6vLJSd4DJ03uZf6WRTFfH9QNM8
lyp3miesrjvbotMdh7Tci9K932xb1uGTMBHSyB5vF5pA9eld2vJddBJA9wswTraESMGHq3jv0Tzy
HC4Jc0/kJPsJfexeRIAOuP4jnaAyMeib2O3UXHAcRbcjbKeZRYCTtth3a5QDzTVNJvTxsnckakL+
bxbObJIjolE5DVTtzfUPfQdk6mMpfwHfjBTIs/WgMJeijjPNupBSNAwl+0HVZ5SJakUNgfHxzBTg
xpdSaoenut+mxCMJUBvBQgPkbFV/yHE+pdFR+vf07Jcbo/TXuQxjw1Eij0Nnb47v8MLklHKco9z7
u0iXbB/zSPVKnX6XOD4D/6ma8lhukWgVScie8O1vcHuyT3m2srvJrpQjkSApaTSVNmvAll3Hf2WD
Ca67LMDRS94ji08Isr9Tl2cCknx2E+pgLRC4m8DD89YKM5Nre2S0V+zBAmIqmOeMvsYxmwUMsARp
PhOBAX767NVw8FQ51Gk+Mv4Mll4JnOz5iF3yAkxIfAc4F94g5FxO/KocXDkudOYcD3POHFynSU8E
Y5SmOFpZmGA4Gc2/P5q4uS5KH9CYA/t2BePA+66Sigf1GxIEIlAdtHFAPrO0u6fwJgPc3oca7Smp
XnJt8qiuXhDQ8xuvh7p6RHKEspwbtScjwG0jlXuAuepmTSm3pPXcTwYPQODEbolXIQWF2njEcF6l
fh/ExBBJeC6Oqbu4ya5+eP62x3KSlQmOmi8gAgAdhxC4+OcPKZH4TA8ZyV/1aCIDTaYktXhW+dfL
avIZV0kjzVqvckONmBWa8581WGhkiOMwyx4AUCqKHrYLNeoOY06o81iPOmpGLB5TQxxpGZD7Q72f
Im+PJcXykCRW497+px2vn4Gv7p1aQIMG9qhFSff02UiQFtk5jM9XeMmpH5F24ULSjL4Acd3kC/OR
tdIGjXfVgvILPzEPJNc2cdO2JOhiQMWhJ8DAstXnxdEwxuNv3+dyEbL7+XKcWJWFijV+lG1HikC/
N05X+S1CEaJAzWbqYY980Bp28tMqGjksFPumjlsj6+g1CVMPPFRkc6AGz5iVtDHyoa60whvQaFia
S2mjc5FetPB7aLA3M96DRNCQTIGxdO9D0oKY+us03uX2ZzFZvhYoSpFRXKcOxPmYUaiXHhshYuL1
hgdMnCzIIBReK59A8yI9Tv1eEhiYcykbsWNbcN+E+r5YGD8+juYqh4wm+NsALHPRQJvjKqSX67Rc
TtoNvj5AKQ5Ln5qRwuMBiJH+7sA2h2vlaSeGvQfeWEyq4fKlpQ7XeX5th8S5lrvpF7OBeegUynfd
6apoY+K1zUaZPyYccreHwIsMdjRthbwvc15Pp1uog5SUIYPo0JLKVGVLQMo7zkH94d94SpKWfL9M
9PLUwGi8kU09m/dilFVFq3AeMkgUhUNZ4evn5zahQUomK6LU6rN+6Ybyv9B4KnTYYaNjLl+pzbbF
SZ4eSVkxXj51nsloV4eQeADsephWL/WlEsfyvR7evQDBNMdyAgrlDarBudrHV9An5XX3c/RBvlS0
qxPh+57hNzgJ45gxjelch8+k200nf81RlWKVaNzY0FHZp8OKVYtgMsvIp+nbAz/xUjn9ENXZFfQg
IpzrR9sGAq4G2722fqX6G6pflJLfEakG6ZEbOTZ098LfIKsNLp8gVvAY3Em7J6NFM6Wk5u4J5fwh
rBsrmFWhafrDYOzGwa2zVtLxcvVjTzuSTYSJOjNVu8t+EvNcHBHsurO6bMaxXw4ko0BTP1A3j9zP
D10H0NiQSk6padBGv0e7ewV8LziliOxt3HmBzxbSF4BJDk6pMBD5CrZGHbaIBbfDLwt1uZ0ioOAj
sKZT7RlAN8MVhlOafAlKDxPtUS3/AU1KW6Aq0r7KKUbems+NDhGXY9l/4K3uzFzU0OAoF/tgjJrW
389JNuRDJoVN0bl6IHWi2UhkwNGGPKtfgAavpIxdmPLEVUB0vpIOPFJOMRqK1zHcKtEJ/d4D1tpU
Iz9EMJjZO5Puua3LbpYwKFo65fbtCW3zWu3TFgPhOaCvV8w//umTuyY4t+obyVCersJwtGpkKp4l
Jnh1+GLojijwmXFP/5STP3Nx1aYPD+HXuEhK2Sk68REevR55NHQMHgqE7QEEEokfC20153kCUieb
qxts/ZRjU9oNGOg1thkE3JeS7/8IvHHgljxhdTJ2wFlHJhaVxhwuDiCNYoz8z8sETHr+DAthEt5J
jLiAbAGXRP7yt62WG79V7tBUS1xhyJ6Kz0GLW3s/+S7O5b7U2Y4+kVWHX4ogTxZX7XfP0dUP0PwQ
bQ9Ne2wyMEvlzSYIJ1YQfkLGkkyvBPQ41tOI5yfoaRRbnQIE3xeYQVjIkQX26ecQTBG7A/TVUd6a
SuJ2dxbcP0q2XWIT3qhutcwQLDZQJcluXxRGxRXOgAWaPY4Rwi4Z4AxjHgs3rtI3CCB0vkZUgqlW
/BDaKv6V8pzetcbZgfwcDPcjwIZevvQug4x7WJLf8iirf4L1yLNIL1phXNXdIKiLok8k4Kev8zXi
T1ZV/8M0MP/L/6UKXT6zu3BGNXJ6AV5nqJYyA2BbSPFbvuhcNeMga0fciJ7Bez08oo7cn7jylfWG
WAFnz1u8p0ebkmZi1wJ1cWkSt2dDxIvX/UyucV6vCXDKJ/nkd8dDq7m0YEcVWdN0ewpCdKtKkv+6
mNJprJIAxG5BhbXIxrmqRPTkQAcYNhhpZ4OxOp+FuTCqLW14QJCpak4mnzjGc/nevH1pSLDIDM0N
/kEIRARMghuwE2zYXoDvUKQrbODNEjUfoynNo4aqggCLWyCEmUgEHpMHGQuQULdx4zR9SfvnlxTO
YgRsutOh14h2x23QmuhBLMPKKptf7uURGbZkRqHBBSXWcjYg8fkvAUyKN8b+yVjyRokujxPHJfFO
EE9vND9JHeFtTZEJ2T59ZlRX3WNS47eFyyBcgoqml7Ykal3PX3UDU5ii7Nc9H65yxIT7kxx3/lLo
X2PkU3WzzqZIVRV6XidqMPNQ8mCWE0xPTU5rZnGqFZcmM0XaabDdZLAJcYu53TTKXeNOwhRMOx6q
Er8VpkdZ48k2fh53KVxuGfvRRLG9duDO+GU9hWzM5sFiPFm99w/JX3xn5tkgxfNgWbNwP2vy+N1d
GoJ3jEMHrU9wZnJRSvhkMrM01OkQ5Zf6/YDynJJh4rbSi78uv7bbJnrkycpXjQO29YD0djkXz771
kpMogEC6Av7oxkZxGnUzSmiFMx6Y+jvRrPx8dmMYPK4uN1Mo5pRb00XL6rE46fkJ8KlvKvqqTth3
B1isTTwY7lNNL/VS972edZy27kZjN2JYRQYYzzUlb4UGcizto5nPk0YcDfGkeV0CyiLNGYv4JJV2
IieuCAgxaBfONM/LQG218c0eIM4FUQ7yMW6awr+8MjfT7IAGXpBJ8F5kMEmCbdQ8ZyEHFQq/LFBv
suJ/x0DsHNDvK5ApkUsVYRmi13okKw4/mNJWb8oxOTzUz+rx8lpy1Vsz+kDf6GYlnUH/XfUz1R7p
bPAZITdtih6qWQ9Zm/sJU1T0QTVIZAjbZ+KFElxRnuZ89yN/D99ziQ82cMF77rlGvcJMFTkn/gib
5qhTm+kkg1n+BlNGENnJz6CkPcEcfdsHFMiM+rTZyAargukeKsvs4idQDOrCap2gibohLQpQXgvb
LnP36UQ0nzRtrsN3wLam/FieBDGN6MYrDOBvdq0eh+k+DYuZlsIU3is846I6/ASZDTy0uPjs9USa
o5h5Er1c6fSeoAImLlZH0tijmxMT8+uZUKEvCaE2Z41l5gldf2v1xt2D9x3HQcHARV361xzojsDq
y6N0ViPa+KtURWOv48tt78+Nin+6z7hp9ugUsthw5zj+VarR/lYPlykmfsV98mtnn7RSdQBfETts
Z0vidjoPNG1WMZkpae/p5LwDFo23cRnsioFlxnCsZU9G0sad5MgYHPYODNWv7v6ffAsvLeQjxeoH
JV7tOCWWsiw9+imnGU8tkJZfl6EhOBrXcaOJ20xV3OG56HMZhc6aI8SafBJq2kFhOihVBMbmahCf
obm14qSPH7IRoXDDhb+42LUNSaxbHRpK9ludL9WFxz+VEAMhsm6hacHNdgeHdeT0epb/Rf+YSVQq
nsvWpxqrkPUqgBAs/iy5DjloaCwc9g6Ft8/R4DWbXG/1W61Y7zkWMT9558Jj9akUnga98HgPuMws
jNZsWGNUq2SB0W4RSJkTFFKUuSmGvKZ6dJPMo8KUu6CH2ijAaTTYHk8uHJaBWZvmrGcQ4cI8YhyL
YiMSXHRG5vVX0HEPLOJJyjKJ6ds+7tx93LINq38fh2ILhHxpF7t5Sd7/oJ6Uw/pcdaXk8B/I/zz+
i9mu/lE5SIZbGVOKrU5gkAFJYkmEYYDfo3jewOYoD4gzE6zEVNxQipA63AmVZ3kgNU4q6g2J6o6d
9x0Q20++nRKN1Ra0do01Sq0iIm/TTxp0FCpnv45ABTi4yp4JeSn9SAmrtReGiPH72v51B6Oj0Ykv
g1PNe7ooh1fS8dPfZqt4kh6Rbr0b7DsMrQfrScSzsItWJ/zyHzp53KzXzctaQId9pndYN0E4ZJpN
jx92f+ZBHNGLOM1p54gGEGykFbeoYRGvuC4jbWcGVGCt7zyfr9TwpTkJi+m44rW60JMwWvnIeqQL
fv+P7GClq9wrXFnZdnZmjb+UZjsqq6Sv7gvm52laoloAIji/YYhNPOvL7B7Hn4gp3dCDQ+1KAeG5
FLQEJ4pJ3vVTZvXWjqlqjV0p+E6VxmyrKc5VjLLeMaN5C8HxqZJeG+lfh5QBTfCDC/9ntc/6StNk
1sDB9vk4K1CPv93kKrVpbDYuAfWtJ/nxmBBusD9WdgDO0xX+u5WwBELirPR1DsWDgKQU9aoyH5Hm
3pyw4ShUmeNmadqpTP168nYN6eZiuFZvRUOeAqVw+CeUc43lPezsBuQNbsb4xlZwH3G8D8Pb6CRa
0vycH6p9G8AkcrxQ3Va922LO0M5564q2ky9sgcKeb5B4MHtLEDnNHEAm6uVwdEkDVUEl2SKCdKXM
T/Ad+dE6ABpYnbogKS0qZf5f3JUUPf+X+u0rUFlDtIbsPbOF5zZ+jqjXE6Tm59irDquJTxKTEqY3
oELXYZCSjkctYImcV6RWJR6hbvM/y1FEFXw8DtxLs2JGa4wjpe1TUDlsByymv7PHBjm/WQns4cAx
IJGplwauhLtB6s7EQwIveavfQeOpg/w0068wFCWoVjSV6WO/TfW0ir+rJ4dOj7JRqNFRVfKOHOgK
aZ07Md8xafn31Gdgswovi6Ez0684t99TLt3s3Iy60tiNZ1Po1rOpwXNeSwRU6Uq6DSVoM+iUFGCI
5y942DUjJ9WRQy0ddyLlK5eACZUNtcPBgEMv7QgeAsmZeMeVoSXpNnfnQZwsx3kgpNx8DHvzHQq5
9IoeCG7oiWuFvCwajZH/d+7mfCGfjCKsF7R/eNU678sU+uzSwnhgY7hs2vggEC1nVY8uyqtEp51H
Xu2IUS7yXnMVRWrZ5Oa9ZaTRm80z9qmnAla+3bkKFwO5QJKnmYhNq2W31oFbZFPoi7eg8mVC7Enz
Dj7H3pmskcgnqjuphx21tuhpHtTWiEnxETT0Cxf+nPYbVRpgOHlW1fDPGfK+AT6t33xDbg2aDfdo
MDlyoMEC28FjMKyAofTA2/V1Dn10v/Ob09Kpq3E30k08CH1Dhd57rQgJMvDO7QBo+kyfM40LxqbR
m9ol47SmLEi74LzUdeAtm8Jocvyj/kB7cf9keKZnniDkyKJNPG1PQ5Ye0deJe7tqVwSEMkUEgxGE
G9VbA8AK49rU7eVAVhvnKJ3Afaho8veVCgM8w/rb+li/taLZOg5iYzYrCbRbEhlUc6Q/3wn7PW8N
spbpvgQdUXX5IpAHIlp4SQwwHBJw0VTDUFACCSyC3GZyL50l1BinOU2ZsnOdAA6y3xJSyVglxvUN
ekdb4t/Fk7h8OvNxMZ04dj+I7dB8+6rzfKc/QJhIGsVqT7JRxQXJ0EJ9ztRX4+zaSNfuETXaPnSK
aY3/PUZAemM899cFv0h2fnz5rIbrYv0DUrYRhaiZHhv3a2dWt6RkIWxvOHLq10wiCiBa8N0KmH4y
ekMCRN1bd6r6S4FyCyCMG2GxojyGjcT875m0/G1cWxMFY+XmGgYYAy4+qjgNBJV8TUBbSbLw951D
zEzDYF7TWj3qlqZnxztoXZ6wW6wZWlUoiAxbugBOLvz1RBeXErnWwIR3QIvXZnr2/hP9QJdMkmK7
d0gsIxQagDaGSwHvBgP9WoUj1iukkgS4OpXlB/NxK3cuTU7DZkOFDGpCvDgmMSCeL/PLpyEKkojR
RMJnHy2czjVsohBsB2CwY1say5JyJVXFnZ+WbUEvE1M1TxdTBh4MgDSuPWy47wH/54S3EWkqpTtO
9xzPxQVYbrZe6D8qSYSJ/UVre6fXF21eHK2jEJFtDlazZA1sM6dclqJL3LS5KnI11S9LMqxbTSY+
KHVrzDnHereE1D6gXfq/OrUPdad78WR8ybcJjyvkCZ1oODQzFTqzS3eUHco0D/tU91p/W7O90pSe
srJa93+95fkXQ7GAdqe3ZT9P0Dp+WrSA8Etf8ogZWt6tbLTTGf4IpSkMPXJCO42ZZULLUmzApVnT
QimusLuMIbsxuVYmMdqbivw9emLIq+RI3NRS6sh6Lpyj/NkiokutGYDwHK5RFTKuKW5JfMoCgobV
aFKjPy4k9/0E6Cn9MgvCHBv+Um2RQxxjxOGpPxY1rlvekCCgagxrCd/3gjazK9k+ceSSNyA91/f8
SREC+flyqu3ruMaVwuIxTM3pNbNWVhmu7Ts+d/33a0u6Oe3R2xHMa03BuCBCTzoNpiNvdRyB+vpa
ipZ+7zhbrHm7u/cD3vV1HdKzAbn5Dy9XUaFH6fpoo0W+P7cboxOet5A6nnPvFbmOxmlCuxuvdoRg
ydXC3THhU0sTVkdNjc8QNVZUkwbMMiyTxHQU75RSh/hltCfewjFqPDPBeXQWL/pigXU3a5iCXA0/
TKZ3zAGdgkC98ynRlde7FXDAVbY/YqjvruhMiPC6mo7/BqFYkkzHlWqbvrke5htp1HTcgTFLiia4
xYS131bQPz8cM05LyoCCp0DdvxyTDBHZNOPShB8AnL/yUSoE28pqF93ygixRN9GVzqlbyxqrO9IZ
qnZAP9U6jRgkjso9mRI7alyvoRH+y3L8RYtxvhkJ4ww/9bj7E0FcevBQ9Y2JD6PpHk8V5szotPA9
HZPvPMN5elb2qUMWFiHPD+LuchKsfVGN2oRf/Q//j0dI/smFSMZMoBevE1RekQ7D8da/YPr8IMo2
6T38CNAhLFkl5BTApcl63UMpd1VKTXcq7q3ND+EgUrR2E8TcaitAitMmwMPvBSNfRqem51pFu+HH
mjCC+ER334plbAafVXSBVZqy33JdsWnFKrESzjMukUfuE1/QqavDBdJk6Lj1HxtoEWKUl4+NjpQ8
JuAQKXJuqjE/FTYfOjMH1zpgX0bwawI0Eo9oN0q1F2GGs1z1SfDx6pttk8U4EBjEczTHuQDvy6NY
S+vqFbJ8lTvZSPND+Bp7IxSfIEmG2nm5cdGtCLGWwf3GKLp4XA+n3YfvZ5wqK/glm+nW0wrtrfSg
JUcbVaHqUhNu5fLuLo9lKcU3CYi3FWtWFEjCoiBQjYOuFI2eYH6FLi68DCctNV7MhUBtyU1AM4DR
xzB9w3WFB6OiuzGfRLBvyjmjv6Xxn/GCexmApPaNuTe76W/4OPT4FEHGRF8utlJVGe3RyE120w7g
hDYjq0Nvvoq5IPqYMS2039/gHG6jRw9MS7qZp47GrAajPpF9//U8e63ncFixVeDc0APpiAoHdjFZ
a2cJqy7AStQe5NdI2/3L6kUFsmz3Ylv4jW9NfRtE7rw/9/YBYRjMgQeftEbDRTDm+LcYYVZR/a6k
wGKxSPknP7wu9QFvD6nUqC/f+09YgCPg+ZKN7iNwMgR77pdAP6rg6hcB3Hd20KKyWQ0y4fgfoFBw
wL+G+4F7nWN9tlcg2nN6/sGF6pGNzmHzYgefuWjOMa/gY+E/LMkf/UlpgMZmxEq/ui6/WQLh1ebr
fqGPftj9P406tmfep23EfF8iBcdxROBvTkB6nR7S6oXf8WQ18bmLjLxcNdN8DDLLiElN+a8wMqr9
beIeoNMo8/UTsWuTV8dbnM55lGlaonCv+OFmnxXKzwc0sAoRszwWN3OkeLlXUFQ++bDUrj9iEoYt
e5WiGNBIupdGnN7bJXkl8sRUt1cC2nvFgxW+wU8LodOnIrYPwkdxJ3Tb8Ug65s8yrfYtn8UlJthO
Sqh0nY8ZUb44D6SIXSGsuK3Pmw2mp9xkQ6Kj0lkEFzkSDBCJcecaAxW9mtDiXyzoN6Q3H82MGGuo
dWNJRX2pnisgPoUXJbV/ZQXWfTZZ1Ep4QRGfUR50b/0VIsK+sh5UlQnnEg6VnNJcNPl/wY763OEM
/mrs3JOfqJ5b5Bxl6h/ncR5mSAd0m6FkrS8oeqotong/3hl9KSSfkr1ieOEp2iBIGslrCI6MVTW1
MnnmFm2C3bXYH0tUyHGOezfCM8oa2QywnI71DMjWNSSwWbhGWojXWMgljhhZOliosnuGsfC3KAnO
J92w2ORdK/l0f1J3SNgpX9OFj1Yp5ddnON2Yqd2qq5hd6Y3CjMQCtzDy8YdrdRERwWZQRCY6uUZq
2GXZltSxzqqlJIX/KB4duhpzPdmRH58Z9Qp5AOBReiyF7qhzSTnhZrGPIquT9tOTm0RrScPav01Q
b3ARo9yXUH8zLOZGV/MYzxyjgx19AAqZoLXEuk65U8MHMVMsmd7NkW826OwLzxg0wwo/B0xrSuDZ
Btv7b5KLQKI/ZFz9HTCEyTOGjtaeWSI3MctrM5w7LcoAKadh9cYP/eX8GNG0Vy/ZGp3Wtbafd2hD
HXvXoy2gaIValMORy1ykP23yQ8UhQEwzLslgHoo8RvloOjcjXUN1hLR08kor6H3wx8QaOybayTs9
QTwPuhU2gTg8w9CPDYnfC8cXs4O/KWZxJ2PhSxjzQrATZASCmt1i3lGtuDMppXSfI60NAYFiI8KM
hmrVPetKFN/72rjMgz6+7UJ6g1/RmQaWZwuvGCeJ05x5Ea1Ez/KTtSiYps5uhQYYNeWyovN/ZwQe
Jf5NDyHOTaj+P1nApdqmQWlXgDIbEsL7UUiCibo2IB/BZxj0O79Zch1u1GAsHloKXsY4wwvhXP1A
FvzGWI/+x0xQqxrL8/Obq9iiQ9oB/A5rmFXNENeXYYIvqjl4BTS4/qqDNA4qvlWlUHMq6RH2gxjq
DuoRZPdDn0xRNCg/TsZEEoW9uTXnB4WhA6mcHr4LMiX57UkFSpSmM0aZ16LS1b9k3JG6liwtu3L2
qmjghIEizcWZlfi1MOlUrkg/cFgtpihfRdrXfYPwpJE+dMyYlVYo67FDA/g+Fa2IWNulQrYCV1Rt
cZar5Jb9OhSADGjWaPkGdO/tU8fOUsRuHl2DmuqbDJFp3P6xFbVuCyduPCS4hxOxI84Rbt8k6bfK
67EGMsoqAcxcSLFh/b81M6QbluAcbQeeJLzK/8jazFN9WLHUL90Im05kVzfUX2uVPPAgPDQySb1A
bZtNAhRmbkzg+VABnqtRrg1Js6MPlvaVfV+D6m2rCa8gij7r0CP4nI3DWKS1omB7LMo5J8SoADY0
+uasSW/f9qI6mb9HWGy7lyT50orikLwjg6H7duQwz0begPQtaxWd5CTBuX++1KMkDtk5N5rWSzvF
r6kberhorhkUb7AIfkPYuJWVSsefk/es0NWrThHs6hrnCbxZCJHuZ7haVLmHNWfbldDmP0lHrT9/
YTHOJWd2brpitacysv0/c146fBXQ1Q+nEU0yMznooCZDdBo0+zS7DysURx59obl7SD0Uwg7Y7EAp
cvx+Nl2pGK/BrY/AFlLjHkYJIRTSfybZPBi2r/zRuXEvka0H9mMEfgVRFd3VZXNBkZ0WQQHoNj0H
rXy+cNuruN+UShdRyZ3820zCham9kMY6Q/8dgHNoFzyhNhLJfBga9MgYsE2+ZkdyP3obUAt7Qxvy
876xXNTvUByJ7nT68LM5JEVVyzmHZmEidMTz5ypU4bt3NXQBuZAXgmJecSSsxXlyaH6ful2xVRsz
ncWknpRYXMprQcj6bxTuvCxW6F39Tvwkt8S+vUf6xQdkYRI7JwNgm3OpduEc0rjN7MDJM6gCIyFM
5zl0pCq5qcGIKRjOmiHW/ebz8En3xAFeweTi75oioOJc1QGQFHpEMOy/DFy2Nm2WHNqulun/oIcq
3NfApqqd32Lv9YPZzhrLv8tv+C/8/5UtbQ7xAwK5fxgMbq0d8Xhre214uS5OgAParDlHfvDI4WEu
nqBCQwomEAjuFBaHq8VlV8VvpN+ouvE7/i9SyCEWfz/zoFFztPHKmfSozjADMIgMtzrIiTQD/wfE
wFUdY5UbZ4fpce18Bm7lKQM5s7ccko3CCbF5moC+CdyMaq83Z4WBHzWBrbli+BoYdAx9CvHdZlls
TAe4YN5W7ZKaW7UMcSV6lELyJmYUbO5ZH0LlTng3lkHDHRXhEO4Ymm9o7JYVxeLNvCdb9U10hlyq
Haevswn6Db/oX/yNyur9NGcWHjf1JPQpMvRcZXqhQu1bmTb8VzmNnlbPp3mJnpSfwixzHkuiHWH8
LK4Ch35Rlu6pnWEENbxvsA/aZRKZmUr1hTnn+Jh9DHkrNJgg2tRkPUtieEcjRp6TIVYKqHHFob9F
IAu7UerOdjOZQ1nF2G58K+pa8AyjUHskqki+bHAEpp+rfzk04TmGPi00mOnrPcbfeoER5HskMZ1t
h38naduHET9Hoq4RsV1xeo1IukFc+DqmR7L+kpRIZktdxDUd23pY1LvbrG7Gh2px2y4Zs61SZSNE
ziFVjDHTgt3U2kgBMApqmnEokUgAL3OtVLXfj08ffYGnE+Qf+68dGrKvXsCqEEgIUbc18VovrqW0
qEx5Td176xoudMTLB77w8CXGUwtBx1x0U2sVNP2uV0fWh9zFIOLtvJu1wMVRkYrrB4PYM9RkizTl
vnknaASgQTjAJKsTd3EkjfTTKXD+/UxnELEPRgDd6soJF7LYql7wtczW2aQ0zWVD41DsCCtdUPfy
HOdg0lG6FGlq5o1SnHiBbYvIYDySqewXgjLWbhTFgNhaaNgRo2rMwdf8ZvQEyrK/QVwx3eRMQlxE
3xH6KL+laxRJxhUPmATGjwynHLw6Z9E2fu9Cf/xzfBussfRrH+upbnkm5QX9l7R3Aq0aInRXnfTm
ZfIzYKvzmPQOQkP+wzUexAoJh+K7FNR7FIG4GCY9zmVT2YOtWgoOIbOcqDd36erB0BGD51QCeWpE
O/FBjQjbnvc4qXudyvbnfQmIlGPMmJUt3FJg+Rp0mim4hhSLvBBWo2z/RKUbqd+9FvVBwfqEw5QO
kKpoOWHPGZi9pma8QWaHOvMEYX03lr5AVOY01rRj1XNy5yQxmgJNMLE+7+nDgHlZVFhy7L5Ptiw2
sqnLrmxepD5l6lhJpm00NSsH8/mxKJtyUDpKeJR0DrWdHlPdoRxomR5sOoJ5ufnlswQ4QIID1qDR
BHu3IYhM0ImwLQY7B4QkLCVbGgTzsnCXhEx230eKOQDuY4LCU89bRMFCzr80FNnINsC+GJyFyjkq
l5FQyqO8Gw91taRqcCHl7fcVOaxpzQWQnBaGXaDbGpLIyESSquFqnJfWqn3Qtfs7772X0C/vd7Zq
QmLb3aFZDN4HlK+YqLaLTP30RJW+sCr7HfB+QwjsuDG6uns5gr41qS6+lFKANt7DljGSvGWGC2Ks
qVP/Vyrc2cJCklT5DvRhh7RzFLSKGcOH4gvTx/2DiTUEwpik9kbTDebDZyCmOPdREBuS9QzKZLyu
u7ByzhEt9vbxlu8ES9HOlch48vm2lSwxMemV92zE1eyxLqHgQztZyr0OBbAq4UtJuXraO7Anm3e0
avZO5MBi4z/y5VUT3WJr8XWpGTzdO6QE9CZNkcpVM+JItEBevxnS60stKxc2/CmZL6qDjN5riV0f
3FWvBtpiW1Pqx43g4tKbwB8G8q2xFq0YJCGLf/vZT9xvuBd77Bgo/jYPNjwExZ1AsDiGSEgfajcD
4DjUIUVmGy+Q6X44uxz3kjigeFHwHgemvAdDEVuEfkr1tbPIokK4Xevv/QsR8xSf7uX6s9JLV3TQ
3vTq0u53J0tLyJ+zvTAkFMimZHPc51zpKewGgGHqb649cn9eB50lbgCf2NNfp+M9sDuu46fzGVyj
tvbYniEwo4tQGrb8Fxj4+IFNWsx5/tfFyqz0dxKhE3mpigvtlWkq5U9y/ds07ZFYVpDR1TIS9XH+
vv+SQzgLZjKcbCnWKDCnO6vYt+j+YYPsEC+7Y84xjLwDwuJ7UKcDz8GutK9h/joSCiTKDSe5WLb2
fYJMBeFvBm2KS0i14sTQRvwcPsv1H0enaXCe4HfjqHMLGzgpPe1GRLex/UMWKMKyEAmI8mOB02Dh
tEwv5gxHSPZxPwykFkNfQtlCbR7laZxMM4Zdo0mk9p0T2dc1MKFXTjxuO6EDgsPNRCx6CqHMl/Ao
FIEQKVdTyJFSEA+DzdLWaZO+qv14FQbeB06nDbfv0XUSz08ojqL6n4vV4m+C2aqmHA9jUHp1DvGQ
k+sjqjDSsQQeVW+ixX9XR7Ls26TRlTEAJXHHDLPvxJ87R4Z/rTFvehZie0NHX4riEATuk2i7hAbS
6CODsl0lRIGS4acY2mSQWkdaaOI0Mrwmiv1CvjugYgHE4vmGR5kkfJFI40leMDWZ7lQtskoH/eMV
O07LxTk4n1RVTwZCQiPI8f0JR8OAqf3dAuXJHJO8QPcUCV+GVm7LaluG1gA68HTnY/dfU9+9PNjZ
RsWn8vZFv4aB2cxfxo/4xJwcLBxF7V+AHCoKKFRnKDm1VcJkLuTr4HhuI7yeaxgPfisnefjETFp1
bm9yZTeqmRViUoUirtevZARER1SMSLIxrfL5UR5FrGd8MV604uR0Cfxja724IaFCfYC+s2toBWwP
jjcY8cFiGj2SgZ1ftFKALQLlu4/YivHjip44XSlo862eEBD9c9jHVjX9myx/Eog3vJMBE1I7g3VG
+2NE6SIBXdvGsaV0+dJHi2lCQCtq+UlMkCcKg9nl5AMVQTJCbA5d8SvBOgFwz8SqW7KoRBQEXaEv
HcrBaZwqexv7XdzJBvCWIqWH7WLP+ZdBhj4PLVP0P8bU2mXz7/E5kn8pM/YwVTAIVl/cbx9tHeFe
3RMOyVoxtUC0+6b+J5wzy+XX1DqYZ2bxsheNrnYT3Enep48U89GhpzOT4Yb/VjXWztgKQFl9KkQh
8gTQBPk8/LuLwv/jq3o2KpMtmaRDnpgEBx9VFtVRfFFqBsBOlJ+YGV0gFcbhQX+lUlXgZM+nrKA2
6q5XCuVwOepaEO+S7KY1coerIqEqTw+miU/GykFAnZTKqz97PYU320xqYrwEV+5ejWoEoHnKUhvN
WmW1we7uHifeX1Y4ai6yIOyjYamhxAnevaKMjCmc41QXJMceXuDNBlwKtRloOWp5/uGgr5nbxXV9
jBHj2C95uWzR10B6SG2w9ngvvwNjPLebc0J/h0qLGHWCUZNGT2DBg/4PuIEJE+D801HZB6XNHGWk
8FblDWbyEvoUzs9SuTUorO2ImN+6skRg1AubONOYyuL92zoZJC29bhxkug8idLKdV2csrivh7YAv
Ts8O6DxFOXLB+MJDKUEuhWHXLEoFDn6IvpNfJSwqf790LZC1ZrDi8DGd4iMNgE7b1MMjV6ksgq9B
f1hsExvBUZpiASMEhMWPklKrFiY1BViXz6HwB9GStbLibXhQD2Z2OvrWMbXXED6Q1tgStBZUtZTC
rVcmd6yx5yPryZE4R2u5SFLDiM1LPmgsru+X6khU7A5HobMJ2R8QPixbUMTFzlOBbi56NpZ+HvDO
cv3dqYmBoSxxciIH6pglnvb8LvbmUin/AMtRCxsawCu4L7aBfydZaoy7AkyPCkpj83B2fFPo/nmR
4Yf8z/wVSM3XMkw9b87WiPrz1qS5H1b0m3hQ4qe2c78xNG8P/rNN3Wtrs6fgnjWSBuCP25KajiC7
6VmZpmKeQrpCbDXFArJichZfEqnuO8CcQdAZ4skTS/aXVMWLxq6FR+0Ho0Y3v/7sHjE5FSr+QcmP
02efg7oYcXn4ZHExw5JRe/23RonDh4jfJxrtZw5e9S55a4G5xworK3fpZUZyE0vDScB+mbyPQnS1
7jsQNeqBopLdZL1S5AioB0Xbn6HtKSvd5HJr0Vtqy2MhjfYFfdiUPnWRnnXXgf7Mgo+myf1NcpRq
Djk2XeX29tL4EkQ/gG17JuA1A2QrBQlpp8M9YJc5gOc6m/Kxca4GK14FwwtmIGNBDsOSN0BEgPm2
hMrvuM6UrUD+zuKRGOsIElsrwE0aJZm50cPfvUCl0GUS40PRyUIAaOnzjo2j/rUn4mfFYiEN6mz0
2hRU337NIEiXMQ8faHk5m795Onu9gppRImucmGTbu77rMmOQ0P/lGmYU8lZ1CiyX16DHJhTIF6PN
7hXV0hXyrTq+iXYwxK4UPPHNTwynU5iaNjdJQm60YoW/s7OhfXIYoL1FHdII8ZspkT3fpV572cU5
9f5EgeQ/Gz1g8oWrzamEmEFcnhBBHqBiRQq0Q283tUX4YvaprMlYaB1PRlLzBaGkrnBvBgSWC6v8
AD9IwQLS0CMdlp9et1FtOHGBGT6m8qm8FmLzeCwzNsZ3sArQ75hzCv3Bexw8VblGsZ/pr+lJwNor
Fl/en9LBjRl6feODkgXn0XI+nV6M3jie+FMv2LXFQk2D1/fG2OlKxHUTj4BGqEDhHc1OTAik8xAp
pR7KHFkAHcawSa/yxkm3X7zUrm8BTi0KBQqf7UdRp6ZQ9qE4wbBWEfhi5A9WElZnUJeELTwXABh7
ONZNcKbtH2czssmMFOrzRHJAbYC33xi8Vi2PMRwZnlBXsMSmdbQolPoBO2MYRKouG1Qd9fXBKzaH
t53mRkytBbN6kNZBEWkkAjir7eSZcTtJRqCDdcDMBS644KpoCIoBYIos0qWPNjE1e1WnTbEIx39D
FIU1ftd9VQ9Gw81FjmzMb/CIfdfbdiML4lrTSk5DuFuAkco79LYOOjlR/v7qVNDHIpj79qM8D6fM
vKBGdmEA8JsakYBt4J4xV9UUEZgqwFVAkWHk7DcSwXZrCZRIgGel7kTCyHm9huAnDBUaQpvvock7
S9c87XPniGX0vznI6NbxaFJvbSBYiyyKZ77gsbHNCED1GwEbdX1CCUDkdalOUAmyitJbucbuggbc
gLPFxobetcZf2qseCpgrwv4GrZ0z2wVizp/XnWnYzw0CEbthIy2kRBzLlJ1qySNc5YE4usqiZVHp
MjAbt8TB9Lef/ZSsPYWJB8FA7410GdS4os60aqNK36MunPQ8E39AAAi0y6YU+GRZb6JYmojdHHje
jD+gIBqHs1i1IoOJv9gEaaZvv8S71IC8qxLSLt3kJAvvOxCkV/LcZehj8EyuLNEFwj9ANHyy7LEV
rfW2IhwuT5LH/hERjFuwjT41STEKvM1ts9mLjLIyOzJvYDgYhTCB7VV9dagyutl9CuTtYK+ysoyU
jD103a3kYn5tjLIub/fy8hrDFSdCiYSgMQskiHlAsZ1ulufT/yRlVikbhkMtPb9ZDXXf2GEV/iQp
LUekiC4k6n2QWrSW9j5UxGInKip0TVCtM39fT7BXoVkTfx8nJ5QE8r4qZLwHg7kvD0FuERVABOy4
vnSf7PgKciPKeaLpxlrhFWgYqiKzof5/bFMb+vjcy0O9MIrrnQE5C+oY+OrTdpFKYpmkFa1vWuyB
2s2D6Z/NsCQpjPrzl8npKUXgy+A5hU0oKGIkXIdafPuM+aGT5f9ckSD2XDm+pFHVlJFYeI8BwssM
s0b+JAMDBUq+81dXYyMzjfC7gKNzC5WJmsyT4mGe9KXtQri7yFCEGM4i4+5QS69gdGr9nG2NS+d6
6OephJkb0Ixd8P5rTcWrLuOl0u09XRgJdhkAK6aROYO5lL1YzR2kY847ZnZCWnb16VN0H8PH9Qe+
FVRiaJKI1TxqXLhY/IQuoWtwUfgxh7UwfNzFD/3fDTgCFB/Ns2TZ2okCRoXFLHpw1EYad2eQCt6s
TyleBASVbDNedfbf0JEaVrllaVQc3JsTtyXCfGj7hYILLKnxEWF/OxOWRXhhXe8nivQHW4qo1pL9
JvO2tPn+SsTSQGLzdxHJ6ymXpA+FtjjXhvPV+vSkR/K2ukdW5ZILkH4eGDKuaa6bPU9gzkZELxXl
f9i/xgbXLI1BPrykgqkRdrAPwkqY1MP1dtMjzpJ8T8PRRidHncU4QPpeQ31mJzQ0RHprY7VH3KAZ
hpF67tE4qRl/bT1kKSKjQqBT+EfALMPcAfocV85aX3SBUlmA2wPz/zj3LbG5tQC+qg2g8CA0Czjx
1rjdIvGI0lqznRNmbDLoOOt0d2yReFwkVs6f7bQG0JAsevBd5QH+J1ZLbeuj+N3MbIy26T1g525V
8pFWWyQ3FI5HIErHaTQTE0AUY79Wukf0Y+BNAVFeUtVElPse2/j3q0gfMg3HxlfExIF/X4QO4wk1
v+kkpjMQZUQLIqeA1cJyDXkRK95L1YBWyRp6mqACsb3ksS/yQnwDKe50U5y5IwmGFMWJCdik1uFx
rwrQvj40bte+DR0UEltc5cu76mJ/EmThZHpmnaXtIHEB76vgZFt/N49P1cxZtpIrfQDjJ9vngZCC
8ZMWpsbCOLm2zlumyNIW0U6D/n2CdCK1uEsBYOrzXMxC12PXGqcb0FKK3gB1NxTCB+2kW+yOQ/3Z
w23vLqTql0HwA9tjPicCaEKJ462LXD2V+pPi1C6lBxeycl2VC9Al5KYsr/OES/S5xNuto3kiZlCO
MrJgkqJQGhmXvTgbBDXAal1D0r+7JPSMzYbveW921+ygCvUyrDCXGivdjYDf52CaQBHgJabSnhgn
GAax3h7aWsl7FlQCwS2mxTOnc/eeX9A8ev/wokcWsCK4R3AOPYEcO0f2D8d/ETi83rpab8jeXBIP
vKFhj67ubKNCBLRZW6yNfk8JYH977aC3J6baCBeWELUEYgz+8GrHz6z/YAxFYXimVPLEEARaW0aW
gD9MlYR/cQWy4DFCRhHLC7qdFPO2GBTsl1bRYOv05u8xgFv2VFo3NMbAnIO2YRpNqIVBcJOGxmRv
hheJsIxYfAbKDHFvX/qfeBb7B9JvmJUp2ZKdzhfFqHCSvINlGyf3w/MZzXG32HcQ9mV056B9Os6y
jZfndio7Wra8DqJlksFrR8GV25JlmDcNFfZaqRI+uQd6sXM/gtIWxSfOPQ9bHj4WusbQYjX3iDIC
RxpVnqEZZJCfsNziYXju2GX6NzPttDz8x3KM6STGKvU2I0i+pvAwaCtpXYqaer3/pQE4egRqAeM6
kbLF85OA0K+n/UOPJ00vruy7NyQXRE8Os4e+ML5jOp/y1o/+AvB6jBSPIWHRw/ydgG2iudXYgQo7
rknrTmK0Qj9PO6EOc3DQYd2r54r+Rbk5+B0q67zaeN/2E5gsPj3MXrSLpTaqVRRqDfWX8TiOM5kx
XWo3jZ1M0VbzcA1tqGN+jWFeeccCiJBfbPJLxaITknDkxucGBmXPqhabgajfOL8Nt/PEIe1uGDJu
nJ94FJ5G67HZUAOYUnp15GhYCq4HIiVI3RMhCNisteWgtjyCCsktrPu0WRzaPsWws0Uw8IBeYu68
M4oxvN2TR3SEt3Wuv50/+lSTW4P7nBT+0FfJKCwo3jKi9y3qNqB4gI3uY9xP4X8nrYMfBbaJ7ecD
Bepf4BcXICRfDUNF0zVjlGbL0awkAB/Wc+VSZ8eG0FTAW+/HGP3TWNF+vjN0wP9hRiGNuXTG5yVK
N9sFXG8kV/sF1i1kKe6llDohgtfQC9JNYLc7BOgCY/jdajqv11p8jnsMvJaVY3ikH81GxF6sRkgX
7SFrfTCRG3INF5iNfpCmYuw9jZena5Eaoz2Fvqv/dHy2Pq1d2GJGJJCKvBWgnPP9oitTI7o/nlc2
eQLvEi/zEDdfq3kEyKuaiFlQktFmIIVLcHzne91ysi+Unfn3laky9Rca0PqxL4bYt5iyO6G9Gdz7
vUK6usRDeow8CJ9s5xF9m5BxzNA64CxGlZ3Y4YC9JYadzdaI364YhjnZOjDk7GlrmN4/oBF1SlBm
mWcW+mNmV6xccq5ybSc+lMIrnGY92WZNBQIQxQZ8btWogAmbvXifndkurJBBlm/zQmDt+ciG4D8q
axgJoexuSmYw207/PRj+4MrV3kTtJVbXOuiIFG1YqZ7i+W2Dyw/oSXpGACIcYz50HKO/li71U7hK
ZzwWxh8eKfFX3XUThcshAqQVKcdBG1cBk5vo0drwqFeycBdziQAQmlVqyU+AInQ3A1k8HKQQXFeM
SLqReqHsELPfMNh+KglUw1+7a58cSkxJgyP2HnK/yiAmWlTKB+eX++uVMbUi71Hsd+084QcqyLF2
VZtmBuGo33xwUxu5m0j/8o74Hr9eSecOZtump6bv9hIWzskLE5qiNPGiX6BkTC0bVVtIMpO/tghh
OR723n/Czah1VSFXku3Vie9UCtrLjBXKm7hlyJ21oMCeV0jNn+C9xIB60nee2d/DfMsWXdpoXyjT
hBO8wGTX078qvCUFKvpCG1VnDQxv74HDM09ep8MnCJ4gNFxDkc6POmLUwNpS419SP6a8u9g4VHze
YDVNHCRgxZlvvu/A1rQR/SjliR2hSPY8Ux5Ia6aPzbVdjJ6fWgOpuOVsysyzockms3CACA2Pmw3o
rnd/bdAFNC7Bv+z5bNZx/XAfojuNtD4HNfyjxjpkaoOxOdn2dSd8mtexF8XwQXz283xHf41iMEex
0VEm+JVlWL/fcQFlkrW4nbMuqTjhoco72TpLFO7rG61IVIa6OV4n03ASiBNmRgMvtIbTJJe28Txk
gukfk+CewO8ku9X2VR5rL/raYiRXJKSK54daqkVmj68jQV/x0p3pIuNC7a5Gf59Um283sVC0obpP
5w7HbPFga4FlJ3583emBHq3ma/G9CmQYHSD/GxLC6/cXeSMbD4srM4MshYplQ4geFMva8OO43wkV
VekzSg4ZcJrwDIJKDOeSjxfLI1oqnitDMiJQcdIghtQDtg0PyFcSL+Rxt1Zg9NYASveSEMdaDcyb
8eCnZz1LfiSbX/Prs8Evp1E6GKiU09E9Y+nmd17uU+tw9IC9v+A6wFp4K2CaQvUa9QmP6/CjK4x4
ZWREHirdh3nnFWFhcOdZLH3jEEDe5cn56pEMiT/JxtHOy5gDS+EwJe8nwzv4Du7rYkAau1CZCiUR
A3ZBkdkEOlEnUEJ0O1iIxbYDZZoTRcu7WXK5XPMc5UfnHjLUZra6O7jjNen94Ya+pv8AViscU3/m
GJNTL+c2M4GHzMyc8EInPKP26+ri//B3kJipzc5gT2nvcAnmWf7TdhJxl1GmH8SHi/caIM6l+94H
pfENv42pVXosvbqwtQhQSqPOir4/vCLHRZzG+knsc4/cgKbRMo/RMm4GCm3iqOva+R7XH0W9cilo
djlGMv85VSvYoo53h4reknb6HFBnzHJ9lydw90pVnRPiWEfiN8VEw9kfKMXJ1Vqg50c5v1JKVIUu
LZI/YoRcbvnvA8nxKpobXgRFF2w5bkqXLhH1QR3ORFnSxJ59b0JzipSUk6YuFY2+VGmtAce6/HX8
cd/61uOSpiDUSFGNuJ25yr4JDXlEwG6mZuLUFf3i97LLE73bMZ2JWKejmm+RJP0gka1kbi2DT70z
vMAfZBEFtshgPKZKhVwuwPkHUMyh10NnnNwq226lZpgTmEWpZsZErel6Kole/bJ/1fLrA54ZxAQZ
g9OuvWUNLGpDeJpGTqVA7mqO1zwGXaiukMRXvcBcIqtlpLXnGTPa9CfmJDTTP8DRX8Aq1DPz/k9t
vL52//3Vw+M9xYF/Qz5QpKKEmXoxb4fmluA53X3XUtnDQL//I4plQdxEBMk30Q7y6Ejf5MFcGJfX
Y+RhcljsyBVtHIx5KQPHkb/GXDa6rN78tF//DUKRRf3nC/SYd5A2EDIFLV/LrsU0wlfMtiu+jG2z
+9nOKe4/h/LeYaKQZcIxFk6MRQd++vYZi+qX3Lu1ryO11spZLrkN9KZgObmaR58xroBnWD7QP5cV
7Dwr/E8M216SXksqQzHtT/l1GNCXA08kxLT+ZFBiDyHRqOIrYJkaKikLKbQWP2EiAoX6o4tfjVCB
SRH6mHRzEnlMsGBpogyAtlT4QP15wMOfUASaiQdXrpNy7GVW5RmNFutSGk+C/J9wu9TZ9NP/uDlH
78cSBHkKoeDGOj5S0ydN/qCj3vGYlYR2CJz9kVtjgiGJc8m735XuRe+87g2o3pZN+R9mgKTN9A9j
SvzOnPUKAwy8uoTqmp2CKZlB0fRpsvRGlh81NGh+QCR0iOx+5bwtjueUb52H3XlXs8SHFaHwR76b
5CBR1hJCLzzO42+7Pfq/XZVJy6VCvO370Ex8PW+L0sE2LtDVzv/RGPvkLmZd2IwWAwr7H5NSHpE3
kEisDSDwoXl1nFw/5hziZWN+LidaC7wCE1ueaXQrZ7I/IvOmnjfJ0aCCjP3pfrFzhZ3NotIxvBHs
ZhNDLjPS7r53lb6sy8N13LlJqZvAwaVt5HaKlm68vS84h44EE5SK7w+UPUWYpXEBN87LLjqFPvcB
VZmxrmOnKBRJCpM+URZ0eYfMSJDcPQra+DQCHhYlnu+rLCaUSpjtpm2S3pWdWA5qaKq9Zo4/kx4x
DyKQ8MKYd+a4xG009QuoLviZr3PLl5fpCBG+GxD97pZN2oLepOENWZytOD+05ajzM1T5k85+obEm
TZqUn9SBnVTNBg9jkVqKg7lBb1uMBR9UgPtxt9QFNDOlyrr2fBcrFiZygDGNglvkd2xB0WJcaPtv
cwwdg4+TdsXHWDN4eyJHOX/jJeBWKqngrKuGfiYPXPaMcjg1PoXZxmp2TET9rXcipUQVMFbVm6Cd
87tgrPGrpfAIIjtBY0DrFGNjCJa8BQWa9ZOy2EjyU4wR9F4ROA9f9fWY7KNfIeoQjrxmyjVnHeNC
jzWbAgxzeczI/BguV1ANRTF4XBc/i7L83N20/e0H0nOeZQylFi8Bg3z3qvsWFdq2wwymB6Luh5dB
vuGMzT2mk1MXmT0b6iS8gVe9zwCN1sHVUZybeGL4Cb4tjckqlfHQ97dxWJtvQVjxaWVMT12Dc6DB
6/nLYlkEhVOinTKzOq65WoJGWwncJ/+glAk/OIQahbSYZup9Qtb7ltFeIoxkjLXPWmBDmU2y91iC
QcTWXRsQmk0XW2SZMCXemeUD+z3t4I38bXOHJbF34+e5i24ACP3v6rNd1mPEh35Yap/0QCc2DH54
Rkh9BsT3hBEyoRiHEnRPMjgp1B4+8CbFgRZvW6oUWXG6aJXuZ6REZPHkTaDtc0AZXeMw3BUWnfZU
9HQN84APvsX0c0v9mSAhR572Gt8QFkoGwtbUljVfGiCVo9IBue0WIYuFuZAJVWKTv9r/ZgBA1SKg
6fUJmmISyxoVo61QiXv2T/fIEpozoWKATfMwvriKWhqyDTWnOBn2IU9aLuAKMY/QPiXP9ToXKw5I
h8oqwr25MLRYGtLfnSJTe4mWnfLbjLmQDPxmErbGycsLWx5AoCU2898icYh5tshnSsPd71GGg/kN
I45UG9jDjO20oBC6J42u24gOBuB/7/EO4s+VhPpegm4/BNztAwts3U7qhgZt5LB20iIY6ZDMCa91
49HTlC0wKMas4+v1ldxDVRQfOYZjDWFMXManc7aXBLVwd5UquS6YuAHTnuTG3Zb9ME5jGxcvQLu8
ycVqAANT5M1bbbMXIGJxWhcCVMM3cZiYvxtC0Efe240YcE/SBdk8dfCeVKbGbOvJ9iXJrxqF7ARy
9A8bWHWw5QmgDvVxyjhJ4/f8nhJZhGi8EByUgU2rYL6J9nYouIl4BgpDArEkvpehaZ+Ba8+bzLIM
qLkrm21p3fzp7mKCHU6zIGhVCkzuiCTDs4TGe6wUoDAYK3wE46QjzHbyzOCC1bCVvhDdyn1pIh9L
5+jvX/veFwbI57TX/yf8KKhSwPL4G/e1gWxivf0bYvXctmUROSNNh/EIOun4gKOeGt/TmtsDs3px
EH88a+LRzMtlJZOY/YhhCRMd1NYJZWZgoacDMyit3lyCmRazOLjcCMWv3VKesMU95kH6l8HYFvdl
7W/VN2bIAO+w54aB3BgYpYArt+02UPu7U8lhZthnIvAAl94YZVva6+576tgrkIZOV0aoQY0xKvcw
ByGwCX5jpL/bOixcS4LK2zuITNBPIRUz4G+jPv46ik8IuAOp9IpK4cIUeLZH9rJMqJCNzjAAKqQi
THtoTe2EtqRy+eeXGPk7wBZcSC4cGKGClbSpavuGc7m0OVHPNotsX4bc3f8S+L/oPLb14YVs4fac
1xESF0pwijPLNIJAOLdSXR//pT1RmLUjdlRe5ItSF0l+XyI2RHDuALOAG5zu1n6OrCxFXrJhuACR
3KF4IBhsUh1366K4UMW+i/ZEFGgB0ap3Jsk3p+2oM1SyQZzpS8cPoHM+v7xCPaXrDTLZum84J5E/
vloNOtgHU/lgv3U5uGKLnJaHzRUd55ovc9MGckMkwGgIKpkOj9ddOcycawa/KnnjDdwXXl6Zrvih
dRL7d92MREzleTHnycartZa+AWzQYIQs/JdPgeMJjGnxZtpSyHwgv8l7h31TrFTRgsR1LynEUOiS
ur9pI4pcewrwdptPNkOYOQMxjt4rvj36Z/BMv4NQI2wQ/MeQguehyW8PL/rc9bfSF9+RFKkXq4WC
mPxsxl51uDpic4REHArZM6iPuPnNXArdNYM05ytAIRkQHLxE1k0DgWtng/JOQslcJKcsOZQxWlTe
dlp7u08299AY/BJCa+6k7zjtXT2CRpba9rS0YpJCwf/A4YD3ULq0KQMYJxW0yl5InIt9d1U66gYy
kTBWdU4EdBUPTK9BL3PhqGwGxXYHvBHIW24XjUakQN0pZ0IH6jAQECmcSKQuamFTg4w2HaHGKQkB
ny9kMsCSl+Jh39+yJ2MntJIzmvuN/D6aGSywg1NtqZMYfZ191b+RZd08/Bk/zGu6oNkrDYqZ6D4s
HQMTEQuu2TK78sTw5vV/YIoMJVbsVp6LTihV5rMMrK6GBw1L421hXYLhmtWVlgJxzHIaXzbSDggW
QmuJzp8uVG0iOvZ+vsU8Q2hzRL3X6RqtzbSfXEB1fiy76T2d2sZcxqv6K71yRth8InvC58eMhpIA
mjA+pyPZTo+r9PiPXOpGaJsebVrSqmfBm8cAqEu9FSCX0uzBk4nS1lza8xqtWL6sguB4jhC3bAA7
N+KO/8mar/gjMxM3GTuQUH96inlFm4yK2pSjEw0ahiHUIHqe0ufb0GFcAAV5JovXo5qHlJ1c2cci
Kw+yZDY6AEa/l4LQes0F6IE4RMlZyLqQwV0z9zGDPcPiP9hvy5Hg5jwHIG7ZtDlHnh9SgEoTnFRD
jnoYfzGdpoAtoMSxdSgcwuLI6OR3hVC8eq4JCrozPoc6pGL2d9sgGII9MP0qv59oEv52KYZ/wdGc
kuDw/UaUVmzRWl6E2k6VnwVqK1cmzfwqgbR46BdvURW+XQNFYAFIN970ySATnodNyl9xBwiLmmGJ
QrH/KlIFh5HVHOPNyIhlwgPjQGJbQh0OyG4/+h3tdNiZX+pc+57OAOS07MEIDHABstpQhI82W+Ms
9ktrTFZbNI62S4SuOuWK0W5/iTixYx/9+8ahjLUZ/alQ9uHHk/yLaQ7xOnOw7R3mYmBqwjhpg62q
ItNgIHx0xNRuoykgP2o8VOCk6fVVDOacadLLOZuznhl9aXs3NCSo7K3wQkyc44ObQucrS/TAM6XD
dTPJhuTLe4sxTPH6imjcVKJOPGbsSL11wIdKEajpqJNcBgNc62sbtgopoetxNERVZG/lpycTQLkF
Zng/Bu4IeLgg93FxVzLi37bqVhhveQS9upxEUtUtTHwMchUgnCyjs5IkY7MTnOAqUNzHfOQJ+SX1
Lj6qzonFf2tD7XcFbD4uOdZ06DMLTOuVayQWaIb4aHhr5ike097o5Sg/95Ir0is4EiRcvxX9q1FZ
FsYG9wELuklpEne5u6na2rCn/AwKNl1ln2d5qCSw8IlGObdaa34RvOnYhJWsm0iqDJClEf1Dcq5k
5SGq9eJCbqvLoANi4aX3mSpbzY+RCK+Gwux8wDeFyCpdYuYT4oy74GvxZyx0G/iP3lPcRRCl4eT/
uJr/k2d3orEYtRXyzr2hY7qUvRmeEQMzHiqyAT2dHekNEjH3e4IPaOpqEJtZPJUpc7yK+OE8Ohi8
KCPJaULvjdMt8nVXj5qoLCFhlsq/PojQMTba7TIsBfeP3QKTURyP5zicWLxHaSopf1amMjkTiDcM
8gGF2GX7ZwfSTN/TL/ecTIlTme7bvT9Itqms2ql7Z0lcoiM8Mh7LBraW6kiRhr3hhanPLlrQx5N0
D+xD7oCQvqYzYzMeP0f9ABhI1xAKqSDmahs/H8VIiZs9Wemuf+VBYiUMkOOITuRa0jI/zbHoonNK
hvB7BmsjdVt57DUkwgwLov7dHw2m1qWD5JHA93Lx28K2Uv8yLTLH+IbPaJc55UOldfqnzpA/022o
tJIyYn3usoiQSMEjyOJmcGbgaYG0CL/ZR4H4RiBH75DFPIHdZyAwldkVnERBJzncB+2KXwS1GWD4
d7WmRFlks29dr1Xhn07iSgE3ntWtJrClVZ5Ey166t3VKr5xNN30QvFEFtxj/SDJDwtDIUHtEyAwx
AXg6ZNE6+gC/XCqhLo765EJFPYYUi7slDsQ7B1GRDxJos2cqU6OHeF20na3s7TU/9EkA64Om+kDc
hgXMiC+StfnwFnkBguZso9ITitQtSFhfAbOXItAPv/5PubkeBkazg0B8sUJSTMaS17tCtBa6AcCY
uRIDSiE1tDKYGDn/EviZemdFhCzLiL8D7n3Op/Qm5wjw3y6jGgdpszSpeugTYyBWRwtzh2UU7rzX
UsyXbgxS1+RJxY9KEJ/sxtsWKGMPL0Ig7tx626VOsCEs1YKYIC4fbDGQpKe+GeIi9LLN7ziKwKHl
a/SFShDp0aAYe2UMPQie0R0/UoA/7Bsk2MX2B8r+NI57FmBsx95x+Kc2xrqvrSRYbZ+XUBwlxwgJ
ySwNcXmMyqXPYhBqC688WFSbrkTWy+FVEgZLsuMzFN78eCylJxtbS46q60873r98Wmin7e8zJhb0
CewvvAn4FZnMFODJZSTNAhKzMp4JegRcqKPw0JXqFDpqiJ/Nf3BDSBcqBirRnakIRxJ77UnK5TH/
Y3e6l0P2fRbFmg+bkvh9jJAn08s1MP4GfqJ5HE6P0KkrJmr1rjlUduNQInvROVxUYUhpiM8cFJEQ
VXScTj2hHJ5jgUXl6MpUWcj+WlySLBo6kZOL3Z1tzt6hoHGGXD0+0d3PUsuBiNw45vIYa3jCMAyF
y7QatdV/VtKMjiUCf0zmt9/Awyo9Jo7RH4HdmXlesnB49IihULvCZy+2WYMDeiiirj6mWYcWV10e
cOovjUjspx6Lf/ptxNGv8tKbLX0BCCOK1/iCzjI3Y6I/RK+mgKZHpcXJb69m9R/qcFdczruA31q/
Ieg2q/6lXa3mssDas20zYJtn7jRWMHA/A2R5TELHOyS1ZvgO+t8zW05v5yzimoERAj8t0XJyE+LA
wqrOCGGiY1Pv+UIcBRWTFpchS8JLogp/oSIsjQY5nFCNT4qA8bBJ7U7xrH6qTXIfEMoNNNKQZnqs
PsIc3GmbtjWeIi0Cw7N0Z4jL/phr3pGipi+5U3l43lmJ6UQ24UYn7yfbIvwfxRA9gohM0uSd9SLG
KMTR8O8aMAy7ZijTU18T+8GeWXIcg49R0xAl5Ctpkw6eFhGLKqKd0TwghIxjuMfj6MYN3gXYrWvV
i1sy2IJf05ofaQ1a8aNAWnjUDtnA2uGqmwxexXJn4hXDmoBse5HeTf+vrKMwrvyqKS+N2J/Ye46x
MAGODT+SncRZNX5BMRA5W9K+B6c+ox8AOhPkL1CNDKctAbMwUx13EjGkvO8/Uu4RS2WkfB9Snl1I
vJAdRheiRFNt1m/iYRdwttbbifstOfwB686vQb8StemjgjTxvFEKP4zthTPJBlymmu8pQvKKuiqo
L5JFndBIjZSUfvPrpCCI9wv4/4aCnMxy0Zj8ETpKVEih2xwGH/zvrQmtcr/afQxGWPf1jIiYyZjE
vF3racy10N8Oi/VU5REpt2aOE5spMNyX2r7xWD21VRPMU9ddnQTQhRuc34duDwHTMJGvc5izEmXA
J4Kdg2dnVfelHvqhK2WckolQB6zbM9g0VrRIGdFV9XTBNPfTwdXUIe3a5IfGAZunQ5REG8HgmSzZ
r3uTEnw5DvM3QJebWgYvPDKSpATfYn6mbQVJXaQVryLJZkpLGnGeRPwj9RliZjz+Saj8RE77JYnd
3aZ53/BcsxbZs/wdKJHsZjOWgPe5Nsqpejme60ixpKP4vDBdnPxnakV+YB5WTuslNrfmovH/U6FC
4BvqTghWzzawiaCt1NCv6OrCdxRrq0c4akU5ambwrpiZMPukaIhVEt44XA4rLBzMnEbnXD4Z7brG
rZTDQ2A+0ha79G3/z9j2lw6aOX0QgD+Cv5MU+c+d2bs0o7p6Uo+Mr5T51fxGqC2GcuM3mdBNNUGX
gel0WBUTL1wZEjiUoYRucxJ6c8ZtvxcuBogaWNcNlxzkJhBx25EoU0CbE9wjlZsigMfnpJlV27Mf
QBmEmEuvLiBvQWLKerdCyFPGBa4tz3YySqPT4ocMKDYFbzX8wGXOg9JwdJwB8VmvDZyVuYZVW9em
t4yVVdU8oJ4HyCScJiGHpl7c9RFmi5WiVWvfLnTCPXGB3Nbfu2rBqSTOrBHuGGq9MlpBqRzucST4
XzHihQfCB8Db66dZJpNR+W+1c0lMx1YeCrBtJlxeEnyi+dvSz7I44B/reBylJpxCoZzkbpr5cct7
TtlBzEE/ZMF5O4oNBfAAIRwLzW2sejR+NnSytuv7q+cYwgTIb0/MEGM90+KyKAFoEd+XdfnqCNju
K6g+HievyUisGOpBPUmT8628O8kwGHbdz3odq5B9bY8k8RJF3sPcgYplWH+duew5GBgEMjGnloYV
b6VirbG+LjAHJVD3E9oFHxeS/iZTcNhtrvHGBUJpVL8FND4fkzmT0laDbSxS6cFNXHGqZH9nygTf
4oWlTKDLR1ofsDyDEVd/J+ZsukPfizJD2GruLSuoPh2jfJpaq7VKHymjjCaTNJU4Pi8yozWTua7F
UnNZ/CperzoyiqgZtLm2B+TJGPGkGvRapxC5BjL92q7W5DBdkPaABKL67Nr/DS1awG3UyI7ODdzI
i/xpwPOZ7TZ1RXNEdyaIyOPl3EpfBZ6n1Mdt05eJ2bfqHKLV68H+4IaeF5XIroEEhHba2k1OPMqL
7T8UxoDwWhMSMaPG6Pr2RSaltjsiQ9jmghso1DE+zjOUp0HSsoCLNhOVztHJ+/Q1QGNpOyt0R68+
IWDL3dXR/eMi1ZlG4D8xZyesJiNpcKNLCq5PEQBlGm6xBIAanyCgflmDWD1XIRBZ8zetvf34VsTF
XOT3ZvCVAXsQO4lXkYfpJdNjHh3L5sPaqcNRYOaqmSpEKVzukAVYEBFNzUyPq4/UNginH3yEHMGM
3hNLNnTXDyu5eWcdTxuNUUnYgP9Ilry89s8Oy/eqxPXs+2MAZnteJFAAFmj5Wlwsd+KIU7RawoE6
dLcBmhauQNd9yGX8VmENsEcJINi3m6RPRe8k83XF4dtqWe+aTu64gasooYrao3y4CWumyBc2GGXV
lBdAzKP3CSMw5rrWaoweG+FFlFbxw1ey+YBnbJlUJEFbOyaELSMTx0J4eEvWPANFF3apyVkB9Phe
+kVXjKARNULHSgrMBA6SVU+egSJEiCaPLPDb7d2d9caHKstmdEufF600U5jysU8pa6CV1F/jIAIu
UwxopPKSpefa4yeOq1Rgqy1L42L0HPU+t9rOdD3zv9ZPmj2AmMru8A/SpP5TbGOiwr3w7i8Gnj6T
cAHFqRpXjJD+hGazAnOQObCEXLBmFnvc1vjrdzJyVCoXaywL4ghCnzu4XZOcwMKUBBlOOqcvHHzZ
bNAaPlzgUIYo6KjFni/gyuopVkleQ01Y4nR1jUJtCQASlQT1lYxPpFJzM5ADxPyBuiv5iVubH9UH
mXO/KPlwjh2UNIw3xjpn6q54PJTQhAhlferz/JMj3naSm/RJirpbSdAVRcim93k+otbGOWbN2PHu
1wimHMU/Grb9KbnXy2pUR/d4+ivkKeMIGhBHGSpUmWJFUxoENrW9+xKEMmzP4e23NOWyQ5pg47EQ
Y0XCoz3HITveJx0fMvk+Cv6/z4cvQyyUAIhKqOAnp3ki1sUqwzqUAdAlNWLFijb3UkfhcsXo7Ob1
Jl7hD2wfOIR3rGs0nD4/ZRxBzxgisfCWhdpNJpSHQG2iQWyyoOGjuclp/wKjxITILLJyp8h46fv7
9ViNBVshpwQmfym4JTYlPVKbZ6wgX95YXrIYSl5NRCjD24g1GDBA8+eSgm3NdiTvowGMW3ZTZmwt
WnBFhkIeQJOh+6rzc2VfQWD877IIDOUEiq36TEcteNOSf+2VQBj1jhIwGQvkf+LZojIhkd7IkOhf
UvrRf8FMX0gNmYX1Ga5uJym2rzuUXBeofPvP70KsSJMYjSnH7b0LwztgWI13JyQ0vggRR9Vj246t
T5qXhBDmuL6hGepcKqro7kGCjsR3rZ8oLjKi4B6TUDU6quZG/bUUc5u+bmKK6cfdfj9vPvlqpH8g
8zPn5uLuXOr50sMAoI1SD5AahkLueMNk5IX8V2uDgQtaMwG/ta05rl14du4DzXWHgeJ9NCYWfAQK
rM0J133xvfaNr7mtKxesU3CtEnt9fpb5X6exykiKo1v2KWaF3KLf3FUjYqi7XlR7V4I3mSs7zj+f
xS+o74c2oqRTnDhg/0W8u8XUc3noxf9GhOYgvpdQXb/BWsKPnKrvPOCf0arwrfT03BaP69tyue/g
j+SJxgawzb1Qk9YGfFLKryYq/c7h3lABTsTVYQkdpaMnFuwhIqf21ACo5pVr9VfQD1FoKLWpRcZ9
uOfd0GHogse1OjaczzmpQ3Q273kQjNNfGyrs/aLbOFDfH7lgPrjSM4FMR9b00QNbqSSWxASpkehR
U9//jcU2A6LYq9Tdt+L+kjytGoHv46hlvtU8mwp27+/2+AJUWJ/34hxCQ/8yCxybM/j8n75pDWg9
eC9bNd5J38HnovfPZnwZ9u9Fw7PqHtfRix+8DCYLtQ5FTJ1Re4PbwJmNHV+uvbT4o+I/dAZDfDiK
XPqOe1mVmB3l9ZTeEA9N+NRXt9be3kTzcIqEkA5lXQ3H1vQHf7LAzBN/TnZgMCV9fCdndwSV+tLl
idWOB1P5IGOUZYqMqp+bm/zTbfU0TEWtRFa23ni+F/mSWqtQ5Tpi00ykRQ5WrZS2jpZNsqJc6BQq
k9duGvbVAXMejoFbRe4lNhmHMIvRA8WRm8qsimVUz0zpE9mMRya2qBothnLWNDnMX91K+zPL6bD2
yYjdR1/2tO+OrXr6uEDzLkK3+VYtZBxiDgqS7iHXVsFbZ5gra1IATFln6H/dQXJbnZVpwGQ0zIh9
Bq7gtqU7C/yZFthGZBoxm8gNuZLKagwmu/ejIXjad92OSwgqsLWVjjG0bllG11EsdH7q/dITIHMD
yh8anVnkaeF9PQqv/owFdWg94I4ZMYXkIM8z8xQxkaql20+wQ8V+GnHqZccts9ESz0uiuxqkM56K
rskrAXrlezhezRbJhOcllCS5HOFYeYc8No8gFwaGumsBBOeHI0pM6ZiLUBU8aQ26YfeeVwNBdwY8
wOtacCJfo694jLmbh+v+S47G+4NrSp+dgXbinBqeUh3lE/mxrn0/zEZ51/ypKA5fqMUiueCqEspj
lzfDrK/mndpPfhOUSjXK1A7LJJOZhtF9FONtg83CZQTIuh05HoFpQ6gCF1JdEtsfLalWUKpEB4TL
sJZloqak32yOWHU+dZKRrx8WjGmOTU3PJRePI8ofZcC+oUswiquWjSLeUNA5n80HQFK0/h9wt89x
cHptvUsFvR14s5tUKQupclfXNMir6yNi1etphDurUPHi3zNQK8HcWxpikOhXn6B0oolaZACE1+Pn
+8hjHEua8B/3muLFL0Brc+fD8ZKHDqk/eGpVka6UebqCVw7qH0ynLnuBavtA9xozYQn1PuvhGTFw
T78w72j/fnpOokLAncRocjSKDoxnvpwBVCyTw6bX0rWm9PRlllTAH7slBgOqq6Vr5CM8zZyFs7v0
ADksNt3wFR9pBLImy7Qr55o2t30TURD1lOJIVLsYw06yRj45ejlPpY4D8B8UsgYKmn/gCACfXESh
KZXjlumSBa7Rwf7sesqGu3ThwiNothfqAkeQJjDAD488NdciGlu5u+Kqkm+ryzYPk/b/hAcdHPrV
TJisWb0BzjB5Ewao2GOmKAvw6UPhdpLSYl2pz3YkEOzKxzBR6fWmgeIZvIt4FJdFLAy/wMYR4QKS
cwiagjIUmd5xjKOIIsZ7dF8pf0NjKx9hF95xWo8B3KUYIMAItRP+JB4xUA4KDKP7bBMJUJdGmZ0D
woqzfvEzEhIkwi4IuBaBmAs5fnMRjiy3122t+bZ68rW/ZAxCYMYs0PkFnXz6OQeOQuBa9f2EFPNx
hRV6xkNY75pgMBp2JuD2SytE2EcdnDGdhjwkcjR5muXxVO78P/Qu5RDZQ9t7rYAHUwId4ilLVuTv
RtBVK4TqszS7ovGrVyAeTPEReyTpyztPXMpBEHWR26rzaBc/Lq2sSoOyV33sblAs+w/9C7wzCxw4
+o38L3tfG3fWaHwuTH4+9MetXffgtNZcIqQy69hP0ojkw0JIA61bIKmKy9HaXCihbB2CcoRwHbTO
OgkL/GeXWo3NDzWvaIW8ctjPDkeVI8K4gUtacnLBL+SmpHfRi+RcdiPrV3l51gMspFEujNe7U7Zg
mt4HbY3CBrXONIyX8TubuBpD8LxGyzPD5VLcUn/dLMnzXBtWYcl4qWe8SC7GwxdTem2GLV1b42c4
pm6nblurodC08gmQ42GCePim+m7G/REVsZMkAuINjLHZZKkXkOp2uftvu+Vsrh1MkS1Pi/7Smwlv
c6jY1F3JZhlt40uRJbCMNYCV1xJti4xgKInhoVyrA6TK4UTmM3EO7uDc9J8MlvhAar5jx86HcX0p
Vb/JRRl1N4lPrBNxpYp8+0HHn4w5imvD80ir64robscsthx2eR1PGDsHPbZa/RTpozA9MNvTkR2e
MZXyuWQfVfFByGrq/7txWaXosvqnBv8nvvpj1Db1FJjARQhKcn40iGg+xAHAbeuM7+toj8/iw9tV
NY+jWHipxOOJuqWbbJrwRurCxiO8M4m3OuExG5TDzRtJ0f7bLidNgzAXB+0Qxmuv6DNwwmAG8n/o
lrgErzl2diiD0oz5Y0f1DW+mPlZg9knqR4hxSbii4kx5cC2YdvsM6OENxA8+oYm1ItSCfvGgRkqz
Lfhh005el0aZ8uGIZfm76pcbp/XO44NGD67ItF0P8yzNnu+QqhhNocZbM8liCfhHGqCk/ND8JlCH
G7MpKSvoXeeCSR8zQTpcVkAK1vaFtW6r1akBM9Q6BevtS7n/tdhLMEVJUo2bjw3qeaBpV3pag9wE
G8O5gmtWu8NHEnRp82p2oC4sGz2/Sp5O74zs966Xu1am2fxsUsaT9eePCAh+eRT+g6ySJtY9Q8tb
ufxlcvle9zAW1LGTQZBzOOQwptOrkPKc9UKKJaZ0a5beF03JsjFs6SyR2FeiSFQrJNav2MknWliG
/2lIzKLpFyu2pW3dFyadhDiCQ6+s1iHFtkC7dzPqgTFwOM1I/hTF6fmGfyi2R2+Axl7yOLUMB0Cw
kOoRElYkrlIOLQebMG7SHn2juOzFeBMSLGBR0j+FLU7ZW2zACR1yR4XjtrWjjOHcOeQCJb2aVfOZ
3mZgf9KLy0ehXxUnemPO2HyCg7mZHoH2ZNoDNEm7vjC/Gf1feCPjU8EdCfveTl3CJXY05MEBjrGc
rdWtiub3o9llCSIxNvoh7UQ+yIUBnL2bcg/53nTV8UStLhezjChXyyCisnlJj9RrjEzkYkP3y+F5
WdHFyKZo7AikBd7lFT5FM7j2fbuLNyYNLXZCHyouh9inBJZ1V/3HOipRcSjuE78svPpLCj5rK58U
48ih8yCzYpHK4S1cN06+V2DGgZtJHH7xix8e0Zda+4EGvFmLu+vReYkmNhw4YQ6W+9i1at/w+ko0
qQMvmTMUsUZDBXa685XSmCf2SkTOapQCaoMHX9uG3buYrlksJ5zovFMkWdVD89EOwmJV4CCjOqp2
IA3vEG4L+9wC5VzgloW23mMRa4zFk0O74XScmQkZ45vFc1HBO5mAEj1afhnm5K++3vl3JrexWZmO
mDS5acXPQUizAR2Vls09nK4gpZsHFV32vJyfFkNQlZ+3WneMSlovDic2XF0rJGDzP6+YOc9+l4Ah
y73ye1TTmGtxywpDVzDckjP6LMRVWKXIRtB4PS6nPtbDry8/pGqlr/Hv5PMXeO4geR1z/1aN8cPs
DJaUWc2Bkb1D884mmQvCmbgx56G/xu2L8msCZXpdhqknzZBg47Ie9O/V5t4nhkOjEqS2L7bpNRd0
1eRl1wQVkEbMNaJC4iqdx9tQc6HVINT4IIbGK2EMmgxdppxIEsD41U1Gq6/iu4iixY7Z/Ox+aV6t
c/1xRYJvtnZQQTzZBX9zd0QD9k0XiK4EDHE/iUi1exkuKO34cIFiQDWaAce46HzDW3sdsBFPzEg9
/mtg+wDX3SXej6drz3WeEJybhjwz/uaJcgIdB5gcxUT5xF6P/GY33tUyhPEo5XCS8BOL/juqnEOs
STWYks7ckSNWJlwmWbngcXOiqrhgKWuRcuHuONtayJmprEd8AuDjOVoqTa+moXtgksxGduwpQlgd
U+6wbrvSHtQbqIgZ/gSraYEtFuPoaq5jn/zWxvGT+705Vae2sf5ZQWEyyFDkEz6DpNRhV2AfHG0B
ADKm7KSF/NXga+tTicPuFqKYKGSFAYwpfi6DyUTTbBNMDi0l3oQjf8IPlKk3QVwu5V/ml1jb9mEG
JzPsoH8WgcdVSkA+iuteWcaa3VIkkxDdp3HJtI3+QEFc+lqtknwPnZzq4n3Uhn8zd5+3SPKBlPb2
sKOU7Sshd6it6bDahh5la9Ex24NoJHPaOE4rTF+PcFV8N+UPdqPTzgT19QSMs4mHBQ3SH/tiWZWu
4HXeM/2Us5bTkiufxmCjuXprIYxfSZOb5sSBFMaOMSpmtaOSGaOq2KA0C/pU6VD7Prgh4WGjKRzv
iRQBkKpyYtp/rPhXxDSbeNzkZsqMSOcx3TCVR8HYkE6/WDRLInohQkyTihIGPTx1dRgAGAoWDwdE
iKcwiQ3b76WZk07wPV1W/rBqrr1y83Yp1GHbSyXXpWvgic1m3+W6+5KXrvfrrNPBJFl654ciy0JB
4cl34knqjt9Ca+HwteWpuJ6hjN81fAAmD5T0S41WFkrSy1xiSSFjmQ/IeAAnhEEp1XdELuajZH3l
zRS3gw2Sx7819jKkvG4YLTi/4BkqNhBPCzWMof+1eoyw9q5kOPYX7QYksAH/fSBHSy7SXzzWmKRj
MpL3VLqIhAkxcWJb1ow0BFZQE+QhDPvSwUI+5yQTVErqfJUafi89ZmANsgiQ1c2CFMYNIpuzHFLe
L1l7/YRinbn7O6pfF1PD7f8+knwuRI7YL2nf3kTb/5ZjlpZTlIhiUpf8yn/Pk0MbjVjLL3EQdPMT
7XBw73klYTHmUcKpGLTBmxLVxeSv5zUs4hQ3ZbdF1L9ypsXDjJe1k1QI1AUTXKkP+fc7r7mrWWAo
uuVNqB6h5Ia8lpVIbcHIiwC1CE3rfr+ZmOYBY6pBvQL5+QyJuJ6503b4nqVi68mVWIKRsltrE9rR
b+ALJopXPPUV9SaymKIplwlapdX7g7vh92bmDuBfVm+2Fwpyh9lIjUjP8JdK1rsIKb3ff5M9nB05
pPPq7xD52jMXRh2ThBj9UsQFhUyPKlZrJ8t+MUAk8u67tbL2ZdeqlVqoun+K12tE54I5dnL4w33/
HiYmiJIsLgZJ/YzdpzcPRjZT5R72cZ110b7LqtAqryTrtL5l+3YXTl7tWbkgdOFYTZ2/ay6iLrvU
/AC94VrIqCfbzVLwshApk4UYrWAhRV8d+5hVCgGDVn+hIs4sA0Pg/R/2znNhRItT5VtAi/bbIVJB
qj2xPob7RUr9HqrOde8eYCHOhO8tE4Utt5bMik/uECQ3pcsWvZOSsqS0/WJAs4Sqgk72MjRNK5aC
JocbOJX3nQ+r++8kcLcJX99U3WNhSu1QjYkp7i82WbTxkri/DG3oHDgDNB7g91OKZDcrh7IVCMxx
d0o227BL6w6VOY12j6UeFO9uRVg4950j6E0Y5b/9NeK7keAVIpwRybq/cx/Ix+T18oykPmun3P/C
K4hoebxtWg2Mk7p0zZH46zE7ilyFlP7G5MgJChYXHJAsMiqP6aCi55WS9EwR2YR0a+eVUrN64u8g
6JF+xVZDujpyoTxs73UB3FR3Tyfk87kPyMsCdJ+RpZzOlxa2EPPDsoHcZpc7hz8VEijCL58lDysy
pGckME6ozZIIqKGtaDhbaniUujB+w2Ds2gGFO59BnZGigxiHo9Wx4jIOdF3tUt/lJMOo3O1Qd5SN
etNrcCbbaxiDz5mvtbKC7Kwv6QXm478bJOdz9unbK7RlT0cRS5SVw1GxkkgaYBVocHYMdkzIYKi+
ER4GgGWXCldmoy/S1f4kin8uu9C+EjL4C2eLiFzm9rVRtPjBWLJJoglozl+c4Fc7XbOBL9T9twE6
hM0lqIHHuB0i0zLL7/JrxCn+wJX4oQswHggw/WWxBdNVJR5ZWTj7H6ALjQ0qrQcDVT0KUT54xuVX
0QlIrq+/CO0WTYTh2kJAqEvAKYqZewFEau5m2z7Qp6zdWH0vUzYE9H/ZYbhJyayEZGHOHfoWZrFd
FMelIPKTXp3Dgycg+jpC8MGcfJD6COSi1i++zhSObz0vSxf/QSVwBMXUs2Wn7DtZ356HIH+wKVmF
cEkb7jKgBbC+Z5F+XxFIOlh8pCbFva4YORfu4fYNnVFw6Hy8s9RKMSSZXLx/TizYxaxdOESqMP2r
tyMXYRjepZXSI55ODW1r6Q7AZvzJQ3EhQblBv61/shNm+Vv5k+8qaNRzbXBmNYVi1SIXBH2oJM7K
SikD0/3DBr6yjgYH3SqAUwKjLSkCUVzVSoXdamEJa1a7/YJMDP5nKVg1J9tn3yWgSr6pja/dHs6q
llp7tq1qsGm46pKs5POZga8aelDe9lgitjOkBmCtPH/nhhuAAewA+vYkESVEGih7LUH/tp0Dkuzi
XSelBb7l+n/FgbkbabmHIA6Re4v6yiEGA8vn5EtRWkAun0cWaUCiiWVbyj1mdiL2V3/VCN3yzPRS
KzN3Sm/NUzpRkvCyvD7+HuRtzLXyG4o4qHPefUvEJfZWGmON+OoKCISYaazgr/x9KMmlkfTWH45w
2pKd2VO4av03pP2OLUWS3mUgsZzKnVrwbwLMNeSC6k8dvnSIQ8X23CuEj8jMtITSWRWtoQsllqaj
iqZd9y7BxYUHXQVoa9ft4qtohuNQrubabByeWd/rilCysMYnDBSO1MSlyeZZK9UdXk59+VBvn0im
jycaoqMmKSEfpzYQ69kI8VQ78LsKWGs2+DMqPDKU72kxuGmodgnc+jPO3QDMnFIRtHvgo5a9GPE7
i034jDLaKbDKk/AxtoEJCEqtRfNegevQ6RNfGPmQqwK+lRhwTxWi2mxB31XVYlv8kq6P/V/3miyk
XsH1sNs5WkMrDjnr2yCzv+IcdL1afsuLT9g0E2t1Lymodn4kWAOyd2BfR5Gef4VGA4b4CX9jcfk+
2lKF9R9y+pCuTpfa2m3J1F5ktf7HD2YKMuaM6G3CLlOp5VpCNOySw9ZnVrdsPpi8cTPeFf0htWMF
g3EzWQi04QZ5EZDLyUKynQqzGTfi6gvcJbj0rn9sOESnf8a8cy+vPwyBwdU/RDOlnLNMP+yL60EU
xaZXlnqp5yTe0oHrW5xTs9wEDCLN8qU3UCVc7h9TfyEWAq+Um/31gwQ0Q1rewe+0z6k9VxH2q4Bp
41RiKwqUT7/dWQTld1wngFkFq86F9dG+0cfp0KX7TgfgrgYkP75JpTusFsC82D7L7HkWzoHuXazA
lo9Y7GBjIUVva1V1QmW60CM4O0IkGpEVqQMIZbsBkcJykEJBcVQPAxmMDcyB+uQDZ3fqdVsxsp1N
yUxufPeOnSfThofDMRf1BTlDPkkPrVTLh9eq+DspFsYPeqnXBN6vYoSBOsivRGQstT5yJe2WLv7K
wnIemne9J8Hu/X0Qvyyp0qeX/TvuVBuuPN8UZ0lNJSfFcijFpMdjENrq/8vSBbZMmakvyKCNGKnn
rrsn44m0hDOVLtoqvw9EWY2zbPfPTycSHWzzJftDctUGwXUw6xMjEkByGtxTCDDVFzwVsosJ76GO
zZKqqPHXOd0WrGHUG8m4tmt3XnROkduAsICHhwHHp8XCSzIrlpboClWOvowdGpG8dQkOWa5hkyyQ
hzTzYD48s2XGazEkhW+4dqzUYFeB6FJ+RhZUrNFL9WYGGeAca3B//TCV9OYkPzIoKrk0Nx9ft3Jt
8vnCPoA0Yzg0Pj/KSs77tJjlTh+3790HTPdb1hZNyB7JXENg3BQGmJgsJADwcCTPT1o1afk3E2UA
atH2rnFT9cM71vvRAnsMWDYIu2ef4QEABE8qJBd6kk8TS+BnjzUFBKjJ6m+2pm8J6Xpq8YJrVq6V
jmJOhUVZfu67aPfEioYGidsxDu/2+NOijqGV7y5MbOh8+2eMs6c7G6YDBPdjAA3loIHEBLyKd4f/
MhqdfxYwumOKk5EgOY/T6hwPcAzMDeY2eSlW+h6t+HE70wLqsVAHtDsM/bE+Xig8BQxSZzF6ppZG
hJWYVCY0BFNK0nriq0LNNLkuPvNRs2+O74lPh5+u1pqPVJ2jeqHzU8Y1xm5zORcGdWNt42P26na9
xINcP7WJgUESNOceJieJCliY5tqg4AOSOC9GKSdFs8J3V5jReBGPjlpFWZHD2wcfG33AjeGKUFKA
It/kXcaubm0zpbRL2Cgt9qxyvI8OzpV9D+Z1tZc8ZjniD5t3peejT3tm0lFf6J6Jec/2LfAIjXaH
9CQzKo4tZPgnCS5XU8I4xx+AQo21W0f8wA9qwgdcfeZz50T4cbc3F+YR/ZN5Q8c4pZSfNA8SLE6i
RlN8dhyebbCOh8IWUh2GB4Rm+jQb5LYIx8mghy55UzYSggViOmps0NQMHHpkPUmEqTWNp81qln5k
ZtG3NEtJV6aaurxV/s7c6xux1ZWs8f0qJq9E88sTLHIf03Xgs4HTA0qr5PXtafTfaCdGR2jd3ME/
QhPcATmIQA9OoVQgV/BaGPd7c8nWf7R2uD4n/6QFSINRpQaAksjiijJV3masAfYBRzeJTnccx88z
n44BaYQcrVYG6SZeYh1nTctg6FDV7sQrmighhQmwRxKwSBXnacro6h0t8Q73PsHvtngxglhfEVmL
kPNBTieeLyTIAnpFVtgmvzNRGmY9ys/TiCmwP2b92gsr/9tYhe0AW0XszHcYKrcX0n09LTd1Ro6K
7LddglWhNpV+a7V8+taaCG2st4rRqKnL5oZnFTRAjDgc2Fc8lC+47WHmt/8SX6u+S/B5ItKIcyEp
/NWTGv08GLMKjWAzFk0mP+tYdDd4D0lW7r/Dj3eIP9PS9tfYCR9zBA9HjUz1a8pMMQMUeFgXOpoA
4ZFwuzbsUpYW3Uk+64t4UbhC6uf6MXkEk5b/7oJx9TnaUY2pqQ8UQSVvVNg+bs24u/tiOqgRleuI
JKTuilaZGczAt1fJJyZfQd4LjYrs1DEyTmAov/+aqFm8WhLSDtXL8ZhafHtIIma+k7bSdTgunjoF
6HZI4sosFlc0D/sn44Gn31lav7v2Z6qRDDaU2XOEy5BwEbaPY6yWysIejn4NUex65w1Z2V0+E6po
AWT0G4Om8h3QVtQloceDDGSEI37eRFIkIwjvQiPLMayAv0QDc7YcnDovWrQ7UTGp04Dp9W6w2tFq
wOAi9WN0mki5Mb/3HUU9i360G+gKu2m/HiLCidnK/TZerNJpqoA0CQgu2aN+cHCBXAQEWFOFnoLc
jpdwxL1Aq2s77xHOLHiQVf7gZnGUoOEHzhlqipD7fD1+uHNNgKpMqv9jJqCOg/BDhMSdZ6Ve4gGt
E5EjxgFkqPwA7kc75aZj1U8QFh7GeFCQBKvnOxQarRSv0wj9pOJQ22kZJL2E5BC153+ilAv6kiZF
mGFiByWV+2GiiIE4N+YJFBDGvJB1+ZHOjJIH1OGhLJHSH44gX1j5xqFyjFR/Fjt7gyMAXyGTGTLu
Fn9HQRYGjjrp0or8fi/W9ht4pkPIVa6GHD5EO/kIupoydGVWQp3D+IYLZFN9FHB3LuuD4rxVuCRd
9KWk5Djq690DHgufbjZTHTKGUoFbtcKToVDoNuGBH3Mfe+sSiJo4CoqOLu94WKVv1SWBy1PDkJ4K
eh8oJFu1uBTod8lVE/vR3GJqPISRrjXEx2GOKIZ8jAPg80+unLSYnzTWKlyz1qbskUabXKnKKCUf
roxjTdtOkQfAdQqki4gG6+Ds+muc4nP4q55irEB2TFrWNrbnlpAnUB3zO/jHujvkldtvpVEladK0
bwcDF87oBxSyEd9vdxMlPWuh4yD6CSMkeVdtYBx9BSwmTBJ9ct65G0ikl35y37p+gQOlxLLZeeCz
D8lcST/ieaTqi0KPOKJ6IOGmlkQ5kqQyJd5/a2Ck2p/GW1xL/Yww16zBtlFfm06QKT61kSzS+QWF
Fkl6ZVtta7K4pys9y0RUuhu0wvqAhjdv8YBry4aWEuG+BxLsjwlad7uy3EBIo1XA1z92jvSFFS2O
9VEx5EyCuCIKE1Z7BRiyZlWTwuMAOXSz+UYMQ3F3d480tpJ4YBPEfwe4fT8Bp7yXQY+RVNlpBokb
ZyfUbPSlyNjfUWPBhR20BSPuj1aDAHdrIasHOW23VztaVvEd2eVABWnZLyPhF8Na2M5vORstlc+d
PCIIdO0xXYqg0ToBDnU7fuyMCeLGSp177gKMgo/bQd57bWPrD4GM/QkOHCN+ANWzeGsPUAXx2rLx
xMgmqRQZHz3g6H2GsNJ4D6Jc2dBkXSR0rBALmetGui3QGCx3W4uylayhDsALyO868NaAmqPAX+gX
4VInEPsJZjnpw2tlkCSJyr83pVN00HRL4pXPGINjP3cx0YWcboQE3oUyoHIvvXbri8Xu9FpYd5ZZ
B35FPaTxqf3kT/Zh05xIe61FXOMLu52htYgNt9bsn7MjX2BYId3xZRvxgr8yD0mPGzIH9tpg6UOJ
GVFUIa0seqjr38wj1ngJBTKnrlTGc5c4SUg/e0qYGtIe0MSsOh36b6w599qkFllY3RE4jHfcE52U
9FyGY0nK575WyeJ6wZ0HxjfDMGqWhkzx2t2P+zKKunKZalh5LB6zjUaoZnC/173gYMzBgKcHCgLM
14piq5FpPBecasTjsJ6AtXEErpq9Uxv3erRZQrIbRK6X7La7bh3s+SJYE6yCk//7lYf6Ozs59Xg5
xaFm+cBaiiIULqoer0KTdQEkkxIMI19iQpHllETVp6Ve4bg9oOogkuvpSp8oW0UrvoioDCmT+dMz
f9chTZ2SeUmq38BlKrmXp8pF/9fAWFGnlJd5Nr4tZKJBJpJfO2Hh2T/u9QjWsnax/c0vF16ELYVu
bnhlK6wK3jt3ESC0r3a3Ua2u6WCu2vJq1wUGStAoaS+rCPLXq2tyynEPwtbjsCahF9ZhmHKxhvpK
koQvgCoCf0CqzFeLGeqnjWrxfRUHUKl+CARmD109sfHmS1Nfre9Z2tvvPUVNXSJO90Uzv/2aMgW6
8AgCN342QXj1wB4O3uYxaBOdI1bLmDDqcLXAPAAnf29F50z2bfQaOSMXfrxy4n0b+4pRxtDSKAZH
dOYAVh0rZFbdepueFwHD/dLNIvtHxHX5abf8I55zltkzn1QTgYrPqmVYzG0AwAB8oMLrdSFHmKDO
phacWWWpOhilyidQhd6SsUqiBjBMJ8L9FPc+p/iMarhxCzCwfvnbw5hVGelc3FLP0kGXI75vqqjF
1difISuIrCI4yzy6gdMD/nBIOS1/AeSwHuP8UPJyQ8iCj4aMMX7ov2t3SY1lELR76069M/p5RdId
HaXZZ8C2z95pqnjp3l6XS7fah7xQo3vTY+Dl7qB4irtF8lL43zGO2mqly/mfkq6JV6DDz4EkJREk
D9EHj+gxTay6jxZiYAp0ay1TwD8wTcm6oFFPQsQM2cUnq3Q2/P76XWGwWNsBPP9YvLue7uXzBdKf
9FZpvKc3gj5ZIe8JslqlxtJ2M7w7k5+6Vicatxkwf9KZU6U96k/NFubQ4utFF47oizh5g/tcHk4j
UfZWlWm6Kp6hNbBN5Fdt08pF1eevM0wBpTiIJXeCRiyNSx7nb3xCgS35S/8M+aTpvTrplDTlO37a
+rGATzF9uK9TgVASkUtwt9LmRHtQ2sVHjmYXZRhJKWj5JiKCtVKDyV3tObCqDRAN2ao5yp2iMD4O
u3IWqU4w+d88FvfD+PBNR4IOz+Y4vRN3MHmlx0o1diNqPoWujLc9qTcUC1LQr7VIsHxDRnAdv6BI
a65hStVupCdNP26zEPEnf0XSfhflovL785avNyRJsHOeLX82vP2w48PX+d0egViZNd3olNjje/Hu
9TkJzY31yZLKEMjI7EDL3n3+A/03b7edLb6T6nF9krFSkB+bl8EZnrsYUTlY2LAgws6M3gRDtGH9
QTdbiBTz4jTlLR+TxEyLIckT+v12VJtuJOviiCrIaA/8a8+S5DMlwX7sM590ai8tpBU+1cq6v1Q0
jnOCN0aZAjyctwRAGT6hAS7WUc06C1Tvr05U0NVCnhR+evntduCx7y0VWqXQ4yQwgWV6adPWxb7v
fPA/xun1C8jWGb03bp4C9reB+aO0HvVSvcMkYsWvnN+P1J8C1dYcvnB83/kRmzyXCB0ofS8XI+rt
QQKZzv9p+SZ9gndhYz11CPe90ahAVHb1qe9QNbGeYC9o1+PVmZFGxQ8NYMTQ7BgTPikYqD/etShe
oXhAfEHyxj3zzP30mN6yLzG2wurbKMgVwjqO09N/Th706PCmIz7xx/zhkH3cfOrj6G/+O6CXe3CW
U/MsqmIrrBWEqeY6dAtWbrkGzJx9L89Yibgvs4/cOy4Nv+8g1WofOxQig5U7tL+s4Vqoipcluhkk
KkvR6wmyLAl7VwOtMLol0gwNE62r+JSOap2+ZPC9P6VdV8mIVBvlM1CX+b0dwWXQbF+WlE9t+lHC
C/EliLEzMCfzulBfYT1qEdLqT73VTjIyTlDqVzM/avKvqFtBpCl/a/6v8uXuM1Zd09AAEmiMuVl7
R/LCV2kQ2Jf/O1lE6ajOr+Mh9U+1JpsdXhlKD44psgCWshhjaiRw5KUEBR6jF/FX3pDbqWXY0cu8
NUoOTAF0KwXAqA7yKyZ364UEWzOXsDVmNS+daNdbKu2VWagauHLinKq2IAUsKL2K2tIJDZIu/hdS
td0sQScuEg8OWYBcEAJkocCNKAqUMCQN87F04do8WwwKCIaxcqRPQIrI3KbHAzaRrdKK9QB8IKq8
p+6J3520raA0z6ZATm4DMl7gqAtIb7y8SXU9jpzDOjF13iCExhUJMU1JTWsgrQVKESFhb9eM6odV
vMSoaXxpoeNFC9lPwWaHiZp71BX7YKwi1hiXkas+ZtGbeKora2R1lyvrp3eOznOBY5Lo//znTxMA
0WxwN/670NgHEkpUz7WAMHmySSVW9teO0rrDm3SzN7aowcDb8yBbPpr/+b3EWtGW5dnwbSS3eagZ
3oYVm4+BPqiWL3dya+Rk1sCXbtk+jS6Ccl5H9spipTJfSIwuvufiYeOdYi54Iimmiw8I7UMDl3ty
itWel2wJtXHdtLllOdCkOBue3xAMBZLIqMbrwu0/KkkIanon1UVlLf6UKitOE/9BKYXUxJG+SVdp
DSB+ujQ8uLUsUTPgFdosU1gN2hX6GdcRh8ZwPosRay4mcXlFD37fmPufYAhRIehN5AJjkq9WPZTt
VGWdGAKr3ro2poVpfuaNE3iK54iYk9YOGq3aqqp7kj4TH8DQsMUJ25SyTOvp/50xg7iMVkmXB3um
gXorb56XRirEN9xCeuXpgztXCzp790ExHYyMvCKdetALD1SFMpho1FOGvj35gDYVRqQorOoxGZnV
RCJoIJ4eg/ADLQYDqGlOH/vEtb73oj8qhsqmLNgAAV0ch5bX0qrgoeUEOeDctm3o6rXXVeXiv6os
KxWTtO0HV/u0tE5y54+h8C9ABooGtAK0E7u+m4R1I94DKn2IrDViIX9BDeX4zQ/7o11DR0+M6BR8
Ot4+dLdOBjyliabYDjr0DtBVXO1dgF1/8RWRZtu+2AEoe2Me5MbyeGTSuz1x3U02LJwx+5jbbuJB
gg4+ad3VNavtAqVVEc9W8wqa4zo9dN8E0l76mosI56rv0yXKRqVb7YgwJjRL+LCRmIdUuRg/Qmve
LtQn76k7d1/HDyMhQT3ddkif1HF4FZFwqak5cod/p+kE0i9KnavJ35OjcSHq0JAQ+9OqhFRR2Xqw
drnQPcETOL4eP0MrjrkqB74Cw1Kgo39LNkCb+h7P+w6T1ScV8uTfJH9sVTMt87SIurs5E2nlv9yL
Bg/Z5B74cLXCECcHtwzCKXH/pdV0YBY/XDB0Y2Q4tjL4iH3cqVjXmmNnrWzcMbZTBRC5XhLKOPAi
z5OSp9nWi2KpodfSkGx5+fmemmu5J9239mysimIV7v3kGz/TLhL0SHyNlk0+qLyHN+xw/Fhogf+V
f5ib+P8jtuHnNtnPBnAu1w5oSRYfVL7IlUfKpTcaO929Xu9NXz7c49NuxqaZWiBGiepINLOyBMFL
iUlHZWzIy0DWDOzFrG7d+ucIlkye0rMCoOTA1NYFLYOeP/PVjICMl92hJWszTec1QJ1iS7Z2yJE8
1GK3S5rvoSa6T8+7JVqc0ERvyY8AdVUDtAm7o/EN5mZEX7uTE8TnENttBpFIEkQHrxHfW3JILNd9
ak0UyHiDyrEAncDxzWCPhDeYTZb5AT+yUrV9EANz5GGMkrCYArw1NmhrDlBTCprMVqWo1bVjRtv1
WymwrhIZsLwNsqupM6yvhHDGIilf4AfLyiFnGpwwV1ijyKGDi/mNN5QCOUb2eOH5k1i5KRI/X893
tofDcctkai70NwOMX5WCB1egG2ozaexI7AOjoir93Epk7E7spYG7wMdD56sj+Nt4wpI4ov0jsqE4
kDwUEyNto562tZG4lCnyaRf4l7jQnODUTeT8gU/mILiA+ji/wD4LwA+/mPu0HYO/+0vr4cdOHaiB
obt5VAJG776IVhEJk1YlQRpPwdRD02a7dhgGQgGPClcp2g9O0MMbDS1u61AGwEngzun6+wK1qFnf
403aINu3TmvD/R/Sc96totr0682tCWlX0o96Opn8ZOHYWgnpyxfET+Rg2buRZydMl8Ikljmju+XY
S2Qka8G8bmKsU3WjNJ2BQu/OexzY06xbJwg1uuCSFXOaRhByYbB0PfJ91nKndTHmX9ypsj1ob8T1
qi5GqoI1hAzATZizkL97O9JnEfNS1XDFA0jW4T/zLGRGz9yhqFZ4SykJLNmeS9/lhJI3kjq9wSI/
2lKU5vFR2XQyfwkUiqodO9Wl0Ib2VkQCPQR9QP55Un6y0mVK0IIbfyp6AJ8FgtUxQDRNJV+M5E7X
AePXRZsRQf7hTL+YIha/gN+QMeqlRWeCePKKLw17ay7GNMAz7bid0nGrCx/U7j2LsdBkHZ8mziXv
s4k5Qrt8vEC6wcOUF9VVs3pZjIJrK9aulKv3ED9eHpABelnehJy4V39ep6BAyzBC3Cn9il1M8yPv
oycdhqWrfKJnZvz468zcQX8Cgz/uuBITtyG8WfViC2IzHCB2ubJTMNIB/jBsUDgVdHlB5OUErpxW
SUhhnGIBVPWnO73TsITnQJ4/xB0gmLrt0nszMqW4kxjME/qZkqDGLlbT0y+yQ8UC02h0KFUgPOah
8c3cJL34LKZyhrYaSSk5BDiQsbw+wbcXxDG7ffYWbAYLOnGdv39HjmhVGDQ3qb3ET2FPlQtgUEOZ
dFwZQTarIkZCW2P9ncrqs0CjaEewLukyuR46QVCWWIdGY47A5NCdomzImi1q0WPKYHrgxNg0p0mC
4FjHGKPvmux/CzNpRcVSthJVzvmY6JWAfRq74nYuEWNz3otxfC/R4QSxMnS/SZVI7bSvFX7T7kdu
atKCp+k/btIJCEP9djJVHgj36DDXDBhZ4486PwH+k9qaM17yWgMvF4UROdAjxtvFbwqrOIzqvK/O
Z+ckNDH7MjWlYS0hWidwo462iB6iiu0cFLpZnQcrzIsoJRbga7ob0fGxRYUXXaib3BJ8foSC10xG
eO/Wc/EMszvLdoPt5q22MDN8AVs2NGQ8cFrvjrpch16vM29ausz/dYM82YV245vvtOv+oiSzhetW
D2yWHPZNdmT4loBN83uHC15TwJAVkNeTjzpeImtTb9n4GOeApFW5iBiNvLA1BOKJvyOQYXfjEZfG
k2Nxfe/lKsGPsqdsIad1yOKPgr0geT1wIxSnFMx4qq9YahOMfBJfp+5NNehsfALpGkCW2INSN/54
3Vm59lD7KhIqtBYcGw+RKyF0zzqpcmAmR2Ogn1YHMsEHrwRPsTdud/ct5kt/XnmtJxybTip/tCDu
ySt2DwdJ4PwJULs6wqnItxxqAIMDd9reHm/KDNQEsRVW1whA8dSBoo7ryMMv52AoSFrxgSmPRtRi
p7NiHUdDIqIWnjWlAVED9mZ5zmCnnqqH/IXc6qRki0U0VeeOwyNTm7wdG2EqwBExHe+C+CmIBZDz
iBdSG1b+HnsU2kHZkJfU+TVGazPOsIYuq2i55JJHy0nea3AHzC6xp2hE3oWGEyzCchkFIlHVtQpM
smNvNQr6HQ+J3KgCvSeOcZChjIEqka0n4Jd7KCWu+xU3HSt4e1CAH7WsfX1McHc6cwzmyEjM1Qnu
iyHaWcDJyfs6HgX3/eDfcAa6BnyjCi3FxhR3ldyrpUkYVWKlD43a8mJBTMA25Wsk0QfkvJp9UZSa
6H+RwnLgLyQQ+2eTbW5VtGrThDNs60Kf43O6us4L76RS1smn7P7FzRldc49uHXK7Wb+5wuYSPKw+
eltlHJi3xuTJr5mkg155WO7bdAI0aIkOZ10WaMbeSu8EGWhbblIn+l2RrerUKf1/e8+7DGfn7pdM
47D0Oh8AcT9/q7NO24dbhQUCEUwdIG9lkUbwDUxGE4rstuYZDGBULgnvlbrnS4WCuimASoqJygBL
/d/SmIOEcgUUfchdkaXFNuFRP9p92BKql8wMS87CwKNKRMjXUwGM/6rY6z4TcC6Ajc5qEeWu1aHS
Yj3qt7yqDbNTQGQuM9U9kSXNTqdhulVQPanFFmkJEnKR6ecv5EkyefFlaw8rCfZtOzxx0hA6aF9T
AiXO/PGwI8hBnIz//UOZmmNW6ii8JOxrNKIqoOB9c2Q780PexGJU0qv6NIof5B++IhzbompieWtn
u9xI+h4q82qQuJ/7kT8oaXHbBurZRSL9OTI7Zy1OdeaDWTe5EFd/dv3Sg7/X3WBJO/oZ5ckz2g3F
e9GZTr+VRhjXJdedSQYwa/s7qgOQeiHkABu4B1earb9GWQ71cL3cWFFn/YEIiBrl6aGpkefxeFHV
2nU8sSCNkDZnwzcFd5ruSo8EpoPk0vykAifm90KECbV0RpCDJqrABBnAJ1I3B3/wkFxSLgDIqAoR
B3IgzSrELr+xpSD94eLI04eZUsnUAmwsM18Dm7SaPrI5+LhxEes4ebFtDeA+zna2ADlrXHQ/jEAS
IfhUjZrIPYBilVrWFmcJ5JwtKc1gNoAEuBojIJiGpxpenltPlpvlHZVJkN3wRXSJ1bcxYAes4QYN
ROk2UxcwRi6/Mih+QwIu2s1v1D7/Wq4LYObYcDuGjaW0oEXgS7ssMHQt2iwjMjtAwhOtDbFhcim9
TVm+rXW+535fHAIUJvHzbQ43KWmkHT82Lc3r7h3VQgiqgkniV1XfQADzcc/lPHqjCVU2n1PUiV/C
nIok5+AqOcGCzEA9G4ClBlZ28klncCWSdimUiooKUDb9XmDLwEQhz2blpL4s/CxdM1KcKyAc6yf/
4u4+WEMlmFAAeT3n0Z0HHBxlOeUuPTnI4uXAwjdm/H/ZNWq07NOr5OglmuCsIF8T8cNKwl0bMJV6
olGfhQyXYjWeAM8Roys/pu+d6cX2NJqk/OeWVu1jYgnh5H5o4NucisnqX6yBF9F4eX1Ms5YKc0Mu
f2eDUrtZVPsJ5f9YTSxcUFGyByUDL4BBNWPVGDQB7FQ8bnTKBXXrAHJ3/dnOZCgO+j0RPQY4/HM3
X0TuUYZTlMVKT0bnOMd/twMFbhN5wyhzNAJD/e+MFGVNDQxp3TVOe5jkoRYNPOUfvUevf0rkHW/u
biFdBaGT2kSizTL+oZgsxobKD2MzylLKYAOlqcyUFr85pNqbcA7FXXteJjsQcAZmJm0HCIvjN6ax
QJ5sETt/iTKySUiBSEF4wJ8hzPnb8S0NKlY71UjajaxlfAxAumA0EOtO/9jQuNyz05w62NhXZtTN
2IE2uFDn+JtO6BpqEe9idZr+wEUSs2TU32IUs0hhKbqvCXKNhMVT6Ga/vdx61/X8OGL+kQCNYTya
Gf+0rVJPE06jDbViYxXNct6njq0LynAHb2wJ/Mr7Jq5mffD6Xf+39XQrl1SnVH8dOc5cU6zhy0Jt
4Uodqs3Gt8sleOObp5jH2UI191M7Gbq1qxhN7C2gf0acInlVoCxUlD+5Ysx6P4iMdw8lhYA5Hdzb
HV8Y7MQA5plwcsYZgBcde1mqR9jJtJQ+2M6JZEvSbPdLkLphU7ySqxQ3fOe2uNUyvtIXSTW/WkA3
M+TX2J3uNUF3iryjOT1aLvn/x2khkI+sqGLu5j/ByrX94wodNh+T3lDvsNUeq0x/qcTNgZLAlP7j
WaIAb9eLAXrC4F9QwTj6CTAznrhyErXpctZmzP+RQi7+XtLwtFd87i0F0SzqhO5QoMqr2WOZEEOR
hiBjiNRXK8Ck8N6MNtagY1uyShnjqS6jyzsvr14rVjkaiaiIknu0q3sYeo0Y82JwMRcSEv4ElCOH
9s9FYw9ou6O4akR7OpvyM1esBjjuVzGtd1nqfcCyp/txYiHM3pjr5H97c73IIzUNLOQnAk83tU1a
rec+7oXCoihfERMn7SwVCCNpjNz0NzDSXYpka8Ajox73bYszUHD8696szjhccZupevRh1HXTQ8JA
BXFr1hVGsuMfHvCcOug+noFqkoyRz6H5nAnJuvbSi0E3Ctyg5bk02KUL3Ric3JzdcXpPukGpWDRC
KWlcxZPECaITdq141X+TZwPTN5sxftolbpl/TKiWs5HjdUaOms+CIJu4HLAYs6XzrxRf/omGMNap
o/2ZrWd4oNiORbUSwnzuw4s/4sbKZc6RwWk06kzTfz3F6suCBPWPP+tJum7nDISWtXuIpz/4J5sb
hAC7kuBzMqqonjzjrtrjj58CDhmfZC0KJSL1CHcEXwLGPEwYkx1JZtErijaDtHLegfVvirBI3zt6
M1/P1mSjEHyxADA+j1Bkl92KxVqCbE+nMAknOzJS/BY/3LIeUExpamPvUMpGiRhTNoczYPHVnxXl
KFIps6huJI3xKSbz83CxP0rCkqFi2TfCWjsUw6Z4OkodZpQcq8g+002diCUJmqK0I452DZjSM7uv
E3M/NxazmZlYgdiqh7AdSfQht/ASd3q48NsO/DCOotEdVAgWJx+bMQgWu7VnfV1ut9U1Hm8LBtcM
zzWOLDSbQzQul1SvZ5E4e6x5JVflCjrHnbzwqmEyakl1KC68LNf7b24lw50EgCPzm3A05KYbXHpq
wa4NcGhgxshop5LnCtC4hQVbhTz+kltpvaJiLw3SoOk4wIteCFkoiPUeqXQiODmkSMlVaONq5Gix
9j/u20zppefEqywfvY3Tt3OhutSO9MOlK0SG691ddQC9AIeG13JqaDc/iRCrXde0vwK9LpfnsP7U
80LuppzN3cIUox3QuGe3rrzsUZKrO6h/LBibRjEBO67eCo9mesAtsX/ETk7Ji+F6ATncMKId5Mq1
pX+d7q1fx5rAWX66cATCERJ7hehOTZfj3yPD7V4PjJVz4AxbXV1DLrvbx7wcVV4C9RcRf38nUc56
hvaU9IYN2s9pvvz17EYv0WZBh5alBPtcAoK86kMrQXm9oXB2JQVTiZo1gKVb/3PWERnW0q5Os+sV
zq8QhwZlP7HVw9R3FY7q0pwf45TSDuBMN6GblsY9KmcxChb7d3Wa4OF6NsQ/d+25sYP4lwpqU6DX
OGjTvQkyTfcBmnYIajzdKqWGp3nFUdN7yXU72WljMgE3yGPB+Zf6+GY7L8PKs8P8nuYjnNG1wuNq
uAadJnPX3zsUJq2yT9v+AYlOi0uwQvmtDSujxNj9iHVzkPDVmOe5QXYmw9EvXj6LagdOii9DhAzc
nS9xN2bNqMQq7qJiKSqu6AMpfFafnzHhcmFS2mmbb41DnLfUIijcdFGk13mUPIsnFCfr8Y1Uy4zd
Fm2gU8I9ycGE2jxppiSO5G7wzGEos1sFGfdCk4H/LB4eToLw+t5V2bZH1qXIDbvWnXJfzwWPpKm8
ZFYoyRfeuwKpKsJxKLjYmGSRpoTP7eju52ZY2ShtlpGypUlIiYgXdv7hrN0rXoycw5NKdPuz4bxp
CF/UlDwsh0d8+XWqrr+1ZiSo9VW7dckibsN75z3JS8EYDX77bq2Gz9JKUNf2vsZ1dvTuKVu6GMxh
SopYcFnJltswNgdLc8SqhKQIV2hXhu0dPts/7AU/mvYnhTWc/0uu3r1p8agar82EpIVskiM2lKnU
1t6JE4GzGjopGfRpsHBTqfPvsMHM91uoerRfpzRVLFkD1yQvb5U2u0yo5NpdclFE+rxdHq7VP/9H
r9wXbdnCzfT8X4OznheAzWFBHe/domtqlmrKhm+UaI2YFiClz1fPuAZQVFCaxIU1VPMKqhcKLZfJ
H6lrgLWOqEuBhG+nTP/sALmrExP453+ip5Q83a1c7I1bJlarx8dMuMsR7rS4mHExPQLmElIczrmf
48tW7pwn1v6aqwS3h6lVQn3DhBhKF6++xkS5NqbnDA6x3dcyPSuwKabOk4NtO/miA28URMUT3LVE
rTpR63P9yp8godHJDIJQa0pLtnqfz0YwsYZh28zi/BL8Yjb1w0QY4+jHtta3v/0PqtxrLU2U6o3W
SS+WyRjCi36WAt/l3VEMaqDq3rsmqwaTdxHYC6QnYQY3Na25utLnai5blTEeYoBb/EQ3iNOJUZvv
bIs7pBncndnxE8l+LJLfFZp+dqVMq5jVCTZUf6BIcjOASTxmABhqDziDaWQzSJPQMXRt83kIaq2E
14KVtl5HgjSyB5W+WkxpobEATpdcR7Cp+En23Nh1+4IplJonpisET+geCUSgEZstBD0G95WgUURq
EJq4penhxtTGma7KQVRG9VPuiLzSvppNAa6mTNL4hLffGP0+OQIGhB4JearneDNhTZMu7TYq/YeL
Lt7c2FVWs+gfCrSTffPGz0DaCUhGTnL47qXOgo/1krQeJvSwvekJVs8CW8aP0crfCUatozveWl1N
6WxzeH7AUJQI880Q6bPWRIH6AHM5TtOqq2KkSPf1YwTNx6tcQEKGSFpKkaAVp2yTD+Mcj3piarx0
D7N88tNf84A78gBG0miN//ZWmO1b3jkpFR9mj6YsTVuVLXJc1x6BG/UC9Gb/POSJWGOnwZ/ukKEx
XM9ZFljb7xM8YSjBTNWX5RIWk2aSj5F4Z3yMkkyUKI+A/VkjRPSBnwWPrizzeZUIFmm9YBWNdQ9N
zECyNkLlN4iRMPfYPjxLi3unWQkn7enoDfNDgN07vroDNYFMFC+ykKdedljjeF6rl1GbOV4THMy+
Okl4Pe2yEzZiZLOlrpDVRv/X5a8AB2p6xJN9Y4byVefiprth5wErsljBwXrOodJEVT1XRAAkxNzR
UTE58SDMjC8tn6kk+WpxLmSvO4MyrML/XJ1yLLkeHBy1zi5PWez04HNz/gXz5cPiCE5PTh5RiuWq
IaqskmVNn6IywtOBfizRJvH+eTosZLiBzmVS1fzVogzIpLDOTgz/d4JGevdpOpBJFoTMNipV42TS
PwUlCO20GzBuqMSo5wI9kwkeF+RnpVMMej6cDKXjDS4u/p+kbj+laW6XOqfFZgZ/lm8A9DFk1NOK
b7inh1ErSmBo8Tm5ZRHvwxmF0v+PB9bHMYEuFfZiS89ebx0UxURnd+fwjcgYxaZJH68cnLTTwfi4
RNd+wnDxlRVBxtGnRlTGL5AMjfhEaIrakDUQOXNtnoSUNTB06UcnEUjqxHhJCqCkT/3c56qr4R8U
cX+E8ZqGGO4Du/hms71Kla2af6JoqhyCZYHoizez32N0aQP1Gl3V018EOf4MDS4ErfH7Qjq6jop5
dI8c55dm1/uI6hRrIgRKqKEYEuDE12VL+Qzf/Sln/Nu6wwmynXthIKj31AFnngjYDcwVZFjbct8g
/jZxCPYG+mZ9N/BChmrdsbMowwVRCrZUZrg6bi1gI3vppX6nV+LYcNwR1UtC8OZrJ3x/hoRFQ9GZ
5xShZ8v8oCqqOxECpUaoNsJpjVvjXs6MpZ29NbgYvuwqE2hyiCRFTJSKz81Pb2PQ0IOoUlN0U0s+
xHyvvUO34J3rZ1U25OCpBd7GjhPo/duDpH8doifedxCIWDLOEqct05WOADH1zzXETTTlAb4S/JrG
okmJUaXldI0Gt2DDc0omcF9+CALY2VPws8CsmPfMLfMFF5ZTQ6l88o73f6E4PrHy9EWWzoY9NDyF
2XZe+VxDWFbN+GlZ/6iCOTykK7IbzHiBpoQkeAVtUPcNmOPDH4y1aUT1BvzBfBsv/2tAjNkD134Q
DyLHQAI7vm6qBbdkv3DxUyHUci0f8/h9M7DlRPLRr1Gweota9z09Bu9KZ6g46aLt6Bms+JI+BE/Z
qr6RitZw0judffOtQu1yN0JHtUaxp0xcK2n1na8lJ9nycuENVGXWti3rSd7nXhPoZly9QG0v5Dqu
3TkvwoSLFYGcxP9TIUdm7uVLUCuUPxTzVeb5G0hPFpEn8xcHtW/UbS/vnlwI+Gl7oERMfzvB4S5i
R6FSwPk+9QdYheETzYYVH6Id/2jJV/LD5YbsSo2atYnyReSggwUUOk91k77+VI429qP6xPI1AfF6
QpkVhxRVWqfBzQZhh2m77UE+i33yldwGNdRUu4axQGMubpcbFuJywSRGcrs7L773c3xKXX/35KID
+nrSTEzxqp/gi1l4e1B6+AGCIIB3rX7wC1Kv/kt4nfbzS3ffAHd1cuo1NEeIMEp4rEpWS/5sDuWm
3Tiai75/tl1e+exHzaoSz4huy1d5fBpwMSPkE6/CM/+yGlY80T9abXDfK5GU7fpYFJ8iCPJyYDsD
2zDWnk2iU/4ipogYdarzfViErIscGybal1kKlqeSjQLHOAktq7+yfJ/2hdSZT0izsRv5pmtfSgdb
dKpmougj/nPRZfPSM414bwsYHzxiyj9/Ui7YqLeqgnjmFbPif6rdvPE6O0zsodhvVOD56UpNZPlj
YDtwkGnsO9r6e1xY+j/s2dJhlH1SsYOWx53cwm06qGElu2HJTRY4jC7khUd4uUjda3sV7bNXhTmn
agkkdCqLqB114FDt95bRCwzsyUkj992mi6jMsveg5sNnLF9Kbs+oYVF06ZRZzXEB3C2/bTCJvXqO
XQp6H1zsglyJrBBegIqDSPz6+yT4+D5yQgVP/M6gZHw15J5rK7Cuf5bpXgfw6crOE3NmfC7534JI
C87aMCdnAM/74nJln56jfkkB9nwSKso4EHWuh+0UxkeT52VIs4eYByvW6HkxM1yj3Cy8yd4nVBOf
JTz2y6IPRwwXimFeEI57YEKCNAlIJpY8wch2zyxFdjAl2lcn81n0/jAgFlGvck74IZjho4OGgMpq
viLIQKyJ+tG+H0W62fwhFYIlpQcm0w+uxw3xp+bXRnRLWpLJUSh0EOEvaRyu9th41yXdHlAdRNJ9
pbSOAe3eFvJUyj4ivmUPmxLtnP2zq8YZW1Z03HL//7+ulm+gl3kBIv9UirtrGT7smzzK6R3yfXDq
svNQ/kv1ScSvjFV/b2tHH6m6w4t8qM0lbTDK/p9jNUGpKcmV36Gb7FPXX5rudpcxnBZU7g5jInrd
DEJfqQeDAWCazLHRcRFdxC/kGMIfizzeSrV4p2yZg/9e3czzALapNLKGp3ce65hbSM6s/+Qy+R4w
PEXilVDuFn+ObKMWqn9B7vXlDQKr1xfjPTQVlxM/uzPrRTb579jFTgNT5JpMh11L3R9OS1QjKBNB
REPavEyFSBaNFd2jv0YhzzIN4fzgHBawSwvfKHKnHc0cMti3ljoHoKqqF4zgykfJxOas+urGKV3W
3F4QO4yjLs5ICYbVkAbPJwrhR7l9F61kgu8aBT26NU/niLTxdmVm1rGTdOAiIsm/GdaSQ3WAjUT1
5yysi9ZxEHuf+uQZl9mMTLLUAdr6t4oyYuTyvzhPNmvGIr5xXRBqUUqE98z3dHqDzfr7e1zK7r2h
qMM6LJD88ALxKve/lLjFPvMK7lqYnsxXpiib01FHZU7XVpdxc/EccjnRIF1/StzMaq3GhzHNeDad
z/wUns8d7duie4AnWwAeI9nTyMXPybgabfXdh0MualjB2R5wMXNiPJIwiqk+jKT39MconjLxgdxd
zP+IwaYgmw+FwrvX+FMBIpybcSXNHhN8kU/m+h0q7z1iAraH0+zLo60F9tMpvRPLiOqM+SG4jqIG
AUcy0WFileQRcukdX1rNrLg7FfxComyNJS7dsPYAWwPtmMezisnX7ZebMyYQkAGg+pSHVfibv5k0
v93ajqcL0gq/msZY1SrJPz1WnoG7tutg8u/HmYiJ79jv7svTAu35j48JRep/khB/oWqg/R2Ekgok
KDSEfPnuWKBUSPB4Ow09epG7Q7nWun1QWf8BHNpMLeAw/YJsol5tWh96+rrw+AIrzMzF60shxY7c
9E7fn386RYav36PAVE54E0yUXQ+8fGShyEXyxrUBak/u0BGuaJfmPy45/rktVQK5h7jDwu9k3NaM
cD5jZLCpO0wwyhwbV48qrlAlJ+0vO+t7+SToTL8g8/Yfmd94yYudVFee4Yh2C7XzqWankczMoYL1
KC9w/84UtJGLpXceI4LrQFybummz19iCydi05ZQFCFI4FD7i/kAEEFCNo0Vpm1Sfx9cyPW4QgJzt
2p/RqM5+2aNGUzLCDFNIDHe6LYGJJk5YTqb3Zk7BwbcqLkgcunw+TG37GRpWrPwoWerJW+AiXjCm
uZV+75qYpRgzLGQnfVmtPjfmOt/vMmRURza9PWuGA88KTrRL05uyqOe4bsJqfdE5TxPa5x8cteoh
1kfkBDePjkNLDRNJ/R5oCAtRfkIRHiqerApJkvwR/ZlpEaL3XsMB1+b26Z66b1VQCmBA91emWudb
PCkZpHG4uP4riRXyfG2X6H+SnL7bOUEu0MKj0dX7/dN9Eib6pN6HVpT8Nb7rVnFt1X956EmCETit
9VlLS3AnakrsC+xzo27KDRD5kMHaO3mkLh0ngiqcuHgdYTIfIJ352mKvZw/xgmNpPgb1dspSpcX/
yYxR2NiB3hTsZ5A+98Set3wdJumO787lO2vegBYqTLwuLAH80EHGcVhDD9a/L1SMebFezxDbSGfV
PxeQcWjuPcSdFrOVOPrWvvUSrweTkXykmoTRU7XRUHyMuzUg1oEAZVBW/ZSqccp6RwILjrhUJPhY
w24/0BopKAJ2TgVL7HEu4gJJ4PY+3z1V3RsyGxfQAfNjHn26M0E0VPbIEPOlYm/p4G94BI6Ha70R
XG6EA+sr7uRWVu3ECBC8Cj8d1D8KHKWZilnYwprMF2/4mdga0RBIDhkDHoMy49+4IM3X957KOLgk
EvSi6kO9A3NyBRBxvxJskBj2Fz9YW/230qDC3/6njIGvrxqtAMmab5XwtggbZLdPEUA5gKlGHkah
NSLeFdXBohwz+HClfZB7T9M/8WEmdUAPHMPpJ0NdLIyJ7uHJCxNMSIEFc1Jdiow20sVZFug36Zpa
/h8Nir/o/zcteetdD1EDMpRxsVpl4jHyLeQaDcyzSUqGVpGTuYO3w/oI9axt/qEo8UQ0ZRtAphin
41DCwWiXFeuUJsSkYK/5GEeRVRHa3Tu7geJN2QZlRBmluScu7qIrK01IT0v/dLW/EXu5TjO/7k/R
cln8oeFGjKJS3TkACN8TVxmJ2icCmL1VSN+idWJcRoDMW5IzyK19gMbxXydP7msThFz+nXk1ltFJ
nMs/4PtJS74rayx1XGyj6g8m6/f85J3y3KLixiiTBElSno75hl2il2l/8ya9JfvF146f6RPXGY9V
vL3IR+0s9KCW3csYFQQAwL8MLyirSlR65rLaVCkVu0l7A4koxQ9+PYgNX/VCjpLBJYhEIdb8Mjmo
JIz7VZ38ZMTpO4x4JmKtGN1G79w3DdxSVcUrvwzZX4YPjwL3V0D4X2YCPWXl+554fi9xRoO01q5o
CQTKR8Ix4u69rXtLqkVPtCAdNMLOosmdffr0cYtsxARMy5B4HGjBGyv+0l++OpIPpGk9tFtJEWuB
MWBiSffhuqkkOturvJhltnyF8bclYtcE9zKCL6yaWvFbhGf9QN1ma7Zno0fO3cUTx0LBjXF1rwAm
hnkwN65hYcyuMNT+MdSKvkHNllhy66uo7SzIrAjJsAVsXKFcJixdZ7w4Q+5YJxNpfOTLRzYTKkwK
B2jh9Nl1CSiYN6jmfMCd6uc/U6VAVLsF8aO1rBvudxRyc3t1RPoNdn6G4PYZkULiCO5ZNPo609yh
6yXruZnMuAzNKkaz++UyForiSq99JYpfRTNW/3C+q1UMjZwsj5LUhM7HUSzsnTtNtOwf5KLJrSjx
zcKs7prOc+HN35LCsPSKzmEgn2IjfBFerWX7bkSD0fMh2RvgeJcWGQYQZFxFFYKOgD99zNH9b6XK
JooYncd6wTuVst5xvIUOesjzBFvP/5psmihdF2tnvlRQtFrbyluaIbHTikOdO5H7P3AJ3ytkOZcp
fvhc9JYcoSKvFEYB65KOGu1Zf40uBF8guNcCUUFWG8UQc/YAE+AuCqdsLghBQEmsVc9xDFrjJh5n
4YU/WboS7tJBDpYgWeLSquKfZ6rtX5QoiuJGBSo/wOC5iLd6J2/GYKUeOUGdp1QFIkPBeRfIuvXy
+LIfSPV6a6rV1FzFIDVbaWwXJYLfSIYYQcf9lXD0+gAsvMvEs00cNaZ7Dtta65wKaP1p+Faxb4kr
n0BLcpXEHdWg2TlDin8qXDR1BORdUqkn58ta72vwa+6py6GWluk5J2uLO+s1paSgxiaHb769jzyQ
LNyFiNH+OA8jh7g+fqbzsKXK7Ia4CqpwuWWVrKPyD50ilX1Nf3+P5EnV7xZm5B6xBJbrbvmWVXmd
Pg7Drj2jHbTWzDN5MhYh1HyGvSbQKamqt7mBJsmcY6xQIt0vuAsTJln2TmLA0t7yKGbFrPuWEd/i
Z3HDNwHZaITAe9dpUmGtsC5WF88faE6pWmJtriWOhuITtKX82leOuA8uGhYJLqFFZ26yiRpVKSww
HPT1X7TZMHZc5SEOQc1GYlWSuk1JHRbsyXt/JL4MWU8AwKOnchL85ISoYS8dpXYEWPMoZ+c0ax6W
0yPT4OInHBHHOb0heByCw/Zuq/ifSd1e/qIsVf3XqR5p7xfSGhbdTAGJ/yKDbY+5dXPqmThol3Xh
DAEi16jkn/lxokqPgEBKrAJBVwSkMksnL/02a8iq06Gx3Qxs/M+mikZc9mq974dckCMDTiHoBvb0
j6cnsSfuyoB4s7Ei22bPY+1XiKT6q9BzCzDOdH4HSulIOR9XyF5JrfHLEFbLD/890ArpDX7WAha9
qI9vyybDYgtvYDz4+k1CHU4jDL6Hs3aoE37lAEqgqg9j5h3Hgyur6Phk4pgmKG5vCABvRHh5OINA
HHc11iZnl4B5fpbsOgH9+y2x8isQ14O8kOzguV9gLVSZKJdOt3sbmmdRC2g+lgpKiJm/8NX4V27D
T929gYmptEd+5OnuD/KHSzXJXUJVEIqNTfSiJKP6oxGe3lOUY6LEXRtHG4/ZURlJlsbJ5lRIRFmu
PyyMY7qATykWyLYHTKnJNoc83/ptcky7SajH5mFUV744OFUvQsWdbv//NCSLS1A3q/CdYV3gWLyt
DsI4IYIT00A/o9EfV/f8FTgw8YjuC0KVluiYwsbs7dfyUF8iY8lS5SL4QKnDfCAHCANOXMhlexb+
ZMSREFErkEyJbdD1OkRzAplJwSt3faG22h3npYJP47RtAI8ii8lKHrEW3vPfZZEhf6Wsrca9c7LM
aLPlwlhfQkMCLqNoU+kUuomH8Gy9ctdzLOfairoN8QLsh8QdHebxt4c/jhBR+sZheBlfWbyie6dG
0jWIu+9K6kggTU6PDakqo+7qre5oqKj2Gxq5UCcG9Gdl4vfdy8LLVbgOrCm3AibMH4V/NA+trqQO
TWvrWgBtp5pVgEYkzShL+UVHX21+BwJPc2TiPdWdoyO/nGd2H+9Sr17T5A99qvzs/+lH3wc8Ug+T
95oqE11Jvmh2J/vJ9ia8oPRMV10nMsl8ibLMxxsPcaqVJI3TZp4dkDQzvJTytE5qzvP+vS+EdbrU
qg3vRR3YD+F9ObP0HSxsx3cJoCd/e2O3gu7WysemcSw5N6n6+HWy4fQu45/pxCpFiR+5yBBDgG+T
L1wP5nqtHoO/7HIARZ+a2MmCBc7sIO/846PH/L1heqkgJ/8+vv05cr/ZEzu3hptTB4lejuKX5j1x
J7Sv//F6pORqDne3r0TnM3FArW+04XVlENkYylhLQsLGQa2KntJelHkdYjXO1jNuWQZ7dcH2IsEX
iSo4KvSHQhPvlkIws3iZ8Z4ZpdLL8xHRNXGAHiFtNSwtqhNnyl5kpyLonRxKNYh1bk6tILyxti3L
J510Ip1CI+cZd/+ZapdbC152pVKiw+9P5QprQBJ1Btc/KCEZ59CMZdLU2RUNpKqG1No18v9SI3aU
KR7bh0fRBJKkLaY1+dkTWdItR5iQGLhDKU1D3ZBFPGZ7OuBVdvNnMt3i6bxltlIbwZVMlh11A9BX
fAYQcALhkDZQrqmhlvA8d8l2yBFP/fQiZctvGkPwF2QU506HHrJxl3jpyZYSfHLdrID+K9ZTzIZj
mprYz9+IQX8mDNhp+WrhIjv8l7xJ4JijoG3d06mtREUfqk5Xc2be4RhSrXFnY7221qFIhg5pmdWb
nYo4zj28ZvifbvsY03XWDVlmbosYWx6KVb7N2bpJuNXmyEM10ga6Z9KlFRxUSEUaZAKuIqkwiBKi
eipLEvo0hptqtxEWcQTmmlCccEJ68fAyGK5xegVpEzmo+Mfr0ILKmqBDQl2HmCXWi90EFkY/iLag
4ZH59ATPZzgNkpUabn1WunSxAe58+rvjiQjB/Z1FLrzHFPahMU0KAWp2bZf9nIMXtC4XLO/YoRTj
buc2VGmsA8N7lviWzwfuJImzajkM/pEv59TQuQRpodkfpjICvQgs+70VMNO6UgR4Wp3TFLJK4L0x
j6ZdGi/A5yCLpn6Vf6mQHOP+pWyCodNjSx1+aVio3D9Sq1VSCvI1R6Fh18dcz7E8nme2DOHHRPaQ
8D2buETsSYXuhnw+VaVhLFwyK+tnYoNwKTrUZSHVAMk5Bvzhi0nSFBfNlz3fTguacifg7LI48o7C
vnwQ3dlXPTYYKjuJyvE6wqhDoWZ90KLUeLP6xZZnI85zDQteBHXlC48y0F3dvvgj9+5YfAqVIxrD
IHPnDXZqh4vL8reBt+mmOX6S05LbW/V6npZ0BLQNZsD2kNSl7vAV+gPu5iuDHUk+sfxtgJUoAquf
qtljlPkGpSAvNihTzHIU7zbGXK6Hpjmg7kvVoKsYD5Bt+g0j0pwlkAKeUMMMDrwK2AFqSlUeZecC
BWBsM7tLORUIlhe1tTXJ3CcUiOG/RwHgmz14MFBvpXgifVkUwo8jEdyc5oTExipac+DdiKZk8Td3
VbF0MO+Q+79NqpYvsGuv9fn7mO4k3jHN/g+vay5qjerwON7KwRL4yuq6DyoL0mrrlODeywSH//1a
jHHs/qjvtpiKMKZJbvSZTINqV+Va3w2T2jpak6yB0zV/Cd9OdZP4nB/4xZuGKqtMDRh/0wKsE1Jj
+qdo8xADkKXXEjCzNdD4XM4W4lV75rWKQxnridWQwr3dxfPeoRs7Q8nLYM3hc9+eZQeU9WJLDgvG
AsJVWRKhCwfnn8+gWdmDYQK0RG17og/Nckp2PXdqxy2JJcaTac+Vowysek8bwzqxaSqHhKWPhXeC
+jsyWoQ/AQe3NgbpFopel84BkIT/YIqLUXmPXx15tSJ3u3G+ioJf51R97HIai6ppQmpK/H4kJpFt
VmeZ1getlV9TWdLJDs7zGSv5G1BRP59TO29GiGIx1mEdCvK0kBrhGXIzwS8f9ZNtgaucck8NeerF
7sFrZjGnwQapotfUkuL91o8+UqY+jkxbA/LdQe5VkJGrK6jzYg3Lu43g+ZpgJZhV9fVQN+CGxJZq
+FiiSWG6GeZq3WRIDFK/UPjcXQFCDQ2MA7qirlkI+3FVzexhzLYsiiJPkHjd2uD6sxtaWXwqf+Oj
hUJge2bVp3K0IfIWT263B+HXisd9Txr0GPwZIMBUt2tLSn1u8+UtEbD843qVlI+y1mxOZ+hcXZHE
s+Pk4rOHD99Si8I4J20hrBd7AL3qNLprogEtQh/jxvzuL8Y25AnZcMiMWHCFKx/mSHFoimxApNi5
sXKLANHbOcxOCmWqUvPobAP2SdP6gZHvIlu5eKjzH03ioHdgiDRw8u9anqBHoeYidMMYYViMjOag
2kMiZOQgbqyLbzdwAdvQxwu/IEocsLarVXcYnOkjbV38wLkOTZQOjYIdJzpG8BpkYscj5Vmf4k7r
25tAT9uKAh37tbWTEOUTdaY+rG0Th8gUhti8jI4Rwx2aAYNNV3L5nO7vUjKGDwVNwhK4VDuEsJp+
3MhAIHe/hFKTDMi4tCfLYEdU/UUdEeciwv5QbYFQ/nJHvwkGdTjdG1m0F3Or6kcrCUMJWvKwPKxZ
EDwQu6MIwYTtuJYrMQGltQPJblu2/sPTQzmGVXnqxoq8zPT5peQ0k4TuR5OZzcFHI/LEaWwiwxIi
FXmSJ6MET07anIddcREq7es/Oe+NHSvtereV/DyZdu3AuLiaOH4BVwovoE9BhmbcSJi37Aduf6h7
mHJsGLz5LeRF0dSiFDlZrJwcDPGkwB1cl+FmXvxVFA5ntI2LHOplofE3AZ+MIQWHMI3uWdcp+U7J
kOvOtLm8rD6jNJr17k6fiDCm47FzoxtW1xAi+ZjO0jlue3cZ5lYukszzg/RNBA+eOTfPxYT8wjBY
9Htz455RHy9DQpUnnnFR2L3i+JcLJr4js02Lw6U7zVBIN5Dk38rCNRWoTw0GQBagHog5fNIHSiJR
/SRSznocqR7+ibjeEyaEyRq0vOAQH5UfW7xhSS7mP25WN/sRoF45UlcxMH+cAfLNVnYwuqaG9vrT
hG60pgBCGTnt5obGNjZbGzRsXOlV5LdaUEiid+vOZ9KI8hsJCSfil+jJNrG6ljS2jHBaOfm77t6Z
5tpdFwe6y6wPg2pp/f759hTIvglh2BQp8CfA8h4xtHEJcblvm82MC0hVlZu+hOIf7Ujc2ZzR9j3l
Rse3uLpM0qZzMxxZQ2k0rhQCeUPJay3alchcdj208xkygpL8MEd5cvTd1gReT5fKHU6p/og/PEg8
kVATsrrWovwRxRyG7ABA8tfgpkHC/5hwwy3YbTMKaHpdhelTgFWzFKpDjUWhORsdSGyUMa90F0+j
ZeZAPE7rHI5usKB+dby/axr1wtwAUTuDbk7H0TR23G9mru5P+LDmljQnGeQwWespgUPN2dVYfNSY
bdBOdeUoCIK+YE/t6lLRizw68cXiQI0fp4NXKsWvf4wuh2nMjNUCgE4oC3218unGkGacdcv2dItD
vb9jm+zxpqWZE3xCRgAJ3CmJ+qLWOVNuriEIGMTnypEiL90coHxznUA7YJ/msD1B4VlcnQgTmrLy
U+TRXRLygHWHq4ewV53ELCeNLKjGd+S0QWABPFV1yg6HJev0dgJnmuJ+jU6yQXBvUfTTeGHUmRui
awB9eFCM3LPbTPQckBSXuBU7d+3YL+/whdh35s1MG6ioHehuT6P+X+MSuVAgTiVMB3n/fP5yhtez
JtBPki2UQaX7mmIw6UIgqR9jjIci6WIVotRLHeshvAlEnm/BEhKZN1bWvQJecXASfBie3/biLST+
43nuOiLN+NrXjLPDG/LJfe9csbCmWNBXywKQpZbvuvMAVDaiHb1N0rCZ2IJBTP3mjXtOtomfKr5X
mgMBkbWnvWAVSYFvdz8HRnGEaSCU2PFrALYEYswazQ1MKcSocT24YV87IJS+eq6XJ+M59l2yziOc
QICVTAh6sJPseJv1l2p44gpSMYAFLI6FK0BJ3Z6xwemDahO9SYtWCrL1S3LoS5IW8Z2wwz4qENFs
cxC5DLmUq+uUoQkDezSLzbS/kOqq/Ltp97Q80YINno/alRMeWjjXV3ljAnY+eT9Kwm00noFOoT9n
ERtFtrDfDTk8NFgbatbNoXCLlnFpGY/D7xbRp2737K4BJdD0jQqG44p12k1Um7oRTvRpawV8ISgk
9eGjPKPbfMyrzGK9kOkPltY65Ic+Rp/+gnel6Tk1MiU2SLL5AH42yVVyt+vsp0zZ1/NiiNuRlrdT
XAPMjjrsOAMTvLhpyUudrDE+8rlLwxihygftLI4/Ou8SgXb+sj+h9Bx019vzWaEHI6XuhiiwLeZB
E+8k6GMUz4+qMbrGBHEanVhQ9Xt0xSfDaAB/4WoSMXq0KIYejrjCLdXbQN9/sjrOTOQ74mVzINzF
/5HexV01wTV3oj7ZcDenJVlghQTScr/XdZoTstTGseZhiXBdPQGXwm/ZLPtVbMjiEiR2GvS9aSjv
K0waxzQPrnOFUB8CzEFPOj1/j5QhQtxH0V86SyVmkoo9fdPLY3awd1zAwsOW8z3uUsCNdCkNlvUL
+d3aplhyAH9FdbthocRUqJ5NMwXfHnA30or4JvmylpcYa1j0dzbbCZMLPtfyJJ6gzD6l/oqzUJK9
Ah8SRZGdwms0CQW8uatCPVtBUWUJCnxluKy/4HFYZzqH/97L8RqjIUy0b4AUINTkXfqYoHq3u7eu
qW7aofytBtHoIfJzK5YSIP9GHs6lDEdX6OAW3VBRf5EnswBwK5k7zWxJHRG5akA1s+a9AiR24mbM
3f+aTHYXc/vj3kt1nTOPjyOkLzNkBEbl5iE74re4IYUrDaJlvvj9EsgG98v9vGGEwN6NKGaEMmdO
wnPI/CNV0HhfcXWAfusJMoMruzCpJ06GyjdVR4OqHiI3KbznqgwJKJWVE4k/zvyaQ9TcFZlsx3iQ
TUcJNe3SNnJJAhrgVCRmhv7eF9sWHlDUsA2lh+lgWFS3sMfG1YkhzRaEdi8xu2Hjqe+eh2DNFBH/
YrqWnS5AEueYFn6tiewsZ5ie4Jde6jjvgVpMNmr/RcGGcB1Kp4tTVUXk7Nwg60MR1qPXRL4S/y82
z5KNezS6PzcQyFS0zlHAAm2qYj/YmXRx822bW6yZFuDkK+GI6HfXUf+o+IROOlEMh98HB+kOVOE7
OXwIAPJn+l/jwxTAM8tfd2v1zXVaMOj+Hp9ml5tSPixYhWJ86XQKGfAbdGbCvs5c3mGfV8CQVZKF
9ozyWxptyVig8yr2FqBNd80XY5RrvMRJ8V04awqXcb4l6VXilV5CY2r7oV6OALHkOdBve9Hw9Ll2
5ly4Km+7Po7vQbV4Dl9KR6HBxHKXDByd+ZC5h6OLB/4oSse3znmCKl+EbaNi8k6P8fHEM2UxJhyb
p1Gs1xcvtFGR1P+yvdf8nRXJ9ZjtYwxQIZxRh9eLYFu0Bf9kqBQsH+AU3lRkhn7U/U+j9gKGDhbo
WwCwo8D8oGrbxvetneitPNQB3BitPIJufD51VI6zo5W9AWV3BQ42N/hE4h2ANfze4TGgOWSjbFEF
xkG6HUbjmiCM6IQBVVMbHKLUPICg6A3YNFtQ7fztJgllGbB9oVtP1fP//nhxXPAcK1XICJwtZxl4
FQ9kjAw7n8zNOMsLov/YDgDVNAa3cPlzPUr9aLLAnINo5pW97XFOFeZPBKQvMi/g7pZxoEzxDTmP
6iRX7zJ3Z6f6v3BTqg/A+vnAx2MM9un5zqYV50HKuydS4vaBqpbPWiUnZQVx0P62egigRdDTF2P3
1dOhaE5T5yKUrC6lX8KDaCQ/R/XpRjLpxF2SZSdjuPzJlNCmx1p0zBzQlWe5sXWgnQJDPOZCyvLd
dDS47V0KNpXCd8MklZ3FYSvk/Yo0j1FxW2oZcYD2YT5Gf2sTJpeGiIhA1EL/Cs5vo9SHJTAo5YEq
cX1yeqGU8Fyeii2TvPqbdeV5UHuc6t7vGbfxtA9pauCe/GjB3COQivYzhqJ/4GhGQlMHyrj6xJAX
+Tijens6Xa+BSQ7qnJ7R4cSKsJrEMs54rUR386b78nT8stKIzuwHCO8vwQrhfIgR4t0a6SmhZFz5
ibe2gzZsuCWKMOABCk8Vxm/44aW/mu9JBxMXohJ02nm0tynJin6iZgCTn1yLsIaFd2+QycGMS5fs
L+9vkgESoY38qaV0viHtut9bCOH6RwiKPg8JJeppZrWH6GABhqIWH+zd8E/0J3dowM63r9LyR/xM
itfZ2p+hnGxjCoWmCoFBIdq4mk8i/y0+/jXvNWV5R6fiS2eg92TJCgixqH3cN4cnT8A7iZxKDiVG
fGm9j5kY+hRBSCWLL9wxCzgTlLzUSNaXpdckRLPVxvuRmJGVU9oTp3Ezj/k00UlYA3tZcqt9HV3w
/eThI9AYZzBDTI1mAG5jWMBI/1NfqnJZCIZh3WSnqs/Qvsuq8+ZUOEvAorTu2W7UzGy5cOZaMyuS
3tJqsaAaUjbJlxm/HlILLcg1i87o57i8dr+tfdEoS9O0Ph5fBvrwzZlcWHFXjTyv+PPkhvQoAlCN
WUam1GBIMWZ/6uP2Un8bBb9xsqngKAOmC53aGN73frupR+sOxIKvTOUa27bE4TIEKTGDHMsJZGqE
8orE6YnahmbKO2woaqEMaF/b7mCkgbJP5ZoB2VNTD8zLTr0zXZWIvJ461HqDnuC0EdsO6che8D1b
qHXYuDQEO0TuqDimcHtt8zTtLhd/bXYb2wpuw7c2J09bwnO4C46HjDK37236TdD4HGcKB7gI84cw
TuqSUctrcRflDpTW1TlWArxzReTgsLVsFZLXZW7dWDypUcYskfIHTwi6jJVGnNpnYawGwJaxo6Tt
dP0fFILhS9A0LHT1nHtp83BUQKxTRc/+Z8IjcLq2u4qFDzOIDFIvma/m7u+ThLPjXZ4ouxCKNf7v
K2F9+FZlQpPsDLZctYPzq8z8rZUXrjSOb9giRWdg//PaIMUlTBK1TNOp2PojIJ6SbxMHGl4b/Wy2
RTFkmNXyzd8QByEQxPzrHXSAjyjM7COn/jgWIaL8kFlcSv74EwWikg1LE6kfq11KsJcnLc3EqM5K
/kSBzkzWbCnFvglbgab6xxD+e0bNAqmqfRwal1rPFadtwEJ++EqPE147lYNMh5s5w490d7IA1Urd
+gUpQF+vIv2uBOFBCTy7eJH9OIrT5+CMfqKzE4/k/tuaGPjrcCZ0tU8jsF/L4630jiswSpsY9zJO
GQjxq9eovZgqgcmIqUDN/gwBqX4y7Td4IYHVY/kdhTQLpZM6Ims30BoWp5cp+GeAV+oaljHKqQJ9
DGr4ISzlBs+L3BKgfHwkUEpZ+IBQ1fEN4lp4c+JQHFT2ELijXasAnYWtv1OgeNdkM4XuRTR53T7d
0GibE8Sudb5mYhgjwpaK+l9q8JRdUWCBr6rSkD72ANK0r0GIYQHxDLfWZEjEjzqYkKDmcIhbTJn7
Vx2zoJvluPybe6dixVIGEOHWVX6XjQ9sv/zmouMqJxqSpOQVDRMD/RXf35ZN8jDtnjf8POA7hMgQ
pHowTf/5O2tpZXMcPG/wRbm1xTrFhEBWIP5hDps/vOZS0wLOunByet3+IxdYPyesjl0WoPC6JpW/
jc2DjdkKfyjQlb8EPPiQcBH0GATfb/DoJjjlEdD2USc3c479+L2tQ+j63BlXyH1SW/runIxekTCO
gxczjqI1FoiEkHx/7BsOzmXxERKtdG1p2En69rZSroqa/uPVodTbEFnL+6rR1iXZ7XS0DlrYhWOU
CRuKT+88sUIat9yqsd1mSDkyoNRskI6z/dmYQwe+fGQPs7niOo4opDEtFTOSZfBvVbwwKr+UPOEz
NR8xxq+eRr3/AI4K3MfTAHzPwGMMxNFW4QZh1Tz8/WR0W+grA8LTlxcollqWKxfJRi3XLVSlI3tu
OgqdJxMIrPbzYYH2Vk3iN40eo879eg+jm3pfjdGN47wuV9QOtZuvkdTwc2zj/KlBsnBy9BHPic1+
j2OALI9fV2IUqKwkhuFtxM1RLMjxam+WhL2pTNaRPLgzPRwxL1e2Q77HzwbCFnzXrwBlZuDQMcmh
pB6pJxZHlfb9Te8Qj/5i2JRvzX8IMdQJpsmjjpT8H4uJ+3dMebhR0DiJ61B8/wc2G9py7Y1xtZlT
M3PQboKdPF7d3gXySut8zLByUSQOtxlKr41tNEV7kc47K/1SkRSJ6yzKR2owUrgKT6tG4/La7cDu
2tdPc8LllBgNxlUVng1QSmsRU0j4UjIoYJImvWromjksAQep43kLgZWBo8UvRKcofGD2N6K3NgaI
6VxMckYQDyLsj7IBRzjOXL8WvSueIYd1hsFn36p1qROf36HOIpkfgBoV5GYeM5kfPKspI3H2KuJ3
iChW9OvjrVXwe0LsO16peT76rnn463ihW0zr5qvPlrh8vcJWvoyeiwP8FQPF+Wy+E3w9Nb7e+5f2
rLyawdU1ytsAOI7j2lo5X8aqrth9afbhkqZL70sgVdmnrDirggxyit7kIWjOYIVzjRYuB0yUUrnI
gAjc2sM+CHlCc2T4ElF1kDMTDlG2l/SDXDJ7C2LiQjzLlURESjz+e2lGQ7iRqNLfZPsGBQoafm8P
ZVVYLaPTPDYyLqsxcYGvU4DKwnuaNSJdWV/9rSHVraZpQ8l1ahsB9eg/a5uBP83pvyzZnA6Gf6/I
MDjwAzpqnbX0Haf8kTn9eR4mfdJU8Sa5q8HvvPDvL0AW5eLc9oaV68LOpS3yIprzI4Pa/DKWLiOH
rbp9egbSilc3nGBrwPfkxqkDIJ1P9KonparA0Lugujq0jyCjv4ctmjfdI1QVL6x/aEcRMTzenWXq
2FeinAyaVg1Ojy0QQppSECyWg0yZi0t3M5Z1c85MsWOndu2Gk6WaPY9YPFfK2208MvgIwf/1Jz8Z
dDD6LEP3t3P/roatbWfqYCBalFzwqaKyO1uBZ5inF8PSDIvrCrfXWGTjVe3CPApnDAqfnC4r1HEk
BMUzGSgQ9EcFfJCkatB3mQuw6WM4H6I4XIIqPMiOt+AQBTFwxQohmhQ7W3/eD6A/ukqw8OE4V2Dn
2BWrDy2VUjsh3PAjTD99hgD69rgXPAQzYUgrfwpoFcc1R3yL6U6KoG0rEg0jz677D0nuTdudWkZ0
pdLb7FEdTEPCSlQVzcJgOdr4IM/u4f83dsUzqpP8W4EwVT+TMSlwGJKfcm7ECOQMa4ZM5lRYJ+Vd
QuBPXes/u+EYl+Gf1kKD3314C++6ajDNpWcpJ7h2snzJuvGMCtW+gdyoTIHgOxu2DSFoYxWBRjzj
j8P4KQesewwPCO6l8SfdxAY5ZosS05+V0us1Eqz0tFzdRMdjVW7I87a/cGiANn+NBum1JsKnHJIR
Hwi/9Yi2j31qXN4p4U5ocn3lbPHH3lWll2v16gidQyxhjyRp0HqUUU92U/CWZ+ANXct+p4+k1bN/
pCsEjG46nUcoAs0K4suhqGO5upZGqBWJEaUl/cqHe+bak2wsbZlEZG+xKfCWpqzJrYHaSi59l6wO
2DfflPiAdkVMZXcD7BcPIGDC2vZLM2jIF+3gsXxyxLbC/HufrdnRrtxx5vNYVlyuMjObbYscsVqD
80rvwk/1L7VH80Fm7SDbklF66XPBKFwLQJpbZXbpcArGurdFnQuEyCfkFsMya/AjS7rSjtj8QXzX
wASkhMXIOi9FXStvoh18APyq+3hAljzz88qtVDiWCHvtSD1kbHIpGP+vRfRPm40/wirH9lX+/7EY
s0bmW9/C9Kw4hMNyay8qWMYfcyfdl+xWf8hQCydVN9Rj+7TX5uJ9Ic8OP+7zJiQ7b3JLy01J3XCb
qUP0+1dlLyimpOrbMDEC0sSufIYDLpQb97iddX6imzOF/+0XN+aKrXMxdPpw+4h0pMF7ogjtm7n6
T1ZmpQ55VPjFesFMfhrpJFCps1E2cKX0TPluYYApnYlzyogN7seXZ0h+Tr+s3/KrrUCR3nzY+F7f
YLOjOFv3ZCX6GBW78hZLZ6OViw0ALqd9CZWrSDgggz3UE5nh/EiNosyBBaYBue71EtYV1/MfHwXU
Ecx9gfIqbM+IcFgTNxuyB/4q1V+UGmXCzfOf3uNielkXk1oNe1AB0ko736INc+NmLJq2LZQQJgzc
heIeSe2IYNg+al1x0ecjlqX1efbntZrCd+jnNcYqdbLXRHUqEUCzjqza/RhyTeD3noqfqG6b/hgq
2KFrXP0OyROgncgbnEYpj0h118BpQ54WqQYcOSJJmSsrpv3MOXbUL+9B2UqTOEL6bR7ybtKDy1BB
Ptg04Q9uwYtX1PuMrXzOwgU9NYQzqcKxesxhxQHjR6WybfjuBRfuiELJoIkUUZ8mAU6Cm7WwOnLk
xjwktnYuAujK1+mMZXyEEtzjSiAfeLPaUEjFN0ySJ/y2oTgKDngR2CYhMOP1BZEbXQBnrsrfX4t/
Qkgzp8yg5CCXnGYh/UHIRwPWoxhuUxQ/UjhJRkQ0Q/sJOaKO/Xyy1MKzI2vnsfWEeA7bFLglLwk8
19fHdQGxCa/OvFtGfbo+cMsfYiLj6CpS+K8SLD+nyb0fghl+8Mh1gk9vbGFWKnqe/ts/nMn/kZjm
f3bL6I6otI/3Nqn0p+6m6YqgK0JCShWYTPS0CCXkfs1tmvKDB5urYIPPtW9tUa+M+BSZi0D/SAf2
UZ56Gy/odpSou2QAeXkpBmdTriah86K8HzYSgQjRAYv2AXV7Mm2Z8OVRQTeDiMi/sFUAxGTRcXgG
oGNUTEL73/N3utgJHVwMBmXbXvuQcDU7hpymPAMUcJf7INT9pLq5nQOh5VDMC45wviLNdizuA+oC
CJ9qNmcH6A6GHTVNJRisLOde8OnfkjXq5uXh00OzyWLNiRfTu1SQttXQAmR6D1U552+WicfN2cn+
vnwpp3NohLlch88z4Qk2mmPIBVvGPhkbnLYfS0wnWji586lcLxVUi8AFN/Jq1TXmGExJuj00FeCG
pv7zL1tYXVj7V1KnA/i7TuPsheWjXjv6XwIXlyu9OkcgDadDY1g+htohJg4+0Wq5yxtdFk59uBQ/
a1i/7A3ZoRlikbr0QoAXbJVv1uXb9aLsyxT4IQFaZ69quH2mLMSyTKQp8m8PbHJCASG+SOSzG3Uf
T0uBsQokAZuPMxMG2eDjwmmkE2Gh4AhaQW9EC+sIlwGnxFLsMiapJbMKyAgNyH3P9iwf4LLgjKSh
PMp7U+4WHeC7nIaoTs44GTLV01hPTX53ZdaC6EMpoJX7rwRlAF8tGXB9SH5x1OouHV+s3bAxQiPX
AeypjkIaNjpfPbMOu2mAiuX4871O831r2lZVESh74S27MRHj25dMB38UKKj0qteM5qBTF+rfq8Sz
v7OEXj4MlOanHJ9i7jF8jr4UimeGazt4L8mJ4XZW55bvhWsVEwJfag+1P9YTgVbl6SEz2M4Ox7Ye
SjEEheJw5zGZFAHhW72fKqYL+voyUVzHkmN6edcZmgv5OaE0Nvl+T00xJZi6J48Vnl3YCajsmiN1
Z1fKmlezMyitxMXh7RMozp7BOzdj3wNavWzwIy/lN/iTGXW6iayJNGriB5CL0IKJFC8uYGl3pnWC
HhvZ+4Li/Wxd+Iw326wyo9tWMewabNva4izteQZRL3OdxQEbdEWdbpGEkYLlxVvHpzhKc2w0/HaW
Ngf2UgSrRQiqhmJ843VoojUkGkv6o8/aLgrcYO4Z8KocI/wUgnzAddIf9g+crYcbpRoS6MVWd6lH
Pn5XVdjB8dAo9GvELuuZKXCI8lxdnBU8jaVnzuP7+SxOfHAnk9u3+ZsvPX6ny46HOFPmIUD3i9t0
CTfvlKKE9EMJ0wEo1CMAQZ+dlxNsy1CF0Td5pXWc7dwu1wmjF+EU+jcQ5FiXbVXUC2673ztAKaLW
B9nMb2IjoMMSnrOgmtvV3Tds6/KEFjQlGF+46M1XCgMgSbEi3kVmIcSF59tX9cNDVFIgKPyU/oew
wP4JDUstcTz3P55qMLevip1gDO1IfdBXsfgd2SsHOC6D8LutzWyR0Mab6Fl387XvyTcgB+dQC23l
GtLCS04QS53XPqtganaBFgWAa/b/NDT+8FMMxaTB5LtkTGSPV3meRhJpOEKfdLvAy17mL8bY87Ub
IepVPcEzX7j4Si305s5HSUDsDVg6GVxn1k0O4X3fXuEesmyPDaIs8KuaMccF9WEGyjurv0A7GZ8m
ZLu0YmjX7FgSmElebR2qFCiqHnGVF0/kKAtutOqqn3GffdIixLWVAONLbrWFiBuWV/F2l5sd4YJ0
Z/Owyqg3D4OOWKJgLGTBvKgUvTeyAMLhFPiwYzU3Q4vA6BwaOtkk6jGuiIIHjSaqdbpvoUFRb+mM
+ZiBmeLimEInnEBUeWyWs6pMjvEJsSVF6bW0MrrkOQ/QJAlAPJaDN8DHf83i8rRXd5QS5Pe8TOWu
KO+Z/NzLAQIRpKtQEOWbe+JbiJHRHV6Cro2OIZSKaKaT6zNWp7KRA4h9baspmkwUyEeRktmKya0x
cFS5O2i082PkLTA9kv9RiAM8Sg3yFaUzKVUchxJWpLYy4ch2k6idG3dSH1CZMhWv5F2VWMDWYoo1
oyaMPgpzO7Mbn8Mk4CuIGvToNwBNZpqq6aLh0OPvU/MZ4tOht690ZZu7yOLWCAqTSwKZxVeV2pO0
6xasykz8dSogJDrd0ykKxGig1ylU+m7EJaDS+R4g6fMjwLh4DOYjO/7gabntWlyn7IEAfSLkJSyQ
MyQOvePRbP6ZzMhZCfRA5NmN+5Y0feQ17TckWTaLGwRWm2Qh/I3k7hw4HH334uK+kNT+kSQLMSzh
x+EMOWl2b7YMJ8STOtr8AZNpRIEDuw8OnBvSh9EBUEs9EMRt30ieOqHDG24f6XieUxBnftVHsKrd
edQ1bdHnRmOmMDXCXbnRqGDRVu/EkocOvrz3WezZM3qaCMoYI/fJNIF1TmRAUoY2SgMcwUPGyDGw
iNy3JbQPcwrRiO/AWYWTtDKWkK5oBImSzPvBc/muWGjl/MwGH2wRwKDdeaoPseA/oizuwWZO5vjE
LqYi0W8YCJ678fsMnZL9KBtS03jdQnQ0uszanSorrC6XwtmPz7wSRGjp4SCOlRpxVyXWpVbshvgu
30TQHbyMod4zjGD1mpMs1NJFNisBMESNon82WqkNrlyTZ4FzRlzCnvalBo5Yy9gTqs39ILhcTYHM
p85oEBGg0K3Ighw1yhVip4qkiTFZfz17pxjFuDZRX2Ycq6H0WyQ5lWa8A4UsnQrvswJoN+El/m4+
7VSO45XO9PCo8QwCyrOC+a78tlEEHoxAXDTNyRQd20tTm3di+Y09r68cl/G7t+Ux3MciUmkK4Pqa
3ATYTZ8QcSF1Ng40sHMeRqPuszZ+/7dVDZfy/FaB/RZY76FnWpWO+dx5Zx9B+cDmLnDW6Q9FSozk
jagJtwD2TnUQCZ+if8l4o6PQ0BkqJy1gKT+GHSlqNuO9dvZ5P/IfM2cCqIvHrWEIJnvoJzESbtue
2jvP2KTklhhvH0dhZRxN7GQh6auSbpFEs2pcRT2Jxs58G2M5Ys6wJrm9Ia8kku9pqjeMge2bAyGu
nv3mnjMU/KiyAEs76mpnwTkwSdvmN9JPN03KvXhdq1KY1w8WwJgl732YErOYObyoj0yvb2is1UTl
bf7sCiCuYuM/WYjaqbCzGOsFNanEY6Rn4aRFEQI2BNwV974XDK+/P7jojduJiUzFajKGrfiYcoYu
jgGnBGOPl7djn7LstnvIwLHhepbxZDTGhz3Ci86YwC6Q4uoIOwx2hh6EDQJGWaVpwI34xCqy2c4v
ymFSte2YCteE3qubl9ECC78w2qykFfisbDYqTBsJvju/yeIMbqMqhmgnsFTMf28dCE2ma3fftJ4E
UTxHFQS9Du3P9HxlnXzv6v4fwSWZ6nrAGy4l9F53iFZvDfvdPzu07oJSKTKZ+cX5E0VgsIInlNI4
nkflYvWOK2dZ+hS6o8vA22JrFh2Uk2PDcdAzyb3jCahGezItDHJ6Qlmhcw7HFKeCFCsyYYA16hRn
n6CLioWCqoEu7R21ZP1OwnxOH5ivYY9cURU/DpgR81cVoqb+Im5IroaAGNxyrHVjNbieRI4/xEYM
q2wp7tX8Fwgxvvxj/Yj5KNMvWOxwVbB7XQILwyLKisBZ25XAbovmm0iZCSo6LuC+eXWSquZelWGC
d3W9in0ycaWDIX51yVYCF7xjBihlK9vEHF7xfrL2vX0F5z1T7zVzlnOlKWBI8e+tJc6D81Xu6og1
zF49YYYLeEPmK2KNHtYTv3wPdSNpUvAjjGFE9JdHULnh/tzQcmfnt+aBdCjOCGCBqs59pt9KbmeW
MooJWIvy2gdS9X5QRPde+X2ehiViqzXgA25/1+yE7omtvDCk07SdaUXUeu+Yl+QV3WeWXlQDUj98
Q2/069/1Mka4AN1oJPw6lhO+snccyJ/7Nv2jJzlPQ2XElOzcwTvTW/S6ZziYD1INw2lqbRPfOTqP
HPme56bG6UT4fhwKSGXBjV8Krkdwp2w7Xkwm8GGW66mdax/yY8pF1vISIPPXA9fSn7K0yydgEmfJ
Bh5+z8pBnmfSLCt+TqiNY24thJJJPulNK3DX/rv75pCLtUENB4lenEgLQEUxqmimNHtn9Cun+cnO
IK49PMhAal3Xg/bCKf9RHvh07EmdjJEuEva3Isjn7kYDI2K9eQTmnREgxiUFWFY4wEr7GXVy+uDD
LNBWzK1NfgUd0W2vz1ngZpelorFtx5RP5rICV4/ICmL3nW/cw6iaUQuFWiEvYlGLGMqp+DK2nFE7
UgmAEZ0RojKBZ/tERrCgLjWaOlMWJ0f7XxmUHyio6UxEm9g7G10qfgEfCO1W2nwhnxPidcxGwXgF
oUj9EINqOb2WB4zPxMucqKjT554vDn6KBZbkJHO6/sHq6YZ47zKbBx/eQTkS98RpsD/XfwDjq1on
qEnFA30jkfGkzVaGEZEq8XYuJyql0NVHWuXfBehskRF8/JScjVwfXyF4QAgSOWa46D9IpwHboALT
uPNJEP6LkQrC0P/Rna7XloDAZ1yBBf4QPj7dHgLN8J6lK+msRdP2oKtLQOILfUYmbToIobl9i+I2
CIs/JceykjBmeJdu7TBCKlI5D/c16J9OV9Oe01r9Z56cPIwBZgmXrc3OLmr0ICkeBdQIlfQQNmmA
vV/MJme0Ewpe4PkKeezpSoSx3KcPXAIgGKdrlqtEgHdSR3WVkOR98btV3IZFE0M8U32JbXI0VybT
V2BwHywhosII1L8QGwW/JHenImtJDIXxyqTheLORmByMq2KarNgfkSiX4LEhtveBonGhnrLBYgRr
LzwqPLwUdgCELKblAjBQ3qEJB881TXtVnU9wzsehgVykJJNE1j8iKBXI0tPaqL7KOoRHzev1gf/+
+J+EEpQo+dkRYfVfxkGEZZqg+mDVtPj2xzhwpiascYNsMTL/0IjWE2uk+fxgzrMrZYyefyiRdV48
3vDzIy0bTm0IpSSBkGnYeBEcZRs2/KQgHVH12bvSnuUITX4A7ypKCh71OnLKox5MbKw8PK8klchw
nNF3zQvAmw7DpGnOCWFlEbJJybHZNziL7yvcweW0i/XsizFwf7wZoHgwbrAZ/OP6UcdxiUWpuyRn
Gr3yRFtv/YbIx8SBicfrpzK7GWtUpiZVJDhE7/cSgIsz7s6wmtGc8fggfghBwXdvYhiYmd3z6zFZ
tXEvzNAOZL5eVYa+W8fvVEkfiiDTeiINrXk49Bm5qw+t6QVlYbkzwmExtnwoZGxSLH54752DVEKA
sxzCvpFzXgWKzHh1rkSaNORpN2hEn1t+SfzH4YX0FwbZBgbfBXTrR+OsKadZTk6XUGBvWpXy5o+e
iBKsnwVwUpy5/WKa0Hw91XsdapmLMO4H8GRZBhVEEaYRK27qrbV9dk45uxLrcUA6J2cpl3N21vZx
Ha5naBQwgGNBUiidmdIibDwCtWXi8vuq4wg0JCNOVPrh4Th/WCrCTWOECZ/TyG4nCg3DgiIrERvg
GMV6sdr8zYv1hs7qRMUZMMh71WyKbUe1cOcb5oRx5anJjZPcH7ssh0t9s+ECicQXmQK8ePkCgfC3
jfGH/wp9Tg55TEQO6atLWVHtCSEt/mZ+XMk3lng0K0YjXOSJhO/GC4515M95/tmqevZFJJXbVxEU
yH95U+7yBSNZ5/ciEbu41Du1X1tFk4O2eufZV0aJrbs39b97ZGOTw2HWJ4BQTM71bMRiY7EWlsz6
fK9i/QnYfQ324nJ4ovz2QxtVi1ZnZss926do57CJOoLfE+bjt5sASRRG0oNUoJNHzlPyl3s0aDgu
6/ixqma6oFiRo5ZlAjWtgRKqJ+/makTxsR0P26HY7t6p5gw1qozXFArmBrdBTGdgNOtXA8H2zIYv
ovyBq12ky0N68J4BWDcUh6ub291njKwcdbuM169FI1Qu0EA0t9/1NnMqw7AeWckrpqfgOf/iqaT4
swhy/Fi4/fwnak+nfzfSZ2m17PsNytaUCg+iayuuMsGV2lDzetsiFu3MUyPc9s32GULNwOhLlUrb
vxYJZE+546GRVzyzNDKHfH1JB66N8Qn/3QXFQXIMgTXtn1QsJkFXdmaLA9VOA3Kbo5QyIpoOuHaL
4/vGl0iTjhzw81zEydSs51nOCFAj7r9EsPCmHZaGgZ9Tb/HyOuOaPuw8ya7hfdjTKGb817EBwi2x
61Rtbcg5K9cxXBafBzvXA/3NC22Fxw5Lb4cfNqE7vEJEZlrV5tQR3sxDVegY5nEahetVn8/TD8dn
t7+FNkgOdvvqx1pSD+XuycoGzC2Zrf5tpgn9BOs305ExPsbWOGHxLWqVWjqdl9OXBNun2MAVVaMO
Gj0RWp3hn1sszjhND/+sqDnR9c72Yyu5vLEHpnuaUnZdxV/C/C0pxx4EdonRJ9DSr3U7Sdj0Cpgy
7qZQC3SKD725bWvwmyyn5aSxjME5lxyPNtl2gw0+/fdN2FpZc1CZgXBtOACunCAOVDdfKhI9QYe8
5xFAmxlpO7+jG/fqYQj3nsiR8SGcFAyEckvvj9kbW1E8cjqEQY8SQ6IYejjnwfHsJtquBgfBDn/7
nly8ia2AKbaer1kWXH+e8WeEyVIKa7z9vXvhY+5J86RaeJGu7pwIKcoE2bXPOtspHI8prXpCmuFS
OURFzsfifUmF1gQPhlOmHKYWCqMD4oUel5rlfUZUXolzotEh+eaoa4prRbr1m94v0Em8k8QTKvbw
L8MDjknUvR/bjrSpRWZHY5rYSlqOUObuG39aOF23cI1I3dp4nkuZ1diJOyd2LUV7fudfXMGvwdJA
dVGrxEhG0QlIVzR3MM3sl9hYVNkHBD0iERdKub77IV6gcC1EoZc+kSgTUKnN6pLCozsJhqRsDhts
Z9RjhpabGcbSleUIDyVXrkCohy3iIVtBBnixMb3XrqgYQf/wVcBzDI6ETiWP+fn0ZPetyPTpRThG
j5q6qPJjT7C/jVdipu/MU2CgDiDNLhAk2Pp1MwiLiRGpxBIFZQNLmV1r88hfJjfRsq7wNdti2Mlw
oLfhVTNT1bvq2cQ2AmYKaLxULQOPbFQ6PguIkswMHnzhO/VjlMmU3vmn5/SKgkPTedF6UAMkhhcm
jagKwUOsPJYC/gi1Yc4AxBAPc5QRrlqEk90uGaXQJpPoQg4tArH2ovo0BmmSqkWKwVMCzDjeMUO6
102/5MrZxgt0MfhjmKqP1IpEk/COsGO/AIGnHmhrTHJWtYjT1tuLlwjrP1ennyzIZXdtx/uGgnyS
92jBQQz5e6bSSMZcUgYQmtTfchblGXGFzpEqS6/g+SvOadO+b43tQky5Hd9s+NErWgCK1iMKkmLI
6PZRwJBr8wQYQSwC81++W/zURP8giyhUPjivMhm2QXZJxB5zqFi42iuqNdy3b2NCwfuE/fYTUYLn
wilAbqBw+YS7YdAp78nd9Dur9mFjB/UxaV5cjxSzHfuZz8n1iSn+yjHHfacZvloMNDhifYGpLVMh
EoLmrn6aP8fIxOqpsq0orICzzRsPeE0WE8B5/cnhvrjSMDE0khAnewhetpf161tvOXI2DdQgMBz3
BP1RhIrXywA/OcRU2+rcedA5E3j67I1ti34AP/AlU/CQpLD8gWvWX+Gew6tJ/iATtALkI7GK3i9z
u/verNqx644NcQACOHWVuqgEYbHlr9h77TkOtUp4hBaignzvKJqZo7bFcrtg1Y8hn/9WpM69LHqi
5RpHS3KiQ0MTAkzoBEgdK6kkStL7iZZ+sb9kGuz6ZQA4bKLZBPNGTFXwiHje2IDiyLRkIH0NE4f9
h7v8Ig6RohYYaJuOcqef0l/zKY2AvPrO66vdpg2R5Dd0CJ7hdCHNrdiwjpKZrCWf7kE2ci8XKXNl
sEv/IpoODNiNnFy3SgEoMKs+ajhim/XmjuGOc2761xd6/uBQCPdZROsJZm5hc5++wMWRa5PDnfB7
046oiEU6DRjjbCoxG3DQ3EgIpe9CRJxYOCyO1YCSleLWAZBd0ebD2xc5jys4uf6fDA7oFYBiqoQY
OHFekloARPQkuojyQvuYv8mfvIkeATHTp+Sy6BI114dXxGRRRiFlpcTI1PB2SmxQO+J65PjUfWDW
wdPnBXI3J7Kns3pWIcw9slSpuO1xjZEwPzfcse9/wQpYlLWJIEW+WdqjQdAQ5ybSGzQShqCrlML5
7VprKpX35tlj2I9DjkcU+gDMnvn2T/HYgth79CTnFIOt4WYffpqo7BJgaF9McmvHej88r6SHlaHP
r7Q7lgdoS7PtRI/Vts+bGJS8+q6MXZA0Yju4bBzm/v+hSSllrU1wMwDabNq8JL1qffmqKW6ZTf+L
2dTbG84Bh+6dSZUcszceo2VylOe+PRlsciNTaKw7AYhj/ykV2r2nQHA1TSFsRr8xluqnIT0Z6eGc
eThJ0DoWOC7HMLJSRBB7+8jDwuXZ1ByHY5SrZsN0KDg/UTL7Kd6HXw5M/LP18WBYU9ouHoB3sxTI
D1sIJJ8Jsesc4qZs2DF6E2ev0miMYYMe4G3ITWRFhLh8GeV2Dm3zZfJDJu3Wrg6761KPQTKnyIZt
KLUVaEJaXAfFc4UlJqOOOEbTEIF8SNvUq/TcKiilBsRl1ziftpExMyQGmG4Er+QT7UWZZYzelj7h
qKu2C1H0Kp2TsmLoc96fwbsy06kaJP/1BwHECeNMcuE2J89XsB5SIwf1nsSw+m68M2/by8ipSFuW
SNG8cXJwuC3t4pV1jxM0w2wkSQmzRn5m2/rD2lG/UUvcRCccsAFAMFj9z9R3+2+Zqe5EMyp7Q9G3
Bv2oUMsBkNIBO9u25veSJlYUj0+GuIt/F0vY4OzxkI1QU7eXlUV/amEApcLfZ72L2V4GiZ+rTg8n
s5Gmrx98oCaeOWl9iZnCvhPZ+6MTesxX1IhSSwyyzrkJRH4TpCp29HK332hNlNu+NEbJK4AR1NCO
Qfe+idvaMsqYW39D9U/mtZ7UX1uwmruNsfOYwQKIqwcltqWmL2FAyVTm8wcoWeycaBeJHHhN4Z6D
fVMlDFVOAq1WLRX1BT7RXSrXfCQlEuH+6LybpodsaysxxfDAFWPkypveZ1SaOcuG1tLvdBPQHQNM
AXdbkyJlZn6M8JztfUfR+S90ibGNU213jyWHgyWDtuvaQXeRgx531aVzkyLB/iQLqyiKSa6j/sW6
sIY61UmkUTEktOfSouIBdV9ALjEn3POCery5Dy0FljQqZNb1cQNmYgvEw8w7TEoWWfZHahyW5zMU
pd7R6A0lNkiU3/H/Syo2pkB8EMMf3TkduW+3/ZYpriCP0QBUkNv9ZVB3/XLmMOh7qLb/IEXVDujn
dKkiYOJfDQ8w/NbQ8+tgphLhHa6x1VN8ApG2lkYglGfSK6RXxgG77M8CNx/pBz3sE7v8JZAjGmuE
cR1Npn8IIzkvhq4/Gzdm19TRysPSSIZXzXp5y+/sCM5chGzlw3JLoMdFkbxHvpDEfNgO1jqZJWIP
NM/1VEglUK6++jl8hTS/NTqAOuszZ6iDpyNaBfm50NfIirnHB8MqAmSUb4TIvTXF/XYharjyLAVB
v22dtbwgIbQ87YO0F6wUh5nbICFXT53LpVnNJEOdj2saYrsk0oULTLR2ConrQBYrTe7UI0VZjLpm
9m9fZTbG1VVT+zDOG+uiJX0ZIJJzu40QreqTZqKwmW/Ww3ts02TfpOI4uD78aND9wr/MFkWJ6zR3
19HrovgeXwalAzO/0nF2tLk76xRzhx5YV2fHwgrxOYyEkOuSB3eg+XaChHjF/Y7uV7OpR8cZMUZu
UcHuLHr/XTHhD+bAhuLJI8UKuiTIYvpDDF5VwqaqLs+1oeoVjeKsHoU/x6G4prnA5uxQRvtFyHYS
7nfnmKuAbwiwgzTonYVgPsZJ2cyMVAYzv1atGEIggRGmyiGAYMHEWZsBhnrAdDyfCK9Qg+cvDkY5
LkRTNP6t8C1rJCzCN9skKTjljhnCms2S8jHXBizHD1xJ80Mx3V8MykZ/COfYE1Qig7qKfJ8nd+fZ
VMXUC1Lo8LxlSqieiiaRGsY8k78szP+sP/90HnL11SmyWDPFlgcCeKpY+ghZQy5KUN9HAWGAlwv8
UNqtLVhqPqtYoXLgHVrRvvDCbEuMhUWlIWKBZ6x14arzreuJPZ739noR7Kqa8mMCb3jgm9Sf3IN9
2stPSi+cuAU8rCyUJm5GX0GbFrdatUsBKvpy7ioYHDz2FbMbBkWDoS5kPyQdv0uKyPv5cGhGUC5k
B3z9nD2XsyQRpPa4jar1eZWkRGw0njlo34bvgyKp1rbcLbOkfaUoXMYD/75Xh9p6AsgIuUuhV/zy
X2fX13sNYSaaqMNe/BDbW5Tfyr5EyuWPU6bYxmYU13o3PtAtlFFoB7mGVMdFC6hlVcTZcSYRj+7/
Pf7wEaAwksIJQbvxQy9d99+BjmE/ds7VZdx2+oCfo1xISPKe3KSZU21NGA8OdHLM4KWEa0jD0Xc3
DDhkf9Cum5Z6W2XKI42DMmbPyM5CgOaumVWa5dKlinN7/8BV+ZydC3cwzs5qhJLR5iVgD/smUjCe
IkQyK4AxZKQm15rQbnVcnABF/5T5e/LzXfVXbvwS5tncGzriLGrDgncToAkcDu3FXiGB15vjRt/B
pxy9rjGJHxpYXraYWKOVAGZNwLxe5BvCW6gDerSMVEbgM0IjndgS7FAiPzU2sqCGuanEiM6IrZ5C
y8bJRB4LKz4xEjgq6ncj5H/Oj75xbFSS0qBFsLcA1KiF2mxMFc8e92k3N6Qg/qhsMyFXZkDBsJlB
0OvJ07PJZCcjqidLbEWk93hhMgAuaV4ou8b+hGOYuneqMvTUKe9MavSQgZSAvmTbZIWyn7IpSwuH
1vwkccyG/7CG/pCcYjo2kcQmo5Ei0fLr3oIZz8qxjZwhlzNiTKUfOryILI8t82XgLpM2T0aYjovu
e5Qja5xDeSZ2+83+9aLM2iEiIGJl6Tce+zLaXvsJJP56UCIYC/9FtuhBs+I+H6Yzo7yFDfVHG8bI
Lm5MJlLK6P3ZU01TJsD04wpvhuhiC67YIOo9/V3hSNqj+XYlgj0krIppRfg9Hr0cdF5ZCMLQApjm
nc/7P7m1czKaKXhUyq02Ec/mUOC8p8+EJ5oIyGyTyZYI24asUJryL9zYlp0Xtot7eCVqidGSUDnj
OG/Nu/izyYPowNCGSy1sjxML8/+pfU8XkzpNpeXLtefB4/ThKTpa9SWEaMMVS6aBFU6V/uUHgQZg
PYObM8dhP8ZGdIEyuhe60nNIcYuB6jGvnKystw/MUKYV5OIDzpOsp1Iu1n6FtSEd2na+lOv3B4co
jdaQweUMirG3dhJ052qqQHXaJgjZyYbVNZd3zwiz022IPDM1ZqzztfyCo9WkqiKTd71XfIJ9knr5
AIAS8by5Xn2fQ+4l+cH9Pzhh6XyUjld9X/nS0CWoQcC50RM8/DU8fnE9zRky6zvlpiHSaFJBE6oW
YEsrFRhnzR23dauklxarZQXymR7JfHL6DTqt6yL5Bmlp1b9oaJ8TsFW0vwT+xhOtebD+6FJfLgoJ
Jh3CNeHDByDGA1FenqKN6tsxsliMJtV8Mpvhok0nImBvyX15JPyCP0e98k5+/ZZuWv5jFYFNuiT+
rmFf1aWdZg2x526R3enSCOxyubf8F1Vd8fU3NVHyqvL3TJ4nniFeXk7gmky2EJoyhrIZKorVjlLg
vxRUyFHjyx8OO+n/Jmabh3g+2e8hRwg/6QjJwRxM38PDWjYPTAL+fv8/p/zJD19Js2NzOQr2YhJJ
Hp/PoypaAuNoGn6f5cdOLNcwJxSJ+bt4U/icUzB+sPA6Cu+LgE9laDEqv5X5+p4vkRohQdccPNQP
Mbdb0e9i0+m4HyCG7u4aVnxrmedvlH781VHHzyRfAstRd+3kVbdEEFtfI0wpbvYgXTCMIJDgV4Dz
D8bmM3fdHWUZ1qzTIiKZyeJNx+KiAPebwhXyGzvFNpkkL1j2due6intQC4FmejToqCNg8YtEG23y
EBwqvFrpYf8XQ9ykZIjwxarAsDpzuof01AvHT3OI0PMCjkUfFfkbUI0rIcZX3KN/qssukidhXkOu
34t9RsZqxGb8nroiXP9LO+kGpu00cnkVX+b0Pugi9LZWeJvsYOo8pEVwxghbbFY94HbRMchQX5ms
mMKTlleIDHvn2MljtzZ67nReUMy4+exnQoKGbe36PowbtFL44AyKONhLZURRf1S/mSzkFWWCSkbW
zJmfESYBMvRWzyoopecNyKM263kxRJ0RjLco1gV37OIlQr1hqTXkRf9zrdH8DFIMHHe5CNmSgnCr
89OVtNN1EVfsp38aX246JB/vF8CbZgemOrMr+R+mqokYfHHNuj9Bgth+K4QH6Nl0T3C7WfWlzBBz
803QZUoAP9mw31KNdVlnqFzLkCim11pt/2rQHdxLBgn19MGZelZdYZpI4/xCYI2/FOsl7kF1S6WU
9A+tarp9C1TuIL+tt6Apj4teg8OiYwqfnlA+HyawBCBYoVQS1OB4x05SkjirEcNGukk0uzBQUvuH
mEbrrUF9IK64GO3SVZVe+fponlqIDXlqtLyjA8x9waS4Ot16nOJyqSQI8LAsEsT/j0qsa47AyAB4
1eKs7UxRzo9RIIGx5FsD5kcKffEOlLyKW0BNBLuzOScCeA0d2dyuE+lmlQcYLCO+YG3eSCKkZR0f
zJJo+YrH9gt8EyQjjvCiyputK+KoJJyUZKLUgIgn+J9liLYvyQMnasmgA9uTysxZJ9n751FcBT0J
4bZ77ZxcgxydekMcnAyYXFwzhl39bgo0sGIXvukLJR4c4jkoQywdUYnrMr/RVFD0PRWxDpaBsiAK
ouX6D4FRffv1ATGnVUMnWHpYoGzsKm70DDh17RtdDVRzxIAPmRremN2eODeOjfInXLCDWyvR1anX
CpqfJ3Td/QWamqk89E5pMQ4et+SAqEKM/zgfp02DDOyc/B53+6AmaW91Bp+2rirfcYGy41KUWEsu
BIGhvSFQMiECSA7PTbDYEwZregPg+7JZnm4KmnV6bjeGhmYtLB/UcAJxUoMDJqGFI85WSTfAe2Wt
C3DjYmaL0769JDWX/XylMA3h9GhK8swwGm3y9c0DhvABmI9ffo6hkqybFJWzLFDPgyweGYUa1nyy
KMzxxwtPMMkgNDoeS7i2RGKkXElmNbgKcBlOQgPJsAheGeNmYOaIUK6/t7TAv+3H+gSIDfBJ/CM3
u8/zSbP1ohgAzMCfuLRyr9tyP9bwsGCXXkt9O1IjZrnaahrfVkZvrGX/u26KLoLg7LSmBet0BSBG
+Bio3lHXLfBaNipvIdnj6Q4/JsldntzxuJZjF1N0ODO7jGNtelRDv9JhKT9ShdmX6P0pPjvBGNu7
9AoeXxa6GypP1PC0MyXMqNrINyMtT4C9xeAOz1arR77JlAjoi5OyfehtsQHf5Hfju4nWG+vOezn6
5YzrEz8ctzt+h7xZGT5PBt2F/N3g0OQLh12ZA7Bx55ijSYXuzPhcbYtoWmqmm7GNc26jzXx3fd8m
SRixQqcCUnrc/WJdo3ysTEj42YMWGKp+Mzv6B427i6wVCFrtdZzGM5JGb7C1x8JITMwpPhyZ0JOc
ou+hcOHFCo5CvkRm34yOLROcFxOHurZBkiKIwZlskB477+RXshrjrMhEEqDrl7jpAzV8GT0h44N7
lyNRyT40FmEVmuNINOxn9ras+V+K4Qoa8ui1xF8wH394yi+AsWz49BobYz0mVnWZl7km+GQIXW9/
8Xbriq3ysSOo7mgqQ/AxrH0gnr1hL5IY3T3WgA3TOshG3rnWwY/mIQ1jvZ+ms5s4mMjlnWnSMNcY
FcEkK+59adLocPTaO2mZsvF8nV0qfijwaCMw3+7WoI2xisbFuNR7GpFQPwTLtj19aI8/uz2CGtKu
Ga4rGpEPxm4UesXUjX/9u1PLrN1zXBq3fsB7LYWtiVT//v+uWuTcbloMNRnxeetC2rhOMJkZRVBQ
7/MOX+ATOyMwOnEfttI/VY8VLTchwDb52jGCAKRECtRS1O+YfGSYG3jejmkAg09hAzY9r5ZoGsbl
Qel6FLj74TtigXDKnJNzdtbYMIFJimxPky+qFQc4bqgwtmaRby+8xAhQdOZuyg5mggI8sIZqOyPF
B9siAwk0QR7wVc7jgbTXJkwvlwwRxqnuCnEilDvD6Bc8KRBRO56GVWGVK8WU1fT7iFSJkgLdjC9y
thUB/yyofGnm5xJFIalH4gBD9iorzb8+JmyPROQCDoX9VaVeazV9hlgmep19UfWVN385/zMwJzJj
sGM2Wb3WvJ1nc9gm+7+IRKVEkM/lq3LBHPb2B7IYlACsmTb4AgKnheTRQcJeun8kjX1O9VqNJehB
xiIAccm4OrruMA9zJrRlJ+3VB39QIj6i8mS33QBJGktIupGSkB5UjYSEHkf8LvIN0c7crosr0/Fn
WNTRh4qRTNXsdtjga9pmyyZhtJv8QcZRL44JoJ+58PBOvKZRdtMZU5ZPb2ADkvfK7ywzVXAeYmW+
8WRnp4AskLq6R1WVJ7DlBJUtdf8iyCYOIgbV0hGYYSCiVqPVTf4ta4Kjyh2e/b3Dz69U2YCPvEhX
h5SjtWH9nsdGfdCo3Wc/QEVa+PrpQiixcZgvsDeZpxrTUTcoqb5kBaSWrfrd1GabMu+WukCaFgMO
dfe8V5qNhA4JPAOx9LZ4Ub3k8luluQsTRDMp7Gqqane08pRRWV7nRI8TQ0o7pK4+Q8WQ/D8esKni
WmS+wojez5Fxnjwyg4fgJMdE1nFstHPQuVLT9KFd2vnrXTJ8UHwGbYury021JuBhQ/297t9Om6zW
HMX5LZBSxaf4XpQwdI6+LqdKCX4Wlvv70WXoB6ThcQozkOufHxRAr0zUH11a9IajtRsIC0lwbxGv
5aIejbm8aWL2gS384pF7IrUlWt+Xu691/KP1oCx3gw1mWyvK231apsuvGlbP+24PQ83SFWdY60Ix
uO2qklj3xlZm61dms7NXtJqOHS3gB9DC2Q3Gy1RaHV3jMLDcj6GuZyJ2HLf//V8IjiHvbMddPC9o
CyWyvE7DU4KRUobrXRpHqZJNoOAffBeLoJC9UpcoqTNHJnZswVdZFa6CvHTiyjH3osU3mY0Q3iUq
PDkuKBdOv+Ke5RvpjTbB0G1L1dlRWUVeTPYiGWmSCDQIaZ58odOIr2WOXxB9pwkA3W19QUvRKzyZ
KzGIhc2e0XuLYKuHlgyCGvkAgZEeSbBZM7OeEJjGmFxfENXbMGNVmhrrvN9SzlqBfQd3Da7yH/kk
lTEvHkNNIUqIfiCn6OUri4kYYa0I5YfQGEMMTkPJYk+H2Ii0221PpX/7v3l8fke0QE4+b5tR3RqD
Z45ObToi5OMhUitz/KHKRUVGOR2//P+dg1Le7msYc6puGnrTdlPxXWl0s3rzC7/Pz9d8vjvI7Iwy
a1BbzmjLCnCNAuznFm5+gr31BtjjRpE13NrL2CKtSn4vjyvwT8sQh1ZgzXw6UOLs71GpMhJptAPj
Xw2ribVj+DlrxHgGMwmTg50rQ0N0ip5nA7NgELBywfDf6qt95x4HD0cdfyOZ6qxyc3yr+qu03Vsm
2BYYkCa8B6dt/bq0cTPEWInfQT62188zb384NLukbaeh/qD5ECaw1s1ve/wJMk9e4mRXBDDJvipG
vmO8C5Ee4f+nD16KgIY8O0FJNsxYRlGM+fhttfxCPDsXawsUpUDcXNd0icp4w+NCZPm9kPdodpIv
/agzPp2LXnUcxW0X6FAxmED3FjD8zXkkXpciYdheJ5KlRd3wN2ngA2OpQgGAx8bWb/k8rvOt4VBA
OrdmHQf9kMA0sY0lWW4K19YhJ2+feKYTfDbo6BrPnb0WwHU31V60+FTLJX091Li5vrXE5+514Bvi
QJvpgkw7NmEpak8kqwUejduOmhX476SbS3375TsacN7Piykt7VpPX1Ou49J286+qmHvgJ01Gwp4B
m9ecuuO4LqA7bDvSaIRHaIOvoe+W4iGscm5e+B8rs4jMc8ra9TT3RPAmiVKTWbDtcsFbupNAKkQ0
am2InX2Mi8YzWArLZ8Eb/FrDXuPpIyPvJkL2/ZYcKU4JB1IK57k5XnDUeKD+bJ9ex+D8m5IF8dhR
DNmwKSvEH7QbvmRjcKUVh1AKCFbofcaJMwOqCwUecOzylMcABkhegeqxRecsY1XAt9nmV8jM76GY
IwDqBuaFVfLAAQalZqRGyG/yAqYo10qGGop6gSgYA21sV1T2km9UTEzCGb+iIopETntFSMLSw2Br
c0B8qR+bMsmwEGvizPmhrOivLfJAWpYCfrfJ1hQWyXlRUeOortezj16HcA2btP5A0iaBHI0zpvIA
eQZhfqtzSTzg7mY6aqpKh7n7A8vvUVPadNAjqnnt0mmzAVmvL9wuxaqbUgp98vq5taIRi4nopNs3
YQIBWhaaERHLzt5NfifHmUnyb2oHyeEVBrbJghBkKPNsPupwPjkev4qbqlRNurHlHgsZmuANwUIC
MPA+iOQXl4hr4gfJAubambQcc2S70H8z+OIovSgu6RucjFxsOkXSRoizlyFf6sE/M0o1SFDkm5R6
kcDqyPKD3PT9L9mk/b+FcVtAr+jDyspdqKKhaFYVYWhjHHfv1hqGr1HQGDxPKGVOU7hJ1dsULiV/
LHvmyw4VV+PqPYMXy6z4fCBVjh+/shZ/HKCnpUVZegh/Cycp2hRRjCQcNGZNYN5wrPOLRVpx2aAP
Eb2rXYwY4UNuuCIp0fP9I6BuBsvXhhQwVyiNPPHbVuD4SRK+ChtUA7ppu32R0chR0CcyFUIJWLOH
/dyjn+vOZwenUpuS9Q4rLoW6Y/Sjj9s1WAtZP0JVu5x/tbOhqmNJH3RYXqi/hv0g5+rktU6xafsd
+XRU6t4P/OI/CG94GFWuQ+gxFiGlZu44XCmCCutkL158NI/RZceoEL+wlbAqvZ5B75jUkQJ5qOIG
nDLvVcMZ71R7ytz/gnAyah5ryMThAUTK+htTur8xq9kYAoeFIx5MM79hs+RR6seimdEYZVMOfcxy
r4UzROzHfV8jto7ufXr7PS1uoVjKps6CbrXU5TGXNeFZujHdCXGd2zEaafJbn96lO9jVIMbdA2xf
szubbj8cqXweJVeNg6gLEA0zQkNRyxI0RLRRWR+c/2S4JvJPKJcpHmMRe2TSCnb2p/k86ayXJHz7
zTzxp+dy+SoOK4Z8W2u7p/k2If5xyHVMa8cbZ1wRKKOAf9dcx+3b40HImrCBZMsFSpfWWjmfY0Tv
dVUUnDTpj9LpaJUPPDtTjcWcYv10VWIbtjQ3A35QxIOKC1O6m4Q3YNMGbdSkNzVRwqpPuGmEV1mq
iXfAKuTdL9555/6arZPEDW2++HS5O3DawpjlvXYBaJi+Tzb8B24mtMHfiNG0prBqdVDBTxKySEew
rtf8Jz28Iehmsibd2hIVrAWpi4a0LVwe0NhsSX8Ij6pohcK4TdjvdgSQcyzo9F/xdHK7ht53Bq0k
8Z530lvBLyOJ3NACjSoCGoNd90qNJpQFF+tKemrxmdEFZuGGsigQRS71dlhSxiHKhQbnONMNSrE4
8emhBdHOCutTLxnSXTq420VfAgJaU3iVJkzviUm4bzCqKsV5/9yS4TOPlcfbH2MTdNJ3+3AC6f1p
sGUELPNJyar4nm7MsYzFiIBD/UdMU5LNPc5Vq+uIKhMcMzVTLoad8S5JzYO3TAUA/CzI3r/ryjup
iaKiRIEKvOxIIKJTK034s0CcytSxEpumvLOTCUBK9DtXLE7gPG482x/6WakdNm8qADG3IfG3hLjL
KtdtwaLXUtyJtRxBGs1u8Pp+BzJqzaxxNmLs1KzYA3N3C9LqHhDj9s6rTA+87ABfnzTZmNIWczsZ
9nu0rxaR7QsWcY87cxQRVm00DBEWzR4gMBbzhi4IgG2VUgz8jlofvE9YHWktE1DLxSeP3KI3/5jL
W2qPpVAEw0oq5mr1IMWecBh0YK2/fydVVuDSFbx1wSEzDSGSYZEfxfua5m9UXnTVx5ambnSMy0sj
B9yL1UoHL9L+yVwydd2lB4FhNbsyISJcnZNZGHqrrMvKHSSf4FBHnWQQstyQ1A31XGu6p2w5Wo4U
ap8tblbtO7CpRZJijJU2hM8ohBHRUKvtLN0mfE8rJMfU3JyLQrBCcgMWcXhlc4iOSEA470WJE2O2
uOfM6S1t7TmfzhSLG4lcCOF/H0/WrUsM0oYvORwwcNo3dTPsy+spt+78KTIroPNeuNSresYlMD1u
Gw83700NGTteLiYsMT6HdSj7tkax7tuEWqDVs7AUd8aJWhsBbfI5G9GJKXwIEeaIhym1uPRUwEQP
UOUB54B/ZmSO00Qv4UaUNJy3wLIqA4/ApKmb71ubZ4tJv9SpCaBTHdCqlttG8Qb3lGWQEtvnK1k1
sUstQ1DPcExAeT+/7+QaZhm/JNI11Fc+h1mAjly2yjBBF9WmFtg1MixvoHz81pHqefgDbSk/tqrR
PhMsCxmNIohU5FcPjGfeZnhF4CkxHV3Mrt33QTrex02RPNCziFPx0HenrgobNz7yoMT/eVJ6uaAr
neHh767PST2Pf9/2mU8PAY5m5ueU89449eUaMo2cc3M3wlDrMwJ3kOF7onHjrlCAfuvCwJmymWl/
fV0f4orNFccD4aiUvr0E+SGhcNnIn2wspmy9P4PGJMQ2iTLiz134PteMIr6ZbKp5OTFKSrBrJ2sf
iZIN2hTVzYHhxbfm0/yzoEjHO8jJHm5XRiUxdyNOUFyaEYkrvtIrzd8WUwuQD4onPbmrWdyof4Wo
I0ltJqVNr+ccNBzwHsFsJjpVHfh0Pq3RsxaGEBRZXRx5KwlKY6l2qkeVWwDPRN9WAnsqontBFeBr
BUOOLBFPs5/KkzZuOAJ8Pg8nu+/Zkmx/z2C0efsyD4ohgZKcR0I0foCiGdMBjPrcyku3yR7LqNOJ
O+xaJ5fsyYN7W+oCRmLc1T8OP2QhvFGtNuN/8YbgrrobXGUzw9frz38UWE3U1NMy7qMBwuGcrGwp
TLMhyrI9l4qAhyj6XI4DQJAs7pOPEQhr/zhov7fRwMyw2Bj2TrRKGAPt6gqmQm0x0dBMmjUrSVSJ
6NPrAO341RN3G4QrMD497jFVecqTl/i+rxn9rkIDIA9fBKBhvxGxMS4BRqDWHZ8ydv8PhLsYjghS
tzxM4YPdmaxVs/4b+D3XszNZ60uHvIfOFvlxeGdYWAXoDXG1lszWKeT2/qoMMTWGdSxz9BbqoCr2
bGa3CEOKQYVOJGKsTHCShMNn0TpjVRGsB7XOIDsIag5rHARn6iVOpOMjPbmjVhk9Pryfc1YHP+U9
jbBvhKUsL8k0ltnQPmvcznfVyBOhXAfKkSF5bBDRnYBcFOBDmkRmFPZkVBvlCxzRGDZgXy6s12ok
M7fBXqpwmTCoRg/0XzatwWSFDVcm/9apyQMM5qccDlcTKfFCksIBMqjdjVojGUrWAaAjHjg2UToA
tK1P7hZKzRr2NbyVeaFdqQqSbpYmspbK2KRvDtk4YMjvcWeKUmxEDq6G1ZLXNxWvJWUG/6it+9dh
jLuNsXwJsKPX/w+3DLPmdAuKC9U21UnPITLEQPhHczt5GY80FemU4uYow9wqwisvy3BI0EBPOOxS
dJ/ATIiTHz9tJ2LaLoDQcek1g1FR8ZDDaL+XYEnguiAKjJ/raIhEDuz9Pq9wAum4Lnzf71TkajND
WPbuX/ZwqN/rXWu4whyIuFIZQHbjAI2761+qI4x6bcvKef2C1oldlWl5u4/ZB5JPpoJ6lV2RmBaW
GM9Hts/JuXNdlzIOQI2PMS/PkPsHBqtjdU9chiXXs0IzZAq7CfPIKm4pjCYLp9ULm+ray3p+WMuU
XxWH2KuN2arGTcbLia3TRGOCEsRBWd7pO3a/fawRvLKHtdC2i9WzlQlsgIrFlzxT4lpFS8ocdhWh
t3bSnG1JLwhgikDeSV7JDB+3GG1/1olzNozjvX4ufvmESDAfIwimA02YqqK8ztBDK0m/8O0s/YKM
sWhKHUgaxigLAJ2glQ55IjdYMmSTUGlRBN6Mrd8mkqKM20B+fgwZa0bdkZG8NS26RCj4jAXPDgLJ
znhXGrA9wNeQiFmeXOvk9309PLyyfxx0XBqhaKvO6KchrPR775z379/dzqkSHeT8QUw8QYJ/cPyA
vA7SAeazA3E0GnFQtfldGmr8PKb/r5MEphYl3JzfSAWFEUZU4YN/nuyyPEnbCG0H5tctawzQTsJv
5ZQsd+8qqWt4uFSRwJSGt6WowBA1KXUKCam+PXnIgtrRuhfgibHgf7LF2TnePd3gjTm8QreIxvl/
q2Ghsq3Bo0qpCmUzsS8bmz5NA2BsxAqnBHqVQ0WK7wAwD/F6PqlU17BhAtxg7McUzTmlHPMrCx6S
sdZMFyaIcimMrJcjvLeR85Xz+nSYm7zq7qn69K8KNi2/zrAQgQWyhJGuFjOjr3GAO6wFmz2CKu7e
nLVnSYmvtbAgxVcOqNluBlxJLdFiz/HKleLGmKQYi9v/6M2wmsBi8LaQs3GeixVJ9ZmuFpmyQ79I
7yU0U1LnM94NaAbiKDPaI/iWOoGrN5QHqM7aVQga/icxGKmRjl6Ejbxed+dB+bn5QB1Dtnn6ot+G
vBxdbUrz0lixo3vJ5z02k8BzbvvHzEZhbhPzyNN6l11EV/vTQGOgFAkrD7eZIkY3G2MsP2gOaFf/
QuOx9ee/H4McdfSSH+wuw9EguKc2y4t09PoMCerWO5YRuENZmEXFzBSgHQVp5VION1/mMdSHxgDQ
tzbOXYsa5Km3i/P7qO3ggBimUwRfj6opOxvHqveZ5WGibA5J8t8TkhysWx/SdM64ER7QRBuAQXwf
kINy4CAF18LPSrcIC3CI+Je3mg0DbP56CSeCU/zDqd4498WXicDeBFsQHLQXp6HfyyGQStlatKpN
f2MqnvfCM9VtMjL1PbRRWj9tN5kzByGuQurU29C1jpTgDxJbFv7xcFGiJzoj0h4fqLdLIO01bi3z
4IWC++QSkFYHPcR1u2QYZHvMLArZ5QbE6T0O41/oCq+seiexoz19TRvzSFNiwk4oKbii5KGVhpyx
q37AgEScUSBAepGVkwmLn2HjWK8TwrVkS8/g/2UjZxwLapeezo0q7IxJqAP1ixAyldjE7dVE7tf7
lQb9aWaYt7KR+uYA96xI0bTgvBsbZA18yxFFEJ2DetV17/D2Z/GfkeqZ8Ee06H+tZ11/cSOQ2T1C
vhon0WN1six+MSksTlYPBIKtOE68lh00ujI5iKUTFEumESA7+GZNqYDm6RGOyJns8vGsV1XmImb3
6LRD1EQmuBOFRU7U7zxPijCVUBnAYkncrrWNjfwNw9vA5+i1IbjhzR+lhi7oRQ1daUD8S4ZBbp5a
HdYNtTPV6iREzdyU4MVC2CHTfIbt2OMfvLx5h4OVDAEXw+OQ/IlUsYbkLPKNlBtoVKIveCyD32T/
XQflbCKNSNS9QB0lKpa6ikvGAA2SX5l/55IFQjSSaInZfTWa97RPvOFFYj+VhlFkjcj2CwbDbTgi
yXjGBbvxZ7MzlzNAqH45G+kQ7UacSc8C865wLGGCTC39HVu20ziSxhm8gbn9EywGYJR2PdhnH/C9
oBM/5OyFcaNRLFPQvhF3puw4W7uHgNtfazw/syV4tLkxGk7CwtRW53dUF0EyszQRRiVvE8YHnDwf
3wKLZFfI2TxPHH8/9vO/yi4Sjcbtdb6FDzx6Es1KetY/aiamREJGSjWJhvcQcb1Oej6TKmbeuspQ
FRaTk8oZscuxGzuiYp64ridgGkW+TnpsHC7wy/cUON+dOn0K3loHfgrf8sLTJZrHAwLpxhgXLlY5
UOCy/gzdtKkLXwQOrsRlhssNTY0XvdjQFvqo3f76/cZYf0pQye9Qgj/fXSD+fbmbhyxrycHlkYQS
OlLgamSKYBcUkJ0IcnCgMIs6hKT3j3XOk0szQl6uBxaS4SLtTmITFOXY2ald/s8p/KFmZjJ5suA2
OJBtk19eJ4oF+7ofU8EQJprqcpBXtX6+zsHd6u3AC31q9NRh4f1ZX9TbTAkWzuD64+SdjCuWhZsk
170OjzSd/0tr22Y07w9mIPqjK13UOcPzAkNbOfstLRSYFg3d6qW+DfWLG7/UVELKcy5u8hdQwpA/
9jE+7CiLXpIiXNn+77A0biyzvKQgfIQf5OZapK/rUtN+1+5Ql3f83SvBu7ZJ7aftwfOs7P7hEsQT
eu061Sn/Lm7xvfbjeSIh2zROMep7u0TEoaP66YEJ5RcjjRbndD+grbrd/catr6PhYp8vKcVXkh+t
+udtwaVzm6tyPfTrllIj1mpVxWxr6acuDISvwOUWL/Kgarx/SpX33oIb/JRLjVWklXS+PctwtS7g
N0amQRbCAfFawnTMihG55i4u4dPEA02WeyKCpmO/Q/zSHZf1N89QdtW37WnWmuHCaAiVUmJEO9J4
64oTDYoluifMXmTFhii2Ca60EJePwc7wI6qq6kmLUQXVy/PUtUUeDXuGoNDqkfPoonzMRcndCpDq
VCB0TGYNmi1hT7pmA4xfMnG6foRi+1uK/1rcJ7kHOGLXLzQaYfqpnhqLFH5lcLSfk3COdB1GIIcy
VI8gwaWt4tlQkZZU69aQFIAuvpLBze0OYEeTbSq7p+TI0iwnhzDRVX31aNVMaUaFfZ/2GfkJY8uO
CqQk2SqxqeDbWEyJ1U6jIUS80pXpAwlBkuzShLRH24TESZv2MD9GOULVfoyyEVfTGIzh561tyi0z
VwjJShRR7juxMawB3MThLVx+O+PeMcFGTjTeqTUKuWsIOXtuISDmE+7VPeK+eSeSIf9gM8o7zSIC
YrVB1r4j6GgSa/vtmtxesRqEfhWt+01fhwlCu+Bdy+OOZQ1I3AL7zJ0MPwDazn6O90Y0MV7fIsWx
fSlrB0k8Hej5Ct1mFkXx3siJ3BvSY48tn92ed+fW+FiB7u35HTFRQY9QGGh1FjU2JRl4pvU4lN1R
LMh0/ZU6sYuZrGXmOJBuQ/haCSpBLb3L+tFxQVzBPuYMwUExlBzkz+E6ni6R2H/aPg4g+T74UXd9
qWtYHfjkawP9iTl80Fs4sHm9RJQXshq7gktfuTZROa3dxi30YmSSqNbPwjBlzKn+nrHCTTa+6DiB
2rd0xEKo4jDp6KvQVst0FjtSVEnaUccZn/3adYUKoaBz0Pj4qdnp9ZcdYIg/e8l2j17lFlezi55Q
NH0HLjoYW9RSg5VN3saD8QKdEkZnRtWk5HRRN8RNJ2XJ4iE9bJSymUUmKUiKR13PVX2cHvTZnUr7
R8DREvJPyjljNAXI8AZiJNApd0L16A3GCyt4mw8DwRplwdhEEEKKfywQD/BmOfJFSZZyVbp/UOLP
h5uefGSwRietyhXYyP1Wz6SCdid4jQUNlzl+nI1qxhDHbyaaBezYCw/tqEdFTqywQiILVjfZzTuC
/w1QGa8ItuoXbyveomYEwuVdpKrWt1EnTGFRVUrjUFkn6tMrNgcdlF/LMkkZKFt8ZMZK/urTX5+/
7H1NMUmAmTHwyld2PT0iw4xhJfRvsex77/ot7gXCD9w2b2VuNrLDLtqk7s+5+rcaGZNFcHcjV62I
WH7Oy5q9dEvJmM/BwpyiRQLpRZ0So6uLcVETXlFG4kcWNdPdV9kanSSib72H29Cy8spNKSwrrWik
z37ZweO+hiIl7vSvn7XA+MhtEILsQGfSuxKSXcNVDbNsbAQm3KGmYtW20H7O1Xj+mmeToBflFWwN
+7HYXsSi54DAZNtTQhXL1zFXdVjMrQ0B3V3k/Djl8dOtNYZfPCkTZLkMcadQeYa80BRc9lzIBkSW
R98MQ2fRPEW3qp6RmQMCiBGaYJrtqHM8NAkJPqMT+4J3OKMsg7qwVCKohvZERmO5s1Uo0IFrOyck
52ROCVNPLSiak/mGKbIKmRsiFbezXfrT2EKH5tQYqMo+/Nl/vEA9dkS6OS/7jniBziZINhSBQZMb
IBSb9GOQKh/yiJp2A+DqBWBDnAPRmjAjM57wkF4HtJwlI87CCojsbf4Gn6SLUk7h2ABjI9Ln+HiX
UsZt1pjUZvtmsmuA9l0x/AkavQVxOep5+2lLpILiH4rZi+78jVvX9J5gKVWsnfFLwsZTNfyN8CMj
2AX75GdaZarLwYyKjy3qKAangYomlv3Vn5vVtbMZhD2qujzl9HBdNGg1A7w+EXtzvCKY83OQ6T9e
WeRm/ouyO7+wGkMq7Bgc13wEp5ihjhZS54HJcV0sZIYBcKVrtfyBng+iETyEO39YixYoU49EaO6O
YRju2vESK8vUt/4oUCx2SuvOERX5qQWOYn+dk5l2jUSiHRkRv0YI12xH6ZxWn7XP1t2R//YC9yq5
DyzquoysHD1oq+FYtzMvsWlhbEvJ6wUfNFYmatMe49bGVbskiYJQHw4G4LPdfxf74YEdUBq1YHG1
C47e6yIZcQZIYyUie3I4XLM7RQWzyyHNl7LWYzJaYmmBo7i2jfGldaNdb/DphIj3xbVSBbtXUORQ
27zIPBtOj/17l/ym1QIg46TpgCC2xm4lZeIw088E7COga7KTC4C14qI+UvSf+O+CQ9Sw/BdpySXx
AZI/VvLVLSpmbCQgWIFpPZ5B0WjM5ERFj0AvOPQYhqlL87Pq1G8dSRx0e65VRUrrur0RZQZzMk0Q
djFHla1csFUqBJRkjgo3/0bYhlhq3boHFAcZM8Kx/AlvwsnyFWs77bqegl2UP1Xen0BY4DiVNKxb
tGBHOOk/WyFuo8hEdZP57lQMZc44/kk47PQv/xfVnj10D+doVfGZjLlk4XPxsIiKCbO07LJ1LuO3
2c+ovHhNDqvXzhbKQPhnKZ7KOeo6ZOZFbRChmhEzBVFjEpDUDT1nCjZW3cNwE07UdfWfJUf8rRxI
TilrQ9IUQDffqIEJmdP8D3FHVxvukCtnXg0YMG81MAkFo8UtH5Je217EV0OzJvig9SamJmDkWLy+
5y8wf9k/NiVlGv8ppQzIYaZ5fmD/qS2qYLpU62QI7fm/dH4IQ8wkJTYMV1/bJty4WwAX/BzbEfwJ
JhrIJFERMTGtkT4FCa1O/l+HTOnIah4q/Wj2HfIa8upOx5iohs0tOpLjQYRbDOW/Rn9tDLAZ52+V
msm3f4fF9nzZnZjIU3tsLzk7t4yXz2YLYd8UOUYUsTCRoSyaibOhiLgyfOTsOI9mmtpz2Goz2IsW
MkLuoGAslKt7w/d5R51KFfvZjOpJBsERa31rpyHuUbJjtVUQ3w9gCI46ZYZxqIYzpQY47zI9X6lp
naEQCr0t5ihDnafWUmhLPlQwo1gA6lvHL2ywiQstoNrn6GzjFhOTSnI65Mvl2UKuv1oA5nvgebJY
ydvaz0RakNxHrcDEsMXQVjPoTf2DidYf1ISi9BDYDv/jc3gxWcOLxMP6hF6O1lQ5R3TiWWPqPy0m
7MwzG1UkdanUe28dlQ9VFwXR/C8UCfIvZy+b8s2sfUmnrBta4OddjJo95Y8AeoS4meVNRDq8zX5a
CemMY+SaJFl+717ZZLh6qcDgLzQ8Dt71oCck8CU+lYmG70NdBL7cpEUYTsC0yBDiUe6KNdBiv7Om
5fHLu7n/z3kGic3dHLnjMQ3RqY+kIGJfJCwkGIqO+Ac9KEdDqHiDSptG3ZHECLXlJusF72SVWN7h
gD9PDHxuEm2x+pNOQZdvujDTQWeyEwdRJ/IWfIZVMru0vX2Go+N7gQnZQB0Iqn2ZkhNw9nyNC0uI
QyjAQRgy/la9n40PUpmutIe6Kpw3J22XAO5k7+8sBu9wI/87g30QmZamYcjcRum0EKF6YPW/Gvix
+OV33UJMRrqjBv36s2L97/X8mQ7nXukfjRNKQryGoAhFIYXF0h2ldkRo+xpAbivNkdczrazoC4oS
EwptIqQ7SOfCGBd9gwJv1k0icPH2WDFkv7JP+39NuWPdhReTdJPYfk2SCrBmFI9rcgCPD32mFfr3
fiqvZBpmJZqvJV0tz5uVFaUX5AeU8L+1fXPN6M5ishXicoo0CsGqjDY1+Fua4mBAbSQYlwlFy6ob
TI5mPS7ypNZPk91Mi56MDcXCqq4upiYIhIcXxwGRDdQcCdoDsgT2llaJ1SVvzeK9Lty5SKCwjTDC
GeMTIUGxlphwvfXUlBmUnEOrgKOVAgFH1RzRYrxRvr60zJfqOVjksMQxAKJKlapQYhaC58VeYX01
69Iy4X48WybP30DKKDpV4yjGNG/822MtFZuJ3fu+ePp6nOs0HoTx5hsr0PWbt8qr1vn9jyhn8w2P
fwQp5+inH6ffj+qeOFoPbUKGDmCE/CwiDneiAoDTWzHUuOIsYIRue7mPK0uzAQyAENTYWh1aQNun
RK0t02DEGHzQTdRv+agQf2EbA0hJ3SSB60M7J/WgvzeBgBN378Hjx8FzxhH+b2XE1B7Cwk9lQBj1
QbG77eyZSJzGMouxUA9wb7rWLgUQd+L7YyeEEjZLrC1DLAD8883FBv0zAap/ALFDdogPWRo+Wx44
F93jK5419cD4dIRpYrAiAH59D0/1GTCsflYmswSGQXlvjCw83ktOq0+hQAmT7Ja2hoH3MGOt9yCk
GbbJu0G5LLqgXTwDAeVStQ6XTJNh8NUh0ktDyOxKx1SQZuoJ+Fn/Mb8Cp9HXSQqm3Pl0/PCRr2Oc
dDculvOLh/ZEEQrD+9ZF6qOiRmONCcZj6rjXLzVMq5kYcUqUwhHnzisZl2wshNaQV0F4huMM8WCe
6tFQ8gJtebYMLKwUViIDWGbG9l4vHNXTlC9rN8e4BYpD2FVeQ1ZaNldaCis/a5Rn1t1sYENBv4wa
w84nmHtryvinafzhJZgyxA8DbKSodnj+KQjG40Y5ztUBOQ17WgFYFPeSZYHZ48ACOg+Ol2M01vy4
6H33gn9X8Hw00a2RZZm2f3X1PAroLVuCP9tH4P2d88+/EmUK5wp7nb9SLUT/9IFbhExFQe8NV7/K
WJoA/pYXbSSxTD31aqRxIOhUW5CBYc108K0TJsmWUCBoqWRHXwMuBxvTPmXeeVuUhsvLbgblEZmP
2Wec8/5mb/EnkzPsKfrJdICGWstuxewWHbyvIOOb1o0Nx/DNPxR6tp8RlMoWkqKi1NpUpcpja0X0
LZnHzgjjqeUFA+eOOr4Sy8aPoUbheXmNG0uGjVcPS6pWcO5aNAenbB3ry0ox9Oad83TvsscMkMaH
FWX/mhfrA+YVlijE9GN2KbciLoX7q+jiK49w2dAmAkt8PzTlUCbXUpEFLvzVPGsjwAk4n2yj0u+m
QWbxENKHBbPbjzJXU3Q0hO4gOD+mkL8V36lWthWQIbM0zF0jRwXK8qHSL4LDuicj60j5lzp1TE/t
hHmPoM2qPL5WCByK2MWN5Q7KNc5/Gncr0mk56ONKj/NmnyO8c9lLcTLzK4f1Q5utptoQErclx3zB
RfB9kJT6Ksj36gFLcZXE8PiKOeu3ZWAFLgtEY217JQgwpF/YObt2fX+H0rcSUGTyZ6HEZWzm6toa
HA8mZWgEbaBd/wdcJH2/5RDyB80psOwoW6WKQ3VOaqdVGJ+yUxhb8pZv28ZLI2TadpUdDTV+J9DX
34seITb7EQkveiHFjRuwIBgyLubk1+rBbjOCwzWS8VdnspvLIbJOLsAKR6BS2wVa9e5fYDTUA+Kl
uzOtl53zpZtTPfzXSfMAh+Mfg+fSVRcZWnZ7BnXDJnKmlRVxfEME5nJhZNgtfRyw+RwHSU36sRil
aZC6tT2oUfrZqexN5vgklmjNnfnUV0gpWtD+pK8RkYErwMQPdBzoYk3O/qb6y/8PBxN890y5bkrd
1SKIpYNiNA9IUEZ3+xajZpdxGQgVIq0nwEzr0RIE7+wDSY0zkO5ezZojLBePGXwgAM5cXA8SMoH0
EVA2W+pR8e75I0/AzS8y3MsbH0XnzFBEYC4jAK60FqWLwBwA+8SC+Uj/JRDKaGn8qgyjPc80ynt7
aNH43bOYizLSb0Hd+IwlfzbwOpZiBJzQtMOAMpgJlGy4iY10Qr9ggLXokSaASjsSlp8t2JaKmDfQ
euWD+I2V2Qj+Qazgsj89ctL8JN+aHmlMsHqYgFNBVns3R3A6k3BfS/kHVEM7osOu1vsbETiAxT+r
LLXuFrwAlXPvEFM9A37vnz9eeNG7Lw5ePMkSBQpEsaH10GvjGHrYqrKrAJ15dS6fGa9Vboib3BmN
TjbKdrZff+qfcz+o0CcpB9HZwigmTZCYrOZErVgm6S139fGQdh+d0LLUOqyEYTaCPeUWcBu7mNl6
d5tPaUYsDGEaPyfrsfyboicJ7Kg+8+qi7DhD/m4p3hoY1I3MCjbvLMuYUWT32MRdThFAeuXHiqHg
MHEUFHwif1Cbkn+FjUQKl4QwLB1zyjRprIZHdV0T+Ds9/ci9vRjqypV1mP55UOn+7Xi7iYqAkdfn
46orI8DjbEw9JkwtCUIbDDyfmEhtcQamOR7CxDiI1jV7CT3/Vx2VSeBY+KTm4wLhpLhS+ONGYF0Q
MoOBNn9Z1mhVv7WKrQqNRJGJsukIaQkIFcHI2ZF2oTmuoDCJ4kxA4oPPjceKa5ijfeoYD+ZN2AkZ
c1EX4+JuSvc4tPB8FQQ4VV63rsSR6u52Q0bDmUMiiEUEP9vhw99SSa4C+gIQN6YRZviCZSkrsZRg
ozuVEBhlpGA/0fu51HZaCN+EQ5pEp05Xnj4SKjPcvvdL0l834H4c2YWb+uiXinO5NamfvFLF8ffY
AkE0tqNTP25ug3SO9VShFSLOe3l0PAqo+omGF+Qvo6HPEfeMkRHnp/r9Y6K1BA7F1aREfsVwVPt2
pV6lth7jUBUfg2urSF+Hv0JGoCzsflCKZ0f+mkUXmleB9ukvBjV0YkY52Pr0KXrp6+9kBeaqhHVr
e8xkrDLuUl1F9RUD3SsLFnoez4HIZML36WQZpenFS0ep1AChfmc8RLL54a4bHQr2XObHIUAzGGjS
IdD2e7HA0WC3Fx+YwrkwV3DOH7+O6VR7BcYziTEZJCWsyw7k+3Vlv8OXUnZ1KHOGHGA//XWv76pD
Blse52x8ER9nznFQaM4TUyPGtz5aRRRfHeHaSpvz9962Z4jNeYNF87QPtrepIGp+Rv5gHOyTEEO7
dZPHWQb/NEl5HxXftLGkLpd9Z+yCerPAI1MAnbFHBzmsq99hAZAXEoWpOVSi+cq1JeNkVh96DnpD
yNVaRJ26SlTN9BWkY1F/VIO9qO0tXGndJT/jbCAPRGPGGwO8tMlTQJD98v0J7zZzqRGx48aAvYTD
ZHr4MDG2H5UfCJm3sgaHL6pYYzpXQfqoUodkdFpR5zYFgcfJqgdz1mJwefq6KVb3iYDFh1vbd8Kr
Th4ka2D6LdiPnn8MLP0VA8Ypc8cgI6baJRmSZC9TtLnshqunwwYrKJ/jYr5z3H3FIGtCnKhUbkoM
kwJwN1yZCsqmI/z3S1Od5DnrDhF+9PfeWpBfipWPSrFPa5GcqHzb7dPW2TYUnxrcMFRdZ3cpGDNy
ZW3Xphk375wcv4BNUHlkGJ8aJnMWxxQLeQOXWGYwQQoVUpQOysVE81s3rVZXOXvzE+Lk3nqiOQuB
1kwZr8oHkLTaWdswqp9HWZOEFjB9frm3geE1zdey1fz80GOFT4BqPny807LZ4OBpGhNylmWuInn2
2BvHGyFEhmFaDV++Spd1iZA6hP0v20K2nigp68crwwTJPrCZRYBFpnlW1yddXLI7qwfmmWLEyT70
CfU/Zm8WdZGDn6dWmBi6F9aesWFErp8hB311SmNMORcjME7RRyl7NsVXGUgO7POfGrcqnL1RhpmW
nXIdfJPIbEtAW4x1PrbxYBcxflGDLdQrOrwvlKaaXORznZeAXsVF1ITb8QCaTc9NQH/4mTzkpPzI
YfvbCLu6/10b9JDr7BEN6nCgGyrHjOcBAFBllkuvXJMg+dueJ/Hs7OT/nbV61IxZWVPqsWn3Au/c
MRGkIBO8GsQHYSG7Ddyhasexgt/p/9aOQxs0t7fogSHIkeyWP48x7tmkHQw+ykm3fI8x561j0DrX
d4GczrZEu8n7YutbGshbMar+Lpo9x9+85yZdIgvI+ovsr+CCaglU+diYgletcMNMz9x31xA1HG4M
68dUYjwkgihh9FBb4fV9swUDIF0By/a2iip/LXy1O5qkRJ9Onok0C6nMR1Fhkk3xxgNNvhNhE+Vl
ykYNGMOczMCjQgvHY/0DYjru/NbPoWHWu5E2Vu4zG3LR2Dbs8tEAo2Dap5kwX4AeRsrhm3N04msZ
uLVIYMC2F+rs4/85Cq2Hr38YGCUHA6IheWSRGaJncvcQhLrjUUNWKGtNwa2u83Xn4fPibbEPuq8H
7POyxugKy+/winpmortnhImykmby7IjoquvtLLaoQG43n4ejkSv8Gv7NSu2CP12tDkY8ERVVnVCJ
3y5cp081OtLCtD6S0UGtYsNrClcaQeIlaje/Tcd/ud2/htL4fs82GSZuNfYvDxzXigfhGdNE8wh0
OEusQ1Bfx6JqAAa8KWHDeQoaIpd1fGmqLPPRWiXV7QWXzTdpmSrUshS3VpKzK+I0fBZuVmH8eAkK
kHcbJQnaPTiRLd7UUdfZQlaXKAGmLYqOU7Wh1UYPTCIZoB4L7yWEvT06zg4sM9UNBAJw4hSx0kGL
QLn5/3iWNgpzMtKkkTfm4GAyTg/LinYvUDIJl7JyFgPc5kO0P2SvCFYoVlQyIxDLE6AJpF1rUr43
TTL4J8mV+gkGsVjRgi6LwMJLuEbLGADn0r/63Gbv3vIKvMKI+qS9rfpM0Kz36GCnVilonrlajYFg
tNX7S/ZLXjvUvjDK8IxtG7WZNY7NMUjKw13rHAahU5xF18oBjx9TwjcVF935jxT6N0jxP/CfiO5s
fC62Khaub0njKfSiKYwFYcBVnyEu6fLRsfrGFSVKOHxfNIvjav3b58tsM9DPqadwVURrMcxNXuS7
19HDR0sggg4O5AHczxx4MFp6RIpSw07xTIijzVkG8cCtACwB/kAdq0vQxiNS6gbp7NHj0wSXBbwn
XKW4Sres8+LXaW1jW+G/goZq3cGLK/x5Iul501SiaKdQbMaZ3bE4NVqVlt4ZO4ByQLeCP8JfzjXg
Juj5pz4V3ouNn+sJG0VuwQa2E+MN/LLqlJL1Mv2GrOIryjsDYkt+atFm3TzzR4oyKwjhMpwsCjQn
8QihTh030eiu6+eixky/ai8QGYItw3XRoYqco03SZxJ2umAxyHO7CgV8nWcjWdoLpn5rQNp+BEJC
V4vpRU+QEnMJSQnUNPuuMn80r2pUx6lNzrpxC23n4Iwbe+gi83AinlSt+afifTr4egD3BU0Fj4h+
FVzdyggGd6hTq64cjHQ6BTFasbveuCF3aHEM09WOTHXaiqyt4yEDrOytraLANM2eYox0XrEsw7/y
qojQ/llTVh1+6TAXb/FWRRsSsa0mPmwa+4XG9sG1pv6w2giD/kgdRcx07UH+RYDmUPzT/USl3ozO
2mdR2eXAeK1a/AMqxTFk2Zw8zgPn2dHAmmxtd+TOT8jLUu3acrpdYRbm3STX18KrJqDoGZQjsMpC
lYxBau/liMEw7G4bSgCH0wZRTNL1RqtRqWg0gVaUKe1y2MK09NPEbRgIXrr+jSZWiKQfnwaqtpAL
lc4aKVCksVMjLxw7pR2z5JedcPe+1sFbHDcOTjc/zE26xEeliQe1tn71nLJx5fFR3oWbGV5MoUzp
PvRyv8oUjPwMW6svKDaX3FWI/qbiO2Nc+Gpx9eYZjKhlCJ7+AOpko8RDrOa82ibl2LD6iuwnSolP
QsFMXpYESpteMzVv0vQi9aDclHqm83PeFl50lBpEubuZd/JanRejLHlGVcEMH45Ro1BlHx1Aay0r
H6Yix+rErpK1uJ/v/6BiODzpIB0qlfne4yG73gg9VeR9P/KuTZIar0jZB7knyPwi0dctKByzhuI1
r35P4dOfzsRHqzS+jZIbT37iRB6VW2qN8jqFB6CinOGiMI1UjJx72rTu06LM/856pyhiomumdA3J
EeX6rNyd4vYP5jlckDlom/M4XEQTI9yqpTHQCk71aNGVi2k8Xuog1r80sjRrjaNEiJejkH4NnV4d
IksGU4Jx9T80Oxlr+oUaW1hBehfHV1K0hKLaZUMeO+RVxUB6NS3KtP1g9FPeoQ8MRniL2MTkmAyT
ZkN0utNdmBEmh3j9N4HevFVYP3K0JpsbSEObRLU/4We6bZFxipIt88O9V1nB0Z00xFHJuDfpImJg
S68uRJ6wAeXXRLToY2nUiu9qDpGH2yUMrQ0xTk+HMB4hX6RD2hYGKwdf5oq6R/uA46rpXJN9Nwko
/QsOHXSPBii17K1xED955xuonj7ACtyGBsMu/YnkxS/gY7jy5ZRDCzQTkKhsV/jMey/+Qi9lrYZz
SLQQ1snFzc3J1rk3cfrX118ix66PPl2eoTz7RM+UiA2OZivNN+Vr65nZjy/QXNM+B3+14BJL4R4W
sY6tMlb6xWMdlAtSDwdfY6VnMWmF81E6857qZMgc2V+vqd01O7JkAvYbjvmS9ke7iNrKdl1drQJu
7udXlf4Ys01YDDLeVyIiru9wrB6vhio5J1/65pk2ZrEAC6N3BmuZArkTaCWBFOWhkZPGGlayYu2a
bisLb8WwLXwSC0hD2S4+/iDRbvNz2TnwHTsHVra1WgI1R1iD6W4qjlh4Gm4vuCJQbx2cvp6s9C3c
8BXd2btkeLsUhrETPn1CDzL2t9U+x9FAUKSIWjSLOZeVtmn26vY5Lz50iwlVIuYU+JQ98863efOw
3i/dDpMRMF5GjywlOnM6ePzj3oB+rskqjv+bH+mjW7qQknecPfSSpneHo9ejXfOtP1FESvxIhRbv
2/5lV9+RIrLFx/oTbIG7zE8uNdOc6wirEBOURWOJMnosqs9NBbYmQ6I8HJkeob10DecA09TXCK7G
lTH/U8gsIufpIK0C0Z3YDW8ejEwbQO4tbYWmF6D8Tbr8gZ6GcNg68ddJtNYLJyEPnIcXkEJsmVAF
Jv+F/zE4nQgeAwwpCcpHei4ZX+Dw7NpTqcohEl3aZgltjj1BWoW1FzopY5YfanKDyIhT5BQ+h4wX
kwOblvBeZexQR1C+90cCaHEnd9B6DHl4FrkFAPdiGoGTtsUYBEi8Wc8/mQq84b7+NxQ/rPSSnrAe
d6eIXRj5WPpSVCq/OKeEtD7hToslrdp1k/pnml27P7twHIR8EpYBrTCIJERpIwPhxLbz0ePCa9Oa
Nx6Xv1FUCFjIOZyBAPx7l57kdwrD/dErgot4eMASxn18KoceVCMbdZWTl7O6qdD5wQUi9ke2AINl
+6ae3lKn04na9vFn8zaBodM6AX5Viz9G5E967TPUxJ3C2B+z5T5ldO0m14l1c7rBpyIdDh3jWApI
xKPvQdMQntA/nzXPVw35hSXMkQ3KOZNDsJwCgJcXcsRBoqePB/5rTSiepMa1nZniuaffXyEsOVpc
wqXiQ9Qpp7qzDwoLf6Vdycc0lpCoTx7+7VR6p0j/VbXpY8/cMVmHX/c9Rw5ohpJxLnL3QJu4KU42
T/MI8ftapRLTlnufurl4L9g+kYslsf/0fWkE9zay2FDU2q0dyIerBHWuCPlPsKw+Izl8ZsUsJIOP
8SMLBBTM7RmXDQekSYv59PaQQ5Jp4F4VgyNdC4VKtJw+iwCZ91lcUsJ2jrdUWzegSyGU30LEBRl1
XxU5Tta0Yin/4g6Y2UMdc6oP3ouAqcG1pFkFBO7UTXIgB0u33M1lGMMw/IyDV3kb1HeEVKmFFcAk
03SxSjcSLHyU9TRQe8uxY8m2kVmNXdSICrnWE31UNv5WyE73Ih83qT+7D5JjYNOvn+cmzp3Za0A0
0EqKbwooMOmv5RTz16mP1/Vf/QBDWKX03i3i/dbiBfHngQwDhjrPdcO+xf4T1KhPDDbZp9M3hpc5
ffNPkjR1zzGtBJwuZQ05ePatBsKvY01aeCQva+UBTv6qf6SRgaqcR+QqPOcCspdjgpeEHy/A3BKV
C2D2IYVpTJ5Xl9cacDJh8qFJjBNi3TI+JUC8Z8mhuN463i0VfSSztQ14xDv0ppIqAm0fvr71pBKx
AKtmkURfs0Kc9s/9rFQVO3hVrerBUtxJIfUeni3U8jMhfMY65mUdXNoutt1ky6aDrYIJCrfEXBYR
jVc/fCIdWpEaRO4Om7Kxp98KGYEm3us70sAdAWaHqa+TFBP7A+ncHOo8ro7JkrrnDT2N9ILsaob5
KMUykc64LixrFjQE6D3ujIeu3hO8SYatPS0dRVoYR4FYci1S3MqvzqoGKT4aBpzuXkEFWiz1cMgR
z+o++t3bpZF/GlKX8SdxaGHxf/z1S4kkdnMJTIWBE/c1zyC4dI/Nm/Dxu1qgCGZXyOinGJ/vrSeA
ZRx+HDqpI6QI0BGapqPsRRdb6iC25e8PDLWF18whztVMjvsdqXZGA0JlhZVhMOWWYshrA/SiCEqz
KVNd4/V8IP5CsVgLV9mKetqkBq56lc4dZ8frLalSkoIcBnNnt5XRl0/c4h4E7wMRflqT76KT+zl7
WyDS2b1pm9kzSq6WwUKOoz4Dy482JIf4Wj3UsF3HKVOhctU36NIOHlWQQlJNU9oqF/ZhCPM710GR
oEsoDzdWiFurmdPy0rZw9Dk40VSIZQUjl9oJJL0OyIPcLa7i0dtpK59XrY4x00klc6vSNq3SMydJ
I530ILJ8FEe0grLf9suigHiOB/zgvpvhLnXLkFqSSowa7i3npvEluZnW7RhsbFATzNGXCI2QLkmn
+lBmE+fWwK6TGVRwLQ1vrTqPUTdXcBMJ4FJnmx+6quNs/PLgClZq9zW71GgTmDF3bgf+KmpDNehW
MMa9+P5dQRafonJJ14ebHoj2WN9vo+rguSf9aVALI9lt8fkjCpTsJ0i0xTYC3RBKcAgzcQ9SLJEn
v/2OuNB7FLseNYH/4hnImm5CMeVfR+Xsc18SQUUa9pdD2T6DCpVPuUxJyiZJDaoQCmm4VqWWH2kS
1LyogGkI5frmtWUfQ3ZS2lMCaiz7o1BvIp4aSvt6/MbJWB4PAFIywMO/OC0RuAtfd/KV5VijtOTU
oIkyZLywfo0v+wbDyaQLOWN8/86kpplfo4EygGevI+gtOrQJaBJWPcoo5DPyeTPqXELWvF/yJwo9
8RtdvX4NFqTUkIqPaUJZK0LwfqeYAbimgT0Ao36lESrITJkvgPk2KkGBq2AY3GEgoJjsx6z2jdZi
Vq+I+9JMaBdZG6duMmF0xXGzAVtCO+JwwTVWN6WWXmsADyNSNqiFtP1+fCPLQ8v5wQ1QUTq87crx
wlqYjJQRa7I/xtSKCgby0Vfdd4rtdwKwfisw/HG9R31XW964LY9i/Gb6BvBJwu3YFbMtA04OgZEe
Qi6shCHhXFu6C56yk3Ity1+gOkJdfZ1tvNA1H7tPv/STcbWlYrqDXc4I+T2Y8c1GMtAU9m34JJbX
eEuBeZO9WfePsEPngB1OB3leJO4bo+X1Qn68Lxh+6ia0QDmkfOJfSrtAkSZCyk5fqWJvKk+fUJmJ
ytudr5HlJbyJExdO9an5VBwZi003mbZKGMiseicrW8ouiXqcE0trSCwmlO6OFTkcXNul5QGeixl2
kGPfTU8dqRAlNEbFJJpT7DRV+oSac2v0R17khjgq5XCMF/sewujHNEl0tE49DIHV34pTwfGkhyVF
rw2mBJXpl3TtbpM5npqMgp9qYuDhAxPZpIG+wzMtWHyDOTrUJUhX4Eu8Tk0Cd6Nj21kE9S+91ev1
EwvRdWxHuDvzo4lp+bBass/JwN6dTDDEPHx8csQFWayXeSGFyX0ekwTxB45pJf1uR3kYpk8zHF7w
AHz8uU5s/1D1yZqNuRR3PzRpu1vdk8KJ3ilQxmsPWR6kty39ZPioliT2n48x4oplXA4NG8yA0YD5
fevTiV/mGuGcSrxgFyyirHtxjSHkV+lEIOFGSMZRrPNbwPhv8aGrdPgy/NBWGgW3xeGHGdwvLtQw
Iz2JHZu6Cn8ZinfEq739lSfJs8vKlvFoqSXM6EBBkjkLBPgpfpFl7HXcMTEzfLEEivmiFoqw1tq7
Xo/OPkITXl5RCvNdk+T5mkmRxr3ujrEUwVsxm8I+Zgy2GYHwQuapXh8wLw4j0y44nWvehi8nyCq/
cEnn5zLJ8sVRAyYX36VRdXoBmq1Dg6bbs1bOql//si2MQOInRvOJMQyNyfKD0VUnrOLhA3u818Y3
45wxtMp3NiM/Jf3uVG8EJdbNPSXMeFd+ILMNgTM3/UCgj2FJYV4S2BxzOmQUTGwdTY65zRtolq5G
CAWtzpq9racEN7W+aY6cyFC+pgVfkuvaIDJPhU0+MvckLC6pg9p09req57luaVivEdGiQRKd8yWa
jsDqAYPWLNZ5k6Loft1CiotjaF955CD+5AZ7nbpFRZT/rzJtCFcS2tRrP2EE71q4fGoMUY8h1Dfz
1bmPZCidsBW1fKrugRwNZl9mh+Li/CScWXSyHCxDfrLUdujk6kmLS41nLEcBBMd++32IzM+08Aku
cZLsydn13aP7LElrV78P1N4lQ8fvUmFY4Z52EypQHCnEwWAJg0CA0gq0NQvbp7Quq84JtpX5xrCo
4oTwZwCqFNPGSdBHNAGm89cKzm0cvXsQ5vx3e3mySC1Xrl9iuLf4RjBhJBmbmvtDFelI12seuKbm
obMeKcWTLCuSQOvpdQJOsKj0hF/TgWrXSp0binZLQIugFl6q4LDxTp1lVG93pRhx1bqPvU/GQ6Jr
bnGoS82AQutkbQPX5qd+5gR8u14InD8M6JEhKQVYf0bgH/EJyfbiJ8i7PANBWHEEXobRzM496sPO
q76pVSu3PQW94YMol8s9QXAKuyaR3nYJW+k8s7u2h86QLJTER+aZhrAtxft1nZnUEkz/a7p4HeYE
HrdPlpSI3PV6qXiaC9kkAtNo2q1DpsoqtSIyORTUJMnQsyvdEOnczao5vSiWL6Kk+/Nx88eNWNgA
LOxwgDjW2WpmolllgTQmFWjHea+zP4JM80lxXMM82su2nk6H1qwJr/BlBAyjNFddGPsvyej2RocY
CEhjRXrtrUsVuPWeurohtz0RIBIH3aH4wqgMucXb2u2Y1IVwVpmrBN2e3GViSLDbsLjQb8ldKIWV
lKSpD/QmLdd5cNy+Nvucfxdile4LNOx+rE0Q/X7FXf/R/PvmwMnNT1xh75i4mZMDPF8F7QeHIfbr
wMo6B/9Ijsxc92eNcOs+7leoi690nEOO/B/aayMX3/FBvLxqifAfdHQ1/ZcGTxsIMs3JAtTtY6E8
XbjJxFoNAlSfh4m3tq5IVHE/J4aa4i7oyQD5NeloeRhJpXheExs0Pf5X8BdIY6PqoaKkMBOwx3Bf
8fTF0NTLu8GOW+venp9ouoX0nDRdql/dDnGWYflat4Zlr/1L3CflhyH1glWvNjq84RGvMo/gn9o/
oLf3GeIjlL+0YJvNepW+wFTtaWURi5X7BlCIfd9nI6R7kb5wfnGJ3LhOyyGyBd1cADlVhZaFISvP
XZ1TdQJgnBtTq89JIGwOakhI6NjOvB2agOv1TXMMxAzWh6gJFMQrOM2eUqZvlRYD7EebGcAnBn3K
qZo/+YYFaLZAjjBVJ07+CxH5SVhtxTh2dDJjVaDrgSed8J85vTNnnykHB4dF7mBjM6uA2fnEpPyQ
vpor5k8g/qtkOXxOSVl9K9wBJsUxnylfgcRlCE8kMcaweY1fmVeOrOtYMrgsccML+NC2cU0XB9/v
wLVG2cfLiKf1yWaxgqk7JkWve5lMhWjntUzZHe5BgHT49sj2/nvZUW8utdXMQJD3H+Z8CmvYPVws
ETdVICPz5h7ydmANQmaDhJHHPyRQTUB35/GMgNV2dh4nCbx4TP/UG6NeiZdxUMCqdCR0XeWw1v6E
7XX6Hodj89Tl63Dx8rzlvdc1CPK5gUpRxaSDZSqzWBh0QICAvsevJLSciDBctJlpxrMLAtTc1H8k
82LG60Mzhuumtp7QuHP5hzIK+uTzD0NLfmg9hZ1/8GmkTCzFQU6hA15U/gpiCz45AKGRWh2guAiP
kPFnsFG8sgsRBVn2WuB4647cIhddVfOH8uhkdptYN9W1XHeTdHXGAg4Sw5ShU6VGSQvq2tnQwOuU
NgzXEFDWyiiFFQ/ZavU4p1SwicSAdCJ+zJ8bps+9Fy3Iyg6ECukobBeXMMGn6L99NNzuvNkuinAH
8ABTtT4WgojfOc37G+Pgiw0QchwyUQNSciZSs+wj9CMcNgNHd5ZVxkNqzUnvaW0ahEb0OpxBkBon
rLM/VJd9FQroA1ZvEvmwsUJb3CgjYgK0OXdFb7zvSCO7KG+g8nE07B8jSBmCjmIWCksxEaPE1OTK
Jk5/o38Y6rKtprAK7DuSUyhj622gSAwMsfhTqleqCY8MuPGdC9Uy5cfhhUdHKw70aHCyKZGkFfIS
lK+xJ19TXsSpmoWfGxODhCSM9HJSk+LpBkYaIsx8PsLUnaztaWR19jvzN/UfaG4Jd0bxxz9I+BP1
XHAcezu6lp6qa4vYvAfGsGTzEKdFBg0pzCRH4SeMKtP7bXjmp0iat6QgqEyc5c/seMvk3LwWNb29
qRjYCk2ecwgDJVQOQpHK+kPneIMrkONhj5z6muBmJf2mlFMynjJmR2PKx3a/1nBDDscVtF3DTQVT
pyBv8n5fg87XivCBwTAT1QgvvI16BVJae0sJqkg4v4MYjO1tpJ6KnIPo+jNIQLFqRJOGBPM4Khzk
VXul7WKIHr1FjZa3u/EY3840rr1AJozsp9dbJTxK7l9Tl8Ah7dQY+gWaY+VM89/wZqQY/Dj3rySA
XD8OQqBznDy4M6l+C6zmGo3vMx6k0d4bre/WvQPXqpvq/iuYcrDNGZgNWqpL1YHlXbxJM+HHFa2B
TOqm8hjUpapXElaPL1IvN8HALNRcNAzqgt49oXEfC53DzCWh3wTtzVruNQle1k8xPsLlvvHTP8Xy
udILvbeyy8ifCGg3zVgWfaaqQoDhyesH6F+66L4/0lS2/UJM4szfg47Cqfx7YKjmW3fFGbu0aBzY
XV8+0XoX3os33V93k/H1hk8/MFBp7UKoIIIeEEZMgAAvdAhaVRLIkpf0nK0lcj14oUzdYtx0VDZF
wHDyWn4Vp3aHFLEJaaCkA/RXsOt6cdz6aqk1MgN0Prku4lPLxaC00n509Z2k5tjfg4JEJ//8vXvn
0+DrDauaB4CpHqNl316s1rUEHepmrZJp4AJkIiXFks4mZe+HiR1/qMjgNxPxkzmcT8i92P64iSyx
yv1m7Tvq0th4J+F9PaICHsuGllpwEx1oVvTnC9oXaj9cYP7ALO0w/aIPJTHoFgNfxn1SM2MVKlLy
goEUDKQWsXrTpXFiZloIwfU0wd6WslE1k50tjJm9jkmskPkgMJC4yQgPdMFeHVu6/RY2G9kjmDR3
M7L9SZa/9W8YMi7AY7Sny2bodDKXw9dnKWnbwIhpTGg2lN+H2yEM9XvbECDl0re32XG4VZ0Kq+y+
L7+mNNsVJ/rcyar+PmOsUNGytdUd5woWkBFhGnOdxpaDp7fYlwstpVOLUXBvYqserXXghDkuD5gv
4WP72VGWI4npjpODNsZbJbOAKZB2QskPPdszsIWfCJ21zPtdj1i0xHzBZ5gHMz15Zon3X/zTfAsP
+0tUCo9OEIL2eGevckVoxkEerjqA33Eh5bix5oLru6u0/5DOlvZbywgC/ZdHLFvlG6W12uyVxPjX
XIuMCe9lWV2NRnPEYDo4FOOwJNmbPhJKeqTlIg4IZBBUwRG/NUaCRIJgjTu9xbL9uH2QE1ykudFA
mJjKjcuzR2B2PWqsQpLJbVCARDXgae4h7Z9ple9NMN4MKV4sddP/rDbPM2DBPpMQHDzXpLOhRFUD
6lRoXadw41g48q86CEwv456Hq6FkEVlheN0vFv9D8cQuU/qCUIr7ZkimanWNDk/DKNKLjJE05m26
BmJnH6m/1RcO3TLmZJcPXjT4iSe+vyrMxccglkJszSodgsWU4NTiI2VAC5V7TCnCLhr2VzImvFKO
JYomqVKd5y3knUJksk5yI3/j1u/tTtbQVnTDYWrqjEQm6hu5vvX07gzhvlrUBy9k+75OElrfP8Sw
PI+YEtu19zCs03xeZ+Oe3mxpNyB1mJOq1A8LA/V1d9zxAqKKaOFYwoppeObsw1vpwPCDj7TBfSrF
aa//p9ONz1axWJJ3safseLDgsB6KKjVCuOsTeyA0UZmkPLyUtdTZdwqzuD9q28gfaBQgEF/QQkgg
G/QMPdqNwzHsNrQCKBgohjWOaObpHjmZStxCPd28CZrHk7NO2wx+7lOWUXzoYjo/8Dp9NKkJY9od
wPhmju7irGPNUO1WBZ8uStE0NCPqdKDvWo1Do2h8ExC09hKFw5CkNSnLV7cQHz56EdlNRk1u6B0R
GPHDY1NDYxcd2uxxbn2ALAnTUThhR4+k0VJxl05URWeQzHZ8diujwtLRi+ZISP3bx+bqUCpsY42J
WKacJ/Uy0wLGGC+mtSyq9DK9K0xqu2NNsjD3XfJnQg5ukGEvwJJkNKcXbd6DCmdqShALKZ/1n16N
3dd599g+j57x1wwS9uqDeOZU1KkTPTBfIsUZnATXgkMWYQmrqRnJNGeumuIFfmVa6UvKhfd0+5yy
BDllVFt0kiG2IKWesoYAVcX3ZYZKaNOxzJjc74PNzhgJaiMz0WRKdTHr4o/5bqOQ6WOTyIV+UdRC
UCSj6htPDV/k3IFVFfdN189wnkyH9MkEQdKgI3ngmgG2P/7qVMIFzJnrOIjm8GTcZwGVx+Betnrx
as3f7uzhNJcrlXNGhzmx8K/svKxjvRdvayVu1EiunsCl/mkEgxx9pXrd8nPjaWQdBqiyRk8qfH2f
8K4TKGqCUeHdRizHdArxx5+tRl4hWA1wQQEH4kPzmEaG8GUvE9z4la83iKZQs8MUBWLih+rXKLVR
CMMuicpdZCSsh3Dd2w4JAlDCDG/wrvs39SDt3Iw4zOZ0C+0TPj4SjzOTTx3KkLgudG+Vcc7MX4Xc
IHGGsFrbF8tcK1Vo8CoO65ZOduTSbkIsYETjbzH+Rmhv54kISg+Nc8o3iM4ciIoNCkAqq08Ja1x6
/KM+qeT/UePaC+vX3AdL9QuL5+dNerQS+KJaezqOV34q7bBzCInZuNpvkHOQIfsMoq+jaAQugvw2
bJf68awZgkUXJfK4B76C7ineu3oHOq3u3yqezLvvUyNCnR7HGklc3eztmdDEL4GzQDMyiN0YCa+2
GYCzn5T124BegXv1cX6hmk9IupSBgNXFH2UAo73wTTiksgfIjhXrIbX8Tr/dB0knBXiwM8GLHZYn
JIjk8o53Wkfs/RLyQWv0Xq572Qn/xtKqAEbVVKVikbfMRTJhP01MY5oRkJurcUk9SN7RGFqPdErX
KsA1Jq7K7dzrGQ8PnP8qefrV2XU/8Vn4B1Mv4X0jwtUy1y738eVfi1J+UFM+2jf9F9uDeN6mVgW+
XqaXzC8ucFa9jZOY/tgPsR+PfhNC3EgD62Ku9+BbHbSNWjHRs6jB7IOM6DoVVVEwQ4W+xcJCew8E
7ZVUj4iwiJQZZHDORjKTEQgUH5CbBIL20pZpMnggRgeRbJLIfbp0iOoqsROjbbrNVwji573koH6T
MUAAHDxxZDDu1wbBlmtG1+n+1vP5Yrp7GdjCFgDcumaovG6nYeKJ1Lr3rmtZ/V5ZrtbSIesOfC7S
qGdfdzDt18QJkVLOLgMqUPOvbpsx/hmC1UubRq6xOA85/D1i4NJk0VEh3/PruZsMYrlz6TdVrgXl
oyagoqxGFp1/+WOI/jgF+s6RC+6RvD2zJkCSpUPjKInVf4ItFCJL1xoCLK9rcmrGger7vVendSyo
qnV6rR6DzTRnKYL9dgaCnz9AI0lb23pUf0K/VfZs/+REwYHtisXlxwfVqYqry0cqVDRc5FPWvZut
oWW7Ln4NgiwXK8KCnEtJgj21TfAG5FEFD1ey3MFl9k/fGER197lUV5muegxCHkif8Z/TpDPBX4Si
8munynTtYYs+03JqaoQWXPXbfsTRPHb/ZlyqUZQ/cr3KW/3DJ5/O1P/vOFz+O/jO2OApcvfB5Ptm
VlBTpj/WSpLdFWsPvfIdjA3tm9ctfgWglm5lGEpYO8HCrPhnW4YUNE4pQxEj3ZUuNbMKDRg92nU7
wMxHEMGUpgax80tvxOlp7/6RooD63PtjBxt+d8YQW8Blfv6KuQqaVxA4I2EZMqGca9nQtX74lpSv
zzZmZ5GCLAlFfQTETiJLAB3GI7t5Vq6mfKdNIPPmkjL0XDRHZn02d9eIZG43KCydG1tnMP+0vqQZ
FavD4yNZ4X11J7D+7RV8E1XWsJ211PKUZMO5sBQDtCac/CcRyojabtZyJToTQyJhfJ9q+XA0I2Tn
C2RTFPn/g1TbQCAJe2dfqjLK2eQQCloPG98/ybfPpyuu/MxRXue31eoT52sAvQPcdh3vyb6DbNwL
Y4iUNA8WlUutDlTNURT7jz2SeLHyyJTSHLQt15S9YqLla282fek6ETvtUehOLWEhbMjzqFzE/luz
ZdojuuUxbYnLtj8a9Kbd6Om+ULJeluId+Rezqeae7Vk+vkjQZmSDcOBQr6+/bkNO9D3z5Rbkq1jH
yRr382daktHLcO/witd1KRgyfQ9K/2nFwTIkiD/m9bNsXB5LnisnUpFOV3UWMTnhsyWzGvWE6h20
dKIwJnBeAC2dU0Eh9zkUTI3RKXDxtn9ZOdZOnjHP/VxcXR6wtGS3eZEjDnKp6/jTbvNC8MGrG6mq
vjWFmEaWNRBeFNwJA0/a1iE9g3q9wQprqQ0ioNGgVKdWzbcC9JnbKyFct3lScu5ILCV0y/kyoeK3
1wc047L1+ryJzVR0VIpK2L9PaP2im5lsjwKK/uT/3DS9XsJ2KKV7ASEVFjcqIyvNEKqpiOXybrhn
7zpDiSnsmQgVTdN0dFUtCavXAwV3mG1ahXu6d5/TaY/95Izytt8Lp2nogAZ5oFEn4npK6wzHMytX
xkm0OASMOptqcVNQokYERB6vXS/h7+PUkkkgIdpjq0MoxrBxIm+xgJ/49PXj94YtWd2/yJEjzG/2
uHPte0Odu3VoN33wvxUEtcndl2g6ZMC+hJ7pauiMVRUNAD1pTsMd2/klwT7tGYqxB9NqK3rPnL3a
h9s4kQTwpPo43iaPJx9FisuuLshp9BD5UhV7mFJhfIt9lZx3dcspcY8lUU8CuaFvg/HN8XcIDwdl
pURXXrx6SdenDXHsQB04zv0+tJRLb3IdL24cFjfscY996XrPOfpB18e6uPx3udgu/wl+OOiDjZyi
Oyynu3D6J5NWE6fiTBEhK3T33YbhTOhXDzxzkjhwZ+OC+08Gc/7UMhqTgvY7bfx7z2k3bm0idvYe
jPXp29MsyHEaChmN0I7AMHGoBkk1ugZ6cKLlxFpQ3CWqM/YmhQGaLsUpMhkIfGC37B/zVP5QEUqv
yMBKlXBWHdu/OCAp3wjo/eUh4wS7TTBBTiyyg0vAOSjL5Qb99BAPcZOtj5SYdZ4Ib8uf0PSI1uoN
QOUl3Sj/2B+POtpdhTL4HKJ3w8YPYwUZzDrkup/ZilKBjDZQ/Ra/ndDc+8XjP3UdUEm8iYivEo/Z
FFCwRWCwiyTWKmDRCGfgs1riod5YQ5x5dCPhIEkFjtSRW8fauMGc8rFRIHStaWUmYiCQNn0E9J2W
GlU6owt/76S8o6OtMzO21G4LCaMSx81qfbbbUMih56tQ8D+dix/OyjTKwrd/tHXPP65FDfyuyu3D
T2hxs8ych0HoFu9FgpbF4mzpTblNvlZL1jamuEL5e7U8SLCoTjOk7zO4dQEj+FJkb/Ge6uPPHDKo
8TK6RIcPZX1ZVFdI892gJ4mRc2i252oV7MWpPGXM9CovDXK/5jJyjB3zkbTxQvoOnq4VUQKkhOMz
I1v/jXYRWpJLQestXffhwlc3JGgt/ci+0g5ztoojyyigM7Fm5a/CJlMhE2lVulf4i43qVZHsf/lR
sIP+5k14l4Ed3BMnmTLjvMUYLq/hiYYNcff3Gn727sIMFSrT0F8+gT8j6G968Hd4qbGO5+N9Zhjk
R15IxRT/833zqvjnWFpLGtZQH0Z+RGViDdqIdgipV0S0/twGBedyv+Qhtg4Q15gOta3hnVWXhd8l
POyRHlUgGGHfJdrW02n0cjUQXCCSsIP0G62jvrH7OEkhwIuHF8ExjXx9M7o0Ztb2TLlyz2c2FH8n
R7GdN/xomB7gNgKLl6LvFb5JwuD1q4SverfUiOPXhpbIh3yh8oNr7d/AyJOnqwb5kPsqxIU1kiyS
sL/hyDGbFVLzIt9T7llYVp4ONQb0Q8R9j97P+20WB2I0/G5egcFiGXydE/1PPojmqODLcOJIk1sZ
nO9XXnl9rLAaL8EyVhXYl5f6jlnZJ4Y6P1U76iUgjgyhmiPmTh4dm41zMauk6xj63hP6Wq/CAzP7
VWDLEp2AKibN8gOM2cDFjhz7qN1YMacwpJtYn6HJWzxyswdpkWMpxzHVxdzJt0z4qWAbiMh0/Drg
hAWuoDuf3260GF9Yw9PNzZXhn7Yam+zpponmwXUpm7HeakS/p9PwRX1Ereljv7//TynmkzO/OjfG
73Wie5ojwouP//MGPFCAqeFaPPE6X/zqnrYDJWjpx2oNPGiROhJKAY1Z7rPbf4iv1PdHH7yTnYT5
ne/c5WZ5QHoOe6KCSI5Vahl33NSgGyl2rne08xEwWn6bvlk+R5GeZrSbHagqVd0Us7F4DhkOXYfT
6faBjujV2hfm0VunooCPLzPAc+gUi9aOMG60Vk26K7hMD8O9y82rP4LR1udKUmCsy5QfPvJ7alWh
rvJ0SZQ/AklZNljHeCRyU/3KXyPtERDnha6uzTZCF2GEijr8IoOEfW2gIGOtOfuwDrojX9nryIa9
DqPxFvkSNfvtSQSiRMk/P0y2Wa025qDZrBGnkflUCeGe1FbywrDPFrOrDCmZSNw2QtK+INtIrkFE
bqujUfrzDYhLX43rwVCjSoDnpawyTUn9NCgKWaUzIqmk6VS3sYC5weU0ixsuPeLeoCRTuqroHU6a
szmcz4Ik/KYgLrGLSu2b1/jETsqeyy0BVzu8FTImBhElXYU4gqE13if6unyUfBTspRRSXGc7rmif
o/QxSTVLxrdd8zKUNVvzJ+R/2BAfnao5s1R/PHo1E9UamOyP3P9YAOKyLvkzlcC20zvp3Yl94t0d
9IDXIpqisuqt28koeyCJlKFpqx/10Z7zLvTSAG3V86xNsmRYCSe38nUVKE0HlM4Bi+bIvXOoTJ5Y
bE+LCk1p76Eo4wBPpb4zHxZ4aSlT0cThjSVMLfadL7M0QUI709F4YEUhrvcxAFLTvBCxIkmJdzUa
wahfHjColS2LFRhjZeWTymH0UhLLy+6uGksqD6lgRq9HpTFXuLqeVSnyzCnJ/JAXNbs0dUnfhEGr
sqWnOkezo0oKdV31Xn08lI3WRAyrspX7O2inQXZfKA5S22NscguyE+O+8sEk4DM9cUArQYTEvqjz
j2zaXGhUL7o9D/UzvRk5dYBulMPq89sIbVWNXtPru1tjcgoUXGkKIpdTvldIvb67mAd187h3ydcV
665tMjAPc1Kpsa4c8iN26sZf+GYL+GP4rF4x07Y4lWBVOQY0whC0bFquIzsKvV7brzjEJqOuNjke
/8muYjoclFon+KkKTL37tEv3SJC+4jU8jxmMXTddsGWgGp/v6ZmDhyFENv6A+aqEoQpf+1pTNQkg
eppg75xirRqUrkBFW4o2mItkBsoYqeb0ecuMB5bqo/ris8ksyhDXNgJOVNbeWMei9oe+QJwrwpXf
gQsDvoq22Dd3MEU7Y1JtCjJ2+m3wZYgsqUfrB/HYl8se+HGJSQOdH38FsHJLmYJr8M+D3hnjQeCC
y+juYL80XgBgcERSE7kjIK4OYTaFw+1T7KolkriM/kY/+LlUN7iUHnE0TJvRGwRuoz4U7pTb2pzn
YcjSunPhT9T8zqQhWbhJW9X1bVaagJtmGdSPV6uVwaYCk7ayFR5UPEjw0mspMNadochTdonzBeWt
Dpu+5yWEanBBRFOvUAa6J/7xEIbiSyTWF6Kuet/RRE+B50UEdjmB9vKNzvm6CQQ0OfC2CdwJKU/n
Lsw+FvZrKoJLoFqtrNZq07qdBVJcJM57qFUY2O/v+TYu31sKF8OoNhPgo3eTi6Gledos1rTtY5YQ
5Rm7nm+sMEQb1eWszlvzpjEFJmvHKhwSSHrrzb6PRNqEbwJn4GQT8rB2V5l3V8GokRL5wq+kkTSD
RVNcWg5lKwgzsDZhs45pxdV14KXQwpBt0DcINqVUf5eeH0d/IkQcKcO61Gex7D5U4/VMrA6mQrQK
PuzCpw69XDgiY+ultDrr9cSPi2Q1cuQ4F4IgvhDa0lcnK7q6SIlGm/LYWCZCDJmcZ4Bbh6rvVdxt
1+rduJUngaLchELv99FYhkE0s4u7sEDD1m1tR71ixSz9Z18RGss2sQ++DAh2ZjGB2/L0tVfaxkGX
CEdcYEw7FO8tXleAcdv/AHwXeuAUDn2QnjgFzWCKcHM3SEhLKhIx0grD3LSX3XnKBOkYzaDrAV+r
s4Q9vpZOfao+TnGCcyGhPngyb1ZMrT6z/mHylbBbtuCzPrzsKskk12+XxwrgxnvvE3g/ZyVR+YQP
qXEzoiXR6ovEKgc19u0t3EeHZv4tTb7GEt5Wp9mNnih+mCYa5kUZeq8uLSQdB5feQCP5NeqOMhK0
RqRUbBUioAPaROS5xitu4F/WsP3Kvi1xxuIKVVf3SVpiVCMr8hXgvFMmU9yb5QwLFql3auEgtJfg
mR5vyqbpkJNiVJObSaW5T/CroOnXOy+xkF7bMXGYZtzpcDJgrxxGf5fMTphXCL75/2y2i9BVgCO5
vReNp8cwmZGAUq0TRXA1YXPlxOCnm/NdjwBE+oyhPtS8UW6TKmnALzt3Of8c0tqNZdTfmkWdr0nk
rdkPYVGoV62/tzVw1SbAX4Cp+iOaaLrSOEYJT0rxvtRGToIBUrGefewc7aKKMfYd0q33JcMOGwUT
ljHDCwfDExjMtlGFezfp8LQ70hN01hP34YrErJ3T+MEy32YVSDtHtFcuEE2fkqaXbJA803ie8Lbx
ghflhVpXbdxt8AIZwzBsAIBBwsLQRk8ELjKRZwp026rH+blBXgzvvpIBBf4Rb+LDx8DEinH2wICy
vNuAGUi2aurqsnATk35RBC2U93W90MG/3qg0x0O4JEX9PxMNtPg8fMxkv5s7nDXCk4GbAzTIGoFe
EdLBJsvNLUtJHRvVXkOE3IJh3dprW73Klawsy+y/sHmvPUfNTTT21oi/SqX6VfQXIUHyKU+5Udj8
NYXy4KkDcmKS4HtgD9krVuQ3KncQuYcck3oV8SmT2LI1PvZ7Qb3uXtYbahmZaResZw0U/FesZPq7
ORhc52opelJXMbJWtyEk7/swM0o0q19Uzn+AwbdfosCZVPqubp1Hs7+OYc2Pq9XUqby5RgjFTovl
seMyBYJuNbdea88KOFMDCoSg+l6ErzY8vYZdCbfe5aMp906PdNJ8OBsbeNhmWZGt74D/G5H2Cb7J
OBrhIOvJSZug+FcpDFWOHlcWUJbuWeT5y/uVYkh/wOUDoZwvTPqPTuZgUH6O1gC8fWgotph+bLNe
jI88u2JD3FTnO5s743jtjgaor8cOMrcDw9AJlSeuEuGdRo48GQBBno5VF2MquaVcZ8VTEU1ilC0a
cSmXu0BE8LXQJAwQDcX5Ws6b1NvKkoaLXZt/llyaNIN47LDqtoGZoBnkWtDhoz+sEsNXuV4zolGS
pF5AEK8lzSHVmBg+V3ZHmroMy/OTSHTvE/hbKjQkRWSA8dnsxknN/ji26bOu6dlv/D5kEWBIB5rP
uv91E6+eofQLlymn9KW4dkqbaJt4mFFUQYf4jQq25qBQZ3W5cuy0/S9yQH9c/aYXR0K7MYkwPUDl
Snuda12iXYd8QZm+arf/ddhNmVLI2N7Utn8a4FGuU0QY5WEJt5K5zNGl1cKvQk6nYQ8T3oCy59sK
pXOka6Ov+P+4DpQX80lsAljejCfOjCevV8dnQ4AuZFTwflxxzSAOerxJwBxsBC7WWEFpeVrCPtH8
MOJeyRakNy2YYRAwy5tO4jXjr8fFn9RaNR5ajXXuRPO15BJJ+tKhxI5u0IYqizHQQjOQIPnqQtcR
6+oZ4oELJ/TwXYj6nPzcN9sI8UsKBJaStFPRvxHdUwB3stxapcVfF3w0PTgyntBZddsv+1ZZUi9K
uUKYvcXWHmFFm/LCEVi09hMpq4rL6WkntI0S+OljquR8N7woIu93nDWjNeBtfZv1cWQBx7AD4yEI
8R3WtDapZx23B9CyQKeN3UPqoVM+CrkosoJZ5/cUykuKtRSE09rUcQDyHW1FBbMmt9kRQ3aka/As
DFbNm5BKUwPWExXfoW7VaZnWC+Dv6+UQJClSHHnobayb/1gZHYPQSjUDF4LyW8fCAQPcowhhz9gk
KJorMNtVrVpxSSaE6kMGCxOm9vR9UetNZ8fStOOhEqYnjSjY3/kYsIkeZ/SeH+9EEqDKPeP5sLvT
2Kmj5MsiAqd55uvTi6n2tsrIa+JK1lgc3Qw0KMfNMZaLLmqnSQlQncfZGrrYDqYMfb9kG9SB48LE
CqDBy/hAuNuULHZFYCVZCMIhUrB2RgebhzFyzOSi7mlgLKUhD4MyC1yYP7uk/QJoDQmodbkvK8k7
92ainBjZvK9Lwh+IbMhSF1K74Jszyvc7WMEqpThFWaLKQ2J1vszMhzxwPgKFxPCSYwB3wC8JUb17
hrJ0yl2tMULUxPdI+O8kdDpR8hU2vE8gIqG/OgaNajevV44xjhc6xOJIAR8C8i1f/hXg5KzMnFH3
/Iz1HoxDIUFe1f/HTZxsZVNcfeGMvFOARPWaHubiHXqvVxA4iLSCm+u4TgmHGNsDoOYESDjzsoOP
tbGXMSsujzqBWNQY/jzpgaITtvk+ZH75FSIG4Qiz8FEyWM5OuxYDOxpEC/z2rGgzALJy7x8rK8ps
IMLqay1e0Gq6njKUvZMnzvim8ovGOVXPwTDcTtyb8g7IFDXgEyknpnwadiFtwA7WpyvzLmZ1f0k8
7aK6W7eGcqK8zxtic5yVl2Cw2z9OWZKctJ0xnG3chBgF+m6sGGZZ2ORwjw2ZwKF1nYZsXSEeaRni
b9zQ/D5yshtPDX9eQorSMZIWnqC2s3ZV8xTavI5P/v+p/sShiTgv4ARWL6k9ktsQGXqA9NO/4Neo
M5DMTj/PG4FfirO+bNQsRPUsBY/vIOLsH1Hkhl4LFPROj46Jy6S4qGbIUszXjKr1JvZxqAC8Qb1B
MjLYCjG9C8vAAznl8Zh/RnlRJhdQ9EYn9CQJvJ9xM81weiUTet257iMtYaftWMz6095mfBKjKrF1
4QNMYGS6ouwVOxZl2KxRtKIYhl79IuA7XDF76ERYzk1SOEq3L2m/K/O7Pvny8Wy6dNZ4GiBxX2SR
v56hkhv/cpyAtv1ZxqOPLU2VkBfP1mZ6r7KlkLKvpouwBK3M/T67K5bPx/MFou9zvxt8P3tFdNXK
M8G2yXX7ulzt6YI0UT2HNZRkml7lP9IRZyppSzoS3p63fCOpwaNJaA8txUUtjWuh89NITUAaQe2a
xEj6cQ+AW/F9k3v3YHTAP9Fy3ETS2Nrg2xzZfHNbsa6liKcfdvAukXdKymtRQ73/AWWg876o9kXt
7DwIjjbRvdNX+RZuoCVqEicaz+rNIYOhcbz61rS8LzRqeHoePx/nU6XT0TGYWi7zCoZKwxADapxW
sCA2NPur7wZNfJqXaR637m0r6V9VV3DtFuPDJUBCxpRS7Hg7KuExEdJ9fLkObGANVP4lF9RTZlse
sADiZH7Zq1gPkc94GhelMs2yqk8OadgeuA2smKxGwZBNXpbAgR6npX7O9lJQn1g/HeLE+YbMvt9Z
SzQNwIQMdHGpKCecVA/kHMXzrvSV7LshSBeU30rVVDCSys3jsJhVndmm017byaBdTKfcQp+KJOnq
MMXhBEmBlz9AXsna5abd8zGSL3VNytnMWPz2b2dFCzullCaeMX5t7zpeMFqbmZb7yQbIL1cnocGN
P9m/sFntvRKV+RC6+3cVdjeBtdMh9oh+MHIWA8EnzfMw6iMzQtbYEU8Lc4f/voBum/r4N9mSoG2n
+seqZ2Km+SQy6wASjW2IrSrlX1Zpl8NtZC7oriTVl0xggRQmeUoaU4Xuky8qz+zYGr+/H8aMgdgh
zefGSxs5JPi0B4811aPDZ8RcTd+5usJ9XnNdiFz6hTaotyFr3kEtHU3MsPQum7DGnIdYJ0r0NJy/
UZ6M1w7LL4MDd4hITXzCByQ1Xhm/X0qN7f+qSZM2JcpKHmVSquA2Ulfgzi7lgirL2izXtcgxp1H5
yMW4vGLbTtRlj9erV7ao0sWEo1Pyw5zNsAsE4cRtNS4+DtWYjGq7uL9/pJ44YfwexfePrdS6fMAI
/ogmz563CWNRz17BJZX8AL9mxIjyzLNZ3/A6YJB+pT2oRyqcGhrJNuF8UpQLc19OhAkP27pt+Qam
LcGzVNMoLDzanZFMMhpoQ5q3LOxM7OSfPG5s+SwsJHeXDKyKfOEEvAHgiU+ODcH+sY288OhoUeAP
T0igpbcgtifZl+R4jvFXBUFi+ixHN/1CeRdA3UJTyGdY0eFquH1wIZmaXZr8tN+q6hGUgK59qcE3
KC/bkXlegJ8ZXoB8FDDbPsUalbccIVaFPcxl8HBAIuGcjNWT8hAjd4T+T72Mnw4wyojCyOsOJX7E
sI877FQp0dRmbkHBorZ421l+HqBJxKo4LyTw7sxfwgVQcYGmuthp1wwG/mfhRoRBpv+Ci73dBQoP
Y1owSvGdKzeJY+297bJaX4B+F/rrFh23p0dAnZVh+boj+pFl5mmPtyS0/Aty6mcgweVtEp7rd6TE
7/IJrx1wLYHR7Wh459i4kEXEAgQiOLQDYZ/6uu14FOyvJBoZRqs38sE7LhTERlupyzLM1eDybFFl
SKxfIsTlvaqhCbpd7T4CPTPWdzdrWl0H1wOoJ9vIvfGt8Z8hDvjhhEPPNIZvrmbYp7qGcKGgaXXz
2nE2wavO0bjfhfMXMOrq2WhG7Compq5+BIA3W0knWkX9l7wmWix37MteTDGM60805Bv7FHLmG3fK
miZ00UnosUN53oGlTV+wbrb0qsAuTW2KTueGQpdJ6kdQyEA+bCccl+dzlvoY9Q8np3AVib0dCDM5
gKzr5uxeoWvqCWdEtVSl6ImqFCqj6mG+dlrHw04LX89HdRi7brE90kkpAMaAQV3nvkPsGiOD8lj1
G1YA4VXxTOOyH4xbRcOjbVdKJGKLLR3MmFAOSWKyiHARI9jIo/psqhKaAmr5+WRGc8Rb+jK9OYxa
wF648qGnuBXBWrSV3dYariXI6x58pIhZxNq5sMZbovO3At0p5i3nJV+gaA9kaiTuJ0nvvS+oIMer
9tRwonIJ+qj+LmaGtxJxN6TQBY3xO75/TKz2p021GfXnzUExalgn2oZEkKxUaGPO0lkbcP/PkLsT
kovtkeS/VM1uzxFudt2DR5nIYnFg/bsP6jGwNjTGJ5kiy2QJNtXzUgbu38JC8UDvCeKh9/3P+4JP
v5mEa6JZfwWYYajd2WBasPLRAF8X1FleyyNofH752KIpiAJrflhkBaqhQqHCILIGwy83mhWK9a77
8he2WRKNSGCCQIgPBtIR8MXxV3GDzRynto8DU2L4tag3s4L0sic/x6ZaOnXn0js5Kye1yUZ2MS1A
GajG7IwCQ3sUCzX5eBhDJhHrkrhxChR8o4puup1LwhBMWPZjlWemCcuXCOefuBFXz9xljAfD387X
MIdlA1SvDOeZmYSemU56bQLV8gKiwKJg4ppMjlzu5cBnY83pXm9pWdYLve9xb0WVAUXmLpnee1mZ
REzWAsX+dW15yftDXKbL6Z7O27fpTw/6AYh0QvH1h6qT//Trmg9TgSKjumYgKL1vPSfwSHjni/mg
n/CI5iIbNrqihUGQ8riIJNYJIDt4EXf7dc8sAY+eT2+J1i5bQ8balkI9un16TT1hVoaz/R1z9wtk
AGKIbr9T4i2dLuAR8J0n0GO9AQdaQx8vcrK3tI2EU/0IpOO421IGyllmR3bdK+5NyCGq6kKrBHpi
Jhlw7PGq7V8zz72P3+9HN4GdgQeh1zDi7jBfsmp9Vib93/GAuVpLPfvmlype5EbtW7XbSkDmoBPI
RMzzwQTnY6F365AMmojCeuWRosFeye3DQT67+9RZsHDVJl/HUNnSIXzF7hnd8zoPheaIji+YGT56
AQ7ba11V9oAnEoL5j6hIifmslEZGtWEyQpGoBUsEHxA5RdKVCzeca5EZXJtrhk9J/NCUob33tMIG
G3bWTlteAWY0CfWbvSumKc6G1e4Y+FzqpqHEclWlNLY3zHoA4zIoJMFC06lcfCjTC+dJj7ocaahP
XG3x7E7NvKYZCGwx1QBslW+/2GvVj4chV2K2uQMd4E1IKTZfnvXovqRjY6K5IFKKIE6U4tWY7ggJ
ToEL+qiOY8Ex7ZVcc3I0bFXccctTvMPbfwRLryqTQiRfPyrJqJzm2ui3O1ZVdjAXbUCIurBnz+Mi
oSVMzmFA+X1bZd0UtXsqNv6pOZJyCvUtYdouaQVgfVOakMlLsNmqqc2nrUh9tO7sVK7XXcaC+IaB
vNnBgQndAj7dtsPW5sQOfirhDPcDgSeSeAjRFDM9f6MNzsRF8zULzWucqRR1lj51MOY9mqdMe0Lp
serQ7tZZU7hAPiwyxpnWfAXqsCP/VGWl1DIx88kSB8g8mqjDQBS5Zelk6VdHfZUlJkVXLzfrkzfm
9TyovKWnnGWTLv9H65yTfDzJ2YpPgVAhE+yqscSSiUeiZa6L+5c4Tkbdlljr4Cd9nIQ/0v/OzQh3
29Rz5htZaXhVHhIGBE25Injz/2opvXD0HvbxjXQKzq+xzHXu7ax6jcYzJEs9PWbGcGxt/jStDEWp
uodPhC3PkxQZQk/IjNtXhlwhSBpZWtlObXzzF1G6LNCLpG5BK01VFvcJ1T0WPlPAZw5r+/cpPD+y
77RxiCqoUe4JHrQSWvg26n/haUCHzDkYh/tSw+557CvEmWgXMzsip6zHb204XBlwPuwwaijhtzvo
sbm8GH70gf2B1I7qqZlOVd0UETSSgm+YIL78LmwaOmJnzdV4EdkCWmjlfVLMgMLB0l2LiJa0mN+Z
l5dH4Wqh/RkNWXm2e9M+RfLH5hl1CcfSuAHFfIu5imSd4TBXm7WTnDSkSYdSxXKKKz80137xrsg5
JsfdMEh635qYSdz89XDSqpEHun2zFRK2enLMxqGPNhjDXnXBKft8CDiEaom2mbIVH0RvpDmvsYEc
8/GZDAdzRU7+mH7aqvmn2YCTW2vNhvQwqlDHlujvq33HMqBQPyyfimYNO22Obt3ShRAA9t4wb1pm
Q0l/8wDVoAMSRMhxbc93RLbO4WEEuqvnoFBfmZJxddOXzdYC1hEuGMjW/zKJsYynvHsup3ps7RXE
sv/uhlhKaaL6EMvv8P5W3MgVh22w6sbFzPQTxNPrXbwfRef9R/QVw1EnvqKQBa8DhOlBvi2quGeo
G+e1eAb0SfDICPxKf7kBMmTzL16gMTH1blIBK1DRnwcXIuOT84rlqHvehUfxP0h9es8LyTmu+4Uy
IcPs8lZ0EhZ2LgoQc7ItVjegkwwn/kD+QAyCUZpQzIijQrfop3VCgZM8a9KA52ze2R6iW+eUNJBw
HzLWPMVwlFYVHb4vF7iJLBeqVWxD+SJGdKriNpm4BcB2DZBVB3+12o1TvB4+zznHqLoD7Hd3K/NB
OkdfchWRSNeWKnCp3Xk8L3n3zRJ+n6aNK+P6WJTg9/XKlsr8Tbc4DjTAnI5GVGe1IsSpVNq97VjM
zWl8xl5V6qiPmX3dzN/PvKwv/YZPMIvAfnHRw/5EJm4qGIOdki/JEZAnO8msfoJETm6hHXTpYjv7
/hBPyyFqanyCzeY0KXFePwR/Sz+ABbCsL0HIfsOrlmno26BnnCRPNCICm+QaR8TehNPmc0loLJey
aT86mxgtYlsqljxG7+q8JMMlqWXykvBVCUHjJd/ah6jWAx21zy748Sq4Z7h7EgGelHh39toWlPMH
Ny7JoUguHX5jdYlRoEflmf3EcoHTXZ2LrlK9QTq3KenHYHUoXlm/voW7nTb6s9XgTciTEYIIS2c6
nIvAQxp4xoSwjnmPj7+nEHd+/EKRzFy9VnY9nv/vSFvPAwu8Wac5gWPdObJ2z9wYffHChKe2HjUi
bAf0IHmfk4jDdOIfYb7YttKm+I8XU5WW/kMcciyMy3dUDnmlCF+XBLoS+gpHeGKarpHU8I7uv/QV
ovMwzWwQPBd6bh+rHm5dpCoQ+18wVU+PveGvQcNe/9ngxOD7uctg9ZXd/h91TgggvdSj8ggurrcq
Byjch9iQ9nx6R2PJqZcV31tC3OidnFhMQgXfAib+ZtVAM323I8Tc2Tyjxfn5gyTZLSXEEc4wjvKz
trBXA13nt1Ce8nPFsiLVhHREHx0h5uuMDbCt06pQBh/qTIB2tLITQimve39mR1sA8h5dnsGypBGc
3kpGKjEYkK9te9H7G1eYFSlIt8rpqapO5KcqH3xcKKtzKbKS/+9ndMPAX772ulDAEaemJ/caKcry
+luvIObNnwToj8CCdGBLP+VfNoyb/Y4yL5oyTMImdsdJ6fV9FE3xgzXUj7nIhRmx57xGvkcLA+tx
dC5N/y/dzc7ZOKGluV3JnO5Gt6qLwl1RQHPkW2ZnrtGZ9TY030n5tooLKFo9Vy1E7OhjcpdpyEve
DCeEbp0ldrFn45Uttn2FEkXlBKs9TtBNwDrZUzKZBDmPL2/uT6ACSVdG9/bSQa2EpM+5nDbcOtFw
ziC/0armyfQSEtatSpw+70lNBOJPdQtT1EX2WN6go+oAHCoYkFnVQBcDAYO6mHaEaqDr5couO08v
dU3ikvClKWAgOe4ygdC+hmBEa0oYKolu2SLLlbd2XbPrCcOk/dsfvDQPSYFbEvAOf1fm3HSrO8Yb
bfg4m9WoY35tcQbuuQ3JhwV39Iz/EXgzEW88/Zc2hmOCnwM5DdouNU6iJcSV8OuNaGPdrsBa/7sV
hMdujSqmPODcAxcc1doikESSgks14QI9FtsrNkHpqpjsqCldNAzXHX7oVlBkCPcq9j2AG9GvhGAR
sxL3n4WE7b1o7zjIIWlOV7N6x7TWqV7CeC6UwrJxrWb1VpQm50cZ9xmUhSGCXf9UrWJ/9tZNv/UL
vJQlQ3ZpygzWeVv7oXZAzgb/ekaDN97al7lGMC6BdzdlDOuzdCogarRLV+I6EVEAQ4Hl807WY9MI
eMQrSXMFty5+YDWWvlNGkvVYHmoHwo7CcS5kEcD3ED4oFrTIV6gFoq2iJrT8Iu/ZGmOTyxqLhS74
8SGHBudyMDW653Xcnx+rrDyPKvAsdjZJYhs9uHoX6WhojCf5QX/Kq6RDkD8SOp6NfXaxDH+sd3GC
IKIau3KDx6xCphXuXmbWw3wkWpSLQ97BF2VQKtI2b5tYVuDCn48aA5mS5kFZPdSJSWMMaSrUCeCm
RDOPV4kE12FdFuy323NEDdV8LFMcez+xSf5ejqRWFPQh94P6ImB8S3DVOic12yFB9/nqOmY657vQ
hFmFj7TrpFyxEkx4f6QqhgfGqBhkb5g6H/4OGPtv33kGs387ouDm8KOy0Sx5s7J2aw2SVqkruUyx
WOtpfWC0gFxfp3x4YwISbclbYmqs36mp7XalqgIOESvE5quSH4vio0RhwVnSh2KYqrrXRhcVvGrB
z5NLAWIGLkfbzIX17NM386Mns9eLPy1AB4NRCKJZI8I551n8d+VlJInjDp1ITrKODqi+iasNdum+
EY2xhPJFrAmCfh0rNd2UYv7Zaf3MSTqJQ7gWYze8bNqDim014LsZUCrpif7lxwa939wGBQ0wRkRX
OpZ97PThEdYtw/sXyYw6rJB+sRAXYQNQvwHQrBKaRDCAqtxl7a6n22sJ8Ql560ShE+HKm7bT5xus
I+VGdqheJbrJy/OadIKALXctjQenU0T4Bf/MVMgDLuSYOxXuZyLJWjUmr9du9XhJppQCpQSgpDBE
jz5YnmXHRD+NIQuXqNUOUwjFNqG60RlmwG7Xln6QliIyC8d4uIQehyOHG6rem/7fOYOIN5z7fMne
W/3sPu/zA3hfTB4/b4Ih0WuG4OAl4d+E+gdNdlnjQcUEfmpy8vaVaHMjBoh4fiF1dfKrs3FzisVQ
jKV3NOlktmdWM+aNTgPn8OBr/N+68YjMgruX9rkbNKXvMF/HUrrvUqm+74mkLWEQa2LwuBY0eMmQ
WmfJXa8USZKJipJlo/i66rafgdwhzC8AbrWL9bvklstHHrSwIEEV227JFRyXesva/rAiU8SjlIHN
LTOEhmbg54BGL8XkJLiLlfGFShCsE8IDR/GvHKdL3cERHG35MjWxz7wYBPuBl4aIlt/O3s4TNd00
D7Av9LCPksF15ISWZM+9raFnL6tuwaJB1bBls/pVE0z/5VxVCDGbkVS8QHScTTZTaeSRQ2SqHf2j
aCcTo+lJzYHk7C6EQiwLKg4sRFx9t09zBclVRh/ypIRI8P9v6/lD5l/yhStPZKCd4KLe4DNfrKf3
rKRS9sZvhiYO/lTYPXenJS7HdJOsbeKKsadAYaQY9kk702jUyQBTtctJFJKI5xi+j2q+9vVUup/6
a5+j41LbkAKgw2NqxvkvrcFJiWpSUUWpsI/cdhOjw5rmLbopDXmPz9M+1C1ka2VhVxUN7w3MmfKe
skIL8/nl9isavaVC+4gYaIP1/JqK6S14a6NCa8ub9L1/92iDFTfTBzVPcfDzbMLTPxp739xgcy1P
Otz/CIP9aOI6SU7FQj/vb87tgepOV5bhqxrMJRktJJoenO/6RmHAJZa6yv7kJgyiDYw0u5ftIxDg
4ZIm6rIfDDyzfdBLvkvMEOhDX4t6qeQ4mzFaO6sc97hGzwtbSBygxIfXAXPD/w8dlvxHOJ4rPFDo
u/miQzkiBy0mlJBVqqI8ehE2keqjojOgEY9BGFx1KDPspD+7w70m2g8qrPy966ZOsWTgKsKSpPxM
xNqBtp/3+NbaupRkEhZoorszu1mhSt2fJjsb2w6txRWYTmbDkb+JkWLAKW93nhJCf2JjpX5G9TVA
1GuzNZTdZEQ6kveLXGp+9rDK5DGsRar+7kezVIqVbzd79ghYhIX6XXr+ry9war1iI/AhR1paJZKb
nQG7LTyXrqALFOYXnM4FRPVLSR17DsjDAIeKUzJUGish1437q7gLOv/+7MJ8jnf0zAaKjrNAQsPE
cyPMOXomiRigKzkEqnOtgdh3dN+KPdVuns6ISvpTCIfC66xJH8N2kjLOlkQtIGxTmRCJFvNwCp91
UOceRGJpnDcuoZFRjYikVtcQgDu+puktKIdISNvAREGi7H1J1DeNNS1A3TyQrHolYe84Trm+QiZV
TpjEN5cIBZkhth9Y6nKGRLIiVMnMTeiGRP2t6kqoM54mLih6y1ajSpE76kIMV3qpMHwfYKRr77k4
lM6E8V9J3MnDXA64HNyyGj9cxC7rc+m6nELtrnREijGZQ6JKMfcEotlgfmJaE8v7y3UGBIA4Q3Rk
PhWh6R5gzwC3PFYFqgUrppdmg9OJYQmtDoyNOk2TRDON0nrwU4SkZd5rDHTFChSx3xrUtkiFboRD
ikCBjzA8efNPs9YyaqqV8ikB75UMG0VRwY1jkLOe/PvAYS//m7s/r/41RMSbpgEk60/LPe8iF+BV
CFGUAP4v58LTBmBLTK7hT8VHZPi5NWiZcVMaXr9M9GnbFzw2WFsV7ZeC1qweH+V6RH5d0QCU3f5X
LzGjBq9NiUiePJF/cRwBqosAkLfTyUG4TF9NVjuCETg9VG8N9D2UIKIvIdJSHdlfIJMA+w063x88
w9BUuM7OmsTuNgCpzTQwvBtkVcFcFmJkWUwNuD6Q4MPe/wZzJEfhma9g7fZ+0OysCSG1wV/KLQFO
s7L9tLEeCojCBz6cUjEhpmBbbKm9EuzLt+V/RkjOZvwqHiv54Q7Z9TkEJEr+GyrPIypGwr9Lx4OV
QTlhcPX17pVHTogVFIQdSvbFjYNsHLu699YuET2yjZajwRUVF7VkuB8w3gEI/hmBSXcEnzQnl/j4
8Qkd0Xiu0NA11cp4l77HbbIKa0lUSA8LplHmJYGIDvxYj53yIfPj/v4GH4nNbJFEuneDIs75oFy+
jSuWohw9uYt3RjsHr7GYGcQXurbWQilINy2MOwwh8MvZJupA5XzCMrWK2oZ5iBi83K2RUcT3djvv
pNG0R+MhuFXLBfRwVVrP2FlrQ1dBcAZANtW5i4uS8LYP1MZX+Xj1/38KHnGTDg+nUNaDf/NqG9QL
vprQsPsG6mkVeJqk1pEJDKGpVTxATfebRXvWC5nkC5DBMJn27sa8xZy/1EQA2YrQLA38eiGIxRw9
bBuaFbc/efTVA0L2uQWIOsPxRC//8bMjBmZ7IaNrMD82EErjKzcSuqZcX1OAPdNhIZ9SS7uHp5Nt
8mU5SDndldG+jZOGXydvkETVybdmiB98KyF5+JORBgPfOaurinudX6Yqahfk26AWpow+71UyTXvz
P6TSOMbXH0L+rh658XRxqUEtKsrMpskk6WYd2WbtKOTgtf/11zh8SYj0glivDZbGI+brAQthfWWU
uug6YviEmPa0HyQk+fYWl8A3ElhT9CltSYBt0XO603iqTb7sMNQvF3NBSpLZ+sPKefqs2wA42sIm
GU5ZTg/1yalAGvXnPptjFoVsgehoIH7jcI0xlNg/tnd5N8ZaEx4SY8MO0D6b2EM2KqXfsrOHfXHW
5nweAXxLdgBojXWmmqrolc+tj0D9FpwUBbQhXUPcZUMVA1nnSrra8Y55UlmNI5OuHpB+zpAX2zwI
abZGePELHKkhJUI2gxeUkmzzKHJ5LFbbKyOX+GrKkZEisGBNikfaljXANjvzcoD0cORA4zN5epU0
5Q7b6f1VfyLar3XpguHJsZmVRXnR6lSKFJSofo2OIAXufAlqwDG54oGaQLS/uRCdySm4XNempq01
Fh7x3Q4moDmnUPC0uR1xUr9SP9twy9+RpNNUmFxGxc02qGwNtu2CbZsf2pnZrTtf/K9pjsekQupS
1F7p4oV2B0Qux4GJq6gBEK+jpnuwpbyhW9erbKsm7XeKv/Z9j5sxNJzG96PeuIy6aEQBXn7YSJV7
iZPfrsnt3zF+VQkPVbQ2V/doItsmxn49KrJQtG76WBPNZU6iw2yd4VON3BQMIuXBwmCoOn54ACtl
VwXPhtUyRupMPlbYztZLk3BfDvttUBiTd3vyV0cCE+WubL9Iw5+teWQHeGwjrXsHxQoKgClUvdy2
nVjEVRcWvak3Yhc92qjnGUGVmSZBHiRsKBVXnvDpD2aGRAqigibaCD9u2yHtcBL4jg2hTB5bS+Id
rg2EhHIqbYphfYvKAmtUu+Nh0nEUWWMW2rxqAtKAUZamSJMnm4hdh9+yya3CPZGviAuA1zY72RBE
Riq5yOqV2bujNgyFdW+20x28JBiKenamVxJGR5Uahu7+GrraSb3IlnhvHcQ9afFeWa3V9H7pJZz4
HglRCmAUuTYnFSkPNM+8XKvEaM3VW37E/9u2jSMMVvAF1SgFVA3XNUnWtE/ip1uymQ64zPd1fYdE
Zs0bhLgD5fKB0MRSPFTkyHTq4Y8Xp00fBvXjxL7kQbx0W58/juUgXyDWaoTqadg22T4U5SqyHuPM
5a7s5riHk7fpQAB6gvuyNl0Vb3ko+k9gwenRMbVFxXt8M7cOGIjOd4DrLMCQcWPirFSuEwzevx2l
eHO4f8tmcTllCbPJpVjTeObVmahDXERXHj9gVV4lJjWA13JrucJVrwkCiGD9FwGJXh1H4Ya/NO9U
YSiN0zArNSIYN1pq/zkwQlJmc7PeKDt3NPe3EHJzrzAWyVbW/i+Yq7/q0f1RkyWdo8HT2O9jnase
HKV6VtG3SoXq5Ia6LERvBCVgAbk/0Bs3TUnGM1+OGQUEaFF4swlkEREiYY/d2Sx7cfkgxHAkxx8J
uuqeO78DK5UVkQWlg2y5jv+/lZjnvJRtaqFJMdh9DMZ8f4Q9JkbjXOJN2e+E+qNqh0olchz2/p/+
KhwB3QKv96ZfXMKNzfmPt9r/ACMpmw021ZOANrZi8HBEkigUzlVLL/hkdk2kXM8mpi+PROxGGqtt
ce/oPqyeWOmaayfzM2N+pyv7W8pxU1q1TjGaqXwCoeF0tn56RLqMZFJ1jZboHFkgjBuxBUUaugql
bTChlahnSK4woD/8CX+qR+VR1lLzzntylBdmjLIztFhYosDDiEl0XVK5rGhU3vYvkBVfDD3mNedl
spKG4whEOzEBFbMBfYTRQ5b0a317KSg1dCdCGBKJbwUwVDWEfOTBrQ7DaYP4WIgCnAPPKL6xgQKf
f7c2m9Iee2ChwGs2ENcS4fHxdOSaN8nqMPhDjNv6wbdKXj4XIHsMgESEQ4I60Ta/yvoC/Ik23onE
A8YGDbYqdtDDC5QWMkDTBvccEKS/ryutqMUEV/8ozEpLlzsAwCxJeXQcsrzU2zUmbcJOcAk0Y6GV
5S6uQ06pJSPoeoxiMIRreWN2C5nJTkxgdL2apv7V+4Hq3EsnSf1l/ilcOqeNYtpG/VxQIh2hIj8b
sX1VUlPS6X85KzACUgJS7yKsNumMOFKvjRFViEE/VrI6wTfGUhHLZSTNnABOskia7//6kRjrlDAp
gDPxpuyXWJjSo43DpRfBCtkkrmDONlDOjQakb8IUmi1xua3U3QlO2HkRrP20PBPi5VPrlMYoZ/HU
H8YLm6krLlPem4l15bmYZ+dgi9zaz0c26W5kRm0IDVmOxdDOPmTatpNKN5Nrg7dHe4+nTWQ36CXv
fdOPaU2d+cgO/cZGJUko3C7l27EX9PosmAzNGsxF8EKAfFEWEnyLLlZumnBJEbO2fizq0NbP8eqR
yGrmO7u/RAowCUS1fA9jEWFoNTFapeT1iZNIMA153DkQsu43ErkuK0nnq8gqByIk0STbnzJheN31
dC3xOAtSCs5L+ouOd69ldm6RzU2jGIOzir9vp6rKTlIN+TDALOJWBr6dyvsw1iIvKWCAF8dW5HK+
MOUqlTooZsXgwmXEAEuS6/tlJ0JZXHo//awtexNNnGPsRH8SHZD4o/JJ0G0qlmDh5yv4CRARv6eM
lM/EafykDm7EKW7ppR2ix3j1tBfd/G8TSfaRhgIUkpIjRLEJagpp23Cz9nzDrgKo03hBfYhY7pny
lpxQ3Np+ks0dPgOWAwS0HPWzb/5osx65CIUj60rt+nQ8YJtuBk7eXKBcXujSKN1xRI5Jb4UT1jfa
tx1oi6mNr90LZihV97LcIeMpvKXvWqHDA/YSsepmuGREhoKX96xJB0PixsYVTbLZUUb2Co6Fue00
UdxIntCmFuWJfkjv32aFhCb4X72zLVPD+CHPnYM57hH8c6p9CRgSetin2DQ2btdJdKXanXQAtAEP
wR2vFdjhn0XKStEuB09dYtAH4DKrxZvktghPjc+udMaUE2SynArcrI5tEOo3sFyh8c14eVpzFf60
zfy2dnnwPcGzlTNkPiJtvfDEwUL7TBnY8QmQ2yMLGvSYhpl389BzUHcwnX341Pu+SX7EMCvxcVG9
imIm9/l24QWyI0C4I+KVokPq341U+X673Mr439jd/xsTfrscJq6P0JcbZpKrHvP7cEamx638G7Ux
ZP73UpBdirx4r8IBMCB3ElQSARlvq7T5sv6zwInOF+aE7kHvlb3QrUFupXFi7kHQV7zM0UYWaXeE
31KzAs8nnBy/tscza7r4TPmDGnwaLqVzOrH6i3KRtA/Th5tzBAGUfYcS8vUxvWe+LJ21XC/nbU4j
hWMoM5mD/pzMzMPuIvHhEnBjOoMNse71AuL+ZoNrsAFPw/pt6loOLH5QMH579ZCrmVOP9meHK01p
4EIJffafC42q9m5Dj2vde7gAuKVDA2UN2HZci+6GlxZGiROjfvuJaNRx/CnThMaXZi5W4rNm85pu
EaMVfFbIrc170a+/4ro/4oCYjl+Z205cK+7batWihxfVc5FSk394SYCjFISw/JdZPrYz7MYkVMsu
IXGxh0O5QlB0/PHXfe1G6q5dI/Rs1xgnBJ6UBqdi87z2soXeema7+8oHBP42lBP9Kic8CzSvGagN
UZFLUdpMcrXjNDnwnJi7+hX7n6OxZaupChXOHO579qEgnnILzOCFG1FugvGhZxIv9T/YlqKTQx/t
b1PPmY28FbhVYtHHH9BK8FFb4/oh6lIwSHFzcbO/8TZsCaxD5dwdIwiCdWbxojq6ex9tvW63OHKm
O88niL9FZfr2cjJGzUOq0hgiW/AtCTSCxGZWTW1ngr6nfOtEuESfmh5a3DzcSr6CJigk2f0EU84f
8Oiz79OGmLxgyMIoCSPgu3vAH/JRogbdo+WV+ia1qudb8UgQiMSnRgE3REFe1LNaiJI7vx/2kfhE
HLpNqlSDUziWdAFqlYzM14cnOUYGgYTEjmy5FMViZxzBzF/1FlJ2JmZUZo6I3j4USdoh3AWl88hE
S1J3HWFg4Ny1WMn6iOvCQR4gqzGCuhVPq13j7xZYOV98vm1xrKwnvMDZ9lYUHASl/slHtnV3jNVa
O/2ZvjdcR8QO0+9P6jqgwdFZYECTZuTwrTjr9HdH+pjsXEoZeWJyhW8ccvJK6ww1NO88hAyLfcDz
8DW08jxKdaqmRZESh00rdtkHKcIUSS3BzXZCAwx3VK7v1elzku69Xc3hdLWsmmcz1xAnu2cnncDM
bFYVecyxENqD4j68rCcuYHopW37Ogbmr9OGxnnFA5RcmKpTEg+kurAIwHRkv3dxLSCQpljAYpuX0
wl+H5CLYC8LkQAIA6miKeVZLbaX78tZhJ/IQ+renhlAG39nwsmdlUGfV3WJtL8NWGfD6ntTx0LeZ
+h9dWTJ8XkCFRxskXktaG9/a2Lvkz87XZr0cjtPGjrOs6EcFWmpiv9qNRKfy/OZq7FOF/DMiuTzF
885oknKn0a+ezRoIt9/KUOoSXr5xmuDzm8sXjW/IqnlQvH4Xn4sXYk8KdTjbBmmMD/i/zqcXLgNL
XsdaitL86MC+8ZNFf+bi+ShR2qwk2TO5amgfwNBSAgAO9D9tQxYQ17EP2d+A3aseE89sIrkgxTGD
LeGDlqtXzb7nenLPBrBXS+wT1pnrjHs5+WpIkFspUUCdSt0JS/POPVaX0zewzxtTVdxoXw44U1+k
JjLo+QSkPleyXmH49zZiwvuczVZyQaHpILXhMIcSt4S6f9ymrH+ppoYFeScdVDwPlFfTn9r5vNOz
QNZKOXIqOh5FX0bmZMwqw0WrDGSOg4BFvBtz9FqnUShKwVNH61JBaseDrowIxsR5RpLxW2wQhCOw
iHQ4YzRzA68xRukF2c+0DdWNBF8VGzjOQBPIQXU/qA1+/JV8ubOw0smAkpnCLQ8Zkv4hM6F0VlDv
rMxyE+nijxdMzmgDAXghc5URc/zxaQYZZtErTqFGVr1k6sJjTllE3Xru6XDXwA9HXgZ8soJzl56p
wqJ+OUzs6ZhnCUlhRmF8U9cXEZ5PKksOl1eFkiymFyq7wNxeMF6u+eWrI6o+8/QwRGmQqn3/3I+m
j+MqzlTUM+XjvKCc4C5ieC3bdMGn9FAvvOdD341WEZAl14WgOgL7Gx55TdD8veLO7bmc54ShRGCS
6kz3RrnEVw0UT3ZIL9QIAjRZFhyNNdG/zC5CM6SR+dpLIXumXEZlKqjfdJjSUm3pJHhJHTfSbalL
xjKcQoLllmlbzY8XqhoxjpBPjnLTXZXzmEH+WmcUaEFBs6tL25kicTIbeQbjTuoAUCHxl8WVZTRa
CXjh4RBE0CIFZdvDdhYPJ9HAbmNMC2zt7eM4FMkT5qNAaL4be9JpIZdiXoweVGu97tBG5mDfilR+
ggEMZZ+97x72tGo5/KgcJtJVUqiM0um3HMaGeDfPqfjkpK+DqPIyyvmMxJ838jOLSzFfbAK/+fXI
CjDQYsDIBEIGrTHWQ7RTDChX30x5u+JmhuhpmVrKU6YBVUwlS74mnRpd80deJzaafEclS8y6QjK5
BNzS9QUBC3b1BmomgZaoczD9FPv8IlbqNdbTjdLspeG8L349wHR7DzlKSMDqCK10Ulbfba3B5NgP
1OQvl9Y5T73x0C5oCRsRPxifGbLE34pPCy91NO7dYl+xFk8WWRt7KyglzsEXTw5LKKqMP/otysKJ
ewOnR5bbcYHFc7rnUFdIlyEdPnajmzHZrF2qICz/NiplnPwDE2UR2EmEl7VViyE49CbiwE6U+N2W
lNQQWU9BPCoNaEPgbqluFcC+ORIxyF7rQyT8GM0fZnFnwR87Yo5ogC5GlCWuiYuf9Th1BFEdBpGf
3isfhD3ahOYQJGLbk544+zt0RxqTev6AyKS80fujAP13ylxjMGx4YJ+2Sxo0U4J3Si6KMs6JYPn/
Br7JNr7lCPH20S6LAInv5TWJyfEPzSQVzC4twtK8S6awGiEpohmG7Cis5Ctg1x9iIsOwANc3+B1e
gdRwua0hbFxPQGUzZ8ItnIbRBUvCxaceKw6UsRPuA25B5JYUkq+r7QnH4MwpkRVNyK1Cb6WhD36L
cutvOaUAsaAWBKj+MgEGnReertn42q5IBLPA0TpCefL6izMWcCi+jQue5oOWmPtm0tsBXOm8RMWa
2ZbEYS17SY7oOFD8s+rkQZdxsdX1SRXN0qpl2UjhHpT0xPXbd2CS4gkhRUeYUSsnhK4aS0d/rlYa
I1iWobez7pRtiFQAnaG2j/fm+DGBc6/YiD7oipsdUBsqoqOCmjoUFbqbSbELLN0BDZcJzYb6I8Uu
w6mgAEl+1Ao2RdhiBCGHLhNrqXIoHSKiG8pSjmYvDPYH5b6XB5CX36qPBqICZ0AHzaCMCmKRfnxm
r9pGkmo5wsWhwvtsnoCH4lvPMXVtnZKSZs+csSXruTj/NYYttgFt9ZPNPhNPVHiY4k4oeY2KeDnY
UgFp4Fycg7trNodnmKq+KZMkRpwc9O/1I1EWDZ2YHg128Wgq9ilJfsDu3SY/hU2exM8PszhZlNMI
M2XPNexHTKJCpbz5y+GMubu4D0QGVFxyOim0bYs7FPa1p0jhMwG/zcRU4kdM+Euf20aVkugX/ypX
wa1HWkz7DAKT2jF1WgOb+5zuMz0ptjdNummaZrnyyCz3Rv7vhsS9Lnb1PMF8TOFwhHt+bgohsjb/
XY8hWcCOfnQ+85NWyvmSEh6Nqh+MxwWoeE3HJ/J6QkepbC2mNaH+mJ7p2/TtZ1l7vCcYCOSPm7jO
vLxE+l3pCIb6Q9W7T7nM7tgMJGMlxbFOKc+quAx3IGI9Vjk2O0ibong5WgRWpeFa8r1Ri19KxFIj
UttHVopJ1aR37Xe5KrIzw2zqavsWBfy5iKQVu+v5XGEa5fAOaxK0R00y0X4KrSdjvv//M956h4C7
8wJeEAxWv/EjZardRtXn0DBpw+g7vxJCrDhy2SBrFDaL6o7NeLRqs076dgz4bZ7p+jHBW5y7/RoF
wi7tUp52yOotWmFkAgIDJco+n0D9xqH3FPLeRHqog/dc+O5GNBs07V4ne+U5bKCDu9Vqo/E7g8Jp
siZDKLnMWNl7S30WxMD7cyBb3PZjrY9YeVtYxWhAcjEmbtg/TNnJ0rDEoyDsqr9ASDz3hFgYp2EX
G+NGxrxEgke4JFo5rT6IomswMq87DbdeXtJda47yJ3USNNxaxiz1MVTRuUYucv/h7Ymhv3N4azVs
TspjmrU5hiBYtc7X+irKFbl12OZmM6MmL7GoKtxMxWllKUAB1/AWvnwwhFE3wDxlQHxp+JMewKj/
AVFguhuL0HN/43f7X5vT9nniiVTruqBCx9MO36E8toGNrslrPGplHtMUoIf0Yg5ykGQQhIo0rCK+
eRik+lzIYMjNlSrYQhFcc0Pua7+gQz2hG1IOcqfFtZ4G0X241htcJV0omHsv6y3NntJc7l1mpdYI
tm+Hy/ZjDyNicoQ3JrrDg7xEhQvj8bbDfeGs614XfmQn/0i+fBhqK9m9JlutzF/fnHAD0kokAu1I
BsGi172jqUNdxIkocKdUZr4WysP9a6vIXC2rOgS2byP6LOrMcXFysZAuXCkw0UKCS6mhXn9hP7fg
aHtIq+TUaMtiUFpMfXz2Y2oOT0/nGTYBmn7vnN3wzCykV7exh1UgB+PSpinwx6bSFYnAe6sp+sHp
vbwUHpwTDlnKt4xA3gNXwIym42DGNrVrSSy3FFMYYw4G+BFX5Z4sMiL4kdqL3mvTFxmhcTpRxR4C
Nn0Igv8gxu6dbybj0Cq5eGUk8ffOoZiGRNMl7loWAZBrge/MbFXafxLqthGEkv6CmWdpys3kZaJd
g6mnc0JZ8qGgpq78JIxjXb0MzK+bzxKgLih/4Ol8WZ2wcQ1rla8jq9w5hea/TCg2h63rZL5c0e1U
7F01tH3xF0dU3ghP9U+c853dCWvqGOk0EKbk6O8LKnEVP72Yu3n9HqzMphXt+3zTopLmc5AtI9va
+UwKwRBb9YmUSV3wK1PNIZ0QAzV0vYUjakcs6fn1n9ZsBjRH8nssZnRB7Xf5+xMBe7HcF9QO7cRW
RD/bs109W9yGNHDxz7PN8RokwQS4JtQssxkc8Lkynh70KtfsY059ScjHoJ5PFpe1In5nvqYL30Hv
yPo94cn0VXgguc/r2SWhx2LmosuuOIywpl6/8ImSujlGzg6ucZQU9PJSIvIbv9Q+4Iu1P9DWHm4F
PSuy9qh3b6vVYzAv5tDfLhv1/eNckgLYiaVGtiTtaucTbUni8bNSVjcbVs/Q/CncO1slKLAvCup4
RmweGEzg8gyXHwkcfYysztGwB6KTqdx67vLbP7/PcxU0xpp1ka+RcctEINTPOLPG79yLSucsusmo
hNrpBpy2AlG5muwczQMd42OAWt17tRi6Y5M4p6PWHIQRcmtswANY5eUDxGJwWdy34Ea2qH1LNIXk
pwAVi9U/CXlR88WabLNbMklHQOW+SCHqhPZqn0FeQS/zY5Wp8qCzDPsgHIupg8/MdyIAnSANwDI2
tLi+TQK0nvM6iVQbE6C+O2Z4GOnU/+kL0JYETRfC5k38a25FCJwCXVk5SeOMv2l/4dojFNipuoHI
VQOmx/VmCw5PCMoyN0No+8PG8dl0r8NDEyWCgTxLiYjZ/+npEVTHoduaCULvsqKNFFBBdGLURZDk
jZQcQUbFNKXpeXgEi9eaa5fa4uhXJPw6yGMw6xTlPqA1tp7Sc7wOoDJvmSvQ9w5Fi3PUZrvTCIMY
IMVP7QTBXWkYRrNgtX68LN0zqu1574EZdP6LFoT8+gCVBJvtZeEG5axN2tkc3c68o+5EiPMtDdYu
9wt/UgqL9QAQldSgpPgvIOaOTvxrMVPfyhMWAO4lnCYFwYdSBYN3z81gSI7lSMlLQ+jRATVvJPlZ
GgkDoDrrcX1SjGQZOr4EowToq6qlpjtDMukeGC1ow4mWd1v5jFioltY3G9gHQ6bNKA4cAFC/FRhl
xKOoPUrZXtUiSKsnmU5674/ehXFvw2N1Ll26Vr5+qIQ/8QW8d+4/Rtx7hmkGpkYmDqkh5KOPsbFG
3Z61g8arzeeH9xPw6bEGeVLNW22fB+/rSXjFEzmz+K5LKijZzx/RTxGOF0+XPmLmtuFsN+cEsFHo
7as75i1S3ksWzDWxrSQVsO7W7aIvPuRAn4XxsbOWrskqARbf4xU4+v/yqM/vIDXY4M+hlNplzpqW
aUrtJI7958Hhz8jF8eyae9NaqdPbDBuGNHrJalACITKg19C9UUZ7Qij+hOo06cIlTxvrZ8WH0h51
qCK9C+js82GDdKgfz1yWuXjlQRfsfE53XXoXnMF6/RXMXPHz1koGaVC5tzucQ+XTXreGD6iZ+X5m
2HvI0GZ7jXSw/TJwyliUc11LZ2hzfuvRK8znOpDKg1yIlT00QRGONU5RLqfVvjHXruu+2qmyL5q0
5FfygwPt39kSHhQwi6SgXliQe+HFWmtNwpgUlSIFBIoByCf/2hnkxqolns3P9i1hQoStTST7Gy7e
9t+2m2O4Rhe29bCx/h/cZmDq6S+yjAHP9MvSSdIFAUg+AkBIRDPeocsncs6i/Dkq7xc+gENq4Cp2
yz4inUgAW9wt04TEcnia7VhTlD1EOd98FEFW6yzE1VNJwu8C9ePKcuL4Z9/g12dWKs1fALfNbGRW
1Vko6RKCIS+7Wqy7H+sya0mj7jqsqp7QAK1gJ/PLp7hWPHwwvuzqGEuskaB42ECcbk+qMpndEhrL
GihhdvsRpLg4dJxPoZ5TH2x0JiiRusGH896G9CEwmwf9fo8Od54PGKxHMBtFWJM9jmLOM/oKkuTw
lHP5pogWYMi+X/kU4i+arVkNNRwi9G+zBb6h8Kyk8oVZg914q3x1A0J3GqhNZ6KkzQxg67iP3cVt
QnINTo3CDnWHFg8sfTk/DEvvz7N0NQowVKd5wf8/I58Wr55J8UEDTJR2lfqNS+KXWZM06Vj7AbwP
6z8jYa2wnv2WKHhwY0vEMGAs/gFCQZ7RYjiKaXJeNQTd74Oi+e5gdmsikEik96/JCS0fXcX/CMeH
EbQsOYW+gF9VKq4A69B84U6KjWwW3aiQu+k2CRX0MVy2dxS2q45uRleyaLhd6lEnplxyM0KGH2YB
P3VrbVlc4tkzScRccdGL8xrJ8axiOG465koQs5oxqo+hPJ05NU64zKAHlS2usEt3dC/Pye5aiRnl
6NOBipAVHKIOjFQp4QVXHJs5TRBktyjatN9yX4bDrZ7nQ3wxNVyJbKudM5LYC8M4tahuNNlp9AAJ
JMZ+y9ZgP1tIvEilttyFBrwfZytw6H0lA0x3FqvApDmMjCahkNNyB7LKqxhUuPvwNr7SzKCDjUfZ
WWbGHNyflfEKa9dKhepgSuHHX1eVP2j8m8bEUUieTjRhj5LA+XMhh4EJyDkze7E22lA8JmHoatVZ
V0+NJW0QETgHn7EGQXFuXRnooqBOH3ZzPubSPunXGs9Cekgw5FUmsFAFoDyg5yW5fRIkOjLosABi
BOGEK9TgRsifwrWlnppJknprCxCJ7pC9oVbh3gCqykuBj66wXSrDRyyyIeTisqB5M5tQ3SpN2Zjg
EVtg4Ubu3gjDGd8orB9xuA3YdkV721F8izdjleGp3X7xegYSc5RysZah+jeC95LeYLR72C2K9Dog
wqKkZSbtpLecvwHNrx8D/69afPR7Wdr74Qt9xhn7OPizhHd3aKo6SXq4Y4la4p0qRWm8E/zp4y5b
n41DS++Id6CnKj/asO0ii+EdiulkEgHOWt+phwLniOqb9vxC+C/ydmkRe9OHWC/ChcnoZziZHFwK
hx+f+pbRkszLxzS5+Wt80IqUelxTvgLJNl1jdIaZi1hfI6Ri37S/JE1b35crq/Dy04aRCDpBK1in
Ax9nhOelS3oar7TVuV/uShd+OSQWL5H7kimo5cceZmXRGfTDXf1CIeE6VmxmMIu+hZHdxiJBf4Bt
Caz7vqM5C510DlU3rtxzZnpKzOBHSFsrhCELd5gjyhTFOKcYo88VqUwoHJa88tgqgtj79NxTzNcc
Lxqvsx9BE3fp8+XlEjvtBPlp0H5evip/1dbuIeZH+2dNzMeWvbzb3hA0x7eWipGiGocwNHAkp7kt
Gi5P+1pq4YqUXzpADLuhZh5In/lAPEw8y94DXhPH5Nc5VnJqvDws2x+dx3mo8ohkubla6mLQMs5o
kh60YztkFY4gDP6XPmr6lJu4TFnyu8IZwk3LtnRFIXtLkcsiJHKamxBHYTMBPVKoDFEgJ3Hz/YfE
cVsdewAykokIocqfQ9v4b7+CmNOst8bDC3i/5PatvCRUrAtW+B0DN2FrJK10+VNHFBJwwy3BEBHA
0ehFq+imaNX0/JFlQOzwm2xWcnlInBRG9xPsNqKzvyUO6v0pYQfZyJxlYitgHCOmOC77sFHMDC4i
0Y77zOCu1ncwargEC9EcA8N8iW/1pJj2EOaeKlu0ng6ATSToNBosoD8TWKHCnqPio6rGazCpUNS7
oGW6Dp3raR6EB4vbnuvV7pMutAWYrTZaTLAczJwT7WAVEQ1HyIooittYkKPut2Ly5hVikXqAF0fw
O93wjRWGfSzq1ztLkeETIp5fyxrjJxYCRzu9g9XypISyrwGShjpM7jbfdyBbs6mRJSXpN9Dq/Y1v
K5x1fjetAbO+JHuFPy0PJwzZKtZeQPc3I892rFUdOEuxNb9bnh2E+Y+0kEEtFcKsVczNTFIftA18
2g7pf1/LDO3BmsyOObGlk+TN7QjKzj+6Q6mTkxaHGPttVUfPu6Jow23pMAKnjbfUKn8XSTxHnPaU
bNFhR11rt9AFg15qwIFQWNhKerY/r3f10N90z1v0txbBzQijPaaByskyQp7GpGmu+LwXcVuw3HpB
Ofz2pDDE+1XgpjCPTHfl63BcFwmAm44NcNFt/ICOLmT6e6dHHkJo9PowgJw513ngGLx+cjun1R25
t92gt7phin/zQ1k/nv7xAhPpeIFWLTgr7uXrZzgyw9F1HmzeHeXfyeg7z3zvPVFLrDgq5kkqaD5c
H5FxV41xY1hEWuBwBRVB7nfk4+dVWs1CMx3ac7ZGhcyMlFVX7yikU2DMOjByxZVP9e0OyYTXgNkp
wYaQ5xLWBFNhVj0WtO7lMXW5SrixGsOjDSgWW8k30KzfIiVFSQKvvgyE1A8BmwcQhrygoaTlr9HA
WpqgilWmc26G2NTzqy8wlPM/ghHx0YbFzRldxQzzZNAc8JaIVvchgCwo0tmK5u9AfiTEExuqZr6+
dJ5gstbRprN+KxTxo+5mCOpcXkJbU6ixig1JHAC8VobyxlQcw52L/wCpDeGg5p01x8L+G2q+SPrH
XsXlGAcaHz4MTWVJVgPlPATbLquylu9S7LaFveGK6RZHFNFZEoNNkYjnkxzVTrRz5D99GKMJc1an
g5Q1BLaAZ3NUgk/1ZBrCe4CEC2vDMqYau+Ghu/vBCO3zYtvXxWOXxPfm10G2JiAdsW8IsHwfPeP5
Oz0sA/J3GWEHGxMn6lJHzwS8fSmvOQkpwnnMlAlczaDvi3VQE1TUzNFSTVsLOOXLqMS1zUZ9lEOn
ParAbY+LYHhGenjEim1JADKfCkj7KIlhf3VtyxbLWdkBhfJKS++tHbOUD8+55msUYqLgCsovf33T
p9uvRHSE73DQgsCJsc1CJpSGjzHRvfqRbsPE/XaY4miGTFE9kmPtv6FdJ4hlRAVwEiVDSFt8Hib4
iyjl5ccZ9B289/BII+RbrNesSnEq9p3GkqHLwR9lAzjaokwlG0A2j/zB3/Xb4RQy9cQUiPl8clN3
+SJwhDpJdPFbTp7sOtPILcRH2o0n4mCxjJoLRV0Fyj6GdEqWEzdVGr2tDzz06L05+lC10Y//jWCc
Ww6RBeEk3WPLRS9Lcy6P6gLx0yT3ViuxgtMLkl5EqtwRDmX8j+t23vytaNUPbi9xLGI10UPJVgtv
mqUsMcZTXh6XN719VOHO/pbkZE35I4SrehejBUBL/JAM4hAooqL/LtF4hohyLmU7UdAe/Ycn2Lcj
OGAu6J31gVLWH8MSm9zGgOHWEo747RWBFVH2j6jCrsaxNvZQ4oqARzf/ewQajFRIKFp9frZtf0sZ
0d4ZU0sbRSsKhvpKWZt+NkNclvH7bNUBnUxwoZCKwWs5WNRzguBb5njxDwupwQQ/Nk+PXbA2e5GA
sfsNnKoynoT0W7o4ipFrP2gWUE3LjMEvs4XRtW/z1NXWN/GGgxu8+cf7w7axfjvByfIpVxGxFleR
NW6GnDLCAyc/jZ3IgD5ot5zQFh5gQmqP/xBFYIUE1amhepKYwe6ZPloLQp/LCzUDpt0uY9Tr649E
rzUx/i8fSKiLVulI9t15Sn7wCLfsn4fcCjWSru1nOTZUBGXRqjrU55tiJawkDDD2qpcT6lm2s0O3
JZT99PvKrZEw0ty3Y2ed5dlNkUlAYSVxp/u7sYmyhAKDQHCjkaprHcRIntlhWkMHkXSeiT5qMEb5
X6KO+I0oew0wro03geZM+GtcMY1jlnen199G5+Dj3cBFTA/4hWNZlAdtqBxM9Go4RX/neq56z0r0
xVjT/xNMxTr0SeFGnAplESPI22YSjnm5C9Ne7oEO2aWt/ZYYV7NaXRpa2qmYPChLTKwwiNgRpPM0
884gP0pa8mCV7+/kUzlh++LNyfik4rfVJWvmPOhCKBvaSxiLKBfxmgD3VRsKnzcQ3+nDcLpqICpg
SgeAweICVX/j+GOEp6EO9isV3JfhOGor3eiRC71pPtsQKM7+oB7OaiFeCdPgNcndaUlc0pRhnLT/
fvpOGhl4SUDnUu9rus25R8wRfqfTmglG5PNBZ0qmU6r0wJeGNSsAzqN5BIjnwx+6WHsEIVWL9lQw
bTsv2LQWQrWBB6bHBSF0hdpsx7whJ0md9Gq6d3tOBXgr3Out7xqJFUiFk8Xffw0sDDxbGG375pdP
qmVVfUqllwt1mgcx0Kbmly2XoBOHqXendjLBiAe+xdmIsAm1WDPkIOpJXWq/N0bfrXlaUW7D+K9g
OA5dUK89j3srA4ZtiT0T7o0cYdGPrGGNJfKvoQtTHLHp+PZV8lGkBs3d9AOnX9cwc3pbxy7kHg2y
4Nk5Y8v5MQ7SIOU5oao75wG/i2hiWSU99p2F0cnkwL5r41id8p1dKKr72NCBKXYQ5KlUZ6Kdp1ON
9zcCxqqk7DAySkcczxmxcetxh0TsnvGWZVQwqnv02rwF9LplWQ2+Vj390yW7aEoh0WLpLz10lLbk
PawM4MLvu4bRQ3VtUfztdnb0ZlTMrZpekLJ5oZIim+32z0VgixrbPyLPbSqetogKy/2FrdqVEd6G
+7tSECmuB/GUE/n6/fKAPWHha3vSiDs+5gpVskGIWS19lwq0qOuygIGhMKif6rK3alrx/v9veACF
NrFoC+6j21ZtXBBS4QpFPpx0XdIND74uvjVt8fw6GgKI/YuU5Gy04qeSPrXEOLj7cn0BUPx6FPVY
+zpVmC6r55Bv7fwZ/JLW+3Rhxv7oTLrNpQ+vJZ/XZw8XZEqFtlS+myFapiTkR8mP9vPjvrLSDAm3
9pjK3Y4p/0OE2FNa/O3vIHVZocLXUWDsVOnqbhjgoHzWsS6H+ajZmk1h1ku9wyQp1h9MusRWmI4d
IABfn8gP8Ux0smrvomMidacmThsMFIxin0ImQqTlxVBzbGepez6W+AqFnvIbgPdEqch3c8LgxKMR
7N0NpvqPo+NHD8UQZMlWOLfi/4gpLsveFBw3IrNLhma573TDeH/MAH7JJRrM/8PebRiewdcpvQv9
XoWYEhUrFGB7K5Fdl84tIaTlj+D1bmkGlO2/DwW0X4gUlEqGlylg5BHaTuAKGmAw91BGMerfIgrH
sf+cB1sMRPNOtb8dnX+3OVABq6Fc3zf5Axg5Lvzflp1kpKPgourVsmxEdTHRaYl3rt35GOuXQSZx
1zqCQt5DPdT0ZDPe/AQYeRLF61AMPtySC6xGsTEir2/y+YYLSmg6PcWGS0Yo3BISVdCDUxfILdYr
Uq5VydSpN3aavahskH2OqLPZFrniNFZ5+X2yUz9Kh1zEzttNW5dqePWPYkEg2I+jS4R1icTBRgXq
Ip/WtT/TUPbdRNW1I40m1fY6U43ebS/H03wVxCfnZmtJlSpwSDGAwqE0ad6SX6WtRaVVQMfxADgv
nzmSLkSiX+11bgPZRYGdTreSQXqjnFoIKTKREM5mhYUdd7mNNCVWnDda3D2umfBjderVCQZ+x5Ly
+BKPCUMeBIS5JOzke/kBoDsH5D9yZB5kp2VHe2HccJWDN9v8EroGeMpdVwU/9KSqrYxrhFiGBRBN
dXiAIajJrTIa1AYBWS22qBYNulvBstsUERu8xW2L1YJZDuNb/+qUpQ9TluqyazNhUU9GyoicfCBp
LtLXDnmX2vlCY3W9Xb742wXB63lP0997SujiiQkNLA04oSfV6f8IRQqZDplvGe1UAgUu0Mw4qPsB
rjxr+169TEHCgP2a/LKVhCoh54sHnDwLM1aUTQ/6WypCpY0GZLXXgT9yfTlTylNfZGhG/Mxe567l
kLKga+yyBZv4LwqWh9lAB5GnZP38I1Rp9VbWM/dyEM4xOrgpFb6TrQcfmU2UYxM47G7igCqXat6p
tQ0wgBwAdsXAvJnq/K06N8JDBJt9Lz5Ef1bCRzSoRlACWQnhy7AKR/y6hrvSro1+a8td8zR5nnDX
pZvP3wEitpMAn35mWmrr2wmmRG7jtAioVOkX5SAke+oWMngw0lBvsSPpmcwADjEMxukAW58LnyyY
ryb4OsK7JP9ZzYG0HADY+oTtjY9tAVYfgD0VQ00kSPG/Gy7UqGC22gCWtuStI2bIB9cddjRXiWtB
SNpEj3in58JNOR5Iy2DyknsCo7+mOtDP7vsKVdAAEHKWjXI7LlB5cMNmVqyY2rpMm5iEn5IkhOSw
Nq+nkzrpCcCMsCzg45d6Wj6BeBlpTQKA0A0EZXKZt2Sosbww7yxMWQJxH9iafpghcz8tRdGUksD4
X5sOrBBNtVYH/PHV9SXA+1B7SXXikhnrpkq/Cy6VonZ2i36WhmK2kKGmBtxX7QJLb+ldv+8Xq7Hl
SaCCveim/OM/j3Z/TDbuRDfxprxdzNAD3PvBQwgVucbZeWUgnI4+vXRTLIBKZH3hBIYicYxG14oR
817/82M29AEKLopoBnEn2oCdo6QvE/3XdSPr3pUTiB1D0GH5+i8R+SI5+x8VROa7bPVqOGUfrEa5
mycAp8WFOm+tk4fDcphCTlXvPYUvIqrD4jFbgH+Ra4HL+cKsK1xq2m4hy0HjdLSMeHy8fpuaYwwd
J2O37tbw3lFXglwRi06DITaMYi8XL1xbOXxwjxlQPav2zGpGveFvHbMn51sq8+LSckKt/GLourc9
fHB2g4YORqD8UXayKvR91tu8RBIh2bYepTWigVT2+oWvPTi4uKiWx57yh02TN6flfjpmY5u2EQa8
qtL5ka+3/9A33LD44P42pE85rC4jEvGlrKh6l7DAN6k0Z/JZehPfDmNmt5XivAFcjOsstWQxnHnR
RwXDQ9SEiK5W89ucAzVuy5o0DiXIbV6TVBmRD/oirg/FrlFzlI26Ds3S4v9wxEKgZXjUUfvyDxGQ
hl6L4LP7d3uBLcXjEKyir7fzvPIIiBHfuh/SomLSCID/hA89wGEKRFnAuoLiJUqN/AsIJnbN74Ne
HI77y6X/X0KSxPeAXihbl+FjvIk+NseXsX+cwoCc/rJnazIa67OQRErhNh0YinqQ+iInJci7wV1Y
kVwiKuPpGb8e7RC+dbhK4nbQDD3pF+6M0kOBb2fcLcD2DIAPNf4ZoTlAb8Ciq40aN6g4bvnS2TgY
WGyVbZ0YO2dsSJKkICxB8OoxLvd9XN2GzLXsgBs9f1V4CcxuYp4t/63MhBTXyWYFquXvHl+sfFd5
vKZCDldd6rAirPAijxOZ4vso0a4mGZt5Aw6QdFCpF+AjRT3Jssdi107/RD3jnUIUe6+nVqOycSkj
JS0/lpq1r5hD1aViAmKllHDVPHb0D/Zkm3MOQVE6IJ7JN9BgYGgOnnPwd7aF8PC8VubnzqylRTEF
8+1aEe8O1904OBCPXXelvFrUE5X8nWSBjECfA2drzWzVK4FS6t3oa5WKGPzKLS61fR0E25FHlvj6
1ug6HdQy/KmitMkXTql8R9zDNgdNKtbGzOW24IHKmp6KaPgL9UKLSlhzAmz/8PExd7zK6Qky0g88
7aJij3btv0UVLhuz8+IlVsbWgiPJuJcnA5SCLErTsGZjSJGZmkjbJqA4K8zsEj7Bz1Cw7rd6p5B8
akpSe/LkM93N8To4E9qSTLYBG8itFyurLLWX04RMTZjBUOD2JZ6fMMS2AkV0duOWjEhVirrQXrtY
Pr+IRj5/rUHcIkk9rnl0BGOC5U23J1hXfu/CgbqWQjRaUx72BN0an993q3bsTB9ow0B5UuxZuOeL
8jh+Gafaj4FyXd6q3TCj7lF/s1cv4hqnUXFoXJUAOIOyzqxwRXxsaYGca/l8nY2P8WwcIy7bLOBo
kCh6M0GAMw7ZhqyDPl6jOE0HdNqjmccPGV06JnJWu/TlX/+PXFC1YnQKWDTnQ6yniX4uKpNkE/K/
41US0jNMYdV8SMn+0/NSZQCq09URgMkw9L3QLTi+qC1wni4ZfKMOa3JiplroYzk4Vn24KVRY05Pu
nP22FgDXnBJVZ5ZBAfVcS1+xIf0Ne/G8dPUEG6PmQP7F10iev67YQuK4HrnVohoV4doj0IKLIm/Z
IbnYKQVvY4o0E/VZT4nUhAVJuhjjQ4gvz5AsGAlwOqDpyIGoGUOUUhhZz/rixCujVVQtjfwOWVaY
ZZ67AxlxeYVnRTrbA399myrLMJ3S9aBPQIHcRWeJcPtRcUZKZdDd/IL/l//AbqplOibrDye+6sVH
MRxH4HMfd/pMglK4HlL7Hpztw8+lCVhMF+Py5kowROje0OhWOxOSU9I2BghuHr/e1ozJPqD/k8wa
4i59GpKsItJZ8Xw29tTY0xVnYxU6LTvWIV/+qHu30k8uOqJnhHltA558Fjtd08t7+hdZzeDLVXoF
as0RzK2MmvRRR3pctI9LGbrKnQjnSCj9GkhYyziockbCkMSGEodzmu7fTjrj0nbGvDjtm/80nbFM
D4xnwEl+EHUO3g5zQJCdPDyoCdjhxY7dVMD7omJFGQCA1Vx7zH807tb2fKZ6mbhc8J0imtZqAdUP
Xcrl+jawRHwvY60QTlEKwOourJBStuBbuuwFIZNQIm0eYBjvui5o5HR/fRM0Un7ef/ffSKe/xDx2
prgeK5mBDlGDeWMUHYYy9NwMLdxOANlCWBD3TP8zrY32F4eufep0PwYX6bw7Nw/1q8fSIeVl4LNj
dFN7qSTkGI8W3IWVvzWzow+Lbi5zfIJ5W1ClNPhUvbK5KMF5FsITubJgd0Va/JvPB/uJYlBLi5ln
PFVvUFhtvSRfhHNmknGGtYiKM562W4e0cl4K4XjztQX2g1XmK7HR+nvUYhdLwqiGAoMhESuBDKx7
TXQMAWK9Hpt5M+SsnafwDy31zrB7Z7wxPNTrS1etFf9t0ADG08NbKY4bcw5b3RPVmMW9xeYhvPro
OOtdGq2FUu0wwwpAH+FbZDiSJjgHOZGKWxBqBSsvnAjygwQYI70BlcNQVYQkhRuI5QnzWndPx/7i
Kdb9KLS0hE7JnNAqpM2lzprxYw5Yb20dcZ45rNn6u+mXf8eT5XediVqhGEEDMvqquaLa2CuGxg7R
6hWZf2JcNKkJxMWwjhoeBlgcTlP/rPK5jQsUXATuTHVCujvTKV5FjSEStw+OYGXaAK1heu5Xtlqn
dlGwW0eSHmwY1TTD/b6s9Rg9lMbYFsAHm5MS/1d63lvERQgNsYOqtEb2rtvulm2JgLvJi10Utg5F
Aw/PlDmpF1mZLEHsq0/RGUYm8xWU2WPdqW25EvdlUkCD0PJU4R1WT9pMqmgB5T5dYCz65GKf5CDu
pnSfhYXrZEJ2QyJFm5bDkVP6YZSpsI4NU9JtP/8UHMQYxx+tjwdiwVjkAU48XJNwHQBEQdreWhce
tJdp9Qka+PmPXSgYwUpMgaglJnJFHOl6YhNqBw4vjCw8MD1nmTTK3XxTG00xbk1tg15q2Yh90Uv0
hKkq4/yV8iCaQfsuJEdJMxFoGx6sAVZiOinFUEsfIoX8sHnm/r/q7JaJnWyNEjlKAPVqFBGlcK/z
Im47Aa681Wqfw3zwafeqan9VnUXztF0Cf8+evgbACr0QeFv4GhZko+BpZe38eM58DH7w6rgDlALZ
WZ/PbF8sHKQxsFzBlMKCI8cvARBXeh6h5CxvZJRbJDm8JlfpYxyO5939QydVcyi12HdftjCWJh3K
QzSBT42Xw40eANIhKNp4C0UGhXOeO6mDuBWeJrIMoOKRKjmSS9hghn8TvVGBOmjKe4bozhLWwwBv
cD8ulD6fBhEp8/9V8hY+PAKTES/ZdUB1NhI2w+Gp/Tfl76/WhUJ0v/0x7wYYs4BR4BcvR4jWwZbS
vD2yn9pgh+4y/j0SbiboVisBqjHyvKESEHF2IVTIhPnCXPIicBZC4PnKmygZwT/bdy2hrztTEgQG
szMl2eWorazCX4UDYw2YzPmSGc3/U2uZiqRgvTF7bgb8rZMtvLV2RrUPTk+NO0kOfklTpNTKzzhR
xvfgcP4z/CCmLJ+yA9h+t/9OetBUJDDCrHGjXLto4+B+h3WjoTMmngxepO3cVlHxhY4rpum9/CK/
LRMuodgc+TWGSGzsNFBl/z+j1bWWiwLwPPptCK+oudej6h9OqLLK09WLEBLe/XgFWBHOeryg22m/
wZ6lJT6Lo+9LDyOoDclJV0GaLPNhadWdZ5sppAwUGrzaPC31hqipEzMIc8fk2UYZqSPI1vEaAvv8
vfZ8ix1+yp2f2zzm7nd8uWyvLvtomGb0qMCWO3tfbDP/dyGVm9eaydaUG7Y7X+dp8sHJjjS/c7J4
ifEDv4Izwg/wPHod8EIhLbTOLJJ9tVaPHHA9pGhAEOYdUezEDD3bu/ScgRYZvojhaUSpUSt2upJD
gxwjId1QF2V7eT23Bm1NHnjiw9DWXD/PHuHX4Yai/YqJbdD3uio7MtUt/rNvN85cX7HiDJWo6YTh
s+oypRzD9eErVfgwHvsGxMQTRw1rd4KwR5vWZcOmaDbjQv4G6fogC8DTTr0H+KmWC+T1VSNvImQP
hl8DC8B1XI3A19/hMwcS8lSL4DhbJy8s+ry3okztuqyHIAl/PyygLTMThHplukb2o1N+zYVkCewt
Ib7XoJEZxgc9A9mZ4ku7f7WWPrcznxTW44E83giS311Hm7hF3fSIaqT/2GbknpmCQhezhTcwfRyz
LnC+v/q+d0bwUKUgDJOjakRjVEgkW5GDC5d8FbxyGG0Yc/gnISQq7OsEM6AxMyB7ur7ftyBp5unq
5evUaPBEz7ERu21U+3bxBfqyrkKyMG47cjhsn2jBlJAQn1Q0JSSYuKLN6EIul9Fz1rO9tAe9GfPP
3oHx1IHmcko8V7fb3Pz/3WF/kHrGN5Nem/ldNGbvN7EfAsHhPgVnR1dEEMsdiSkgA0rnfv+n2JYY
/DaKIQEcLiTFH0eRdBYd9RZr3qOkBNLI1BMSbv9fmskSaf+xAKXCV+G3Ru5ZpQ31kGm8aWbPK6Yy
SEww3UkzBJXslA3OExxDejkdFTT1eWfc+7SJo1fxwQQg+QOtSrndqmM4Rt5YwXDsOTJcD1vwUreF
fIS2zsHIrZr4f1ftf3e+4NkqkyWjk9hADPnMUeOGA+N8bqJm7zrp1r2HjkZ8FwfXq1VJ6BnnpQKv
yNfjDBPe/ahID8/RpIwMVsUaXwt+/+TH+Oi8hYIZQ+a0HGQIiPax/fcd+zf1gDV7ejSKkwlElZN8
iH5VfTmukfGC+ajCFqAfJYDmcUwpbN7BvuNKR9XoUa391pjvjaxI6OR6eJnKtZYxGZ9mwHDDlMio
e5kjm6i+SHSTVS+StKVF0GKfeLggP23wCdzpx6gSAdDEb772qFEfQqRiwfufDL+a6PabQnjUTssy
vDlEiOyDJLzUAzMbg8YY1kcm+azEEWQR1vhQQtJO0GSBtQt4IbWqvkOTRxOiUkDKjiXwlo3ybhzs
blryMaR4AaM+W4yROzzupsraJdeugGsJ0bCkXDuhgXhwSHkDRWOWrYODYyt+hqbVjX+y60Qz/jnW
rVRKLBrHzWAqbj/jDgIOHFknDT+0cqSJGYCwnumUz94IJ/Rc7WhTc3KFMlyWTvu0tNbdUm/p0Szi
dsswpaP5lErAM+arP4p+TAak8SQRiAeAPoPq41wb3oOGIYyrFyShY7HoZxvUVzbJ6BHRrM9UaUP7
jBgX+kpW5eJSNGXCgKZHEW3mDMHsQBXPraMDPjrIZp67oeavxcezIbuM37uJHxxjiAuEO+oYirKG
s6Ny7G3u/ujf0c/GY1smzH9bAcREP3qFHWlfojQDjIkq0uuViziM+PjcOb2OYM0u/8UdTqVLB3O2
6Ez2NSxpOdjx0vt+JIpY0nPkENE6dWoX7v+qgoSOQAQ+ism71ezozW9e1whTQt+wKkbmWVql5IDX
16XDYBYJ+mxvB8e9gwmjM8qxCEYllLYknQrMkvNnhIBdbrpJeobvaQ34qae6hE9AAif2TIkkzFR5
eow+5tClrfodOJfj4SzcLqbcTA/hBQh+UWYZaKu2JDU/4icND9LqtUFYNfOZ1jcSB44tQyCFQ0xb
sYRg31o4cMusFL2TteUL3OinUk+nbKoKFnUQAMfiMZmOf0R2+lLIrUuhNZSQgMslW5iBEEQ3dsgA
shdnzSoA4RO9gsn9s2aNR/hyRr3HsOdXqk66ZxcSIY7HOM5i2uPf5SbfAHzfjWJZ+7YQvvN+Zp7/
nw/nR8gtmNrFMuNohhhnybyP0rNa/4E8WmU9cfxWjWgDy6BGMoX2POAm6T4P+TdXcxDLAdAg/68U
o2+iZwpZHvWHrSFPhAAi5Fvve9ZTBbu7/8i1oQYcLvUBCHqiboWpsinuMNDlbijQX0Qpbq13buKi
igw9vpfGQKnUbaH0ScAIKoQxMvhXRkCM+MxbFTj+lHycnDnPkvBlhyjfemUnk57KLhs/G+7ZRhOW
AHnnZCB9LoX5a12CgBed3xFRSwwT+xaUiLfsAplkxNS/rM1UNmqFGnkFoDuTj4qLswR+hGYPuypd
HMgXInXlKmn28jvcByvGwXQMmUvrsNgXUYNO7eDi2omA+wC+ORN7jhZTgJVsRDlNyEojtEoPjkgw
4c1osFr8fhfbw/8RYIBcXkiFHpoHLYxy2/iVacu4wBKe/FMHqtkr3YF+4NuDlmP8465VUWOwf8kD
jYodSWOYQq+R4ciWosKonozzrMkH0ezwQz1SRfraSPoN26g2g8OyD1BZ8sVlPkT0eAIZCJuoP6B5
sSS1omohPYz2lsJmV2N38rJvtkB9FTN6e7FjvjOyevYxlC/MH7ddZ1vFNgza/NLETHG/dbsVHeMM
2hTeS2uRhrJ2ZLVpW83bl2RKilYJ/x+lo0ZQv2BkPDnHaR5MvL6Ct9P/oExMhc5VkpITfGDRMasU
D4rGvTOP82kWkgLXrL9D/RkyZVP6pJAGxRixXfBkDtq0bTx/lyOKtDg0GYY0rGarODKMYZ1OFpYo
kbiW++iocKWJYhp8JqHSBdkVdHh4W4KU5mF/mOpdO7jmfSg63SYb3ssJGqNtvP2g0n6Gbgp4BPly
Mw/HAV1cljOmDZMBQrZGp6b/U+MPEfoj4F0YpijEO2MXWBdaqA0mgHoTp4q0W9PtNeVj91WAISE8
RQmcaCarossg4oLgEZNY27l0Z0ujYQFjx6AAbDD5JgRuk+WAY8pPfogzjejFX2ZzpYngakAjLs/y
lA0EXFTzqa7jdi3uVOPzN4TpsOXXUuDcenGXR/Q1R0IVtU8lj21vVkbY73sYYXFfjua7cUxH4Al6
z5jMUPLo6HOZBLWCzTwdOZINA9mW+SsGfh1asWWgn6UdXpJfFGesFVgCmNuZ0aoMpmjz9sqbwpvV
1iEv5nRqoz6/XO+O1gTNW97fk7Sn0rAQ1li/fnfCgyXovAIQ9LFKy4i8YOwaRzzXlTddF0USLLYq
taEfNoSF/RKYJ9428W9FUEOcNtmObk4Bc7iocMP5NJl/ijfKfBaQxgaAGiLIVtFXtkCXNgYA4BZu
q5AcWgfvR950xHkZvDw4K7vCJGtXH29Sls95gJqLJSamEVtQC3G+eGNhaiTgIBYkm8alabS7BPtw
IhsSOnqvV09xd+ACBbm06qdwc78JqZ1E1McfXujaO+Y4XxSCwlktl2Wheyn0wrAAs3qZ+AcQM5cY
NWiUs6DebfyURCJCQvMcIGT/IfJbyJcov2eFVzJikajwWSqFsrP4SsKn/b0Xx3+11CIoGodakuid
nPThKWvUhoYAtQCy3Tc8vd+Bj9Bfzgbw+Dgoyo5jkwzQM3sJNwq7FyZRXwiPLmSvVbCwV3ADrlpr
2XiknLjPhhr36GBt2cmVZJILFXEb5loO5QBDNAyWXKynr0tUvwZy7Q3vkYmQvdNMHCogeKV01y8a
okn0wGcgjtRogLpuhRc+j8ZcbKQRmzUOWc/Bi0yIOsEpVopZZ0PxhseyLNPyLy7hO5J2bZhknTbG
el+A3DQVppiJ7nka0VZlugLzxi8dHCnoB/pAXBFFn+WjNkv1tr1uW7lZDx2Fm2TQOmmKAXCaFX70
pGLL6JPwlDQtXGzCLUnz6AfSU/EE46k0Z9zWtQ0EDcX/mmvla9dna5FuJhGrbL3nFtgOuJ6lh+x/
o7Hky7zv3RmVKenRkE/sTU7D5ik1U/EUMde/HgO13f+QFJziN7Qj9oWnHVrRj96ORYtQbHev1o6R
3koO0Rf3+4gD/OxfIwQyrcHCPgSA67KnqSHJ5keFv5FgL/do6ijhLDyN1Wkdwp+vP+C9MFXDNDxN
oSnmlPaK5PhHL1KfYU6k3rBqyrQHppTla0VvciZMI7Jpv6QIjTKK2E97Tn/PZaeIUsLBuTEhZ9TG
C1i7bcPf5JB1EkqtG4Io8elicHkqLlRNYdSLJxFF9cEbCd/NB57mwNSA/1iL/xO+J+rgSdqZWyva
LcWxOOTF8qVUI8+Gf5V47VUIuh+EVGHTjA63Hn+a9jPyELOHZ5spbjoMVhe/Ot5WNB/EZqZBF8zl
uD11VaBVTeD/EJYmsMqUtGERP/Qej4HwckXAtC2OnDK2DE+iSAA0Ml89NwFcwblmgyA1Dvc61See
i5S9dixgwjvKUvt1By/8Dnj9KO2vKuyY6VJHx7+/2PcQXZXkIc5zW7n4cpBu0sApOq0/kekfGIcY
D8s2IYjmG3AMg5N4TRuPDS8DAS1gA2NYVqsgUUWzaySUOSmnWF8JwErum71LLAX7+gFn08XIVChW
bKsOjnZktDRrV/lfrpWvw/q3s85pBR24nkXJbaUlETLmGqMWJgBYNqZmnLJlo1HHtNOZeSrOQk1j
y112vCdOxPRKNJqutn3s6QCaop6zN3dozGw1gVlAuJeDQ3C70kMa6aRRYeJvGXP4GOeIKL3u7JlT
uw9ZjKRgQSbGx2pY1uUB6b1QUbz+tWBrbYGOfhSoBa+fqExnCUccsWsPPjhSMILuOCk4BvD/FhLt
G131exok6P3/n02iYx1eSDduAlZtyjEYC1oNUJzX35UODmQVDrU0eJAAD1K4RNGCJ8/LJ9gpWpW8
oyDTgkuKbiU9JpWkSn+n3P/9IQDa6bQsl4GQsgBFfV4+etNaQNywoKL/vzjtdh7ZfHDNOTvTLsRv
TUQNH92TYrGJS6JjzJNK7wzAMdI4R+zum3YlaoL9OYPirJNgc/RU0kBcV6fesMX+jSlS8Mla9mx2
vJK2Z+wH+nENbmdAS4MfSX6DGpLtM2+I+tERcbPwXoezZrOCHXdKKVJSDPE5P0pcyCInt48eVWcH
0rDGY9h3zNj2yJgMifFYvpKUVp/KLV5dVabU9LFf+N+umxqeT+53FwB5FmQywmfLcqN40lcWDuGy
dekBf7kplDo0na8zXcbYRD2g9RiXPsnfveoayd+rye9hbHv5btNQvEOhf+O9rf1Ybb78HiiOjQhc
FHbJt6M80wPYHPya9+WULd1BKD//NR22W9QTj+HXBNpFkHntj5E6Q0bmbMLPY8GCzp7NKBYowe4/
F8gKAZIrlAgCmiYTjS5PZGmoMS+T29bFE0XVtUwKUkGCqEZ5K8cI6BKB81Ckk5BiqDYfgVyEcTZw
GKWN1i+FTyyhsQRqqLFLrEbCrYy/Xnx7l9tjHrMo5H09DLIkUCPdO8ESUsUBCMWcFf3FqZXOmmJd
4dszap1QE2fxv9wE3p4JA1dvv5ubaH2v3i4YCmzKeZVwlX6u+pwFNocTFH8tRqLXIihFjRKGCNEb
W6f/k0xerTJ3DFM51mTJ8EOBERGMzvliMgjq2vWm37gT4Q+EZivZZmO6erHhYcjYa5kfGqDbgjNj
8MUuwDbcFv8B2Q3iD9R9TCKDtBZtinfprPFtvKsEb06HgC7aJSLTbacgYoC96bq8SU1NqetyWdKd
vLKDqTBM7EoW39pbpDrqJQ41Pkhk3A3NAlldTrFFUINd3cE/D+39mkHW3jwl8yWflNziSh4WKTB3
0r6fm2NpNaVwkIGEN2Flab+PlceCuk5qtNNPm0/QqOIFbnVdCOnU0WXo31CjzvWDU3wuv33qqwWJ
MfbHbYEaSxBg+6o8vUHYY986TgON3oUEOhyMAKOrKYNJRHM3KKLm0IFuAdh8YKGHJxZeHPntikE6
PJo0PnSj4y5YhOciyt8z3w1XoCnWtBVBNMo+Eb6WVYdV26XNRY/RLAtgZVcOHwOf8Ove/9vV7/jH
cOHJeNJHn2+Ek1gZw+wiRI+f+TF5zUkmIajT8OIIi9wBjSNoZ4iD5FzLAp3mv0u4AZxBUgcyJNQd
XFGHtbVY++sTouJXHCbTQ2to29ytpDvoOZv54btrkqTOsvAkMi/UFTh3DEPsjy80VQ3F2HTr/M7E
K3/RlX9H2TEwCvhfMQUNigsWGeu6WCXNoAJ7+Jjl9YodCUToW/rbwBfPqJv8PPkDvu/SIbmZfg+4
H5UiHVIXK5pDede8F38zShBAXAiB6NkxANy1oS5I8yFGTLjENds9uHjF2v1XOj2fXB4OnM6Lphbp
hppBWwyYTjSLw0DpuDFNoGo2jnGSYdUKjnNAbiw+Yq5SM6ifB9UlHrnzp1YUMULg9wkNh0Hn20/A
OczxGxEzr6d36B31khTlwOVzKOPI7tN/cjdsfDeicEUaD/o6/F5n9ijyXj11CJQc79LCoTFvPQPu
TWsfLu0BPSBQyzhReWbPXI5a1Cf0AUKSwxu2FhvbTTsJvJvNpMrH6pvkNBTIl5CmpapqXITebVJu
M8BOatxRa5zkGlW+JADCgiLDttvR8bmTib9S0aYkXB6fCgqX0G4cmlIv0icR7EECBfuxaG0VoORd
g+Cy8LpZToriKTctCaDWjAeJwNnV8LfqX9F3mXtvP/2gcsKJqDoGtNBs31176vt2B+jMldBtatnd
4DBsDs1EFFtr5a9s5lpT3XJgLmnhBSpNVuVZ8qrnAJUJNReUbNOGq3a/knH5fV4C8aiSzB/hGyie
xud0atjWDOzQTA+aDfZG7HM+NVSzxH3fJxVagvTsSH8yEqAIWidw3kqJ7qK+Vhf59ci+4q47HK5j
p0qYRxJdkbruLWbh2vknsz+HY35jXAvorKE7G6z1C7MZH8FlWPUdI1IRtW70KvtPIn728s3OOSAH
KTSl3KXRQRKqmsoc4cJ0BycU8s97iSkiRHkbHNsEcwpeJPOhZU+4WGdmqUm+F6Iq63aZZ2kBeB+5
VFB6wo+j0LOPc6CeOoT1stiIhDDNjPtTfNqua1WmKktgAgk9uBVHslG4a/BbVz42YLVcm3OXc8/Y
6btInPUGP05X2vm1fryHtlJUIeINBYM+iZ0zcdODu+4PfOBi9bdj/T5qL5cMcH7cD+aLqY6K8WWi
cze6hNfzCzZaMTlcH4KiVSnEniRpr5NobSlvVfTmyx6LFBNia1N0OqXxB6io6cAuIZhC9j3y+K/e
oeIf6OQtXO7WRdCiO7UWwsQvqn/jKKPlskvNwoe0PMZTOO8fIb9WMJjQJfirTyYJ0FUi+HZXM9DL
CsVLtnUORffkk3oUkVlX1q/Jj4fDo3sFMU9l2rMAiAoFglJO0zdy/yHQoUzLRdJ+Otxw5IL6A1E4
JHT6f/9OskeFUKx3kPkFcuF2+EWi/c1u9zNrsXFOaxuH6ZkUOn2nB6YY5LkXim5iCU5AZHRsa7rw
3AeU9EIa4RJ1mjdw5PS13RVAzI0N9XHwbCfbN3syF/+4ZAtRwFmz393K/yTlr44hVQG0LHhDriU+
norjGZA3hIAsQ/2yQmGauS2zBOHa+3JORUdh3ajM2EqG5JuncNKWNpJi5da1ueRy5Zep9jAmJKw9
LJQAaupTy/HYY+/fFO8KTQU6CGC6UzKJnVaR9zmE434u4MKWzzORGICM7EAaVl7HoPBiZAhJIGu7
MpBU7FgiNn4P+RmI0ySw7zaalNLFMn+Vm4UcS0yWvlaCFHkNQr1uiSCv3NmLI/BD2WMNxazdjvbd
zedzz6ciDxP+c/P/V0qqLdpDrMxLh6RL6XwiV1vKmmhWpnmrpEBPbraUbnb3+TC6rHjo5gFPZV2V
AbPRjtJ8GOkmtD9po9vunhg7/ttor4xV5fKJcdMyqCLgewPhB26WrE6XWz+pSdrym1ttqJAlIL1a
pLMun1Uyq/R2fhJcoJxJ+tdelJ2y/76miFyjOyL7+4CRkG0P17kXtto8Q+95ktb/7OBfsHEzjyYS
I2u0p8asnKs8hbz5jleKjoFbJntHhOvrstmgCpnTB8na6UHwmt4rIkpZcP6Bb1xj10EqdwFvmgJ0
gT1B5OnbN1f5sUU4Bzmm/fHGCGoeg1ZtYLqqdOhZW9nOThmzu895zPuXBTozjYolu1xHnM37A31z
pOgKeF/8025r/+zPUvd/45J2r0VWA+jxgJaH9bLvAaI+Y8Nm8TAWcD7rfmUeKbMTXl+iuWfHBQyI
PLSxVFYSoOCVUKZZ2o3OcMydx1z8Cr8QEVC8ROr1YNklaKRd8VTVVsSfgxxeeaPBLt7dzV97Uu3b
mPvBeT+bhoAQZbA2eHZG0E4cvbbsGzb7munKVemR/P/NUM11TytEAnRpufRZEZ5yluLOKdwZ32Kp
O5JevBaPD1XqhxAOHXSiOO6G56ZtSuq4NLv0FaykUN+/cMpqzu0EMa7g0L5MbwGwIGfSeNrHE5mJ
Kl0XMybq/SoG9Rd70nDAUH/JTK+gpdWU/qtbnC4NkCHJa1sz5QuGlN/AVtl809u4Buaqwe89YmC6
J/iciB9NCrXQscjroGnqeN6MlxnS+FLB1S87ArQG1KGpbqB60ZxJmG9bChA15CTZ6th4qaP2uQHk
xvolyoeS5xJBupnVNUVW1hxB6zYSHPkooQHjwgfIGyYoyvrLrm1VApm2ybQ/xdtHvDwXP59WcQ1A
WNx3iJkAnIZjNgwMzxLfEnmuH9DiabhhZ/EEbQquMB1AOXh6Ctytk68ykZcWttZhMzSdvIMMzjLl
bv++DoFVmqCU9+jP9lqQAT0jYxuiSiBOeCtSTiw+YC42UX1BstmyH2UGvj7cMCOljjI5fv5MSGE8
tYOvB7vtEAHDTl+MwLH/il0PqWkIZVTxH4424xdBoMN+ppNm/Qv9aGX0bFHV2zjao5WiE7lmbj6X
6+sHH1hNjOrUpuiXwGnvl9pfRKU66ekKeNGbVMx2cruJtdlISGdWaf5TSWcIC8rTLTprMjfq4/uZ
MInrNnKM6Tsms+cdvvLWtvgbwnpz2EVAyJF8dvLco0aqXnWUFrHznoCKlc8mk8ZqBNEf2lMwzjXa
ci7a0cZTKgGmzvCN8SUWXyw2yDC9jxCyvpIXnNsT2JkiydCHnP1lb6s1NaVJpKBRGTjoG/PAlzwC
HRi/4mvrf484sTalPpLrsjDvjl6FvKawQenRznZbHa7aXjJFdNQTjskKnHrp0+pguund/LoeVHvD
6Spvxap7mLRaI/MSfPoINmkcvVwHeSHJSaSDtcFzezhu3DkiiiOyNl2AEiyGg0BbLkULbfyfspgd
v2VvQGPpxoUnb+5sxNEhEObWp276Sr7w6j2L8XX3mL52hyzuZxj1mjRKdOm4++kCwulFCJKUq1EQ
0XyHlpm9HPDn/LF0L3o3iYOaL5gPof/WQejDXRNMLWee2+/Ax+U6a4dd/Axbek79BL+SrXtMkxYn
SsPnfNLch1ESteb20iYhZmNCo8LY01KJ1LVwzH6Yi+l5cdkGSHcvm5dRMNgdIHxigU10xkS+no4o
7hu2rQoj+gJStcdYxbdn0vAQ5lO1yEsFGFZ+R7Lun8AK8CQbw5JqDfsomJLqBzSi64udnJDAkTIm
9DcwFiIhfrh84YgpH/PkJcno0jL8i/hV/q00939ahe+QTRxFgk6UW34DH8yOhj5EDTOB1KavWxFG
vxsbUGPytdYNrmkn032Cth6wbedD0ek3BBqzfhTR++R9CB/ZxtYtX7cNx8sr+w9hrnDT6SCLDRla
qDsyPwvn3V47R1daZTjCHwVrGJW2k40dflEjhp48SG15Lhc7GEIUa5/8HTdf+PoFIrJNXgeheWwS
zYw7KfBYm3ZCY8HAgeZUt4D/TKZAscSBl1lW3N4bSGpfPGZPb3rtmCNiEbU//ekGkixiAiHpuLGx
sBZ+ko1N21/DLlOboxFGo8fAJFo549z7M+OAJuvQhAYpV6jdFHkuFStXEXqT57rj6+nW74X8I8pK
8kI4cMUyNtOwYctEpv6nXB5vPvjSxaHUaSjzOR/9aS/nn4Py0j+ZKGVSxIFTa1JC3I3HOwUonNHy
xyJWnOU9+55uRRfCiZO62JWexRO4S1PFg/ea9vBo+gToGYpuoPbsgrw8J6eBceB1sTMtPLCkWHib
mo3L5lQC35sRwPYeIwpdlzlg0jhmM6bb08TiNORp+5d9xEQ1dUOfA0Uu7tVZgvXah2HkEdv2R3XP
2XOCJ0Xra3lk78pNZZEVcfzdGiYO2giNGLKm5xRhb0OqGhREYwNSChCmOTOXN6MIk+Zgoh5f1RCM
ocqso2Whd3xRfS9kyGPGZE64wYdaaklM7Rfmu+vqgD8NVRTfGfVvhYRojhsYbmKJ/UASatC7Gpmp
uq2agFhoRPetqgL/bvI1dKLXMHXccqpq0uClKaxg4/5goavp2vFnBeLCLGKvWYDkb3rby1avBApJ
Iy85MCpelQDodOUq8QyVApMzRSYzMuaJOYlbTzpt2ETJoGPzdZ6x8kClv/6POWg9EGNwCTeX4G4j
FK58FgOc06bxxBwfZg3rAer0UTxNPBslZVol6CiXM0ObAL72F/l9wvkcm+xSXl+2PNbY+X3XiQaf
di8acTjZwHqcr9cityldsSnV5D4YpF8Or0m1tvk0HURVaPkHwP+93cTcJEy2sfI5NoogZ37qZC6k
LtS4etC7OscMLCszpBU0r7O+Jbzw5PR2+yaFc9s/YhjzrNR1v7Y7q4NXZKnslfACnNqJgTc3/kY6
GmAbgF77XLfrCZmMnCUJ2H5Ni1LuupfIT3APLjC4IrdNDb/dewyv2YhSXIaapV3W+Lh53U8Hif2j
juMK+o6ZXSCZGAja3DBo8mmlD2ofdZ78HPyMWpV7rRQ+RF2V6I7CzgXmSFPhsQVfqtpY5okut11i
fIZUOfVPdOZppaHPqQUgtfp+Tqh6x1mWSOPTUpmgQGCZqUccbpQwItSt3lFpEbyWrfiVxtjdul7A
EMBSnouadC2AwF7kS+ZiexylropmpH4HWWpQpGg7NfbAAWKYbn/t9KDGlrNT3V3aeRGM0B+5Ga4Q
fx3f4EFrnpiZV4H5zGvBjSiW2G52JNnTcZVpXPPZojGXHAVM9zeiamUifELkqHoc1LYUl/WT795S
EpS5bpeUUWWSfIAJ05qILqkz5OOY+0DIeknoA7bXfLoN24aXEnF94yaGb20fyI3ZXokdQEWXaHfn
u3o99/4U64TNU1uV9b+TKBwMug070BMhZL4RGZvaBtuN8lZteBTkqsLqb6ZFUnp9ZpoXTkZiC5UW
hag1T0wLk9K973zitV787pTpbrPfOBPQcyVQ3ZDq98KOlXQwRv16nGTs46pxNR73QsuM+dHS5zSu
iqYTOC522ZDeKsV+Asow4tbfB+KGqBN6sKqhdJMQRa+LFGeVkaEL0p7QMxAIN9rphP2nW+VeSYVW
35Yul/iycuERBVS/XLPlN9xo86cCd9mwrzY/Sros5L+7gF9FNAf0Ky5rn9V0rXJi7NwGVKG8EzEE
iiopiI9yXvf55t8lczBePNbmPL6HHxSAd4ProkyUUS1Nzz4S/QuZZYBzDCu8Im5nwwaMFSsAETOO
/Rq+UQLpkRpL15JsR0UwiBYVwOWldzwtZaLx3kCMDVOfzvD1YF96Y/TRPiTYL6G6d7sTuO9nfWiH
stzHJqJ1xOsRhqOmWwJY2MzUW6U5YVrokYACOkMQdKOcN3nTmV2TypyEnMqiY125hgGYaFSQ9ue5
blnUQbaxRJVqw02Hh4rDjMt7wsbGhMp8WnB8K4GO7DPswREmxacyUO+pknqufyH38HsYbXGsfCeI
okIcdNFACFibyoGtJPE6mALSLqJpzXeau9PHUXI6w7Hnv3L3dll7voKq9dXIVAr1njORcBugx75n
+GGT+6awcSvV8Qb7o6KL1oAxAV+YTriOlkhAGWUeXb80J98bKvf0XIhMHPbevQd7Yj3iqbi/7NKL
mxMuYorMe3A0hntS27DrLrGCoXYmu+KFRYd37U4akwI05MIjCn9ZIq6G+S8y5+BHHUGvJCUIT2N9
3sA2KfbC09Z68+zdyC/N32+pQXwxQ/I0J9CMmUg52wTt7lvF8tKr8OgKe5P5jsG6GdPBUbhKaPbF
hYfhFhjFr12ECfRrCUN3WQXr1TsH6NRsw8CS0uPNRmaxKpHMPVCSqvBolrshEmzu+p8sscKgf/7B
iHSdbDCtl1QYhTTehBcV9LaaNlpNnNBc/2TSr8ogobhyRvByPw5Gf+4SF4BMTP8IL/INnYaYIsV4
oKZu62eEBaD+p6+ohVCI/43k5uyCme1r1vydEPDQcH6u1Uad5pGmvxNUClFPP8ZMbqyHGdPE14zQ
gQ/5E25aUQO2If/bcY7EC5w7h+9WZfpMXMEDaDOac+12lg8tEw9d0YXgx3nsAV7YX78OztqkHoB1
7QT4a7s0nOV6k6E5FQm7ZNBC2fYVfy2MjDHFf8Lync/26bLf6oX8VW7M5eu5MKjky/iuENtv0aX1
T3rhkMZKpZQ8fTWMm8Ggdol6iHHfpJ+HtWu1P8GBw7fauEIagvZtjCrkd2ZJDJxCBxUm+x+7XqH7
loWNX5jBhfkxZvxoEMOnCeJJsCSUW6v8xtLefmcsjhST7N7C0S9HM4JLRiejlfHcwVtS9x87Sbzg
8bWxydSiWW8bSRGS59SxW0LxSH+Yz8LHAnhqBuJ1gOEb969ORZRNdcrcGtCf8l4QUFdbkcxjANdl
iF/u7JBzjdX9+eLMNwqEvPg0vyzOjPQtA8vTcjEc49O5em94iWMSVubYXUqOnaHapw+xifE9X6Uy
LZXTMPlgbEFjA0ZLyNPGnKHdlw01Wl7HGo0YGwOBpFquYH9n3KYYH79jnjuFoZdpylIgB7KPsQKI
If9ktMyfv5tJ+WNG0Re8SaYy6ff4wLGdS/+oJynbNed/dvv28UibtS/0ex5zfBL8r8DZVQ5N+B+8
S+7wHskivFkI7hKZ4AhR9p8qr9wij1wl7m0XFokWcErQ36aKA2FKFj7WiHtPoXjrdnDFhM1MEqep
25/Kig6Ci4h+yeHkRYybFMNTg21MUlsmG56jTbjEaqPJE5JEbF2p4+5Zk2ZkELtkKsYUboe7U01J
m6D4Ak0Q+1qtCYLAxCu9mmQITZWIRMLVSzlMJOEaOcWy7vhgO+WEwWxeNpIMvyVo4HHjsnXPtaFL
WMLi/GI37v9xm+4z22RNVlEXXvVKxIocjDLu6p5kdyf7K+2ftLkN3F8y+2VYt5QSwHICeh0gzuut
AEsKG2It2fcyBwTlIxE+/Jg1TUpR6HjqX3yP4pCxGnSERwbk0Twa7LnntICcrnZGm+WGrKeK/THe
hL5Px+BPUr077o56ktPPts+YkfNmVC6GhVV3xPxkCg44etu3irzV2lns0cl3UWxYj1UIwXkHDlIa
S0YhOiXaTeEa+TKEoymDPYWqSE9SqS+WfBaoPYAcTORb4V7ufxwGgw4Onnb2mhRcl4zwPXunsjDM
9PvWGf14DXdxFCzE77pnuydwhuzRrpr30U7/gtX4vmzCggGBfDplcGcS6iIekWw6SfIos4XaXbup
hilKGjbbNhi708sEhLbSN00i4AjLhtPdmQ/921Qduc9WTfCU4lDMrr34N+KhSY4BV8jVbMeYjgaB
fcM79ANdKjRUpW55wpAiZEW/wwNFhpp1JFDDUe//yPbgLBpuKbVfus8BC2RDYRbc1TTar2Zl/cJn
Rgt3TECaMaqQp/MxybuJz+u8zr6klmBWLFexPyc9R6wIGAELzm5D8MJoqLI2Vd3KThN43E9PUCR7
3KcpzZbGjbc9mQFx5OT5c3I/Wj1KCeasNkbeGqHBy17arh4mf5oUIpC0V7kLTwAvTWUCL/ETqAgn
uNliXMvkOb02O+hfPe3zhXZH4vgZFSUE7uXYDVspgd4iNwm5Rz6RZdpi26tvZxiF4PXk+U2ElLV2
v6bbkUKK/OgyLNJoi4dprMG0sBgiPsxiFzBDJUHIrz+VRbbHIhKGVyneB2qzT8wivVO7ZMdqQxGk
+XkzAKklUNYalHwEdOYiqo20nNPlzU8BvmFmlh5F/20HHUEF4S6rhDzaO3kW6DKp+n9QYV4xu5D9
8uVxqeh58cAssrIUOKbCzpSfgf+0kpPNmMBSOHAUlZ6f087LU3W+2bQFK9ATIsXZST7yQLCWYp3D
tSpxcV+zqvN5j0AKpJMRwq1wpxvGI5bcdk+hC41S5lCoeVHLXY11tshm7kfPWenBiZHUlOpl39pI
M0YPi4RG1vHnOl9XRe4PwdfjEnqBTYS+faIhFdBfgCacyhsnIvJvNlPJGnc/QSlWrXSns4hTwrgM
TCPOaR5SZaYxLQ/K+z7ug5KP7lV9wul5bVkM5S465rcNPUHW/T0ZmK8aSnr1FchioWE3guWsHOrZ
HTkndGEaHOajWDHcnYFq3aI2SvCsxRLLIMvjkj089B+pYxnx9zGR4/lOgl0MmTiWGvQdUDNf/DfD
FDfJlDTm/faurdPXr0ku0DAL5YxFUIjnjM1aYW54ovXHiVOkuCmyKF08gZ5iOhqXs0h8Byq9Tpbk
ev7+NITiu2Jtn3u9tbTUOZ47h/oQOvrTOo8u9ppDYJrIT0Xs01rTIvbeKjyK9Tg68X5RcbA5bfxv
3bhh4Auxx6lSqKI223mbbYFXZKyOluHYZmkS79JwuEo++TG1BzQLrn7g3S+W0roHKwdYtqSXRS11
dq8wUS+nSZnScHjyH5pqPmEpHYFi0g44Wman0EIIn8UhjeZP9gPe8xr3pY5iwGWBJGNagY/MT/Yv
vijW674QKcl7KBqx0KH4VF8SVijyZhYHMxJ/wQtwtSNDLLZdp36ALgzR/ajqalvQKdoL50NFsPVY
0OyvSXXGvr99iD+PfV1dD3tG8nyM8EnIvzUXtyugmL4BkwITpetiarTg0GxrqXMBxY4z2tZBi+Lf
nnrVzVWlpkwKsivTdSblgTpEK7/uhAroTmbTgMqEBsOpWB5KBxrVh57Xyacr4jAnYLmq5kD7ssEE
hW9gO8soMJZzDiyZ0LpHVyML5Q2dtv0DTUgR38jSzs5iJoGt0mvXUFkdiNMZAEBiLX+UMFi+9nzg
GytlYyh7lmrsgwEOxcFDQ8yvJf2Qijbuc0haX5Y8c3yy/vhv8TcI4fJ7+V3TxIQuSb8U+tkFYG5h
4SO4Pxt2b9gIbtBdQhO/SlKylAyyA7O+KRFAwflB3XVKoznOZiHnkQxpru7nw5M6DYpNJgHHSLjV
H2+IWGetMnftYTmuB5uzikH3txmPINfbFbYJP+3tnBeljTsj0fv69OPU9STf5HvzpI+8yK535Zf9
W3wqN2lWJJaBo6pxpA5NqNZW9X4Ki9iD8xByV1r5cZXt7qp336N8yVSr7mq0FbKjUB+dTMfrFIVh
3imnWhkwYn/tbJ0qleeGDwzm7vDhI2ZEtg4FapKCLXcHlUdIyP4lxgq0TVnpoXheioVif61tsQeu
YfPbV+PsrWZ11u5faHeSoo4AmChzIL+QiLpbqgUnIrmyvJ1yFIrLgP2T4yog+CCDT1Db9v0FJZTt
CZ1cDEyjlkJtClrcEY6GKNjbk+UJAWibGK6U6PmmusIFZg9jVoKD0VFEfJ4fJsBCgj6K6JmE86Ez
LfH9pwpm5apqAhVmLG1nDdMikd6xc52vF38+iBYCbf8OKnzMH3uDDRITkYaHJZUPSEu0viOy4h0C
GG8LsOp2JnZhjBgiJByyXrK4hrOT3cc1nXEA0PHo+oxS8QcWhpaM61dt9zaUtSU4jY/BoCyEZKd4
qb9J9zv0Aa8g/cpXdI33/PGrpWIjy8yKDxP1qe0v4PSCC5185/FR3E8qauCspudjAV4HiL5qtTYb
pr6sLqlTawgafwsMKoAxW8jhtbuo+hhvchP/ivwu4rLwUH2zLceUqs/u1sXx7FEgLyNH6MzEdkbq
L2zKEFyUW2DMW7MHgFSsJH96FF4G+D3bapdfSjUHZAFL1OCptoSE5sO8jMHtT1Vfc9R3em4ONXU1
V9S0rV/WCQoMlZ8akq8dL1v1PyCTooyajKvj8IQbZmDci+kE0fZ9hiCXWFJ02XN1Bxc/3rPyo8nn
I0pPDM2a35/tZz3E3pYGoxT5kC+/t3B9C9VVMFNlFSP/GBx6niWo46fwUWHSQRly+yvZqdXVgpFq
8Jx8AS8mFYN3Bt+pzw7cjTWNII1piLhdUhP/VngqjvgS862E+UuaYEc5KgxpjeeGEsq9xNn+z//+
PHDOoe8RS6je/JQt8f6Rz7NOrKLwxNWu7jBgBJwP6jcr1XXTu4khu2cbVY4w3yNW5fMgquLiwF25
50jr7CfXS1Ij2VztwPWkpS/pBmkTMkr6cnXDlM96XVHBqR8qUu7MxVHu7qrpmu50vVd57F71i19q
WU6f34rTTjnjRnwfpfQhjRfn7CmmsRCaEqh5EiiGD3yyWDmCSdlAC+IyVbzrb6Tup4FgDRAm+IXl
rm2ZkqXwk60t2Q+3OrJgzxu4FK1pmZz6E5aoLW3Pjav1i9Jy7CyS2JTY0RIbTS5VE06lJxUZQ7qU
sFZWFrqDD0T9tbKV4MiNisxKuPeQNJ3Iy44hK2f1vu2vNFvWHDgZKvwyr0OrblWVRkw5yXgEuvB0
E4ZxhT9mor8AELyiCZIEXjh9k26inW7QxSpLTrHa+VSM6nESsVYwB0a/Quuwkl9cFruPlDy7AAtd
5c27HUAPO5Xd0rmIgW9h3EoAfgTWUSqjFoKOUXCAfCe4dR9zQrwOg3WU2uRxByxyR2z1Y3bXZ/zG
90zgGlFvT6tX5AoSABiOnavEAGutoPfsphGb88ii2upg7kGe9Rp9GmzGNvUyqDyPUunQaFYHycAh
4Wvr9Tn61cEVrRtN9QIAoXBCh+gddTtnagEEtrYg2tvvUUPrJtWOik18uhkOtUiqbwueW7KBxaCv
PKfgMBT2+GEMe3LqhaKXvT2iBk4JrcL3A4ccBsCpfqWAUNxUTJpqUpWAn3pGUCiFwQ9xzAPRqEGY
OJYu3nAZjUIssL4f5k9AK7aydo7VXWfzGnvh80meoHnYtSNFDV443VTL8y05R6NKXrWYSPDoeEOq
k6P2/K2y1eWYmBizi9S0/0XP1SQwM/juTRscZ7fmnN8MVxSf541smdWWqJdhg4KH59+K7gPnoG1F
fX/Dfc3ZtaIw50D37FemkGl4kPYcGowJncc+O0Q5kiRWbbAzLtpCD/WrBN0fv6UOv8JUTNFk64sc
52VgT3N1falrrns1QWh0CmMgnfhpgkPjKkgQBjiOip0229HH6nuInpRbAPl/kVgNx7NHvcrXFz2J
TQaMZ0J1fhDcYHKhbahULi1NhOKpjJeta8GZi/RBQtrNp9cHSI4dycpkLc+rB9e90mjWqno5lPvi
wz6Ld7eE0KEUlhUcGwovrcdmtEqPICV9JH7+a5aDkIDazHCBPirvGBIpON2bjpHB2YNgY+xC5noP
0FiX0/UuTfL0EopX1MidEry8cYUSrYyLvDUFLbYQufWchjJlUGWjE+RL/prsMUX48cHFOfyHOzMm
Bs1i/61ExC6IeIuFfPrCfGtxrZ4myHdts/LhMH38Xd51JRyWqhi6r+f8fWmxCbG4Em7TIFClBYQ/
zONHy9c4GMkNFBG0YzxLvtRA8vuUW61niAIbR303Lf75tcNbqiApqAQfCrKVQ3L0aNFrjpLWIgC/
B4BYHH8FPLQPbu2vMm3YoUlucC4LZ8DtS05GlJJBhq9yyzo+TCMSfaDFO56zB9SH4Ra0s+AP0ipI
aCx8ixOYPArWXSruOOgMew0ZgZplgVxIDJhq3+C+tkmpNV0QtP5bL+OerSay8ZhsiTQIRrGjfEUN
zSvW6oI80vDee8P2MIvPkicmtIaIhngtBrlzl1NOHZwUGnlrOPH9rfY4trEwADsvmrMSB364OC6B
IHxNSmMhiiPWYNq1Weq4ah5oiedIod6NB6KlDJk2kkGjUrs3i8/LLGtYZv7OMMRtVTAXlmqm5TlW
soHXOEk0yUDkrbe+W4ylbsKQQxEwrLeS9pwCXRmSiQIFbF1VeW0o2u14XgzXhtA6nQcGDlQi+zLz
qjExdj74y8ozTLyJQDYu99ZqrSWM7CCXKohcw5EyZlKAB+yP6WjlZqOnCuYyKM09ki1FBWpZzpom
igb7kEZnuYdEXgLT8JIEWXoM4iRVYsRP/1I7S0FkIhSU+rbl6b7oxJwnKcw57nszG1otrkpLTytQ
UlyiHLeWjJMrG6ZeZPZReYJHzTrL+9QaCfvDR+gSBqxLkOh89rxggvbrN1t4Dgwh0QYMCWZFE/eM
o8zvteqaalAZJm0xMFLBe9F3OLEz28qEZLqV7hPCF5rUWaSz9ZV5W1EqiBBUgSXQIqkPhL0mK7ha
LBIoDrniex9+Ztgt/Oer3jb+LdyMxtYFsmfW8V35zu6hFNXzO2eS46bF5DWGS6ZapwcQPPzNDtaK
mvqAC3CYh55c/ZjL0EvOUFsTCF9buLIG5i8ooSpRHmr50a+enA1xsgP+dsKLjltiO6InQMg1FXmy
UGhw3XmVog8LeD4jVChIAuYd+kNWNjUbRmCXA8zrlI6veClFPnB9qxbluhkTwO+oCSdjGaxxyHRD
q3TloFgA9OxGq912VfZIsXg6nnlen/jWuDNgxLVjDVvRLgQHf21ifhODgT42uRDf/P8edr0/l/cM
hAy900PlcteezvtPBKNpiEzyoB3k7WnBydqM5ITAyLC76LQhpHehfhEXGfbArP8ePnUv8OjHn/o2
Xq7Y+gGMmeSyR4Fv5S4iSEfSPLvdzziczC62UwfByxrqtgObm0HqWf8HeHtnLFslu12dB55uLqQq
Nm+ipNVoffQVrlfb2Q3DDPy0r4BuZCy2N83V+UZa5+/ObjPPVJH3OoN9rI4R+XddIJOYQQYS2Xrb
7XhG+Z9yTcAzHbYEdpGYA0kQZ5YxEPomOlfUbLWJhS7PE0Ghh3QUrWzhlMyRiM+R+CXf06obTTYN
K+kGftL5LXJ0lhGFQHRUZDHfLx2R+IHKh5zV1RrngDC+GyMuGRNXo4MEXaI5raurdDfBICJ+r4QB
3r2fmhRROj7AApCjc1ylASG6I0cI9mpyH26/HM0eE0VIh1OMHwze6eZCpsCRHu9ljAedDjdOrIXV
U8L5115Udm88HjTE1eqTAAUU/bD/Os83KihTCfiiNOoC4v7iGAw4Y4BM8GRLX6gUILrUG1PvSM3y
OMzFsx38oxphB5uXf5+bJCK4vOoZMlbY4K22qL1N9wU7mHosUDTcAA3YEwnHHm/MQVE0/f4mPNdk
lvwEgsmuotgUsvnqlgS0e6u7qD4df3w7oveTWk0E3HsutNkwqv9Azqo+3YrzehkveLyCi4pxjgIi
rLldQwe7AtHWSZDh4kaeN3eTyOJZb1Vme66cSv40wrDV6d9IR+jOKzmGZ2x2LK1156XqRhmgvmA4
TzM8EFWYGmmjfuifu4V+Eaw1ghpF9RN06KcbcGJMaiLAGYpAfZqZYCY5pkf+e4uV3J7tomkp3PxG
3zCqm5ytwtCzQSvpX1jlW+Tt6wF1f0fcwfMaQXzyEudrsOqpNXzdTfV3IumHtb4XtEnFmOzqRufY
/m8nMq5FuMaaKRDO3FJpLIi5/eSE5TOaFVHmlRwRXd8Ji/rO/ToOXxQWGUvA5BdtgIY8bzVc66U9
6X+RwadDAux37I2uPYVv2Tl0uJsfzLiBeiXcu9xV96fFESXmPoHEj5zMMyWMUS3tJ+XMM5vfnn1R
GpP4n8gLqNJ+LDM5GmlPzo2GPbTL0QBcG/2S1ZbTW1x4NM/IoW3lkMQFpPiYTl23zAGHLhOU7esF
njhf2rEPAt6OkSw3a/M2C0TMyR4BuSI5NMCJ+YkyF23M6IrOp5BexrCUlNy1/3pe1Uz8fu7txMb2
6eDaGFFcAx1FH9bACgG5Pw9pzEvbVBzZi6ZaXmDc7cLoq28A4OlpM4DHcpCFvVLROwo7SEvqyiT/
05X0Khu7Cn8b01UxbdT8QIzaNlksN++VfP13Pnme/R0NeSlDw1iBnIY4n2PoDPmPyuDtXr0gK7te
UFswo09IRrN5HNxuAxGy2p4yaId9KZGZRZPHt/9Foiiw0bOfR3dC7akBmQ1r8nlQR5rbwV8VmY2x
4vD2qy8r0emFFSvgwkqjYiizweqmXFpo/Psr+W67EcwyTRR08SN3ApAycc6XeXesVNIWCePn1LR6
Z6BtAiAZt1rPVBK16KQGd2fu6PgY7V4NQPfDlNBkemSFsDoNlsJamdkMq+rfRC5BWcWaqlowXO28
KzsV6/mFE8wbSUwzK8mkJho47CVLwoC9O2DNKWLYtVS+sQHMgiGAD5QPo+UY9NskBdPOGHAt8o4C
fbwxZk77fkiBqJPwTd76PU7v20GlGjkdRdUi3nX+RqqUFDxTCkpc0WBQACG8qxZxYx1z6Jor05I5
86No6dY0fu86SpUtF7KcVdW+xkvsFG14txoyCq9gUF7BS5S5ph0G9n5thofloF85p60YE60j/y6L
k6Gvd2FayztEsyup/0rgCSzsuP7/3Qe8o3chubx6F/yhjGX+bL3tUgV6HT+7al4LuxrIaqEnP9XD
ER5iKgMgZYxgUvEb3h/pvDhUo9zZW1Ye7H+HME9HiebPno6m1LCLeq4v30jI2SED5yIVrbzBRjHn
jMzPm4ajEzeC+8b2P41xWCD+8YAE35eFPuS9FCG9R+KgjQNrJ3P1DfmU0i8y770DQIclTTcJs21m
yK07LrCu7GTBjtBdt/rsmedR+CVXLHKm6D7XHBTlWzcvTjvErLL1UbKZRlXvqQ7Ma7NQtLlBZaay
vzloy6+jGzQxZN+gs7Novdxi18ke9a2+NntMIMESlQqf71sMeQaxQpMghbux0p1QG5ERUzvKwxaJ
GqZidmUz6OdhwfyZVotLlXW4RYCAxmlCO68rcMwSx5GtRkw5BoG04+PnU56XTLfPEobxT/OEW8QR
h0uVqdRwRos5HJkhRrqJMZ7d+tzgjEt8vKENHZeUWB1X4uUJmQZRKx9R+p39Lhv5e7Glk0gBvPOX
dGDMwAidXcstlWLC7k0Q87XSpIiA+fJjgz4niV1+xjTXBhzYxidWUrIxG2D0OTGfPO2TAqmt6LsB
Ic3SFL12MXlKJ0bU7ThaD7RkwY5uT0sr1E27D4z217yLjeHJp8icGN27bXPbrFHTss24lm1UzHOh
CB83WcpvmtJHkGpSfvECxBcPTSVZJmAJprFAjRhjJTF4npWBswYyTl5+fBWKh4WI/eJub3jNe0vq
8KX8oN7lpIMr7WqCyG8vOtXHZ32QJcL02y64/81k1MH61BEybnEVmrf1rc0HpMb7loxDCBBnvaRu
OOtqn+hBz/k7RAT93GViG2l6Jl5DuTuysRhfXqm4s0wsF6gf9phcpDwGH7ezlg+7b8GGdgYex5S5
yhCPVe2hq3rbzN1C9plnrrkwh04rnksIoXPWIEn8j/65Bo3ZuQfyDslxQCGlasB1u0p9ro09aOXN
KrlgBw8uVsX7A0tB/qihyN54c7yber4FOOvkjpveRuxsmkiG+WMDAjqVJfBiFGArQDrtO1iwfzr8
9VI8fq6kHM0SMEayWW1hezaE1Ihba2aNbZ449N67+Oon8n/9PiwqPJ/lkGXbVm2pbGrHSggJiZlw
IsZoCS3KDujPTmob8bNLVTQ2gVldh06X5g/h695ZC0s3PDSlmUbPSvEbKjkixBShyy0JB0riyZzd
k6rvoVyraOV7D6JYQf5vXP5yPycGCA7s7+3wGpbdnJI1Wd/e9KZ34JKltUa/DCR4oNEaLDtf5ehq
qwbrLZGSUPJJDtfOFoDDpBAnbW3irhmDowf6YHVMtFgdbhH4oBz41xovYQcs5pZ1sPdkTCagUM9p
CyAeRU13ZilEvcufIVKR99/O0DltoNLn7TC0bVmipiaxDjd0snaBFmPAjIXaJoyekKq85/qoPm12
GCCOV7e5RYTtUXqpUZoP5GBk+OEcta/fHz6qguBpuPCJwzmglCmv3Yvy6UvuTiB8ewRLfuYEJKQg
Nu1MVTWGHuBpBPhGJcev9XajS2gkrhi4vKFn83jmK0FiAYRykCcanTy0p//5snoE/XNKSQUhVf+4
MKTx4Agwd9/CX7jJ7lHBbezqEfQAkZBjuS8+d3ZkRluvMDvL2ZSEKrNtPI3pA/N8dlOMaPUCjtc1
XAE/5p8qXOo3fPSAY3lClwmuuL5P8rOx2DC4tVdw9ltmaKQ0Ksslsfg8KnI4uvzKh2XpNDZKP6WE
TUDipbMZxQXP35juDPNFzN7o3Diw3TGWd8p07A/JP1Qx+P1toAI3XDxBxlOj9JPtz4b96eP2WAmY
/ekh8Gi7Fd8GynIom7JYZUWFGxexxMiRfCZKC5opI/PV8O/yMVJLBLyw8FMqT+oqdvFTQm+Cy1nF
Xk51ubcXrNJC8LVQjohLOEDh4J2b1S5MP5FRlBBfoxDjXJ9pZA4PxL848KLCtSfjXX8l+2ef3IQr
s/ZZhxRafKiLvq2VCSrYCPLWsA164jbnV2DVMZI47+BhL/9MPjiCzr5+Xer/n83Eju0hq0huBOX6
Y4pODjbJsY2yZlfw6kZzQqayKtDr/qNuLZrBQJDWmlpCMwqXrDKLezJWcmheGXryeGGjRYdeTd7X
pRSVNaga5BIQv7yX+hU7BPePKxGd3Kqvc+2xKzVr3xzOCzIBzxSxLZPppOmelqhr75r4vEG7WHJ8
lZ+h/jEcqS96gZ5vZvKYhkGlBsOQr/bQVUdwDr7pM1Hv6C734Uj1lmdde6uuo309tng4GrUqqLWO
capXgBZksPvD9Pn7qfx/pwcP2/sNPMKmGq7iOfamrauIDeFcBNLh+QDkjblvJHmXPh2FSSheQyRK
ykLtpFKHSDMgzU3ScSWg8DGQ4swkLpuDZ85hD/VLkOkT09kd2sA6oEnJo/DqwovrG2DUwDnuDtk9
S5y4BUi71Khd9jBDNPicoOY7y8Pn+X5GxxFv2Hxdx3vxiHFpxGmr6O9zOe18ZSyS9PbOh38guKCr
XwoWOJbR12/XA5IEOW3/oB1USyomxNsWwNXICGp8EmfUg5JbqU+sAt+fpSRmEsImuRCAqKHtiexU
5ipDaAXTjYSKnvYvccMkIrNGPtEEB32RMMUnoGxWjkta93g0ks3pxIXbj9xQpIU38WvAS5qZSZ/b
UJKXcouRCPMEa54BRH424/SOR85L6RLiLW1A9EyYh/3XFQCCxZh6cCujBaSawvEJXEzcg27uqk0k
8MvTwKFicb4pDzd2zl6OMyNzPjsVgcZGjrlPGi3M5XdnfZnM9gbPGSefLAr8QYzqVs5+SzfHEcJa
hGw/Jy9xYOK0Lnlnd+GBdfXKnJm6Ilsje9X5Z0JR3pVpyG5AcSD6SefHyYB/utpqcuP+oyc6XxV6
jpCUOi59ba4mOHW2hNa2hEz2VxMcmXP+rGoY3cm7azGfo11O6IOVlIUyc7sEtskS3U9uZ+3zjTxp
5D7xhqA+m+G5F+ojisJEqBTO0j9TDRzuAnursoiIJLOdrJjhHCsvZ/JERrt9bMo21VFrhnv4EB4e
rTN0l5k+Dz0/x/nlrj07wCWqTJ/bAhTF3vKMCAhRF9JBVhzRNq1RsPAfoqsy6lD2TkKCgnc3QNRJ
8r+QdCbz8wKrxtxBDpT/dEpARlLgGCLu00OLa9D1zPlTXFS5oQofWv0ePpyhCiVMVZnzSXYm1K4l
2ByQ1g4QMu+YV21fvxTIDLqQClzT4R+qMWgn6qR/wDbnRBDIltQRMXpYWMwDhJgSRqgyD6ZKzL0f
Kmi2/8SHmikWUHMVwb/uQEsQiknhc5e2JQSIIjpjnYjwF0hLRIN0U5slXihwOQNe9kK0rdomzHDx
eIqyv/KYDGMOpUytFFItInMVk0FZf96na7mwPuhh/MrsIYVODsl6uatJ3QWnGyYd5ECkeK4jeuPX
7eu+EAAgngK81Do3Tj2QxFzsEgBa9c5g4hiK4QteCSKYTGJoUKgLBif4MpnVA2JY5+L2hqtm93f4
BA37teFPHLMTuFDDuZKSJhbxX4WgHhEHNR4ZKvDVo3BGE2iZqqsyZ7oHbepyeIYL1lzhAaXBKuPT
nE1eQ92oIMn+B5bAv0cLjtMLXtAELL5bRhPULbs4D3qtZ04Dd4PfSfvC0SMvxBr6puAkFIbLE4cH
9u5lAn4jMf3ULJSr4YtAmQrga8FBx4eFmrpTBRMwwZkvZmZwhllvbSxX74vrA8aoOz4P0cI8HDKF
1JNReiCVUyNtG4Mj7l4o7qWNlsCmM7XLMZ8SNCphx3hTr1VSG/z2CTLI797MtB8EekqQqTV/uE9o
raqJFYm3+FmUudO6Gy/GF8tw62AvumcRHqnjErP+U/7sQbas+le5jCr0bDXhnMrJR98YzVhEf9+n
h+TvPCT8IGxed9NVzAc+f3iVxBh9UW9IAnY+wsOu9qS7Rhz+Mn96wUN05Re8zbjPLfvKt0aAMXTp
VLc3UhZVuUjGdCl87rvB7d6QF+Qpq/SCyLhTglhCJD+2CU4s+3N1qU8/vWQML7EFzy3R7ac6HM5I
wFyUkKOhzJlACyO/BeDLuTKsBl5oC0SEia7NHBGQA1ELqnU713ANoqGoIZqWRdyZzMfKDz6AGoka
pfFoFHYIejca+n3IkS4iuPjzkUaTcErmedUv0UixeL2IIJ+3ELrP+xhemKolsdUDEGyiDjoWc3DE
TCQSJzqG79qiY1vxb0k42cCoWkgCBJ+aPkhQIigMXok+kyQdJQa/PIG7V8Ea8I1goYSruEywtfs1
QW3gAQClIbd0B/iPL6XdY2IeltRWdiYm/ho94c9LeCFDQSuOkXoesa5mbrYaTQ4ssx/uzkPdGB6E
0sFAMXxlHZPO1Xy3w4dMvVCOsCXCfAsGSSLnuG56AeHvJuv5VGe8XwR+Bll3Q8nh8NOZZlW7SJFR
6HG/uNjok8CKyTahFnUANj6Oh5Gc7ATQIc5VeQPirqk1WTTtrH9pvzw2Yk/qQGBS3r5lPw6CQLuR
PnJL/9/yXo3MrtGbLcDyiOOfBh55WYHI4JKoPijjJ4HJymBLinWHYUjqXBWqVrlpPOo/ML+AHaLk
ENaS36b4DnC8W6MtwOuOXcUOE/KZiMm8DvMf6TmI59bCQJyOnWGyAMAsEKYnbYqlgWcDu0xIlMA7
f1VMiI07KTqUT0GY66S/bLnJBRceEPk5AskQ9WwBAz3ZPp50gap2I7aW5Becy+k9dFa7JVg93VlW
kyQtBwurxN52KoDeCQBqAaW4VSwQwESFKj+6vJ3o9BZHHshSBCpjB5vSnoy59nqQvl0Hv58KGocY
Ekf57PzozoKOkqFwte6Jxr8woLiBUGiTrESj+4+KuE/SZVK8xAzuqxmIpxLN74j8BgfEUhXFGUV0
byxms7heIHL8KII1zF1mMYYvqDPFqofVXjpDjWc2RkLZweYcccymO93uMykxsOGO8wTzI7res+Ug
nyZgBSO2OZZxR7Wol/wyLhdbcuhsX8JNKwLbn2pAgOhV2qsIwVcdJiYvpKEM0m87/n5A6Hr07JR/
YyEtx7GOcT2640FiSxLih+Ri9QOpkCynPKcProNGXq8/CKWl9Rgmgq+6JDP+jrwdD2u2IcM75fo2
1jYN3cyn0fUxeAZ5VlasgJSX3f+QYEHFAB8LoXu4NJhySi3UL7lpXWKsi3LMeZygYUKgCOyj87K0
6c/ixpOa6lMwLSIhq8K5Tiqnp5krMuJud5GBXyEfKPzUjBmwSvzr2ZbvzUIGNSDI3tMEbN0RgKBQ
/xqhud2pHn8xSUpse4DXuYFkGgOSSUECeQSuWsTc7I57nPdLyG2eYTL20ro85t2U9pmGlEKoOXd8
S7ITZt9DKiUNAdz/N9XjYhlnZJlRJ20j9odhT6t/YGtJz1zba5LhKYOxnKGYiPuiDeeBE3xuI3hh
nSLtqDwd467qsZqW3rd4uQaBPiIqoYHwxmWnf1cqt20sFM06pqtcQWQY1eRAHlNcBkMr0+puC8lX
EfkKjrUS9XRHS/jKre2m7zHefIgJLSivC2x6Z3ANHeDb6cZKHUe4/Iy4k79ziImcHc6/Xqghd0O7
t4aJzxK7Gtk95AdwmLf9DbHP+nU0qSWaoWqlRQgep0AC9/PLyyE2cTyvfaaNDxSXCu8W206UmCz/
GfhTMa5UinlyIkTWbmuBjXE9UyXGJ7dAfOZ1KkySnvds04GWgPIpHXH0yWiR7mchTNYv9I19Ckuv
SsqeYgpYIbEy2d4sNyE7QqOu/hJH1q+ma8hyPpyspUPkMSuwJDFJs+viluY8sRUzzyhyjYxtQMk7
sUmZH9diaSRIOVLI3CRwLuaUHAGz54ROAu9P6QhHIYzJIBH3u9BeOf+2QT5eXb25Yhx82gTPWMGf
p2CmdTWq60CIRNEbvVeAMrEGa6j3i/CEWhLhc4O5YPEuuTwFtfAaHuWPxeLNpJE68p9WMUhCf54A
XUGmPtdIsvneY2JvpUzUEvxvLqMwi/jZBdOkjB+wMumqPW2K5G850UgQOk8wz9p/Hd4n6pf6Wgci
gSWs1MbMZ68H0XOa6yTq4akWHF1gD2m4Heo6tjrrp3QPYjvMhPxAqb5JLliEqJ8TcWj4OEBTO3pT
ddgqxYpBJfvIcJ0ZICzAmc1whI3UF6gP2CWeMcXtzdvD99u8SvsT5lgnQtqC3WlX8KRdAsrVFedu
4xq0uK03mp1xtwR7ZcbHxClKHZrBBWqZhA83aFRowB127FDMFnxh4gsIu/7ccs6YpzyNOv//2Zc6
EiVc9QwFcFU8bvoQTI6ekcaZDNRB+6oQ4+CU8c4uMRbRqx4x6tAj6Fuog3PsyG/zqa1mHM6ttwGe
8Xquf0g2oKLjfhnsskZf/cQOnmfDRquc/SwKyEPd7NpbnbVN+DLr6qYSAYrNBWZkqaJ9Q1fa3It5
WjNIsbhUaRbChV3UzhykHpFluezeoXm7jZLTEQZoWaM8wgdg81A12OEhQhSoQQVolV006880E3pf
cGVfelfPX4q0IAHMQCuixzzNTgE2wepsp1UNRtDl4COW5L6parXqF/upQFHjTqkNAUNPw2zSxuTI
dHCg8RbLw5OmyuaUbINCLxN/TrDiMk+AisBQ8dnRqI4if3RHFlsCPZSmS+lDXApxTeycB+6v2xzS
aJUvhaPjHiD4tA4RsHQGAUBL/Tr8gifnMgRIMGa08PsoGAokRKD+Uxu1YV95WsotVI+rKUKxdAVB
xlgiR3mIEKXPKojfrp+v9WF5/Y7XVg3unKhp+lGP2tOqRSxb9XnsMcXDrZYv9lSvpmmeK2Mhd2NE
7gIvT937IN2PyD9s/o+v6F5A9PtfZI6CnDtTbIm1nnE0eIJFlG3BZmJaNUc1rGrtsxuILF8fbCK8
fsLGtjTuHwbuFbhx/WmKMXBBwYn+kAD/OeQ2mlvaaJIyjr+S0L1+UzAI1bK3DaR17qdNlOnmQRtb
Rntot8uK/R8YeGJWMbW1BFyu8griGHPPOT55V5L62JMu1IwMIYIyh4qvBJ7JxcEKWbfzx/riaFIN
IyuHkzqiOt8tTq6CMuK+59EBD5f8QD52Bl95UwP02SeyMoT/bi8JqHdn/eihGKL8rvgEwGUGvI+a
/zd/LbyTYTVj9hap42+9sTycPZX+gZfGEC3RigKlg6jw/9pjv0OkmE3xsyNqkSHX6zfSRY+1nC35
5B1LqwMd53JwZEwfm4ypbTtLhyqfTPGZL6v6IDuAsK6ylZWHPI1UzvvWMuZ3zu0pEGQFHX+aXmeq
u8aw2YN+XMuru2jpGNUjYnNjvZL3659QorHVhtMgMGSKvZQtlWg2ysPzzXkcmXk8wEgkyWZCNlPv
x4viNqhuJQT44OQclMHLvbJL0sRS7gDIKoitrhverYuh+qiSx0eH6O5jYagtjzDV+xKENrSyC1Tl
QeAMrM3hmgxCWxiQZtTzxegMjpnjWMw2Rw89V95qXLkJd9x8u3OG1/yP92NVO7YvYiy15n2Pi2fC
/XaXaL1Ep0HjpzpPm93hgcBP6LNmwyllnfU4P0MzZmty6mM0YBNCXNd60OKaE8pAgZ9uBf6OZ4GB
4aBMQViCEiXLwNrgJhem4pIooIaub64t515frdVlkzCsrZTa3btMnXfVlEv1cASQk1jXkq2bw80k
QpPlRUdADuI60M6/1YkBZw184lKc8tBYYPFrEI4ANmUnxI4/8w8ae/WTW8gvlt4WdeKv6Skp12sh
IdcC8lQJTrSvDrvjvUkplm+Rj1z1L8Sn6ctAtzo7lD2tVxR1/L4l3YUAN87TfDChi9/TfXKZhg7l
McIWSjUT5oZy5rrsW5gHMnyn+cYDVE3dSvXCRcwT2Su9adWHzD8sHvm/TsXm9CweTV+shACEcPBA
Eyh2JmNCVJfF8046k1h7hNUWa1ESZVCXjwEx5XKnJGl84xJw2GRNoU0UZNlebyrDPdRm8AblgUe2
0IdAyOt4zVknwEH14Wx0LhHv/mGlTrrxcKFixfyYEJTf8lLJVRBTV4GGYTXIjVZKfXGk8O5UgSUn
FZN0xAcKyM3vWeypF0E6EelAkDXI3cwTK/E7Xw08LQMcIkJN4EIFm5f8wbwkZmBxAOF5XqvPDa51
W+Tal57UGnYBvkZC9TqlQFihYsBlvlU3EwBz4x+j32gYo/Iy0ZJHb6D31d12bavKARrYHibwjE7K
42+YULUVoau/QdPF3BtHGFzJmlwIRnHx2aP31G6HZgGsIwz9uFuXrm7ZVYH9uOqvsBRebfoAzWLf
mX0LWwMQmxt+wow3MZSAF9M3jtW42ZrQFqjEQubOeSoyKcPSAuuQKBsh1lWx4RovKhoGLvzTW6lY
M9CCr0qgUCuxnv1ndKvwK9vWmQD1JsU8WGXKlAuwrhFbapGiKPLZsEoPH8tuS6inj6zt8qL8f+lG
qRc0YBasFeIaydVWZJJoQgpzjiAIaLCs3iKZy84gNL2zRSru37PYvFsLDfKczZgNi1ad2/rjUnTi
znyVzECgXVUSOm0vsaqx8U4R6uvoxYdOVftXFYhwr0y0FexErTmk+LOAHd2k57tvPT8iXX66ml4+
LgfOj0hqQZiraoZy4Sjk9qifn1Zdrv9GW8bLO+ovFukQfAFxAVRv6YNN4k8GbIfILvHOwMq6RdME
MfFuKMM5pDujJd3P+kO38RJOF0eBavX9t1HreT9XngbWBZtSUgb9NZji7VtN+a6IHo2+ESqakB4V
uhIUjInkT3hJ/Nek9+gaIYy3k3F9n42o9gYTy8WKOzPVPA85V2AHl8tKBhERfuwMsZYVWIV2qXrC
ZD3zdXRLLLoWiMLrCWWzD1bHA3ggDCYTpgBbrN9NNOlvrfarxNxMRSDyTUyd5LDJT0nkVI3OLtIq
/3JJRHIcpzAiaEhMrSfoL3Wiuh6KQp5QRxDJ5jQDMbJ8QDPNv41QgWVJFm5uT9/cvfjx7+QXlxzL
eVjykJGthJxeyp0hMaBPYFA8Niu98Zs7YDKaMf1SZxrgQGzGSDbz+bf11KCDMgD2fjMEYs3v4feC
Lt3AFhH1Awkxl0Niixh8VHwl5jK3q93DSbqMrxkfWKwDCeO/HuJ2EohgaAiYpLFYQ1QY+maQwnB2
ADvGJ6WoeoPYpkeEFbDbUciwoWmUyBmYONzcTU8ly00Emi5SFepvHptWmodgeAdf/j6GF0946zxS
Y/VlE6SH/F8e7E7Qn5U7bT+iRK8XxUw2MD0eVRb0m8NNu/EoAl3OJqTGKYCpxGR5JdZQnpSXKK9Q
iotTweQXa8gASbzrUD32K+QT702XftNn1XeHGGPl8BoM8HKL57rIpBX5MjRI1qgn1d7O0gP0o2MQ
UxKMnZBlIpA28rlIIjs5Giohg08jVxCY8xg3j6kwcUhhbCnEELFpHaJtCU23W8j818eOG7xl/o3x
nkUUyMNHZ6QpHj3lMO8JmOdBa+/3aUGhAuZnPIJv68hS329KCQUFyeUOMWAZ89nVFXj43LZYqM+F
CxbhN+1u1zfMbfy6q4Td/DK6YHh7hshYhbdYDT81NPQ2a9onAfnYIvbIYOQjFGyvD2nQMOEcubCj
yT0oHUtESoV7Ui/fCFvmevQIwa8/HCqtuMsfTfywiOev6LMdA4lNAl+oN2on1Q40Ch5tyvzd4VN+
CAlpzItml2Z4j6Tx51oujrHJcsK4V2HdPdnTVL4zdXahF5wCdvrfeukGus4gqs4fHKCgjn4h5lHN
luoSYR/1/ZYKM9naZyzoIfzbzkJ885yzRo445ipnrCoBj/AFTrqfWsYpaUyoc/77DByvBuwf7hwt
j2PUEFr33Xehgc9jKZQhFr0KFf58ks3N1EwkaQDY5MlRbKVn+Z2GfQP4YALNjLzbqJTwCidrhRgj
vqcyMMqwQyhwlVQ0ZgtxlOgc/YJ/maYEU3H77yj5GqUoB7YKDHUu2vd4VxB2kI8svSWADPTHdsv1
CuPJ0GFyZfLOxs/tI++RgqCYhtGKOT/dyrl93cR2iHXFqg3eOtTkxfKaybp8ba+N6CIFNsgFGZOj
VoIG4n7+JWaaXpyyrhSeWrwFeOkO970kJLirUiNvRDP/5NMQfnPSOdhVJhFsIRageZDn3tNuTKz3
72rBMvtgMqYIrcL4nc3rX71nsIuobQpjrZmfSrZVjcXubY8RmelzAMxLfno3dcTiwR+9fruQvIpA
U/C6TbT7kuob1uk60t5oVy4lT2u1Pgz/nRH5Gw5CJQY3Vv41h8F1vK0Oxzmh0o9xKkvrEshMMVCW
axoSlGz7iQxxWG4g8DrWV72WLBFUX8cnqdMCPux+6hhtpQkNS6F86avntucw+AkH514pM9ZD1gJV
gGT7kI6xLfiFLrP0c4Ynb1DAQXI/uhMXSS/XD05w9UG6KEiXlrCU66AaOFLVkX85RsKsFF9oN7Oc
ArddqeTnwGq5whuSFQmyeOpYQq+zR4SROmQjn5L3A/0XwIdPg6QQSgsiTmNW0oLGiecwzRtYm3X9
mvvM59EGXnA4k9NjkkKN4PQfAAIVAQsId/N/Z0I4nUYS+/svkt7B3lNflyU/tMnXOIvBYO5RyrXc
XFwlg8ED1A5hXCRb2LpJ/yUcyxrzTedWbBpNxysDh7oFTiGKDI3j1hc8TtuQS31mU5eMwlSTwQY1
NycWtOTwM1gHgokU1Y8BNWvdSGLbkoadnsRzWj3l/r/+V24Y+8CTUGEafGQQ7LAXINNVXmv2DHoj
xXBDNgVZcA7ayjOzlUf3qAKVEmqfMAe219URRUcgFO5ybws5ed+PzUIBjA/6+xUVHcIMkKM43P7/
ozWtHlC9p2o5RxhF97r/yUqPQ4QoO902uNqAgYV8M5M8Gmn2vBMqp5KP0T7RMphsWnPS77QE3Z7K
3kbQqgcbuNuVRlsrohGuCULWwviTNabiPdxL34vxDNZk1z1yYk0F8quXA+kpB0vGBkxzST1hrDi1
A3CzXU46h9UtfBsJAkv9DzXj3uuP5T4xfwqsCvCLB5WzD62dFZqtoUdXrVU/9yemSNsbYpSHtWQu
ro0Nneom4yDT8tncCO+2trsookaCFHysG4ChrSuqT2BwbV/aGQIQ/jzuDPk4381aiQpQwfIFZLbN
tgSafkyNecXf8SYIkr6lpAqVUvY5Rhy9lWQz6lfU22XjABxX74/KjD3FlQ43O9l4if2CZU3VTAQS
B387BLYPFHVzTgHmRRyeYe3hz2eC0KT6N25QPluzt27r298gJwyefY9XtsO/Th+vWm++Wzv/A4dS
D+jRM0a2/QFKVP9R1F+W0E5VphP3U52AaH8xm7p6+f1gZUCJ4PqQHwIB/k7GM6NauKwcGm8Lcjmo
uARH4hWIJEQm64tAXc2zjfLTmql7iIu1A6SY1UW8NLOUNvz8hp7ySJXt0nc6CdK9o7aUxLjegHQS
O2oVv1IivzL6gNVhcbJV66DNcFQCUsTMYM+lkxSvHiNYTZcuhlHuruIUSmrwhddpxvsJ1/Ogdi0I
8AeUxChJXNyYZKzKvMmW0kvZg3PAI0ex7wcGgO1x6laoA03VBuQ85UpDF39Tvfmrb5FJ8GXboG4d
30dwp98ELx1D7QViTmhYKAKuTKpPyB3v1dfqMfBMBBv7raF4g9AQuwpx6vw6PhdgviXGErVAI7aU
JWfnViRz31jOlHDxhcEjt0ZZpmXLayjRBQtrMN5HbtmL5UprW4LuUhjH1Z2hQ0G5yuf8GMAs3qQ5
R7v7ws2nOJzUf8xjGDhZbEdPh/c3I/74ezLHreGs14F2MvTMvEIED3YPzLN95XS7xMOxS+iqJXKy
hJiHnO2VEB/ZQrZyumkExinrSE74rnrA6KrLibzVeLwmTDYZF+b76ME3bxtNEsReRQx/acjTDG2B
sHQvXn/EjRui3xtMFM/oD0oyPSZHIktVBCF5GLscsYM+mG1eXycTiZX8s/EX86/YfXgkHgvSzHFJ
nF06FtSdp3AhL2KAN0UUkYFGLeFFIPHcEvGv3Wf7NIWNH19oDA6MBsLEr80RB0xt6YWYbSXNTd5k
X6Q7e2eplaBv1hYTwjOAO+uAhJ4g8solEDAIsXiZg7cBBbahdumpchQP9kNEYZEgGm6gUq4+zDIe
8XmjsFvfQfRcM6AiMuLi51+/uW/evlpPTooas5l7JlE3QxxtPwXfrtsvBaSTZnl77nQ8BAv/ZEQq
rM2vZu/6P/OKBYOljxiXCLEuhFWWwkvRrNLInu/Y3U9Kvrer5OKBf+hNvV/HnLwoskV1e2ommCKE
Apb3UOQwiy870xkpocHeKg5yzN5bRIKcTJfmFqrY3K846P1rodPL4k25JhI3tBWsRSu4j25/RdCN
ChDbkar2LCO1M3GO2RQhI1/L6qTncJ2xnBZi1burD24j1zd2Wgj97wOpMHhU6Zr+LU07XlIAvFiH
k4Rr5J/hCmls6oSjPVKJn91vqFkNNONLxKJMaUxR8fczSC0W1ZRv6lBVJdphkBhmlsUwMBkn0wYq
QoMkZDKRSUi61wDJkpJvZDB64bbC0c8A2hmJKZlYYxgXm34hlVHn87ZqtFUQBu+wxNKyfZcdEJaW
DSY6+VJo/feRWDrxurDt6Pzn6TTtLEMdsNlS9PZgcZlvYicWhZcCrQVW2tS5UWFvcY6bhO+oDOzR
zuEwN3xZzFcDsIrbroF/6SuRNMeQbBOZIFnTGCWUztr8Q/DBDnh1agkci3HFYawzpZTfLwm9ntJu
x00//IGT2mODqRi+gbBgM5jdI/0D7RQVVoyWwc4tTbyY6NnBcvZb79MmSfwGiVhQuhLLH+Oj7tC/
E2+QhiLpdkCY5zwEphpH4cmt83YknBJpmjyGeMGIZL9N+38gnfwNDm8lk4Wk20ZYluNWl7aYGKK3
VT5iebOcj5623Rv3I3zFb8lkEpHEqgDwiGFrveluPAwR79vMY6VSRETKfhJBBa3RYpL0Z+yVRIxB
iXcjGWSPMdt2hAND9lxDRIUsskX0D+Q6NdJUtU/UCE9Wy8gR8r9g0dqTLrw8YBb+EqUDtRi13srC
iUaoLDZQtUj3spDKlf5C1M+sRxRsZ4qvoeLRjsdmzXeoW5i0Zg/mHoPbTawIAJ88kdrWdG5xsxA1
8DKf7r0HkMgXNN+IAZrogm2MFX+icgKgqTfr7iOzCrmLqGT3912IIuqanzZdmyrgwpO4Z53M4FR+
KA7zmO0WlVso66bXyS1HxQyULnzfrmz68Wo0Qn/TbgpaS/AkPoDsWW1XbTV5/h09wSFw87wq5/a3
Lk1MgZvjG44SLnGqeb0nFMYWjlKL5Hmx/wozzxs7XQuGbg98qiPAJxGvTYyZAh0WdCx0wvi2m+7r
HdFVp7Vm1gTdGzi9ewGC/TD+WDhdTtIU8fofIbrWuNeIfPgsLS+jZRhVAHy8uhsCHQPryz6tDKz4
+DTbnTX11w4W9lURmrbZgdX0lpjdGqoH5YD7d8BRJ56pnGfThfJz1jUV7keUpUNOOa4376ML8g3d
x4HGJb0WzTILoAQoX+MOTQ/gNlIOKJt2L0jHEHh2+v+KEGliBctOeXNkTA0AbISW35Xa6LDqV1Hl
g0PC8SZz1q7R2kyXdnfXBFca90fJ97BB3w9S4/jIjDHqGzEnD8HKpXWd+A8AKF5x9kjgVWb7bFTn
WY92K4WCPlcas3h2w8wSYzYtWZikgdaRHhi5vj+zMk0Hj5vsaUYfKfJ6zxWv/POwXrrikT8tDIML
abVLfGSPTzISd2oARTsEp8GpT1xGkBDNJptxvDlkthpdqnMDmnT3qaO4uBH1XojH1AroSPo/LCuF
JQxnE6OCiWswkY4nAnprm7G7BDFb36NqLzy+hCCsyfdI+jamBzNufHZtJ7h2QyKaaeJ+feyDgATo
m0UbQmAPvHhOmR4PKFlCPwjz8XUDD98TJgDw16l3X34C8lOWYagchq8VLufHlJH+bmp3U5nVEX6r
FnjQkrVyF0OReZ5as4G3l0iGuJqAZ8mbjGMpKpLI1j5OnfsGJewDJE7+dNUnOpN41+3LhwOsEHPc
SDzFUwSK4jjjJs+zaRHXwUgi7uS+gATCOm1xVB+P9Df2qU17tmRF6fo/bc/7vMtfsIgbalxCRp9b
nw4ipi6d0DLOPcP8hGmWOg6KrosnCAbvwKieBm87jnqRJYREj2l4HefH0mK+cUu6AM66xuq9MQBG
rJawXkkNPQHj1Z3mtTiTqdVkwt/D25xwut8j1A59FzOVicmBr5w+mqsKYxntA/AzcemeJqpH1C/6
qLVl/Sk+7eQLnXsLffJqywq2JEnCb3ud79moZNwxBjiZy8BZykFdsE5cXH/5dmhp4x/oCiLTBhvb
7Aj7f6jyJ6/Sr4cHlNz8w+iuJZ6NBFSElrjcJyYNO/kBYIrLvAyebzvjPusUyPyXGYg7vypBMIra
1RSljAvIpKQe7E/TraUKZ3YAW43RXm0/QgmcG1bSpqgwsn0kM5r28mWEyPEGtEZJ3Upjj73gKYNJ
iwyxh+mhKMNJ3w9qKHU6nC3lNzUf6cvkQmonkWy6kkSO97ChBk0lUu1Kv9E+VesxkvO+CqabZfRB
Arm5jF0enjIQoqVkbWXLn5m6S5obWHD1YLKPQhr+vE81PzhcLEPxtjazjw1o+KRfIG0Xqc1eO62v
Wx548+yYWLXo+BiJn0EWKc6nfpUCh48UY9hwVKT7Btl96V0W8m7VjZi42bYqAOXe/Nrw71Nr9Utk
LJOOSFieCTbJTXBl4WbGi89jSf4nc2+2S6y3VLWY4jV53G4pJ4CPRK7bji9d3gM3FkuBbcZ94DKb
Xl5KU0EPxIK5RMd+uPt00Z+eMDHA9cDve/NOq2igPjziqoDbitagy0XM1n5LFk45O2X4Cg2XVeMC
SAur8zs6oWgvee6fzP+xenQ5mXtiSr75Ilwdm0dI7AWATa5ibjgkQMzVyQsEgvu240XGToUspKuX
iH7TMCv8kOVvwtw5jgsqg4IKJNhXArggE0r9uXrVQy84Fdvl+FN2F48nd27njiA45MGHZvKDrnHc
H8F40S6og+TNzeXrSBPxEc7uVprOgEtUfMIlkVfQUonFBLqekd4XqLoagBpNfc2U7HNdLSiWpGEb
T5/vIhJPOAoJOUUKWZPOFzr+8GSotmLeo1x6cRrTP/XIOOEidKi3jjR1pFYL+5ZlfqX6KNySoHSq
Qw28om3SDeSbUmu9eJRHBGPp2IgizKt6+R8bQN+uaG8UmgcaIhhcP3hGIV3PDtz2jfkXadfX7qKc
PT13bFfi0KbiN70258JW4wCPSy/T25PsNj+SB4wIbmTYJLmJMtsAvxDE/xDE6+IZha2VvgAkwQH1
ti+cbr6U/V21GbG1WwpUwXKEiGerd/rkZO161igthdIqyX0P8ID6FAP1ZttN4h0thTUIUtNZ57xP
f8QqxXMN/JYc7GOKDfyUmlWgy+iC/ILx67BPkBXRq9ulrcd/lArkc/6qtQ29szpPt7s+A4GTL4ol
prcEs/VE7u/S5kUpjNqiobXSvTLc/WW9Ni/fobcGhlx41dWp3uSISXHl/qVMVc42MqyLh2ymNVhW
uOH9YxT++v2XZv/ag1nWTS6ebDfza3DFTHgsUMqtIXpAepL/3KfCnRM43UV/iwwtvx0z6U2FGTfj
dzrLJ+nG+ZrruG15ERuqPW6ohRMj0VJ1DvP6A9btRFlSAwVNAiQsYNB/NPy4mhQPzwYf6D6DiqNm
kLtgNcFRVQr8EWSVPSArukz0A9YDT9vu54rNuCuMt50Xh9EPRjMUwvsdP3eLmdUXjt80O6An2W9h
Tjm4JEuZuro4EaY6Ym8yzzrmBmzMrkrtdBYXOVGo0snIzd+y6WfMIeJ5PWPEmSV78wgF37QIdBuR
2yc3WIlYvOuH7nQGHq+2W1y6HuWTI5jJ+ENm3zEwOUrqIG0OQaOu+XQ+3f0zSuxxw22PCZf9Sfhe
Y2qACfd5yR2iBUc1HlGXToE629+Mxaf2y+gKieR7uUku6pVAjiG2uNMAX5t2uXKOOBWzhx4zcxe5
njmFPg+Gl26Qv3s6gfcvF1Me860FJLrydrhIPF6w6+9+/PtuqhBm3BdDv3CbSfzFNR9QdtxWTpmL
WxMdPcJyQgTlkTkYVVT82v4f93fiJvoaaNgzTI0CUmMt2JJ4bgVdM2O54de6Qt3enJrx88mBdr3p
ukrT4Yhqsy314fNRo7Uxhjh5pIw9DU4I+KoA1Z+XIFNpllHgBvfebtvEcEO/5oAYInvrK2VgBjaD
vf89lHPJ1QTtnW8aWR/ODyIZTF3rP5XVxa2r/ivy2hKCogFVjjerkkEuDqJFVipgtjQ7wRlMRJNx
Wi0GKAi+5XtGyiMsgJdnJ6O3jdnHSLxnqZDK+m6z20LX/wix5BN4oKRBn/duDPiOo76+syKfKmTu
WawMO/J8qnfnJm1mhoo5anIfSxcyGNlepi0MOB/DtGo6mQAYd/EHcjtFL5n4FwjVERm9mYhxqENJ
WH+A0P1MvP0DmE2+AU0NbwpI7970KEJ4PUlkJZOBE3bMBy1H79Vq14Bsr9fdYqsp3MnFyY6gYSa3
8agkwn6cBC2QqZiVE8kv9YxoVYmh+QRmPWhhyhk8N7aJgpDn8Lo9X8Ce0izZFw74r7ppXCWdQC+T
FUaCCtFd1TtWY9QfY5Z4D8mMFBJGXkA4BrYDeVeOqEi2mq/cw2XXjnfufKScqwPHnaBc6HvHO+As
nqDkoInWVNZQbfYSqJJFMebvJKyMB+QZ7h8iLUwRd7XOi6HkBhcp5G1+hf3RDvqyxjkSJ4fXvG83
B4fNQe2G1wNJW9DrNf0P7cYrV6F6pax2hSd7qaVtzEaPh4NoBrqub7zqSvR0VFBXH+cZ8VGjfCxU
pqlsDoAX3dHqEdLydWxmSoQKJK0gdTv24ST0LmeSGhIxj+Ki1WN8JedUQmYOSztGqyk3EcCYOmYj
h16RGX1cyVUrXBQAyrcqLTRsEoeONFq/iZFjl3gKzHQlIaooO61kBvoLOkAMXhSQz3DGVjtGXi9o
sH8joexXwJ45Yzg62DkE0jbi+AgmhNxpcq3wwNRBScoaSkO3eErPtk3D9yqzbUsxdNpUAewLefRy
RT+7cf5Wet9ZO4qnt5NkMPUGMfO+2OBYwo5Pk7216ZuJtlfqJafN/87pEjG7I3mTkcBTmkOx/ecV
5a+yDOwsp6eRXr22WfHvgDzJpFQguI597U8QTlQAiBBdORvX+hvQn9M6LlQLkUUFsIjTXPI2/i3g
su763xALdwYFriWkZFHolvTSVtUYyEDx1V8jyQR1+SVGPxTdvFY0pT2nj9SdqWi413SvLajoWoQF
5+UwzuoDJMFhAgzRBA6aK5VLVq6Ae6bkFA+CZBlFDvkf7Loql2Q7COKUUs7SqaLG0sxJBs52Mr5T
kVZiIIp5bJB8QnhWoufh/Gjam0jZNNXl5tL89eQ0tdqrrd0nAxs2Qv1JEcD+cKm1WelljGi7hboJ
88BGWtuu2IhWgAtLrU601LHx239pzm8KKxWxyMawA44icYeXA/UpVdlA836Dh9dxzw1G3loYKxC3
GnuI/g52G3VCLm8+5kd+d4zROjeJgkh8FVAfvZGI2qIG2TwwIJptpFgJttMFjlA1g+6cPBa8yV7F
FdtyBzRUAlhsXF+kO08/sNx7WOiFEDJaUL0M50DKCfwI9PPZGeljc02B6yrTOY237zhVFI1T/0pq
V8/7IzW4HeekDbphI1+uB3egpfHbvuhF2LdEavNUY5WiPvFNRKQ0QhrNE7zSlX/Uv//ZbNGMPXfA
nAKbNgROdP2NlcO/C5kEPk6fQ3U/7Xgf1Y9kMeTwhvQJf/9GE9qei7VzBgPOIZsxZWdvUcMEII93
RXwzzoRdo9qzpA/xlarP8pW8Ds5GuR3FbZPrQR5sbMx1K2bEs9C9vpj2zIKULlY9/fpR3/stj9+z
nkOQDyR2DFySZB7gw77yLTQcFFOnAzCoGMjthAMOK9EjsyxojHPx8XyUjUmu6DxfnbQMU45ULAWG
YGfABbkohU9L4/Zyd1EjWNiLSBKBdbTmtBZOgGP5xuKRpT9zYaFajaCxqtW6inFUITVtUtK9SbmW
7kUt4y9XNEBWB1QwXzmcuWy7G3vGAVNBSvXr1gLj4BTUbvYk1cLC0N/7vCZV4ddCY/KqbW3aFhrX
HW9Z6vi5bkMgbNVtdSc6Zpx297qhb5KYL/TBbvMnYk0+xLSsFNUZZki0QiEix0zS+7tjwTzd9ZlY
DUpglN11DP1KxkFGCy/o1cc7sDxy/LTWx6qQqb9hfThaz574ec37JrFQTTcI422hQE0e3SZtzCkS
mNAnSvQ8AzwkG71IF8GqdhMLPje7jOPR/f9oCUTDIBt51V/Uo7bD5T2hVjOQuZyU0yJxSw9N/8T9
TtHh46wvv4P3Pf5Kno/05An79piDIsoL+o5ShWjSFL0kS7aLX+uG2zzhfrhc7pTDvJepxhAtzKaP
Pc25bSMDHd0LOdVVsYIEelCfJfVDcY7iwQuNMOFypx0ZyePEKEQMUNyCezxx8rD9Pqt+2H0XDDjk
TgByMrDgCCponcBjYG8Imel7Z5QJpq9RjQ+24qSlb71eYsuPczghM0whdWQRyTaf+6h9BXjE147t
15H1ZXhbI6Ik6wzP/NP4RQ9pxOU3MNWbB9KbaVp1pYifjxtHe+eX7hbkw+51xypjDBA3pcPXHxD3
l4OyQ2x9nmJvUgrrtdUnDKo2DLsEreKSIuJXHM/3+AfjjBGvqh76DiQ8Nz7z8yxLXVCJWaDGPNZS
udLrGDk7ybtUB5bbeDPqXHStFWnToVqwpLHWlyFZmpygUX6Mdh9yGdxVPquKYPoYcdEd2uQqeSgg
x83/JKssEcItoG/se5Lb3G+rrseyZ0G/lKJJRiVOqxv0/TN9CpXGGqOIYRIz0YttJvbXlRz84pqU
LkziAAAQ2kYnrDoBZm7V3YfexjbdHVogKgzAXDTLiVY6vsR7bAfvQH9Bt2QfJMVaJECknEYXkJZs
84+EvYyQ0qRtQjTil3jReAG135eqCwT7PlgVuFY0MAgceq7b3mWxkDVxL/LQmO9HE+/IrLjbfhut
BFil2VFI7F7Mvmi0uaOiFuLSrCwBzfg3kcBv+gXt1+ednHKu684HJBt2RKQueG+aFZocvqkjtq3K
TyG1wVbcLJBnOqh4B2zrMR6Jq5NHU3S0b4cFElq1ocl450WaaS4Bkr98AYzxFz3XL8J8LYjxiVnb
cc70y+k38H1vUnVu8ZLW2jSC+czDlGZ5fwmSVMfyMNkTGhDCtGKbO9ZJWGsAZGoqhxMJj0TBXU0S
9fgCaudyn/z8nfBi2UKEVbjscJ/krG2c/rS9CyQPhyGZetm/+auV/U5cZs0NnkGHMTo8hA6J2XJE
jXFWBC+U9RJu34xN53BnknnQcIwpb+G3mfCP50FwbbxMffh6HwV88Y54TZGXX/QfZOQMLAb2Y0wk
2hqfAPA3TJIH5Oo4kleKqJ8KXwsRoN6Kft3HwJ947m4Z2d2+eJMHS5Lve6cW6gaN86dICYJIpa/1
o1CyO4ZyNxwaCIa6h1bxRIGh3C2DtX5h44ABx2g3HEFL7LMl518hWc0Cc1ZC1L25JdGUqzb0r8pY
NpSfkfwDIyodIfcR6sjMV/w69oi56+V+2WzSWsdQOLEcqfxpNbl5AsHnwsEkJ7VtQ9GV/oe0NMvL
fRuL6+zo2DWUfYr4jSUri+82LgYVpeYnzOtyfLHm6UzfqQYesGBXZ/W1VAEVb/g2CwOlfOoS0RnB
4l5x8WZy492rJGlqTHV08M7Mxk+eZdc0fSD+e4hA4fU6bJ9Fyj9Ie4cpPcMn4FwI0b5k3KahZGwu
zTSvkr0x3gL1wPwWP9h8S9uORKEyP385sPiiW6yF/fjJofyUAvhciEhZztjEdN6XDdSnkxHlJ7XM
/gpxGXjZys9qQkbDWswz3Aiqx3SX/0nIpCgrBN0dQwFyvyBHASarajaoEpr5kdtGpWS0wQG+Jl+e
9h/h/u0+ixA/EKyqhRjIwiooQxkGRqr6cCW4fYsb8omLy/FydeZEek1Fw6EFyhRT3Oj43iIrZ6ba
Z4MGZuV9scGtMFpxSAQCCrAKG8j4kABavDNyAq1kHtlBIPsLopGjBdExvywH1JbLrhliVsrXPQRn
HMS74S0GKCT5id8HMI+5tQEzXMXkamCpZJP2moUaitm4DIDu3OBs3YeGzeXa3QQuRtfHdCdPjEvv
L8z4mW0uR7517v5Lc9DZNEWmKWmfELTsrE7XgzmRN1dhphoS3U2zdnky5snDppW7rVENpoL8cTN0
kBnnhIkGoY/DHixnXUm7/Har5E6vDwWct32J3EdGecdgaFeR/Oct2/LLo8QQ5RllWCa+OCEXFNi4
a0CtByBRxPBbJ6TR8V6baS/j7v2lNnPbw8219+r7AWzOWg2riy0IkhJLW28zkBpR+V65IP/FCKqB
4Z/Ep8ZJRXK5qibdj+RafFvPvYB9Tcv65LoMyR6Ojis/v4YhUOwrqRFsqHOcFfQ1FWOFxFuhF2iC
gnVcmCU/BOI4BO1+nwRF1bExmCiQw8TYVt3+iTlF8VVo5obVeKocF1gKeZuluN5+aeoA0ervXejA
GWNAFeAt9XE9vjyxrhpSZmn0rRTtw+lFiVUmAZQ7YRXZB7NQxC8Y6JiSGqPLcTnLJLUoApD3Hg3d
IdCIL+j6uMjsIlPIirfyiUyoXBmb8ijrhIC1fRZ7s3IXxm05MRvNQd7U83E2mebaFgqPRR623QYb
83F07eXx39T8GqOkISiA9uAGPTlUNCJH32Fs54BjWPlPXinq89fggGYfAIWXvvJAge5enjLZ7AQZ
3qzCwbzwVr3IOJrW5Q6z6+CQcDMBjEOGGz8svWdOfbHqMMBj53nkF9SIGHjXtzgGtwfTkG+kpj/6
h5s0jAqbyOL5hBNA6ty3/Izkc39NXZzF1KxwMgF89BXxGs7qblwF6onzv001s/5/GtDuewN2resL
2J0zk8biqf49bJQjACuq/4pWCnRBm0riWAdJvzdMOMWCO/FyAGYKCffgjTlzsNhLUpSdnDV0yIj/
YPXlkNyTtkNqRpLT8qnWHH9Afi79GdXsAQ/PnjMVwXYbYkS7KfNVTBCwdF/qhAvWrNNgyubAlKD9
Othz1ykbMrIdFLHphbJu+mLGv0jVPLhBgwSpFsh2Ppa0+vprAGUOwnBns62gqCuP506/REw8vIKm
cwJ4ElDCW/I4Pqu7tHVo3VktIbi5q7GYvcMrn4HK9+SC/h4uNQabQJ8hdYgQGptFAtYphfnUI+qd
KuUwYbZe7Pw9uXElgxr39u3LiOqmq3b3D0OfwwHhhSZfntWZGLCxPruhAxEWXsulesZ4LpqKLC4w
ymKXaq1HJtNxNG8hyqI2/Xrjic9oTRNfGL3I7pskKYOCQ+F58vaQL3L1ssfz9GL1vJD0MArbUjv8
2yx0YzV+Tkr03npoDV3XgnlZQVSDdiVE7gwl5fMANRRNlJyfXJrO1CR9/XOIAvCGSb5aA4KvOBUc
1hVfo5jCzlL4DgJGNtQAkeaRoq8O6R+xPwRyW3zxJ0ZejmjwRPETCZ3YlLQWib3WsvE/T5IN0wnG
T2srRrMRTR6Lk/EgzF+5hou/dliyETqlk2xTizDLW+Xa2bTtmNFVPeX/pInImV1wBlfGlk3nmhPX
Jc9HcMODCdTZr/UVbV1My3A5d4xx1x97siMZA2eN98m3Z3KnbN5C/523twWGJB6lAk42zhZAFC0t
6YBNTg8Yk3J7txJdFikq/KSR12PRP8KvTW+wsMglgYyhG2lMmMq5h4eS/mlYP5iYVOgROAQ9DV4i
6mGIdICHElB8iI/Gio1pdQ4zl3wBL3CWc8Zydx1Zo0SsmB4U21j3OZz8yUEw3p4efR0xsikvE/eA
nRclhbLKjgWote5iCbhNVvjRriFWYRwtgJ2dqipw/lx+MMrNo6ENew3rURantQoz6hxCT+64prcO
XRW686+bWys0Brsq7+oRpq5Evc/jrskXiz2wSCcOTx0X9+9cW8hkncHZP4STw7+l7M7OA+OD7Ewo
HvE6JgUDtvsgplifPO526hLw5a91azpioOp1wLDAtL+p33hb510VuecQyqsiWmmlg67GhD0AAbps
Ds1qbidlpNInLrizMfwK8H2o9pygfhu6AmhCPi6iRinXdDyE/vGeE1OqohMvifj82SmZiplAwSS1
1zmq+t+ed9/dmfiNmQqAkYRzO90wSwX8gCu5TyxlfpOCN+xLakkjOhY6TCdh9F6jOos8pJEEdRDj
uftygyguMxskD1ZHVVXDEHU1QOQm84Tdyt402FblINKfUPLDOIMIqpUdEP3pC92OWR6kl8oxD/aZ
zM07OsaeCEr8VVRmqI5AIO/sjKLutsGBGMvguBN0n147lA9Uo3HNjsFDmvh2WxKtBkWK8IU2oJrC
XpkwPXCMHGeFjmZtaq9Z1ai/kNxvtrLLHVh5HNopWUy0itSVT6xqvSPvvvecrxKkPsFXA3QOECqX
BtovGDd6g13XrjiQA93MtSewh5M35M8qqjclkIszbUY7DHk1Ab85OtX3ugnCJsbtgyT0ywuLKfJb
gDPsuahBI127oqRLuHwnmhd4/pcM76rGZo+7I/jf4NlGqztFybxnLD0vNDYS9cXTztaiakZp6M/P
+zrLWXKRbkKoMLG7odY7y+L0tgskVpWTOt84beeWwZABoGdTs98qFgroKu9nHl2ACjrbu1PvHpEv
6CdrEPtQHsYTbrsTp6ydLaby1ThSbxaEy0e2KIT53OBEiwijpKNNvH8qJwoHv4GECsEIZ0IwosSd
uP6XXvueR1sMAx0oeyRXpnt+8kHCPhC9BqFOMXFcONzF7Rt/1qdQejHLgGbDo93/lNOtQ1ToOfyH
1JrsfdPDnJafQmSk/9HmBIY2yieYhml3UviKFr14JhATJjNzmt1XwDsnbWrpd/H1XaCNrGeSsvHj
njTXSw+FgAIvYCDAFOlXexfPKesDsKUcP4wFrd/F08rPPfuTSB9BkG72RMDW0SUrusaTR9KdoZIu
vKyBHPrCzOhGKQu3Z/mpQpXDOiHLQkOE3pd2i2zKx/ZZLshZZH6UZ+/hKyVUqZgkUb7Dsu3eTsup
oiQHr1CWnHaA4ZkKskg3NUNdLqyDKipRUm2TW0OI2xjCX7by0NV4IgEWpi4xjMpllrk1lFtCEoLz
EzwdIzM5emL9e3a0Wh0xDQ17yTEYvWpfIHUmyXOlbb3g5tVmwdxC7oRAb5n2Oj9sSP0Pdw3andhj
1iLXFmOQjoFAECkCQOCxCnHgtdILqcqjPL7UoZiHhLCXqpJGZRp96mz2FiU3czvCpj9pL66tD+Ew
x58KaEz9OZEqjjIMpwFotKXuwJHozbE+Y/ViirQiqOlBi51/HRJwU1d0giBKMYyzX1B/mpNb/lEF
DgmxKyiv2kOYGc96578s7O9PhhLa6cpOEEXcofXYlhShs4ara7A0TpvWGKhi03iE0bOfg9+RkaqR
TB3P5tfEhmxQ6Q237fm4r+X62ryTiwEpQMA4jYUh/IOtzRXcet45V0Tb60e53sbOmaDV4j0cYzzV
hIBRCMFQsTuDnhFVkpat/+yn9sIfZCclBXKUs87KomtwKRR1/8p23Z25snwm5eoaARiE8V7l1EyR
qrbsI8mPha4qdZRH8DkGBeHqmLyz6s5kNfPxQAd/9AL8nE7r2uNC5wVHDrGN9j+8JPx3y6ns+0Ws
STFArurieL/58Am8F/di5RDnvrq4IdU3Sdl98DRUpU+JCwDRHhv2Ymev+93SjXZUkMRGeYEGCjz4
HTmMUNgiU02KqLG+pNsk568ZC+NwGGDdiQ+Lj9gJmiar5IuCWhSbeWerU2ewMEoKCGtP7uLnEboo
AibF+R0DoyUGyCTGCb+nbYILtkfMfO3cqHbF7bzeo/G8Jyao1YaTZf5T47P/SpibvXhwNZipkkbo
yfP2H/8twWoF1tOZmLf7fAbyN0ShstXieGYKV78xR+Vm6TkexHDgn5lcOeHYTSINt9n4/pxN9Xvt
0fbAgznkhvMAcLDyfGoTsxb+tSrfSxDmHwH5tkAZBTk2d9NFy/2EySZkHKZLIhuQt7LU6Q8Ou6fl
MDNdMbKIEjB/uReyXOgRogOgAbfkhRADHdlrZdnRofgM5Kde12sH0wRKDquHho7kzyJ9MSzJE4oJ
Fue73fuzLkWO641CZhCRvcYoSVlRIDki8Afvx6Uk4xg2HybNBjZpukGPVixhY/3TRj09vFRz3bX3
FCvxOoGr85HFM5PhoyRwPmKA8Zj/GW1GJMMT1JyIkMqTbd8eofOkATdJzrRm79ov4Fh/18UN5pqA
lacghCI9QiSu4QyAfZBIUGNx+iCx3fkcgrTMK14FkSbW8gnjVlHqNyJOfsZtxd6Gjceqaxz9/cHY
td1BsO7LXhqUl0km/roJz2wLiEf8iXvzsBa7j1bBCl3VfzaNITPJRl9fdKf8Pz2OedcsJctmaSed
KgJTyPtY+brt0EQ9MojdCuyGDAuwvaF2B3vkFOjy2XiXui1yTYrgnRtFlbYXKuTKIsBlRtE3dQwQ
9a+11C6nL6ko3fsP4yX9RbuAs6k8fvKUYxV8NIcA86CIqsxNr7ONM72wNXjbdzXTiYYAsY0fWnwa
K53OKigtKhmpCC75UkFwJyGRcYYERaiXWzx5llnzYVFUz0Aa8Odym/lui8TXXWRMOoBuNls9lsPu
Q1YUQgLT9fbxriCKKiQ7Z1ZoDEYko5uo2GuAYjg5NGDiB6bF4+H3oh68IuEjSKAkVx1C+cM2Tp0I
E9LtjVrMhl8KUOikbokebot7EsiY/k6szGKtlTFVQ1cpCAFCXWlEK5BDWIe8qY5T8cEKUjmtI538
GLsZOFUr3NXt1XFLOc8NGdMy2kJ5WFrUEmbX5PpBXyO6+C5JIJNT00sO9DKbT7CW5T81lYlvscTQ
Eyn9bp8yCfmCNclKe/kyJFu/mm+q90pc2P4hryCz24ICQicFgFdqoeOMaEORQDoJWRdf0GuvSfQd
1PjsgRW+H83h7+4fiLSDK7rMkuu1AcosZ9rteEMS9CR7lk9S6LwuNP06GjwnU60kN1CZlMm27dqw
ryI09pntv39aYzQciZeYji/+JBmCzZK6/yu+qlzno2lH6pKNXfoFS7Jwf3hcBpfDDhQJUvftQD9+
3labB0h8eA/Equ2V3zdjBznSdib7BDmNa5yQWcxFFO7QQ12s07+80TfggCqW9WBiTvhCUv4sEY2W
e+0EowFJXNJZ7meC4PVZykpJ2HS9ZGS3SQc4p8GwkqJXlSaQ8HmWawaXlS4gvx8HPCo+P34YkajY
LIdN8SjzfDoiMKqFVQmSRWxXiKbLbsDkZRoq76fb1Db2/XPiRF2gTvZoRF5poszQ+RdM6K0YtW4X
NdMMmwB9ChvI/H2PjdyWnyYaUeVDs7SDMt39n4n2oESTFp15/DwQLG9p7gm0e0N76bDcOErOTstm
Vk3+KM37U4qsGG+fEV6aP+eYIFctjJebNhvyQG2MtsHPjHKR39deqntxs4VevWd82ctluYDKX0hx
AO6ikowmYfxF2UVGZsc3XeHTdFfrjq2Ju4Qo+fpvBCMwmoY23JHvVu7CrwKZDBXUvP2uVDiOfC9t
BzBxvE2/ssyyBIGe08z+wDr+5X8QnwOzrvb3Q3a0SfVqMWiuH5HM2pSCoxDJ+H9xgbxLSlkZmyH5
ObZbcqRwbny8Xff/7cogbPR9ah5dQLx97T3Vhrm8Ab3ErdvJTGFJfI4774CS4gWCeET40qGe2Zkb
QP1zwcyfDuBrS00ZZQ4IoeU2CaZVFgk41d3Oh+C+4w49UWt/3qpSePD/D7mqzMuAQn7nFCX2iK8Z
otd4u79WjS1vcR6dFTemNlixQzAztkvRlKwXnWp2wVN5rUBnSpYd0xbhxKyqpMaHJDV3h8Qbubmg
M9pvX/zkF4ZqCcpNPC50ErxhWoAr7i0+JINz8LPp+BzZMdA1HeQ96tKmsk/x5n+hTvVBejRCST2s
KWvSKVKk2/WzAmfN04ecZFCwUJxSbTp+j0W6Rdfgr7OJq5bxJWG6FZYYdhIlbkuDL1Wd6mE53WkP
13fv/CQnNbCWTAjNbAYXx6Vt4a83mfMeudVAVVd6oRsRdDwb5+csvF7YxRPMaGbBCF8SZs10OLzx
NOjtduFvFKuV/sq8JYMUlcGbYz665AQxDei9JBl/VhiH6BjRN5N0EiAdLfFOci1QtOQTX6cPsqt/
aKGO4OzEyBjQgR5UNfg0ucX0GyT5eMRLy02LtEGxdqmrizks3wgvgsYKAakQ2JBaOJkbjRhS0QK+
SMJtIf2MOXfePfHnUyCV6Ej7gNAGAdV9NsPvx4X2TZbGj/ylNIPLxzN57Jw29kkdCz491lweeYaj
jG8tHmkYTCPdmqSELRsNbVmP0GPfQnUeiSd3KXzVyzchJNU8dM+d4JcZ3zzBlt8pCADxZ2MC/Owc
ZrWergqWYNzdtjuLP9FXpE8FZmHeQ50hSaV6cllYGqVmR9UM2crpRpw8cnlA8byM5W7v+tJMnPP/
LTXAhCT2BQh257l+8DAKC8xvy3hPASnveeuG2XEWJyfET0ClY8Z0m9Ft13Pw4qbD0XlzbSZCVxjC
TstD6g7yoeta84PaUjWeeyQcu7RkDilf5HVQgPn2jqmBRgrGDfVhJSXlXrmcoyFXAPnl93RmSdLA
6mQ3b8/6qZ0dWDSwgSlHgTiZt04NGQYZUMO5z/BhWAZJIjLi4giEvQ9nrTFcXzI6iEzmzUcWtuhb
ND1cz/P39Hl5bXD3556SxLGdJxq3V+Q8FzITLLiIgSQlPLNLfhSb/H5cVx0JH2jSwgvlg99tTlry
kGc+5BuDuKOoiN1SFZvFpxJXBi6eCnWBokjFf+Pb8zQ6+fGIKF6e+kKyLKiU3dSDYZldq+hQG7wn
ES9HfXInaRF3BhxJCcIbCu+qCfb57eoikynbRkdE0aI3pyM/xwDVUWGtYnFCFex/GctHjzg9NWju
cCenW98vM3/XK7YG4gxmON2c3HCfVtqQrUpneP89wWFWCY9O0cJbI0nuXXlY5G7JG4kxJUssesSs
gg7HgKFI3oTEAc6vpOznODTE6z3+1lx/uoGIKsvoz2hn0bgQ3AFdtphVEGSDknJZwOQdItaVfVGW
cewsFjJ3rRQI7vvA/3KnwXd7lI9naSgNpXHNSMOtQ4ZP4AuVGj6W29KhWxNTLikK5JKlyoGfhecS
pWfjBVS1Cg8HMALQJcX7bWiVx6oOsTGiQZMXbuDvuPmJ6bzDXhOUg0mPne7kiGpXOpc1NuoMCS3N
7piP9H4q41T9L+e2wRiDZ+ZAEXz9QnduLvu//i4quvpwS6zUh3xoilWbyHUxnT1+ztn+TiMjK25G
HhJrH5+MQkCe2snY5nO6dw6yFKRqwKpyhdX2e7L48yQ+j2+kx0RONdR2yU9b51WoD0tv6N8Gwj6m
HX8XoP9/f3GQMQkSos2ZMVelr+FGQdQ+gMYpK7N1pyfcmI6FOZqw8zgp5V471+NW4No9dX7DZWvW
qjwM96k5TWWfPms1IvrBKt4CLWwkVuE7ljrXxDzuitv7BGUBZrZEZAVIt942Poj/DYp2grqxWPBS
qRhWq39iQlVY4jgMPW4wVkoOZEHf66PkLzW001gw4wJ3Nodn+F+LCT6+h6HuAiou/NDrMBjjVgtc
8jP8QmYOYH2LvvPx112xP9bRB62CFGfAx5CIu5SAI2K5S5ABBUSJYiavwPE+KIc/vkRycbETGiV2
u4A2JliSvTXnyD0Nhyl8pgTto+UtqLeICqVyP4l2x4bU0qyLFLG/2anF1h59Q4mAWhkatJVb5gYl
+/7/TqYB0np0e9+adwcZebHhLj/Cb0r8hB5EwzIH9bH/pMDjzcYSyU6+5qYJrHDTNV+rL5+aCaZs
ZMzvSNgUzGxtOYqL9m8tr8jDyzdZxrM7n0aEUPpaV7o/hio/pEf8t6W2ePbbl+zZ0lnd9Z7+zPT6
+Y7HadN+ter+I6NVSOiTHGGDCRV6iVx4s3dHf/QibpFz6b0TPSMlWZREoP3dkKCbRzj8l0VkzXYG
cYziLdRGcU8Wgylk9kvK6p2zT0PXb2AzONaVYyM8zb0XYMUNE724/1t6U4vCVEf/Tsj+43eL0FFl
UHbCxVGWkFHk2GZgn7cAufgPFr8o0GCJOQRx7jYjNrOjIBoBjOeRb10WW4guy/SXz9VvKJLmNrxv
U3j5wT1tVBwkqqS3t9vDMby9iEyduUBTz7O7nNnp3ykLHxkF2mnkCxlMkjlDeTqKrCoERn8w+AuU
bnVZVl8x5J4Q5K50m1fwcQhxNartb46dfc97MduSGUQhQ6hEmrLaobw7HruOwu89GvXfrK9JJAe9
hGsmoYvz7ceskGMhlYaF4fo6uUNAtg2D9UBrb51/6ohFXIIt4c4DHJFmDBSkYAck0WJTP4a+nno0
2KJ8NWPLyxUW21UjrInj5ahdKR2f0V2JK/9CcyeHe0zEW1KjqfdXdeGqkGjAVollp60u3AvekGd+
w2RyK2i9XakzPiQncpYU5QJsvzy2IRky+Qv+WcBqutEznOBZgMbORA/4TBj3ETWDINhT8SvyHgmg
BZQVB6rsvszzITihIuQN1MhcZhzAuW5EhlBQ3JDOT/G9lZdmOADmzXrCKvgkzKvDYXminPXGath1
4pccNAmhlTOXHebUlQuWU9TxvonGFTQFx1Nnob2vCPTFb9QRXfWLmzw1VaYdQ5ILxCnsy9lnIJpt
tEbO0bSYfjYoeGSjNrqKwT77KAU4Gr3g4Jv1Rq7G61W39nBHh1RS7AL8iop491n1DCTyzn7y1Wjk
Ju0RHqrJ7V7/tbq9SWQYYjUUztN9wfNQfMA1xMk8elYdDFtsFwYxNnl70c2QWtNZsmJRPRmoQ9DE
N8PWUNtM0kcXLYl1uUu/HAiXHzkxkXsbkoHfjTR2mb5ogGbc4bvklxMtItqR+djbk5WiNRUd2WPa
7osQw15V8lUW5CFSdAndWnCwtDvdc5/Z3sjJVU5u6BEhcflei09x0vO+UKO6lS0FBqv6sIj6cx8l
VB5K4zVMr2hfaQtfrS3FnbM1JY+8bVTiFTCJfQxk1sdtH1dtVQMQBpKVDXc9AQTqJ7uCUKtCN5HO
HZqOqpWFw05GvRvXkmaTB5g3bti3JrBioQYjfS1zsYXzlCXZpyeQpCeKv+i0yoQItmCKkoIaMTDN
0wYGMdnWZMhl4dTXOuHka67wP0q7pXcq7JTfLqK0JyUc0bVqd5r5JvFBrziM5K71qlTY1ckH0Lpt
Uizd19bCfy5dc7rSYSrmx+SsB1U95vIHjkV2ffo7wZbBRLczhx1RtnfJB+zPdpUB5F46mkUCsTMS
QvJOt1AmHlckF9hBMiNeghwxdXeNHDwP0hQIjXrlRZbmkjaeGPvFM9BFTvb1IfixkFPMQeDZtgKx
lIgI68vlY1K+UhwC7OSAyT/f4Ww7YUBZCEDYdKtac/GK1/2uBVMlGQ9mFionJmlyJYcloJ5wXKKf
h3FxGUKZ10+3TpJQU4hhXt9oeyasIqxWm0kAgLD8mHtvSoBKGom476xYzi96K/nzwhGl1VuiKass
VsS4WMo9NU1gnsmujLQjoZjl7a5mEhh0y39EKM11Mk1FpKiLSrphhgf61mysjM+7j5CX5VI3Wdjl
+oN+ofSu0GNHwLXdP6qBb181cTlUH91cGg5SpLregTyDQyTZy94DStQdrpLaUZ6ZB484xUATlMyp
hL+qrh2leTI98I30aVuLu2yMD9bzPpFAgNroWEbIUfV6D48oRxWBupT4VkF4f3mOu9OtrZzBVNBM
CbFqqZBtme6jJ5N2O3JvQ/yKvXk3Jm/Fm9+E1vK3B6sRqEQGZLXG2KRl9OPLtoKsnwwbYLNgIbuu
YsDCOdiw2IMlN2YHBDGvtYgu2PdyHyRCJFkmtZzbWQywra1kGkvim/P+vbZHmLjYEoXY+p+fohVF
1nnkN4SI8BuCyRZzjAI00NUqrND7FPeYzvcgvKSLCCfor/MpF+7YRQPdmQXt6IvetdJYP/UMgIKk
tj/Cw+phW/mlFQi+TZrOi4yvjOBX1cTpUNHf6/OsZkJLdw0GSkkyDO2i/GekR9mi9Is4EQ/fRYnP
i3VkBZMSBZaTdE8/4nv40NAlYAP0d89jyLeemleRP37uyPbVKtzTU4i1FyVz3uK0fEnjkcQOFVbD
BxBTiuwjwyUfKuAEW4GviveAXMoqm3DskvJ2TgOnflonXVnOdZ0S1RJ/QBj6RvT0mDZalniE9y42
wNfs6haRSADi+3kLiBFlU8QHgN2dA0OB5IKuqbaceC7l3XSbWh+7u+BVPLuxlA1vCWZxZnJo4GsL
qhE5XGsnUP0iJgAlFoSWx+4bTk7+om/qB1sOtWEfxPiy1oZuu9TEdIYKi4Il8lzeHJypT4hbzQzS
EJcpRkfQn52tKywt8vdFaV3ZglmCBWmWDIDw2YNYYql14awE0mHs5q9qDQtDVo1ILSb4P0SEIqXY
Te4QZadJBTqjsWqmwcnLRd2O8gMbvLQppgPUIWLgGlXlPakLy5oTIsHst47JDt4bL7cxb0U3ZcjY
BuuIfxtzUeG2HnPeqhmRYmF2tp6SjQ6UV/IMDytzSo4Q0I5f8rFUt+tYdEF36rMH2bvxmygBx8EL
+4Zgh4vZNSA9r8MAkiYrXa8adBgDwTU7VBSPA3D7VErUKDeRFjniR0BdDwVdNYBU5soLo8rNrHN4
9rOsTAjKM43xw6UvTWosFQnOoWK+kvx9Mmm1QsHQ2q1IDjNj/E1ApyfHI3zTREBW45W7wLIO0yV/
tbGYFjECUjasKx3B0tAMPqMR5AUTY7uUaq/86Fsdkj3TlrJ+CwbT2xKOAo5bjhQOnkSpWFIN9gO6
VXj9VvWQ47Cgc+g70Wo2H494adoNlVFPMs+9MC+4qWn2EmqSXhxNGlFuFClk8snqP4IoxpCHBVKu
rtWKIXnYekjdLkeVxC/phBlAJRA7Ob92xi7AFXIGk3OuWBICoBBJ5tAaSbIx0/9vQpLCGWcQPRVN
87JVqksOvtMLwZGKoGMqDPw3T6HjQy6KhninlOm90PQxu5birruQYJS2uTFnIvwYVRVvxSOC+dSG
H2gTrG2u9YomVU1Ou63rhIMlGy+eIzU5KdDiGfBDU/mMe+KCTdyeTsKkHjFDDVwZ6nn1IzeqmF+7
cnNQjJKWVAeGW1S4fcSiI68m7AEn3ElZlf8o2Bm5MaYh0zJ7XS3Ze/IYOudRGTvN6f6COSiuW5JR
2plgg4QCQzh8HA3UTixprjIkcp35HPqjjVojz0eBwoECTZQx5vKSu+Obr8VLdSDRqVlI09TzlBwH
UqFAeXo1AHD1yfbFsDg3roZXMTh7or2CXcqCXn+nEUXdkDQHcZhmtcD9lTP45PLhlgRaUS+W8yXa
esPPiT0Io1BL36JLlfMw4JKnKZqbLsHWG5qkuPDa5jLeJnVCBHbD4VML8tPtjlpEB7YkvtVaExw0
buZPFiAZgOnssJG/v6UdAhLIQq79zKVA+NcvEmJ5vODnmGRp9Ow2HCNeTtwEGd6gWa3PlN54nY/N
Lx49VKuV3soZhnBMc173m/CEisF6cybwzsRzOp2Jbhv24t+lFlS6fL3etmrRPs4uoIxG9SyDwLcz
DLiGuciKkVP6kldpUCXJhh9hFIfZ6O18iqS2saQagpaH2ZaMgIxpcnFTSnijbiZ9MxePmFNxnrEu
14I3t2XeV84AIaZLIXoBI1ZU8aERFvOQpIlRxHEdGxvRJbKYQFKSQbEE1SWtRPJnuTozwx0bKAF5
Ba7sCu+5PafmNiNRJ41S8f8e3EKHNwSMATHiP9ySG3a8CzuXEJnBqITcpHAvIBHYyCjQv21+1qNB
1LAD555b12tSIJZ/CuXuka+Iww5ZzGv3D8cXBpAFoPBePhQjCjlbq3XrWVB3aBg+zqysJlXdYKN6
6PJQoYCi2HolKBV1FZ5VqjhrlfhCg8SZP3Vn4n1yLMIKZEAnHis+7x5CqyKsflAwGCWZ4hkmhTeB
ZkvcGWIx9KFYLPrWHQSjK49+tNUpZu4FrZbJoVh9nu7wV+yIAIcWu9u86ZeSLrk3Rc+Wvu1uY6id
HBKBpuE3dEwzrPcfWfIe9xEFq0f0f0ZYGBOEH/dtRmeHR9MKyX4jc3C5yvLMPcOwX4uQq+dz/z8Q
+U2PVq6Hlsf8XGfWcV4/BbVILR0y1nbwl6XgXYALh2vRLRpxS6NjrUitLXhph0WVBf8jL/66cYkf
Ts4bBNYgsUZi21LCyPBxt466XLJWAraDK1veq6KUZf4CSFNdGquVQvQeGtULixoLxJXyt6/PfXd/
oCaCTgkA7R1jBP4OPj6nCMGmm7uSOZdsi50IBInMlrznckBlvxm9FgSrDoC4pfh4NuJkAEgfvakg
kRDPNwVVnGu8O0h4byNVSga5SJt2KlPkSu/Wbn9tMW1tbXHjh2oSRH/apaDCvuHnsbTpV+3tLtz9
bI/L65mVOf2+0/C8DBh7m6o+v/9NLl1ZRtKX5oIqPdC8xXGmOVrF5cWA2H0P7KPhIdHRZyEVM5Wg
41Fb9zXnDX4wZz0Tl80cCCRlZJyPXonjkvhidU6/VZGeVU2Pu3oeS3jVvJlEZLygxfmlvDKUUY61
DTsD4V4hHuge5Cc9sNe7CcLxDKX8U23T2JZ9zZEjv41A3BZhfEVPiSKvu9z8lKGJHW30pdo4qLie
bY7HShTcXYhf28yCKCnZY+0zCQI5/5yqgdlz446jqm2boJ3RIxkvNmrSbwWMk/ExJ0nmLj+X7qqp
AFicKR8XeSw9sNgert42DDDqOIgtsG6lKJs+u7XW/1q2wniHVTdTpbzIKzMbGpVZz0hIXY3knW7s
2XrVbCM4qkzQjAstj6aTC/ZK9KfN45r7FubEeGpHpsm64Z1stWlh2yZ+RCgUieiNSLXijpcM9nuU
4sBxtKWpDAFMbw0ALjenAZzknh3XRRqZVqtskq+uR11FJPKRTdDfxkv4ieEXRN+9XGI7T/S083SL
tV4PpYRJdAyfbpjHSw5cqk1igrbY/YcTUT0AHSjWoQFXDu/yCDpCTGxiseYuAM+VJJvvMtBcv3ts
Sq69pibJJZW4DUuL/fmM0mY+4tCxzo8tEy3I8DGo1XKLTkniqGMRH4GbuoxImkKbPr8vO5pz2mYg
5/WDqtl96lTO36iz4LyP3sWzcLdqVMZwDDkIVoZbcZcnYDJIO+rshTTgKGGI5aeLQWu+IO/QQBZ9
QABniB1LIoHzKsN8ducrd6UhSEhYoCkObObNWkltr+CK2fxociPO1qhjOi6YgdV/M4i9ftLWC3id
0vATEv0zgZgrQH51bTmwApf07YleVQoUqto+PR9uWp6ZoBROtyfoz8V+6Bt51esiEWRtJ/u4ScEt
XKjy6ez5Yrip6cIcVgJS15u9kJQ21/R1VGJEXN4cOBPOKJmqchB6E3YBWBpiOpju1jVwKTayYsFs
tjv5+Y+EOR2z9mal15BSsrF4OF6szC8risbt6TfyfhkucCX5+Ffxqp78qYAzu2rVZzHflF9bOnfl
z9BfJAENk2n1IVzWuqnJ1IOLnTmlc4m5Y3uP667TsH0ECx+osP/a03FF809oGwADj6AhP4QDrXBx
rwFOVwKJFvUZc4gK0n00ncWsY91QbXkd5gYHHSYTiQtDr6wpkaa9SNu7U+YE8zO5up2BYr3T/s2e
58l3MLyWxgpJHpL4EruqWWKqp++6fYUGnNpu7JqTtbYwDv3PULAgJFLo6pNIbl5CUgVON7ms3z/B
3j7Xg8AmLfxs+V8gvhUdMwJq7pGCOj/88gdmsb9HDa6dtvmxwxBsAL1d7CHi4q3dYHVOWBl2irul
wpsNBVvObonlKscKb+iOsTRUn5rtxVXAF1n5NIddTHF2T6eWIcpbUfqFrwIYJSNuV/CGWaRgzDTz
ZSeQl9kxFU6OmQDhOyd8lYzonmQ4nDBsrvm68JqmGNB8TekEPR9oeY9z9X82DpXb/WbdvlvbiujZ
yeiagxGzHlOwWL6+kPho0YopgJ1lgBFAyd8DOLXpTtV1EBoRAailqjf/9oUxhn7I3kJAMWqw0eWg
OsTs7qi8531nQDbMn/AmQ2W56PQIpByUvcmLN6caF3TC3iVoghbMAQED+vDCSAPgq3QRxKou9JrL
g2y2gTL2thtQBGwXVGo8UDGykHnnUVo+jMmniLciieu5ntpMn1OZ/q/gI3rALdU0slZm/zGOU3Tn
oj8U0zlDtlMwbHX/b1prsoL1PzeAaLEWot60KLdUYSQpiuHFh7MtcEysK/enCz/lXeypNTY5q3rZ
9Fued8zV1to3VRW1vAZQxyljCcqLQDCekl71STzqReNb1Knie0Ek8RL2wRCoeVREkFxayF0aWiRd
TgXmaoQeYUbD+aN3NdjzAmjAJie3jZKNx8bR7Sv607oD4wbUncp9R081msf1W6Ogz2h1050sYWYn
E+nGHvNeomCQK5w5qn3IUupE677DRp38CfR6U4b/VxYtNCvgNZ3WiMMo9XZMcBN8rEHPsLFeQ138
YRwLVZGmw/uKG9p9Vib5KqEe+HiM/75+Otd6HCsGk5tHKNRQrLyBggyeNjfCePS6xVd8BpvKxiWK
/0kEOgNlzuTsXA3MRd1MqtSiJft3/oWPGij8nosN4B/0K8w1nOF3/fs+UycYmb+h3268+pns/cYo
piZG+XnrrE9nuxu0totZxo/ezXATesX5K8BQPe2KevpnFm+/3cbscVKaQrJOfmLPC71fb7tTubhd
9b/JiZiGnEzRVNQ3wQtvwaW+8zfJM2Wm4tneeWglyhueKlXdjFAebPt5wuSHXRm0pZqVJ25syoul
oXQ+nrD/AGtww8EgCcmrfNGZPbM2hizfI706DFURG+sXruHg4RwPFAoYAWizcXJ9gdNTx1fxQKMe
KKacLnz4Km13nmu+a87SBi6gv/inkia9N8+rHzcR0HIp7TUBw+j9V1AI6aw0yu4VcGTaXPIUEZoQ
scZK/s7+rgPBavoOnmov1flS5RCIU0au5gq0lVX2cUUExNh/L6qx31StI/mnsT7BI61SFG+rdSFi
oH2Gq8PbmgxfTND1G3cn6K+jBGxh7r13ohG2wRGxhIJsWMbPbbhX7P0wH3gwm1TcUDzUhV5I5EGq
/Kg6tUt7pErG7+p4QK7uMnNLZ0Is7syxKgJnDW7MBEJHWr5H/mv817N9C3cJhG9u/xIODW0nWsuO
j7AhqCbuage+7klMgwwBOHrT4mp3WyfA52vL7sdNNKcVP8C8q5cNwrqyUsKnVyxjYEU1wgE/R6BC
AdF4Wf1RRHVBF5HQErJDtTs7ASJXDrbMzDircSB6bDNnVrfdHryJwG4Fx0CB0MjiYtJKxUYB1HIy
4F2PfoYuK9aWY+wLVcV55bXqcXD2ZrEPZxoOKYzRZV/u8X5ZmBKJhThJWusFs7RVWYA6Nc2x6Dhb
eAw50I+1qJD22yvwjExUpPcjgsJIm+khBc/t5x4p32KjAVZkgDdiJ8q6p+OylGHTWQ/MR6cg3Cke
xgfwE2ifL0oGJKxEcLzehL6lVGYMY8LdSICTMTD+gKUIQ40kNCWN4LUKm1zo+kbtkmx66A3eWKiE
h0u5/7t+rDxjkW6DdUhZaFpNff8DBmwKDfgI9j0stYV78saUXniGARg5sXNvKl6zijtM4YPKy6/I
s36sXdcomfR/39XR2WobPogtVNgSrkWLv9ud21HnO0TJT5Bk1EN3KAnCM4/2dD6393UsBapNhMbz
G8UadwGz1eQ5dFh/hTBfN0syeSaKepj8F+avpdGaDxi2ZMjFQG0jarqKI3im2Db1oxjU9q6qQNy6
d4jFXUgA39VUJzDOOD2JUPeaOkCHsUiNOh7FCUPaWCpsncr+p9Jk7w323qG3gXkB7PlV+PIkCaDv
0TLTD/hXrahuWAPcKcpDpmM9hjcVSvEQOF/W/ZO3UMcFZw1PxLqiX45jHBfzBEN81Y0gxDSEv/Da
06AKrpWvYs/HRkfCq+9okZoV+hGD2GaWmigmp6ilgESqrkFqt4yYUm2jMGXb9GVF4Sr27dsZGN/y
Kl+gb76x2YwHmhu+XrP2+pH6a5Xksm71E8yvUdzvPwJsDygoFh1voMMwIbjb7m+HBNN0lLVcix3+
Ep+99YMOV975GstedprTfqImr9B/xX75+zbb/uMp9e29nBsXaOfLuUQVNoYPQqvabV1SeOCmAEqm
1NjNCpf4NzusGD65jJXZEd+FP9wNNmHwDAe2p6wuqq2noOstfc3wlDKwBK3a6kx79OprGRvNYFVH
2dVvAC0Nyx87HOEx47FZD94u4dx44EU69aFY7iMdkuY9QFUgEVUDgH/8QGRj20ucbrZLP/BuGgPj
dDG15siLwTtLPv353DXUOuxbGIhpFDE6vQW4eavss3YjKeq6TuhaMyeThMgwnRbSwCztUczVMos9
JAVCdImRtzpAtAOdUvqMUxQIInY919M0Z0IWwW0WHEGEX78t0LMi/DY7gnyLzq15AsYDpxLG6Pgf
T3TJFEggSqA1PTeTqsxVwum8m/Ni4urQAIBZAJlObbVp+RBSrEKMQjYkh/e+qf+De4Y9giHUlm+Z
oFEY4qSVuNcOy5T1AiVIZhYmoIT2gwHek0VE2SouVMSxUENnt1g16G3E65is6p9FgPblGKI9AGVs
2VUn+v2MdJNKczbCiDGlz584oR4Le0e0xKxThCOWjc4zY2weL+S2NLk+KxUi1XGl/EyYZEE57l4N
y17uyBbz+jhtKWKEqtw19GHfBtIwdDovyC91soRrxQfFRaOiAoakid6GdaTXXDMSohQztimW299N
mG9D+lQTn7GqbiR/rKJJMBre2OKBSsxz3+yFhpMUXsM4K8p51+bFNqnEFeQ3sM5SiNlP0BAI7vCm
LpWoJvFq0RBdcmDo9DwBuInxSxCxiQcC2iwE2H4EyQ7RBlkB9nxa4Kq0+dAC+PGIu5JMxFqsUkrf
EBTQoz9gEvnHJisKGqrE7qG7+7xA9hwdrfr8I2RR/yCS+CzfChnbeAacKGTB1GZn54Nlo9Du3Eeu
neBTdYFyIaTydElOwQy4H0ejfEM2sKDLs9F1enF0JiYFH+usV6aGWT7TZ7ugtzU+oaukDq/pM1k5
tltrpIRlInx0T5KuIHArvK5p65PWsIWIkNQfE+RSj/oRLujNxADZnQkxLS9TYcZYyg2TE0uyjFwg
y7SfjyjBiJ5N8BrGfjdPfx2wEyqeW0FOw4v0li4pt8daxfqTWKaoBtr0E0BKmJH4xl/Lwo4G7pTx
GHps8EqMvzsxRRHMm/Aldhu8Vpg4LJQE6B4XMBo0wgj/vQoY14tIz+scy+uOLhqNJwiSJBK/Qqw5
iDZxAjRuyuGJdzxFMebjyFAGz+4IFMN4QuN2BWhMdWVCh2Ri7aX6LjH4LJKo7xpI7ZOql106FacK
JRR2v1xommQepPUgWFI8+qKBnEwv8KGwdMh39xh1hACSNjdr00/EvYQSEB41SXbNVpdTx+wM0K7L
iYBPfIkfDi5d70y+D4J8QAevnQI6pxY/BPGX2LDeM2+5PcgZaSK6A/+xl0+U9/tdq4wNhFyB/Q3a
KexHq3K5SewMUiqdQ2PLjfskP6EJ7lABXFMKcUILKJZnHGsNFbuwYMp+GlEWiYPN9rJtbWoRTIyE
b9MoEeOm8rcUrCVuA+idM4+P/FNilvOOSzZXO+WrRwwpogtdtqDPLqSTkZjL9f+ah2BNGSGeXWdu
/ZyOLQdRvTNEJcpaqwh063bdcdjHclOl4j6zTAZ8Y0F6Mg6xIcNxIybOOwWVjnYP+oURcIwNiq2N
6pVvK/Ripyz/0SlnPS5gfIrAu65+zhAU0XykKgXs8uDiYaW1iu8uYc1YzelQvv6mY67CKgG32cVo
rc+vUQMh3TDb7UoTgqo8rvB3YICWIT2UH8hM+el75RNDLb5aVsidE8Xe3Lfq0xE3m1OOhMloQ8So
d0d0e6/9TgCHlmUEtMrZHG5TTo6oYdNjf4iLGJboge+R2+V2m+Uw+/iwi+r1nqsZmgBymXPgNlf5
A4OHgzc7D0aYs23Pzg+7J2ar28F7y6xG0Eif17Q1yZPup92u4+U/tyzkVSZbiRRCQMoW9fSSTWdA
jEP/Ew8bYDPBjyTBxd63FaqNHdeGXqxtIq9UxkC+YgWUuEBE34W5ZV65H7mwA1BTJVYsrrfiGow0
TabAXqjXMmWtKyUe+XHYx92PSDVTummOymxOfzy7px+3s0HF/9zL2jSnmko+fQroX6RvSi/S/hkf
xJeKo7g14KJA+ncB5HLLWfBSsTHbpXxIlwuhYFwefkxVG9QkAxfPFNZigampyz6GIrkGgjXG7Zvw
uoKcxsD9cCNubiTwHw0oGXT9Bmd9Q+qSUxmYygU/DCdb/kRInSWDZHsng5wDkkjCIhMdrtXWcXxg
JI0VRGvPcJ09DYuSw5C17q96WA+73y7ncdrkdra9l2uRsJO6LmwpoJiiH96xI6hVJUP5tDZ1HJvL
UyJr68i6tn4j40XDnv/wzcTyKOdwwbmFCKMqBqWIWZK1zwgfnb7SwR8YZixULCUhRYCfeLx10lfw
CizBq7IZ855eiUIVw6f5+JfVrh3c60ODptEvceaji4z9aynKcbKmW7sNwk+D/6shvsJkQvNR5yXd
8uWf3JNNuqlaJTZhpqL3T8moz74le0KUyPb1Q3qk7oaJrBidK+MGLKrqjho9eSRRK+KRIaw8fkKJ
wIPX6LaX/WS0shSmXIwaO72hzwQxtwyRG0so6XDwbtQFCvNaYsNsjzpdfHDESiAVbsgojC43DBbT
PumFVBDSgSBAKSJ5lmJbcqJgypPlEdsuLl2T5Hc0vuNvtArwwy52IPVzqK5bZevAI0WDWOXsw+EM
Wh6x2fRZl6wzGBr0iQNTkZr9oy3852Y7kkJ8OK6g8kjSyyKUVhouuSh9X9UWtz8I3Ar5LdiceIH+
hEewuGB59HZblJt3uYKcBoj9Vkb8sK746qIr2OM6/s65AkTb9KJTfMXBA+lyQKYaDlT54fE/Zdof
CswSSTV9SAFqoSb8U5mFl49erczaSgntePsVldSUV700SYPYjuCL/LyxtFIjPQVzyDq9VhbHn33y
ZKLlU4jUwYFmkZMZDB7IwwdK5ZwePCS9Pbl1E/QSwONUzbvMNlBXdf8J4R5pyDGYEQ9sV+2VipMU
Uf0ny9EHUOyY24MPHpj0zrp4IOEYF81zKhQG60GmE2TIvfScwNb2lkEkhOvmm2UYq3wqswhZf+uj
dFsQ1H/sQ/KWXxDN3kQ7OFhuQ3VT+bT1rOVIwHszl3WxVoKy0SXF9Y/KAUtVPa8pn1V9QPfcjjyZ
PcoCVo/Q3zYQy3F3pIyknSBjNO1CEzhBV6q75VDeFaDjMvopT4V/x1qIUpWZlHSa0hMJloIjPduc
RuRL1pPTLXDeFbPzsQsih8P1mmgDlR8lZ0UbuzaWV/TG/yuwrViPUU/vXguJz98969KOq4WY1pYE
yXsQoItIix/9Dj4jZ9TmmvC1SCGnDaOFw1LKhMjxL0uBcn5gsCw9fmnmUnq5TOmXyUCh4r7MEs34
HjG1DpdapNE8OJV91ioBRcm66tpHPKcIsZZBMT1fBw3Dpp6yms2H0vMEBor+q0oVte3riXFy9h91
BJ5SRUHwMP5OWPsR+QRl0s3YC/C21qDWcZrS02rrXyI4f6+u9T7PAjJm+IMAT7fiKoEV1Ot8RGyq
WSOmxeVvyQXzuSdgUrqxHGdpIdcXc+DVqlYUx0Ff/TgLZBfUIwenHNhv4XW4Yv2W4mCQbcLgFbuw
Y/J69zuwoOrJLyVVb9Xdx7TatCaI8vwsWnsyrGQoWfxSSlDDw1VHEJGxHj0UdgUsiZsmDeFHt2hm
nB+ONUJCQPJq5YLR59g0iPC4nIvN3S7xkVsqq2YEFGOGhCPMemo/y3aJZvK544VY9b852xjEcmGM
PRCc3ZdjJk7oBaiqVfbhbv7T5J/Cb6unce4+JPlEUZ+1ONysTdhqtzt97hK+hXs86PGyvxqjKnKI
lbeJMRn7p2vF0w+J4jXmuUTwlBxUyxREZrCpCtF5puuxfcQvMv6UyHFJIQOIx+C3RggN0KNbOYWg
xQXhl3mRBx1N2jWvzjFElcTZgfpoCr7vurZPIYfY3yGK/9rtU1A8t9z6MXy8M70mToTVfIAPFFL0
0X4Pv7sRr20qeQgHw6BmiHy470yJq55CyDFmq57nAdV9d24UuTPMoGuvf5Qy/UQTSKTlv1dqHa6C
GIbKiKTfe+sRyAZgUX+zqd01urjpKMtk5lhFNBHCNTWQLYwJMciaXk049nEWjrIZ3Ue8U8x2DiYt
0rSUhZQF8aIyK5AYlABmMrpxpSFOfesPIm62ESCGHK1LQC8fsp9sSUaUEfkMPj5dSJnS9O8mYJhK
wTrHI01PUlAjgtCNBMP0/O8RrpLppsOVTZbG6wZAz+bSPloLHnaM2vj7ZIT9NLjsgR4pcHFDTvG6
jjVzrbhREmO4PQW7POE0kZWTuPqvCn0cCxgW6CNpHRu9sQOFGwnEZ05X+FcTI9Pkw9xAMUpGifMK
WsktCmhVA7rmDUdMzcvNFBeGFlD2Xu3Qynv/SKAmZi0BGWxliorcMjwAoeIaONbaSXBDgbwabvq7
rxNh0xAdXrEKD50cTxI4cHpLXl0qvCRNfB3Js0MW0lgygIGmojGydMlRxcibM7FaCCZyAXzLSGfl
NiDRIIZ3B8fQLsA4cNaCB58Y67YyTBytcb7XYJfmKY1jh2r7ASwNKui2YN3EMQubxOtvw51aK3lD
7Vk9LbWv2J4SaOZ/FQ1jvrA9IhJERrxQf5R+Fhnbs+u8mCA07p57uEeSMDXIMn8Q65AWU7rZzwX+
UL1IcJBXkNo4MXk+7XIUG5LnIrtd+AVhhgoLRXRQEimonFmi4KcAUx9IW7EPYRftgRqDBQCAGaxX
eZTrkeyUH4DsqjlxvK+Yr6WLiwUWT/ptuzn2h84m/Ux8xIJJTJpp4HONtVGUFKqeXIy/ybkn8GPH
v0Z/Rymo10FQtj3oy2upIqB6uYYrjN+aV6xe4WA6kF/zopvUxFkVncVhjmZaapWPRrCl6GoWrTlg
NIZBjNQdFSCDxhQHlIYyhCvf6mDclo/aLG0Cau17U5H8u6HC/lZbCpwT0pES/SfcLPrIRzNW7g76
+XcQzL7a0H9WqYMYydWY+VQ8U/y6b5TrmsiKnisY86AsDPGHVdNrGrsLVKG1s8h3ai6++0fXxqXS
OvUeJ3mM+99eKRUmRjRz2/tYV23rDhCqTFDGsn+K2lmnTwTVEYdKss8Po+p1tydoRYnmhfrQQ9Qh
R6dn3cqIaM7nGbHkFkUs3IIH84p+Xc80/3gQXJlOYF+EVoDOGs+605Y3d4NcMaoJ4NPXJfrUfpH4
FsdvAgUEd9SxkiWYPpWVnzqxVdZFtJlt6hNbq5H3xUjXC0KEfWM0nrfS0YqY+OvRKWfzVB3IzYU0
m9CNC1zhUy8TWPoKxUIGiM+T4Ep4wrYcbcCg1psclEysRVgfeJXZite6qNpgCEyVJJsXItlqcuBT
G3gyq1hESsMr4iAXP9oM+9pHXhP7TDlbZNnv20ztSsLe26RJDN/rCbbNwd4jqCCATcYx9vG4txdd
Kq/8kahpCMXrpy0gCOcyYaW2DJnLdgLo78ajHmFxOhwm92JhAc0W8obPfCMpR2tlCUTuOl1mRdpN
n3PLSy25lFwP0I2gVFLlthldvPaayFo+esthhucuUk05H5otFqGvzuBK29pwEYWo3ALf0Nr+qcKf
DmtMovBB0bHxAc6ez2VSpuBHaN9cN5EP8kgWfM+84POXnxoS0cc9yCqhyY/pLwzMqim/0Es7GNta
KffvilmcSxJLSCSOdEsoHTvO4JF19CQh7id1ehT7BNew1pqfMbJa36iWvgdZ/PwFt2TcYxepW5s9
3YmZ8tPSplzNVRzGCOrFbCjcl1N5fVX+8sG82K0zv8HDL0AVGtkT08z+2wv/o/xSpb5i9K9QPHLy
GKMYC4gpNb6wXedlzW1VVEd4pf1txdRQVvssTqPW/DfvEAwgo4Fly7mC81dRL84bVoRelbmrsPf/
rofHi0+0i51+LG2U4hhQL6B9/pYxai/9R+nwywN+PiVFFOpzCyVF0yPAcYc7vTMNWqSIebQGe1Yv
tgCiVXJd0H2cbch/TMxl6gy9r9FLn4KiLOtLr2yffnKXk/2r19goX1iXmudabjNmFCVzGvgUHpfa
wDI/c6XwNWqjI4UqpXzG1paG+BMXQlXB5wOok9UGbVOLg9D/tdxuB7Vb/wysT69u/e7kpI9Xzah+
7bNb+F6mTZPtaFx2dooQDiHnT5DNnjEqYLScPoxdj66YDk8noD+9pwelCpKcmtTa9FWi2EeRjxXZ
9qH+AvVsh+UhCZ+ZQIeqv5V0h2TtqOaTFx5p0HYiN/f9RdqsTYsy6zQdTAly7n4ipYDQvZ5ANsSh
b4DVUt8Io434wN5fioZz53Tn3ozFX5DkrO27xvFLRdil92rgsUUB/5tpL3+CnFgetoB3BZty1p5j
+P0WEWUPv067gw82ZjtbwE0g8YSc9zLu379qzQFPFIb+r+1cOc7qfJzRV6tnTmpJE64pk0idMq7R
4eQ3vz0NLesDhDI5h1exOYsM4ct33vRS/986o5ypH1oR8tVsNUJagzlvETDa5ke07n2tLf6LG4un
9jYKnNZnP5yp2v9Hm6G7KK+sb6yLXIZKwUI7jbh1aL6FuC0WUAlU00TsdNrPuXU5nXw89HT7ocn6
z5/dsFSYjvNUjadNPqBlAEEGiPn6Zf/qJMlcbhqg4XtZWOwHA4IlLX1X45SZp7es4JwGFP2gd5pJ
Hf01qjnobx21yx3wmh4Om69D8dY6F93QYpwLGDvzM5wEuH1e0VhpDA0WvMOoikQxWNGjVOt3N5iZ
TSmT8CdEn7tAcNJMkfS/GVFGu9+yRvokDpiE38XzUQBQw4YB3Z+BYkfQ0MXc2rwikWZU0mkradYv
fBOneVB9nrcd6pgbIq2OKgKqVQu8ZcbeEUwepfsu8CRq9TkEp3Q0F9MoMiSfY7GLWIx99P+5Du9C
wHVbJT7a6hstbVTJDx+HWxMtIpO1o86/YZtADLGip7zLXtyCZ2LaEh2NywHmroU6dXMhSxPKID3u
cq+VK7jme/eup9OWhomMjkkl806HG8H+v0bAQdslXLKMctA44tqU0CuQ6U3wbttlGWaARCt/TY00
C5z6b/K4cbyStwZFCwf6Zr4L3tjFtj6ZUvP6w++rrrNxVx0OdLIxHHrxcvHW2BauTAUyguUKuV8g
fSDQBe4S+Jk8vwYL18T87ha4zB9Azh9dhwmbgoxP18tvH2rV/HALSxxd/D1uJMI3rneiot3xR6AK
LW4P3HwSqssdjosM1NM4uoz19iYW1843Kfy0V03eAPtB8YeJMAeIt12Ti22cg7lehxlRPw6ibtth
OPjeWAif+msDGCteOTyDxG+a10reYcp9/8E9A8OswHp18n65rU3rWfzsguXxNmPsZxbjwDgw7rqS
F8ADyobBSfNCplezlTaf8BSUYLIo8UdKybPMazuhRVUXYgRgKhZt/M71ecerv+SM4FxU/j+DwRnL
0QwJGRaTd0j+FyAIdyZfbsWCLhKnFr7HRYgGHmNe2MAjWGnkP8vx5o+2hEe3jYCYwJeffoUQV7nT
Yf0Qzk8losdfj5X1Hp65sZYyZ/nWU8ct5V2Jfq+lNVOW1kN8cJ6QMIDZD0ljyfloIKK0btZa7ovt
aLna55s8nAA7hbJNOVNGQds1eL9cxoxtaqhW6h+TJSl0HEtqMHqYMIXQBble1oYMA5X0sTKakm+e
Qqo5XoGVah+M5hHrtRTQdUviy1iPIjr+vBTwY8SwZ/Q0P60G2aD/3E2JQsY/FIwuz1K5WNPrXiII
4T9UIkO+3lmXFXFNx9cPwLEL57WQKVK4VLkxg7DSHm3HOXBvIUY8IwKeXzg4V2upKKt8fkkT/WOy
LEAQvXfEBy8x+vRX52aLO0E92YEsvudAOkVwukIwpHChSWMbuDHWhrGaZaCIQybEw+/0MLGnBQSS
DNkOQ/sdYElpCDVle/os6iPvKnGcjSXZh7FnSaUYlPpvpw1dkxo/JGXboBbl9EQIDvUtR4iS8gvS
m/yXhRtZ4mnnMFP6eDzpjiG51VlkgiFSzuSbtsQEwrH/BZaUOeCmV+6orE9bf0805I1QUu8f1Pl9
q5FOpFH31NAVTkhwmrpNTNjD8DSAsI5LnPqW6JspyCdIETklgxe3s7M4itNeF7MGp37hRvJ8CZMj
QwpLo/L40wii+IAIp5ueuO3TKtAuXB9fx6Yy/MIRrNbcsk8kXhV16EaHeIPILcIgvTHdiyGFRUdy
LsY72/4n0SIS8b+XiFXPF7neipVF/vwqYvcP7EZ9BV31UTMOCv5Yo4O09AQlwEz6x6vgNNi9wDE8
dujeV6iKnTB2T4PEzyamsNXA71L5YJZ7zqn5SS+qX+r1acih1kCqqpRy75XYJnzVRVzn6Sk1RjYH
oE0jeyuwCsNgMi8QSpEL1UCD+sbhJmcynBWgTy84yI4pQKc2X0RgPMUVs3uP/mjlzExxitaBxHo1
lhzK4VtghZbZgoITWG5+ZHRP8YPeUJdHEohRuWY4JM156oAHyAPYOxZARmLgA3kHYmww60/sh1fs
YgXQK1n1323XsdCTopBm88Nc/lvkPkk4uKEnkyaKjlNHw5zw7cGhTNkRGj3Qq2ty5fq2TT+FcgGg
XTfralyf3urpxTCnPqdTLs2AE7KEvNJ8ArnZJdD5616uoOjLeGNEMTeGLOtwtxDaUopR4/n+LKws
/7SVTnebs5PorEv968vJVZDd9rYpECaggmXlNYpF1F2Bi8bnUR9EU0ZkicWgeyPxf5SPdGg3lkSw
jBELE1VLOq0daEnAdTJ2CRhpuU8OZ8OWEQoGzTQiPfBVX+n2VmFjsbkpj1TU5qjouGEV1P5dZDoX
q5ZMczTUuQdSP+VCu9/3TssHmY10KoIMzuiTLD/dGwBAxiEGM22UUOfV1UmshauxP0DPqdxyDQtV
8cIEIK7iactdyl7iVLBvmKYLUSvpHSwnh75RxA395dMT9DLgDeLak7obA9q4e4MoNSONmSm5BF49
vJumkm6VQs6uawW3kN2q7AMT+UVoPG6FCO1twPLUGTPz1LU9pnSiK5SvAZBkeAN/cpdotsBDghhW
ulNBlIw+B3K0FfkdT+QA/+XXxxn/bmv2e4YNHMdd10rItkAm/0V/5WHRXYzEREy5ZFFNvpq9UnZg
ohBX9lMW4YGKoPPuWmkeCOLW5XyAq2+yd3/uIdY+uafZAtmfXmSOfc5yH3AQInt1HAsiCYbH+s67
7Hb2Lkjagyp8XrEGwUu/3YvSfwI9lj3L4iDB8PqT0+AvDGW6ZRROt1FUjhp7alDpzNbN8+vu/rd+
Ll9ly/jsy4IqYS6l7bAD5Mm53qfekzXPaUVV7i2eHWijrqh/4lWpUFKTY3K6Rk8AmAAD7xJ8Uv5N
gVrd/XxIoVhmYOxm2l9lLOoDzjrsccqOgHhsmsYmFyg6180fAPI5n9j6YFDNiBVZM5z5wOLv/SFt
ue/PNM9RN9jai7gxSCn6HHNmxH+2FaYTSun1W5ByWxq/kBQE48KEpV8M0i6dgH/yHFGpI0AtU4Ww
0tftMKYBbI7Awivgdm3VIAxwuATxf7TgpSx/2tA67Jq1vgNgF9gu7pE7QEA4qJz7jZ1SAosMhXXV
1PKtiYBgBNsv4yCQIwwOGEQqOuoO3Ygc7FlqTkCvKHasz7fS+8nmlDNeibRBMKU+GGsBVWY9J7ux
fX6DEOAGldJnE+utqcxnltK4Ovd/2jTj85XuEsPy5Zm9bMNQJn0JASc9LseXTS5hpVgHgq87loEm
iJwVG/xsQjnkq9mYZ+wbeE+XQ4+odpRC1aQvBrRtwmt7yOB/GIQ7goGQA6yegRKoRAqTUBZH8Oi6
esXjqlNCrV405Hi0IuIBABUBkpLrkH1IOR47Rn0vfLQ0oJxga0/ZSyl91Et91CkFimeh5YOOV6Jj
2oMwigA9QLmWlRaeZG/iMwh0SSOnLC7flrMGrJ/pXiRB0PCVSIDV3qswCuBr20IIzxQynoYCKzDZ
GXxAqgyeF8tBYfj++8cIJAAC/Htq1xDZGLQj2k7vVAjk/0EySe+oLe2RKV0YtpW7H3QiNXZxpQ7/
Lf3J6vRjpzzDeJAfz/B+nBN5YjM9JMgy++zZL2mG8LN6yYIKps48N3lKIAwGY7emY18g/k+nYOGD
vrERJJaw/aUI6EO3NLoYsyaE1WXpTjumRPsOtHXWUu+5rW/MmVp/5FAyiYHJ4CsOzDrJ151iZE5h
uqmdQtKD5QOU1ITyxtEsdMyqlUG3vOddS3L3uVer/pxAIX1oP5RbCyiGzRjw/w0WcxLxYUktjHGt
EgVYjH6SHp1cLt8ZnDXZDQ6eiSQl0wt07TNv+Y7r1Wl43X/zp7UHy05Caw1umXAiawIS/YPPefy3
AzlHNiuBQXjYlQlT+JT6dyUZvsrIXbIWaoV9kT0IRLvonDVcfEwxiIqNR+pnGIQghlTnelURfKO0
mmT9qgNCyFVX0qm1ro1tsG0rZrAFcTJSdSvASQJwr2rBc9DcvQkKx3WCGd2zU7MXYRvJoGpWgUOI
4vf33l//XBxUdk21tKZhALrSARyi1RrX+hMj0zPTU0rANkM/aFAQaIoshW6L8Nab1Lz8KJAOAUKf
Y5OwN7eRsr7crAgUJ6sX5iagIWWQh/9Vwn6/TGHOZeRfIs/339o4T0wPLGkMZKuM5rSrYebMHD+H
UA9C5zyn4T7wCGCsMdl6q48yDbuTGFo/s8KvYdwNZh+gqhriTJJ+72ybBysSv6Z8TCPXf6XqSsSI
aZB36Z4ERvxmCwsW8rlm2AoH+3a2Vh3C17u9FRNM6aM3nb+TKPo0hNImsqy1shC9OIEM9P1i2PO/
wOa5U3OmObwRmvU5GP27C2KYeZej80xSHzkI9nRXHO8oI5vm1NpLzDCe5yvuB2Rs93tf9ZzrRP6W
l6JQjrTKESRi1ObktYu6IVM1qNEtAilKqBJ5Vb7rkzY5njFTpXSZzF3T8/ydsosib8dy3QRUKup6
7bFk6EhKD+6rFtBGqlwgicRA5ZIqv2iKtPd1cry3/paNrPnpt3XSFUO1l5SowtpzQ0qEpYA34BdJ
xEH9WrERl1LgV59zh/otgfniT2UU3ws+lcluGLC9lIeoifJwT1j744F3WoZT+ItrzGNtJx7UGE6c
C+i9vYWmu8xwQwOVMAVBj1mf0jWpLWb2tPxGD6rD8zElVAMxMw9Sa5Xhzi790jrw13E00WIUefY3
+TSO0K48Qnmo+f6IXnQNy5ZHKv1Avu7+/OhrVIz4ifs7iCkLoFVEiTzAmrECXO27NYgxVhUKHS7z
GMc4++g3sn5b1Eq4kpYMSjXCzVZqkfPi3Vs6C/vJJYI4oFmxCu0xfI9VDaJed6rTnI26o7baxazl
6A2hEonzFrY2WNus39EsBbg80MyeXcAVs02YKwzBGsIY8teVocXBPoGE6pK9JGoCPbAR7hVU3cek
oRo8ZZYC3fMCwpci/KFXf+tzIgH41ZJaUkQ12Es+7s3IjSnZ13zJxh0X9zvUe3Y3fOibx1xtnVkb
EZFUupJYBujjoQK+zOAxQrwTM1TDnXRN6SY5/7ZIUqAwFwm1lZ+qiXJwOmgVlW0eqn1edjYsQtDE
W04F7R/m3hRjB2NqAJ1PH02W/IqC7vtuAoKn3SGTM55LgDJ5hhlUF2I95lUE0fNDVxDC7/qBJrwV
pXtQP/P3QEaIDLub7+9yaSVrj3EZ+z/ZoLXPqqZQezNV+5xOuUKp3dK7ig6Tzh2d6ALgi4d44Znr
Lge15b9mbL5Tea3b1tw74s5MYNj2qm67HKcsBe/e6JDpB16Sa5PUkApMzL7ZmVUdrTJh/B3Eb60X
YQ8TL2N/OV1YqkYU6aYT4sIbG7suOqj0EDFW/f4Erjs2EHGRC+hmCPRwPba2ZigaBeQgqHUWihhw
oXZUwWtxwTnJeOyJAKbukbb9muj3vOugU5+mECIAeZekHER1ikgL/x451/vlfLx6YYVe+Ewd8xaT
Jg/4IvS9OjLOtsQvOytIqI/AuYqdAao+t9DGyKSdzpiK6pxgzvHqH+xoC3P45WUPrMu/Q1sNUH85
dD/Ox3k+TK94fMWCTU/THj6FEEQRlznDTl94qo9FK8OLNjVq/XmMKjeBpNAlKM+K8UODccEB55hC
m8R8aihYtSzYBP6cLofC62qg7o6j5e+WIKFFeGwzyP2PBPE5t5piwWbBbjgCgNnbItGmxQVvgFjH
MUgeOFR3v25gmzmH33AAYzeG2aPlmHQrpNQmN/gMoAFZWFn2xO0yU2HbD6AbPexs3SBI0pjgUh3N
G4J2E7v1fcafQlVYO6o1XhGqfQkI2DG0v916nkuTGFPsl+v97nEdlbLCGi5UIq0c1ShxX1Lf8GMb
rHX0xZdakZ7O2/wDF62sg+WwtezMe5SAtjCsNIgYlLaXMgfkiw+7f8S1mmwFW2/5M97gWgTGxJoB
CMDgqmnwXkMRGc/wvhBu7EUhp2/iNVO43nbfa44KMr2VKW9pHc744pAT4Fr1rvp52PKzvB2CG0dx
RTrb3QeBhXv+mIw0FGqy1GrpZt5K6xhpljd4zz6M+Tw4rOEJ3NBrWgEFm80ue7wKvz1kNYm2xh4i
bPGV0j+serUvbhH50PVJOvGOA2jwkvPIPN2BFku58gaEdQuSfPaKZPGbj6X83G00hIeXevj+VMse
81opjGGJS2vTaWk6StnW/ZMe0FPBVABAH2XrWX+wo0fnFmJQiNVo23uKjK/ejSKNYZ/gYHbFv+fR
fE5tk3Lp7b+M2Uh7v1mvGYzV1kiW6lBwdJkHyrKp5GYRUpcli3W1rvgeRPCuUWJ2L19GNZgBH4oX
Ilh7W/19z97Sq9a5lpI1pPB0SfQCp/CmLZWqsOcKGR3PBD+XHenB0Ttt4zeDhCRmE9q+X+BrK+dN
Eliwz3UfALEf60hmYcD22A7Oam5CanHXROc/9KBXH1KfVBJTFtJLk2m0rVW/hFxSXLXCAtYO6Nzv
+fnAl8nvl+r3Cmp72qfqaP1bNh5LclKJ4FiLrD8u3Yl91YanYPUpFHlHxo1sE/Ic/Bz5zHcxdH6r
oTeLxpyS1kyl/cSeYpxbNBeTyZOwgy4IET5fkOPghkTyHNyZ64w/EWduCsZFUBW0tR+t/8p8+xbA
myueUIBJRUotVk2elq7uaCZpQaqN/y5Huo1Tfscp/2g/ypm86kRu0Yz6UoVAI0PhpA28eaJ6Y3kN
20QgfguIl2Pgp1+5hEVLNzmaMSdiA22vfXnp8sByQ5rF0Jo8UlFceNvHjXYd1WqZEOnyOEyz4yk6
VwnwFl5unrpJoWTksTCIVLU+AELN6vt8XRIL2ayTLty359sOdlagQCmKF+wSbQJ4SkvXynIuBR+0
0q+xGHgRBDwhtFEFqdKlaQ7QYA8PhVeZIhlmCR3WPkImTtGUpwUcgI2dMHyNpagA2BblryhIOHHR
aqMklGPAivlpwTxMEG7QhtyP1Jt7y5XmCFcb7IetEISbzZFpvNsoWYsc5Bgbf9BjHezxgYSy4Z0+
2dw/JbUVq+I79tF13UAd79SAvnWQ+xVB51wODZAsi6WwuBdPo9donbPsElNK6QRDuyunUNcDW2g2
UIXs/w69a8CR66edHY70sta01tccyuqFrQG0Lhfl2AAtvMJRDniHuS0Zx3H6KwrnABHKOINptUC/
Inad2DSTZ5duPt5YvzoYgMToj2FsT//36YuOscpDnrqpykkqR+bCpFG3sEAFUiEsGa7twZGEvm7r
xexl/diFmbkSYE3iWs5+a+jDtp6iyVsoT7F2Gom+Ik1VuPC6evOr5dS5d81fXSkHHiAu1JvwQ+Fo
R1z5tL8ovddOUgpzzQVJUBVQWzfAe1VMfHsRGyCbB3dzTG7f+c3U73uLFg1L+dJPlomhWoyijIcd
RxJ7O/uk0x+xHTx/+IQueucXhewh7243Woa5bFfbCwbXRywguHa2Bd5cofwYm1QPqc/VUmIwboaF
FqE3dYf3NitEqfgeGzPcMfUO5ZAKT8MaKYaNdEMLGY+xJmYyZJBj4viP+DToqctp+RH3meVeaP5i
mxIRSESKlCObslK9ZJsnz9fMl6QpGB+GQhtcjfBGs74eXs+uDI8tid7p9quDOb+PYHC2KmY33An/
qfF3VPAKKWu+OeFzZ0n8m45H7NgmHJCSbEJl5nnhV+eQ13XVDJNpV0aTpBfe4JT1D3ZA7pcmb2OO
I+uqpB5dsJCPDkFVjLLmfdBijGhfHVc3AoeDHmne9vIs9CeiBJVBpeVJpG1+crp6RQuesLwpaktI
2gdZ5J0Rt1FW6cxdNXVP240D5Gn6JzGVtRq9VO7owZRgY6iE4jWb5km1Tx6+MzTxf1C0GIH5SrwY
wf/oj12k0eUHTP0FUKOMx2gckc144msxrlYzyum+oXgwXQOlf7AwmRwYwhgRzZvaY1Wq/GxH7cns
jEo08J/PX4uBBhfEOTwQoVPGfUIhXHR7BsmTGJeZqF978E2el5/3sK+ZwGP49B4VjKp0XMJcAz1x
b1Ef0lFDFMi1O9EUpsawU95uocsylp/KcwKAHj0R87JRE8dhnEmn3YB/FFakasC152GzIOjjmZgz
UaOamx2y8crC36fd5J1+yMwP5sF++p8GvMPnMdZpgSR48bl5wRnpyhflQxROOd5Jpbuqe1gm8+Ke
A3rBNcM7O8b1YPJ7o1rwuRG1RCXjKy/8NH/YQYh5yyF04LxjES5pGf+zJQGgcW7YxSZG3ZT6RWZi
jL/Dw5v+xQlQc+2Q4D9tD++Q6DtbQgb2Bv9YvUG6tznIPRIFAaPeZoItr69a9uLwKjv3J8ai6TJI
OyQNDDrjDv2OLFvquw78RmZ50P/qKlW/YiYobNXZFQ6ScBwXPvzJwZ9yc9UDvJroyqTzw+RmDYdR
Wc0GYbN5WIuQyRc6L+CE4qoNX/AkTNBWyH3dZ6+bKI94SV4hJIr6jf2XE9rDmd6pvlFC6IQ92pQG
CVpihG4HfETp4qxiGak63efFznOJbILjf08A8xt0wMoIk/HogaO/yn2+xyMzGV6so3B31EFgDL2p
KfW7NB2UDKuTYlkAlRxQ58tz0hC3dGj1qo4PGjPX+FhFCJ4HGVsBOMvTNDQc6mQmg94XwY6ow/Sk
xOmg+RWhZXPHpMgCfwh5IuDYSQyveIOsvGBrsksuSrC9xSW4voqI3OUOoM4GHUGaNZ9n90+o0vC9
GIZSUw8QGEwcwCVoJGIWkYx2nMdDYX9YhWhbIgbCQoDyTDg+yCXpYxX71OFIvYvv2NCpS+5sFi5p
Wape3qSKnK1lRLRjz6FMbSVb+uPZlCiFJHX/T7FErCIRhrL1x0Yniui9XRQPix3dbkdWf66cpNtu
3jkC6PmL2AHWba/OMHW5l8DJKo++IChbsj0MpcyKntUhIMgytVank4BV4r6SVzt4bdSEooizygIY
YG7+LfW90429dYl4+tigABpnap04QZH3UdPnH8OUZqiCZjv5xGeY3UROmbikVKTdJu8db+U37A9I
jDt0nZN4wpFNO9kTKtneq5LFgiQfq0doliXoIaGUaLd387Nq8ThAxOSf1GGyREXPuIZr8YgPuD7d
IY/MRXmQGvHrOToCv9Cml05XcHiTR1wEBGGellGVWWrvVPs1p5dQqWZkl7QMUZt9uIG14aunmMdP
yrd9C6kIOyAiEtiF9zQMAjqV5l5FonDUPRHLrVZrd5VQ/rCp6o9AFf8G13IkbU/C0aYA3yn3Dx8/
vqXviuPpymyNxDmGPZqEjkCGDUwdXCnoGvi12yD+VXl2CB9+QToCHw3Dryw0nSBMFnAUT5hIztJw
ecXQiPklSYj0rzMRNBnvnkfIM1bAaJxEzRHrYBaxkZLzY67eR863wFpmFRiaJ+Kjtd0E9pkZ1vmE
ymV3NkVIpdEMQ5r8zD0TG9WLKxeO+MjBtN6yK4UHhv6Vr/yZm42/HBNihHX3CnKmoN5q3exaYROW
iytK/vTisvknaRORKHndYNSEiq4OwzxujjKUM1lrz2wCgbeCZf7IFt3bZaBD75vQ/cvv0gmgwLkp
06LDBKlrfviqlYPxjUtOqt+csJ25M5VsWqIfFiD+6vSX4TbJlhpwqzNsCeUkhyKS/KggeMDhzbsK
3fdiivY+wJld7S6y/euBO2Yr/OLkAZTbLbQ6B4jzXhguhLBKCcbL7fSGoVKY2Qv3X5UosIcGKRec
x2FTXyOdh1SCL+WCxWStahWu19eTkKPDtd034mygysDA1O7+mh9qBX9kMJ09ZGS5xrmAyZ/yZbPs
IHQgmIVDMmj3flXHvatAcPM6c8EUzFO+bY265nioBJjiq0TxkliEW8n4Jzh9DyHxa1smitPbptHD
FpKxwVWSrD8pKLhaPMKf5VQOs6HMeuoxmm38s3woBxgETb7q3EfkhgfDcui1wtkBHNAEBrHXK5rV
c/Hu8li3EiT1GIuN9A3OA+4CCpRaJvO1uu2VhRZu0a3i4yyzhxSuh8Nmhig3rd4FZT/CYRlp7X9F
mFNUYGb3OW7ObUrpG8BQRHLSTKR0FKfwpSy/o9Q+OIOaLeABYrWoDHEG09RDeW/cW5xVTWOsILmi
0CP70X6tGpe3GMm9X12PxI0zgVLE7zONOcqLnehTwWU7E1a9i7aag8E/Df08wAmGF38+/bN8ygaZ
pbQX91Mz32RU+j2Z4fsi7Oom7osoZxL5a2sgbFTWczwx4fGUZ6xDDTmlxEzKBg2/+DVBX6qN2GrE
IEyZ7HXsLKPKEih53X1tB/YcoGQMWyW0HIxX0UGT1dlmCtM35ZdQXAN/PhZM9TkDw6rD3H+uZ7ll
6LgvX1NgZvwyVAtrzL1VM//a8hIoIiX+lDaUb/NZuPdF8Ju2GBJ+wFu6x3fV8bVT0+syjhVB9Gpj
7dzpFRjRv5FWbQ1/0MibJ4OrBMWkNmeWeJuF1HotCFR68lJNdMl5rw/HayRv+jopAw7L8odJlaGZ
XE+FX4k36EGxx+/S2urhCPf7HpNpRmH3wRUYYCp8L8kNBnfCMFJshy27IczeDp32ISXTOOcetkhc
9oEexa5h+z4Z+uCCePIhlwddIOMrLitlUu+PZlx0g5mFv17NWKt5WW+Zz7QtIRRouguJSgfxxN54
chb/ED9SYUfAk0ksRENMpBxPtMEyq5TF3trF3YQNtrm2zdZc+OrCDpee5L617Vvn6qS93khtJ8q5
yosof3v9Br4RvavX+Tc9Lrda+7/MLF5cnV5HJwUyp9E4eH+yn4fEpyYa6h7jUN811I5wGkP83yOs
gV7sfpfmO0fjBNhaWAaYb9YcxYmGfea//qSyTPdJwlq5TVj6e8Y0TNHVNfqSgeDAAgQlKdsBhv3x
/RrQR7Ki6VXvMmFWPfzDJUwyG6dLCoHPRxWzfH3WOb4BeGw0onJzjxN24olfiIzQrtIUojnx4T4t
rkKAd504SlR8aHiuY1lTGyZqSuHUSV8grzN13ruP3eclRlARIGj4QZMT2dNkACs0mKBDrPeA4svm
abhPbFXZ4+pram2Kml8Rf6ESH5prl/RrPaT4HVZbm442JsrtVOqIOZOHGh7xOy4uPghMMO8YLtUx
GylnEaOTpXb7M+72iuyaFXB5VrD+dvc0PEH0GG6A5fQvKzUSQ2vrgWm1Yci8VvGs3VnCnY0Srloc
JolPla/6pA5IAlt/IIOysJ8hnDdTeQbWjBkVDEbdwKdoChKu08PNEFHXLwWh30yaLv75DOdGGqZo
5QqApqfJI6IsMFAa75nAfaCH7k4nSt4mlxyCtalMC4+XpWtA7+ZBb26KBP5vA58920ouAfXrJGBR
59GC8Y77e9ooOWRZS0miJ3tQj7B11QVruqUN6aez+ftf4gQUNFzBCB8dKIOx274Mi7bea6+8SGpO
7QrLLSSjK8hFanzq4xZsOkoBvxO71ZvcozlS3BpK95CN/7x+GU9LYDQ2Me6J2casoo6UKutFl/gC
4KTj9wgs8HBv+jzH1KYeN6XNLINEZ/ZF79yTb3JLMSIJq4sbp7IXToizSGxsE40Tgp+2tk3zaQXn
F6um9XPicQKUpvAeMZy7TZTX6U1s4nTujLLqR7GWBHJTWA1iGb939G5u+t3XROIPRDiqgo5KqabU
TuB34JY7rQH/TzsXz/C3Yf/JZpO4xuqr5yal97sUhNL2p/L/E0k1yiVCxslc4Xog+8FcZNw/Wgwt
1QHfhP9CyQxZ+fKBqAavJgvshdSETjHMP3/SRde48aB+Cpbqyjx3vtyV3xnBLeirhBCQXrLmaz9r
K/22RXb6iUf8KZxJLVpB7aleY/9Cgw1ei9IdE2x9Y1/H6/T/VtGgdYXYmyt86ApG8SPbYYtEOnbB
BnqPQjiZYoUa7TVSildI9KHU1XgJr0QIrrn4hY/AzfvhH9bQLr6oTPPDYPRgtBBX6KwB4I23vKtJ
Ok6mcnvV+A9Q1DitIXcR+qQ0yXEd8QQJmPUPpkXggCpkFMsBZFM0VmunZQGsxZzlt9XUWR3mQlQG
LdGelfGWy16dpTepcPAi2zjrEE258jlyvj0k2YK15d8Eix6UJpirzupTjy1n7sF+UaY9jF4MUT66
2lLRM0vmk2wLk7SW7I/NrWLu8pWZUFxx6+FSz5HS2rJ+gfquS5rUihpcJhTjBG4m1YcRaVRyWokK
npfd+zpH/qk48k3OOZwApQQ24Q7e+BOu8qh5VSBs7gbnYa40QEA3tPQNaOyR5Gg5cGhGdONT5B+c
TKhfDdKORZ3SmcqZ3EcRGqaIx6WsKbdcz10i7ADwcGWeud+XfS1iUIzSjN0pa90rgXJVKGGekaMj
JWnyp0oRd44xm7B53LdEttNhY50r9uucNThZRUE8qU0WuWs3Iq4zwnHsvHMJ/UYowLXsxjb8n4dI
3zdd2X5r3564Cm238aUWeGZN2QTCuBvC2J2KNRH4rlxPUT/qYsPUdEHSlgd6pTXZRiRjaGWAGhDu
SrMeAgEnR3arUxMhHa72ny2EkfgBYGgJI5UUM+OhWO83ts9RQZIiSqDaJD1rUbkQ8i2yKUC2VFLN
qv7SDxQvy8ZP+DcjyfP+KYItBlIBK380ms0XKpKETRmjCfymH1YWgHmH380aXWXYJcRopY+w6t/O
I5d785ngu4VwVB0fmM6JNWw5gd2Me8j1Y+PZYsw8T6crtNywiXyC+0rv8bgnKI/D4XahD2/6hKPi
EN82lf9yKhWHEa4B5VMPaI9Nk5yrvNnIV+gn6O6MPN4jza/es5g3T1LUmVJH2o3JQc0ujXLk7zTD
NI7yqWu2IDSDIUJpFGCkgqAwSP28uwF83wWttBFws5HbACBX1nbrPwul6IvB8xpR0QbBGjw8dl2C
bd0DTK5gpE1R6lKxpeTp6Rz3Vbyk9ZHpKNYc04h7IIaSIUItek2/A2zNgDKZ9YX/emGZbEAEeG2U
zv6we24Uy0JKO0p+C0sgJrHQoY1T778jkLO3ctClm7Xkm4OU1M/gMSrPmuwpO4SRAVjTt3/XY4ho
SWI6bTtITFV6vyNMln+3sVhq3Avdz3HoalErz+NKoqlkHgVBvGA9JncVmHDx5kFN/r2Uu6ZkLPNv
dDaSIixjOglBBAhzts583KwkHG+BynF3dFHytXYOyQUDJXA9bIZuRUZJdvllt0WvJmye2yA5fN+8
wcg54qhu2m5IAbdxksBiac2DgGtwaY2/G2ym0a1hEZoRT/T/yczelm24g8PQwmeMBRrusoQGpvoW
ecTolCOYi21QhC9IU0QzuVdcP/otsAIVKEM+X8UHcUiXeeGdJ1fL8iD478kFEKH2AglVOwqu7BEh
VY/xHRHJfhiEzzGj7S2Hjv9wK4Xudb3XGwMNBaEyjtmAb1dYG5fnjgk7JWoo4jKzAjbXzvOoi5zO
1WV4DFOw2cH4glyzwxhyQFKYm4J08BlwXspRohcvTMBA+Ig8WYQgQ4i2QSEDW1jatNlIThJRjt12
Ys3iGQMZsn+vP+gFXadxWa/3YeSwaJyMVqC6WGuJr40sqsYXLJsVmUk8i8Bt8oIgcHyJqb/Uqbsd
zdAWKFN/Gjb5J+my+nYMeb1StgUeFjtvfS2xBC7qTXPn42DjO/J1irnTkH2Ru+YDSDEAT48qXEUM
7Wpo5R2ggsZqT7Uw8utpwpiS4FHfcIww/JIJFzW82lguOOtMKUbUijeV1B6V0YLw0VNk9NO1AKVF
BKOsMqPidGA9pmEy3ocUdS/fzawxdsZ7Bc/YSSn3cIUjN71kKySgbTW6mPK0PzC+CSTGUm3f3i9P
Nal6HiQMPioVuglohPO8qncrIsya3jYuR5ETPKYWjg9sENScRZ8Bd0iVoXhjEubLblOM/fQiOx4x
guXP8xz5pHHEtUzevDzwgNB9bHfB9MEGqRN6uRnfd7c7cx+MIrRjPSl/tp2DhOUYQCrIcPCYw5zZ
COMguH7DsxjJFNDrk70C63kezzhiGwKzh5TCWp66KJZkLV6EU+HTUiDvC9Vbc2vZq8NO+M0q8ugU
1q2Hx+jiNTrcK9roDRnjZWJIO4PEDAMi1Zj07+i+nUI2PDx2tJWIORjHk7QBTg/oh9ug1vrNiNBh
3chRwqkFUvcu30rwHr9u24WKcDPgJxALqReDKtzSmWgAaf9D9825Qikd6U9Ffox1daIUV9BpIQle
kJvT6V0AIE4rYUGGuURhvk+btzzCDrhOFcHWm+LKZAYIt9UmjwVGZdeMoKmqoG2bjPTMWxr9a613
PGIbkBEvwEe7idWz7w9Nk6O2MKYyigDMwB8dXonyQhRS+Y3QTcnWxvJS5fsFk2A/7nU0dQS+C/Oc
7my30g0htJG6ireP/0enQiVP5XP0W8e0pZFpyLbq7V9Ulr8a/iyeKBeYRFEEFhPT7b4oRYh0EG2E
gUPPS/SbAjxmg4BVSPYvlHQqWlU4AROoWMRbMWH9gO0BNhUBZQ3fIEomJXR7zfifX4BfVbY1HUO9
kW3EAcA7XumI+RjLojg0fqqdE7XLjoHpDw7py/bHXsEijoD8RQTX03XL3gBBKuBPpZh5VU9dUv+Q
wbcg7bMAK8JKUwjSBv0HLDDt/X3O1mssLHoXzhyoDJManwbyI1R6oXEwYfHT9tIDLUyR8OwPn9bW
HUuWF4Oej8wGR2O6PaDVBuvRAlBI9uTzh5jlgKslXrI2GxNEXqoev54Q2uJ3i8qRAW5F9w9+Q3Su
nm0b5tuqH/3cc5RCWJhq7ut9JN0OEabRUso8NR8PLEcLlWOfr+KwYZEZt0RDg0VBTFzbsUJvkFR0
/PNw4sUC1XIolpBSTgfRjtyeSaBEofTlEwIAhVbkSEP4F2RZNJNitgZCc1fJ2CtFt4Ot95ptdgUo
Ddgg9PjU5dVZIZJLjRvs2s91JtaruyRfCKRQ01Mz22eXRQMErFDaloLc/+fe9L8xfRNLCbUjSKmb
ycdTacTcdQnFxVwomuNitEp+PAAek2hBon2Ve8SpOKaa+OxDRAdPTukpKMjWJc00rsEj3tWFsW4x
jPsXAWaXqkRvEK75kgTS7qvBQ83PpEN+/mV+K4lqf609u4Q6UBzbdkfp2+PzR3aFVqwcIWTfLev9
R6/SlsFLnL93Lv2jU25mZ1ORgXWeXxgomdGDnUX2zkM7BwoY2Tvi0rCnTPwr7yhm0AbMjS9k7sSA
q/puajJiq9qUR3/C/79HFn4xkRx54/QZSSyWYRd2f4av4eK1zrjcmYqJic4Yka9BvlXVrlc6qFzC
0r6z6FCFfli8AWAidJBt0DXnql87w/f/g6oj07E6AlHBnFGon94gNkYebvYCVhRjP1nTijYmeHwo
vHbg4cE4otmySAm7rbOkzcn6HiMUqybh/uJ9y12NUKIRM4Vb0gVF8W9aMy29B3DPvfhgM2mJf3dJ
TUpuPASqJrLvRCQO00mQAawuI/xY9rCfeQZxFcGlrLha+kYpfXuIxRdfwlLJuSD7VeYHOA3KOyea
zW7dO0459DcRDE2/LaBCCWHTyeGh5eOq1IrdJ5yi9W71+sNUMU4TQCzC5dmCwM4PR82bFmpaUwVv
FFVmRVfIhgOCAWgmIxBlIN254gcArXDBnduHvvckfnAnp9zE/k5wUSqOb1gJisGtQdi6arCnsaC9
SjnyT/F3um2mxx5IoHm5MHX+pjgRvFytsAgGEsnlM6QEDXrUDqsDDoqkCgm2K+QPXDq483rdQSmx
mA3o03//2vM9epvm9NTUGIHLAjFnofCl5gbDqx7Eli0Qe4h5kQf3smTteTVeOk3SNU9aozVvN8Z+
R3QLNHDmJh6njU6n17CD0wJfke+tYYhH1qRIlhk85QKqimrLVYYUInnCCHOR2bnZ86NJ665bgVUu
yeNLkawtUgXfO86GvmC4mqVBKJk5/J1Qz3QGfdO5707L9q7iAVMuH/dVkecdFsqjHfWgD6HyrKUC
M32G6Df9aj1U9ikS4PkkRORdDqtKawUwqbcoGOdFvA5BwFbONyplInvN/JfDGZ99hC1lXWsfdan2
j12EqAOUScBLcbSv9aVz5qaTPPLl6TkkUTz3QtbR8x48zXQsP//kjkTOuYtJEQcBX4P1fe2SZ5LS
1kZ6kDo1kOy5e249d/QXbE1m6/Qj/enzlDqdn8ZMOA/CBrgx81NS/ewU4OFZwBcCfs1g0ZcaY+Hh
/7naGDtU+6qI0d9hrp6U21nCWhKML0mNOUAjfckjmaCEuXeDeapqbaYcn1Cmi8KQ5QNQXeQZERod
X/WU6HUKgRk2aMKP7aUiK+VNiNJ6z1IfazbsmI7qKISygEuFNsgKS6iXTpz1YvM3N8s1I5uo9VJI
uL473prgyV58Hv04oR/LqJIBmQhTn9eOZCY8QCEVIxWBU/VuYnnQqDvyp3GxWKijhoxsngu2gEbk
+AjRAAm2RfJDkAYgNXSaerVTy6bx4c0IR6T0NFl8eCC9oi9CBeL2pjqif7T4hBLl9+ML2VDTScbb
7t1SGnAg2N/Ky7BBqPQeHD5jC+WN/6gub7jQ0UeRpA1Hdl4NkKZmXNbo+M92NGsIYVX02bn6PpSG
2Vj18uVJWaLapmkH+nVMrpwCt4+17cXYek8hbZpt7xgqRZs7SCTSYGwWDRk6BF8ncwX2HQt8Qtva
VUQoMbc//pcYk/vQnt/DTv5A2FvcSTw3koHqK/8egYP569u9qPxhoh7sLhRWFFAZ+XM+yryyZHaq
NT40svcr1srQzyQVejgJQ8NyPXhW4Znnj42UHnzoH0z2ZZXZfIQeFFy3Or4qFWM9LjeboApQJ7NO
keAeffZyFsakwcULGiGA8Nug13dDgYOwQLtrPZAEwDYY0b5cAbIeOgjQ/pQRKcDXS45rcsZTgfc+
zkPPzxaM8PBYvP20FBV/kTLSBxBZiqeaxddkehTJHTiRNmRLID8lBHfxA7uJjN5CGY9Slo+Tb1Qb
allZQd8MvqalgZolhr+7nmriHk6YjGEjhXVmX/VOyPPlzsg0aIgXLFE/ZaS/C216SivZCvY4uqfJ
lP/s8MBrGQkeruyMxZMMYClCGzzcU8E4ngxh65MBHqmkJAsWs5mPXYTgxsyCIlPPtN53M/dobzqo
u6X3qAO5s+yCkuJn+ZfQ2Zvq3BjueKUdhFrD3TjkpSLszCwvWALIFmNo1AiKPMcQOWtW5a3oAM0z
A6w+sGuBeowxKR7R+eLc4zpBdDvD01gdsDadxKSN+0KP+mGVRafk1BUJfr0Nwga02bi9nv2smX2C
sRjnGy5EEddaO8rjuYlro5h8ybK+yEo4Zd/YWs7ja1uvfEwYDVOXOiCuL643aOtISKSWRTFbBrcc
82ugCfimBwIjs7vEcNJFCqzsWWXTGfYuJAnToaH9XkakGGNSaa8191j8SERD7Did9pA6B7l3G/EV
uHj2BgKBr3yoXV8f0KTBIBQklNwwMiPiUDQkPae2qS9tl0cwfeSaTPY8JJQvJ/LmpCKhRbfo3IFR
rfED1aQYsKiLW9ouovwt1IhvW8Kddlo10i9yal6QEqRm2NU/zhNGu9r5a7f1GG2stayTLPKFk1yX
0FQlqgoUAAp5N1nDkvytBUJT1uD554Pz3pfeVJ/NS00hUMF/1ZCvxM6VJYEvO/o2+l0uDXQaELXp
m0H7luYzCS3F2giLNxF306/0v7tG1KkHSZ+6cNKfqpiB+wjx/m8bUHuMrzaU0P4MRPoDPEQ5AXpg
fMTkYGzs86n6SwIhL6GAhO141CLUoAe8d4bF1gjAvMrP/beFKVKT5O4TwZMqT8fG4y79KjjHUS59
7WXA3oNK2SEUKgatiXm0MPFeDVZVmpwCIPYsQkd0Pud6tA7lkc797CdFSeY3p7r6xRUpBYbAT3m7
Y6SwS++RFtMIVOv0IMHPV9Zm0ax5M9hzraQ4izEdYenFMOgLkXAis6APf7NHibyHvyKPix6Lgs9n
1f6QKzygJfxQTUlZtLd7fMIVdBWMeMniPlQ85s1aRXuaFWl3taCcgOqXSAdFHxeo+sKhp9nr7Hyd
RRbQt6svwnoYXKFHdDQED9W5dUcW3ut5SNmSD6vYQ8mdWM0hFS2eyfAkrX/BsWENw6rkN0o2pkOC
3LlOQAKAfoxQsWxtta0ej6O9PEpOAKdyXOmF7XpF7ARNSU+afoau5vRPINh4wYWkZrEspKIFbt8v
5v+S4ESFvtSP324A92ybR3CHW+9wQ69ZmcF2KOr5N3l21mVolwHhkBsptefkPb20f8gL7eAaA9YG
dNaK6GTBgF/XzlJlb26ss4uzgNYhpCoAyKFYXUdWKh5N/DjLj6s1am9sMfIHY7tq1CqyJRS4sQ73
WL9zO3+d3kEw/rVFx2GFqFhDssQTO57aunEr/hrvwbDwe0Uy6NCEd8gLQ9FUZMDVgjM24rachSeY
TF/ZghfANVs1HDd64iiyVlXsbecOJF0gACtVBEmafQ+tdfQhQ4QX6+QEsLKkbaq1Yyaj//ZGYhQv
9WfiG2/kTFWy46oLd9or5x2jqgovNhl+AWJ7WLmCzoDVpVrMb6E/DUIU1UwvtsrJEcFUbTHE8JcM
17TEsOJh48wAnuuHFIiMjxUARGJ6PeQ180bnQZTfjXEk0AwdfRIchNEQ5M0UUZ4D+ChjccB+xMur
fXFd0HTEDcmDHuIt3tpteCLOVdEuQ3uFg/kqQQNp5+uqgqps+XrcOSusC+33t3fyi0kt6YxpcK3U
W32IC21QKafUnEkKa7fQWBN3XwLvW2K7bktWGi6YLlaDtiENRsoAqMHXrNrXMvnp7bmqS9SLSsOQ
K6JOkyWUg3+ycw6ohEWMB3w740jSvN2uig5bmmw6tfKKOss9iOwBLXsT4Qi7jFGf9/erGRmOJBa+
WY/Ap1pdPJTVXVDrkxAg896XAAILom/CAH4JWBdE0cC697cex5sLABJnsBDzitW26rakOym7Wiy4
B7iF5LW+1pF4SRU2h/dLXqVvyeTwFcC3kSNm9jxfle948IT6Vym5cVkcFyMnTG3zYMmGGSCizn7p
s1Ii63WHCbNh8mkCfD6ElVDqdAuYElmJiHJTHluvrOnlRDBa1hiJDU4LhjzlfuMG4RJnvLQm+V1H
Weuyl2q9oU2LubmjPbsXtPheWQrjiW0ZeSzhPhHCbKE1rPSfIqoD0umecM5D1JgUJyqlXhua6/XA
HB6/xjQnlaWu2lJxvFwwu2fZO5znj/u3P1bSH5y8HWuhdNCDx0ZCh3caUpNS5/fdAn4moU67Mifr
AU+J2t+PBNZOmge8e7/GzTvNF5/XtjH7XFiRBhBwF7GEkdGKP04CAPeERRLV/MaLS4YaBteupzoC
qgxz5wPIw4d5GBd96OYXL4l4hHJGlBc2KRuePuGWGLgyYQnrM6f+C7qjo10i84xQAKmis7OZDlyx
vsIodtpwtZvAwuL2PaJRiYjAFBV4WWL/QYtgBTTOatdjqtFiNhAH/Q+FPeRyr/DBsAsae/QvoVkk
/yBkJz+sgyuvC/B+ec/0qNaPSXKY1VeQFGJMjUIIduic32xGoHGPwYVrsy/si75bKpyuXIpRxqRq
6+RgZXVbEUQE8tKocExnFwAoBX3ZlcKewI8YWZ2QmBvl+LkgbUPmFtKnAkbuDxIMqorcD4i0Jmxx
/m6nwAcqxN+Aq1WRpp4iGRJRnFlyRU6nJhRkeb8EmSMVo7qDRO3RyQ6IMrKG9zIDdSzj1y4gLGpL
36t8v4EKFnXJvNn/shrQIexRPt01pUv4p/PPFAOslunE0VvmefKHG3u+zyuyvIbrhlp7PVQt+gog
pMUxWTEY4VPAE76h1de5FfEVfXRxVBy+/Jz29xIHvA8VN9BMSLUPQqwDk614TIV/sHosz23I8DMd
PkPPbRHGgTbxEzJrUoILuJaSfX6zuMNjeBS5JIWcwhB80lV4dGlskcdU87DYrZG+4VUB+0iFfUT5
w2bNfkB1wozQ23ows0tW2IYHaa8r5cHSJlSayAHSYMuv1KjBG4iievoujqBUtovOB7p3KF6WE2g4
ZRFgGhJ/0f+M0vYTJt1E6ClfDsAp2Dah74c4jlTNe4OubS3NBogbQ1tvxEkC00OYU9Xa/DfWSNYn
rxY8mKRu01H8ugi9Sfxg7dOiKALzD3Vf8cf1LHkZqNH/LCXlLTGYOc+UEYyzxyIg4YtaWeSoFIpM
YdaXZ+LQNH7jroD5UGDUH2bkGG0KXtwWdGzz3PG44fNVUqFLj6zOPc/KqayLjyBZxgTb2IMd0DY8
XvPdYX2ee5HXyqrozGYn/eB+LfY1XEzSHnb5n9vX7C+PBe3S7GPoqNR1llEkoBSk8ioilg+Tcx8B
CwuLcHJm9B3DTnTfi71OgeaUkb3N2p0vE8dblbof++5CJUuP6s3r1beN8tNpuKKvyaHppHAQGS+2
hMfWcKDSTByrHvSie6ASKVhxnaZKnsrOUpOvSI465sr9eSVDAuZYF2gsrQGNcIt7+TFzSFEaJrnV
G5Q6JGr6q2oLdGN4i1odlSsQxq1djH/l4gew6g2XNlUARxZ6zJmJh/dQvmaBJAxMbrMhcBTH/m+i
0KKjWBH0g7EVcHQs4pgOygYcJr8jrHPmSL9ErxpwlJwNGXUs4rq8bLgiaTZuarOMpx/85HS991cd
cPIQ7DmM8yWypYWPVl05Y9Hc7nwiERdY96pAYucQwI/9TsQdM91TZ22OgHPtlqGT1zhXBFndtgeB
yAUs/GbkkCT5rIlcRGLravDi9SSSEXNiUACWeo/ZFRiDGhbLlwvfQu9sbDNdRtpCFr+rLpoqXn/+
AD4OR4FtpWR9who6EbDxVWJSxzNECUbAnywJkxQuBuamQZ1jk3D4tw6Van+tg4jG946z1pQCWoV7
CGSEjxgGXCn/DQW9tyPfmZK1BGZU6pWlt8kzIOaENtSz5DeWBxqBNyuK6gyhD8bEXuV3N0Rob/1n
Btx42mDCw+8jUR9dkQ6xdAXt8PsQUXUf/T2CtxGj/rQLvrvRPyhFH3eytucNQzlqJu12n1ouT5Cd
QXQVvXahvV4RZ/DG9/MVp5eyOgB0wDb7Udkpz1O6eeX/Hcy+8wQJxeSM1ZNJPTNObWYxh5Akk1cD
socvThUegmxfmYBDoCDqpCaPbS+bBDLr0pwcsTr9THdx9laCsP7vgrZxt8jb64JcnNAiksNvky4z
vpspbKQdrPydMcklGOc8OQiSEdFMxJuvHHPACaJSuV8oIn1r6suI3Sx6fXTNJNdx7zGKjZyNqKUS
OzAFQOKyFIXYaAPr1Nj2ZvHH2oYjn0XaNgEI34M/oyxCyGYbacLlVOnss44SakmWehk66mlsyb3x
68ifg9c3HnNci8+W//YSmq9B8iUQXCG8oKRWNObThf72JOUPHpnRGqTrdJMM9/3k+3lzjUsyOTgK
6aWmzFA7Ygo8ed5HcNFCmjCjkH7X+zms7JDLiaNeGPc7YOaxzt6zgHeT09Ft0F3stYvadDUyieIh
6+ZfJDNbX65N9ODqL9lF5FjvZg4UQxNuz7p5ivIkqlHZc1lihWbx20QZEBcxbLKg7Q/FdiSIZ0J6
/16MEruyTaZY5HFZ+v31KFmNr9oPHgS4nbZAuJ8AeIuqPIgUzOYPjal1OC9XoC6NF+JCmLrvw2t2
wFU438uZpEaPOO0L3C6sQTFUAC5otj/EQT1Yo4hA3ALodAmc7DlmdteDuxA2//9Bs964RkwHnGP6
uP1kONKIaSWp9+v/gy+IKt9lJx/B5zkN5KvYzhWYCQxG3diO0PQvuCHRThfjbVl6ezefkrxb7zcH
STx2OV4Ue2om6pgfrQXl/Xn78g4NBv6jUNHLST8piZk9co31IL6jKtGGka0luinZStDAqucKIyTx
cI0mKF7ozzNkHSDWVOn3EfG8Ru5bu/kSHMQ6ah23H7xh5KAekPaZyzDgkq+GOk74xMbtBu09xwvi
NZ3g5ty8+FRyYUKgRvxEHdbXbtXlCkFZBOlutfNn1IsbV4mDpytC0Tdb7hvWr3J/L0JaEU5o3wxN
+F3NsxVlpqZzZh1bDHvV3FdnVexyVQedX9rR5PWvICkiXMjnHHvPT9OgHiiv9I/PBRQf32w7In4x
Lq3GyU5kG/uUfUNldV8X2/XN6FY05qbefdQpZF5KKiHNarSBfISA4PSOJOhV198ghwBDsPo3ehk7
BTM66ffOQAxnI2z0D5r6N+J9P4jQFEZn6CaCXifmA4IrNyeJ2uXh0n6ctxuXchNKmCWm8QacjRUc
W/T2brE7C4Hpt50dKAzl8j8kKXEYxTG6OSUWdJ+6rNzflCXAITSA2oXIWMXqmvZjpx34Wl05+DtR
MwZByP8w+3HrHe7w3trD1AxRFunlpfcyAypEHgL1AdsX7N3NOGcMmXhZInj2uBSL9QUwL3qIWKQV
fNUSHlh4qd5Pmv1LKmCL+L07ghw5tVaXmrd6c4Hh092xpKSRF80SF6MqAEJ7ze5XwRoSGDCImBvT
ryFgzFS1nUGzqvwUtKrlwxv2fdV/cmb6hKl3hpbDKysTk38pxcFN9uw7nJ80IhnT6RsdQltehFdD
oMi8+Jr31DUbjj/GHty1EO180KsK3t5OHF5JJckVmRNBWGiK/VaHw6xB4aQNoD/vtABO/Frpu7ea
Posz9vaUZgJrmpLl7dhxut603eT6lbcYeKzndkwADYw4svTKR3V1/SWw1vcmd9GxbPj1xYyDP4hu
5Yx1rJIzr3uPM2SuAlt4VCArHN8QNV1Unq5LUJTPOj0t114jbs00XwqWowGmJB7XHcAqEr9r1ns9
dI4nPYRa9pWgBMo6UvDZ5oZN0hyF3In6b+P0cfw0hj6WAl+//CUodwBpOKf4rtS07fVuFQlQFR56
de4kOkaP49suq9Y2TckX46A9Tk1/X2iVQZVSpLe7jXf7P5XUf9Y78VtBWMhUI6Zb+fRT145UnBAF
4iFYEjo/6JTvv1GVnztIqgPXmJKLNNteEgtHnk8owg/WScczLBW0ApZ3aqM1hsZBq+9jZGgkSbwi
KuXLQoXj67jsmg98dVAHedrRrQgmh2y5ZyCPAVgEizdt7fkYclcKREpVKeFJe+HJyEefmCGu7POU
KfVt+S8fN5SIdHn38Buz2d0ClhfsYprkrywbwfHYHg+8Nhdxtz8BYQM52u1+CNckjQcRjO5PGbPh
Z/1kmN/YD5Of+6ItNHDcsKoQPdYr2Q5RPPy3ZZgv+kr6C264d7jkVoNF67bkXC52O251eVhRz1PB
zsciQmmJJlpUITtLrJhmusj8oVQUB/Km5+2/NHfV1NGV1yDODVd6xzLtb2V0QNFhO5wlBQFKEWQN
jwjGE5IVYOZLW9+STy7MRTSWWCVvYsJuz61Gniee/crUW1XXa8juJTx3ITnYZsKnKLP4KZmGgFPB
YBbLhWht562nJH5w4FXsdKl1af/Gi+7RA1LS7pfFhuQr6QZSX5PlWZTJQKVeVo3xGccDIsnS2YQi
gVxgtRqR0Oq16INxFl2+2qigvQnJlz+t3GbiPND5ORI/S5Hpx6k2exeN0xi/0/YN2uNDo5ZiGoHg
k30UPuBlMe82SP3UDWh5PlYF5a3mEtfWDXUj8WhuxdTO33GN5T+D1iQe6PzpM/HIV7mFZV2K2kfE
DI2FBi5IrXVoPRCfHBLfD65fHI4Z30aVvO7itg1QXB/UbFbInxURQFLQHcIx6KasKIwkhqrkj4j+
gxvOtMXdLNt7/J/wdp8AuD2zEDN6FKn+oGG681veDu3iTeemWn/5k6WosfVkFvhkgfKCwPESXig3
CATHN+Cjnfbi8u7qT3Vg+xa/mcGIYreg1yC3EnYQG12dbXBy32hpcnkPzenODykzP4rQ+zGavzH8
QS0IkPoUTfJH3mDVMqdfi6uJR7kmhy+tjrnu6wnmIrAS5Qh/Z03e8iEKzZAjsLmrQmWQzXJOE1Hq
vYPt4EgizINF48hcovotP1/CRGvfy95oFLBez/mn/K3qXteMQNZvE72DM0vRV0RCXM6jh4/8cZlf
gLuLRxiTTcgpLNtODhAeNRl1qfDBfAmHdVdx7vjAMs/OBwCdTrqFSJJZ5rPJl1UxhvhsrvCMYkX/
Qd89xx3bJYd5kj8y3YQwKviR+vBSME1V+x8aXNIwniB/Nic6qHdMoijNas9JfLYDWwLF/IBCWn5w
NCyua2pvtwbogZwbynwRl9J2ZJKVALLdZd3kpHqSy8UEEVsK10Cm1d63RtWiBZ11tFhRCfb4MQ1o
ZIllBzqZzrxp+85tANx+r73YGB9aq5bT7SpcFh8u4FqEEYOo5VTXG/nXYemRPsGsucp2f4jawmXB
UbmoUFUP+/HI8Uz3OdmG393kypIleaytUzRC/b0wIaGxOR1W7jbpacxR3hmAxXO/cXnrnKLxZv+p
qRFukLJdychCu+BeJrXmwVeDPpbrAhhHd7vbQOma+aV61rLbHslKRzX9dP6Zgl2xcpT9i4PCtJby
2GrSPbaX24gtcUug2XNFCUPxvosRSuJ2WXm5vf84iFsyvcHcDvmgu9iHvyvI9lOBKy9Xk89g3bVi
K3PYkFnCKuCu1APAOiNQr+B2X+3z3uuAe1pOSZ645iTZwPNRGqK5C4572xYwNpwCS++MpL8p3Eim
lTaptDTja7rGWq4NFMPDexxk2lbaR7YLcJmL4MokKcfIcnlxU/+06yg2aqlSUtKVA54tD9gQ0XFk
7GiVmM0N/XB5C+Q/ioU8AH67PogDfHD80x4dGEPp0NLK/l+W22/XDUPpqOUVNMrKUsoel9e1aUwt
xTg/WphguQP7Yj9Jo0rzv7dC3mBJCtXZzXTp1ECOrK6Ax4+QzQ8Lbx9L5pEUl3wzUvb9G4mwMlhn
AuLOqLwDIJovpm1h7X/BYyLQDcLCvDfgNCXKDzWB/2uFDN8fEwTwX2kxzFEYT8k6oplYal4FAYd3
bg0/jRwu1eeGRzDyjVB8EwLlrvKPntKX5DzWh+zGz5qEzoB0AAbtHaPfY/gNATl86p/02TL/M2a2
tqaqxCnVLtE4j0tJrS+IrswXekKdMPMJWbGm0Bh2bFXESH7mj7TVjDRmmYAEVOVDGuNpFt2SywGY
9jlq32K5IVEsVHQe1Gu67qldqTM2sQwaBAZKqjQm23DEKDylouKJPLLjU0JdDl0GLoOaTVFN1sbZ
xDUFhqzH4LZwabO0TRPEI6YCDHILyYTL14rnMrXa45QFgNQFBrntz0t3lLi8Tdp2CgQnHPcU9Psm
MvL8hxPsk31lARSo8MHNhko2HmZi159pJy5ywLdfNDmWC7EmRbm9+EjUPKJegBYD5E//Otm5fbZ1
2+eKOn3ur1AEXRgywDumQRadQ9jxB4ZDz6VsvqPaC0TUj5nsuVUUc0I/S1nr8nusVXYtWWSYHaXl
L9wmo5gQjWVKLINsD+SGXm6tx5rdRNbLvdyh173sI4X0i9NBVgZfoSmZVc2g23pmwRMhxz37l3WV
PRlYMMNFmEo7wMk8dffPKcV/vrGlyUFpWMNBYaUhXFbHELROD1MwDipySvrbRwtKtXXNx4XpCbtp
2h6RsEpI6b2HmaCQmAGu1R9Nf9YzuZkfS6bOPFd54p6I0QxlqRwvBS6+bxRVuZ4Zi+dIlDixKDiL
hz8YHHNQDlhdhS6CfWVYg/fFeYy2BP5RvKYFoaf5upAxxjvdzBoHaTXDFM/x0FKzP6Mg4uM6i8fh
KmtkqrXrdoVraz39rGChyl7sHj80izTPjdzrGJOddXwYk922AVFX6WmJrUsqOzO/wWx+nn5iZJr1
weKe4zprGRiUztpe4EP1r9wgvhIfGAMboAo9XPFpAe1n5WnGmJwbOLfydTAOx1jQgFvBJ6Vh8X8c
2XSEf5TBtsFTJK3P3uxhVKFPzJgKcVdkyVrC4S82Wg1JxhhEuGoHnmebHp7yxr3sfhSShtMZJ5jN
3TK0k5mioM4xoGL6Hd8cqP7nMi5SwME3ODYF8rAIaVVqkBOFu24XiS9TWObZIfc4TrzF0SyfC1d8
hFjtsNAL9qsu/7L4Hsud6Q+SiR6PEqJAmrr6tV6UA1dVeAkE5U++2oJBr8lsIKHc247NOM0HbAjK
NzHgAZFllBfdVn1mpdcAb10wUyTGFlbMMnpH2CgksJ83tGG26Uvog8rNSDx1DA1//RvLfVlgxOp1
Gp4y6tp32WDeyqQ90/xual6VML/u+a9u/LWvieOjpy3hZID37BtgjnobfZW5aTO/0d2I1MyLWXco
eq8pBHJeZJ7f1/XcdKM4Z4/qZX2mAn+bHUoesCBApoP0vproQjQIen1s+2LBm22FwOWm7ZmDiP32
ToR30GmJob1v3aHSO0ffk6wjR6sjSoUJmFKkK/xIZOWfIB/hDyH9veRCKRh6lCYud45jqVZXaWMZ
48kKMzLYh5s9RHyENO8doLk3IZbyGLoArI+rSOEjhAhouyJFmI3YNGf7nqlFHbI5tXVk1ELYPIky
2yNM+zzc77MDBXyeSLUv/zTRxgzzrnxWS84iyaixibDCdMs+8P1pQSU/q56k4cx9x76bi1fmK1XK
I2+d7A/Ld+LZBlUj76O3vot6L0LtRPc4pUUj4wK3im8cU/ZHHoNokcy0UtHf98UFJmp+/407QK8y
EKMbBsjCTvV5uXqAoAP4DdEDbZYicgw25BTXohvZweMR1Dsz6VkfDEAAyG+QeaAdoWMxoTX0rYK7
Mt0KkAmbXoammx0hc4Zro+bLtop/NaNMa3VXfKpG6G60+H9MINM+7gJRnz0iBK/SQ3d4Q8ed6jgw
ffV3nYtf8j2ptT38CbEr21PqFAOIAVemvC4OhHddlpqmqNZvKYSGBLh0I9VQVm6pqWLMPos8496y
ZJJJW28VSxm4Ehf7/uFrQ9wRaRay9nfBYpsCJiPib3wEa1iappt+eCWZXejUJy2VEDYC+ofr5dRe
4d6TZqCFrC7AZiRSk2ZnKyBpyXPjgEMPDT66dkqhb3ytxZxP3G8WcBPg1+TA34S3mpZDtViyyB9h
chcFNAbN0DXvvr/PUsVpmYWTGDd9pQmpZl8eZmgDcqLCJoL7dXM4v2yNynE0truDpZ8fqXhZQUuA
MHrKyrMEgTuVjSlH6m4jhz6XP+L2Zp/RwGQ6Gy/O/AhIXgWqKSpk6ayklCLboPjXm1qxlY7Zd4Vx
nh18X6nUSJGWZl5nriWXD3CmnIygGcn9v6OHjVZ3FHtTpqSLd1yDWk73kaH08/l6Z+QKnl3xAOPd
G7MGd5D52Snk5Gbs5hzVvTo0BUYKLVSNBvIxAv7zkB3y+mTkBFicHqUGeMQ/n3cPgyZzBZfzlUiR
YU8KOkqeqvGHqFtWniBwMwzEAUNBN/swcyPsFVbMDm7tOyC+bJquUAEdOe+jwDhsYqwIQq1F8KlV
8LBZ6DVEoggSXxX7whjw7lgwZsegQebrjeRTfnjbI8ic3UPRK182R9D3uziOPsT6KiziKil++PD3
K5c5TEdpTrlUsXeJuEtT6oIL357jmO4N7peTxMqTvYcU8NGo8czFmX1/z2ZmcjLCIdGkg4emZz2j
HanJk5hFUL5rn6A6OKf5u79edDavKbp2IpVU8pn6kKeX/vpOBvGSJuKAGz144sqbgP+dRIv27+FN
VvRefvP9MyQteyH/mM3x41KPZu3v3Xcmf+l4x3Wnc+njlgI3dVrkcHvRjef8c18W8bmZ2icINDCd
dtaVptFARzw9xImSvxE03Eu3oNIvCXitfuK286s76wMD4CC1Av+eUuQWc2DBBcGz1L6vNV3szWX6
dYiGbYylQ43ooYxKqAMS5VHKdI5TAt/YK8JzgxCowBrRYuMVhMzDpZ2Wkj5mxnT4jYgZblQCNP+f
p6Y/DUPYR3MBzOhDc237tRe1SqNF7qmeDM3Eo8G4t6EOsufl+4ph6/wS0pm67hjnTq9GprgHTXrI
+Zc3veblMQ8SbLoHeOMRGtpjYfLtYsmzRaiHhPBZ8aBrhM4G4pX7Ditmfnk8/ZAW3kwdZwhGNgk0
NDgx3N9UC4bAF8hONl209QbF8dWkO6znuPjhL8wtNnTMGsX6MN+KZeMlFnNNZ4uaqizKP2/QWrC2
o/Qltfvj5Vde3/XfOdG0PIKgpSMKBgNAAFp/9JLrq5ByUsBV5QdWVzez7VezzEQKH+iH9E/5j2Bl
3bbhKgAp2p7c9DdEldA6jSN9mYcgQI7Qy8gk/3Kpei0XdMoOTdq96ab6p+7keWXUstMnyp8D5dnU
oQq+Tr1jt+riMKaDGdTaN9UEEnc9Xjl1gaoDaTxEjMYMEIuqA10b2ZQGpxsk0Pg2oz+Fdk4hWRM7
Dty0SOHPeyXcXE5hnzP/5IZYWgR8/uUuEPXVItwZ8eOVbS/dHpGHvE97yGBQbCFRCOoL5cxvb6lV
AH8bU1s41zJxCd5xPHBjdB+nGYmL6rDm8xka+NVIFzEjOr6GHit/TspSr3orWNdlb6BNowVYSdqg
ym/XAyvu2Z4fXuTOdOxg7vmhz9pQGC7QCmM0SLCZOEZmapphW2Y2AvtIs2GyDhsny22DgjX/uT9e
Wb1FG3AqnAfycv0XauasQLsm/yHb1kFxPiAYU1thj6Z/x89M5aIxxR4irK5sCU059uL02Rn4jGFE
0rFINZMXBuPsnQoEtwGMSHf1ybURBeM1lZh82A2kmmrf5/Aj2xjzY2iFaaCCDaFLvwuxlEVxMN53
bpYAbCEDBcyKF81aH+EZlm44rKyUMirIJJoACW5kpA1IRRi9663Jbch0BzuPfZDdPFsLZXSMkNgS
KdqU7Ze0IIm0Pbkt2gHScr4IbfuSgilRIR7gXoTMfvgs1Utdl5qDu+6VI1bcC//0CbPY7AtkvaFu
2imXNyOwW3Jhj4qqb4Wc5TTcmOLNSHVWcWkhLyM4Vyv/zz94+8blf1vl2D9p7QQQStovVU2KjBEr
09Ofzi7o0gVKJPvuQzbhvcox1NO+dYpH9/sEp9Q+P6tTy9RTPNVpW/TtkNjk3Zov+Px/xJakoWJ6
3AupMbEfghds2DVIJk2D8KVOKLCVyhzZfsrZDxUo6vll8Yo2EnVU4u4OspF2Am8VLYRzKs+pVs4y
di4++C6/VeJHQeVRPbEX3t4dqmZX/xurcsQ3rnLGyHRQha9OaYdsM9BRsdlYaFD84c+MnBr/+sQE
c/3cL0ibcofYvo1Rvqck+VMYFGlku20aRy+RhjiVUQDkp5RZr+vq8Y2EFsJw8jiO5EWsBZYP3BTk
JMV+O4hvN3r0pu+8zE4RnsWoqNiG399Nc/Eu6BSb/Hrk6K4mbDVWNPM6OIdLOVQdTzgOqGE52uwr
V842VCEl0i0krUza3dO7PO6pQBJPsa8s9TOKpooj4TttPHGTAAM0XObBNFA8gpFYdvyVG1Dd2GND
yoz/VVzk96HzUNI3f+GPm9uugX79xslOYAYP6LA05B+IErvvSA60LRzejDbSCSeKrLmLBSTKWARD
Lkr8wsJTO3eHDjyB3EKv46jnXOe3Ux1EQdqCFjEs9y/2Si3eAq+7PwYC7b4P4XkR3NNvRS4DSrWJ
mJq38Dp+sIF3pD/sMhd6rKK2SHRpEVkN51/HYNxrYilocXrH1oYOavOsEGAsJfU40XpiI04/KvFO
6bW6hcrtxgxVO/LlfZZCbn0+6hqzOHg9rnUoHlkFMH/LIudyNQ5e/nNmlPfpK5dllveP1CJ/fDBU
UZPfLQeJVuXSosxrm9T6k3eYRxyjPwzR2BcNwVGTavOJQfPDuH64ro4qW/GD4UEjVku1/1JYJkkx
JzoAk3QiH8tdo9P5YQHQVPJx8lpXhZ9vWO5uOxHm24plLKTAOiJcbXBz6PUKSFdG+PNPdnDBo7Ab
3Gm84qghWNNLCZDynoRDBwqPryQZwG/n3KLIaIaOHf7IB3kiQYVrZwsv/t/2rmoTPqDh/LfBkM6A
oWmcJKR/XYeySdofv4jkStQcnNpyUWWyEgjG5Fm6337iP5u2HThykIo179R0m3GLH6nzol5W+XDj
5AuFRsp3RsiVAK31ZnrYVanoBGwwY3EC396E95w9KYrAq/4ny8KUMsxDjM3Kzp9RofHHpNhjckAz
VbiTmY3yfpNTLRd/PgFiBo69lhsICna3ojLeId8M4SbOKu2uXZHsf0N5b9dhrW5tPFbsJwk2+9OE
4n/teMKE5sliZlT1DaegT733l0m9qn3eljnQmIgleGfNCQYtJOd/poNT5dTIOwsRxhK9/LGa4Evh
kszn7swnM5zvD6qUEXVz/c+WBn2GMQ0/xaYQIkKzbULr1FzD5bCNXvTMFu1mnrI+3L/HNpbBS8p0
omMOhhwY9Ohm67WECNpR0tYJ1DmWtErO9XI232fG26PWBvOo8tRNgnNUV7VidUaLUnb+NJEd4j2C
3A6JhVxvECn/uqvGPIrrt0sVr2rCoJJ30MbwnofaGxdyuThyCEN7Gbd9RMMrDQf0GhIV0wdfV5bM
N78iQ0Z1hiJjnsJtCFTCZOLQieVje601rdOZ9D5h/Ge724fDsYx9i4j7nmvnXp8QDgxkBNfd3vJv
oBknq1rY97ly1smkYha3NihnoHD+J7b6S9GDSPxOGEBGxDialn9zY6kgIRO89HC6x9bKitesQL3j
YjiRd/DRvgQd8Z7UF9eocZLRlo+N5I+gJBQkUt6fGBpo9MDVmQ4HzqU2/ZFlWKdJJQ2e8jpF26DS
I+XvlJvxUpbGpwgw+sG1Amsxjkcoe4vl7/VXpB+GdZYW0zkItyNeGUvf7vaR5HEbCzaKq+RrVHH3
WBpdDuFFtm/12R6+1Bq5CSQc35rlEM0X/CAgvv6Y1/+cjvz89B7sh7PFtdVFF4Uz/AgygGKCNz4h
WBZB7aHu+ODwbp0MPTbcehYhHryZp8EuPI4rmKA/Gj8ERUSjo/4MAOz02X2+0A89CHUNziSngfOZ
ZOSaDQjtAKQfePhPaWp3///1SYfXyptbPTvgJdSnvgn1MlzLdLSegAPN4UhSEDzJbny2hH1l2MzA
IMAGstszAJ5c3gYxED7YrwmcEBWd/5YqmTMdiXFUp5AM8/BLiIsb/oD7z5qyHroxMegsM/b8AY4q
O33xTVpRYxTxAgp/kuSJnTjbBPnuX5qlUmgDVQgkHwYlJzQqUMs/rz64flIbe+jF2GZsHG9tUnw2
tpmgzNsanpbdR0djJaSvSJR639JzPygCn4toG3Nzr8HV1LkLZy7dEeMsWRnuwUkWdTu4U2lan5jr
y3KGNMwlz0mZiWCHztOW5CA9UAvVsz5ha7R9uCXen0yR7aFmNZn8yXbfnEgiZSwwE8gzTRA8X4tY
sYcGpDebf0nIuWOuzsIJhtiEm+Rc1/7wX2rpeekfntdhzeLCauxPN8q14f3Z6ySpbYNlSGWo/UEZ
0edik6w1G3gPd9qz3i2Vhz0jZachbTIipwGlhbbiB3gQpx69E0REpfQMfK7HwkuFDhindNuN85wa
7w4kaf+hu/FMoXpSjx9nStVlVsdPQ3vHoJTFVYD4n0m6oa4VDU4rW6vRcgtKJrLRIGjuud7v2VBS
AGN/3M01ysM9WmzbVh8FFirRUbxymgt0ioZpBSsw+v2oAywbvhGenl+HEzgJh0Nnxb+vky8VcQeO
DkQARG6VNDGQ4ew7oJ+A+LLR/cmXVkzXwOV77eTLRp9BviPp0U9ADVGwqBq0VcMpcGd3OZCDJnI1
6qG0ZEwwXkwXgSviYxbgaCh8ZX0zT1QAha2x7RKexS9KynbPzDVtTVsghqqS5KdBolavmyoGIKT9
Wh0pQwUUR8B6I6poBuwmMpdvaphlQpVvs9Lihy6L1eMycMwHipPDYmLPSe+yBi62UctBVpFtuAlm
mu/OkpOE/35wfHeZA8DX82AGaTEIa3nsAKyxvZNVLnbn3ZiTkFs4pQKn1ci5cjPOpja2CXkPokLy
yCXxpzVMTdKmnYNAl47aTfOFsV7Xh1pKZKzLpEwtOuyPvdF2LOAWbF3TT6NSEbzg4z8Cn60yIagz
BtxSOwffhVd914TGWWWxRbOIckGWb1eyvKIjNhgdOda6dcjoESxWXrCQD3numD0ldTyUaRg3Okw6
CrhjyWKwCRP/uir/pZO4mwLmBvOz2oYwhU7RMZCmSfZgimQCpHUWWTcKVG+qizOPFaSTp0BQrCsT
SUWBguMvRIxMkxeMEM5+/fg3BmCec5BnBHIeb2bP0UzGi06NWR5etx6P5b3nKa7g6LjumJ6sJln4
Bsz4qb8MNuzRKp0ABo8M9TY+yQ0XWBD0sDDWEKQMc/zg1AMx1WoNIWuXSE7Ml91oBZcW7ho9fo0L
lKALG0q1jMdsYNMQn24paGkdU+4LCW6u6omDTMcjY4175IHBJYgxq2XGLNBscGLfCFsLcf6V9btH
g/j0BjK7q+0IasD+MPssHGjdGxbIUiPcgGOnH05l/Rz5BGHPrJQ5rzGFamOz93G3BIOc78lbXa/j
Z/JefkT5QVgUE7ra7qf94FkoHVhswodjHj1yij4NG0K/G9lfu7PgH7VE7w1YQVsJTApfSNkovhHo
ZaszI6gKc3uT2LYR1eesqiQlGgZHGAWRbyz6dgi2rmv/npS5pzu02HLpaRyHxbdl85/pvljTeE+F
H08nhYmaB8KEA7Y4X4SU7uq/1F7hpv5NbjZVPKk6qrbqMA8PglF/qOwutVwzee7G+lqwsH6QgrAv
IzNgaA/qj1kQxgntQrUvWqmw1qlspO65z0ozOpD7VmJXQ1bk7AZYFjXEar9ClqtNZP8Gz2gHR/hu
LDFR2KA7HqUYhZzw+0y/N0DlM4szk3OcU5eZ6y4APCcW+MAEt/AV1wEEsfaWTxTxjxFmlVAhRuX9
ra/y//jcbOK8hxqry9YdbMhvhbOmi+V0w0gQzG1tPvBYpoT3Ko5KDyOXd8Ybw8cwEmqjQiQ8btVE
KG1UByFr3BXpuiDKhOZHSDsYKW6ozrQyjgXFXZaE1zL6gvBis5T2WNnjbByzPiLNFu3+Pgfol6yb
I7dMlc4005M5VbXSNJT+XS6gPW0rnQF8e1JtlIzP/coT1KGCrWsqnFaiw/8dALeyWKv5QFzfUf6M
NV8XG/l4DAaMv9+LyU+ulhE7gxrfAT96Dli3/79eC1lVAkmza3/qedAV+PujwrDKZ3YmF6PwEBct
9R+JgvkWTmS7AOmkQfnQOSzGx/RRbMCq8xmE9femJPvB00gWZ2zipiebk/ZPyxABs3TSroIZ+Cea
FHGzs9EPmjrLnitwSfFC/XQp4tI5fIy5CzawIIKbHEndbQV14uTvRFduSOF+Sr5J7YG/yhLEGTOx
9juBM63Y4Z5GwYxSBjAZiT6e8SDfmoR6sfxzkAIMwKgp0l+8gps39gtAlkc71Vsopr2mD59ejtBZ
BkZppDVsXUpBajrRdEUOghMwIOmOS6eX8GRDPqx8Bkcy/d4eGguss9YRB4+FrByjn6J4X0TCX12P
n7qdCd8ilLyV6jwCjfrbu+NAvPqhLizuRrV9UNQh5qUS6YWgfBQyUHnwqGc2E+C94/ZdY+v319lu
cKFCi5T2SYzvQkj1jHN1h77m3+lS0lMO3Z2OeBGSIdy1iPvv5vTChZzJ7LAdQ/c9zkpouBR7tV9m
MKNpF9sxLarO8fbalf/BINXi6Gm/bFgB8fEH0iLoIC1iOjBKKC9AupaGkfRvpesYgDmdLHOiiNkL
neguwc6S35kn8FKyjWmkdDmyqvSRMWdpfDZdNl4qFTFqq1TNhCpMhhmH7/bdzbiIdKofBmjtCwU9
MnvyF7xZgA9NYZUOhmePqNWPYaSdMdKjHLWNWECwOV67a6+x3jnV3mwwVkhy5u5CKu3rtOGaDzmp
6cnRmcwhZ8PwCNuQEpetQ+Th2ZeirTh+bncHcZ8u6YuO/7FMsw5gjdZA/ecU7lVN/cFvLYEI3Rjn
LcPsC63axmKt6kEc3B/ipRTW3O/xdKfQpcOHZ0T537HiTb/5b/8Qx7sgkM5yjOUXCpYwQsBkRuBi
IuDvepSqGzZBtmWcw9OT9UpxmIDSKRXERS195OpW8PzLbqkls8D90MMhe5GTvvIv+r6cc7lVUy6L
2jPv0g51XSIfj/wAzzdu/OKpeJRmBtuc+wMfRlmdOSTHXihnd9VMCHNPRzV/jKf95MDtA71PpFJE
dMgi7ARFwVbTinydQYpLpAzqSDBy8FCaLLReo1a6cWabaVCSdeaBnLV+gkYjhy7CDCxB55xYTFUj
Zkr3p3976wyhTZ6ZjiqeCx2a0+fhPM5jsyZlaPdoHKf1Cp+IK65BW+dSegWn3s81/X1V8OggcYG7
nI+XloUxVy4jGwNYI0pkLFxz0fI4TlPW3woWbehFg9PfAheuLQy4hFsPlviv5FmwYOkxXqNxM4iC
K6UXfHkDnvsR56uZHWAcLFSqxTl790cC+B/3vu20/aM9o19GmO0pZ9NusBL94PMm0yTdb6wtUdXo
OfxFhobhfDhV+wFKuU5reJPdp5Q9Yh3M6HcSGN/hguNWBOXR0iYK9IvjAI/Uiz6BCxXVstA0Uv6G
BBQRoe/g63Fj3RKQu/yAJW9xhPGAVUY2A+dAEPWs5TsmCHYFAT1GVZT3YgoK1XCAB1araA+LQlZM
nZLW4Njc24qAe8ohdRg4oKN4PebxaWs0ABcdGRKHVQEXtQFbuaDKE7FOnidA6pe/raeig8x+wX8V
AoTJPd4ggP0xgQaDrvyq9xcP9S5ncPghuH4/WnTZb77P/pjnG1GV4E4eDDef402wVZGlvAa3maNs
GEdf7y0oNeIcf3ZlOqyTFabG/w9JMEbKJs9zeFf7efNHDPusmDkCka6v94QFdapfhGQnxM4o7G42
eSQWBH3ZYmNk4/0T+zYE2M4lj2wlWRYverV+aa5AdkmxN2QzkOwtFVaXCq06Z3XX7TsT4ITb9pek
qAdrqm8P8hMB9h6PMaO2L9fVGy/aTFbBM2WTQzSO6bKln3ad/Yvy8ckuivyoOolHGwV1Hvigm4Dr
am07XRclFRM/0Km6aoqfal1pQj6Nh/uYpqNw7dcRvA3n4BR1oOe6FJzXfaH6bTt7ldUXH9xK/xjc
vWMFu1KBQw8xUGyIhkjn0PioklPpeJCqwkQy9UaMFsbYbWgUkwIJRcErwfTO0T4OnLvty8T/O9de
z3QsINWjVSxfucZM1WD69sfKqdXykUlLW8uv3ICNzbyFG/q3HRcGFv9cFm8hRuY/yB2fgavkR/r5
O3mecQbS25LyD1ZMz0CE7YwMrPpYc/oV+L64JMXWgCH4Vu0nKDCvKDGmDqwqfVj26ua2j33wLnSG
RBSszcV4NX7W0YhhoHzqgeS31lbolRHX1kODunHFP8fAuOt9iN1KJ7PpUCxrMTb1RML/fVpfLilQ
oquW1cdU2JgUh9IRH7PxU6W7C+V6KSsXmYrtg0A+pKJTCiwAjUczx51UQIYzKljpB7qZm9WfZqrd
1P8xbH1g2lZr1gBTvKa5kWvsAX7J6YlPtGvcwwFDk7w0AKY+Jse0CfoRXxpLWFnIjAMLWw270SD5
g6eb1mJud5eqvW9YP3xdLGIRcMYsVtdM2iGjjZFJAXQr4SOYGBSAUqkAzrXPyyK4P1hR33xAy2ra
5ZjAjORCLM/QbDgiFGWw0AkquBNBUfyIlRtsqvAP/XpZb6UZtUcHhIWiqp50oaFQoBrmWTchuoMb
v2ug1FeElHf8pRKPrK7e1to7Hj+9bXivp76enTOHlsQf89Z5CBCjUWxGyN3mpdlBPaPzSqewytR2
XOcv3moFkdzzFerz4L0nmELIPANtecqWgYWU0rKh9iMLlbYmdQfkTFW0GPJ87/gyTBmbukEdRFcQ
k3Pao+GceGizXV0C3p+1hK7ADyVj2UJccBR739M3Cjxhc/iOAJjMYgYT2RplBrErtbx8s9tcVtmw
eesS+vyNQDeAAYpziDzCVkoStevuDn16zKGtOcbFvuIBkEFd0tdkWWMygy++UXCvnLxiUI35Du2n
W2MxSpB1tcE0V9JB7G07Ztr+LeWevBZKbP/G70/nWxTA77f+BNryUEBImnwRRBZEfPC7XLdMflgz
r5aJ1QtkUPMwnOGzZxAen/Tj7S1+gBQeQGhqk44sy0DHpfqUYs17CbAdFt9OeeSZJ3PUvMtXEW1x
IWT9r4WSm0imfUJZXgl6pYmCyUINfkEv0OIWdGcMpX0f8UtBUuogvfzxCyZ7H/npE/nZjAcbt+8O
jF6a90N0TtklnmeZvIbCs95+zdB/cYMc5qi1aU/l1urwWry1ZuAXQavaE5tGAKrWOApM1lOn9E/4
mAACoouFXPrLNzuB3Usnlq5ru4tPvNu1/bCic92mepHAyVkvJ/BmUsqJPuaWrAT71WQCTrZjm/BI
tzPk2A5mBcSZsVNhyHSMXfE2fwm7X44WJAdmZVLH9BU3qxRc6jSytZloCRfr2rBD1tN5736eIE2P
N1ZXvex8V1JD6tdWQPLay1tvZ5LV3F3lWjevMXvpxkHGx139Y9O4IjuHAvHerbeTm2Mt7IWzGkV3
DjEmdOV5trBnmMmGGu+efXLYYIat9gtsxTdzEIOoq968zKSoqEEzAms1fooPnJ0Nc4vakCtwHG77
PZQMjYSCtrDdnrrk1oeIZwo0yO0g04jpbdOSaXLBj2/R08IDgTqZ99WFuiszXeTtEtVg26T8Ahw2
ozrgt49SA40PQd3DgrsfcsiZ0o39ecnp3HiGocq3mUsWUAmlxEXItL50LuZnqrteCeFSp1K+PjLN
brFFqnwSFowIUjRNPE0+DRpBXEm51rxRlbWm1wmX7UB3YIFDS4AevVKdTGJyidIBV6a4DrvIM3Bw
WrInjdUom8CP31prYFi69qln/cIfTGSEDtTyUdmRJJRtwzEdX2SUhrs4zSc6tsOodP39J5oW/msu
cNTyyV+n1tbLPLXSoIAC2KNvKLRyO4Z7cDQ0MZtko/dB2zmnOwh5Vt/HdycInzzoklJLfhyBJP0r
yhGqZKOUynUpRlZccVfwI4kEenTR62Hn+vW3b7/BDTD6sqgBEGbpwG4CRLiCqu+ybVBB8yqVm5SY
/eocnW9zgHbZ7NlG/osDCLTFvyF5QdUyFa9h/xLSZ60UzMmwAz1HyrbWOuRPtH1pVMjDqWToMta+
7Z/O+yJZYkPJDhcjreL8NRQn/blcuqfMqDQC3a9DOENozwHpbROD0VI0TBI6DtOL3pT2vtguptd4
hKtq6CH5+SX9RVc9d5mOtk0g9FtT5XQBXsqvpDnQ2KNx/S9Fg1epzoRAFoxlFJfD+nAWC63O4IGz
pxXWkNp9TV5iMaBnXNmRyumtgrlnFE+egC8WcJNzuZa36wiA8qR/q6gzLMNDmd+nNLrg4MWQIEEd
/teGxm4eh4HZXH1h65qEOUWxSVPdLptzhsnHJpIvIqLsdQ6lLZvKm5Qk/QhnYbjMrqsb2jsmpS+q
3aI71K3SsR1Jg+0/+wBYTQXnptTB7zx25qAhu39VdsrQaQZra/LZC5gLygD6TV6AipXPlWLD1TRU
FsSg/CuTxnZTnTew3Gs8hCut1uHIiEZkT8m4oddHNdtfujdSczjRmU1PUm7LsTrTe0LuA1MNRCVf
JYjzLG/CRajDAHpGm9Y4StSuY6AKnqWG6iFDMwy71sw/JGHw4r0hvRtn4GvJQ4FQ3FCEp52FgH/e
uhM0NO3kmV4kAR0EXDwToUJKek3YgSegAkRqlbEOMQpdzY0mpw3UyTMV4GomUnOlezrs1LIFMGpz
g9bAjDLdQ4vNRdaTBZoBiHTBm7Pw9nFbyQH/4dNP/qJb/d4jtVVh24RFpaoeMCrf3oBsUP/Ay4AY
4dlsTVRdVl6a7SRXzpIpfk4OX9rnNl8LDknopOUdLM4C6BThxOzmUwILqKvYTsO+aEsB62V4i0w0
a2PtNkoBHUpw5BlUo9BPmzyACPWBS7sJH4FgzVLR7fC+04rP55WFcLmdHSAszSMJnCZBwtCHjwdB
YWnfdQHLwl7AMYLB2zgfdeG66BQXmXBfa686FuV+gU4nYNHKjGRVI9pkIcjC+vWl8Hm96R8iy3fK
YLdyIw7+sGDitq9WabyknA4n/EGvi8TBxYyjXqAwo5AIFpgFAfRg81zDCm5SUVdHN4B9iuCvaGL8
oqHEPoeFxx7081fPZDXVqcbCWfExJ/jOrwzX68vhTarXYGUNhW6pDYo25GgruXywwXV0lInwmJ67
Di9uJnVG1ZitnaVdZPIDqX9eAJ/xGP0c25OkunCLoSp/6xNNJQmRVlPUlH5oXtFosfuRkvH90HK2
qjwP7TQqFm59MWanUFL3obZEA2YTAX3JCYLod/LLzvSZ4iBpa7U0NP595Qn2L0TgM/8Xsmvl7Cvm
LlBhxTZKWf8FeTcLVouag3aY6RpxmFJ8zB+Lkim86oOhrYmeu20JlicN6Dt/XrM/LpkmfsA69Ngy
HZXrtln3WHSvzgvzWxw0PmUjkAh44AYZwkt68Jwx9sPQsUslw0hZzDW/pGwdRK8dv+OkmlDMPPtg
xRixOyE+AGtTWxfQR8DNvvgmwPgPFK6RJQ3EUguP7TUsZraPmAo0tk5vjs6XHUmb9zCKL3sXgI8h
5Ypnhk6IMQSyGdGV5LgBfgsEIuMT3KjO0Dfz2SifsnfHcJYvPohDu3yI3ze1ZgZ99gCMpDHaWBcP
jbgzt0ZOQNZDEFWo80QdXTM1QyTmNSDrNZ8RNIaBOgwQDxiquOvoHhe8UUnSM+8mrnD9MBJEzEhG
NSValNMEX6QfDFXptmAjYKxuua2h/9M/krkaZ54mVa224SKonGMd5iYDSsduaBgcLoV2RcND7dsq
150h5CVTMRA1rSeq9W23v6JrLvyUnX3z014Sk1tnPH+LPuJNeJtKTp1yBeF5FTLJ7BHKQAZaRpMf
pn55DK/LvvL3ut6ApF1oagtt7KO9lg/RLQHSqovewVhXDd5/y4wSgP8C/cq36IoYfis651agnd8O
9dIUF7ZiU1k797aw53L23da0MB3hBp9qtq7Pe2rdvuN2gMvx7Ath5mL3jzyVUIwWvBVeah6jocBD
Kl8AxyqmuogIzhPV72eZoR+eytJC7yPc2sgrfawXOWh92Mag6tTIjHjTiY4rpzb4yb9kzj4atv4P
eIphZiKbhsV0p5JoywabjnGosfS9QD4u0A5L4bv0QeacfXyFaBMstOkDgAZkqz0/AACP5HZF3kPM
gAOnR2NNpq9SojfxwBN9BRxNIudWex8KIoN6KwaK/9PA2xtQIZrw0svzSYvd1XTaG9TVI8So8+7w
BHhpqeEmvxCOhMW7XWVR8tN46AwefR7u095o1Ha3BiHgRH+88yFiPCvefnGrPM151fw3a3+u7g9p
H0drBQi3Dr++6uPLsl5bvLlhA4a5F5e4m+/Z94VB+AQlyKoQKiG0Isju8R2j8ZnHIrANZ/ujRY4d
BMbfbBPv07dYACXeB2JoaKyYRzTzGkn2o6sBzQv74f9g0NPLkkzCk9g5zTYMXW/tKyFjZQuc+c22
Co93HekrkdhA0p3zfSUxhuTJXAQzJXrJzeYj1JrJUUfEFKvzGyEhN/GK8sDBWSFwtXCtdU437rSg
n8pSOhj8cfKKpq2Jei0DedREXoov8MXjino0uUCTtzCypi8WRe1HIKYmRxpX8jlRCriFtBth83Vq
M8YsmnCNn4LDQF72y7WR8SJ3lSpWCw3kvC1vAfHWD2yWzMwgapH2Oh/v+T7QpSU65eRRLhteYqqs
yxPCv0EpOKG1v+KmQpw7rl/aolsRpaqqkixv+u0htadJTDPoADQg/S7IAzHLHBLE3gkZaTons0Hm
fRWS6wN/j2EBvGxqPU04LSRnjILWi5LgSKJmDYxxKvj+/mdv0nvQdCV6umZ5HJMrWRZ+xEQbDL3m
17l9x0YsH3vlpbz8h7B6GcN8T0G4PA8ta1vr60c5TvULmU1DpqJzsu6/M0jWfBwsz0okwiqo2bBj
xSefFnmoa3gI6e7bqNk+8/EJyDYQbWjwS01z4zp4Y7HazUrHKSlLeUcJTXipL3BzmAI94QjiipEz
Y74axy35YhMQaR+H0o9bz7eMKlTC8pp5Na7MX08OFA8qPEZa+9nGsyf0reU6UkFaG3oDgb4etK3+
qxO/TnzGAokRAY67Kw/nwAagkGdaU6UjhASy+9atc3Vkc1McCSH66rMa4IbbmcvLH6C/uRSOJ1zq
ScViPRoZlyhEfYemDBxhpNT3ef1+l5KYkgAU0vogrnmY/EOeuXSNQEXH7iIviIELhIDfHxbfWjHx
HJBZFP3KCChxwoobstr1G8P5tvDOm2Idp32HuBIo+5RqdOjgew6RvHTiVjGKEcmYbuuHeaKPP0IM
gZYm1e57fybmn+MZrzutLbNLaqnvxBhflfkogD6kvBNGaMEV+cmN3Af8WSy8fx3niF/lZpMJUNxU
XRETrqRE8VHV1GaMYGpMioFERLwc1jPqbMddh9ytJ4bpAKLNPn9BucXKIhy9hfethWs8OBHgh/Do
y+5bPSt8uAf8Y9NZEYns8OiVemePb7lFnPyYdTlosU0tZ+k3l0pQbyiSVcATREcqOBzY/Ugwjlqo
ar4wpFLTar1NPpLQBwn0gX2v0HPmH3b+2k18vtbOuRaNgdv/4EyX+s3db/3YWCa/atwpM9Ku04IH
eaZJuTUVEU28Mme2RS7SpQ7jdWj6R5dBADzJ50ZUIj7iFikq5l1T4VFj+HkQ/+64yStSad0trVQj
UKQuOSadyWtvQ/Zq3Vuk3kZJM4WO5IP8NuHxcHA5LHKnW5BPSEfLzG1xWzJbVc9ppyh1CLCF+il8
UFBP+l5Sbrin34YSZSSLlp6xsaLSE2VuBiCxvHINGUn9vG/b8nbEM2k+UPzPlN5SK/p7koOzPa9d
6QzonhnIgmdwcX7Qa6FWCvbdK4b2Yv6etbtN3+oxVKvNXX6UlyF8uwm0gYP/KiGh3hhcqEfmi78v
lPqzdrMY8yFoo5lZfqobrqjOGr0zGcSCD98SFyW1bNdjIFJE7isebhlrG1wU3YDoZDR+bkC0/6uB
Q4jmBjlILTPyVgOUdYRkYQ15k3xW+T2DfoVKY5It4UmspSxKLCg5YzXJ0wCyUR3HTTy+BK45VbJ4
rpGnEs5/m6zjvwOcGH/I0ZAweaVHDUXCI/G3pp0UkTvhBCVwEoUnE/LH8Bf1NVHfSS8q1HsEQrik
mK+R2o7tPXQ8kkWfQXX292S8Rpn82RGJIlRrP5LBhsTzEqCu1bThgRc9g6Gp3OZnq+HaJ0XC2mGt
1czAw04L3+cesxofT2OJb7XDklQW170UfQRRHWK7gqvlKmu4j7Gxa25UIwFsy+2+OfkPfBL5b+/j
rhsCUEOP8l6zIEHJaAId7MRwcfcAenLO74N1uCJR5LyVqFxqCvTw5fAkgqxu3wfHcrzU1ZG4lmTp
Y3M5hcU8E1OP4EwSJSEvVBFH0Zxl0oF80kFm8HbZVIrWpQy0R045/eJ6Ugb8bhosJ4BwZMkrbrcf
FuQk1EU7U4xxNTh63W2BV0+mIHcvPnhb9Bgqrk5Jw6jnW1jDh4TK/qPYf+7zolIjQ7kARfPc6y2t
1DQz51lO+N0twFFnpKiKiEOhT3A2bIXYucz0Zww+prfyqIXgBkr4R0dcEzp0+02+yZGeIflyaEGy
i/1scKxArgM5/NWDnkHNSftSMJ+zVY3uhldRpQODiGmYkyrt7jc1Ti9loCvHhIyyiSVAYotHi6MG
LKeDVhq37gXiQJ/G1pWfniuhkqklREnbPvKVJr5x4inmeFrJFBAzQUl5c6W0KfDJa6821uDrsM6V
1bTF/eZegWnm01rXyQCNzM4BDb02XBLhsFtqtfXJpjo/8ivJ6SILRzddrbPVOxcOoZmJ4rDNKq8t
nBdVIIRhUTgDtpWq02ySGEHZhnBe/Z1qSeOZwc6xEaxL7BbTo/pE89858GXo7LF25kb1KE5hrheP
nKGD1vgWTWPXQQOwy8EbqzzakvqsgZTuraqlsTjanpFswMn12PHQy6SDVdB3XMVDuUSh1+4d66hj
sSIXuEWT6u9KjAcwKrybzUjEM5p/B0amK6xnk/QLFQ9sTT240sewkAdqdxYkMQbSQe0ZDUeT8IGB
TGI8nD64LdX+Cuo5Hu9TiRqmq8WBIWOHV6AGrbc9VyoW4YZABm3cn0EeiVEtgEx5JFWyxqVtK5Wm
OaSTc2nrB4F1oMnb8ovZVmtBOamboq+4U1FtrD/IEAXLN3KrGev0l08bS6GKfYxepOfzWUUuKHol
5FqZ/UmiCeZXb91lY3gyyq2qQe5fTkYWJd/llYB4seaEsPE6DM/jjqOX1sxll/u7UNPW6HQtRoD4
D+z63yrgiYSwTP95UgqTCsHAIDS599CnGWLfx4LLkve4ZKMxIFLs+hooL6gIWJKPICUGyvKEhULi
/HWc95gdrWDezyGMrmeXCwtYe+S/zh216zQHIVX7XIjFF4zmbHbVXlsD1khBQWPY+NMNNoiT6H9p
clbKlLZM/paL9A/32m3MP11akxOx3REXpmfmsF7vi5bePYG2Pn1JB4iIVSZj+qJbZytR5/fVPLvu
1I7OfIgWW0afEiRdhmbPxi4ZWvjCXi08yUStYSpegdigyhblW8eS6LGoDkFGNL7eR/WtC0PJEf2H
Zm0xiy3yDNPn1A5ToS+6xDF0reenOdDCUK2XZa5RxKYFnWLuvSeKhic6EVHV5wpmBFVIjplBoG9G
NuVIdEDk/9njo+wz21C0NMFmFAbop+NhEW5VDrjRBGKvKQ/v8smL19ngG37iGXnokpxPknlMtnFs
T/Mf2NeF6SzRH13NfpYe2NKwvZ5fPkHi3loK4RdQr3d2g5ST6ZY7wb52piy5w9zByg0rfpL85AcU
kBhL9KHfEZFpLhMDyGv9DuOit87ekg/VNv/Q2AlGSPReecFiRQmyey+4F6qVpBoUTsF+nmo+J1MF
BVRxIg/cr89nrRiGppGjZHvJrB2sILiSWqvBM38Ym92rLpSEJN1iUf0ZtNJOooihUWDbzh+RiKyP
nil5zxoAnPprEi89YRDduUH9pC88dM9U4tyqcPuAUdLFoQPvEqNsVqoOSxwPYO/WxFoheG8AJkVx
fmLURg+zdgK/zQzQnWo4T8zn9ei5a5XZOcGSSjEn0mhj1PvtwTA7JYXaWtXvEJ0gRunoQTjhVGUs
l3YsrQDIImaA0Bz8usIUFe0x9//sseMRb7FGdPItgMJ3MY9FO38EAodFyhufBFiP2sBpMMj2kj+r
IkvCJqICGucmFo99Cunx/tyevEUNeWgNPK9ApZBZB3ISdGywTrS9O8l3G6outDzaKeIGG5S0gMx3
X7qa3r+QvXODnHJRrpdcgkvuLC6ggQFKYgVoM/qRMvhg6lWgpJXIZXheOBbGkisYqCmcw7mnDgLv
rieKP4TLkiiDgWaL/XBFLCece1aEbpDXbKKfFzDEOApOpQ3LvArHWKxCJ1nhioUTMPMbvet8XATB
w+z+scT4K22eN3HzTVGA8NR9ezmloNO7ZQKvTxM2UHw8nbSm/8pOSl8lF5QjgX2w1AFjptAsS3RP
mDZoKCjlU+ne2haTz9MHyk0i7XrkeoQpT6HYanuHE0wU5MRgS+CFmWv3gx7eebDlu/nEGxrT1KZh
TGZ1O4dvZDS2QmbsLYEXH4XT0c/rEZbxNdd49TzoYRahh/GaSy+VClZygUVo1K8H3o8Zq1YCK8s2
IKMY8pSjH6/OULeC0UTrF1yCRKOSNG8ud3QG2u/z1odaJYMnDX3uszUODYCekuyZewVTvp/NlHy5
3R0DMX6e7hup4OX+muTBiFPk4sYjKvYlQUKWE/EfcZfT6e2VJPJsvmVxD2XKqpqFadSB7WLXgJcu
zGFEwMJog2/g4W3i02VUGWDivshsmzV07tkNNKGwQHEVhJQgiGO4b6UxrHBn21OWbd1BPXio0M1P
wTjubR8tBRgvCmMTG2BmmwQxKrNlLViLcNC7JA15u5NUjLBxUfdqHLPQdzNRObmvlkof5H0eVRsb
ttLEqU6HpWwDAU4BWnoswu0jELD1PTLHbvPc4nY63aCUmWAOBJalIQ3ZuVyvHTxGow9/dyTllLAU
sN8MdBdzI8SQ6JF6vtcSNUhS3azTtojioANi0vhauxJYwUmqw50C8ZxGmhGnDsd2A/AvW3wKKSjw
+p3Yq4DCCgBq/zviPUS6++PfF7+N2jl7DKLuO6exwkMj67GrziB3pJLK5enGJTBEGeeREJQF1Aj3
I3srtHzK3lCtMq7A3zXAENufE+2WzeZ73oFhMDzHZjxNHSlI2fIgMttxhqYqUaktUfQ2v1VbSEwD
jnZEdsu7JuzrSct6MTviSlwBQGLJDSNOGW4OnwZTukzQ6OM3AINdmkG/7LVpRHNvvNHj7/lZzP2K
NQDW/LJT27XI5elJa045RruD6hUmvhUEm8NrGDEnr950Ce58J7o4EVmap9M3HmwBTliTqszxmHDQ
vADcKcUXSmfju+yMXqYET6VnbsoEY2Tg65oLsNfgGOhqlURaEG/2FkUB2NxutO+aqeEzLzSUL3E0
B9Xnv5Z7dH0XDQEfT5KzGqVOvDB1L6oW6Okc/uBXdgHr5as4wLY1/jhbBYtJGrlCZ1cwi53Lax4m
2PNMwCbPKLjoZUYi0eor88qMcqkSIcKS51Wegj3qdwUXZZHuiW80u+Su0zo7ioR091Szcdo8WIND
HHq0s/d67OaxVckTryA/IXPszYQ6bvy5c09UTKMLfIZpv3n+ml1ST37R2zTd1KnJIK+w8hA4AQ+B
8dekpC0j8JN7r9iDFyvTEaaS99d8ugtt/0mR4EbIxNVUECtexIcg2PWqGpmKt/mP8xBWy8hCzRcW
NsCpJQCG4j6uAyZ1sAGoeHiddWseueHgTM/Jvv8owuf3S3nHbL+QYbuFdk9cQ6K7xiyhsKsuEGDU
5PETG0MErqiRGZp5IJp2X0P0RiWtS3oOCi+mvIpRYmdZ8pzJnIpK+5k3gAAucZaEvFsHeI+lHGz9
b+ibF4b2TR6q2BWtjJ5GhHDK2plcbEhJFna/qyuYh90tO7tQ6ApQLR8P/o6zV6hPLwiYMXddxY+t
gjJH0v7JwtlDg0V6BKVTrVpCeEF5i35n/ujJo9JidkY1K+EswxF6NvcsHQaQQMzDjKAqEFfvWrn7
rBBHMkYWmPZ/MQDJ0Ict7Jv4cAW+SkljyrWeQwrN1ekPjLRxu8o0w1+ewhCNIyZ9ZPcVftkAKWbq
uxMCO8Iqkzy26Qp+SFu0qW/hrFzMg3UvJeiE9cOxQ5qch+Ozc7zXK6FXD6c3lS8f/jqc+upPHV02
E9WtgwqxGJaHGSBGzazlFyKPbX6o9XUVhHtA1U4Y7oZ+xFghfuMt7iTUU38apacsgM69/yuX3xcf
qi7K3idaTdvUtrL42ZpXvmjR4nS1fklZEKzWQ6qC7+ZHTlO1IBwZ4XCayj6AP81SeXGp7GE0xTun
tq0NpCOoqvRsmmeqFGQGetXifMJfuInPMe8yb4weSW9PB9FPyBRnk7RqUjiGOdbvSKZQIqGTdPMt
UlrZe3SPpxqEruipKa6nCuOfLGYpZGj2w7nYjr6o/DsNAR7VfwkxCEjSMSOHSC0TJ2cH6W5SaxWw
oQrnX/RXA3R0poONqd9LOCCJcrDPVPmAfNK/BgXvE1Udun+6RqKF5kiVwabmOiobBaut+sUmFwww
u5TPBo3rSSSIXCVcQ3ObaAwIlI/TZMhjBZZ874uWQ+pqNqfHuFwdoOxEQoUwAreGfHJF0VWH5RZ6
M7REUoe9nrsR4mji+eyDWhLWkedIc+Yrn7n5JBqo5Om1LM9Avq7vETVPT9iA/Erzi8pj7sBB/4Gz
OYrGf6DprpjMuqmMF4x0b0PlVUfyArEA9KRgTKnacKwbaQzL47c/ZlRLb6K6kkKApIWeU0KabJ/Q
DmsWH8xTW6cyZY7X0pYAyPOcCZ41MEYwvbJgoJJLs3pVghDouzhdU1xnTpNEcbETqC+vw3zyJjO8
Y23HopyoJOd3cAI1Jl0CKaFNHkwm1s06TR3LpSVWqBoqJ78m7GVewfCwfAr3r9Z/1kmK/qS5N4zp
1oVgsVGg1yAvJSw1jF7SEHCBG6Eh5o4dCsdPszl7UcELx1yCcj8fUH4MyKAej9rGeP/Xxcb8iDAA
CeDAdDhSoGMOxtuvtL7P+AAnKlpuixybQz5jvcUWp6x9Ea+N9rPDNUV0qIjFb4WTjliKIjCCW12d
54hLOkb5In/0pCtQ4ROZ2h9rjaW5PN9qjl2JEnk5i1ExVv2IyKeOPhETAnEi8nz3/a3WLquxAbsp
TfJmcnFSEpOM9UqFfeIvmqZ1vw0dgoMZXphKu3o85FEM2GHi9hd/ASAT/EKF987i2WF8zYyi6X33
n4Qel6NNJA8zOAYqASHDXjGp6/QSQ5/Lg8cakBI/wG92H9RsG97WQdXOwrnwExHZ+ZQ0S4XInMA8
Uj2Sg0Y/Dkq916DJvhr79+vFE20M42fZwKPC5MbiQa/TgVc982TMawRiDH00JaskYx4FAs2tUAs3
lHxjTGm/PyQ/5chvBJcQq1ODkXae0i8Yqrqqt3xWMSS6ylrRgblCy3DvQ9kPWE2Oro0nemFMasxb
dx0tkFHZkLBuwnfMIbQRftudo0lFF5MQcVCBsP+JPKSYkqACiuyO8Vhx6JrCcG33jKiCf1cpAsG+
F8cyvsppnuIlCvrlW8PsPqlW9d7xu2q4lis6fPXX9JJHLE4S2UyGwbHQcALAAMf/xKjyv4hRkUus
gkWi1bGfUKv2+QnDuPubu1cNbu0Cr9QOS1JQsXBw5S12t272ulpcC04kebO7dufwlPY98ibnypQG
kqdz/DqEhluefdiq4PgGaNPuN41q/p2Wx0y46Sqlt8tPliun65VlgfWvp40ChgMwd5nSgchfI+/4
TiIIPt0nLUJ0cyUgnjd5tUzWwM6Gqq5c1aALVVjUKgG3ks/7TXkHwEIQyQIGAizhXat/6bLYLTZC
GM7v9HAPzEX8HYAKhQ2ZFGRSlqXitoVcBkbwbjKsrnMTEsgYEBeWYGjZkTxIoxYEmJVKfMkq2fdp
DZj6OVN9Bc8Vu4ihl4qdf8NfUCFn+08VgQtn5KH50vK/nqJeQYd5dfESrFwrn5WqQA8cI5y0doF6
uQLAwoeYwHuS40P3P2YMXzSlQxKb25mgAxVWJwCQU8qwg8uqgF6uuCIbuMFhK4rskM2GIXH69Mr+
8AsIksyXL7r5t1oWo2jFAoZfdII/qVxVwh4h/EB1pw8aB1Xy33+Vcke3ChR0URymrHYa520uaAVs
0F4CPdVSOxJHktQ5F0Qg1CNE2wk2h4MquulWjY8WfeYRW8y2oftQ4NFKEME9YCd4+M8PXA+N0FAS
4k7fo0rsffm0gxYRvw0tJMoPYRYnDNhi7MRY5nY3SkEcVMfdz8y8ejRAF7Z4n72UocgDETqPe7Gs
aBbjJEKYsmaSwQtNpB0sUgBK/lUj7WW01k//scBpRwCf9+pGiSXoKB0AUixjHVVAiB6O76OpJttU
eeljSWqppb0mB0g40lPI3aLZzh2n1hZPtMNegWDFGBOXKPCOq2eJhVBWhxVCI+IEJZ5H7RTkn0kY
mLBvR1sSMpUwTeIJbZy0OZ2fpDGs7AM6tsJ3HG2MpSVZ4UAyyuobWa+rXunaQ+7uPwTe+o7zX9uq
cHHGIaGPBn2IVpDg2qQQBROvrg73FAs8N9O9qJ5D+XCZ9k6a0KrKTdOtxt42iz93CzmJZTGmaSV3
Y7ZFMpiVcbtXbP7Y+TRuY3lM2LzElqnGXBemsN4OAFZE1hIShMsG7JJ2egvoQ+egcEG1oIdQeRRS
GkSwKdj676PgTdAsHCQRPWacbIaMnO4TQuVu2Z8hIt0zBx1zb3S6F8EDAx7TPFkh6baeLFDdjXXs
LlYK4lQePxOcdSkXlrqbfD3XDDRmx3gFFS3sZhwqR0ouf1vRnTmLk6Z+7vzijn6aYgV7vGEicFul
iIEkD9Va9wyRM3fdPMvzYy2ffEWfTdqJapanZn5XDUqF8zUk4q0VWyC632sUI6xxVLJX0kKUrM7G
SmLplSloCj5lQgc3lMXYuWWzEDeTMgGqTgwdhZ9LX3NUEJzNBstwuFLGYZcPLdXjuFiCXlLAaWkF
9o/Dn6rgV3gnpj99bcTzeucaczy+cQIQCl1Vf/++OWsz48xGHW0ILNDvPBCiFrRLQXYSjI7NXWjC
hZM7bOKC7n+XkjwdgaL0WtbIXnqxEU0XN/D0ixo9hujq0SWVz6clEU9/0bbmYCBv0SDn0rmwOKaB
2weFFg5IKUe/t8XX5un8iI2ub5CsCdyhyJb3KEpuf/xg2+4md/zw8m7aYsD0Rt1Kmz4NaHbnSDR4
lIW53flFiv8FqMZ6i+3pOoKMNFt7kxh7/O2+tzCnx4qpoLS3o3W/rKz52KDAqRRFqV2Tgxg9/4GH
pzWLIxrF1OmVgi517E0caTFybOqfM/5x2hfs0MMh58wRjl3UCKRPCNsn8Dn2wIUi1EOiXIDI+NYP
F1sF4ohIt8xEpdvYYPtL8QBt3wQK0aK135bXlmWUEXYJtChYnRZXxIIyuUprMB82XU6Htf60NT/K
1JEM5G35+zFCFkh4i1L6M127sD97JFkqg1WlKUca1r9V2F/LE4+YH+1+WMJ+iCOFjPu0mduzWlcn
ZoDVseCKgeO3U3p4nV/swlHKrKyVWPW/yUpOH/QPpRsepxH2xhra4YVXFymnW06phL4Dpm/3GJdg
KDjY7eveazMioQ1N7owLXyETw1QZTM+h4ssCu9yxwXeTdeGYICC6G3t4xYRCZShjj3NayZcIq7xH
lILtCH29Pz0sNBPwHmkg11Mlm8Y8WFVzgH0da32C8m0wtdtdQWXGrCpkaJy3ieQra/k8LMRRoXTv
Yu9o5tiDT0rbNiAJMBleOBRLWJ5H2ldVHLAMv91SK5+NbU2JUEsyYEitV6JA0fMxOO47HPYCiQtF
D1J5RIfTyY1Vzwo53FpyXuDqjRIlePPy4bf4BrmUPofvgZeEEVe3WzFdmtpSQgIrYA3QI5+UOJoZ
FneN5+0nvjer6+ODSjbGKDw/U4u6FihLatr6t/WI0In/se2oV3Fa2+SiMubw7hMepOkAhDJ5sJHs
y4GfytpnNa89d2vpuIjZtaLkv7clpD3UB1uF3K7HmUAM6nDRqEHMDdqo2xb6oitUOLuLsqBk0SNs
Bfn1E6qxRz0NybPTYa4GIRg3+XCD+hcjqji8ytZ71ZKjIOYJ7RIQGR0tSmd4NM26TYYv8UrUKPFy
6TicoZQuI6BWGnDbRWhNR1wExtq7Y25tROLx4cHOQNAnfPmYPUlU9oueh95qWQJQPSs3NPnqahdO
HS9EBv/2h0mx11bw8rZw+u41PlWYSLcWTQdMoOz3GIHNbyovb6vy5gweLvspdvUTl2IW+mrKmEvH
o5nJ/yHQrEuVnQ6dTscroPJuexq0KsKxseIXMuyD8tXeKl00m6Q9h+KilRTKK+WmG+MEIlzvcm8d
PY/DBV/NbmpTnN8zssnbeC4l56BdBQZvKfet3g5O+1VM7G5YNgbddH9UIJdBfBTOEF+01PzeNpAt
WTZaWKcpxp+QcIfFyg0UIEp9q1rKWHVZaKbQvdeiLiGNXdRIvzzuZuDPGC7CKEi5HpE9d4Aldxqa
1tmGiDNSdEe6To2jq1D6262huSuubZ8dr8bnGO6YKBvMfluurYhxNZstQc7WmTdNRVLGsGppmuKZ
N74UeN/hC29tGhohsEr7RaG7OmCMi/WDRDThwEfeJ2bS8D9hb3KE2wgYKc7dnvNP9ztAFFtGbB0X
Ok5+z+h9W+si+RsADOWWszHJ9crszlmWyoC6Xy0L1DkV58NPrtDBD8gZihHBHf3/SY/8BNh2nYQA
oyCOAnMmP42FpxJV0jJ5PgEph7O0aiGwOFmURG0wJOOpeSWorCxn/ITpmlq7oVCz5OPABWsmmb7l
cslMVGetydlgxsx7h3ilGPcZCkQyEXyiyLmU5pYKSQHTfhAVwba/l45Pfw/1tl45/6NjJgSy8rF6
fI6LOBcbdjLOmES+9ax/4bxkX17AaZayHxK6rFgyZiYDEDQpuRvAhu1hOt/BpA+BVSCZmETv5wAN
gxOg2knVsckf1LE0OAwRssNl/6dmNnHcMgSR68NYG5jPHRehgPC7G4mAH77d4vJ9dWMHdyzTwyGB
uaTffbRUU0xoNeGkPwVCybZYSPFLxiEXCeSwOufRegFRCkewxr7j7PdKRRKauzfU3tS0qYQ5dt7h
0B88U3tQHE64yPolBKjRBsR7x3QhQz91k4QSyZNreO93npj+HaHa7Eg0Z7Qkt4XXMyu7/ayOvKR4
v3iym+8WqCLr8uKMTZJ8PDv+Q9n8pzP2LMWVrMDXuk2Wh29hbd+DzDsWuoQpLLuWym53JBSeOkbX
sJ4hw/HyM+Iz9Woys0tyxSNTmagyhEwkqNWPHRYTxUXRtjqifhP7k2u2h5pyuEgup5w+tQ/ooIDV
0aX2M2crMJMMJ5F8Qx6CtWPvsXyjNBL8HVJ+MQybBK6EMAqivl0e5N+4kO2JkMcDSJRcVaJqWYD+
WhNcLytyIfOEKvNfMZ6eR+hSNSJR/NdtbNeyeLMn5FtH+yBMKSXy3kJh4k17zOL/IkAXSjiGuYvK
qnqppHWrl7FD0eTwMMv3Zhva9hWIv69YhW7CiVCUU7MsgEC3lGM5U8yEvSNiB5FMdMtHxymFV+VM
7a8AJ/dwCSSUCNNMUJCL/T8BQabnl3fx8ChGXQi0uo+dbZWZFCWrlV2MO5pjVZFk0MwWIm6XcWxN
2NUqFKTL27vz1iLVQC4viaosBNnjx8Fke5r8EVyiXsVAkoHvwwoQQq6x6AICc2PvLyCzB+hxYMWt
4eYhyQyUj+5TFU8xXu22N0dlHDJEpy5YjohQMiyhMiBQEnHbnqRAEYHk8qQN2Bi1HQyedM9l9CNC
nBDqic0HxBEWs3ijERoPWyXNQUuuHzwKJmbrf1OwOgI6LdICdjJKAjLPj3/jnNOvtU6IN9OH4V4g
gzIe7gsNoSVfklObMj1Z774IFkrrPjtRLzFPaz0bbwX8Pqn091+HqcdKKhD3gehNnO5eNJjuu1Hp
tqhoYpJnVZO5TOHFZnru2BFfWpE8GTuTGFwGXfetelHYvauUXcKn1egpCsByqtX1wx8eBaM77ZVG
5K43ImcJVtBx8g9PHDitK5Fx9kzt1OUro9+a0uuLWZg2hqQcusEzXBtTTNdT8k03WRPv0Slh2/1Q
b9St0K3mNuC3GPB9SCkxluroIoGzdy5KnUKBA3kHVmeYQfifFE89xyQZJ464tmqtsozBMoqqSimB
HBBzcc3MtdhBCEciyBL3zFZ5tg0DeEGeTtsdvnIilshNUaXkDYmMA3n0ws2A1qXrxxHs7/igTL/R
H3xkL0m/TMISQIqLhqJLoEhFK3LGREr8g+5yRIgNF1ZwseryZghF6JAf/lIfOTOCf7r98NF2niVr
OY2UqV7hQUEpmKntb1cHuFlq4j/LEsJKtsikrg+lJnCHDRS2oNTVCaZSlHCe02T9Fj2Rqq3jsCag
1Rr4Vt/oxUMivR9ZnJnOVgCS16DN87R3+S8e9Q4DLy5oK79OpSTmYA+YwBrU6ZdCpF3P97M2iKZI
7pxQoOQhlO6ZSJQZ6x9WeqYGIn3DKFFtv7eq8svC4JKxJt16ntdSbM0QouVMifqbEZZC6uR7RIHm
Pnrkt5rk7d117QxC3K8G3mVb2dhrXiSoXaWso363BPQRfyGlcEFPg+mJAho84TklsVits29Pxu7q
DANlfT7FE6YoexPjcc19e2o5164FQakZm0WfPD+TOkbxvyWw2RYUN5ii3YOcY8wt/huTYS9Q5Ai2
oOY1PNc7SaF8TvmKyhz+QHXFbHcxDjNdStPqoig5+MEZdC2Y+mLZJX2jCYHUhgtI0geZRcfXUjrp
O/AbwCPTX9FvMNd8mv1HI3PYNiYYTjozfTn0aW8OKNTomzRpQW08V2b1aR823JvNxRhCDazk32WI
S09xmkRpxpUQbTC9vCE3t5RcJW9QIrkzpYU7Odm+3lmVHIDu0skOlrO3M8mKEW1am/VyTeJwSppX
hYiS+eb2Lhs4kskKUs/472+e5KypFo7whl0efLKgsD2Hlc+UyUNsd3jH61I5BXM8rW1P4etxhYcA
kxMl6GexfVGEuiiF0nsWWpHZS/N6Ft43H1RKgk88GxoaDiizcKLlPnx1TnyegAxNz+c8VmXozTHC
4/p5UlY2SvDAvzmRi9as9yJ2DbUnbM9EPAd6l9rrlWKoQtLdxMVrEHXlk2TWey9Z1zWHUH4iCt23
4o6lD5o5GJeiAfRPCfrWyA6jtHianNKrdq1lthIJJL6VNGOTlbB4JOtonk3tuR0KT8RuZ1kg/A8m
lTjEYN4AAq9KPLkDhdKQjTmemZwtWY61Qz6MmVhJjCh7FHNyI542sCe+ehfg0zUISqF2zOb/tp2+
yS+I6K+JPvNizq4wjIWTbpv8F+Sg7ET/3dNbp3YE1KjbR45FjLZ9+4r872qlNzQ3qrLb2ir5exPT
yw88ZweR4BdwQeQoghuWI6hywozfDyoA/V6ffzC7x+AsSvS6oJx6mirZFgSlAvuraN+2jKGNgu89
tCEk2E6UDzYY7kjFSal3pb7da7/0zS1FRJH7JTuhSxWr5insnj3v7WfTDPLfqLeJ18JM//+iAXpk
jB/fdhOYVI7cA2aPIlI0FfHKREs+ztKyF/ZQcQmKpz2bk1gDaDjlkY/iynog2OKFJPi4n9ugI40N
2MM+ci7/ZP8k2F2NihC0/M3gjctNsrcIkbj5nkDXuJB2o80F9LKeZC8i6NWjmWrTQgcM8cWcX2LD
w+Ll66htkhCXWaGrh/6Z4XgJgRGyiu5mfjZpvhoSEUkzFY5R4awONABntU4sJFPj+tjYPGKOgpTT
EkAZMXOCvWBUJuSI51+UapVV/7Wj2mGWOoT/lEMcvVA8Yk8NbNPKX1rNTlGeda9KVlGyeI9jvlkl
SGO0S471SS5pkIELTDtl83odSzWoSwp2hf2dKANnTeaMlZrP6TYmcAP5PdTT1eWfs5wK/tJGXmMK
RyFBFO84ol/QQ+L9SysIH/NyetALFfu0edg4L9445LW9GdzOLAMFDJvM+D5ol8jIPmMpGE/nfwq7
QZSWe8KrTCs6hVUEH5taNslNQByPFY1/pFNGDzimI+GppKcr8kI/ExLZE7jMtiBIUhy4s9ouCgZr
wT2y8uFShr3LPr9zPOvf7+gnOjIItuXW5DEw8JUEYVykuiukdEaa8RbjQqcU2kqgxm97+6ooDikZ
9+Tl4Gxeyv083XnG+WJuru+9ZwaK/1fiMMqF22JUZayhGl5ha3TJjWxaE5QeIL5zQKIU2UCjMcJ7
ClxMeEAoN7oLPsVzEeR5JfyrF9IctyGKfHGUWJOJAgvA+GHbBp3S7tFxMHk1uzC+BvtZenzHE9U/
fjLL5PWz44VGFLwX3kp1EDR2hco7kkNIWGkJLf0vYPiq98+76rMZsyVBbrcCdoJWWes6H5Dd1RSz
ZiUSOLIw94xDtUCpyOyYA5E44LZzyH6ZmMOPWt8vbNIokzN2NL7yBwEsw/iPrslBDZ+Vikd1GTf2
fyJJQNQaPXIaMzYqHb27zIXYm8Ekp0kybnC/qYJ2HGW7md1jRO/xyZOUdFJyDL+Wjlz9nxrF0Lpd
Fh5khvtBUNItVjiSCaQdc94bgcAUyr+6bYjxzW10lvUAnWsSWYvew5/7o90nfAHqsP5JK6SHFLU1
AZDDbTEQHima7QEOjhFSVv6g4DY7DkAyd7hSNQIKRKRSFXOLcJKQX1y4FRb43Fowop9a+BTSFhYA
O+wRKo4C/GX2ccfoWhXEFH5d1m1b1GYbKD1kyaM7gcqsMRWZJGHRr/Qv5z+4RMo+Arwdt9S0BBaJ
zM5Pv+T3fZ8eQyhlpLwcc1ZseeNFshkqRDagV5t2my7g7IUm6b+ydbgpLT4ksXfSs5o0XUnhW+ZJ
s+wJY66U4Txe0rAfpMIfB/kA6lKM69AQICA9Oego9lJWsLSIjDhTyEx69mUNBejbC5bePv1+X4hn
cL2+BP11v1dDt5/g07W67Xj+kSPgeu7ewgk6PO+yTzlf5qBukYDuRk8ot1/rE/4kHL7TMuIIfcWP
rPJ3KCyu0zMWrYsYE7r38NMPKCoPCDsZTWo1fj2NmaRUf+o0kCMjgP2ZywnR+200ZwR/V2nTdefv
zpWh2+4yb32uIybhM2ZPjjERazr0sZNCm9eIV93e9N9oMfiQ2nRpc6PLhUxGqRUXi1S7PyeubT02
8fxNG5a76lpy9ur4p9OxhaE5/LbZ7vvgTMpAH52Anrh1iA1kSyEirglSFLB/vau/8hO2LMyTCWYq
p6ZiKeV43g63g/yLL65j3M/iPBbG57J29c9lHfyOtTi9EBgiS6h2sAXl6QptFVZ3xaSXAQ+7kfRB
ofLo5G2OAx5DbTFHFcBjhz7d8MFdT2u/5FKkmBdfU/y1xEe29VyS3V+Xw9Sk/vhEwwmLJp3l7hht
eTtKQnNer7d+v8gFfGSEbdD18HagRqwj/6ueLWwiTbjwIIzy5IEd1m2qlcMNmZVlIPTi251y80Fb
3+Kb/ljTp6jMm6/5hBgdoiWNqlD/LqaMkGkgzcg1W6Gv9VWYUhq/CUsxkduyhGgUTK1tapIzcjv3
fgnnmgMtfU03ifvwLI8q7fz+skpISV326XbxyZvKHUpHV7ESErn7JtmZE9nBzR2Rle0sr/F6NRSj
JIDz99Ttlb8AFv1W9GHy7UjQoWloglJvAbMeEbDOJMY7V75tJd3xVhZnfpUFVuUNfArawv07iSYB
u9ljND7A4APhhccDLSpCvsZmefelRp6Tr1wB977q8ztqrGhI1413PVRf/738QjCB+6iVSnIVyyaf
mUe6Aqf/lkU09ObkElS4ELyV06xe7KaGBywZ/sdvFg0SdL6Kp491hfCnwwOJ2oc26Fsr/K+Ana2T
dZ4VYclJBK4V8M3kw+EYWKGfTsS7x+547X/62LvW7Q9rVvCrEGlv7MSwlVEsWXHJv8y2ZJ0+PYWO
PyCKdmuiydgpj0hzguI0VioAnhf0QojNjO1TPkX5UKzYSezOxW2tAJpBBPgqDrAMAUEUbc9HvWBb
AgsWufxjrvwgLdZgjq0pHkBpUlDQ4vtXUyzeaTbkcqTpLKX4XQPmBqKxz0TEYpTCIiZH3+jVTjN/
cGoPbn9GeF/WZxaR0Rw5HnxQUFyfZBSrhWw2CTwciEWHHBAV6dXLbreYyd4ruUbmVZU3bCPhwTH1
UQs+Hu/No8tVptt5o1sHScoNXVGnknzMslRCCyY65ycSbAlB5Z4XXPbbK8aAIHSTZ33sm74DsD3N
lGe2oporLYyo6J6PmjvDo5Djg8wBhrWvyqdfNEup9EF/CAfdGaDkNWWvmtCj0yOKBAKtPHB3zvc6
9XZ3eZRIgqyg82CxHZcuzV9ikAdLci/NtIXiw/iiC8P1qKmEKgvrjlWkuHTXnudjn5Ne+c80KJ04
1X1YfultKw3JJ4+rp5vtyb7krtkgRgU9Q/QqJL2c7LmvTd7NP/6hWug3Zqc37uPkJ9ImCPoltHpZ
ln6iugxp25Em6c17kdODuL2aNyJ4ku8UUS6fXPXHdQUMbKbmv6Xf7kXUQZhZ9aEDwFgfKidLKDya
X2LQNfybqQi63C9tRCewr3D0lkeYyp53jKJDvIO+rXzGayS0KSyZg0kWmXNGnGhZTQp8vtNUjBLB
JHj4xzHbAWa33r3Hl0gsCBi10l6t2X6dtNFbU3vN/jtDEOW+5/NrdLIIuVKJbwyKj6u+GYsXVNYj
jAhheZb+EJjYXPbNXEn6MzIYDz/ZowukeMhpNho0/nv7OL0ndlMo5SEIXdnaNnZWCt6a21zPgaV0
eDd09ax+ZiGBPVtTSC74TQzwoA6r0/FxshXQoITDG2J1D8qT/AbF+rwVdKGAh/NznmFML96RkgHf
iUY5Vz4yVjBHmLDa+xKKimX06jJp/qEGTVMbh48t2Xz8UXemSdkyq4+oTV5oq8w6KFfh4cKqM8ch
BYZriYggq6eNtNbABjrH+YtROkr+qUdEQgrZCvDpWMh/kDDzfn8NpJkZOrlwTdXIykjyxC9K41F6
KiRv2+RGe7KpB/KRR5vwX3oBG3pE3CMrMd4xENk39ONa4aHPk4c2jjpH5S15hKsGnH5HoHoBe0kL
t5kCiIhRs2PS10j5cS8M6IoIEfuv39HDQQWAlPggngNBqrgBtBt3kP0f5IWwK6wiT+7tE8BbyOaZ
KVssu1Zy09Kvk73shC8ulJSrUfRZp/094wISusYeoXvcpiuRZW/1OzJ0foBYOhubcwMcg3uFEuey
dz4PJOJNdQXbV7sIMsGnX8sQX8eg0LzxCs5RKhyIOj3a+JmBMLDfXym/oV2k+cSzBFncp/bMjJXo
YXhs1OnOFE+drJPpw2JGW1ittA4+jQmEZVYM0Bnl62h/IPFFCNDFkC4Q4ousaWNMro2Pzk8/8zK1
Pf2wApixDDMw3kHaWQWGkLzjht47ujiB+uxuBKcj2NkH6AS+bEjkwwncjUocFBA9uqyVIseJ1mvM
rJA60n2hIifcNcTKrTpOnf+WdBshn+Ck0Pxop43UNbMZCh1qfZgRoEbX28vKoLBQ4ffdTdsXncg7
fNHRJwBeFICBtHgXwxDZhOijpg9DjkY0IeKEU23xLL/OXxEW3c/ipqc+SVWJ0yJ0PHaYgL65c5tD
lQKywNUJ+x6NplWJWYKufs+PGbkcL5hV42Cr8jHr7uQArb3DEfPXw/nksQe96FRvykO6CT0h7lgr
dU1cUg5aF8lkfuk4MXmndoyhUgsbOrq8+NYJ+TKMpKVdAE3EUBB5uH5YJB9wNFz4A3oRr5DhKlHr
TBJy54oidc5F6Rzfur+rTR5EwNbKmGONxutzvRqxrRc0I1y1WYxXTdNrvlOzXpXvpnUigp3PN/w5
UL/nOXAG6GgA72qF03KeAXRRZC5n68XU1O494FM7wsmPC6PSZ1meNxcxh/2mlww3W7r50QACyALp
Ex17BEDHkNP4nQ8ZJ38n5JB2VOqisxYtD40duqZ59jSC3RaiZ6ObM7EsHeENyTCk0pzGvm+oliLw
OUxUbaWXV2pOWOzFILh/bZNqNiPYKaztN64ez1J3lQ4Hwx/L/rYfAN2ftqdfsIinCkIFEMJxlU4k
0vbj+MO8IC0oMsKXJW7/DCphH+piekVMZi3rEZKe7/wQpzJtisPZxsZr8UY97vyz/hnKpryHfck/
XhuiC4GonCeZK4Zogf6h0fhsBmm+APtSOKMcvF1D2345+ETZLQz0WgnBp5uWs5WekA+UZMauVFht
PusxgnnOlwnMrOTg0vnMZ0Hm9KCOteqL8UkfuDcOlbcLflwZ7/kcXZ3mnjVrQC56u1joXHVwrwor
p9F3ubVoojbUH7zr5R8tpY8sN4eXlXCbCi4fDh2t4OYWZKhm0KpQrQUIdpf7G5GQGdSCTlh6/98m
LMG1QE55xO4MzCFcCwk8hAvUWjVCbf0QNcoffEoI5l+iTPB5EYnwKYAnAQ+ifh8UjYcIGJcSCe0E
OWpo3T7xyUTbbHzYPbk/+EI7BYYo9PWbLfnaxs0T/1mMf+5FBLLCrdwMG6CgNySzywDWx7Q2bB+U
QqtYF1P/X4eLKoNmO+0XWPoBjs1rKn2y6OIElgE9PGoh/dfGl9+KGzQLEQDfHsuvtQxGFS8adn1C
oXCn/aLeBy69+XngEf+WR7BYBkToy1GmTPPIpoHjvnLvvhu7+eEFvrgHd/Dti2FLLLY+1dG15wPO
xKnU2q7Kt0TyCVWZWL2PGJKS2Z70n5n2TYrZXO3Nx/sY6EJbJ7t0O2Xnnqs40JlZC0SYaaDRyKms
1Ec58Rad2CfvksJWHFAawmUnh9VTqdmL0rfLbddTA107X5tdJqMbwRn4u/hxDAWGS1yNnicue45t
3FFTHpFOh3xfbuINPYwF+ogCPNBCEI4WVpAzxk+KttepNgf411fP/3gLOjLUodHWBB+mhKkaFgYH
fJum7kQ7YrFkxhDZbJccnNQVwEHOoIFoP7OAZYZa4x3+rrocjrM0470egoL7oiiktTw2kGgZgDCv
Dym/lbCuDKdvUCzzg9vl9M/kIsMufIPGcF6zVdCLt3C4OijbuoL6JkMRG0e267BIbF54A6hT/b0x
mGzK7SgwI/K56iYS7ldnpTtFtEDTIyfj6UliBXUdHlG2LanjVV1XAoNy/4PA0hCIrLaQsjxBufmo
jeV25zui3PRkgvW7IMbLwNcCqF6AF6HpKrPttnQkVSFKEtmqscgFBCmsFswbRVMFg3KGPtjFE/Tx
6vxplVcLtxoUB/F6rV6r3088KaEbKAq2e7dRdhCRblP73UZfnjIMMfcIWC8C4YSWM3U4LQOWM7A7
7QfFFt6msLIREdRollB8wKoYc5/noJvOhScNS+tgOWxZl9reEO33hN7FQZGcFRbFHkoYA2vFqtu7
oghVLZ4tuODXZUPmAKK73i7m/f45FKei2W2CsHK3pl1qGTYjf/74wTA2yH5Kr56+X9zjiaQQAM6E
X6olVW5qMfUh7epQbgfiY/uIoFV4C+M0x2GXsCYkJUF9Fk9wXoKxgv7DyJkmgxac+67GZDX215fK
7G5Uq/P2H/AejdRCqq1ZsmguyX3ULszuZ3qhBWmJj1fJXBInF+A/1N0A/5G3Kn8FABNeidYfkfdn
nMAZwUDHJWfpRUvjhsnvrll4/vncgBlbeQjoLL+dk970gWUI05puJs03Wuv2hDNXyJlTJZ/yTsgo
CTH66TjG2MvphLsB3wfy7pLxXwDpcHS265eRUumpcwqkQjVG2GJJIBF7Wx69ewutllFKkkm8Z5wG
v0lPuR1Wyf7PmAmbgExF6ON0eUVbpuP7gMIY7dG1Mgv6kAES8LIZQtaAawraO+uAxEWqW/SE2CJl
yGNG2CPSSVHMAl1Lb73kOd5Qe4Sd45MkIzyBqgl40Q1LPV2aPAt4TLsCDu6Z60dew6Y52kNQzB1d
Q5K+JMpInQRvQm5zNiZGFg1OHZoWfcPwnTZA0tGTKwVsVeF08pCpBCc1go9Kmj485QZj7CctTreY
EeZJkP/kI8PNE8WbV/mhub35Djm4LycaoRdhKUO6EPeqNkNicbXO3rMANNu/Hg84+z9xfLwOPldS
z62TLEu01WW53KmZG5+FxK25fPKFA7QfxC1dW8E8Fn+Vvg0fMWBEq4k1Y+1YDitI9Ng8H3vDr+Av
g3FZBuyyrSxV96Dme4oL9yneuhRcYqY7SySDXvtowQxFYuJqNRMfjui9ewrRhO9XcPY1jzdye8gY
wRmbFlyLWygU7ew8I1mBV/w7wkHWFeTxRjz+K8oRY9lx8tkfVTkQeHrABXQaRU6Y7eTlOvilTch+
66/LQKPNKY7Iti7TJYBh6colYUrKhl5/KL9uEUrgtDJIFPSdzGIi2w8HCsscERtAD2RlJ8H+d1x1
W+11qze2FcTLzgDTx+3mTXQO6tQy+g2xyWz+9/2bz76sH6flE/j+73DuG1K9MCVSYHW4OnOlG10Z
mm4MVcRTwHEbuuGpZfSURPMmiHWCAIoNT56vhhDpTZ++GxUEponJekrGEswEhIufp5WxW7DPxiQA
rwcDlka6fzv7MQ28IPvVu5Uuj4sqQ3FUJ1DPM629Ld6jaKMj0UNAM48E4+sJs1I9+H4XFHkMXsLJ
Tegjca9596mWmu+FExdeqHTOiWtofamP08QKp4qLub1AGpOx4TT30c5CTG0DD+HKqXgu8RmBVdcu
kro4lwURNIVV1W2daXJ2c1w+wIgU1/Gsh16x6U0PU8YswPKQhEPDiVziGCInrI4q7odpXJBH72De
+Ixe7F95p89nr5m+KrHjh9ULEE634ssLiU+t7BN4gfGZTOOROzXpPsDWaoEDm7FSphdrnE4GfZxf
b/j/amXTNyJawl5mcKJ8F5/a0Kmg8q5V4YFv1b4ZLFuqlBGEjqa70ot7zAfbxumyjPimCzj2QhnO
47gnY7hCotUvobmA5AXI7M6evnQIugw3b8CkSUJ/+1Ofck6HyTNg2mQP/ERWPnL9m+BA9jaBl/4x
1rZOiS5V/27UOEDaUv5Cht9fo+vFQlH2yoVgimVlRqxUVfiWEuXLcu+3CJKs6q46KGFfd00mN+vM
39m7JmdO9cle1OuGcrsUurSdwjd+trsi+sINIX4utmQUJMJhLNoeMnAv6l73MLMhfNb059ndYRor
T2gq5m2FlmPUmIWNTIyWm/RZoldSgiWJ8TgctQDa9U5r82BlWg5dn9ZPECafpSJzO7bQlzBMm4A2
FhTCdGZgddJWOik5g++C1hDhSn8vi/eo6WnPMSBUGHJaYmTnrfcmprATBWuzacmiOCyvW846RhDs
JsS254h/ZZy08XUkVjpsXeJsmimPvpwUoR9PnDGN6chkaXUTlF8y8PtV2Z99cLCtJVYNatPDo6CY
QB0zhr5/vK9fmtQ2zBuaXmrTHaKD4xG7Lnm1ObTIScVfOTBhQUUVqN5wdzJ///mhTuqK8u98P5AA
A6z8l6hrmWFKtsBE38pGXbNDo/eGkwEBASi8YxKq4xKyyLjcuJnTT3ZJBIHYB1mmn/QrrSyZzq/i
eb6efElpEAuj8wyFTJIVaWCHlPF8g8IRssbQ6CVFVTNN3GANi9PbNUHZwhRTldHxqXwcWVf1bUgs
P6Y0xXQ4XbEDYfVNuj8PtJSDKgLTUG5H6t1XfoplanrJ7xzXLvQMsHY7IjpJRzFVLiZzAjvSd3PQ
807+xKgWa36lo7o4KLb52CjrIgNyo/4KKxK1W0JqbQkuldHI2OnfaDTdCjMXDHo4R1nFkJeSl1BU
tt+RL2vIUBGd/WhVDsE5uhMUapUv9nL0zbTsicXOarSGfDYSkwfgpOiM+WYH49htc4jLtTUbKJMJ
wrKfvx+Jnl6zg8+4OQ9NxhMkQhnmYR3XMMVXVuCQ1ejRpmvg68+36xL2hxmOJVRUyZJ+SR+PTHDC
agpz50tWy5aXcAAqy4MqgUbrBIVJn0p6C6uXrrnloaMjiLo2XGIRP+MpxSrXTM5HEyanHqUbjTWK
9JfWp03Kk2zBaO2fGW5od2Xji1Pe+rHFO7unzKfP9fPK6Wq23t9Iw7g+WTBc2q6z7/odViv7zGiL
WuFBY4K3IvfWN/NOq+Of6I+tQGCCuCYWPnllOEZkGUMlWCtc6qzH00iAISq43lElxVgdm4DyuY2i
yTaHUCd7wEH7LAITrQlNKm07813HKP4n8JnqNRuUNHWiUJAypiOMjrO9lr8BBB4in7wws+Cq2RUb
ok05nsQhO+qRkDqP6r5HNF7+YW9i0g8ETupCGgpsU5a855mrUBSYX04CR68aHIsRFth02ImUd4QF
jOWMg4Q1Q/jPwZoL3ljADDuxDTe5eyQsl/CW+KUSC8UaFA/+sMjFbXay6p9i7C1JHXuJdUtt+0oQ
XMecKa16/db37jAwg2WqblmbcxbGlJF4MZ5pZ7GPlDWhdIWmVsgSjwdVsdAjm3xRXVyfyggVRUam
BTGuecaRE1SVolvAfyt675JTAx26EZRyVtcRjudVI2Fc2450lNfHHJBSHxdj59OA36sxIkjAfv4N
V30IUwLwCG9EcbbLsSHCwJV0jow9IMazRpaykI6tv4M3K7bGnZLJwWlZ9N3543Xf7toZT/pjVnyx
Mpgo89N7ateLZqH2FDqLHzwFbjavKGfjA/uq8sjdK4UnwWEcBldl+89Nl7/w2rYfNTk8nwVlSVXl
6jbzRhvP4w+kGH/Odhfal9tP/8xvGvImybSUOse1mr1iDmlJS56lvmx5MOTjRv9dqpIvVos1YkY3
Evaw15SnRfXmiXX7n9of2PVrgoKUcJMiK7B2FOAk9yUdmVIwCCK46eMQxod7TamboH38Qiecn9YZ
sLLoxQ+Zl9dfwCLMzOpuxI3rkOEpBLYkykZkUjgsDTFbXwvwRXaHHEk3/3Lk1uIaGad5dTDpu9tY
oxttk+7BXyypheaUYDwq2OqRXdE8/fXBmb+7kEJA8/ZmvlquGzZDwe8jI3cOYUESbSBq32fnNFnw
L/4L4zqKO3GpvMn8YDRAHn0i4cIn44cOFlxbu+vZqTjsEDI1YYbuWOSNTV5nbDYdMa3mCzaI3TUF
5+9e7iaEs45svfxyVfv+7JnTrrwNyPk49K0dqbuyV2TPKhAGkotStA94Vb0qpBq7OOx7xjvz0MoG
nVFM3Hpf/P3OxTRINv0PTADt5x4LO66gRobS7oJU45V74rDXTUeXMUKQrowy0n5nLi9MuDk1UCPq
CGNs/BzQ8px0ntEcvR9EoBuQoljXSVgfnk/upr9HUjK+Vs2T15+Rfby3y1THo0WJ5CTX2UPAjx61
G14LkX+s9LwTMMILuDgQe8CcEwuedHxclbn3NvVcZtKWhoNM7U0LQvRugmWslrGOjxpQwZVi/Un3
rllfYRbELYax/pRLhEkhlEE71XK+lOoFLl5WKFZxvxfSzze2jq8KnuWmqASHAWsIZRDa/T3QAbzz
NAsLuJWJeuecxaPmnV85S8AB2UtAjWc6UgV9fIxzxvwRZKg5t2Y6Me87ExWs7GqcSapzsjRDsRr5
tUcxS5+JGHnhyns/gvi+URUeG5VlnVq6336lkVG/WBPCHreWBgJ5gP/agx1gWQJ2uL1Dfj9ZDRdR
EzxVzw3cUluD2PkUZuh4oWeiIpgC2PhW8ggL2KfmLPbg1ck2YuJOKYQ442qGxq1jgqhAAashrPmT
/bCGcrLrLrfUhjEdzdGnp33X1VBNMIjrdUNGZwVPPsJJJOhLNNdApdJLQNlCuVsz0niMH7+y3SNX
IvkSnMPG5WT1TDJTxs/tcw7p85CiGYVfjbhbG7GzlsoKAZUnclDFnXQ9OxxkYIBCsmL0vCvnxPa9
jbSUpO/g0YNoU9/nvcvA1H90y3Twp3K7ybPfJtMASrUoZD5lQed3PiFiWwRRJUNFHqSXOpCEC6nK
q55rUlWUR9ayBgXxZ0FcaRgd4/mH+V1miRwn1RtpxF0MIO4zVYfTh5wP3cS4w9Jzi/UafycQRxSw
nf10Q81btNrdD7bqsb5RGkavy9nyIBdMPlGvYgt4Q+Y102GFzrHKmoA6HS5fl/N+pHDif6ZxRWMf
bsq1eLoo+6eZqbIUdAu0g+N7sKwhe4NQKbcUe/Ej0qk1FBgj4iqbATFYVhM/D05uaZbXp4v29dN8
EJnToeQ/b2bjgyZrxoGM34hfvX8ePhDAlFbIwIrqfi1j96sXPJOSFPlPR7i9xV1VchA4iQdouQj/
oddC1HcNrLIQe48Xk66Nrg1lo3r1kOQj2bnSGv88yJa0onw1L29bXg9FphqnIucnzmDzU45qZrhg
D3WNjHiBY6E3Fw6SM5tcqZBVa2GDsXZLfBO/ujTEhGiQuLGz3tqRKb2YIwLyIrDCSEsnp0Nc7+FZ
r15IkerB/0OM+zOc3xMKvKBzYDwjXWBGCAb1+Y4WZnVZsPlceW52RKE3k3l2yGH8E0QURfSbROSd
+NOr/u6KvtVHVSFN9mbKGlU+Wnx7f9LdLS21zE2D8ZY1FY9JmzhPL5tCEijmL3TatQTYSVrDh7AN
iKOVz+RBvQKYe2ecrhHEirWiaHt19H66Caumpd8VhYYkhBxWgvYFcudib3Rp9MK92Lmr1LZHJtb3
uZf4njrxwSW5fbdKKe/pHXUUiUGSXkEPNiGORbT3llLFnjuaYnd3WKaxAYuePXx8jBeAs7jPI8vI
y9YOd5eOhtUJTDARZfcbYTFbZCQLdMX+0zltaYCEdNIsUtFjMF4vjYmrAuGqo4UpAXWGjpckRmJw
uHYRuD1Ch8mEpk9iA3/qcaRErOQ4pkmeYMoe9b7JvxrIacpeNtwvz+Iz/BZBBzMd6cL+8nYmYuFm
4xAQcN+cZTrU/twuXDQVdwjsYIbDI9x7XsXCLxmsTuRFk+D1jjFQ5qFHSjdxl/agNVEnuXE9GBlT
CmnO+sACMGy+2J5OEDtfanNxN1Tm5Wx/AuchkSLCHpzfsdTrMWlRmwmr8jM/eZXk2HfwTGhz/zn2
L+gcm2KKToO1JplMBKg0phXTppy5A40E4jiuo4E8sCW1ok+dtNTaHHJ6vheFaSR72obxQqDDTuPe
izwtJUcB2r+2OmaPwIcJCBu5PW+idVns8B+EnBBNmcy1LbWoAJ3lBiZIcLNCUypG8srKkgWWKRTJ
+UV3uTd8H5DMVsEP/t1RPzltIVNz8IuFfsbeFu6q2FI0jxBhENXIrXSg6pPTnzsBdOjwzU7zS9fO
AS+fP0P077fwYTyT4+SqRKnbrOIEddDnq7bkO0+ZUYOE3JR0c9KmA2f5fYCQLpV3OB7DJxx+J2oc
scFIvLQ0XveVmNvVF2NpsV90QZMtR/YXhZTZkM4uWv+wMSCliUd8ztjfre3B97/tumfGVNA6KZvL
E/KNV7HUCxynI+j65PPBjLUyAxi2jO/EyThqhKM5tUSaQTnAaaQEJvjudxUXhwVYukezYXdaqG9a
hzrR8pnZ/+IO6oma5OU8m3RfsZux62voTiXc+d+Q7dmNxmdhmNZXllng3i/pKdc4rsOVlhg7yF4k
4iro03hciKXVdlnFs7pCmfjL1dLiW8u8e8AmBrIbGgbHnj0zVy7bfWapb8Pqy8SUg3FMGxUGkc0p
JV/FvWrm4MYvtfERfGVWXhLzlE4+owN+LMFvhFX7lOGEVJobr5WhiBdeFI4Rq3kgd43FZDBViu+3
tUnz1/JvY4H0k8G0N9h3l1ppO6PwUEpldNWdEcaEs+qJC7ni2Zk0m9QJM7BI8cwYQcsz5hNJJJKC
QddjNMvh0SD/kZmjS8ALBURdYQyN80Dg+tqi32g1s9/NuOmqRZBbE7DHEACqN+jLiw0LH2pdaSkA
WLgtQoAWsIw8wNVelW70q75L5uO8aIkl8n/VnHRTXQBWpn0qYmUUp1Lpr2hb5nGiDfy/cPPVTaoM
F/l6l9MB0rjFa9VUmhQK2e9akmu+nPBpm/N/xW+Kt8iH+CDkNZUCt2+/YV+TMc6Floanm/N5UZIF
KXsncirnV/p5gQbFR8JgFtb0K+kMBT7OETOvZixhGl54DVZbpW4z6ZSZV0vaB0O7h3ajTHrtkNZ/
ws5rcm+7lARHzkYtsmhD3QZPhOYgiXi2Q3t+Kb5kn19aSAGovtyU4o0vSL7ypSXiOJU2yq2y/ZfP
X0VYjdnvb1KmFYRclNcOmfwWGkCEOqywF+kSQbZyAbugCxoxZIudva7daP25SOGF1X8rLab6QBqd
xM88h/siiB6m3JIZc4RcWlUWq/SH5bjliyVaqEjXmwy6Ow/Bi3QgFA97FIL3FSVYzzY2KoJAxZNi
ndHcptGcd9PIcEsJBjU4Qj9cTQya6o3EfvPP0EkHQmaKoid+yMtTNlUurepm9h/m6ae21Fu8Pg7o
qE9MdhKl1NDc/LFuTfzYrCuwMdkXq0yF6mAsMN6I7tBNGIB9yE6ayZxPQPjuCChgb8SuhMaWmh1z
9nShf50bRp8a2bw5P5+fjtdZZJFHfmU/SnRICQ0B7OH2hMKohKpk6JWujmFAbdmMe1yzk0N45Dq3
sCBL/1Ba+GicxpMzwHItRR5IN8TeURsu74GL8I8SBe8PHSAXCCDAutMbmtiI9Fus1nSgtCFf1xFu
YtEzCEqrAVGn8s6/wS1H7UHzjg+DHPOK63db29Y8s/8Ea0j2+XIjHaZvOuYjmd1Tuw9ed/9ZUAuK
SGkbpOxuYgRDh7QFGQYdjEyCoT4arNVLtxKnapxvfuAoh2NX+8k9y58jXBmOpGeZ1dHr1bKoV1BJ
I0m9NNGnsEbfkwgQ751E3hvSkmMYCmF4PWaVhk56M93zDJ7jnCzMMUMTNLR3C71Z1MRGRuRAzHqZ
xpluw5avfQ+nmpCOAwgUbph8O8JpYLUw208avYU1Q9X7WsIzUOoJoShKbc1Vd5YP93GhkRCgZufj
SAf9Z5GO+t349sImPDDoiz+69vC1rmQaNG6JPCQJkLdv4IxQ2mIicT5upDughO8eyVR+IbqOug1G
zBvIwspyM1ZsEDLFEwODIPvFKmqoZ5j22hRanh0sYfZ0/QtPZsgfIIl2PxL+EkPTy6mL4lY7w2uV
DdVMevbDqimTncDkQAqBhjX5ZjCsC+tenUP3BAi7b0B7MLHpuUSNfxP6HERQ+xLIo44MGrLbI75R
WeW3alWNge2VibaiBVegy9ZbeVIyeZ3KKNdlZR1ZdPQibJHou7zAERNo9j73b09fywHhQ2aag5DX
zJLzL10KI6ZOhiaqdIZQ9rKG/BppbiQQ7GYnRycqK2DWBK9ZiZKcYjNyqVfPRpNV3lJRG/BAJLqd
znFjE5+F4AwHI7aVkm7Lvnb/QdK+01+ZR+6AAysUd8R8wnEGIMBXcpnxFjB2f2bK/9nkOax+bcKR
vHWchMmpd3w5WzDvAoFrKYqDlmBgCz1ZFcrSoKF4+EUB66xj9iWYmGGAf8nfr7iHxe9V+bMs1Jf6
rLbFJWTk87fF7l0wWnUcmO9tNtPQsRFrzAb/ccbSVm0//BDmJen9aC1EdOK51XLUWn+R9aku5co9
K7mRTVEzwtnhBObIquDXgIhK27c69ZdhsniWk8qcbt6wh1AA0I/Z5JQkNNdUna46wG6Pg88LjnSP
grxpaPTErwZmA5gqiFmKDUVbDM8+NdNykH1aMmgzk/WQQ+k6lKw8MpNtHDFnqVU2y5d8Xkhoeu0K
ZNqckzVHmdLfbZMq/2y8HiNYh7tp1uSnQGc17DyY0vVAyOl60UCO+wNJP0EzI0Coliq17TNZJbRk
z9qmLdD6tEoo3dou8eiVQPIFzxn1uG7VXm3YBJgdcT3aTMZr58nFMfYqIwnVySR+IhK+hUY5I9jj
IA1P1JkdYKJoz7woZpm6JjOHlmyrwuILL4tUuW1/4gGCQwNEJFggdpXbngUqiBvrgXf6X1v/j28f
7fGj5OxrbwA6H+gq0d3lwi5zBAS0nyh9ueR8RqKNOfaCPq1kQSx/fBGMX/2FCsRH/42SYu+gP0W0
belyCNtdpemFlBXOjP005zEkUU4DyLiGOhYcHPNe+7wJNBZ5jYzKyg/O6d5lQx/EYxAIOqzR0c8M
OEDkLV4zy2jyXyF5vajR6fZR6fIoM7xm/IPQnY8C0qiBfwQT8vH/4sCkEGg1ievLz5YQsBeDX0hy
RN1dOiNR7jBG8HGIQLmp1GvapVmpdzTtrsE5TAsoulcFYb0TXHgPhJmfasyKzjwkpRF8jgZsTS/F
vYJPKrGebTpL5qxJ7ts5gcb8jLfxrWpuwpEGorJeGJPSK9AGcGGUtik5fBQwnisfGjQ4TVVs1xWf
NzxjsYeizWKib8NN3n/Lc3E+OEqOV6vHb9UZ+x7S80P0AfVo4Hn4SDaVEOlrJfhfCZ8StqDft5FQ
dcOVf4+zAn7d0sVE/Hj/0CsJW+vSnZSJXbmmD0tk1MUNyUFKwz3QPUHt1Tkg874Yllbd06woY7uZ
k/pvVF4Id1S2oDrCvbl/2KbJtvXqhiXbe5n+kq4vTBlQLUTA0uz0yHrWn52M5FoLq1k6DETxkI7v
vaFWR11uB2rvoU/Aturl+Azt0qBqhHxAu6IQE1oeKRCorhwPpQuwvUd/z8rR2pxn2fwm+m4IH3Dq
hEwQoJ22SKs+69hJo9NpjdW5q8VqAvZeYKa7BNLnKB8uHJgK9VQwyb0cp/5mQ5MVUGz6YBGD3yQW
1UevCxM8ZF/Bn8UIJpy3f63lo7S4pKQbmaarEfJtsZlKjHCzugEqB5MFVcOVWbUlJYb/+Xp1VM0J
A4B141mBK0lDgDQMhom8CyEjb625gBhH73+HHN8PQLLV/n1nIt3y7bLp0H5oalArKwJKAY0xNuFP
l8FAa/b20xm1kuet8ZSRn7B5pVUyP2KAVTq0a0iD9iyi3ITq1EFofpnHqUVAc/QLXgOpVNTQaYgB
yXaburHuHb3N9ibCHgRlQQUt47S1OsSiGEoftUxyPRD0ve41sqJDkbRYZglYguKpEBwN56ym3r2f
6TrDmMP+6Zdt5VJCy8uaa3K3UNzI6ZHCb2Uiv/ijCXmjzBLAo78rFnJqzgPgMdyx+puJxLLsDar0
dOUg4EvNmmyIYi5rgHbbji73ocwoacctyGM3yOLC0eT/AStfcC5+N+Q680DQelhUm0PtJkyOM36P
DhOs+Zq5Hiu46KHFKUpBRg6iKeNi83ahYoP0+ELeOfsjfCU4I5Xh92M4Cdp78+xTqfKFgu+XboA5
+ihkbAM6E27BRQ6bQ5vhW8N5+g1FmrzHM0/D82D8RLmeTjlYhQ+Q2eWFsZdIT+HpvvY7aX74op4z
HkDFfoSf7Z9Toviig+meiH8PWynFWT8+BpUCi+hOrTDRvBZJsNtOqaYT3k35Y1GWCTW6fMhGGi0Y
kt0OqQgHJb3ICFIvtNPEllqD6dNYj3UTcihuzQJlGW7rGQOprJvhrXAUoHAnqAgClIf4T3g2sKN9
0+ohpTpxwEhjLIUEw4U4bY35G1spMwhtovKJTnVGkfEHjhhtbb5S+zCKJklpOLVP7ZqWqXIKU80S
wbY059NglneCPdxCcTWpTwtth0t1k5ZG1Z5b/GPbT+6ubhHqGf4Indf580LV8MqHOvf+OkuIgLCF
ZPgq77tHxsItUxYd2LAG9etVPwkKIocA2zo0K6QbMhDJr9T2FI6TtB6c6LLQvAf45+ydMMSpbdoC
Izit9KzZx/7k/YswVxigBepDWwkh2AqJDc5F6zAZI0xsqi87mGCyHxh5gGb3ZUDEF3ZPcD1lKNFe
pA/Eo08DNTm5DQ3e9y03OnDuWtFDfv6bZ1yXcgh7Q3iU8aJRw0q2FU/k2JQElL6EGCOtyF9ZaOrF
vlrEmzZ7zO2M0M+4NZpJTsWbZREHLLiDsvNf4LKGoMokbguP7PPatj3QDI5BeCICVWDhJs0kEcJG
WFxlU2XpKP4LeVXzLw8ng63ycwNP7+lqMutYizWHJJ4goOsNhXPTF471pBEuCIvMjaMzPQQJBAGg
NqioCW3c3+cqz5F3Kr4edYQ2A5pJxxwaoL3RP8erNAdZop93iQgPaCiN1Py+GE+kP5yb/qbq95Fg
L+T2Yx3KD6YtmO8rul4lNardOjVmM/AMP5+a1n5bKPH1h3lViLRlny+LXgAxILWX+xXsIuCNfHJT
ZO+ZWHLA/XYGSNnvdX/VzHYBWCmc1Ae/H/vDXIgeA3ZgWsTiq4SoTkkH3rrZ3NBbrJFhx2caooOQ
QMGG6GeBx+pP2Nqy3rAfF1Eu57pKMYsgC9YUeC12qNQy1In/b462cY6raUE5taBZfmvaXJSSNrPo
63iQblHEAaJFsLRLp7HL9q5Q/50QvBCPMYyuQ5lkO4rPmIDp+oJoLFTBhsmm73dArcpsnF41VCIb
2TSS8+QPOW9PSUN8Rbxc01zgYABSAqsYu741Vv5j+0M7bREaMm/FiYCuklwZxBgDXyMaMRbvOfPD
g0UfTon2Tx54qB8f36IfXtIKFtmb6LK+3a99m8mp6ObHwVw82UhHBf3TiRWbaXQkTr9oLbFXhvXM
URoYrSPu9iSzm6sZz8i4z9fkBW1IC5Xa210daU3xMzdpd5aeZ1HXB/14EZqenXJnxMnYMhAmBhvn
chfnGKbgwv1Ev7wBP6Jn7Nchg6reA65uSldQSR2sgWZjK6iPU7jrUeQe0Wkz5XgloseuPlbwg6u4
aJWy2iXD//i+HlbvEHK8NntvfleTbTUHNcbtz3qcS0l3HAC5pbPBdL07cwkjgBTwoRPJ8wfdOTsU
j2ZXVlmaZESIeydhbT6w69zxvU9DvcFm/8/yHEixIbcsQgU1LI/55QaJmbX5cZ7eG4bYpDlhZoD5
U6I55Wv2YN8zu6K7O+ifw7KkZf9CXlrZ41GPSQNfr99p6H5ZgYtMnBGNQF6Rg7eTLsDn20YeRcuA
z6q7w9aYdpQBTFBO/8FPyfzP7LNxxqgPbU9l4LealQocJa2vFkKjuMifupVEZDZLnyBTQKx+Idto
UPeFeWNFEHDLP4Ltbnb2RmbEgCoIkPZoIC7D60NCrriKZDWgivyBylbCg2Towg4AD+H3+eUZIoW+
SBW0LEjmVGO/jieOUZYahlnJ3bdbuaxRuZkdnfU1ewFEjyoS01dgXZjBgKHFNUaSZKb8ef3Fmz7e
I9OXtUoDcYHtLjlRM+52+U/VCYXEKmWRQATH5mCch4B29zAXYYRD7Pgr/6OhvD2Dl9DssEhNKnMZ
qd3BlxDkEz39WAfbpVFSTYZqcSPARO9N0S+P2bE2EaN10Utu6+RRQXIr1xSXAnEWJMLg0E54o6oJ
ERQSY0VqQICEg3sDtkstYaT+FWeKN73hKwbdRH2RyrDKjaRHeZGVjuk9mvFugQ5+OQ6tdZkShfK3
82AJ8runwjokIDxAO/YR3CaYGC0hdC0vYvf77282dlZ8FUMnE2VXRXoUPaSXPj/ZApA1VRBLmoa3
9bQ8WoxZxZFBhAEFARgjFXPMi451fBLmXJAl5/k6VVk9kuARBTAARm2yIYherbBFUlAfppHRDLoA
X12khMMrBLs2NI5HMygaQVer/Kp6LrpVy57IscAWBYckcaDNO0SPnyH1sp397JyA1n/DYJar/wOS
3kq/vG9c7ZIGuR13a8zpXbVbZlxDnOVnZx0jTnvXuB0fp99/xkMcxGfjS6u41hBI02ojrTjpPpUj
plIvryAWUU58kd6E3lsjC83lbTceqoVvzRaTiWGa0BmpNEtXXDGFxBOsEOsp8T5b5N10Wdms+D7G
+e7kIQTwFFErfIc0KcEi13F1z7jMSiOEQ9by2mT/e2OhEt3NZ72P3WWXuCL/ZP46UTeLNrbX5fZW
Cr4u7oDGNb3B0opmxvnPoBSIVQ4kYf40x7u4cgP51lPB4XQwSwSOdEE57EbpbWJuF4if5yK97Dj+
UkEJhlvVxU2afaREttpiZFLQzv6A+DPBdfZFYtIAJKPXPVgyles3qqohCziag9zyvkOaLMthC0Oy
GPhMGwgNQlWtvVjpTnQtWgsznyPiMCrSktYGWd8hedRLqTF97tTRJyXR2U/43ceMW5OLVNV563P2
3mYTYmAfgh+552UdMe3riUzvFuzTKy0o6iC1U05jzEHNMyw2Pt5Uaup2cNlUf+QKWXi92Arn/VnJ
g6ZHQPoPBQ3ttSKLywFaFow4P+yWMMxQlS5t6aLGqm4BiW/7zlProSZeAw4gvShvO2mf/jnN6Yxf
vdSSZhdVAUvxmCVGcva7RKBmehaB1MLj2K12y4z4/v9hC2QMRCTvmlE63/U1d5UkHQZmMwQhaa44
77aGtBl9T6vXbEnUWCcRU6aGVSJ0hO7W38PB0Bimm6gdhUXyJywjhJ3uEKjEjazOeN3ED05N/xUL
82+jSnONtu4QIklxkM2OLLpG+VHUf/QZDas8Pd6Nxk8wZDrULAaz6baLviYtCMyyX2UIitZtB2zb
YG2ayAPXGry3q7ILUGVvKfdt0JNDlSE2WyNVzm0NbxaN64Pwo/th/qNLDaQXtKbCeZ0D7TkSLr+4
z7ufp0WzDHVBjokfrKn1hVJQ2CmWwasm3a+JCJekULahCBEN78eeWzbz9WHcGE9qkwEmAfhCa0iA
I1U5Qr8AVrcPYnXJCGzvC0ZKjOF8KAFf2KBld0AFYKwdwUdj1VGj9KiZaeCsPGVr1gbCfqAVeLH9
2RjAz1tc14uUo6CJzSsDWcHlF1dN17gpa7KorGHE9akdaqz/6Lu2wMFFn+qOdIC/QJ/Zlb5r8Zyh
RVj+Alt0/dvkz4TpmEv6ZmrxUIr7tA+Gmt+eIj1H3GLd3zIN5Ec/IWfEIJb+9JhIZMlAO4d6N1pe
p9ES2TGQu6VAzRK6pDXn9Q8iB2wgpBbG6RXpXvyCip1F/JZ4Sre/CUQQ754i/wgw3lwIKzCGYXuI
llCctE7fGpUSl6HYm02FL1GwZe79V1u5QetIlj7UJ1cLXZZWm/gMSzbNQWWqzFUUUW8RJTi7qcaA
Q0hUDmcpmrzJYcHcS2xO4xv4NwUS6RHbgWoPGgp15LGYPR29s0BENzGsSLf/WoGnZhtzhmd3DrS0
n+xZNoVi+gDwJ/HZTLMpoT6TJudCy8Md/XS9MzQIBpESNTNADeoLw+kf2RzC1U6eegeaDrbNxWqJ
pNsX5g8oqoeOyzbiJ9Hh97d0MsJr1lHTYpbva6Hcg7VMgGLTaidZdgXOS4JXyB6fkosk288ZAOzy
J1HiaeNcjsdynWcegTq2zMDZ0XWftRpuTdlGasWt18t3NZr/p4OGAY1LwbbmHo9/oq4d97k26u8W
2OeAM28IyyZ9i8MEtR+NeNm3htk+c3auVCA2Gl9Em2WA+Nzb7e1c1rhkHujuRrEpwuBJ9Zx9CUyh
dz7rfWvUNVKvOvbKWdJiuwaUooWqYJy8/pngcnsm6SSEal4LIQZqyAQ/iBJYwqvxXZ9l2LjIpneH
3sMSgbEKbF1NgEZEhBS+46HwPbSL36V78QntaJQuhuO8jP211l8k5JEkoOchAvOlqzTVauKWgoP/
FY0eeYP9w9/mL151TfLDderxf+q1Z0jvF0hY4l6E04VdyFyVmeaLaLxUOwoYWS3k+mBurEZ5/l1L
0yL2uUsOLbntID+xxI0HvSqr671KPvBEtqzUBLZy1lHRajvlCSZwdDpXw8TAgjlddgpv6Qvl+Bi1
uOtQMGoKfsOGh22odmOQbjl4rhOS1eespWvsucTddv3e3fFV4F6HgpQ+JBTctEPlpFmTetmPv1J2
+gRR8vlQhuRKRphtnyAF3UHI0Yw/t3pyh0EICg8NomtSFpW3/916Fs4DxF7ad+BqCgRl9F4G/upI
YiTy1q5iqbu7tukxUKDWXxjYZsH7S/JWBgbmo3ag27Q/XBZY4eYZVhu4+hE+3TCdVsYHh1ewwxfJ
42QAJLJ+amTY5m7dEGAaKL9G0bnAcBYJDQMnN3MUVm1Q3PYO6yzKawgQ/gkyGk4mtOAozKd0RJrh
JCbQlc1YAAADkOJrms98byDWDtPwqDKIVW6rSQOTzt1WwFy7NvgmLZ48JOJ/ILL/Az8UoxXulYmi
9W3TJ6iLlPLJemH0qjTQSCnRonVZ1APHckDuBhuluNSdMS63cXUzyoRJ7lc6KGJr4SOZ0gcDXTVz
aG5n0OT/3o8oWqk2DGnIwGpOOquK0Unls8A+uBbX+Uwm4Tz0BO/NYf8IovRwb6IKfty4tQm6749F
+aKEpO3vqs+t9McjfzXdo2ZWcmo4VxJpzMMCWydRKUoBlFUE1uRVHvA+KUXxoVPp9hBfOUqNTClB
kR7j+i2BBY8dcx1lt1tAavZu1lRv30/awqr0WzqT8BJAf+im9vcgkj5dXObHsOHkATXb06xlwrKa
nWCGY8jAiZOFH/KfYQfBLcNpR076Jmmv215mAYWwT3GM0c4IuUGv9xycVD3CZ2KXsN/CVZ5Ai4X7
0UldEOX7sKM7yy2k3WoOGk+7daoQuO8TzdRm7oTwp+InmNKGxt9CEOO0V3XGawah20rPm9PAtAov
PPj7lzMZ3P1Qt7idSpkRkiV4nCcGhfFEtCD17Xt9d51rgMTVfVc7j0x+C/ejtDr/y24s8VBTEogz
IPvynfmVE/Hn/s4bJTFg5oze8V3iO+LLmxWHEbNveSI5LDxwFt27vfjisPzSOme3XYiumOWjPJj1
+6aD3v5B+8kN2cKS2JR1KBAHLBvWkir56OqVvL+j6ZlMmL5pqVtzOrof+emMtGYAnWQ+cKMD+e+J
lQw+3JzII0uc70ob2l+GVxfAwkmYtffONx1IcIppUPYdPb6xa5impL0gaolTCK6IYHQZzv3M8Jhd
z1J6gKZLOkwwLuOAysdUrGdruhR6f1OHEcVnbz9nsHsnG9429rYUCc1qxdMlhgcTKM81paAb52UT
LjztU+ewT7Ez4F3KObzqyMJgRfJiBp2/XkskokwbVQYT3ymqYHMECvtxtnghPddzF1MbFXNGxu/y
LKtKjNle7ywAZGAT1k/WU+jqAkDcyttK3zGZmXmjJhAjHh2hi8fAFHnnB5ZugSeCWOpmEE5L4IzM
t+Cv9dsL0VXWoJDFUT7z+Al518k0llGHDzkEmTX29xbEjPwXrszvq7UArdtsznfmRxXVAYQQGwnt
mL7ioWF+t7hdu6aT+BNR85BBBpUfCljvCo2fdrBq9wADplM2i7kldKMYWFUNPaIM+5/3erTw63U0
NDi5WYw6VG07ocpWZ/e8ug3AOE/tPFw7FLCo6xWh3ZJAaK/vjrq4GT3Mn9Ll/TTezAFMIJ/NQoDf
0/A9GF9vBKdKMKVNxYAhmRKtMm2Kb1dvktVOOcRN1t4bBgJis0/8zDbPX6K35Ij2leVQd35kC7g6
26mXp5w+WtvS8Vx4T2PhXVJYgYUnevvUPkXk0owl3eJ2Enlaw4o+NeahG3RyWjIiuvafl3AnV4Ie
iJK2LyI0JexXB+JCsg==
`protect end_protected

