

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
bq9Fhk0/GLv62Kdp4GNmJBK3rV/b9RTXbbI2h5PtAqSrglrGK5Ok7HwR6EEeSBE8/Z0c0P+WbAFD
zyx0FKROuw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
WpZf+3eiLdpJYbqiIrakT29RZMomGGTcm6ljLiJjEZQDt2IELIyxS/r1BbFUtcgZxmLJxhb3YxI1
ZLQgzUSVH6XgupNWv1GXXxdLr0EH6vhei903utbVt3vE+VmP2fhcGsCOfq7QGSMKGQCbkUjuoTHk
bXwjRk0AR73DkUzgVfg=


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
g2wu9JZ45c6wElXuA1w3VVJRgE7B9dKqOKpad2hq1GxrRtt3DTdcBe3Ja95VDOehTyoDY2JScfeu
BNaERj4rPSpz9eTqvn6ni1KnVzm/5chkJIYoybqMuWD9eHlpi/zQgnmEvVxOrgtJdsQMCE3wyovm
0IuHig4w6aydst4EHxU=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pbjreFmgi/ecPbQe97YwJwHbQ8xErONB3Xw6d/ORb3Q988wgyHCGXou1S+3+vh4Kh1db0kJTEYjB
E5fSNU9tzR1hDPSMJIstpHpTcHO9iXQw365z6oTbmjybdRQMuAr5MihCb4h/KE+rwVzTl8H2WWrd
pchw960F+s92KoiyyKuWUCdi9kd/bF1/5AgMHBFmmvBFps+aNCe9LPZdRGrytTha76gKSEekPpxS
Gz5GRAHIZ50JXkYEpXHxydTz1dTOD3s4qJtrA/5dGreREmtZTngylAj970vudfKhFqPPCjwtcHjm
DLlTipNo9XUMZ7NgeogyQpq2dLX3d/n/5Fo6CQ==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Txl0MWffZrHu0+NsbiOnDFRivawQWjfEPbRTTGQ9uMjcR6If8fL6GvQnz5IAmuNhxhUrNILDKLz3
rBzxPd/PWPJnhGC8/slYUx1wuWNmRF9kK3IEDbU9ptyhPEdUaTI/16ooL9z+ks/bCkgiet3tvCmT
CcSMg+tZGwpWnV2WBteWnPAy3WQTgJjBwAiRWp1JgBCeuze5NtthzTtsilGfdFX5f3xw3Ub8woAk
lsLOCTYPKVbgv+XU9+U/xCPXEE5ZW9ttEy4HkBID5ad635hs77rQVqL6oWJDsLP8RPrpAUS0Zvrm
7brOm77sBE+J4yPgHG0APhrC2Dek348JN12o1w==


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
nNSZ1VwZJdDnj30H3FwwsIQGHOhw9ZnJ+mY/NxGpUOs6Q0mrbaggv+/DD0EbBeGcjM7xGuk7YzRL
WrbwM8iAAhuPwl/ILc9Q2hToNA+s2uK8WQQWWIGPaqLTz+HK2991cPdqD+G4CFauZKZrSuPRlMwO
Vtgsabf7HupMXUf+gqkwQxJP/Z5m0ZuY6KWiMtgYtPhmDusRrl6H8Pcg8awglYP4Rqr+qqp5nw4F
GSQqHtfo9ryxAaJsp70Y2/iK/iuqd4agSUt6/XgDmbQshUSvNTFr9ZX4tPkrXy/noz3sGfl49/KS
MsZ27lS6owSlYD51HcoeSVd1lscGtIs4aZat+g==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 551328)
`protect data_block
dKl4Imr1OZc/qgqVFq63ijwjLBh3pzCpLJWkTtfoHn5pH8vQ/WSEoagBUIphUUNGDJx5vkWN9lTk
VPaQtd2M8ZTozmowG4AhYaPuFSrVZ6D/jfXqJjb0uSHnUyow72Iul0t3oExlTzIV6urquEYqSLiQ
/oGOu+c7pbu3cuzlxtzxidIgjfIPZC6htinEZgqc/Yj9CXBGpKcozbgXwohIAaVObS0uppvn31Y7
rLc9cEKASvUTYgtT62PBLhGXRKFGkYKWs0sLef8xooWuWIsldu1BzEANVzKWPM0ulF3E+CfoMXbE
eX+KZlfTJDm6qspq7umeUXUOe4IS8pcQa5ACfnad5GxYgirK15or13ivadRAYBzQp4cpTcWYqSQU
zovvQKSkOaCpmPRZpwlTSzmWcG4yW/oBU8RmJoOGSnkR92eH01qB4R/8hBRDy1ATuR3IkrAiGBZV
BET1bfaEfujpjNw1INi5zuSXwg0XnEdAjRs+Cl+Pi85AKn9dVB19jRUU5vs68BGr6p96aDewzhHH
03FcgZnhs9OVm6s0pclmb4couhTU01lXscQvUzkI7OW9hgHuuYaAG6QJ0X4f9J9SXUe/YRlSSETo
b/OYki7GxXextnAzSV0gj4WO9+UOimY++DEKNtc9VLhpDKzMfaNL35Bahk+Q0ufXbvT5OPrhBChT
5pBQdTXex1PoshJII9TUm0UreCbYfXfsAI0yWeMMhhFgssoQAaIRhQZ+uxAaJkZHWWD39oPiCvTg
FSiQMGK9tMQzniqpfaUxKlGwiIizGU8KAqi99WczKoLN3IO0VENo2oTNHjTmC6U3vs7a2225qyU0
E87C97cMKMa4l00FJLjZPG/LbMMgjaAnqT3Z1HUEUutkmpNtlL/aA1kgGlm0hiZc6KsAKpJ2xrPe
7an6YrmJuVtQssHrFAvKsGKubb84UDzLg4wYLGAMaGLpsaDH5RXPYmeK3jd4gtdpY64q1X6pD/Mj
itrIvrYr/zKtNoY3nzOd6n6B3ydoE2ln7Rhx44Dc9UlzBgUBz0AUuBEkYUsr8LN43d9BS+X7BRgz
67kXRWoaZtfgwZXMZSlFK2lHLsHSwJIJJqesKGe06CGGrNtgYHVNZY/SgArPnchIX/fJwnN/T/LH
V4KT2vc/+jYXuf7hHvOv1nzZsJmLJamvkX3iMVN1x9LcoziLKuxzqm7GUvWRg+07CsCFKGvxK9rL
bma0TMH5FMDPojp8HUSYU0c1Q3CfKD8nu8oaWA9ah68G43lZFbjaAvikReemKbsRako4sYiKEQrF
S/obPaa1K3tDZxW1Q5SRsAhy6E7DDYYGPGkbkkwerz17yaTPLR0rVWPWIZt4RlR90dn1e8TmyIlJ
oDYWW9tyTbbJnyC4fyOPDi9pfK2D5PGFeLufdyBuUUl+6GwVETtavwfTZ+wMqpNqfuse9oIycRcH
7U+wPGL7XHXqfDh3pLB0gX3lpD2K0Wk6skIE9J6uREyyy8uBK7A/7mb3cRsIuuurojVBNEzCT6T1
8ODoUcw3zhHmvaLaYIv4hUYMgXsKuiNcfOzvFU8LlOFLUX7FTRAR5p3Xme6nOlU2IfvHl70nCdk8
Hd1KAoiNkPvNKsbWFW8EP0YHwrLA2ngriMwNBlm6OPOzJPyxvkZCERm2oWjVs7J1GhqSoyYlsO/x
/x7LqkWZG524iYjfOOi7ZWv9w9DVSPOeI4Q/Rlvn1wE7GjrbooBOIC5EgbppEWHWxyORReizCDo3
8un9CsXQFFSO4dkWqoJoXR31AqSbIeJWVHgsOqlLXITQgZpywcjSfPF1+QjxSeS0mZ/aXdrzlEWf
p2aeeGi60OFubxV2VuIhTIsZmEXT5BOqwdf/fWltf1Udw51mdl2rdGTy2cYRTWWcXboDalqem8L1
HYMe+J4QYMuyfqLBVCmDYWAurNkVc5oPneWuAih5D6/cjg0kLcuDtMIyPt8L18qqFfH0xqMprLzy
mheBTL5JAlVsHtqHbEojL5TD/drEqvCkwiGfK89ZZUGAnxw/GbWMRM7FbPS50RFyOI4u7ac7q6Cn
NJU+bZUpH3adz4kr8pQYIn7kbJ3ivRu1wsung6IJqUSpwM/pKgU+Uz4BPsj+hvmrz/JaDZ+Phknl
H2RC2z/zULxXpMNv1M4eXF4ybTTHr3GSFAzDhoXnygacUm5LrwW6cwCc0G3ehRl2xvQI3+KoL8+6
iY3H3YuSvmJDbGEQAf0+le1s6OTtjTY3bSVki6I+E+nRQglYJ/3wxxwsndGGAPfO0bvWr0hXCmYZ
1zgBj4lNjdbjTi360L2kPu+S8LtrvILqlMTKTKyHLGHibBIb1ulYDPuQRxF88bbC4tmRC4SrNqWJ
aYrwbETTp0uDx1Nz4HWUZcd3b7YobpoiVC4Df8wXTZpWjbIu1rNCWhPXB6FctuAPLwfBtfEd5sVl
TiLzNwqRp6nT3DNWVEBTMg2J6rqtapUOCkOzhlfDb2C9Lzup1l6VHyCjZwZ6NmXeupOFbU9T+xPi
Iihl4uKbWe5vHx4fGrJ3D89ZeMJNxb4Qc8u4Q9cetcr/QKLwRoPY7yc282+VMn5V5iPUJ7mN1Z4S
6Xw82W1N9Yb3aR//HxQvnUW8l8N3wDODJr4lUwjsczSyWuhg1yXyKKd3vzibbPz+UzF8AURsVi5R
Bx3lX1BihEIGuXrTsrikgP3ckSqlZsQ72y0AJq/hAVIMtWz15k5qMyQbdcfFDpdkWTU1hWUiz1Id
orXs1bxtavV2564swXh4TeXObaQralnGL5IvC3sKBYbEWzwpWmG2vp3s/XlkEN0rp14KptT6damn
+yV43snF/nYaWctydM5iqgYoX+LXEGzVdtAR1kDnRcZyGptfvCuRG3g4y6wooOJ29yJfy1+yqoXF
e7CEAZGbsWLpbjXchkCLgKuI6oLh7KtqDrdUpBpZjpnOsVCCNmdal0h2LyQqBOs2sylcDsqM69Vv
sOwIvo+EIwMXWpd4zpfgGcA6vvgJFTq8Blsa71bHeiSwj6qYYRFAA43+MqGGzvhveQMGQ2vwnSdN
1IAsR9LjF34Omsx7GlOuIOmcsIl6usNHqc1ZByVaqNavgw5YQhWN0vFh/kGg4Ob4cg4U4P2JYgVR
atatfhjt7AqEZ4tayybTnGdkeuKtoACqPXatqAZS/T9Nw5HFw2vmeT3pGqTc93bDJmXiwgR3MwRe
SIImA1vUHQO4oYSG0MR+mGqVoiVQKrcyK3KCCCYkSej1Y6lGg6cnWZPQAlh0MZA8i2HrIEFZzA8R
2t7Hf/muMbYqrRw1+g893pAxTAVHIFYZkpKi58X9OIz4iKxl9fmJXiReiBn9tg35s/V37+Ck3pCO
bkGoBILNX+OaO5rZN9/4FLmqF4bxOymi5u8Opx7IwxSl8Cpi6cd+6kllRVaI5oDxLMqE8CvBRNiI
2I4YE5+9vXm+32uF0ikG4AOitSIi7iHog+bGPI6glyQHlXn69muwdPNF25wshGvrI70im9LGdHCX
TWY/ddylZYwVVUpmmBtDqpnt0o7/f9vXJD9es+wVD8mM9qK7T6iszSW5PtHKMmkpVBF7Ncnayf9R
3188Fu32XD1RHXO+rNODTwmtrAML+dZ862G3sIMhbsAlJUaiKdCMMUNxQ/youSZyOzL9yLq4wxtd
IOor0erP1Qfw6H0uTkOfuhZ7qvtedgoi5xUZgMSAefi2SO+dkHx8U1RhxvigPLjjxXG9ZuuN86aB
wUyJuY9dMKya1tBDPAy7S478/CBi8Z4fdlqyMbzu0APeXmgDbd4KygR+Dnq0uZSpuhhkiCqtxEQS
/uGYerz3TbBU32hqHdrbFV9hPOClAt2kwXpKvNh3JXvHHr7Bip52UYzuHlWS+b2AYfZTvFsDJShj
TC/HJgS/Yl7kI/j3W+z7b3M8I4pg6RR3/ZinqpNoetFlc0mQ5A4QezDBLJ4hU+nczrkUs//RIflN
dbeybleZwB8MT3Opyeb2GFWT5P2FmYZqTxRxqXp9o6sPmXo8kE4b6LxVCswyyNXL2D2hxY90FADY
oEya7Vxp1Rvtjc4oCu110WLyIB1iOPvmg9npPfQ0hOAGl/uvY6YE+vO2K1WNG+g3AphPu3CGT9zb
EmlVWtBQgjlmchB7d7ZMJ6h+DOLH8cJoahneuQcA4P8MM6q7E7t3f/9bSD1lkTRkxpkmBlvVkO7a
k+4PHjuj3FLpFG0rJRQtp7cwYRoKDnK1h1XMASq9g0GXzzipn5oZvxAinpGBdPtniiCF8J83pDOn
69V86GjlNBm6Dz6Mepoufxw5jYCt22iW0egQqtyVZ1lbiYhGyucMsYuiRM5lQugCepbONu5vaeBO
lVF8XBZd/Y8OQAKJl/rj0fJuuNw4weTmS0U3dh+nFXmKavzsQUltlXvuW6TSpVg8faqCUaqC9y92
IUG+sBy7MYrsDstbx0P4wWkx4mAcIUq0IWF8VHVO7YIL8+BN8fhTW8RArSqxaQs4a1jZp4BR0rG8
aCN9TtG+NW3VvN11vyibNDKA9x7Ds72Y+eoVWQ2BDPMSfvRVXgGLbYiNYqBvBHjHeamw2gEZ3YCJ
GGerfX9gnKOb7qkoOf2cLcnyJmGmkwB/W0YEJMRwgxqvIyle/qBDrgpchWvgOPM9ASjpjOV7+mWs
gm9c9rsPv0vPx4bkCb6eUBfrSUyAa5SYtxJd9mthVbyc9X+P+dwPjhBa7UA2B/7jUksX3jQgbFKT
TzOuYbL+fGYthDr261gEqjEaWWS27jrWAzzXLwReNmOGpdNji7lwGwkSxHm/RpA7C0vi+aVtUggE
a/MwitpvSm1F+AcKwhKgSlhYs/32v9qS3fOCIKfSYbGAzruMK70pFyuhPmBqr2BTi7Y5HR53+aJj
Z6i0CKhaP3nWYqqN/HhnKbjzxc0Z97u5VsmfVZGjt1MBg64ONLANc7sjH0HLOTtDj8KdKca5VBkx
1w4D0COziK0hRlnNzWa++e9VEEpLGp8ecnG68tLB32sloWjELw3cRbQE2JG6700lfVTrD2nQRX1D
xi30LIvAX58ncc2VKj/s7JJ9gttOUe3oSVbft9owl5b3g7wJOXs+5JvDMaR5A6tKZzmY3b0RXuiP
uZ5NnnHGdLD93FEq3+H/6XZMVFFY7Oy8gub5PNiV7GxZF/FRoFPmNppkOP4rJUVZJAo3wfrZIFMG
4TTP9PHhVZ8L2zB7aslszAX9SXkhyS4foZsKIfKK9hD8H+mrp9awnQ38ZyozoO1h2JwiroLRwTuM
da4RG0Nb+FUszWJXlff70UhJuThp//vH3HbZFfqEb58LqzjREaV249xFVXBXhSEXDnbwJ6vwmjdk
60991lmzO4II7AapH2Bk5Te2Ge8os300ycDB3W0DZYMomcfYNQIOGZWbINU5MwoHLR262IfjeIl/
/4uzf90TjmF8O+eCAMsn/iSj1vDgsbhWnyEt335dJ6GFmlFBsrJ4IBDaO85pbiCtrNRYWc13+IQH
nDLYAvn5iQvVcdr6XQKi3ywEU+v2Kdk8+tDrjnsXZKNzznORd+FHYMDTmTKwf1wi2eIyqLtHXx6I
PQDFJnvHCs/bENx27bMzq5cYwPGcPhKkqxIZP/pcD5We0L6XQt47K2PUcFjw2PMiPTmUG2rVpJ/Z
44gNOrscIyOcgTEudNCJvADhRLu3vviYDMHQNH0alBW1I48uUlIybobiMg7PLOOjEes4eIicKjtj
F7rKycitA1VBNANgziL48nyvgvqXWDhHbDVD/FZC80ojJu6GELyLqkplDAphqOG6kUV8revycEAT
ljBMzquk/74Jvpe6yHYWG1jNaxfpZYmZ6NU5tDLyBpOxmW9Ha10d1ImtUAGkYpvC4lO8zmr2aXY/
onfJFJOrRVKeRXbPU3LDEMa7zpypVKecLD6m3BJ4crQjEVf4GgscDioTT0z2uATnPNKlPUIMZVZ5
DWVyfv4uoGENQGeVuWVuCQA7T67CjiJJf8iaCoGlwFoJnp+MVsMSAruuIaRU+/tw2Fvyv0TqKJgW
PAjWrQ7l+QLfSla+NlpvtYLOpqzaDeh6gCfyz5B5stap+RdjMFGo/Mj+0825nEHv6p0EXvKBFA/N
Mh5dqTEKE3NeBEOegQzG8jxK3VBpDoHO+8JdYAVzsgm1TiTn/Z/l3NeULLl348aTvSZ1rPliYZoa
1MIFTqLMQwk8qH7nwJXIzcznt2Vgz/33cPyBZcP3elqq0Y7eJ1d5cdkrVdCFMHN+9Nk5bB+uGl0u
FJ9pb0CsGNWsS9xEqqe/As/nutIZWdCKXAtC1wvZsjNhIwQ0ZbHY3Izzg7JyIndWd3f1No2OUg+A
i51w560oAbPrsI2ZWvDjW6a4LCYLfKSMxew18NF1dPAN7NdGEmXZ8Nw0rlypW0A6yKVRNbIZ1tnb
7rwno/3nwlQqCQfQ7MEs0OE52NNu/yRLi712CG21XE2YvPQop/umMSPeLPUU7rq7mftkaBjjh5Li
yilzrRcQbSp/ZsWOUvjRBhpkVN0gR14CaPxmUMMCaYbl+hNNcSKgpLriRP4Q5mfqLfFh8MJBZrmB
TaEdqkQr6Oi1Vk7EeULt4ArjrvFbxCF4ibwVWB0Qz0pyhDniyvqwV8iGUAVgBdCuU9FdPkIWGZqW
ocSUQy85CU97ppFRZ7fcRRBss/v5UOOzpeTiYmHHLCigwO/v4p/0Xhn/ZrMygvzB6Z93ekXDDnX6
+VdQfb+MOiNRaYPkLRlDo2u42mXJ6NgdTRgfqMlhF1exHH0vuskeT7ExG0qFYi1neumOmK6PGVmi
SKmY2g2BPanyaHvZUpcHIvBVi0syPSIdCW4ixZud4eF7VTAz4+wgYQL84pkx0cHsShx4oSVCyzbP
eXuoofx/ls/1j8Ab12N8wNB+iNYTH2ZA5/zudWY3KveRRVv9DqB9DndMri+Uod7b3TflX3vgbfU/
eHMsuvK4M9Jrn9r50tkcQGruNtmetIXeR/nt/tXyRacHNybIXQihcsoyST1KtaOvm2/i085l46Hu
tV7h+AwqD44KfcWDXt+A85Tk98LZLU883R1tIWLuNMy3MG/2mHMQK5KPoksv6ipjQsW+mTXQIXEf
uxkrwKdg8cdVTp+ZMxFbbGy/BHrmWB/UvjdtY2yZuWwXA0L5qWjcXB3SJ62hDxXyNb7ywQnt/klt
WTKwf1CtDkNIpwSyt08kyJSgOORyU5Kmo65W+iI56JOWqhS9/XXEUjXlM1jF6Dma/3SWLpaj3bY/
gLYiH5UJlI4Ty74w+2g6cx61iGs+pm3jTgs3U8sp35rEgX3zAKme6AssVI1IAJsDV9/Zr8eJ4jAO
LhNGGRbzjh4SaOAHHU3hwo+kcVzjTgfmxsTsv5j3io++8ohf8XvZWdKMaDo/axfMhHBunwJx9el8
KaXwjUeEd3s/Y6CNPRCsxvMOxadRnnU466qgAWbz6iTaiwsukFzGRDqukXRlCQQltMiP/EK0WlK4
9UGqEx2BA0iUQ3BpF+TfKobwtUCLf7mjnXorRx99llvhF3omn4aBDhwrcgZZCdbVy0NlE/zPo/54
KDoT5id1wCODs692pdieBxTcclo+C6ZW18/8rQ+vxBW3Qf0jPzc7ls34RYdECj9J7ee6qF+/2zMV
gLY5yjgvZJQxEMF+YRBLsYAWnmvaJAEekbSwVL0n9u9rStz46CBerxUuxTNlPeUHjmbcOVdcztpk
W2wYp+ev15lUlqn2QFogVNAVD4eO3kMW8QWwYMs0dZ2Mcb4HY/2eOtqS7ODDHPhGpRpbaRbHv2XX
TIi2wkdsK/k6aemPIAQXS0J0Yh8Xc6PDj35uiVH21gYyJt8JfscXf4YfHxER9AvaCU/7M3oH0+9M
gtkYHQn32zbKYjoj5rb9P+U91k78r/HzS0+J0wp9Y+WeKJzChQJSHG4pqj5kx6fqsf9xZ3pNmkbB
aR7lKsgjtcNw0hJ4vY96ao+zEdcGf4bH9Wx5+b6MlSWIpTNCPMxVv/XgKQxx/dgKMysQIyZRacSV
7jvp93MudSvmRmaBFwq9FIoRBB3l64vJIvk+HiQjt3nMVXHACvApX7jHKNman8l0BnBqAnA7oQZW
zgEUn9O3vm3wsDebmKatXsgUelHrR6mLT0a7vDHIe32iOBhiMQGNPrc70D5KoeyUNu1mAn75RFLE
Ttg060Qv8qsoUa3zVndWlGNj5JEYVm/xpUH0GoAbHIne8EYiy/onEpUgJFRqyPJ7kxym3shX7pUr
RGh3HdzLbuw4O8UqweN4hBSntRYb4c0tJy7PBRqYMBVJM17UzFPDpS70YrFioR/qEGV/2/xRYtWI
8R3E3JSgii5yAB/XHKTR3lLp6KCDfSX+DtHmMRvCK/wAgCse0zfJOIh7SlrETCNQcnUBfhfOl7BM
hT3kSB3F9TW38WaYZWwgADLyw+DmtGAmaLFZ5MYQZGHrjaY0W/49wblZJpwahivl9wgXM/rUn+vZ
oSbQpxDMTrBXAYHR7XR5XiEvapdbjnB+IvLBTNEqTmpz5nVDNDn65BYLQWMv9ZBgPaD5j2kWWAR7
cpu/gD7n+6dYJy/YJsCAOTAt5J+gvJlX8kn3CLdPrkJSQJ7qTJ/fwGLJ4+k5RCF6jnm1uM+98W0k
Ulz5ofksfyYeT+l8GkqP/VPffrlPSZ3JTzRgsQaY/NMlhyIknWCU+KgKEYoMhpUm9AlYUmKGP7JC
lZNnTlHXo2Tg7DAls3DT64zFqSZGE3sws/juNOud90oP7HJjvQaiIyzyO2v/S/7aPOtXDO6h27y/
PtVDv6VteX4xDNVzhsDyT0iWBwvaEuttMWeJqupZ/ujWiLU87ooc4jz3JZ9+pswsdraWslkQMbiW
/KNjhwSNmVQLSUbzVQWoeL1U493Tj6bCvh5mUQkB5Xj0bQ8iibxz8N1CopXD6UhgcDBbBOHgU8ic
eidv1t9ofK++Pmuh5V7KuMi0Y96HJu3YZ1R1deDUpinrp0p/zT8XGw8q84pbXGf7HzLYeAzG2Fk3
QT/bqThSzRmk9YKavW9AVdh8K6dJ/86FRrntXhIFrf/uJI8J4QAHxKrcuibzas89dMgBHSooNndD
o62Qcd9KfQHtWiITs2aaUnZUAp0JSRSNRRCJtrOIURTSlICYmDvJQzfuqWJVL662096G52KhA6sZ
F0iZX3RlDB9RVaQCJ321iSiY14zdKofWDeKF0jRUydAHpaiGOkHn9heTbmjQ0wcf55hp99QqnWQF
ogFLn0xtBbYB24Plu4g0XcIcm7C33eKpzS7oR158OvbsMeCzjQZrc62vRUR+820Og354kF0pBVPN
XRhFhRNJWH040SfnfGGcPVOHXKamvbWaKyCzkO+r3F82y0ZSfKNQVM2T6OQ7CNFzwcvsEbExAMaU
YK/4lvsBf24+Kpb0kgQpWKI0oq6WXpdAKWFc+HBteKwCiMppwQR8Zzt6HBX2mny4cqnqtduPg5Fu
klwaPtOaH4Tcg8zOxHKH1apiYh8bCMOSq1x7wiTLnRdqbF5P4DSDbb+jnu1ZeEHoi2l8Ev40UnT5
6JKc0ZIXM9RZbxq57We+sSSLd7HsalPxcnVCrvBeWdHP/UdFLSpGbLJ+qC9eqG7fHRBf8VAzy8I/
kOHRV0LNRdlyCr35KMCCmdi8BZ0YkM65704v1JJCcOx7bOuYVPIu1MQxcWf2qXfrXND2DZrr1bnk
94WdaMmbTpz3dxAAkgcC64OoA2NJL/+DI3JA2eMJfquwXPCRR3RK1QDdPUxBmmXVeP1L8Fb4lux9
vRF406zgw0kmaKCq/ragoR53PJzAjucfC2I8uKuAv4DN07wO1t2zZjxBpbdsmCNE7pqk7TLX/uQw
FtIoON7420gLpUhAmCBs+c6FcgowtnOQ5FftTa4Mo7rR/aWVD6guNGaS8/Tr/LpnpwMypjMcqYqE
37EJ40w3NG7zdh4+F/h6pNv0cKaV6bOzU9/F0rdfMwzrMfKKPWvcaeJGk9xA1BYz1/0WfKyFZyxb
bOWAMRCQs0msrSbXw3f4ckMrKBYYS051pcJrvEeedmMj7U0ju7ahUe/AhYVu2cT0i11J4Z+/rxt7
mzggBzSp1TPSuNo7NPQym72i6/bkIe2BCmhoWpPHI2cxQHTe9QKX1K+9zMTxXzaQRJrvpEyo+qCz
Ds8p5tMpXhKwou3nh5GsMwE054c52THWNqSy6xzkQIPTIq4eLxcYqB3ZCLuXdexZkEvVd/bIf3eH
CB4xMwC5RVbANIdWU04nUtIxs/LZCabJxuefN8yLVwS+bTxFz2yfoLLyOTB5Kwyf5lBfXEWIuQyL
IGygr3xC406Gj7luKxUfkPxk/pjpZYW2sDb6DfEa+gYr1yrPGqKuwVyKN8jHT0hbMTIOY1qrVv9n
VKpPKXdyFm/Ve33EAJxlD8hJ1yOnwORQhMRAoaVdNpfNuCvJXa/QXFwninE/Zt82cOQZpyjgkXVI
IlTyQtQLl+epEANOg+qu0eZmPHWp1oQu28ALOnKYem4f5rFP0Vh025YXUKc9x2gDLof2uA9YYK6Q
Cja69j3jIS4I5LaMVimTqwqG8B4XmF9sP+aBoYTTuKDy+l6ytJuCfib+8DQPWmOxFOCWfTaO3W46
ic5E3/jwsil6MSoTb7uNCEu+PLARr4Zx/ntJyJcgxCKSXxozngM+Ka3pSIapx54VJWvfkTCEOUHa
pcMMb6E63GlBL40syatWI+7vjab4+kgl+ByfBBQFk1N/P2a2h2AF/k/BBkbK/F0KGUnqvvy5Yoxa
VF5Mx/6ws4+NLltcViaNE+jv9tAV3oPtXKhaalh5lEMVqWOHrnOTIwY2GjHXVun5T8peciSvxd84
qHvl6n0W9A5d0Qp1JJdRR33px/9KAJWDcSbdZCd3oqi9tYrZfF+CRU7uVKto//t5x4OHgg3I/0xT
5LttPYwrj19dvh/82lpw+F6W0JnW1ORRR+SwWX5r5FjgqA3m9C+6+WE6wIrH8drJHzZYB2UFr6KA
n5tx2Plm86qVkVgVjZ8zGEnN7UtJMLLxFNy7lmmoTLl9N8pLELD8dlmLW27K2vEAwk+fHI+A5RbW
OSbEojGm05ZrqfoM1jUdaZ1HiWOPOXU9r219nBwU9iKBDXzKn9ZBQQ7LfGp8TthKCCyWezF/M35w
KFtvOkMBqU/iEQnBATLdw9010L+vhG6oYvD4uH5mU5N0GY/ytY3kcZSseVlTy3/5zM9HXjmI49Bo
zChTmwba66P6Wpv/FGCef845VrMIpVRFKh4yLdTY05Spl0OcSpG0JGhUdmOY9gzbEJEHmh5SJuYE
Y06v0BF9Wf7LFiwxqRgKj5anGefPwZfx7mwdqbi28kEYMsS1aUFjMFST4LSCaroPihNj13b2cwDy
ZlhR0emkYMx1b1ZwnCf5VfGG5XYBAJTNMoscWQEgLA1xi5ZndCa3pDmGlq9IqWOCE7ZQyQauV7dL
MCUC/cBOCPGc0ie2AimMfZg5bTEWrNQoKLlZGKJQZWQRmUqac6lygoIKpIDHFlAwPHOx+SridDd9
sMa8Fe74BjCj/uPAfgCS+8cVRDk/5NZyry1iHwMGbH1KaKI2L0P1GnkZC91Pj7sWW0R0T1uWUAqi
1xXrAmrJBhUUx3/eF4vNA0mX3E1M5LW+sa9jgD/YRh9mOS+cwcqITBwWxjD4UV/00FsaGvtd4XEL
VYymqtG4lmrEK28V+NK+k8Bk4dzjrqHoNGxIcHBWSzlGqJsNxTcsaAAp3Xk6knsAYSUe/fqmOFnW
YisxT3jX+I8WKD1DBdmhfr5pUUS5e/TYD25fKoiJUWZCwi+sf2jLy8UnVHCdzBwnkdTgzVTUGbj5
d477wOmVMda2Hz/v14pSuvqIS3KV0E6RkNQO9O2EeA7g2VdLqHH+e6BJxPb7YwUVGl7MAVecUSY3
QCYYVChZ1z6k9inAd6GsAP7odvL5g5XjMD1ONVXCg/dNrNHINFBoEY2pW7lFaUN+6Nb3TlD/o8L9
YyH1ER8VXX1Sqmhd8J+YO5gCbxhbGJGNxANCX03uyY2m+AJlftRPf7uYVGbCWCUSq5N4hl4p6E+8
wyi0R4QX25Xas0IerIBhsNvn7gfnHk4yGf4m5iYFb5pbXdZhVGmrfCOtX1QERWteeeUZXKb4I404
q4lO0Dmi8KXGZxa7+fX6A0HeLNuIrCdVZvkrzGy1bgGDPZggP/mV+R2JktLOE2kP4O2AWb8+G4D+
T/fImM77K4v+VDZ1u/ifNMo2mHK8q4tcKRGEo8qBK5+oEA74BQOjV77Sdpab0GMZUmmE5Vl5WxHP
MT6Xc27fq4mJXItFMXf+Vt1FMxDePCZfwzFvCJnxNYehDNERAMPru2+uE3f/Uj7Y8vBgMkDwuYRE
039e4t6aaSnF5XK29DUy0pkGq5ZfkBRr4xIusgCNXH2pFB8ywolfHyfX2zk7BoZB84/D5C2YXHnA
KYnNX6zHMlnDPNYkhwqoMctUU3+BGXQ4dMNy8skKvdOYe+CoX+Ai84KIVjKhQ+FP24VF84mTnRbX
YLeDhGilkfqNa3Yc5R1BmCUrVUbQhzFHfhn/Sf9j8NT18oH3GWLxTw0JwADh2m+KbSY429gWpIcQ
ZMBdUI2FAtp1PrdzwiSDXDd3DwCxsGtHRA95LLusWTRHaX2YPZZqhku32FrCkh0a0yLYCZKUpkjy
n2r04pF8DDNKJX5zShkbUfurRE4DzEMlL3zZm8ZhtqMgTVnbPkYLO+93vz+bMoG+6aSm2bB9k0KK
WfC3EXMpvjEt5gio9AaKmtUBmHSe659hfd7232ZfywNCv6S3m7QOuzawuRrvMibuqKSy+KdFTazy
F2lIbNYAhF4brg3XmrSjWkow5W1s9E7C6NLU2JysBEDxFechqNcDl3QRFTgokz3anQSy6efxG9sm
9ToZWcnkrK3iuS9eemDgbizFu2MM3c4YxeGZ014oRYIhTPFV12xxGhfqcCnSoOnpYK++iKhFWYDy
Xt+3yaC9IBZcugWkUarU3DcnuSfmJiEic/mosNMHt3ms5VBKdm/QPLmwGfdIlz9wiPCGxSgBalZ9
16tf2ELGRsXFyaoSjw5P63xG2Xs2GkD7iI5FJuUnkuFAVOxmcYede7EphJirPA8uXdqdEGvg1NAe
vjkGDgL8TdgHTwshkuDcsQFswcpJPuiAdmjc8NIym8+M5b2ZnWgj7qOI/BkgcfJcnF8L9V92alJF
6gA4y5Pj/xXbtX6LWjq02mpQgfoAp53GS2lG6YhllwNkDDfAphPI8XCphGyRE2LAT6VJKMjhU6zj
t6lBKktd6kejDBJcD+CPgwxRYmGTzxtMkzlZRgdCbKoEpeBd8KAxpHoghm5FiKeZtra8/C89dhaW
w1yk5LHeih5p7PVH4y/ZuzAV9pDD04xB3wjDTT0+Asei1Iwt5sxbPUMy597paP4BoAOC41IXF4H5
pgRLM3P0tFPLrhW1c7DE2n2mny+fFxs9kR3wIx64RAcSFv1tP/Xy0BTC9UeHCB4lRf0HLbCDg0HF
ed7Z8fvyn8f6czMoErPHHdjW3aGJYWagnIY7Nd4i72Qm0GfDMDRkCjVD9aHFT9fLQSCcxM4xh7op
fH7X6zgy6amRt0/99SQLIdmcM2oaiYwXNw+z5gDgFlltXvb/6JUM/obZnzPt6dHzYCij503eyTFm
lJFMncqiAed+tq9YgRETNNwZ4akNjHy33zay1W1jGQTcn4a6GkbIOWXb+SMDdFA/zsIw/SFcKleD
ql8WTV9cDk/rmqkIFyhSdOQz1EIUUJ8sbJyrwvTqJTd8eM+6R4FL+PySBz92oPtDhxSNPAOUZVnm
475cRBu80vwAKCsESud8AnvDj7rAEP4z5epyzidvSMSInQQpQjQGKb2zZ9APuo60plhcY9m4cHdp
V8oGdeW8hClB0Zap2anjzUjKw4tqEif3igOcGQzI+rd1lAobfiFtdQ4fhgHt30bwHXYkZbWJs1p4
6sJoYqCJ1ti/LE51sALfb0cC5ZH+VtVlx4dcwzDAGsniBuaeB56QgyF9by9+dphDUEMsucmfZKLs
etv2tbVW/0PWabhv0QLq9uTkUe8iNZE1Z+hDy0BiOp0lQDJ6luvCjBTpk31JxXZS7BN6E6qJ4ZH4
TRRuPVe0r+m6wIRjRWwUGxNP6w7Ezt3VmnC1qaMkRJcxqpOhN16U2Ai9d2L5iUbI5rshiWDTvgKZ
76LN+dchnv06YxVI9PGbBR9d+EF0sAKmABEUncpG9rjvMIjxc0OWLeyPpKcgw9FpEmsmTR1VvV7u
Nn6uiTMKvhUM8j+bsSc3X25ZymLKMXfHwXysy0S/I3H1Apxwx3psb0AY9BrXeoHSEJ+q5M1MsRSa
ZvApFtCczv0oLP0n6uLFlUn735/vG0+5thAQ5UUEMUtSZX4jVVD1L4tP3icyrtBeOZShBP6aqB4Y
92/2s6ukOxLiZQA5zXZgjg9kRIoQlJycxBYAZAMBcI+n5Bhm8l6iXW5JUlV6ftk8xkvwbEl3duqM
7G8iuZWWpMghs7BI1s/v0xjM74jDgTxGWn2BQ+O4v4C44r7Gs+7kEP+CiGhiVoiXl1Itvf/A3vxw
c+UF7BJaBrBqJrj6bCrCE5NUUQHbIu0V06UE5jg+HEO1SkMBpviLhPDGL7n87TyY+yTtqQV1WH8g
CUbl4TbikMkp6w3YrJpTImyLqOCwbbli5PbU66glL4MST4fKKjkKNO3To+cDdyPAp64YnVRqjjjG
zvbo+OzFiJ70xukPSW+B/iP02QTBcYzf2fxHsu2iOgVFTzbPvef7q0/7guVtMdGucVaokVbCW+sj
16CI0VizN5pPDOWs+SkrTIurVsunsr2VSyTAsPlE7m7JerEksl+BRx/CgoJbFBlBcmeETZ7nbfCp
jpUlvJw1mLevuI1OAHDApCJZ1a0bIlvxBUu0Oq8lPsGIx2bTgElxqNcIz42Ut+998UieMQp5gTjQ
8iNc/aknb6Eo4NcKh8mAwAc2lTDXFfrUq0OO1FNkxIQouLG1ISRfbSxpjX/IpgQk/mmTj86Bkwmu
t2gkTAV4ORTRHHk5vJmHmjZjdNTDtzMQto/pYuEc2LpkF0H3pcKAp/rR0vSQCwLthOrRvdxI7XpU
f3llzgoKxJniVfhLW7jaTFlLrQ2xuMXkLBfq/kUH5sXurs2hOnxN81Y9JV/MkreqPzNQg0XW5CGP
7DAcQLbv8YVW/JXiNYBs0XzvW/ZgDP6tQT0/s+65uzvPXz4NbXFtPDAlD0jNUXbrwCrRStmaA9gP
aHVxw9cZgjOvezNpN8gfJn7YVGHSQVwnRjP1O3e6Igq/iBFLFCiTAOd0iegRrdHxr1N3tIVXEtQH
vDTIY1w28kU3W/r/iHUMPYVWQDlSRx3WIsLcQ6Ne1fYQx7xjPj28w9RuOEoB2cqnBLMiiiWeuWny
eq5raKroIPJrw6fuI0pfhPS09MpV7a/d5J88lwDhhDbLMiVeUhYm59v4PaZswoq/N2XIM2hgBV6V
S/mpjuiJ4CXxbRz6z3YhYbTOyjbi+r66/bImEd60dNiPGDuDOV5j0nCBOEMjhOTBWWKiO0IVkvJR
LFKv6BwiojbQ/9+G1JM4zyLBh0DrVWA1ZFawLV8dGnD4LLAlJGKkeXVgH4jMH5TapcWWC/E5cObZ
ZL7GCqYJ08trN6k3Y1n6wWwd+1IoE0YMNiqcf7C7roIfoSvJeStln3UHnpGO7nKm8QM9fO7xo2pb
SLxSreMsLb+i8uXhjdBctTx8ukHWVwR2uXL5PvBngcAaVWj8JUNjiUKrakwpkyDDL5aFDs+hy1UU
uKPfPIrXgGtHgEfSGjwr8M7xyJycDVa7DvxDu4oeqV1jDV2P276NkWam2ahqkwCjZcAuEHg93Bq9
HMxJTY/Y2CBvLC+flpXR48X0KRNywdbpDqsChZENEZZMq5cnR2iMzHwuoQFtbXMDfp7riqzxBD/f
6koxVFSpETLxNI4Il2vKRA4LVaSoaRJfQGVFOHyHXYUURXz2V4KfxqIQaRT+iVCgKT64zdyy4t/W
a4s3OT33G5uzYQqxTNmzDO5fWrpQohUUyexnApikoyC70EqYxP0YOj4KHnOz8/lPIJEkWP/17kTv
PU0AUZ4flxicRB6kSaSbzG03rmlb8/yH7zXDyK3aqCtPX3CaqSUdZ8aMUlexwu+OHuni5qxXwnR4
ONgaACiEf9tV/I1f2bS8HLnwyFp55G7yj79qEyEpLrSF9+5v1RmbHAyHIqozeDHgDe3I/BrFS/PH
nnskVqCPSr30sprQGYqEBfKWzX1wiGmPMfXbJ2Rl/Vbcen/yTPwUllAAV4kZTa28y7dmIy+uYZJR
iwRChAy2iFUVNu0g/3Xhg0r1sUpEQvQssBbKUB59H6/9ER9YBS42KiM9+CwDRituemgM4mm9JJPt
ALYET7X4pI3zAQ6rrBOqyGkuWX5+mmrnA+5B649SH3C1s+htFEeRPYGj85VNMYOUcuoyoZs/yN+W
EMrubYGY9qM/T5u8Ey5pA0rTa559qx5fXN87yv9tLaP5zLcKlIy079b+sezctqHy+/mAq2zjhmWk
gO8j4wUEJthf78QTV3VBm3Mgubb0xhSO61944ihDuFs4fB9mKDEdNyAKmCPPJhMico9grwgW4612
lMc+ogZBq7PHqCVJUgovhcWP6SnRAPNqmO1wn/a1XFh2O6kdvERv3HTqFlpev3N6gDgodNay+gnc
zphT/RSTsWx3cv2TvWIPcy3/YJUMYFkAY5Kk8UNDsBKlMPLyOK7JebdJPPTK45ghidjBH66vrq4H
vAbsuQkCRoRsf9vG/MiU+lfOhlBu+kRbrW+TMI1XTl7BhvhPkpz5qgQAvq8+pjGgl9qcKyoiHeQs
jnNZ5fUGdi2M3u0KOq/2v5p0CAW4nQTDOveU2Ron2n12otyiD1jUG6SKllruEqjLyKdkZ0v24ggH
VP9+jVZo0j25jXMRyKrHBhJNweOc1aVtLDdkl6BnsJ2Lf/arw5Idpm2N74BEPfStK78YBXgRjHAy
IRQeSiLAOHkzCWSXB9bGDCxRX4WEK0h+oxKCZlDxaDplCtgooNxTiHDcbbSuC0i/pVqFJdzmkW3R
tBlivyDjQgDl+NnPtudzMp6rKK+o04oCcb/L+4jb/DyPMlgOemMJwaD10f2lBxFTloS7aiQVZ550
pgKgQw4o1BfvYVJgyGqvtw/6MVl27Ijm5LwjeuXffxtG8R+Q8TY0qOB/53bCBCQa/hDe2l7RIICe
PuFUWvxIGq1ZjRrwTXW3aGBv/M4xdCLp4eqAdzCb3ugnH09Pus0KyBTA4oflA28PSvPd0F+IX5Vv
DawmG37zxoVlNdH4Lwx2IaaZ79tC/ngRLo+jJvu/lDuVCEgdcucFCDrUTKQfHg9sxsHsnNHUan+S
RKUXoKd/R+D6V7y267kCooLRtxNpWRIXg8QM3XiouQUaS8ngGwboe5jJBGzwBzQ/Jf2OB6x9yg+D
hnmiEB9nI26OyBc0VjfGjO8yMzsVFzZ5nYUskjMrYL90JTKZEHRJxmE0cFbbqHjUw6F6TdY64sAs
LRHgkqosdhquEWuVFfha5pR+G5Gbuvb+7YsFnVggf2FYUN52QnPGq00lPERWszD3A37khWMhN8g8
uhfFHpm+g8LREt6HbPMmS7uPaptDj6OVDhboPxF3a7KYJNnl3iQuZzIzNkc/v979CEujrk2nsJHu
BPaxKBwhV//4G0pUxmcTnO1U7weHwX65azyEJEhuwsiZp2M/cu+Uqt0MKN4fAbs0CGr6lGbQry9U
b9lHABIHGDphK1cCY8Hq7SUV1l8UQbDk+UUZ52NnYKjFH+4IkDAACpYJJWThaGbWsPIgFDKexvI5
Ef53WepPRgUa+v84mmbdKdLXnDONWAArSuLyEwN3Brlf6WjBLE+OVZaiki52DtMil6bl93sZgaEH
iWziN90ZoLeUHPWvTS1bJ+5B3tn7CLf2iZbkm/tDCoX2n+xhT7VJk7zH84SPU0KZ6IRCyB0KfKyL
u0KI3rCYbeWc6LVfHYddUdIcZUv8oPmDC5arSYTzzH5dLzmAQxajkmiSiaqwXs/3FMpYLdcV3Mwk
QbdTmijes/kT6mi+5+HxnpRy9jVjQ9C6BN0JTYQyh28P+lJJDPJDLwfgtv11tm4gEx4HYjRaRitE
F/IzzYQJ7lgFb+Iqzfu0Ul2WGIhgCM1LekY7NEkOmsp3Z2RV3t13vMGofGTQOGEDO8Dz32nJ1Ei3
YgBeRBIEMQJtvCJsH6VzH8YXzuE8PAqMJOlBjkGR7c8TvWDKohNPuFIp6jvgNFZjOpqIs4iHxtE1
IXDT1sy+XEdj4ieeE1cPXpkf2tNPaDcPMca5kUief8MRSKgtKJ2rKgGwZDVODOhhySOFSgTAETL1
Yci89Cvf/3bjxPHk7Q/R328se89ZQuCsfXhKwLQLSGpoH5cYsNDi1byWhvffOs5wygKEqf3yj/Ch
gNxxNh1KrN/M/tYtZUqv1QIg6tryYGaLu5K9uVIlEGM8kBTRu8NzFt0umlqTwTw9jJ72dl11Kpnh
4SND+R2/LJ6gSCxxwnemdvMW+N9TiwBdr2JShvgo2/yKNMeRgvh3wnxTaK1L37ijmSQe1QQcs4GT
gWJpfzhMa3S1mlrtMK/XgpKfaO59i8hUfC1qPebDP+inkrbdHvF0xEAQX2iUWdhoo/tWA3gaAo4i
heQzZ5vyunbXkrEVfqk+bOIgHqovQf0BLNcHlPfAsfREgimMXx6KKiyzGL4Z0qjfevJGU0L8qIpt
ufGZfJL9bGFGz02yR2YO2hJfZ2OVReneHFtab2QKXk1XH29z4vd7/QxTPovwwLTHycb//9UxNpfk
LGQJd/+VjC2JwP9PCwwytf/MUghqN7ayRCSXI+GCEGhmscmK81GvRKPGEIHEhU9A23wxDGS2NYu0
fUwLJK681XmA4q3bHicPFrTyrPmzJkd/e9zcXwP13E2BuROvfxYgOBlK2jW5BlpzWc0HuuQ2OoWl
F2dBLVUqZwlpPVtOjTQqJk6NGEwDHcG2ba/bS2JtdA7bPhmRFW1rs13kiPpVXKhinolqajaovXZR
4dhMkjAjPJZhUO7vkrTrt/jr3wR3a/dXgN51AYetp3g9yYypK2xDDJce9AmloWUH7kWrKNFgm5Ud
pmpeK6kqmz3dUPDGMIHGsT42nsy/zFYWjYEaH1jUmjCp5r9n18NbovLeQurO1ue4eLGgP3PXTmDp
aMd1CXwQ3F1bYqzcayxTRuvq32y6wmGgq7AbImUjuFxTX/NhFWmFdwAbHT6OADrd40g2XVCpVHg5
IHd/SwVp25OPK/GnOdDbgli6+PNQWi49i3i/hIMLHi5a6O1xE0u3agmOt2tpUq0Vf+uYI4qx3XyR
S/SozsZURXCmiw6e52ytfO269QT+lNbBWdbXqDe/PXa6m1lNi/lqvKAfnR4mXEWS4A1LRRfqPRo7
G9mMbSSeGTPLHLY3CP5ZpAvuHdKj1ZFheRlIZT3Z7aWDCB94DHGoLUogqhPq1YKQ7962dDzhHugG
jpGSZcYYDQucVN8zqemNAASPAdNAzqAwVMX+B0uBgNCFAmQnrn/c6O9USWMIxY97PX8Dpod+GzKj
OKeL02MzCvM7E/8bVcvDXOUHu0CDH/gnnp6rUrUqMp01Oe5KUryr6XDDOcyNiYO2FoUK84PvFTXS
n3dnIILna1wjrYOKX08fA1YJUcGaqSjjH7j958ay9gM97DGSMkkbu/ysp8QPRd9h4cHCho0n/Ita
DnMeF/5BMBzdpON9vC60TYCpWiD1dkk0qyZLltUKk8Ojgv52kiMXvJJRS6IGFJcI1jKBohET+G1h
sXJIoGBUVLj6MhymtUrdRQVp20mNjV9cxNYSdxAfjyfFq+rHpUsMpuJNJYPfeGwULmcNFfKuHViN
/5nEu9JXDlf0gHAAuaf6cTT/DMNqwZbx6sDDKvlLqtThNAZ8CXIBKjpbp4LjPvrYI4BJUbX9/WMd
UZGD7H5BJGSeeulKtBZVof9YvwKaTdpfrvKdXQmlybSxi5e2t9GB+oYySmZItLwd37Gu/QkYPjXb
4FUTpy7mNMznF0Wm3g6vf5n15PC7d8KgACYA6TRIbQ07+YEPgHyldqLjreRLYUogovfdyFzm5T68
lv9Opy5QVaouG+ykumoeHA+2UnjW8Eowks0xuSGYpBeW5aLibhLzCl3c9DbGbusXgHsB895FCnYH
cl/hHPLckIXKwhc81ru7QGC1pIoUWVrjatrGezDKcaSAZWU9FAWRd8Pkua7jNbJe9buWJwJry6lz
JLiMF42p3k53+sfQDKdk760nufxTfuQHwCjccnNYwfTfUVWPhFQm6xBaUcH138EKTfAcI8BSuEAJ
Bqz88pz2mJN8ZbdQ77S0UKpaH7jTp4HfnHHUoO3DTDKWRR/U+Ix3QOwTQ0OyR5dAc19meaE/CA1O
lEXc/ALo641/AGs7ixrKbGOO5x6hEOAXbDoCDPzl7m295I0bttIqWABeBRakpGpxYtCjLaldaVEL
XEVlbgpuMiIO6pi7AEpNDX5FEmzrAcnxt2HhuGzuwsZv2vqpDej2HUA/ECL5vVkFXbH7dsaK6Ker
shuozFo6trAljNBK7k1mdfxmtII0nNviAzkeZruIWRiGmXfb4Ga0zXR0HaSM5kCDvCfMapuSj214
PZUf3zs6nhFp3Lx2SeOnnd1DFA76TlV5MdDugbUF5DB18MLM/EdPprmqJrethOGaF6ePXWsxgvuz
EuaoazW8ef7OB9eZea7aqrZMD84kuMpK1t95psPmwnUhDlhJKrNQpmunlsGjIuvfI2EvVvTAnqE8
qvJ3QCTLRpP6BHU4yTEdUU5u87Qr48bS631zRsZ/+y6bI3Tz0Ayxx4mbax0TSBG/+XacdaotcScu
86TUNHP7slGXurQ1KrIy4YQkEWc9hlcSksi/1MotjBiJ3Vw5h/gH3ESUWwHoAGUcPdKU12xigRfd
TRQUfKaAu4Q8MtWNzfrI8S5Ehk+kBcC021TnmZ2Wiq60gasmPJ9WsN8rZaUnlwXhn3Jd6F7F5e+4
tNaZMgKzHBkFkye6IbDn6xNZbWAQ0MydhtoS4VWp0uQaC4eMVC9xCYJZptNuxInUgkw8ggjBT1EH
WNOKgeW8flHUO2egU9/14tHJ1wPiZj9jU9u/1v0V0LbFkLptXpt9orKOX/RiTEjr3wXf/IHki5CT
JjyEv07uONh10CeimsICZ9lowz1NlPOxMjmR3rVNibgfvHt5qVRC6+El9kuFENylD2QeOCTuclvr
ofQ1IZVx3eLWKGHgwX9I9kxiM8sKvikpf2Pxdh4WuzJE70niqiZZIpDqFvD0jnNxDLWmQJVfOSgF
c269vbWSh9jkz8KGtNi4RGzZ4dsGNC1emkf80Yi2IED+FRkfzipJgdWipjRkTsxlKxYlWQOONYNM
FPGEijYsQvOqD5hqKeopTfWz29t6RDvNh2kiKrAvqLZyIaxE5gLz/Zkq6tSjRb63u7I1x8UZDH+7
K6/JnVGWYsjup+CVPTivOPud7JmGpKGHARApomg1RlKCXgjh9lvO1cdrKcUcOPVJMk5tZ98xhlTj
11aPdcBty+LU+92y/v1TLM5yKfg4LqB2WrK+25Q4eQfDF2bfXb+hJePusY9nC8fUXvROfAObMDGa
8hlIoYq506n2h97nQVrTprKZBOvDcKVbWet5eEb8wc0JOMMOKWtcqXdVx/T7g/IQ2FwW+4J0X3n1
8yh5CvQMR87yD4OqGBoCDW86xtJ9cRfBvPndim/KlIM6IqEoggVwm25x+zD4Kb+hZtJWmsDypE8I
sB5TTiNMP/33zPh759uCwP41048nFdklP7ABujz6hRq81oa/Qt59X5LmxirfVr7bkHm41aUOhRRs
wa6SC544iNvtxfumLZqlT4VH7u3/nR2O0hfPxto6QCIIO38W/TLqT2lZnu9UOwzi+3V2rnb0ld4t
ZLzY1h3i5UagA6qmhCWPR+SiXURcJmfAANVYMnOwdSTf8iqeZjgRdAIREimxCrf0sErQVS4pm53b
/Q0GES+EcRI3YZ9B4XjNUqHzGPYxuNhuS6vRlR/Mq5/3tOP2YuX2T82L9wrNhSWj25I9N5h2ejy/
09Gc8KeYYKmia4bUWui30D6qMNWFKrFqfBNQJZNoxmKhc8tHSYEoOXxq2C4hMQmqAnr88Pp2wq3b
xeXKZaOXlT5ElOu7GspSRjwaysp6zlJezX7mf41c6p1g/wHRYc6vBEix3yTv1z8UP56zoyMXAfo7
1NeoVxSHjvJEiqX3Vil5c7Fz9FokZRNRLa5jNnIbBffyK6QEuYwZGe3no0w0u9zAeXwmrHpMi8E4
Qym9URoBBFznrSF8MibvYkJ25QB9ecaqOJMff4IpMVGyp1t4nb8z1rj0KwSJFBlsrtyu9iG6KD1Y
EN0dzta3L2KyXjM1jSnSAFqhi33HRWTrRZ3E7pSOijtNkJb4X2tKIkU7XQhPJsd5H/FiciIQNe5l
tYW41WV3wXa5XOrIz6mdkyPPcAJFqd0ibyo9f/bNRDwUBkE2UJb0rpri6QKbulvxsBU2dpb62sul
hV0vd3oo1GHhbLz0UonVVq8oVgKMWcaiv+C/DTMlPgMI7xKl/BodWTNpbj8nCUdT6Yyt3oATkJhK
n+MvBlR6CBcL84GwAr+GuLcfkl8fcqcXTLuBWTHt4EVUD4tuO4W/nyQJrifQ7Eiju7y/gzE30/ix
fRd0BqM22+O6U7aK+JjRpT9LSF3pv6zmctFNdkl2Ccbg1e7OQv691c1VVAMVrO6qhPZpuhhyubrQ
WOOID9dJZEtkZYVhMMYciDPEVPl4UkqeHutyW5m7ykHKg1l4Cwgrv+ggc8AAaVasCu5+fKbawZfE
4N5mC4yQZv1tFvFwOfehW6hV92HrmG35G60mtP/pf9PUn4l7Vh6823WjhCVuCdXyyxQlk2duKufe
pk1iO6g38qJ2/7RigqHUp+jxUwf4imDCs7VwAKmb/ecgtc2lCRMPk01B/q1ql/xzzeZOS3UCHtWe
XG3YgQIWGNYPRaJyxvawOHOpGlg63ODzeD2/I7az3uUNbW+1SuDRn38sxw6IaO6//561JsiHWSK1
/DxXuNgpki4onoQJGIILwBKihiayoAUqwaGGDXiRbp2N+uzRpeNLgOI/sthN37dn/PbIIYHsFDO1
OpKRMrS9ScMB0//BQ78nwYxzcoXI4uQyt76EhmzGJHM/iMagHf1k/KOKJW8E3sMZXfn0tItuniGI
gQcOQ56UYqPIq9aYTshSrIB+CedWoGnO+V4MZqqXUMpxwSfwKerlJxKiafqxX49K7x4v0Buqx+7l
SyYxdmlROZXFuyG3We4+YMw6JkUBVGtBWTf9sFYUWEOgtlntZs9pUbTkuHNZ7+NawaKhYgfoRrXr
HLomO9egzNhWARrvnlsYpjJDQsT9N8BXihglNvDXK8uUqrRnEzVhFHUnaeNXrDfJ7REaVbWnrKMP
Df3yI+uE2XhS26tc2QKe+VBmrGgO5jJ03mua3PhRpBOBljML6OXy40Ma/w3ic2yVuRlV0GluulH2
v+dIORO9x3g8j807g/sNXFDZ/7ZY4WCdgq0PKt+s0+CvtxEOHGgJnQgOu0OQO8KKdKD5EF71Qgm0
NoKGXkBHeJH1uMS4aFbLojFVP/wdPdC/7QBg8GkYTCea6CSNC/Y6u7TTdN0j4Miev/xqZDNGX1AI
fxHLejKvAo8zczf+ypqeUY3KBNd8Ub8O5kZ8bY5GrDRxnyT0L5IQdLNv9TU/d3Jk/1yDL//KbK1C
Gj6VPur7APFQVg0kelGW7bcjR8YDsEzJmmUmFSfji9PO5bzgsme2A5fQmVDhRE1iEPhsz2HM8Vhd
AhsnlN7foI/E1ih4f2/oncS6NNny1Eb6MlWrP1ngjZma4dnPY9ARW2VCwSqjQw2JhY6NBB/1h9zJ
I5MmCXgnowvlkM5mFKyxPkzAVzotZKxdUL6xRjjzGWa6xZ2X97Yrm65MnsfLNCyK/xg8xfY1m3Bz
RdY8srnxUXZggtCaqsikbcMQBWUlayuhK4AQd2M8COx/YFIpoFi/tUOE6zJ8cwekWCAer7XfaNpO
7bLX48u8H9b1Y1eYci/sM70yA9XJ7Ob9uqMaUU1LhJBdTx9nyXHBPvh55HVualkFi97ca9tgHYKt
p3CDHFe4pimTEQOeKYI/rzhbmDkg3zac7Ulb/esUJnROTtOZ/o4zldVxpV16AVrwC/podW7LzdJ9
ImDIBaMmUsl+oWnDinN+i/q4C1VrkgrzOS8fR8M8nOHBVPEyQeqxDiA9VZudD8PJvIGWG0X42DRp
m4Xs+AtIuLIDEMmcIx2J8aip5/8om9EaNX+I+FJPeYQgBtuUlxkJDqtp0HVNNu/HaGHZFubpgZYF
OKqkJsxw0c8/hS0F7F8iD3fjm/aK6G29XEEekf5eDnJB/YUHi8RJp/QMnseb79bGIqJBL/btK5Tz
4zciPkmJxbpTF3N7ccsHxoFxpQNOArjTGfwAfxLf/27183gw/cVGUtjnpWDd2yZJX5T/nSPe2vO/
Fz+ksNbtdrgMwdtQ1pX+pUZ8uhttKah5LVcuNUpf7kVEid2d+KAUK3WIghYAp0qHDXWY3rOTSfbX
a1Yd1ZXxnDYFIf8HfAxo5y119dW3yNCIlE8QOtkcTe3xpg2Z2aknpJiIVMeqjHnzdOzj2+VBejp5
qBdD9g8T7Q/6eWwURVvRAUv1ehoz7+W6eu+53lMmZH4NL240+wvuxixIW5kj84Rpy1++9g7ufLaA
dIzC5bsbUH2wsttkGZYWfeucf3u7YEhgDF50F6d7Cf4HyMb0bPA1sbxNn8iO2hz6rt2x/9b6+x6o
aAD1/jP0e6zJXY2QfTLk7STTSVHO69hEFOjSgS2xHb812aV8OriCKoe0L2Rd5IMDme6OrfSTVFiC
Al6jysGnPFEs1EzD3uP2gOyrigkaTcji9AfaDbRQzyGzCAOQMl0gf7OErlRxWBxcZYq9rHpFqI5R
KnUYa/l6Is4Y0BF8KDkJJP2kQiueq3SELLtFDRrlcX6fOTBvosynIG+gH5S1louT0QGN3J/Q7MIH
vUSOXErBeP2p6UzGIi1WRGAnrlsNFLHkeRiqAbO7gcMbalyuFLS2jWeteIcPDy8E5po/NsZknKqq
vsfOM2VwSwU9mFcfD5/RjU2gMwIz8HP4AWYwk2Kol0TI/5NS1lVeZDAJ/YjB3j22gcOfN/sde13I
7gSswFXOqOYSPD4r4YQafzxtG8KEXS2swcETk70RDL7onOWlR+ntKS+iyeYxmXlm1q7KYYiud5C/
/XcGIM6pDwsTjzVMQH8OQAAEEkIojQxsGe/jlNEX0CttpM1MOggbMYfNFoE/7Syt031wA8Aanwo5
YfLUrCm7e9k3zWALIt/bAifBpa5N9fLT4fgcAVH7U0LNgSvkZYD/h/Qxge4WUU29yENGwgiinCbI
bdy7GSKYplJAoHgCSzH7UJWovP4+0KfDTjPgS8xCHTGABbtuP/V46ZNy67aeYpotdLJ1iAMBDK2R
qBFee10EbN+MWfef2KU+Sq4HwtDfbE1LzOhMlF6+QQ6eq0fDSmWSnCS0oTgTNVfrbN9SUAoXlfGK
uo7vca2pI7F9JwTSsk2pinnIzgNaGbrH5ZuFhL7mmc1SZTp6ZeVfaM6eGOwRqNPWraCEiiykzYry
yk9yxeDcKzVhmyeml4/p01B8UCTuKtXDAySoT9MWaB/rSt9koKjC8w7/SbER34C7lOmhM/mTg89t
A/BHIBPyi7CcB6eDuU0RYC98gwrfnoJ/oGSLfvKQT/cEY36HanmZSIw9cdPYNeYAv9pMad6WbPKi
39b9NqcabZgvyWH3Ecn1j3UAc4Nw54SZ5fFDpwk0FTGZp4QgeoaksooV33Wi9PJ9K36+vBllCD9P
KvPZ7Wnb/aDnOEuaZS27DP4Lxb+V1NMQA+AkiWgKFVweLCPGgwfRwCsYa1cgUNC9SygNOJ4fwvE/
jOiDpOfM43ESddEpQatycflpqe3pVx9pwclzRHGvo8YaaaFwO0I2wNzpFyHM7NGNIgtO+bpNt/AI
9S8hnuBdwmd3UGgZVsw4qtDgPIe/7IjF22r7GcUmf+JM89lZ4g9TcqaA/o6VRlns5WtOvjPGAcOu
cwzQGW4+DVqrL0DUO6i8dSjXBKJUP/+cz4xae68pQ+fa98awcJYWRNJHzKXdZkgckOL3IFg0kRyy
tUhtRHaVy3nziAxWUOgdjGoVtt5TLQvzvqRTrMIeQg+sASCyKKoiufjpdm6BKd8eDbvvlLZNEcAf
9iukzKDpgYas+ccpnUvKCcxcA4LaoFO+sDLuGAVfkRpPZ96JixHAkG+pNy8oH007l21+uJFg4wk+
Aye7yNG4HnOftPRZgeyi4f8xC9Q0SjRwbHE36lxLdTpLFff7Iqq+NmrpVAC8Y4pUxiHxEnKBWVQy
eUE3gF3CR3iu2jp2H/GlDhSMzMPox3W/nBtMmJf5fpMrJpCrktY/vCgJYf7BphGhz8PkfzZ/kUas
HvkvPGQlLNaT+OPgIs/QOhwxaHQScT+W3kybvXYISJfW1A47ZYFlmSm2sqLr9bs2OeVVfytSRieH
1DsvWTVwxzNvgHo/YHETmeIoH8uHz0PRvTP3k5vaTAtMAGTF2dF0nswZdb0lu6qlCx9M0QJ/hJtM
cixdMPTbstUe52UPAefw97LAdKXtDV+BEnLtfJCaTgGxFJFoNMxLCk3xxeCaIlYzfOXHikICwSV0
w46dlFjr6KWmmTdQUPmcOJSZKO6WzOoY0WcJKKJjZ0ewTQlejfkGwLM2aL2gbpoSGIiQ0sqJ1sfc
W/M3Ooti/LG9zcFdHxhWbEM9hp1rFcnTuywkb8wiKC3pIzkozDGvkVXUV4QuoakotwDHVcqmGn/O
KRCdFDyjD7wXILoCW6x6PF+MyhY2/RAtH7cOeBn0A/mk+uKHBvu0P6wyAg31F+pugFxbcIlOlrEP
JhmYiqIEYpaD+6CtlA1bKWEdwvszcEDwCYrX038qokwKpj+YawON896KQOxMbXt3yC/hQfHzDJ1J
cHthy7TCHR4AiklQ/Vl6mgmARyODee7/RD9EgxWtCP0FGBFs46X3mGpHbPoCACmvFMH7WXfCUcDL
JkE3fhHJYDWCeTRZ2p7czFIJfwWkxC+1jZhz9KfsH7jc097FzP0MDceY1MdvtUlTIubescTu15KD
BLzkLHHqSqZoEpV/v7qPDK/wLI+2TX2/MEWZwHH33NDpLUNLDh5jsEnHhNHLzrFEp9chMT6GWWio
y1NM79Hv5Gz8GUQlkuZKcRjnKjob6RUvFTxkhA7Ey6gBWpJ8dT4dVZ0Uq98WtTrnjFSpbt0FA3Um
V2jihdrqRbRKZZqhg5gltRhQWL98ZcH/cGOy1+n/lzbRlN5t+/XlUTfYGaSxxrHsHQAsrZRoVVbZ
4AOiFK889Q2wf/dNiJqMd1hNViE+JSsie25op5v/Yrm/aWaWa/fchZ+eDposwvuTeMCntjcNmlaT
8tkPBQaxC4CKKwV0JQzAX7ano8pjSLQJd/D5Jf7tg9mCI+U+YDgaQDZmBu1/SuaokwNffV7wFfUo
9yiwryOY31ZT2O/fcTHimeg31jhD8RQDD18xCVpnubLy7UPm8BURJ/e5AcCkiFXXy/DJ+p8aSQc2
Tth0NKpiDHieCuc29X5j3OcaYgJWz7QD40Of9iEZvXwVsIhQwPietFs7VyBq4KfFgUCO7FPz3t//
zUSWMv2dC3e+PyGJFTT4sj0n6KObMzftI9tdJX0BxJSw4TxL2/Yz1M/IWOE8ucD830roXFocBOLP
Oq3Lkz+hjJvUQ8eB3CYwCH/N94cDLABjwDSKh2ObXav8rL9gl/grBUnGnhBpEO3Vfm0bHTN4JmWL
WSeUGTsdqfR2nfPXZWqFeg+zxv4taTDXaE95/uCf3zN2b3J5G0LjpuDIw84rvLoki33QSfPYE+MW
lGw5ivJi36fTMKrLGKqeS2oII7wJM36MJsIKbE36Gm1fELdGkAYkhGfDh2271nsCK/p94cW+/GzR
kw6rkQarI7q4XwpFDKvNlZOWRsurg6K/bahIK9aTO1Gox1DsrHnA7YRiffTZ8WMZZfsrkhyYozmR
xSLJ4xk1IX67oDH+Kod2Pzlqi+s9rCrgK/5dE0yMNUAnyBqbrshR04G1UWQiqDZDdbijNPbzUsbh
58Hyff2KDRlHOaVID/mrYMnjiCwu2PRRZo25htJrcSlKTPN6TPQj+DNzlvuZFWbTYeb6jR7SNw1h
BZheK5G14BkNMrQL7TkdkESuPnfo9EW11AEfWcFzQzxgBGpBPldsTAJ0IQ7PrG1qq+F2UBHISOBz
Ef1Z+8awcbRdEOCINqfMda3bw59UiUWOQL7woJYeAMYqeAw9CWKMZ9W/kmbNn8RAkryJVDU6QI1m
4Q3vY1vyFt+OFP9/vYtBS5mfUWI1QKJddqN6zLRx8M3/rZbGfQWCbTcc/aii+LkPrcGNef4mGgKj
DN92OTiWl6dHeMOKecQRHtvYPMMxNB3HfrD0f1P0AlHH7YEunHPu1nYvHb/gQH3F8q+y4PHLQjSS
c/tR5EEM1SDoGIqZjJx/OD1K/F40EfqWccU/YK1TrFuClsJJdXRB/63Xgp5B65UppvWqnN6rQy61
LmIXjhFRxfV8CNJTCevoL8t6X4GpqI+59BCOOIIWQG9pR4QACwTiT/cvx5QkfZvUsIQmF2MRqg/Z
vMK4jlrxf1Z/nfNabPD0lsYH6/+9s/CxCXUv88t6bdXPu1wZlhaCdTYxcq82hVRad3Ip+hC+9sJT
7QrDhhNDHjXYXFV1Vyt9+IH0TBMUyP54Jjl55/B7VrRgBN+DSa2if2ytvVBTeEEZqUcRz2Sx93xe
Lj+uWuQLqMKmcg64l3SH5fmyjc5XZlfHBxAd7G2LcHSlMUgv09QWFuY5/WIICXu7N6OSqX5DOh0X
Ln7XTevHkKEgaTkq1dsrkiJBK+D8MO8BCvl01wT9Wpzc5OAfqWjJxk7eIdIlPpQ7aO1ZPGUXN9st
2DlPWbsRs6gfTREvcmD1t02tKBm8eOzsAm+7MOMYC8xElsEK2v6mSfcF2M3bK+UraZr/iD6zjXrj
7ExDGltGsPO01AftVbj1B2L0vSfPCsy/SMxVFfX6auwx+8rEqTDiTOLvNxFKrwAeoPoQqf9V6FBe
sBUHH0s8Lnbafeqoyhiu/qiYTU5dZ+heWlqcaTIxkYtEhU4YCK36drhisZkQsJQfPPeCno+cQG6X
3GvHFd/95CCzyJlt/6vely7BHzjK50atf0OgM/NLT9SgsbUXjpKFyjnDVsuV92hJzLoV5Vy/5Sen
FBYa4Bc099YTQhMjB3SMXxF/7p5yEJWDF7ljpHHdBmIu034H8f4V0+Pk2nVJRUJkdoiUkCq4wSE3
vzrCEoykH9dP0LeCb9RyQ476dusdQvx0ryLtThA5/ohbAM+2f+pg01JF1wtcLzLtQ6klhOSrgcX8
1cAhCOUY6znp8DJbxfwRFdCeufoesYmHe31DULIMHnOJ3lS4jjMxe7jUmuuqL2V8dZg1botOp3wR
3n23XfAnj+sxsD5lSeVth6TwbZ6xhtJRnOx/E440wFo8Wjw0MljacnLOV9dFCBObpGbgbtiopVCZ
9gQjHMzGSynkeBWJruEEN0kmhXX42F4s+98MtjgxuWM2amQfbh9O+nF7X+Hxr2un4ca0SJQgzIns
e3awHhe/AxdBPNEeQV56M3fO51sCyU8GysTdVcq1UKJtq6wqpnWHBZa12cw3IS4Qb45D7+hShMpm
Kz53n256ynWWbVUa5sR5rdahDgLOol+5mZIeEj3DaMnJ++GA+APUnG/wf02JIqhjeze2PJwqS3sa
gOtLDFjVepnSvKFj0Y+y7aJQ9SNykc7DzZ3rNAbwcIEGzjapePVDplrXvT6LomFIxyQ+kAC95icE
W8QvXu2Fdm1UqKg8BTgFA+mGL+UoUTkSDJcTpfW4aC25qsNfRSVeVkMu+pJyQ/pJF7pJJAIaHRUM
rKGF23UVDXSvfAsSE4Kmu7+fXgKhhazNHHijHXcMlUryGYZUlxUeJsvkj4+Lks74VSsPj5/pLNbF
3JOZYbHOxjG+8FWYP9cfAxZd9cLMlTwRT38Q0u8TJ1qeo38c22BWWCunuQcsmfV4DOmEy43nPLZM
w6v4lo64ORdGC8KAK/lcx/JP7q5vvdXmwvPs+Na0XOVetrwYYs8E68jBbuOF3dL05Ij69W1TiHRG
4ERlQEFrv2vDBRIPguABIhmHpXEDOEknB/XghHNntaqmYVHMI4fBYJ5kQY/Nc8NsHF1hSVr3b1qo
/Qzjs8RLAcP/EsremjQ3412/htdkuL7oHeI37nAYFavKvgDIoXkzyqBXy7Ryk8PmrGiCrnlv0KGR
aRqKLkBL0jSNPi4pxVJnDtulvMkFK3JZddwha+2vBQ3AcDSerluqD8bSJIS+PzQly5EFzWGK67cb
Gz1M/UWUjSO1KqbVjuiCbcD8FCQFFHHsz92zrbOx4OnsXsSepps8kvnMUfXgVqDfzxOINdTYFrzl
TdWkBWA/UslIMyCGXVLE4k5CJuWx6qc0tYdAv4TM1DuhW+a77G7ftiuMqnkR5fT8koj+JU+h/e2w
5EeJHABJlrloMMNSUIHl3s29D0E1eqI7jo4grrSmfOL1BEWs50l1sOqUfM59NsixjP1kpwt8Hn9k
N18ws5jC+FJnumAe5gXPsfHXhUgb6MmnQRDqswQ8xSIYGmIPFFibSzwabe0GCSrH2ful6xpZx+YK
rUTZI1PTupJf2pCOkfV1GfUuneGlrICuaoa6putU0KrINXxijn1SzUxmmsOR0AUOlpsPrGzfj7w4
nj22Pm7e97cezhDj6k5Htv4EPX+WYQa36CvG3n4ai6AyKuLSo3YmaTVGM1PbZOlkEoOgtnxvMp2n
a/pYmHB34ST6oqBCoRp4Z72oVtnFXMhzrwta1jzRZOn77flePWEJhe4D+zgW42xBgyAEmEbuCQgZ
5hoqmJgfmI+Qh9c2q6Iaycnqv/FE4Si7TTZqZqg30mFOLXSkjIyMhrOtMU7BdjbaCK6Q7yyui/jn
aWgUFwOEPocLr6hD/WMY0RzZKLsTekGhHy2luhX/1wr353N4NCH9aYsCwD32/kI4+lYhwVSl4FeS
PkaXzPTF14/nH2ek/boGl8FFlDmKl05nxl0sMUKazjYXeyBJ/a/EaU7xDV9EPvB4/2YigMqzS1N2
AmiL3dwYwUPvXWh+ZON+/FxhdNxMlntAvE3SKWi3BD7RZxM9kLczq6Z0rMODOP++CqSJt1rpChoL
DpOT1vI+4ffaA2oiw+6CIr8YrXCQ3AOf4yqdmBaB5KKpFDYN0KuKYyjZDkwCWvH5Ck8NFtq/y47H
x6wosjRT4KQu8sCYtrcTdQI3cdCd+cdyxpkEuMcJzvBxDua9ADpdVPzJeo46UOG7A/fhNGAFK2Fa
seyfYHPdo6mW5c8XWETvYe6hK1T8R7MF9Ej67L+H8+nt70AkddNIEsbhiBFOQTl0WtJIP0FT8JpZ
euqzKx0sNAOsoqM60ZWNYX6TuQTh+yP6dcl+vrfqgvh8o9Y2Ut+wyAt5TtOndatweHfrVk3N3CgU
B/OUZrpGGvNerYhy5OWH6eg0PKufAE4NN/RKS1XeBkftCwuKaQajROJbRZQ0nH629nrM2rNJCHOS
XhpaO3g37GvAii1B/8F92uI9vWjN/JRpnUwTZUdeMmftLNQKQC34k/uQJ0gSJ+vsBghe1VI/rOOz
k8Kb1Hji7iciG2Wf+6NnNPaSvAj6ZJhzsg8jSWZF0DMc1OdaIBzNlqELBUYyZzgJTEfW11oRnuKF
shNY1PrcwjbmN4gCbVbIStmKTzxZNtEQTK6/9/uuhbYra5wg7JgUPgQdL4mGnZgfKMkjpJaGKcs1
PXY81D5yiOiksu6O1mIVkMdF/CRj2CiAc0Ovo1GwwbG9mhGpF8o5U+kbO+FPqIXICYyBRvff7lT2
ymnZuM4gnngZOe+xkEhFseatRqiJUK9Ccv5Q11TEcQrww0A//honuWyJVxyNZ4gUsGyUVy8UfBov
md7iO3vc+XabgO8ZOJUtJkkvVCmdkFFa9kn13Ka/R3j/YoU0GrbH1Wh+h+lkZSQpBrGu2HY5tUzX
7nI9ypBkGMpp7C0mz+/dAOb09AVCw15yffPhMJmY2PbEUzHFBmuzUhnNt6tRjK3DZj4DJYqoP+3f
kT93128Yec59d8ceRA8+NkQcGh4ifZaOabfk0SpEFrlR/BiixR9hAW3Poz3bpWFGQoSNfOWX3tT2
jYQIX0DQYPyxoyjveFUF36dQF3ajAOwbp3g/ffA1phMxY/F45sVaSaVEMC6JuJ5+4DcLR0tDm+gX
+VIPrcsUVfHE6U6+GAKfMOo2oc8PvJyBVGXfhLeRkbmeY06blr4gOkSfqbo1vFuwP+Ih65jP5hot
3GCcBKbctCk+7poCJ1+Cx5TfRc/RLXtivNiMRHYWy+NUen9Ceqh4M053G300hPu0cBU+O+5UQF2G
jFyBoJ1J1NekUqPx8KV5Uq+fvSxSIUcGZohni2uqIpzF3eoQyK+qnNQgA44rLMKXX86o8eQ1mFvA
NjLDNI2h1faas3X3Rlk2Csc6VRX7ct4/tVuBENGefC8oEOj2UhshijHCL7LTKijvKKPw0UPzwrNp
zGlPgvbSGIKChKb7/Tx1KzrJmLGRbs1M6cMmv8WdHH5+loexUsPU8KzQFN2SN/PEYE+9rMZKXrTE
fdqL8NtlwbXZ+2n4S0YVG9+QYBNK4eiRMJyCEygr0CIvw38HYQCxcBEXMIwQdGH7tJ5KXA4tjbr1
yVKZUv6rQdoFPotrKSOKsQRcvWZtVbvCi2Ge2KiJECA0SZjjEWyQ8jj2tszajBinFgfKrTOlB7kL
mAnMuikJ157zYTSBXmqVWDQCkWzpMy1c88NviOjp9qeWfZ8+ZtpUdblWxCxb0clfu1/wutH5whWF
uurt8XAjdbK+064RRgWEVo2sIaxgOp1/smsMNjVQ5p74O1JAWIUyvxL4sAadqp0+PqttxcVfID5r
mV5yzLBnwblbBoRl0KNzFyQvfKHCbTn0Zg5Gj78IAsn5EZYT3VTkuou4X7lGUUMk4/K94jYmsmo8
A/CR7pf/RSdZ4sYHeqlvHr2Vm3NMcr3ePTNCh/cc3doJfZbT8pNDbRelbg45o3PAS/RyiA+WsJD1
0QXNaWUWyiu91Si8XhP5OYtFkEAgfmW2q2RCknu9m/CYTqP20/rfxHoW9/A7UsZAFXkko+JKqUT2
5VEau0TwWWDeuF7+0uv+FbE9sHHmaYzeQQud8AzHrI7RLfAPRodU0MH7VbWBe7r1vsMCYw5o1ewh
kLt1E6/Av/33bcwFWMldeIQVyZvbfjzwlp46N8JfiNDLU+rhRi4Rv1F02NsKK3EjGbKnN1JJMga4
IdmEcA1MABYx7SH2+53P1IVkVowR5eMCqL2fQV8e5qIaSkmFANND+if9/gZ0+pRmHy0Ik2JXS0NG
nJjxZOypG5mvOcBEZlbcrJ4M6PgqNeyxpmS8D1oXfgyLCktsk40ppQI4z5usjvfjsqH9zyy2/u4I
HvSdG714NxOVLHL4Qjj8tc5f1Id0pIcRSruMKiA+SMlYWQWuxOl+NWlZ1NeIeGnw7ECx4Et8MQsM
Ovk7F6klBHlmm45Hs3f4OPH4rQ+tPHhz6TIhRcyUgLtIdOy6R8wl1ULs2VSckCgOcCbPHgFGQVPF
0Inh4wSEZrMI3owGYUDhGL5gtdiuNlUcHqb7hBhzCNg567gO/69TOtc/UFtGMHFv2p6e2G1zqIeR
R9uhzQ5yWD6+X+sNCZGl89xhViiOui38H0SQ0zk2nEMt/h+R2zDFFIfcXeGqnelWDM0f9UHFHFyu
2yzhTCFdP9SNyNGHT1DRTOqM6KEBuj+azFk+nvP1h44FTM9+ZZe3dVYXi1SX6E092G/Tj+K3Su3A
NttWGwkacod7ZejIDdbWZwNdmChpTalKL5hDoqNejDMI0wXnEPjcvAYBrwN3EIy46B2a613OsVSJ
jbi708oQ7bUDKUsh+HM1EnzKVP30oDx3tpfYeRPJbd5XLe7rZFh+DmncgmlnGd4CFMe2x7d7385W
PzzRWAdhWTKVpx2+gtX23H5tbR88te5FAqUyPGT8W4UuyBvi+YTv0WbHdTLbuG3n9c9/970pf4CV
FtqKrMBN79DbC4FWM5kVKX8DHd6rZzwuxLWfBymOWHRN9yIx0IDqcs1LdpHFClhickz8gy2wdAfu
lbWZsKunSBtjoXXudwRg9zMpWQsawaBYUOyqC9qL9FEXEzKvIbG7grwt/lMSezGceNDurrYR1x08
wHFWliqm2VstVKtzvc3mBbFUdql3w9+/AgQLdtmWLNkhm3ti0/cNNtltlK8Trn611zcKqb1bDG3W
i58AoixgYItb4dfEptJad1RMKhxhQz44AS7QFkoIHUCSa+6xA4Mi7yk3cDT479nayxTwjffbWeuh
ZKBW8NX+GSJIKGCX56w0Y4dWz5rD2Nn/zOS0+6Q60I9p8AM52Pz5evmnweozY/3T9aNUgWvlg4zf
kiu0ulgEbycFhjUj093JXevO7YcbpFU5VqMnSTGTgPLGWVOiZmtXC0sQaqgGSpFG6UxepOafSF2c
mLBI6cvdUXUUbzBE9D5Os0lJ4GDGonTSezSsVtheJQneTj0gNBYPbOxvpU8INesjxshIxYk1LSSm
yYfJBkyyMUY+oJjHsw+SZx+c97sBFNTjtchjK5rgLL5FvDwI8CT0euYN6eGXngQLTVxqqovZ1oPH
L4fW1X12csQUFcNkT/UhzOVh5YXkBcW6lQzeNR0yWTd7OLWGraVzJbthL8XJX+tbASYKprV9m2ok
eu3uvSvVPRfbbSd63tmsF9b/SlvmgWGlH2SmTqb0CkFImhf7z7TlAjz970jZzpqcMWtQzifzhyMq
sEXZCUPsWc2142u06mrXeLDkXu+XpUzvj7Juy4Fa8iGAfxeUWp3JYQ7yyZivAfxrm9fPpQWTYHUn
ktbSilf3USmzlvtq/gjxU1X9tuLRFU3/EHXFj1VHSUwSZbTI+yLD/a5az5KbvMYNir0U4ytzpUJK
eP8bv51hHAYTxgi5DJOl9x5AYpM423jTfg4HWtK4QD/+4lhIpjTwoKyGsKl4YFvktevP74xQTqMH
a0YL9KF5GmVQe6XN3xXujLcgXbBdxnu7sb813FIuNHHam8T52fhECXxEQIc9Jow34z5yLzEuOw+Q
QLStvcx2lIMn5EotnwaLPFJNaWuY2VCOtEV2/hJ9KWRJYenxj2GUCY1NT4K57kzrvmjJl1prxzkN
omT4JRZMCPp8rWhMhH1/FjREJFNGNuYoa/70nX5FxPsIJPIu5jK3xMiQuVYE38uZvXV46TC04phE
8GbNPCg746BRdOpy8vFKf9SE0kBb/+1vRcEY85SuBHk1fHi1QaqyxAzghtTeefiMNi78cNJtvN+V
e4BpNY+H8szdBlbXLGFw/D5M0+IdwhFqiKJ0ePwxB8In1XpB1IC/ZE6QeqhItMrTf158xP9dIeFQ
og4z/ouFHSzm38Kp9H0el/w1E6NQW22tR8gFLU+QqJGX6eX3+nw2I9PkTNRYiGNn/svrAg9Ruc/l
Y7Ru60QDs7NT+OFT85+ZAmzteJyCie7XvYSD18V2ofstsbIIsETdnw+uocEDiTZGcXzS81ojcRVR
V0LDP+yqUU9By/81G/rp/IRuR/tG525yZYQYVwinlYZblimKw83CRbwk1VO5wmnaD1Fot6jh1yXN
AKfuyuFvtPMoptMbtu3QVzunEDbv+M81RJbQMil67sBXcpaENNl1/CQTiN7vRfLJiEPNIUpWP5XD
v13fkek0kaTL5X45/+IgnKEofH9Iz0tyiMIasrfnaqIOUATKPiHkBCF9s8dyAq7swHHEJz28hlUH
x+1Jyknr4bYGj7YnN4oQTi0zcA9X9yc1CnWDY0vMlmQRNzr7KO8ECMULOZwjC1No4mdIKbb6gOKR
MG+4ld9XfOlCd0YCdFWbQ0PAu7m8mPKzPKnw6X8G7yNCoV02nT9VmSpZKYSoDLFJynR5foggGlJV
LKa+3PWMD0ABjNUGMVMyjE6v9mXoEmHR5nBJYxWKXIM5vHPNim53hicx5X5uWdWatXzLPFLgrCkb
QIDzTWTiVEy6xEHJxXPUvLNmvJYitSWm8lVM37pZ6thr2qJ7C1Duewi4TU1nI65HIAwEwOBnTDtf
LjgpSJBbFL6grISEG7jFsCgOluiIUhr7hRSvA+1OtW0FdIcPYh17QJvARUEt3v2hzh6G5dmESVg3
5LzQDrBAb3CxIyiaQibGHfA+IdUUuoAEKJUIf/RLzdzJ6DgD4Jiv5AUZVMikgMuOua14Shzvc8Nz
wIWttS0Mo9k67WbyYQKI6HT/QZidy4gT134XUcG+kTbNsqZ0CVOFrh2f9kpl7qBs6KbhqWjCXGIS
QfQ8/nuvLtVsPewzrhYV8Mn3pON1Bp7XxYnUBycLwAgPe1xdo+aPa20fKT6zeBXZ6Ta+6eG/Rgtx
Roy2VKKR9WVvGPZFpvrh9VWjfIvem/J3Ppo8fTTrP6BzthTuctsvW0rUNGVuHqIO3exkEZy0R0fo
9zyBUNWymv/Qjh/lhgp3Bwe15SNBOBzj3amx3Gsb13xNjY4C98WD+kJIePJkLevbkQ542CqnAioE
0uv3850a49RS4h8wBXM1Oo85TkOLilQ4YZI84aEWtMMErmhbwP4AxbisAJInR8lPewTR0hHdDK7r
+pj4ykxRDL5MOosrXso3WfP07AYPuZo9LRlRrb1UOjH15NgP0z1GLBdzYV8J8oJm64dtP7vDusjI
37k168WgsgkdAlPoSgyABi7zBlldmmcx8OUbAa2ppfGaLSTRF8BcF3a3+xul9Ndpyovb5qNQqGrf
2qAqPNWdzs07eU5gYUmUPuO56w1akJy3mxKx1JM2Qm9292t9+AJ2aA1kR41zeEqHWIoma+7ivM0J
pU6DDeXe6ZR2ttnW0rGupZl5gF++Ur4VNjnOsAWX1fdy68Ed6Wqo3v85AnVrrl0+J3mL8YhUqQlk
wMaYggB1hAQixbufSz8K+f4iVAiGFPWJA8rEydOcEPd4gJk3GT81TX/q9w2KI1hf1cm8WmO1DLf1
/Ixb8aEUFwbNA/i6RdhG8YmLlVh1u66xkstd3H6nosHyFVDnI/ypzS4itWwfTUy/pU2gC5atYQut
uS9lttPfUG7BQYVSdAREWwH6Y7WNUCrvO3wirvntvnxHWRNViv4IA3TGyyD5AmNaf2x6g279AklH
r/KkD7pWgaYVdqESTrO4D4EZzyovGLDSI5NCS/HpQl0FqNKS4CGJ5oov8HOHXWkWNxmxsnTC279t
LZmSneZhnK++n7jEDGKtF6sn1C7VhZzr/hHXnBGYthNOqYmvlgG+AUD3R8Uu6hbjsQGT6AWGsGp2
UTipwwetu84mPEgLQv0CRwaLJu+Wn6fXelnKusOzXsGG1k699diiNhSFPYQiMgdY20UmNMXcROax
pDcYdoqPPj+VZ1UgN7bJL0fH+WjpSs9Uz97ns9xlbwOxRUFKsK5NYqgIlB3p7vHb5QGNwR+ta1q4
HGNiY4OHsZWjz9G7736bWGyVkzU2r3x/N2Dv5E+7bq6FbB0vlh2ux17p1Rs26ptFqVhEw/kgJ71n
+M2Mo9X0eM75RYfu9o9YTpuRF2rbqT3q76gaoNJIWp5LNZ+0LIwClW9GJxZyakvGmkrGKHCUbA4d
hblWEDAT4SemVjh45H4WGnV0Sqk2Iidgr3RAGs0sRqksygI4DyxU+32GIpyqtiFNwOUelr+MHL0v
ztqJmhr+kycAy6+TOHVqGehr2eL8r2WNl68IuD/fgEE9PoRA7bOMdLlEalYeLCAn8BZamDQC1CSX
QJGHa9jx097OWV0owI5/ljghPih82R0u81MZcaUJqA9bJC8fAD0KNN9O1dbmwB0XSNep5maKR9qz
QXzGYUaSgcGY2tXYz8kDB1BITHyiina/Hw6qe2s31n0lDFViNvrlNByRMtQ0hsAMsWIATfwRC51A
1V67LplIB3C7l+K4NTftT00IQDLfq8jBRlCOcNbB+wiNSKQuEbRwgAAE5zS1Hdi0ZeWfXX1ySaRw
muOdzn1a2pSbVNQqwZf6bpq9NnMDWmYHAqy9B8yi4iP0Gvt1a8K9k+y94FsmeoZoiMEajqRBUT5u
ksNNXT6tAMD1K+f/CVjNulIf+9EmfoIsD1enXMWAzyHJxGGRdclj52IYhr6GKjLFIJ6WTylQPE4j
Hcfpn/0JMNpYhcUc5mjjJtDk4m9T9/FVLluiKkWDlyCzbZHthoGqDTyt6/wJ/OuaXbDcIXPHjL4o
shG5xzVtH+uYh9V9WFGukAN0KNJSJlVy+N0Xvo4jdsVmobo1DH183ho5EDNy/irRUMb5YZCR1HnS
CqCBHtM7GsU6tEIRf/EgthXhq6Kaq9OCmwOoYJDgrJhxqdn1BuEnY17AQewPzdM8Z4qz0v+pBsZ6
8LljOQClnIy2EsepCpuF3mI1O3rHTh6s7GEqwPEjBHdvTP4vjlazQqNKMa2c16GPV04BJijgEAiT
kUulejm4eYkw0VZZ9aTBCf3f9CCg552zJXdPeyqk1r1gQBezb6fI72ihSWTJhUGlRpB1oI4lrls0
+vEyBbg1qUA4VtS0BiO9RuBYNZkkmOw9cocH4e4krnC1NBzfmNlayPOmUxIzhyjBHo4IxHEfmLEB
GhzvZoGGXb7gz/iOIXbzTMfNgrg0U2UceJ4nSmW7qu908Yt67b9GKoCQgo6bntj9H8c05lyOv+65
q9FqANwYkT6m32cdABu3cEmEpD1Q40qt2jUtFWywUQHOau5uLfKQYNDVlX2r2fxEACd+Bz1K+6ws
m47Mn6fAJNkm4wv4bbQoh7T+vMW5GDfNJiOJQJbB3QkW06W7kpRazCRoTDF922/brRXVJ2zmIJ5k
B47ATUZ7IDgtSKVON6B3dx3FIwN9Mba5pRO0jbcRXsdNNmbS+9xml/YzODCCoBYOGzSuTVJFdfNF
kPH4Zq85P+LH2xx7LmF3Ze4VBbEbFc+EqXjcbMfF28mhdL17nFeG8CuOZnbsZBUjQ+hf3biYlBfw
oYksbU1MjKC0aeQC7lN7ZpgAaCo3yh4/BYYChcZYlz8m+V+i4L1Ys47h+zxEIAlL5Nvf9trbRSt8
BKKTjenRBuXMlx/Nh7yLapAjdSsTWOU7VaX5uS4IfUshoVwhgn5/vnjxxd70KikJ9joI+JDdVHUE
YLo1dAbSe4qmj9jO8dlnHPy9waeFywXHbRVK15IXv6JBI3VfoNwtg6r+SS+0Fc155GUrGoZgO22c
6gz+Fo72mJ9eEHHoy3iX9NKzFW+TEaIckIDBJJXfApEebGwGD32IA/9W2CGUnHMmkISj3wgW2MQK
Il1Y6CFljxfR2YriNZBSMiHSnbxDU8E9r5UBfVMj2L0dHPcaqDIIhz9+QUUYAwqgRxthJYOJfN3Q
AqbGD67/kHjdI3EModw6r4t/L6m5BplsR0yflc+9ZXYNZE9QMcB7vr06YLzdTuXdjHqfiW0+bEM9
st+Su6mrvgMF9qBqPO/yD3ZGksgGVedeZPm5FRMZda0uAQrRHp7DofQLcrBwIU8H+AqkRYIaGVI0
V9M5oYnJG7ZCgA/YQUFpAJ6yp/SfwhDuhkYw2oAyFrkHx283ohdrhle6JMI1s21XckbwoiGjnPYy
/iQ30qGWi0lAcQdKuWsIFsENqxUEOS1truW8vX9XeruNPNh6j9ZmfaJX+vzn4PwAlJdtKnkAVw4V
0wExzlehCxlVDvjIetnLxw2tambRxvREseT/Q+kMk5J5u4+bouj3JHYR/jncswLcxtvjMdwsUZSJ
2SqjtbBqIw8PAxpSXkEoMc1smqMwbIKGxuRRIC8bS2S783QsoJe7jdDKI5FznBGUci5dX1aqM5+R
YvIxXroczh8X+ADsYKGJSACq9/g2BlFtd4P9S2cQY9VSqUL0kAj1/0mJjfiL5eADDvzpQDWT4Lou
bDhraY/MYwpWheM5AZ984kpdJRft6jPjsBtyaHFXpHwgTug2yH0y9M5QV3a1BqjrnPGqXI+x2d0C
iWBGsQI0Oupo4ezxnRF4q7CWIQvoPgWM2Hwf/XVBlgIpluKj1s5DJOifE0PB5ymCxCWgLW24rvMj
CsAxN6ZGgS0y+2LclRfES998G7jp3kiE28Fwi6/ICwWcbMzzlixclnXaXeHKiPap/mK6EIiqNiYl
vuAsLGcJl3LdhPrWguvfBwRcSDmTDp6VnQfVI7rQYwPBSBI3bZMgjGFbjsTON4hLOFLFIhYBLyPA
FFY62/PcLxGdCn+Cnk/hzlPtfW31UiVJUkbZtcopO0rSb1E5surNizIJTw+HCdo1RFLrRFy9HF9x
xY+iJyK0immWEJDy3x3vnetCkub7xTWliKAKIhEhnyVc3lMIQIqSaNetfL5ElTMK8AjXuco89rEG
XY/HOWD0mi6/eGxZRgLaBySDYcNIzox8BxRwSHwzj1eQ6r5Jsw7+vZrKrpvWfxVu6AtnUxEEnRH+
Y6e7yJUQWrBHhE5nTRWgx9LOihRyORsAkA2ED2Y6NFaqwhDBNoWXve5VdXVsBjHK+/Pt5PXDdHqj
xDttBg0qVRgSHRYStSgL5qEwhHCL3oOzFODdzzDUZgY4RLo1w+yCiZcNGe5Hu9omaznV1HGVp/FT
jPehk/u1AEOl7UgA6NjliLLxHiEUBJu9cR9ukZbUqlTCvO+F0b7ZDH/OYFgPqiMbWe9AKAHNeqkk
bJKYJ2UgpqtP1g8ZhBDzPX9IHbLmo6UOjjIi/KIYLibqngD9WvOnabKOqMcX8vGjzGfPD3pt0H4b
eIWRZGQU9Z1Jv+oj3eXx8XHTLD6vwXxnf7x7gzJqpn7+1lHkJbPjmn+QqFTPFOTKaI/iye5fevEr
2X6uHTNk5cGfaXarfy+jJUHNoXqaC0BAJJIafiWzcy38pPbvqa7lwlFz4p5x02SPTyhc95jJlU5I
cuZInTJjtnxiem+LINpyX668in0RuIwZgCW1Owydy4EvH/B3TKmtaQOgQ1SBH0BJ4SxNlehGqn3P
DeWGCaPZHql3dxcdxAtkNY7VhMFaTSPf1+JjSolnbOg+PaUjj7P075eH/3IXLh4PAi7fIaD8FsqQ
MnYYgV1ENBv50iPdC0zZFBe1Bg4CMYAbwoebSMPWQJ/cTR/bff/MUz5vPoQPMsU++TfxmcBn9YDG
4FIpPixeumqCd4W5CdNTb1nJNG2lXhx8/OJkxjICCRRKU/zbUB4ZhH+CRB9e7Xip+uNlsD0erIIP
2vNEljA2T6+fflHCB2X9DwQz4evePgcH+krjsvjQjtt9ERkO2v90IXSPMUr2Gyu9W62YsD9YR7l/
wGOi8S+inaa5CR5jBTzFgZXgY3lUtd0EIHssJYFzAghev40vnuvNwAj0jqClSVdgNDK/e62FUJSK
M7Cb1z5Mrn1unecw9BcslJHUp9cgMJtwvTn4fsd5d/cr4nv0pJcw9nD/CkgbQjt3g66U3RZ5faVE
8R3IXf5iotdpTNvZx/raa5TKK13hoc+FdzpLxZmVyn4RcxO+xBWALxRQ7xrYQW5D+v3G19xVSKW6
KhWT9ZXI87pTF0NEeWEz6s6CWbxS/CazNYW2BAYuvWGDJxrAXqP3lZ60+y19ettQla7c0ZqOca+g
AbmySNJ+sOlnZjT9I+jo4ZfMz9O2jYSppT7tQb7Q97vypO1Db9yNqqrJ8GmNf/wGIcr+m9NPUB5q
wQLopPAyOeuw6iS5o1MLfFU43kXyXxzTiy9TN/AIQA8D+GQCHpLUzDKzg/VAKXp7r5wfuStR77PI
Um0AtRSXOR7ww/Hkhu6yCprN6L/uphLPILz8C8eKSERKPHVB/Jjah7mF5yUJTD6J+y8MIvDAoP5r
k6bzDNHRaoN8D0Xn8b/ZWwJUpiIjmatMGnYKlYxj8o0jQwzRQ3doRl1KkKZk2vsx+lV36X8L5Lbj
R4cd8BLUCU3mRAaYj+ZC411D/XmHKW9stldk6g8LQvRCqaqSQJ5+EXgEcLIa8jzR6rkNaXDr+VI1
DAz3eQmn9ouRnE7nRd61kSFRf1TdKyI9WBVxWvRRiS6pRt217KtYFL47A+fHDPzFRak/DizJI6eQ
fU+q+gfUFFF87vEnURNh6HiiY9ogCW4dBS/Y3gXwOdUnHJiYrACI0hunIePRZ3TxcMjCxYW0Ms/Z
Kj0aaAUBLsCXh1kNQAmrLurr/tdKj7lk7VfcDl+9TRt6sNZRuwl2rxqvzOp81RIa+xsnK94gVPE9
6lxibxLrjQ8yVUAewz4DXmFVno7n8kwhiqJm3cBrQdPNaAVs22shiKHRG0jD48vV3lBgGtXHfdCu
IIEkoT9Fji7YEHkX22UbtZDG5d1QxX7TiYU68wQaggvHibjJ93s+NWex6mjooHAaARJwDwpU+C6P
EVtopSWbEMDPN3IcrS7PadS1cqda9ZYy1Lc7WJp3UqN9ZlQyGr2S4+WPNKraq+hCBM+vx+qsrrJU
/kHSGGg7r1qz+0XRUVS59AxtnJrf7CEEv7DFVUCi3Ue0LoLvTq6Ihb/0MCidzi2WxNEbrooxuHGr
9TpaIVNGZ5gDSL+ILWF/F8yQ7Z4aoiTki8YfnrNxIwo1ymjIkcwNP3Aqz4EfvXkoqjqk6TQDqfLa
mVTmxFiFfNQHeQv435NmSxR+6Zgjc+6E4IeT9KXA+YvFeNRQH/NTb9khhQR/35+8L05OXRmidEFk
RbrsnthX00Mm90wedXcfQHHbpkK462UlR0BPzyIP0SuKybatHYYjD6z100WyjXcF3gu1BUIuVDef
+qWvZL0icEbnAaDydvrwNtFhjDThyeTc0S9WTqN07Uyp1Md9u7YUj64JQhK/ouBioHVCt30IseAq
aD7sHeY+O9jrdmSgB+T7t8ECnO7mF1+ygLB2cPricriasDtPSbMqrE6RPrJAx+xhjuGVPZ7hKaEU
Cmy4G5k6SWX927cNVlFr6JfUjA92OHAnkmpNrgC+VIJgZ1qfZB3KSAbe5aXF4XThlUft2SNh1UdW
k1E+5IKEO+YJmE4ObpdG1KH8Uue01XfOnu5Gw641NsY7ebFTJ0mm3Sek9yuPg+THPVOHiykFMhxu
xXY2kKn4hlTvT/A4gHjF5EMPU1fOwn5IKFITbowI4+Lr8EIyDRGv4C7ZedtWbDeg3I/rjfICU6sG
SKFDgK/b1VQD0shMPcNokJtXwL/0Vsd0NZpvOlnoBgSVhbFXR6mUKoguseKf1J+c34QbilK9Cm4R
ns/DZr46PoBkjxCZsmLQPkuNw+18jPd5XlnOR7sOWtTuieQDA9Hy62s5r4hwnsXcDSpX39zermx6
ESqNMZlhwGarUFezftel30939oLqefQlN7J9Bkw9HVjvgecUSeXVKn46gCCHu3mY5lNE2pc+icKV
Ky3LhwF4SWLnDo7zprxgKaPiCgRnZXYjp3y39voT7vul4DegwPC04e0u8bvIWjvqbGRIT3yG+vEn
yP1N6cMcc690pxu3+i323eVH1DdODz5wfzD2Z6W77ZBGMYEWcjB9et1IQ9RSKUkz5pRFxCrIVkwH
rnY6NrxwzT9gPFxhIcujIIPLr38mX8wFXfFP7p+GFea3bPiUb+Ak3bPv6G8m+OtgtHqdyxpwBuPI
1XWB7sEdWAyKgHMTiVASr/Jbmk3GtSrMP25+o+eOyGtkmwMn7h9RKBAhZJ0cYNUL5V+VH+3Glp01
DDb+XtGCOWIV7Au5/pbqDUG6Sn/rVh6zlfzyZz08z65IrSt5nNZYaj9EXy6QvZjH22IqtIev+w5d
OPQMb1q0tVIFOVJzWuKZQSzdiB3h4Su4TbgakDR0TvuMuG7VaQ2DjBDozGDOtqfXVdj+PFDbo3E5
p4hwxGhYUTjhAWXdJMFQx/zBdWwBs2DnqUHiePW8Ns3jH+nh+p8kuqlimyCK7oLixd3Ss0ey8Rwh
NQVxZNeRnsIjoExm/zVkSvoPJIpMnM707QFIS/D4+RMf/sRRfTeXc2KglnLvttwMQn5juYvwCy7+
Lxk0Vs9+NA2WHSW6jQBbj9mkStR2Yk0KcViYGGnz/C92H5PeeeM3B0HSjtJX0UAR5EdPLoYuOm7j
eENUwUKfWrUch1BYfEq2cD7NbhzxTpTuB6CeYApC39RQ6DzXwYwIhzSNqoU2AROyXCfpIYr1eMpH
lxPT9GrqZwwr/UoZlDZGM4PhrjKpv9RIX2dkJdD/wc31iYS82tgH7h+ofTn4InYQk01SC0yiVl0j
rJ0cM5XhOkUz9lSHoSsaKen6Zhql0Xcoz3vh/jM8u+3wPJ23OQ3h/dcuRZTUB6n4s6EsMvICOCdz
32z1p6cePeJvN2HiKaVgFY6+IH9Y5OIJVjOSxLoj8RHue0UytQubXz+17jYLab2PAP3vqDkT9GSq
g5BWOy9ixRpTLun1kbnr0lvDfBGcqE9iPUXMtOipMz3AH/RebQsBai1H1aVl+RFeim24UtYr7BIq
jUN4CdPsbcREmxR9cNKsXTAsa+QdWhsz26vnT1Iw6JOmxvWh8arFmkbc2P4P7zxYxU42IoXmlIyn
7+uI4CI/jeWLv06YymBUCoGtDtWlBbWSa9ufxU1JJc70pdqUhPe/8nEICSV/0sAaUcVBwBs2wUB4
bqHxc8oCsQXHZtRpEM6u22qS/3y/1ox5+bjrzQQG5XWMet7AiIEMExfhQl4yzaR5piHYSamca7/y
8FFyfjzYJRmmFrBr8Mu2Co/IC++F6R+ypuP+XjF+2gVpXmniTCYxYHN4ZBuaQlDpSFneV5DUJwd/
1ZJKHi9wjBQPdK0r4MAT/RrHReYtHDH6Wyr6GJ2kd8L+rufUR9ut3kj2MWjtyWHt1l7xV7xiCc3L
K7gHa+fhIPO6INmgo5ke0jBijp/qnNiSC+QJbpHDiE5fcyjBUkGVgZKYh6v7MFOHfFkaK8cznUbv
16LouRyCwzvWDAj6KvtWOKmWZyBvIflF+s4IEZ8gGjixX83PpHWU59Ypd3ZfXmTIXjDqB41y0NbS
4m3LcRSANshSLOxdmmvwMx9Tk3ndtMf5H7uKe7hqghmkYMF7bIXzqDe66y7UHnz4kOzp3t2S92vR
GTEmyJBdDZSNt3he0wN76PdPGWpQLCPdvUihQH4gm/NXgjWzl6SmbwaBeBA3xeA6KRN2RNd2aEce
Qzlx+XOk/cLT8ye9crvduoK4eMIumuWqVFmOHteEk5vttAILi3rvGEyy5FetIR/a8REhIxrVhPJp
bWFhD4xvwouEiOEAz/UKwQPhrTWevGJJYL+CnQKtSqZztzFbhQVNjEHDDrxG9t2ITQPAcPbxsK8P
qJZIkhabNVZPhg2cJTwdTG15FP00YEIhMc72u1Q3KuDZ82iGUXeBaBqMo5QBQudHDfFTHKa0wx6f
RZyH1OQsMWsD86dU0yUwWbPQHXjM7osp7fj0RTFyS2vYH8DNRyPMO+/mPd+qKsrOg/cS2Nybi2wp
NuQ+BuyM+QecVdbIUqczU5hAhvXTaobSSMsMDYXFdiWt7KwdO5DKTA53ZbABU+aqW0eM4otXzxKD
DWX/fFAy3uc9UfgsDS+eCM3lhVNIO6pJHPlOGBs2kCCbNiejUBHkDoO+bEnT+pdXo+v9nBQDytKA
+OThthpZmuLeRBm661LbnZyKLl+iTYttugn43gPtCAmLNlmfbwt0QiFyoqj+TgDJRSec5paV/QuR
LJ661j2eLKizNrzA5GBVp5Oa6+dnvnqxI6pZVBDRbbuTw7RUmUh7xOl8Y4Q7UgipTnyq2zgIR3FL
Q6I+uWxNCBImHFQYSXd9Dz12oG+8OykDA8VPll38us34wQcipln1FVN8A4QcjTj3TX9zmweHO+OF
q/rVKmQENYUHj7GhIC8DlXwoXQrT1Yc3J1/azzFzDz+dv8Tp9PsCPqeV9RMJN/StWjDr2LKDHbwH
Z2o7goy59kJCass40hZV2ewCHQLLu56BIxTguRC4LjzpPE/Ow1M1FARlsp3mub08xuEpbqrMIG5X
cdRLE1ry9NaYShxFbprXusX8xWb0yNtUGfm28PbGY74qoXQZPbrI9G0GeFriYO/rfTe3nUjiTjLo
ZFsM8fznJUFTDhYV8Kul68x/srvLeWBfSpOnUfmz+eqGpgcLvwMzYjhP9eJtC7JGbHe4TCFLkXk8
7j3cFBUpETO3S9WpGy6L7yUO8RfDBcXD3jyBI0mi8KkhKMICRvduaKaYTzppXU2UJ2ARDTLgHRHu
qZvBwWJ+U/GtrHUcu6o8SlYeQUF8EwWPhME0bB98eb6RciIYffSUCKZFRSuxsDqwYPVwxmy+lBQI
4eFO1D+a5by7aIaav8FwolX7FaVgTmkko954eMmVReRQ3Ssow626onLQqurNjzO+Efn/bX8Pxm1R
N/H2hFicYTn3Ia3XTIShwC24BpXfOBnHVt5On58QyfidR+/Cuz0VpqCH8ZocXMqSaus+1urf1gc0
qMhDj5oBQ1UM8OcXHnvcgg+kGjjjueaHGpYiJMeBo8CyWebXOx3eB81SOpSkfbfzz4dzla86Ek2b
PMKtlZk8vCVlYGKZ2fJ8vcDium6o2MALt/AkEXrsDoGWIoRcj8yz8Z3JFo+qtPEAKXb/1+qFlnry
25hPYm0D4j2kEJ8R16QlAwO+WdBAnczohoQQdeeAbNLgO/xdELvJAFKWyF/S9037Y2+a/z5syqi6
0kiwx5NcqLnbQ/rSlXMfVp7nxYooS28pvsnFJlJTl8g4wJEa1POVWxVA+VnrH3rG+9bbrzlImGs2
k1DplEW6mAKJjUoXkgUAW2WyDcadcWZnn5E+G4bj5lV9z0BGvQqx6IcdnIy/yOWMMsZTR5OgVpZl
ldlqGp03B82ZywcCtgf2fCIfBpQeUHCplGr0ZxA8WhFePOxAd/sOGQ/vLhyJy4QqzLPRNKFiQSm4
UddIM7Xl1/O2o0EyCSjfLJR0YHzek2/nwYgc/ehDNv2TvA/R12jEsvlxWcfQpWs5JjkXh0UM34jJ
izplH0EErLsU5SFXQBZ2PAi5tqkhdqQF8lJxND8s//TFNjnjEM+AbqgDo4Lpowc/05gsAgNnwajI
PFOVgPw+wKUkryMk9Hg/fbtCjjpOLekMwp4rNxC2SgXeRdCy1SiGLVSR+cWOw/T3sFwQbtY+isr8
bggvpnqIR+Kj3wM1SueJERq0ys3qzO9vjH0TdlEC4fE/NyQidto+Ez7gpZDYM7W/9RySPwYvwc3T
bcz5+SOP/IG7xN7gjIvFZI/3MCRvvKCQNY2KtYATZbSzp/kCJ4trur8n7fGd7N+PYyqmfhPdrU/o
g4KLimIgtte+cSLPq91SxsCJ6yeKPadgRfTc+D25M0dAl4bA9d5tNXFkCCG4ey9P9KDt7SqKio26
htYgkY0vb7EQ++EvTz3DTwLovERht325vlhca+/VAV9GxQ2xDq3HTA4q54/j4Om4TUsW2g3A7u1z
XJMjb5MTRpDqh8Yd9iG03qsV9+HUmJ9ynxithWw4JUpehCTd53ekIsteczgvbYAkT6vhjWX47ah+
OfRqvIj1d+bKHOpYAjFR2SUCRtrCk6wbHeyMenA5hjIes1FO5vR36dUE9pDE0Rf5uiI2Rg/2Vw4m
0KuEFWko32GqBtpUPx6CBscBH+98KcBFUUoBedhhqSH9Mo4FNPSiX+muqcmMLG5woLSDFbY3/Lij
LnwDT3YNuRELXK48GYdgVjvYsXHYJkdPhLOzZyc8KsGC0FKQwR2psE5pA/wifGNILcWzaBTYNk/O
/4Zr1YUcJWNdDdIIrW0jIaf4Xw6JmP/vronvfzJ/5Pj/5XSnBX+N2Po74oV6Aim6EGunYZpb6USH
PvktequjWOMwnRZYduZTcuylZsamIcSYaTQ3bn+Y5dMex9Tryt3D6I0tgoTlhO7UZHkxm4zHj/7K
QzWtdr4Bi7xrA6eC/o5EIcyPQsLS0gTPvxCbbBzP8MWai6ndn5qYH+824j0qT/P4aHpzWKIY2Aq7
V//5qnsCWrc3OSnEFlgVYCuiAJYSSn4jwzVwz1WZdZQqfRwZUidL/98s7SkYi2bjUsMn9dhYSZcu
Lu6rLedkQn88afcwUqH4SZ1bkvJtjxAzWp92u6leKocVzuQvyn5r0Dro9Xs/ZtaNmklfChhEZEIT
LQemtPbJoHrKcCfShj9MG7CQDcj3eBRtvTE3FijWUKGf+wBFYp4/b26PxNm7ERRCWzbS2Xk6vGu2
RPDJEKtm1DC+P/EwJ0MAu48Uqyl18ymCemMhrTuscy5k5kiV+DVUa0qaYA8nToe+XxfAaKZv6Hq6
mdsV2OAHfIWii1HWxg0aL2/OdVnxtX9Dm0mOqDm0y22RnYMoWUiRxntgDoDwvyNdw4xaCEIx4vTo
SA2h5eMVP276L68RKE+o7eKccVSxDip8YyM3EXiOlKFngsXHiWUPfOo5jZtEeyh0pdQxGYlH+Mvl
sgGpuoMP/Y32X1BfaIAGm6vcrOftLJ6tpV1CUQsRnco3rXoIJfNsjQx6gAVcvzv5mjAEn8JdtfS2
/ly+w+m+1MlwtR/ii8VGygSfQVeH/9AM1qjkhOoH4XoAtS31dGxhG+MwdYNK9eCVwXmWjEuEs9r1
YkQGgZ+ZBfHNIgi8vuYWEPJLMxx6HnVgn4yBpJIz79wS0u/f9v4jJyNOf6/w9BduEcHDRcZg8i4B
DX/OUVL1aPPhLYZ8aBBZG0fdmZf0+xwccfojrNg/R8mLJED8P2uGVLlb+7DvVnIJxvrpwzrYvEBz
7xa0lq2iR1PzdUxpZB0slHTD0SEGekARbFsy7n5e0z1q0R/A8xZ44K985sv574gXJ4vyncjekE4j
qmsiClY6Pf1tzqPaBBnPBCzbZUq2ga/DHN+J8CeDuTvVB6a9tnCrGf55fxp4BsUeHN4qoum8DKJ3
mArICUx1+UQtIiFsEr8xYFQDB32xJ1BbgU/GjKJ1oYead+jyeHjJPj/6gwzESeYNZaWyrqjI4KUm
7d+j3UETD+S7oqwTXguu/XB9fl3g3Ij4ZmCWtS/Osvj8UVpJrjJhkl5VYNDa4aG2npEZHSD4T8Ov
g2zIpYuXXukqHv8PK3hIa3ubSxrSm8iMD9Gs/yfPPCcijIYHIZqj6J+T23lHhhf+mZ8ZqFWZcXd+
Rtgm/NUgGhUnAkbczzwwNWPfeDemnzsG9zi16FDftGAvZuJwA0Gkrh97rvM7GXAXKkVNE+vh9J0q
OvWtl1bD9bUH57IKBI4LdNKl2XuOfv7OvrKhwEClKlHARAWW8Ohg60rKRVf9jjyjdD9JaRzJ2aA4
scgo+sFgiC+QvMQ9zNzI2yldC4FJX7ofo3f9FDYCoG/YVIPIHaAr/ibiD+jp8EwAHkonnGUTkFhr
Q7jk2qDsIGna119x2tEHIpJg3/m6cj4uAqblA4Cs++0LYRfSCSyMeU0XLIuA+qjl/CTPhT+3E3GL
QeIVtZZ9No2hlFOaIy8uiRSYGbjiaSVFKgtMR2+cfih5WRhmafE2kvyqxRh/SNprxZDyO+ml2L6v
D/qoLXmbGeMvLWZ1pSFxxol1I5McHGjWw1ckqcYNPr5N7hYE4BqPnaUcaSXFI3hsFp4O7YcNXz8a
yDxhXsTZ1MbDYcxhn896PgpoQaFr+X4+d2LQx0A+u0d/2EEA9Ain6CIiI5A+URkAf60C1wdudxLa
kNwRAidyhyrTx0WZW4lHJDx5N2BTnTq9vjCmly1Y2v1RUXf0OSWIiz9G3J28xbnOQsT5tAsKU8eQ
w+PspbPjgCA3xH5HRExza+OrGVqPpOSeYPcLRQLAAi1Ekc5+JA+FQeoURSQpRSzCu2UGywPxcFXD
iqfaq1hj1jqTugIXvEQbDaSvNLtsRH1PzOAPAPa2LMuBkJ/EwqAnTnKJ7a+yCQIIiTlzU1Jk/ltd
CIWhnTYChkJ09rbdaur4lrHBXRqeW/sclYaOwvJEuH4wmCoKXU27ssvekRHc/AekmGWQ2TE1O+RO
I6gE7mI55lFVcdMwvAb+75KJc2Nu7g5vWV6t7Lxdy1AQ24AbtIJAIp9DqvduONWTz2gBOzi/MaG6
Mo1XgbuKmgwD3xaw/9HwGkd8/HPXiELhPcY5JQXyZ0a95kdxaXIBPLyS6eyJCpFcAeyeLPwEoKRU
cyLFq9TA9p340nYqJpiuXGc2VuUkeiOoDe2h6nGQesRODpsFOXxBZGVqdiLeuenvTTqzPdT9U8iq
u9IxofGKTeAkSGVhdCmxcVSFRic6G4jH441TmL/3iVKJ+Gd9hET2miES+zKOz6v6Vy4DVsk+wamf
A41rCByd6bexIzEQR+b2KDs9D8nJZnbhGbabdoVuMVAKhV0KGnXUozn3k0LQcvUD1JcM7YGgazeK
MmK+L19HpS27vRjw5xxTdFnwI/aAtlvrsgEUeuQiFsJ70G9GfT2qV8ZjcGMT/HMaCxWCXHst2s7I
mLd3BOYMJ6GpE7zgVKi3wKt1Uews5o935CUf0fBXqj68iKSIoZwlFHasZVP+Em3nJBl7JNkAwyBv
tsYm18JG1PN3n5lHJZvAeBmLMEB8uuzY+UP9NKsWN0H9atCjP6dTiX/txcoYgkVqkQcEvo0uUpQy
vgfSbhBQhllCRNaUEdH0TdmTqqlbmlcCH/YlHU9+ZnhHecWT/vw6UzowXupuG53/0IV831p3VYWM
pqRdMKR/d0ch4t1zDop529qOEBAGmOlgx3WtAnQm5kXDufnGbDMMgEQwVvYIINrrFmBccgE1SJWv
0QQGQXJB99AExVIbB0IEeFnfTjOMQZlvPAlPwI9OYVlq2La0ObNY50y5K4o1stDjYKmq6RRC3VXY
oTpP8lvRk2l8cHQ8N3QLbCRwi6xX60krYh5nEbKaI4RumzCksBaaSFSdkFnUnH9V4kDfJaeyovoO
Wn71qgEtVwL0r33UfhHCK3g7TwQ4f0YEMe4jqPGDuTZnv0vZI2gMRVYVDCkP4w1xPNf2zL3+o5Oh
tPOcItpxOoq1pS3WD7KXMVNr/39wuYj97fbmahuFcPAvBGA4LjslK3T+FPo+OKYoAoII3yeRhRJ9
Ho0OAtGIjGD7ceDLn4QcYiMtZK7LRfCp+Z+cBGGeyTYAEttRYucvYez6FbdKo//MTloNfjsOA+t2
JKxSHnnsxo96uohnpqlVXSMFbpXMsB3JfQ2U4T+3D4rAnskO8t9YAgtxB5LL7V+vk4cIf9sHh7HV
MVNf40pMbaqzoP5vIUR3PRtEO1s1G4XjNsmZFg/q0brT+lEcNMdmBKaGcHW8rrJBT5JHuH4bx27Z
LE/efdUPoCBUvQjBkf0DdZKOu5xIMNGZtA6eT/m0fbUWdGtujpD/uAdNBfE9ARow7Scl/CXKc2Fr
SqOpC6t1lp2YCT4i9RsAJZ/R5Mb1qmVzKhOZDHpYMUX+w0tEpYDRGo7UaQfjx0ov+3dDxIY8z8Sp
E4yIxaTkapkXCl0mb5hjjWdkp8VrqT0puUn+ENyOe1ree5A3dZqzJuSC9/kh2VaAhCNkuRRjW+wI
sDEDfYG+V3TO6jFNGTZLPSMV+71qNpvjX0L3FqUQfEfZpHiuFZenYK/uEfJonRXy8uSP9R8+BTxn
YX1auIrlSJcsh9jXmuYjSiuDY3D9vS0kmcYYGkXycRsOuLVJwFSywMb+ELZE/eEztlLwSGUHOv4W
Jj0ID3ZNQdgJmWlBb69ShrqXAW2p8dHTYx3bcSFJov3Y4hgaVlxedbhoLNhdt3+omC64qS+fqwmO
LHtKAmP8mmRU8cLqIr5adlERSRepeFy5zQIONzWhtgPMKWE3aIbDbM5VFXWc6Z8Izn8rcUOFfCQm
bAQ3zsrlp2XGtGcH5at3qEeVyraMmt8OlK5lDgzizXjKO84FvjCfJACtP6EJDGJIrsGeVFwjQcOZ
OzImzR+1wjmvbW+WkHJu6Fr9Qq7sa1F7majF/CbJ7QHhMmoT0hZ46ddDewMhtqzBHuT9Le/qhSLu
J9MlJ4WtCi1RxeRIjzyU2ojM0cGFRGcR624Gibj+wP5Jxnz+N2irQSQuw53XUKHJilkSXkH4qrCW
o27uQrOhS8Gye9uHNpVfVII4YHVmw6sB+mhteo2idnwuvOPvIGKdussC3x3RThgKr/WeU9j3V0C9
zA9pIsDL1LrKZelocNleOPP1Cz5F9F/yjNQSQsMlTQwnId3/UYodLQwry970aXBUU7IO+6LwMw2N
JVZeR1yZI6tRBQKC262NHnpp/sFcv2XY81D9Ztvow4K/eFzkmB85eHCKsC3HyMr3XN0kFcT//3sZ
a3lfo/3jjqVHbGaKgjnP3E0WO2F3aYutcTiECHkNptmg2MiapbCNkvU7e/+mZk7LXPLFn4bW/c3n
kKWJeoxNAHPei5caIgyXldaxmpZ22QBbn7KwLriV5r2o3xGTlcd/ekRfxS01rNegoJ9b6Bnr8SYJ
GC/iExO0hugixh2V5l7DxPhsyuKoouJMGrqeNY2In/4h58Plf2iN1PBe5wvl/5DpOHdF+AhNYNFO
qggmVVVd+zt8eHr5Oi+RHZdAbFdM7W/oG1zry23UwnOYy9XIj05CTH9CwsUx7fR+XM+7HQhiaU08
BGvyRpM6wez53R6CxOTBgSWIlE/GYlQk43bKguE1D7klqqviRqR/z5z7ACsNr0K3FB2iwwYE6MQ0
zWYWBlwtvCkVhna+R0NFNm6NUKxrfmWFNAhnll6IM/RPgN2xW/xkvOP+CSanoDU1ZhJIcrwgU0Eh
mx6hocut7wgDjZuqMfilNmPrJegJ7jWkYgQHo2Bimc2elkoi9FNnapK4XqUt3WIYy/yDOnV+Yj9d
w0EU76eDD0cJv5LdHLDQaiyX1bYr3Khe9rLvm5MfTo3XG4ECGWEmNVGUmEjRd4o+qOaR8WEQvugh
4sh2wdDuK+cHAQMtJMP+EmcUY3BGa/z8UblE8ZWk1P4c3pZXf/BFJPSygzyK3sWULglCgXZ4RUlD
LVRABEYDgnxHSdb+k/wzMVT3mLOH+zw6G0lxCCFKXP0pY8V6FhoKKzCkU3kMwa7z52x64C7or/G+
2K49KhLTbe29yf7S/tL6gkq6TWSigfrkM8GQFemcNRk3wXl9wYQR+CNoG/JJhLm4BLFmXRnWYz/V
WopU1sHLAoqZmZdJwUUUE0JtUDL/3KJ9SUMTIqY/UkmO3bCFs9Wjz8/BXd2yvCIDVgTmK1ozo9zc
ETB4DNhFkI7Mz998qBuxunlI0sa7K87LtsiblG4ACCdVOxWfpzU9GCpfdZC6GrdavVUMN4iyCLTD
nIGLhtgjw0q9j25/5xcC12U33ZNvB0khoqnZWt8VcmTXAMRytSs4mfEVSQX/67L+mjKe12oY6oE7
GhUrc5hMELbbwSOONTHtQxQBOLyj/B5hzEkBL3vVLxPrF3g5u6koQYeTgmFTUjswkrOT4Hzb/RNM
yuyFE98wKcex2JHUq0D788OfNaenzejDUVez2+Q1t4XPT6T0u4ypp1EIO8R/vHERWho9fDy/bM9k
hmvvll/dnLioVr8Vx43CPgefI+7YNOczQCIdzQJETx0ziWR6P6NOOjkHooOZRFENiDuN/hsnuRTL
xnivqwVZW87JEAIbTGVs1XoTQuxB3KVqWHOo/lhfyX5IIrXx65epu2fTzeEtCg156AWaENytD070
zIuv7CKS7ZvKsBCat5+WUzzr6qerQ6QCsukK6KIi86yRSxV8oH23dUY0vYbZywKD6IorcziSgeRC
Nlac4Kv+wENaT6KRepwRr0YkItHeunR9cZGmdrFEDeTETnGhNG+kf+rnpv9Axtz5oikQ9qGo+KhG
lZSHZy7nidYBhp1hJYKsE7C4JF4d092GHqSkbdei9a2rHAmFHe6N7AAh1qdP278u11S1orEHM4MF
frLuMnidSG0VknmuOLbfMdkTAvU3rfCvV/73gmSDC0jZcZYznb7Koq5fz+znlZJq6MHDRJ8rmhn2
FKqIfdGiPD6aiFfWi/Wey/YKqHNsRTVUtMJgf+haRFtOjST2/AV5T+93qCUBir++YM1aagrgrAVg
r+PBFsSpLmsmqneT5ki9nHe2nC9xAEJSFK5ydzrxVZBtBvtx3IwmejEUjPhFvE44Dyan1s9DEkvD
X7mkQgOu+M1ZptSsixUEHg12oubiDp8cQnWOgZxVJESNKWZuzcyiEijIbjBFZpKiF5YQdaMt4k/v
dS50MY4ZtjRisP7rYr2x/jqPDVY7tYFYfTQRropb6C3m2JJmT1RSFSIOQsd2tPHPi+YsmvrDQlDM
IrAlD1ohIhFjNSoQwb59RWnjbEe1ZrmlIABCKRwGKMSSmhlfbdsWTkYl+vrkfsDMOHMRXK+M/JGU
fR6NkG6G36KnJssCob+pJ/nqAAfx11V7EiY0mjoLkQKwxt9B2Y5GahJhI2t5ltJb+UtqcQx5nkEC
dLDMBE8Kb7yQB+Xan0eo221tqrrNMQg91KDop6nqp86GF4QQV1mXhQvEetgiSiCCwL/ScFl8boqb
HRSkMSJC+BguqPA+6Ecc7vVFJA3awQD2fHt380wZVWGfIj2IGHfqVTXaXuoi5DW5RLtG+qX+rZHD
K7J/W6nchKtWbDlMtvVbR/rNDkDQS+DQdVMHrEAGjAAaTq5bWmK/dipDXUnLd7mdsXAIAX4iCDSd
Qgsv6hlrh3l6ybPhFb5aRY0UDPwHqQ6Uxuf+/6A8fItATV+rs9NaZ8gTVP6Sa6Qa4mqU24X4om4H
FLxHiWWHzhN8OlJOi1+TITJmVoKFfRfqF1ec0R1Ibz5fyr16jwGPXAGY+OhX9cm/lW+0lIio4W7f
b8HEZrKXQD1vIFeRK/4SgGJ0gZqaV2/r4yxN3G39z+QokDBfJX8rmuW3XBEENO/iR/Gie35R+R7g
NVmHc2TeM5u8jIX1i8J7FFgGykh/+OuEzvEOHl4i/9t9o0K2wqbOGDLkqDA1SSHEhOKP39FddyJa
2CpESKSW1ICYoFmsb2J3KrSxK7e63w1AmjY5ITk/WVkLmKfl1pCf7dPWgilRfHpqkc0i031z7qpg
8EfP1mvi+TWIXQBmECr5cBzXXQIonKYqZu75HjGsbuDLQXs91lyVCTHzjNnv4WAB4a1fqeIVMMMh
fARNZ+9JQsnoy5UOgimP5MiWSJxeiEzVyY+kt7XzYklYU72fdbe9tr6RCV2rDz64YqsNsJKImTnt
mHlEkmHP/7hC1kkaifdKK/FUSOhTB61Zfyv0B1zF5MXKaaK0wH4xHZ/F1tZg8bX2Ut9NmcgObp9U
ELGne0KAKx5VEiui86JZU+oOSYMEEpwsv/pHwhu6eNTjRBdOpT+IsGitaNGsX2MGqxXsMSLbOcyZ
GbmIBu9YCMVDM6kosRGsRHBD+O7Mwre7jmF4MHUMZhoYqp5jq94qrkSwlRfbt6Se3wpjcFR+OQOM
K57bVRBaz2DRP+1u9X0L0L+v4nNaLy1k+QXphr+7Lpn9PhJLcmXyokaqp0FFDOHLCSEs7wAIrop+
zYfnTlSD8w9wQQMJS/Tlx1tVBRNsODpvYlw7hW7cchr8jVjUPYL21sIy4GDhGArN3f5bt55wbW9f
dcWaQ6cTbAAQIkBGNaNpwOnFiACY6K/CDuCBSfdbRG689xDWQMyoQUxybUKR53sgRhasRceNBADj
gw6XXM5lgkuyz9t+5w1kEq2Kc+AVUejmEBu53ZBaGqn9l4IpDaT9ROiSTj3aNJ4YwhJYkTEF9yTX
dJ1zrNxP6Utk0dyj8a5Wz0jdd4qFnIs0JkovAlLUGp7c5wy8TweZFNplDEugHq3qM3uK+oMf068u
x0bOuLfqSP615oZkTslLj014b3rcPlSwq9ogsa0BQvtWuJ3rTPPwXTk7BG2nRBRTHTHbJ3wyDgM/
1o1RCPRYW48r0PV0810zcUG2nKUjbENiVNKJPSZEpLab+c7iKqbp+FOzTd832Z+a2n19zFA5rDfx
HOzp4KEo7jW3yLdyV4OfFd8L1jVxb9s/SB2IZnZBkKIPkyzX5/vq33yuBbPta3fFScYZIL3WPoRg
RMKjWVBvxMZs4uIwDJLvfrgZFKHL4Dx5IeLcQmW/tPddEsdQ2CbiRQzswlR7sqIBQSPdvEkNTfOM
+YSvQpAX8alAVB9NQBItyNNRjiiLrmcyrSP7jFZ4KjsYb8+2bs73xDqFBLmzhGnYY/tkBPriqyf3
W65hiuNPbsm6IJC9lv4SPWi8XS2uWOGb/rWAzq8UF2jw7eR5H/cmn0f6qoQXhyfp7LuzoxhHjrI7
btPVFClkq6NCTWlhC++lt+t8ujE9ue76VinjgHy5Wrd2352Ozi+g43Ty4F2iYbiZyMBqish3ba2Q
ecd7Uv1RGkzdHIUDusgTo8i88vWbXoHyRjab/7Z552iLUhYpmQnnyDmztCM+bAAwPCspNdmryetG
0ONz5ffNhlMsclNnm1W/BzCM5P5dyUKIlM3lVC1ZSxkUvTOoo9RMi47D6bl6HsZGbp+OyreaCVbt
urv8euW37849oeuj3ruckf+zmnuuhjfiMUOGz+K1QCRhRpbSoWTnRHVH0qzks1YefITKsKrBKJ22
EaRiwDbWxte41gWV622BwhjMxuTrYhN4xF2Oi0UkG+DGKDL2nO78i4KiARo4vsYLDXZqUJiZkceg
+it9k116zSSWvLG04JIanFq5HuWmWKptzREvy9pfUV8Ti6JeHSd6RbkLI9mBsa9lM2IhcrZmlHC3
VBwVj6yIsgS6T9ltKCP4qkGlx07C9KAib0J2JxX/ZSCBAmQvXYd3vcRJK7uyMUFMeKxuC1tcy/7j
isDXRcPWUYabcCkRLYLDqSukO3sYzft2lPDR1T5vDrlNaj7hwDQOmsNwpm8kVPK/dcb20tvp+k4L
rBt1FWqyFsv4oCeBjlZZzDjav50Ane+9F816lOIK5Fg5tfDhyUfnp8GiiFj3PO3Fq/J1YaZ4y23F
/m7S1qRuDpxY6G9K0rk0oRF0syhUZ6Y4bTmft5j2Hush21R7TgmDxyHGgfY4Wja7TkT5w5E+VxPC
/eznmyfYCHLtG+/KiaL7FjK0Nb8nbRt9Oo3IKtkqeNL/F1J//hEHU8jnVxA+/3t/uB+TfkO7oxdd
m+aJNuZat+bC1dVZc0H6+9RR+LijIZBw3R1XqfNbgL4ZauE8JiAt17w5DVD6Pu05tIAeX75OQWBo
8Ev+B52WQ6e69Y9aFbleFRwiSU9BXMfjUvwdPpGA3VvEaNPNd0mvk1lhoJSi5JHYLG0Vr3ZPipQ1
7PiIioZzf2aU+liKRPzONWfJxFaaBCeuDCcpJszhz3V3RPyLmTB8ZCLnYOPin8jpt3jVhbaL8quu
rq1fcZS99aQpXA2Ya1zyk7x4HNI00Y/m9Xm344hM0k6bC7X4BobOQDVX2V8MCLnBvNnA8yw2vIRy
ovarjbCvGh/irVQz3BGR3RQPU8U+6vNfAbz1RAT9VuWQF1jrLbKtOs60zfv5hfjo8kAGf3oSLhyn
tpAXqbcsR6lgfjIwNNLYDabs7O4Dxdug270u3slFGHca6J7Skh73Y6hrSIKm15Z6fL74pTv2dLFD
X5APPqG04lvm+Lox6GTmZG5VaonFIuoXz9LqcH0KRyWUo7G6M8UShTHy/7qx/xyrYhO4kCw7cdZp
ORCvWi/XDNbiAFsYlvVnFwG2CqBBaL3NlcLZaoA+KvWuNtjpkhqpHhzXGKoX3Ac7hDbvZZzFYolj
DLSgm4cp6lpZmkWiV3oEfnN/iXrghq5K/vZbXCae6vsFpVWciESQhW0sCrCfmDBw103XNHZwDC9B
po5VUI9IjYx5PCxbOOlUX8kUyiPLia4wvcvPW66zYXSsHE7mp2uSv05Uz07qvXfybOK/x0e1uoYG
vEQ1nK5EuNRW63ZsEYpAfuxL96gBDed4JIS3m/QO2HysO01j3AX+U2wNdWaus2YrIygcFuuX2K2S
KceYpVbwmexDizK9JIofEryzDZayLs/b3Lw25LKSN3FOIQzw6bqAKIHxtBpmazigjpUMPUnOm9oM
05OP2QtjW4LdzRgCQstMgPciORlSQm7cSzgBJ/mx9JGlx/pcwYVo9fVVk2hhYldGkuqDPlHyM+2j
AuI9tU0bPXEO7I0Eys+8owC0tYb9WM4t0FwqUaxnETn4DcHrZPtPWfzvjvhZ86zxbMo8TO3aVMJA
mnMdhGvsNj/9j2JiJFjxn0VKltbj4hC7denCCKw3+F8Xf1dJ+NWXz+KJKOb0oyuv/yv75xqkV2rB
rCG4dT25lJ1bOIE4uzJvWyZDaAYlSCMjyRXnwMsjEFsysl12FSL1rt8SjQDldvY5y3keLN6hRYKX
rM6wjKIADTmd+SQPaRElNYxOlVRFvBlV0hrRgcLBk/5S8btCVBy88wf3veq67KE9urS3otFzsBar
BH+j2n0ObidO3QTPC3oKuLkl78tjcM7sdK1sgtXwplVr29K6vkvZELstQq4P1i1PFZkUGpEOBmpq
x9g3vt2l2tdmse0svqVH6FJdYsUzFogs6G6EnfqRAwVWVXNZMffvnC1FxlDensg9kXKhhiDGmcPf
kCrX/6yaZY6K9dpa+Vy738WC6/tUVv0/bWoqhn7zUqjpT01wE9ylAV2nHuSG3GyNOqcmqxUhyPPz
e0vUqO2edWNf75WD42TTFUj+np1KAp5Vy92yXpIGBbRY7kqGf48uBJe9CY4px/OllblCQ8O1Kntx
i/LcRWeFIMue2OdbLihGxvv0e7OlcCw2i8mdWNA3P6e/Pk4QPviBBRSxVTVNN31Uyl3XoNk1p3D9
NYSR1EeEpKPS5y9q7Uj6fHU/DTCYhgX6LnQYV7iijWP9SOwk3YWZk+IXGGDW1LwZjL+0Z9ynAyYw
O5FZHxIS2xD17phAvvPvvCMSaFiu3j5Tx1Ity3tlRWpwvNfrnDjn8uGqxx+IQuNVDY6CWT4bgR6R
+fy7I3PTStrW4uRz4jB1LV6oN3mPdYMsGbF4Ypua4Q+qbtYFbBSLhgGnpHqpVb/+DSrzhEmjbn0u
O2fsXu+vTur/Mx6A+49ilAW4UT5dS0dHe1PzzOrm9DKrGazdIdyv/7BFpEx1XoWJepq4E2UaEXlR
w9eMzOTn1yE5Tf8PK+mQSUuQ70Eir2LmSYJlEK0Dj51JOm20RqNMf0S4uJxnzag8wOuuAF7URWXW
lyqUygrqD53hDE9HPSpmGXzFT7PToL0dr/0aBNsUPO86kdETYzDK3S764r0sAsbcmw/ep8157BD3
Q6BE+nec2rVRpzRCmcy+16pcBc/rrZLATMyA2/dEEWzknJOWpHI0qkTrTtBOOUqvx1kluwohdp3k
WjpMmBfTB0/KcpkpLO+COPhg1OsqJn4PU4IGKOQByYk+wRPMNwmeJw+OdKvlbfIInmsqWQNBO8tD
8exJrVkZ8NFKe0bQ1zTUm6UxkdHkaZoYIaZdftW1pHs4MysOvTacMNj0nsSWblRcEJMn0nUEU7MP
3wkLbIeASXcNS2P62BjDYav/yy4DAn4y1PtvC7mRFm7fOUTxBKEr9BLDRnV8siu4ynP6jgrDUhxj
kRzBCVoMzNl/QcWgnheivM7vbBeP1xa0mVwngfjFbTBO4WZoGhTafpqO7kUftzyem5z+F774nb9F
KQZ7Wml6Kn1R4fh9221Ro0vVmHhohzUVD+LK570/wVASt5+t5V/SPaZFnjF6NovfAEaFqqjfJD7m
uJVhcngJmUAoLYfWOlwdPBbU3VKbfDNFqzTaaddVA03cXYrkhwRsvFo7LAJD4CQreDYD8A3RjN9R
C1Y9xgFUjg9ImcK6slfG4Cmux9+yRBM260clz4eu4GGwvrFjNikrmVjkPg+Tsy5wQ8fPqfu3MoRO
O0D6Lpq0VGEf1hMMwWWDWFiDxN5VzXOFDpfhYRGyefSiLv3nWlXcF8h+AN8GyRMz1nT58ub9pa4Z
MpwFIuYiIl3HOOXtTELkcZ3YeuGMeOd9Xpv5SuLxRlQAybTtV36UpN0i6QMyrHhubOHln6mdQYav
mBAFg8puorScNsfjjUK0xX5+RBKXNFsuHHeKy4aXRlnAyBKMAL6Nol0EoruFnN8PpfV3+MpS+AmE
Y6qIOh2sTAePwdR6hHlkRqYCFopflqOrowUrVZI+EOrf9kMrk+Wd0a6uzEOJ2WuV9COFR+HgWvAT
2kmL7+nrtTK5nFsoINGHufJkh9LemV/nONf1RVYVP4seSTe9gY82VKRgGP/pEmpohkT3NrJ7gJPG
P4DK/Q525VkYeN7RfLusta6bc84AQx3IDVv+w1/uG5lMQFjvVek5QA/05m9Pl5Loxpg936pmSjs8
D4EpUoiX9HBi66SGba4c9t7ycqgKypl9HT457KhrlsRe+72PUjTmHhJJgWpUvFVajTx2l9gvo+XB
X9tW8vcHX2f5KOdxMa/k0MH+Jg2TNpyR8Md7culZvz8KtMVjT+5LvBrCJoVyJr7I2sto2IFrBX5V
86K/1raQqc15emSt9QiipF/bM6ZLGYvrz7Ga1k8T0Q5Dd8mgxGQyfgnAd7TGEcZj+G/64U2bBULy
tVsFwzJRw/oy+P7vjXzqCR9Z/FlG0Oq9TIBr1tHvnoWPbDrIAtVkFyTA6ginBecoj0arIIpWX38U
xiGRyIQWVL4/A1GOCW2OGb2vhlBUhXd8rDyp9Pe6o2/cdPPimgnGCHhDoGNUZIKqmltzey//4eFO
OGOa9FCxz9e9gzO4Nt9iRN7FU/qg/Vs5oPZzfJ3fY5LUzIdWvznlmo7Q4DWUu2eY6V+CEyKPP0Cp
5p/u/kb9xR8KoAQybOBUk0VfjZmQ507DEl8obwRTBnnTJzaKAeecnnB90+4lNZR+1AAJQgy9zgdg
kywrzduQ/dGUQPgPH1yIYxKaGR5gkiSMqj/Jj4+sMq1QCBVxBRXgtgx+/8ax9UIEF8tS3ISIlOau
PUGzNHRudwk1hlwTZyPsSEndZxevQvwN2GNh+TawTYNcVXtkoSK3XnF35oZc8YxcBmuibwPhUZ1T
9nr5eD4zfKsLiUMb+CSoBgKvIanh+WgFx6NiYOZewxtzOiGw1AAyt9kri+V6yrtUpY9FaOP9yFGj
AVdH22lx9rANtQv3vGm+wDRPjKixibdxmZDSxduzPWrXNrkO4Up+4wpg3eam1if2ElTRb3GwoC/X
VYY3XzzsBk3rCYlZBdfMLMOCAbBDu/hk25tsBMrIPodkVdaiJCKhBmvLeNHYVpG8kxpVhMKiOnnF
cZzRicEwqSwom8Qn0ADlmbvMChShOI3G/L/xEtX1AxgTVaIUZZix8W80Ox4CYZTRe6eYD41ujTdC
EDflJ9tP0krZbuNEu390KjCmIpL8aECRpaln8Wr8l4+FpoQqMDbhSIVkK9w/Zl3cDIcQIphSPyjh
0ccXcCVpBSuxubBLbuHVT0DID1R7U43whTXbV239p7/q71RER+7Y5pUBZWjx3fiBJxbRdHQtphFS
3Y7T6YmQvCidN8Rv6lOCjNuiHaYfnOcezmrhl29DmSW1FM6x69rZhLbDivxLFcfctJoofp2jdUV7
ZUMh4/y0BDQN5yGumb9MzpYTgLQUjSuAZB1uxq+7/165knLRsUuq5IMM7Ujj16PZDy/hE49giaFo
t/sm4e84Mvj9Hgy5n86Lwrua542H03ycCAOqKTnoAAO9/5uzt1BlXYDBHFBmbWz1+9RMODsSGqPC
pkSDG6LNlzlAeL7IST0WWIdoWKEu3peM3HbdC/sXz9/o5enIoFFTqQf5nQrSP38o7o3hD0woTkMc
llOkCZz7EDKjRXVmlMN6e1crYjkAe/qY9tz9N49J0ScbvYKqjwKAqcJrt6dX4EjcMX35yGbiAoiM
3d3d/MXAzFHNw9S2BW3uP3cZ+B1z0yYT8cIyCc2cLQEoYysWqyoGutVYn0Z+3+kQVHRZnhWhsHc9
F/NxMYOUiIV8LuN7Es+LZWrv20bN1WUnwyj8/DPCnJ8cMuTCPQiDKave2BzUv/k6h4rDhyR0iBJ5
4KymIVdLYNqL7jJ0VpazIFgXSD3zScbcPrcjwx+Rd/CNPRNfDi7jtGJJnKtvFAkCFBpQOOczIzKI
7l0T/d3QvIro7CECt0ZdvM4bM3TL4wO3Q2j9mkH/e3pNnhe4mH1JaQitGAJKO/26E5lfKsB44AAa
fooP1vlIuChfMd1icChD67yMKt7RSXT7Of8IB7zcMJMo4oDh89l2jZPevJOV4unE+d7eOI/FRePH
NIXMFzU9yHmzGxEXyP3vBwk/C/RPyHoL2BzQqLOD0Y6m7uVXrsyfMmsSLgLc+LN0hcBV/tHaDykX
gvrhmzfH/9FZ1oQtk6XfPVqF0ztGx/ae6Tw8OC16c2tdnvWUvDkuOTj3JqO03rq59vlWdq9ObLC2
26pFiBGzklyvibICQH+tQSnYf0aPlZ49SJN1zvHF/VQMVYa7yBd+cSNQGsdsmSy2B37o5M5W1JU8
1txgQk3z7gj+3ruj4TxvKZtEA3t3v35cx4q4QAFt194wDEuJWu6ChwAm9x5OxlpkU5/oCLhfP6AY
MfOzKBFy3TEgw1gANT0cWBl//QYV8/K5SxU61CuRAA7qG13812Ga9fd4FjVbiwGN0HpO5bMmeVGZ
/0vDNqgTpBrojjzOImPdJnRYqhNceUnE98HdUhm2OO3cDba6mTXQJCy+29dYdXlo8H80DbbXCYGO
0D4H+5e2r49wX+ZSc8UuNdO+ifBD7AW/8qoJyefbKltqbqJCQZ6gtFcxsEXzW85zodgshZQlQvp2
io04Ts8tuKZbiU0+yJHr35TkPr5orJ7uI92+HIfFFLQrjqncMzaIQrdQ7iMMUQnCITxSDvOwakT0
6wl7vqxDImipNgbmFyVv4mRijtwc7mDFbQpMu9Q7PKi5EpJ27d32E7ry9tJB1yGjoxarixKM5rL8
8Rnbh8fqR9PtmyPe5yrhzaabP9YY7qwQy5ykn1fPDVX2gzoLEIs690SIRgHYq5Izd+Ht4L9gzirS
L+86B+pe0U4w+K9zg6Toqr5h9qYKlWPAzUO7EtFSOmlsi4Hi3myCDOxej+W18nU+gBuHEVqnZwhz
K/C36uXp9000TRhyCdh0US0VdRCL04EX5ZWGfHSp85IYCvq+D2VaaXKMBRRzha70O4ZLe78JCK4G
/u/Nl1MVbxAe48Ipj/8OxZTefp/hSFp404SsfBa87Y295Ag7R/VRt3cOIytwBsqym6wPvtejibn2
bPJS6f/4t2dA2MHtVYk/DPkLmXF3ju/JOMvrLc/SAiETjFMTeIFiHTbATY7sURce1nsiQA6leDQb
GGhSgoc2Pkga4jC6gYMlJH8xkhrtovskk92TUJPeC7g3i7lPtAXl9g3kpbt18Qy2192QXorlf5MV
CvOgMgklIzmqCwlSEp8zkEdTL2s+FY+kvitGPhTOXCx0YHs2tr8WOXd0OgM5nMp0uxVLs7XjhFKZ
0Sxh59YAiJg7xrzqqKdpt8kyhTn9Go6bXp2pxPWiKj5pjybJAD9GBRJXsblbbTCgAY8Om0sf0yvp
6Vhv7pwH2TIMJitwVnsXVNzIlmWvsmK5QZgT61/KyEz5yUhBasv05yfpPfJO9f0OhOMQnIa1+Ptw
EqqD4a2z3p2tfZwlqUO/xVrGORYOQQOIa2lV6zsvKRkIEjXkeUYbZq+ejf8RT0ts67jeiQ4vuKUu
3Z38NIoxv7aWmdgm90daTvKv5Exs0wYl1uKWrRstEo5uZccQBC/VlhFaS7RaskvC5bVcbd9k9CpQ
QwmOXw8n/j+JmDNnqWO20CCAHv6kbkb6qzFdrTGHE/ayj25BwT0mv8t88eLISzblObAi3E2CWqlZ
fSBfY87BNqW2OC53NnbRNBgTyEt5YI4ZN9EJR/rnZjdH7org0Slv0mk6MzAbJMRN0j4QxgppYjAq
XNX0b1rb+qybJ5hdCgEL7G9XMmvE/DKuMQKdqCzUpGCEgvM56oZCSXJo8vfcFPLmue8FcyT1wk84
fEyGkrGrT+gchybk8N7xB1YCkjLSlSNxwHXTlJm639gssp2jWZLu66T5Bi3NwfX+ZqEz2eLUWhlD
8g32E9nptShYa8DinWCylX/Vmzk3GQBj0favZCsF+w4SjB7oOnulo+5UjCp7o92ZHGGcniHFkiuX
2l1Tbsacl7hEjKFzR9IBpM5f56Sh5yd+HbnGXcne9Zd/mlTj1ZK8HhqQcut7LVVfpB3m0bT6wahW
D48upb0vknMJyPuxZPYxGUMw4TWNcEno9CI0gchmfCnvPe4G3oDzB1Slrochz7Ten25b/3uL5oUu
xSfk1oz762HJxkH2uTTXPspV96VEZJ501l9ewIHDzEXQrPdI6cJAdxstEJ5C/Ne7I2aZc9eJ6Pzp
0PAqcoSxZTeVkmfQS8VhbKyVyIvfGFUIavjJpolY4vQhs6FndNTyyb583i/GAxSREHROIM2Rc3qD
erQoMgsJkFAI9UWzFYdZzL9K+/gsC4PWdirPNZgvTpFBGsaoEZQh6UUN78Zo7sEAU35iOJXK7PWy
VBsPH2EOPw1Fdko91TMFuDTLZRUB+zt0Nf3rlYbMPAzy+jTy2Enp9CVF0l1uYhPzP1GQAeBvLDqY
ocM1VcIbbQk4N4uOeT8FOLFZdWJpQk0Ovaiv6VvlgGfa7MNRv8vbtw+ooEgB6PwztqGiCKPE/q9M
J2ZgBkYO3avEAjNbG1vetGLlK1h/LVG/WITsPHkU3TnP5Jd+c50/+LlEkcvmQ6UHasTvKtmn63GV
+mGYOj/7ymaKMKp5HfOqEeUiZRnL7lB8lDJnQEqiovWmSDm/4gxtsErMEX5/pxWugpZ9WkxFTurY
B6WYbesYMTgJIWO+VuamfQ5dN7J7+fWPHzd0gNQlu4Y/3PlroeNe5PK6MMBCTg/zHr1kGuexl1Eq
qy59BcCWrxMUtnFgHOTMkajzQCJ7uwkxc4ZUO344QXOX5EMH3i98EW3T5NTgp3r9+U1EW5GWoFr3
kMx9EmdUX2IihbIySPBIYpBTfysEWjhKZf23NXdff3Khy7hhURck0jmOXttEGl2dtRTY2TfrqODn
LrQkpZT+mf7lXOy34UAfQeA6HKLVLkFA8+Ec5jsHnDU895S2apNIvgTlq9k2VKgB6Z46VGd4jH/W
tAz1RuMjPrxn6uUB05TysCApacQ8QZ1HRiRMXJRDzbI+1CaxMMV/hY4xax6cVP7a1Ll+GFWBtH/c
4bdQ2DDwlmXn+OzURCLlilKYxobPcgto6i8FOTJqmgXE++dkfoiwBhbMkAwwOGHV3cAUlHItzOqW
X1BuqcZ/tAaVxnlRwZRqrDbt1BbsCkPgP0ZM1bjTStkmeYrp2ZuDnkaoyOzZZOvYTgBT/DrhHbCk
RzVsRF1Cj0SamPvzqHeMJqOgKrrKb25lDhqJK96w4CO7289JPThDvfUfiI9xcB8sHDXLQ2wBmzEs
+M1cvNiDSlFHFNBDH3fI+ktlJQ3J7p9MpE1FScZM7VaQ4d36OK7dWID0/GYP1wPs/C1Jh+CrLgyM
I0o4C/N4avpFFUnBBsRu3QlyHAfRghSebRwVxaGlTsXhC2U2S9carnUHcCy9CPqZAwfJEbe66tuR
WWBuI8FeyG43blM1ZNxn0pW/+NYO0er9USzPeGZe2Gh+0yhc6xRHP2X09gnVrNcEYg3Sj3GjYcg0
5gvACsU7//k6NBSBBHV6zFIPiGxqkk/dh9xrg9i8MOO0hiSCw/bcWY81LeU7oyZ0yj3eE+8BCGPX
YJp1DgVVJy6SWEUfS2tuzJ/oFdTj8Bte3+YWpTjNdSfHhFQy6rDUyacazG52dVzg/g18mNZ+P9bo
G7UpsFNLTkm7z821HtlAvlFzrHustW8yMTEB3fhPLgjvnJ1fhAUZuvcPIZ7bdQ9zgdjKzJRjwDYe
iziGfn+XsJMLF5Vo1UX/s3lOjbJ3u/Sh3BP+DcxAGwTSfNR/4SdnhdWdOimJVDYDdkuMca88TkSs
OmqeQIWyeDWt8xHV/PlltopSNR7gL/3ELGzTyiQGjWjFfK/hSKuSzv2bsABTqy2vK40PNqDRHE9X
Ouf1+dTQIj4dvuwCfebl5YVuXnEBzZzk0om83Em8695v5P50Opx73TN+NSryAfjlVfnXSPACFKi4
VW0hk9w/pRULjNlrXPODiGkHwxwH1DB25wKaYkFYtZ9zCJ8Ip8fvzp/WddGAwp3zRDrCmv3d2mD/
HbjhQsuTCUQyRvYsLGSQBVzgqYgcPPiSccUC8Hsfu7YoQq8FSzCSDxMoDpo+eEydFRhJpc9IQ3uk
kA4TD5IYTEB68GT57sH4K1E5L1WgckQm6mt85+vPZZMKuTlAxLemkReO20Svx8HgV1iDVGVYl1Dn
LLRtUGwFttV37syZv32G7I7mmYUyQFt08OjTI6VQedVq00mTalav/vIBshHnsIzh4xidjbWHoGhN
tBMb9ofVzUCmMtp67T1nKszS94YRiyLUooTUJHYoDlL2QOMdb0d0WFQ8nxfK7BIF7sQFYMrzulbo
RiO5W1I/+ptv3LCH+SOydZgvRAcsT730irV8fi5TTyHENyB2hmK88V++dFJVYznUMK8OSC/6AAzU
jWcZRHExnuscPwnHmvrfAYyKUdfEy/fm94PYLVJaYMwRtpffQgugLhEJ4e6jmxQF2aePqBCjQqXJ
oFPUuq1zIqGCuFRGTyASETkU7Yb8P8gmBS0R2jmxRklZkV3sKXNb8FUG8N1RvUwlKpN4ynQ9tfZR
UNq0qEvBz7rPQ4WyAy44/exZI94bLr5nHEnHuaaBuiwXgIOFS4wRVJQZy3LdpQ4HMacyVSSytgn3
LPC5GRJuuFbNOOroZ9Ycr5v5v5De+r3Zw+5zRIfTewcmvo2HuhRQ5+eyz/rIZIa2CqpiSwMWE4EC
h9yglccMBgxLu5XXjkaJNGIO+effc986BkS7b7YLuzHnAXxY4KcgzC112Q52ZVGwgUcrbI7vrbl4
gcDXa6Mlny2s3OFx3oZbfCjJaont3Jw19if4m+dMjdxYXD+7K0KtagdSavRjvMZGR2LaT0exQ5u5
AefXY8QvET/XSuILeeEZ/LpMCwZ9LZoFpQU5rTG4lq6vkKae/90oPH0RqEfCUeb0/g94U+PyekGV
6jvISgOuemNEzZyLJ1CHHdAIFLz/HmFkhvZq4jMd6Wd5Ff5dUVEg4Bs9nYIB2s02pXHEKyk1xdA8
MYfIpAEn9l5MR5QOv8aAl0RMo4B8x2szeVvOezXmEr3b6r5PmL6IriXpc/5eTRULW5VaWFrnBQkp
iib00QAC3r2EWEmrGB1BgaeyheNdoO0eTiWDVh1MbRC/Q9ldQQByXRjdoAAe2mEh3Xn44Jup1xMi
jlW+L3ApM+trJv0/YY0dhpgCQKwDt2D1WGwZtZTrAW+OpcQPhM3YCkACg2RbXeX+VgrqzmAsFDU1
H9W5A30uDMNP9QbRUL9IrQgxym5CaTnOu2iZeA830tWOCKA1gQCHooZIrTjWDPkBxsD+2N9/8fbG
LFQKhl+hTc3LWJsGiHHdX9tdICNbeh422VPXPVmAuHvveFlkbuMRH7J4bHlwTfEKyv/lg9lWNbZf
T8E3uIZNy+8rb3B1+jZLZ+U+YQ9XWM/xhCWbVh3KBDTuh0sloLd2aj+NRUTlqoeBY1SwYwF30lJS
DzMUm2Mlqu+HJIkudCRW0563iWXsxkFmKWle5HFEU+KVt6S8qz9vChltZ1gfsA9KOkZPOHQozePO
fxsQK9CgXGa1EwCeLArNEmL9cx/TKcfDt4KUPueYJAeevP9opAFe1AebvHqxzsNXB9xUBbUv5RX9
warmfSaUFKfofFVUTx/l1/ZIXcwc7Juig7eE5JnBVhWeXrTnF6aVWuvW28uhSQgKXe79Q8Amu0c7
dApavH7OecYsveo/dwC3MjNVo7bU3Y0DbyX+OYhIxK08RK4Tq+vmO3fcFi2VVuOIAPEv2ssL7ihx
Wb5Fg/N9gp0XSSinPKC036pT06DRoTb8fmTI70wdiidzdKeQsLknujAKHHkFnmCiTj80RSG616DQ
9awVdO+A6LAiEBo9hBDDBEb2iofw6Wh6gSNNHy1snSP4u/+LdA+v6B2qM/dk4IEDbnMtkQLHqgXs
Rf/cbs2uZIhAJ/OWHjpFE2pShuBerSINzbdWgMp3QA3D6hhCap3Mjkpuivi+CFD95u41J4MG6eiK
n4dStwGkLAr32SRNmyJpkK+Esp4LcqCxnUMVhQqPuoGc47xOvWE9cAMX2fGDYmuEiCLzEGR6yGbp
V0+G4O/91AGRnXweiMrMkd42kmZXvEwEF1IXZJB1Q9PVIHvEl2IaZZFLhTLkh4p1B1D9OK4k+fsu
qE8014KfEf5Uioqtsv92x5jdBs2aAHzbV46NlqFUUeOpuOrRtRZmHu/YCUiCMDInrWuhXg84NZj9
jqJRFVFwtGOlo3AJLj6Caj3yKWvvmAh0R5Qwu13xrhJruhZppC+b2b7nYhXmhEopyVoUi0jjKdRp
2185SuLStcTT2wE4hXC5PcebAJ7YB+NKBFnnXYpTiE1dviJ9f2OMwED3gIB0byRmMb3Uko16W74k
aY5rC+ekhznFqTkWA9B5xOiaDfDSDiChDuY0EY7tP2vCqTz91bk/WVthY8KlnL9hunxExuyIHVTa
91Hqg6ZEYnWsIwMTv1vCotLj4xDRh+DckPoJIA/lMhQefyLf58OZjrK96E4wS3lb1B8rv1yLCXpq
ulRqNJ6BTm51Epr3BJGnknjwHK6GvEQZ82oOSqm/6bEy3zKIjTYexzbfexibg4MyrWsxXIXPqq6E
uX+QrK9O+3ANWK+0V5MO8ipu/rbXQ4My2hp3C1/wqyRZfFlemeVv5aDAJGWTKWh/sXyKDN5Q6V8d
Kt1C8QnGznRdoqjJSTYxrfEDmpJm0+SA3Ze8wG9xp+2AAQNAi1VT8Ty9d3XeGt2TZivxP8fI8S2R
PVASilHGjiqrrjGoPE2JH4XufPn4wSW2dGsOXkZOwu2A/8CJFjLg422AYAMYB084ZFjR/9J2nO0/
3t7b2fW+An0NjmynnXkJGu+VzTYAxT4XtXHAT+MLsGS8rw/GhqKmJ/4ueaIsM0Xlyp6Tp7yfu5+t
RSV9RHPzcsxgDmKbRbgpv6DbXqNf4HKEnoo4xlgpmqIw61RMHng/Cpk/dz4SbKVeqkL9EJY7iQ1t
LMn+Q0W6Q/Lw7Jr2psP3e8TuzzOechT3W+nORBmKaWYM2AdUlKobYkXF66fK3Ah6c9tGTHlWcK1/
HqVwvDACQ8L6tPqDs5Vs+TRY7sIJJoaZjxBwPKGgvwmSgwwlYPKaoH6JTLaeTp/hqjMa2AvdCsMo
W2yDtEzFd8VVQzG7bJMpKFdkVr01xkFvItNjcW6rjvGculLIY1xqqtZJMJUl+ytmmGbZX4jMR2r4
JqP3cgAoptk+z51iTXb+89sJe/wfCfgsykItoqiZ8DbMUuzdn2c8NImFcmgbcUQn+dQo9b7H1DNf
OJSF7LdpEedgH8UybUdZp2Ban86nLbTGAUY5Zy7016TiahQEWGgSBAEKYp5rCuf6QGsa+fGZa4AV
acZm7K1yIKEIpmviY1ZUaVtkMCiHu0rXI4dY2BGJQ6QPYUJHujLzzlWpqLfpoWb4nYm6Q+XIsnEU
pusxt258mVM7jXgMP6xXKLQ2GRckIB0bYxSqRlhDL1jFfP1EuYSTXGgxJNs+tShUjAHaEzLQy9Fe
2kv5tz2UrFuZFEstZ2jw1ha3B2NySWy5fZa1+g5E0cUaftWNRGkcINcSmkzmBfXUoFw8gCgPnrdC
9DOHwJSnMCyEBaiXN+cudmibUwDwdlZbBTEd/CzMCzEkoNncxFNgI7D3F4Thw/VS77aEVdaloxUf
hTl78X82t2sGgGC3tzIgNpwZ3778bRKjiNmaU8+/V1GtmX7rkpL2Xy19Qhw69EIJHha7FmtWbvEs
bC7mUMKhAoL+c3d8jhT/HgYkEB8ff3Au0EDy+uo3JR7n35g0exTr/PC0RfSjrSURYf1jtx1EB8UP
O0MZMrgYPxAjYMnjG2w4H4VCyAH0bkRrvfGjw7mhzwRdaHnG5SXKqi8mBZvuQQ72E+vxZZmShy93
PkYhnZsG5OpdlfsTpeq5jY5oZE5FFvgj9agVJ2Ae/mGy52IYu3fNYqu0+AStqd5ZOakmh7cBDSaO
xSetSutUEcVE9YF+1aKGx9aYQpY0uf2m5ejXXQUtMZuc6o/MrhY6LctF9sHS2RlAVVUjlglnGgdB
vaRPRBmtkMVNsadaqmRWca3ZMc6IgXhbEP00wbIri+sgaI1YTsXZimU7ETSY80WqRJnxToYeefs2
ePGAf5MwzavF6pbKql0SEqmkgt0eulXojXtG+Qrj6EiBfLOgu99egbvacJdl+xPkXyhowjhkGTuJ
UiF++gLcKk9kG7cOiWE2AbXBm/XeoxV3iWoTi2li6l2tIzepurW70901//8LrJh/EW8wJDQ5ALgq
y6/4chX+gkTT/JDuqyo5qxyplWKmy301rK0rPNGqRolgx61T6S+BvmQacFOZ7XYei60Ls3+thRj6
e3rXanIc0dWSpi5xB1bD9718AHDbnHY6ME4AJ55fSzhAowSSaeTxeX2yU3g1QkJhtqoRl344qDfL
h9QHgMhHpwMOTAVaMsyXzsd7QCQnUe/pl3R8+Kw/uSRh9kDj7afTCG18PXF3q1RKJufz4xYg3VQf
q6wVm9T52pig4birzl45uD01irnWouL53I9plnlOgNa+HzUkSurzEqURLfJ4fF6M/Exwk9gVzcF0
TtA3DMCB1PjbLlKfz2e7o1O1mERO3UdP1ns84+JXI7f93Je71jx+L2fJxfBcyYCe0yXQPRLey64G
MW3dDHTWSQRV6YOyt/M0tbeKTVOt0tVLTK2vFmSnSipRkzcNZFIp1pHxB5PwDOrOdiSkfsE55AjR
RXIf85z8Ye7WGWhmqVDifmKnG9QmYbIQE7U8hh56A2jwV6STY8LwCvzinXVKF3C9JP4F4TZBm0BL
w2uz/Swl60mJ/PQBkux+07iF7uh8V4UdLtBYuOxwU6uBC0WEaguW2TAdOCLy0xiMnJagmgE2fJaL
etGU8ZQ+h0o0wdAyTrtmKcn4BeyUpj+SqrWeEox4rWqdQ5hX68IRLEQRM1nipzNP14GH7aSiTKaP
ual7sV6Mo6v+blgG7Q6XHOdGxNYF9sDu8/HadMYtKg4yri1yiTFtxrmBZipqr/9AWgRbZwW8nGh9
12M/ZVqyCBYUr5matzhAiwt5wK9AXzc2H7TVNn2u0VmerwULUFP3Tc9iXHL0H2QQeZuo3psX+hu1
72273Gpzmtb8FdtatV1FyijUMR0L48kELT44fpIUjHvH61kisusldIXXYlZ/1Gr+ah8Rod8XWvrH
vVNh/0HQlEgaNgxiO/RWFJHodH976IKJDMxC05N9CpmOUnDCzDrLXKHHuWufeNRcNwruWsT/iXwp
dng62nPjz9tOzhn2BOxkVRoC/c9ZW+b+RfEIj0Dxcsz1cAdIEdTihB+phk1M2aV4mJDeLDAxGHD6
SnTFxzLHeW+q58xGbQOFH6i5ZJNXSjfkETw/c7ORuK2VtTEj7xmVuVfOUGNFI0lCUHI7iuK7Fu/7
axHrMtjhPokF4HOrzAdpICKKfhfoX3goiTYBgmtejlxsJ8S1hOAICczQg8LSYe8Q2dETBmFuxqSf
iGlk7D6koNFuHr+yLyqEm271dL2pTQf8t0+ZE1qZIUfBPFoesxpxNu5+T/H0j7YkVHYzxph2INmS
XxilR9lUvD9KKTrVHk/63apgJToNWT3hCWAf/h+WraOPb05XmwOjWstHmH+QY6GKMTueUWfAl3rw
0gqbvpZ2PeDv3hIZhra+m7XODlIeUE3OJO+KSUEd+XIiXq8xWmy2SkGcKcsNsBRUGdo1GKc90T9o
7aFgPtT6t21/R0j3UzjWCpiBn4kNbK3fim1/svCrAEhFyArgPWAl7u2LuRFJAU9RjnNNWjH7v/9t
p+Vex6ubn3aE5bN48RO26tLwcjVkf6lp1eJlzoWljSnlDgwA/GphJgHqRReGo6cVjArz7gDw9X9s
2Rxtx45VF4NFDEY4TvIzErof37WNeNEEpXA9yatuXdBXYYvKKiwB7+nznYRzflamZbPuTGQ6p2ES
03WsHAPyg4eY5mp99MOk+GYh6X0ceti7eD7DgWP+VLGDt8XJZvYe7l7gyovCK7GeOa0ruu9YLjSE
VsU6M6lDuoB4MCHufNOgDR7KtHevLfuloxYzOHodtXF9GUYvDbdryMYRO2aZfbLMuavg0cS5D5FQ
Izyb0XPQjMurcrhOjkFHWvoVejtLOwLy4Fre11xnme0lC3guMmjQo7a/qGdYGSRDhli0ECLta6nI
A4hnfu7azzlqEkke5Zjba4RPC7scoZhdugRMsPSCAbsXLqsXx6SnNAFU2qm0Z4Pqu32fKFzyoWqF
ZoxuNJ4BA6VM5olM5150Jo4Af8bL+7VO+Y2yfkVM+mjI1LtG6/uTIGZPQ9CGt0eJ+Cpo8gFGfWcL
siIqJaMPA2tIpy2tIo8RqPvMhNUYaUK/eL2N8aBiOSbuQjkFjpRjLF9ypZfTkBVQAOA4e1GQLiWV
/OxgzOtmHPV4qnG1gbWgZlgFL4MtQbtTmiEwgyDq1xkK0kccJPnR7/ssLUrpyUgGgfPMxyjyBPsj
oz69YVzu6RKISPXn7ipBTRGmEig0qJlePGr2osWUsROcK7DADEYgCet/KR+VX9MQEW90Zq0FXtGw
JVlmIinKL130giCkgill6G59yky4A/CeOoJ2/39pxRcrtmWZ1N8/SNgXFEnvhmiZAu+eqk9w68Ee
EqGP4OD4OATdijMprKKsGSkMHgfPpm5O74vezL/Vsnn60ySLFadl/MWtLauGGIS3Xf3Fc71mZV83
plaMbw6ds/fa/4rwSYZ3qaw4tAvt1dX0R9Y9pUEsxh89ubAmKFSLCdHW/287XsyAsyY+Ej4gJABZ
EzBjx26gqkqSW3uRwB4n8zV16ixFeezOl64pc4QQCM4oIPy5a2B6yuJ+nnaqPXqqbDME5r8AAWBx
vess5scBQKxGaOnzrCr8zyOjxa9PoR3XGFfL2cYV13n3Jgudatm5e/ePkugcPyOKs/h6vhTeSqIP
7hDUzdgY1OcgyLLLVoh09G9vytEzJEsoHVaM0oLDQpLUhA2WPM6hGVv5fJEvHzZJ1ijroIpn3ctr
14wmu9gVntMeFzA0Ug8E8d0f1dCHMZRgJNde93OB1julVpLq2mlvAX7fIXi4xtOhoU2FRkTMysln
RViirxpzOBgjfpNPQGJUCjC3NucaA6Lp6oZdGYIrbwbpFZPTPrkh3aXU9YGWxopLkO2I57LL0Yff
93Grt6U60Sz9f+oPTAxIPit4HyoDx1eZD4f3DbBlMthnKnVPei8rTjPc+OpTOzUJIXPDkOj1tUpz
CRG7mvvYKbIJImsXxRr9GUHO7PH3/L7TOI264WsDd/56xbjrtandRqC1ylpiYMoh22uYPS2WBcEL
fdkwmAsMVunBM7xJyg2m60XGCegY8n4x+uOTvkt5G9qjGLgi5k5czTsifDYhsXRYgGJJ2ng/HFM7
j8ORqnnAlCU6OuhNRi3SaWiXD6momgjJYuHnQRpoqlffOVxkVHVn3ii2JrAOLDKTTJtGGbVE68hk
ggOSVd4jmn0nMV+Wv/hng5x7xhAku1NDturRhlHAjUoAquaE4ai6MnWAng/m/UuRD6OavOr6F0nv
kgAjupIb7vJEPXYoq5lh3oU3tYb35i9uNxrMDV0oBcm75E3mEeFz/Q+RKVvUYENQUsoZuujxooxo
LdL9V+2JnJ9p378yiCXMR40Jl7zhwKKEcs4mXsS2fTNsu6qO4KmyAnucK7rGD8xCaVMAVxlohaYO
ZJ2HZqlCE29tpEEI0WZYcVSa6EDu9QHoRFYrxhATrDFUnIXpXAXaTiRIS4d5iSHGdv5tlNOvLFCa
4FfrfdpUMXyjyUdSA1OTMoXbGh52oMEsdpbyjz+Q5Aq8ncMYyhEbp2ZWAgkerRCoi3KNjaqjIkZp
oB8AjeTmkVnl96uSVk5nD/Yaf67Klv7SvaneT98I2EwRN9eW0i4GPNXiogSn6w8JBztc7AkBA78P
hkn9D6GskHTEnn1snsmX6ZOdJ739p8YLijII2nfNKJbQ+6R7DUFGzPWfForHlxqIAOzc/1sUt4U7
mhZjrxtKXzcBvFXiMHqTGJksueXSYrk29gfE/jVxVlqCsy1C0h9gP1hB7J8xwo/F+tPigIVVbIU+
xlD8piRP3+AwmGW/g43EjBMYmDXpHv0emeM7xx0QwqaRuk+rk2VPRAuZHHruClLnbJ+PIErgwKwQ
G8S8Wx2XjQjH5E/C5F+ICQQVlh70HBZ0fGgambCkTB3XSMM/YRlxPrQtJRHMJFAh/Qiii7SvMhY7
SX/Zqk5GM3ZjogeLo2E3fcr67bRk7AYfq+EM+Gi3OYUo4K9AQ5YzO4g3Pw/ubFQBL5yo3XjIEsxK
51PT+G/6aBvd6xpVjbEXZlQeBmKornBl9R/H5ECgVe9qJbqaIpvQaiIgTwgLYH7RA/iLv0ugCvpX
ysVpXIBWmxN7J9UbMj5N14/8aXOIZ4/t1ZauEwppLsoQL/x+CC2BHthyD+L+CACbpXSjXkx1b+Da
rY8MF4gIH2rHaMRxAPmbJ/52tmZqorlXSbtA2DfYuARDYEdJbdFsnXBLESAyA7nb0rVUC6+jMwyj
TZ7zYo0ToF77FuouSJy99VOqii2eXW14s8Kb1y0g8p41Ghq2f4Sb1c9DLbsBmjAujP2Eu7/H9g1w
xlZc4a2eyRw8mru/S+Ja7g9vdsOLOp8EbSgBb6anedf5bWzt4VMdviDgHVQMWfGJ6NgZdaQKJkDm
6Hco43+T0oJYWyU+3g1qg1GULAVU8WYeb1mANVhjQTcm4I9I9uzcYXn3mbmJD7LjB22BGcFVwTru
MVWm+dripL26wjicn0FXfNoDCzjqlHJQD7bFHq1Bbix8m+HUyFNCEquzbRCvHNnFawGqsUZHbi0w
UBRdjFCQ1fXv+W4q9PT40/mo0+Z0XVfRGMkZpJKVdbZ5/K/ivm4DbgPiPUeg3qrOO7qCZ5jc5/37
K+KYgC4wusMFft8GDtqs5KiSz1IEf4PDElUCTXNlAIZ7JICSfGwflLpn/iGNuo+2/dm1ggz2P0Zs
iBPyz8Q0VgaxJSX6nDa78ESNGL5+O+xGNZxsFubH20ywYb7QhTzst6N5DSmk3qT7FSMLJ/n5S9BK
ndqfouG4z56ADq9g2H+vKfnA1HH43bzYGtzap1A+K3oRhJgCJIoWC6Myut3ZGaEt/fr7qS5A48CG
0nQJRt6Z1rb7K2hU93s2GfWjsO82dVDCckufF8F4cqiNYK5gOA5RVFCUbHul+BEYrx5z45VstxgS
LWTi9//9yWu5MzViS73hCdESpfCuC0I8hyl7BCotbBQbzUWMkjpdGRYKDpmeopEg16ppC97YSX+m
7k6WgRUDiphzH5qeoPN/4SciXb2KnHqjaXvNDH0QmTC/CbKOCZ0oBmO3bMjMcf2jxwyjRkGRnjM3
lS2MeT7IKCABG7m6tBueEPzuK8jtYGowL/i09Z//SET3jju0tWzXk2S6WNGENeYAXdoKEKtsU8Iq
dUW6fesVr55g0csIak2sSndniG2YkLHXJifvHa+27zKS7/A2cgGVGlemhp5e2EjRINAgY7Jwa8kl
EIAAS+DY5iI6QdqEpl+zWCne6G5DGtdeu5XripvqfLIaJcD4Q8dq9G9/EQpz3dHl3+IAijv6JGiF
V2jeqYjaxJLN/1DAGWRHoxZYUmOihFEaXvGgmKnr6vXURZTJwBOVEpOcrZYK+49iwYZcszgLNel7
RcIsfRuqj8HKERbbqyq48McgqxsYP5eCxgSscK5zVpYtir9UJ8Ol+Vm3pwxvw+W8JhAop9mcsgms
qplm+dbeLXaKrSpWZOyDe/vYPI/Dtnk+0ksxprs9agJgpCaZkEd/O9kWTGcaHS40dI6ZuhAanA4n
mRKPZVWa5PSMbFG2G5sUCDI3Ha2iYP10/x+d+kDvmQyESP0eBFyRmMCWnVa0L1IoPKrNedBKJO4q
IOD9O5mFIAGDKXC9S6hzmHMtrYmgWEHwcDZc2oaqdp0gepWURWuINhOINwRrzxBjqZTqm16vKEpN
nSVkm9sIQhhcHznXRORqZPzCPEQOq/jR/6Y1k12BVP4MYtANnPSwt25/TyqWy7KGSUIbuPiDrajK
Et+XsH9LOmhZVyoE05JF8vV5y41AxnRUDY2Su2jaBHTq6bzBV2UKHLQcbXbDwWVwfQyS0eC/TgT3
JBbUwA8WpugLQsWAMk0CKwn6+A7A3wHpicqPIpcb8hqPOHrfsdnOnf4pMcex9VyqYU+NwQJ8sTmV
f8NqlvZi87zS+hpKykSeA1izrz8qUCWT9Eq/1eW/1GZSJUdoEYzwyqjSvYEuHHNK+NFXZo26hhXc
bUtiLGlIcjb8zmJdIey6pAoOGG4Y9YniCMEERv/+9rCEyoU2cNsAdbO6wYoDQmqjXqNWGiGWlgod
/9URQldGAsQ00ob60s5bCXKDrAAu5hMu/PBk7cvxAcXs+KtrGwJuXONhlaokc2Bp05YhlEH2P51/
Z96lApDN7gjxzRs2/3q6mpK/8yctQh0ENuyJ2L7PbT7l8yxcebLrDiOaeSZOeIt5tBp19xIvoNHh
VnDl9LTLHtBBB7wtYvLqzO7u8MIHogU2Frkrk70jKVSXbQ3WntzTBZokvzhigWj6mkLXjyHL7UQa
MsHFTcpmnB+l/yy7baoz82PvT8w9VK3V5WAx5A5T9VFPWqKTsJdFiZApn3mS76CwWS+UOrTMEcE8
2PGuO0lbhydiepQj0JfhJWd9w9MFZhpUq/LRm5nrjIgVRZUCGIOcFMNbXTsXulztIRo9MLkQvdj5
ZahV32k37ZrLttrNBqIRwnexXvzaNC0D7pbgje+iJoAdw4cyXlM1UUlLpotHKRWHD030LzQQrK1t
7FSPK7fm/DqdA3e22F9ZTVWDZ1IzFZZBlOZi9KVpbQoYlyrXxpnScUpOKLr7v9wEqYQgXBxEnZBU
MFoz2iPcZNZdCQvmgMKanLZPGZoVoa7kbk3b6OvNSVNTi4ztFIVNxesKaBQPkAh4SmKRojizqjqq
holf9+Y+Fjlbuc4IKNsxz2zA0uSABVopzTmGdvBs7mdQ3HGbLf8PLdW5uAlNwRlmT4e9H+IHyQmh
bMjsGbTk752U9flYYitybAwKwN1jfXAsUkeSalz6+2aAHxSzMZ7IZYGaltpAXb2nXuL+TGf/1thj
EWJw3/S604HkgO3w+FL2bKKE1P6p0mFp3+pbNPVraf+bkTHGVkYfu2ZIV+mFRYNWyyW7M22wRISh
Hm3+UtSHhp9TGK1cVGb9QQIwB3D/eYpYLi6wbzpsCBnl+tTix4MllCQG2fZaA8qnWA514d+3ZHmw
cuEfOz9IUhJOSmgxmX+gl2r23z84DyW4tmq7VfJv8HsXUzVA6AmYECAck96qq+TDCByATJcSktti
bBMfg8XbrgcpUo61/fYjO6wncfWbzAmw8XqOa7iWrD4WzMgaYQ5hH9n3c1l2YQnBuYNfraP4uuE3
Uw8qucWc7wqde8D2pELrpIbms5vzcRV/ugVT9EoYRVZ5BNXgIyvLdpZJRyCuZEo9Vw+uhkVWahpI
6EScRCpVuFNwYSGNFcbIFnBL2GK5mb2Cd+UShHQc63J2dC2Bype+6WFM4P6M5aO/L7u16/vyJvYe
7XS8NqtPaba9zp86V0AV6/DIsTlxEZeZXmBxZgC9j8s5GXu6l7KeOFlb4b3NtgklyNywMVB+yyEE
1Z1nDt579+2MCtriNLODbS65QcIgrLbxkbl6qZSfqDa7x3ohYjnp/fD6SZkeZk4xAUBIgaM9Q9Xj
GP1UdMib6/nwOsTaJvV+V4uGQMPyL8czEs9pZ1iOlZPZLD58a0ITnH7DQgJtBI6VnuqjU0pMKXht
2UzH8M1/UsIQRAxEugZ8q1gZEsWpElRTlShVBjhV06NL2IiM68BEtf0KEaH7bDE6kS4o/Ath91Dv
k2xn24KNEfxBECL/NJx4/8/xcsRYAN9N/Q7EMUlnzpPbzdGuHKT88bGoSw+EJpP8cOdMHWE+Hl6X
o/H50jzH8kWCTEJJmDWciAqQhkcQMdcEdor92IVvAwMwCW6r2xiZsmGXPs2ukpfh4jqfNZcgyr6k
8rKZppthzcu4C5VWCwK7+xpG63CTvDZc+RZ6HgQ9A7cnYd91YDX8eEJOSAmQvSq/47JnlInNPl1L
0khEkSzMS4rNJxbn1q62ooeoqH5eZyu4/gx9D4qTiIgzMUdeJ/naBGZTU5HIHt+W18Lpy1+Mp9/5
LyY+qL2ROKeWrt7heL0kjHny+v5zCB7Lq8dyuXKchZA7GNgvN2Al6qNaq43CvG94mOtneWIYojrm
uuBjGTRfMXtoEEcyXbbGHiJuqroE86SZEx1KO/m19ROXPfnsvDC/HkLlnnmb7gUxuIO4hOUCLu8q
naq3JXlgEBrMXY5ZoALyt5Hte7OYKYFAlx9BPnJLrIyWrZAmZv9axK6waQWMmCC+wkiAV9eG6KTt
L2eUnDhAmAz4xQczfk3eE9iJZVmeojZ7ruSw0DyCj2MgofdKLDRQ0gOO/2ifHRTYnV+vkfl5neJU
m1NgjMsW/Wp/Ttvjz34kyY/yDQJvNgn3AElV66JYj57b4y83uxg9fy6uhQIdjlF08hacB0GVD6fK
3AfI6A+2kjayMYj5vgEXsu+EMqfrM6FusKcWyTmgFlBmGxM1SMCV6N1FbzUrWA0/oY/NfvzG5A+a
Vs1yyjAStrciEMuGb3xbb8PYQF+xYzAbZzrtG5pElgNDO6Dv5IvOhe7ySWe3V0zahO49epjT1gMo
9L3Nfa/zb6pk+5XWdL1d1c+chbcnMx/PT4FxYpoYJKHe8xVRnM+P9ZQ9+Bqbr8i6jQO6mH7bslO+
j93/On0E4mZcMNV+SDxhytltYZGZxqf6qNMum0Js9UqbCEQJKgReZP+vln94am78HdivSXw7KgqQ
W0z8lgz/eKY6IZwa26QMFdei7JhPMTIN0qOMMtrGEDduCWHLzMox5AoDeYBUuIGVvqMenZtpabQS
Fr0zWw3AkEm+IATMwMXrnA0aClNoMn7UR/8dShsepSRNUU5yfu78Y6SCLIV4/sZHRclrYbMx8DdO
i+daqRqvr0JtY/45u2eC989VF9CrTyAUUdVz4WmuuBl7WWhFX3KF9CCWpXjNo4osQTH2yRswH01u
Pu3V/QkazAkjUuflTpCh6ptYKkiS53mTLaamuolm6/4oNuS96OvFRfMYnXHQxLiniDB5iVgIigGn
4Ka0+GcUMaPQtgqrbsFWO0JEClobsa6Kt+91Y5mQCJrQ15sf5i4gk/ECwj0ZcM/4DY5WTFVRzl4n
LwiyWgvI3d76+meEWWylxw4JC06MB+GP5w/JX+ad4Lv87mQKQ5EYNG9Zwp+WYmPAP1YEuaqexDQL
ADu5vVM58/ag+vWHYOjAKjTR6cmOTyEkC9f7VxNLMCIzrO1rp4+pgjB+zKGQc9b6iECXUGwPOBBi
j4fztwWrlCJuXfezatTnkChiWvNyJuakvLKHO4vjPg/ztRDpwZJnlfVgXaAHIX4ON+cU5pAqluHJ
d7pst3BXA2OHyTG9MvIPvj5pJr4EJFss3mR2Ou5Xew0m5V4vHSi3ODpI2tSz0fpxKSsD5tFuf5aU
KzNcVy7Lv1Jh7IeoknIXXAq6Dd2CDPIPKWF+lqmeT0GyzPpEeMrZ1whZe1FZrFqTbJHSEFFjU95+
VrC61wg2GxwPchuaSTcB1wL6Kc28lUyAssu4yMLc4ndWs4zJVhEnh8T1hyzY+tHf5PxMiecwWU5w
x3a5yqz/EtMDi2w9uyAMH6vABL4qsQs8k2soGH+pIO2+OnIPJAFk/rVFtLedbQT/4LMfaW8I80oT
0UnUrs6gnLtgS0sljQtaoYJcT3YbcG66qS5tZAvJ3wA6tTUd0cI/ZDAvHzSZL3nsY4nRQZT9nqNR
13ZoJNXfC2d3khBBhFe9XOiQtTjwSiMO1vGeQhaufEYrFLLUkXmZTihfiQtclnhSnsMGFhgF7nqz
bSaEw5vN7oIuDIvLc+j0Un6tIx0QuJu9Xc57Ivh5oo/QE6nVeiDO6WJ1LDJ7RRXL8EeQcLD/lH0Z
vcEOa5PlM6biTvgy9CJlsPNi9LHKB7mWnPqCl8mY8fnhCNBi2Tcv4ncQsM9Tp/N7p1hHwvBlQrMj
5miS1ddlvRN9ZAPbCSPVbTeG6eI4gh3mWTF8pZTvNx8ejyBAPsx/esklBSJQKoKEe26CQKEVdhtA
OPHffLPGito+FQqaZxZ6IqETq3aAICmLhIkuix6f/+iELennOZ5WTzliEKy1/MlbP099/Qx8trms
AKcI3OnECJOZgyA9ndGs999aGGMLk4lCPUueKL5pg6dO36i7IaIEecFAf8kGiKVE++7OoKsgoNPH
upVCPjgahThtkpWBT6nP4ewwVXwy2RjVNwfmXSWWV9FD45/SabVp1Kpr1qiOUpB3zq7pw0DGlyFD
2tkYUGLqQ+nzvhOFusjgNjFXprGD/0iaq592KO0zMTbivnEuA+07smrkyu15mQOHCqJfeIE21lZG
v5mbWTa0t92bamHUbyPnYyGXO0Qph0Cq3z/5Pm3r8qFqh9LHNg+9V88j7mbG+vG8i3xUqCL3F3lP
j8RNWlz8XSeNqhjbQjMHkCOajMPzt5YOUn+zNqSkwP5+MnbDVoxuL4Ld7R37GGgVMGu9X3Uyr7vA
H8ttQ8kG/5w77WKbW6JRqK6m6dp+LZAjd2PjV7y3dLT9Ew7qC31fx5kaqsDiNyiRSrP/cUmrJZdL
PSvjZAo63knLsHqRtNeeOXLVo/j3jh+vJJMr53And+enNAexvWC1ukuBYL+XvWv7RGa1vi9vmWnQ
UulTMHWqtH97eL8RLHuer107Ajm07gJPu8/WNGsZ/L3m2OSTWpyETCscDpBPK1shtu8TY9XAicnG
3SPQD6AEKkzFloJep1qfu9EHpyZaqVGZOGSNv9dRMi46IlDlG9OruqJCQ8BkGu9lVKgZD5wizTKh
wdmWuIIXqzpj0y+A24S0ZlUk4QoYIIKxeJzm/FIhEy36VNqXTFjX+wukcbqS0nywRVFIyxctDC7E
W+j3Bp2FWSlpcj6GgsApQyzWP2M/xQ3qhCc8URctKkyN/7HuVzc8TC436NlfCopd34H4F82s+R4G
zv69FVCMbczWWuSLZTShnjOGImJLQR/svy6ShBRB+FtwrAPBhAHsNp0SPQ0NpS94hfgK6HEtQioN
SYjm9cMyiLClRIw47iSMO2Nt1ZAd5fTB68CxpglyqcAzKDzq+4ELkB3MSckuk5gPr5HMhLBpctWk
vMIRBqZs9Qr4xYQYz1Gkhyf1+9I6+tOE+mkJN2cMbHDvvx09/bG2jrbxlLRW7yv0DNwmMDPG+6hc
ZdNK2Ikv61bNc3ski6ZDzKhD3zNb9Z8FemuuhrY1Vw5HqDEhumoJFN0xyLg080XOoIE0C7iAmMcH
g86vo74CBJ7gQ3CQAjaWnDc4VU3ibMBJcVqTxWkvU2ZHwL4EyffsG75wFoIkSM9Tq/mVpmTTGpc9
OfUgMrsQ5j7WqzuArEIHmk0tbbRfgUawF+yiBXcPNdhGJMvZMCT0d1sDcDWPQ9OLC44CnuFzNC8n
MFemRwZ5bGHuCs5OdgpE0ArQ56Ng8/JvZ9qrXHlFfW9KDPNF6sM6G05a5QZ7DbAdK5HoQshEpjcl
JgIzZTAhHyakVbfB3ZHB+0u5qzebdnIm2JcPsIhyFWy7BAjOj7Wjm1xX7YaIEiu0GC4P7STkJ9oc
IPH+AmBSUSfJzcO7a4XYIRUpTBs3hEmarIJbH0BjHW/yiGZ3mwbdXx6HWLM6lLaYkcXLmiBVm66V
Lw6+kFQ/dibXCf3PX0KeOng8/J1KMDpPJPY/6kiXEQ2ANsPS0xDzcmG+ZczbbMQNBWUpv2xJcLTS
/FwfCjIFfjG1xliKtWyPIGkpvSfefHfrHqWDiQDp8g0YBH2H+EWN45og81aA8aM2K1P74sFvIJbM
qM9t5NfvNWbc+IBajAvyXGqrqppRhFB2pBLhvU+bnffWvA3awWWfuhq26tbWEjY0fUBE6oJqiQZp
9VsxUicC51LSCDD/s8jcyk5Z25utHpVxaq/yu7WaK5mjidL+ee9JBbS950JzRj1l7tRGRPtVfSH1
K0MIR0c9QnryZkNrkJ4cn1CdLgkk8y4VwEFbV/jTBX+iZdTnvsoYVP2fxSyIVVkheAbYcaYqMMz+
pQerjyuBtnFlqNiMQJSVT9LrkUtbAvy8yDgQb3hXlo47N+9EhwGggg46tiHcFd7CIizX1h+wdbI7
HlO1ijMNMqvuowYQDgN9JGmPCVn3iyWoPdkSTVi9wpdz5+ewlxyWCPq0WFr3QkRXlt/q0ohobl/7
bJeQPKLGnrVkmYFO+t9cJCyYOExetDBqkg6IWKX5r7NcixBe6lvKlBrM6LO3K7IOwFDSgYbVYpa4
bCZI8EFgjE6EnkcQV3e0c/xgLEwvqto8gvBvcyb0DFvUnZUXthmSJxoxkorT73WT4f6cpFJDF7I6
HXRH1z07AoQ2zKlv3udmfAQGZd6TCMEW2MbZK2guJCOYeID21fUyx4jLHCPCDvpXEsZ9jTsJKKu3
/M3RC7bXazT0BPXf7/LGFmStZgiE9BPsspi7/C1BL9hqGfbJeCOZtSpTU68DegHWv3LqvAQsZnD7
HckMbQ77xJAXLf8ySed6o8WiZIiKZ+N2NhC3MPGnIgeAe+ABC4v9dk2HglQRIm53r9C/0g6zwJik
Gps0bipMmXS8agttf4ch2hSxSPmiCJ+f1GhtAWQ5513BhTlYkwr2FBt5BKpeZ2VacWNlXf4GP/ce
ip+ruIyIciBW+f5x8NWM+Aj3wQEbc37qHQEi8ZGZlierX5bsKZsF12orRR6iiKiOguN7aRrqJNS2
sSH/tYOF3qKBwHmyt8DPM0HoTarhf12zmCAaY0vwK0P68ntuAYahLoHE/FHLwzKs2mzNvmWlckLj
vE4KdHLBEsrCp4fiwdXjjbMuqZ3Is2sTatjENzqUAJoMwCV+EERqOerzg5h8JK/MwL93ntPTe0dh
TBNnDj7rS88DMfQlgcS4MRx33qjGfB0Gzwy5K2ddOa3klMUOtDAmMjCnKaXOOBJ7IDJkjTWsBpTi
aJS62+oPuLd61pRTa4F/cpWS66miyNnJ9vQA9gmffoWC2b4t6k+duPU3Nci3jU1JskjLm/MuJAPP
NIuyFiHb8sOWXpbj3CUUTfM07THCE04R/A/wiCiZdsg50bu5T9jjlpLPv/of05kgFLy+a6RKH6MV
J4kWfch0LRK41AGSYMdaW9ZW+UDi5t9cDBTJP2FkxWXY9vMZWsycMNJjOEwlpkPBDYgeIWFGCxnZ
+A8GwnR7w/j6h3VZHfMyxmAwIFHJm4BkiVteHzObBhAqIgAu41lGNJRrvR16OqK4my+9/rhf7U4s
Puvb5IDymUtPzVlM2eXnyj9NgfXgszakP1VTOWCBdko9+x/cl+DvOFz8HbftS1gpJrHkhUcqVA8K
nABHKJzSlt7ICHI/+/nVGIAPhYVyRz3w+BZ5BVZ+eI1r4/pAuUdYlUEwxMF9WmRSCfvxUPcqNO0y
uotBXNraR9U9G/ptkCeGmXh1eBl8CKQna4CZ6Ns7VX3vHsbUce8Ubhijw5wYSuxD8RycjdQe2XAm
4vih9UIaHvUzdmxJLmUaofupBmAO7VuOteEFCjkd3K8WVPxql7PQXPqfNhUvp/JINwBHJD4kuVHF
SXGzt3yeqCdVZ4MbALG0gD8SsxidgmWTPvjLFx1SHVFGEeFQI3T0UyTbG/sqeaQa6agtVXuz+1ff
goI+OCsMUfLrQo+UeeFSNuVnnhoNeGoi+1+om7etoq5cKx42Quix7jYq2XC5TgOyLfW1LUCu510o
vJXT/maY7TYibXOQpprrOwRdXaqb+LsVWgubxTLxffuD/akvT3XlnLDNoih0je4vD+M+cU5NyHIQ
sJdsJeIPH4l/X07wl/5F0tMBDA9LWnADb7ZVMVUwqAYuhpTX50lP+brhHGegmAzL9e4IRA9l/gDj
5zJQlJ17wDU/oQ5DLIDA00nefoaRzeoRL5AlNkQjEky2U2+ZNUnC8o6y9A3Pwm8QM7fly2kq4SGY
DfDEkOnFZF2w8w0VTXLMAENuXVMO3T4NkqYYxqNLoF+IxeVNI7GNJ4AhTvSk9Fa/3rOkszpSy/zm
rqFKY2OxDdqYTa3OXCj2PmYbX98o4NfvYmCUfmDkQFmEhHhVtnMty32INAHMRsySE0INwFTJWm4g
6c4efSxl/R0QJH2RYCTaLJxT4c3rhHW4EARahLAABJg+3EywtFSklNI9dMvRwluSnbZsvg8bnwLd
jNrgVD2h9o3Xw/oUt8wEkCB7HU3Bth4GrszAjdWcVBw0zgM8o3L49x8GHAhtSOMnn3qY2YHcCfPL
WDfgt8XDZVbxoNeAGuPo2FmCyuRXhkSzRjKhuAASNRU5o06aJr5QWxK1+fndMHVZY1y0/QUkd9pv
HtdKTcb8UWYkLTpLY1wi1gUa73sdW2O6uzAU7bFYQfyEN+Ua8stl9IYhKUCOY1WvtWUOU2mWWgfM
P71q/7hwtggm1aSyl+3EKDHWmRqfrioZ70IhvWi6a9/7pFnClkBuBbC2NHEaKMJQTTL1R2yaKnsj
4tj3eq7tDyCwsKHIBz2hdtufTFBqdF77g/8FBJHGdzyJbnsEzGDMLCOJvO4VFcaGrU80ujLtMqHj
Ntgml8QPXjQUcwXfy0LtUQ8D8sCnQfe+lKIL1LSnUbChCDC+x3T5tqD0IUGFTZTyFSXeyc9D2UeP
ciu86d6vahN7P0OR4u/9PxBfswDVJCgOBZZ2xVzIi1+R5d2dN130or7IrOTVjV05mSUPzu5esCSk
1uf/29ie8lB8xFVKivyZk+zVeooObWfXacQquSsXHRvz/IS1ZppaOwUHUTh6FSbOAixS3ZJ6gahn
vTveDqSddTKjCWg5emKkQPrM/8qxLTPScFH8S8jg0OnwUwcNl50dCHtvHZxMMZtaJO4A51BHqvoX
L1/pwVPi7El2+BK38NMtopjD4hmEesJ3qgnt75sFVzeIhgucfKSpf6IJD4SNbpf1RVNBig5BcsGa
BIW/Z5o5Gv94MjpDAToDWQ42fxBqSWEFgZQAHc44KkTjp8/iz3FAkJrcAip4cE1BA70WnBnt0B/J
sLU27SnhFXbUnRi67GreNu1hVE1TENg5E6fbwoN8QboFKxW2YjL9mxye2x8rIFg0uGo9UBnOXlJd
7jh2wGv5NFZ+o0oJehyKr3azHf1FyXospFf8PdNRLn8lEKPp2KQQe6q7+jYv6iV0T5sbIJAyZ9Ch
dfXV1MGpdvunNBEFgUSoC4xvM0mR38oSmBfqvGB8kjcJkzAh92i6OkmwNCOkKXY2ver4CuKQ+vVQ
cW9dJEaPu3qPXYbCd77ErZ+sCZ4tdYKSg+yWiZyJpZAu7gma6k1pZJQk1bjcEA75O7bfnJd+JXqu
nEvMnNfGnuNMO/0UEVSucObaxDa4xcbPWO7KCAwnjMng7eGD7WJSfj5ypeCnBFpEPBdbEWYp7+Qz
M9USMHwkI+iQxbz4Zp0yFaNOZ2K10RGBC9ILXbUnQ4Qj5TAMs2PEOfKp8W42YWsP9jzVdlseJA/S
k7tdLUQdZc+2Awb8VID4m9+mbuyNXRhbbUQ4fQO22tdVAHyuT3+iTNzbXELmOkxeqDZaysOJJv0H
ExB/9/ts1l4EzQfPIlK32mwzQlJapIzB9/1Q6aF2TRNAvu+bU+qmHPmdeZN6VIHU5khQehP4NRfj
nXdKLTwi/1LloonybYPL0wZlBRt5uO20YTyq109Y85vLcH4N+wrqHa6+QMOn18YAQUqpowi7KoAM
JbxaAbsnzL28W1+41QoNO4G1efktl3phCCWqSIMAdTDcgQ8EAzSHbi0MlVvh33ZbANh9y18UZHht
ABPIrWnfqcgqlB1h+7T1vFSXc1PnKdPFkrTg0eNt8+hzrXRAsBxJP0io7BgVYtxYRG0peIj/X6OP
YhwFv7SCSm9WBdCNGIAliqKtxJYesVmos/383rexUPAnLaG1QBa8Om9CfJf5zRnF+NedVY740/CV
8W3zqk5K8T5kWXsGN9XoRqDdgRiIm8O51f/mcLXeI5VIB+kLbowqaLHv5qe+qf709dtKgMPRkALQ
I5en4RsNe67wNmVGYHlAPjmZmDDzBjgINDCoaYjHPIpPf3BbgGSoKguGcYDLPgtCFidtcK1edRiQ
C+y2jNG35ydLFmMfOc9l1L7iVtMFUm/OsLO7d1ayz1tqVp/amFjgW7v8c1qJYBjhqTnJRyv5Vlu+
Py8mbveotqBii6eCNjHSqhi7SlJuk4dAHToy3SY6AaoZZKVs8IbOA7Tvez5q3TV0t9dewPC1Axfa
yTJsHb152+xifLUASkuhSyuAcJJN0+cycWgHUyTV9uuy57msGoYxLl6CCMNKj5ZhRNMQYQnZD3zR
fvj7EG4BmpEMsfm0QHd4KqpAdevkJfqCQR6lEXV+2tcB6NbQQgu/gdZQ3uA2fGwE3IrR0xizeRGv
hnyBRJm7J+e2t3VFp65cYgS5rjgJDrv6l7tlcoMLPDObA/SkSOJfUi6WdLPFuzSXl77CQJfpivkE
QyDVl5Tb+gz0yEW6DNd1NagxnZvdAF6uhJMwT/kf57wvbmOXYaocfd09iO0EGkmqtJ5IvBAfZvKr
a71G8V6df/BufiAgCkSZET5dmx5h9b2eOVjfz9GvX2Jbd48acNnBuki0ABCnxZY8CF5D+awv8BSG
WtZjkLxAY6gEWL5hHHWYCfF2xcsJWxU099kEaVZ1Ls05QVAsWRlhc+fIM4jCx2s4Z1JyRvZc2338
69/a6ccnEy4iS3mrF5D0Tql+1lp4vfTdBjOl5z/hSQytAWQKvTVTBPYq13SGY3IMlyoB6A5zo8jR
GY9XwxI0cmBZ66MhdQ1yEXoPrUsQTN5XUPZKFi8rPbYJhg9C8okT8xXdwVoUUooEztYje6wutkED
3UnCc+T+UYnMeDoEq87rrFwOC8SXJlmuYZ+DeFFDCw13LEWGpWgSLjtZhw02qsDfyHr/4tQNNLaw
8BfozR3NKONR0C5O2fQ+YzMMmp9cBu2PGMyvyKT/37HzyGWDXiuhRZtFqOxNehEczxAfm4Xe8azj
+AINnrXaq8xZXjkJL/ZoZrpTGTz9/np9jVpBlaVaQZExSnDmlq0rSEG7e3IdUq+K9xx9KZ4MtkOt
B0KKlGZTqzsV0vkx9WfxeHB3GhPeNu9tcCmycuprbq5ZMm0s+fz5/hTJv04AOqEaAxocrm1vI0fg
MVfHc9pdpawSM8i95k3HEeTR6IJOM/sBV5RgRYaKkjtvTNmBUPWWJsjNJfhaaOIRVSUYXLjsZpKW
d0EHNz3iTy0Zm3fUZh7lk6GVIJSVDesOVjcRTdol/aZLAk1nvETrB6UTGwSn4oOA2XnR7KwbgFBE
hRb07JblJZVVcY07iCQLAyhOZHF/aomwjql9GcUcekeRVUKUs/UaFK8ASJCpBURf1Xhmh/ew6712
Mu10qy+zPdxiT92fg3LqAfPU5ek2QmNEciAiF85Tjm8tVl+k26XUKMIbaHQygS4a/fOd1AXvJEG9
YyxqGmuiS63RGE+3OS1gMUFsICrLZLp+9tQNf3ib9Bm0KdRimWZCx8V+tEJWlb3iS6YIF+/Um6KI
5U5iN6NQ5aNy4xDzKHE+2OZ3bag5xYgAyz0V9QVYFb44wzgJFkxyStFRq11Dvq/xvpfEUh+hQcWx
2KhpMS5zhJF49FdLqg6HK/GKqR4RRn2M4Wo376JuaTMr9FnYVE2Huhe8zzeNhuF05QI6F6n1gYZT
0fMhFlnvFESVqwbkfNgvBYu9qOLlLt+L/c+nhBHoVAVN1QGQ1VgE5zF6Kg/mhibkzAN7hIfVWGRn
JNeDgwK7kWEBHdWB+syXZ4fddzBGiXah/U3jM/Q6pGnHCZk9o/PFv3OGwlHWizQ8ABK3ZT4QeHS0
8fjaxAzJJwKCMhM57NlkwvBvu9f0vfbEzikob9G5uZIHSrIowcjBw1EF1RKxbvQLpKEB1EeZhf39
5GfXreKAnolCZOTVkDWimrcoUDQLLKvRC5EJdS+/gjKtXrgS0oD2Rm5CvGRV1jcT5ziAb2rSW4ye
xZ2OMTfmCsP8G4Qau4DOrzfK25Hqu+0vVNFctZ2EAre2pF0Opgv2aS/4gsvxcgqgZ4ri0lNRe8OG
//iYPEgkaHXd3R4d58ZkBo8aJkKPwGA9NAXcMYhWdNEaicsmkDdeReT09kUZmpRove954kGz/RC1
2P0agMHYb0/JhJPzFQIdcYymR+3RLNF1viWiBkqmHeeQ/CYgn7868iG6JNXg9QBllRdn73mRLsTq
vtXbOF8+X8b+msqnDq+6nVPbZpFHMD9oLELbLhWowvu6N2qCJJF/pgv6NfJdvzlXDkel7V4hDvS1
WQK9RH3gMHhL7f+63WLAIbTQZZz/gzfa8x+JOmEpBGAjRj1UaBfrmL1yWxHCnxw6bY6fJvWIFAE4
XXC5QFNIHJ9IljAiEwAdzuEO30L/iowtT1RMwE73nzCiBR9zVLbKn5iEAuKYSSslvPfKemLdH2l5
VOrtqOoYG86lqWWxAe5sMjTHQJfdfl9MRcwAp6CTNbsQAfo9C1b9bZ5UEZuAZauIFKN40OI4K4BC
quaXdwfyZfrLrnu/9nKr9TeZlSdomfaZX4BaY0GvO993ScNeLcDyMuE25Ortg6En5HzIw4OC0nwG
3bFXOO8J/awMY7vCQTrO3GUlk7bPi0KYb/b+AimIwYURLWy4ZZigsixq8U9RZ+A1GPUPrxEj0XXQ
cqj/TJW45ca8lTigEnZjb3pBIuDnIY0ooHgyOkQRMAEqDDNkIxVjkdSp8mIlQiyrrWqnWJK0R1T1
b4KxVQA48sEcUjBtFi0Kkp/UQfyaTILKFyzzUManIPWu23H9okUdJMEuy0vduH1BHCfIkgF7Uid0
y006y3tPasMUnQxWqY7wqIIImkVK/mkY4Ol+QdFLOfOnxgtm+6Wm8ShjwfH2Jr1O1fK7yRyyLNr9
tZ/gjzq6SJGc5iU4zOJrtln00660ZR7oFKXrCGyfGxltCoHYaEKomRyg1VEBJws82lxaAdqIy4fn
n5rKTg7Yeb8wcM/gbqNH1q4Jz02dY2PAc3smCdc8mv5Iwwmn32Ev16CyzftVOlJ4DixVTwXKjRpn
fAfTx2WSWAAhB6HYzrgu/bD4duZbUbZJd7xj70YvPePMcJqeNj6/jl1/Vb8WxG4MNKDz4WzlrDr6
BLfYkqLloAghWvDCrQaZwTFU4e+4iNbnckYXL95gk3mu2eDHvl/2ugs75oc0c3rGyYli2CGVCTJm
yJ55G0meod/58mypmzeIRVlF4Nfx9nK/oGw++wZXMHTGlBaLVquOnT3tEsLfx1bxU6JIS8TiyXdU
fXJQjRpptYR5QyD8D446Thq8UOonFHJ63y1OsBsFr70GheSNHAlAqxpIWM/LQarRGufOjQi8yd7u
N+2x5SoL7zzyJMK4R/+/83nx7oibAthIf+tiM2wSzv5WF08eG+nF0OkSkHH1wAUYbFjxlUQNjuuj
l/uF7SvZM2G3zxQUl8fDGr6lMa6HEUBjlzku0QDQvEK8J1q2/eXbHTKpuUzVrzf660zqh2/DbELt
T3Rd2X66i/4Lx0oDiuHcm5Xtr9vN9I+YCBZomb4a/eQ0KI2OB4lk1g4tI8lYOGlHi0Dyfl2kSNfH
O1EPZd6CospYClLOvg9uEFYvAqxvb8fvJUCWTB9TYraFLDJOHuiMzCSdtuxTbuPuqOLuot850Ahy
HkrWmFurZ1yVNlhdCSNlUkzkejkvwektvgrHgp2ro5tJ1AzqzFF0sjBobku8VBObIfncjS4E1cz5
GhBXAzJe6hrK83BOETcolHpVH6MzG4hWbIMvXIeMbOG/IRcI3yPLl4Oi5Dm2kyuRrW076OK8V9nn
0qCMH7G6kv/0McDiOpJlauLp3kA5Qqm/8d7v0MxzxpoGs6VwxMVRstVo0suYOjTqsgSCW+6oCzTg
jvVINw+zgXGunEWTAORqwGRKmTFZyDASHrlGrp5QV63+kKeJl5hTnSy0JAfuUEroSVhf04oEaGrQ
1t7173l3tyuJX5L/OmabpHmATDGsFXGICIAlWLYjKHF66WHPkZeepAw6wmx7QX3Ad8CWqhmWJ7CP
Tjfod+c1xihbckOAstO7AEjwr4CiO4E0a/e8kGOwQ9f5kl0iWsnH34aAfQDD1M7Sg/IIo4yVBc3W
gFAuXy4sKqsVl4nSeybsVhUPiVgW22k4/RiWsYQFza5208IGJYZuhTye+AjlqOWS3c/8qT5Afacb
IGOGqtcnv/oTxVmi5q57zpZYpStmtPzyyEcfXJ9dCTD1H15qWS+/I7xGcE+d68evR86fXuhiFjJu
VXs4wtls0ZI5EGpNRVLVZFZWd1/Tz00vycd1c89RG1AZnqLtR/5OuWQ6Z1oVi0azNJQ3IoA9wGNw
oFDy05O93kPE4I72jc5tiO/s4JJ8r+PAK2FIi3c9Wt9RqPtT/w5dJHqXaam8CYd2/5H48WJGL84k
bIMEPtGE0JyxUXFewAU1cYvWZsAVtwSwosIJXR0NrBUn2lBzAtG50/1OlVF+PemWikf69fLUW6Q+
QSs70KV7RkzNVf1j4ah0+OnaLlUrXLjICPv5AnFBqZnbz0iv+C2KYFLSEtZTaQRFe3ypT2BDxENu
5vWrInpU3Sx3aVo2uMU1/iErLkcFp0AuepFo/EanCw/xO6jSrclNlYJUiySITDvO0PHvtKM8a/0t
YQtYyi0sWMbc9Jb56yxrzLzOjR2fRsBJfQymbB4Zd6SpG38hYHhNKimBJir2XAMtUBO0AUK+1FpY
7ChVwvPy0EFjX9u3/Z5cLJFpQDksQ/rnRIro/ENAQ+KeDcl3Oc8p4Nf7aM44nW+6oeg3fKmlTLtb
YeXTP8Ys2yyw8MqrZj/ITM3S76LOcRZ8invy8uQr2ED+eIw3PI7A1AiHp9zxeE3BNu6aw9aF3i6g
iilV1mZxCQkDAGYirC04c+rvQmiWxRnvnGSw/RU/vfJfIqarx27qwRS3I0JdyXsE0RPB0NzVxtei
//Hj0OkVg9vNJiWlHLA+QXp1q2vv4nMr3ZtkgWvFMAg2A9xM60xhEUAL7IukrbMec6CtR92lXmB2
1WVOcIr+OwvCIpCOh62AfER5vnv7Mb1J1psDZUpiOdRvjzTLqi++VXl/626rHBKS7/m+iTHEByag
bTI4FN7MRqTwAteeqUSnQJxAaNmkUjxCKrU/g5rX64/kXoCrTdrMJsdUVRUStHhKuaxRkmf16tFD
TZQVVjxbUu7te81la1c8D4gm7g2WiCV+vhYxQyrkpDPR0FYLoo8LPRsB/AIY3oq5W6x7sk8pa/wj
qdd/lMI03NCcqMYc81M/5+kaS/pfn+Hp+FNoXI0orvNQfJsGEyzdJhtAo9jI9Hn+atYIWQcGDqBG
6jBYWT4w9hyGiiQHA5mGA48Zp/BvH209T+w5aN2SCvI4FrJVshwxsn8cYIUK6QsE/CXpdyu9ospc
ygl4rDIUhmL7ciYBW8vEBJma+uiDgLHbG2slK3suJzmzc3ITHtVhmahZsqKmI43vivy798Axkkdc
WF2+Lx7losxm2QqLgZ80oGg3Rzuv4rkoxMgDfhtQPKP5uc0BuE8MviRAzfshGm780tx0Zs9C7/CQ
RP8SxPlQmVjdBdBWrxHGVPTL0Fjr0ZH7w/MoJCJUYNGa2cDPsRCPSInD+83mGRclEv2UhX0X1qzm
QW3bhoccoOebYEaOsTdE/kB1C/cgshyci6AMi9KP9gGAienrFTECTLc4nmrKCeIXnrRlaVKL7Qo5
mxwKKd72OPHmW3Izl6AOTgax6n/kcAvNEhcneENX2UUSWVAhQSJA4Ru4AyFJNI50KryZPIVHXOOS
E1nuQ2Soh3fPNhzxCkzFepYurTtS5+JIrjzRaNv8fno/+sI0pz1ghGGm6WujC22qEmkQ09hahA0q
l0bT7VMcNQkjcvETrhM6mPQs8y6OcowGGb6QqjlzL6H+QqB6SOpURc7GfV1lM8VvqQiriUjEPOX5
5sKSdlhyW9jj3KuQ/EsVueVRmJup3iSvXgge6odSqKJhnFVCUjPa+63F7j3lsTCyIyD+jKcYO/2A
ADoFIn+8JxsqEy3JlGg20tK/bXbbuGlHUPAlxBdoN6+2snys3vHDyEdIlvqt1g89CIMmZNjDMx6Q
8xtDV7nYGGzo4KdgrmKlF9622ZSnAK5mh7npXOyNLCobAuQo/Mzm3AZ3sDXNWWdwQMuQh32VbTds
VZY/GLBIMt+InPKZf7GX6T07ILPSMIfj3chohIwD2acBSEUBKGU2wEMqReXjILLGZnTIOj9wmuKl
CZd/PK6Ygw4zSUpIZsw0r/ycZ8lpBZ6R0+SXJHDfhLwbDPecgo9urh0h/gDCOX3AueeiMQ+qbQWO
s8OsbPZ2w+5PVzMyf0k0YmQQz0wJ5mKlkDT4wKpbZmnyaHdWTgqpYz54walRIWS+ycS/rjb2icFq
gFyVM5QSHGfl5vV/pJQAPJR+PKKCXUNs+Pn5Z4zBLmNaruLO0e+1z6vo4LLxReK/DJmxlqyrTJfC
4QCUXj+3GbfAwYjGpsRGbC+Hb2/zJkm0oXswtFkCh2F5Umji2Kk95GaOXjerR4glHDwxAw6RypqH
bnHOapDigfQGfbJ+7rrJVU/chCxO3Bp+xmnrx0FmM8H3FIFH+ZWYXxKXfouPXUo5rFWqFbq1k9lC
11N0hNTiqGdwQAuwpO8XRdOiWMRz5bXNYv+4wxNU4iActGtmNXPD5W0bnyetmqtG0Dr2WzqiF50R
zsVBCAw+LCr//TDA2L/qjUPRNhbsUiBuMS8OJ1b9OZaat1yhLjIdsZDav2yMBP9sXNOu/vsZrKhi
qEfmPitBNht/lb832ffGm9wZACmDFEnbQgmPVrSEOUZfGRLvoJFGjxW2HXUsATT4rMgEYq1wVqao
5JFNlhyqQuhLqMb+xj0g6CE9OifdvQGsKbisbJu9ZvrqzKjES1gBDdnw/WqbRHH7HD98azPULako
f75o8URkjB0/8yCamCekMO5yZGsUU499pZnqn7ui16aFW9AUzBecTRkSkaLZ31zeWh0TGYHSEfan
ifre3TM+I9QrXYSIcGKsYTUMs2UdwGl8eElXEoHt/ZrG9hH4+jFJKjSxGU+gXalKrc1uniotIxcM
uJbSUpp9SdBJWA/BLP2aroXHCwvtwk2G8iGA8XO14hPyB/w8ZTJNoMHyWlef+deS8vQPa4M1dfEb
35kj9zR/wEFuTjPyBKfO7u++gwF0gIJPDDRLKfeGwWVJUFD4Tceu/1zhzTOqJPRLP+qYfUORcwS1
jP70f5+vDYUYzLJKNCHQ7qLHcKdRtP7n3qf0H0528r/OIfjEy5nzOIp4qExUVZWfQGRlEFca5zNX
DHIP/5mObtaXEJ7MJjzd+j1GsPWEND/2qU57EGR0ceyThxkuYejb42SEg+LMZxgXMD+KHZZ7+z5j
heIDVM174e0h9K6hVAQnInVgPpS98RK9pAw0/WZNeS9nqN2uUsu3FjLZ22Orn5hYali1EkKum4J+
+H99sEQ8gnOYjoTXIZId7dwam7Am67EKcJI+Dd1TqeM2iNblr/foIVlEEbUJ7uio80O7Izdc5myN
DOeYmMmaN7HJtQoRAV/M3v/Jd9ZyaTLpwheOdMdu36meqLyriDAmMV66tqCrpXFKt+lF5G13tihj
MJiDcLHBHyb9cNdED3VciP8v+N28jR5Y5A2XRwh10VGmUZQ2KTyjAUvC9+4e0R0QbQdLQKtezkYk
MhzUS3ElVdP7uG37WWgWaxxv/IajWof/+obMDzfCQWRgOHlbaD+cfm5Pc/viN8vJnZg5sc+K/JM0
A9nwXct3IzEr2pUNDR0UhjUfzeb7GhDyt4wBNfw5/e1XvNKLEv1SeU/i/O5srq2M+ZVznqs6/UgT
WFE0fc6TDJO38bxwSV8i/alS3hkDAYDqgPyyZWAHk+758YdAEdFIgAkNNxW2kegNryAA9BQcy7rg
eUGqEEg0tlZDmUf0KtJu9COnuZoyd3ehglIUXuGC+1nRc0vSdnL3oDNCb+sUdoQzeEMe1IH3+1nq
27Zv2C2l00VBSN1Edhz7RwajwDf5a69kgl6hYSsR3DLyTd2er+sjmLKcZl6sHTSy8uePbRvM2tiL
7wqptvb+n8i1IYLWyL4yJYCGDtE6kYXBYD5CqJK6m/bHuxgq3/XYgAwVDDFHAQ2xnw/yhD+ZB6Md
pxtVVeYIXo1w3pzrylXekV1ztbsercAy/DpjypeZ8bIjD1ViFI+HFkA7MBYOd69cx4MRIBlIHXzn
mdhb3nEK+k0wMAl9A6LLF3DFCobtGqHUbW1lTdADOQzBTmH6Emno+UumFW7ojdt2k2HuKElG7fuG
7yBAJJUoSkEY15wY3AvgBZijZ4Fi5zjSwGc75uqVCswo9qBgiQv6sE8uzn2hUhnEJa2fWxucvx++
fkDVb/3IWlLHNn09XasBKEWFKaLeuWAM0hrLEiGRz43nCQQCzcbZjPM04nhrSVwnid8bIXHTFwCn
XlinP7lbpJQheYITu5Od/kXIORFEqSqrfGfzMQn9P1L0HO96k8L9KftNw9p+6SZnw5hk4BFBTBpe
kAK4J94b9lgyzqYGlBU3D8F4e08zWjTu06VFKzGmNEWru4Xnh9g4piKPMdmJkRrS8+m/3b54IBpF
n7tPiV/QWq/OBBgHAjfm+RZizxE6sccaeCQfcCTqhLQ5npNK7tiP7A52VoD23RxJAPhuYurKXYIl
b9gzmZcS8QaMB+JyZCvTBpFfZhercxq2Qr1kDIGLkskV0LFPhCPkc/8oH9Il+YrJkvlNjH4NMlaH
oPkOTMnp+a9XqyhS9gf63vYkl7yGULeXaBZzjixtbTiaJv9IK4JBVvtvzLjcWhK34bVWyYw3Y7Ot
fUe9AlsXkRKoqzaBKhpM4hVN7DVlg/OMSRXaFlznfbt8OgzUCrbTT39UeXdAV1KWSJbagw+WnSO/
5G2bGH17+9ng6NJbxosxbM9acvXpZpTQErPjN+TfpRVDxVfIlAvKX+yfqmylqNidWwQuDgXBuZ32
40XTHqwl71DyLKl1OpO55hOlmtxHbPe1j9E5cFTvOPtt7G61cVG4GG7LhvpzuwgyVPuqdVV7dDYS
H+/71kstVf2r0iaPqYOTg5UCxTA1xyZ3hMTBo9gFMM+2AWYHNLQXXlM8GgNodF64MJ7qTHJ4Rx3v
1iyS67L6GcJjS+NT4IHutmARUlDN85ELjoOA9YiH+qc3MpzTF+T4ih8ynAOvKq5N+p9mFPVxPbiB
c7Ym+ljNyz8WBH4C3Cr0QCMpmN9OmSDHo3B4aMgGGE7Rk2GIolY3Y7GIhBWkKt/C87ThDFXwqK6X
ZPVgvtK/VIub0ETtsdOuiG1pf6fasnyRK8Pr8DzxnIJUgW9TaYek18CJCERjpndUqIaPHimQgp6Q
o9ttcSvXJogdo5B4PJnTdRFQyYvXQhDdK5mg/ySgQ6+NmIZXNTjRuAkcTLDcWPzm9t636tfipJcO
+mQaovNSHAhdY25m+1/zLiWYLNA8Ofith52bF4OgU2/GTC9TU9H2zvHM497pC3iVAF66YTxPC14v
qOAusfD02UIV1H1AGxD9YeqYC1/1EMDD8b1PxCXI1bT2pw9zd0BqAR4dTwzgNQLo8glRik6JeI35
3aMr7ItLkhB0GVIM0J9bxNukp9o5pNhZ8axjnojPEIyW4KZqrBC1rDcqKRX/L0SuklcRkjfyhYDF
Sjyt4D9ALokhyrLhEniRbbiSxk1/uHWIoN/sB6rdXLrE++WU34GfaAIw/wG3jHVk922gLK67MDum
QehJ/+YFLVwNHGpnryrCyxSV0AyhOegS9RQ4DbBp73grhOQM7I4DLfz9Ji33jmUbeMvQ2+cT3O2K
+Z+klAucDML94oPJsWnnhaG9ZMCc7Xo+FZNCyQ7DzjKBHjz5tASR0gEU7Xh6mp6eDRfIZQsIdZWX
EsADU6ljfIPD5BOHLeGJ1t9j1+htndcpf4zt6Z4iV5dTLkDgzdWXKGTVM6hjtIT+B/4KG4hS7YlQ
Yo8vWWE1q7+18u3xGwolEN51Hkr+KrJEh7AWCuX2bO0ixc2qRUPAxqySQl/DS4sS9V1ULEV67RI4
BLB3L6XbVV62m2on+gZVpT4CglJLoIjXKNAn8WRHGpCunD0lNoWCksNsiGDNBEX+lWBKwywGP3Uv
4uxml+sQ/g/D5Ii/SQOnFNvS50/9h0b7wYprId2E1wYHruigMbhnz0gtWUejzJETlIklKDR2mPD+
ZpqRtqVfSWF7tTGKgUrDhaPNoO6VTme65r2Gu7QvKjEQTdZuwTBKw4/FXby8+TAfUlQD/eZyTxU2
WjaTTAYN9LKz97K89MOg6L31owbNY6ywui8nQvvnVagQdGYHOy92cQNrb1N3CSGpUYD5ZsezqH9a
Sai7FxCMVZbqcAk75BRCcBemx/zgnKgfWdZDoN0plbpJ3DSUjBR426qwgXXwy8zGdx2vCGSHWAF5
q+Vut9EEZYo5bGJl2pM/u653hurZPTLHT59L83YHslJoW6zYinrmqCHYX56r6TGTCU+yyQ0ehc2l
z/RL9copZ5jeX3M8FWy8jrfzJQA3BoWFBnQTC6/XtDlve4GuhoGvJvlQTcQYoMho7YYWzq1o0UoA
dHIoli/SLdru2n97W6Vp7HSOnkdILt4ZnFmiPuQeusFptJbXlPtmTBr4VZfpBmF+Tt+anic3s7Ev
iWtbOC6F6WkyJN0D+nLzRsZxh4yVn5qGO4sqxTR3tob/rSK/jEEV7eEaoU2dEADH+Jub2Q9YpQya
VdW1scycvIluw96tZ0OuOFF7hWP7YG4ToJn08Bv37zqrdCpb3aDz7uulk1pcXAoz4RZURsjbyFKs
6/Xz31CowYI5FDaK8mnJGUHKl08r3AmtmKH9hhXXAnhERxp9PcimY6bt1xPDh3vZg5aAdissK0DY
VTS6rX+BPItmKsh4A4fyRrE+hFjuUGfCgQOONDZsjZptcn6wMUn2wh1+bZbiEquU0W5H62UqqKlQ
lznEITUWEUnBn5st5T4MaRcQHPivOc8LD/vPL2GbIBBLJiqIzODYKESptiqr1ZaGs/vgrYsZdmxr
9PENCUuuZgmD6S3NrmyTIxi5iNlp41SOEevqy9Bja64yiHKzK71HfQTqDrNHhO+qm1jhVAmMsVsN
o8Z9i6jRdLmiAULzL4J/B55WG9olRGI1597phaoBzQ7IVoZoi95z89Qf6BcQ+vRQBR3y1ZAvaAYT
7pbc8X2DwNK4AEAcwqGvmZ35cQ21Q73g5accp2FhXDei1PabrvK92vx4+DPslYojLXc+uabDSyM7
J0vwFd2iCgcJoc0JCTGt2D8CVr8DloedzdlTKrEx5eNEWR9WjuiuxBKNBLdFftB6WTnvxkWZ3HV2
ZnF5AqkE+C8R6RwiCxH0rubuDYxgCutqv4FQaqALEKYSqtYr8eGscQYIqh6vntoF5vP6bpEgq6FZ
vkuAxvpb6Rr3lDQeh0VWboKth1azHoJvQppixpfDwD4neACiDOWHg3pWs/of9yH8DBisuyU5WQH7
gk73PPlvgNhGED6WdZKaSS8gwDuRKZDEPcf2MbDg/FO4ePrdv2s0GiG4iwlMrPN1x8PqccWezEJ0
7ug7UxMBIzsLKiM1HCZbxFGkwm9ePHXB1MMxEsN9Jrsakhew7k3T9d0VzSHF5Ernbt1kiMmXYBZR
cy1amJWrjlk3Sn659r8D++sifwVMEEf/ZXIwHYbtH1kKHTjLRSN7ZutLMS+DXDEGMA/ROSwYm+Ub
5cXH+Bt07IMeXL1+sQEpOLs3r0TttoUnPOJHmcO2Jxp4sco77cL9P7ghIvEFJPyljBzv+lL/+r26
lX0dm6t+rhNcJXdXU/oHtcVAodHX+Llg4tK7LlFs4jg1sg2/MbYdekofSuytYHfr/ebGh7Y6kWAp
XP3gA3BAkU/F0O9tFSaG8cXgdMWhWe+GQTklfvs00kFiCYo/FsQY+lUvMSPs6SudzePfLIbhYlUd
yFP9cCnsfu7sTvjrhUSLKOvwDu3KWfFdej6CtYGGxni7Xj3dYZLscse+lQ/lVv4fuKjtzi9tFix3
9xYjgBdNCaR0uGLAAHsULgwkWpQIDVowNh9WqfcW2G3ODJE9ZWoONv5KztE3AQti3E1aUZnD7T17
VLdqYEmxBULd/obw7F2Zol/SL4D9vGAAJsltT5Svc8Uut9gwsmEcPKqOcaRMdCkeYqsgztJl+JA0
vPXl1OErXC79CVqjFHBWGfj7tTTz4vBvQMySqp5uURgLqKcVsh2upMas3BSrf8eMIHlunltKSa0E
OigBbHkelNKxwkL8zAyCBHIcivahj30KU7su14hn8xO2yaCoSptCW2DbBsp16pzn0c77DU/T+MTO
scAvk1PAwa2Ct3U+sBRXXa5oYR9ZOE/VM2tLsrRMWGRMsukkEd8041m9Wx8qJmhe40XHsnNb71yH
t01mMw8SwKSGGQBg5decALlfUnRBwIY8JzTy72wwtGO9eVa1uQyrLXB9LMiSW1kmATvz9Rc0r/Hv
PPZHM8MOmFfVu/p48jQ685FpfMFOvtIPYDU3/LcHViHTDl7Cu2KcaJIoPJJxlR5mP8mGkQNsVl8T
Pjwqfd/fqv7Jjnh/8qzSqIz5qUnCnUiQ6+KSfGZEriJqqQjPgsTny+dUlgV1JtA1OSA8yGLsmyd9
yI5zTEfSKOHSQxH7vkR5SjShjnlb1LX+jxIor7eRUR4Pdcsb0EsREXkoERGtyPCq65g1bJ0FQZ01
bMG3CW/VMj2Hwlg8tecfWVO/rcq7qup2m1wgrl9fJQ/KWKJ4U3zN27OZM0AoTC/9Qf8OmuI0xoQx
tY9K3sVrn1X/hCDUQRMaCtgrRaeV4Z4UzpjSvr7UHagW7d36JYD+4QCA4ycx0BAGLKQ818zepnhH
AvswGegUTn3zXIf/pHCdR9IgVKs2b7Z5XDxBjPXtlP3Wn+GDkCjjUSlmglEWgopllvXlQPA/7l0q
VyCSgalnrVxXLNz1oMQ1dkwnjqNdgp8ffGVyJcl8fNL/EX7/Ewjvh+7w2wwMdiDgWiXGszPPMlhh
W40Nen5FTgDkFHwhrVb5SM/eLAtjQSYSAx6vnBWZjgwJy2DsFF45brMBwAtzkHWzmMM478Ex+cHa
TAQTTGVnS0NMdXYwMWUUyXiZQtV44EmKSG+6ssSzX9QAzmZYH+92O9JT3TZDhx+qIiZE7JeIi7Jx
L5JcpSXWxvoLqnJHDx4KVjRF0GphXcoZu07qerWuq3HeKvBr7XDAOs6yeIbyPIR6HXR30rF6ykK6
nf4WaL4OWt0HZin6RYphipaUBmriEeQk9ORCG4wL2eExGpPkOmMNbLMDvs5ZnyTRXDdOkR27voUn
fDyuatsokHCsomBCFcW0cvNJOvL/Hfml12sINZdv+c98dLKazWRiPqiQoAmlbu8hGwEoDwLTn1Wr
X2ylxZnSnMszCcPiycZqWLWgF/6MyViSRVkYWdKmOmPIrWZdeEbx0Vw5iOJLSTbocIWIOQaNdC3v
4580kW+lVMT6oJrK1bTl++OqerDpNV2lM9bVECZnR9i7lV2AylHOvaL1aySZTUIFyOz/a9BM+soa
OApFfmJMFxDhEcLoKiSmNTjzvyRVfCzrJmIT29WmYYkG+eLRAA2ViAfAWU3a8P18LBneyj2PAkar
HLo0C0kBX8ODPxnsXPpXgQqiiJex12FVIMnjVdV/tuAJbT3z6RzRND64r9MGywmXfcKNnl08YfrD
Ottj9fA4EcO2qpJphuHtDyTf3AJEI0yxgFKxOtOdLZ4HV9peO2O5qlvc/7JuhXd4whe1jaXtnnz0
4Ith/jGlN7srCEVYzKhr1T9wQfDiT5INZA/Goy1UcS31eKLyfT8TdRY1wj5p1eZFmafHXgaVu8RA
A3oOqe0jjRkhVaDoerxJJkjUwx5wbziDGZZc7Z1234hYjyNnWd9DnmAlXnO6QDdlUQ/bbjTiA0mx
369sS35PQMGydMxFwo6ffoPX8Fc5yyNC46XdS2nY+5rp9I8cdRiVSOaweI7oCcRw3d2UU8iwl+iJ
PVj2RkWlop3qIlYsvGZ3+vNCmLVeKGGdE1bgs3t7VKZ0UIkIxepHizV9HDsRRvX/Kc/Lk2jRVCds
Q5qmIrX1ShDUM54nRw8jDxZx0loR2Gu0GJYbqJD3bDdcmabDDn2jfqE4JSqs/SADXlBLoUxFyKFv
jJOBd6Pc2NC9loCliGqjzrUrC3bN7HnhVXwL/sQ8NM5t5uAX5fUkSB2k9RxQvE+o5vOpyxlhpf+t
r/zZA45Zl1XNRA+RO0U4wMTtNWx4mJ3dOWGBff4+HxUZ9eFr1wVAe+KgI9rwxLtqrZfAsNjlcXqY
tiBz9ZXIds+BuDh5257EWIjtg0Ne5KDDVdUq2ZxlwYKLMfkihyUaGMuCUUoX/TBHjVIArGOirklg
+RXB3tBWAKtXpIEpWgIwOqvxnGT3jzs5YV3Pp0SQ7vrU2UyybK7xZLebgg2Oc0CZcpL/zQCks9Xe
Aa+bLpxYzqkW1j0YypLdiUSTOoA7MS7EssHq4AWHk4o0RM1odZX4EGHjwO8Pn9nQh74LBJIufwVr
9qsmRdgK4GZXB3k20AU1CnApyZdH11SAuNbvh1OwfCE/U+660wyPKsRiAvYOwgOazuI3lPkz2ifi
vJjwXhNvMXUAPfDgLLta3qIfq55yGUz++ZOW5kuZXKtr6XvlFFK9TODUgPbqyCZCdx2RM5TLkHj2
tDGrJFgevUfhDGH4lgeoSX3jSCekJBvpSMPRE5WU+TuItMrS0kK6+kPwv5rPmhHr1N0HmlMVhwps
nheavpPRD4sZr7HF4IwBecZOR4SbfrXDwJUJdbHBudUv/fE4pYZFECxXTpfw6UzzvkoKwt9MGGqJ
WvDb8g8RQer4GVoY5SWup22w/TkF7cMRyeJDgNdWOioxMi9t2hE3tTYDk6LVWqCI7mTXJLP/rGOV
Zl2UXh7NLkPeQKiqYsttqAcaH4jQ28Lnv/OB/anl4iIKIeO4w/jxPdPlILoQn36XRQFXzN3wpqY2
Pg5Kr/1hyCb5msfFhoCoF11wHu4sRGVT4rIs+N7Ys/MYBZ1uuVcVeVwdm1h+kCGcEm4HsjiK3fLX
m0MCWVN4k0V347j0gtCZWpCdhTaLGu/FsA4sYoQ+64vVc3+pTJlb1mu1kPhGj8K9ykfhu2Q/vUQ/
x6Wg0Lt9hLU4Hur9oW31R8n8reyR0Gx81Gn+e0wnuzE88MUuHUy+qSzk3QLpYYSr9r3/ouIV5hjD
4c80aK7OEEYrdZGsEoMO4TjYaOHb4PeBjrOHTpZlO0GiVxg47Vxr9+UwKw9aV4d6ijW290faS66W
4eZ7+l5HkrTeAxNVzw0UoMnYGwRaz1EcunhpLrJHsC1tA0l0TFd0Y4i07rNkqa4Z1Fgndn0YXeE4
rsDGWB9B9QyZ6VZL/CoX9XR6tdxK3fP5sM3lbnkCJaZByr4kmgk0MTk7uHAKwyCkoUnVC8iXiJEG
fTwS+Hz2yyevweIGmEVq3rPrQS+Yojt0Cl9QJgD6AcHU3EsNkRFM+dUEdQCl6a0duwpcwl4ADQS1
TbjJSZreF8tyHroua7NHEcw8+4eD3AQVmR4XE79ZEqdBBwP5yqE1Yc2Ltsdscj48y3/tsIcXMl5K
BFMnD19cjBRRdEtAsnOeINKqFMOpFBwOuONoEnYxwQdEIkAi82gqAp3syyEd82dodlhdd1UEvMFw
2RhxAhIkrFlbXKrOcAT6P2q2Kr0HWlPrhpe1/tuAgzJM0XSdmQ0TzNy5usAWKUSFi6VSWFKe8EAB
qHIn28djpWuJkAxYcWc/Wfncncu+0i3ZwganfFzLbQ5nF0sCFSq+zJfPc6cGoB59jPT/j4N5956b
cjTbYU5Nmxl7vOhoy2aVANW8z3XztUHgppdHr4HF8I12RuRKiNfCqKG/quT7Dz8xAygj4KnrNysO
9tE2kTP3avvbBruXO6echuCrK4dHfHRmDcfYL7Qx7wWF6S19HeWFBHLLhZHTfwq/c8ys/ze0zDql
1SDpE/gXSewthSUvpzEbZOKmOcZNgUmLRyz/KMuVLi/30RhCxaLx4Jp2wps4zuc834Nxb0ciA9K1
GLY+qkmG/WQIF/+3hIQG2sFT5RbA14qKTGGt22bdfJIJpIKAjgYaIMHYcXmNNxL4X+o7fBM/y9FD
GHtPJBZs1WeG/PncdBpuNqu07ZxJI3uUZaAqNgnMnhtAlMgryWdtqBf7WDZbUr4qchpH4tJzF0o4
TzLMRJ2lGrgvtvWlCEosjQabej7m7tqEAnYzRKxgOwmIwDCIi5JW5YkaF23BZhrSJYmJ/QTzTLhk
yZojq/nAu+yza4LLC/hTxAPRKdi3OB5aClddC3m2rpVZSRzS4ieycHaRc1Fo2+Sal+fEurpDy46I
cQIvFxO3BaZvcgtfC63MSu1EoKaHnlPla0bz2ntJ0WczJprQfoy8IJktFXtqH2XQmU8gbht+hNco
aeseMg25GHviUU1NliR/LFUHfkzL2adOYJorEZNK2wz7hHl7IdjqsU9XlC8V57YbxGBPB8P5gwo0
8xD3rDdXDarBuCd/dpBxBvD7UCjU87C2xcvaHeYFerJ7GKOt28NwPvJhhiYMHZJ+AJY8LWHF51oR
gOewwYxWd00ZV5x61AfkhVMt+nbVCZtjLBXXuE6nMxrYDV2jlmj7qoiFaHGJnoMbiyBynplQGXzr
ApYx9mBrUlxTK/vAUaEYYBFO7qmMSCtUaZcbDuZNUVdpwvUlgy1fqMLMJjhk1znEYF9ExSUnaCrN
zSyo/w2KD/LrtxA8izdrV7v1JVY+V3D8OEhPz1D/sXoSTbUrYokQ3Ggmka6CPw46A4bFGIUs9GT3
C1VcLBon1Ym+AuDYC2ehPbTp4kAksrhwe7Yln8YbN0nPM+UdbjPxTIGwI/88HWz7kZTUALwn/AK5
qIYpu15TxWHrquBvFxXzbRmbnqlF6eq4BH52VSeaONqYvzViqgT/1V+jPtUIW5Oc6PG7qnnInsC8
9DT5pb67V0pL7Jihd5afquHRvKKH1rwsHl4AaG60mVuDE+vVQlYiKVECL2byebwre3fAIk5sw7Vr
7jGqKHrw4FvpC+/PnP+l5yd/+VId1R6PiabOVKr15cY1OUp53x6AL5mdEqGsvkoNhBIQxrDf+yeo
LXTH7ktkajLjYmqDturHmD/Q6iJrUhQ340L4KxNC25XzluwcOAPFM5Q8DZzaW1Kn6+SGB7sM+juD
f80jYZSI38UH3RDGSlcZtk20IAAkoOA55oZVz5qOOgrjg4LyxrB00qRlKxAyRxk/vJbEiNQ2BR7r
RZ7QVMsZkL/mwIJ+aSs+ieofgABXo+m3yx97D52Oto5XYvMG5UlDrCVXyCWGEeEoTpmZGow7ykPp
ZNcohUJ9x7B9q3H/qGoyVDBraCianfHXLIWr4gZSGBGMNXazmm/49VnjLsd7u9AAXT8GBWbXo8P6
KbXHtdy71hVjHVz9mshHD3wg7NjZQoMMYQqQQguk04Hq61zudYiaaTAGb+1kH0BuJb7vCF6FdNZ5
s3EZOerbyaBe6rmkkttAABGqRv9doFmuw7LfvPG0S/tBRYVQqctQc0gYpuip11WVGEP2p+3iT3fh
jf8CCYaCImKpkhK641kYDPEkMmQDQXNajL+TvT6Je3WgDaEH3dNK/4a1vyXxkMWPeDtfcf2BKZua
4cQ71GVxhY16tDYr5khPVTsmnRikGeMBd2DqoqWG5SC/0Jh19/iUgWuAO1FD7thSJhvD3tgGA3w8
LX3Cx/K6OHNvQh5eW2Wo0NUCbmBtCpLChCqgLYmyCWnLLbV+QGN1390iZNH6RooFAWuSoqOkFKCx
F5r8wsloYcNibBDYSz3hC411D6Kk7oLlKRVGXrLNQKZWjKYHvDr72XA35EOnHFIhRZXJOHgDg2/W
YG+Onq33sILs09YE+v9ZUYAPysLhjSLOMT/zdXjtTSUBAgVN5amjsGC8figfvp86Y0ICOz0IMO+Z
gWc21Kq3K0quithweYO93ZlkOf7JwC7Mn6vEMtu2gwOsXIHF8Pp57eeIfAsKluWG0Wn2N9AXxKQ6
XymN1MnpKHGlCyBd39FBaLL5qLOutXrqvB4aTk2Ki2dekax8141bHiMym/Rxi1MdVAEO3w/n1aCu
xyRPLoeO+3BolvKXHptdfx0rtty+mSqAbfmsUHZ4YK0cXLtqdUdTJUjZA7fzVzeBKKMbc3S4g1su
kzrA2z+wjsETJFq5AjC8rvIEHeHNPHRsoLPyMZxEZxE8/i+Wp4JOTrCVI9NlJVIGpQT48/HqD5ha
BTf2ElsISZHSw2NaTtdN4GB7SAvr1lAn82XcB08xMUbvZfwVAyaWQKrkfbaaiUQkE02G503MZfmq
CwWeHMGnWQh6J9Gzwz3wvDdnOFJ8yixcj2zNwoMTQgVRINbQwiDYYuQK3UlrLZGQqOn/d7ctGzzr
r3f4lsHofh1vC7mOGZVTMcmBqCxzuJVIvA/UhbQ7o9KeSF2EnQy1WRxUCzXMifm/NeyWSoVF+ajJ
FxyVmXM97Is3isfkrgFKHy/Io8J+kDOrkM3sxX0l432lD1cM9z2NUqMN1/VmZWAzCr0+VKKVJJ+7
TKILMIceMDZHr55ZUFnWN8NDIskwtGZBLvBd0WpWTiUyXBAE88byPG5aSHhuYCJ44D/nqk0GUkAq
0hJn0LtxG4yFNvP3WzBRkxustGPMcGP5X+Dyu32SPGpcN6OMHf0Fo5bDvelsl43TITTk5vLGdeum
hZ1H6B0Q/mdpd0VXfgTbYobqZYfrJTMP6dMRDUyDrMt6WY6LFxJWCrt7Jb5Aqpywyrw56e8/9dBK
G74c8O17gCfKhklMdcLocWK9tIp35G5jGBU+naNmdfmryU+SVp6CT29B13icq2A8mV5m7QPblHwy
bF48MqYEeEzHw5Wsy1KhAm+f09WuQTUdoQwim0DZ/ZWXCHJQZSnHkuM4xMqCScJ+yTYJtxOggB8d
IYAnO6XCc3QjcbcPdlptFJij+4yozVh6MFrg1CS/jh63ET2Hx8iwfwRW+qcpBxSpR66dAvZFp4uG
kLwl3YwYXPb0yv1LDa7pJqSE8fgd9vLNtKmSjXq7j7pMzcxsohkn30n2Tdlcgzk57bZlfHc56Qzw
VEAAZknsP/FiMFlNvoxJ8gXEbn2H5EYgmymbugVCkoxv42+FuWT44AXBNUp+DCMd4pyg2dhmxkZp
fzikRRP9Y6ieeale87IoH5p5oMa5gvmMoAAvxlHVFZAQQUDP591vmqtDLlXlPzsoVjXZilIOEWJX
UbTH/+4AhpVZyrjH2/9PpALxKkJHk76qZFFvWkO4v7MBtBdqbxHTrnSkieiy77FL5taQfHj92KuI
epkBk6Bnd/th3beEclM3Wbi2BOwtymfEc5dB9wgnz1NWdAp/C/UKyIDk8Dc/pBQjQxXVICUhKIn2
BagK4/B/OygHQOBLS7A3+M8EjLOMfupSGeQD9ZXccVlbl73a9YLi24t9n/XqL11YDVk9j9mXXII0
9IxmLdUQ7HnESmYesCpJQiNPfid4KogErSTSqpEhfgqXceesC/+72A122+A0q1xBpoupzzBWqwvB
t8YZQfHyDKgO3RJCRIPa1k2BWWmzQ3V62ZHEqfL12wwXSt/QSpFStWT1WUWI1bYuxe2ChRc3Ll5E
aGqgN7Ie/b7OzwlIQs5AnhXRGKihZyo8phAmLPtS7buRXlYBZc/fA4RuuLF+C2iEuu/DZE3l1J2R
kqubyLwPykQVaSQtoqdSDR2JQ64i/sEzFZ2B/WRGrpe7b1ckCRFn+tUfK33V2/LBrnzArje3xTAl
bHP9xm23gVnVq9rv+YZqDZm6rMMH7S0bJB8K/R9dKnLyBLkehbt0yr8NeRI6J2ZRUgETlp3QZtiw
FPzadl27tYwfMd+pVNX5JfcruTv4DcXKRS3ValR792FVgqsN2fyyGVi4Sl5Rf6eNlaEAr58A6Uv6
P+XG7fdeasblHOInghLzot6lKTHXVCtLKUQyXm528Prwleag0OOBCzR4szQRWo5kEZro/TQWsPfh
d95k0dzxIvfkpSSamPualSY2o4d9BUVmRud/lyBhRF0Frij/T+B0SP+1CEw1M/ixdzUumBFJx8ys
/ZnOIJrJcQOobiuIn2hFVThOPBbaVCCipREK/PHGFuEUoNbZLvy4p9RuXGhxkxpC3jG2JduACPNB
Pf6PwoGaEZqVueGZg7S4l9uX3byA6VV4geWrhGCIhehiGPQ99V02YdYB+1Wp/tY0HSRFct2tZk+6
oV5DqBSosCiS5N9U2VUy2SVn69KFZk2Jw5kT03+VrB2XXipnfQDYnDQ/+20nmqTKJNGJ5HmlXwLM
YzK9hozFPllHOFExQ/ORyjc+m78kEP6pIE3dQMsEdGc+Fnja+RI0lOXG5hkEctqz7fQRXeK9q02H
AeTM1MVep9AgQOzBfEfRlvFElRtOh1cmc/qLuJ6nqSFqlSUpgS8F2opQ1wz4/vv6wbTLANHTibI3
PZdYJURTNtv0Fzsgzau0ovXhRvqt+hKoRR5X2e8nHHNOPaqDBplnyosAZLPTdC3nSKeG03gnKIjp
+DN/9Bii8ON9wPIuLGb2vN1zJDARyGuwWn513nPq9Vv+OvViIv6l7mSNUtYf4T5eH44XJqlSsVDi
QQZAdUfwOOtshzfKuBBQE0/3t7aX1BtWSwatfCZNOW348rGq8UhUoUOAl4zYghxxKTR2YmzecoNr
HhuxNiSpIsOu0hlOADNDaTYQ/RTde88TshbxmoUNp54C6i7mqkSnP2/R6lsQ9YtCjqdu76ljMraD
Muvs/1TXicpdKmD0Pp62EdJCATiGLnXZSGFz+1QtfC5P1oXlWAtE2LwHqPBXcaHB4cE5XQUDmrat
+3O0EbDKjZWxt9XeUYvuyVP93P46YkEfQxuZ6Af6OWCcnbb1PYsr/MjHdNSnGvr6sqfII5wl62Dd
5seL1Tnmiuu2r7U7FyRvq+N+s1IpRQ4INHCvU/r22xafNPf+FqYI74bwRlsfWWzYPou6DBqrTNQP
kSSBgzfz2/cN8iNcvsq8mHXgFfhsjHlpx7k3ZWSecq5zhxEo1ZYOygfSSAiKd0uugz1TFoxVFOKI
ksL+B52i96JAKd47q0tkSsAwlhO90/NgYX5U/BASdUI/BQ0t5Y/URKAbblV51XKsg+BMXD5bdwar
iamhMaT6qrXPEtXOqTtD21eOFvIOGTWegmERFjVrt1/FgztjiCj8hAYb5c4HRLZBCeda+yojnZ+z
nyOxSHFT/CmERJXiZQjCGN9Gm1P5EACGPODDGKw7Zw7L+QtpfCqE97Bx1tGT+wJP0mdcGB/JEb9D
nfFdxTBoB5rvJ/O360rgwl52SUyOWedCDl75yO0QEY/FBEMzAP9uG3WaDYrL9rNaSRXzS0NHhUb5
zl7SEEZDJqQW7wc8SY4q9nlA4XPYt8TzFlt09rdCfsZGKhHAHEix5O+fnlAGb5T61xp7KBGbjSHC
HxS7jXnwhTJQ8PkqS3EiavpptKInHvP4XfaHJYcIYQKDrlWOF7YVq2rYlBFcP/5ThvZehRpIC+z8
GLsMQsuS+tB4kBcJT3O780zzEzgDLwxb7/700o4bdFUdVahN2Fz4SsRt5Uj3PDrDVAcp+Tdhijxh
DszozTzk7yK9UfqfrRlR9xR3dY8+Hlk/DxuuTmRKve+BksPAVS/B7Et1CEJMYx5j78pR1EawEm1E
Sqjd5y9AsnxdM7HoJ4AeZPn1mcojqOXWub6P+SzUp+ovk5KowB6cKLezpth6tf9W9vQeWjAJJITi
AL2i0IP8S6sJCiZDr4RbybEBZCaykx6opiE4F9+fZUDHdbTMTyVkmz59H0Jgfsric//1ThhegP5P
i86x5xLOAmvPB3rqfioyzocOilzsAMHViC5t+wTZ14E5efLHVGzfSM0K8QriPLU6ZIbkrT3VYe5w
S8pSCqyf0wchowXqQYqEMOaCZexrukaxTex4r/D7vKkjW+y9yW/Cn823a5kFNFEcMJzirrxBJZgZ
0e7apGWZrs0n9/N5dWo5Hibsra0JxkHAl+bmk1TZRpA1dmqW5En9CmaGgfuJYuZ78I6gp73kg3vG
+N/Ma/cUDUCsvpWGlrPbFqffxdqc5zt6Rx6lhSN7/YAgWOrf3FVN+xvgwwBJ/6UX/TmAHmcFlLK0
MmqXqWDPPE7OYRSrFhT1/u1SgNxLgyHIXhcYtnMFwdyJ0nqtmldKaT5ZtZ1IpvtG8Y4ImAYxZPZw
bjzt7NvYxHph4WomhrzIVC4PcoWJkjQ55P36Qrik3NmZicAoNZbe/7l9V6YKdWwgfUPDKL30fg2m
xg17tCPcQupa5HtMa/+KlNIwo7jHbu7+6ZvpMO15NRqvw48CveT8Ph7nGQPB5GE9yxJZ8xhqDNhl
K9LVH9nmvntM+nMoxiTLyCcMpmlW/JYHsPuPR3fUoPQPZy4W3PDYCOyN+JQcBs0sCioMCv1B8d9J
G8ZnnTNrAUAdFAHTUBQNL4m7WcgUEMTZBhZP+EIJwX7d2NlhgxKTAlsKR69+I+twIt2VEn6c7RcS
KGJuKB514zEN/GD1wSB3x0pVgqnhS8ZAh6pipalxsCJKyvnZIVsfG+HFoHVM1aYBoqefPBFQZqDJ
uzO8Fa/TLKvpiP5nsVjKx5SoCwAWFUUrsTuXr9b7405+C8EpNrC9C5lZbrJ4543nMMMyCZD1VZnm
VcWMTMlJMzO0GGZYkeQCSQU/v8BAu0Ei4Y1TnV+Q40t/OFgc+81Fj1CQrG8UX+D2MNJv4GdubMMr
ZsDSA8gcGoFgSoKvU1c6nC6A/HXTvTvc8qtKhWBCV+vNlRZsMpCsiJVtSApKhevtolnM0GMJZ3eK
Ya35R5RUGUIb0PhFYKNkuOAn7hKEgktGIZqox9jNIZa6RRTxYmpBt7o6I9dPybvRXK3zefxE7anS
4nPbbozMI6D2vTwXsAyX1zx+nKT2/B5kdKxVqNWHSuN00gnuTJ4zJelWG9ZkgyxwURwGYwoPkRps
slm7/3GE4W3RfyqE4OGCio/I4KUWXUGKlQBRTr/Nn9+C0o0ZBuR4grOhN/67Ci/J5lbe2zzus+mi
bqpA0/FnSR/jlrVTLrxZ1iC7RkGn6v2otSEdWAN2vlVwXJX6pqlQSjdi5pXy3qvOUdoO8Du02BRh
KKOET2K+iyM4/owi25HLCh91vft4jxiL/Gf5Rx+1/z4x34Wi5o15FGPpIFrKB8JrzxvM/lOn3p75
04Hi9/OBMoWqIPp6IfAcr1fnntlAfpqGVyVHXtrjpMFvOogvudwqWPNvXoGl9kaDquv8mIq2brUK
5SLRrCgkFIdzFHxdPGGvhdS0ILds/LsVZxLAaeVD8vE7DjXZuLqu4KRGgU3tqAH/QagZgb0aFMgq
Nad2tImKuSU3cc6b9Z/5DKX4H98ZIrEPwndQUmkV2ZfRDWaPTTmmxws9dX6ugZkVP4vOrzE8n3Q9
OoysQkqtbEb+GElj8sHEC30+P4cMEdtXuI+g89uwvUeZJcG95xDhZ1LGs2aB0OBDXBDvbJzrh2ZG
r8/0L5KmSlxqECalyejuQ8l1GkhUKqH6OWLJD6H+KB47Jsf9WrCUsz0PM3IP8q3Sy3RnIHnk6zRP
bYhCPuqenjSYS/xBw/sWclkdox8lfA1POks2p6ewpNfCHT50XoIK7uaOP5qbs8t5tZF9Am+CMSxT
9n3At7U/NyINYnOpcvf0ECBDqoE00aRdHKDaXn7OTF1sq1pbMlfawlMIH9G2eVXvKTZoP3E3puw0
WpC8XUON9odzJI6OLirY9W5iFNQvjh7LzXrwJxCBHniuOLw4dTK3ZkT74h/tqIEtLXKx3tR6nj44
I3+SMQcfzsMVKc2kIK62kI+H+7385N3A5mKVMqJud8D9cg0EC33CQRLweCtgT1ZgBAEj8QnoSBp9
Ik9rCd0HoafpatGDwn0tQ4iR3YKy4L5CMrkqigS6pDXmmguR3hCh5xgR5NgNstblWzCGNu1J6lCH
mgnvBNArxoanVsmPHek4ZGyK83/WoXz641B90CoLBFiZcfc+jfqZnFbEPfgFDqRlKh6SR9AX2Hhs
A/RP1qJFIV02C6azzWuXvjvIxxOIaCQveegoigkI7AJ9A/Oiq+7qO1uLQ43t4XaS3fbOSy0+Rlz7
9Eusp+beeo8dDG/mAkDsnkUqWuOj3I/idHMzD8pJjoWSO9Qwuu2xij3XCi/jPtdJklzyWAvN0OeO
mKPKd8Md2XHqVE0i0TomA3QJjczl98JooqZFHgZlFsgefr+yBQL2PqzbueCmTIeL9CZZ9vUa7YWG
i22Nst9v7I/zB4y3kIvqMj8buPz43jhm1iU6ru4x1YSTbGnx+gRiSATOu2hBgZxuKQMtN+IRa9cD
WRnY/XinNxYLInuMBQST82jsl9P8phaqCC6t03/ZiCqlpvtpsKoYjkXkVuwo6oyZuJZn9Al7kXAl
yaslxoyf9k9sO+AkfP8Dz7P9cgEB2QhpN4FuBi1lgdOe+J7jt0OJvkGjvgW+ZdYgyQQqC5+OwziB
Ds8BHAbTuQFiuQedq20qo+ZQBJd1qYvwpyWYJ0MvJ+qQ/qpOp91p/o9vgQir80sTOFstY2+8p09N
q2Wl+eUzLYD0npqXDJQIacv8K302wLltgdSNGua6xtK7Y41dfswSEIiHADTockZWqS/a7wcFG3vh
YPLluFWOF7oUInwfx0xKAfBj3SNl7Zf/DTUH7m7IuAQURsivy3/N+Y76ik/HQGO9hYrPKrpxF5Vh
/FZRAyJrtpEBERWAvDZUtVdZekdQYeVXic0H431/Il77vfBksLyItwjEIWgoQ+ZZ+u0Gzqk48roJ
lfLQR0xLiXrbQRt+G8x7dltxOHNVcE7BXZQjLt8mpY18Vj4lpzJdl5x2lBTT8WoZBbbRswmZUPyy
oH/6Rlga+j+Tw3Bvhxk3xY75QtX4hRnfnnsh+KxF2INRSYh5PEkGHH/rRiEDQ7wK5us94sVjHc4O
BZV92VI7mjCxU/jkdRX0G04Lz6S5DArT01KzhrHGe8I9Guoct40ifEZOMrIuzg+kimmI+J0t/Krx
5EKH77G/GwCIAkH2N8KoOVnUinui2HsClN7bEC8Yh72UGnrN3dD3OmQhPXENfxPcLjMMsQX5R9gE
zDijqJZDsD8UR1fADZ5s+zIBiS2AMokeTxphgcU4BogEx3urSgHdJc/y0ghF9t0z9szcoL1h9Hmn
O4t/x4oVgbzoAWz4nIY0uMQfl3hMVuZkcvrvtX7HTTFno6Hg21dUXhYDMbThEJvKn9rGV+RZPjTL
hDfPXU3oJis1JSUWj72KOUYI8XJRLiFAgcssK8HRm7rXM48sTV1thi+HWphYQmrX7jzeLSGlPhC0
wF2rO8QfWlbdMPj+4lxodW2HMLrVB6Exsc7Mv7XoXvozH2J+OMpKbIEuHf5Vi9W7V/MfNejvHGbP
HEXJCeddJvLJNAC185npZzEstRkzlyZ2uVV19srtXuW4g+JTYCbOxDGmaVA1VcFMjkNlK98P5Aki
ElSLDnkG2sSWnqi5sJWV8CZ0fMWmwvLJlArpI4rhG+sy9uC28HSl0P23566/HF75cgRVeD8e2N22
gdiO+BSXyo0l9oxvKd/sdW/+DgYjWURKFk0IlSNxEO/vJQHmXxs+F+iD4YCOkK+BY2SY9Lh6nxUN
LouZNx2MGdlC1Aw1eX9HGgO3BOEcfBEUMvFPpf0vHxVIR3Agba/1jw0F62vCFh9mnkIY+kN69HXb
qYQykhytr00mDuasB/ZtDRcG5ya04gAUxPmOO8odj6aSDeNUFLEQOTBDPNeVtJ1yo/hnQ22UXOxO
K33GItvyyumCYPDk/zaIVoX9xXn5ZrB/+YBCYypuFE52zzmpU9bEw2lgxM6LkIz4vYPXQXw6nwno
LjMLp9lCXwRsT5Q1vqvCsj/fll8nHipWIGbwvZTfPqkhYqW1ZIIGHl+pb3KQ1dEJHXi+7otPD0fi
vWMBK6X/EgHeQmUQtPw1q0KXfzSPuUV++xn53DXJbMpSBXmEw0R3UxpHwna2Hsrx1B8Td+TUW8bm
Gq2ha/u+t1N+O2RGifim0yO+UsK6VEJIksHKurb5uQVlqKh8gsb5uNYlHCC/b5ytLvEMlzvxAUdL
BYn7pHC1UUQGzPxf99+SVR8V0hIQYPGMIQDU0gF6RcmQKX9kT6oVKtOaE4ZEdUlY4CkqkW/jtwx8
lVhg7BHKz7euhEyG6OQLqQr9voGkWa9E2dRw9OmoTp4+eP2GMHzXHgB2k0DRNUKR89BF1jK8TbKZ
VJz9fo7TPjoeKmBPZ2AN481N51dkOiMEdRyoUP/rs79UTuItprB8DSnH/kzSA+LtJsIKsISEzFWQ
NSQMLHhYjlFlCB4Dlr1FAuQ4hOyVNNGZ3pMpO3XgZyAgLbc2htLL1TYVJj5zq1aAbYEUYuPEcU4R
us0D07KUxxWk1LhrjfUeMbsPDiVs83d+mP1w4ftyi9x6+fBiHtwmmTOc2XtSwJWrV0QimvCqxAUk
R5pdPyFZOP7b1PJ5gy51AI/SmYI5T9Kx/AZdfep4E7/8qvK7hPEpzio3ct05exdx1h0y6Jf3AXgP
pfc/imWZJic88eNCwRP3Zs5aI4lK23Fy49jsG6+usptDSFoYxyfTTCtdtxsNjHbXUfn1UCjWMtaX
ORbsaa1E10QDDdZBkL63KYQRwqP1E+RSqX9g6HWlHVvC3mSz/YNPIRnCxGxOo6kOnWy6Q+rYXTvJ
ZeiD8uwdyHIejd90gmFH6tTVbS09VKiDcyhHFB9G5OITa8Y8b1xBAvVBb8H2z4WeL3LDOB1QjdDy
APSJ6zW1aqDCLO3ampuHcwHHEfz4EtUbY1+IL2cOTXJ8Dr6uvxcmnucrlPp6B53CqrLb4Ccwxc+X
SNu6wv7qPAcm3N2K6mNI/yoI7lY3dxHrkkwygxt4iEH3VI08pfWZ7tViDbQHyA9eLbfAUwHJt5Jt
L67KGWWFY/2C65VexGC6SQhrJhL70Ty4QUKsCf10Su0NnWsXkD0Cn+1Kf9ZgGduN5CpVkwIk+PcE
2cpjgQ+4kbcT/oi4cYPFT1ONbO7Ew4F04x6x6cfvQqXSC0YNwi+Q83tQ3KIslCNPOJ7p5bRI4cmX
J5PwCzbi9d5+6FxufckUBHjA6AB49PY2BDbNSFy3+q4kfjL3J5oNJ9bbtGTUrSKAzX1gfoBavUH/
U/p7uQ0Ky42TQDc4Y0HCyE4FPyQ8WxLdki4EVoqeWAMFRlDJ4PzdgBRXps/YmMZadHTohWJtrOad
+CJ4YPdUB4WQCeSGXWprAtUFnIttt7QqTgBlebZvZY7w+gJRoa5enyfLZ0XEt/eAsbuMFH80nOhW
fom00+47aWlzPnXfyqx4GIvoDJ35KEReCuAn9NWr5N3UQwthBDRWUBYqn6krU1sANTRmiD4fwUbe
tHkRbiQDDeSDSoSUcpYwHWtI6xXc3OtYjYkSvi3blE+62MfODa2OMHrKQUY18O8ttZ9Y6DR3KXXK
P1MHFnH7PBp1KKkTS5wNEtinuEaH7lj9h3I59fqbxFmbWN3X6kC9wkzsGHpKiqL0PS7f737wwTwg
6+iSqSB39XtCGITVViQd/P8pYRq/7nUWn2jNf1SQKix3gsNy1O0SwTmtTZIKSioczqxKyMqgfur0
ZDjorUtiA+TrcyUMJUCZzqzZ33k/nqUlP1CSATWdkAsvMLHIOInH+bvtbZMU9x7WwstN+84evpR7
VpdccUjU36RL+g7GSyh25o1Q09Mrdp8YDeSNBAysfzVqQAs35KS+Q6tg46IAfEkhTcdw+1d0azOj
KZPCUNa/kBVoWKFc6ZHEnx3biAa+VC0r2JiDg/9t6XF9s1s/NOYaoQMfQq3PahdniHgJWuZVAYzZ
aQSdC+OBwljc98UYlNm/84DP+g9Zz7t4YUTpyyxB/eb4U5I+ifNGYewqAMuNQnNviTxVOt2wIz4H
liLqBBVFkuwwNjTiiVhH+W2ZG0FxED21/Xf7sXF26IbC49DfGfBTn9GtJI2TtDZy4mr/CkHjSYr/
Ot6axGVkEnNeNz8m9Yvyf/p6so9LCocv8E35hkBWwqPVDiEw6CiDTiKs5Ae6dYrsq0PJn/hL2gHV
BL2nheRqHs4P8pGFD60cxifG4V7HUyC2N4RYpeyMTNwQADNRRk1vOuzqXB0nQpaTew4/9+RtsO2/
49V4h+RDLqGFzr2rgXXvygmfKbWWb3Xu5H460PS7xYwn3WQmZB87AYcy4hmnay3oss2fYpwVcU9S
4i6MlO2O2XL1KP8UZwtHpMukFtbkbk2djHW6tUTJDsvmJnoEgFGnTm5s6zViqNtUhdb6KUhtAkwd
1ktzR0ttQMX3RVaq64vggfu7kbR/lCK8CqGuOc9povow71nsyBOsya3LHAqVCsnbq89j/SQkVUMc
O/ymcrqynSe4BTcqd8A5Goiz64SLGJvSRb482Fi26npRBLE2YJkLMdBLOe6JO4UjNICTncU7jLmp
tI+g3hJH5dYDFq8tR0ow2mkp6Kp9YZl7zawLzUTV0q2geJ0I1MXrr2zP5W3whh6LKEtj2hueuQ03
sMe5NVvBDMacn7WjDGx0KBBQdWmAIqx1axqsWZzJpeK/Ih3NVsHd353B2cmKJg5zasSZKTZiel/b
UoirsGLxN1urdCQIkxRiC6Oz68qd/+ar2iVq8xzceGf/ar9FKOf/ueMJ+P2WRXXYIJ6QcjF2Q67T
tozXhD2+IrrfjNQEesIjCU3VnIQ3a+qD5tb0TBn3odZtvDQ12KvJrxATmgZTxc23wOqfyrvUCEdv
eFCbOjSFFxoO9ipeCSaEPUy3+WiCtKjRxuDV+VLwQFWv7lEymTIeBYy6e0l5vyh8sELMyK9ALY9h
5TYOo7872NbDhniirb/rg7C3mJlA16odgH5Yu3guJvYrmz3jFvDAkRGNx2eaULymn7QYY5qxnijt
HQUkCKEhKj3tkv+XaqR8suIdKkzo7kehzjgxB4mNoT9WyuXD6amkSJst+lBIFzIQVUy0OYdvu+Sr
BuBswhQDo6coJFmtcofnFBxyNTvXSwH0Z8mHCFM7Y+RDpS+WLeyGOIX3rJ5ACzLK0SuB2j03PZ8J
pGTLk71SEjpHmGemsMr8SSEYIp6YaCnXky3X3WiJeyvqltaEzc0HZIhr6BTfra+esplo5vbzTE1l
kLk4SsEuxsmv+DAzmvfs7X35HPyc4WRmHHFR2W6RjdwHkQQ5dLkXlXX8ZTQbxcIwP6/Lo/J0dYz+
9fAyAQELJ18fkFIzssB9diJRhZsqYpUtvYnl2i4vfXGeW2W5zj4yCVV5lpoFpiGL/BSlQYdhILLj
b2ziQvcK9o9LjrNCkZwHdT4kzjLY4e0bY8h3IMMjiZGRzsjjN1gAIeUJK0tpIAE8nodSwBLYk715
zDYNWFSNrnReh6rGtswQQl/WQgMHXoam5CAH8pnx5Q7vanuyU6US6sGmhS7BD0WTF/nMI5g0wGV4
RcXyKYNVy2wsEbe9MVJlAbFJPGTAmhFdk8ff3Z+rfE1b8Y5k7N166guRfcZYw0BiJYbUQfIzpvGP
Botz1r3px8BmtpcrM/QMnLGbpucnMoiK/MyQfnFdpX/k2Ls+vNtIqFTd2iYp61opMJg+lsKgkLe6
ufg6S4545YHNZ+FiFA/GRvyL6XIS4WwVjyQR2mHWZ31FpRfkoMvyASEdX/qdLkks+R5rR3EszUNW
RWpYRLHbA8Jep2oJMM23mWaF+N6FQck0Uh098zhZUc+UmMoMVAF9ecMWJvF4pUQ6lTTBukS7093Q
757WbwOAcaF6+TzvFevNL3UXUSb3pO1A5kGHSsXnqDpJJ1ScNjGtbc+X1UBPY2jgLtlUcY7+gY6r
dR4MxMeVwFuFxOBT9kAYK1EqN+LrhdBj42LBWBwbIDGU+4ip5UjmbRz5NSdamexr4EDVqNezIGJw
QHhc2VEM83VOtDNTJcbl2Dkc0M+UEY8aZMoHnKd7OPu51e/zTNmdkJcY9mO9ea2eS1wHWeWxCEav
5Df+bXYLXAuXplA0PtegbHJ35zV/0vGfSwB8D9h5Df/nUqvvvT3EYFm7VfWdaGiZKnEQT1MVxVzS
0YcUvxLsIQvwMwtIuLya9D7Y7JvkV1WPVVRH2DH4Y3NrZv266cMsWN0GZisxjZDskkSDteW/mZpe
OXqWBqu3wtvo6uVHJaSOEv7smf4CqROyd8nBNgaM6UTUkFFYCcQmI9dMGXdhRsQw/eg3lBrwN+Ow
/hqUVEXuaPdb/7BkeSjftaRELUPARMw2Anu+UL13DCpmMxYcurTewCJ1DFd7DUR0Phl09I06qiEr
+QhCRVcKma0sLNzqAU8faWoiOyhb23e7lGrDUL2rFKfwXAUVVVyme85Fq/iUxRchUquVKJn/K3MU
fsSiUUqfiYX/ZVw0s1oLLCjoihYI7N2S98d6g7ah3zYUnqPAm8IkYYQ8d5+L/Kt8T/bHz1NpeLC+
2J6mOfhxsS8d+Mjq4xSkKhuaSdwHGzj2/UHp9KsSERjURz1qcoYBBLpIgksW7gMdOIHNShGsr85E
uTg027UmGYvQNKXUwZ0ngJPlWk6WIShXs50VJlN2yQBfyuEOmlOYn1Lm8xL3dyzdo2OBxDW9mgkJ
pss9QMbP7Ruy0sqlG4SQXBV2vY6zdyeh6PwHN5REmSDujAsfyUY2MPwGMjJFZ2z5wv/CtYYkV6Qk
b0dF10mkBWX1pJvKiDOHPSIdPM25MpFi9elrxsDpj0xc7B6YE+gDtkUGk/qzNGtPzB4JBjYil6ci
yRyepR+3ySj+ctgzmfxM0ZmV66iYgEGcD9y5CLGOAQJN8nfmhlJtxGBvFsQGTqg7csZiUxZfG6UJ
PgsuEahlKUgbVWoV/nnXXn3nnjc/4oIITL0Av+QR0ly8kZ/0Oo1tVxzGYJWLySpJd5KH6SOwNU+C
GGmFzghdNcRUwpNvCmc2rLsEDZJEWsWScCIgXP/BRY3hNkDNKAyVZ2zCFkOCmJoYNs9DiuokkxuU
oGqGvSPVPutKPdopW78rswPN9Y9jeoj1O+oSBFnXeNfP2kedg4h/I0wR/065myNgT980aEeuWgbv
r+ukPp3QYb47umC8YSJThUlRlkFmztIEWDTB3IR5Y3NM8YVfQzoJbXPdzTq25W2YXxOGaF84AH8P
exQ0tzrtRp0lBEU4an4lyHwWyOeZyRZqTOw0BIoiZjz/g5B2sjUXK5QZZH0HseCg0FxdMJY2TeZs
K2FehjY/OVXedxbjX+3RX+GnA4e5+HSMjBk4/dPB6ydSrDYRpO9VWHt1PNBRmbXesQxTdT4Fb7LK
rQeMhcRP7s5i4jmChP/nd+F6Ku/WtNXUuP9zbL1svS2AUV6iRn+mjSNL6cT1RpTpqPJ/StlpJQhW
1tOZ4j+juy083z/q7810MolDb/dOXxyHcHp2GOlhInLAYk98KwrrPqGOy4a9UXH33ZwZwtZKY0FV
UpHuDE2yM7oQAjD0w/UBkw3QkT4xbjYQhvL8UoQs2D+g7ufl3xtiAyLy0muRuQCr4Y0oGH36QTLY
HrtmhNPPgqPUucAKoE2Zf16UWTICwv3ksBi82/ofcYuDo2VhwnY73+siGWIJg0iIKy+11yhVjA1Q
a0Epwaa20kuZeM71qgl+DfJ2gc9Oz2pJaekcr2Rae3Iwv/7inRce6CFbEDWy7EjLOIZNYaB9+aSr
HTZvOTtuq5kaTWjCq+7vGyfvd0gLXy7RbKENvkdUHc957LqpguASWcMHnD2sMX1mTmDO+bZk3MFV
ov9FeqEBuX+Zkb62dWp7Dmwfzay7i8IkylEbfxjCNcFwb5wWCV+EBwJ63dSa5vY5ERNFlp4Ttrc7
OY/eQ1D+bNxPFoTEr0eTNzF0XG9cpDl9Ya4GeDdPwHcCJh3x6ylC1Ga07pNAAZ2nK1PWegNhkBbh
cgT6kSk8yRvgorB7KuHa2HriSeMltxvLiVizVJTShTecFQF8kzhdmUeKTa1L7oaRc4Xt/AGNsPvL
ErBv6gZiqQ+9w1WNbtLnIPzjxRq+YIGtlqxOC/htqVddhGBVwQhwqyb/RMVpmuMUEpnRstBwy/4l
7iF/OaI7SIpv/QQgO/NLvP2XfHN4Fct1hQVzH5AERjcHmSHK5b7tBzIkxniZX2dhKQGnY0RkQdOY
X9VLLkqdxzJdy7AlQBXof5vPUSo9I0zoO747esISEIOMKT6rOolgzcuVtmmToI0dhYjbxEFF93WU
5HcsF+AQ3MnzNHMEnIxXMHPMniQyEFLqPFuWtHTmbkmNrGUZawRrL1wczTR8oMngvsYjYCiowqnr
xoMhxk4JhL1DACymDJakl03GoPNQ6gpS0C6w4oytAF1XG8J4aJ0nMmfBrmsEUwxGADVK7Npup+lq
EXts7+/rupdmfIClZLxux2U1Gf/541wppjZ1FfBwaBdtDa8Zv6XOz9gnfeVW9zmHPQ861FjUpsOB
Nt/kDWI8Incq8Oc99TBpAp6kPpp9Oj/N5zyi1VQRLRgmjtGrfcTcuG4wmNoHKX63nCjiFYd2Kdv6
igNad1qj6DeIn2Nzf+npwPvjcD/HGW7Cue+AaqcXKq+ghuFvApZqdTr7/WO6mpfPMi38ay83nTN0
w0xqnvDUqDoD0LyVGWDF6gRbVNMyHo5bglI9fjC03tSLAjH6O/NX/CoMELtJU5FyReINfpZmkOE7
5VNJI5iJxIlauPgakLs7S2Nbz+fgzoCBw54W8Jvt8xqySV3dDEArlaQPzs/NYTW9gc5dQ5RHENMN
nKJwFl5h//Ny6fbQtDnCkHlU1csAPG/trrrc86eNf/1Wp99g35iVhWNCxQBR87E/ociRGDm1koza
+eGem7haXVq5FEynA15oSuva1u9+aJAVDOo5wdIHyfiyOjZKT+K+fNVTNepubYsMe0uD7hfIVAXv
uvq/dN2FdLDKVZpCodonPr+TP0DuevUWujXIqag/xOVU84fHlWUhRSVCn709+Kli84gIwRlkh2N7
5KlR5O52Q5wba6b7YIlsYak68HpTNDH9ODfBwDKA6+Sc3zmdJlVmS7Sushvpi1oFYsP9gMu/7ucj
HwKD4br3dvOfx9bu7R3jpYQV2Vp1kMMXvhsB3/0Hc66zNXTcWxUO2ltVtkAPOrMwasCoTMCEqxZq
s3sqxBHJejeBflm+oiXwaDMphKaBnlWXftzFEUee46iHwP7OsuQv2oMi9w6npG6Xix8hvIKgF/XV
5WUmzVprnKnM4aH/E7DfqmxgXgdD/qeYfDiDC4rE370b4gq6vnkPkn5XRYSKQeZ1iGYrLn38AwcW
OBI8e2Q/YmvgUgStr+AuBdSeueddpc2A3cbG3CyZlH4Xqmv9petnfWV4rp8VghS8fIHCccsOD6G+
IMF0W1dHHWPOjGEWXDPZwDvPwgMLJdLwQAYOLjTOmp5TeeY/7KQAbnNJ71czFRUocob7BePKa77D
2Cp5tQhmMQ55/k3Ylb9sjAcTs+Azz8QXenZp7zDknkJxgoEnYUoRJDXPPSH8N+vvaKJaORE0q5iC
Bb3SKiRMqGLFuxHnEG3jNi/dLIurRa2T3t+PPhFb5htUroLI6f3aT912Qlt45E0uBKIkikhcZ6/N
WPNoQxgSk276nEh/U2U+WWm0QZWGTF6bEodoqH2dznA8nQ1ADnSrFCCCEL3xEOFx4oeF2Lk7hDXD
9L2XQjpyWKwP78qlYRrYyBXJrRPaeITiU0yFY3Wup/zab5CaRuBQPAFnuN4aFhsNJCG9wZF/VNOQ
urCWzwejl0g/p9X/zS86k03+4t1UQZYjLD6e4vZ88bf1SqTcYOy6YXM+uK+dHYVh92we7wIDOszI
MILsO0GC1pVVrvHZEvUnshfY1AFuFJwmpFdVd8gLWW4GudtjG+OLW9zhRhUj90on3TZjADXvXXQi
XzGFfL/YLoQX2LGQKzJ+rd1iYiMRoi9WjFeRqLEgy0W5CNfiLcEQ05kTYK5NzCxv+BwxnaqvQy+S
qGBB1NhofaVMRciY3x4v1k4XDZAVG5oXk2o0lzSuYejESpD/tncwvIkz4gaandHNLSl6R+CyBlvT
RhMtrNwPwiDxrriPxpzmzX7u3oLYc+jMmFTLMVGCJvlO597PNFV+5e03P2reQ2dyjwfn2gey5RPY
O1BcORVJw+bvv3e/brFgw2QEdSnHlstULHKmPm2uC6ypwadSModsE0m7j+sP3tpvQ74kfHdfc3Vs
EGHQPD+JMixT3JbH3m/wVTGq9BQN6lF6YkaOpHh9R7ieNl6H8Vrcxl0w81j1Gc10SOz/1/mUqKp1
QPr8a8msIFIWWw4KsQ3N4q1iTL91OlsIP06mg2vtcVq88m7Pk29uH9kSNghL+VM0LP9VfXiS3kij
vz0I4rLyyem8XEVnDwOizn8r6i0SvVi+Kf05KfjagBK61TP275rA9Y6FKMrMdSrbynfU1CH0Obot
IJljmxJKzxI2n8MD+IHWaVDu33ak/HAyOZZAkWJxXMT4bwFWiTHuqlCXdprqKWeJEmcIb6HYnlxV
5xSZ05+s0tLDH5gwnvBnFZFzWd4GCNncMVJuTBbEI5+teCL126/8TOO8di8ukUANhIH44yns0L7I
/0QVkYD86eEX3KAdPn7tr9EjBfTFhj9viECv3M+ISztc/pmG+L6eJwtVOsw4WER79yepMezEJcS+
KKuyAN1r1rsNor3+HYBaerl6b/RqEIpTuXc63GajxLf3BvqRQaEomvqQPTD3atBGPBHcAqf1OEzz
AHAP+Aoc0u9hc6X5h8fjHLbVBYosDDG9W+xSadH8orp/gv0u05rifrplLvthHBgJAo0dBCTJd7DV
DvUiPzqd0VMBjP6h6Ghb1CnbS0AMYrbWb0BUzg+OufxAe6S4pIhoa3GFeRWEn23bCooKB8gQ3sRV
ZTOhcRPOhAUX3U+LdWGTbXDInYdje0FxhScmRWRqiIBfwFufA0N8MEtAXaCbkSRd/80i4Y5/wIjT
U/DjkLVTLt4InxWQbShGQ4VrzlBSAQtxBh5r+ieRWhMXXOX5fUg5vU+uz2YPAqEZl6Oq7cwNaTi9
jXejiLWR3yeOOeIMvFRaPO1m3W4+xvaTggmQg3g5BhKEaekaEBJ1mD86bVb2QRjZRBf4VaEkF+kx
kkVnvQIfn6t8y2Sdjx3ABM7ZtibTlz9y2V5+pURaGVpMpzP/Uq/soQKQm+1+fPKu1o6MQucdOJWv
uTeIsEvvnHCr8NIXDENYGAFALLGPmeRpP2WLA33GViqVEtfy/DWM8geiPmGIX1sbdXW4C36jipaN
5rxahBkO21QtoPQtFY5dfidbSzKE857AoYokC51s8BLPAyYUIgguJLcSXPjiH00pSPrHqW2DxRYE
SkME0RVSB5BOM5OwhO/jtq+hsbPRKWSL4W/NGAH7+aRqDcWyRj7i8kJ0JG9ZaA5Q9YRvucpna4Bf
iqsrlQwIQXFR6b8S5vmWj0/VMQFQlH91Bet2+MzSBTRm5p3H0gm9+zCGhLS9wHR3/FWFFzrl69tI
r1Tffpnyor5PsdlZd+8b0kzp5UTtz8OV4KC53aqqYYYt7uiIQFXGgmvi2tm6GySeJq4FY9G4SgVb
OLcPBrUFJObKPXt+DLowvJm3+rN4ihrLHNi3imv9uyXC6WLwNO4M5MBQYvWSNZ96AUaO9mG57TFK
1NqCLQ/+naMdOpgXYHzPMIgQmMv64OURvRq8GLU5RmsQYpLwOdxjgGb0GKTReV86FJ1Ebup4v+FH
wZqFtIRS3yGL+VJOdU7lcs2OCFnhjIKpsck1GvZMSvGk7BE2HbOF0WKNzwXDhyzezRnuhUqz1izO
fND+b2/41EJSrQb4XK5TFPXEa/fdDtn2uAtO9sX2pvT2eBs+YsA5WDH0bcwXToT1LBCdse+vRdTq
Asqps2lvOPE9fyVJO+cafOpi4fWkf0JZ73SkeEpYirTuggIStmvUo1nxSDTJnACVz7w2ker1Yo6p
rEpHofagi8Hz1u5Kx8nl8KHztMEmiAjF9dHLt2uQgfpGi+JTxsV1b7qU0xmSoNt9ButB/XScDJv5
HdWYGI+jyWetUTsJCbNSWQgaIj06F2YC0CUNBdQqaPYHfvsMdovoltx7kX0sFtON9NkI1V4J6awd
aDpZidodEJcpsmHQV/ngkMlRDIghuMGdH9q5OKO94MtNdysFOMtPBR9oUEhDdKl/4Nhr3SBBClha
LAYQm+PLj3Itu4mn6uVEsdk4p5l39ctJdFyvkGmIRhHekuW0WOdS+jbG0u9P5eYSFOtCBqEfV6mb
rp4vGhoUpA5KWt42T2qsTHp7mrEd3yEi2OUvbXtl7nswO4qoEtMYiDpC+8px0KZNotWvu3RFXSCG
EnnNs1uaZoVK81j4FF+aJn6/cxcXtSm6VpJbmGZVlQcpG24GCZw8xFrck00IsD1ETgxsjW8fppUU
sdskELQPVb/Z0tSs8aTXU22OR37CohQMjmWdqvW1pmtatL8cc4GkEXCeLQZYokzChY9Rt+8FWNAn
ndPIVhp3bD6N9qT3tjRtBmAWLwJ7gY6SVpIlOmCAMD8JKAHtocMRVQ9roJ++uxl7bVbMJZlIwSB5
NxMDXVAXyAUgaW+VEh7cKjNMSRKQnWnfFpi70psWV0ZRCFyybihOhPAzrsTnbfsXjRxnSSZU3+6p
+5hQ8omr60tyRHMPOH/i798oS22/cbC8a5WWLF14JO7ogS2EQlBv3km417HvkZye8k965eyGCtK7
6kw3szzQLf5K1yLRdefyspnbGzivfq7Th/5GCv+76ZVPToBxUOlyVM7E9gArUOhLiluEw0WHqUd4
sBzdwMOPobhOp1pmwxOYAOuGiTv+l4hWK4g/YImVOGx8nuSMYX004djnM33O9JkFH8A7uwKaO10i
ONa89uUmZNMlGwcDwHIn8aXE1PTiWHgYADq3STFf4mXvw0vRVhnphMaZJD0FYEMgDqTbLuDV8gir
m60l4A3eUbqLk9Pl5YFKFsGiM7C8HDaFvv4dD1x0eI8W9P3u+3UrXFOgB79nhEAmNSn2uxnnWT/I
fvluLyPoYdL50KaB+9x4DCGVl8s7mm0Mko9l9NXJitp7dM+hsuA9tJO6vttDKlmDKUfn7XZazw+t
oMs/duFTan77n4lAPTFbrvsI870nURn+1I7iS9KH+iUCD/guzdFC+Qv8XjOqOmXe2g03YHlfniqG
KIBzN18dy/2l6K0bNF+K5b3p94MICn7vDLNchrPVZmHVxUvVEK1x48s6KQrCZwXp1qdso+zsXa4y
JSfV2XdqXFYAPoMj3fuOaykfr/6iORCZPwdst2Y7gnjGv1wS0JOJbtwR+I/0IY4rqCr4rS0yM22o
dytvDkwQX9wiKFJXcPMyyFb/ebRHAnUZXGvpy5Loc+vcQ0b8O5G+xvBJFz0l9+E7/aGxWh/XAwmp
QauU9iWkekL7KvO71D9HYzjBYyUOdcp+WtOIyh4gXnopjzb8MZImX9MOmiuBkhKHq2HqQWefAPs+
rIZ0o1vmWKC7P7rXFEfcHnkOS9GZz6uEMfLdhYTZEXnImnai0bltcaLl4uij+5Vdf3GHIjXo7jjf
UzLwKzdqG77M/lw1bDJe9MwtdWTDuQPB6Tj+EROwi2Lt9I+xBieRbx7pzxYbay3yKsWomyUYSFO1
PljyGQ3h0n2QzRgcIxBYxzPL2lPtyUItLw6hWTc/WIpjGvNm1PdZVZDtXPzanyxveotq8BZOtM/5
ftwTZvFWSfwh+qK+lcuWhRzreLchgn6JtZmLKnL0oyV20JC1iaOafAdbp9G56qW0a2y6Mo8mE++S
+3F1yx8vAdNfeLN3nEAQaFds9bkRjpqUPsCXkKsJ6Ugn0EpdkY4W3jzBYEWoH0vybcZ+kdm/QZRl
NsfI03fBkKvfrcRDi5ioxbzZTIwZyGXYZYftZ62Fb6P3FVhEOaUmJwN35XpS5hyfvYoj89LfL4ac
+c/OFAptW420orY5DLnkirWZi7GyXr13rdtge9xCY/VfIl31U+sy16Lx1mZ2LWLA5MSVmGP4JExr
71GwNjYTQw8n3lDv+uNU1Hm8dNgyWbDmFEbMMqOcjYig2JmbbyrST8ezTsFFYKOqwFtMM4mezkn+
H6P2g2gA4f6rN0AOTF5gaE9aOxOOXf64c05BhaUFcmrHfSUJrwW1LYakAS/RSiexciMQqBfiT2yA
+6olAOHVTRvRrgf0DuMBBrZ0UBV1E2q/z+V/NH7fB//kayPSL3r1THVTaAm3Uan4N0EKBnG7Kxkf
KdOjNA3WaB1ZcIX8SXidoD0U6nxrOk69LfeHJkANxCaxtrloYqTC6FCoxpYLScMaJ6DN+/bK3gJI
3iECIZ3kO9lDEG8WiU4V2l4ppcz7bKlYeCzGOkQ2YxSkUHVHmROVO56K7Gsup+FXxSpMD1/+YFTj
OYynToEsOvu0gIBfpzff7ULfCzPQkJg0LSj1/OS9zLQrxwJSM/PamMn1aF2GXaSOpQrCI4TNMAop
qrFzdXtQ/BG/34eitzQlDFI585Lx5xicUNyXb/CWY5e3SDTwgjJ8dQKjx45xoWOWUznAN3J00+T0
VbeFVTHOhS7ET09GVob+4fpWv9tSSiZMeyxm/iJDVjAzEeXqlJlk4kKKgXQWfLi/nrnqsCt0KlUW
oVSdNj9A5n9Dr9FByFFmJpG74JlK0rmMPtoH7awQlAS9wGIANfr42oWttkoKVgPB7yj7a3V8lI4A
R1rAw6lRyLA9FGVA5nn/BFLcQoJMZ1oWRrg7nOAozbO6X5pc1PsH2CiozbKEFoxDTxj7J0+ZQgwU
Jt6qfbjuqTnUZ8EoUi6HlJyOORzSfcMpWh4BO0/q7tHMdBqsMY9YUpRXIRrp6lB6ug7jFVppQwH7
IcraBo4sGVKkf/AaaXl2a9Kl8K2Z6/qxeYO7GweIxIyYq1Av2F/lDf3USOHQrMnoCh8hRa92Bf4R
0/e3+70558UEJgUrWNVAAj6wG5Dp9P/1SI6zIHbB3Mzw77DrxXl/LDUkgM06tJ/bPtwmt37Hkaz4
wkCxofUR7PQOzi1BFmem5c2rM+AIaI/qrQ1AhTGnIs3z/WRch0w3DTtm4xfoBseQOnAGPSiIUYGv
Al34/wLtzuniHFi0RcaM0GwSyfrlG8j/wYqKTpIQlpoCPcH3CuKSLXJTzYyihcmkRhv0CqGjdZMt
QF6wkGKGUBAH3tGqsbcPBWlrxgvs4TKCdxBdNC+h0cXvPcPhgI8g+9DP6cmpbjzsyUSgbpLpNZ4q
7JEL0J5odzQeItrMwbybR+BThto9Jr2XoloeA/gJ+J16FjAhEyYP1ha2ziNwlo8vc2wfneWPT8Vl
tc9J09gZSvCi2MibMkm35zLY2JH9R6udzF2Wl21VRfh7Cr0gZRBJjxwbalFT1laVXn33sOm3pnSE
0zWwjdqiCKXcVUa1NGg9+6R/gJcnfnfJND1DkjwA+E634ens8FSrOhVHCT8Mpn6dJplQt0XymIzr
fEi+sWFCmBOC7fQGUw9hgyhtUd7r9cx9bS3Bfh0PGyXdJG7LOVILX202r/pDaRm2p9SgYJW/Iojv
As1rsKRYoLlfb/9XdeGhstQ83yx2XgimXqvrnTXvcB6RjLd7MdhYrNZLHqP++n0Ef5FZMcS8dcOM
cZzbvd23ynfW3thgiicpTS7c8GJaICCJ12ZMNxcKHjyIvBgy2f3Hy5E3zGpT6KMB6qsy3ATaYsxG
oz2MCoV0icb+3WZTSy1UN6JpckvuY8ymMNClgDxd9TWTv9n53rJD6yQE/bWOmk5U8lm9PkNM1w1/
fP+/d40gT10RT6VROhn+LPuzvi2smRBkU1iNnDdsntrDYHotliHLAwkTqjm750qn3seKJrSxF+lc
l5M1tTmDjM/YeiqQHOnvuYTYSvafIy2oTJhEolR20xEx5Re6aqI5iBlvj8Z7DggFxoz38SHBlfIv
oIwJxJxJaUKE1kzRrcIg8NTk9Il3Giok3/1s2KtIeI1k0Q1yT7A4oXJ12+q7Vdsg5mhfjesICEcG
z/zFjmMpD02eQ7rEkLH+2M9MxFn8Tw06DmkfBFkjmXUvfRmdSY/POrLbO8ol8OfQjbGWeoXzS/P4
4erEXFQcKdbSwtczj/XNfxpriWnImd94hT5BjaQWQI8IFB5zkswVb9iQxCbn3OkOwcAvCIPQTzXX
GYaQfPZP2/s6A0+SeOVwj5qWePvsYPLCX0Mx9CrBG3Fnuyf3NTZk/hUMJbFI9KrX5qpNyHMdWw3b
KiGUQkmZzCuOBSWehUzPsLp8lppf6FSChSlPxgoNTXBSJvjsefKxdeVsCKuL40K48PHL6c4jNy4p
sS/xdfKhC1I02H2iBq6vElJS3J/VzLTY9NPlYpaxvVmQDjGFIel9HmvArPOoC1wlYW/+S7n3r4Ui
aNckszEJwD9yIhAuvZTOCwP/lucCSLjvQOrbW5OGK2CzLyd9VHTAtt6boxSF0vi7opWdXciA/2Xh
0wnTkAvrzn9ycaSCmEP6DejQ6CL8P//UtqvTgMDq1++L04oAUB1ovdSN0x68S0ECoa3atWbQZntW
sfyENpjM5tN1i7bxilbtFY+DoaCLnBAUr0ZgmK9KS6uPyyfwnwSn5t+R7bDOXMjM8Js9yAnqp90M
FR5+/piJMtNlSMXg9yirsKyHbQFiamEl1+u5W+rczeTwtnlc/Sr//C//tkvtx+DpUzU+rS9847vq
fBjhB9ycXh9Axrb9k3n6UBUgwSb7HtdMhV1ZIXYFrF1Xwy/45j2+vw7QJPmNozsCrm3N3a7a3XQY
+azrDW387GP39GQ/RJe8cWI8YTHF/pp3Hw9t4dEPKprwatOZui4XKx8BGrOWWDjne69PQWifCfBS
4jvUAvIKc+Hg4Q2OeXdxQ7Ul6WW+T4D9fREoYpF+oJYdeWxGFNIfqU6g9VnNvzY/CjK1DuHMd2+x
1jwqs/nER7xbX3iqz7loYb8xnJkaC+dtKyDDsep2xJheRIZfnHJLHiFj0ZdUnHrs853yKNTEox65
6kJQV/pkCaCcyic9C9JGI1HrOaf+HrgELkoEGufGB4860T4sX46A1YC5hdadbDCp9Ld2yGbGsbaa
1YUG0Flyw5ZTQ5rhBK35Oapfhya+iY+8HiLNZh/Q5GH5/N6zGNR4VkPbOipkFwOHkPBNnQ+F+aUc
LLIvbM2nOJ/myMT6jWeK1PgGZn349Oy7BeSP4UJISGd/3+c9ofG3SHXeff+u8hFi6RFWFuG6up+A
Cc2rFb/sXH/t8x8GJGJfyTK70MLOz1pbYBavfouZKykVnSjtCNYa+oXlf9PBzFF1thuMty6oMUWs
pR6T7sr75FjC53cpOjdAI3+gGgq+LiSe7sqA1Vr5m96L6ZIPc4+fM0iCTuVomsMRtNmc0SgplodM
RMD/2iSTDuddYX9SWDuf3+WNrNowpqUUmasWEpKVvwVvBkTW5HtnJAq6u+y2LVyLXMV0R+qQ7a0+
tCvCrpg5QqHXs+bmf39aMBNZROm4xtoXWvsT6pPdZUhqnHStf/0BVUCEcVS0H8CDPN4F1uxgdZjF
4tLjWv9KEaVtaw2ihgyRW04BSb+W4TogE5ELilSTGhWz86f0vv4DiCAGnwUkMDvCRgiIM8zgygf1
5u8U2JjFCvMeJ8VokrV9wwfC6fdPPzV4DcnBbsKPtUz8n7BtCASj8w5dTE8vc8h4Jhfokx+t0ZsE
B0lX9Ut4QMLTJCSwGYyyrj7DwLOnzs0ZtwV3DffDMk/AfIdlEOMM3ix46PGrxebQaWRGRtTwPlNX
7VwM81mtoeclfCYD/yDzpHOc/KcFNLJZ+quKGWEQGovD7jtdAfRw752ZkLrJQbdmMeiv9ajwfTkP
R79wcS3VIf8G8eGYGwbnfR54mptt4n4ZEQ5OxLMiFNfVXnKwNqYpaV60rMS7e5yrXz+qPvSGCG+u
z1JOzRjGOw9lkZQDo7xk9BE2m0iIu0hygQRw7Myy4XPGHcPKmlRPBAYlrHJ9yXikkdM9Xx+jC97p
oHUMgSlH9kBDEw36NShCcm63h2UhMzjnuqxx+2ptbS//TW7gCTW7bIjU85d3jIec8ZrqpBCGBZi5
ZcHbv0B/0riarOx61rz+ATI32ovARA7DX6rGl9Bi+uTYH7ZYis4CgJItNh+07jiFO8w1go31lZ6G
j41LUjieP4N032fMEexHgcQKnAqe/40NqCv7kkpi+dLeIA+Pkk8FdsVD+Q1jNtbLeDQG/O5Zuu4e
eloc5DPgJtYNE+7SCRwxQYb1dUGmxrHSlxTLEvpae8cKoVbhvoxSH8Gm0939OQJglPZcgMUouKJG
LEET5a3u5H1yi8/QGw3AhHbjEA2yvF8B/HnR4fRZyviiSDLuj0TT+wz2JKLikaXEPUuhySfVcAEB
R/Gkb2bnuWOaLXmwTi5A5wwYY+z3qkYbWS+QmCU51mNA0njqI1o4/sTlZMlznL8D2AMS38vRpgC7
5dHjd8lv9XIbveogh38LUSEMpj0mAtl/jBAJ0j6b+unRF1pl0kIwp8FPpHbA78DFAuWkYL38axNc
pueusMY0Fy6RCWy/RuirzqO67cstYJDjQuPpYW5hMhFv130dJSLUBnQXkZ915ui4u4YatsLigZCE
BelwcGoAvopX0M5vef9qgzYc6DBE1ACP2KnLIWyM9jpeKtC5GwEVKpOyhCpgw1eSKQee6l7vdAjX
GHsAlaQM2VUpO6zENF0rc4svrfj+wzAjqB9qw00LU4DpT/TZ+1a4w+EdCv8n4Osx/2CmoFEtLINM
ZDXEdMNqCQjm8C2QLwggWsRBXG2piXi6AENXpkc8EqJ+YWRPq6WMjnshKNVvJ1zc/U5TgXKWz4D7
pMDgf/uMwG+ja6gW5LSqzAvFpuB3bUTu78lThB9ORpm7lCelZHcW9DWTQ07poOJ1nJDCm7h4tx+f
ZxJ3ofFos2suLES+sbSqxR8HSVeIYhRUhfMg05QDd25yxJs4MdwIdv2IbhlpIJ0U3UDPe3+tMJ3i
P4pnDwu8EmwbWZwrc8JdB2WSOR9OVwF4pbpuYXmmUahLhnRO144YZHdP8uB6trDYWRbgeoqm8Xes
RmLg5lhYDpPHX2ohaogGYKTrSyaXWEQ1KHKPttLDAMsbpXn+dm2WbTs3x8XWW7jBWXXv16UVFxMe
gux+DdfNg8jAe2Ukn7PsVSRYcQWt0ZJ6NA8+hgGltNSKGrSTLHSRlQNxVhOf3fkbzrxKpLvJFvcZ
jN06/cUQfw7OoRi/RG9sWPoKZVePu83xbtZvZ/bETA4S0h5haarj0ifNNF/PCRUqsrLQOuJlzC01
laVm8sRw1t9Cf8Hcpi2vlhHINwi+NYE715N60ObwAT4Ac9CfZNbpWnVWjjebCX9Msft32wLhrp5v
NGQM3dE0xgJobyXR6BpQYkXEo/8n020CdX4yqasGwAKMQmDexIVFS9Rov/S5R8WC79daXg3oPq/h
gyE2sKQqZV+SGZt/EHvK8GPvkWmFgjwxSksJRO/pef9OuRtqvKNM6iMeY1j1hjtWa9dwzF+plkxq
eEy7qkE3ujxuAEm+GOsJ1+7l8bK60L79whTshxXzvea013lbbXDD9fi7/A51GJwIodTfkhQ1zZ6U
VXzvHOwFH4zgdGzs4Mp12LSMK++9fTEUpN1FTZrIRK5yKomxuIQgCs6Hi50vKBQ0WjtLbSBePw82
VGvN/g42q3XlEF7uDnr4RCNTHB8jDaPNHN9SLrX3Q/R+ZWik3vwf3vbtTalS5NsL0t004IQZKIQy
8bz0pBssI4qTntS77WR+4HTZFQbOVvN51a5WDwIPi9i3CyGOHtNL2+8dzM3lzGXKO7bhGVwEykXY
qACoqJKmTXjooxIdkurg6hpW3P6etLzc94y6j09NdeKahx9sMu5vbNVcv84ZXCB0/u/uAG34w5ct
MTeK/xuJg5sZZKFT4BtyNztEqrB9EBMouCexRp26O+tmwzu9dBaBxdlLus3J+ZcM7UqYIcsFtnXs
qhg0J/OZ1YmKXvnnd+IM73oWYnvZlr2shdVxsgWhZDcAvteCOqnkSnWr3QbT8eCDP15CBXPRJ6yr
1x36unpPlB1RlBlN/II6Zm8aY7SQIk3gu9HhX9Zji7EcJ4ZBu8ie2FjVb3BehRXOZZ/n/4bGsD9W
Weki4OuALl+G3ulL7hSEPjS3cvjs5DB74/d1zJyjDHTmLkPF5/loY0rXVPbrCE6+9/8DkG0vaKek
0Q/7pV9Aq2TXQPcpy0SV1uN3yRFmJ5oY0nAoXZvtA0yeV9GXpVjCbN+U38q/fHYz/UxYVr12/CI9
l6CtgvFME0yYZ9pd/dWXkrMB0PzY9nmjMNyNSV9n1W7fsKgn0go+k3kc9iGJMuqUWbp93PLvhWzi
6oI8G4g439I0U5tIL81g5VMOOa/9o+Kt3KQdDLJhCZQnXhxbW0JjBzIMAEPYUHdA5t0O8vB0d5e4
yGYnK2OQaDEpw8nU6Mwi4xpUuDP+cCBipi51s0/fVMqJYwdpjOy1+I2pi8g1gZlFSjc79GXplJzw
5fr37c5Q6KhW33LdaPQeP/lurlWTbsXlEQTl9Hea6HL/aASU6+b70nnm7Iw7wNLJ6srL9xTQR86v
w9DVvT4IPRExBL9Erh19u/sYNYG25c0tVrHqVZYJQnVenqbXtct5maPvUoIwTz7aixHXPE29AVGm
XaUdox7xgJI6kntI5teFQr5WP3ujXZ8DEr98/nQuWROzJSJm4vpUE2MrdclBz/wSzmQ1fBqOXELF
QkN7jkxoupknpzasTIzRS3UEC9X3iIkHOKYknnn5DzOkkgxYyXKgiLwOk3GzD86WTB6hqwGJ4Dqe
x1CE18Q/4ykvhsuuHJtyEnZegmg2g8n8n8ezbLokjQGynXDJVKUleSBnbcyL/8INY1Ns8NVSvA6i
QDmvqk9mNRkWeiiMZldxzzPuCs4YNZOrUHFEX3EVqnpVSHqAlVlrPiJlux/VZfjdxT5iRju7dTyB
lSBN5UaaOp8f3UWqZvOEzepJck798nUj6slkRBtz+k/S+5Xjwgte1teJ21ieGJqchUtvRQykTJdv
ut5DMlEr0zudEQjOyVzswYOmfhkLFCvTv3BvJD4WlY7piezs586WiIZedX3sd5LUhW1QhHdaaS2Z
SzvIPVgF9vwXprqgRJsZHAVW/sOQ9LBjRl98S+0I0RqRLh05WzF6S0duerZ4QQmjOPcLiaymdueU
QUJyTcbUw8IsoLEQl+1P9CfJItWdCQ7G8tPERyJKe7BwsPTuoZSE8KLj9N6nsWqKPcmPt4e3qzuf
Tk+b8Q0nK9wwNNyUMlicb9tCPcjN/LSuou9T2lcN3XytYFW2KQNikAoFVU28L54ZyORuzuqGOWa4
KGGqTha34dvKzIKVhYT5fmDQZOehzLDJ5zQJl6Z8cuOwG2+QC4RUBdBwnYJS06Al2wbW9qOw3SyF
yI7Elzjrt6i/WNFtQEuflMkRp5E65kmMXyjpdA3HiUTOkK0XYVzVHUAmZTyvv/1P1PDl8vR0htk/
dviRyeeVAbf4OOU9livWE+wh1VHCJj/xeqFMX8MP5WfNH30Y1AR+ZjLGo6e2heorVcsOvXNvLn8V
GMN1sEHuNPQWYsavwIIdw/nsqLLvkAOXoZGr+v0IBLLwhCorPaoFirqg+Ad+EhTEoYd47/Ip9mXS
y1eWlB1ILSCWVhkkaY4QtgUSVzrBwZP9/BbrKNeFYkrGgFAOXsdH1py0HgUEMdm+SVGp8IZ4TTGb
j+OeFs4ZfH4xKrzml6Iy0N/MeAFAeLEjy8MtPeN14yfZxd8wwn7g6ZpqMnn/YAGWxRggbnb5LywA
p692TMDTKvWmOguLpejP//IS4OLboavltQES+OHH1ZpsohY33hyzpyVSGBRyAgjOxvIGZD75if9a
U/NiAqrfvUlthlKFjcBVC+X4HepB9o0ACWHEnIRh3bFzy7UClt75dPba2sq9Wl5argCyyHCKDQ1b
t9wfm3cqwJLadFw9OJ7qsEN0kepINrWef2D3kCDSD12S4QN1AwEV5/PXJc4UtNZtGlzg170AYqBY
TH2rkIwPKmvQncsbWLJwFPXgBk3ZbkxX1Lo7PXZv89/jcg5FgvM7NokKLCd/ImyWmT/32qhiIECo
fmq6FeFj9zqzmr5/F+6yNrrraSmyAXfIBVnWNch1PiQluPXDyvjbiG+lR8pLPfsGhm8gGcRx+ML1
2V/8NXyX8NGceGFczpKQgWpBY7cT+oK5K2q6S04Gti5uOOt+3t4ed7KsA7FoCXK6LdoEbgwM+z4K
KpJVxOf9PIjgOh8XxTfIOdhVGqqLhRqHh9aP+v9WquXqFXJRJbiIR/yL0vu/eY4/9xilcc6FfKqR
x++EM878VokQK09stbBdxr8o2nToHfLs3p7Gr5DYgVUOWzqh5PdmgtzkhRBizG2k9ng1QZZl+Xd/
wLPVhwHhkWBX0fggvCc2CkyZsfCwp7d/IF2N2lAyI3+p/DGPwCOnyaqqxGQqQY4W0FjdzUIOj3If
XF7asAyXlFukG/Xx/GxM2Cz3EHV/VdxypQWtPeDoSUL8H2Xa7nCRZt7ZyHgP9RmmRlsd2/lelE/4
qQXtmJvN//mgZ/oFbSksecUl6ZDuqR0tmeznchzue94TORyo2Jsa1Si7yf/U9N+rVvzxLcB8KhNi
C9fDim9gFh5ZqbxThYIDJIH1kvAYKhWla/sOFjLti8pg0jdUGZgcHTxi6JG/9ghvbaAUEEI0Vcws
uu9GaOJrY7rUew3EowsNhos07KhYy6pzQKzALXgfqvT5i2PjcIqe+vn/tBWNSNObche328FgXLzK
LaL+SMC57tleD/40P0b80/t+DUfwLthL4LpsLUYvugEahLWSAUIVneWmRFEZIQ+R0NvFZF4kIiNZ
QTVmRilUhgXBx75vaxygF+akydk5r//gfGaohSDTXSmo/57su8VkeN1JeuAa7+/PK7pH6etFnzRw
t9s3XVFkKOq6HkHTFA2Nvu7VKRVZJxrn5vPxsiPQZGhrXtaYKTE7soh2zvmaC48RjAICp3lqeMae
5ZcT3vKsKyXHNpG9u2apSssYVLUtDmysLEgO2CGYvILtuojOY9bDPHp59L4WGRc0OeEUoMmwPwSH
fEUi+rUbqCbXb0+a6FdjM7ESmpXAC1jZdJGh1VOmANPcFOq0tRxPNWBEVCcBnVYx+VdM0GbitVsZ
FT0D7RBZ5U0zEwW5x4Q+tSyrjjOZnRYtTiPZ4TZev3VSShPQj40r9YOAPKmPZvMLQVBLdoxNcStI
mJ5r9svODA4ZWf1JcDGQmOtGVeVAPkhJMvdaRmxUecW9e3hqAN2jd9eUqZwHtl02Iu7HgWxqUFVk
3mk3MyBOi40jAHUqG2GTJ1Ln1g6z4ONrsMX7yHjxBDYJZhv553HxbR9CrgeIApt7BegyDh8QsWYt
hijcQUMe+PhKlkfomk3AwwQ+vzjpQXcoWOihsUW+DfA2pvXgQJE543FpCD86xyDBEWOTYUPHCBLc
s9hUvZGRYhexlpb/VPL1tu/4GlWO9zzSLR8kgTf5EoYjQsXM2P5eHYFBSfvcpV3nukNWO2CnRmBs
XD14IIKGossQHwpv6zM8jOn2P6304SRjcmQqyw4TOpGVqG5mtXEEY9dZCwTUWSyoWCLBjfVplyQE
FWmLt+B+k4rxydU1KVMWYQdjEQI1fBvkq0gFQSCkC5AoVBo/BheXLywwTA3IirJWKdJxmGQubbAM
rbF0l357nIvF+N7uSVs9NaE0opewqRRzd1mzHEN/YISVZtSeYn781pX0kse1/hVIqdcOqwDh/89c
SZwf0bUlwY6881krcYC8gdh7We0hCEqW7y8xoaa1c6+wRCHE5zP5aPiXIFFCZqDUyukLZi9WJu0O
BgfaqdqtM5eeYScqbZ4/sE14wbcIJh3Rz/+IN7Nqi9Lxlgs6Kgglh/UkGfn7Q1PQJbFktZso13w/
ZOYZlPY8QwDRGaoV4WpabGQQkaqy7BT906wXlFXFbuilqIl+849Pxx7DnL7j/oC/3m3yap4i8Fmx
ejAghpIVD9ZG4iIuKV+R+cMtxRJm8SlgluShUrSFmkpIUQ5/hu1WhvlHGBtytd37X73UAEY4FjZe
lpFLXang/PVrRrV0v/p35NP5RceQ5yqo3/lAsm+GhR6eaaAIWpBWAlgwsVGW/CBqROiLCqXMsEf0
NMq7cf66D6a/DPZEL5uQ0Wf+W535tPE/xOw/xCY3Cm0Z/R7qNTsax1T0v42tH8Q4ZlM/Rx/9m5l7
EXNVnKP8YDWcLA5aMOLrht++WKwRYFILIb07zEQlcSXWFx5Wu3nGq93qB4ydnGFYVwKFom82SZQN
tmrPm/Z8THRD+2Vir7Fweeo+1ic9922EWtDtIbybb/fQRsHBGYgGdgFrH/5BMvSYMnwoQnIZyi8Q
fvHY3xOJskJwnJ4DV0uGIdimvfMFFDlx4zAsDZw3dlIQwqoL2ii3wvwR58NlZ3TYLFexvus+0rVa
EoxwwsI2Vrq2OJq+QZkAfWPpJ+ZI+/IXWSIXZf8tv1NMA8HA4MI42UUdqrtoA0Lhst0JRXiPZ8Ac
2mLUqUfLDMdGc/vKzT62KdDJL8yGmUfKVbjvS/wR5zBu9D74dtJHuCeaMkQDWWE+95pYqU81ry50
AP/ZUuuVUJrAH+pnrycb16nVjs7iNid2IhdkvOjWdhEVAvv2uZOoD4jkj5XSzGgl1DaJ+cgUQnzr
W0SJkXHFurib+OsotH0RqkD6DlpeRHQib9wEbWFsScN6BrIHOFIbIdFY7CJn5gJkxohZegbCEbGU
Ovb9YU+3iBkPdzBHH5evQEHEju/9AeayIlbujbZB+GuEzjFU8Z8iLTOc0KpWW/QvSqvOjhAvzrn+
R7cQ85QtVXimjYmHfk/Ok5p+NziPXHuIrTXFFjqR9MbWAT3zsriElvrpH+070wKY7G99kwtZdkMo
g+3s1Ft8PqDJw3jgmn7uh6tD0qSa3Vpm+NwPX/8wJ82Eyeg2dFVK4HRTlXjLPrTX5hppDTM+Bb6v
KfzcG4lzCys5UIc8N3QKSkYxTuRj01h0L0wP5I1P2xwGmWgpgZwKY2B8d7mxXK5lFTu/+1XEXAck
CPKFNzfyYLGAGceb7LVMegXTwtGvO89vrhPw4OQdg//HLGoEGrptrqmVRi9SQQ1CZZGe77FMESrz
bNneA7MV3SHln09FZuA63VqIBX/X6rNFreuJMovD9q8+4ElUE07DrOZiqWrgbJm8Z5BEbJyP25k3
1+7D7iVT1Pm0Igy9gvXDL9Hmhwzo3lxxr5d5FfBlmIitBR62mRokj+6HCAPBc4hS++3YItycFSeX
QOHFDS3L7eGcE7IAb7ae2ybXRKF0kti/3VKwmGGetnlrmVk6hdK9jbhvLDGTxh7reLk4HYxOmZ3B
rnhY+7C1XnWRPeDXc1tzhsGZAFsTjzdFOMTWEvOobc2t3cYpHhJ9T/Uv9sNB77nx8dd87q23M4ny
f84/dIodU0LJlSQb5ElqNV6z5qq5ek7a8HqHuauSo7kBvIcC/aR0oXjv61pmB3GBEmZqPOm5LUsA
eATuLY89+b0lq3X9h5Lh7cSFNvGDYAI1wLvodTR09QH7o3ujxlSBtftHuitQn6GUVl3ZQdz5oTVI
dDsXtZD/+U0FwDM7A48Mcy5+NXeL7lY2GiGMDZEEP0chz8zR80k86CwQ21dRaKfYB4w+MtwmLF5W
lmI0tMqexHI5l95V8WSVKYSkQ4a7Za495nNhQA/VWFnhs9UwakMmDJIG7GFNT7cIQpjtfcRE0sJE
rdyyI7ZF4zXm22WkElSg3M1Fb9sLaV9rNq4+eQvkeMCC028sZ2XQICIbQciBt6ZcdDbBnVEnqFHa
LM0/s+6Fr9mG6nocrgV0qIbdS9wgHxMbYjk/70kEl9kXannf+mKSQPVoLSO6Rz71iE3I6YJWR7pI
nchQP48ura6Wp0Vsjd54RGCM1R5yNnYGOGvHQ0aFNDq61yupu7057/rM0FqbhuHtuVDIROcx/n6v
KikEhinKbpREyEPQ1ofa4NiQJfPyr+1++Rj+CDwizf8jJsZegWnkHxdDH3AP5DC49Fz60FVSoZuW
Z1kJtHKal94zu0/9ooVPWbfFXqdye6OffpH/ulA3mVnjB3OGcEtVAvN3AnX/42oPgyK6hCTQ6Oo3
zEzVj4KIWpHMw8Cy1D9yusAciahYY/W0DZMQX6vuVY6zbmTC/XOzDAAyDAnnHcaoBZtZezJi7o5Z
2s+NlMOPVjowGjRrKf940rXN6XWpD9aG6iCF6NHgzkDwhaMolKWbr/ozn+8zCiXo+kp35lE8GOBc
b/UA0gwX7ioc6OIEZb5DDrI01LCLCnhC64IvyKxxYNzLtUmCpNk3TlA8AwtKbMVVOEg2Eqz9+HW3
hcpERwseUKQOm+ml5xVYYMdeF9L121Mb1Cv36PRcMpXoneI93KvHOZfdWBePScPmC044/PCES/Br
YEuYQRFrSJS7yrIkTTZs5F0/65dRisbAp5TdlBgtVGCCWyifF7DqeMjvra8mJ9MTfxXLgzVl2X5D
2M8uVkNJ4vhfxHUZ6KoCkdk4YAY69eqZbsKR0wMpDz6oBFYt/gQWsl3neRUKxp//Fu9pFJtO+je9
b9bXHMlxalpwqQd0SZcPBGL/eVjXU/FT4UpzWr2KLVu1BPEO0FOD4Cvt9ChfIQzTspf0JZZ0C4wF
OewfkGs0k5ecZSweeZTJELhe37nTavj6z+pSIRQ/PWHbsCNXiVBRuwLq/j6gjTYNP99mZ0HGukYv
8423WT5GmMz8MMK4qnxbrEAJsOWqXgkf7LJYmqIvAQO69PXK82c5+x5x6gEcqLs8fVGAzEiao+cH
VmIQGgOZCF8qJ2EXRjhgYpNjaHKoZZYW8us5oDETZeadXlDDqRQ9uRzQZkfgvB/pIKg/+LooIcQv
xQOFNzgg0KxlZ8OWPev+b8mMUP2L71rbtcFjdNRtI8KG5NEGkxGYD8zlqmgui/nno6Ytm6wrAgJN
Rmdc9zyexlT/HRodUVUBe/2XBKji6jLDp2jNEDIgHQGJi3XWIOqszh5PWhWaItZOzkZLqmYMHjRh
gqGkeKkm0DaoEHZxgGmX+U5HjDUHas5bGpcwRmTGI8tjakrbN48eX0U9QFfGvpD6u7Uz09qxfR9R
cXg/6awauh8x6tx06XuH6RX0gn74Bo8USbSdYdNfd3gWjaLxEClIPj5lN+O3NNx0+Z+bWIonHvz/
JRP8XgxICuk6IjDfQTM+dVHiXqZIoYjXN7zHlEK4E8QLXNdPktBfPi7DUuyOumY1fdyqv1XAi0Tt
p8BX51mw5EEygZa970sYJ7cZBfeBbWnHMGBNv6meVTrhOm4eD8Nxwuht3j+ghx10jvJtCeumg06Y
6sqa1GBV5CARSD6WL6Xhinjdx6ZZdOrwZXmvV1urQDzwojvLoZM1jYwpfOnB/tgMTR2Rawz+DxmP
JdjI4KZ5kJyYDFj99dUWqv2vkn0JzOrYC+E0dZBhaL9o+dGPpf420i3A776uWSA2aZvHOMBebWBu
4qdlxvPKzPkq1LL/t3fDlCkoZNGBrzUxL8V1daPPK4keQN+u2Ay2bgmi/HJJj014xAKKJR7uKevN
aiMP58/4DTe2qin9jl5OrG5QeeLiuWdyPXDx3lNMHKFHxusz/YMYRFZvnTCeg7zG71+FAHrcHx17
+zAQYi/+qsacJTXXXQYiiMTOCJ280e9IUSZFl3Ld6nIiKWvyne6aygfP6ZjBtAwp9tFfXrZG+UTI
9cHTm5x++tNr4NVHB7+mgdHX3uPydcKRn9ZXodPMcWtzgVPXjaNGMKCIgDEbbE0OmdLDhoxP4nfW
Numot8ccQR4GhcmHQ2IVRRb+fk0+hkHNxGgI62XeCFbfROt8dWrsbJyWWZQQhtgRT4ahWk6ntyn/
E7OzFKR1U4Ir4VoUh9YYp1ksVLKU+U4+5U9uyV6jmVRjvjgzZdS/GPH+k3f9KcChhamUaTEmtIeb
TkmVkuSrNXiihRd1z3oyeQZpK3ZTUr3yAA+a/b7YI1NlcQp0tyvGW+4LgYURBnQrU4r57UV6EUSS
7TVukNQ9+y2Xa/eEDIllWx06y5KO7PgKf6ThUqeQVAITN0p4OrgzmusB6WbSFOWrVFPLZPY5x61q
1YP2Tq1yk90HD/ayiG16lFxb5ciJjZcByZNPq39SwQQqjkpSVq2yqbMN2wblkv1yfTcYfD79JtKZ
7gqwQ1OCCquA88dxnpaLrom/kLeqzQMMfruZm+EkhpKrnid1ffRO2os1H5A9gFBzVMohw8dyhjhk
2kZ58zG0KFudd0yP3ZRxjAehQZ/fkZB6Vd6Fh/haux7XO2SH7tE/CWfM4Qdyevv9IZPzsFbHtOjB
ooeaZes7h3CREhnu6+vJM7Rmg5aJ0tHb6xibeukZIsWKEJmcHj91neDeksvU0Cj8xe4iaHWsTOQS
uu2WvS0h4/8Srcb/5GeOjv1F9FLNQphi7tcR//PDq0+v5TQwp9WGcjxXhYTRdh5g8cHDvJJnTU2t
DZOU4b5Xfyo9zyl/8FqnTOVLZQZ0Gu4gZQnSRe/p+tKAFI1bdr+twpVzKnOcbmVtfBNJ/Z0Hhhqz
dfneM41vBQ3kn85M+lo71cceygQNHjuc1iBn/YK8/N+bDrPqjyXb0FNFA+GZ1ajvoOsQHFIHGZSy
1KY+tibnSW7UDO/F3HMm9OCfNiCvs4DVQlQgNSs3LQPlNQ8iTv3KD51mjYB97SBRX+YR5o8bK+YG
k39GnRNtF899xJQBxmm6zgB7dGs5iCPrpSwuXhDtgiNKD/qbd4PsFvD8poVYECGPdG2TA7IfBG8r
3EhZlMcgdIvayh7bYJnu2U6r3KASxS5E4seXWAT2FBfPGwYnQ0BIG5UTTJiLWD2M7ixHSC73LGoB
UxO98lIzuj61Dof+JKSdPf7jPiT+ZtZsmWEVPn5b5PuCNGiaXiuUCJ4uD5k1NbjpdMo/jaVaYSUG
jZABGyyKwRDmwYz7ytw6WFiz3UyzSXydUnkBEVmAsQ4VQ7JZcE+bfTu2AkbfSHmofQhb/mcdViLg
XHPuDX327k582lW3WIl7ZYpBaYoL5ziDu+Y88RxXGwLs0xqLnnjlSFT/do9TASt5jHoBvSini2eT
0s/NeouLBXnO+32K8WxhSjwA3jV64IaApamRKoOYdpVW5s+418bSJV7wBXmCphLFLchMVFjvQ1GO
OJ2kDxZCB43wFQSwov6rvqqxSTrmRiAhqt+vLLdkuHjcMOIwLgNmPHz8MTIt3b9B2PUDvBJPfw92
PmdmCBEOdOuHVdZNcTuLmzcy7md6irrwCi1BI9xNPHSxlqd9ZpHEnR8S9+04OtzaQ9EJvJM07K8L
BGkZNEabt6oWAjM5JGDzHyTx2Fuf6+TgKL0Eanzg5SfOVR5i68EID86viFGuBMYWy76aO8ic+lye
Q7fPFvBnoJZLUN83tRHtZa7wMrwY3sjno/JdgiP3EVf7NqlRy+MLlvUl+MDyqTqiq+Hfnyn74LAZ
MLKKeama54Ezj59UrJoE0AHQotXLSQNdEtc+jvc9f2N94krgVUtT34lmnDIJSGwNV3SRZkZKmF0T
R6EAkHW+ppAF17CWv1sUcdzf3qW7NYfYmv8Y6FxpIpZlOVDY1lNPwetUWK4AhQG+NlTALVy4yAc+
q/Z+exGbbe9fRS4W7OqquiFnqKnIAmScJBbQWzmDvQNmYx6uhuNRp807wpgHQjwLq0u8UB85BaIy
Rw7nLUFMqZ5UMdRN1vgTyhBjWzZZEAFSAAV61xtaEujNA5uKSa/L9hNc2k8gB9GUPLGPKIhFdlLi
bR17TZ7oZcrC//2rA0vUdx+t4DJ6YOdLvI64LMo7nn5vfv527q6w5Ac0X21jgXur887naDG1jPOw
ef3XRZNKdqCbfc3zsdZjIRidCzVcZyGM2SgNsFNJ0jhNxUAd/88QgFVoUMDkKoYLWjFfm9kSQhqy
c1/Hohf048sIMzqSq0+DyVnZXEE/O0CS4tqfaCZUIFs+tLq/Vtz3PQ3/zZYZR8NBSgu7kRu6nWTF
87nEfaVtUfDb85R4XrKyuiV+VufBIp5Nj1D353sqjql6vPwFxYw60xXKGI1HsdfyeubCB3pIJuup
68jb9eyBeotkQurCzCZ86ZoSWNsGljEo1y5UWWIwHz38R9ivV3i1svIzwnYz4bOow9c3Ysh2cz/N
nevpzfNwnZ7XDv7SDWNoRc2bNNOWA7zN+eFXM/zpsVdfLab6yzSNRlHtp/1wqi23PwCy/Dxe3RXJ
4P9U3sNvo/gBIIH1GqUmPThVjZ6VN2u7uvH3ztw1bekH+gYVlJppq5wG4VQea2WbT2WMkZdPsZE/
TebLJGNoui3CeySXXzvW8mnEbSFi87F65OVLUF+yqINRLLyynDx9kIysIiParINQMDFOiXvGTNQi
R/5SpZbRqyiBanK76tUYtUNlR6cse8LQ2kCBiFeBQHQhNjCUWQcVGK043EjvKloUefXxlzc2a5EQ
2RXVGaJQRLzrRhoQrvEkyfIqzBJZCxIgwiqPtt0GmhrvXUyYaujitTePAllNE22nmEQwqYAVPJRJ
n3L9xHoYuF4b+ZL6J0SfN6Zq0qfrjOUIQPaF4lgisGi1EGPD1hYse8gz2RH6MaAm4UX4v+2OTbNP
F1KC1kZVCkOmqbK45/wJWk3N6ioJ2hMzh/cVrD2OMqS0xzefOgB+89spmOXQpiJ+T51InyTrDgUJ
U4HWj6SFH8mG/mWsHieN6lm84tUzxaaN0TOXtEbkOjiDW7abtjMfeuvUicVA4fuEQSr7Q8pE/mhB
VapJOlNXZiCsXNeU9bcYV3ujQ8FJ9TOIfOEc6w3BfSfkyRz+FKayE7RYxZxM/z753zjjLRCIjUlO
O8NtOsm03+BCE1VFBdEGJFNzlujln5qgQSAwQsRbQ2r1KXof+JPNoM9EbE57aNyu/crW5iH6lG8j
9IqVlk25kfacvBmjjLJj2eiX27aLzVKK5em9z4GI3pzA/5cC4Y6BFcfO6hHG0u7EXR+epT1UcZ/G
5JNJUpYIlFxPvPlZxh5mvKTZAkfqa7LMA7sg5rpbxFQtyiQrJypQaXxMtaKOV8CJIk6I9WMzWRAm
qiQ+ZPFWnJ0Sfo5ofMXpE9K3biOpwQwnFT6/xfiJLyowo5B9cTzKEv6uUzL31haUwOmoSApMrjx0
fueAHgXYRc+/J9SMDXt7C2jLeu/SZ0eeGORWge/A2cS8MnIjAQAEV91VewBHc5xY08MRUVu/b6tV
vsGjV4NQo/NTrF04CV0kwAOdB9Xvw1Dci6Uo3YJYbuMFs/fQTosN34qfs82tcCa0zUc6E9DZ0Gfw
GoaGuTJR+XN/Q9xJzjCHwryXjcV3Emhhwqqp/vUypCcdHUxLqSYqnWTWoHQB6Y8vYCWh+LU9PJZA
1ZOSiFacPvGN2YitBj1wLp1jLkGAxLa4bcwFsS8NB1I8337JKRb309hD2bBTz7ZEx64QCUzEiYwS
qIOYhiVXZi4VrmunLIw5Jy4mVS3FSe066TJcgghsLRjB6tCXh6B7Iaa8EUJUBOZ4334EpyoGIM0W
O+PCC8bE7ZkhhDV9iPVXfZ8DGnVaUKkPadbo4hoVG8gqwgqScik6u6aIF8/Q7K3/gTEIrfW2NW75
QzSZhEYw+Uak3BdxWnjYRVBBHt+jasRiQHz9YpKFtnR4Q7rqJYw8E/BmIFiMgXS+/9RDMeDYwAfD
M6jhYQJjW8EdnISymFtInQHipYi0tMH0fkvFHjnHIbqtka80WARUbY3lRNcgdxuBkWMkjYkmIBlH
ca0a54b7FD4THNHD2d5EeLfthbEwcN3Mwcp2o3anBbvKtsONbled+H/jCbQxMGL1SrjawBGeFkCC
lbTvIIW3rl2fkjdP4/JbNnaIpo6lh+qd5XeTQdi3lsudc0+Sfn/WNS/DPmoOQ1bVjil6hSw79XKZ
29cj6DxhbXMDvYnDfT55YzF5txCbbx9CM9jN0cxAwXKS+KuXP1NBTkddTAJ1XiDURiq1KKzmoLj/
CBIIqpL/WxEW3hyH92UczAfxPK09stqLY8xyWw6edig3oyE1h+XvAVxGcK/SvCke8wM54PcKao2d
VgzfFMe+8M4xInsjt6nlvOxO1xwUgjCr71XgdgUWDfOyUnvVUwbu2nx45QaySNYq2X4T1ZSJTVj0
TtVA87/G1yAqls9Xw2RPPFBsGlqURo6oXto74wCEM1Ei3p/9IbphQ2sgNbV/q6fh1vyvA6fp0ZF/
FRL7KiFlwHGn7S1MQqP6wYIOkWLzBDSJNMVj6E0Nt0tlcnila+lCo1WVd/C3usv33q68KqL8o0da
RqmLCnpF96fKAojWB0xhf3LPwzUVKAw1eNYPplNroFFYn/DlacIpOkqrXgLuW4/pv3PW4PDkRG6e
EzE5RrDPBk8XBIlY/1gfPCBpxXBqvDPEght24zlNp4L7izBhUF2fxS3fjsetgGUn2sikFzrLM9mE
jsj3qFBvTs3GgQoLfGCLXYIEsE0+nBiCVvYUOcbn7RmG7UYTWFOY/jd5hhB0u+FBiWK/Pm+ZYCXA
OglZtteYHMG0+TuMkM87d7rlLOHJkueV8z70Un9RrTH7zRy03weUn3UeAMpY28iK23I59R1tfqTR
VyJh+owXJhGZFVlS10eCF12E4AlK/zYokCxVqevMeCA0uavTagKIbYVJuzFmL4t/cvRc9pClSchm
/6FR0CzY2VQxh6OiRuSoscYpktL/U8SoWoQrrWlk+MKDmmFsV3uGIZ1gO7yDjA0YkLbToyslt42+
Lx6HGTu4xS/VLoWLJxOm8x1wQInVMbpnbr702gfsUIQejTaCMF6Ch/CmyDntYlALpJueIzg2QAPc
xAL3qN6zrw9YmFApZdUaI+BX8Qf06vp4rO67/CZKc8ISygjfurng39eAETxQM+H2uzqp/gXBx3SQ
PfTvPm7Qx9SRj7ij2ok+yLqazD5Bo2hAMkROUudE2aCEkSrCHSfFDhHZAmGOPnZQuOznbWC1HVwb
jpUg/dv0RheyaFewhaw6WEyPQPmv7jyimjpAKxCimSBICzh1NpD1ISE9MB444HjpZ1Xmco7IRGtb
VJ42ENTPnEIzhLarcDu4XnbuGjASvIrVD37CG6LZGhR23mv7vpUysj8lH1S9T+XFdXVCjQPGvjYi
CVMeY/71V5oVuIsWPUDbSc0aBlZIIhRVKXYLYLQinYxp8uuLPwTmJ/Qli8WYnXYcP/+PUQ3Yoyyl
cbEhDcSTO37gYVEguCMp66S548WSjcI05ddquTHxHYc0EMFqTsaZdWaNtpUcrt9Kkb9cvFB0eeOd
raNnsWCODNNjM+Y8UdaqcR66g01TKEA38WgDB2JSKOe5+El5lLP2+eZfzohWAeZy423ov10ZhI66
k/8Zll5IT401DBnDe+upQ7nANlvY75eAZDc5xvKUnanlQ+7CXWItVFN0CB0QZ2FcyoBxHLW9F2QA
F/APpSZ3jYdeVYBeCBtjsgwp0l3TmLOpWWuWDS3sGbv9wojFl7IYUtKBgxUGGL0i55m+FciUxaST
0TEF4ivXMXWu43dN3OqLT8CaGZ2lzLTb2ZpCDawTUE+YY1Wjnl+Db76XjY68FXPPrQ7po7V4jmeW
qOuFX9q+G2f1lbG80ctPsYy/zO5duSHc1EIp/8E9miaKi+00wIDWVzmzJJffZ/W1jzAcAheWhu90
/aBcKvOBeNTiotRtjMphQPqpzO5jaWOjkTTN6MJFqx+7nHv4GUdB4PAUhHRsb5NSiwtxXgErRju+
CwZcv3ckATFQWjuHj9k87+x4QSEUDDDPoVPpuT/rhi6c053HAGo51tQGD/hU9F8tNSLW/GU/FEqL
1ZP7J/9R2DkGdPHVrwKWMzxxDyfOG245idKrueccMWLenaNz9rNe0HYb6nmmb8hHm3rplrh1Xwhc
zPutwSPwWGwkX3wJWyxr5D4t1B0KGwes0MiE2D6Jt7iFBHEeUkfbC3CcOxRUImDDXS9jpyyrWKqJ
g5RPtjakfR6eWjRG377IAPE4S6QkIiF+XlfnKuZjaFx8dQw0uYThgCUoG/NEG2IQt3nXvyxx9/Xi
tUoAOsgnxUyQqwB+0eDKUbOllD89/aKAKuJj1g7YUAey+5MYbSAkrWs9rYIESylJf9PWqhOEj3dK
lwG+Bd+wkXnOu8016oeWh0LeSEWrilDuP0jUIat0ycIAGD7MxhHO3w6EVK9pLiJxZ+x5cafJDWAd
3ZehR3SFhwYATBI8x5RXLKIvUFO1Xe/Mlw+uT350lbvtnvEEzDZ4hoonxXAxYG2m7JqGvC25xRlc
RyxMeQ61APx9ZmbJpuY0uaKd9+ws0ekEhwzIsTnlEPL2lQdHvVW6mLqSpndC44xbioJivvos+Wgi
5eXfkbFpg1XrW0euKvB42BR2nvIH6DQbSDBPKoZ5ug2hqgEccdZ6zZMj/1GYZmUl00Uu6tQAbCQM
RKciOYFDhFkP4YPiy+bnEGHVSjSGyf7KHm1nPD89eI0OCMj1UuVpepLqNI2dfNtQHCcklSjFs6G0
NHou91rEd4G/zktiiITHTCJ2T/THs9qaBB1U1Xn4UJGHYPbpUVDScIUklQHMhu+50Rlv4GUr4KJr
RW1l4JsPMykGc9AQ/gsUBpXDkYMqaREIHWC1JmgtP3znXMNaEX10/7F+26khOjb8tY/bYckRnou0
P9HpN171v/L4gxgqaC2y/MIS9gHCPHtlhLc/y//H3LQVyqx6IyuD3GwrgF8g0NqISIiMf/clmubI
u8LB+fmTYbg0gmUChMvVrDJmrFetL3nwnIqMBIe5PiB5chy64w3hK2jqWSx+z9f6bvk7fCzyUJ+v
/S5kxcrmNj3bpkpafPFwMVyHu7IPtYrc6RR06wPhdawNaG2Mf2XaS6tIp6hIyC9VBOlMgi5Xacta
EinnbjRYpOadZNa9cMEsZCWhNXnt5UTYyyg+2wdu9RGT6z8oSOy6uUZVEPmHePXN+X7lyje60vHp
pYeHu0pei87hClKb4bqZRGMdSLkKCGgaftXPGt+pPYNF58vB3kUVyeF5JyJ9ob6AlQiPmHpeh6A0
hUX52LJuNwugiZBuCQCVTQ2goBWMajwIuVhobiHeg41dCbqKvx8DH2LbHyGQlqoTWYT3DpQdMWmQ
EMg4vP9hK1qi6HgoKsXzDJ5SyTqWVC0L81ixuz7nlm0SIoUS1JyKf6G1of0HcbjSdcr4ow1PcwyC
keM+s4TAv3G3RT+44DAS0oWOoTy1lTye2vLcgqCWsx0gh9UkhubNlbLyp4Z3wEjQtoD94loC9tOh
JBhVvy5b52Q1HHymPuL323Gd/JPAE8waSP+RgPfSFmkeP1BA+ZqyOXw8ReeBT8fJozBRsK4EjMhW
XbbTO9iu8msLFw9lRRWQcW4zZ9zyJuQ0pAoF68zMLg/5aB/x43xLYlYFqZBOn3Z1a83xbMx/RnDP
PnyGrHC8wnqpoZ3GfNo0qt4hDPwdCRkHv0RN3CkVD+nZBDCPU7MfQtyzhmaTer2RxSCHV/AMZEyL
SC/LvlrH075DIKZs+Dkrn2B+mXjGkD1FwHfr+IKzdfyCD+hwIdZQ00lmcQcsZCMhoAvFOPOnlTEG
a8RGGbyFD9QMIp6CdASWGnlFVLHXxUfI/6pwwvinyYfwgVjHY/pkMksh3TUyqdUb3GQaydTfycpG
TScnaVfbKm8lapF88txP2HiQst4xif20TDcvlW3cCf7DPb1El19EH+lffavw9FTVktIwEd4ctuOK
HbzGMffJug3RvvDRHkpdDfIAcITtp9Nh94v5NT1axnhXOFQKMgLIls65fHwISyWllhiH51csXgSp
3zOTSBCjGFp8lfdi5uR2f+P50Lg1RjRwYgxXXduai1qvag1ZYsqm8F0gnQHowsZr0G3M9jG8nTec
aS+bnK0sV6UoSv56pjLxL4xnL49iZPN+2130wfuxW8gSF58HADYYAwvKziAOwSJAmO6S66diEgpu
LgF3BOaAURDDKRsOxCbo7VjGSWcp8gA3WWYkuhbcSn/4XNrtjD7vQCIL905xJnVSv/lOBQR5TTsy
70vYjp2Rvz/iJIF5h+UiwwZ0a3h0Cd5TTInZAcImckh/Ytn6paC2lFY/AlndfdTdd6hRkYjn5vEa
ufya8x2Rz8d8tw5mADDTV2pHkSFHMzY5oEDt6wJMAvqxH14aLR/OSPVPRpeL+vo7Ny8eYPjxRb8j
U/8Htd7OX9HdsPJ6a+8jRI1RB69GK9fBfddknaBMuMSRFXXYSEBiOLCqYldvaMg8oMXzXOboaRBb
jjaiZnBemFGga1CtsaKKzRu1QspcvzpP74taGET5YHRNSRBB9oCZ6lR/PAl0Uavg5e+nsqRkTVIw
ti5Ae9FoOGElxBMiKpkBLJ/zcKReG9fjnn6NeDBi0uinOJ2aPMM4OwJj5u1Ev0nGg1ef/xAO+lwY
eqWgvMMxi90ekVABEmzNwGdL0QkSFniAGAoUbEfXl0ejHm7VXt42/dEgUnWZpz/xq2BjaRKOFUWr
FqedKU38hnDoMWoQazk3mXfj8Wk9/XwUqn//XviDgJMyNYBgP++SHiQMbkXwoNuGOjEo8JRMyGc5
BCa7kmLRG50RDDcb7+PRmJdQw8/xwAOf4XQkudKabe/6NZwJ49K8HkWxmSMG7MNSQuokZo4x3pGq
jBFI8mo9AIlfMLd7gVR2JY+WurnCsQz7nmtLYLkDWHN5jzGLwzHkP9kGdFWQyFV7mfl2Uga9HefZ
Va4bHa23ljEZRq6/3uaQwLKFj4Dq+I5b9knU2gBlP2d+JonNTIBpGcbDh+sP1fEZUUruERQ48T2q
Q8RkPspO+kXuvA9KnUZaBWKmfdFm3t0JnNT98hwREU9ih28ZYCE7+zMOAwuqUHYy/UKdV73v0aW2
kUBBee+bVH1mE+WGNpI8bKK6q41GTThjsIN5aFzLIQhNbU5TpJRuXqRI+WmwoPTgRHKAAbEmm0Zi
ySGgJOh3WrUhn1aWkcS4maPf1MlpHae3Q1v+Q4driOHyQ9B7fVEvhI5I+F5twVn5llIEI5jGnyHH
6y8B3KyZ3UUFkZJrr8Ur9o3pSYwpr9pObnAVkA4YCUiL40eO63JnsA2nC0JDgQx9TCgckUlKtveY
nFTUD/aP493i8l77UOONXFPuBp3AbFvWY1hGmpNmhLd1x+7VZMyLiLBEe3CZ0ayrFLzPO+6wkiVh
CMvJ0RLKuVd/ZQoSOMguLuCkUrr6XsjORAtgiQO0sokabs4m4BcOw+qKwdZDsYJ+oyfcY5hbyqMU
W+/jYQZnmpCDEHDU39EvLFy4vzslQXm5kPG9AYBcITiQk4b6JKZ8MVBzt3WaqQhni+YvyeR9TQM1
5ylr85zc3H2COQucB4BLQIzMt3LNCxUTwDYbymfX1J90Uv24jXutiJ5flTfwZyydiaSqqkA7Yw1o
3lXlr3gBX3Q/5lpD/j3rLWp6dHlgvTI7e7PbVlfXuUZiLbMFDNj14B527Bf9xrt/bwyQ8UOItP2G
JmeGzK4y+taAyUnshJS/JjyYWS5zI+ApKzEBHUmQtoiUu5uC+G9sqYCHBMStGL2UYii1u3JIwK9p
9104rZV4FFcGhvOEWb7JaSptBlOKq7y56Ao8Snm0TQQ72s+6368KHJxf43QkcenOZVdZf2p3ufcB
rOjrx3tHz9KVbRPaNnWe/Y05CCP6oECExCwpZUeSo+pCmnLbzyreQbJByqp1XWNAaufqz7AMvtV+
oEL0WCoqKVqIVZFHH3hHp4aRUFScMq2rzrui3rW/CYV9wwCNMmfeGCRJpTqprx02E3zpAcsG8Q9v
wpIJ7h+ofEfH0IU6DHQHCjFavl2+ciO60MnRXIF+sjvbkP31v+ATtV+vW0Weeqhq1AD+tOi4SUZm
4J8xQWyARyTTfpBv7csBTfzo7x94JlAXYo9CSdhu/Hd6c3j9+2RFOkAdDxqDxYMzhxnyBi+TQ7dX
AbAOwOWYgpUpIoRMhh81TkF3adLwtb45xDeL6GZPBnabrdKeyI3zhVVk1Dr3IK5KmiGVjCp4ker9
QvVj5FBOz4ll9oRqxCys+0VbK+Zc/yBjcilldwtVj/WFlhvPHxfUsMpkMVdf47UXkTDniyvi3wEN
9F2UzXHRrBsjtL9VijjKJXkaHNNxdYdUOsDeTtFNyLW1gk3ykVN1ofHwO0MqmaixMh9rJC5L/vzx
TRHDMa2Mzc7qIXNqVh4NZbs93PDhq+sMHKEFhdMFLpKFfrysyQwGaL8uTpKX62bTQHmTbWJpvA0d
QWxCRCm2DkJawx0DLfPJyqHWygpG1yDmQT8uREyFUdR76tgdvLgYGT8j26qHgHbNqDVdF1bKvhfX
1yacod0j6ngyNAjWLrCV+AHkmMzGiLEjfVXBgvE2f+AjBuBHR/KFqJyzpHzi1sYeCvc63NnEn9MP
tQV2x0kEuFb+GamZ+pF/AAmNsEiskHNLHpo28eOOkUt78925pdGPjyqFUfdN2t0Jdy5p5N5yJz2X
DgbOHOUyt5JQ6llgQ2Sxy03CY69SBEkLldKE7RP9bT6plhX1W7yQG0jjzwyb+i7l3RGfazfy2+iT
p9xhPa6H8+Ny4zGyvtXy8WNBVMKlxcftX6Id4eN7EawogOrSu4UbZrOU5tP/Zu0FeHSlI936bqvE
fcUOFtfN6Z8yt+PSb7hRxbm31Uz33hQEEmXntyMjdiYT4uyd/uvsFGGI+wFVUZZ3ln/4g0L9iXMo
Ti7tYc/a67cXkjznJtq7IBLVhHqHZYZZe/wojh5gM6dnzVwhPCY9Rb2YfqDRDwnOJjsErS8Esgo7
9SUu7jza/z7GAx+AeFZ02E1g+gp389O/y64IMahevxztJ4bWUXBs1SOXwO1jeRB540MCBWbSL1Uj
ahd51a+ZgsOM8KaNckn1gcWkNf/346Jim95RnCMjbYKIovxDkjTCviUS09rrIEly5VzkEh+XRKYN
n4b4sesNYAHk6RRC16NpCBfFfU9rZ52Pwd34QjX4K6zhxlVKh5xG9x7Yfr6Kv/1O6MQqJ57XruFU
2N3I4z56VyR6GGUAdLF6xtoxwpQDp0FGF8ImfiAK9qbN5ANsMtIecjEfhrCNXXlYx5dPvzXTfILI
KiuvBPcryyUL3+Qq3Hzv8H/JxXCd9mchwVB+bbBNoVgjXjuwpVJZDCh5HOH9HSNnZiM9dpWP8O39
CbDYjWHtosyagb7JMvvl3jkmEVWxnFc+FK2gN7Mn18BaeVW/g8acRsVv/ebivs6OdHEEsvFIU+cv
O6kjPXDDPWYyC7f930rX+J7RcAjxPr/Otkhl5bzN0D18gSjpUPxHAIgs/bgPVJmm8VJcVKVHmInb
jBar6lG+6T2G0hb5D38rTnu+9yi1GtiqywOdnqP1rjZcz6yD1MWx/85lFtNUkNbl6OsLCUMQf9hB
GRSif6guJmqgPh+enu9nfsLK2r9xZrTtWmTaW0tz1uYKxaJ1e0G2zk+60hM/HKPz8jjWn+teohS3
MzqIhmEYDK0wvUbGDlIXyQK3yBObCLlgA4CYqXiglCOmLwpMCRbuOO5QVYllQ3wajIXCqwLPLwfV
n+GJpFHrRlPyUTe+uA+x9wGLcVuET9+DD/gpXB9NWVUKr/dvjJjnhQQBXK4Xrp97TsqFI5X66tN7
8PZJ1sl+/0LVHX0jF9iYpH699E0K6ssqSzXnQA6v4qZfra/rrucOPSYsTX+BCquMHhjsoKiGuZwq
Y09jyziTeRMa9FcIArmEuNsfHhtw0JK/NxtYCz9+7dFO9GZzbiEKVNk8Kj3MCaWkUhhN8K3uyfLt
ByWTeR0Irl/ahQ3/+XBr75SmzTjAtlNj3fFj3QwoWG6HEeQjhuubdRRU5KJytAhk5K4m3C/FcR4Q
76EaL9WTzJx88SepFrQ2WAaQmh8TLWuhuhsHJcwJiWCKp0XAoCUf5IhaXALpuH+twQLQed2WVei6
UOwgL9zUD2W7DZwuLeHCgYOXuuIZ3+loFB+JTYQZrL1+VBBQxmeZJpmyhKT5KOomKKCiYF3yZ+/1
eMbva/BwuTdVWcb/x8sqMHVTnJHDIWYExUHUED0JgudyaeWv1UfIfCbHlrkPziEOFyD6WjGzACmo
EHRRBwCwhp1X3/IfyJ9Rth868aZat2An7NHJsmmD4d323mE23zkL0jbHB9Q5mZJP62HUZRSKOra2
GGzNJBu8/jjOBn9gR2v3dKeNykwoie3LEakTVpphlZ2Mg098HQx7P2dGk9WrdlaS1dU+xyZBEM0q
GdrBsUoJ29GQZjjrhQxl5TqlPSCOFad46GcAWMaAzz0qIAz4eT/NzaphMh20xaG14kwLVOwCiBTV
/g8uriISVekwKgUnUlTDF9XuZSiqWNJa6igd+y1ziXX2UlWPu2aWGUrkUbjCyl8JTpQqGmQ7aV4u
2BPvPujnAPGWNT6jjiZ6ELTu7uO9iS4tnaMshqvxhB0UA1N7gutldI+SoTsW1IB3tS0Vk2Vxlh4a
KjwxDdU5qIwYYD471QuXncvUYkL/sok6la8QyAxFZFiDlnR64rCveaJO1+4qmyypNKRfLKwzgEuG
LiXRupXScSILc9MWRPeZAKdPkuUnUehIWAAXco6LSCsxPqxNMI0Uoe1B1OJkLkT1/S2P5cO+LOsM
7MvvavMdWG829LVAJF5VLTzdAuvHBNfMahD0Bv5TGRe8ExFfZwh7SQ1FDmB/YEo5UuNUPt7uzVYO
VzwgYNvF9iEb1F2/1jLwHruoHGHaTCF8OFkXwfi7vQrI00rItQ4hLqghr4SErGNcIiTXxFXNgobt
NHLRJk5ne0vwFmRRf2EkxglVZCm+ZpDPzO5pEzaKBsRitcGnd75cERbHDd0sFDpm+k0qX6n8s6rM
xq3Xnp+su8n/Vl7bq2sgwOLcNIhRR1lWcStBqEEYgR8ilJnk7DMDfyVfLA68RQQtdkSHikVm6+gX
g2ZgXMlQcMOrkJPbUFZc/vgr+CIE+j7CIP9HTw0aGiCz8pFXY/RcNQvzrWUkmNyFQ+lIHjZEddp7
LHgA4Hcv6LnOMGBj1n+MwLSJUSg9siTt8CjPOarJxlOxDfAwZ721Ad7SqL2ufakg7sZyiEbEeDhT
vMOA3cWtZDUytOPHNR9ZH+VBSz038edQtw0//jePRysX4G2IjGoaFtPD3qHHL/YyPGJu05b8qTM9
m2QMQ4IYqPWlrMClH8L/+PClKqYtrVcmGhSQCxIh1j1GZpZ6IU+WkPjZeEPY2j+dSaixhiOpGREp
7tz8+HFpyDHPhUllXse5SBnN0UeuG56vFC/KdWxOIR/XuoPQE4TDqVRIDuEblHAbdrVV838LCFlX
oozIAdIuN5PZXCTfC4mYKQC508xjvddeowPfBn91wIjMaSRL8cVAUx7LEBe1FxQ2r/zTJXdz1q1p
LIuiWALMcwMw7hw6guSti97xpjmutjl8jzIz+E437j1pGHbl23LdVHqK5mfzhLiiONcKcgUMRh4O
uivYFdz6Gwt3CqkfZD+JjLUlhevYx+pTBQ4kPwnMC6nZweBHgEfRIgYPb3JWtEb2uVH9VTI/zWQa
PHPvINWCrrTxxebbPf/OSBMtarX3n5oRVAKy8B85tPLy+Ci81aqEeEUpzt0eAxl7u09HB4uanuOI
YtdBmtrWW85mRwuox2WpgprlERJpdMLJ8SwlER2/iCUqn9DVW1FL9Yybc4pqDhhKisD430EGQCZu
yJwc4/jNmQ4GIafjQK9tKo1y3fYB5dleXqEc0fFzYt69bryuIIb9mfLQRWKJaxvjV07XkWcp83si
sa7f89h4W9r4G//MXzY8D8qftkQPQFpOr4/VYV4oZRIeCUo5ayioR+aZuRPs5EwcOVaXOFYsaVVY
INaKZTsutIWgp/ftGiHEPe7XV2obN6n/pN7/QtgPqWr8N6iDCGYv5DCE7z95u50X4qaDDqiT5cHA
ERWSG0PknBdzJdYOzwM5ytumrQu07myfzXu3svxHaidNcIhOgQnftexPaFCtGnZAsfTIZrxhIXCK
YPXLPWgbEyH8ZfZiW1DeQAwe+sD+kCrtiXY9uRoSXvEUpxjpeZPWvoAfEo/QreL8SJm7Cg5YvE9B
TKCWfs0Kjtc7JRcNQHxF4aqUQVxPlLN4CNgeRqc1rz8cgmTHmZKUj9oc1Yppogj8t2jhCNMQFliN
4w6SN9i+Xzhr+gtWt7a85/S+8OOCH8aiOzOcf0UC9b4gTcmdde60vXv1BrOOj+NgplhxUwQAehFX
rC86IK9z+1NEVgoU3T/FUxhEU49vlcWPKRUkJwDxBpqhbTJPPhgJLU0lq2Mn16hji/+rElCglLW+
fRGodaYZHFTnjYyYXiIAKBDGX1Ru1YYcy5jnkp80tRHyGjlbijZAvDn7Jg/eQlf/ej/z+uihYhA4
R0ByEG00w96bbzLW+jz9nyFN4nf4+dRTmXeRH89K3/6vRo6fH4AYUIXFA+5VZe5HqCNwJDLPanAe
2Xp3K5AkS6BUQHmXu3DMkm6s/j/euGpRrRkbYIIpIqVaX7wTzfXRmmqiihYLc9xc2f3jyeSHV9be
frWK1dEjrf+N4LnVDP8BAPxB6phA52zVbEzjyqBbHSKcKAGmtiNuOJJZZ2ri7sj0X1qWxWO9Sgl9
cpTJ8xzlsIHW/LI+abV/oAAkatba+aDRd3COo8g7sDjDDKdLsLiKg0zTimy1DZEghPMCz4JhA/52
vqKJu5gTXau2Jtg9+MxqLr8IvGtlTyNIzDX4yfsG9SGkr6i3iAlLRRzLy4o6i/xJIgroYyStGfVC
tcNZKF22ZVaG2pQ1bJR0AE/qf+RWdgMfvoNYL/ofoJpKbtmg8dFNbN3Y+yvqDs2x/OQ5QnY4JyTq
szJsig/urY8RT8JBA7ZnYYeVIHkEE0Eg0sRWQB4VzUv/3K9UVMhPtia/n6AzYQuRh/DktSmQpXmr
tsgmE/WHHrRdtOexc3pb+Xh53OQdSEuxlyszYq/sOF7XBI/ZNzHRMqL/aeeHIOWqu5Wjf7HhGpGO
N5EhSqv0b+lzs9BvuflWFqS8lPUrujoAMcCWTpdZopHlDhl++GxSzZm3GB3EEwxp/YvyAEv65Ytm
wfkxFMywiZAWUIa+LP6QWefELcL0E1DE3X5OVPv0L119K/VAMDjFkBES+YRQdSTAKsSqcI7Mv6AQ
dArm1rsAv1q8fP3FSCET90eadB7qdq9xsYbUNP1c3jQjBcmnE3G+et1lgBzLYtrglBvK5vcm/KJD
sXgknl54vzwygh833Wz/B5E4UDAfzXPtIjvl4WxsUQyLGoiU16nEOAAQ17/AhL/WhfIQvmHTFYU9
j3lmmLlB9bg49cgDFZKqSL79OuvLQxBOoxwAeDkEgV/SSorbv0XXprmg5f6+aAYLef2JsqOOdKA+
5Pqn+2yt1kPVvo42V/0tywjYXKdJSOV4DcnBYSzLT8dIrvDSPrySEZnwXBUOccldjltT7vpy7Fk8
tpLUa6K3Y7BBM+ZW69QG5aio7RZG18yZQBtaEeMLYNs0NQHDATqjC/HomiGYPDFFsbp1bWNEQV2h
b8gLYQO8dSN43vTujBnhYM27L2GJoT21ISGYmqYb/Lzlbzmp2xZiteKm4mv+Yw6YqCDvhvQpeeX9
eNwCDJV/HFyxygiR4q/r/ERdV1dsolEgzI2am2Nqu2SeoeSNpfc9423hb57ZidrRVh9P+ibcguAP
K5ueG8Mv40tebLbXItVayVmkTGtc/9MC2+4/6jKitYDBJZ4+dItsm/JwY+gbt+007/Lk8L02sK7W
T/4/k0BtcLakXytsN75KK2YyW4gbjTQcgh2xTAm/gEea0qmRgQ8wfqRAMG8XGbozSWSH7utnsPaW
m4tpEaA50627RnPYpO115ADAlaJAGLQS6XyTwdoSz7DOPEngN9Xhy2ombOMyEn74gYQ4ew3nGkHU
W8eJFQnwOJfsRJBfP4coQ8+tU/edoSD0Li1Sv8DpnwDGQjXHTPKh7QxsFoEKrlgjDaJDr+TU1PZk
vxmIoO7qBQNATw4E6ew+RrjlLSXJbqXJ0rUyPtQ/fkOqV/K6oWMehZfK/nRkNmEi7AcG3VLVggrp
pUytCVzfHQGR46Sza6xiuAvfLz+8xDNDius4eQirLr5rYwfhn4Wg3t+DJnNvSEw3EA1lnDPBuWJi
NOOWBfDCsNis89qCrdP/Z87yUxidAsM/9glefCeH18j8sxfHMVpcrrK9KWga2dO7Jz2G7hQ/IW2V
7ZvDJQj8fNTHa4UOYx9EkbaINmcfkIDlaFdQ4F65FHOPXOHN6n+RymfLzJwl+cQiY5kiR9h4TfsW
6e49bZ+W9sCuoFTBvjBS/Hn2M1yxAo1pcYdmOXk98bQFSiwIQ0LRdj/2giNFJT/nZ9fwUp7yNvIu
ph97aN1gfv9oMsDwALeN/KgslyloymtK2HOCoWTRUhlvYSVJSPlrW7b578k5vEiJmWDccWE+yav8
m2DIZGN8mGTrAwCdCFZcxMCs0aP/pR1AbyIVNsaxJA5EvFx/KXVFaR1b9Ly2xDhzGu/Ol2SnQMXo
SKFUVxHYV85AzydG0vD+6taI0XAihSLsrYf6a7rSvTMwWzZ2ASrBH9njooE86bvS8jIv/vCN0fPU
9K9AEjsSkdwT8vHzDAJBpjG1/8KLXBsOhcCZP4VFE9ACzktg2joImOadSX4Pio94A/GuGOPO74TP
EwKciSUjN2YerpZhbuEmUFFpV1XOaBTM2SR2b9Uk3QhntwllTPtQaT1kAL37+uQx8hUHLqmzMT+x
Pigs+LHjvxiSADAQsi98uXgjc+g2BNemNE+OJ1YBtbc4aRb1VtURRzQ4ymOzoN5ExP3RToiRS4vS
PaHUjZcWjt1bOGZo9iGwCNRo3jgjZuYFgPRGyMzqdMCfRqnqjpnFzEqyJnE80rj12+O8SMVBI+KB
HP9oGAGf/o/htfwMm8TKTBqktJZW6JnNhU6beDryqvL8lysGiV4aH4RN1HT0Yq+MohazBneHuMQj
ZojHY6DuZ9IeCaaey0+FDhApa6A1zktG5gGk6WEXcIuZu+MFN8TNjAo4aEGnOP04T6LpRcrBCpNO
AVhjSU8e3uVC3zV2ofSgvWJ63M43xAeKxkabH9Q3S70QswPE2HsqWGwCdLkYqRDz0rnPNKSPBHxc
QaIt6ZxSpvYQSz849zg3mlJ2xW0qusbIRqaHe02o7W/nQLrN/E5yxvAL14eOBnF9W3ZxxjxcX3ev
FljE+oUKuy8LePB0rib2kfNiownDfTGykU29F29TqNRxBWuiC0IIAccvLSyYtSN6hu2G06CYTBYM
w8EYz8tU41uMoLyCnfP2qVP8DZwW7QccSeg3U5E29mAWB782/S0cL571a2z+bsKTlZnactAkbGTi
dhwj3ZRKgBrAJs3swPMZI2NjMBMg6fd2lFUquIFJmggO6Ev6viMwiYLgnh8hCDHcYCeurk6bVDaq
hLHd+jZk4r+H2FzZwkAcJtYgP+h5QfMjnPNzOBD45AP4TN3nZgF2iny6XzXUVJQV9DDTb1ZcNmCQ
9AOKOqsDWd12Uvyw0cXdIwyen0qrvTlWFUIWeXdzrkWUVVKVXoBeZldXRCmIHh0OPgWosg4nF/PO
5QxZWUpVh893Cisz5ZZf5Ko0WSTc3PYwWjkLgmP/xVD0tu+zzY04Sl+WZrHgMQ45xPRQGJlhMeeN
ap31ZhAW4V1m72OPfqURjjpXJy5q9Ee7/Iij9W/mbLHilpLNHW0q+MEjkAZi2mDZ4tQ0/GJxxto4
qVuu4Abc13EQD7CXSAv8A4falq3IOJ1z7dRSMt4tLvYY6afOkBKasvmbPM3eX03GD2ITK6OWHHpQ
Pbmw23ETcNPNFAq2Ws4ogFEvfb7rgrsa0/2k0kKwHHSeddUh6Gc0WWDWtn6/boWQIRsRfDT8ok8q
oRBS0ZSe7wVrKv4/GoGQeB7pe4ctcJ2HSOOKtJ6bfICe2eqTlkiJDnOf+TbvH+pWHab7lVDMr6tB
uMCo7Pp6Nls3G9kRqYsdwhU0DuTdjzmrn6r4tntH/3sCVcyP0WwFrPN8pdVAb8hWkB4XBPXlJUIq
qw2GRPCyMwQaHwsB83p5aQ9ri4fBKTpk/SjIHYW4FaSlnxmyBinJP4l+iVfhZY2AjoAwuS4fZcFX
XidW+zdr017ZLQ2rXcOzR0xlCWGsSJVXl9hNAIi/hSP+Zn9EFL72YAYIT2zn2tgyWIRf7brbsSwh
Qjuf/uJX4L0cAi+214DL/viFf8xWO5wXsVAozkXSAk1aLqECScfnQxlrcXwib8t8zjC2z7wXJTGT
n+mNecY2nG3LYtMsopC0YR164DP0cPK3X5x75fKbZJCmg/7EYEnsVcEuf1wCrXfjgzKzFoOdV0g4
PlQ6SITd7zVXbRnOsXRoixeASNmMUUXkirohIYdIVowTSv1Mi/i7lXwem0sQJ4rjqb7keicsDYJ9
PQuI26rKGhP1EmXq3AjIjlCnQirOlDKxl9Yn03bagY3VLyKqe2pCcXZ3D2BGLkNvMyq6yhDiJ8if
Jsnibt3JDq5xGWkXCCD6wxloF/eN1EMYP2j4vtJnbrTvJAPexDxUs7VanGs6ZKxTT1XfIO7dWz52
bfIhxzJ7NQNJuK2S35rgmIE4kQBEtq7tE0yatjsH8uxaDwl/Tgkz5OFlBmF+7210UJiMzf1xZkdb
KxtYK15QmP0xfjVB+4FfvuFST3Ac38RvjD0jwYa7k8j+iJ+tpScfgm58wDgUdw0DYrCQ80hwGA0c
HzqrDnjaK3x3XhIDrcG8XS2LiSnKXwZrrVYges2hBve/AV3GnhHK1MQDA03IqidtCV1EY41/VlRE
0/+35veIR/pRPsmme1vBAZIqb7NoKenO2NNXl1Rg9zLpg9HcYM2jnlx6aGVdoq91h0SgEA7kNmRt
3nQl/X8tL+kMMx9uXqa38Na2t6jIZLdKgjU4TLjgjWXhNRFR8GV9oQLyNtSiAnYbHy7Er7J0jsYJ
InmFEIUbWQaL/oDBslshUn54HZX3Otn6Ey1qJLXy+mlqp92Q8BTp1Fcuk4AhqUdIMeYgPLcS4FJ0
rCyKS9o6ctA3k3NYxR8NAyyfT9W+DFV0eT3Jgmy2qP++Iht5uqWevdJnTa4qVHfkcfBUnigtYPY+
Ir7meuvCyF0srRAze0QcPghgbwGVb7/uCa1yLmIFPDYhvnKy6mVWjmJ16j3Pjbrdidex+LTD+xaR
gznRt5tiecgQzOSHwAQCO7wWa2/vuraRlLqPZU5OFSqDnwqkKDqY9RvQrErEQTcnafvEIosgn8vr
6YoU4X9vL0RcpLOiy/f4M/jB4vipxZkitq7GppLnt4IO/+NPk/xx0ULLt4D2Y5JW8LLRyyq67liE
VCetQG6QzvcIVg8ETWyv4BsDXanoWr44IG9N4+WMsUCq31wM+TrwOFGPdN4pG4v6N2+PBpbnh6JI
veBtJL4l9EjiOyW1Jz8BpsKKKvXp7n3fpYCBWgPA/zy9M0Nu6iVaTiJHEgRGc56jXQjHEWcISSvC
Fw+xXwTGJO8/WVxs1yT7MKLgKnIX26DIb8EWDtjvPDn6FKhXRWx564MnIWstusTH0VOVftCCmEgX
Md4sB7MSV/8lLRk4a/bi/vW1RNwpKhh1Hh6yyUn/OXjfpG40OoL6enCiCBXJ9S0TjVDDxEHJCttP
Fi8JWQlkNPTiEG7RbsSI6xj3uWir+4rBfBlRanH0LDo4AZn/uGRD8ykvCLYtPeXH0tNA+/vJCekl
o728dBITZR4VCsCPvsAleIA47ciOrA/jgVHORg/lHIdQwekvkHT0vS4vnvVGJIo9LE/UNlnR6+qB
QxeC9EeJGNNz4vgEa3e+df1n1Zrtfv+oTiVoh4cCbWPgG+ZrM8L4eo6e/ulu0sd4pnThUiPxa1ZU
TtRLTMs7ZWP9oAFBRLS/1US4agIkAXTHviSGQF73s2RxBRMS7tEXebgk77e//7Wlmlqj9dXlScTd
Nu8CCccOKCgRUT2Uxa4ZvtRdryHZ7JVY7SPwmMNfb/NWSO2AwY8SCVdlQTEixZ3qyxld9uIzfecR
32dTmVv9ts0UX5TdwyYgcPjlfLaGIp0nYOq+qS0kN2zKzOJpjw2dnYTrcmWuwS8ql5mfoD6D/fEn
sSXadQc8QoVee4IddxHkHJWEP0b+wADzV7fWfZ0yO/eJDjVU0Y0F7NvYWO8PlKI+ZtKycNXakgfJ
0MMPjjGef9DTZNEPLq4pI9DWe4agW6oBozSpUtXaFTjplDG+qlqmC9ax/ttoQTDGJTti4CtnKr9e
bu1oLtwKGwIvqbb0Qh2D8M7aOUvN9k9z2ye+mMg/tnOLE/BsvkTTmnJR7U2n5uvfRj7ugiCXXVS3
8Ejxlzr9EwtzI38WZVF57i31kwc5X9e2SQ1a53KpR3yid2qSaTjWxR5/M7eaqYzo6G8Pd4HWrtcl
JbTSAQjlLePO8XaBQvwv31jbOfvtJTVjQzxGfi5/LBixcLRo3dEf+tzBAA/AH3InNRuEOitSVmxZ
eoKZ6wzUCNSdvNUQsXlrE9KVaBlPZ2tlptGnEkwHvDsMfUls24hEuoFC3alRy72reeGOtGeW7Oes
FFg7nkXG1A76er1jTfjpM50C5iwRwP3ZW/ps4Ru40urtpKh9zTdsh7N3t7QRyrRNMiojHZB0/Tm8
G7yAtaY/T0rvOfM5O7LSwd8JqQ9rjck54orRNPJCTsyaUlM05HIyWSuWZZ6ctT+GN7guk+tXieag
TM0z3stp0H6jRkhk8/OHwv7tg1jC14g5I+rtJh/yF0dyCUVmF/UD85v32TBOqmd8z77Tom+XIn+m
eZ8scaeEHsGOplClmAIvT5D9tXaSKUdb5Ir0bH7G4HZ23dQrEMNLh5SJBghjxJL95gfHyPrGxSfj
2PB4ry9m7rEt+lrBz7xi7b2wx5rS2Qu8lLyFEcg7cX3MclJhOyEn+D4c4cpHZ3nBCRUA9P5VW3V2
rQye+O283anzAmDGU3NlN9SYuWhcbqMpgYmIUIBfhWhMnFyt+zA7uI+IDAzHCqyolCZVfgYhYOCz
FCAUA+Fb2CJtheVr+1bD1dYDEHlkMXsAC1z3GP+0uIfqcqqr4u41Kj8YHRqxog4pIqzg0nYPZaN7
K5nX06+tsorvscc1WpQZZDNw7I/El95mW1K8p6PB+H8uOyYvAHDXC8TmUabPlLWFN6kEY1sU5mhL
PY6EGunX6bM5bJHMIVI7yv0GPsPwhPN8l+m1pozawSJZHGFEw5qAN3B96MvYSeSDo1U8PyqWBrov
psv0jtE0sH1yYt8TGWAumLUbuQmfwa1MBvi7ukad2Y530Qiy3Sp8vzghSi+XtA99m4P0i4fYMoEY
DnUgMUTbr3ek1L0Vp5/wFb5N5tHc2PAWuMED8norowGRgOxeiS1UBOxPJEOHrTjfIPN/DF2oZygq
oxOhNN0Y3ifkPXdSNP57BHTbT9cPb5Bp25UwZqNAw4OrHeFRGS8Om+gkFADQheVhXJbu7oBDYxv8
XxP9I8R1sUZrvYfjh7FI76A9piGXOgZQ4Nm8BZYY7SLJCGa9cYhc+viDoC94zTgQsk+IGcd1gKtC
XcHYU4qUST05ax6lsEZGFRVxMEtb7R5T3wfgcnqdPSveXgHfMToZfe+mnY0OZi+jBU1Ylww/GnEg
sFs+NyNfZ6MaRmzxjbYETqQeCKbaeFRBRl5NAp0pj5NYXIVZdIs5wimoTctspedcA9vH3J96ZROk
E82F8j96i6vAV0WkjhKLeFqcMQx9nFPKmXZotH0UIzNTS5XBeCQuwuCxJZXaTEWGCqJketXmhzdo
1xhPFexzTMBFDv/JIZF9PdEuRsnLlpE0lNiZaXGxR65mBxhaT7n32sIshujifAHSU6ufY7E9sj8P
ddkPTEpZ/GN3TYGKlNNfcHUivBeRRMx/xoEWPcZ41CzFm0XbFlskCQ3LFApSqOENQyNANq0+wXPy
9mnc4pYEftZO5IVsu3OhMrGrfUfRU7Vel/uZ0LqKbjor37IlTCpioBSFx4UbNQe7foaOqPTxLpzw
B5FyWFwI5fQy00OigDKB1HK56OYZNLXfhnL0Gj0H4WsLxqfRWkyEu8Ov2LPFB7qS/m45iuuvs1Ah
8p1ZTGz/n8IFQ0WOBRt7E0nfmqu2T9bQbVExga7qPba6rGcJ51Wouagj62zVB9dZ/CZ4pE+gBrvb
ycAdLqNpg8ejP/4r/JqccffinKKrGx7BBtIvTqJp0pDkptAaupF2sYQbMR2wS9RdntV+ujkbKrxx
Wxheal+fueNgG035bbpsrO8CkK8CvenZ9bUVZ6hPaTmlNBGXEN0sEXzQW4BKfOmgpA1K/SCN4zz4
DOUY8l0L6qw4OR3QZtolXPb1orjyAaiFyQqfbgvO7muOS8PTDqT/BfLfWbW+Zlu73Xm9Z5Gxw1HU
BixJjQyIDg2MvR5vNLQI64NxZGwhiUahRb0Bf/H2Om3UZdlbCIFJuwzAk7JZpqefbJKsp8MdCHGi
+meplB13w4FWmjk0Ol+Enmt8RZrCfwKqGVsmcoeTqGrM0HcSMtYdGkl7V/YEvOKqL6GXdxvEejhT
WaXb+Y0fT5sgPTh9T+OXPMT8V7vMlWxnlXisuBi8GCImXz4NmGLX3nTUp32cgxcEw6gkpGzymAUg
/NHnWKrFpziQJiQ3MGdLahVMue9SrsYP5VGasBr/M1/n27LYuQFSDixthc6r35YW0o4xbA9JIKq9
1XoR7SNrfCPa1p4kF4cLAAwaPfinovJ0s3SLPlCwJxYDwVpelxr6mrOOI5IcfDFtdYFrdMIVUFqy
NqZHHQsWziuudHdwBlOROhg2202NjmmscczLgis34TSedSC7zEzYZbJjEaLR0otaulegwC2J7a1b
rG1R/eIurVyzvmlSZ0Kg+GQ2B2XtAnsc+NgmJzCGrBKftYNaToPYHG0P2qeZf7bKLltQL7FhIsM+
fZ1HEMgEt9roi4yH0KXHMhUK/xWiT2yQwfmTXNyiB369iq9PNtic5IQq3zqcmNTBjQq5lA7kbtx+
LYQ159aK2TfPoax2d2Rr51XKmNibewQB1z4lP9Rp46Cmm9n3bsGHthb+YKL+tzPl0qqwyJj86Lbf
xUFxlOo47MiQqVSaw7hu596zrsCwPKoS3+Vgcb4VEvTTnUVgiO5h2lvQdU5pbPxFGUiq2tGzAw5d
pisIA0PdvFKYa2WAWQ4mT457dlvTWLbxrcx0VuROpL+fUMHKOWykbtGQ6rN6FPw2RJi5Ndts2uFm
bBhoHNDvSFZQsZCL5F+1pVPylqkicAVrlJNP3XW6b+V0Paqjj6L309vXXH5G6SiiHGoxCLYnmOI/
Id7mKHxwzM769KvsFoj9yQeunK6oviw5R0T5a4P3C7MoX6AR4nM/7qa4a5aceMntXhu30GvPmavs
BCR7BmJaubTdpiEIL4Vfrr3lTC12irUNhWhDy3Zn5XPP43VJMaLUd+D0CuzME7I8ywMGuWZy81aT
mkPkeKHgVOV6GZPsZxE2Q0scw425BqUlBMXLjCHtMEN42s5yc1Ha7lN0XjO7OmqRE6L2icHhQlXI
hh8G2/hCiQ1ItEgrmROc22mHDrcghWlI73a4V858qtmewXreursgvXcKY6xDsYZPiGWGtSBmDNb7
WAhUaHFhO1yCSCM0XcMS0xvNu+oKTtE66o3Oo7gZt1pSu/0mQ5AGJ7tHjT1vdwb28roYWjhMPD//
MFxepFVgRNcbPvPk8VamtPo29WKxU6tL0HRN0iTmLTQdpsaPPI72wsykQxDxH6GkErEXdprL7kVX
gNYWUny1ZoEH8WZsfT1KZ8iSJ1U75DdT6d4CUCjBvx5pPycPlVaNTtjoaS2OFrjZ74s7+UJ5+kuu
e3gi2FHMGeJcyWbxk5sqTfLEnzoxyK25qBpccIEZdkoEdWamkZz5plcKRtOrNe9sbFPYxlvr4dtY
SyvkVD1zAoYD+M/nsWTLo7hhGHeifqhylzPM8+ge8OtTbbA1eFGp4/bGFO6/uLD7vExxN+d9Xi0R
A6EwsbAyG2BcBRVJ2cNHUIj2QqIQVCDGZFz5feKnOEU+vf9hKs/mS9HZooluKn6SxlWroQBi1IJc
fUhlISSa3/AHdCePxk+G2KuyGJ3QrIE2O9A6VXMSXeBQRInR/o6yI915JzCfBl5h9wJEPcCoQ7p+
2Jig0VFxWqck14iQLbV57418A28m5kgtapddub/6HYC+bvGL+fah0xGWApuBB57EFvW5wvlKr+t4
FsOJ+Ip/a1alqQUKprhL+dYFO4REAsl5ezrDuSmqlfx+htH2+Log0GgM3ac+KbzQBteiwQWh7FRG
MRD6y/YA+J5YHk3iLpIU+Ew57wAbqH03WarQDayv28pBD4TOpd5/9Z8NgqDh/O9u6JgxbmGbRgC+
612XSHm5hzivNsJoEOunSqdlj4om+24ja0uWwk7mYnuhmZp0R5upa+XYmgiVBHDasDL+0lYrkThI
r6BWDMhuo34NH2bs1TtWzJyq0xvUY2EnC86GAaB7R+HOxZeyl/isr7DuRL63wwYdL/0fSxa5eZ2M
r8CajXxjbpklsP3tXkxy8000aAgtux6t8WKcIhq15ud4HCzXkbLvCuDEiKmCClW5G2Tlw5ZPH4RF
j5qK+I+3DVfM5lfV2CMisrqYsBHPc2uJuZuKpMZ2dxENe5mD+kaUk2qMswan/Ktc4OuTCxOcNunr
UBVw9AXrRe7g/3XBplFMEZ1bnVxiv7uIADx2swm4+OL3yjzH3CP+ezaxIkR2nKO1aRoRuDNqexUU
FOWbvrK0rSlYszrV5FziU56N4RJmlodrWCHWYXF8g+vMmwLGL4VfjAK4g21rexfd1fa9+ffFBYEs
7zqyQObu3eqRgNG0kU14K4+vZVzzk3yL3nrYWNMIJV0vVJephViDCnswlflslbhHDxXt6zlVxWTr
YzQpjlx4JqYP5XmZ1T/N0KiNqlb5dbDh1rQfjelRi1kix/IuIsxOf+fwPXqfgyUsPCrN7xDN5fQM
smivxotZkwZO33U9l8wVfNdMJFZkAeryebIoSe28x2+xlevcTj+lqTbCb4GpC07/bCuZmAQbn7YJ
VK1hdRghLOjJn3+MrY3FqmiqC5BPiAra2iBtVKo+fkZIav6pG59J8IlP15+Y5/K9uSUPIhSBgvEF
WeMF/uksoekb9WxLca0K7EEi64yDkpY39rMIOv+seqtisn+wjqKUER50eiyFrq30HyafBe9rarBS
uYjjNdZk+h7Xgdyd82dGuQBvhKotVv3tkj6HVgXGnNT2MxcI3xt/jPw8CxrS7yp0voMqE86s6i1T
rG2XL8mwh3Vcx5G4wUA3sUxDUyITbWMSzHzH6qjFzCovhgXQ+rocA2TaA2CzPRz5UfM2cZrZSUnm
BIO4R9GmxFMqUPw/ngLzL0dbC9Bui8XiNGJsHpxmm7vjM7iQCNNmsvBDDwLqXr0BHlcOJIhB8hKy
XClkYgt4spbNyX4Ul27aRLmPavED8XWdQzj2eUaozkoOPw8YPIoNCMft5it2pyXH+KytWgm0Q9Sd
6LPhGary6PPbg9AXDkFhDWQGzfUi8voA6l/DNB7tjy08dOjj6C8IiSMcHsOSkD1m++SHsYn6GCvI
0Upw05BJVT7+vMX+wEtkGJ7aUm2skO4JogePiQPSFswqlaRC6+RN7+YKqlJUtdF7FlSXZJuokQhV
ck9oWXxxQMcnqWTemGGV65PTfHw/5ahUz9PEednuGn3rxWRWVtXFLp0OOnol9V4BHHN64ZZajP3o
oqHPRThsjOKnkrUGsIS+cSqKOlzkVBIJThL0dJSp1Ap/t9AvOs6BVD+3YEbkjiLs3pg6XU1YWqET
JJgFMYY9qdLI3of4azUiWuk0sYPDuSNX/dbbASPWdmKj/EbKrxGRh0vKzFXTtrqdmVvpkoqIo2Ue
3AJ7ISiXYohCUP1vGUCdfQFe9LUGi72aApe/bvjDJugx+Lnt+1daqHw0FBrFVQj9kEr94rISqunk
tXDJQqiqX/uOFRrQzOLhEOPgm9SojwbA/o9YN2uiZbSPHMgySzyGq8jv4CDfXjEE1L9Jc8I92IwL
ZeP0hkihZws33bNUbEhJjFtuNTQmUyU7C/NsFVO+rRx/veNZvSVaZGDmXzBH24Rc7xyjCmHnBYLO
tPdVmtDJrHbMgHqlqaJVQ6GhZbyL1P9CT0u7H1TMbQremUGGQuvk7lOrNsw1Vak8naRaQcpXAY3m
cPWq7jFvsSSQpdwgA4g3KT3V33azSYMS2/9aIwOlpD49f5H4yz0sE2JzhEmFbskvgzKN8NlRIpN+
/FtKywnAZKKyq+Suhbzjwb79t/4wLgf/i75kXnmbN9m5BxrqaFKWryvKyTz2C4ZOxK9nRzR0Avbj
EdqRjYUAj9/3UumxVkvj1hbYfx9NtEV703KOf612eFWzj5OxiFJVNkbuRLedc9xJ0igFMIKblNkT
H4ziNxv8TO3vAojSRRo+6jtF4j6Ws7kAvjFCL3ZAQ8XXPBrYWRYfP3+Yg5SuMrb0/cyke23mjtai
W99y7bjJUii+BUDc72+L12cYZN160caqxE8Tr0DuTahebFvg56/pVifntt9QcI5iE7yKrOP/mLdN
8f8NEIitNI4VdQEkzOhfuSSkjaBepbWJirtlXta/LUX8ZKHRrxIW64r1T/yMQxU0AflAb2Xsr56u
6g3mPry287EOC9eRZbAS/VvlTRw2oO2VhBLgW7tS2z0pF/H4eOaZUPDUNSdHWPanaEfCXxrJu+TC
9qYJi2+Pcks+hTBsyFl4cDQ2K/Yk3uiuLlHoOBkc8brm67kiVcsSx7572UTgkaI1RO4eQOxwxKnt
8Q4YkfEc6OWxQdwAyq3T/N6LWLmYGZynGI+npC9AnMAn5jsjTLsySriLht0YMHAzQuguXt6QCfXB
aHDFcjhRONA4hQAutnivAhYzTFeWixbao3mIN6nF53HOV64O34lUhu5jggPiu9mk1lkn4N25wRVE
GtDdbp2lxdyzmUSOoUUlHAJxtS3hYWD5cS2NVDVQ3mK0xdX998aCy1Wb4Bai30wwki84LmZmJMNC
kISGDfmLegJgzxPB571cqRmyI1+JfIV9XrTLre6BbTiYxraUYwwybs4tKXGrMqwYT/on+O5LPp3T
9hUGaF8ai3t4qmUF/xOghW2U86Qhm90JGmAzRGqDGmYZYhkWdmkIXgvBVv3r5j+R+tFJvJqlVvFy
J+Mcg0aefZIQAGuF7/EcQBHrilz63A2TBiTsGSZDR5HA+cAXSkWmUC3+Xb14iifOIPPAqGc87JAN
c4PjqLT/nGNjZT8xwchgNoyXyRFK08tgA/U28oobIZM+5Cr2NPU/9VpJ56xBWTZsGiu2grP/JAIh
Q2oexVuZ/Am1wOqla3q3omdHFpQ8no/XwNEN+g780ZRFWrYBnjdqfzYn79a7meSlkEAEs+YUorEM
LQw1KZ9xNgkgKDEOstyMNe55iPQdfS3MzQyDddP3n9OwYLd+hLw+v0WZVuITmLZ7xbMlTzsVnYLN
hTEaoQheHkFqfGw+6Tsgc/50dOUXcbFs8VycRTn+XAERPUM8bQ1sxbjjeOoN5e01Aix2qB0Kbds/
Hxyiloh/doDs7kGaM21YaNxsMM/A0nYECFwrov5EGqTvkzCcIdeWB/woPaJooU4HRA2bvnusnWiU
xRgoABCOGYZm/zgan7XvsovA7DHOoDq5M9hFeUn59jdiMT2rpY+7zth2uVlHhs9gJE9DxqooHKuf
xkDNDbQDGLGQP1S6rqmiJI+C1q1KvpqWC3BAHxh/tA+NTKNYjpAZixxhhe1zNhSry4aZBfF49tEn
q3a5mrIrwotxgJA40ZRhgF0PuQZtS8KQ6fISwgWOEuNQIP75QxTIXupw8aCKVi5iKy6qCH6NDBw1
0UHsuMy6s2UvdOM1GlYsZHOmLRGXs10RHu10rxFv+NtZiCTA9Oj8hUQaL7u1mnzmd8FwOkknvxWU
is6Q4erbyWVfO+4Orq7q2bhEwJnHlB2VARmx2QPX/7q0A9GAZjWmh9NKhsVwtv4H/mvWq9FZ9+62
1N3l1K4jwQAoaD77z/EfJ/FFb7fWkzV3G4NEO9DpWUjOzhWKrhu3Ci3WyYijAft27bkwjxcdU73M
RaCnm0Xw1wOdnZE9jMDS0td23OJIZzx3HSIUSk39DQ7RD4CYIsem134KstD9Fby0/wGvTHL6Qv2j
fmd4GlDnRC8CS98rWp6Homn0k1F7S4DH5hBchQD03upPu/GrMicYzSee15SagWyxTIhTj/2kRk6h
99tlgz0ZhZG+kNxZKZQIUwogyJDJcH7xdZHmhV6nyS5SOWNrKHJRXqXpFq6oS44+QkjXu4sMIVnk
hZ2TPhHN1UNa/HxYUTtX4jIpOInRYQwu1hvuLRy/jlqsK1cjxlEgCsgP/0dOpawUJA9+FpYX6JPP
qFToniCZoIRbN4q23o5zSHAn5z31Rcl9pw7DA2KmpTvekceixdpscH5plDI87XiO3PVNpTt9cN8m
y+hSgwSIW9WFbIb7VHab4XJEFn48LHXB/M1wvpoLrDs4uo1N3C8UjfJI2+FIiZGPWJopgqUc9ABQ
O1Ndnourg+JD20RaKE4xYGsVI6p5lCcuUp6nn/tW5vm8UyB7nTl1ibUqSnRiZ50FJljMfNKaINGe
TmXnGeuXuGPArQ18vokiIw8a2YfNbEse/Z8KgRfXNdYqN2ioLbQA3eJ3UHj8M1/mCwbSMapbT7Kc
3KwGuqcEaJYdJ4LO7YirVcv1NPYIg2EoHEF+uoZI9A+9LBCqmj+kp4UnIyj4RvrgoUVpy42cVPNw
0Uf0erN3eZVZNHvNxh08a29rqPOGX9c8dFPjhoZhLyfJWvB2KgXZ0Uu+k8+0lhklSO+z/vhMFbn1
8FuJFXTtpqnv2M2r98Ba+qnlT5aOA9Wp04AVt2XVuOas1HcITooZGJ1Slt8aAKsTmcWdUYIVkSD+
bzhnCKJWS4HGUFScw/A0iJsThz1cXWUVhAyxt0TdDvgm6TJlyHlG2hXNPTIiBlvO7ESVDD1M0Hml
TUkjyKpR1hmgZnXx2Hhnxoev9ex3iFUHeaVs1EkNpcPiIOO4lI+IuB1lr5Aj2FzCOO9prtjYLhkW
XvrwrRM6AfrAxlPT8t/U34dpTBNLHsG25HIt2jcQYWbwtiwVnEq1O/G61BYUMZVoLvUySGK9qoMD
+82PhdJ6jzFpyjEFAkfXCGatoqylI/iGtG1VClyoaZ5J5CySkHbjp5JJzBiQaxGTA5MV/zd+SqJu
PzxFTmVRH8tSzbyZ1kV2bSnLn29L8BiJ/xjwiwNMgQ7XXlKJ7iJaOyySKiKHUvgdtXBYCtIsDclk
XPopX/ROm1B2UA8aCsKZ4BU61fTmKxh3fYOMSUQw2cGU8TRB1FfdXeqAtaPEi+FIYdRaiO7I1gvv
zXT9DjnTJ1Ow8A67MDSnbc3KCuII/LJMGiSJgDCiPybBgKaEboVM7exql54HrIa3e7q7pZVT8IgA
7MVMigy3/j3AYOkA8zbB+JmWpbpNoUHr1WdhTVvljxhkxVAC5lZwDVJyfYNedLaIXl0QNx5dVQyi
PTYL/K+7p/4iDtC5rOSc89fP+564nJMePVweEEY4D+76FZa1xhk1n1foXU6tfoAIzUIwl2AkQiCJ
vYltrGu1TB9g3C7yIghOSXWj3Ct9xKGTPFoCQiKVbdaNHZr0kzicc4I7FObD1jQrrOh3lbRk+lFw
GMogYyhSRaAA9HUoZPsZX2cT1Ra3K6YZ+bFrnagUGKjFjhHder/IEJMPojpfogclaZJ7VFvV1k/y
Miq6q4JXJH7Y4CbfagqZcVm32NhNHsZDvIp6wHkmtGGLkqKXWB99x20fwYm9aU2YPS/e3mIxigMW
CoR7Szx7hJ5Il8nrZttr6B1apbyud6LgZO3FT7hDV8PAT7EyjAQcKCW9zS5n31VTHF9wBAxJdhfK
Nn8RKcfdOA5QyaTztFoQ/4p2QtMIdGfXREniPXWWFVVh5Zw4LucYqDAVW4jg/M2e+ZGNHiSA3Pdj
DkcyXaZgiu7Vek4825vfqMlYGI4o6pU0HBouo5E3bZa2JIadUPYGUcMaWf304Q7lpg7efIvxynhl
FPg27DlOyKArTWvDdf+bx2TJfNWbx0f3WuN+CrQwKv/KPBFHlylG5mxPM5lbljFNXZrRE9CWllzw
npk8vGqSHUrKzNRq1K3kXKU+1+nc9Vl1coxIJ9LEuAk5RCUbLyDeszcPEzPiRFx0Rh38Y2g5FOa6
Czp0AbP6ksmH1VOrRRUavDYj+w4LPz1fh/nSUFblc8KSXQH0jcXvIAltVyctQX1Qf7FXNpr7NoIE
8FhUILpu80UeeRFDqD6Qp2aTQRsld3Aze9eiyOhn+skqukkovgI4K/NYG+4Wp4ZRyNfWHw4lgnwt
xBl3DCECMHg2Sfq7mhoWUcrd+qODCOnEeissUbSqMSrTmkBNMHES+25NcC+4Yp/TIwQ4LwLoh6T5
cj6GIO5gYtbv0gnZGUU2SeMh6TmopZMyI95a9uut8IX/5ggNbKiRKgbtmNpwMv7EZWh9ZmVEBWld
iyZ8Rv3Fi/oCPREHYMMPgeBeWwRta2A/0BfKvpknNxAbcLUGzb+CH75Y8uJhoBZPC8eEkRj5IxwI
SvZw0gunnaStsGvbkxlQPauF86utVI29EGEF97GZY52eQ9wIzjZ94TMAb8ZQVgUHjdRJrwcNxqQm
80XBzwB/ioalVUqtrzoRSWz6fNnfETWP3+yGl7N1xFsTrGXrnE3i+boYOMOqfM9HH/He7cV2O/Kq
w2BLdI89V7m7Fiage74Pby+XywhOsq9CNIAg9qtyEC3W56rKzwqaf1vlfuzvidlLbUNLm6vwQycv
1ugxUK+XjHAWrsOnpUbhKMwjW6PbmUU+9CGXaGoqPKbsdXb/EyagTRfqEmHsFXjxMuNpUSyt+KsJ
0EduBL2wTYmicQGtwlzQsK0sDLqtk6ryzBc1kEY6pWO7wabpJonAVIEMKugQGNRfhpPxnRIFDOWr
ftAFzXmsRqhN3F2+NK/VYMEduuRCikvmHUbBODqmI6gMIDAhuamWySovUdks1TsCxXB6hKtG1NSM
FgagmYTXsi7Sz/OxnEKW1YWi0xZq2xJjyPBTna1MD2AF70yUrPxdBZMLMxils2Ce+ODNhAvUKFSc
G7YUWi0OIePlIjGYNqB8Y4dCUyXzfs9n7oG1Njn3CVPPYAXF7xqlXpkdQ/SgNAGkldXYELQMXIJe
swj8mwSw8xhJXSEiAaQmGFRVkL8SDudxCTc2A20KZLSSfITzZKXERj9weSQqZ4cHRdTDeO5BBuaN
frN1z4JW50gHqtzNvFZtnIthW8npwQsZvh86iY9325UMzo7AoQx4wsFF5ooN5JwAuhapiGnai++c
OUV/AuiuSU/y2kYZh5mHoHs0lrP4yegoJwqrUReqUjKarfd0+IKEEAPGA6S1Kr1auG1kqI8ifIbi
tN/YXKifiDAjNrk8kUeRAlVxFoELf9T5U36OlVzJSwgGL9+Be2LxblzmqoZz5KYlc12g2isK4mJI
biq1/2la4Vjx9mALT9IsvusOOnAHOIe7duC5xBehHYs/086ZCkMG+4wZ/ffXIo3rEkzx7mahHLMH
m8InfJTcvDftp4gXuMnJkSwAqvrbHCOvC8XeDx4z+v3FtkX3eNAj4QB1OyXFvtL0Q/dywGlXLwYQ
QhYvbPSiB1xERapmEFK2XmoGSlDF0ZzOoAnLA+aYEMYgDPz+oCxSycIoo3uVCrIN9cC+2tlWc3KM
9AfQe8pldAGUtpIR8qNZjbxAnUSVTvQ8BsSCfjqAFfP4MW7djdeK4wZAMNdCcoRg5IPxp6T5hrox
b9U9o8Bwrhvb1XRHJKkj697h6aWDIU+jKg+BXqX81BQUqmuV/WKLTpwPCgmVhX618yf05R5h3v0j
mroDJ67d+HruvdVpu81F/1K0Ax0ttAkviYuCcp8meiUoMaD0IKjuVIuh6RUYb1zIg3oLRwgZfwTW
yLdzBGBPeQv0KyS+ZxvkCoh9l0fTzgXhRl2ZhMabJmyaIZwvdBFAwoZwuCMZG7VxiSV8JCpSz9T0
B8gp3EQARA3wAn9LEkbRBr/o+Erfk6Lm/nFURBHmoryNxhlixzFM5hp+Y9KIUPiEHAs3P2kpagad
y3zWjacjJK2p6S/cYeCPms4P6AATyvyrwP+N+zS6EjWC+cnA19g8UiwBcjVbd78OpPuaa1YqU8qV
BP3Db+ZWPcSzxBdsGX7kh3Ai9mG9mzd7ido450la5slSaL93lQUEsTwPy+jrjUUNh/bpVEwJQLQP
S5atlPff1PbgGHJRxGslkhefYJshSrUIwsuOXNGAbKlsnHwZflfDis9x5csyQmsMgE+julZ8CTFj
xNbUEVQZXdS6MEUZjvQPBiIFfYhakmZGoNzods+YGYx/h0bMvqr7NsgDXFF4+d06TnlYpVMEG/fH
yf/hM8L2M4aKmIsoEPjy5xVEiq9cZuiZKJ4SG/PZTVurCbkcdxSjJ0rcA7Zn+zrzXL/OA7FPpiRL
icNRPh7qJKz5/7dwsfD3pHB49kgl9fLEBkrSgW1H71Q9Qa99NmHt/nk61PoH7Y+0kpL/D1KgcmUW
SgIbz8VY3JmJbKBpkO7wh2kKj8E9LKeY0FGjHrtyBgU0fpxmsiOcYbsWT8197Mdwrg8tQAL2pqt7
RiFrCiIdFDD7igBW//XxcDZXvggUyZYk1lEqIkB/fJbsVA5Opcgz00vtp/RvhX8REmGhctSnItCX
Q3rh+XRj9B7yw30lepfHECF/Q+uvsoXecHsC3kb7F3LgJoD8/CVD0NMb2wtSHqJWO6TZGl/1U0cF
hGtlTC3tEgnGMC9FJP+EmYLdpSRaroj2eoUIQexYVQonwKHKYpfZnQQ+H0geq6KQ5a2pC8WtwK+5
GA8g9gGEr+hOhs1UI3AK3jXox46YQEP7SaANAenfs1qiplilLsaKGxRrLcegKX+qXIHwJ1yJWe0X
kWdItR4R4BNs19nPEMf7wo+Hz6aPJvp8luitwYLz/SpUoMkEp0YArLtGsoHGUkFWC7MgN9S3HxK/
WeLs8/vOT3HTxA7BrK6uHdQPQrEGSqpv0pnRNxMLsLQrCBtg3xpaxs+UEr3NjSA7Y3mzhQDnD7l1
go7WtCg6qnbvE/vZtCnn3y9ruOZP0WMdn3G5uFMF9CMLep0Vvx/el3WRCteGUGS0xlZN7D8BxorK
fB6bT3clEgP1p3IwMdp8yiuxKf6rsSDj/UQZlYN0GI6ps9RO0d91271qWjZmxHcqrDcfKT3F4Kas
Cw1tFUkDpfc99gWudbS5bnI64sN+BVWEawwy7pz4nWjal3tC9+PyfAKXlJoUOMGk3uMqgdZCXPNN
G8C37twi/DFoB4mJ4t56gqdm2fbLhntCobWevFtir8PrwG2iVHuBx/uE8YJLv3LzI3l5nQZlD6dv
UQ1rwGMoEnyfYeahOAVXRjyuyoS+3KQ8hAr4JmPZHnHGFmc2vitP9HSsw/x8JGpDuAWxNkgIsBJF
fdqUHyin263M18Kuv5WM0Fn74F0e7MfbY1yXIyzi2mQFYoRJVNcnPo1DOlYJijB0Vr3YY5ft8fD0
+ak7GR1SCZ8CQ4EJey+kZOukCEQ/oWjOXY2kancnxK039aa/sTVf+b4YH22uJdlYGtVLQIVKW3lP
IToix5i/ka1BxyWv+BWqft/tjQROtkSAv/+EjnrIg0EfCDL6GVnbvJQpUlH+JXLL8mFSFbTjiYJZ
OIbiXfHnciylLTT8p3UGHRT/ur0B4OXCssAWZymYk6Ausi3JadWp60cbVDujCcinJ1xmUHRRiBAq
txFqR/S+Cf7Pn/KXq5hwW8z+t8FFVLwxP0R8H0fPwARjP2hO8cX2YkTmy6pbUDxz5tCk1UvIp/cV
H5BGKeDspgI60rMpasHgUEYamQAQAmRwh2betLwRlmedVy0gbhRrxkozOeMadZxtX0jMPFAt/2Mg
vKusr4W6NU+/ZXseU1aSh4AwrNU8+Y+jRLLLLTDYgJsDpEn9SNqVcA+YPXB5gXKO/A7ESgsEx6iu
kSJEdEXjF4xCX1irXI5yXLnF/h5XDWujYQjLpyIXhu8gUJpaJMZyGu00Gr6Kv5B2kvnRJBShfTfa
P3kqklwJ2r2xxmzl29/DuskjkazuWwSBQ2Yg5O9T5/6KQXv6xqDaYJgUr2p5qjptThBEPxICgfwL
c52rZl43j+S2EHi7wEJUgYxZGY1DSf6m0S8q1Lr1Y1yBe5531VvzEmGnrPRZzhyF6UhIvACELe8d
aSdxDP1WANqtL/L7d/MtUsFaf5EYrDsHPlTnJaHfRl5rcqdIoLw0rg9W/FaePAcjhg5V10dZdHBr
WjjKa8zYMIdsCgPptRnWNBin0own2V+pk5iddeXsgMPTXmvTT0xCGZpudJMpVzCLwTAteLaGyONl
n2X808IkXDjzz4y2U510tm8FWz/DsgLdTpRvj8TY01iWlSDLbzlK+/j3fWzxlOwO7EymVe3YB/oQ
l+KqRrMF2X9f2MWfEUdDQOCcmVMrTo/btBWCppO9aYcwM7FkXWuwjVT0fbUTCUV71i2poAyeApNS
hZ5us+BHx8efjf1LQkRjCNLthqg3NCfDo2jCJGqrUEp25mY1eQclFKHDG1Wrh8MxcItV8eU6KM9w
9EJVRaPh634UWt6T8dt1LJ5xEHDomTxeelfUix9Db4SmWjJvubi91xZdSx3zq3oHy3vQJchQNXVh
q2b5zb1ZBSr0QDO7PjmK0goVFwIBkAQuNAnzHsz3YSjwWibb1P23Irj6NCVPVpEt1W45Q10dm0lh
VkRRjzXEJE1gHcSDrmwh6khJqPVjW4a2Y8tA0Jia9X3aTy0VHIDeakHP2PDms2/82M5YZVgVIhEx
qGJqksU99IONYmjppgOMIemQrt5y24YzDWjAbfU1cLrTXYW8+0kYAUdaoL/R4/VXDrp1hYF1XuxV
KJiS2yVTuYC6BnTVjEN13KLnWRRuC6uKnf5h8KBQv+HTYMmFNyDwNi/zC7AIqqsAmGx+iGVTLHVF
wWmjtBTPR8G+jMRoHVmX0AD28djY5r10feT/mlGj8myc7zs8P5+P7Ls37Ei5s3H35zrfIvQzvmMu
Z3maNZzDSk3hyeFsMCup6DR6ZsysK0eKWH4fVD+qJc0/csOX+xt7crW1rkr0IDd9Sb/Qqs89QSfb
bH0aJjErkt+fEJEFeH0VyD9vXfNG4L8LIqH/fCtZyDmdksFD40LJO32zpwZDxTHzEFi27g1vPwPx
oynS0MprbaKDk/yTEfUneUPKyjIc5hG0pxqs71to3RIo72fl58YmZVY9/XtAtrNo7x3rbkOkvV1C
XpAb8YwRQkQbJTpeNDDhuxj2qZZkRzYB88LsOVK+lT0pYEbTalTQfoUshNn8zWkMnERTFOjs4sHH
2fh+R2Q0XsxJW3TBRcJE40gxrf7iDVWukOJNrW7cfdxHDPBuydfvF5W1dqSlHQQ1y5WvGmwGfvxW
iiraEvJFuXyd8zcORKeE0V4U9T/jLnmpQ66t9yEBFFJ4JblSyu2ytQDHZ5tv5BrW8OMbdOJ3rHuE
XTVws4c4QpaiLpIlCgsG2X6rY/Z3I8T3cWXWtVk/j0TgBsWrB/CwTM/FfXuouxdhsJ3PKNUIvY3w
h45bBoq0PtbUctX2XWRim+mrWk2ji15xedVC9u+th5I6HnVoGi7/e/Am+7+2SuMVYf9GkglcU+Wo
pOW4xSnCwSwuFayPVyuISF/uS//0jeoZR27AQi83o2D7awCd8W9qHjGWZeIlFyyriJaxDFksRDq8
gGvMySbclz6P/g1sYUrjYg0vvwqUQ27XYjY7s0jn4gJUToyyOaSyDyHpH8y1WHeX91IjUrFDDl4Q
JCt4QsxFw08Y1Lb0g7Wld6V9gX6RPifya8B7gALTfEVN71EoPlo1gybpGofKK9cCRikNK2RP6F6z
xMf+CMQkFAt5UQgR3g1ju2fQBzCa+VS7p+GqGItMPupkW17BDOcyknB7OrbCUH5Br+uGVHRiNR+U
100o3Bo2MCrt3Oybx5Uywl6m6eGkNvkqJRIKvvyNFJKz2VfaHoOPbTLvgNujjMljK5WbAWju8ysH
SXIk/XWIM4ht5xpqUnVvempvP92b/42zuqWnIpNEQqf/vmWkMC/Zcbz5IPSVRLm6QHzCg6T/zQG4
AyUeXAOsvNgJvwFYHQfdiSuA3wehTZH/H/k2Xi4Bv78L4SKF0MoO4pF76I/lLjcywXusnNgt+OdL
7M2H6mzQfVzk6rG6qG48mSUylHHV5/U4nghTr5Gt1Z/q/Szc8HonOErBZhjswVPmX5xJwwhKRZ8z
tMoya9RmOEmgX52FUQe7iG5xy+HP2QqnT7/0RwYee/BO3O4MMMe3/CwD9WLLaEIJeKZbXbdmBnuM
vedaXmzZsta5skMQNj/evTxzkkDJ+rMN6kT3gwIUEcV1keFhz9+zfA/M1RLklr+sA4UA9ckHK7vU
l0zqdzsOu3FhCtZUjoUu6PQ8t8UYkcAiOuU7bYMqjAJJKQReeV+WFD4mREip+neOdE6GlxtiSGPs
vbyQhuE21T5yXUMmrcgXHzN2+36zC3eMeDw/1nNOnp6OiflTHAH2hVlmMX2N8gLOTpkRrhB+eP4G
rwkwS/5/hjwrJEDBsI0ZAfIhyep/2oyx+b9NiCLW592ctiLPeaEIKEP4dN2ObRfLSBGqHlnIBT7M
QkBDfhqgQ0eFkuUwOB4nTN3/0l9FNcA/aZpvfUh3ms+COLjUM+kerd1Dya4PXebYMRDCsFREmBmu
WKZIVFF3qZ0jbgTNJ+sUpMG4RMeVsZ1vRBwymzDtlaE46XpdHnqlVISqxuCbyuGxR2C5znQtsHel
oU12sPfJh3Jf6vlywdGrGVm2/D7z7QNrvRy9pVEhgA6VH4f7a6fRF81R1U8EZu/2YiBbyjTPEjhy
86yIiPahzoHP6sLDonNE0XUUbJSkOxWLM0MziQ8swChdE+6tRBKimVGD9Kk3oIv/e0k1JkiFv52X
kplmRNtWVa1Hh1Zsi9a5NXeDsBsOwlNXdlq/4zNUKiGef/xnrFAaK7RReLqmGkIMYXOhLlVTwftd
6i/fQHXipoHqaR3Utpk5vgmQxBPFEkt5uMtHeBbVeXgCLajt4He7qlofUuisFBIPKwbMoOzkhjtb
zQrho51yb9lLPfreJEViJ5tS9/fwCUAPai5v+23S2LQeUf21+H7lNuQWr4vbefmrEbPWsr6YBCHh
hDFQso7AbdAwe2/mGn855UDuDcuLlFm0o2alygtvAoT17PUW4OvE30SOBYTjslJ2sBOC5FiX1X3Q
ywGb5PC1grKoUo2gE++Yu2KdPhc9BK7yocI+AWisXSOMOm7Q7mnDXR+b4ygYnzuv8NeXmHvI22R7
4taxS0r34G3rbZtCKFwJvvDGjBDPY7JxMKPYeZ/ZTH9ptKqaDHdw83AxCzyI1roehEFvjBzJuszu
BkjHM63GJsW+qv2JESXnWGzJJUGBLNjUw77OlbBhkvd1kBxcHXI05WnpEItzeUa184vb0O+FPi7K
L8heqa3k12X7gnsBgqu/dj9iGsSoFO7UwzVj0qgPviJTr1QpygdWgumhB5AYLqjB+B2ukXDa0A8Y
kyjF1OD2qV0I2Yd7T6IeIDEaP1lfpEcYsAV97Oq+uO3xldgJdrojyMTY3V5r+fuMhwQ3jYsdSB/m
2aPLz9RshZmCNsqD9wmEMU8YVf5N6FPBeNUM1EYyVn2UCwUelLAa4FH6bvqxrfYPKbwm41JQMEUB
jde592qX4ti+cw7F28xnLJBOtrXCB/uqHxP8xhWkKFktis+ANiNon+rXhViVPLFsBiP2S/XqKCvZ
EpMOkKv5xt+LPGbcNrT7b96qxehuXBjpev3L+6HqM6ly8O4GyLRQopeS8w7ElPv9lc339n88rX4A
ONEoVceqM+hvZeaicQEPU9ecK0GoXdgu7ioxTYJ13cosRH/urWxdfQaoUDdcDTKuvI46t2Jmg5M5
QD1bqLFaLleCGvDIJ9XRavXmtjk+LAeirpyyZJqugCzvytp0Zkt6R6WTUM+PQ3oK/mi9QcwHgNKx
MIZcZ5ZztemO3UgyYPHylY/nGIgIVVwtX4bd+eO+LmMJj+p92pDP8fziAszvAhsmRAYeo+A4n1/n
mqCKFf97RQ1v9460WXvuZEg1G3Mx70P5Rfxau2Y5+X0rZX2JlT865EHvMt0To5EQLkM9wg4yenXZ
kYKtUpl3ERAREcdCaBE9O8XAviwA1L2gPIMkOtGRAuVmjEYD3UjHhtyu8iC6dNqYQ+nsWPr6CavQ
6kNJ8xEUkYPB+U8Nq4vhdSo2r7qZYAh6dAdY4ciGJdkg2CmjtrfUfZ09iFi6/YtlYVpyP5oByFoK
a1N+6b6xfkz2RpaS+j9HLnV2xYMB0ckT7RIW45e/c9mB+1lAIKDU1x9fERG57HPWsS20MMqcA6Qd
4JL+6z0M7IN+eMfKZMsMrtl+v32Sv00WXK1B76stM76rk7YYDpyrhmME7K3Esa8MIU0QjFRs6QGC
H8XaIK5GlQrPsh7QB2LL4P5n//5dBLsSASu+dPugv/kcGVF1vCjCmbirtcwf/j0IqXHbOUfTgs2j
ZVPJFK3hP4wjkung1KXZzUiSIBsgwGHPHaC2/89wkvWhkaKohq6pt452xg8u9kjKet+c9tATxs/k
tvXx/igSCVTyhxLogawj4iMI/Vv43RpUReJyZ61Fw6Img6+ksDeA8SjAE5wHlPm3UjvZa+YA66dD
TiZEr70SDRGodqI6OAWmrZHil9MxmF8NpvZj4zvFbuvgQNxb6qHWmRRYkb8ultQsjL2bN8z2Z08u
xLWnVpxMLzOiUjc4f+Z1EbblQZAo8kH61MYw9SjdS2YdVsv2r4Lc4Xv/u3hjsB/cWCMF4XNsrgI+
0SJYM3QTtGNKxUi5PdVbez+CoVpakjlsG9XhnCm+vURcYlUaK4t9hIGJhe/ZQ+Ns94cBqD0mbgzF
3K/36bScAvbStc10d4Y39SxVWRvFGWamuQUsxszSMSMFfYBdMV7+q00nvRJhg3Ootpq3rOuEMeAh
QVXXpqQ2sVz/Cg5Z3mU7XMT2fW0sY7PizDp2wfZkxi26TMrDjhICxLG/5SRwcY4WHMLg8UQNtThj
bXVl2cN4282XMPzALoJu3RnjnMb7kQpsj/nVgVyaSxspJJseDNG9QMgpxfOosdm5uhEZH9kcu+Pd
j7xHsza9z4EyzGZHL+0eFi+Hsc5qu1u6v1HQKmXGJNKlSjvN0aV7dGKOLFXrHhf0B0GWB1srqwvX
j9oY0RBTnPuzcyvg0+AfXh2dHiHD5EFZPV00cKKKcinRd4NOoPXEJbJXbPbn9p7rBPTZ1Al1W9d+
qAEgKcS4chrMgjYQHzXHF/JIxR/hENqj7yq2x8csr74ZHqTo1Y2xjlaZ+WlS6f0DTNQlYBeRCWb+
K+nWRKRGOL4UP8IVzoIQ/ui+yYg4ZP8+U1fToUYYuvI+MwkJVF8SdB472g6CwQJLYMBMpka97QE4
u3mDnz7OlQ6xD5BxlpxaKK73Zl3mhs6Am/aCPycsDAI8dRbCUCZ7awld3e86Elx/4vvDqYoFgtIi
utyj3jOUUnUwPRLbax5PVt2Fy6z6YpENuHWUxOQUVG60foBvkD0g1c+yXavk/n2YdKtngFVqdM6t
lNp9kakjsCO/cPjEEiOXIHI0nuLnpPDqbEaPqyusL4sNxu+P2kyl3RZXbKFG7gLrJt+UAuq21iC3
WcpMTFjWqctJB3mKQTsivuPiRKq6XPSfAA7pDxcosNO7ld2bFceTwypObcu9zgZmdqTO3NyMZl7K
s7txjWWK0k8FvYx6gKsF01D7DnlPwv2cjofU05xAqzrhzPRHdxLuVCxK49a0mKZq2N4P6QOtw8Ec
ZEyAFgIrIbBG5GA9EvdE04+quRgm9QR2F7nc3QNadcNHGNxRKZQONowfq+f00j+3OtsRu4DmOusi
PL9ZZk1ytYQdeBswJ7b7GyxlA+6zvM9+1D88c9IG/pY1+B5Sx5iiRrN8fdPshLSE/5+FMW7hZsFz
J+Ye3Swaxe1qbcH8UaGaaBD0IgADPobD5iDA2HUqjbT8Wck3dvjUw8TCgBVZROq7EVu2D4FOMlEs
IZAQPkRAMuWlaPYXMoLTdgzEL74kuv0ylM3F3N/Tq91LqGnGMe3ToO6OnoKPgrtfzMz2NeKKpvG+
G5O5DTUT9akReLpWnshJoDC4+J/e4wwbV4wIK6AP9YNSkXvmnAteWEvgI5xZTGJXTStldVNzBUl/
XlTwTCi4PZbSIaK6vylXIJXJUI6akU5fSQwFbRcswpmpAYoTRyO1tVUGmmQchFWYw8hTlLNCL8F4
PrU9YAm4P/lB+ySnWUlpo5JP/3EQGQtwokBgTHve1CEGySyf3z+mdeNOG6OaoDDpqNnynukecqKR
JI5L+3JgHWmxz53wSpciLJQQsnxD00C02F+ZOpRNOU/Bb1VoEpOKyna4B2Ux21cXuZ11HvlFZr2O
lzLIitLgN027eU2N/EYlva1gxL2jsAZUEmi7RxHZd42iA5e1l1MuYw+oTa9cyjvRrPXhZYMRYCDF
aVs0rObmu7dhC+78f8F5LkHHqkS/HROYZiN5RaAsQgHmFJHLEIZYrPbWCpmoviPCDn++g46OBpQ4
j20saoSovXqhiq8EpPaaGd5ru9bvJN3qP9Hk+CG95WTiAc6lWw7aHb4C3NOzLOQboFRz66XtR302
OkP4tv3sFv5pgVFgJ4i/2Jl/6bF1dJP7m5ggveHb/FD5COc7IoVM6sHsOfDyw6zqr7i8SswN1mIW
jNC9Y2EUPhJdlwiKf3AnbvFPvNFA3FzAJXvM2B/G12UhGehx4D+brCG8S+/4SdZcjGXXq/3z5lvr
/9dj7gmxOz9sAc8qULQzaKbc5PIGCfIBYrLeruTMTa2TDIHx2GSPD3NUn2l5kYD812RzRe3Micv5
LXr1Ppj26DS+JLd6v85y7FwqMiIFpNzJmFvJwy8GrR/b1poanVdQkL5PnH3D8NDT/IKS1Kkh8lVA
XxQmkv+aRW9ssfghYY6yiHcJ4lAoQVGsWkZqdeRzE7cWNlcaJIAick0f5ssJWtxeI6m+mX71fIJz
ASB94DUsXeQiUCi/aOcjx7TN/6ieDvs2O+X9pjIJs+6URHk4r4ygkvpJulvI5x9SnQz0okS6bl6p
znDsiWwUeWPb34AQe1y0zV8Xg8NI7hlNTqhmGqbBcQmIEwhHh9pEP7Y98QLH1r9JBlsIxNpPcIzh
NUUT0Te4pn4Js3h1T7QUWBWHn44jzBjm4MKL9hNZs58FXSSogy4G75SZelR0Lc0tLch+9VH4psK/
c25mUn14mEZtgUaClhhts4LnJjUgHAV4ahnUZQ3P5Q8eOEpHFqL2S+RDs6fAdpk9F+m/6KJs6bqp
+nXeTSIVqeMbcqk3C5eXg21OQ+rDPyc1eU/c72crTnR0HBQCERchYxhOVhaCAMKwcWcJXMMNiAzq
hj7wln83qMbIE8H9f+Ld61Oo4EMBOkYV+mU2w6M0gLzHA0VDVu0/Wk5w+xyOKm31Zkrj+cNev6Kw
mQ1gtg3nrgZlaWC4UdG8brfUXnPRc9SIBB/QWTEJMiC6JZ4gOpub+fkaIoiPEPhp5+CoaqBCORLL
ERyLg5maIfEKEEeFtQ4Rs1sdgt4i5md+DS/tGFfMQ5lyjJkKO0miipxDlm/BqJyli4DT8QCy0AtA
G4AvW8Acx+BNF/EqJtUbJd7u+yug/yMleeGN3AGs3jmvpe+LXgDbdMDDf62Jsm8alYfqQpFxxtMR
5Uo3EqwurMe54oNe0Yol9eTRdLptTdH6aUh7GgUUHvpNYD/6EU9AzU7XfqbsYRjWp0JXlWfbHRQa
9I9GmZWpgpIFdTmE2TP5wgmQ/jytoG6I3j4/OmeU3rKxInkhvas6hbC8QtZEnmqIgD13d/p8RQLI
kls2mb0VCAqgb5IyggheH60vS2peEMbZEzNHjW/In9LKhMeC1uLtNcGsYrBjjXjV7xJ0gjdDzD0R
TlOA1SPBQQHbbTCG2O4oi+oS7+436YgOXjPLPd4ZJWH1gkfx822YlPUKsZ0axeokrFCtZQDBRVfQ
wi+tlCSYNyk/xY+OVvkVXg0AKdcKkngf2gLrNGDBAFAwUOpaqS9w1225RnDqU91/Ovx8A23Cs+LH
WTcKDTVGowDlTlJiq2yDlnIAzoyAa64fvcdKVoMZ3cqvNq/3US0DWbJNo5wkQgMf1SWzum1trzQl
iQ9YvHFTGITwZknrv7grdn8Co+UQBeYblsInvF2Mew5Mv+bUaWME7xW2/wgTqR/MWo+0c1W4Fpme
Ly0NlcplfvypUetMsRglDmvkkLt4hbqegRxS0DDzMyvsR9Zdfv6ng+9cyexAgnA/uPWc6V5wKX1Y
NmCv9nqiO/Z1ZTmeFs/2uAnziBXiUHSEL/WCFQL0L85XzWQE1d2zgoc3Szcdlm2UP2r7ASV/Y5N0
/0UZnGvyZuqKKrF3dY+TNrBe55eRq9teyO1Lzp9TRH4Wb0pqGKp2A2XMPL906JSa8jcOuKAS8+0A
SUSugqXEeFSUwaRMaLHC86Q5p7r6ei/1nw6Dko5tSboj06M6U13W0bT678iyajWotUanLbQ6fnm+
V4H6zRp6IB6l3n/BJdJXW0wCvBwrmwGGpvNXHG7Kw6H19ArR3AgAb+NeKSS+tkOiD2qC1lnXl7Yz
+6ABuxvkdKi4JOMn7/kT9I6RVfV2Zp8Zu2MO+HXdPpvQ7Y89TQY03o6ESP/8VYOkzj9Zz8RODytu
FKDrjZEnCBVlziXR/0DtIFVlHr8nlSDlBQ5hFr2L8DAjiHVnoH7d5aFr8MOFx5nuzTMDGNam6N6D
C4wYwxE5rNEU3RHOan9WjxZtSe6KrDyD5zpO/ZFsAOvUnOrzQ4n4zVEk3cDiUavm7ET9x/v1rS4+
TjpkYW9wFz383UCvvns9vi9ePnNEv+E4QWBBqDVg7WahfPtWrZ1JS4iKghDPq2YGsz1umUHFv21w
ZyNQi1Stc1lb2ga3LwV76qdvgtahgIaI9kXZTAdlpP49YKkbSq7jsf6Bx4qVQrqRH+NM3NBf2hlo
NXkXH/QUVpviMLwEbtthnKVGrHf4xM27tcYsWa4NTVB6SDH80gG63uoBwTonSR4W23wAP3PkwjnQ
rvdlMYcqRKWAgqdR8EmWwqyauNNk4P/JO4p7D2ab5B8zlrAKcXdWDlYReN/gv1Q47tWRfMkntSVP
5RDgMbQFAc0vYUA56pA2EVCF+PEb8KCG9tx217qT9koYzJG5UT710TexgtF5WZIb60gglSVJGsSR
jvloTCz9RXBCZN+1M/a4P0fNWZQlB4aqJ8iqM2hbsPCXkFoiLq8JwtFlxQwRV2VhuU6odTAaY5X3
b90sMF+Y1JHFmKhyl9JeOVFsSZBHcAT9UJAWhpEma9rn3J+AqEDxJeHhNBdXN7hHmLIpltD44QLM
vSh6xmmkXfuTsWBp2vUeR7ezJz5CZPdAl58S96X37WnaUk0pgP8f4PQvoYuQW/1o6xqGPYRgxZdZ
Ip0bcr9jAJPMxAZNk7J1VH86mkH6GRQ/JsMh18PDcB0UE689MqFgZK8dMik06Lz4iUp1vCEdowrX
vhj4Y2oSDLvPl6xvmT5uo9UytxvAQX3kmBFUYn3AM+M1z+oJccoPFiY1+tQj9VNqMjnP72aJy7A9
oybNC9OFW+UdJcBTh0fZEK1ySKZ9hDM6gaXa0Uy+Bgg3TFUO5XyTluvT+9NY+iR+FLJfWyp4Trau
5dvcL6TBzliTNNVlkgMlJZvqB7eDWlmeNoqDELfUjN2cPaJ8pe7DOkmFKzqyBjUMdmqERSfbPdbt
JcddbJdx9lZkb6MHwPJnvyX8JiuK0Jv4n07n5AyjupfSwow7VPBSk+GbBGM7Kosq+MLsf7FsfZJU
ldobTxFJk0NsbEiV7k95G/d85Mhxqg4XDnfOVXyL129hsAcAuo9Wpy0U6c5U8iwtOP6ODzEepTY8
VeK1Qu8lEWlr00s2fPP3TD7i0pQhsKlt7UCgce4f/jghfCaXIM0OHNJqSesAwiUgmLYxckv72Bi0
BNXZ/GJ/rrZeJklwJih+uk/9PcItp1WUW5G+9kqNpz0Nj+Kz91ASkuTlhMPrvKoyyGvvzJMTUxhU
KtsNG37/kjaBCOIGlaMUUNeWPAJzOkpQNTX5bRNmt8RO94gKMJ16igwN2hDtXXSKXFQr5yMracHu
RD0KxJn0Ckj0Rdv3w/u0oZdmgSYwmkakk4pmSZRbyH/hGpHbd1wpTEyFsT4mqB5s063uBJgKnyOW
CnqHsMIbl9qyZ6HkKpHpK+Ex12p7eC+0o68Ttq1nry6N/8lI701CDYqBm6EyKLXvhzdY+qxFjuqL
cw8nF7jU3n6pJkJgJNMiJt7/q/DAj2n5BZ0Tkbr/IG7oP8U+E3qQJp+9ZaMZ5oVdOfejGfSRZjdi
X7qADpfAgZTn5230J2fzShItxMDjon7jsQdD8jH848LdqswwZqPMlA01Sr8OwaoOz8FO+h3WMke6
tM98e7pJ//FYLvdM/tHX+hYDlsWiQdsEb69HpEZ5zXJ1x55AVR4+s3dotcsRXnKEQwB/uEXTOAHY
Z7DwGqu8g9KuyxLN1gFYBYxPFlBPmMihciUruwfJFs/61OJCXcuDGepxaomQzZWo5zJtn5ZkR0Ri
YdJyLCxkb1BFS5PWz5o5mz17TTWAokTHKD3qHCtnEFE3YAKQbIIGUVwhftiamOkLUKBI1hg2/Alj
gVFnhzOoRy1LfVf932Ua0XF/imfNOqt0hPR1z8/vXcL5251/pzp3QiXIUwumFS/A8LW3e/vmb4CR
u/rY4goTrzMLjKEG6xlHBD457XfbtM2IGKHuQA4Lt8nwIfMkEX/QEg57YZr1z+0CRo0HPr6b+T43
sc1aYudeI9zHXQf71bX4gZ5j09oZ9yLbq6ZKxDdvKGU+OejTL1ZvctVL4leLNvdzgrGv+/FAeBmt
UM8Jv1KxumXc7X6+iejbuxJbgxQvfgrJHH/73K9SsF8hLpuLF+2rLMscJaOtZrMirLheNSlMc3c0
yHatFE0C1BM07W7qVLffhqpfOGDBKeFirRlH8a0f2cZmY4FNv0JIwUJ7+xqLkn74vaE+CPMWdi1b
HSg9jZGJ0TYIoP9PkPjx/3hZx5ISLLU3aW6/EnhkRKb4VQynXKzBRBUAjKzua5WurgZFljOS8JQ9
/FyzG+OjX907TG/T5a8UW3BJ1Qr9HiNNZiENjBjuB9cM92Bgjvdw4WXXILa2i0LkWp8Ho4J8/Y6L
LTmOTByeeYFPxrbDpBGuKkr0Di1VyMtnHDZJaU97ZMMIhZJ4aymX8bgrt77dBZgOU1MpfM9ri1vi
Qy0nTC7Tcd6EVA7pr6RtkeStvUs0T5SCh4xLVaSJVXarUN+TIN7TAIfG2b/xct13VvpYq0xiENXm
xjt6T67XUY0Ovpkmhj4Sv3MdfoCi/thQxq9xhYhEP1kYJCWz3rtZ8HCkAn76jt0JoTD+gcmzhSMG
KlJ1/FYXcx0+iS9OBIaqLCGuMGxraadwo0tlik9PNVOOHpPp8C2JYS31kg/tz+k9qyuw1Iyl+L/2
v6eufKTu/N5LCwLRR/C5Ck4Wz51Vp6vpZiZOdMEQciF6MjN/UO7/w4/UK83fPkZSBdRsFizgCBW+
d+4NvBYKjh9GMOu0tts4sOzWiZa0Q+bsHkPt7gn0mkpbUVebcsc1PlEq/fmGhZS78odet8lQ+lmm
FuYMi7k2aTOaUP2QQuw1EFjIaT2XdnspecWpuA9eQyWjcqvH55Ubilk+pr70lQtsy+9YryhlQ049
S9HLgaiJliZwZiXtF4nYT6jSr2bcTUSe9Bc+BiXv0DuWArJoYYlO2SqQpXeIAUiVST5eUmpv56yZ
JnWK+BEFFr9s+XLFekbnRP08GcCWt/H8rsXHRfRCRJBJ2skfG1bGHuertEf/lgmWkp4cLNa/vS0S
HLWHspeRs89iVeNarWZg+aL7zfHXeyYAogU5+B0Ed+f3S4/dUN6NN52xPWMYGHJNWca1gF7j91BE
2QJdXrN5Py9e6yWMViYpeCezDQ/T2UGJsy1irLsI08/iN8Ld7ZkV7UDdoEqPPZ4iuSNHq8d3RwRj
5sUSrRwDEgm+Il3qWzFuEUVjWN7w6MdboSf8f71FqVE1yBaspcvqNMPJa7zHWRTCkKCsnlGg4j5X
nt5hih8RL6YLhom7hSnIj0oLc404oOuEk8IAinCjedD6Y9ZubEbHhzdkowsr6VWOKSQPgAiJiy2P
fcR62rJsAJXfz5BIpK5Wd2yyLvOeyttyZC9MwrfnfPjp+fjx05crM9wifoJwHgDwQ6ID955P6sgZ
tV8md4D3azwQa9JMY1mtiikpzOMS9RebSGWP/WzMxeqdiTE0hUNgOSTdBDHWHdyTDWpxuBv0einP
4LdtMO87iwDhzPSiNdlBj4eQt1BYq9Qk7FVtX9ibmftgkHfLcLejquTxUcBq1AbtepkyTjwq81et
97VDnXsOg9tdepOqWfax/HnjCPEmprqSpKtrN4IKdG4vfW6Pl8Xp4A55UncKuE4GuMh6FGYjkwWL
A2jfilG88dWPs65otGF7/fKoYeMdJJkQGRO+T5xaIRLpjy58fS8sRB569UQbkFVL29vOuYDfD9x9
4WFqV5nJSN/IM4fpaF7lcwayx/58Iu4BQmf9VvF3Vr4SdJoE+AZAmN8U15YqdS4SrGF9XdY12t+R
w7XGaRfz+648FnUq2TZdoVJLpJdXUPu6yKvF250et70Xm8fcfAVGUmERhWiS+GtV2swqpm9YJQDj
3jvlgtTmtSBsqGbxwzP9S+Zw8SIt97wV/R9xhNktNwotuqgJ0O6xkbZOnlZ1YNItyif3QUjrBDKu
k6/g74AOcXwhU6C5E46+RR4+bHWEkE8RUaDckMCepGrV/d1u/nTAdr5S5rvOg+V+1sXSqiBAHsxv
ldlugpZwH40A97VF3V6MCVLsQkZtjZ+AGECtbokPMNzHsrt3lwXXE39eBrCDKIA6xhbdhb1oFCkt
oiteTFF5UL3t6cmaFM/nMXHMrU8NiPXaK2cqo91IBb5XHtK1BEcTQDPhZwnTBdR/keTSAG4fh/J2
NI8Q/VEgWzIkBEz92R3gmWBNz2gqDv8onbG/rOf1b99/TNj6BqyGKCysAKUUN3vR+tsBL3FeyYe6
6BbpR/RoGNy447usYWw/13k1WU5Zw89etn+9gB8johxCTrGfzWsstoyqp9oqwGm7jALzM9ced9BQ
BRMj/rwT5pYw8UBbHRIW8BrKI5wpbK/RdNme79hNE1Fop9wI1jsJbkGNdcLyWbtP974Hft7aepSU
V7UCl2NVOoQEEcLbp2V79MR9vX52hJdDSu1cWoEzmHXU9xEG0uIJxtHjgoJI/LQVfVCBcYPNrMMf
s0bszKVyppTesluLXOoxU5LU1nO3nNg3OR64TjUm80bI9oGS+pOLxMxPKWRca/L5meF+1wgw44ey
WmVhhNGfZhkc6RL83Cdcf+r/WEThY5Zkd7SZlKQQFma5ozxf8f8zWbsq5Hr8VDlf1o2YjrggIKYm
B96ZXq4jVQdB86RLNfud/d5twTrJIHfWh8FSQrKXLgBMQyCjE++dfsH19IyGU7dALGDYhx0J7416
HBm1rlbRRfoYP0YiUTOskb9v5JR83H5jGMOX3t/UikntVZgXCTLabFEuQDzre6BD18hg5WNwyX9U
h2G5KBBW7uC0eclfgPuVVOtn911OFnIViBA5o+soKmzCA5BsSn3hPPlN7QPcpSWLCOmspxeJYzQ7
JtPbweQrofamMPxZX/heC5ukAXVBI8uZrGSdU/qridiJlbTaMPEpRZhNjrXt5pEh3y/TNiPEWcOC
mku8rKf9aI+B7fMqQ4WXb8KNPqZ/6cAVy+xH+IOR8iiWW8g9gguOvPz6q12IfpEYhACY2P2Zvidm
wIy+sBCJQqz2d7MXPjWRMZegNjCKY81Fbmc9++gMfiXbrgu3G8TYp/gfY6BxjvSdboj4YpiA1XbS
/yftMtQU+Kgzs/RHPyRfzDB/nWaWPhpoDyIXlRNaP80u0/Ua+GfFrGU1ZHSRa2tZjv+hoKXPE2z5
pcIGLAGILAjezqQApgqeN80uzKrGboRQEAKmuZcdN8uLl4lMq5xB2owwwWxc2zNzBgsjau5mAB5C
p27KSY9AN+7FG69EUJgpq0Dthn7jSME65TaSjT5OL72WhwHKE/h4+YZVWDcu/tR5q1sl7jcjetP8
p4Uo8WpqWT6Dc9weaHQ2uO+elUICzyQIU2lvGFUvANh0z4PwpSE6n6svSln+21cYoaHz25/psvuM
m1K3dTCKRKK/VWzDRu+3HmPX2els9sv13vD97KjV6o8v+6h3elKL2lCna3+duti9c85DEhYwejsl
xZaedAWiQ+qb+HqXcztXYT6vf8AgdTb1rGx/pTR9OAprH3j5ZjUgqInc/dB0mosvRPTX4CKyLgAB
1jJNLQjRT5/JoFY2xMJVV/N6OikYxJyn+d2pwgVdCLq+RyhsOo965ysoRhkCzpS5OFhiaYzBPN0G
7Xnr+wVVxPxlmaUMq1ffvbYwNuKSxqCG5KsdD/InSBHAPaDWo8RC0jBKpheQLiW/FLXpLkFfn7fc
VK2+aUPTNXE0eutwUxm279IrazjoTk58RaU5Ap5Z7bsLp+qYV4SUfVuQ8ZconYP60MVyDxHuSEK8
BR641ZXan7UShiUA7P2kcH+zbW/hztacjI7WI3zCtFbFuPZR6mnoM6CHaV5b2DS3azLb9jTUt1Es
xkRZmF05l7T2JFW1q8BSDszarxdKlccB+5i3VOwCCq9xV4OINDqP8SEFAM8wmUaYkQnp/6LoDMR8
VuJboDLkbuaVj4s0Y2HAdJMVZjfQS8QxMqpNXAcAkFAAcKZXx4VqRci/726gVzyLVq8oZmhpse6X
uT2CfikFZyfeL901QtYEEbM65SHHLytRUkxoUxcMwg2RV8f+yrp6aITvJ65SAQ8+VGjtlAdbuMKp
aLgvLoGIGN1XJuUAKqYwZREW25wrcgQllOy92JFi+aqh4BryfWFyZ5vF8lOxAjBmbwjKbWbqCETZ
Kx9vNFzPsR/9+QPrApuBuLZtTMZFX6hOdzD56Co80L7YWm8A1bjg/b9IgZC7idarunAkVgP8OO3B
1VybhCCPqn8/3IypOWo0Wv3dphJkspbGHzqxYFYy/SALYt7YfR8dTwj0q0oa0DmgJt1o4nAAP6Cb
ct6S2arZzdKofLP8z0kTqbq55oAoA4xGyer+KVB/XtXqF84x4Xv+/442m+clGaJyuNNew6zhG8NF
th7UVGAc2Oe7j0T0H3Q4BMJS6ZkNbEFso+J+Y9Qvn2Ar3q37cd3QXGi68Ml6/fFN3/kbZPgmACZ4
gK+BIZXKkFISpyHLfsMrhniFNnBvpi7QKvaxIhhPwaR7udj1ka8XIY8tq8D1AEmcTbx3SGxVrebb
NDMj1Dajv6OOa2N08anJN6Kencxi5ql1Yye2beVF26GnZMbXgC9deT2fYqjm1VmuaoWqYZv0zRuC
hvq+Roz2aweMV45lvUKJ/1vqA86NPAygeglzI3MHQvsi1n0oup1uaWoWj91q4dMOIOUD25ZaTRSN
6L2U8VyBMGvB94dMY52ZzmWXklnlq4OAPhRMl2pAzNxmF8sApbh4HO4TH0V1mXqq1jLO4bvb6jQb
2K0Mm2z30CdcISss1bsjMpp1NGcDOT7SVGl0vIUw2X9P7nQf1rM0CuWMzAV4qVq8kl62kxSCcumy
uPc+vvIamh7ddtlPrbgKedRWA2XAuldyVawX6qKPLalmWQ3qYKqN9BnqQVY3+RAwKjPl+1Jz3GZH
/ruJ6t1tpIDE/aFw2dVZslxKbCdSY1JokCgNsMJjlYnOLWd0qZEbs7AN/AOMMNisjibuLttM+rq4
wdZAr2PVLdIqNMDlotanXFbzHz1m69JC4e1BOl6n8bYfYpNHJcSLp0DQtvBlpXWYY3chvgDmzYFM
b6Wyrq7maSlF1V+0tJafbym9XZsAQYERBIYuWbCxdSUWAIq4JWptKWLhWQySvxYaTGlCUAmgr7MJ
ruXHVx3U6+MQixeP052u1HPsFDwC+mbAMxHPnL5sGmdITnbE50bD6QVs51EmLPrcon57GHocMXlH
sGm2DXp3b5EJgLnCfsgmhJ3EYP6wLbn89P51YHQMW/YbzN73sYb7uhZdFUEKemYh/G7slcio9zT1
WfKCNNS2sb+YeaWtS6F9/2HYSfVuCnNOSiJxdJ+viFeMWhwBoT9TFSsuLOKDbhRnC2zqnOcURW4A
VA6TVxbBF/cY9uzJc13jt1cVQVoFnjHJLgMuLK68l/XYqkKt3Dy/5yt7cukLZ/dkj7pVjXgDJSoy
5Jwxc16HPNYbqrQw1lMseBosLhHrfFQpgYO6gf5Kb4HlrFw7GIedm8Lo9jxF9+pcGKkYR+ueizQs
PDsMWlKnXk5s48kLfivRy8Nm+kGwiLlYRHFHy5pzoayWcwZpdku50kSWWCNVJMBwoxYeayt15/Pe
DmKhiQ0YbdGsIBCeWBIFvtdKsOgjALZ/0l0HgrTD6fC6mP8XA92PMJT9IT46B1YKxXDy4hFs4uJA
51/PDaz/k3YySp9w7bL+G7cMg5meQIq0CeOdIwVN1iHHlq3iepV/MOQ4dUhfpTN6N3dLT73tnMwK
Gq8DanEczkx8GffREjU/KxLwnMe3sorZ0JxPIGDxcLo9UevbxjQ0fPVKoAaETWdr/0Gk12L43+Ao
8sJJBkBqImqPKUfv+q6d4UxYdk7N4OR2B9+RNeSV34+R0o14Y0SdwiecuHNXwyDT4kgoqFf8kCS0
EpMSOR/7dbytld/21/egm4Ru8L2W6KSdzUvKG0DU52iKf+IJfzdvdxZr0j5yxtoZeI83uANWDwxX
DZpgndeT5hsDRM0a5hVsiuY1O/XZGCyPzUOQ6uXj0trNF32D60JtOeJeeQ6NkPwkSIY6jLLbIG6c
eAcCGlz1998YtFjvakUgnCy7jXS9gTE1vgBlN6nYCNp4toNJNY9Jp7V9hwtdkPjJeE39ngICk/Yh
h9zBMsISr0GHozjSXMt6l/NQNdbJC+PGMjjaTjgtfTBVmJ5ctBU63ayDJsoTSakRG1b08a3hbKDi
0PWG7yReQl/UJl69MBfPkPwHGmK8o1sANpd5efXynmSHBd5s+HVQcKPw0eA8nzvcDu30hYcG9nkQ
Nynoet9c3fEqwxlwpoTh5ycNqGXo1bvrFWe/a1thBovFs2O3EP39StqQGMw4URw/5JN0q4iERdHL
1696CBzooKCYeldl5gG8DZBGwfwMb6TyBNH3aBoxMpaQLTVde9+kogV2DoNHC38pDnVA4tpKu7Er
FspU4caFu7XCYBFQNAd437A8QTbiLymPfBkXyOAn8orxSK5MjNFt+MaaKGCPDGNfpqn6BhUpc9lg
cjFsLvWIXizfXgGBvFdo8XZzA2yDD38D7vEJc+7bxdIISX4ab/rLKF04hTfZYwSMZV2xqgs0zX/R
MY3YgApnAzP8gjIixIxjdhHJY2rlr0TkhU347GLuEYJBUMKva6CbglawTUm9w+cTM14wpIJFHPfP
694E8Bk4x+ig00qGvHZc2h8QyRI0+1nOhPsUhYiiH8gKEjhwu+D4z17qGaC0QuM3RDsRzl30Il+8
ZD0ougSFLVvCSjETpkZ51ZlbmYGIFX2/Bu2gQ+u0Pw5ZU+VVGlrSubevOf7RtrUPNRe0+JN2C8Mh
kujSgPDsfLCO5tfCxoftSYGRTDgANeAiG6j2CQoFoggu9p+OiLZTDY6RMFMNZ2DjgF4NsM2/Crm8
/5JraOAzILsq5gEnFMPZnsNsebzalKyDk9dzmKVQvKgZgarxe0JvuoYjETWDTBnm1CWitFT9doDt
oDYVRr0MM0Xmpd/0XP55oMY96zdlSAb+2be9tfflLkehM2Uc6N+dl43pRzX6Gu1r5GdmF75dbqpO
fMHfsoCYQLxgNdtv/oyx80KBdgCuH36OnfSutAgzfXNHvFKafFcjyLvy7SFFKJdH3iwTfO/c9rY6
2i7DLzY7LGJOZNPhYdB/imHR3F8vQzcNqYw9bz0B++v8rfrZzA5nKZZy/P8pWIcgKuzep7fw70Fg
ZSWrFceqSKqRCr1jXRqwxeMDN/qHri5KJxZ7GsQXBot6TO4cVu7NniXjgPTq1rcrJ46CPsvULauy
pRACqzdgQ1/V4xQkb0zG5t29/QA9wjEx+0tDMG772DzO1YuLQJMiBg0R25tDRgexQAe1th7c3niA
mUN8H7WrPe+9E4+EQS/HUm9wS9OdiYvBPdp3arJUA/RSO5899UFINPR8Gyfx7GiT+s+E75vC9WwO
4Wi4WMniOO4vYIXrutaa6Xlg29JpiEtsTEir+V+oZ/45t4Xpi0Www4GV569CBdEb/CkYEtE3Aa9S
aT0umSAyPvY526k77ivgOP0AmG6RPhZFVwxn6VusxgkhQGE578RWfwsL+VG7aTo8Xu6Vy79Cvtyw
cZJGV6gPvGMP/jdt3csNOPsUyh5SXYttLrRqrSUkswHFH2yvzmEDexsdyGax9TUYCo58qlGM/Hpt
xk54R2Z/TWip1j9biVnCezw2qNNdTo81P//y+wj4pQMu6jqXfpVSl0NPackQAzHvI34GmFnI3DUM
SwI7lBtN01ggPniOafa3wieAoQMoXaDosc6wgQtfAO02NBinrXwinIiPm9G1lw1NMgeDNbL71VCV
PgEUbcPIDFqP9T9OdoGXwyEtRRTXOVaYejxPf1HbPPMHWpgUMd42Fyxh7KcYGVEkqDmHT3kZO5t7
ol52K7SqfOqLdW6hwqiKhp6rWps839hct1amphEmZeMDF01UCX6OMtNhY5J+Q94bKq/h9L9NOBLa
J/5rFHcTP8CctXKZzsP11kC5+g1cpnEWcqsn7kA/9ZWfZ+vCJgKTT2NKitmUHntm3P3OCMezzdcV
tjT/f3FSP5ecAf0QhPb+T5Ce5btiHril/GhUxhuAET28syoaBi2jAilhGjLyVu/NMq5jh6FT4vbJ
LeDYjvCJJllWYQNSdNGGv3yvZTf5T0JyZRot32iyCzbRQ/jKJD1xILlVuk7LunDpYuZbXnkxqefG
0sKNjHz/I5SMRPtUUk5ffo/2k6BAKrzUvdNDDzUwBT+gnAJ158nQxY9iIu6jRwAFZmaj6XK+l+xx
SUVEucudilW53kpd0Mv4Hng2zefg8jTMi8HQayoF2vmwWkOI1NoK3BsD2L29pcxq4YA5CtfcI26N
Js/9IpV4eL2o0gjhVjYqs4bI/gwR+qm6QbT+M0o3V8dar7lc5i2252UJqKt0O2fmzL0mVwJW/qE4
EUtqO0G0M3s+77/MlzgYHBTheon6oJs2gFIO+Va7PYVfxQuFDRRum7OH9ncSn3ajKMRe0JNow7FK
+C+LHxgYWB9bUOKMfqDankaZRyYPqfyxsnUNcqFIhcyG5K/Fk6HfuUqXfsM2Pe2kOd0+NcLDkvVu
jBWwocu/8GEDY//EGV6CpBSXWu+0jIrnUVha6srlCEXMg7jJPr1YAo/HqUfkr6zvA8DEMtDIbIGD
tkfArjMsNz+eoRXT+vnVGYcBYjLLBYlxX8+4zCRWmfylmflKwrs4A2ZUETfv9jqDjboRSEKLKwl5
BCMq/P2IZInvemGXSTuMLbwcszHH/1fxDYSS/okFmlhoAmu7Gid5zrV4YiWEFVH7Dq86YlYO999D
fMG2ckih47RQ7CxkQzLXxumNZRIpu5E9G527t7SpYUO9nTnAUMw4b5A+Y4koru1Y+8nXWitUyeTK
D0fanHu1inREPCaVIeEiHUhtZGUfg7RijMPkYU3OZ3DThVBkQP5oy2pgMzIIqGKAnmrFIO5nWo6D
j/l4Ms4+7gcLmK9uface+jpDOb5Ctn052GmoRJ9BE0jhASCztaqnGnekMYLOf65DJ4zld5x6ssaV
0dWbLKvX0qxzjhi5v3/VmVx89tg37TQreINwKqgTqlwQgHHg+7onKzck6UjkRJ55sSfBIkVgFxjs
ARBvDgHopcxi/6k/HzxqH9HdEi0Uv+Jh9mUHgWrR74/LXgADzgP/DIjrBfAYM/nKVvdG2YSsioHU
NTycAn/1qGMdDMYBQQVzlSkFOEOPi88RALXTPWhu/zL9btsR+Qf/gFlQlc19vbvRZMt8FN6AirmJ
I0422RYrj/LEPLWYp8IZb6+KwgwNGWkLeXyLlPSLuLw12PZJs+yfYYjpC1s4TGGl9zCnNoxZjWz6
b2IS1mIif1fJlQC2xlxrQ6iUw72afIhWCA2Ug9Veej7PPczWw+SvVGz1HzuECLyna3CzLfZnZby4
5aQu3t201cxx9v8FhlSDeD+dUDkHktIEWu+sMu0vNHKl31XWTVlwpEAtWlSUZGuQ+1rWIVth2BC9
iYmDPMNU50olw0ceWW/3KhZB5LjKip/APZ2dithh1LL6iJxl4gn45c56eBG8uvgL5UV8otNvmE32
oFAOVY3qYPnPSWMFSFQaBas+0iQTSa8c4tBFvLj8iL5Q8ccKC1ZV+TngvK5kGzsz3OYu9/zeZ4ib
D29QXJFc4RIfidUfG8YOiXUlo+EzdjzGDRNeO9T/gmoYqFEXcUYjt3rnJDLSGL+stbpDzU17V7XD
cXHVMt2zV7ACt6HKD3MM0A449xK0n5z/CJRQ6Tu2c4Fc73irkxtIEHa8jgZuEVWp7KLCw9mntF2m
Wt4cgpkIsg80AHFLvYbIhWeNha7K9Qg+QPzvNALyP/xW5IEC6qgFWhCZU8efewgArbMb/M/QB0gO
/QUkzme7la5solmH0fq5rUVa/B6Z/hLSTMF+4CZSJ5pdo2rM6tsz6Vbp3bGFxzSaEEPYDLW2Gnqs
sFyehe6CUv4kj8KD0NNkQoUD00YZh3lJcJAHj8crf6xvPM71CAMiM3xWdjcuT4kqlGmcEic/7sif
j0OkHIbCfhvLEf9jqE31/Yfh0QG0rzSYZ9GSnTp2GIU7g7rLgshHae3ejpSlZhL000IE1KnBS/FL
ijB9ZoOj0T6KPGjtu96f+MAp6clZXfth4kpcc/0Fwb/o2aS4S17WJ0OuYOOpcBZE04qlib0rgLVI
GxECcwQUXieOsXNt24wyUcrIpguUUUHXcXZ6adG1Z4WpSbwfhsZBJlaQvVzDpYhPUoM9o45Rpszq
8p2Ewor9NTde4fBoZtZCUgiK5BNwh69dqk2Dds5UtEkfQG/sRGwXXEkdqy1W+0B+v3zR+Kn8mGcu
Ic3ySLmAKUsNnqvXY53gD4mjOHWhiKgqqzmqG7kBnmAZrTnVr78pcCcaJ3yryR0cGWNJ1pnI/sX2
Zp8AX521bGOUfaW3KaWKquMP/nlisxGcl+GGva6TOS8aQznFQsFuFlgmeQNRbwtOvx6/Q9NGEvbj
hM1R7JOy12vhjsXQxr6Dua8CkrTTgZRIS+T86pdQjG/936Gcb8diCIkRGKyh/s7E4pFJRDvQRnX8
mdeD6E0w+PaeReWeXOKY7BbPOGV8nkXYiNS+C3HQ7auf2CU2Ai2AulJ9R64/0vXcAalZB1X5ssun
EzZziHEptqMlizPdefLpEFvoR6VJKEWz9pG2rnTBc394zX2vyQzBNIwoVLIyzp4c3Y2/kP1fBxNk
26IsOFbqC3OIP07PkJ/5gUWDUYofoGGpda2ZmKTtyo37chYlntiNycY0y7uILQgQnkHe+D4G/ZrT
DEAd4jYDhxar2L0lSwcy8OW97J4mAjVbj5bX9y8c013LtIEhrZdXhRe6jB2qTcWZN8l5WWQrUWQm
cG4k8a35ADuN8j+7hfVC0IT5gC+sjYWOulo/Rmkgi0CrZkTZnWjPjsy/KZsVEO0moSS70ZieAXgv
WRC/W021IIaDowIp/2Px2Pi2JOrPwGFZ2BqCGBBmnNxhHPjGHpFSwj90RMggYA2BsHzaF8wPVd1T
s8cZODubxS54rRTT9BRntBO9CbWUywBsJTXUrLWv0jOVLPWJvEUfkQVX+p1Cq/kXfMZgcMy41GI0
Vr3ZcK+/RTtf3jHizmPvh8HwHzjSMtel2Vb0/CTL0OgFigP15vcpZE85Wvuh6SdAksDHVyIZE+vu
OHqaagUmV10UMMzZelQwy4bK5VCz0mHOsfBZpyzD9hQzz3xdO0p5unIb3EVaTEBtNNkkOage8WhI
jymW3nB5uQ21OYZ3dftZmi2US1oR7/Lq4Do5KaRmsO0QWQEQkyXm29dQaP9hHlVhOb1IkMAd5EGI
Ftauu4Uqh7m8hC7q7m0RBV1083GeeDpZoKzFl9/aISTZ1uGjW59X0VItzDeCjF/ouhTzs4hBu9c7
PkvxAti4uLa99lXFXqkTEDeuNPqtE6F65mHrDUC+R4pscGO4deraZdEw3k7DFz+TyEn+EZv1BNCb
dKVTAkxRgNOimbrssS1elqEmzcAWJ6UopMmzod78SAHBT8x0VnDCHfkmqW4zKanI/c5Cxp7J+idn
7zNiR5Iw2B3Iu26DcZf01tWiVqqUbeTbfjpa7AhR4UmeAGSUm9RLJGyuJXMxzhH7DqXWSnCTMLhQ
xpwlgKYjMgwDOqAb0ha1jLp34ymRqvXPtaV6Sa3KknmkohnF4DG8I7u6x0XFPTjIP9jbhXpZRHg1
00WKcs52+XtaMp0iTCQyynSS8dZc8K2scEYkawY56BJI85l5kS86OfaiG7fLkN6rWdn17vVb/ucl
n3lLwnj9v707f8QXFFFlhM7XbKYoXl1g2K6maL7NTo78bCgVLJGZkfqkVonR/3hY2aZsm3WMSrg/
Tet6QhviXwVIPzNRlNopTkr3nGLyTBdHky/gpiJuL4nTwk6KiCN/0ieOWHbpVR+3Nu6mL8alZENB
YHZFFRnDTOTYOATl2IEX9gzZJSbHD6+0N/LFXd94ipTYSeP3Eq5Rj+Trwm+DIGwy0+LVp56I6uyr
ewCOAR3ESvNk3JDLttydgPYvwYVGtqyFeQLlJfLKUsPvYYyjC1/770n72mBnO6gLqI8vOYEkJn1N
oFDAJAvsslnKm00E1bWmf7GwdSX4Fv4TycllqLlo7NlTbrvKQpyb/oiWVIXOvctpmt25PhSXi5wf
aCalAFWicr0LUQKyl1s/h+SEx3GMekzciejmrLi/oqa5W1MmklsE6buhEfHGVlAzsxu+VQuixVkK
ut1pwc7GjdcV3S/QAyAmm8XKHOm78PnCp//waNo0ypiVxleUixRREYNFiWv/ZsLzfbG6IkTmDdtN
GJiSbxH1hs60A7l7wOcpkWYwmHVzyhG59LmpcVVGPDY5Supixk00Eo+fl07+hKNQNZ1QH9mt+DbQ
UvnbSdxN1H0k84FAI8+WTmptthhxEeRohah9IjF15Nj6aQwSBO3H/gXasu1M3xjo2Q2GJFsjpVGO
CVNst8LM8ovUaroxtbARbaxvoYONjww/N1ljbOxGZhNEjiaOlU1hBiCZtwcupwczFHfzuuJ+fsnh
W1Fk+6Fdwvsk4EpmLktLdvH7/IMZ/wiVB6JxsGWrfD3nqBRe8vM7Hp2ti5HkAJmj1fz3t/jfc6gW
widMhGakLYT42/GuSV13C6LkFcsY5q5NuBaUzmPG7kEgzfUF8+COtVtUbapsCLimroh/vI0Qbf+A
kixfXSjxkudLj6DirP6GqLtjeBXy7H8toCklUg8HdctnpRAbom8UlbVjogAmQ/ZHpSw9r3Jb6LA5
z+OS6Be/qI1QNeYPQDuCPo3mQt/2eLy8+ko9t2wG+stgA+XiNKHpYAIorKDmnYL+ectXrseTSy/6
lR//u+c9h9e5T6wgJNClw/Y+AxPzVG/wwX18sabO8oHMwqEMtMvo7nQTVuNcGbsc8MY1padKu9oL
7yNgCaoi/JRAxNik9LJFHZYwW+2etp/l4oQhBIOuKd27yxrY+viMziM/p8Wd8TB/2NlRnZE2TS9+
zd5Ecym+miH0WR7doPYDU/frjCZTgH+zLq37Qq0vbI3UEljI5dovU1ka3sy1TlY87XhxkWdDt894
/JR0wXsz+i2cqpEj9WqEUAmR+65w1V+vfuRKp6J/XLAXD+VxcnBaVzEbRfkTs/S+H+O7GqfUnNY/
21BFGCDVNoIpFT3MYUSwEtd38mseJh9qhz4L11f8kEPtcsAOEaryY8x40gBU20bAZikJ61oZsHfR
/dz9l7fHkrZbFGDJxrcc0lNR4ofb/e5nb02ZqxgzIgWYRGrQDX558smZpZf2KbrIEijrcZJ1qOBi
LHgNVsCQIIkxateVLfzgcYdWh/cVUnvZfuJK6rK2J1rlS+wtVbUpU94CSUCqitlo5qf0OQy0QJay
h3RC+Uz1ClLtmtQrGLR2ZhFWOrTVIQRHSRGoNf2FTryxz4wctv2GNlGoj4O1DCxEqxmcTMGW5NWv
XFBFNHoCDBQzNcsY4Qd8RKgk7w2bEdjEQNAURIk4PYZOyfsFURT6iiSpFpzpbiRUmajb8TrK2e7R
Ba1+wNCreneFZyeO1bdHgnp7jUDZSLnZJqB4DWLuRuuXj3GSwXkgQlz9y8Y0sEi8Qs9HE1F3l5SY
kUccWR9sOAg52u0PJfrSO9ldGZYEIERBNw+QWg2y0nuX9Rw6J30KgsMxMi5vvLUQ7Zh59XFm6FPq
hCaFm3pGYVx4qhbPxAtBhCR4ZX3BAhJKjMgGcwmBuEbLuA3j1ObV4gnhbIRpU9ZhtzrGCXIVdOwx
UGgM4L72DsfxTCC52htcuAgmGTyxqB5cLyrjFvr1HZ3ZhUAhQZ8RVwuA2UgwqjmXakUykkSbnEjj
B8khZdrxvMmfRLB1BM/aQgoavFGDvah41mwOvi+8cbjAyZo5hLmXnlecGhS78XwEbcIzTNDYghOW
dgfXSxp6Q/XsfGiHxrLbl9l2DUkIIu/1N4W+ywTb50PP4S2zWudk7WMwUuNW9SVHevpwL8anyqcn
D2mznM1YyBCo8CSUmwp10LWx8mLUEPZOtpwNtXp/MwSOQwMJjkrmGuFqzvILpAYFNulp7lU5mU1j
5nJdh/wPrbCj7Ib/EE4k9VzEDfTcviGl+82wbslWBe43A5lZZRPCk7gIwPglpiOQY7EaiLYhRl8K
bxPMMqkLcU6LnVtI2/ktdCxQ/XyyIOqNKpfGykaHEzfU98vd/0l8n3yfBPX6AEQ1xsM+w/I5Ycyh
7n0juRJQA6BPCFTslA+ZkXGIGmqW901iSFu2c0N8fC4Ph7FuWK/YNOHD2vZ7GrtyR/4LAGMiL7Dl
1IFEGx9EsFAXZEHnluFP71/FGtJXPNq4rbVy+zWAN+F09C8R1bhGgG9gm1fZsxfSi8dNnHHDu8CO
TidzRqNqEC4QPnUJGHfwkF0Qawbl01jUxHjSnBbodqqT6qjtl4PVx6Q9b6k1KfuMC3Twk/qgpwIk
nCb5AWjEm24vs4dfa0OmdnenlnT6kNDvYiq0gOvS1NoHRk8RLHPtWAS5wbYCTg2zIaunHkhZUzK2
SaR2M1lao4tYSxFG50bvHLyHUS6Lx/XuXTl6SaPm451M8bh1gRgPfJ/yzguUIqO/eQOighJTnzsu
T+9+nOCHdlgu2kXviDotU1y7XwkG4hkBD/DTtXQAM4umvrvPyDGLq9U4xiFAxaR+IsyJbMF/95wi
Kr/OD++3d+qwbjDG2Lpfi/SYc1VQ2AVLC63lT/YHiQkmYsCM2OHcGY8A1Z4UJOCinMKRstYvMnlt
M00177oq22xBp5QVYX7QnJL7wugeNWveSN0hcWpxn0TvUNcK/2EUU8Nbef6uam7LCePvDcOpZKrF
C4f4wE77WrScwFLbky8apmSQmA4HUPYydxoosew81J6gEeIdinbX+lBcqBv5Ze/9a40w5VmmILin
pHUKXZerOOXiJDqMkja+w4qrwah4cywa41UPzbJq4gI9tRcgJvjairI55wJFRR7IJ71no0BXNafI
CKoKceK0QvqWK1otUI4ef7z9r7EnRcir29GE+Q1SbEX462nPYTpN9RsJikWNUTHzL4aQM2aR+Hhs
oI+J9cyS055wDrYuXrXdZMBH1zpmMMJcr80asGtYJOfoYUn5vDPKSJVwTBeqpxgb4x8AFjeOz1zW
xO3HCcycIaK3yZpH7UK0ZG3h79OVUBMfRS0nMPJiuZjkwA4ONnvIfF2Ducz1h7ywbqz1y9nKNPk/
ChY8D81Lyk5LB10t4EEFojruQT2aItHbBQB6DzQUM40Pfsy8aoh/M1hMXqg+qCGRyzDd57f0pziC
8tufdCkFxalLrxJMWdtRSc1rz4uB+RFxjbz4EXAxgSr9jgLsCWcgXjwzSIncp8MnjzpTGqWTYZOx
e+h/v1V65jo7vdHc0Vwgy97hn6FIpoeYCMGoN3DceIa+LDs5VQctKREtWjn/p5lYB8K+eqiAcCaN
2Rf3TQZP0xIdAAPkhnACn7o6nP65tS6LqObpecRQGDeMt9SACja4xLPt43Ui8R4hGADyEE7bYPB1
gcXoR3F1n8llqkBgOosgptNzkbOLcA3TJsllssmJNIxwBnTCG/AJUJGUxzGMwvxwPfVSh8tiT2p+
PTlZJqVXbLEc4y6By1kyUhCnIz30owUvfn5fW9NjfA41tWvUuPGJhzyco05JLxttXa3Zyk0f5Jzw
E3DyjqSWyZ0JJBca0B7HA52dlysNnz/TPFLZhlhhAR2iTgCpZRnJgE12MYrZcGYDKNzRgVmauIeW
pM8PYPTMWxtfxu5Cwrw1CyPZ740j3N0/6acbvqFwK5L0CXmiMnpCUj6KPzY/0ZdrVdhvjSesjZUR
v59JIWb8i6QYCU4dk2BIKvc5VvcpAJvRAJ9wohcTzu78MHJ/s7Tlk3t2lTKfyFp25ZAPEugigNMe
TmuEnB7ah+gXgKwe+ioqiHcaKqogfXC/obL5pPnT6nQpvE7AclOWJqlzalUhj6Oaf+pKTV8JBuz4
XawEn2kvvdn9hxMQNxG4JVmi9ifZb2f8TWWfrWr8lBg0YPfdPMY3t6WDrAclPbIDfdlUQ6tRWwY1
BBTmIXQcDqKeCGWpJuhrv18A9KLeKh+s0Od0tkghFjdz9Ty4DlZe3cfHUD/Q5k+fs3mx/bJc9Ea1
bPxYmg5uhER1fWGvhJs0PV2Pi8K5nx+/M2EE/TKAZWwd492iYi5HXM5f1LT1BSDYr1Hmu2raox59
EPpxkuySdgjkJJdVwoUQrSmW0br1+91ao3wEG5NfUdye3OEcXanG1iKiqF99L5tVF8JtmCInE4NQ
Uo3Aej19QTwyGKY6a0yukR4nGmLNQBip+Rp0Dk9YA9VSAfPQkZJzz8Vd2aFgAF95O7o6QkclNOr9
KJmLjQISaRznrqV4gaUepgtfSW5x+rUPA4B2ChYxAamY4+UWT6a5YMw05axPHbk8Q86pJJ/M/Gu8
VVnxe8uSWopmJqS4B4ry4R7o8MPT0ynxGxBEcuGUeJHaBHU88ziQ4CEQeOz/NPVQyGc7jH2xRC0B
Zt+IoBS3/nJNrpIe9003NiJvl4snT/+aVVp+PshdAg+kGiAWVhzgPQszeZ+KiqhZgXUNi76VSb/J
xZDmQav61gkkFn/OG05Zp+zO6Odl7AHxJsxIH0XNd9wZGMvhq6A1kaT2POC/z4oOUfP5p12IuWD0
xk1+XMqSR88n4lq0RRZtYKvuvyg6BJ7xlYGJLJD4o1dM5pPgW+RHGK1eDGBrEQL+eKHRuOTQDNmG
mtR1JUkXJFJifnFyDuCEhmdwvizCb8bCcPjD5oD5KLd81s+mxQRnYw4fiBbCSmmR/tI/rrlG24kT
d6UOO7Qq+wvRZNFUV7PIOiDTLrUXeRBdrp3NynD8Jl2EjYMCMkKsNwvGVZXX5cdB70d/RHKrlOeL
39SvL7yvmj+Iv2YJJL+Ei672YTVN0+MK/S73LIC2+HdscnmVidqQulrUsjZfwSfV6s/fT80kT4ix
KgLdNxbmQjbABs1Fg8nuX2GL3HdaXsbtcrpusCuN49c1c0KxxlZbPO9U60wWtxeAe0BljhP62lrX
TWe/IhaqerxZOZEk+sDLzzKmWN8mVTBrIMAEezdA9PdfK4w+mKFM2gwb09CLgXlgtBZRrl2ORuPX
AkrQRbn3iRS448sGZckxPZPbgttY9cVNcgIQXFhuqe2QdzNM7mV+Sasml/HpfUGnHdmowvwv6Csq
MOjicHl8nfrSvEAbXesV5FSPObQBS3lg4uJJKSQyL/gviB3/3jALnX4SRnnkKn7aG8wzuZTvcTfq
+MbENoipaRZVqJUGhcXWOP1BvQINBuLlWLlD6IW9SCRXiI4TTipmGrGhevdfIe6wug5NkYFzcKNW
9VXW6jx6gDLQ8f/1fTJ8QT4GgMYC7pGEE+lC/WclLHgbMsH8euRUTlwYud/RW/uOxd3nYDbpbOoa
LtQzUFqKAj6H7aRLEjQUpBwmlF6nu1y70PR/HP9/GSRshk936RUPLSi+ab5YPR7EUDWIrUe5zbEc
mJO6XC+EYOZVyfiDRH+pkhQlJdGHtHRhGkH5OuMYtg626tjA+0w6MJeR3/jk/G3NrghZx22kxGIx
wcxrmMholTXRNcBEgAvG9TZ4eiNuO1a3e6IwQvLVvkdIm2o8s2lx1JanYOlxaN8TW0Z6Gm/F5RQa
7rRiMki5Lfdci0FQUPTsp0+m/sZxvALApK+kaQKv2/wa68ryrDMNm027eLi5lv8DilZThivYa4zv
Qo5QLK+r3rlmwFRe8hGiJs3V9ubyUPBDkoabjKr3wyYV9uYcSOOtJSPi9sUOBglhqy1X9KgcNv0t
7bguzXatfpUR5OVhhz4Ixi9LdFkTVSZzSOiTUfmuMJFe81zxtk7Z7Urccla5H9TbdPGNWzB6m7fc
xOW08hDfDVxHxpcBPTdcpABQ0cBwgMfkDN0c6zhClLUYpK1uPPoXPKsRw7PR42F8UYD5FNM6DE+f
yGvPVSnHze/HODiPzzmW7cvKm2crEriPHr+lKLzeQUpNbgcKS2o+NhrnRArF9N5nPTegypJgcA0K
O7KxLyDTvM8XrD2j4hS5UGoRhTpVXmnviOHa1OhS+dleXOBvaAuPBZzfuvW5ccPM+Z5sAIQGT82L
wVJqcE89zAx7kwN2dYbsEqqYbaTbXiFZFzgXB7UzIzZ5wrtf3CR2AI50M2ndp8650fbSC3c2T+rg
xb3DvpDeqgY6ebldiEX/4BQXXhzVleSiu1BCA5+DFKCa1gmbjt5BVkbTAt3Cf2BweqCoZMY6iXnk
aXDwLyvB2ucaSpNLFVGfPFt/ueSE/kNWgq5WSHaUBgeUbW78ss0A1RDEJfo70Ji3KNokajZSjC9f
BvKX35GSm9DTRoFkqCuiieSAyVJx/s+uRvLEu4g8nsRagG2cLnQWI3RULZM+O5W4WUM45fsyO3HH
8nTMHzu1funAEA+8k2JuLn+Y+0Vy64CNsO020vTnF8o05GIp6jU/I6RxdGBene43zrG3XMkU+XYD
o/MKEJNtIDnrbQ51kRyfru59joGxTfMt12NEBztGjt1soP6y3nkkiQCAEVMyb8G2+nqJN/+aaX79
TnmFcx+umpnaGZx81xu8BeIDl3khMYEPYhBcFfnhtNj82vK1Mvk7AKawNSb1WTQ8+sn5V51Hk5BK
VjylaEonerHwvQ45Dpqg4IxlnS8JvlsvonuRqDjdFLgxouXZ2x1gHEtCGlIOnPEc9PntZ/wllcFd
9hHTiKpugvev4XLk2brZqeI8wUIRe5lnwSdb2G15P4QJpLqwH1K3Kn3m1fvjhKOCVsBNrJvFCUVq
sUEheKB81QMXvm9WILHysjkrB9mIV+XIDNl+93lM1xMsUK4B472iR0xhzJ3bOxKCd8mbXgPDFIPF
OGPTGZP/w29y7/mHiOZnsHN1FvqdTWeegTS0HJyLRuyGIjwF4XOVGG9+PBCjo/dK9SClfgHm4hEm
qNQNk9+RO4gN+jX4wiacjqv9vFOnJINToV14cAS50CpsbhMwol1kZC0p8fqi2WCgSuyszcZp6l7O
B7pBTgd2PHbkhK0QOfpLjdnDJqn+PtVFAwLRS5vJ6UUa8nBAZUoKl5cWlltgYS+OXe6arHnYwggt
3uM+qq4Cuqq0BpnsXRqjzHXyywAOvOmjrmAytS181rP3Os2jR5bgPkn+9AE4dCBK7TfWVIhZkCxA
kQiCt0l8K3fxeNpVDpvCDOjU69XU0xKYRwgpVovZd2H1Tvomv8zMq5Bsjgsjodcb1dBtd0xsmmGU
9RaDXPZ6687op1ld7ivJzSRatWRnKB5E/lrBsGKhKfvlC9c8WmpeBDAbryQmwU9nchD17jJZznO3
eU5HofWvRQVi/Zsp5hrvmsjxjForXxYgI5m6IldbUyFQtamDMKgFPnes4xiVCIWixBmB69kCT39B
+T89rdpaeR01jBkH9QIJQVeVsurWivWLI8UvFLp6LgFv0AH5nI4rYRfznFALxLCTm9qYfBN5D5w3
BbK7bt2d0ch2rTRxDWJvNMlhv6K3iPed+fJ109E8/ZuzQjYDuPbWKinTyhfIWhVxJtRoPux47IWw
FdtFph7ufnh+0rM2N1NhHf7wI7b18k4bXohd8QscUfJ0ot0tokAvB9t78IeDyjrQ2shzw6bPNOA7
nNqgyjdH3FYDCw88/78Pk94oDyNB0r4SjmHAPN5GZV/GjP0oJDuTqEslLKjxeDUWPu7ZovAYXuxN
s6OLZAoYutYwrukL2oUQ2dMR3NgZWtiJDp/amioannxi0t7CxHkqg4Vq4cz1DLNV7+nF6zAAUUTv
PLbUuL6BFA6n0TbNN0pbrXSbVaHxU+qA4yA0UaGHFF85U/sHRStVOQ5/+qeMu9/lsCs7uCBOg5wM
kd0/aSeb4Mu70s55ecbudARsgNWZYHdNvDmOZJZRVbQLXpM7y6QLUWl/rCSxMYekT0EU99PSE2oT
PoBwOEvIkguA+8pdBpIX3vVJiQJdf6HU7t8hanc01O33q1araOTFwLsIbwnQBtSsVa7Wr57/uw4d
F7/lLW+qrdprQKDeMGfLMUsvVxGWODwpPpZukYEtQdKeeQKEEeVf7c9dd6N9lfVnfQBQ13p5oRT6
wf8ZTkZdN+AIFlgNvB4Xrip6IUcfq8NA5Gz6wUMAWBZ7TDJl+xbY8b4HSo5iT6bo+6Yy6XtMZfVj
iK68kwTFpl8pSSdy25MKfIj1dVd4/uSMSc55Vmo8AwjX1meAoaFIKhjAZKoLA/1tYUAtUN89LYQ3
7h75hJizYbfMjVusl9i0F02WhC7+GN/8dCNiyD3dm7CnOWy+utqHwJROgjLFxbSzVVpyVhlvvKdW
hKygexMrvZBAITrWH4ptWnntPdfDoLMj2m/30wpiJPH/OywQWUNe0c2wMM0GCstLas5MDfzgpbc6
eWnnUCB0ytMGY4QC/HdNvTaBvSPJ+8HPD33qnTV2LrsHiUDrH9gToExRfnJlemKIqYm6e8fhRr58
OX+V0TKAq4qSt6r2MjKplxZ+z8bZV/XoeyjK3usQDGzC241wKeaESqd08dYwVghFB9lfwFbQbykD
8Q9WTScCIJdgWdmQ1QE08BMEr4Io5+ji/n0B6e91PW2ojtySH1MWgi6raVtWhtBXtR45WaR/04ay
S+8WIaTuzJMJYCd4++wuQlVKUVReZG7s3U9X56OGp9OjM4ETeapDIb7y9Ce8v45heMy95wPORsKf
Ok8bAYEzOHfk75hRFv+lgWfU8a01BJrLXTiI0FE7mFpvNFQSiJuwAQ2zRw6ADcxDfRtHX+jwkOhW
lBMJbnSyODfI7qlMjY+hHRYXv4OJIB9IloQClGoAw8frhceAQw9NzOXq8c5vconNJGzPom7QEujj
qjBbeVZhzgjG+qB+J9M4Jp2JpwrRdTGPe1Nc9XlKa4ApqiVH4xe99/xBpX4VxAXEj6Pagg/4Ly1B
lgSn1CfSNKjvcTdeIpZreLuCZ4lamPBZFnt/Qk4yMxy7h64BBMYJ/Z79jLCd34Y5CaIaw6FhRS1E
ixeDggJ026lcZAoB3pE42qesXydswf5xl2i31CX80EZAF5UtaGVevoRCTUytgMkm8t+I05OxKOUr
1yXVNFTrKN035tHDCY4XKgsBjRHQsWBeZTbk77GpawtvdPbBWo9vSCaTNC8q5bSEGw1PEdhoY8sm
zOi5gnN/y4SqwWCKwPT0oLCYDsmpvp9ZXQArYcN0Gf6lPLdltBAOi5tMRQoS0Kqy61WJrk19sd7J
vgxwSvZ2iGIUxUaqVXP05ftpm9nhcP/dwGIzSJzRcDn1uoV6wudDsvc0Kss8dGcQuSC7hcPc5YuD
w1qZ0g5H/3+hgsjXxZqlSgNXTKq2gD9Ra9LKJaS3c+xcupQIJil2nltjNsV0Z7RNWWCQRXJ1gL2u
kbJhebWQDbr73yX5tN7r2foJkodq+FSiHIDoaj7CmZxvuEh3TEuu2GaPqLc+DnrBT52qZsBALXus
ouUUGpXClyiFsY4QMdUNzZpGJ54eppNvOktiJImKqf5GKEGA5sE1qrMSYGi+O3dEb3wv6osYD3Dl
wxd5bUxWYtCG47OnjSDZqganMra8mtNZggpKP/Z4y+fvG5bEFTyI1tXPME0F61psH7lJe4Gkecuy
CpsEvoszxf8JYmM2w0tey2XSkd1vV7FSIf+rR0ZEhMr+7sHHA7GfJluCBRoe2SFl80bTPr9ejD/l
hh+m2QlwrbyzFuBT/YxO6nE7u8700hOUikBkg2rlzWPWPf709fncNEhC8Sv/Br9vtN4YYcSbD567
gqinr24R5Tw++3Jc2oqGpqMuX/Wh9C4RLzo6whZxTYpNOy3Vpa76Bn1vyUxWjceBz373j7BOvrMU
kzH99EhP2HY7ke0kbG3micLeu9emRhRp56eLQjycIA3kpiYpcv1Kcr18n3hIzgTDr6wo9obOMwS/
w1SoB1gXTBYKBRq18ifSI7IRTxHsHGr4ebDWJWe4dS6Enr4fw2SXSRnxypiMWH8TJX4F+l8iTqE5
41OP+bfji07XiRiiFVmsu8hia65+2i0BzGW3dpShKKZiNdrzPyaj/RJyoEQkwoHXccXAuQ+Ng+gh
UnRhzSYDjhsh93ry34EB4qfXznNWEBw2JgLPKyljSHwvHRLh7th4vgjblQU9ujj7oEYyMsqIprZ6
tR3j7hJekWPvldifL2cD3aBtRWTTq6/Y7z2E/s9xFexLIFwiIIPp+darrngIkAc/dkayKE8yvD/O
7GZEASn6LwuBREOGxQQpXOSpSYwI26KeH6BaBDZUPJUoqXdtwvWwAcAHzNm6Z3VhnZfm/Bt2H5fJ
fTmO8WEQ8F1p9FL7Xi+xyKYZcjwHASItC/FuCOOWM3bRPwdlezoQ66wvC1iaBwI+vDZbHToOVHwR
rv2Hz9egs8fvpsyUA9QJ8+lG5XlHMezJIPcAcs5He0wK3usosymesPJJJ+96lPYJjXIVKNVB/GiP
u60efnba9+5G/0lXhWaRZwozuvcpvolCctd+DXDLPo4cUEnRjt+LkCgKTtfhummnmWfP9FYzsKvA
N6obV/S8xUp6+2BK05k1KcTrKH4InlMhkkdo69wh3Fbk/jYdhnTfEXibeMXvg+Bb+2BgwVt9iN8S
YMHBKjqsbciN3ZfafTBwYDZO3rykqp6Qfh6DWw/gDCTjpRF68mA2x0/t9/RbmZDzRc8jAv0XKcsS
00Lf8McQLR+21mZFF4AM8IoEpfTflZCwJn+Oy7PNfgPz7+gH9ceTZmp0MVRoOCDyiLq5x5VFRNZX
JG34fcGR4MZ236H3e1u+if7ytVraFeyf1EC6/ZDhzrljhYZzD6vi0BM2Aqn/8Qnpwq5Q5mxQnHtK
SqqRnjOp8quM7V3x0dS0+0L8GkT63Vp2cEJK8PsfitMmlCqIdR9m8xfYpQI0bKfhaFa8B3JbjaRE
W3/Otmx+4exXDlidnd0BswzeyU5SwRpLzW39bWyyFHwvpPc3OJZ/uaJDS5eaOxHzDN7sf0pdoV9X
Jej6tDQ1HO/4hvMnz5sPcbxUHO/Bh1D6sAf7gFudHe+33Q3TokNqi20odecR+9URmAqjTHZ5Uz0L
KU6cb+Jg7011d8zR4+RvDB3fSjgcTtPqC6u9cErjBTvvtL3MOaIpUrY/SVbpa9Cu8oJCrvbxGRgM
R83GE6HmQUlfbbu668s9JRAk+YAzP4cxfTTWrgZHfkUdGHWQeGnxU/tndqDGsbJ7hs/khZsYZJC+
KZcHMGeDqNlb5zg4UfxOWFa+KsxnLUsXoVeTuHVkopayl2CGNk6BqdL/s+qaYZGeResM5dMhnPtl
1dpL6qDUBJbAV/NXx8hspGs9O1OYHrAvB9ljKyXGM7/LCQopiIvy9y/H8TAStVzCYR+vlk0Zb6Jl
zsO1ghHVbCLSNa+kCrK+2w0gHYaKV+UhGHd64f8ZSrRNFCArPVmETde4H8Fyvh4r2oYVSs48fpNk
JJG6Tpo+Acrsd2GGJBHGDN70tqoNrxKMw7IIoi0fGYQl1hUYT4llcazS0T1rGJuv/xCMx0h18mWg
ca2MD6/8kQcqQEWSYKRcAkCqZn/GY7tRwvLcR3f0/AmksRfSrmUVNGe6Zgf9t/orglU0FKayg0y4
J14EwFgARiOIaGruzHZvfQjbBq53ua2SHBkMpCCD1s45o0Kvd6X0CrqbH9ej6z7gclJFDsIOiP66
77GCTbUzFy22oGWDHy3z9UuxKdSL4cpVmrLmqYXGVJyGcJtPkx+uActPYBdlJgb3FQrBLFRxFVFL
eCjZiBWI3OG884i4XRqOI0hiXoYJmkOqzT0S100rU9XcsB36evU1buU7YkI1r/NCqOrUdhkOdtC9
xmupNkoUUptmiJmgITAE9KUu4ycVgew0+qgiZXU99+/kbPOsUfVQMLsJcqhq+ml5oWiqZR9vH3e6
3T+eK6rrtZ5qE6JXspDhVQWttFCp4B27b4RVquldl891XhmF0qyQWH77Qe5CZRlK3zjam+QlIgWy
XWovz+tiUiBEa9518sETuQk5Q+NJqdRpM4vsIdbv3FuEz54Q8LOfiUVOu6tTT63kbazfKYhjoeEp
TWw+Y/aO86z4IGsBF/slUDRTkOlNvB/0GLkpF30BcsevaQ6HYbYtrdK8VqilUzhKhjeUJ3YGKdTB
uiSnl0xpglv1TAAAaYlSB1hpR7hJkWuxX/5vKVqoDlFOast3jnUrNccgD0eXO0s8UpyHvjJVKUw1
V0w32Hxnr9K46xoSWOKd7Z+ckIT4mQJLXm0iwllIrz0+sK3f9k+jzSX8TPNWs0BqvmHmKgA5eT4M
aq0WZuAcXpt1exxB8N0sUn2eVYEcbH+W+R3vZou4sscayDCZtd1Z8OoTKdl7Famqsb5p+so3drzu
1uI7TZ41MdqgIUQmjV1Fli+9e3GYX70X4D7bf9WbN9bpnHvaxh2Z5RuVwxyppNknNf3jBXCpynbf
+4TkzZ1kraCjaQnKE3CiCrkmS0UEb5TmFknUo7JRbr7MObMoGBYYPg2RdtwsfbOBcQJ2Gs5ZDUlu
szbFW2rpOPoa/dcSjtkGHh0hm2yGrYlAEdC9WuT4pK5cunJYzkbOJdSPAkhD26P2A3Allo6CMszI
vxfNE8jMA5oQ5GfoqdmoLhAb2dWbwX4w2ByeTiSM6MvL9WSnikQghIAkCj2kR3smdLEGT4Uky9L4
pU+n0CnP3/noPBYxWMLUX9Sfy8+0KRkrUuU4OyzNJWrmdzcp3co3seGUYNcN2m/Dy8vqQXaCbGRG
hJbMmc+ceOHRBz1vZDw+U6q38oEeGtwi9flHVygqOXFVfihbppIuqKGVq7Om4XF+0dCgTVa7neNs
WoIJP3aWPUg2aNINLlHG+59FH41jKSU+xTpaPg8gjIupJSHwImISwGifFq8drDNcgKPoXeF+Evrq
RFMbi72CkZ4awK/x2wr+Z6JziwnahQG3JhcUdwaIZbSqUuTs6YXqnFMLPSy+pyzZRhVqpiHXsHbC
wN6HqHQDgxMFwO3ultl4emdidShL0YYd4LGuA2xs3X/bKr4chQRRBtXbxC5w6E2Yt+uI09P1cRMc
Ie94RCvH1bmqjWPsxkSti42xAGFRee6NTdDbKd8FoIkkOTiafv09Cy15XViBJ5NvCBp/1sd2nEK4
wnPg1bMQ33DCLbfF4aJcYq5O0fHY/EW+4g1tjb6GGoLj2eDXTMTWD6ZwJ8s6PdCGVaxkyxlSd5Q/
nXR7RIrH2Ms+WLtI1RnWfsC8hcqhwFEPDZs4MnvwuaO+lpOQ9dUQkwwsLS0v7A4uyNAX3l86M/5R
d8CL5vQ6qaJ7Emtp3HiFhlfB5tkEasly1jUn5mhWN2RvntgCDVRiUbEFvbzcoJmv9NX08DJfNoXs
LBVXkTxPZyGNnUBS4eUFzxGGPtYjbuBlR386IsONCbETCRiPn4t5cr6uXz4jTnzMZc7FdvHgo0zg
Q3bcFwoVhxN30UCn4ks53DpyYnGo0P4Gtu70nle5Etu+fJVBCzjT8gA85F1RjWFGcPiO+OvWJqIR
oDMQ9fYYIA9TTvA1Fw4szzOzM1vZy9dtu6hCeTCOZu/vwtuggDD5MzmlbOZTsh0GgWNdqBxwzCJm
Y3e5f+dhY2w37JUXnh95OnkgnVMNMrgQmGCB8acFtpGnN53BcDVeQVXo+MfmHVTlhrEEwRFSz8bq
gedFgq+EnUDU+stcuaCdAqYVY9fNgaeJr/fvqxArcdkbxZLN2CnoV1LFtaSwRnO6072zwkrEWn8G
XxK5FungGeVsZCqRmP6yBg5+tbfPS3yorFmBXZnkBvtqFImJREsg7Yc7ybiaJLrk8s1a5TQrDLjk
K5ifQ0/WkIGUcACtu+XHC9kFolyDyUjxyXfEhMSHvFYwFMJcU3oAKZsV4oEcAZ0jPegRXUqsP5cr
PRxy0U7k0PRYunI+UrKSxpvb2FXifsqoEX69EsciUNYq3mOGakqEb8Hb4Kba2guKsKPh5karLAmo
WOkfSzpMkavKgjYfswgJhqOCN2BVp4y5BkGpRsyLi4OU2FPLwj6x/zrd7S5lDtzxkAeQfAb+Yu9h
u+15dVRrTHQsrH8xIqL900PbZmNrBXDlQU62ukukw5opAcFM5cW0eLE4Ck2nteRfiTacO7qkVB4O
1pThb7bm04OvccrHU13/71b4Y9xPoRL1pe+Kz33jlPF0Oe7O9/JBnm/8F2L6RjO+1UbYkPztBGVE
RCihpLOI8Qpc8jQ8EbZSmK+i9Po6+cqEp0PcPdXMmqrxmtJStdtdDYvhUozriL35vafafBhqlLyR
PWdo5hi2F7tTyYStcwA/xaYFNllG8Iu21b1wQ9u7jTqw+EKELGCmkFpzlk1gFCPU5gefOlfoPqd2
aLx6GV/ZTC94tI4WJ8aKd2tVJPxK5q2cuGw43QnB2OZrXZHhFAv2GYHuVT4iRAJh2XNQ3dPfLr5L
Q1TNh05cZux13Lln5FPYwBgbBLAVzVcfnoBr3z7JHnSGB58Cg+xuabOpNtM6dKANK2LpQ5mlSREC
hH6MTidUHWKec5xNANsY6qy/9FVUEeztWt6jJhHlIQN40xFoAsahY/1U3+ZFM81apatiAS4K8f6z
XtziRdb0HQ6gSDiUPk6p8xaYoCeDTSA+YVNHhJJue1ZD8LGRqOmb5WLoKXifVAvclZ0SvbhK6fVu
f1cUwcOEzp/VtnOl5sDDFSIXl6Taexd69OGYWblqwdnCfc9cnmxJnAsh0ls6xoZ6lxz+TIKUMiLf
e4u6MvZREJHPAtx3RwBLLN5r0qi8A8nOThHo0TcUOlkG8GhAUoCFFUyXaryeS/OJaxM1T7XB6cWH
/N8IixkuIf624lHzIxCwRiNjLTktkgj3fVhmXsES1SSbxVWz5yv9tTUjOd3+dxchGrWWsJmeVHpx
1ppUsHFXp4kOWWaq5UIdXBdjNSXfsKYuLUPCf7/3t9UyTAN1olyHObBSRGNNu56+SCI/DPoUXXGu
Uy6xZPuROK79iFmlTg2/QPMB+XaaBMlv8Q1sC8y00Xo0sHUZbT/vuKhqJeS+789qpJboTGN7Xt7L
o+QiILEtr1DuaHmfuKjlRrnHngq+xK+Af9b/ZmgydN+IWSrrSd/YDHZK/wZMmHYwAniEz2kl4BZi
QObj4AMQ0fmYoEzDCACW4pl84H2AQ12mG04wnfo+ABe7Ik3l2SCSibWyHIIeuJMO4cfz1SrwxQJn
3mLQuTxcAuOYTQ+oyi/vD7vio3lm6fKEROV8EFOjNW1l4vVSZfDT623GfCw3Ytn5qDbgK0g+7TbU
QWkl/64ypydgBzZYBigjWhtfy4PhHqpsZshVyMiLp4D4RIPfFbFjtZZVzfMh3vaEaHcYrSw5Hu14
DyrdRcf3kLagIJhwwYBSMLeRUOBV1u9uAebalCE9Miy1YzCTdW36jfuh65WHlrJYBN5jxy1ptAq3
LJ2ScYfaVa4CqO8XiyMJSHup4pJsyCeyL4jesRf0l3TY4p8PhZ22B9/IcvSGZ1miHktw5kJBm1M9
oJRFEK++BfQthi9h3zD/WDZWYWMK2xBz3IKX5hwoDcyxrvK4Wprv3loCFzQ2b4UdInu4TSW8zR4N
VF9SAYVJ1OIMzc6QpxhqTlp+9EaF6TBCRTbULYj91Mlh6j0OX+ltR1z5PlEj//cvBoVNCvUDWhy/
wu1macvBJs/IYMXRTJ3mu7N8lMqQgE+f5cf0oSSPYITgfid+Ni81U09rIVb2eodvFPkR8UaQSUZd
DmOuNXvSBBp5Z1F/aR1lvp33e6GgHG2gFEhe3EMcRdVgmDiQnlf9SPUAlNAeLrH5JueyZp5eACec
5m3Y2hvv9t0Y+w6QNtAuwH+n/J2GA4peW6oPvZA3uTyuwbY7BUl5zRbNIxJJf7/2bnQYlPCBXHDY
Az7Viv2DdSQp4DAtJwzgffDPh/Pr2T0FS2QmTwE7plCMObgydI9ts2HXFHg/h0zMl0m4kDK4mdhx
4yQjSljZ9TK7NgjwrjmHv/iOCsY0iPQ2EICSwzLpUHQCsbRW9I4tl6roQO4xkZF/jC5NRxvmiD6U
t64jCvAsaxyUH7QyrC8v/M9IC0FERB/cjo4dg7cNo+BWR/xfnh6zeJUxtGUotBk+Q3l1vhYqUQQx
WgEXpgNK1BkIdl8COvuSXy+zouKkpqbzF0hpm8mI0r+fWP1USzPbJnjFLAH5PBzo0SJKpAlBdrPU
Eh6xzpX43muNd/movVccbnBzR0NFydlur/iKODXJALnKNsU/Pi1qGXy1MSxYkJOU6K1H8b9RL8UP
6YwyU2VieMBrt8TdXFFw66saJIlid5axOjkEDfhz8Owu72QCp0eReqzaPX1CKL9kWZUB54DuuPM0
2Py/a2X9oAN91ay+GImzlkXJuCg2bZBz3PVSLb5WlLK9sCobz+3JhJHfFp9pVIMAsjt3wU0ej0rO
dKm1GXnUhvRZ1mTExTg94NdJAuwjK38rWaF08KXq6FAqBNMU76HZn5CXaL+jR4H/Fy1otqBAAKfD
6SLDhyDvqEe2/yrskX5H4OxdN9VhWnwH1C6tGWsvD3j0oqmvt27wC7b6v+/KPUxxYIRl9Wc1wdjT
cc22dvA2cQ2pmwsrwhFlnipetsE0rqffkI5c1yNdcW7+0OHmx8eltbWyXTYwBMnJ2hm94l0y2NEh
l4dVHf7hHjg/FmLkFLHMuTQZJZTFFZIU/24URUMwE8DEdRfQb68m5aStenlZABk2HinnV6JdnJSf
DwaAdmnQ4zT5qxs0gpaLmAdYlUoqYI6Haa2GPf5zEBD99/O/pLqd0uHX3uqldGCtyZKr7tm1r12l
lJHdv0WVnuwc85FEiD9lWE2/u2aurkq2EgtyFtukKvW3bjlCmp5oSIwyGsi05tdFt9F/L8FOWQtr
Yr/ZWtwIM3vrPO6XbOyVuzQ5KEJALUppXrBZg2im/uEaOCKXd6zJM8WSVDQe92WM0xS/3dYOK3H3
UQuki9tQTbtCfbKfVOL/DV6E7dXS7c2/mTpRBpSEExDp9o5ay5q5Il1Hp7oDfus4B7Zz3VY7+Xy0
Ef95AIO5weZ9aShMJ48UZEYmJ57PJMnz6HiOiSQmrzADYZTfskczfdKU2kWAmZtCeyxc36hBycdH
RLtUH91M8AOvxmGIb9S/ShddFNpnJwTF0gpjtepm674oCSfWeE2Y75ZC5xiwyhiPW/maz8clQyTl
YiZthcuz1Iu8HYQ+93zdrSZ688aVS/MCgujkpRn4eQ36H5CgJrQYhyz60adZ00BnRKyhd/9O9TOS
ojVYdCT43CrF3lcdTih8vqdQHHFdrJLMFT47x5HIW++l9tNC1X/mcahlUs/VA7yy2HaQgDrMasJB
d5PPWK+fg8fbr24ps013xvDcUET4bvR/vdul8P53fleekK3YaSboPuaqX93gERJACHoFA4UUnQva
8x2Jq2qFnL1rq+t1YqsgHDSDnIRlavCPqdkiQ/rpY6n7QW4fCrTGujLc33iIGtsWY1CyaEwLtSxZ
U+4Fx/SVHsNX/2tnBBB/BgvkSUtibVamWwFbA5mjwA8FrV8lpXDQExzt0yxN1TQgEr2/lWevemNA
2ojnzmgyCHbHd2ayScfS6h3gVaPhZfl5E6Cj61e/Xfg+UAG7jt0KpZjcosDz0z8LytIhcgw2i/3T
T99jARbs1Qd8KcyCAZZx1l6K7kdfDSqN561mag51YR4FTEPddys5Qi1IEmzcL5RK3JXG6w/s++0v
ucw8xEH2gOMvSWK7oiq2/ojMjiBh69g/2MMQbGzDbDfw8fJyAdHWeT/mOWN6Bafj2UNuehXto5cZ
hjyuUXEM/2RLAkyWcohGUBCw0/5/LAFUfC8xAne98bYvoBb/HW2hEeUXwZpjgdLSF7JUN3NV/LGz
nKYREldw2AeCs2ZVm8od7rVtoh1sdsDQuCDYa7dfVTkcvf8nxxCUON7DmIyyYYLoEzTuodaGlaFo
jjrJVQbJkMnNStKHRoaZT367G8QhCo8FEP2Wl5F/c4/UGHruooondT1oerOGUOHdpCyfu4IWRYmb
J8AJ6xev/M+a/uPX7Ap26St0GsHmFBlHFuJhv4LusIZemfGD4qcq1NeS331jDQ8LUZg5WbMbYUSM
dADVnYws10UmEeQRdRkTC4WpUXkk4ct0UWLfz7WCnKKAFDNdszU1L7bQfDcCuimk/uSEJJS5jnKY
ljURNE9ovtBOTCz3SEKD/zcDcktmRGfKHz0BxtUw7EWwFYLddecQhHGNXmCK35lNe482Ldy3bRH9
4WPiNV/wboqJQ5njcIqbxt3AIR5kNuzpMxop4p0cRkdsww2A66PZaqvb5Z+8KxPEkqrfakAZWxdu
QSwJPKX3/hdo+U9DkiEbP4p7rLXLoGqaha9idmLtFdWfY+JF5uN5QYlcVZnAKmhedbLMdCcKlX3X
45J9nODSbmbrGfgrRhibpM8j1gUQRs3wOnxW0x+pExlZ5c0SsCqq8iX8BcrqogFfTNZ2igsEVc4d
2nYzFNzqHopwuJ1cFiMEfGRzc03RtkQxIA2OyDdMT9rftaOF++OeqATzfvL1GBXKUcc9bJG+MeL1
UeVgR1p3oOMPauUlwD1Hh1m45DZKhDAb/0/rdNLAl3EqBt8muBrQpV3HO+En5paYN9C9DVrGXhVn
tGHzO1dwmpqO+lTGhhEZaGqNRGYEj1L85Zs7iX1ExYD1D1hVZsT9kBPoiHKlmNXxxOKDTtEGwPks
b0YZ2+SIpsoVN/C91jjOzlZbLfizcYZRiYYLuA8vM4H65TPbWV+v7J9O+NRNH607s+6HebkHf/4n
P1UpuuEufu1+TGQaK/xuAt1tv5oRBEThKZJcTG2+8O7/3mLiqYicF+JJNjX0hE3Kopy/MAIJ1/Jb
SVMZaDyLSII/myTr+XOfY5mx6xvWeSGSjjDJo3yom3d8liwD2UxLfCE6YfFDbpxeI1s8lbSxmVTN
Kvqn/LtyJ5Dz4M2H/ov4ugFEHJ2FXQnrAiziwcusj082Iref+6OTM5eVYK+laTJwlEFdTvle6S1k
W1K3ulBfjYcDpKypO4PNDERrJa+uthhOajjww2gnOERqoqDJFn/xlb+d6eBZeRQvdL7d0C7y2hOv
gk0p6oroRwpiJLuTh0epjIupqzxbbwZF7H9HZtaNxDGgiXSmpoAcJfN75vBxLriuJqN089cmU2C4
9toar7tYOlfBhDHhSdXoM7aG028JxhFkPvALsQTFBT+srFgbzlJG93/RPOxgeAWftNVGHMs5Gphd
UPKce4ooVTtl4UvntbCw8hiFhAwQUY0VhL+21xMz+iUCJlSyFYNwQSDpafwN1OPQJxp44LLR6evc
W80lIu8+1qgn7r2CKOg+WCJWYYQXeHPnaO1aW5wCOTUp/2z06RqEUrQi/jX16n8rVS2KW/E+AsW3
n8jFmGxpOKlWuvJsnocLsjW8RyfL3dk3CtHNWgreN3Kiq09/BZ51kiWaYyXnwlj+J7R+u1LqlnVS
fY6iVutH5u4D2uezlvo/Lp+ffssCgaW25CazgeMvnyv4YRNvRt5aza6n5eTpdeXnOUQJkVPt5YK/
T/PlpNitaaRykNoAht8dU8r15avN6/vUtHoE2IipYzKD4OIaCA0zgbi86aMJEQMk/fdLVs1m97mL
6O/a7S6UNkHb6yzsfcFsG/R4irpSmYeI+U/mcg7J9xg1vLyAcYZGFJ62xCgIRGUAggDjAMjKozBV
ZHpX8CNTzUr6tECno9GcVB+ZzVBnre9iBrtHrDWSyd5emaDY4K0JKlYytOukqP6LlUd5nr+3Yp4Z
oeVauQEUf6phw5iuqnvaviAL4jmeDBNFdDhbkmJlWivdE2NMsVGlwUI7S9FYSHqKKBgTHUX6D7ZA
0u4Pu/pvwspmWGBDtGNXI4/0Wz1YyKIBJ1U2Qizp23hesDhVRHaszdtn54BKyM7hf1j4q4arLMUl
n41MMGQZfBDFgMsrkbMfoZjKQqgE4uoNumQlFLzI9Ft80/4BKD2TpHpnHKVQRmEIout1+wBdd1/P
/sHCGVJBrt4v6sTi9AqD1+s2pPyHzkMSJ3FmQdHEfJnrjJrpvfqzkfqAjKP/jDBA7DWRuYvv2ooO
VR5gOz1PVtmElcL9Corc5RW1tNPUKHr142a9RcB32RVuZmNHcfAjwdp2OmqJtSyNlnhz3QWmrIHw
rVHFdvi2gqnVg0mWQ8AvfVeXhz/4O6HgpB4S2KBoWwzLaMK1dO+izDH9vLbWTz5G9tzSzf4v1rDr
jUMLi9znZhI5GXby1cEXOwGzE50XthWt5tKoTED34MTF7pqSmQKn5+Vmz7yXFi5/G2/cOivfytfc
5vZ44BDezlKZbqy19CdlLbKBuTxjIZTFoI8zZqhf9wMGD8u+XiZTRjtiGyAsHcRBb+He9AGdws0c
tmpJRxF6htBFz5ExCAb3LJ8Sd44TdYe20sC4C7P+QFyR8CLYj4dnelrR8lp0kTKUUO7G0Ee9gjA0
ezHher9q/GqFX1YUCbmfSkUBmmXJlLhSmpRSD7tKC3Z/N9WmiDfZE7q3ic8flrqVqjkmg0ar+uab
XwxDCxejKTuziA0HkYlGVxvQRIuAgnzaIrhguvK7E1ASfT9tUxBZVhHnHpMPWqiKz3bxGrKwWfmz
2Uv42fLiYCZe8/XXa4XrEB1+uO6mAIluMiXMCoFvO+ICQOVHeB1UOjxR38/lowb+l7wiqRbEpEg3
reM9GHdogGT8yrPL8P26/uzlxpuUnbRWefvLkOHn7arBUQ6zSPfU/+TD+9EFfMcD2vTA2FstpyLP
8PfoEe/jQowE+VV9nBIPRVnNbNf/c1RVctjH3aaG+od4ry+/BgyVr42WwkFgJNtnLvNb86qVN29j
bcJj2NaypY5rTn6YO6thenIAtAIL2heH1Hzn4RXimx0b/aGMa9PfeAtglEfjbtystU/uw10MeuNd
bWDJyQGm9gXm+Zx5EsGoy5YehP4SKXmJVbuWvO9hShba0i8n2fZudST4trIeYR+YjrrD+FxGKDxH
hLLXs7sCe1b4EbcDUYvLZs6L/naaPrYg0ZO9qDJirh0J0ue1pXXJZhsDAiQc+Bl1pZp5nxHQIgUC
lWQbRRWL0jp2++5lPDuoAFBdU12vsTVBuyPRmvZXqc8IBPf/ovz1wheKz9rSzuaKbggZc2Ah1aeT
ggxM68gK0sQwAEmIXwr4fbQjEH9WT+dmnJ1C/Nrr4mwS/UqjlqwDrzDD13AotbkVpbTYF2o7B335
Zjv/gX7c89ZEF35SVH9lYXiibF8G5zd1exBhwKd+TvdU7ezKaKeGTnwUUMI7ZxtfC0cYJNk0GcGF
S42Yax6liWDhzjKgo4P6+yJhhgItrL9/Sb5FuDNvQ1kkskGkJJqdfBdPLJ+vTrOApCoiJ28i46+X
Vndl3t7hM5V+t5UTSxYpt6vZSIeQtjN6/RFbB5cAddv61O2spofAgCWOAjhmvRaxEj84FX2iyAg4
9WgKgpZnR0vDFodePh4tvakZsYPC+afj63lcYcd9fQTBncJ3HKR6qIsRnvmPgIsD3aJvTzt7rUmO
5SOOpDzzUO97uK6X90N8FWppLKzKXKdm5P+8MjTNvIPHoszgye2LyxKZ7nLqCfU/Lq7veNNC9ARZ
71PoIRNiBxC8ypRkDQ+3BfvK5I8XKGwDk6isct79NYy2DXt3ZdqD/VdLd4FIngxbfUoUu/DHw4O3
lOp6dZrVswVorgm6fIxeeRfBudDizanr81dfCzDMDturIL9PCCBtfLBWTinarhifgJxZ6L5vhtfl
VeU9a2/Ckus+I0AoYyew1f5mdvBNwFtYx4FFYbNeSmv35BVLQ6fM2/PRfW97VWfpx52rqd0A2Pab
tSJ6/sNlOQH5JkU/2kpy0pRBYvS9IKmqqFBLhHWfTEVmqXYkvN4cyrOu2eibVbXLyjdQwHBNwkry
YNI4VCNwVGHGKv3rUHDkl3bIGeGz7ECUdkoIJrKieXfRCCd1GNyvzKxi4gSrcuELIFLoImFRj0j2
NUPusCq+iuH4ahf1C/+iVq/1kgjzkx2XapuuRsE7MrCnVJftH5Nks8wlyXZje7haSaqyO7up1Nuw
B0hiqRG8nhfjgD2GkDuNFLR4FvSlXm0SnNzT98nxA6wt/gSkF70veDuJzkEYwyi+ctT2RcWaWJRx
qqEBt1QM6Fs6PYCIIoXA/hsJcgCYuDr0XaL/VyLUH89RGs4wmELlm9ThiHKvMNHcejk0HQy96cbJ
lSvYM0n6K/etQ4d4liq3uqEnob3Q9oEYnCk0fwMkvSF58XUloW3VqJV2rCfRm14W3oGWRTIj4QCV
4AEw2Xg/hGUxX7X68ZmbpB4pvNagXjjwsJotF3Vs7U9RfTeMlcgthLMoIhSpMeQYf0bDd6Gu53Rg
8UU7E26A8Z5XNzVCQQJNYgoy8HVkFaSBsg5bfHksoTp6oTXAuBVdey67/5WwkWcVYWcG4avJ7IXN
sGjPiYxLrwxxDc5s3Mfz8Qay4+uWBSmst1Gw3pztjmVPLgkicT33Simcx+k1BwfM0I35avj0puvk
ovw1FqYWlg9nGCCQMnc4/BpQL/ViMMtY6eKiD4SipFxpQnoLa022UaodedQpomRn5qYab5uBPqBP
RHMpzRjiFzIkX4S3unx2t05scjx4/pT0KHv4jIvXOExSxiPa3HwAiNCe6ONQRfezr1UvFHbhIRtj
yKCgF+Eq5AK9tPjxfcRpXH9NSA8HJevzvhKS96msd9uGRDlyKwVrJQigZtSy0ya0pE3SXvl+eHV7
HjAAGRxTExz5L7b9P1zAnduDkpRwb1wR/EEpTl2pPO4wvWqpiTVG0RxaV1YRkLhNxRpTyE9zO/A8
DP4Q4jQEcmj4vgsrtfbv6oKHXSwAlRt/73r5R/o+6I9NOIw6vRoG9bEPGbpgumZUd1NHYFPh1N7x
ame2Axiax2InXq7bxWBzmtMN0U7IisJxkwdH9eOz3IjwN3wZpYsO//v8+DsWaRh7O5y0XJN9ODrr
we81kcQolXpYKI0N8ERrpOzfwDbZhSW5R50w+4TAelyG4SCnGYBdxNo22NG2CvgDU878QVG8PRHV
X0PN8JphCx6eOlDec/7pvlb5YhjM+CufI98HsjDMIn2koMfRulh68B6oB7cEvcmUO4+QVGLCzJxj
DxWq48iQmgQmwOSngZ5pt3l7oKtSimQc+Z1jXxvdzO21dO+gt7NTU6AlDu8pvBuj74rOj7b0UWlJ
jBP2/58uXxM1X+waZhce8AVSmjO6ZCCwcN9bGI/tmO7gdukWl1wZoO/t3WLwFwaL74xJ8JdXTYHC
n3sTLtCIMcoiOwWXjLM0AS0EOrfGdljbhoIqto+LtUOwq5btUKjk2ZMmyWoUwQQdzvV81suuUeKD
TWfC00Sk9O5xGrfdAwIqve9oo+5wsr3oHyy4rnz0Mw3OiMfi1RQWb8HGmS5CjSDYYbnipLuBVN3G
QRtuT1/miXA9JoKU/cRSz1UEqJtAGQLE7NN4wyFeP88665/amAbtfUuzTPM0jV6R76y19ZBzigW8
xkrK3AYNKrZuPPLhvsLin39yXYIXIpPfdhBiJ9/AP+bu0n2GPh3ioZ908QE1NRr+fHGNIDUmFdpu
C0kWiGwaG6A0VSBrrYITSpxgECdDSfpXtuyCZ/SIwvaXUSAdruGcxBUZmUW8ZettHhHGfZv4YKHC
qSsYdCOpmHXcMWOsWXEefmI0jmVnZoHolY9E4a7uh1Wmn/K3ZiWX24Yje8LEbcD8JeoVmccSvucu
bo1o7dOip9/BzZXm+FpEJWc0zPuYWxKGeGUDFUGQ4B1Z7wqed6N5sPZu+vZBEvd20lmfORGf767T
c3JWugkawGsAT8wLXbVGEIF69N4SGN+S0TqusANNGVAEz4kWQgywY2TU/2nyg5zBOcWVxLP/gblG
PrZfYjuztISRAJORaJR71GBEGZPlH0GdO2BfFMYUPz3coKcXng9bglJEojyS88hkSdh+oQRGgZl/
5L5PBUXnz94i8BvdXpl5vr+qTSYgLDb8reJwg4zkQutFec7J6l9aB/iNdcV51RqibC7tZ9O/bm3e
fz6viBTf1QFbP9TGWNhqEfEr5kKwGZKWN73IneekGMWqw6WTQ7XQivY/c8cl93FPL3QM5zxAwKgL
1os4sSYXE7bdti3BeNKGcKmaQ/KNin7L5xG2ELYKYi3T8y9FkhZiFP5PRqck1aIBKEhkm3LIzkLr
1Yvl/8CjvXAXLpUpz6tKGgGLYKxbP1WRXU1xJFfQefv+n/dFZZaztPSvlqTWE6VD8Uuw+YLgURQY
ANJxLFQb8YKE9Zz/kWgFVr4fRFMmqDdEkeiZv6aWKh4K5co0NZOtbG0zypazclT/xWbqX2N+PG6f
9swclLq8zKBCPykPJO4uonFKtNOyoLeA8g9VfwyGps+gseGFQZr3DwfDltmw7lMdtQWVtYD/VSqm
u8oet1m9O06GNferJ91Hu62vCEUslAym31RmgLODsfN13WbqMOQ1OJPwQk5ClbS4zTueGOSzbAEY
WTcY3BUgbBKaGPEqyjKhvAe/bzA/4KtMM0r2Y4SiF7V/PFxs5mQwI/HsPMFx8fLGa9EGjxHp5RPY
zuSY4HxeXfIypUm/mQsjFmh9DqKei+k3MMwQ1J2PA2Mh0Plh5ediEDusTEcu02Cr1ZXRqL5XTsOj
LoQPc6dOglcCBTwPTQrMf1MHoLJhanuunZymKAfEwrGPrXOcNnDRoNxnjxIEiU5Z9nYhSLC34grs
/x9lVrNoLATQ3oiw2gCstHnJObr6VR9OUGJEsWNxWdxDzibLct+GS0N4QecwoiioxKpLd3ZT+i+y
zhCKFsluP+4XNbl72/igPPGTjZIKzLXFT1uQ3WEFr9veHTjJlge04tjqu0heiQm6Fq3C4MPtG5TW
q3a9MfCaEWgybA23HhKs0ENeWgxE3Y9QtZbWyz0gEiy2sf501Fy3NQDeBFqYZpTu+YKxGqUZXGVE
pi6A3VoUvfYgoLoR2l6gyHL4psOmi3PpokC6vGDq6Uldrw6A/n1derqTRuPXtgGmCA4sMVN0IhVz
N8bNE55TSgxek5mOmOMozJsyY9xWrfFGB+jf4H0DYGK/NpmhMjiz4AoydjTvj7gmRjgBAi5p6MKP
W9AJLTjJeopLvl/LgiSnZtR7ZfwJYs8iMByEFJn0QmrcEINKDe99aHWSJO3yG7xUJ3os1YEet6b8
fzhK6ur9PVxfKM1EvS34ZXlUcrZ7ZGmP9yjOsU2P2atWkaSIp8ufG/JYl2zG+hudfEVy5DXk4PRZ
TuefJeKP/NNaYGn9bCZ9eh7z5EXk8joZtkbsuL0Lwi1R31/GIgs8NCEnfXpGEv+1hjDFNXIefIeb
GKdwjMv9XbQ2IcZQFL3MIP6X9KCKNcvc2IAUiAuENQjFT7xoDilrgRoVGF60tKHPO3n6At0MruU9
mE7uwOxjUYbcXxPubMBou/2HQ+RTHB6UEGcNH26dF72L9hUhOQ+pzm+GRUKzAMtFLr+mC992y61N
BobCJOTtmBWKjo0n/DSR8+PYGYRW4qX/RjM9pAKrZrh2N8G42uK98uy2s0kjkTVwlPPJ/GJNhQ+O
I36U2/RuCpPz4htkICCGlkXEA7UyXpJ3GaDHOhHik2rYeQEvsJX49pW/pVyMBJsOeyIRIgjwx/DF
Rc6ALdyyDglUXe1LeNSU7nlouh29SUwYPKDG9jD9LO1cRukRKYjpuvDqflFDTfaVOhb+sZz5d21C
oI60BF1/0Hlhg0ELVF0E6SoflqSoRYjpaQjhbD0uRwG7BlFG+1Zc56Rw481TS9Q6ej5bemMkl49e
kPjIDWKpeC7jSppHwvLOLxgfqhMlpKmvk3rCFJiPS+ApCiSw/mh0Cmplyj55l5b1ppImfp89v4O5
l+0lWAAMUBhjdLuMiFvQEgco+M/vPqsEEVwz4xBuke7fGUvFOO8E27XB72zXzSiQlGJA0SH8xvI5
gC41lNa29tr3RV+lSms0/+EN2vmXeLEu7/IcXsHGT/ty6QC94qZZv00FMdw7inbgokd7wOc/pXDP
Ij2Fx+wEfsquPQHbpTla1F5MvdAaXutwwxGAAEjch2JEtoFKkl+ZoBL2vnBxz+MnY8YH3V4l3O7u
ntrGk0UaHT1GYgNLjLR1FzitWWFfomFCNq4VXx97j7AqeoTJklOeYqMpq3zUBedlKzEFTXOZ33+V
qChJWJbjUDh4QAK19KjJxNACx+u4oQrEAt22yRjut4amo38E3KpHwQ4zFYOJpR0AucCrr+hYk2VT
JlMf16n/Qw/wkkr9XKZrb+BEILyq7cYOv05xiADPexTd100ShacWSqlmdWYmjabgoHMHcLtuJNci
kV69jFHZDM+pGigSotHz8qDGLAanYRS2MHkpMi/ZjYErOIwxaohQmEUHKcQBLFjIwIymSthsOfJc
Az0N/334/zNdFR6jDocHZ07hHHA0aiqoYeLFEB+fVzCifnKbN7V3TzWfykRtfixK7WQj5K5EON/W
4fDCeK1sTDojW6m+OMOejB1n2VRU1VbOs/p+R6MsLCpxPV4uoNkWbBl0UsyQ6EmhgZJh2Uko3yHD
MglrPnAAzFn6swRiS7s0m9uLexZy6p5ksAJcdXCBhGtqHGXbY3l2sRf37cZYtC9/y2Earo6xS9v8
eW81wkG7CPkluwrDSO6c4MWBB3yxSPy6V/cM4b/cV4s0UYBtAxeNysOm+0gEIhOWJtjs6LS2GZo9
QYQZxDkR+xr5eJPCBYv4WF9fBUUoWzVKah/31ioK63rJkZ9lS3s0GywForrhL+uyMpgQsB/eIiDa
oTdsGRl/WlyAnNFgBpjW9x42NilLEoAvqPb007eBhAI77BBZgFTdXL+DnFt9u0u/2my/BI6F9APv
OOot9CVkNwsjFV7YDqywL/Qs8mHf9eH+1gvurvnd46E+6LiYt7UbAD1QOwFaTB8E2j2PZp4PbIcO
7cajpO62neK+TYCCWOare9VvYGkG3DXiMOE/YitReN/1zoJ/bAsB9xiaF+liBcSwhbVACMsXGem0
U06hK92AlbGLeYS+234aslkjM9MScFwE5ajsvPZbd5vRmlK3AETm/j/enKkM1IwXhZpeQpEyvoUf
miA8B8WieQ9GSBxTwMDvSTJZOVOU6mqRwZfnIDFDF+s8RVlOdG18DZPkSlId/Y7F5Tc7QADep9zQ
oGl/FPCNAOfUS2vhW6W4Bbp6rRf1WvhiE//YrIpmmZ15srWqs9ItkXp7H9ijK8Q+ZZ1D9jRgvLid
L+74cM7u0QkRZfFQgtt4Q6eY+DosYaI0QAwIpRUUWJVcQAiqY/cfvkjqb9n+Ckq4agwbodp9t6ir
4Rm32TWlPzLNHJwESHvGJf7MQr1bkY8rHC2wHFtZTYkfOgWN09GkoGKlHg5SkB1q2SxxuutQleMC
e+nMmZmWCfs1kjl3cbAWBXN9LQGTQ182hnUHKHow5NKA0uivivwvWVUgvzmQZT7RAxUiI5khpu3F
avb9fAr1YvDmA5qC2G4ZBq0Tzo95a5C/1VtCdUq+ppws5eAAWKgpiCyQm/u6berHzNACJD93s+UV
095Lea0xMV+5ohPfPhdsEg/wbvGh/U1wuId6Vi82MQV8K2W6k015CNYdq/6yeyJ/jxBedelSRKDw
Etv1/i8UUblIsZJyGdnFL6jemqbwcnRxLcPgJeOgusdJ8lO1TQr/ng7Shtdm2YRXd1dlj6/95so/
+hZ2BuUX/Ya36pArU8M3OXMZPtONi2OcRgEFVjOERkCFrr+WknefUru8p/bPzzDNNEK9dD+1NlMg
SUI5KTtaNWmVlwo8VQZYmKLHwji+61e8KHuPyfONqJLEu+jw/ALEOQ/DgZwm3HxVRefduatxD8lv
wPjMqpKpwl30hhozDqh2kqVbPOpkFlnT563DfrwBh99wRKI90lw8g7TMVBQhgVDnXomEj3zaj/AP
xfO4zpiPuVIQNHvBNd/y2q91KTYKGq7H+l5MzWHA56FWefHusawcwb1+k29rW+tPkGkclRSDDDBb
OFffahXK4LLoGC4Pu7MfwgXKm1xBnXLen8Xw39HA+kk1TPJvpkQRosJTiwhLzuF8pANZ5fR9eYV3
Pivs6vvE475Bgfm+UyfmDjIn0Og7mj0qu0Vd4161rIqAWyVStADxbLZpv1sHEUdGSx5NPl63jZcj
4AXgAHUluHh7FXamFz5tbB4IMoFEDcfOnKU1OKz0a/a8g0kWmNuXx3CCA7628DvR1FZeIyZoolKN
K2jls/39uxo9chh5490VBA9UAazLiZGjUhiWVFb2whBZ8w4FDGcuPIebKv0UZEPuULEJN9qFUlGx
pZ6tMGP3b3bWFVnqyODXm6cHhafgkguee2HoEFGqYlYJH10ws979cJld/gOs+VnrxU0jMEyQQ8Y8
J3zpXXByha3KpwWvXIMa6LaS9V4RNW5ZPpNghcKkU+IBpDKI+6Zdq/CGLZ8bqvKZ+bNth2hjSoxX
McLOWspGicV4gmKc5SRLs9gwTrx9Z35uH8a52C+k0fAfhgN1D0Lyc3pw88G0uuYsfb0sA1fbR4TZ
VAelFZ2EYIkQFYhNQqrO38E9lnZyyc7jjomHrQT/GYGLJn8sgFL7k8iAQ+96iYvBykYGlsf3tSmI
oiGvnoW8+RxBxwHS6JZjULpB99A+ibldA5354Fguk/lpnme9NET76O9o9ikZB2lWj2Z+iMaJrk/j
3Y8wkv8+jqauHNdWSLuqRkUPZ0eCD6MuXLY+DuHTA9SQZTg+OGnBvPdtxv2T6Vnd2x/l/7TPi7r+
xoyOfOBjQX7PMzcbMaqF0Qt0a9gHWIbEXkLTwZH4RdT3uWWncurDWnH1jEWq39cvMcYMj9lKxsrc
cHxFb3NH/jGdwPi5ANUHjx0dkhK82Igx9zwhccjlvSn1C+VX6un117bR1GZQJVA7oPUUno+OuqnL
LSUpF9gZF0ssV25YUnWrJeAhe/z/o17Cz/Gdi4UfDgQnda0ttis9bKOWV1rdZV2cD31eWpJoewZu
jCysNaCERDfSxBLkdZYT6/9dsOye4leo0SRco8jsSsH4ng1uZ63yG/gRUssR5+WAyN/MrQhsaUzF
XRDB7VfbyKrmIFfVHvhFS2rmVP+3bifsCui7UpA1TkKYOS46LqfQGEv78ODS3Mr8MTZqztRZnjPx
AEUr1bILkfMooZKDjf+cPRL4CI5nYs6KphPgopEqA7dYagqhMr/IZ3RUL3430wIiJOJrrhtjjmiL
omXG5Hp+mvm/zh2XSZD8TjI5BmayOp+iQbrw4oBDuHDWmiVitTDKuDBADfB1RKC1Q10l66vRgQpL
DKSC214s0qWlHxZYA+VpMxf7oeBW4hUgdPiyuL/gOFv0jjXe5ETxhPYbC/VWeyz7GoIlDgssI0zI
Bci5l2rpGycjhO8NuxZaZ6rnxNSL32PCjKENpeV4ftMi2yAOy5DhmKl1wKmZGH6Vy74SNB8CV3TP
tiIHwb6eAgvTyTfNFnIzHnNfC0Zj8MwmIFKn9sNpJyMiDvgBTSGNUDa0gjs3oB4VhWDKHQFGdiiR
rY07anKu99ociZTs7pZoPHfmw8hFbyiff8VEyWCLHqBrJYcY8pmJj09FNsTo67BXC+sx9oUSc1xn
tac2pvZOIRJ1HN1/B/yZm3ykSKHtrjSXpcWpMDNWOjS6Ys99rszgO28X1lFaPOZzimjfHV2Z1sxg
Ffdi2R4CEIeImIGhKrECZuf+iZ/hYBKNP3WIshGvyovgj7W2r0fZv4H6366WsoUEf6DmWxCC870O
WMDTgj850GO7x8ujKvswuRR+33OJbNmxHPxXH3umGZYxkD7EW/1kSJfaiH8vWNk3gO3/VG51De5K
6wL6TkuVLXpEutX0RwcF/LJOAQsUigAFIRkFv7bC9vWW7enS8ArC3J/mPgW1aiDW21ZOUXmFWIHT
KSQxhC1j2ZzaJhga2DD6gHEt12yGXZT0zxQQK07JDxpXGatL/1mU/Lt0a3WayD1GTJFb81fJzpDY
2joJ3snHrfPH8P5p1pD/qR2IXoH50s8OJxRJErBmBcM2P9lo5MM8Cm1KeGwiyjH9bIckc0AaqLnn
VuHuG9ygGC/0qCKao8j8ybD0y9uzJUL89uUvXMMy9aLGjRGHT9uZS0R8onXDCRBCiAzaNaFym9CR
SAyj1lSKEmSTa4BxQuVYFLe7mcX9Lo0m7pSzp5C+yETo+K6WbDMQP6O+wcDmOtzXAW/54UzGtplV
LUK5HnOepjRNJlhjsWo9ipviieY05sI1h/TV7Iw/3ANhOm4+7/Rt1F9CdgJB67seHegejMs2h+jU
BWh1pfSzw6gfx+bgJF5P+pr6IvEoe9SVackswM4twUoQK647c7B5xoSX+TIEOq0SmfgpGEzc6nDd
tPhYinKMaXK3hH4fK/jSDcDAjQagQhIppceJpB6rMHAKkmYx5NMRMMf5uYP6csANMR8fzSEggW9g
jYKlYVPZiumziD0ioztZSS4nZiBg7Y/ZWv6ysoJp531c5Agxl2cM4abgLbHKv5xkiwuyVcTdVx2y
QrkJkYNUJd0Cnimbj6rWqBGgV4zgcMNyxequ7IW5irA3ZL6DfSnfE+gLpOEq75fSUl7gPQ9OJQ4d
KG4EyGM+y56W/hdnzXQBQPUBKWeI9EaYv1fuN4I7yoQbMwYLDfB2TaWjszFNLmYCl51CIRAAHzox
gvmcKXEQqm4gJu+5xLDBquDEaxmb3Nq4thQNcVPEVBVQs4vfRxgz4TFz3LHwIk0/231LW/Kzu9Yc
cOOjBG/RktPSYMzebPgTIhji9lT8BSBI+znvmBVAjZo+8xjLyR6kXqbTDVpsih1XwdNP3qxqLAug
abQwJWIxirPIpch4JIGP9uB21eXmSOawm3j70yHwH6w3TQr09dDpvLpZi7WaYLlCIUcDbZx2NcDo
svYg1PdLETQDE092/GN+3ERUXkOn45DP6uWu4IBElUuuqB0M4EuGzRtZIAZCmf8BF6ygSnjzU4vX
t4IE7id4FfGghGREin6vqcVCPBci4RCJWmhgJ/kWc4EFRrCUPxnX+wJuVKrYv9oYp9EIDTbQzMh6
Kd4k4DMCrF/SiF5+ifzuS1EpDym+3uMJqotdkzfg1qEF+TlSQPCQgJI1ha4ZTH32+vXlt4Vyenxy
LX/Ayy2vA8196BMbbWP40pAN9bEvYzxEGhBoCE70C06gvhCHhsc4JbAvpur3qgG6q4WsZZ0KQoRr
TxVp76wPBaHbqoUNEgFE6MlcKt920Q+BBvTDcslVrktWTRo81U8pOl+a+r4UsjMutvaq6STKOhGt
/yaOAYwND3u0V8XEsb7gmmjat6u60vtzKrbzNQGAKpFy9vu9Rh+cIHfO7VBw/MAxx4d3d/245UtT
/u8sBawPNf7X6uhEmLxIPg4968nI45AgcyOsjTWBGLlqHqfu+H5+DreM/Kqy9d9Z4LMl99qRy1Ra
wHjNL3Ea0xtgzIfTOWp6Noead0b+LJb6+GeWtYjJhxlOQvle2D7UZMRSNOFh7D4g/GkEsRov8itI
zRcMZn/oa7wwTlY4UJ1cCGbY1kZfhyUL5tcUDeRmpveWgdY4XzO9cCnxcks/TafHwmp5EreoPzQx
JyFbEbZ7pSuwzKdHEyYBbTSNm3yALtGUThU7vEGC6iBfpLfqSA4iTZDz/14vpkcQ9unW9nJatCq8
8TRbrepgqBkit8i0k8if0U3ZFDSpqQZCQC7K39vNTEJeqBIqZmVb15Q2Nlis4b6kGMnVcY4wyimP
GLMtRw5bRsJSBf1Jv579JnMkiFZE4FI5U/ZLhfm+6UjbAwjfluuN52z9vQQDITArFZJ51/zRhISj
YNxU4Cny+1OhG38Yn9w9liCWJ2eCPKE2z4khxs5g65rk9nURaQJ1QUkziEPEo8hkLMj18NSixv49
kRqph0xbJbpodkD6wochONcP447AfLWTBVHq4uuyZW+KA9xLJd1Umnsp/ip8reKolVWjHrXjz+Mp
g7aLiiyzQkn+lOITY+/dDpTO7m9FKRBKVodJBVwv+MNw16foMC3j37vcZs70EvxqejbV5MCnRWiJ
JxOmZ0RA5YIRHK5g4EQ39Uz0wZGtF4aP23hWB+VUjC+cSyJDzhwdJ7wTjgytdeI4Amn+uj8skcZc
tr6Pv++e8iX2K8xh75/1RRPoQXRDQ2Xc+LO0pVBbRrn6utyrQEqHuadrZ0kq4TElH3PN4AsMJ8ot
dr4N7/rp6Lth2BFiRron1Dzgg/sKs7AeAhnPu/kHoyOc6zm492jGmRaMT3YhqGcqCVUEyZcMfqsY
7K/PWm631FUbWOM7H6k8aeuJyL+YbBLtk5it5+LTYJiJ/2lFWwx7jMrUSCzqcGmyHBjy0SyxqeJI
jPditA5RNoLZwr0Ot3qMGEXpe4iqfvQmEmCnoAi8RsfNrEkt6YrLnouBM1ksJi+fSI7QltWHZe9C
BTnPCjlONq3vXiuriUiKoEEAwdTIQaAxjPsG8bPYiiLoDaWnWeU+T/DZEuFqKPmzslhCUSq4VQ/R
laoy5TOXTXTJohGUCs4C6crHbEPQBL7dU3CJDWbyQaQDjNNpKZsF1GjZ3FvoQFsZ5CO9Nwze5XHe
32Uzvg9LWZ9AHr5ZGf+HPJTorbMp/4ZY3j9qIzI/6DBpPMzIVkxgL7gmvnDqbYkJYN3V96T+lvZf
hqcO03md0R7wuMiemYOSs0+s1YdsM1DorlU+PUiMRynE3c11r36XKm4egKhrh4MDoNTunAfAQI71
p0leF/XFJoqGANVudSEoBlFMTLJiNIaQEZYmljiW+SYpwci/3vd/DJVku9ATd2ZyLHtuPwAt9n4P
7Aom20+9CQ14QUEci5kXyVoiGgK+QfcHJ4PsJhB/klKB38Yx1KNH92V5V9drgcNmZlALvxe+3Hou
ZBOcp7OiyVG20uH7QsEHRDXWfB+ZKScg3yOZ35ZsFXj6Y8dWxVivrEwcMZHWAravs21qyYGG76/U
aJ7+0mcWsQVi8mYxVbaploAsMHIgICQrZ30w9FB/MfVmSIkzCnk+wiqYn+PcqT4ldTpeALtdnYqY
U9DTsGis+vhFITukFCgz3g2XG+qEni7HrFgY5uwSCAijZMcZhbS91AFYMpIoC7PCoHr01gDbjXLE
oxo130pQXxoC29SGaqql2wI4SdomZftQyYesaYySrV0cyzNDkEQ8ebPB35LzS/Fsi9WB2afM4xZ7
oRc+BT8ROK+20bJtHMRZ/T1Z6y2EYCcf7R2NpRc6iy1With17Z0tVGML85zf9RFTAAb7d1YfIHu9
253p0XdtvzWZcY4pBvti8eSXxV2ullyLCT31vDBGIgNZDeLBFEpffVCYgbF14miY/Y+juUA1BKSa
FPILRKTzuNONmAujjoOMmyJebFto6943scUs1hDkm6JFyTDwAlyRWB3JmSOl5aP22GEidDVO4IgL
rRwuG84MEki2icU3CVvqXKESqbi51MWcnv95GrrEgIbOmzFc94Yip4qz6ePkCREtohev8z5CkNyg
mJ51Sik2MD9Np+R0eHdaUQayjqGjdNDkSnxztFKLUbn/AqhlUPa5tzncSpkc/ivUAbH2o+ikTPg/
5NcVJNOSk0E60OLJgB4U8jqn9pjPTL0cmEzNOkwfnSdyU7/2tNeg3sV+kGajJUBL4gU1P3aNU022
CuQAdgDDNsPdmVr5Sw+n487eiYhKOTxUfINu7bWgLmv7QC6tZ4bIeU1BCUA42RJsC9nrCaByxyFs
JqlYMe4OcaY19mrGL8Mgg1ocmuZ+A2A7wv/q793WE5IaXTeE3VoJDW01TEA4nEF6JZ9ecxWNZKt0
2ql+AR9oHPejSWz8idLwV9auAHQF8j4efvVM7zhSrOcZ8H78it+Vof24FHCobE/EVy6xxsCkXicA
yopsKY0jdZv44SPqRJWng2xUwR7k95ZipzFkxlESdlwDiBzYO1jIrGu5zPtk7clDWQGMuz1gmIia
06yP999t+8+9alAhx+NpeQAhHdeMaeWkuWwdGFfaL7LtJ7XaW6i5TxbSr4+OO5acKMY4ydAGRuqf
90yXEpcupPhPa+yvrzoMxYHTnub9GpmwAHOKYd0nL9j4bLJCmWxd7a76smmsyNWn/Ilww4PynYuw
hXc1/12+vND2fxpK+LdZtsNs7vJrL8a1VV2a/U7QHM/JZfuO3u1FfM20oZt7VDJQPhXH7lgnA/Vs
tj6tyNeOZKBRNcK9Yzhv3ttR+Gofun3ePEAIRP3sGPD37l2fprPLA8NaU6KKsllU9GgLQ4KIXOeJ
bVWZzuIQRw6nxAK8ebe8szGOTN1JO+nlPocnQx5CxuvrZbJ1KPxkWqrJ4Agl04xU3+Eax7g1Dwmz
CKPyV7LXghZyaqckybsLxIO1LeNieDa/lhp9YGRJalXTFI+7G0sGMXbGaS52uELFjtmJkVnvaKBy
ae89HRzhLdxp0qQna2ZgBydYKAgSV2pE3kAOeAG3TU8OVMNTsKYuO4VMIhk2/hHEs9dXGQhwZLuS
yi1UThHYnvsGC9J9cCDFQIQeEjWE8bIlh6MW7AoSynHifL/rEqL0xuO69ygiawni7S69dJvCW/eL
2Lk+b/E6+8GoL7Duzne87s3uej8RIP0DEUyXf6TzHJyhUwhAFEoeoy1qSO0jIJBMbTsND4v4AceN
3EnQ7m8sCQgVC6QEJUOKmgtIZygdx8Alxg3eCDk2yfHztxYzbsidQYJya9yWw1NgU93SRO0dOMOc
UCOGlaUuQJJc9Gic2LBsDCGZl4AQdTEEFrANg0NWCw13LY3g/MH9GR7uY9X1NImFlWyW2zIGBy3+
/7IMrTOjZ9WlhSA31bcC+phWUBbY1CXyESK62eExRULgJ233g+j+NN2zuveCApCsJSxrzNA+Xr8m
B8KI29N2VvGG7T/O5TjbEHbAM+jjgCKZ5r93/gafQJ4GhCyVCyzM8wQCuRE296zX4v2bXM1GWJhd
F9vtEVthIneYvKnLuha/zLyctBjgBza7m3sPmxu9jlIZjOGK6r6CxW16y9NJo0qByKTTszUB/I6L
6V834zIcQsgkRltrpnvA/MnR+kMRYlbV6dNctLO5fK9kM/hCrnjqvOdWjgWxZYdPbtPQTnv1EunW
jvgFWPzChq69DnkgBlL9Qog0NDTD6WykT+tHa3vhvnrBcn36tSuA5WdJz6wwcHYx5KNNytRcYQpJ
YwLMevg0HqZ7jLX0LMnpQsy0SsS836hxNd4z30lFnVWeco0iia0olRf+GmB4MsZGG3jUGsegzdyw
Y4qfR6GyL6Z5C/TP9+uStp4Dj6XOlLWXZFfjnT14MOKhZ6qnEwGeLfFeo4Kmx7jgsuXVnW1syd4H
14shBfhYUCk+WksDXdAkN0BYCm6+CidOzokpi29fk6J7ouaLo52kPRVs9CVc0dgodd4W/j5WZ3qP
fffiHD+p9KosNQO+VtnWc1sEnqlBcKnke8LE3jz5Yd8MnAr53nzvaVrd3dvKwKVQHxCtiNFxk3qm
CnyXUbgZrByq/UsXb+Q8+5VQId+/2J+vGSYdWV9ryafj84kMqTK5FzXUBVSyh/RLLWrHAjpfh0jy
bHAxdDn1tIJR+n1CQ+hsZyO4K+OosrdUmWTVMyidPPLK9vUGsiYA72wUE91/epDROR3rAk80mzO1
n8d6OTNG3mSdWIczvgganvZsDsnnE2t5LbN/vaugZ7kJcnJgK0jdRLJprTZNnBRbbT9a1aUv73yK
FfsLqYADpvkJYNBUEIhbs9WRmqCmJBwMe01+X/xuRAMZpE2TPk7a6ugylMquWswVeMvvT4m0c7J8
ZgqAms2SjN1NX4Ek0S/0pA0MQfV2yPHxB4QVJXxChh3awWKtBWsJ0EfpQLQr1u0J+aMqlrDqGevn
9G27rKIQ805ZG7V5oFQrqJe2RZwLfxElc8/UXVrl95r5KLN7kwshrwOLQbXlkyZCNX4kXCAnYmOz
OMF8gVJc4z81UmTqNgyC0dR//BVE4YQXg58DNwyRiPv4toVjV3Hvspf4zwd4sP46AqV2Y/3yqwMz
xBx/BIZNj8g11B7YSfgmkZauZPNcWOiuZF+QA+Djqwr00rRKaYjMEpXbqXgLmQdx4lMf0XQfkjqU
6RimxkDGR94fIa6g6/sXHsmZk7MDIO4oABuosTKjx3eSaI3ZPzd28DItzTcXSxJ0Hx+tf2z9nVXy
lhOlROlcFLw0tjSCb2wvIGIQ4c9WtX8ehb9iwB/NtqIjDMDtuVj737IBeH55Yt6acGfWqnkTBLPV
wzJia+rrDSyZGOYBbmPp6qg62lbkrGos6AYyLgHborv7T7FvpYRhO4rwwAc1/oduogatxDAJZaFW
i80B0KePLpOhPXTUQfl/tZEfz4056RtjqwxWwEe5jokrU4nQIJzoMvfxEXCTd2ukuOvSyrZh4MnG
4+p0kReciBTsFNRvYmPYEvoVkuo7mA6rYNt/jhT89X5U/yD9ELFZAjBctZuAIp8nrczOF6gsNzzS
UYivbvt5+Bu+Vy2pmZhyhEHmQzwzm3/vslrCXo0MP22M+Q3Yvcy2HPcL0nJV2h/KWGP9R4XYFPM0
HZzmmQLyRpUQPuQFO8yUbNpYFIdLOvtBjvXIfFGyOo+veQsR62ALNQdMCXOEXn1R9F0O/BBgfumB
GgKezK8zGuQ2VIPkzWQTooT54GUbMdWeVv0qjlI10P/8jVvZwdWY122D6D0or5qyGp8//CPK9gyz
wzMpzy1W9nqq0vAV/mRWjfeneApOxXu6rzKdb6al/4j8ExTTHs7Bv2kfBxRipyhLVsiJHprNmfJ2
YpOzHXydg3a0Rv7ed1mMDVrhDTW08eXwptduaUno7kgJ8f+4QSB5+c2V6u/aSg4aMR2K4yI8tuZ/
7IlI/SNg4fisl3lkZyaVk2n4pkmYKSpIOrihW073ACYNpJ1MkugGe+eFuedLYJe8DedHFL2wkvd2
Qj7axOgNGd267hSt9nbbmQhQY1P1xyf/30+4LK12P657Q8heAgjzjGXqAScrQYXMD4t2QUNgIxY7
tQd//2ZQOelXfhSOp2OFQuLVsJOhkNdzel2TvEYCZDZYV4CziNoLRTam1+wyjtP+xRuCQnsL3PCa
jnTB5LIwvouADL69T7DmSmdotuiBAsSp7W4Ew4h6pob6fG0B73dcG0MjutbnwvcffVaeSX+zNd5A
7b9i6XL/WJoSnMiUulkUFGbGKtRHdwcSDmPAhjphPu20scTb7toNQBtwFiAd06war9JPkJmXO/4j
iE1gB8OAtyHbqRxQ3AAnUAkHSvoxeqaakWvw0TuQEYaLIBarPXJIOqJiLmLpwIHtSl2bpEDtD2pV
L0Y348obOjk1CcEjTZ6MatZlDW41Ya3UpHfKX8cQUsy1UJpZfUwnejN7xy4LyRB1V+CqA+Dibdao
gSVz0/UdOATQiXkm0AURDJ3MDwSJ+ewUOkt52rwx9hdQmrx5bCBq66WzjZMIhyboHUQuDEjBYt/E
eJcF2Zo6W6XA5F10xspCMJN7cr1yd6HY+XoLFCp2rEWMvaNX4/D7Z1D1pgoL1KIPVhhc83NxD8lQ
mIr56mieYj5S+mY+x08omYx5g3I9Y1p1+ivZf2PxVcvfF8R9ZIsKqERWxLF799MZ0lrAZiVPYy+n
zzyn3k88mHM7+SzPWJ1b4hUiHAbx5+Oy0rV+xlhGXP4z0MgigHvmDEPHNIhqNPTqoBbOFUwF3ZFc
aIrKWAfMBJTRvogk79H7yxyFC6rFVBOk0Fe0ctOmBTcbjO+j9h7DQA5BVsmfGaKhj4fnABJVxWfE
SsjLYdGi22Yv0A7DjVVb3CdrKc8HhRGQbg5A9vCEs7BAL7LeiL4JKly4GAGzoftSiH8NMZXoMoXK
pg5cBhJb5e3VG89OwzfbNP00p/YUNTz4fiAoSUT68frFmShiNDl/krmyr4dQVHphnh+MOoElonjx
zhQRJb+UIBZQhZloRi3m40anX+a2lKVDGSfcB8yCyQwtRpZzpbPHPVJbCegjXj6ACXO5yM71LhKd
aV1dwKOMuiciNEDOJ25v9G8ku8Zc20kufck1Elkgmfy5w7IF9Rb5unLZMXP5aFYEwfi446WayyB7
a7Huq6XJ8E01SquaB/LxI8H1ZPV5HURO6g3BoitEkiaZSTi1B6tzBAsMrfB+d4N5ki6OtKTyGXz2
ae6FspJF2NFpVIZlnktefHcHSKV/q1rFyuCgkV2ngDlUBMq59oFjRAX3bX0LHeYrw64dOdUsG852
ODDQisX/p0gsJL63LmAKqYg8w6C0E0ah2t3xkfzzGtfndEtDL7csAVFrRcpYCgU5sicFCAtt5T0B
sFaBUreBjwHkRI8DNI2ptDxu07Oy6ct5vV+cmLRD+H/ygtqX733wPFGQkUtn1Jf9BWUc7jnd1edl
G+oShOWAKFH9XP++/WZ3pzJYfk1Y9ZM88dsiHJm0RIPSKReW6t6NFGXMyKPqW1hMaE4/JdPIG+tV
RaR3Vz5TzejjLWc8QCV/M5htZfwdUoJ1JNV3Ocg0GV604yiroDZJ1chC2+kmdlknaFl8Fg/Pzf5q
FaTMVlQVX1DNu5k8KDHLTUwfQII6l5RqcYlTU1wsSKHCc5LTUlQ9aYQyinaUUg/3fubl5dM3idev
HiMtEFuNzPdsT0LrjUPVPJQMxvP4i5W4NWSiw5FctfHGQ2gVi/OjNNfy0womjlVRcLjKa7g+8Gks
8BDr26C/+27uObQ6peC5A1IqZRCFjxQ3Zs9FupJ0sWMEl4vD4iJiPT/mDkTjJnzfkBCg2gfrn8lk
gyAstGAr0lVyjTSy8rlVHIfBGlHCIg6O63B6zivp8GjKCrr/57bsec7sqE92fNgKwr0gD/soRhX9
P9FNfRFDPFyztl9iZZA+I1LpJH0pQR1QJFj/UhSObs+8gJmYfvsEf/hcIemQEhji/Ghh2LKMZZQF
ysbCK0Yjpb2rI0IL9AJ5uH5VYKjmizQsH9LizkyV1zzk7JKAEf4o3w5DHZqCNLohbU10fwKoRyAV
feVc4ELTf0pfsN9AS9pThxOZaW+LSqa+u5vhSWEmK7g4XFVblwVW/tE+uRPMOYp0+cvi+VjAV5M6
yC7E/F6WBNPZPyZ0u8fpx0XLhPFdBHQV6W3DZmOvvJTLRzaeGLsqxJ5LS+hdSjvr9Q4YxdNvSe79
AjtHy3IZ35glXMvxFdZwes8FYug3A9GZI57inesatbiB7pIARWoe2YC+diy2qfObOOKObASTfRfv
NP8nuzYI3gTaJJlQwt3I2FnoKYmF+hjU1sNM6W1WR9rEX5JWuvsAZLWfdHB4v3G/8sjBj/laFxDB
0UiWY4eiKFC+RlzjMY4ff+u5bqOr2sF2r/WTjNzY01TpuVtjED3WlKTCHVokmg8uPxr2aXfZksEo
o/jJz72OWYWIMaKS8t89X0dG9LOpOAgHHx8NDrOfpEtPO/KAFrILDQ5CTjtKAmn9A6QTx/HW31BX
pq4dpXlRO3QkfUibXW9SM+MZnmiaPdmlax0UKWqu1mqjhD+Bity7PA6tWElGVYY0WWRHyUTfA4HF
4prdjFWNsskZdycwbwZvbGX2EgTJoGNgOAkrR2SAKlLttZYZGkN8yN6gmx70LvqWiTbyPjUkeBYM
BH/0b2VZ+alW8qHna06oZo3xcDR9If7Wtm7qTLCdPmxtD4CWCmxxO7Vtuk/C6ZlZQm13HJLYPBA7
oBfQXI/A6r+VYtm9t4ggK4ybGlFEvpGWspkty9W0SZjtpLHHND/Ibmjn7x6IKGqjS01Dq26kOzbn
Tg5T3654gBjWmJbOXjha63qtLsQ5wlRgtn2fCheVd/vKQKTLlHCpRzYnDiBjA+JA8nqowq1vgF3z
ZgSUmmNO2yp7ztlp0+GQaTG+vSSyVMj4OqDRvYIvAsk9lUkIINgCL8agTtEBLQyC/w9OTyxAZi+m
qnH9BFAS9Gb2WSRqgkDKhzy8DTXYNDXpWZTBvweUqNUioFxBbhdlYPjDFtN0MlaWV/73xAsD6utQ
9l5Vng8tkSlrfk1dMkd0s8CwKi6OzEhJ09fX7Y8xmFiwXh0IJPKWL15XcNtY8PSirRE3iiwewhei
dF66a+hGRy+jdZ4dBmiIxbsiL1Z2OEqfnblfj+SdMXYLpYHOlTndzX9iNENl1u2xiyh4ib0CG/ES
jTPixiPpVUtsRQLbYbi9OIhcqTFPPiISTBkb5z8rkP6AlcmVwkaqplZWNBEP7teruXWms+b0icFc
z4QRCUmpZHy1JfSAHYc18uTwgf3fwResf4odrXrolQ1Pqy1ZDGQ9ciYWEnDVvFxmA0YHJ0SwvLRi
BSC4nw3KGj0rYALgeJn2b5SSdVYpske+byg4iQ2eE57om4VQP5DCbxjhVspt1IcAHdFrKsYndi3/
GqlL3QLYYPrkFCkQNBQf3I8VdI0cBnJ+GaLYZJw09HzV/kWgrUq6f+LgYA0bIHuK9qAHM57Mdj0S
ZRbuppoRDBQ3sHZ6wxESt0XkJK9aM7ritHZZBG5rz/kQK+LQUd1Gdngh7H2XlAzGY40nG0HIxHul
63fwkDIAvSEyB5A/0Y2afbk+CbwJwbeb07vVVPcojYAb8yGt5aPaJe8mMD8ujqYtMatEzvO9cUqc
C3TxdnPuT9JsVO8GJzQlvJ2lTj59LPLq4t8Py9W40PLOeawgE1wwt17SvM9Ua7/tYd4RJbyPUzLY
YvUoI4mGAvbs1re+dhqXIPjvMl8bLDmbAcuWn5pFeeJ5GeEIcZ4JKThLd5SfYkRlCIGGddj+KnUr
KmNevTxU1PmIx6BkfupnBZBrKnsTZYxN6kdUMtxejsqqZ6/UMbCLVCopzXRIahmNNYWQ2n8tN/EB
QMM032IWU/ByfBcJ4oYTzlCb4yecWy51KeNTIIfkIBL/my91BkeL3FnotKXMuwDa++De9UBW1O4M
fllY0WL7ZwLYr9a1tChERM1ksBpeOIsumrGzg2wjSszExdIsJYuRzjgMyCysHk/x/v9ZiaY17KeP
tUhnml+xeWdm0Z171O+bnPJfMQiANafUj3cpQTniuG/TFkSCGHSG2LiJ4xXtL04nLcbp9sAHibui
e98aB7AyJYPKbsRtRuJwdSe3X7YAPe9npLGv3ScRZAottwCe3ZtDz6oDNAT2qOy7yLxWhPmHZaTt
ieG0DA4OKl+ExnoAf5WZySuX4r5jjUpnTbqLNRzBtu8QPGHGq+uR60DL8Q/nxYsCBm2KG5XyOu7Y
j6SOra1ynomwCnzTdDaMawi5tpFeV48ckxbPOJWRWJqPKL5dhRS0ctMDpmRgzCnsMrhCcj+QnSPY
rM7GijBcGDdDJ4aCCfbniWA697hIZSO/FPQjfyFA4w7xikmPjoQe36ZoORbrGp5bqLpdrV8X+//E
TGZ1NRSgndXbFJ0wBXGFa87kOtuKa1e5xtV6T7viAeuEr6aEuLbsj1AC2S6kqQRrgleMxWCat6Yf
LzQvBzV/E9dfK4aIvIZD5CxmSk1dxWDcPyupDYCcfhyObOiTcomZxdFVgDsk6AAXtq1+zBzVzxpO
pWGjQF0KWP7JsQ92jWgomNEpm3hUGcU0H4LN43K6YbBuNBSLw2RrkgO4eWtqkhMoJSbXnfecz18D
/2wlQB6ioC0GMvYCZgQyBHb7u/cIecPy69eu4kX1/zw0FGrfVVD+sXOo4TvUo8k6ORJmC9oNW97Y
ApZippWitI9Uqbn28Mp7uMDxf142QI3qfRvI4nMnMJCL4WDespGilR76qT5ZgAT4UrIArtHprPWA
3FKMLX7/K1wTGzAaHml3Pwy/6ZxpOX3MXbcKFcPv48X8trTrsGfoXY9BZ1WyJcc8WkUwb3Aw3Wid
P7dEt2LpYgSMEBzHjfB+49v9Ty99R/IXarhVtSXEmbTUHvp+eDt6VqZbfVtHX+GOgKZmMq5VTjGA
RcxXMez4WtlYsEWR5TgRvgLfXBgYfe3tet84Weua039d5KXmIb6QIk2vFXJPRnQ0wMYQuLo6HSwB
Auxy2BRYthizknKE3CzaV7ExhHvauLIyqGV1+IdsjrwEaWXUoJAb+xLM7d41A1znyfPYNoFKvyFZ
E/40buKXZ/Yfp/LbgJwidKpAETn/WttWQgUfLphtx2V32e1qqTU2Dk4X8AccftE9wTA8PAYFyo+s
rvYGSmnF10K6mdaDj+NCMbCi9PMwrOokgbK74H9uiNLkNVQ8LcL97gfRj/MTfHa2MLBQEsBnVhbx
HkvHjjgkvnyzpbtKzENgum71wvnfFUNTuxI5wekeK831UclGzSkErOJwionGBdzehu2VSBTftEwN
m4LelWLYvLgNWmGIoBp1/EHuOpROg/6i+H39pgVAxAzKRt4PdZl+b0NdLuxL5DDLLXrhlnQ0uKBi
HBlaznhm+E0FIu7rDxYxPLs9iuUHf9vBNiIGj3AjkpZoZz+LDTb1O5TknnRlh2BUu/ymozL8Mgnd
JplPHW1I4ZhzSRGDrXeEUT21xECuch3dlpae5T04FRg+5Jo2ND7p6AvztUfPHtVg0nkN5n/T57YQ
SG3fMPkpyOQO2y6zpaTFMQhaINJO58uj+FnkcodLqerigsA01F+k1MOAUbzrU+fJsQxtbha2pjS5
EwVBUvTVI2zXsER1nzrElAgRAxW1FiVoSAwHcYqY5zl2e5G5ttHRoSyRnzDhOJI7kRnhY0rMMEMw
9+SVqMQOydDHYpBpzxd1gnfYKjsnFhKjl/9UX6uHTPE9FBh1FXhQCsPmH2p05hxh1STdJG00g3Dt
frp/x26vfOaCpk0QF6iqA5QycsyfQfIqhodDI6hOia5u2ica1H8S6mVC69yqLip0pMUYSMu5wQAw
N61XVBxYsa9F1PZzBOEmxJhQHriwWLTfK28+6Nv71tQr38/YzwhHcENbXDuSdw8j0c76XtkS9UCc
kg53/B4dR7VNZthTqhK40jXH4AqXAO1MNZpCelTUpqIvXsaYGqvWUXdLOYL3v2xaCGu43NevYU8i
yElP+RxDqy3CZeUyq7iRKbdiuNTMA1GaFDxYIHRDq/hI7AkYxXAjhdThylMvSMzBY7cigitGANuK
o1164hpTFkfMuuk3Gu70Udmqp7Kn0nfWmNArlembxeFjkvbXzK5aeHlCmMFLO6zRbndd5yvQkyJ+
gd5+FarkE+jtiSys1lg813BkbYKsFwaWd5u4BHMoxFVXh0mwxvQr0FXbbFowl7FHqjxeGTHju/dg
RBBebMhrK36wIKxeObTgCxBTuwvs+wERDA5TZSr3GcLN0GGd0FngvDAMP7wKDnqNNFc9wTShg6Cd
5MWTklzdICKs1bA4KYnWr8G10AOfYxp1Gcvemi93R81GQ1+147MzmVOf+Xz/7mdqENBrNinU2H2o
haSX7FYxKyHMfOY+z639rIRv8eDBtSdqZ4QVQ3vHXWChNc/4BSNZme4DO3rBK5oL20p1z/F3n5mi
K3pgWk0LopLFj5RkhFvAE73Uco4esFpsJsQytviGhla0NEm0KfxHgzrod8F5e/HyfX3WIfOnDqR0
+GvKCHpKxV9eQaj7H99/8veOugt9UVJE3O9K4Qfq0APaCRqngRtVDTI6XF9nznPoRpPwro5XqdUK
9pf9QSo7ksiCnFms1sgsFwxcXgCQMNPAJDGBr5OFIp+eCMGws/BxzFfpZ0CeoclfmX6vLj54JtO7
dgDo2YzJGw99/zPszTRwoIjMW39lTcF7DXo60+ujCgjjSYkrK0aOT3fbRrprZIdAaIAcFSFj5v7s
PQahItFCPL906u1VOXHOfhVcT0aVbLI20tgbv28d9dRP6vIFMEJJXplF7hWmzAzViR//Aqn5jeic
PmlODXes/pRmo7VjVna6hc6T9TkrE9vxPftnxnSO+sAwUd2CiAjrw1Wjk6fIdweSDKKguOvKr17u
VPPtkcvDoDC/Xhh5e6aBplLuiKVamTFf4rpo7GfZehmQ1qqDGqIICRUfhyMqPM5dZHihFUfBrPbe
mLrcTd8FYqwXEmv8s6NV7Z4AUEjgQIJNZ0Fkw9BVSKUQCOKkLiqqdyjEKPR/pfwYi4e6YPh9bFzC
JgCEfoJgEc1bjrRR/yqhE8PMU3sqy74KbvEq/P8j+Ftd977xwUVt64IRqnd1OAkRk9LaqdxOVdBs
9FPWaYymrOx9h5PRGR6ej24/ZjRrnEeGWw4oRwvHp3umK5giEUFgcdlRWEley7Q9pyR1EB0pGk9z
K+BNel97PcqTtQFDKNbT9V77Y+CZIQka6p9BJ78NRLNaCEKEBAx3zLDxKSiIZieuJ59Zn8FxTFLk
rAvEybvNOtnrBmfxeqIgWcqAidKmUI1EOBVN4q5fuSHbJ0y3bWuniT7At6rssQy2GLCxLMJBcv64
UXsjuDi1V+CTeDvE2jnW5henDEbsE5dl9vn6NjxVVQTMoLV7BH78uh3q/LcxarXf668isQdm2IVq
A9wZTjts0OZDrVzJPLkbMhutX9t36DjzDREqTO6HCEHdTbV+XT3fPp34IY2vgufuMaQdKeVH+vW8
/QzQqvkYl1F1HvC7vHsTlnLXKwpOoyserZMHJPIPHZ8VupIymNp/2R/u6oRIM3qhGZnHVZ5o2PZp
aMLKlWE3bTVlKlXTcygRsThsdSr2XPLlU927hHA3KklI6r/iPhfWtH3+wHLa/wHlLM3/O1v9Hvgd
9IaMQnWh6S++V+mAnueP2YirenDOoKnXyUEl4z8AL+1/XSEm6O2xGaDrHKmwywl3tpPoCookVjlT
B3RkTj0E2eBZTYx1YHIIU7PN0PHUl4QDTjE+n6/28RzNPwYcvXg3E0vlVRmWx9oWPzDz77DRvUtW
hOD0yUkKSn3uhXKCjIhfcClfGqG75iVW5g3wIVGywR0rysmcKIPQhrvtMjr0Tzfq6vmxVGrqOnNQ
9o8PJEyB3tuaBMYqhTNJTwfjyVuu9BfpbdVTY567dWJgFnN3bAWo0jLvNNdJ5o6ABgQl1STebEZH
5bfaqAwVuZxobCvHJltRpVWFeLyATEPeShsNG9rSJkrG/omyo0+zYYk1Fnskws/1eicV9MZciLaR
j07pzxDaK27mZX+YBbjyVLTa89mCqDDNeQJQJl7U2CRdq2UN0sCSWBSSrVEBWOUw6WxG1qpVJBCS
8UC/TX8a7dpRobf3QIqCIVAY23m2EtKO7kYTjKrmni0AhAgpd4v2142AU26bIzZg2bL3O73YkwaJ
xrvXJSmMfNjI64jmWwq5wnPQWelf1x4Q6m/4fOmpzVwXn0Fx3z7tjGDcm4VVH/KB9aXUrxGz27iY
Y+/FAVMXOk38/X337uskPxNCMoOvdtVjpeUI1Mp890k9LLtQML2mfpphcCRX9uBLpIXwzaegwFUY
QkpF6tmfgZ8tGsDQ+sl0Qy0l+TJiGZl+994vIYy6ZZo8/gef40pKrwxBOLfFAv1TCta8lhA2CevW
cfZhyZB6Z1RPHavbIZ6g+WAt+bye1oqz63v3CLgOgN5N5/Ix8dBQWvOqFbyiMjdjl/Pajcp16lK5
XgBfulAIbZFS7a5/W7wfnfmrtEy0Lnkyk6rFnBLsoPRHyBFJDvDDxV5xyJD9/CxjT//3dRSa6dNs
jBiGdmgttreOPV8ynUGV3xWV+6yqtjnWItSNPbbtrix/hVv/qA24yqRsVZRWanBJT5rs4Ebc6Sk6
zzBDqRDY2oXO2nbRXDKZ5m8G2VtJWoppmFBvQ0NFxadO1vMHg4NUUMDL6ZauMvqhH+bCp9ik2dQv
9klTgzEsczySstQRhzcjLptISLeti4Kkbw5XwClXUQ8r4kPXJk2GsKsoAnR8pAiEV5Zreo9qKJY1
50YgSpFTHCXXrehy9GuN5nmcT1ZCzE9y7nKCBXv322fJZHo0XlA/At8jLmnWLVCvRjaThzcgIp6S
3n8w0Zc8LGv4YyBRY6xbFVIygtVo7eQ+9BR3BveSWB7gOlfWH2L+wGD9wWoEChmGU2yp/DzLP4Y3
bOeRNkKXNAW5Tuxqpp2BCEJwQmIg4C6l5lLAMTtk3tIv41CEtNiZxTuxk+R7THzhDn5d8CczDT4f
j0sONPskrStXLLX1IDF3rMtcilk4Q+Wo0e0lglQosDPs5EAD+FUBM2S4tHo7ahFJVdCJQoTXO/aU
mD4D1Ed0LGtBbYTRPM6dG2oU94ZdCGnT0Re23OzeUGqC4x1ZmLsCo22o8N+2jxL7q/WA+2pZ7vI5
OqhqqeraTDu277ROaNPnFj16OZJZc+5Ub4ni9AGOc4SstuN8LBlLXFOD+5EoSkhfoaKkBVzVk1lH
bOQHTzV7SbiZT4JwpJ/haQ3LcRVTbpj0B8V9r4gNn0NjRyEoty0Dqa+YkNZ0OA1hUt0aaqHnHtaV
goIJ8SQrtkYT3pcyO6foZjbI8d47/EXKAEUcZtU5Esy5vMlWoXHhMKM/qDkZfXSi2gYx3WPA54ZH
p1Ymb5mAlJYCHfvKSFhOkcfWNEiAV7G+EOrZPXlgxvsgBEMd5JFXg+OSlPjY2EKf3YaPo4DQo8vx
p21h6XIWJsS//ovIjBuUXdElM67VlvzqmWcujhixiLdJ2esml6g0TGvKAJUonK9tM+B2F/iSuptA
UYgnhFGhqMGLiW+xaMMEPERsQF/8+yjaVLQAbO2kMEKHzca1dO7BCenfxE5oUTqW6zQDwrQ7yRVq
ZUbkRglFzdGNVdK/whhDaKnMj6LXqXPnpnqKTyfxa4o8iWZlLs6geSBSIQhwGf68iMQmV2i3dJoy
NcjWoAn1upGX9Bqp+cKNQxpv0hSV6JFn1P34efH9sJBcnjz7Kc5y8LhTI1bVPG6U0k/bSOEDI0xV
mdYj/F7k6Es7DvE6Ex6P2QfxeBcKH0jVGv7Su3tHazRuT4xd9LbCWb2lB0icWzPBCuKUPPJ4LfhV
v9XJdtcCeXK8TvKiszYpDpWfeMLZ8F2zxPMnnVqvFRv16IWYb9cnG/gy9MrtcRj2GjJXyfDlwRB0
S4s6UVDRpC/RgtnFM/LNoxQ/+Jj2cCshykV+idshjbpNdPkFC3nSJcb8x8JeGic9h5rbBlyVQGhO
YsrfTPxAlpSovAAR6m/3D698gtWOEqX+FAtt1ksgUN5maDQo/1u2NtoL6AWlFSYLi3AtI4duf9Hb
6kdt0D1GgmcDYozjZqTA92cAuAuGFym1yHx09jX+MadTNzlytdBjyDAdW1s5oisk1qsW9xbEVBf5
UpjEA+vGZrZYskxe7Gb8IYEghTTw+DSaDPpi4ql8JWqTH9OoIxNxJmVZHcJHpjPvy0tRKzOsko5Z
u3QBtG+d7HE0++m0xd8O3rsoH3iB5gW7P2TMLKlN8N5rHuI7TWvHL0L4Yo/twucJyj6gMZPSoQIV
YNcW4bKQRhMDLE6NvHe/chVId911k4OxReJghvrBHsq5HGXVui4Z/Vi3ZCoK0FFix7YgJgZCR/A/
bOkSilY/90pzXwkBbkMDPQi639NSgKE6VvIE+hqIp3CIT+XJk/odYQw+/wOzXwGUR/Z8tJ8t+07z
feOLpxHp97/2Bv7KbvQ2d1BF7zx1zI93lmekl8qDYeqDZXvEIwuJF4yh6Vj18835TJjm96J2UVkY
xuK4dSPGIHW7JbRe/1e1TMtRIhKZS1F7Y3ifyN5PW9VSptMmAgIUtKA5kvUSMp2mDjrs71zLTkAW
+rnU4uiGA4bA8doL2Q+8KHmu0eyVD9Pjw9R6C/3Tv/h1a3zPwOwU2YavT9/XbGs6OWVAvQjeScNn
89hOzR+E1EOGptt4CjIreHE/ugmpb6M/F86Y55Pg/WpvkmvMx7+QQUQjziFQ6XufsuAxgmRdTAh3
4hGXyIetTCHV8e+g4Qh//KcZ7Pg9nHGRmw3ZbX2y+zWNeA7OaHGf5ABFOJI7bxBceGhcc1TDuK25
NgsLfau1CcbFgTl279ZmfIDTQqNYggWcxCVWjSplUvih4G6+x+vRCZO9zVHGCoEjJymXA6YkjhBs
AwtfnHa8jCmPhIf/Ync91K0bK8QMMJoObvbe2sLIeHIAiBj6jxAMv4Yfgyv2r5mbvMdA/EwCqqqj
N0IidIxxEi1oqg9hHZG1gklmJit4s+j+SUUEizkY1jkLehQxWDaZFVdZNYTuI6MtYilARaIKmXl8
M2JuIP2DIDdag5MIFTgR/wTq2nt4APNdDHePCo4vakw48br4PeODZJ03UNxI6y+W5fZ8yFmbmuXw
eccb/WUPnx2Ic04SwSIinSOv04rnPadmSUGxxN6xDlA5hbVHvlPniOugBPjEoF8HUZuouhdEcnZG
sKZIlSRc6vuZA1vYFMObXV+CopdIbppnRkXooTGEwown4ayQDjJKSjkXsEkvdRI/pqrkN9Ch6HoX
sp09IXW3M2a/ZE2gVmxyKvLClGgP/A3PAQsh1kLJJiWdj+EgBUu2R5tsN9juLVu6CVw9XL45LC1O
B5JMHxo1zzKzilO//Nqai0QvpluG+IUIh82KmOxjn7FNXS9hVbv9umhQIp1RSNCJkSAP66nlusFW
bPsiOIxmWyLM2skO6PxSAcz9exAStW/pCRR+hsI9mCaa6fBGzGgSwlUUE8rWs6uHPYIUW1VwrlZO
aOJc7d//StELdSItLy5372u7ln2YKZ/65tr2tYo9Lx+FfbJd4bnug0jkOFD9+/tSnuOXSFDFObqJ
EOD5jBhW3Xf1kZp0wsqwk42w9nYMJgbZbxlBWcbZ7AG8G9Q12Y5bSnnhhtjlEWO85eu+C4whmO3/
RBlyCOkNROuprvI8SNCmnaslxB0uUf9cDztj5xQiri/4Uh31IwnKastE0824buh4GfxSn3bebNDc
Zyv5AMZEf4BM6gplG7qn06MoADr8No9fOqlRIQu8PTx2RoUc/tZgJZtWLZlJUgYpO2dlE+ELm4B/
m+VHbVm1P8NnmPBuuTcXizPsMRpaZZ5jV7C/ns5rP7TjS3cZwyPm8qL86wVq9FrvaW51p/l6ijTM
qZz/RNCzocLWAnvyIGAzuGjXKEW3VXxvXHFzyWoQ6fqP2e2tsA1lP66JNTiO9LyHPr8xVJh8beX/
yCk6RMNmYkvvv39e3r7/esZZhQYDKVPH7WM3bLEp/m7wJU4EDCQ1kQBQ7ZeezlN86ASDCFmTbRZr
9z2EGFOU9AKbTeEIu5i2rkWF5yP3s7nVa0JsECvYz1CFxVYrd1Xcq2nqftPYV/CrbqXBe4+g1lSP
N7f+ePS8010Pfnxf/ZD0LvqTlRqi35fDA1fdb/NJxOon4DAp8lJ9mbd6v9y4Snjga+uCLR1igrYc
STiEIKxtuLMPa+4cei3Y6VSQ38ka2aXSw9OJhOCeg8lEi2CGloN2xT53/zB7KSXmdISOWk63nbHq
GHYnQ0D1EKmIHE6CsM/BkPcVuhbz/A0BfKVCRAgp+0pNiNetlEPPctt3TXbHf84g7MZiRlY8CmJr
/Lb0dfgy6AVIZVW9n8f8VjqVhKhqE29IR5hyNL8zner7supEhWRUCLCQ7lVgFTcw6Lr/AsAHy7uK
LIAhp/ppefLI4aVaqJ8hOIps7DYM1XeEyR55QLj5dtVK3KqaxFF7jLrhXGHOJ7tG0nvxMnNTF1P3
qtUq2vKigvE6UmfO8MUdF+dbf9hW1abZWrgt8pIZ7PqWowR/50hciVaQ9/Gc+QCUQoVto5QOQYh5
r3h9M0Lxp97iCz1nf1I2YmjMTBGctwNtHzADSk1qmGnv2ef5RtdzeAsTDRLjDbDq43WpNakDpTtn
vQrZ+9neAH5xVhdPNAb4NJSJnRezvPSkdbtB1BUzuiPDprWNxHT2XOgsqhfK3WWGIMAMWXoDceH8
hjqLxPCM4lB9hvyhyLfD3WFrnan1bcVr8HOx7SFs1WBFA5zu0i5Xw9Mh72Y/VV/E5n+1mg7P444w
f3bxM5gBV0sCBvY7euhU5BuwQnKU2Z7uWGQPREA3qfUgqrYDav6W6cZIgWNX5MxMk8qyiy3iB0a6
FQ1xq2fvOGUKM4XOqL6NR3xb5dT6aVTdDhOUAn7iCL2T4FJZfzfCeBfT6SYguQXaET4UVUO4M16Q
8m2DZtS/eVpbETVITsTFeAB5pjoFHFzIUBviI9qnmh0tixFkFwN2nk4kTcFq0ixCopIrnFoKUaDY
qvcDbWk4EIeP4e7zxJ2qelY0VufbmrR8XrHyhV1HBIrkNdL18ljaScxtoSRQKZkRm8HZJ+3M/nwD
/v6uH1sUTRzPYOI9Xequ88JdShswPQt9dSsy/hYMHA1SGd/JEPB6oOwwvHDq5xs0MowduLzJqykl
XCiHpGk8rZAAAvlZ3P+PEZKu8P+X1rFBxichTxP5MMsWOb/a7ZZ5pnU41Tac6auCIcZ9IRRuzlOg
2y49BEU3tbb4uvi8sEJmYUrzfO62TGejfK3eSWESM/GfImo+3QKL1ZiCxyIX5+JaL2i0rgSszNYW
aR42hMJfw14t9k/AWU5ZHVbb7ZIxcJv2Gscw9ES5dCX/JsOlnt1RtFo/n1t1w4tBeIZwkF8czFjl
abKKXzRBZMRcsnNUwGUBaTv9od+juqqxS7nJyFm2LoNU5ZuAGXSM7OjLDBgL+aG61vAPQh9j6Mf7
MQJtTNuZQw6/l+SmbVMKyydjHDxpfHxxtWCVwKZuhdL1kPuHJeo/ZKmx3JYy04R2nXUzLuB2jBeW
p1XNvVlMuhH7I6M6PvdzT81bySPSOnHlgHnZvE0zhvjRYESEAAqgK1dJ4Ror7RpTNQimaikEug31
076jiAGqwEu4TagwM9j8lAv8hvUKhtBRwGFGz5UYGxwmFJgEtDB9XQOOEB8OPYysFTV7PKwwU9Sc
yUko7yjY4vty46S+dKC+miOzp82nlTHkgIRcIW0T8QZtjbO9tKUPOT+qZ42aeDRBSDIAe1DOlqPn
bdhXoxalpVe/NWgHg4RSMkyisDAXx939OQ2qsRGZQA3/XAtLCY59WE6WbSt0A3ybmuvMELDgqdav
bYtDFBbxJJmGczwx5ffC6nvkCmCpC2syGeeo5Lm595Q5aoyc08TfK3iKVsW/wPMpzPo3a+Ckz65K
+slBaAv3N0rE+6tOI9zspATjcrGMxNsyTlndWKX4TY5/QixsEWypKehTKFzk8ESXCYz7odlmbg42
36xyUzT5nFAeq3UvjbupomOMVUrZikERKkQqSbMShFx5cTdDNtUUZHO6x0xZKB4CBTcDD3Np1rMp
QjzoHl484mXBUXtqzbEI53caeytjb9qsElpLPsxlXMih/iO/TKIBAOEP1zlegQLCSiRkZvjo4PE/
aJudeVuu+pEmSwjLanowrjd4P4ebc3h0gL4/ifq/AQ9eOKKjan8pSzFXEvH3ZF2M936uY2eCOAv9
uba2SNq1GtaLK8NOQ1gicnAyP+HYroC82ZpXigveB4J6rCfwMk1PcBW9BNCITC7qWYx0qiLILlzi
oAcicPMsXuoWfCBpjrZaPNq6bQnrO+fXfFq3cYgqnPQVszsIcu4qhlyNgRkLoxGQxXNQ4UUME6dX
6Oo+7jL6JrI1EXrWzOOb7+c69rOf8cOLNeVyFdlW/iizqB86foB6x2bHcnN65fr0gOpawWAiTfbB
Ru+eChc+JK/B6kyI/jRCpCAIVp6dJkF7fhV1X6VP9pgqgF/vQs6i10WPc8zC+Z1IJVR1dF9cBjNy
GjReeVUx+DcQQAV+bqELm5How7C4CKU8s8fMiOuL48zEE+HHw7SFGltfXvHRx+1JQReFk9xc1uaQ
tivJc3z41a605knU9qOLwM1cWqzN+94ggTgdxdExbhPQRps1O4QBDAaGBrfZBtakfJMyLFGTAKEw
0gox4d5ysTGOuEXLobeLvCNEQ+i9oJx770RBtPQdM/9SffEF4UnqcBQY/A9cUXuig4A2cgGBUWBc
wTuhUibLqgaSknpcx393QTMnZ+YzlJjHiTLgF00awKs+PrvOHSTchOq5Ks0WhcIN6CfakR7frXo7
jBHTc92oi/InX82tSUySvzmIt39GjEC+dA7NqrcLquLqCe2wMKlQINEq80XffwYZmx81FuXyY1Ul
T3l+xvCTZvtbKPQxAdn8o+YCN8ukETiXHMJDZtU5uUVqITp+kh5iJkU8XcbwApy3B+cNNlR2XgXi
j6HgFbfN/vj4UWe5GBfSBBbN2R0Tuujsa6LKPr3zLfE75K+TnBLw+JniU2+CBUOC5aSpzUH642y/
0OonihSZ7t1b/HBAeZVqGblFLql/O/5+HIFTYO7VgZeAaHfgx6lb5fUTwSxKxlE7LOv1rGIzvUZF
/fyePOzUlDbuOF4X0aXQP3bjq1G7HJ2EYHduvLuPxfaWprat7i+dEcuEjefhLDTe32G39EViG8Nc
84zMPc0knyyzvhfw/e/OCuQDuPLZm5QzQ+RnK4G2O8zfAlP7farLhoHP3l3CBla/Bxxu0kjefsax
AP4hwtYWd6pNJDaiw2uVJOlI0xcLhrkt8m3xWTvbOuwKdOUnI9U9dvBoHeGob3GQ3lG3shiTxWp4
7K+XP6XQqrWgZuv9zNptrPW3PCMxAn3y7PZNCguFZzkKj3gET7apXvopTjmuOkelcSqDXlcHUYtF
69yu83pFNEEKH9WeWnHXv+DyglF+TQRS0luvn8P16PZ09eKA/qB31ef9SDIcWI3xZnh3rLhGLbdu
CjGPGye6nom0MjI2qPnGaiPmm/80dKxDtCefLW+EOX+VWjN0V4DAO4jpHn+Y7SoH7ju3czSmOLLF
uFXOs2VsegEta4ynDGmyr8kUCZ/lkhgixleou2mrLmDkvSBcXOuzBy2KB8XsaWbpzQbL2AthVmP/
q/9t8bNcJUX9lppuMXFEzFmHjGupWZ9CxhOFCvYODuRZL8UamRP0IJd4yCeG5fxEyx36t54Ozsp+
LjYixnUD6CL/NR8TU9yydRJWM0L6Gh6xsgGCudaPRjVR8KWFbNI+NxaX1PubftGJuhhqNSaHI9Ra
gFioUzka2r9TgxDP4/sbJolD7MxrTqQzlUeCjlYYIRMNKgFDNFvzOmWAeyoxj017esUGhiud/huk
x0wf7VWlwQkzleKBcorD8820SuNGoxKAI7MSpo/G4N2v+sZ0JKfYoA5THbYb3/aD0lBeD43dNprA
RLnMme0/NpLSvQJb0Ci7IICPPVz9WnxB/AyTE5I5PCW3fjA1HmaQxJpfLecydPs86hHj5sI61rpq
NVm4L3udMTTNQzrB9L5ZmFG/kg+tFNUPCar9TcO8Ob2mTrenSC6jjivbGR5Q65kO64s+AKa01OtN
kEzFTxLGqfCrf7dK1Gn19wGfdwuhDQuNyvpcT+GR4KZTTrQ7IyZDXJAirtp5nz239g96rSRd8v1g
vLVzm9P3porY4GBWMWQxAolOojjVnLp6spcoNZ2SmgU/FNQx4VXM71pQZyxoAj1qgQXFTdta5eYk
Nd48flSjyBR85KBPp/mJ7xE/uGY8Z8TZT3VWjuewGrq3XSOmoroqnP4WIugzbtTnAKQ7FIXTJ+Ap
Gr+tONeBoi6h1XNtW6g+SX44EUxGs/Ws//nINz8R9r65ZeL41ui+fTTKZc98ruOHhn1jy9x0evob
fCEItcGEjrvIj8jjVrRc8AWeiMKjueexl02bqZwjLQAmrWC2FWVbSwTl1ijqhU/gxb4OMTlmGQvZ
CmJAV8BBROIsaxy85DfLi7ipUphSYBbZm9IXXspgg/+k68Ax1X8e0rWukKf79DCwiJ0jhANyJist
TREM/M3D2djPy6QjWYe1Y7maA1Og+uzZb+1a6hY3ckomLL2s/SrCtEbvfAUn9ZWOipFSbAMemejz
B1r+6OzTMSbY2FwZb3mhSk9LgRDmPSKrbjkZ5O4VKIGfBQssSbXHkt9gzRwG37k/HgQe5spRKqp8
bQxN6m8YNObeTY/ZvC+mrOhlcI3ZNVyA2BUZJR/yvj6vxu+7d4hMuHxWogJpaov2D13mXkym8Fdh
fVCbGccjU6bgkMR08lFBRH4Jph0GqYXVwYtxAXzpJKIa5VtI9T+6vMgbZZ2M16oz48ms4o6QIiPV
4QuSk9aAji9OZcG2FNfnZ1TI1mGUXAlMxKYsENi2DPBHZ6SmNsL2GgQlPR9x48c6B0eH0ZIOI+vR
fFrKKfgtpJkLzQ3fhZPwgwbuoWTyRMwmWbBCp2yyxay4j7JSHmV6hRuhmkG9KzOQUU2Prng7rYjx
EXg7Prf2NpidV1EwcQSFCjMP4KyqmXrOebiAGdi7ueUMm+rSyYI/7HGAcA/aEBOigdVq9fy0Ltwd
1lpu/7jimOtkMRwFg/cst2hyjTak3KYszetIScTgTVMBPwJWOkZokXxMjXTv2Jk/b/bLDbbW2LwF
P2TKznot1Jd7jsGYUg6/c6mOnFmfc+tO+Pkpr412SDe++4cmsU6aVVu/7Ox2o6wHNk1yxjWBALpR
z95+TQhNZ+u1yuAjWDp6pZoL1ioipomAxaIZm70oEUy/63qw8a+Yp7Oliv9bC/NUfAFlIcKjRByM
lKlaqu+Bwnnb5NHF0MCX09+N8244kPGhARAkU44mb+K4plYKSGFmSAlXJiTDm2Ro2iTPrIeFg9z3
bJcn2IKHBwpNsduwelhbuNSAtPbko8zMuYW1/XdDONLPQW0Hja6lNqj9qAzd+yfa4DN84yTBDj9G
sEWo0EoNWZ0gNPrcriEU67pUdKQFvdeKEMmWQDHFNDVw9umF8QByFyIRUAGNCfO7X49R79M+ioUm
mPlv1KbSWb2GJGdoBNq4JWoKRbD1J38yy/G4c9+Dr5N0RoGRrNtOFUiSxtn2w2cTwsmCZy8MAkWv
TC+li14u0W+YGKbJ8T2p/lh3oeSgHsgNpLK2zDECsuhH0W23/t8CTZ6w85WWeUh3IQWyMEuFDjJ+
MGmUO7m7F43UJ2/tYi4lkCI8Nl8U8uA+fv5nJLAfQoFb8j3REqQCp96Ax2S7yYKtm9+Yqy45wypX
xuPpv7RPinwx86AOlJ1yXEMrgaTkyMf14mPD5amN9R5L9TlqySw7XkmflUgiKQAGPf6XMo9ZZe9k
WmTs+YTXf9OCvzX7vNN13zsxUh69okrhFhBjNkTV91heMJcgVtOpKc1xvM7XzeYqP/dUMfCQFjkD
5uNNl/ZSkIMsFWeGJa5+KZMf3Fz0U+zxKdZXX8tQTOcKZQdFAaEV7YKls+/6a2TgKLwKt39dZ0Rp
/qERTTh5z8mg1nAVD4+6gR6nlBJMxgTaO0GKUMvwsXeMT7+bzYHWiC3o6+ofruHvseZnj9AzRwME
KOHO7aJJVcawUe2+RTZMGt1hCbjjscWDVJqPGCyW2117cVtK1JRQyRyiwz64r90uBcDtOTKRPXvb
+pj3eKk8PPc6XP0j+UFwbeU6dW5I0BmWvzeEj0qg0qCIlvFFKwdJwg98fX9Ug4wcgtACuKMeQDen
qeMpAoT9Wqsx9cL2GV2WsD1uhisCY9nJEE10jNaB2pbvzSSoKASIGP7tpD8pqZ9+tVYMippSl40T
vLt3uqn3hdP+7yOeSy4nSkZqRxfSXZrmGQDCHWgTZPtoB6jngPpKc8eWabU9E7GQctfyMrN/PQt2
HdJQy2tDYbE3ITpnDI0OhQ8WnZSTHt3+QEmPw4vd5iAFC5eQfU6kVapNzLnyd5gOPatGnnoea+Ui
+qLuAp20TPuFwhd8o/L3fC6Mex/CoBL/q8CmbXUs7OtSgzkuXka3Yik5Zuk+khngdKbfa4Avnjkl
Hb2y13kqUiTd35OQWTs8aTekxM2SjKQ1IZp1tArR31tQNSJ3/9ePiqTfmQXBBMvJjl2NNWnO6efH
q6WDYtPUQpg+hM5issQ6oOk5W1YErNUIH91cijxammm8EH5Pq4ejnQYPEbvtOv++S+i5V+eBxsVz
9/hZWtkeaK+rB1GzfiHjXW3LS8aal9tSRG3b31DBScyo+RGz6vgJ5jskBsO6Zc5+nmDHfmKIoLg+
3BA4WPTDI6VnmvfxgTVSiqHJvXuyJIAkQNF22zArcrsMUnLgYep6dCMPW8bE6z3JW0E7hp/CDKXA
55bem38VoDJyjr1RF62i8fsI4cuizR0tGyu7NHzIsvq13I/kxin+ipwxSlaX7nr3mFRI+A/meusF
xRMaG8TxEQZeVfFmH9Fax76n1qkJFFTR2bxa2EUQoFDIPZEvpEhltootNonWZeiwl30c97egO31k
GwZDuGYIj6iw11dlFbvTFYgJ9FV1aUcE59HlgmgDYIamb+haX2Gg8aAHgGLObSR3cxd7LBlAlG2+
pA4rZosd1eIGXICM5DqUl5Mm8yN1UM31C5yUxlE713DCHNtoPmL0BTaAECSu7qG4gvcw3L3SONoM
0EJF4VVZ2Y3NTds1NSaZh+Xp8ZOm1FIhUT7QAwG/le3RFOQCUSW2uvQWDmCK9v0yBmxc1pf0cFpe
rXDDWuazdjn9DFp9vALDb+ryt0s4XgI6k/xXnYhYvbeiRjfn7GIz6z2quu7Fiw79z9UsdOwLNCOv
GkZJ6SpVvhKGG0M4m6Cfi3Z9utnIRkltdeE1qrTmHHFL+v4pqrkePCutMZGjYp1kTI0KaNEVBXJH
uTSu8tlea8waygh0r8l7roIWXqxwGpoIkXtZefRLWXzH/312vv2hSEMZhfG3Olj3sEyYu97fdH+6
5y1vRcmgPkCScK5TwKW5LpkBULNrlEqW2yZ/lLNQ7l38gRuemqaISpSmujGCCu6nIgWT8FV0+tql
A+XMCCqpd58nFl3uZKTQHCcsKgTASuKTmwrYepslLARTP3PNnacuDShnVU9jO8IUpazEAqIZmE+y
yrM/LC9m1sCLghHrGVf92erI8d3k5+6hgQbkaSsw9LB0Jzxzb0TEFLi/jgV45ionFdhRSjkiFBVZ
GVV/pYWLiTJYTo8lK5F0FZE8hqkHNo6UDA2Nh2+skKttbBuH1N9Fl7OmVR/1y9wcmzBT/QGcqAiO
LcgM8+KiZUrT4uHKDHdCHIeabzYoQJr8ogGpW+gK5FiEhKZn04Niire8RkYQIB0FcTOfGXN6dg2Y
HQydvg0Q8IFHEU84V62Z/4eHmdFyGp7ZkcSOPzQxCjDp4AFuFZdElIzj4dHP/VgTFs6Q4AviYt8z
tPftiZLYmYeLx6h27P09jJ37Dd0ewqxaOO3L223eD9c0bDI01xoj0p6GtfCdpTF7DJqi/biyikEe
ClHOK45Iv/M0Xd1/mTli9/HFKddnbxBz8Ma4eWkYsTJmzLetmiyYZn8RqG08p7v7s4ndwKBOZjHp
eaQeICFtM44RkFwU34cIijDlxyxDHJ8lTruhMXjjix2FOAh2mQwIaH1rUTp2rzUeQtZcgrPj6NZn
FAsq7gtoJxzKQvu3Ty0eaE73zSIV1wq3WSU+wp9pbH2zTN/b88+AahoRX3IAh8dom8W4xOHAtlqK
DWJSIXe4IjPzFMtC0JyFDYWoEXMko6ksJ8XuJLKV0biqYJDxJb2odmEPNIymr72b2ac6AgCjQD/m
JpShSU7Dp87Cgy4s9bE5BysrJhwlSKAGOWfDKntjWnqW4CoAcR767EPBaMVajDpT7cqDti0YWIn2
eD76BryTE9BfQ5LF+h0rQar4bJBWNQsHSf05187iTddJ9xdW5H+bWQCAq7oEbTt2pXq/IuDXCG+o
sqixhUbrBG9Acn/+6+kiHiG4zKApRIcUyC4EnVw1ijwsAafwbgYB30lt9QvfY+1Wd24LdezG3G/s
u32GSQ4eeGu8VK4qVCukA7ADdRN+LeIMXS0LMfyzpBhECHHT9Wuer96pWfnEExTUZeD8aRFOCYPW
K5uiVnDUQOOrvkZc3wWGOX3IlCCd9tuzMtN4qkX26YVoxU6n7WTSAN/PA7+AFKpZxCY8DV2mEuBa
9IYIlp0NC8nPbT/+bk2AeVGNTaeKOL169DQzbAnsTxh35uL2FSodARkB3enNQ2Jx8Q7AaOhjZQBb
mxKUN9fAVV2+AEpUUhRCckhe6i+KpvT9/4LcKdhNO8gK5Yv11fnDlzSqfnzuw7EBPwqWke4C/nlk
gfEX3OLVLF+zm5JmBLtzw9rurhjWuFmp3hln/IyQU2kg9/L9kHcoFBjIb612kj3SDsTtaSopwft8
o7PsSVPBkEvpUfmYEnjvdxo18A8oporioBb89ZKA7t3TCXiS4gK/tnPe/RYy77Adr8cR/60Uzsxm
msz3H8O1g8qRpPpiPJfM64ekWwpZK7TIkTGmbFvtzUznvQfvOPe5VCoWqAJgz3hB8r4lga2u03xj
miSZKjJ3X0ge7Rp9HXNyswoFV6cRV9O3FiTVDfLf0fD5zPlm3zu6ausHXEV1XpPCSwtACVleilRM
BwjZISLnAKv3Et4mmkvlkoL+IP+VpuzfJMb0uk0EJW8uAwzUYSWkr6t5/BdbDNZD/YT9BKzaOlJf
oYe8X/ffMS9HxuxoVzD/W9KFlt8qXvCdDlmU/1NBvRoOFlmkuSwMeYb6svOQMWYWxPHRD8DxufYG
DnTc9KPKk6ZIs4Coykw7DM2vTBKPE8T5FJGs2v/s0ibZtjAOjR/9vmCQvhHvwSQiouzMA/75X7AZ
WNZ7Srs2no5YW+UU70uuLvJinBXB1DlL9/7r2T/Pps0wI53fByipb32m+jwrhuRGeZW37tSNZweS
e6y2RR2tFwWBHgcJJEkWRVdaJPj3bfTrkUxx03z+1wUoNWNXxNM/i9TgFH5nszN3g9TzfChpIcWM
6JhCNYadOTX5BUa2L8sJTxiorJhd0IA/eoAQKYwRgqjllHoekHGwIYFcWRG5DOkjNOEd0oTtRjNd
g1K7aGrs38ZI23vQVzzRbjiRD9bU2l2zCPgUh1B8dHav9uiEQ5BUF9PTe4PTFIFhucQhxyomQDQj
g/sd0GSD23/zMS88w6QTpQbxse/qG1aWCGae5OoujEnRqvaCIaDER4jFGgY3uHBDHhziQVVVchjk
Q+NqTPqaJXl44zazO+qIVO0t18Vb92B+W9UyfsUCfVJrQhicEO5oAnXQIqZSvwDkyNLf6PSFhlDy
u8Nl426J4d8lwidDdwJNwmO8JN25QbqtpXrHrQp33Ngs6SixSD3gzFqEdaGOkDtqsTT0k06w3yyP
mfQJZbQOsj3CdrbUsPzhHzEjxGpX8I4BE6lYYNUQ/CGlYYzL/5e0JKc3OpvjwPU/Y2oP/Yc7+V6c
jS1JntPdKflzea1xVLnx+sVP1nSjUMrBYOt1bcIbCI0gpam4v0Soo6aTMClow/U/6lMELNDS7VKy
5ORK36Sj/FectgeMu+tM5V9ujs9i2u5P8B7Guf70oOJLEW1/Cq3soP7YQi64Qma71i4T65lwrBbw
OKgTrdZwTHfQNubFnvGVkILWjQ6oqkDeE4FWHELdZqmdMFZz8TgSW1VrTcLZz3WDhAQDw29ozgzw
XvlwkbywGOwtu6SCyas4F7RYykTGoZI9GXhOMIMBnTOj4lWxgniIUv3/MqXtuktb48hsPMiOsBrj
mKvMOst/LwCBEHOX0Af/1NPyiHEyuU+Wq4XxRrl7HQecpsQ5pz59idHSw+2LG+4xpJHoiv+Uzyx8
WGZ6Z3iYYdELgosxq9BgqmOjLTdfKzY74th5n/3zkJsLfSMn1sGnzoQzFgOFuORKyUXX0Of0nuwl
U+1yykoj4FQQiQU/lrXYGLRlrYFKquxgxP/ymfelRufNOYcpGuDZwEPBZiBZiBmgSn7Y2ZovtJOx
aP274aNr7s/nFRTJgnUHYeDGzb5ULKOscQWccgmLJnIlOjScjq4CZULOeZLrXlPtZ4ETmoMsiO/u
sWaqREpGxcWnY4EmVUB9rIJrHORdBZud4x7y5xmehfggu/bNP3HJrN0J/iUP1/fZtbae3MzrTXYz
JuDSeM6IeKDZHEmHLxRBDhzmxx/Ra3hh4Z077sPZf1hJDfbHmhUkG0AIvZmW5oVUNv9UwIAJIwT8
QMwHiF7OSz/B5ZuF67aGUWaRzOeaBDlaiXDESFn15Tk61D1n5Non4twv6OrQhckXMl5tznCyCQ9c
8R0Bcq51rplk7fg1/pIZrA+ImXScnByk0SpOshhhJqFYoCuSbtW6IAy0WlNaMppdWDj2pIftdq26
41bs3hrFB+hY5in5fT8bxB3I7rPOCgsvUA+/WPYOg69dzgEuaQrcSiid/jyfwNYNckktw7uVcVlM
yAnIZOZCvgdxSeZhs4Lsw8IMKGeXPSeAVEozcNVINqGqzHcub1dRJaxi7Fq4DENl81olI7oNoIsr
UYRlJbeHYTS0yaa5AUKo4tUF+S0ClNBfrKiNCbGvv+Sf/p9p/px76y8BZvDOf3u0rY0Xquecko9I
s9waoh2NNrgL46IxWbUzGMbMx0xoNqS+w0A+YInraVzDr5q3j1mvP6ORhaufWj7Bn80tagcCFfd6
7RmNVldPZmmBkUrpDOzi1h5yhuu+JRhVIOide6v8Oq8c/ThA9sFgUJD5pw5Ohz3AP+PJR1AMLTfT
9MWkZEcFEHEdsaBmR76Uzv9WL2r7iQxcFEHN66zByQJO8h1CmHc6PxVPsy1uP53+RvZc9d9hqP4i
NZuT+2oJUm5sYeViQKSRaBpxRNqGZMfBhQYibxn3BYC2/OuW1mNEZvgZnwssKMciA1jxGpbugU49
pklWcjiQwcJ3FLb45K6l1D4GKWNvCn4lIztZKkBKa22sTK7XmNOAVwqoMoMRA0RaL3ImlFipK9AK
amiZh7qNtNAgClIagdUJ/ykeJlGBzdsLVl9ezfKOWiqpDO4CGHKILYD9MfChoNpx2kGnqaI0zqgk
kT5dD+nGsZ2VFwu/djTrHKwNd+YLmU+Ll7JJe/CHXd3/5uRsDe18xUMavb+M6s2VlNejhfx0tpBX
GMF+4ZU5uyNAYNQ+rSZaNYSAjGsKAm4c1BXaSDuulK4qz5sINt52vXQ67KR+HqHFW9spKh3d9gOR
t/RM/MoZZDZYvwNO7GA9o32SQq/cxqt7rlepmQYn+kJS8/z4b5M6jKM4GaAZLo9ZftoL+hoMhM1O
Lq4x+sUVkruFsSMlM2gFGGAv81xPUqPP6x0qLRBypvXHzFMcBdKV8ZZX4HfovwE8HZATQjp5lj60
ouMjR2ozBt9xCZ2hNBpU7JHssCuNyBxXVDzAgd8gXZXgFTx2u1shKlez7sG3rRNuPBB5HvdQr4H6
wxtVK+yPgXPzQZ5m92Vjoku+campByAE8aRjjrnkQuv7a8GSAgV6uJggFpHBMIPd3SSMzCVoTH5Y
7GdgABSsb7cWW7ZDA3IgUFiA8hp/OdnKLBtqIJEBazo1ljR7soL12Q+P9oJFQhMGtYKAF3iaj8yQ
y6nZ/aypskKNQTLBb5HpjPDJ1BflGoviqB5AJMZC3sfJWkPQ79VxBGwqoK0Lv2zFUx9sUyzQBc8g
LApCGvTAdB1D2UIWGa3u/4ELQ7B60gSjIiUigaQpdewwPX8TYh0WODk9Um6B+ts4pqkIk5kapYux
+WZqTwwcGC8Mtkm1U7u1M83V+PWdmzLKfyEUDiL5TbpDl+07rJeYrHe8CSWmllghQ6P2GRn2bMNj
JGZ8QEmxVJVKFPnlei2jgcXWA2fYOrwL9+11rhr5HzxsDSNsMh918lf386dOxGNK4IbusihkIIdv
HGcJL85LUAVsiAE9D3eisZST+h9WhxwEWW2DExqTd5SWvSmu/vzGcc3Dg5Lnh7sQo3vYlmt6GhX2
BsbyPROvUemKbdVZgCZySlb4FqvS+ABw5vEv94Q/s9CIRqMz5StuK/6Ej3D/nobMQpmua1S9DmLE
QObTiG++YrcEUsSKCQ0TjGOjiGU4tSAEwry99Ew9MsYB829B71/ig4TVVnzZsHzaCuWOyZ2E48CZ
qs+75PSD0meX4C8G5Qs0mMr6i2zqifajVnpI4IU81yIngzok45cbSRzH4/E2wToykn0r8VyAXe2N
0dcNnB3IQN+D6n+t7yGNORuFwqhl662sgpPH1D0Ug8TCf+a4V+C8uTd0lO3p+rI+e+YzJiLjlgRi
iOc4k5Wd9qtk6Mn4XIWsT+MVg3xRej7VyL3V2DXJ1JONgApg+T5DYDb+4UEvZkIpRSZXLDMDxRX+
jkMg3wxCuac9FIfaGyPMLYBUz0Ecj13R/9tv/QJllFweEb5965V9/T1r8zcKRsVLkj3hgnMmxBK7
r7dbUX4o7NRb/1+nJRLkIRx2qmg3EIqbhCxpdjre0tRHXZS75StY6fEHf9/4WGvJBLGTk7t5mLt9
9HHpdrxEkPJadz506HzzuHE5yDqf2I2vnQWLCC6r/9e5F55d4pUPjyfO4E+xzD6U1c9+Nt3Mk7Rh
YdDEwbolZjeP9U7P2LeFoJJBQywiZCdaQ90HORH3OcDmWl4qBTjuWi6I50gHqbun7K9WhelkXLg8
cLF3+609sxDeO/7ZjyK9wpR2vtyj+5oO67lMdBzev5IocKLP9QGwmYaLhBrtVczSzJZyDl/Tqj/S
uDBY0RAO7q6rt8vcwsBRGqzIO54QKXJSfU/RqAOu8iTfERMmYkMNxYoqwqb2SewfXzLkh93/xkFb
hAz+V2J+zbczThTwgYYFRqvUO5//3M0hXydeTBh8T8PJ3I05AdoHbuqM26M/h+bkXO2dXvCxLBXe
GdxtJhGD2gAMYnkJOlNzjLzzlSlV+oePS1fXoU6eSZ98BuNOriuR0Ce6BXG/2aQbKaxEx3eQ19vG
aFrP4o8rwnc4jQ4pE9V6FFmJiyW2KNw16cpWJO98Q5fyfDWQnZy/sP2HxQjaTZfX7/rG4IVBXL4I
ZZOxc6iaIsIDNIlLAf0EUPMgsmaMmGryx/v0Mbhq/U6lB3wGvdF5uTGUy0xU0u5GY11eddV8Qiew
0DkmZ0vpDGuAQQDSY2Bqcq4+v5ZoKmxlJ8aAHOHB62Aa4T4Ie18iMRtsqQ5gbbp3YyGFbpwwo0zt
P5kZA4gP2rqb0/uDAlrfpQauUiEv45MQJnzaXjlTisdrv8dEaOfgZSbLm2gAR51m4vAO7eN/In6q
LLxsOQDfwVEWZyt1hP51MomXHul3zlWNHAK63ZMlRlTKaeZqRp2xQekl04465cYr+mOFYVXKoTTo
hSdsWjPeQyM5MMG1SJD1/G6NhFVaOPz5X9+PEIecrOlEj30kdmkZ750ubB0Ae/nk/9AVRtb/4EHr
hC6+0reRvrx6sZXwbmsJGTvnCv46rOsieIVj+ZhVN4T73yAnwhbwDdROdSxJ4RaGw5FnMrw/vU8i
sBB2l6QvrLoBSy+UjASxWDSGu9NtSTRMQWCA9FoMawbDNviOcJRV3wKsrw2bjuvt+T6+LL7wturL
gh7inpU9InsosmXQBUWQx93xDj466L5to3cncfbFT8NhBrBoWwJmMbj+xfBsDrzXqhqxsgOVG1EP
cIErrj05CFTz/Z6cHPmnCcZLWO1ZuGcOlyyRKGGJamAcRUlui17kfhL021PSUaitQ5cXV0pW7kky
d4AM8zJ0+yxnEZabUJ4uqylNCfNQxWYs+iDCQYhdFNY1nAh8pk6NR/47b9LvAxBbqDxI/K4fKkwk
dhGYlfKRar5JOVEt0Yf2LxapVAvweVrEmHFU0gok2K3ngM/b0fEet1Nr6KFio0ppJcwNPQLJpq+u
1BYeznfD0sFEE/0cdhqf0iAMVM/EhCr2oG06ovmwfVjKgtjG9xl7UlIvybGcPuSXh/Ayf7PO2vL8
7kuDv4ZkolZx2ol4UGRYvrNsZoeitxHIaa7odiLAhEUjxJkNw0mAM2C85N23D+HPMKLRMbfmwS6w
ENKNF4KrmFzwVotpS3+vWscep6Wqg6BPfgbW1ip9UDLOIO8KvhgHImNKMh5VWR7gaJsjpIpamz82
0tfOfBSB3HiU5NuS4twAJi+HKPKYevvQuzp4n0pWMB1/XqEZnlf0nzrSGdGDdOOq0++TnxKmMKtl
RZUOOlBqoqSD45+W09uzn2C9PPCH+hgNBV2ikXF9z4/PB8Ckl97uk2KDnE3fH2kGOgMBdYG52Lys
FUioQ74hwY/C/aduhXDkpOqM5hNX36IAEhPBkCGUsZq5lp+ZnoS1XonODqSRy5bhU75Z13DN+ije
54K3VGC52uF8eC8ODmZ5kgXmhJEf3rD9qT4h12WHMUanRIdrjHqAbDImWvG/oCyKdqd75acAeGSG
qBTOpmkBuUANVkKStcqRnt9ih8ri0TMRn25AUggGhRUBTPEYvyT673lJbAlVNgrj7j3k2OV5YkTN
GEtRBFbefz+8/toBm2IJ3OfNBJ3tX4W7fPEInutkmFH+SnyA+g9YP7MgBBQS131VMpyB1luvWcXZ
wJT1F9FgWBS3XSUAaGCYbahfWDaeTfNgPPnh4GCrxwPlVofKXF37LPAofxTyjKK0CA05iVTdCcCm
ONfNeyz9ZzkeORBb0NMGyMv+7aiB/XV1DCG4qRXunLIjEobbX9YNilMPN5Nfp1H+FkkMXB9wRV7a
Z9rU8edjAYCgL539MLKogWwzAsLKpYeL/0P6ky/74LCvBt6dxKVY7V5vAhXT/wY8CX/5quazeIjg
C7udTx8Pyuvh0G9++pA6+nZruuOVNxNGCTxmhoWSZQCPct+mp9IW8AsMH45RzWyni34GmCvYOOzT
G424Wg9JlTfBVw+2gAsoSZ2vTAHWt4TNEXCXl/AJbVMsLF3S3dsWLJ79E6RHOLbN6Yrp7+Y82iYN
v33F/zZNNFsVNRvG92kSzlsIkJiqlvSqMMz/84gxQdOwofyYOIGMiVCF0lFrRdjSM80LzPQnqK2L
ipyufgDKqgl67lm+VnQuCkymlXaM/q2pUOWRpRBB4LJsd208r6m3e03ne7rEl1avBdOHxRsATUWR
nQCK03ddtNuDz89n81EXwqG2sG7vKoMQRkWuOsrnWjOvJh8/vGmcFSQg/D9VlZCyO1lgOIIGTQ3s
FUWfLgEXfW+1hZfqvTOcJ8T490gr09yp6qrm3LLurGJor1vk62jBAmxjnF2wMlDuuOC0SDq+vW0w
hZm3HvevzxxPaRySMfpNsWGaG5XprveY5HdQBZPWpYzXtcvAN7xBkI8L9Qn8KbfoYKygiGVO64yK
IF4LFSKidDOGVELcZJ+tcx8JG5tGVI2o6qqArD48FNj4EJeo+MHoFP89gZ6cQjynpLmkoecossgL
rVV7jIy8qGIWAtB7nLfW2g7aNzE1NfMbDF1p9+XBp1RbyKiV8sVUkQLDm5KI0vOSSU7ERkX2XQTC
VUSOxBeUvRDt5hHAam8tmOmvrsbe7gw6VFozjuJwGukKITQ0H4UpXxC7j+5jWE/grZqzb+SgaVBC
8JksZpdzpW4jj4KGfNeGZ8f/XRLCx6nxsvcB5x/3EKukAVFfzpquFFdtOu3jdA0uo9ysT5i/4r1g
3qatymmH3X2ouAVSZkqgy6tn68CBhStePzdaXUFHmjZnx+/j3eWoJ2Fdt71P6lf+ofxJybhCtVf9
RKZHx3aijf68SOpR0MoV1olP59DQH5vKN+8auTvgfVQ9di5wMG/qUf7BfovNvC6TZ3zNuKvGCVYo
3bqkbLfuKgh1XGBKrPDIacs6Y0xVQY755Tkd6w3ksWDh8abILVEsfV9A5ykDXxsN7aKSfjb7XTwz
FdM76m/+lzVF93mg5fFxr7C1Zd60xJjTe0CX9a7mYL3mYYOrv5wjHBy2mtOfuHaNIOiSy8XmigTi
icS/2D1r18cO0gYFmTUsq3AM089W9DJfU/LMnwiUYXUwZWNhKD6ea+dOOVb8zmvfkMpyqsryR9co
S3L/Q/gfYoWgls1PyH8AxBJNnBzSxY2cP/f913BLsAj8tDRVBAaVSLHhLbvxGbFEXtLNAQgo0G9U
Lss9LJBdrSyrj5QHs3sKbuxtdOLhydPaAYYPanD0W91BCb/cJypBth+rgiFewAS+q+72U1fI76lP
tXdHOokiOL0EAiOeOcm9by+DVzn7O95hhMEbCYHW4Xi5e8zyklLMk7gfZjgEtMIHHeAmJnExzIaR
KqZHjR4f3sgjr85oY/Cl4FjV0kW3ln8i/plvwfV47QOIvWWu7ni7Eo52pz/sjZnC8+eJkY9ujqYW
eMM8W6GouoaQ8eznpPQ4m4/p5auR/OE6s7oc/dbN1TurYrQQOoCgmqgoIuLwVSI4e0Tpq+tuwC9l
jSEJkV+GUDnqPiZDfXtu2qa3yIfKCNRQw67dhiQiK+nLuwARPwxgdkKwjB2tiPTYl5Ggw/CkvK6b
eui1dcZvrKkOP6VpZU93IQvuZMCoO/nnal0sX2736MsLbbsM0IyGGAVy+uWwkX1b8o1M4ymtDG62
Er8ZabMOavVVJnzKWU3y9mcZQCqmPcnZlAiIp6qWBIysP0CYtnzBN9n42VgGd0VfR4jAOFzbLGev
rv0MRAm5z0xU6ZdpoVqsY16HgCFdzo6iVcmDN8OdKgMH95fmYdA/nO6oqkM1EhdH4bPGiw7LzFqL
dPCfPW+QzmWuFejLk6OymHrYcISU3PNyH3SZ7gQT88eZG77204aMwoTtj9l/4YrwpE3ytBMOHl5I
UJ1fp0U4kFwnM0cW35K4kVFY/T6DnQ5YvqP9PrAucxUmQvDA8ZFxyW+UStEG+pEHHeVtaXlD4Ka/
64aokeP4oYAFzHeSl1yqbMgXDRkqjBel4VBA93Dq3LsRjEPtUOwNTx+3Xz5b2pWcw51W1SPS815+
fy4y0pxtKkPUJZWHe2DlWukFfRE0Xs5+4uybSSBjsLwVOBFDfETjKd+efm1DyUlsxxIM3Qfxh6Ov
atgTdWB/VH+rnDnNfsWbVTNrCsMPGjYM1VhbDkqc+KoScd6s0YbKafnuAKDmPZuq5T1FW2IIIdVj
v8BdB2UgJ954zsVGdRx+GCWvLkgePU7KnrWSmD4uHx4AOLOcyLNVAL7eAunREjk+vmrWF2e6yEYm
NzM6ANrsjbhXwDCuxfGhobzUrRtGZ11XRYg3xmphvOSomEyUK2BDYWkIXGe0FKGQQYt1aHHYiD8n
84C2r8/oEzD6G6DELtiINpXcaOnGxyN3HgVtV9nX5qN4Y+YoskZrEoHeupN+Er+iFQC7H9vylNKv
E+AAsbhmsfTqfz8oTXALA/mM7/vIymkhPtAFTPWAuAtQSgsleaK3QNMgKD89V0W/DU9fYxOggAkp
u+hUq83Tj88LYDFyhhdmEY+BKwj/jMGVMgZZdDeMLInX+VwyxyCl1F8CDb7S8daQKIlHHNd0aSbi
JbY7JhnXckfljJqjfXw6c5SLqVO3nuL4PnCrcJSEQWOvlkjfJcHg5R3Jh421U2QMxIHsWLcEo96Q
SZNfmA84voo/4G71pVSZsu/JvMn3fyLEUa9jxmqZeJf4J6xNpAVR4DVIzgyHhyZ8UqtnFJ6XInbr
1NlcVTlgh/wyA7vdABV17FDpL3zAuYUoebSq3pgVkcym69uYsm6D2XpKIYRTDqOdcZXHa1b8Jtzs
401r69vyEP2MU0jHcyorimoyiiy3KG+J/2AiaeZ0hGlFtf/3W/9Cbya3pCRhArdtAbKGLgOTt4QL
UDsotGsDG4rfZFzgdadOGg+xma++EjKeVRjtxmFgAPzN+o93YRdmSAzKf/z9DeR32MThXxqWj6mW
R3CPrFMUK1A2yGO29pG8Y5gIUydL79IKR4b2iLIjojAl2FF3IBosDLoVuwV/cDO9GT+D2RO5IWPk
Q7d9v8DgwVsmHXBfoRyLTqwC8r95FcUou5xmxIIgnRPOTYZY7fpB6XJkLsf9Z8TKzc9H1AlcrRoI
xkv3Tsgu+gJZPbTKPZUzqreRkN2tHUGhMi1VXu+EDECMdGdKDDWvvhzoHKkELbIBPQ7bCBY5Xf8h
Hxe2IoUEmWN7vwAGoajJ9ebhW6lEyGGe2HIzpOGxReB8D5EXWm6SgDF16XLd66FlO9pbt1EELV7d
RwLAZH9EZJn29cywEeC/+Lxp1XcQIGxp52ODyJycLBUZzBiBo7fY/GQSecovtQqNcqf5OlafEl24
zpmAYBkXV4NLEhg3OV5//jmgeFdvKKEBwVWuUhN6w4n+f4wzsN2cfHJAIuCItTWW9j3brqxtgsYg
ufhfHFQOgLC/Kwo0XnXJzz4wlNeY1iz+wLbrFHergtQTlXrolFg3lt2195yiChCcHu/29ALwmV9q
wz7UP6al1r+V5haDB1U604ada1YI8vBoJwrv7zD5un6VXkwLRvDDvrtwu2DbjI5bcnd8/+1wtYko
ZVX0GTQdnoVpTQ5xKp3FRKvGmy61kFpRtDpKDlhVczRo8eQQ2F2PLNYC2IZ2moyfYhDKHLoLf212
gTTxvTdJH1Qf8nJmukl5EeZszYrF+Q2jAHFkfKkzvBKFPb0vfrCnFjVsHLoFtXxixX48i6u+TM33
KAQgRSfL+miom5cHZL+BE0whNgAlDvnbbQFWB9dPWWvvg1iUnnaLW1sKMM8NlGqjcwL22LSKGPfJ
vrj+SY9Tq+YkW7fBrycwxOO/61li6t93txFIZWSVrbVni9ZmnpCrPpXxARZRqNPx+zYVWNB5EiXO
+iu76f0q7L9muLtoYD9YkAzJsEuAX3kQcVCyKfB9ZzyyCaqBxegdoMmFmRxmVb+gm+HOBIadFyoU
rOA9DY+4TZob657nlmkfGNj2buoh42qiwLJYOnqkx281BjquSNfbfGrvcmFjjIVuKK/h4tUQrLS1
bDLeIS8kqADudXvKWDm44AHcggp8NJ4aOhGfIfSxT4X3MfA9CBcxSZw1MnKVzQyPbzvCJFVBYJ8g
nWOr+aiRmAXQhvyP5goPJQrz9hbtTMorAj9aLKkEd4BJ//KUlFxUUjhM4TbAC1uECoylbqNYhLZm
uPkOhV7aU9uM2KKabMpPBr6nkWX49hO/56m6DBniiukWWMPb65Jgr0tFzRVOzthf059cJzDLNmrg
jsC24w4qU3qMTNTWeEDk79fyshbhRcPmZClHOFyUw+zTWJWSL0D97D/p/4p/mvUVkTX05hAQAe7n
KlGjxLLXq29/k1KResG9kAYaS5Xfucrjp0Ip31n4wXQUfBiAJ296DFSMV0pn2qdPr5hdHLmOOl2D
X8S1ydbZBrWBngtgCL1TBnSyGXcrlGF50uAD1NRv3OHyjcwofEUy+exubXzEFXYIkbqaTmPNTQBQ
GRQ/lH8NvML6ybfvJOt0ZD8V/RR+2L+/Df6YUjh7+v4f1K+RTyFXaB4JXgZBtE/OdLQqoaA59a46
G+SLfm4ilU4QRNxQR9y3/DvrD2hWJTklIxxY/0wXAN4MZt4Mf5nUo7HqoSF/SkRDgqfIjHKuTjpU
RDUguPkveMJLx/9v4Gm0gjI4vN8NqQhrnN6SKbmXsXiu7Y51X5gUf4O0N5ukORgFnkEqoecsig2Z
fxUpZz73R8ZgIeYOlrjAy7k+yNsd3Qpl5sFiUdAV5sWxG00hP5+mpXJntNhovobM13hGyxY7RdRp
pMEdTmLwy/CE+9EL8q/1l8CAafuaB5RGcMqkjnCSEa1Wuk2tjzqDs4SmcJ//FVWeF+juMnZFJkpt
0jDIA7Mv7EBHTS9tWs+MV3mOcFQphcJeYj4TpkXBazJqEijf5a9+qrXRTsn6x3UVJCyec8ALWplo
XiH2t9vEh699m7lfgiNtyydITxlG71yg+VLRaUvfwwOuYziebn2Ysa0tkKhbYIcwXp0xfB7Yy93J
pGAH0btI3K0krA5xomg3u95i9eiALWL64gMNzK1lbAuf1L5XM9hWGR/Iygm7D+WPOxlr9naBQBD2
t9lbsuzNbIbPWxIyiXOFDChExX/87ZwrJwtjpMf8OfOl5myVJfe5fBsuAWvtP2sZE5ckT7z8DLmw
O/aOarJQLNkFO0Pmyo/lr0z+yQ2tT/pS8pEk7GSeP18kIXXGBvXkgxKf8v5dyLzk3syYHkA4XXf3
qKsvx0W61DGfM5gt6P4D8ewHfIFO2wo/b1AlMy9unUIAAXJtcjWZVc/bMy4JTkw/LXEmhfExrtV1
EWraWeZyJxIX1AfEmpmaV+mj/lTpNd5EjIZ9QUcTkbMdHFtvzBrLMGIFmWNNRsor5kMst9wQRiFE
LT3cijEd2qETvvTkKOIqqL5NYqO8RiZcTlvH9ZYNdIkgsdhE0i5k3IsZKNIkOJMORPypVTOSskES
5MUkcQ8zjQOQlSamSbmUuhAZP2l/7XklU6IUKfpb+CTzuUnIrZbHQ5eKLVgZKPj/YD4G3UxbOh1Q
UzucHQLinP4Q9F684fhHEnHY4mHPZ/aUAF+HHaBsqThuekQ7Bmtzyu7/Y+Oot8Bzhv8cxMjpTNh1
E0q3vdd1IqySox8QG7LokMpqiNkJHKPm+mLMgDJGk0ALAxHOJWhBlVFL/rtgIqsQ0YOBNw9ICU+y
cyMTId0UfY2jxCp8ZHAOMQWZZWp/237w8buZBVwfyzbdXIYYl6xQaBZMvugJG6K71Yb6odxwCw/K
jK41LunhaI5kpZOawsoqYng9GjD2seIw1wPXjeo/MgPhH+YOgIWfSdq3U4vz++kXyxwRT610T/wG
irbHUMDHWPNilkjwZhna2gL+NK16chyiLBxX+22ODhdlE/rlDJfsM/9TziHJtuU5ngHAaWutamAr
gx3UgDza9HZZlL5e8X/OlCzIAFLDPgwZgTrRU1QsXy+C0ORnK1WzAch8KhArEfjWd80o2hf8nrBm
bJ/l+TGwMrs9rI3Ee+RijVSdM1SqrMaLOLjy0yiyiuRtWslQd/tNrAWgBVwR2wr3JA2j/c4hvyEg
PqEc2GQ41r5G9/vAZxsDNchd8H59kuBK6UkL1fhEmwiGq4+e0SzL4BD2tSeMS0txHXxzsM+nYC2N
LP/MXvu63DxVMWMJTf6LbOqP9xmEBmfqZhpOu0dU5jlbPkLZruP/MWLjddbzfWKh/oBuSy5m7vZ4
YKeYNEuFpRA+npywpIQPlQh6Elj2sPNhoKp/9JQveeNDni53dxgjfSmJ1ynLDMeadjte2Qw5bT9H
lTVavRH5oDTlIc5s4XKUSuP7otg/Bg1l9KtNtrLcCL27+hOXnbivVWKF3SR6bpy4Kxl3MypUmZCE
OLOEkwYyhXZ3XHqTDw2+hSljQFieJLzJqM60x4so/l6m1qCX3Pvki6faHuGCpmZX+1YWL1oeJXrI
8cZurWbHv4eJKzVvxLYyTqamolcPwhwsZiKRA1Hi5HEmt7bvgeKHaFaR6WspNm6Ciys3QHYDcV5b
8jf1ii+uZ5pABp22zDWMQU8yLfzDGcHKyR0CCW6RyKl+lhMAMVreT7wG0StZr7DM+l6Qq2RBEWNe
uV1WE+D35d8y8yxRgQcEBXd+iGC57qNHSxGjm+D45Q7gF+U74/TJQ0h1F4Ix7bxBXXwRBT8zNAYp
XF73C+ui5G8LchZ9osXYefAlEnafD4h0SEF6TOOWNmvbO+hJnYxIiBR9Wx9AZ3aZzJ6Fe157HbVX
2Km4piGwz8YJfF0ZGG8l57jgEedeLDCPQzNHgscJD19k++QhY1HlJOVPxBUohRZIH9/ltT3HHbse
XnVTGanuRObRTi4Lp+UqXnH3+8IDFEEHI2HSHYCmH9DVfFq5lrSJS3KFW7WBxeuUas+KDyUFfnbZ
mY2o4tZDMFdWtoQlv9Xys4heldCPxFL27kWsDH1l/iakZd6aRpTY+k7/DyeF/ckcjGZeE0MN9mMj
g+pvPSkIKoXCIjmAD0y40SIYRuEsdDZFBSrU/OYSEqqPT6DHESH74EsdWUj1f1EJ6pCs3wXUjZww
WTlPDQiR1Q/oKXZuE2BEvoJLietnUv6cgG5iwzDVqLQ6JgDA67t60Vxy7cnP1/WWgpe76Y6KLlha
wXHxfR1uhlsrXWkUmn8sx9vbIk+SQBbZqJfxuZn5j2ZMrsrV8V/HZao1ttfcwcSPAsH+Njmze82N
9JnjIg2azvJx1jP4ZYf/GPNyCN1KVEnSedizeedF717nkTFeOvHCmUv/xNmfkpDBOAl9k90TeRFy
3xADvbFrx+zlHO8kFkiLqrqr2ynP4HPov9Vul1uV4tuOHoczlEBuq5zTARUwtD4LLthu3jU/753q
/bSVYYraM4IjjMBo+NWR7RHMN4du4bnxKzoSakZzPTWSWWofwGBZBb32J3Onxk67ebucS/hKxrzt
QA1hviaj7EyRLArIv+xMc9qLPqCoZMxGoP25IZ/udB2Ame4kpkeTm7TTJtMYNhyyOUf6yWFAkwW5
NAyHf3haVlfmac3bktdWdCMkhtkiJcSqcsFxngheiMYOBOhU3dIN+w/MiGceu30nfsmqFCGdb5pl
h7ZBp9hEAz6WkiPtcjriXSLwv9PpYhGODIbnwA70phPWrwP+vmMcRuSclh9nD6k+JFnGzM474lSH
unmxt/sdOKvEFQKVbbPrzyoK8FJIK0lCw2eRV1qUc9MPxmb4nak4jk28USaf+swM9GTCsBWWmmZR
o76D3ArIfHgXDxgsY9Tgyaz1ikzHe6sT+wB6Coa8Jd/JiKyvLV/zKTaRFdbB3jc1YF6wGbKvmfxz
xrlwVVg3xAMyPUj8gfwJaN3Rpc9IjJRCOmeznNkKCUHZUQm+sKr8CJT5+jQP15AT9FOAotshGcZO
wVjZFCGNVEtfD5l0UYwq7YP/TFWgHsnnFmFHW4aVafghDB2fMRDIpjeFzPYfTfi8g6phpKqc8lpL
r+Z4p5nk+6/RMOWJrFXmNjArgJPLhLBFdOb83ra/6+UIYi/aYg5vzzVEgSpYpIZQ3nLGXBfTBwbn
KMgzpCVJzqgFRb5IgRjGC9Q2QLsTMzPPwYDfRt92BmmPw+pRLbtJp4Jts4246Ze9nM6fWEXkrqeV
ggI5HzXRfzUCBEPSUvnbgkNVkEUuZbCCW4D5I548VGH1ejUS6zxdQOoyn5UV0Iv1EmZGzzqk1NW2
qijsAJFmhbD8umAaahPkAgbcdhItAjdcSrPs7PBTp6VgNU0m8mZVZKZjzfozU+7L1xKuVhkw5Fip
UP6tuI1nto4Ii6wRQ3DJa5aRJ4GOzJMDFyci0t0Px67kSXm/W4Lm2bd0sazsinLgqrEdWsLX8Am0
cCK+DhQcJ0tetMb5U4B3E+3MMmXMdyLeDR1XV6mSVYzgjV5eCifT5QLk9592biBCtJ7kQTts8bz4
rrp67aAzEtWiKQkW10POnaZMzMZMpv3y9HZROnNX5ge9AjdR8tRmUbEXVxwB6qEOoLrBpPg8sjsR
x4Hqen1XB2vCA7X1XQ5vhBxCgKg0yPzUzfxjkcC9rDX0gCEN5j1z+v82bjy9SdJpiKBpB49bGspw
+vkWF1eWncdndMRebUGHz4Zpl0hWepDqU1MSuRv1PHdzgN21KOKYA+UuJ3GWa9AkitcGPAVCujnf
wXFfz1Ao9T10D+GcnM8o3qrrWwd/aMdpm9zvJ79QO8oFNexGjx08JY9bQcnZtE/hy87h+5Be99qc
30E8Dx2Dr3GwB3YovDw755GpfLbT8fqqtTCTj43NnPa4XNgyvpx35BTXNEX6qfS8/I/O/Lw+ak4L
OR4B0GrwxXIZo6IQwP9D5LVLw5SFGXNXYb+igGtEqP+c5yQ9Iv1gxixsYTbuSqKwLZuwzUXw7Y3F
4kqv/2sgA1ncfeaMgwt22J0RR+MAdPbc+eJMDu9cQUqqWW57viTbjdndBRqSGldrsQo2HfAQvnC0
8J5YuMz2kER+K9PYu4Q4NO8Y8MsKBItuQWlBlmzRgioDDKBJPr6BVjk9Ol/KAyD5vAD/cdgbFoFK
CRT1NxZ6ivMUvr+y0FF/kb0W15RQfIRGue00padCgwFLmYy7Rsmdw6wQ2sgbhS4pXkQ241AM/dBy
eCFUO+ZY6eBd8DM7QXLFS4zGYEN85gm+6gThLnjahWAZWoCIxDkuLINy0gpTl2oFPen/youGFN3s
Z9WHIM7qiraZnvgdh4NYOn9IvL0J9ozbKfhDu3pSJPmnFCqmDdNV0C+xIqxWyGGFNP00GsI6/LQ3
yfJknelwHSoM66dxgqOHeuMOOD6tX4cujOl0UuUpEW0j8NuTK1s6TV/M+kkt5DT9mXsUCeeMOA/E
Pc/XB8bbskMdkwTq2BetchtMLQSmQLv4wxe/WYWmmnKK+28Xr+1AyX+nHwZROsD+jQF29gRH7nGJ
9PdXNcSqDgTPk/csr6w77SXegk6Sgys2lusJTIbZO5Oq9pNEi/+u0uRQy6a/gqdZozzJeia/3hPw
40jJ4Dauu6MHn89dIwydH5jt0mnYMlgS0xtDPBKuahU0tQzuByNYoUZfGouey5QWwhe1IlTXlsgf
axPz2psGii/jpF8rWX2u+L8Gx1FfZcndmcrjZ97rRgqkG2ZRGJZKwEGWDkPBxa+LwBArJseQHLs5
JPQqHBjZRiNGJcrA0xZW3K5gzVJ8cNWpiOIj7OAWJzoE1XGUk6hYE71psTxunUSUJVTYwJ2hPIpj
3+yRvpe+3wgbpIPbZfAsM61uC5Z7bm4GQvSc+clU0V5YiGX1y3Y7X/zDXUmPtbBUgwCCR66AhHIF
+UBwxPJX2ShTjHsmHPDHp6cWalIF7rEViReUv1AwXtM2AzNpV6yPl5l7DFX1cO3J259ZJc7/8Kwn
/jT5p3sUmh5IXuaAKp3ETh3KBTCeNUFRW/SriAxul1nfYPJjhXlIJr/HW2eSwKmVxuDqaDf/rMKQ
7rcuiZvOiSt7ZBnunLKbrOXBEjygvFId7brmYBEHETjZoH7aITZPxHiUPOmMOlMNWynPHJjT/BWr
UtEjrrn8jCAF0N8xzbXJpPh5Z4E4+1PLEilMh457p1Ysx/EsNih/oT68ZHeVFnU63Y+vRqYzLJ44
UrDF3ki6SX8iAWnx+KD5PO39dLt+0SqxlhlT3ZzvxgTu+vfuM5dkY66cSHlXqa90fFNcLawNMk/O
z5TcPveAVrOfjK+NWzRrjsUCo6Xhr+9SzCBujQwEBzYy4y3nQKQEElbbtoMKkpBc5dGfXkzKPFhQ
lAg5WnF0w5N/qDIeVw7iPl/u15B2CCjJ94/O/ov5aZ3/DeyPsSj0IFSpB4QFywDoab42L01VyYFj
+2OqisqUCz1LKzuBCL9hCQzjWlwWEan+/qrU6Qtsq04c2lrStUAtf2s97iKHKJ8UwvQu+yRY/XO0
AqeLSMyU2gm70y+NI5UE4N8T8XqXSSH4NQwMXoWJ+N6Ol0sRhin2aTYgKYoWSsh7vv+Ujp100+Dv
Hbhu+AhXYiT5msw0IuBVGxyHU4ZLCFuzE/zMOQIv30erkGmQ9aJLlAd6/ZgB8TQGqRXwHwjkof8g
SwjUt6YJxRgEyFNyb4l+tx9dfaqVroKDzU875ullc6d3wUXXAZloSRYolXNuqapPY1yS9UGqmLbg
CXJ8ZiSnxUm0TX9T4FIre4Med6JPUDMJ4qUcsqu1LEJrRl3+LP9YfWV/hne9eiccxohGSiPWKrB8
bsHS8Bzj865R/gYHI1bzrFvxxUEbfN+bPcfOmMjv9W5k76A+hTZ0dTWjzFkswxiAYfGO0NFSwKLk
O9xZh7lqlUtY6s4qL3vrVIqBw/q/3iANeXCWLjIYOQwQskbnJF9N9gZtZhQ3CCeLaJXdpXGp3J+t
IkKJxkARel4p9fva6QmV9ScMBa9+o2h5DkQ+O959v2LKgbOb4soqyYDLOzRXLfBjRW74q0qzkM/f
cNElFEa4Z600lLpSo4h+0czktNnHNj7R1QKgaWg+jSEoxo/2lZTPuwDG3+rTBlIu1PFp6V5W6jK0
ZGk4b6ksGx3ZqCKClGkRQ5T+cg6sTgGyF94nXbUNo3OgzIhO2EzhFiizwFsXlFB1zEQYOS0fctpx
yhpd58DvxsSrznM2+T0Dtw83vvbhp/EkAnSqe19QC/xInHRqboAwcncisCZeJepb0OPQ5A+WbpTM
BPXQyEJmeK84AK/+jwepJ9zAW+drIyVbIVQY5PP1f8vmJIxIWDKnuwt2jErXi4BKktrUOhQ2Rhjp
6Vszw7A+JMTaVHTH6gz+nqDCte0LPLz3PGQqJrXKlbotQrglZsMPlw5TL925SRsNsJCnktYrGyFZ
OXrR5FYgt3Ro4f1NYRJjRV2mhgeg4krov4sT1gLeCeiXDvrThTuwv84aoSgJQHBLkrGEEjR6rC3d
zvr0EsCG06MnHczVeUb2OFlSWt6C2jcRoEoEUUcMbW7QdfVaM8z+Vt/rodMVEURELGWlTnrnQ7VU
Y9dFw+X4fDcQSCSeaF8MdX7ip8q/B6mnMfBaE5gDywpZVkj4Bx1Oc+sBEe8yq3EannoPHWHqwaoW
OWwxHP6x05FPT4FLHs3M7NCozfzWu8MSeQhVLbYAj+OORlLJLjllRYhbih2ToemH7xJSL1zZLvyy
l/6u55bbt2BvjpLhsvwqac4t4AAqBlnzOMP2lFE4s5cv5uPnflvoKfUVGcy1BHX1aQ+hw7XcFWgK
Di+M/KvrVd4CtRyenVG5kx7BACTCQe0ayrs7GOsodsX1c491tXHqwFAOJ4UtD9imszYjr040B/y5
x8K6tpCuzjw7EYsKaDACR9N8qoAgS8jmS6Pi6iL1dlyMQ+arkV3mXQOwGOM0/zmqAbYQBxBS5/VV
16ZBkKMzxa3ICz0rvM7xSsFt2D7ei+Kyl0g285hKHBAwlW9KlZ8R5PIS4yMq7+R1u2dA8RCfQhSY
mGo11iVhJfIJ8Z2YhI2JQXK43ceGsRuPKFo/SbVoYoNvNmStulwz8wYmKvbt+4KVQifm1zlwa7be
9Je3zbC5S16UEA+3xQTN9zZlNl4/fYne6EsAnDbtqUMQQXo9Fih0qzYbf7k7IOZhBy+ShbOd0QSI
Z1Bvs2Y+ZO4NeDiQk19WA28V8eBZwoOllmRfIlCjw/6EqxSCqmCeBvZbP4uvqeyjOca3X1t3X1gk
oZ/rytEgu+hWrQDAZ1goKfxnd0sD9L7VEUYj6tYZkdcLu/LwlQkbYZmBDLu4kIkSETK6TCKDjxhd
RwlWDYpv65wbKEqIsQFuIuiFlPgcMLr4cu/TPZLcgNfZ5Uy1KaeWe6VdOjB/JAT0A8aAnPOrLyny
OThXN4b9Mc2KMtLtkbl1GdS2kbsx7PGP7y7VmlUnBr65SbPly3dVVXunKPAKpAVAplsKbZ2oOKYw
wkhJtUVQvlvV+f7BRXhp05Os4Z55DT+REJNT+p71IU/ZjoBWCBVyL+YxhWi/K1ojXT8JgwopWpwI
MoewjtfUAaoCY+iXS7vUsPZTtMjQ1CXcuCbp/LWtAhguoKgflrhXy20ImN71g39H51QMzunFPGEN
wd3s29lrxcU1e2Mq357yZBEOdvMOv1GzVfXwxW1GSem+O14rWIk862GIjOGLFYRNlI2OpWw5aCBN
DH0ab7Cb+rePAsrUkkDJxOENlHr3kTEiRVonOl+v8z5R/asD8CLZq4JZEW9avps7A1b+6dVXGBXA
UEt/ILgPF7ZKaURSjt7OKnpZxNjiYJb/2UMM8Rwx/GS1Em9zQo0mxcZTeBafkNcWmMYdtSOZMQfF
bv9woVaVIuISTXtCmu3rnxVn+gv3o8JUzvp1EeNFUux3Xgx8ok/NeiycmpdHPnznhD5Un1u56Fp9
Rhx2kKQ7wxqqurZqlW7iVc9ha8ytTa0REsfkpAl/jxmTJuFSeFEtCxvAQufBXG3JCGVM3y+XpcqV
XWV8aE12yfxrPZxjU98i+KNDj1I5mXEVDmggY2EM1DeznJYpUBbijZZPmFkfeN+dkGkjxuY0GQl7
ao6gZ+UNJ/byGTQwtpv3X3Ggoc1CLGc6MTOKhPwEksO+TFHffX+ITJG0R9axuJrtPAUjQQywNQR3
rtQZb4D89z19D3GcPoGHCrlJvpdgkoRtfzrQsLahgvbJVHrjFnPQbU7BuiqgPyy/BPUztnQjYUe7
EEyxLsw6RJDQ8ZiIhiDL/xyhGccd3vGBGfbIpjQJskNCrjzRUYgzxppY6OjCBr+k1sm5toobXaEq
TIMkzKGSNW5dEWd90IIw/NWf2hB6l1QRW8yXOERmfhp8pTAnzgsLtInwQgdhYdm7FPrddbJmi6MU
28gqrAOOJVYfQNWaKwYjl8yM8tEuC+OvP2NfDEPi54VFTqaOU1uWRE1qPyUxv268LwuNxe5kFsXs
6LaswwEPrcCUd92SBl6SK/hTHDISQ2cTiT3LqOtFWv12bJgqatwFBijqPGJWpfgRbqHC7nXh0WQT
Yt6VqZ07vtqkPDZ2FlzWnzyyQGOchP10kJwPcPiizUmkxabrjSxXkRlaWsou9ykT0h+doS3Q9CH+
bVf+F5oGEiJ78qfNKF5CuHlg2jWJ3Wx5QhP90uAL0jyXJzGvaW+Pqg0dm4dbG2wBjY4X8Q3d66pt
nKlTczsLlagWeLq5mkS7rmtgb58MmXM5T5At4rFL4K6C9oyguDVnN9GW3sPssHRb5lPyb4aeytGB
cW4DtWX7CMcgu9B2q0GB9bvc20bWx64uPFNxLcE3Fc7M7/kd9DkHUXho1xoT+OH02ByrDeyUPSvw
NZLfvgqhl9zTp0Hb1XniY6DicJDNluAA+0DR0BAygdOumG0vrKk6KVkXmLqr28iydHgauOSNlf38
nz9bqKuBVHWmqVCCbYwv3vATGX4CRL0qvi7c3NGWQ+Dm/Ge+7D/h9sXqNBsOHdWhZA1RC9Ek60N5
j3lirnoLK47WDog+Bl7hERdqr8pXLFlYgm0KlD6z/7bMtH7HgRgKPfcEz6MudNLfrwjsl9W80FwP
sBObLfCgTTpd/ThpXm2sC8sqnHjPdbkAfXVL79cdeVzAstWf2+O8tlXPpbywn/U9pFN+7H7SfnOY
VDZ2zfOtLXtnN2fQJ+hCay4y3j6rsHo5VZjpMtnuxL9MM7Lbcm076OuXyMOwWVR/rabB5st00eI9
Y0FfWsh0JVQwA9zJzZECflLgpgaRAINgLUeugxlo5fSz/hCY7ohKxw+Zx3cjoSmo+PIQrIRz+YH7
oagRhCtEibW+gn+kgyMoWlNwfxVlK8knNpBPaQ1VVfMksFLkRgJ5FERQYG2LWIdj8X5oyOBkXz4k
LNkk/MA/t/fM8RjWu18hoqMTIHchgtS4ck2Za9A33CyfaPI8ReVZoN0oP13JhdMgsmg1AcDilCZe
zdK2vf1Zd12XVZG1TLLT7FEP9CuM9Jn6pJ6qxARWVTogfmfLX85L1lnEL65etlgQOk4/1iIZn4k2
qz+iO8ldthFexHLJXz5SNAwLT3AQxcOnkGBCP4FvTYBtRD7Btg0OjTjvioucfEwEEFqsGKcTO7qT
r5+9ZFGpXr/KTvh0i2UQjewYrDu8ST2BkuQ8c7X+BYfdsTEX4o+IxFP7OOqCzurZkWKoCmbwAMPP
2MESgbxVbLKLDwBlhTSjMjc/tXx9opXTVFsky3QiAaT5NcNuOzbI1lnGJJVNKv/qNSVlMo+7fexh
cS/JYtcFbVB433IsojTbTIy9nfa1laALdBvtyv8SWaRrEOzSJBhTyyOqvTCMg2e62RCtbqyOX3z9
dOfxa/1S4IOnKH1Vkk3+T4pNiziSMQdqwLyBLTYFzQb5PK2BTJL4Pc7FKumVxD8WjEbw0su+T6aH
cUhcK69vApTttLZxdUsjrdXSPX/L+DX3KrnCGLMi7whhPHE7upXB6VKkTdF93pApzJpw+fnQRPor
9fAk79Tss1YylnLQMifLpJn1P3fMfuwctPNuZiyqYKYapbUXzxDMNEaeEV4yLGWNZqYU+/T/NlJR
PFpxMDYbWn3dPumwAhMO/aHGKkDJr7yEvRI3juEuM0z5G05V3UDmCfB/8QZiBkNVToeRdVnArVyv
LDDKuE2aH987zj1RjeE0Fo+D5IhCipNd2kPlaId5TOL2PMNUTIzj1KdEwnjTMZ6xexcCSWXk/Sus
yvDAuoDss0Q+1sY/ipDLcCNyaZ+q5UrTamD6urH8vEmJ2vfFZNkWKs2IaEjgcBmr5/um7SQ8zjwa
UZNUxXl1Xe8sPUwUKpn3QvlEtvB07ukpvcqgyIW7j1wqJVxrlrEHydvDJfEhBO8oK4YHoNpTau2B
T2f7GIbgp0TiETTdLY3blkfpPTD+PG/0BCNEPWm9pZwaqwOozUiSc0qdQna8aHxMtpQFN3QLopen
jfnI77AqTAOmB4RYqviOAqyNgnDypYNMRgAu5KwEWcAC1kCG64hLcsT6vPIIpKk2WB6A8BJxHwEk
mqIfC3ThiuKwNKZkb576BbFuu2dPmPKb9zOR2UF1EmxLisahA7CGqMTbL0r933mTE13zoPRtI4Ac
PDHvmdfy6WTeAKK1e+PDMQs5j46R86ggSaElJScKhqLDF4d/vgjfN4DUCS69GsGUmXfXjZPzxJrz
nfKpSqBiIbgo2BmZH3s2a+StTgcTjqcJs8TWf5P5oeb4jXkbujU/aEYbTB59gFdhn4M6lcgrrC1N
hhtwkyivykdUyKFz0cMUZUrfVLM2UvMClWENhQBjtdXrtMAM7XbEnA1Ke1ruT4o2gcMfIYr+FROz
+Bi4V/0iAflwqEUXr9v6UnRLp+uRvkHC2shqXnPuZVKXv8fixPG4WXTWECxdz7qyYlKr3/+abwJb
RqaRAJsYzX9Z8mlSXcSufeGTt04gLwL9vuSAT4ytagqSP0Kn6qQm/2O4sewFI1/DzT4zJYlKigeN
3zmIlupf4IBnE7B9OffpnF085kG4icBlJ8BtTpMPdoXWou3TsJCqZBjAZVUVpT2rBpeBlURr0elO
XyIoe93yJ6s+bHawciGjN/p1EYDSfPuSCDU7poUcSZNz7c4Fa+SEsPsGTIIN1FA3WTBqii3hM/D5
E8gul2QhGDW3mD3WxjnDwnrs9rbI4jYfwpJyc9C+pg31iEoyAWr1vD/knNaw+VDO8W47gSiUpG/H
nT5nEZRsxDcOoOq9egH/8Emd6ptioCR/5HIccj+D5MLy4b11UefE6mVXvVmdIF6BEzIu1aX4BN21
Jo2QayS7D9XKsNA2liWhhoGEieUXcgxqXZE8/qeMWg7JJyNUPgDZ1ilDfTI89jhB7AzCvP8ACEL5
qNftjP/P20JOA4nPoPmY/kWqFL7diM8ysz4t0C8sdCamSQkDBJq1jdFHj4k7ibvKr5z0qWqyTA0Q
shlknkC7HVezYaiqK7OXxjrXv+UUxg3XW+AD4lUFdm+7AXDFGwN+KKF286PT2WlOlWOrBd5Q2Rws
ijg5FT9ojekU2P+lLWRJTOd/8binec8SLXHzMLwtgLbDKpYWO9AiNo/H2IbxcTzG0PZVUxHVr8ye
qXu9LS7jO5BpaaxGSq7fSiMP4gp+TSiP7nWjOO7GJitUu6R6RgDXMEUMNoWUOrn84PdXKD3d5JgX
Lr8svqymecAzUWBUdgzEpUj94OoZsBk/w3dpkUQPqkdlj94fdTGdFqZxaIenjEY4WRU1+brsejmU
K36JMIINKtBnmJJsMN+PPgaXzCmAiTFmZMjZemrtOw9l8gpLugv4JU8nHrH20fxF9CF+RNxCM1g3
69rBYuPkOHhEWaXIzOxwQWCh4es42hIl6SbkTyPy5ppe2j/H1pwxqPM6O5B0F0mzN3Qn0pOQ71XA
3dVVZnOghKTNcxHnvE77Bk21BAqUraJe6kzlHKKXjiNAzwZLZBOu8mlXlRMVi8bOqu6j0ezvZ7bQ
9ee3i0nb9Skq3rCcZ1eQDZ1jFAa20Wh8ck1L5EEbGWnrMROrMKOLXv+zt2Rrz56VFAwEsmTpH/xw
Gfz9pM0AbdHV2ukU0/ySVWnruJtz7dPFd0SJmM9+uuReukV5AkD5LqKc9fxl221BhRuyk464MUHX
xNBdrWu2ckiOhYaPurj9WXBvzFMjErudB35dARY3WUlo4lvODTUkSoEYIp59QVInKhDmUAY2IAyv
qTEiL566nW02CGksDcvs61Lccfq8Dv9JacJqXhXf5wcAsJKCLz9AJnbi2tvzWGcaUD4z/sVxdUIK
kE16HpIxal/bmu20tSCLitfksDq30NM9TxlgqvWeT2JMTFo4mL9f2ZU1PX8TAHaBlDg+qQiBLvA1
hl6Tf06cVmKvGyxJy72BMZFr1pV3KuFQYgCX29F+4mNrwEU9IkGBT08gIhdHlxWq+LBPJMxQOSd0
D+x4Fjr2pORyAF5ipo6GivMYE+5ieN6XYipBL0NFtfjhZIujciSUsWGD+oyddEeG1em2ToDh1YBf
llDpFA6jGvKU1BNJg7LiERqcOyPggRw9VCyLmW887uzVv5yJ7yNvJLaG7vysajSm4geSKatV9PwO
1Q8kU407HhQBzrEJVwVDPr9anhAejaUxxdgR7KAsZp++s2dFoK5h0uY0SrQrHm3VRgz9StWNi9AP
HdnY1/mr13KbIzXNMq3iq8s7aVsN9IUSDjqncU+anLEgQbaawk3qikXDSxmL0MiDqIiPtlAk3wr8
x1npuK4d7XrcFFzitSCdreoU1IbtSGduFMvJPgv1hoiJJrXX84V20qN6j75jq5BW7Qf2VATZ6Qep
kCMpapc/xE1W8JSXwg3NOmyEruhlQCFXFYM3ETKkaZ0oj/y8kQ4b++5XaMPq68YZe7aN/1T6f2hz
UjGYSYA6vePGSY03WxnnQht4DZf7BjJeyP8rWcm5XhPWzktXGycV5zAYpON9oc5jkWCIBp75RiqZ
fosYDahvQWyd1LAYEXa8umFzwafaTQiuEaCmUM+eXymWNyTe+DqrBrcMIoDGcv2UKKP/BLUCwg4H
CxXdVTTUI9fUkA2rsjOWQ8bp8m+WKODOlJecbRa8+1BrzeGj05QHE/5peD7OQPo78PgqPAhEyjXv
LcYsjlS4vfcUtRgVElIDy3gQMrauT/gLkTTve6DpNZyqwtouOWaOYWbkxEPudDelncqpPWho55Vv
u3wJL2jtmOeg2IzbSA+DkFBWNQAspvtRiqrIiJDg82UkejkQeoJVFJ7xiWCOboNiwYJUOc5xDDbG
CaaFHgrIvuIBVJbglr34H6Dp1kgyu07MiRm3rnNAGNROKL3aK4VObMtFrnqC0mRpl7HbmPftlIUb
1AdPhqNfnf0Bu4iJNd1A+psE/uTs+RTk8PwmK8YNECeDoMFtiL3eD91JlCcchkG/mgSqmUP5o3t/
ua7h+nr0vqGBKq9+P/MDFlaRdbjb7iRdiHyZojtBe7tZHbKUZMXcoG4dDgr8PWUp/pcgEWzb++An
KmhohTDHgkKVyot3vZNEfQ4XFWmJI0r1X2aQu8vNwlSYDBhULAexzyzuet3HMYJtb2mapjrjT8Q+
KtrUbP8MQfFj0g7is6mkjFgt7A5Drkwli9VmMZuWehB7LnoJa527npqYWDhUOm8/fvLht0NufGbd
GfmnMHDoNE2OGfg2ppJS6wpwQjlnnzQPmygNyR9bOGcMSgrcNe+Y+PPsPb1rhbarupc0xO1FTuEz
td1+OsztGYgtWgs570g8u8zMMDXXHvo5/Yh3VuKjwrhUTyr8Vb+vW4xa/BY9txtYS7H45TVQufzn
WM4pzBvvADGR8eA9abgqnO6X9I16pqtQpt6gmy098WpGvmnJZOz7iqAGR/zZNXTZ98IcyVIMx2oT
XkdVwaw3/qB09LT4fWYD7oxIirljeCuj16VUH+ZIfO2Jqi2jEIT+tvFj1+hTeJmj712MZOjR0gsE
XxjgT2aAhCVIkLj/8+lIdG6klqLFLhT1q7pgWYyLfaUk4LfKM6V4RLiH4bW8/LJXmg4veZzlxY7Y
RWJPmRLTVFAnB0EiR0ARuLaAOjiEKrdmNjHyNDDOp8GvFUmHswLiyDNTrcZuv8fGZ7naX8Zb2eSn
mI94LwP16FD3VwEjpfVu3XR4+/+QhEyPiyZiH2reiPcz02rwJ2K51FOxfE6mtAV5YyQXfw5Q2c88
yOJQFro3Oa62F2O2YRMl6RahoJ3lLGRLSwFm2ujNk8kcHTMeLlY2t67M7thEaU0TXZEvwPXboXEQ
mU/MJlgXWsDormwfQvx2QexcLZUouiM0OkIEOOnpNe1jO8HseS7cAkpPBCkJmuXyySCw3kNaxFdF
ibuqn88MNFC+udsE18t7wYljOowQeqvkQt9xBUIDSR2gW3athHQhDfgWD59RVAnnFti4kxzfZI7G
337hqaPxnIEDui5quxa/ARbmJs6ZI5xJqceIOZD71CI90olfSo+kPSVzKpSckb/i0f0iMYmvS9AN
xDVVNlEv2DA1Ag0OLRQo6RznN//z83/RDUSP5iAMpyJgEOHpNkmOgJwu7RZ9yqMLiTkKUjseM1zk
nhpk9zKiJ6PfF6TCdZ7ZGlXg0a0OKJyxaS987yvNAX6xFG78+ApU5r5qSqv4zct5Q9ejjsGqmSCQ
ygXjhbp9wB3OL2elkH8AgoEX7mduZ9ItyohxP6Nb3ElhMGbeIV6MmI42kltIKZLcrJhXq58zQmAX
tQAyFWapuFBcLw2HmtWnqlKO24EfGyBAaqjIySszzAnCWDmnuFnDP5fqNwoIBpb5p+7uLD0t4B4D
YQr+N/q4Do3D5m+v77vdIAlp1J8J1VZ8M7HdFyp1uIKLPrh/6NF2+QOLWKTlZET4ULVDallhQt5e
kM6DaWeAAt3WscmNc4aUo980NF4tb58Eq4pbxrJuKmJ7Afxb+AJlBUdZPm5CvS1SwkUDNpuyKTIf
CFHsbE/gDDsUYaOdDg9puam2VBoN2zpapEU/37qN8Be0FjOGkRpTNGSwZYxoNSYwNPHqVaPkFS5k
aQtawQTIUEM2oiuwWvU+JnycIzJmPxw8ZKvWcQr45HyHjjNrUqbRe7m/lklVAfr6I8ltVhUq/1m8
4Y7qOXbeKAdefs0b0t4X6FPZH3ldFMDtPJxdIlykKbpHOBdR031kAdEacwdegzMiSZH+IaeBrSR9
mgHU57Q4MTZtWUdrfR6Gd0Y5Z22VYmb6/oZ1YQVKSvEuCaagdKUJ3t5AquVeiRLWOskpmSX/g5B9
hibGxIVMcvkxofnwrMHoROwHNKDduOd39sbIC0c+XbCiporXMnd5ScoHoEqOR7zvf2Xd+ENbgS/a
UoNa0fv/cdWPJew7iBGzgHIajKDAD5ynWkZ996DVupsCQ+GaNMMvHQhAeB+XzI0u3YIzTUNIBnp7
huArywb8VnFcePl5ha7FYj2SLefcs1r2YYylZ8oPre6bVWCe77gj66fYKOQ8KTyJPf/Vbh4k1Ms0
ROsoe8Q6uNJMVofbVXEk4a3lp2kDWcCelS3wKK5D1iA+HrfjM2nF2iqJMQbw+f4KYVYAj1Mjc/Hs
yz0XgShwyEfD0gpMVATrQ+yk3tUbkIjIoDF5V6assUJDelN/j163U7dh56fv6qReZ3VWo4jA/GJW
qdchvBeF1hhOopT5ioDFgRobGHxEXuf8MoYDZLczptmicCMw83QN9uymnSl4EGBX8p8ixd7Mrozb
sbs8w2zNugVtp7gy5vYGbWNr17sX5arTOXG9LuRI+/u6LhjFzEccZLWtV+5Ms21eOfWPF/W5O50b
QfDj0I/6hiAIcJLrD9WFqZd0ZmOem09YwZAY0enPV8DTo852/IoG8M9ehOxbHfeV0lyC4Plvn5iJ
pfUTEN2TrNWRrOHxNA3nkK0R/J3/QMz21SD9sto7hjOYteeVejFNVDYuSydHoz/6O/3M1sPrpu0v
O0ajDSa3wbvRTdO25I+KAHx2q1AsXSb8W7WvQ0ARnYeulm6HTpN2LGM4k45tims0pHKHHjAObmJz
mTvI5Zs+/1NC1Olx3fKdExl6yU7pk3TiZ3lnZlXdVDfblh0tWSJfXTSnmdGdVPnlp+FR9k8ikj8M
4hiB9tVTvZil6tff8eAf6Er08P8wZ4aswH/g+j5yWjez+ee2VKFemET9md7NEH322ojlTm9tgMRZ
3Ksd0nB4VIlCaZxaxnhFfBLEw9nIg1Q3juSj/ypkYsWh3UZgnQ+QHn/+m06im1uPc4qI7CXjShkR
eEOQ5eK7fETYSvzNFBfZXB75S096ShrfUbWkkp3LSyt9ytZDFSdFU5V+d6HK9k+r12aNN0BzOiOP
PRg3SFyQ1c5DK/Bs979Y+qlJhpSHbcj1IO+zNAV8NCUh6FocGT8XhAVt4CmZxdRzNqzCm3ARkmAh
wij8BNBfqlskS4MalPskWJDJi0YoEQ3trs4OW8u/qUBdFPQKrrI/XDynyceJQQvonIx99zf4YvmD
cpYu2L8u/VlTSCcLG8BOWTthbOJXrnreiPkougJVM9Gcba7iDnCAlBzi3Fkh/Qt+Sl4uzhAp/Tz8
155k0EOjrpJf4Q6SvPecja4MvoVzkNZ90FCg45XadUL7IH7qhrYlrTS1rQlbxHUL49oOFn9SOjY6
c9SdssYud3DQ/Gq/6HaNy6rxCjKUDLws8O19Zmfgt+UXx85j6Jy3olinchfuzCiGXCTsY+UELlfw
qkv2zSIEe0sG9F2sA4B1+iBeJnA9sSRu581mpOrgqymUWW9JVpNDIHFMFmpgSYOCOhwwDfJ/9mbj
hKzgp33qWT+NMBCHNi5lN2N/qSO+kaSXTvaN55a7+/VHtxAuBe8FpEAMKswDHWjauyF73qUuoPQU
3oxVAMVJus/rvgFMHlf+/VrpbzsHYmnuy5LjB/ah1PuW7ASHUlFmVkGX/1W5ZxF0o0tG6FWqA0hM
7tIT+zZG49MEiSOzua1z1NbWkYSf2wskmoln8hyz0YmwThc/eL7vPDEmJm7GZAiFFnSFhLTymvDs
4TFot6poRFmd86SJF/UT4yRTe7SqeT2r3qpzJ+QsUZR6tjDrzieXrzRMBfdcNW4gAAb4DQ0XKjbF
LU94mEV1tKjov8gAPLdE+C3JfwiujHfEvPIYf+hz8a9laTWIPrw2g9hcifEEtRDI5WoD++UCw6E4
LOZK8d2GVYXyqJeLe6GjqXRAR41ods1X1nOu/p0AJbKPEb9+t7BbEaphx3WyBL+mEHS95w0bQHEL
MAwOFW6oDPsJ6qyrDKtSXHD58l97h2teks8PLfFQSsjLzuFjpn4irdgtmGl/nwOXTmzX5KEvmw2R
J+PStjheB95s7+Gy0ZAutBxQJax3hG7fCG8WahHhJOZsXSsK3CyNyfW5W88Av+ZqccwU6gF7nyia
7QVt3hOmwZGoGKCsL0Irb6qP2fz91gV9UnLHnmvA3GG6gUm1QRwxRwejSmV0wX1Bo8hU5OLGGmI0
jD2yVrZIZ2s/a4Wp9sN6DMsZzp7eZjeLL5e9nqLuuqY6mKHBxU1BmB0GAqRewLw9GVLR2KkqU9AU
1L1aKl8aCUsQ35QRH4+Dpu98N3qS5AczhK248xvYzzGRnyu0WrWtH/ggvRfLsNCkXCet0TVLQb4h
3W/FSc3bQduyStER2vcZNsRhAagwASRO+DRcdEGpu7Jytkv5g3tw4+IDzrVjvoUJ5uuw+x6rBqqB
CKzGCFdVWBjfttM6LkeF5IWs4+hcxMv+3Lyvm5JeHUvXpifjCngDCmD5gyBYL8hYun1InkohreQr
EODCOqljWTKUT51Ciij1YfHLTj/WY9vQ28LrYrHFNS+7CR7m3noXB5gjniAf2zwvrzvFdXlG8mWY
6WM+sicFTdaQEeeIh6BUETvylWsfFTqZPek63e3F0rVlYmLd53pflNF1edAP69p3de3GrPE8U2Pw
exhs/8PhbA+fFdW5wyMOkoF9ibiFg2PUwx8vJbmGv20PnnMxQfy0Ak/pMRa/zzamOtbHTxK+WlOK
aRmaTsBDVrA0b78crPul9lNIdZf4OfDvMcvY09XKB99QYIgVKjNfEQZX4LqyH3AanFt3W2Ys40x5
8K9jBuY/yxjYJdkMhaXbDwlFena3uQJxZ3ZkScPeKfCo2aNxWjcbtoSBvAkdS48zDOkTBQcTTnji
aaZZTgwkYAE3pwTZCLi+uYpi3sNuM2Yi/EoD14ixzMDREgRUcbhAWWSRUlwuWnRIuAhZBS6l7mfA
Bdty1XocONnI1OE14W6ncy9pQkSh2L28+S89RLnx83VXXnPNnVMOHevYyrLmEkQLwbAVDXJ4bYp3
dyJZh2btlb9J5jEPObuHlZa0FUauI23Exv9Dq6zBsJygV3+sE8R916KmKLTrBtENzy9/Ff166aQw
wt5+wVCic4/z7+W5ZGUxFEbLXZzSEMDQcTjXeAhKax7Aqw7va9Y+ZKR40bdTamJAHa2hfUTUMxJm
paclMOqwKIw9PECWT/JLX4zGLVWLaZIRZ3lujfkHMeRijgrF3teiTEz8wS4vaEQvNsOofDemF9g8
GytRM4GzRkqosc0RrRyZs7bf5KWVd7zNEb6VapSx7+1Y1dafDHpFkHG7rS7uQ8igeyzv4HDpCbUR
duncA1R7QaCSCZ8t7fPPDOZoGlVwsUGsBpup0HhCvWU6+D4Xj3Nwfi/MFKnUfDNFrF90MNRt0SS8
X+J3nMpaoSoSdPhKzi3Fvs6KR3s6s+bm8E32PWguIZamrP6JtxSUJMeZILLk/UQ2fLRJLfrW4MZl
URxyamT9VE83lf+KQiBYRTYQ1Osu1OPRWF41U3AncMQVxgsOSszYtj2lYS1pNzShGzmeGTHkWGj0
V1N1NeNVlpPZO5wW+L0oFV5wXWqY64ooPVs26VeT74YsDgmuLYbDKreiR9dLScISl3OqbnSgbWdd
Hl9ElsxKWBuf9wu/JEjylByYo9uJYruZ3RuXu+/Z72vxWQyi3ZzQrrjGdlB9zwVNp6SjNJcfuwlv
WHy7yVdkBf75vu+pSYpizZGfTC9w6AkIwuXEtEEQFOPB44tx9kBGxKVxk61R008cfTZVth/qjaH3
WnCKUKTA6UnLbgd6a2+DYHSk2p/7mkBLGftTwmNUi5SG2D9vu27ptdg3tTrDdsXmZwh3jrMFIczu
rmbpFa8Rr34x50pjbbICMLSEUBiLn74szfLZhSv4/4gc8YTkamA8r7Px+PkYCM2bEbb8YlrJKXrR
7/5t77bk72cwaJ6tPVj07T5QMrAsKG/qvcrXOFCh6WSNpy9odC7hP/cRsmgtAnmRm20w+frSA+c/
ttpF0i6Yge5vOJNEXpgXKFtHcnJ0GIEmkFN38pw4/j7bEBBjg0E2fiPGcptuM4wuz4kdNk2LICB0
4miTeeZLwKzWWpI2d9/m8doAoqzGfnm3mEzLz84tNV3eX3h6SvZyXmC/av0edEljmwcpKmMtQ+0w
s6CwLMxGOqfwlM/YNB0Jq/QfDec4+CakezRLwVwZceL9yo9bljaAnqZAsPgENv2vQGiQcA0j0o28
WFqcPeMBT41y+7y1mDdhAfC9h5mS+GQ5WHAfyn7unqabLHo7g5mxz7lcpLiabQXkR59ZDPf3+6zu
zZvVkBQQS0j32T6saYcdAb+VkRUtrV/1zbDp8Z6V2maz6QDi90iLfm3bhBCHL5RG4bVDGYYKThIo
huHDHBrK+gwpNdidfLw6n47W+1C3Or/6Ve5CDvx2T/OneHGNOEr8TDSPVACB6zDi0QoKtiDRwrHW
04vrvnOnzG1z40XvttScRjyZYzoT8zU42MRF7YvXqb2jCeX8CAIsb5D9yykMZiZG7KjeD4kooilE
AXMrQsHZp16KLgn7fkYsNapUjFrqdKjHiiPOhvOzAeazH+yTileHIAygZWCC7QcVRUvNq4ZddA8T
K6xch4NJT2zxW6DfZHCRluPK/Y1LwjLy48iUxKKBYryY0+8/BnlvLTV1i3RLELjPUQxSbqQviDD8
1NjQ4O0uIpwg2g3WTyjWyEaH0DOa+rVpITLYau62DOZ9p2W6s+MIWSj+v2j8WM0/vsve70qsU8qd
vLrIN0SwQGCvAq5hgh56wAJIa/7N3TPEQtZ96tojFGdG7n/qHBPyOhvBqVlU1po92cSyfYGdpsP1
FoMDovw2DBdb6RLg/b/LDuYIdrDynuLq7T8atFiQ5zfuDsBS5pxxRDWAOW6Jn188+PEw0WzWargJ
JUn5U7YEqc+AyzonrsCyggKaZYHa0CdE5rd0giTdMmVjYqVO6AN4IznU1MtHyncoTOIzc3rYsFGe
+7G7n3wM1e8gv9qg7vKj5SzVIsPM3eEU6uDnD0d9dY+l+G8zDSilUepyWTy0GDr+ZCeK7Gif3zee
LGWyCN1Tb3PQgvnAMidfVuOR3rsOkY6Dv7TM8canyUsm/CcQJOhFg0mrxale6wfs7rL54v2k946d
i+i90SjdjCGst6Wh49EzT7T6Up49sAqD7CrrPs2aWI6Wc/SohwIffxx95+LPjdbSfOCcbbwdoQ42
H3uwUo+V4RR8V1hBMD8RWISQCe1LvqEN+C7uHyixCQMf+jzUbMy8pNXkqbPsvBwQdxKIVYsVXOvR
K5c9MVCV40RoSIWSIT0DkxdhL6zaiqHO0dQqDE56M8hXb3cK2hw35Zr23t3fidsgaAnRe57VC0/B
ta6tWQ5qxKi9RBuqXKEuHMqinE8iO9qsflkha3+sGJ6cwecuiuO+6+fCAD/YmjHYejdiv4koeBVG
S+0QzuGPz/z8zvK9XKuJI86y8tRaoNYtum+tV8QuV9+FNllLjz/45OhpH9ypJJN9M7zH5UX2mCLk
ixukjXtEctdH+6/7q2pRUzGPQs096OaFpS4Sgl2InG2vpGhLULQo1yf0vibBRlSaWzMa6LG8BbNx
lR+qhTBeFIXWW5Icxd0KOXy5LQ4E+L3JLm9UA6dNRNN3yR8nGbm+oe4wfSm+Y/++aaMVGyS9otE9
jNzXE4bEIanK6c/JIY542yB2FYn8Vg4AjqBkfJAbKcMPQ7MpX3axVK1rEnfzyWaNLfKqETw6kDq+
mGaelVaWiCRbsbmuenIhg3SVdEx8DPzJdyAFFO7U+LLVWbhc09vXoX8jDFXeapjt7gwU3KG/NSK5
0PPRMej2U5+lXSGpS0oxK6eAXhPPwwXaFVrFTzPmUEnuXyEna3Kqomvp1s9PsF/xsWMO95h40ZkW
RjifaC8KLv0iqSKbAWA3Aa/LUlbeagTtMnfXNcXQJFNBuRSJaXx31uWTw4v7fFYuGRsI92qHQOPM
+19JqzEBkc7cZ5xXWP2MyF2VMlMgGWd4hC5Ob5CwqZ6I5BIzq4QrH6f67prMS52X7tvjXOeXCqQy
684Xk27F5LAhoTlG9Rux7rnFnEwYeIS1pZCj9rshTpa/snYEJV0jVhmRq3KudKVvzuoIYl9K/zuR
8zlegbOFQxbqIprTTn+sUUKUrKAKsgS+vLQjLHTanj+mlSCToH3eu92YBjNvT3UXjJbHBwF59ZM3
WUXQ/YoAS+A2H3gG6caq6biKTsuUwzwZGzJEosP6dRQGC7PcSc4S0ELbVq5pNmzpx3SnRDbBMjHa
J/E3z4ULGkSqJsWuI8hMh8MXktNqIUrv+9eEprQeKFKbMnc/wLAV+AYXQmPgOL6frV/3wOeh2fby
uTUrVvDPgXDJhpu9TQlQUv8Rgt7V00rvbS4FNER0P0k8TVRAlAsn/otk24zoeDCeSW2bej1okljZ
scuLZWHIX0/7nXHSq5S+s/3T2OAqc9IjrvBm03FjM2RsbMD7BjsYZmAwvlV7VW5mh5I3fBpBuFjD
AqkGDMftf3X5r43x+KIED6e1FlED2QK5eTcVFussodqi4pEtC0z4f6Lfj8eBala0i/8lCvgrzZVd
+pyVEZlHwNRW3c+VpqphTot+U8jL5lRiNj+qknHAG2/Eb3OKJJpbAR97x6WIgyWWQrvLnuD676OM
Juu2po+GbzIjB7E1iXeeDVHTsHAScXgNs0i1pdznCAyzw0RxXDhAwWP7eFW2fMn0i6QOH+fwYuMm
b87ff7V18sSgreSjcUC8wqHp5Rl8RA/QhF8UgS8ht91OZIRtCINlbriv3dJBLKhKYCFtxIOhhfqy
C3aZoGZETwQuW0kALIhYhUxG/tzJDm8VjiHPIPBOQiwnROHGX38L2HdMfTMbN7738p0sFgjLVcq/
gEn6RHgLFqAoTo0K2K6oeYNvtig6b1cJkNP0Ttx+XF84AV4bIJGUzKzyvvr+RxzLgk+vAq3U94eX
bEk6c6xCtMSY5KL+C6Q5WQNlX74idfJjuRTl0WNo+oTBmknHiTF/p5eqehRi3TJHUEVLSPtfakIX
0DsJXgt6m4nGmnUEECvZbSCje87O5UBQFi1LkLoGGfHYpvg7fUsuDhNoR+UwW2WpswLJwyVRSO2Y
Dbb5bSNFNVuU7cLcyGIJWyLfc1i4/eQQdn9EtM0iXJWV5JajF4K0J6HFpZoG1T+IUEe4m+LV6S7T
kAGnWtD+3HwF8RMy4mmBO1BsXgp9m43ZQSjPMb4C8Kn4nlymZqgZMHQKRXTH2WkX6ybgaBwhre8H
kJX6rDGDQ33D7btx+56xStLqGww+eGYEg2Izt5TG6PuP9Ax/hkPYx78J16j2XMu6w2ag7WscLTHb
S7JoHtqt+dUfpdojzawSGR3INcmzYYBNX/zMCZwMR0PJKeAuSlhdVCNgT8R0pMXd2nR6F4zr4KPL
MXTGH9HQ6nScqTeEHBZxcywRLIn3oOeZYJuV/U9CEjdw1CZ3237FABuPmHTQOGQ0pYHllku2mjLz
mZyk6HatFDestESOX3TKi6V4IjWBs7OIfWvA92l+0ykn/9VgHClpw4B4T7Y9cBiuRxEPocEsTd3B
CqtTKAnXp9BU9DVA9CUExghBTdTagcuYfY7STIv9qP9XqnXnh+5vDU5B0oK/ivpMSc3oxq+ehF7p
p5vVGRMp/JeZMX+q591Q0g3WsE/zOd9bOd3FEt62BWF9V27Pr8LnrgQZ53uF7QhAftYJ+OYoCOuZ
wQMELhfqfCBuuACIeUjeUoidAs6V/wuxXsEjI6HQ0NKlXTuXanI7ii+3/8cuWUajn2NvIKDXH6Ih
stOdp9JdIEMHbbj5067dR2CvgWv6HzTU4E+/us5DntYvasGbd73CgOw54PGrW/UjpaqzMcBbt1TE
OeiE72SE5VJLjwerO9aLgKQ7PPd/C82XkH2YtecDlZZbTpZehSBthlGjZ2zrOJ4K+m5NRFtbNErk
GIlLfEl+C44lf2guBJ05Olx06WlDrfaC+O0A4qGHffQ68HwNI6w7Zk0I7v5vsHF1SUwabHXWN6BR
C7FErKILuUrrLIX1cI8q98EyPSg+uN/ciBJwLH2YQgL5ch2U0D3P5sBOuKyG4mRteRbt6TEGUJPj
qdei201e4MoUSLIr1IRy3MfisoH1FIKGv556B+re16pQI3a2QUG8EWJSuSC5A3xsiVx72PdE7Sgh
iwNyy/ML4y1pLfqGFxPBf9LqX45lqqkT5MuP2kQHGlgfiLxG1t2ZWyVN5c+6CPyEGtKe5HtePGQc
aj1Mzavn/sxUGCvuSDLM8Fe/xy+cFjgJoiFRgsQWwWaz9HgpArwOoMUSQ5sfFLHkhnLY/slTo56u
FXRhYiqGnvJjsHoUNwh0F5UCtwbpvkJwvA6BizPJal+wzhqUvD0cDhw3zLYygeAfvP7yqXRM3Sbn
G55qJfIKOapLpwDCuNNV2S73XUNjnLVTBdgb5tyZOFn2kqIFUHN/jcaNihiQkPc8IYvRu8GqG2vW
RmsQjApEsIPbelPAMb0DJ+uYrGlnj2bF7QW9hG5kPrp06DOXcQT5l+7ZfXjuDSFEswohpe5n8o5u
yyYa2TXoVt1v995rNFAgv1zK/hEPZp8QrE+B9Y1mYHWjWJPSCUByahu2ooTiyx/koZUS908+Fuze
EchJSZpd/ub/IXLrtMM/fhEcRkwh4w85+I5eofoTjHedtqTpseR4P6/6CvLwMeaxleMVgvAQP+NA
fuCXeUgot8ZCn5VE88wqwDjXLBlqTnNDX4a9K7cuDg9/ePBRbjpw4ahdQeP0bMO9e4LISsq4M/m2
No+HTvenZvPHzWJHV3aMTcaxiuiYADcHuSw4RTlbCPEcR5/GwCx46QTQr8uXd4W0FdjmDPnZtclH
8SYUDp6d0mkJVq/s0nPcsHBqgwoPyGuuFkp0z5lYEaIg2eydk4XU8NnjQLg0KvcPGLLftRcC4KNn
AiwW117CWP+QGEECwvMKnbKtU8gjTxuoVTK6D7gJA+FNxwqwcUHMx0rtCV+vnXB1JAAnEcO5Zrr6
luojm4VKAgje4i9h4iTVQHsf7AzRGRShBl1UUsc1+0Y+Rl4bp2Y9tvHC7vp58QpcC4N07rl5nCtY
e3e83tcshoHN4hbkJd8CBgAXD5l08BcShu+hjUadb6TfElYpRL5dAUwNDc3Fs5V9Md5ujtqkWK7B
8cCe2Hbs2X+O+H+X9ElUZk/L42Wp989XbVPxl0S28CYSfdRo2vGl63i1mBHQgz8bGBtatFJ5wrT5
PpxJSmTo3FuqXLu1ON8UQuFhWZwNwH/lmaFQZKVKVoreOk25JUFeVyIpMCsbB9fb1119F8goHuxD
huOqWCFPiIN7htj56X7U6UnL+tMkwkDz3Z8B8Ea0qQXpTncqoSSRmUK9fDhHGpD3IywqrHOtNjUH
SyBOO5A/qIdbQVw6GQOz35RRqJ152nNLfYZ16WUbkyV4I/VNeUtxK7Zr7l0tDlTg1Je/TCXdEImv
EH+lkdFah0MDtgawzyIGDgOpUYT37AjxB8bmqeyhDrnSPSZExkp6phmAJr+Mz2BTnA7vX2xiO1KW
/eAK+KCAMU9ihiGUwckNmatLU9W16BQmiuRrzWHT/U1KeTAuKOmovWLK9fCja5KZ2bJZW66INTb0
gBi68MayFk81vrJSvu8E7NK7Y7o93mG8nPzl/vDyiBQ5gfIXF0ChEOZmqLF/8bHdPdilmd9gFnRZ
dte/+yqKI0yeghJ5dt5DzNUhHyMgFZnRPmUaw+R7oKjuX0ohNUTi4kHDTDsRGDR6clwip9P8n09A
sY+QWqNb9DwGjmDGRDowmrhXGNK2SqI0hjpkOMLvvILh/pFTd4kAUVbln+ysv/+QV9oCDXWEwtVy
JbQ11Z61Q+2jUCaEhxs1n6ItWSYbVX6ZCK+GPrrsBq8lsrAiKW/euwvhuE+zr9LS4pdHbh2Bxqwo
oDDaysE6Oyt/+unQln8toC9XhwIZ3r4Qli2JPCPGz8Q6h+j8aUEBsEpifNjQCduYFQrB+mswKvFe
0LRux61s5sHKTJi1/LUPDO/fu7NpEFUVdtHJbeCkHKH7UYKQxHagF1B0Vuy6XeeFnyEvwESE/z+k
ZhtQPWJtwFWoS6BbYplVMiLZ7TC+YlahfpHvjVZyC1iM//hCyAoTZiKXRTIQQHCYv3FI+s62m++9
+FgKfibZWgZY+OOgERUWkF0U/nOvQdNamp8EgwUJL21PZYrALOgOB51kaazIwuKgWs5T+ecvKtn3
Tk5//QXaUrh1cxPzK/bhtN9drDnR2ZwA1fE9RB3K2HIqbJp8gJ6zLVPfdWkH8TRKSuLr5iG6u5+q
RIcHuwpZDpyyg0UUfVUtHdCs8mSNHeyyxx/SBiumrRNaKi7gwJYvu5csZSRPsTnS+t3/dkbMJCV8
Gv3oqAjrlmrrJgCtRPJaBo0TpGbPgbtFCHsuFBBbigzEuFbLNqKJrN+1i7Emjc2qlxr/F7Xdj1vb
yFSYdhVvt+4cVAILqVYz68jHMw/9EGhFe1rEPSd0L6o5H0gef2Or5LSLbN1H9CFYfyMy2cRz4tfC
boy4xGAuJVZwusozps/h+Sv66UnX2kpiB4+6HUr2T4w0j04MtkCqL9Pq1ZepXdKmcJSvpXo+4MFd
EtW66fowr23cBCG2wuoUDCBuUHCtOVhWXxMbNq/h1DRHBKGx0HDl6Xg3dycUJd9gqxjOz8oe2mcD
FSrUtbwr2M1Vterd2ybW3jnq0StZt7NIJjJm7aO3wR2IMUuVcwqIc2msQBtnwqjUad/qldVdPArY
vTsZGaXbaHLouQxgqKu32y+INX9uoo26cQWZYV99VDDET5bSPmClEOr5csvGCDyaD2Wcz1iFXWmo
fk+EY8T3GVZWDJQ8E7KF9Mi5UMc6+uDTuKu5vx6/N/3WFXaZlpXMJTXw/mDCd9T3hhms6LsgdKOj
aPZ1kaQAB0hx8pApO/hZMoIFVAbKk/iHNDTeeVFIUKpMkZeOhnt0YFcQGJrCFQubj3UgQsLSb5wN
VFuPtRxX8dHmGILeaEr9vkyJKDRvijMaPc7PCA2nNMpTW6zKDScRtV6ulRuef2E5g5eFYAONuicJ
TP0oX73GEd+TI27VtVgp1YESZHey9pb6Wl/TrZ61JuFDKicVSTb0l7qc8MQuX1wRe4XRLrfDOxGk
as6gGYcRl3rTcoJC/ORfJ+Vn4LiclW4okUvpQhjDfVJNflgMI6/TYYG7QtTTo3MJODA6yMeqI+/N
ULwjlHMidpDOteV8OTn3fHIvF2qAJdkfAG3i7pVAD689Tfwij/4ZHuky1Kn+PXceAbOrkRP74v+6
EEolu54NiHOpLGyu9QGD1CApvRstonXVsnS+ox2OJLEnV2WimM/wi5y0eBkjjTZFRBVTruy79oWz
rlFIKTYtFWmVuTtnnamJ/jw+wIz4OKkt2mFQ26SPXjrqktcaJPlryJTxa6R6fdqGF2I1eTtdvbGe
VB/iXA+TDteg0q69x7Q53WeTpu1G+3Ub+EgrhbKCxwFdWiIT6wSn5dXJ1/tBo3yQa4k32mhLbxOo
RRpeb9mck4UsnLXXNSTcD5e9WmLsLTe+YWChcNglt3dHbjCzG8/IM2LkOHh30F70WmF6hfNVM82K
WnqEHCG6sp0Abt9/ulzxe5y3kAhkTvruJ6CWw8cPHj8TXCQOvZWysi4qRoRlVe9nS1HIZu2YsSY4
1qJEtvbatys/u17VsuuziDHyEnKZXtaRzraXLkU/pYHiwWiEa0XxmrB9DeEAe8ivW7KPnJTMHd+1
q6vReVkiDkBuxGVO1YtILrlM9O4k7EJerB5XdYhYKCb0exzJQm77/UDVWVZdId4uohwe1OVyZ5Tl
+wEQHlgpcIrmiqCe8CaFCOQthkpQw1KFPQlvS60D3cb0oeN8ghvqkWljquQK7Y4+mvsgm1kX/tta
Snx0Y046N2GfOECyYuD495X9fykbl/ZJYfoUkM2FDt1HxrcETjcq2PmZ4POLAxbEbzdDCl9WbHUc
hp7l5izdoLqw123XKL60+PmFTcCfUfqXWOPvD62wCD+18C0A9wNfU1FuIbdadBvIIqy+M6rqy90Z
jNG+4HX8NKiaRKEyHWxe2hiEI86Y8cNoZLhM1Ju0lxUpu9UsUOOCdly9ucwNFQrbuSJGCpjZ8XXD
tqFPUCxgaZHeUhbWg8m310cvYi6ZDWp6robp9e/naxBZlQjRbMbI1hAvRAw2fYtZ31IB8iJieoH3
V+FvJUCJAGJW89gbcHp8utp192KpAP93OC9y5kYoiCVNsv0ApkRudpLUZMxJ53qn66nfiE/6Ts7O
QJAEFHRgwRgzULkmSmnK3fPaZ+h08Q8qWt9TEzsW/y3DUgnKGQbW7AuvFdDy4ksZDt6rioOJ0SfU
4tebNvSV4W5OhVQ9tHs+pCTjQHwCBqFF+vka2nSBFZcteO2L/PY4J/sAEQlmOgmr4onu28kZFpxu
mis5PlqxA/Auob0AjQb2IRVICu7IGomOpTp4rY4Skxn//TAHg/JBq+XhCCZxezR9+Nsa066PURD/
8eyBxAqNaT+5fbVW3awscc484CpBWrXgTbIqMPbqD42l6oDBPyO/5OG1bSUYuGHtYebWoYjkZyJA
DF3k3PjPQCbOFQ5qxvS2j7qSJ7igjy6vPLSIhxOQpQT+4lGaNnqXEM7yr7HZGdGyxAwtU+tH/50Y
c8KWZ9dea31fvGN7KD+HZgeLhWov3oMenQrFOUI8FFMtLVVMKusrBqXTX0Fpwud/hkFWgOv335LN
6o+WUQx4ZXFJjcGyjdvXMl1tny/2K/2J+aMaS3uRxCNNtdYXbJBxLRxxlXXX6VnCg0ogYzmCXdXg
Zwdyp2Buj/OyTGTVeVFPTDfca8zdTAhdE3jTY1Qv8syIqRiUg+vn0kQZjDUOLZRCK/Jc+isRpwXm
2nn9Q2I3D6q13MwKiwmCdrQQxJd2yxc4YSPB/8YRn6qmh4MtXeIY2NB3dJytdCPV8jK/xTop05Yp
xkUPsO5dTPHbAEsiQ62duTZxXq7X9D7RHXs4iX5tciIb/4A9LS9q6/fMK67+YKEbduW7FILETwcM
tJxGdioAKZ4IoJZekIEfxmkUn0fP8oyruY4jM9f7EukEcljuY0Jjs/90lIgk9CVHqqSp4CMOvrHT
jdLqfArw/lHE37CKcCLGN2q7d6RbKmMjzz/HsczKd6qNwOse4QLyiY14u5F/lMEJ3HY+MCARtN1y
njpRorblbr3IGWJEXRePFelmxbko6MbX3A8zTHbh9EcMu1ibRul6sNJ0IH4KRQp1u1XTmOWzTUjH
3EZKaQ7mDEVUG+HR+IFGw8oRHZePpGOkZJ35RCIXkexFiDleq7Wgh5sxOzMLDRjFBN4GpIKKr0d2
Owa2udodupGhHmiaKUdS9Fht0sj3rOfTBNde2v7hNoDTx0vE7JXyrAiDfZbVIpSvnfHp6IUwARqn
9c9Z0bSD6zWrN/fQme08+iOaGWGk8WvENkEMM2C2sVEde8BF13PLYrm56vVGE9mn8w5QeDVdbN9p
hCDjVvL2RN18CxblAzc+wUooeELFM5BATNbAYrqfp4TsYJWYweg/isOblJ4v8IvRUnWXb1yjuN+v
d+R1hapSsOFNQT5oW5YhtsYuSbWmGbFdD9yx6oCYyqvUoQ0FG7lkAk2xP97VB8y8W1kdQVgXt811
o/TiM2iioH+qiM/FFPWBYAth5vSLLeXQ2aNPcqPvYcqxFWfk1IWQtL216baiEZrfYSlxUZScoYsN
L45Rn1p8eSoUgUazK4JLLijvEid36eRMcphLp7iQH9hAQVTGTEPYCouY73kP76TJOWoH2pBf+JU5
kkErXoYVS/MJAprEYwEZarr0Z/fHZCSpshBkrUHuRE3OIs9q0/03C8z3FJr2/R1l8X3Ti2l5RUYp
QaBkE2zsvHDdGdPcbRMjOde+3LGlt39Ks3+80oWO1umH/9coqCaICYBnWHspdERTMGoDKd75SlC1
06DsUO/b1pAm6qKGbdCd1atwEbgWgNjipTk17dS+z8VBtaLMziiT5rMyI/eCPhqQ65HyR+FPflQA
rGm3/Vscp76roy1AHNX9IvX5Q9tGwmn23An12JmxGSh04Tu/5qXbuStuV3xX5V7xKgUV7xcks3BK
kqOT2mo/OnRMhPLVXZvA1z+RDs/i6AhUeZ1l8cK+buutQsAboengpAiTOR8R9xVfSCqu+72ekWaC
64xQNsUJ22lRjHAOagmhTEvaol/xqD72NyelTTwVXHBOG4NVmP1FtCiqlEqvewoAa3rIy4Vbek0/
2XVhsIxtnGZizRfc6RLgvp3zjXhE/rwa/rMjIdMfpW+luU+8nZHdZ/IwEbWzHPufOljnrAkjPICU
AemIc3VmMQBGI/XYf/e2o8uTnu56w7CUxaNYokbsHffa1Wn5gAp4ZS8ZFDimDoF2rbSMcgEwq+OR
VQe7Cjq12Hh8cHGxrpIzdkb78Rzb2RCTIdPFOR2e2tmVKEPecrvC2kqFCW8vLmbm/OLJfuUAQCQV
FJ/OIBP4FOnS777y2baPSnxwrkPmVNwxii3mwcuWsakhrYgdtNisItXl6vMxks48a/xef0D6fmWo
AUauIHlrk3mCMZOwR11RwB6RRCpq3gfsoo195KNm4/N1aFbE9fSfO3u60MFx3OjiOnh1ZwAnxCh7
tNI3OSsm9vQPgscaV7JbMPXw5g86XcE5uRHjIgPI6P63M7saduqjhp2+1xSy2xBQUrcxr1uf1eco
J0jwb2gsqjMuyvMc0VRme8BqzR/yL5ZxzPkbKyLcTASjVZicEMvdSNUgFmXfuKtMUwqJbNUjm3LS
a2lOHhyOAfCKgdtgcMmqrziuZjr3Pzm2dc5EK3OY4TAHDGst0Yeo4ZWMQspKvqzEKwFoguRM2MJK
Yj8c0/qbJWuSeg2nKg4vfWOlE5WfPOGMtwPe77N59+jckHUGo/emzjJcV9ZILfWL6SlfaWQhBGk8
pTmpVWazR//s6Lto4uGaNfiWQTGlv1SBgzpyTj3hZTLk+TTdsX7w2z6jh75NHbg2YW2j0pn7gLEj
bUNhyBQulriPPW25lIXQixhaRDADUnTSHc+4uldD7bXY/Ee/4quNNbBUAdtjm1m/MKmYnrsvItub
B/3c6yU9qPMBpt9z0++zW7NW09nMvJ1fTaalyJ1UHGDE5PVboPn0901FstALsWBbmu4NGQvpGHej
PMgT0/p9eo2BKG52xygwqPWxyPoojBzBQ4SA01Mbz4nvotSsUrYOuMw5o9OEQCVo2W35y7f1cO7B
uP/667LbKG3qkKHEFfT68CpMI1XO8K8WHqpMqZmvO7peFXySjwYIqHbeEjDBeSalPYoYLbdUCLjB
4oZ7iMXvo9FplyxWH7QjINJwimfTN9WBLw62UD8Zr4FQBkG+zzK8FdfqfPmVLZ6G88g9IqSYcrrw
dDqP+avSlqZxaULjFDTAU546POKoRWZ2hio93bi+qZ+6h6+I/pFvAFusnUe9/4y+syN5dwHWG40v
iid0yZbEwNzZK/sG/5x2506+1q+SxB30GYHqHLPEXVoFI94A+BiMa7e0nIRghedsyfkO/opDteFC
ykWHI20N7/WyZDSA7B5Gi8mRM1YEmUVOKJJY9hKY7MiYdBN4cGl5JQWpEHL1QkaKzrzWe4V8JJLo
MMNDdXmmvelCszuMoKNcd2Zmzm8ncCd+4zqY+AXN8czFvHqfCT4c1++71Yxfbk7uxWn2ezFuoEBw
sjcIQRKv1MX7t9FUU0ViiYnrnpQiyoMNNGp5zveOanx5LktgNp07MD9AhzSXMVM2wQ6H1IlwC2n0
/Luy+U9ib56FJHhQQZqmi0ASGsEWZQX4tSGG2qrw/MegnmgjXwf7NpSd2ZomhdW9mtOTiN4VxRm9
wbiR+sM6l5br81Zu51ngZUopLJIzV7dEczZUG2Aqd8ibfWgZXzprTFrjCqBpTRBjRR1/8YJ89n/m
4s8Dxv4+g0MapdFKqYTm2qDOxrKp+TTAeQt9ok52iEmuGfEaRN6jxNe8WFeV1OZCerpZ0pw80XCF
HSdiLHQ9l5kGD0SdVRG2ug8hsSi9TpRl8wERWXnvm6cCeXwx/NuWi+9AAO83KPK3FokOBal747g9
JUBSik35jW78da4RLcoQ8kgDvV5/H5k80apCHB8imOdYSRdtIo4kdqESly9qO+D1Myy+xU55hTug
xEzV/wKGni50UCLgxpETEpI42Pva707EwYpFin9kLrQuEal+tOi+iuKIG9dGU1GcRyXyYMjTpMVl
eyCnZo3xU9p4yFBPJna/0lL7IZ688Fl48bMiGBdlK9/TJM7idwdwsL6BsQxnhI5fl9AgOgcoDWd8
DIXEsjTG/vjrHNhwFAM3/RnyM+rbr0hG/zqOchWrv9wnCTMi+vEfawSyc25yFWlxXmcgdbD2JR6c
DO/pTUJZ3YfT9QMYbhDJ3RAEg/3Lwwr+Y2vWozyhVvUxm1SJABB5tBQa2A8sbqe9aI+7YKZZk4f0
2B7DE3/ZkBOovVpr7MzTgMvLVmyEUte1D0mYUp9Mx0zp0QQzss3pLqL138zmXSmKo0hoB15N5TqV
kZgadt4UWbSjikpBVE1fDn1/Mc+rclsC/1B4kXCuD5nIb4win3OQrnNOcuQYX/JuZndKes4svjgL
TvTRm48SMQdj11k6gKeHR7a7l10L0bwt100RwIZ0YFlaagd5q10x9F2QnxutyyrrAY3Ksoz0iz/f
Dk8eTndPMYDe0CtWgpcBU9NulgMHyeiVHdxalqZohOBolvqi71+5/3DLCE2NzO5tOPQYFGLcpki4
2FPci9f5xA6ar1C1K5JcIaS9Vp61T4gYNbLLtDWmvkHGjB48tER0ws147M98LthVXXijqmiLkKo7
endemP4ZogMv1DsXV+w8faHse3wHoMwRNwgexUXHdVesofCV5qZdkQSe62FucZk3bJbg8TOIrg5O
XEYQcfw2vdddSHMCk4XBFVXHwiqw0zAda6axsZbw+X1h80BOc44T4NOLOtlK1o+eC18wxAbBIj+a
K/J14alLYJiPwnof8ZEkPSB2NWSK8W6Yvm2VKYK1lM8UeEzu4m4nYkZOUoZgJwjuxwe2bDY7Xv/+
X6V7AIjAJ/8QFJH3FIa9l8hazBqBUl7Obp2H6kILJkuqTAtAhEP4BX6d6HwthrroytH6SN0UxGPW
Hw/IWpfDVLrQVJq7lTGdRLO9e/5OIMsFL++Py/huPONmGuTjoVfta6vIhpxiurYN+TVD4ijVKNVr
axLPcVOkJ2DKH9WZHbUBHZRtydQo72WvcIJyeOmB8l+o7XK4FdhbeguHjT6+Epcla+jePVW5Xux7
80UPEsXxX90jYCA5ZaHomW5l4KGuPbw3UzVikGrACKfwbO2M7L4U911TZJVAefK4oa2BlwujrO6d
NtTGluhpIcTn9dhWkzqJjsz0fRM6zUk7MfjUSFikdbyC+lmeeESsxGeFAy3H1vciuniwomAjcfDI
FQq3HtXI0Nkp1f0xnziaT1ucxxG0s9ssE/8I/V2nRVYaGNQg2C05SVJyIJw+/cNlav0sy3Kzhkgn
HURTOSdsicQWGleLAmJKhtt5qmMfLaGtt9XJ0ibU7JcO7YwHG3Whhj+xkhBVs/DVJeHASL6sPXdj
GKW4B97rYhtIlW2VxkLLxQni9D/fRXM9Gz2XdHaHMFBxyjWzlbMjICXuKLWYfQHh2tXnoSonFSbz
gkYQMZJN1/PQG0lQVS6aOqQmo2liHPcEc3wWlJp9FeSqymrCBcKmpNhifvADbiaTUjTcUjIXRmCo
AO3AQyraFf3SLvzMXenOmnSPaBuFd+9FjF6omkmW/xf43PNn747AL50eg1+idGLWqzYv4S+Pjsuc
db2nBorw7aLFJSd11aJS5vSFOBakEkMcrIgQdfjRX+TWaH36sSLZE9wEIGP+yDZFpZmxqMnaJjJP
XlP17Pvjtop/5vhgafoUs9JnSXsvOlpaJanUtG9QtWW6niUrWbRI5nffhU9iwlYAb/CsS5L3sodx
XlsiimqSv2/TTM6z/guqRQvgzSwwN5j7Dq/E0treaadzM6pRem2yi8IhopAZKB9fFlN+DG94SYeO
/eJNtAwF5AulNrOIUJ26YeIAcmCGVP6bQVELt7cyy7JQOlMoDa+FeD0LVPyK1l+Jk3u/q0T32P6a
vI5WLXgbXCFYLKL1/3PBfSPrZw+sn0+RvfZBKPRNjrxAl13xs/MraNOJJ9JeEhQMP67ocMKbaHUR
dzsiUbStq6LZnVHbquzeHYSVuuO4Z/FZ93y+A7phv7q79aeQDDWRMoOmjXY5m0S2rn36gtG9lcmw
5JqN0/V5JZICRK6di4JAc4aQU7muNl1yoaNAG//JLJSq+5VSo6t5v3FASRfxOnbbnGHdVFQFWQBk
Lk76GuMAh5MZ7SeBIwtcraUM8TSOfy+I+PR6Q24WYkObw5DbqfgcjLzgfUZ31EXChPF1VIhIqamZ
C93AerMidQ6fQKJnjPRUXsSEEzPgo+d4r7paLxCRDuRfNqfAUiWBgDMABe8qqsoblH2RaBTctT1e
d1TWHlCsdrnKkbyanoT5did9QRFHImezkuwsndCNCjE7CijCemDAmApJRJa7BIbDqV9t5jPz2SlA
NdR+42FCsvpCDAZf1BBjCusbufMe4hDq+ZHW+TfRxZ53Sya0mV9xwpbjkz+z0Hqez/0iGJmJMgWk
p9fwbASvB9BxfYONos4hBZ+kH57rk4nIn2GgX7aAIIikYwBluIDzt9h+n7bugw4CDUhnwKYlMqNr
cwTRLg1Sr262I5deTwoe0byhbmhDbm1ghsqtFgctAWNRT8SGEKEC6Gku5WjIV7T1SqptlfMuVFNA
3jiqYclyS9X6udhEjcu4qd1k7T8js27BImQf35MOtyGPEaiBQgxBW174onVPVZ6DRaKlBHQF/d5C
O2F2CMtPbojz5lHrKMpZinQS76P8I4VnRr1KZ+Qmw+WWIFtuI3j2Qz/y8989EFOvM8fGkBXYkuEF
XZlzWe/dq2kxXk4tb/0/2W95LfvuraaYy2rj8bajkEAP53ApoBnQCxxC1313MT9vnANUumQW5AhI
NzsDJrdcKJFiExnau+bs2VaSU2fTV+zQ/B3p+1svkAqkO+e8JJ2SmCAvWTlTY9V1ZoFYDf1VD5NE
gK1fJ72dIvleZz/bYPDd+7/52nSv0N8JrRFpdnTOXC7dvUTH21Kr0hETvTiSyIOBmRR0YlscKaPM
z8yNE+bC464v06O+966luV05AWwTungx3ri5Mr3RqsAAVzm4Tm//4z5/FVD6lHhCzX6QmCvwFAji
0U3z3GQl9926yw1Vrq3St8pO5S7BGE3r8tYS1r9sOwAOb+H0wX9W9zyvZH5bDQdFRVce/X/j9gYj
+KG917YS+MRDsMHs3yt2A41nHTtV6pce0eetDN75ttBqjKK1MehmyD6ID2Wp+PpeLtysV0xR+lJB
T/HJB9nv9v4FeaOel+fRzDiRa57QkYtg7xWjo5MojuvhuatF0iSMfHxl6GIdyki1hHCic+b0OwDw
jL/V/cRQn1l28/SXidqKlqHgHMeJbC5Y3XCQ4TdEfXTS3FgXRnd0YQZF0PsUZb7pKINSW1TPFbRR
wyFzpmOphylJzflNEHRr1Clc8FiOh7L0LjJA+ZE0WyMKT0JOT7/HuZWfI5f4k8kPk2mwnC7lZY9j
xUoYx+ssNMp3QLqr+a4o7IGS3dqf3Ac6Rkvf2VuaAbET2jmTbNM0C+ccMpZc+7XpmCN8EWVESWW6
um0PZBPTp110knB8JnpcgBLBCJISh+Xv/7SE/QJJBizob8F+0Stw8BjLoisKypWuIDFkeA45xFDc
Xl6lmrsss0ZlLmKzvvjSVYJV8/Ms/CPMnszEFOpZVQ6VcDrJoVhDmbpFPzsf8rC4TtSMHLktm29X
LVqGfBxRSUmRx13VA4QEuydaWNnvP1/KQct+xQeHe8FHTzVXYg7rGKJyixLKeNrtFik3BPF90ta9
Zm5c3iUCp874z/QHirElOyvsbqErjI/BP0mr9AU38jTj0rhfKRad4Wfv28a4biqSuaakvNiTVuQK
npvQ7TwQrRVSytM70Dgom78rRgbZhX1t6scOOPkcZJZzYUBdfyyebt04GppbO8/9QNTFgqp/UL9b
BQYjEZ/NeJAca5EJGauxwcZ5i5qSAZA8pUn1gCxFacn62yF5agqk1iOoS5vQGdTpzfIWISGPVG+t
RMrwGt/AW9cgHURw/6qZ+ZYfNZB4S7g3y55qi7g909LozZfJgfjCT84AgFuZQJvuAZg6tdGd0Zzl
Kp8PL7718mGBpPIc8AyyTRUfky8wsbgywtX9oMKJruLathhV5aikoOIxA/YkUXblDbXaTtl0EyvL
e8LAF2dYL/EpWgh3L4x4xK9RVh1UVKCxnzQh/Euqj3cSna9GuOo+jZak9C9MFIHPpAnP1v8vOQxP
rQG2k8luM0rw0MlIC+tZFCjdMsqlW00BSMt45mikCBjVd1KgeBV1cuzMS9ZkjFy/lKD/jWdlgu21
9jT4qGgI+ehfy8oXfyityWf/C4P7qcmf7MPr+yjXi3Teupp0NjglPSmQKua7mMeF46uNgqbXh1v7
VrrcG3lQ+l09J6iKZUUMANBENWLnyaDSxdTtX2u8p2JRy05iAcbOEy66/6jTixgUpIjupMa2cy9n
YHDc55Y+SOe1pQP1qoTL/8z3uJ0TFjtd5WOc9/u34+80eHxNsVoCSiiqicmi1RrwLTrfmg5LL4PA
EdxZ8I7WhMVTn97+vMmTipHawcPo2uVu+nlCs6hKLwLz8oOUkdFJVtOzVzUXAhW/FYvg5vAacNCu
gY/PFttSTtPzk+hiKkC3CiA8mihiPpU34efA3S4nf6e2ssuRjGe/VMxXJc1mrTpJMf0akUciIPmy
nQhcRbhYr1Cai+g9wdM+Y9oZZ1J9A/TuL9I3SEMQUTBk61oHmQxOnAYqZNf7SXlC6d9EB3cA3HzE
TOwuzMnlqssi/eZJCkHiNJ/GXmDdp8vACJb7SpQ+EuZ3B7VAn74KnQgnKaktjHrUAsqxD4WVIS5f
AZZEOGmwvlkn7EVe89CDHehh2zGXWlIKkwU/iYJtffjhmSLcWHDgs0o9KaJYv1OVY8iWu8tCIOV6
HapVdt1fKCOrJc/IQbP5hA3GcYM/5LbXjYfbu/mCdQ2Ntxtl0ga02Ze+dTwzH9qYDU4O9OMUKzqX
N3J2My4ItRfuMxrlcHK7298oSBeRzKNnuLYAeT3s+G0tdt987yE0ClLAIGQTr5vD2pIHwqLAw3EY
jGOC+0L02I3VQkR7qTt2SX4JtpexyH998C1RC8eGq0yASXdFPr8bTPAsUwpuDE+XhnSLucYjtQIn
xQkr3XJttYf+Zd8g04W2jUAPfFfIoxvzHjhfkcluoLF0viN/p5Nd0COueDdSLkpe7EN6GsawjmZx
3I+i9Sbkat2w9sCe6j++H3ezP8nshgdAXNmTpNkQDAExlbr1LZqFyDOII8DwoE9ek1x88VF8nHTn
SL28/XdGVzFW0AQxRVc0Yn03ZSMYY3f/wOSzNKn6nTLK0isTkslz+fDS9B27V8Xc3ssfovXAiMxq
eundn3hDgtHwh7E3NA6fycfX8xfREeajuVHk1neQjHoyfvCHmeDo7jjh+RjLqBvp6qdy5lW2pnz1
A1feP91E3HIXy/4fgJX27cFeDrlJFEhOVlXINZ0l0fTlqAOLBDW1SSeGOsUMumfstQ1pXioAaSKD
un2YwoqXgI2CHXfupBTCckOCciBxmjQK2hs3UwnSl8Jc9i2jCWAOpeB6dsh+OKmdE7lR7fIeUfPU
xAqUBnOdpVPQ4EglWpkPsi2C3frDnU1Csj0HEwoObM/57TPtKAZMbgQdyIGc4CI1u+4bsB+LyV2M
UwlCF67BIvINsJMWMPJkgvqzoaPborTMcJYi2Mhwy3HJAAbE7m8ouPfSYbUbh5DSev8aedfPK7i1
KCsd9HAS375yVTwAolMdWWvSceB5wYKggZXtrbHTPANqycZgsIf6sYgxMzLL2sBLphYNXI4gtEO+
zKRq3LyjA+YrUrZg8caqueTdzYoA4bPTxj3X9RtS/Kf2sC0cudGXN+P50F7wBbJQ6uCFGRq+BBdm
bdQEQV9gzGdiA6Qnv245nMUI2LbSZdzGhrR0TP43zo9Hf3o9k/n+QUnNoV2vmnKN1EOeNp0zIz0j
qs2IFjm+ee7riIsuEq3QO3h+JHB0vjIyweHBIo2w9/htpff5Lq5OvSwuC1rqhZOpjP8YknGfIOhP
QqKryRm8ul1PnVxRvhA9mbOYEB+Y8KV5lU0is2fUOPCGg+Qg97mPy6NJJ9AY3N//jf9Lglq5vz1p
8ojcYm3f6wiq/h+c3rJOqFoHGD96Cai+I2QDG/yDT4WlBbxIoZgAs9yK8BJpLyysoPWI/gL2rJrZ
ToS2b4pxTuwSVXkx1rQR2AQ9swaNOu1nJ34OYV55C7EudRnTDqqhlTqbD+P31WtOfmeFS79uhoBn
1Op4SF6/26j/dStuforD20cG3/SYHx7N3ni/IPxcrHpXq8HmFAXz/n5x0Hi5FSPCIZz0RMkG5jPn
LZU+G9YVFxwvq9z1TLpXYAfFe2MuYSma2llo22W+Uc2Ln+i3jnOA0QpEoKsasafBPg8F6Y09+xOP
4eHPZCIV8DJOfYVOP2TwT8qIINOHF/+4WIBRcNb7H50CN0b4sIy4P6IY95z5Udk8gclnBhAOcPOp
S4YLzqTeJF1cj4JxJElotKKo9zoIPnDfFm5nXdHzLTiHdYmG9iqNa9/lo/1tD+giJBVkAA3TklHt
8kee6udx0QcIAnpmVjI/cGF6n5eI9ijK9JGzOibGt6MO12rFt+NRCrWbE9BFaWb5P7IOvbEPqDzE
b3ptY9FyIO7Sry9CMGZhm6aFOa+qD8RqFOdK4aCJu8AZWM8RBhhaakhzO+08DNl8hB5/PSOceVYl
MvCq1pfDUe3gnh4dlZDq3aXZj1K7HlVfHb52Djlw8MQpwNjWoZJ/l5GNbdVD1zPszKUIPpQEyDTO
CR+Iy90hmc69YmX8vgCIPmuGj1sKLb/JzQAjQnxzfxhEvB33Zw6Pi3UB5ZJgANOm9r6cYH8jxznj
qhKUYmhSdzcjFj7IX0mZrky/ntCBq4ndwwlMaAl23sitsXEcKWxKOfOAQ5uugLQIleJncUXJj4bh
cEEmVNgBoT/B6oi9J6Y4WlP0/KLDxQeeR8PbCv3RK2USYYxX2hcyJf87o6chb5omIHm4lpcOYYiC
MxaISsdTdk8pPhh8GNhnlZRnaEmCzwAtX6K34A0YR10AunT6YhNP+dWrypppXOgo0htRrO31Se7N
yDQWAYxrLcBZUrDI4Xi++YskLDHouPK26WYXLnes2FBhqweXz1+o2mvUirj+Mp1g5Db6KO2fcLav
q6mcvcEzWmA8xNv8Eu10CTG5NmkNll32HShVTBqmJhXlF8BxFw7njhQD3pghI1VwBUH4dJ/+8KtB
S4zs/FRfwBBjgh9QwFgTN8wwR021jsL12VUL3xvzfrlKcygnBoco9Hp0K+vpb1X58nOn+eDbFFpS
osKXR4ELnRYxNs8mfUbwclQtfYabLmTta3mZeCfhZ4COHBrPCLK+7/csxa2PCWOSFD/Wv/XILzEY
fnboPTBgHveh8mx9DKRCIBgatMalT0ASAR9riRvYmsuR+1GoLlvxM+bmdAHu1yH8m1OmyWZILoIl
F6buiHAJq0IOF5XKWQe2jm3vbVZHVdQrV0Poq6sNyvobT+XUK4WO2jcKA7m1Szb60VlObc9AeChY
RZ51y0B3hV4zsYP/8uQeBeryneO3vcSbByp796N3iwbpCxecVvVT/v8JsovwruCFJror/Rr3mI/N
Faa6FuMH5b6nSIVlFyWUMQbRn1bGq/yKeL+HMnjOjUaP02cn/xFgweu1dWEQ8epjsrLEZebaI79g
Q+KmuNB/NjQ0l+hErU9E7Q1sVlBNsoUzp2bB2bu4GW3RMfNgSOvmlub2gVlkFRjsyrwO3Ug4AvX3
m98A/8MvzLNPLOY0YaOiheOeMEr2ir6UfqeIFki/Hjiq14Ya+20hNBlvz9iWazwnWn5Rssp8AGCm
O18igOFx8KoeOrO/Lfo7dSgsuhNSGPOpnrekAajvGaVjqM3N+RYQiZUt8fcCWjyvkqv10rrjZqm7
yQC97oxZaq4KRw4I3dGucCH40Dtnnz9x9WH7+kq2cthEthSvSBdTc2HHeSwPOmHLAXUotAcG42WE
FEet99DM5A3zPLfgwSx5+1UB2TVdI/jmBJ7txk+WMy65NGF9wvymdA8K22z4WrAgyx+PR1urmrlq
f0qvtmDrSWHIpbdBGo9QYOKO+NL7LWehIynLEr2zSPUoSsAJqqSQZZBJardkoMVK5nukSQr4I3o8
q/ojzvPm1iHUnZsLXA2fScAsQ3jbySuTYgo+KRFu6kbKUo4wZHvqUagEkz0tYGRARAhpLH7eM+KE
yXFwzv3gjAPe3+VTChFbrM3JYSalv8zSpwGe22YcYOOdC8m+IgGL4SHBqNL0MqnqkQIYHKnuNdza
8VgGTtVgPpzsdAaNjyfzMpGwj78FPGUPFm9nvZf79/PhW7ozjaB5bj2TFfi+QSEjUWS/GCCmlZrW
kTFKSF+mhry3C20lgxXCYLVP026AKK+iFGuqSfJoOuwT/J7Y1wdTFfIXtwRRL2kyPeDPFZQ85UY0
FKyYTG8KvGQoGMmaK5zEvboo8jRQw7D95AsMMSmMEHjeQ0Yf3fjt2O6EpfLjQRQPPLkEgTUYDJfU
sNfUMhq2Pn4whZwm3ZNvpDAGcgYb/JEjY77dSgpq5fKDoGfewPL80TyHVPBOnNh+mtSiRCUdjpit
lAaX4qeK4rAmw1iHD4Qh7sg15X294ZU5TSYJlPAoEdqAvQJgOqVtBXGZjhf93649id33qTnE8vMN
sIFA4p3lIdBkyFEgTKBlHqioolC6LoAQNO7OelvgMdVPsJyiU8CR2faIJdumkpP6hmzjfezwllGR
zl7N03iCkcGe0EDo8hMx3Kl8ZK2ZtllTyawGfohrfo35IamLrgld+wXtR/DEBVkRTbiIUKy2izn8
0RN8yj4vLK/+eWU420omTs3zZolOljT4meM5CuSeAzT/Jp7eDVSYZzsarP6VrVOAxMktuz+uheca
Rh3PPxNZQX8gK+MypIAiaKczW9Z1t7uTIKqXb3huZkvUGnWn7YXLJBiIdAOPy1GMViiRYwd8/Bv6
48ZcCUpsF1M5YZiKSCuv/txBg8PgaddVgf1NfIpvZ+cha497173I1lCnANoIfzoWB9aWtOMOQFXL
1irnByT4nEFfBazBm8ahyvr52WZBgBXwNvB3jwu7UNUI7Q1OBAZVHuzfuq0pPuBkUq11Q2//rL3S
mtfT/67f/Fp1QdnZ+07iN1r2dvw4GU00ZuEfLTGp3KvmK+Q8sFUvwZahvusnam+XJHAVRNQaATX9
DhzrjdwivQRh+Q3hce+txL180CanLj6dI8PSX8myHmZKzIMjVBJpKSaKv0PCSGKl3LfKGOr6/IJ3
oQz95Zs2On7sEWQCdStZiZjWIBFQPy2OqDTyUjiYUXIMGYfPyTsMRo/50IGK66sKXefI1EuYFnFP
QKF2sJFDV44Mgu7QpDlzROCpmYd7nYVdMbSsQBjS31Wi/31HjqoJkLg5L4XgItW4LY6TO5/0dm1T
whiJRmXwLKdQozw66WiBxa/tWX4V1yl3J76BS0RSoJd63i6B/hJpNL8GneMVsohk2DYsu+0MN2YJ
2nkT624MznKfMBy3hw3lkosPY+nPWrcl42T7Nzsa7rhAcO38GFSqZ4RtoorOL/RQg3w6jT8XHYcf
xBh7yDRwVMBBBxuoCC2HVf/zFFsfbqhR441jjTr4lPXo7IZVB0gwtFd+gm89I6m1P+u2F0ktLNnc
Q22b8lDMGk6O1hR4DPzPrUw/lx9WoPuGN8y/3TMN3cyWXvkc+XlyyOGUse1ETxcHrFQ57Q3DfxNN
hGM1/1EFne8kSw/F/cJ4lEIY9eaRQmQI9qwC0oAQdVUG8MD7b6UlGjojrW907hlgFJ7QH5WkK0iM
HPDkxVTCx066Z4B6O+GQOwo3pMPCIRxynRewdTLCGbRIXMd/lCcEeicHZpOMr9F3eifXu+C/WEQa
P1OGb2OfFWk+tCQJYLJViSrUjgU9wtlqMDpQzVwvd9KA2Um6t/mMcOGUevRV1LzYHcS7T+V8qglv
6tPeALgctLTj1Z2PFvirpx6karvF/ScmANuIwp6Og56HS9xJWv6QKbcWrmy4k4w45dm24N+Ap7fJ
7uVaCvYHWdp+O60nJ9Eb8795EWIdw/S5Lq69Ohtx2sLAVg7YgFmIbspgdRcE5xsEwQABmYrjBU8f
chXs8peb0oqcZERTRs8gqJzyhdYnlXkDExpGS1QzfCvcbo4QeewRsglfI5JtyW65AKoxfUKo4OWX
5rw/8PqX4KDgSeF7osIfAP97g8yn8+TfrRyqVu8yGCJ9hFr3SuIWZkLE2sjQmMchorr5EqDEjRbR
hWKZiUf+eAkqQO9Ewbgg56KDEWRiD7f+twhoPdLlFgqrShHnnim6Ms90zb2aNb2cUFFapNjmPBOM
vnI+m6Ho3OiR2C6kVCgggNilSnhXSqFgsrV67bvvzIdUONbByYQYQJ/8IgCh678vMTPzjN0vvhYd
Kgez4dLUlm3OdVllfmn10GutP6ObHTNRPyktufpO+Ti/KhUb3LGjdHhKqU1p++92YTO6xckwjMdN
GkMN/97i4ZnFGY2ZgZ+Ey5nRMVLcTttOZjoc/BAlxa5JCiwyJ+QpVg9Nn8BjI5dvBbjW3WdBC3x7
WOJM0JEq+D5aYmKCxxHXrGZsVhVAOKuAyKSpOaKwn5KIGvApecOGTSXTcyF3/sIRS6y8uCyUh5oF
76VpNzJ337uV8o2LnAVTUxAZCECtQylCJdkNkWBpKDnPB4cw3ODBPKGuNBvTUFEMungzGxcLEX9d
7ERXpmXTBh5GkP1LRnd0C3zU++/S/0xWSEzmMuMfL+pqRYtFmU/95EuKoOpQjtlvtY2r4m1o/Jia
w3EMsRHCDtAwBsQrcgxo7MLXWlq/TP9gT0C+17WxiDFCk1QQ1xVd3uHSXNSg9LUkslDWrrlNuzX6
npoMFK4/xHSYPc+iBYd+p7AUuWQXopxPZCUU3Qh7H0h7aYUELNeicC7dGfc6NIMpevHCxc1S0gTs
/MhFZxVCSGUFAd2uz5hGe5MCHCAs076aw6fXEIuj4n1aur4FJKyyE2EPBQhDAA1QTisCGNhwzbVz
gUzM6cMECc1AisgmDBHQ299x6jmriE8xGrvULDzZ2adLuTF58M8tPidVWSI77PWAH3nNw1cwWyEr
OXFQxQ4piMX0d1cdY+54s1vvC6CYzL6lcHWUAv22fkjI40SbfK9Wd9zSp6OnXbEOPr1Ge7NOXGwq
CVwAhd53JK54rg66/EtpAABbgEFe9u+402XtR1XDoHQjp+ceZ2d3Fp3jCr+wNN3suwRe0VTEqn2T
xTS/HCfjsYBE/3XA6O5gK/zchpQDXt8nIc/jz9hZZF34M+q8Zz0r6rJETLi7jqdtoL1TpFk2Gvkl
XcyjFDWKQzOiAKSX/Md76Zt4uulpjqdJOZ2nQ1SJa8OVbx5uQIM7FvD/4/GHxZVFaca7Na6oOYxT
OvKwZ4gGuAjd7byirkFOmlKu3dqDzs77L/PfOgrX4LXrQEXtee15rtlSjacoaFBsoBMxvbtKCaea
3tqhdHNEDZ+X51Bf4SHBq+cZ5gLz4Qv0A6dWAhpl5MOTjHlB/zmBTF9K06Q3tcL51/3fD1zumkcB
4+RUsSKuhsa1LOH3znSUOP1PTFkyX9BnWdCLfyLDavuQ+5+qvB08qk6+15ufMM7RVF9S/M9WynK5
+Qt3gduOgPRWALTq8J+4v6PW0HAApW1qb0aYQ7W3j2ov/ODaZwXd1SsMCFP/GvPiNqIKUNs/F29i
se48ru1+aML+mWFulg0MhFD2q11CFbrz7jxV8bwE/8Ubq90AtDgW5wGnRf7kNlMrdL8GIHFvFL1Q
BVGam0Cw6vUxb+1MH7L3/d5EGfdfy1JMF1eMpPinfU3LcSs3n9z7m8pClpQBjq1QRCAEoZaehs7J
wyCp9MMuDS3xy3pixjOSoU3tpuLBsr4UeYQSDW58YAi5U2VueczAKRSgcVdWeGVe9ytTBoDu70Th
mICVLNBEnFej3ZjyzNFJiD5UlH8Z8ldR46IPh8C10BlsjlNkm/3O5fYcqdbyCs6k74KS4v3UWZ//
dk1hmXGFYn1e8Fu5mDBUL33DIRIPQrZ2bdXPKZcwCpMeoGWbmbdMWskKafZdiVSBqdlKnD/iY8/6
6sZcXcPiP8AgpqB2O9QtU76WV/HAMAD1SrYfsQgn2P2TX67K8SbpYig+gM5K7e/kjjG6yBjEHywI
PWofgnOYtKs7Ktq2ktN/TGMhLUT2Hbl6wg/WsNVBPTd/rd1oZ5RY/O9ip28ZS0XRpS6zqlqTXm6O
LXduUjXWEoVb03BPAr48r3pTpLOtDX+vDyxG6salUFOckxpLNs4ONRumPfCPR1/aIbzdioARgIKy
q9JQWCnuCTyD9IhyKyhYwbDVeKmp9Sr63QysS4oKqU6I+m4xi5jzfesh3506RK5zr62G1I3NnIcb
1l97n3L4Sbtf7xtuOlcGf2HQF/KKGysCiodNQ+4fMLepdxYqHUiw+CXdOm0naiXS4p2RmP68abAd
uwyzMKmx36oZIHQMqPra9mMGcftyLtK39yqPE2liqlzIxNQTx08s3EiHRJwHtbSlYwzfmafQtayP
bYAUTscDEVUdgbG6EtfJrbN/6lCww1aXWGl9l1CT+uTrhsvzjvFaCxTiibNwGYqcIS1zRCIkFNo9
TKDMGYe7lpO2ysIuVzjK1uUtT/dS35sh5G94igdblgA7DR0AP/YChVwT/RkqUS6yXEvC4IeU8UOi
Y2LuX1E0z9VekTvsBojbVzdqYc5KtMWCuv/MEHZoO2V2UNXj9C8vxSnN7vcKFLMbmqMS5c76kDT2
kjoqk/vg6Q31ymZuJVVcXXwxUAowd//D7qBlGVRBgLFr/XlKiSThqNl+iztyG7HNCC0r5xMbF174
K2NjcyxjAo0cbrrOUk8p8pSkEeMPcudnEX4zBFfTXJZCGdkfsvTXLPoDHBw1fkekK5zYPPCqS1TI
jeugFHChkck9EDU7NP6/1X3n3KP9Qivx/VTIqwKF9vHrDdTOzy25cye/SeqVt2TFwTf2x+U2S77r
BrUyXl8lY4+KLT3aMFy98QlgJxNvIq937s+/4Ix3XesYdA24HRpByvhYO9KpPsI22uyPy+5V8fmQ
yvqml5ABqLw4dqliN6tcNIBWat2CU284GHJbKlvAijSoaPoF7aeQN/u0kAPoCIJA9DlFpd5rXiir
acc4RWprLNJ/eu2pGGFn/x8c5r9/FS1vaxz3RweHqSBHd/MchC3VZgdQ5OC6yde4cZckrgYXXNOS
08/I+0k8dkUpLAziXxVt/Rl0sw+fPJb47g2x5d1X0U9ZNt33ib+YO2nbLpwDVSjvSYOqlYjdtUtJ
k0QQ36C97zRVx9xFfE8uSYGHq60fa4G2YlklV3F6JUUEgzQticXO6N9rBGij1qVIduXwjKe7HUDg
j/vqlM6AJu1ANpdK7loAlEELa7F91dfHsbeIKSqNSvuOBDCt/IvQcXa2hWwf43B0KabWDvXABZg5
uuJ/sI39qnS8D/NOh2dQSgy6cXpGrhRDHF/uS+O4zDWU6avrKNF6dB/VGTbqF4EmyIjQqukg0bkT
XFB8Hvk2kyndMZpHagIIdlRWJ3bK2JCBshxans4p5pCe0vBCW3Q9fgTNLySubrS8PsbcFyptFnNP
4lCuVzFniZJorYIP1IsmEtJSdC7ZKKxBVW4wbFDY0P7f73F3+ipZSIEOhLOmxvEbyK19+NuWg3Sy
qdXv2T2+KBUag4COzq1A+zf5SrNmYGvL/60B7tE02SP3GIUNnTquyJNEUAYbJWrvMBFQKK6lsVNQ
cs8VPPwDTHRsPmmk5Z983oiChJwkuwZL28e7VRGPL00eS5BnMhcI8+ip4BADf3y/SwR+kVdV8Y92
FfvmKwNmhu7Hl2OGUILEI57Bz/9lEVJJtDGw6ajAn445ARZcxospjTG9d5Han7W8PBiGQyQMvalH
nPSxVNTzgxB2JI5acIhpUzfBgaGVH3CalaOqOwm9niSTzXKIj2U79Nay/l83Dfervkote2Zc832+
dzNTMYc+rnleslLY84SN7MRaJCf080B+IjnkEAZ9dF/WKKdz5BrMywhM41kqRzRe4OgRLa3jv5b5
3S/xXUfsY4jvzCP2tzUMpxrvhsfOwgx2pofntSnw9dVGM0kFNgdvgb6sOf1mEahq7dBt9BNUUU/Q
ssnRHuZuKBUFbsOHtlNRtFbXeTBXvC+VeIdceLVhn7aMRiiGxs6bR+2Oki08AEOtJ9mH3MoMhypV
VkNj6Y24eDqqTLb9XHnb4CW7DbqP9E0bDN5aaPcGNPTzxOL8R6YWlhHBbKoAHiIwzH1iffK0dl8q
g1vHPgIpOAJtLOgRkLpyJ/UghcY0JiBR1moiLzfO8PgaFciCUuZrDRGYPeoJ75L7ve14UAsHltPU
0uJfgSO+GK7IwQ0yxx6jIY3rFIgsyekdI0CJVfV9nhJ1FRI2ZBKv8vhyBuFYk/S4nuZMffFECo+V
OQxAUthTOITZb6F6do7UXbyaP7dCp3sIFvMdrwbBOlIT4Wa7N8agYqkCzmqesHRUsM+gQdSIVPNh
5+syWcj08BbeCHQKZkcS7ndHr7iArvKlixmvrHLeExoNIXYocKig4JJXgEDeE+Krv9GQ4wByYzX/
Mr6VUTG9AC7tojTxA7rSqk6QjQxHXi9l+OV7/BbBuBSHQjOCwSCz95XHmKe2ktuBVHj2JAT8HEJL
NPGOSQ1PiCCb0EwyUnHtrdnNkE4b+ETWfQaHuVYQZrK/U+FWNj7gfWuaqbHNgTRDKEx+q1SxIEqZ
fp97rU8xDxBqR6mFCHvhGogRphGGNPnrWwl2cIE6F7CqZI7ISQwGBuxgnVGV3VwbMXtZZqqz6Wbl
n/g/44MajADOUSxd6SDoubTAhHJ5fgB5xZcaPxo0Ag0gJqrjYdGAVEKuqMm7QKZXgme03pxKvh6F
hmUBo1vU0B90LLpJ82MJbDH0BLPp6N4bNZ/t62EOSCCko0VzMOwGpMJKCw/NJDVXW1NwVJ/j3fNv
VriaJeuSGk5eQbrdv/5QmK5iOl7atPP1TUYNG/gZ+kX0kn9ks6prU4JCqcXerM8P0RKfgNjxXAXm
eTriybpeBIfVg2v/5nBsRjQReZ099yL29l1BdNi4rxC5anzWrQw0Pj3YUY9v290dUJ0/m2fndBej
vrgYKEdtTnR9xY1pGjLn13USQQgGHa53QKDuTm2S/mpMOFaFzJxrBnlgpj2+ouAFDs/qrva8lC/K
NV+1JKPQZ606T6N+IiZvHs5Mdkr4I8acpBVKDyNqpNEkV8pIVnahfTaAF/YVwrFrZLrmQPfjZZDg
A6Su2FEDr7tnRidwlSwe4gcHLPUlMDF03rqYumjl2glhPFbndGJOGhIILPneTGyCesXKnl4hlnMq
cZKPs/DMjT0cs8BgGnPe3HlB0zQ1GAnwBvTNCA6xeZn6ckLreyj5PniUy2R1tjRhemcpD9tMBtE2
nXtFgvqx6IRLpSRZfJSP7K8nu9aXIW8Qlzai+a4wAfZghZZwD2qozfw60+byApYQrwaKlQ22UmUK
zRqapJ+Vk73gYtGvQ8yGuRmXeZl1p4Z2keCB6NYAeKKSFyNISyuYj0CGQOx1Bkqe++XQhhxpIYYn
+5SKxKJXGTVOQ9vNaH4QOFZmt9qdLBm6XyBEsu1KEMPg5V+SMefNthg4lskgsvvmrLyO3WREX8l/
XgUl71Ed0l7tF3ZM7DfZvCbGjitc+JW5PeqSt4UjuKzxX65AeTm0BzMpw2+J6is+WQzevjQ1PCwp
q/VNLcbbyzjsOT6OdcjoVGhzHRYYNJQ6zJIzn32ERN4+mnDF/eGUF8XPdb5Hbio0DmaLMJhPIlGi
vvd86DBPJnHcJ5ZosqVUZgXO0SGAvTOuiq8zbjDH74abCsg7kCKc7OizW4IijjlpZqShXp6bju8F
ENwzho3rqXkd0fLpWa6thJMYfaRo0RuIQRrI+30kjx+BSWo2bLcLzb+Kr1WG1aEaxFroXsxBZHJd
2iANh65qJW65M4PtnJdQEpgLJAiLoOQepzwu4aj9I203t5ZVe1CTIsUV0vUauQkLy00P/jNF3v98
U9GV72jspBVhqszay6hGvDVL2b6JdoED9JDSmB0cetA0wJ5QL7GaB3n5TCSfcqd7ELzRN7Nug4NC
nwd3P1/u/qUbio0TEEt97siRcEazrwsDZkd8b7LYD29kz9ntFsM/eDctKI3wyetDHECDC5MqzSSg
OCfRDHhbxM4OOWjfMd8GB0VMfsBJdhcp6RIOwQYiY9DTiT0xN4evmWUnc2JMzTR4Weu0TLojzpE+
JW2We5wUAtRNAmOf/GmgiVRjfUmmoS2nixLxyhFlMUvMxES2ZUzreZjOs0Yf26n9+LKYoCN+3RRm
KwCTefnGxJf6WWzY9XAY30Pv20ibSk+6FmB5n/JLbZiADjZdoTvtsPY0tGV8xLxuvVrhJH17/Kxb
mqMEILyzw/nzHKlUOF6HLFJJozKpVkhP6T2IBUnPOFpq17aWwRCuYWvLvlstZpROAHmSCoQGnWQ3
j+FMYVfE3AsIwSP/slLLEj7Lre+GwTvwXqFbPoX1dAglsVn+AlPtJHvLJPDd6/uzsF5WkzP12+Y7
A7qWSaYKjUrDeHIJDwKZFGudP4OVR/N523V12AyCSSEcqbwq2+lgeDJw12HNeNHr1h4mRujNp0cu
MHT3m8zr5Zy3oJNDvx1m/8GmbDGTIl7Ud/NAfszFu2fQEmhAxzrM70e1m8xdpYpW00lX7Hw8ApvY
EVbqp+jK82eQxMbqU1xoRiSFl7GX+aKyF0YGpXOAXvaiBSz2V7OMEd5M45+vLMoRBWsFZNihFCJN
/5E/pUmG/ASHW27AzBOtexcDpbezGZOOIVNrOqME2BQgrdMsopqlfHrAnxjlZmN2o0iBDP7nrZSB
crMh9d5t75zXIne2fNa3IzDZMSowQKU5lyS3QWXe7C573HevxQZvhdcHZfdleOY2ksJ356ZVPbsd
oXmm9pZZGhj6+IUe/Q2cOBXx0vTu+tnVfho+i4e4dKn4biXqz5nWlhk2EeKXjPFSkyIazl594Lgv
ZHIGhUggOv6QObZPNEvd4bq3bWPYtXiWWHs0Sf9WnTP8UD1c5kfum2LGmieDFcQZZYapg1RNhWY/
S0S6FWOSNZCji2AsOs8gER1pPxAgZ2xcP5rTO9fTRbq+nRcqUxNdtsv1dFzH6L1gjhZFpn5gGT4O
Bbd1YldvJa+FLWuujUghJ00SjUe106BdKuyrevb6lbxAFuisZpp3/t6SHiSYVGIgpaPWlSTB7MCX
lthJBe13M17SS+xF4DJ5Ty0ViUG08WauSNB2sy4P86QsXTl1l80rvChWH1qC/trMILBLw4N/3ye6
f2f8mvPN6b+dh52cTYt9lEdrl4QTTpFAt8pdz31TwdrxtS7XCaGGa+yCtPHo+TjJmlN7lEqBpcnA
QbcBOIlEQGj/BkV6lNsXViMdlEG/o56Jk7RpttMxYRqS2c5PQ/U7bTvSuRrA5E5SmOVCEilaeu0V
3kOiHtk/AFpSiQGn2pIUkfaRoYCrvH+2rSLWACkF+kEV9KDwP2xy9mwI/l/zl83wk4+Lrb1fBWa2
XwQ4lzJbt6cGW6tja9tDt720q1pRcjqwrdQXsU/ppxZr73Zv9joFkbY5JhDItAI4IJd+ZDqneteQ
cCuFAXo7H8BhPOQYxiYpnD8fsj2L03gkKt9n1Y7/K90WBDC3F1+EmADVw3FbjynEUCLP1/BjfMj9
TyTTYyVydBBVYTzdKSYVFumyyez7hM1HGZvXvQu32tKBciP+1GGukL3G04PxSs9IXDSkw1wxxwqw
QwylkYZPd7aNEOHuk066K17ijkbp8g9NnPD18O5zWTRS+XFl/JVAqdC0S1T4FlI7t3RtNd/XEDN1
IASL2+6ERchL2GutJCAha9YNgSjGBXIsU7NMhQOSUoBQS5Lb7rJAfTJexiv+MN5XNbuTcre9aDMv
/yolqgorb4alt6N70xH/u+Q07yx61K5MyGshL323f8Zh1gC5c+txelwayt2KNA156J8OCcaV4s4z
bgVGMiRkGbg29SKxdkXHJZDhB3FoH/DLzjliMLRNY9rnBE1YbzZwGMJm0Ys2/4nlQ9PdZCjbvPTK
6g8ONNCwoDStc4GHc+E5rP37AOm1kc7h4tn19gs6sGBgx16nqEKEjVFlcluAaYwUAsP6fN0q8TzE
M9amKKzqzzMsVNZPJABBGDihpO8GpMADHTRTlX0z+8NBrjWR2Mv7ZlQHb9Q7fx2KnyTWhYnWWZB6
UCU8bNggCD7CE4PtlcOqYNokZppW4pVI/BjC9GkVh+t64gIs09sz1lxBBZ4I6WfDj6STz8rIMbu5
7ttWxkMwGuwnPY2Vdy5L+veWFt9BsvNuRtJKa8rgHTecETLFDsGNIPuWvgR1c/8z7vRBefpHmXR8
cRWaJ6rVpHp7BzpK/7PCCUw66oqm/JdeuGUrfjC8fZq2cDsSwB5jxleoFVl7grOtTLXnWiE2TIqr
1VOr+gFiOmBAJQbUCWPJIJHpHntH0UToxysZ1fpUEUJ1cHmCezW7OkXN5b5ownNIS4LZz7z42ebY
eyQWeacksOrQWniCEEhLqZMSyuoEda26gYYsbxJHaSNv4FeD8t+dqRfhEu62S9Kw8C+Sx+IfQS3o
M6mLVIoUxcLmTGQ8CPtbyzMqq8p/xHJQP3VPxzVAnpGe6VDTwFfJuXACRaYgBRXA5CRuYKKeUaJl
HBuMXvHoNDVU9J76yMm+GA4AxYgp2ohxYjWjyzZgiI9Q8CLdnVZjxAUnKQFrsqXk3sMSgY3skEcA
x+ECxOjbyEyNWoXB00Yj+RHRiUlJWHOpWcplID2Z6Wu2/YIZavq/WTlG0lOvf/ZwNNDv48IhWAMQ
x8zdDRcnBslsh/3KAibAtnf6R1sXNKMizPOIuNIok87TvXGkg7Re2ikZexeV+OvIkcWFrOpyxJeX
xgLe4seqQZ3SHK9hsRKt6rl8JPDvXKpK22g13o4GfHAaRgxK8b9tfuxiAoEeyjXNlkU9nQchY6I0
CQ3QybXfwWTeCR6N/HLLqU/T4lxcg0xFpd8MMOKeu6ATjhV69ptac54wQCB4Le76fR8dQYSmTKBV
XVTqwVMugHkx90w98IFFBfC/vCfzycTui2fifdEu6gdLco0v6b+ACIAPbWVXaqBNqJfRTD0htfpu
fuXp3RA1uyYu3kWG8xNZqhEc4rjVBM44cCaG6jyCcEPeDKIsda4qt2j18zbdvR/ALyiBV+vc9BcI
rVnioetV6IHCobdrsJYj3vKkEDtNTqbFqqssNyqXIgk9VwZz1hy//h1riux9XC9eUVSUnbt3Cngz
h4BSKCFfja5KsKkVFFoLsB3VkOI8JMhejnrsXaHzJKdr8MufEurSciSkuhrRgUfJBTDuPZHtD1OZ
XCwsRsZeJzSm3/nzpBngb9/FuXLtGsoscecv+l2xkR9iWXM6MVmIjYYWgra5GWGs/xgRFdASy0uy
FBgRDhwbHbWvuv0tJtOjxz2zXdeXcsPiN05XxqOF4hSKEXoNjzMRnpyUnz+FgRwVCvtLa9qcihmQ
ktN6Ok02u6VeNK3OaR7guU89a+/8OExJrgUhXzDy7x4TmU1pEi8PnIiEzMxU9NhUS09pwfofhbEW
FIaI2caAms9ryw99IQKEyvrzyGiKdOm56LZ5BL30KfLZOE5NwD5WQ02/4TcPONdHfjMSOq1vzyKc
WJ3QQydo89OfBNnaIYOGwnqEeW4nGo4frrVfllHYGUY2u5wue2rZ61jozHqdvKuu96BitjgqpsdM
BhOdXXPLkAbkR6UOelp1zEVe/7tMZNUhhaNskk7/G0dBxQNq7U/Wgs8osdcZx2g/WrBwOqqs7PWl
sLbSEqGvpTgErNu2Ksk1PZ4qQ9VeCFCWZ2SV72+MS34WW8nI7hk+OD6An9Cm9YHodTPtDC/ZMCeI
t+GI/jAqiPCqytYVn1ucsbEAhbuOkq9WtnCoLpZGpc5VpOZ/i3m9kMLcxm6Taa1v5HIobsouPQOD
8YGaV9DtcmmafUen58ddDtGL6N9VHM4COTCNyRaN6jD3TycPxERkqZcUHvsBaiM7m95tl4WUHd8v
MJ9gBvHlW+LubP470slw4IzIws76zxDdEOszbY/+7aQN1KTVcizwFuPG5JmDhwbaFk+babCwh1RF
SUgNzoKvHs0t6Rg9GNSdSQXln2aVI/3y+8wbg6ssYYcrlO8EToWMT12Ok0hOE/ZfZamgnAs1EunE
mVg7FryLQNXGb+YaEYAdzxbdcEDYAgCTycPSihsNX6q+M9WU/RgV4EzKe+i3K76m+stk9d5kqCMk
swIGEpoAzaI7E348QuedlVth+SeOY1vvUN7Qr6FuLEDXS3qkSqih2dUq8MiddUea126vNaTnCbb9
2sovoCNR0BRlpeuOFKAu5+GhWz9XxWzFNREiUHHXunESJ2FPdNN90KmIJeuEHHVOSIMfvhIHfRPT
rHVUxI48t2A3osUbC0Stsd7gQdKItqdFeGCbq2IW8AoV6BtBsXcuo0ocjlHnb5usewC/XJbnmgbs
f9f/xHiNOeb0pOcjWwT47ixvi56WSAYgUjAkl557HowwDX1AYfUsXMhsX8VrIL4a4P+bO+ncAqnk
ncq5lFCo9Qi+9GULo8uxO746xQ4giyfE91KJL5eMkVY4clT7jQuP1P4EZe46unw73TGbYKpQDEHe
f5VgTKEnTOZ5slSFQL4LhqpVohx3K0g4gvbJjXpBGJU5sKwjYWUO7kFTGZZWNwHJyKTHlTG0Ogw8
/nVRA7guBStYlCQNznyKNVVTJ0Y+OjvXwx7RILv0eF4bWgsL3rM/eAxEUxgovg1RbsdLBTOv17rg
wQMCqFgPKoxAnM6tZEAwAYAOJZrnwZher5KOHV9TH8iAa+h4avE2Fx2D/qRmTc4ZLhuCs6IPp25z
OyYZhPPssMdy3E45mtQRLwYkT+3wk4Q0FQE7/bMShu82s9BurFnxIHPAN/TvL71oPxBF/VQeXFye
aDqPD5gO3BFxP16AvXT2a0bjV98AHYkBB9bWsUXUFfpcpiNbjWxknASXNRgdR9n1pBtOVyzTBb2a
FVlc1RattH+cuOWy4Ek7AC9Xt0oQxVWE7HKC7cl3KgGV4ZOeYYNXd4/rrDBPc2ioARc0Uc79keAQ
dERim1tgtg+mRYfqh9J6gwuIes1WDrp+l7CO6nC0xCsI59OFpHiPgb0/1oOlv7ffUzuRri42U7LR
W0y3tGMaikq4jiOkWnSP8wwhzQ+X87Mn/0B5LEa8P9lRo6vinsTT/HMPBa5bU7B8FHg0ez2enPgb
oAY47hhNp3WHKpNqffOMwQby/J0bbIkCnM4LhUqvmqq9YgEEThGdvBJn6sPaO8FbkQ8p1EQWxRSZ
Yed4R5OZwiNAuoFu/BarntwX2WgfVtYYqwyndqlp+NHwxCwAKgw7ZU+insqZiAPiSMkpNbSmmNUC
vfWhX4+8B++WTPVYmbU1A7FR1/7rHf9VcYjZYlLN5+9hJXVtHrZ++uYS4joAssRzC4mHsPUj4kbk
Hq3mN1b1MlK0qfWGC0VvEbY9ksJoluuHhZD/a4+sTBF1zNYIAcYBNWPpZG/l5jD/ThM8hNDcMZgA
WpYQzL/EqKwabhe6clmg5kmzJgehs42ZtKpkkuyPAXnP3Pbxs8Z8KE3c1O8Ua+z/w1O/EXFMuJZK
e77sHIeEYn7PZc0lycpQNDTvofCEhWN5cCJjBxrwMUtmUUkB1OqMvaMMUBH0Jpz2mbA6DURgJ5iq
gzxRcBtC0tBtv+BQ0e1XKTXLQiq5MDkRp/YmQScdbFd9AMCXz+fRGYBZWAS8jwuz51+KQKToeO5D
wOBEwRBx5xDG+kAag8IuqoNbW1ADSXBHXREkhtRRnYegh+mSe0BWb45+6fCptFxxTDcajLi3V91w
SX2VCUsXJ5bkfiIVdKio04iGg9RLcpfJZu+tC8CHub3f/Lq5uo1dQHmkKO02j6vPgTPJ+GT4ugsU
nGdRW3GsQ2ZoBkPkUKFi+QeTqr2dGEhemHfq/1/DulEGcdmy+5fSe+us533aGCtqm/qTxJ2jdLdg
VJbNPFoAkueDFbKwaR3OYLMOB2tsVhDv77UO7kuZJviwr11bwoN0/DMfPq7809dH+Msms3VT27KJ
Mf7Nnt+/A7mCBeEN11QdKVWnG6d+KWF1VceBjIR2UNpWQHjje9R2Wdkr7l501Vmue+tXjFvbsrt5
YKwT7anRTue8I/lldotn/aW9ddpG6q/OPaTedvL72FCZ9fgeYkdYKDe+clrBn5kogcjLIpZ0I4N7
IjrupwPJjxb2fmqVjIgs3nHcFsodFsF1+ATdaS+taOZ23taRlwIYUE2+gp08oFsxT1STKmDch1Az
1YRo6lWUcmF63TIUJc7rWULAbhoNdcNAN6RsntiAtTczZn9WKf8Kb3ILBWH6PdjYaXE29l72caZZ
SN/nHn1WKS8rNN6aoGazrOPMmtPcHI55TjlOlY+SuJA3dTq66TmuI1RWcQ8JQODXU7IJpwkqZyeq
h2Z6KYqe0i8X+szVzbkFREj13pxsYIQeam7KavGCl+9n+jOCzz1PwriIaBP4jFvffhDYU6tDxFxR
yhh8Le4ZtfNnuLvTQfAhVE/2bC/JE3zYsOypbmWHBaOZQaxpzl1UXBhoQkpOgJ9OFMM6Rg9t5Bd/
3wcXIgPT125bcTbanQEQQH68V6JMrletSbxk3lsCLGEpwbV97WWtTpVCYKNRbOn+5299E71rSXGn
tRtQci7i/uyvKxbzdCvDuu0Tjq76XRwY6JU0hIzYQp82DOeASaZkoSZ2xL1tvj9PdzmukMwx+g0V
LnCmqy0JNC5hVRUYNetVfQ3anAn49Q4BEdyrWxf2RLArb/x48NRsSEclqnrPQ7Uw7bXbsGoc0HCe
HDoZkPmgl2hZmu4lK2bv3sjShtgQqe09oX+XhgQibXGPNmnUusLRVx0HorYNNz8Qs049LccwOwKc
qSX8X8siQDUZRwXHwckUHHBiLpTWrK1GExgaqQqmQVaPQGx8KYSLij2GunExJOT2s+JBUtZpAWJ+
P5MXYoCPi5JBVFw5GKc/REvh4GmswmOjMBrU8rArjuunc0xzu6YhY9dip/clO0fnVDn8vee+kfwb
e/8UQmwcDj6rid0yActzFQgtg1M1tsZtZUJhT6tNN7RJWINb1XiWNbz1pUJmFeOMbihqozgkAZOM
9Mt13pbktbIJrq/zzIVldYi59E6A2YBbfmDLJOgXrDVJWfsRifQBVflxSeWqDxphP3PbwvmkdHxx
2ZbiYAzwkqtIr0p505UWpG6nd3ZVOf5owrkIfMbr4/EANLVpUB48gAokH6ovyOpkZDq2Kwt5bkki
naz0dca6g6gWgm9g+Xzr4zMNhniBMcn7IaZngUXhfYccWQU0/XQ3ACVObPktQYqUKJMFbqkKBp5v
uk3xbFWHpfVRO2/dOgahfwAd2+WRZx1yVCjJQTlr6ozfzkB5ldZsU81LXkOoH4gzYSBrInpsCqfi
Hz7qOtS3HwwdJWibfVh5F0DaMxE6DruPgBRdTz8/WGFsLYoAB86hiDFOBkt4AS+Yw53pta+rf86i
rcLjcWu5wUMBs1Ywff5iiOChvZU9aw0SYzReL/9buVK/iw7ro52J4+81wAHt4y093dIJGEr/b1YQ
KLL4DHkV5TjkPc3BpzAGruI2pcGGEbRkUNDEXn1PT8mpoTG8So+H148l9d0yVGyKLexFyI09++98
sZKiXJ62TaRzB6EZaTcpLvFKkJo/t2em1q5JE3SJGS7iWtGpVdsp6bviFJTzumgr7+Nufj/HDEw8
innav60xuxoSmvuwcQBupZFZILWzLQuVk5o5re4ee3wk1vcUntEupAL6Cwl4ALSjxK1SeM3ruhtH
AfApAOW6XXuNwFEOFu6lF0W3NSthus1NLV7dV9MvaFH9+hjbVoFCNXbs+HQRvzb+JxeNxjPLmfdT
JEhz61mee3Ow63BQBISz68llY1JviGiTJp545LQ8Xi0PGChsEx6OV8V/mVHqaMaF2ibtyIhZddD9
6Yb3gqhBOATNwfQMRnB+hEwgg53vpysQvqSXPxaChWwXhnMZDFDlQWaUuUh45cCd1wmXklysefeg
LRwd//VPSjpVjwHXZ9PP+aX8bQ4tDaCukOdlJB27t+f9thRcnFiHGpzGaYNOxFS1N/qSwdDxg3Iv
BseN4GqzLeV/JEr+FqPbJ1gaABhJpZU4zWyh4i4sq3lmQdGHMuwOvVn4v5x7fiydgG0oc4KWjwdv
O7fd4JMGFhqvEu1Z9KPl5ESza6Q/vneGuZNw/oFffYE18IgqgPL8eWc8emORctQJvN1eo5tPFjEZ
F2aSSTo2Wr1eg/8L+e2VtyQI7dIkjoP9xW22vsVjL7sVZ11v2McewUKMiUqSD/ECg89HBTn6tcd5
GWCLLy+ht5sp6mFnXBlK5R0a0iu6HmS0Jbai3Dl6FPoZ6T350vXzQzYjJ1QOnL4TtCrZ0uqZ/w5O
o1uA9JXgQcIYZyXWTzxKprS/9Z5ZUYCMtyVCS7IXU0FMXco8JI6PcceoI52m/33qilE1tvLewyXF
fMo0LNGI9vL2y66yrRN3E4VTQGwFvYJ4Cm006xqEut+NRILYwNJfmvSl5rWVMD86hd8x6Biq5+Vf
VKtVEMqxebnjLZCJsHA92IhJFLH4taBQo9KFQ6v1l4wkmE/zM2bu+RIyWOUAUqufcCa4Yz/+/pGZ
XQkumcItLPegK547miJk7SxiY2NOzEOZawHrWgo11i7zGB0aegqkzuj7pmqK9OU3adH+r2cAXpsB
wjUnCXDCfjLi8GiCn6sxCJnW8Fl0h+5PYa8aKjhdklGc9yJ8ZRtSR9pf1+GXB8HvqwPO5cLOFwTn
Z64RmEeyj7WHZxReZ3VZIjenUaQ4B09Gp5LgXYmOrZuW/oAo3oIOQ9zHj3mSNHVrpMK/hxMZ4YSZ
Gci+mmO5AJ6YeP7ZCzY9GDBaC41cPKZGPoBK/cK6ZEMWtE41dvx1sxirjJUdUkuGnVy2TxqVgfR3
Dc7hnCSf8Fl8oQboE7WRbWmniiUiYE2Y28Hchha65K/upmkfay5XFiUVyqDm93x16spl0HXM0Cry
g9UIF3apxnKj3lAeJIvtLzDr8ORKWlK+6+Ry3kdm//1rXZkgoakehdAOb75Rx5LUgqhQhw5oRDFw
tSOJSBYE7KvqXBgahDb5mWs+Zu1utni7f241OY7wPyhsH+POG1ke20HPg37CNhTb6yCKR3oYgXaA
59y/O/CMVVJW6gowoQHYr9JXkrBXDUprglybjB+BJdFf7Or9YtO+3PJuszDaTyiWR4Pn5mf19xUC
NVjoBx7RTOgDIFWSXfufCYI8SKDf85PkCCnkDV5iEarXTkBxTO/NBZFkCJR6tRzauvl/SGbKc62m
RNrsHMWqSJRE0oVruOLcpZreQ6iC7mjt2IrGzt41FaJbOrkyK9vkJPMI6pWrWeVQQA+PLj6gBpU3
Ik13liTB68dksFx9cnVWFOJOUF4p/dmHkVzx/T+a2c/AzbODs94eR7nSLgnDnT1yHmf1L4t2303H
2NbRr4cggU5HCujFVRXiKcRjL1puQ2k0bhM8Rl36AJicn68PT+hF69zGbRMmSfMQC6xDwzBME8H8
IWTPpt7rsuB7cvtDX2BmmIb2iwwWNEJ2LW+WpfuVTLOGI36dLSuGuJfI2Lf8R0wSxQ3vedu0c+SJ
5SOSmOd2RkCMac0uJ6aDM1wv6gZSHGPVgfYmuH7iHBmpWc5FBSGDe1BReV6rZxPHzhghWimvSJsX
SmoyUXFOOpEscZjeIssAyU/3+6V6uZd9GMlpYg5i0TJeJIy2JoZ1mt9FOhDQcV9VSo+D6au5+mYG
EmBrzYzj17BeKmencj3Ep6FhW2qJin4AaWz0FrQmo/XiPCdMbMK3TyTc3rX3Zf7MlEeeGo+P56al
vY/mGW4cyx70S23ixQ5oa+vxR9iM6cQ7D/T/wcmGV7KVUFu7ypSw5nmFf+wJ3vaMzXU3o63RP35O
R5Yr6LFJnEoGwYdCTCf6AybB4s0SxthrXvmOjHp7Y7rFERBc0aYrEx+H8TxUDJEzG13PoeT6K3z6
M5P/HBUi4M/x2UopmKbjsuzpc5MRe23HjfZV5J3vwWXX5U+S61kP4L3+Gnop0kZNq2BkBvBP2zrC
UK7sedBgEr0zBXbtvWny8a5865/K2gOLrCTVRzA4ulmi1Uhm/aCco833H2etj1mC+U7Iu7Et7OHb
uiLiIyP13xMh6crpK/uRBXnfAofmrzLw0qjkDo+18jSXSWrakLO8zuvomH2TViy2D5+JJOUqvwLl
SAAk7Jg/H2hsY+kMQVUUcZ+12Yscvoah1JbpXeeQC4Vs7xNSWFyozWZwrwWFIbZoTgn6I3KTVNCL
6HrYY99yhbkrN/x+02Ien40DfOt9/Za0/+RK4Fao52FXNcL/Of2ru+qRlSYGpvRvAJT+XcP0c1w6
I5zAEfl89azXtb/wwrgOLWVSYpSOgOfohFK72qG67JfacHgJM9qn+CodTajrN0Lhkuzh2eBj5UWl
xhHPXiasAdmmMmbswbXI5sbwf3FfEukQzZQJDv23D9fcd9AbS19wRz599Lduyy0WJurWrmDfRV2+
sjTZwznl7Bn1pGqr9lFtLg62TGmp11EGFDlKeQAtBIWTFJ4DZK9movGUCefkXDyo+lvltrrLzHMK
hE6VWPnbpovbv0U9RWxrKh1inDm0wy7jwAu8hq7W8HX2GAxReCmbvAnAS1yjc6qkkslm1wEVGagF
hGP5Q4bbLhdRcZNNV8dsWA0woz94P9iuj+upLHYKOJ+LrECuWMFpT6f7ZqzjzJU1TfeXJRrs0A3S
zR3KjO+GgwsHsXKcZtvJG06mCcyjz+R+MxvToSo184YOPPcDWS9433h6XnPMfT/qWaZXRpk1K5VV
w6AcW9Tcvzg3MAGq0JmWB8iz3BnuKTLL2nSybtF9LVBkOU9Og4b6jvHRUgsaQkQkbvOmbSluSuy2
jwR+z9OrVmFCAtqb7E6RgFoe25XS6/899gsSpPlQEeZGgsdMyFxraBzYm/DVisiFZoKd+gttsdyd
4uyQ8ohuY2dF1pjYoCr0wOgC/Z2vgyxIgJD2QBj962PdsrH3UKxyWecgAAYcFS1gaQsJyIAxdvp7
Dk+XQ70iWoNviV+G6xvTaqUOkjx7yLkYP7zMfLgmp5kEsmFoNUyTwnWKQpoMpJy7DstIRtwuU/RU
4aSX4B9z+6s3NrI2BGr3HSxnmvE34BfnCD2ZhL3IkJFon4bXTM4+L/4AJ038xP4OpIwWaB2zs0P/
QEYIPo4SJHdenTeFHoZ6QUeo8INgwHyhfD/nbsV3ceLqRa8yKS0vDC4qciv3IIUYOikDyWNaTSNz
TXufVWo0uIDNo9xugg1muwyNnYafKLoxgN5CEJZhI6zrw+FZ03j5wCu3B6uN/CS9g9WiTH0sNiOx
oidfDToNmKu/CqRA4eafVdMqgpMTDooYxE/X87kMo3Zb4Fyn8gweflmYY4JhMhiKwX12leOtibiX
rcwaawByVziEtkXrnWvo4s8Kzkq4c2VfOD54SFEg6HBYiQT5Y0+G1GZoTYCbtHJ5n2l60b0bdU4k
l8hxwm++Co/OkuteD5vNBtgK4MzvDWqku4AYZTDD2q+b2eJdclEFYINVHlXoV6MLVIAnBjvXO8xZ
Wm+qLeCOIwy5qUQ/SfPwcaj78oJ3mHswt8zPs88NxLFX4hVdyjKNRo3vDtx2neiihepRJf/IZoq0
Ugmpsx+45im3nRGxzpp1zEU5zHdZfNX+IFJC1W1jkU/U57AxmboKdV/GkFBZxudN8Iw2nPzKHItt
aeb4Bb+xVoCDETG9b9ZLAT+uXVkyavhYqHkT1MLhV8XNHYYJILl8uYdvCGYWFmvEY2SQbE53k4RX
w8wmZeRZsb7nntpIYKlzC6ZwqiLcO7lsW0qPNftGq+2xIf90k3I3Gs2M0grA7vm5OqALScD1LQPG
U/l6f+WmNFXPIVz4iHc/bxuQozZs6zfqHsxm6ceEYbByE+xqtIW7JrKGZVVT78KfrlyspQu+t1V6
D3VWDAVeoYshE8l3s3U/DaAY3xJwjGT3JxGm+0ZemGlpL25SXPWP+vdzS5/pNFCVHqV8Lhu1tWYo
7LCV1t1jA9vMdsnW9AYiTuJ8j7uCKfTmWmbisRKm4u68+vMJ31n2fhg+WCOgeAGzMSPXKi+8bJuz
F3bX+oS8BTy7Kes9j6gojCMCr3NZ1bQ+ZJzYH2BgWEEg1suf+Xbte0rvVImcd1iXmBktUAPKLEp/
QQkryDXZlbEGlao1rAYe5GNnl7FPP1ruHRWrlfE6L4+88RDu9sdWvS4HptraWwbaBHeJ09/3nYf0
JIlsURPMBWHqCHTMR9IBFob1/1uUMsO9RcLzJObWkIFEMyz8FsYdCX6B9Igy0owB6ggi2jCSgymQ
8LkDyJWtGErvzrzu8i2Glp2nOmNvJ6FKu+gN0lEVqQxEBHJY26222WvoVR1L8/qPQ4x+bFlnrvVB
JvAVNyM2zxWprzE2mw0vrByZQ2nk0TA3bDmC8cOZyafgfeXqa30czPKZmBtSuFEzmhNS33NOhT4M
bxZhlCnmeZgCdtc6aW9DgDgrUBUwi/0wUl9vLlWiWUXuFuQrzD5LnjomZ3ZYq1bcnpdp6QWlFnIu
D4IxnMAHxEm5mcPxXCilvb+ehm+7gYS+wEIo20xqX37RNjvJnlNSvD0dQjfihU3aKZMf7ByjBp+T
WLikAmhXqI4+k01lHoY5Ev4yLKF2hLb9/qeF/CFfJ2nOmNU4+xbujmp1DrGJr/gmCCP+FFezSvgm
2Glf3p2tciRWxdLfo+iMZ+rzAPxiwOelMkpMJEOKVb/HCHgNsvSCJ6TbXHWG0D6DFfxgSeneqE85
AGwgxnOSLviS+1v1mUK4t631ncEkn7m6ARRjFlzjNLZVm8upDqb5EB96R4f9hzavoRinjPw0I7HE
UZ1OtN1k9Ftd70w0JQrH4fqQTPeVWU9w9sPoWYehFzHPuC2b7C1WvQO6bytzXRyLgYoq2fIWs4T0
tTc3pHs6RuwTZ0rko6xI+L/i0EjyoSbYceuodGkhRGgIuW35imORB8l2lkTtyMCthOC6qVgZdcaa
+wLCmnCgbAD+hdEpiLcXRLnqVpdBDnuj8JrSFl6vQLWW1aU4kudrfC5iaCT71zLBI6DWHVUpY8xT
xpeqsfmimvHt92Mf7oCP6r+85DONE62Y/Qf1FI2ALNZ2hwH7RAPMT8FaWHieTNys0xZXl2J0G8kv
aaK4H5Wi82xK3KvSDJ0foOrsmd9kTmStoGJw+PiCThe2tHPoqrKhqquEkLVi54VM3XEZmJ2ImoLX
iyz6Sf9D/A6gfaOFIVTwmT+sTGaaUT7Wzs9IHwVRt+tqTA7YezG0v7fkLc9TxbMIZtK0h8szGEih
HoxVEXFzBpScb6meQlYDKQ/s6aiDnRmYs6WlTmQkkqAQUkCtlL8+W5/u5a0wJXxXoFOzuPY01EZt
UcvB/+rOPgU40PjGDONPPV7iSyzbiJ8KmljMMSnGw82ReoLjjSjzYnVYvsCocJ7wuERQxIeCpp0f
L62XKaBQiHydvj40hZRjCOSmgAYAD/UkOiY+YZHa0UAgRioKdULy6BO/707kSQtr0VM4bVFoi6ra
+L5lBpImTDNoD9/Gl7lKJiCto53skYEc1etCqUq8rKfZ8+k9ies0BOpeQJ3+aF5bRS2v7PHDGfvm
x9fZlGrNXAIcuCODzt0wd2MybkkzwYi7vmjRRIUedFYQj05EgjCYDGcyP1+PUxmkyB6ZAgrudY0S
i/k39uk2GxdlGwBuaOyAljLDzc3SNvz44MY455fQqpdvlwVQcx6nrRgSKbXYJ8/EOJY58YdSlWcg
WkeGnSUZZTL9tZAGisvALc77mIX1juSTIdCevlJgk+JRJ8Wt6gBEqRshTcRJ4mMpPVIfsGc5u6op
IeIxvB6m4LFWPhumKmaTDOg3gEqVHNFpO5U1IIgQMYoF3AJf5b7jNOQWrK5+TVm6sZVQMRRbkZ9p
TfpuNrZdASQv7zbK93J9XAW20AqXCbDQWC0C1OsMdlCGAUiSBfszzbuL/843F5sztnHGzlkFTo6f
alQ5wV83incBD+VNpDskP6w4ddiP83QNkbqYklD80K6kXQYHS0f6zIoCB2Zah8wwZhVX60kKfstM
FuZPkz1P69balnbX83IJ2xJ5AGN1SGJvZuu12Or4IAzpyPZ5IfZxbJk/2mu8ST79oKxg5iI8k56a
Z+Ne++U5tbm4eYz/j10oAUsPTr3pT16ABnfRujtMoXRn8jyWIbSXQbmOoi//E4f/qWVEEI+7TsL5
KAsogse3ZR8Bj8rh8M8z2eaaetTrkgUq1BlnNuSFyws5tqhcgTVND8XEWenQJZZCv6TllBwm0tvy
aSPFaYD2grJ9Sau/7mA4jbcElJDL0jrVNUN+ujAnRgzTSxEMzUcX9wb5bmNr7EOUs/BLNwbmNQoK
eS9x3vPtXiVHXMvA20A4O5uZRzFcnplWwLKsUnyd28+vCcuhq2vQxmaYmEyBV0l0Pzty8iFSkt9a
TIaUROaZ7R/jRC2r8EUGSS0uQeLcdnLsnbxxujenRT1P7NrgX+oiekQ7FGeA+cuZ1cxIzVHaw7YX
Z3Mv/Oc175ibyacfc4OU1qvBtOHmOecG5VhTmWWywdMyWar2EM7AkZUVfPVarEbTY80El+eFHauy
ptf23Omlbj37yy6H0j655A/C8maWgIAd366i53IXp+zVsJHNOLQ7S6yg7j2rIBIMiCIi78gSvip3
YGH/Qwe9kFp6JOhXkRI85FlKsZn2aQ65oVQZH6bEKuvSV7yXMrEIf3Tw6Nc85x3NFPCCg0U99Kmj
4y4gImYRtY4InII8l/2DNAAFKUzDrHewsnmNEpqbn54gwnECMqhp0XPg4jUvKleoBe15lIdKR1bK
yTW6MxMqSK3Q5keUFs3D7q+KloxEd5Mw6N7l7rj0UsZxLozT93CzdoW99Sit+coSvXq5NwmzmXVZ
Za96xKBh2Cidzl3/XCjnTBJSxYt1dx/7QrIN3sCKn0uFBEdb2YJyY0DSmM4Hom4iD15y045d58XC
ua23CrE6Mm1cLvjAq5hmKTd9STZC6+x6FiWsIbSvo1JYXns4ldgPbPJ5XQCVFV9RjLSq9jP5g1bU
wgtulmzXPZ387lMcTdOgAO/lDJq3yM7vO5KBfrxkcxkUGmUsb5g/pCQy//4aK76P9aq3c8M7WSbd
seTLjtGTe8iE1IqOqmHSuO8xNvXT2r/BlFZSOcyHQkbENOh2i2+pMzfSuYohSjl/7Hod6DOQLgsC
2A5vVICt3mGjvtgd+j/zbWaORfTzmtDz6yCOR9CX2k8h8XmzzIEwIJgGhq4tbIuiX511Smvpi/Vh
WDoDBCg7mmRshzIwe6kB1/4Af88Oza3nC3Z4clerLF6v6wQ9xRIY87ckGp9vVQC4TKV1GqGtGGGk
EnjLGP5WrV4IsbXiPcHQVSWboWEELktlgo1K4YjFkXz61VrXDkJxY9pRflULhP9KR04mqS7l8hDs
V4aCWlLGzG6TgpCk0g+/Kfgod2q2GayCrp8D1dGpmSYtHDIB71pwQsCrgGInqkdFT625hnJLmefx
mP0mKAr4xO4Nz8iRSIMnCbO4LnK9GMKEKIsGfGhcLVB6NRqAMbeiawG5TE9hh5bTxn+9sl5GPIBd
Bpmp1qptYe9dVsQEtZ5bXWfyIaL8T13bJ4BmFqGO/c+T6VGxYA+pseK5nonUnIQ75x9YE9CY0lLK
PmwEYWsgeSNawLUTP+PZVaEFXHv7Pti5DwSkquscQgltpn5w0apT7J9FvYDz+XRn2vUbOvVCQDYS
+blBWGhD8zeVDucAPs5Fs8FUjsrooH+sugwM5omUFxKbYco4MIpQIvGsNNEma45Q0GD6aE96kfUG
T7ZV/17zmlEyYSyZEFYwyfxZXjqSdQflHSSwvz2rb0dVgc4MbOcS92Pe6W6Xu4VLY9KEYxYcrLLW
ApevKKFEWCo99pkQocIG+Lgt6G2QHdCQxK5tWV7QZd9OwA0BcKY6t33OB93ReT19EU75JEgD+2ug
Gp7TEhZe0ZzOmUkKJWHuSeXdD3lORXnDgFmbkHpXmb2RqnupTiLT81pCy8tYnZeorsgqJvWL3wWg
yzd1lSBcY03qPAqz90odePp2c2LagqldP8CqA7cuBBO3rKbbd+D19yXz3rL70bHnO0hHApc3NAvo
OX4q7hJL4W/q/9qYM3peWGavNh9hslEGxX1LGYXSlA+jucbsqdbZ/z8xLbPK+Ef3opojQXitlZvO
r8T49id1wRcxwZxlVe/cU8/x5Ui41h5/Wb7Qhx7ScMrazeHLq6SKflJJH2oevNKqK1NwKwmM+2B1
mLyYGJSNACjbsFsY9LfCVd7BmY9yJDBDeVWYEvfnRfqVWtqIRkBkdPXGTo0C7fUOkbVvvZ5CUQQ1
cqTjhXt8mFr/QLnVZQEHJb2Vo6X0nqNMUop//D6gukZzyVxCD22i4HGhmx3m7jG3rRvPnNfpmz1k
p7LZPVuFZciwSWIn1qs9MNDKe9UyJnERYOUtK9EnwtbcTbQV0rJS1lPlg2tFHxcpAj7dGUS237ge
eyu7yGo/419Iug+nu+TeH4x5f9I7gAyMlP2qcpS9WMM1KTEHPcpFSMCYN5E4JScRV7VgsIIkb+6K
Ak87Vl1udJsbk6Pwl6vvsvm3u32VOpFmoHKweflFfsd6ihXguZf+PellZoHcsPhNTIVDochyXj9W
fNrCgDO72QYgo/W+52gMNgIC669iApHq6xpEB+gcPcrPBFRDludTubGDZaOp1z30rFPt985T+M4W
yf+vwlpuZTVKqzI7RP8dIF72ggv48QXaMzdtbif2eQhIXuF7rctRBL95Ks1f6j5GSLezMZVzlYZo
czaJCCBXM5cwnyIyorzuiooTWM5w4YUNdMENshC9+QTVMTG3mpp42A168QxNK5Jc9qVD7pgTBQtQ
nh5YaU1YvSe3ZurTj1m/0CvY6Eo2HLokRYt/RmSX3StKo0fPzayhkrUzrxYKefckQ1g1AZuCwYJq
Xs9544iExCOD6RI/kdeOVmeZWxnZrHcqjtQBaId1t2YiZLO+OtAeOCtozL/fg04GMnyHXTNAHzJS
sCy8Ain6Tn0P5B7Z51J0vZNuY8e7Rm4riALUXWc2TRowF8FBUZN5W3arYL73Ml/M16MuWQ7dAbM/
ux6WAW6oRqlO9u81zJ8STukqRxpSjjR/gdHRu2MJNhWBBN0wu8xra0eMnKlzTzAr3aeizff7WR0i
KYUnyNMucpDxiHL4b92XtRPoJ+X4FiN67T43aI6qR7n3HWGLOTpFfnZVk0EtWy+KdmUdnalIU9u4
SgfOiujy7xxvO+UINEK8Tz9pNw3yYm4nXJR17sbOdXXLdb0BJz7L6QfHRSAQA9dfOSTCGx/9+Dh7
LIUV1lp6oNjhFo1cMrn0qo+IEoQWjqZmZwRJGV1Un8yb3milfvV2F2Hpj3sw0S0h1mVF0r0rzGHq
yA25gJc2OarcHNEXntz8b4mFq9GYkK3hbSqIl/juH/QRJ09P2zi5DlfOl+AJ+vD9FG7BgMzm0C6X
FaNF/+Ab4LHZsJbi9pgBPDt/O/X+xQscXAjHXLsl+JK5OXFXmrsoTVPSrAY7AMZWjGxt6RtwBSLj
2sJSUHlmVOjRTWUG2+1gGbzef9/JKurcEqVZB4AFB8+aKyh1Vsyr5RItRVoDnamIanxz3Yugzwvk
d5hJN1eOcE2sQiGvfjhlhIIbPL1hLp8j38WpajlecQ9xr6s4rF8KL+IFEwlyMSMMbjd8SsoZrqBi
mAPLQSvMMXIfPKZrT0a6wIanQZNvv2GVB+trrPiUtLGMpbPudS2v4D7+f6ISZn8vfMW013JR3NfI
zP6Z4cYDCo0VgzvhdPzyD0MS4HQsZbTlhnZKWX2aX4PsiRKehYcTUBVsbfbpIR5+f1PxUSHv7vie
s2bNuzvd1NbMgGgmJa5QFiFourZK1YeE02MACa+RB2LaBRDLco3o1bf/qPc6TyoCYVsv9amzNbkI
gZZi7LgJRcjRQEOWWf9E4y1TJNhYq/raXSl/3kHCnIJN+LFgVnW2en/+hGqcDCWa3FzSTMzX8z5/
Jbmwc9r+3UXaoKOH7q2lqAZcT3FQdqJuY6ttqwmfFGkh0IUfzbya2MAvgLIYGMXxS9gg+YTAd7D4
Ia1saTxgfEA41Ci/OdBDCvEGcfkbLd5kO+WGCQA/ZPkTko9qtXkp0Tphn1VVoiJfRHVt9GSaalJE
wxT38gSjSOus8hTy46Di1CgHsmLsEiIZpFlpDZnAnuUvJhFoYjegm89OgLT+E5TUs6mIvf2YsLae
TvSjSWv2HIkGcCvnTac1P7wQS4rfIjySwZZhFCAFNjIXga7BdXcP74pyvT9PLh73CTuI5jFqOOtY
1jrcyB6pH84mnGhQOWeUvwPRBK9bAn+rM4HOVOCBURqZW7dMzJdaTxB+kyGrx8N2Q9kW2DVkbV+a
2r/U1zjZfGiVvApdu3FRn9f1kc/m7dsW1dNuQt6vbEYKubZabWJ1jQr16yveDPuuRWiK41a2QK6t
NeyuKH5T4dMuYm/qqxY6LCjlns16qSwDClMgcjxoV9Ajq6l0JdynrtK4xouOgrzCdY7H7wn2rNvs
x98DrL7MQRoNx3sgKBYWgt2ODzHch3BrSGwozoZbPyvQE1Ssobn4uyenzHBK8kw+w0hkMiOgYJ7w
H++RHcMnNix9seMJ2m0d2GziL9+w9OdpsP0PUPsPaK4PXLVpC8QsoW90NGljid6/mQgcRfTIzh1L
JEyiMICb9UUyxtWLyEoSQjm19yY9fu9qTUWk/0I/DBsVzICod0uXNi5OZk5Px0AAZ0SiS8o3EnVg
wSGeg5C10QqxIlRdDZR7/jWXwUKOiqOLNJpl9KtSAI0C5/OqcBzFFkLEtVxQy4M8xw3EXSRrKRMO
4a1lZUd6lTdkKB1axrj2fOXcFh8gRUVYDAn4/ZqLE1NeB3pXrmEl5fyGsLzfzk0BpK856LdWunJp
J4Fcv0c7qZliskqiwI7BuIoIWe0fheFqJ5sgabQOBN9yAmrMEMP2jq8+SLX6aCbXL9ryv8SEhbOv
xhRvQgw5UzTmwjDswcJZ/YkBV0UYlgQkOMg31G3Eg0x0s4oM37yha4hUM7fETc86loL+jwWrSva1
rJ5UUJsOACi2CN7X9AnG2m5o+CNONnaAT0rh/yBIbYFsjopQu9UUAGZKvK9gtW/n6nfh4MnTT68F
kGD3blRRXnBLvmnwJS7gj7nv21y/Gs1s+3KnsRlJaiYObK4KE7IgR6PvfL48fUCs5ua+Hlojip3q
bq0kINrMee6g/x7ieJ3hqyQKDJtzp+gQDlO6mcGSTwtk2YpX0qLYp0NJmT8c+iwj3pMoC2DvgTy9
bpQAgLiJuB8A1WUhit6lwA1zbEniUs3cfeDPQnTLPz53+MqrCHJ6g/qiC/7OjWD0GA4KL0wBtVXz
u/TmB1a6fhklyD/GfSWhwVIpp4Rsgny8w+7JA4+FMwWflAhKislSRcH1s/XejSOuw/SFf4/rDtr9
Cz/VGL37SH9H0TE1AZwDGJyV/P3Is5ubXC9WdwCqUaTeoPmabd1E/bxvTvlc/71XPao89l5c8Prd
meXV7mo6dNuXL1LlVT+vwCNOlEYSxMzAhN6bZBex7KvYLUzGpiZMfx5MWU3I1O1I/GwF5ff8y3iU
ayu4u92jhv22g0arEGYpVEywsBVQhDt9EEYul71kqk3XtS6wZUCBE17Xvtj9uwSV66koIHGz4/pQ
QjHo1IuRfsGR6evxWB7zWbtw05FU6XVM4Xxyjm3c1CQpwNT8aCNr/yvypF+Ra3HmLarIJwACs4kG
VojmncwvEiqi450Sh2YKAaSS3sGFNsk6udD6ukJ9ZG0BFat+p6AlHBfkOE9fYZP0PFbCOUi3eL9+
0fBomz5aNFFshFMZTLQBeVk6lCu5JWjMPS+K25PhIHHpPD4NAwWskWx61DJ82WzCE52Wg0frx+1r
i67FwSGqWQq+ErVQV8EhVXb4mJF9VN2MnHK2FEHjRE+gmITYE4raxoA2+iukMUfIs9TMpvMC1713
kKGjoJdL/9tBlHLUedtSnHFaXd0Qek6GeQm+ynEEK4V61AQ618wJNCRCL62FttiWjNtz3VZVWG1P
G6lDEJzQNSCV4Uiu2WfnxMgTXxTmEdvHAtI/rkZy+blnbWsVqy8rkHMCTe0v4tLWrqD5d4OUiqb5
YyC3Bjc9PGI/swYhGzprX2oy6WJ8L86IQUZUEBFTo11oRgOSy853rn7VGGtgwamPyFpL0xFMsUjq
U9sx1cVEV4oaYsDzh0m4PKygUyM0DkTBfzQcfQWovNg2nAgsHILGNkjChPkpGj3hMt5+9KpFLVZl
aRRn0VyBhUfqN8o/HAd63I8XUnUPHHe5SbizZAoBdlz1mVDo3t//xsXua1OhMJyUm387orcchc/I
1pdH7m3SEcGbFBVdQ+ubmacAJO1NmanGMCl7b8gg99ZGdbn0Hxbz8V/KxRKpJL3J5oEy3qynRQj8
kazWlS4FAM3iqlwJ4Fwib5wQpCNalXK1wFj44Nx9w914ch+TU1KYiZgRx/fMVVZQjjjZA325SHcD
KlLqEWZHm18o83SWUzwNWiIMaH/2y2YJmTMT6aMp0nwjXTUbMoo0bX6ynara6gLaozJah0RKw2X1
bnawiFw/ZBVgWVxtICjGlwbESvO0Ts+NBhE4QK95NlmcRO3PJhVRGthkiK55cgAgQTqmzpNdzi5n
oHcsBg6Kxy/ZjRBdnqI7+1FIoLGPxYHJB1xIxqNxdNYFmeKLuqKNHXNT2Em6sF5jbTEp/Cx8lqSf
DoCaeuWPL74AMG3g/Qb0UB17tIE2pRrWLn7GNQwml3J6mDACqZBLankTZbRuS2UhyecGYDYroagV
9eXYIdtdf0MShvUA5HXb7m7V4m1D67Sr7JOF4ZirPV3v7wicSVJRU58c4QoD4fsZa3ttos14rwrx
wKHQYl14YEQXlwU7jUjKREpPqEBYGpRUC8+roxTjYMjb+DFEt39ErObZP+AQDnAMFMAlxHfUnJ0p
ykKDBjwwTen6V7C8TmuvHhKEFiaZuaIaAWz8eGukgxwg0eqwgcP2HzPka2HZFjh5BXdE3WfOpKJB
jxLDn/rXm1sMcvx7HqbSTwpRRB5iLbePNU/YGPBneB+jbHTv3Vq6uqLa7dyZ7cuQKLkmwh3MXzoz
ty8YPIlXcMs4aLHTnyddeuFPbQVEn+izhVRJ3BgQof5axyQxHAuitiffvuQFUfts5ERQHHD1nrgP
C/9W/Y9FgKR69NjgyH5F021mZWa1icHnkoT2lS/i6kTgiJ92aFK2NtzlaHGo79ImIB6FSgpR4rWq
P0R6N1R4nxMYj4zw40f3YksN2mBxaIEytXi46fRLwuMMR/P9kYh9TKySLHvCmdtD2XDKHnLCW8UQ
u6Bpw8TzMMlyAZnc6r+7RdTXZQ3m1MM1DBTK8V1Vi8EnchGbcYTUsYCjhHG56oA6ibgt7FBfczhF
acIrPs+YoxXa1MygIS82BQZmI7rv9W0MaSPN2a3U0cOAgdOKBhNUhafHSbyIrCI52uzGeqVwrdnh
u3zbWd5AYJygqTq6n2K6NhatdpcKOqUgrSRTGGwmQA2BIRpkAF2Aa6tUUBFaWhKHeNkHGQ/t+sCm
t7ZwmNdXJ9EM51izys+dnSMuWyVdysfhNwKg/I+hwnebjSkJ5TqGEc13Dkl9O3ZB165EawL2Y13e
oRi2YXo8E4+CDvXZc2UyKFpxA6TeTEroyPDmj1GcL6ewJbty6ZqoNDE2tW6rL7ltCtQCsn1XyzCa
4t3H7u57WboHizvxWddhDT1ElATv9WQ8JrYY2ZkV81addB6xTwGlsYgp2fAA1ONnvETeI08br+IS
Zj030RBa4c7is35knikU5mkdn40zZ5Oow9eYQMbURBvnimeWbXgtpbceJ2L6ftx+O1NhYaxyO4wr
WlRkyJeL14svnDcjnpKzKGfqueZu433v+fKZSjMa+F2/I8+TAWblzkMCM4wMfC7BV66TbfQvZbXj
695I4dhvLcV758b2ShU7aGHf3aW/9lPK39FpRpvAyVEhbd00Q9L00NhR2afdt2Gf3+P4B6kvotaa
S8VlZkDDuZh1sD7L21MP0ile3qEWPnQzrcfeD6EaJh2qhVghWZM/QwiDOfsEulMEAbvalZbFI2Eh
MnBNJlejpq/hqEYh1G8lfzq7ulsBcrUhbp2pi2py5OoRF+12XPeOVuK660kKFMdMVUrYhkp55J9i
4IXX30fMvguToXXWR3YaR353fbloqQm2lI9JzdRYsT8U0lpfcXUodRF+dqhSTVcnca2rFdtGQQrA
mojDCzC3CoisgSeeG1CLsTGUlEyXAmgQIoRk0oRCFImomQ/Qv9SyE2+/Ko8ScNCBD7eGAHPuTfgx
7eLijtOQfOa9ZdkR2KLAI9ve3VN/aju1Gxk2X1ypeVlx3TA2iWz4qntIC15/XCyIHEzLZcx6SYpI
R3nHVi7knxomVF2V+VHZ1KOl+GmADwJbY/czxHlFtfwgbXdcbGSXihK7Nc1OqSnkh+9vZtIHgSpg
fWgbX5STxomAhgdLxBMRLsla/q5U+TwGf/F3uazX4eUjphyvkGX1acedvGnnalfp2lT+MgREvhII
jaGbORHq+ppOBVSNZNKRHXJaZzRr1Wohr9E6Y2IfnMoIlPxC6xXgFpXrVRbvUcJGitRfs0ShLrDY
QqsTUoqoYlMS2zlyRVIODOLduW5zZH6HiXjZ/JoLSP00mFun+4NXFQDzg2rZ69Ox9aCrp4jSOGxD
+JmZBNMGOGtbiezKzH41ZGqT+g80nYl5Hovkgyd+gGhmRmofxjhkOCQPyP7xRt53f3yrKlaSzYrY
hR2XHawkfan5n0YvYnkDrmOBVRZCPUe3bgFJqn15/w4+oVGpEOIJddt8EEX6v2CG93c7446xBhnn
sVmPlwDHt1vLCsB/tM3oroevy3nkQyYUt25GWbbX9p4pAzsyHJPPTvjQKILblXUyKR763678Yk5l
A/z7cjsjN+8LLAbCYTY2Ko/Ni+SmjH2JohUN5nrapqJB4ZzdQOfJXrt6Rm+wLIViKaKvAuDR78NM
tVwa5HJrGzZ08rlERzONLP0txcqB1SOoa2kmq61Uu+jL0QWT9z42VAxn2SZhLVtNFuH4ZxS6rQYm
7hnclz6vzsHkfMYDT4FbSWrt3qW8RBKFkjFDu1hnUlmot04g/3733PHb03BBYhGo53hrzq6wC7w4
uVHQ76f+xzico6zRqOQTLG4QgkmRvtHUbTpHx93lv/PiWyTqiEe4vNt6IHhz3rA5PGBQtyGZKzP8
an8v7DbwLn/RSl9bwt/6W9dnAVqGi+TGLZnQfWY3Dvqw9jO5fTH/0FZ173dGr+sKWdDZ7ghR7LI1
JscKGpQACJyRdp840pQY147rBHp40/8WARkECGQ72CWPHscfEhWeP7f7AHxyrNphMsQU/u1Pxn/4
+nyky1N2hWwLIyp4I5estuD+Coo4ViUW6SLWAMu+lqphXGzNSRXLlyWW/w8vh/vqcko6RwFWBBfd
WeYebJ1fUHhIyoQtMHdbTA/lIHzFw5K7zxY49mEb/0SM/9nMWN8VhC9PfK9SYvEcDDkb6D5zZRxz
jQhTG9RV+USxtW5w/eGGyf0f1g/Qy9Imuif3ok6JAuZogvQtFRctatPQW4JdZZDi8MY5EU+P903z
TCGg/Ep+BGknme3EnDzRS+Hlny/hUHCMQ4MNwLBJS+vXas5d+wrSngMQ0JIQdEO+DSvv8awtF3am
MWygELnKcckity+6paQ3vsLueGjpBUsrK9JdAraPqNRcRd/3e5jwo7SuAcGEmLThK7Ih7J77fsSX
KXpLO0fap/hlmeabqqekNaiG0jMJlxfbjHSZruabYJRdg0ZPtkLmm0igoxazAJPXeeR2TIwXHwNk
OUkEyn1tm9CEMU11jQVWH2o7vZxRhaqHX2QLhT7u4rdgtZBAT0uOKBh434TVVtThrlxET592Ffh6
rmab+uFW78k+McFtVoFBgI//oJSgMvVAYNtjG+wRBZwKqW84BtPEwOa0IOzCuA+8IDREp9AaouA1
DKFycks00ig0T0DWyMKyM1zMGjukuVjIBSH7e7pZrX5q2mrx8wLM0DLxkDOkHBHEsuK3yejzARp8
TLHibJ1n0WyeOqeUyYJyeT+YVKyoCUzzdzqxdnz5IxIebOEqlW/2LmDVJPzmjtDOdE32FIhxs9oz
oGEuJqARcsMO1kSvfcFSRiRay9/GYLMb1Jj+V+QUIoGPlRXhTqG/ZLbTQPrvPhM0e6eb5ZuhztG8
9mY1iRqoMevdc3/RloLfgmpwsQHC5u1EId39xuqUCEPp6NSA7lFf+fZmYei0WAq17RBCksGbSHKa
+BB+x0jEnCwOwMlypGVOLSFxIkGAW4IASyQvc3tvOjw1SVV4BgIPOVN0ZVWsj7v9dwAm1N0h24kz
MPSaBNEd6ruOVFE2/sgZAIr+S2CWZI578MYHj20eGU0n7c6+bbGvpC5KnfWNVvDQOsLNQhXYwNc7
uw5Zvu5HJYYEJGQlae6Z+asTMkB3QJmuLXB0LCkYsood2ZHUYb9O6i2hphAgiRkZkWhiRlvTV02/
SOwRYZyVMV29DqtklYdgnsBTI5W0Dk9Z/9jy8Mwzf5fpcD6WnAUW09wWuBEOomC8PqIOF0yjOJWC
lhvFTik9P2o5DWOEQ+Al61N09W3eM5q/P6LaT7pOFTT9eX8EbjaHTXweZMCdFbOpD/MQRz+gMTd1
t0VZ+/bKz8sw+3JvSMTvMFL30r8VntPIOg7nJ25GTIeaDa6tQZmWZkBalWIdi7WAPdTFc/KX4JHk
yhStFyZUxryUnBJaUMMgIH4ExbrjzQf06tCUeMi3iRDo1nNDH6ZzS6hxoNG/qKjW75SukVd1F++t
6jvZlBVseDW21gDAXLpHKeVjhf9o29sSTnhNDE+hwmdgvgZRmG+5/1rMl4tWL7WRqR6juQKk+9vn
iiyoyoHCschbMzQ29VeJ0GKpR9Vj3XGMhBasXIg4yQV+KMz6YRkxPdD8DlaMIuIxn7P9Jlaj0NI2
P5Bi1dTWXQfYsZWu8gBuIgIhjcYhfSxNmhMoKxq4o27s7Bc0wxVWxtqpsJ3+zYp3kOyeNhGsdot8
NuJsyzr4ZCeNZb75fcE0BGrvx1c+2dnAtmDn++FwRjwZinoVDQBpFPsA3US1bg3ebYv8yJKCm4c6
efxAPV7sRDJ4Ir3SpSxj38V0nchLCLkof7tcKJVQLsXadinqfKwDtxgjm+ktCpEyR2v23Qis7wZ4
zLTFjHrW7XStlDXew7UKf2qAxS4RYFHzKkXPPNOsU07Rz6PVmATU6JE/pi6pfCK/fiSyL9rCeIoP
ZPLTHprmHRl2KVFSgtmFvqBteIEfWL/+58hGi+2r1OP5uqM3VJP4SOPf9VdIt6asQoqXeRykVsnu
Mpd81fXH9es0RB5tuOl8gnbFVQJ4Rw4pqJBj++P/mrEbgCubLCndHzwKe1Ejj88AHCyk5xpKcrrA
gmMaw4UfFz2FNqlY0Em0KvX2JYLQ+3IsDsGhlr+P08XbNGVmCEEq1TY8VV+rChomPJ89+J0HtOcX
soGfI+gSXJnVjg7Ig9J6WI/l5SLxF1Srn9StVbVLQEM7DNhLp6ZRXBo3gMZhZ+9GVAkZqbpepccM
JgfUkj45kcVLFn+gcL44aTZ94L2Dd96hXSCyCTfLn1nzh1OK2HHI41Uy0utQpOn9vvJFuC/gJUoL
nqgLbioMNrWFlu+Tgq9ERFuaXGE0q7H5P4bnN06WOP4fL37470u1bFOdzMA00DJbBW/UuEQhPg4+
NjwxoRx5HA4RbW++0PsS2jZMPea34+DCXj872eMB3HX4OMDRc+O7dvSDDze7F4ILFR0OpWwVszh8
JsymT6cIyw6118OP222lu9Bodi4WczA+Fw7ZhxuxyomDNZLzS3S/FEgaWwsaCgfHWrx9hVZ7nmSW
gf+tteJn8vE5Q4xJFUDGH/6k44PWZpgBMM+FLG7VTe6dnhfd4g6d483dU0i7KlVvLjh2szYNrnhs
zue7u4aTcGxHrf+FJC5T42fTaa3ADS+/pWw+a913SbISgfrRfwo7/ELgye4Fn3UZ5z6ZEhiLg1Y9
R0tGDtHVokpiXmteglQ+wz+8r6zIWM2hohh6Eq9Xcdua9fTfValixbpHL6C4/Y5NA7W3/Txq7T1b
AGA+z0Xpl7JZM/YGUzcPeatL+dvZlMqN2VcW1zYF+nAe6J0gBrixn9DlNjQ7XLwTcoYHj/w17BjX
cS2QnOdl898tfRo9ZU9cn51HQDahraDA8d5jhPOquw/xOlRlNl3vOQ6SRRgzpumr/fiD0GPUvxje
dxxITsElx17hGEjhHmhTIU4B8GXfEy1ABwD+/Hwjj6jLSyhqLv7PACZQrDrJnqYnmBu6hALUqBSZ
N5k6To8Tg73Tr9+OzNaVq9mVWvGJx4z6wxbrsPUgAxrgJBnza/+MqQqs8VsAZdvmAdu63Tu7QnTu
p7irLINjJL8LqCiIVmNUezd1HK/77j6jwm/LKETI2+CsiXnhj1CCVtl2pNgQ5Xn/D4Uf9YQ8SPnt
x8vnqGpDA1d6jDtIJx2BD/9bRFNR5ONWQFN3p7GeNeggPlEycdZ6goJjR2MhhBeFcneHDUDDSTTf
GwPDzbT8rSMJ5e2bw0CCDexmEE5eKw3IQM5cljytb6ee+CMffMG4W9U7h2Xzpo/Tjtb9HajXgu6N
nwl0I5tBHCK94jJqI77McIIrMjwKCI6AJtV1uHT720vz8fBfD4XsaOJRJWzATbZcxYVU2z0HBmgX
rlb0scD9RHuzUCYhVqz+CSYaaxTxLkRwxfoSEh7J/ECHFMzzvZCsGCnlz1iSSzIVm2tQntuAp3Sd
RnT9sfl+Voxau4ePZoeDZzpYwQ1w0o9y+Guk36fYXDIAu2/R7xiCWV6KnRhDxIx/yKWpiuOtJS3u
DtZrwnc7lmMJ+KDdp1Fvx/l4GoCP9+98liTUfn9+uJM9cRsl1Pj5i9Za9bmGj+TZl2iNIBg84EPp
2s6NqycPRCzUAzIVeP3G0ZU5KJFRVZN5Tk9r7GTcd9e9GliIQNMoWCBeo29l/xMfWEqFPGWBOQjB
uqG8JAMHwR7rfSdIe9YHpHWkENmDi987nCf1LQUxQhP/M3TdGfbnkP7jpqstQWctL4QTbQ1tOBNp
HjAvXrvLhyKW0g/DLhc8Jr5nv/5SOhaRrzgawIg8xJKSzkys1ZEEXEz3REn9YfHciYScdE7oIba4
9He+iz4MeqWxr6v1LUclNKjZkZHBJz+d1uw500yByIoRFN1tIBv2viqdzLHEBa+ES9XC13euf9jb
c4gmPRMxBeTZUkMYj9efc2vCSziVAi7fJ3XBJ6WSrXBXvRd9IGSPgYCtsXXZ/9LbSn7qh1pAyaML
/oCvCA1YHHCVXv5xPW74t5vG7RYoltSwRjd+t8GqBT9w3VwLjv9VHrjsyBienRBq1s4+QN0f8euC
8Yc0h3uiE8XwQiDmXrqrnybluqwpdQ1crnTjmQDAbXqDwAb073/yPu8UWraiwhxw8aamq4ctMW8K
vB89c69U82dxHXOsuEt5Gw0Ijila38DjH00s3IM69JOTjP1faZ1+hxjRDTkxFVYckF/RLFbQOupv
fqyVSMVty6J7HZejy7gLLzJTDbFVwkG1Z0CXIilfBcASY60UhF52po7/+7uy6pfXLhA3LeEdLA37
PeWsKpIQC8jJIEpymXkkVjlevG0VKp6J+o5bWnx87E2SI2iVHBtpqdkRJ1nbd0kOYJpfoeN/+loa
0aCq+IRR0dkVhUD/kTQZJhuEz8TPwqovuc9FvhQwop65bQ7p/P4dl/DS7Lka179rafG+DesGcWbh
oU11m5MCajqqAHJ1617jMUSqb4cWXTZkLz2f6jwNS6ieKO7YqC/KAmCS7fvQc+3RtRJLYGn6PNuk
QwxPBluuCsbqRFXcp/IpY+tNOI3qv+0E4DBnA809cZthzAZYmj84wbQy6nSpHvuSbMRTi6YH4GTU
vLceGUIoZ3Q/sNZcWqpvpx5jYJOosum3CFNimsXPLdXKXR2XsEes+F83zYlENbXWi1MFjLQxdeW/
/UZ/lB/sGPiz3ueCsnehPnywmyE16iIs5T47/Ey1tbZLYJQyIPeHnlq7lzwLZTCVr2NKbNVK7x23
9XhyH3a8dAuzNdXtrTwvlKD0F/q7+U+VDChEIHyzoAnq7qB8aGhYBTXXb39nHoznOuqlmUL14Tiq
bAN1tzNcFIMClOc9Nqqm39EACG07E+L5L3IzFbyVGXA5W3W1PTwPdL3SAmD5Phm+K432GiBh7seV
R+IoAWzd7olphEdo7NCrPzHMLk/ZSljFdeTIoabPyks9NQaLV56tzPf3kWzp3meWD3QkK8q7J8Uj
AzfbDfmoi35nwXSHP5hcED4KfvSFHjTGBRl8436ENkuZD5Gx76YZLF17ZiYhfXFEOI/+LIlLYPRV
ptlnNp6Wo9b3qzW4KnUxZ+poAIVQV+GBrfvSek9xWUPsscDfG8G+5u62a6Ti1MiOHH4URgHxxVbs
zOfC1NYDtB//lKd3fQ5sG+0dA1EUcoTGtbB0RLC0NupWmGjgbr+KP/ONnBYG0jyB/G9+F5G6mfvu
FDgXBMy9sTFH9CCYz1jjgRaJXjo5FbnFgyE3qLc8T6S0TNKO6S1wqkwXIJ2Uo/i6cFRD1zyDlq9o
aDyqNOOHjGt1QmzzgVnkILm7DsdASANVdiwJA2ZT6T/qCSJS04xxx1U7ggU2fOhzFQH2enLEaFz4
gmvZ1T1bLByoauRQWJjlgAkAmX1BT6IOxx0GVSXJpPuhtvBAGTRshv+hm68lNA9kUSDSrX1jhGSp
G237hsdPkMnTXYZaOagGspbfu9gO8FOOE0Zs1bjphn5eoiEeJJ9cq7EI4TGYGOblXyHg8ZL+Zgdm
ZCiEnHnu4H8kUqEroRfzBZGsvgC80v7hGX8G9Yhn4O82f2TK8zln2UKAcDTgwyXn3jRFPgvrwB86
CzA6LvApSTKueGLufNQJUOQePAKIOhjxVp5dWZWTaIHz1XWARTyiK3RY6prbJXlvdYRyNvfqCXOR
sqt3m7+I8ERmDsGunLRb9YRjFIQerKSIkRfYWk+gBD3v6YZyZSsHwxlbEJF9E3UqjwFEHtmnyMZA
6rMBS+i7/WTCNyBNS/qNai+T5+USzw7cw4K7FM3iidnP4yJICrksHS6I6J8MPD8KUviX5hRAkqIJ
mWrhP7c7S33FfO8fJjTEf4OHJN4oL3j/lS6R3hHyysBFeDJ6fnuDk08I/sGqX/eh1G/Q1RgPkujA
wN1rVOjbMSRfgz3cQY3+I9FuiefCUFQHFtB8T2whWS2UGZTpWdJ2xVoX4pePyDAI3S7u7od3v1pX
FzVoiqNIasNAgVJcKJ7EPRTJ8qMqO+lz/yHPAume/bjW7bz/LDPMpyjVYOHCupJfO6+iTLe6hXri
337UL6hZ3a3miY/iyy4Vv5cpEbRQwJK40FK3I/zAlocRC6cSeoXSRMbbRabkThI0XV2kilQ9grDU
YpXVBkB6aBiMQIbF6hiYbuwPsXM3S9o3jGngBC7t87YBMHZybokqk7gcMWdHQIr/tw6AFuQ7QrXo
fqF7sx4EA6JbQUc8CqGZfJiDb5gSSKaF2Gj1DNYIUmNhZ3zPoYDArGwUOfXVpiAMv247O0O1519r
IUB3KeVbAFGgibsCjX5p1fF8rqYM9dKsNwI5e4F2HRDo1bvC8pk1IqH1yBLUqxJVwcSRU8vN82lz
5q77HAf8FJtEOhLbg3ZYvPUkWHk5b8vl9E5fvAP75x6++I8FnmHh/QJO8IRPwVfln4wlZmaHwieC
Bnz2pLbqL8v5npOYSxBMXfv50bRzoMHED8J4ld0Y2l2+Mszc4dHUeXV++7K/LsUGrwsriyETjLRn
Abh7hoWC4Danst80MU1jjf6MlIDJacJ0lGFTOAoZit4i5IqynJsAzFs50I+mFF4vgHqXr/Bx9k4T
UtBBJLzaeDmbUEqpl7A3S/r+k//7Keb6R08Bt5aPpnh5WueMmDpMYokLeGF1B30BpdMY7SzsRub2
8nXJ7Sa6a8zWR3UVNBjR8lftG3coXEg4xFHileU6N5TJThJI6sYRs4DAnmajs2p3dmgrydUo815O
ktc8zZK3PyNzh3FQ0YXneTDK/dT03G5ZpJ27ENKD0Dr3/g2KaqeDEdrmySzVqrxmn9ntCY6tu9VX
fmyJ3iQVyP/PCODHoJmjlLE1GhGkjDkIWlChLGJSl3TUoM4bGzdzgUg/gu2KDo/VwftvS8dRrRNp
aMR7MrzQebzh5azGFTCZ1Y4WC3YwGAIDxwwFT/5eIpjbF4fg0Wc85xlAjcaeA4XTWAKrdlZcRf2d
eBvuOB1yvlHozJvsG78iag/MK9mos5jTILlIxu5Z0YSN/ZXkN4Cg7PPbgr7Yvx2UD8hRv+UuEK0A
WLH/Uxz1cD+3JirjWJw1FHdWp6dEpleBrcEII9JUayYXXwswchAWIAG2AxDYA7Qv6osx0meXll99
cSVZvagbU5G5i63WZV4u9ybieah2h8k4hOZp2rkGgi6sm4XBIU61wcS4ThH6Ow0Z2DavNT62mch8
QIjpz93qrJnIqzhjy4ZpNfwWzh4UMJ2HtjFnYJqBDzXPsGo9mrb3Ntv3jSu7xMvIkYAHTUHCMgto
PDGF5dbEgngntogTPsYEWeR/PnnSRWhPRsbk4+2M0D/jkTjnT0Bvr+OhrNZymO2IhXWvv3urEDFa
o4ZH4tYBVkB13UKqW0zjSIYvfCZsunaS4kHca1Ag9BhZbB9ZD2h3MelNXtihnH3ccP3YjXqz4A1l
YzfOvULPfroM/jlymwATEmAOK1dSBTJCngIWr8eAIDcJeTi8cp9VSmj53w52jQ/FAcPhg9NSVOgP
t4JKLDmt0v/zj48wBA5/X2HVFgvFBxvTGe8spbRg5DEHf/gvy3pRnllGc9oV7oi7Rli5ndiugNw1
A19UYkc/qE2s8yjNvi2dRwMDGpg84kwmLNsolvEPA3I984Gzp9+bpmm17Z7qrjGrLOi9DLWqnnVA
Y30Foc4Gp9rhGZrQNQVVnduUi/xRZx1JPbpQY9SeKlN/OVuX2nWWV8no7HwExyksNQJ6fQ16YMS3
OXYtZy3x5VzkfHSSE01T4CJz3Bc4rRJUfGbNt/ylw31sRCaqhRawTW8L1bc4MF9+6cRRDi6H7BQr
ydQ3sd+h73PFaQyah1MTDSLaki1PV+1XLTxBLjqDlFZnyqh2rIf/XbHxMff3HgSwWhr+X+cGgJNh
TNBAGDAgrwhfP6p1UX6uTNe+09bHpg7sIx0EnnsK2gdFqBEuLvlAlfAWiHTjKJOoEY2uwyUHpbn2
jnm0L30xyIlgJ2myaI6GLs7114YX+23hNHbV6XmpJJkHo2wuHgxq3f1RUQpKR3y6swxrIVVgwnMy
AUh15rM0iPWg2DrPdRTweLg6n4myIdWa7VC0ViAjeix0lfeuqKU4ayD/j+HtTY/bqKGA2CEIAv45
UCxYpNDu/CdTvucTfF4QvUSK3sSgUy658JNYbZY5cvrU9/SuNIntPmSnoNY+ZRQOLbgEsA3xt+qj
K138DeWQtPZ1yK9jAGItrSnafc/bf16rOy+cKB1eHymrVD0dxgWRgYagitYXD0cEH3VfwhXKkw4C
2V7aws4xEDQBfgfmld+2SD/1Afz53kqevlu4rJZFGJAbdE7sgDFmBIZHB9ogygsaYCWElMsqmHvv
JErf2wJOTvXh6pggSF49pGyAkqnrIcYc7L7C8GLUk+y3RqpuBIRnN2tE5EmST2LjNLlyHjPVag77
ih38nkrxtz9xXZ5lhaMBX18wMdB6gONAhRm2jOx8kmdBnCcvmkyIpBDr087QExJc7GIUWM0Q4EiA
69/vhCkpbaYlpGZmsAf9wLUuwlyD4WTIvctL6ZTpTLeBybcUwGcgBu1ia4EyP4qnQsAGq0ZCi/CG
z7QtdUSuuSamjHY0galZVE7IJDygFIFw+/8BtrR2YBpXbT9mp0PYGHI4y19BegaYLZRriM1J/pyW
pmsYaX7NhKjauQylyzTfX7GI4L6o9Ar2Bl6bRKPuby3LHQQtiis+DYWTTyzcbxI86JYKUGgjhBd1
bt7sNEQQVSA3ZxQLdDv6Yt4wBrSMTQvE94cb8aT98fcvbsTs7rz7C7zMCgMoHE9fngov2kvwhfUc
zTohF9gsHFq7pcBVjW5vse3SfePx1yf3A1EAXJmjwhIodToVRIcJQmzMvSBLtbawGgXGI8HRBUqK
YolCRoe5sLhscKc8vtsp0uhlyHNBjLD+jsBhXnunLAGx5gFYWae3mWAB4123NDZG2NA0hJKuf7fX
B1RkTh1dhUA8JHkCtMYRP2dGgsYJFdPnqSTTH80ACYC+S6l7nBs6JZWXntOhBBTPW5QXMlRE3lNo
Tq7tsOV+eC5o0NWmafXVLDscn4xPfVBy9zxc+g09qfi9e2+1Qlvnxdq++Ir+pWPiuqEKpypBYCy+
LpsWt6S9zZ5gz6GvVleAYiGJRu3RLR3MyE/GmRo7q3JKMAmS3vm2XuvotI1s3M1vnqNk8E1nCXoi
N2q+UgnHB+zC6EqGQ4a49SdnvgAdHEH6AYXnx+Ef5dlG/6oiDsptCEW56s16nZYCIqX19reuZG1q
YagsurCSyb71zD8uj4FZraS0vMy9AE4mChzF/ndepoH5KfZa8leral+We3KgwxNIsVsu/rou8vmJ
qlCqBmQVH/PtRj+FE+SRibQ0uzMF3AOXU2MIczvtbq1Fh5JjUddwOlBUSipuVoXnDGXAGrwk0qwd
pa2L3WD6S3Dmkt3EFt2qoaXdtki3UtCtxGNn1m6n1Y8U8vS7H/HtR9r2i/pPkSX5529mvnuyT4ty
ZwhOThUK8CnxvVOjtbS9woUr+MJo+/x93iDmP9RRz+UigpauNe7ks0PnkpB8Ug6am83oWzLGrX2f
1XTfIvQfu4aZOGB1GWFx6jx8zRaMULmw9deNYI3CVy9lG119Lk9PEahKHUnzcFpW8ltN7AFYk3Gq
Rsq3MiWT+I03bAlE+3ctZtsiGQQWCmolZcsHgTEPILt5mtCzRz85ABYsMclGFNzXSGFNuyrc+MIi
CwGGhB8NYqgxCsCOylrlj9Fo0XvrSADz2SWor1YKWSB8QF1gEipAy9NVtTxCGDamNfQZjeKqogzG
CyxPph3og6vUGYaUQydcSPp9D79yVz+B0P6DZlnQsNv3NTulOVq1vzAnCzW26oBIi0Klz/q338bN
C39+6j45ej76sgbLkXiOaD8jU4OU07ft51TSR+LY6l34+YXySMiSGmr3cqlPkffc6MtrlJZRJQNK
thRgta4pNLk+yCX9BHLXKes7kEbgbMpFmhrPsWNgp5hNIRmeuNp6To+egcG7bTNXcCXCYFlgJzAU
xjyE/3mYcWWDNixe+AaEDTpBSID9QwOI/6hGpSTo0df9IV6PMcFUjIJCtlCknnPEOpklna2mUTvP
gc2JVlKkFwOurlkTZ734GUVoB/Tj4diqLaZVY/HktKuD53vx+E/Irx3TosUtyN4Tg31xcKfAF1Pk
tSkdywuqD2S2N0cJUnhbcvhm7IHIrdQzS70AnKXLGGq9qRm95T2SdkcZ9YZY4+EPkTTlibnpbJmN
sJsFkRQ6EgdUUkSfCLFNtYTLzbF0a3HniwstImMvWetQF7nX+X3kSL6rwQjOgMocXf6MmwcQPGfI
dYewL9j1uwgDp5hreiVEFJOgGAHP2ptUt9UeaW2bi82MbG/G/GtaNqjr9ZPFUYoY+gE6a18TwQor
EwLGjY7spwWzKui9tfGFGpGKPzulV3hsEydWoaXxAbzrY5UTv6tzlrdQ9w8jnC29UnKsfdOglJVK
lPyTsbzaFx9PrnoYTEvNlcXYcgHmnvMGkX5tn/mAYni8k2dzdWzLmSBLsXLOhedANu4lRZmFyPDo
7cSEzzdMd0XxZ8K9yhF6rlxbJR1zTm2yuGbp9amdhasjKlX43mjUePRxn0pd2HRCYxsYl4/6vyCv
X9h4r+vPWZ3Qm5LZE3vrS3XNxgsYv5ijzAu/ylWQAY5FXHAvPMlbxkeicnj57pq5lcHh/QnWrB2A
JpEexeKhQR2gy7HaEx5g91vMuKCWuSGNkE6Eb/hnHxLDsahAvXkV36tW1ZyJh66T3tgk9Z5kRhAy
ZEDW4o/Mt1LLQGxuULpUM0saNjHOybVH3ktwqvADVTbTV5CVBkynHakkCDoP6kHmZ93DbC2fMmAv
MgcKIs8KFjenw/JJjUH8Mg3dVERN5DWNfdBxTxlMsgsBvEDYgDm5DQ7QhT7A8YA8/YfY/h/8RACF
9o7ShE1gcXqVE1KcYp8jWw6pEiyFpvJoV5G4h72F37DUINGjgxa35HLXZupZdTo2o7VCxOlu/14n
lMRJR19AfyZ//OetOHL+6RObX8zY94itKb5qjnNNghw7Qer18GbjRKLQfC2uiFnSW1UnozA8fnXK
yxfJIkSCilJh9aySJpwWoSd3xY5EHi7Q586UjuR3nQIxoMdf60KoduJav6+XmpHFLo8pKq6e2qyP
PLLCUsv2FJR7SjCuVHVSvNaacsMevkAAinn7KXn3i2Ya4cJ/P09It1xV+Synw3wkvhBKMaPduuzm
C410b6a9U/FRoGxw8PH/7eKQWL7aG6Cdb4f4k5boHzlC07ZD+WY+lsKe0gu6EnNrKCQEF/TYg/n1
I8a9aFh7Dga0uEuYpmUSq4+6uIJeUHGhTtacuG2JM0zb7yp02rq2eaUTeAISwsXgqKebQrnTdy81
sU3QGUF1c33ZC4vgrRDr3McYFG5P0JoHgyI5SaqjsUOhTo5Mr/GzP4V+LZS7oL9GSULzaG97NL17
St4/SBH68t4hnP0R9YAccic4e8wsIBYQ1MLghWxi+2kPcHoQY9ueT5FGx1lAeel4C1gtc/3HXAW6
m2PUjh750wfODdBPyrFfHRwmNQVhwWrnFzAPxN1MLnqIqTNhvTfc+e6EiumkO6OdzvLVRTpaSz6f
p9L5sGjcfl/k6FD6U1PpToAm1RnAMKFl6z+G0YrprePhQsqwyEyFqebAJYCWXHZQhWa0X/GAsQas
K3HBbc37QPLwnucOlNrRXBN4iyTLqtyNVlcENlYDXyB6UuUwly6VFaz3d9VnEpzqbhxAlj6i9FeM
OYp5WspOkp9hc8S2Qdf0+f3z080KsYA22yYzBcNojvq1Y2z3TM2anWepOx0mWfq1jcN7xtW6kPgh
d2kErvBqseJmleBYSNwkciXt0oEnZkXNs2ukW0jLxAlsAxw4KUQX1qP3ePiliDB1T6vf9so18lwT
skb+i3jcTZSAeho8Jg7ohDYrcuju4c71x4LYZ9PYZiiI1bnkZuwHw7+UwjxnsTLJ1a5zspVACVHm
UvwrvY/q4VkMpq9GM8tlKXlxt4/Z7sI3SMVaJ+aVSIiMds3g6pHtAOzEXgUkVJ/2/Q8/cRD93Peg
yb9mGOVLdjzw9uEL6faPeKPxk62QUzpdLH/JkWFS4uFB3QlPEKTI60KyH1cLgsQMYO0vft+7HtCA
Iq+pHvpQR71MKXAAfNb4cSqhqxBn2PuZdUWhntpQMlNtFMXCoWYqMAkKeUBUV7qjbwiy1rVfWN8+
PRgwcqhIePtrAx/FU5cBngmXfSzZA6rsmDFpyHnqr2KUBXtV7NCDGdcu4GHVdMFodI4cF5a1Wt2g
gZ/5WY8MdXmkVmu9NyCHzeAixuLYV4vuymHC9tKbHdRZmLXsF78bEZF4Sxf6JLArlyMlJcTYGtxT
PvX5cTB4IJvXPbAxLFVb/nZFyK23rvT079akDH1YrEVIlDZL9HA42lOIvPE6V6W+s93ABoHE6TNa
x4dSRN/cW5N8+iJi38l+NnAF+4veBU3n6pf9sx4baglIja+nK6HD1rsVQLc+AocNRm/cQyiMEdDG
9jNFRDE00lUudvJHHxwbIas+sXSwq4+I7t9kvvoZPyflAN2DI2ei3BjM4U928a/it/nPjVUh7X88
v1K6lDKBHFOPDTXtXOeYhzBtgPpwQsSEXvTNnZhCtv/Jjy5G0ETbxdNC/rJBMXt9OFJsxQWzbxP9
6bIzBKEMHp92Z/SaoG0EsEcfe38LPZGfrsLwOmza4VNo5DFP6WZIIQCPMHXQxfb4x5W4VNxdfSN8
79jgDPZ7woLKdmx3J/CgYLJ2fObOBNUhHjXZDYgGQWDlmLPtK0QjitWAx7p4JXSZH0pxqTUREQQf
Jax7rdA3BRmtg0egfkPlTviI/W1xY3YG67VHyyZKUvK2hJxbrWBhhvjxNqL/PtKmYvnexY0qDI0m
eJhFj/ZyIiTOPLNxJW8Od1yp7ZWp3CcOuyEZ4ee6BMFljlF4JKzU1vYe5Oabnxs2BAi1/lyeBeRW
FjxzUMFwdF+v2KniNVVQsf5Z0lEstWHPVX70cm+MhkI2qfRVhpTgZ0sas5+HwnQI8IediCJ0W+xV
pgP8gHBW75jj5gsOaJNUozugGcwN/g3hWoeN+9zC9fzvJTwU9PvqSigwKg1ShuNLixUa9hXWywwr
rUvwOWHIS1utDa50DOeZ/JMQM/KvUBxZLb2AyoO3teQ+Ug550lXPFwddQfT/fgzITQA+s2yL533j
I4rHwodoZdj6Dl0vMEKx9da7su1Y81oPjqilgm1uD+2wFrgWD13+TptDQgCRCRZJeLHBa2XyMhzm
yh8hOFPw7nXiYYkFuj9m4MKBS2eAOZ0SU1EA5SZ5SY1yltoLr1HDvPP4LzJ+EWpc4E80VPfKWWgO
zwSF5BEBzUaqcxeZzKRFm7Qon1PeLQ9jxWEKGLDIeAnBx4vb+cKmSkuGOmD/UVUxfyYlReDB9BLX
Rn0/YomiEOxfHm1GNxBASgAk0DmAR7A03QcQQ+nOao8Z/CciivZsqbUX39EXA9mdEPn1y+1G0xXK
R561jMnDotFOChg2EsQVEj+XcQEAXWD/0+S46QyNCNyOdVbCCyWYaRA0PEz6vhOpt9liSEmnglZp
Yw6btZ1goQ58oyYORa50EdimKUjXYL8imXXMx2hwNe2p4nPMnEH4+rTpbixDiSYZhRPgAREXHK0Y
/iN1qVfPsk4us8PKPsM4L1Af/k7DpRukHsa4eu6uCTKVakAeqM1zasBxgYDY+9Aean912AgCp5hY
Tjifb2e6ThgT7ngzXwqgtSWy46JS9qhWBALwCnLbZrqRj89D6nqM9EXVN9wG2cSVrh29lsAobIpl
l3s4gub8PhZGxUC+HASxCa4Ubj01tpMCeun1mTvZOzLWG+QBwWcDDkqm3Nis93XeCccRrkbGNqRh
bJ5fWddnPtZ4ozSc0RReppUSgcI9a8cz/1k8RjfjaOVU22jGhwdVC5mGPlKtMI6PDY9/O7W1GWyp
/mIyQKsxQcepvHz/VV2cd0ndo5joSi8Gidpt/DPLULGhZoLaCwV9yAo9+3DrlG7w25iUGUO9iX7t
ajDxpTjk583LgaAj5SPb55uyf5jdp4I/EvSkUF6+FAWpsyC32Pa2HzCDSz7roETdcfv0AX3dgRUe
gi19sWXItjzQINPcLi21c3sNXpkw6ZWyZW/qSPEYLdkAgNC+lm4w3PeCU4+6EnkitKsY6KgJUXce
XZM6rjgRtZfklAnSnPf9zx8q0POZRXp6CEbhe53n/5LEBPgqjRJMrj6KAL7wU06wqghJNk0bcn+A
S6rJOG+KYMcT/zwAr4HWTi/p7paQ8BE8BQuVZxZX/qlqiPJ2OjoYx9bjYJUdFBoTI9j1bk70Ouon
XWe9u3FZu4TeZ7KWytApgDDz+tQTAJIZPI0NsWd0N4bascG8P85p9qgiRk3i9TzpgwU9Wyk343pD
tqR/a0Fx1pMtTe1CsS/2s22wLevHgBY5zACWTEN2fhuEw+LDUPMmEPUJa0as7SxO52Ggysr6Cpxf
Dm2QzXUfF7siarwyB9nBV3q3UZsEt2BAR9T/kXKHmNazC8EJYWBrdHulAwjXelKjBlWcoiY5UBpm
HkSAERuQDh3BjO0obMgJSGntPsX4Mr4aTHKos4BA/rkQRw98GIHiVaU8VDHKVyVgCPLKwMFzMKpC
3LqIWK44carG5KXgmHa3syrill6gayeyObwUVoX5F9qS/iWP9BgCCSG4fqioJwpw1HN25yxGus2v
k+P6vYJ2AggfEnAqfTFG8k+VNnXKCiecF8IFWbeEVLQaG4IouaqQlZ7wcG7B4C5CtJoMXI7oxL+B
lVQG1kJDnOOVnYwQkjerDfCe3RFkdCjOMQtbR/GsaxU7llMpCnP7i0/uIXBsiLqGn1rNtQUaFpO5
I0AoqeftJhZ+sMk+FglpAc899xkyX2nECZ2sYwv9mTe8MhF4NTbDkXrJpxB2AmTwn1MZHTreRJHt
1SHSC6BjIwCSLmwgZGlAmWXjPYrEhAV5yLe7g2Dviov0CFzOLN7m92UPMUfko7nxuF53OHLzAjrz
WZPEEJz+Zygcgo6jPDCNtu2Q00xEMGWjS0/m48VBcomy5KN/T2F5mb8jAn9+yB4PwWI455mi93oB
D+DyiDFeX/OkBLHV5M5KNaXSpCy6gkLxb54jt3qAuWH0J+SuT+A91nIZNE8rRJHK50ENNGb80qCO
lJOWyh0aCekySIobpRHvmJnX8gcoo3IzTIWH3v+P91YL7dlbuNs6xD3zuAiVrFPs8ZuUFlOd9kUz
fipORB/yu1SvMsj06J1M8GKFrM3hm3rs/VFzyj7ltUhbCrmXMjIWq7gR7R+z6bMabZ4ya7gWCfrW
A0iM/BBBjPbNrKWcTMAInKtUBSQCeDCKSlVV/0f6aIglD3qoimqM4PJm1WhkA2WEA35ObpQrwxGN
OVw2dtJxsXl2T83WoRILXXolOdiRMjdvpLQz/XgB+4CxQCVWmYGpXbLH3ZfG78uYxhGSqXC4VbXD
w8UltP9E+Op767xkpI5TppOs4+y7JaqSUvNSiBttP4y0145UFWkYBkgxJ1TJzPpBsWI7zF4qfOv5
LhxMpf5QiieqHWvfGgnDL+4gVn0ufh7VVKsS3n6BTVmQljLgK8MSvzCmrdM/sZdzvW5/8ZhtgoVG
ve5qy2Ejb7APgbYFb7l+O6wri6n68dOulNuFLQ2pXFQmpk5eB5pHGwFiBONpmQc/oSONa5zgbsDW
wc4+dytx7kCXr+6rA4QVkzTORkZn/Y3FIr62mgLEMmQnkkH5YTbZXohVppoPnwfGJC10SsyQRV/J
jykeZmGB9ac2utFdP31FyvgztvD5PbtMK2nZ0vdgX50iQ68tvX4sKOzkbb3temMc/6Cx6ZQTgoa3
f8Jhvza/zA1gbscFa8OPZBA4x+JbFAAnbn/HLr5p0GMNukCLL3DnTSYxLTTBBEosO0E3iU0ZaG8f
SMXRNeo8KyqxsW/oI4OIMQiF5Ghh1wdNw0ookMm+7qDw/KQwOwGG70ZOcgHmVTLiC12IuTB/mIq+
yaK9LX4mcRQJP7/xza/uSxjywn/2hBiyj7KgXPT+Kfsdsg5MocZn82K+66C8TW2Saw3pp6vzQO0J
IK6jZ4CgqxSPsHHyyhPdtb9Y+SCXojaDpbDVhcmhFh96chYHpl4YrlJHBOi9BY/U/SDrvozN9gLX
gFZnozBsCt7cbx2ghF07sDgQpKlLBUcBHEatIC/v6fD/yjanG9UDnUh/wdCGvQU0OCfsu8e+HJc0
kq7GXy3kd2b2xPG098qZ+UAxiXTI8tMOWHZxU01XIy0ikG0acz4nZlxzVXLCSC+vilN/a73UUlc4
p2RX/9rV4R/W7CLnIfEi+LWklYHKbSVHuI22n09kmOEK0pFvNb0DBs8WRav+iV8qP24KLwZNU81u
78leTqa87TWeavY/gT8eBDKgve3WVNqZsnTuAogS3+Iqh7bTllXExIYcvrtjt0EnuwI3vYoZO7jp
fnEVlVxwuTZtf1kil4W4CpNKK00tmBMjpNFnALpW/GGUfEulQUuvviLJmWa7E8ZGTQshtli5yImr
cZuP3luoqSnxWL6tyxEfC6pDb0PBI8ueehiLPlZ9q3r4JUKgoN2IpzoZ6NJs6ZV19spE5422zpxP
lg7omhI3WR7nXUqQemXuYpXXePDpdWHXf6a2cWpUqjRz49NLD+4nUAex/1wit0Zb3oUyXQ/8oOMV
SyNmF2UTgc5dOcYcaAiTxiYDdmi/+uw1Fi1Er6BIVe4xCF1HzNCCdmqGjoaayBudorY0shah2AVW
Kas/IBN/Jkk7+GCg/8R2dbxhTu69oxUKVB8VjhnPTVh20roOr2z+60OSAhIQKT3LHBn536hnZs5L
bqupXlg7M1vWIDZA8b0QSyMke++mJaG9qEWtXSWImimENWEq8+5m1k0TPnmksq2R1+dq0PTEmLqx
GNxIFDNQGMqraU6BRBj/nPwBSTKcf/1t78GL/QKqJNr3CmmjgdZV38K/K8BufFgc2wf9NCpcxxRL
xFTGsjH4M52Sq/hSsTEl5ytINM0O0Sp7ACb5yVNzuDVMY0o/AtAbdRer4TZ+Bs8VUK7Nca/nGpyt
izDnwhPglPy9BFypZxPwAnWFfMsUnqA9Dr/TjEO8jHnsmGdnB6XXHMYxd5BULPFih94o6NuSBL5l
uhIBs2q+Z0oLAWOVmHCs+bWKEGUVpS5DbpduIlMUEUrBjWvNe2pT38mKBEECcYd1vC0WtWrWH4JQ
ZUYRMszRF3UH/acVAU3UWgspGsaaaYeAjUsQmUIscCnhoifX97IHpsqMAFAITgATlcAq9d0t67vw
2aN8MLbp6VHR9N2osl5cf1Wc96N8Tl9xCsmujZb+DHyManCbbI5kjYr2L2OkDu+7OOjVHYMzAzzd
H5lBjkiFWusR5kG5bFKRcOvOepZ7DItts0RhVDYyJcMCDLa4BV4OiQdS4npyQgEeaW1IGPjgy56L
9syNA35kWEjxmotJNPXV9y9sGjLo4mmf8L3YRm7l5HIj2JbDIi+xkxatlcl6iLsu+rpGy2vw/T+B
QZVv/5AOsj+jO6SVmN8SulVSv9f/fcoEKw6RuVIdzMhvKbGd2vo956Nsgs7Df6JquPqWqzPFFWrn
QO9YkBwpcwJ3px1m6g/OxZhBByF0AQKo4UllCZIQplvPK8Jd9ci/oiRTu/HjlwDwovUbRnBhwVEz
XxOE9bJtMHUcq5wx2sKIajdoemABM+24mPepBsO9bevSQqptyDCF1GclFyBe6iBFxEV1xQjfntbl
TSLCih086LUSEIWu06pkX2PmFuMg6mewO2ElDOIcPnVLrBkq+QjgBLPHTKX/8gwNi+W1GLoEwthy
X0kKlvDTkbnBx3dez6/Q3Lz7wFqJcJmY0wsBgwlMvqqVBgtcEKJMZ2F60/46JrTOIVOUHsMm2nmQ
yImG+AzF1Q2k6uzE4gk45LjGGmQbCc+3/uwSMc9dl9iuuzvzyVM6ZcZXOqH/HUVDr4GIfsvWprbk
d6wU07uT2oMyKPVvtBQ6S2fI50035pFVYrmWtKami5eOZtC8emjgE/1cmsJf2/jmNysOXoD4mv+i
oTnn5vXinJtE3njpOhMzV2SjoOAzB1V+0V3kzKPuVdcOuEeTRE4EA37Iytd1W2gmqTT2a0ZWzggm
RRtrDzQyg17MTuzQa5zk+znypu8gOkWpRS+LPuX0zVjPQrhIkJAkLj3IBr7XJR4tr/ysdTo+qR9Y
+EdOf9BeWx6sWIvtNPijmGJbTMxRSCu3TZXOA/kpoO/GP5SRlHm8mOW07qXfN6gwRp5c1sRrC59n
bd+Sjcj7OYCOnfmCYIzEMExBE7L66RydEszRw91DmkEOw8ZXZDr0C/l5xk+Ei7DRQPPtsQP765Ig
w3v+Rju0wuFlTsM/p2L58SQd9wWkJSKnYnVJZbKs3+tJom5BFQeran320YN5PBRWX0V8eeL3gM18
qpB0ZbcVYqUWkkzlfFYZ9i52eaUVC6JsYcIo0t8205kANlX6rCeInui2i/FVyuAy3InRo2q3WY0W
Gm4pkQVaz3kgZq5puFz41/TnC75uJKwFuv879WwXCHiTvBqedjM9VkBmWg8STvwh6BjK7SXteG7Z
TwQhkNuKaoQzT3MnpG/kI/5nd3v85T8HKhr8l+w68YJEKhwTDuxRQgmHzb3A2klnyPUKSL5cJfQz
fLFaWV1KY/n82CK0nHl+AV/lFZzbPsyO/NUCQ0Ztbl8FcQWpK1YerqwGSig+YXRejiRI1gAIrbJv
E5VBoYHBOQXv5tR8YpU8iw/IKHItqdrpX6lNKYiN1Zhw852VRKCQbWWYkIxDcewLruIE27BVyZ1c
raifwkCLIexGmID3/fqY9x8Vzvx4g9yb4moFX689KXIMKwwoza4kt7BZk8w9jkrtdi+5w7ltN8sc
YZ4CKIn3+6OsJSk5sHlTTLM12gwTCpZcY4cGkkvkPLNiGLpGoSd+/t6HsXD6Is2t9gE9EJH3UorS
r/uPOrK5CV+CjneWmbbnhivY2wXZo8j+3djn25zqyci6XQMd5Igs/vWsbbFAGqNEJ+QovacG2Sx2
M6E6pguLyLmXWqZistck7do/CgF+DTxi/PSdg4QCQ7boEN3RHq+Ldm0XVydAZmh1YPjcGZLuygve
iLsEYiJnSEu6+FyByDLWjhre8OxDhaem5lQC54FC1K85SXDZpQxbzF3L8jXIKRa6BdNeEZ8Pv0aX
g3o9CsqnZ3Ut2avHaC9cW7ZWM2CeZf7iYqvF152Eclni+Zu8Jz6+a0wU36AQHcjnbNGWF0N/Z5z9
gRz5R10wmDRjKGgEVm15oDkrYpfdHa2Bs8je3VUHRzdOoysSJC1IX5DfGEA1fwotV34+MwrzNvTf
vcSJJNRkfKQ2CibDRr3IskpUsmw0ANisJWBh8eLfMDs0Ph8h0O7NQ7yK62BRGyzpvcc0Ups2kPPf
QHS4x7A9btwkni/Fet4BEQhpwW5Jo+tYwGXNrY0/lVbdvpYDxdGQ589Njbf1gfWRlkcJKQHZNj/O
y3hSDzBunTZdKVDMvXeBFzbzHIvDQ5TDrIe394obcWOqFW5r8qdviMat7ppZ975NI6jBhS5Xqo3p
zCjQvxtNsKwHWIN2DKNkL06Myp/9ntHDZofQcT1rTUC5vFuzna+iJsqUwEMdfKrEwsw785vVmeo/
2wSpw4NtRGBXUSgiUf4a72KauTNaIXc9kua/mTcr3okuwjJ0K5efuFPhhz4lLbolIgnR4vBh4hkp
pdB+DTI8HrFSe2YPUPEZ9E3KCqGWa796rVPnIV2oaYuy/4nV9fTM/YDECyc6ctcz1IeyCIRubosQ
mtPKN+8h6I1Dz5pG7VZWHfBtWR7hZSv00rhHAsCXuXojiYeMKZpiLtV5GltOIQKia7Lu2TBBfOOF
uOt/VJ+7eI6GrYHSqPOvsu8Kuv5om/WIdY3UUo61lC+FmqLr2Nr9cIqaZjT7nPGma86ARgTGLWdN
Kms6+qNedObQF3p9U6NhVDUaXC32M9WRzFIsDyKEB3lgOBvTQMnomDKbpNHzwy20WeqdOMWZyTfE
uDawdf6AedFkeP/hCM+yHiGp4/50RaP57xgveGdcxLJEY2EKGdItjhVClUdUZ1rM8IN9396161Fk
C0nm6jJgDjRS3NL7Zb0RSmQ6vAYUtFPeqPq0tcx0xzVpGGfMLZq7o7kJYc1tyAxB0pySSDku1oYk
Sw7CWCl5py24C0AIj7nYvdVjEVT77aFx2/NZUV77lzMv0EF8WIWhWLU+LozxR9gP1ASGckbKSXdN
d2Ravng/Jb3R+YHIWaKoey1GZmENPt3KEX4M3PtWsYThDaFYTCg+oUa0QEl3MX18HWyD0m7gfpdq
DraO3lefbbKU9nYjQMWS2neckIcmlJhsJjv5n0q2PMUJ9p2hRzYztMgYRzPk3G4YOpSNdEKuQL9f
JSovwMhfnhpnTogdRePDzynX2rwDnBKhcH4WXe9qGZ7xX/J+47YGAmdgqIFdB+eiH5Sy6DshxoQQ
Dh2Pnw+fWT0MMrtOICDfpzN7X3usXb+qNu1timRYz7itKlneie4FvtujjqlBHR9cjuFxQmLv5K0W
TuhdifDt2qNnR3Vn+2TQqasoRkZIsjE9mF0hV+Uf1kW9yTt3suTjNM7bjQz2MloMTSP8L8i67AAK
S0DOBLgVutYv/Js3jfMZYLMw1+wrVPT0JM2Bzjnqd2Okk3nmDM+j4doorBI+G6eX7l8kuaI/gTKN
vkDrsWwX/NYsWwgwgM+/D1Fja62glWKxuWZkT14TUcuHypp1FXG0vfdh2zVs7fCJIQgeU9yTbx9o
I5HBIqS9Y8o4M7PShqX37KGut/HzRBntKcgU8axZb+KCKMIssU55Xr8fTwAmR4/QeyXYBYm2KV2h
oIwUFpbITV0k4mL9g2aYD/WESbRJk0xy9ZZmujf2sX8Ost3u8qEmQUeQFMNGPpdgzB+JTAVAVXrv
gpJ+MHTbbsZvO0gUjw3WgUJWipeuhIaULoqbGn3QSRs5ZeImBO7hdHrEjSxZ+Y+To+imRxIw600v
A93r5HSe+G3qOLsT2CBzst7My/NOfToOh45QgQinCdto8cChMx+qJaQGfK53ECgmSKHS9oAty7Wi
An1detDBOQUMlYKOpF4U7o2abBbOrMUTdJuQcKQQ0erEHhu65yUFVO/3gtuGy+jmhwHWkngnDNJF
mDfMkLl1NAcNntmFvy8VE0zZML27Ty9ZO3yyvyUfoEy5YlHwkcuXQqs78Tu2q8NmenxeYzS/zkJX
aObOE5h3GWDMQY6X3JfzGiWMhIGmLWj1hVqX/2RfWr9YtzrjKoRMg1P958tYQ1X+DUOuVZBUjCjr
as3s+HLMdayx8hCeTT8MljqfUJLte+EDc94QRyV86pdEiZfhV2vvearPcFexwHiGgRft0RBy2YOD
x82F5hHK5yiygL2436+p18gHiqDvDqLzMi4q+qpvRuXhiOSoV8udubR71KD2s50OtU6horlzR7bt
47C0B6hAUSX6kMPqWT6trZoUuOTkGuDDy5vLFh6I92Kk91LPUGjsCh6dnf6vEpnnUz0ZQXL5sB1L
rNmJzvhNv2tAhn4oOQhGHiz1/AJ38A5OTFzPndRNITFCPnqfDlvoGU8qaCpHkJK/OHp1kvvrjNXO
YcLLHxpPm9iUS0EsM8ru6HHAXSVZMEazfOuPi7vqcAXzM1ac1zL1mvx5NAwQYGYkgD2urSbwYIl6
BvXmMfb6/bneYa/h/0LZSuIETF2SjOY9lYQBni3yAkpqbszimbvJUVprIQCUo26YuqWmzgkJ4IUe
LJm5vKTuHtwBfdeZCH4tZhVbjLEFkGq4jO+WSme8VrprUPH/LwKByGGH6FKVC08eDpFt3bkyJRX8
BF2kWEp/s+b1H4kTwRXDKZSEwd5L9JnD0wvpHjMWl0g5zDVkFWgqu/xoR4IeCoFleWNdrcgD0hMB
9vmdWAPhu0K0/+/mHreok/uqCMgS28KegoO1lYuoYfrK2FZxxWHWi2hyrPROl6ozLZtpcw1BRVhT
PDtHuIF1P7EG6hR/szCgQv+J8at6bijz1Kd0IpqqykBznjFRYRynWnVJ/UI35+67xxi1q/dVxVu6
p09vRmfbUVa/uTrfhPw6Bp7RyF2y1Ir68WQcb/qRh5EzanL9dkYA19ZAzv/dgSmzZF7iVsRHXpwT
Qf4PeNVYeB/9+FbRg+zyxdEhJQo8Uk1sV1R/sgxCdcxb33ezq/TtRc2iM/w3sAgat+owBteJObcV
SXKZt5wDgPWvGmvtYmh41IYP+vCsDzVecxSmsb/wQNu7MWLLVG8SEGJCDT90tjzDGEVyciouVwAx
KcgRVUbr8g0fT8Ap8o7/8xFrgEMxqPiEq/ZdlUQmcVpFPcFIyh8SqOMnAvzvABU6rowRM5V71tfJ
769BhRV4/A41JqLqLNJyVvHzhEV5JhyCWEGx0nU/LqGsmOwDmDHHW9RTNgIT6eG32S3gCUTNYtuY
UjB/edxmfkMHjKTQdYmXRMBKh8pn+JotvYE3zEPq/wQEDNZe/tqcXX6aH66CVt9jlOOorg4/XV6S
dZkDDumhuRbAbA7W6xLm8bddm78zFsQHMqVyCsovk6KCXvMCsZXmk+cfVasbi7Ay9LvJ5gsDMwbE
ZsIRRz4lKYNgAq9aDpiiAfkdXiBkhnHLp7X5xnS4sxymV990Rq6z9VB/8nMxeNTA4Niu5R9kapiv
tK0zES0hinqt4VTucENWkgurbQCwSt8bzI3NMeL/CrEI0TEgvinYA3ikhk1t4AsGG/muhGMzVS0i
cHpcSGWcCslSk5bIDb4L0I4MafLt/FqfjTDqVmT1DakPJ0wMLhawo2m5AvdjrxOCqNADig/R3cgS
0EjM6Ge5raGwIYS7kgcYLTNkXZZjM50Vc4SBpUz5bR7UzcNlJiAJwIoxjI13ART5x5mNX1mAv4gZ
9+Z20H3EvSSiD/jUdGfCMaLujnmsRM1LPcOFetg7wNUmkVxhB/dWhs1mHIcXkZEAWKmi1Di6djof
mZgDIAne2oOrxzPdl5X003XXc/uDUGttTFUpVTakrO3gRShnwf/6KkRHeitEMe2fz6x/JXsY03Sx
sSOpAg/7pT+uDZFNUxH1e9+FbcMDxjyrSb2wOXZnzAvuG3wMEePhvL3a4PyUMoB+FMzQ9DzXlgr8
Juj+d/8HtaRdkProKYHGoxG1WlF2DnKJEnuGNfCOQ/yvxjkreEKzS7d5nABpbw7VMCI4nsq34DWw
LzTzruECp8MyplgkREmLss6+8Bc35HO9HfJkV4NATeYWeCyqIs+IQJvlVG3DQ6+8qMI9NlRQ1Esl
ID0CJMjLfg4EYroALznZIw6xpmlm2+XaTuk64S4zFmEB7k3OZHTsj7ii6VR68R/v9YxImfsNkgJD
RmIUgnTmeBtkEN+9ziVoc0ps6Jln0v4XZAFnIR06crgLaQiiXtO/9L3k75aihyGnkq5yUNdVXy0H
3YiR1x1ynd23EYMcP6uM+0yGdv9x0LnfWeNby8h1kqDVdRyxLbdnmSOViH7WFocwN4JxfSTic9LZ
1L9eaZxCpWIZrwVjm1V7JIu3S4VLKlghVm98MhptZJaf9yVxtIbF60yzvBbsH0BOFVBdj/OXSzcW
kuvSeEn91aXsinS6gU80bOedX7zrxNZdcr+4vHLH5iqFyOkjhkRZkC6COpnckD+GxA5XxHck6BMJ
tMWwg7crX82kVnikJiyG4MtCb04PZlj9f7Vcgz1P1AD7qACtcnscowhyNY0b0LXrpUpgtTnoB1qC
y/L6WD1bkOfPwjwhNkuT9kEIID/fAteo9sEK5rWM2PO/csIlCKdBjVji3d2PTnWnU014JXFklR5s
LsGXgmfmQ+/Sts2Hru7zYPFrYwN5DSMnWDfJO5OSg+V3iXSlmz766mfxGLpEFGiJIS4P7EBtiXjw
ZgrxoWXAn2zJY8XocoyKhSAD6mk+ICUXwWvPA0vXlXdgYD/d5DA/BISQGq3LY2gT1VoxXFU0oNv8
SDQbsVegUDyQfdaIWektFAEalPneapx5YlZs9bdDVEdShrCDuCfkIZRDtKldbNfdanQpas8yDb/X
7HGouszz1t3drHgNSZiprCm8X0D4uhUt1T8QhaBPJxNYXjEzNz9aQCud+2nLRralRoVug/Dn9yoE
qvol1RrGYyLqwUf7hto6aLR0XWmlcaHKsKgzcJZZ1ym/ySwAM9CQarHu4ZcdICPB9BVA8zShMxVd
Noiph1lmDGOCCLgFsrlJ7LGDu0mDq1OZtIZoO7lfJPWgR+Ji2b9tLuiAe8R1exwPI+b5v3oip5N4
bBZb9xufuKAicDOTefNAJ1NhXEQM1lEwytJ6AVQ9Hzdj8iGyo/MNOBaS5cQz9zHK6QI2jFfHZ4ye
L60WKfiDNWE98skOA3h7EHC+PwtOwCMi8GTw2/bukV+TgWUlbgohN7CQTbAwIX4duzBhFLnE0Ig7
gLubXeY29gAjsiQj3nUVXkahjNWrfjNBxgEGZid8/hXUR4Wev0jxN9yhApjfXZuwPDpy3oMW/CrM
FBpMYRwuCdd/2qzvOjQsL1aFPaCG85Dr38ccMsraBXvU8RYa3cGGG4Y6eTD9X7nBqd+s5hw+kmjg
xB35PLzLxNLF0FIYgHjxR1YWDmWTaOZfLv2sGm4iBpWZ/LiqtgSDK1YzYEaKUSjHJfF/c44tU9Oq
gIwkZ8HCET6M04w3Bwt4UrQWx4mxDKCELGPPydUWUxJeKf6fz72SMa9vP3FF6QiO58qpmdPmtjVP
JFToDMLeY0+UuBvv8P+dqjk99VCTIXrdWXr7FgOy+jHdzMEseiBwnK+7KgtK3Hfs/5sg6ehKAWrZ
1qNypSGlyvxJvhYnlraNoaXamSTAHmRTVniKA2rJw+Ec0x7NH30qXWHEYXI0KSx7ZjsBc7+Wss4Q
g7+fJtPhr2F7prLsU2jAzrxpqGuNlLIR8H7jod9FEaISxebysehMGIevbkkYxyHxguKlClc4TsGn
cTaDl2M3IFQLNqwh2dxBSWOMpMTzXzQ5NNyWv46XIOafCgKPpJsLlweWV/22z7Rml9XulNyywwez
E7ET7RAd0m+kqDurjqiLk7wFIl9k+pOYi0DS0wcM4yfBTC/aTdcSIh7YDGz9gob9uAAgvNvF+MVF
5v5XvigKqQgxmkvA1QoeurlDwmxgqgu3Kzo8zFSDp80RGEVIFeFten5GgA1uzAHUoNLH+DN+MrRy
0cRzuiR+nwyM/pUO8SNRaHAhrfNgrAYZ2CgzXRdC2HrNE0/bTJiVlmIdkcEvbjUYH0479VX9MvnN
t7fP8EqjB/aEFCwlYZQsRs9i0iLPQ9IYLHJRVvAGh3NMjc8hLh9VgBikp5ajfjDbMYcyMGbzXZpp
AppPKBZgCcqqc/0Izy4MhtIMujMOKteL7Dnffdk4ccTV85fZgY0Gd1uq46At1KaO6I3WeciDAkBN
1NGELDbT8DryWa4+5lImykXLtZjoO7ZoL7l35bg1a7f8hxwydvPtD3tJKwAiCHC9Mbeb9pPAvNTm
DVh2IzZyuy1/4aRQeNmwW6y/NAPvNR1q/wQAOBN5s3o2jffK0EhJVvlXsKuvEV9j4vw2vkIRERAW
Q3ospOi/NCGjDSdY3GNzouZsWhrxt+QjuRK+N1/jtCzYCIGcG7/gdzMmGF9geELVITKxsMKXN7/g
HWuv5AWE3AQoeTTQOy7LJoEC6GuB+Fi1HmOSvQP5UQMo+ij7S9sYccQ+89E1gul98SK+0vpaXX7I
sjf+waqo1IQjBRZgCt2p2Eg/SjABsQXe3rJJmuDKBk87t+FAVlOwGSGN6SkzbxDrjN9QBzDeKjMR
M0J1nwdtDOQyu6OEyr4xcojh9VQ6sRb8YRQt5U0ztumj/I4ioqyCXR/O/1xaLSMiw5C/kLpHMNSd
HkOtLUc/kNF/8lhhW30TrQY3783eS90W3cfWTULvbsSfH65B5XAWj+tDs/dC22IzXs9Fbt+tL5dJ
0BxjXPMal0hUlelWrhDMwrctn3R7Cxs8XVeCkDvQV6j8HWuql3iLWLxesfO7wAfvdJLBJx+oyYsN
dyInXQNLcNhp4rfVwv3agmvB48zaOHyzEjLDPlHXQhjdNsoo/WAVOGJUHrKxK4x6oiwnSRH6q7YI
1TyOULWqXvnIRqYoV60JWiHkzN8gEvBfD28NjGf7s8i0J2DQ8xyNASad45coiLgTdQPD7WQb6pSj
TkF97m9nMKqVD8ZzVX0aqApvXbxMaGw/uCmoT8ZANimA8Wby7BzMnH86HD2nKQlSx0wWWhWoBNTg
vDVJXUWqgZ6bhYKy5y89OOzTeu5c7bGzt1z+gjyw4xNtPKCC3l9o4KO55jiQ3ihDyr4eGj2VGLn5
KuccyPmfe1u6hLKwHvmDxpGlKkSSzESDpOadRKhaX5DNK3Xb69N0x1apkfDGrrWJxKKwuD4zqgwT
0LtP1vkQBpKOIvFtnkJGYUPqlhvosLXwL6XQD4adWNUrR+Vu3HWRInMS8SwfrwrBqSQ/zD0xNmY+
xSrhxE3NdCJ3Nj3iH4RmyJ7CDPI3FzKfWrndBtUZUKO85VJ6Fqqg5mMWHvw+zAbOmikC4+0DXSwu
BojjV4MdxV20Q0r4xnz1fAGu21DL0Qv4Y5oSzCcWhIudrXx08WAn2um/O9NGLinbLvR9xidIHSAL
mCtKop6oxYaIHQQkLkrIcTJwqm4U2RxyfNPOEPJnGbyq/5SEyU9yXCXkME1ip3qEtFgA9TMr0bYp
abVVThjZi4tzbHLNJ5BptO89hIeW4JFQRD2ZEqaNAuWVk98d949xUAC3vpuOYC+c53SQD/s+E8+m
yZNLcjBCoTyhak5j/ylNjfpAiQ8sKNkvrauBdpRu1ZN1v0JCSR92NrsydXfO7U4WGHmI07ByjFMO
Zw/C454EQXKE7OS3msJqyTj/aCt1t8XZfp+vLGr+iHW1FZejiyvCIeHAejyzDUeApJsv9GwCCXte
DvwY6JFcHMv1D/XnJteAc4BoM8+a2ye5PaVyVWmbPGGQBAGd2CT8yg72OaOZzvtD3JPhjWBP6MIU
1CAkTUWEKYY4OS6rm8jsfB0cyQjIrdq9E7VPaiJf8Jk02AybMTQuy5dI/GGu24Q/5hLcwmeTN/0j
fJDsdIeuyJm4EYfGsupLMRBLEg/t8iv3vhiZbGumkmsM0ggbro4dLFv6u7cOAm469nKNt3WlmJsj
W1OzeFgK2S+HpJJzaIkWVfyhNlRivdibB+Q+IHIKDmEAuYNhP+8WTF3659NQTUqoVyE5nW3YjvtA
pliO/UZsbrC+3Es7ecOesCwv6kRWGcKAHyOVauhygBK9JZiwIqNLvsBaTZ4AhunUUFhukQFZEKic
7cuoJmmMRZJCsvCWzbN/s5XZFtKUmc/NVFXhm4VpmCqRG8mNmrJyyWHhCnJa86hm8/PpGSi8czzt
sLuQYCZyugZCVOGGHfYGKqHD5ObvnMJcWjWOBk+n7WhIb3EaZk/crYdNqz3yo4J9OqHUSbj5zzob
Z80XwJIkihwBTu/q8miOE4CrEbHjqShVpFrHDuv2VJwL25XmsoNpz8BzOlEDc12FARyvOD1tPrNa
W6chKrwY+wFw86ZXasgVuuG9XLwV/KvXrEENNPjFfspd+aTKq8Sfvu+uRXlZRwY//wcO69bzrE68
06+VYrfukqv6nMHEQ/XPB3iXBFuEdkdq5rqgI9CwmvPrGsZ/yTE9RfPK8nIB6oaOU6qtbxqkQc+s
dFHxEYhs8ee9CkKLBX/mmRrdIHF8bRo2r48DD883XvKtHq4Nl7Z7SFVViZuDju50uScEYquPFtG8
unM3L/+0o15SCvUmqc+IsmSJ0PNWNt4jvKIFXnI1oKAufC71zN83lFHmpyCVV2xiNP/tNZSZYGFn
pQ8toVwOAMnHmJCTzHGe4aULyeZLADAW29mfTtSMUpFL3SdSv+5Mjpe6d5hF+p0VvPHVXvDV1ow6
u09lanXWeSSz3ut7BkbG7Zswf9hTcqAldXsXtdXma8c513cIaLdwcLpP30PzLztpTZtp1PLVTl+7
SgdZKzt3L784qeNv1zXb9C/dcWumP/VIOPz49aa2jF99DgdZvxKMPH/xi4zEH2ghOMV/Jri9rYf8
qxqOWc9qDHw/zP/WdGG0oE7unxp9t6x4hkW0xhWPrP59PKYsHs8bClJBOiMwfHNE6FhhTRbTNVKP
1toe4pthqviPVWkaeDcn26wtxpdh3CjOZ7HpIFBshbxkdImCBl86GHAjHlTXhTXR2aJPQIlNUixt
YqAjmB96EwDtQprnk+Nu2QouZptf0W+SBiN3nf1CMPcL0vKdLdv7ss7tBEAP1cg9ahCI5exwtwDw
2xeYbGJ9h581iDnxYRrXbp1qRt3JNmXlXWruZAoX4goXzimyxFyp/mV201WUhfV/0GCBsTJguYWc
VJCROyIMJaGta0TJ3VHXVxV93BQm7k2evm3/cnk6UE1BYaOb38KhybZ/Er2CZttVRiQyO1IgeJun
GSq+3ip+R2j3QzcyKVRWcaP9MuRn9fIWz4H3heBxQzO3zIR9ZLZ6Pg+QitBDhXe/VypA4Ocjtne3
XCVntUwNmG7S3LqvMCyxqEx9dyB+B3JhhBujwPlXtZwsqkV1XiUL3c7t4kXMKeW5J+/Oxkb54l34
7Aokiu6VZ6zY4adxba1M/zaUwoY4B0iFTYENYYZ3LVfa32Ff3hQ9e0Dzfpi5nM9umqpoYoPkWmCJ
v/wJ9utacUTvH62BiM3lYCodetRtnVoYtS1VkHRv0KhBOh174eFNgTMRF5wlcT7GS9s00Uf721XB
nhfKBXCs4VceLtkKPQqN/W8A0dStd5xgaXN7LjhpxhTafIgcFoX398wQtfqxNrtAXKWIE1Vl5gpI
9HvXrRMK688br3kQhI+yU/eHSZMNM/f+ahEKhY5izXTfEgIl0+9QKT4Wbmlr0ufyU5DEh3ShP+sI
CdtOd7wlOKezGlnhQ2jpzgkjfiN3a3la9dF2+fXn+u19NwQZFoVdN0c4CLLDNDmRVogKC68kR6Lg
uQqOfVUJqi0/8vW0wrEF/wixOJrU0jGEW1xaN3XCgfGvdDSN+21wAbaQyxkobWe/U4TTY0eXJNCj
XlsTHHq0wxMQDvjFl2+fPK+Y0kLsQKOxlYJVjaGd/fy4Q0XykI6vBmYTdJ+mo/ygKcnMB5f0hQxE
peN/zP+E9ndnZs84K98rGFYJ+s+7FqT0VsTafYf4yVZHgg1nQlVvJB03Yu6BDLnw43t9yVHVCvZ0
gsR5q8a12RdIaw2/bzmI+Km/u/zGdaGxaRM0uXPOc+5zU2/X7dFbkVkr9LCtCTTrDAEryTcmyjGK
ZU/4Be4esTXVSXYn9rDkKylc44M9JKsrlPh4Ey0pavMOoI4sVpDSudCuyzF9GJ15WUaMpaKJdlRz
1UqdvBYyUW+yp1QMDpF9CkiK/kEvaQZ5U4n7EWIM7txWHumXhEyDGksmyaZtS0zDYKDxSwo69S2c
ssNqEN7V4M80A6LMjKZzE049llZtdWx8PnOJf1cfzvQRLjFUwsrjeEiV4pu/bdpqAoN9TPeBQYvC
MEUn4c59OK5zmzpaEw3F5GHWN0U1NE5inUp1Ch6WV41acOH9EjOc+H8KbFGCyT2dA1mdp12+XGLq
tMe4tyaBxGUR/7Ds5WwEqIu2bHo8ZUSJcUvOEUu8HaaPwxxsNuePpWZYfoOzhhN5TPTWepnfv+tn
BwY9/pnqDqVNejFhL4PyZKeNX06Rz1ve2d0xhO5yHR9cDd/7nycJU0VLHF39l5V2Hw0l+YUW01I+
Wpdw+vK/T+AW8nwAg/4gQDXpNJh+Angfc/6/9KizgSNOryAUotSu2NEaQKhNunuXSVaoBbmGhMn7
6EcGdlfiHJlXAonlKzhNg6ECwbLrISc+s6/m8kDDSk6PF9GIvEZi9t9MP2muqnNPnk0CzkspQPtc
3wDqkpHSi90e193ISjSVFhQj2QxxvD9DXzd1F7ESt3v0/B39H85jLr9iMSieIqqmtnX7ahbBtefn
cJlSCMkboPli9QhxgJxPYJnq1YPu7nwujI2EQDnHKcjSTfdxXPw+QJTfX48Dzqy2R+l2s2hd/5xM
4NzL4y6qicLXyoKxsuTT11ol5SNWi0Mc6/kfEPTOoDXXnX50tX2s6+SXj9aBuK9shnt3xF3V9bQI
AEeZzLQ3lkOs4RIwIwd70JPPuzntD7FX+rJR+qkQXVABTmEyJ5NrYjMmPpnixuXFcoYS0vRDfYrp
F65/Lo0PtPrYYQu3FENCIk5h8zfKAh2Ry2HBYBHpG3OvKN5ITFC7cuzv0d00e1C5DwxbYwli3ywx
+h6FIlQ42pBV9nQanssDGWYfVbde8Rf4d1jNqVyAblDyGKTQ14W5I8SneyqBPU1BslBsj7UaBi8C
PXHKZLBT2Lt+lGoWjv7MS5tMaDAbMfVvEX53/b6/QEiiTT6Re9cpuY4YMSCMXgH7Gc8AlzM4oOZ0
vtLD7HifAsU1TKRjRPPCr+NoY3Rkd2rLqlP3ScL9CeS1sD18rrjT7E60UJhO4sBdWsESAwhJOcmS
m4jPtMfgLWpOoENb8lNB+OkMV2lluiBXf/5y0JEqbzGFu4Tw+Eg1LDFAqVVptpIKS4UlpUqpM1xr
mN5SpCHdtd2yRHDQ/iNyoGbYzXNznVHnrNgmN33/HAI2X9nrTkeg5oi0mWgY8HvpVfgCW5p7tE0l
ZuMSknhW8h3evz0g1k/ONtQqMwNBPGWdDq7F9vvrsuzNrlGrgxjcMuPDunUXDmgFuQ4qfpIH4Siv
W0mA5pCdJYUCUlUqg++vlZTOFKKTUcR7b/S/7xtitSHQlQdN5S/aD2315uo0kCtMOEADNFJKjgGV
v/CDWFsbj6mzpR+/7NdzxByAhJaxVzvEIStnBmTn0gkn8Fqv2E7EbIH02OLehBKHLucvsrHpihjU
Tfs7RnfnT/f0mx+QBmKJV5J3yzN146oj7XgPCHx3GO+ieJ30kxH3N4HvCSZzSVGsqrS32v65dxmq
5qR1PgvfZG3i4hqjFG3GH4fyVhnQIkjyS4Hza6NXdb6VdkHvTN7qH57C8bpDbr2iv9ZPnF7Ae63Q
Sh94A/1Bj7sk9WlWVo3qkX8jamc0N9xeJOZ3OmzmwzP45NUlIW3VgKeCiTbGoS5Jb5TJi2/2ITDh
/WfKGE2E1jzF0WwgDVpPlixCLa4/a1GnufyAMp9neEKVjz1P4FfaRrSsDAbZ2ePy+wJt/CvXZz5d
XifFSX1c5oEcVf+TDmKllGRbbG2DcQa3OpMoAM9tRoVKGPNzkl7DRqCWkFUPByXx/YyrKKjAq6Mc
WjH3VfpRgO8KC4BeCpPQ8kffECEcz48SsamyolVTgwkO7Eya0E0Xxa2kmuuDgBO/ANXQSS701/vk
93m6EVhpFVl3Tz+TkM6S2tA2ynufAFjql66HmTjc0kvSG9Iw1MiXrH3/N2uZJNyEP0lx6YZUpD+7
7aMAyOgccmnkjeQuXgNF9pDQrGeNozXq+qvKXo/eDjXRw6ZcIdA8pBpDqvmfw3gewIwZKDDAoHvO
yuZcu1Wlu4p/y02IX2Y8w6L4ukdqkayBR6ElZqBnvNPebgSRYRU3E4tQI5O7Lu5i5StRhTxcr8au
y25Oi7O4whAaTKPMU1UmmzBXmE2VPKASZ3kkgOe70CDivRScCa6P/98qeTJ6xMCw+6R15Uysh7lh
94Yh8+Q9La5CR9OZT+OGO4i0G1oOwNP/hsiRKwa8cy4hTFN4HZDHLqS0URvKekldhhdEpvE/tdWq
W18uRWRPGzIGEn0XEqRmvI0zLMOrdb90dDQMYN/a16+uJ5oRzpqwqxMZTQDwGGZyTH7dwGnAf6A1
zHX+OZl2brWrDg6IyKB3Yr5UK/J3ADayWaMYuHoHglhy8k7K8p8tBlcY08nmS1E8zko/v0oOznej
GlMrTwidtq7vyC2mBqnoEOUaRnzGZhjNBJmq7ld0+pkRljuh7bFT1EUI7iWGArxiu/13B46s1O60
iQNont9he5Lo4V95wUNAAkv9mzU/0M1liHHKWzgf7asW9VbH51FSpNwn9KJ27MQlzJIdX7kMEzgo
Q5hlEhdN9d5M4pYeh/tdoJX3ClwIkAZ3blLBoAPtZhyQT1N5E7KM0sLZ0cXwf+PVpKmLuyWbSI1D
2X3Sxp1feWuzYSjjn5qdndSbP7yJS0Qn7tmDKThjDl9Ct6Z1VPevnOl/9ymgMZQ8HRcMzAhXsgHP
mAaosCWc/eOWFm4KxGkduLe928IOSFOmtIE0yf2lfXx4HYX7KJz98hfJMAmQmn+XQ5I0BGXMZglI
lO6TfMJNtG8G85eRyDYn4CHojJFErIlmmwRGxlIT0TvH28wX3iHsFqMiZfCxVqop1YLzKwMGzkks
usdnYKLog0NOijxcll1fnYR2vJkgfOkk5i9pdvLVGLVYciv0XxLlD6NVbiO3OMC/igP6k83nl6VX
7PEPOwZ2/K98u3nCDb7oyl2kOigDanOKSPI5g7WbkHPXoJ0I+RCG2d2k0yI4VDj85YA8EmVXNlj6
V3VUj7k5SUslT2Kr1Q5fkZ5cjK5rARrk29YOhVjSm8MV5dZasi/OwlYdHDitqiel0oHLZ7Gd3hWa
mHV9Ucb5yCwD5RcaHqhpVlg7C39P+yYdAC3R9BEBBj3aMp5s3shTv9QZN911EY7gQqmD3Vt00k5o
ZYv4KDcYAE59sr2Ac3J+0UpKK+xlXylPyUftWALPh4aAssD3vDaNDFCrD6icDEoLvv1JiTr5t/+6
oxK14IptXBGx+imgPNiIyOUtvPH80cRls9husrjzYzYDsMtO+MbhwKjcIl64TOqMCPAPjqtAleNr
72cXgVXkfIXxbwSFr/UkXKN+DgaNGoN6iRiqS5ZjDflWosMRC2Ki3KxfBXN1spNhH1GtUOiqReD2
vQF+TCxv8qPvu4uK6KXgw+CZpJNGi4iShGMSXZz4RMWZ+ot1BKCRWS5lL++afb1hNb1rECkpu0Mq
DMuZ05kLoY64xpbP/PB9TtJr9l2Wrz0ofVDo8RJpQqKQjNdvEF4tdCvTojX77pjq1hJjiHMTvoJ9
AX6rscSfvW/DvUMJYiWLlYMBy+gr+Ma6MZMcD1Fgmk3L2kHtXOQ5/iVPSwLV1olRPR/5MB3J/EEV
NfwN3V5xlt87F7V/zV3AioH9uNnDWNWUGDRaNDSFED5yuaq0ipOsw3yrH0n4P4x5cSOIWaek2RtP
Q9cpHF+IW8MTZ27g1HPjtks8LWUicVn7WE8hI9j8yiB0y5uyNXjrIFM55tu7WN7rLj4E+JQAyc80
6YDmgXpm22N8K5hJ7TJlK8S6q0Y6U16T7fcMluSWDMjw33XS+zOTq1CfCm5ksyfos2LatswuDXfI
cROv4U0efrSRAbF6ZTH/OPkp6fPO7P3fz0IQcPrQejV2SPkIQOM60va9kVEb5AOuRELKJnd1VLJT
WtNM1qxvuKeUwcndC8gAZywRmNLD1CbTjx0mbNmrlRzL3yvZVZKTYttBxVQhHJLMjL5HA8Uhxv8M
8hJBzfpp0C6iw1b8jOYFM6ZxR9L/IWgfVdDRCnX8Mr7i2hEZqhC1Z0EcjTEHd9UKRP2ExQ65HriJ
hxvekYRDSMLs3tQ1h+nwVeTKZEHRQWDvsaC1wDUEQgvVSFqeb4hCf8ElZx/4X2gUY29xq9rEP3GM
JvcCLb4K2aVxNKWJ8qcJPc2oTPN82pP5SCzG6IdAExiAtcDz20U9ugZp0tR39QI3JHSJQCjRf0gy
bGW62U/reB6NDw0iYVin9SZ3DCc6KhLEJAHjkuFv6gxpXUudbbiZ4Uq+YSwMRGJ5qdFRNSaFmfft
zWEdqjSmAAaYGiNb8eHDM0yhK2mStOw7Y5qcoPukhNCXqRicveZeHJpSTAdCKVFPzRxPKlW0qS+h
uNJRNQDjSTbAjOt+PR9PC1y4KiJf5plQ1eHAjewjoHDTDcDqgWtuVX83Tnq0viJu5ycqW4KVHn/s
3w25PzQaYqPUmiIFpJmMbO8uKsHoZlx0nKa6TROO21lVlTgqhNy4AJ5MYrullrFL+4Ym8DV+enIZ
+r6bZjFodTncwdlqvVvg6+xs+On7ikPbiOVp0m5Ed+v1XmKnNmTQBYPVkebjGgcsKnD155wojXlF
rTMet9FS4qSn2VhazRUb8XTSU6n0fgQ5HNXh0nKXINJE8EiCEzJz4UILXVP+eW1le+vP8ISpAKVu
aF4hxwttGM2D/qUz3p9xt9h+SXrI8aJF9iQsMaLYAZknA8xNgTP/+ZAram5jELtjZmt7p9fC8nPe
eZPat9X4iwhuZ4XovFO9HTj0i3b1EpaHX+W+MQg658xsOlhbcztLKMX663tHnQOcAkLmolMXb2Gx
vltE5/k0MbOFrzvXrvUNKZx6Dk+1UHpdIgFMUJ0hXtrv46aQkEM+Sb5IPV8N5UfdT5/CK3nNpJ11
W3sgj4CUEEyaxvaPWOyNozZzi1GCGY3DaqM32kwrhdkImmk028wLTL/ra9XJD8IiPi183xu3xOcL
Qy2lDEYmwiJNjakFVJVJYzWXWa7zGugmks0EO+fouKfsxVZPWXRFdhgXIchpOuBBCSX25CZKyX/J
IpbF0zaqxnhh93/GSuQXftrKF9iKifTojKfAVSF8AwHJOPb9jm/fPC5F0fDfXxNLSV+R19IXl4oy
gdDDOFpuMTYE7WVi9y3x+xF37dqNSBpr0OTq6BVi5d9hk6Pjm2vIEvPYTCxbCDrrOP4O+Ys8K1Ae
RGK9HhGRtIRXD4vqhnFNJ+ZTGDMKrmKwQAPZtbLgmEkfEz/pFY6+gF9YiB5p/yIKaZGY+5pVgmRr
0OsfbDXXOlYR5rxdLFvYQPbhNFTPrebxHv+bEX2OZKcZRoqq7GcMVnsp4oH7CeJMIeJIGUdP1VSn
lO+Pb7E7VCZDDEGwRhI/AvWZZXP4cxf0vRfHbUfAjPTw4EAwOnNWfpDrDueqwIu1y4ZNxicQF7Lx
wlzYwJ04jN4Kx+4chvP3RXE0561UzZZgCEN5+5UAkC83NcTGqqU61aBzbhaOJegr7EFbwOSoHXOT
659DEgUCU4XBlzy/UWaqr1enfREuU1nDR5iq4WCPN9coYZSQZ/r5QVqEZLG+8DEBCpy2BUmTaV0b
WK3sR5NGxa5ALRZAL/m7QSx55t2uk5z0a7qrbvjqfQuMlm80RUTlsYn+fQbN39Z9m3QD/oFbWQmN
Zb6+5jeg+znidFU6pK9re8zawaMx46M2V0iurnexvBd1bFZcMXB8D2RIBQvPRFfpCKp6ivkPaZMK
xjhj/7dRNYKJzDJfeZjXK3dEE4bE4l9q11RmoVASI6RaG73nzx4S3NUwYZFHqPWKElno69gGatfV
FbuI6jzKNE4E3sESkQZVgsZNwhoadq+N7bD0M4/7PrzK+aVL+R840U0vX1CZ1F+BN6DNiOvPS/0x
z2qjubrsrD7spxna2L7QnLPdM0+tVGR/BJziVx6tRyxbpoGfUnHF+IZ447W7qjxbvLr/1F6wjvU7
oy1twNsnLx+xE5wdCtO5pd+Fwbx6yg6x850PxiQGdWWpy2PmOV4j97eXG5w9Pjky52tmMl6ZbEug
xT+STmhAn70Wni5PsP2Cm3sCgJM556w0wh2NP7H/3m2GfrOJs21GRMQv/2c7WGMbcTtqUdcE6EYd
BpqdCNxVasZTUrP8r/tvW3qRBF92Wdxdd5jQA/LgTW/ibBBio3OaSJXdO881/9uRBUdAxPzxggCA
JcmHX590cJNLAd+ttDvyK0Chr1/id9tfjMuLKsF2mXLVkCl6b1v1NZ0Kn8/F+7OQfi1QHHHY1P+I
2+aARKqZNW4Rqu/kKZm8sUJSe86LS/+va6z7Z6sgXaWTePUdnDwe6UMKh7q/yo0M7jDlaBqw632x
gdtPb+ZkpQvNJLqHdeZ3tPayzXKexIUtX38+DqliJ3Vr74+meV2kda4px8n4VdizXYYpPNhXKxCL
gUBYLYvGcjl+n7S+LTEL/p0+AR7c+yxl30ZMqmZiuwkez9Relk7rKtL5jGFafM8WDkSFrVyd0QNI
SnWLYFXw8IJ8W0se6oAo8Hkv1/whVwMmBfPI4w68XEcCPMZGxJUs4e9LPhzGo4n9y6kEcoilyniJ
LlDOo/c/mUqEKislsoFIcxQqy5+w3Cmw/AhZg4+LLs7PT1ov/3kNrvX3J1xkmsQhX3OqvVvA/dPi
HH9vk6fDJQDHW2xESb2EQUhJARxffgf+CNvc3z/+hlJgpjODMCEIgg0g3fyWsB3AynEkvqawuDcS
JknGlrAmMmwnjSI0IUAG648pY3uEfdOStSVWawzQcs7zM10w4YXtrykoHC0PmiFWwuV7/5gFy84b
6umx0ugD8nufbdvC/rIJ335I610nLx+QmAF/QjrMsKeTG0Yxue3MI4Ft7lET1a6Vq+jHEOvRCujz
zjtNxd2orqhuZYcYQR7/dL84EZpRiPBPdcVzYzVH+xHc9dxdDonIC9lBwVSpt+ZpXAbSiuyaMlZD
wzGCP2QPwx/j2wEyjNvQdqtz7WeVkq1CfbTfE58nSBpe0i8X1wvypg+1nvSX63AXUHbtFHxq32Tn
JeGQe/4l1en1Dev2bePv6GvSwUvzkmX60+FyX3J5O6P26xeGrfrcT2aC3F/HtjC0lP2fYOK5V2Ok
vhXNLHDH/R3r1UCgxwHbzxr2l05k9vjmXg93A2eGywMZ1FoiExjo/qmWXlmpWfew9+fOZY5dnKj2
HWLf62LVPGXXbYvLiqqNeGvm9IE3vEUdzyT5XAOMFt30CafSaf4gs602+kPPPpHIDwl0rMnC0N63
yMdWWw9zeGcROBsQhY2CI5+tbGZLVqmCcqjomUVL42eUbihRv4uX+9RFSJsDTQlueuyGI3qCr5Kf
AqGPpJJIfWAn3ZkWPOo6sA0zOhGcbH7crFvPdiOzPcEWGy7XcmF6D1jTa8o2dNx9idcIWI0jmZ7G
ZFOtuIMoYSd+NJneAKy4C8rJzCfwlxwow+f571sccrPygVzPYd1rjYU0gAyj81IGiduUj0zF/MSI
JGMV5u2nXBNL0I6urMgfTv3cgjUbM7Xi6wVyp86/p5rsK0Aj7u6wrF/SCqs/mWckTrneA1De+9Fb
LvWega8MjhurXwubitV6sVonRknTWmSOM8OSZAbo7idM/adYmq2K6tdHnEQKu0P3h0ypKOVZGuKc
tA7nhb0TzYxp9NmvR8VRwNmE31uycwqM0GbXIV4vgaeTtsUI/wGMjg2sP0pFFpGhza/0ilMZOnWG
8xSWz7NUD2nDp4KmXrV6lpoWKdZr/NdaVtuvSPDqzBnmKsvwURD9kQacdD0K0xECqbaW609qVvs+
QU0D2zUvfge4USzhKWJujpXEw2gbN3N3CbHIoHth6YvQl+8OtY84yABIyGFf/YwcKVzcuPxzWuy1
CzQtiCa/kQxjwHpGMzNVJdyfjqAmMlNcCRSqDplAHDCCW4TPnW8EIVMdb6j1/luWjUoem2SwibYM
pJOupG5su6ZM9kO/+K22m4sj7TMQDA88bRFPX9AaAWpj80OYmDnI3nFMHDS3ZGMYW9lJyd+L+46o
8YygP7OZFJGcL8NPGMyKB74BCBmTfcpOzRTYSWnmdQhC6yQ2aHVRMVo+/eOa9P27Y13O7QXRypl3
X9zif4B7dc1y4qvkHbr9jH8VodZDpnNWwGSSgnnI0EuB3gFNnjMNOpmi+rvN9i3IeLi2NF+GPqnf
o6OtOzJQ6s2E9MzdOFX8SlsE/CVVratU+MhHHqF0qR6ONyEd4w68ajC+oCslGsChd0f7IUgdJQ7j
CPpzqbpHF1aGipt6sZZfObB/qKrnWLsHBbe4a+kdMnrXu+cl4T9owM3PhiORPcfbptnqRmtcXMOa
yCC30P/APSZ/51aw4UTm+rb3LUCII70IyoO6XZKa31vP+3IpmMmjErb1VL4E961lTo6iQxUnaXRn
GCfrQbecNpVa9tQoR4tVWJiMQt70f+jpv8+pdoeOfFkcheZRYgOMI2wklSRhzz61H/8F/YRMY4KS
EVCe1vsuszwtRYZ6lc6dYqRAyRiqlo+ABUcNZxRG//HGY4MJ75+mLQM3tI64PcX6zVzvNXBjpmr9
RfduD5I3vyPfX1avoXG6lrYS3KoH59GH9MCc85fQVZDKP37RtiseIZP48Gt7uBHtXU0p7LcFkau0
v3Jo2MvwgHI1+hpN4QEyuyhxqhKc+VsmPaETsPgRk2uJ6RHInATDrFOFo2uVMII/ZWCtrF60CNvf
z0mpS473GaAvozhOJRXY3ldDBmK8PWF9xHom9MMLkOpNHs5Qjt5yEZd4EfoGzPCCR3PPGpeQg9Qc
gcu072HV1zNjGISGN/RV1fdAFkl24BA3FhZ9pYo3ADBEAy+4DwBLc8WPhH8iI3Pwb8B9uQirR4YW
UOPu9pwTtvB+/hKqoNMw7kikiUzYDO8OUhC0OBXiLANyY7cGMO4u3LQDGS4Y9FHw4CQYUzK+Cd/d
AnjVmZaBmk+pIasJLty9n7H+96VRPnB0n8iqYI6o0tWEBh9YJGqRmz6eeS7DPZP04Tia1OOJkQHG
fum8cXExj6VNkJg8lI1z7iIeOo1+LH/+5IgqVQbRteN9ytCcbAhrEMvBTrHADwkAjniSf3U21l6J
yy1+ShMumchBbAv8A67u+jKWXPGz2UVbDFHGA43CZul5uoMktfbhYjy+dZHG2AbMR3ybYtCiMz9p
0yQzxXbu5ioc6+khx7zGY7l82PenshBtTtU3GLxP/YeZyRcHfdfSlx6Clj1fJxaiwdDftN9yME5P
ImrFKtbeRc9LYu9KXy0KqCDN0QjHAPL7hB3yHqD33ZSFDp3oDyZYY6Ee5lOeV2uiujMs2r0wAr19
5hwPoz73EuqaNsmTon0hPmM4bOxLIks+mArYJuwIJ4zhsPKx/XI1xSqlMFhzFFKQYy/4OGc3GjZN
nPm42ypkKZguQxWTAlcHFS5uauLgkjRjHW3NqNe6ls8Vjg9nNN+e5QkVPO1yCDAod73FZ7a4kc5B
1n2S9Q+3g2hCslvn7/+X4GBp6A1bUDbn1PEWo0MHYNzWBYF1DcNRjTydOc94HE07FpZyepPa1qit
A+dOxenn/Sp2t7sylSnh9wogW4xtJRlyq28vP/qvwMr8ao3rBg2XdsTnp+ofgpZBS2PfVyCHI54a
02j85mKbJjsCs2TW1HpyARbSq3gNuO3tO2BvZWhMLi8eMXBPuQJ4/kWbtW+HTEZBKuNaUIZsW1dp
GBwwDTU+VOObt2evxuJEYS/zX/PHNBoghOXopptOdWsKrGW/JurREyUzPZNDf0IJZkmRSI4yeRZd
/5hgkztMePSGuE7Ssx/aR3BKFtA9sLyF/B57UQZOuXrPe287JEBuRyd3CasWimHlivl31psbXFTL
PgyXv5p2K9JHpOUSLSN4cSgBwL7/rs/WkhK8l4P43t15oXV3OY+lCZov4J/tF5hSEkzyq5P9gSpA
lWzeRTPPmCw1KSfJKKiRYp9ZSMamIlmZPP8RjRWSSjJg9BUP/yoeSvlTHhhRrICt8nCw2a33OnwC
R9k6lWrWRayLAjIh5YXDcr1v7DZjKmPGRV80TV0+9/6oXYjItr6KOogMNaKuUdYfvio0JshgvKyJ
hYQTK+sHupML+lfLJ5Wh70ZYohwLGpQN5mPrpss71b7+gIOKXsZlUy//1rAjtxbuVo1nDmgtyP/5
bEE2R/3tPscGHPhUOXyUrseYmCXVfdTrTFnqkKQIoLdAqcK8fV1X2cI5dV2j8JHKOvod74Fjwzs2
XaXxyu53I8qjVwdb/uVVlXmHs7CJN8bum9PV2Y8vO7BVb9RJlh8zSzqIypcyaD1G7SvNTacA51sI
qkmPaNFrWpPwjfvRU4cc1BN5g2WetqOW4h6ufuZYbuy2OMnGXGu8vkPIBh38O548GCotCA1W0zXm
HSQPP8Y5YO09Ri3jsPI83MX935kjgLtcuOocnQobuvvBdkt+/xmRT0LEkczcueArM7BFYl4xgFXx
TrDYh8MnryC+6zX1AOQMxSbnlDAKEGdVO+EZ40LxymLK90Y9HUjkytX2eX7RFf4ZAyLCyY5pkK7d
mWkdkwrPP3G0JTHQpwe/Fb8jdsfotRHvIJE/s3lUU4N8cWX5hgS9bKmqW3uWTeFMS6ZZWfImp1Hr
vtBwF6oicZ91QERxPoK8NbrZjCcMLJi08541zatlLwhwHr5wdCpjRs9r3ZAHrx0DxkxIl89pDDVK
Asyckfy845JXKdqaUgmRUJcGtH/4DpXb5Ze3guzxXRFKLYoHUshfQ037hiDSJcUhDak6wWltjt6J
ZHZipiQVGXKnCQ2JnzdexXcHi385iJm/LOO5eFJI9UXeSOyVDkTkNLXxnjA/4LjdYNcND9PCyARb
YlZB0KcePOV6FQA67Xccrbt2gXHTDvP6QNkm2yYJlRrRZtWO89gdw8dfKRavoqmYmTufiGCY8ueA
K2Abz4ZyGlP+D9v6OhHnF0Z3OfM1axtieT7R/lKMh33i+P4f1lvueuOcqe2JYoU8iyMaLJ+73/OT
3fpdhNITEw3zirdUzBGRpVYHPGNRZcQhLHztwYCLvzbQuJio9rHHIO4t9SwTKep1zNhvTvPw+A77
RBG5bpgoIFl3c5P5d6ayH2nRFYxBvwIuaSgmTBJ1Y164feD84oDToaONmxTgzKi/M/h5N+FGhIYl
FiompaJGnu0eqc94rkN99Serdj33dDw2p5pWkMtyIiFDYVBTi8B/oAmMy4yTEah2sMe+Ih0Vtp/J
OBeOThJdEG19alcpU2tD+7mZOGAAGTfDG35uqDhY2XZtSZ8AKcvmObIGipGZFL5iF2aQOHAiQ16E
bg5O1SFQsJJoLsNwVbH+6RpcDSCas8eb+M1wE1AJCALd1lYcMcdAlXy8S7k+3IbSMdxjeaEokc6X
Y04mExHjrDYJHUmn7dX56Edxj4secc1jntQdHBuUFvWNJcUeU+m4EyfWelxXAXwoqxBBjbuHJkPD
O84YM+qO9uj0rIoUR4jjQxuvq89AAZYc7LMUS2tr4ABOEFVpWeO6zJ0x7p48vog+SzTheywDVsRI
s205WiaGxcwve497nldUTfOxUnFc0vceHLV3dnb1mY1WoL6hzuFM9d2AWLNAUxvv7sQGsOtIRoSx
y2KPYNAbNbEXTZAOihN8KnjxpMLone8jnQHQnmmtGamqneOZF+Xmjh139IhHI/xC1JS8zgsPo0mV
wrICTP/5F1ZF3L06BfYzCNoSPPeTG4ijr4+6Uh/kxd5Sw3mJaIzumKgUoANzh/j7DTZPHcRxMUli
MpFyb7xIBbxGEa889JzJ8/d0+HemnbmLg/+oKf5c4TcWhXzDRp9VlP4hNqd3/USt66T8+ICcgf2C
IrfaGl8WcnWlG693UmEuOnPMDRdFdr7IvwI6RwAgiWGjQQSXSJCsFkHBNAzb8N9LyykuCktNC/KO
MtmOLebmvxYnY63cEl1rwJpZ58L6T4L+zvlL4Hy6Btu+/qqbhMIHAfj+BRI7+1GFXnXHXUXaWPX5
jbRaxnhHPBiWwTtAu625v3vqtIOqSPFicqg+P7lJ2pRcegaF3xk9DjNJzI40SHGbj83PdmbzeIcn
yIR35IKqFGJr2DrMlJjVtY0sfSykuk2g2GhmDHBnFAsjupZnn0RQ6tDnwbc1hy18fXTIfDr15MBJ
oI0ehALNSiKkgMULIX/SzYWSNYj/whCopUkd7DbtRdRfvKjxBMyzlpTucwKJB2wBNKhmwtouH7OP
kmfhHgzzo2MwehOybuBF6lUB/9Yhg2x95oKG3BDzIgx2oKqOvprGRzUcPcdZRsj5UF6Qa37hjo0D
cRE/BWy35ZQI7CWLlXX0Rgswhk3weHLWk892m/5pYS6GYgG/KEVsi9tlV4Kmz1CY0AJIrOWjCYq2
FffiuAoEk9/jiD2efzQQVHKBi6yK35MBKSHDewcybUY/ejrNdhLd32Q8OjK1qzgEPKVD4YWJORwB
sELtdup0rL9+c3F9Pw8wflrCBBhnhmQEDfust4jRafOXQ12N0px6Ao10QtQ8ieCoa9prPU541wqu
kxc+VrWRO0WyOllAVY8Um3fsnPg1Ond8BBhrrEnqOmgWyPNxsq36oyV0P0FvJPen4aUa2uDCrkrx
FSfFKIzho1SDENNFUbryNkkEpf6SBBqNLUT4v/EM5bbYDpveFm+8y1lhJx4mj+i6WT63P7JTIPAR
2UGDqDLq8snQPbR43Z9gejF67nQ6gU/VKfDoy8lamRTq1kuPf6AXfH5pvHuA5xp7DQIrAigFkEsW
jDd2rgbYb5oSd9zQP8QEinUrW8OFEghX5xwUTDwYOxGDkKlorL9mNcm48ObzD1j+kGxr/ghlgMfp
4kZo5+qCJXDajHKs4G/nW11yAOVI/tqnmMkf22W9NojK5ig9PjmWbmjjdc3a0qn/kkWV44sfvsqT
yu3bQo5dQ5mU5y2ZyTi7lzIDhRw1FrRYQBNJQDh75HNuUT1QD6Xr7rS3AEQy1CxBobxSEYEGsmn4
0fI1Mcr3ZP/UYL62AMEnFQtJRNt3S1Ve/I7Xs64Z+DiUPnwKxjAsMCcoa52jqPFGK31VtCTsx9Nv
PCrHdjt7MA2yDYtDp2s44f2BFEy0QOOxSVwyRuYZU7jhnUJBwGfwbOTUfA2pTFRQMmUbqdJV3IJn
9iRamo6FH9FI4O/+Z0TzNCPMPcz3A/Br61bpugllGcCnZmTJPaVuARSoPSIAZPSuMeeCEFAzTaX9
FZK/Uu9i2vFpDuZgtIwegIeUBX4kfl5r1a/Z3Gg9THSOAI6qGHo3oVzy56145lMeBLU2eYfKJ9Sj
y1JP5L7bClPoYAbdmMZVCFDYoKmxfRwppnz5J0mBjq192uBAS3Y0XdBlHyeEYEoYhfjei/SoDb9C
CaR1zZN1lvhqJLdVc6dQNR5/HH9aZGNRwf3859v4YGFSlsp2aJXemLa5joOmbeHqSwzHDh0ie0ua
bZzp97ZmeRx/80PPaQm+FoBNgpumjGp5lb16Y8qd2pYF5GdFonrOsXyc4GfmVt5gTPd7b6LZQxGi
XjN+NsQNKoKbTCmedlcj5f+2A8DCvtD1Ag8onB1Y6Bjlp7YTp7p6b3fTiIZsnk21YS1f+rlw1qWJ
ESGaPQGLA3rBeDPOKlvKiDmpkYrv9T+5MfU9EmqYKip5+l4RqzACavbuzzucVh+qs8X3wm+VOBet
oFmty3SU8zDWCYHOsBfSzM+/rMlZ0sB1K71WyhBsMtYvE9+Nzanf3xcc4Q71PXdsd+HwwcF/IX6Q
uUxCAwdBD6SA7kQJdb1Ec2/y+5CUflYTFh8slPm0/qTQa9vKfx4L7LCrcNMbBD1x+cxkrM74uVz7
1BYIo0VAOuSzqE6kTw+30QgDJYDr6QUGQdHBoHXQ7dL2xDsgy/JiMnqfnMPJqN9Eia3tiUjOOWYo
R1jbQOuA5vTmu2LSqTm4IyZxydw9/TqfYuzFIAmOIEblS+tav+jQb3hVrR1OJXIWiy3uQpAm6SHF
St36iocqmLkF4zYx1psUXCyHD3wW+ktxtnywcxCanH8PQDD/PXI8UARPbZ/a9ti+SQRMt2Z6ouwA
xELIJq6cUESuUmceX1ToojQ7WyphdmqDA2ggkiDafXJQ4RMGK8iIF+Vd3Z1Y6Au0L43YvaQ2UQbQ
UMBEPlfdFlyVK9Hw/B4SQ0ic8T2Bjt5WNPmWKqE5Y1pn13H+8clJ/qbA/TWhIJkeTEbs2Jpx6hgi
peaQJGqdW/9i3TExteKcDzlMivmCuwjw7EVtNEbd6h5kaihra5Yy921KA5I1Ixr9hHcwSZWn3XQ3
TUiKRd3S5s3vEs3WijPTNp617HegutmY+w/8szKX0pKjG0WVi+fNc6z3Hqj7Txje2md2+YdCfesp
Bq954OYnPItfijgudryikFmWW6R1Ucnmf4PzVeCNDDNhW7vlq7vPoLxGP+UoiKjMh4rOs/oYofvP
bTrV2/wpkTYeJ3zBQnA9kVIxqVvR/cgOTOKJ/S7LzvZznVaQ8ah9/dZIZnewqVDjDvKlCixYTpHt
I3c4FwBCAARPaf8hUfPj+06pShBZWcVS3iccItAFoonWz0O6jmdwdku00FyMd4acjSCIgui1wJF2
/EP21Av8eeQ2sWTwKHJ/yL1TQpzvMhYK6+HLzIosFg8pNk5PTVIqHU7djImXgmauCE2s5rN7qDvx
Oo3OaIHK2BoYdZsVngMx2JYlvrkg2RKzdtP2QTdd9Ebc3/1cpVgzYW+T4/MZ/KGxWzL9ouOCS66J
U0CkIBcljtTaTsa5u/d28R29HFlFia0wF9LuvV1F94hzxTViCV3kqc7sb8VUUbljohZzXQNkNhlG
2/+IIpWx9DIKDOddt76eLcr1AaHtDi22nuhGkQpB/LZZcQJM/iqvfCI4esZK7uh4+ESWbvlKjlxN
b+E71aw45XkcQ9TfYrqZZ42fsKLfaBgVca1F5F787uFmWPwChga/3l25wGfGo5VxPMVyAi+7Ve5y
IMr+dWXlO+B5YZiRihjEW4BIBd3deR8lOEcvd4bAiAg9t5f/ebDTICE/l1kZ3kBgU/1hmBxMhYWG
D88upxUStGdsmeNw/17RRuyB59jZBjq6qGXlED+taKk9JB0hu+vR2D2MLdRsNXl3RQgV3q1WhyU0
uUeF7dGd/qx0o+KFLnIJIwicLjOGDa7SgwowKId5t70/mCmDsT/v/Nb79IYJ6fTR+Fhr8btACYDd
PrTbR6N7+kzQaFdvzSj0cX/nlLQQSm+8f+ZuQDWwtahfKWq+XQWdHhViTfdL4v+6AeVscTzmq6Bg
iSFvAfoOfeIViv0/NPhpGDrbt77LswOL4fEf/DhZXmebk0Ze/WL3GffSyG34QYcE/C4eHKAMieVd
YrIqNnUTCyzgai8OqD5CZ256DzAlVYNJUgJ+aYlApPr75HUag/NLb9VseF6pAu4J++Fz6XuJkcqC
YvWkqyBH0BZdMWlodU1Xzz7U1ALTcn5Bz99ApocbhJxXdHYk7aXfnyB04KNFoxeKmfqQxqtNmaG9
GDEHTuIw08GgZdeLj0gmWWjmumdQac0mSPLFZTGe0QYyeB+QEqK+6OW5BcAIPLLU91ZLhAU7+/o3
bvARMLgjZ4wxPln+eFsBtZCyvrGXu6ytPpJuSXqqlL1xvr3me0ixHT9E0OhaNw2Jq6veTplwIdZ+
KTrz/V++6DgEgavsi+Nn7fPASXIufgXzQSsSXupBtMMir4+usoo16YXs/83wFUMhaXL53S7JbrXs
ft5BcPVYOcTC2bhOvazj3EuR7xgJMtAFjiCcQOJHN4c/yvIeFYnRKQvpeOkpfjS2cDJ8k5Ljyzlr
tNNM2H2lxOdbWu7t2vLhT3sbGvwMD0TM6V88z0UKqsNJ6d6u26oqOvs314YG1Do2l9ICCYeKTnun
pwpaGIGZOuJ4yd3Q5p+7lxs/WGyVKroOG9nkfGtaZ+O1iw3G7OBIyLIByiD4g2BoDg8lqzhIVnzE
9YQ9QRWaITRJNIvqxmVFvU4TRW7Kc+6psyhWb/OvkwYQ/SL/2NVtFySwosmeUlhP4rq+w3YV8jLC
yjWIpRL7QB4G+yvTfvleVIyltlU9Awd3UZOk6iANEHOR0gIO3mKEi8xiI+5UTdkwUEkPoZ4mRl8V
2Hq6bVRym+sYKxIFisvkvwGxear+ke0h7L4p6Ddl871wW68g+tFwDLr1mgUSp6GqVEaEhCUT0C2F
MDIOWj3DvwswMGkHdwYPLIAMnkBHOMpg16lJo1bjF+42ApwL7HIFMUpwpPlUvlxWtjDjFpP7MdQ/
aUgAjmsafmBtSd+HgSf0c7AOTarCkG3oAeWyQNszZSXslCDpahXKeC66RWI5PEiGvdphe12lfz8i
gr6k2njxuPLop59TWpj/E0kdSHNrYhJA4URzhnkYLpcr6o6aLb/n7nu2/Z2TwI40Y5LRIE8VwHlA
uyZ+38T6hv89STeuIVs03mYFrZcn6X1NXlLPAtadeVzRUV1GaXKDPY1mF/OorW2FGop+fVmnifE1
rvkFUcLhxDJK3gPIqQZoiEhLl23TNdqAEd4H1+E8RpmWCsSKHprs5crtA0iwB5dgfNXYIfW50jTN
F3qgn+TJYwMKeHHZbj4tP73V8dNZvFVxK1TyG5qhRAusbF7sEjPBODvDLr9R0ctntNPGe870pEDn
K2fPXhiHVnoLZug8W0kncvgx+Sq8RjfLlsuzmHljEe7QYq8TrSn2SabxNZRR1TsTPWhv+TaZ32eW
P56rHys0X6AKXysPFvBq1/rE4HFidLLgdKEAB34/Nrpz2/cs4l8lSHgzSraSRCHUrc3OPmOMKKhi
P8NaOH7+NiyiLkH0oI4hVtB3urcAjVKrUlY1K1XUGegSTt90MEurMYsqOWZDOIMGHiN2qDwSWHEd
++jYhzcXd9tN0x94gocTUwA/U7p/YHxMVJ28cuWQwQLICPutJdt1/GSH7BsuBqdaOTcTVyNlq6lR
eml4AvBD6KJHnIVPn+oY5s1+GHL0BrZQw0GAN6TJ74+p33cT9d5/N+imbws5NDVEzeI6w0iMZZsN
avEj4LxVRYxI5ESwHLtPl+fRYbkCNvH/7bsgNj0c3JB2C0pJHUZn6d3YDvOtCvdE3iU0M3bx0JIP
E2IPfxtxU34OSX8KKIpIGSAEKyRLLKz40twt5Roximnb0lR3OdLmHLhiiUHAX9S9AHfkgwU71EmW
Bkq1uuqM6xCXqwLMbocFUA6j/U0G/RjUPQ8OZi0j7FqOHVl+Bkaz1aGiUcYV5XmZMFwkTJFi4uJr
jK7qs9rg8tZq4Udttz9yWsAGUjrTPp4K6mL//P1lW5DkEIuW0HhDWmC4d6lfEowYEzKat8bbiidc
KQly11ISvxeALkMBDEa9b6NS2FgqLFWriIvZeMRkj7+zhkBfcvObyvP848Wl+tH6kby/6/LxBtkE
I1lNGVuYRsZ/UYUO9mIDK8rTtEYPIXsVCgWAoFEULxbws2tPBmbtaImRnz88/jxIKE5eGAJczAP9
NLnuC2dlRzk/+mpk0bMqOnMyN3bysBPktmzAwzaTmr4+7zw8fYiSq/F81jDoNr9i/7gFyyFspEII
Rw/NAVuIM90FHDFpEsGdqXhKoKPmtLrEes5nxhWOBy1nFMEHkB5iSQXUJsAezagxReY45OvVZSmn
o+49hCwPHjWBKK+c+unrUYTISKfm6SiiUs9hyuc5qmKYY4QT1sgFty4CUNWmL92keY0arIM8BLmS
JRofw3mNATap+1plYu9Ptlm4feet2cFVJ+nXpnoB6JQ3Ky3JpCTscim3bRomZQ/pnBRk2BZBU5KW
0PqM7kW6GM/oME3PZsgPr1TDagODBaBnWiKOgffmsBtc4PpfM1m/4/uJgbaxXH6tHyT8n7y0ugh8
NQSwbwnv5skhwq7Jh3d6vrVcw4rx3lu+OPBFA386px3TSkhCHo9RcJlZ3La1wX8mhu/ejUrI7tEU
L3x5VEjBOX5SqIjdb66XPL4B7F/dOjB511g0s+tV+6WoNoql7hmQsZOdSCXY8WGeBPQqDDdqCM8I
69R9j79d4kWzYp2JKCtPNa5PXi+9B12WCSPLVwjmUuoBCIDf0rsUOLz7zPGJgudbZoTGUAmcQUPZ
kr1sPCk72xe0NpnKPZ9GQMZP2R7yvWsuOeNu10j03Jgzs11s4KNrc+jwspQeibPBGuJCv1YTQfBN
/fGgTnjgIvQWe0O3x2GaLmd83YCRt0jMLJ8C1oDZVlH78td54206dfizXCTB1KzIE20qBYobJeUL
6KZm29qqhCTR4psqBs6rxs1z+8ZJ/ySYW0xNqrTt5k8Rcz5VDlO9g1nI0uWCPpvdXMNnzYRDsX9j
wocE+sEIAKrQeeTNUeEOt6a9RDGyu7QuAJp3aEDEhsZNYv2xZHVP4oaxJdMK3KbtNzuQzqkYSOZN
ot5hLZtGjCaijeHdJnSAul5qcG2oYWka1qPg3FSCnkfh5/4lwrngh+qxUzPkUDF//SKhQYz4cpx8
wVSzHsLg18e4nuZtG35m0RS9ywsskQO0OzG2oDn/6mpVa26WqNa6Y66YoUUQKOZ8H9LMCTsFqzDe
zC2h7zYnwkndCbik4BXeHm3y9PJFt9rnuKsezzZWd7NWlnSFD5bWr+s/InRYMP1NvMhCuIAYyp6Q
7DSkiXH1JEqUEjQVb5K73StjUmjvc9Z/tePVo3eQi0TahiRIXpjVzr2AWbuSJCAgDmXvg/0BM0m2
UqrzU88gJuwo+4qBq+z94t/yJPS5wNvuwlaK4jc439swzIxmOOfm1Nx8+OWZI1j8oVqPK3Bsg1yg
x5YDr4CQKvbiLbGdLeyTS3f5GJqf77GIf7TEjYSHPQurJWitrovY/jrfsWhOUREk140lCVOJyyRL
ulzw6mWKKNTk9U58rWhZcOWRT1Ft1YZVU1bdpuGRulSeagX1H+9vmyTT4hkX305SwkkGCJxzFRl2
vU4qm5qfmjKfFb2/wUTLKm1kahQvQvhXjttWVaYwe6Eh6fdlkZfESs02uO00e2YyRq4DgEqihGuf
3kO7X6dMkrp2ZU94q0sTkvygsUwvv1Bn826q5MdnUnKNGEWGVjlUyNGZO3wGpxJDTivtYv6XM+Wa
EhbbNrMkp3cyHc0wIndBJrEpSf1BmqdI7KrH7Uz8t0a6lYLTtw1QevnqvFDZJi91jjoG3CffL25W
MnkyKwYopqHuEzQChFE1bPVWYcDGp3vbYbVTyMtjdpEf0I8r8OIFIjlwiqZQ73TF5nWjzpwzt+Aw
K/5h58f/qjlsMgHGAfzMnQp+4WSNNTplIjLvwC3HhutjT3Qk9CFjNBmAoefJGZoprlH97RUBELyQ
dZ6ah7CzH/GmMyY0MaAp00/JUOFecRjRq0WMtF8MWRIp/svXasrQY33OYmEvxCjICF8w3Z/vr23r
YtuqFo7blIdsOCdo0LaBZrpTJcl4OZIRyRQmyJrmLHfsoEwccMTbwhyULybFHoYMS5lAsbg9QKJx
pRVdOil9ODI6pMqPrSYT7FsAT9NafLjZGRAs8hBTGfH+16X5zP1a8bq/FQOd824DyJuc5jQqG5+K
KxEjPM3Ss4qkM7PukAFlw7kp9Ad0UFsNQZLRr7Rbg4QG5hygC+6BqQ5WH8ss6zK7BDCyhJHEHIzP
kGSR4AXOcWFVEHSmZ9bk+Sh7+GUhacSZWxb+300jgC5G/JN30pDqbisghjm0RIFNSmbihDAeVeE2
OiBv1OcRIeRpAIWcuG4Rdo5zmpe1FAb2dpZdDYol6pRr9Cff6Smbf+WPXDkNzxH/XvDIctsB6DLI
DiktwynSN27BrsDagrEgQXzxd94UjUHOEh9M42lkHGXOC2PC3Nxsv00LCnjm9DrJWI/FpK8nCXbE
g9dASeQB7QtOLf68G1C0xnHHD/IUNLhNsSgD3pDBWk3qqFC+atJOk+Y7esEMuovx7PzDyv0TVKa3
neyweS+9nZPguTR0km4fzxwkduZGZVa/RP6l0l3KA35w2zCyD4R1dGFmIZv6NJ6phEcwnkExCPNI
kILKG7JGhqmKKkRrpt8PJ0Iwx2qSkAXEgflCHoTr3gGH79xzfIuPPURN80VHMfp/+23nZq0Sdhuo
TDiFfxAk4QjdjqniTxyVXG6Y7UHNrXMYkyKePY1LM2hS4gqjQgy6kI8BisQuQ4CAFNIK03U9suUN
PHRT6s35+k2fcIg2nZ2prG0ierSfQGaT82SlfNiXy+8KxFMtJ6ecOkAfhQyWSX0jGHW41nqFY2q2
eWe/WTS5b8c1P4M7p/NZYLyH805PQBqHpO/3c7EKuBrQtH5R2ozaGqzy3iFeMPvhmljc150Uv+Vg
E6Ukj2MXQV1RA5tM35BgfcL4462c7w6VVzpGq6Hd+WZ7W2X6Dw7Dlxx4dtaHQeEYxBNbNieXjMF3
J5rTGVxydQ1+8HpbQn+Ik5jyUBqcQKhF6dyc5OV+nbyeHh8/YJQnzVII/V5NOH+9PmznVaoMvaW4
Lh5KXQMy4G6AxxIcCcJzxu8Lu4SmVEZjpAbe0vPdy1aJ+y0cIEBPukuAhYl842sIW51AYYqw7Eo4
lVF1JVtfit2MNVhqxVmlCU8/1n9uakiSn4dFr/YNxjTGbI3SiDuzIhpe96ouu/e/IowzzRrEoue1
cxOuN6znNjewaI54yf3WTm3xB/3UcsUZ7j6pOORqOBLTxKG+3FUS62g4cpX7NfXJOOScA9ytmFy4
XMtIV3Y+VMnhICBmfb6dtaUl8tg9qsBQ33hdmvN9SHVJeDKv3MqiAbXGvA98dHP7FvzvGRcJZ0nc
Es8fyZEduvNAupL9G1dwI4JNRtaBXnnxU+qBxA8UC7sYnngTmaNPrDbNRSuzEzLYa374rg+GpF83
mAcOu5KQK/CvxnzE7yAgDlh2QN9NUHgM/wGb6mpX3MZHQZKzOy3c9If4r6OmPaSVEOwxzdnuEMYY
U+NWP1e3tguZOnApV8ZMutVM1iPH9QLwcJh+Y/e1FV1WuVEHYYjLMH2xrwRcZBIW/jKh/pmBFfYC
J/6hrkejgTeBGeGbnZmFjxqE5YBJYU8YKj6luxk6/V1cSkwwi0moR7I9C3xgmBMEijYxW94GYQUf
beCu7AqBtnZHifRnXFV+uVEeiZP7CNLjG/zYGb6X4qZtqkI9VUR7mUm9Yv3Emsl9mtxPZRY0uX1S
mE2+DZQ0mnd99xw09s7FczIByLMSHlan0/SBiwT6w62DsyySrmlYIUeZvgCSRkWW02S+FIzZSEZ4
eydsRPJtI1imjZtAuqp7rlbvgdsoMOszoHkoOufoDZcQVkFJRt+92h6ufKFa2kUr8WcwY2CeqNBE
/S0oDfVyWqsgzMTSOWNNjKE0Y6bio+IBpMbj7D2NAhnrQmgyPcopYRAqdprMDpjV2AETfjbXhPUq
Au+zA5f5Z+72uLFm1Vn23D06K+6t584g2wgEaYAMpA0WzhsAug7dOMlxp47JCGyNxaUbwaNVA7pF
wg/QsCmeLIRsL7hVwd9Cm6aftHLP3H+4YPPBc1DiTwDJsZPJepKPuGvLdSY6n80ruEVV/JlCXs4g
ZSJEvRaRubo0n8aIehygSJqVc11mHZNxSWWqCElr+hZepqQBHj8bejbmvrIWhhP3fkFmu9aQDjsj
dyBxuZHUdgn24B/4ws+5yFgMbC8WXiZzfVRb2fD2PFF5mv6Zf1vNWqinKpDyR/08hoCShZx99FPP
HQhx107XVXcHzC8i8sBii0Xx59Fpytyuquimj2+ejmhRlpj6CglZB8kiCJhMon1eY+dEEpkjeytR
CiJQOATaPpDFlN2U6i3ES0ouEjEqpKtR4qJiD0FZiDQP0ICfElRXflztex3wCHNMbJNkl3RvoCHd
IbNW050lJniRiwpibxo/acnAiSQW4RhyFNbYVvDosAWZWWaEGQzQlpZgujqAHzTx+HDqHwdOjin3
rBwH+7VZb3pOh78d6CKipihbUGcxB9Yw0xG8lGxM8QxCpn63v+b3/WA2m3dORwYN+1S7uQuNXh59
nhX6H3e50fjKmpjHQ7Lf0Z/G/y6RkvBQ8N48pWPX/1XJ2LGFrwz2zzBUp037gGdJ8rtteWpKXEb/
yPf6cVXPZMjUGWfV2cTtgJ5xvcf2H/8X6WXLxbQ3RR/M1ToZx267w43ZB4PvrnZkUKPvbcMP+fs+
ODe0XhEeTeb6XM8b2E4CdnXhB/JIrcg13ueqklOuHFgqXcyM3fs+nAmO0sZBu0X+FH1u9LtM2+Ok
Xm3fINKmHPimqDGwgN9gqA6ul2+UAV3Ly4Ao0ZjJN5PrF3IA6pX9S0paBoV3N+UxqExNGQUYA5Pn
yf9XSERwcvm2RPZ7MYa5xu01uj/iqNn2q6GMv2sFD9sMr8btdXkghtiqgxLJ/j8oAGUnvJVuwpuD
cvxF7UAysABApsnFqdCV3PIcnwxR2rD/42w7qqVy8J/svZzpl5VtOV6QEJhGQWyITnPYQzqNZHO5
uaXo1IDiwjyebtUmLKe+a1bkU9Pg+3MwgvJFgsH+Da9vtNik454FgRPjhRvZeOFj4Q+MzmMpnR5D
rdVgpPMCYYJrOOAscpAQp5T6Asd1gRGPaWig2TiGSuGnnkHTmngDfrdfNriqycByZmAan3P1eVXQ
sn1YDfexfVMFf2QVMMYcfEmWQsaE0ZpDtfF6a6thJ+EDPPTkFmddvBPztX0MgLRjcbkUGyRiMtbi
Xrx/6sZNASR+AbIzZGu1uduj26qZEpNo6Sf2qK/zENNwOR1FdEglzSIB+BzPB1NMa/52SMBQCAe/
EvfyoPge4hts8LaRYauOi4z7hGcmGLP8jP4gFEoEzq/XDbk1GIflx5BSW5Weyoh8X7FofUqW7K5J
EI4d5KhmTLRszXncPlCTFOJVUF+4cCbEb0ctVjPCcV5vlkREGz1fIgX9hU9PsMBpWK8vX06Xv/cF
WiHKRDhXEL4bU9rqscEpn6nr1hSyD+AwmSf9gHiz6W3zdzqMkj667pXPboP0ygt3CGTeb9W7wLzg
WrjFcC3I71iOWduD7qz35f6SMDnWSb6YlG7w3vvMoMdKV7op6mx9BW0DfLNq1yzl/9TbpNcp8tIp
MCj0e0OwvNGH6WYilWX/1IiBTBo04sTcQZp/WB4s8c9s49tA/+FlS/X3nfi+RZ3LAaC1P+LBCrcA
3RzBsWwNmQgkNwS7jkPePHN2gGN0Hsz/NWaCkC3c2ZW0acOCWb2dUvF3MpEUzbGFcD/3xXiaP0Zu
vlUzh6oSZCqrUiX7Tnp0vL/qNy0pZqZMZQR3uhbpbSAapr2Z/qXtXMcpRHAjm4jab9ydXPZuvFZp
t3hNue4+AcsqUmXnNKGRg5BkpodfUoypvD2hW1LFWHFGJjUa8YWAT67QbZmRK+wmQ7n05vekmq7z
dvhl41x+rE6aXJlZDCTomr8/IANRd1wCs1qkH8zIBNJ039Iwnl6/aAz6UuglbBD23NO2v92EhkRf
wq7QGsxbc5pJq8MOGybMRbLXaYNKuAJV46UJ14BAkB5TkrAD1xzKHMrQ2m3c8uYSZMxlVyY/COtP
/8A8twDhoAmnYScTNylj5oN3xjOpN1oeO3KaOs/bcZEygBcGbFuwux90ghkukI4i+8M6Dgj3Jc1x
NX8DA3y4BKgnDyCYiru92/fVlDx4j2c58fgcvbxUgSOQJTjdbczoYAbApJaseNP9vgqeulscZKse
WQck/G/v93ouG787ccNI2cp4egLRYPNHBfmQS5omhv9AXrlhUrKgGs2jz7Frywm1INq2LzDPNMZ7
GT849a7CX71/VxbePf2ivq8rMvYd1pn/SnOCYtlT46jxRQ6Mz42b2DwvwDFKQ1JurQoodFlRfjBI
ME8V5j9zB54VsCHQUEt4oLNuuTiS1OjKwIgj4OOgM8SCifSDVoRpCXJQ+w5AXLjvC+LoiKJZuWdC
s70LrLlVAkuxZiibWuWwU2JpQxgxU1afDTM3QGH74Prc4CKzmEfwNUi8YpPDCXbv+v0tFH9qlIqi
wTaeqMLxounYbS1wdJhlfnIT5OaQHbais4+VqjB7wzxitpyY2jrlfd3X0C4DkzHTwgMi9asc9+S2
YoD2D9xvjXC3BasRm2MP2KvrY41S7AdQo5Ba3mfIuHXiovQPdg+CiTYyjRm9ijVg4HeCU8LAiRV4
UAX7fib2U5W0PUkHRwGRtYz8aB/PXXTAoIQoFoZa8epLatoagdZWk5+J/rVko+j4FQUnfoFna+zk
gnTwe2p2uQr69TLNBcrVtfB9OJ4TIR5/UQaVtDypAxhPD3N7csuoeopHrRAmrv8CATP2tSFTweHB
WMtOw0DJaHLIcCTY54LUfvRZzXQcwtPT7o0ejxyOly4pJKuQGE+f51KvSrKmngCKTZ77d4/Slm5M
Ux9CabRE82RapoTURSxxicajceC9tXwnJAxHQLp2Ch7eH3qR0DXppsrCb4G9Db2YWCle+oCZoJdh
N8JgY11YVtsy/F6NCbilehu9R2fkvRJr6xnjCd1uZoCqIoqVkWTuK2Swwysai9rjyVajtXeao2RR
ewjcoRGsIT0IPFB2nRCjt6/FyrXRzhvDPQ0Mw6fUL1C6hQXiq2YUtYHGmt0nWqZHsboyff+So4Q0
KcPNRahMlIxIJicuS6aq44CT7y7iFmKAedCUMhJQpDeBezfX0bBreyczLV0tPraCpOnstSJljSkP
76OyXudgvjS8W3yfMrbk4K96SRRtB5P7qYw9RjFK3SikoFCMbH1YnyvwytoW4LMqzdFsrF/yIr6h
DEKqmT7KpUnhxNfSZgpto6OAo2AaLIxT0CeOiKpXKK+w94sjomV7E/SRlsKnuhYDuE9a8WR3gFEX
Hp7Yd0boI5fgGIVaGaSrC1wf8nl8yNpkGLBmAY/s2iDhUeBS6jOQBfcK0Cn7Sys6hiVnX9TioHqk
/39WjJGuHtOq5unr9cQC84BY8rwTafkIJcRKbt4POVpeNCnXLUpugmlHNID0aKnqqyF+/aSYXVPn
g2712nsqac7IObD6z/ymwFSuasL/FZTGCmck/fdbtfimWEGb4fXly/wefMnT0bJVhiSqHEpcxLRY
tJKz6q4/In2pdbXfUcZgNWx9FPqlkTT6rXVQ5Nb1Z53hkDqBmOH2SkCqwjrBYKlPJPJ+rAoj+oub
EeIY9TAIhbGZx4tL1FeVTD61elShPby2c7/LxOcDMYynXsZDXnzn3siWikStokGc4udbriN+7PYZ
aqMFPvCo+nNFk756rXuruQ84EKAj5hkOe0vhpVZboFh5ex5SYi2kb3L2ZGe053ylC407ef8H540b
la7EX2FML6bgh83d2TRmYk04gTf7lSmDmRTZgOyZS1zJd5H3zlRv6/Rc/meiaW4WzRcAUQ03Hmvh
krJWsIip4zyO+LmPNz3/mkl/CN6fzRDj8viPTs5jnMFrwiCbZR5802toWDnJn2p7Hx+NKyxT2SAJ
1xrGm92y25MSFEXP7CINt6eoOIhHnOLyWGSKxgnf0Gk6iQNX1LIPQJLUtgiVEdtubFazZwYKLCxI
mq6XaTwTfPcuhSZnEIWSHjCxPk54i8sE9oIqUavZJnmUWmhqKZ8ilk17AM89Yo87s+xZvp/YgE5s
2GZR4dIJrgUTtIQyPZ0gSbQ0ClN3xbSzVfhGaaLgDAsLZYYaj8J9Cl6E05JgJPGdZpbIbsJfcs1y
BcwpZ0bb68FCsLyXfwMEXRe2Z8uIsEHNjGsS7NXmtc92jBlZMjF1TI9FBmUrhbyBr+RlYaMOU6HM
rrrvaeEvur5fHpN7apIn/znSGiAimqHcvjMRgoYqm7/hto/v8puCuJl/6x2+RBpbGo/IhxOjfgfq
ftKGA4/cKvYCCvQSVu9BQw00q+KRGxUF8UssHXUSKGD9wOp6tD2VkWv4OEbD3S21gSnpNcFSOA1g
ocoX/Jj/lMOTVnn6gFlIqY+kZMETXFZHGGu8LkVDioPbOOjZmBFyaEKUV5XAUwCWMi5yMmWplhu6
3XSX4141fRV/ClDDHUgyP+KuZAsP3ikiehFEZ6US3Nen5H6NiarWgytE8YRgpqNquHaOu8sJ4ziE
7l1mjN37041cI75yz+dQgCXXEjRngzl2d3LUyCrSrIUTzBCgpSW7gurt7rRcL6xGSnMDbpfTflbW
tsHzUSOOu/DFiRDJ0syuAvnBOkApY3Mf1fVVQJi4vhPYHvGDwvHkzGFAIiseDysNsOr7nBFTCo2f
MJSq5eefd476oVYmV7dfYRZ5xkDmGM8I9WgKNhWn1JZO1OKsdpEdFhT/5/JkghD8tglXrf0TxCGL
/nz6nrV4FlslqAQ1h1XB7FKwN8B2oJgO9lq6vryCbU6PX03SOIrauDkke5iUDs3VCl3uvtfoXQiv
LQKkK5WeGojQQzLs31b9oBimsN4F0gS+OD3DYvZgx8mdTdSZBtDOhlDIo0c3EhKRCWvye1PPuXL7
LweRZd7fVy2jvqQcZKTmlVXPUak7ASczlhas0L07F2Jc4kiPwYlEWzLqdEUPCxwq0EB3rIyxw3re
KrBcOdOpWWe3MD9UxPvnF1PFy8LXlmvI7wnXhrxyIphdJJrLNTuomRq785h/nzLXPm53ys8N9wzM
4aLHbLDUMJ3SdskOLuBqAWam8dkgCAnqAJVkaUbnFvE+bsh2Q615JbuN6E4iVX3GdiqHcFnYQcV7
40f3I604i6083suT96fqazG8evXwTVHNhJjJXfqNKRoUadSEtKzs7QpWQSL9ua07IWfpE1dwA+p1
li+ESUrtivEQETu+t2dtCPJ7MjmPr+pK96FysFDi9NozaMmHVCgCnGs3JH8fdRaaWN7P5UrD2suG
elxJQoNstF/Bmc6TSwQEjftzkM9I03Ijskch00kjAgqZ1Gc2nOcDG545KCO+P6P4vP+IsjmQxvnV
oIKOX4rZ5SN3BnPp0Pfu2rctIBfCRIC/T7mNEU/4wCpQxRwcVQL/mwZi/fAMKy1VbebiWFJ02yKS
7ce4fEfN6gXE9l09rHvB9OCIK8+DKTigA8nG9GnWC1BF+LBsmU66obUvr4GJv9upTGHYYOIOCcN6
rBEx1YK7ezaTS8bCCLbV1V1c8h9hiNh6U08kFTRPOVtzGad+bvNv2HOdUO2n28bTrMI875V//v7o
qCfiOnKCIPmPhgnM+dbRqS0iNDAfQCrS+cwjgxtJIAL3gL6jJizPw8LQz5tlAVnrD8hQcZX9qzIF
a6BE1f4SzKoIEApr/90g+ZRsj3Jo9MBSX75IKT9V0B/WYsfMzPbmil8QoBkVQCscT+g96I0SA/hA
dACXSJCfioJLCZkfttHPZsmn/nWN/3ARhHz28dCsKpKmrata19auC8RgaWdCoxC95ZQJ5YLiC8m2
1ahrP9v5aSSuI/OFClYGTcmK+NJvvpP+QnFC4Vaz1fuM/n9eVokdKLG3iRHaUsFYGzQlNiZRVQvR
Rp02r/Qj1jDLlP1kHQRsOPQwCO6mmo6KwQbLjiwRy6Hm+i0xQqti8J9ua3JozLsfaP2GRkpHSPCc
QIzMzF/O3m0hRqFzo1uV/lni71dMxlyAzQeMkod8M1Q0Q4LMdKtyWfAyHWXyf/X6nb4650efMh3s
WV2HVqxVEl73QZk/aIeqh38mrmSfqycR8ELpDV6Yf9+mXMrd8beODGAUjJKcp3hzw6CDX0XjY2ej
XoYTDOKcntFTdiolFJie5dRXBbbGlfkLk9vh1mAJqepNu+ukuGdjqIjIB7mubBBLEEJmz6wIuvys
CenMdmcR+9F/a+HqX23wBX24GI3ygzqInWHx5Bd+3iHZ3oIlv4LMHu2SNUwerqji1AMdADMidXig
XKhCvZURXUg6bh9QTS212Q4nxNIcQNBrr6a9SKGiIyhFa1EI21UO3SK4O8P9Ma6p85KEzuygS9qS
VaWcDiFVjkAU+fawRgtVs4Fsg6DwOwviMuDTS04bBoKUz/mmhD7nbrGUFAFA71IIhBCCCKP4UvBA
sbOpDIimt08tPb4NQTYQE1O20ZIhZs8MLsLuUXbtgiXa/farHKZ43IdagYuj9Su/SyiXuqUet32h
jNiDplGr5wsyXINjKAejPMdq0OSaSTID6Xb0fu7NX631kIPbkq0x30FAKMFAMLeQxPwo54erABkA
n8VNkuUdmQJXT4OLVc+Gvspbn0tXGhFD8QKN7tijYRyBxCbKKrykwmt1Uxx2bWqvUZPJu8GAGhdL
LJsM7Ci+41qcTRzeFqDbj9JQyHeGGB4/52Dbr1IzjEaioKbk/6zZtXZs+VZWsDob4dw992zIBByB
1K5ksPfmm+lJwn4icJoR8GCXh2aNKLEtrvTOF8vTaWgPyCVXQVDyeCjT3xwdwFXwbrqqgrXTVBin
ZSSfFIik6q/PBuy3tlTy3ELXVu7KugH9xJwWdNo5fdOu1KuRJa4GSeSCrAxqkzKXksYYNbZ6bLcB
T7tvP+rgR0QX7z9NZC2ICFphp0JTdneiDTMDBmggk5CWtF1YHyxq8cheuNNTkNf779xxdKm2vnBH
Y6y75mN3R5VjP6LqHx/ZW2kchvBs2ou4exbDForI+4zyJi99awPV2DhsCEqcSMI0F92twk76Vq++
6yjfSbAIR6C/Z7VncinX69Aat4D+R4/ii/dyWob/FuuoiRUytU5jFUimluwO3xqxjVQp6wiTgKuY
znyzRLXYfqJ3Mnq6liT5JXaRM/RhIrHNyhFgCizaogwj7RdAYA4SGTGvn6KWXqsS9FffobMwQvCe
P9wb5VlchpcaVKnUaI+CQygzKL1kCeQG0AO/VKYyI7EbgrJoeDec36ctHqYFM9Mq59j8dHRKLOle
yGQ71pp+MVUstwmqiOKh45ucxvm9q5zapSm1+FRJsgs5R7xSBHjMb7q81rDYYVxoo4skgAZPQszM
Bc30jVS1XZ2KCD1rpoqdbxQR4+uE/Z27UXy68/NXoFYozpvzoCc95H0gwTlVt/kKBV2nEb1gvEoG
Wuc+8094eelKIcQLfgscKQ3vqXHwaeQoQKmIQ8llGyQc8QGij3hK5A1dwsMpOozpr7pTah+xYCu5
V+4/ulCxo1TVgKk8+tmx5sgnCt//3OOjmICsSexJHDElN3LepLU2/etB6hLIKP4Q94nLowf6Omnz
SwVvrsv/HTEY6n1kkcEcfPgYqzkDcRTDRRUQKtlTXoh+rQ7XLDlBxIFXGZFS1c61kOM2wRc5ZE7Q
34E+q1y0PY88Le7DlJoE+/3r+ZfNlwrCWjWU0paHmvWrIpRmazz31XbrH7XlcA7Xxg2v4TlNixCh
YVi52WLkW5FI0f5t19lJx9kFELpB5IJwqLL5eHgDYdiV5KJwYz/FycuzEGEVaZdBjdZe7MoOO8rI
41lfKRVrmHSJZvX0+BS2PMraohf2nTcHpgF6JCvYHO5+fVvr+fAwMrZKz9Ck25D+lEoOvF0vfc23
RHA2q1RIlFWYHLs0FVRFzzKjT7tXdXl9FDCq0rmQ8yBjRjtTY3i+RJQ+RBC90IGRYBgFATOAiSLI
I5z2U617z6+NNIjfz8lhe/qXdE/7dGo/kPT1gOwFMzJCJV7t3DHi7qzhppAa7Ry9J0ANTiLO+pKH
on4sNiQI0Da6ti0yccLig5GS8wbZtux55xMafZg1058qqV+KZO89SM1wFQLBOorfEPxNtMGZZ2FI
60KKt3WgMBVfVT8trkqDoEknYWWQPvH6v72yfh0R4tzcPnTsv4YoQaTBxMbuTa868Gl6DydUB+OP
+gTKWEs2FSgiKkU5moJOeIzxUPgKMmErDTEF7t8L3VyXCbV6tjYx1OXbcP+SYSIQrLJ62YIUsJQR
pz1mqsP3w/NuFrkJnT5/bU2VPevh8lX9qnXq7s+oS5ntQxF9iAYkEAcpYlszBIQkzHd4kEYhJ3fh
oeun+SfykrYDCwLxs7t0fCEZqy6KhExm870vhgxFxskYGMc++w3Uw8XuQ7R0+kaL8TRoouiDpxUF
g9U8Pja7DKzU7nW9a/Pqu39V1O/uvyBC3m/TjdaBbgK3k8ftmnT11AETpiRqVIc0+eVoMt9xdHL3
2TS53YrQJdqwpdRgefHqN7iYbVTgOxyNcnUgq1E1xzV3JSuswAf84HhbldsU0T2EpHIUvbjaa7H9
A+4FsaV+/FkTwI0lAlfvK6lZ2cQEe3psmY07TxLXDb+dvN3y2jg9/jSnKPGElsjxyI8e41eoZLlQ
A4Eu91V3yKsWvSOuUiHGyBNSsabcQ8S1qSS85DDjQUZa1vioy6XdE/vHG0CSQn8ewzoFO1hYTUsS
Kniom1mjaH72uU4saTDqqHqkSskJvi8WUNW8DqusdoER0ToiOS67KP/Hzm6FeyjxFLseXnQtl2Bl
L/s3JhPOGHBEr8LvnKVW+TLtF1ccfny6JIge1Ja/VwbrX7+7lz5O/hsFKgqCe79BLePASH06oH/f
UBTVEQg+bprpALe7zDYbbxvuoYrtoyjmGwz797cqDfz/Q83y11Rhf5cxYWzWE/E84ORW+mWCzfCG
pkUQPcAa+lFXry1aOH3jbtWhepSCfxudSL/mZGAYasZXwYMTlQD2lk/ZukJv5281y5M0mtgpFVs8
7DGblO8VkHffQ4BzQTmrcTNX1N+5Y4/gBrCBGs0KQeWRyRO9aJEaZZy0O02QUBQscieH9x9Lo010
7r2pQuY8S8AMafu9u2ZwaAf1PmRXc33j7VAv40dot0jyzmLUROMBud4w5XQ0ZIwjJu87mgQBR3M9
dpYqiOsCztlhaXpBrMoAWCjl+1Z/M4yZrbWMW7R1r8S52a9KBWi0KGbIOa4Tc3J1m7zL4PUrGVAe
7nsBN9rh9kDbcKLWEuU0o/49iPLp7iQH6QVoEgQeE1PWkGn7RAPqxXgy0alNWkCgezy6tfKjnifz
11yivn8oAPEAzfI6OelJ2olvLqCb/9tsG0HB9gZlBf8X6F2DyFEdNjnaWYD6L0MmCYZZQWUg3Sd+
UAxn9Z6dCabhw7nq8r0JfPixa0dcATv++XfEyeVwW7x80w1xTjKR3szmxzHGrM5YQ2X6Pwl8zAKy
FYSDsAgfJsYfJ2pxBr0bmBIKRYbEUUWvDk0P7YQnESZh0gMdl5vAhYWcoLWvnQWA1njNBRGPGjBm
4OQMEv728WwfI2Pw556LTzt8MpYuTbySec0IuDao1ndQntEWaa0uHYOvVHLYrBFSWjlUOTGrIJkw
8pgC2k8PtX/xo5VWjo4SCB5Ycqr7A3EDRXNQONQS8wf5f1T1PSK+HJUUhM4W5+gRlPlp8QltCCX5
x8vF++Q06Z9KCku1Q+JHWehcshGvrR+gorO78/wfqpbHFeddAHAzhaGSZQ4dndwNJDqDubKolWnT
xwBcHuRpyhsuXT/6OeDzTgD0PpMzqIlvpcrtRfYlU/iwkDZqNWpaLYSDADYU29MZWNyC4kknW79b
W5LQZAYrhtNDbOfE2/4tn7edbgGQyhg+ZEhEJXf8n3W/AMn44WXr5S7hO8eGp/mZQaoBYCG1mYJb
wL4K01gdtEDYtfFBClIOrDYLOuqC9fvo12Xw+oNYPxetdz0H9gFjHJgeouHO/6t/Szd229vjeNB1
9obhjPCVubtNND/2boP02u1yNX/RgWT1t/E97jXn9KoBqUdE30j87EfDsR0rmA5OfDmlslzPv0Xk
oRjM1H5kS7Il1ADVhp0Ugj0F8MytGtjx+9t/ta96SpUnqhAunvpBpJHEoogRPtugrbALcPOR2A4y
Kng/MY92CLGLolnq9VowYk94gmQ2+W8YW5T87AvAQpIi3kkHaqzh1AdxTXNPBnIBnO4SbBvBKAnE
yJ7febtbmdS2kCxmINi629/2qTmAxfR5yQZllY1xHbDAZ4XUQclhEdSVThaRzuRMra50ZYD3tzgV
xRxXsfIUJdI74lhxqkGZrRD3+BAUNCO51UfvFKUAeqj9THdsug7CSJbgg9DV9nJV3W41oEkr5MP1
bx1I/xsz5uphUNbgGEn9WoqXruP3crpwkAQWAKXhTODycO4CRaM9H+VQFStt4p06SkE3ePmXTfZa
VUpBIFbKG/qal4+v3ZNrqRs/kjyaeIdzr5DlSQfDCkq3MMIR86M8LSpmpconpCrxWo4JyTObIpte
FIzzU/G38hQNFR3R9Rfe7PhEPuei4WnCmD1+pdAau02HKnQTGdVyN3mx5Ctr1sxFIVQdUPQBPQnT
8ZdD39g7vqWuonA809pr25fSA/Qr4Wc75qUo59iWLX+qh8f6uwdF8gzf9Xe5oXOt73R0mwRt3NVf
QqPudp4SAYQIGKLoML3LAfvMtNVxIDPRdem5Euw5ujB1J1KrMh8mTCwASMUGfbvafKmuUSlkfec5
yilK3j0qJJ4Hgu2tx+QUiWPXgUO51NAVYp0A9Gw0sTDn4ml7y00iqA+ccjHeA0z0UAc+TL19Zz1e
/EyTcHHUJ0Gkw9gEuWG8yiIFTu/JI2Y7+VjwpOnCzDp/ABkV5CtGaG6qYxhPSZrjzTWMB945NwdD
62/TW0GcTFPaBaz1XWRAx2NJ1txFepMTS2JnOPCSHvrGHPOynik6H3ry9ET3/mqb6osZUkP9zuNp
YOUtjCDEFPYRD7ZwliKto43EMG6QDeW8DrRjuzwiSXNNqc3IX8UL/P+/r55+Ez67DqAXEuR0fthL
38gJ0C6B8BWE8Ogth62bH1UHrqa4BIOSSdyORGxuSECKrw1brwCNDXEnpUeR6GowGk2+HdAJPjFE
7DkSDvq62G1ZoVphuP8wnCPSnW5ZxJrxVDTSSIXcpSgr54AdHYneRJoDOOSsCAZ6vhGpUferNdW/
ZKaFmhn7Knbju4L7knqU5y+EmPzIrmBNhzeTGqnCM9tL3gOuXyehv2mcxOm/xclQBxInGYXVJy60
lrAQy8Kt9IQLRhZIBBe67zyjScbRKDCAgDoVv8Ze4KixYSWlV1Ph3v98GvjJqy3sIVjWEfThoPjj
5aHyUUo4pldiN4Ad7Av9wGZYQ25B1uYQMSrvs6FSQUK95sbCo0xY34hV3TVWguJV9frO2xKfAMGW
dhf20gBnshHdVj5JSYtgl46CgfM+Cdu4zG6qaDk2QAwUwkbzAsnho+aqkBQSsVND+0++VoaiinZq
aFj8Fn125NZJ7bdnWnqq0ANMn4hwtp65yobuo1hqggPp8zpRsBaVOL2Fg+owwT3sVt+X2m2wlE6p
RvCxBDxz4m/nZ4kz5HGqUYS73g79plyEJEeFcYF40yMP5plIPkHlZwk6HbVNyT79PrNWAvQH1Muf
BBu5hClXKltiZJEhOn7jMH+01aVY4YS4eE3NkY7EQ+3PdOOJFVkjMpDHqPSbiLq9m8TP9BvYfOJo
+G1+zke2b6mfbNp23gnkEZManapOxELeyuzbRs/d5l5RbEnIuj9k85UsIEU2Gjkzu2e8f9AfexUd
+9VH7SWj1v702JhCtsHg4oW97dsP5hEziAxy+YXgTvVZWz6EHzUjdm1uyQx8Q4RCCvxFKDGYYq19
f3EPg2mWpLrsINFDF0zw73KETYaXZE604tn/srK4lvtpKjx/btoZwZkNlS0NdpJSP55VIHcBHs/2
dHMoDypuCRuzBTGycFWMTlDmJ55BHyL9SiOKIkAuk9Pi0R4oYuMU69mHDRjxusV5KIBXOpdHDd4C
yjc969n7kr6dhP0yVAK+eOZUjRc4lQQ+xvbGMxb7zQ4fHJ4vZdeAKWo1zXh4OKSLoeZjQchi91HK
wCtmL9bpwzaMUdd4arYdE/DAJGV7kcvLdd0MsvJjuocIkmuVH72uMY85Zpdxw//4ZjAOYuLBG9Tj
9HxPd3jHrSTA8npozINMpQG0FPVKfFuzKOrac2eFFIBNwmOdYtGQTxqpWKJOmfMFNLo1TZ0mrSxx
1efGk6OSX6qdikZQ0vxD4y3zYVCtcpCNWMz5PLEtlfE/cMpug3zPpGkjKtwUo7r0O/o0GOd/z9yb
r6D1meDinAqxDRi9/ucwD4rzkIzIVgslBXSEBzIk8RThG/IdVL6M1zdDZwC8iEoQDu2qnBdYfUfm
NGdKP895DPZjTKDD8DlT1OupO+Q9Glkhk60A6xIJGC/z8nptnCcMWqkF1IQjMsqmr203cfw4ewSa
EvFVd+5Z/4bu8+6qwhsD9rmf8zxLhUJCCsvk+fQp6whYxwdO57joJEu7JnpfbvlVP2mMcfrdM0p+
Dn23DEYE33zcH9qMXwmN5ibM6DcT+DBGz+5L8O0afRzH95RRig+rznRn9zd0yo7TMZdpiUZvrmQp
eYj/6iAnlW/3ueW7lNkR2LL2ok2NlM2c1LtqYcK7ColUKuY+6vMmWsqI+4O7Y6ZNJhHIg0W+qAwA
K1OdGqNPEDVhGxqLatte+VEqUl9zwC+gd34O5Bwlk1O5HVtLjssE4c3uWmoLrS5FcZBCH2twzsOa
vbkd8h/Tp9CMtKxy433Npvuq+Arty+dKHrGXzEat1iVWJeveQ4vB6gf0sbNoqCYR06+PRdMdVjIj
U0mH+Eyozfty4HVkvRIKy7HyC8oebNngPCwkrhPQZ0omx45TjZ1iMF6CBzIE7mOni8XZKCbwWzt2
8Q0qp2KSgMttyUXdI/cJyHnm9qWvD/6u7rrm7yDg921BZzo17GXwpizx14/crX5/plxVMv473G68
/4vVjrBBrIQf1hrQMAhm+TxlMF33tpGq9z3EIZC9nAaczTu1ymGcqZwGWFNz/TI0cT7RP7422vOT
YX3uLEMtlFwEm/rOJ/OLCNMWNA+6LJNz1uv/Q6mEqXyuaX4EOF3LmHjPa+VfvwTXKt27+o0gNSGK
PwVDo7/FCGyLzz0LZXjS4edHIbeg0YzDqersDcBX57oACaswxZwAfkGA9AbOFNH0ESmexEExbzgM
JVyPIaSLSLHLdT0FlGrfs+24klV5E5VOCgGNd6p73RiA1k6Z0kMgkF9A6J6S4zeWkNtore//+41o
5Q2qXQ7zXsIGHFPNxbSg63EMgRS0BtPbdo1pzjX3C8ta0Tf106P4bCMNwloUvSHsZZFRSDEma6Lh
GHhQJsElwzo1gZIXj26Ync2eaUr0/rR0zl383KcVyMqpHEehICxFmqqj4U+aqyLEhis34vD+8M7j
E6pbfKllRk4FDWCumunzmmp6XJS2OffBTp5VDFM5JlTVmDZ1Ntd2hmDWPMYGBOzrQe7UfEvKw5PG
FiC+K0kPZpKbe4hZ2zdrwo2cfUuDhdC/YSyFJmx4ZGh+yAGQQu72ad8PdN9Vb2thODLds7JnNXfh
d8JY7B5YSfLomrjDZQlaQtZjm3xm07CxFJx5xUrvWTlC+6lVWICuyoUQMdq9RRhO1PoPShYJ3Ygl
d3Yesdcr5K+5+Ma+lSKvORofQR3q3WtQy+cHmtWvZQtsedEwNnpk3cA50i4Tb/q2lf4Mm0BLrEZU
LE4p5o7zSodGyAMHrQGzOdcGJ/HITy3nLeYG+/02sRG/W4/BDkj7bbwvGYamga5f4fNYYGCDhooU
S40W0Famv+cI2hVY8WvtQ5s+L4BIPeHI/i4tbN62CaXFjkaoqA8tvvawZ9PqkmK/NdZ//WITUSbt
Zr9y/Wgm7E0+IUJH0e1YqiCFH4Y+wwK1Q5a9qadN1r1p/mpFDLckSfHNNhYWp0WkUKaUOXQTXlKa
GRfkLOeW6frbpgrGV8s2MtmeZKs388pYFPVr+JOckTRiimPArhH5raq8WIqlAu0HGWlbwhUJME2s
zaCkdPYDTrgxjtBCHmxtUi9OO0KPHYNRv96EO/zpPHtl19sekfquwEO2QPf0ScoBysqfCNCqKN/z
ILQa/pQ8oudguNM8c6ziddiZGJVpFcmF3eFqXAsbQjTI55PlBhRyTOYQoWxUELH0j4dAkgb9DVqu
19VBPYXIVvDNXVJyo+SjWMTr2MFDem5RWYIXfe0fhXOgS/M8VC9u0YhXrEAY0UskD/UL1pBd1qNC
dWrhxLn4HbvuK/Ny5zFzZt2rFuwFx2IT8YlJTf98lxtfxxVXA+Fvpymm1EUbvNJ4FySjAO1XZqQe
K7DL0wRyRuA9onqtTYjLHCUSKt4sUsEiKAiiofzKdrJy+IJjPZgskhRpsmDid/z6AF+RFcdKVdNM
7850+KN/swfqRBPFXETxB9KLUO8kDeh4WnsDxsEKUClhg/aA7i8oTHGzNc77P+z3k+eqPOLUKdjg
MxqmxrXwm13/Ijv9M/hAZO4nFhu+2o3OJmByxkejy5pJrvXUj38mxATltFT1X2Ss4mUnhhaQzlya
PoEDGECrWYX+tzxU2pn7iRJhR92GC4o9Fzf7D3sAbAU/ai5KcT+SOvAfHXYoUBX9jidKWukye9zd
XlLpAvHivVQbnxz9Lpp4C4akzSeNSJvu2xk5SA/jTrwEIaeDa+I9jLNkklAp6tcbqFXN9J6mr4oG
qsRHgjxyDPFUoPS2pD+uZc4yVYzNFibRMSRw87HTqXMs3RlVHstwouHkQBM5zlNLkE68VhiTJupT
MninRL69fXGyKT9SIgbnJObWn1ziEqBZuXLC8Khr1ZOOS89rYu3W4L9M1j9z+JFICbhORT9C5kUZ
ATb0DjmwgIIlYG0oBpzlv0FT7GBtjfc2cnZ9iraWY4iz/ZMNgFx+jDFUAcmgpnfuVfmAOt22F0Y+
eixEOzWBSmZ2Ko1ZVmmKaC29auI2ImmWt4mTEemCTEAQ9JiP9X8nP/5hH8VuWAvjKdOi2jf5+AJN
K22GuRlCrx3Iajbkd3PPFZF90NBJkKoH8bkuZLwtlvhN1p29st15rkITR5slFG8sgLCPleDsNf68
UnXIUOkE4pVb62riGgu16dGzQ2IyZahdvCahc8VeznmwxlxHeZlcoexxKgfes0xtVS5J5p4hwGKK
p9dMdqPOqswmatow27d9qHUs2ov0pHejOpiglfTtWWlzdlusgb09gXtj0cpOhpZOy1YLtc2Jm4rj
sI8Zug/kpfXREx1KnGqLaC8YhhQPYKcY05RJbpz3UaYEz+NS2Qvbmt41IFI9ebQnNvTV6alMY7md
BQJpZcWGHXg/IrMqp6Xo4VdnjfKdnoYatjlqkiHvUMeMnKUNbqOTriQPTK2dBDXMdJZJ2zIwDI/1
IjUzG3Iij6w+aeSOgVVg95Zxf/uOM/ZsD2ncvrsMFnlJ7fhVP6faiLG0LcZo7zEvqVeyDLl6b8eO
Tv8mV8L/EUdLxks4rFBM8qgLuwYSRAzKzjdRkVYDWILcdo/RCI5j4W5WSwNmrsbBghYCTWlLWZ7s
efJgQW6qg6Ju53EEgiKWNYARTzd/jkvJK8qJcc4hzHkNktMVygJBUaryQa9WktAjeuVZElMREIoM
h89dH6Ki5EKwKvs7FMRPpEf3dgTK1uOPS2Jcf2V/3+Y0eG/IBVMzCWg300g1z5ZVJ+YUfPPMPNZx
meYluJAmjfSnmp4xesEa3onzCAyTrTEk7u1qCjzAdUyU5ZJuedbXBVhwZKJZDjzN27AGAXdVb2bR
Rg3F7O9iQtnAAmmEjm2JtUfy/prhJr9kckDHCjWq1pjJlquMyVXQW2qu7Xcx2cW4F1UvfJxLB8dY
WN8xb0DSHhGlP/I3mQd6Bw7mxqyoNe5qo09lhFFRiK8tJACOAINi4j99pFeQO08YEEXDbZ+DTSRN
6PeqiMrGO9citTEHR8u4FjyHh8k7zOaYkinwJqSP2OdOn/VS3+VZNa8P9CPQLPgsjKN1B56MwDEJ
INLOInDy/t4jWbLgCkd0Fy/lemSjkQX1UBoAQFHyAmomaIKCzH6+DHUlqnhc8g2yHtZSC4ia5K2G
z7U01Psq/tltgQ3b/HXG0iMMUcbNCMPjN/F8xHpZPnZxiezgyxN+kEJEF/yWTji7rsCgyQNU6OmF
TfqDO+TaZN174AhvDhyCtthxwSWc4I3WQMe09NWgJksYikkw8UgSOaDzTWOjzbkVcmycZLtr234y
snaLV+VQJX/FDui/Flze893nneIAF+L3E7VwXUUy/yEIjhS32BxYyX6tAK3wXn94k6VE23zOuR79
f/+ZIi7WwuJMcCJkkt7THlymt+i78JsN/qW7Q06D2ArdjbKebJr7ZuwTb0san3/58Fe6pD2h+WXz
0YRELI7S8ITseTm5FuAjF3yr6VyOJRnYt70KE1OPB7RifRBSDi/05LLJCGV1j/rKmp4ELx0pWfdF
ogsOI/NlIyTAUuSw6QYLfrwvX75xHfoD8jD9qIGcpsG3BU5H2MqmlKLb8aUZRWg38sawW3Ic7mYg
rI8QxrBrk9LiqfP2vyYRMfqPaeSCPe7sofdTFCSVFwIBmUEbg3nLdI0KMSZdPOZpvVNyNdbppyCm
U7yIEounFRybajROyfs2pk+q+fGjcaOxml2ySv5F92+wPeh4iTrwXXc6vxhKkj/0D/D1Yj3ZoW6T
N8zgrd8xsE5yX0lpzmJuMPe/n7Ap45Mf6UGz8hTZdKaDBHAB1VU1YDa71bImcVn9lQnLm0TnzhyA
/g07bx1j6R5G0drOBT/VhfrIM48r9z9S7dGwoffXc6RBX89ybvwDitZhKC0af38QOHu5NmCzjOhf
5cL7Ozmw6LRbALzmHtENfMsXyW7Pm/vWJzXtv0kkv7Tehq0wZonBoUF7aAt3JJellG1PGxEbCi92
LyIDbOtiBE72opR8uTiYWCzEuADB6exQSAzbdhz6so0fc8mnkh/IVK3WVevN7XrgZ3Yy00yQOVym
qG+tvvE/UP/XtEyy5eH6/PsC+9Tc3EN801H2nl8fkAbee1NUl+PVsXKlGYEVy8PRN+S7fjseVQWW
8uMFTst6hLiUw1KalD5gOBjc635pncTzAXKinmT1BgyMcNlCvLzHeuPCGojLXpzL33ZL45qKbxeD
DOnSTFw5BeS9vvcbMil3+h6M5oQBexxKvYEA9Gxesfwsq8toosLhR0nC9KECj5p2k06jmcK68YSI
eb4L6gtNcS7SrumY0STflmLlL0uZ123VjWXwa4xAH1jMOhPuTmyc7PSw4l9lpJ/jXKvUmalIcHjd
8eRKixVr+f5fjgQcN9qVeO5ZpQUw51rE62rgJASe5vfpZj2Boreks9RFya1DWHuu53S4dFClQfjl
Z0Aa9gOOviGXdNRM2YIrmI/kDywqzbgMPeVUndBnsnKZ2wYw4O0mjwarmfi8E9vTS077xolGoJP6
UTtMoC78Ce1rw/3tzu/WgspNSsPszOYt5LZDQ5zVF+5qPUWT8wIBehOvWcQuxnBL8fLQi7BIQrOt
hdJr3el5l5oTnzFC9EE+fvYEvFuYpVH4/YCV384/gPkWiOiN3Y5VSQh4x9Iqt6wsefSe8yBG+eOr
sIo5aFTidjE7J+3/7xNDZ0dC8Q4PuZU+lq19Yyh37yt/BwCHkfaTwWl081OFT/7G8HAim46asrpU
OyIjnULRRTSbywVHv+EVCi+uwpyv+LeZXP5+AX8fJIiFIQUtkh5IKrP+s5Z5VUVLGyXwiyfHF+Nv
FH1mtKckpg1jJu1jUH2gGpLuHYlD47eGgyAmp1E6L5n+sZKtJtQSEuktyt0e/veiyEdfn9balOjZ
qlTZgQYJ2vRurcyvi9oXct9PHuKtCHuCwu/fyTOZtODkthIuKjpCMtcHTUEVyAaDpAoS1zbbuZU8
rJWo+z+cR/34Z5019vKnFHU6p8f2BiM1P9Um/s2jeK6xZAq72p2kz5jS/7SCNOdJQxfZEd+717sV
s8gS+nMEl4b4bN8LM9TZtJLq1+gfq3f+hg7sDbPqxOqYG+R+F28zVnMtE8Vk6fVy3x20snNc7uR3
AG6xJDZhMTyrSKgCLObXl35O41GWd+ZU2q3+I6hOagBY3pZIMRQ4KEzduoNWMY5ymU4l4o6RQohx
qG/5hENrXs/8q8qYNlILqhzw0r0f6FZKclQdzpvf1PoNrurD21uYCJ4ewfhhVeGDGYeEOq2wkg1u
Q6Ppgo/bhipmCINg6G4vnrbIGhRf4SbxiKI6+L6nHWKMfVbpo2485J++UjqCyhdvRWGrGoLK17fa
+bobnbY4RTIPoJgxGTU4JXgo1EUHe4bga8O676r0BDjOFJRr2RrcpeJEdpq7H1wSyY3rMQVJ7uLP
I+rUWeAu5vtxHAeh2eaZFPhSPPXK2+0Ps2LJ7t9FzN7BGWMFz7L3kvJOeZ/i0uN/GHOYYFOUfrzs
9eFD/c4cmhEiai5ET72PFI5pT9ZwCD1Ejno7Ipz/p2bMSxCRiomUVRvHHRB+hI4JaunS7Rg0Wj8U
fcNJDX1GAmQtd10oCZdORgf/thCwxAyio+kwNd+mRGiJRqcn6P9qCUXG/scvifLZVMtGVHTP7S+E
4sqVwtE5yrYNvdxbApqj6w2QNkHJuaW9DFxt6YAgg5O89lmbgbUx17EZ7MAoe4EYbMvqeaDw1gxg
nNdKcDhAIvrK56eV27klhqrlReViDO7iaWMPclqDsVhtFkRmMigTV3or2K5+kilcycNR/VvU7DWG
ntmHTyCzoU8rMwbJas7KM2hjsxjpqKGj8qldq0qx0JMh/29ljo9W/1WJEwdtpAtQl6F2rlvMfSXy
U51kivPOOLmHtubLyXGuPSmGExDhf3frAMZEsyx7oE1ChG+y+oVVDbLXCZnftWYJuqODJ7OmJzl9
cDtrBGdEXCp6wG7FMmP4MjRyfqXJtdQCtchsob+XAkzqZCo7TV0Bz0+vbffruhgVDwDK/tavAqVn
V9Kf/Nc8v/cdccSizFbRnLIJjC+xvJk/kc3A5RI0DRewdhZnOdleuoBfntHvgTC83XuIJ7lJUhmL
bL8p9tV5yYRjLbfy+dd27g23ngCI4PLs7UdH5d/vRUBiBscOtuAmK0q6Byl/0IW7xJMQjLQGmM+n
t4T/kAFmWjGIwGQn4OQ2wM/ORN9ZRd8uelgXILExDsDacyIsaJlOds9EqNII/Hv7ae8I1IXE275c
nBDlMjdW6SdlBYJi4eiZLNlx1Sx0vsqP0I4ZcZribznPTDr7q+7F9jNh8qQwe61+2S3/5hNpL96J
nHT9LZpTvKo0+ULe/LOqc7n8ld1u0i0qYXg7+xsmVMOQBXRM16NK3OIferDcS7MgyViru7K6phc4
znMbqefEWAfCtXHfvjrRhsGBRKMFQGEWCwSWCwfqNTWnz8SXN8KkDpn9l5kO9hm6o+i0ly/0t+yO
EoZWn2pBQkUw5yfiROpXlmkahOcLgaqBJe2oX2EdIlB3cJBy8+anGjzAmWaO8uuv97qi4xM6lrRN
kwl43yFOSVZf3AVMYYDGcIG6jcIaZDeyMAxVv2a7x36w6H7bN4mK8jYVhETwcRfjdeUBVEOa4hV7
4vZSTP9hYEEZYzL7ssedO14255IBILxychEKnczZ/UOzk9V3eN+Jvm2zux03USLn1HfT1we+CvGQ
sJ7lqtndKeG87XDrMkjAnijyWKs6r2hYwc3HHPKPa02DuqURteaUhD2RIBSxtBuFtKHCvM6tRmZR
1FmdT9n35qcEwIgJY0v3NVuUezXxf1S3f/u2kU9n6S1Xr1cMyRno8SaPRlXFDrSyqHItf/q6g4Fu
qUWaQPKcwMQhyWyk6dIBKuq3Rb+SBswkLyAvGdo4AZe6MUIbQcaqyrSOkD55lACyr9YtmI+zzsAr
dM1EAputx36s7wut8lA6C+zUF+XMtsTvwwqrpXV5ldwtZJ7B9KrZrq/Mn3pQpPn75JWyuhnPGexE
SIxTHvg3lR5iuQb9SUXo0a5lB/kF92DbZ3WVThE6EAPhf6rl6haHVamzG3kOQTLsb60BbHfkbwJB
nKFeff+Yz2fZJ5RTHmYvJt8huZMSQET6g5qDQX6fHJbS760iY0P9I0jEjs60kTsbAcYvprt7jLlK
rajacUyRykfKle1gM77JMqpBvLA3E7eeiLJT3PWB6FaKfuadSfbInRp5ouROlMNkY3kzprvKZK3X
430rMjwCVkqk1i1/rkr5xqhtk2hqoEZwgF5Vdpl862LVKcRu90coAPOGXlYGbxVO+rwPlrmU+Tex
PqO6++/ZJH/wvtepd7LPJ5jr0yin6/qYzZpuPMmWjA1cnuA/t99qge55BolvcWD4UQgXRJhyjFa5
5RNlJQnN3IFjS0EJ4+mYrk3zhlFJVseRcjblKUINa6pEbvuE2CmwXlFfBZRGcPMu05JU16FJVsBd
eZM47Mji/rLN+zSJ8fOa2E4lpu6Y06uCJviz2kCFV62M8RxsQePzI1q1JXqn/4b+UoTIDOVAMVh1
LYihYaHkvhs1rcVtNzO9Hxaz/2CBBiZzsw+NilF8N0yzT+2vV7o/zF7OO65EjHuzfHsJMYESL/fz
aVXOg44l/1d/pgMe8HXBZ8iqsxmtDWKsi/BowhoVnuy4y1gV906xkRQpoLFqz8b14n5ylBG7VIw3
83DQwaO2gHq3yxaWLlfGuCoP0xQFhqWFxwTtEX7mxoJ1v8b3LdgI14R2xdEogq0YrSkl5ANTUQSP
63V3ay/4HSFTvMso6S51NfrADAlS0WP3HCHD1dvIOQmvezarhfAJddckynlSx7Xo8hKGo8Jxb3Af
DHcfTKpVPc5PUna+qUEF9GAAG/3e8mxzcMDXMNSrj5qE06hL27qiLyxLX4U/HTTOVfnPIQiuc2+d
pEpoO0WaIH+D5yy3K15GylECWNLuhhr0sYYIPMn7dkvD/BJl9ZegERoeiyNHUhjTapETqckKb2v8
KCI2PPCc8h8j+aFxZz5RNXC5g5iD9dRWMTErzCOZObA4fAYv/0wWOoOpHDRYMVJ1+WZmAben9vjK
M1aCc32XhX9abXB++lEcb52rpdw8OiOqIUvTi5xCkvUcmEfsHqyLMUDxxU7AFpEhHjCZux40kMsh
PPnMZF4PnP7LPjG0laAA5Qn3HkKLB9nM+p5J28D/+JskAzZQBtJWnXnVRRf5v07MPNxexlobR4RH
YItiUOKiu73vA84qjwVMxIW3dm/v1JLGQl+ziUF87Yucvddf5yAGuVcHR/VMYifkdd3eIlW/eur6
TVAtkyRIlBnYU0QBNOoIU+GHUBzJhVyHmyQHy5QglQFNL+jltnMACUYxsAswRNBJCGe4bNAtbnhN
E+O4Ur4FnYiwYirmargyYgbQq2ZpXvQvbbTsPXRLeN2ClKQMIso7jkTEQn4RsLgeHVDaAkUcwwSS
eRTE81zHECUTcmC6IVW/pGdhZeOZjwVFa/2OnmwHxWp33dIpxtziLTB+HzgLodU2M+bWvY8/cNcN
qBrhzJVrltzh08n7+JEcPIJsCEzTAeNzh+DiLXLE/K1DxMG0VcOHsywajB/HlIBbq0RJw4hWbCCy
eC4HFMTFZlMmjZ4mEWku77USStyZxOG3HZqmsF1wMtkNx2QwUnUCJWdE25S4bJBVumNBZoQ8Ri97
rSRe27FVJGhljYoiI27P3Wyo5dEseB1bwHb+5wRhrej0ZJmhtrPLpQPqrXe+EcnKOuMdbnOKx5aA
S8VKakRU6chPP7ieOb8dNulx5n3y+sA2CEkLtwWqqxZWuGh9koAzcP6hwKFWNlPZIiDGSXl6Wd6Q
w7LWBiABCu+GAm6IWuugiPhYzidOoBUQV88/u5uhMVO92zPhUjmiieRFgXySQVSHVJ9WE8V7CCKG
/JkznYr9QzfcKdU70NXb7x/LuENlHcXqTcdxsbhV6opLSRlwC+A3cSy8b679jA1lAhCGg/h3LQuz
dPAtHI7uQR41TSLOtKXgbmHFTecxLQ/SBE1z5XWGcIxh4VsPt5q0Hn9NjLwJtPJ50c0zyvMEukyH
bqXV6rzPRcQG+SGjfH1d91mGJaMhzPItzRKjciOxhqlfZ3sfQqBJPiR9qcY9q2pCw8HrQqdJJ32a
yAieWprqS+8MeCSa0phqpTztx2bSoGw7i2lc+7JhXA2hk/NE9r+29NO5dbb4KCS8w99osIWgrApx
kOKCoOGWQq/gxpOoL1D8vnundeq9HHYwXqwlG1tgqIOav2HeMdBu45QmWijLeftWKxbgf+FAQ4NP
A8JPi5vnYlV0ym4Qqtdn8u5eJ0izwp3m1e+uR+xgvyZ2UOoigIBrNzgNc+AjkRBYIlCR2TbkemUq
ZQfSch/+ByWmCTIe4FpaZVsOmwTGFAigLvqhFMWuunDxdAGrHcIVK3VoKW9dnDZbhKoQvgIwSe5R
wLsLx0ui9I0K2ekRwmASiSvp/ahJ6pXoUSq+jzeMGbeqhqTktErnSikR818wh6GksDLKH7bPJyBG
y3xUnGalKYGl6twbEVK0x7MTM42JlAZcZ5t1g6pGgT9C960bJgZqwG8kak8ZqCBiIo0ND0QIHV32
qScF/IBcR4w/p5THdg5bGM9zMzRV1U12J90zPIQgY5Q2yuX/0ea63DXqtw88aEflYQb5giQGOK29
RV1EVOXvdRp4IyjXQGnfq2xcnmt/X8V1oqZLF2Ie4prOy1f0oC2fp/KPbUghsKbyqrF0bN/wHYbZ
vjJsbfFt21ab9AkGx32AQUWNqrG5XK745EqQ+BNh747YUyYMdUJk1BzcchfSUXUqNKjoBaGbKU2z
wR6VH35aN0bSe+H2op+EBoAxjaTQr2cNacisPF5ktN3eXtGG/dzQ6TFto0T/BGwn/F6RLN3doZcj
7LaAH2UoZgdO54bThmTgdCYfhzE4U1Gc+GgoCv3bjUrM0GsT2V/YzqMQk9Iv+EhOl3MmeNBz+Nu3
xAvhclLkVEFC8Kq0Bad6FG/3H+XizB5i1oaPwnzpUplXGsx7d41OFArO6hfFXEajNGjg+/8+OAj+
qfm4JVv83rmbjlS2GhGStVHOEBaasbt/C03qxw5U2/mAx5kuhQkg50vyI8GG0YpxyJMSROFkPgyT
qSXyAewDY6hkOVtiuUo1asm0YARIubbwIJzVUjlMN2t+6a0ch2lgMcO2HwiXvzYdBymGqbwDplKm
37EOLeujUAUJnRhMa8fweQd9+w0h3rQFdBFjKaFsRu/RJdPms55iboDIx2b8lR/832FWxOjbWGJT
yGC5NqJ/WlDlAHhpGr2woq0tlTbv5134h0du2zkk/fEd7jVLpmHtYj3CbRiCNArTiaAd9vwrk3E+
zm37eBgjvxvKt6T9Fi9t5Jn5qaqxSCrJXOabeu4+An3n2Mqat48dfQzz/fOjbvU7/KZn02/4Ux4k
2tFN6TPhEhHSq2D3NqMBxVV0NSGVtJLzQpP3zoaGLArSXbaiZLjSDmYkDTwJocr6q60ehSI5QpJK
+k4QPVCowcOzbOGOpSin8MLcrlzhRCySyhEYXG6peO+gudAyOrJC4qV5P9omkXPgbvCS4JeuLm3n
G4Th4je26ruU/XwF/5reAAV+K3fHTl4RLF++Q1AU0A523pJI2mAqmtSESk3l3g2ctpOmIQW/EfcD
CjfNF95fLCRQiiCgwSahnBrPdzxTpYe6TDR/WgSAf/MZCNNelNfkc7+ZPpBP/9VB6ORF62bmdMUz
g9RKgobDQejY+0HvJVVBg3Wwwp0H9AisL9p/mjGeEfk2TWvAxpRkdqrzLddax1Ov34kVu1mb7V03
Dnbjh89XICnqlDjmMJGch4TYsbd7ClMl/672bcNezhxxWwR6DOMv+5qO945KXdR5RgvIwqsOeyPR
F644FfLfzp9K1ghOTIART3It15sgfVC50HebU0lWVYLYxDZbKQ/bna+hC1x2u3U8O3jliF3XRm9r
pNqm1kiHGLoZdc8+27bE4K4ElIPvoGj/xW3yxvNn3fV85DBGycYxYA6hkKijXv/OyKp2Wd8Ndww9
CPWiy3KAg6i7+QwWRE+JSwQRkBYqnad6xLvkvfsPOg/xVPJWFOnESNAuTySCfXPp9BnqTc6A6n0E
dAl6sSfKL5TidAYi1BYW5oHIQMT1HqaKmNHTgBthaFCeaUirG0Fox0KU12ePlZq2aUp0XhUIfeW9
DnX3pFCMihAfYKDBlAuin0XgCR9OVPwGGiJYMbPBTXUixhUJvikNU2vQGitpdEZTXD0MqMGKLDtD
xWKaLq0RiG+SfoM3carAOyNwmoNRsrrPpbmeBKLwwK66LQCN0TXS6mym3ZCEJyj0+yqqkS21T81O
64gx3jxG1eQcO25foUuaDU9LQVXmqFYg8OG6PkZyJFosYw4QXKGb8wNSyEvS5OopCQhHKibJW9Ah
8K+yh85mQiYZ/OlYPFyiaqgdeH33MKNxwZ4Q8nPdnMVSxtwzIzwKY+gcbyfVgZeafyzhetu8qAw0
0Tvs38m3NSvATogFWOe3UUD3ovBVJEmSJyHttTXYLiGxfVH0DU/8oc4HtecKrLGNw11l00dHX8d9
e9zmlQyFJxdfueOMbtzGHst6H/g+M51k9RFYzNAMnuvx/qqNXR9doD0cXTKf8dCqKI2ENE8XHRbF
PZJoqfES0zJLaLdfMOs2kCEaKbJxpLbWjH2SQUXc47KfdjbIZZJHCWRrVYciWcwF7f8I4kzp1m9M
/qCdRzUx8rdEuJl4/lhHwmKoH2TsaUH6lezPw/lV80aMVKJCbKyDqyy2j+Eui14X2ubdLI7nYc2b
3ktV32AwRA9p3RhWj0DPgqGQbqznukSKG09n1tei61yID3zbxxhFelWqd3h9x2f3F++Lj8VLB0pO
+BkBMQ065BYzQkLNa0AlKQi4ZyUaG0AHko0pnRHudGwcK7O2gNvvmmTBQjMXDMP2oWq63CnmyF+9
H7Qfs5lS/jsgz37oE3cLCVYK9mXJluXzIvVt5FZW4ze5akbWqMySmHuNHkLFOZNsNNLdv7dmLuwa
Dcjrj/ehnBkEs0lfMUjKRLC5uQWX6q8cz9JLJultUjh6Wufuxrs+u3SVJAZVsWNEH5IWir5dOduI
UhQfwcpsmMMxIITyjFnPIIbt/OiYOsV5t8JFrReYkio4wXzPjgeBjK+KyJpCOffuU2AS72Y+TC76
rgc5urKUmAGrwYIHR8Z4At4pYXiBT+jJv5Wq3g3es2PnN5a2po3/aSdU0WZzAC0FDE0ZdiGWINL7
sRK+CXJkD6MPTC9vCFKg52Vvr3Tt7rneYGl6dJSMvwwM7vibswQnTlSLSX/xkyWS+bDuaENnbKd2
rT/FR1gsOKgaqMV7IQI7DxAJLT3wh9w+s91AL/Blfa6DCQ1i/itvlzfKdO3f4wLjwG4tbgWhiuvu
h5gUs50Al8B4sBuMd5pRHfVelzP/Epcd8NMGpIkZUhSGI3gBE0kTaG/94vFVF8EVUU6uCTXeQBdE
Y4UHgbRM6zAQ5F7kktpYiNhRrg09AF9Sli5yyKT31gXmihbjpZu0kK/62VxCL2R5cJI3r5cG9wrH
9psl53mr1XU6CBWdxASlrwZ3ks0CnYTucPAACFUkS+gtON+wgNF7ioL83PMK24ssFUDRrt3NGROs
kyzZHiiBCd147jrrfPaqyCb/uRGzZHn1DmulFRGjq54t6rJSkbW0xv8/CAjjxZGDVC8isjkCHZzh
HGn5bDUzaeTuALHgFO6VanlBzid8oTus3VyTLKdp4ihbclOcQw4IJ2QsmAtIo06LWtOP+HMWcreN
oc+aQPe7bOYvyFW1Lew54YLo2/+x5VcwRMXu895JP/fdFkAI6gOS1dHCdN8UJZ/skMBw86NCRAZ2
lOAh03FGQtrFbrZtZt5gIdQBOE0Pm3/waKwHBRszA2+AKaGUSB5I8j3hovI+5nBDELBvve17FAOX
bVu0Cc7uUo/rUOzWVOxLdNXcq2jDI4QtNZpHp4Q1yiilv+v54stW4NihbwqmbtDUp4RrJClxZZkW
WPSmKuyMkOzQ3YisyncaNfuU3CCUTbaP+FJNXnDUeHXLLJbNTyeJIDikBCPYKDhS8SbzRWg2IJAL
JR8fjItr2bOA0Z+dJMhmy5Oll6rVFKjwLpKIXs6RrgiQsxqneWgy4p7r9ZU5G5OIxBOeuLa+RH2q
yZvr+cOvkasnKtPHY5VSuuaCsD5hByLMteBOoBE14UDv0eiH9NEbULmVYDWiCbioQQLSHIiGa6Oo
n7cOD1dXq0QofS2BQ2Wolcc/P8OuAu+XJBWC8hs0uuHDOrDlOwMNIQs9bVaMM7sBee8MgOU+hc+Y
ppSCUWsLIykB2Xq6mFyAp1IMQqWmvrIVYiHCyTUSPYMBikvdzncDd4AmszNHxGQEbATPK7Kr1y2q
VdEN6eo187JJT6EldM0KGdcE/erDpQnydwJebwNEG01wQBpLK/yJdSb7zwvKDRA0FIEKVLFQTPP0
v8NtKDY1rXmAI7VD84IUsWr8NLJafXHql0sqcbCa4hson9PHBM1T1CCSliScpsWaHtkuHZaBn3AA
L8vsEQSLeVjaXPNao5w12lgUtgctuVHf3rO5UgZe31L6LZDC88gnhPo3V6c40m3Qjg8yZnB7yfkZ
jIfu+foY71zS96gB9sQeFtPTp7u/U3kUfE4G1KQqtrqJmR9vSUBsjwwS6FT9xrNUKmLKzoLmCQv/
360YxPBMjt56ZBMX6ft8xsfkELs8NUA20NDkqW0WQTVIT6Q2uQsAvkA/wBGTJtRm4K/WzT7RuCGz
ZvdT2M4WgnhBjE6w2wJO29Sg+7wxLTn50lq9Zl/thgza2opHZ7NTTHjS7NapXCIaKldxhdh9biYx
acH04x2vCasNitc481sGp+b7yWyo7uLncK9n4tOvKwXsF6ee/HivJr38BF0H8931ZqfSxYAU4QuE
aBz1qkTQ2GhB1+aPliI+6lN1Y039I4Jzgy/6DmykvnAVQygCWl/XhbrtGMCGALWB3WYWVk0Cuvri
PkFfl24F/0HrKyXW7CpvH8R3J9uBpPS5AQsF/oLtihGBPIVAcKKqHbOgTDMLe6meMCC1Gae3lzV1
pmptu60p279zpS7eEa92fgUOYB9Aw6vYu++5NxRJKX8WvlvLdwHFrBxDbKpMpRpzlfwRTZsrsg2c
fGqs+f5R2yOxxrrOpp6kdHXHC0EAjjfw/MktzYqQY6DviNsV2QLNtc2UC+gTKNmjC2olcguHa4PD
wGtIJBsNBZeE8dRp8UAgVruwFILXdo38MCpA5mty6gPbC2ws3NnFh1pl20SXxDTnQoXb7TuJ4cSd
sXKQWmApdJi16wL4tjjAYg1G8eyOD1L+zZNGdZbXKL5RtFFHXezoPuE8HG7nZDWFFSwSQzD3nYUt
5416rYTZKNX2Xl3psvXdE//MGWMh1L/mPzPvUsT3xVOfo8QojF5YTEEVLlWImqCP35P60ir/1yxA
f5SrC/3zjaTpDCe3pWPZT+hDcz37OUTVvNmu3zzgYykpgVptrU7TQaQ7tvpAKbxOr/W0SX4mENid
BjtL6f8ci1N21C1/8pvoLz25OJhM8dXi5XMmMIYiPESHOCKwNx2S/KlMYwC5lNd8x/BBWISfmYZl
/IqTi0S8TKAmu+yWVXFsxUvrm6+JUPbfoI9H4IEyjfgu4gbLz3/XRBxc1gAK7tivkvbFkc6qSAVJ
M8SnHunhDtV6c3Xz8LEiSgMwgKjfjNuUID7WbJFELX+S3uRa2Q3GsUqo4nj4Tp7iyxHHz6mY0+B1
CpyDkBxLHTvFJ4SgFtcKBXv8y/YU/INM4rG0wxJXUwJA5kgnBz7cZhRz00gmyQT71Ix9n9GPNUW8
7n5HnLiGVpdZIMsNbJtSRIJ32LHkwK2VPRW3str6SPC1RxfkNm2TZ+ohxwiqRMGdGr/EhbpGeG95
zyZNnbCZcgzL806p2Nm4Mt8n3NzYkfVg6/zkX1MIeeq6zA54Mu+G/PXZRtAD9wkgvR1Ild/GMbxM
vShcC4oOQzDVvnh4m7jbqG9lytdblIKmGi0I6FIJGSRzxCXdzUm36UPxaGXlSsxUEj8QxPBeuUmi
CZJS78qFrZhJ/qbnXAgQCAv20DX5F6O0FdnauHXWjXKQEc6BIAzshtkmnWPzy+uHNsACTcRbUra5
H+hHurXSqJz1wOv5LSJV3Oq4d2TqgkM0iHrGfo6jK0VTXEJW2veEoPkb3i1FTn6ezl1lb0NmrkOY
FtYvvWj4NANXR1VtP07g+e2xsz0Cv3D+Oe/Nqg4CviFVPGa6WdcVFENG5nVmDKJOmFoFcCpvkndw
PwgKo/rMHURNmuBLqK1Uy5+/xR6sgAcD43kQLQPns0gig0iWZC9f355kVe/hMQFjqITH+Fzc1GRN
eN/xA8Ptv2MojAjpna3FoU+EvAYv33MTJUKECFnp99eHk/UwTMCDBlMoFRWd49cifC7nfnPRlrmy
oa6as7TaliKwr9fxEFXHdPYPdoyUeoH47/D6EkY934+I4mXsM9hXz6bwmEdGQIn0TLyzG1kIde/d
KlrIoa51Nn47q4Ib60juZ0ApFupCalYlRZK11N6doKljpnwO2bmXabCoY5tUXlKm4mri4wTpke9D
H5OeGKeFcFbocXo6137C4anxtQp650o9JcNA93ZZi7ZoTlIaeeYd7eEFYi9Ye/w6qVjZqbkSzsF3
8MC3nfvmmd5OL5GYakdosK5iafSRLZejpU2P6pSGkjGbnStMP9yFqZrSHGNBgDq2LMcQUes9Vq/Y
eNYbewRWCNOr6uayLYa5Pg9ljAAp+9E9r6TZiVPqMWBbxVNo1xZEZPSGt44DQ2hz8Q7+wuwv6RCx
d1jcaRm48PWuFqwxRMoucWqnddYcqiWtZxBTQOIH0FBkBCs6X7/GWdioVjesaUgh3lIEn4FbvwWh
BQzX7GTiVVpiD8kfARVP16i/mSc8pMr14yO/09wxQq1R5dboFX7g61LKGrrUKKvbHM35NO3pOejR
F5zpZUG7FgsUbMyViLNfdxpD8nD534rt6E+RMbZNS7FQp0ghS2Q2ew6VZiRLYprp3QNB1hf7///2
M+6Go86e5qKofqLzKnmDcAZyLypJW5HaMyJs5x6dCvFnTX2gco/hmGxNThB3xB9ezoS39wU9kdfV
SF/u8pGE3v6H1i7nrXugII9x3fvRBufM0wkm91Tnxi2RbkgWVDaPFKSW1EJU0ny0tLsscF62cpAW
gP2XiJhLd2g2s2dOL1/fnONXH5wSXkwsICV9Zv1F72JRZYpNHTMi029LZ1q8yVWRJP3iOgSJVnwH
SxwsDWBgUwZE9HqKMAvOUMQSoXn3pa9arulrW9WncUUMOXfyXWpx+swQjKUnkRmVFK1sRelDvlqb
+x9NwTqjyg0aZdgqNz3GPzR+4K9ma9QSoSLibd/geQkPDTQXYmKiLb3NeFjv1ZumMgM+ZxGdiZ/J
OecYmAzFqk8Reiuz0ngqAsvFHSoHcxSKn9eZ8iEZ+rYi7lzn38SDEWwwxdP3KxnYvPmuj0VGlob0
0jS7osUY/SOyBEG+V3bU+Tmsw/uBb4Q6hEvmyQx3LZtrjXY73OEbDg0Fpll1VzqxwM8pAzkbkUiw
o+R2YxjBq6hbs5Dn855jhABYMW/u8xK3EHIk6NrrWLbZBVwC6mFHFj3qUwBj4v6BVMGGBMuE9J3f
/xt4eeSAng54gILtkOen7u7B1k1AGMaOkCkRRbqyk4KEXbdHB0SreE3fjJd/5JDxMJlGmheBxObP
eU4gyFjcRb3J0us64Q5n1DnMpozWvVQFnDUl4iy61UUa6YeFRJJ5OP08ReAkoE0GdtCyHIrPQeOH
eYE7zpsLgr5PWVwX4WjhCynraQ9CTAXwfdbVFYI6RfHp27X5xjZFOCQXUWr/ZCKNjiKWvP30cAtT
eyPdKQny6rTZK3IuNj62aRgBnSD+nNcdaZzCW66Hhe4rlGqA4/9kb2eHd8QYliH6+pcOALpcb9ZI
7Lg53KMafMhv1Q+X5i7o/zOJkDCYNSrsFOa44EEXfSbjv3DFmVR/EbXAh5BWOGeQyFLNDhOkTZG2
BkLOQDlaDgb+aVdLtUGvJtVDykuanoN7LkUddeAFTMsFzsBlYNXyVWCEiOpsyQ6M5r53QBemUiKx
UaFQaCC2BZ+ScCSYYrE16y9X6X9SLM6mjg1URQSWqzJVmf5Qy9l+16X74nvTK1wpU7TYticGeCAd
5QMjvRhQgQvm+cS/NOXa7kCN/VgCcAbnsCkPW4Kfjj/oW/GZmcInAUuRH4c7JKJPRFBkSWZkS0zc
qgH9x2RnnzrdHMJLipqEPJLqQ0qjq/Fk0LIl7QTP4hsgrAk1mc57HpJRpIC/DomHzda5fSTejY/a
p/JdCVSCXlFPV174xrjRTy9QQ0geDV3aXd3bcYwsUZWhbHpkjsFHA+FTluqQ6syiAUd84FmhG8Le
yqkeV26jjoW8L9b4XmeRM0VFpwmma7uDhF8Y7kdxeSHzhkk0IiruInx8Bd7M7nOw0tVx9cZ9Xxs9
QwuDU+7x38rp+48gQ/dEEkckc0ZlRll6G9G0rOJeh2NqJB50ouHDtigdD9iAcSeTDskXoaalmBC4
OOE7x1Y+9SOlml4Egd2E4K6M8LPAj44brrcOry/ZJrEwVFEkvFWKP7k8PmVRAb9Z8nO0Qi7gnr4n
q8b8AfutzYym5Kg13TTRScuPDz6h9UaJe9zlpEvOZt25A/uZtmdhOk/GOeuxfwHM6w2Q6iupHXyB
PNi1Q2WlSU3fQxJWz7bU7yanPoDKaifUbZkWkkpTjBHPJwIqFFOscMt2GyzCKz/7kAngTYpTff/X
V51Qkq7sX63MIokcl+cA3rW9WK9TIiIV4Grhxenef4y5e+DRuanJH582M9hEdTNe2OyiLgROTvF9
UeIDztER35X2XVo4ZJ+gtAMuAgAkVd0B9YubvBGVGmRDOdnur95jAXjXwsIgQV7Kw/GJmKnfFnut
OiynBYcf4lgu+VW1qn6SMEfIfukuEzCT3S6XGCKtpxH2OsNQDOvcWGCq5c7f97lhEK7Hr2rY46uF
xHhsbs0gyAEZoOXYoZHMxJjlTOecOrGBBoFGT0POBjfGdNtAuhrQ04q0qD8TWXZI8la2TUdT7+jf
bt9uNUZvgJSj5mj69VEtX0EEufCXDLLos1m+v+ZdfuPhJqe7sffq6LL0hbJ3zNzvxKlhbzXTkhDL
QRZ/rpYAI9WAi7IynEQ5khs6EnoNvaimoaa+9xPvYL+JzH15rb9wQNXyPkLm01ibTf8zqG53zmDR
Au4qkTPR+zxfGK1ydgBQupM8JvTiokZZGmYl1ybLoDsBGopkWAIenrLPzgU6vUcXEX1zSSfjbf8e
OHFeFIsBL0UOTJCdgB4wWh4V7o4ZI8RXFLNJ63JdGOnEl6I6XkhEZYCgs+eV7yVSCVvRHfwuesU8
4/0wE6RsE6Mdq4YwzI130QeWJSeYKCMUPq+nt8Ac4yPchzrPFKIhQh1/YOpypfhEF81mgoweklYr
DcPqlez5iZ0tpZgJCrpMQmhIQhtz70tL/wEmZ5eVkdxNMQHx4709u/NPKsbrY+BL15UjkDklIo7S
YWKI6hHrWHFH9AT3ztZhUJvp2WWN4nne6xusbRF6e0GKnqii0Xskq51Oo8EZ/SIEgacW9wZ0dalj
ZolXUI7dh0kiDIFGTnYOhI61iMd6ocP1xnbis73TpVagGeUD15IKhplkuW01g1ZB9mnDx+Pg+ncS
qxAxorhlW71eMsUebFQ80MZKX7doqZvtR6KWrZFQMBM2kgV6Ny3KpzcgdCRkGbMxHs4WputUoeMj
WtXpSiZhYFMJqkGtQzV5KfcpPueZ9G9coyHdZnUDqfuGzO8u605VAs4LktRhgFxEZ77UwtKXCEVe
PY7oWTXqCaJsHogpgHeK5dQ0FSpf+4SbxQuHmPYf7kNBMXEB6O/oIQqQTmgdRp4bCgUbw+4bjEZr
aETsf2fkysw28o8kAlx1aoXs+VDLZIcxNm7VCYA02cm7ArrT2L7swgkbq1Pu5wHngDYuAs7G/yVe
aR9y4y0TzRxBpCYS34arjGUECmN7Fq/F82YZovluH5nlGmO1yKGJH+5l6AbmhtgjUBNnJi/R9b82
pPFaH+H0/h73PphPoMl7XBhbe7q0p1cdMABaIQ3/s56Z6p7c7JLCFZKV9/7JMWpsqC/XzufLe+bf
1OzlDKSvKv1CZe8UocTLmQ+ng6FLAVPVNUu1FQDwhzBdnczwHZ7s8pzFfc6bJXeCtvxf3WnqPtb8
WQz93dLUMLdxfsVdzZCnIt5zkRqs4yRrMZy/dUsAYQQ5wnhCu9udzYB1RWPJp+VjzJpriCPBZZ9T
XNr0LolL9/s/8SMjRc7ocpM7JpyKLsHeVP08yiIouwdn9jlaLE7gtVle2vuHijQE8q+puSicM7Mw
+A2B9f9wrIaoyOqcphXakEcWiBo4MNIhrHtD5I5GEPM08b5IRjJN0K79PGc8lh1iWK18ozQMl1OV
cju5nDvuSjWXyODBUjCPShpR8G2TobvpG7UxtjbL83eQdrP6DLQaY0zRMpf/+SG02f7gZE2HTdEL
7Ju1jn051+MwfEsqI51PsxC4zwaPco3s9otQXInfQVhnAD8xehJWOjmCOWATDM+cdRpD+IFrW48K
jS9QT6MstB6K522bCJEoHPxlKJNO7zXQuyOVANc8jaJ43Bqm7KDx9DvxnIBEBBG2wnIPuOuv35iw
UI9XaYwIHtzF6madrQZv000QCrDW1ih8cTqisNzH1hBfqkF+e+toNrNKKGRj5PMBq8Nz/JUvTI1X
ci6rquql1V0UK08sdMydrk/csjcb1oYlSGiOKUfZ+Pqft/YEy9kcQklV9GmVhbT0w6bHmQ1nciTm
JKtuBZKcnj8QTj/LYwWjVt7+uUXMM7C0qfy4259c0bjiP38BV996yMDL0tU40TAANqRkDzcoDf4H
RgT/xhl1NzMu7uQBkmNAOLpKbaHDjizYL4267PC6PrsyfbB4+vgJuQPtfQWUelQwIAf2NqAqb87M
Ucv1foLUzPEqFd9vWgHnNaxx4ZLx/Swv0+AXIuzlH19JGARPx4/QEl6EErC6euXbFAumE+nLJHIG
TouDFwnUNXYZLrs3G0mO748EYdd4sOMTZ/LImhs2NmMCjRZ2+pAD9JoPBeVjJYjN9J0oweWZ6U6y
5n/4+CP9+aAuoMJmlSbypuT5ia7iKEeZmQn+daRZaqMRIn6FQWREfMKVBKzPBF4tdsrJrvAQCMM7
uu8/kASpUzWsYwYVpoSMX7X+Xr0pMG01Bi0iW0lJ8gGkxh0HnoXkOj+ffhAvQ0pUDSog6YGAhFTk
x0fuYskGM3pPwE+8Wr7W3iBoJmAEfxIqq0+JpfC/0Ln1QHJYhnH7UTPNJgW/Ec/bRhCRBZHdtC7E
uLQfpw04veA7TVouraUyxHO8UsPgdxKgobjDbZvEOW0nkuxbUnrrK2S20LIjrXc3B2IUz9EKd1dM
a+1IeqCl0WyoHXwJYKk0T840dKAFCWvcV2E5vojm0mTrfXQi2vDJJuf2zci5C/CNrO2QdWSKCnnb
jU7YTsE8UfVWxaD7JcLd81pgGXx7fXUXLP/7eFenWzpxnE0kTV2eXpOmHQzbXKUogNpVIWveF5tS
dM9IAvexzdvvhkK9MXFMnQ9ncRT6yJci2NsgI0QYvbRPZjnoRUqXWIvsWkfcRHcyt12zAI4WG2CC
+ue67wv389xhxCtbcMGUGupHoaOEkuS1y2B0FGNWHH+r+Y0tyIpE60pwp/grvXpH+KM3Y5pGGpjO
1zpYfAtIN4YeCaGq6K6PG9Fymm0wLvhVvp1Ymo2oy1VSxxZv1oK7gQ3wZIjahg1ERgmjlmOJyvvk
mkJuyD7K5vVGSMBp4FF6e14rMo99i69WWcXxtp73UprbLIysA/UFi0xnrChrs2C9XntlHf0wkor4
7eFJufihdq0Twyu0WkVJ1sB8Av3zKO+szxW6U30HDRsyvdJF8crGbz1/qdHQPA8mgcVY/sH41HEl
taraaYsevY5o+pv6TJ6qHZHei4ARC+WnMmyJythp6gGUkvWlf4/Pd+jk3PtKGzH+PZdPPztZfnhB
WwrJK0M14e/RdKp9+C9KbdUslvbCbdqYdZVYGbIGfIwNfcn5oD33Bk7oMQ4sA/N5OzqkwLKUkGdt
zxPnFTIIXdtvniIeHHJoaRgMiea8oRHu5PRXQv04e1/vHrvYqUQDna5NYYaGhkAwd95VdL0cel3T
gkEM9uYWOhcvlMEqQgyFPZb4r5lIFITrFQdC9oYB/Z4nThWXgbn/N7oJPwn4ANxVkLzlbEdeWXnQ
z4GIn+bibzlvyHTf+dYD2qVNSwWSRXZFFvEOiD3kOGRLs4D3C9R5rYvMYYdu+pP97S2xWhQdZwze
Jjn+kJOc0h6lrixDesdhoCUEv0bQf91YA399M0tLTxk/CYMUlwXfESpEkutQ1+FxW1xJnpPX9me2
eXMC5QHiRwauP32AkcjRuDOi/G4UUUpAzgI9Ep++Ab8spDQO8SCAWAb4Kw964Hve7OgKjGmSyZ0r
X/UDpLhcqhyXZssI6xUlpiPYAVkfLudDQcj/kgzENPABQPuvKiT/Gpn+htRsW7oBXGIS6UtohMaP
xNzy6Xz8bGF4uB90rC4rAG06aetER854JSk7FZlBQAfPOu1hawgBu0Aew7i14s56S+SbPJ+OlBCK
60lm1EsPrlWxsG+XMX8P/WJmUILbLcC3/BFhDZJtNsvfzIehOe5394+yMrBUlgw4kLyGnpvfHWOm
qUfcXxzl0p0LrqvUufZKzh1CNNX6DILSXMeu7Lgf+YL1Z6+n+7wEg7dLCZ/FkMm43og98VIr1w7t
L47rla7CdJ1ccr2UcCb9AX1H6P14NEf3HBOAR672x0CXWza7pTJI9XxMFK4yWzUql60OocMXuuVL
3Y3P+7YWl/NZxjBCi2Ie28bo2S4AzNbDdLWafMgVp13D+kNG4sWzwW6zwyav+aCnjBfC4ZWIW1PQ
kmAXz6y8HoHC2inuCkARFXkU7uwsQdB2r+h36hqjs8o3WsjOuQThnGZTo80Stio0x3ZS1tekheMD
01hpd/ytmHKE/yVCKFoZ13ydK1X3iLFFH7idLJ5KnYfWXpbi5pP4rAZf32/F66eirZA4cniGIuQp
ohhREYK48LCUBVYyGAOEWxfStit8iKEexD2AwYSlfXP/3b83o8DinDA+x07Na+0prKH6ABT72Fvm
lj6hld1Sft+uX3WSZrSLHtiMol9i/EAJoV/hDD5s9o9kzAiVs7ol/9FGsvMgGZzlYPqQYlBgIdHD
TV8dz4bOmYSbsQhcUd5b3zxx/WYPiRAEidxZ/E7QgxhBRXrIL/rESdjRByZxVo8G3w15gqe8GlPw
UaiB+0vUcqigvfdDkQL0TlU9rMiyTRiXDUvepp3GaGQz4TxC2lehPiAdUZkRWjVuv7zM+MKV0LJZ
tatU0cK9EI98EfayLzgrWaxAu7uhc8eBPRZXHP57WeZNoxPeQjPN2Uo12TRG/oE6CMff88mGiDB2
CKi/tvM010d7EQzuqJQmOIg5olBXnKLE1VQK4VeoUhUwRaloO8C47msK5s5l0jzFXX+1s8D+SncJ
ilE2DkG6rY8l/6cIeXANenlGFZvNphuAl7Edb3+wB9gGfLVu1T9enj2U9PkzhGCeY3n1lsmVZ5o2
VltX4iDs4LWNXC2+DFHInugbjBu0wEmUX2BjCWCVXPBZKeZv/GbDPzBo8xKgJ8F0byZuyB75lhBz
JW2maDFENUy4ipIrqO3VpKzkY2ezU6BixrWWEbizdyqwCcxbVkazpgmaRKFmfYjjiDk59jpwhFXU
28OruD88ZWuvO0m8WgGMsykb9mRjT+AlcqP7E5I2i0/SQ5QtiQGkAeB4Tf2aR7sges6Cs++aRdqs
+tgPVfrzJv6q4SzuZClwOsaq0oWyGzWLPAXXd3RFCHopzz5fmM+DyomPAwTgsBo8cImUbjJZdKXs
8SvM8bOfd/vbbgzHwnz5NzxSoGdCL635Gw83uJOdG+Xk9H7R6wrQihzUAryjQuo0PCx05Ss+IyCZ
WtHYtPl7GB0iRWMiuoiGxMXWYDH5DVBPGGX0bEtPBMIK48ETnxfElI7WXGbwCvjmfONsaeJ7ROkK
WJwC57xzHr1REI7dpMifgqAfCS3/J9AqxNFdHeO+MjXRVZ3wA3onfQTxTgr83Zs+FExi/bPg0gpr
ADAEm9/NRIqDpi2MyV4VwJVxbah2637WbEiCt2x5crJug9W+eqBsx9uCmXMD5Ak2Nyf7++7WJLD9
Vy+vAYxeGOESa6HIcL/1TVZc2ifYRQS+OeyGiqeXKv+fZetkbQ+1nmjoznv0BaRY1a8kUWuKdd2Z
rcCwBSa3osYdQOMdKILjJyVhxseWycTtYYVRqo6Tl9+0rhp1c/Zg8uCuicGMR17ozS+5jdFCNGLR
ExtEnfrp8aRr4q/BGha6DgLtb09OtIVrGGv18z7smbCvFpk2n2mst4d3vGJpGYpMo30BSyrasLtE
A5DgXPG1Pv+TQQ8gD5Po45MJGqfrvk9+RCytky13pQSHcHfy2Wsid//cBj940se56j3zal+zaoCq
UsS8CuDBkt5MmZdi9KC0Oi9VPQNseLeRVMJ2cvHYqDybRvRZD2I4RCRyq9crKzMTYprPiA5Z6eHJ
EA4eKsY86dqPiPZC6llG98HP81+LPucoS8/5xQq4YzVcQQLkGMt4WK6FbLEA6VehiyhEBe5aHsk0
pqqt4aHy6OcDC22C7Et00ZsCMZw6ZOSc5XWEZ80x7uLAHm6vOhKz/5IefbkRv9Z7TdMZjPF+hMVr
D9GRxIZLn3Md7sSgQide2vRMUX04AANKlxpMZW9bWk/x75tw9UeOvNs2C7Y3wSVC+RtQ5T2VuCsn
ENnuuzkxBk5KQS6pnA+V/xmkPiWLo8yjg8HviQcE0xXzQAD86FyAw6iYtLVQeSuol6ZwGIdooNaZ
0K2KOlj1aXfQgUv4m1ay58YdIEA6eOBVh3AK5pqwusj1eDw+hsw83cKELZXr/dZxDAGgGQYLhggB
o5VpDUa7I57M+XeBV7Ci7couEhsMNdAnenKgYyluuYLUaji1pa8EH2kIrVr635TQnjOIt3/ZXPJi
brK51xpQ20r8tivDwinb9Ec3/qlSEg7jZrEokeUj4wKGjzGvUh64bBq4AI6si51omT3eR+pK6HzU
0KGzi+sEv3330JxeS9iuiYuGSSlLLPchdYJ7ADpebN0R2mIX+X6JLSX7z4YkODQ3HajRmTsd0Mpo
6QbACp8YBpuLgMfAl0HdQO21kAJFW3IG0+Yn2UWdEv8igp/WExhDz8Al8COGyVEHx0oDzNDbBykH
V3Wo3rWe2Q6/fYvKKn3hDeyMLQ3VWFyPIWrNoHk3VYJYyUYgw1HLptH4xLL6fJ2HGVqpq5Jhp64f
rken1O+zuX2RfNAdkVohTU6f/0i+kGSxWwZqmPAgRhaEqfH/TamQ90AakwodfdaJThi3xdnPC0ad
TVU1F/TI0ZwbJugBa84OsijZRKbt/ihI8jcyn6E44I0SUaURy5Z2BcIePZ7zEsSz/JYtl4HZ8G5M
oCZQ6o2wVSWT9Wk/LE1zU9+uL/20Y0C+EShdbl75jeE0JNxLRbNMfbJc6OcvWqtexhgaHMjOKjXT
39Biss2n18pe/Ncfx4dWgIH3MFjQeCbbAGUgVDoyADNGkcCsmI9PjhNOP2j3/NPpbnMT64C2U/Bq
3QvCM12XIijOPowOlP16XZ4ZlJBs2q/kNZaPGPuY4bVdesdIJKN4zW3p/rRoEslnE8p7ZTn77ed/
bXhEBPjs/sFqRCrrIEPTn/SlYEP+O1ZIBbZ4QWCEHYHYxb0J4n4f2N+iCW8IFMMBC6we9NtnsSkf
YTJAy62c8wgoSAveRwZsimWuaVQIVW/t7jRuJAQJWzbrXgVtsQT0fj2k3PRPpY4Kch8gnSVBF/n0
1Xwoa5wgBseeeIPjrCMXAUKb2MLgxKwV4ZIRuDrLsNGVUyz2Mdg7ehEDpVn5mSDG2pqcYaMzxvZb
4V8T7mpq/Wi4aCVI9ky75Tluc4vCZWwN2mdb+9Pld69/tpY60nusph1r0RRIL1A1gSTi0gvxDDLt
q+tAtDEBnfsCs+Oi7JLK6FbJMD2gCF1oqHoOxYytUWf+QdPKCWaKg6F+zQ/G9arT9uBttjvyHclt
DyfIwA5nVPA12nOtsUevp8CqZiPJUGseDgIXTeYbszC9V+WH474ajJgNg4D4gY2lgRcNuGLZ7TG2
VNW4I3881hxQRy1xUkElxGEERq/tirUTiyfWevei+dKIpxwjH7CWgQBD4nVADauL5vD3Ny03MZQW
f+k4TwJTgIpm2W4F5snNIOBn4JG1QOpK6g84UMmn1fGiCw35BZyvV4sHpv4KIwvF411cN37pXZcv
S6nXO1UapBW6XC92avfiVpWduKBvqFGEZKwt5zi85aA2Bhd9nurk51Z/ZrXX9glSfVUZ3pesN1Ca
QwJz0NTwzUtAOdPsaEWZUkYSiZkYxDmTclukiz9T3S7Md7nwpzlYYNJd0d5uIExAIA99x1ItA5sw
QCRIw8FanaRz7Bp1wKdpxhkSwgzS42xwPtKlx4lM2391drX0e+z1reihPrBKnev73Pm8y1Aw2wwy
Lui69uNmVOGSvptLHFlmNq05S+ccq9rvyVF14X7WAFr0pE2Dc3s58Au/cLA6/4d4xgW18cyM7VE0
2KawdSEovtN+f3HL/v/JKrJdj0M+Vg4b121I8hlWaoeOXChT4xWas70eYNiklSq2IAOvOacNfvL3
0gaeANmLHDyeYFynHd/gWcJuWL8O3IOJY/xlY3yShraJq919N733cSezj+zOb6inyvZQfRSBIp/B
2KNgGNSh3SAfZtneQDjC3TR/pTuBWmCvY10YDyrgdkBwu9ppDTw1ucAuLPs4vwLYv6UbvJNsgc20
pLdFe2x4N3tOG64jz2vJlodSFlc7hVxdHXiS2Z46iXa6SxwGi8++grgaYnzNjWDH5HcQiW/hSJKL
YxumX3BMKcryPKhP5Nex54/RJgSSHdbw1bzdqIfhx4h/lMPQPoreSFTZlSKUPTnsnczODrTIw7/d
YqN+yHrlWhsyRjKyDNbSVzWX5tTjfYjQyh+gT+zJfYOblKLAv0FGJCkWXTfpldM0l/fT+JiXkfRP
rdFgReL0SjV7dG1mA0pzrPnqsX8a0xtHJIEnENdIhqNF+hYutq4oIwlZP2VErNTIf/2tZSChoqvB
mxe+cViixasqC8yC/zRZcfLJ0cOsm8dLbbgfpOLwSh/zTqFpVkRultSPvL3CWxUDZgwFvzG0atGE
mwNouTN6tZpOR3OENRS3GTddGBnHtcq9+SucDmlPC0EPF9aoJAioNOtkHEUTY0Zzz4nGmRhCbUqd
UzjPNUhDJC+ojaadaecqMbNSIWSMM59hkpH4X+s+bJ2/ZcPv258qSEUiJGYCLsfM8uo2MsvdPyjI
v80TCqLgJe8t8akEXGjoZbA5PabxFWr+MupdpJiK9R+Io+6QCf2Q8c2sl0VXAR8kT0tVm9yrj/Bn
RHuDCRVWFhAm5D/0ztypLotkynux4B5+S7lcDOvAgXPODzJimUik0nimBH/TIIKosyKCs6kO0EiW
50Kb6GAyqQnB70AZNBdtizNqFIKsWtrGPkkHlJhBwW3TM/eeP4nkn17M6ulh5KC5kij/ZMX6DvIk
4uxsKtneTBuD9uVXAnhMebpEQE2tehB0O7qS+Cmhd8pBb3B6z/jSPz4RqncQp51IIDZCm2DlNPXl
h7G8LYHkaNFvg70reulgJQxbfYiEFQejtt+Fmm6fpalepD7NdqAs2tGN3QYidrPrk9I+qE3seVGw
DN/8aCjuUy+hz/xWP18FMbxk8AemjOc3F6JRNL6e4jsGVREehZeIr+vBLhjIhw9tZX2NWyi1SEGN
4KBCgVYJWQNErFKP2BSeOgGT8mageI3q216qntEir6/V2E04nS3PMiMIpSGvc6M9Cu0beYDtBehN
o2VTrcW7pJ/Jsm0NWLwBxzdk6hdLas8pQgQ+kfbXD5meQ0M8NkQ0M7CBL5ny6W8s5eGOEoi1Aq7y
1bqO5L5xR6/AalAFHdNBUG2ufDOjiyKF60GIIUPm9cWfAWSkAAZr5mvRRXtXGaKOaRSAUmtdE/8P
vaZpik1tkn2uLkKy54KbfY/7QAfy75PWXrXVlASVXM3S9uuI17S857hCNzjmAuksv47qP0skn7EC
yaHMe8Kw0GV61xrShtfsRvElvQ56mOu+pQ8v7HgEMuqHmtAGe6/hdQV9HZ4TsxRSLLJZCT5AzlPL
TxiCE8iDiKS2SButdkLqfNXS1RZkcu8Omjbb+dPLtWfhZq5XALwGcJP3TKrav0SRCsv9iYDLT7+e
zeu4VbrnStFVNFeLNHANIXMYP8wETqCvo1/9VOUWNHZuua2F0bv12clxL/bkpWj5vu0w16Ddm8Wu
prQ2qa5IrYjSlnQxLgPqnMz0J5B8nH0i4+uX5uJEcb6/xKcOm/jtdWSP3g3tSjIDCxO0oVmOEiNT
vhu8plUVeXJkUBj6kzLsPZ7yLIxcp3Acck26VqyDt/g5J2h0Z9JYMuYhYjTAIwN46ji7pdh+qEP/
cMiFXkVYWhrvGIb3DfgIOr4mb4tgBknK7nxOhHER8pJNBy8Iw8Pw9J0XBAXN1MwrtzzGaSyljAPx
4DA+hrtfu0wAIzxB+zekZJZhso3tI/BknPFErvT5qbNtVa5X5GCrJw0FtC+cB4xFpLo2qJ8p2Vs2
XXsyCz1OlMLN2xSgWUoI/vZ/fgYI/cpRi5QNHBs2Y175HkNMMXSpOQZEhQ6u5KGNaYUhxnnfi6sk
cGyJ7rNmsw4VP7DrzGgofTkIGOWbYBjjOpYD8zM4PpZwvHX4+ryak3+6zBy49sfAOg9qNKYRWjKI
Y/aQwXUee8IgISHubiyzhBnokLntLW64DYM79zFeTxHYSB+X0WyedWqEFCuzuKL2WYzhCclIrEzQ
yvRAdw9RlwxcJ7Otc6mxHZ89r8DzB1LFQhrUn4wc+dE9tkzY6PIcXbiM983X4VjdN2MqssaKCMOU
2vCBwGM2mYz+Q/7xquJjMH4oKClRy6Bw9A4QEMpZpokBT0QJ1a3rj5EAM/0FxD12zW8ip6v2Ryq8
RxX0XlRZJcjzB7PXEKe+EhQ91ZsSm7l36yrocB6MAqmzXjeToyW5zCbybiKjjs2Ujb4W5zid51ps
y+ChSepBymHNtaLnv6WE3u8vPBAFRiZxQvrms1FnFXy3zfO53TM7v0/KCEAAuXTWXH02CQpAq10u
XfxXDoOAgX353SrMBn+PAiIpsmo14AJnRkr5VnIE1d0NRMZ1NEeuWXSVynqAxJ2dvvPga+QdrqXv
jmaOA5NgstokwNLUnOrPh6GIXR454tCWNortKy8W9V1Moz/8xBkHaXMg8meqb8TUlFgwcQkyndRO
yAU1u57ZpX3hNlYTJqclmiE7QOYSnQbB5Dt2fRgQYSvLA0TRKUtTHIw1LabAUZ2DJaqzuhtEEV/0
mFZsR56Pn505VqCnL+AvkPp7aoReZXgAzH1quDHvyH7WH85zMyewITb5Jw85N0LN57vmVw8VTMrG
JnODJXMZ5EFNymNEn+yM68vgTDBVjZzyW5Vq7l9PPyxhg6+fLgKTj8gzi50mac3UCJPlJdnjZ4Lo
bJxeSA5q6vvF4fNa2XuA4r7opg21VhB+9ZoELyLEBee9c0p9gRdydG0yRHQCZOELAMmTrAGPSsrp
PM4ZJb6x0tZWu6JlTe283KV9sjE/DP2+/sCifKK51CK+P2mB9MuZKP6W9A17VdGFN1cUJ+o1xH+9
zJV0rWvXK/iI2bttK9BauuAXhW0JY8TTezMNhcRlzitfZGLrWc7CwyO0pWoejEPe1bk+985mLzMO
wG9CA5alFnussHXm3J8vR+opuIZRFaq+6danYX4yVdeXgqw6HP/pQ6upg/u7/z1S1mPAbM3KwRvy
AfXe+ncJdtXjN7NNH5Z53c3HV69uGusfC4WN04ua62g9LidHWigjm7lSpll311IoU8qFpHZPlyOB
VoDF2WSBRAV0ShK6+EBhcdMYU0Q08vdXNecWCFi6pVK+24fGmwjL/pY3hWOeBrU1/M/5miNQkrGg
6bRqyaGtUphtiCircsIhha+OXmMO3NTHl7QEbqPJIOvXR2ndQYFEm6yvJAT/67TanLGyHBoJ3xbQ
3ePqgt5vO6Roll0IHlOJFj5DLLn50Z+fRFwyZYEWKOzG0HCy1neHaOqp3Aag9V3v65cN0t0AR++O
OKc1LKttoOrxrgeS8EF7IS+90fspmcEAXXB7PAovIPnk3wuONAsDwYwSLa19WguUpQA4KDAZbpQ7
Gm7dMMz6AV/wVtUNbh2bxpN6nyM5OMWl6+im1fvFvux6JOnIPF2DgjNf6BTzGTBu29XYKTVOwo3E
lA64UWMFXnOo03YXDPWfkVL7DNyjr3j03ElCFdzxGe6dCynYgF1HwwZB/n4lKT2YpXEBesM4oG/R
+IL9iM2ThONuxRIwnz3duk9R/XBGKMeFj8QuNpI9SQDrw3gfXkQ4RVacFyE7d8sl4Z6rUx5n6Ws2
JBOPxu1jawV9xznk0c5m0E8hutnInaQJ3SP0CKMfHQdIoaZNlefm/5PN44cU79qffVS6Obef0orx
PoiJ/ZuLEcQqsI728qfXCoaCBofmWP6AVUKvndmmDjV9oyvXJcDRhSeZo0Z3bHMqRe8Pj5JmKqPV
6yxRpytHKtnFJXnA5ReZNW/2lOHsVAmGZe6kTFKVhnLiOGLrXumeP/NtrT8lFcOX2FAQgGEUfnUl
ZUU6tC9c0IvrSqMmGTrvYBRN9rEQ8Lrah460XPjfOHRrVkEJ1S/1Cr8Ejk2FO2cQ/si0rTFWvquu
c5S5IzuzSN5qYDuNkETtwpc01WbyVkhPLptYk0Gh7hmSwMJmoc/tCgBM3JP/VJKl1NhIPaja7pR8
omGtUAX3rPIDTERfAP+28mZ/g2Nb23ord7Y7P6Q/AtJ8bM7bL33TXJ7SEtAcGvGSnDxFL0cWt5AX
XwXrGq0EVmFyC/pfzh7RQZnYMtdJX8Lda/+fRTJLD4SnPuWBmG6VR9RpmmoXojocFYqZaAX/IzQ/
n17FVTCsiHr1urHtWoVDPlyWyalSW2Ocp6JQQ1ZDN90vGBu8w0M1Dad6oGrZS6GJvI/2OjE8onEC
/z2PUC8aGvhCyjZcZ+FFboFlHuYLrUS5VqSpnaDFAIW87dlLYVNLB/STv5xwMhav4qKARoRQ4Nsx
l9se7zK4N8p4OmD8UoI8q8QKI8U0qRcCb06tKh8KVh5EfIbqmdWgCNZ9moaNBRghFlnfmKdukBJY
7Eq3yNTBPB7U+H1u9/s2pfnk/Lh6Yq0pnooADUTOJ0cjKLI5NDP2d7X1j86uXAEUeULA+nGOMOSg
pG5O4Z71EkiTeoNsFP9gUXa51LVNcZTz9Z/AyNIy2fJ+BJoA9naw8w1bWvJSr9H9VubreOuSsSYM
qSzwquF/ajYP6Uu1KXcsCu8YhfT6PqVrhU2pMcgPUdrkXHON9v0BHtOJ1KBM9qssH6h3UT1pQCoN
dGwrybwIwrqA1MmUZwK3GOsXmNumGCgearvcZpiGcqdJCoheYwpKzN+iTFMtCAukvqcZjb03CuS8
8ykVSDeEs3B9aJF9ozw+GYS1UAHc0LG2Dhnu/mz6XGKXvKPLdj3ONahaFhxmcSH2vXoxf85kGOTZ
XBUo2t6H0UfeOvIPmljsuLTkTT83Azo8W7Zvp5P1i0qFd6FyIJ1eEQBG/9kyCU2/cRxy6oP9y7+/
w9KLIQMjuOir2mHlSabOwIyHr43mZW9uQDwYT6kuQDvOz4jUcBvNebzRSIHjAKRc33iIsyPBhLl3
3BsJFdZyvId6djK9xTbyTXddmSHPNM3yFUleW1zPireriixn/cbM9TgvIx2Fwsoq3YRviisY1Coh
aK39K1actyro66dSHBntq4nNJeRfZnXsqjGQ3Pce8ZIlyRm3NVdVtfR/HJzHNxuam5bEiIW2Z/fM
ke00UVLim+ZCMQRv4cyTkQ6JnN7ApLFnMdocKYZxpmr5TCzzP0ZwqIiFtV5EEHN2gSnffZuirMHn
21FCuFinl6vd2z0UJXm6uE/0FDMIE6uei2bld9fWOCpNlnF2mq+pEqFWaI4AlNhp6xlc4RSSzSKa
EFKnNksKhmdjPJrkwTDU7HXq9LY5E7fpZ0n1U6Luqqu2qq46LuZj4D2U8MS5XnuuUpqCu7cOi8dO
elzAD4oTZecVE1tHxPzcKoqa22ouPaQjkuKzX9G5WefDv5xqh27fb6h4zmdDokonALplZH3BRnYF
QFeWKnzwTlMxnA1m6dowGlg02qwJVx9wOkGGT/6UjJu1G3AcmmCIqsqSwUHL74tMn5G6AQiAQAxO
rtOaDb86z/u/Jk7vqn6L5JLW6tfXF4kCxp1N2irb4jl1f1dAnLccHLtoVcFJwlCw7Xa6Rz+ahF9L
niED8l6VsQqkK09UxCYi26Od5k+uK+4CIT+dwpyzju1A3aj6Pht2hIpY8oluxqMEYelBXbzOKdP1
ZL2kSI9WvIokvfi+uL8DVAO3wWDuJFJXv3r+Hlc5iy5JBT9fF7w16nohQa/rzmBp/4FjeK1c4OIr
cu/dl3wysZFM4dD7KqFzDAZK2ug7pXMZIOZ2AA88jHiCFUVSV7aedgIJqVQKCg1cDb4TbCWSTjw7
6LndMy0cKQu3gmElvOBHZIn3pIknVoBDg/g5xOdg2p9nojNcoe6hTeYsMGf1lyaLvagK6pXSaNnp
KBFw+LTSUpJ9DQxWShx0KoRdZrv1uKr8Uo3ULj7KKWBwEwhrGCaKjB2rS4SgOzfjDaVVNuOuRUzz
HmnIlIXSE6a/chwft428zT4ik5BAKr7BZ89PsB+bOd7T6geTP1SZ3yX0eW6HJ2UYUlQziNIk0Y48
Jhtx1v08oAd1KOKNwN74CKPAjy8wr1uP2GO/MO5aki93s0pWMl6q1UAXSuCDSg1tm2GQlnmUnFJs
pduDTHPVT8C7gOtUvErkqZv1kc9KOnSRz/tAgpToj7Q0HObmV0c3AjNtNNZzfzxBKxSZYXe2yMez
ZjVmwG0IFEaBCcLCX773ANBlYl6SaZgXNeq20ZH0jM4QZ0et1RZRhXAUb/fM0tnXUBQa/DdUeTAG
w/ZgxDiZn0HWE/UUYCvqofrBpg3R5mBrvcgME6O+LEiBKV55RQHHEY4LHNPWmC2Hw/mOYATVATMm
bt8W/chS9WvdNIIFY7b5O1WitFjl1a7rHjbzUo0w3mnsT4fq25DTmGupNSkMhK8IDqjStMlor15t
QEY8cO5DJAYyih5atWv3mm1efP+oSqylW7L3DqllGRKhE6/xRnK0S0MN5kutsvzjKSwVfJI+aXGN
trSY4l13R+Evh8kpH9IJSn48Iu4Uk7v93TJDNuHpuTqwYAYnKW4a5GfKNvTBDPnIpdEa+wGBCUAm
cwQOYHhotjm1G9j3Xs+YlMPf+dzBB9MF4KJjpyYdGUtVEKO+29zVjI1OwpaMOn84brQ4BHIqt7YP
OCEZrcNpIzA/NdHYVwwzmhjvulLIjLX7tcuxsdWqZKTwc4UwcYFxtze7odxZYAnyfaYffdRdMBi+
bVS5QGkOWCSbmhcJM83OtfzlPX1h2b3HwUzwaGu5Hqcr0K6n8IIDBoSUhRBuJvOnoJClGlUA5BcL
SXUt3ghyu/dLhIsqExTEcIRu2Ih1eD0rOpXXOg/E0jC6IkewqeeelNamPDifBToVHC87VNYJdt4o
VWVPTHlVfaRT5l+bU5m9MsyEf/3nwmB3frVoGGP1LcJjKqWLarejQb4MGEHhWgz/DSdpHfR304WK
BAH4ySuB7troiQ36knHNAxeFZVvoEwdtXmSXo1NKiaaRz55e0cs6pR7Nj5/rb7TcPganjyL8tWpo
bS4U87DguxYR0wFD4ndjEwIBZ6YAlZJ39ZPep3XldcxcNHXVmr+jI3LdwbM4yLXpqHefk4NQpu8G
b5ROpiTCeUJ7Vk7LBoIWkbUwUXsQ7fsNP97Lij4F4//BzkdMZAiuAueDLWqumP5SrxIXxvRSeKUQ
8/nK2YxGpbyZxuHzjY9TPk6Lbxa6AKkBC1f4es0TwyiOjMyudcP+Wj8kZ+He1h9b1WnJTOARgUVr
lFWFrlU4mwztm4hHuG+wThxgvQ834iybi2yerg2BLB4QYdVB9bjq5JGrVWny9bM8beLlDWhrbIFn
yfPanxXHLYCCsAzVJKNdtzOXMCj666I6PN555WQlyALLqJUIKXSbXn1gSRRfgODnNR4CvNWej9KN
njVodGOnp3RYFra+PbemsxjG94nslXs4cYQrEHvnbcMTM8/gIJ3aat8mM90A9MLk5xbetr7pFVbv
OL+jwrAkBLXnpAS2Tnc2E+0muCWZ+AqS9GP+YBaYj0r3DgqRPttZKoxlArLppjGbOPbt3Y5/FX68
NGEdQeoU70kx3NLUZ08ReAC1TT2EOnb7nEth4Rr7ARFSHbHhfhjvQ2XWahvdV8bsPbQ+MW+TcZEk
JYcQTpk+HhN+AUYGyVb8t5+UO+adTql9jgOZ6Jcf7tvH1+7BESNqJMJgIzfS6t0zxdED+Ky7hpe7
8cjfN1ar8400UBbvo2Ak6YPjdL9VnELxq1vOlMF2Np2NqYPHbhCN3bPv0jMcnIn5PEMfFTZBXKmu
0un99v9aSiqsoLKuBvKDGANwxSvU0wIr44BAETYGaCzSgDphn5LDmTazXP3taGDThlhtB++Y0tjr
K/rmQGUdWA8lZehPR65DV/MEvgQyfn36P2DIn0rxEVn7cmQfpD6iEPdtTu+cE5VRuqX40185Hsot
LSxjmQFeSZOqOPO2OTpWwiP69lexzyGEIHPRbrLnx7Wnt4Xf1+s3Ixud1wjH6aci6htE+hjSYCxP
YCvD2v2DzDPoKHW2qHxarbJJI8mc9N6ffZRIlDOyy37KofZ//d+dnKGMU8Q7RPuqhLgu79Z/pv7d
RD3JYDq9GJyUTcDir3lqCTBw8AoR0twyZfNdd+rvQ9FbRbtYqE1j44LCeDsVuVBL8ZwlGm82vMM7
BOmIp/ZhGtdsIrIE+tKVBq3AyInQM2HpMChRTT8B5fOKHYADTadEBC2lcQazZ9EN48bPR//Ep24J
jcSx7R4Rjl45TKwqtATrP0mCtHW3mNzrDLS9fqP53uSeTSQBZ4ru1AKSA1mD8+pH7F1xLfurTwn5
7Th+W/ZsjzS6IMl7/WeuOWkn9yb/TJRFCQ/kE+8FvFWLqqpIctsdnOTMpKOhpdFjcez/wbICUQcd
8sk4Y5wT4sHTlsmuB/7Sv42C8fc8ehXscol7BQQYI4w7sK/CQzDIhf7six0gB6mUqK2Uqqbufdtz
S4ZezWTFaee0vonqvI64WUIQRM4CiivClER/bmokkHtGLyYRKOTjmEL59AOPV0ORti+XQNMWQHuX
GovWb2pD5oa0HPZKK7Uo78q+R5+QbxSk0NokICkwkzkcty8zDBJsVxOKIUKQfB9NV/k/gf1s8mgt
k53g7wNauVGRTCsTE00vxYgyk/80TXtIQdy9NttWO4daZshIZ/Ff71SEoJLmdiqRogbbwRE47UWp
bLWisof63Ku6m4jQXKSTpJ2zOL+5vUYwFJ27PYn4am/mrpJDPL4QglO42J4L09UQO0qF0xsEkiID
nb99oKBVdB2s4CjnodsVNnXsdZB4eGlbVi0H/yiwi7Dlnj62Cl6CafolHANwPttHqH0TjcynEPKp
ySoA10AF4CAXxEt7mqH8AIrI19MEFIVeQ6DWbtV4Qg5rFtBEHYenXZNyy5XCE0WY+hiFBOPxMimv
mHi+XiN9PxRQxegYcFxknMPzWc+Rf8K06ti0nAHd6a4CPYrvD0ElbldCWoCRS5tIu1UOYSULgwAa
rJB8ZKwImSISIj3FVMhuf/WUJSEm+jv6XVzp/rHgO/hx/Hap05FUQgBZrPJ8UcwfqpW/t3MibQY0
ap7LIEkJT5SIglwWf4SNWitMpEXC/M5I+8lgjO6SUScVqGLA+CrYXZqEdi7MS/ZbxnSgTuGf2JmP
oyyeZytQcboEDYipPwyZbBTB6rth4weXJSExkLma3HvJsX+/VsTOgF2LOEsGajZcO18S129DbJYx
4RRiTJnwtc6mqXDg3AlRNkqn4MLQjRBWwIC29CtAiP5oERbZsJoI19vdrcllXN/S8dt1cxhqrTbo
Okcjs1zdQIDMxhAIHRyY7gCps2jKcED6BRcM6UzvRX73YqBpreAyJBuDLSi7rxXuvKp1iG3LbN2Z
OYsyKD50hOdHouoypO7kvqGQtm6D8QJuiGr5vJrmZNYluXJ1U3bnB5PozKWvHyJgJF6nW1rU/Yhq
9/fbYg8R4vv62k00RSzq1FAyujgAE/tCUXk1qUNAFmJ5aWoz9R0sll2k1AdemVG1qXPNP0unaIH5
ApFbF1pjb0MVW03MwhuvNPs39j87U3C5Nrl5ltnEO2op3fwh8DEQw7HeNxvY17JYjOKrjQsF2ovR
A77XuIe2pATogCljLpQK9D8QZjhpui+7wWILZ6Yhd90s0MqvPAv/lLkipGF8c93NLXVRHW+GyPNM
D6DzUuw9hmwGawBGfL88Nt9mhD28y9tAyj1UNABPxthvay/0QeaoIMELB6Ets6ShkrDL2SNC1pH4
FXiLO8BgzQH99LLfUWPeFFLlS24v2H4Es0aTh8BujaplwLifhwp0wiQDd5gVvMO3J2yc0lGHHr7r
44DLBeEW5H159Kcnbsgd71Zf2tx7KftQRp8mow4ZkWb9JoG6zr5+kXI8y1DAQdSc1sklM2nuwnR2
TvZXgCaJRhzcTYk1Ki9Z7YfvUt7LWNHwVb+zP2BU5DILdCoYMnoBq5OkDnhua9QLAQgZsyC636j1
qB3dAYTprR1tD/tyl9APsdi+ATjS2uPmnCnQmqY4ePZW154i2uRWmrwURJdaRw5ttwJlXquqNMMs
TUGSruPcv8txV4yFspUZY+dGU2pj6zNkmyGKS40EITt6WG4I1UtXmvfu8xkvYyoxR+oPSntLnF6T
Uus0Xf5fGh7+nBFsiYnqp2PksickdOZz8hrHR/8KpWx3AHRJoA+hQI4HhTYDyB2i/UV0RxNX1fgY
ETHDqJydWUxCXDf0TEXf+PhhxzZg/ZAZvi3rqvtjzUAE1478zfCW0Fqr1tThZGzwFOCVA40+td9a
Wj/ifiaPfsQUg+ITivTSsG7SWKaNy1Ppjig15R0O/IBkaUl/0zQvd7AIPSOPIT7iZp7dNlR39e5W
zkRqd+JQBbfKwLJKtsywq+oyDuLsX31vLgWQL1Po3jH1N5hifkFbSYJyHjMAnKP4eky+GvniECRl
1Ld5soR5kIvFmAOi4pxjcVTzdrzDnALX9cxulPX34Tqe9keRIpllqTIZe4X/nD5ZhyU3L+RRzCra
etAkO2WeM0HZCohpiZ7ZOVyXz6Pewv0Pw0AsYvivMyTz50ap0NlWWOfbHnWt5uHgBEMXscxowIRy
/SflyIZiOMtflHYJ8noNrqyadtGfH/ujPYQSWuTo437K+ZiqIazzAZ8v54lgOnQ6mz9jfQ+NktEk
DtAZx6bCH2MXHQlX0KiFw6Ike47Uv7Vj1kuQyQd6YcIhPJsN7O/ACizBSMJyf4GXgA3+QXr8u75P
gzUVoig1U5TGUfkSSCMpzAqiBvANy6bLQeFJn3aBNg7oUhcxptNmm9rukY8Z1EPyzWmi//mq8YAP
vNw8JCJJpA8Z4GBnkRCYrNTUmeP37Sghd0A5j2pCB+pz8VcJ4lhegMFcY/4I5wwLiI4btwF8gCLg
TWbs2J+lycjNRbxHlEAAygolNYYeJ7cFtHu5Cf5RKPr4P5t/Q6HY7iuz2yBy/vvzPuu5FRgF9bCd
1lmLLmyyVxYWyjEeBAc0SGSyJWZHnhIOJh2IFa/1M9HVeRMPFGwqBYAE19r5RrNAtvKf5zjfQrBQ
m4vii/iyZ/sx7G+c9SXmU1cijYW/HLbbhrOeUU3lgQbJToAzOeH5EOGRASNlMw2/EwMGhSJ1GZOP
VJLHOV65Mx9EzY9CgZ6posFiVr7kp+iCBcyAFZ7P67C9qih097F83+GETDxcnnWKEEUz9HlJYBnT
32JBzxX+NmVYl9CGam2qW8w2joTxtC16AxnkzSg3r2kZJ3+TrV2svMXUk3Wm8fUBLAzdBiX2yvrw
xwwARdZEReD4z00s64za5TSVlwYXRYhIxKes91DiQiRXsb+99rzx5gaM6IHuY4++GRMjk1WhziUW
vYFvntiMOtN/aB6oBt3krcTiAeVJFdD64N/lwi+DFYN7ERHGUjYs+2Kio5LDKdHBZHIFgBJNhTvm
UTep46OGSef/iyx1lTIzn+fv/a4ZRI4zSBILulO54oR8DqWEPorFMTznKH+k3U6vDagAi/+vxDQG
PCmcWfiodnrCcm5ULCwLZGsR2PKfYgi5ZroslJdpLdQB/ojAMczNRpo0yzCHJqeA+ecR3dJ5UEIO
iJl0uEkYc4pqlicjbzwMHyJAiBuXn2keRq8iW5D5NTvry1TNUByYJ4wlK0U3MtuolMrJKBN7ds/B
x+79e7p9q8rNCxhwrOHtJ4y7Kxnye4ymF9OOc8WL87v0sT2mw5WWBbx6SFld5Gyqa/uJw3oCZJoe
/6WIS9vJAhP2nwEKM69zt4rg15zCbfmqNG9f9FVZjUFZelZRhb1USQ6Hct9pQCBkXssWSxJ9mDH8
GImqU1c7LS1tvwVP7VjWVZV97hIki6uzBCNRfoZyu3KpYj860xE28sLCDC5ZFJw2vuHH7ISwxAq7
uN20hp/fLu+rt2J/uLVoeCjuqE2jSToj72fpsEGKHrqR7WcCyyp5TRozieAuf+GvO6VUtNLhnSM9
CxOWIm7om0sCtngu5JWebmsllQOF7T1vDq3iRWK2TU+7tqq+zhEDc/irzjGEOC3D/IQI4aXC8GhD
jsTk3Sa+0OdZmP6vGQtwplX/slPAXCl5fZljYI5rU06M4opl04tMM/iTy2UT7sFj4W7hK0hlDpZW
CQz9x2YiQlnj5JywBzRUf77AlZlIR5p6/ekT2vs0EvawfvhzFwoWPO2zcDwIbXDYhouHUac27Fo5
tFrUmnDdayX1BohBixbS2pPgbNrtGXFWghcXyBvI7e1zoKzHRgXo2fvUBEwvygmvIS/zoTaNEnGD
Hy5kpzT97o+Pyt0NnWHXPXYfiom6lXeOZOEpc6iZA036tbFVxCSJLJVp3zn4/nLb2rA1eQujE62b
CDBg5zSXhxlMKf722f0AJUY+vOCNvgk+K9WEK2QY1EKrce1jDNqvnd+fV40yq1vd82FuHrvS70qv
f7mDD8gU8Tmb+cJ84GlA7iRaX84MgLiLralTkpJU5f1qT9/euZKJKvr445EBB3+bORJkX2wC6l0Q
zP17I7e/vV2WdTnaEFoXmXTGxACIHVswM9QPxgvANraiKqEPCsrIFgiIuSppSQjXOo+fieRoJPhZ
TNc/gSbR9nNKvJ4/oYxg0Qj8eGykxgqJfXAriTO2xyanMJEXyGxM0edunSOv4zthbt2tcsoE+Kel
LPQBqlXy3CmeLXESlkaKLsOwLeLUfiOXNXFNHrkQ7F1VrDLHGpgsVKn/pgBdT5Z+4XpewTx84/mg
TAF1DMORMSZnWmVDc/Gl1vRCDFxYmr4eOMsspzghv1zU3e1dtjQerzJEWBw2APOq3r0edRg/kpV7
8mrpHecNN6iLVfTZpVIUtZuuSterBi2B/r2IzXjF3Lu+hWZ5oBFg5AlTdCi40H11kvnb3kCtmzSo
fb2+uqj6nImrsXD4Wwf2UbuIbxDpia22oyR+vMHvvextj2sjXmx1IcdjO8FjbJtShb+KrUZ6Wudt
ICv8Py1TlJsIhUP84S2Qf1G531O/5Z5xLy3ukqtqC1TSPKN8ATLGgTFfi+JVj/5O8DpJdC3ya6Cb
wYFmNG25Cup6xeU/LzJbmX8YZa1E/exunhumBBEbsZtI/O/YCwyJ8WN8X5OGt2GNDGu8yysh5rt8
I3HZeAANyDgvMDDRke7C24oZi+t7Cjy59Yx9dltGHsCQ28Edx4trXi0j3HDIq3G1obdrRWhJTyXf
+IkyhGGTM/RfNFqCAfAZURcSk9RLzN9Hbr5Y2H1YcJd6i1kPfkwwSC0UaQp5kpvLM/nOwFcFc55S
D5PxEKvOEqQ8hFYmlwTZ6/wJQexqmxD9zGkxsRFeqXABHGl5vs3JRhnqeKACP3J/4L0H6FY7ccYQ
A3wBOC37qg3IKqFK3+qaD/FCQyzHDQU77sH15sUEzCTZtRibYL6B11JzNC/Fh005TCHmDRQmc1ee
1QsSyBH1Fxrtq9iU7yI7D7agMNCpih86VhKhQ4V35z2v8PTEoveiaYDnAdQX18G86OHRzDPerKUx
bB64mFeO5U/oDnpwK71dyB5gfKNJJUHdLbIe/bn3RCBhs4u2t7dgz5LMX/SN9tdQCmgh/5Q77wXO
LNlNgouYG3dZ7dKQNVf2Hc5pKzJX+rDULQ/RbNLTT62HuUZegqfp8H+0Yqosg6hKMwQqvYK509Cw
pdVdB5WddG5AlrEpXzvd3t3z4YVauQ+zCA96z6TZ+NOGWHB13rC1tbJnKeCwHfFfBMoMi/7adK1o
uu25LYwW8CuN7LclJQh2LDi32sBm4e19MYgJCXbpNhCgZvFKhd+3UHZccr0klIfM+jFOxgMv0xKs
LosIBdCNw/DYKGr9D/OKYDJSJJBYsrgf71hgR/XC7XadI6PcJQzuyehhed1nULrAZZSr1RrRUvzq
/VDrACJHqbeyZ/0bEKfstnl/ry7R0uB854Qzm+1Qb+oenSr5ZT4EBbAtL0l13FEYfLRAx21z2avJ
3IvXOxpEpnXOIIiIvkm8/7Th70yy3udX9Jx4up06YUCZYjqGlDQpeZS8F0/iN03BOple9Xy0lGrD
M91UMq/Hm1V6BFx1xbCpJcDorhdnbUjQ3pbPV2p1eIwP7VcBn1ZzVVRtEQH8XGZCTPh4xGYkYPFK
nBFZD4402E009GDtQEeMzicEtcYVKFsz7Gt+Fwc4IghmfJDeaHzaaWEu9vJ/8ZuSikTyX862Gbb1
8Vw1RL7C/0L7vSyzjbVqYLMudSrGyg24iv9nmpYgyPoarjtHvMPAbGi0XJ8x66KvCNhAuqiDiZMF
ibbMS+05FyJ6mz32kqIHR/xDyM2rlLjws7TBVN4OhKkQi53NVHqzWUMIFlXLiaYT0EUEmUE9yFkm
G5BMIZoFT8QD4B6z74m9St2O3vBvUi6uiHHq5IIhGxYIym4SttHoVGEglDQzNfqil7RJWbFHlN/F
NbvhKf/xt/msFkI8deX2HV2PDgUvVZVgLg2z8AyAfrWP7JmnpxA2kcJ23Pp6ivBKj9KVXVGGBUZ+
cr6pvYXdQ2HvOpzcdw1587NSFjLJXHmLEKuDufEEcludWiOCCz5ZxKvlKSi8LmizIlqS+lFkQBCF
hWMon7TDaX17WEWnBoparFT4GmUa9Wq5KP1XzZi5eZBcEjfLEUTWyBkY6ELiQcD1mU8AKonE5SNY
Mj6Em5njtTAcWUKRChbTtVuBRNJdElt0C9SyqhxwJ6XTrVl17rLqu4/8XhceJtuLvVH1MG2pJ44M
qPSIc1iEi+6auMm02GOpCrORZZIvk96lAud4IfLCH+sDO9tX6d6tqBhD9HYU+gxvpz0Ql0LB1f4b
7Bep5Wlk3dfWiobURKKQELqq6KfMTHNOyR28TuJ2RxBte2FAKE+IRy9w4d0hbPruIeCFe37fxcn+
P7msr+vxapsO2tiid722xIA9PK6DUKw2poFJagtrTgL3Bty9eaZooV5LkT92o4lGNoluju9v1Fpv
URZgfuLDZa29iZj9ZGSvCoChsOguiX87dRZ4yk1dwAwIkrtVwUP5/l7Kbdm5AMpuROsqcK+NzVkX
umvOTpHlanFG5hBRDCQxOoFkRq7fT0SEa2q5S/48EGBC5VsgsGmqA4JjjAUThA5P5XKAdA1iO1xq
bHdUpFYjsoqJbbAmQdassCzoMX+6YrnDh8Ml+T3oQGqo1eMsQZYV1qWfavPU0SjBSAlM0OvXQ5U4
pUj6WSRSRZ//Ir17IXkkfRzKDVgn33xrWk/5Tf1zTCpQicMTfoefskqs3v9vCvfT24MCp3z6xKJd
DKIF3RbO/c0VcVuxjvwLtBmAkOPMYwIJqpDWNDfOap9skyRQJUFeIYbUaJo/zhbfWpM612dkWQ66
GM4z2z4nwIPAhfwo/kRIXjcCzgUKfnc2URNKlxpO8Jn2V6MkdQhwpv4Vf7130f8HBDmE9nfTs/b0
xm8ttUG6nPwIuOfIwW09yBdBXBnzm3d+v/1besNbFUvsMFFmMNJhScXzXpef4lYPPi0KfrHBkjEt
UR6uvWU+eedmTnB3U8+41TfZ3+YeEBWgyRaoTO55xFISvj4/du5dxRxVmNXwYF4TOhkxUYjUZ2re
J9Nt0jiy8x4uJfhKNfrfX4m7u2q4YLjFIo+9PEB+mUn+uMY6cC304D2rV6oZ70w1QfGkjr/NRiM0
0iMYCOExQEKpuEtTQ8rSGhxe0O6FwnfTYDrOswTJwVQmadVZDNK3QBI4ArtP1QLVZxrh4FVcSWKA
am9S1pr16iIrD/SjvDu/f6cSIsAy5GDOuQ0LXutxytOXaXjbPK39LGs+c5E4wOb7BxaOIo8IWUnx
vXgune7wblhDi/ZEj93Ktaq0gJm94jKwyt0dqn9e/IBsqGqI4lTqtsyH/j8vtjerInT6ra/YZiHs
7XdpkTy16gGkk6IonGL8rnsSDTScPpfH2ecB5hpSOazXcXcWjSXiyxFprmvxkv+P6vzaUiai7xnZ
88KSJOvSNXLoVYb64A3RKBmO+9+b3FYnATOjFTbs89CaqqNEo8U/EshzJeMdOYME7n+Q2pnoqAyR
jLOnDzB3+2KGF1sZ2Q9rHvsT2k2ff4OooyM9bk4fO4vbcFVJCS6kn1ZBMpf7MLhulZ0H8NoCWQel
SbyOBiEvlKbzcnwM2RgdpF2oqPYeBKrFQCUmpbX11GgdKJe88nbdRvf+qaE4dpN2nOydc3NdgU3i
Fzr9tfUD1vSce6LUSgeRbpXxrKARp0xDFfQ0j5/XepiyN2Vfdo0wN+9sMxvOVrmY8JOtE7FAB/k0
XhQZ6g9FlbLwVZWYYsNg41GhF5IUmI7R3wxCLo/iiTuWwjY5jaEWTHnq1+jLkTtRQvHbK+YlaCME
BSCUTHXRHM4E3YWxgei5Y5BtV5dQNwDIGC9XusLveuVphlS5sOlAc+Sjhu6WegrA+bjzHZPq+zmY
ZRBOwgjx/FwPAbrn6NTeiN7enwPD7O0mVQYKaED0sBKAiS3J2HZPZpPGh6VZa6CQJB85C3hugq6/
/IWTatKT1BzmjVSinT7Ei/eAaXDLM+8LOaUi9KNbwBw3heEzwaSZ3ar5TfLOKeKvxxT9qlE8mH4/
iGKA65njOsIZXa6UGA7lO5VYxZZCE5vAi+Go7xyZ1+yTxjZVIQYj72ZQpweEtsIg2/N1ETKviIfC
tT4Y1UpgytZrnVmGr7p1J5sZEFVHICe905mwyJT7LXiVj9ln5ouijZy38VDyAq82oxaoATTQkx7D
N3F/sczTG17s15RRIFhl025Sc5cBWihlfLMdY4Pm2qpMtzfqnXms0Wg3zFBQ3VqqwbZ5E8jxyxHa
5eQz67yTaYItfP4xyfBZZZHBuTviSqJG67W73qtAtc/m/g1rf3EnewXpPD3eIai88GeRwbX/htb/
TtruWpVhtmXGgl2BCKkp7yd3FDnIBoZxkO0l4HHwesYUNJ/y2+Tg9nGaziGwYdoHNQBBd0Pc6Q+V
JuH3bLhwkiyazue1mizsSrMINaft35zeX6KCAIN1XIrLY9bRFlyqs1Br4q1/k8soc5YcJbF6lZ8o
jpFFxhjAxHXpal9ZhhOIIcc1IkEPTTIVzWOVwQ+MdLcRtB9IPzwB98GA9HWv+2fV1OsD/FDNoFXv
2TPDsHm5x4Jz+IkqYRpcTqmFYB1ShT+vU/EDG8D2zXBwm1o1J+TZvrRddLvVKeYgCkrLQCeSHTnG
VsawdgxbRD6e/1+Q7mbAJTeph3diylbISF+ILHOj3eyka104sFcCdaEy3apc3jnsOQHCP3TC/P/E
qBLD8V82My7pzqvqqJPKt3hRMWetX9Dtm4jhRCijDdcakUw386pRr0ZqDDHwZYbf6eWmatzj/YkM
ouGRTIb07lZ8O8cZZxPKoVMF2pR31h5OlZaio5yxGUcF6nbS7JnbQ30/b94tOnkh5TfqePBOq3cL
tOHu9nWPKEW1l2NRjbLIz2C5eiOETQ3x0F7HcWyOKeKkePTozwlPmUdICzMHINr1w3dfqHA4fLTN
KML+zKNWyGA5KMe2aHHZXYTXdWWJQTv3xby00JD7o8s4rxbAszhEqAo8a6qQ+s7tFAR9k5OqfYQP
SUE2nQfRizTyGpOPUv+R2nwQCa5B8YYQpZZGq/sTgQb1b3mbJ/Uv0QvTmsgfFZwtKEcI3CXL5MKV
9O9LYLCivaK7fNja4dBU5KgRaMzAhWrMCVSgGFa+xG+S0h5/c5fO0ZJcBCUAGRDJJD6mwLrI/Zkw
pVZh23NoVCeGwMykF8TQSXoAtmNp9BpvZB1r2rXj5lQyFgHnPzs2G82HOMEQjOyzrNQhfX8LTUPI
ML4si3VOL/UthqCLepP77Kg+cowyx/mBXVYzk/yfnW8qaGCkKz5YZYc2m8ZWQwiWtX7EOhbH2KIK
xR0WLaxlbkd9JMrkyYTJuWyLzBRCmuL0MGf4ka+/eS1N9G2CatxyrbOcWv20ms43gqcJFI936Qvs
okSOj0SoqgDICNpfTBquQwWsvp7BP6JRdWBF5scj7Wz6ZDnSNSMZglrDvM10Fbi7bbEBc+dld7eM
gbEwfKlMBY21BMRC1SVPA2u2Sbd5IhNOfuJB/OYJjPbBrp+g+gtsiFtOwo+TIRy40fcJN0wW1p9I
0oJ9xrs5OP9p+GW6jfayUD4dNRHUdJQ2w/hD7CY6nXk6mQwHe0HFE2kF/qzjqa5+6ST1MjtYDZFF
ZMORQaVvlp1IPwBsYsdBH33fc9Ib6TsCuccJ6A0vm1ueBKT8R4U6ra/ifKELj00UOrCPk2UgyCB0
xmv6wrXKFfnXk5TRZr9B3tIZRi9oO/TSzJz85dWizvr510qvbV0S7BG8HPoBeULE/+8SRxU5Y8V4
n6m0UEUYA2eBDLFin0QWNZ5+aCPOn5Dr7L9kAvEqyZJF0Hgrgm/yLoeLqsIdeSqEVm5cb6/vCZCl
66Ul0l4fwHwY+kkMsF9CejLnpOnkBjOJtTzPjmNiZdv8F/ugEMMEbOhCg7edUyBC0BZ5NbmxE3bm
QMTPK3pamwYEVaGnbIzegMk3ME2U7mZDabUgPdw6/du2Y2WQs3ebbiBG72jYfXqUhdOXFAD+ZPMl
Nef4lglBTgj/Q9P8NyNNBOG6lAPeb0nPwIspLGaxk6eg4LjFo/6F9MwQbYK2eQEQFt0A/7ULN/u4
eFWNOJ09hxTG5pMIagkfHTtLS/A1fEtPXtQ1CorLr2XWPtb5l5TDBghq6coh9R/Sqst8FL5bV6Tt
7Dyke1KLjC0w3S7fPrQ03QE2zQ1EmtUwovLFKYiZc7X0NUwmKh178sLLvYzFf3DawUXXgbcdYky1
VR9z4IZClGCWbeGLb23Cj9XSseX4kj0jXmYWsUQQAHCxpsdI4cCvhk8S918cS30g2h91XCVAvGcg
3FYWvGEpgO66XsEV3o2L2NjtPrY/AUmVLDOJHkML6IZ7/nhYT0hl6QhhGAi58M0N/01ksz7gPRiX
YQw9mn1C1i8HXBxPC3mTjgnwNbVpBY9CCY7UJwFpF6umw6ENALO9BMrNjhOQN8KogOGzQkqbrtbU
e+TJ1aCFS4xs9JHOMbjWWfTLxvW94qgwMpn5PcLXVkyuGMQ32+LV79qxCfx+l0JOgrHram9tmw9b
BuLCEaU7vpPl4RF1cxIimY7PLFb6ltfWhx54ebbYJfBM2vkquD8UaF4MY9oaw/edCvMCtGH2wBsJ
Q21/ez+KBno0gnME/ZFsr4urt1LQ1hF54Vq9heQqoqTXTBRxmWC1aOgiU8NxExZLDl6oSTVwnw+Q
ocoIbSD1dHtkht+PF1vr/vIz/cKehXrJVl5ojZHY/OfKXVkHX44xJ38Cf9YwEjQRkdEar2v9zouP
cP/nUMzdntttV1LSPNMHUc4W2ukEfw7WrkGG3uU5EOCrdAHOZEVTV3rg7Jy+eZo7eeEvuDWQmSJn
NTSYklS5MRs0S81X0rjK2L4yNHq2+A6FHWhCsuCtYwBh5wJL95Bry+7+9EGVHy8qyqo8xvA1P8D4
u6567tyjqceGVyzu1GVcJts/SOXrE+3yqXIiLKto6cVFyUZawXolQMyuaLFjg1SInetslCYCvdqY
tPVsZlVoB/EtMWeu/Rixdl58TarSYDD01qvW08OQ19W0JKFljWpHbGYsWFeaE0mdDWYJrIU8qFUq
U29b7TdlIqGPIJ7mcb8rCwd+LSS/JAlK4BdL498RJkGinhmUF4U9Thk1KGln7qv7T1WMLWeq8SHZ
ti7on9y3p/cfd5zdF83HO1Xbb2d+oECgZf70eBgSAm6G5B+B+4EeJQV2L4aj3k7nrGwWZaHhk7U3
0m13czEPFEZnik+riTG94NKzi10/mHNe+KabgLzTLOpEyqJT7u4SYdOZQeyblII1JvN0YsnLAhhh
PFZvhtzT1fC22BZDLMqUV1+arEpVS8737E2aIdXrnFR6TCL/zF8SefTIXhThqoXgnSvkLP2RDfmM
hsD1RGaJTm0aHFeD5y7lbDm3L+qFiJ/NMrbpxFC/l0yOxga+bnUbM0TsV9trencbby/9D1jPGvk4
sKmRz+g6ymXCNWuSK2xPCdf1yyWmaxsmtCPR+yVv10JGtLtZblQybTo5kY5BkNFQzOunwa1apkI5
v4Usd7HN/MPJDPzPqhLCLu5c8JpIJTPNyvMNaQcDTi7EUXuUOY8lmbuODooJkht9PCf/MY5zZApd
SrPlX/tibHavFubywySdM+trOJCE3DHpoQPRSNq8mHnYSkBCmO/jfYO0n6BWv2CwUe0mR1GEeELH
Q2zm463lN0HhEk0FTphugMw3y2xAKBVsYQQo5eMFVGkq3XqfYOI54YDu1y3+bytshxZIT5fSXmcP
+qQNZ5yRoK1zt5eL7+3dAsev0YBf8U6zLnLZi0l3ZokI+1wDArcLlrT2pt5+UAo5NYYyxp1EsMQX
Uj5HoL/nVnoW4Q1bCT2zqMcKSRNrY/Q2YBPcZV4UHQT1IklZ4g1RAU9gJxSKxOn1y07JUouA0XJP
ETCr0ek1K0dNexB5SzROCvprW+a+7jZ3thJxrWFIUxAaupQBz9rlhF+PK2tMiPUQClQ7ILPI1Zab
kSMObqf5ulmdJx0kQwVC0uJUJxbc8hq9i7dYODbXP0h3PY+DFeysjNle7/6/LVMtWDidqlHU/CyH
uq/XGXs5unibULvVM2MKBNxoKuwia0C8FfaCTdjFn7ghFls1RCUxh3yWPJTymak/t8WMdi7Zjh7Z
hXLcJV2RAhXoUUwekuulOokJ8ycxesL4bMLaTLAKk5UH/B98A+Qw+yI2KyM4+CcY42JBN6/gGcfc
Q8PA2OYDNNFHLktMdqOZ5JXVurI8qH68LDXsodXLTIVRHsb9pcIl7EKPr0wo7jGmUnp6/0Bsiv//
cuXBvgjr0g7OVKywo09pqNDX46YnMmYHbJEzJ+QMnjsZSUD0m8TZEw9VZu3fqwC7L5rQ9G/bA6yx
MudtuWfUvYKzDDV6BNhtQT+WLnRw71Xo7kBxTgICUj1zb6ivqqrNdR/bUeQHeiEDfVSONzeEwMo+
QmfDZf0yOu7KuKvEoNMwvUtkW5+euUdVXrYvxIWxkN/amWjfRhOckZsrmHPmMDgpzsRAsa35YnOH
JHvw/P+jlxh5ni3W8Nt1leNDQ8Qnkul37Y1vQ3ymcnCwnw7snv5gHMsiXE/zZk6u0oJ1NnlX6OuM
7jXLaISSx5u4rUIYhtB+QLNefayts0bMBGDgpoq6TFvOcTL2KpM3cfRYBthseideGCJNeJw6UtHU
BkWD7pqsfnR40Z2CIL3S9SBDQB0NRFefu8qAq9th7WS0XluBQIDCFR4Ep8g4D8fmkTw1hzvfluZ4
uP4VMPxtL3PPdpoTrwcsVY7no2pMRbv+aPUITkPwqs9h0DfDVW/0JDp2XPU+7SBr0LdXNyCkeWm1
wArYYMPrxleHk7uWPf4nutoHStHv66ZY1Dgmj0vT5wawOAwCBT4ilCfeXSijf//CwZ/4R1w3pBQX
iYVanLj6wkkuz9fjmIQmRYoMOUAXMSkLzJ+0jnORVFknEn9Yt5CFl5EAyot8pq0ONfWXs2jLA1w9
3TjmKsfARoUuTAThtMmzrjSKSdIDUfZOuDxE0mmV6s6wEQpB0F9V1y3UFIO1FpeRdDKOqhEzDeaA
ctsSqRtZ4V2dm9V+Acqy+9xYdc6XxrofvO19swlLCtp1dnPNzXIjzVlW2eRDytLp+8BcHYxHk8ru
IF5Rli7DbYR1Rye5T2efSoekJc3qm6MUgIjfR6dV+hy7NwQKdH7MvGCxKrPbqpXO7r324Z848zlQ
d+ejKr9PtayBPSwMx3NndZcovftbeFL2wNE/KwFJlUfpecM/SUnSAJ1quDYtnQMHsqyqhQSsGIQ5
PLLiMyquvs+hH2qjN6hNuU+Mccyu7AZKereXf1S9f6svSFRhUsWd8ICIC2RNjWsh5bx7le4wuyuC
phmSGayig9pXE2fIK7tZ4f/mFsPUyKsu3t6xk1tgkF5kLIHgfXq/Mkbo7TaWjpMTrhGTXT0C/IAj
WuCXmKhqRwCrgfJpdSUnrGD6bMkeI+8eixeru+EYyK5o+W8bGn3EUH18u0PyuaNUuIKkMkcPo3+G
+7NX/4PRSVzBwunuLOl70AXMfsT8TKierlD65DtCeMCtgFaTA9N75lS6JfTMs5ADrYVo9Diu23Ie
BO0eL3Oge0kbjsnpVJwpO9AOGZKdtw9Sf7hMkK0VWSb3rNadx0bazRdN6AKhWFnFhD4UqwAgJitD
Gndome2y7y9MLMHon1h3TUqHO6OjSBWL5spFhHrBV4aFBw4KCWrYSZfd9XBw6kti0AJS5N8D7Cm/
FnXP+NSI8XOQNK1y5mp1wq9fE3wJ1oM58+33aGJ66FivflNBOf5CtfYzdaOzs8ufZwNCnUWYIKAO
cX8UH3tzNehTWRLZBWxx+V2wgvbHRzAljQ83/jtZrpP91J+LGS6qMmqHMvizqJtO9PEhMfysTmuq
FViyAYhnsTKqwzwEH/tljiW+cc58HP+M+6W8bJAha06L/Q1VkaTj5d6quDKEZb1pGFEjBjF31WLv
yduLlD2ADtz+8p8shG10t00a57iRJ6/YMu6Wp8h5pRkmQ7m1On7FGdbUjL6YBJ5eacY1U7PHUgbu
Sb8DKAHNRSUUygJEBHnv8igFJkPeVU3FcTcPkwPFR+1izmfVXC7KFoaMQsj5v2+Li5UjbopEjCZV
fZ4TqRQWQhQ1ryQAOFBZ1cHmfVhkm/D69qDfvTHKgMf35rMvhTiS6ZUmmK3+t+8Gb7Wllq2QT4VJ
JAAmMUtq21ngVY5Ow3he6kKjhzIazY9z7iQVryTURhmzYe7YtaiqPoWLXcjUL7JfEmvLUBfH8aV8
pzNZohPW1XbK085/u0g2PZ7yxeiC5dbVdG5Q/1J9eRqrypfd614ckzNWfUey6/9JpbduLpkLsSGK
/eGa0kD08zn73Jop6RxZA1i6t0/qr2Z3wkT25WzNjbq0fuu/V0wXVXY9cdrwh2nCBhuw+NclNltA
dp3Kg9nxGnYjv62f9DPXTEXtOudL/J9kuXyJZeoAtp+IAxqxCBQfSr3qmrHx7jjqHOcUBYMkKEhB
ERi+WHzeDMxDJL6/UGRFGoifEzzhVKASuEza89WKbDEnW43BXFA0jlXzsdRzl/inAfnARKqAECb9
eBaCHOPRLAKJJ4Xxxoc8+L/qmBsMTTaCUszH4si3AUUdJH+jY6Rw4psJ5cnK11Ac997xXffxKb5i
zC8vm9xjGTexUDmseccPhLS9F1zaW07a/+b9dwUrYOI4MiXje0uBU03t5Sl55IgK5/G770VavY3o
EvkS8Alxmqvu4JiKnpKBMW/X8T9aJE4gK2WlcoJwuF9ReggacpoaYOJ125BMBUMHf4i1yz24StrQ
TsQrApMC/3qChFuaB3WyRk8f//2g7VodTp/J9epnWTyBaCpjVyZ4qYcP47vI29Djv+E+39okoA9M
sSkVe5oWLNXcaEjRjEwyYAIwlBz2RgmEuMXo19Cek9LrmvL+r7KQARvxi7S+QHmehaT50HwrpW71
o+gONhM2qv4zqCz7I/PZukbii7ZeTFR3kZgS91Z/M8OfM/hCEslltUHJjbpVCFqqamltFL8uD6RL
c5XG5Njkovv44+vPSG+UFjnj4G3kyfW6JWsBf9gadxSTOQKT/RnddP5ow5G9KW8wC/MKKaZrnOvo
bVmGuixLBG2JSoO6SBF5o80lAi/7ldZXVJk9lpNVWbSmIVgjApBqh7u06qzT93vkGgUyEj06YSLw
05S5Lnnr5PYr0WYnC0rSF79N3uEUu8WDTlPgULTQtG7AQY718RB7DKdbgcQf6dEWE/Z+yu76JDo/
JBZlyqKxlUa73zM4uYK+7sGM1Uxiy62uKBapaRUunEA2Y2pjvGiRLfQQh8upl3e5Eyow0jpEg42w
xQMhYO0a9gSlO5X/U+ilxdW2D/pZy/GIY445CRgQH0ZjIj7iRTdTK/z5LRZ4PaROzODAqpDswwPX
eERL0ay0XUrNw5Ivwi9RpRsaG/2YWDAtL8cNuLiqckED7bxq2X0CqKuq8SyhXktTPfsTW5kkVVEK
n+N7slaYWFJ4FNkZ2CU7QiGKUuNXXQaYMD0rxhe24yT7+evQ2iny4n9fQx1sCVgMUeOiSAMgCexE
sR0CM7vOULBDGeGdwvH+SKr3ayen6Qxc5OHFmbF6ZefQ9avcfKgYc7XT2DTSM0d5+qyY2Xj+EhJl
Ix+3iWnkiFaXU5mNov0e0HE7lrwFTb7q1gaDypMA1TvdWvvR4Gj+Thp6BYi18/kqdmsQsmr6M5X7
/6U72DQwwSrWCR0kPc4YMGYLyzx66seHkoEmDGjlp/FJyEjrZJIbIDGi0wfiptxqXZyy+6pyqy9W
OvdkmJC2PjQq2qmAcjbKX+uY+XT4hbRimT0VW3ax9ZRQh0lObI0MsdoiogmsdwQS04dyKu5IqA7r
TBG+oNASH+SL1B++Y1R1iOzTGvZraE2OjosrjuXTmBoNT6iIj/7oyNGvCxPkmaIH/b0rNbHVeNIe
icgA9/uoi21PoDCqCGB97DOBHEZEk5fCdp3MNI2h4Q5ZmtX8IK7YiBqmZYyQ7Ew/bFxMqx/xKfVY
1Uc2hXE/iECO/DrGFDYdQOmswqJ6xIghuSu42zspBI4V9twnwGetaCDXaqqlL1wx8bNquzTqWNhl
FXRBe8S3d47CuQdGAMGYpr2GXqvNMvzLSLiwhzy0oORMX/+YOW4ZaN1lFXm5rONM9rWckOSPZtyr
7yAgZ3KYsgHz9+rkJwCmjnp4yeTd715sN+SmLKQzGR3lAV/nikvsN9rLK/YswXkQfDZybg3ZBxVn
KoQvsxKfrmSr7jgsnFlfXCIG7ahMmTmIkCh2EFtqZVXKMvQqnQ+GM+8zDQQEHEgzU/nBzSPuR9mj
ZJnZgTJQyFF30B3fMVpAG7VJQ3e+DLjDdBR6XU2RHtmws0FcQBxugy+MdsQxaWDk0z66AZZU0Z4z
lX6AOpGbapv0uT+T0jurn03iQSghxg0wn1jSjxqGRHdTehL4YL8xCKvQ/Guiz2hC70Xfoqk9sa56
DNzpphbpLoJKA8cAwpoShPIARjyOJbIsa/izcliS8nN0e7l3rK6OgUf8z96t9ZihueX62iKYKfMV
4x7H/V/1kcl7ATb3FVorFs6LXqYbrblbUUjmvf9oduldPBRrLAwMLCwCKFDbivR4RdlSQ9hxTuC5
nVl1jRHZAvH02Z44FD/UGQ83oqaQuu6ct2i4neXpYm92uLW5kQHnAtkLv5pSD2EGuC7A4M6vcx4R
E7/YSFoWvPMNhNZgT4zlzlkRBd88TJUEwixSwkhFQiuXkafa+DF8GuzfnDySHBDsz6YxNFf0IsEG
KLEc/53Pocnr7J2THy4FD6ieMIx9H8PSjmVRLpQBpR/I/sd7DsqesCZaIbvsNPFF0V++1ewNwTZu
iYR2kgwSWt1nm8rmMnl3Ev+CusGdEbu6piuTR90a2KRvj0tB51cXfWlrWr3wAIpwt+thdF4he0Hh
x3d6dIAMgRszvS8NtNwqoGJWfGBLkC+/pp5uq2HCjQGWnVkhzVvU2363ocHl1fexb6WXEx6Vpwm8
a7BmB2pnR78bPWXgFXkC21zfzbi9yHo04ldykh25wqOPWiU3m93QQ30vW3MH4LfpV4WA1HTHqU1y
/5n3CK3khflw6kiGtMlOX1Uqc4HgV3Bn4YZVeXKyTILmzcs4rNk8avDceImAD2rcjdFo8KAHx2fW
Kreg0/o5b7Hc6EoC0ZIFKOBGVgGhVioJwJh0rmVdGThWP741dqYPNm6xuvqHI80QAYOB0NxGACCD
aUPNZKFkuCYuDArfDlBQEnQadsWGzQ/ws38bYbq9KT5KCGUXHGABV+RKa2WpgtZ6GwGBYFzJcqgq
SMlHipoA9K/MGm4Ge6EUzHpvmg/ZgnXU8X/mLnuEDthG+UUP0JYD7VLSThzzLXCqQdQ6JS1WQCzP
NGEZPIC0j3fdzuzvZ11d3g1kRmVr8DZ3Z/U+/3q+XnCIzC46u3GLKVt2ffs2TcE2ZFFwhaoFaCHk
0fin9Gfpmb/sjU7E5KGnpciFoK+DyG3Zc4K+98ZK88VwB4AZe2/smnPniKrGp2s0y6pigY3yoncB
+bLmh0lAk8IfFpjbz/WrJw2gkDFKlqARRm3I7JkxizaTSN1KajytAVC6fkgqxvBepbKmJ0JClQhQ
lGRbmkFmcaebYb8FgAu+wJgUdYJketMb1FhMx/BZ2PjyGVYXx1e5bI8AubVjTHYS2hQbtXj+YPsv
m1nWiGU8A0kvmmagvoa5kYWjbMMzKFBZz4YCVWxpjpPmvqzEdE1V8szzqAx64rZWTOmQRyECywSW
dnFXK6xK+DDk/efdgOUAeCSXmiy58cbmtuorN0FXhXmiTZcEUECvhPXuZlgQvOVghNdu/ZsEtTrB
Dusox9qBLEUz4d+3NJ3RAxegu5+Y2QrvHKohYQe9+teieQBpr0Mkmw6+WDPUlFX/4h+ulS7qmuFK
4iJQosbnNUVhm2LHERwRNvamdUX4aXEtSWvMMbPOxP7VYt5vt0iq7HF8XNYqLREl+qWwT12ssgp1
+viW8a6WW1EW1u55s2yDmLynTR65tQC14oYC7HLlB7ZXkuvte27/7ws2ls2/yFUf29qZIetGE6yN
hFj3XL7qy9kWzpVnDnilo0WGtGblj2z46nObJvpGp7J5/yuOri5cvQ/SFC7gn0WZmzcV8JatKSbR
DbLg++59qCA5lXRl6MvsMlCIq6LfkXYTuzgDtdVZu+IS6rcO7Ffrt82CgeRkOPLsfYVTPOHDX6/w
5dGGqmMdgxd9mFiuyTP2OMjB7QKTQt/3/AC0jxErpxj+U4RySdMxUe2qGVDGD/LM8VK7cEAbsUcC
cO4RAGXj+4zASyvORgYGmBw2E0N0OqJoG6nUyS6DST06P/du4AoTJrynhbuHtcjsfhNXnrQYbdeL
3NI2HUF+7zDrmkGLVngCT3S1sksEbIQnzUiOLXAbYhbL3TRj6hpXIqiAMzAjIg0np9bsibmnM7AU
/PIpgzegDlvhtiEWxs+xY62uGojvNNB4lfCb557kU95K17km89lyUjkxAGubmguojLABTesvWR2K
iakamrZGtvJHku8o4ryLM61ut1VZMdJPqMvTDR+ftGaiYiYt5uzcT09HYEJqFOeTJj2JiLcp2GFB
dVf+whp1tEe7YZI0zhDghRgtYnD+heOExW+PTA2fW/KV3cq9LKtup5zh3MtpNEBBB45pJo4HcSdI
P4IHSNYLn+Rslvg75hIVkq2ROBGF65SOXi5m8McN9Hb3/kCe74SzAJRaBB8k4sTlaMJFdlIo6SZQ
cC2ekYcy8dma7OVnumq+Awcqk7ZeABGkhni0rAg3xGu7LlViq67CQxsRKYR+q2ZZ6jKPt8Dd4W2d
bMytdrdGHdLPM5VTJTb1F0CQ98lkZvrf0dZkRnxjs0k4rOIm/cjwPiz+q/5Qt3MxaZNDw1ISWNDz
UTmuFNqck6wBPm9SWXhik5f5pX//jGYK8SeFCrLkKzxUyLep4fCNX8GtAYU4fiOzuzvnfNuVWqUo
IymywewtNrAndsocYVkE9lEEL+hCeD+Jid/8kDNqiTFmMsGF7+XqBNXn4wXF6CpcoU/1aA89gTko
QOZzlEjLPJvrCbKlrWBTPcLLtvsKVqup0MiMWqQysMV/AeKoESDefaWAOYOiArneD3Di7RowJ/CC
rAWGh/uZjTi0NKCkJsiyO+vzZGPgzwKn51D2g4+KLjiCClW4jVBOKC02hOIYG/NMM3HJvrteCdg1
7EmTvuOX3O38pWMEw2X+4AG7RROYIg0qTzWU9Ueh2ozjOOqYnz7iiw7yZzkxmn3CoKS+mL76r9eK
RuVI+uILRwxgoo5tPbXJsL9AVDdOTqrdoGQfb1iKyXhqvgGo6yGynJSvyhNy8hpn9R4jBr2Lp9e7
94g0OzuB9DeSdfWehGaqMvKXl/izG7ZVeYpWq3NDW4WMLswu+PXI58ZlzWfEHbHDVj4j+8q49vVT
OK3YaQKNnb6EjzEgisKcRGfF7GPJpuaVs1sOLkJrK6a8mciJJN2GsBsP1ZYrhv+o7ImhRlkcansl
wPqdd/n88XAJJ8vNrbjuplyxmw1n1lBd/kaY1UiNwVDLLxAMmbxH/sXDVrM2ESd86BFuB7jtKNPA
4YkiVslswqLjg3BinaeaEp88H/p9ZvXVdIbepAURvc0LibTyuOVQ9x7VUg3f+B4Q0tLgoXOXuGOs
nmHL8X+0tOqfJk1PTbJsWuzdhvsjk+vWgokFSmB93lCiRZIYzpt7d7mGQKQ39Gei4ji5RpyVf76t
QoNu9uIc5Ysm6bqNT49gY97J7ry/CzP4BUUAwz99zRlu3na4misnHvHNt8DcOgJvl2omgGVkxkZ1
XO48ssgokSMkA4qnIzyZe9qXXdK8jvqv0ihTf2IrouSVjAS5aNfeP56v7Z0wQ9drXKimgmBACl4V
G4DOKp9Tf9GnzBZjdMCV7MI1l9eA6YDboa/di25UVdukYcCIkw6ms3Hv5s4cPOKOy8cT3vpu0Lv9
A4wM/6ZZRmrdR5VbENKX5X8aVg6D3T7KtsLvOGritIh904USZWnyHqLOBuQaF/IsnUpJz5/zCinN
Pz72yh7rwcKSSfH0a0v3g/2d0UMvD3TKfHEy+CA7X8mhhlPh0GJSJ730lkO3256SDQQirVmsNz4a
/skIw+95I8LrEptJiZ/xQ1D1TeWfRlMsQCnULI22oiMpG8WpAQgwtC3xkup8itIY3q2XFopt1cFa
WijD2MGXJreCUhaiv5TfEvkNZvwiDi2g2iy2yKQThQR7hbIUJTtGwuyna2/j2zRaQaE+cqPhEfUs
/rHkENrTFbmPiP188hTpn8URTIE+HvN3NndBDFPE9hqt8+a8mbLsmjYM5VrzOvXrf26Co7WYYO8f
T9PPird7YmDNYzuteqtGMswwJy9KCIHGKf+vWHhg6dmCqKXfa0gFrUES+lVAQq4hyzxWjbB6KVhK
hRV0PGZYWU612dPKAyXL05H4/8w3p7Dn3sRzarevv70qXSkmAJowH9vgDEP7axvPU8o7iKHKsQy4
fcusrsqdDQV/em0GZHh0rpeKmqs/9s9Os63vusrBKR8tVe1eWxgd44sEofkJ4KbRw1hT62OwA057
lQBcbqRw07tqSu0AU9iy67KQkJLPkkZlQmQ/VI46wrecsyRDUXYHCzLBofexQvmkp4pOT3lb4eF7
UzNO+8Zo3Ws+dR3gLyfbYbJU5WWYk4qF05wI59FYW10cvfAUFyH8IDtU1gC3BTxE3BQnfM2RSt6b
HvXi3fca6ZyMAJ3Cw0Rny9qflNy1aQJzec++wEW83/CaswGRyNDnNBrHCgnKCAH9j1DKcZbBTXWw
MqF4WSuznXcc8a3MUtiB8e2ZDYzysKwauJEBJGQMUPP6gHHhoUE9/m/g+26FosN+dzc7CZtucp9e
bWVI4tpJsm0o+5rdZ3d31ppcVZ+IRUcnyRmtSr8b1OVWFK9BmO+iLqxgNHueWdoJvQSM8JXHWKVI
3mtCGzKA9vFbvxkGHeWIsWEPo/pWguFFIOpiH2ZeFFwEX1FrT1mxwTVO9LlGYknntwKhGbJ0ld/F
DTTARXzYK3dMKlsqHPnJ7yEq1jR8YtRg/I3J4p4DKnvNbggPT2sEWKXF8offPrAYFviOXTFecCrt
aKTh22F6qzvYwnYI0ytZNl/cbdulgbu4U4yCpsUtI99kLX1anjQyTQfnVE5XNjktTBrB9QZJV9OW
/HE/LxFSx7FBgf4VBIc6YOrek7tFt7+Yyq+xUbavgJJxqMlK1CMQs9DHflJxALPFs9hI54RyYBjJ
iS+jxC9UcUxm6bv1nS6j2pxnEsvPJVCePQY/QWyZQy5oBNPnpu+pdesAAx6t7QbZXLxW8aMQJ4Ju
XezVQBotpd45O82fm9NDxtWc9zTsLiPp5McSMKpnfcGLsIhhePAQlscONb86RAoTSbou33KLgW5L
8kfzW1c2u9gHJc4ML5O0rpdUSyahThuYqBg7BVpVF3JIdohc6VG7TB5UtanFRzmvJ1J9jx/6tNF2
kMBCkv94kjraPkZtxR8L0Ho5/PkoTEVbT+se8mtiWhq2N+Lxol3sTGI3lX87sgVukEOETiNgv3gI
YhiuIC3DbJLQmgMgxX4Hj7pI5yudW3JBAoZX7A95C+u0slkViX49fkO9uMz70GlHzLsTsXYfTsFU
dLTp7TJTiklio9vwYenIKdRn0h+/0rC0PmPvoReegUvYKSXTjJI/c57j2aKQ7z9aQwjDdH8SRmlA
0dcWpoXnuYAZpcMKwCS6CvlXGTQsxZbJAjYAXasXw2rxAWrzWCztHcNVkYX8pHYp5u37RXTTwQvz
R1uz2NsrI7Pa9qaIPQTdYiH75OKJ/tZkIUJNAV9Nnpd2jYpaKXk4H1VYZOjGvNKBwNR/n+k8PD4s
GhhLKK946X4oETO380YoorbVGe0iNOynjTKgvDTyp8rzS6Qu+sLAxukp8lWFRp878O92hFpTbKZA
PoqI3RVRLWDd/qT0zyKx+e9iUJuzJpAGQ7mOR3KYAypTbX3Bdo9pe0eDBVMT/6nC6pVYjgIEvJC9
Br5h3HI8ZsonTfA/9k94IH15IFwj2vGsP8E9jgU34tD002cxrasoD67egOzyX0du2CnsdKEAw7Le
oRYydBTB5fK0shtb4ap8ld0IwhvvFs2cGPoYXC3NTRXhCyI++zO8e/dphK3pL4JvMg5GPU1pQKC8
HKceKFhl+co4Ix9JrLQVwjcAaT9RRJoXHzvobrQpv6sUQZGQACrPwtceBPOzw5HZiif2E3lKMOK+
86SORBt4Gy0GJfTvStHzQzltv2yX2JD4Ytm/77Hnc6MI+Yjc8gnSUp1XK9NS0NNRHOSSZsy2NVSA
Hvx42DJZjfTXcz7qdGyypaaLmsy6gfggve+oPDJki4jZPoCK1O58pETWzeTJVBewA0TY4bKAboUz
U6d2OZy7cq72hLPtRNn0sEAzk/TNCErPCfWJgm/nre4Kdu6xujqO8RZ7b2TFNyE3QkLqgr2xO9Og
SIIXK95lG5RhgBXs/VACg77hiorj2A5foFiFzoqpO/x4YpgsxzItlWVAvsJXmVrcMzfd1Bf46m8g
9ZTMiPjU0IuNZsfZZ3pHGr+w7QVbA8jUYoGuQzfd6mnXuImF4yqpDO/jgm09wDim5L1hyK1C00zW
O4YmCt7zAVuARIFVDaTnf1LCmKRd54Rau2jf176/MLVif0L+mp2qD1aqM9zE29ABoB36iWdPvEGj
QbHGcfl9+GgWH1sk+jO148hJkERgKX91J/aYWEqoiPi9NDWMfACjY9ZpoFzx9lgnSVYgF/+K/+WJ
HE1ht4rK1SJCWBu6LhDcOmWwZS4vAzfZeV4Fe1znTzJTX6pugFdVtYxWuS061yYKC49oxHMwsCRR
xbTw41TBZff4UBYcncArwCqdxGbEfaCQtnwJWyag1shx35tCT7F/+elDI7ckVj4MCWqpThTtB1Z3
Z8N68m8GRmktgc2bnL7FBXT0JbX+BTShtmzeCy7S6joGmMk0jFXrAv4OCEFGjMDF0guHnVa9eZvO
u1AHpdFEEmVIgIoV78Limd+CyY7eFVFnWlu2KkRBZ/8a9SmibxMFRsXY3VQateLXv0dOjfngQdD3
vZodFjRqmNM24V48iREujALiS0lVQNfCIsDCPQ99MBxfBA6pkMiGQVUP1BkAihKpse/hWFl4+HDU
gPD0rtbbZGpXdpmwo48Alo1uUIUKcVp1alwaIgyPrOjh+cr5gsq6kKO7Bb0VyG14MDtm+ev0ACAh
Ppe6z+tX1Nu4YKlyn4vTmxkxD4PgNEoi5wlfwQvjWxTKIUBKZM21qGKJId4nn28wowQVtuz7iWM3
YMjVI7Sj2M0Lm/wWAFQ6cU9ZS/7AI9Ea1LxyV6dq/Kv+K5xu3YdeFedPly1NFynwV8If5RCofzgp
74bbbOzk7ClXTZGRLz/xXIySQ8iTlQCgVcpGZ6zuU6xTtYtGlMjlgXXXRbgjFzSD13mi2aqoldny
PwZlTR1cOXh5nGnQUTWtFMaYhgK8eQ9Nj7qvp7i7MHfXMiN0Ckz7/J0D49e8WqIBvH3EMVIY2nHw
ThIN55MaOmY0+cV3WMjYLMBboOoOOnxK/+6ktR4AZy0yzEimVKUILY+dh4yde9ZqStYFEh8X2lve
e1twjoyS2qW3aqO40ll/w2gLiPu2LGOGBIJBCdRzXjQwLws4EYtPEvTwDtAcNPBJhYJOdmkg7MkS
JwfMLPuGYgkVTk5jApQAJFm7IYdqiLFrXvaUzQDwrWbcDBVou0jh5hXabtEJuy+mB3CL5xFPwNWH
uwtAX05j+Ifj1/gcxoMrXcuEHL3yNzMHuvF2+6ouI6/XQeo410MjIYwxSkv/0wKekc9zxHfgGYTC
6MfWL154ENSxr2LVyPH9pBccpupvaQn5uOsBxoAMOudWsXJu7RgEjjIn06EcK0HA7LzdM7MyDUjI
GtLUDRMBlLf/+QLo8muse71hthh72Lgb/9NYDuh6tkZJL9d3IwLKeugA9AUD1ISfrJTnARP4doFB
uSvv5D3ndtfiAAjYvPdzjv9tyIPaaxu8u0HCVYAyKa9dTUSORqeE0+jyVXEssNmuOVAmehouRfo9
kWd2RTER+QlxJqgPVDjsIcIbtgXU8SVdHiMCq81Bw+b8uje39mWOMo4eLdI/1mxcQT7YP06SIwer
jw7GOgmHnh5DaJ7fflbuGXMOshARrauNJD/PlkOXftxdshxHXj0iKDC+MamCxI1KPh5X/Xu7LWZI
fn1QiFQ+UUHPHQLQeM7YDvjfLnIn7bdQtsmYWZLUlaFKvoaMGQKH2drEWnmOwihRNtnlDE7gKz0f
VF4aDRWOO1cPOFXLwIyUCh+yUv4oBrNPAXQT9iacrlLNfbYt9IpDjN81JO/ikVklaR53BSx+xFNw
tq/JhuH6BxD6idr2slS0pWvN4O5muqslgE92F4ER2XA8ztggsTexdPWfuDxRlziLBFp9pYHv708i
8qMJW0EBHmNcW3qq4jazYozfbAB3rrlyxc4H6itJOvcDgbJ/3iE5xC3EI/K+TWu5fzNujG1Sz9M8
zhqCGKk/BBKS2L68Q4Tku4roJcV0O3zQYZi7/6bhKJWi3vtrljW2mraCeBuZhXKfLc+MWiBa6BeA
gvb65x0S4D7+4mHTihw+5pwQ9M4Kjt5XqXMIWHiQQrKOOKl0562lo2zK0Y2bxq/N2YgFxYixMcgX
c+v5kfkx7Jcips9qxdCWYvS2amDupcGxyksZyuUpCMLDzeqXE36VTPCM5dSI3qnttE6IlrHJavNa
hhsoh2uEw4rLTGbpCQi0GarkzVgn30vjzcvMN43KDFBERN4I/f6l31L21c1UPZkdLJtqxTfiVSjf
PoI6jX9qu3tPdMtOc/TxWPWex10F6WjUrQi1sLPRwu7JA4Y2mL0nt/bPMJuMxZpEh/n99i1sMgeF
wSppIfjlteKLCuXWP3IS8xI0Tbm0RgkGVbgB7xRpmkTmN8PGynxOLjvJqjvdFW/pLo8di0WNHlFD
SYRrobAzVs9EtwlkPNXObYBs/9RLc5gAyo32EmJPRy4MSEYs/cUXY7UMsoE5cuOIvpk5QWVuD7Ky
Y91nUN9BepKc2fm6Rie4AXjGx17+bnR1t1vLqLMByTXLkRMZB9tqs5smVlN1qq1Q0dnEqaHS5w+w
YvNVnBt4HWtMU14YkyVHuiD13Zgj3ZhCO9HaZDAXUwZvFtYDRvwJS6ZtvLA2HmfCZ2DVs4y9zbDR
hbd299p42BOb46zrMlmpnTiVYmMQgoJQFoo79rrZeEJDkcu/hLo2pUWSjoCc9DVaNRTwhg3OOk+f
I4iNXfVGHQ5BBEdEF6yLfQuiTkFn7V0i/waLfxEKvS0ANdF4qwW1dcETRgVpaG5eUXJatpaJyPZ7
KjX7RHvW0Gfe2SxyMZ3yumoB4VCS24oLPsc418OEmFz+8xAtz3dvG29VDN0SvWfGYrdUd4AJSgZN
Uq7Chj082HqzAvoWbnh6tOUGJTxhfcSs7R13ecuA9z5DVN0AjEQBIxMvxhBG8df0ko/10grP13c3
+cEcXw4MrrUZ7OxpGwTUWFknpO/uUv61gUHRbiZegVjlwV2+erWbb7YeomJe8jZQHP01MFzZ6XDe
9JWEuv9pr/5jp9HAJDnTUVEdtjJ6gWal6lTbJpV8ze8V0MZWBd1Kzlf6Yx6svkAh0ksghPXQyfKG
1fa3sNQHJDch7jZpjS8CT6sKjMwWRm4F498pI1hATllOJXEgVn1jlohnZS04FfkaPi6DYk3FI3ic
gHY5hX+p2R0G2RS4HoHRmv1encgg5kMmf7HbjJyaX57KMZ3IPgXg0eftFhhno7ANzpHHVaSWlEqX
oxd8JDcM/OkzjqcPSXaV+brzCYEwYhiYfwKFmYoT2txiLrra22zL2+ddsjeekr1vY6pAc9Nvbie4
QdqnkK5zk3ed4ofwwQ4kqIt9eg2o6E4UkkXa53SVXuT0p63IgDjOXxXhLpwCZ3Xp9gEPYcLrcvwy
gjU/E7mA7JQVjJMUmMyjRFTVKQeoESvXF7k/pxVhAGT6/koKHRiP1wNRUcw5EmxZ6AJYok5DDkKz
hlOU4y9JM9SqYqqQVyD2I85IZ9CGPtAfSrMuledNb76s918w6dtOjjPI9+USU65JTcHlIlTCo74M
ETY92TrRfWhUDHofxFY6U8OWkjUzbrG3tBipdu+YEM6M4s1O0pJ0Y9wRsZ/lZp/qHfI6avKwNJ6u
1TA34mN7TIesx94wvP64nIO6dkIumn7j485NnYGa8K80PdmpwajG7EUJBNkKYye6fFXD0Ve0kzan
jc8SMCHB9RbWEdtj32N8HI0T1FOU0UTPBpoIgHMhKfk0uvykU/lpEMiaU4cVKvmkx8nDSbUuRmpR
U45viPd2jB7nO78LaCspB/a0HLByYkrj4Vv+ztKMIq2xmaWMAr9Y9mtpCb7qib5JdHJcPWrxf2fh
3WWDSYyEMW4Eoj2BY+CENaDdILxK7SBkBBMf97/61B7+c0OWPslrjjDbziT1Du0ZaBcCe6qKhI+L
P2wFl5ezFo2I1Uoh3o26xE94yddToF3OdsPbYJwaTSGW9BVI7hSGSMuEbDyZqQgtJ7uSIBj3Ew+M
uS/q0+jtBUEVzgXoH6L+1zfmgc09gbbSQizYzphe6gmgcqtioT7WTn8MziM6YQHsZFoXrFhQugVq
8R47QF1ekea3ENsXY+GozyPvMGQYjOBVx2OEvIoGO9GOnyohnl1d1bPd2uOEtJokf3KMjUHEZmjH
2HlCnnpA8WisXPdHWySpg01SxhFKC+brT2NJ0OkcP1c3j7s9e3NLCU4Bb3G3M4iMPswc0uDW77Bd
uyBjTIqklFZvEtXGbfE3XybhxqTdbtU9c6xjNS+kDeS3Kew9jVdfBKodnLowG8svvg4XDZphECJe
9HOvMxv93girDos6ma0QtHXfs1LnIljVSUw9j5UdFxM82HtISWEMtPg6kFc2KSlRHjqlQ62Xnrqi
WUw6YQbsB4sC3/QmOXDbouXCbSid+UvQcekUueU1C+DJjplZLp6TxQEaUz9ZPBAOUzbW5rbpt4s0
bn3pDKqRQxnk7+uIrJbE2eZjod46FwGk1pDp3bzf9c347Vh4GyzniPnPFUC5opdF+5VYWEnvGaMK
PYYG8NIyLihC1pT6sMsRcV5+uN4Ut7pctsCid/U+J7GNWddOcWU0akrJrN3FGEOoPIlhsTppEDS9
kztawCQmublf8rQ/CP0q0attRutBKdEiFyyUK9NaFmwa5R3ENPH1CPpSRlH+En5bELwpgvtH7UML
/9Bw0R9uRcM1F5NgvPS3q6aUjbcTHz7L62epuvOiPWG+smeeXU5prz3oABexQKXYReNmIkh4L99h
os7WxX5/UsgcWRhXYY2XJqdNASSyQC/8rkgRhLjucHwB9zrGJx1k/OczRrrEImYL6K3TWxEf+oz7
CCSNu7IiFG3XiPChyzRX2s8s4M728Tw+BQt/RG22QNMj6TPHNkR+kuub47lJgQ4jeeadDwc39E6w
4AC93VCc1XmYr/Fob1ZvxnTmjeSzOMv1HQMoEsTcGte439c4OJYRSi/55YWoZ1x18ZsnvjZo3/Xw
qTgOfXs6U4KuMj4vcQrnasP9r342Tw3E86Qub+cjV4LGFI/TyUk81NLhijAwQ4z0CAiwO5SlFzvC
svhe3kSrCGCDRIgz+7bqSJZLLEOvrvweDWwDBNwyHHODLZFo3dBjSlCjTQr8XLSLStmAIVl9ZLn8
oVz5sYKBoeqceHF+5qsG2qPc+G68eITCEHy8RVphaj/3oef5zcSyCBhETQKqJlWBNWINMguQAMIM
V7bX3gbCZiaui0iHoC1FhMJXKt+1WAe0AHHheW2tzP+yg015T1/h2AE1dX9yWNBpYwnrJ+IplYK/
bf9QJ1/ha/FyrKuXzxk7epfAQ9PZmtncDKmZ0SwTXHNU8lv0f39iHa4pCFbVCxalsvtc1WuKGO6Z
vlTWS/WYy8W+Mf8c72pZKVQT1RYltGjhWKWjTim/+auOG6nx5I0mLhV3naF3p7nUv20iQKdma8Yk
G6e4rjsNSdgYFQs4tITkiyLQtslYrvhxyBIoIFQ8cktLbr5ZUTK8t6hJiFqOUrUQ5FdBZGhWyBGw
6ac9kbdKcnszj9bGOeZyEDVklJMv5G24yuUgv5A0DsWJ4TE4DRN31/68c0Ezfu7OmzMW3hg20t/v
wa3uR7O+zD4kPgGNQF/p16j1i4Bc9UG0ZTbQZ6rWb2rVp/+dCKXK5jJ74xcL4rfVdXLHAnXAFwHk
FiIxN8nE1tbI71YkA4OqdgItfhYszyZQD7ouUQDnQkyk+Tso+5MAuwVAuyHeBeogkbJMBmawJ3r5
NmX3R25eQM9nKKXzIdFeZxyn4KkVnJZ1KSB/907KhtrQWKDBAfIkod4ijFIC9n7GArmwc2bckIvV
yQswVrNxO5q/0jPLIHGsC3EVdrCelQtWhqWNd9kQ9ucIOMo5SgYZmvBN/QiasxC+otGjpjFux0Wt
C6DGFubhawVUSS4HiLsjhQ27tuXopCPHuroAOCqoNPRh1orPqMaPquFf5yvUyz78bUe6Y6XMtemQ
zKi0REia4W+NoG6CGKpIoTbgOG2+4jtovkmy0mMuE9jqbzOPr6JeIO+zKLNISAIeweRWQlfqak+p
NFBMNLAAA8ezFicuEiqrRwiP6a6d0d3ua7tSjG5wSAIt86G3qhBNQPiZCZgiUGX9gn38ao64Wyp/
LBK6Ixs9qo2ohauvWaFhL38f+xHcyzSfFhZaluFQ1975ylKtss7rGYAoiJu8eaC/WQUla8kaLN/g
oOEMqWvSEIgsWbmToKmIhY+i4UjyQYeGFyxPCKFfsehTK1zy2Gvvnx6nNkJoA4VfeLUbehpd0+bc
/QMYc9ToisRcu5qBBxCj/PFmFTqeyvw1Rj10izrXFweO2juqLKwHj0SJV/x+46D3dEEQ7eSGFedD
C6ka7mzOaG7QaHnL01AMCe2+tG0GmeOSkRFJJY2aEPtmlSJtPWVcvWsV/OC51UTAhK+OpgVZnLNU
7sZYbnJfUyirobuZ+Q+ibBg08A1YqU51Mf63CMqmAWeqwe8fgOFEuX7owwQO+/CQj96wxJrtBPL9
s6f65ECvl4hoB814uiD5BlZO1JE52L787Uzd6GZR7RmF9/aX18bsC9SwNUo6oRezpTOm/+4PPd0G
VeH1+Idc0+RUSdSusyaEB7pW9WFcmL2FQOTUHFik1bfqd+bgHoZQnJ/nocSBNRWNL9TCnQxTVUsH
tZqikiCBjumehM3+z83xwgcFWwfTL+2kC7lAQRm1HClm7NkkkhjItSCJvFQV6A/ZLKCaZ/QntNCs
s/tEpropMGe0OsbVcxQqWrpbaHUD8MmjO2GnqdOpbqjVmvyTSsnBxpwXXDulTvJO2PeshyDDr5pt
tW06ChIKYkse/YxVXBTua5cH5KGAkRNI25eEhnJba5+V2tF8ZSP8SmMnw+VGd7HLyMCxYX9o2LnC
janFdR0BqpWptRqcl6cPyGXH0HwI13hjscllA/LD6qfyD6wdqWXggc1+cOzjRr8LGPbcdd7hg2rM
+KFUg/ZW4h/C1hMvmCGNmJF+xjbZmLKFV0wPLnm6a+1Gv9YvukGF5irOwri+/lCnAX/mPYI6OYEx
POO13Z9pCCV5ULkHWSkhIclEt1UG3pI1V6Fu3LsFDHEj3+tV8mNucVMiiGkcTELVn0fXiiylUSiG
iGvMnYi2MXo0IpAbM7fgsBlXFTBWNexXa3wTAE57+dIMGrl61MewX2O8yb7nrswzDyKnsePsS6eo
AnNFgYDVpVd62sQ6/GOipH0A/D5FO8fEAMeE4xlRTyxryAfXkEBiPnNDM+vOmA8HicN4Ss3Kf/s0
XzOdYvpDU6xjOGfVafaQsA/POsrSxQDFqLiBLEpSmSnlXx23+2dnqDSkVTyTJwoEisNQOI9sKt3b
NdHGD2gB21ydofUuJj7CfFxn2TO7ibBG+aKvp50bEBls4ACskqKNUlKGbFyw04RKP2mQ3KF0hgaa
tyegx3dUq8ztRSHBdDaASAd8zgMeJditdDEQRJEwSPZRcYIFhTGE+EXzTGq7uMKqp4oGEh1nLC+N
syOcGt+Snx6aGzDhNdrBHrE321LXPG5o/hS0Vf2w2KxspvHS9jUloL4+PvsZ92OI3hB1soMRYtC/
hoCE6pTbXrKwdeZZ6xHbYR1MGZdXusfPR3c14+FmMXfG0fe5dLSdpSHtssYf7iheQFwWcQzBN6pR
fnIp4plwZkqFbUhrRB93tDT6HcZDYEM864+SeqLrdE55u3t7AQ/WgLocq903J09DieHRC06GGNn8
wG4Sx/diX4QjxTQOX9r4YMlrl8Szg3RrMJ0kq8b5hzAdn/Ge+KGNS1mb+oDhaR+JVa117Ik3uFAg
XjmN+BGSv2elN7pNXzDqcUu9GGZcGopAdYNMZLy6UCmWA2hpRbOwfj3gNDnxOczLPUaMcnRe0PtJ
rcGBJckq+LXUHTVBDY7pjhuxTgdpeaJv6ldYGpJI/lHXmjIcndEmXyY/8idPMlQeNJnAPydVKAZz
z3v/jBmenSJMcXOVtJvC9BT76K6XSJtFww+4EAzTOsB9ilqyTv1f+dG1gdu3CkWcd2TxdZKkFL/n
DOCXY2RTH0PD0GDfQzT5hVRxKWxgi+g5eXdTzD76UcN2/ZcEmVbr5NP7Xbg3c8lI9BnV8bVVJAfd
yH5F7NNvqj19vOiPPMUYU03FgvgADiBe6gc/PeCRoTwsrtnqxT/6JIBbW2xeQe9Vu3JBs0fXT/y0
B05jacz2Ss0N4RBjPJZVpWMt9Jme/6ZpV3QV3u4C+3vE4JvYjjS23e8equjiDdhwXInNNe+kJlnV
8uSC6974wKln1hUsMuqs9y2Y1Chr/gtkw+kiud/wBzhj9HuWoC2hKPqJhP6vokEIh4T9LO5XlUIa
flWWFLKBUrShsyIKWPLjm6zZq6El/RU67+4H+KRgVFP85Xh1NFURIl4I+lgld6Atc3xGukLO2Afl
VZ+05xSiLttgeAghvXmHlOFBg5Ar/9sXjGi4X+FnTPEYddGKq/BU1tMyjyk/JzXqhgT98vnqqhJQ
oGQXvmkKLnUL6lnj1L9CalVZi5zwqMT3F6Sje0beTbw/xtgS52nGeUw0dy5B72tGG66ngNhsbdZH
3w6R03/Ca80g3qh4XrLK4a9AOS4hLJc2xNyzxr4WthknTCGWkMkHESwxIQkMAiaCW8h/bQOIeNOl
pNCwa0BtOCtCCCc3l+KLrI4lwkcwdr/1p1fX5SxX3nOKB4NN3bjEMdT9wyLelJaJ6bqyFneBO4uA
hZxh2/RGq7S93KFYLUn0oNU+ERMrU/gYqUlMsF+b4its5OKxvmvB1chQwPNEE4RVWelUMd9AyCvf
DD60iqpJhlU3zfLuENIMdPL6aYkRS5eDoPitQ9MMg+4lnVTWKH+a5f1yu2l8UBaGy7nQRem0lBx3
yu8tjiw+pvOtEFQLqt785aX/fGuMtqIgZSRzaP7/n2U7VFA4ssVk8q5hEoKSvGP86JsP1VmZo1M2
Q5diQtyVbX90jB3B34dn0btAZyuHYghOoCpYZ8jNxH4s5F0OqfuQeWaB9VFdBo4Hh1J+swxic2gS
LB5D4iRUxfFMjj3Go1SnSZPrJIVs3sRd72LSNh9XgP5IhJcUqu3/HsT3hBgLkCSN/1zs6zx3p/XS
KSm0NnKPKbUSjevmZ7yihr/eceyi3JH2Lat/hqbogbTswyghTewtcg/qdF3pJn7+SCtHAd4HLKKs
zD2hlTQJeyUWGV2u1+xOqEUT/bYKXDHNDz/K4CgjFwMqJMMsi4VcOK5nAqA6Jmqjs6zgCkC0RAcY
NeEnYEQu9Nto/DQWTrP12q0DimJeT5VVmI3TvkdWM6VvkrV8K76D5LEbapVu5z7VLVSPR7EacSJC
Lgc9eP1yRpqnv24oh+o57U9QhHT8+QcYhHEjJhC9ixqQCeGi1rc6lxhKmloHabvgAzOIVb91rLoC
KbeRRR1CEkbil2LUQMxFktYUWota8rKyNc5+ulOLqBuqJey5/OupEC+6sKiLVvUh4KaHPPWbZgDH
ZIe7AYh2Zj6djgpL0M8aBu7tX2M+47lD2O8468BodvFSAquRGFLcJ1U+u32n6I+WvZIAiclDPyJh
uPCWKV3C5TQh4HTHIUkORPILbvxWR0byXkqDDXYhksiANF/L0Ek7PU+OXHD6cjYqGhRr5vV1paY8
TomRAHa22vMyie9qTctOM7JZKKgkuT3A4dM6Y7e3/zrH/LDdaPfZMZ+ZzNFpfwVAAbKenD0aserN
YB6SH2WNaOfOVlO83oG1uE83Rw1ntHcyf4QXdztuznSgjFIdTHtG+bP80d02wa8iUocjuKFuUZtT
zEg1n/KyhBL9bj6FBzkvI+Vn0qvjdQK7rDRtQTJBc0PLHd50/WJE2IaXDoNKwgq8NfD6L5r7BkJx
LuXkU6Vl1ewFHY2rktJvsDsqeVyMWqdeK5E3nfCOC5nhiJgOiQhY1Q08A0QVDNS1vciQDGVwuFQX
ub3sxfnO4q6SSL2fp45QBmY+9QA/ZKpW9z0EXV/MC4aAP9b/1K4dj2Sk9AMSzwk9r6nGhceiKCy4
QC7KhD20iQFhZ3WGMLWQH+UnLqIJhROB70MGDR4QMEkMAN9C7HIIYTgOkR4wvPDoUHPXv9l2OvrM
vuxCsWEAVtIQnlEfRl9TxTQdwcSNu443RUS/YsAuWJpXnpUDS1N1nhj2Qw6Dnz6lNumyrQRBsqzv
AZPA3wFImpzl3P46BBMDlWg7FyOSh+VXROor43BduURtxm/nErUjbdTM5fkFWkqQqdeePEHe+qtq
cAp6ZbWqyiBsT8RphqhaHphMqdMLXp8B0W3/cwGRncGRuYNdP2oAegtj7Aj/o4xkSrxcuCjmg2pz
7/9i5PQIvofFG1xihdg2d9vp57nXwm8tjQ2p0a20TN4UVoZIXO3izZpfkViXpFhYDpRufJF5nzX6
JS5u6hwTdFEbgAFmjjsqqsgVmwsN9/kK8gzPd6xey9Nqf0HVL4bCDS7WLIyeiQKPFvxVjJPb7QeY
3jn/vHBgSZ0B33L9EdhcpUf67S1KR8RY/vLiTvSBvUAKa8b3DGt3RrTO44Z0Gj2rtD3zzV8zQUUf
5qApFa9IdE8M6p6bxqT5kNjlvkc1cdRrAYN89xAGMmN3hGbzhAvvxPzuz2ezEe2+qSyNfTqyghIZ
AvD1IDUdqkWq15bF37KYb5yAguixGHUv3NyCjgy+vIvkXqOXenQCh+Dsb/NlRg4NhbYnl4q1mwP2
W6CZ4jP5DzIegtlsLTGpbooADQp5UzIKjHjo9AY5GJZgDpEsJ8JeutjV8LBD2AWvwEhbmWiRL0V8
o2Dhtv8ZAh152lGbCjidVT+Ky7Yw/CKOb4XvUsONDUx/kWzCzssVFB30O2lbAzHhRg0PXILciMU1
t5OfmumEONznes+XsCHGDSCOqgCUED/Vz/Uqq+UmQU6JJhNvzl/LvZAksKp3VnMoTJ/NnfOIfA2k
QX8ZPeOdHiP8gSiqnTIBWJQD29ZU3CzIgoHgyhE+ObsYnbAFVTFZ0eLUs82UwxGN7O4OqvAufMI9
O4Zig+cGbpheYnl7lLuoj9I06LHDoWCLEotPdyma6bap7xV9zj8NUNopK7ahqW/A5BIAXdfvM7Vm
1nNAZ+jQf/xGr1ZpZk9zHJEMEfGBatp7YoWy/FoKfa0HXpBRKdQ9PSGryDJyr610HzMlYWbkalKF
P8jMNpLTD1jvqljIrE3WVY6t4sRYC1FwDbMFYg/6VFt5x4ZlZ8gp1Hsy3gC+J3+Uve+ec1V2srxV
OWOBkASUeUSqHB0aJbwToXZ/xvfnNVgybJRILpwLuZtIcMAdrGabhHd/mQ4JxxoYCg7bzuUeHG2f
t9k3X7VQ0kZ0mDHrYNNVdac28u7o+zCbXUbYn9CGoxWQXMjdOig6jI+Y3mkm6zK3bYyTHB+OGX50
lAuVxnRHKxafNnTi5L5LY8nutl8ho2qJDHxHkMT1vxY6h2dOhtaocKQKSzekFBqdKgmZ5qoeLAse
n1VeshzfXS2yUwPLAJTUXYgn1azlntRdk7HATXW33lUIkJLnVsxIYf216FUb0wYXXmYAklJWozqP
qcwcDvNH2NkoszydbD7g6TewU9LO1WPNXDY6UB/Q0J1on9CuOmaMMUzNVgbA7I2o6wlORiVuXGTv
9uYot1/htwoizJALlGwxOigQtaxQbmEIbgAC1YxUF5xwy/okddxuoIh+EykSDfyhwYBjtwEx9dKJ
5qG2nkJAq6wN/C+C6xhm6xPn/7vWF3pOBRN7fmoMI4JDGXzIFWQ0+9xTLR27Clrrh8Wyg+aUCOc6
aMtih5eBtq6HbVYXwU3rIWLZqqkhNwhe4arOCbjgMDZO5SZMN5sPbRMWVyYIAEemO9HsaNmMdM/H
fHICX7bVU9jLmEls0Vo6EnVAGCs8kNeciqtoUHLpNMflrgq2cYqdDPECmt/1XFDzpQIEIFLaYxM0
AnmJwudq+jn7N7miGe8KwXgBmasg3S6odiN/frKHx7Fv43Ki2jWdvgSmT25POI1axnDJWLa4Ith7
A8Cz1AwFHL5iDwrZkYicb2vXLkmiyuoOGSW8bC5Tdw0jNG31z1v+r4OCuVoZebsqtZjqDgp67E7J
he8+27HDR+EPPc9S8TX4gdbUT7bRlJxeA7kdAmXjGXtC/1gCPV/LJJF2KOo1GixWgRhvo8JBahSH
TMOP0PDV9rTyiJxGheQjfJ7Deuni8EUMgTVQAUjGOA3RN0DEL2P0WUJfmPLHDkCvL02Aazhbp0Ek
/S7tCcUsjXyS4pX7Mt4nYyRJMVSy26GoYV+kK0S7tu1B0Cd6v7dhOQ5MrJWeJq3LMjHNb4og58Sf
gJ+NlEcPbJbyWEzQfzQOEKonC6Gxnz7OFOEKOFJLYQv5D+IJfYChHQWFko/fY1rq8mZSRymFoYr9
dvIukX5B4oS8Y5cCPC1xrwkNdX9MsdjHuB9ojiHhFTZCjmB5VU/9HSnrh/rX0Ld7iusAwrtqTenp
tlDQ7ev31rOWpLhnzQ4dYLts5wjRPUYviSqpXoDXzhqHH7XKojMWhAlLwyrmNlr+3rnMYkTpCdjE
SgLFePDXNJUYq+sfaoAo2iASbze+haEff/3cQQT3hc8SsW6dE/W3JocxHRw7ccDaL8cYdpI59Y/N
62fy6O/fDsSehCshg4qIh2uzHh4j9HLW9HuQoydjnVcgZxPWYiUAOTWvsV2jHhwi6PW6NF8A320B
rBL40YtDKcaLzCR7OdRBeQ8E4eB5GHsayVxsZgHrUWHMzlxKsh1Bfh29C2ONaCHgtPCplZO86Fb0
mbUaVCz3KEw8scn12KZc7ukBlMQYHWLjjzH6Ja89TusVjFbm0/SLSYnBix4bifXvnvFVDRgMP+KA
kLl+mVRdcH8YVZvRFykFIixvFaAaFN91uu3OHpA3NWwW9uE77vNXrNVYONWVqh6ei39gndIhvgPE
MO+9dhesopik/cOlYJ1L0S3XSWV06LWbIxy5b2mxl/vIxqqHNCRHlq9UE3y6+zuCmWPklXd6zlIZ
Ihhu86D7dlABz6rOvEwAHZMjz/J3qhfW3tdpd602T5FZpftYaZMtdXTDdJCsadRtp4o7mD+CdU1O
8GqDJQ2VfCuW6alYC/7gOSsVKg0x4PHXdWK/vU8k4GP32uDlBoZc3wxgRVVcPxLrSl6fOG63IBr+
f1u4x6i46oOQGsbNSqIXHiCGp+Eg8ypCyXa4pML1eRdIjCoH4sxLahhLBdu5o25l/eIt3dIP9mrU
hkIadOrCkbH8NC0hJZx0ib6osHzVOhIvskT20Z2Ca/tWsnxRLkNDvhMMM22Lx4IWc1wfVQkTvF9w
ZkvRSZ3d6v2foZnw/5/x0WLbFpJpKUDbD+FgciCKEPkWta3UeSaFQgIe7qz2YiLl+JUr0rSJsz1g
Y40j0eiZjZKX98AgN+ag2Mw42tkMW2WbeDZZnvp5H9zcY2rYvc6Y+0fR8jmxwJTve/u6TYnx/dEb
ajzSu35bNMGXS2aaGuruv+KdPWhp6I+m/A/eM0mL4dpy5qXvt9NDFpvt1VYUuCMpU1IgH8xrgJ0i
1GIRq92eUfDF8Zt8VWRQ7NGMzCsLwxtBNfV/e7iB3leASaj/RptyCj5pxbhbU77wX+pSMTVV6CDT
wbkQ/YfFnMZ9DkMVqfwbPOpB59zl1hgm8AWxLMRHHFR/LD5JIVSl7mA4Ho5I/A1lFaT9ltw3LXOB
02YW1D1fisCNiJNc3UMqAaJoJIANjd6PmZMtedeXLsZapV2b+jY8GaFEHjC+6g/TPSv7l4XoYsdj
N0b9Q7FhO3qN71ovXxBNUYabEN33xLpyGddJX1aWh8uJhqIn4zu3ww5U2s707OfzO/ST7Eboja7C
BKbY4AZcKF5c0raGtQ9EJKtEZjZVNKRgN1CyhbaEyWG1GE6U9N7/BuuSgAkk/R8Ofhcl9X8XCC3e
4iYLbh0kco/mSbdFOqPpDwyPpJhK13YmShj3S7ZKJBOdFXvArHjIJC6cNisRqS/DNupBIgLN/MUY
dSpkkhCEbqQ/guzHolhrD2XZZMDTvuFs3yCfb5C1doP79JaR+j6JwjxA6OJxFIczi9DGIskfZFXY
OiimtNMZH8VnexNwjOhNS7Y2QTxPEuOFLShONat6GzRbOFBBccwdebj/z7XMAtLQIvY3K8jYGwwU
9i0CDSr6+hf2kzNk1XjmsuulJDscTHLZ5YgN7q0R9lh3i/VprJDIEaNzR7Sd8MXodrHamxDHIIPB
tA/x9eZQ4uD86gWSFfBCw02sLGHK9ffBUPO1td1FVO9ApiRSeqcM8gj9OVWQlJT9IwrPybFwl7mS
YAfug1Ip2WcQoKV+OdtxoRAS9pbAS/unAlmX2o3elo6fRUb3DXPEjZ4/vXfvqllptdToE/3RHfzl
wdckUOdqxCdleYY64n7unIcil0I8owiz+ceVEwefgLL1TT2iChwGTq1lUPtRPtz4WicWwcUuASoj
STp67Mqm1Bv6EwhP15CmPC7Locdn/Ks1r2uo4L1SrGZwL3VEWQZPz77gUEl/bJgkWxxhpL8n0oKR
taE/8KLVCM7EFQCIVFynFzkKUZtsHM7xWfOhbm1+HVtnodHHe9WzKsH8mdiJXh7ilLKTl8qL7XVo
BoxeDxnJSSqwwbSuFiMwgyZ68IyrEU9o1IPn2paSnnc12YfYm+D3OYb8OfJFQbjSMprbGZR2Y2Rv
aSfT76VWWz/nfLjKmSSneSe0bZFcIBOTcQh3rPVwP5NvYp82OLiJjoqAV8yIXwg8E2fgXgCOwceI
dcpcYUivyeGcgoTz9IZLPtfXR5PMTIr0ULI0wsE9vfIBG37sSaC7VLzp70aUtnSC9YuKkquzsxxK
Va+8z68pAJQXK/4baVpwQS0tC3x2Z2wJJxiU6B6TNdpH7FB3cWSJVcHnlNFY4U9Zh7kUQqSx9rtl
fuq9lOoR4jYc4qScHc1yHXHKXYCa/9KcvyakHMRDNrsGgYdCuGJAYHDFHi5ZwV8FEyVQFZpICqld
Ss9LJKgibsQ5t2m3q7x/S0i2WLmflhd90113tBRjglSDHp6Qblj/Oaa9LgC2PFaDV6uYeQ8w3O2j
/s+YgDMD4NR90UDpBxSD//tw6Rq1a5SGghJpW0XYfHXQx9XzK7dynpEeXxkPevPjGQGCb+qDMTo5
7zg218FBKlgq/eV6DPM6AUMD2BpHe3EQrpw8LKfFZgX54rh617fP/ZhFV9LDedDOu/nVG458H/qB
gS3xmTjJxpv4ezccuJnLe01OuDQUybU0LlDdUXpMZys+JREhxcu5oTArAVG654qAxro7mxqf1Qqa
BgBCZJBVTUgu4XZdRUT8EAAPxJIpLrQZoqLjz/rPL+H81O+ztWwOnUOELed4YsGotHfo3Fi5Ya5z
BPYfpN34zrB5BL8/S/vBmf2HsnmKZzyXSmuBlRujq4nC4z5XYTN2Z9N6r5QSvMSseZaekYF3zdTP
6rSxPeQaznMBTfnFE+/Yj6iiEMT4CNmytdofCm5vVt3F4Wz00a7xqnv9tuUuTyufVuHBB28ma9i5
lx9U82E2KgZZvBRKd5Zz7L8BBJoRn72wDmoZMfy1O69uq45YjuqgGZxDu4VrFb6Fpl5LJb++tDkK
wd3YMJ/nfowmRdOl5HTq3wBfU1Wf2KpMZrwPKK6Gl+NCbIRyRmlmd/4JyMVtXZ+pNP5AqgNVR5pz
IsEpd7aD5IruoWb8CTHpi1LXj+Hsasab5I6SYM1/2UR/NoS8/SmDNGXLafUH6VQqIQZHwUEeaKBf
qqqS7WC0i2U10EF1rra2GtsWUw0xKCJ21Tc7zOOnT33ZiHiAduc8I7ZP0WoRuXnQG+8/+jnUnzFI
llT0k23ZE1CnGj69nOoZNI/kjvTGdqTpzN24Y5ORNT92GZ1jEMqRRheug2yfrTuh4fnTieNMEeIj
Dc6iHon5BjT2qQB7a1QVZfJceDblX7RAmDLiAMSHfUKEKC44d3sovjKZu5wQ09pc4NZGQkTqa89E
RrMvHS1dOzaqxtuLhtM1B3iOsJWTSz9Um1COZw61fgmxb0FWvDCasgqFwzQh/K6eNzDik/TikXE7
OzqYbhNrdlaEIDHMTIbbFeLtahMTVA6nE7KYQXDr5HzdLJP39Pef0zDK8GGdnqwo65FmhPspULap
vuwlT2uz+9k/jKSpKI9VLzkh8S38usT0MYhye9nZNqGWNW/yRPNs9JXkg9UMk6vE8qUxXSIJuhmu
B+lsdvigQwrvbR7POg3uyeBpVGFG+oNy72FVxnKe6gjwSxfjazujxEvUv01HyeUzcBxK1+2W500c
7iFhRk0iKDaFqZBRi6Nn27zPwXbDR9s7sgAMehFtJvTuwQNzPwf/dHzAdHxIUcf8LSHXzknYraYs
GUPCD7YcsBC42sK1MvMDi6ZDY9HOFBLHq4xldXMO/nM1c/LnStq/Y3yQzdoM1BmKuFN1rJzpcyWh
jfrpQSm7faI3IWxDY6GMO8PKIX5ho/U6gD8MXzLhYbxMn20tcI7kOUJ+F/8HCVqbtRsWRvIxkeI2
HaLW1jMtZBikAEL8FvJY/Nv1e99CwqGloK7paRPfUppya+K+nced7MbIW+b4/dvmBTOB0GH0IPvX
vS7ynWa0rDfq8+TKCTFtsGHC5VCNGLUASqB81Zez3wYakBwgBa5ynfOjVTFzvRtbIYcgpC3vrJP6
H7AS20qyCEydKFVGesiZBlj3SerjJo8NKe6EPHC5Jaq4Xou/Fe2u69eNMSrK9HOhp5QP5nMU5dWr
mY6RiQRB0YUXpDJlvA04yG7aJgSZxBb9fchrWrE2n6SIkbzw/ZbNHWuUEsXdYFpfWfy4UhcfbhFR
jHIF5xMXlll/KwvdXKvmOrhiEf+nArRIIBdmvPBRo2ENpG/x2MrjoQp7DQMfV3bgvjcFpQVK5XoO
DzK75RJUWV2IhmXlzN7zfAMnAeM4GmuOf1c+byszxmYQ783EkX8DxHwYn7tTUsBKuW/w8NufRfEI
lIQZPpgEc3I4+fEGINA7IEPuZAPvmg0Zr9uLi1hPzvsyB/LS+MVLfRcoBKcZF5UsG5vV6hVrW9tW
0uiOf4XlHshbmFeYlczwa6heL8dJfVCA8MZSQ0TyQsrrvPHrjX2sJzJD+k8pAWn3mQ0mHatNm0uD
VmoJY7Rm6QmW8J6UuM3cYc2yNn2QTXJzRf1YZWqvU3yMzPUpUPAPXFL/CNNquWs2MMIBOxdUnpnr
IfpEjyI1leTCwWsQ3rQF+ds4cxNle3qD0Z/x9ZdCLDHA6wTz7tH6F74B8yXQ2kkTjlQwJ3Qbu7fE
fXawgUVMpB6a82/W02xrHGngFjwrJkknDkxI3E93sdqHRaRjgmzvWPVAmAL+34O48ggo+AQrEWQY
zJIMKFnKd+8n/C444MXI9twZNl5Pv50KcSJG2SBOkLdqua3bJxbY1PlRSCILlrRO3bPlhNQy5hg+
CFssksC/LrawA9tAljDj92N9tSt++GQ/zlb2oCSFJ5vDs7SGDPNpFyC9trUb+oG6FELexZ/FvPND
lxfh1Zt4+BvJcQhaJTvASmR+teXndPR23IbJ5TqpkBTdUm0+Gm410Cwf2xFKSO0DpDwD7X0xdKdq
DAaFbezxp98+AtTwIe6xh6CkPzm1udpUJLvM7uAM0+DkoY85PsBeCwmuiWw1PVolitgZ2QkcpWva
E81XvPnX/sGjygvNK81GUeRdDsgg16ckGof0ME3vsMaCBCJyvD8qUPY2xto/Ow/unbDhNxU4al9/
3qeaqSIolsWs8TQ7PvOBa0FIcFO2kSaMwlk1vHOKBTXw6qOR1F/s9B59PUKEVYG4MUc6QxKAw9EQ
QIiC/KvCGGtqQ1feAhvEqi6y5hW2Y2FGaFk8LWHhKTIo4zZ5G8agMTNcT3Sw1Wi+h1cwo3TrM1gJ
XYMbv5eadHCvgTpstR3qkUhTJYalYEctKv/dz7gprE1PuVCEvAV3HL8xIZ9tEPQK7iEIPkvdxsw4
g/e++5Te3Trca1B3wrI2HNj7y3QVEBjqojocdwcPkIyyZJsgsjfs/U/7vSrN4qOTlSqdCSNE3n7K
lFYGHFnVBx9B3aKFtu9ymSmC7sYS+ERvOjhrd0slJnxvqKA0X1L0BTao3Zl+BB4mz6+ahJhSP0rd
RuZe4NctAeBENKArPp+ZGrjMlhUK8MWoBUhpiO0NRkE5MbfSngU1MXpDDKe9n7+BtASc6VEbtrFY
eJqBTF4uNdamvrCkxMtzke8MtiiDBmJk1kPhoL2w26BgwKcomroSqOAT4MYWwJVWquytxZmur8SW
1ZY15DGc0GRe3rtxRZcCS/5350+NcdBVR7uY9xhy+9mNntSc8OdJGW0kLowBxSi5KecX2ei+ANLM
L+z6p0xdM6rnm5Flt+BDL7cRptN3BDbX5mBuj2uuz7sFfXp7OfleanT+OkwbylyM/kPimRjlnjr0
Re9E98VHxRVi9MyJ9mEmt4Ddo8J3Rp04DOd/04RldtEXjHryS1bdjeuoayrcHYOT1hHS1cjrT26U
268Hd4OYDA+CvNyD1Fwg7uu2rFP/jb5DowSkc1uLT2VAy5vGrcdIqdZgrS26qmIHlBRHMeknn+go
kDnTbriSnariSkOUQR8VD7UeUbLPC1T/JUtmLIUedvTPVz7rpVTOwShpW1l+TUZ1OnyqCbYfKvwu
loKa/lta14Bso/XUN2OryvTASPLiKEaxCBn/QeS+QdbEKW+duh7mjHuFm7v+CbammO0RVfH8N2CK
cLXOt+AACb4olK4Xn+h1cKZfOtmc0FqFXgLSOQYKLQbolJ+f4YsfuwQRUEAnRBJgQWm2jg/cnN2G
epnc/VJW0/WXJYk8TjrftdJamx3U8ZgwOkT9sjlHQGVNQzzlkPMaQwZyi79Fmqxcuuikj1AY4Yl3
aEkKBr9bWaszVJVJjclKuL0bfsVzzyrf0sHrjq2qDzxb4f3phEqyDlbfPvOXJxCFciBcoQEcqlHc
Gu6LSkePcZy2Os9Hv8LirIULwvHIC2WAlhL3m79e8EUjkbhEZWJ9yDq6GMDkzhUNigJSuhCLFIT7
I3cQciY0tfn2qJzanZ1XMU10xWx7i6rQ2D6/NWiDczmdvi7hWrZfEhongKYBlflRb6hMr+ykjZzE
NfNDGpVY15dyzYGoj0+5n6tXAMbLJQWV4RzZzWRLcBJZ3jG7sBJgT8ZAjeMNy2PZDJraetefABxH
nz6OOjmFcepXAkGbAlwz9eZ/1thupFK48ArbfznW5USrBRlZaPIr8df8WICQsqMaf40DSadkOUNr
xS5X5Pawa2k8xuMfI9Kcxmijblwx9xTUuqladPhVbbxWAeprDLxXpDVEVZrWygCsdsrmLF/FPhGi
OfiCcpCWq6WFS6m0be5rOCScWpdNaoL34o269NT5qx6BssUt5GY1fiehg6iKgC61XEUuNTgdI38H
QEqYU/Vzvx6U4MNzcQQlsPOAonocmBFQmJpMlK1K3lWdZ5RxNUrLVCS5kW1TRmnXXp6v9DU1k98Q
gAVS9iqN3BwGEfdBZT8g4C1CtokQ9iv0LT7iCtzq2PW3Ttf1uxLTQYyrXQ1brdIgluHilLsDrtIL
cYDw1qBaGBwgXLSDQkcKAQgqLJWcAJzSWeFpUx5aya1H8XNw3TPAJNr7VZ+0lOD/Y6U01i7OdP9g
TbyCEpAGJKbGpwqgMJkNBGCNuDqln6h49pJ07SOmRteCemcCb48qrUkP47uKLAxyn0LAzKQ/311c
nQTEJIAwoN4lL3ttSLbs2dlAbQin6gAbZhK13jMk6adApNrgTOpoRLewskG+wIYQpSdlTyTJZvOt
Vwk4xxwGNkSARpcXIIRWYKeRLh9XYSwNNpndECTZIB1dGE08mXrBXsfFite1Y5O1yvpQC/9sShuN
GDtN/RZ4s+/CbQsiMdOxYv2W+8sGk/0jdc7TUa1udeYyMxz1aD4+6rfgadHv/RItE2Q4D3sAlGpe
YPBacwnKte6bikLpXa4OhEbfJjIVW1Vbgx/XrYWg6HjBCE7ZtOOK7VNbqQ9x67+jx6P1/3GPR87W
ZY7zOb6bXGoBd9qfZzdmFvbK1xecgU0cII8NlEX7hjVNj4Qeb2dCUyD0RktxKV/AzXhK2XkedyDE
aW1J5UEFRecZLFpzYZbQ+cDGSwctbWIisxh0Vvv2XB8Ft3K+zO9SLCZRkXKtDJZWL/udGygPuzNH
wESady7g35+gg5qeJRSLh+dvs0MXjHfsSTlugWJzWRqi2J68BCHcYtySV4ncT7oaFLMFqotKEhxx
U9noe0WOTgGJRh1jz9ze6iokfQKMu4u4B+QCyfet5M8ulfZtfdtMjJDywcPTQ+HsRcPGXoLkAh01
hQl1JwpnQbRlwic6NfBG22c8v+d56rlanb78N3slXksgLUr+9AUYhPjiqSxlQ1XAdzaJ45iYrM1J
rDqIYywqWbU9oEiHKNmPHak73qj0nlNxNTFPowVU6Smp62UXR7kZWRmjIWmqPZ+VJiDoZNTnUMVN
e1h4gSosNSctygJHIEpczOqzrJgxk10eMANictYZaKNUJnaqijup7CD5+SCClCv01ju3UEPNkKX3
bQ+UEsTAvsvBI1W73GbI1Y4eXe1hOLmrPsXnJ0IcSTMKSj7n06uGV0gOhd/7drI3f31MK63x6UOz
UIO48SjFNUmKVAj21nZEPSVy7CNRu8dBO6rvBjLX7AUefBB1hFUPWbRqQEtD/8ujffWEHpJdAytZ
c3V/axOQIfSblelJa7/UnW0U6tgPVk9t/Bx9PK+UFWTGInnrWMns3fwfAx5uFUE/QjKPwdR+nYOT
2yhGFRyUjIFp43Prgj+WYWczYybpvQEzraW53HUhJNh9m0A9W/ZsrydRpzvjpO4P8T9fMh9zRUnJ
rtsAEqqk62LpYANlu6XxjwBo5zvLIto/HhzYtA8pLyfv5f6X3hLq8TLftM1hGiD2Nx9eUxwiyzmX
ECskaC4BnwAay/91ffaIsoqiJ6cGSeI+Y5P1ytrhjv3je7hXF8pqqVIK7CF5PTl58EXe5VdAsVhX
g4Lc4Sdx9xsbW5aPW2oA5t0i/d668SaSuH6cnEUoEW7lDGTlSaqh0akMd0xCqgbcx7EUJG+5bpQS
DGerKq7wPvWdwFGcAFtvIPdzw7E1g3TinAAGiBt25QodjcpULZViX27qcfWmrHYWjCLZ7YVWwa9O
w5jK1vXspP4TZerqXX5PI7YEyVlfTV67X7CBx/AnQM8ZIbyOKCLCuudsrlQCYzf9FMflOvCjaxnn
Tc4TEGWJNZd4s6jlGAtN54X+hKISjwFSJx4FBRdJUwpiIjIWEZPITempWG4YLjCH9P/XALDjMcif
XO8k/mPIb2PrXnRXpafo3SVrKx9BI/ED8fLs5QihM65aof/3t14GQ7zub3KgEdoCsOxMTLjxXN4m
SnIVq/FTTSj1nCMjUXQhw0fsBN8cBnrb8haygfhPSnblFyTd7AYouHBpr/i+RQZDUs6Emq3G71xx
uXeUnUccm3+8mBp0gzWf1xr1Ikgo4n2keJxkopuKtKmx6gYTGtkkfhtR5JlnzDnUjZznJzfBRFsn
JNNF0vaAaoQ8YrcOBj6iTi6WHdPKsqF137/mKDtvTZbAXH6t4LU41iXH/5AjwDXdxQBIkyupyX24
gzRUNuu9DQSXegfP46w9v9lLAKVUWYploi7srbdW1Az0PoiuS9sEaqyKgYJewizMFbCGnFWUu4RE
Enux5RMrBH1bxKqfymz5h5LV207s83Ictnm9hsaketC5HeKG3CV7cetKQfGHcxBakO46cMWF7k2f
ENyatA8+Sr5r3GQDEC7HbzG6ndo3bSnB6abl8Kdrp3eUYUdEbR83F8s8UtPvjONbojPvnHj37msL
eFu/m3CwgNjcF9wu7Q7czRPXJkww7kS1HW4nw5nNpcjR4V1G5ehl4c3nNW8PNrJ+S5zfwANae6Bo
66X0Tfe/i7xVXkSRlMJ9HRsqgBQv4cQaS2vjOThK8Y2YtsyVMt6UV71G2xyMMeNDflE0CWDl35iH
4Px9l2j6r9+uSLYlnY98y7whNxuRV189WkUKg++xWnjvMjR5JdFxuUBuIG2AjZ5hivqBuG5fg/wO
6+8fr1xA3hUE6saVefVB12JXoEyH325vOCTnlRRvTqTUo2l8ENIA+tZ8i9o5tclYiBFhNJjug3zT
4iqwWQZByDjaaptSpOUmPUupm2RnTCOHAYk4iQGRFEPDSZ3yoebXXK1znwjhYZAGuLKcVosoADMc
1L9R5J6fzzFoxdEpOf1WOpirkTypiWYsLZE6fkP6haOsoHqvo663wIeLuksvkkjZJdewxLJduvbn
1Z/JoYqYhz1B20lSmQvMAhVjgGCy49+ifixnBnEgvr/QHHZXz1I+DQ4FZniT/NgInNZNPnt8hpeX
4KYA/Og3lt+qYURSnD46oikEJmRcuDp347qEz/ZeYaYTBFEuQ/QdLS5WWs4UgMAJPj/A3bPC8IWQ
xv8fiAE+ICFu+QzWQQQqHHvtmPCqyZG/svUI5WNqd9Or8rGuoTyZqoMVJTrpO22jvNapD38LrJLm
MHoHH63XaUxN4Bkr8OPH7/eEMzPB9NhcWQKR5YIxJmCmMZSfwE3SQ4/gcIpEFNj9WIDUP0wSSLI8
7I71JI21vwfUpde1qcWo7C6DE4Ist+8StOg7KhTiGhpJddSXcq/CM9WH7nwgneYDnEWR9juBJdjy
/rdgLwlCQdtmfPQ/w9XFappYxgEBZ8UsQMCNLoDQ+9E7W2O6vwWqOMgYX0k8ac/NPCgddyWl+sU8
UJfWlpRT6Vwn9Gmhf0HxqWjYBnq8OnW/GvDCJ9NiwPZSr7hLT07tt9EEnnMdwkenTp/WtQg3M9mq
8D1scE4jiIPGc3YM+OW87J5aQ9AaPW8+fM1kUv3ywNx9Fc6KtZpwVH1dwGntSSmkwP56EpAUqiGN
jmTRKDl4VmvH32rN8Vd2seDguSSHZcORS5VqLKW9A5v49WFc94JHg5L5JKBIYabQPURrbV0++SES
8TWRxgO/8hP/YExHMlQugOJlFbfTBXMkuTDw+5fHbev/GREUAhX17S2iIZsJdsjVH5RumBA+NhXu
xHBhHjatirsF5O4i9n1g1RaFljKrpd9XLR8sU7wPFDEBKT3SQyBMgJ9zG89NR/49mRgVks2Q2gTE
bE2oyni+1LwxQBBnn4eNqRFwBp6EimRjORNy8csrTxaec0ZGVWtaoZABdczmeHXEYDoau1XlE/Cg
lqbRlWgzMrOdzGF7zBkkxmovlSzokAmDExs0zTedk7yq13C03UPFqMk5kT9ih6yBmIKUvvZTMdyd
c97uX5bNuuTXFGEcNGasuRYWr1q/GzhF/Ce9J0uCmlLDhVq2ZK+qox+Pp4R4+J0eWVIpQVl4qFEC
UVDtZ6kzCAT7OUF01Q3p+NL3/fUyGpBZp3jKwKu89f7ra88vo6FroX6r+W2ceBylLnPGTJIcm7bN
ekVuEYGlb78gG4YaVIBJfHdxYeeCEGUm8/P0gBgl4MTKWAvtk5GwMx1JNFHLRAtFU5QVEc+ajVok
p4GCl4c3gJQcheDjKe/UnI0uW6jGJoO/rLPZ8u+LbvqPBE3tnDjbwFTYgS2eRHDDuydbQrVVps/R
SjSWQHt/V8fxMf2YOrDYvRFr/tKZdVkI7IGobTTSp7iJuVbfD200kIQ/hCCDpjYb92TPY5DpW5yX
Xdgh6PfOqqYuQn4B0xRu1wMyu67bgd6l9X2VYBlVhyV9EPCg3hNvNeXN4jNdphdYKOdraPZMN+q6
EMhPJIphwTvbmeTgYvm14iorbqYG4ri+fAtuV+Wnch0amxLTcnLBBT4iv6zgGbrJv5Uj2359Gchf
GgsPlodD/7gZnOdYniFQzAhn0KnzTmPDNOQLxgzuAV/C8NK3DLv+7TV5PG1KqO4VE+17F6rNVn8F
FDpXdLxHK2rBUVMEHhv9nXt5HP69ViaLx1fb+F0YaW0X6vz9Yl3jU0L7UvEjB76LKJFM8VJyOoN8
IWkgotQWH205N9nhsENfxXN4WAICVEoELqdAOTxkIDFaHt+ltAxAQkAPNo9Pj4ZJeAsnPasTYTrG
x6xFxb9BYqIUQkU9L7lkJpFZqRrkxWYKJ0kbhtYvmpgq4QG9Anw5U4U3DTq8A6TrUHaC4soEaJyI
nrUSEzItcbY0zOmVT4TH/0+X2QnWRe+YXOYmuNJGYxeC4NU32VLL3RlV8yj1QZFNZ4NDdY7VzSGc
qICscWV1QaV3tOTHAcjxHyTtM+7IPuBdIwmjb58q7PDGhO2XW1CRBGpnXR2no9d5DFHA9XKwmNPw
YJi8z3ypYle1s7/WGBz0y8aD7fsvXwCc230qr7nqigG8U6xhmeValkLtXiYQPY8GzM6FI0G9i0oH
GWvetwdYc8F27prh0ccV1qhHCmze0q5U+1XWjo4otY0r1PTHN5lcTzZj1ml91gBmTDMWkoglLo70
ymnJZV2fCZHRgOs3Xr7Zei0S+Lc8xRYX6n8dcDLmUdzIJ3ROc5xq1Sg+/tm+qhYxQmTiaxZwhBRA
Otlga9dRNem/4C+Lqpsi4LECbr4Axzmr+dLHHJOnGj0pNm5jo97hF92ruI4zkb23TyyVcE+3mYp9
KgJLPNJeoD8GLOr1fcx7MEASuoyU95Sjg2i4FJVyAEy0wyeCnAzwxyzsHtLtEZmM1KEIUYDIOxVv
PiaQeihAOK5tTgHzTq5gEVld+1Z+rwApoo1eF9LrFrNKD7EzB5TdVOEesYzvKsSE6Jx56l7LZfum
tcPAu4JgKDiXbSP8+3oQIIw3AJka+gtw9YnWDZmxlx7Ztpid+JWB26Tp02NyliJ3cSGcfqWyPs9u
RJ4ih/SF8CgkC0iYzszc3q+qGwaw/S9dSi2qNp+unx2I5ZIF8enfTYGRNboJej+iS0f6uShLYqXG
hSP8cYm3PPswqa1bOFr61FCinx3DKFeiPYjKo4QT+aziWCfxI98aFI+24ISyjF4IMuvIU8Pgk83k
joDWK/7RlEH8tTbO+u1jpuX2DkVYZWjjd2CNXi0/PNk2IX8BoChZio85biEw9+/GqxECuzqPzyUq
NZlhAHuW029g1jB/WLaU4Qs0dpI4126E39P4pxFbtNX0faJCLuQtu1JA/kPVVTidPW+exypLKRW0
cMjMsYO/CFMGhEAfaXjeXyAWLdDHU3LnH2eUjFAK8wtoxCSyvDPKIQaIhRcqdXQXXUecPOTOnve+
yZfAWFcgyHiU4Fi/d1IXb1Cev3DwhHvQ2Gz5dm7e8JxRzLfCqhL2mMlx5I2ANz7aWpxfRFO9MuXC
ghXMwooesn0kPAqr6oWCHUDFlnu3Z3pYVqRWDxJkmilXwFbEzJ4CKXuESQ4sx3hKhs01mC1KZBBX
WZshiHLV7kVnAVL0ckoF6uqUnnCb74v706g2lfhd3Zt3MH2Yjxr+xOhGukbQjXOQ6eGBWsxYACb0
svs0ciH+871f0tD/C+tBFO7uGjlY2lfc0FYW4UUyn4pi66TGAt8+/EWCEVjA3K0tUc9lcMztDqu2
wPPwQz2efdvirL4XziXuZor3rEOTTsbbuEQR3lVdyZMmVwCOE3ryCT1XmmpThF083Qj8fzg6Zn14
G9qafB8i+fDzghUQSQL/Ls26GxE4Cv4GwQ77X/3ayGk1r7Z/hW6kdtdfmKd/9OK06IhYlh+Lpie8
neaMqnQj1oCQCJJyL1dw8jVSrYlIaP2Qh+NiGUTWgOnbw4kZKe5ou8FFtpLdeFa6p/5ynSisnHcM
qL49ZAKBO+PrgsLi74rnL6LIG5zUsmVE115LxzxWPqilHsG4qI0wPrcpg+G1OfTwn7V7UlrzcnfY
QJPWWNb7Xsg+AvouplCpXZfkJtenZJxwRI6AWChhBtX2zuRiYAwFJVkab3qM/Q75xOghOLO6T/Oz
6M1tGR6Hw0Le4FZxTuYQ7jA09cC1lbZs0tL6kjPjEkrIn4epNhhsNZX5/kQ0TDOQI8p/uvKwNNhd
Xr14C3ylbiBW4YIdAWGu4avtCSvibUsKlxbiTISuop+SeAcyMp8f8dIcX+RRMaJBRwrQXOlBlt+T
f832v8Gz4s4QgaW2m+irdJtL4WUteRNTXepIHc8edrCfWjSZbwKIb9AhG6egNlT74saHrrPmBYFc
SqmP6wjPibQcNO+cihWj5CtQYGj3AmIHL5VtIk2jbCOi2bekmWW7PMydGoR3+jxhETlrZAzE5ZE2
g4uObPuhosZX1uu/lrObPa5pj5s0JQdnVUyZ/X/1jAJmgiIYTzft2ceL6W1iiOgvWVIK3nD9zlRu
g0u/HA65IPhzx8iZUu82HvYJrMHOszHF58FqtqjAVDM/v9JS+boMdk/3gH9tzH74X+ICX0MKDWrR
JEvg5MlrXIpgSRv3jvexi8tvbAmpisU2ytqJJTTMuUewS7WFwJAXdq1Zgm9a2qIcbVv3S4pCRLUo
8ljVNeQxtFBON+i6StgQSNQZr3RE6oIqXf6L4PHi5do7b4ancnQbaSbi0sMCaEbhI3IrIJ1fWOCw
sNiEarYen3qalHzyy5p0PBQxGB/bMRNdw45GNsF1K7b2bUAmUSoPIvuDarPi8tuGFGNlEVLu4GTD
bKrWS91WAYTj1w4/9Z8n8YmEruha699F8fzUMwpPqSy0GIkGOCtMWD1u6SYbf99jC+WwsoNuPSQi
I/hRK0GLRgOI8XlHI8dX8CBtjliuaVCPHo7BNP63ilkVhOc9cJE6Mm0R46/bjMU9bGMSX1yDJqHf
Q4QElN5izmitIS8024Z/TZJUU+Pav7bDMQgRN3EGKyX6WcTdKYgtEWdnUem9sl896pD+9ltbqQ9e
mAC9wDyXs+gvSHVkXwG5GPRwjGx9uC1GMGElawIkqmFHCFT5qQEX+GPfEyN+2xRJDn1i7WhVlHgT
NSCMPtBgapJ2ZFEgHK6QoOwltiJ2ivoy12TIz5yLgewvuBCNUlxzi6ksg4X3R0vfTx/prGznpOiS
VdRrwLyD5RRhGcxh0IbPF8uoQx6agnkGKmo6yW20NejADKf7v1EvbIrNpsauVnMRjK/T2oIxHtl8
6u0K14gz97OXnlxeAS+zOseMkmY26XMrhPDcG4e5WE9Hfg6iVzSM2nqCCI1uSkMPq48LzXVnxUO4
WjdW+AnH106lZdMKejqTI5y+vsQwp/20odef1eubIzfPjLWwBtgSqSPUgpKaVYK/Vtp9LhnY5grq
eB37uepcSZnGLGCPBOCABpqXZK3NTe1iG8Qq7DnecT1kYzTcRXig3QZGTqUJCdRlxJ4y8pS/zjkf
lnbRApkBZfXyw7jXTyzY3j+5KvaKbXmOq62b6mXpMXn+ngIVMV/IuJio3NYYh5KBMtpuTd6eaX1N
oBbFMyOmv100+ZwpUTKmpU8Q8WUO8j3bKyAeXqapT8l7u37SjSCwcK5+V6s6g9fH/IGuOUnpmw2v
CyJ2EioUqB4/aemWwhh3N6Q2cbPgEwIfsNHftDUC041PxeGnpJTzTBjIEssF7p02erJ4hDm9Rk36
ZcXcb/hJck357CG8qTPVm4SGuF6OeHXcmrMZxl09v2EjOH8i2wiPLF7MGqrVSP0l8xPFUm9bxYRx
JUe9k7fGeEDB+omqJ3ytnVxkAwjK5/YCnZMNhjGFe3FGy7fxAlCdTBmTlZwSEKm1AziSmyZuhEHe
QTupbIsxha2eVAEKEwNzXdm/e/+tvdurztSu6Y5b0N8kuVYgiH6bYAFlxB/Vqbf7Uzz5Sl1Ceis8
cqt0ENnPeNvunS/3myD7lu3z/UmxPeXC3x49lfGHUp/DdQgQdpPwT3FPID1dA3h00MLyVXRhOGUn
qmMLWyz/ojLW8ku5B+LrBepl71cIvx3MbeqSD9x0Hjj1sUzmrfu5KeF9+W4zd8Wqm1xqjbs53gsV
oJxRcoskp3QLcMH9WjkLZjyBm0Z/XV+Y4M54k+eztLcYQJoZX/uKSrt0TsekX+ppmCgJbp9oOuwq
MdMQZtw/0d44Ou03+PZNB6BQvSD3D1/ubzqp8OYt1gOfZUAy4bAUZVzd+i5pIIKSijF+wmziCqCY
TtrGBKNh1tPmcYN3Fd0zHJwqjsKs0I+5D/hsZXeXAa7zotFSJDfijGp3Xn76Pwzdw68SzTYdG6rd
uIzQ+K7qSFpbigVtl84TaTaA9sPO5qOjOzvroMoUUlOMA80uqqU/t3Lu9RjQ6egPJuHF/+llPC8O
BgCU3aMw8lKeyby6fRPGfudPZAQeNlgQHtmghSIWKbWfss/hQfYn0kX/X1iS2bvHG+LWsUPLznbR
m0BFJAaS0ErWU8JFISfUtINM5MzTVkVUai+HVQI2DpGpFDjeq8Fw20ojBaWO5WNmxc/1FghWnFJo
xo3T6UASCFwL3X2sdNl+VsvmciMYiNhMrDzchtMyQ3H7jESVelt537SvOclC4uWPvsHJWvVFGj+k
kKQXkHK1dVC8O3raP66zyVx7YTe4285uIwe4z3vMe1c/pi6eLDAcXdw6qMS2JafFIE3uJwio+WfP
Lqk9JZDHT/lLpbhr554wA2+1DMIyQfDOpfXgNm2sC5KKuRxXY304qi/mqyhnuPqk6EM1B/A8PJqR
NSxY07DQOZgPmDcC+ncll1NAkQhcKWV7biItcSHxrSb1/a7+XYWY37tg2MTLHrJoXtw4WbNbrJG9
eAZrPgLDY1a9C4Qf26htDzMcSAPBVUQ43/QsDijfs797XCPq1iTYdU4x7DfgHBQdUpmzR/yf9N/H
eY/3/oaE7TAiFgvoXMWWud5AQfG2EG0urXQBG4BWxPwQDTQY8q696Z3vFuA81VF301wfyuuZR45P
Ae6UVBVzJ+kpGyruT2A/HUShgEIZUXGMZTrPp0kJoA9WnDzXum9Hp5eRemXTbAwGr2E1+ipEPL9l
C+J4tE8BMoSdTayGCB6z2Y3/jJnFUgA9tOg+nd0/TxlMmLNY6W0cd+WJYAKHUQwbB1cXWdyLg/s8
F6zdEVTtPKXgfLnvji8/Z8FJzI9MrD0w6g+opMrx7m1KHeEpjjrV8nB31sEwQsDs2hXEIjexclE4
r2adctmlJ66SjUeTDsIXZfcItdr5Sa0CASaqde9HmbS0IgqIJC/dzjIukDGn3AWKhFfaag94Ckto
tf+IjPghaYXM1tBo96lBGmRNU6GY/Q9kTLD9VPXBlcTeCuveRxoMNG9Tu2Ly6q0RZuin2tblYoXw
hPTY4crvLR9tYe7tms7ckDSPPuqQL/Ih/7TR48PyF/NmDPVBOLd26Usp+UexxJmBymRi8pPsk896
GdlkiP7yr90O5MTUqI5xmCAhgqpyD/zQpyhKIa17x9sl15EKbF0ftwYTXOPkX0bSiKl0i9/BZX7/
T26l2qRCt8rk0bUKoMXMaKrAEDTy2XIAdlC7wrybd0VG5jM/SmFMR65xOclh65fbBXHxLSIC39qA
0WsZVPsdkUQHy3se01vfjDJfHSaZGao0B+mMFFV848tUsBImRkkjx7wNDhQoJ24/MIoI6cDXuC4R
OFZj0iZUIu1yrxCbVoojDj2Sde9UgI+S7O11ZMDvOQeAZwUToreyGLp2sS5K7slpkPjYdmSTLpnY
pqsAz/nSfDmHdJGambAYmwY9P3j9C3evkkTsfAMd9p42rCDenQOiPYU1BNxBYsvcOcaBesLCLztP
mAR6ahjuzHlqTzzBsp/PXv0DeMLvbihvS0Zix1ux/hAhTjy+PX+v5+dvBJF2An4nMh9TAek29iDM
YGVFrGMKixtwe85EMpPKrm8bkoy6zzKfOJGf1oDLOG/+zUvFetmitKD1nM7pXMRxUUYjenaXVX8H
jXxcwhyPQVPVZXhs/RlDBqMhuXFYbFrHk5jwyT4tSJfQrBzahhrFnjtgm7gFwMwH9s7WARZCKVwA
LUhukaMaTz1Qvpnsro1Al/UebVMAVmj518YqQ6y4apVEwyovLjkbrr6iujLcjwqwS3SA+VHg3KSR
ZLT7cwv7OmrjoagQyiyO8EY/5BMU88qkRFNBrTaUdzmqqHdJxyojWAAEYO/XulGkDMYQLc9fIgRt
ps60fJNaF38HWn1XyJ3syaOV0Wp0ROoj4GjBfswO7I5idGR7rk60QMitoETybjbwXKPIBk4GZQuE
D/zf7l8pEim6vcFgzAWsvZdJbdlk/tTnFRRwSfYrs9P+6nyQFMJ+VkNRzUrFrs+7tDvYEUY1SgYy
vzmYgNiWGY41VHKbpQ86ZhS9c8NkM3xRXaDq8o+97UQIc3uehfWNugirnacyF4VZtE9ZOd8XX11f
mABW2DJirsT7vfu+VCNXXMEzSmDj1qJ2UGMUmsY4NB6eRLbgt3mfyWg5epsFvzEKpNr2O9Yb8Ark
5ZqWs+rROcpb+JMK/tdntFn2fy4NvuwzUyX8ru8ONTG0vTXEe3dEBWnX+N8VgBIRDIpML9Kc33V1
cJsB0Cs7c19Z28dqqiBk5/7BgZS8YKjsbjnxcOaIcCGn6t8Z0E69tgJqb3InP+0PKdB09576pQvJ
efXdx4QE4Q63UE5I0E8pHmlaPJEk2KPNmYcdZtlhjwGQ4kFkd/B5u+AUP6lCRBEa/9FBu7AsRkeR
n6TmFAXpTNVXJpztwFXXfjP7M9J4hl10jxqcZPko3XTuL5cBpIM4jltnL6SFV8JbQstBlG8TvJXp
yRkMM2Z63RayYbHtTf+XqNtL1C9hFgfc87yNBaUzHC5TbBZ8nrmpNaG8XXlBf30F9dMUpTChii5Q
nDsllcBUPM9eTzrBzgrXLtF1WXxI3aP6NMGyTVjbJoj603nJep3OuT8VPMz9yJ4WEDdNWTkS/RfL
I+67u/51P8jat0TOEapFw9zHGrB3btdTqtpXWdVsk5zNi3IX1Sx5xoNB7ZgCexOs4MxSEzxLyUql
8i0sqpETbPyE6dfpxzXKx0Q3CgjRkj7Pj+lu32ppbd5BnRvf3eEbUcRcaXrsATySS+j6ZeEGrofC
px0/mG5GRfNpq3VZ5mG/OMZYLhQNGKJsZquIzWvNdwM8wPEbq2Bo7i0xZwRrtR3snTFOhSPOCIkP
XGZqqcrbmmUTqOMjaYCdHzzVHuqct6eZVBgbMkH8uYPQSRLD3UP+G6yovstHRX070f0qZDDxR69R
ClIiGmSy+/OxEadbumXDXRCZBJqh5ErWBbzU9EaS4Bush71jWZhM2Uuqm4DWunvqQsmUxxTsVgXB
Z8FUTrGvWLG6x7riEA0QbKCzEVEbTGtMbirSr+iwYk8tWQ9Kl0DHejgtWKAsOmTCMmqCOhEsYlAk
iVCmY2VkldImaHiBkyoNk3WiaH98Qrc+B2mzklTz/I5TYz2r6sTBVXkn7GrxKzvnia18DAqjf+Lj
eA0fqTxp2IEsRq65roAtx2h+KFA/j5emlSYqi3vdHNa6WL1god1kGacF/U/NINHUKbcXemXsct3U
nLmIFmLZa8p2i1DvvhSlD4Glm77iuNvrztU9wJhKxnMp6LYKFnwX9W0fVGdSloEZeg7JOJOnVSb7
Ir7xD4692L2kek7IGJIA9oaXFvy9VywiY/az0w/wymzsNwQ6kd+TYwQxA+3ZNAvU89bvZe3toWLq
QeCt/tHmWHpUgeH2T7bFRbBAJMNhGwAzsmy1VU4AU5UHN/K9fkpexvpfy6eT7O00TW6m+y5VTw3S
7qs9vzdMikWnWnp9bQGaZ1JIn81xbtPk9tYCqdwVkFH8bZY5HWJWFWRgAOiEaofYT/ZOyh08iwXz
uN5V24NbHKECIUFamGnuJKSQfYsbMP1oYWlxM0Igq6btdx7D/k+ef2yfp+DLkezDGuOAsmlmgRwc
pjlO4xvA/VKjo6PlIP8UbXRUPgyQC+/cwzIWCVZbo7yra4uQEL1f/iA0hTLEmJJ/s7W//R/Sut/q
kEnc85MMAxSnp1dg05LPP+5s0s+42gnvwUmV9n3UY46hBwG2UN7OY2K63Q9t6dxqlzKN39vJzmHl
22Kgdha4fg8+ar/sVuGA+L70bb5GHhNUXocq7Vn+JqDyJSiGsqdj2xKt4+xfEc5QQPiYBvVLWiij
zDLGKrSOfbd2R9eqWGTwJfFKWUOvRk+Y7V2gosx9JgTGlIjwfeHzb9cyQdZBqhGW6Z13wyAsTVmp
ncgJ5/Ds7DNOvcQvkiMMg4Ke+R+qLmeEfYTYaXE7em72uxLIfwHftEK4z8MboQ/MgQNVSa56+lWO
XB3W4x5aYqQAU3zFx9W/gRcd7iLo5niKx1m7Tsuhw+EOhTUgAMGAlDmV9Ak2V2loRBX+ugyzsoD/
vnpm2YyTKABaYAyutw5pOrTrS+6S3SXuvak1u0foy0B57e94l8QohKodHaEHaIN1qwgWSpZi/bem
fQ3934Q+FvNxkTC0+gdxPMGPnBx7rRcYPWQiHYCZDnIIH5WefTbw2w5g6XE9u+5QyKLqZzwklueD
/Stj9lU6c8h1Rz3TJ4A4iDyVQoNW4q78K4vBmhWTzLD/n9vw1GYeDDy2P0+gBIqbN35bSh+RsCBX
0YiXoG1aiKqjEbZEXRpRg8kn6LnfNSqu2LqcFIknz3E+wRgn8G554v5t1ApbzlNlTINxNYwK8lis
8+PM682d21JGw3wCqexABVY65D8MEG7cNSzdI8BkcqPvEuC/AwYrcUmqQbFS7V0GB30AYJbaC2+g
Z3ekqi99fx72j1kQ9+Q/j8Br/hV0iKdTIItjwVaHm0azqWmU4gAikaxi3q+qfcRe7pRfUG8TRCKh
VDhCyXf1Ic/70CLTwLJ8/bsqpXwOBdQiyx3NYzaah6olMbefS35+5FzKCBInNeCJjtUApsP8iZbK
lyf2LRZPH7HbSGRT8+6w+iEOBYJHYUz7KB8zHhyMqeOBtO5etU+uFOPNmoBo43V/xyvHSIsOs325
QVvQkf5r2M6pjR2K4AYuT3yi6669/v48+7/JHMpgBY13hC8UnHixSQL+LqApqYzvId2VK4gwhxjU
By0BNQ5OIZPfmkahVxyy6IXTNT0Kni/iHDYil6IlfRXnJjlzDuNLhA0Vpn7Nv0I+E/ZpBIOUftoD
ave8zkfQeuE2b1eGiCSBSXlj9V6z5JVs23uWKEOcnGDTeEkR9+EiGyWnWSEShIMKwvNuLC+Cyd3C
SYbe/bTN3fIRPuOhcfKvDf/JqIPEhRw2dfxxblaGif93NGn6zIfmslCxxVD0eqII8ZRt35jDp3aM
KOtlg2SRJDY0ZZJ5aP41ueaTBS3qmFA2JkIOF8AZ9FrDeetd1HX+zUMEl6vwAWcjtZnkp9u5Al0y
uwOYh4Dq1MeESaOTtAEM0RLpbI58iouPuBIVJngBI3lgiJi0YAJ5xrJ/XzosLfdZyqgfed0mB5QZ
lMB4rt7Nz/wEarCBeOI1BGtRzXwJU80fNKvlO07u0b9gJcKCh5WwQ+P10ng5Xoo/KREUNrpPsoBx
On1mmqxKrBLKMFSF2x4e06LuqULJuS218EDzApwJ1eU8gnofVi7MSlxktdiWC4/34C4VcCtAPSKV
F/Uayh2pidzA6+cEaIxHmN43ufpr4ZPgrrUyJt3TG6bkVso3czK9eVysGVCmsy2XLjQgGZ4SmYU7
jxlA39p7FtNwsKTYLWdYunJ/bNvZRSDDOw2d0pjYVJp3aazoxgig+AgA95A8X+rIYJLVnZJqG1+T
hZQoAH/f/hOn8N22P0d0AKvUs7MqEuZX/FeVU/2F3JvKaxV9pa1oHG5EXGWi67Bg+MBmXckR1WCj
WPYaELni2rsnJ/lAMgcz1k0dBizxcGkRbnyB5NY3VExAt42Xpkzraok94dOaUufLjJv+bMKGovHt
p7AJ7JGRyHK0b43NeHm0RUm4cR1sxPGxAkEWC1Mj73eX4d0AEPbbIKao5Xxi17AbEHR950ViQlLn
/CCNa76JLl+MbM/UOmAvwTCojitJISRUnzEeK+BNs6XNhCxcZAs1s+MdmLMsd3osz7jOaJmcKFG/
OGbJ7SJgM89gsgAl2DIAer6R8+pVLj89DMuks/XgT2oGhD+to5uW/dfK1Pz5Bh70u3B2HzJehsfH
vx4mtxEx4FUFL820o6R/w2xefeyV3b6+hw9WLN7Z1mr35hA/aw9ElFPGvA6WGrmwoPmtX4E3LHkb
jxnUT3OVNDLj0RAok4MufNWBRvAWZ4pt1Ch+dwimu1FXKCwxwtdHtrY+6ika8ToSFs80kFvckxhB
h+ru5tPsW7XLMVSwHhtfMnMiFx2BR629eWu8y0VWBN7HVTJfzamCW+fM7hSG4bAUL4a3gQGDxE4Z
Y5MWwazylu+2ZO2GualYCo3q1qLx7J2iem1JIi4fSwcO79lWL/vZzCZOLGq+K4QIIXBXgyrp4lAV
EZOV62D/vf4IKQSmNoYrbjh6Heyt5uViRXiaR5X45FryTQcb8GjiZP35MB1rMIux1d0e9J36ORLJ
GD29gn7kM68KSCTM5Y4h7FYAKreDWb3AI1yarV4LAtK4p24z+kzc6CspUHKFQpohC7QM87fN5JGZ
lTgXquBeLMc1WHcf6wZwuQKP9wZWa5TpNFzqm6qeJhcbAL6kuivQh0gnPvXe8msBezuxh7vnoxyE
Evk1vkfpWAamwsizp6sHMSgVxuogFOSYlDTwK3MaK8U6WteO5QPbbnnvlDwIA5bCyvNj1o/aYzhs
jmVa9SuQJYDzhVFk1cnMh7OhC0wEfnkbw0i5w4YI1pdE1d7CVI6APHHgQoca1dqAMZvJoK79bBqo
lXKKb0okcfv+mXea577QAzmeIEI8wCSrTxcWaxbMuSm+R7RwrORFrJZ4XLUPZZWDvQykGxpxJZga
PVfoBkYLvEfnIiRxOLPW7v4N3zr6r6gYRbw5zzhYNrJjbnlr+VEZ/G2thHUIw5YSZuAQEdD9JDBU
MZsGJDMQ/c9zvlcUGyCXTRFyCuj98T4beEeR5ZjtfkQljx2YuVx2Jj4WRBF1w7h4jryeKLtEZZRl
kyRwaVX78ytdjhR7D1wlVNnqKzigOUHxfXG44L+eBY4opeM40hjOMfilpev2d30NJgrhOwlFJcfW
lIznKcZIIOUVCJrlV9u0irna8vBFpTIAz2NKWs07Cp05lP4442yXZQVb6hp7KzfRH8fdtM8uF0xo
F1ml424qCeLK8lCog+JOaFu+m2xv9y9j9LWDDfYN59jYglPWSpcIzTfA/Pi530/AqZ0jNs+GDTVC
j/3I8bwc8jFNbEk920moYyQy2cbtwzjZpJk4rGCfPvsEY114b/Ae1dPUTfKw2hlp4VAFc976Ixza
c1HeBvPX0G0H03VBxbTJhom+gqkTN6PO3ViCH0HPQ2D7JwK6+MYbeBmfu7hVVL3uc/X1HO4UIoRc
c7YYxmDaUbm6NEGaE0P5cx0mnAkm+l32JRUrwwnoqgYkp3bcnP01Nt5kv/BFRbhTv6iaxDwa0OFh
be/UDuDk4oL+60TlEauaKmeJUlkAatNfHaXSrV5g+bb3IqKIGB+Ucc4kV1s8yshSxvXFd2We7Gdy
To2p7Uda0PYxa8iinezywP0cSe29b4pH4xBKaLG6HovEUNbCROa69ArZtnF+qp76LfvskPSI/OjC
OyAJW34ahe6tjhZC4eW7xnzlyaUUEHf2b0dflS7VVWFva8UwQ8uwSQmVNi/ltF4iokEPAS05tdBY
Lg0fLE0PTKuB7VWaoDV5Y6H4zjGKVQmbj4eL9TdjBRX1hBlGPP2F4b0tDPkh2Bu6LVmhzITUM1vE
8xSDA1qS9f6udoaXSNMaTkGwWgTuGFLWwTc/T4byms9XIfIpeYOZF4QgSru5HX6jX4b3I7ZrSZqD
0ntTwu3w5z8p4ZBZiOSc6SwFmHjbDlFNFIuaj6J5DJ5BCB22DyWkAQReVdQsHrYOaOxQzqhesp6j
I7NLISzQ93LJaF0jTFv62iBLsvLLmi+l1YzaaT/Thzkc6Cij6j7dQnOhMPYEcl8esjAPFWunuFI8
Xah33IHk/EpV5WkieTtHtNEzzltHlhwtb3Z98zwiAHddfDFzfgDsECcGw+0J9mJ21Q3kexW4pIlw
BMPTfkehsjQEYuTaU2aBr56+mcEPjF3nLd7XpITsDU/+KUZPbLSfnr3Oo/Ni9GyEvGvOFlGX+4pJ
VrZcYPf+a+U4cm8YfSMflXxi1gEeI+OsXolxX5vElvjbaRuRUv8g+57UbxFBF4Q6WWeyODfKQQPZ
or0zOU0XJIWvtASQsFtBaDaELhyLJ/Vd44IqkWY5hGH53AYUL1EX4hUVsR7mbadC7/J6Tz4wPF7o
dD6+2EjdYNsQCaqL12Bk0bZb6vNkbsN3lyM27yJ8BIfEW8sAo/6jK7GlaMRHVbXqfLW66tnZ6Wgn
OAPbatNIimJUH4EAwA5UAd4HrtUBpB4pwYw+wAcd4ugS5arA72ERbd4089tXl23FHL05AfGGszhh
QOw7SxoBcZRY4VzB/CS5gV5vAcD1oJxfW69Go6WNJ96joDOrPOVbJWhvGJlbNUMlf9Lj1aC9/Iqe
avs9cBWgLCIVRIrZ4kmf+rMjr3siETYiBmCh4CyHxeNN4rnWhycmhcBYCeTYgmtvv+nsN1QO2e4i
OpRgwV2S5lxAAJ1G2va3YE8Jq1jAqwNrjhT5PJ02Qa6X8JQFbZ3B50Ym/RYRluvc/03CchrJCtgX
NjpW4Ig2zd4iAruXct+TyBxzy2okfdzL2fZ9EFzXfdC+7WCyvgA/8fZOvq87ZYiPb4kWnCbtufv6
4zcKWukqgSV2QLg/Vg3ip0sUxyH9VllDZ+u0RaF90gDJt4sxelhGOOe8P50N8IZt14tJmTKdjPuZ
cFnp2T0rXvkmx1JaSnkZJxJACcCRwRYb0ZbK31EquPWAD49KNr5k9EAMQ3Lq4cgUs1d9u2bN19yZ
8hzy9giWnY9O/JccbKkP+8DtFbdKgGAobrsCqndf5BQ1MwNHcePQALLMxlLjN1ntLUteSKDm0zlu
WbHP6bqlTz1B09c/1P93UHahO6YXT2bpnJnm9AMASXukOCl1WwGOpb6XL8LgYWU3tX+dore/Asfq
9EjqnzZs59h8+zPMSNE0WThnPFv/YkJByYR8ele+6wC33opKPkyXH9ZzTLyvdrrroRVBJcPJtAI9
ePhUBGK+J8dASiYDhcWekZmFRBbxztYdrUGdVdNtF9vVNSANpQGTlzxm41tih8dk8/wJ6rkYwqRe
OsYepwkt83MjWBibOP0eEfWPSW7Hmuhrh1z+rglWXJAnsXiGrWiq/bxi/P/LwC+8zz5YFnzA+rhM
imwfMVMqxw7aDRsTqE7EirOScrKgOHFF04d9uejP3voHe0a9fHWw4GTrIFih3ffNAJ6QnoN9CDTY
hmyaJIrGNgllLO4bnXuhHGWJREhdEkIUBQNpkr4qCLqp//3j+BHBK10q6bweOn4IQKoJYQmo48IQ
Gosj1VyD53p2PadFpA6SKPgyyRBKCKuv0rs7nY4T6mgK8UfZsDzbT7Uw8RTToMZH9cyKWHWKAwLA
a5OBEg2yTWCo6dfgdD3MFNU1gTRCXddWXWanDewJAXJoQddhzNm1m01HBDSDncJ7yLK/Vknw19Qk
wRHASTNPGwiriUJIYN5XwVcXz6JUV1+OZ4428+WrYvJHisTS45BgvUUpCg9EsBHt5c7I9kl4vb3g
83VVaaiUH8G4Mie4BqE7I+7ve3GU2lHH1nHjr7nSVzh8GQmGjE89u7k0503wSFPVj8UaPDftcjeQ
tQg7m/LY/9GIF1qc1bwbBT7f4G0vqPAoSWUzSFwrAOzLlL+EHlXwD98JK40XVwxelVMevhkWREXf
L5Bfw1SEuS/1Vq9yMy9F9tDRR5aYIRBERmUHLS6DHf2VxyNXTleq1TfC4UVmLmtxt3R8JN/BC5du
zZp/SML4JlEkrgLbpu/OZpauumQbJTHcgW/W0ZxRWEOBxRx67Cj0268iAn+cml3K9g9e3WCxv76y
cB5OjZYQJoOBz9F36eUH87855SaNngUf68mCuwH/Msl/EjPN4MYX/NJLQxyKOJkjvyUiD2GJGr35
D1WcJ4YkVuqR3EZtSSj1tPdk7HJ6gqsk8hWb/H3Bamizn89YYjRwiFzIPnP736jSS38v7YOTwK5k
HeYamdnSSpn966Wt2OJuqBCAczA6xfrW1X+OyR0bhhtnbMpSXLafho5ibpcPNi3W/sXG0ODlIWES
HQYI1MbYoR31Aan2ie364SYwqPW0Uda/JHJi/dIgevCOCJ4B2C5mewQbhuMouaW8YxNwiXu9ffx/
b3Brqw+OjBnGwEHsdDfSHu7fgt2hPgw/25TXyNW24Pv18xSDj6esx6iBIt/vMy0I9/UXr+L85Ilw
7fZbI1wZ60deYegfr3I2f2n/8DZrndX2PTuyjE5fvZ5TxjrovWYSjeIaA9JwXG7d/kMh9zwvEIXx
zAyyZxVQYd2REnQVqdWJA7vtl8UcN8wdXPKUBrK4KC5MCmurWWEp+EOaPusy3BsvlvBHB5RhmlEU
01FlpC93kZQpWIucb18vvAd9NK4PKsF8cR3hmHskbyUv/ICdilCdNsu+maJ9YQTI/SYNR263e+Ce
VJ6AKlF5l2Cs9DXd42ynl+ChmItidVbBZMmoSHVXecNvaDZEP/hyxdwQfYPHUeGT3dvz6kEmOJzq
hEZySmYLEMLHaVeobR1Bt/R8gm7B4Yugq1nj0AVqU61fhqdx/AnZD5WgpuKumYlJeW0GlcyCgcwl
4XaDTcipaHBkGQLEQgwZ2d9kH1+R43N4gnmTHM14oErLvD9cOkKpX2upCb7himP2CPwiTPl4qaJY
tpEKFQ9HqgFGjVY9V49Lq1VJqVmvTTR7HE2/XPSzhDxCYvnBNOgaCy3OqmshdJ9VoQuwsE+jfD2C
168miGnYMF73B1IMV3oW25EjxyJlB01vHn9Nd9xCoo1A3P3MkDDhtEFh3EiIdUqiI3b9iWZ2YMuX
GQOB5y0dRvJNSHDDn6w3Ogis8zboec8g34J9ejgiAn1kHtOsLs7GFhUZT1UXtUYO1LOxogR9ZDSJ
5+CBDLHf5/eTQ8FcxRlpOp2nBx49Xe1AIWs0fERdmEc1juzURQJnp4isQ/BXTFvJPf7vmjHltCAE
h2UPkPZNP6Lbbp93pzMyQaU1J1jGGrVDHfOMSl1FBcPWXiCs1Cv+Mjoa4I8CHoT9NPAnrTrbAXGg
MS7JTCpwUa2bKC2J1JNKxv8E4VLw9rv1igWcW372Z8Es8nhcK57VbEJIg6kqWkOBmWKHrHneydhY
q8kWmdMTegBINO4JDQW6q0f4kjv6edvr0X2bUh6P6MDNXuO0NEa4e2BtOh9MhlrEgbm3QF5nueuS
PHa16VoU+N6vyl93TQ5r0V8HpGn6GmP4pgmeDp5T0ZDh5APmZlzfiaDIfTWQSxXqzBrKFwvcGSAv
EhSdHw9Wn6RNM1FsOr14RiAXvKF1jJm61+D28nVWBmXQMSz1HwKF06EiEqrX1BXOTEaLHOu4corM
ZLTI2cWkVDrJt6cUUsg4EcxH7T3QE6+qPK11lf12uzLGogkmh2A06jICsX/g/iFr8g5pezFuQX0V
A1oiB1ndOmqrgRAd7CRkJksfxHia2VuTUUXwwzhx4dXGpBdJaHog4iX21J2TIGIU28KMBfYIuzpQ
U44ynCcLxWqykskT+T7ijjIoCWoa9P3xsCwgLKY7MXL5gW9ex/FlT+ewLfkd4rh/dbA2u3rPVM9N
bofhQeJFuq0FQ0g0anRcHKvbBVZggFJiaEwpMi7qH0Uf0XiKcHd0pq2Eyh16je5EOfWlq8XyZHKK
vSG8q0OUlZe6/fDiMu66ffjurCV1WuFKpCuZO1pzcr1KbN+QmKj+FLzAuU9+Uvwdv+2FdK2wTLju
RI+eqSfedB9FA2Ov//Bvf8rOEsWVJdO4YQuWCHn9/i7biXhlijbhMooDmjuaDncOs+I89G153Cpu
UUkwbpdub0QlFpczHxo1vucswLjqxV3+UADWpuRWDErt4/zU+wgaGWnMnzF33d3DhKqNMFeSWzkb
hwBT8JR4A0FOrOavmEzr6+a//r42sSfKX6PGQEDeEoQTrxDiyA1O/E4EcEXXh9lGumKhpUUm0B1v
sk6OSCAmAuJAXw3IA6oRZHn8c22XDSc0ytWUIl7zByFVzaWYOeaaje7wAQ4RyidAM9P5RU+6xdJi
u+60eXllmtLyk8IsbrHNzWZkdje3bBuXUn5KqWLW/CitslD2bPJ1mXqlVDBUm54veCK7HNF0/ujJ
vVYkPhW2JugCjDYgMOnhkD1ioaxuE5SW1AuGzQtQnn4Z190NTkdz79Cn6YqJCJnGa7eF1u8v4ciL
WgyDK8tSYs9uf1jZh3HnnlxSq366YfBT1dgh2/7b7/LMlIhb+EvbFDpR+hL3PEv2zPOtwPT6vs1q
Ac4uRLdn34L5B5Qz6WMb5MuPMfGibt5qgmNjqXcyCzslo8jKLzHm1dCmcOtoTmN5+oV35rcvKm+X
wyPhaBD2ewEvqxo+um80OPsxLlEZGWVC3CgGMl8xrOJUwi7j1ZPWKjrMv127jvBGr5tNuRuNn79G
SRDUbTZ/XzS4qqPGqjtzCqGLQetg+YJ/ayX012G8t+7NhgRFe+2w9zWq+cvqsezLpyn4B9G2as8k
9Y5NsXSWQuUnGv4SZ3zDXKgFFT71U04qVbLRai92ACMY5Y+QLD6Yq6mg1Q+a22HT4DinWROT1XLB
JSEoY8qRYTRtcMMy+qta8JVLJ/P+9iqOCfWAt+TrB2m9ltKEluQPBRolY99ZEj1RYJXKBNYQWlrg
wLmfBGtTHMESJhtNHQxMOZYuPqvY0fSSt03SNqlpAU1yucKM/hfNNJWP2WMRTbkmTLXxBV20Z007
cGbA/gR+954Ho8RsObBpf8cMM+g9cPhI8kD2dhmBjdwrWDZN8qCGkM5fJnqe4ghQNyOrs+rD/m61
rI+FqCFjy/aGcy0V7/55gh+66PAbL+OTlUcgVewR/EHiPWvIm1caU2kTY2nctS48fHdP1bgevgmd
bH6P0HpdyigJNtnTLZ4DI2k5Xe3gnxZATrPe6uelQdHPnT0CriKP7bzA7k4hTQZeky9+Sp9AMXMG
Shpd3tWYHv/4iF+S02ph3YSSjCY87FK2+W9/ShQGhRVzpUBUi3WtVuJ6t/xA6Sc/NmbawgM/+M5w
hPuh17F+Jppe4c3BKhk8Hynbwol4gGh1x0LUP5sJgKoAGY6Hnnty1YdPPBFdVquQ2z/eIVqte+WA
SKpIKfqgfalTBqUkCodADiIRFcSbiO/IBYVljthN1vlXq2Xen5Y+J8qOSJXki0fG7wK+18GLN+HI
2ZCX2QIB81jm7NcBIgLnKus5+8GISbPkEWcJyvHhzqpHbbjGN3eoMikur0GETU8MuzVNGHRitiC9
q7kLorkoSlkcUJF9oI2btEIXCaks+1YvbtPzzv31Oc9CzLTsMWLoibZwL0tJM/Zva1R97qqvlBpM
oAbb/lIpDqdh2TLu1at2flemcIPR0HxQp1jYcUm6hwYPM/OGpJWp59Bq5/+GsU0viF69CixxkZsk
sUhNTCUIk/PRjpG3wBTqubifq3pIok/kVNRZAB3ahzDeQX4/Y/+NTgxoRXGdJPnLmunDXXT/3BAj
QKeEqfCojpgZYjQe7f5x4yNFD0I3y2ZAgShtUrEf9i8TGbMwbDg6oUQlsyfj06jqecNHCj4SxzX3
oPCWmXcg+VUR1YUL/avvseoO6Jw4fvZtWxjbqd7t4LFw37cnJHzT0A7pM+QVdlAN9wMv4R4Xfvze
pqyLzyzMwun+WnKN4AYrW9epzs8UeyGz9bA1AHADnhAFGthprl+e3ZsBvy36QGPDdlZLV98X1icd
7EghWPxX1jZoA+2LxEYg4s6Gcne+rMIt4e2Wta78YzWOrsyqsF8FqqAEazMcoeIUap5ogNQHIElC
XQHGpBhfK8rSDcmsyFQpF1PdlLqRNMnQz0pJUlCX7t0r5LS+Hh+MG9VEgFRGby/+WVNpnRjuZrTa
WgW98qUfE2okojvJS6Ust2Q4S5j0lGZoNwIV7E4J5ShxrzfVkU61WUDLWCTQvB9fAGFVGlf+rNv/
mKVp9HT3WXlS7kDeF9nkR4l+PQ1aQ7HV8Ot9F8zNYboaGQc+Drm09VIo5Om/DZcVMlvZS3tYxFPr
MB/vLRaFu823xSG7Rj1yFhOS7/MdvKChTNa5EQzvjtSTniIGw9QsppBq7GhJ0Y0DYdZ2uaHLlE9k
OtbjsVaZ09ExIoJhrSX0Yq79YieKkBL2w+lkk0McMigKB5VRJQEY2Ko19nqiEEXqnym92hYInIZp
7mnjYl7V93sOHaOUhe8PW4dipHsEcEY0yqjGf/kIsUnZ7/RpBzr+jK+xB02gxzUD7WoWcVRS7v/i
tiBKkXhGO85qmkq/b7htho6mwJSK2pWJVylUMLL2Ty+bOI+BtW6svp2b3dgO9ZZdAuvjzyY8W+dH
/1CIKNUqUpuKD2kHb3eALcOI3j30mRmTHXxvH/jTsLgNqU0GXGhizfjMzptl7pSH8Qvy1lgbstra
8tim/FFYstwqJpQZf1x2VktKhoHH7uT6EIuORM8NnEZaNyFonGP4JlMqlYnoxNYsaaRKZE7hm39N
8ltMuQIBFS/hjtsojyAeOX/XsAOFmcw2UPOgXsYjL+b/NoZEt5tJ/BffzTOlCx/E1vgG/kTpE9AW
NQ+IQUxLQVJKcC/DDZddk2ZGaSgNxqdDMdwAQiLoAVY7LS9IXurz8zqX7KLlldvjETKlZcSULuoy
RaomCDcNDct3Kv8tbMyhvQdKaJkNDQB7UuJai6Ht9av/Ed05BssqEXx2uuZfnpKp+RJcsNd+Do1u
MZsQzQz+4tbuTrpTpRgb8rX9ZjgdSR/gc9oRX1NlVGiPpaCkR3m3aIHD4jj/9jTT9MTk8fCr65po
s8YXKHxZCQh+V/EuIgm/tWK5RnmHLp7/U0f1m+rpyaMl17QhTi6/7VyIhKfd39s5I/Ctn4x3CO5f
avNFeZWBQhRs52716M7NY1R6Uw0gDu+15IO6yPn5A/dlZscvmVFGdhYbFw+oZv1tC1xTmKIy7XfA
Nabwy/7neW83S/jx1dizte4g0WB6fXnPAsXlw3M+Z4sSatB7pUU9G5fIBMg9mJEUG4rRD7GB3EAD
QadXHKWA8jnGTEJSNd3DJbIrUGxa+lhSGXqHC+7gvMfGBWwSQBQrZSFPfIN3k5vXS8NOR8VhTdAP
6/L7L6pkPjaSvjK92NIEP5r9P8kCYTWeEbWKDp5nat4LOh4oXXw1kui0uK4bqhN5SCUPl4UAcAOQ
uCO6SceX1w/rBijDA7lWyKzOjDF608E4yNri3nC08yJEJPGrEI5asCYqz4DYVqogyJd6xCpHVqxl
f+oiMxm+lpQzQsGv9K8ZZLXTUrc+Db44FbxPj06vXCtbc4Ghp69XXkSH+oEMSYLjmLJPQfigC5++
o4PEawl6KrUAQZ8xEEP5jS7rmcPf9CWe72rpLJ8EB4giPWCfAybosHhu+rKRzWnAStJjcjXoppe/
KQlJNG4HGolh9F/oFmTIcgARprq4XNzZTsDY8IqiU6gmPlluJhVmA+lSXsqKsfjx945FzhKaCPbF
WaTPHS1nEr2Drt+FNA64eDg9G87HAhT2/99bqg2dvScpmbqNRthHQBR0ogQpbrRJAGoPeJ2CtDOQ
D1aYQaex4J25s1+hwajAAKoMho9rgqmwzXncof17orNNmVvBnciSaxEjyNUXvrj17y64capQw296
OkMLz8JNsVMc3eY5d+BZ/MJsFF1YwzZZXE01D+Vzuf/Cl8QDHgeP0D10oAI/R4BaAUbXs4D8cVY2
rQxIU/MH/8iYNtJSAlkUNgkqDZ0U0DONpWqBAyD/Ql0d6kDOsxCVymJnsaXF+boFbZrPrssvDWCo
k67iYeX7er4o1BLvRKmdnE55BzsnEIynQQYzV7eCcikx4VTozpQPf+JVSUqj8XlYVSmFpHZVDCb/
tvxW3xBKuVvM2RSw3fe2ujHp1J5usxiKGK5i2mAS9rBd2MV5WOTZTs6Jbk9Ms0yJLfOOVZ/ScCyL
u4mrvR/Y2qQYV7t301lLJGSGkuz/8ntnq7iaUgSnI3wFs/z45h2MU8Ig8OaCKayNyI/Q/JV0lAsL
GWU33A2m4++rW4fU2acrT3/Ff/DculIV7wPLMSTbCi9cC8jBjE5qGTdImhwGr0GMj2xHWIhqWq1Z
Vw5gGhpctG8Ei2615OgimTjuLjWRN1JJpqpWfZ11BGdwXrIse754dJcfVhe7Z55UJB38oTsIW2Hc
8oAWBLPXNbFfWocZaVw8kpsmk+6NUgRxjKKUx1rPgpqaO8w/bu4lS51zAzLl9AyJQnV1GTf0WBN8
Usagr12eNINzLuVJam2/trCsd46yAD9c9JEi5toxViHl4+jngNPZWKA3/DcrHSA2AjnrYKfaqoTS
eDKg0NMyfFW5uDRHUhIEhlzO7v9IlVfP3u3JJgFi432ISkm0qtF1IPK0oQHPN1kFT9mEt6RHXB5g
IkpG8TZ54LC1+AdSk4AF0s2BHImx9N31y0vfO0PQ09z/nFotBR4G+0b05N1ec+0PM1VeGeAVYozx
FK3R8+hpzBDnjaEQua8SIGrCjej376dAQ8YihbTSqAe04LPgEW2xsci/1Ue3nH63jQw47e96QkyO
sI57qoLmwZoxd3UXQqT9Zhz56f2JtlvCdMsyGZFsd/GxxKZ0TJe8XxOIE7Y+QILWu9Q2uZQpJjrf
3ta4rp102YJw8NNrFU/OEUgUTMQGhtlgpdCDuIXPPAQszYbFkcOn8Vd0Abv+5NU9ddseFIj//fDh
VaYk7sF7Ooh8SwryTU1hPrab0+TMPhmSn/Of+ZHr1l02akkWqGzdrBq1XeoUSvwMkWzNPHCn991v
uMS9tH3NnpNQFI09V/fH1xvYIoEJGuu9CnQQefJTvQBT2Wg1lZuIAuyDtox6t3UYF9EX+Q7nx6Zs
dJBXC5BKoNEjTos6MoZ29tgQGtdIN+VFd+sutsaw2Zmbej3JNzGp3MaWbi/0UL4qiBjVhXEs5Z64
zBrUSqbFl9LGurjXYKQQEpHmUVdnbhZU8NhDjL7yhroRIoTYHkUBuhSOvPcFL+FGYZUaSUAedPeq
sHuAl9EBPuKPAmLO3EKi6mDuhy8KcWoy+uYG4VdZDxghWDQFl75VPng//GEbQcYsVtbmrGq/C5z/
YLUTKiKKLHndpuOq2Fi3F8xC6bvBFX1NdqThCr0MZcI+dv8Ogxbkq95g5oaLA0s+cIpiz0B7dJGK
sclToPlnS/Lr03o+2Mw3e4D+Yx7GPicT11TKKlhwpmqjLIMj2SJ5y3xiooKztH4WHEP5PS6q+i0i
tnqcYAv8FyMxiUdpNzEIkQ9ME5zV0Q86v067bfORaVBkTTij0dmjNJiPpzX50vDJaaZoK2cjVpSG
GnVxFtfzM3R+qssGx5B5KAykH6MoQM0ZUG2xkD3SaHG+AL3fTdwsk0hBMDoVZH88cyA+Ym9w2EG4
ISl3xM6R/T4VjM9BBbf3e+7ytHt7CLFcAkOGjcfgGScJB/5P0W1MjW6QbhYwgkG13GWxwm+ccRd8
4WKNm2vdniH7IN5bejJPWKxHO6ZjeD1QBzv3wF28gKklmr+o3Mb2uxiwsu7XjS+Z7Ze0454lNMNx
FVrLWGhSZ2c7JGqQAvsR/OODCAa5JvqDHVytTFiG0O/FxX3HVbJpa2x63bY+9mLagiClZPCXmY/c
LehCaa9uVpyELdNxca5Afwni+QwRBAnwrS0o34nGJVWJZiSqXg07oezc1GimtYh9LJiiVcppt1TX
srEVBgc0BResTX8xG6csFz918CtaNPa/mfvH/dVE0IaNSw5HA/+LEVfhl35o9PvGiekU+Is6FsrY
CnLqB8yT4E9Cs/LdS61QiYlqLM1gUOBkNBTfoq8oDlhMiJDYm6to0+5s49deE4pmcDBWNp/cfnpb
+pR+RZPmAqgLDIIerjQM0EU81w7aXQaVHaokQ5YrJqyJmyAyFB1yJ78U43M84K508hYlZ4YPyZPC
RuNO8omUoNVA6rbNFoTMyAM1vX5kYzf4dRZh4w9mlsQxn9GO4yndXDW/nOIVn0lc0LE9/RGsBtiZ
1waHqFybqle7lTly+LXhaJbY+BqlM5wQD3Ph4YfJ65HEp4RhWsfZeRfe5sWTV5OV89VqrwuVpuU4
MJe5FVbIn2xnELyx17wlsOdSvbX/aQfpjSPfxXNYU7AKZCtTJ2Sp/aA+99JZEnS4c6eMArl/jPWA
lQl2+NWHIicpcMo0FAaYHMgF01w1V7f19KoAulxK9K1GiCs4r5vYDx/Onhm0O86dwFVvy0aPp+ae
UA9IsHaMLdKxVUxUKhzXAPdfp7wjjePk7n/TyAoKjGBhObAtYeatuoTFi3vUY0XaX5lx/0P1UbPA
1AunYUiV0QW+ETqdQ+4cE267h++dqSZWK2tN92eSkRjsNUIOjb20EYXULdTY5N365eXkaE/6skiI
raVHO+bjgtkNCo79UEzcdixbs/3tg5sqaPFD8zV1cPVppbsVD5uFtILyEjQEKOJ867R4cEF2OtO2
1J5UE5jrpKkrEyjiXWkZhd6teHIifxihDcFaRFHy7Mx3RMmVdKK6SPtYXYRi8Q217jdR542O59U/
w0gpPCSu/5NBc3ip1JbXRMs9NaE/ZTEideh3p/vGbahxHavSMhoDtNHLUGr1qO11da/hwpB04rb5
q5JxLgEyjEHSPbAxtOJAiZH1M89u7u0c002FJYu+W5uXiaLlzS/eyRBhQ7pjz5JtUfPKwyl3T2vC
Og41UWHWTfOEuckps6KGfltFir0/avmCxJfGHwZ9Qr1gkk0VHZyf/WpJijvrX9Kk2n8hT6SvlyXz
ILcFVovq2TqPBp2KiehZMc7z5xXKA66m+yfALaca5mgogfLE1EwG7T/W1xl0ys58dYl6ZSnMVBlM
NvDb8DdTxdu9/XfKdN2fsU+TicBSxrkNrN6vtWxDjxzBbkVAcBpTPyB5UeMp5y1RQA6OlJZ7UeIe
+5VPeHr4MXDeXw+obb5ehX98bDQM2JFbbWmQY5S1Nhp4xR3sBvK9ELhTLPjvH05QL4el09SvSVnv
UVl3wjeE6GvsIVbYA219v4z3IkEk5PjheMp0QaVvxIiVICNz9DF/eFssDbpSfCWCRfOs58/n6uco
vOjJsHfezVSMV9LPo9IcIjqUmKNGhQv/dVr0Lhr0uoaqFDnjX20NMqH/e/pSgPouyceKdoy1fStg
IEt5d25hoyRz+IY13ZIVopS5pstdS+ZfqBmXO+xkxQXIaDi2NPY4ZC5Q8AZeu+e1+JdwuvXaVIZg
zHtu+QETR5vhmDJ5X/EzkxuWxX3x6G4FWlHXjGRT+NyYB8un6AxpLwzKfNYyA86QACZCR+EPvOM3
8+ya2up5wz8rc62egYtsbNc3PGyYF6RMpizwo2gNKOB3AHin04foq0yKpQTerWbbHH3s1HmrhWUq
EfTvmiv3HIi0yGZAtCL8phvq5uPpmneELEpr2HIM7cErkcFeRpbo4ypVjznwPZ1RgNypo+EKNcCK
2EJWK+pDAF4ilO1vwPSususw4mDUYadxDwzrUT6WcPBwsr1P6/fEG3v3teiu7gkLeO6BMLyi0Q+r
aUW+4nuUkK3jjt5+PZa2Il1ypXJx2zFGncfdYRkaULiR9B8eRAp4QDj9tZr9WJLoLAI2VhFBjW4K
4f/L3BtubAr17e0bZJNxZ0yIrTICf8BBqYMYjJpAgu2MzdEz7gygYk+mn0xFwDqC3CP4crGlovZE
u36bU43QEGyM0Vb/OIb+NRTskHvk+Jp2dy/YRqer1LdrjqPOUfJ6H1lNOav4EQEGDVaHybRFBdnR
SDb5Tqs0tNGjqVB7cQCmqhDWIokPC6yLaF055KUr7OfH4SP10q9ag+P0AU096iILzx0jqXswpD7S
tm5nd0GM6VdkV+oLlnTHVZXqSc/GYDtOCAtkIgnqbqkuKOxX3a6F4MlNrO0Eb9+KcaSYLj6PH0un
hBTDUd9BhzMp8zam6tBaBIczatDs1Z1aouig2RZhwiux85MBn6F47wNQDVLiiIQ79exHeDswWXQ0
2EWO2LEHtlvdbmJ2YJ3/kO/WTffdaZNZEpGXEs/DjtkVmHHYqRgjYiNS0mI6i4Y2QhGL+z4F0iyY
rjfPMnHWSSt2tz46DTivKmwlaDQ4kFCWGvCiZ06dDnfHQZ+OkTJ3zrmy+VVSsRKWIdZEgaTGeCRA
3YV8paJC9GixSrPmPfFVIDShUP8Tjn1/PrTiPLJwcDKq5woUxfacsO4siH1s/1oJ4AMjAuKQhJGi
rkUBRcQSlMyLE5JWa+sZ+O9+DAwrIcR0d5nTGiRGgkHt5il108uZ34Tep7ibHcM87noa2ZZ/6i7n
4dWZFmqgC0bbA+Ibymiv9xuXq85aTaNpWDHFbO7wbnasdMf+5pUwzBkNLObtl2S1KcUtY+gW020S
uIjujJ/hS7yM9SMJGi2LCIbywi9fH/+hsg2AuZHdtbpsUwev4tj9RAMlmcJCui8KmgAVjr7ZEJAC
w1PZrtvj2BHeyFma4IC+L3F7YyqqXJr+D2sF7Ch36W+ztetP9XHpEQsV0L6TK2PZJ14KmldnJYyU
txqeWcRyKNuKGuYK4ZyyDtUQsGIuBLchCzqXQtd5LvhVheQPIip3VkLUewcIrffqyM3RnI2OxK5/
R6PoiqbdZ2vh2WYWhZNh7LnfFP3+2u0M66bMxg9o8w9X/YtT5cNYbbw5Z7mtscfnIG3WNglGbV7E
WS1NlS1a/q+aXGK66lrfCsSbhwGI1nnlCmQXZAFa4UfK3CypobSDFxLtWOJrZV1PMcNBTV16jfq9
E6A7Z3k9CFz1rKHc8VRsVd/ZfWrl9gKjvCnWcxdOqJ/RAAN4yEiWSgECY49ZUAmzhh1JzMkDfmnN
bBIXt4NLHBHQ+8zabr3ADN07caQ/oERrAs3kMPuSRYNNl3TePafbFFAA0WTG8fjCkra8YTzS+VYW
6J0JBphJP0eZm2EWh7PaAr3FS5JmmC7vJ+U7om6aqt30mAwcJGdxT8VooMCtRlRrENIfKlCzzWcB
eJ+TFQYjYeLR6jkXrZCJKRbEkyx7ldpuYOD3aTByALojJdR3hFLxnRltTEcfs+F0K9zZHKWUkNlp
8FCnAhvCTqYdfF0liG39uQvTg3gBf4BBkVOjGgFm4xa+OR4Fa71ta7MmloRLgB/xJVYBdpRVoquG
jmpyR7NnEsU5vas7sIGWS0/D18wes7wh7FQ7QEBKjw/wpwyCGeIhiOZ5NuLjBVbteaJML2zR1g5I
9qQJ/zvcBFIWaLLlHOXvPyvw8iW/RUkVpjiM8e4dcC3NTHesk0dYydPuAJB0jv5RQDy9Cj8uFFan
F03Fpt4VBPgkVa+4yMAypP6UZkKMCm+/1wfkAuYjW5r72tgCWkqzEqzA8nc5qbhtttO6R13g+iLt
8ctDRUZYzM8v63KhgPqY+7mFrKXYxRwEpurnfDonjtksfnAqqMDYcq1+iuiH/zCEo9H7XicaXMro
cceZ+GWM+Npgb1tPy9yWHSNUrRnSBO/Xvx72jEv1A9a8v5zGy5TR/r48Bx9nJoOoJJuyzoYerSUz
5qf5xUvetEffu0ZNqoUHIOCE91NN/3WGj9fZcbG2DNbCF/YqwuEddv5F/drU8F6nLpLEB0QhUWhO
q2SQ+nAsMhbSFVgQcNbDOR0c48IAtSQ+SJ44YXlTUYPfqbCHL20XHbVNsZqReD2AysAC8pLCBi6d
48gPC6M04T9OJ1WX7OOsO1kblyBxwj7by1Pgt7ae3TidtlAee26VyDdkW20ghV41rwHMTI4aUSSl
sc5hUo0169HrM1RYjNV447ZJZd5Vem+lhH+kol720wFopK328ID/OI0CKZhnZaxbSklMVvLqapz+
HlySJncUKzDB75hFlb/Cz5bpyUSULst+2znkioZoZOJW5A+c4Wze345C1+RiSWVVBBLdXf3690ja
DB19V/FdN38tjhQtNXNCwCuJxq3AnNu1zsAah3G4/ywhaLMMOoHzOMxW3ph/OPuC0XViaW1aRIkN
CDWas8hzjeODEQwDHvJKch72y2t4eltgIAFLEmHDaNqM4IwxLYepOE00h05ZoecL9Fjos96+7QHQ
OBUOStQulCEyMmOerB67xG6q/X9vRLGsFeDAqIZhVJXwAdsUekauLcGmZYH9F3ZD+YbbZ+bQ/uRK
PgyXc3vjXSqgcnWxPDmqJ/ZiCoVx8xuO3rEsb3ak+hF/0rud1qmpjzk67At2e8zx8xzykMGmpwFJ
3RJ9I2g1MAwCQ/mIRdKPp8COjexHxOljEHuAYKPYo+6N145hKb3J8PAJ9tOEChXqPe6D+6UfLBIm
tcz0ZiDh4plewq00XvhbwzOkIo6jrBHmDcD6HIo/1RKRF9wsETRud1Ep68Z9aB4BwCe0FG+LnQsr
l5od9nFL4ggnmFaokyEQ6QKEp17Fkpt4j+249yfevMNyG00WQC5faPXjO0cxoyQA4EtqKjBZbSJF
4GUZYSUZBemnXVtekk4RPluxeCmHVWLOk/IMyW80lzhJwbZv3fj8v1xyVNz1LTn26S/KKxcx5ivY
w/Uk7bdBUSRSLtIuqvoYvvOmzN/fOukT7RmIO7TQtmC+mxaNKyG57BDfFX+nwV/3VW4Tl5GJUCmJ
ILeL5apb97mrRpN+rC9/s1V6W2E4bYBTlby1ntTkMSecnqaBi7PJYH2xdtyNgoJt/tYo8tRVyBdZ
SnHbsn2/Ub1crbby30rWh/as7hziPAgIJFMA0T+FrqyAK3N7ONMxFdJRMvukmqN3CFMf248ONb+S
KLiCA9+iKdv9TH2hLCHbpDfZGJTQ9nxJqseiCvunA8ONT/NDl+CHmhNpm95UqtwXuAi5AO23iABX
fkSwhztNq31K9M+jPUlx9rxwJuWOPRIuzNv1bkRV3XOwV4RI16E/8j1cKJJnb+CPf/hA7Nts3uM3
++57RhuPAl1H3gF6GhOykkO2q6di4eI7scHBGkNl1Y1edShQQrDR9+TN5M0/TQa1IJJrvV6pywP0
n8Zza8H3BhvrXS7SR0kOtV3FDLTriwAnWO3Df4v1P78v5gXYOrnykAGv+BRLzL6Me7xh+BUN4AE1
EkgdHGjoa6VKFFs6pF2N/ZEYcwQ90gso15UNQbAJCZtvSrmFQusCmzv/rvN9+ub7WScM7mPoG4d/
Xxv7RTdJwjbQWCjg0FgdhdjIJtYKsnckbYvgdJQSn0udWAW5htqVoojFLfysJVrMUEdeTGLzsze5
mXUgPYor5Yn2y4xlm4lSJp762BNf2OIXrA4GU2PywTswSgsqfdgOeXHFfivE5P/kdBz7wBjV6yEU
c4ZgmGJFJPdA+WgVlzhuImumWSGPHrEG3cWHpaazex1D7Abq7mizMn0xrpZl/wZAWP4iMAlbkuQy
m2H5dLasg23ar6G7BDmXwoCkYtZyKiGHLc2az5Z06DYKfiZK7IRs89hNUma/3H6Z7nQFwc6tg7f9
gmMiK9FM+bSZB44ZJH5PoRrj3XVHYd+mOiHasKk/OsDdzcQp8ork+YDpUGd2s3jO85b1tWsk2LQ8
gCikIWe6+cxFwvgcHNd3wBOVpjPy1pG8jeDkqEp5ZmvMo8bSAmKNDS+89JYoWuGa+cnPnZmXHacQ
zdxesqU6ZktSeYx7Nx9PXJO+q7nrKA8xeJaLFvXvgg8bMGFPhk7HQLd43if3gJDOMnXX+qkKb6pv
VYtmvl1X1qbp7x3Mjhy24Pl0p1mIsptj+7cmiAtV7xKAoCAWTdNS5wAsuQkk//xaXkvpWjb8BfEW
/0vaGG+thYhq9cih2akOR+j8y9fCyyPjy66oaD4BnZhUYYmwGjwY9tdfaWd64oGiNLMO5bDzVyc4
1F8iwlf6f8cdApObYMzNL601H0fOQJ8HGsoLoNwc5pDoY3ZjjmB7+ClUNdY4BUqvoPe7iQ6ut9A3
0S/k0n695rrA5rK/XiD/ZZ/8fDii+coeQ5mC1hMFTNINQNTrHF3+FvZi4HtDJnM0JjFMttMvIXMe
on/zA0eKaxNefiWw//eL2zBQsUH2f9psPXfOiZV6l3DMQ9VySFTMNUJTsmSG7w5iWt1ANLFGa0ZG
oIcVL9WyrMtTJQGb4yxEuvWNPbor/zU+y/67S2pfQim28vzIu5Qy4WNddyHnaMF7RHczQU47PZNC
7gOUXa//edpD/o6rXuCr2wQ+Djv+/Bub0UiZUQSALHg6fumEYmKJyIAYxrr2TGnvzoP2vFiRPAEz
wMMGFeDbHAQbOfACsOy/z2EDidLTmYyTgC6V3UpIOvYmuXOIhSL+7bcIH4j1gxo03Le14xXnuc5k
o0vyhJjvlNn7H8gUleVitQ8lwIOtNi6m1hNuC25QBSJkNW1cj080s7bYInIPjACommZraGXnUhth
aT1PN5E4Y7Ueu88skpblJVWmFroZ7fNOJHQcdg0vr1Oxx0/QM0DzopsWwFwhByGHK3cszPvdTCNG
+8U+Tm54rp7K4R7D51khrvXd5ox6L6KFhHQ5WEk6g4flPTXjFc6vw/hjOb7uqjQJncJmrErcfRhQ
6PwAmFJIQpjWH9Wvvy42ZEDTGdVgVx18uKsf/yv2bbWDsrO/yuOPVHDm67CmXZSkD1CxBK5z5cr8
DWwAsXcrzfECpld4LDf4w/W1DFU/GJlWhb/4YQIfWsC/raPT61ZYu/0YFkKr3KzucsKHpzWVV2Nx
KctRUxf1Ymuwql4JO8qzmNF/GR134vyVhjRVeJR4Wo+A27cDjHY65PmYLK4mKBx3Cd7bg4eE4wNO
kCVyrVP/H/bwpGjIQopokx3cufDrQiFZ+HUJyZH2wtJ1FwEpFxAGXMMXYjc4hriCWoAF5BMKdqE0
ZJFPTKzsSVibhVJWE9kow64D2xIp11HLhTnNFo/hABYwiCHUJi1VyMzN3z1S7sY83l4NvSAKu/o+
qjUxFAryFZNT2v6NC61mtWiJMlLLWBXsRbN6Pz3iDb5IguLu7s066bFsCnUrO/iReZ/9i1Si4rFY
e2cGg4kRhDrtkcZdsD4g8jWevvtnsdVu5CU4fOm685oJcEMVVrDzxbgdrMqySwmNw43Syh9RRDNl
EqVGy6wX6X/7Nyov79+Tsmm2JD71euBKGjPvv8APHtsCLm3UiZJVA6dhSJ4BRIhGjQGO+q85lk38
pB6ml/RFW8MmgilcWbTxNJVIRD9UpebjYJIGcO7mFYdo55tMknuZgVU3ooVbDJyILgih/RqmYXVP
x/7NC7t24oUbWFqNEC9cPkjd0D0sI8M5iyJv0+ABX9mQUAtiL97cVyh0j9vzbbBhLA5dI6j8Pva5
zZldHwhz831QDBRZMbd0taF7Ziuc7gEIZVAzDiDR5xmDFeOK2Z6sBqy6lFaTooNFF+RFyGUAqFrX
F4cPV4sh4loqqZQRlrMCgpgRVteTDDGQlqwYTAaVoSrjbzGWyVRb8xlAp7qMYLV6m3lYpeB865MI
eo//w04zNDn5twfqcT4bTOOpGVAdVBHyYu232y111CoT4zBsA8W552zQ7pKFpxxf0B3/uzKC18x2
C7b/JBLBuN8HJHE9Nf3qdNNdATANhCyKeQ0IAGeu4czYbzPDPTZoSqs5e43KUycuNZtJ6pkKY1MB
on0iZL3+xcpfCV0ymPzF+yq0+gaWGuOx5vssqOyxS2XREHCNm4sC0YIReLu0jYvfugMAwOvEcGHi
81DT0VJAvPvwsdETNduM1vTI1Vk6jqq2SFjqun6mc8OSpZw/y9Q5vBK57ldEL1QU24j2lgYikCA0
hchpgCvuviEohQ02Spo/EMnMtQwr4aP8NrCcGK/mp+1yyZB/jvUzaHAS4/knuc5ORJyRyqswOJt1
kZqKUQ8z1AwzNZerb6/ky2hGNFg7v4p+60CMsLP2h0yIpua1xGw+rUMifIl/HJOBRB70qzUNQlEL
VZrk17BEnXsH4yW/WwDAOmrAHVeTza804FwZWF5ERPR78cdcRFKkM5uExTlKnRcVnkgON0mxq6xv
lSWLcsShwalTK0NpZHqFI8jVxTV43mCsmJxpG+ZoJX6pQmbQu1qFZdwulCDHXJwGnx26hXOhPwS2
FvqvZWWgovwsaZZhBDBCxF8CTpSUXpxn0cpVAIr3J8ISaaB2jtuQUigfKUbMqxz3vRJhE9odK/76
am0YM/m1oLDE8/w6ZYjqFiiFchA8+789gWwvbwPPmfYWj0sjz4xWHBI6ERrNXVRvb3bXKdwEtWnu
ljalJb+n3njwk1fmuKuR0ca4NhCWkoJ+kTkb4FLYChdOGp74mJ3HhdVBbFb/ZNZd03BVVCg42WCT
EMdNJkNMT4O9byRRrIY6U10OevZe4Od0FZRofn7fdk4fJwNzT/IIxMlRFBdNFpSDzmCBHXcuUets
baoG2Yxn7bWtg3YzVcQ5+CvFgDEDUaNnqTL4u/VDDz4T86FHE6gXQOtHHmaxo+okt8qsOxwEm+s8
gi/QPVVAOaQEegQwaYYp3V73qfUPc1EGd1hw9GuoFrdhaPyenuf1jKdx3VUELcQLIEtKKhhP8pnx
YHfknbwAITh0Pu6gTmWHQmoZTwAhWWrZ8VzanGQQZ/0j5bOpJFLUB9P5ZnMMcC2PDGxy41Vxtb0f
hO4QuqhmJToUhkHt1jZaCfjt25YOKX7Ic/qPhoCWhb7VCKKLtiaP/v+p4ylWlUtkQSEPVqdACJXD
mJswlOUbmGMJi82vCjBsxqJOKZpuE9nebUe6TxxW3u0udd4U5b89hL3XUeqQ3RXjQdEOT7SE+Qq+
iIHWhc5jXyGmQea2aJsUgTdWbobgX50r6a8534ArR/K4WRr9aLFal5a7wemOGB6jk3jVoxxpDzsA
wioCanW1A+pS/gD49Jk7faKyzfCi8Y5RR5yiWX1t3bhALrItuq/LbKLCxDQIrhPrzbn4H5npSMpi
bpL++MU0BaapNjbAZT68lyXYCI8GgRpEkDT8ZASrWUctpaAMsvn8YskYXVlfBQ73Uicfet5cjmL7
RAeTSqOhsLl2o2e2TedJzrlJVnLIfWn5l5hgyEGgcMBvRSyfwIKYv64IL1FMOqEAeBi/ab9Vx3kX
EPxOJ8oy0up5zoxsjeRr7i345+M40t8UfoN+/bgkH0+2LvprAne+0+GyppDP0aTjQWAqZ4eKRKTk
6NQ2L9UF/fOzC3Os6GKLlSrlmMsxqPet+B0TET+CB7x4mkxQB4LV8my/XPuw8VoJRK1vAa3Qcg1n
0FqPcsvbMwQMqZyizwvFqlA//80cRnS2jm0awhU1BR7FMoMjJjCPZnxZ+dU2UMs3hDB4XF+DrhVD
gOefG5MwD6p015zjMUpXlf1XeVUSufuLfxOZzlrsnhFv3ZaaV0kZE6lS2oWGfV7zgshhFKVWLtKv
FGX31fat+S2gO2mnPjlsNxwCss/SbHHEeNklEB6NYMx+xRkp9Y+wh7XTsF+Zfftm/bs5RPYw+Lht
MXjcqp7JedE5vLsJYcrzNWyfiQPQLCquBWGq96JPRyEGD7rivGI5bCI+rffz+9OQ5umNOsexYnpZ
ZVc0Tqjms2FQtnOc0X2xazji8SceE5EdPxNR2Um1jtYiPRALycTFvLKyFdPNNE32er4a6iW4zjrP
iayWqn9SW/ftvaq+mXueGNUDfkkft2caG0I3itL7kL3tGqy4dsZhb24Ol+i2UkxG3np+pPn82b9o
rYbVRHh36Eo+xreNoAbcLw1s/65lzSGSpGGL8lDT5pRecaKSts1D85cA/396lVRjxo1SnUayP6Gz
NPI6UxQLdxDgOxIhlXknmmPPvvo6mDFTrL2EL1gJW1l2R+XUJ1FlG2PBX5hDl4ka6JRIcAZtgMsQ
x3V8hiISw1dhHzDrR0RfaOZHDrZ8mbO6ZXTVP8+Ei9x+88k/X2Yq78eKkgkjbtge0wMkjpILeGSu
Kt/SYg0M+NyGuNKV0wTvAFbsfQ+HhHRlke26c9bJ0XapCGZ6pdqIQi5hvVQURifcWQv7PkZZ504P
UHdxWqhvAiH5bMiZu2v5vWqAMqm+i1dkn9lDCdc4/QAhXp39h7cPMqqbmvHHKNOrxT3vTwNU504/
thxyq+mNuTWdeyyWJE3UINcrmqprPpGF9mOG30ejXiyMFpI9C8nKPMdw+Q3bM3wL3s2ldJfTXsIr
Z9idL9+tXfHfClrFIWhh7jTktKaPBR1zLrKKUl7/9TpbR2Qp3aGmInrf3mkytGGqRXwLeLXRsgxZ
u8POw+AuUWHCoae/Ip/5f2YgKoO4hweBM2hKTeLNzcqjeD9TxKAjGbB4d1RK/vYoggl+bRThJ7X8
0P3ZdcHFdxlpyywidxp+d0aO+57CC1T4SOjobYNGRgtAlG0B6IjzcsNUktjkVR0GaH39XEY7lc2s
2V+0CDRNOgFPaxVj74Sb+6dPimZ04RUmwfoyLpqO+w7ie6Z8Bqy6GQw8C3fKouzzN0bx9K8As/n0
BGANToi2CeVA6sCafJwsFSQHyLHsuhYqX/qUKpwH1Q7p6rkVOO0JwxzEMiqnq7MhYM3KykvBIAPh
DbM2SAcBOF07Ia5kJrVNWLrDAJx3SD4N36XOlFlfzqlRBadfddQ2batEmjtr+Wy8tKYD2+QnrSrW
CCVHzXghcd1o2v2q7rpdmIe9VvNT0YCkIbFzXCmotGoUf33Il5UZhjoPQRIdvn+fKW92L1qJgph3
3DBgUuCsEKkIfXpy3flLugFJRoKleSyCN7rpaLHwHbXe2ZAM24wjXRvtA1dr3th9IOaBMVsr7bsz
ieN/Nc0DVwgvMDF4wxtL+2vGc1Sk4zBKGBXRXU4lms4qTP9uM5raQ04BQHVRKpvPWn653cxlZGlb
u2M5AmgmkMvActDtFYN+17J9PW0L7w8eHG2JUDFcWhrcFSIk1AwlCMekCgkBpE1dm/2JOEI3SD5V
PQHU+zIjfttm9LdoLLZFREJ0b1ankhtdLVXKOpsYrfZlwFKmybWhfZmsq6Z4TYk2lVMyMFa7HAAX
87WPiSc7N5FxEoQBG4G3XzJlFugT7vKxya+0gVXosEETGRYHAGpszYWLC9MAXFtwpH7gVEEGW6UG
dB3cQT//6O9fv3fVphIESHJK06B/KubwNewzQx+ttTSJcGQkOv/gp+Bk1aW+9sIC9oYoFPvLdvMV
/+a0acCdaVctPGP1+gaT/VQSir/A+uxxZX/XuDOX+1VpQfEJa51WY0244fBWwAynTA079jQtsHhD
WF1Es8pVzRpe9Lauir8+tJXzEw3Uzsk9t7Ftuw21yRPwrlgzUa63I5BMy3jQGYQKqxVBWLsDyvQP
d5KsIShzLRbGcBKOq7i0MULzPbCOuOPa1aAKje4I1m+ooXGc6khUgJPqWBS8zTWAsqBjzqZxT0wj
LxkSD6PvqllGbdL9EYhOHOeLXybsUiCNYCQ6l+jZTgxfFGTY0tvXe4kuQHTxncE0luUUr4GPPl+r
fjU7PlM1oKajGhASb/d4rY8hivfTrNU8miIoPW9yFSQPQ76jzOY9cg/8kbr7WibXgClbF9Ct6jb/
f75+4nPsoS9+PzQkq+CLflwi6q4wNglkDfKQXs8fMjch71WWqd9n3tIWWbCcW6u+Iw3x/yko+bm/
LePSDQ5K7YMqGPO9fQxg/P3PupyVa5fsfnSN/pAQkUHiV2AasSVAZ+mYFigQkIMsHAWKCobqZOHx
rhigs6+oNK3IWqJYyxO7ZEpz74KkNzL3VWldteoChqeaCN7viXxTNUgfyMlwmOxn79Mujz81dwCT
Q+XhvmQX1sDYWXf6w55U27Ea+Gjl4GZ27ZLUSn5yQU9fC24flPHi+wALJieSAXYmSVdo6EWYJGFw
2dtFFo25+eyBinfE79ErLd0+GuAg4w1w1Ez3TNxznsahDyFtoAkNEBInDKWa3+ahJueFGNUVr8cJ
SrVoEWQ0VxNsWu81NpBYIJj1dbQShwLD30I2yFopLmSvLD2Gml27S+dcfLI1+q1jYB9sRQjZ9LOO
soowB0zjFsY7awMgUhhEGcdSaUVPRbC06ufsL8bRkhk/Knr02X0EfQjSEzxgIhzH5seD3JGZH5ln
kKWI8bAPZWOXQbDxhLEoAvYLgi2+IVXR2FRlMc9Bn55baSCC872Y7rDcoTha9aoLENQOgs3r+glx
wQCxBJRj30DFTOv3Y6/pqujnM+/rfRWdYFVLjBV7yjpAZsDwHiObCE/O51QG8nyFKq/shGGGWEP0
koKBEfpeiI6w5Za/sau/XD80UsCHjtUkXIXzvFYtozB9fRJ+eDm2mnJzgzJ90qIbY1+fK1n/Z0hq
zEEtcIi5HvHsUG1Drmt8mqlQoIuSwSwyA3C5Fa1njqy/+MQTyFB1UjpQYr6vHO0E7kJDZYl1w0Sy
dPA/AAOAkWxcvg0UTJ/a7NZ2z8WB9xEB6+kDww187wjPns3HH+ZnSCP8jC7lRF72Y6TBDUPnxStC
k4GLL12bDPyokUTxN8JramprKNIQh3+Z4cXVFSYpN/5JXDiAeOTnegIWDOIc62bAjxXU98GKs5Vl
F1Vtda35Udj9hdnf2Mfm+UKLtwFqp9wyLJGrnKwwFjh+o+hVaWNetJSkCedtEuVx/F2P9QuEZOZE
6sfYacshXwCMeie/NkBIhAkAenaMggJa7Mgwfa/R1Wb+jIlciVnnOwfcJPyUZlHTR2MJaz5uAjwK
G5//8Um1uz0AlOjhFUlLdzyt0m5QAzWkClHnfCVrrJdMuYmY2B0wJp817hsG2WHrsmBNLYN2pncQ
Jgx+e3fZFaqJHQuP4px8HoToeT7/PlGqovqyqAUUGQiazlIAGWzckbHU5IvTNzcwJc1Wkc0Q/wBJ
+i84CwenZUd59+BPjWnMBUbjTS7HSfG2a+kQGxslmGfooN59KwaZFw7EFPPQvt3UdF/jpdIJfQzE
0GCIxq0HoSKbBR9lek3h8O/idy5jxpRXfV2zDUUZlQnMgBOSiZMU870rBa3hzAWvm7hCjI+ci8Yq
Ie5eEq47FqlUmUYvvHiueP8XuejE0BVLDocEj6LRYBY7JxUQk1vlr9yYr295seCrnKQ8TYYe/8DK
WnzEH45b+HC6H2bvw2WFJ8JLowhF4XZSM7reK4bMI6+chJy2JvlUltUtX7sFIhWGk9Gr8DeUGx3Y
/UVxAVtko1ch1jEXOTQnlJ/KSHOokyAynYypXODa5dCwFIptal2tl4uWgPUqyELU0iFczn25rkSq
7UeFpqXjnToWI9EXMtIc7GrTgdSDEJ9VWs/kVCaOqjjFuoomLZHgp5aocYByzxfTt/HMhRX4wWq3
ZZX/aZs9OWpZp8uPF1DGspjUeF+xlIUtD1Wb6NXxsFvcWF3dN7xHD11rSbpQx+JyqUeCtc2N0FnO
zwVaAxtGs+nDL32j01+EO+P7U9haxFm77uaHSILi8XNcsjtVYG1+iWPElimm8vDWoG87Kctjnt3+
FqswD4GhUKnDwSXqF4Gvj26DF8RpzgIvf4AuqScOvdZOQCyCckKzV1oQAs7paxCGGNNxS8SfsI5k
FZblX7T+BWrIrhl6VsYyDLja5kovEAoxog8k0wDTB0VnXRMYM+rk3Af/4KrgZXwR0YiOHDObRuze
q/EvMFhQMIU9DJeg8j5Du2W4TSkWZaHxn18DIAkriYuX2et3e2CvZE7zppbnCwv/tMntAndZB9Wj
Xl9uaxkgCoOn9YxfRpZrgODdwCE3BdkfDHpfBIXLbB71gKaudmZ6Pu+Yzjs0A5yO08geB2Ax4X2/
I2sS5mAIByIQnSy4Y/7VcEySJ62rEX0AU81IiD+AKcXxHkS1nGhXOjQroip/30GE0EPj0R3koyZR
AQPSvQ6ciFWkNoZVB5rqHQnPmcxAtBJese+WT3RKrJu0ESOobN3iKl5G/UEVkorb7JR6OA393RKH
rjd0N8acLoCkoJUB96obfk3P+2c0p5C4LdJqnu9laB9ZBhpZMOiF9eEDnw85xYMPI95UUpnbOBI5
UJYO1i0CyFGgnlKd/p56JpYcDb+A3QK6vOupQAzSzmQgE0jNF3DlFpj4u5Ml3itY9QfDuT3jDuLD
ERAzlkEBAfT+xWFJRaYWyWWn5CDR0r78XqL9jVobhAJKpxuqGkMy0veCLYmueYxyH0wBZrQIhpWE
xe5f1LgtagDVeToBLCD1j3jrgjWboDHLAhOxp9+6ZcFOLauJaWV+hUzIsbExNKvOWqYJNepho7FF
7SXbD3KJ93W6xA8v6sGPH1/Y1jJHIyQw4Dc800fDgGykCSkykXKgqJ1/8UV0muZsDVfKBFIvFPtd
T1tW7nIdU7x0++UNcQG/Po43t6qletA76VGUVHCShkTv67h98JqGItUFPJ7IwSdpbOZjqkDEmWmi
IbZb4ethDf0TShmc0T9KBP5s+wDkPVscQDfGIxQkktpAFgkhvj2PRuUqK56xA2ISAe3DVPEgTGTU
ku1BEPNYNYHG+FxANSn+W8roS+j8H8z6Y2XPosvRyzHMtC8JXt/6MX3iYYGl4sacW4upuCFC1h5U
Y2pOXHak0hqsLPDqj80YM740dGUsxoJaP9NZEHSrIvmoYlFa2/DLIZjxUJviil2BJ4YA3W8TxLbG
ajyGlBvEXh1DtcB+CHaGIzHGjOmiiyZ7K+YtJmE71BjyW826HZMkOGpsbE8fTJ0TrKAWuTKMSjcY
SrS743qRXhjvTy+GNY4rWn9P2a4C6wO3/Y0gWnciHi2GRJA2zTxlFp3VES/Cb/eObAZ5+8P/KotK
UhYL0nMwM05sJRXtb46jyOHlWk3otKPcfckEEYQtFbVThqjP2+ge0f6+P1Wz713Xurco8OOx5ab/
ZbUJf9jeUQr94A9cvsUxLQT8YMwLIDDUsCeXYXl/nzUdtQsGwOHCmgDVg426Kg1b4A2gLjpcKKeE
m8hla11FsRIN4bD3m2w0DMqhZmkJU0DsJ7kvcAcJklik9lWiRhkHdPrJUFLnufFGSBubPNJyvANE
DWnmYQGbWIgmmgaI6iJw30i6eZvfGeK0pKBDJii/R4jMOk0rieEwPhpSKiaGKlSylfSOEyLO9wPv
RsceEs2RrhjjErzCJk82Tjmgn51ALlCX3/bJOzgWjMjENOB83F6hRmewJ6BsvACFWPyZOJnbO4Ey
fo8Lyw+g6P2O1dFyd1d26G8n586vII81CsxXHTlQe1crm/yd2UJOizEPi8dmt84noYMoze3bQqQ0
bh6JryBaTcFq8xpDqZNWsXJulMBVVlnWZXbQN9kDq1vR8GNa0A9bdG1t4lawZlk4yhwvymHF53NB
Cg0gjC6zlvI/bPjNPrHaVZLqaEqYfsiN22NmrtQC/78Zvi6NBvOEOlkBY0u+EZIcbB2DNTzkvd1m
MI9EeOEgR9WrknMuFpHARijR1mCNaFx6aPv5/50TrIePzneiBBYfkrN+GaTrMHAsowBnUxDDkSjm
aH0g2IOmnQbBVUyqXM+70G1e9JfJfCk8GwzOXSriJJ0KECkXIzu7MfDYV9Kmg30/MYYkA6eBDv0q
pZQHGRxawHs1ml1uPafhZeVTSzMJq8un+Mn+rQeBJJ2tA7NJCMiOp/MiC6N4oiS/DBMAMM3mjorU
EbOsp1cUDIT51m0Wv3e9+g/q8tL/UeDgTgSS1PWwQxg8KzLuwKoHI08Fk75a9KyMLbc3SM39oa7B
Mn98qMRgV2KD4mgkraIRjf+dbyAtCNtGYZnF9ED9Ri+CIDkVy1u9rGSNk5Aq9JIaXJV+0UQDUXRT
pfqDSLh3phUs64ViMlFa2fOgJap6nnuoZhl+5cXUvVpoheQD5IYsH2Ig3ScRmVkCcVjiDZJYABqY
GBLvBERHPqVVfUJp7lUa6vvlQ2VV8T5CBRMs15SdxtKukk3WQRrQwu5SaledA+dulOFATDyWaji6
Rk62sNiwzuZ1GZbaj4WExO0s0pCXacEGqYT5c0dWWXH7NttxKWhedUCvEZfVhmUyKu5ypLw3X1Ra
1gIv90efEiE9MIsUNM3nwikQ+E2eYXRcD/0TKdYSZf8iSHnIuNqyWdK5fpJ1A/C4DDeJTIw+yvZv
du2I4W82r+DhqDmVtzfXVWjRs4Np2LAZjI0niWSxM0owT70i1syuKgDcBuIeMrrUL0QEvrpIwQAR
QTNuCwcQofpTzMAaRATYAX8bl7+TR+M3GgcKF4XA2GFRxEROB17wvvuOb1a19i5PKdFJ3llR87BU
jNLSM+aePXIeYZNs6eVtT5MP4m+UulmN9dEKlMck2Kkg6IAQwjHZ9+RlQmDlj+MCQ/awLWG99Cdd
otD2nW8r4WznsmtTzumfNPsduQIFZtz6Azrnv0/Tn/aE77Y+wyAZ0DA2ko1RuaHXT0HKFxbYvMBy
wTZZ+AGVxbY9s0z/uXW8AGTRHxvspIGm22L/GPj7+OrUJfP3CbCkO9nidDFmPU3j+aGfEIoEGbPc
MzVML+Vji/V2/4KszLs7xt8N6y3cioTHBfZ8wL76VK0oO9VNqeWpfv1KvRk3t3b0VpmK0AUU7dbm
fA7aTxVnoA7fgG1tiX7gzdGN9G1bYgySg0wumHjO5soEqThUIz1ZuDLzrLCcgjh8aOic5j2zjA1h
rZf4YdqRr5+3hB/kNP11Sk7JQ/M/56OKf7V1Vz1Ij51/S0fxRwOJwJYY55WJy5PMs3qfnC32r0kn
ZSIDOjKsU/aeRFTmAypiTDc8V92f8Y3kNTxd0a+7V+j79JMtwWP977gzw6MpzOqniRlV42LeDZyI
c7RXGqUVUH1Ws655k6vaOZCKj5CKFdn7OTuMm4KaBn5X2oPLtoUB/jWbCZGVk4i+50b3+w/qs5s5
9lR91wJJoT/FsQPPPtk36IUinQKP1aWugLmYtCf9me2ZgtZskaoGzj1UjmxwdJeJ6aGM1Edgx4cE
J5Ex5DzwHp/Cf4QPiXDLnf4fn1gu89DdZ+WS8+jwtEhOdIFpnXOw3lxAWd2VKVN/d+QcETQqRUoh
PzHxrSqs3UzzbjyDIcWblOzAkG1kv5Y5LhSAD8QtDQWbP7iu/bMsMDhkQyzcgErJCCfWOw7h43Hl
DfCD/Pgcx+yEP6y3/R5JYEk3tiGXgL19eFEVRGpKiheOt/K/L+feF0Ftno0enIiMnScucHJgf2Xq
cUden1srRCmQ/ysVZ1RYOAFzBrbNJAPUZteQmDh3hblSoF/3q235YjmAizW+gNMnzRN8IPZIuplE
49MFvpTlMk9FaHauw5vwe8qI4SDTqxZ0LGf+6v9Ku4KtsRUxofFUbF3enAml0kQ3ocq+MbCwBE0A
MdDWtq1WpOMHR9Aqm3WuCiA0PCjnh1QBD1p8KsULniEkKRr7dfTkjWVnsbtva7eZU1ErHRH2qCy+
XHnIhVrU9sukp2BfYr7OSRVw4DE12mjOmZIntjYbsQGQeHgK0VQ/V7kvQceYkv0XwGDrHy5vEAmN
ulenpkbnB0XC1/W0JCUlXKcoOk5TSRqs3xLYrIfbBEiqPwefflfDcHHe22iG2W6g1HVCwJTSDMNI
cJT3w9PwVog2KMBvsNXCJOTWjL4K02hIVzI1D5oMd5NqrsZiGgpoRBiXjNlcYW85xyUqdbwejVbL
Tj1mLtgrItpnAz0gHnzhXXy7+UeFT8RpdWguzcyenUyisIzdMZt/elNVF8VnljlrJa3+t4yqRXc7
77uz0uXVmjYq4ojI5SoQ1+RCSTYc5UlSp4KKbztW4u05BhWp/aMPbpzzaTKXYBXx7J2/lvWwEhc0
AaxcNb/k029vQdftG1RB3XkNIbJy/btVDv1hA+zlzISVSFwG71zsgR+I1w2qlP7vsppobJldQ+f+
TWg+GpHiNEbGBMmSoiArwJjpAYe6xtO/LaxWyPjdsSKte/+iT2PkuwO4vKM5vbcM/GVfft75Btc4
69loG49hze6o7M5g9Y0X13oExaWkgIsIiAM0bfAU7JyoBK6xGwVJqqLQ8lGFU3v2Kx/Bdl8QkQY5
lULjTMOpy+CMvACGr40cXiMn87cvpn4iujBQdXaKE7uiuz+uqjl9gEQc3EKAYq7NWX0DjIt0H88e
v1IXyFgtQsM734sL6Aq1nl90xm7Evzfxj8VhOnnN72HiW3PYHqmUn5FZbFiUX6ApFsa75r/bnbCz
H3j19qtABEGXSHLip36HL4WR9PnLb/WrDneAYBPC3d2TCLKN9uNlRa6aXw/Tqg6lS776rcBVOFrt
a9BoXyg/y5DviGKTVm+P+fUWkIsD3udupkh2teBpAWhL2QtoNLy8F8BHwiecNlE+ufQszKtG/RVM
r14EdAoavVappJbtnV2wlVISFF9qCraYXPc9kDa/aejxV6KwWXwtEO53TFeJJmhDSKr2/rMepRTJ
RWgqxyNlV+SAVQ4qF1aYDlpSU3sYxV2BgGjqie8GfIdO93F92vJv0LAGSBTEsSsnB0FzSNsrd9fA
mB+SjXTPAz0YUIVKdERkLFVKlguafi0J33Z/gmZ+OP1KZQsqL+u7Mjzp7Z4w5zr7IMJr2MhXEjJB
HysRWhudz3k5mZ5LoR4D81t/J2eh5zz16CBs43XgcC8yRDtq9NuS8vd/fdzDzdxqr0P4rvsHoFDK
jfdRdmhWT4rL2zUXCjBkX4wYBycrCBctaAQ9pBIsCWaOJO3in+I576qV1BlsJ0KIHWBTvU/4ftPH
nBGvIcLXdc1oxYcAO67m/lHwnCMbull+OQpLLXVYq/ifnhyEQ2WILHq1MdtXhCOi6V3mRp3wXyrX
/BWTYdxkNygaZUtYGISwrcuAeVldRFloC1ZrYii566Zwi6SI9SI2O5n2NV1QvY1eT3VcU+HxnLvm
Zbmo6GfwT7EVK7CYAcPmgpDX9aYR0RO2W7miSfqQrxbn3EDNliH52SFG5UqHToh9cjv2LcSnKaJQ
iW3+JA77XIgOSXMPhl7jCCPWUcmdCaVqwT3yDz5MKNXrpgF84Wi55QHpJ157MlhA18mO9THdrKNK
sQOhQXacY0zGoCL8MMTQL3T0D0El+zgqBirlP0aEwGFXXymkx6ItIA942gjZZcW5UOwHiNmgVyCu
zaMp+85ckqhUncQkxfQZPDRdso62RMQmUl0ABD6BRn0PQtrucj+NkmEetaLDLSwzDv9SATAoU4L6
r9I0hENchUGmyzlOovJHEnoeE0FlgH8kT2860nBRMO9qvo11HMeFFeC8Y/AvlODbg8UemZ5dcbrg
PCfQMAB5VBaBklrdK76ef4C+RqzO8XCkvUw5uotkJ/MF/bwQXDsdR61p76IEgGGtC+X5KaWVYIW5
NcDQw6V7q5ZuMyDP0nZHHwKNJB0wd36X9rw6gtEUgTl1HaClNuEcMWI/nviBoO8+U+YhpNRPL+F/
dKXpPb047jMT/qQtTYpLi5zZCLtbY2yAXlUv2CliBghhclMThrDZlX13FOaf9VF4cjHvdFQNRRVy
S5tuF9z+0uvAhpgyFiFRIYG+MV68ZxIfK5V1mBYYdOhPlaVKl+sj+cWbxeFdCwMNM7hV757pL0Ct
w/PHPT9a+M2WDSlxhbcYeDZW/PlIs3ztWw+w3NALBMf1fdgnvbDmHl23dM8rnL0jdj4rFtMQPIUQ
jSGWxMODyvmpEUANIQn8iorLftfhejd8rLcbvQJYzMm5syGTfh1lxRDDOgW3Yc7pvJRxhrC2Lr1o
qBJSTd432wninVJPNfnIxw705X0zzKrZ7KYg0w6wXURmVdy+3VUKX0adu/pSooDwfZa4SPkh4/FC
4K7x7yyTvYLuAu1vvEDlm0r8i3Xr2f1wWjkRxtbSU5nlHHrizCzNjG64YfXNai5NtBPKRx2qPxwm
xMqvNJlsQWGlxsh87LwLEWLi3yvcmqvzlC3S/fveGuf5QXSYXMBRoRGz4XAqgBJsyPbA14hguTxc
3Te3coY8lrG1cayNChymWStfGoqeo0UgWCdudOZho91LGh4aJpT/DbKEue3GHZnLh32cMEHevJO0
2LzcmyTCI00le0o4f6RiLFblZt9VcawUv1iMwkOcP+TygyPOxTY9syGJT6V3DDMYeO6UHy3tzIro
w9XQUHfwJK6oe42X56VKpyHDZ17EHzqr9tL9ocf40cOiL5QkHKRtYA5mAyHNHpWIRJynMsVs/YUK
zs5G6yA78GZu+Hhdi2U3PZ7Kfy/AvL1ypVtRJ2ir/CN6GQZKFnzwcBhlKgtXmzyrSSMETwMVLzfm
fjTQRWPQsEgxpXQsUQfe4UTT4vJ2wAzE2kvIqqmOAx/SkaWdQz59fuZcsUh42pB9+q/oIMYOvIY6
EzlzAehWmq6fjJcnGl0WhSOXV4mA16a6u8ftvf3iyx0ZNrIn8GruCQaYLFPvYBrcQur6+goFVo7O
KymR/srlFUYtOykEzidBF+W2vySn9fcPsFoJwLs3aNtVZZ6e5d8y836EiwqO24JpCUSgXv3SnXx/
PGSP7Ap/bO3jX5SMafKaHb1ExANOOKelLj5Lfc3HWr3/o+UEVGuxfV8hsyYbJW+IjyMDE+93YlL5
xmGowaVwCQWVY7FHp6PvS59vdNdJ/CECbEQd7ZZfV+rYfJvMpv21Hg7Spq0LzgIdigei2sA+jQz3
3rq3BQwRS72EHSR5DNAmTeHw7kcYVDzn8UY85cFrguyTV+kPTfaD0g3zaBCja24/pK+4118ke5fR
MiMK0nYwHs51X/NM6jmS5siVlNhRzGWfR0mQ66alUdS3xaUm3d/FWs5y8OmHfWYiAriWyeGCF3K8
kG2DQ5pCqD7yducavkRttYdPk68KBUl0qcpUDF57d8pdytXrfd7IASyvjO9ymgjS2h60PwSJXWqx
JT89UjgKARbStzGziKHdO0CvdSvSV8jSKKcn82Rf9MxskQVd+Zi5ul8zzfWJ1MQlmRyZFjME+14h
X+oTIFTX1jmLuSLZik9N8lSQvJpuA3Hre3cLIDK381/PveRrMqxyMDdL5cy0tF2Mh3aPMtwJdPlm
CM7Uxg81j2cufVq/VVq6vLSF+OY17vnbGStz/dcMmzGSzIDetMcCBX0Pb8uw7d67XkG4L+YZkLmy
9j7HMCXemZrXlngY7kfJaoefSKLY8PvUiFBjWGjKIIoghCCsJ0TgpuJ5Hx6Gdx6WuXnZqofIeaob
Oc7rX0LDKiFQor1gCocdteptNx51UmXyGCDhtYFgzzrrbag+3W6l79/rbh3zAx3Lmu57Im0oQr6o
ukMT+a57SPg8j4bRa0v0JlUVSHyxN17ZJAycBSLv1uwKmsiJ7TgXRAxzs4ML4zBnI7xs1QpGqA/w
g769umKgdX8MSRGTJhTTQ003A+476+JGljyeMBGZYJfXa2TWJIKhZIOIMmXpCnrVwt8XOqDNHugr
jZyVcUS+U2ucU/IqT9Ds9jxAVgKof7a/c1MEkG0lUS4WsD3A0biJcKCfoFFX/Q3KmBwCEoxs4CWN
0/9+miVBGCSSrcst2W2W6SOkOcu5T4VUVCyJ1chS3uO183AhFZRHAr/dcMSreD6GpMj4s+AD/tqy
20SrwC/R5Jq+29jZGdrL+kCli11GsWNZObqND6MZBA3JUAL+PKwyTv+DFTMJjLIGhM5SNrk3Sbhh
FQbJjy/d2ha0clkPiGy+XqiXlsx+XjHMqb3JXAS9KETbke3d6AKTJ36WOkJvo4ZUovVfUuS5g2x6
cYmUq0Jpm6pWVCCFKhuL8bYsRBlFGJMedchlyidVLZ+Z9q3N5vRnpt/gnpXlQlXxe8s9E4Qqvpnm
Fiw7wqWOzlPewxw3RB82FyZ/jwNLRwq6c6XWlsESuHliZ5ib3ifB6P4zY9DkNnaMLOfcFYoS2PDc
88s3aHpel3SvDpYsomvd49APhix9Prr1utPlEVYNYVBftjDXyEmTJjlsP7t/ptEsreLFBnJnjfnP
6q19YwofHCmhLkeBSIrfHGQwVexJX5Loq6QGg1uMs4aUhIxdqWnFWZu67SQE/UuaZiy8IxBy8zv/
qgL/OkOqUjMLiJHavRQkTQR45kanqn1C8O38AuIgXJ3yfTIcb+IdwEdwvydj3TmWgyNbiZsXQiFK
Ei4/6uRGRICLrvdI0xsQ9O/46zvQdYKttQB0rDiqFUjQ6f005Cm+yjp1EUe/St5JgiKVj4/SkYlH
glLV2YtYrpPB6nv9lq+kYZMAd+utE3TIOMpFkZGHoF93Gi2UHgTIwzT3R3rZyOszMk2XBodW0FTU
1cllkdolFCf+auGZ7kRMb/Q2vdYLs2usOcD/UZuE+yX0sZ3h/LGinOEfXV10hqiGhjqvirl5q4Id
2PhuHur+2ihMEH5wEND4QIE4Pi5PO90+5gQZISESKm6I7F18I4cZQt/PiID/qgIab8LcGJTnVkNd
TXyl0mVKQ3MYzKrXyzLNO/e4rwnvzf+4oS2Trv7mf59mUj3OGV7fgWvW0oZYrtOLkQzxm7+Hs/Qh
XYdQXKk1cfhtL8R36q7+uRhpA3hAPvkSAMAvieCE1yQk4AiTzgf66ovhxXcwGjAf4/Ri2HMTqW1t
7ksODJcj2TDUywjZO6Ravbf8Vo/m91xaK3JPBaKTsCm0JHA3ed13mjI1ey8c5F4U00mTWSgI99mK
joOFZbJD0DRCfVab6jctxUf7dNe+KuhrLgqirNV6m6e/ATSrDEtaDU3tD57DfW6obIef9uVe06p5
BP4uZ2l2x7nZio33g3sqREOWbeRRG+jrhfKTWeXJaLVMbAmq1m/jznh3UGVBcea473rWc7jQykat
gcazG1IeCh5C2gZUnN3kmDtnml26t8HLGCDDbeXegGNN7+ONm0ZycCxL+e8YoCapR1v748wn0/6A
VlyYVw/gJP5z9XS7KdtCIvP45inE4Zj/exsUGAeOqMStZgscboXz5adi2SHfPmBUTDUS1bEowwy7
b98Sk2CKVi+SghTm4uY1BSJgVQWEvFEfpptF+zCRFiNwsrWhuDEpz2dchbfgVxv7RxH0VgdG566o
NXBnzA9L+qtlTvJopqjEWRmUylQ7qFJCD6UTrTnA4XFM0VozV4Z5cBpGh+2QPUmhmR/beea0QelX
+jdv6OJ8BC7JVFsgclkeJRFCmyyr+JArMnDqeTzFa9kqj57kAueMS4571Hv02O+Ap0PQmmDRUIjP
eR2PnMLfdllnRewVdBvMH0oqJb0tZxBaLvnCQXwAI5FtIduGgjwcNI8RMm4Fz7dR7D8k8C52jUil
8MDCwh/CHfDWwFD5k3DlWTdplnkFFRXuO+QgUtPVtUMwgRuzGFlrLeFfVk9wA3uiEfQDRtdmN9y6
0F5GUNUCM8X03BIuHJJAi9w2QjwbL78CI0b9Qd0lq2EApDwLBhYwNmbh/KkF/GanVANs/VaFfGqv
2QqDej7OyLSNIveCJtSRn9M2WRClYAC6Dt3lW7sxChm46wx4Y+I/dtf/bBC0tqxOX0lXAi2vr8MP
ssJOF0kEOyBInvjfLkJPxTUqYfix70QRA9W0uz1Ftuxlzxiezw5ewNPd6W5Eg5CmEjsyIHzhc3ux
bFGrYc1QDP8E9665fA4Xn5kqyAttP7tQ2Ej9xDieihIf7tWFdpGpiBYQYW42VTeKnsk992n7NZqG
50NJdq0gbF7tZebbp8Z9OA9tH18o/0i2APtStQ9MH9nz6Zvu7QCehghH7RTv4AkObuoEkjHSeci+
EvMPkvC7gPkjdm/bmidf5F8Z6Fj+ERnNaNTkPGPhoSlhSBYcuprtQo0WbSGz+RASgEi0UCFufKO6
GV2yokiVYpxkRaREg1zie1F8Weg+xzs3P69ALViOGbYznmWfogrQjkbzioYaIvq/PBHa20DfPo+y
qDOWR66QiGzFZaodRfykJRbEKqqXgcLqQlSGHn1AvwjJJ4TgK7fQeoHWhJiUxTTwajBsJsoKPeUZ
gLh8rCHjmT8+hdfEQ1KGpznFR9inzuGvU1UnRt9LVPX4TXf8KG1UW5TTDkY71gaPdLuAzKagoVee
sdZ2xkP1PRhkjwFg0bmoss1ll85DfIcvnvS+j9qx645sFyAZk1fi13LymgOABRj7+77Bh091mapv
yj8VAU994S4oLanUi1Gvh3X7Mn2+geaFDip7o0IIGxg3KffXBFhO1J4yX7qsuekRyl1nM1gp37oQ
CuSZlp5uP73Tk+ly4G1ZYAdf2Yz6aE35WTI6/rfIU8wNdEImmaFc/UU6uAGck9YHUR3mIW2IgF7f
djZCbCZdEKf23gXJBrLqQ3a+31uQNb5JyBieuliVr9MDpa2kiLjcA1+oXXtiRX8wxlgBsVCOOq8a
II2vsMbM1bXtdRI/GEw9qQUR2m3WsaD/415uYAATG8CeSinnx4+kSSoWl2T1Nw7hNAVLHScxFycI
Nvnhcg1gs9Lp7SZaB2zR4gsow0ks6X+IdD4/bZ/7vwvukaRjlNeGYVTBCLSV1LfMqMXSJzGU57aH
rpcL26CGiuAHVY642ERmyI6wjPEB2vrqk8UBFWvoJV5pPgbkqAgXM9YyH0Ywqg90BYJfPuX6m7cI
tuprhVW30YTnFPU6ypGFB9QH7XxtbYVHU1d1p1QZUaed8NhUySuSm6IAizElDNXqAve3oGZH3R8/
Ihnwmp6HiUMXhGqLmhPhLlXjzSnYC1eW4OKWwVdgHfi7z4JLkyQJQzURPBUC2PQNuumo/Y3t9b/t
oqPxIweA75WMcqIbC/UG1wQL1ac5+tFnnGpQ1FGp8Bb2GLFb9L8Lm2cbtLryAcaraXJAthBjG/jY
xdbIlR8IyuS6NgbwbINwUHFGnnlRWgNOw2XS+kkOHXK5U6uQodpXcW09FNNYiA5pIEmDBeYzxZ1Z
GvNs0wKbsHlfEweo5CUPTwIUGqTJ0SCvzvFV4m2bx8+tIgM0gsYZR5YNJ1CrTiTEiCfbeg2UFomk
bbkZ0AcVbclbAK4fyvv406NlqfgBK5yMgjsPoBKuLAPU5wD/bVw/foosrzA1lXzgyaQ46zw1hhiU
NIKnQ8RLxMiAPgDCRqR1igCRpe2IAN+WP+a9zy3oQUsws5WZzwyZXCRkzyNfO2mmSf4dUGkhsSS/
WVzaHneOPRHu0QIJFVx0K3bJOnDLu2wYIuepLfoshhhx0lUZe9WMY4bHHixzVi2CiiYSkpLSHbUd
KIoUmdt4Ni8aHgSlvZeUv9Os6UOitC57czqLn5a8y6VH4VKK2PLH3bESnEZINqPeg4AfM1Air4+a
FDZt8SGtlDfTIoPZSC0BlKkQ0i6AOoaAN2bfezoZfoNV6QUEm8eWTCIg5WVbRGE729IscpTee5oS
3kbZwH6yAQKZpU1AftaU2ktIscfsAYWyB36MhCUZgpT2dLe5rhV84RZzToNpx6XoNeUrBWxGEB1T
1SYOQq3rmIWRojn/TGjeCGf1LUBAPm9TFEVdjDqGjnGS/V3NgzX5LjtKqqLjK0I9jZqW5QyvEYz+
lFwMGoKcrfY5SEGSvN09MtFoNmZNd46PxvIlcdi4T2gH6ead805LbQlziFXnsH+AesnMWcypIEM3
IFreNBJGucKzhNxRM8hxW8k5ZiXpwX+GvmhWqrPr7DGPxu8ss9zfQR67negc/jnNzuC6pW0c0SFb
6aC92IxeVrFtgUwBdB9E9QNYyOk9RumgdwLMaB1eU6ExR+VMDRm4zycTIeN9HCQkOfmdNW/j6GwU
aA/VmpMRb4zj73mD2rECQV2OzE3SVlmzRUXhsyKMqk+i8Z2UVVuGmH2zERax/xHm0EnkLIMhWwGX
cWQ7gOYo/SqdB04Ny0Xf3S+zwXEDRlym/lQzkUUzmVEMQtDlnLqHJH8rFJ5dsdHEtNberLyJ+Q4v
qh4LJyzLybT15Ce5qfD+Y/nlhAUFTCXP96cz4V4kiWiOj1wWkGIkX2hv0wKLYaFwodElvviB2ZEM
tNseL/i1kEFaRg+kyjd7bxRvxJZDZSU72kT8TelFJeO0FCBtPAxH9U6c27xIVFdFMSLG4s3vWxiM
YIovD8fzEkYBvj+UBTQN/q1nFzoJekU1gF+AS2I2ZbYWB8lzw5ZB/PryMvAoW8jRpgX2HGsvMhhy
d/bcSLbMjgg/QT4RFryaXQgpBSh/TtrFZ/jNkS4dE9iy0iYWH5W9q0HadnIRYZWc5MhjCAORmf2R
4nVsc9yjO7fT34gc2Cr15jLzWqHCpAajRH5lls+hoYNrj723yCTYYXmD1vB0aiPmHeLgTTYqWEHv
1jFHI56bSYOMGctD39ZBXF+3KPjAX2OCapjHIJXiLnIMF3OTl5OMo2KAOSQCN69GfRRWjV30mijG
4ejM53JCaUk5e7CDrSoDgaN2jLbbFaNjZGPn36Pnht4XbTahCfFqt5D850Vg3HvuKvptuIvKynLX
+sxtQZmo24FxGnjVKLYrZR0wfKEULZld3U3rlu6QWZ+TqyA8GY6sGYmwN46uT03x1EI+KQ12g3R/
qKJetiY3vvfyYUbZ+Np7Ca07xw/YcYAPrP8ZX1YxE3j0e1YIMHmEI3yC4WLmjUQ5xW0oeIMq2gQE
24RQev2Xxq/2TWc5m0azGLCDotwBlTdCucCo2iHYZySo9meodTD5dfp2gh6wPxw9cJIX8duYin8F
c4qWR1y5YVxlk0GcS1ru680C53UmCuVrMwuaYo6snoRKH6ED6t0741fxVEaoxnZCE3vhNDeD2L4E
X3EDjwZTXT2cohu0Ezu28BSR/Jprl1ubw9hbNxo+chUu5LUKicEUdG2rwIg2GFbE0n/aqxwIKacJ
j7i4G/ke3YjIHk8/C+LPAcYFTriqaBg2gXH/Uinzv4q1WXsXhA3kbMk9t67FHL+Ermlj//rvGlkm
sMIX7x3db72c7nK8C1XiYScuwkP6ngv6rP2ZVvpWsmdMtVb28wAG1PmSYR/3xhu5eaNU8UY5G8Re
9owNe2dHqH/rhBOYORvup6gO8N7hzHLOlDrBExYVQwmuj640Z11gc8rkct+qMIVglcrRXTAIVznx
LdW9vqNRQRuzYnHu1fnnuSXn8iuAjz7bzn3iu9Cu+iJghsv/zca5kVM94993Lhq0keAYG9PkocYm
n1+k033/Xz4pBERSXBaIwpQqoTwI8PeHgwPfcn7Svr1dDRQ2X8qSLPgTIUyGol4ic/f7FbUY3867
klEZIyzxpbXdGcg/dAB792jD1855HjFy3OtQ4y7fhfWbKSLCid7FLXFLgmzyCSnMyMZ/Fkr7FbfZ
hQce8WxRkI5KZ8ppBPdAnETmN39G5qxEkPuCVN0FH4F3rxlgHSWNWV1G2js3re00JEo5SLIXiVGZ
m0xHfysiDMYNXHfHqZoeU/1FzjBoO0wtnK2Hmm5/ZJRuSg050RQaPfSb7+IPV+lUdISJiYsGy9yM
bqBHzhJ5PJyd2zr2YT6eTJdBbu41Y0v63CflEy68j47vfQAONA40X59T2+HBNYeLYEy8U2Z5nyrf
Ey/Bckin6NXpBkcGzLX48oRHSI7OJPYQLPXUtJYPd9q/S0i2C8ewUpIZ8acwvCp4QKjR5uHWy2Fc
druQr3idJpl6+tuqHTFB2wALfJ3GOVJ9fRlcSgB5quPFJA+crl1lwxoTb8UGGAZdzmQhogqXFaNe
s9EL3N7gTvmS64GvpOegAXMix0Dswk/cKoFZ0CnnppunJ9ZueaiGk8UyY+MwQShvrLuf6GW8gZTa
9wF8R4DXc2nLhuSw91ElM6c5aAVxlZTbqZnxWu/+46/viuYITlesNV2hptbSC3LgUPx0CMyMnHLy
2KbLONANURg8cARywLWKrHiYs76BNNGGYNb0lrSztJZdixGSI16mtgek/iVhGQsBdenBWNHZArv2
TXhS0FqbXOrSGwNxt+qPWTV5s+ItupKzM08HjWLoPNGlahxMU2TKiCItl/FkYiJ0Y9XyCVAv1lm3
Hw/mbZwc6wvfC2EVkp6C+SeGGQC3+IeyGgt89HzbYLWVakiJkFkxoU2AUt2/osRL3l500GLdXz1k
hoY2fBiSvefEEgbwLkuk3aarkcDCfLW8Wz1aG72EMpOjzypQglngh/+jWBVqN/sx5MNZ0lr6mPK7
/Cr0M3wNHNy5m9WamTepDxFJNkJwLOj9OkYq2DUXUU7jNypr+JgdTa64wd+sHIQyuNd9lDMqorZL
tu3yTi31V5/wu9rIkcMTOFTstdUt0P9nVChQFJK7Cp6fO8t8gl1N6CzjFdNdoQqGHHxB1jHKhi7t
h5VhwROmTV7K9rv0b2FXXAAM1eBBenDm/W0xnlHtEwOWwIGE2qwk3k3ZRDP6LpV+N1FIgIeUYYpf
NfUAntEpQEQRH3dTRxJDvo8Mye2yzeHoKOwqnCN3cI9QJ6bKX64n6CysQsqNpxKAn+imExOcubbP
X7GFa4S5/9BFKS/O/vqHey1Q8RFzL6cTNC7JAzRUCv6PZGmD4e/7/Ps/opZCs8cR4QfvXMPFK4FB
X9GGDqiwghIk2U82J9BbJZ+vURcYIaGlCcGdggh8QNmptIIwud7V6WmZxqdVwtw2XKj5RC2HnKA8
ebEViBxeOH7Fyt9sKNVPdWYksgf8/RPQP0cUq3Hk9z+wlvWunnQ3sjj6sAVu2fEHdFu5xIl3Q0JR
4je3l39cNlcgm+fzuI1iijkFFwxyh5vhy4z4qV5pfqKY6zKxudXjXeMatgujlbwrm2xNinQkaKrv
d9WIw1b6fqcfC7lcJZBCmR3mvGDorOxQ1WAyIgU7SXuk225vg0QJzBauanldjZV4Iajp469k7bC6
K4wg+fgm6a2PFjUmGDiVZrhwIYPhDZOwn4oHUCjLYWQlv3kpVy0vaEPZtHDBO49cEk3uZZe7Xk8G
w9G2VTahFNcF2UGgRZRZsYQSS1V5Ncyj6i6S/4In7akzoVbgZw/8zFxaoI4PAyWBoOIip3mNtZ5M
eqOfMRBeJB1HgN77fNGtxwf4DA5cFlPqc0snrghfumfXh+BulwkAScZ0uvJP+2+FpZU8tsuRn1uP
H8lAGach/LZhPdOjtLRl141VqhfTNoWhhiA2+dfzqBbesrIBLGQHxwMUm+U8yjNGopHqJJariIwK
qe9bTpL1jmmweNzIC21RigDSWpJS/ve0G+DsDOou7D2YEcXxxf8yILKbGaQgj7kEkthYBJF2dAO6
Hryn6U1J3R/BC9IfVa6giOI1HcEwHfMY/67faBYW6++siY/9hq9IkkeWTP065FmECV/FjRseYoTj
I8jzBh0NlCfqv7LuZvthQantSrPSHSkm6I3VyW9mvdWCHJZquET61KE2bRubepJOMcAqpcu6l7sT
+532D/vyNRNkTi61YzrbwzhcHThRIbVb8695rHIHCkq7RBmDiaHPn9nx8+ZbNttpED4FSFxBmc1S
va2H9CinlfGAnZEHe+Nt9oXSUgwMYlmce6RES4KmXyjrxpFRJZP97CjMNMHUWu0S3Ol7qKT1Swy+
WTVrdZDVcWgN9O/jcv4xGsW41WYmNS/fWsJmzQ70tOZ255KtOQhOWCCWlG/TI+g5D+cMddcUGycx
92jZzFcmXZ7w/44jcyapTaizEyL75ZJ4o5U7FZBJa4WY6qIykjw9lIOAGu2qTzhQhPfaqxxJ61LN
ox4GNbiX5uBXJmk7k6kK/MiD3gJvDXlQlga4LnHFLFMh6Kccr4RDJevnje82NEyQYHcOMK/njCEP
tCxRjXHrz2AMvCrL0u+6cXAirLzvw2xwoWSjeUJXmFXh0kC2EKOHqo1d2sEy/ZkxhoQIBz491d4K
sJwxt6Kj0T8pNZH6+TroHz/eB6ySjWI9g1BUkxvUTQdxlJUK9kZQoxbgCBQpZerBDV0VliI5Wbgz
eeeEsu/7e2sNpwTL7fnSWPjbS8t834im3lotbruAy9ruo0ILxrl61bmFpvyqkhheQnYGQy6RzRib
ejYerfq31nGCrxeR8I2UjWiWxLjZ9nzmTttUEYR5ABcWJHuccSIcWcxRjh2nDIFg/qat5yvBq192
6FRth7PAnrdDEbSI5F7mBbZEyKWkb8aV+2S5GgTJ5IyuTf9SAvY3U2e5IxBeOer9EhPFyuZiozmB
ffFRe3XGFHQwRsY3uEMZ097FDOfACuR4vcu77802F6U/EqgDzZQG5VKL0UaPCWKTbPkpXWPvRDh2
flQiOxt3QvEXFefTJLYOwQn5TPcv6RdKUgN3Ll55OA6VvOxtI0AtAFSPoFMsny/oww4MUbo/iIMY
wUa1UQouxzwdcv+yTik2g1SEfX/Eb/HWMYjha1IL4z55lwJvWe5vIko85svfS5pyF5oijpZfcX+C
4lOFa0f3DE6RNHl7aoMKZHFG9Ig5nrBbOenp19FpDQb2CSkF3KUGKjt59ZuuhbiEN7BzyyFM1oRZ
PEWK3S3BUDgQWSMFDr0b6ysHzKlGDUjFPN7141vUno/3+YeRS0mXbMkgO22p1ivo3LBZtPPVaZMK
CQsATzpQq0k1bdO0fi4fp6GyoLJcmgqrYd99mjI/i/I9uRTiUaNNtfzlM+ZDas4QZhUliX4FgsFf
KL13wyQgj9d4CYIS7UNCklhiFj1aATUTHZ902AxZ09dcNCzAel+2Af8xcFg/XOlnUWnL68Xioei+
zRhAIoB5D+KAWZT6D5RfYUiQ0zjgnAIz+CIpBYfkUMHDn/o7lSZiNlUf2/zeHBsJvsIWu0Saxte5
q3xbpYficn1f9BKnzsvmlcQMh7ABEtxaZVUtIEUvvudBD4PbveFWQPLU94y8zYzr5AJ2X9XMxUiU
vXMIO8+We3adsOEiZsY8+VHS+H0esW5id1HO0NuSUHEe5IRHi5dacujqWmkJq/AKhiBm3hvOQqhW
T0QpDvqq7Z4vrS/Ve+JEnhYk1n1DdSiPqlETnngwA6vjWbANcGS6lkYSNJ1YvFsPB0amXAvlb9Yj
/3Hf/MlgWbevc5lq2n1qYcpCW7pfuJRDVdYXimy8LSN7WauuIUOflTtKw+/RtTxRm9E0nG713SV1
8JosPShNd49Dch5KaDXaKzHG+Pe28OTENWEPre0PfVvLrLj7gOKOWASWk8/wdiPY3En3DPxE9vuP
wx+J6hVVPD6huqOaCbN8zteUHvqrUe0Er63oD10RP9W491D2tjtGCah9Kd5LC3ACodsXGkAveyVs
H1bLRbUZaQNdJHobcG5Iv8YHJ6tb7VmuHlaU2y7AvNsIAh+tA8j2JO4Qo3O5JrVOGLwfu5FpPFxx
qVn76JwiS5I0MrV3MBZll8LWg75fOoHNdbElB5g9TVEHKx9kXAFBccAJwBKEdFNlR7XOSNYtNvUD
g1Dr/iOsre+Uu7fmSn29Nm4/WVklEC/DO4wVnl7NfvFwJptwqSUFe/X374zu779+WgKp0KCRr0Im
6u3pyHpaoFY8hffcWv+P49jSpl6fWTyO3gWziAc2fHxUZ/5UReA3+32T7i/ioMLEbg8FJeyej2FX
ntIWFLkAtQSCsJ4LPx+E7v9wXwMmixSgyaT4FOz9pSYAYk62ZVoAhqJV86H0IJRJxpPeQbw12DW8
X5OfVjvYcGLkT6dBOiD9u16bsYJhgpPdYXIqS5gioLqiC4gdeSWp4scWrEVoXpeieZ5xo3TiMwdj
jKqv8WliGglLPWUnCiY6i/orN+LTmm3OI/edsuzbkc1rKPfUYq7N9ANxCRjgvr8kIwj3zZKtVPRz
mNHg8Iukutu/y2ksW7QYutbEVLWEfztj+xzpoVUeqLR/wOFQ2wGrMJ8WkYQ5mOItAkpL1zpiBUTW
SPWJazESXRmPOAD/s49AumCDWJnL+70pnWVX4JaUpCd7rljxJmyca1WB16a2Dk872M09O4Iog8JU
6PqnoIur0V1CPa5aiNNnpHuH7fhM73k3INe9cdyiTue1CE4cbag7OYyHNoSbEvgp1lXHWHMTWQHG
LaKNT1hV9IYRCUCLftAqAjj2B0mbgD2Semu1NK5JmvaTeriip/lh1zLEG8/tAVo5MPSsbyPJCH0N
g3RdiV+MGFEJyVhzH2Nqw8m9Fw9NTxg/u48AiL1kgVbPXdfzynWGtQ5BnMJBh/AfedaAQQx6cB6V
mGNZQg5EVXGDEekr57hBJ4gEwv0tU1xTRr1fMQY84N6DAOq/ZgXE0F3og9nRkcGNaIPidGiwDj8Y
PJdjN3N7Hg7v9Os0TJ88ejPP/J/4GGtfpjk44WNFPiz+AV3nEhFUmcb1uKCDHfVM3omJbkjolzqb
9nEY8vu3VvLwRVaDbLlJ7w4/SuEXbH+ukSj2pSoM6LWAT3rda8YbVt0ncWcVTYPA79aYXYUHBA6I
QUmnj+t+DJkhpvwmMCR4LU+4L/vy+Di35S2JH9GbDInRL+aGxNcvvEsVS4bDN8kJUUHgruqjiwam
xrJQTQwmEqyVov/hHrAovxp/R72PL3rRB8cRkVpu1pJxYZIMzsKZu0R0nWbJO6GIQZMIejrVna8k
8pteB2AMenkthVr9c8gDJEwmF7kqisFWhJ4aHvH5UeIPGueDqZQER+ImgOPRoEOcHZxiSmEXsTmW
KMO9NRCaQQamX58yDYCK8nLwhuf3UMYgznyjT+XLl5uoL0WFqH7fmqCi5/SlqeCFdb276vblQfR5
aZR3DSt8SyQ9RttItunrXdK+7WAbZsPi4ks6MkwQTCTD5Q6Y5OJOfUH3Ec/lem+Vaq2+mo8Xuep8
hN3WLCUZ/xFxaWN4S/tVs8dSUach9mP2hw1lUaawekDZn3nyeV2Bfs9LxbGWG2iChgtXIH65HPdT
b+udu396Ka0oxroZAUEwMImrKlOk6GTFLmpoq+ef0EAFpkWVrjcDXz1WxWRdNzvrADHU+85cUXh4
nVrPHyM0rqwk1N66kQKP2z2xGmTRpASG7CK80t9gS9eyOiKPwtiYUnCZFypED5xm3GsO7P6miL7w
k9v0+ubtdqsWsSMSpsUWHGs1CJ7pEF4uPPtlxLmEg3wKkbyLagt8LxyN4j9O8ssoTMiGGaBmQI18
aGLK2EpnS7NyD2vv0UK7lpEoxJHo/CSUpIA7ZT191wJPpCFiGo65a97FST09C2KaMcQySvSeky7w
XoZcUKYJPllfEb2yaZirokAyoKVmDKKhlzXvHqLK0Ra0tijs+K1S/8WO62Stjd4upn0uRWR4cxwJ
EN3q/jVRCojtGhOjUh9iaPCPz/V01Jq6Pjhqla2KciLGNn/dRMmg6vmybV9AJrRweSMwA3eOIhO3
ZtEyQNWivZ2TspqqFZ4kXaHi9+m/q6jYOX8RHuav6pYCGLSxK39WyVYrHWm01o7rdcZDZ9hG2wpR
SS+NYErSiqA/oI/DXcycSxws5kzTJM6eyJueleU4vySM9ulycSk1dihD6x4vFsszpP2B6/1dXLMm
jj9KglJYktmN26iMOkcRjfchzVIaB22CQVZW0PXbDn4Mf0gJlZ5lV//xOOu0SOgS6tta3jzGw36I
JRXnmfVxMJ6nKW3Ns5WllHEHjH407qfd+Xx8WgqgPqznXwYN3hdx194wc7cDEFElLr69SwFoNd41
o6TYAlWaEJ7Amu8fdm5hheHinyuyxxo2l7kA6PA3sgU9oJUS1vUBaK6d1d5gSIqs+fcj+FIAdiPa
Hn+nX2rokXnsPhTBI3AJehcG4QkYZ7eh2YTF4kEn8KA3Cg7AbzMaHT24ADDrZIqFYtgHBP9o/+Id
G3XjWa2IiKRrNeNfUFavnvDTnygu+sKrCgx4Wp4W1i77oByxiXErDF10l8neEAGQGkqrOYaX/KNq
AHOy2wgUC4ZDb8184ocTHeJjx5RWDWPhpajjZAKoLAjOXR/gHaDgZkCXmjAzMPWT1a/pMfY1gssA
T+pjwne6fukqqlKZ9s9ZPTwdfCrX7/ItNz2dXGPB1EI/n/QLARl1jKoFrIIZc6QfPkJKDnIQsBPR
cQfgawH2u8A/23J76DWFtJXQMrOgi5lV221n4Je5TxK2+/iDdKQQTtf07J56Xqm+DAYMR8goT1/i
v4F1nYu3cfMJ2QMKQvV9kkRnCwyhP7448jMZF2vTESPKr6KVWoFe4aCLWIGArVcdLCp0jK4Y3FJp
xNhJf2SyC1DtpF3eKTjfVLbU3UokDuUU4v/jQlw/+6oG+cZsNthTdn5smMUMWy+FKWN2Kd4DpFHc
A9LpOBx+BoqzA27/ahKLGMnKSEx0N1mA58P6WF1bD8/z4udoCPPbysm7771Zapt7nP/B/Wla0IHs
Gve7f+Vo/5hlP7UwYu2yg9/Y2xOR38ywt34QYqX2cxoqE8H608KXTEvD9OJpgO1M5xkJ7S+b3xJ6
ego7mzdOUXwbmwXvmHR5a8ebaBDBfo4yIm5DlwvJArsspDewc90wVWUV/jjNXGVInbCpnnddOxrE
w0up+1K+rLGRroTJBdbj9M8eqW+qmShh4Hy1WQ0obq+IuyWM9pPZ63AzvgkSZxNT6Du/5VPo7Bjs
YJ2k9non6jGFoksVtkVVhqikZAbu/R1DNCgRF9Eaknl/CZRUjb/q1Gv8a5+6Ae4jgxIPrCXwieo4
YFNSMkYLdfJj4w2tmmHJEFtNPCRfL7NTkliVDWstWr9jGxfOfqAL0Mb6kcLzelcXJc0Xk4+3cMFe
CeL8Mv5aRjz3D3k7VNHOP9k2zE9rBhLpKjoclkT4FNLmeQf78lQm4ASHx8Y4s7a1sdM07TlFppqD
aLl/BtLt4cgX463p5I6EtE6xxbUr/+9rm/YHZnbURismcfi2fOTPLokGyY3Nwwar04Wq6Q85vc6C
l4btOWxZuDkQDGyePnXCLxUKx6XAuNT4i51JizAznUNKlPVXrqAX/4d457n8f3jYVUrBFxWOmtLL
PDAJKpBN2jHTTjRkM58TwhHoGNT9R9u4fEiK4irGVtvi2RTuBeQ0fitK/jSyYOJPeegcH3AOzBdX
X792DXpw0So/pe7F0rHndCL/y9U77XteJDlX1cYNCCIByH+fpbEu4vinjDnVbR9pt7MqbFQwUka8
uu2lI7IP0IezuxYA6+ya7ijGOyPn7dIoLyq9AgJxuxq7M5Hv2UauTTY80Pw1Zkuska15SYPksTmF
HD1/jVJwqvVhxmzLBz1g8x1Cydle7HxkF/fMm5TBxdci8SmUUXyZRmaw4TVktTBisAymn+vw65dE
EbFwijfP4ftg3ZCVhKnrIWemmjeoY/y3I1K254VfOmc2SQgiewWYNtStA/ZzGXELaFEQramzlSfl
3QyYh3vyu3BUUYT47G6RAqlouoLSxUcwjnQvqXJMT548rPe8XhMkzXLgXQurG/cXZTitJk20kNqU
EUp5QxX92kFk6asGjLGD99dAX+mLhrEkYQG7Oq+Iz9br6rgx65ArGJfDE1lzGNu8moBIO54bjPfK
STm293gm7ubpfTJMqgRfH2h8Vgk0ReTqhlTMCrsxgFOW62c+AL2qeAMpSSHk9I/awvkM+F37N8U+
AXehBiwYDEhI4TgIeYZLI868daiG0q1M8eH+c5imNgjdpzz7oNQCXT2Nbg6i9QJxT+3JVAFlJkOd
uhk7EC/6uc2l+JrUPAeA1ltLqjUJM4TJ83n/i+yKWWxhKr++y0mXd40YPZcjt7nVu5cs4irhq/wy
6qcZ/5HOIHlQMNsMhWOC+TWiouNeh3PmbM/9yITokNtWX6NhSPJ60gPOHFFwVflJLf21TgRN5OzI
LhsA3Jrp+h/B3Qc+ynTBjbpUlXRiaKIcqVkk7slZT4huzhB9m/56FN++urKumHAswxplSxsjOot/
zujUiNiXWn439gM79A7NtDenZHhfKvZOKZAOv2dEi3tNNSrFm/Y+4z9kfxhdnwD2/Tlaye8nysLo
5YN8AMR9eQTyBgAJxVWL/6mxxGVEuNGt8EQ/tD+kBVbUQWLEb6SrbL45UOyd+mmWJooqnxyXP1Cb
EiJfTQYRZvOdQPShF/SIimjxF8HJ2qjqdlDIWZUv+VCj+l/jq8JHLLOWYUFbnA47PANYgZRCf8ei
dORKhPz8Ohu5xnpFKmV1Chnr8wSv96VufZWC2zowdZGLdAAHuViYv9lDFNoZY4cbanq6lSN9B0w3
1rYdgjzegDLI5htOi7CTNfWS2HbNaYDpWkQOnAMYe/HGfKl2lbcfWJqi+2v7NTNO0r0LlAGiQdD3
xsUjmToshIjkKJb7jTaMJkOnFgNVr89KO83jjXsLnUMeRyXd5WcvxeByEDg8w5UqhceVQPb2FYTE
+dKOSsuk4FuuDshOCncLsGjaRbiPgGVunt2Ld5ePejxPDBX0lahsc3CI6YVgjjtnKBwjqs31s11q
CNQsng0747MgcZvNQQM886f02Ln5QvN6z/Hc9xkwotTS1jST9DiyK/9Y6fGwhO4Wx9KCM6Kv6pAr
s8ICxH+DUnBqzK0jimYS4K4WPQ3ZZ9mWvaXBHF7XV7Efr8Hhw7EUKiz/QZ0c5kXi7tyYb7Ejhblt
tnju/5o1gBHkhlwCYYkGVI7aL5Rahk7SPSyNkpNGizvqx8hBRelkwy/Ms+6Z0edJ2FYO2SlwPYtV
shhEDXhQH/heOL3RIVjjpHqKPykrVSCa9jE2SflIoy+7Lk4+J9rvbdkBsP4bCFCOQLfjVYvSerHE
7rRZvQSoDplj89WOjp0XQVzpA7Nfa6hof+VVpcg7DG54GINfeQK5ZnRcOO9S5r0nuxYXjbwGfrfX
4oX9ZzgRAB+MeQkXk0YWQoA34oRw+RJ0VgEQXWZAdAFIxFdBGLTS3mxvSBV4hP70X8GvdvSBKx2A
+48P9nd1m92unHv4/ayVxc0NB9UvW2zCvvFDqrN4UubYxltW4UlYajmR3lN9taEJGgzq49MaThbe
QT4pzosJ1iT3bP2LJhW/YiEdKMzT/LLx+GBEco68WVblERKrvWVJkG2fDrv2/dfqzqe4WLb+J5Go
rY4EdkKtV09JnLHuxs5L4fMcA9HkYqQu914wbVRFcsTmskaKmpHGFxxLpxTaM4t+WOMfDhO/gFQk
8t4lI6JDtuOuG+nZcdJNVvzdC5OrLkxGpRMQ8LqkAB1nwrCc/Wq+LSWRSL5Oe6MsrycBCbWG9Rb5
cLPSedaKOsGWckmuUg68n2gdIowSMVg62pXvPFBJK7vsjNsW146XUY3BMMA/RDbeFk4hIZjnuEgI
zAKLCtIKv8KZzP2VRH1tmXNMQ1kMjO/tVxNKx3gJNvdd6JmwhNJKUN1zUSQh8UbJzb/Ti0pGYgxM
W8pSORQmTXc9bo7qby/aWDA0UzAWdMxAaod405l1BnMJrMQqe2w2QGnIQ+LvNG0BDk8hv5bzoEEJ
Lc/BrQoyj0RRyjyX9jiA1hPSo0BbHEYRNssVIh02i57FE/fdFZlgppSJiUihzDTCgry5KMqs/sUj
EdjnAqP+QVfYzkk1H1Q1RYZRWBt90H051TbVa3hg532yqlbajUYSzKMkGGJ3SpvYeYwofbOqYRnO
NiBg1EDaG9VS/m0+QVS1a/Los8Ee8GuxRUHdJi2XhEa9PlzXvX1Sq5jnfxmZpnoyNbUDr7/aioIc
rJ2jdENFC2svNh7WfxGEk0GghUCbLrnAUiaPQ5nvLDRLe7KE8Dahm/+iRllQLP75+VnWytQlJr+3
+MyMW2HYgy3k0YIpJShF0gMV2naPl93ASJ8d+HKhyf1/L0SOT5iYl3bdex+P6VQ7uV+g38qhiNks
yfA3FEWbaSpBLCfCoVwRdwymlW5OB3ivShfdhWGymm5oYrumFAgzmxK9w7jLudYYkPkFsh6aeOeR
YAH1s4N69BNYp11o9onLnmJc9e04Caaydb7dj7t/eBn5SqmU6VsMWL7ujZuohUaNSHBpjyHySLCg
bKgVzBau2a1lO02n18RJHOiUnoZ/tS6cfqEP+vfam2lgrMpP7uTjCJeyjuss+ey8TBA7bcKIlHso
nMbwzVLRxGJyNOi659BFDyUWL+9V1q3zYbGRuu7IekQ/F55RT6OGxbdhHTR+cD60nEtE07y24ygn
OAsLhwgL2x96PO6K+gzwzpSB+Md0OnZpNoqk3dCgHyLbqNR/FXojTviLN2+Yc7OPozcTvXKwZvWM
caEGTObRBTivxLhfOJAoxYPv9cDLphoxhf1x27PzLWHYHHv2Jmz580Doj0pMy0LHwjeOTIQ7PtA3
zUIKXYDVYXkXxrt7V/IxFkg2gRCZsOwIJeNK0YN/4YmS3HkQ33IOdP6DlIdtaMgITxcVSoCz/Rbj
qz3kdZZwVqKp+xHYvdSPl0mWj+HrE4Gn5dEQqLADIG1yS9xIC1uRy3F0gSyW5ltl98HH+HG7qPPD
6KtG6fs6d9+cAzaPgLHmLe9DMcE5Iw8Oc0MvWiUaR0lFVl0lmqw3A7+6USEpdTkiIjPwRYzuhlTg
KTi8fO5/1Tn5o75cP3jcZGII4DDWr7Hb9PCX/nWFIkNz1yPpUILEfuu37F8gchTad+jCpjrS3PHs
wpFZwmIF8ccGDEOEuYgWzQXAfelhzlXwt/p0thSnIE+yYGomav0mQjWPNSIIzZZZ9XiX7ITmfRs6
I6ZJul+19p1GV+5Uv8ItdzU6lZHP6FX1f26pCTT/tKf4oJqlrC0V14Q+Z0CfXIsqt9KRE70wqQMA
1YeQnUvV21ahg2iYZThXtAnXcgZ3AXJl2gTk2Fulw6IrCsagdjdOzZ8JbIPdT+UOr99SHwl2S12i
eMLs04x0pyvq4rFFDpgugwCFCzsKmnLaAc6sIcVwMzKyAnearr8SzkR9N4ibS3w/sQbvkXu2fYvk
6WGS6n71CC4Ti1iCnHxd47nKegX/FAdK0uvdKpgUM1jYBNltJXqH5qvEI2JQLvOaryqpAvwjWEYo
hT1uTCID4kBvlmaVDLcdCn0IoE3yY4GYvUehy1Pjk+UFYkLIbTLSyYMFHOyWA82vgouBMGgiBxfs
rch6WoPbO7DTyhJtn4guqCMi3F+Hn7NaebpgGMAol7b8GmmqO7Ct5bmNsSLlJw53shi6NAwH+U5M
rKdmodGD3f3AumNVXwJTU+zxB3sGCPIkMRmpr5q6xV4D4F6wgu8jPraJGt4duks+Yn6rrnQphOfx
WnCIr0ByrSpGccOa+qScPlpLdiL7w8VFPeGqNwxSuXmGJHsqRkrtJSGUzNqsdGpj1Q61PEdWGo0V
EkvhkMaRvrVSPrFyMmEDwjrcZrvyIQLsiQbSA1HZ2qNctmtwqjqCwuptyR3H5enzvJYfpQ8yGAW5
uh7ia6rHTsdlrHQuaBSjEkNFYWpnC4Gbh6cYwqwRMqSmg/IJsHFM7NCaMeInv8Vu/UxSfFR/aclm
M2/Y6NfcMm+smVBcNRGTRSuv7oRfvVUr+0B6km6tL+rJLxGmd7U9iUI29OngwbOgClYvX+Aey/Io
vOAhGCBB4lW7Wr/rSOL4nAHMInzab2Mu7o0fs6LteV9UTxyqozZeys6gh0/yyjfvQ2wRWCpVofUR
4BeNfYmdQYse4POMgqS6GIcKKzUPVd2M0s0fV8Tl1+EjSHYiCuQIBnSBLS8HrZ/srCd2HuE/6mvM
RiIaI7KalEGG2FELv4/4EjueGIbXRfAO0xeeq41Jx/hf9AVuGuBUKb3xj/iTUVLla0moTGzrrJ/g
Bl36BFyzqT9X0o9apNNZE6P/CK6OVgH+0QTYOFJ/SmAcjZMdks7eebXHYBT5plNOtiL988enVEJW
I7jhXeOvpNp1kz4XMKSPaLXMaoIAbZpATNeU8esWM7Fsjwibhz3hGj35B7KiYYTQOstegmyUEVlj
kV0Bq1U/MHPGHN9RksIn48q0gXnCjrhFZHsJVsKI+kxPVGSlMBChZtbHkkG8xGZU+GkvStJcrtaP
z+krz5hqVAUwTCOjhdp5+6tlcwcLSVBbIa5XPMrYAQe88/UMQu1prd5W07W84fURZ7jBuTMEZKFY
S9OBJw+cTPueVERvAz2Fh9V4qIyVKPsuVs4uyg37I4sqg13oBjASBO6qgXjm8DGtBtHMDmuU7D7H
NqrSTEjAlQDIHOP3TXEXiS25gx8LFCRU8s/cDL9+F6VjPNZXjGC4g0apAuif3XvifFA2R66qpS5t
MvPplu0LfM9oUaM6PugVh9k1xDlqNg/6Jx+hwtJSEIaOcogGsoUBukeWtBDpeQQCgDQHdEkkjtC1
Npd5oIcqhIkDpCovf+x0k80gkbjXxxQjzhf0P+HJuAp+n7ugrixbwnn4FrFUYcGZyeLsFlW6Dr5P
4CRPhVaCUQdx3x7SGpiGDA30pJudWzp7kpUz/tYpORvXMhyVKrw4iazqiKn0RyPDyXyja0I+Kcwg
FUeeiutnpenyjgF53mpnOj6bV3hFiSPVKgUNZ86jF8b39aMVAwP4FU7UePCJmGtcc2o/Ak44WQv+
TeQHwxzOP85NuKZsU7ThTlNU7MpOyPvhKODCR0jOgGKu6B8kNialJiN3UwL/+zaX1XhYMmVq3857
va9ar2/w3ZhKaN3+y1w+AMV5Mp0Rb98FziIfyBk//CfUWTeC64WWlb3UEcC3utkTlYBKploDnJLq
U0QzfAU6U1yCk6wlXGMFfKPFpXe9DG2apRtHdzAPL6cNPGmuntY88gfXBZrx/zC3V9dks6Z34loR
UboefbwqYDJGKw45WFlTPJZJO1Yb2THJHGqA8FH80dk05kBoAm03sH5T15EpSdZO0p6QB7ReQox+
9bLCo3xrsw8tOa0kCq/Y0gSpLKij5WTiTdiqoKGm0/RaYyw8qxmdOgqSslZnN+dXC9ekuN1320qG
VyJmQ4v170YqoExKEb+Tt79YwZbLVd40VhLydhOmaGYhNMmZ0qvdj6fLo4NYPQCqtmnv2mnYLX5V
5HXEDXbqZABQcTBdWMRju2bqffppICbwj4UKNcFAxEvWdoiqaK3HQrB5C7kDGQRLGPF6pbQaK1Na
Vbo6DeqvNL8muMMjKHjClQxH+y6lSgd/pPGZh6aeZyVdNBai6GXTPdPGF2DHb8dJNON+zGMpsX0Z
QOfQI1tAJ6LNtL49FFbJyub8K8rnunDJ4Oeb945nWNF7uJ593t+IV57F/XVD00Y/uEOs3cWvez2E
wsosQx/TIvxCllVdUWk5gdo75qeI5Y99ySHSYnDKpm3VJYVdl2tV7djoYYC9G3S6HcLO+Nunh2RM
kRhj1OM6WSKdebSbYLVfKolA423a4HzTAdEBP0m2FGlJRlqMjX1eAz5G3/dMutRBUYw3s9GauOZc
eTIOTZQ+tf2sOvGz/KyGJp5dfSfUuc0bT+sZxn8q5voy9m9nVL6U8QK5krva8Vd+bDz0VKq5x5BL
mHB9KddnGcvBk5O+GNYR5Krr4j/YkyobFmL8529kx2k6LOFHOsmtI8M0kaU7pVRll1ByqDkK/XyP
1pYu/tkpvoLHyNuZ9BDOEA6VzQ+Tjeo38X+xfNGu5rjH2K/aQ+vK2wJy3QQtSPHtGJXlhbjGQcnD
LBS3MugCDjQAoORq8uFaJriiCSvlFz0Q0/FvU05jI3D/bp2NkHoGLeyM/27Aod2ElK6JFWYXA1ZL
x3a3EI6Qi9J1pUoeO+G8kY1efwkCjIDbjdS/DUaTS/u1s9lM16cQ5q0Sy3DxgBWUavFkcYw0w0q8
7kb6oiXT1zZ74TbW6CsATzA2hMczDByfeJIkJ7rUtuZCEc7MISvQ2Khbv2noR8UWLymsvJ7Mb2ng
IiLxsGNDXoE7XQGGfmNDhyR3FO5PSNr2SZ+sBJ/dYd6NyAcx6kNx24ByJK57HHeVAVcVRoD+IF6+
B8UdDcofDxj9A0TOsH/ig7UkZgYxVnJ2pAN+67I/YlfnwzrevU8SZsUuIZqcBKZY3KvD72kKBmKg
aksfVXWpAc6JEs8HBBWCeB1wNBfBC5m1IXswad64n7QdCUnh/C9IOJJke60VvEBeUGeFjp70z9+P
8kTcrqcHbErjBbPII/+oZ4xUFGWBpURiAUCAAIgd0YR0mzEMT0grJUChu4NS6E9lPW/jsIOQA9oB
0f2pEe8kXAMY0l0eqP2osiiQGLkzD75a4xjMMU+fG+gCYSultIQcXi1q+YKarXanrgcqrMGkVemf
1KxGZvWqKDDT7Gp0jxf9Gl5mwx992ihEAmV3KLALVeNFhg4f+K2YscIj6bXsDo6tMCD65kcXRlA2
ZA7sJWiwLE3/yjkqnGrL5Mgfe3+AGmGUgXZUGZl2iIosbwBtuwYiMD0Vroz/aoptYAGgcf2Su4c8
lq7VyEuXZqmC76j9ojkMNTDC3YNjvKRStlQMtjwc7KuuS+fjVfBXqza3neF5WIauaNIsF3DjKsE4
Z1ydBOuFoaZpyPRUXh3kZIogoa19EnNBOZXpwdo6fTdZvyjXb1sviZQU1bXCVrK2D9NHnoqUaFxV
6FVBQtUC0idpc9fyqRFmzfOs3rtgYCUalejEgK/HsorkvdkISykCRfPQxg5D9DjXxirYV/MH9I8W
6D2YGj32dKec0I86bcxp8CmiIJxy/muV7blidD2/UttBRdvqJB1bgdeSWchYqGa2WTeAsBEv+1H7
gPYlscCfbF7xQDOCRgGAbdgix6cPbjrkXi7IDRn8tB7BAnRDt+0wUzw3Dumm13UnKaMR8xfIuFmu
Imk4ZsbUVOKKE1UMI3ksBiI6sgsztORYTb8PRIywdlAsgXYw8kHYjsy4kAxCb0yex0UlxyI8DAPj
2yQ8PjHldgZPa1ZrO0ex1pBnj/R92qBtu3APCp7507vq6qmPDn8aZpu/0mHV+bCPyHMiP/6JQhoc
HD/HSCW8jYs6gSH4AO/FRVh2D6LNeBJsnKD+eUIbGa1UT6cO59uq/9MfEpi5vIATB24325+ZFzG/
FjJXh55af7Lwzvi20ZXpzASog+SLhY2qVUXB2/sU/eAcSmyyjpOtg9ymuRcmkF7hvaomUDnAgD4q
KqQZnejJflaDGvAP4Df8zmBRH68X6u+NaEvJzMLyNL9RT5RTZO416qpEUwN/ketjZv65k0QKp43+
HPbE4eBfRGSYz99YkjYH2wJd4FvMb7PYVF6A3YQjyA0E9J1GwZ5Q6WKBRbaaU2Unuk+aUuUCkMac
a0PamITMiQ0JUb0ds6BTlzOGywi88b97D1viELXduBsqk6t8I1b5ut0Di1A8bSeuaunIfYI00gvG
ZsZjPC7OuGvp+34I5M7+U8TTw0Vl8WF2MLlJI4u4zYhy4r4M1tTCFJon/vTqWzejzJ2KxPds0R6P
RXptvE35idkPcbv54k19A950lNQcmNdoZGUIgQ8nc1Yck3x81uCRU9XPxbi+Y0ESDAbltutz6Xai
iMAx8jTvf70ziYoWhJNBxR6zbsoYUvYFmVBhtIXTvxhgPoG86ly5QpIxarE5IRx4isGz9Eje6C7q
ppE0NWgxL0rfz9wcIer3oyWSpnyywRPQb3BGD/+WuMeU8CQOB0TyQ3UkrkLvBM9KcaE5F+H6wLgl
1Vmwpj0dICB020NuLxmVLPSHFpsl8bOpZELMkJx3+ARGN1p/gCEKfqO9sCSXnNI0Fie13yKfZxxy
nMZtPZEjhtynYsQn6Q+cypMsP+Y9Rj59fY6WzPGYKZhwG8S8vgFfqUGKcYGMHscJoABWHsgJqBlB
7rXCKwonOthEwV4Kbpei66V77eLaJJtMOG5IbOHAU6BTyRAZcn2V/Cc+KHqAO4AkcLdco2V7ALxR
hm28IZnyqGKfAaSh7IyWv1JCwJ5+cbpbaGqE2Sny3f9jr3Ai1ivAZkEtF/ph3G/qVJsQOn4H04c3
avu3Is+pMIqTRceo+0iuc407WvJzr80qLRdbT+9dm1qOhPvuGgKtVfgGScELvSASEvFi0jfhA9Ev
lWgyMtatUmOm4pfSKvmY9/t7oQSFq1W6WQgfyT4KGEq/cjwxtP/q5aph+2nJ/d+gyEBSke6VmkPo
3GgahGN2q5LWncn7GMQwM7dUuQEdeg38tfE/edsB6OtAw3Eioq8PcWOKPeZZxrbgJA/Y9axoEYjX
IJjsinku3wOdQuSCcVnXCry4yDx+lKUgqfnmx9wTQ7c3DYWnAVrf9xWmsCy7FJi8FNu2F5UlGkkD
nRAUY+/bSXCjI/p99wKGk8qlYiWd4CtaN8rZx+n/qJfCqty6UG0XU20wUSK8I8zWzJYqQgLAZXMn
kVwMmeRoXoeEcpDlmu4/Ko42liKslBqtVtGqbE2HEUKdOsPoobmATEVIbVgUEuuamKLOLw+GiLwY
dyKll9aPRHMpbCIbrKcyvQBaW5zM3e/8Ck1vHv/qPlUVqDfAA8KG2wP+bIvC2ma2O92XhXE4W83y
/p40vOxGy8O+A5wVHLKKX3My7hybOyX2WLr9uoxIiP4hgaNLJDCzTFVHhiJb/DdteidISOieltxH
jkb/WqBkn+Y2QJlTlxtig37BMeOCHQTn6qg2iDhvqdKl56lD/yxYpVV1tAafylHp+DcDgx1Ur0B/
KplmyDuurLGxjBWi11966NbumJLHlGuuUHXzq7O6pAsgyjwZO8NVY9Y9oCawCqLsTFIcSSomYy1l
oL1r/eU9TA0lsDxB1BzkkuN+0avDv8UMVgkhvUeYcb9zUECgkig5Zatj/PxPLhpelPExEZElak9/
fW6TSGmB4iRkDa0p+5rfJEuQHYwKhoy1fVbSTSrFh+ixWOl4mZyIvzDXLrirLDpHv+BbOi73rRTY
bDC6veSVh5c7YyvS7h3STJZAd3HwGQvrwZVxFZONeAPEava6GzTzkF0tGo35ibz3/RjX54FONJQT
Zh+ngYPn2BsWn3uT1HCi+mjUexoRW8BAEXhdwRyJrtHSePj0d//zBsCCZD7btyGmrPYaRT+H0y9l
T9PgEJ0uPZ/vh7ZFOOW6P5TXc/fGls/Soync9/C4QtWhk0Yy4RQB+2VrVIptjFYtWxP3RtD7SXqm
NVVKaGIih7rj7dE9gvn+8Ul8KNYo/wk3WRpt2m5M13GfYiIU+gJO6SouVK/59wY1uH6wkEpoVg1X
bnYJ4xYdSmBa911DvnGoV2X2L/17+3adBBl+YIsHqXZaaXzysaVaJbfrOoqealAEfBZZ56fVf53V
aCFQvg1DQeIsLLiweL4vr1nxTd774IknTV0lgTp5cZaULjTx74kgfq8cTtAigyDY+59AbsPPqYAt
xWh9zngu50vSt6CjvIhU9xFMarhRAZkdZuhK4akCDcEBhs8CHder+kW2ICleajKet2dum7OyDQis
K01NhXocMIQqk7h2UMPBCR6gnKdn31AAsVpyfcZBGrShzuN9xerL8mpgt1sJ6eS/vRK9guIptKek
8Y9h0CBMkA2HkSSQ53pLKNTig03QdxdnMBuHpK6iBEQ+wVhuaiM0kGzgybI2fUf5TVLuRcBcwvFt
yiE0TVwdyLYhBzWuMrE2Dg0nsGDUUw+P5OJN244+Y9oyZAfniiemz3WO5fkoKdn5a/dBXrzxczC2
1BSl40FNqwD0/FLhWWkseLqAqMOuNnfQVRzdYZ7DNTRyHhXQL0GolsNzd1tuohD1RZzpTFrIWreo
U+0fxmrmIUZBFuNBFsutwxLboSyGqyHcb4jvFcsMR3Sm67R1KsqHRbaz/TKH8yspR7vH/TvoXBTe
au6gPL/xdR73YTJv9eMGAfsg6HQoTNug8ZGXZ8tUf2/mF66+b1VQCZqI8B9YyrYgrKG7eiNexyxl
j64Ewe/eE6oq5Y2/+j2YVogGr5sBi+2PV0g0M6+VOzAP9zCjEJ5eal+yppMUlNsy3BgZHofuw+Bt
OWno/aRhqMWbw8opSwxpqNGI/1kHbdQBTCV6zFazHgIB9AL11twqKsOGJEI9c9ZMWWRsh/ce/Dvj
uEM7RtEOwax+UbPqV0Yxl3HtmBpWj7cAd2aU1/lBSssDkppc5oUsXnB7TYSEpybaodT+JX5JVoU7
IBV1Cal2DOL3va9+ynv2xNHKgj7mGYc9toLs0Zpw7kmR4jqOzqKGM/HwboK3aarhFwJBNuCStG0g
aV3oMjHuEOS+HqdwexMT+F6XlVVjMfkKYpM0xJnJ0WL9UJavgiPlSE6Xpp3OwS/pAoR1iSzSNECy
9HGc1dBdKCxDt24h2Lbz7WwdIP07i/RAKXP6rKprfGaKa3e5E8348gvnUxH38HrFDabTJA6mx5RH
q7XzQ/C3RO/d8gzoPzuwyUgkvf2ffgp8ZxY4ZsHtqUMt/3gFz0uq88XlmzNgZKBLSCw1GbCCKICl
4V4G2KVLqDt/C9N53VctJwkBr8wBgGATJHvDMLvBaPC4SrBSozafMUCQhIjtw0baivIlIXZnhnFV
8SiYIZVvbnhitiOZboFq5b0sCQbUfak8J/DPASQmfy1jsK5x/NaVaew3hwWnk/9e37w6YVIe+ZJK
oaEa0W4ZPscFYvAXGuUShORUYkLnVGm98JdiX30zOw/qd1Y2+D2FI5KgSH15Myxx6afX66pB3SY+
yDYD/rAwsbsoTIJKHVxP9nzMhkhVrcG+n+r8hVRvh4+1Df3zogni5VxrTmpHwg819/M2VbFR5hZO
cGvLEEfd6A1+2RQ6GgamsFI84eOL6EYjAusXqutOUblMttzUktGrq1WOd+DTRaCsY1gbRvkUygAb
+by8kl+TmgWQiYoQEI89pFgcz417Ilzmj3wSwvA/3vCeybHr6ZFk0W10+5MAS0A550FWKVC3A2Rq
AjjQYbmxcb9YYiuTD8h/MgZssOPI2aJoqJlvlXj7ojyM85+e8S6E66imLSGZy3o4AHz6KrTq3oGa
2QcQBLo5dT/Jrm+ktBVR6rZ5dGCVvjD7Svvj0KD4z3h5K0PDwACXu+VFe6uPgaJ2zW5BL2yuxgnZ
SelcXJJXaQdqIJLh0wjTgFibKJ/+DVzbmJ67qtJaF9rnH1ti7abTtzyajciNSbJpXuyQM3OupOLz
tL7Z7sbzdu9jhi1IwV0q9ZpRODXARB121tSii+98hY9ZYtPBNmSei2aW7g5OoszVxAoWpp6cQMOE
IV8hzpXIRMRNCRXiJOFzbLPb8W7I3qIKTUQXN+yZwJcfLoCy3hE0+86JNjLToNbbYIQlXyn2EEK/
4wGzmEs7FyaEkOVJEzsVvGwh0J3LKBXRnR4temsfifog/12O3ntX3jGE6hYZNTBKnoKClsHkkFZ7
FZBTFhcWB655yC+1eo6c3AxuZp+4oX4Hf7ZckNEXiXq81fD2rMR7Q4ScS3wjvsH/eVbmII1fTQ51
4Xa/EH6w4LnLhqzgsE2SastwVS8U+VRNL2EhO9fpwVTUuM2l5TZP+e/Z9lTIKXK4K93506ydbYcI
h5pJ4r5BD5H8Olh+q9L1Cl3f85q1e6iO8RhbsbwxZEijVMPx8FPLHeTcPtoENUHT279E5lYA5i0h
5c5Qh/uq7378naDXZRom3vnXPp3THqceDLfxNnxDX3aKYksVakI6ck54l7QeZeNGsW1sp0ynO3Ey
M+wxgP5RgWnfBOszdAn+ipvRjfLjz1VNtHzEhy4aS0ieHUNedypJve/vXSI6oa8tjxj7iXdLt4eo
LbvopaLCz9en+7yD07FHEdSqZg2EgXT5IKvhFJ/AT8GYSJVKW/F0TuuxBzixcB3YQU2XpZf2UQVj
pxoKKmKXoKLa1cZmKvWHH/7MKROKl2Nbf/ya5+7IWZl/3tU/AMmbxJtzD+/Bf8G4SdylI9HC/AVn
ef54XdOu5RaHV5w61Efni421efQ1lwYa9IFYZNreKAZTziemTwR7JwbrAZbvFOo7E3Z+/zVcueh6
25HtHjV8Z1gN9AUy27ML97Jj96rCwv6e+sV99olVgvw9KCrIkopyX2Y5IvTICht2idLFZY/LD8oR
Nbp5zEi+Fqw8HIi/SwwhyNwagIGmYrFlu/jTKvv0pBlO15dhGLzw49795Mo4g0BdcyMTn7AUCThV
k+TykGY19wpnckNM3UzrA2AkskEZI9vW2Xwcp118zsUUlOC6mBIUQ5MlK7B7OAqiCJRomzGh8Xwo
uWsMKSP9Jc4FVs37Q2Jx5RTXf1NcNzQmwx+ZbYhpr75bzHAkZAZMI7DNB26G3+0Nroo+MSX5MFx7
aFzjdG4+M1LakHbxbfNZ3deUoUVyi+bYTk8pWfxLBrxEL92BVJolp3NlJoFhSDrKr1lhWqZCLkAV
9+EBogD2lEGbqLbqnKH9NkSWSEh4Zfq70rqZYZix0PQkkra0WegVjcwaihL5RFvI43Ah9KMzivi+
od8Ov9yu6bS+nom4YVLGAyADqJFNZhmiUMf6YicqhcPD5r6chq19B0pkhTc35ZZE6y25RVac+EQN
Gk75mCaFQNCaaBKOotqfcP7/vpvpHYwIKQtQvwFHD3S7tgIiNrjfyKOPBRXFh9kxv3S00KYaYiOk
0U/EHEFeZXAzFkKpaXoXX9gD0DAiZDxro+KH303EQX0K8tIkJJzgSsgf6/uOlZXldSvT4wdBJilt
b4kmvp/fqYM21fWiSVdtACcbGd8PqDpa5vSqQ/WceNrJPJ0JWABoQ/S2gCxq3hS5rCGt+ljRndhV
mq9zYdTM7/ak3stKtHZVoYSuae1Yreq7vCZNQQ1HdjmLYVK4FnYi85UXtnhegJEnStPo0U3AFwBs
oHh/iinRCV5eBHqpTW2gwfBlntb24sftaWwtFgECcWuxuDTBva4hgIN37AFYPWHVcnEw6/jLhDF9
QBXy5+Z1PHCqQF+mjFHaBQQCg8WQ1ceDQIBDt+vI7F2SglfvnbzskJW0ZDGzI5ppprdPnfz6up2G
wusQVOYMMkXZ5tOBq6raKoNuNdZSsdw+RaC6zC/dq3TAA4PT9W9YDtfX+33uDmXazn/baIhJekpP
LyvCow/nh9lCW+3Wddzc/ZK6ZShW/KWKezUtIhDZudPwRNHe2XELujtG2ogt32BsfDy+GRI0y8EH
jL4AYhfHdhN3Mk2oln2MlFoZFiKTIgvOaUxvNRo+H2q3IcYDpPgJmITvztps/GQ2llGUgtZISVZX
xo2Fpw2ujV51VhHNhJ/IqJyaDTbmNdjz2OaKJV5SKPlkhTemjK6vlDdGkYpnsYTTBIVnPid0TWJg
mFlbFuo0mO8pEqKdKi3FDKtFMpgXADvaLP4lFi6SseAwxapd8pZq/EdYpOjE38rLYQLCHKmlkm63
ELa+9+VpLzqZbjTGMkIaCHeKvrxQHT4+4NRbx3TTbDwvlWPGwX7aG7kHYKpBw453ZsfovIg8A0LU
G5cBev2ok1rgXKuzCATZYrsC7pGYXkquNN7FTCNP1o0zkwQhMm9wZovl7hyAzs0tAWSMDNbHSMmK
BTe74dz9ahJnSAmrz19i/b1XE+2rV4um0PBaeE9DWjYWASYYWPyN7m1e+W7JPVK50s0EeX4+HyuO
/5dFAi6ihPBlVBZuBLKP/u6tbdNGLUyVwBKqgEa1hGYnnpvRtNhrtRVCZx6x8IlpsOrzZfOZm45D
lBtzcEeMZafvNm2+OBQSlfkv+zE3XDVWvbt5vARfRpmgS/AOcEYzBjIB0xEBrb+oMOMwkIx97pIJ
6+Z4kjt4jo3NtcFlsGM70TJRUF/6rOjReoAxV4JSi9x2hrI4YXu2D6YnYxz7sbDI4wTKBLsoLkog
DvGLXS7wcBMvL2GSp6r31gkzTtceCBvtFr7dax0hVdyTVKXA/bdK2JT7rxCAYxF9TC6pesMYXIrs
jZi8/n7Xjiy5jQp2vI+Hpubem1SUDHoCuSyqSGqy/k5boPbXJReqcWWgg3Ob5c3DRiiBRaXavrKy
++Dpm+SD6yL2ir1XPwOtnIWG7sGRRkvv9IDdQnkvyO/uus3+UDlrNXNJ03Rkm5vndXnZPkjjQugx
nMI4SWwcDpAwi4wKF4AD4VCwXDI/nIyuNG851i1KhnhXd02vBJ3nFdnvJe0B+CbvzudjGiAutJrA
Y5xHlpFOsKQENuIeSHclGuQ8AN3uktiEviKsddvNrz9wYE8HLLjSyeNt6eP6F/n+Hk0RvQFwbSnC
FKJJu8DMi0Lhcla2U8oB1yvTAGoN9sytBVzcQUnvzR59hfiS7Aqr6ovJh47Zsrry9zg5nQvA6ftO
gpNTuA3M2E8UtrVGWBokntGcmPUNAWsUdid1AXLF49iROlVQj81CKQB7d0ZlST8MX94N9mf2SMv5
W2zLuyTvKpLEpXN598ksc8CYjVHWxWeHonEkozdhTepaqr3Cj7N18GMfm9DR2khnHF2wOttPiaNQ
StltcuJFSz1soGsM/JPAaHoUJWh5wopIPyEGLxnWU0Z+6YBpGEdY2+89UbjSLE+cQ1WS6+oCAIcf
4DvnmWF0zzb/BhwLvAmoMpHkshIo6qIGcyxzn1/VrFC2D0yKhc63dB7MuvdfvW+LO0t5wHQFpwFK
LobwW/ohwR9ofAcjMdmVAEBYTeVrgRJC2mLYzO8CYscLc7clh8R5FHfN0Yj8wMEoQffvDoljg6EK
8E0+qWdVDH7UEfcyfxu34lf4ZsKtnX9CCzJpL9rZ9E5kBOTazL5X4kMeDM4xOPjLYou+EIIrQf4C
6Eyziuuwiux6QVAgclg1XG0IJTSGrUGvGCTKYn4N9PzIxmiRhVgV+xod24Os5KlWqSBNUkpKLOBm
5mKTVorKC5FfOFCARq18Y8tJU5Vr7kRFnW8jkx8npKAXa29wKzwkKgjXBp5RMe82NqgkTQL1HTBm
+6MvB82lR6W4jrAyU7KWEy15uWkDvrCPIjatRzx9FCcmEQE6bxUrpz/i1aUgd/YgVYcbtfhGhyEi
qqjTxrIpQII6VvjrZIVqmVwY3QlES7wkchlFGa7eV0r/03/si+KSW9nTfWiT+psCieQW0CDUVXJX
3QZvPdZTwDKuzeqnr1HroJxc74ht1chBQQiFdaTQuyDxajEj9HJ8wdvFS0/0XIMJd4f7brNQTYNL
Uf7o1FSxoDFGPDAXZLQjuwADloFtfY3NFaUABgji04qMG32zPnK4wQDi+CvfWzOO4VvEN9pYw4nE
oSZ0aXbz/WdAdCXZ97gAy8BROI0IWjtqT7IykYXw5e3xJnlAPZTTSck3KxJaWxY5VLskQTA9qkfd
9V3lZ80jwHjYHRSH83dL2OhFe9jrV/Or/Ra8h3IKbO4SIa4gRjjo7xlOOtgIanB1p0HUvkDc9r5b
L4rSt0UUwW60gd4fX8a6e6chuUD7o/G72Q6PDZi2iU36NVeFBmrbYkyG8PeCw3OqepbDNgcrWTfc
fc6tF7kGu9+9SnN76vgIwAvxWGnN4jLERq0ElGJjBISRPRSGT8FaDE+2g04rMUje4lM95CGZ021j
jWhyrHMKz7Lzpfug/nDOOgGMFP1pDPFLepia1DJ5CTWGwxjKVkBh7rZ9HS7deca9X+lsyku1rY+3
hBFKMFzJkXVFC1OCKYzVspywrD1EoYZMjhrhl8HXjZJWj0V7zuEKGDuCt63+y53JkDqRcx3RZydY
K/D9b2inEltIpXI+xLLKC+/p6vAnHZnfrFUJ0+w7q0yS1dDukKn6H1BmHwb6o8gla8+iVLDPK9HU
V6fjjcxaIzxpGze0V1qpm+nAo6yJOuwz5U0C3TMJm8+2F4Ai9wkX5zs+1cp1st1+76IXDto4vtEO
UEfgSGeKSankkEoiV4pNU71feiPfflxu0BrFTK//G0vwEToe+gO1WqDAQKQbm71RWLmItqU1cv29
e1u7DSSwcSIDV32+EOA4kIxJo5nihZbyWclsOVRtVj1EbpJQc89jpTq7kgu8pW6y3VJte8h6TO0h
C+QR0P6orEBfaN/JvmBmXh7sp/xlw2SAk01kyP+aeaIIY7o/kjeq4E2nbVO9ELOxbktZraTp7DbP
EONa8TjpIM87f11+qF7KifjxMaad2v+6m6cCNsDwl9oa/nynwCy0D3G2qH/cTmjZPxkKzY8oe3TH
PHH3FP9ku3DK1JnE+CLZJhQYb1Bx/wYWHYhmaaNVHoFAreioWfmfCDBl69rtcvHB22KdE0BNmQvF
BrFGAZECIgt9qjXT+aEQLJDEokHgm4EWrRqiOaA3NYHm9os9sg2MVq8eBl+1fPX8unjJu5Bq1frC
1QMbFMJWKO+xP0pT+PKZxIg2gO3k5djFOjKvX9UqH5JNaptaFTlGWv1n7Tzjv1VllV/XUo6sZ01d
dVRW1iSwWrjtT+w2PLjaic3ZGBJxTp2uRIQDy25hKBWq0oC85h6RMRShmAZpaLJ2lKq/NtB2RbUs
8y0Rc2eyWyorZ1yjj5CAxST6Vh7PPZM7292UnTw+8IxuamlM/tL+cyd62jWcGHde4dB9Ji9nNw/U
Tci552mewLX0u0HEbCXncou5qR62mRVFzt7QEwzMohmNDmkm95XY8S504NzMcAK6ApBQWLAcZLZh
Wbu1oQF0u1FyQliJw+N4VlRR3vPNbeX37lNmwjqWWbzhVLU0aGCD0aramDfgTwVXeKH3xhFySDTk
jop0WFMDFqwARRMT2PVhm/VbbQht0BtJP8RCLDeZG9mGdsvos4Ji5X6IkrQWibiAUHyZs4udtxD0
wzjbVYU1rL8Y3afSUt75apAA7Yre8dS40DS/dGfyW0rVhWdxkLSvUL7ARBNN5gLS2+ScRS6s/Cxd
NcFsI/hmMacdoSM6tW8EVF99l/iTY6yCj56R0wKkc+bK7pmHLdGN/y+YZJLG9MlpRHOhHLUoMJjb
Q7doNBFc4uluUjlTKIIAYD4CirGYJc8PztxJQebhJgI9biihCJLcZNXwqSiX4hsavXhTAgmrzIRW
dGdgmp9/6C3ILOoJDTsX9MvON/JZzYvvXGwMbKKYXl1NHP0K/sjgmLj5iI7a0nicuihRtbsPgW0z
sGyDTOCb393pJxhkUZfrQ3DYPBg8m1UObOFdESCWEjVKltPfzlp6ODeJeGPn1TQjwvNIjzTk5zit
E9CtUKv1c8fV84KvSzXcJDT9D8jUHE2sfGIfAeoqD0TjFdByGZrwFfl/krV1wZR0F3bl3Chpc3fX
moMucZL1UBsSt2nOzxQkYNWytOtyYnNxkq6jGs8FWViCa0mU8Gyc9g1Bs/LAEvfbv2YDn8tkW8CZ
v8PuD1OI5lf75kPuUuoRP6bLuluQT8vUnmpH7zDqqSsbOk6SYCT7XcSzpqqNru/odpHDSROEhtll
Pw7817hrfeThJ7FrAexRLbpD4L0z9FF/cYwJirbuTEH1IKRnhTtPOnz6m+JzeBk/W5Z5+30z0hD5
eFrqYTS5d/JOhCPIYeT4Df4w/SjUnRy5Lw506nMwl8ZYCoj/CzOgXVXvNVZGwGPqYDmU0FS9xNqj
zuNjSOADcsyYRaut3F6bLROuEK4BW0AQiHN/o3r2V0f/y87PdN30DsDRiWW7XNUVfmE0pDkqQ9JU
uhPyD3L3O2Ii4Xc9I6VO90EryTFRXbyX2hUZ0ZPAw105SHPMAm/5h1STi+ZdN+n2FwBIWXY26jKL
UvhSRU8MWxBv1HC4Cwf5g89mVbnS6P+fQgpAuJmQHkjAz4GMxArB17UcJyh7J8PGi7eJQPXjNMIw
5b2Bn7dWfH8fhm02ynKmiSl4oV5e7mEqXlwevhFlb4kmo/6KUI1VYgnMNH63ibtjjf5M6JHKGCTU
LX45Rn0YZW6CiIgYFu+W9TNcnR1BG6O11yz4QT11QPGLzraAjIXYW2T7QOzJbpIDEmXnNaBhj9ej
afQ5OShshI77puWXhSizh/iBXQMwfdrcfPwE2DfuqHtucekUkFexTLNfV0JMTAXWYqsNrhp4XACU
imm3zvIqSZXgSSHsehEqqBwJBusRN3A+oEaAOlibcmsdhF+HA1M5y5IRrXwMSsqtvtqiPzX98JF4
p9lwXk7m4818WCqefYMa18vPPlrukPof4Bhgaq14ZXz9oKRIu9NS8Jxr1aIYdbDMY0vBC9VAd6t6
Zu4BTBqkjQyf0O1jWgYc7LbsfGu5rooWIGYXiNGbwJv1Z791efLA+PH3AKUvu8dVnGjP1qdNsdCs
2LsouTdbsQg+Y4yenJSCub+OIIgkMK9Z1b0c30Dcg72DLtoraMqON+hRKKTHpr021IHHzpBRdBS0
NE+K52JUO6dR751wgFt0zagVsvnpWxkRG9ipEMUO0Ud+UUyakqtibuuTpwwJ1ghQYqdTQbaFlHWG
fu642HWtzf9nCRkqAYZ4r96mRQsvtszeqn+f8PJmHn+AJVeFwSLhJYHv7FwqGbCkwYlDmmOSAxal
9akaT4+m6uimmBNk1pI9MWcXD41zm9jNmGESqw8wNbNA65o4Kp6q1BUtl+5tl+gLf7Q/cCtNZ4t8
+jrPpbC7xYP8hGAIx/McSpAPhABKeL1mMcuqS519XSD2Lvap6ciZk0sdPcERyDbJszXTxegX8Fzt
K65Auj3IsLjA7xvs0OD24jndUs7zo0mfgCfOW3yeiea2dnXXsPqct97y7lvRdd+knGKxM39S3UG6
NWpeO6DuQcfKTJ3CBZQi8Wu+7+MjQj++fp+9kFAhNz9DcjXHVmn1vyjxOXW8RR1JIJWghuxpDdJZ
fHbYTozv4W4qTp3CSLFkHhv0SvkoisRJJOM1zmAVXYppHdUyNjKsiLbOu3D/aQVszCl2J0jFTFtN
lulHaYBRwdSXJXTOmciftZg6EwIMVkGCUgn9M1ICP+9PMWtgKEbp8FDUjiKJMZ1eJzjEBI+5EJcH
Fl/F1ZX3YmzQFP921iERB7ZezQGUNliiolUVOoi13O+ZT1FF4CK/mQMUe/zlt8gJcjM9/waq8aTr
vQpYdvM/LowvFluyGp37u/QYxTfq+7NNF+oQ1ZNbi/Rf1utALaw7wlTImKdxAMun7bdWVoA/if4S
cUfv1JmseLXLJqnKK4EO4KOSgurVauX2cQd3L6r3d9QXLK4lBxZwpvS8G5yZY1bzK1eRMXNQjvie
tHxw3bEHTyc9KKH5krdmGRwYJ3OQYT4BOPewwEbC/vu8KJKXKRKctssB4XqP1rdlf6oRXZubDl/w
/Jpcjgi4hcht40f9QdWKoPNZe+I7nGtU9LrlbdKVzv/8h0uV8LtTTf8vphN3m6jMcSQZW37VRoCT
9JeHTLUOjU08m0zeXw3bGrsmikCa0ql1OttnUY7S36bu7/KAHMQpWbONeXhlmkeqU0m2iQXH/CDS
YD3vWH0cYIM0R+Riqb0IvwcyD3ZdbDIDy9lxSzPjX4z3+h0q2neyiUGBP08lKs8LsZRawca3kfJW
bv6800WflnXvMUjbALs3tX5+QaWPf1/Vn4uEPncve2MRa28VFatXs60Q4gGObMzRzSY2RjbAfL8i
lJzLJ2xUWJmfCOyv5i+qrx3gusMWEpOyXzVhVsfxErYHZtlELGq17fFK4c536X3GYR4ZTmT9fhfj
rbCMsZYSquuUgdju2peLRIeYtyhlbNCXuDNUPsbJys3ktwjrtgj9x0QeJaWqtw9xa8pZmE01l0aE
uZcuzAhY1HfAWgsCFYgcx9FzIqxyssKSH9V1VjZgqlB8jmvCP8+bHHnXO2XDYwQygPKP6MKmqcQu
FK0Zg7hhyEdaM8hPxYQjBiyQDyfit0GaupczeR1ZtZot8iQh7J4PF3TtpjjjI2jCMfNDeYOy+zK6
A8Uwz++Vnvr2J5tfB2UZJ9PlC4nJgBTEb6q/Ktb6RwsVkowwulCxzf1rn78uzlSr7a9wgmdE/SHQ
wSwvrVOVhwh5wLvIMn9toRMudDsb9a27MuK40hGZSYhEP0GUPgPYm+WXK13SGQhBE/QGO6hH1SJ5
52VNUuYJ26MK4BYpLiOgporj+BRLl3rhFa5TItk330uaYhdfr7MCXWmvJt8Kw8NwAoWx6Bn2pQAF
aqqlA2q1eGjcT+gIOSET+GwyPyK5LgoA0Ox1LYbRIcl6xOejsglb4Xiq+Lvv6YnenTHKfRkn7zub
oX0kdqD+Y93FlB1NQztCS/35KadlCn9q27BeGtlphJURLgqQx2N3vRTZ8AAWrHqBY/hiAUx7wr+V
E2j8IRseULF86vyrFRyLiU0PHD0hP3b5o5HPbHG2Q/HYzdGS0qKEAxsbGV5cwrngqxA9VCRsatHy
tL3ycP6/p6ah/CQRrpYcjNXXxhgVuU1lXf8YFFnxLxGGstSlyhoyB/QpZPCGbFF2U34R4ODNzQc4
W1Jk5J8xefMbXiaY1MVWB8M/ljAAMfMnfmXE6C5MtayceELkgdOzaQvs/aBK+IHhLCM9qyn4GgAI
0obJ6QH3QyDsehD1oIQ37RaizIskn+UdbKLU7FyqP1MvREPngcHX9VnN1PjgNM6PF/AHnmBu6yNn
0Rt0N0x+Bhwk8oEiMWQY+OxXiH8wML4/gGHAAMkyi34LYFlO267KW/6jkoFvTLyGvi8sxP4fo2y+
3Pt4mISgBKKiYBJL2m9etcKI+7oIIhuuX9//TCS03w1Cpio3wqUz4OvvHzx1c7w1x7cyb/PRV03+
NYlY5CAMIvJqb5IJi5Pf9mvsDZntOpOk9f0SlC7f5nX3u6Dmpp14qt2zQ1GuLkvBbyxBxkQ5BjrL
5W+KUR3dHD4K/oL3NV9bhE2innGiccfP65dhvvmkJpbh5n4TRMXPmQUmGSQKG3inc6JsP8CF2810
frmWDWze2E2fscT//BuY6VL7nvjV5bhrkWmt/cteWQsPSQZu1rsiv2ndAM48f6WFYiodpIKeHQpx
u291x0QQG63g8c8mFPRph27Fu0mtktxHcS48ZHSNaohJciLWTSxb2e6ynG2csVxLOCBnPd6Irkr5
09u26yfGyfisWVk4TsMZJa6pz46K/TvRq1RsiRAQPccfgIn3orLDbosO5grJ5YB4zwYnLg1Ryjhj
mhtGHmJcxB8cErndbOENFeuiPXwlRxOLrwFQa0x1VjN+VXiEviaJj+EqTHvrqsOnujWK+2d5QbYQ
7kINwoqaFSnPyDOae6gvdJ9aW+ZeXOx3gM9e4GehHnuQsbxe63H6epseOOMgjZuLFBsJ5AqFk+iL
LSsN3hyvDa1NwFLP/qKMIYeuaYGs+A28JAoe7BoIcGZvIEGFCC2d0g4Fjx+qKjNfdje3y0dOj9XH
5xzyLcF+6ZWH0xWSFs+VfK/HWmgcQrqNgolhagni8OqaJidNmWucPeaYeFEx/WzlTNMk7qhUpAa6
XHB0Z68QCqEvKP7CYMlELHMnPGSW/wizok35q6zXb3XLyIMy0hxIcpuaJmS4Cf914SrpIqOx5k0I
kPCppgZqSjDYxKQg79/R2cX8Oy+pBDWAhhLHxo0LPNFCmbD9SVEc7elht/vz8WWvN6mxxVI2jnFl
6zRLTCZKAV+ybPADN9n3jSnW7g8ZttCJ5dktmGZiTO5ZwFkxkpRGyjVIVFStR3IJNMdYiJKXBtT1
WaklE8CAIexaiEQBqJgLdPKpBeXrfKk6TdaHM4T1WHMumBeqno/xlNqddKa2xk0qL5yY5KucvyBS
1LLcKi9oUnNWTG9OKtYdWihwl9nlDxzRR7fMNI3h21KZYzrTL8q6YUP3ZAWjG5S9Jwa35X1/3e3T
P6rv2l1gWAd5MUei/eQXsB15n3cPUwxpv5k+46ibsWs9TySAvzPENyWThj0o64rIg96Miw9LrJ5c
ixs+l8P/NvdX5fWCoo5Ok+bb0dvEQH6iYElyWlG/D9Jjc6ng1XWV+1GaSoMuIAFjxgeSAmaxvFGU
gszxHPfuQw8TaIXsyZAh90jvR5XVDxftQcGl7DkNrCPArWVKVJhetLf1Hu7tHeaPETsCba7qhBgu
aIQSMAxQ8IhKW24jny4YYP0/yPPQrko95H7/D0VB9dHOxm4AGcKGGKXjs5XbHNSI0wwvcJ+t2aU+
Vrjs8/y+8JITxPtNQgMi9QHIqrx46sz+XwIql8GoHyvMEiFE4F8x/cTe9daVnJOUKZstzYMqMUUq
JoOis4UoH9dSSKp1+KFEPiTZ0BrzNd6wBxcxxo2sTyRuyu1zx/z7AyhkboULRQFxrxz0A4NcqMs3
6la0ML2IBhtjtG/NjOYw/96ID41cbM0eJY4T4/6+jHZegOA7cYKzYpca1d/JgVHOrkDhC9xcAKUA
HrdWZkxpu+9BuR7uJxe6jaelSRA9DRcL2461f9KPfrAM8gEVCfxDt+4zSJ5C0cC754XeZfDtfqC0
9H6Zc/djDIIdVpEAO9K0sGxyOlTxs0vv1AES8rIFrkjeiJi3NUd65nAHKO8e3/nHd82r/Y/PCirp
45s0JiGBkuEKt113n93+SCOnk3iGeIJQs8MHyU4KA0KsUzurSwMZaotnwG4psEeG5996NhkGE07T
d6XJCWZnDPXwPcHUydlzFnjeh+KZtI97QfHDLii9b12dBSRzCAhD7n0DUgds4JYmE7yYYODQIlti
SczS/pP9pcvTag6PoSaLFPC7OFN0A5/uVhdyI6q5t1pgYx2Bm/QDKRtg+Fm/3x6v+2tdUhZCrPHD
IUle9rJMrWkg/wQtMKo9WRO1MQ190bCt0YGKDfbCWfTXTTDiFkVaT7iqMtoPabZ4kDX6Ut9C4dYT
uewY95ePPy8/FdJuAhAcjMkKx+BtC7ECcXOXtXZiSYq1UYpd+X0JzXETyx+hr3pUa3BlSAAJwtLU
0mNBOZ98OjNM6+LP3YFXGUeAAw4afbsqHlSaJpyg3EaSfYvdNe4uGTTgrG3T8iJ849hYsZAsmiQD
oxYdkNnPqnyBtSNcNGQDNcGTYmvimlRh9c10QINoKRwsaN8ronPjlK2TVgiD8u0xSN2EMVZ/VNkJ
lI2PNCXiLB8I4nru3RE/3kqByYL5pECTDCb+8twdFGGW0fOMSDeMCkbS20Mp1mPFtN86Erxf9FeW
BfUCJMo2sS69fiDRMVFlnKG6MnUX6Rb2whbIfFUANrxFuJxWN9koeQM7T7YEzO83dxdTys4IOp+S
Gz2uzzvAPYPpEFSkq2sIPL22W5ZmzZsybVu75rpBgt1cIAWRnCik3ZZVdH0r5EytMk6UJfdFFNnQ
ms8o8zXvx97CV7JykraOEXBTjQyWA5dA+DgiRa/bwC5UTlEdJq56wtR0uWBFnQAf2y0+jDkhHlq3
OtTjD8m8rIU8XZlo27xvag1i8PwGO95sO4Qzlnhp1N0kNlvZdijcf2TjU1XNBF9Ul2+927YTOhTz
3zSM3wQokiC6M8ft0Yl+TdCgG9vt840v+1K0I8JsACqBKGzsNq0cOeDVK+JcqJrAZcKGSFJdMh7B
++QNmThlWChLAK9X0FlCStSuO9FI0DzqzFFZuZEMuiimi8Fqt5C5isaw0P0GFrJ2b+8+K2gGojNu
BPbMNgzo1a7POxC/Z++RLdGjQLVPx3L0bjBFxFVoXycBwN3BwS0JDtTa2/9PyFxH00QkHsXgKbjH
UV3VgDwKDOZTBsQ/ICLWntD3gKwHYrXetS5qUYuDrPl9IiwI/F9ApUbyd1V3QIy0OrpDUyHgDBOD
LIIDpSOy+TPF9kxQ6sV9tbEhXVzwtQHsa+O8aOdekmjCO3varzUJ4tkNLLQTHlrCyBOsOzLkisEp
K8jQLWrDFggPuOrFC9yp4prHkYIkgRfvrc+D1uJ4crXEKzoj8h5JazhaxnGhpD6KCImfDMKypxYH
Ug/sGovK8lQ549Ssk2BwRF2DMjAt2vGVqYv2kzRRDI6G0+JC3EWIuwO8VgX/Gj7xwCktajqiWWkE
9Scyc7pVsHQ7rE+bFYYLKwnmkAzLhwbIMzs+Ax4Ers22Xa2yeWTjPSo+clFzOJKPYspfWHFTuPu8
3ongAYHP/LjHHSrGqmcBjbCR30+B3uDuo/m2nldObS/48Q5T4rUljzXVUhSsD5XsLV1XrA2E6u/t
tjWH2rWtygOJ3hAuij2IEb11nrqp1Ye28ZFWI1CeI43J0wssL2+YfIqd6GtrbW9y/PLFu2J6nFma
tZxt3TUR1U2d3qZFWRB54mxBaXu9RLtyatg+OMZJhzs6nTlYMXBRoS+5TZh8NAPR0dQBcC+loFNt
outk3GHLC0+okXOo3biDwyQuhQf5iuJ/xQTDgx4kDE8VqK9ms1pc10gK3alnpNn4myclOVkdkSrG
ut5RN5lzValCInKedlLdhyG+1uPeVmZuGVsmVHwd/lWkNPCkCYl2LB+tx8xkaWRuOk0Ose0JKHe/
OkXAd9sgtS+9Mm9xD8lSJF/wQtCO3Ik6TFnv60RkrBK/Sywg80TemSSzdF+2CVOqvuTPFb6vm64z
nUd4Ri6Qs3DW2Ms3OcHOYQERxDm0ACj9xiFm8bAHYWZVgplvPsrxCqDM0atBeCgH6zIsT5CIsbK+
ussG1jRK0sAbFly6Xe6Dc9hYSTjSNnJhP7UXYBX1ADjPkdPIfIG6uTpbvk0r6QpBmCkbPSZvMQk2
wdTbwPCftql1PbtJwQEOlyAN4W/K9gNCZEXtCy4EDcvB8sUns3sFDO4G1azbaUOxfyeN37immNvy
bF2pAbsgYymgUVw5/41a1bnLvcVapsMoAIE/7LUE5ESsg9PpBggJVoZZnqtNDScbmwkafLcraQAc
al+kkvEaVDBIsxjixfg2FhiAUh+Hs7Ht+xftI94LuUr/eAA9hLe9x+pMLgo0p06/JrNw5vzQrk7K
JVXuP6G/YsgYKuWKOe42fJK8rjGjKC4V5jUE8TqS+amjV9ehG9PWpvrvN80EROa+KtcAMvr/F7J4
LQiVnty+AacAAtXmfATxZBuC3zkG+J4MOSuZehIsHglM8JFfBMkalBG4K69q4Uv7AUDZ8yKKeLe9
sJWmv/PMA+3onAqG912c68LW8D2wqW+r0YGJkY1TqpsEZC2jwyjaf6/cgjzW/NdBXFu7EuLylqBa
UEzDxigYRy8kTAgilnNE/Qb0JAYIezcyHVDJivJnjiClFwtDMeLSrRlY0S0Y2OMPUvI+wVLLGbUj
uKwM7RW4tq3gyGaI87Yk58JhGyKvksPwD2SKL0yRVTdmjFPTnldv56Tdqu4zlOlT+K17RE5OD7xp
K4BZHqlrg3ogFD6U5j/v0LN2w0uqYmmFhpDf37+8PhvkDBYqI2rt3tdSZMIeMjm4jc47PHOBK2rE
hjjt9bHtro7C2NgTxF2S5q8Bc1SpnMhLIRHctukSFjwGxuZyuwZcz5LUrBeVkNQExseqrEvw3v/c
RDBypAGhqZk0xBb37yA4icJl5l4og1EnsakRK9hZXqa4qN0b2HkZIcguBJhWt//dVJiM+mJwftle
yDXyA+YHf/7BX0Qj+IRENY2+6b4lPFaQlf/t8Pe49J9yUl+vbAyZpNN+jHFlwXq4uBOEAhBxNJq2
xFtnQQAMvhzYTLEA1U8kM+UL95Z+wsUbsOxHo0UJDMRazB9qghLsx0dG8jUNKebUkITuHf7AYKOe
XldwOlxDPTaSQavr1JEMQt/1Pl4G6r+aFZ+Q5F2xp0tDEa9pTgH6u8O5o7xAoBQOEHpqCxB0noO9
2QL1b01MWexkbvu/GiW+MwjWIGhonb0cYDngU6/RXWZkmpOGffH+0UXK7JEvcVUCRkm1nXmRTziI
OZeBRtbD0hv4qGs0Zn5MfUVNkxF2yA4s3ETlAT/hxgi31WuzA/ji6SeyYL+nO8bTZ78E+aAhzxkP
O3OaO2tPmn4696ojG5Xr1CsoE0QgOnRJtbHQ/T/Vgsrf5NuWH+79qZueYJFbmdkYkgIXieLdETXm
ri61U0yYpgU7mR0k1dg3vzfgWo2SDHvdVRdM3BQqjrmpOHhvTSLs7JC293uAW2b55jyq/oalNTjk
7bV4UiKuHlwxghqMv1uY6aMZDW4FBMK4XGY7+s1xZoWYxSkCxs2ikivKOj6yczuiSBxJVyFFfN3o
gLTFFxgCV5cOyIk3WM4Q2Lef5//NgNpt7kViqs4j2PrIUKFTH5tqM2eE578gnKt4iq5Mr2dkdRvM
GVXR5yi/fgzeMlhSC8zMnvbOP+05SuvgBFLZvdERZD9sqbjkCF1PtrUZQgCErN8K+7sBRDjGzEvx
VSYvZMeu8sLL3xpZ1WXwY4HcXCfChDmAW1cInFMhCHzBNrw6iHOoV8ipLzayANDBmzkfnyZbd/pt
nqMe78KRStLbrEPFj69/bBN45GuET2bcHa4JDSnB5yg9VdMDL0uBjIvPfgZedF5/5kAxr94Rezuf
z1RlRMVQ5iUrOXorVjwV8cgtRkknjCmcvJqS8t+wTcwZ7L+RXIYLjsMCV1r4KkQqUJ5t7aT9h3+n
cRcsd75vzw972Jw52vVHtqt3+elm4aI2P1CqBD+aehRdujRiC2NGuYeEYpD8qgalQFXTgnPSe5V/
+cMT5PsZktS/6FtkIbcFyblIGDmEzF/qRgJcYacgJo/VhDHe48UFtmtN0PPQn+vAavUOxixVOMR2
CbezfH/s8XG1FsN58IrlXtnxabJh7e7X/XJvCkeXDmfewYRn0sYSln3AIEBdnoYcRp/xqWDERXUp
Q9deZCxKcsSxwuv5MsJyaoXyz/ECjwL0vbPVZYX3uy39lUizmdfBYAYEePPlVNHy+6akS+d3nh38
qCvKm7UKd55UZbOj5A/a9X1DnDZwQ57vfHorw3E7VpXmIbxQ51eIriR7rLEW1dt4hglhKrHu07ZG
Xj2pDLNYKNon2l1gmHE4DGF+nT9FbMB+fLKuAg2tpV5Dm2LZRlz7vKhf91J67otrGgW/cu4WMFce
y43L3+WqZEF8KsAZ25lJ87iKPrk9v3jqINSucYHDJkYUN881MzF5xaDFuUxvN72YGKSfZm8fxEYQ
S3PoPJoxcc8G7TgHJ7F1gkTx079mJM6zjIady1BIMmkKl3l0MoGn8wPo6/2YyvaQC2Q6wpcfWMYc
5OhdxPsGD0AlhutFt6efF0aUO8kI5hd41G7/QB5cAi2VYwLnLHFcmMxGrB83AXvRBOAj6LjF4CPd
45ibUD6vUB9HGSd8ojD7JZVEvW/gdG5hZIFZwqg4i8g14feP7Wh5m0waF92lcIREzPq/nZacDiIZ
RX+02QI4MNLXbNpQNTxQ5ii2GFk2WJLTaUjSgtLAxgBXK38uaKGiwSfcNAl+oip5+OKkUtQgQW+O
cWlh9lVUWxqJ2BnVL72w30Yg4p7zz7pz3un/7fGacxnMPC1YPoUNygRfVMKMIswWs5xvJ4gL6hv3
bOhFxPdzqSk44LbmyMv2JQ8Y9CvGn3yKFbjFxRNEb5SPOLDwInUnAIxjTSmHY0R8DO81NsgQdMpP
VjgPT4MwEFzD2A2hSzLxypVHMqEyutkGEWXydcKX48ShrRm3wprUZs9JtfDL4m/dlq/kck0vkJ94
Xy77AETu9U1Y4h2nMQm3kCEtPd7G3oK2zgZ1NuCtUASLVsidGHtVPZRBIiWmon6/MWdLZ9442knW
lxPkKkvhOyiujF0oQBXYj7nzWerfRhjN5OKTt4+ovPBZo9xQ7I4M+77A0CC2EwI8e//M2twhyMkQ
Pnn0yUjdv00mZEQZOPqwGsMexuK6DCTuvHuhdNvIUZSksg4pWqjSAOapqPneHgYU/dgjnPEWQtlR
wkkT9bdWpqSICQhVCtjI2AMVe2qaOFG7PC4fVOyMueU91PaqJiA+4ByqnKWSb7Ik/0KQxfgDTfVn
bdurQb3LVUqukoQHTYb3dywVRgQqXPnMV62wkuNOCY8hVZaN7Le6D1CptwqQL6zBno1kI/kmcoe1
Zn/XICUpgM3m/GrkmjKrLimNnIDzHAzJ2otNgafKKjgqC1LDst58sNPTbMCQamdntk2k+rFTvNZ0
yyNog//yKYqSO9dLq6sOvAxyNHqXYQU2H34j63XNuB7zfG0T4HGTWFju6D/n+aw/NwrEACDsOcHR
oYQkWYFPu69d+8n5V87lR2E+TNw58WKPIPsursUrofkkNZtOlGblNT+MPNgWa8h9ruWiBrlS9ikN
5wR9pWzzjVWWxc2I37S+mE7EENTMjdc0mktsNXISW8BaE3tQfC0IlMPLfZckn2re/u5hmha+h/BV
HvsMFMkchaYl/Pvt6msotptdgAeRwrItOIRRireq1cXyPU0PJd/Mfhjg+szkTAV1GLjg4DZ9D5nc
2QZdKrjBgHSLt7bYcZ6MwuQS6JSk7kQbnyjbGyDYvdLbMfRvQnHRDzGINzWtvHFQk3C4kdxmzkZU
dNo4J550qJCJc+YARPLbA33hzkHUpe2OOZo54itTxWd1z/DpzBxnYzOT/VQyAdmMkBJgEjmTWdWK
4O3iwWNJ9j185RqC85sDULB1bvqnYsU2Y/2LVAHsYdwbzzQRUKcLW9UqI3mNonblBdke/ArWxd2e
75Fr35/deyk9I2VPE02TrWgGm9QN+BEl6q8EEvHj1bmA0DtR7fUJN+WBf5wd5CEoQQCzHv2Jbnpi
9V3zBtErTVwachXCoeKxK1zPXvBy+QvC2opJHD/qi7eKKk5cHw/prGM3Q9SpKFDLQNKMnQmhoLms
xU1GQTEn0N8lNYiVO/7HEZCosl6J2t4hAhARQsspSIjx4Ton2S61nA3Tz8oSFn/VACoFJsZF4jtT
vl2ZQn9bHp6U6SGkIEFTglfr0wtqaqzz0E8rBp8IPUZ6BW4SYDKdNZYsoy6WBrDkStFyBzKt60Vi
BrlqT9GpvtfIMdh7wJgsJGIRhJndFfxc8wEfIz7ruEncBU5+jQNbfpryClpjozseIKMBG3d+1g5f
7mXVGJ715jsPgvOGuHtJXiein4UP5O5icOAYuxJ2vx59ZJ0g2jOPkV3nx364+/srYrzkBCiZxhxY
9PQ8rvhMqoTHluiAvo0dyAFg95eRm11OVW+h1eTWKoNaa6jRLmPM13zmSruRQ6mVj6hQTyviI2BW
tpkD9zR0xMYOIQZ/tSjb8R3Mtjugu2rAtbVKWCIJ5VGv3BqFN4VpsRvcqexftoyjS5fyduN5JCq7
5qzmVaPORIE/hZDl5A7abPlT3wqjI9DveWZTKUW2gSAcbtrSm11FIWG0J5GViRKadTxgZZoFLIPX
BX+HZs8h0F344TkjdM3pr+ywGwDq/F4/l8qsJZc3kmq2d/7C4c6RTB0+OwYO9t3BfGiUNsEFBili
reEeKC52ED5dfrgW7ZS6OX9/DvUl5iYYGFCQKkBj2nhIfTQSFtEoIYnBMQ6/K7MQJ9x5Re1kVBMN
C3+BVyBKh2tMWlWeLlGsiK1aYJikz60vbCgaGs2kRANAwCpkFDhgLik6cZpM7EXNDd1IitQODuQU
xlYpC9OgugZ9cL1X2ZsmDuJX03CraVIYDHICeF28vQFoek36OW0Zk0KjUqb0NvEDWLYGrUvayGxy
fyO3Z2WayTk14wzlyt9SyJuyk55dJd7GKP/OCs+YjDMY+tlXYslXLZaC5lmy08d+bjgUR96by8qx
9zzjPQ+loKzBSy8TXR9+ToOI0uNaIacGxwggPmeHxMW8viR6JbL66hb+r19rqXgoN+8mJ3k+Trr0
0DJocFQGQZRpOgq0FFtRoP63rqI1wrDFxksevMIGluPcz6cce8Ca5d+6lhjBPysVGQxUMc8mdKs/
B6SdTIaXL2okNSEQi0S/BRUxDvNnR6uxwgpLIQEf5/iBML/NCL6imCj8GbIhF101ARirUj7L5eUl
a8IqDEYVjRUcYA7Ha0dKH/H4Iv5vsN4fFAVSggVFOlVBpX+Rg6eFXBNB3X6rw/CbrqvIQglsqOW8
yIanhAnL/d8Bn73gR+ebES2qn3MROnWhElq2A9RUEeVE5OMDtfHIyew2I9Ao1G3LL7/6b5F4p+6D
OoOfWhJQfvQnRy1ToTZRVvP+GI74LnxxIw8z+Rh0I3ejsJbtVANM/CQEdvqysD0VgmayUHETVZX1
+cH6J0M6gek3/OI6JyIqpX9je3VeOhAPeENxco3hMYIzb5YfIUUNSPDZaj+m2G+hJTdPn/FCILzP
iESCv4qCn4ehns9zPcJNyLhCoREUa0VJ6XyjahNsR1THcKp43Vd/mhckR+KWPz1SJoh0kDgQ94At
iPKbvkVkGJr87voZFFrF1yMzuaO8+47GvDJnlhab3dDhJQlOjn0dg0/HvmBhcLiq7LH6ATUCQCrN
WjppfiZ25ALYyJRFKZXIOIRL0nBWom04U0xBa0EU8MK8/FuIdPz0s58uMkG8hM80aKRq5PTzXYjJ
7XrawgKDjdrZJYfMQZ7YHmAor7DTKrgG3ZoHgRaZDmlAzLpFNAhS/4oLwmZxp7i8zw2hi7Qab+8A
OWxiO5RUQmZsRsz7ycNs7snEIPeBcKUT3RacgSYwTOVVNb63g+eKfP9u5h1qrR6BCKKmpiMyoaqa
pFW/PuClE02+tCDBvYAArZbgEn0VLl3N+TsVMwgJxDB00rhKW2U1UahFIWbHFmrz75QS8RJc8vEh
qCOXdM4NHAvwavDlVFC81OziSPbEH9nOgVjKoLqXnGabKrf+OnyPDAq3Bm/lAKccLKQxa/Pdx27m
BaYThK3azcrTYXMx6huBlbZn1Do0296GqRwzAE2XHww+7TzAZscDeASlqw4WYN1Iu/Jg4O6uISW2
eL6yCCN58L/KxgfHQbak642tetAuoGF3c9vujfvc0FvNxOrV7WBPsO+w0fjc0NsfpRtsJBbKEPSJ
oNFizgQOdu9jDWhXY+nv3UiAmoxRQglSwESk6TGPYqPLxyJEvFZai19Prws2vxS8SsHexRBDdD3f
f4UQ1fiNxztanOui0X/CkHqbUmdA41IRF2b3NjGNzzl9oGuFjFkPxgTaNvn8ZBvlBjN5OTRDMokL
6CJiT5k+8qjzWijv6q9vLcJ789tY+hNs3zkYkfgCFSOOFkPXM3NAao03POMGMOiHC0MZFbbHk7au
UtHT+2fJ6qbjwaDFLSeSi+32FAfayZ94sSaWb75rz76hib+wkRvJZ4+7ckVJvsoYjADdytjYhKut
RaFoHSlUn1mJlLnjZRcpS9420MxXsTl1Z31Urx+w4slAoaJ8NvJdIAn0yBa2C6xwXt/pfNWZgAbf
BRbN5+H7e4MimAMkJllHj6zm8rU38tkyy5wMnvlcY8K7XZbUkQBhyKMrMPRvHdLMy7LPw34es4U/
/jAO2fLxu5NwCQJ6Xqxie6fKdjNVJX/dfbjVXYl3t1hZbpY/YTw9JI7Lol/ny+AHRqXKNMjOw7Ik
3sFYsG/KX2um7f3KtNpQWotmX/i48bL2szHZTYHP4ryBlmn/gqUSFh45Ov9jc0zyw0MmaHM79CJv
IP5iQoZbpIWCsCZMP/Qn/cjHFd1B4RePRcUNwBtssoC++SCYExb6QongX/T3oCzsSPZSAlynbfzB
zhvHsalDlVCsFtSFaryMvLbQteRwwdZSLJy0K/23EX+niYJolEPOIVW1TgTMiCfaS4TWq6uz7mmH
5paXzE1FLJ3MnN1Hs1jkEFnw+YYt8Zwtf8atbQ+LzUrOP8p11bJmgLzdgfHsLv6+GyFIW+JMrwSi
EABHtXP+hYcL0MkUziSGv2eW4oNYzi+G0JKRsN83pT+CsVQ1kq5b/UqrYbgefuM2xAL8Oo2dxeNI
OclSzw7fkLZ6KOGU1EkWAwqs/8NTAcqSEUSbs4hnM6ydkR5ZbE57i3fROt+nPz6SAkuKUwaMqsVB
5Qm/QFZbF+kk7fJFx5zTekSzfXUdT1ss5eWPUKjjR/w5+im37otnmNLy6jwtjKA5pqIBOyNLGWXn
XqfeSWmwxe3bzrqjSu3FfinW8A+g/Ncf8g8jVNwrqguIDesb+REjwpIbrC9ZrvT6Qj5Gp16RIwp+
QDdFLsKke/eY7XYj9b2NKWIDXH5yaPsY1yUfPPi8FdqkvjK8hSL8Ajl2sbTpk4cS29tGbU+k4hM2
OpUmhyO8I8Sz9L1EIut7Ek1A6i7XzUNdO60p7DrFmkQqC/kGpDZkd+B2XMyJmsTBTBxoarZMShO/
gAvwj49gCtuhcIVETGgPloXCdpwenMudsTLdW/0sij2uXpwS70q9gXVdN324wcvPr9mO7AMjV9P0
A+/u2kn11ToqcQ8fzkbH0oxWt7qQiuChyjYp4p3BgYfOR685PYDxI4ub9E9qyez9P+kfY7rQMR2U
+d/S4rwczFN/tn9DTDtWLQuSxVLm0oFt06UQJkBd4tTiB5rx1bikZ1kpGNkl5e2F5+sEXwwYlkWP
7umdwX3nbKd3EFc+zApOnef6AoENu2Fejm8kxPK4e5T++Dpup3v0mt6WOa9NEqBlkvYXnXPIMBpa
OhjPKDf7aqaw7YElW4jqSNuROGBF7+mEgEZXwSRTMZjfSuEL2BxlND3vwbrRstiFfBQInVeRxvTR
doqFlNYR5DkQlv+ettGZzMME2RVVUwVlSmLVyWAQhWGR+HiyXS/6YKn0NvFoyJ+PiABtm1hDaHoc
rdi9ZUcCaOwsvNPBFCZKsh8pUaDU82UsXCzZkyEj34MFwnKhmi/Ww64Mfq460W4/F+jiJy77tVvI
YxxujRj8jZbHGoGZ468wR3elwRNfHxCxsWRTkC+dJlvSA4wCdz+QtVmT0GmW2CEr0AOCi1sTZXAe
2xLxdD3f80wHJhZW3exQ50/xgQ70Yw/N9AdwzuBkdCxZ6pvMPZCsS1cKkjeODEby9vZVirKCBztq
i8qtXFk0YvlcTyFIY+6MVvwuzTntJhZGdRRXK92toG1/03UaA+EPFZaBWPa7sI2JPaTyBTlWjjoP
oStnHv88OaeahppQf2kct/uDyxH5bnVrwYltjYhnZAQdY1GxIv9T6mA9SGOfrpeRSYZoE4Upp+6L
FyZd7hwK8o4uJFaQcuZj4HskkqCTLDhfneSPPq4I6b92SjWwb3Aox1RIJE+7FthgGMo82ccN/4ax
L7/ZPQKh0f5Gj6WL2d5Co9b9WPEBGqkhCS6bKITaB2JMmmQXV4U1JLkQ5QmrzklMqrRWlKVzMJr6
dceEg7hdlCPm4J+qHUAgZmDvEc5Jlbs84PGDmWTUgOiJbA5L+gMdzfAiAQYXoexDJvZUjdOd87FF
wHOezvHl+upgzy2vurSihHHTwuZ3rq2aVoC5rOwuyIPd01k3UlvAEvJeCD+OauWN+DP+gOHPd+hI
x1jsjR5cv/A0CZYnJvwx3Guco12lh2cOCXKHiibSwoPabGxP+QdRvvnuByMqi6HOESbpc9dy+kif
DL+wYDIwNDje0ZjpssusuIkSvlmgNmeTwFaPJcmN+Gts0kJKejJIda+GG4U+LkPxyiT0f+M+rAs4
pmUmmO7JGIx+86dvI9bZFMuQ5HrJ4x4nBrKG17Dw6jKH7veESVFOx1Jr2T2wQ0IXQxgsxCkRkQoL
yBtFLWnbQ9e/MyR3fcAFAtNwHfhhrZ5HFMo737ogbpReW6aQY+NpAd9EraSSPq/zblLwCFT82CqT
ZFFnYC7DEaxHJrTyzIJ4kZm7gqvfbWekZVvxWjf1S5Fg5NM3pkj3tRmFtGNHSaHUufe3DrYZuZ7p
U3Y85x1mkz1yOKnU7J5mmCjk4web/DX1XZFLfY3mp3+iLcNMoLbo8zeH2ZbVxt+nHWgVkm1lX9eJ
CyOM2wgICbcUBKzOzYGjPJ5Ab2HJpyQKffnPnlgNsowAJId5hugL8L8jWU66WuXzfqMbPP00p3iC
V5hSw9A8cWNp3VaiCRFtNOZ/zotIKL16OOwfRA2i23WDdYlUMHmZttSSW1mQ729WmCqc3LEW3IE7
l4EyBDLuIExjDacBmXvKS7fW5kKzjb86H3WlVKIw28TFu5wy52svow9tLK/EZbNskVb0Sm+JCPbq
vRVngkJN9qUTmzh2oH+gOEML/kvd4tYL96F94NB2HbcLEXC4qlZOLHwy0cA+vp4qhK5fIiCVqj9o
QbtalDbBYQoZlTMJ5y/7K7T8GGKzSUchqA2RBKlkBxdmih6X5gUS8F9HpmdUnoA6YvxfLr8NHLjx
/yWfFs72/kWdtllAhdLjCUDVkfvWihL144M6vzvV0HUSEkvR/0ZVDiNHjt+I/PgsMZxObYRE8Y8k
yrcqphBxgOiNLtvemKbL7o1fhJevo+akBWaJlLx5iniPgB8F2CHjiE0C2Urt/Q7wVMNeP1v3APDu
BMJi3cCOJVyltNLs4F43qAH3I+iLwaYnOibywG/Rl5nH2oRTjwZQM/dHmhC9PpQVCJQ86k1/TLJz
nlQeGqGLhZ2DNc+V6o7fgq+sifmVg/eptT1Uj0u5PDkVyhBSQ8ZX0PRjlXb195IlTI9CJ6OKAYyG
JBcvjd1x287SL/Ub2+CEzm7Uw0j3RL++zfR2TRCoiX4FApYd/6cpu/6lq/iI35j7+7e41zc8pyUl
cObuctzS528FkbDXnkQEThB7TH8IRyBzM/VJboNMRSgaTiZTBOOzB+yEeqF2MKpRmKXiqMOyVB/a
4nOlugm9yjmo/BzT1fromNNlGcPWf120G8COoBi+FafLHi5PVHyJFo1/xc7nDZGzdAqLVrRq5QFh
namPf8y8VwuNwl/pgb94p0x6W+JuxaAfdX/MN+TMXX0DR/EmDv8jFCTwUX6nSD+x87eFNJB8xmdm
WY9YgtjOnFqdSxFqGEjPOsGGbDeT4lJ81SV2SzfcnGM8DqN0C1mBa+4unxMlbWU8quSPE/GiWCvW
Ux8TIqQvRUy8aP0pC72N0L1a3hKwhBl4dyk2ZuALBiMFML9abdcehpyKqVjg7QRkYRz7xEuq5bbE
AUP4HCgd9Gsd+A5CZ/Yy1CuXdsGOQV8Y9SkyQUOWHhh7eihUpMh9IEeyv2C9/dgAAwDbiJyah4C8
NFtgleGkK1ck/wXTbmlcI64ZLfolpTzqkJn4nR64JkWEo5daoY1F+i663CQcKk9wnUoQL3tKQMud
AZqwjD/YOjF8HRZqDjftzJp65R0CfWoP76s6tYlEG2k5H9tCUsKCZ78+y+cWzbZv34PGrpbEYuh2
Hx74/yfWnrYoTGYXygyJvk2YzQs7t3/iVs6DdAfsx2fPFuFVya1ynm+s8sXefY0/2HPV690C0aqL
nrI9kS85kbYpW4rr6y2QsB7DA0832cAtWCiT238brvCRgO7FAdfy8ScKqmCbhHONP6YC+x26DI+S
18D2TT8OSYYRpxo5J1Oheyab0OLEuHiyJ/tbctBoKz4ew3n2Ya/2/E2uRA4XVCOZry3kPMunzc35
fwDqRJi9SHHSc3G1LY6VVjLwELSy/ZUPMkH2CJ00tLFzZz29P7p4MwgvDCzfuqniyczkaOTah/KJ
sOzEf2k1TtAAbnjeTh7WvnfVfCdChl1pFwnAIcjVGGglLnCLauq1RBTbjR4C5ehoYt0Na0+EGrb2
cK7f6uwdbFJWXHyOwIuEshFUsTZCQeXRsKi/SllXNBUn7l0BeWtphjX+V+6nOAeCq5pbpNfot5M8
NPY+/87SukSC8P2OfnWa3os8/wOISCZt7OAsPEfz3QIUmbSYRzJILzBFLZL771ExjbBAtfmct0CM
HstUk/XPGvnm/8/Z1HesZ4Q/uZgw3GdxkiYWZhNvReecjnBTUK2nAQjg1KEoOA0Y+2Ps9gnZcXoY
zbz0E0WfUz/UxOERlcBel+CXrbHTfxJkacLxcIFgA5bpHgENlc/gUWQQ1xHSZD5EktGGLOcpPPBr
nZtj+uolMa+gG/I8KZHJwuTgtdkvL2CvL/EGIH7/vMcT9unkRNk7C1k1d17mwFhTv7ysb9Jm200f
GADpYdZQjaZYcBzE2vjVIQTo+rKxOoYvyhjTG6mFvdlYhvd7NOYsddonuo74+xxCvuQ6c20OmQnq
Skk+BJmqlUo58JneboI9IXGIynBI6WFE61ViV/OOaEBTjXioobX/7+Lf/I2fDBmKmWbQoP6pu/U3
GBv0p/aDTRnhECceznVIx9eTgqC3+rbkLcjAcYY5oYPn8S2yEs4UhJpJwTOHZ15lg6KN0+FEH5a8
JLaHWTDYNQD8m8A1LIHb11rl3b5isIa0tY7ELPrkL5v5GtXdfGF8LKUhBnHhFZ+HtPm0kSIlG42N
nHDfMxm++/QimssQPfX2Nfz7+yGUDsgvBz5LL2S2+XfkcoDkCIuUpvbPSUPKikBykLKX/4EceJjq
4jgUes2STWXAC6jUUSiY7JgAeLcc5VoUazTDx9j8ESol3480utNW0jgcCe9a/3odbn4fB2ZnG2rO
6Y1U3GPmhACJ2DMYSvyV8TdMasAz4EsDSPeBjm/clfAI4INooJcTAUu6hIVNa0u9kYfrrV6TKhvP
Vhsy2sWyLJHsKmeEkNzDAGXram/szzpK3cePEK+qoEtYWrdiauaeH8guJZUrh+4KvzU/YAdzdLZb
opiQq0dS2644LAfiG3o/hX9Zn2XuL82mSnu6DEbIn5wKHXHTG/0zkp2FctTRWbEwpazI1ABsomMu
aU2HFFO6VpAtK8zGg8j1hru8pSwho1jQJVNTfVkY1kcLUoDghZg6oCALvVNMuH3p3HxiCYbvAqTP
MJ01o7gHVd4ezc49bm726f0MVb4H8V+8vOqKSpdrfE2SQokdju9QScqVlc7UD7THnGp1f9991tIl
w/ELbQ3rCm9fVtvuvIydozRRzS7xgNZ+XTjZjCPv71SQOxYvZOQAJDl81OmFE49m19c4n7UaNM5G
W8vdnShqfbt34pXNY2IFg3JSWUGnTn8e93EdcQAZGCCYLjI/EB8m2a6sG2eXjPB4Q7oAAcT9ueiT
D6SP9VlbspsklxkYIkbHg1lWKgIAgXhObc9CXwsN+ixtm+zvm8X7QwubJYpG7yhK9avva5FsSnw9
Sul+v+fbID13+FeNKNEGbK6FxtEdsfJVtd/9ttb4lotGaV5KE+UXlk4DoSN1eqXagYfrSSucPgOg
I32UxSIogZMGkTLteHVaYU4Dg31kq+YtYK+oC2AL2NXy5JuE/COmwNT+y9XqYPJ6iTPOM5V8sycf
zn55/fxlO9anpawydNHN0RUvof8s0unhWJ5QY4q+yI6T6vmn98HKMNN2njgdxpSGhlhmCx/T0hMj
weCW+QCEzOgQpKm0qfTnCxZZCCg/Cg2yRqaEGu5u2a/Yy/QzX70EnCRovzw3ulVwkmVn+Yv/0bDq
tvIZaDsI1koTiSrTv94wmR3dcBpo5MXVZWqykwElUtnLtZcQuu+nQp9leCZtxVmy2v0zJk87pjx6
hirNWHcA9tyHeNQdBfWWKfkgQfQ6oHMMV+ZJV7x2hhIDKLnl4lt1x0kT+pQ0bpwud64rmL6MVykV
VNcAM12ZRmEWU162thZN7SVPlM3xNJfiTQHXkZMR2FRq/rTGmTHH8rs6AGw3LpP3dJGeANE2PdGU
JR5QiH/RXaQZFaBOR4FD181zailZGv7FXX30pibMEsIgJnSwsHPBXvI3PvnsTaeguYj3ZqWzcMvc
nQuDfv6WKMME3mOfnm0wo+65+GdDwhSSNhMHmD7LBOdNHRsYRqih0uPvRzmpDf1DTyU9Gpc9XJ62
1elAUfjSClS2B7vBAoUONzmJVTrAd2mf4+k7fcj4yXjBMzSgvIaRRzHKO1Yhd3DRbXxABn8dFq8L
yK3503kNLWgzxUVZ7Spp9Bf6Q3XjbE5R9rsm9NaiMlr11TzT6XkcES0pmVpRFJZHonV0UvWEmQRI
ag4fx4UtnfcGd8e/J2efP6lvJTSK6L3Q+i7gx3o8knxjh1uhqc1ccmVtbqYRYHtEyN/aAo6DAMg9
fkmQGFtTMrINmjDCaxmaIb8Y15zlxlRo6H6X7iSAeavCLL+Rxq4xI2pqghr9yrF2eJL38LAA6mDi
Sgg4fFEr90TtQBWxxzRbd1xzYQnlNWQJ/kDfcSDKY3SvouEn7v2ZO5IOTq8C1Po4yEjrfHCu7Sbk
EeCL5BxImW9Fb/mweSnQyOLh1G2Ae6MjSXXhsjJ9HZqQJ1Xg/3O3VEikQLI3/uU09r2jc94/1z75
UeJ6GaJcEzekXOVSyfC6Xwv0JCX+G78oKZ4AT2QkV6edTph+c5GluYC0/DVqqnd5A+fYcHmV2d1m
wGGDS5IxKxsGjvgVSx8S27lxmZ6JyLV1r7jMDe7KHalGSJ0nPK+/vlDjIFiRUMCRZjSC0YwnXMcq
+eNM14gDHjlPiYG9zCH1vthNWP63J8gdKzSG8fsj2B+bk+NS6Q1rK+I+0VmQdtkeIetcQF/JWRj2
jE/QX/1qPOl2XwI2+pbUKECbzniGuXCaIYj3zXa0vSznnz/X5MWYjOAjtKAaFgAvf2mgLAgZ7eWN
pQA3ezE8ynKgJeAkfcv1xixoe4cHtZ7IUqUTCr1xabd1nijSktmszJx4tHcp6oyPoza1ayU5FBTT
7adlGRWe6YcGDn2TXDh0I58UuX2wOAK0EsO5hKPuuZJYobzI7L8vSCGJs1xnfWtYlcc4LaH2R0f4
E5G6VFfQJbHAm0VxdyNInwQWifi+JoYaeHCq1UtbUoLx5/4T+ZYqxDrawkFW49Tyx/pJoLaOob7K
/aLjhDsqUtmgwY9UhBwMfn65odeM7g0pZWliLihhcVxSp03uveCFNGJ3CUxHoPKVNd64/woMC/Li
EmpgzTtpUEg1dTfL3eaw8ehxHmo37G2rbxIAvau+mdOMUyPZx1akzTfP21Yx29HO56f+DtMR1+wn
ujLrzKcmZadWhSc95nQu5HeYieJdqzJ2CIG1dCsomDnlFYNnr0WnPo7E5JwsGWjW4jNPRHDlulgX
NcJqGB+eGzRPAPtMHGFzg0u99SASHADGwsni4pfWivHMOVJb4fLkLq6qKUzMnlePCyobZan4L6LF
EEvdrwRtGpGwY+i7xUvmlmNcsyJpWghLTWzDRuJFNUNvF4deaIsOyqKOzYDW8N/qNIawsxRjhGU4
6M7y6spw3eoCpG6P7/RP+EmD+rKNYT0EF7RwnlSbs3Hiv23Tuy59gqDhXhbh22hkR6gHRUTB9iq+
i0MAj+dT3ojSvkrXMK68R96guyouIbFMGDw3HtQuhMH60aOnsH3udCBLA9TKTqsRpAc1VCHN2VI7
cSPfFarTO6lkiRlTkU0+ixrp2kwWg4FDcbA+fsDU1H1tT8ly/gBhWL85lC3MG7keWR8+gLJGdXMA
pl7pP65sLW8LX8F6X4vQbVh77xI/rWCkjKXcrlkTSyHbJDPBRQdMyhBnIF6+xpLlT8M/54BkB86W
ehKczJSs71/RGXplQvbKBrcsuXojfpAMZZy8iYCpvSU9R+4OPWJuZ5HEM4HNWqcITjKvmUBBQHLJ
q03hFI2nqJtzPbWvYA7+TKahNWKGhkc6cBvXMHYE9ytccGhc92xqP3s4FwXzH4JL4Z42z1NuscZk
JTrysJsRCSWAHXEGvMIsNcDEa9lwsaN7cJoEUO98kbgIp287goiGRpYukm9VzXTDPlxpslmUKYRH
j2/BffskmuxscAcHoPxv9WUQbElo3LVg+fWe+s1ItUZUe96hNOC56wlcjkQaapmY4G2a75HJOxSM
g9eSV2gDQbYs31NflZgQgkqz4w1Eqf4bW9CqzDN+UZQ28QtT2dxffPNLqkro76PQoLro9baygPqy
RXObZJqjGg7g5RRKq69whcT3GK8euSq7qiV4It5dboSBYNg1T0kslzBCpgTu7Xn8fb7HpfFWM+u3
hoGUs11DYiri27V4ayFPBr3clL7Rld0g+hvaKYnX27MzABVr0I6YYzkghSyO+bzpFMMGgQP4Ir0Z
fXAbGgNYpKVQItAqmZW3PqzuHlFF+2IuY/MT4uOs/nNW+1HfzOpJmp2FI1bTTtot2bq9C1fJRFJm
j/X6c2eT4uzuVEMGykAQUoGvWK6WvlDc2pxMw+lVsGHXrprMjevxm4PUTLbN63JpOeQVpQaggyzM
Owg/4QHvhGyp5fS6Y6B/98V9A6vZ+xK8HY3H2uQWWHny37QMtTkRgHImCiSRg/Ke/ub+k0KhJ3qt
Zxnl3K1Vs9zBYzLrYbHBVQWK4zxn34et9h1Md6lVP+R3xOzzGS+eMErg7guRQz6S9rwGLLdHEn6K
c94bwO+rYpSO4446KMN2DiRisHXn29uzrZDAlft4T8wRo1OuLtT1Z8NLnUkKQDJotNikBAB+q8a/
Jc5JA8Ov+3IopSjQWcEqW/EQXuT7FYTM1SR2ZvLhZsb4qmnY4RVS6c/2ApAHdHh4MNWWSSHmKfRo
LFN5x3Al9b/3vNBzfpZZgu4jLbRKx8no/imtcwY/+464PVHFQvjB21tpxMcZe1wYb/phod05/CRB
k7xcl6H0H57ElC7xdwpwcsmG3rH8VEcW19dWw4lC5b6qEfYLAe0Mwbxlm93u1YPKMNPWZ5gf/vuI
YVBEg6k7unoHnxT9eTX3dcaVWLqdr4BHbeuA8kdasFXokwZlgItsdQ65mhIyYypzIZdWMMoTbUsI
17W6uCHbjLNgB6Rm64lhKUGjpR8CrGe35HaPtGHfwmTJWSG5C5UH+sf02SbScYY0ItVb96MQ9E8e
iz1jViLv9UQ10TNzcDMSH2rIzQa7Jte9Ie5yB8/sUnChZUYZb2rFfNExq7xuQ7WdVr8jSb2FjQCi
jJL9iTLyfiwlCAK7pEDCp+ZzbKAvJ0CiPq8rAkopaL39xD7fdx4tQSApuYcl3apVOMNzHZ71L/vU
b2N8q7L+/0KtDOsHTbh5ChPevYH78ia1ttNn1B/3UJRpXGCdSjH6Kgo7N1JfToPaJhsgCHHaLuGR
HzjFEh23GpnmwdmJ2fVBDoR6f1t9v2rl9OX6e3p6PrJV9WXTiJzW1s/YbXa2p0Wb34QbuTg28JK2
CCGO0Cp9e9QngLGpGAuHUcnMpwR3GnNGVupGgzFq53BPdAhx2Z5QatU3+5KsXigTRPPRt/fY4gYr
/wg0BCx2xvGT1vUvMC6++k/A1OMjI6iQkG12U1LFB/88kluD0KjyYu5zAj8GkeuUPa7yOXXWl39i
V0EudxWJ4d27WKwDtmc4Zff2PrKv7+ptyzqGuQMSFCre4ynhPv/4BKyNYK/BWZucbFL5U4eMf4UO
jfgWbLfXgLtV7dI0HZ2w3m56APEjCFotxcBEX/T8huFT/s/Q5hezb9Mry8POySrvLzokD3AwV5pJ
Ug3oL5uUual6k57uVnCTWeb7Fpcattc1A8Qv2ybMFPFhWdiVKGzEiYWigXG3hcRDLg/zIEw0ctMC
NK726+UZyj8f4bNhipKtId63Bm03z6yCrdnnAcj3OoruUl51LTR8+ErLV/nA219232BlVyFYYRaT
wv58Wsdq3VQb+75Sa2wYYFcsbmu4e9cFUH8NRkJazoV1AYuH9h09tLmkIGd+zwy5ditzXAaDbPRo
Cwd7OnnG5TXI/IgEMkEJCLPsNHGHEVQvI/OzBgfBn6R0YTOw1Nla8amNnKD2c4wXdrn/1D7lPi76
HBAw2fEPBz4x5t9BXMzZkJyNG0O6jAURfqIjIaTMPi6oTDXEVploUmVPWwS4/jLNNgZxcheyULFZ
lkcBZ8efo8ZpSIE+uWjtNSCQkalFX1pSExG1az7C19/FtcR2RtcHiw4Mh/Be/tVqyxjteteBVKC6
5y4C2XQHZF1iP7c8PquIcMHs45oHihIOH9iXw4lQgEvoq1zAXqoD1SxEOofGsCvNc7X5EHMHa58N
HBYW7ywO/MW4sisgT1pUSGNV493EpPNEbHKn3T8PEqNbdF5zE0PC1LRaZKToTVnfbVRRB3kFKO17
xDXIWKgphSLoQZqurhOl4N4aVQ4Y5CStz0bV8ZYgXMDqmtvw6SQ8aVX2IslH93Ey0dgA6Jm5/fNj
Xgr841X6LFAvDApRnih2GtV3EDq/aVCmq5Z0y4EhVd907ZzxdOf0HKjXKJ6IKRBJ8WOcX5bN/QXu
rblP1vmALeehoq287PH1zUUpI5xlU0eEaZzPOgbHvIItSwK5vgzCqp3ztsZDhCXAVTeeY0dHA3Zy
oZttJUSXi+dVZ7YV4qX56guassM0PnV33jdN8bcQgX3xhDw18FBssyifewyY8QLJcgbtdj/v471s
BHOZZBY64GYTIdUz3BAeZCrZU4bRlv4YmGq2PFinXG+uT1EvAF/DKWKTcL1XtwdnfRv6b/qALSoC
cqTxpUGn1OPlksOdFYaLy7ZcQhbcuDkZ+r7TIqOLS0smexvV1cy9hoZmnD8VbRPbYA2D8DNqL9l0
QfdVj40eYstpBvivBAbLdJ1GoyeMzgIN9Yxgzi+3JPLEBt37gTfE6WMgFy6y/dJDN2xHIxGvXsBM
K6+OQYMN5qVeoQt5j7J3S7/dMANrmymxHX8pstod5/3jFEtegh8t0UNFi9iudbLGcGFYyOTXhpCr
PY4Tk7KYzmNjqzpLM26p5GOP+3ipP0Ls8IB1fUPQpjb5HnoRJHZuO+70sJGVNSca2ZN0axkC0T4O
osY03FjvDYSFmvAOxSsubqLKwfqs0tuT5kywviUZqgRMbV75CvVkL4ky2F8/hXY/bTIoryLR5ydZ
SJF+U5trhSMQmb0ukbRweuaIi8WQqSWAEUis1365GF9ffDGYf8mozCFD13o/mG/fFWiawm/mRyYc
S7lB8jabbRUq2MYWpLP8Q4IgTx4na/s9L2Aj0FQSv0KD0CttgyEqGGLVDdzZ8vzM8RRqisEPlpQ4
4+ml+o7aVA4GrgZ0EldbTcNWiGj+YoYNBZnvyIJjpdzk3PI7Q25ALP8vIqpjWHRc1ZlehOabH17n
w4v9IO8CbBAkW8zuJdOaoX40YP9sTZIE/kPHzMfOmit3XSmpJHApnWrJ/NVecgjin4bVVrgPO10T
d+Xh0Kaaxc7NVOmRkP53pxQHbzgYNDoY86KmGAhD1f6H3x53niQWxRCQE6xEwXHBdGWSNL+zAg0i
40145Ygox31Lb+8kVP/g/XNZ1E5+K1NIuLbg+XcV+fYpe4km+kVAJk/vE14zMRyFniQjxfV5c7qB
mDID9aOSCllJNamXg/qLlnCm22RE7bu7ENgtV4faCRNE2RRw0JXKWR2L5i4eXBSVIJyCiR6eqo/G
DrG8h3Z8Cym69iNiR+mRKn4xp2AYgqhp0+5rqMykH7sL9gor8WkOlZy3Nn8PkOyUEWx835LEgJGa
gvxwvGelnFxjeYYAG7vclEzMoLmzIVrcgbTBrIvMmqwV6QWqmlfiX/s5OIXO9xYBoZF28vo1hdsT
U+T5M5CfL4PnqEryKSw8u0lOWstu5OlVBrRr6wQdDP3Sz+YFi1MrkBU56sVILytBw+TCbR3GvWBJ
ibkIFI9x1hTds/j63gi+5/5lXzgykyppay1ooMo2TflRRZ6vu1DAie0a/dTOPvyAoX4H4Cv+oC9P
ovTMLheYVMzRwz5vyHq2NmUJmDr2OMZcmiLE2DBaJTLDvxaDqCeu/X4QW0TVL7EEEMsETyo2f+L2
5cYY+iLBlbGrU1snjcL4fRnnslWy2kEVweFReLXeDbQDqs2GG5u40MdE9Zp9/seCMVue/NAK0vSW
mEGT7Pwlcku9xYjseYcBWlq/3CHTjKoh4oWW1nXTF4yacZnK15sQoK+DwZaIJqvFS+F+epkE/aaW
t+bQsh768SoppZEHypoSbF5/nZL8lcMQHCitxuFjTFeJqJQNq7d4drI2QuWBUNx6d/7YleUUyxnP
a70slt0Syn3rVQEa7iwMe8rSft9EdnBS68wFqO3/WqurZpBwodBPWhEpS6XV0M0C2p0+AI0T9Urx
oj8P4+ui0XaVlVUSQYm5XW/sfrYuz2tJ5U0SvKBp+j/GfmiJoIm+WcgcMbT37Uj7P+cPTmLkZil+
42ig6Nb2Rnlc57eO0gmAd1SirTKIzUdBzko5kcGPbGMNs8WLjlaQgFcy+mLgBXu9+GzrAlmO861G
H8vzT+A8/YIHIVtE1/IDlXemPHgxB52cXq5vvFjf7RxEA/GvOzYYzRYUIu9zwWTTyI0xOeMvu2LC
dMA7MLfNH4yZgbGhL3139yB22usD3JuS9T3VmZYSavFvbq0i1sZfmrOnwoGmqgm0NXwu3Squu2mK
yFA8pxxQVaWU2p+FNu/Cggzx24FDrL8R97iiVAVFBw0pFMbN+atWCZ3QvQR+8+ZNz+dNSXvnGqx5
zpGM3Y3tLM9Veg6V9wWjbYhInxjr9RZIvKEck8yqs4LyObgCZenozFNZGz2S6J4XmyT9Hv8Xx8IC
pFKUWlYCFgOTm1wlftCbWZso0Vn1GIoDhsMlEnvBj41x1MrM44pNwCliRIZ4fkiO6ksX24zO6cSE
5aDbOAttbF4aOrKwoG4GuOci/2FiSWOFpHbMWdh9n1gZXtjZOY8LWWQjiDQmPx5MKC2GZoSIIpip
L2t0iWk3hVff2AIvhURdwer/86de19Eo7uusLLQ56pLcxE7FnJAGNaJ151Rzb4EFF2gGLt1vfgZw
+cEBcglxOEicen3J/v09w8a7CtvCGOcwgBivWVtTgRDSBuUBB3Kdim9tzG+u3Q+9XohVwBQx7kwF
uCYTdvHsak4ksq1bXp1RsU9MPFlK9WorTx/xHhOZo4TK4tc3HkZP4oLKE/jve0//e27lZIZ8kiCl
NNyuM3A/T1s1e6NgJUUIGfNPAtrdLiuevrE+VxaUq9ObfLwIlolm1fy6fpl2R/g91ld/d6C9a1zr
d9WwkKwaRoVYyXqB0k/3qZSClct9665dckjMA07tFHPLGZ3pT0TLlSoGpiILVFXlNaj4DtRIy4nP
vDGgVeVLeG4NM8iiMNIiuglE4XZla8sCGagOrL/+OghADw0lgrEc82pXUB0z9BVvucFMZ5Z10KaS
9fwas3tXZmUUQEz9FuVDzwJAAv6nolRfvGDlZ4NZtZtPxW6uXGdTMvXNdb9j3/SoVLCMXZ+4G71k
7o+awfZ+GnI4H2CVz8MRQdj63H3iXRc93IICGpNYerIhIg8XWYBH4fHsyoRMLsNN8eZV8etKIpaH
TTvp2rUXr2i0hNJMsT8P9exXAM7mM4Wu8WsiAQsQkl/npRwW7a30QRzeBgWr5cZ3bMIItmCPV/PR
v0VsyWv2DUYEtzotozAmjBxT6hFdAPYfM5HeMp+fewRr6diWGW7G48dGWKR59ieYbapoHeF7O+WP
TbK8Jbqvk5kXn4v0ENb2Og5PiuHv8f0HM2sW6k8Tn0wzWc5z24s21hkIWlnpAY8ZcjqBsMe8n+ye
y9EcQOvtY6DBHawuuW+awQdI9CmYvd8vyTKMpxRUFGHL1IGq+H8aaXYizkc8npMwbLzwhCVT5k3C
2SjzDAboD28lWamU8ANUgbqnLLE+JSEWeUszL83rYq6J2rQ7x464UpJGZ6poHRwApv0ZjjAaO+k9
AfjjPdWiMDf4EJg6iv1+xSrZwg6ROMXibXeMNFg6YkZt3OkMLBo1GPew17XKFWASkZhjDZEs6aFj
Rq8Mpxuzol0RnBFTMMrz1+FDzvkIa0tY8XsC1LsLHyf8RkWLV+pTv/9Bl3qT1ifqYsoYQxZoBOm6
mWYJo1hkYxURHM7ofGbvDRASOWHReTKJDzZH8ET2A4KrguflucLOL11U7umJARreA9ET2dZKlmoL
5bdEUzG7CI2Is5fnnnZev/ZQnijCm2eSt9fPIzNf9JGTSkloQQyEDm6vtOTtMzyNGFcy2Uzmr8zx
tsF4ndo8pWlajm4EUjARntwkFeACbV2CqXSb7XRRUpjwoG9Xwm9aPO6eoibYApcfx2I0NK23elal
46FhfTScruCuYiRs4trUF9DP5fg5lz/vT2G1hRYz0+oR+4JpDYwf7mHhJs9nEjNJvAjyBB8zEIuG
ZeMxqg0uQVwHDQb06Uw5KfvJugqAIgbDuPry7Q8L7hRZh73jHV7G60fxVux2tK2eUEigQCT2fY/J
FBdJ+cT8iZHTDMklnQrbBXo48+U5rHk+ccu2Y2qYJGLwwREctWXbu4Cx5/ATy49AtYGdp8Q59T5J
LhSclzsDdFkGqva8pGnUPkxA72qnNlBIneTmEjwNBDApw0dYwWJQwo9s45m3YYKN0HbLaihpgCvD
CquKHd/KkQsv+RQdH8Ya2kwHXzkb7YUnzC9NDGfP/C/3+USkea2j4atxVdYtB3MZP6EtyULI0YSq
v8ME1y6Zj8RQeM47woutQvpJulnKLyLW7slMzZUzaI2rxG0jrklKjUPZVIPnJK1Ofkc3B/MCToxd
7kqdIIJ8NAqbvnMgG+42mcuiwwJzzx3/PcfGOIj/85CqGomNhnC/3Z0nbFCo3VoRk2SAC/xAXKmB
4t2SLFEs2dlV8HAMEUCZWMg6sUL8tMXtU054IYHUQfpwpQIFfh+IjL8uCohd0RzfzdvHWvophj5U
ahYH86qpGDkKJAtQk4Jh+CE3qBqlIdJxt4uPwSF0Mov/erMPikHuBDUqG2dfcgo0Dq8/vopGbXYQ
1qWpFH7FoiSpbtI95FrxEzmfCvv5EbEj7/idw3SpxNoX7RKEOqu/LFchIdE3LZ+ihg0JiSFrppxo
Ga9RNWYXXO8t1LSQYZa9CisUFeZTutj4QxTSs8Y8FntrfcXarYt0OFo4iBdh71jw/AKC2TDn/uka
Oe3lisHzpvmVqGFkSVZh3ZQ6xJNjNT9QfO0ZHSgN6cl2f37JnV7B80pb1HHKFx4zuGXWDK0EAidF
zn0a1BqFNf0RX3TSOS27tFscRTYNgi4RdBL1caOVUogFgpqaBV8hYCzJOnTmoCezlzzSIrVuhiP3
yrkEjGquLBqVUFCpNTveYMcSIkvNIyn3dUzzu3lWTuGoGCmDKv5qjUe7vAnkk0QpLPvAYnDV/Ave
QymdWpscuLV+pcGLdVduFOWtP0lagCsePIcAp29rXBG+UXncWIxyJYHh/YQo5r24TVvHUgGSThBA
yNuaDp50UjPyC1t7hCKQ9VpU7/HOhmeVWycdPPDdNrwB8b+nP6jLn1frU9Unin2+Ww38LSu9rJCH
xlfUMD+fHTOC/+KNL5QRbhKII6Om42RvF2g3H+FklGZh4r7qWsDROPxQK7/Fwo7sZamXjAKnYUNh
SG6KzXT2YRS5MgCLt1vhAeZrH++N33XyUwRIEfOWOdVbafnfaBIMh5Da4MxBevWQyV3OkvvMq/33
qfgjHMjkFFgkD/dnpqC7wbEu6QwaIcaFG+6hmBY5JvEk/ikuyjqwUZKSFxe5PyGgQjjh08zJJ7NW
dnJ3wAUsdsdOmhD2w136AAPnhMkt+SbFfLWmnhzvNpRjP/mjEAp6RO4Cm/eKrTVnKN17Y96oXZR8
euRn4wZdQlWZ7ownKa59bHlwb8Hgwr7km6vCIw/v2EmaJ6eq0SeDZKXMnHZ1/S76mO5jVQxHysGd
dSpG4BQa4SESOPhJkFwH1yLYyCoJay/GNigjVJqQT7F0NbHbQyr0MAqtreUvqZ62XX1tDDP2FYEx
ulbusfdcH5oIgFoiJqhDPTlFAtORYHEuxfyEgYQmW5b8nsRYyUNG85SqN38ZnSoRZ7IDKlw0rWns
aYWUhweXT2w7QVDTupASadQo7pNw0G0KA3biR1ggDNWDK1qkuTarfTI+wsGwqVNC9W67I1pLuD2k
Fja4FLH8fwHPbOHiF8mV+87JEAItYbgjUf1OYQows8alJGZwE8eLPEQHddO74xS+tvjCi88exP90
txoYWCora39CY0+QnXHUWTSdLEc1K7cf4gm8vfhuSBEg99JmVfiX+MY2m8mcl7gFWnD52jOnwiPu
wNR6KskX0E1gYrDZ9EaV1tY8XJrcRqlApu15fZF6hWfB1tT0OZ+3MvEgLyCENnJxzdadZVz4g8jC
7uTwJC+Cj4Ng5EoGM2RLa5JgjlEDw+Nern0Xu+267FiDyIpxZbowMOcLeygMD3Ka0AD038NgRgCe
po3L/Cicp5L//ZQA4ho8230CWZprQpbQbhRgf8/cJp3fj6aY56hJ7CLDUOByvW6R/D8ukWcfMusr
joVZzphMgrCRzX2zKHcZkwVZVQ4BESWIuIkagTM7ob8nKOnwhBMSWtOscBVwhiHiR0USY6huCHsK
EFmTPixKWPAOK0/kZuaqRBdN6QE/eIGzlLo2Or/lyQwn/2fCN7SdOtf8ZUwZxA/GgGZZtGKntzBT
XGzBM5GsQ927x0rE6glWxf/uULjyADbTJ2fkYdeGuRM81mVIZQHqHf2aY/z6Ye4xyf5phg2Q7hi0
9wPF+vF1Y3vtHNYnF/AsFTZ33GWJUhybF2WqOJihTkNuABMISl80XkcEvbqZovV+rjNivlxCAbqJ
BP8swHgbCbGlb8kPVrFW7lh4GHVNEJWWeOtRz8/t73DnaNx6jLaWjr74x88tT2zFMDZItW2GgvG8
NwMmyvK/34+btTYdFvf+vqc5HdWbb5W5PXJbz5u0Q7G7fLSWAtxeZRNIREqJA/cXKQoWjL0ZZ3M7
Mqt6fdyiZwdVx8EaW6wjuGtmvI4E7jflqCeFcUm83KwCC1sQG4F6EG8I4gE81DfuiGDTcXIFt9l6
DrkBY3ZlsoFzJ0rAlwfjWL+ySGYUy45TKF7V1caBYb0yWlqXl7jQUr7tMRp5CgheW4Z6NH7SbFv1
M9H0g5eZalA4tLtmJi4PJ0rqPKer1DbixfWAWbFzATZKcruJeH2Dk9n3Mf7roWaEjOkWQ29Mr5YE
wrK/gTNkknt9m/OmLftNvkyKj55eRLjkDPUpgGt0trGX5JEv4gm4+CHzpfo03IRMRvvbmgk2bDqK
vksf/Z6sEcyu2/Vc+AasvoxbNnYJdLPKTxpQV77fxTjampqi5uEqlkxX5tWscd0SbRIBA8F4AQDm
5cJTtEWdzgaOCFq25mQ9rvj9nyTH/yBcoPTtilCKzXSaZkFryscxDwso1f+R7ac+V0Udks7fQzm0
OOHB1ZtQSd89sCXoRf8mlLkiDdJj88vkaLFA19+BAVRaXWHzcqNUN8ZQxD7TSHODmrMMKojbThal
Jpf4zcZcu2CeoZo/e2EJMXhVcQK4iSzlabw0Zq+nIKr5pEU0XQHdAVwnfRWhxD34vMOg298kAk71
qxzxjlg+7ERomt/Aa8zSlY25flBWSE7fxmGYOBuLZIzY2Htd1nDcDrunUqfP4FZi/bDZe72S4EkP
RhiH06qahkhzpxfi39Irw0hsbvRuACC0artd4MyO8lu3ta0hANYDJdVDncKMNG7G5RdVKqhaXvfz
g6KGk16T9RTpaKui0ri2Ik5L1cpCOGQncC4EIYgJYeYE1dxZf4NI9/lBqnepaMh27dCHLJ1QyRaA
lqqtzFqGxy2WQKHx6rBwyWRyV7G9iXQwk61H1zC7BaGeZp6AN6800ppd+cxk9qHtHQ0mj1yrG8Jw
lfRtq+nRVNjLZaFcKslARCRYvumqeI+FwPupNeLgX0fQPqnNIzrMnvH4xR63yI6VTgokTqDec+Uc
NtwAAg86pUDgD34u0bpVNdVslluwAijaa2+wGasHE1v9JsctZeKjdnArqLz6bcIj7IjPZ8cJ1KCC
E9OTlU9zhy0em7Ho8iFQ89aBDCq6Qvz3itzGWNhdtuZPrUZdalySZVhalULqUB32MxaUc4M95g0t
+NGKKyuW94JhTUM8YTlXp8woigatYHJNonU3xw6Sk7IqWm2hQ2l1AXAW+mqMGJn1NAjcsjA9X3L6
tGM9nlicX9CsSRsN1O5i1rZvXadPXOmAsAIxzZJzNDrdUbsgJeTAh+BlUM9lj1Pn+X6zOajHDdBO
khYJw/pEAyHEkqMaQLygyjDDa3HY1quEkp3bSd7rFwCpgyPCTCtb9G1GUN6CQp3HO7QbCf/ztPB5
FnAlOl+U2wu8mAgU50MhjwRhKwu0BH93MGNiu9sf7f31e7yvjdtNKj7SYZXPUGkOQc4k8hPVnlcf
j5m9Q/A7JxcrZAWI00X4qNNqY8bHtsBhE/EFsE4yUPqtKaVfs9mXuI9+B2UMVfbRE++9DGXh3Rm0
aB30h/DEEMkz6esTXU64idXdlSsKdxs9prsckaR3ns0Y8dHy33+t5BbFgAO40vyb4AEFgDCAmbTi
pobaJbPoruvgKvHC/eCVZiAPE5P8bVikHNcmNTQpzdUpQpd2NA8FBalBKHDG3MDf7lAkACwQS9Ts
fGlYNlkTN8OBlCcGU3NdMuexR9CDlwN/GsZQ8UNSNPj+kUXlIQKQGkMzC4jp/4DEsQVPBlMX9yHA
5w2vIcWBvBnuCASkq81Tv8onNDshwqu2966ZSrd1x6hOweBX0kSi0Zz+c26BsY13m6NfqK5yj/yc
gS+xa21drx3DS80tzAFu0xdn/GqYfhMCRhZI2l3TCje7IkCY8bflDJWOt+vXigs8uHDVhh6RdB52
TkfFBFER2TKZkN67ZpxIJy1TLSp6dBmUWnaR/1DpqChtlN66Xm5JOnavzyUjO2HIT9/ZVZl9uEQC
cqkjuIOrsnQ/goTxdZ8pPRoqHHHWxZ2mf5YBiuR35ejjQzu52+eSNKM2vzLab8rxrtg5mvnUox3J
DDVGvbWMmV2TLN2wqdx3f/fyJ4SokOVi6Cr2jMLdGap6D4eVJn0MP9P9K3Rk0R3TrmkFsw9uiF7/
oHsSkP/lC+RyGCCBqnlFx4sE6ayoVvYPOUhAm8vB9xQ+ciGxEjXFqR+3ElmiBbJUZKUd1z1XWxEb
ARvC5IV99BPoJNCAi1qzFksF2I6wvl1CToxq45B/UBU/sJQ45nAOEgG1xm7yiUB9yTcb1eLdTAwx
aiKgy4Qdl4YwuctYtccgOqrQZzOx8kYVHiJN7M97kEv55E/3uQQdnO9DvnvEebUfpOiPBi9pXINQ
XZT4funDiSRj6IuR7aPFtr8BonQ9rkeNXcnXdbCN49UNOxG2PnG50FwluKmLnfLzcr47Lzs/QxnU
ivx59BesujhYY1Y0fPKdGtSywbQBaH6G7iYvpq4BwVJ531QrW4oSNmNjvrJGsI7HBR7GJbe+4SWm
wL7vexSGk/vNiZraHJRF16e4fWUzCOMVWEQpnBqbguTmp5SMEU/S3XcC5uMeUh5C1KwmRYPycYxD
J+lf1YuMcwYTAOWO94NwlLrM+ot4tn/De9iOyGHAe0fUKK96kVDHvu8sf4ygOmo7XydMvKZ1p1w/
ANQREJb7M3btu8lA+BSWa98/H+S0PEJIRKPye203yiGRXlm+0HYZ0rFa41MbxUNGGWxlvpthpCIB
0urZot5rTBP5C98e2xEEhYuu6ixXSqBArLMKI6KSv/Xjig3WrXL9mDlJhRyfmyNmASvyQD8abavu
EVeVChXdY7OOs27A1OMWXJJlLO+2qIKu0eNUIR/s2x/4MlZdD0GbKuiFm0+UgdYXsICVni8mg35t
Kh+sAWpbZq6+6ysCWvz9+1JH7iSLbfKUJQVsuYYDU4tEGuM6dwnjZg98WWTWF1wI9UaQP1Fd4hBP
YNSA1RxmVmrzjhPPVGkkW3m9aZh321gHcdBa/S830L1c6Q8HU47BdM9pZ+PvgNGXd8l9muYeEPxi
KFdjuVeQH+w70hp6n4atjPfGgPqLdej0i/p3ufyOzsmkXFi5nLcMdUmXQDE08V/1Z836pEm19KAK
H4cZpwgVN2pnzHT+NELiV4VTF94FeGSj8LwYIhrR2XXSLQrRAPEKi3B/s0654WsCLoo7wxQPgz9l
8dolN4Fdn5ZuDIooj9jHlo0CPY3CgSG8YbbYD16Y4QFursfmPTfueJcG5NmkXCr3xvbnY4hBn5nM
zjlZXUBojClEAk1Q0pqzs/IQMz3pSkWkYvaPM8R0y3/cpUsLD2LknU+lJavRPTHvTnrCXRKSTNMG
3nOI2LUZ+5N2/HgMLihkFKtDEQtF4U9sLdnacn7AJ4cTtgMMGgS34Mx4/5H8bABKmRbZG696ol3z
bHUq5BRiwcWhkffQUfJ47tLxcBgbePIma03bLw4sfYniRef+4SKdcNFJMiKXrdEPLQZP3aOUKE9s
5xIGbiFY/QUBl22iqXCsFL3wUTx/zid0lRp7ar4jM+Yz5ixJ1ZSO2nCGrVyv0l+9p6t/SYyFCTbe
Q6BNiJ9AdUY7TYYeULgf5ZYP/v/4lSRhUTPHJF3r7PGaho29Ntc7lieQBNj/laHLjuHRlr6J/yvc
WgusVgrn8o0e4vg/+Ewb+DFnmlNH8J3blozn66wi7v3p4V0y7fymjYDS09qlZ4zKZ8AgAXBM/2DT
vkRaCTiIyDu44eYqlm05OVfxA/ZUDpStbw4v/mAzuYdv1cFwhiPnXyNsLYFgTt2CApTv1JFKr7Yd
gl6JrP2exO1Ap8tEsp2vzo6sGhrgpm5uie9JnBDnnOBmPzWWhfHf4UtqidarC2WgemFtA70yFxxz
VK9gwIMZ1e1r/lJCkBE1aDiB6vn+wjNtxWFpsL7aHiobYMJxcCppSctAAQqeldnFcgCasKUPfF5x
3ITaJVYqffi7vAH0IXfomJu+FMlQEGocDeBMcR8cSbxTRWQQIhbZv+9x1nv/y0bQ2ZFvBcJSkIer
Yu45NDKAl+OK9Jo46lBbn7CLo922aZ5n/RSlU52pqg73VrMOzMFXwRPcMX/wSV1/2G/g76y+TAOV
XOnqOYA1IPFbPVuS9I5LGWLvCDmwjA713hzhyxm/sGJ5ba8mFGJtSxcm40qqVrYU524DBFK6Uj21
bJogBkurA6scHyes9F5PP4+9nArXutq3o44PzQLmG5URTfvWTLinHwwV3/ihck61hKsmrxKvtin3
0Dz/b3Sc6hM33q5vfa9vite9fwU7otxl+W7mVd0l/L2VfI2k7tlMWlXvwmErHxo7uWoM+Y5wwsXz
hP7zW4vJHw3zJaxsJZ0NC46RdoIHrjDgnD3VsxJo9Quvx9OCcliBiBNAoxX+wZOtwbDBya1T95wv
YNsG1ua5YLShwqKxnuv09zkHB4LlpbKBVAf1HzalMItlEn+0aa1+AO9Nf8liO9uDhZCO3uJeoQu5
67rxacwRzUC+lo+O8H9RW2wt1G5uJPlss8zF5oVqeTeUMTYWg4IIDJsCWIWVBphWt42n97VE0Aup
lTt34qtqy4NVbBtWi5NR4fdF2JOVQEm4ixHHHMwds693uCcT/iyYE1UsVcVAe4v1n/lN/FX0JWmQ
CIbAoxe4+PrEAD0MGSQCbSRhj79lEYco5RFsB7gw7nNyvtsQt4aDF5CcxhJvhzPLdoKcnmMdiUSK
BrRI69OkYE+xxAlsjpCHIw+rsETfFq3Wx9iosLEGtsKA9r+5AHVdpC6VcnJKDk+CXH0bjIhnTYjX
SuBayMZTgV5tEYU/LFWb83IKILSGqDT0pwKsNVdjIBAQtYtQCo4sf6xm2MaTznD0x7E1ZHziWYZs
cUnCz3J6L/RWYwT3Nmx5zYu/VhmYcZA+7kMqqN9LkSPBaV/6GW1Rz9KAjV85SqlxPIdlXdWK8yga
wtW04tUuj7zi09hgkCxTy/rKzfFS47tHKxAgNrku9RuIopYrTqlF2T8gF45wRG+ntDi/AMzg8dX3
Q0mL1zY1yix1HiKngqJ3X1zuoBxZUuNgdNWl7WkGILIWDZb9iX1XDZQs/dSwjpx1JyuLb/ajgW+/
vLSBkW9MuT7l4ll96O34XxlQpVjTX3wLFThtQx3BgPZkLjBaIKaCwl5cku4x+p3gnqY7c/II57Ql
eBaWT+kp40hofK7VxIg8m/uvuywpm5nSb4ZpsxAf+81Q6YVexQ6HpxEhHZc12K72oAerOUVyO7ko
ckncX2z+yX5GqKgKPKHpCazRdUSQQ/AHtUeyqWPoBh+W5Dpta21JDIUh0t9MyAs9L+SwHGw5L9fD
Dp0GAjor4l0ZhSNxvlMv3Ee8QlD8O74dwaLw0v6SFbXgX0KTzQlR4kGJz4I2k2pbsDlj5IzJwsgm
vAroqh+Pvbc9k4P3jr9/yGqtQI9opjoDebRl23uuq4uDUbNe/EHy6EqH/DGg/l1sh3EBDbMBQRZf
n8d2Ru5EDW+k8ofELxDzfkTZbWhqo5djCV0vaJpHSdlnekohwrHplFndMYjtVXdztMwTq0y4G3Rj
feCck3OxhLy//fok9F9cs6rM+CX7hd7h3aVvY/2Co9ow0Dh0qsYsEULNc/xNPTSjuy4OBcv3BUHi
wkumi/YTKZHIZYdOJ1eE7NcdSlo57A+3uWh09OLSV9FQw1Pi8b5OUPMTwHM+OX/LQWibHHLcQhJ5
84JZKvUZJ68yXsqUfOKMtZjOp5Hp515ugNJc13MgBrf+Avzj7xoHTEtmTC9uTx/G8ZwwCQS5jNfa
9WLd+yhIAfGnSPSfq1eeXVW0sODjxJG71TXWtxMKEXBPrpN+j1ssh2s39fJyRzke/nJpyOGkVBDD
cDpRX0Gco3tdley1bfjGVHrGymS+ifUBF68GHyAGPqIHEyzBxQzgokZKX1ZVRh4FgBScUjDrYc9J
guU7r8sEuakMVW+Ssd1C1iXf+gCrUbfJwCuTmVtsqsuSdula7nD3mOv3/lyYI+J/yb1p1A3bRt10
UiiUOhXhdPMdY01h+00gPn0b7rpA83vMmK0Qfs2a2vgOSDccgdJ5qeWGpTkYJmoQyFcSstXWxt3m
grvUtkCMzhyj+dZhVBmAT4PgM3iQ1d4QG2egqddSXHBhXK96EiaJvYYT9kJ+tEx5O9rMqJrR8UJE
j+BTlU9X+0NmMOPNbz7CnB9raOzxOhb++vyR7yuZcUPjtKxblo5jzqBIQWWLLIkuDra9C/ZW35QK
vynHaNIuikmAacVfvq9iieFR2e3Gh5EKBc+im42gDpW21xQJfl57Dha2HUxeuoZyyrPBUPjEjKdD
A4ayUHR+qv0Bz9aa1z508KqH0DR4rOI+tDtqJCVlm+gIi7B7Pt8UhqQdGNF8NNDe6kpeCqlpIIpE
57bb8kL5XC+ADrIt8wREBOEj+8JcEpuinO+secE4oeA0hEmXLSPCf1zrVYozYk2TninMQM5YtZVe
5rBboLmtfUpT0/nb7xyVTkoro7BuxQjoKXklrY6G/tjpw5aNn0pKKCbJKylJlsahnmKjN68RFW/3
bgg7PGEU9z9X6aJZatEhb/aQE9ORNWie2iaP7LbYEll2RGxiJZ2vcBuex+D3rkuwu8sblnDcozcl
LXq0iuXvCpDLOAP95Lug9GIiOMBvwCMsDIdFFteQuikLrXnx7YWWKvnL0ZB2upeUJbuXIZtgI27H
b/vEoGUqbZ1RnuE4/zhOZrQu3t4Ime6LGSO8TfG6qqQObdwRoh8YVpiNOB3+fOI8gLWF8nthEciR
qE+6iCwy2eZcUptILznjGSDyg15AZe3o9QLO7z3AB2Xr2U4diZnwCaPRCJ60S63Cu8m0SVN79IfP
CXwTEvgz/4730dagagY/FKcfUs8knK0WmY1+XgtXPGy0OnNaeIBAo1N/WFdpzjTH/DaSGVVSqUAU
hCEnQjQSpNqzMtX1Ec1gz7ETeEbKCf+suy3RD8s3Qle3gPQAFY/iLIYKeqIN9kG2R0P4fweIPoW2
fX6qOePTN+viGA0er7ONlBYSQk9KWPBWydbp3WzYoDwsgJgQLbVnum8LVOz2XrbNLDzkFgXaIFU7
ThZWN1iLOBHTgO+G6Q6FAERTiPyT0+KxtrAHlZQTzJ0MyaAWFxzbkq1vyNGUzLSvjBogInGTJwRH
0V+FCKaM6VSWe1D94pquyNCxVxNECGPHUtLbxvzkuloIZ/C+DlNwA27vj/Cy3ioZaCCVcqeR4w14
zg9GL7w6A0oU9JnNKhGQvx2lwOeCNPq5xgYXyziKODaEcVBFwXwniILDpAg05fOufYZC9c9n0QeI
TgZ2U2amYgGxgrIqbjo7TSx6HSlvK6fUyCpl7R1TUWZDegELRjDPtD59wgiYYNjfPWUyiTYaoXT0
x/JMQe1p5Ne2CnhKGQq3eafzNuTrA3v/ogi98l4TLRVEWTojP+mDGz6onZYGQYx8BycS6Cg9inP0
GpdtLqjWaJrtXrtaBYNypo7jVb/LwDK9PetMCnMVNg22Z+Fa57UT39iKl2fJVFAD7MibDcK8HKU2
r30o1Dq46PgTDPGLeLxqSdhbMv3OppVWzgYdKl96WKzgxb+3j84313zefhGNH2ANwS2Dj/3W8AA9
qOIqq1m8jNlYsoDQz+53GGjZynDboBhpMfGzPVAMIJGyiQnPhuruLhgzRYU8vX0tLgwCwEhyHL6R
tB4Y3DnGoTNhhGek1pmXy3XgIo5VFaH4Awsq9fHTwLTyq8UC63ynw3eQN7sG978zdhbI817bwVI1
eY4bRW41uQ4+1IaKbNrPxVtn216zKG9eq5U6ybRze6WRj7QPIZY+0UpVf8kct+KMVT8kvCFDkurz
qCHpt/u+s1+mpiM1a4MiwZUSMlhgQFcC2LjUhX6XpemYY5XW1qdVZtzj5FaiY7l/98mkzU9dZQ/G
OGrWiBuWbX3YkESYCU7holCb0B5A87vMSls64nEk5IoFfQgnQG5SPjYjSn/isyZI7jcDOA2FODyq
9oqhvPVXrnGiBAqEjZRGdsBYvWa4COVoKibQBmmEh8BdPJvWG77Yz1aEV8xfTPPB37qF9V7H4Ff+
MQBaMUl0wqu+gU3+qCTM9qoRmLaZGeRBo4q6RTf1FuzXIyS32kf8tiYdgnZV2cpvRNOBc49kZmvP
6prM0dFkuHX0PCC692FSYkRdX1FtxHjT1MBGFb+6y9SNtwRfKzsQmW96V1brgsbPa1v/kCGcnZqm
MFuNGxNhsp0bDeMfkIIy4+ZVPokzwftNMYut2m2qatHsISRvMSkNHR/jFNVkIpbMNh7EroDWdMmd
ReP90VItvpmTEHDjHhr6m5IaCrHKqtep94oevCFjvYzFlXrpsH3VNDDK2izl6daWt4hTwiFj1+6j
8A+gbxh9Pzb75kP2Wdraq/3H5M07kS0PH6rXHNRpyq2Jawiq5lxD7l3l0tSUigpGG4d6kg49ymXN
bXtNe2gDFhetaWlRI1bHOiGvnjOafuJk5lFysHRqgQaVIk2UpkAw1xZu5XLzzx2fQ4oxzPN8BvsY
eJKaiprk+6F4gKCP96kEAHrLzDsdx1nH/EwKVH0E82kNIsqNXN6prjKiH3vNTlitOyNAfvccHXxV
WeqxPpQjw4ItwMfHRgvDBlTWQzB6LPDvnskKLm/c3/xztWFfFEdTrxi4Ysdpp5hsESRPVBBi8rBJ
Bx2e1iHetIj3zpg85IuMu0+Ppz7ybHrcGxN0FLuwpNlaF+PLinfywyw40snG3ookYHdj4/dvmb5d
Sv07vpeOLtGYN7bjRm2ugBx7Lr2wrwbcAG0eWqsb3DUkRxX7FUcE+ZvZpYdtVuloKf7Vu3TeDDtI
AXZWfzFxsg01KKxsfJ0S8hx/irLD7BxTA/zVmahxbvk+Cjh8SY1Xh8Aovoj3IHHTUKIa6HOiP4DW
oZPvf1K/dtJip2D3cX6NDPyqJViIIeT8dK9ASrBYC9f0Pq3/cqV+G1lb0mf/zYp1UdzIlfSBJ0Pg
0gx4wcgvKzhfBIPeuzt8C8/djaFeL6c6zXN6Zr9QxLxlbeoF34g7qyiGFN6eXippOzStTOfMbZj8
TYZ/ptmgxSb/44HxEANIaCgJi23ppuHd8o+JSgWVHqhAmD5N7VyxRA9uN0361AgY5aTtjXq66kbd
Hjk5Helxdv5mkTNUdi8P9VqETJf+SJIOV8VFb1Trv3L2J7dqHsmYRzkkEf9gH820SMwjEN9A0axX
o04pbUo1lsWJwVMd+OCq3Xdz5qvObHtZgYqewK2DSD+U7BACbaN7aW4ekcPR9Oj9efqAcQ/3tfwK
taNPoHgF4GPCM70m/9f8IW6GMvLEzN3LonEjDZyGTmz+yGhIJswzmNGzDonHe3Up8N8bYJQFLplK
kGEVyEg9K1aemsfv4twNgWWfVCm2vvJrEe/+tPELDdalzNCUXvWa0WzDOAR4sezBf9ag5SgnEVF0
p16dhgj4V59hF2nxap/r8ji5TI4ihDlxkxCT4EmZwLkrfeptte89OBAsqLkHqf96qZ7UuUUMlc/P
fzmhW7ZLitCa4RHxtX20qWQfmRaN8MCBh4PtoR1QV7vRK3CoK9YfcJQryv8vR67JA61f4tinDeZx
BPpDWo3IBrzbjokUXOGGo+2S3SSvHS2E0/N+2smdKgsSMo2uyKCNV15GQzz2FFTxygkaE0pdoIgB
/ukeXTfSOykoxfI86Po6/k7/7isFf/XR1ZyAWGPZv57lGsAyMgZgq3bg5JVNUxAvp17rutX1Zzrq
f2fjYG9m4NMkbNXgu74vUZGH+nLZAJoU9EH55VL4hw3DFutyjiFrAIEcCZQnFV5Mp7PkDsQVMb6/
r/4skuRZ9Yvq3Biaz0jpqjz0Ijwzq9LntDXosxTJ/Df7zBPzALgzvd0scUMq2rJLUjKvMzEB7FKK
c2ex3thcePQyRd+Ejdiy8uGI6co1EQa3zsgPSiIJRKZsL4nlrHPUe7xktMh517K2Hn4XuICd/ZQD
DfbTE/AuKCK8/nUy7IAfqVm5aEPYSaZNOQ9c39PrncxQo9PbsHYKvsbHffDRzqLVVaublvhcnSNO
8PWvw3XyE5vWG8BxR88j1TRFIV+wIM3RHCh2ACQTmHsvYLstFdN33TMajDRr2Z5BH9w6jR/p2jzP
O+0O63wn8mOxnN846QrRPh/Uj4+HTlaCxjIWr9frYu1uFmLjka1EUZvKSxKgZnD7qqO/oOiOaHIn
yWJIV3ZRCOW9YpgcGBZIWQ43xJUhuWkSv+8zGiufvl0v9ks0XCAPmUOD10PGTl5OUupzDoe/z9ER
bhtNc45OTWhGxDRYG+QbDOLKNTKwWxXqX2GfL0DWdhKOU4qrEvaR5bGKopXtwi7zAlPZXAjyUZy5
F0cTWO6y2cO/WFaIiSJNhOpdDAn/3gDCqus9/klF1BfJIio67UArmnyXbgZOxHEmh/iry+nNiFFt
MZhRsyKgROqaC3WP/9fVB2KjgDLBvog/6wAmsHSN85Xzatdj+G3YJTpHs+SyKLtkSG1EvtNmDtXh
69ZlqXj/mvuXXHjYv9yCDV91cBJ8/MojdDbxd9orqYigV3L34X+P1mv2jdoEdmY1ZVNDqS4C6WSx
/onILJmJuL9olAKnh35sTjA2riQYAXJWI3B69ipoLtaBII9KLhCA9W6Tb+NNZwds3d5vxDTg02Xk
UsOU/KA4BHzvNPNP+8e0Vgh66aanZP6/cwYnnoYloLKN5SzP7jwhoyXm3szF7njfVev+jzmztYhT
62WOaRJnFvctf8iclmReTl/fyfdzaOzFWhW1ynGp+v8VRfIdZNbCfWDXzzbS49LSPf8hdmvMZH9A
YJgK2mg+Cz+GcV8YgVIfd96N+CyPqSh8oXlGe2G/eVo7EiTouKm/YN6a3GiYw9GNKSWJ6D5Jmxw1
RDvil5oua99KvGFyC5MbI+9T0eJSMWeKYvdt15L+HijEaKQkuZJDbLM3oD421w3Bzdl5RIfx39oW
WdbR7WSD6pDVgGRiBoUQsZjm9cMCkS8QmmaPqeK4QNcjt6UctVtgmF/6n6Lw9M2fcWMb9Sn5Lfd2
SRcAN0qkY9sCBKtdeZsWfPqoojzJdhYb/8Bn76lNzHJngYAGD7YC25CTQGSOVMx+rtfZQjkG1B6F
o/g+BWzB9CUH8ckaWo8pdeBRSeaKWOPvifkBQDGPqHT+SRUKWcQjapROT4yIm41hSJjjMdOvSbt7
wFclWZapC0bX5RSFvB8xIBBTS/t5hIxVBQiFD6N6WGwsimhmNiOpEVG2o0ILJhaA/CBnBKLdfGTU
xLEYhFZ8L5bjbnxKgSQjyp3Nd3gaqO82Shb1JRPeIkpbf1cakHgndUL5nCxpF8J1aLMwTuJ0vIz5
1MuNgHUBdSfjsKX54iybweTIX79X8MK6Azz2u5h7S3dWBStc+lKCV3VO01FBb9UawljErZbm3o99
iIcFf7N/ciCBb9tF3/NR7UMMyAghkAdafxOHiwqQ1Au6nVb862NWhitTIckhVHKhxOehiE1K6I3e
is2S9djwUi3J2h4RuGdTioYot60AuNxRf4LvPfWR+VlRrgCMwaFGa+uzLbcFhva4yF36g5Vl7p2O
SfhSjroGeWgwUDlvCAsvyb4ivqiU5mrq6Sq178rmvqO9cujUYNmh7gHZJ+H5QIiDLMbpLyGaItlR
VF9rQReVSTSS+YSEgP5NstpNhFfuT4J4G3ya620Gx89/lRXaBp31ORui1nZc5C1sKG/+Fk3zHpxH
cjqfdETfwk46BIsGD+PKMurAi3dSrRXhT6gwVhi0ToXgENmYTfPmmFTOc6i50Pza5nQZ8UFiv6nU
W2c2ZDEcRLZf+nvgYU8e2lw59Tl2/yHLan6BRMIOySKhtHvhix+aBIMOgh6UyjADxN63GsdUcdHm
PDDgV89mtWjOZE4Gfr0n1qoakk/ERaq8mkeebecMNyGaiLn6PbCRsTGL2srJuahO0mEA9FwjWFy5
U5FYzk61JOY7wyU1V/0w0LDSdL/OJkrUSjTNCLYVe3JCYnUJ9loeqQx3rHEKV/HeUezntnGRw57w
5yNfdQ7RTqJeySLP0RM5WrbHru55b3Ic1Et1jqthJ2xJlZiAdAqyZ5+DEHeDweTS/hzOIn0OZNVE
M6ut2RqrM19mlYPrz08K1Tqxz2QQc2h7rkOy1NVn5dslSALwtT0MLXF9irtKgRcUtVSZbujgZw1Z
V8Mc8MkcjQI40nyMLTIDSPMF7Ei2Ic9ASetIdHVgq/GlkmzJSGmgn3Nourp1AE9pSbFReQXYpWVl
8tn6Idi8Gz4pivsPR0lRwtdNp1M+70oAI2NJ4jqnSH8BGaaWJ75SZlkYu+AKkLjaqE/llKephqbR
kVEFZhnH5vbR8Ven11O4KJohlkIAMiMq97pwZutvvkfrx4s6h8ykwXVhyaG42ol6rU/w2ZDjUbrG
jqh2gg8o2H3OhR+q7Z5sBqQGl54keZxSmstYBT6wP9HFKpReSfEb3o+p3r4G8asZNCbYtipAZCn5
eRzz8DC3fPx0PE82pl2YokcsPO77CyHdZpOSv7j38ewjg9cFw65vfPveBjIacwXPqWQIst25vWk7
kTPlwAn2R9AOx0cM61Wk4N2vyAxU9l7sEZSfId7IFflB2Nd3fWrlqsu9n1y62VQjiyTIe+EPpznp
eRlJEhZ6tPV0TuiOq/YEr/6Om9cS4HBh7nH78UUbSy41vzqzT8uDJyULk/QCN50LdYsYNNh8FVRd
uQe8CTehvCa3SmUsMi/x2bxXgzUOd/dpxC0Tkp1+9ft17q+zC3kvG5jJKAqMFKfUlKZ6mYHw+Bmo
GrmC8UD0lvTaTYJSQs7nT6LNtVbKve8DwEnfpG5BXUa5v/r8S/w1QGSV10nLib4Am6Aj9Wesyvkf
YIdDKhimsKF9TW5hQYAUY2jEbfwsHchEZqi7pA1+EcRLJvDGjFjIoeWXEbzFY005JAXYG0yF3K8z
a/95fX1XvBcW6D7Yxql7geICsNmUBUL2UWDlDDQTcl7Gctsnt+MOdAi7qA189GITr8mdyIHxi4Of
RdTb8rSbfTXFycjf9yuv7HM3XkVUEufqi8944bc61CocXaCbnEOr70441Fiv3ZQraYKrcMSboz77
5n5Z+dSwpi7hZJSxoybGrr7e1VZ+h1fWx7j4en+Nma6P4OGNNQtabWnpw+tKvmcsEAoqx4fSWGcT
jyBby+trbZHDZrXmJtOBmF0JTOSZe59svxwc6D/B+byd06aS0qudF8uFEl/kOsicB0QzFjNEIerQ
RTUpAvOp+4igNJykCf+KCCUH0Fx800HFJ3AP6zKJOjcfEWxBr+WXuz7vclxQroF8tYJYumfLasud
AHTCx6ZdqCp5zQGUwHPpBH3WnYKFbJ10i1uHS3QNG5pJrvtJhFwn11lQJkivy+KAjYppprifKN7W
h7xj/vxyV9Z2N3yC/p/P6NYlUwRkH2VEe3jCvJaaFSggPOvWcy+AV4xknxUorDeN30s55ASA1bBg
pHpaE5CoKehK0fpLlAIt6XRTvqN1QnIl/+YlPAUQyz3x+PhZHUU+N+2g+V7Gb9yRyA2Hz5+i6wxz
J94UtUiHuOjDjvCnQx9o8BZbN0eC6mROqZ4KZbf+EurMBVS+I5JIhw6/CqtmNxoo8hHYMgEpbw46
YwTKy8s4Mz0tARvcHfi4OyJxBiToaciji8PootNGdpgViZYoFUQrmcQ7Ap6Zbm/3nR587X/8QoRI
nRaacPhJ35UsVCF7iwrD8z9enxaYZa7iNVRi3On5SEVRaOAxyT4O+ztYQXJCKeywrQMZ1Pu+4kGP
cjmgnmoN2epWnoAjPdTOs9bCGkgpmnIamc44FMhBX1O8SHFkscmpJKw92BlitkRRhFq7SUXjq3BI
x2G0JiVPgrlNoCJLGJ7AZBYF14/sRRb28drJP/zXaszbNYHWdBYLpP0/ZE17BtxZD6ra6pkVlGjk
ptAHRFO6Q6QMzyB60/UMdlIRWHmTYq/6fPJtmbXnlUigwvGJXa2I1U6lI2Q02Z7qqSx0QzCQ6g8H
uASDa3HcgjDarT4ENPu71L8HobciZdlLxkpIkhWBYUyxzuF/8cluLlc70DjMTPrGuTjt6GB523lM
XMCKBV2nPh8meMWmyBR+WSdZZAUZyhSRn6h6sMqKTllGWW4TAiNAEbUwVafaaNnJr+BuJoFNdBUg
wnQRxbaQjWOL9wxrlsG/FMshmjSSKY3JnKOgfpIHtWbjY7ZlwaPDYaC0w7libkTvePN30qstrjyS
nx4NvTD0hvkE5n51mGNf47WV2nNELXsU3PsrwDkjtzufFii3SI9NUTCtQeH9NA5biXgGU3vhWcae
/NelgtCEYxcFV370N24oWV+VGCL3HV3UU00A5oyvHrR6yqA3kxgY2B6oGki5fiteX1XRF06E4rxM
RLiJz7HkpcV0hsNku2gJULYIUPz0TcoRsqSKp1U5DOOMpjZZ0hiHKiLnt6D2C6gDS6ET0zO/+FoT
l2lOUSI2EWtGEDnNucSinEdz3tTNDd9c3MKmGvZWjL+ntYaJg4sIHxEhVQquCsetWrtkS9CmjTem
tvgtbMGjyV//pCZEbwg87n/ionqDNqZA2gS4dKDB5q8Hy1rRGYTnFLtdxiP3FWlb/Zt46r6YAzs2
U/U8fVngrfdQkEs9fcSd4VaDcgMzyIgwrNfjCQM0I7T/KI4lOMVG4JlqiZftN/T/bKs17T4AZYg2
p60rbRqY0ZFdKh1hc8hYZBdI7SkZogxbSDaigbvQs5ZgoF2mEoex8teHe0UAwSPpbXgOg44LnXv+
toa+ImjLYF948vkrrInr5/m6oYBSdwg9xd/e21rTFzZhEstSsOiUpREh7YzFkk3gCofHZe4iHPsS
N5eBQ9LgD017Cw2L/Ga0AzgH6DZgTMLrnioX2NFzQKoyEFDD7o8AKJlbyp99CAj1OnQMsS8yglGw
uuUgAeyxEcIc3w9chSrEjx9mO6uo1qUMB+HEqx3ZL+PyMszKCcIRAINzWzu65spkm51Mb5PdOU4C
2DVwm3exANc8Qt1nsn7/B1tjrkQMw2R+uQv2MXwMnKM3UbkBE/hMpJ2VkHB5rN6sh5lrY2rMX28x
rviMQTH24wJ0/QjTT2yJeHWhR6VM33+BJcovVefjV2jRRt2bx0tXZJbbGV5Ux7i4+IWtcXg/zoWl
83g8rd4q5ZIw6ZNLQ+FNy91tufCua6lRCuLEwhiSTDnvJjT0SU6SXsuKkSLP5v16jrTkwG+5ue/+
COMw3Kjno0HMW7UvJKy07CDKnxedcl1EoeqSE32jUh2d8EWq3BEkViISCGV8mn+GczpYw7XNhdnX
JcQDnfzj7d+ZkmwRJbeN12HlQd6Jhp//1ApmRNP+Jl3Zs4g6xnUXf9hjCitZ7BV5xbvbW6PlN46f
vMJpxWEA8XnVcpY78PK1xJjColHQDs2CBgszqLs5SZLEWUx9Jd4m14V4seNaEmLedwBBo/oNWzEG
oFQfBmxDOdvFvYqxPq9+Dh3ImjEFvKUIZrX5chaIG5257oYqbdFHU/B6sX4I3MAJFGIWQsGUgtiY
u2V67wu+iOLxQCtfcO2LVe7D5aXBFF288x3IEBHoZH7+Os/150n+HhUAP2JBoOMqxLaAkve4XRzG
BtQ6VxVzQ7nAr6UH+cgw75ptzXlpkb4JHihj0pRfNsdYxbLUrGcStCI3NN61OQRRJlEMvZc0bPzU
+1jSIs4R+IEQkJxz8bO/LyZ+h3/x6RzplwX5xSbWYM1fkBuwBbGK+edHte7mrzSXEY0Y77dr3pRL
iyKr6+kl7fTfo5Jg9xm+Li3PhPUCVCHBCTJuhFn3r6rRcAX/Q2FkVDpq00uE21+53Swp8Ne1AGwG
t6O+00KH8XlBzT4/w69tuEm+DPa1kWyknIzE6fsmto2E7pNozKms6QdXi9047K1CUi0TO53bdgWc
N5rhMv/7yHjLpzBm2tH6yAn/ZJWB1gdYUP2AihNdcvpHuFb8nKsaBJYq4mBb3ZJNEhTN4MCm/nfp
uJRoQiqHvO/Tk4GkeQc5Q4/aLwIU0UHWR7UbZM3/xB2rtRayMKyuoyeh34jRlN5JC6Ell6qBN8uH
ZgcF4n7R7zmZuUvcftdf2S1P1Rvvj++YFKvokknnchtSNr//WS1mrkD7TuHrG5JIDA60rmEkU22v
Kw1xOR6owFkB5H/cbGUgCVK+CF/YzvaZ4yD2fwySyYDMEQCv8swbaEN+yCDHp2T2O5s0m0Uh3j4b
W6iElHURbcFbG/n3SMbfUPpRqP2G5r6lnsENCmw3fhSb2K1BSjrFtZXeW0gcK2PMyMM1KOTbLrMk
S/8YSLoIPXcB//6NMLQZO7MPY8bLuVT3ZebKp9ScTcxNN2BW79Ne00SCGK7lhdNzFvdJEYxgRoyz
l3s+Oftzj8VKdFZG6ehyCtJH78SADLSKEjtbByipjjo3gyfRWRpUPv+++OdFiCoSLc8ElccX8Za8
rgD6Ntcv2prtcUcfYBk0ulqyw6Iz/lleJ8Uj9Hp6ISdnloiAjEByWV3hgXSBM+1BH6lZ0IyNaWTV
CDGFulqOh6V/u6oEzMQlwt8yyxqNaIugemzik0EcHFQLi5p3sR/ZmeBlrp3BwAW9sWlSiVmB/EFr
FNMoEyqfV4jHXm64MN+9rl7JtHvhUHr8VknBxUQi3Nwwam/MdcnIx+DpAS45nA/V53twgzhnkd00
L+rQr3ZD/IH3BzERjMrilbqPMa86obj8FriLYBbjiOyI7mYxXyl/q65KO+DoKu0z45XsGVO3M9M0
0vAujTx9WK3ef9I8+oSfht1mo1/Uwpa8cnaJMHw2WO8AYUMgOWLO/bbLqlAqVEREPGTSPuddvBAX
riuUSYwT51TRQMCp6JlbARgCyx5qGmIPsno8uMGNRZNqJ9JdMA/N1Snd3deqRBKJ/2FHkXHlsoQK
tyD1v8vdCATPv+zPDibCUAinC05iwRd7zR6yokgXMY9eaoc8Vz0ayDSzsgCsXHas1yR9J2cdNM8a
dLHwOf0Z9L5dttN2vHEP5ZSoucQH6a2K/7YpdYFdIITsm7GYQspNcKxb+sXdJ522PSVmW7T7jsUY
f8CZDJCovK86t+zLoG8t+8tsuzVc+YbS/A4/uk4/8juKovKz03NCt01fr2xEg32A6WKwxXZq+Ev2
zd+ddwcEBqfmIgy6kXq7rmr2ziD1MencRawcfOABvOM9R4Pz8vvw/yR+hTm6OEbX/HSVzPF7ElA3
jI/jCYBgwbLf+GV3I/oJbKLtCMUG6Y8fQUSa7kAGBgKwbyG2CO9YwiSLkVwZutMon5+ESb9XZUOe
ziLso9lPCqhtqn+l52g5Hqw4UapJLpUqra4pR6lquNpx/ZH0z9jgg5bvEcJt+2Jc69u80onh1Dqm
Hv/mm3LQB7JisiqQKp2T6Ri10rHuZqkulBAVlocAgkb486cAtIXGEHAdVRxSGVDg9rJ6uZZyVtJZ
rjCosAvjxzIAdOkR4zaU8Q2uy81NXGm3MpEPI+N/w1ruRv/tanFDUEFT8boaji51Xl4Yn3euFHHi
KWCsZfrwC+8Lxt/F21H39vyrbY7DABxM9drLg/RXOGkwW85hMtHU5fKUdQgPaGzgZyQ36u6CZNEP
BzAd+2MkAucfCs6LiUVH/RpS0kFKYKVRYwD6/f4AJqwYTxBVzD4QM+NPRCvtgV/dlMqAXFqKzIhN
6+pgk3OcQN8h5GmPfGZF05Agsqnw8Np2OaeWdWFLvcTd66mIAG8au6gJkyNvkVf/iRA9uiFXwxRk
b46w1D0AQno/fAS5LHaMpk9vp356FodsVJxzPynDKFfImKtzfE3t4s+F80vYZVh2qV/vKAdk/0u/
J39DQ+PJZr1X//5E2rWNBpix5T0U0o3dSqAMitvTGsNVCNJz2+6gNPBqDXP6y0aDzFnJor0q1AM3
Fodp3RjdfSc2xSFJKgMIk9vS+X9GhIPjGBPqtqr+KLplhOlPS1Q0tDsBbutsgpjEUfD/hdQizRWr
ogqt0xd0tWolr+6jo2S0muFJA1S3XykFPrSHVazpQWM9aOWsmBtGRENVb1FPZesvh7s81uLUUFdo
hQWj3DdgOHK31BdzgNnt5UHsrc7A8DN6anbL6ki/qL1SQpZQscDnUbDqWyO3ymfiIInj8ibdfF9z
KWQmMh32xDi4MHimD1U6f5PN5qCHIIyPN7IpWB/puDspChkgxr8ipAyvfeNU6ir54FKEO5UAHpuG
XrYwbZ6vuiu+YrRjNstInO9g3iOPiz1AtQeY4iNMWlEJjwthlOpQrw37mwOed7yIQSAMchi0PFeg
fvSIEpSk2UBNoF2lep8oRRGazCGwBoNyFanhlbXhAYxcexaR9q8GsOnTO2iPBgcOoMgzUZuBNZEk
QgUd9KrBSMHiBdbRNBXhq812Os9BTb8XWrbcqxVibL3Is8EDjVwDH6mirAzOXWUPODDWLXQzylXc
fCz4vSe9AKJCxu0bjXSV0pJtNiOgHZIVkpnWKVokR15YyP54ehjnB97fjHGQz7BTSuOg+eiB4VQI
bJO9I7t4USZwOuew27sDHksfVKWzM5AZGFTwT/9nKdNgD5Kv3M6Y73Uz7f4i532BarBYFQVtztcL
v07YtL7URVROxNFQpoyiK26uVm4quXLwyjhvfrIp7RW6dxNDyXxpnyL8eQVk/kgkq+vvy0v2ZP8k
xFOllW30sw7EAQHcV7416H+5shPxKbZin1uJg8JQSeCklclCCzq/PJygHsKMvqnTit1LNVB9CzJ/
MWe8VWieOe22bJm2fu4MT6x9pQt9KF5YMXd85M/s72GToQkeZ91cePMY7xPL8PqzL8HblyPPxnVh
8Vt4k/Khk2IdoL8A0XfSRacxnfYcJMNM6EhABlubQk8z9aPtlq1BMjbfwwaxKWqDDK7L4Du0WPjd
1GvWx8MSZrOedeJZhRRbL88DPrS0zh/plMqz3KhKgh8SyS4dtm86Z+bDgDMlCRQ8745rTvqV0Cs5
8GkUfIQIFjnQKf14FbKPf+VBRhG1tWU+AVlQGdNnPoWkZf7EG6dOwKAAF39Z7Iekw8BlnQuSkmj5
5NpV54i3Bw6D6VnkjA1OLVLp7vApMu02j5N+96y2pL9biGt7xiBzi9hw4WQ881Pfdxdl19hAb3FK
PT5SvqBA7Q7z1rZfUTq6E3fl/wg0c1z4nvm/tmnuM0cWZkVgc/CCj47++QDIbXBD9fiXKs4agzy2
vUpQHBZ2j/TTcp+sRPPUEr341aD6WZ0dAg2UvDrpdPaS8AztyafJxlQqbjwcgG3mKCumzlTFFgpB
ztJF+U6QTjPRdYYh/T82h51pUEqMLejHzaRKnytiCrp33B0Fi9IW8qH9qr3m8+7NwIaVIOGWAgX4
JSb2l4JPtLRzYF+KqqEinxlMY/yVev6LkDmGaEf+SCWtm/RybiP+Wu+9VTLdL6PxgvZ6en/CqUt4
zzTYHldPXeytsN8OkFW35VO53d8KUpmlqwzF8APShm8SGMrhIYvyTmeLLaHiwWb2W7AUmGA+rQFI
JOpDgyJeYYkVSUAVLDLFcq5DxNtT7ai+W1qnZQLRPitAxCXT9pEOyNqnw8XDYsB65h1rlCuMGsPN
GHmTR8uZQq7LZPzMvAjKK/pxUsDjZJfw5EI2VLBbq1qjdMMffnyb5jH8P9ZN2TPQu9HpkMVMMLFu
mnMD5W0ug0D6FanKpdZM7vZb4d+SwlGXgRQ34lFWXn43RSvt28oHBHWPSn8FFeFlSthA7/EH0MNW
YiJl/wmV2Rq1X8JtSxu7T03n5M5LyWCsZ0gHpnTgj7UTB9Q0uLXdiClq3PZijYKVMAHtDWNkvFNX
L9Gwty0oTc+kV2lp3mdgTRac/Un2bMlMKC+0b0D8wXe+3fjB/631LBXmQVo8hiRr/839T1Slc8X7
+y25sClsx+PN1AK8UY9aPKfjiLWI+eneXM1vj/rcK9o2GmfNg6F8zmJugBUFQMWIPAxId/udGFxA
wxzeZ56YWeyCTbtKNmwLQiSIiu7atJtDg6HkFbKsqvLHac8Y/LePB2uAxDbBDYLstLtZo5YtKgSb
Anb53cxrL/PV3TlqGjL7D/WQdWMTTJFR/MrfQG/A1ClhbvV4ALZKnPcG+8u2swfzjPHeMt3bZHUU
+yQTJJbPpx9XQBH4HrgXZa6g7b4faHaxNmmz1JK3coA1BWSbu0iRbah0yPcg16BB/3fwM2MpSX0Z
naxQBruquXEHjLeljXP15Nc8fadEmQbmNdskwjKv3aM3w3N/zjQnA6Qmku5GmJGBhfDxU+wOrtwH
h9eTBZgMvuZaespUH2nG4XCpjl2YrIFRaEQYeRvzFegO3pWu4ENevlSGwbefN+7erzPaAyfyT8vo
z+HQLOqfNiNZW72x4rs8DpLy3T+ZMZGP/rlAGE7LB8NhrUp17q6q7gbcEbiXGbYQPlpaGiYaE+zw
jjsu17Pvv1mhzFicyZo+JTp5mfmVO4FxK8Hfs4f3wlGmXmbiAEODWG1pBaZaIYcpQGcrOCB8fkJc
+JVjIdSYluRwNBVx9XN6dEq7ViH4vbdxUZV885P/Ok2QaXFwkqRwU5HYA1kPFIFfOuwLKhDq/aPA
jD38/hM1nQEhFHZmRnYtTbYJajreV2QBZO9kODmvkXElDz+WZPK5tE+l0SIc1nOuM6qablUBMMBA
HKCUh0f/QvRNMfJO5KyJ7XNpTeF6ieDn9fR+yf9P9P7cKL/gHsTKZVbeI7qwqcpBKE8RWWeD8lzh
kXczLdYnvWAzVMqxFnwSVPq33wjOWsJIXbFgk7JELH5dErTKNkFliY1bUZQQKyKvxvO/nlo8mjXl
GTN0yV0KMoP46YC6nU6pu4KeNkdFskS67aPX79IHumfBcdCgBXx81crFNkW0wltr2or8BTzJln4O
ClYIyWyHeGACJaOGNElkcpVVjCkdzYahWBoutV/hRPAtjo0JJMaHDtjNKkGikBL/x5ER5Li+150P
90o+lgz/2wTbMco2M6dH8l4h+Smw52SA6geTI5Qge02TLrCfmoH5Q9Mztubfs/VP4IeSPc4R/6pL
LrKyiNp3ycx91RfcCvSXJW8OXRTybG03lDxUoVuTU8m/orhy4NSzm05yFcE2sYk0qS6/ytW+hw9/
0alBh+nJvCiy2Cvgdrdpfadydy8id+HBhyCiYEaGjVs0kBBPgWYioSqJKMY3VIsi7+tn+BctASa+
OS3TGWwzGk6nEW6SNbxV9kkf8kCqP6nX/gNJ02ZvEQUY5j7fta1tD4jui3Ew/5ceGDRh55SSXWhy
UsS1Wa74YXFM3AXfZrjsnzEEh7UZBmtZ3l21V7BlF1AJg7azW0wQLR0//8zgrQ4usrW2cI74Qc7Q
uzXZ4cGtlT2wdI4afQf34URT7lq9G6eKkklVIGNq0tdicON9ZRq8JPnoDQnvlikdmBZU+SYB5+yd
sZkt8Jear6v3m4u6+qPEBzhQQIWKPkWIU4YogcSSnXZbwa08I6IlTatR0wAS/077YgnwXXJBOF80
/swlEI3M4dxsN8Us3aXQAtkR1RQv3gcaQDWSkhFMM9fEn0U/L4fOL5MWV2GFScdL4KAPtIi98sCh
3yZIYtisiD177A41gnwjywqiF1SwtimysGCrP4fMec/2ZHttWYZ8WS9ASSpyzf7e3CMXh50Xiqk8
X1i5GMfUspIpqYzzrNO0dFAevf5qpM0XxYcBm/q+HM3AqmO/dvY8gDvy/N6Lj505jJuh9dvjtYUo
KeLaljHULWtB/BdsADGJUV9tF5X5jmqMGERO9rmzLEH8UDJhgyacvmRZepcF/bNbSgd8StSDUMKp
1JSVmB8A9CsYWIWgEUU8cui/MYf7F292gQgUddE2w1OU3CCu4+N5dE669iqgXOx7lrB0rYcg1jn9
6XyBYur/XgvlAHmVAoxZQPW21t72zKvV/i9HPGmXhtpeRKCEKpRxEnHwtuZmqkLnDiH7XxP/6k6Q
h9TyUaJy3zYZICodLxl4rciFbhpOhKJmR7BIpyilV9amb6Pu1UfcqkXJqxdWu+XlEyA6myjhR/oL
82m5y3rsZmJ3nYk3I08Vrzol0zYDcuanQUrs7LaEBsybx1xTUooXL2vzk4JteXWXBGlwpHwDhfw3
PrFmqzKMfDZ0mnqHiMBymzW9RjGN2JZcCdxsQdn1cYGQGhN89U3FTYqP7GeSZ/aW6jImQtVdk7hH
Sz/OFIDuYmJT3mhelYqV2I43sxIZ1CNfXssSW0msUeREqYJeFOWjh7/nVDYRHeFQo0qLO+5dHppC
2OmkgRdW5kTbvS+lp7Re+6bMyG1pz6qDHKCGF1byw5OdtdhLPQUSS4KpNS6VgA4kI5UABlNilGrv
Qe6bXNLGdNonUVD1JWNMlBmq9D/9BJ0+YXN8sGoKHUN0pqwwWb+nu4JCHR8gMwSv3uMV2M5AUkiG
T5VpbA+OJeTk1y7pDjHR+ghMWZRQuT5OLRbADPGKoH8ZBPeUZp9mvjtSaPNxPRjGfdrmFWqMueA/
EzQL2VIJFWSX4VMYDx0OZ5UBhOorc7pD7ukxnBF+s+++a7Hr04XOHJ4m1hYCs+8QHRO0Nj0sK89v
dVCvnt1AWNsHvBY2ErzUa6yDAMtx7T3F8uYGTt97gNbHMxWdU+ykKNScEzF5zS6Le0Ro9aN9kONQ
7SAleP44OgEYDNJt9xz9utncwSg3UlgKER2GYDLqQMhivo/36c6QfhiHxJ5N/ET8yyLsSZQVK4QN
ZRbjU7vJ2UfE6cGHSxF9B4GExVYvOvX4suhWfVJ0UW08xrINtzuogWJLc66fe3rhE0jjI59uAOnY
O2E1SkPdn+L4vum+o9kT5UnZwrlkJ+zmZUc9PQrMEkGB/33YDACZayXcR1G8TxlD5cBjzdh+j26E
1jT8bRm+p2n8eqrBkqxUm6uX/0ys5/fHm3VFf12Pb2vfi51tMLFnrvYT8vV7HNDxkaWlKjfFIPQy
/MUuKYltaHBwEpvGKy2ukotRZGqS1fpORr2ITawbWkVXbxK1FC7UhKN2Bv5ynfbHJrTre81csQa+
GJD049SyYnKJZK104zU/RevGux0Dh3QTjeRsko/vzsyXaC+5OuwXkbAsabvQyfVdr5NgU5gF0iqP
OR/fCxrGscWoQwLamrfLziuHg1f5RNs3KCfzBm3dsJJwVIIlssRYATu/xG0j24FvFyPFuGNtufCc
DVB1I9y6VNjhD9GKY154mTAXZIz9lZ3fZRWQBrW7kcKbnHXVmCCxUZ4hqzMTIikQyJgvcIQcFP0r
auMafpjOK5arKaB1RyMkc1WnAbGk/F1UyeN6sK7to5oUjF1VCltCwinrBznfX6NyGz4v5xV5u/KR
1aDakn9657MtJd7pM++DvZU84frsKLWAU+EJnhATZfRa3yHm45F0YXYhsx4bstkuV1SbU0fHKsxS
d7gABwy+0Gnqx90Iytio3gPYG2qgj4iBZR2eU5ewsMCCdo6qlIttzVo77UrIfFHXHwqURn4Giopo
R/p3xWu8I+6Wh7kDYhNHJzWFZDL8v9uh04g/tF0v0bU3KKRzVkuhpQJhyHp9WX2p+kI1BvNnU5fw
d7ei48H5jNR8MV4IYVkbu63DVdOylJpd4RjIv10Hk5O0goK5cVAhbE1PnCtlaItlOHj8vfmHaCDz
dLyeHwXqWnDwvQkPP2pJ0CybUzwjNIgqw+NjbNEo71BkiPnPAjzjLH2fhJWvxouCLwLKRvntmMfZ
hgPjV6zJ/ojjDeOUvMW/AosQRbaNsfAAI3NiTA9mfR6I5SCvugjT8/cnqJpYtdhbxmXWMW90xQMz
tI7qCWAe/cN3NqKH2UXkIZiYNtRK8TAIoAzxDqxORXZ6EGC1dMWxtZ1c2ea1Z+HP77ow6FfFrBJs
ANmgZmihe8KbYurUMTh9e/acvgfyF+/2lZpz2/V8E1mLN2fmFAiy+/lGrv9olSBOqV35jcrHV2Rg
luupzJ1kJ7SburVidu+1vGMK/o1qRjnyl6MMzkKXVudSw/PESx7n6ABia5WHS7n3/jupvb+vM+d6
F0pNAPNlNPQ9dYdP6KszB3h2KQWg9/4bIA2WQFg0Sg3YorLWQ8iqYBdfv6gxohUmPpnhLy5BMIMd
ydh0AyHDnjylNEWBtpkDZuVtajYuJ1WelU+tzuP2ObQDKrjb9KsurAJrwON3UlanFvuLBx+P0Js5
7Q9BZBRqDDkO4zrHNVrCq4MQV84GetTDUpp5K+Bay76MtMNA9v+RepFFsKLBPpXOOCGskuTpK0Wz
OQMf0f3qMUjmTHtUd0bBKE5exdOW5MxwEgWFz16KkOsXPI5R+/jj9V4irJQyk2VbZ/oJ8AxFgEZR
AHK4EoGBqw/X2JLYrdMogzj3pssMnvIg9S1Z+k2RyOtb2ZVzhh9wuzboAkCGDoFSQ5zsXKHMOKTW
Fy10EMyvchdyceItSHSjJzYut5O4Klmw+ofL4DjnyiZphKlygXiTUN12PiY8eBfRxU5ne/0NKieF
0kcRDI4BNWBig03CGu6rxaw8InrDbBazaMuka0tBL0uON+xeKFtEfLbbG+7DyBroGwnMSfTsBal0
ADzaYsUCs8sxfNCW56qhf1ljh6W7YXUVvTCtc1pv83jURa81aeNeLpHq9yW8F9aUSL36E50NJcAG
18lcTgLCS5PuZL3gs3jQcX34b2k3qEwty9RbrMkiGBOrC60a4zxZZ5WiA2zRDOOXMW0LW7eAnGnu
D9MF1XyKQRJkjCi/kzxdxv6saeAIcbeSo6sunz+J/sps6fYODg1uyQYN2FyRzyRSHJSgziERT3kt
petLzut9PHYY1OlRJmvnxzGToY8fChrMAW3D1sB7pFymiFUB/JC8MweoxtyMcoLEOovPbC+x60he
G4vIUuTwJ510hvMfyR+0z8HB1l7V5GVJpT6YvgIHpel4dJF7LmrpEjOlXRuukXO/+cwsYLd22FYC
PCGCZ6k9Dt1lNsDb9ElmRPVskHUHYgvFRdo7KrRpiXIX5UR5BEJLrAypcvkmwJS/6F9UjG8kN8V5
f23Jl7gTbXRq1QhZF/9/zGIjyRujiZYqDClEGjcYT9EjxNcJbOIlndzHarxzMzeJhc4ClFCcDHe+
CEkWMddl6nK6p4HzgA3H57wrZ94iMB8KgF7Xr1G5BKCW92fUzjXu+L5fEb6xWazqhUsLZ1y8ok9Z
XGv8Ojanv4fPBoDLuV98+8NPTLXESV82HXadIOqvRcDWzo3fdrkG4E1ISOyGxspdzcGcGlXV8C2z
/UVZ38aF1qmEhYaQANuU2IbtHnldMTYx1rTsxz/48Q3fwShcUtx5CDl6RedhT1NUigrYu/np6G5T
EQVQh2pCymnOIUYXxV82//wUtGOco2hNCrpkGB4YYJhuYWJkYla5U2Q7ApWjnzOzVFgWpHZa6sAO
XLIr/M8bEWo93igWUEubTdN4qRJpB3XhTFJWfE/uL2xvIV05AqHPtbXers4aK0bue4J+pPSXZDO+
uVsZRRndFGOAAkOV5XR217NpU0B2hiDnPSE8eLuNMnY4jbu1jFbhemfKZheBbn1hoYvBw+B/zjMM
ZjAd15Gv+ebCJVLmMcCA8jmeM33sp8tGZtpyYkkXRxuRwql6baNYkCEKbvxu8CsP8vt90tXfRADi
vtulpLxy8l187PleAxgzOzsLRQe4jyZxf7cBe9cvd/Pz3GLb4wkcMWEJcfH/zHxCWMQbs/eorAWc
zJAbwqMXOjtpPnVC6L7/A1/cLSgixhhZGqJ6EAzjIBy4LBFcDVEAfvS3oMxY5DdMOH7dpQYWCHqJ
qTzmMMn5yoZjJGrBOPr6ExeOIWtkR//sRb8SbE0+4JEy2Kd9kMj+Pob+NEJ0muMUlMJvl3CELTPx
3WQRa5ruNAXfKTyVAEN7bHTFgg1jbbuAIja8qZ3oNxdL453XvI/7lZ88yK0WLYgL0Y7e+iUlBw5N
yAMuAstMa+pK2bwEyfXg+XhFytXP/iDHmUbrTQhx7HXHRqwJr2KnmE3i4FeZ4IfQDsYjQl30AfdC
hQTTlBcSVelUYU+F896JHguyHgwpvCpgAnh5vjCCvjXePAjbrbEIx3U+/e9Zio7pNm8FLmx144PN
jZtJmuTIR3WF6thtJqhhAxQIvd5zz8XgaseH28l7+EoRC1bQv7JZCNjr75YRjcixcmhxXpz79Idw
W6gD9T5N5Yhy7Lqzi1YjDnWr7K/TA7yeGqn7YjMoFq9nIKUfjD/sBjO93rfzgg8U0Hk/x9kAnkaT
Y8XCNC44BZqU3GYx6u17HbSjB+hh7/kUihlm0z4mzELEh9t6uhmTZ2Crx4IpNkWiMi3PT4z/5Ny/
Timh9Voxqs229r4KMXBVebxgL9xwIs7Yai3YPSi+8/PNYMhV5JPZ1TbkpVwbfStnOmQr3LkYpDe3
/II9yAQEDpmmHtWXgn4JnrZ8ufyDuSTv5lc0egMYOwKW0XwvR+1+rJrtoIl8k/XpL7vZrDuUqao8
evkfvQyoA/DaAGYnbrPuVmO+BRAVoqkPM3VDqA10zQ+OWqory+ldB1Mfn68H4IZkCK+jP8xUaXVt
cZFRGcvOOuj5NBmlbz9Py5wyyRyUKTALrZ7IJJhwzPjdQFc9KsJRUu9OElloM1aY7lH2LpWGxR1T
z4MCJHb/kqjZ6/AYw1alHGIVOD7Mmo8V179/uapRxWMZ16LFmgaXWbGze3dW32ER460+8zkVozsj
+cYB9yLuR2YVnP4A3YTLok0s7qrWeEQ3zhWSMc7iYfofnPs1pFgf925ImnkkCKIxyiXkpgvH/cVO
I2b3i5jeRFCd+nQYBWr63082HpHkQVFZIJfWQs0ZkwI4U/cA9BfM6TzYqy06qA03m2N9ylaD1zds
3Mr4Ya56HGYZPJe7m72Xr0u36mFPVdveErffQam20b8k0pjI6l9eVMa+bgesoAE7tjfTRePDHLLO
nTsk6xDJmDiZKUaJoyNt+BQXQOQ/dsQeC7LqVOVfVNrWwtNdJaQmK9QgUKLdrDb707Y4Fdx5awJp
8FIvVQvfnW7vWjGrHQfsNdQbhgg6QYcyufppugB/dXP6PF98r3yOaUkdtHIBVLBH2Gbx9ojaenoI
tTsnKTokNCw0rAC70ckJVeEKmOq6mHkKgDIdvSwh1hCBkpLDNpHxxyUM2SqIZQeldy41YEjLKice
0/FWjB6frIIhJOyt8zX/zT/dtLyJjCBlUw/c31xWMq7bfrcrZhx+39iFVv503hDI+xQkE4zQbAzw
68c6CaNwaZZ6PCg0a8cUJB16DXtzu3veoJtoewCdQhXd3JWhsmGfuiZGEnN8K5CodVUJdNu7WO54
VhwLfclL62vKo3hAeqYN0pS54P4wFpMbshTTsy0t6GFZbFI3XIFmlvrrrLBZExsRe+htU4KoYa3R
fnWUVHE4cy9hrPpqAE5Eeio5KWanKkQAXUsBNXdudJcARriMMOjap7pAZDTK4W18rACgzd3jedQd
RLzhh1m9q/KP0RH/25hNruUq0jMDwsKzPcqR5IUbYTvn3sYJfjDhh6goE6paDIpM5k2dhoAY1Gc1
b2hYKg3Xn3jZ0I4n4qXdsvFbSld3wRBeA1QA02VipCI70AW8JCTNwwwuY9dH9t4xTN9WIEI3FGaG
UT3CzGKI11XDki+RhVaIApaAjKA7JFQ+8WTl0QITidm4v9/GyGF4m1RPqOUY+pYhBImSNqD/e9Uz
Y4k1ZrRiq89E9UITvtsTfHPLVol3eWYSQPkpL/r/h5XL4rBxt4H9Ki6owa4D2gdrgH6qDrPVFPQD
fN4YL9y41TJ4KBtYqoz4qvHUpfDT7s2Yt+iYM2XMPHUYKEU6GA7EBTqZP1GCoE1Yojeu6ZQPVzrw
aem3UYpa1fXnVpu8xqYoK7n2aW2yDeCsxQd2jzBFJq1lIlG3JmD0buRO5hXfSTFnr0Ghc6Ovyi8P
myOL5juDuUJjNUkiEVwBKTt1+CgZ4fKRDh+y3NCUBJZ3c0hjGz0mLr89izu0opyzQlDDCuz7dB0N
NsKVICSxlgzUbGyxCkdd64Dxeh3l+4610UTqEG3Jh+2Yi9f1LxOAvoAzCj3F7XyW/+biYO8ZUblT
AqN2HrdWv9tIsqhUz/uP79f5K1D5BhJtd5lcQS2t2a3GsABh/12LEtLtFhbYAPvhhEm29UnYUjHC
FkMlYTgF/LcN2XeuDqtuZm0yxdAA0N7cph4VhGtqapJlsTgmRfScKCRrR5i9d0bIc9GX1FgrqT+D
yKX4ujLporK5zAJHYMkX7n8qYFM3u+hAlAblYn1TF1DdnyZWuhgyB+G1JTN6CaeVL7jw9UaodATc
JEuCWEWYM4dObpi64gCtCiKSlr3hEL1Xx4V/ZzJavoZ+ljl3LiQJAp8gPUfWtDGnej50ydrmY3vI
d16DJhaxbJdLA7LCYePoeIwdDnAYyRZ7d1FMvBWaUgbHIlPMirFo3FT0mln5BESHd7CaxOLL9AMi
yFziIukFxrsmCBsu+mqjHHLFE9gC7kM0eKCkUhYgrwycf9jQV0xUQnek+JqVdlvNlswOGKDkkBVY
zrhYAmwe0hxQtuuDf1CauHLwxusjYBHkPZRwP2HQvDmJ7LoU4+xfC13yNGmqi6a8Tsozrvclet70
RzOG4tw76RmEG0X86OHkfbtKPbbYZQeF50hP61aKkQxlKozMH24WOkBVA5LavjGivN8UF9EDMY2A
zat+xcBl8vfoMpz+u0KMMuTdArOeAxpCRfYvLNit2RjemrxX6B3lQ3K7c8EFfiGT1pVhz50fTDzc
hJgJ4PQoIb1vIyV7kkOeFKOSEm/5WMlBw+x7VgHjc1M3DkU0SJafeY20B82RiI8yd+LigxmfGe3M
QnXWcRJtJ0IY8T/gbKVmIZCz+Dao7LbrBsbmjiFmCVg/3FQChmnOPuucQOaq4KZgGdMXcqF/z9xl
zHFUJsUnuAaYCBXrGwvlWKX3Q5Y6h1LZrcdi47QFeXsnG+2EtCMkoWymYNmHJdxt9C/4Aqhao/tP
aZxsDxM161PKcr4Il+ygYf8HSSz+/QXCxpjs5buMXUSPaKyY37Nu+t7vteYZE6RxQRCjumYbcVnx
NWbGNTosaZZxTjgFBCRitaka69KhFADsAOrS0YIpYg2QjB7Dh98M3eYXUditYI+zgY5NS3SYKXBz
wiBk1wB1PfAqiondIngLEf9CCYDYvMnR3OqJ6+GyDq73GzCCVLMGGn5bVbHMiebCSAml0fgXxDn3
soq/9ILxf4XJ3uvVgeTFhfpaVaBqGHaxJTxVNznzb6+8sRi6D/LTwhz+Ss1UzxZK50hmg+AwTGY0
YHzxF8jvPSmXB2JptU0TzrSLAGcSLde/LMNWvnOtsf0cyD+HnYrY0fjVoletLyb70BOFEY9ulgnu
FC6Ddy1MJKHF9pcGkq49hW2PzI6XcJpUYIZKPbQdrBTaFwmmchEMpNRZWKwkThXzIRJmfmDVJK6o
yfAFOMWvrTqtYNGbQh5sil8S6iGcOKFZyhdSS2gy06rEj01I7SmBfHPf0NljISR8mUPXb3EXS/yE
kivPN0YcVnPMAj9EFFnl7AuWuZjfboOSjWoeiKWzCWGloVgHLUmJpodtGl63ylbhWjN+i3aBW7ox
yBOIW7OyySZOnrNuEdollurPHjktDXjTykL7HhT8yAmAStjQKD4r4L8qWoFFRyhETcJFQN6dxRHY
Ykv/DaQ4EsSgV7j5kTQuo0xCjKiWr/VSghfJ2Yeb0EqeEUem7QPO9SUaiYXStAQy/P+l4QYmJml3
5PR5qImdvnLNkPydFuE4TPAStbMweUC7xLvwfNkEEpEPQkOe4VtC1iv51oI2a/W70JmP1krCi8vv
132g6hCumAJPJiYM6a9SIx+wDi4w0KwIwvg3uzuth2GIwjJEBX2Dt1wVvbez7lIl7Nu9Y0WOXuN0
0RsX7MdMDNkHLNUFDEs8QxxVz5l2u7O8EGsKMW7rDzv/l9FZ/7e6tHSdxjMsb5BeOgZZnA+xB18N
Advm2u+pFB9M7Kv7C/Edxv5j+LdIk8/iH7aMDb9Bm/+tkucRpfJ4pTV1WTGGL5I5ACz/LhzQRwLz
4UMoHnjaRE9IZmC/6lQi2kcC2KK2Kq+SuCbT0M8HIN9rBFl1iOiRvL3wM7eMYtIHfIRO/cTdzw87
wyakJcFPvue2sQQ132v9UefJlu1RtpHTRsPba0Dj5eBXV7wyNveI2wUyuKe5CxAJATXlUSiyn5oM
Q4CahZS/fxyQv2ruwwG6AQeJoXZ1rJkdKipf/Tqq88hkVtZ3x3xUYN7M3GhU+Y4OIjRMUNzz5KWd
GtN4eEns1cI+B5K7FmdAdlupO2M1Fv44r3Hi6POdLDFxNs7DTmSreZaNhqEz2XxsUwky3WJxHV/B
znsvfOenyLEKec4L+PB+F1z5xdUMKHQdHk5QzB48At45T4Ir1OKj+1e56E86OFUV+XGjmQTq7GF7
oQ5gpQODr0/JkTT8IMkj0lDI0RumqGeC8/wjKHL/voE18SIM8tfjHS0+gAsq1pyTRKu4VpvkjRbT
jHXRxX9uHKLK1v2XU67mvgoFoSbblYnx7qI69KvHVhtF45ePsQY5Td7kJotldow3GhdiEwRbm7MW
AfRAmkr62ZNGmi13nVutAc8ZPWmhDwb+puP7uP/F0UHM23sgHfOr+oOwHhYLog/gUZ7pWrrPBCvP
luK1740k0o+kCjQWyQsGo5eDxjqCZ1TH0xrRIeA4qqNJcZ0vEDJD/PcMbredzgMP8YieSietGa2c
bAL2wCdGv+TCXOvQBXigDWUg5JrMLG3sG3e2GDvXdBQJx0tLEnzuU8yhlKaDXp2cAvdfrdk5Gum1
Gfioq1UBqW9I8SBob73lsouKTaJE5Rjq8DhWNI7xkK87Wg0Hd6xMnrGiyH0KJ9+faNOM+hsAD6qT
WrSLO3PxbY8JqScZTPuMxwIke+UAJLV5guRFXRUvYdEOVKv1pnMOioFshmg2ZaMSyj20ElUVn4Vf
pL/Ph6+KXyvFUuFe5sKK8K5cs5JiYkHb/Aij/QLPxu8uTpPqfoDN/QFoqKJ0JHJdVLONtlMBneD1
mOuWcGGGcDa+1MDKabKeXC7VaO+VF9cut7mkrjuyYmjFQgvztEVg4n1oNaCs6MoOikMtr8T6fNJD
Y0JZ+KXy/JMsKIjPRFx8Lb6fp1Fyk8lhfztKxdnX3d4FHhWq/ZKJ3u1cs5WpTKbOS00KtBOVFypr
3ORmlVmN74O3KfAMYkhELb1wgzpMeAfL2CZjBXHVMYQP+1P/49MrluUgYwMhYvW+QPA2w7wUko+k
en5bQokRR4BKsqkNMPPNO9wk+N5UgSubA14UX8mOzmxTHTdB7SosWOhvC4L36YOhCfpCvPeAo85e
lpLDbJP0r/ZbcaMBLDlDFalWhl2sRylrc+2x9/+IdaGii0UxagOelX5puJu21F0N7UAF5fhDpjIy
qDYxsTOKde1w+YjtIjpJkMcjuMKVTjWCFYuHg+mMELmCILx5qeBoXOMONVLjtaUhmpD+6x6Rbg3s
9x3atsXyN7g8/ubKO64VNCDn7LaBSJxdAVhTgi5CT5H4KwMBYjY6AVeqH+UjgJJ0VjktVJHFZNRS
cOSfCe8412ShtUysmoWGLPliU+vTgjo24y0gNeVd/rZw5pGyfMYLraif0bzOD93gMU7URwKZ+jLZ
Cx4z8OfcEf0C9p8BPyK4C0set1d2/CSvKnWnZCP7HJW1TFbo/cgRTCsOw4WtPWSrjWI64wJ0Ays3
1eTeJLf3fAxJSuTMThuSqaiuGBLKckBvraROZPDcOoumH1Qj4IqMhtKfTY3vF/Lj8rO18yvJFYbC
HskAnbuQpb+Z2+OfAiSKt+rx9jwDJZSaQqCV5zUakE5i3+cUDKcO1ZyLIeamg0kOXWyYPM1LM3um
K1GponyIPRhx+HfS1ookv/t/L7afxBR9jhGaZCRCkSDy1JEghwt1+Tsy4tB6dYhrwQM3ZaOdxvja
gvaWDRf2tj8AQRNK2255hfdwBf9WU09xynlVTSWryATY4KMTv0R0YTM0W1/PJuncuaSMiG6jE596
rPvNMNTFMOwHwcWIQgBS/KOfkTQP4d8E0wkyocKQCnrMF0bFE050TjFgPmrDk53eBpDa6yPnt9CZ
dmuv2K9P9Crc1/h82P/0/V6Z6eG15C6IR1Q76tjR3q2ZAHHBUEdq0mI+u1atCR2uFZHSU5QXYAZY
bX6nuY/hzOAzqg82NA3Rx0ux6Wcdo8+SaLmuEg6OJVw9dgN7klqTn8TONu3YGELc4drgX2OkLqOJ
xyDfJyfeV/Ut12ZWkilG+3VZhmWGfRzlHr7a3HQax0e+xvOV9KuGxNbyoVAjShXX1B6nJaEm5rqu
2dMH8NTOegzDJo5PCFGAE30bjvYLNXo6y7WPh38zITEheU+nXNrv9Uo8rM2UOsiWe3lurd8ov1Na
Bj8WDse0Qh77/TrjvhvdG/NsIOqWh2+R4tSYqwNt48fvh7JEeFytBFNT9uDMNCN0w/90MXg07iYd
nCw8gt9jaozJgAy0zWFg1k1ORnh3yVvWEDWyT2KuJoBvqkZMQgCAZITXVa27Vs6pT9T5s9iBiw0U
ytdmKeREKwCgl1WbuuWslChADx3tYYLiKaUE98OzbFLd+JuEs5NcsxkRq5f9oyBG1lUBQ5ze8noq
4aElt+ifeZ4IWFo82ubkb7MhhCMxtLASqYOi0buvRMfiXSH5dljUAmNMjU+zqo54KY7j8hz+tZdk
7IDCRczG2hBzd855aPxU11s4yGCFn1a++hSG/SwK0gpJYaMTbG+uGvvSUkUGcfVXaZRETa112Igb
h0dbaacwoq1BawXNUKnEFNsyqqj/vnFxn1zYVmNu5C0s+WYWYFL8Ob2TeNJ+aKArXiQEOSgdUPRF
NMhtlJ6UDJeQ8MjBWWDLkHPm2eXC7+b+y4Sehd5/COWl4zyzWtLYsA+GvVRu7RlBb+G1aLy+YgWO
l+G2kJ9pDP13cj4kl4qP5JYezLrHSPtQRwEAnpLYV+5rKsvaKdtwVVPEqYvqKRzFitc5yb3G851H
idbM2TR63coBHajsnD0pR/I5so++5bueewqlwdnvA32/hbosYpjZRTFt6K1xVUS3u95XbRO1G2qs
6NHcqGfmsU+tf2p4D6FixBSzU4N5xpDWTQUgWTeeWCnHKkdd5e+S5rrCmYHHiGAC9FBQgLybhzYN
TaF5IKUoTEh7bNJiI3ufHdIwciVv+JEE6vOyOTGyolV15qsUdCWi2tLDUPhZkZQf0HhMHogRe0X7
PQb0q02/wFN44SUd/3He3WMnHcRy+MGwj3/8LSZOyjaKC6IveS1py5urPoNs3wtU40+MkcfQtR8T
bo98acAYcVc0bzs1YQ2Z27b4UZTFQM2YbYcQScKvOzUXSpW56Ovh/aNwnNY+dLRBavFYrZR/xsku
xJbMtDdVueTGV6ZU6M3eieOMNUQDRTrRtSAzJh+bipWRuybJd5kQYjRZAsuVZS1O8M19tYaheYVM
iKOBmXHgsGYWeXJ6PpiayolDUU3KJ1ej1Yej40psbsK0YYaPHg1OfQX/jFljQNgDqP5j+NVCqvyH
ly5UvXor0sqF5fAl3uTxFvwKOgMcgDbWuq2LEsovR/S4BtlC8zySMHIoeoqklrnckhYlhqE+xi++
Ysd+uhoOjEx9+jWxUb2ZBJd4oP/psK94lLu+gbOJRtbEfqkxZmhnBJTBc/DWZAUUqN5KxKAr2oGI
nh7+4cVa/itfPux1eIMk9OVIuYDu5cy78e1BKJN3f/2P5H7ce+FVhw45WyG6p8oJhpIHU+y3hfD+
wmVTDoOi3eDsYEN/PQ25gUyQeaP+naNFHv3zxtZiNlguS7GVFTu4q9Ye1RjdhsZzxWJB1K/qIFj4
sSIFbQOQAXM6AAyiQXXmW+4rX9UoEm58NMAFE0vUi3WflgQmEf8XNFGYPahaWQHGM4UgGlBH2o+A
v+c4mISgesHDRIT2E4AtHD5bEHJnen+aPO67GkfTxIQ7ksymLtP23O705C/dcJ/h27zFJh0TG3PQ
L1tRQ4uG7b6UzZiDHe5jFbrHgxaDFinrq+TzlV2dNpyGDegPagH2gPtPkSNw4yy3sEMgDaehtIDf
8BdqaKxewSfe2ahqQCK/LgJp8jiesMIjuodKp0obE0A/51Nnf2rfgsTo2KRiPjH6WtwPe3MEmoIS
RQEQ0Dr1DkGRTmHT9erfCRCyqSf3Dm+MKRhbnDfwfmJ3Q2T9GupEWtqwO5gtLu7eyIRJbytSRtL9
0XqaSr+eVv/kgcxc/KYdkjn7uV3Muwfa/pgsWPVXrZXpuqalkxDSuzk1g4AGFnMAubdg7Zmiist/
fiZhDMxubK38OEYz6lS8KthAwmPe2vfff83SYRRRxIbCywitBFFqfqw7b98CH+Tmi3fsDkCqQ/3N
hGBlt/pQtl/wOmDWvtoEp2QEHpW1pXBme+iKnjO6hcyxiCIPn56mswwGEKotfT+RGC0HPGNyXosj
4edt5ohNUPsJZeKC1TDDfXt0wqyz/3nTTDdUpGKxlsQe9Zj85DOCO0eWBX1QSDJiIDqql/fhGczf
G8GuQWV7vAS8XOfFnl/BZxNDGY7VldDw7vl+IqbnAO1//YVTs/uj2ge684Ca62c2o/0T8lEWoP1J
KPftpJyl9gvq6698cjUOiO1KlTPbziMGMIBFhp9nyHNy31coUYoXFlp93dfQr+e8fK0BvMic++7c
clAfrl2lp9xJCg/m41FiKAxUPIkgyEPpv42njaCcpHf2/P+TLcurO3Aaawd/FZuaUcUATtPHiw2z
X93p+Lx8nF11RD/ePrRk/7RKp8i7/88fv+kv6HKgVFfVD5044bS++3MXZV2U0WRsZITqc36cTylq
UTNTS+S2xK0gGqEixYcFM+RYMBplQtSPXrHs/81kd4Zm09REgJmhmEVFnpH7d9KecWz09B/3c9gM
jGcwBZQanjHpfwtY68ugfdqarL1ceWXyzBTg2YFJFKSOhgwvKUq/rUIVDBr1IvjFoEGU9kG1G1uI
KFzx50CsKLau6kH8xrp1rYuYzDVAb9rw9VpYwbkzkeyWYcUne6r+dqFmJ0ffpmQse6Q6QokE3Opc
GT90SY76jVQrEoxa4Q7pn0kMmOA7mskPwQNH32X+QO0lq59yZfVus2mvcvJMvr+Fc5GrILSAX9+2
dSkPD3x/3QXYS7GKWKac/sMXsESFq7/0ILcAZ/fUPjWsAZuJWldE3c90KAvQ8rEjpCG+Eh8tZi9Q
blPmBNUsrESE9cjCGmEoWGVq5RSDTIILgIjcn53zaysNzC3z5wdY8QoFUh4kkA5b6MwiHSMvAPY+
NNgKl30jauvemmJnZ9ORRaVZcQFXaDkwU1ljjYlqoXGc7QA7qc276k0il2KvLF6LUIXs42rUZrUY
w9kfJYivksq38Onrxv+77ZoPzrifbyUYV4BGKpEgFEqUlLW1+fFntNpfoMNiWgbiY82PJ2ecLWCv
Z/rMDyuPLTN8vYy9uVImdNBkGTu8YHthOGh6neCJGZ0fwLDnZcGoTYrUOjBOYm2Car7khfCnpqPr
XzF+EGmFTRAWnhT7zBorVVXtjNRq8614qWk4SS249xRYBQfyqEGSb/0V7dzs/ZpRLw/VWxi3ZFxT
YY1gfvmmYgSJsaNRg+3lCgpYJ1rUct+kcyXc8/VD18tmXui39+Gws8XeyqhB7WNuzbAd036oG/R1
BVfkPgCqEFBMXvm46yDXNCVHrHJFg2NIxNUKHY3D/WXCy2wLONpdwGKq2Y3cUdtjlwUie0YCaooQ
BNBRjBTiJZbVZ1KTwU0NR3UOJ5XFPI2wxJdbRpPBWW1D3JkzTCjxAKUGfwAVQqwB5kc9+cPWrhnE
GmLy4ZKDhmy94Wx7Yk1W1Lv+fL0/eXN1MFELcB+UHbgHygf3c7UnI6Lp9F4lBvpdO3Czm25K3FSO
ICKNSWZi9J6jZpomKNFTEq9ScEbXTXRj/NyOtvmjGNCU5ZBG8HaeiDnUvKGLwm44emQ9SJzCPeBF
dV6hywb5y+ky8Y6NlF2Pxi1cdqMsfraTzd2zI8opS0kFGW1ZrTFTWIKB+XYiUi52wQ8E1dvQ+wsR
9e7lS0E8z0h7vDWlEnjwoMqvMS/zGsbKy6jRdAxyYzKtGPDTr/yIGud/KK06fgphM4o7U9Vy2dDj
7FoJZtxtOuWtTaruhlw0vd0WuIcSiOR8bhpNaJ8hpHyGlgCTYbyZ5BCnSFr6LMpGqcAqJJJcsm8U
nrZXGrvS7sATUxUUSynl8PBznW3snI60YMb8V05IJsCqoCdPIKiziYC8bWJ2L7gBCAd9XKlyLIBo
sabbyOV8b2+cwKzbhKykgqvsaRcriLoEIh3VpYjdDiWJq3c3Lx999Wz6sabZdGacatT4J3xtGIMX
g+an3RRO0FNzWaLMdlz/VqEOi3U6C9g5qIXCsg4OIm5MRgSeDvxttZFJz19KkvKfQm3Qkfudqq3g
qMhG+GdGqTLPEYeURkQ5r6KIB6PLlhBa4zafNoo4nf0ujSbOcYM6oKAIoDIpT06bzgNHq8yYVpSd
uqrRizp8vaAXVA3uuzzdavG9P99/1bYKM2Eme7yunYojBtEUruXv0rFjk6bwD6t+aZdhyuvbT50G
N8M9VatH+oYBlWOFuupI8TfCN6lwwzg124VD87/S14vDvdZnlZLUH5Adv9THwh5BbUAOoQN+CHtv
+aEKpmHS4OnN8UB9GLIgRThHSIXa7ejW7vlh5hcfzfR8RnYlNObgML9TPunQY8FUIDA8wKkj/lwD
zZLhkz5UXxeo+S+rJxEDADu46AzKw05WBQGqBwhjnRbzKKoBVe4FOEzQL+ma6ztKVPsmU0tcRQFC
Us/2IL9BaTCvhDSvplUG9/4i0xoQgwcx4scAp3FqyLaJj7dtQIHtdMrE/164be6BTzXgFNA8YaEI
eCCV8T8QaPyvGHVCLYZYUSISxOzLw2/P+EKchKt+CW6hMTQBQykH3ht2tReHZPtIpNQsCA0KEaBa
Z+n40WB41LkLaU6EiVsBZyRqtDJunb3zGO4DsIwFzANvlmyBTyqdNeg4DUlXrDqlehm8ppMF68JQ
BrBeGFcSkmclVZfbpRdWtX+gIKLK2HIfmravjXgUuc/8+hu2LDYhPyShkEDAJ3pHSfmDKD39ez9q
Bv2LJ/7YneeQHC4vOpAQH6znLuDf8bhvHYU2RSTIWm9iRWw7IiALFB9SHqCx8jYNkGLV3xaizR5O
MtBpTX85d6wmYUBXyZ3HVnxRl0ZAWSj6a/EX9zANvnkPzFTGdGtIw5VvhhrMcqH6ajdnqLZwGA9Z
+Yt20eLf7Zt6bDDNm5F3CYFBXL2ulFqAWebCQ0NJqssYB4IIFyLVFU2s6SmimVFxfDQxdlJKHpuw
jaaA7hDbpPRUiYTSoVhqRUxIIDi9pnuHc94rCH0lM7EKiNLIRNxgSd0GFh0/iZM3CAH4L7+q2tE/
YTF6PLYZTo6UPDC9G/fk8mbJ7xTtmIwSEqUik06wmSpTNU5SxqNsKkk9Kq2fw7l0RJdzaM+uw09L
006xlVpJS/U1YHQvhWzaecnf5yItKCwn79D4hrOSygWY1WXpqtHnLYm0TXN3/aZrvhn2PQ/zdeYr
TblBaF9wpt8SaJrKijXK2BPthb3HQVeIqY4VmmJ06J0w1v6tWjvACRxyJ0M76eAWtLTyaaZ5g9jU
Er4tX75l+xSCyFraVkt9++F9xBa8vR+Jvpxkr13I/4fvmJBblxh4ACeJZt6pMyFCKmg3QIZCu43+
UHt/zYs/P/T8Pc/6GND9odGTAkRyLfp55r6X2fUg7tFYXstptrdD1Zzvgh+ScSdGlRZaRboZ5Avl
/IUKkFZjekYyxskzyn80NRtC5Dy4ZUfS1gryVqETUJjtMyBGhq9p3Eu7hbAYMTGA8RJJEUQI1XXG
t4GPYCqEqjxDMzCsbKUCpdhTlB6bp6lO/H2c0HQfF8OxIk+lWAG0iTYwV6eV9CFdKvVRiddMrb74
N2PkpjC0H5YK13NqbU3vevK9K0agSzm2z93b6H8hVm/++8QEs/TEtAcxVh0ftcX3HCCzJi6b8Xau
nx3aUIeR9fYkEnPbe8gOTfc2w2ehL57FqpsLXOctOjCeAmOk6ttpI2tiUTuXEcFW+m3ublaohukw
kPZ2o86/Vz6zpkqGXwGCBghnbc5xCJs4mK+dzXGIvMNH3zH94b+YNYZsVWKfpnnUPT3EtZ5U9y6M
gv5H0irolVrcv2LzReat3TbGIkRl3buqC+xgVGw2jbcvXZ3W9494M646QRJqi+J+GjRZRHiO5Boo
29YtWYWY0+VjpGIOZZU4jyBcjUsWS9IRN5QGS+OwY9BKxTGVH+F2JkNH4Z0s7Yk9gdNYp/DN/ofU
93DJ4af1L8kIuQitvf5GKcSBRPDR2TXzFsqaYjlyBKbegowNHYsXRGup9ED9nUJW3quvMM1rMRN+
rwqfz+Qvrjk7NqVy2dJjtWS6GXAopq4Qt+uT4y9z8W3WgIcWNm/C40bZm6ATe6gR9Dvtc7VLndNW
6FH31P5fGoQB0ymy0XfWTw4EywUbH7l2LFYlqhaQMQ6IoBUz+G9uOXtCFSr47QKW9IU+R5o2i3In
Os4EYII/x3fwx6XQt7Ty6NUwmAr6YJkt3nlVJxGbkLaofOzuwsKlTXelMvKIpJ4qnrlFQMjQLBoB
KY+97dQfDFs4MFPtZymh34hAqOfGKfIchke3FIbBngXkN69y2OUNPJUfLHLRARK0qro0ZCpIJ5wH
t0j6NKXtU7gROFqs1+wWsO8cLZcUy9WteYihF2J0RHLazi06mnRur/kjLCaRf/1RUCM4x9DEtN8l
VBhI5UwnxLnvgCcip8EWynfNdKnTtbkxcPY57nkFBwDe8ApKv9fMdtQf21ooNNUG4k4SSBs2ZIc5
PIMc9hR5NFP7GkzsPCOTieB3tQpcIS3zS6vF8OQLA1mECxw5tnkTpF6wkWjnR+f4++MZLmrhg3Ie
idbrB5QLt2py0h005CEXaI6d8zqYsbaPHWNama/ucdMfmtKsBP6avMXNbU7+7bA1CmC28yRHEeWg
psku9bKNby+0JlgrJs15U5o2vpmd4pARYX1XVGnJMima369sEQw8fSIqXRYlnL+1bmuE40QU+gbF
RiXMawaN6EC0TAnCscaqb/EZcmSG2DnJa8uLtn8t6k6XAMSSgx9SONU9Gs1c9RvjplPPimf/R+RR
JVKRCwQFDogH+u3sFinEcLwnDl5onumzlZYzS7MhBodtGgfV4rCJOl6pIZ2+AdaKNEME2589mBfy
qPK5Ihb1g3r6ZmTx/uU3+dMddsbcPojSU2VBNXJAI+sO3tcm2m2dYRsu4IhYydY8UBhmNhN29moP
SxMDuoYTOzC//1Jh2EOoQ6HJtEe0PlltBuTImr4jk4zvwEbw4Qak/QFwW2y61tAu4M9JtVMfZYuZ
4wk8PIXiAonxJjudjK1vUqxlLBHQs/7dBNhkD0c3tKZxaQUgw5EivqvkSGnxSVV12LsL+kdGs+ER
wqKZAzFmQP1/t2+PExm5Ij1Z+y9HvOa6sK9ADz6fI3qOArqrIyi6uwvg7pCOsloshVOblyKf94EI
BbdDkys042hbhGz4n2Xzg1SM+UeAshHmOIoiDXErXXX4mQmiDbE9GQGSV/UG9HOec74ntDR3ngRN
Dp1yavUW93jdvJKVctGgEYAAyD8L9J3Cca1mSwdCy2gV10Meif6j0V0AGdtuau48z9xBqGAxjrSX
jHkJyv5/Fyb4ChXcPG6UqZMMuU6GEaOHii4PUnOe+jra9cdF7uUC54WCYm0dyBC4Wtf50MnK2rQ+
/sDgxxOK3ZifhC3xcKnoKJUBXhp2ros4ApOkzok/apGCCbIaGZA9GvU70GfkGMF2USrRWYmaXO+X
5DMNi4nAghpu8H08aWPa74EgZHGEv682DQC/8B1b9J3YlazMbrlBGCBXgtmPwdiPCd45BJ/TDMTE
wIKCUEnQxtSDGmjULAPqXs3xo3ucA3+S8s4/9kBo3jJN9nxIzIurvwBMFmoUj0O9C4rS8tpMRUTz
CKcwuOBPE6G+3XndqWZ2OawUgyJ99/+xxQuQUmmX+88xfnRkVLY1KzCdSlnHXixyVPynTwWWe02m
8+dAra00WAn1P8iRYjSqvQx6TAcMasdfXfjnMzP7oa8IicVngQeIDEms3Yt9xaI/qIoJX+SpyDKY
KDyTBGtedMFP1Q96MVqP6lBJOAaUf5PlmiFPGs0bDlMkXnS3SKPGEPMzzb/HoTMzZXCjarpPekcz
vbOrAeNRFeWgkFvyAF/OGQ07qKFU4JyToDWR0oZvD5DJGSzl6rB07udRsVa9BwN6HggnUCWIlZWD
3Ddrkf4kCiaoe/tByHoRnvXPTH8donJIHj3vvk+hWyjhaPSiy5Bk4BxMqkRLxPXpBmpGGKCgHCxG
1akJKwnQg2jc6HhhuUXCS0x+LRqQ1KUzSZFdOh/GNjaIHVQY1Z0bocg2Tcva8709CT+wQmFNG4i3
YcnmJtLvqnq3hvaRx3JkhrpjfwA0KsJz6CtTeOcVH+fuo+xC3SdRTDfAzaYMyhPhIdAgG+XJ7s5r
za/Jja9ey+4xYF0qvcdX5Q4z/KdFJdKxCpP6HgZ4N3QfL8qIh2XTBzRyD7ooP6SQtETUw3f0C5UJ
R2D2dd4WKL7g2fhREBgwENPmEMHefmJl7vfnQSjCHgBMxPpfZq4yHuVjQJ+1/S+t0Gr8B2Zkkbdf
GB5Q4vgbwnwgnK+vkhVNKjcyyJ4WqK69hAj/y4fw1YmVlzOmWfCrJBkrggeBVup0DvoOUqPxJJnu
7V5AfjRc0+kKZejZl6duuzfJbm2Oy8AHIEfwUFhDl4oZkgzYVbLpPLieS28TLz6oy7j1rA3QBHHM
FRAKcTxJp2aiFcWMSzAGgGG4QyBj7+l4lHZUL9bFzj4N61rF5KHP/Z7eGrlWsT9AeCJJDEYXleGN
1TYbQVbD22+aWneT1Cb6UBJOdBYOFyvKmKrqQEgcUQwzsmJEMPDoTFl45jHLnzg3DoZStARBlc6G
++nNmQIBk0EpaZ5WlVrvnI2W7yg8MqF5epBid1vNR7vcuQjcSCcQs3SFitmfJE2KX4szJ2r0g7E5
FtB3DXGAfnlvRWMpP6WzPxRRLEtM85Ew3aJhdE9muhjQ+RQHZOynzN3Ie0JrDjjgHiYFQJ21CETG
QqFn4d+pB3b2GPTM/1vsJCr3+GGBs5grnzbIViM8jx09o/ruhB04Ir96h1PjkPHm1DEgvBj1Q3Rw
6GJPiaAS6TE67IfAmhwEcMkhLDUB9m+M0f2Ya2AfCWKd08h/Rr4oUquoUHPBsvkuP0abCULdAkpk
xyYdhMac7gdMTGKk+d4IiQhrA+DZfEjOPkKO4om3EsD9BrAAFBsA7yS34zPC+FdlrypdZOoYVk6y
arY6Aj6F3oC2P9pjGk+lsUkvCBg7vTexDfIX4yKNcsSWLa6dZDJULMOUB7w/jyI+kFfh4A1rA+AL
jGNlEBicSRBfJMjoxo1Xn67RS2OxiU5uUpIvi0bgCHJcNu6IfRoS41wg22GoYtNkWiBaR9aZopmI
Eim9CHaZTigZlxkFB0wQXmCHU0Mt6aJ3Sy4W5ytgdV7C0H7Td6chvP4voJAlM6OGUPneVlZy1omx
3Mh0W+XfUiv9d0avTYjc61O/cSIhk4UOTe6aWupH1QpLHYOSKXBK3eDH0yEFySuL1kH9hAOSiZzU
yXcnW8f78jpX3K4/Mo6Kq5P0lkif5uaCbwg3kgrlyQ+jmZI8qLaiVN4SRNo7oX+DIBeqdnRjv67v
Xs2MjY+Py43Fmq6azAqWRblgqkgjj/fPmDo3pJhHHCR8A+C71/9ToU8FA6RU6ojj3o1bseMhTDTG
/Iii2+5jc+dWiYvFzwQsJSLDJD9bYyYVqoxcYjpzJm5a38we8z4sqL7k2AITqhMle7ynBipZ8Vvy
uejGU7Qew6LNFeyPjhJt+8jB61PjLmq5Ghc8xHsMZLeHi8P7vTPphpbEWZeTddi3DCdnK4QBbNYH
TNuU+ZrmH1L162Ym1ilMmMp24mADBHERrriKlKvtGlE0KG2v0EOukAtxIQ/b3/KO2t2taMst19Hq
ZOJ8rKP0P0x6Q7iUdiOAcVH0/qmIEmVZMFz42lO1sOi4MxvmYH2sgN6D7BZK5Z7shTv0cymCtoHz
zCOMjYE/EXfsuZMSOS/363hg/p9RRsY9WFxnH4ErK7AHLbqYLdpak71UC1K+EMGBJffNYDRY7r+5
BDe++jiw4rEiog6os6nQc3begAeofez4Kblwu2JiaztG4ZGYb4xMjcAhLJx7x+ye2+/EIIx0LVbL
OAzwrIMKT8Tvti02jNQxc55ZCy/LOhVRqnxI+zTwT6IFjS9UICFC+m3tIV31GQfIijA/uH4JlKtt
sxHZKimWmrhvMtBro0cb/9vZofxSiC+gkUSe7JuzScmTbvVh7TXAsZrXYtvx3udaDreVpAY9/u/n
6ZQg594dCiaiWSgZDJAkwy8L3zz4jQWTTJufHEu5DQtnPcF43yR5c+ZEpKGXOjVxn1cm3xOVXWnq
LZ0MkbMBAGxTTjmZ7duN44xgcrpmNowHpCBOLHHih+eIGoxWwGv0weF89aRrs24tYJbSekNqX5Sk
R9cWMvMtQCA2Sv9zV3Wqha0SdS8ZRaLNmiM6wh2auOZOnEE66a+AFYdXyaymc1McggaIZmKU9zfn
8OC+cbfhUkMxiPAUnNEjR42XkabTYrS0J0Oz0U9oyU2I74Oc/zYg54kicDz7nUBWkikhQsiBgJ1i
HKi+0rnp/bnnwU1P9UiSJnHX0nwF9rDmBy/PKiRVu8oYpWsc8aruCZDwtX8XzqzI6unX77d7NxTq
05HrshDYs17lCl8nstzAlgMzwwTiuvwTYZrATMeoZpalQB6rCvD967NwmZtdbYXUFH0TcpOz/6Tt
wpqd5f7fDMtuLzjdvHb/fgMQ6wT8Gi+35gzfIw8EI+HojEs3L0CurMemGnKhehOyn/v3Nldfm1h9
XJFpQ2HRmS5vc24y8RazR6z66Yd99EXs3Lx/TG8KyN56Zm1AQRjwS9IkiKWCPAzBk8K6rLcEOkV9
2u7A2gB3BoDH1PDByQmUzB5HnqpgTiGVIAdR1huROwKy8uN3A7s9dhb9hk07IuYqgFQHd7zOUfd4
zzFLzX1DMTQ0/bFlthFKYoMiYFhX3TUNWIBW9TQ1UM51y5qTpLoFaO6W1TOe1894KE5b6pJlcg5G
HL2eAfd+cqzyMQHwqaZI30OEjxFx3YI33lR7BMv/HWLhag87gdnsHrtKfUt/O+oX/KqvZgpk3b3z
srXozujb8af7Qxo76gCqk9utE/aPu/BWn1mb/hrgBlLZ1SLRAjRm5jNks3RAfvRfUNmjKnBGgiw+
YvPTbuUZO4wKVsLYRH4QMqzow+9+5V8i3xgcNz5wR0ulP6tRRL2NQzOx6QcmNMicpPSBPPyRRl1n
8wcULuDAKtePSCqnQ9tRuWtviQCfI+m+3G7QfQucpJehZsvRcd8HwwObFfBg3zqVaFZTgIA2RV1D
B53x3FneqRhOlXFfQZcSgSwZ70BJd8g75HgC7eHYg0aJT5NJdMUqiS2gIVsz2BMa3sZdChPrMxfI
uazCRxfz8JZQi4XjasAJPpyGLFUgj4VrB+DVGq4bXYYYsIUl2HuaFJyeTNkmI87x1NbIn49lPw73
/zbZqjxIUd46S6P6eCZ1Oet8vQqLzNpKLSKPCPBEQ1TSx2caw+3yzfr5qzpoOIAXv4gFjDYNzagj
93zYiGFXkF/wom48q166j50RXLbQD334hYT6Us8I6FPjHRSiWdWphVeJoaBiDuEWSj3IkIdtGf1J
YlCh0x7eTF1urQgnWWXWKBk34tGYZaa0081sJ3FKgax/Az14qJ0bGwmzNLiwxfMCRLF1aEcWuLOb
b2RI359GcFADS19oD5UIlSdTTEBvTJxf9r7ekVtWcQ3pNBiuC+PU8q5v3MszkZtpKdNYVG8snfnF
h2gYJPsbHIs9LMFAAiouEgDrNf6ZjqKttqEZIANzEcijLAijqsooL7DWg56jn8wNMFfK7+6nGjbQ
kvdixgVv3c59o40nUPcYCM56B3wg8CDLXdo7D7Y9UQGm2WNQX037JcCc1sTG+I4dfIV7B/PMikId
3A5BlsDSNqzNEnleD/jm8v9I20IMaAyakTSG7z08DI6ySUobxUT4u8DHf4g43o5q+ZdvhNurgrJH
MKtBvRlHOVGqcOfljFqTBWSc60mp5Y2xAkiApqugu5AA0feaPssj1u/H4JkBT2Fh3yBPfyhZqqt2
jujNJO8bwTZM3Tzd31irtEkckkIUtBGopVv+wXuTTCahp9CKaZEhjCAvi6MdGO80upSqfY1nXCSF
naMenvoid9qSK4t53GRjbkks6eQiL3Ke8k4BY3umNy/lj1OAS6j0QmxU5VyL8uReKLhkbDxpzTIT
UkjLziV6KS6ixSgwG1AcvYv6klTZxFk/Pf3QkitjXJDzdLkdCjct8wevaKZupRYvIHb/AmsiBDWi
/U+QQyF0GAod4C+ddwIs38e3ChMt8xL617m9F15usdiAqnJDtTvKjgR+JXNooOmdbZoXDJxQgB7c
1ZURO1GfAwU3eL/tRg7EExwhi084fmmLBVJ2AlM0cViT3QimsW/OsbV05XC7U5gORt/yKlJJlkRO
8IhdJDvYeRRfwmnq5fylZg0RbciXvHy0sduBKs3c3YCZOBEYAwXmJobm8n6eJ6Hl9/whsJ3C/Omo
SvaO/3af/L/QKtVMGJAzC52iTLnj7UgNRxu8Otf9xUFAYhnL+13Cly/vPkUMckvW1/ezhHr9CnTE
JBMPtnZmJa2Qe0ju0NYAXWQVh5aceXtrBqvlzHwh26TnaRRe+pI/c0qt13zdwNXbitP+DYvtAfIC
zS3LyVwTHp6AcEJWUVplgVIZAtPe7Xh3OwGG59rIFVQn274GC2Jdjh42Qum8D1lwOh4ckRI2CUXP
p3hr93OeKBN43/eFAXOGTYsNCy+QAyauq6yYDs8NNkrAnYqFY98u8IvlQFuODJxtzvDCfQAF4KaQ
cUVmaviyEi1qqzj5UaDxwWmb/j0gZJWYQ1BhrQyjbybo75n5BSNP1gAHKHKj3ntLGmkrRUdcEyRp
MJC9zqna1jXyrQRUKSF9b/d4ZN4qWyfTSLvuo0g9gLJP7j7gbt6JjMD/H5rprIn4k8GevmJYq8ri
4rFiBjCRAvdnM9davHXDb/BqL7jjhz+X7VewP5U7VdKEWWLKTgZQWJ7gtYF6JnTA9nHRP7ZCLP+t
109lbvrABgJ+WnPbu1KGENP9owMV6Hvsh2/SlAYIm9zbC40M9mIZ5IxczHAgCEa3f27q4yk7ahMm
l2wu4PwMrcJ6hXo1O+SgLs2yE2gRO6U/vbSS9NudOBcUHSA2X0l1bAcmXrM2rqKxK0ucx4xiQlDm
K/tA5ZMQ2tzVIKcUDQ204zA2bd4wzdEgD4f8m1yOcL52X7OGKlUAydu/Q6hose968CSkkhez8I78
PaVb6GxrehhZTXHZXohKM6JajON8AKBihQkRiEFePzDPrKAahm/p8IF7u6H9rOTzGvZzbAp9o0M8
83c4EZaC5+GakxHubf/rhz7KGTU6v8hT9x50SUIX1SS7AmORd//WR34qMc7r1mw3z4wA9Dwirf9S
237MYWrvzlxxSLyNEYdcchC6/Kg/k9ba6zi4zWVTDYONtpg0E43aeSiXkXad0lIr5Icrd1/sKpzN
vUuqfRLWJjL7WN2xSbw6nbOWu5o6U/85FRkzAqkTpz82s68P5jhSOjasA5RCYD7DEvPqxf13qgDz
BTPsRXYZ3lNRVaoFDqK0BU93JkcHDLo84SpDLEYKR/CadAdOuCBnxieJaPVQktj4yG9q0OIM9mV4
fmHzAD9PMZpwegxd8u9M4dkyYVqQzuwNiifkjcIl1WGe1fVd4mkZGodlnrS1m9K5ST6SuLw1IU8v
0dnlwhG7hHc/FRMCkR/IVgfeyZgTO+lqHa73lfubj26osDoa31djDvyIahBTH4XuIjrjEnilxJse
Es+35LQEQOktP1PAH32dg+ViPCIdWs9tvEjZ265OJDAOufGwBfYrulwvKgAPbOy5k1lEBTYU1GZm
Q9N6toRPITcQClwB6MhS7sewsQjHS5tqw7gT1Ub10fxsZ8YhExDKBKrJeNZAs0MmVKvIupTRyb0v
OmpZOSFZ8jJJf3l2r8j87OwyYdGbnfUIJ5yJcVdfoR4Rr+wM9AItYZeXq3eqx/XeRLQ+MguMBYfi
sWeVIEk3wmsnLetEHxaOdtNDjT76CfS2MqbB/mAQIYLNWEN/h2IFRPE0Eby+6+75cuvGMDegpmvK
qRKwcPr0rc1sO7dHjfYGW6iMjRDGFhi/IfIml16YpemiJ8bfLaUQvVJZmK67+UAZvmFcByVXMxUs
k0ms956/Ki8ZZq1TzkYYDTBlAl/9SZOqI4VETRcWGkRos0ZhUznEVFJoPS/Z9I+v1BzyEgfcbGtU
dlVZJ5lyMFnciKZBO6VanG1vk5tSyUErvcvjp4foWM5oqgepXxYOYCjgIkk/QjKF1SPODprz+W5z
2d+BgNDls6JbFYJEU+AYYerVSCgyWIiTvdvAzX09gYiY8Uk5cZmSGAD5MgxFp7gajOufzunCXN4h
LLdmH6zJ3BP4h97uvfDre2vKpOp/j9F7BZA13PrfMUtt62MY9iK+bnzAdksC2Py21zvi5dqBweWG
brXlHQ0MCUSEORM8hhALCmbFCDeLg9G/hjiYyNeGJ1zxs76eeVSfHP+pd0G5FnVEakMhn+tdNnbk
fq5CVZUIDY6cMtkpTAgYU4SqOTA4HX82CXRjhsSsH23bR9yZRG9xtPUHIp3nJmKNxCidB1np0JV+
Cc9srMshJ/1imdi0babiN457X3SH6NrxAjLgqLMJBTfcJ/UfnQ8KSUs2R4YtDqYbAfnJZERpWNzr
JcaN0WMa2/UB3Aa1F3Zp+azWxMZgWi1PaJWyL9D9rug+cG6lTd9BH7M2zHjut+1AD+ORrx39XopZ
LyL2aYMXOQ1V5mnTPSfrIPMOvECL0Rlu17Pi/xA1rIXSqGK40GCwX+U134XM63007apa0d1mFa43
WcIN/GG0058T+m5J33m1ujcERkVfRhnpc/82QTLOYZV8B36yJTNSlxhopgfNMUmZsJRMoWnvF8rF
QpytFYCdzYNXXmb6aRpNodtM9Wxids62cZEmnHaIBxA0wKQyQu8vXB9/X+2aNYWynWDCrIgeSZ+w
bh2Kf2w7c1PIeQrtx05HkCE2oqtzn+QwBUtpoZyCvSwGz8BLRQpDr9KKjGPZ9wHiZvplKQ4OSzpo
n01Vlmk+2Zc4l8+8xVsvZMexT8jUm4Mu80aVtuyW6/9RJvBoytAJPp/q3Wcn0JjTgWWC0h6zRP2b
hzXj5jS+sTfx2fdVL1WXDeaiqsKS21v3lu585owsxamnZcLutt3KETg88M0/+1zF4juvHO4YIN23
aFDtnweuwMHgqRTvvXdhCm5q0L9KTRAk7sV6CMNA594XdfuPDO0tWWoPNj7kZJjOIHDxgSfWCcx5
1FP07FdGNiba1NkcQ9+Bengzp+PTrfPzGvbwdrpuT480U0Guc4vktib/wPR4GUEScGWCR8coREfZ
NpYtfvVLYfNJxxfhsaM5P6qgf9B+1jUL/ia070DOQIl1gnS9CcO1T8xjYoxifsLz8agsEMrzLMTy
81na+TeP4Ju7TFzWpqsbSTh4bYjROJIqCOeU0+9nkpvQDFUNBwWq5EPc8gTZrGe8NAPSM51p/s2S
UkQAkmtFGkuVo5V3JTVrJjVNL12tRTepR9pz7+kJF9xR8BwyjHdAuYHpLCR6wRFtFNG8g+1KzYxO
LLQP95khuyV/WKSAGASZToK8v3YnanLuraPsqiqB8rTYCXmzFNiqNQjGmc7GmMH8CdhaFUAU8vXZ
ftNsjp1yWDSZkbraU8+jIbHbzS0p5zkiCjxWVS3xRCwsy96FULxRgEa93SxGJJCO/Yc8BB0hImje
zYqhwBV+i6zcGP5nF5FciGz76EW9RE9WwJhSFAslUKEJLsv3NtGBD4x7imSnn0kyZHJsv2Rxy94G
M8k50umrFWIowHxIrrVvELYSVy8awAHVzbxZ2IYQx8IGgEzQUngdDqSkxPoVdZyZOUrULlJas4t7
Zu7q4DNJTSRrSWWEYsqrRNM0UvPKYAfdm04Gzs2bN3sxzKlG8kyOSoRrwQFCVtnQM+2U9vS9YOgr
J46V41U1YZIC2vEPPW+RXPQU73kSc32dIqjZcjjiudjSISp4mGIGDQR4EtyC2UBdGekzSHQwO3+G
Vf4K02ikoikV8pEfhLksJ0lw1pMMKnTugXM9iMRtFmK9SaNKY311kYs5OvMe/HohjqNoOutTo0JP
JQ+ODsg2Km5fCUfE4hFHNru5fvyxtNf8/fG8FcAQJku+ELOseq1OQhHI5t0l3lYgov3Ei8iuSxXo
wB+XYsn0G8OSzFHqnxns/Lb3uzZ4WSJ+6IUGl4YFltofXr6WcqzQMFgtfvXL+Vechp7jL5ZyOK6b
DSdi3+EYiWu6YeFV6tHjAxRsFR3kDNJhNEPyqC+YWZ9Lz8UqXpFvPbhqx4eIobl2qzV1KQzuWf6a
SBm8YBt+DGP1ae/VaKhNpugit0V36ZioGmX7S9DJpJhI/fkwtqoMUvii2HTGOFxAK7mZqiv0UV4X
8S3WYKQSQ2FcAB7Bm9PTlO5P+311Kb/mPFQVEmrPljLx9rXqafFmW1GTmkLSiLz+X0yPPWijBXut
wFmgkQpOjAPM1ZP7mv9/8uoLk20F2460bavX5UwOFbyW+IVCMfmELpPlDCfpEnqf0UHHDWuNMbND
PAMU0E3pkTowPQW5XQ/xTts5lgt6Sy4rWcpqClUkSNwlNIl3DqLc3AV07pArR/K3dcUUjEAUUoYm
CHO50+fr6TqTURoulUTAvMhsHdaV6iSo48h0TJoc0hCUm8LklH2LXdtdt8Oh9ATWY2mzRpUoxBz/
o84P9bwBhNDHPZqr62MKNFjSSN6jSPMHhhxYXG9hbPFhNsAGPgJ7bNDGzAdtvD2YdcjQgRVjoRPt
CfYl+dAkyd6q6NadQV1F2n0B+wSLJBiy1kXtTQSd6dtC/l+reIrybZWqxI6ATZJOmXehKEGzbmiR
eWnkQsD7UDcJP/8N+BV9n4x/oE0GZpUwYD4YTdOCRnbNGh3POO3JBNLdAm1P6/ZDZ3kLJWW1xNrq
zDIKXogaYq05blkbgR0MXoacdWVNAIKjcbka7dqh6/3FtKI/bdRHzebGkQbbhM1KzqbrbG09GuMq
GmN4f31NNfbc/W9s9z28RqfCMTm6ow3pV3nT4JdPmbc6BH0Iw7CiEQC03dZ9hsMYFAn24OvcgGs3
db/5ecoJe9gOjtxvQEbiEyfvIzlHWPrf09xdRq+jT/4l6BzZAT8w7nqibekERWlDmI97Dm7AH23j
C7mzINDsdEt/5FKDnx/mYWkoc+hNO7b2FfDPwyFy34/4Mq37GKLAYh1r/LVE5/FEy10IH5s09bnx
QbRV+18Bbwq6EnKaUI/WeUOJ1tpbXzD6NlNUZLyNblSP7QLvmQlo6SsJo3JCfulUOq3AoY/ASDi4
BBX+/FwD42ZAZueK/9lTEDA77Enz3hf4VmqYMc0/mQ2S86g7DQR8yqm/NOfZD+agzFFsFGpdxB6q
EVdHskdVqFacPVUEvQvJdVSs3r3E3CFh2YLfEtEdzUkEIJcxKzwslNuOailrpVG4Of7VzlAiSVcH
Z/kUSqp8afKhnKqgAC32fs/vayIkgfDLPCyxiWsBxLrCPrcGGcoasS3dLsNFLs5p56aV9m8v96wm
LptENAyCIRToa57qD9RIeEZu/DEwo8TLqQGzfZGua4SWopHYXF199sHHrEiktC7QjYwDw9lxdsjq
yziY9yZYtIZFYooXd9UdtySSWC1ma3yrapgeDDUTvJ7l+rN52jYpvjc3cA0tuBloHJonk8c2yAWA
PuKjf//G930QYeu3zIXICrQQ9VXmJ+LiOMJMLjPlXefyZW6iRfy/VBJ5mtPRsEzqufd2OLgqFO2X
L7JIU/g6zNU9r0EB8KaB+COwb67vmiaf1rCzSGENsOk+RCpvL/p87bGzTau18rP10uLm7JWTfEax
1Q6pSW0nBPcsLmx2s0wtCmf3tw5+vfgfC7RlPQTgeJGZrRSVT7OKwGqZfa7M8k8I8YwZYpgY1648
N6xVP4cqR9rjtBGcgW16BiksWQ9lsGUp65azsCr1/XyeXjHFoBJ7zkI1Hu7Vw5MgxoloshoCczcE
PNv3LbrGg/XfSTCVDZJ+xc91F/L4ypvoJsyATMUy9PE2xqGMYAPMYzLOki5PX6Qa5QjIUvUVt/J8
yhTDEqDF4cTJfYrkCaaTou56zji9Rh2z5oI1QR0Rg3vP6SM6Ly3nMQDDeA79u6xgSxWavQFO1jtG
Uv55LaUN0yK6yz5xPsF5dCcERl1COgytsbC2iu2KiMggt6UXUuGN6KJciuFUSRfhKwV01gYd+awd
pS1JUooDmM1aF0V5kGUFLL0Gn5p5GAF7d+kujy78hd9D+sS/TYhfVsVwGUn4nGaJQtCdxekP7nzh
IIznDehGIpd6L0cU+IrSy7Cgo4DsiYFR+Y1tDJiRtEyr+kVYSnxQa9FodyAdoE+ETPsCwSQc0T+X
U0hrvOqC55Re5hkVQ6u7bBxhVaK3QGEUvpgM7mQFTPZOSX3fAJ4c+nU9xVH1ndIDEKtB6cp57SbT
kxEK18SeAYOBwcTWF8SNDx5FB3yRzrF+Ft9/sdmW/J6m++eLrmU3OoB7yq5pQ+AuEUerme2fWRNt
i3A76x9mEN76LrUWJ0AMT/MxvJqkTlkw1JnCTP7JeLY55wXmNkTeJ1BKa5G2eJl7FtWVrk5rbHnR
zlkzFPDCp7bRY9z01QAU6/V4cAjVhgVa3dTy1h91LIR0kYVhDndjWo2KdWqMgizvcFoDBo4puMA0
kR0h7kbElCplsl4xluYnkrMhoImxjqGbIxqtzS2+Y34LfO/4rx3azNtqKRA6xJpgAUz6/lG7KWnN
Quwld9UxtQSqKshDxR+hl3OJgLPSWraYWPHr30u2Vm1zzrIgujwKBnYMkVREbjcgy8+YTHACfhsP
ecLAMMtfVKPVv5Ui8l+dCSKJHIY3i6LlQ7RlmI0UcL73WCnbk3d0MC36MBUqLUfTiHrD1ogZ8TK0
KHEERcSfcBmdmQKRA3GfhYEPn1qe4QyfDiVMH2VbcP/7+bQ5rwdclyAajqoIvXOpeppNxl4xykBs
IMb5eZHCW9+7KNBT7enswsu6M0DAsAsUk7nL0M6ifp6iwKQKyv/0YvoyXshKKLWs6HQd5E8eau4H
vA/FuujP2Fg9IIKmpCsBSsuPujN+R3iXGhAmcDF/kg52QiaO+y5Dd2DCoUup3nv4eEhRJZwcKRS6
RRRf3YiVz9+YlkYBU1A4UzSwpsB9ryMF2g4WrMAplOhkgOzVChcjs4vEIZWOKro/5R1K9ee3GiLy
OOXENLuU+8DciIr1Cgww39y1/0gzx8kjLjG23GEg5z4mtEd8oxrLhUWkeEGPbBafO0FSW8h/kbFZ
LhlJ1Vx72VSpQKcUKS6ST4Jj4i/Nd3/tmVIcm3jFwBkchMPctV2Daixl43eZis9Y41bpUgCDRrEQ
b2wEA/2Ge3R11C1k6yU04Lc2o502s52xUn/rEsPRMDOimbZItVnWo4PWqUpGmHAlFS7/rOACZ2W2
tF+n6FfYBAs53fMuQjC9VwWGHBe2hF5l/lKDaYLHvrnkS/8RpgaLwcZl15vvh5yf/X7l79dFUwjm
RTAXiA6GIYmLyPdeaNYeEZXXHK3V2jeTkhmJf56NtZq3me6o1Q2Fgm6Urd+3WPyvFReM+eeNPSmx
Aej6n/yyQaGwj8ECXf9zuh0MvyCIQn7fd9L0CVhGTBJsbxF4hluJY/WlZvwwadrodsna/pMUaue+
4u4GU3FFCgGJ6aCJ/Yo+rgf+OeGkWCBuUGYqnoPg4U+7fWAC/OZzyy3/cGffuH0QdLYaBzO8776M
DZizSHQ319tHqioimwM50RyzJ2v7vVhYtxy/MX1TdQ3iu4a21P+7Ho/31ux8nATz/Jzc1tAH4XCh
yKe3Zs24+tmGiGq3O+qVzlUXquvt6A1iEpdQKFS1fBoM6KvQ5eSPuJxTNCcJNJ3eFsSoX5QJaXJD
7gCnoaqer37ISceXFjsR4sAXXotdKJ75X7pw+2UUYR5l4R1YaQ74wrCyEvet90ZiPJyQCE1vaFpz
KoekrlU6UoIFv0uhEt1A/+5kLkOUlbRNMHwMCUptgOgMhkeAZCeq5D5j+nzylnlWgT5CucG/R9Qn
9/OfT1vOs8I2toDgDQq4h5M+6n1jg5rq5qT6ht5ipLDwqXoPnjmHvLvrz0FLLa+5F2KiL/7Zrlzm
4SVFonPbkwkWBcXGkrADMKBzb3jDaTVg3SKmL02+tH7SUBaKtzYtdjZROwtHAKibBTd5ilQtpOxY
gqbdVny0aInw46TfRVpvJnX3FCtbj3KMa4z4R0ixzyJJJ67K7GultiVTShUp3aYvwVMIXyQNUYsf
xF+DbFtE7rYj+vrtkeuCG8TlTtV1q9M6yhCkk0zRXMQ0AgtSZDeGYDOBHxAYyBx8/sanWd/MpcvN
k/6RIFXJAMHA6UmIiPptu0nKDEVd80K1m0EnBuU8reQGQMmARpiQQdscjkShCKF2M+dVNIAl7pcb
CEDDxo1uKTCIN8JOXlRTzNlXT/z881Hizf1lvgzABG5yYxJjQZ29aFdtPUdXjuiFcJMy/6vGXb9y
zYxuYWCscElRKGELxVU2sneRd21vHjpyfCQ0QFK2nhx2eBWVmUlgQFqtrlAaDOrnFSje8Vpa/S/m
iV8iZGgAAlyczCK74hUQfl7QNxg/unKU4qtfp//bY1WM0KWU+pfG4wdZY6wHpzqUdAsSkOYFvjGI
/R2SHTHiaMBfEtaSpy5GWXXwjBs+iplGalx7CLuAP3PR1SuN9aCn4ndZ6CXiODJLiZ+yWVZUe+j4
q3Ke/NwxAsy5X0nW1yIgEjzdHF9NqauofnaZlI3qIZyRyzAboM6zHjC1xOsUxPQHduXarCtEA6+Q
DaBaQ8eDSNYJySmEne7+Ve3VKZBhj6h/FhDGO5kYq+6TMpMG/aZQcNDbDtVtYEao4xDn9EVN7Pj3
6vLF5kClV8dANbsvJNQfLBJSaGqJBvx8DEkqIONHAbWtuV/Jl5CSpp/a6K77wDdYf2/LodJoJlNz
WJmU2uiBX3k0uF1PfWB3eWIYCDcLulTlAiGlI3YzJ4llrlK4dNWCLoOs1gSmXzTkIiMtqPxuXU8H
ArNASV9xu34+neUw53NLcwQtTGDJPuB8IJhXOJPL6G/gxwVFy8RKCttwRps3Ci6NKi178gy528eM
rpakjxJ1Y0w1TsV4/U1iPrLuoX1UqybGIrE9gJR87lTBMRLxp741Wf5kfHG0eT09/bpHF74249MH
OHwmJIHV3RkUFMN0GG9MAIIqXilH5wEt9BPTdbwb7QqnBIJJv3VewntXedPE0ukfAWH9d2lGF5e7
2V4pbeWB4m/T55BeYzepoA/iLcHWPHXNdy2BPnJWyy31wXEEB2dMiZaocG36MeqqQ02JLK1IAuu9
ACW9rW9sXsAh5WvttkTVtM2W3n0bL7jU3lh0mSUTxDHFcjdiyHJSF2ODZnABUJh4OTWHhCKMykMA
jJSWWKiWm0idUaDSNXb8amaO7zsETHvvwygkfOHLbIRDDw3tGN69XwHtmZrtkzSCYEbwfDhSIOPH
36DxjI0sxaGp484lgucreym0bzk+BhWOcQTFbF+AGiYvbXtzJxbyPpvV7L4ItvsTbjpAOeCu/EqT
V91SlBlK5cKOQnKH6lvKps0QHyuRn0fjQsDkpYf3N6hA3WsZx8j2kKrZzqjNs23tknY18gjntoQ2
DgGqRI9/yrIQqE+m4rvIiYorPxSX1Sa911tFAUOujU7Ub2WeUrlWPyzGAoGt3vsP+HZUana4glVV
wvv2c4O55SDVR47+3efZhq6Xehd+mIVhW8FKLdlUMe9iVX2o55H/nV0fxZZr2dVIMjRbR9LCcgoQ
RtR5entTgMQydh0TK+A7d1ItAEoz8vsd+5Nx8/+Fjo3YB+kOXqOGo8olvi32a66SJ4zH48D3hwQQ
x6Z4SZ0fLFAGVkxjzBytLR5T3HEDsG6n335sd6NMJQuO5Q0He3TVy+eEGlwZwwD0J20VuSflLCsL
mEbCAPs0yWH/cATvans9NKUdVcaVa3wOZEg8cOuqL3EONLMIvfKM7PypsumluIQT6Fan1DqoJG9j
xqms7wud33AWqHPlV1v2gmlyCYDWWPraLahYcdt6IEfU8jnJYYBUB09CfDEkoRigvlCDrpR9cKui
jmxtNORKzouXPnUvn6L9RDdMoGu47T8CGZRwgAtxNiQgQS2V3aWjiugFBsYp1vhXqFfbIL6gWdCw
xSkbCNrMT8UebMB8qDgNAV+wt7OIkRS7P688gHjpewR0uQFXNb+jpFIdhV+qywYpqmdm4tLqvy8r
xrGv898r+KrJ/sgkydOrYyE9wFk5ebvGVJmzEVKb2BmyvLNpZLug0hXD8NA8sym/Saiw5IwxyQCr
s52Qr8M6KFMa1Y+aGal/25+xY8SWeEqhpKchhEl8MfCWuixieru3crIgl8OHoZ9Na4uOUXbfWMsD
LXFTZ1+G6Dmi6eUFGOvG/aPrboYxMWb6Kvi881G38dty+XQx6eTpYmpNzPsCH/x59Pu7iVGox/bc
wC4Uh1g5QD87IC/uNug+clw5p/lprQQzR2IweakoQ8ad42LvtkITWUkfA7rwQCeP1TgtYwAPuH3A
9FJLvVhA7edFAJnRqnFBoBPqk/Wa2Z3pD5FBpPzQ5SUOpnzeZcz2DNOpYzHO9K1OH/bszemmj7cP
dj+xZJLnzdGoP9BpJ4z1Ov9/c0x2xkmc/XfXUgJ4dF/RFZWyqD1hxBUN6y1Q1gqkxXMNoSwgum6L
YjDD+7GZsSeU15D6JWyTTv3ccPnawHsD+x7xiJT3QTv7NjvOC1qQMcQ1KDbW3Cqs6ZY71QbUKqyD
2na9Ilu0tbnrE8OshaUOe0Bebe3T/Bq9fZMjzbGMM3GkShPRm8jYU2pDv733PQ3A3lNRkM8EuWQz
pYFgK3udXRL+VWCNPdw7UCogg4SoE6xq9BTeCTWNFBARlNmLcoli7Wb/uKwUBOMR/C7Ehzaffa7Z
2pPropD7pHUoeMxV9kE77IkMKjUCrUDHjn5G9aCRaIcxhqtJ64ENViGvg80uTNMHWtp9TlsQlHF3
wxj45PFuIEVVwdhxOCvpk+JcNHM0SYvo933XeRQPW/uuhcIOJ5tMTom1R3iYIauc36vACbB47Alx
ZUk4ldJfn3DFwpbmOdNpCFutplOjCSHndH31HlSlfSDj6wS+Kzx5K9/Hu/4M38Vm+qtvjv6E2F6W
RzXBao09IA3/2tZNMdpjYxzzlqP+YxIqml1GNcHLqtuTEu5mGnGTSwnARfQvtCDo6BRG0bivpyHN
yxxbgsN0+/d8QcfO7dmsdjlACBXdjb2tm3yOyIol/k5YiUdvnumIzoZeXvqP7DHN9brtnXsLSVrP
/UJx/HTCIPkIcpf+Jo/Ph4SsbF8ZLdNwDhvcNvo4uRv92ZPzUnM/G96F3EoJWzTWSsjTv/D97p7c
tXulefSLygxUQ5tAJYynmlR4+NN1TgjvtjfM09VVyg64NZUKg92qepShWzW+1jPDykfsBeg41Etd
U2psZtkMe+SQC1fRmLimOlQTrEW4HUa+DLTIJs18YIY2dZn0WhP50NmeIapYZCEBzRNhjt2iB0VE
5pJ1fp/4Ma/0fOvdcKc9a3iVXuKyp/zInSj3qo8rAKtQjoIWePYNggxtukSirliW1ktVLrf1Tkip
7HpuPRwIhJQ7onUokAcQ9eaOy/+3tAYpByjsLg9qKy2DRDgEbGumTNxfIhv5PMnmrVlCBW4BvIB0
6wa4dqyb2YxLRauyxAVe+C0ncSamwdAqfkPon1dlbxUQcqUkHI2JJZ9q236CqOh3PQgXsItAWhvU
byx7Rs4fs7JXD8IoXM4ESY1EISseutrPQ4aJkY8NxiME6ZvGpKov+7D+L2W+jpdCNcPTibUMAkit
L7BVXEtX/gMxuOkjmQx0JxLE2ec6diCYXr+sBOYE3RtYTwZAo8E//SPWEfDQLKSvQNRybvkAulJY
K3iYfXE65rGkg63IzKYBg3Q2N8Ny4fTa5Mx94BMDj5ml7aPeQyoj5ZNba8FdYFIOoAJYFmNO4ARv
4niXS6KGqLi3T2JHYlEeRGvBx6Nw9X2bR3OPJI6cgHLjsfYg8n6YKwfwSHd2SmeIbHOS1LH1EYd6
jaGxt17cPlF4PNHvy07QdOAMfuyfoMBhc5I2FB2Dd6xSO0/xel8TlxLPXYwmKHUvn3kzNoIjlyYF
cnj+yxmBSze1KSQu6MZoP6fkmS2NeDmOUT4JRvTO+gSBXBkWHneYerAHFgY/jagfwwnmSqATDkmB
l+BmWpZ/gXUlayPGuFa+yatZBDV1peCtVu7EwnlutUz6/GRvveGGMkWeLyDsjqtcpYGbgtXRxiGP
4M4RY/F7yTXssgLWMyA6T/2BQigl38ZayUKa0FZ5NxuHkSUMOcy0uasKGu36Xfgz4g9f2SHAG0Dp
yr++UaP5kwyuY/OWt2hJZxeSU7tTWAA+VAzddBzlTJbTDfFNMdHnMluEYmPtZPhcnNgnqvQXOYlh
qfMaQmxaUuyEMCyAJVZTD8pwsZZaqz5gySaAms2I7/sKc6k+xuaSF26t6cKZVgolNolsOkAjxQ3f
/vI9bnH1lnBGqOoC0gvNRQj9BHxOUSlmKBld0RMYoomcJxEHyhYX+uOQBYt6KW2B7v2sLSLJunr5
WYn0lyOAu2GpLFsgJylU7Bf0cQ59ftH/Ldo4ABhHmTzqzX8Be/bVkR81eeJZnuqrJo0DHRcFfX9G
nu9OUOVIj9r9syftyolDe4wKQ/FdL5MDSFw1n1iJzs0TgaJy2jSkUDHIJOKsQiA2oDG4RpRllela
AuBIqbXbrCfcZvFUr9cWMgdOQovw6pG1aQ1YXl3qSMWL32ArDBv93ZgAdkSE173mFN+yTzYRbHIK
Z7uXzLPzwlXIHiJLBRuKD/u6K0pCBecCK7+YwNOTLcVDJs40A3lQ38I+HPv7bG4w6qw3WYoVUce+
F6ieRIAiqWnngYQFbncMV2NPnNleCR0yu7TSiQk2WmRkywGPyZJnqE1IL8c75jCjNEz1NSg1LaAQ
9JNq2CKYh7q/kjoOKIfP4OpvH2KJnn3AoYeQZN6GlRWHLIGhwsITKySNbMqpwKW5E8IiPHHIUvlF
rY7czJKUSgM9FXEkRGCeZgt+NLJz7X/KjfgXGdBqJx6cXT1JH82+jaT98AnN6gcdIa4waRNoJ4Mu
1wgBZX8NZbr4MTQ4ukKyjt48iCTacaxKs/5at4UuAJ1RysJFfci0b+SY6AmdLtDr1XyX9tTEM9gs
v4yB5hPc4UjIwkIczAHtwfubonU+gOcVceMv866jiNd93aqWjUCLzad2/MBi9v0iu63i/MKEgJ6q
FgB2QZBwAbuVZruBd+ufvnq3d9Y8a8nTWn69JmcSuGOPxYq3mqrok0+apk1TBI/7QAlDK7dT9cXj
j2EfWdjjwdSGUEP0AqHdI3TrX7kHx5kjAjc1mE0WV3B8eKoMOcxN5+2FKE5+AsUC+iAr4HZGumCy
v6WWsYkRJQjFsyraNtvqsK8gbw6qeNluZ8U8ftpGy5GRRwFp+Pmfckkeg86AoDUg0Us51X1ntJEe
mNOxC/NU/CX+2YUpyeFRL7BGlxW3e3taAWf5TXBE812oV6JijRsqzHgatKRI3TR3vFaIe7k6AGhR
/axQUjvGHD+bUigRqhlO2tZhqSQDHoyoWL/3t916szyxysDWBdGc/ivsrtbAIDr9CT8ogP8sU6+7
b6yThsN1KM/0pVB+m5CDgP9w0d9JI6Ox2/R6JIBHCSIw/tC6GwwlpUIdyXaPp/5rs12jYKfy7YWd
/kBDePl9G6ST6j12NDgFZQ1x0HpMR8YnrWCEvOqFmh9GWq2Yzx15dttZd1O14Ay8I+/mZdNvqAgl
8o9dCaC+qczf8Qe28NWf2ckgluALhtuW9PBsPfFtrqQlBncsZbgBaJKHKmQel8l2aOSYLzJ4UaX6
FR8uIhdeivOXq++n2RY2/d2Uzme8xSd2E4V5Y2+zXpBQRQS2OZRhgQ6jFeL9uPO549FHVClQ/4UV
TdcUFBvHj9zznvwcrzeS6tw9zRFpwJ/bb8Kg6iJ3Od5NvAJcLI1I7tfAraW2Sx5pbtMsZGOg2YPy
1C/d+zyHGJ+cXsRH2kqWPXxdXq5/7Qo80Z344VsRkXGGWb5sI1c3kEG2lUFSGrYClHNDstgSC+K7
UipLtHid5WS6+aqF0JElR1FyR49LY7XV873AZGywdyqIrFPAwwJZv12Feqi1j1pGUZmsXvG2IttN
yIRc29SabAbOINdsNNl8ANKqpfBGbmt7XhMwBrTwY9/0I1T3DHqHEEJmRC4aB5SXrTyMWy5SH2fJ
PQZ2kr21I40T2FCQPCbcgfNgnNTBw4FsPQxHORYcKsRVeoGdfhTYOYH+32039M8t4knc8zgFX52k
yA4bTmalaEW/E2cDfMFb9jHMDwxtOyFVTs7AOfEHyEd0NZwNfkuOwCOpEM8ZtuLA03ZsNLbzVEQg
wKXP8La5aBK2cvQiIgPI0UW3a1mIbipouno91GHp0JdhL43XKS/YgfBc68O+kYld5y+LyI12SAIX
aIwIYJkruM4BU0FsZ6JCz8NhLWPuB5ojykEFFQkDvqH5l6ugCumMmWLrhsk6xPzltlMOIgN9HaYW
3PtH8bCm7zL4Ct/828dFNmZw0r9AX4SwmcInLWwAV0bFX5cEtxzH1Lq1E+3FR/QkAI8cfLCMPLsZ
KuPHz0lMFFCl1gcODsJLO+LhvKCiT1IlqkFfQAlcOSfvxXplQgILRlLToyL68eldxJqVwKxjvX7Y
R4Q47PbG9IfdcRA+ngWL2ZgoVCQT14Zo3VcHY6kEgpxh/N6H29d9FdMWG0iML1Rz0HQc+Ftv2cEx
nlzY6E1Hx7Af96s+5QZo0pBXv1GbmpAW+rJrAN+RQUmhbNhWCiAmjNYTkOOTltiN+zVLPRyUfzgV
bzUntqjPWgmMqWaYSn3lnEDOG1PwqWalI8AqY7U/zs2QjZ+LpwmzFM+WzFvV2BB7NyQExLD2HOp9
z/EJTVDHCQ/l3uT697DzGSKJ8tzmkZEPEMF8YzupI4jNAJdHLgsv6GhATK/+UAjkbRgswMkX3q++
jlE4eKm9PL6XYxmJqAErqpYJdrklJRpjTHcJvrghJrhNpNKmL1MsCcCNvgnTd5oLHLByIcozgQDO
OmcgJZsR4JYE0YBIWXDcVDH4wHuJZ2D3AE678siT9uEbnhyHckP7IUzlFKSLwc1dLhjU5ew5B5Qw
inGh6/U1GYqRjQdMEVcOhZ19RGGa/HXPESlM5GvDp9ANvQFGk1Acil/ZcjaAYeea02pcNQOpLbz3
sqnf/VBqU5gq16cODX2/XZ5oo11InM6EvdlrdHwaQUVqZyjDcKXhyvnKLIpdDG8ojdDURfnnsJpx
AHfW/riHMLFTzqc4d6OLQB6MAodgo9xQoPMkHrmUalHBrXCLx8eoxZmONWfEs+uqLbeOm9g3HWdc
0EFphGR3ewgBCzPv5kEnC+iba4f7JUWQREW/m7O3jDVDmhMIXGsuwss3/LWTVNc/3lbhmBFZ5IUN
ID52jBaCb+CnZm00IqVkHN0tLXEKjvf2n4JRIAzthmYRF+d/YuhcTGdN6fW9hP/5FjoEnAaKgevR
emR4Ee14hOeXWhYBoWrA7hujBQoEUkkHAVaj/pW5AqjUJIoL56bPEj5cePsVwxWM2dU4Yq8sF8DP
Zl74Zfj+b/Gc1g3NCCRnkL9o6G3NftjAA68yeRaAzuJT6NkSmcBiWJfm5V7AmubYpzpM/hpaeOb9
bJFE3muMPx3BPzCihGIYfFogwLf5pT1/O+FrdZWN9dbsB9146XpTdU38o/S+vpZIj5zrrIYq3Z+e
dcdCA1y3oBynu2j0BecVEh+mt8HjL8iUdlLgQPxr38EYoI8vbycoiszhAL7jlWoVag+0fmQa0+pI
CHJDK6mSlDuTbjlFomG2Qnq+9EZeaKnQb6sygREQcmh6JACtDaQhRF3Z5cIbHIADrmIpcuuclUOu
YhvjcSf1m+2hp9UP6gazMlnQOiTA9byCrCtxuh8zUBI/GIutFuEfCluwt4RtCtC/Bc9lSdvhCr+2
dt5I58h20OAnoqG8MCOPfluCfvjOKYEHkYTkP4BhpvuHCM8xVP6yIWT2jqsatbIYgBWmuVckCOAv
9culWog3X/P4itu8mBF7zbqQOQ0dESllIlCJCO38NjPKV5E59Ga99NMvweELVlRJM+bJlBGvGlcK
OTspbgfAa8+zk+/0TAh+HUWYznZgiQ07mlD4jZQPpx64XwX4E0iWwqMi6O4hLX/zISZcFE270Sw4
7G1UvONSyfbJznJb9PucmdePmMRa7GHHGFv82FZkR4mCzNoA6ip5xAGwIGWUXdkGoJdXDzHFDhLq
1NAIC7MDpJVwc4yUq14mdtKXIAeKajl5Ut0Uqn9jkMqyWsHKBE+5Ym9pQXW++4uVmbbnbfIX55FE
tSeP5J6tdvi5/f7x7hpKfRyi+ttaeonTWZttQVrj/2Ls8l6713EppRvX/S4k7F3x6ewzwqU4iEJo
jCyTJF3HG/Oy7Koe0UWbpRSgzgZWWGw1wNi9iOD06vLm92wgVSmrNQl2y37MdBs0rWhBdsX0OayO
Mg74sQb4tXK5jtKlCXENe+gevQOVV9MC6sV+r/sgy9mFIW1CIFn7O4gB+kKHD07uc3grCKkeR/9z
yAGCH4n1Zw4f31XTUTSC1YyWgZrV3kmdiRCa570knm1lXMExBvvNSbrwlocgHe/2HPs71ezDRgRE
D/5jC4HBXBxxtkwvnt4Pdm0s7rqEneO9XDroDMcUKUqaJ7DruVkBbBbhtEGeH3M18uzNnEpC7NXw
a2EIUhyrkuzjVW9/T+w3PunwOThK64BKOJ4XezXlmVZ62mhxi15mVmk2WWtg9E+L+QzC4w/zKeqv
6xr1yxb+nOdr6R1i2+dx+oQf3FgJdqRZ3onVju4WA+ZV/r7SCKs6bOlqwmiOIGihYdKtkff03I26
FFS8h3Nm6JtKwv6QVJgJcpZipA3fSAWteBXazFTYes96I7UOnyd/DOJ3gloiCbi4jUhrnBrqxLFo
0NLggD6Xnprzfer6yZ7HAQF6zoHh6LLvcgsQ1bMdJ8Mw7TVKzVzhkSfOhcvgIqbpOpZ2KNkOkNdk
cE9IXKUm2d/cKxaGjRiwNWa4wXI26f7ykFHqeTF/im5KmN37opS5aFhCVzrGmIBDl8Qkxwp396YB
PlH8uoQgGoRDvKoYqsF+NO7q2t7NTS4UF/Ik3+77Fvit6iV8l/vJ+o9uru6yAkydTdDrxuNFSVJY
2e8XwwlOrVS3MF3YqY3GdqfIie9SRATyxYSgrVunCori3HM60LluPWnYg2JouogCw4dD9t7lJ+P7
5rFjqG+581NuSViqQW0aNj2Soze6/30GLE5HjmpKoQV/bpdYxG+mnFI16+5bjAzxsf47eWN/65fx
6jlrE5hpgyM07RVPsHz/23IPQQIqnGBHW6luMXQw59Sn4HegGqEGBkPeafTZ+OARQyW6Uld1Ik84
+MS1BUbrLrlRnNMy/45leWMwnCE4y6+DRjqRx9cGZ7+3U5CtfZlkRW9qdmhHsYHhGs7NgyZ1TFj1
KC65i7SWIMM/5iIl9xE7qZ0t8LTNdLkrfcKfz9w856Fov5MHRViBoaWLAzOmLfZR5JBjeAreIeTH
9k0EfQwBP+rnouaUYP69CC17aJ2ChMwYjELNkCOD9DZmn69I9509pczS4zLToosQMafUInN1yHzm
i5aMyi29Wn7k3DuRRUBPYmxpa1g5OfdODSbdmruSmnJArLiufzjOv4cmEvfJUAi7I977ws06qnoz
TULPLcz4fsj8L+ZCS6MYS3zNmLLm9HhtaO/7ma7eXtzDQqAHkJhBbsuNMHzBbya/D4IOLhHTiCu6
kQ6vrKVB5DTS2XihNNC3NdGecs7rUaKG+V7UNOKxNqw9Nncs44rCuzsfIxT5pQcYU5SEGYJ73M2t
2Nylxs+cHyK6R9XZG0Dzkd0Se3IvcwUF4MYljxJA/JICJ1RunAtw2aAxYxe2gAYJz+zarfOE6jG5
HIKuoIcs9AaxX66Ryr2xCNNua7xqtV4WEjKxma0lPL6Wkq4/oRT06VjdgVVosdYGtTOQ+cyk7+W6
s/obyU3xT+b7+IUCr/pZ0y6A3wzbfryQGXUiy63dmlj7EViek6ectKTUL5pEAir+oG5x+09OLZcJ
S+kI8Igjtq5a7EIDcCunZnNAoExMDwr77yTYdL8Sb1pYRDCEpkGq7YcDIJhBL8uEahfGR2vw/qEV
gChoAvOoVGMpcYLOeup60rspFlaYaDFaNtLh09KqlM5hL0G53j/axCgkrVqe4ziYSAHf7Xy8pc3b
viRhTlAQW0BFCwMTLY8uEybvqo6064lWlC/7KRyzRcrZ5c3CrtGHWDKdJ7x3Pz5Hgyr4r86Pwo5Z
zzxl9Yy0jnrCzlW2UW6VRMdx0COe+qMf6WPXWo3O0WEfKYLA2Om6d18KBxAmtzP3ehPzXd4SFnyI
nlNjfySkzZcELEj02d9eQEH7yjsm+Gvp0FywkycPhjsc5MtsUKBolJbdgG/CTtVM/0vdDh8kx+Bp
CVxMxvXtmtaAPU7VMwYkws0KpjKE5ill7yM2u6pq4yVZZcFqfJO5ypkTiqHGvCa1kYkbpi/OHrv7
8TwspDkeHFfw7YFUNhuXUieEObFv5oZpALcYCLbO6ct7r9oH4cqCYwbHGasx0oHrO2s0iUUiKVMv
MGL1PYUycNIUev1/yMcxJoDUDCWD4A/Sz035d6wDLlcV0N1Fl9Qu7XlCHi4a6DImhL4Vk57IL4HR
QrcKqNfKnozKtzRQFQXJdjqlv9PVmp3I1+fAezh89h/ptglyhGXl/WKUT6UdzAzPfcPi5x0yPUAw
IPxlbpdVfdiA8XNmOas4Hpf2lPfBWK6cVrcKIMOWxn9X7I8Moux8QsT46PahQdAxB1qXoXx8ULHP
YXwumKrWVGJr3nJKwA6Y6Vdf24MZoUWARihplnrcbCRaJp4L+m8pCQsNMAnu4KryVpo+/6+A2D0T
h5erKBx0UP6gKEyemjOrkOfEwioX9bYJPppxc53EK9F8VVH6Sb5bv4etSDVIOQRDUXOv01AzaVQY
S9EyLaq831pHVOdPCuIIkDUZY8qUReZx2PoHcq942G9t8IABIjzUCfR1goKu3cyO1gdOKAPPyl7F
HLf5VOSL+0HC9O80yeZVNPyx6+gzDClOMuXbDf0C5RTzCScU3ih2lKUEIO3XQf/IDLF7YedTJJ2W
X40CxMCT2mjBwYweQsHPgD195apbXf8slim0PXJZXvYZ/pVHe3aN4JjAee2TYZXCetlpxJP1ftvR
YlsYmL5w7X6CczMPh/DppDYFLQhOhZtAuIgBeTHFGsM3O8VKUUHq3gNeruNCOUo/oN6tOJ3lVmIR
rDRboX21Bg3TE/Q4CBfVfv6QM6XjkKmQ5lrxGVCHpcEFSf3bwWoBo+6hb6R3suISAT9pQAWjwsQP
TL9fN40WRoGh0QSz2WAo8HNWfuUq/MofQ/MTdcSyqtovCR+XBjtIpznQz+NkMLqu/xddxSXpun87
FYn3+f27EbcKr0/pchlmvX02m/QP+uF16OJTQcEB78ql0mYA6i5JEZhnmiyhmnOMEiiQInSBSO+q
cqinmTDXi/pRqnRSqIG8j4/IQoUv4pn3DKPXwaFZzgdnOyeSXsw+e4vQZjGGCvghSuHYOt57g2Wy
ZSLU7NsQmUfN/qS3+2KNVVsfw6Gr1DxQiknK5SBDwvO+lq0iXFLYbK8gjMfVWy/TKRe/c7OjpXUV
Kn3WA2SSjoBnJbagOj3nGmCoO/2VV62i5lgglp+t5WsdNsKtnch0UPwCaGU8rh/w6bld3/TRQYEe
8Zypq0VPkkqDkvCc4scLnpMIEZ84BqGBUyZwPJd8hiSFv7mP8Hwfn0JNXpvGd8MJhKDDwgdIIXfz
buuRhh2lQvecusbU+Ixq8wGaDk7yg0F4PetCjkiJBa3b7pgYeWyFCuEAyUf6rbyDxOzMKfkZrzWI
c1YQntryBDIxHe6dWsZm+5m98fdTmQ9jJlv2Bm3ymvkiWW2zTYLA6PBajSG6w89mcanqHMzjiIPD
I9fAJ2grtsuTwLsG2YiXlBW+azhBZJsFEGa4hAvqCdWX8OwFI1zdOBNr8Eygqabx4SXMHsNx9wlN
v4y3m4pSzJNefoId8zOTqWxTEb9ybRRTtywpnzbw77YOMEQYP8wuyOSeREBW2rLh9xy9SgHtSc9F
nBRLipu5Xw9/RAL0IE1MCgB0kRNoPWNjxB6/RBuLiIL90gZrFb+AlZmSbM3C97iIqdz3lzWRhstg
gtEvaxC/uegYEyjlymA/dA5g2TPuPjjvdI1hA2tc4rggommQMrgv4bM4RXSFFtdYz4cEz/GfT/1/
uMQK7o8rSxJmjhbZanum5su+2yTho8VmjrRnORVpcnV7u5gB70R7Dhx4GLAFaR+GDnugQxs1/Ztw
gktvvbY9aE6x41/j1PYfjVagyf5Y/DUoyDDwjdtm4xa77uPWmBTZD6FHyZgqqkpCkFWpBWB5+GRM
BTYLsW/bJQ37ft18sf6Tg3/9aGIxNmVDhsWySYK3xNT0id1W8yG6XCEhxeuPJ/k+6xMbMZTcqz9I
pgOBhEan9Yb84mR89zrLQECPF2Ek5Y1nvjHN87h38kBhJOEbjthjqYmrjWb9tFODMXWuf8eGyreP
DtwXv+Y1RPi1m+oOGSuY0W6t+Tw47grwhebzJ55RA0peSpnuhI2TF1Lfaze4ee5oaD9hxG14KNXl
w/+IGypvnd7pOkd6thcI/qmr7Kg8YM/UH7CTiYF1/SFUVifUX0dCmD2DX+MURB1TwJ0GpGsJ+nGo
INcaWGSOYKULcnM6caLhPOF8sb+RrzRDFlQOGMC9K8N5j8cvbrmzLmr7A/hTXJY+4mzKjuoUNLjP
wmOuGnJqfknSHvCvXI6oLDAcjKODhj7wJLDbBxd5evmEEkYHTe84m6+/WNj/Pv/p719OVuQ5Ex31
MWtpDk6nAUJf2YWOdphTFq4BD9tQ80dClb7nUkIMkqW9bif7hn7/WMbruO9b7MLOqFLqniaXXanx
kAvLRHuODAa91frjHbokh04TiGighOAd8qcW7kOfmP21qWfozIslbPknFRB5ehOCQspk15/rA2xu
gO8makSguRYlYHhhzEUJ3Nak2RULuSqxjAz5sBhCKpz6qpisM6oAlXQKgDviPsD78hglkj78dyZn
bEZJrEEM3ywznjwyGfKuxRh0fmuHePl5ltAvwXwT5BEO+TT2iSIHiwV87vjyXUyZ5LIJKo+WENBF
UeBsBmof8IGa/qMyB9ZztFQAJz4uHRelPX7rCrn2mseUV+Kb3HLgqPs92nOQ7KA/sF8W7o1kbRN3
Fo489hrP72B7W9xoLwKF7ArifkLAAOBkUj6699MntKcrrW0y/FmBrDZq9xeX1wJZbtVhYrdYAfCc
Cuy/xAIyCgZkvV+fPxd4SeJvzWMgtJvZD6pzYYt2Z6OdSk+jj9ZRRJG1wDRTX5Qx61k/pnlLWcJk
K+NC8KYOjiBnzbMM5RWmKJdxGCsmdyDsW57Ft3yrLQmhYKKYVhxyHFDe3wzvC+YUZAU1SOkI3rwW
ig3HGil/ne7jgJZ5BOrC6gTp6pE4DdoPX6P60zPkDx4dQ9Q+2p/K4YTs19Rjnliu91OO8l5jpJM7
jYe1fX8kLxUOg9/jCmuvmYXEw9eHgecE2zR2rhQVMhNDZVxIVToP58uTBXKQj0/RdFbAcZsCffYo
3TjjCDwi67eL2fgtw0GPZhew2AgjkLuG95YEYUozh2FrPKrhtikwlbPSUMrP9GsPClx8bh4/N4P9
WUDoNtOJhfStnPV4j8mamIPWY+jOcPY62etGDlKWrcc04bBg4UM29YNorUyAFSQXBKiIpX+TuTwR
HwoXrNr/gA3FEKdzIr08hOefUQWamFrNjF8wpjGvoQaJl9o6qu8wPur6CARSCI79hHhPHK/y0CCd
7MkbKqsdhTI4mQRZVwsUpUn3EAFToXJ2+H+A/2WjvbfIJe7ph957TY6STzpkB9JPPzEYS6O3c7/F
Pzq+KWBOXYwWjG2Wh/MJOYmRQ17hLgr9O4tT2CAYOUIHXuewVjkU3N6PVp5BD20tbjlfvslVjbZK
1g6ELuQu+4xHLBqNgGcuLsxYERXfoO/rz8zo9PPGjZnr3zX0bEwoQpkdH0bREwFwartet77p4w7r
miJVPdfaRhMpPCnMjpew92Q9Bdq6Lvtt1fHBt2M4U0CVJ/oVgodtJrspoERWXoi2QWqYZiyoPd+G
ytUNIcit4ekqwgSL/bJ9kpCdPYf8vebqR1HoGCeTUVPKQLtynV5oJp/m5ft177Aah0y0KOyxmSzN
XZORYTIBgU08DrWApBEHUs/v45xqeInr9lJglhrjer4GqhaLrUyohP7hTRBwT4GIn9bEjXultqDT
PclZ5tXktZsAylXGllbjo+vxE6xMt4F0tS24KQ0fMAJbLPNZFxmtHoaloUMs+PYKRLr/IjgeDsXy
mwn6RZU4g/CCkXp/AHJqYT9M5OxbXQjeE1VgVtt7GSGnRacjqSLDeGAa2zV7Jbyla5XFGh+dtM8/
tpGZnEKnD9WdjgYwQkKp8Y4qVMnTZCZtQjRiAPJLsEUY7e3Hifl9cA+navjQoJltroQ19ffDufK2
vY9IefuzHWq8dYgs1FQPCuSM+wFiaWF0dc4kGqjjYtbvzZZ2OHuj4Z3/u6CHRyK75Dh8R6wzeOi7
6GZaHrCrMrSkmSeAYwrW6U7jt2r31H3/X2qQGX+DpYtIUb8QgpYdfjZEb14xjCYWILLDjzUhCKJS
mewAX2p2xobz9RbaKJLFrM3mFxqwAzp4VyGNIBLgMDObPMmoGRcVS6XG7f5lXBjCEhnsrPSHuoTP
9xP1G42zLsZqejnLijrdMOlq/8KdLj5iGKGj72L+/uC6NrbeMQyzYmXjASb3bH4qmAofsKgpKIUO
iYX1/+zgMyh2GKhg2N0CZe/coCezzp4qgh4fygOmtG1Jp0iXg6PbPDt7OfR+3k2KEKrFZ8kK40y8
z0ol0ausYB5hBs/X7pkniKgvx5Gl+Qu9+Q0+eNug8rJI2R7j1Bjjwsw/Y55+y+eCwBVw1swKg9+A
uCKlWn426rC1bNbwKqpQfGgT/wg8a1NAh2xxAdBs2nRdLmsqcrk5Oy+hkdRtxorKsouyOIQrl73I
y+xsIPWp3xCntqMk9XQgDw0Y8g8avSqw9vWHrXIgUb0wMMW0DK2e9Xhdmn8hjD1z2GTLZ3xLT91P
CzNaWcqrOgM1Q6UwFUlgW2WOTu8H5ACkrP+jPMzwuZwaaiGnRWTBZnle7F+d+HMB45srHBiy7I4d
XsygS9tICUpyc67271nskd90SNceMTwoldmUgO0hWsX3nxc6w+SY+1bu9XCeb81T5pksTcqFzs5M
MLwxrkXHVZ4UhbEpRfwWdxwp+BvV9OeGxEYC7E+QHTBQtdEMKMWYMpTH2IMsr4q5YHdD4fWnn2Nm
g3PjXbQEya90R473kwZtwpzZ2RLlHImknHu0npGcPPh8rJ1XG2sw21fh2sqyMuSC2DxvIKiidMfN
yd2nv3OrVnCfTktEkSBER9hBcjuKEmJCB7SEO+wWXC8JA60S6Xkcp34jht+OqROOmb8pMIbbGP1w
2joARU7GxF+B9MII/aGD19/UYg4MyFmZK3QGZu5oowoSZRx4Z7qRDfSG68s41phGTJvec4xuReV0
xUqbxkkLiuSPmMDoxlmXNWXnhIXndcxc8FZNv7zVo4WelguRjXXUmb1sP48LKvemBlfFxdq9ter1
ZNOV4g+8JCBfpYXqcEdWWo4AiycUK6b1//XMriMNFzv6OlfSkwnr9NcfFF9BAO/nFgJMyfR0FQOm
9as4CMGJI8w23bR+tgq9nbQXE1fDRqQnYH5kX2Wml8tX6HHjJOlLKl1gBCYETMSW6U1EHYHBQZrU
Yp1Han/Hf+Y+UXBYPUgt1InwjIieO1qT2ug8xws+McESd5aS1lE6QV1kxlP2dehkngMTpZML3O9a
TChRWH/y+Y5Fq1ZH3rLtin+ev7KxWPkdbFNLwwbvzgJMT8d/mLtwNDH1s4SW8s4oS0XOUDubCZfS
79Hls2EfuA0MoBN44LhpXf6DVrRxFh15vMSKrbPHjjjd4iZu5OkR/Pa6CilJBTsU8Vk68lz/Kn4Z
H4/o1s6PfVi/0Y5CMo62vgYhbuMGNfyGb2KuxYCQWRzDUcSzG45BGrpc9O2yronUZRxxHcaq/lKr
kzw9o/lTn1Dib2W+zyT62lOkbHwvTMQpni8/jUw9rxTqzepKbMlF/hiswj9ETW4s81EwbDhKTSkL
ikgXuHBk3gNM0O8NF7Sy5ELjMV/xNzue+NgcxA2b4PiIT1GXVJG132W3rlSdB8Jlz6wM3Vd0Y6ge
Oif1BKVHN1kO5Gl7e/IfYLk2ZMjBRJytaTCWCv7ZXOiP9NVk/hK1ecSbgCeJa2PWFMsnsuUr9g/G
hCDjXIPV/oIC59I6iaptmUiDVZ3zzFKuYkyP7pkF7ygvMejLTcfO4SVSDDVaHZg9P86nQYfcaERo
mh7tiSM0ogTaYJD2XbozmUWYMaowJM/jzlysKOq1rsWk6nCnp0ohErRdmp++gWLZrGdefAUBu5Ra
IUmStWttkMuErcvu6UORnI+dBm/C2+WC7YflrSQCu4naLKLpPhgBi+tNKpSytU9IbLhTtay3bNTD
WLbNTSTVUo6DEphpI8mgY1Glf6f62mCUuEEykFaZjgF8NfjAM7kiiuJ5ukHsM3cNDanKNILKR9Ba
7oNN+fopGHfOw4gtUgZob3QyBVPjnVwo7cEJrbzOw4RXlRLAmGMCyFTToSyVEqGHZSvMxFjoskGS
EBGhUeQ9LqtOC6MEfWVjPggZLZsatF+JhbJjBhiUkjvJQIjwIzPUEieHdhn1eM1bNR6ziINPiexZ
GpFxo2n5G1QfYKqWWeA5XtrnU2MygWl465cSxnb/8cHYPsLz3tmEoayQSd4SlirUgsKTDD0lUhmM
thd4uLarPW6XZZPfeoB8u7BrU2JUGXKwoj5CuEkLbZdXunLfnsJV0cGjEI5fZ3+2s/W8TJCrLM7l
h1NUKIqqTvL1WEYFYa13bVjZOpTfE+jPqWZb3djBiHZqQ42ENlggwaXSSkH6tf7HYUfxPU+Hyd+c
bBgksRD9HPlUk3A7lp4e0YEe3YyRsAxp79jk9fXe5Dr+ndhYkbe9aSVl8ZMPZ5QL96bldyvmCAVi
B+iK8uA+8bwkk8EBWh6DIhRnKWoCV1+Pk27PBzE1pJeUNjtFBcN5lrqpU8N8NAB2PncoWMoMOhP4
SbI6VE/RYarN3aXt/O74jGCWF4+pgYsz9uzsCZM8gPBTwYcvAfd7im/hPbMT0ZqRxiICVq4fAccp
2XhB9ewJGp5F4bd7SemRSJGLmlfDxl62PAQjlgkRFzpwUBo0JRa+gJq+q2wRYSprou7m0mYVKiqD
stZE+5fbhbsJGyoMDoYKepsRDA4Uact2y7iU5h5w13kaL+zyQHb0VqFXeK1lUfyqIUtCLzX/UiID
UoQnI0i3Qi9ph6dXpQPj2IBUabzwCJ2ggimWTVIPz9nj+mLXpvLIaUuYyMLdp7Slzx0zdj8DmE7k
F7FwgNzwCf5VQ/NcJ0agHRhKSr23BySQfzavcPbxr0l1v8BMbTtuN0pGalTjecyNx37SLAmuVxPP
DIgvrZY4nTc4ImMCszzIvbtvGyY0dDN5a7lYU3XCB2mJsSLyf1H39pREOTG+W+bgTykpb/EgqoHu
sfGazW3DPe/Z25Is8ArfunYVCwduNCDBoHFJTuABHHhmhzlkSDG4aIE8E1nwZmjJ5mZ5yjW0C02t
sCnONW0E4yluBtbij2B58RZIyKnlxHXDtesZz0CnjzbLrnIzjZXpOtezPxQHxWmYjO/NiSWFy4zv
keDytpRgl05Cu91lzOeYUsiDs8/0aFrxhTzhopt1AThOjsKYeoZZQXGHFqYh4DkgFySANJ0RZRTw
QFT4lFWvU++FQMxtdtoahBi2gYY+RloX5dRqQGxNz0LbCZbYcoOHKBWeLXdy8v3QFEmpzV77tga4
n4ahSUGmzZUoQPNGffg5ix6o9eXFtwYzxc283H4yBvq7yI9zpl9ngz04DLHsOlvPhsI+17NXfC/V
E9oUDVLyKcCQVrlqAV58IT+RbsFrrWfhSEVxU4uR4MPYb8LvFIZbQuPDqQ/jRa6xx4sJ+6V5qeuL
YdJ6GS3atQwhRQF3kTO91fOYtHsElXOPpe0vdbotOCNWDAMj3fIkfrvK7j+uVFgqFfj2maJvrkCM
ZXSspUbZbcZy6uWdqg8i98L4E50srdBybihgPkOOYl6okEpWhcupYap+sOGrv5oA39KhsswkptMG
MJX8lwrEfL8uwavbRzWvc8R99SnrtcgTxSP3HA1IiKYURGR4h31dEb/EEmqFkVw3IY4PnQOuQg6T
Iva6UXjLt/I8I4JntjnZHEDNKHzV17xCvdGVcHsPu6yrDPUV+u2NtnaWP0vuzNU+HRW6vycactA4
8sAQUA7GbqnNeVBUzB4HP3Jl0/NZ5/F+XzpyBrck6Pfi6Y0nQtqoMo9cL1R71XKJBQDaLblxiOUu
UAwtm60n9Vk3f4Br/2FVkBPvENknvwGCbPlqnCJ6O4sBWFlTURIidNadtJRUQdPzchMeSrfokeV8
hB9J+ntpYbg4DdkUTfTrZ5MZM5lHTAk1tATM5gynXuwAe8lrEjHHpmj2dXaEJt2opVxu61IL4zOL
LEqATNC/BZQW7VI/GyLFBdMd2SfQtMcbzLmwRtlPEVxvK+T3/bllE6Q2oQjHBuKbnIvLFgkGp3xT
ba/Kxyz6IUmKDHFXX0nr+EMSKoWDrz5NDygrhdqODNevv4zTKU3pHheqME4R67zU9e21z59z6mn5
0LYo9JRg+Hon/loNx0qc98eHfvgxvbejcgGZlqbFuP+smNp+hJ0kCkbvZpTtMyrx88Euz6KGF5nN
dE/qfU544GWEsL5iHpN+6l+/1NP7O85eZBUfHzoc68nnKkl49tjfUZtIW1Tm78hwHKZ/V0s1TVzA
7P3skTLQ/3IPQ5LZP2m/4YCRbt3RvqReS/K4QjS7UUTmyfYvE5zNDvbrqLLLNAEAkUQjzyq7JDqd
Cf6mTkrbvEkEczrqmaC8OoHre2Y2uyzTtT8ISBxy+PZRiK6KTkzRfOJ62LLl3xHexvPyUQtOr9tD
Kclyql5uLGnmyutkVi8exTIg0BiCLqtQpvnZ3KI4jhUun9bTR9gQDUCa9MlYc8oJhveFwOVceiKf
yL/prnkNe60t34ZhszIbarO78a3Bgw4q+DZFEzTLZy/qkda1Rw/5ytpDW5HcqgbShnXnpHmmiEgF
Ve1LTiXgKvxbuYekG9lvTGOl1AU++2cLV74W099VRxm6+KfXeWI1/fhEGT2K/oPuNSj+yMBmZJcl
/nlsuFMeJOOoike0gWagExpJtIZ+VFbMf8SAlkXTYe8B9rhZxYNqnVvbKNEaPaIaX/Q0Szx5sDsG
Kfgg1iWx99bCGLUyWBELG+RCASThcRctP/jR1sanO+Y9Wn7+wSFLrEoPH6bEUs5C+EDj/JWBKO2u
L167Ukvd20tq1Xy1PO2wxxvNkGdsQq4+IJgkI7LMG+y5rbjYkqtZI7MUSNULNE1pvRzqObL96H8+
lXKqymzi9AgyKzYyaYPOlZLkcDDpfkickbkWFaNXzxcMHw1oxArcZriHlssvrP5YEigebrOI/AHs
pUdr0HTR5DBazZY/rbk1Rp4noA8WjWKvSnAeS1evoHu6uF3qqehN1DiT5xIjpcx7SnSgrlFPt09Y
mj4pDXH41MeVhzwaPDFjfShnim7sm0+3pupDzX7kBKWSCyIQBpfGe0LEysugr0JT7SHEHMCsLeLi
KWMDr+elHNcsvf9i3SxYvFnZ7qPZYW8Akv+Hd9reKj0LnGzznJezfSgcZ6wkeaxpV/Grn6I/vcBe
rM16IYzzrS2LglHwuRIQSj7fQBXaTO1DMNCogxFTcTpuYAiVp8O1m3EXWdrHJRIdSG23s57HXUM7
mtdR4sUX9BJL9nd19zoUNghMAxYaUnImtL4iIkXJ7Zy3ja+oqms/ptv1quZfkc3d6GnoJdt9aaWm
dmo1XSytU6qFYKiT/pWP6TJp/7tFTK1S7ehBu3+1O0IRpPbiX+JAV73PFnVMo72ZiVkKlL7rUfOA
HTyQoZiIghQj3Ktk0jDcGqjRvTD5krrcDIU+weHnCOn5UxsIPG04fxHRAluCYTFlGl99gqlsuWyq
NDwVTzqL9rrNIicZa9Rvp6G4CT05cndD2au10jfa4eHIkx+wYfUEGTCXO4HijDG49S3+kyAjKZAH
sNypuAZCSOyXSZ+CHTwgd0ODRM3PU4+cySdJLG42iMbBCqGDZYNE5vXATDiffUrD3ws2Z/Vq/cXY
NeGm9b2Un0lAiRduWw74uq755vzm23tJv69Lzo/W2pb1i5Mb+i5PI5d9TYPbvs3HFpbNt07GnNy1
8hkS+xV+c65C5/WapumVy7L07CCd9D0qp34/xmp/1lnPNsg4zPOBrSYz9RPM0O5ZDsl7TV7Ygs8r
JUbPxjAeufJJ3Jv2U+Sy3K+yxMxqp/vW5jl+ph0lM/p5luda+f59V75PvInLWWOBdQh72b9Lcp12
x3FFdT4VBaqDWLnRnM5JLnh9aOK+69vGiGzE4LGo/ZtXnN7F8Nwi/4HkIFNsFpdE+kSziLu2btyO
FXyMFecgpvLM3q6Vc2ywLR0DYmITozLij41e4s3v0iFrztkywyIsm8joPArTUYJWtLmshwTUy137
QpPoVTOIj0lTmOpIta0jP28uuhHsAYM91WQMJ3Apt61GRRkswM0bzJ9zM9G744ksYDx9g8oOTTDU
0pl5t+3SsFIV5YZxVlX+hwEET4SQT5YKRDM+mTz75lKqxQS4L44HYkZX0ydEggr8RtL+PmmDqQDU
/sjbcSIPcMY4ZGLN+hK5GIUQDzal2gShh1H5UqGrhPyQs6+kI2fy4wSgFqe7N6/P+qumcd0sG6rK
qCKr/AltTEMeu7OQ5x4s/C1CVckm/ZmvZ/Qjp/0lUQcxBO9bERChlCQDZBXvqbichCaAF67/6PvP
Fcal0IkdJbZyA30Qyxttjjl3z5DrcTrSown2rhOaCFl6RF46T1EUq05MF0P25hk4caTPYM5e4Uqx
Ze2nmtNk/c0FrArAn0UKjVIxJX7iKKBVvuLRetymE1TO982VAd39fFJHK1BxMSEWpxHBHHypbCtW
+4+XPH4qUHqRVjcRdmMt0Ecp2xyetjDfwB/FA1ooWxzo59ZnsRUfll9muCSOzEIZloyuiD+6tLD2
ykQCOBHJ4bgwKe2Yk10WWTMoxY3wtFn+xUOuUjinvC0gl2FLRxDBqBc4CWXUFU19448IoKGr3Wbf
H1Z308F6gUEDHlu8CEzJw4kb4cAf8RVLJRx4vSbLeO7xmZH5jaFJ+JUvD/84G0css59iU33MhJoa
CP87WggHXmhBAcXSMSVTWAUf+lSeZZiFfVvZS0aGW/uaWuP6pvXmGXM28ez4SFzMiQhlnm7KKulB
xbINPNed2IrqIpFgxlyGK6y4PH9SOjAOtbn0/IScfoSmt86g+gEXasyW7lVIwusrltzVbeCYq1lB
9p6c3hgXiLEgOWSXpRuvERIz+o0lNxIwAjQfky90wYsSWgmRL5vo1vSSrVlAHuTmlPZxuhlbIAu/
G8JOAwieBvesl9Zz2Z3ZYu/WpiudpGmUFgNmdkeyKV9k1E0HoFTB04MXyZRgnChjvFNWWACnCRWa
gDgGbmeUu3VDhKIp5CM72fr3VvYq/jA2YRfh8W7zzDxM3WmsTr0wnohZTfKjddJvDOMejim8C8Eb
BOwfsYebKJFgDDJfv0bz9suCrBTqEykJWoJ0h2O9F2o3bTp8KNJXUsqEMc3/bXcwYY11kjbdvYlQ
cLaV/kgVyTZ1rRjerqU9nX+ao7giz1kNnZ4G33ke9ALiH2FGGDCU5LQuK5mXSCOuV2KlMu28rRxH
u5qdAnpl54vsu0n5kYLj4WOnInRGELEiX4k/m2AZAwX1nAbs2SI7YdsIls8Knl1V59N73rOJSqLJ
XN2Kn1p6liUVUxtqsbNcNZcvLaZ6Ziqea4nDeobkWEYmyXpnXbzFD5/eK8wtkzE6MddEy83xg+wD
6FkJR8asTmAPuyF+u3yEf2FRx4duA69t4EbBDgUTSUmsh1UdAA2k2ibsaCi1Sh99qMZrlQ4uvZaM
ctbiyELSK3BARM0rlQYGMLCN7oS4B2ZkxQzr2g1DLuozVzMuKAw4gnok5vXxxRsyQNxvkeiLhwr1
YDD0g1UUPeXbAc22pm+arfBje+TcASCu/B/SBCypyh4biubQ7YIewSXAGVwT7nnyvyeMsTvykSck
OS2Lm2EmRwOlfL14XrU4MAaS5U+FesvxvvbmvOi4VGeSzpFI4x+NUmJ4FCPE2jwDsOBPcaAC4K1g
opNaLp6EeDVMIVTqRsg6XdaaJ5/Rg127YGaIkAl8lbnhKlbW9wX85+mGsQEAANLjaNIyyEhtQXc4
HcxitETnpf3Zko3wcoGuxSq0L5w1I2BG7jeMxMzMNJVAmdqL2MGXCCOZz0zO7WBJbQfjBaTsmTLm
ESa0yUQeXAdlZe2vQl5bImZhOLOLKgZCqjG+ylM3XmMjsOyCDvXlgDgNExoe6QHpS14ml7oMQ0rM
NLZcuTPVtQAtrHlAp82f9t/On2wEXVucu3pGR2mOsCXqdhmoBmSPbuPBjF+LwQMVOKRnXNxLKVuq
UFRaxEo2HaixLgry62lsyG+KhD1gEWaZZ05HEcE1zTD0G9+dQpKYUmVAJMjO7PZuTiJWmHt31Jbn
nUgHaZp6rcxkT6Om/BRnM3uGdvu9TNf9DOtc7M1CjYYLz8zOOxmK59eIbNUzd0UsFgndCqBzFqLY
I932tM8EYdkFoxfyps38ND7dwPpKDrNhWR5G/v5142ynijiypNsUAqxXio9RQdlSqJZZRkQRRr0j
2ApeCxsP7qEnEFuR/nGChBZpk0CsjRxYuPBpuXldmx0bxS5f3PmZG6K9bCioucv2QMiSZO9pNj2z
r/HqkjsXNBzN7JjPfjwPsK6ALZEdKM45vQs7xwhYKdBBXKFTdCRwQNpFQuBaSyInSMuQT3fUnjRs
uhqz4XOH6lCPAWxaPHQCL9aWi1e6UnpRHRpYsyu4UgchAQA7DhoVaRvBT9JF8Ht3LBOFExQqsMMP
8rpjDFBiO9DPHdwedmkobO1vUaoQhufRcPE9UjN0PeZ5gPxvH+n5G10QDeF2jvBTyMs615mOpcTy
vAyBpCC6vD71vy3EidtVjuODYpLWfQYQ/NDyd+1vJd+w03o8/b+kle6Iibw+Dbb1xHfB0Baz2WjU
31P3ms8omRnHhCGfqh2ZtQShx1OZeywB9HGclGkrvb46n2hUTgalGk+ZrXZYbB0ZRmZoD4a43Xtg
r1kkQONlvZslT3j6TDmdZ3Z0V1llUFWuKvbjI+43p1pd0ss23SgAvbxs55ORBCYJ8N1xP6BV3K94
YpXvppuXIAAFDI9ytmg9DBTrlMt1bjJn0VvCVu4Tbnfo8lIaT1gOZ9k2F4XxJZkxJMSe/ztoqHQn
c9LC8WS5knipFgOslPyhGY4Gz1KfUJD/ivgBH+xI8RYzE1L2CvruFP+ivHs+hwcfX+L+BVZ/H2im
jrt64Ok7WoHpIQbh1j020abcz+Idh3Wf3WBj9x4nUMLD/6Lp6bs2WAkK7X9TUFjWmgLlwsREcYRM
QM+ixtLyypP7Y/MWW3X8X8Rlmknv4E0dD5S67oicheR4ipZ2APabpiglmDKqrTYOYGapBP0YG9ft
qZP4TA5jhNFjqNewvYRpv0rT/fzBlUZImjSoNs28ZV8StWydfcG8Fq3njIit6gZAySWZIa0oxqUs
UyUYwkg1LG9AFWLSDMtT61+6VhE4RCR90iqQJbBKfwu41mYgO4N0zPzRbq6wbVl0DXLRmDIvhOjT
o3Re9CaC57OCgWV73JpMKNfGIZYUDTN2+9S5WPr7gX5QVJsPyGV2F5NOXFqYe8Tq16YYvhvPXtKh
JdkGEPrq69EbQ0pmJVFDbL7l16EcapenvenoSN4fVlod8l2qQKqx1mx/JWXDMZSmMPd64rdceizG
Y6k97B5oHnOL9KH9HOmIMX9Nis2TGzvp4tUpfN9ZjBiESwycRY713ol8uSM+C9J3+/zvajH+qIeY
tRnA9M3edOqL+jEwv7+bFVgDcPDmt08hF2xJ5zOFF1gqrxxhnTu56Fbcg6i70tkQelMrmKbzrroJ
fJLe8FQDljID0yV9hZWQe4Y0mAAVkG+pSqCWKdy5ZMC4lu6HXkI9KQLNZAr8eVLT60mBwB7dlaGZ
qofa5trxD3PAInDeqiuOnwQdNjlt5daBXLRBwNd6dYEQ76M8S0DdVIogfeH/Z4AOWpHcI5Rd2WJd
hLx7uJLdb+oxT8nSGMLjQkzxS0kaEDox/r/WnKe4+QZhjBXb6kJnz3RHua3LkckWr1icTNrkrdiO
LisOF3sLrbUdcelNjAEhCYciJNqlSsirIGPRU+2srH2dLIwmQoklMl57wXBFKEjDG0E1nwm6tKdS
BDg/mudcIphM0M0nfZA0fIcXX937zdmS4rfIZZjyOg46/nk2xkB9Jm6nbkkxcgL0RF00aSYdzT3X
vtpVKDc9sMHzpRWgIv4bquBDq7bB5M6HLSM4k1DE5rquMg6M17cvr3/T34jF9iDL5eNEkFlhsCTr
8LqsmBBvOLAdN6kwdjrLKkzDK2o6UocWWUXxpNrhzaGyWgol7Z/Bl8WAa9zk8UuRlNXPVFevQb9A
6h62Tn7wdlU0n0BwCDnTecR8jVYmpYB6SzGqcFmBpwKmkX2BlhiuzTQ5u2IejiLtx1cCI+H34F8n
cdP/Ryh2VRBXfDv3sJQB0ngaRvjNw2vjiisXQkxTFo8YU/dULd5GfFORuKFj4A8pPPfpCCgJMydC
2tv/0QFIgqSLNpgNnbfCSOlXDvf5Fnnla9Fe6KWibs473moYe0H/Z6m0QoKtqc5VsSMFWiO9w7YQ
bDPF3LZYQ9HFrIj6HtV3hQXGjC8DneeAi0I9LHCfbaB3GhgZURXXZDT5HefUZoYguAFzVak6rB59
t3ewoUM+yeYJKy1/XsndzUyfHHhYPc9qzHQJLkaNGT70BHYFfwp0k1k0I2s66w+pRigI4O88k0dB
2MVtQeVRnOhLQRbQu9ELgOBYpHy5Ot9u2hF3cx8Lvv/c9vNHBdfBHay+c8KadzByi01qk0X6LvQ9
oLLUPMIojKUQsLS6nYUViH8ZAeSLZNvZuSmGRLwNkcgdZpHMR/K9/JxVtPcY9s4kjSCUjMtz9ouV
NonmFKPzkB1iHr7jY5VJ1gj6T0bdjrfd6cA+PAQ2BA6Q+SPnvSHHv8gDZQ7d6dEAgK0LhGpudNbX
upNLY60EV+CYmwXV862E44u+pYe8/QJ3u56MHAa9wiycFCBiQomYol8nVYUTC7cNka2sw/zy9Gv8
H3pkAymdkck6l7g7KnFoOHn7/fDpQBMC1BJXvy+OiH6Sf9Q9frKIS7bhqLhAwovdPTq4w7vKrdDi
zmkumcxt7SGAbKOc7hBNtpVZBMElgN/D5co748XwYFu5x2esKuBBTTwEbl4PO4WgscfBEFFB5rxj
aLkPfvnpNgbRKcmblh78VCpsKGGZgaP88IZs1b4nhbuaa5fhAfU4+0fL0yRubIiCpB9EmsmvE+Du
f55zyVLqp4ML+mulV0nyysQE1Pcd8B/Jt0GDA8WQhz9mvYZbhGpXxM2PUP/ahzfZyy/3hcM9V9D0
ZmlPmHi7cB7LXTIRTuAr4cA3mpIvXVRxs+6l8VcnGep4WFlfSDa94G+lfl0koICXjYFmjT9ucmpu
1oFxIfJW5Qaf+8uirg1IhD6l9PQ+SuG6rHuGKZsoLMvE5zb/givOWDxE6t7nc98A0IdnMFkAfyPc
PV/VgUPMd7ThpM94Y8op83/kqbsCXa4dCaOaimWIDGHggI8nHKxMIvgzRW8VqD2cOhJY05KiK8q8
F5mjqMqUIyRMCfSliWRVHGpG1mtfo9Dm12UVT0XNHYgdrAlTNnjdA22cC6sVNfK0s43vdf3CpiXp
rbI79ayzrQnYB4g1Fqs9UCEfenmYCaXZJTf3cg5ouL0W4wPt3NSPiyZDerWqQ6blpfSOuu9OMAdv
gfEHMHy6UjACslh5R/9VGLiexE8CQY9GoXq7YvTuJKpcr6U/QBR88TdV0CVKGiwlm/HpIWlQrYgm
BlKhCvTUJUJW9TN2Umo1XZvJoX3rsuSctwyICoG32MxAgV24Ap5XwOxXvKOEEJ4OlsLM0Io5ubP/
ITNEqhbIATA0MvFt6Ojti88WgDZ/C9DdBbf9yz4OC+Baeikybjho01MooRMnzYUMjhxbzL1VqZNI
uX8cblDfvR1GhlfMFfistscy7HQ8I0HmB8Ar2hnNW4buEeSRktWdiHYySJJICNDinIrnNLeUuexr
83yOresMfgLbCczHhHsRleHPMS5qJ+VJmdht+jkzgPfGb1O0ziWfgMxPMi3r60fQgU5dxF6XmuIe
foIKyOo9JI5ITUqza+4TflUXs56eA+GciWqHAWlfoltCcQs9r04i7D8rS/fVDxh/1mhgZt9zXdLs
a+veWeq56t+of6/12qQ+e3vs0GlJ41dTBI9a2Y69pfSn25WGnrnJocD9MNiglQcjwWyG8NyslyHX
5x4nYkYsUD8PywgY59qprkSmikEhm/lwMS3vcfvsEPhxI/O+En+VqaVKe19zegFSnvFlFpiYl2wb
4CETfyGLtHa3P0PnWsuq+3v6Zb3n1jYl+D0wEn9XJVLRV2XPztcdeIYUiEHP/+OVj1OGrvWdz3Nm
LEAHQEYxLpcGQgX5K9MKJZRV/2IVICW4DrWV6etCC5K8PUnAQJAdonUKLqPQ6XGG9L2RYHx2d/gV
ox51/EnqIWNeaRPNSoxhOE/FDtvz+nhhZT7JU9s+149EDuwLql/Pxf14P+b4QRLmJpP9oahdbOZR
gPRpKVjiQfwUChJ/0bq/TorfqTAb7XUp0pXSm2hfaX2YmTxAxQg7dwFAui7+Ty2CtSY0QVegr07y
cIUzYgwyW0CTZYNz5DQObWjGYtTAmNa5U5I9p27VeKcOVI5ABWAJkoHOpPaCeyNxfEmSunMQDUsF
6Wmo5afMsUYeaMYeKQngAILRDpx4U6UAFBlNhgcsHOt7piHiYynXiNpwl+X8tFSJ7FMeVM4ezwcw
SPi1hbnCbhTGnHIBCUGZBc85fiX4VfZOjqv7Qnmo/vDR+iHDAMwRMgRuHNELvLNyEQsmzQj64yFo
+IkAM7KuqTbq19B8aFSwJfHrm42zzGWwDEpvIcdM9hJGPxsLNtk3ix8P6svGcbWvYJdEzzF4PZCI
yJNq0I6bnetOD5nVILVWn74oIQklb7YQpFULGt5VW4JSqdII2Uvke1uc8txgMGrY7dhJe1X36S/n
p4NUQhrR6MO2UA0MHUz5zZuDnoyBmfurJrPepypdSRiDiO195z1kjNhnMRe9eR6Q8d/vCsKkMMQ3
BVARu0rSm4bGKQ3fkOoUDSl62OW+lX+yWsAYve0OQkypBOE/D3fKCdag2AN2LLvhr93N6cMFuxxr
xuHIEqz/caKsXu5ftnry5n0+T3AaKM+OxsN3tjmcrAlwTDjtfYwDkk/AwLUmwgOs2/ui/tcI7k0a
ZeWWq0Om528CgCHIGj0I/haIxICQEVCWtljaUE9Rhd0UIU0FcM9FVms0FUTBGvGrbk3i0RWjGC2F
OtaYw/vJ/D1Mss+M4i+pR6INs8rLzonoY2+Zrr8pa+HzQd6BwmOjmpwwy0MkpLLIVvRjjKrMoCgi
+Ab+ltpWMtFm9I6C3fhT92xVKMu1pMxjWco9BC4wSchy+dif+jlmOIR8fx/v7wQtsaS8HuM0SR+5
pb5m3eZE1nhucaBiPicrHUY9nm/Oewv95+2ZM8q3Q1E/fZ/WAMPWDb0J5tWGAqe4V7//IdxJjknx
6aRSz6RSuim7cwoH1l8RiBUqCVYe8UiWK8LPbRaIJgRnurp5moLIBlW3VhegIkZXbqiuU2bXVdpl
8vBAiyLJ28HJ+VpnCeKaYDzDKQnEewc6wowUjhxppOK9HJ9GdJ2rI46oJ471OfbM6OK1cJ4CPAtM
GsazhhWl85XF73+LPfasYP2VNWdh42E2dCNYNR8JN9JnP5fTHISj069COXmyqmCz8UHUxA3BDVWq
N8MSy7ZOB/oAh/mQGRRWDMbYMhhZeIrDUrrNQQ59jLcI5u5BLKhiRtRqFTIXBFenEU8lmSbdbrpG
NZDfKcfw0oaqKfI1Wga7rh6FWH0gFXyJdSAZF9/++hxL4EQuPeAaQi8zEXkV08KNKXIydcectM53
iFgJh9ZYubsX028zgPb75r/HnkptPYYOjmIApsKA6nB433wV/N76cmVRNFYZMq0U8Umr9WowIG2G
ndFcnMnACFek33aFnkYxDu8SLxiid5yN0Konxao85wfQdI74ihrCUbYc3VXgE6QPI08zUFhqK109
W+FWjiVte4Cwry0lUsbxAcxmfKorTW4jUcONVpBd0V6mN4+0Flw4PXYihIcFUTc/rBi4r5M35HLk
VewDXNOziFBQQRwoUj9AL0uqqEfc6zXDrpvAN5uXFymn7q3xxRNTAegVGiFiXZzNiJXXShlG5YcR
cFgLb3DjwuJhy4pj29wGHhRhSfjmG3gzq15ww4goNO1oKuJw1LRIosp59amgMn2uCyw8k4atTJRB
RODxJSfV02KeV6ij374yDC1YKtqK+GwLRGyZ20Pi84YDqO/FwPoMj0prfq9tRndjQdl/qNnk5jmM
Nl+Q08u9PkCnAjUtFCHhTNWO15S2DbCiVsyv+tjV1WEfgQWpu8fJ8ZnbFXPUpAgILMdwoAbgS5+k
wg9M1RI1bzH0WmB1BLvoZgR0sfq3pBEHZ8XQkC6rIM4Yf2JKsLUBIfMIXTTQRm/SpqAlC8ZxOxn2
YoxuFlieBCcummuxy7nMGGB9FcPp5D37KQeluxwA49MkdLBF5llQSTD9Gdl0MoDdrJYigaO2D9Oj
S/yS1cJURf/SO1t6wm8eeByM29qyJUet4muUqvrWPw3qo3i5fNpP4aOzBcRL/bTOCBTeMQYfajrK
fXBuyK0S2ymrP6RUOKVPt1WuX4R8LrCA+j38nyAVFNi/a5GutWWA3oInbdYwyiJiQqQLFdcID9OH
SezSnIyT+DTsugGUkoFSzmM6ikbvxjGmy20T/6IcjvExnGNLUCwzZaPMK7wKSp0J7oSrW9UUqexS
QsXLuI7cD1HUlAwDay+tM8w1BQs4azvR2wE0HkHfbegv8ZaxQCxszaZI0qB/TQfv6lwJGmf3Bt6z
SfoTpWMoEkB/NnzjNFT9nguU4WGPfAH56a5MSCk8gWuUcIVaLvfG6myK8iVRnr9x/JSGZnuajHZr
M/AAohnU5maaKHWvC+HtDIMe695+bnda5WN4JoANOiGH9I4R+I5Tn2R4TqeRHC/K73Mfj3fixefM
dmFpN1aHEa53e0Wzlgv1ifbe/ezWzOWDdaocS3iZpnERSEfQWIk2/NljDmcd5QwQpQCAT4gupqII
8zn4GG3wkQPE3diXFqJ1znglqZRlZw1J5U8EM+vnTikgjtdspfu4MtFVtzDOx9XQ6wm0OYWF0YpR
Umg6GnOSQNwQfHYIfLby1AzMRiBib5+FudhJbtLkhuykCr31LVBsejWQzoSYZjHK/ioZiNr9gDaw
aBriKmBXNbN+BvLmPd5iLET016sgmQsLw25ags5qHf6IUkQanVNeNMAKfmJQHcwIXw/jIVV0Y7nd
ZC81WlNm4+SnmzZai1ywhDaWD5zPKXs/RRXxzZ0zhzE6maxvlB2yVkfk5OD2p9sTyDDn1mNXhqKY
XS5h++TBTULTW1TlUspVim94EquSCPd34035bmaydFQpjFqnZZTqA4TdmjFuIMNsOnbfKJQLRUrc
rqinEGVnbkxBczfRXL4wewuKXHOwT8mNskezRdQry2tpdPbBinLSKB5tLgOIS5SpdOMOuyosMmal
1NjqWg2zYvrXilYENJq981BYX9g9wqHR8d2x9wgMH82/kRB2W8GSgF+EPd90X/NQdfVaxlsL4U6x
qTGNjz/+4vUw/31gHWOu7V0E6dHfT2zLNvW/5gYP9nHwackl+6hJeh3Diqn4qXJe4X8kQEdO7xiQ
o+XWEmADlBfeWRJoW2kBHxq5hgNgKiUL+Ko1FvfClA6INzOwJJBrjw/2soesAD1K21l3dv3hMgtC
P11KKv/blAfIKH/kTcdoilAYB/xATcwJZwuOYzc298VRMvC9mcjOHP4lb7l5Og0sRPaZ1BQCJpPj
G2gvlMEa0VMhEqMhcK7ccfOXg38kfUsDWwshZKwY/RanPpwEqVbGNuvAC+y/2FG8qzdlyQVEX/Al
0ri29tVo3I9aS4UvUU/U/qzEdBXyDcpDzE3w4TiNNBkmIfvZtJddNGos3iX+nAte7ff2etij8WgS
jz7QhvEqP74oGEem1tVp8VAD8ddkPS4UVKAkJFINW4HsjJgfvfdqUpWOYrwSI0gCdG2Zj9wSqIwp
HzFxbEtMuj17irUPxltTkoNNjw/kcIX3570WMCVD9vwGqiaGKDblQk59weXEfgZlAwwNIcMcz18W
8aJ1yPPARDyqZC+MkhKvpfHTlYPWZMOEwzFIBvSn7vAl/zLW7GYWJNcrAClJcAFJ7FghiXg7xg3N
rJXa5PC4P/UCfdSxiuo5BAtUz39eZDDYc/wFGvoUUdOoUrn1EIsnrMcx/txvlQ9wP6/RzlcKosEC
247wiAbUCLHAPyEHNyhvrqc1QAuBV1cka4TRV0Q+zdi68roBU1YgqOGfCz73lKC4rfZtpc6uUpDy
i1pZFJozOYrnja4QJLAQtqdZmjwqIUB0NdMCqtgwoKCrx54vFQpXW4lch+WfR5Xx3LrEDsIA8no3
yhaXIqtlpe7+yY9RHvEk6JznLwhEcSJk9h+XuhbWjI2NqrgfJz7E45PxjkLrdGrTiQid+1fcga/c
DAeGVZ8bvruIXm9zNfOEJHh0PjLYWB42LZbzaBXQvyWlY7okawyAJkA1iUg8vXABsbrD2qbMymY8
eIPPwl2IGF/MkhT3rg4E4XZ8cApseXPH8pNhrCzjbjbgdWy7MV2/bk8UjBwQq1MizxbkWv04eJXJ
3DGs05V4kykpbe5i6UB7fd6cvlqSlY+48Bvb8a6zOzcdU6WJlwWyW1Yqrm8NyamejuBHm2CvgW42
7qTjaK1Dcpui2ZN67jHqYLyUcWntt4oa1765vwfP6Q28O8wI/JYOqr/GHHqUCvqnxijAUxmD5tNB
k/3eXYwnvTVOvkNlo5UheSR7y8HmD0E8NhUItvzkROxpiP23cbjR3PysZcaW9T2kIKZOT97Z8jt2
00AOTZI7mn0OYCy5KmxI0xr0gzBAOzODTrFss29GRwkZRL52CEKwcmPrMIvsiXBCXmEaoyAIHrUJ
MDqKwCtmkg+nlE5QijRp+Zl+q8Ck6h/6HI2x1X8MGRgMjW/K1qZoN1nSuZxqRhxkjprJlmnBpT4F
C8A9LXEo1BbZPpuVZ61JJvpXtsjfVkfa8ykxOvzA3LcJ8l70I+TGUa1HvMcn7FvGaeTjFWaomAqa
xhN0c+/EA2nLiMnP16/i6sIYebrkDJskc0x+YyRLjkOjDr36k+QCZ3IyfgRxM0/CtvYoVlLun90v
DLyZwpKlNbfbjb+1DOJ/D55EA16cnwLQxuyx83YU50NrAZ2RfzGJd4xgTIP2DdPfUrvczY2N6PUG
m+UK/MXo+JXphP7DGsm59X2lRQBARLZ3hVc3F6MWXlajLKmp7AX9ZaRexmwkUvOzQZxdfM1eVeB+
BqBIb/7vU7C+D7DDb2CYE6MV0HDi6m0yfB3IaRL5aVkj3uggpyQX2NMoDpDqibeZZATIHQAMFX/p
/OeKOG9rAq/Fd5KEXdoiFOguvbSN3vD0CLMvhagNdrmNZbqFLBzoRQYxYeQqeHvb2ezX2xKjswxW
a0FjNYi9D3sm1V28xfSb1aLU5+jzcpCt/DhU/Te1lHlStxcriGJF1AmQWFG1y/qSsl7CwhUimsWC
BL/QCdSpFvHAmnRcnGw9RoLwPlTOi6V+mJXH0fJvNbRq39PYLT+YdiaKQxpiYUQGQ05JPof7u0Cl
EnA7u9lY+WkfHpmFl6YicwSqYhQyQtfzxc4ujpk+JU0hT+HyYQSFamvOTvODVkhkvYAzpzCsFNRS
D9NL27wW3h3Z2XCZPp1xQnTBjrsC6ojzpNRfBRd2k7OdTdyjbJuCGN3Vv+8fMZqDC2kkSoPTQhuq
NFsOXG9KU8owjdPweoc+UAy7XDA0OM13AoAgF1HgsvF3IvsYVjDpDEoU+jTllUuv3OyPvmxcDTGD
HckgCZWHAGY+VBse9F3NpqQrl5/ggq9Ae5JYiH0nKFk+9SMJfEpTM/vXxF+7/03JavJo2RLlLhrV
/o3lTz8VDTCyCXFwQ3WwlDA2AT0Qr9AShB3QIYDlQMUCl4M0JeBBtRA/SktWsVFZPlqs8AqmRCBF
Sq5Go/NuXiitGZCrqYe8eSJ1EIon9MGBsHh6oqljIppSsRtj5iJgY9hs/2r8Z147OyKi6xqET/Of
eY1Eg9IUpCTM7Maas8OU6ecdFQMCanjwRl3dOEQZpvrKLe57A2K52CUbaVZNu9wG5UblDBoKS0xS
qffjqxUgZvUzFZ47zSpXsWPNGjyEbxZqvfsLWRs6DoH7Zjaem/w4VQVYsZ/orMc1oXVjDyj98Dhx
R6W/bhvDL0zXhvBa00fiZpnelpswwO+E6Oal0fD5YY63F4HfNC42+fmrHatVsN/6Ix2KoX66n+B0
Ig07+FMxp2a+f8HrW9a/BnXhd2stvE4faw7eS3smyawyslxHXyOL2VZJLSidM2aD49bDcLegx0KK
PHc9wIVXg/XsuDzq6F8izFJ0CzDBbTyWB+jXMblQEnVhZHo056HgFGj8xrMe0W+6OgR0qTUUPfsB
kxIfnZRO2ZZJo0OB2rVFB+FORKz5vQ6hMV0BXcD+DhsO9ZMgAq4Y4n6+50y/M61aEneHxQAjCqmc
38tqjv1XEVfhpGODwI0kFlt/JhCp7cKV9+Y6YvVKf3ptc5IWBc8adODPNbaIi1BVf8BFH8sYYSDh
+hAIOSYJ7jzIiq+0FPR85tpyNuH70C1WYNS1Aa9B+ZpOjLMN+fvTOjY52RVA6N6MGmLLx3OtVtoh
WYSk3DYfm3MkHWvZLsMFe4s0f8tsjZTgLFg0RqTYB/oapzjgbzMiZRPWVuD4GC7yd194r4tFd3ZM
6tnW3M08JrUOWF9STvokgdH1A2+j6ldFSoaR2GJbGUel7ULUwg7rnEToDXElYJmUuX31sKPcx6NS
8XtsV9ZroVkweRl3x5MtgJ4VdCQZxogPH9vS1dx71YQxtMerHjx8XxQbJRJKtaBCG0IkjTXZ4Kro
dM7B595iYGjZjX+vOxPfJxqtTaWl0HYM/edwWpowyp8DmHvdflD77eALGT5AlwgUBca+nnA1/2OM
SJXGzjD9pUO2HB8gehDOhV7C60QcTbGCJVO5EcAk5SC+L8ZuOWqvkFnQdYnhB7JRICfWecCyGU4P
qrGyplVdfazzMl067rb8/wOJqUeZEZDnP7hv+nMgiqYgeWdiucQIRjgoyLXlfoPmDyl+k88fz5mn
7YArzxjSJKM+r70HQhVNdN4nMZcf3hzLrjwe3DaNYq9f9pbmepbi9SO6bajvkBhqTkrfH8V9Tz5v
IUtIHHkOA472fOCLWZc0sEbtli6p7HLzQbWn99ORb8BfeW6gIJCS4QLejdvDxom7CL8u9slWedS7
uqM+enXHUmAc545fCJ0Lbn4OXRywOlcOj/D0AisVxDY3U3Q5tVr3MBGeNdd7CRxUYMTTUGdTa5aH
2t/cj0SpwiIAHAdcUTy8IStpm1+dsKg1u9XgIQYJZhaVKO0iCpNp3AycAesHgwtY9ZmbS5rZcy4m
H9g5WlvyUfCny8lW7a5tX105DM43mG34sylirP6y+q4et6jQkNWf9FT510VDh9IDdqNuKs2EntmQ
KzKFqKdFvp2ZbJxXCY+8aZ38F3IBmV3Eo0OMGcEsdIKpS9TdzSQN66ctNS/Kg0yKyVaNsZkxTW29
piazcbIymTyWct3TAnauGCOHpraMgFS9x1iQZHkaYZChqzpRsG1mJ3K/TmcTOOKFubfBTftjjyXh
Cck2w7yn4m44N9bhfWeTiBEXL9Mmljh/tH4El2G9tWML91OSgHJ60ItQl8ZwOTWYgm/7stXwFF4j
TUFwresMQo/MwtYrpV2e7eGZ9AW2I0oYWfkziCpMh17xEyjdirvBl1wRdFNQlhvCIm7PEP8EoZjv
6pPZdOdHtkx9UvyWH+3leB6hZr72DZyerDcu4dRcN3F3phgq81snqwBNeqq1NEESfZkBnr8n7Tp0
Ku3+Oq1FRZ8wTuXyl0swLnsCyPwEpMl5v+4YSHNQb4Pq5O6tx96uQhs7SIhSKeQQp5cbmlo7l6vA
ofXBUP0Os6l2cTIdJ5hmoEELbY0f5aR2Y/o0HrFAvc1tJxI/wrb164rO0hI1Qeh3vl6txDpaamta
vYhLi4P6KYmXmBW/zUY1l9VIkUs+wJf2i0wRpVB34dyPXo47tFukCoNyN4ffvG/KdZ5zmlg9wd5a
5E3wvCzsVLbfg40flUe/ZonNKFXECF0sFCNKVfmORs7p2Q7aJEze0YaHvAOAb04UE4vgFS66/AUU
YyRbGbDwWKyzIpXf+SwzyQoTc1xRuButbUBoEWYGUDoCh2r78TMt1OkLsbVt2+r9n0h2zXDLyPXx
pPr+0irXnK09TKkbQR2/X1UGqjeCrxoldEyuQgnsIw0uRsG3pRY4oKujjJeZhRduLPPEFtsVW/GU
0oxOjUX6ZTNGiZABzdpfSa9497HkqPiGd6J7ULRm7qYl+tVzK9LNSHS+FwNH81GJW8Po8lsTitjT
1g6+nfUDVXDJQLpwDYuGpoS0XouxO42TpDugR/YO02qnE5yVQw5hW2qCdcCkQ29YnQDEq8doprYY
5gHgE2xapsYssxBJ3O0rQhwwjp/RGH3be0/LJ2nTb37ROLRBI9fGR/tFKoBdqXxN1vIlQOHdMp7m
kgmFXzBH5pF/FeJg1frfCVmwEVwhHm8hkX04URLXy4juu29JgIYuEMGLHCuVzHSbjV6lveNUchnE
7z2NUvYrjlg+x6uImH86IgYan3GXKwrGgSojFB5F3BSqKLnUMSgcbcFDnhNx0HVdfLhIW+ntvObL
i0vnA0KS/eGyR+d1kVQ2gWORcmhSE+/zYQ5rcSrg/t4ftl6C+/LK80viqeUPfXBvGEorr66dDO5l
B3Aftqs5I2h++obp3uPQTPeF8oAIisr3a5mIt9ao3XoBCuGQBSbpuVxDUErcOXcL/jLm23MUKqQy
1OGWSBVMxRQBQw0TVBXTBQX8KQP5W7Rf73DONGU9fiT5OXinnBmzOnv9WJE0ktiSEag3APS83qi3
LtYqQKXekdKHxrDGlO+RnjU1XBD2RhhTwJ/CYh9ghUjaZSWxNAmZtrKG4FX+S+XgoVPOJzooEo5j
+dp1MhOeL/ysUKwHA4M8f+cwvRhUqBiIm+Z2Imipm5AdMqoXpmqrf6UXK977O8w3OGrd0msrlCWV
bIzorP72D+RGRHMy7Gi3mpp7s6zZFKyLTA1oroNyKYVlxkxQZjX8OR3QO+LPMb0oCuDVFCIevWrF
kDw1R1HZyWA2YgwLXlj02Z4ZVF/Gt4jPt9vOVSHFQ4hwuzx4cz4TT+CGwnOMw2OlMA6K1dK9Z670
5pdZif5CDX5cvOcM7rNtE9RHncsOMyT/VtYkFhyhpFePT3b43DzDZ6/i4kpBH8ylVHky4//lGmRW
2WBC+becPiZSaRJaZCAEqsnntk+nA9qmujXwInjcRAvQ2oG8EMTHEqfi2QifEliVNs1+FvXHElno
kKDofxJAjvF/uz2UpSw3P1Pg1rzOJlqObs+EFf5uYNyH6jGfPHvH0hxjLblD24epK4BLaOCzRMd1
ZgWGIUQ/IibnlZTqnaDpsGmze3YK1LNHjnE5OaTBbmUkQKhN4G2zv6TtEKxmwT64YNeZ8s+sYlzp
45k+j7eJExT3YKT2azZKoi/Th0uoxwUJEvIO916sX5GmiZAsf9gzgBMJuXC8ne5i544aQANNG0ml
Z8m52xz8urIOtqg6FYkzasT0QLhl++b7QlbyUEt2XUZXgVcgeQGugxny6UVPPsljxsA6iJNp1u35
6R4wljZ6jJHdXmIFpjFfI3jFhmjxc4wFZEvVV+xMt4LkE8eAf5BjgCB6iRiOLRURrOitAcMSYjxS
sEL2wrNCu/u47yEBQryFYTi0EPjyUnMRRiKRslviJzDJ6wiUmojzmPzVgDQdVNzSFhKyyxAQnANe
rHI9tHauMHP0yTVhiZAjpxsuKGTv4getoCKwwO96klA3ZDUXT5CbgXddw3TGXAtg3RbkOXoKPx2g
jXP4FJQ+bkbsCNgNNZDdmA56XIqUGDLVm6z/Sa3PLaINGARQWUeSwHGdfdQ+I7qQGJV2kapzKkz/
OFTDWQ+hWhbGSFiGw3F2dvW8H7zi+bcsWwKB1GRQFIZebdLxGxPNkIUCUlBaZZIFo+tHhv8V/ynE
1HZkDIvbSGwEIEx/LMwGbYCZhvOdAC4h2ch/I4S1IZSiu5giMiWBLq6mEH7/18ir4eoHU5S0RXUq
CoQYwU839jigf9gLWQ2RsqMmFGwVMMgPm2c+tfOsDsKtLdMR8WS65dKEf/hJN24HfvB+xu5quyXr
jNvw9KOtnkpds8vpcIJXJlm4AUJu0ZGziXH2sk4lLqVQh1FgWBB33bzXfSb3ILglfQMXyDahyLYa
xbqNAHbop/NZK528wLv3XMnhMDaoDosMoMzDT5HsjTLXvYOidxM0C14GDBUieSDoIJ8ZFeVtH4E/
cukNdxn0ocbfoAWSo7kAIPdB0SXuL2ID0T1rHGGhhxZQ9N4i17w7hLAFVVbVZTSeyCEI4eulqtKE
K7DrJRm2sYWXHe85YnxdDiWpd/QqDi3DXzuGMzqjsrdsxj/kocYNmBZLixutbKcy3WeVUBtRChgc
kU13Baxg8WG02XOvvRiZHX2dkAL2p+5pL08HkYP1OleYv1wUhwYRVYWuadNQJPrYaQ/Ot1U/aT5/
vF/ZtlPmkVlokieL6uIbjxFGscVhDqQ/piogles6C3N3pFKIC3fgeOVd44EsnSJV9EZvpgUOOVVJ
KdoRcKBzFER6D/FRFyox5eiTzKYy6i+wBFmovJK6vTcOWEErFCOx0ds74nRO2w2tHI0XINvJoLUM
lW0dPkxhxyzQ5oOKuM5j9kudkWDB75ufDQt879APRJkSXk9vKveEBVqybXvyPi/QaWIaCQPQvhrH
eHD+hkKO6PA0+Nqhq5bS54z8MgdlS8L+vHnBZtgB/JXZXped5YWwAwhu/cSPkQ13zf9ZA81EJpx2
+n4NTz/UH7GQfVqll+PMYlT5epB7mJ4InQJqLmsaZFmZMVQF0e+mhcxKWIYQs+cyyoVok+WSId2n
ZsC1CFgEiAQnTIPQ9LnUSyl86JUEOxMKs89/3yxm57JFq/pil/1s0yXusZMZBT82qyKr5aNd+UZi
6Zg5fDV76OAVdljzgax7+tt73UYjyMpu3XaG9Df9Uxj/s1pRd61AhxrcGwklkkLsH9sttsPULOJG
hE+Hge/tUb6mGRewS2hRB8eRyMwnp0G+Nn1LEC7ZI2bUMNvgKSzx5A9R7fWkTUYT8hrENHhw3KLT
TV1aENcWSZNr1XqH5cVvFdVrBnUzORruqMx8oC+Z/GPaCVKQKDwF2EyEk4eDXPG/U3XUYqLKZ1eT
kgQpVPmBYVvCrU1cf941m/e+AJjWZtI033H5/9eQXU8dFJAT1Orai0I0mxxkAUC9UUpPQW+ZgLyM
IeVOKvaCJwi/O6dtnjbtOcuikuZcJKAqiq4yVNrsL3LKoyZx/8lLRnnr8bH+SAGOiGYXl/LPmnDy
I1BBwiRxpm0G26XzIRAfMy+dFPDgs8XpwsB7vHrxkhickYEmBL2YK1rAbeU6kjYDk2RbcsI/fnBa
w32GZNxNK19iUZsbPDAS7oiYiCGCbHm68/StRQr0i+mcPwcmrs2J387FleBh7wUNt9SXezmYpI62
MkzPLrMDdxCJmdk2+ysj6HQPgZLQpi3qa3IM66/EW2lnkkgsexmjEyDf+CkUC6MoN1E+lGjTz2KT
rFXHvhDdQjLlvWCSYBB0XwJuvl53xsljABbNcCHzyB3eOppA5g8+ThjLmMBq8SQAIeCguAFB4beQ
RW81I+eoR7+vBxlwSgo3zVqvmQLx/io8bchMh6YTIMiD+KuPeHPa9TbDXBEnp1/XLNfNsVar+Zw0
qDBY3I5Na/zYgPVRYtLsEg0FFOKnXxVN2V/+w925c0AMBLa8x8xAE/1epbeMOwyeiD63sfFrB/J/
WjrhxavbNX6jCuKgP92gZm6xf1Ygy7XCkBkR0xZkzEg605LJ5WRtYUTCXfv2ikl29aHXZjsn/9du
OUy4MpNt6yuuTq5ywL7sS+DtnPWkBzrO6FWlsxK4tqSbrEqnF0OhraYN2jgRjXHfXlWBekTR7RtX
u6PtB4C9+P+AcoQyXm2XbSbEKf1P1h1fNQSwYV5HSRibXAkjPpbiv4RnNp1jGamwyQYbhory49/+
P5TjmU7u0A2tCYmJ98zITkelJPkV1PHNqv6Q+6UtQzOM9v/TWmMxiw9F9JZOd4Dch4gAvtKBwsyV
O04lLjn9LaAsftXdPtIc61tmEIvpECm+uBnP//E3FMCLkSP6h8ibHFfsXETfUL5Z1Qbg5c7Fm0dI
DXxzc5SBYjZbmZ8zwMUNBIhpFVsQ2cqdqvyJ6hjBab99AyZNKBDNMgHbbocidDOfiKBPg28wQzu9
NQGL7IM0hK/yjt0xG4Olt/zkcnJLLp8wtROomTAGjMBqY7YP+Jm00XWjDSztRL/5ZCYGmiQfDgns
oATQtvbaQuhW70fmwhQymrUnCzs+5oIFTiUrBqZD3UIpbUWalExqqsawWh4cORDnoKocCaCSHSy3
8X5pttT0OmZjk2ptheodl43kniH88yMCslR7Q53PYnKo7EMd6uMEAAi7tYRGYe8lGqA6APiDiexu
K+VWJPXtwWWSIyK0KfwWCoYLIgWdFNW772pAO4w7t2TEZ/1MP7p1bhiLhZs0PL27GRlUx8wDYBbE
NwJZdXtwveq2eX8hI4/CSzvntBk1de8qj3MehLbrI/YKaX6n/KHgUgwxWSYC+zY4YSjswbyskqYN
yVmBh9+KsuYMZ8+8hAPMD9QtS1xBIe6+g/yXn6QAvlQ0b8B+lBuY9dHMT8pUzV2EbR15zsMwdarj
adupkJyW42YdIx3lyv6F96232OWZbEnaGBSbvucwz+YXtqHN3l0Y7zpvJMGocbCdHaL7+2Ut+8Pm
yCPTdhoNKGV6AAlulGImLT7n5/N7CRdW+4tWPj6XzRfgRlhk5aQVJePkynd7K2OSvuadqh1Nkg9f
ZgDoqO/ya2OTfPhxl3FzUoLDUHAvooLIXcXNHS5hrn+DdQyENL35JO4g3D3RCFLiZk1aCSkNUG+9
JfBnope6/rBEJhLIJJdumludnnM4fSy3Sk3m8pmSkXgtwe9GqmNxo3HDykWzNg/pP+hQsz8K09we
6OsfIYMmfsUeR93rSzAcLr4hUjq4n1xt4UVnUALYYMqlJXuMVpujX+IFykairh5eJHf/VaxPEoVE
0WIyq7Wm/cYHqjM3BA5MElD2IjprEqqnTcECgIRk/X+fNE3SWw83g4hZaUPNkszHJzItwPAvPIIg
FKa5RF5uxQfzsbfWnPifpyBxIY2UVf1eNpSsHAaFkh70ATdhKxJT3+Y+34MSwGWuob3BAfND6zYD
zM7W2OI2AqK2nIyMlsGrVBl1I8nBNirKVCI4wMyE9sMuiBChCoBPRuZX1n6amwHgTmvLbXzJzd+V
LokRe5afDdxT6rx9Ab3GpWlm/W00qlsjOYKDU6phPIvVWt6GwN2O9gad3mNdR3qBoxzRwUJ3r11L
V5hpkypdziI4by6sFisXhFOzKLU4yLZEXTElfCz/2ngqiH+JjucIjbTxKf16PQz9nvE0LeeTAuYa
T1UJwfFL734oo2rCMvsjydNxNpPXK/HPwkk55KLlveK1SpNgW7NrLrHyd0yTKK9Y6OH340OPme5E
D1IbA4ZUw2BIuGe/EvkV0+h7Z4KMXdmKDxb7wnPnGEq0lPE98yUS+h0t6OI8SCyVtv+PTXyYzqXr
VR7yO1lHxNRGNyMYo4P7YFZiajkhkGhT3UdF04fTmt/PwdLl6r6r3AEmOPm7AtH3zTN1clsu0BiL
HU2W/a/0bg23YI+C19XmORHhLW+FkYfY2PuHx28pFiTILqVE3djbClwv56haDzvfYd8koAxL0EN3
Bos/nPUSrRYOzNgRfBHuKN1XwYJyiitZ/z01tsRu/3fQIAMjAvxmlP0f4/ft+xHOznOwH1EGXZE3
6Ia/8ij23XFYWDJLN+BwpTYt6CQGR6HtttavWWfr58LQUU7P/0/ahygMI5iJOlbi5T/OZ4Fnur45
E5mmqppfzrjYOuOF85P+BVaO04jMZeTuBqB4aCl9KkTp2XZhJ2aag9SlifMtPEVcasR5xGJhgHeA
mww8+xOd1P/0M8lwrfTTjoIsVrmAm+dlBeTkaXKm7jAs5hAFHF0Y9nFFXXO9cTLhYJDw00rSHX8N
khTe1Er1twM7Kj2oYXOxPGd8eYwqohWYR0ae8mQkuwoSpmndRaIpSI8Qb7ihimfWnF0DYQsv3Za2
AO0U3JxFClMSJJFWkPruUYZkLXFW5SBa2dQIGkIzeViBDLQKz/Juhkto9xN306UtzwndD69pSs8H
QR2gY0nd6Ncp4IG/gvACfMph62Wco3oaTFcfXtzVNvcJyuaMgx0ktdcxeo+30EreUMcbvrUxbBof
V3GSPUd08VJkO/palpJAXfBnRSnw8uk4W9TbSXj9dAKY7xuFsYxl10yfSsCksFrlEyymbwLweebW
FiBzPH8js9BkibravZ3nwc+6TLRYdu/PHKDx2rZhaobFcpWbkNwV+oWiz38tNM/LiAVQ+3wWCkHw
qgFqcqJOO2Gk6hMTc2ElPrQjWVEQMyD/GC2507NMGxQ/KciaGETKZNIdS5QP4hs+0yd4PZLjWMxV
X8xdqtlLTOnwoB2BMieUYO5FUVva+RlEpKrdSBP196VySD+92q3dcVeeAfmGFQvc6LS1hXDXRhEQ
JhVp1OysRaUPTWINH6gv62t2zEXXPiY+YNQZk7BlaIC7Zur5yIkVY6YPIA5gh5kp5CZjNatF88oP
kzrB00M6aPwEImCtqGMpMcTzRBP1wr/ngc1l5HED/+xy/Fwo75HoZsDfL1j6UnhU/K8KYPHCECqt
XC4k7lxY5QrSvhtGIaqD0UdetZzEOx6IsFiDCTRBdRIrHyQa7U3w1W97Y0CeV4pSsbU4nbHb/GbU
0ZbS0JAGkRBbANQn8sFDRX+KpLn21euyCGY18ePbSTK2zJwIlq2yqgFwd1lmiU3WKXviD/2sF1Ge
fy+XZ2B90LiXaSTtEsITsXZ3CRBAOq/zfojYTH4b+zHxbcQWRqA22C4djqwn+RDdu53bVb7bDQl3
Eu5QlR3nvP9YtNuyh2O6nKhtDT39jAmw8Oh9qnPq+2kE7Uqcp4oNc1YvcSlaMXDCVB7o8DgZ3fSn
518BXk0A6DuyLhBXABMv+SBdnBb+H8w0YgmFI0viVJyCn0pjcaM5JprLE3FYuQ75zwHoNG5EQ53X
ro2Au3RNs2QvGmr1wiNjxMZPl98rZWtRQFX+Y9pYYYv8n0R8qlMqbVJ9fDUVIZlM3nDGuKP392uh
9Ip/cpmJTAGWFQGcyLBADi6X5fx3tR7hwYAjofxvUyjNsOLAE2gCYYqQPYhNycFGyzm1/t6qyUpN
0p9Fkph6CzUyw/qK/e93ZGwQtyq7PajDyJEeTNiwedgF3ceWGAH74tJ4TJdGEMcNZf0da+BHRI7a
z5Lp/opHBzUdZieFH1Ck0eHSJhj8obFwCPQnWyRolA4pfUY3FcIl/GlspGaZpKgAxsj8wBWSPcTO
6W/FG1BNMbI8NkbztGIGj+MHc4SSlfPCPh++SZBakOHlWQh2rnYUIux8do9mo/Z61SSi+ynFHwSM
6iFcVmy+TBA4VdMEn5pXwX+JBcHEllZxpt1h0IMPmjEhrChJp1qZRxeBAUrpKJ6F+YtH1bFOIos4
kuMbk5wlWpCIo+eh/9ZF8MqpfaK8S2SltvktP5jMPbN7+ijKXItlM8THjLNSkZytzksiLSgjdntd
V3ITKryFosrcyC6YKeJ3BiBPbovsVtdC2xCxpURYG/BjLfPXVzyEHeKIXZe+Bv0u5104KgovcNgG
oczUJ9cOrHbsLK5j7A2aVcRTvsZ9ZOM5B4lXgUmfvcfMOTCEcBxU/yFST8pCXFgeONIWJjmeIeHG
3oyEF4oL1XqOHgm7pw/FKBb1/jiWOo7HsVTNREYpQ8bVXdOpRUl8X3nwmkcI3wSCpIRTbCZ9L645
Olsw2Wfwl1YzonMHPNP6B/2+hhCdb+UvmOcJkNmAwTCV2jWyX5jmIyeoWn483DawulBibwC2Mq5Q
akzXUM07W7CGA9jW9//laO80/H8AjbTe8RVkMY/Y/QDJfqUV+YHXyh/JI/6HDQ5bLdHWOLu5GD+T
dIxbipAnGgP6dfvgZodnjRTpEmet7DO8+3wJ25zjBKOEIfP1ZAu6l+3XSR64IAxQIFSfmsUtnId3
TTociITdTXAbQEkBcC+si+mxDx6nZ4qc3S+bzZiX6T5Xfs1Cp9Ri5G+q8jPsBKNA93A6K8Esl3wh
MmDf7/Oy7nyRANW27EtYyjsnmpa0jDGwcoq71HACbkwreZSQ6Kt8RUR6wwpqO8y1wuTba02m5GuC
5zcm6JCiY3EdBfkA5Cf+zP7VQfImr9eD72hmOTujoTBX1rLcxINUjgIAZ/pBM3bPWK+8p/hyWUXn
/nOhBV9CR/e4nNHBgdob5eNRy+GcXs7aW673/5Bzi/4ZKanunKjhmsnUyzQ3AF2OwHQ4ium22GFB
+MzV43oi5YJA3VW5mTEDdmJ1/2HfL0ST2f5ztTO/VxhJD3YfWCV9FMZkKbWJNXRhoLys7gecn9bp
9simoMQWuFOYvtrh8y9IuOKmWWDYDEmsX7xkvZcFeWc++SlCjNsvyZSrkuY3z0a/J1fXBQ6nVNbh
lDlsj2Bwv77ICMiBwQbY9h3rQeMX7/6viUDaSsv/ZIzyYZnZHAPZI8BmXteXOzF/GIEqnEBFPbQ2
ddmLBE/1zVKaAiCCAV6vNFuP+0sAG9AL2O85pYGZEOLjIeCvsJ9voGvzonGYySCGsMSnQdtWPC2l
D0BkHPpQwutLOpTX7rpYo0Hv9mE+IYajJo8HzTI56SrtevuzQ/sNpDzjjl06XW7BPxMhM5Ar5t39
U0wUItCX9tULAnZqhZ0L2KSjpnDGmzY9Is3i0FJPnvSSAU+zvdpNOqzlwYuKTI7h5EgBDVsAgv17
VqS9csu04GalNWKVcJ/IgJq3kqmZKYvuWd/JGwXyc9qXD9vW4mt4saDzSFY0NrXEJNOmWt9n4ibC
mbYKvHu6cXj+WUwzg/WH0kUMouETe2Z5TttMK15wlH5dyIKKs0j6jSohdmzpkEjU9ngFbzgK8CQX
XOh+vf7MUMSjQSGx15J4FSGaUYRYvt2Tzy7eD8D05RiK9eZPE6JLN8m7iG+zTtMESI5Bs7vuuqNY
2FPlv0D8DPo6JrvxSlQ+c2qduT0RcS6lb69rfNzUAEm3+hwkErm0MzoTgP3soF6tDH1qYxZYAauf
KuLKtWd8Y5SXUBM4JlnJx6D5cts2sarOOsuOHyjMDrsn/T+pMFi0/mVx2lB/dapJ41kaZOKQRsUf
mGKu6w27XAufPMnI7ByMDR9nMHCIGAPaH6zfzH/GhPpT25qAaAh+taXSpcXgGbgeoySM4FV/hc6l
pKXbyZrACw0OjZPzJa1PI0rcE+yJm6pDpwjQywHKzgFOcv2nZj6CfMVG+K+Nd+TSRUcAsDq9eHs+
AA3NWegbXHamJYCLkDDGtY5EdVXWDjh/HX2R87lhoJCeAS7Nvume/+p/nc6aVphCi4RulgyFG8bv
qwJQoOIIALJAgANxmdfULPHzxxalC2k/hm/Wd/Typ7hUvxPI55/7PZRQBt10c9ASmq+kQqpH85j8
4+xR3V0k60rsieuJsnqUis9kJ8fHTv1Yc/8avPyw92i+bhztooxXelYsNX9lG0tKuYt5erG8XTMG
t1T1SgtXw4ymslZ2esDn+nUoLyQer1JEeN/bt7ic6ZhxvgkX7uPqh/yJ0AtdgU36EepVn2vp5f8j
gM29NhWkMrP3uszRisV/+8oHf1/lJ1kKTUCSuqUoyVHMopNrraKuO3yWv3aOwmjwzyH507DuIQVw
yQLBKg4otuFNl4RjIcR0zPszPSnZBexSPZzIZhqY+fgVk2tZUpYsJOUW3rjsvqDtA0eFS6Qqk1vL
1bQsczqfNn8of3wYX8SAwzU28HQ1ZinvBeZBmkKe2zq/PeCjH2P2Z/sqQEt6eAyI9lEXlMMOAm1k
4X2Heo9g1gsj4Na3qpTFEtRzNG5XVMyCsH3vA/esFhttKGK/jU44ei18b+k5DG2mas28FTb1utaP
Od9bog1onFl6ZI/yOmuhdx8Bac/udHFM0TUNSOQxJtSxb+3dSCpUuEkFutr3ULSbFw0xsxCjJPD8
gm+c/Ma7HkWr6O+Lg4kV9dvxe7wSZgkH83dsR99Y/izuuiJzQJ2yvy8N5g7oja2Ou6rzyL6RC4Pc
883FotuYYFIMnemKHUpZJWlYu+oBWf+ncOxX0EaREs1maHs5W4cxflyK3ZQMJKdojBPVtUdAfPNC
hpeSDGAsMqhJItcpEtX3q2+MlJMzfIQ2GileQ/d5S/ldeWGZ4qrxZJCMh+Kv9SvRTETg9V1CVAH4
wSGixKgPwHRUjwKy5AKkpx2O9coqJSpA7qVgzJAERLa3TkS9Rn7Njc3M8sAm6XVVqlLhnSf+zieI
jca984jfwl5Z9/KzZUvOpB7LtoNzErPgPoZfsXXy1laVR5NkqRqoLonE1jKBiSX8Rnp0GCA1qnlN
rtWLvHrTyip0o0A2FrcLygknvEE5ixKRWz7szIG0NhXVc1vATwc61A8YLHwtrMAv/HBxL3pNfItz
8NbowZ2ZaRapTMk1+vEKF1arQ+oG7tVr1t1s1Wwv8Cs8ZI/Wy1C3mPuDyDgZU8zIaYNjc9EDivvL
vx6CZMVh+5EsKxbo3lM85jkUErPjElAxzrv05KndXcqM/Em/rkw5HyPzsBi+ANTDymYisTelfW+M
CDd0jxEWhsyu5cYpj/DasO3h7HPHLOBIpuHQ5ui07xTedRdfWtJRP+5bc9wXqTAFn7MdX42AkZYl
dSALG34r8dLE2WlocP/Ut52AFUvLEMEfx5x5wRrDib+mwcyTdaoFP0x42vhctaINvbSjgP6xLidV
ybY8hRl2/WLVNIH6YHCT2/40HIJA05BR3QfBZeMB2J3VYDkG7/2HoTf6Z5EPmhhd7oIN9q5PZmYD
MGNIu1Fw0Cht9AsLz1rPmEN/CuIAkWhIRDqUM6sCpVU5d3/xgPN0SKFSc+lefdR51iokvkFUnK1z
O6S/garbB4eHXC49i6euis1E5vWo6sIrqQEKEfaCvN4zV7Rzmo5k/hhazVHZvYCFvOWHu1yNw3YO
IU8ORr20uiwy1ELYSc+1cGVirFoomTu2rey7ugggwtMAGGmKadAFrpXrtqkhE3KuquqFmlqQ2v0S
Gid4FOolw5LuWeT8AFih1NHclWtqBkzhMxbXP3uV8bW4wgWHjkmpdf2FwjeQvVPW0Ym2IrEq54dz
XfqBkJCDo5e4W+3vheaCGK8QNLDsgZZ3YysjxsFKYXpJRADeNwB54mS/t1cSCU8IO4xy6fWMszDc
SPcGBjNptHdbUJtXPHFiKGsBuHKSy2R+aeZhicR09pZTOB/fuAF0oW2aRt7u4/XpVnv6TUNqEuL7
emdbgncMK5Sgx0zChf0WgIU0ihrO8vTL5uAI2uFAc1WoKtFP74Mb5qUE+vauwXBA4hFl9BLk8uq1
L2EFE1uvK7U9lyTrOnoKvzsdZSd/ZDlh4CsQ+WUU+iNtnjPQGkSI+ijpTIcxSppqKQ8fPDqtya3e
YmpE/FPlpDjJBrBqcjh76lNVBIlAv97WsdOxNL6qvLI5V+Cz3UO0LB49yfmvxBpKP9oXeAlKWbOf
UjMyrhPTMw5uTB4W6UG9KZe8fAoNuvMWz0fxChF7TOUU9QjE6Af7MZq+yQp5Kzn2O3puiZg3bvW3
M4p+3fbRfYME4tB3ciqxMQFKQR+XbCzUCckktwfJuFosJ04+IDLCqvPQd5fHon3PlhNA7F72HahH
dhxzwaWbVij4Ux8cTeiBHK0AIxJIMy4jJN1r3k5568oIeIesN+HQ4eKsE8GRMgck3j2qF1B9Lw1y
eD67KzQCHvJJ7E2eOC3VCXR+y1tVHHHGDgxU9WUh6eYc0DYOHpiyl5bLOp5XcFOJgxIJ6hZ1oQUY
RAzvyAPDdqkip6K3J/lpb1EZoe+2ngRtS2ak6Wnw60DKWatThnAwjnRAM3EmCG92aGJK1o8IfCJR
1+2yHj1X0mRAEMdGH2cBy4vsRifdXvvDfxlotfOrdQSaGl7mlDH4VOEnA7WRkBmoGTIdG7N2rrrg
/3YeeXOuBbHersgau7EqpOf+FeHea7Ge3Cx1ImYYODjoj1VGnuzCZK7E2J3mUWx9zuo59CPJ4HTP
asQJeOmKoDmv1xwdHZH9WMbzP4dKoGZ4y7CBbOFkvDJD3oEihr9HJ1x64GZri+RTEHLtmRcqjZfP
W6ayaPkQ/sCZFgVsuw6Grz+wvWI/MYHWUeJizUrq16oOOBUWV5JN4sAbpztCLxhrlyEK6FZaQJTn
Jd81TE4ynjMKscpD0sRJRkVXnN30avjAuiS2FqN83F4TXV1EqAg8ILI+VdSURgyMwbbQlg1nM8L+
AetN2g5ZwNJfkCmCqR7/MTTmVHtJ0xXiyjqBvZfAugd95Hug13i0/YiiMEsbDfcwQVGHXR9My11L
/QFlzp0YlkiBwCvGonUmvhZCa5n7FZMET9lejkUuJbHnjl44mj/X1lg0XhmQd5qjf+AkS2Y9COIA
4d6LpEW0yu33/Vk7kFpw+4fvorDoQGeOfpraThSbNGoj4CIzM8AAuBgdFaedHHFPOVbet/rhq59E
Yo48+TpMyUokgz6EolfybHn7cbc29K6HXYMq+LQref9qo8Y3HEyQ5/n6xnoiJWMYYM8rLf/BoCCz
daemx9u2HrotmeD0Tp8Lh1S+yPmOyLD3IWUjRxjIK3FuOwvYDXZifRMoVtmlfH7xbDMyfYysgCK8
3bnKfeM9xP1CDVz9/4L7s0gDpyRSm/s2RZUWqnLm3jdNGrcuDCHoqfOJRckSSScQolozWzD430q0
5ssa5/VE2WnqMY7yBCamYDF8tjrefapyr/1ks6U4kenejo+wSYEeexOMU9NiZvgWR2L7yotHC2/V
NB7CIdmVl61AeVc4ROKn05kf7jhvj/ZlTiUjauB8UjGSAJLjIpY/CnrFV4eU+uZ001Me9+8vrwyo
IdjWvS8miiejcjDW/z0xY0iUyivCfwNKjw5sPh55s2BR19Lm3kclkihp7ekUW5DilM2zQpdqO9UH
bNLKPs7YoIi6kegoGOdzji2hzg3IJZqPHuHj4AdwYx+BUcUAw2xTJCwvbrYZS/UpNGeY4EPEhRRY
z2cVnyJ7AKo07X79/09hXdiKUSCKY/+qo8O/+SuvtXg1zYt6MOeD+s/apLRW5Jau33mfjvJB6Brn
x2L1HniuQ+miBUHjFSk3iCnwHMECA5M8ZEuneuIMEQQhGx58oq9TowYDVum17v9AQoDw+tFzRSwt
JDbzl6mTlKWmILasQfkEqeQkFzGJrkc4n7i3ASr5K1T1E3GmDYj6nnzySmUi5/3DotUW1CPgeQHu
gY1vytmMsyjK4MLlRDv/9WkVms+JujhqZ81OJTSe/AT3qfD18fzyr9W0q0f7i1narxpmXOSvLkHt
3Z8i1piArOhY4X0rgdWCHKQCbjLQWliMSgpvh+yNq3lrm8IWtU7kLNjqtIYneYMM4nA3IqwQXNia
CKI+kKRufgLc7T/akz4hDgzdeZwJ359jWArS0rft5TxFiZqUmDJC8KnWdUCsruw+WYW1K3383gRB
TZpw5YijeUbkTcckbVUPn0Ab4xYbpIbGYLiNt/QL5yX1oZsNEyI3SUZXnz8ZN1F4oZ0AS9jl6zhA
IzQkV3rrdeAfyvFHELKvb8nzHdHBFyHceb6i3GZCT+ASQPRNSQTVBK7P0uP7O8IsYY8o+/qSwth8
8/HNY8NG2AdstFFi9/qmks4bfooe2nc0pdbxFhoxy37XCghpb7R7uDDpN5ehnM6v3G7HN/6+xfFl
W3oqTGhoP4TAJOfVkCm3i0SwSVpH6AdUR7jT3mDwM0dSQhmhTvzFdFc1UYml6Wt+H/f+KnUYchcU
CwclWkJEjsRnPEZ74H6MKC3dCE2KjF8KEV4xwMqDZoEYGLaDQ2Gtk3j9YU4LeDz+h+3bIzVZJhwu
eIDft0IymHHVe+3S855CxueFmxDoEW/sEwnBHRgEWKEXOUeH7bVA2zexF6yO2AdHCUQ4WK9F4mKj
akIjtSGsAUyZY4DMK3BIpSp68DxWvDLCmXwxFGirO5IEfilGsp4MleSmzGgubaY4g4ca/hyw/+ts
yoRORNiyAvq/5osLWPJs4YH58OVX3QNddKNWnHkLbmnvniKYBz1bL7HmnMiO+egaBbb/cPvAlOXZ
VRccfuVYD+3zebV2HTa6KQ+879Ls5GKWDazpXVC+R46Y/ieJ6ojM/nC3aDGeVTBTwcbBc301i8Rw
PjRbn3ofG00S/qhEzWdUvd6bl8RqePjLf0iGGaQSyNI+k92OcjXc9MSRmTp9wqWYXbrWIAbR923x
lAtrZepJXNAInMcjOlYJQcu/0H0JJyeT9os3RFVnSKweC3LoTmwxIAoBSMgW/UQxAenVMHT0r1Th
0BbWtJWrEsQ95yKex9cWvMF8vBbjGxcZi9JECEkNr9z48m6BRwz+jXe2SPdtT50GG6Q7bInDkq6I
gOyM6YpyXKiqzrBLUzYVBlceZfj1itJTAvCJ8GpSR7jsSmhJEbss332xAblM38wZ0QfHZl2svtwF
0x4F5x6+cKHJHZFXnxQfk24Iwytr9yHB99IeOhyRCDiqkm1LiyFLdGBjxx5ouSDOgnfFOz411/uc
Sp8SYca+Bjx9LOjdegIh0ga7cy/NCRdwbC6i2T6WtcE9/asP4LTMdkV4MfskV4FH305/Abdu3YXN
MYWk9oKzwVMe/4VOkSqfnVbtcoxaDtGil6wGh35dpDqKA93oVWkgnmJetP536DIcZvCKT40SB56S
StXEMgYgc3o5fc3fanTre3KbB5JM60/SYbWI1JNJn5yxcen1qzHSm54pXWYBqFeqz2J+KloQ8RAB
aOoDNnMOtlUzQfx1WdpV16wuEhGPlGi5OqBbWTSODDhOBl6H77cZ8QkNI2uu7UfmfbJIme907nl5
bk8Ro4jpdDjcSksIBu1pRT/01tbPXzAYc8UV7tnPLvGGGBeEeyWokHMlUrGR0oqxNIFQ86EJINjq
5EsGaxByfh99Ax5jPAyVvF4iLGGMxGDQWUEgw9xOEgZPuW65eCThB11GwjJUpwo0S4Svv/hRKQ/Q
ZQ7wD5ayCr4NBS/fVSwLwBYWwMAxVNINXOGBqApXbzIzoBYM6dHip/LdbZ/2Xq9R6Muk5Iuygr2H
d3xkYJ22fCxtU8eRwME9SupcYdpvuyGHlT0Jfc6LmkvutXFujptaEEr9OanEEAZY+aOc2vu4mDw3
oGNCJSr8D1sqqvFp1uHiKtotLJQom7DoX3gDUzixZ6FNkzqo9sEgh9LkEPaYvFKziAfU51UwFp6F
e/RT+uSBT3BeUizKpIC2lHl1ms+y6N/ZMHsAX8MUaYGBO6Xug1UAXQliTjHh5iHc5Z+gRAUx24LS
2MO4g9iwoVDFvmsQj3yhJje6neCSg6HjCTbpfEglaU6MIr2bF5cogkbIW1BCQ4S9YVwQJmRki8XR
9STUkptloRj/5tt21xc+nGxf6NOPsKzpF9aaIx1kplyHVenFVZwCT4q7ZTNPvepXnefOy4uUmG7K
8KRRRLlkbZBibjCLhW5+jxp7Y+7niuPK5KcO9PD+fZ8aOm3vlHgIduslUOLVV50IiliU3zdSR5dH
wI4xjTiDFvJW4MWnBTXoneje0t0morHCId3VmUYs887hFue0+mP32J1HJD0zXk6qTy061Uxe9i5i
KlOo9jpZj+9IcTA2bTVr7oJVd0MDJUa2evDiIKr1WrDAFqN7TYAu0kmB3JNXTYwOUP1kdyJr+yJ8
I5VDhkVXikrkao9/yqCAh+Houb9KBi35fsXrweIz0aTZ1vZ6J+dU/Mhvoh7eJcHinsiOfXc+QB7+
nUKFtdhkDEMatgbN6P4f+mqOj6DcrQ+77nJF9vGTcm6/k5Dbg+KPWUnvrR1+yzPkWo4wI6JaWo+v
fl6u9C9I5QOG1DVvcHoupvC3jZUTl5zlX8sBVO98axJdxNRV6GCqoHexKfvbcgYNzE39sWbR8kwV
W4Wv1ehfKnwm06xhxIm03ra8FwmtRfC2+56sUo9IE4J/G+GMq9eetA6/Top1zKqlXN/xaxhrGMG7
JSrSmJnw+e7AC+jaIL0g6WyA6oSAxNaIj1m17m4hF+rguAsKMbtl/GrWsXSVqTTqNQgI5vEGwuqP
FOi9ilOc52451NhA50hSmxvtrsvZcMB3UfwPxZ2nCRdnIxhbvXHkEHQ/q1IDfHLtSEKBBX/hfRCP
acecxJXqE/Hy3tjiqasr7FuJpLZh+QLQ3ZVZZY2gp/kKJlbl+3F//lvShvGPWrvRTCjsGCG/Wkxl
4INgKoB9QE4CP2f3c5XT2xBjM5xtp0mwLLyEnzAM+z40lr6S0ZNkElrszP/1pa97m0DNjvENr8ey
kSsFzzDMpEajkqEyBCXM0WkJWYJ5orZ7sGrKjqmUfa4YGkvdE9h6lOEFj0ENWobOB2lwj8Iv0jLL
WELuM5J5KREOg9AxqxlB/+uxJ9DI7CyNeIMGAYDQiTSHEfbkh50FCoNzu9n4JE6DGndWmAP2TbON
s4sb+A9BWOM8FEULPePxl4hYVrrdX2TdT7pzhIL/0Wa4LYilJRS3Je9kYf/ji5zTctjKeJ6HgROv
iHJpRSRWfJNQ+MbTTrzEaTyJngrMJgxIz/gFZoTgY7lPfR4ijb88b3/OyqG7qz8Ftlhj/jz7kJd5
Y0s0EDr0A5hqWEKMqbeZV+yFIiDAzjSi7CvMGfMlp+dCQ3f355Vg5eEOYu/ItndlwYTGgZ0YUwvf
98f2H1MeJJaSKBDkhkoQkV9AqEU+8u+Em2g0TGscdcvKxuvII/ipK7guNSdNaiZ1nspcDq4IAi10
bXCLQEWs0hElb/7CLRViJ1emWILNP+JQ5nA2zcYKvrcUC93obKtOfw5imTh9d3US2Rws3ZRDSCse
rZ4wQORcSGCG3A5MyRUxsYjoaVJ8vX88q00az24x9p9SIYL6hxlde9mnmKcAVzyOdVxIzRNYC5b7
2Da5YHjgJk8A4+dtnyPDXGP/oujoEeKsvL7kKH7xGHLXUEo7Wd8VZyA7dAfiBEgT013F2VsPAavX
KPVItoJ7CyJRWd+01yUHO6CgTdkrffy1w9uVncz9ZrGwXWbka/Of0+o4lkHpNe5tropiIHHUp225
iQAlFGIVVwtQAdQpbo5DVEu4puCrw28GhgGAdx4mGsiSMP2sj+V7LnHf1v5Dmz1TmyqkhafJkWsy
ivln+xwCmqttkpIUChtYF4D4lga8DYKlOLEDlo8zXwHeXHXHsSfVqK0uM7KatawFoS9C9OdSfpsb
gFTo1yyFIqx8RVTBvQhezqEzIB/vvf2sEmjOPkvRrAQGxKo8Wi/9iJynodHw01cW8+aXHJDXABiI
YlPGvnJrV6IamCL45mymrhVh1yzJvnSH+V/qq1/bc8EXMKPaHvIBh2bXN6MUD4pgunerVy0QU+F6
8yCK2npNmovMwOFB68nzvU3S4NEUiQUFeXnoHgLEdSU4NWkrDQuWNCV+yPNyF/nvYQcG6sZ3XOln
ThbsudhV04Zi7Yo/2eN8SeWmj2rORkmC03d32hPjPaNETti3nZlmLeZJ7reb3EWSzulIRCQ+wN51
M7Q+WQa0MQL6NRKZo5hEWzmHAKqrg935ThfDkSJ24ttGyBbi8YvOgfGoaqx9s4Cu77H4EPVMTEiq
2CMnfZj1IX27eIJJxMQomoojOS/ZcGSKNActcwpBMno1fBYRNlLzW49kE8ipoErbi9v2fuF8GJQG
N+JtxpeQrJsycgkn6rH1dwfnhCDT+MS1z9zA1LADzwYzeVe7zugBUivAgl0UMQAwsZWim4tpeX3e
ucuLApSiv9wz1/i/x4+LxO5tj4rThOCckvBWVwpIbHhDk2/5xMvN/RY6EnU50s2x4Yuhh6pmlyl7
lA1v+ljULubQ/5VvW7i+TVCOKIZN8WZIJuEmhcbrEtUxOiFNrDGyybD4Lcr0NWDyCTcFk+6tJSod
P0PvuTEuFz9mxtUH9SRSp1glQWPK0wL+TySut2O0ozAZ/RjnCKh5KW5XBpA0O9G8OISr//G6YWxY
eHp60Xn6lAIMXbIdzYQCC3oi7HjK6P5Z4T9TqiwPCej9NQQN1ES87jZJDAeFshUcOTWK5cZrOWMs
1d02OMf1QfUDoN6Cx2e35bTX510r1aA8hU/nimH6COEXEuQxhoqY2zSvHDQhxIlWvvCKhFJDawWG
tWi+azBmy/wM36dCpCHOx7ceXRf52/cg+cfQklE7wnWnxPGQ4F1PO/3NGixbNTrHm4mv4HkCCHq0
XL/dpKFq0mucmHfZYGMd/verLiHq8SxCaxDs+UAr1TS04WZaA9tusWxGeb1h0ArKdgdgn9ey7q9C
5MfVuNHTxfkyLsjDPt7jiojQ2HnD+DJpmq/Qzgqrm041XkOir3gp8COGGsyWqRSgXPqkVueNP0yA
SNDwvoxI/D47YbnKruBvzA3Av0OYzZMN+T8gnOGdWjudoMPUqc44uPnnMTT6SluMmay7J5OPbZ9d
tWuBA+H8M4FLI5K+2Rye6DcJm/kGJH0vldwUgPP0QeyZHzEzXx5uRIlD3RrMJaJK6RiIsYFc1LV5
tDJlzwNQfTE9XaMX/1N+RM2ImN4s8ehIYNyITXB9GY989Q1WfW5AEMNG+tqszrcj0iC+p2Yu5fK3
+4ADq9LD20MpguXcnBvtVDd5XD0jmQKfDfhXb0aA4qtGQKYcXy+cANFbALhOrgx6aOvXyCXI9iMK
8UXqdAFesl3dFf0Ie+s5Jco//Wfs0CRkdocy8G0L5gKiY9NtB+ICiZ4lDjuQaRgEIeOLIM20VTVX
1k9ITDDnFwzO2qNgfmMVkuU5DtyMe5myHGxpWYzGUFL3sk0xAPDbUpzBpkPUChqnFkfskwyIM8t0
rob6sGaOJZAqzoQPx/hPCfdjWXUf0cGMqngzllnOUY+UbQWcQRw6XWdC0jlTdeJoqwBAI83+Y+iQ
0D1CWIlF5Qn7OUCbv3FWpJ4wL0/p9p3UPM2jMBTpqm/5GgjjGrx3Funa5K5te2kmWSm1jD9yC7ec
TDvBZrJWajT7vh4zEFpv9mVCTaHrEcDvBeXmQnVTzQpBKW3PG9DBWHtVfchABGSWAWfb7BoKfhnh
s0dLjJvro9WfpvRVbyQ/5rrjtNsQDETQ3vm/hCq3xgPcZjX5iCZh3k2ol5uHJ4IQ095md3+DFCsR
U1JeND93yIbEGNe8efsL52pylCsU4JOFmLs8s/yDvsK48D3jTySQV6udaB/Zfu+MXxphRmgfpAcQ
MFnPPnqz9Q/CClU4YPdHjicMf0hlYt0EBnqC7EDLEWmewCNGhZVYxmnqegNFYVXxUNmhMpFrTwrg
uz0wtWZKlts4/b4U5nhtMguDlpSBW0Q2Ey1k+NUCBvomkfiQjVf4jF1wHMT+MVmbJsf2OXi10QUT
AJvKuflzUwB7G103aT6PDwzaHdgEv6IIBaAV5i0B2zNjYtJescRr44RgAKGwbXZzqQXAdGxhsOs2
IV2zFnuq/ab0oMwEyU0rFu48cWjScYkTAPUoaJuPvcJw51EPSE6c5oRTI+raFHHV8F40V/XC4t8o
Q++0jDMWnVomZ3RBWv++4nIU2ymQp7e18d2H/dA+CoxuR4pqddenVmU/axQ6qKeFTjg8fguiYfeC
LFR6jmz/w0hwz3xldZhG92dovc5BI5sb8/xWxfG7ye/DIA9bU12hnb1+sxFovVjgWQ3CgUwa+Jya
Klgx/AahLiu08/oalSqV37HlRXKplXmdC2sNOBhLWyAmqxDfQ4PgDUtHCstD8UoeMyr+v8CBrwpY
7A2qvD0aOetiCiydi30kXQZFCM/Na0rmtoU27EtN649qKXYnynirb5B3IUwt5nsfWNRCpyw0/g6V
dL9HNN8btknvxTAHtX+u4r8lwnUFmHC4CPF87pcgQ6Jt7nSnJMimt9zU+qZdGLJnKpKQjQkWuJZD
fKpx9cY5eIlBgDoGUt4RiifAs5BDZWBui3ARG8F7dpRehVJ60+CWASBIGQ5Vmko3wcou5mONQFPL
K8c3J2RBwMsT0Z9+7h8O1ram4gGpmGUioocHfPXwPXNvNj5CoNtiegj9MHY0CXSDQq1I540j0BXt
C5KHt9VKs8bvxVFfY4j10WqqZLWiScIuul/L5mGkogk9ZKK4HmBiWJ5KB/MInCRoekWiUY5bd2C5
JHLabZ5R95xjOzcDNgj29gzXQhOmqPqCNjlr2N/nt/TmF0NXnM53XAH7Umg3SrnEXaajAHI4LIEP
nF7XQDxr9yHnv9FZTAsSn2YtwMqAa377pSvlNoS+53gQCBjVp+UfFIc9y9dlTa9ZNm78KUYSoEyt
gn7Ns3T1vqlA8nEl57Af3bGCqnOAik/SNT5nvNbhTDLrcz91jx72Ed8pWswGMN9ttu536P3SV6yH
Frtn17NqC0W4cbPmyVoMIVxK50blf34cArksdyhGywHInGZ9evB1ATQxJzCkHpljYRaNscqOTHKu
7K7l3CwptzUu4ouJKJzVp0q6rHn+nvic3PYgswPE3X0c/lAjuci6Uj6H5Un2Pp3HIj3N8yZxsug0
LGwFHhJdvTempJ/Sw9J83MsbPKoBiBxEVrO1VMDQ3Q5S0w0UTdUIN31ja6Xdu5eMBNuw2Zw63Wyb
SzFRF2qIko05uPXoMnS5YH3NipnYYEfczFbsRVi2zt8CuQVd5s/d/f8GYPCeT0v7NpGwoRtAUAJo
0DP1IC89cTbg+pUjWeN/Mf7ev1w8MB1VvH54DunVc+cMC2Oy72/LgZZu1CfDnVN2Ah8y56yAR3jL
eANg0HLi298+gDZCseEWZmJ2aGuRyPcWuYWeYKFurHS3DT0Lh1zeZ+NhiWkYYght45/rL4Yrv4Hs
AmsES+JY9/jfoG2POBDT3ENNOeoPZ3d0ZsszTWfqizXd5Rg0L2okusmYb5c7ERtpuSLP+yn/gbwI
MyBvZOj/fWC5esiqw61YfBJIPFOmneu3WHozdgFGvv+kFB/taRl04V+zQl9moYrvXM2goF1BiTG4
qLETnVgdufk9AQrbIWRhPZIjc5kSsYrfsqtZ6nlXsUIcEiE+Xviog5BR3DRee4Iuhczn5hclYuv4
weW7wKiNmc7KRGhY1zfVsBZj+UKApHabl42lg2IAZmm+57wRwTWBrzzi+DsrdXXca8PG7pe60RCv
CWInfxz17KljWuEMFffhVsAxXYOE3gJJTku4hxmDgpIL6PsOz2HnaWyh+kvxjIqVWw7sgo2bCLK+
Vye/u29xiO2DjCeYPtcN2mAq6KltF1NdI/68FXCpMFOPyeg/KRcRSWgemZJwB3XVh6ngOqoAZtVT
iTdK/2I/OxrM62NP+hx+jdHVfj14yJNCZW/s0CWumcLtaJiwOyZlX+G+kcAKFc59PxwjvoKT4vIb
tzBJLoNRXC3KJNaY5qd/XghZ4LNNrvEhdOWYLbOcIwCiDVzjazC8/T2mwxmVG/ULU+XuhIctdXQC
SlcDUh9lV4EtDaC1Eok1A84coLiCEcQDVhjEckdS10ZZVSrqVihW6TeMdcRW5w8xWq2eBM97pzlN
HSSFIhVAfWdc16MOUhdcUMPa7saxuEbwMMiEVsNV0FTMMcDxdJ3B87eyJjQV1+ZSNrgdPTPFRufp
tuy4NAznX4hbAVM6ymTOyDj7xOtF/x/UoyWDB4xNMCZM7/RoxIVGiTzNrcw8/5hCsfRXr5yVHCFX
/SbMo4ZxwsW3yENCbJi8uFxh83WEcIjVUlA8mXnYJjqo7jbF0pjCmL42IZ6yjlbejhvz3rulPDRC
xJyjg7mZi8ylfZfyUBwkjyfg3d1we2TLErvbuEu6RbpoMJhw758mQvlihwTEK0eqIGtHZYRinAgR
eNYinv/9baF/tW/qVtagZ0SVMAgUqVmoB8VauEmKuKq2HWXFm8TvzCzT8nmnPLPjnxG4dROJCzVU
BQI5TE+EXQELYVfSOFgqPHCXoyeoQRpF5+uUgwyXMJqnFwKNQ9joCdolr/XFM881kraNBnBAI/Vn
GZgwcX7aOntiYYsU0yXNVc3Y+X1+aojGu0re5hYAQbB8Td5XFpmRx6kZ9v+V7PcgCczzALc1HWdp
2nH64B72nDw/9AOI/mT0WGqQtmdUUbnO4nNz4vC1en6Gdb4KfjecMzovxvdCiFg239TJgEZ4EhV/
ny5gqkhO/iWD1uUwoddidxoJF028fLsK/est3j8Y1MOejQ9yH0UG2iPZuQdjrV+3wPFgcgdX2l3P
JVP/TW7seWqv2q4lbyDNNREOiUrZmjk8LBhIQ4t6u4mt+/wNCAMF+cEASVHbFNrSBBMs33wq1b9U
NYPHWcnkWUwNOTONdHIZJX//WgYPGpTXh/ysM7HjFUUTeDe/mWB3HUgCof+WLitutCL0/vaNFRU1
b9lVCyKNLXQpjMRbByT79RqlAIp+VG4Rm5aa8ykd7zs0QOuNVEGMnTB6ZSOci5G/nJdXPns/KuT+
b5xdYjH27jM0PqhaVgGj5MbLTUWPmabrU2QjniYptqx5EsCV8yRmBEW5x4BUhyPX377yhkXSDWW5
ICeoPZ66dpaI3LjyQKSNo/6fMKYyAd+zvYEau3Q5siEK+tif3bt8ZsU5RUhOagw0/Yqyc6QHt/Y5
smvwJZFQnrHwFk2/HR+CVagokYOhxITSawcascpms3h9l7iVcYueW6lo9UI3XNHXp0BCoSvQnPPD
bAe8o7lcYA36AKvO5GmyVgm9UrTVgGFWAbCcRau/kziKpHMFdntMtAzpsRAI0zyszc1/c+hy5fhz
BFhR6guXQ7HmopTtoThDjDSbjL83FpPo5WEck//p1LOfA8jkqv3jLSDJqVgqBgIcmEdEHmFPWqGX
IiGlKTNu1+r45Sdm2AQzxoaJFWqRbt3gYaRHqcKn4yeBTEUrNYfV44E2pAWifnhl+5n+4KQOLswX
Et6IdCtWd5jJ7xmLS8PRlluAKCzyxjkx4oGdBs6eSz9UADLMoZO+o5SM5v+j3SQwoPgnHOQshbyw
TC/EXJJPJ3h2eX+87Pzlsj03UQ2uSa4B7Z7eRMylA5mfSSAsb2O3PXZK5iv3LfKX6n8ILjRVycXA
0NPoiBaZ8qKaTHH+gt8SkyplpSIeBWFjqdI50YTagzGQ3FcJX8q/Bz2Kaal81HHS6+y0GFHqq8mn
8zKvGWnq79lHKZuDee22BvqLil71tduRQFtfgCRzuuGE8CILMLmyBRJHgDHB9Yg70QQy5XN6pESf
jR5rWJRX5ToOYNHEozNqrmLjNEXnjob+/2dGttS3bdCHIpF+Bp33tu5dM1uoJ4PaxW8jQWqXFH/v
8uToe4AgLPfgIvPqIiXlSJaCoVnYe0hPCDTYv9t3+ehZy+xVnay7FZFt5bSRwMz3KIZR3GNP4p7z
0gtHwYKQIlyU7bmGibdYVc/g98HX8r6tgXVO1MIR90NZd2ykWURVkBdHwVlDiaUsNhz2Oe6nNekj
VOhauhYD9tXTOzstRNjDVFNMBHN4M8s006nQE10bT2Q7fR27esMnfRuL3TUF22O1YXs8qayNTk0P
1ovCvVFaCS3mUhMeW2JdbRCEcSEqYNnK3AgVh4UNNAesAeEaBGt7ooof/ocXPM+FSflQBCgmgcMe
wcJpGmZBESpIfG6h8amK9Sdy7cKgKqCZFq96XzS7NdZ9lYTjfN75n+c4wAx9OvG/I/IK+vBrpu5p
ormvNfNMW94NN87vOPYhmn6/V1hWvUa2Ql9B44rxFo6pJCM7/PBKTuvRbtxBja7uvjpNDTNhH8o+
aihVbhiwyx7ea3m//la7VD20KKB4ewOY+tRqeVHLynyaoHvtxFJ5XNpQRdUs1LpQ2hZcIA1PZOFQ
pf8LYmADW4Naxz4SqaKIZoVh25jMMOkd6lNxiooIz5XK5lZ33ZH5/LRCExbk0WsBvYQixD60/b5Z
xFMPrGkzeJqtCAYjT4gujNlH9qyRP7JYP+ks6beJebxHT8xhRKH1rQkxRXYmSXG6440Pg5BaybXC
Kp1vsJZpIpp/9fjbU39RrlBzOUkFNdTsiONdYyjSbXWR04xfDLh4eyUQotxke8umn0jTDr+tDkgO
FzgCliLZ9wt5yljblAtVP/sGJV2sW/NK79Xn6L2hixcyCxrRE1FF0+CHO7R5Q1OIP4rWMae9NPg1
nEXru26X+q/lBPssXI14R/ER2lpfQh3jEzm2SUxMuJiDuVfdBOgoAnO4OCc6sJ3/6u9stlqjPMX0
BxBSbnZ2rG6vEXMb6hcE6Cea8iNXVF3FFzjl55GCjVbTCkisMVf1FBnRCT2BvvpJA6rXSR9qM3Dt
ivMPoxda4+qglXN9V2LNIBbL+AE1XScyBSRW9h/g/3h8aaGuA4DMTTvDcNo1likUHA+LgPUwRl1v
4fiwYG4DSs31Sb7AaHiriYWJBrk11pUu5tfnpvsj1K3pHvG+Zu4fFrvLtogmEEUWk8yg9qA9TqA1
XgoxvdwbWW0Y+vgrI63mcASl3x6h5PqeS6kq9mWKNmXE3j6zguT+zBq2qYv/lOw8uuXYwy2Oq3Cs
Gnnb/HKoNMC5un8sYsL334OU/5GgAxdQQ0UBqA3lRayiAcJtBvZWqsTiKf0S12MAw9lUEgv70Ec0
3UPhd/WQr5ZCZ3S7mYFnO8ovV4P1SJURXo34KiCp4HQQetjmqaqPlk/X8N0fN5kRA0oQi7Zymxf/
W88iyLjx2GzPVt5iaXa9pdGBaU9TxauaGSuZga5qU36qCELkYT/x2Yk3OF2MPdOkYa3hdU74qiE7
dJEEOGhcMY+HGZTIiIPo5EkNvqX3md/qwNDPfhdcfou2jvfww0qamQjD3PdvCCyxJtoKdBNFHPon
JmZJTDge0Sspp7TboOAI19NhHp50759RPfv3SYtJJMZK0M4tvkc4mdYAtHEc+K1x04Pgfx8CaxrK
Rios0N/J/IyGPljKt6iCcdmlS+WdLaxH6vW7nODfY/LD6A1wPuCZyk14J8EOr6igbR9y21OuRzsJ
D7zC+Y8kysCoUHe1RbMDYu/0CU+rg7/O6fBfXSt+xpikg9RHY6XsGUsRdBpyuYJ5RTap7pNxX8g5
6saqn1oCemPMekl4d5vHec7u/Qe5gdb+LX5g7IiKYak+GU5l1rROIjapyS72h4xzQoKCGcQq+lBq
6D6KkcaFx8lyl4VupQd9szGJR6ZnYOixPGrJyaGWYHvlAkrAm3tbD6GcnVhwX6kLu3aBSVeOYcfP
Pxadll4bcuzd8qswN7OgPFnFjRpr6jxgy03dMPkfv68HtKpECve2ipPhxw5wjwKrgxHv6eONHq8a
AT3J0HYWFE5hUMBQCabmICnwRurJwhGfcQ4+44Kxa8GOnO1dS9pSw1WGXROj98YthBfdZkekIjDz
Ajvk1DHEXGgkFP043RDQe8UwQEjSqOLUUfErYgTDpGGBvgvT1WZDIfMdvWqyeSuHM8nOsj2Dg/x/
vE+hz0gixr/TyNjNC/hOazIg4PlLGmyCki2SdG5fzzzo9mi9l9aa4z05e5vyVI3Hk+JaFqEnt3xb
1DFlyNbyyGKGzgsKwFTGvNCVrEyYwFdhd6/ilrMdFaVe+Fte21Vim3k7dIpWTOWJqdS+4mOx5uc2
OnAuDCDY1lGivDHMxN9nZDExWRKnencMcftvowvUOoLKtzp8DE7da1WvajfGw5WGsY1E8bX1kGuB
+ccJQMgQiEINHE72gyL1rJzUY9nFBDgO3LqColDS2SbRNscO0Hj/UkTSyCGxDYTtDH6Fi4NKDrhj
HDsOklY89vCf7HYAMvOsUO9YbVrzQCS+F/NDJUtg9u/Z+9R6+a7RNJpUY8TwqNYCCkf64r7CNe6f
3Iz9GlT7u+C1X/m2mny1OCFnIUcoS28qDc0R8efo9upaWGXvtFchCV0EsGQ66iaBmyM1iVz8Dy7I
qvmrQeZjXwXIvA0Huq1h2kDcKE3tLvqmkTPIRMZU6Dm7Wcfa8cIllXwBm9xQkS7O7Fip58cDVwYz
z0r4WdtK/fV1hw9LxxShlmdIGTUhHKtK9e45cIhamptYUkgVhWwkKvRutJ+ldN9J8QbvGwog8Bu4
riPQm6tFGgWH4GxBf3uC6JMHYHCy+Df4rhpmNLjcT8rNNgdHFFCd3w76VC65dGZpiCHrY10EASF7
Tfd4PMBeXM+fndFF3LnTo5Ne4l59dxEWdw7IP8Um9x0YQfUkif+2oRkgq5PBWyYpXfkWjXZUOzp8
7dJi6pHW30Skeby58TL8GEbNDrM4k5dWyEhQdZexYHEuC4wnYRawEYtzcTR1ImlYkpyKokJgAFtW
okKiRm2LrmrlhaRyIS87Iun6NOu4p69+HJ9pjZxpVY5SqaR+T4H9XvEuKPyfj4yM1FiVlBfN7C88
SU3v0QM0Gl2VkwCAlqCf9OOizGPdo4TahRtxYfVbMQIctIIbjPjLW1FWjkBr4kBtIw9L5KjM7BqX
ez+uwPKY6jADGYrU/foknG/nU8YdTu3ICujApwVZkjVKQfhuB0zuWv/vt58arH2ARoO04SZBXBdy
H7XhrKfSXXZpcb4W79nLntmMvbYcShIQsL/E8+pEbwiWFW4nYVEuqm4OAzasOC5GYacOqc3YvQBK
XMlf5JyZLDj4v6m0G4wD5aEvQDUZTmybrEvCz50qdJiIVduW/hqimW0aYxMh3Uxv1xXd6FdSvLlP
nYZwtp6pJK6MoYm8weeNdEs7B2sAf3TrPZmI4tbBnfpXUDBn+lcNYmn14lQv8CP2mbeZ+Qi4+WuX
1hPTQyKfUSW+SyIL4i6yzhtMqODOOflPFrVpuqX69ziGSNraFcHogAyAuz4otCrgo0iu/WLu2I9F
AneS23GpT18XB+qTaZBkhSjgrDptUejkXWk5fJZIM0HgzyEVZXcLONJb7uSEcbrDA9tTih2v+UEL
BOlSyz6ruXQqrEHhZHFb/M9is5vedFIGSv7Nm48z9NnLetS0SYD+9TIOE3RAdEBjWThBPhURNHJl
wifYyHUo1NUzQsEP/xKgGPZraHfRvMkB9TzqsC0CTuM2TGK+3s3XvDCcvk1fnVADexQwQ30zQoFE
ZY/vPTMj1iKy+kTMS38V2OQQZgBw+1RxtXrd70EJ3goK8H0Q6JQUeJf8tj6MyXJUut6acEt2gXbv
IZa3DH2sRxMDZPCm/HiFPYyR1EdnVp7VXn08LJbF+fp2MfxPVGInwVSuq5DufOMvNKLz45GcYWKC
I9qzYr2hmaPgbq9Ebw96YOS+H8d/W1zvLvAhMjYQsqMWziGxdbwNylJnl2rRFfVWQA0FTC7HtfKG
XLL8xZkZc6HJvet81FBRgRn8SrlvfpEpJq2sI9s9p4WWwQmVXyTtF7kRPnE/ZyVmCr2sDiUOVJnu
g+/6D2klQfHG6y3XAJlbJkrutIu47rhxPnhL+YQWnE4KLQQDLc5Ou2MzGbs8VIH1SwIrwCqqSFgB
igoBXQyL2y666S+ZNC5eABT0rRjtf2QD6vNEGLGbMjmiWrrDuFie3TbYzEiElm7ZMiuNudKlcUOQ
aNQDDzyotU9E5M+UW/VurfVnUbK//o7OQ9PzEFVCcu5E2Zr2BzUj5tqSxkYuoixlF8rlCj4gGCxP
tsmqfyt2A2KypTgCaHIZSb7JF9YA14j/cxxAzuxkTMvPF5XlnK9yEKlBA1rYvN5fULiFo+j/B5Ma
dexaXBel/aYH9DSB3bUx2ryzJCtnC/zQM6Ys+ZciT53fTqydds8RcUxQrQdjWkpbmmtIr3luQnEx
djvjVAj/1flHQ0O8fw2H1YbW2CvD6nsR+2R8FyeBrLmf4lS6s3+LmpgYP4oyvIwMDsVaOZMCpnHx
ZlogKYv3kggYpuZeYUwJceN7ThqmkFGxzmm9Ai4SHyGHOfCPKjbOnPD+zoRGbCdjNgxPD3rrq5mo
uYR777ChrlUDD3kltjMn+/pstDKXXmexQav/JGnQccBdlf2k5O7ayKz32CuWwU2n2WBtJra961KD
lC8i38Lq6U+K8yW/3vgqKRK85ToqSPzdY+Ewul1NieGudBVp0l8FIzm1uWZTH0X9myRq7ivu3dDi
Rom14h9qC9cAQRGrAVmW0uLR8xGN3uu8haGgIaF1dakRrbFoImaHjzFW8feYizRomVsO3YYjBklg
PFVsDnvTC0S7bm0wJNvGv92107VZG0uiS6ry2Qh/SuBUqNSk5ikLR/pMwR9su40f58ZaUoFA0dvY
Yj2TT4xaaGFoOuw+1JWN4MqnO5Aykn1ovKma08KxbEKc5cNVzu2DNPIHvN6m32f9kzzIh7NTLtEf
CI2V4lgMChfEnDVNQ1GZIp4Dd9ZTLN52BD2XtO96k/iuIMLnfHuqLp5dC/j3B4JQutYOZNyhgYI5
yHdYzBXjuNd3x7ZIUG2DHIHyJwIWiF8UziRMRFmL4vdsyk2k+K9S3oy6Hd9juJbLpfqkIFPoe26w
HZO8CzlQZeKcTzRM+aBcTba/w7/FfWLhIG5RmJ66YUN1sOceSLdn98TuHzGmlJJDQy89kwczYG0m
cSkGxcp6dTutWNjbfiYu2+Pz7xXdGLj/3UkO2KM7ekSHndjm04Bn2F5CeI9qFeVgP/GQUbNrJKw3
QHaYj/4Yn5F0lcc9/gqUCE2OSvYB+uCJSMXfCZETCqONb/syEqY7TEpdXe5NQ/5yWjs7CWaWZCfp
VZtuwsgksq7wNhBqmSnoCANrnwy0k4zv+uHBSdZNC9qesmOpag0eCrLoMfg5UT92PfNA0s3qGgk4
1D187Tq3Gf9Zbq6A1641j7o8Jq/iyLCFuiR8a6Z4/3uasIt8P32uaXPj55re26X+7pbibtSFjmvJ
WZ7QTdyWXyujxL9+sPfSwnaVCkZBPkVTgZ0O8Kr4tm1aH7xI6HNOizFO17C86gS2zFO3kLGbOxU1
aH3KcSyNNwIWFDGogH6vetsuIk6KL58Z9ZxryUx+IW0ySyUikOQkGkN2zULHIIyoKokmtnypyVzV
BZLU3CHrM71hQ1tuIgZykUvmMqRZLNPT5vDB5NVhCFFLFfIkIOpyZP4YWVX5ilIG5HehtxswcOLE
TqLhVFY8rxJjfJv8yfpG/g3ZVOxIj8Hrpco2/KgTxF36tUSFNVCVWlKq1GOqNJivqEwrJTyufrQU
7xlvuCoLrdqRk22jtqIqPYbN9mxjY567J1NtardI/cOJoM2q5LJV0CDxPBWun1b8x95I4Z0fIjOW
tYH1NZE3lOnnCzwp5u9XdAFR14zpMxtbCoRanwouvbf6pBDxbPMMIb2gaNLcVKb3Lna5vamcgKoS
xoImNUJce4mXf7WaWtt9Bh3qylhUHEcSyR6aBSROlk0gGkGlg2/wnw/M+6IEoV6MJ3IIa4jNJOcs
UjqEh8j2Q4pfOfkNX2O0Pebi4CbEhLWkuxz63PiIe8idJqg+qTc5PKEwjx8zKr/Pc7sOkQTZF6C3
0m7IJNflvQ6D9qS6DCzDZ5xF7sVj10RdxRl6oPJ++znQRuxPVc+yb21qOGFoM4q6Jep3KmPcEOC0
trDzOopQiqL17kMpT5KABlguMMOldSWfdKRZT3Ob+y1T1VPctIK+TKctVcYdrqBed9h0V/xbRl9Y
GjscRQTrDSV3bJvPoau8lqeSOVm70t8imQAdtQkjjbjln1EGEXlDADkzhOAHl5uB/nt4ygSXKUq9
+ueQ1jJVEFLidbzknouc73/2en8YCQwOXoGCP9LDDfEx991X9lflA4khC7/qYUS8GU4JxiwgltTU
4qE7C1z92Xr1iu0x06ju7UhC/mlGv6nyG4SFEl3b4SLWpd1Wb3+9t/sWBjMf/pMgCH3XyfZrKOu4
lfvfP8ZSXugxo5H5E3lj3R6XXFTRNXTBf4qHqy/SkMrpCr7cWAxT/Vprghkb9ojNwmoHcmBiltaj
/cVmhEaBSayNsyBvaIky7BmfRqAl0l/KzQqBJE5LpQ1y/JzYk+WEiLdja25fHK9qmxZq29hl+bP+
w5WS8zrYH6R46bzqTD+61LiJcyiMUY/hK9An4HduR7115VJlI8Chm0Nd6mOVkl/seZdaIZZgVweh
rbf2VrstBm9ru5FNjgcZbEUWAHT8urc1AAz1jNzADRnbp+gr48KuBjkzqetV76huDY/qVvl0kB3S
NWuV/9p1XzcE+pqdG713XYlSYmToQoQEqU2FJQfYufgoQWpCuHcs4Jpmk7ypPEvgMbnP4dWvpSAt
2Dx8Ri7bzB08d18NMraTRV9wQiDPp7P4foY5D4xrm8hQ+NVMT/K0GJcHX2g+Xz7gFnF1vD+6vMB8
NFL37VjkH0KOlrcEnIrqxIn8NL1j+vcot5t2HVRjC3gItbP1ytMx/1aXUvFepnCyL/CciJK4MFGN
smd4/7eZ/ID59i1VV9zZiUytnnAHcWfL0sQ0oFVFds3lqy3AEwXcbBE451cCfFWfRylC+Hdtf1wU
Sti6PtqE1XWrJPCUekdCXG0m9DbNgtS8TYwJNTIvSw2byRL7b3dTCjUrNTV7idehx9TueYtDbe1f
wv4fjztkrZAlQwiUmzhKKlqnXoriRV8FKaPxfK3UvEcfowiFm3q/6I8VI/bFZelHm/c7eGg/8G1o
Zg1FfQyxKcz6alQfkWVRBGoCOd8w0w6XFXa7f8qrZXqqqImqrlxx+9PaoIgsm85Z1swDaocTUmcF
5SJ7tzg8XfSYgEugA3vLbQqQdVB+uBvp/kJU1cYxa6UaUe/Zxp5R5yT96ilCZ4XbgkEQi6vyanfV
OoNbCUd/mjFNCmHEGm5KYaI5upTeh1dqAaZbcMp5Z0tLAotz5MgUDuCNF32uHz499oHkZlJKfWWB
lGVb1d0TAV4DqnwLlssVNVK/rz6kfPoTyoc0nIr77OV/+8YcV4rvBpWn5XZzlVA966ZW+q9wQN+r
4OZFKwj7ceGhYNhzy/VBqhhXgoZEZmIJ7RX7MuAOF00WC6ZTS8MxXlnFgm/vXhbAgKSYJg9ZxJb0
lyHkE/zZP+UcnSKADKVE+xYcPFjRmIKULMrTUFqATW+QVvhQtcpNLL6TpOrNYdQs4+HexgWbcoSH
4UrT0ut99HRGTtfNcwa508gtj4ite13n0IgeRhwwWkMj0NOQeMKq+YtRU2fQH093GFrh2c85CGcs
M/LuaA1RKqyRj6kbGOGarymBfbR6nNrTnD0YxwGduUZwylUs4DMRRZb79IIzbrMpd+xoo1ZXVb06
xEzCVUBKQTc6YUvYLlr3ehX9Ji9h5apjz+4MhDbVhHVw23GWVH63jtDRY7z0iKgGYLrC8eYDDmFR
6RXwFtUntNJK5R5r4sdx9kw7P0m4656t0wZBJrffSaHfslEVEfeg+VaH8G8bCPT0CbKDkaMp0YSa
j8T81dV3SOn+D7vnm2tBsZuejvCaDe91d/tuXRa02n385+1CWWI6GqwzIgotsBwmX7xbDFz6KCXN
sGBpk3jTg6JLZqI0JtkYyI5IUFlazD7TOyHVr0bzjfveCuP5if7eX2jvTc646rXyJ+PqvnfzoCcj
iWYrvqa/B6l+ZYKZLy2B3i1K2GdsV9O1H48j4dfgEekBwmVdyeSSYVx9LsnILYKv/380kaIvKEOl
/keQ01HzsWOME7WacrBQkeoIoXX/9GAnDYBtu+eg6YXrAF1U1hhJUTWNyTHmtVsYg0Ncrtas/u4m
+SX4O/Qzg+OE2IRj7fVhH7AOzIBYA7llEcu5LXlLLepvms+3Btk4DxhGNxdZwYUefRnRO5JlhRt+
jPKnq/MFLma5vLx/+4vL9duUPGd9dOoZIl+adshUvsh8cQWag82i+8lL6I+eFP5ljtR2gloTsb16
n82QvwOf2zf8vzVkFaiU6wQ/7Vq3Ygg/NfuPWyELARYjiGBOIJ8n0tCWyuxbZwa8DVNec+smksjZ
7s9WrjaTSuOKq5c81MjQqafM3/gXxmFFr8pJUCPvmR819UAYcQA+HG8UpvgDi/ZE9d1e7+nhCoyu
GCdpfMTeq0pjHPDcAt/Qy1tLXEsGYyffNAP2i7+gxiTVPWW/osr5xn+ZGolmjoEHBRiXKFDJCBCV
tonLNnUX0/WqfsauO5OawNX76sy7kBScnaua+o+Fu0LzD9SJahV7R32vw+p9zm2Lw4m/MO/KYZdO
kikm4cYNCzKJ7Ib4PhmJ6YO6VflZ88NTItu6eKLZUF9KdF7eU+45YWX2CahhGAKylGQTm9xNf2BB
tuqvxL0agg4kQOd0LntNW4vIwfYTDz6SkPi48NmrUN7j0kU8oOqGzze+ELQf4Bk1GiDoWIxZnd5c
41mJsWpoMMb7yHnGKCOebVoBWuhZ3kIBol034YP2EiFtV74LMyZE7zT7dLvFqF2AnAFBhXfCdh6D
lN/McWw//PSNUnWdCZfTIbNz6BB0LAJOLIsdFkquxhRM18u/tEZHZGFbCYQmLCNl+OgX2dD+igyU
weEu97qbumb14cl7RHbYXMKlXO9FCO50+yV1MOGPL9z0Cl3sf7piwS4+VMZMjZnAVdZB+86d/NV+
2H8HDWvdFQ9qwpYs299tNhw6kaSOMkfIOlIwqFJXaLbm1mlb/Uc+QJGaYLzccFs7Mr9m0srAgs9s
D1oJU+XEBfPKgQ1N9pBuOdFw85X6JpDvTL19FP9dH5YQVw/1zmvuKJUmtgQdFySCUP1/5yUkTpKg
SUDR2CfJB0lHeWdhWPA6Cj2IlCM+Sm2N8VUeQ7EvkNFQsZ4/zffKN1M7NXrQEaldgzLVjgpZ5cXB
o5C4UdKvUvQkbmMk1jCp3Fsk77vdFZNJ983zA7Z2oWD6BCey4F8EKloZIQmL0PAPcissPA0jqeOS
6XVzKX6zDW49xja69tq1TOnGk7O4CVre7qLGpjO0L/0wGerWm7CGUF2Q63eAo/ZSxtQEP5+eki1x
CO8ptuvsFjMfvDUDlF4YEjexk+zNzOtzm+ZvVId2egf7mxQ7VLTqXVwgRzjkSI0yDz7BlSJM6Sgj
gnm3VifE/HpKDR1BDG52idL0tZzR1QSN39qnUB5zOEzdhSwKTmqNkpHbG+eNW//omxEHdq/c5adi
vIZ07mia0V0tJf0/6c1GxMgSioDltcJqy3iMJLlt9OIqqH54u4TwOrd5sxkdZw6UQ9FbsohsQ8uT
NUKirCs61PHejug3snilyNk9h2M/j3bzL6jMPmW31cuRG7tskR2mHhEWOWIMQqMqF/pRuyktaLzX
fUymDX8Uc7KCMzDwFF6YDijDtNjccvb3+rqNmyX6rS7UQxtjyCLrOPCNhlL7x2PKrlJ/AQM3sIQM
hUWPlFG1CeDxxfWztsvU4bYDj6fHk4a3Xnqp7FTu2pSnIpRo38C+JgwhluRagGBHZFl+hNIxWSPn
Y5Wu3YXQt/PsMIVasa7Zpt1vtj6OgnHycLudOmb1ndAteT6eQk7U8wangE9uHXD+wBBWWR4cwe4r
zV3PRLoWO12EGZHT8Ya/BJrFSLFQCNofZ+oYOfG10nqimdBdB2jB/oaqF4gnyZQhrH+kbV4rPESX
Uwkrh8aoM4mZxSfrB22+DSKENEtGkZLHVI+x91C7gkDm++iav3Dar/pRLgIu7YVnEo1QFJx2tgcg
iByuQjRm9HGBFeUsmclmdICD/uxd0stKJb/2eGc7DlIfIRDs/vVcvO4aW1J+61sgk+9ApxVbHcZt
st5S5CHYFssIcGewN7guS+kwdlXtzs+0r7swjmRODGsyIhnIta3FbRxG22XMZVR3Ncj9qD2o03U/
H3tyDo0vQo+P1k9ewmnoBKeFjt2MhjGzEH8eBh56ZXRa+fNBOHsqj0dbBgKjdSr0xfUO5mAI3cyK
4K87Axdhh9xFSnnFjMy/rdxIVBRE3PNudzhbRDsFAc824cHzt/6Y5NbfsiW66NhJwHevoQjoyIIo
vPVlEnHrxwe7do8+S9DaYhXARNf0L+MYUHHu8WF/ojCT6pcRicQziGURXfgH0zl6lsrnvpawD4zQ
ChiM8ymB8cSDlo9ORcP8MKnY9p8KGt3Q9B33+3qWIp2Zvyw3WRa6SVFMHpNlGmjZ4ihelIG+hp5E
Rv8Wmq+zUuXkJuEMMSd3oCVQyGLLKGkJeHd/6KT0gYQDfMAxHf6E85oSEz/3hmwg9Bnrh2VdsJDq
35e9tzHfU406IL/xbwXGk3Y+a0bYIexR4siqa6MX2yuDqzTzKb1GJ1gaZm//GYJru1U5YXw89/Ad
zx0Ktj4rllvX9gK+XHTDpSm4bZzIBi7eXozRfCcnosfLeMsWei7T4TglAr4hp4GzMUMSw2s3dh6+
z6SGp6U2gdy/vsMebe5PhuIsLFGpRkW111YWbWXsKhR/orP5LKfbFOr1vkLs1qdFIBSMYzIqExhH
Q963tfv1z/B3B5Aiic3KNXsJOL9y6I3Qih5HiOqcKn5WBcUT93qzKO+vGe/E9WWHlIqhFGpSwBni
YK1NJzbXKgGmXxpx83kZGLuAXjkMTCuPJ+ibACJRx2k+SLaMurtJG4SQnIGZuGqhrp9JE9zaPFAl
77JX1iPNrRrisunnyfEw57umEi7AC9wHodndBsJESrB6YJtxuOLSkG2CCiw9VKtrWBnZo7BxBd4C
PKsHD9X6ZauhF90s0FYhmYMYujg7/Mk7KZTL7LMQ+hSt0PI1bS19SRJd1i7dejFYOWfIA+9UDV7e
tigD6cWV8bbBCdyNtrsxbBmG3gUgqzKF0z6PtkVwb9uQoVG4Rc5kIjTysiOhOFYF5jWXPgILPiUm
jaaj2eeu3oiKG78ehDHiLB1iIkhOUr0nHBtMA4N2mKEq2BuNulSmC2EfOCaK42pqdYNc3uzLsHT7
cAz1bCSSB6gBJfgPgMxs+3L6GGDNe3h5oy1PoDSDnrbFZoaiC9XIQiQ7z/Wuo35C+GPcVeZO3KSV
AhI/2O7Z+IWCTaCQKLO3EHXAKBdZnP3exA6movI5+HfdTlnxhgW+/boBi5oCJT2PwZayfqD47OVS
EmjuuO6Qavz4f6Hi+W1A0d4Cnd4cpQVEE+YRjJmC/r2Q+A7s6Kjst4Vi4xDUNg57+hT2oU1ON59+
RzM0g921fJma5prlsFD9M5bLUqMITHYyoLAFj/LBv/q7poHPfpONRXxjDciLObedxCnEeeJJ+kbe
sG9gjoE/XzRPBTw4OEK46HrWdB2Z1zZQw2KihFbIcCUiGJvercWgkIa8+GRVm4xKXkHAZUenMBSv
61dZ1pvxlHn7g0rvZepe2bxsVQGeeP9jFaSMddnUU/pOcKNFRFH48QnZJ2wbFJhiw+1Nm/f0gxuW
tDbeMfwz4iOaCmWiDX0+oKDW0sl1W2rKS32Ub5aQfqN5AQNyCioDmi10bImbePHDoNWbQxys1KqK
VsStX4OWT4KTDzYZbqv/NBvr0PbVeA8E/GQPDZr+eaJRr0ja9hPo9gxLta03L4v0oTRBttKlTjXe
zjIyJ821cS+WXcevjLu2a6t+A0yS8nHpvWH6/7UAsF4WTBvIrE3MkyfP/ojxptwDbfOrI6LeXINS
TyO/1ARX348xQ4KwAXDaTVnb+iBHVV4OkpfDHtYbSbmCJh1a7TFC+fcPKAKgn3cal7DEl5xSDGsG
xDsGcxpYATIziVOR1W/v5w1v1Db7Z50Nrqmb25jqZpuJvc7yGMurKYwUq958o3HNmLar4yseJ6ZM
fBYSYW125h1+ROVtPAPI5uJYopt524ewI2D6/R5tS12pPXdkvtPGPbpOqMpXu48hCjeCQoC3/q8w
rV0YxOxYeF7TDzfL08/me+D62rFmCpzL5NKrwiKYilGgniJg1DDvp95D0Ort0kHcD/FyNCa5luq+
OgLYGqVuRWJNsr2n94FCQaRCGR8Ybs2vMn9wrlsGlzNj6AVPXtlShjip2Jstk7heZis/dmUekr1V
m9rvxElV7ctNK9SKWl+6tcDq2/rlafyn+C760UaoDoFU8Lkw+Zu6Zd7a96wxizIJmNJNJ3ELjX5u
GgMmCLC48kN6wumWlJpf8ccB4YupmsB4NdScmLQDEMqshfGs3n1ybuslzNjPrchlhUtzi4Bwyr2o
8lLpb5e9gT4Pq+id9KtW2BqOAtRUfsYHD2FvnGW1OaDPB1o+qBIrGVcq/+DKt+/PNAyWGOTQ71Qw
/PjZcKdmI+gIeabmYSf4u8nUEyRGRD5kzQBMmB85eomp+AmSuR+N17v87Y7YkXrzR5QIWgDjgZ7P
dLvEevMyMOsQOpjL6gLNCP5u8CbRMNocboBcJ7az6hFHUt9BI7fWqFK6RudKFNTDQvdkfa/hzSD0
44AGX3t0ce+ph+rM41HfHVkhdZRZQamC36MIKZF+DKf5PeDq4yJ2yqkRLQhzdsNUDBq+P1O6GfVo
jxtcbwu0Mx30BzPhh6OngJYRzzAgFQV241LzmUsXp5LDhpzfWzZTJhkXur1BdV9pv3K+OYiCVel4
tiQqtmUMAU86f0ioP67a5/SzFVDvUK+ZkMomgXGCvw6harT2mON9R/FjIC/TgLV9orIVBnRmY0cm
EH8LD5YHKORj3XsTb2/O0gPaIuf9hOhhUb72phXiBQgF6FbAusnYSBd+L86Q8bIhTPvI4wx3dn6L
1zBfxrmRKC4sKSIzpORg60UC5tbYPJ71O1kM60OvVpU7rKVp2vIr6nWCqAPxvkoRj0xtTvsnQ6dU
rDjjdZv7t99U7mVXsYUEDO41mv9KtI5Z2Ozxph+31K6qSgDi6xsdzpZvmplXc8rje5jAyRka+T1l
lAjr27PKgv7fZK2IougZYAOJN6p0+uoGgP2+jqgl6QZ5rZIzpGxhZQgr3pN1AGc/gToTNWpSzO6w
YlUIB8E8oUImTC6npePAoTsxCH6YT5b85IDJ6up0bwwALzLvx1CRz/GCoztqmOEE7ZiJcLoHhYfT
/drGd/3tOzde7S2CMwS5HTQF1/kQSdxsT54bq646R03babuR2HQf3ue3Z1j4jfnUzMW0W7Ktm7Zo
zGcNKWEIjBmi+aDCHXbdLAkjxXHoO4YYg5oN45agTZuI/UkcAUQSXvj15zxfntpC+q+htr/pf+vl
63BfaD4eD779uNBKImdMrY1plPQ4cgCV/Ps+gpf0N8uakdxRlkeZYD19cPENycF/uUEkhM5cUDl6
Hlo3ag5O7oe9KtQ/HynUIZfVBBl7ss2TY5dMuK1V1g/ZEkBGopzNUz3o57w33kJ2fMkoQR47bPFz
P85K8qz9oaKe4o0fZB/R0t1IwjNbgMm9q6jpeWYwePdKPquDXpv7Q760RDmS5eMI7x7DxkA8QNGc
geEK9c5tof23wLSltD/rSPBbqoBayvab2GmkDIreKEqX6wGRMDTIqFxnMApeNl4GVhrN5UI5gbzD
brvGLQIq+kB5eN+rNVAB1gwAk9ygO8ApZupSOIToWZAiIVux7X1KpBx9hUIW98x7IvPu+PJh82j/
vgdPfAb2PV2CysPkoPxjXU292cFkLOv/pdYJhQCmOcGD736ckQCFWhV8ulEsuQY5vqU+uyaK3ioi
RY+7Js62bTejI3SrLXhpjvKqbO6STMReF+c1HIdV85KKG8drvhZYMXQN9GCxaBEzWgHuapIyw7VY
SEd0grYvpRq3RRpuHKgXOkXPJehrlGARPyFiBDoDr2JJ7a/jYHXy2/OxVv3b8tAU8Y0YB7rhWFDQ
BGFArGDYmzreA0fRFDMlc7jHIA89WxYh2+ZA0lVZoZRfpGhqcJo2M72k+npgWl35GwO3JzNSJsXq
sOgKMjegIJhhJzU3d7uB+9ZGyIt5bK924Zt/lfIYc/I48L9t2zqn6Fwlz/5aPoFPIbtnxCtM7RRv
461rbsDE9Pl0GMAWpAGMPDxzHU34sTgAPjtVLhc+2dXwMFa9wfJs+PbQ5HQ+ZROrQLATUKFzzMWr
/FH5DdszoAOpLqK8OcUBlgB0QNfMPMcIToPRvQdJP3nUCBmp2cI8AVm7SnP95JPa4jgIRho2DxJu
/CMOHVooz3e6TC7nX2NCR6h+ZuijrJE8ichYGJbskx4Z5lCycycZKY//G2xpH7l11bvFiNGQsHyv
d1haDd9jmjImL34FNdysWJgEpuwLY+vlxbu4EkdJrfZhiVGFpH2pBQNdflFUeRhzjYC8map8g7Mh
CcwmEmxfShrARpTEz0tmi4QAN5VfuQQ/AGd+zjPris3R1DhXLrGMvuTar4ETBFFU6Aw/WBOe6o8w
WxlwOcmYjTExuLeLqQvbZxViQytq58i/ntzYJeo+5SmaZWHRvXBrn7AoXKIgI4gMBSGq5iG/inQm
Q3Td5hrUjoclxNrpzuU4VlxmEyI9PsgLAeW5pxDrzBj1S1XuWVPyDOLbP+YcigcOq+rAMe33YmEo
iU30ghpoCUvGP8C0mbCWdEaJ/GrIqHFc3ITKi1rKd3bZofTz4i1Pr8NOHHGUU0turJotyvV0m5Fq
OGUnZfPeMMXFGow1oIuInnAsTXeKmhqq57zticrtzbJFOooN1hjn1fYND/m2C9mqkPGCqxndJ92I
0M/lW7cZNKvzfGn+3YXXLpSOaqPIfBKevZNVrkVXDAO1+rDEtsA6uoVFn0Snd2urraDWIiNqafYD
TwY3OvzoHrjxSpjNWo8xNXUDpuoU/FYGi9V7NActiPjRvnu86qlvklCrMhsWAOhHHsJm8Pbc4u+a
K76Gedku36d/OuxtZUMIebbokcOxjFgDiqSuliwRaqRReNS/SEQ411cqzh9u1677CeoAb9Af6SRk
nGEIg+MeWbMlPjvN3mlZpyYqYla/VASpu/JgIufU9KSg9uiSZiLP4gOZ2emQPiadgG0LgMV+jILu
XvCk8FTDA+Ll2xJMg1OFq1x5OzERlvIAXXyucjLKUx6AUJfuha47SK8unUY6LN6PRH3AY2prgMhq
uy26XdoDzWhT1x/oP3eQ3+E1NjnCNUnnPAzncVEDXLMTUVFh8jeULXsOux6nBVe+ZgUVQqzV1/Di
QkelhW1/VpCT+BrObvQYxa4CxLaC6d9ICKezSVcObeeov0vJZS0q9HNWpT0lkgYoshK5fa7DcWnu
fm9x/SCddjeIl5SuNW+brKJngyvOhx1QWGvVjEwAC/TtbfJCV2iNMp7kbVnIj3acVC/EHyoXkbM/
Fi6p5AUJUGmWWraxS5bkeoh1br+2mpLNhPRSlmJZX8UwvaonSvHkQkTV6s3PzVQ2HMlrR6RIo4zQ
ZhFaaACceJpAK74XKpPD5p/Lwm6QZ6WPCB5jk2in2wiIClp748mIaAdFhV/BO0iYNkBuZMSvGeIX
lz+E7g/y2VMZbUOrzcWYz+dlIPybrEEQ8JnLwvmp7gLS2yugbAjEt9al4oId6c4xQ6LWU0tqdsHf
a8RH1xTRQMdvZtjtkQLp2bQmVpZ6pcqArIpctPPoJiR+TTKXVJnq2w+i+MPA9CIAd+5atNZ3Wbtr
zL6MxsAIZjhZWskFvUjnMnC/TQ4bix339nJJ5nAJZp3t+VjXsDIv5eelIT4P0fqAatnPmMtBMSrg
xQ3vjrLBt0X2z0oI6hIswRhzQL2XMGmDV/iDokLZBoPuyCvYlQdOvca6rmTMcT6+gaaBmW5aYAEI
BILVU8EMLHZ71eg1whdQKQtbKD2RaIHORColX+eL09AxKHb2+A+wXwe8dxvai+SpDB1iu0oz10Bl
0T1CT1euQp2B0VNVWgshgG+zYm4P/5VQF0HqbU+YBJwIOi5ATk6A+SXmqFDooX1Ynnyx3hmMmDYt
6IS42CG0vE2r87XZtuyESl/FKOyibWSRAuVZwJwzj8gB/DcEAAGfeScI3yQaRjy2LtgjWscC/uUA
uuie+ULi6PMGl0kZjXR5NP5huBl5qI+8Hfi/lvC+U/LTG0buIi++omRqVGSD39herfDmYVKh0H9z
xwpThcvma7HspQKMPgjK0oCNvFkyakuFXCYpfBeZPSduDh7OKc9FVugC1mvm15JmOpxdSeyJORWi
tUi5MBW4a2YCiuKY9EHIc0Cra18VoEa1B0cXmh6qQEPji52fkdtG9aNCdSvSsjol2doSweBJLZHL
u9a0SrO5G1FSMtvWT/BdTZhcjfZyv56FG2detMWnUFecnzBHWYa363iCJ+/RDYutk1dv/v1n78VO
758LKGp3AkFJTN0ChxhhIJn4kAznjUWAObJmy1uDhlYQALykwcj1Vo9WL3Y3lME7EVUtsDBz/8wk
so3YkWB2viHNHNnwKBVST4XPO1iZU3J6VlSYSFtdZzTo23fFae0MBAvQdjzlLKEAJu1WFbdqdH7Q
xR1l3S88NdcVLAhMKqMwPwZMLBCAdXYUy/4oT+N9kJ6J4is/U4p+d9TdWUDSdDmLdHufJiOFNrbM
gUTkQjeHbJWK0WpFgm/XXxs2IqEKDdIvtKmJLNUkUdkwssPpc9fqNiKTsee9GCxWmeBTg8tvUKKF
YPNtFPf7dw0KqlDPeT6Cc5PM24/udJHORPgigrTz5p0Pyh/mc1w6FhfQ+sYEtIWUV0hIYNsl6WHM
8qJDd/V2KLxX+TDV2xMyGXXwGxhxvBgSPP8YUJVoQEb2d99/4V5U61We4Yf6ydfDZOB4F7M293zU
cyD2Z32qWnisZL9o0Ho9KnyopVMqYT0StXjapOvD8Ez6T8Ua1xskoiOp/DIweoU8u/a7T0GhcQp7
XxUOiOxMuRfkYr/z0cuz+m+hsVNVkTPlOzh+An7uZznUG2FlXaf2ev5cE54ID4am5Pilw0N5XFqY
1VqPpPs3xSaSj9YbXnCSbekrQrza3Wa0aIOYTkKpW8bKO6HgA3D/Aj184D4BMAtuAe4nk08JvOd1
KMmDg6c+MJHgcmecXVyfr/84LF2MnJL1F77HSNVjXYs1CRfrU9XjLzkutGahireok1KOSnaaRfnB
K5t5xzLiY2K1/EHEietv5iUDLzhwkgX/AtF8FC+wxrxbaMnOeTVx7bJ05XAm8xxMYyURzWJaJhnN
7702O5DianRqI4sOq08UnlOtY68gH2rNsXVyU+tOWbY7VkCuwEnOwS2Hn0kZjiB5OrRjYPrDcYf9
nawIhChp1r3Kis3n2VEh9FprwhYPWW++s264v2X5+EAQD1nmp0eDHkWMJhMoHuffAl2pO2oDUch6
oM5wchKlCEqEpyQe6I/BAwpZYvNP6WuSQaZ2ofXkuJGhKTCiRxDUVQWDGtc1peUQuS+PCUvhSLSL
zno+fvi3MdP7msOnXaMvIQFr1ah3sIYziyXTsgLERJ4dl7iyQ6A9UkKNr591wXTKn9raIH8exW0M
q9qhkoa5sYeH09k8dd874resnDoi6ICCMDUrBvo36xB/mYmbBKANQAbrWbmMzUGO+cfPH/oHDb5I
vcXCKFWQIBOzL2iakQh0xQhq/LFDAihzT307PHClBZn08FLgP9Rkvkkk637NedlVW0sWXHukYa6H
jSMhaFqqUbin7I4Il8xRpgijiNBmGorPHU3XlgQsyXmkKeYem6MA1lJ/G7XEqe0ZXouJlozgr4mv
p3rEyuO9z3Zf0BBDkQ2GlcHSs15RnOa1b3EwcSeysf4tMmw/OWcW9xvy1QkAOS6j45rl6+UuxGue
x8m4L1Tbj2wowazO6Zw1hhPDKfFBACvmyEczyV1f2N+LS/hNiVKkWhEe+YMvqIz9MwYXK6IAAM5d
NIx+TwlBGQPLJf3TrnvkfufUJXf9gAc1bWxEM5uGGNpCUQTh7HW4Jjm2ZXvyVHlia1i7t49CVFNY
9+hZXIRMQ8E3ynQrFe/T8DoOyBiAPmaFhP68WY2xi+ZxWNZi1wTi6yHSnX/wHpn781pkKCfPszvj
vKDarhfLzsSM882aNyXPBQIZNvV/CXu9P+/6jmTDAH1bIGjexqB3LpcgWbWY34ZL/FTZq2SoRZ8d
xXaZzQ3eazaYSxf89vynI/iS59obSrDsqppIMESBFJNO9tKfjZXHOtzYvdUphubG1FEgQIoSvn6e
VqqUKHhbDv70RfIjVC3KoPEKda7sYRHwTCBq0xPAdPsYtfLKW+pGa2Jo27dXmZ1Jh1yYl0qbVoZB
P8xtQINjaOnxBVoAg4pgx9y3QnYRk3mOv9J+5INFoM135ZMDQJ8E5Wh8sZ7m3rCx3QwmuEDVor1e
8oKsjpiM0U1M+xd/HLWDdnPPiz1OtWk5W29BSCMMuygKH5+ylLRKWi6YcG67y4ENEf8jE3NVm3c1
JC1VTVwWYyxl3j9c6lZduLb4YTLJaUZkmmPd4HAkcZpgSEMDboA0o3yYTZxDtlr4fCQXZFoszTyx
2lwYS/FTVzT2VVGiwI1k6b9pIgKPr+KG3VqUHUZqSOAtrCCIk0Z8i2b0OVjoK1vM/KQwRj7aZUcj
I/SOiRO4ugxt713VOz3fteAXZbpCbs3boc/Db0UrR3dk9bjIOyI0kDHqlJOnCpa3XzvvCZlbV4nJ
aiDWcttK1r1B6m0HPW0ObXzIFOtYbx8M+sNPx1Ze6KlPym31nIszl1jePz445Q8F0tVISFq4X9+K
MgJg9SY4Pq4T3WvjvPGc27HqZOKM69L4Zad81/9Py/BQQh86f5le5GSdSbbj224ylssdwEyNZjMt
fcrgI7B8oFqAFhORYjO7vlsHUqQoYA9ghznJm7tG3Kq1tWKfSu8xw86dgut6ZQhl6jUjWqLKZsWJ
TPExHnfnM0iFSJixmoVhGSctAdg7QTYg0YFldThhmBubRif45AK73mnfOHBCH2XiRAVk/ZtGR0Y9
TJwO8N4t52Bj9sQpNjUL0vHB9So0Jcgm7lT2p/4PatV9pVWgBz7DygD5kweHOrgIvlGTWZSgQa2o
aTeAv11JRWikDGtXln0R3nZztzQSdu4k4lDobxTOgJC8UQet6mY1fsdwfe8PsDJ/q4Mddlqq8e0G
a9brpewp3uJFS4QpQ/c8rFSI9uYRYqEqYM5xyOEt8ihPceuJaN8iQF2Vkz+iVVQyQL6WrYv0wekV
UMKXFi6xTk/fIbvEtRCRD8noVAQ6lQyscMDbdfRIIw1Errk+cqq8DQIoCQpROfXHu+aUTVd6Dq63
bJTp4vAY32jZhDURXB6yXl1AlBUujkGjQCIOjvZTcLLN8cBT0GmingoiazUQKjnkl10u8mAlfIxz
dtA8/EbV58Tc23TRm0sCKgFpZwQB3EY2uJSrqgn0rUhuBc3saLFH8l1lf7XpdAWzKyBQNlT5TyOZ
/8EZwy4eMDRNDXgSF0NTu4BtwHnvFF0kK3aO9ONnqWlvKyDuT1gH5ZzmU57l2xOy1XjunAiIOWMk
M5G7ZatL6B0LSo9ES6ZGPd/tAnae9FScz4bEionVWLkgQZaFsbQYEi6Sq4ts0ZeydytQGb1VtRut
1Wd3dAzC8rjZZMXKytlhrmCaflkaCN8o744b8M4Gd9857aPU+DADQHWRlCQ5bJWDLBUP2BzHHjMl
BKutil3d62jGNjU+V0ri2J4oi5fqKuEDZWAbq3kJPPhu6v0jBrB38AF5lPeChNxExOaJ/zWxjis7
HGO/DHUGmkw/hdsCaS2odZ2aXKhxdXONm0ekKyXY9nAZGsySRIJxGxzpkeabJSx8oPnwEGrVTQMU
Bd7Fl0YD6gAdTp/MkxRR4HnIgxE7KHaiVaCbI+JOfT2KspwsVCYOAuYqjPQpRcL4a3a8D6kj3VSN
+iBMJxpVJJNmu1yMT2zOI/TMYJyaTdZLM331xEccQDm3M3l9YhSbESKOS4UwzfDQkNCdAt8H2CSf
iiewZm9fTkkKXeimRXXf1D95KbAkMLErmOhZ6LVjgd43WvL3b1cs4/d8w2xqW+COmobxecKteda0
1rdaZsakFWmHqnyroeXHPDe6hGljW1TEJ7jrqZXl6z0+jFNZFOPwd4d+0bj85DrCKufAZYuwvegm
FpEdTg8dn36ofgYTNfl27K9/eVujGKpw8yxIscYTzhCyE4WhfgL7Wnr2y8cyYY15UZyKLbq0L/Re
4inz6Kgm3WZsW4kKlypGpB/6p5uyxubPb+TZWSVQzWri+4tOYIKftHwjG2kKhOSDEkPIaJYY/RdZ
q4GnzuiYin+E2l3DBMuQjRnmk430ggxUmXVAVst6r4Ucp4/mgoi3/y2qWqu7IJh8S+/PqtPzz89w
y0W0hrY07G/KvPEpNIP4UiYwP58kbumE+h8ERqUvHxejoBRTkapmufxuyP66EEEYsJrURU850dhn
OXpZbjoK+KTLWpuJm3DZa+lrqPtQDf+ngk/gc9ORKGBuUl9a4XHQVqM4mC99+en+jCv2p4/nCPEK
xkhaeolC6REAtyesNmcsHNI75wa+ITjhcBkcevNy07GaggwkBSAlSu89K5mWpCPeHK9cBmpbANwk
5OD2MqTTnJgIZJ2BwPd3Xx72IOsJN4ah082Y75j9f6Cx1sgt5RLGfk6iQMqXIS7wi+eoX1FYVrwK
RkAX5gRWw2lC/7A6EMohVIo9Y2omSpO6n63zyCiFNKwpql5cGBH/xdLzJV3VT8HK5eVhZTGbuIOv
+WE8rm4J5HjOxQenfaZPfI6ARi1HP/2tybBaNPdwG0ZjwrrznowpNBOwtK4pG8Z0j6bn8BFuDdW0
r9zzKjFJyZK0fgA0wwBbZ3Atu7IHjFRbu0zrdb1HHgO7tAF2FxvzMKX7zJZ89uQdG1VSRnETZYUA
RWccyZoEB/N6GfRi0ZtJ62HfTNlm3Zf38T6GIIwEo3ytkv27pQqKdcGo4NAf/itMlYzyG9r/4+vs
M5P8ZX+V4kAi7iAbQxL6P8Ohyv21Q/0gi4ELTY0249oAw71I7S0HIMrgwYg+vRy+An84EP6oVJN7
CEX3GB6F6J9TpIeMF4OyDFn0HK0QG2+nhFQL0Oe/SHnvZGPJuNBvPyK9lwX7C6tj6XGUhwXvaq1A
2IzH2gwToI3QvlCWhJ3RpHWP1Mo8AORAOv5rJ0S8KQVLzYz1AK56W5fWD5BM6TIpYORps74HgK6x
4J9JTOVS+TWTR762qgbd7txMbMqvEkjC+FLB+F2vr/s+nLPCr0v4I2ZzDcCbdx6vgaPODlzgA8A8
OzByHnQTomeLIQux8D6JMQDM8xLojCPNPAZIeyfe/KVGUpjJKuZWtjNmaLP7VdLsNMjFZvfm4OWj
z866DHiNF6pq2jn+gXYbcRB5kS4TvPXOPcUfnVBskLn8jovY4GmoO0Sp3HaIMJhrrQixKUc1Vp7J
y6oTE+aLqva4tF99WKJGcztPBIM81j/uuaCgjC1al2g4pCrznWQiNezJU2G/u26gOqpmBSn7Honh
cRx97aBmp29gteoAJrvPp7ozSo/ccKMoV9+zFucukcLsiCeBb1dHQzB7Z1JivxgrkeWYLBKVBzaa
pnakG1x3NRZDr4fWZxDwulr38+o9c7AMAL1ur7+8cBoIsmcQf6asL4mTt0DUjkmhyWuRh+rIFv1K
eZG4LvnRzk0rpWtGRnFSSD4wsKd1+CkWyWRlxtNzHmt4qR6zO7qtqicSl0h+9NZ3YY8aV34YGyIa
1NY3kU7xJxZ3x7M6cCjHKGKRXjzYh/xHHFSBMibccrc4fEU8+55fKDn2UlMKPtAhW/gjeDHmqsEi
7lVEOaliH0vNY+1EHFZrja3WbrtAgUfhxpsZ6j92U7Y18g6zsdw+ExOH5uhzQqJPfbL+VL1Jfgux
jFCBuyUF7jiIgQIExKgaaP7B5t9Z0EZ548UGQ6cQoozFlYqhJjuElCzkofCna72JO8dPQKGCNSwJ
q/ntQN7LKS2kao6JfvshkUCnRvsA/pqZBcKgLwuR4bBKp9eXHfqwxbZMj1kqocI7mGMzHR/2xbgX
O2HFvvPa1pAEP6BBLJlJ08y25PxjUp2yssQBbktanvp2NrBEHSrx78fIh/gojZTGJjSynWTbapB0
6uePDGjaKVwAtI8OFmVWI8c7uu93r++tRrQgPrNgZDfKrbDlhNukXNPaUIuIto/5apSrEkdxjGCV
Emca3Efc5r4ne9JNbk7HiDWE3BpM3XYYhGSjtmQgsPd2gDq+m0D4s8M7xPx8PMuw32DNAFRnitsB
oq6/oTP7+SnR4KqFsahWJyiSLkK/N8/ysttFSzh+39LmxCXx34O4ei1WeWuXn6RsripTUAtYEUzz
6/64rBy5I//E/vp9U0lSOBmlMpL2HsqISTwamPKsUTz+1e0mqPILYcKyj0Fa4vZZHEZpRY64gH5Y
jWAIF/vCJHD2ghzPm14pzo2Q5TJIyEWcXe4mIMkF8eajtnPChGuTUfm4vXKoIvu/Xc6uh3v8j7rm
+E2SaDvYzWqIpU3+lmHJwyyQfnb1/LzG/CyCdF+jkprGmn1nbU6Diwhy2ZVqGICQ6TxOTvP54gP9
vML5WMJG2/U4uVAz0SFXGYzdUxIeeXXTQoQzq8G5GIFBmCBz8hw8qWxai9oth5I8BnbKoesKYP9B
SJlpl55AQFYZiHsmXvwDG2z/199Cdl0J+NH4GTqyyp+73jEkH+dWbeJlJM++W2b0JBsGuzRCQf9b
90rVDg7ck2sBwW9kWhXRlK9vvctPPpvfmCFz58NWmv6FMMWihc98H5vcSVQFPqa7bnjw+RP4q9oN
cyokDbwRPydiwWcEqsvjtIwA+2lpqapKsEbkql52Pw0lBNBnKxyCIuDb9S8ZaHsItSzlH6LgFkG2
2OFQgAII90jeHAGM+ZmhKD8Jx7FXilGMyOyl9IIsRdg2DfOwgxK87EdhHwcOLGYf66XL4Q211Yo5
/TMg9oxKajER5xDZ7w8iJ+uHbKNBGyR+F2ZU3hTlG29oaOReCmRzXgpdVoPWbRJUw3GF3mkbGrZT
nKZiYeJ9oM36gnyqsy5IfP5t2FixfjjLS+mjhb1m0antlJZRENlnYMQpHssMR/1TkU7yO4Hy90BN
sx3SELPgZRclAoyJQoXP524ZR2ScyhcdQ/Q4RnjXwReJdeijOXPb5RT7TcfpQzOY7BBoHeLH2O8r
jJ20ezaqfb5SOsKbPcgh0D5cm8HFHjsTif4Jmr86qsIkCgGUP8U9pdXKiGuPOlhzlFa2P78vgg77
UgbZRHrA7lI8lC9W0qR0cnmIF45xexCNmdiJhElKtph1lcRkN3y4tlcTSnJLCyxdUIhfuPKtP0Dz
L+DeeiTI2xdB9ISFfkNfXkbn6l3mcvvN+HNtZRcuLa6OJBK3sPZiQXR0ojbpQbrs85sLRNLqtEoE
Uh0KmWx/ATR3TdPHAB6vI1w3Nz7MQZV6ay1HnaoQRKWpASl0VCVVY191wvT7IWrBq5wymuos7KQi
40ZnMVSYRfY54YxcWQhssnsm1bgIq0VJLf+zp11iR77djxPye8WtYJpLJdBJZM2Z61ROOhsT6fst
BO4GYpKmc8foDT4z11Jr/9udBYhDQK0v3W8n7goHUeAP9K89Qk2uBi6lAzrveaBgKeLQu+LkPpkz
CDdMXHeN6D4TothxZRm0FNQwo4kZSJtB+hr/8GCltAC/xlyAXOzbXqSAr4jtpVffPd04OiXAlPi9
og46ETCXaiayFx0vSb4wJrBsFrf2RU5efNJq1WT4oeDZBEPYhUrxwZ/znKQj94YMpyuD9Mve/VHA
aBRI/Pax4ocRFH3e8QAsgcPgyWWZZCthDpM3OL8Y5WXLTicoBFToZCklKTLDu6Di4FhXFwhLuJTB
xQOC/w/0BH0YmE5HFxw1HGFpxlouoRn2+7NFhuOewqCAKrHx1bi9sRDbNrdRFWhCFAOGtzsmw4ez
7VXmX9Jkv4gQBw1ndLLtjx+wCOksnXWK0cOwI2UjSm4Kh5xHjrNUkMGWEM7cs5aO9Y+RdwcQXcdG
JXF0eS37P1FNqujPUb10ZxR/tsT3+iuJkFaCOCGGsa0JkK4S2t0gSf5/cBZCxImWPZB/ex3szyJj
m+C3e6WtoVItgwlfv8unNAxyBuwjOuoljs5/Gzk0TZTHAGe+xXp4iwqmQLS8VIXJuYOMJ0GrK7Tk
vRZubNYcrarA2wrAkqWicuBI0PKHdTImn6NqQ0F8VEbCx6K2tZU75KfnZPOkr+xAt9tjBM9DKpRN
SxmqEynFWxoSNnRLGb4UxsUUSY5n8CY5CASzjl1A4jq76CoCb9shXS1XE/7Soa8Jn/+HjnvMtIN9
g3hDDq1hGRp3OukGO+TwTiaISkUJ4QISU1qVQiHNXVgT4GfbFsZPM0V3ftftE1KhXP/hszk/6GGL
zSX1bDYhGPXA469ikHWyI7qSXkclQUb1tw7e1FH9m8+vz0Qt2mWqpIMLCKRhSmHAL0EJHy2eg8H+
N+jtsHpmAbsK4VeEa6crEpjtHV/ZpPTg1HwafpuItcAY/nwM2LiP71DxKxLPZNW5eRXeo9so6diH
Tgi7yaFabV4W+9qjXLSxVPSwUU/N4yzws9+kfQ3qu9JL5AfJ0jPSDRsa4+enehMMuGg9q/Y3qbKS
Cta8JEgPNdDlFNt9ggos9mAFyfxLA/4MzTCGT0IcX9pwVy+IjeQTj28sBDSu1eh0D3GR7RUPQOn4
cIXxP4cyAuq33YCbn5n8zNZDpeftFhBq9oeI9sqAxivq4FLl55mtyY1ZqyQnYl82TZfAOigk073l
OzhLQGSQ7Tpycw3OQ7czsZc2HvAXO0zuIOF4U2ySWERHY4eFy8VXLqdlm1ZfvRmp8FDEigssqta1
ItcGB81E9AGnEVFmVfQl3r520xTamqcOuNkQTC3ISVDWlcKJ1+Hv4LSgSRv69yttqa0Qu/wN98Hd
2VSDfm2xJ5vtzSybA14LZF2y85U4+6KwXaU+h8+EVr2aRtHO3KT8l2WHvz3QJzZ7lwgIgrEvYy4M
uOEH216NOfmcI5D+mXH6bLa0zidPF3nTciezMdmxgxdXEWn01dt7EJBbIZ/5/ZcaWPxwTlUDCoR1
s4kBpENjzAbvv4TKooqMBU5CB7Fiql61Jc8blW4CBj6ajjzWGOOd9K9Ung0cbtpdYEo3WcsW+lHE
FhazEeyFGFhaslPWHHgWCZp5PActXuR2IONk0bG8d6bpd2hTKBjVZXWPkmLL2/qsnOMeIReGA++1
MKXbmb5wckyBnLjk16bMbhP+zQ5nYwDKczMIDKhoTMFKgc75YnI3GXzZyVBhZltb1awtpECyHBe3
AuCuylJ4z8Je3CV8zcV9RUG/zJ37ubkJ/8erltrhOzwoFpJg01rZuBvux3aONvJQcH6+BjC14MRd
xMKlFTRnh2HYmV0ogevQBX1xBGH3ym3nrkeiG1GR2ykjReQzW9lTq4zz3ItUMt8vwESyBkqalcl9
GIXwqPk1ncsGb0jm08fj8mAU1Kg4r5HyjFGJJ1U0D507SQPaJvq3iG+RZQZY2z3jGSbFWK+5ZZFW
8lA1XcNG2+m2/JRzsdS97U4oOwG+EQqBFXUBr91GcY384f9pXGKZvnHsomsHglnKWp3/v2Rz+QhN
5Uj/f0wwQYd9xABvsZcr56mSncqLlEQrVUyHiCu4icVAFH37oT6U7d7VayLYuCKE41aKV42LCUQ0
HXpMYLA3OIc7FIH73PFWAqgF/IsKtFQIlGoMzjtSYph++JESTtMSQmyLwqZ7fHV1F768HNOZwdPJ
mYmtNaA3Lopl9ztyLtjw2IlrdehWT0TeBeBaMU8bhZXVRIaPLe+VLG+gjBeG4sQdt767GBk5MVHy
SuV1Ff4iw4VuqwHDQkC2qIzKrKe3A1jx+h3IcC267NsyS0lkuEZuGFe6nWMgnavB0yBi6z6k4OtW
9PTEKPNRI5Bqe9pEYsJ+Oh25+QqWJNKKy4R2GCR5UFIuGWt6D9d68K2VKTOfjnFaTTRZLGq4a0R2
vnhEtWQD4zsBFldvzSJd9+E/naea3BFUKpnIbygNkrqTsWsIPIdv2yjdfOVly2SiX0EztnJlgFRx
6cKzlfQ+xaD5pJnAuJUnsk1/KAoBnyh/o2p3S4vxgx6+UBpbjttbFrZpLSmvYJooMebVLgkMqUgk
UOBVHmQKSxEL2Pz001FE26xzh3wvwpyrNkmxZbvxAXBU9xVCT5czcobW5OBBikhK6c1h9HvHG1up
pn7NgXsR0XaIG5KLhLRVgzR4Nlkg08j+yPQp3il1Qwlka9LaZh3tYweiCqK1OeiEaAhSjFyu3jvY
kLOQpAiZ0Y7Q2p+znfjgEqQFWIQqDo+rYtMOVZdvkBRPi4TdrRSTW+fh9pvOb7BN3p9VW4k659S8
IXUCbZGHGbXyD3b5MrLICjL5nTht/Upuo7Xrm4eRq/CzfJ2tP014jMZ/VC//+7ZaPjLLkt1FKr7m
IdkLRq+uyl9nP6gS62GZ2OhYA5hOYGJ2vfAxb+1teDarBigKFgv9b2VZbyoYyFx5pr0rYnhQ36Q8
aVDkNnrZEXuntoXXH0SE5n0NPCYXlcyD5IJlRdoRQ8H7OGqDJ2HmCTwbRPi5N6powByV37USv0b2
AsGzu/Qepdw7roFG3NZm0YuSBdPXrNOicnEIRbF8qrpe6hypEb267iITgsH/lj6bdRtF0AlmitV5
KlHUpD5rozMoH5vwg1unJ4fKPpimDBAsveQO9oG2OcyfplR0bllm/LfVzATeovNFcVID+ftM41rp
bQCNiY8bjdrPCeYPRTmr+cJk9v3xsrZzem7+12tA0YMtW3+2KEoo3B3+rM7KJNQAw2O4VuWNk4SR
SoPz3jXl4ZRQe9WsUBUS5oOBpJjVtjTkXlt663RwncaJz4Tdv/m8bhCmMcwayFCoXpq9+sPmWGD+
da3TTx3jjw1bVe9dco71S4OyP36ADZusKQ+5belI9+Y2ot5FGHjQmbBR4EoYwi816JTO/XviQxMW
mtEHFMQdEtnRoj0L/AqRddr0z9SDSmC14eYwC+Hsm+UInyoLIsrY+OIN9QoUKwIPxZ+0mXwj/b+K
+tOdccZJSYFSswnzTNj09sHei7udUOsPFVjaulWbPpmA1+r+8ayYKOdAYLWDLEgK97AN9hIw0782
dA9duWZVm2nMHt/FSDXJeNiGW6CEuPNArz/KQo6oYNL1rKiOQCYSNNWKUjhMSLjUOVmqZOG4yB2w
1DdGvvvI0hKFYnOYsEiGM6YtEfIgelrHMURVOAAfSr743oxK0bloeSwjaYlnq2Mw1F3xVOGG40OS
uGImcfX+9hYS+zrerH8m+7gm7YkLK7eI3f2Uh2wFPc4EbBKdhUs3kMJRmMYh2+hFDs0GYWKIFHQo
87tEx7i+uo4mK+3orobqfxgQHr7SToczsV5V0uOwYZOvtGOEvZgLwE28UTwo8SO0C7LBwQ+2V+3a
z751Qojl/Lb7svH8X5sDgzWvMVM9c+sTiqX1zGyHUbFxABAoHr7u2+3qxK4iNDeudmrApt1UTqH6
cCjI/bAcaZ6Pr/FmYWoB4zDa5tSDC/Qhiw8MAFZYZPDxOcEtAxgd1YPstH3VdbQPHWdXESHtdm2l
w4oW2AOpI6xbGPjCKKG9FRczhIn1QzctpSJMQ7CPTVWVvnUz74ybsGq/WhTBWVNMSIlNet9sBLk4
rx7e528rG+wgWB/4S6lsdxt77TYGl1R62Fb5+9ECWFtmmUz3b7KFPFkHN6b2vSyOznDyvLNZCQYv
q4ix97KmotrxnWmyQRLujpl+592YZLI+ekT0WxIoreDQhibIfox9vWuAF1zoO5AVlWHNW/uZMFEM
c/mVnW+o/fW3Iv+GPZc3hk6aRNaNqxdYhOHl2kY0QRTmP6OuGB34iFrbKBKvWyOIztwqkiM/gW0j
5qBbXMteM1vlUte4E6FaN915FJt9MWHojNpAa1Vd0oZD9Ef47gtB/++UHIH4wGqVFUDznUuzuYjt
MHk8OTC/xBvxCSHdlYVp+GVG1TFqE1hTsZTwbnnt8TqInfZQFuIhfIbg0GfetiY/vQxq43H9yj5J
u5F0R0fbpyCq0U78XC5SX1T/KV2mh9P0BT1/4R2PsamGmt+qQd3k9c/2iESeq1oSaIusbPSYQuaT
dOLA88eJ5iRhsvfZbOwWjlcqkRfp+OQ0YWiR+yc+pB/DpC0+3/3tAPsMUSElqUVXu+9G1cCKZWhA
fIVn7CmU39fBlEtw3wHYuAfmQYqZ8cWfPkAhQakyPOGKl1n8Yb1lc9t/PdkyGN5XRnImRrxL9bz+
DnJXkHDTWNRqYkJmGxH9WM/NXSs/ICEG+3VNXxS01+9TxbZHVCP/5T4omldKfUOJeqklwRIgL7Vk
S+ursuffAaa+IwRG9yhS9hlyPZLUbIVmUH3r1MCLj2NqshinWjSsH1lgaApymGN7O3zwTwrLD/wh
zCW57URvjYeV70keOF4qmpB+CHOboh7MhLar387/fqA0cVk76heMpB6PBJNOihRdTtwtsLC5lWkI
utRUhz26wJrsPyrfmulh5fu7HVWLbbpnGSGbGIMO2svjd/PVNXFnVg2ZS1l9MHXnGoEasBrx5myh
VRY44md9EC3UEA1H6ar9ReviY56vA/f0hTZqXQ5B32xQtRA4ZkyUl3SLB7zZ6W93N5CIg4wgu5Bc
DhRZ/JbvMSFko4OfVW6LcfVoR542bL12tHph1kVuwMYac1SgCb0Bm63qUNcorTJk0f6oJsoioF5x
t/Ic5CHReEkyTyMH3iW3LCZdebmc+z+s9DddxCZeOJKPVaEKAMzyBUgPZ2y3szjdXVt5WkjOgae7
H8tuMaO7uGLfh2IZBh3wGBmDlNCQhQkePp55W6BtchxHGA68jnbjf/Qizg5vHl7qt4xwcoS/EChW
I+18O2mR7yqx7o6AhK6dQ+x8409QPmEwSz95HfKNDIpP5D5lR4db98+CwG3cBMf6bip4HV0lsn0w
/qHTQNbUh9POxVSMtYDWm9F7qJucfV7+vyaX/MNyHLDZpnPnfGNDGVl+0nb327+jkNyezqbEFhhv
97AoJtjmoGXlbAbpgmT+sHE7tWoKFwDS+OD1Tw4o6BK0FyJIDeegCGhv54N5QSDLR8H7ch20wNXh
KeM1BMHOv1xVRF54yxtHkUTaQaO8Gc9b9vF4aho0PV2TLRlCZqlKQ6pUaYXteF35qbX7eiSEv3Y6
qt/zlMCdzNTYoDxAidABJMilkweiHOes/dNx76XDblGlCMOb2T3z4fsITRazt/32PHTrnhcKo7Pd
DlYTjtiZ5IuRp6ipIl/TZdLy0MX4sFF7cS5Ye/sT3cZeJIgxEKB9ipOEFaID/t2lKgu6RdipbQMp
2k384jHWFsgZi8SzMBL38b7zk1+hO7QNExLG3+x9LK7OhIfrrDgx+fvdG2Ujrde/ZwjDYwh6i22B
MSVzdvc3t8bFjO+owgNdRkzIHugIiYBqJ4qOsa4QNGzwuaeWow5QXSmB+Y9YZ+ewDYjyFphKyLXd
D0p5Sy1YfB5OGQ1xjluthVaryz3Kjuhd1eici5nZPxsTS5820kPoI4ssq2KoBAia8xMoD4WSGNGs
GgzRzuDi6Xy6WICjRCcRFrVsjdccw6SnTOyYddIeE2dEw4LPSRAsAi2C9+gmWlchMzmIElBVLW8G
fP1nPpff4HfJYj1mOft2UI71BBH5n8GZA/c0/2n6GNzwcbYm8QFrjU8Wco8lbgkRO8NVvbp3aGqQ
7kRzQnCmRA+N0AS7vIrJJxgriuwiYGPRxhhVbLIT0VDIAjICgs2kTWlb7siITXt9XgGUN+si52NX
vIoTpj3P16LAUDIWHQF542iKMf98xci6/CRBGHHedU/leftoWx4UKP2DtcbQn4J/ajdsbVfKoeY2
evYuD+dwsWSygWQB/0Ld3h0iD9WLN7RzsGul7UgaOG10inSY7mIYf8VrHphNzy/zl982Q0upUuI+
TGnITMV61JhOdplhMqTKeMDk8Q0vRMzr86WjsgUyAeIBtHpsquztjyOAmZHaiPJN0mE9nNXVFJee
05AeMntPMyGTsfDgKXlmncHLzhtCjIGoHD4GAML0zQAhuarVLJdZDodtb7xwx+tK2Iyq0ZasYtZI
y4y6LnLKiIpoTva0MABKw9a369swsjeo72DMJAUqRgvigVb4Cn1Dgg1mD+BKneoE7LMcaF26Rc7U
4LjIYvoor90CAk8SXpFCSMU+t7xci7IuaVfurY6hYjPGRywPRVkx8lnFogukYgaciSMpKCa8HgJs
rXaLQnQbFtPwEcN9lsrYHp1NQLgfCe04kPyx1q/Otdh+K3QqOK59//o5qEwhPxUz4WDxjclHCEk1
/3rhBUrhF4o2GaqDJh7D+rhiztZNBPujjo8yeG7yLjelEEpmepV10UnYlhSozR1sLJOfUq04v5E2
gv3Ff42P7bu/x+MDxlof/ET/LLdPPZ2PvaF9xpd4DEpwbZUGj9kOf3uWtlql7iGk5nsVNWX3oQPU
AXdav70rBzPlMjkEpyvE3lJSfPwMWrhXI6wyAfUwA3pry4bEJtITTUhgvhnNLCa+ZobuPCIrw/6A
5rZec9Uxhq/flaMoMZa6Aha0A64u44PlunYRXL1N5RrIY8eIP9YjNloJ7/m6LsELlFA3Hu1FhwhW
NlaI5ggFvzDxMR7cY/AJGP70jU1dOmbJsVI58hj5Ced+QPTIRfSE++HmxDg1Vt08TaiTNI39LSAU
sxifOJ743vCtusbKECK+oEOF0lezbXB9Msto8ESSsQ3Iewa40b1kRIXSU6rzlhp08osswf5kG2RG
tyqBW89nG12IoC18s4skdvBg/3+QbtXDm6f2P78wMQR0sVSBy2kfXVTOOHsRcdm9rSMQ8o8fbqum
G3pXjMtKuN0p6DGGbCdzQ9GPAdehcGgFOScIQVufZJPa7tsJzLdDR3o8E2CZ4NLIQlWMlZSOONvU
ajcqMhuyAx3yT2fJwIa5y4EqR34+YeUJPay/Y+2DItaYWXORaeZh0y5pLXRbazR1nElvGCFxC7PA
uNAgE7aLu9Fq6kW4e++Az4XXc76DLZoRIDijg256EE3Y2hSjDnYErCpzKzeegzeU2AdG3J2OyU19
Vqnb6DZeWOlPhQPHTGXY6/9jmx55Nvvz4BATdnMe8W07PjUwx8Zf/dr5eNMJMPfoEXycMaKn/ELT
CnXAqKzDYotKWlYzw/QlgyLtuitbefESk568DYdkrS0dUp+rCLp+1nK/Tp9H3ozsFVUc+hpKKACV
9TFVZSlpYViynPc+2OdceO9jCDLUT/8p+6padPOOM8054pHdisJPAclj0PS9JbRpDMgPuh0M1h37
3nK/Yg+i5hLpxvLt6O7v2gNVMVmHZ/s+u/ivo2V88RhkvyoiWo7QCkHdN8OqL4M3DuyPXLIiIBK1
kaaIrXPjykSM7yRoTH8WHdDOOjmpTM4Hz7f7dAjGuX/iJ+sprR7PmtjUXX4Yt60JLWi+RhmQ4XLv
8GfPWHCcVHBgvwkoRQIFPDkOURy8KI5R11qRaH0X+UdSNldk3fs66X9EfTDD1IBK+PP4+Qvuhli1
B/28T6B60X6wONuhXtZAFbV97rvuwUmVyqcxgaIYaGxtIu+aF2WptcZcozuE8eMPEhHKUPrz7594
Sg6VXuUTMI5Hup2kL+PZi1ExBD/BX4gZnnYdTAcSxKq6gE9v9Fu4cluqJJlI4uqvPQVqIuXwEXm1
NmQ80J5awTKnTo1AcY9AJqSyAuecX2abCOoWAtZTVzjoE3/HtE3KUflP6a1ebuPKuLQI/WyTU7sI
9UkVcERcBt7lJm3BGVgK7Nz/4vC+tU+NkVIrEYiw2DgagazqHUB/d6W4g7TS5EGXN/5izHP4Wpqk
dcVXm7FvudjU7xFzA9cG7JGMKTTo8tKHjUZ5iRlxkr1xtyhK6NPZWTkT8PAtG41hdZMdYBman92C
h7IJvWm/qeckohypA8QEhZyAoH25mGdLXwgFP3XVhbeaX8XNwdbKIK0AUs+Xc7G3VJT9WVLLJX2C
6a5MMZG2ktOkTjrLsiFy9lTGuuBfL/nzLuqAe9peYYZs1jsmTWD2jb3gY4r/MDdOPo41FLP9IKk3
XBl7ySPQGZsPI539CqhP3Hq9/p3hJlAntZrgLrosZPpF0wHB3kUJ1ypywgxD721R9VAMLDm93TS8
g6wh3Q+I240uwZ9zL+fdUnSrszSI0o82lOnpPun9AbSKAykWurQ2RpI47DHKeQAozl70fBRxsIgo
QQ112ueHwFxST7fwY/ifJEoinZc3tXj/MWpVQtCty55dWm8S7PFmT9J4DyM17kI0ytSQmbCH3lMr
8w4ChOQmuAZPyb5SoPMKbKlc5nL+IaST/gDHlyWgKauP+4R83oPbJSpd7bdJ4qQ1D47mI9TIK+Cu
ld1nJ7Ci2nuFS5UNCa5TM1nWyzL5+j2XjpDT5+QMt7Ub2cpC25If5qLqYWGNerTg65ry3O+1wenw
fxFn+LejBdS9wCQCkbN7Mxgv6M/oki0im/ekO8yXiU/BRGJzg8xzOATIJcie3uwa6ekixljBHA8J
IILNUfpi1rqps1P+kTzzBwOlx5ZgfqZmPaMmgVszto1nQhwcmDza5bXi1zNYCgg4gL1aZLp0Xgcw
KIBs5wAMsQF3vD54Dl9LD9EWFK5uZUrRR9rZOvt5rSHwLSKfbPrA1+ix+wcCagQQJK0+RxOA9sET
otidrZNjwh8sqKOz+oVlIouQOKH/lWfnzyDmIkzrTi8NVQJrg078qjK140q+Ygo6yF8kGlp8Wb7P
FQISegtbyVfE3tY47y4tTKrbSqJH0e92Zzs6wxibDG16jw5sjdH+rJlD5CoNLtVDee/iOtJcrMBA
aClBl0B7QKkM+XSpiyVECVw6LYPs1n65kNsH0nr/BNP7E4xXYGwO4KeKD46QsTwma1PpY+OA/QDS
4lAhpVtFRafoXDwlboymTbX8Wp55QgTbXhIQdamIOUg925yYst03QX8aAcG3nThgq94IgnSGVvBn
xvlMNDy3MlUTx/SezBzrPxDURJrGjZwYV+OOG9W5yKR9W4yIRactA28W9zYMZQQC1Np6Y4z3d7kj
bXs43vx31bOylhB8kQ6iEs+nksk3h0ZLFHXkO0GWKb9iiU7QOsnqigtJVqUNd2knXTwgqYAb2WCY
dNhRzscTLSLpN4JlIwyBZ4v/AlrW1tn3Q1GnDst+PtrXnjLmV45eZ9kf/HYsVCNa0BmDf4LoY3OO
TSI+WjPHmZ5Kg9t8nKWnHUnUlUXPUv4ynhH2HVrZHwhIXVcXIamUO+zmkBIHW6jiuE/W1pkI3bUa
oAnBcHltwnkPBDQSVhJW/vPb/RidI9Etn61I9ChaxZmcIT7clOcEbxmvSokxiy7xkCK7hg+6Yv3K
/Qf5MIBL66jdBQZb4r6ZRAvCu1Mt6Sbk4GeLfNaNrNriGK2E8kkFBN9lZfJ/dHhPH4UNFuiRjFEK
qRB4x4rYoXPyCD+hlnmjcQOn6fopT+FoN4mbbaTUm6b5HEgRzgNYES1ZCHGBMXgDY5JUC765J79d
UQ1xdGR2kh8F1tg64yZ7iQoxy3qcsy3NKNB5yLue0isLXNzSRqCBiSFaoFDKZMiQaOk2lQ4i2G5w
iAsKDp5g7ivF5K2gpMrXpGaoNrNzwLLi9YPVv1U/hRAxw/JYBWrSF63RK1QTR9weErE14Tm63FHS
MB3WnfG5EWBNIMeaDllKU3E396/2VPL4Bax3oAwSYzB4F8kUL7mTQSab8cYaL1I4N3Mi2+Q1tlb3
Qj0H4ZDkoZaU4ith/sHB1Lv1NkhDp/rwIESFr76mLA3OgIXDJtlN95+ggGexDNVg4G4RAOMaHfXm
uuOjlJ5f9cV9i/06d3V3SlKIVgUW09r2ZWmERUqdGQU3SgU5aWf28QEHKtopJpYmNfR7/M2yKOV1
71cSqIHgnKAJX6oc0r2QdTvK9SPV+Xyyg4HUd1WLpGmQkYDpoQUaYAT+oNRaKC2f8Mp8R96a2Bpo
O9Qu4BQU94TfNwJG+41sFKJg+jshzLKFmun5T4OiLWzsW0dnWCYoeBUXzRpaiV6cHoGGTNnVlReN
Rg1e51Ds59m5WqdJCRkz0UXVtIAyI1Ddbx1cS2Os0lTYYlwsDm4xsqiOI3R0PvswIgcpsTCq69Ae
14AzJrlBeK1SPD2ma2xmdbi42M8D4zgnWnV0TImSghfqZpKaK7C9XWewgHGpuemLXdizkhYGEhca
jk5WuPJhZsRr5i/58JV5xcfBij5NWZw5NeAQAusZO3Lwx1bkF44FWktCR1l6+lIBHgp1lV4icigQ
Z5iPV6hi8h8b+B3ri5IqRoDgQgSg3OBkMD9J2/8ztCmzI50ho81Z25SkAeXtOK8ZyvmNqZ5moATm
1GzvtnDvpwj1QoF4Kgr7Rk628TlUIrBgTzVDOb6tOhPv7Hcoz3VU43tUgwaRI6shKRDxgQH+twYh
qYk2QA6b1880cwb10fssQyjKeDUTuPhFUcp4XCz30WRAhD5Astj8QKYMFM66s9s4v1Dv58x6i4OT
+PXnvPYrdm5buIDtkoCest3GeKTKjGAM0NzMAEZiIfyU1YQRZdcwcqm3tUm3WXDqJZ8kLctUlGC3
VU76n3q7njRJi0BsbrPC0cyRZV7zZeWIsX8AaE9usGP/xwUcV0gEUG5cKGEkUCOQKWq2byTj9ryg
EjeP1Zvk1bvPbUMaK++9G6bCyb/vONv69H1bZHDEfjO7E6GbQvv73F+C2BwcTb5l576/dAIRY4gE
eVwjf0PmQfpAvsntt27Ze2bY+v4L/mzDPvyyeaQTzGezyOJ2Ml25a5zLVmld2xTxw3JT+lkg76N1
flpyIX7gAB9J+/qcNbxheKNRmEzLHSS9udprJNaEMRD4d8bvVoIwSGeN+uIXlNR2zbxMCnlebJAn
fNvOWYbTIfXiW6RMwk3ystf+sIzkoQoTk+8Zkcj+nCMjEZRCa4o2wEs433xN2Kl34zTjZitp7cv8
AfPd0cuCi3r7SfioDm2C5go5ZIAgGejwKdrCbldXPqEhUO9wnTZWwxF2Uk9bWyP51GbyTUSCFSSO
GQzaWRr6kbHThcnY4TwkVOD1Bbwv/T6P2CsPYPC2GN3/vNZyVDny+s9gjbsEmOvSqNVrV/+FFQLf
oaVcn9CuNKbDaKb/MOmrYpHsx940B/JmU6Q/+dZ+VyWeb3XRHiYtpZ/QHWew7jRcYNd73qRlEqM9
UElha8ZS1egBgcWutcSfjbAwhUkx7aKpgj5LKWs/2LteENcnkkCR16toLRKGK3mxe7uBkleaNWNb
chxvlmXwJjDcz1aZr2+SDKOOUfCu1ZFGf3kyCcpGD7NBSR4mujlu7llbu256JNrx23HLvkAsz9WA
HDhgWUmigKVmx3XDZkaTMGXK4H97v8en1X+6lF3kMYVfBWgi0maa7ctdmPETdiwh6t7JlJE69gxB
3cjRUTrMB31HEKq/p9GT7dJ8OyW5tkJY6QiNvpxBnAQFo8RX/eiCe746YTrewy9wnhfZbTNG4JPZ
K8MraWf2ZA4+K9JdKSkcBMmJo2N0ACEoVH6dS994BCNtLlWdfOTNikLp5ME7NTXmvGkQcxiQQnyS
4taCTDggZpv3M8wMFNmFsHaNHaPpZB+E1yEI34k3lMWks+fTKmwBo58FBF4iCzBo3G8eNZq1gcaW
EOEuPEDkz6/qb+w6/FpT3HL7/RCl0V4aVGqPlNi4o0R333JtMqwNITU6Kmg57LqYMhNbkxl1+yEW
DjAOFrreZqiK8jhpS598im5MkyUwbX/gGP//QsVZtgBJpl7GT7QRseEZnEQyNZFBQzeExXYn9p26
AfblJS+nwyYsEiTbqeym+vNmRvBazEiieQTdsDUyzgCYwnu8Wr5KYGZZChmjqJbugugUuBD7dR6k
av0HFqDoAXaaGvm0wFdZMwPGiFH8/QBXmnYgAUY8sQRjgZIDdcaVhXcKQD+a8748RfLMpRcATX7D
c7wl3ZDwpyrjt8PG2L/LqL30wG1HVn5QZUf/uTQj3rF6YyCMkxR/3iALO5mmIN+QPsu2J/E9bGIj
rBVjjzoPJFBsXtpPYw7/0rK4stsKgW1wObjY4yj52OsNBKyEzrM732K7h2wd+VmwGH2eZfsgmolx
Wo3UqgJBDM33Jz1DRh+eY9OZbLL38qLJPd3jSSjwszjj/A9qqk8uMXRJnochkjjAG2+D/VsqROVW
FJ90egPLk2Ruh5U18S64NpdGA50J3YyziCCO4uCl9UiLM8f9q47Znj3nDlFjXDDGNj336safWWbB
AWO5zgKKQY94ygm0nVjs+Fahs/Xp7z3guTrmBUFvy2VWzPHkOZVth2J2tzSnfCZM2ydTSVY9ZH59
tgn9oAMMILAgEatQjPIqbS5qU8aBkfw6/uP/+RJFfcZIdM2bElkRUHw3yBYMa+UPLpTckEuvBCkd
ojU4wPt4x8A7FoC1mSxOnW+lc9Zbb5HLS3ztwmEFTeYrZYIvRc7FT4w9u9TlT7L56plC3kM3yY4o
X4eAkld7auetYAgEdnnHnkEISHzSCRBXWGqR5bC/4rKaI0Y+unXJtTnkr54hz65G/2pm74fJNK+Y
Nv9im9QLnVrI3MNBWw2XGS/dcrP+GYqFlX/RhYrOtbsFZAbgArocyQ4DVrgbCP4BiGKonb6XdsQ2
S286j13sEVsz33AnQOkH/I816736vtvelorbmcC7A7l1uFJOdkYC0ONyAvIt6VFpYnKfk7Yan6k4
Z28lrlU+tj8FpwundatCJjB9GHgS3/em3be8FMAcCXewQHbsP1N6KEe4QZdTH+tj2ublB5qy/YDc
xNmBtHBIZLd5MytFOgJ/sG5MJlm0J0/cqzKB3rAfcIZhAKAwawFDvoAZsgdFOVtq80b+eXDfbvc2
fM0ZCnA7ZyNUtuTQKoegk+eFuidUm4EZ6ro5AEYcogo5h9k2XyIOX37bSVmzUYcHRbK06N7XXC00
iorYBPZfoOs8DlAjTOjaoXpm0ztkZEeEVR9SsTaoOBIQbvXvs/I4+wPN/jADiI2fcwqqsDlgyd1h
ltyD5SW/TG1g+I52HsaixoKRCab37rNCC42f6OXrH/erQLOoDkLdmi+8bDBUqhjuTFjsfjGiKFLI
U76SUAvCdBssoWq4zQGNX9WKmpMndnJOEUcG4pPRGJofaeo+PZjUoIg2vPz1KZXNZ3mjAnKCGMjV
W3otSLk3grxPrvnOpq/4Dv7u5jI2HIgu0E1XReil+GyLqGKxmDSBhwDcsAbPSGa5a+npclJWmdjI
1pT9KrDixkJP4o2H+dMy8Q/0Muy7eFUKFPv6nFvjvtMhUIZpxReTeXARP38p/hhtjfeqd8hWUozr
jl6Rnxg0AeCC8R7fROndq30cKmcas7DnGUflZ6r6E+crILzPtE2pvmc4N35ctUM/tuCPuKbjUN83
hV64MmQ+rIcjzjat8GuHfVMwDoZfnlkhpwUUaSipu89MjnmmvaJhh5g4Chy+ROK1SbZSjIcBVD1x
ivLSviIm6af2ZJqfZteDqdD3WPd5DMdwUPo4iYoZZ8vpwF91XsAyxn+yUv+QKnSW/RY+bfD/bdo0
8e9uNbINqDR4Df917hF3WJRNP6du3Qbp2rVnuqeTlFaXHGtIP4pZHYPIkox1LSdUsxzHHGp3J2nD
1JOkmsuPawX5QYIEhDLJ2YcOSbxdV6BApaNN2eBGr4sazm/nnn7lj6H+nfHoZUq+5Ups2MLELJmG
YyhQMcVpJPUAqU34FVI6wk9Fh3M0Bl1hTm3/5bX6d1c4NCdc580APqEHQOcqin1eTsYOoejSbKHQ
VX7W+rp0Yz7jWBejq9xMRuHWgFfTrbrCFF/3XNuwTJfcrM/2ErOJaiuT0zaB4N4Su30yEUbP+he/
mkHQs3N94r27yYM0X2vLDHlVzYy+ND8ro5WFHAtOiJ+Nbn1TmMx8ClWTKyaF6e2xK4k9ajcE9UuZ
ti4F3z06/6a6TXGM320ygnH8dczqn8mchvGYvejcf8Goa8T34ABiNegqrmyX1LNEVQ55lTXliuQd
aDd+VDBqSLpt10iEV55Ar8U+EvfZAgc4voYt0CndWtjxOs+JEMYI7Visyw9biawtKEVHppwgx2H0
cHQuQhhqdAASVRUGwOnyjvaRDnPVH2tT26WY5g0+ecxnp6ZVDbSheTCMl3NwY8cuHl4iqvBDnaW5
IK7FGY5Hn19eiAOlGWgegsAlFLH7QqMvReSCWWMHRD44KgH6DYs7P14etuH0TkPB9534XOPp/cpA
RCEw/lDQVRVB8/RpQrVCrq2yOZ5/nvbrb+m2BUTkcvMiEgoyrpvliaI/5u3HrgCFFcS97jt0DMHj
gW431zTyTj/m/WrhDGpRixRP6Wu95d5SRkwDfnbGTTG+PIao7yd7SBHV9GCE7yQd1W1EMr2ZFGG2
DfrcJFJ1I5QQrTVTXf/0m4s4gV1Hgfngo22Q1DTHdATrqH9PXyCM6LKK9Zby7HFpwcOfgwh1SWf+
yWdUDiLzS/K9Bs+CMCv6WWTMGzwsrk0ZjI/Ycurq0t9n9bpPS1mtqCE4Zf1khXlbjnvhasS9wqOl
IZo/eLV0mfritH2NBymFwTDbOQMzYMyRYt/xvAWP/ElgVHUjhAyCeywcXKV1BfV2anpiHYyrJu5G
NesX4Os4FJ/ZFX9NQXXJZRpihAFOUJuDDFB/GPG7WXO7yk4o4UFKSC3QsAw3YSXpTvUoqIEGMfEv
7t1fC0Lj49L1L8C/rcfbGez0SxHlufctJFzN3g/Fw9ZCmzV43xLhNXpBaLPVcbXIPTeDQdRH0Zde
bXAmIF1TEFlFOq7bkPS3UHntHpo2cUY2RBb4/trDR2Ja56x0Wl8hEE8V5JXzMtWG58VIH2MIipc6
Exh5+MMeyl07CyAEmak5i8/py+ippFraKFUD1ncEiPkRTG33PWf48hX9f2Frha1RssqKRvAHpDJI
6YjIxLdeNnO1RGlsIm+yTFfhhKxCKTUDC2CdzsYlZHl8OetpSHrn2kMimd96YbeaPN/nFLXTMMIx
cry6ljrMxuz+x+ieGNDWvNBsNxUS1QculY4VMvtMLbZuSG2rT9A2xbOA4sLOIev+0UaoZetmo3dW
tX4wKvCibVrORxJ2DN+2ItzYikvAMfQbLVrLBPYveAmBV2/jkYbSnkMiFw+2u1GbThdcmUgg+jJm
RQuQm0PEkSS66u9rkSFMOu+eH2TynT7zjtddhsxSXZCRf8Oqj99Slzdekc6SHiJciKu7p4Sdc33c
V8atagRQxSvTNRV6ypd7Pz5WE8h99pT1LyErnMLM1cc1iBJMWJl3OylL7nbO/RUVPpbUlfSQALrk
mcBn1qjle73MuS+eFniw3dYgNuM0gL5g1fv8ZXwUKFwJOz4FRlvqZ6GKQnosaMQrxu5Lm6Vnenew
biu/nx0/MRHYbgzJodt+EFJmGsESvFh3cNNzO/XoSqXwisKaJg3waT+pRVZHc4ip8VFe0lOm6D84
Fi+g2boMP0vciLkk1J8XdfI1+zQqUZHYgd+kBQ4YEa/SwzKFN75wRo8sO2YiZqI3BPOwZ3Cjwj6K
TVwJQd6oAHTG+zQdP5cxzYNbQgnKdKhyJRacphm9PMm+AWnp6+mriXhotCwX0pGfDfVaRItkmprZ
NKrunWyco8xCXkVhryZdCYKEVLZoW6Gn
`protect end_protected

