

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
cQDd3XIPPlgRDhqULvYHvwCty2ZrVwzfefmANvx1dZIylIMC/SlAcj88wfYJOEUSOPC1U3p3rRJH
cF/G+RPdfg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
hcwXqOGXIKp1yMXglvtwKNDD2csTguI/218BbAfP1Qe5YaY7t7J14bh3PN4/sY8v5SUfs5PPhYYF
AVoQ7+Y8KyIAkFOjVjl8Q3cizlaMAyaX6UCc4wmflvCCOjy7mkT0VJKPELyiFH5OE1gTiKu4NfqY
cLpas2QiSAVn/xZw83g=


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JJiSVarYWytdLFzHp3wkrD5+jxEb6zxCxwIxMuHES7X4vO/81ppoMZmSB67P59pBX5Chyu0EswKT
bCRha6XDZljqkcBWrrqj3cLRE57UCaEr1RVpDNBMw7hjNrwCb9eTELEwb3X0mZPKBqVrRNroBMN5
Mb9o7SPJ2GKhIDEDF5Q=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
x9rjekK3vn0E248BFQkRU8rm2REs1XV6NiMfscimCVnt3moe1QOgVJzTLPCcPYvThLcZJXwVyFUX
J1k2lVxuHKaC3FNNToKLX7girUcVANbS6jS2AjaAfdpYmQXF6epSjXy+KOWM7AfrGv2r7XNIcV6T
P4He3ZDDIABlWanBaDiVD6NYtB9SspFXaifjJ2faT9Et8gWmYJogYQ4BjXl960BUcxWS5faBudWm
MidcfsfVFpzH5bJ9L+thBkdIh/P3Rjr9ssCSzEagp+1l0DsZGX583KqMaKiaZiIsR+KyQ8Hrld0H
vh5k+kh3k9z7ewkJNwM0LCpa2Y0qGSJOxIauzg==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bMGW+/GNxe7XIGxZQsPwYg9NhBUySelE4d3DawPwcsMkcAefxMJ1JdlslSvSp+VjxIobQhkauqfs
plGQEEjRkhr+3m8iz7uiwT6s+TtBZQ509t+m12KAHsziCshi0m7JEPgqnpkYUxS5ZbKQCRgudms0
J1TIIpIIdBJiHjiJWPFKhl2FSk46olekE0MQ/LvS36IE6UC8sP+H2MLZpAxpzqHuZ9TNFvVcyr9C
pc7viw1i7pElJF0USsLWRjDFrkLdXdznJwKPhjmDvq2WWhH0UZss4B7FZEDrUrjB/HO8EjVy2Hj1
fpw3eQ84VC/StEBHWhh2/ovbE1xsoAsXeBE8Tw==


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pp8HZNaXt/evJqKzoiOa8A1cmkUh/1mQf/2Vkpam3N+hCoX7wAAqGU/zZVMPYP16RpMjeC5zeSin
YvUeVcdgv5x+e+joKUcjexTi2LwQorDqPIl0bCwYx4LccUexnWG6I9/pSM85Q6QNP03F3dTfZ+nY
q8I48HLVTNxhG5xD9+JTBp8D7rjXe9TJGi+hVikOsYhuY2PrwtvuAWhuicAfJnsIE23LJrp0i1cL
6oyVsfKsx+68L6qOWniySUGZ5yDe5zDF3WoQ1oHIZl8/tfnTJcGPsIRyeo3fpk/6/w5zWnz1pHuZ
HvGPaU9zIF3KNoE/3qKTDNhAcVbvP4+ohJfKxw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4784)
`protect data_block
ufGjJ2eQAYu3yVAh9icN1gNsLxeVXpp9NuTk/xseCFQC+8+W0u7tp0cOE36mFJSDltF16UJjzO4n
FtQAy6aGGGhVcP8UzGJcieqSw6gXcxSbhHYNeYWE/TWfYMGyop7nrIKsTiBSkqzfwq4qBMBEdgLo
y7wPvobpdNdWWN5xAz9qFjr6UUWUDoGKdHf30X3SRJyT9E0hKle99/b09DVzXVfTJdb2htgxr4e1
/3RPHot9GUu+W9SRzZMIiFkCW2zAe94NLUm35cVXuZvzbwA7myvNcnBO6FLqK6jSEGtdYXIRuvyR
/pO9WtQUtTb91HYk37BdbkysOaDBErGll6jPGZG65bcONSGeYKEVovK0mQ6V0SpJ5IvdPNsZl26L
ddEzgUqa96EFSkh/x+JUY9UK/Oif2HejUOPR1AIueo9a6AnhyiU4sTXH5eHDBjbgBOKaAnfUmrdf
ZMNaPIIvyErz/EGyZtdAJfb/y52LejtSmZl2pBq2NM5Jw1lHHHxHwSAhBSx7f0ws76dV6xkcQUPJ
ECIhukvIlEKtUo4x2lSwisIufmDAF6d/8IN0G+sCKbNHpWb6XirkScA2A1hoHCIBCQoAQhpXyUdy
hHwxDb2l88pWeI+S9g5ZcvhduqPn3Md0RcYXeTlOEXhYwGU9jP2XwAHc5I6V37YvmM1T/SJwVh1M
YG/HImfMjn2vtq9FRJ2M0he2aNkxT74C3Iw7gk34iFjAeH9ty7wTJdSzcjxPPJp/BgoTps18VL4x
1SZ5f+nfDV/fEplypWJ475SNyrpAuA1EpCy2iJ2azm0Zy2Rc7LzTsw4Qg8HulvhljTe/U6HBm0H1
N4c5XRKn17juHtofyUgMhC4KAZBCODkrRoB4+IaBerwaz5UjkgUxd7/qTROZWFYPQMnnPJx6yPcv
2I4eG0AlLtfiksaFJneKp1QntP5RIa/E7c9nz4BRww8HFpLTtLLaNjr3YhRY/LkaXJwlS2bT6xPE
bWAIY8zJ+27G8DSk8PRL9tFQ7cx6ali5I3gEvq9Bw5wK9Kl1M2/yWCat+BhN/0GMDHLfB5B8bcYC
H8RLjZsdmyXybsUtX1aqtBObT68Wi2q3HkbdEXQ/jmibYl7mn9S4s6o/im2Cm1hmBX+sGZsHEHgk
bid2p9fcw/DbI33j4DOEOV4KIIwPFwj0nqJ4tuhICaoiNKqkRP/VjYhFrbIWTqjAijO36aCYmzcV
N3M9pqWSDx6EHEmrE/KZvSgr2x0vEIKl7ENL4arV97WwdWfy+qfjWhpoXvtsMB4aG2GBE66p4GEX
7ecXcaTnzhkish2kwCnJYkvP61+LmSI9jVpNo7RXc+IZi0MR2+cCDGwQmBRwRNkbdL6PkUFKr9vC
R/Uzx/MI0f1iTng0UuP50ngxtz+wz3GsNJkNNvIrculWqoqKqWJL36z3kddKOTWrJpkVYrT4lLGT
1arUvhFz6zS+PdSPq0qlW6+zT/QZLnfoOE3na+R5VcAtTgaWkX/BjRLdF9oud2MKYShPStHA228L
qjvtqZmRZoJVTM6psO+YuTyKzDvedIORtmOoL6Kx20ugEPcsqA+LGmeCuSVb5ugFz86cE/kCjXc7
o77krm2HVlB3TDKOsj+v7BsSG+K+EFL64p2p8m6eP5uDEV5bwmS0yGgcS6QbWHMocfJrBRXtId+R
P7NhJx1PG0XuamNALfs561jk2vguBvupNO9g0WMb0QZGZ8XxiGwcR+68ihmEpAdu02QVmyF8MUTM
U/2CkuHwerwDDnf3t0XB40VpKFK5KQiXGFK1TSGKWn2RU1sEbkPzQpu3haeSJ1yjOCFLYMvbFA8U
rV/BGfsnI+g9bYlQoQsB2vXTjg80036GMpVlKROHvsgTFMeqVs1sEm1kKx1p5tdNGbwarImmMk4a
/O3eGQ+i80RsBnKMyjGkMmnawiGi0QvEZF9aQX52iaZwrFvweJy3Z4zmnfXkBr191/f+fNmP9hy3
ZxwvJp54dU6GMljYY1xvlGQ1VmdOusnDHR2TrQND9dnrzDzmhPvid6RD2pTQmFj9yKB92rWEgVMF
V63Xb3nPPY7DUh2gFw+QbUoGy0SuR6njLh2vVSBosKADBIi82oGDRkY6SR/gx/U96ShoVxsXT6MS
ZkVae+l2IVzEO6rLZmLsj0fglvjnesPldB04ADDh21DVFoTk9+5q3sziEqPC4I6/zxT3Gvib1HGR
RJ5nKvgiq/foBsnDB6SN54sVySKb8UUPwryMGKFEpPZ5zEI8IFVHFDoipcgbXp9A6Epvyp27B915
yfnwyzrjfQen+NJuIyPXoubVqgadMoEBFcsfc868USX39eCUoLI17ZeIXmPq2AKeb9sBGdW3EDaF
VAdNNC2h+TlHTzw2uIrjDW5B1kaAjqyjbuNr/KBhAr5gVMpsd+ZjFN4cbFaSUkhNLuKBs42ZyAWb
AJ/v66Sz9Qi1rZI4QBNwjQqgMEcx+KVnKYChalrSeVxqP2JNLjwmIT3T7hWftARlgjAfwVPAnNNW
0A06HXNSW1GtFLYg/cuccuot6vJl4gZMwTawGnx5ZNsPSaxvM++dOles4+2khT2GHFZIV7vr6ZJU
2BwpvvSM3aOBZpc8J3jA4+I3VoEJCAolSa2WBbuvHNX+hzMmHPjJag8ZDoSLKyDM72v29lxK8S+6
YIvEF3O+XJz6pXwmFr+NgInT4O0bBNkO8BZaQqzcElwbz8BKhwm8WYUilHR22W5ebZPiUMmPbsZc
KFG/0zYk+hir6A6L7yEzhkhj8wv2t2Ha0iWS1fowMBjTSi7pTfLfb+vBgFGR2mqDb8sYM/0avI7B
f3U9FHrR74DkYD2W+jq0AvKBFqN3POx4KI569C3SeDXxQx379wVEFDePVxITQbIKe7YFz6+QMU+z
Qt0q2yyaUbgxGQ9UGK09sYybaXtiPIdc7FfQWmvT4ALn71GpFBD75W5ubdD3P5gRRWbrcG3ht+pg
G6+LEAr10h5L9HaKNNtdBU8IhvP6HNfQle29gtEPyIdyCsywEVpZt7RGhqxMUXh+EKl1eOT9X8Nn
qCVtSOMaOLJowzHFxOfIr3+84ag//kSonZX1HxcB11rwJ05bl/YaxanZx9nE2HYkRuMIRZAhrlnn
lOcxLebSEw2O877bVl1Mn6Ut899dDjeUYfOpj6swDVC5NHrCfHfuY29STp3Pr8zVp4/lo+2WbC6A
5SfYUb9Fnj69rIaBTqZVLjlAmXOUQYgzdaRsA8+joUzUTwHbi0gjv12h/jb/RhfAUCSv/gs7MXIJ
TQOkq9jsEySF2jYAIYn8tvcCI2Wvwi7VLpxNuOUZjsZ0Ow3qOUJVn6XVpAPy+HxeH9Oiq14UTzaD
Oj4HQkIb3V1HP/2FY2KiE4PREjqD30CLhLk+B51h25h++PIFwUDdya5V+/DO3p6qH6kWjL/5sVyZ
QDkw/M0jfbDL/BiKULpL6dIxSb/377vJyyXq+8S+AnnfQZflS8352S152uaAs7EQhZBFgrXmIwxg
2Xn8nWTR3rqThBQvUUyDyCGKv0vxrtc5/uGKs1cteh+w4ZKQB/hI+CxjMV2vqb0oA0CIZbo69eaY
oRSOFhFaqY1kcQKb6zMKR3f/JA0EYLnsVSnv9BjN8YyGqP75YGdoZCMtTJdLdHVBd3ujqGC2yJjl
ewBwFjHL0m0nje4BX/rSPNS01Jsxkb2tWOyBVEK565mxQibCUaeQnFV9tt5kz8T4MBRgnyGPBKhB
bN2nHC4P8xK1iuZ5swyLaqmeHfLU2pGItkYBNm7vZLROZN6ykFAZKt4EUQ2e7ZGE8Ae+LcazRjgE
0NGlkZS+OBHzyTjSB7zilMW9A9xd8dlknqadnNqbPdOSTqY5n2XS15YT60fzHFE6Gt3EUHo/FKKf
42csX1fWpeu+DB+JhLlmDIeSKDiDi7KURnQEdxeRlfsY06ucuHickXKdaCB8vW4M2f6uTuZyVneG
2x4EJsWZ5oG1vuq4Lp16fDlcqvIRdIx3XwesO7nTlMpKq9P+POBolZlUDbkoNm55k18PDbXcJ3bC
A9pe3quk4lqjMadqqx/bbEGAL5pcgMlZ2iifU125a04Zyoq9zHjS4Dx6e7UY0LMFdDqkkMlvNIJT
HriR51Afo3ENLESE5FYbaIU5B6D07dckKIN+oLyw9CW+PXDe/v75/Fy84RSgLgmuYM2aXfMyJthr
Lbt2zIWIKCvfDU5LWFVDeQZ/6F3nnaxpdmY49Q+OSj1HwRKITHX9yHnRH4n5KEA6rc2PeqQA2muY
CGnAH1AD4rvYoMP5GtlAF3yJFJGAQ2HXJZB6TChBpqucCUXvu7nWHjzaOBqAP2CYAybHqtz2Fjpw
Pyp2aNXle7yIzQL/DTWm7TCOlXQFpmW9OB+/Np99LIL+GAPRmxsTQlPqz5YycfXlThIy5r/nrhmX
Sm7CdYUjfsGu6UjbYZqKPjsdHBP/RIXRU0hPCS3pXqiUnNcSPWCYW7C/Ju+AKvBombZs9y65JEj8
1tq97OFvOKZ8K/CO6hKb+e+6gdLpIjuRtLbTqZ1HEd22Hn1Kp/M8Z20+oLbi0g8pAO1RM84dBLv3
N27/q7DRBFlt9rCkZg3KDf3FVqFULsc29lWSlknbcgPQsqLllae5CUDGGKErZlizCWQdwTZE5xun
S4RjQEnuZpZl2T9SR+e1PnSbDvjZpMCeLgTCo4YK7i3XetY5LNIVqnTiznwSKTb3qZFTzbjorp8Y
vznarFF2FO2k05qkNQbopz1M72C13EX/wtLPTQH0jYhx8I/vTad4k7TJsiHe6q4+K+VB8T1PM5+X
suWTBSebZcwXblcuFWcmVdp0PaGhyHJWFysEBL9E9O2E+teqLoBdoaGuhGe0bW1qOlyagMedn8I9
usedHqWm8RWYsmfCL3gRr60NfmyFsrsaWrZrgopSgbLHDtks+BS/nwIMrKZJCUN1XZs8vA510DUq
bNaE/i05FTF7dBYSg5dVSVgQwt5NHIhMG3QhspDItm3mDa8ofk/jarlalAXcAWXEacXqG+L62Jp6
TpU7jtb+giDzTdSOcn7q1m4+kx/o7OF8nHDIkEhIXLhW9v9u0stZfAxaVYmfTYHteR0AJy08gYCm
VPQ2fvnTSm/PK8BuaYLZEaBgBHyUe7IFoDG6OCXsDLBK2uh3PK5w8Vdaph32wWfPmAJtugahRca4
ga+UAsiUfgatzXESO3ml42UokhshkVsnhsH7MjoVf/prMDWdKkW+SACPU8HoudOFMVXiNuDKqRXz
EdfumXBieNXz6TPYRcOHJwGYpnY5BLIu8cwy0V58AHSrF0t0XiPmgvwDefUk+86u8GoMVbiqoRj5
s4lyXWGE+sljW6tTMUHzHGrtmGyNNi1YEhTho9N7dSQ91R3bcvWa+BAONUyXUEFX7o08DEfWYlgx
B4WP+Tvzq4S4rLVaKMj0pNo3Vxkx5B04AEiumQkipXbNoIbNzfrs8mEOjad6yImAkpg2DFUOT/hh
xLr7+CZ1VGVZK97p8TfrZgkCkk2cYfB7JcHH65Sw6vKSsGve4wDDHbN3cK/UCVSxIiyKcXCSrVFU
7cNEqT4B2CfFmE9dFQkB9gOrxhHUAbNRiYrO1DewIC61g6QyjOVPM/obzBw/aonmNla2wQ7pduC5
wOlqmiuDtoLi+i2JAcFR7tGcNLALwdNzSMbZHSLnJhsvKlu3wcZD76vOYDnzjxeVmFedtfPKDPK8
OFltPUCt7HEPcsBaJv15SLXyCSx71rnQ1/njyxPC0JYwX22rO3LHwpJ7hUDk2zssY6adLMUNb5oH
OoyeuseqvrmMjnu8BrkSqIgT+KagLIZeOnwxvb5BzofDGdJ8Fd/fQD7AgvQLOI6req9gIpVqAsK8
X8Gndni+A5E6SQOTaG1V5tI4RFXb/9vGobARD5IDcmbFQp/iqw5kdXekdyvfbRUhfPVCbUlUB3Lf
pwB5EYdd9KAIoHKRyu8aSQPw386kBZOsSaajPbQ8stVAWYuUl2B8WWDACr/6EFZ7w84ZtB/06ML9
zyc7iHA1nMMwDGcF22XRBq/S6bb7m3RRv1VbrgPjHJ3/dPGBRsv2QjCA+Ctsd2QKGYExZoZ2FSYZ
7855YiIZrCksS6hxVBVPSK+VyR21ZKdz2QOUxby96MIUhNy46yZ+gcidlQrXxvidEFr2n6Jh2pQP
84r7Dbj9IB7tJXudeUgr7jjTpt9n+Xlw3Cf5vQwImkX9zhLZ9/2vE9bVFB2dc/mgMYi3knDgfLLG
ilalWn3mHYApHVRjSVjPKPqxvXsJasIJtOfotqMg8xkKODrgxzTi1V0ylqcV6pEixD7pHp6Bnhys
U3dCVFHnlL2odtbUQAVhwjtjI+SZdUMQeMYgpTpGMvg4MndHzqToggaFjSO30ZCOYA31BCo=
`protect end_protected

