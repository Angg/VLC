

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
gD7l84kB+WAh1ATog3H36h0/cMgn9QL5jGe9p9PjvP7N+FJAVvGVlrxcgBw6dZaWDNZqNANQuRFv
ZSE8fsSCFg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
YQUcxim/tlzHeVlJ7otHN7u41KO3Yg5DFb1yF4GCsbXGLtUvWNlkFjY+UPIlgYImR4Zo4dTHJQ+j
3BaUNSUOqAVzT9CfyUelv2YD2ZTfAtzIe1Mboyb3+StKnuzxnZmIhVPiZlowdW5lQ1r7BjDPOsge
ztxOfUTbvYcTUE1ABIE=


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
eu4MFD/NMz3pssr62VCh1XDd9mthYydX9VaOq3lWUwHi5/7e5dl2SAWHtYwTnBgGPY+jCcMycJhy
WSlkhQxVj5BsMm2aAItwXFvH2mSbjlPggtI0/+DNGQ4x8LQSFLTDYnnQbBrHlJymsS+/asMkXACD
SJ2tF8LF5tMhAlMPZZ0=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rNAzbNlIFUMjdhvgzZ2FokzvR4AuFtV+1AHGDKa9QgeBsZ1e0Fom48uKbJ9iakvqUoUcKKAvRzeY
OBkbx9P7Imx0gvIgzFsgiVw23cBYWOhbhSqVb7mef9aKx8yeF8T48n7gKldUkwBHIPeqaayRI9/Q
HCZO+k2+HCjRZE6L/Gzd+IOdEVUFOg3NtWFPk2JFkfZkxs8X7Vg/xxtvH7uvp+/EbVyiMbnwDT/p
NSqOyA+rJwBJYD3xRIPTFDI83XJLCF+1i4E8hyu7Y0F9MtjKugqEHwAG+JK3jde00nzNNaeLVUQ1
OfFMZJpkk0Cg66d2cvJY/G11oPkmvTq/JZ4+5g==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
apuTRT8aJu0TR7Ciy6ONiGK4AT7TUEiokS4gFf1g+kDg6PdKk9VRun4HKszIadRtahjPQo0of9uS
yvu3GS4EQo+Y+T116wnAIXnZSa8EQaEsDkziOI+rCvXv8IgaPYN8Cq0aRlASFL7IHOWNI49V0c0A
FIG/+5U7ZyNQFCVwuE4gCgK/pA6apm5kY4FGJft/EdZ5YAbR/nCTzK4P53+XsKHrtGfw+/MthFWz
tI0OtloKqc7laKZWKOVFqWq8Qmq7UL6utFODtxEQqzczH+q+Gw4rkUyOosIY+cbB67hX+GlmXXEF
jMwvUcen9t6c+wiH6rmBDcUIiuUHHz6q+jCwJQ==


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dfDj35aI8y6zqcW/IHFxmCDw2mpyex25qQAUnsL+tIRxivv/85PqpCOrf3b7NWnwUKMrsxtw+JBY
mtlPsVxQKR1gn6VkaHwbEgwxXXxFe71Z+1nWQhfF8Nt55jGvq1joWKMrurSV7Mo+HkvHMSszXj3v
8ElD0S6sN91oml0nObejOhxzHf0ybK+sGag+CFA7aBr4k4rYglf7AzOYrPl3nNoCkyrFDQFa46/w
SXJm/os7zUHbsDI5GGUH3BU+NktHZV6GK3iyhtHTwrMgDtpGk6vKHMKULM1Gjv9g1/jp9Ao4cUhr
bCVOXM1v2e8A3564rmh3if78zTzCKamPRAB5Ig==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5312)
`protect data_block
716GM0+0QFfhRz763sNyjVc9nfHih2iRatrw5kV06KAY9a+CaZG0mGeL4qpiIemzx6CxT9iy46rc
P2StC343+Z8czkhq/DZxPbx+EiDoRXY4imhawVw9LfyhTsrRZjPMLAu1lsDkRumR/JT6TDSdXKbP
5VqLCfUNT8m0E8NhoWCamQRCr/nczbVDuJfedUxBqNYzB7BSrWJnvkkDTT4fhODNGWg6L2Q5681I
Jk3yGtDBNcbDkkXO/Utd048SDfVGCy1jGcxdMZCIN9enG56vUjIC7tetNg+Mklc2FFhIyRWSfceJ
fbFCLfn+czWVekhiWnKQvmZN5Syp9FkrzTfOoC0jxKvdmjxXK+fin7mXPOaki9Hs6jJwP9TKDkB9
cIED+7uuLAOh/2nPn+NyHOe9O8/GYp1UW3Sl1WEVJ7/2Zci0cG3ybiRaq4lYzi4h2c9ehzAMfmqz
xWCjlHILYAGGvhhlfO1O7bI2IvIn+JvPxbb8RcRlteCBIC4QsJQ0CwwjqZX6OOz4ivmCyJFGaALM
6ZmmnpDsEWwQedt+hut4k4gjoPceTVk1hyT4iA3QX+W5rDpXETq+jpwfzUwA1Y7JQi4w8W1d9+kH
MAQNJQIwawdrRt3W5CsJxA4iTfcEMBatcO643KdBV66rIJdk0JmIMBgXnzzWcS5Sy/e7tVXZBBJW
oWeN8QskRt7qSM25DFdMNwPeqJm9QxugSUG/TnTyGogQdDj6A7xfH9DnlP38uDoDgk9tEX4X5mf2
zdFfot5/xLfJLfYKdC8s7ytbjpi3usaiDEEk9dAnwb/vhuk81RIp9E5qlGQNNSlxSe80iGDx37Ys
57p9LW6Csq7GDT4ZxMk67bWIsxYmAIUEykl8d27UdKwAA8L7rNSZStI2vHZp3aEP5tL/BEwpMfVK
OzGlNLj9cC8PnAU8YrO8jDe7CJMX6h7Kq8x3UMyZ05PYOXM0KjYzF384/+tVb56pijIWxJckj33a
yqR1e0ecq8ayNci4HRUhazDJ2yARcU8y8JRhtBeyHpCx6SyNnSdqdDskmZ1jn2nTCy6DmVIgOv8k
GuyWnCCTYM6oiMS8lYd4C7p44/NQ4MiHdl3WSvKeKWycRWy9ent/7NFK55YMe4lwMpLs6K7CFgrZ
ZZeSPrrsQpVKjQaX5hqhF/9tQz2XavAIU6A/8R9sndmp6DTviEyf0Mt2ubKAK0B1o1Z43P2+sECp
1GVpMFIhng6pLrM5Q1XVaPoTiwwOC8HE1Ut7IM8uY/5w6JsraBTIWvOsWlM3WizUVnyliCR+tU5D
PuQOG4XvWP39k2firr6ZBFtfZxVGboUb6UgK5L73S8DuIRHo1TojUYKs/aPc+lt2IHsJx0AhlHeF
xAQ3C44OuExejkMgk1qtMPA7PZiR6tllsnyawW0iXie8RqsCfHVVOyY39W0kG030BsJk1jT+wcBc
mQNeG0X0BumThjciDOgw7HkDdMuOb2M9T+7GSKX7pocIH1d6wlZg3FxGHGIVP+iv9dZZAxH2rtHX
W+HInvuv0TI5Ef9sW2jzEbhqoujqRGohTUIowB+Vo3ueTX8eYLvtHqaZEFViPDf0MhLrMHYhk1kA
2jaf908Ps7af0DlrE56ruW/GGXn0Oijh817IM3nZ6397MdoNctskHdodDC0xAjtzmBT1HivJ+vu/
vEJn62Dz9nNMsrV4HZ5AQa43XUkqIC5PRG76baCFWasNVos+Foc00UGqJqrTZJCAhG0KPPy/cHhN
IRMov7/ZyFwTMZqPoY64RPzQ8zW1LxJ5alAN6ZaZYObUzS9lxMdCxTHQySNPPL6G2YsbKQNwAv96
JtqRMae/06f+FDYsWayiVVUyqTlfuWsUP/6chhfMhpS+M/ZVGxUW4dqlipIG6VVpxD7tvG/1avTn
3an40s1B5jxbwcZE8WM4LhHQjgy2skgIO4ExkN5cDyrdkaJo6D3WROI/8c+34jHRw5OHquu9d642
RX8TMks2FkP1n5m9mWuzGXgyostLoh/VxAy45er44v/ba2DbpuIIdUoGzMzW7FejMaLR8L/yjFMN
7lyA3RH+fB5bdNFluvg0aFF9T7K8cD+fSb+OfjHD9/kRJrK6PIX+BAF2WwVEfMMwZdONjk6sdhYL
dZIrLrWyXc+eWgFjjcvp6Ny3+AbVt2fF2PViShHc7gNJpJrv2htiiXml/531I+fb6/vHZSFwBXUA
KAaf/avyDNOAUPCZ7p07Tjhi8qWX+P3CggKSuvNxU4JOFb4bO4iGVTm3PwxsDJve6EY6ZqPiu2QG
F2BdZqiPq3fuqVWUbVh6NIXUrwMtJEIdCFbhh2kShuWTuiIx4N6Z+feFDzakd1DQdvzJzmHpsrv7
uo4BJMD5eIFmsZaoSNa0eBLMtX4e0V+3N3GjU8sHtBUTan8RUNRYrSJ3T+3864WLvpS5w60UMwfb
/61+cR8dXV6PK6M4HMQ0oIt17DU102wf6Ty3lJy6A9enF19TElTg8/LfvAqvSTD+I8o9SrEX3ak3
leTVzyNOmGJx8uOP/5dvCIKf3hOIUMFPfiNYZ/SGbCHsdljEWfll68XpBbG/wh4vltuFmsj2Okjv
NsM2oDOcpfEum72tl7kg6W99LlQGhwm35I8wbxNNfYlMx1DC96SUk7Lwx13gDtmV/GGSUCdhQlIO
eVWsZ74xkOylt7FJNkXGSmQq/S3w0VGFtGjDqajrbvhvcFtO09qbSwWdSWj3KHoqqdbVi0HHGnhH
VemFrvp1rDM89JiYlIgu15Hm4GTmi2enyUlWtRk5YswxMQr80Y0I7V4bm4nUJeR9G2cwzIPBK500
gslNPZXDsXu6spczvgyJ5P5p2TJDZkDgpxwjBXvCQrMR3EJnBdOFJk0kIgSAPWhMxwfpogjHHMMT
GLIZ9YDar55uYYMHL0sN9RxybLPYGP46+EdVVEd5b+rcrDUcaSZUqkDx7PuL34HNXd4o0w7dCPs7
GAv7CzB6LCOkDe0iDWQyMBSEP/BoNFPM/fibIZZNePeIgos7b25LcGMWN8Sgh94NQGU2fbvsOgAn
U+oL7f0zmLQu3tpbwn4zGPOquXkcovE6KfN2cpy5sgp6eL+dKytYBFs9boU3GAx3X+KqnLpvd2Ho
KtbNii/YERDX235Nsvy9FCy1CsBTYPmoX7qdg+rnq2NJx1dol3rCsA3JkHnMwCRC2D0HT5OGV4FN
h8g9u74iHDRLjOZCCFLp41+wv3bntcfNPwrKn/fkmhN3wEKahyTxCup7wWy4XlbIsqXkNLiEnCvf
2Auiq8bkeXBRoyojd3ChzCvmocRetMyzdvAq/2NM7uZbd+akc1L0j90f0gGwTN2rx8i5bl3qqBcC
yLMY8hp6w8kwOsnsQphYxMoTYl8yRMBIqOJvkjBTGAo8fm6TEuiYkRUG+kcmaGElsDapxAtg/Ro1
9fVgnezEuqeywzMoikeUZgh3jB4VgmOdeSpvIp8sdc1EVSDUKYE+EYILw/ik6lKq87NctO8Asu82
bFrpg0ZISM0cWlB5OLF/XUJ9CNjQwgDcfDR5ecleHhelEuvVlzTFWYV/q7zY2v7s5lvdU27VZ6Ww
AO4/akjtIVTGQNAUp8GhSs0QDGdGVbHnbwHseTbTWRKHxbDa59QTFHePax80NGF2xzj05wLBxNok
pS32rWWuhIWxeWQGUBAq+UxHECDvwTVVswAvcImWx2yH66VxP5OK4cCmH+1dtBvP2dmiGvlODzjl
+gVW05BzBxrcq6hC9sT049ZEbDYzugpHB8NOf5P8qIPEgJeYtcQXc88jgFndBaNeKwVT+HNjElti
djRH5rAG6Zm+CzWC211nH/VQmzn6kmJSgVVFR1ZAnGL0gweA5COJg6hhVlmmtrJHrOJ5ePO1hVLl
iKuevZN1G/DnzQpnGChs8q7WC9j7iJYbjRZiR4pHLIwPAbGBXtKfD805JF1j7Xw77IygaicDTVxh
R4cyo7DE8+Uk/d9DU2SZYFVGFdk3qV2R5ln8+GtLf1Yp7cu6POfBProqgTctOFz//D31BB4O+Ec6
7IKLeo7IcpJZmu0ISKv5ZXpENuyKFOTOgkCjy3CWOOOvjaZBPWx7IfDYWV/Zpa91zFQD92gA1BeI
8rsCXbRPnbn7sMC/F7nX2IsxzFP/RQeuPRqyI3LcnW4uHzt0UWSIT8UVc+D2t2zpUSd5St0zzaMr
4tlvfJXsT3QhBb7eYv8tYox2x+hVI6UwkBCzkw5TODXFDY/x7NHagoS2JSCJKo+bPKm9UVE/ikWr
II1gESRMLZ/fCqjUYYECDAuPUEzLprb1QsY997McCVXztz0R6Rl1ki4gfADl/hzUH6Fyz2z0oLle
CbfvmcE9NzTplftJg0k7pwYmcVm4wxwsdsspyHeYKNP5u8z2vTRCVvXiYmVEH52bM6Z0oVEynZGT
+EpWw71Xlso1OYvOWmlQc/6KrZlOlL0llc6hlsYuHfaH56XX0NsqFcWTYAadBp+SPnX6otQhkknd
6GIKqCBGr3CklcQD+5jhArsV4yyi1LY7TMoNXSslTfSjUxYL0CnrEGMKQ5KTXlOCM61zMYoED3md
0Fy2lsWI1wyDlFGU3LlC9NPLkMpMotFNfxkLV4f7minsBbibTqiPfKXeQRZZwSuJbQ9ygCEzmLGL
iDQovwWLNB/JkBoEQ4NS4UisynLbGOWtb/X8nET/uPsu79gx7spjbE0WjaARBb9ofbFfmKdXSgAi
VRcVAkJS5TFo00DaOrSnk8UDa0/auq4znly5kliBBKYsptpGdBvsxu3f6Gv+wInG1Z++6cNccPXX
xJIhk7gV5nqoGzCSCnH3tn3TUY2ee8kuU2usY3OgelB8yzXxDmldoXVMDXpBq3o/uSsC1t2KOaWD
HaDQFXkAQliRuN+taG6jKyKTmW99vVLpCdFeb/8dbgpJyw9jxldy9e3UKUE9aGvxG6rnvPiLQ4Wv
ZxcyBuDXSoCJJrF5X4s8Jh6Q83Ge7jZspmWzuB9QNsKZ92iGTmoHkDeMSa0NMr5VbSiTjAFoOrd8
kaPi27wIFJ6A8U+H0WbQeWpZBrc/OL6Ao64AQmK60L/TosNNsQfm5QhPXKbHmqlSXr+/xguK7Ttg
wE1eh5U2m/br9qldQSLo2/m5NHyhY0/VQmNFUQJRmrvZxXOGuWwYYccyTTU9gTE2EOXsmqprBXMU
ay3OANcaEF9Ujht1H6FO9wXejX3AdsavCoKOgXWKk0FdoGz1XrOnZjFcVg51oal1LRu4DcChy+AX
reZBdAjYfqAxrWzDg6Sa2NDBlG26GVsBKMoDXjhXi2t7QjAy0uiJ90/rrr5PY3XYTltjiXeYTbfM
GxKBNn0Qn34aQsccF/sTDlsO9pMN11k/rgWVqiHZVE0fRQ6ptXozi3kfrnr9a/L7d+m5O50rO17K
dvqHcEJB8PT2fdyD1mAYjaRrcmko89Lm9xaM6a8wCF3SWZZDgzOCVc57R84njWKla53bYq7rPnzZ
6KxtJ9WAstQCcMOaMCRlhUHLQec1EFjPoBdiUkT9o6/4zRmhIeDQaoJpLI5l6m5aQqSdin4He1W1
/ybN8vcjOqEcQqNwTmECMwVAmRjQdkw3XGLfHAXqtDESAbU2+R3PE7YEfVPxpGsMdqDXW6Qt0+Kx
2T4TYSkOmKEN+ywBDjPKsyWzDMiHiLWo3XDaFEqL8SVXuja8iAw18nh3Glco7Aa7Kgp90aUiGLv5
XTZRTqyEIlZtFw4wS5MGVvYL8fXgYr9uUQ7RjBi7BBNnBAGDgKmjor8SVdMTKxpPCjtlI33zAyW1
ka9+5Gpi7hG5cNthJG+ortJ5a3eEqQFUQZR55f9vDck8GYE2HhUviXBQ3zRoysIUcTNfqKO8Ijwc
lsmrKvVT4iS5qIAVXD9IqbHy5tKc6v3bt4THW0mhAi8IUj8YU1Uu/j1GOiIq2lG/10aAbynGBIYI
+cI069dPQPpGAxkhWV9FczjF3KcxlJzRms7td3behHtrLEaGQ4UZmu05a+zfpU8kQ89O1ChQBIMO
wvfQgleoYy7WR8JDmmKYyKIKpYYw3DA5zsqQZDIl0lG552wAQ8yH4onXDaAjIkqBy4nXYcxRMdYh
g9QI+phsL9SadogvKoRIS3ub0KLG7VMtJe1Z9/9Xbg9+3ldFD+rU/z47PqbHhEgmKqcFMEwRFlUT
uVUofYlSkrBHQLXFeVZdT0F7Veu/zJnSBf0Wcn/N2CKY82Ep7WDTU5Xc3qc7wU/q96IofzRQ2u7Q
5Ym5JtVm6dDH2HP8Weo75bIkUuFbNeMwGwuC1iXgBhCLdVDLEFwMCBk447KhY+Jhgd5s/o6mHxJT
G/WRcKPE77DOop/ifbnobz6p3MUfQtovtfhj3WSYfxNafFulHDzPKeiQAf5gjIJgeTyyYRFX6dax
c+QJ8JUXueLBRjqapImC3182HzRY51i8VC5Ps5Eg/sV3/w2WdJjQjks4aK7nMPv2XfsSiKmebH+I
Z96Zm4p6hg/PXHabQUQg4EYCrqlUa2m/0wMkvNAbg0w3F2COL6ZHDAVgbJz2F5/pUiNXvjTU4P1V
b5mPbIkQD1MnoGq3evwxvc1Cj0E+k01V9bTAOwDbwbk43Yz1cKoY3ZzOtmPUX4L89uy0pg3Kop3I
W4/NsilCAIpPyf4RmSajHw/r/oBKqS6nMZhXe7KHhk5oZer5wQVdTdPEWwc8Qvi6vi/mQ/XjctBL
QHdfQ+gC5fATdU7svhghv/hg5/BbBobuLg5d6gLqXj9B5z76K7LBqoR04UKQtDUYsRN/LdDyQTTe
d/tIU0+Y9R1VLqqd2tvn6rxpiu7PegXZKJZpA3UcjMTZ/eRTbKaMr6GAUG0xIf3eQxrB2JvmTAph
v/CtQmYMP/KG/mv7YZtSLcakvKgs7wATY/Wd5zqo+IsRShQCrjXId+R8PQBmfBwD3Eev4TWcTFaV
JtlA6PyZBJL2goW2mhN/atpRyW5kFGvck0izEmJrWAfnNxnvqRvTdBe/BrGI3CtO94lf5q4WROoC
f11hiZnXIWrf80ITEDVhWDKDv8QFCAuohiHy57xhIMmTo4n2Jtv7V1fWHmuxYHU/7tGeGRLnlX+/
1e9WvsiW6R345/A=
`protect end_protected

