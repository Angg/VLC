`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 10/20/2017 02:39:10 PM
// Design Name: 
// Module Name: OFDMTxInputBuffer_Lite_sim
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module OFDMTxInputBuffer_Lite_sim();

reg             aclk;
reg             aresetn;
reg [31 : 0]    s00_axi_awaddr;
reg [2 : 0]     s00_axi_awprot;
reg             s00_axi_awvalid;
wire            s00_axi_awready;
reg [31 : 0]    s00_axi_wdata;
reg [3 : 0]     s00_axi_wstrb;
reg             s00_axi_wvalid;
wire            s00_axi_wready;
wire [1 : 0]    s00_axi_bresp;
wire            s00_axi_bvalid;
reg             s00_axi_bready;
reg [31 : 0]    s00_axi_araddr;
reg [2 : 0]     s00_axi_arprot;
reg             s00_axi_arvalid;
wire            s00_axi_arready;
wire [31 : 0]   s00_axi_rdata;
wire [1 : 0]    s00_axi_rresp;
wire            s00_axi_rvalid;
reg             s00_axi_rready;
wire            m00_axis_tvalid;
wire [31 : 0]   m00_axis_tdata;
wire            m00_axis_tlast;
reg             m00_axis_tready;

always
    #5  aclk = ~aclk;

initial begin
        aclk = 1;
        aresetn = 0;
        s00_axi_awaddr = 0;
        s00_axi_awprot = 0;
        s00_axi_awvalid = 0;
        s00_axi_wdata = 0;
        s00_axi_wstrb = 0;
        s00_axi_wvalid = 0;
        s00_axi_bready = 0;
        s00_axi_araddr = 0;
        s00_axi_arprot = 0;
        s00_axi_arvalid = 0;
        s00_axi_rready = 0;
        m00_axis_tready = 0;
    #10 aresetn = 1;
        s00_axi_awaddr = 32'h43C0_0000;
        s00_axi_awprot = 0;
        s00_axi_awvalid = 1;
        s00_axi_wdata = 32'hFFFFFFFF;
        s00_axi_wstrb = 4'b1111;
        s00_axi_wvalid = 1;
        s00_axi_bready = 0;
        s00_axi_araddr = 0;
        s00_axi_arprot = 0;
        s00_axi_arvalid = 0;
        s00_axi_rready = 0;
        m00_axis_tready = 1;
    #20 aresetn = 1;
        s00_axi_awaddr = 32'h43C0_0004;
        s00_axi_awprot = 0;
        s00_axi_awvalid = 1;
        s00_axi_wdata = 0;
        s00_axi_wstrb = 4'b1111;
        s00_axi_wvalid = 1;
        s00_axi_bready = 0;
        s00_axi_araddr = 0;
        s00_axi_arprot = 0;
        s00_axi_arvalid = 0;
        s00_axi_rready = 0;
        m00_axis_tready = 1;
    #20 aresetn = 1;
        s00_axi_awaddr = 32'h43C0_0008;
        s00_axi_awprot = 0;
        s00_axi_awvalid = 1;
        s00_axi_wdata = 32'hFFFFFFFF;
        s00_axi_wstrb = 4'b1111;
        s00_axi_wvalid = 1;
        s00_axi_bready = 0;
        s00_axi_araddr = 0;
        s00_axi_arprot = 0;
        s00_axi_arvalid = 0;
        s00_axi_rready = 0;
        m00_axis_tready = 1;
    #20 aresetn = 1;
        s00_axi_awaddr = 32'h43C0_000C;
        s00_axi_awprot = 0;
        s00_axi_awvalid = 1;
        s00_axi_wdata = 0;
        s00_axi_wstrb = 4'b1111;
        s00_axi_wvalid = 1;
        s00_axi_bready = 0;
        s00_axi_araddr = 0;
        s00_axi_arprot = 0;
        s00_axi_arvalid = 0;
        s00_axi_rready = 0;
        m00_axis_tready = 1;
    #20 aresetn = 1;
        s00_axi_awaddr = 32'h43C0_0010;
        s00_axi_awprot = 0;
        s00_axi_awvalid = 1;
        s00_axi_wdata = 32'hFFFFFFFF;
        s00_axi_wstrb = 4'b1111;
        s00_axi_wvalid = 1;
        s00_axi_bready = 0;
        s00_axi_araddr = 0;
        s00_axi_arprot = 0;
        s00_axi_arvalid = 0;
        s00_axi_rready = 0;
        m00_axis_tready = 1;
    #20 aresetn = 1;
        s00_axi_awaddr = 32'h43C0_0014;
        s00_axi_awprot = 0;
        s00_axi_awvalid = 1;
        s00_axi_wdata = 0;
        s00_axi_wstrb = 4'b1111;
        s00_axi_wvalid = 1;
        s00_axi_bready = 0;
        s00_axi_araddr = 0;
        s00_axi_arprot = 0;
        s00_axi_arvalid = 0;
        s00_axi_rready = 0;
        m00_axis_tready = 1;
    #20 aresetn = 1;
        s00_axi_awaddr = 32'h43C0_0018;
        s00_axi_awprot = 0;
        s00_axi_awvalid = 1;
        s00_axi_wdata = 32'hFFFFFFFF;
        s00_axi_wstrb = 4'b1111;
        s00_axi_wvalid = 1;
        s00_axi_bready = 0;
        s00_axi_araddr = 0;
        s00_axi_arprot = 0;
        s00_axi_arvalid = 0;
        s00_axi_rready = 0;
        m00_axis_tready = 1;
    #20 aresetn = 1;
        s00_axi_awaddr = 32'h43C0_0018;
        s00_axi_awprot = 0;
        s00_axi_awvalid = 0;
        s00_axi_wdata = 32'hFFFFFFFF;
        s00_axi_wstrb = 4'b1111;
        s00_axi_wvalid = 0;
        s00_axi_bready = 0;
        s00_axi_araddr = 0;
        s00_axi_arprot = 0;
        s00_axi_arvalid = 0;
        s00_axi_rready = 0;
        m00_axis_tready = 1;
    #60 aresetn = 1;
            s00_axi_awaddr = 32'h43C0_0000;
            s00_axi_awprot = 0;
            s00_axi_awvalid = 1;
            s00_axi_wdata = 32'hFFFFFFFF;
            s00_axi_wstrb = 4'b1111;
            s00_axi_wvalid = 1;
            s00_axi_bready = 0;
            s00_axi_araddr = 0;
            s00_axi_arprot = 0;
            s00_axi_arvalid = 0;
            s00_axi_rready = 0;
            m00_axis_tready = 1;
        #20 aresetn = 1;
            s00_axi_awaddr = 32'h43C0_0004;
            s00_axi_awprot = 0;
            s00_axi_awvalid = 1;
            s00_axi_wdata = 0;
            s00_axi_wstrb = 4'b1111;
            s00_axi_wvalid = 1;
            s00_axi_bready = 0;
            s00_axi_araddr = 0;
            s00_axi_arprot = 0;
            s00_axi_arvalid = 0;
            s00_axi_rready = 0;
            m00_axis_tready = 1;
        #20 aresetn = 1;
            s00_axi_awaddr = 32'h43C0_0008;
            s00_axi_awprot = 0;
            s00_axi_awvalid = 1;
            s00_axi_wdata = 32'hFFFFFFFF;
            s00_axi_wstrb = 4'b1111;
            s00_axi_wvalid = 1;
            s00_axi_bready = 0;
            s00_axi_araddr = 0;
            s00_axi_arprot = 0;
            s00_axi_arvalid = 0;
            s00_axi_rready = 0;
            m00_axis_tready = 1;
        #20 aresetn = 1;
            s00_axi_awaddr = 32'h43C0_000C;
            s00_axi_awprot = 0;
            s00_axi_awvalid = 1;
            s00_axi_wdata = 0;
            s00_axi_wstrb = 4'b1111;
            s00_axi_wvalid = 1;
            s00_axi_bready = 0;
            s00_axi_araddr = 0;
            s00_axi_arprot = 0;
            s00_axi_arvalid = 0;
            s00_axi_rready = 0;
            m00_axis_tready = 1;
        #20 aresetn = 1;
            s00_axi_awaddr = 32'h43C0_0010;
            s00_axi_awprot = 0;
            s00_axi_awvalid = 1;
            s00_axi_wdata = 32'hFFFFFFFF;
            s00_axi_wstrb = 4'b1111;
            s00_axi_wvalid = 1;
            s00_axi_bready = 0;
            s00_axi_araddr = 0;
            s00_axi_arprot = 0;
            s00_axi_arvalid = 0;
            s00_axi_rready = 0;
            m00_axis_tready = 1;
        #20 aresetn = 1;
            s00_axi_awaddr = 32'h43C0_0014;
            s00_axi_awprot = 0;
            s00_axi_awvalid = 1;
            s00_axi_wdata = 0;
            s00_axi_wstrb = 4'b1111;
            s00_axi_wvalid = 1;
            s00_axi_bready = 0;
            s00_axi_araddr = 0;
            s00_axi_arprot = 0;
            s00_axi_arvalid = 0;
            s00_axi_rready = 0;
            m00_axis_tready = 1;
        #20 aresetn = 1;
            s00_axi_awaddr = 32'h43C0_0018;
            s00_axi_awprot = 0;
            s00_axi_awvalid = 1;
            s00_axi_wdata = 32'hFFFFFFFF;
            s00_axi_wstrb = 4'b1111;
            s00_axi_wvalid = 1;
            s00_axi_bready = 0;
            s00_axi_araddr = 0;
            s00_axi_arprot = 0;
            s00_axi_arvalid = 0;
            s00_axi_rready = 0;
            m00_axis_tready = 1;
        #20 aresetn = 1;
            s00_axi_awaddr = 32'h43C0_0018;
            s00_axi_awprot = 0;
            s00_axi_awvalid = 0;
            s00_axi_wdata = 32'hFFFFFFFF;
            s00_axi_wstrb = 4'b1111;
            s00_axi_wvalid = 0;
            s00_axi_bready = 0;
            s00_axi_araddr = 0;
            s00_axi_arprot = 0;
            s00_axi_arvalid = 0;
            s00_axi_rready = 0;
            m00_axis_tready = 1;
end

OFDMTxInputBuffer_Lite_v1_0 #
	(
		.C_S00_AXI_DATA_WIDTH(32),
		.C_S00_AXI_ADDR_WIDTH(5),
        .C_M00_AXIS_TDATA_WIDTH(32),
		.C_M00_AXIS_START_COUNT(32)
	) OFDMTxInputBuffer_Lite_v1_0_inst
	(
        .aclk(aclk),
		.aresetn(aresetn),
		.s00_axi_awaddr(s00_axi_awaddr),
		.s00_axi_awprot(s00_axi_awprot),
		.s00_axi_awvalid(s00_axi_awvalid),
		.s00_axi_awready(s00_axi_awready),
		.s00_axi_wdata(s00_axi_wdata),
		.s00_axi_wstrb(s00_axi_wstrb),
		.s00_axi_wvalid(s00_axi_wvalid),
		.s00_axi_wready(s00_axi_wready),
		.s00_axi_bresp(s00_axi_bresp),
		.s00_axi_bvalid(s00_axi_bvalid),
		.s00_axi_bready(s00_axi_bready),
		.s00_axi_araddr(s00_axi_araddr),
		.s00_axi_arprot(s00_axi_arprot),
		.s00_axi_arvalid(s00_axi_arvalid),
		.s00_axi_arready(s00_axi_arready),
		.s00_axi_rdata(s00_axi_rdata),
		.s00_axi_rresp(s00_axi_rresp),
		.s00_axi_rvalid(s00_axi_rvalid),
		.s00_axi_rready(s00_axi_rready),
        .m00_axis_tvalid(m00_axis_tvalid),
		.m00_axis_tdata(m00_axis_tdata),
		.m00_axis_tlast(m00_axis_tlast),
		.m00_axis_tready(m00_axis_tready)
	);

endmodule
