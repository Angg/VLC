

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
bq9Fhk0/GLv62Kdp4GNmJBK3rV/b9RTXbbI2h5PtAqSrglrGK5Ok7HwR6EEeSBE8/Z0c0P+WbAFD
zyx0FKROuw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
WpZf+3eiLdpJYbqiIrakT29RZMomGGTcm6ljLiJjEZQDt2IELIyxS/r1BbFUtcgZxmLJxhb3YxI1
ZLQgzUSVH6XgupNWv1GXXxdLr0EH6vhei903utbVt3vE+VmP2fhcGsCOfq7QGSMKGQCbkUjuoTHk
bXwjRk0AR73DkUzgVfg=


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
g2wu9JZ45c6wElXuA1w3VVJRgE7B9dKqOKpad2hq1GxrRtt3DTdcBe3Ja95VDOehTyoDY2JScfeu
BNaERj4rPSpz9eTqvn6ni1KnVzm/5chkJIYoybqMuWD9eHlpi/zQgnmEvVxOrgtJdsQMCE3wyovm
0IuHig4w6aydst4EHxU=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pbjreFmgi/ecPbQe97YwJwHbQ8xErONB3Xw6d/ORb3Q988wgyHCGXou1S+3+vh4Kh1db0kJTEYjB
E5fSNU9tzR1hDPSMJIstpHpTcHO9iXQw365z6oTbmjybdRQMuAr5MihCb4h/KE+rwVzTl8H2WWrd
pchw960F+s92KoiyyKuWUCdi9kd/bF1/5AgMHBFmmvBFps+aNCe9LPZdRGrytTha76gKSEekPpxS
Gz5GRAHIZ50JXkYEpXHxydTz1dTOD3s4qJtrA/5dGreREmtZTngylAj970vudfKhFqPPCjwtcHjm
DLlTipNo9XUMZ7NgeogyQpq2dLX3d/n/5Fo6CQ==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Txl0MWffZrHu0+NsbiOnDFRivawQWjfEPbRTTGQ9uMjcR6If8fL6GvQnz5IAmuNhxhUrNILDKLz3
rBzxPd/PWPJnhGC8/slYUx1wuWNmRF9kK3IEDbU9ptyhPEdUaTI/16ooL9z+ks/bCkgiet3tvCmT
CcSMg+tZGwpWnV2WBteWnPAy3WQTgJjBwAiRWp1JgBCeuze5NtthzTtsilGfdFX5f3xw3Ub8woAk
lsLOCTYPKVbgv+XU9+U/xCPXEE5ZW9ttEy4HkBID5ad635hs77rQVqL6oWJDsLP8RPrpAUS0Zvrm
7brOm77sBE+J4yPgHG0APhrC2Dek348JN12o1w==


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
nNSZ1VwZJdDnj30H3FwwsIQGHOhw9ZnJ+mY/NxGpUOs6Q0mrbaggv+/DD0EbBeGcjM7xGuk7YzRL
WrbwM8iAAhuPwl/ILc9Q2hToNA+s2uK8WQQWWIGPaqLTz+HK2991cPdqD+G4CFauZKZrSuPRlMwO
Vtgsabf7HupMXUf+gqkwQxJP/Z5m0ZuY6KWiMtgYtPhmDusRrl6H8Pcg8awglYP4Rqr+qqp5nw4F
GSQqHtfo9ryxAaJsp70Y2/iK/iuqd4agSUt6/XgDmbQshUSvNTFr9ZX4tPkrXy/noz3sGfl49/KS
MsZ27lS6owSlYD51HcoeSVd1lscGtIs4aZat+g==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 551328)
`protect data_block
W1E7nu//xIqjlUDl4J/54/uZMUIan1zQqbzy5l9xMGT2L0bQeODxbxpNYVUJ395qIGCpOzgONe02
CJS1NtVw9LZ5e+LxDmo5qvjq1G7ug1nedVndE8ZJC5/jKeyONefmwuGXzfjzBZksB5GlI1MjBG9k
Cs2aIDl+fGFBgixCi8sPmF0/dql11KOpJKAJZGR95oSdw4D/nUEJqPha7QT/qVO3rjOrFk+PtsgN
69WP0i/k74iMdfdVHfqjjIXeB5eEcBukt+pgkR8/nqvpbM3e+5gFf8j46fQChiCUlLGofbQzfVyq
Qk5SZbzpDUipoyyRYW+aApQu7J0R8c0JsrvGxQRd8T2wADBcSbPvn2qIS7VXPsulS8azsS+hcZFJ
kkYI3vLmHWQ6I9CnbpVV3iYgO7myv3DkZ6JUHDIdzoLM6q/keYTVdjqTsyxD5ylEKg3h/MZd4Ucn
Sj8gm4Gcd34q7vjkoT7zpQkWlhJJps3LVwD3v9U/Gr+Or1BEdyEaJOA7oA7gHY7LYDTVhy+6DUSR
EBVw5Kz9MCl5X7rdI9gfW8EVdkyMY0siZzDvUJbq1ijx3mYgMOPztTFGooVfiJzkSRNDkhQJVXKD
Nys7Exm8re4NYim0eJySonq0o8O13kTgIbEF3h+lNGdFZiBlVGLIG5BZtx03+8YYJQMciGItS3I2
bV33SItUIP242xxqtZSzqfXSROZkQOq2LoSM2zwsMJ69T4Tj157kdFM+bx6AoDd4Q1Qa5SGfv0Dd
/TxgTNWtExEJFcLvfxGVZzTRsJK7Wh5Ii2Y6X8cywqG2ePWjYAuJTZsBFzOgZ8P4XNT2uFvxcvtH
xiGnQ4ehmKyQ4w2GLAWSSf17mYVJGzN3w2sz+tjOK/iRVSPW0U2qTxTY+CzdauwDCfFduUd4oh3/
8lhTYT/YxdLsbwP3Fc61iaMJJRdDAfg/Jh9GsE744mjfZjYJPJQ+ez9WY2OQKZM3M8q7k/1a/I6d
QaZuKDGHDnITFbAjXmbnizIc2CqTIqivKbUdtuvuL1slBpHZx1um/EUItRkCg4kfhb5jDvZUa3/n
8Gr1dRNQtoC7T25Zl3IuOqR+Naojt8ZN4BNm64x/fK9KJf+2ahhhbM0ABXJlTUHoP/BkbdIVBV+1
0L2k0jRwYh61zRXYVjhgilH2T70zmUTfsdXEYJMg4afGq8tWfp4g6vxbi319VWoOohwBt6j1lz9z
EtAsqIzHmSndpQYA8rgiM6EYb3RoBMcnnmzfIx+L+qYy1JwjN/G+IhEo7YIybMsZKIwB2/OhiFty
TIoEElWjffFr5MAYXOWtcUluc9L7mpufqi3j+DfVt6rkiB0zmZomHwhIcAsNcevgyfFau67jQT6F
ywLMvQuXqwRaoLrxyHa/4C4ANcWmwy3zCNiqBme0FIAfmbCtklKMnGrZDfQJ4uKIvaTroyiLyNEr
YuwQpl6c7uRhgyfmISMFgdptUVeGRaIjjkyZYQlpmOkM8jsfX3ZGStEA3TVpLX0TFjm14sLtqDCF
/nbllvTYxu72a/kRntCImT6O7qzevs2ky1ty9vbDpRItN7Y2qRJItwGHBDOa/d9hKEv2sNTpxs80
LGPiq3lxgruWjiRDBZrJaMYk4xqwLC9SZAq9jS7yLMTENLaDIqyb4BVdV1mqj4WKjXSFbSZQlvIr
UnxLLWZluCFXWIp3ZccQlh86MEZJQanty7M+HOhL6e+cu8xiD06j3KmcQt1/1W//RTVK0W4KScKl
6S99Wsv6zW6ZEmRW1pV7bgzQdSOJCyE12AGBVOg3mYlEsoVgvoXrTIgiK3MV4CAKBa3a9f/Qu4KI
maTREReHxpwTEDJVlIfytmZhkFtjR/SLbDY/JjmsY+juV20w9+cvHZUVBOkfasjIMHtaGffBL0/I
nuVy4ALvz0Ysd2ENCStLVjt8PMawyOug29IlfMSMXBGfoXt2o9DRttdycsLvDssJwUOPAry8uWNl
cLoLmUM+rmHLXRAbAXVY4gF/xf7ElUWrgqX0F2zITo0jr8Cpw1IBXzDc0rhrBBK7PGpoHchzUuZC
hn1g5NDzeHl99Zk3tZlKwhRRF2vPifiCqSLXmKuJ5bjFU/oq5l5Z4ncrh7yZFIKmCU4phvfw0fWP
I2SMK28FzOW2u6NjzPfXhL7FQwSPKM8WFwRF/UYXg+qL2s2NNXhiDXsQusXeSsvt8JZiJXF/D1jx
eW0aDoiWNHym8COG2R/CJI7N0kdAimDPseThkWU5hFysWuhQedPpLAGPTlDuswal6c4Q1XmgSNxy
MlbtJ6F+9vHzm0tHBisClsUzsdBSo3lETsgbJJesxiqkToAPMzW3q2VKxxRfODe64PTLEtsCihLL
ZnS792CpvkSXb1Ppqy5E5wcWxf9oAp6QzyDu1+3hRiklvVQ6UWX27yr0/qSx5vlvQY/8mbqJurHE
EDytXnx7f9wOiPEgIfGZukwFY8NvOCZCCcJA258+FWivhPiVDxu8l98B+RKXcCTitGhcmRbcBlex
CJ2m3IqCT9MesW/e8G4L7bDZBASmdwepAoxyyHEr6jrjGUsDAr7oQgXWQEIpEu1qSZJTR4+mkeCB
3+vk7T3XrYwKotQU4BVukGnf7LUENQP7DV1TByHfCVSnfAjOsPmu65yp+qOB30960wjWc/zqIKwF
YowK6oAkBxUpnYRphmGlu1Jd8EXA3mosbXWggqHLWTsjPBXAwrv8M8XMxN4O6e118s2h3TWlOe93
WVRSAN6G9sG3pRomdpVyVYdzzjqXBd+mcu05IQNUuFYUZgf3C1oJnhlpaD9OVWSu/C0VuaaSEY7d
FTwZU8gVwe77zQ1yvK/Pe3mGKDeMchyRcggp83EZKzBeCsQWSqbPRLsf37zZTT3RdfQbEOtaChId
nCLcGoXBUe9OsaWJYk21HvYxyQ7p1rozRGXeq1YCaR+9P4uqYJL23UhEQ1760BgsZDfuYGmwuCma
y+KEVRFXAZ7c323+FgwhDQ7SqvswVKi1UthnoYEOeDvCiuqHwOYpToxbGt0cavAGL5T+ZVZ7zsvZ
p3IsCDPVMeKCp/3zsMJabCthGSoIfNcWlB9VKZnZRlzC7Xf5mNZfrddNtjBgpGTMAxocZn6zp04F
2fvxUutKjM2KCZ86UafeD/IEXGy0oRERt60FzfldqmFfMNZcykmqnGNNug9A4S5VR/SQyiJRAwZC
38iIxhTeDsn3ihH6fmTqaaBWrHSWSiAiXz4QaG/2B6VAakkpLNdL9YC8vV96w7FI5bcy5tzHteq8
cbK9UR63ykQg9DODiscbrfDaSsk2RfhlMjG9PDKlI9qhEqzK/QTPfYj+SsgdLuiua/jDpnbMtQ8v
G6zSvZnqOCrlptITzePGjOWUygLNg8aDN+u089xRHAMa2HvjaYRM3UT0JGBvhHQ6tn35eS+sIs2p
hEMX/PSp78BxVpUNPcK//QhjzwDMPxkXKttIhUU1bZtuhKoL5bLfnI+xIynZj7oM5aCGbnE0fyvd
gLnhmPnLO9xs0uppdIyGBzA1uAzrZtGEmcSNBE2HGkLxHxHiuVM4k6rx5bnVY/Iw98gX7/g3iV1P
ErVafCurU8YcCKRAacSeVFPDbTGdP6Cb9Msg9l3KWjlRO5sWxL1wCVbD/f3uQj8OVEacXZnVjCHL
/xMHJJu6UKfQcEWL78RwoThyFys8BUfPWPgeKWxLS12FXVNEDkZkPqWi8f4ZL31AYeljxoAVHO3a
nhDEbAf4dWXgwFfWQ37N9hmbPc9o1yQzX/8MyJCE06qwgToviY/vyAtQqRLe+65amYPHGh227wHg
siQ1N/5fXfqTJ3RpHu8wpS4ynDDFJU8to14uFrsFaSeHJmqGahP1OS2ZQUj0IkapYqKCZw7Ia3dM
f+Y9aWm6My/d3E4t4wfnxeOdnNmnmv4b0DOKZ3cQUZH7hJC4x5dqZ7O10HMqit11IeL2OCCbicu1
Rc2+RX2clyqPEO6cXUmiDDjpe/OpJhqu3RIRfq8OyOoG0k3Ub/FRb7PfEgErIc2ShM6mPrKij37O
KLsIXjQYK7TH9E1RhbX6V5UMuT/x2lE98YR6M7399LfeaiEnlDy1WTsfKvIEZAQFIeMOFXa+naTu
XnSHwqsjax0O4jzkvtu4sLkrbWDrtzMDFVL9oBJsq6dSCOxvM66YELYnCwlYXcNteLvxVMk9YI5h
HqoPkbX/7bGeckUuojEsgx6Ym6CcWBr//mOuUlJLzH0C5iiit/bizYJk02oZlQIJg8jVLI5Wi/eN
ieOLtY+dKAa99VrNELzRO4pHfGPf1ajZwARWYxhB8xgJTB8yD0N5si/QSEgpVHMDBLQfUGONTbEd
Ar3BZvsZ3apbGKfx2jozL8kY0TBl+GbvZQ61RXWTj0mGrCA/uF2h7iU0ug/5Brd1SH+ZhJYdwwCp
zI5cxNPNx69fAED1+f6jCzm4PAUKID0/7j7qVsehLMBY8euSMEFWuWFb9tScfs6ltMruGFlf/mek
iRGD2jaSQfPprzZNxOdOGrxopo37Ic2+8rxe1fI3wlDfAsi4AxXZKxum3nflp1VH8SSY5qccxbI3
EKPFmUmw4WhcWdoccmwyipmnGhkOpsZA+txvOt1CWxQvEXCVQ4Vr7YUB7rRYiuA8CiVVtZjMXYeW
zVeUijPfMLTjK6qZ45MWnP+EC2ijFtTfVZMGwlebFFcw7tYdV/6hR+PxE+3sWmSFh00J48KMVwVU
arz4GMBRVx0Z2wI0odsdwPfB3nNBjKHI5AUo6kL3K3M8mXCcMupEIgWvqGIfd65VOQhHliXxwWJI
eeA05d0i83NYtwEVAU8qlVlOG/jvU6nNmIqZf1LM+/kQgSx6LvfdDiFvQWCZtIoc0kaW5Lu5dR1Y
pRy6utbtJCLOs72Z/QFpHDW8TbMGB05wSnzhzWKUEFY+9tKHAd3781yyrKccMCv1XzwRUUXHudJa
X1EHFqvxYu32p5BEdjKDdfYeEx/iM9kkhhveIrqYXFeoZRft4ZplCuCa6F/vEJBHXNMhU+IXFM0C
X+Vnu2IIUkRpPmtIOZvnmlXXmBIItIqGA00LeY+ZTwfVWWOm2cDkoWuY+npZ7gfozBKlU0BfwN23
gNoINRw/aFLoz/9J0fimoiT6NhvgQwYs2/RHYC30FSjUi0/8kUbkRzHh9BwGRiKq+WQhoI1HK9+Q
/L3MQO/LaASmj7i2nDX0Uaey+91bQ74iEszY7T93b0hwmmvsxdpnusN4yZrb0xQeHTSnqCG8PCso
z1BfmxwHsM8hcrUcU0It5WBxTe2KYnBM3K8MwH1KX2MBU5H/s2ycq49729CKjfjl0mBmkqg71rLR
QNWb6VDKYXX1ObVcTz221pnW5uPEdgeElFiSI0ftLlU7YD3p+HCj6HS+yRy3qtuIvWEF8X1hLhxI
0jFLcS1lsoJKR+R3ILggl0HRbur3DQQco9YdaB2+mGtg4tT9FtpzNRMuoO1sHy3vPdM/Tl2wQ4lz
hSpq0jyvlhIixQ48wC5+60bOT1oMJN0vdOzcTcn1QjSHo6L3cDMcntgUGEa/I8XrFLOFYqijmI8z
WMtUePvDFIup5Ubm3eZOqMgfWdsPGxi+5WW0JicNjPenlCvPcbZIpmBu/kLDIyjyY46prVWUMs/t
l/HoM1F/gz5yig7FsSXCQRcNMjA+clDU4XwqxizL1xLI3kDyjKd0q6r319dxaKd8w3rqFUkxPmMJ
PFyqitUlEnHQw8U+QsrqexprRnTApOV7lc5ensztpZ5x+SLzWidz6wnIaOYbSc4RZaUPYzhJcyXx
TbJn3JEEus1Eb6164uIK3ge7cp7Mb2rhERB05zCre3TtR58ObVxYdwtmTat9Zd2WqYE0UHC2l4el
F6w0Zj6YHH1zyPFtKZ8fGfGJti+A7VLG1ap/aJhwY0fLLAJhka+asbJlBltPMrHh5xQUeMyMKkRm
PsCAWLD1LwBCRxJCGtiLS/I369QBh6lVgYJYoWsJIIOaXh+jyYxYOfPRoujOcvi6Hvh6ASaqiKnC
t3CdHTbfxaOQ6oxf2+dzCmj/d5/EUE1HIt+wkifiGfcdcNmCM0Q91ExWGc2Q1SE5TmpCHou55Ltn
TwmLx50SB76Toc4mYmVDozb0V4QT2K5IAdD8f+695lKkzAmo3V+hwS2jogjwQhh8+FS3InXTkAsW
wXQHha8L7H4zKB9ohz1KILjQ1e/Q8cnLL/3uOtw725bXPFfH+B/Lrj/bZCx2cDf6sirCHEfuvU1v
cd+4kRf47z70MGmu6FbNi4lUnatIsFtYp7TDDRFqdyS+EAm7wwg4Sl+0z7rsZhaydyZlIw1HKUQS
LulsgVYPOk7q4EpeHzOwsY6B4KtqilESO7EhM2B9y0jS+UjEtcbwJdB2jOxE7fdP2LW+cwDgSP8w
A1HXOvDDgI8iLDw5/m96Suj2MLGUVaNPWmErwi7E14MFMeA91+1weLWm/ejN/lolID4LqUKWbC3g
z1PwVLIQARzv4ouwdAA885UqG/WkAgeiHjAD3YAmSuUerFz1t05pS+DXE5NRqqCbNg/1+CLxQ0PU
Jyak1K+Fsty07FdzDbEdH0cSp5PSzark+PRDbKxNOjYiGFhPGp1Y+jRiiR/igPdaEJ7lgnDwQOIH
ovLnmcL8B57lsgNf9N4x1frNeCjCKa9JW4n4Robtam+2dCq2dk2Hq8ClKcxrkTA4ZgYUuuh1cQN5
D43yj9OCWPxIUjX7iYO3yAV0YfRlu8QVg02pRJjAYXcB0q11wkYhI3WM1XuHUGlZWgYuVWg3e3h7
quror49ffb+AibVCOvm4wi6PYq/Il2yfAQC5gfd6gBDrfGy3/+rqE4sb02eC2r3VaCmLI1Ah3H5s
we5eH2nx9MQkeDVXH8r1WGSJi0POUBmc9w17cZ8BsVYCP6CKtzf2757VIAork2npLOTQfX9UCGK/
WJJvxHgcfwWHaAKBWrP6mE0kourZlU8vvY45y83uRPaGfrEj1yF4pJ6/2alyKXxSAm8+iz7EUc9N
M8xsI7ox4EYwK/6DIHzRiDIEACf/CGpa8fGQe+cq3MxB9eABXMaknl3JW7W/fxlSgg+ojZs+Akpz
KBivzAx3JOdhr0UOYAvRgJyBFnWjfM8sIGDStOCUq+iKM+xHvg/mMTO1/uYRD7g7p4N7OCLR+0I7
8grKmVN8TtoCq9xqSmFu6RxBatPG3oTA34ScTr5/B1YArv8CLKY2He8cfJvYlq2QVXny07t0Xc5h
PsqBCw0hF8PSolS953/a++k55z2uAX/6leUc17GGfV5kRegcubp4P76JP68naACMcJNfvQOymq9p
9s+/c3cunQUHwc+5NvRulQyuJqdbCdWdI+knKS/dopEXptWDSt1lNks28EhOHckEkXCP2V5DeieU
4FsUYdEWaRr76BUjSaNL4AIMDeGNJwRQJFNMr4evnnp+swrBxpTO0M/gWm/athFxzrA0r+Jz8fzV
C/vn30EN3i3Gr9RlKW432AdOtNsHR9h+vk7NJJgFZuGIkVswp7Xnmn7To12hM3eqE5OfYBEOX4CB
wqHDRZgrDgxLGartjpfu0mTPpbI6x/4/eLWCZeh3Ai759TAi4FVCyxbxh+rkM34K4h6zpUa7b3wf
ithiykNv4acsPpYS5GXYShFNH8bemfh0i18dqMRv0q8YcGg3ktWBdC2GI2jJMQFlI4LGmexXN3jI
bt6clQRGLfjZt1cPFakE6xrBn9kSIOOhnMl7RRu1hL7x0vQSlkQUFqKKq7ZT2MY+lFYqKylW29y8
q+BPUSqBAzMK2YUVRZKJsJJjDuOD0XGHsqvIXUOAhGUh5hIY/GLRIt+Kt/ZZ0JFvrS7WISLPMnK2
+CsM6koHk0BIxMZmWYu23BQhw/WeZ4I3E76senOvUpmvfI+5sTRc4e1GmFCeYI55NVMwTaXd1hWL
BDr2HfD8BD6bz9WFA2rW9zfsjPZwMICSBFLBwVr4wJ8wXJBYmhaAOW64wtybipmKS0wL8aPMDIF3
D3H5GF0/FOaWFp4K3fwPU5vaoQr4+0q3UUFudLZCX29sCkb7EheVSr8q6209za3GHyNjktt+BrdN
PDPgIPQzrV1bzyb7XLkmKd8nFRQwCxs6gcFuUv7Qzk2l5v3hFHsqkrFgpqN6Dg1sbO3xh6yCse/v
jwiES2nvdxAnnzW2NbwF4Mud8Y/DTVYTdfnheio3j+YA2inpzd2D0O9Fv6RNviBJiwjNvQ9e+nh7
8zIIn0DMb/Y+CMvIlioRpTuU5ifcAqq/XEVgyvVuX8H2PQq/n1P81JYl30fkcKbb/HmD+qQ1QY++
nPfGoAxDlfCKhATIiDsRWtwXC2BoYgeZNXuM/N2BhMcfv9znQKIdbNTbdyKUz7Q/x4A6j9nG/C68
Z1Lt93oVHTvGkv3xIXOgMtpYT83hc2BHU4uFq6MHF5wjlfnO8+RkrM7HaIsBiQJlZv6q0B4/u9Od
PttsTfAL6XsKnDbUG0W8oqCGkhprZAkIWntAOeRifuFoArXvAvOyQauqKV3NTcAoj8Ri2/3/WrDa
5/VThPaItIeZa+C7UZkeFFtxFM2Q6v7d04fap3FNLxWohTJlDWQUZ9BgpkAyHfTyULP7I5TsgCc+
PAdm0L7e4ToV9kNGQQPTSphvjdw6iE1AfkJu0s6K+lK6uleISsYD5GuCnxJLhi8/BLQyCnWEb6YF
KbIxoDq6uX+HhRDb1bmn3cjmVXfHFkjyFXKNVIirPifjxlrUVIyj5Pl9yAUMe76QH05n6YDoN5FV
x5R0BuFc9K8Q+KzWkjRvHO/yTgmyJWJqpkZjM4moR/CXJwIGNZS7R+O1TBRip/W8UKr7h//K9Rys
ZfB6yY/DZSERO+jEvNFpi0p07dTTeh4jiERNubuIXqM2YsNHSV7Q6ywanlFNGmh2SxgjuQ5cwkDv
TsqGojjFYYmmgLcAJqGPMKG9vYQcJ4b5weq9UPBybojfDESlisWqcrWXbRCX9zh9W9uAbTMQJXZJ
42+gJud192H9OszbMlbI28y7ro71uo7JydJpYnn58v+sVcC9Rv0d7q9zhimuF/WvkKe5uLANHiOx
sB73imGuB385fOV0zj6FG9RkdRSzU/dj5SU+XQ1P6cWhdYJedZmmNPKdc1Jjzjk8bXo5PJ8DsCkL
YmBs5qsGeHoAbLFL1xeX+YsT3AuPahVsIQ1Xw9/F0/SXXhm1ZdNIp1RGOiCa8pz/yMv970fiOQZP
3WIYR28wmW4D3uNTUXnMnBHSO4Gynn7OsAy1fv+RT3MIUD8ObXv9H2IswTRTv2814GRmkoKmznlJ
wSIgPEK1Z+S/4hpalOJfReyVwTX2II6IsU16/YmIm+qqDbzI6V7W3AkoKrokt95HqnzSsOS/5BCs
9GZPxuWxku8xsn3TOF1ZGKWpdXhbdpFn5rOez/cECTwQrvooKVqWCa0KYXNcLOlu1/2CNK5puRvn
gAZYefFTPoS0Izx8vJHbd8KsxWg8uKTNQkUV/1oRzdmmwJpITKUixI8JceU4OZPIDV/ia7ij8UZy
HPtTP20jN43KfmX2tBk/Q+PDOvlYGXAyvhQB1eRlwI8gk4Xw/BL+3qE7Ua3rbTJewhIAAWGx9IDD
mXE4Oq/M3fZBh0lGKCNIExZjkMHEHBqByNR/dRqBiuHP4EBqLR3C57odTORzpadSvCD8ujpa5+LH
elpR/slB9AonoblekKsCnThNleN3kFRY1kTRmUke9ILOrEyowfEuP57bkFM+9I8nswYBdDD3PH8V
Y5kyR3uXZcmsJ1QqT9+fPK+nIkltF7HJ1vrRHF1KqGZaOOGfCw67jdzE1wDGm981lFgoeBWkUTAk
iGMnA+o7Ca26pJFzEXeu1cDhSZNiWl2GV5IsoZLdpfXDcjG/Pg4+WJRO4k+/VmyxxIfI/7Hbztup
G14LzQNEVFFfrAIyls0Widhd65OlS5X1wK4r+LUBi3TJJm++uNNo1o2nGf1fdowYb0nOIEZ8p0qi
wGVBb6E/8B9yyG0TbDiLnvxrwwDour/ck4k1z0kb4n2nHueq1c89I050PJpvVYsAGD0L0d7Sc3MN
gqQYA3kQ7w1Te32lAU8RQRq5vZe7w0GtYK4GOv03Bwz5Puqvx2pLpcwx3ZLVxACw6jCjc21SXs57
sw9opdEsYLc8JWuxgHglYygTU/pgKeOmveOrwXI4I6pwDoYPXy9QyEwcJ7qNlek7xUoTi8AiGTt8
tzGMTHOgVc6hICRcLi22jhyy5NtRCv/wc43RiQ3s/cTky1ArQO+6LOiToy/ua73Dsu8kL/yrZagV
+LCg/yXG25Lryh6zPfJnNkdYR7Z4j6pwfsHKRqP4vsGF71+aa19DIHmHI0KNsZ+JD9gKS8WhnKVb
rl1PGi3CZyntofF868KwvgslJEL3g/E8nsi8mhcsBgGZHam2wkoOvB0k9ZirNa7R1vbvenQFwOzX
N7Hsc/NP55n3dEj17pG6q0IMeSqWDz8LhBN+52TiON4c5hjG3n/55uohf0fUOqA6MsEdpBrLx3ix
JH+/Y5z9ZbpcpIWjNmFcnGyy0W6PZEUpV/3JlM4N14DH0WmKfUEHgt0kD4aea1GkB8utKpzgmPhB
D1R7eEO7454MM/RdgROWrP+REZtxEfdHdBo+pnbMZIwVWmbcru7HijL3Ed/1B4RtHjj/5BJCYZvS
Q23T+/2vqgf7qvzKYLKSgtVU2Z8DShRTZiZ6o4pGtagoLZT8Gm8GtSEOqwlvtUCqYVchh/6OF+7/
SXZOtntLcoKt6rejvTfQMXEHVPTmt3059Z2SvF+9YRqlF6yfPBUIcrHiSy5bABO7lp7ceqe4hOAy
tXjZiIek6mtthmmUcbIGii2tdYXCuSXZ2j0ZSNz5Gy//oxmgFhS/wsmAKuJtjXLrbkIRAQx8sKDI
JfUl0si3zPQ9HghQR1tC075U+GE7UXv3FLgmpJ/EUyyJdgS/jbjcrP5dO86d8jzjROBiPVwQdvDW
sxiA46IAqN7YamFxibwunTOZ3K0cgiQ+g5k691sqzNP7WQ5MsU5YuQV72jS9rXe/mVcM6HRc6vOm
8tZOujO76akFNngTohDGp4zWG/sqA9LcclRupjblSLfHlykB+TibspOcPx4tiSkmiZemn39vDs04
Yp70S0vdCu9GOSFQe09Hw5P9IdysfXv4nT4j95hAkh7FggJwfi9wrq9KaDQPVVhyi6hhBncDk+oH
D1gF4UtHzHViPVvWiHGr6VX9pRrPdmeN1LkGr/D7KYe9MIbsBF4irp+pENj1Y2VVR+vqrCVOiFq3
MnV6+PtQ47ediUwoxfYxYDQXJNNH2eDiFHgLJQPfwBmqkCru9PJOYOntEqFHEbVsgDYBGwUGpbCb
kulUfWmKYjFp2W5MIOXMup+Z6GvQ3azLwExZsOjNlkCEksxc3AgbYqQGwUBzyTU+FNCgYhr1IJsf
9GkN8mlYBAw4CSFQv1+iAiXTTUSObRd24BbzBhSUrU7V5TRkWIjNF+kxsNmklS0g4uwO4QHzRykZ
ojafIX4RqW4xzDxcNqT+u7LR0kXRMmGvX0K1leXCRwUM5Mqb8qrIv3gXWNn6fwY9xMenpvasEDLd
23umFE/MDwvr1mhEIde7ODygvORPhG2KZCYxfK6EFu02o/EZXdQ0xAq2ywpDCHX/suC2ob37eVvG
iGJg2877azfSbzX/QdiWl4NtVvAeJZskG6dn5kz6j4OiEND1uBsZ7Rn546OsdLy/Q11lWeCvIUgy
bpAHB0sSHxzn34u6d1PoguN36c+a3dIle7zDiaOn+IHplb1jD6IaOQd4sgVPRNvr6RzfwoBFMOYs
o2sfHJRTBBmwA8OOb77zV6OE0DUZXfiHx0CTHWZk9htQbQ6xYin6OPJw9uwMdAQreh4f0kxY6K1J
ImhON1C3aGfZMsmQsmpXB/PHDgOO9blmn6xOSWxAab29qTovYxCZ3pK+XT5pWFK5Fw2XEtBFSXcU
zKDFu6XxbNta3RIIzWpJRbUejp+EBu7ysj+Z+sC06p91Gji35UKqKmz5Yx7NMp0Zbhp6rd8tG5p0
rbmvi1uEmL5Jzj73dfTmE5kb9ugGkSEKVLA8h+ewgDR6tMnpEgbtJVAmEkTy0Fe7dG0KZ0f9Skv9
HvpkoCxuAIXU7YIu6gMF7TYtdU1fYfkAS3/l4Ou84huC4t2BqemhFo3pc9WHxJc3hi+guaePPNMQ
uQeNXfs4zF/m/+DLHfgudgUrP23LDIfiLevzMwiBH9vuzMO5Ztud1cIVghxiVLF5okOJlisyP4BM
0GkzmvUpWLpoPdoEcoG+ln21HdjtOh3BvyWlgkaMZ9cr52I0gvl+Sc+mCFpv13mZaa6pjDVFcI31
VX2CSHv5dhV7Q6CB5imzTF8HTJ/4jxm+Bbis9/TDJYn0xWYcF8IPrwUzHxFbHMYNhD4E9uQ5aMwC
SRsjaAJRk4k23oZUshvGhBkG/RfERED61JUKyDY4lIzfaPsv6ehyT/dtPlqBstPzJ6o8BLlcd6pw
kLXyr18uQqGU1vbKVFn8NsjJk2Z+eYBeCiqIDwrPqlwl8tz/JFz/X+nlIOxRumjhMoJs0W74s3tA
9jhDQewPHg4Ztou9VZRe2O2+Bt9u0Dulfu79nQhB1H6fTgmxmMmlz4rFsLAi0yJZwCytW3V+YF2I
V3h9OdkOB77fDkW0v61evrSrT+vy4Yxe8Y/hJP4bRG6dfLpdNzNIsq88uhyGtPNpPrawWElFXDX8
kQO8qRA2GJGcanlSEmTbexh38mnTFc05DYas5Sucxkcqj3fq7zRA7Yn+vmhqkZJif8O+E4s5xzHO
RrAmeks/3wEEK35tvY96vMb+YIBqZpjRU9sjewDgVRqtqknqwHaff04d+u2SfHFRAhqL1CkVm9yB
LbS2U7JwwEX4IDY9jUSyD+kLqE3qqhTOTNPjUzbTF16spPmOirJ/xk+SUVwrp/tDtil6tbbh0l8Y
11cAtUnK9bdxoZV16+xNGJ39dsHvL0enfmAwOScxB+nX4MVZICZUpUvqhyzdYXVxUZzRb9Poh+Gy
9U/L19ybngB04Q7u/Wtl/+zd51t5UrrWMcb83vXNggO2dPQX7jNwC43PG24Il3ku0Qil94LqVQHI
uRCJsp40Be9snNvVpl+cXkgemUYZ5nFv3P1vsTYA8AIoLgHeFjjNSAeVZUtV5QVE2GeBuy8GsH2i
abweA1lLlI4IRZte+7IVJ/z8lLL7TiJi11FjKbTeEAXK+zSd7hQAylDXgQKY44LPy7wSRBePeVl/
ItOHTqY6QJNhX7bKFurRffNqfzHTaFfB5El6wS3dyhMeoM/vTEfQ2+iKSDGdynuAkxMdhXKDavk4
LCDX6cXrW0YYbnFkvQx+nTyZaBAAvk0nJxC/5lMjIiwyPOA7fpa9zFLm3P9N9LnpWZc/2NXBvO+e
JAMTvQE4Gv7CbCNebxmUlDyKHqTPRqH8a8ElmKOB6bVmNAjX4DI64t6LyqCQQiWvI+MuZGotXY/L
IuTePDk+BLcwaam35MKcwDSksszmtCgbPVPJaW2Sxedcb5BpopUDTJFpVyFKyCv436tFAZv5utND
MZ9vE4rqPMtfDinRdTRg99Eq/JOWh5ke+b8dfbeaHhkbwpUpn6/QVXG5KN7c6CjIie1S1dpSQ1EZ
aRB3kRSa0KF7Byi5vq4CymdjsGet45vtiF6TpXMvptrMaO/cq+vWThAQdZ2HtVjllCJd3CcjB+L0
H66W3LUjPERWiXEUJ7IqHmNC7tJ0aXUiAvGzpzLAfA0G3QQZrHf2nChv5oSDYUHGeb7wY0xqQUb4
IVz0mwgmUlUmjV2kMUNbg8AhXTqsaNAwF1jtp5w8K4KlMY1wNLD/X4dakiSWcKw1D2EZzd9ll/fQ
WqfKv5vJdnZAP8s7CWG2JYz4CuTotEzR641bxTlVXHNUI2UXums9f9FCq44DomfK8ZTmKtFNngn1
ItX0hIN/1kA9v9leFS3Y3Cr3LtkbHM72o7chzkPqRi0h7dKNvjunVUrMNVL+MJzwIb+TlOaxaUjc
CvZc5lwA63mpNXmZGrdHX4lT33Wuq5UcKPvdisGB8oWpkU/gNWWKWJHhVobQMUQmSLZxDs8gC/5N
tWg2s/S4KBwpL+dUMdSrYWzHoseW3F8X/nMbhd/73tz8IPWVMJoYI6Ft/Pcqx+pVYYg84SwsPRYA
yKIyMdA+JbSVYMFUOt9x2S28Ms7o1I/Xr+35IDM5DWj/Uwfwh+p+C3/7+q7hHEBgYTH/Rw2QeQKj
i4dichIyEIr4s1DnhuVwZ8m+yeJzsS8g764JqTcebS3SWpaqNKBD+1PHVNuzOEcGcMJYschBS6Q7
h7ArHA4FnTAPVCfRPLxT/mhYzHyopgbKKicJnSyKNU3rIgpVBC1thGp130fzK+wgnJBxiQ5jbK2v
s2rJ9SHxUimEc8dlC99utrLK4EG8yhDwj154aAoRliqYorx3nN3W5rILuTjZL28Vx+xXlYowCMfz
gF04bu8azAPVGr63oE+vHQI+SDImZj6HR9x2VX7cNx64agFkZxv4j5z+lcrwDlVKR8KG/7ABFSQQ
skz075JCO9H3hn/M/gfcKxMiRVQ0hWF4jDjFBhevc8qWMzTZ3JneOeWo0t8t38FX7MRzd1HbvszM
C2xbAMTPogA26ZFEsn79SU24gJNcLiCguHoQLZ6WvdlZbLf5A3tA+9FrELimfne1JH8v9MQ+wK7G
UZESU7bgzSDnSj/5MX2AtA2fX0HjbopCtfEYJaVQKLnGIJGtbTpDc/RuhiC/BfLneo4bPzIZjZ88
r9oGwjLcM+HaYNelAhjAAcTI1WKgpl70GSPojDDX8EZEfI40rcFPeUXqrSX+/ljttt9ER0qh6aks
5MpswqhHEcjo2/cVt8pIIzqhfk7/NWMLDhoeV5MsgDFo596LNksRADsQxbDNj9OB5r2pBCgt/2BQ
JKrI1sAANYLHs8zr9FgpO36XiN1ronZ+0qLN0hmzmm0TuJ7w12g4fHtccUvgwr7ysB1HNOmg+bSs
dRwBAny1lljO9ex94c7rWy+hDiqBkI6jKFl5yZuofk3FRdnnCAlo8HsLc9Cbsiix6d6OdGLpFJ2R
ErLtSrNc/g8R2tZg5CLwyrtWRJIOLTgNTOhIACdJnCBR0P33uwRFHkAGPcjwjzdDgGz6DKoPL2fI
XWx5Vf+9V8OriUA8VqnwVdPCdNsNsveFU2nrBRYBSkPYd4Q7mBAXrbdRpGPDu58MO3mQY+N+xBbZ
Vo3odqOpI7iD09sSFkilM/cI+rZmLyzryZwo/3XKxQcyPZfU3MG1mAXi7i8SqUe2CZWJORcDlG5v
E2bDrXJ6jwC9Jo0DhbqRGHzkewfCaaWYJHH4BNIKUdlEjXM4GydeyLXTyEpnCuNqyQu1aWqlS2Te
14Mt8J+QEYC2ZzqTWnLvXBR5XB7S/MqqgmSdQ0zpuMFoVWpN8IGaPaAEtcj28puwQDrWlYx2C8F5
gtOAJO2es/6qmYnM8MH/I0VEOA0Ot2hHoz/dwt0pX+zzhWL1W/KvwFRcycjYu7NQCt0sC5dIxJsb
RoZpjet5ciY0/Mqh0GixYev3lbYU1unfFnszChr3w0oAc2kLho1VSIzI8xtJgSkSEpXMvKWBCUQb
mDo3rOsOgzrZym/sgI7C+e6RWmUXmykoQdCmthzO5yCwllgIddSXfoIS8S+wNF2kcnIElcWn30o4
OL1Hx5ttMz0yxwuzYgl2lsfESLS3Iimm2zCzxbnZSm1T2CMxC6+AhSpAun/NTW8tDh+fqDTc+P1R
e2Yibz87C/rMXnhQ0Hf6OmoINay1cv12LwOZhXGOv51dSSR9IYBtvh5MhumdSG9wNIpquwV5/CBZ
jOFBLCJjUcaZgXl0oURsd+TOdf23ip1Z8N8TvSpgrDGGZvWLpMLAd94mAawGyfFYz/0CDHKRgpWE
cwVYAnrDcHeh1zq9jTysEO8PdJLU9E1ICMszbhYaXR8F2OPW17pQ2ligY1Kb2L2bTMC5+ZFw9Hy1
s5ylq1fTmobluPs9yM80V+7ZSe40DAtPOjOCsKBlp6qzjWO5ZFtwvxGWDkGaFaLPdqMHkcyrT8Ux
yDu2IErEW0cyQclZIi6X4Jy9AWT7sZQpsfGEqYLE2WHWkic1Wx0FKiCVWcAQgtfH0+oyQ6Ub4101
nx7Qb9WU/zod1UX7Ygo3KLAqcrTt2MqRCL4HpplrA/l9XE5Ey4lfqrEnOm8nOZzxW274+hvZonKi
XFdQjs99xztivqwjMU2hzX5MJdhxxHpYhYmOM8Ini9YLW63DVyPveA03R5XnkJVlaAEBXPDDiKe+
36p24TtZRY9H07srOpytbnBNQwNMdZJU65X8cYmqKibm7ZAbEtfMSvTqmQBRkb07yZp1GwWlLch0
4QiMnCkfg4xWQkJR+IqOj0RGHxgSzJ6DEDofXRmfc7qZE6xNPQ0PAUlBzitLYhTm1H4ka/t/itEm
rWwUP+U8wiUUvfcZyTnQBqaTvIPEbSZqJUSmdUa+nYoK4h+BSN6PnYVdt0ao1eEZU4JsiwB6xJLC
JRl+G1ZMpJQXcSvG95fbu7RoT1SbCLyzXkeUIMoCxDvSo+xoFntkhULIojTmsiPARd7MJIqNNZfr
3y5PHAs7pYCzTC8qJyGfJcNKWe8Smm9WeAF/jqE71H6kVleZGePsd1OCxRtM/c6JKENyKImeV2p/
cZOiRwpPsOme/M22+vqS9sUD67zUZp5ZdsYD430Ak0PPtE1tY6dU6aXvdXALus5/4tVCXH/iiPfU
qB96btL8j9r1UbQ4XzlAiZHwswxKjOIYtrBiTsTrChTHA+RIuk6fmHdHIAg48B3om5EHiBvs+saD
ifVKvMa75l/H6Pb4g6YDWM6TyB5GxbLOsYLlRlX9F8d5SgkisNNxQu3LmCjH5eR6NHffXWButvUY
GMPdYt29PgcqTq9DJsRCSvEv8cRHSIIlCLfGu4299a3BROnev5rm5u+QM2CkWB4lFuAxA1OPoWJ2
Vfrkw7uTQGgyrXcp74/lWMwMtCNkYvVpr+rH26BhRS9EGFT/9nJ0e8BLy76j8kGeEyBRUQOFLJE2
BFRr6x3gmpLyV7C3qaIQxGXnsU3UTtJqZO9AgnVroOHPnuDQTjFlyl8MHetylG1U8Wjr2LYOlKdb
QJhiqWNAdnGSlkGbAig7e4odiUW20AkSI4/JtqYfHm9C5Iwa+DfN2paYR5gLZvaAftVGDygviclJ
JM3IabIbN0koGr1PwSimp+P9VZAKZkd2EPd9ltp0OCj4uI6m92/s4Izy8TddrNWUXu/+CrQEbynC
BbZb4lo6htOxm/7J+Yy/wq30YnYIRG/mBZTURd7mDtStzWF6GytoWf63B+t9pC/ofIDoz6Hff5oE
+jTvUFfqK67y3g7+ce/iPiQ2W1O5HcSRlSdH77kwWuJ1dUshdhhGRoBeFuwDq4wRRoO8c7AjQ/wK
7ypBOd8F9DpF8jjdEGqcPR0Vf9h1tfOWPiqkWry7uHXz2Ns1xxnYkLqx4di8lj7z7ZL+2jpyelRg
JFt6DZR25MPxEdALsX2XLsrMtCiPzx+QCmAWe9WkXGEcsVTbrTpoc6M1PwDDHvjmXtCft1IjeZr0
ByC7gawSMcTTjzAsjlapIemskbYdESgJz7cJrf2smPxHXtpN5OjCtOemTabLzn6g9oWBU4whBLXR
8cVHrfkiGCwWLPchooSyYDoaD2fHG2o60ItLRLCZG4HVxCz9ViOLBa6EkcLcje1eEdkdST3zOBkB
xU9SY03D/8XK4BK+V4w83h++9QS7WCeorvsmrF9iOLVMUZq0WrHil02t+4A+DTsXUgv/Q97Ed19/
bD+3w4ON5jXzf73UXn3C0e8Eea73OVfjT/SVD7LrDByp22smHBnzQST01H37mEs68DctjbvyA1BC
UXg01TDp1mv6ZH9pkj+7WUFMwX9FaC2Lo1G2WwSpUrsTxHCmFIYBUEb+ys8HhN+zMQW4C9b3rOPy
qIHqCElgvSvyUgyeABvWOemPi8u+u2IVrXk5cHb63i0axthc/BKPfWos2H0JLt707XH5ebsokWFE
sGe5bnjKgNB7GbcXVFBTP8IELLaRk1bjXDdQBaJRH7uFRJdWYyBJ48L5m1jQnsKp8DcJNR7prH5+
axQ3HYmXlMHAEM6I/Pz+Muh6FG/T9UDn8LlG6mH7siTdnqLm6sgqbHyGYl9UoRirM8WpFJOmJOuw
2rBLOXTmd4teYytc27rT+oXM8zDowxA12v0+BjphVGp/710Hkx9Oufmx2sFoHm69Qox7KBuCMEUw
/TnXxtOuM3hAIF9heBsu8DKLn4LkxmYHUhW/U2pbVc447THAj06RjE8Uy8+KoG0juW3kbqvMU9ah
l+Zs+mfj5xzbCmu3+IbptpEKfGmIWJWL6bL1qP+YDmPTPHchy1i7TVY1vrJtLXBgZGvskLqX/nAq
OJRSaSWqkVS6NpY0NKl0kO/Rgb/nKGfz7+2MnOLBWXLsiWTIJIuCt5VROifGHVUP6io6pzVc57q0
AjUN/dTqoaSEhSYr1R/h3SMfGYDkM7M1U8IntdSm1+dM5t4INq3sA9jOJoiJZFHqtwYbL+UdieDJ
LwQStSVMLxfOMgd41R8Fkwhi30aRSATnyn6ZW6cm7bvPkFal6nt3WYqAiZs0VIkQw3MObcqPhxfU
M7F/UOYa0tKi5AWFSyQsRLjvlN8QYKbNcu2KnRODKuwlHYuTOv6HNCNYuqWFvC4qagYXxutfPSNX
sAiHstNAVKNHsXLLEM6wUO1lPaV7ypkjbEU/6jsIClBmXflwz65EY9P1B6//IW3wpgygWeYk7jdl
d2f4baQhIF9gqj0xYr8oVG+DRiOpdsDfMgX1wffrmRVFH1New9whqx9By1LU3y+IvOrOnVKhDSsx
lUGwSDDMJAfj/D5GCAPgSsdqL/1HS5OvDw+wjEPsUz2E4RkwchsHdlNdNdrVdvngvyUxCILl8pC9
EaE8e0vP2bkK3rIrrA3UAK4tCGp0x3trQd/2Jnv5VRPSTl3X9p5+yiyYQXlaqIUltWT47I7xxFWx
oWDtxIKzI5PFeF7gea8Qi+JSTzhuPjYpEx4+IJL4qHv5xi7R6/hXdc9kIDNE25xBBfN1hOSzA8WZ
NVnMnglQB6vQU0vaVhJ7bPLBSitar0/iI4orCthEvR0ywaes/3fB0Q1DWgP0omsbZ/wiaje0cpY7
BcX9gSpPiBxpYwiXFFHXYtZVKGUodQWvPWDoI1ZQgpEmyVlvn1zskbskfLO3Y3CmbBGZB3XRp6bN
NgoOWThLslRySZtWRGzd3coHERT0+cUku5fnuJ4O/tAvxPjf1qUiejM8Zj7a8p9TRU9fzGv7/eFC
MDv1jbU/4UQVFR000FzfTX35/CTRdrRGW0X7PSdYX4pPW46aIYb+x9QFfcZa7+LN3gQJ/zXgZrwO
XIwuOfRVduf1kvlCyPQKDooeR1PjThonwTf+tVt98Px99JbSxvDxaFPy17Ko+qA52jEBfLO/ZGKY
nVsANhhgT/5B0xBZHwdksTbm5CBDZQK4efyYSIZ+c6YLuzMk0eM31J0FvR+MXyUmM47TTw7eaa80
ia8MG0UG+cAd/LcRkIVSI/KVscOMjkp1em5Ixvn75BqiD7xJ8VjovWzXGXark/i5TFMinl7iFcTi
u13PwyvG4x6fyVGq4xOUrjRrCmuVC+z0NQAL2ET89vnxiCxTsknrnU34mPDqxabdwpbLTDg9IrG/
5+DYKgjSU4cTiUvPMaQgawj+ZE6ea9bg7P/X5E7lorZZziuTj9SZRuWKrFa1TTM1hYPsUylksiXz
4XVMBfsOoh0fQMfutUKHtrbzyomKt80vCt2t/+MonBHPPRmY1rmanzzrw6CVlqVm93XeMykT57YD
cBOYUP5QhHDZ2TTsB1PlMMTcCaZO9aGiQnvktxhIQnN+Wn6Zc9Qfkw6WvO9JbcDITY5FYldUyJZU
CVUGvo/CUH6rgscZ6wjP94wPomLSRW0NwR4clQ4ZnwsWbILZ3meVzspFh8pP04NcytfofeOrWZYA
Kb8ulTKccZLCITyE0/EQ4Hf9UTnpyzk343Hn1geLQqOGShnElY56jlfquscRApnEvxytf0mzgAHe
a6Pj2okLYftHos/IthDvHf7K6JfHMBFv5S2XZJnLbKdrC9rT92UwFXyibuYoeqqh8D7m5FWrTAZz
sMCqsf/SyGSPUfP8Qc/2hE+qMFFmxQriHsJILt/ulf9fDxzBl6ECbc6xoCBWDvYT067d7Co4hHRw
Rvidgah/2zuVQhDyqpFfPl4tt/nFmxBXpmhG8qa0+LumhA8LPNXRG0BnbSo3+GfZoF+cfo2RvWFM
Xrq822lI7++9GketEFsB32eHoUuvic0xAo0vPPArgMzUf62MlH4IMeBHsLq8lYCexmrwSvfHtNI3
LgVbTadVBJBHyfevuTtfbP9GKlrpDw7GWeKdl7ampLm8e8XfywDQG+AXVuVx0aQgVjn7PKaLwwRS
Se7VBYUGdTSuBEZd71U3W3oFsz/jmMDj31yMN1/DYZE88AcDQUSqXDe3srHo9vj6wZlOB8qWjryX
scZC2WoFsXfRRBrv8jbhwiYkci/j/M4hdpLhGvWcSTZn8HrFgbupZ2JLtWECmXUskLrJY2Pzp8dz
3XFGEWtwY10N8zY+0KRgpac91wiUNCw/RUI0MRm64XVz5J2eU6t+eWJ2FrTPuc+n4UO6qi+XWhiL
EWGref9ZtDWEf55FSyX+DXamrRy5HQ8VavdGvmw+nA88rhsjiqpjr2+X6H6PsI0Hpi1xhoBgvKby
ntgS/Mx6bjm9CZe8I8WqsQ7XmKBp7Rqxs4GCin1nTIyBSfspj/oTMyo460Bh60NVBsv4ypAvda29
6BAOrqNVfOd58RoGUkhgKth6+yAPkL3iA8JwrvxbrpKAzJQcy8e/UQzL4kzgCSWm69cg1cKxBjF8
Y93Umb69sFL6TJEr/OuUoBcTs9GNc5rMbanrUnrwCLS/uWRPzShu/TN/flEX2mOWz3h0V8yk9WMl
hzajpsoLgw5w1t8JtlOZxvFHU1jpo1k6bS2Z+vEvaIpytrZVF85i8D6+S/kMgamkPXtkdosy77/3
2gugNgIJokO+bIy71kBrsAx16T80psS9hmm3lH9OW7yXVJWl4qoOpLhCLfDfTtDKAWz3C+2vuxvb
AcTbCzgN/o6HFFBmzaOBXwYLVJz5av5/yOE644K0WnvaoNt5A6k8abiyZPIj7z5S0+LXc6nb33WT
Vd5HfxF6krToLHP4rMjeFmPTonYuBWLACC6Mv24mqbqGQfA4Hqvm8L5XkkTpvqDFamOm4vtHs6GY
IlmBXekuWvDYclz5AYvHTlkRXKr9wRv6ZNFi4GQIDr1cducA+llFgbbgsDtNcalp9yrmOJ/6FQfg
cSLCGgmSqCRFPtifVPxfo9mfDhPVTOK1wbZc548zDEp+G+8H3FEchkhjIGAEbWQ9mSz7zdtDxNTZ
4Qp+fOG5oYTDZakWo/FM96/rRoDjN0K9xyGPTPcCKepvyaUC60xgOPbuSnBYkDFmv2tVp1rNL+Ei
4JYqlxIhyS773Z6jRE2/Zt7JVhnWSX0Hp2PkmcevJ3AVVECCzISXnMryeTSQmNOcxMq3oOMlNBok
tHGGq/sQYUl20mKSYF3Q6sTPA7GbDolRI4sXz+wYWoad2P9kr6uv1QjCpJDg3o1i0NsL9O6yW/Vi
MjHX5+iuBPYRvtkjEr3eWVMeiq+ecZa0T6qD4OjypXzhWj0+Z+vEnjR/HRjVe3EyUG7P5+AXqB2Z
2Ho47oVLIpyeWlpGl71akirS5CbBjlv5l+zKr9Ncnjj+oiZQCFCmr+4BiehMb/SBYvOwrFoymYr5
el9OD3/Kg9fTXUwKcD91wb6p5FrYpG84CQuyRi5XxjfLTpWOZ8FWdwwFZGKs1f6Sc8kB/LJfTv7h
VF+/BfNDdWwaWqEHvqpjzDCTVxnFLfXR6ULODc1SMkZJRtAltdTU8kt7VNnu9b9/Qj2WsyLsF3hb
BSiRfZnAbrAQWtJhu+QMMfKdwJ257sW+YUqoIyeToduLVIufMGHZGy/Z3kwCkTaLlH/Pe3Fs0IVM
9XvKpS5uzYkDCHdvgVh2MvRx4g0dMsGtup2KZjHQ+Ahj0qQPmlvhhgjKezY2RV2cfsEll0YwmOHo
o7YQJbB44hFHBVaNYY3T8heVqP/VOFUbTzIictZelsIpq/5YPpYBbMugp2OQKSeRRrgFGnZLDeiL
Q7UX8BcZ58vIXw+qJzyRl5ligry4ZOTdB5W5TUoRMcKRZiPdTphTIwYgo1kb/mLlA9w/j04sp9W8
DNrTyqIq9XHlKWN2TBDY+BXjMFrOEDo+wEMhyoK97rj6F0ALOrhENrUWVTYQcJGp2y38jb2nh5iq
ZRVm5CTj9V4PKfXvX9xH8ItDkZihPvQoV0TigobVxB6OA2z4RP8pJiz3WGeqlOcfjCoYNrucKYoA
1pbuhMTtE0dY2yjT7HE4hquAZzrb3tarW0Wxx2TJ6aTQneSY9mQ3jiRZM7QyW4FCNbZJg7LNosv0
3RIrICazsECgS8q9R2TtIKVvdwWrK4tjzh1wLxyjLxKOYQlNmQyRfDaCIR0qOzwBJmS/zxxmeNAN
qfByls9EcxejNYKBs1lnRc4Wb0IuHOe5pEN0PeFiwhhOlNH/rN7u6M8343h2/Bf1EfxeKuE0FOah
Jk44tKHCUznUTBjV6B3dBRjAk1rG8WlZ+Bzpoyi7mbsgyoaTs0+mS/LODzTMnNUg4Q/eE3bmnl6t
13TEO2i5LZ3wPQ/dr8RfWCFJFaGzMwiKqIr9eSX6rEKniF9/dBBkUvSDneqKaJRQUDPvAh/sQdXz
n2h00rX9I9rEpyWLZsGsqaA4V1y9iRckLKTR7cxzL0vBJr2Xk0iaFEx8DcB6j0gAvJfTbRQoPVSH
YpNRV8hoH2+B+WDsZfnJgwpK6ReJAkDL+N+9FxlXJn2ZYND0TuyQLK0XcD8QoLhTdLPFetPXfsN4
jI54UtDNGw2yfDqkk1bZh4FjaLoClBFDF55vTidvSiVpz3A2zice21KsKxtt8ht1+MDBdiuXvbOo
GTQaohynlNwdPr/mCe54HI0YS7M0lhvtldi32v2PykkjshHeT5iiKNaMeBRnVtweGSafplQkd0GM
s5AeSBSmfvmy0hGLIiXQq23nsh/ljHmR7tVqNboM4NKSR8lJw17/Gkc1b8cQADSsN9FyPU5Srfet
zB7xM4mo7LqgvjbiqjartrQFcN6R+7cxQ2kWHpZqOa6E/ic8URurA5a2YitYLXP8kNa8gtEYOqfj
GgB3X57HyU4rbvAGiCguy5vi+jRnTmYcNbcsjPzAj9Pk+lf+GG9FWIkPiBXMAp/L8TEUEy6RD3OB
hQ4YLfHb8LRKa4vWm8rS2MFQntX+1J5/QSz+RNiBM9+mboGvaK+9NRrvVBROPvo3xI6r75w9F4kr
01eezVT8Ho1y9WL+cHydMp9Vt2fbF2z52wFoc1tWs0m+pGCX5xJI4WPktB49P6QauQTqnF5wmTXK
jnUWRTvwvyT9KGXhTbeA5d32e7c18tyLgbqjTPGYsSfhKb0ruyjLGoKNOLbq7hk1ZIQ5pZh411mi
rZlmO7wl0ur/t701ULsnPcxlYRU1GdvkxTFATYXTzuk7BDnut3XYxdTZ1o30kVuaBRGc2zSZBANj
8CAgeCXjwniPfI81twt3s4E/srVxwZlKSiWIP1ax3rhK5qp0g+ayMQYmbM8YSKH8DS/ovutW8Zx0
+8OgvbVCCj6YxnqaUfWIyUKwwjRHkRirtxAkeByr6cXZ9Yj28u9eWCr0be3xK34LXOdyXYbhqBeP
wfNDOcEmtP1g3RPuMjno5oDxQZhbAAYTSjrSZCmVzRD0ck5Xn3Cxr1dMcGpUPcShRNgOxi7FCg9d
3VMEVA7WydivIQF6d739PD3Z551LzkoStTWjwYtLxWNSjeF1uNAd0MdeZ3kJhmeuO7Zut7mwR7Mt
etsJpXgQdokaBd5LFsyfopNjS29glplFQHCVoAfCzPb07yLY+Is6XoViRtcsN5oNPFY+hV5t5RHE
ChmHq/8e9jjMbefOtIhIXP3RT8x4w8FQ2HAmQr+M/SHdiMzJ4TdnUOW/ztNQvfHY4y7sqvabgIop
IcdQLXQ+n06FqC/KnHzmj+S0PKlvHZ/MSx0L9m5BuBWW46/sVkFEpAjuogPtc2brfJDCYFjqTj4m
TBvXdbjwzVxj2CkFPlFEAEw1Oa9SGXQwJ/85F1aMMZ0IcYvrQI/aH3SGWS70yjdl3r9/nZuI2TAx
WtOOl1LpWDSdTPZvv7Eo2Yvm3/FIp2waTDoOI7A4M6YeQVhzfQ4ws9wVcoKzwNwQS0u1YyyKg8cS
NaYc7L7rP4tl+Knz+wLdJg/5wP1VJJcPGhDfxg8aPnnLxBJIQI7iSO2UnkXgWdxsLlZwc7qRl8J8
XR0Xl05PTNTgWE8xo0/OIuG8JVVo2IGIba3+3n9qZDEEfg4GvF+q+RvTL7XW+HRyJd2p8I/vLjkf
WJBlWsyWn0z+0UUq1QlpFtjQH2D5X59u4b1ZiY+A/TBpEYezLknqn0F7oUWgN9FEVweAVEHLs1f2
zFAkbzQt5I4/ONKf9z5j2FXEyMyYdZzPhGCs4MCfg/iQMZ5IpmrLCyiPUc/1JjhvzCROvgdaCUID
JjTObxZes7z0yFJl9hJbq0fEHMwqW8kx3xH+XcFjjxjUKLwCrkvNZ61zG5YWqVxEiCBfzEo+U4Ym
sTb1CtX05EtVX4PCn/tlQm0Icc+/AyXmVeht8Ou4SYo2uwgQNDzv6uydPV4U9igJhxaDacBp7XJb
XhJtin7XdF5CVO5oO2j2g2LCKiV1zp1P+7E6wvvu6xAGOsLL/58Wq2D69+3kv1laIPsIt2V+eAob
kogxwn/wI+fayjRDkg/mb/VLT0+VQpCK3ILVcyyTYjEBL14GdR/RHEZwgiQGTgPYJ9E5/Fr7gSFW
QVwptT+cBG57GGTc7cv2kCAkECNCgZOkxUUIjd6iyMxVjudIi9HJseqsyo/hP0UPQR4T4VtfL8/+
SEXMRFYcB9RWZ6FyVQnYdOjBz6jdYjEdxBI62R9/TrIG/oWC1x+gQLpoQfM49Ox7Vde6C54hlPS1
/YDDjqR8w74orfokTti2ybPqZ6cEiUIOhJMetnu/AVDF9LhO6w0ex+EO1cUQb1p0EmxyZQhE0YdL
VmPioP/yCVfPF1x35WPgc7/wexjwB3yJeIgMp/TxWgRY2Cx/HBzzJSAincOXQMGlDpOmZBQk/88P
X6iw5thJ22MxBs3M51cMeFNmyVldrqUWaWWTA7jl0uyTAXdoDE1zVE7Cuqse/8lxrTmNVaZJR771
zoVADQ3aa6HEzIpLWsbkJB80RM6IyWeNFxmId8dr9dhfG/bl19ym1tXYsy1xMN/FN+1EL52a3AVM
ZANJBTNIRw9JjjrSXXW8lC9iLo5GewguLpa1yYLre4d2NC6fNzYA4OFKUPquryjD2BeHvMC0+Wml
YJrjLygThe31AQ442Vt0EVTwa8LDcFEJucBhA+q2RHutouyEmCpsYZgLB8zH/4rjXs6GU57C8vS1
QjVx5w9ScmVvu7GFdtF/QFZYv3Awmn2DWIO6Nn1bMieNclv0TRJJZ9Z1lcT7rPLREmiJ/evlcH0F
kIe8WufIWRsb8ldQEqCu1fA6u/to4lU6Ae4sNkYFzo8Ac/Gq8PAjIealImgL/YziUl0Hn3b+QfqX
AXvD1bxUfOQ9XGHsIZgRdf+ZNLhECMjuCTBdybnIH3fpStAXDYIWunQPvIdJe1ATPkI9J3OnoMHK
Ac91pVN79wtnnCYSGlk9S8389EhgupcnoXN6pc9gkPse42Qwgp8kx+0sJqEbdYXdaFNXEXNMKW9i
0twrUPt28j7isLkPY89pU9L50WYiEj5ftZI06JkiNSGXoUvEqB/Wyeh05RRmNzwJB8YLhFbPpnbt
yws4g0gzh3OmJOhn/UaK373Rp2kkiAm+OGc6ZjRiU4dNGbedybfzjzhy1A1lBDgmhsj+zneOCBFv
guWnXBpfEMPHYQr6JjD2iYoCn0McenvuwFeTbJvJwxYxVnB1vVVYRLio2BVFAQZoM+/Cs+bGr51t
rSJ+Hsota/O5CWDU1oM04oTjfsZMFAMn4b3c8L/m/7+rc0xeF2sej/kyM1+LmKz8W9dbmSgJDmK7
TAPRWdLbbmiCKdQPj3YdqYKKV8FLvKnDQufqZPkbiYIb+RQePeQEzwFC8kt0V2qIQKB11ik6IuIs
2r1Kd+dvqZEr9xRd6b1FUE7fiFX+rMpcX5oP+bwcJ65LXYOn0bA91fbUlbfkvyxOU8ib7foks2Ee
FcL5WLLzxenaK681NlH/XZN3ePC/3QfxGaGIr8zaNhHZ+qhR7si2qEJ1FwaPHTuHPpfHiC9HpAjo
tR6tcvK60jYcYyaJ20uVcMYDMhSnOp3iItBNtgWbOy2Zy7nD5CAN6lzFDAQQB2VDo7z0pe8xkcYC
VhQYFxZdDct4/R6YUqxx5xGUT7QXAGnoTn0FUoqIT+jPKGv2Jz3sXhZpxmHd/fKt6oQ61+Z01nFy
ipT9bsV2EPrV+ordiEOOxA7OR7vz8IxiYB2MuOLqLPM6/Ldi+GdFCp8HNnU/nyQXMDCX7A0tVcU4
PRdKp5Mki9dZL680yClMZ4vWulIYmvP9EapkHA1chAkpd6bODPwffbpBhsdU0alvRARj7IniSMQT
4hJEZtgYxGaoED83YjEfASu/qsa+MpTB/3hixrjiTBTTYK1KMkmAgGGvv0RgX6Sj3kH1gb87+jh9
q18nkwZWwcBFvaKkub73PzszBM1aqmXolm4+MbkV1am1mDA426toN47a0EfhBASvL0/n6gRtg3q/
36eiM2TEkdLLFJIPPQBQbIP77v3VnpG+ELhU/eXJYu5s3+g1OZjmDhffkIZ4UQe2UamIbWdgwogW
kKCn/4pSpfaVu8b0n/cUuepQJ1EeU3x4+p/97yQvk4kxC1Y1NRfkJdxRnynNF56hA8PNHgIOdzVN
pObRODQpKAZr5gAyDRgrEUGz/jdOMoeDBiKX4xTHB+mqRnOFDXF+UdrZeS66JM8f8fWEo30UR12O
d1L5PolfR4qEthOa+Ex+42ZXuuuylT90S6BIMbJBleHUpSynGbMkV5syZIxLFBEETW6iijTfUBFN
yJuf5p7O/PfKFAVj82+F7hvp9uUhQwsjeNsWkV6pQYmQZ21r8XscPjtb6wu3/tn+9nIS47EfchRo
4p6AXivKEipWzEfKc1Htm0bep5moX4VJSEUf3hKXSP7sVFTa3IHTVL59hBxcgzTdyy0RWbuu5xdm
LpvmP3lzxsmLcxkPuLUE6Yir1Pgoul9RW9jL8HMWu51wXfCDbx5T2XTIbKFdbhogVZLWTlM5LAdc
WVvLwN+2d/TxODBteT3aLrYhzatlE6kKmMs4TTTLIUiaMtV1OL2nBwG8ww3TlsIhCWLDRVYZmUtj
BUTZw+EVTl3rJ2IV5kww0U6jpJG3guqnEmbCKFrXV7m2ew8YSqXHtiUMcS2S0LcgF8DCKLedvQ0J
eNEOa0544rY97OAEkMiagj/tlWMt7nB/HKC2f0Asi0HDrM0kM6D/Qv+W1vLr9EJwyPuajGRQ8nnS
dsYWRybvSsodD/oS1+4E7ty0Rc3AenZ5NgxsERxyio5JBtzL5twE/MVPT9lzvQaHuExPzmbtp9XL
wgQUzT35Fjlo6yFL0VzewkKwbUzSGKvXb580tZAH368URcOXuB0W6XhSQAdCzigM9YwymSju1G4e
mOLCCcgdPa5/nX+67Zjd1Gb0vscVXPZ/uC+o6TmCdzQCP42QE8MkCDHFnOt0gIf3iEfr47bmPuUb
gz9PZ6DKGc+5KwSH9+2lnOz4NUUHT7QBFFYI6QGN0T4FERK9kmnOGJlWoA/POp/BG0jUpfgqfjNy
99FQ4UV9vpLvpriZX+n8A7Vv7sLoNQkJ0fqgPPxvs7QlvMh+vfOnJRwkNPvbcBJMwPmZ1EsiK6ge
eKYv6w7/PGh1uf/Rp9vSHhdOkBzlTNllBgAZ0YFSwT4gW9hjQOy+ZHJstmE+vu9wkKEaTHFaEdWD
rfzEbS8lYY2cul1vTE9l8jdVM3oTMuAD/AQ9gxaDoPMrFG/8cDx1PFH6Y+eHn3td1de1HlV0H8ks
YqMErhUkThWCAbYvbobcxDZ/A2P1r2BJmMGvQyV9zDoaE6NVqKZdhB8AL6sXBAyufKTpEVk+5e1S
VGukJfIWBMwXXHEkbUYL/Bv73DIvvVomIYVtnlY7d6n0h5/hsQKJ9y7J4Y8k0auVEe5oZpeD46Xr
2m84f/DN+u1knZe5Ma7OsuMPOo0eov9CkmS9Z673eDz+vj3A4i8XXb1NTGSweB1x2+1zkKu9CSql
Pl0l68b4d79q8OU2hAcsNTY11w/WIK0XxJW+QjmnVSOONKHPYo7mtgddGbR5y0sVnNUaB41HxTsW
8RCOQhIzOqa16eQodk6qrxs6AvNtfs46eHWWo0GZRDKWy1Y51GzTt1lqF/8Gi9dv4SlWyUD7D3AF
yppOXCPT1jJGguhJC4IqG1+XnBTqDBc2gxR2O4JDSZvhSaG3a/pSkb7G8XUxF56O+BJIF4ibN0Uv
k3BGnIoMSk/abCtJ+wXWgWHWutQPkzhM9F96tL3x+a6iaoZWAAUjVM8sIppb/igRJox5+jHcpyBl
kbFQUhBHSBIT9mZRnYS7iguWb3wcr4qu8p54GpMgbJP8CWXLoNoN/h+gAXad76ow48C9kkGJur4U
VAzu9j0n+ZR0oiSE4TGoKG7GPaDDx1KGqUfJgtMrJgBsU1nfMf6lHMD5F44jEqg28HVStywfwju8
JoxelWNA0vtt9XMTQojhaOSPh2b+d8bLVUJ9OEuV4mNIR6w0eXoel6gQh9wvKNmPOeT8QfP1L0FA
jRSHeIXRWv/jyw2z6LYOtF+QeijPohMHtgtbLpnJjk53XDMbrvv/JmkJ47Ono9wQR0o6KMIkYKyW
iPiGRrAcvltQMIxC22+2z2f/Djzz/IENPE3ZJ6+99zfZc5rydVcUWi/C/tWZTuzi9/zdU/tpPAGg
OeTHQmnohgzXby6zShYwNSBeeL6VweFg7p5VlYBqFcXAkyiJv4FheM6ifNNor3d2MOKA57d1TWUT
wcboNBhOk5VhRHi6kxSApDVdGQUVqAt8ThKVXMqzWVdnEJkmFSI1Vt7Gnr1ilHO3jARERy1wFcwQ
gk+5iHzkR8EWtvFxetPNIn/pz/0+C95ztH46VpOlFdIgsmvLulXYNn6+daVrffg03dsyfbRIrn6X
DngluCbk4nlHvf/mfSQIBk5Y6xxX0bmH3n7gQFc15YQx9GaFdtPXBQ/OyJuIr75zI5izNNxi9mv9
eevW1ktA2RoUfjPPfpRcCu/I2G3r6At0zibQffwJd4+xQGICImeQ791HJ/VcNEGExbqiUxLNRTjS
d+2v2/yaEQBZsVwoB4IxgIwCTd+zO0iWGCHC5bfG37MEXr1Vgy3BydGb1l3xH/8dTbi7NHuSLx88
et137u6Yjg3rRUabip5ZngKXmEhippQTeAf36ZNDX/hXb6m/GkFkJ0wYzx3TgRJyI89aKl4/XSkQ
JR12uomoy3XEB2Ncgn03MIcQ38lP00iKmwBDhtoUwvnn2S7lMLn9R7MegGEIwGKpp8wpDVyuat7A
rwcT11KxuO9li4qT/c0+TMgkRAxFMqg+EEdaaxtVYbG9/E8+oWtn2PlG2T3MPix8wxpl6q7txj2n
cdy4zMpTB3b7d0vF+NiscuCLrcDhjIDoay7y8/MUgRzEkSiWRjcGSWBcFOKqAH+T0mf1frJ5z20Q
tAILCGoDqkbpkE0afCMTl2cujjfNyz3jz3u6htuiHKzE0bLTUJWoUh784rA54bdCpw1XX9j+3/yn
dDb62mBFHZtVuG3RpPgpGmN2tcAA6gUKluPrWhY2szTeC0cq9Iak1Je8+P+fGVf8Pso6Vd4ag9ar
BmPpjAUmVIRCH+FMomOwSaAQszx+jHcbhiWf/gZ49CmE1ZQhqJBc2dqSKolV5QFSk0OXM0cYJwdz
ISkqESgJBdiETyWEsI5A948TQvygbneARH6N+78xTWqL66unyu25UVmDVLAp5gu5B3ntAkvDeKcc
zwcU+jgyZzDgPMGxbkvj1Ce6fxpL229F4W1oCMMLlUd7CPE19hDmvGVKN7yFG302YJQQHNk/CHpP
5sL1p1VsmBRfcRc8tDhT+kkA+NWJmN+T2YTTLjIsPS3SmSd1eG9bQRgp4SiidDtZSqQ/9+KQZ9Bj
fn846qGo3UALL/OT4lPNDqXs9BsFoWek48mEZpqtD8D7JMICRkm+0HMd7GkiCG52Sa638mlh53+Y
XJpClbM7Vlrnwg9zUOt72njCpLG/WEXTCnbvV1hQrKH+GX6XF5HZ7KkZBkPuz642+x1gYgfGQRws
IV6XSnJvJ5O2Nza1KyBpWyvwTb+V6+BeIvxD6t5XYp87/QNJUJ6Fmr1ZhcUzggvjkSlLn9gJVMFL
hAAMM97KrjpUhgo++GYCZNXWg5j8QMc3IeMHKEmVqnJeaKMi2TVL6p45CgRDlDhbQYoziDLbJn23
uZumuKn/KplB4ZgtaqMSslRMFXqo43XJ77ZQ+8KTxxJ7prAKCLjVmV0a8CPX/50ytxgEf4HPp9dp
rI9YI8dtTVLYk1C3p8vQFeLgdc0CDMAz5zvrhskrMdYKNYDqPrFwyd2gBbaTn1RNV2Mg3g2iVeCc
k/fRHxhZimySf286ifpei3yA7gK4Ld/2dUp1X9kHKZtnHs4YNPiWFkC/ksKFK8RxPMibYHtlikji
mSpwN+tryYHRUItvjmRWG2lGnP5OrapH3CNMiDBMI+aYkyDVSV5srbCgyRMpSVRpvRLQdIy23HIl
g9M+EADYJH4/X8jaRledYVUoOcFc/icWbi+4oar8GXsITh2+vEG4sW9Nur89PDYo4+O9Xr4kC8ZG
QOkZyU4AAewlgFkVBwQojYFIPnu90AM8eZ1fk94REIWm27UINn2xIJZLmYD9hJVjl89j1YhwDONw
Lon2Jwbh7h3Bfcf8mmOiCACft2WU/Ak/Va7fJk5MhGuitA2/DuA/VB5LkZ3FbVxqFcY/E19xL5rB
RFVXxhV7TjBmXwgFCfflfHChqS1uP/ZagxhEVGuPfkr9/h6vd6sDZGWEIla2p0t5jT48yKYLrrJL
XbzUNEOPGnzFyeAtHMLuPJvmsvxy5gIJb8e69/VaLUjBPSvn4XeuYSED0ohCLS33N96p4/Mm7Gez
7DvdRzTFJn9Hs53z5Q+vxiv5M7ouGG3wBgoVwW7rtDzZYuZ1C04O+McZdTBTcPFPgC8/bfUfoaOA
JBX7gl1tjKrewaGG7xHlbyNoEsv/IYTlNdmnxYjDi2b1u6jjnxNnM1AY0XCTlf3VET2GIAtC0WIU
ikSfsUkxfh/J9FzzkYbsX49hKeLz3hoU/w4MF7utn1Vg8WXCvOJGg2xRPW+nyIM+bbbsSsKAE/mT
V/gyblAkjcBsVaSW0UxYP2O6sU037YxnsdwI4YXPRtxv09LsjhlKJPXED/ANIhENM4ki++BmY04d
wzw1iX2X778WuWOiLN9VZMGgNpLFtItqSnFQb82c7DH0VmcXxlDAAFsVXh+tJ62rnidHYwbY5SPH
fRsuDbIKCS9xuqA/D+u2CZPxcHuY8iSGvFlqlkXQvtRSwqqtl8E8wgr93ga6ocLPzWGJt2fVoeJ6
pfK12cLBqMGT8DQESkK8wlDvVva5Ozv9UhiTFa6XD9v7XjjU5DnaNZEP3QQ+UR4vf2n7PQK8jByF
SYADFCZIfuHBB7F8vuMcCLuLFiOu/u71PR+DN95AkFdL+TylZpXauowl3EM/C6Nkp0bYdHXfQeoT
2hlH4ybtsVAXI4Zc19IBu4mpUZ6NDI8xsd0aPrbF+o3HNn87tJx17wNCDjkt1H0NgqUgYdIWCe5w
x7iEAMLoTvlVbi8+0bhBmxdDB3tjdL3m7UpZRMaXYpmEqj/ooZk8r8IWzmXozuNCDRadrcC3VtJC
cq9LT/hGDaA6o9c2G3Xd4XXrsyEMTeZwVpmSQYArtBMFuCEBpalYbkwvFup3PBjD4CcG/nHAqwJO
YAGW2tvBLFIzucKZvInbQ9cbPFjQRG9c9QzGB4bUB+n+qzrYtJnen5alyMpguvhxJFP5QEJo8Vo8
RS/Dpxtuyqhqu18KYtE84QdPF0Ok8ysNqsd5/Su2D0ExIs5zTZF7F1N31YfL/MM9BsFKDbMv8wN+
3U/3ORJXmlBE/PiKnh/oN8nYxUqWCftSrnd2aQljaDokI9bgwrxTZggkbA1XChw6ZokNc3C2Uw0L
pDfRW82MOTyh9D49nmIttUrwbA2ls8DbSSh5+NOys0awFqGF56l64xQb/G3zm5Gei9YQVNP78JQ1
/+DN0IU8SK6pBCEd7cgbh7Ip/yREdP/ABKkKcfJsykdfgCPaYpSKRLAflQFHKRyBDG5X4CUtAs1Q
e2R1bX3zTIdjofnH2MIzMciJ/9n+Xbp/tsOdP772xCd5YJcoXgb2/PDY3KmVqSwj02pD2WMH14XG
GASb1G0jy2QoXUqTGWUg5bmckVY/Ohm0QpvnSM4Wjvbak5hZh1XTT9ej101uUi0RFFrNmCDH4m/C
xE90+sekLP66VIdAPpfYdN75hMx8akaS9zJji+49CdUgJvwEEwIS/+txMGTg4kMGyMKYGMwAYEEZ
ksVU6mgGpNxGqT4rRqKaQq1NlxlkwP4tZtw6p6noWsFqYXHbKg3DyQql/7NIj6MTTFNxWN6Z5jn0
Q3pYC2AT6ax7uJVfP1S3OPytYDHl4D1IqgjeubUHgEr3/UE0lYxms5a1zJ+DYbWJyDbtM6WXKbqI
Osnj0pHnDI8hBxvl0tS0aT1yNlNcAd49qdIdA/Gp55rrreG80wtSfzYP+WGudXKNXCYuArqqgSfv
RldUWG1G5tDkoUIBfSsuaNbUXn37H9tcnXUqHvb14txAfh31vOEDcvyZ5dibSdYIVA5GGThH183C
vWsS4ma7gE2VVC3ebAD4ituec+4jr5ylmQFl2oc2kSJTppiHbBVe83fyL/YTIp7rZ5eXsNoRCQFT
eWpCERa9DiHUbz9MhPeCRibEj1TMmftwFTyZRaBP7jvG4TxoawGFe904HVDjLOtI+s5u/1Fc9SEq
nPW/M0Kkg4IqopGPnaSbU00Plqy9sW8lehA/J9mkiRevLS/kcq4UDRMtNJoeI1BBDN4BO7FeqZzY
2K+pSjvLtzmp43lCEo+0nsVamy4owgl24YO2TCafchJABRdob12oOxy5IpWh0MbjooR0DFKTCKaT
JydXsQqVO998Z3f8wKkDmE5GbOXo0KL2tIaxwap2l2nVi9fejHDGm3yIyKS30lg7x1+txOjFMiuZ
Afs0IVXdBggp6zyCqvdojBqV247FUF5N1IJq6MvtF08/1niYA3PxCnEqguO6sfLIOJmahBYmjnk1
azS/CtDrN3v97vWAFPduS8BjtUeMLkZEfD60ilc9K+35K+yG2IH88bgExN9B2Lc0HWwtMbOYULDL
AHVZ5P9NA41R4uOtXLlYvZXfy6TAkfN3TK1BcvTi8geUv/bc/ISpQxve/xPSo0kdeMYlGx7zixCc
R5Xu2eNMjFfogOGKphuXX6je2QeW/BojceeVjZhkT5/68UCxKkp+dRftIZrk3I3lyNEFGJQccrr+
Ff/XNvpt0kuBOhP4Z7uDn+QSPSRAoYCe7HhTuzDIvbQcdOaLMNtMddm5yAd2w1hyE1x86iBEqn7n
HEGk3Ou0rc56k6rRLvuyB24JUKa7ay/8ggDWoxe3c/IQkT1S+PmPpzfuKYQ6gLpYmolBrenN5gyK
4T4J3Hi4NJCe4T+a2062hEi28v5k7ipNuPmDovVBTk2woayhBYKzjCitsvCAnfovzI9D8sfOjzP5
Nr9B6PXloyqpF/4yxFOQcwH5sJpsxMoawjglReUAsYutj9JjAx/hHYz+fq2vrq6qHe95GBhgk31b
+ad4xIhQDWArlxEDXgIJvsPoZ8J6y30v7X07oWUtwcRu5qd+GE6E4XVPHuLXnO+luNMoDG7uepuQ
fh5OjgwC//TUcdAfl6/tLiFXY8wAgV36i0SvuCotfNIGvkg7pXFhINkB4pan6NWlyDg1BNqN3QlP
FVONAbljBE4rH0nLZAW/epnAb2tdH0D6TAhPDdw5g6X9jgqC56pP5I0dHavGd3OfZBCxXPR+cyNj
WiQR7uigcdN7CMiGnpx2UtjV7tBsq0vu9Zq2KExVa5IWdTdbP9Jtm/0FmGCkl32sJeYnuBKqUWP0
LX4J3P2nltcyJ+31nfGp/Drf8vMFOiNlZwNihXCULmBiaIejK1p2USNqE50DoYVJh3LbGwB86Umn
0kXOcZK5f45VmlwBcVSWD6xQK1S1JEpFU40zVHOcFJ5gsHQ49OnWpEmC0HhSiVr0yPgS2Ydn4wS6
gafCqppQu1N6aoylPYwJeTxyqnrYAtaZOx4BOz0D33gYcKM1glDwYf9QUX0Zbo/8DCdJxT3uCM6c
tETDTs2SiVWNyTY4gKktXbvcUfAegWdT5NUlxezHyyYQhiFSKTGKxJfIbXvhnA74qJQGKDkeUzOk
JlluyrMmIov+G9ztHMy9feTFDXNZPBipaYvWIzi5d7oFMW4davsqqze2vPf4ZG2NoamnES54vbg/
/QOaGe17GbpF8XU7MRqhgD9ee2HA6Tcl2frGZTpUEmwRHQm0eM6xRMRtgCcpo9pp4xVl7mYRVryA
yHMLJ3BEYUKdtJcVYywlhk2AhjapDS7w64mNIJcwjhBcWYPuRDzugUxqhF7KvRu7V5VcjVd4VpbX
//6gerUCE1WhwhnJ3iKVBf5VznWFTtOCVwmjYLV/gM3XYn6wYZygEuKi8L+hV+mJChL0m1cHS5Jh
b4rLQ+wOpy9J/Q8p6RcFgJJdtkRXKfBPXxQ3/QEshtNKzBYvO68ehS3J5uTWYfTaa/kNaTTbJwuT
D+jA48Wsrjf2Q4OsAE9+V7P5BIqbOIXzbiclz2UZAZIKCmTrTjsBiQbg93p2hjC+nPwpBMXSZ2x6
dbCwtcsxy9KkxWcIQbBfslr8cY7ckb4N2iIWBgCWR8SukpbcUr2V+dDkm+hNfeWzdAIQmxcDPdYy
7Lht7XOHRYApuuASC7Fo30yImbbPCX9PdF73FVlybJv/UzbSW/K7Tn0rhoRc19JpvaykJiyiFTcV
wTQlMU8N0TE+Anavk56Kzpif4aRWepiOqs/2plzenAQSgmgWxDLymouiK5UZYOwVPlF2D8BiHWxi
prDWZkvImKSxBfM584y9ado+Y6qcTXOJuvbWWogOY+QRynzai7yxMFQiRKQb8VCp+IBuaF/oM/TV
2AT26/zhkylB41b7ND153i5QKZGuhXgGPr4qt5Ou1fwu0zZZYWegxE0CygDzzQRYFPoLYTE85Ssv
37bKonl9qXDtehZctIq8wUcmGgcWlC9fupjNkLzHR3+amn8oDj7PxnPDR/0MXA/ODfiTEEmVsUxa
1Q/V5pM6ab65oDb+lPxYMmWkRKJXNJcAC3cjdOQtOJRliIFJB8HKRclTMqaxJD0JLMLlACPuxVqe
hpdGojcunAxlZVWzQsts9ZWpWTOXzAsNSH9uM9Kl9r5EBlh90/LiTEVSMtdUjw7Sx5c7uuL5MF6E
zcPSWdleKlE3LWCJUwIphCPJMO0uVfc+8FTx3W4WVJObfE3H9KDLA3FiG/hSLEh7W+KPMZN0yaar
U0UkR7ExilizBuSn835VQf6rNwfjryJbFSKx2mqWpgDdGKVGfGHTGea3jvdCIGl5rcd2M3us7XOS
+dDr6jksa28wQv3jqm9npcuL1VYOxCoriDC5XkltaeN6At5Od+QqGgT4FoMJK+ZgyRJQxYxhQDOm
XSfHRB8kN7M+VkJHJTvsVHU4W1eezH0fcHdqxChb6+sxwtjQROWVrgdMaB7iKbRiaJRpfVVg/lAs
eHaYEVIKc/SJuvX6IIDOt5phu0RzcGzKQ1+dSBviv6LSKqm8m49HVTcQ541q3j6ctvwY0xDzTt8Z
X7BjyHf+7pZNbp9giV1HusEx6DT6rk7D3zk7vkXm3P5dhMAv8Vd9QjY+k7rPuYNWp02ghhwADRam
m61ksmCeLhIzjpZkm1dVDeSf5HeGPQqlxL5H8G1WHhnUhgtWsnLypnS/F6m7Cj66CN8H+ltndJ1Q
8lppyu23SPpSbgm6GBg82po6QgUPl17zQlBinh8CeOh1Hb8vwXsRDT06TH2ObWQqMDwBnqmhlWi6
UJ2MbIPE2l1Jm3J7y/H2gIpjSB5FZKVu1BhXLt8gjl8ipL/VNI6WhoxOJ+brq0Eg6KLCB71R/WaO
O8xGMg8ZZF/6xi75yzWZcUa7Xt1BctUaaEbf6MQybUHWlo1C61xMEglZvz/jO3i2WxAfpgpxeYjY
y/lJrh8vzCba7z0UQkqSgQuiZB6t0k+uhYkIebxJN6fN/LgwCiQxVB5Nc3UyCKZS2VNs+QOnhXWI
WveP7qDa5eQHsXA/6aoDlZBe7MhpiZg1QVC/hY1L8c+48wg8iBpra83GEuARYwXuiSo7KeOzQBzX
JaTQpqHyGeAr9TG9sqCQzGk2jGnj8r6kE0RNWp7NOM21RqRCzPnPvKegFEFzX99VPQ39h9/qNN2g
aCRgnTE9YltQ7HhiLIVA3Pu5q6t5X6o9t/cZtSj+f9MHETmYAdFiD9VWVgC4zk0/4Q6pl1BvUd2E
U2mpZqRhOOq4fpZF/vDwr2QixAo3SUOQPoPCNTtqY0nXjk2MaQiIci8MY+1ntadGvO20rYs3tRin
nRACQ+8TmKf6qI8nWC9hQNaqF7HIeVk5J1CsEJAB/ER/wuI9662DVXIzDqPTsvKnKlghkWk0vfB2
dHW/eq6jHBkJ6Yfk512fGrwMT+Z151b3aWkLsvDnjNId8zfFGz5rzlbrpZKl0X9gdamIxo9OubSq
C0G7/JTj+h+Di1NSXP5020aiOAod6pPajvd25SNalI/DLrs/+Wf9noZqvi9cjFuRCbmf3phEVFJs
/yrjcoj+hk/3ujxeflrkmsXT8dTYlntLPh8Cby09NqowfWEdnKxU0gJ4tmnZdRABFmDWmNSuGM4d
MvwNbpuQ1lEbBL2uCCMx9dId8k0+Ynz+4f4dMTKWWsGFUh/NDdL9TsLFJP3axY4ERmKQh0P6EP7I
2ClwUb5411QoI+9zBMyH/p0Kpki7i1SRrc73YN8Zq8yDb6gbd/iTz+X23BmUiG9vzsJE896b3sSX
ulu8KSlhXBj49RrW9xWnfdODJo6pY7CTUJr3MeCBGGBueuAbBpmmgqd1EYala3z34heftcCCD7os
eA4npljyvuaRoJsJZpRZtHn20520zCiJI5eaMWOmeqg1oejM/R1ha8eNqMGepK77/+fNuI3YtHQl
su0ZUTD0k4Io3+idePrMGRrsUdR6zac9fwEfpDesBu5f0nTyFlm4CKmZHxCq6piHOtgctxtnOd07
7LAK1GR0WfuxNETfBhxw+gpAeTNq+f7fSguiCFe0oA/ZJJUx63pP8KpbVO8tRBa2z4mWPp9XdIQH
krW4KQzUkGnAi4tA7baN28PqT75y8ek3A0fun7yQOMJCFYltv1079FRW8lVJAoxnhE6IwGecopFr
6h1lPPtLuW3BoCrjG2HeajuXWeyB1x/SRZodzOpk/Dh88qbbXjfALJe/JzJK0Sy3KFJYoyeU3vNy
OoCACgQcYlZQj/QMdP7I0xkX5Y55z6qBBDU3LGf/oD1n7ozUOnqn9u02MfvKVPmLF4MEO2CDA4b3
S5ZKnQ6bixXrSW4T0pLtoMhSR5DzXmyy8bZEXGgkv/i3KJlzxK8vvF1VXuw3NNyFVyZY7U8AbpY6
+1WK2yyyl2n8D6Os17RdzB3i3vVs9dJtSKxaxrG8RbO1XD/LdN+vAyY4F5Enh5WYmnn6OOD6OuCW
uqNDo4+78aQ7jy2ICb1w98BceFfxdu/izgXEz60iphHgscrPjpLXY8+FUfjE5eOsAQT5b61BIgRR
3LUBDG273YkpQo4Z/CfULqic59PLcocF/Ul64vYBGr9W60ChNYGSIsQ9LPYR8vX8QVNhLnNoGW3n
/5kcpYWABGWO4SNaBxR6S5Ht0QZhyU8+LyUct/1ZXJ8YqP5FSxk/hmXIsDzZhHdYj7QvFGHhs4rt
Uc4Ovc0YRLqbFTjXaIT0FIJvJ2DH/Roa8tOZGuUKp/yfKtZn8DDcljZf5LJ327Qh0gQJahZKszyP
MntAf1JSP1LJvPqP91j5WvMGvueSemXSQGoAchofS0avx6JFXIpFH/8kNgPjjBYdir9eX3uv0hWj
p5EKohCfzG28ErGK0BN2ti2GZ40xT1kC20aD7pCiklSnDY4pF84Kudh+ntb1XJK949qCn7hwGsdE
tUjpG4NwUfQSjRhC1uZfBZxfTmiSZll4vY5buxKFJvrYGW4Gu0TZMyn+i2DiLDmMpGwkQQ8cGs+j
hHEY65NvVP8gutnfAClZ6tvnepwvmuUifrNbMTcfjyXLhFxDoVn+lKzneR2Tb/U5KGM4taXkGtaE
lqn3Sev/F2dT5UueLJiHx9KM1IuZ/mG5pz1GgijB5vzHBHtfHIeL+2hV2nzwntJatHr8x1aQWdkg
25Ep++XlhrVw7JcP0crd17qJal6XIT328c3MijUPfeyRtiYtGk8SAyG1+vdnJIL3CHkAiJlCvTTw
RroZpZYQjun7yH869bASZiDMYJMvaLOYQJXSNJLNgXe2WU+z7TTq/aLSF4PGpdGWLs4BTPy3jWDC
ACvPe7b/tMCvIcfiyrdvCoakuBNrUURjl0xqyZdEwHifB2hBnZR8wkxA1B4qPwOcwcpb7du7vosZ
qXQxJJJkOcHJfe2yj4264fD2gTukHPjRQzmM7XUG/+IKTI8GXneaAEIewezfG3hrhwXZvdkYNEk9
B37eKeqNlgl51xPpKs9IyInb1SgBcilp23r2yOA4lAQZJGPDo/6bKC+2hl9P4LcEWPcZ5+Cn48Di
OLEPfVVzWe/E3/c0Oawt9mFa5ENamLB/5VE88D2T8nkQ9HKEoSs5PckRwG2Nulsq1BR/k9sFgNsX
rOJM3jRVHmgSrN+vy/rd03qQuICjgPPqWiXvEwJ5UB7V8fUjyXUswCne2rSr4Oc2c39XLJsH3034
VOv2nl/NiHYW/1Eghn6YRYVsSK/RQBn+15s3BL4PU9kYohv5XpWkw2tZBOiyWcfKjF9Tamzcb/iq
YBrYxDbCIAeiapC26GrTTuwSOxRBVjyPO688atfxFjQG/lZ/7qO2H35j+MRREUhhbjUev5uPfI+6
vlOhoAOsRNC1zEMou/IyN5nVcn+w9EFvfqTj5K75a7tz+90anWxLDn4veSkglZ54EAtf/W/A6aTi
qja/C0ifRl6+luC/wSYDJP2eWfWm/9mkLZmUw7vG/nkUXE3Wb8n12wY9ZH0tRlHQGqnsOzYTbL6R
11IZRysHqJiam6YuUEAVYEp/p2slzf8YVAdO4coTyhfRbOvw3c6CF8/6FYKrqIamYFF2sZPZpEw+
fMopwwYjn7XXlm3QSfB+pW5oo5/XEr9jjYbog3xusqxxZyCvc/NM/WH1+ZzdZaf5mqc0tJdrocho
ryB8uAuAkBrWCZwq4jBuUP+e8KJWeDdHNRS+F6urGSPgWHdmu6ZvZzsjMStJpjc2MrJ6fZQ1kmVA
LvyImgDcKms4pFytbI0T4H8WV8Y+/m5ISHY+M5zuoa0e096GO5I3F6BQw3f7bZX/8vSJBUMqzKfQ
OkekGb2NAHrKbLujmaR4RRuMPAyTAanNbc9bJqUflMqeS6NwYViOM0MX2ki5eWx/QYST0UJU0k9z
xyF49SjN8EyaxSKm+PM5H9L0ImkTnFGh54GZOLJRK9snjp4L4g7xVYtP/X3Icyg+nzWyH97M9/UQ
zwX+qG6/MieLSFtTxHMwBNCx49MEHD3PEXBDCk+aAfqSFCBy2lN5P4ckm5Xvxs8VideAIuX3ti4T
yZRYdBnJ6qXCoJpZCEkBbNLEm/dfa62tcmA99xh3Nmg7Cor/DapbBCosSNo19izhG8Fj6Vqd8JyJ
wgsPkgveqssEOmh1/Rn2nIBcyrMiOGP2leitDXTODMnXUQUDHHa53lyXLH0ueXTrQmiLkfN2etl8
KpqmjWKL+Uor9SSqFB/HxI5OO0o4Yj+ykeTAsuNBJnADDSdEXZFuR4eHZTqSMMI9WG3uo4pZf6Qk
O9v7NruWQ7EUyJYeEMUUdjea3O6xC0apotbD7inqeEYThljDvmB/fGMxGxl/HCPnQhFzvmyP4jRT
1PYSheV/CWs4lyEpNbaferVZ9bEA49iyikllR9XJTTfY+0qcK0htGYnpaXpyLw/fc1U4OMgOEAxj
gNnmWzq2zUjmM6kJl0mrjivvQGb8UzfbM7aLZ79ST4Q3ddIQPcx8phaATqNUzVhUg5gaIOD7/mrV
BQC0AR9Y2i/XSl2v8u+cCP5sHnWcWzf+xwkcRebM5HI5emTkTBfgd+0iNt/kkR4szKWMladdT5N7
l0BOoMnLk+bRgrx34efz7vbflxszXgkIUCCc3H5c4TIDJMGNgxH3VyeQ3xAi4/O3Mqvemc106lI7
zTA7+YkRG9gKV7TwfWZuCOCY+LIC7dJ46kz4yOdjPVyYIlEi6c+jTFJA5qWSdqlZd4WyyV7+fLoR
8n1Sn1JuQ6AueCEG2k53sZFWccXOBi/8cIFC5DoPyCE61ugxhbUA+VNOlPXlMpZ4+EHrN4E8GUvj
eIyfqFo75wlQU7H6St1774/DIWYHW+HfT3avnZUGoVT4AY8UbTk5C2SkHrsToI/kTIdEvdocMEvC
AtZYbj831BrZXhT5hpLRmEOSEdj8+D4y6zg+/1WxG8DifCpMVlQkoAnAOFl3u0ovX9eEv6Pl6kqz
Gzud8Ha1+mBaJP17ansRMJVX4wM8+PHgwXYs0W33DtLQtTHVVnfKsR7v7/BE4oHtrxxTB4O61sak
GhXdr/Yn8ek/uuvBAdgaEkR2qTrQOOD3bFCdDiGIGEuzRt8tpkWGzaSYW7YkUpz8YMLmLsRR4aC3
eavO1aqKOVkkPOwINC2NrSyIhO74FhxhNAe/0Tm4IvpsCC+tx5iDfzY5cvKSz6COFserG08beVzS
/Hfj0X+wOI8LQ7VrgWMbM7cpGhMfwlopobu1W/sE/lj99b50mEMuE62z5FfphLdN1wCNUJTCzSF0
fNIs8b/n3WV15uArQk4n7VcaD9jVMGpCBb1OI0ybc7ZKg8N1N3bHOViMuyrZfde8J0AsK8lk7/Kb
qoyIgPuVHwCXGoDYaJdRHNJxarbtTuSRrvrePGyYpXGny8Vlf7Ofznj/n8ukvGWx0iSIW/TbnHj4
zbBxBFtzKo4QOCq51lbgeSWgT5+MnqY4BNIXWiDdc4Y1vO3RJSMu8bPPPB7eXZ13zYzpOVq1eJQL
nStTt4Alxh/z9mwj5b7BA5bEfYPNt0Mnb1W0rY9jqdIqpuwQXDJBBKNw4fQ80z58dbcAp/SeUqGF
GP/8FQjTv0JMKlQcjPbPU+5Y5UOaSmuBLFJjmK7CVmOFrbs1zRK8LC4PksHRXnxTQGIviIziDaT4
hMLDMo53vQtw1KaDqjXF3z3EdPK7eyy0joMLhH7VdbSq9xwwDRdcbNymjSNMarRCser7+Ar8XYox
2z/QZMetVDMjuLVDvMn3aELipgO0RIbQXFPh5WiHxGTsg40ge1yeiap9GFa1Q1WcDqta5V1GKHVl
jeLmpLeBVNE4y6nQIA2tyoQCLCvES1pfbqOONyr+UOoj0b7nECMAvYQEAJORqufLGz6O7lMc48rl
elL5wSM/xgQdfCvRNOtXyAx8WTFLQ5j0K5iSHbTLSWbuWd/Jq3HO6LxZZvRlKg+QBSDXXyB9EQZV
Md69dpzevQx1LsSeR8m2ej8ffYMGwsuoi+fctgxMVRghnEWXlCjIwg4MUDgtqyN+PcQ94vFS488x
kY62HTaioyK1u1jn1333q14BtbUXTkxIsehIklq+DcfUtaUKwAZukaep0YSWsCk+GooAte9Gftlo
RYDoaHZbIbYV6O9SsVbgkkzIWjXf24PwNBlAFvwO3oSwp6QiZ2HYRsEQTAxZnWQHoErPioQLC+Em
t0nY2zg5XiteY4Ch7HtajqX7CWTWVTDhEy6ei04x7aOkz307h/FZCFoQD/5BNJb9VLutdIf9JzR7
sjC4mTJ2zjdUteLvW5Mxnl8SCqlJu3hZLDnYFlC1Zfq/ziNnhHWqSx+5O3zGcQdSWiKnj3znF20N
okKV3smyKUC9mHpf4f7COtcAwpvhPsA7Yg1W/StSvY7mZ1v9atJbJt/TyptF8TRbSDF3LZUHyGSM
aKH229hU8WbOhAsWYpptuCsRwPhQCo3Sg1McUNbLPTQ3a2EIoA0lWhXc9u0yo9+amNqtVh1p5ruo
xS84G5Qkg8w7NusYzjdmnrEhT6oEF/2wCTLQYBov2IZMlMZ4IfvjY5F1rNRGU9CF1BdIFp0t8h76
1ERoPFVbatajnlHSUGVxPvyQTffpqUElpa7t2UPa9OQciV1MngIo+4SozWjRgZaHuIXzHngS5nVU
TweXK07pTRMk0pNMpw4OKzr1jaYcxlPlmwywqugD3s+16BarnNoG0h1iE7NYqq5+se6J8lgOi2tG
U1WM6QbfQZfIkslXAZajPMUfs97DzWPqrmvVIuy2qgC3/M09ba7l7XH3zfYQgc1717CRHxgLxDbX
MI8IQ0Bs9jSEivQ+e3MzVjhKsYL/LAcvtiV2LRJTorGG73mr8P2ym5BPd0ddvZWfNGCquzHBd74z
/iXyhV4QghrCrQIiuc92zQ3B83uXG1m8RQTmszYx0EkmFJnOZGozIL8AZY25oKd/pFyWWtR6h7Zj
P1lvmiXf2FHpNYpSYzri2JZ1tjNcjsFanxgukm8qA/AprhcjJ0Cqjr9TJKvh+MV2xjYaYKoI178D
wx7g0x1x5KzQyYErohmt1eZ1BDPIiy2XxUu6RGHi9jQJXSi8F9MOtehbY6IJTxqKd1CGvg4SxgXS
IYP3x8MDfksNVb/SpGuuNnO/1qW5+i2ZNvvDjV9dZaoPBNZdx+6sqoHBVFtUQDqna9T8nlHIl++C
s1Lt64BO5N1zesTiI9qjwtEApHs0mi3K5GVFlYZXtyD1WhFog+gjXwffKCeKYCKuMUxkjnPwkx0H
gEBwPjZ2dCTg8mx/GVRg46LbFcymiQPf2AeoAq0LOvVYiYLGh8FWuwFO0EJS8tvXOgxOkoYG9mkP
vn2InfyHdLhq2070eB5MB3/NRhba7SfBsubH8iiXLAEK5YtJapSdcLc7qwVN7uGPWPPHadSNAYaM
h30Q6Bhej8Fe3V/7ORY/VKo4bAyUStU17GfVKwwyKuSaEqwd+AUZu/1mjBOoNW4bnEWr/nBQxP4s
dUAnMa6Bg0PSYZ6MHx5QbfVGKntcYfwoJ+XEeEMnY9vgvxCut1cYjJ/nZcKeVyUEltWuACbpiPkU
/RYf7iZjKYZqW+CaoWZR6h9+t+3xHQ7yWN1359tzyfWAk9skETZY/SjCqFUJUEo3vuCfW+da6GKT
glj+askBaExGI6nA7xtpsp+PvEkqRGrYwGtU+4QwbAWgE3cO6ITjr34fOl5ayr+WL/qcCNjz1RU1
iIW2V8H/BW6Guw++83TxWfRk/KUJAxxwt9quwwqs0cYVIePsGKqsdNg6ofKZh3g+z/FOf4bCQgnS
rC5872VUu6LoZ1sqTfskOCZwilxZhwqvRyfPAyCIbWcnzZZNoMwIHVLW4RIGUrDqGdWiJNcRdn69
PJZak3OYqzobc2r+GqnHbEmOflpHiI2m+bWd3r4PtJxPt+yKKoeXzjF2QmdZaeU80NhYBZ3lhK8G
APFP7+nGuK/Ut3THegBErLm0xQD5sgY83Zo4ELrtkugVqjI3d+r2eDvrjzErpzRDJCdI9pUOW/VS
RXBsSstYAsR14cszp3TdbIxgB+fzEJgJDSIsRBGPiGdIERUM00edLFWzOR4wG4J1IGjMd+w5rl6S
N5e+mjjyD12TrOD84/u1LI3HR0UNGE8bQnd9RTA12ecjmdzi2gDRubJszGhXxaAFjmeTDuKWxrY/
vqRroP0Jq9ldNaWEwbAhxsBt8e31UrcMQZdtR5s2BS7UPe99nlq4zSR4tVELPTRdE6B763Mcak+O
R5HCIGUo8/9DlflZ1d5Vvh57opmymkXCrGBvLwyWr117DK+csbn2NuZH2+rrVC/tJSVfkAPcW9DJ
3fr4kOWXW0o01ucGC7kKUIVemMaRs6Cwxv3t9JBp0NNwVtbQqz122kz//+gdP3NW21ok4u9059cV
nFb349Binot1otf75MIXstp5mtqN6NxrAdmC1aG8t5Wm/LUD5ylAcLNWXuiNi/JHmlPZ3K6IL9BM
EmqxCVCLbCD20bYNUv+fmq62mgIY8oyitINr5THwoE1ViuIPribEH/qDTNmL0tQpBag0ZgAh353J
sxjy9DWuqLicyUG9hcFwRqfCd4FWKznncPI924af3JoXnBSlail/wHyezlD5GeN/cgstwjqpjf6r
q0waGwdzliV8/Nze5UfGkHY4EFdyVuCo+LrQm0NwxTLy+KulRaKjEcj6u6z91NX0xYIk+4Az0T6O
b51QNtTiC1Bi49Ly7mmKrQ6ZbYVXlAh6bXZWo1Sma/v5txh9qm2SEnMe7rAFB81li/ZF7Srj6tqP
aEkzO9VGNeubFOX87/n9EHWY+xIfzv2yFmQvPQf8LPQ8dc1pFai0mWOBW4edBgtk2Z5VXlw5jw6B
Owew/lPqDlgiZzf67I6KdeKMCc1eRL/iuSjKZ4NLEIncDYq+s8EvYc556jNLNTilMQCWvgkq3nEC
K4HJ2pGN+ZfoxG2dTeYnTdu8G/Ip8zO1vTGL/qIF5NQyIxQYKoXlSKTURg25RkBs6LTB7X2J7qPF
0N4PAC/HzMl/KQgwgBexImreyUMb0UyhpRlUAoUSeBY0cde9jembhmctKDOk5tBxRey0BQKuWY7v
x9OFCl/gP+T9bXf3RUhVdySzwJYD1a4adotCqTxzhwRMgCUkmzpXioiYZNJiFoYgCjcVq4qN1gWC
R/ou0o8QDo/7/OxodwMWmao7XLfcVzkVADe0vDs4V3Bv/lpuyY4MTfWtdnXGa6i3lFKH2YJN/XXR
5hyN606f5E3iyOzBmQC2QGWr9r2EwZXG0EZpfJ1nVTPFUQBZkpkXn/fTVv5UXJGA5VWZbhS+u94i
6ln2KvkR07rIfjbpaZFK8Uv0MZmeKZhA3+QBg0orRwmUvi2Fg56DGC9cvYvgRWnI8tpgj7YxJioa
vm09KEdkK54H8jvuLVKOCKpTG/T48s4NjcCU/KMvPtOd8/y/OHp5v9iREbQmXc1YbNx3uqs1/rrL
DUeUKdZBFnK1rhwtrvJl1Oy190WE4VRvKWu4A0v+tFUnpj3igT7JAwvKoVvxTcsy6v0zj04QYcXb
+6BE7WlJD9f0cs7sN1ch1/0VvwofAIosJLQqLA+X/YBIX5S//tmQNVoE2GzmAil/wNWSfVJOAOET
eG+fXRwniAcDgnHRtYCaYHoYkElvgS1RuaJ9rpgXTb3xR2b5uwb1e62ezg1obp9zb403IKwSNyVW
Hyx11S4refrdvdH33LPEeNNeqxu9zbe5/OdQJtKmmMVbnJbooZg7ZQQayMLXld6uQNqJ/YkSHwW9
VoQFX+VRgJQJQF/vrYB+8Gw9Jnnv1Wy8NeDvB0di46UdNs26w1uC/t5STk1EfwOvHSo2M24ONBQ2
RZSHozhJ2neuZVIH8zzP8UFEZk7op7rAgYW5OxCi/qKCLXZpUGx+LcD1hWv9rby139z2CYuDAOh8
6wkEY71e5m0yYJ+LyRPrnsDBBMO8Kh9ihPOBhHJRZ0244jikGjV/cUPp3xZzYEL9KqgHymMUfeqY
/U1Xou7nT3MoiB1ixh3NHucOD7/skdyY46CS9A7RTKb5n9KMQ16TTukltWUCXkm6Sju6DNG01hbz
58ZKVPgJs9t6iDbxY3fDunmP13DQSl1bl46kWH/6pL3Xb7rTA06bDi7GPOIuR3IkmKSNz9yEJTaS
zcBCL8/Bm7abUmiq8tzaWfGCRZTZfafYXvXgrOpkCD++0bRUhKks5TVeTkN1GBJbHjYDAG8d3goC
WbcFI88Q1pAYs4AA0pie2I1zYnU+1e50EPlQLPdAUE7Jnzft0dmtXyDefUFW376k41ePO/OavhmO
NjhMEOtlTjk5PwcR+jC7d+9QQ6sG40ZLTRh/SdoqAmtlrFRNN7Nv85gpfE8n+zlO4KPqQkcBvR/T
VC51VdSfaYrwSFZL/T8fyIVVVPtJPixeqo8oSkKsVmBfR1ppOhgrZmfF3bV1hsHiEpBTdj3yY/pM
8K+vtai8k0eOPS4CrnwDEDW75aXMA0J9VP1roWIo6uMaPRNbTip7iKVmo+X2j38s4OD/rBQRzO+R
vfGQhX4EAn2VqHqRebF/GooZuZ6+vRLLbfm4r6ccMnjbWYBvUHYvnb/G35/kxRvLbH37dTV3tNmc
I+SEOlShvpq/7js8Su7P+hNzVvEiWno+d0neymh+LWYqVEBMbIC0IYQl8yKzm+mHrpTGIRCfnE5x
ObETryJos2Awj7tjmaf8jXkwxYbd2dctvSHvMzNJ+CEzeUFoKo3EdzcseZIN4SYryJ5q97hnh11W
ElFZOZFWndK7j01s5KTMtvm7sii4+9JB4lX0RSnF4SnjZxq+wWCp0CtQM4YFxn2QX+nm1wZByE7b
rrvYV1jrdowH/77BMP8P3Xq/l8tdrOsAUAkjPcRwu0EQVwY+PRHxEJwDPlL1gIUE36vtHvSTo2lI
LkFwIQbF0XJ6tD/qLHPEbbNY/jmZIDzq8DCPnSt3VE4GuateIzOczGvC37h9XPmnMsaIV/srk8Yh
W9UxyPMQKSbbWASk3N6dUcHQ6vuGOSrqNDoD1yOpJC6AzNJiUGi2mT/Rx3a6DP3TDx4Z2fzDEzp2
N1/dHAJK6qaEdh+pF6vJx6+YGR1neVx74E2/yvcTYaLndeDMW9cbofStfsTrSPs8uj6tiDFtbFe4
OMz/Oq8bMVv/vssA3VNBNfuQJi7j7F2RgG3lJmjZE5TKNaxoPdaV1magMNMfhUaaanoSly0LgDVe
X7EqVbecXdIbS3zTmlhfuz1Cg8uBu3M0+as3A+RTx+3rNtDNDDfSRPelXLPjt+LpTHgVqIa4me6V
C3nmwVlrXMIq1ihrFERqYGUOtWhYspT70jX7WekNjWdijGelmMO3Cza3ehKruoJVrWgnzHgoa4Mv
IMFLgDPPmnD2IxZtmHRXf1BJTot61t/kJLWo4UZ5PtnEVznb3qc0+IFzdze94LQBLc1BbwVn9NUt
/hNRYcTlBldJuQ5Ey8gVudvTtVKQcfS7onHczAZPjnruZSJ+O3tYlrJwy+SrS+DvOVFtZmDIghSL
cXS91oxF+NAfEuW4KjQsil8WJY8xjIvrXQi6mTiVxSGYO0x4sWPXGADo96FXufRvdV6AE80kKgMX
XsHBE7TVu/mvkOOZaBgx2Cuh6ewKI3QgG2vhavzwgLcoH54Z5fa32CTKJXHF7ODOtudcScyPlbgE
5GEroNA3tKJFPGTvC7PF6AQmMQ/qhKgkQbEHISikeEBYt5Q1mdPmempQHjrhSjqhdGbdGtp6KCd7
kbMipXkMHVLSBwln3pkY1acrq9Xf3VVh8K4pqiAD3YvlMZ/qAulBEng2J4Oi3iSZ1Qr72oKU7teq
9LXwjRedQ5AyN/BATZR+bwJA6hApp6EuVL5OmpXdJt6Zf9y3Sp5cuBdqI6BogrOgey2HFFHrxltI
2SoOSLF3QxFjtxopWNHWKcjhA6qUALjoaDj+f413D26JnCOUfqM4pd/hpOJoEMipMUwrmGEdZhnf
Lpa1eZhQgYDSO1WhM0WZtdRw/1P+4o7k9LnDBhI1kNARQNPWD4Zc9g1G7CpjnIC5G0/JRxOVEx91
dZqHZvv0VA6t4pwEaHwc1I+wIYgjRalBbp/MfpAuPrQekCWemGAMOHxHNvh4856rlDwcNWSaKXuU
O0Op2YKxSzjv3C+liodkrhzj5wOW7Qn0TgKk4c6DiTiC7G8GU7th4dJwKq9aFurBN9e9HTm7bqIx
7whhdfk1pXHQA8DgfjzRWcRgM/gm+pgJBcC5MycTFqiWrof75XFQkGqFhEyy4e99Rp2zwEldrtj3
f/l2qDCRbeCs+kiRmSMcSH6uCMpWeSWkeQilBoPNGxSMHGQ4l2XIRYXqw560kAT1nLF8ifp69uQP
P27oWsS7HUmPjoTs8Zk6dFi98qdyu7CF9A+xYICVvP1geobXLy2+G/3+X2lOw9VPpzPYYSBjEOhE
P+ZyuNY2iyZFCldZ3d9E2eoNdOzSEoMlk1avI+IJoDuU5H9MKa8bT4L7SrLJ2drkMhgKszW7jl2Y
xvngRMwmo3zBWkonjBNo7Aw8xEltKe2uI/thXgsVbyz3IYemkaMQjrBgDBe7hY8C4yDUr0byqVuA
t0sXpt0WB+3VMPNBtE1nqw5aBkyo6JTmiGCwxt2XBso6O4WAmFJ1m3YG30cnaCs51D+7P7RBCtVe
bJrNfDkO5wvXoa+CxVmFG8xP5pQm6t/6KeZu9wlkk3AIdoVxRwXI7I9y/Eq5r6dBDps9CCkz00tx
Qa7ds1I9S4/ySPXfOAvvv5fAgDZLLhXebzXopti1yj0HrjPg4maVK4KS39C9M6ZFAwefMi3yJ+Qe
9xUUQ7P5W/P62PuAryWy7Gvia574+w3/7ZvcB6zcK3wq18C7cpW+KiuUxo4pZUEWR96XQ8r2rT4D
C8Chp8p3qLvvr0qPKZF4umqS3+nJJ0EmYlbBPNryJjfC3GKHPlCE7UYC+YPuz9YL32ZI7Q3TM0nV
FigMxR+OU1i3+/GJLQ/gMEZWkB4Dk1jxt+MS51EGM1f1XkBa1gsL7SJukNoINaVmC4RuscUzQ9VU
2x+v0O5sqTA4ye1D9JfabHg575SAPg4Y2jxgGNb5l3h3HiGKGMfnpnuid/qKBNgHxvMS0XFyakNg
v5CyGwkzaB+jzAtdSS+V3T3fXxrgl5jDj7wQrIVzjRCVJNGJyGTckXS/qc1nwgtaW1FnlD+Evirb
SHAdhOvD287e6gvs/7X+u0FnskWvUvsdPb9XVvee/a4V3Jx1YpbviQFQg9AOzmUQtnNCFGWbwt+9
RKX45KZyLMQBJ6dwTsik5tVegmT4yZzVaX4fECXZ6Qcm3jtU4XOtUcY26XLq922fP+vcXBsL8+Es
OICPmm8dmq4ySBS0nFG7GoxA/Y7NV/EZyugrqdrb9C3/IgeLHiQjdQbj/gb/uMYZwKEjzp70mf8r
TwmG599zO5zz+LUMS4h6D9AOiWiy3Pn9lovZOqZfkNx4BYeep1XZMpJRkCyFAp8pTiAiDnkHU4tO
CBZ5u4Q3+un+foIBgJHRTVIL1M8QYmHBQAL6fJ+Aj3jipFhov6B3g9keWGVZz2ZCGuCiW7fpylsG
3ZeJskNcQJrwVTAck9WVIEPg9i49H/sj5Sj4RyBhtA8JCSTzyEEWIjjovs7Jx53gJ3UF8me/Ni5t
bd97Z5WZklXEHJjgisqYmPyV3rsk8IyyLLMLbuYtftjNkFccNGtheoTqS+f2pgSIF7Xy0dqSTZco
hGUs5wBM/Ii+rTdA/FunAcTgUp9a1AHaLdb8rTuhDquusVdFRTsSqwLfRp5DV0Njtvn7DmIXzYwJ
bVVhQDGSgEUrw5X6wlxJfS3rvCclAx5DeTualrJh1emfhgu5bYULPShTB0xjRmRkF5quydBJFdlB
RQKoGBIb/8rd3U8lXDfJTi/ipsmjmR1SvxtxNhcaYhxRaSsAwXZ9UZ9SKVNADHzUolt3HM2xbTev
ifxtc1seDU0OmSTiew7SnoZq+mWPlbnurYJWm1sROkQOwa/3WMt9mw0HXFpITOuvylf8e8YRz30r
2KgH+67o1gFUqJkseeWy4YN0oIg4PKCONjIfcDH/4yRGCW2QrhQdNFDrmDAiFMIWC9zLZqZVZduQ
nFUnS37FLa1geOYzU9GlM+3vYCwWGCWqgrNPjbnHVY0DARZ0f+VwnaXto+wml85XDo9TrTLhpaKP
II4plVQE7cjsZJsJTtDHUk5sbd5m2LQeH3vVQNs1hy1iGeNXUo8zS5IWRB4mSQD7xh163IClactp
DpPuMcH31uxhbFE1BkoSYmh7HAD1O1jEDP70yRhAporvDmiLXHASXBBgRbmyIbzmI3Xcoyp55cnK
cSApkxLtWzWaGt7vdVpQQZALP3YKQKnjfbkR2GzcVv07UKMx7PDprk1pSgAX4CpYxX4z8mP58nHH
ih4U1HOyPxoQKY+pzvF1DUOWw+l5bLhQ2xgxgT3mU4H4BK+sMcRRmSlQmRu0GxMgC/febmCECq5r
BjsxhhadbLJDIFeu5t5PF8KcExFpo4FsyJTwEW3VzttpAzHk/aG9nvghF/B/xdzv9kFxGnWRZbWd
b1e9U+M16uPiMWBIOPLgLE8+CiWRLTsmXd2npfrRsVZrWXMIsNK1oL6q6Tm4tzEd61hoWRGI0pU/
MEs3sUeunzYXjnN1QUZEMYtwYu9iHDCBOHjqYM9xV6WtHm4oWLoZyuNAJCw7Fyb5aG0gTZ1vuaz5
UuVX6rT+RZ/ZnYOboZAQvnye+Uuk6Vtqtyzh0MiDGeQP1o583LhSuVwObP4WHt8OBdiTxExBNkHY
vW+7O+VhPVLaJSNZ4kf1Z4sQxFL+hZuTP3CpkpxznUZzaki8weZIOgf4iI8iJ3plSfLwB4CR46ip
qQ0yWq9/fkX2umIVYKpQo0IrHXUZajXCgRzEmq55vMEDZVLwQKH0/9OK4Qm1WrV5gZiaAF0ZqfBa
ypLBzsKmUNlHwHJCG0NjjVpMuKX1xS6UVNyvYVrX2rsQmp2MEpodZOCKJrVuEtU1y6NpaAgTdfMZ
5lBd+6wHsiFzShLY739lQsrLQ6q2FkpUU3VnVW9gGOYip8aH0dF+2Pzs82x0wpm8SwK1rqWLFaBu
BX3xHycoOUqhZIO5OFkOg0NqLbgVllb3oxmco6nBUAwiV+9hsaLc+jgl4yCAWN4VluzQRVE6Lft+
e/mZ0UPMX5eoQSim2olgrB0rxxSUxLo2ufhTQUZOnmJMlcf02ivQrZXQcUMVCBh2vOCSX9mV2h8T
yNgWdRH22ZXGk5MBzqBx40PHDS2QzR5ZGM/jDkfvoipFb2HaYdJ8BrlIisYzpVh3i+4lnR2z16dT
F1XJSI8Jv90zvZSEVXdAoCccrX/t7O6HPHC4wUNLEPeVAMMFuTyrpmiJEICAkDSlP8xo8cezfBym
442QVjP1X2Zd+5R9R3QaJCwBftuuQJ8bgQ702JJhdjdOEW5LzkGVi6PL9w1wzOiIGxb/EDN8P/qw
SG7lvHxJM9D0pTn+mVEunTYakqTrcqaKDgSMRqk/c99rXs7GZC/YQr0FmdBitUPeH31x5h9xcTNi
VTWouzdTNBnC1xHHJeV6Ti8PIR67CIPFH5iJO17Z2GaOJId7pgQTmvs6xl4X+eofwmlOX+F2J/OL
mjZ5DuVOoVMI4L3outuKFb0mQP3vUvAFEh3PN9WXxb2MIe+pRM1Z30D6YX91AhdGPf6wrmvHbP0d
fcy3HG2YTF65N6AiqAhSVhCkZXpOJ7fo3481ryZbTncNXO0ZMyjkOAKDxBGfMt4ZQgexmLgMOE5/
YW6V//cwWfH2HnKLWgOe2/mSa7/tIDQ7NV3fkh9ZpXs7Fwua8j48ePR1mZFunJW2Qd3onHwku8/l
vJ47rNt5uv8Z2k4S76JVhjB0nD9K+X7t90gYcAqOXyqwkXPdtUtwma7ux8I2NwAeELazAOn2oZua
1DRTtn81umOmroXJoDt6bOOOsvsbHaC2z02YhBmy72r2ssFcIC5+jN52FAFo7WtZhCVyQlImv/JM
RIuCW11ZggJom9rOQWSEJKbHCcAJK8QoMuuztN9Zsvdx2ezWMppo8d4MDymMEZe7eYZdwySR99MJ
xbfejbcHj+PHx9Pp5NGluTbo3ORk3Jl07AUvg+UeZdE4Su0Dv6J6Dird0cdCefb+E2MEhaNAr3VJ
8xQXyVdc32R1a3bmU4qrErUYCS1nlOlSOnVj2gVprvhvyyy1+73QbBTXzoNnjsykiI39IYzNfhJm
+UrULuRLNcdFqEhPym2dRmsoRd+wjWNmAq32orDagefTJLZJgohZQjEiv4DPFIklfJG63hMfI9b+
MtYjQ7+MnZuzHcgrbTqYqxpLyfitAmGzDkFBlw6KRoP9a3eloWGwcMKQhGD1Zth9NNrYLnUVQ28E
29PSseV0XrhBxo36eFzECB9ZrlTMeqOPtlf8Dui4rIW6L9xIHe0cm0uEZon6LdGqyZZYvmJXnr6o
IptyXiPndX4Exm2pvDnsvwPkGbuXui0Y+FQDOnGUvGeG7QbIEbyO04cuC7BPQ8jjUhoZCzq9aJKI
mnrapeLJSWtubOKgzmnjuH1LOnug/qLBcIeb4qCFQtKN+0v3Iulj7NX5xOgc//rsSPLNXQCmR15v
8OFJZys2I1SQPm2BNB89AcbBao3ABecr9uYekQZrX0Iu5Cfbf4Ss1FK7pC7jE0vWlzdpu7dZmH0M
zg68bf1g2nfV6fH32PRtl0alUcQjJDU5kn9e3lnlq9eIvXBdcOPLL4bJS1T0MBMQoEVFC19iMxrv
cyF0QZZTzf5GdD8Bf2r5sRmeQtSo4+iwnkNcAzthancpEHCW7x71TvN/BtZm5GYnf0GF2bdGNkPg
ByjLxy5dMehgjhZQuTm4QCSQZfRgbv3RVr1lB0GfxkJRyYbGY0NniHFBLYj0oqz6EPKT43RYwt9P
r3i4O68s783SizGaPEYY5fzF4yF2Slu25Fp8a1odYgpV6o115LZKYFkAuMCqB69W0Wd2Dn0HIK3b
29oJ1trHpus+8oolIXJAVJx7Jih8TkmQUg01i3YOxxbyzcVn/IxSuy1KhpHSOAcxmNbI7ZgxKuig
05CPcMFic7k3qqV7qWHLdTQVCcSj3Oj2qBpy8RluqLvzMLbnWDrAwVkGYkbb2j0zxG+YQay3UsZD
+iMq57NTF6zoCiPYljUpjCV7kXRSCv6D5RsPPI+6P/QW7eQRw8/jclyZHHYPIj1ZUc9mK9zuZmIS
XWvQ+Er4tiJd27WhDuhV7qpkVYcbIHC4N3cSm5As9W18r+C/n0pWmEIHe/a9SpvcO0PqHhHTYXOB
Qc9nayt2ImDFgXdl7G2eZ80fI33i44ok+abGlUrSv9xR3yHvqQjS9FC7fv3cRXiueiO8EHF8+Bx8
6WLs88i6ZCy5NKEn4g6VAAQ6ja9O1YaqgmwdazJKU0KbftAFDq26nI5kGBa3frLa8CF0Hlh3a5Fk
PhZWv2o78ryGWVtEhgAzRDRjc/OmRf5Cp86HAZYWacARPdfWKLWYzQyHR7Z18hITmLZLteDcKia9
4750NRqY7xQe++e/FYc/VEbXDVOKXv1mxawcGJ7Svj8n4xgfzIRCzHWjJl1rhi4GFTKqTLg0bQUw
d81Yn3ZBDNt5fNPI3UgkvYRlU/fg0Ql7MOPPdhNu1ZRzumsuTheau5XjL7cuEd9G7MbhlfhwcD9T
+0LsiULpDC8+uYZQ0QLW7ocDo8piw3Ss2RXXoC1WChPnzH2IaZRFhcIj/n2koffNaju/AvmhGqof
NrnmXyvEBoffzw0WGQ4RrsSNHiSWmQx1YxQD0E30ZRvMZhYGpDZtM+mS5jR8FF3kvVdqgEA4deOl
fW3TroRpbQWUaHn/5UZ1fQAYYPWr17j2AiO0ase92QSzLxm+bSxgzNp4vPBvdI4Uxh7kfolRcchu
dgvcvDfBl1O/DBHwCAT2j3x9Xm+Xvy8xSrrvVR1TqRwp2azYDGA+XzSpMPRy2reMl5Pa9QFSO3FE
HcMQGD8O9Jmupzi/SgfDVpWAW+6D1PgLOE7X7VhGqOgL0/hQ7SqDLeJMZTjEFvMat7MqOrwlVwRw
ixwmlBCIUGJNQZO9YGIB4a1Kyq6XsCIdP4SJRTEciHwpmK/boIpsg3vcWQTccZBzn7+RquQuiMge
7bHgH6Aj2GhsJd9HhsJofzJLgWIb4GKAEya5WRKY5vm8zbAjhdMEILYzkGfNaMjLCrqXivsqfQ46
U7odCqJzF6ionGzoGrakxpwaxYjZocb2wZN95S7sZzYzKhtfssoqDcXulw2YFXADHUCZ9G9i8pOW
P2xG5vm7N6R12zC99PZcY0hTRhcIOx2IUKFMjFijl+pfv97HUOF4l5nXmvJIIK+VZCDYJ8PRm4LA
dJDeXx2woGIWcGGuRIGHuY9uU7JI2l2RivdyCkDSF4nVkVyAnGspfKG/kFYt2L7T7Y1hbmdBFbom
3mQReEQYqHGh34iPMvcW1d6BZYkiWdIHg2N8iwf35PplC7h8bybRU94WsUrFM8hEqqCsgx3y2S5j
LXmVeGfVkxVJzhrXGKZgIDfKihnVXYKvdQ+9ZgbhdDwnGtXAIQdp4EpmrumyfDc2GNp5TaWAMAjS
dvYDLqxZ7+znuLdfu1A56I0F8+/1zCsfYLiiNhgdilMVW8kYQYbsOX2vxAvQ3l/Q245xVQGRP2HM
ycxxd5Ki9zr5TkghKD64n/4bZNSSFZys5kl3yiF+nq3iZ5fKqA0FK5aKvpzt72qKr2BcGZ4cdV25
QyDs06p59q37ELlFzQ3lrz2rmeq30Z93auqOR3o6go6Wr/QgHyvMy25b0hF9ZCid7/1h09pbt7Uk
fbt4y2bm7+AwMNMbD0unQzj1PpRwX4ClphQCeSfx/xvmzpzDCEIf/jIBSKAEAQzP0ijWlsigyvuR
tfvO2P9y4djyvNgcBo7VZvXq08L+Ng0IP/UBzEXfN72VN6DQj+YbRG66KVfdyB5gYQVK3GNaRZTt
PBgxLpwlLBzdIS2KhBLFg1lzYnvStADQegMzYqIcZtHviF9MyMv59LlX9XbBdQOfHGdZkkl7hFMS
DvoFaH8+fPKchiok9dIjSuM9Oz4pL67KeMxD9pK4do852fEC0ENzg1kZi8eD8yhTnKBjPRqVuD+f
iRVsoET9Qo1SODcRMgdfsY87BWXrKKGQWCElAuWR3jupp+g8CtJg7y6Pso/M5cB2Uf3MFaZTs0Yl
/BqPq93gI0vuzxmxPIwWC/bFqAazAN3Ixwm5O87jeQ5tddzdlNK+q6rLyidU8lHAAiuKsuHExlaX
XkdeIbI2qku4oJeZaHVcJelQWXWRsfKfs7M9oC/AUhnSZLYWNU+1fD01BV62mQcID306Cg2KIWr9
+djRxIzDCz+ji8C5gSpNg0YqW5vpgNgH2PKB+MkNopsit6uayIxcht7JKn4+RdwapJIetD6m2qr+
2y1QjCzOrJbgn+55PEcYU253RaN7dcgnbwrgde56uSQ93GxNWyeIug5fEnHItYiwJEVK7MuQyeOY
/Ssg0eDFYWGPtDxTLLcY+88HBWFmHNAdBUlH7/a8eQoQjlmIzMnabeQOGiM3H5gALsvZFEzLLe6b
RPgMkEtXZJDX6Pshwx3Xv77vEGXE1NudQ7Sq/neylGcH+MXoA+GkTHQyzKuYQ6tBRcghNcoKOBfj
moljDjFMkMI8Zg/p9S/sIUKDtwQxIBAV2egYWJnN/9sFEFBqTwSl29q7J0TgU50mclop5OQ2Mw6/
mOf2MdabkO9FyM3iOdRcV5TpQguU6XK1luMGoGix3yv1Hky2XUNcyHrBGeJM5tO8kQ3l6j6I8q/I
4jxYHm27GreNkqhkld9g14wlDxzkKOdmwT5fZ4tgQga5IZ5X3Xs4V9Bwz2oUXbv4ulrxwhWe8T0e
Qj+m9K7yRXraqHacbLYMZVmrDWLmFdNcmCZmT6u9bBAnwXx9072dawa6PChciGZJUJPh8Xyg8rwc
6vVTtTXJ+2UF4lDtrl5ZMz7uoFyhTkG8W3MilW2+tIdzGbeHm94g/mxJOO5yzxz5TnPO6VtjB7Q9
ojpUVNBnwXg+nXOCXvigDpssNztSV0t7esCUdDYMWZ+gWACok+QPIqJwOGqjnfB774NEmR0sX6y4
T2988M/48q/WEARYDXKEQTecd1Wim9q7mMTqL/mrGjLoI8aO+0SfWX7rwTwWDSUdYU/07Nm8B7jm
SD5y/I5OrwpS8cK9bTR8q36KlawDYZiwEo2atFsaLYtdaDULGMjnU3ASBiEqKbjN8wwhzhW82UtI
CiF0VWlehtPCkQyla53aNkUhz2pxPjVZVVRkW/fgUPjGsU4KutpDWmWHE5tjBPgMZZgNp570YQN4
3ETBRMTTHqRVkSgjniqVyIE7fdOwru9WKBUNxZTk2+opqFsuV9o9mEpK838doFPZYC4/ZBoMTdEu
AzMXY073bTPQ2BesmyXdEky1zpvA5A2RqyHlVTmlB3+AvZExMpRgOfoTqGJQnwjCkMdwWtN2wB1j
Rx8S8q5SsxDRdNxJzg6jdOe7Y27tUenvqD8rwQqYY7j6dyX1OvdkQ+xr/rMsZA4vShVx3cLLZRND
iFskE6HlVZAkI4on/m9kmKo7hkeR6SSe4dEM5SvET8iQ7iR8ai45sC0CD3g558dH0NmHgQzhJ246
P3+lADZN25JucC5TeE7xSnoV+WzK6z6Hj7B/ZoK8pByToYVtxtXjykq269Y0wppFITtBw5+C3mMe
xRQyUa5brXtY0ufZo2KMQ18Pajjf/3w5EYYuRX9bnyTWMo3pwm0ZUDfeNoIpZMxpo+C9vuvofUlk
J7WhP4pprJnj2mKPDO6FUZUJk1xHhW+X7rU1fv2dVhZSRRAyvSa1zIQcGo/EHv+cdG98SbdlqJJe
BGiLYjwFN6X7q9lBSjJpDU0/GHlXXr8D3QzLQS52dR9cl380i3Y7oWETH9jGIBgdB8GLkCYWIYaH
e1nNjV/tnNpaF7h1S8yzRq+HJ/5ScOwDxxR/AEYy+HKk4/NjvVjUrmyJkzreZfpBJPWiL0shIGZv
mXcpTT34DGm5NaOXpOQhOEmVDuomQ5dINhHAqmA1EFrlShUA81ED46a8aZXCYShBfNyQ3wB40f4Z
r8cnTK9KuqGSI92/4WQSQ2ROBS/BgBhOESGOyvF8P6l5Kc5dvcqYRKLuz7S3vFYzcZfBzGlSLpb1
FBBFsK6EQ7tsayFJonvLYs7RSWyb//TuCfWQNHnZ5NnPoHFWb4WUozATuLhRHnsjBy+vEt8im4Vs
tbROeOQdSDc5IKGjwrVESU2zTpt7/uEOhuI0MNBFDSwdtwmkSFT+e567WLKUTPPf3y6gcYkfMejP
ZRSWjg0qX6fVdnQikgbMTRYyjItJQUIKpGsdBswO6jDDmeFCnRIjB27/DsdwGPja9k4iT7itbTqw
vRjO7jsDLwtrfpZKRF6RS1BphR06gbyeJxAGaNMvJqHMQqTfLC1tJBOq/CUdeFEg8pQkx17NULk2
sOdS/XJz+GPhWXKEapVdfiylKqflqzYelrLB7Kg7RBJfxh2YXY2jFDHj3f7hrmbzz8xmSEMYvxob
4EN+8bDjnoRUI8tBecAkeVmxqNDkU5O1B8IA2dbEz/YMPzvbIollEbw01bi7tHram25kR6N5ZVuF
TElz4Ix9uyhUBpyl/PTl59+dfAmAOKHEoDd5mgdjOLJqLiCoLoQ1UjWozBcChwJXAvzv3C6A6RkB
Rx8e+GaXf3zc8IAztvFA13sx+unLOyp2Uid5b30SbtB88IRcjopWubfheuzGE3r/gYJLkZ2EyiMu
nH8ZheySV49XyF2L2w1Pw93ZUynKPlwjEzIa1+agTh5UeVLWR7nevjJXXhGKyrDGgumdtP9W7fVV
AY8usB/XXgG0TxfmuPKvAGV+NDag0doPVMEZ/uWeBlsSoTEeTINo6bXmA8HeGPDa7IyX8ia/xZQg
m/4KZ93/qmsni7BkmRDb3MZ/CLlb4byf1O5hyE/euNwWrbRsbSezvb7qVigcexrmr5hsi4PyhlIf
+jYj7caA0S/ZRHE2pvL14kGGPkghX7O54PZL7CJy88D79vg+XCXXUxIKeqwS+8EUQfUqSnd0nhSg
kb5PM5xWRk1aqXXWYfkSnpfhBy2GG9jNmUNhnmz564ciNuEvLT/L8whs7pXNYKbd1WHF0zobJAnp
200uPnAwGokoyeFfrfuIxIbfjZoQ2K1Cek23p3DO6n5Q6IfwBZ0AhPGdZd4o/YwfBv/Hbfgn9lFB
UmDrSj6iiiIzqB88Gzf0WCwffr9RnHj2q3wJhL/wbFLDqWT8Xtec6KM53Z1o5Tb2HCPCHdd7xCL6
FHaAqjKTRPN3BzXSdbA/4mHEV5vEmvlgIbDwrUzBtHRijypmEsumvjtyUGPtcqr+VVhqLiaJe+yq
5syNfAc5GW650c5FSSF+B6yfRKnKwlYdx7EJwm5Xiuhh8CmlxMaMA7jLRrkwzGIyOlQSP2YvJ17v
mvaiKWNy1FKqbOaBmFnKVam3u7uyLtU9iab872gC8N3ek+ILI0uOkn9nKX+rmiI86Y43LmFct/TL
tjQqgqlfSKg3aw4qkHq4GxJiI6UELHgpSmL0+Tvx06PkMLU8yDbE81hUn5vKhfxXhbqXTdei3m8g
66on2EYmw4cZjepKPfM7WWK5IacExHWshEZewRJL5BdvCvLtiVcHSIQVcsVXnxez+AIqCR9ai0/b
e4hNhY8/s2+vUE7lmrjahdBkPUL8fQnGmUKJc4GHKrYLJwzYoTu0K21LbBGllZ9cGVGhQ7az2TA2
77kea9M4vWeMearRh3LYEQ8Iugqs8GzaLBVI9E+iLo0H+/EkFnBQkofXvtthOOBtw1KQzDBPNMku
RYSppZr1JXkr3nMdGl0HnaOh3gzE4Z7h5EbyJEh/QupCQKh3VsIWuiVLB+cpGFypEKfU+UO4MP3e
qjQT4p1jrm1XQBvhhJrjrET9VrprTsX/GjSpjBFE5q4Qajq6rCKU72I9aE8jKdgBd/9QQ4+u8xWG
L7MvhN+Aec7l/4J/BoeKENMOPlv4QMjrKXNp5PVPqfD2pEgcDeWTJSKZU7Rriy7m/XvPm8m8JyCm
B+R+nqVdDV0vt5xkSVxxZ8AZpSSu+9rPzu6VeLh1/nk8hOx0JzylNZBPxroS3MQI7O2PP1LGYoye
g+E3n/fwFMVpZi3bI4VyE34GQwoft4rfRX9liTiF6Wnzt6GBTAxqcv9IHICCyQmdcvB2Q0M3nM8F
Sn9KmZyfdRVmjXQhPL3HW8NaTdz4aKrP3CY2yzhwX5ZIIUxBNEnS/unNnYhbbJuREvoX1QWlYcms
lZp7d3356IM5rD9pg4n6F5uHZTzHcGTMZRlGfQ9Zhchm3sjbDBXGAjxCXIkIuWQhnBbUJJZ5tick
aB7pUEB6fkqhAHhr79YmAQ9+ov9gu9cGXY22Ov0nj47xrv+7KnhPQpGoyzmmkqYDNZQP+gTk22C1
fZun3uf//BhVyFJvg9Y07Xajj+lRclOi8WIOXi/B0RHValP7Jp2UiiNV3tM/tMGDEDJVHzdpxwmW
duUjVNEsPgaFLFKkYpzRdXABRd3HGh6gwV/I6sDJsuCUw+pSnkprtHEnMO9e+f1JgWw4dqX+NrPf
EPHSIDjd1GkmCqGNa2QjD4JZc89nGxLklhAQP6Vnf9T3qPKZo9qiSVlVak34xUfKxeIyt976uFaj
dD5CmLgPMYinJYGMQCdnQCcPYVpU5vqbNb8Vlr3raEQEltsz+LE/+EjWKqFg44Sbbr9K17bTtJtA
Ju2e/ha3g5vMVrxhOq69txPv5JDIGT7im7Ae3wFbZGtJaRehh01eIPSqJeviklnyr+hyxhN10w92
+7qYAuKMgvwZd8I1UCCtN6W0oiednGoqPfc+jtN6ctvB9WnJn2Ul54JrJ13xJf3ihM3dgYYk0k39
Z+du3+K2V42JKXtQh3hzsdC5dIZVgCQyDz1xsdxqvR/Pgz0ejsePkM0+qGZjXoje6QTgGs+kv3WI
84cBYX7WVZFWPejPKJMI3AH8e2rdECsGfIPis2vdJ/T3Qx4CbzHE6QZw4H3nnjeHkBihnFLrk8h6
23hKnYrS74wij5dVzNKECc/rHv8YCzT0ZZ0nF7ZpBzYVJZXa2VXrZAQ7ztgB7nZU3yEXfTeNeM0V
jOlAXQe2+jZtez48g2B8MBnPttLGf0XoI5DzeZO8SafjttqnRO/BMT13ShbyEmAZbtOc5pfUpvr+
94lY0yIbT1E1lPd3ytwuDlKSX3x+qbq0Zol2LYE+QJLaTiE06YowLH672xsd6zUc22bIfdbhMpQ/
mYzwFlOgWYMr1REu98aaZVBRBGAkbdbyVUKb/5M/05L1fUfT/zT1IPm7roG8LUOY3XHibgkr3N7I
kvC7EbOGdFhU3KWZ6eUZboVyAWskJ6sKXB7vFypS5yhBmKNb3KYdBtcI9j5aBOpqAW9A/mcWO9Fq
2MhXCOosrSAbCQbv2vyQPG+XCOmEUX2fhup+TQ/0Jf1Yk0yRP0HKSeazracgSQoezQTNytA1HsDy
HKh8Ey0Swu2aoVesHDfal497kbkrN8Vh+oSrSxktDJZ6p2d+dBvMGKr4vUTscawESGUukqqmNugu
h/fUMJvspDPMXIujt1UItmc3fulYzvsBD+KQjoxIqy+DD9wEtjc4xe3LJixc0U5khsdo09wGJj4o
169LruR5QoEb+6FkzU8+8hujwOxefuzAHlhXU3uc6/QYAOUjwy/ZBv7Qy+BMxpVCWB8mJ3lNU9rk
u7Oy4LBnur9bO35Md/AF7QA1FRt3EFaxmHdI4xVbrmq2y9Uff39Tplduf/uZPPaSdMt5/rJ/F2bK
ebG/6WEEYy/dxojEiJvEdbd4HoKvB2H2uGri+/ruhYjiBdCv/9YfFta6uU7OffNLEFRzz6C2Dcrp
sq6BzB8Bi6ZgVCuoGNgEVzq9F1xaLsM0cVBGu5nB593dXqBdjTCJpHMyy6MwF3SAwPlAVQ230dfL
vMOed3o83xWIMftb4dtXxWzD97pUHxdCno9Prt67XEPyMNxJImwFZzg/iwFiL5jtLwsIfo00Klk9
um0yPBM03Y0UXryOtgND1Igmkr+vKeSDhpMpK/Yh59RN6BTdkLN6DoJ4gIFCrxVnxCe3YG0yFErs
W+5WwKavRD9rI8kxhIbLwFmxieacD5aoDhn2+N1laGRrrHDPerDAF5q0Z+KXhmTId9D9zTImCpoX
snclZjye0vSeNcheNMi345xF8yCpR4P/czGpDZka2q2MiQqu1RzOvIFVf7hox+rBEwfU9vw8f8Nm
M757l47CohMdoktxRd+qAI2p8X/BtOXvLzbf9+EkgWVRM0eij1SlObJ/H6SOjL+lkBSPl62qJ3Xa
jV2p0t8xQBztMDf4u8wHFaN7TBt0WGp/HTcxacArXjITwuVU3Oqv3tb/0L0vId0O22UbXcRzDuTk
j2zedGj6sYS/KwyDXlhWsZ8trYjFF2YOq3b4xBFPSCWdyxV5n2A8HMQFk0gDmUA3myGQNTGVjcS4
j0VOpO42hoCZ0CEHqW2qvi4UAtZXR4FEebhjch+r3N3y4DVe9FxNb18vNxpqh7t9NbqFnU5r1Dao
HR1ZY0D7ZdKftrnhAhGL6abNYoK7JrkHCUjD9DTLc1nQ0kWCDBlf6UH18EOcSTpobDyS/K9oK91Q
VWFb9/FnZl80B6QEAgfmJjcu1A12WptlJ3oF511oT1gDli9AGHe6ckyvkYZcGpz6dlHi2SKSMJHg
jNMbGpoQ7IfedM7JiWGg1w2F3Ta/YkzKLYQl3WtT2NGexI6WIJwgxelWQhCUdRrUqMJyZDoW/jbb
0UfbwjVYe7pYtrbukRaXWlxtT2Um1E2FFkf1/kxxs0ndP6DgUOEoqCAgTCPTDN4tfHBlCfM61Euo
SLsEVasuH5v6oLjTwFH4CpdFq71MKzsHiPXYjOCnUjkHOlA8IScR+pCoFQyMflT/VYwqIcD3MiiU
2O97meEQuagCrYoOf43Dnjz3/kVB9jZ0U0d3eYzwIWAS6sE7g0ZHLpniS6PfGhRkyAVmPXJDbhA+
/UlNNEIrdFlx3NoUCrYLEKdBwJNRcG1JjxTO7Gmc43se30deagQ04ggWLsUdVRQU2OdlkZ+Z1XtL
/093RFdY8OmAaJQ7zSv2kQV8UBq7GYaFhNsl546jXHMXbqZtrhNzZcHZOkcpR7ZZ0MTkT9ohvwV+
lBN8ET+NTjp3emwweIgRDcEf5lKgMpTuqJRZ5Hxh7N00futvb+WGLODE/8PyIRh3t0UD8drOnv4n
Ayoy2/qiFh+jWAnUF/TH/x3y0wO1ymUTLA4lNS7tENrjvBCQ2vEMQsNvGAGYXyrADNnPTITHHoaH
idRBK6Gexdbqoe1X72EzzUBio6Zghcl8aTGD8x+rhsoAvgI8/MEffBVX+K0CPGy4S9tsUJG49Xx/
ZaiKx8M5A8miq9ABmyCE6n1rwNO5gW4uoMe1hyLtLaz9GSF9fV3JZaKG3O0lBDYid/iDuU/1P11K
wHFO3c/a3QrEUH85vx/02AlkXzbKLxQ2UFH9QYuTo2V2Qdy0lb7GNCJDus0r30/TDFMcJjs5IKll
LbcmdtDSVPl4D9lIAx7sqyN9cqTu/megWC1hTvWLWDBZSaGUEjVf3dnZo+wwswpx0/O8MzZGgDZj
0N28NKwVAYJp5D2EIRC9mtZvx0YXivIMlUkSvo/DCBFjByMiYRzFGRi6K75TnQGsehOcujHaJ6bD
OulDfYiwFnnbckkd7StbPM3RgP9LhhwyyRD2N9x2SEMjGQEhSWuYiNXTiaG+hZxHRZyKQKgHgvet
4vNv+paXPixAoF3jtBbF7HTI9odTgCGrgIqAM2BFe/+8hW0ypaBd4ZD4uGwzLSJ7+eKtgNnpPoc0
GyNGuhGOTXIrCAj2PxAl9MSAB9etwcbOAherZC6iDUhPuhFHW89wS7p3ujMI5fgE7MovQYqCQCzI
sSw9NvtMjRya5NdCC0FtKr0ICCgFeDbctQQtUmL1xqBHZvrmVs0Sf/loYgJG2AV8hUAQJTmTS6YY
8xudNRg2sgpSXwgnVQ1F76hexcdsncMaq8rl8jM8tK/A9Vs8IwQhe1USv5L7y54I0nd71MBXn31b
4CbwNQh5AGvq66XkOX1FbY3YYKmDE4b+yOGGMPDtfc7EbsC5qqa2hXPWaalbBj3s7XoOshHvDdL6
WO/kjcuqZGvcp4UWNkyCol0cxq91MqEu16UgwDaTGsfqBrMp2ard3Y43gw7eqqSk0NK59qrSG4dE
MHRAW/uJtFUeYMwuOt9l89Pl2WncfzBnDapdqt8lHATqbT9Wf90qasqgTgisxDOZ7wUWovc1YLsO
pi5/KZI3zOj0NtJ1LdxNfSdZXrld2YnsmXIs2wm0DJGK4/BwpuWhMhrEH2aUtaUezow+9MzMDlgc
RKhg6lp2BqI4eppdw694y4z5RyVbzEkBEdrnYtFj91Sq7t8XSVgalHe7/8CfpeTVBrTW0/m4CcOu
naOowOrUazmqDfkjA3MEWqC0VcBfteVvIv/P065RML2kbLX07/CnnPtAyVfwJ+t7U9+0pgIQlvRd
4wuL3+1hRc2Miez9Y/5L/lw3uUBMklZg99SRz1OnfRPy92itzevmeVGTDzu2gfGOyfYmC38ElKq5
F9v6RjerXvXMDTCypu36HvIo1Hw6qclgUi8Vo+752826PGor+PtoYqkfPvc3bORB0ioNKuPGy4tA
slAWYbrG/dmBKctCAM+5e9ESctmn/3HwO38jZ4deUp7zMwT9GcpJsOLHTaya+yf+6pGLFLEJqn+j
WlTzoumUu2C8J6nIHpiT5vn9zyCX9a3AeoGNXjcIriw+uwjzZETIXsbc1XL37La4/kVePdF6P7t2
7fSgXO22+fO9jRUvcbNTZulw/vWSJC+9iN1Tz+LZTYR0lseSwLgOqx+Mb2r5M6DeeK6xSvcEavpa
MMDa9kKhPf7eeTfHop3v6L6ACYHGdcb/te99RrB4IOzvwsWQjwrohlhZy2jTNzJZBwBS+zo/M7t9
YfNRPkY+NpIGddDafOO/EbZeCS3z4DJ7OsxlB1UGiKt83uECK/q3MXXn3KCTUOHF2Y4jGqfHVAkj
QlW2+i/RfTBTdkmxyuDAwctfGM6hnn22EyFeSm2QbENnp2p3Ajetza2P69rzIsrCc1NUB/jrnciO
QixirufB9YCgYvGT9p65mlXJnT10OBXR2aFjzjA4q0xnE+IC6SfkQRnfMvPvVqIHVmMjq1MXNO+0
qVGmddanuYGxUGs91U4izIUxqrMzZ6JXNyWYqdgOEem2eD0yaq3eFv6O5Nw1ATnCXnGV2MoZqipR
7orosHQY1V37+T+qJuf4So5sYcugfB6WoIf3cu107B4jK+S4DGtpkGqqLW5LVGufGWl3MdrlbTK8
YM0mVpxl1v1pG97KdLI/dHzfhl2Z4I3SPJse5sRfo1VARJX6FaQAeLNVFOWHo/fz8nqyRi1Gu+eZ
d+7I3JpHx/IsiT4XqT15Fi07egrAeTCbAhflhiD9awth0dK4183XGkh4lwXufiEyXEkHN6FDJP1Y
itTdQn4eVwGzzSVSUb/XZ49nE3jsYw3bHs9oSyGX7DHvDd0Lxzovv5XNjL31gwBMg9sDapZZpoFS
UUM1R7g7zhn8xlia/5djVb4DvaNp7VJJt2f3TB4Ryrzg10L/anyflGVuoLxv1RJOP/ZZQNKxj/ke
7T1DvLMDCJ+vNLFvU2GPlvFf3q8Lecq9MEzt68g15Lj7CEmbHeYX5YpEyyHXZm5fwL3K73qzRGSx
Yl5ju97RVrhUcCxsjdd2qNnqJeB6aBP8RNZSY8tlBXHiFOYwg0uTULsMW1oYsZISItgpGa26+dwO
/mxvZzZMH94u6lBvlsgnY4HfneLiZ1R3gXAeAQ5/5Vi/t3UkyMLTYeagfIDTk7UExiSOfHzCqOVL
niHHscOsLiDGMsT96qG0fyB6NuB583eid5x2KqS9UcCFsdwWbJaP2N8l/eWeMsKvXdoEFe/6MQJy
jlrMVWRM2v9d85rAzRGLs4YsYPBjvtFhyDFosgsQGa58yppbfkyuUrQQ78nLpGyuBm2YmK/MNPwS
VDLAdB/saR7UCqq5nLJ59+DC4HchNdFjJ+BaWBHF/BwzAVnrFMTrd5Q8xnr4s0nmzI0j8nunKOQF
UhRYxJKxXIst8Bq49RDeaRMN+WtSu+pwGEHa9C7jeTkttaRGnkQNxOHkVvomR51dv0Va5MmgfDCs
3cpdg7/1TehGN45kBCAhKNWnfJEpx3iO6YpAfP9laECdS124CRyPl/x1uDMXoN+5ea0KOYJe626V
ZWIPlpO6f45/9BMpkqFlb53Q0k5i0QoGTDaSEmb/1GSrO/RxKLtPY7urLBcDp7eUGJccwagYE+Tv
iWr1xRp85glJtKwJ6htuPGYe1UmsoJdQLa7mMLXv/JAMHFGKoY1peZaG3wO9CBMTd18sAimpQJca
jZ8XWU4/TzpmZqWnXttWkk58UASaLZj5lCJmCPeY0Se/h78Q2zHdZQId6ZO1AZOW5fkg9ZHYCGXn
NPMhcqSmV++jxEf7WN2q3Pg6cbojFzKgFhAC5ag98+4QZTzL2nKrJb/AybdEik4ef+DIz42NGHBZ
I40p8XFrokIK7M8CPBKYKcOadsKNQuDd2T46e/rTO1x0gIC/9l+nbM15rrpPCVBNC8G9MGCQe1zs
WzFH8u4z28zN8yDdq09vyYra9+TYUk46D5zH3jiCXRttpnZHEMzp4+HhwC/nD4lw7rTpPvtdLKIH
zHcKBqllQdBy/oj4DIazNMn60uNT4RHePj88a9IMDi6Ne/SQB71dJxZPTMcgh8R90BFazF/YsoSH
NFSvAjkGeulFAscfJWtQHEHdf/b7y/qVoUBt2iX/DS2PtBw9WqBoTXbij2KBWTxB9cPZwz8gNbr0
G0lilGucX5qak3bMbviC6vt3zPtaAT9Oh65GcQtJd+nSQdUm5mtXAnCa37SmiWiFAI6HdlUFeJNa
4ynfotQ41bhaltRy9Y7pr/dIolGN9inuN1xMsGiWt4nRZAzmO7n3ks04tVmCzeC/B7gf0qgSo2jh
0nvUADQp7VPLmjBs4nJPmdE8IW6qpjrZlWAKQQS9ddg1x1cv+S/HcyyrypJCJ1t7sr4uK/56XlGL
KbNrYoDUPs7bijQDGisanzfUKIJljEcm++4N1f3alcLtxWFqaKo/AYHpN1eDOxs44u8kfzoZCdJ+
7opqRT1ka20IGKwdRuaskSImQ7Xeolj6yqlsRaKFOdLcaeHQMO8m4hrpb4Zm/PfWaSgvC3qzgPeW
nqbEFeYQvG95yBzJEicAEJDmpL/7kaRhq9af6hCzwNtWKmLG9ytZ67k/VnY3GTIZqp7DvjDe9DeI
s4fU6ObDh+jgFz3PpgEUXUZHLOU65blQK6MTaEcbQZ7Zy4Kybp3doyWMPZC8lqerjLuS28BH4cUn
/stnGujrVKxgRlDiMSz6okgWulXD6XYfYkC7bAR5CvDqZVX64pbqROxF3OZq2G/2inZEtLoEhOZE
YXyq+2oqLHCkl+E5cEW5WZjJu/xnjnbNQsajrOr9rGk8VuHiGe4hbiRSevFXaNE589mXqtjoVVdB
GBhxGF6iHo3GUbSmxwf2R5dznMuLM7aEe+EH/7ULp37GiczK1+59H7Zd8dJyKziy+GoEPiwtciez
Vj4YcWsYinDzGnIeZACk6FGP+ZY5myhsy16yMtCkdUUx3ab5RcpHF3TB7LAgvOBTZ2MhSUjpT9cx
VueXbHYkx1PnNIuhkyYk4rm0ZYGR0muwaXF9FRMGhROXuJTbZE1DzdKVC/RcCMQ1UdjXHG7OzMt1
xarsnf3T5QUYqBkv7IwiDHFt65iF4pasFQM3MVMkz8cKPG89g30QBwKbE1ZLjHr50/pArj01X36K
di44waDbucjWVyUvASdRz7veXuu02SLoojJDAGRWADuCkYn4DGgV5g9KkDVBzGvPLc2KV0vDQYrz
+wTrKM5V7GJQODo8ZLMOdXlV0bSp6TaSoJu2AQSGU+ffFIc1qk1e67w6j0TbN2uK6LyeuK/mHaBV
ViKNOb2o126rh+K1deacsZu5SXpAq1dA573n3Q+52XCGP+t8hncATOQT0cQJIIqBoSLUEK90ta7x
0SyIxEfagxYWaNG7JF2s4dFZg+iGqmOzvuXvV5+cgzkSRMj5WiufAbJR4c3sivqmRL1EAWc93lTj
bTGdokqGVjT2Tz9XEknTknANpvG0rrV92j2atr0fHDnEyjPKsITJ3KyZRDOe2gv/yna7luOcbX5e
ycW+6go/Jky/da+RJXM7vKIilSA/dlWMXi5FHMNa1My5djA0SzsRiqR+c6Kps75jWhbYmfYFKChh
NJqRVuR+Fbs/n2CvpCDL+FfoK7LCVbH6CQafCZST9w1x/DdCKHhR4rUC1wkO347YSTAJvcaJ57zz
WFEt4fcoZEJeufd9+S0lCpRGjT8wCFjJDQ+ItM6Oofub9e3n/0oKP9YdSMMoWM9yTZurg8fbIaBy
K0UMC6V674Jj+l9b93ixdqgmNlLAm/IUT2fYGzc5/1Kk4L08NVUhiojLnlHCJhZyY5uInbYZPZzD
blL+zoB6Ma7qx7IoZZPctuxZEd1o+E3WeZ1Mo+Cgj/djfUiQI6sBx4sYRl2kGnxabsiFt1WGeB37
ZMOdnvVrilDTJnWKKJBUgZrqpUN8EViJsfqVCfGwB14ogzr4VLg/IOxbNyssEV/BKGk2wYD6DKbG
94YJNmupc7RIXpU5A9ndZYsI1ycUVM/ZSOj2FucCN4K3gSMD+pbLs3gWcOw2LZFZdnGyFfS1Rt1/
H11DFyblShwbgeq6+UWHBIfPv2nKSq+bgDOqn4pQ2ks6kg2ST1aFG+GfpSyN5Vfp3+z55KEJ4F9A
NiUT/OYUHi3bk24XXhywwQBA4Z0CyMLMLRrFG+440qf5onqmqy8SI16PjCQA28trMVn0V/nPjm1O
RP8FNUMFZLKew8WEUWs7v8oRXtzno5yAxSUS3edu4y84SKkm1REx4Pck4SlU63RdDCeTrW11H6ZF
9NMlTG8yFrGekndYRA3DMbMkc0vx1YmU/7nISAGYeUnVf/cQrCOFBpMm2QqfK6yYCPgbnUmNevQ6
BcTDUfNMHzGIXwipa8jf9jA4nvqA7ebSI+sklvc2e9J5f8bmZsbRXEuHY9DAZWCbf73Qn5L6JQxy
XB7EYm0UnjSAOsJDOj/DKAmSEbDUop7qXRPdMeBy/Mii1vfs/NeLYjFiT5/S4nPtUN+AlG3ZCo/V
I82lJDfdWJJGjkf1hK2kWJIqqi5uaCbhIg9sedHnnOR9+4n5oroj1Fh7WX60mqAR+5nhqTLcfpPY
MXS62WS1i6w4agWlomiMHtADBNqlJgz3yfP3UQ+xX5Cwowu0cBIhJCUQhaqvIWwc+TsqjPLPtI2i
rpYhdHfFUT9BPEPreAx/XXbumQa6AnhGXpvJh6FqZizqLzKNIZoyElWJaNsU2er/zahsG6Qj9Or7
wDIUhJFZNx+NDBVbtb1zGbAg44C9rTymJ/4nwGbE7Jlj9BuYeAj9G2gxo94YGJOkBoeHI1Y+FV+S
tarsLt+T9zbDQXleHi6iLBrX8l1RiJ3s8oKudFzdLsUqgY66HzVrGtAMuBzR9hVL6330dnj2Uy29
pAuOVgSU8YvsrB0qoyviyt1BhdF08nzdEjs9NXkFNiC9JADcXfcGPGG15unRssKRcBNPw0owqgv2
iYCB4RlCOrIoEi+4Mk5egpMwZLEGsH3w+Tt+BKGs7ukyk5PssUcaKsXyVIlYW+L/glXt0kyJkany
E10268uN0lb356eeQ8NOqku2uKvkX3Zl9tRoIuiV8cWIK/Tj3mzTQGNY5c7G7kaLi27287Ieb09P
wWbc4Qp4CTKY9fHTbW3fiHwIdEyQUJ7d+72xlGVXmmGhQy4PchwzEUA/xKRS14lMmlGUShkjSN+8
sbpvViaVKzqFO6Zr+2LvBU8/1xAFJSAbpOUOWfUtC8T8OgzOPJHtbZTkSpckO2oMW1uRfDlvOI6k
QoiVUJrSrKV49GeKZHxIDnFQvTVnTSJtovX1mR0m/IXM4PcMLHWYyray/yK/Tw7oW0Wj/26xlZbd
5KAm9RexC30W/rkThvJ7++bsjv42sZ8dNHxPGA45RQb9SbGVUXs6XWLFEzFxfUNGzOjGae8ReTtS
Oloq+ETvKhyQkc7NXsIkXBITr5mAe5FhZrlbC/s5NY3raj8RFPEraWHobvOuEaq+atY5bykSAU0M
m/H18CBe0umCx6HbXmq/iTMWWIBnnoajMNn0sjc/+WW0uyA3BhF2By7maRSwtGU6UeuHbkRK3sZn
KsuqijlXLvpFK4JVe49k5e5geZYevbXWZnqFwGN9yFu/t746BYNRGi3+77fo4d+vKy+NrxVdwHDj
+zbw8KncXdxqv2PZbt+/eeyKuN4zCxxAOR1KIDSrccY2C7VE2BHCIO4Gimx0OeSeC9jpGVFTM9SM
/eqWManRD2cgdEmpWdq3l0yDQ+zg9Mfrj0K19C4/U76Zf+Rc3HFl2465lJ/DsAMtAvOg7Joa3ORq
gMFf5muLbmDRsfN+63f6UcjtgCoHXaKMSsoZbxBFIjYgEwsl26Op9zotA44kf4AP86q+1Qolk9Z5
KlHPvTzSSetMBHhx0knOfDAQ9OtZ7TnMkhhtv+Szl9EnDZ2bt6m53tjs7zLKg3q8Q5k4BThgApZM
0z6dMDi3HydL5FgNzEf/vPa8zXAWvttzc329dQy7iAFu0ldHXpXu/DjOhDBPgaFgBVgzww9Ziu9p
zMn4KErfO0mXJZOp376W1dtiriboNV9ODl2kxWyqeVHW7l9OQBW7eW1UblT+vdCJtoEeF8En7Ga2
Q1F1pz7rOZpLU0eB2NgmBdxlj2/KrA5vJOLGZLybJYI6IqA1dEho20xiCv+/OM64zNwjriRUTx3k
RqNhEyAnJZ9Vu1GvoNd/i3l8ZewSnxwXH9ITaFillpoU6LVkD6wTaKDkLzTd5MRayiRhaaAZugso
chfx/3kqB8pSyyIdGPxadoGzt9qe6HM88CXj1B4k0Z9kX+AAHz8FZSymfg9AILD3MwtAy7T9W1H3
iDWZdDNbOrSNmZjmkzqHAadCgwLNrB1DpHVnAyrAB5DLNc4iKjzOeMHEG2Uyf67vqK2c9jvqHk6Z
Gj8ZDgbvJAad+LTbXco1kbwQxX69sEhkHqRg4KbuHtPOZgRe0j1MgVIPAfbgqoKhp4+FmMVNM681
yMECgZQp0vm28kL46UKoFsZU50XoIwdJz4ZlLo6LYBiQDp2lRB8/JzegKYGIfm1zA6YFDpMpioFS
+ZTaLMTGPmNX+IEPe7QrCz2GXIur4/oIORP0au9Ed7AeQKX1/sZWjj6OKNjl4y3Ic0w5Mb1HUuwW
kxOjytLWFHZcyHk9eQzcuK9t525vX03hFrqXM9jpMKFvpr7JeHG1+QwxnjW+VUNekg6ylsmMUWZb
sgXD+lOYcuiAW4u37IoLBrkm0H3+t+MvoVdKri9+QsZfrYyROVYrK02/25X928FPX3TmqQWiNAeQ
XVHIDBaAc0ujIJCixohkGZA0FisRswisp7IOc8Bra0C43jDgoW7veK1ps5ggXtaYCMMt6mFzLFpu
U6uGZDMTty62fzJJ9Za4wm41xljaUZ96ItohKj68rvXd+7vnb10KzBE56EWvaY1uJAQJ2JpnvMKj
8sra3LJr+LwbQgrchJf5B44tHG4xcZp8PaYlntYeU0auu4erGsP9tCzcj9DiTFRdCiQT/n5CYj+Q
+1zi1HVatwrpz6tm0M96OeLd75S/1buuP7VgKWSG9GrvWaIQ+CroHy8Gtq8rtylMCUojn2moNnBs
aULa8gOy8kPlmnHsQhrTbovyR9SCWPlLXSAMSdXn/mMxbAT830McofSR+VaSxgH5MzWUBzO8GLqM
Y6LZ6cS6YJmnq4F2Ue03QKh1/3G4jolncD7voI9JZBn7+klg93r4z5BbkAAYIhLitPO/7pYyF6eq
CUfOedIu7NpukLmuBir95gifHa5qb0OxkxG30GiXMIoKzI0rq+T1q2yCI5rNu5okFbkVMdT5mY0Q
tRAKzVNLDaej2pS+KFloKIoKSE/HOI9T8eBvNQKCakdshmMkOZRADRrrbQV7s4cPwdm+lEYY2o5c
tMpYAJrNn0z//DEkBTn1Y4J4f7u+qk3YzZKAc+G2Fu8A/yZoasUPyqkbyHVnFzkhgYEBBO7kQ77x
IEsbf9YwJRYN9JOX9IzNgUfgHZQsdWmWHobdKmGIuhNhMyp/WVE5JWfH+WnUV7bpM+aV8zqrT/Au
0LsQo6iwFfQaNN1vcEMMjchKk3zie6Pji02FjixOyRMYVqXomnAudKLziAB/Tn69itHGlgat94nH
fV0dlURRP3HDmmmvbJi8G/ly2LCKMcA3xDUBxV15Tofg7Lz5h1QX6Zm8Fb+IEYTKkoaTWv7xfbco
SMMRyNmtNZcbufBgC/t9ExUuKQy0vBpvtA4tn8RtW2VhKO5kTzL08l3uSTEQ2jkFNXImNm8298qg
J5Bkpbuf+snXLO9PU7CbqjAbuvP+RsUReHEMEVf+OSEK51g5kge1U0kLeuf8djhDHObN8HHKBnRj
l2Tjq4MhPYG0XOrP44g+utiNtxMfJ4IoOo/WtQehHkyIuuX91SGBsi2dcLJ/gmPB68wk0vo9NoYf
GWB1OCLz0TajdT1JrtsI5KIqKTbccGpO7rI45G6astl4WKwVmSXXUdpCXdjcPb8j8kkUvOMPAnJ8
Mj1VkV5Si28t/K5gbiq6Wufst5XTdiwqv6kB4eQBPomWH3vnXdaJRXtQxdtZZpLMNt8f3qGAQKU1
jhtXGlmN9AP0uOLGJz6kW1KfOAWrn9vKXQjyaK4nDsHgYnBdYuU97+me/WoIbdfC1g0hAa8WWw8l
Ff3ZzfIoQtQBTukUoqcmQQyuM9BeYxmwMcLQd5mWYvVsINqwUADhccCqA04JS2erQBMjfkREfDsK
VVBBOgoStzLMRb8Fgin0Bnue7/n7uyZnLh0iVLqymQSkRCv6K7FKHTjmMwMzaypqGKt/m5iWNxvm
iFHkY2XGo7dSDoPvBqy/VIaRvZ1nmIvg2/4P5nDUXCCLCHPHYkH5mL8LrPVJ7JgoVhvuLuXPOnGB
v56sgbHlv6BdfJUHwyTxKgQM5eLaBdmpAEsBis1e236uWA6QXLl5AoqFoVyX0NzJzQvn/ULqY9ra
IWF8O6G8qUawPAF3w8cARvXR/tlQfVXeMGK9llL6oLZUdazLzGfIzPnA4hO1yipG/rBR/kvlP3bI
uUiEn819fiVnsSs/z388r4z8qUDklG6aWAei8O0HTAToUBorAi0hFDIBo3/jGGv2zo/G5rspgfAD
esjilVzTXrDLHPZjSLIS//pq8PKCEROM5COwZyjjkzzL8iGb/4EYFmyKdifrRSlaaHosvwqZn5iw
QqzGzqXN+0kqhQtlcWHtgP1k+dIFAp98TxFxwiiJqmaoVgYnvPJdre6eEVry25FjS6ZiQxZdwHut
4kGrPpni6RYaFuc5jcCNbZeyzTz1vO3QJj5gQrLS9wH+JZNDINLmaSUabP4reKJVZly8AOxQ4ImR
ZFdTOh9LN+q1R9/WHtiL/A6m3l3Xk3c/TXf1CJnhISYTVlHqm3WrbcDEH66/C60oHRlPy14Zyl9x
QdCy0Bpww82HfRMUb1L2QYFMgoGk05ePKfJkgExAaXj9i3aC2ngdD4XEDdJwJIcbR2csP39KVuy8
52otRnAJrxexO4SmgMI8vfBqZ0WKFGrdCwjb0ZCSYGTNtfg6WvCRcs0FS046z3xGGJp+gM+SiJyX
EXzepcCjiRmA1qoYBtnZYLAWX1Nm15aEPD4qGPkY2y528LSTFuS4O/gr+QptzlJvRbyUhbM4XPyx
9SeOpaqLlEo3cpWacPgiD+jITkuBzXGNqzxAQED1qsVhFbj5xEyBra20rrqNDQtlKJvbNtrPBbZx
VmO0oDZ9wc4Vv08ugxMKve8BWeycYWgLfU6CBJ1kcdgrWsc+QQZ2zVx2UXkVgvQn+nVgiXIGjfA2
f7xn6oui7Z5BK/FPa07AuQqgIg55bSwhBo03YVxhP4moW9WjCBX6/R69UiDq6CNZsELIu5hD832j
KmrZIC48sTsPMdQdUxaxLC4bbdpcsCFj0hiiENgNYUwtY5PaAi+c2bOi9csvDV+NJ+JIXsV1r1X9
vwBzOgXymje+HaPL0sLcNaaezrdtLzTRV8s5xKnAIOApvLAhzYTbTN65uQvq5oumm9TphUw/Vubf
IoNYnx0x2EPFCMdL72ckBbLiLDAfH/mchEln7rLOp36DcUwk5pvhibr+e7R8uOZbAMQjdO665bPS
gJbXzDspEMM2QAwBA2SdBMHv5Kt1Pbu8ILlUW4ymQtsKwTS58kD0icuLGOSjKqYBu0GIPPi1zSsk
QkjzrveQcPDmSle4Ag5uqlt81OKfhrq12BUcET4ZFSxdBwDuZjGoYznqZEKveGhjMU+FJ0T6NiDo
6oGizie5b+aKW2SQXfRDJc90US4J+IofxWQ+UVhJJySjl6nLc5tjN4T+kui8M5ni+ErX15SmRau2
iHebe43l18SAdvdB1/IVFV67AgfGISL1hoYuWQwSUs1rHx2fEvdIgQYsMU5sDVt6O5Vu22C8PUtL
bs9JqIGV+dyMygTjfFFv5cGrtnof6VuaP4UoLyq4BjrpOF4XWLstF0m0zcezyc0RatGx6S2v1PHP
QeCoGoIAgX6hZRTt2AADxgykzviPovE8KIx0tluaN5ARNSP9VDMIKvvL64aG3Gk2VF+fNAWFr+36
sHA+icxCCZXRgCWCiNXtxf5fiTO0O9HocJBt8+2ucRo/0Ch9G0kbviNyMyu2W/lUfMkl3inkGTAW
1OksuDT7ybUYh60IdhC5m38+aRkfTOwcT4W/qWO9UXGzIfdJSS6QdHZgeyZbEc0BAWgmSU0/h6Sk
gVVv2QVWjXsZiSDHfVP8Pf9GrppSGNy7UJ1oAjrgEq0mFcwryLj7VNpnM9rkjJLOZ1UE9YHiOBJK
jyEsS3J5Ww8UFsRvZq33seFEatMtlMCS7M+TR3m+CoN2VmxEygSmOadz6vlJmGO4XP870gmw5re5
PgOkl/MhyZf/AiMtfWZWMA2qnVtboempasxn6XIgNrApu7wMxx7qSQx1HFg5vsUrSS5U1LD52qr6
s597BUbcHiiqbgMx7edi/72CY1j8Udecfjxf5rTXfWe6+BnSDy1AOHMPRhb9x5WqgHA6pfWJUuGI
TVfvAsrrGRa4XYdsJqSRWrqkxL/nyVkBUNSUHsusFS3F+szHS6yjDTg+e1I7yi8Xf4T/5ZEj8T/S
Ru3MN147XqVgPxGibA6UI+bIFAAkzkO8IrAU93eTObJtvNs2GzPvV3pDrnngkk3vEIbPjjln4Fxf
3jQjmGi1AgqErmd27xM2bLlWkGaAfkckY6JO+g6Dz+41Ecb5d0A2E88XnEEtqAp8tdyRr2VZNDYV
Z/+nTtSM7S/frO4c8C2btG2Ks/uzPh9Z7rclwydmAQokwmkqeKNMGrOLQIC+VFObzuOWGSxOA+Aa
aFI3LMxFJGrgOTAYHiKrwwYRTy8yMp/oRKM7dra2vtZ6fbS1EdBdYKhcxGrhGXtCdhlq1WFIQ6+A
cDvlJ1g3Fcdm4lw+7VblXl2rVErotVieIKUoI6OnT/Ke9oywagkBCwu8lkH7fI5AJ6BbVf0t9Ivv
jW5sk9wIchyOyC9vAbIwH/+J7CBd5ZLNmqLLTwEMM0W4/cqA4Nk+dJorx5TNbXGlU1+nDRTtGMPY
iAKBDvQ2vtyXzOLO/wmONAjhSGpBp/JcP691WeRsNHekA0Mr69/2KoCIAwSMCmrycW/j5yH+mXoD
5pzzx5C6gS2/7Avp232J6mFYitpXXkVvGgl7ofyNwB2RzuriSSdZjpUwhT8Vpqt6Me7hShlAssS6
XCGZTpbW4aCxB0m0CEHzyAFhEBXYpGN4EnMUFukGyqoa5ldRDncZCgHkLGSO5HcrAURBBir0HGRm
24JMSUZU7m6axTGbV0Bd0U4xempt72RfHaCBKzrwb6RaHpGDeQkqfScVbjhiDohKsbx1KzHdG4rS
TGQUGo4EsfIYUMJZ0DSCtQQTajSSiCI1gFw820JMcrRKA4GBFRSTqhaE0P2EEBW+wEKHvyuMvfSe
yB8gysB5pm/m6cpCjv6Q76BQz4WZC1zrHJQy+2XNR1hqkU6Pq1UR3YLFaXDpPGrcCg82VLRYeXo6
UGiKXGqGFl48U2D2DxPn7kzXDOqQUzWLEnwHVj2qSbq6NKTSKrVoPzxGIKwkMkDEaYM+sX5MgfeJ
b6LHuL/hLFfo9tsJksMs0QR28V193pKMUu4WqFEKMIsYBDQ0EltpH9Nt+Cvy6YLzb07xxGLMMhhp
22p7D+m46Fl7DlecFuaMA8BAcfD84qzu92G0JOZOx0ItDcAsM7tq9/rbSuypg6thaepjXsd+ZeO+
vwu8O5ZMjQsoMTuiv2RJHXrdRe6UXQjZ6cAsxBRrovliKfSbB+FcAkCa2f7quNR6fEDG1g3eGg9k
La308xSCXWODRFunC+QWzRUp1/CMxrg/b0NIJxu5OT9riyX9HoZM5dhDKNBu1GWOmiNVI8zh9Dc5
OJmj0XAykZOLpK5vKsXovPXEmRDlBxRjBs5Z68FPPswBfOsQztIVqtRics0pzqgj2aN1rPtmUamR
FdtqvL1Tofh91vc9vHTr93jex7tKcKzpEaaJSGrFsAM1m4K0K4pAi0pI/UyfGUMLEaIyPZ7PFZ8r
IYVxH1gugVKcFgEa4UjBSGPoeX6pof2a6e2mcxlmTZjbXX2km65O8IFegWkY1FoSKAOiZK525B6b
oqoQZ0C8T+pUUukh0zkT5V0ebCGxIIMsyfMBT2TuQ3FMphS+401XrOCmXo4RZTIuZo+GxS1GKbUi
TfNPMRXxA62PaD487h1N+Dk2Er89jC630CT/hjTDWLRhlH3Y76T9LO0nqXL6UZelunqhCkerox/z
8BkZqSBwK7JcOfP38U8No5IFxXh9MPjvGbnm/MQrGlY5U4XSI2r1/qmdeFPzbzTFuKRSy34oT5j8
LyIbNS7w/8wvC5kSZMbEEkXwe+grEGl0Eh8CEcniEIgwlkvv2RjrDOnScsm2Z65OFHbLb60wFfW3
17+7H1MBCROKsSoX6xrRKiTz+8FPK8nkrJqMD/wZ4RWMqoQGX6qrFccLkwUrV23LPAKYruMpqvEA
r//W+2OFrrbZn/VAAmiMQorMPfYm8cT/sgfdHAoO/ULzk+Ec5+YHCsxSgd+Y1s825eucQzpZhrdG
6p61hW1EBHXkH/yh60YA5Jffoh4p28qF/QDnhNNThNkYZZ8zsYXx9M0tAC1GVDiT6LaOI+XKv1ri
h/+NN8zrX3Y8Ubrwteo1LWQuPID22y08wBiHhaLVCznzrIHVJkjoyr41YxJzhcg+6xmABnLdgocq
JB1AcK56lfK5HrK6ZBzq9MTEC12/9G6bn9Rajxr1hykUrUP+GbPLy0WSjuiwLrhNWrCzJIZoemka
ipDZO/q4UZLw3X4l+7viYoYbeEodtSP+d0IwTtRBAFibW6VJk4apMZNZKs7RBEkpn6lXpsKACc7p
QS6qo/sEu2Axpgn8lZla8wRGwfXl0692dJuRG+3IVy05v3fgbq2mSf2sBZ9OeSM6Ecyor3FIylT9
TzcYIFRmyHjdvVMWxKs60/2RZ0YWY1OThC0Jijc0PIFDsaZ/ICvQMVeWATJJJefALbtDFg3b1haT
Nw6eUnGzkfXgWK0hkw+sBwo20RG0sT2oe4TNxS+Z7mwJ9VFT8OH3eS0kAQMvJ+PKIdKBTPD7vnKX
MKzaO9dvnlV3oHwwmBlN4x0kx5IesPxIWAsH/9C82qlLnNwTy54UPPwpmqhRotJchqTJLr59EvbN
n2buPMkzx/xohSmYdyrPGL4Z+oLMJlq8aGK/EM6LgYLObMIFPyUYR7dMMF5vfqgXoLiHRrK465U7
cZAiGqWckprjBOyt1yVAqKWB+q+SmZ4eE37e6ZVwXYJbXu2PuqZjR9LX0aQE6wm7XSRwrhn+UDxc
oGKaFaWwbyLR6q7B56CwoGoVCD2+w+3OGGSlKM2iOR2fpO+gmXD0wM/RZosCd7TLLtqtmMKn1rxE
21GMU3Xi7v3qmdH81n66Z6RuNe12vpXKXYt/qhAc0+em/0UBHX7G0Y0Hu8CXVHDEcHbZZd/oAflo
TQkDUQc7zRhAxPF8aqIiAZZTy5QkV3brzF9A/10GC9gW2pwsWiT6mkGa5u83zpbpsescvNxnukhT
J63uyZ8Cb76Vi5c5vHpNSo1IgtemV5q+mm5sscZ6MqHvD/fjQn7h4lDb4To0SyXS+igOukMf4kn5
z8hLBolIrJ9USloyaNGby62m7AYfBtYtsDR5q+lQu7rLUKN04xK3aYsb/ko/vFRmbdXFhmrElAWs
5qrOz1L9K1LdVQb1FHqBZp6CGFkB8iKswG9EzWYX2ZOeNXg+MZ7Rew7rDa4n3fDWOqJXiF/ln02E
SGvIgktsengdT1Cdp0Mpc5inJDq58p/PcbehTHOuYJVeKx6dv8dOYOTjnnhZ5NomI5K22A9YIN+D
nt+LHHVSJ6gnMAVroqShIqEsWbrfDegw2AGpIGqvlsYm/PA2IhWNsesDk0PWxhcO5vpzF+fScD17
AjhHtKibETgu12yktHfLokrTIuAsH5MuahybkVfkhAZxoCraHTPfaYo8hyXQr4v2c7Pp2AEziRMC
rLhfzJqyUboyqevuJtRzPN+SPKn/lJ6L0cCzU02qWHYI4b6/WE+cwC4lSD8fRAJJXlEZTifpeVCQ
0Lfh7n4HyVQ+PKBmEend8f3pZG1rVOJTOV4AUguAmiLv5wZoXaPiUTR31Rkz9TLbELBqJD322ioD
s8rYq3gnrOWO6T7YCize8hW0+U6XyEaxya7Mu5Ltg/DcSuYOq2RMBznh+pNBEBPso9w0C9/FXvxU
onYdFQow/BPJKkc7By8OK8Sg/3MF19v8MuHYG1d2UkHrYh9oT3QNwosSBFaSG0RhpUmIcQKigoqq
v5M3iHYPkV9LGJ8glAAs55LpRAaQX/g6RmJk++HHPeQd8rs0FAcVrAG4PkfqwV7GFmRRdxtB99+g
CuI0ap28SEdiZm40DhF9NKDEfR4t/Yb8fbvhGl83sLme66rABh9P6oeHIWvttb6iBGp+6/kA04bL
g3SFxy4z6EH1QYuJH1sMebG1DnM8lKjlGNULhFN3S7Y8+LvdFHqQ5f2LRCcNZJXQXbTLeGG/8C4S
irGxd0rbHmZ7h/0fgJaBMMIEz3SOCleIWOFT9jQ5J9XjMjCbzdfUXhs9GQzve00u7jzSiavbUAGD
svPCIl8hdBuMqlh5kDBpiLwStZvoAtKj0A47imXjYXx763KUU0zY6ERczH2XhMRV7Y8eSWrKEaad
W5DoxGYwNRoa6C32jimjb5GjuUS0SmGwCC6JfQeth7aOI8SCJfUVwkamyyNJb8uYHORBUOubWsIe
Ly4u/K5ZrOQE/xhdIuT7UKnXYWLi07Q5Wv23AWWi3oAsJqaSz5T0BVxDIcHouOhgQ3SY08AxoUTZ
99m18rzhWsJ5RwBaaeLcwcx2hY9WNMCfWXS8/afgZYk5NlkhmSqKx8sh/J4N8Wmvf9ocndcJfTHI
lynfwWOMuYK3FPiLAc8/mjL6CXP6PeavzjPSrFswVJ7p6taKmLfsrpeKN91+fW8yV4sOX7npB8Ul
jcNmO/NSdOJ/CbBENp3H62uWckBju/R37PU6vRhQu0js6DDC2I3kOqQ0Salq4WehtTdUuA1Wr0h3
cVxRrTwqWXWpHrO2763L2upMve9oVCdetcYSuA5DEHLW2ON7TNQUl2OIn/9sjDcBZMt4IJBefnk1
NrbAWingMwESyAbvQqYMv1pfBTZOnQ+c3GJ+iyHdBQmopwq501sD3oModPG77WitizT/or74LDcH
h9cEUwRr3s0otyFe9C1qDvBxfkwBk1MU/M+Q2M57qzx8q6zKP1rdRomVr/WEyXevSxg81tlUUFXG
Oj0PznqFIRZJmLsmmp1LEykc4wnQ2/ibejiGq64alWe9EdHGvm8p9I1cOwOQM9eRXnNA7GOT1je3
pi/FJhJLo+hTjHeuefTApqxp2VVuh3UXM7pX2RCZxtsnknWBDqdvQmEUOLif3BwO6T4Php738CXt
0U9sqaYz9XZ7icj2SDKXOimZuoB8POx2uq+Vtt1rBAIBaQMn9FBVuh8/LcZEJme3XJbkP/VGnwGI
PcM/cbLJPYHJeNqNcCtKGaYV4P/JeqrNbKIDQbBToxM8MZb5gbeQpwqOF1zLXLfdCA54O0yasO9N
7kRdmh+4eEHk1x0IHYuXuTlPW+lc+5CJO555/JqPlcUR3jpyaWP63Pj2o1ax6uChSJAEdA0KWNEg
PW1wi+/ZwZQvIZ2HFPloQ4bPc3kZH9oflkkTkUbn0p1L+7H60OoPXOFLO5QQE7LCNjT5kxbIcyDI
jdGi99dM+MSXn+YFFAeCrnVyPrrUPEE7SXGfbL+KUgGwOg3WQvEnbaZEkQyy2/k2nHxf97PIbUrf
CeB8XcNmzr5+f0psINLXXyYaxYVQgtPb/bUFtCQoRsAkSzq0O9plod1UIDyz7U3DVCCYVi043s1w
xINmmNH6OOI7Bpa+5xnSKXQoIJRb+xmCLJQbHNNlhpVqYpNCWM58NMzNnnfbNcQ4mQEb6p4Aokmc
9OHm815/x6YmTnY72cyss22Zjja25FGJBVJiNZoAgIk/Bh+qkOGRovHbC8XYLX6mHHaa0nJv8Vb3
nz7geTv5JiNMhayB4/wEY64AjmvpC8qnMuVOqn9ic5+yyXE7Zy2TUd2G2JIRvjPTfbGQy+Se//UW
dI5us0zZE5HcDj4AgpISGDjz1fvyL7GC6VdWqRANBe2a+22SOV0kn4Xz8LRNrVVXtFvsBj1PnS/O
dSVOdH0bUB7kG/amHeo8r2premXQSPaL5P0OKyIyiPj3xQVie7BrwxZjBPkQJwxtafb8avWudrdl
umlqJ3rckl8D/UnBzEZlXw14x8ZQh+PI7djYp3HP8Lg1rspQZieDHf2IINCzbXQhVPXTZCjoPHxw
0kfxSY+GvHuQ9vAQq8AbhB88F/Xvmaw6DVo/iOi6K38miv9pClpDdLWGztOkMBHIUj9aODJj9U20
oE5pJrK6v7PGcPYkih+kxPZPAK0qQqFXMgLZCpQG4Rnq9LtdH/xkEpmI9D1fb1qpkRaAMHCnfzpB
z7dcXT0DxkiPvldyd80UrgfoauY5a//FK8AUzGYZ9sqfG5XFc4R2pF4VMloQkeJP2gJTYIOXptqL
/Nsm9xqxmlDh5FiRqRMJgIU3qBdGoNBUzM+Eaxy9o9Zdyvjv4H+SFWNsgPr95EfIojGAub4QSwuJ
S4+x6FHOXKAZcicYtTR/6D2mZo9K/K3Z7kJGTpVwx42RZJnwy8no80xpuoS+t579uRvW+NCEYdNF
yq0Egfxp17grwf8lFUFy6gyeysKnSMON7yjSR+lUEcVb54QHKUwq2thfq9gOOqLvGoK6w1VHlVjO
TXD5yIjHgMVfIqxgALHQxKJNB+PkmZ7fGd0MPZBBEUmWIeRwKKX+quaw2Mp7IYAbm+VIHbQFToUR
V3YYQlhr96qTi5UNVUUCFkyR+cofFP3i4Tnkq+IVrjlqpQR9mzrf2xwUZIFaD/dAy7p4TcKwwzF7
YBCOCYEh6B97WSqdBZXDS/8tlHos4a9VhbqDzeHiIoyOrD5SR+R3DgraK+4kg0mjO95knEzAV1fP
9w/iA1tzL6W0vqWeZZOXmta6JBgyYej0EFy4Q0vDVhZmfRraFRey1q/rjYorVods5libJAoL98qX
aKiM0cabem6fLJRYqhq6JRZKHjT5JCtqHCNTITQzINi17XolUwHKDXBTOrc1JLq9AzttCdjB/21Q
xFzJukp87zjO0eRW6VyCHGWCDqLJ0+qa8tsV7QgrcfGkvJMCLIf89bmeBsH4K+zp4aIvY6bXS2zw
RS/p7K67qPgU3Q/sHe8iW/pCJ6NZCLAxhGdczSGCve7GJ/SNLBIyvJHNcZXf4BB5XVZFCYGFQqh+
PRBadLiv6ok+RwBMw1FXPoQL+BDGCA0fsw0MulZsSGKZTOcp0oittCVDsJ13/Hb5xTTTxDqM3hy+
+x6Sj6WAm1KTcb8R5HrRKLIKOHVVj6uynBEgfdDiYc8ORJsXvjZwm7bl73STRDMlBH/tcgfxujWp
e6796+4Ey9sh63RPjSj8WR8Db+LDMOMyhDdHwsQ1hg7nIvc6e93Q1NmjrUUoTWIeUcpdWu47e/vF
J9yK759XlefgBlphxRpCdBbfNWgzKSc+vBpWwm/h4Ccis5xiOoe9xmh4TB3v6SVdxW880qkjpzQS
5JdeyD+dBzL7V3JTmc5CybDy+3lAu3YP4OGkcO8NFT+iCW29yJEGKj9+xYEhXGRtJpShvyQeHJAe
3tmUcTaeSCVuiB7u2ALkAp4mpalAdZM2D7k8gg0VvS8S6/i9wiFUkQL+Tkh5wcUO9uDQO01Qw14F
nfjfKXzRa2/hloXYFcV0AiBGuyAVS39+Q6VsoWdCQQTLtKTLtUfKgDZnTzplSN8x4ZtxakkDPEMs
/lmdpNHWWlFFogU5ztjSuQ+eGQia88X2A8yKRakI18T/mlqY+vA2XI9Cg0kCyDOgopSQM1IYazpI
2/tLTsFo+6RyW9cbOyy8C4WvRI9PKfEak8f70KYqQhb3ohktdOSlc0PjzEGkD/hH4KS3CyppUOMT
E6dMHd/EYdoegXV3b7dHft6cN5hRd3pz0BLJ6/ZIvWypyMOlWfGFkL2n4NRW0803imK2zuEMj+aN
kgzXujwse/w19nDPcIXX8hy9MgwzlGNbSJrenzKpVrQBWjV6ZuYvf8mxAoziZ/IbtGJboniiiYkH
f4ZS2YkKBduSzMUKLetEwPhMaaF2ZsgcHHFyu8nRQDzC2WLlZpLTCW0CQ3Wxijpe3DYZW66gP0Dr
HH+AQ1j39lPJkdD5Wa602OMid7RA+OW4MIeIIDN7Koyjm0DSxrQjxj4Oo3pP57CuMaAt+9lxMpMT
V9nYzJigchQsY+C0rBcBht+RtCO6W/W0ZV7Wcw7SnHtys9WwygRoA49Yl5KDQTtBQsnpaJ1Bmo2d
mOc7zEGmS7QU32DS0kFzGrfiEGmFbfXJcuOg1a2p7HnBLO4e3MP/EhSaNU0ujpXHQPvTS/utEWWL
nqH2UdoXdl6BUEI746c4K8BYuMSwWGFhmnPueGws+o1VUK2yLlK7P+9jpZDgXjktxJSfK8C+zAyq
j4I/54yId+RVMqtbR8nncPokpEm1Ql9MqniDAZ3vBAGfG0mHqeDk9z0M41q4ZTU9PXxTCXrPlKa/
gd0OMWxxrG4fWe1UpNtNjAph4oA65QmdbU+l0xDsC+/mCENfhxYOwEnIBYc299X+jwCKnmcfu6MS
UKXOUUa0U7iM2L49aSw6mO1MJz+gwn3RCxq5cOyGfzPzrFOgdIFxtRO6HUNlUmGu5AoInKC4YFOe
hxhfu/V+VmQFWxDsnsGrPXTBIU8Uz8b9/Cob8qRA/0fic2SSajS8WQUnndqIZYZoNdlWne6gDHSh
5ApUKyhYCMKbE5dkF1z0HkjnQCpnI7b2uM9c9hcUZ4QAOiSJ1ypj2LNDZSdEx4zS3fg7b1oH55Ac
3KkSJJhnCMyBTYFGWPIvX1VeILTL0sfnS6NSD0WlY73Uk2SghDkld32+KCjFbXgcb4Vx5S5eOLX9
U1KN6gn/RAKLdBbS4jkkzlYvLbhuWwE80jto/fwstnFbLjrsACOSF0wJbW4WhXQ+MwpN4yhqZFnV
yKIfVJLJ8K2KKnaWnHO68NtddHvf2sdRO6gjpQU+X33l/JmWO4HS7EyCCQn56EQrTNZHO9M5Z9qR
480tzenXrelGTXH5fHRP3TCxBRUyGpr9Ylqq3nejgzYUcC8avJ9OiB9aTq824GkEDWsPUEU0Pm8L
SgWYIJn7Ao5bKF8aCbz2yqDJlflVoRTEgG2EwSlibCyPg70YaVjRDkjbIOt+sbB1fHwUmjMNGF4v
SFFveQVs6viPLY2YIdxl7vFtyA/DMmoFnuiiSlrCNu0w8B6VDfuwqdq+qjQ1NDnhKt3f8gkRs2XZ
YqBTPerNWtxvx/q+TI4XVx+xHiDwd3ErxWCjqvFxBtuBEeevM5XiGeJeXwvIB+g2VTvU5zpQlIsJ
3mGDpIcriqwpo1ruvRquROWRqRc6k1acf8p9+7s6FXimBQlO2v97AiMycavzZwy2mwrNh7B5C0hW
xq8Pkqn9heYaYzvP6x0qz+vk4dMZbAhTq/7fM1/57LMk6R7+LX4L3l0v5vlXttntMUMrmbf9T/hO
ZL6VrhTYdtAcm8KLZuNUWf4yGkq/pXKCrFVRYna6KDLT2cJXBLKuxgX7LQiIBkHXThcwUaFDEJ81
l7GUMBMrFUeKwVOkieES40TSXNv9ox9SQVjVDs40NnsKdwGWsXc/ERsQYYvnepY44uowLus88yBs
hjA71X+skGZxowm4pwPKrw7k5NZgk8RFrVH5akjD5MQhWOEg+mRdD5uDxEn8UOu+oorLAtfYXz7N
OS7+Y2i3A0WAK4eSwhhg3wMigCScY02V3kahoQMBV7Gi8XWrEsmNUMoHB04WycU70eX8ysuf6BGO
HvBt6jiPsc5E1Z5qFPfOd1ItIxg+4WVFC5CdlsRu3AGo/RicBW416DBTDq+OYspepcwHHLqxPDVo
YzbQYYcmVPDCNIJDsGIUC5XS2LwkJnUDPwX1kIrFo3D3gCpKKYF57X/mq9/1bOQo/cph+LbmNkdK
leVVUdDSrGTIlkNQt6kHDG4hZH5EAD2qW9RKZ5/I1vn3u6MUyZrYtf7TfBogL2GaG1hsR03bnn0m
uzZFxcPQYW37kMJNZELbqAGr7J1PccG5fNDZgMSnz1wr57rNdBT6JjHJrKOQZgfGbv9K/N5PRX6n
kVmmoRndXmMfCSlSxjfxCDK0p1b40KLELEo+U88l2g1XuQ8nfxJDnoCdwQyRU8Z5np4YtjjIL5YT
0yTW3Wo/HLK+KJRsCD49jjzcY5hVfEjY4VS7xM4Cc+TATSGqgRDB1UQgLhtVmIKqMRf4fL1J7hUP
b4OHvyMKnKw9x9wr37IehwA6S9T4e05WOSAvNfoytNGkUFcXyWKwaFLKFkai/uinqwmEgJ/EpP9W
AZ9+0FiY2mbOlTELEN9ek65exrHo7W+zRCibstIFy6acD1P/wtW4Wgdjc2aKNTo3K2oAug4p8gHs
9U0DbQiXjLGxVMgErS+sTHqu2AM1xw8FCAz1CA4SWuaAmfFbdhSVSCq79krU7KInrQQEdLzOEYaF
j1HOEs7C2RY4r1sE/8tuY+whvLZNYUQOrw5+TweAzWH3yIBHvL2OWvFLXIdqkjQOYakitPhPRTf1
qxHD3iT8tuMjO96x2wtPRizAbUay73WmvM3i1Ecv28WCn6yiy6KX2S271NhfbAJ464JR4ht8Mdkg
ENfKhS1wJq0/+Se8cL0bbONLwMWBSEMZ08mTYi68yR9H1yuBKX9VGrpA0uYmDv2zVP03GFfdywE6
Gc0p4lZTXIMLJW3hs5TmFFVHojbB9Ew8eRAUzzGNcrsNxPcHR4/7mqnOJHgVzBvG53ArovouElYl
VfBG9z1EdUKTL74zT705zDZmTnCMZvjutj3UBZ1FFAwxRGVhhObTr4Jwwq9X40yvp+l9ANERl0K+
i3YrMCY6YcMR/oKyhN5v86bAB9dfPSIRv8txig4Q+VT1KEuS90PZpR4wQu+kSHABDtrSj5qQp285
+KTfIEB4jOeYUX9oS/NYAKPkeaec1eRnIzDEyD3Gz2IkbAP6J9eYkQ3RtueiE6StHKIPDYSa+Q5h
psEdo4ls36/PBD1wEhkQ2a3ckDSdwB9aIYfZoKr74luYNCfrri8G7E9ikl7f8kT6QzgMep+3pmmR
3fRzHA2Jl5D9FGEJir8t2hE62TnSa6VvEoKnLR44JakMRLIr4dPoISgeH0J5AC2YREAEmle57ojR
LPAcv9q9gLgF366Tt84MqlHFqg3zZcyO6S5IMJP4T6csGUhcK7+zVd8UUAwRahAw0ywWCg/+u9d/
gjQg+dzh1IF6LwyJT0hyUBgr/Nm2KZJru+PDQBDOXx06jJiwxerG4xL09LLG7nb3O6NSz4+0aMe9
gYbEcXC5HqQViNRIE5GWzXx/GAIpasfBR8jr3peu+eIS1OmHFCkFaGX+nouoVHhrCoGWO9POC2n/
PHd6iy9HSeg9EBT0gZ/IsBS093Eo0eyQ0BP1bsUtw+NzP0+P2P/I9QPtob5hT20KXV8VZCDgQ1YZ
qXNUwkWsCgFLdL+aUlvFWMxWRFn0GwkdP6YEpZKOQc7BCdWMjgh+TigkwpNVd1VEZysVHl4SiVid
Kehf3PH4wnnQ0HSCDU0u3A1Hl/n/4GoPbHkXPN4aEGKCy8X9NsOPwhyz15KlTiVhV8bSq+tKrTYu
j978BqEkRte5Ex/2HavS2k6htKgd3F/2jQ8AdL39XdxdnwZ13jMnBrrQWo8VxphhfTawO2CZR6O8
fnIocQ3uqLjyQgx07EhpXNLl7UwGT7Uk9gVwy+VVkSc/LkzBdt6MHVnjzGJAlLy9cqTqPPAV68iT
CZZTypfwmq3zc20AC/ZFdEz9zyP0zjeZOgE7NKe/Q5MMJ9T37sja1VA36twYXDBEsZEHyD+OZy5W
XHYRwQSIbdEgnBrX7/XxfXv1/B0S+e81IYxH3m2NgRNd9oebtVXsZkT+TNiYnfFXcTujPUzgU9Zy
n6xtdbjSi4Cz8TclzbjQ9Hr3OENujveJOPGQNfAj6Pr/xtr+uVKBccZtqrGbKD0E7PUO+2p2CaoM
GgxK16CUbrjsHreZU3tO2njkDV1IdA4Jzq1ooeyPr5sBinNytS29IvEaUKPcpbQFTsyOrzVaKPmx
UCPGBRFHuE+yl8NWDGLF+7fUcdmlesvrmaMhwkk86HpesFoZq6nwadyQt7Qi4IsR8JYg1pGy0RGa
dLuUk/7jHz2x/uRa091kRmgT3UMVJATMsBEpoGswQYxsvvzdCGAihQiafVTxje/PIr1Xf/bWlod3
WT+Ei2Oozum33ZczMmi/f57Nwvj2h0gP7jOb+wAhjnz6K51ig8Y4Qozpao0rOGWlYVXDXWBy9yrg
taVFa3xxqJSV/mv9V5UWI/O8/JpbADNiODgzp+DZTgXrRDlJta2ejc4vCay06UjIBOdM1rt+OT3T
DDBb+NngNi/tYeudkRRwekvC01vA4N7xM0RNo9ZlHTwZnp+9xFIsTeG3993JN31xWmJeGVyT2eb0
SLKGsBVVePobDR5hGfJebwROne81tGWjyFSyccmLmYH5SvPR1d9/rHwW0C7vjZcUF12iLoI9ukh8
SM4CSYaoqfFQTXu/a/0QpuD7UjbOBGX+q9GCW+ubE6hmrNNrl7e84iQuyHZOS2alLkuV8hAsO5O8
ef1PMHa3iU7vSKSrLyq/j3EBrZZpDnbY1sdmQh10NgFcndbW/Ur/VAzZc0SJSzF9t2VkIdy+z7JU
5Okb33gL9QD09QpTcwfFYzoXq2C5V1Ijbi0pS6PYaRajlwtwvvoAIpsEY2MJE7JAmQ59eZ50DfOE
7bKwkdtXwIgeqoKGF4TOix4p8ZCqrzEO7nr7HSXbribR0ml8AeOpVsXwjPx9TZ5KghZP1vK0nYXP
71RaCSxVtcw+3kkVFTXSKoKVRwdNvkfGIR1yvp2TNVzfFlStRl9X0hbktIZ3oJ5RbVdh0/fkEBTr
uMHZ25bfsS8J47Xb5qtbE/QHFeFl2xRhzK/zomNUcqrV1nOTGugJRYrQqPQ6T3XW/JAKULEYgtT8
b8JDsniqhnjvk43uFhPWvoohZpu//EJgL2yDkO3oGl59a0tIlQzHSW51hAeRwKFVFGwTu15vMuxM
jtXWpkOZzh5wZPty0v654E5BW4oVt18P3qb5HJ6aLn4qBxctihGrWIwFEqs8ZHUiGSt4+VTNAe7N
vIKa1dGSl2UFwsu1NBmGRCVDpqmAtJSMTP2l0hvGqa5ST4kF2O+ORQJf8Vh6zmMSUaj6WsGRmWZD
2ymiIIU5RyjlI+0Tga4H4WwceKyHcUXVtcbOnLy263zHLsnErjC6FQyphWXJbKuFRUezkRzlFQbc
vDmi7P1ScdaQBZOCc+T/aq/wFpSzTF2ySlU2aaanIFSwF+xXtZUJ/w5pLZIFnI2YeHUi41mieshy
/xHvsMgs9b3S6OcGORNw0wmdvlNUfiUjMg1ouhb0xewL0oYzqOvn58JPGnTyrfmCkphF6cbczMnx
NOUouJFAl/zM1Oww+x6CNxLmCTRQFPcZJa3v+PEzsY1pqlbcEQ38qDGBggRgd87DboCibplMR7Wj
gRxP2CPOBJre5eIAaSq/7HqV7mw7+fAbwUBz5B1riRW1a2Dl9TC0W4h+ZxKAl9Sa6hdWXSA7UfEG
e/PmzB/aOKj1OEeSSV47PAjMmcNsRia+9Dntzj9AWHDAohfJXjrZfw8nQIofDfnoiScQ5fyKTmkm
TxxrOBxr5ghUR9rlLFhcu80mZ6M70EDsg4uuV4VO35adGEX8eIkkZVfZtdTD56pRMoLKs/t9nSKN
On7GwVjGdxpDZgVjySYJ347f+PSE/uLI3H3bxzbxTPJP69OlsEap3RzUi7zlRaNf3Sq3OPz+aq8T
l2i9Fpvqr4Mt56KZCtItNykcFEw544onX1CUFEzzrH5s5aoOT2hmsVhuISmKnn+hUrW8xDPj03Pi
uzGCyRV97Qivt8YHZtW+tb5PLVcv9zLj0KIhb2PPsL5uO5Zzwild/69qwmRQ8iqRnk3/RZyjioQa
tx4KQitFWvk28hvYvoA07jtoDEFAACqeiR2G0UMEGP7qINMxzqzCMSMNX3+0oZj3rW3nahAeISUY
ILx3JCNypFNdmFeRfhToUP91hHqF8fsX/uWLek8vdsCvMOU3o9Wkc9ELbBn7kwVxt5DVuuuWMJY6
ALmSC05GOdiGcVx2Jqt4wlburrHIDYvvJMBRD81nxOFDnZMFemkRQy9vgWJFSmVoeab/evsw1GlR
bZPbkaDlfzidWo2Nj+1zazkaWyMQhE1pEJPG0RmU7ypNeE3GemYqzwdCmqihdMKMBKqsFZLLJnC9
Eoag3jpc6OhRtSG9ZlfckUaHoQE4psl4kB9fBXVu84U7pt9TXGJ/8+I2Kf/lkkfJ2vaxHM69oSEw
0cWPchcbeEAT1kk+Nu0r2VqEXuymLaRalusykjv4kbTk3lIXhbxGPcpT2LgsYTv6g6LheiACEq+9
zkAypQ/tFfXTTGD+tNnYQHUfEujtYR/3wybLQqpAAEZqKIOgGD378Y6LxINWxyFW2wuEijKMxfjG
j3yJa/IR8m42cRyoj33MmKppaTBvy30Ry/9yXzLsAcDpmcliMJK5bgDNfY6XsATS9RsrEBPIbNqy
pd6QhxceyZB0Gy5Ls7/Ey+olf4smzUP8TFfAWnXqnB0sSc+ueHqNyk4/GvM0RUL9oVwmtfvgA8xf
vTmt2PH8dTkVWZ5xthbVT51qhb/8KG6znDiRk04nn0OoegbOuEz2S3T1Lq35Xm+xiClx4LBhjRfR
nmjz6Mw50n2Sj/vkxzSLp4OXAjvZdSlF7STYL62ITseabB1jgKr0blhC1Z34kpPKteFEffGkNNlE
m9Vm4jBYL6KYuAvUvxwA5Lchm5LgsuALrwTgQuzfcyvi6BZB8IrrzTa82Frj8qL0bOJoiR73Nz6G
NTgegNmIkX0vNkcGBr0ZOmmT0g4y/H6Od2Nz4dZkoaoHlRh8sVyIx4AzwUTp5/imhaG27a//2KAQ
XK9+ov8Yxo5IpQFvJuAlO0xepY6bRDO8K5fbE1ubmQB7qLn9s7F6B3G3+lS2cpdJ+6MWHgbspawg
1lHpN5U1padsem8drwPi+CS50m4vi/zFpr57KnHp/XxcvslxBnxGp6jlx//hicLAfen83EANBD9q
s6y+fhoWeYmGMBhJp0LwgbjYlAWjC/hwxtOy2mV5AdJokWSJVjLxNtJFj/HYUfjcjmafj6FqjL86
62DYhOIjpJqZrjFehD/ubDARnGBnIwgCF9FSz4JNzJh1a/gBatLCafwR5GVoDyu04VnL5qp33i3/
89IvV+59cECIJ+e3TKMul6P3UpU9+w35POyOBnTSzURHVKEEPdQGtLdhNvhT/Fh4LkqzdJntQoH3
PXy2Fw6OFUWK5iKT1wi7A3H3ObbMMtsPtzRWag2R+OMGBg/FkBRBFmteoHQOmN6xLq6uC08caDda
R0jZaxolvH6iyvZNeGc1yKy8IRwFR4x8tTqqzqfkrsy89U6xzu7vo3r7nvaUKNfJEjuazy92KOQO
pwepKSjy1GZpUhnw1yXeZAtbaPNMHurI8uwN7gm9+5zlbW94aPlv1WYPOVcL/tI/PDTJOrcl5FWC
WZxXs6V/MWXnKWv6bFld3IIAAxT4MW7xBe4XOwwaInxmLMhePgfKYkJA2zE9Ude92+NAxakMrv5K
kgagGbxSaRV0JaeMDoZ5IWjM/UyaWUnG1C8TK6gdspSCcUSklk7aPZPm3DQHKZ/+xjAmN4ZRX0kZ
WxQ1bWNhFd3/nWPwmhUceQxN+tnQ1ixAB8w06+bvJcWqoq9nBZB+pmYeqkBJv16RxUsXuymtLZ2O
CdGiVbAWQ01NwDB+erlIcMh76qWSi8KPb9gEEAK4ceLee69j4d3ysMxooIU6/6MpObYZASnMaL7v
QlPuk5UvMYEzbyWiMJ4coeSCZJh+0GrzIP44RfA8jFJqsAeP7eY2v04SK1C9ye34ZiQm9hEeey/k
/ETuxj8XJluHxvCUtoNkS5cdustRmN4cL8WbiYMf+sLXT46zYNoFWRAPqjNfnLgXb96n1U3cqUI7
0pF5zSzZ2JiEQBwCvwOUd3Wd5bKE6R5eALrQ45NsnQgg8Twlb2sAuPxpak12Vh+CX0aej4OHXySu
YaEnZedhBXhQS2IpI2o5jM1wyk4GMlTZQ6fdQV48E88Q0xB/MvbVSH92KWjQ5AI3bu/XsBq3YgWo
vyPML8uFcLz7WiqrKoTCT5SWmnWsU232ZO+3BMPF/doRav30h8+uhQmiwr4dOobNFh16vD3FWi5f
TUKbzZXKjm8lRPdF8gkGB+vJs0/Z0JOXS/10pOe2z8uPzINJ+MssGWDKH8d0SDZ7Xu0K/Nauek43
0U7hUVUmqqPDrvzChDobzlQMU55TJNnCi6eQ9k339/PFGCxAjEKEe8fXccr0hTOoed2COfax77ns
GLUELIiI+ls2ffsVbpPdrAHX57D4eAwiO4OoA4VRPZ94Wub2zoVPxiXfK//2MF3OI3k1VYD2HA2m
YrlhYUNar6mDn3vYup0xSyk9IigN5mBENy6dvvpZxWwy8Bv0Jjt0x3GcOVzjGPMxCIbnapcpNY53
VM8w2L4fZP69V3rp1BoCVzF6y5WKzfWXj4FHNVtEfqRaTXuM14Z6hcsiK4OnwTq2bD6NNYbPmktO
1Mmz+ejccKiji9vbggxgu8/PpJEbFJCE1EHY9xIEFjl+ICa4ORcpg1W7DYpGMRNUxbnUfyz/0sn7
AZhhLq2dTD7ZunkVKg5gKG1X0yUl25X/zEWFCj2PYm3j5v5z1duy7St4kKqY9BoPQ/5zLY1ZlEDo
B2ftBUCPCOnVEnb2eppo0JmBDODbT15Pavg2AxiXAvNCOan2n30RYxZyiE6wfhGHv128QQVsxyx8
gxRTPj7OWK1qdCCjfoScJ0RSmVNebTmSl0G6FafWq89Icd6+kWidm8db9yXf4NYqPPK2hkHYFZyN
KwshT7YU7LTnEDZxme/ScJwAzWpOATT7Igg4Sh3AcK2RkeApSAl2rp5Jv8u+QEsErU07vBNlch9i
BO5UljjzOMor0D+nvXTllWwuboayPUZFbxTODsawhDaCpe9P+Lrc4k6NLV7a7+xEHr8ZTCR0gi/m
Nf+HoVWDC6mxiwFI1aMxhT0SUNfXCaeg4zYxYiYDTOFY+/Cdbvj9nnRobzmwlpNrWBZBvy9Z3X8f
4LkqRCGswh9+VQEK7sq0RD7g3pPBdBzn9OHqaKf+06VO8dh5LPph65plUp45WUP1gRZAtAZAPnEq
Fsuc9Wr3HSGC9BfYClYTJxDnAoeLc/0an8X1WBCzid4qRTPToaZgzbDfg7YR6Vi/VR/iDAY/A9wi
MujJL9nmBObSKOnE42QSJC7LYNL9RGknbIiECEw5F/rpKJ3ClfsRUaxhwHAcX8rWpHOjmiOfoO/y
vcFfmK5Dv+4nGezxVKAo6MlxCXsX9mrD6XXVWW+giR43BHg6H7a92Uc11s0YMJq0+cC6LhyqJsJK
QfWqe/PHDtHg6yDwhELsc0NcRnALdMBL+isSQV2I4isGpMlfGTpBSnPBZRXlttoRSKcjpfuqU0Jj
OnYVZx9HKm8z3jUm3ZPedLsIESlQuVBj2FXM6DM2DBdcYlk7blIE8BVGNF0mlq30zZPi9RuMJr6V
JQ2xIEnCgv+jcwoi4+AgS/EyNDgFQlsURINs2OYHw6cNiaPHg9r5qNNwhI/VcESmo8O6aNYVLqNZ
O2o1S0cqlzfbEp0R3B3rAOjGOwMLFtP0QZpaYaaJH+elY16t/TbjQDO9OxwKBkkYS7jX0Hu8pI+G
PWexitRP34TdIZthMc34ChtExGg39rUvVxfIhDERqnScfgYkB3kIfXbRup5jSXA8qAsC+Jwuxz3R
qt20mCD6h55bq0qnu7jCQHn86n+XRmMw19ygcNPpvEUI2Lm+zX7LeLnMHMFG5ShnhRZt4Ysv9lsS
JydV9gdtapvVefv9rFWh4dPLDm1OWIYFiR9CaxkpTcxpYiaiTU8gL8v5U3UecaUGmjhgCNraXod4
3+H5iUpe4kR7NWApNjiJQaRJjlUZPqoAGvaZoYf5FX25iJ2j2QVscJpv+NuPC9FAxzgr8xmdx2e5
gt8QhgPQYPg0LD0iCOOVlWGXLf8PvDWOOudiZdsOwi6a3fqtcCUwvnuAOl1NYESjGAvTG3Ys3+aC
vcvCm0tvf0K28Y4E/nVQiZccj40J4IBXUxeZk/3Opk2acLr7xYUV5jQQfmkoVzToJwKF3Yyt+ZaQ
ky/La+zt/TwexzXTVUDirLYluskOUkIkGbsJn5Mu33kXMLBWJo7HZsA8i1mGZiLyTcBQdvUbmM1B
M3cQ+hwR7108y0fxpXIDs++2r86yhhshBDNj18Bq1r6obSkT4Y84ujegjuLcuAivJGleRcZBuslE
eelf6qV6Ah3OGSj+h5df/5P2ddWQ1M/++AgN6wlVIenG4sEo2NDtD86YJlHEcLqkAiP21rjl8XyN
YcSUHMRuqs46Dzg8cUH0w6xZ+kcKjuVOrtTvj9Cln43oubRaPkPrLRGG4LCk2Lj5u1ZaO+eVJVQb
munY25yFNLLaLnnjeHeOgMlPcjpmWyev3wpKZKS//nzeoLKAgsh/2GwwJjkYelyZfHiUA0nl5PRg
M0nn1vh+ZtzL+TZh13uS305NiQLseiIRxB9xlcGF8UvpoqCX9BcODSTnmjJooKYe7Py2XcRxIe4L
uSkajWyt55jqwSQToWVsp3Rf9c2B2jsDmwOSk5ISR+gXJpWlrkPzsX40ZM0ZcTLee9vPY5rGQBeP
GHNA+rHyGMU9kObcwANoWV7iWize6oOAFhhT/wLlXvpGxc7H8UMqjA8dvIuz+MB+E1AgfT8hDQIw
qnWq+dPJqz55bVKlbR0sigxU+izeJBixQ5uuLYgG7lVs6c4GEVkAzjwQ4/uui2o8EGu0vyVdLlgZ
+miRdObM4/ZpLgaQ8NxuYfKc+y0OF52vCEmgpS20ti7sndqsFfNa3wQ+4iUDkicYnfqsqAAeoAt6
LEmegQKiDSmtwQ0ztZLcdnQkpjcmlCykpG5gcIoNj8odOtruNuIpikb1TyKRii2NK8sgsNYZ9Q0n
W5UB0ojMeE1U3cR9WTNtUmLI6M0buxxkLjkntAxuwQ3VqEpw1hGToQs9xxj1XjN3POjhxDe3r+CW
N6daemo+Tv3ylp+zj6udkhc3fYVL7+zmmBT8Ubu7QdR3U9KCaxjBzuiEusNGF7Sx//dWDGfyuk3l
kDOOBTAze8kCKEeOYsVBkhQStznd08EMZu4RRbt98WBq9Hpj8sFHRfy44PiUqXHsJKEb2iIRNhc1
JONQ0dObNpTCCrhKCjPCU60tEzhEKuBgxkb2YnOVmJNnmmHUy2S0E6iefyqH2dWA7Sp3R0dK1l1y
MidSbfpeuPXXNW7FNNDOm56ewgwVFQCtj0CxP9w2T4iGzLgiG71/dV/BE8Pu4UDZW1WTSVUDSeTh
DSsGvXb5F7mQf9K8lxUJwxoRT9Mw+Y9d7Ld3NswOsOjMIxVUSdO6jn1G1l+4c1PGcZnve8vM2vgW
9wHkkykRyJWTRElMwKlq5kR3l0XmQaFzyOiSCGqAmA8v5Y3mQq0vywIPSo7B0ZHlKtScHmE+S925
tZNVUjBsAs2HAW6c9BmAOqFYk7A++JosB+154pT260XZ5/0vDXp9Z+sgbiycRAepa0YPffdOc4P4
ea/Rzb8ykxs8YRDv9PdubqiFFjV7v7dEYXyLO4Esf6XGO7LzcXLoc7DzB8uK6FYxEcZLX5Vmf188
cFXgQv8Wv0WF05uZXVdkaeudlm0EoOsL6gMbc2tzDwCJuGOJTCArStth6eGJdwbmUp+UKHcmFR1a
JrtjGsyjT3FSKS/y+6LowsNZtArh4UgfH7k35S3t6SvmYwn+Vwv/+ruRVsv97yI+A9Q2wAWOZc58
VkiJL1E5tZiwekQ8RkVeRmo96DR6P03OUU+7Ssh+FIFvfpgV4/Fsnd0gs6IZLzzVkQys2RSET+HE
4uZVITmLi4GxUzSBGLWCZtryHvXTtpSzPnsbwWdOXm1nopwo39f0dEgQOrydzxpi3SS7C+aaQsa8
ItCIucFJC5DXM+V1JlUxpCnRSbEH4j+NDqfS05f+GPJvR0P8s0Rz75xrAxCA9QIeM1kqOzjY3+c/
4LuI/Y65tIdUtg2I1jTa6DMRgrzkcCXzFoscYYlC1sbkK7cT05wjYOm5kwmEBHUH4+OXi0MU9avR
8ACv1ieT499wH8x/C1um7eZRirWi8jYs+1Lj66BOIcN4lPxaw1KtCNoWZiOdlzodNSdUsnk1eF16
LD6vrvAdvB2KI7B4n4CIstDc8hKnf9j0b2Me5DAL2rfV+9YEMJqqF7m2+jjQTCyq3I7lPqoXVCOv
EcdtWAPVTGYrZnLQFRWiM4P9Vrnx1UXetxTTFDIjBpJjGF7hWDHnYZ5ulobWQfUIgIO7Kpei7Hf8
ZRhZ/jnaBCQUiWqvNdNCM2BOX45uJ5+E56Bvq/IL1JVfM6xXBh/SnhPOTyioGOo0XEemx6uC3P94
Bu5kOrX25KASCMVLaG+UogNbEdOV7yckgl0v4Jj5/Sfy46FnNPhm8sph22xg/LzRNe2P9AvTKiGj
/2QLJ45dgY1PPjvRKGhc3tt1QfuKdhPqB7dXMM/T2834rulayfi5M9yILAoCvSudSvjTQfU9FmQM
8Z9juEVnzgWJhZSkum7qcrFk+F9f/Wt+Ox3ISRqee/jUIr+KaRkGG64vKVFsOW6kdZF+NOHVrZwH
bVuowGDSV2fZ5M0OmTYZY0rbsqnEvd5iDgykXKPcxNNiaOaYH2py8Pls4tHr1sopmc4ifrupqMAG
ig+TP407Xre8KNxaWy2w3Bkp0UvfCSRsc6KEq6wT2c9iZHWqiljAFU8iCKtzyZ72tUIBd8sJgvf0
yIRhWSkrRjf1RqErVsHjBbvTxuN1TmIOjotK0Gd52G4mGnoDlEZEg2jOEM6JE4RXVCdgIEr4gV2l
hFk+pNQ+xkei90HCPQvngx/0raHRq6VSjQe9sJFIzxma0JQ0PNOuleINVz6UdbRDczikDjg7lDR+
Q4HQu2Ie+Es0rJSwKsLfrydk3YwMDj3lzB8UOH0UnCXr77AhbXUzpnsweafimArfZAShhpvwSkcO
QN8knmz+GeK7pHqf46mJwAfUComrAn9GjxiQ+IQaKwudIevrwSD4mQDON6axcEKeYqAsZXOhtx/C
hUS1vgS8ZxFKM0I1vJ3VBpN5vylRbcPuNQBMR02nCgjfFr9NI4Q3ZGA0HX3voV3i6/mP3Z2mJdg6
TK16sIPv3ZCSSdcXB+ASLj8W9YhuEo8jnGYiR4JxkjZtmd3isIKkYbVTy0vPPCg2WXt1D7UqYsiF
T8NY8+krIVlg4+53yy7c6kNN/5U6WBN6zJajBHhYDZ4nilNfpJYZ/jKBIUj10TvhGi+djXoVdB7I
gZa7ESgCciPnWCuP80ojdWCNGc5BR0Z9UocnOVFWhGSdi161ypL/Sw02rkMx9/fClH8Zr4QvQ4we
uQkcpLQrx1xLg9LlAWyYTR1yyxhYIckUBSRyC9GI6zLE7cp3UrLv0zcC1Npz9Ur8OsG4WXXXkaB4
ZuJ7QzOjFAz3JMyV4RZHKHXPOKTQMweojgwkY9bTgEAfWUijgYclLtTg/Ies+XZvH0r7Qt6Oco4K
FFbsSYECLho1a4aR4hNWAY34gVg/4ReXdxcM9/8O4nifyOj7eOu7gMu7QZpZfSg+qNDLU6f2Es4w
obEH8wnh0SPuPv7E0RvD93pu9g2PHqhtcanwlabsMRLdUh1zSOY+UdLp4auwjBgrK0nVsehoJD4Q
FDP2WUdB059qisnmyH3DJDjmkvo5PBoebKO9SmQFdpHB6AyXbG3+a3BSCvSwYIZxV37QkPVh7Voc
7wKaA+/pjFExo15stR8NQgUoqzIwrpHGDOf2GHv1Mvf0HjWTIqo6ykdjwhE5R97kal0SS/VT2Phk
xRrF532tnOAw+MeWh3w25vn3ZQQXkSRcnTmC5+Vpu3jmdGlQ8kl7EO8yWI7H0R/TPkjl2CEni1Ov
E2v+vDSOgJ1FBRnJtZc/aMKkEwInoc6QNAqbKG90UQbvASVWHyI1tJTQ8AdI/sZP1mvPYRkTFLST
RXeUxKNUZuqTNzcSYWG7QrO3CxkUJETo1PGblYj5SRo0NWgh5S/nDnSG1yfRTDfyrKda83V+ATA+
rV/KNNKpSUSL8h3w/HSnjVwH6Vx64E1Cj9p3iEARVF13wWB9uIszM4Ad/yJbjIYOBMFzLIDz3jf5
pA6IhTl3EO8etc9EHRVyV9FD2qD7KaMbQmnwygwMR1+IfOxbVGH3tafXq67IR5xYaHVTPlRahlr4
AUyb77ffriTMhZnlHQajf4AzjR4sv2sNcP4AxAsY1LDK0bsl3pbjY6cehJllVTCkOLjA88DtQWtZ
ppuxw7B5GTiCIbcq9XmriW91SW2VV2aJW7VHZ6g7Bk7M/UBOPyUbQ2YBBNgLbbRBVB47RF41zA6i
TfxlK6gguVuzrO8yTQC2VYJlOB5GS1/7s6135mbCRBss1Xyn00v0EgvGEgwe25zIRqOZPx7IdO8l
NNYrdKJdilkCRjeLSSQVquwIDbzrxMwOP/a0HRjR+4hQvp0iKozmsV5+xF1qJxPiZ/KOaAIZ8XZQ
Qqz/VBaZLFd6Zkplp/+i+pr068zKLHxG84NAHHJ19el9vcIJjJa9fCLLiW6E0C4uLp7AUc/FxV7U
re9TlpQDb9rFBjlCBX9n+4/5w3taULAoRAMf1zsryBYhEG9Bf478w4uUCUt7YEzgX2kj0x8lTqze
erFBjAgwYLdFjPq9svAlOYgngul3FJlg0DojpmxP+l8T9Jx9IOhEAqAfSCBDgjSb7/1uC4sHiSPG
643tHO7W3wRdlYxzkdkkSaoZsD/TZ5RF0ja+93aRM/8t6FLdb155i2hMbMnoZC2ABfWAScZiMF6P
1UoqaJsNLn51gICdIbnTWmutd/rd+OV4+usPirjg5sw86XCEsoPmpp4La/GEGq/X6snH5Qo62UGY
nakRSMZdeZ9YH19h7KtoOS9YUpSIAXGBz6GeSuFP/jO+Hjr8oxh47DMnYRij/2dN0CYi5eXztIqr
A3VAwF5UUNdsi2GVvqizokiLUStsBQd6ec1JZh+tFuaKbkfAISPo4iT0/jK7kv77KleUtKOoIsxE
5gZa54lQ5g6O+ilB6CDlhUkDKXvVOpzQ5mV98LYIStwbDttagRgpHoLCLRl6LF6yC6SfbkaNd0Jr
xKEgBxgs2xBEmkHukfQAETUuZdHrp8CMPFG82ovYxuhWwyH90+rxI4mT8SElohyz3fXdX1YRamIu
G3BfSPiv0Bn1Js7+1ozeIWwcsoythUmYP5vRvqroRZ8mhrg2lplhCNNym7B2v8UhgOterXjgVDZr
bmztI+49E+FNJBFy4guDWv2naiIOdaS7hOiFx+hR9hZ2gSRXyGQt7ECTTmD74IbCQvm3nzXkaJ9B
vyXdD8QGvRyYhq9cAPmv4agjFNrCc8YgM3epQ+ML3xKFapbe3b2X3D2/KpQR2M9G7sH0AVGzVmuG
Oj9JNmkgFI8dx/yirWWq6MxIUKFF3ou2gsxksRMOa+/uihfuruqYiVzSy/ZS+X2dDdginVSnRs+V
2RSEFKEORHTjQhHHVJ9MltX7YmGCSegQvKTF9Kji1xuyNr3UkArqNd4QyEAYVezYEnmcZ0EOkFRd
I0gosg5Ytg5s6+/D3kgXts+mun3tnjp2TI1dKcmifrcV7t3kg0lNl4vu+ph775M66AWa62rVRWwA
ni32CkAkWLuyN9vgfL4KVHc2gjPHpvMQHAcNVot0bPmAY5+FjT2GqwOzxH9laTIeyzuvPmoE6RPL
F0VsL7gfWKFgRLmi8c7PE/YruQ4eTY9QKK7EaUB55S94aZheHFIldQKgLs+k7ULdD7WwTda8ZPgg
IFRd/p2ha+nC9+/FyKrm473WZrTqAPlSlOOXvRAPu6g7XyVli67KL4iRmTaO93sW2oBy0nTQoLgU
vL3hTPBigMvcpyKtiYXtQovteKhoy9BhfxZnKVSiMtrC3fJSpGB2dMP88HC8spAFJEai1bdFLEHu
3ittyReuisH3R5yVxPyV4drg/TfwUsznKcU11YJySvU4xBBunUKOI+aTQiX3IncwXfulHqN65Oac
JpYXEgwngQSWyBx+diYRtCPIacv19bkBofYDTFqTK0YDsf/ZsJmYJ+V1raEzewFjxkuOdcqRoTh6
2rhgX26skiceyJfloHiNomfOw0GSV+PQ4mlfXUizoD54GwukNd0fnXvB7i9kwb6APEMbe3wvAUd3
NYeg9EiUv59F1EBiadmpsL200uhLxboZ0dak0i0/jTPH3BE6Q9Z1Z2cbi7wdo2JjnrAEKq3tscCe
WR3Pmr7IAhyxJnjgrBOgHtvsPMvBEp8QrH5N+rQobseSGvmeAbm0PTcRx9pz5K9uj5frY03hZF9N
C5KDLUuqnGK6k0sSL/8STHJVEjmU5BZIIyz+o0ZJiu5VwfHI0h+604KVuDYj2rfGL0Kunti3HVcJ
uHKSqxV9ebrf4+FzcKYmxMrWqJJ4rS8HaRvfQj8Lh2wrTuECXmksIlJntKjCwvQux4ketdQE2IEN
z1fCPOMYpWU3+ag1XFMjvdL70AbBNeobXKvvCxZtEt2N9eDSbKdLoyxYMrTJCGPZnYUrv34soJ5m
aIlCibm6A0FlskwpqAqMWXQhR4TSRJrkYMm4PriqqxcxpS7gct0wSEvI83h1GZaVHi75VgdTf7Zs
dsgxc5L5vOXig7rytCMQOGWnqlRLNP7ngnTEfNdfMxdskPX4ii/8kGu06KHsXlek9nVv2UTCurxO
llUezzzr3P63gcj41R/BYy4o9QUGJ86pRaWdh/S/HhR3hwY0MUYSwO9gPhteXY/iJBWDe+xF8Rjb
35HgHeagZR/BfoyShD126g/QQjAZ+0mF+qNljJVHpq2GQtHK4Xftk3GIg+uYUUE2aaBwr6BBUf3m
/Wu525QNtfYinBfot2+rkRP0PvFIr8/Ezp53SjW1WvSSOhoORLKccQ6oVG5KD7Oazr6MB22QfnQq
ruEikT/2O8V9WFXWpFayxnpNM8+nNdcscESckTHD0yeXpW1L1WnePW25w0YlzH4mRa46vEZb3VvP
ZqxicXmpUjwOQEcfLSLA19e/3E7jvpHNefGntuivdEHpxqtb4CkPCkvYylgiAE67zC8/C4Lli74T
B7mW5llsQFZleAMmfekqG2H75WAlhgPdQlTZq8KR0lsMR6IwIQPpg4g7msuzGbZUguyeUF+dfNPH
DVls4TRVzcRCz6d6ThQd4Fwaf8qbqJaTtNC4hACU1l22m2tiNql8m17kSQYYaEOJc7xzVrHthXG+
9tnHn4o+bHiRBfE7PU7VGDZQDG3BvB3L1K3H22gfFvSJ4Dma4JWR7Pw6tKtmEfs5ifWiaxLMA7I0
hr06CYd+JIoqGFQwCeMF+HTZoCrpNEzP3jFIHCG3N3+PKqzppJJaiMOj5BNUiP0sE+5v3wMKbHB8
a75345LOePjTad7AKbVwHWLQtlqKybLsCf9/A+HioKk4nPkQg+eW7tciG667/xY1s9Ci7UKweqoo
j+t9MiEddOD1JCC1H791y9KeHzKsteCZCpvfYcQIyhEa7P+QGQYZShITwtCUs2aqnIc5z7IuLqMw
1/XjNxHVlm7Xs+Wp2Mlyo+2B9RXMq4gieZG27vt1QT0GQ2I7jl/i1na94NKHWwzkWadklhEzrqrA
ZRi3h21i9thm1tbZWhOGrylXjdnWH3rVfEuK1ml9EO43p0MNDfSiDi86/4/B6CKhpyxHn8KnJfdR
X7BGjveHAB+SF6h6zH32pGQLY34W51OAHAf4CvDPuyn3Ryey+xr4Dkr7NGU4/kz8fAndrq/knDDL
10ZzgSrx3d3E14n7LHZ2EUhGGfPXTMWfeBmWGTOO/7FGghgRX8SkgcKfZr1oHELtS66b4FSkZa0d
DggFAVLv4xsOH8URfEOP7DxCdvEi6/wG1K2Ndh0my+PCRwdZ8J+UcHxZSGqj+DAdaLO0grAX9kT2
pRmbZVf0Q0RgPKWLwZWz3guQLCJYJDqMZY7KHz8nMuy7ncuU7TM0cy5DTt9n3eZNykEFN8a86LCn
JWdjuvmBgW/gCYOWNRNdNpgOouMEavEMua+Ny+gmLZC7F/iQbb9iovVmagx9IGCQ9vt1jnnfIaQX
d1v2+4pjPkZYBdTRNd974yv/zbfaTvdkmYbOVKVOS4VDFbXFHPzSZlNUyJhjSgQbdRhLhhVE6WID
3f9FZtjZU1V+iXtCS/JYJeSAwdQwvgPtSauInv9jZwRQ8JieNFTQ0t205GWQ9KFNGvNwOVe07+g6
UbNRCH4691J4zJCUfTYmXElm2xVDUy4ZZL1TP7z0dDfDLxBaodiQdhwYcS6PL2yIL2cWcbiPLCfQ
GugaPNKlRL05WotHS7h9lwebUT4YR88De2FoQWTV/5qep9oBpVIaas18XYcNeDP1F2zgjPmaF/f1
9DSO7vR2HqVVGD18I2VWDoJofW3ZWrW9weYUj3clpLp33zcxXlJzcLfF5sOOCHAKE0Lbg6Eg9hGk
lG2GPsDWdadOtrjEFvuXcGjnDHdqcumGb7T+xQPgiB2tyvL2kFjyxZzW/GeNoYsNaVfma16Gfy00
HRBNS8rNtkJw14i9ujokpyFds0Lg06zHjuQN96pC3J2W0mwTOG/Lw5T8roJza3+bCEi1MI3vamz0
371Hbca6h0GCKoIzhdeeWC11cWQ3R+DuDF8NaDke22pRmQf9gTC1mzG5K7mtXW3hMUT5CqzFRFjt
DDfnNZwHrX5XVIe7RPGu3cqcU/k5PVACH9LYriCDyWFEN6XjcZ0IltE94eqbQ0jxlK/TERJMH+ks
mpq8WJVphCD1WKnZS86HjlVvWPM05+c+msE1FTcKogzVKUffoENi5wtURq3OVCX+pQiuVmj15hOZ
u3j/JpylV5HnC0omC0w6xlJhRaEV6ysql/jgmJZAkxQMOiMjLPItG+8/5aE2vmyQX/X9XgRmVZlp
aDyVAM68WtNNzYvxwZjDeENSns1XKy0P3SMqNK2YXjX3FSyi3AKXSskMYhvJxd7NWhcwSTCQtvtr
HntK/QZ2ENDYRGpcJDGdYzf9RKrz/NJ5YLv1RvWbZvUiSVjslpTU9Gde9m+B8yGgkPSms47esIgy
POkGENbHnE8jfJDD+Yh3IVRkL32ouogIG4hEVJf0SN+GPQ1woKUyz9uZ/i+2w3VfTxNpewPrvtiC
+klOM0Pd0kf0PWpslBzIJwsbzFW5nlE/Xt0Af+2hjO3jBRuEoEHConqgBlU1hpXgO90+PILRfylH
2mUy0oq7jjQJFY3WDbdtVyfwHvlzUzde6DlfR4T0z097fFMcuhPMQcUffabHmy+EG0LxuyW4ayKv
ea8B3mYVmn00zXcWK2BqNagpF2c6Y1/M2xlRkZ4Oa5KfQqN3m3gnd3yeOE+JEsxRpbcbWT8XKRAl
sOTj3T//SrkVdfifXbHGjGb/npWpy14MUN8HGR7x+Mn7UFgy0iP9Ly5pJrDtBnwHBmO7cYGcMteu
W5gJtsXaksbqE2p+in23ZKOd4Ngrp0XGQmycl+GbeTo3MgcEwaV6gDFnII2d/63oWZgT4N0kwB0S
JAY/6+dEA6YL8QkYstaZoYxB7EjRNj96hW/rDqqobM1Qb3oh9ckz/1M14PCx93Ji0kSjIl/ZcHVL
5yKXjxQHe0eIOJg31BADh5BCoUenoZswtLk2DquCrd8T87l2E+P6BEPxXZp9Hr33cXX5HRW3bES0
UWXRvHwNYNUANn2gFGce9X5AO9Qd4LXveC6ukWRoEBLQC25IIYrjTMLncU4vyPl/sU9//2mX2K91
6UnID+JoHTukz0pY0ZNZK11wlazgZFu9xQQOvTrom/2c3XvNDVWCaFmFM4fI7FAtAW5yPPDO9Rxt
+s1xQNgPRFhXcgUI0JoAgcvoVSnFtTeb1iJdSfuGJDURPXQOLe0oNlM2bBQwcNF7OSA0jEIrZLFp
37MNYh9NyCSMdhx3jnp7hX1YohPWot6W8i4bb4tOrnI80TML9J4sFV34LalKtpjoAr1Gmyp8Ddrx
uTRtCiC2eABi6VEuVYTI2JWNXdx57Y9yHlZ2hqqF8RoLL+WA+VV2QHFiCYxGquyQa9Dof1Q/kbTg
923jVxwwrc1FNJbHrGT6BOGptg/OM+B1sjNbduM8m8TTm7bZqa8BOBUmyyDDau28gYE0ohpvPGiF
ILEPbGEWlG3Fb4/+G/1AGL4PVQr29MalVJvJFhVjp1zW9r5fzK83G18Tw09kVp8YdK2EATEUbCxq
d9WGAFNZCMyI/lcQp3bW9p5sA7gBlF+6fN4JV+mmPToyTk2UuUv6EzlFhs/YNfjkaxCeLK9UPQkJ
QRQWXQclxmhqe6koIOIpdMchJK4DsrYieQoMFam6ZRAfKtglbmsKyLLn3pPyN2T5Y1Rge+6jdhy5
MzhID1wFAoeddgxlPmiNt92kF5obu+vOD8Dw48KT9+E44rp79DOEXA6Q8rbA7jG6aPLD5HhgvjsW
gaxPUFVYRPf0+yq+i1H11E99Sw4O1uy1wAQwLl7o/xFTOXEhEUDshIheuiiqOt7o79ufXT2Kp+5q
WGW+Y2D0TWNIFNk5OS2jXrEqndG+7FTuMYbUVcZ9OuV9DU/CIjb3u6EWwaon+ZBIdZx1dCBM1IUj
QLg6Se1sRT8bIGFnBpgQksxd2o9WHNmu+uDtm2J7DUD3XVFdSv2ofxDSR+jQZT/aIaoAvs21ry7G
4RPw4S2eME2jiFlIDB5jD0t4cAJWyLMHeoXArDhcHhVZ5NoomDmU7UDucQfbxytMB1HNX2XUIQWe
fQ0EV4kLWlLhv6LcdkN54Y4yJoI81i6V9jMOgiNLDpTlmU0enF4ubJDURYT+VNLTNXuq1Mj5IkpN
99ugjK2RkgykLSTpCV7JL1AdP5N6lVoorPLlu1VQiH06Caxdoj84OxzkeLbwOAqn/yqkFq4eV3QS
kGV/TaFBwk4xmXdYXLm5suctHyRQ8V6JhiBHXiYFRGBg/kpDplDD7qgG1QTZ1lvA7l993o/U5UwL
5VTVfnFZGLvnFGVzlqgTT3lTtifPFTrH+yqv/xOtiqm5WVZEhvBFL/tFdrwAbHdDOLWykZQp9iRB
NeYT1IwBpxw3CBBF9blrHxSNqdSrceU2FLkRUcCHLWajvKgr0aKphi9v2fl/nqjAbp7ug2FQUChG
QiYPiDqUQtgplxB4anbwPnLkheuUTfHQunEHUlcA9evUwlnZ5y8lh8AsrYZzAC2LMTqzZYTyBDa7
uDPAcoyA1wUwYdhLWj4YroIGRZnMaQYJD643iQDZFFRlp2PUf2EW8AEcHP8MCCOzbWPm77JGhvRv
w9Aw7NVRvwX7lRKrP479/zVVhFh0UnGUNQ8jHg8dPxTUjibmTIyRB88GnXMGLasAQQHHT1r3F+a6
54dBFrffeLM8KzEranUwtzQGliSXXah+ILZomalk/k8onRAkjxXaFpSMKrVH1sGWu2CtFMA5/t9/
oXMSJjEwILNkQv/3Rh5OuYWirOrGRyB1PeYt7SD7yhKNh7YCLYdQ0svRQ2bJ1pagdxsyRj3Rzwoy
Fd+i6jtBZ5PHEfO1C1VxVDTU0b6xcX+ER12WsRIJDXWRpuRsYb09KJBjcOzEyU/54G66xPFf6ToI
dtA5DLxe3PQuFrWF6eoX/Nj5YAh/2uVaPaUUf5Dg5tBbXdiWjQge8kiYjoa7sBoAI8ld/xTSd612
1Gvhb4IFmnuUFxZ0Kt/Uimz/rbCo2GqEwCrwKYhGEKXLtGkhc8mR6T2UafgGZgMASMiReaJHfgej
vL6pQJm3fYHbiu9Ab/Wa5uNvgJD+u48gRA8v7PseN+8JmzpavBf9uCQHNQ/TDceE9UikFtG82r0k
1sE72xx5J2SF5ocUp59tjc491YyDonoQIjogSQs+VpHStGL8vq1hMGjxRDeVBFjJkW86JwTml50z
xBv1Ffbngq7QiLS+EZKyUBhYCqKpUbq7vR1/afP5dz/AwGP6kUbdtf58LpSA9eSkwl8QVWSNS27v
6UxC680QQyZesXSEBMZfrLMtbVMNezsh9UnRjCeu2o49TOPhYj0wJpcDYWAaafdfIjxI5Ot2AYSY
rl2E4uIfyoUyN+Lgk7ZzD9xJOWb58oyKCYK0OAUnFzqJu7Ht1wpQJG4W9yIRjLJ9r8QGPwyRnZPs
PVdghtXwDbs8iEiR8CIcua73R5y+RoxK9WVFP2dYItvWas2hwGIX6Kvhez6URadc8g0UA4uvSsyB
VW4ot7TasUgaxP34NKF31XtVDf8WLVOb7+Akt3utdSs2Larh1fYEB1KrSCX0nf2blR6wuDJYdU0h
O5c/EP1pLPb1jtRmkPWBEcjSxFKaRX2LT7wKJeHw6kDZSDIIeB9RF/55o4mhSMhBzofHABg9j9Yl
88xnWQuTANS6Za4mNdfOUl6z94Bnq5Z946PnQf38xIcwF7vXWfMK9zfrTPe4rvn3BjOBWpQCYBcH
0sEMtrW7OQGBAeH7OTriNKKa+tQm0haZxD8r2P/6o9DTxT+EA9o3eSpgyssGPJezMD1PUHyU15D2
HfARHkbC2+ykyb3FqWAXCe16ZETFh110DsqQHBuLPHy8MR7rgGt1cTeCmEW4nEzNH1t1VO2NzwLj
9R2H9UJ8uUQ/pt/fCfJ0AlRnFB+gXQG3gAvuVk/6QRmfUdnt2zLKLq8eoSvkfLHezmqWj0L7+dBd
embfEWoLdfZUxDKABm4AK5obP0LTjj+QB7GeGHrzAq4Y2SZhWwUABv+ZR9iYLrg7iCMgSp0/Ncob
+N0X18I19upDMq1i+zqux8YSa6okwSSP6WAwcyOZSroBs1XUKoreC8peM3wAYQ8YEOwYdq34BcKR
pjuktzoPMop5Y7S8eJ+PubQdc9XHR33lgX4bcaotgr2DzXYkZ6JZC0pBV0+7lKJKvSZpcdyDOgEH
iWFqaodcplpj5l0Kb1LSxiuNZGwqk/xWoDE7vg0IrX79m6XPjqXGb6MyAyAM/HHolGrY/UpmskG0
nJ15HR72nnpHJVg06OlclYRKDeMvAVqNAt67uhwQOvr06O/ozWfcNTIi9Xoz5GwTPfPgrpbaNtih
LoV8cHuC8EPBPgGfuwm/TmPJYhT1P4VR4sYmPzj3D1Mgk/NkP+9QPpcwoKXZuzCrV0xPrjawVgLe
bvogfhkCXVoP3vcJ7i+lLedtmTW/r9mHkRV8rE7IwsbOZWnEIx6t5b+5OtpnB710xLxxet+kZgi0
clIptNHvG9Rg8gbKfH43RyIjmsWehfCWzv92BDYAYp0e3B74JJPpk15G227P1W6AUPW1iEsJ+jgA
s9CPMXr/rEBVVijpewHBDoMTPdYDW7VRhkzs7uVEK1F/fzd0kDt/KGircRdYuzKMhNhvGwfBAcD3
hUP9UrwD2/zIIYkvn2qVaH2jHw7ctsLm9YslYsSmDukOWyFO50XM6DxMdVse3oKCWpgR6dcZgcg0
zO2DCBb4S+rHJm6aw/63sh+D15dOuPgq3Ej/KIgYuwcl5muVwCDEpQ+PeIHZ9N/MQhPDUbYPr9TH
PmrUfOgcS3T9I2ttLBnPaOWAqiy1v4sIeeTqpoU2fv+TjVjeGLX/f5pfQ93/4gADlINSY0tjMHXu
slioK4xVWyNux2/McdMeYQ4oAr4q6DvppUxcFbWgkDzMHO6VvlJlRJDRPb/F2x81wP3oGdkO86lu
WnEKs9ACGPXY6YPBIjJCWePYVJGPB1tn9tAlMwk2DrgGrEdm32T1pvo1x+iEckmEnvSGLZLR3Xnv
II58Z7X8CEIiEFXBTxNoUP/2y5XlDbwJiyBGDL2VenA54877JJkXX+pXQwWl8aXYaOFTImEEgyr2
90EPfL3OjiOSQH4MuC1kmsRvLijapS0SLCZNm1TsXEbwhS8GXkmyKJpOZwbFtuqgCaQitm35QbL5
Z4FO6GejHrPnLhdFl1h1uK7u/BLVyUWeFIYfe1dTMAKqsrA0q28frOBo8bxjtyG7eIr++LOOiQvF
45UtVQby1+Arvksill1n8PAFGbBJlcc3bRrxWJvBreYIc3mXIkSfEpy9W8G12BeAZEVddHI5513X
ww33xfMb68cW4VyJRl/nC82BT9qKn+JfiTl+EL27k+vR3DkGjjAqHYAugT9W37zHS8xPmzmZ+l0T
DB7cDgk8109zfPncKii6rWmZM6PmMRX5/nPmTXmzkBD+YFioQ1lDrhZswAughhgZ474BSdnmEUYs
QtbUdV0djPb6v1Xs5IjTRIni/pV/GdjyEDrykCi/c62E2aymcYaMKvFRFqtBSLzSH39iEC7pUxbF
9HjCt7keumLd+Iq/ky7/5+/HUdqniMtG/vCXC5XAiG88B+9dtHUn4GhikiyA8hAxjJUjW4P2nXOz
bxvHpq0/mHrCFTXAPRnrUVGubg9F/ti8B0vV9AeJz/dYqW1RQZjIJ3XSIVpJSzWII4O5Q3vtCaJh
Ly58aISw7Odzg77B18ECVQoJ5dGZxvUvfYmDM57pfI4Yuqsftqa4clx4jEu+l9OU1f17kWXVGhOo
kPQIFckNkZNt0uiAYazKvWDWHe6VRNPXTMAduu5L/TBFpFm4RwB4ew36ivNjdwS5mbJ8hV5M4jNE
ATXcHHflbouBH+82V1hh98BTmy7MORmrkBNzgac5a3bMicjhP4ZfiiuYhX+bU3YOD2hgYHbei0V9
2XqgwmQnVV4J/l6U2OYHiivepUVez2kmhCmyWkvicqhxg2UG5cypJCehzpJZBUzIFiA6RDVuHB7L
Do94KrS08EQnvVD4bkClW2MGFm1YZlOjVfxrTsnaGpO9Lt2Cm/TaajSSRO4u/XSs3l6GF0li15Es
gsbO6u3HsQHcM77U9xtacIK5unHqvJ2wg9o23pZA+8OMoR+TFihVvb8BYqijcwtXYzkUK/ek6UG4
HbNKZCpPdiJy+ZI9i9fPPCqLaR18dlp3kLNtaQmiiOB2cMNZ19W1pa7T0yF8B/G3mYpda0D96EhY
L9VSey+/NQWAEG4I3XnqceLHyOe1Ira/yJV8esd7m4qT1LYKphB9Q9FLtZPbty68CSAETJT0EOEy
+d/jeo0ugI0KQTD7BrYYJJ29Itx1T7dVEdZ+sYsdx80RVW4HoV9R0+9guHA1e7SEZHcWMAm2m96F
WJGKllm8bKLHXTkiSLpU/Hgtcj+OS+nz6LvqCilPMosL0QhL/Q7Pbr6Ulwyf5ehrpA29ZVnxSM26
BayYe6n8RQx+iWRW+Uu8ajsIuYnKXsXVJ+1VZB6fQ6F/fFZDz0nxYK/0Nw8hH2pLYssKUj3av4xX
GcgYDD7gwKI6yDMEUZt17soggEo2uEeoQfJah2f+L99fxUYbfDB9u0VuaUFPsjZXRovoWwewTU8T
+WXs4ed3CmUmY8cNYUw9kD1VqWh6FqgdqnnJpPXhKUNrvRtIJYg1jMELCUK7Gg1I6MdBXDqP97sQ
/GvuC4F3tizu6xn66Vjvbcc8SaFx/4KNrTpzi3L+z14AG4u0LYDLm+UNvNaXOV/jj0Nk8BnbycSE
saaWr8GOvmf+IEieQ6woXpsbJuHnM8Xtj+9dtdLWwm6dsk8q9Gg8GfIdlzSKZBxITp6ykSaZURGT
VOr/QwFEuxxSz7NlMwMI9oYaTDlJYl5VNC3YOJ1XWHw7/+FrNwclkvbIh7tPZDle/Cea287UD/Bq
OiasC4K8eMdESS8TQ7SGcohfAYyBDJ6zulHTwuE5lWJPlKTrv3t/rbv1e3RuqAiIa7DjVjx551mG
idq6Wl8l8Z3au5ovkj4dm2vpCoxu/FqL54ynqq+yuFcIdxBhlAsH3zMSA7UrnX08cExLT6lpA4uZ
SKOaPKOKmaBkfWP3XvwOjEDUNjttKgdKIKapHMM+Ez/tZMmDxphYA8kKXEDN7ddOQyB6gUfR5+QJ
yl0vUtGb1zPkXgNM8EbsYPPTUtbwB4RCEO0lT/jPVZtWuqNa21wYTy5F0Vim9IylgbQiIotHM/xy
3CvZoesthiQnmOKZfkdmxfxRe/cf5sW2Oyeeor9B+OGCq4puHWFd8MeJ6BHJ2Be3NpLd3gZujN72
qdUDs+2Oq8HVkaLYHdUE2NJEYNM2z2zEMvi+Dnxrh3eNOO1JecQrY1nKBQ4ybPodl0JH5xaS8Tpm
46xLTMsZ6pllGf0TA09LmDo63D5K1xOZKlCMUP2cD1mJ2CoGzhWGE5mvHFWSBKxLQe/Kx//VvmML
KeZ8AMQJP4xh7QjhliJ9KzGFoNpSm7T5qFMCWYUhMKZ853ZOThXtXh4Xn0w4sF69BmWeg6BlrGba
lUx3Mdg6eLomloKgDhywe54XRmSrs1yruITsVpt/j0mU0ZqVkKewWfuEzEMvRMjXy0UZ/oSEgzhp
DkQzdcSPh9TPNZjrGEckOwn5F0gfoRqRX75Wwo+mgRyVksNHTmKwbwBioOPnTVH94hFpn4JjGpaf
cm2i0fJwDnzaFUMC0xGJPSw1thznPkohraPT8n7XBMpyOMejbNZ1QWGde9y/cx8WVdHfICnysmZ6
aq9OKHh+0571U2Luq3AnuvPwMq83CLoHjFkEsZ7h3mTCP2AnGV2AV1xmCtGYMgOLJXibRG7PYMmG
MBiw4tK9vlh2iskI2DXfQaAb9Xe2wULGBQPDSsUbotJa0VDrfIZTc4Kipp9HDQrjaZmt7ViUNqzh
2OeRd0CLl0ZZQHQw/PE8LyHlp2PdgerYulpZET+8/3QM4rGTIU/OrGB1sVoTmudtbByNicUO5hB3
lU6ViEDNH4bb0Zn9u7cU3VDkzf0hBONvIi+JMEA74q4E0PswDVuiVkypQbkWbGjJsx3Wr+DZ0p8T
ANa4gyhYPUhm0Kzd09kNYBCj7VNGRSEQj28rUZyglFyFUSan5bZoKaqHn52BHd+MBR3gAqynxYeC
5dUswDQTGibZxv1zQSHuwwIGOKeTbXK344lNVq3zhH5/nIvlDrW252eokMajGYGBAXUrYWwOBAQh
Zla5oz9osSj49MwI7gPhpeJfSor+N9xC/u3ymdVlhzjkD86ilAH1jttYWsqfkIPpzR6oU62tnN0e
eCVDiL+SAlQHMzL/GAsjMyLRsv/KhyMsaBBwjif0Sljp83vazyzHngmlWD2IN8IaT6YdzOkxMEHE
iF/4n2kDvnlpWF8nR1XQtGMOW9gmJV+8c0tJvmEruY/54HTnm2fdZOvDt1faNJlb5nGmxGatygLF
M029j/CLPqd22TUkkttUTYlkNKUyWekyU0TlTvm64O4oRojt2050kHY3d5jAdcRTMdxCbTW6Jq+8
Uz9glXZfT0rEv+wwv2ki1BxFbs2yDV67T9Muee37pvn7F5GG7A/kvX7oiYajEsiYHT2ddMYHyju2
BuMROTfY3y5aw5NXQQ2RrnmOppRPAqBXDTaJCtz2Zlcxv0BgzXNc2iR/A7D4Mu3BrMlW8sP90K6v
fl6ihrTEYzHStUIs1H9goa4ikqLQiYjk/V3RC1MgwrrgyAi8VlvEhcGNgVmeb7GFxMYOxHwegeb7
jmrjDyI0DhmZI72xpn520si9wP/+dJqPsm5p9rtw0NJ86H3DKrws2A91HSvyMRP2hQYx111LAkaV
6vB7ob2m+qKkcgDl3tQcBFW0fo5/wBVpKCGQAYEHf90UxPIWZJeweYqGLMG5atnEgtVyiUKG9cIt
C3uNiz2mxpFsvcb1gKR2diX0dtVn26lnF/vfNukvyIY67pw8wUf7crvepzcO1lr83u3MCec4Zwg5
FlVQtUtrebDj1XMYz2fUAh7t4tkxh4GyBAGTg0DBhFcZ62tSYCRPxJ0DW11bfJ6dfaDk9o3JBRoC
uvuAmKeFGq4SkkYTjfYnpabhefUX87L9u8mmhpy8siegtCQI2Nvmoyv0bvSK2psmOMRz1ByVqv/J
3JZ+QzMUvoG3q8sdNVKD4zZbdsG5bPrM5lUwV60AXJmt4iVNSTmC6PWpjbkSYRxaxyPIz1x3OkC1
wT2fUtKwX55OcdZS5joOm7qGDT6p+Is3sDlziLGo+R+KY/tBisP2v1QRVSNRwvrzUJVfGQ14b70Y
Q9X5+UIAGMTM7WXRD4X1+jave6+Xs077ivrOpwiniV6h/q0iQlpF6SVsP24ObPsJ2tStXzfqufdO
yTfngUTVHIMmzgCgiPD2fzvWV5gKq0zOnHc59TfU6pVarhHYBJKHK7ChoI0gSZDUBUayxHiQb9Pi
XjjrSpOSJfIp/aNu+ElNbA5ReXr9sh3eT3TUjyyb9LehQRQrzWRWuT414prU+6z2PhhN69/HFa0h
mEK8xR6TaTi9UKNx0+Euu+cyPSf9cUX6bIro6CjUkshY2SGVsoZulenoOPf+8lwn6Gn+mHjBKaIO
CuoGENhGi44VJ28aOpcNuRu6QdnHewnX5jUGKWFjIIa6os3XgaYHOeGbZgSrvaUygNbo74BWnj0l
0ditZLraAy87ispzrjh4z2JsektPnpuK2BGn1P5lVwbqsOc2CkNuIZqC2XeYCsj70yYaJG+9daO3
5mRdk6D5e0htbyPFZeNoJ4pg2VayH+YbnqgLcCR5v5sdGdlQDDom2RHK4TexEVBUJuNTmle/f+vC
JiqRFX6hUWmlP2tm9Jnk5jNxCKgMKxM3YMTMGjFegsWdePMJNdtzLyVk6NcBfawy01RzJEVZfUjx
J2tjMtpws9tPa0gBkGdv5g0mVGw/47sqlCPFvzrU6YKKN08iz+nfHdi5FHj0KyF1EaH8ZM+WX//q
w9+e+Ko6/SXUJrj2d/lFXqyNcSzJgtT7uiZvkD6ytW22ipmm/W69OauIBMQhCPjeXZ54fC+jN7Ru
2PpGbpgOrYLjM5f9fAruVdhLr/I3LJS/3UmJMZTFDRDMf31jGUqqXj9spTR3aRQfwT9kofQB7dfB
GdOfzBUPmPqbICVlyCqfMCRIkqmg9L6CvsF+sjjHU9Js/nwuO0nfUiFHoKWgj6IdjM/UIC2veZAi
s2yhVxnwbS5WJLXtkZwHvlKpjq0Kyu8P6Rh9jd36BCc353PnsLLkH76daq3/shzrg1/JYcWkRXLw
EO7gAC82Hevd20yK9o1A0ajtSbOZEKhALYquy18FFv3st2WDYbcGKy8ya8Tvl+Y0h0TGAHMgoq4D
ZnMGYax33LN3tMsPg5cFIKxfRcmvNU/0T/knN2Iwq8jPR0oQDb4n+n8Fy8Q77MiX5SN4hgOISGOz
xk0jSt/Vw+WRLk5sQx3DNR6k3nehSLmnyAuKa5sBJVYCfVgVt3CqcJ4GSZnOhAyqwMtKn4wO196r
8rQ0Ke52tciBZX2heepXJLPEqSp3h/EtWPw+yQpPsuhFsE89sN/jR4ZQyMXHO6a4NWpHo+quGYZ5
8vx9fRI1ggQFu3ED9Y0rnM/aKmuJ0RE2db/dHkOjsRL8fTL8RyjJwoHKtYrVTXkBtw3bLpiZVqfy
IifzpmO0ZfR/WYjdTXpCNgHncTieYMNHZynllDAuIhO10woZYX/XXu0pn+I/i9gqvpG7f56aNlwe
qGj4Hx8BbF8Vybkny1TLrbMd1ZnErbm5coM5fFh0WOP52JxGWdokkfzAy5M4Hphayhqy77i8ACBa
qy06/jLCHVRuv8nZuQM4yUltbYF8mi5xRKmLZVC6AkRd1mRTFfWkiTYz5WptwQ6pIbO5c8iranFu
rvzPO+t9s5dMHeV27toJGMrdbnxa4pRYdFoCa00xwP/D/WPdrvr+jp9qefV1Xa9knLTF2gO+DP8q
gl3AHLci8ynUhpBKr8VNEzp2iasRCVm6njyZk+VDsE90Xt+JAAiQFVwWCteydO7XqbVT8PXw4hZP
4SCh6/qX2VsUrrXRO+wVkUOiFyJ9b5R21ZAuyuEU+OpYHA3jaTkW/lMh1xa/niB2s1jwxJXn1uGp
Iw7UD2ZsEomcDhoI3JnroDvJgEesEFLVoIXwwpbE4AupNbScMI/7KZsmnp3GUQWZg9btC41p3Pa7
c000c6J34EJbiT7tclnQm17ms5zg3gJhZmKEZ58TFW8d0JqPWCCCV9CGUYuv0VCnRzlMdWgiL2W5
rtOTJ5FcMI4G2857VD5Sr8agc2VlBINxusUQIRk9cuq4Xz/ODo2F9RE3HA2uIDpven+li0DMoYUb
y7D4tVKNJ5LTA87kgSNtB/5UR81yMP65X9tV5krVN87ChKA4TGsEXfAypHaYAD4JdhdC4Ko6/YOl
9vty58Y6dHFEWwbdF5NW6S21B46IVBi1U20vgvUJ/iPs4CRTWsivIxhWzNyykzFihO7qGham1Zi1
uE3FsH02yWEEInJjHdZUBnyrq4l9CP+4iH/DMnj9noyeqMX7OTioYqC9SXKVik+AmuEPFurvqxKj
UeusEIVmn1EwR/Ml3FB+kM96W6moc3imZYzvdA2494L1Y/qBAqx8tKB+dFyeniA6f5AsxSca9gYE
HXKaUQ5N4120RQvez7Tbh92mMntbj3NVZQReGfCeE85O0tdnyKe69G/ftmvgvCaRVYNx58CUEI4X
gEPNC63HWK342VP+y7e8PFCuKR6YAsPxpiu8EPcCdOFpnsl9KO4LMnSLde27Hqi+l4Lu2Emc5bD0
KZnsPi+icGSF3/VjodJKJF0NjctwEliguPfB21c+WMrMKgHNuFAYpU8Sve7k7KNS1c5LpqWOEiUg
3Q1wUPr++lcGUOC2WSk2ZPbJdaLLW2ZUmkb/cWl++oxuTAOgBCqPBKO5mE9JjvL/YtIxItC+PmM9
wFhMJ3DaFt/KGPqdBScUn4fluK41Q0CWXWnBUOcX7Dbiy8LcsCgYYMAQi/Ftb4HKUXOhWa8Ddnym
LFYPBRY8wMpBlkBLlj/Slq7nFPrmL2SR6aN72V90PqYaap4IXM3YbnsKjjqxgFX6ZXdwBhQmHk5D
oRLZOkGklXF1hEILkB7eB1FN+c69ddqa80UADZX9FZQLu8O4hI9cLSkw9odhIP+/GP55PFzAx7IB
r1g877iHS+b7yGkWKOr0eRVOGdcWi+vw8IhOo2YZcKBMdFZe3XsY61iPphRgZ7m05thAxDl0zIJ2
tcaeRZ+PzJqw8UyALEEWVvFS8RMHNJSg8QmG+yFi7l3+TmvseXTC+1sGIqw6WHsnGojqnnf3qxsJ
4yHC+x1OGgnmnUZ/o9OUGw01qRMmfJUBtCSVeNB9NFRPADla2y70kbCplK9FdAKlKq5NxPG5p1+W
ueDR+MIwSbym102tiCGj7/c/oRUPyAXIREuMnt0sSZSLnjE83RrH9LcwYOQ+mECpRl0YW4wFbUuu
GN3RWu+75OLKQRSCYCt+faHJ0qUcdquIhE9Y6CX+5tidISYflNqYn6rTIeUO2S23Q52dwjW56wqO
udobK1sk9cwLAaYOT1lL4o/rnOKC8AvCamgAKEYKBzViNw91gCAZP8n/t1CLrQ1WGEq8Uh/dkxnx
lcLHrUEuD6oRKSFuaR4kcJP3LV0Jg2LqeVtxHYeqgpjtWM+ys9ZqekDvGWFyHUosjKrQk8irxSSq
LsdE5TglHA6G93ymFrqoN6vuOYmggOQ+8KG5gxzevyrfkyc+jpUze0e2gNx4awb66M4nnzp9/EKE
0RA95+ldrxczPnSbXOgB86LM9Zu0CMr/o7lyxx8+4i971r/CnI5Azlx+rwgkgRYWii90NDu3sYVv
GZx+MxTtIPvlAycxw+3p00fhHKplDHbaFuzPEUjBWFE0L4TVo08vNfeuM0m3QaxmUoEQ5Yl2nYqJ
ohSOku9NkW4ctkHs0L/36pkc4/W0MUBBzZpE7LEo2gduoXlzJoDO4U8L0wKeMREoKY0wqFetm1L7
SI1Wt5V9iT/3Aj45uSkP8wC7KZS6/N1EFjhO/KsTGQLTMVIuyfLFQlwg4CAhs4r9k7FC47/jYQBz
YQhDWbFpzS2KJJNqvbQrGJOxLVNamJDArEkwScu96Q4zay/fsRigsAkzwAJbbVMddop7UHm0Ya7E
lTONeGNrAzvQNdfgjpfam2+2Em5nc0N9kUy0VQJfi0eZIuRS5lBWU9tKGQX43nMSEjnlruxGkKkN
wsYGesqxLjDRVGVpw7sh87rjoqcyh5wjwtPRgDNFC6ckt3JxY2BFst3/D7vcunVXxoY25D52EZK/
itr9YfmauxvsOf5jAcU0JxF+fOQxWR0oMQn2fJuAAkq21sAzEtQ3hpLFfWRkse7/QBgV4S4Vwr11
N/6hG3SFZFRWO1mhRaeTN0omqFvXFXVXQZYmn47BdkrM2cdNgGCsRy1sdfG3mcVXN0ozZ4ml1F5L
40kwH04AAqBPXn7dSjVWRYJXZveOavtDB80fWlE9kRFWrUrT9O8hFC/5QpTqDkBBGE+7rZPS0kQt
2ekgK7TIIIaie78Swks5/yXQdymlV+/Wvl/4OKtsUPUkzuVMZ+55oEvzIGvJYd7aX8mfB0eVT1H7
Blu7FpTtLiRdmCq19LhQBCcKD4drYHOfTLc2S7RmXQ/ChsnvK0qHL4Ckc+VOBLpMTBHNosCi4qYx
y99Ix80/4iR7jHySA/lF7PehyO23fe5l+O3zCf9vRldAIJz40RAV1b6yFmOKVCMXEUSUKt5RP8VQ
wTj4dzylclpGEvjqPxGIT2aN9CG+dHLac5pz4MfFIB0s0WRob6l5qkYRGlfM2y7S3DAkdbhvbq3e
XC6C7wIcXiwnAV8KWimDRLpdmfn2xSX4SxQHadftpBVIEyCE+mwt6mW2d4fW7F7G1FS8ZwIOu6OF
iCYJaath1ftJDKzKAN1Tvg7f4Rpi7/+qOzOdB6Lh/EdxIwvIe2YiXJlC9KBDYi/2x+3h0JB1///D
V+uw43pCmQC+kmOfskTkM7cv3cPf41IqJTbAYiQadcooUEXigUz7oRHwJU2UmiSWm+T0p83VXsK9
WziKGZq0c4jmTZlLwatSFZ9P9dTOilZsXoKcDygYD2sPu45lteK2fgpSooFR0u4OBNP0rfNkXJ7U
g8rJfdKT3C65ekbTOAhEIBaUdD81bo3t06E/ZGRGAfiu1S1JR9xvAG1PHYTxs22rnI1Dg6G7Ki9H
hMCSQVJxAZrSvRcOVdPSRjy4BMBnnYMzxIjrjxt+aeOuMofEh0rJfHAneR7kaAXCnU0csVzo/1Yr
oqfbqLUxWZWJ44gUreld4syp2h0Nss7UkD1RX34lngqq9RIOntefPy8rH08Te+64LAM0bbOQmZyQ
K1J1OvtKjyJ8Kn/Q4C7iN9/yB/cySwBcr5AeJpWuxk1DFZOZ5I1I0AsMzGnCjMHiFmi4amHRIMrB
kRS0W48lTqZrfXDecOmPJ4qJWGiWy5LDr39aM8vuNyZlDKv7Fe9KpTwZClkKXvTa+OWoHN8HHvO5
+Ck7W8upJfiRvpe4xgMA2FzK0OL9wnD4AsUzUYd6JCtMs+IL/eQKT7O9iygohjksIzWUdqGKEC6d
Js7lqf4yPcyTBJtiyWVZ3J2VF3nof9uGEX/nKuvzH3baO365R0AY263qCKsp+2hn+OqtGWpB0FAW
OtKR6IMBcCb+LIGpbYN2ux39TUtkwnMM47S7PRIoI7hbXPMFnuK0JMAjrLj70pgCs9UVMd0e4H9C
IsO6adV+spuZ9IT/yMpkhsMfUyS9m0RC+cXIZLOJYxe04vyVz/usdRbo3LXFgMb9WHJ75s7ZmaOG
15hyN1zF2tT05Ff7je5zRAWGUJFnI2sOyKrZO02a2Srr4vjfgdg1MWFPpetwxhzU+vzS6f1fmsYC
iDW3oLcAcWTTqHEQ+O6hZfHV5NnGDcluKmYXYZb8VcHqd49PhSVw6/j+V1iCUc4McoYa5cUZTThh
/TV9xvkxJmJPHhQ8JOJPFdFXz9FpKz9WTmiSgrxN0Pt7/kLJF5B7/8KlRkOXZBzV7qDDHPNVvXJ/
Z3eoejNWa2sXICBivTr5dPacIkYl8K5Z+3MhyZu/dTbq/u2+6Qa02qcpCQy2jRdPbPZvvwZv9sec
o720SVZQX1s8mrbBJjltAFu+ThYG8ExI6POjpZVSVPIHuqlD8r/sEeAHhdnmmuYuPzE+tIzXooIG
knW2KfwwT3GpV3KpvtLIYCOfYosAKEn/Ac+k7gtryvd2zLbMPJbYdgVPTBHGwJ6pgMxd37hpho7Q
FYb/XS/ABD45HYElFuNzgz7Ukg19atpKosttE575rxLpRZY4wM/9O8J9Rh4f/7Ri9TJeQ3WLUKoD
7JDQYENsTU/bF60SflDX/fobHPDyFf4Fo3InOyw8xt2n5zgM5YuwOSb1UqX/6IyRk+anBSBsR18c
z4O/HagSaI860Mcp8yh/bMbi3AqcoWNC4C1fw9iGjCWfcYimVJS1J5TTwfZKOJOTgpjXGPUCM4K1
VCmiw8uKOIYWAFOw7UPZeehjtymOUOG2m8BM6tN+neR7ZwB7V6kY5C2wHoOIZWhn5rwSib/OkGDE
CGPwP153/VEFEDXkMbqAQlliPRAOWAf8YUkhASfLKtXXMD978MZSO5+SftCoqF0wSzuhJp125qTA
uAspcrcl6PUOpOLdVQ+oLRXAayHg8AjDKfx98BQ8ZqcYkv0EGBFV58LPJJi05W4WDjTPKq2eDZsy
dc/S6+g2rGH40KInZ1MidFr7KRAHwLV5BqpU3kHH6TT7x9Q1hPyhzR4wD73jmc/D0KHXgLu+5igh
Bcze7aG1E/l9kg8jsWmZ/Rvl2sTRAoHq4+fpqOE8xHw4lrekYOr5De0EmtyA91PbexLfDxfLYDQ/
0lMDsRKF/XNDdofuvkt5dWlkEecrQvaDMm6uL0jcAxWLnNuiWEijgVi2DvqWAn4EPAJrKLaj+cDU
zxfTOL0S8ZbdAwU3YWTdQosyCZjjwpA+tuv6WRthdG9b3p7+waAl6tcxK2SpTUx20fxj5eWplxaI
Cghg2ilsNLQ/NH4FpdPPS4bbGUOWdU4ory7LvVL6sQonjJufjxM6g+Ep1s+2TBOLgLxaw4nS1+QF
TI/NHBNnPL/L8UVvyXWJasN9HWyMRNy4AQixM5QSSi974/ULi3ueHwELkItyV/wLPLs80m+0YYNe
oLJEUd6ZwrTiH3clR8wIAHIDhDM0sEn6yaU69AOsiXA0aSWrVe6k3vRFQUdiwPnmAKghoiCqXguN
sgnHTbItPxsSZjhDsAFJFUSmchBkoJmBpeb/v//1H31+x9+6VHVd6y4ki55n5GSeEvTU3s53mGoU
0Q/IFNaZx9pxNNDie9gWqiepnzMrtF4FFhuCjEaRE3EwOqNcfBEbpkYXJbQUL/obcggTNGERsuP/
UnV4gPZmwslbazFSVCFdasP/1bt5iu1oHCVMjqDNKCa13r9pP/QhgtQjHnNPLtw77mxnn9VXhEsk
K+cCp56Pgk6+yAnuyIqwk9nslr7XYBYBNSYfp0OH61v59d7vthoaBFF5Hy0UJ1WyFaicaEWU8YbA
cXRRvIE3TKn4rVRedroXaAEh0RbP8arYZsbIOPVfX3+bC0Bu4v1tSXZ1u7NgF9l06IfbebSiGSYE
7BHQFlRbNqpV/ehSFSxFqcJwDv+cThPEqIjukfnylphtBLBXZw0sGSouPPxu5m0acWkEg45fOKr0
S/4jbnqCsK84dvKxBiQHhwB6i8bVzC4RZzgxLf0hDWr1MJ2JoDDqjwaioTFDYgtbeFSTd4drM4CX
U4vzqMIK3hy+ZeVaVROV97944MUPa62yVp2QpxdzKLNvEjVScox1r2ahvOfGmFf4zYhRaIotULD6
23ulPS8O70xy60otGcgYY9Z/oO86dENTNwQGqeLL9ubplJL9NhlEnXiZxZXk1huWAL+hy6TGltmJ
soKvkiBCgf3v9vsYDHJxd4kl6puUk/uu9I0sh2rPGke5KE6VNL8JCs2XbErNEHZ8CwjY8F/OPFpf
cDzJCUNvvgMIwuvFO+4pv+pPfMiIHItQv7W3r2Xmf1bxTE7VWpwOL5NkxZYqXzrBy6rddpjXrIqZ
MxUEbLT4F3u5xHKLQxKfTfNyTKahyaggnykpSaLtzCRDDGJFGEooVaFeoUDUo6yuj0LS0NHKYN99
We4TD/yCz+WL0HB1LV4bhWSkU3ypIwXm6YNSW8Gt29hq3u4iHAryGtCvRkf08J0LqHNCDIkkqYUi
tjstsgQgcK/aTHvt3FmsD9e6K32dFs3O+JnBVc+Ez96gYCeiz6SFo3PmkI2pMXyEvgddIrZ1AjjV
/97pkQGG0uT7CLb9cpECUuUORDOQJHdJrky8fYqYDuat82mr/nT9okc1kzMr4iFQjL4JIhnQNXxJ
sDRPAOmCrhCXZiDt4Ay8g4I6cfJmecbfxJ1Ifn/ZVKRgcD1+1CZLayytQyuW70RSmnJbVVEfWWtJ
Bp1VVSvr4ir2sAfWV4a54OVhQ6dY/sAz4Kr8UJnHA8dXH71nW0rr2f1HW551vRkMG9tLkP2WrOx6
O9a26uYYUEiHWVQ/CPNQHdTXjk60I2lyieIMhJUupjPH4doVrKiPy4AcjowqIX/zfL3KwagQTnEu
cVJKs1ICeHu2TRpNzcDSNhhlvmr44jDrHDWC9gsu782i6aqtsq0PsXzzABpQnbYYVFhPn6g5wj+I
GUGihp0RSe4FblxRyIXEr2hTbf7Aj5NwpJk5Lmf0PA9jhJdq02f57SYbDiMtLjZ6By0JD6q2HRaL
SlU4t5Gv8hYK0EbhVaiP2mOHI0o5+BEhKd1XCdi5R2ITsvMMfhAZjo89rdVJyd4zorLgQhq21YBA
hKzT9n9jGneiTq5VOXqbvUoFKzFzFn9OFhlCMObvbAbdekXE3qqDD45bQ2ZczofRwwzuE+PdQqtf
26DBYCmQXFZT8/pjHrJf7IlCjfnXzAmagoOlZIkVuoV4u1uf5YF57UEpADnrp3l3aTDQZ+ciyR0N
JCNHxA2Q/Lg17KCci9p3VVWQKoSr/Sx+Z46GNwHHosdwHw1e0XIEJ69YNzzfUo2UfWmORusS/x5I
A5GFR4cj7Dk+Ha4tPm7XhuLyrs20qu1qZEaotik8u5NHejzKSKPTlHGA+4iENZauNEeJf6FS2sBr
ybwQeQC6kWcZHoXm/lWpfAQVsQlPmMT5Emx3T9+6LMPWE6P2bjJPrCtLqB4dc3EyHGXv+pRpEF7u
pH3VG3rC7F06/bIeA3sT5/UqBJNfCTzz76v8R7adkPG0iomkt7EWN/vA6EpDQHpvo+EHgqNpGC3R
DTLh7USW5xVdWU4TKPEhzSigTqxB1fR4ueeaCP/aJ0vhaIWo+bb7UHwn+5eJHxNXyAo+UOtcRsOb
QagaDQuzTNcWFgAvNj2yRTnYIQvqdRPWVNUy5KXttu2KJGTyIZZra8MiXlhqTDTc3gE/Dmf0Sj6k
3IAuSUeBl1ca/+HjpYNBllMp3TWBCt5SzAqtDAJc6F6DfSwk6vYHjPZxBOxWTS6JmivQgpwBmGRa
Jct9ceTiHp7rFXgCGWYQe3F1+jHmiq53PCPbfqic0E8cAcFcYUlkyPJw5jUhWAI7oJucN9pfCS2s
Njld+pUF9MP8MvHDdhbb+HpcamHDyx2Wt8sCX6sq7kx+WCMM3AKFVWbEn5S4zXwXnpGK11RXmCns
MXAtwo6lk96Y69PIdcSI5AQ5g5Yda3xnKvSp+RHFV3nOaiENn7KLHoBqoToQQNizn2D06zWHNqjJ
dsWaMyp+cRYXZiaaRZl6EOxgQlEzMOKLeKSlhDsPBhMRy23lz4vWH4Uanc5TODKYKrS/h2heePsN
U0O2z2svZucE6HaNZ3m9p3E5dFGLW/Cf9Q4fDYIKYKgvU0pk0lpSsFsNXd4un5MbABW7539PYM9N
0RE164Hgq0HZ+AWdQIlX9PjAQtlXYKiqvwui+wjd5VqEcBbJ7LFEJmGqqjCPqVh/BAfzR5kFgT8J
rOLpAsbOwIqxHVTEEH1PE3N1SKg93EH4vwJgzejwlF8e3qcmbuKOx+hidlb2oBKdql4Jax8jvvNs
a6FPw4QZBElZ3rtrwVwwzARBYzASJ1aN+fmT+EIMgXk/Z3azFEnNn8t54H8RCNKEj1Zdo+izkUdY
vrEUaRK+IhVcG7Q10+Vo1P5BGVdQs9nrzrluYOL6XWNP4ACz2iM4u1Z8ua7xuL3Mws61pdNNaegI
Kzj67lWJOqVVLGqmqkjcxQu7k2AcM8tdAH2dO5r5j+sacOH01DZLx5zJ2B4JCWbXDMiNyO0J4Usq
1fvpNVGJZppBMOPjtM995l9Uwvvu/ADAsjtDVqH36JfCA0xaVX1MgicKYpbmqSg/gH9jX6uNBtaS
oXRwdNYmnblJeGUrBcDbtFkPE/MsDo11ktArmYPhoxKDdhMWNroVL5Q6m5pj8cyNari/zj901/GZ
uKVHGJbxq/Y+wFSyiqbP/jlGDK2LRmR0p6eS3kjTDMXsV/DWMqwAFaVUHaQlMP6CqsOz2s7SBB7W
2TdwRt9LOpvDku+Kyo1k+FZt+sjBAgoeWNJ/P7KMULTyXAZuQbW0JN9zo8C+O/q1S0Uzbx1UHLg1
ab/PhBujaVNE428Z89fS+Bp0p3XlDt2Pi75W9dsUA/w+KqEw8egovi1auq2zBhS+63Gz3Gvph+7/
LiCTnx6oPSlNhXQR/MCy6dLPVAvdL1RjDfXDOuBuRygN1/GpcPSA7wzJvxZ9dEniYVZvAUICBcPj
sRrzsTpQCCGrDxlr4apl739Xspjc7OtDoMdanXvo2WU9d17lhS0YBoV8yEmwQc3unR+wdZxmys1N
n4/PIkuw/Qmt8a5aI+3jAAl9F26vtaBGnPhXD48T20DDzmu1WbXhFNV8Vg/Z9H1u5p/r7TBFgFvW
wnS8hRgrA8Za7NbcQtcDN80i/cFCae8VO8CbFFjFLgPYNkOqffzpoa6MzxLht7pJKGjdO5LjqAzl
eydTl+AIZ+uWijtcRMplmJvZNIgNIYSfSdvLqAqDOC1lZTMc67gLS9jbWxYTCaQ9kZ15x61PkQYQ
Y31yIvMcKamzkDiIHlMHTW98DfDVhLbpuWaN2XpOdjnPJyhp375XgJvVSTqL5oh5daiLU8wxHttj
fOY7CyI3bwbXhO72M4nkbxHDRNoP746A+ylJkdS0/+K5oEKS8Izwl8S3ONIZSaa4+m8PYYSC5Iwf
xmN5s21tEGoFCkdASKstqB6DMcqjkgz6n1EZoIOvbfEmT+i3koWhdv5I+mWpU9f0wVfZ95k3WHV0
jBVrGqbBsnJ7Ykkm9w3G3YyGM4gmfuEEELc/6Jqd82I5FB2O/f45EbjLiqqFb9MlJzKCXILB3Db+
MapGhySnmYAcfRmn/Y0rs/2MKXkeWT36315q273twYJsw+jT/l4FOJL8RiA0WpK2wfK2QjVkIIDf
7mC6zQp5SUN1RQ1a4N+BlgA38/qxXDVOoXYWbb3yCh+KnTjNLPvGJXYQxsVCPiEa5KFmE2VShuNX
0RHNfSvNN4mqAvzoLJ8Pv+IbisLlrwhvEwSNZFdMxxP8dQgu0XDRjYD0lN/SBHsELNxoafQkBV6W
4xPi2ei9ZMTZIvOxEXAb6/gRbMHS1wEIWdlwGbrGiUbBuXzQ4aNalF81qCTE4oFh0cQPZ35ds5ue
5/k1IoFu5mTuTH71SZW2nKCpi0cGw1L8hwjxrcq+cRK5/P+PusyE43mxAJsIGUZ3jljYqHy3594P
cPLnFhvlj9mybe6fiuU7knp2Al0j1707boIwxe9qDta2LM0Y2jnv6Tl6xJl3UCHCDp3hiHBAkaDQ
1UG2zBaERD4jaKtGUzpqSTg4YRRZ2aFp971c/N3BdUQQAsWVpkZDUsfd+1EZm9ou7SuG0Je8XRuT
AizklS1leDO15Yn/5lX+JISE+e+TyyzLKlH0tPjH52IIArncueEecKqLq1Zj1+kXHsBBdJp7RtpY
jKCG7YjQtPlJozPEpEImknzVfJSZfGwKWCOcszdsihw3h/jCnPP022amKkuTsIL77KTZoZ53kH6s
OefPs/mjvbOAljSxu+QCDfGDM1UczgLYnyMVtJP0EuLnODLnNbrYG+56YJtmwT3WzbGgTaq8N/EL
2tirajmhgur32xcb5FBSTYuf9C+9zkjoFu4ip5p1v5qHfWCAm9sitqSCX+A4ceR8CvpJgby/YdmR
I7JJIQfdXG866iPGGqIDm7M1z7lImZGxKAKvT/4IUJVMTBXE/AMJcVhugz69p8SCX6c4ttTfrKZz
xyxpH5nt0xp5mf+DDcaR80dxozfWYTsKvVm7LsfVAcemVc1jkWFV9wobwbaK6ZfMGIbOmayUTNM2
osNp1XAVAnvzpqufS1nD+jEx3rxT+4F981JNv5p8wEQ54c1sYhW2A2SsUfTVANq37i315ADnrENf
qWkYt/NIPwwErGvJwsxyhXuwemxHc7/HZArNQ0arVyp57S9qbXR+gZhUdwUn4xay2hjRHolJXHrB
7CGsAwLOSO7X74nvSzGJOA4O0xfxiy8LkeR39j5RcWISkrfuuXAro+SH8/Tf3u9yRjA6r8tBxOCn
i1WYGsoa3+9gbwQ97GtXEQ++htDpM1sqEv/no3hKq4pkol6Db7kxy/kzY5/+CupJ17WT0f28S6XY
x5OiFa4npceEVGjk0jhungtFFq8pu5byOPxkNtxDHRDAz0sBY8Sk1cG7nX7U5r0hJ0/PTSiecL/f
Ne/ita98kRZWwY+DeLWJlpPSH8HkUmkB+gWa+I3KmZ9aVExAYAFf5xqsvMWtuC1wwzuv/grp484i
m/tzxHpwcmLA2f+r2qHB120spUpgqjXg8dVMkYZsNEaYyF9fAbBzRS9QDlauY/nldkhAlQ08SAvE
7uxtTjeUDzDv9PC4y7eIubJUL2zjXKUtdo4OVRwvyE/19dL6oeyR18cspvOgq0+h0BUD5xnbbJvZ
cYKXgmM0vj63ety3CgZzWNxoklj+cNuKudeG8lfC3KA33t+YUe+v4/vbYOY06VkDnrxMVFb/8jqE
7wAUJARzFa+zbKOd9kCX8ucHWrrQlaqjrvYpZbKyidlRx7hvIT5V/6t0lOV4qHwzSFrc+n3Yif7x
EMIBU0dPOMXezaPebT+IdPA16GbLIja5+MQNkZwsBi3jCAS5mfzM80Qt+iFOqw3ccnDslNmAASBd
89TJLCGYXIIckQy8NIq7STUHp4PkfyicoCwNKni1mS0M7kPa/4iv3TStVDoWKnDcdUzdnDOj4XB6
F8qVxJQjZJkfSr/EF27bIlycR9fnuBFt383ANnWucWmPqXzE7KnfrfcV0izBg/xrEVO3rVXixGrj
XDA2m+lS2GftqQE/XgcIFkx93WUiG3Pz5qlOs9Y/X2ZdKuyjAsvzZfb+ZywRk/gb94ZHql5fLeHK
pr65vobYZySpHN3Lo1/HEGWMaFrZhPBrcBHlFKGvv7ouSPB16nN4jqIXqvElYg7+lNQ7+rMogz02
OBZuzTx6bB7DiZdQRbLwBc2c0zKH0THTGDrkiqhsp7nD6YU1y15kD9jcf6dU18nlOOTCDOFXpQoo
Qn58mOislMK5YEOzSgR2W0AzIFeTFnrEHiAyr6Q7tits6RDtdQopVpYEebgyDhkkYEdfYXc3yAc3
sTJmgomGKlnxOHLb92TtjX6sXtO36RY6DeqkCCz3KtaGQwYvZh/VgQcKmOat0f592lesNn9rBF0o
ZBjqGGvYT98vkv2JAbmbrprzM68pIp9dhF94I+/w+5URzYclNKJlFxIexHFVnqi9/9rOA4UnTrPl
N830US23yvymHKNB1+RQh582rx5fHaT+KekNNeCTOUeMSgNpSehxW/8eEB4ujeXi8R1OTd8Reirb
xH48ra+zqYQfgQhHRsvoAZlXEFdC7I0+ES5Kzf6dC9WGW5WONKt/N7UizBu9JCvHxrvOr+HNB+rV
K4MNmPFjygB71jQSMz5sPJcttoshgfCQ1nByrC2NYjhr4o3xJr8+c6GrmzMbSaKUR1D+2VQFctgh
mEa6WZSEY5iVPgWIdD7PNxO+UjxJ5xmwD6+zcAa+3huycbXHxDoexDX9EEBj06SSWXiE6aaXXNzx
xUsnm8KAMml+QXW3oeXoqvIk9yNJFutUUAhc5VDf+JkLReoUpUIsGaRMKh+1YEv2uLfJg+2ehrNV
e5hyoWAkXwDFZwY3e+JSDGd19cq0eNakEEe+bdSRQHXPx2hQoePhfzg8naEI8izLDVJ0Xlx0dhNP
6Kqc4T7zr9JwsD6GXw3iSRfN1SPJHGWYA9Y1GCRuZVDfuqNrijcPNRXMNX91ecBL4yJewag9QAzt
ynu/MefEPWE/OLexX9iZjcOrkcpNs8OND7SCn+YlUIwomEhNBLrEQDIG/LTWZC7hZLdleUYA/e29
YttQqxQcaGBoN1DW796pCyGMh9DGose/+T/L/hBGuzaxRMHCIJwhFOvAXB+pqQ6heyTxCvJIL45x
EeNJ6lNVYBHRrIUw7Wn1WRXBpEaocZoui0Lyw1AWs+MUM3PslURLbzpabwxd3XuGLEAlaOXI4nPO
lcCiAOEmKCej823MR7wIQLGWxlnuBxOL00bDL/WX22drZPO3F9mWe1ZVEmXldr1DKNrka35awYpl
Pv+dYV+Pha3n4KzqO1i6f2MIc3RbsDdUcHHkW8YAEVvkOy5OQsPT1UniXMpRwo4euZGknthE+VMh
771N7SnqdiKlBErWGdhKOk1CtvZwQro9UwApRuVfL17JqIMVQZESQzutT2lZ0vDbufORorY+dvar
TQF8zrlOmuf74p3J9w3oTmKO87hCdfOTQYkj9xW/vwC+ygA4bnQhLkAxd+vivTXGNuGrXRw9iH42
52ifjzBzJh81DNSZtqmWqCXNn5USW0XFvzA0ERsqBdS1aMJRcGrUTtS1+I4dzrz5L4ALv9/0DGj8
YiqHttWCAoOXAVJ+y8kKdALp9uE0qyt4fORfTc8RTWHglqQw+7+YAApXM/61Vn6K3MBeXBwD1b31
fCc+1ix82TbbBPujcN/jJjzNxtXZa6iFSbxj/Lk2Jy0NQ/aDxe+B4RhZuW3TWx4nsgFH7VEKEAEx
JlnfnUOLwCVDGz61WmuGu9ETCPs3NyABaBxsac3ea9KkBkewkIBgCZA5Wp4EszUEgzFhB5m7+qDF
0J1xTR5zbOojmAfqQgiwPcqFlxnUrw23N04rD98xOljLQ8pORK+Z/M4uW6aAYP8l/L5d/dPpoSxB
ujNSDljaS+UFp1sMXfewJBiqsJMZVAsEygQgxqI1N/J8V5wXDCsXxL7lmmBsWQuU1f3jTpNW3UG3
zp0rbyHDDpSler7RHTbkdSKVSfhXU8d6vJJZWifCveRqOtKtGGkMk2WjJbhip3M2oEd+njX4MDQA
AwUhaELPqTpvVmNqQfhkFa3UwTyHEq9QB+DPEf7MrPn0F7ZQrFRK1W0v0/A4uR0ZMY16zqhEFpyy
8PI4HJizwAY0IME88VhOeGNJcEW6FD5KYz8BCB9cU+ORKqNJXGePvE7HaH7GrpecU6bH7TJse2WF
nUd2KU8tG0TLfiC6NcjvhsvPoZX3+4vNgvINtHjWK+Pg9yaDzMIsBydZOrp+Y+KBVHkiJo7mE1v/
oPGg82ccUrgGTcS9TseMzxXQfQ4/v3DgMpHj82H1Xwt5V5IQtd6amLFnvNP+5OAPFM2T+rUXJI31
7UM+NeuMTTAuBB2zh/M8z2us6SKan2oMcldXPNGmnOQ4G3yeHrc5QCRGNB6chyiMKcQr1sL4fj0e
nbkHP3izUTKmpc7HNt7Q3FbYes8mCCoxYnNgtc5xEoDAP1nZGOBk1bkbH+blslXGYrB8q82VQnPC
29xp2UgLdSLDHky/B47Wz2JDtP7Sx4Gszq3aKNHKMqYCKUfHrRt3LPC3FzBrtXXJgWDo70qS/vNp
or2lH+brmjThJwh48EbRsqe5gLgmx2nwBhkG54H6Vcvf8q5/YOuVNezMl5tm7chRbjIQJG0l+RA9
UMemD28z+9cn87nBSf4o/uUjSnuRCuP+K5EfD5SrwsJn+568u35namh3czgBrGih6cj/fvdTIaOj
YV4cnttTxe0PQc3a+VhEkwt2mQhHgQ4xjYVbtVmVX0OcivTNpZl3OmgcqivEfRo9GxrsmMUVK6IZ
K/qLRzfT4Mwq8P2GN0nans6zDmnnmP06jbMp+gWb5fCyAXQbr0g/+Dk2rBnYkr4qGa4RzsKURlep
Kvy6SZfIaf/1a5SSx/5gVU8lCqK6bh2eKUI7xyWbhsEikRIJZz7xw+cPoaapvELhIn7zi+XlKW33
ocKqOM9v7FNBJPSyCemFLswNCHLm9wEdiaqHmFATgRiUGCRcuNUfWROyYju4uhvTu8uucRnOdmqg
7Thy9NumbCUUHEK1R9S6Uq7E5WqAaZrEgCIHO3Ti+Xk3TyY7yDJ2QAFZ010iAeQjX8JO284FVGpx
vwt76BhWQ7u2/KOdfR1HgSYxCNzmhuL9YEA+SgbkL8Es1iBW7zt+7Ce9e7jINjdiW+6smfgvlIWC
5zSyJ9mzzCApIVy973RHV5eFz/Jw+ROLGVHsU+a8PT5bqhrBuTO2Ptb8+y3atDf6HAcr/4jhuXQQ
1/2V159jGdD/gsVBYK1QW64P8PAkv+RhUer6ipkKJc3wJKxk+ffQDQeGcJ6UEg2c+GQ3UST3HaJr
4KsNk0DfZkHhcvQVfQWHj19sKPFEmxTMHsa8fThYx8r5613nCqts45AIcLSbtKHgm5vMPNy91GlZ
aqhuKGQCGpqHOvI+BCvp9S7vWWoHfzcVsKToJYgARU+L+ILz9uBLg4eV8Lgp3Tg+3fU6ikh3dH6M
RVNXb6j9kBawVnRM0xWlffOpd53ckVI1Cx+aVw7CIVyqnOAgCglG30Vp3NIdKn1+INYO2ibU3shD
AccdPxC23tR446XKGPW320uzibC0sFBjFfIyMl3YOjOWLKE/PbsbIOONtpdb/lNRPdk1y4s0FIMB
6SmayyTZ+gsr4jdONgtGmohjLQZqjzpvCnmIky2ZQrO4A2jn4eOKqt987RSsiALdbBDU40pWKNrD
t8QqTl3czOUswlg1eLHdabY7LGX5Mamwo6Of3o8A9XelJKAuxlrZhURtP/H2anXtt3mO8GXpjoEZ
bC/IxF+7UExJ1fpQncER1su86kLtj+U7pK7CCqkN21ApoF71Tm2exgOgJk0UtI1KF3mvdFMi963F
pfinhqBZksHQyPpcb4z1RbjO0+n9Kywz2gUC2ziPVWbyQhPa+x9i9rkKes3eMoQuLkJjlZYjDXbN
mi5xTRmCGQVjt7uKYwcfKGj1dNs5smbJo4RjnlSe74mOe3eUMJPuU33C8m5u9nc6N7vif+8YC4R3
bbvGwYyWhVvZFTbztzSvE0mLy0HAtRQbxvTNiq9ZTJDuA/Mej9rH5laCJqBIVogfH/FNJGSutx+7
FKfgj/FRof5ufA0110vVGeekKSAHPJUPaOdrrn0x612Cr73/DkPH12pXVhrXDl036x8/XibZInp3
HJYuneCQJ6TqqNKNod9/YRZwD4UzXsaIAKqogOPAjSWSZyaDWCj7ik8iTqz8A/oS9ehQIdxcpPZj
T3y4tpwJBh1icwg+/y7wocHQqON0pAzJZimHYTWjp8iNe65ej4W1FS3py2tiRfSGxVFk3YS58tRu
Ejp+VVwoyROUar4+mXFm/sUkxRCuz2cf6rM9HxN8SnLaXHrPRQ7EaIVvyhM8MUAB+il/BdmHkFvZ
fAfwPnUl5jSuU9qeO6EYUCEzBdI8RztaW5HFmBk6fV1piYxUQ+LV1wn+uNRP+HaKAL8R3Czvuhf/
mzDEEtSNDXRhBiW9Lo6LLJlhvSLNDFClWGIe86NPIVr04IOjSmQevr/XvgjzdssjRVsMY5HyTvyj
V8kJ8qyBOA9foAIDR3+c8EorCFufFOinYXZuDO++rOS1s8x8y+FHGUsTv45niMFUHczUcXCDizf1
xJ3a610SrA5Tx17uJr+naDW1kmwBSuazuIhmrFiuow0Ch8MroMBOmkHWyaVjpdw9V2SOgNWo0u4e
H9U2M9JfWcM2v7yXQZQKxCmN7+1ormP6sG3N2axNZ/MVmdpz2Iu4prH6eWBRba3EBjXae9H//Lvc
yPeal/jerpgRJhF/Xx+7QsupevVZYtC4FXhSGpA9TaiM2f5kaH4ztgWRO1ONA7kEAffb4fVS45sa
rLzPgMvTUGlOjq6N83LPl6Gigbv5kfU3UyyjJRCm3W7X+n9XCx7SR458txEOb5sygLdMFLtlm/T+
dAMfrZEuIY/OlJfgs6N9VukGDFlOZRAHfKWOiJMnOJTp/R6L2q3xbWGQ9iFdgUuaXOdgStzJ9nsV
fdfqwGZV/KLngYu9JWMCbnA0zliysVGB/+Wl0Km0cbHwH6+2D0vClRoOt6O8kNkrx/I9frPmKPCz
Lw0fcArl3kU1SLOMyBDOTsWcbQ59lJBnrgwDZ5LUPmnPrjUCGD+dVUoEwrBGKLw9gCGR8FMSTVeX
uoxzfYOfnnFqMpDv+5I639ZcXyo0fuHXjXhcLCUTCVkeAGu0ZfJZt4RUPjUlC4ap9D6G2kAQ3qSG
YsIx2s/pDH/ntW1+gMsNzeVV/UPt0B9x0qvHta4AAjyZ/Dm46ZjIVxoP9E6LZhCZzviZVsFAw+Xy
XQ2pxXNSXOXZFGDlDH8PG4jfWAmPD3lq9a/kf8IVQCbGwl02XDIs/YTVLEey/W9rvzHKQUgb69kb
RfZGWfV4zC1TNn89OV5Kjqts8+piZFLFki9S+Lf1R9t2p3AfIKIfbhPFS7WfpM8JbIDDEINclc4v
LxaronrppkYi2fS/syA2fCNw3v/+yKTDTP7mYZt+bv0ii1HxCLOkVwtG05aharPvORISoZySCXJm
93qt7fVnASkauQSEVP5jMU7kBEfCc6SAlkKzkVuY6/acdBm7LXv+MNcMTZziU54HuMb6uS4MAYF2
z+w1dL7u7uoegurkESPtUitCO+tFjARNyrSHIVV66abFt4DvodAy15F189Y9GGapn6tJAqpD3WXl
M7OPGAX3il2P2vgmxOCt4YXSua14lJy7AXrgNsff7lu+51Kg3+b6pjMaLPhjiScVkznIk9CY9eBQ
fSl1lBf3sxTyiRlPoAC8wtvQn7VJ1yKTaPTK1h1ojsjgv50L8TnmvkswJpkTsvHEuo4BLTvRlY1S
XSv1EPYv12mE5gAAmwIggYSjNl3wtEfW4iRFqHFHXX/k1FGyB0EyZnbA233YDFqCKZQd0qu6lDci
LjlY/CM4HsHzJ3j+KsuaDUqrRSdV9FMv91YST8Eo1P9PX+28Wc+QEnCFxRlEB+y6JYEvQaLSo5rr
Kw1VyFdDI8TQ9P0IiyB8nBAlxHEjBk3k0p9CUn1ItvDeSZejG+IeU5cuOcE7BSmfzOojPpaJI0ZO
2QIy4xeiLalym4u1xIRXsiWTjAz7B3I5g2/Bo08iKOGnNGOJr/Niha5cEQA/nmbp2pKfO+OGMIt8
MgPSTOoOwq7j4eSAkynxPUoS/4McXRKV8/n1W7mwGhhw4mDfj+Y9BD8NLTi9cQ/j96Cvw8xgbEHo
HyMta/dqd6TjYL0Lyxm9dEdn+wzyiRCcb5eim4j2QdHEo/MwmvRQjj0CpupuSgrZbb5nipSIruWj
7FU8w0W8dU4POZmh7dseV0DUP0b2VtjZgZurY8YYrejfvyQz7op8UifpsLR5nz/sIDHYIbD55pz7
BixDpb11coylmgy2SveexvmiTIFGZnT9SEGIjyZwT642lKKFxhQ1CjqkOgQhAde9boMUTAAk8DYF
pBvZhpk5mxSm3NIDzD+iDgpebFtHBL0lVgNdHCGTci/FXiBvdvpG/dNvoPx+AMPG6tkb9+TLCdva
m/AqiFs8y0baFGDR1hTlFTb/euhs9EU5ACqdMcGYkLv/p4dCnYOgRH7jvyl9EGR8nQPRacR8u7Qr
LJgCMhxJppZEyFhAvrAyKFiWQCTTNUhhwxiL93+AxVgvwsM5m9WiO9lmZw+svZsbsa2OTr983qIE
lFG0h4j6dSYYq4H2AcoZY0+ozSIuI9mSuN77KWV58Uqzjlq5CtkfXFeu6Juq2WT34xf/qMFB3X2o
tpQjlUjN/tpf0sa4+ohtBxsood3AZU3JqDHKaMYk1Oly3tJf9Jq18DswHXMU8obuAG7mlvOJKEEo
zLNIeE57SJCjmD8CkkNRFsfB2T9uPwxA/XhoAYKSVlrJOTE2p9IczJXDPb/w71IRtASJlDQ9u4hP
uUHfJKuxeaEJXbiLEQlVifs1HZuITJqCypgSV1aY+qcZ5lWYmTXDb87ch8AXNHBOJVQ+l6R1w1jg
FepK2V7h7DbeIpJN2Hb/FOK+OHZWgKPUn3kvl7951tJ78reqrIAyfKI+DFuKtnPvh8loIz9ySylO
tUUdSgzBQHG7VgJu1+xQMIkUAEPi9+lKj8n7lnnOc698BZiyONC3QxdVQZE80d8zx8hzp1edq4qM
1lAy1lFx9E1ZGaNzJe/7tB1ye7kHeyH3soVBN0fk6ibjyPSjNx72MJH/BqYIo3NubuY9oobyZVS1
yS2BwYkozkAzxl7ubSduLoMKrg3OfrDFcGJE2zm/EJkkkc1Lio3eFANwgWTUFtqnuukyIN1ddzSh
mjA1EQz+r7W0ROHLMpQHKESc8xyUbfeDwmtcTuYT2pK3+n9JFyOHykwKpIWvp+zj+Dho/aT07QYG
yqGa4Q3hJdfGmrRa4Ixmbh+MWqGN4IWOJQk6dK2gj8kF8hekzNssJakvhg8SR3uLUvIlGy4ANQhh
7jiHfqoK7mrAwrnrAVMzygSFEa/76qa6fvj3zkgdD5M99RE+sYwBsPQ8D2cWub6JHBwiUkUhqj0J
joYwo5ePEm/6gGCLh2wxIrbF3Faq+Eao76ytOIfBqxWkWzp6gUBwar92HC0XAI/5Y3caKMGfuE0V
pY8siOfhfKp+h4mUr5a8qm3TPcXETecimd7JKjStZJ0fJzQjxOGYlrid0WEqnGbHsBiaDhE9/X49
qRZEbVQK/P39djbY69dQGoif5y4BNZ0l9KnS55dx20d1/EE/hSfxXGzw7rDh/P0rehrsnIMmoaXN
6QcDz2RKEXw3Ak7lB5IR4d1PxfgNA7RJQOgaBUV3IzmpJDm0W8kItAeCOU1guOm4J5HGP/lFB+dO
QYhnJeVIpKmgGGsoLadT2Emm2ggFbSsKcMhRWrsi6N3JOWnXJDsAAEHOZ+VUhT9Ot1KohM20VuQS
0sTKjmRRmFNsdW9mdWv2WYtPNsrc2j1dmE+awqKy9gCdXKCjqMTvhxEs2pAfRgKyL3AzmvC3XY0g
xvcxSglzXW6VLG+riFliktDF/3jiMiW9k28gSxhhwNGPUw9n5cvzTCRCFgqBKZA9HgAjlTzdFjCZ
w95e0VAOBemQNsROpAeZ+IsqMs2e7LQY8/93oD7vWqihEYMgHnXZUWeTaFNObxFW/qFTXJ7h6YdL
tzxbiDZbqUoUlIjxkIH9JNs/A9hhJbnkDOAcmgf/3y+ieyCeTVwung/f6m2nS18BGXvkpKsKI0KC
0gFcNuR0SAqdejJqrXseNUjHvlgcgrxP6sh4Tw/LhLakLH4wA9EaGSknpUnJXuXe56agh0fJInqu
W/rVl+xP/pqBElTIaBK9617oaavxJDNw4q9Rh+19ICfPqaCyudjGCavevYA+98i4GVeqJodUthXU
2ilfPizWw5AFNdSle5ERTR21AUaA53GBM1YqMNpQp2UUhwpwcHaGXRYrAXnBhTvwYscuKjQTP4jG
/e8gzzDKNWOyBDpahVLtYDKMvmY0fC6qgbs0wAQg/0QcjV+OiTu4iBlVL+bFz8yQ307BEqjMOVDu
Qc4ABxRE1zHo/I75vsnjSl43xfchSP0SUgkyAI3OAzIU9zFaMdVceg3UhaTGn2+ck/ENu6MtS1A7
DwRzfHoyPctBEYUDZFiD4UbxUyapcir6tdmYNK7vWKQT5SVwJsS3DbSlMitp8VfkSQHoEzytFlNv
NiYO4MMYsnOzH5zbRPaR7PB+TokhhZU0ZYbN+KKFVKH1vgN/gvXu+6tKZgLUMUhsGAmkwLdGPGiu
Bh9bhGXNmtOT2jSgPmXLfqPnrkwGhyuHXEwOuasWRFezr4ctxKx6Tgm64VQoLq6+ujnu3hvdp0nT
die9I3iLoMpJ3hR7V26fXyokJZ2Whf20CQh/2VLPhTH2Yf/7EgMI/rlk8aVlPiX0QgtU17oTESZT
eKbrStCpj6JVmEQD7ctH40BtPeFS1yi9/d7b+s/oQ+IUusAz/0mMUdSHEUpgl9IYIOh26jEKCUWU
oKJG5D3nlWW3ThP1/7qk8ItBcSNk6cmQXLIPPlU22BiXpAV59D5G2+YrWKRIvBbwvSxbnNWACkgv
PEzbbmLi2KGg5Al0xJLNBkcYccNpNzGZlZ+FgQmJdPP7SWszemNnq+dnKBU6Pcyk8XtuvTKhJoEi
t3Gd6+IVXzC6cAbBa8odC9bI31GPM+MUsACNlPGVQyk8pJnk42eMFdJ0q6VayLiQC96AIXwX8PPO
jxYxczd+MiFmaiKK0rxnY3rfDFIo383yYpcTiZ+rqMh7ZELtlT2J8N28zZmtZFp1SMrAe2UL5mAa
xUZgDiwDvX6qFCzpcW+jM/TyiOHAxe04nvEYJNDu1f7vGA1yAGcveJ9Dowf7S7RMqGnv9SM1PlY1
PSIsnkBVoz0bLVlC8m579aLEykC1iLkNyZxIIyYNwfIzkEsMpcl3QGjnDH7TAUlu+fCc6jMHswgS
D1R3ihLWRqL3JKRrFngxNqQ5NAaD7BLx16W7wEK7cm6NVK4XT2u2bMEncxvbr+gSm83FnL5xGUKB
05uzReXs4dpyUn3qffA9OPzPVM9yXFE78/ooV1tBjGdXHKyr/FS+GvV7DALnhnt3oDRCGiBM6yAg
RCePufYSE4L1v6XgsqfmLls6eIRbGTP53i4LDgUF6kXml1WOKd5tiUnhnrMySsWVY9GkvEnjvcXm
obaDFzaWAxo/0+lgWpDiLTO4JyOUcxyV/Eic0SwGHUWGmgY0cPsLfTd7ofMNmYYrVAZw4lGNl06j
9i62l7AgqMB9DS3l9QSOqvRMEMFyagJHo96/vlBLLkoQraE5jnhbZyJ1cyGutM5i53okeeCSLAcZ
VBFcf9eVlP8sVBRjaMYFFrxRnsVX6yhlyvxugnu+fQ/SFmI3b3RmqGTh3afIADMXQ5rg9wb5pGAG
8pb0mtGciwC9g14EptYcXCvCu26gVL5YsS/HOK3vmsNmJkUyEUgRNcye9iCAO3axiubmSOtGmhRO
xyqcvBLfyUi08YopWGgxZRLn0QX5fcISjiwnZgmnmpDN2YNGOcMd0OIdKT1y5VR7vs2VQm54bqqC
EmMpORekDnS1oW7Y0DeelstrfuK4w6uQnwRy/9HA8HuopX5Ck1q6m1SKxO6hBbbML8PCyjCWh5n3
WEgtJKie74/vIP3y6UT5+oiGH91nE3QRmpcRsrCfNBKdaJ3wrPfoA+xTu5JyvGUWZM6cpZSLzKXs
cbZMXSr+qunvmtxo0I5uxSCbkEbW13TjjtN+Wnwe/JnPuNqOxxH1ahTrvubxGTvjUBoUeyRq84s5
Yjj8nf5KTY7WcFnnk/r4q8KdNc1hbUDyiW0x6ITkkuXEM/WOMSVV2LQOXT9iF3bC7KABqdQYTwz4
63E08SitZ4XovEKM3pNuxPJ3lpkg03jmjzvEBlbZkjzRp9igKBDxpSRE90YrzkQA8Gg25ySBaoC0
mylZn8WC4CfHXW+bMIyvanTPu6md9BzWhzwkiP/NwosNgZvFzVvxUlMd8mKvPj1d3aAkfWDdwtHT
z7oa3w8RtkZDqUhB4mRXaOU2nkCqBFhKJDCOSOCJCCSX/M86DmfkyFbVqHO+2tI3ghaGi1ACWUss
oI/lG5AsRSI/K3PeIa2BN4tcx6osz04wetmQEfDipGJ4x1zfi6xbGLfNEQFAgmGHcCYDGJAfv0VI
+sX326Szgrv8w1zA0r4hEW1ypeBdXoBpI1hFi56Q0ewvEG15vtmaDOnoDXd4DfmY6qzTJSTBvtGB
q2H3+rG2+9K6fheqIUK7knCm3wAgAE8exxDjHXU0TJWPotg2qGfDqfGXWnIg9/KrWcUpCnwfc+Ij
1Hek+M4qN7BRY0dUkXvs3QbLZjDwH00kJcalNNix9mg0+AaAPt0shnDC4fnIQFWofbeWWc0ueXzy
nBWgleCuLC9JMQuRtSWRKhEe6Sf7pV6iacAHCKLV5saI85AiNVAE0pB4IUMynN10GylBphcEuSt1
i9x112gV6eZWacpxfawtAb9OWoGCunCnoiZPJLmY+24wp5Mywejfpi0TqwjUmlGDiX5WeWXQgtMJ
8kQroxgEgranA0L8pfN79oE2NWEfUfC/DadJs6ZKUnrXk3z2xDKQMMt3oGXWlZvLNXrXCeQTpe4E
6CcMdWR9c+rADFe9yHr2YoerxOJHcgdcZewH5OePzVUjmddM3KS2AnT929YYEYayXayuwEQO87rq
QM6pEg42G3CuqjvBwNXtbR8xZ+aMRfFlkN69GGv/OdxGrouomnIH3hyj4IrKyQa9aQyyLzobxuan
STM+zIWeutK745s9QFuiobE+bRZPD9uHzPwHe7lgQ526m4BSz4rWJ+Hq0l4WnE9kZ0t1q8jXz2xO
WiEEtBwKSkYZQOBo11EwbWLyHKxlDRAovrPUA6c3ghP+e0DEw9w3yKz3rC6zG2JJ/CI9Issf3le0
qJKigZ3zjLQWp4n3XF13O2QQEP1uiDsktH9UXL0L0hC9MCzbg4lEnzDvHgrltLJ9yayMzfhI28Bm
Mlb5W15qFl23fx3M11bOy7DGVap1h02FBeRGjkomCe/sm6ufSykccTdenV1liXupUDI6DYt+lUpR
PeSpeR4U+/gYJf0AQXtMu0iBZcEwGifDhdxIbeu7dOIrVX5jUl0VYcISLmKHDQqiOPFx/NWQr3Yi
iYXlkvpJXyweiWdVXBnU83rfDt1K/ADh6smtRt4J99Sur3XIjgvdcuNQzXSwkO+3uoeLfIpm6IeQ
Vh8614MrFPi6DfvLUDTXoKsa4mHjVtQJo0QWHQ6ItoHTzsNJ1PoUwqUtqP/KjDHA5WbSbkbp5RyD
p2Ide96wswL7RNSkSUt+qIB4CqCJuKc3VGyh3RDxsR9QKRmsmfkGyaBx4FVUyW432wsdV04zeQJG
vpxu9GSPtQm24GPq3GhYiQQxCO1BYEvBtSAr2dKaJFg7pTePtnGO/os6ix0B4o6yVtstsNd1wRj2
5JDirpU+q65c1TaE5wEKCv6+jA3MeJ6IhVyyxAM5HHtqa0mMATqwHao5c1d6x77JXPI+B+SbQbPQ
OAjfwdXLjNZs59pWiUSSI/oiytMEafmsiGrr4FcvJleaYmcRGX2GsW9u0oRAOErRx85hTgLjyfF2
de1q1IMVWNf+fmAG1mXjNPHhuC6h1Fgwp4KRtgksoTz1gizk+LBUERWWuGbfVWzkZVbsle06rtvv
MEJ0i7EvpE11/5LTXhfI9mhp7x9ZbLJNzXOLu61qPs2gnX2Hx+l3mY+HTRA1fxw2J4mIX//HhXvW
VKPttWziq8SjhQ7EXAR2t8PcfhrBBp/rH/2oXdYS7KJ/9Ql/7Vju5HtJnPc8YqKRTg5ARNiWf7W6
nrzK0HH5AYh/eFrnnAwDlpP6fCzON0maUbb6z+D46jXclj9wABgAKDIqaR67wthiOYv64i7+HZCE
cJ667HPKS27EpSxM/+HBgthW9pDDtTPgql04hGEzDiy9FTTNKdiz2Rip9zU6s2L9x1fz09v+zklo
v9pgkNbgLmi8+CO06gDC75ilmFydPF1OIJ6mEsC+mkY2L4JuQfCZnLvq9KhVWb8lChvZ2C5RKpVm
xV2arga5KV09NJSreDIQZOyGUpoz+Lv6FOlnVx96f415lY9+gXr2DVWqxd4xReppqR+O0++d8GHc
eJUX11ldXpVwAf1Q80PSFabWjeMvwUc3Yhi2/2nW04BF5Qwu7vnCPTg293blbXCqt4G1SyXwJAmP
fnu8+YdnutzWhuofzBGTAreb5XFOpxYqfyhyFBi0HPy/xvRDnIu9r47cn+kMh3YJsJR0OrIoRpee
m0xMFwS/pzZn57/pTJCyf1Z2RGCk3r1mGji/inSHOMVz3ka/eyvMk0wqa9eKydNA204WKi819j2Z
UzLQCxDsQg0RlAEGbnBuRKT4j0Gvk/WwBWjifzxn9lWga45p0DRP8c6IdX9BThPb8McEJFOdYG7J
OVvXPgDnoPJlzBZByVp+z2TE+AW7w87XAWcG8xY/2Jyg17+Tw8+Q8JnVtxf3GuZoNwG3telXcDdL
D1QVpI9t1ZdiJnkIEk6ru4wMCWZlTdt2dI9bNlW45IXZVplCHlDg3TqAoO+WvSqj+vLUaEvsKfXW
41xn4J8MW64UDljme+m5tNn1TNS+oCspmpGT7OrcdB30vipfpXFzevSshgbHVaM+xOjGIt0nWwKp
9gCWPqdOcL+uLf79pagVPc5RnX7x0QKQPl0r5Wd23wQit3qoEayK1JkMmPftDv6JgzKqwcyKvBcd
vTqM6PWltuMn2m8oihx4TR+tjbnQIdkPiJLOIEWrIN6vKX7w5/Tu4G3n5GTuSLx+LdpRxm2JYOFs
LSENUhYVIy0AXFe+CVmRj9weBAqo2UYwqIzwybLXzIRrreYmJBtde4G5SDZfIMAtkjArOyvxngmg
fJ5MtBZM9CJ62V4bDDQD0KjY+PVVkz6gMbq444Yx2nRp7Y3fZO0z6u1qdR2pK+OMUR7cHWC76Hgg
/CrDkMvPGMWdDybfL7AOJH9Gt0oQKkqHO0u3LWiE82bioq0uKjaTHVLg2DDFLVMQj7dw8AIX+4dq
yJvFtovT4eipcmPuLVQIB3jj8xKGky4nhIKMxSWoLRHcwafPLBAtU7a4iIr72sCsrL3Uhb4ffrAU
7T259Qq24Lff14kPjsrjArrfpzf3W68fJw8XlNAKePBafquCJ/QQ4Cx78gpRPReFouzhijocBtuF
bwPAoEPuUE0BXIImWRoS3COjGwneV4J3sjHfVQbtJhCNz4xqkQYbgAgb7VweSPq4Pfmn9Yv8uZuQ
HRuiiA84NqwXCwCmp+Ry7xJWvr90cF4lRNiflyjqf9DVkU6gD0UBlVBt6D31dHjx4sGl/dkztZNd
KH+JMX0CIepQnOGyOL9o5Eo8GMbqucJd5XIHbXCV+pAlE97cJb/q97Ec6UvOte9TmW6Kp79c3MDA
JJT1s4wOPLytyhj8Isl+EvH8pQSYEtYiT5tdlvkfx9sb5pPzcF/AALCgJTUpFUaoj0P/hC1yzVqA
45NS3hysOBxDVmh9xV8raQ/+xcPP/GmHcQsMmARiuml6hdZ1ziNbCUDIiVjPo8lsw/RhMnDD69d0
0c5nGukmzuPhiDw4hkHW3OwJM0ojszbLthzr/KEb1bhxGkaeO155GMXqOlydkECVPaSQ/qnmtqpu
5WkVxcUnGT9wbwiaSiuWtx9MgRWFaHETWa/OpLOiWldISr2ojXNngDPa7i8Oe0PTEMyGAuv/ECbD
4nL8oaedOjz1nilvypniytlJTQlgC2Dx5sdjC4jSh0MXuGM5NQ4mWChJSWC6NSGFpsgTOA8we1hi
zgVYzw9gt9EIvSTdyEf1B78eEGeYyTLLF7qhyPC2PkcgPL6d7QQWGdZ8q3i5HnUG0Kf13Qfx1WwC
MMJn4Qgpa33rP0Z6vGZmRMuXHpR1AVCDnjRWuOYs+NHiy57yZtpizJ8o5CkzJ19jJrhHB7KYYeGA
1FQ0jtZ4hmcvI8O1jCvIPT9wVtPxl0ax6s+vMpg0kz0PA2U3vQx6CqnHpWkC0Dv9GVkL7gFZmiBj
o7eQYlabPfLOT0U4Da7v/lPkNwYfAi5kcS2j/W/PVq1qFg6fUWaMEEii2so6HyuyfJgEoXJIo8Qi
AMa74jMwbIIPExUq/2hT2GjUNj92uDHW5C4Yk/+E+KL+D/FrG1ayGItNDXK1VRlPlEXuwh4/9tmw
cT67dP5eDrOlgFfNCTgBwqwiqQGl+HuWRZ/+GOP4KpiAlhY22Nt+Yl02jgXPiBwCFjNOkCXE9UbQ
OKehakez6vh/TRn5KArLa++rbtWr0fdcJofOpgS1OVgNq2PCBl6VYpAw2efqtwz11zVGf+/zoqoM
Hm20kuIt/vdYczUo7uDjc9rPa5GOV2m9fjWYPZD3mj26MIG1c79ztoqrjC1zLCzScU2pAxtSHGXd
jHKlUOx7NAhQuJZlb3ach3hikqB8+cpktEn78q7RXMAudcwUMWL8WTBwKMWjbKCUyilNGMPdAk7j
eOYdilEKeJMG6KOvV91CDGw3bPKpWnKVjnHTbUP3lqbWqrG7fbVqaTv7R3WaOM1tIlI4YNTWVBHm
sh0h/WTfPqS52i/lireBhUeoK9A7BtlvIfllBpva2mlUWEVgB5uZxyhha9ECK1ex0PSPsl6bgVSr
LB/TfYCErbOd7J5HezjPsTC4h8vLlsSevUAcvywUfX/3MWYfVoJywJIbmcE+I+hlURfp5HL5JuBN
2FYJgP1YjmBbV86yK1Ghz/xyTx0iLZCVIBBM4R5BC5RgsoUeyxEosu5dI7OUnLion6iZKKXGKH1N
ScZe2OiQsBubFaINbADalVbgQLrwdhu53/zE5nIUu/MzgbNFd0E2al1Zp6YOjMl0dDnwF/uA8Xt0
F73l+wQbfV3CT3swINiOR8Z1LbE5i7llHiNrzSEVYfHP1OBksgQ3SFa9z81DiNPV77CRdEI3d46t
n/ZZCvhhrNO/vVIGG1D+WVeGcKI7k3nyNeXBmdvIipEdj5ATeCaLvOQu/gAXNc8sW370twkkdRgt
Nf/D+LLqrEJgw0mlVGblTlQ7PLxcyOF4KlUqM80iNbaCUoE7cm7HvyYnRn9Y7tTO+IymKYKf3chp
wQea9DE+N/THHoYWuBUkbxLtwpLXyITrFv0457WAuFARTfG8sKfsWmRNYI/Ny7rKqCW2rawdTFIP
nCGYp8DjPhCStW/oOcT+8fqrmdPJGusa6xjHbIQC8ewovx4N3i9JYw7fvJuDhTgPoZXu+mt9hm0Y
aH4fDImcl2W9HfRf7034t8ttuu1oYr4OdXX8pnk9GQm+sirfToxsuYVavw8QLuFJNLyaFHsDgziP
MyJ0CvBFI8hPvmck+XTrYvV3EmxyJNIoup9irdUSGTrec/zvCPfEfFHApgDNnhjEYzAc+jXeMAAN
Q945YCoyyiRoiLHz4LoQkGP7W8t1nLUnXqgX78B9g1vbWKYlAYVROxD4o/0oPyPuP9C/7S06ge2l
4do8co7mDixwvjSue/GFw4s8wiTt2wdpenrZu0mWNjf2kmyd5CsWsjURixMxL+dnKzfUydsHkNPm
G9WFWfzN3McA7++GFhKz8mXqRaNdmSTJqj8GOJkfpkkIX/h7pDnlWMlECMdkRzCWtdKmcoVKRPPO
NRkosQtb9mXrgpOtOKy7v8wYCx6KdbtCbpW6U7sn93ocXDnMEq8mNZoe8/SEs/7lZWwFzo1jF339
GOFQq/TUdEByvPG1TzDcSSwpH8965M3qXR9nl37f9JNjSWyIWdRVlWBt5R9TuF/VHArdBPkSXxUH
0skKiEgGkzWy8oUQOu47k2cLwxQLLIeqIMl5FLzwsmzzWct5rak8CjvjZNgF/JIJZma8Zvmkoniu
pkWJ0cQjQLFFb4VS+rD/y+oO+PqhGxSVZLHNdjdbynMkMpbgceKAVARwRqWXbjnxpRA+Xh3sD6KA
TPJT/sArz/5ZtmW7WAk5GF8MRcEc/UgyL8BUuDoXQYb3yzEyPHW+7hX9qIhWCRpvBi8s+PtzuufQ
KiNvjQj2H/PlEzkVjEKh5Gu30CQeF3SdKhhdKfPopWmcZLv3+iNBIpiD4G0pk7epQsdgYVlDcApR
B6mITNNZp055Z8w7UxyFM2/Q5uI8Y8tRJNiUXMNXmg5SNHS2r8vr/8NtG6skYV7q+f6mqCC6YND0
GXd83iY95yFS37mUqT4cDfGqgrlWmD0Mz//cqZsUvUaJ+Tf0aEh+uWcz/5slpeEqqs7yMqESGFkU
BRMS+DwWb5RFBnTw/kWxzReoMkrXucf9cYWk0Yc0IGga3ikpMBty/jVEJ3XcH3ccJ4HnVfuZhPHw
MOR4aGS+kSHW59YFLAC4ul/pKwpR5e9ud+4mYIgvOdHk6K088sNbdg5IqKy5uAQAdtLbaWCXYUcy
SqrSs79hLOWPVuTP55T7dIGZxbgcmzOfPiUlp7W3d50jg3s0Oove/6qL5oBDrgn9/oCtS25UBuwS
+BOtxBKnxobNgG1H2OPvF+yZeGceliQAaKNRd7KXiRYSKUxHAG2IuixQDx3Py0N8vJJYf0N7eF6J
NlpdqEef4N8rM8ogL9rmok8J6m48WPHvm4PN5Q4wTdQPaApmT+IRVLCKdbil5hePKGDyvVfi7C+e
X8a5O+WH5rIsHVVFnsHZVtFz0paOJIMAjDUL4bfvPcA8ulobzaxAFzsMGwQm8rI3RY9KGPZDd1l8
bp/YHcMq3QMJcCkOD+XI+FO64MgbXNh9f8amVwsqCYmwsNpS2pFVL9Gq5REFh7nXBojEwugbFEFn
ENyvmFBj+tJOA+ZxNRHSDQwKDXMJFegfhnkUbYj9u+AK3rFJ+7GbWjGTsVGEMihkyjQXsaBLIe6M
7RlW7Ghx25EIZCrFPRuP6XH/X+oN/tuByyw6FrWuOf5Gnm5K4tX+GcH2zKG7qvVhGays8lwIxkrf
0uP8hpdfV0MTZS2OPZsJweFDni5uE9OZGXcLRTZIbM+xCZQnA5KbWRgYASOBQ2qsF133Kpep4mJI
HjqSEG8ftFbksLvAOJZa99Q4ifQRRh5lWRaePyrqUPkWhJEcgZhQ+Rrl2ixfiS1wMNiFPdNCkPxd
FWiI1ghuI6WIMu7yaX+NGpopPPoolxP6kPajJr0oglJCzD4vY9Ny7vfiNFI7O/XmMdeGo/QNfr2v
xDUwFNJhJxUJYAOqTG0MXB2PpNoe43+gn16OTWbdV4LBKpg8kw3Csp0Ue8aB/csghviVxTKtwprD
i2T2YbbNMMeDYNC0qzdzlfqrkOw4GR0vrLTOKTbv5H0kdbO8LdQpZDEIEO2YBQse1deXo+OpWT6m
tlie4m+ll6Z1f5MwdESfiyA6K2ZheynMiy1k4h1LHVLIBGtOOjhtgb7tkcfmK9WRWCuQEZZ4YOid
3qwecVR+eSWtxNRSBqyesEC+HwP7+yFPQdHuCoIB2Gz83XYgSLolXFWpuU58QAc30SZNyxuQxOo6
Wv2WvNdEtos5jQDHd9A4KdIsSSGMw/wGuN4nJTOgqVZAKdnQTDwkaapqV7AZVB0z6WKnwvHFnJr6
J5f7C6Ud6qiVqnUv8srgEozpnPWBECEzzb3+cZd3i/ap7fr+gDwtQrzJUm/CUTlEv8YSCO+DLqbj
a8kELuGq/yvPsHU/OynmYHkiOUCNYatcoDTm44vPRcT2CClHKabFzJJMjA+O6NDqDrlzNz2ft/IV
iu7oE4mJoB3QdTwiShzJ7QILPl4h5fdecttgGzcrExsh8SAIwk0/dC/R3mmNYVmG7E9toHMNCN2K
6jejF/Gw96kdC0Jdzh88uIQotpJI8N4HmD2s21/ws0zR+RLoxS+DzVYN/la/oKAw5EUVxnxT8+Gb
v+rrp+vWrJ9TXwKCBzasb2624nhZ/x3vGzc3QhyLGTITyFQj6vPxSC74SV1dE14/D27r5wHuDlbH
VpUeQ+Z93aHEtdrqjx+pPTblLxoV73RxXU6tXujr0NtgXexr1khF//ix9JD20gP1XTHsodD1j/Gd
HQjOTZHpHaUvN1UUkzq5dLFCr8zuWAnf73s1ixkeuGbI9qX7nUbGJB31mFC3Z85Km66N4p4ndCr3
EdgUBZFmoK6QW5Ubq+BPtArPaAfHcRBHSBTwtDMCLKbpdbUrU3Cm8A+F1U1MoGaaLTw1+zRBKQQ3
XzdgIprCCKxZXyUc2yZ3aY0TReUXDPDHHpsh6uGiNHOJapZLD34k+wDX50n5yH8sjjSMiiZggfX4
sqyQuoMZa6AGHtZmk5qq7vdgNQGrlLl8Zyep1EUyIfHnJl2Akta/KwjAJcJiTJPeuS9LwlHOXgaj
KRBuv9911oiOoDZfz1VN6yTvX2Z9ieJG4h7mUtUR7/iGE+XzbE1Ci4RAXiABIdYsS6BpoPl1r668
hWLmDBKD+2wvvxeOBJs8AGjuxyeMRhzKg8PPg12vdTa/VEpCdfa09jPBCLDcdqpr/A7Jxbx+soQS
jPa6ZGNQSTZP1y/K1e8h6RhjyvE49mqcMmyIdxRm5/ZywQ23XoptH4xStLhcPGGlnwc3aoBRe+i3
L+/TWApNXQzcy4V1/9hKdGIzXbw8uIlTDoS2O17fgpPkWjmqy/MdxoLxUuEMnAr4TWUVwPWegAaY
+0amaBmccVbW0uflw8I+JsePXLDRkVV/71ZXv0TMu79a+DGRemuCAYCAXA0f/S4lyx1QPJ3qEdb/
Gyy7rNwK6YRnxK6d4q919ntSy3Z53sfBXT1ZUlDFTbsPRwgavq/nTZ6cGYzR0SrRU1p7bsOdVLeJ
SfqxMy4QYQCYfUf0SvuCIb+3N7MTZm10pB5V2DcCUsQG0Q6SpU4+F8COOAJCfsADgOAfuxtvZDqQ
8ISoWZFG/vMJ92Uk/KJwulA5FoaCgQ2ReUclG4IRlvHt/t5c24zVXWkHyU8YIzJ+vKmj61CCjOQA
OwEJaEsqulQTk8iFo1YQW5touVxjilzmMKov/Xns6EJnftjPj94U4gcI2U2jd0/CXxJXWmFZNIET
BpHtTotK6ogsBlzKfHaMHgWKgj+TGnr9fKPXZmQAIL0gD2L5WntTIZvKPEah6XVXl+1CVyGdX4Pi
1Sin9zlQmgqJFS7t8ORHB87pDJ0wWNkyri6VrCwZNN23tH8SFb+NVaidqIKJZj5m7wynC6W+p5Mh
QH+eD3XwYiodPoTXPggfeYr1lTe55qQMPEM6T4hcivd1/IHNuWW0PicILesgwIxQHsaIGooS5ORS
Fk/v42JU1NqbyRm7CfAqPwt+ceO9pOp9rD9ehKFC0IGry/V+bAvYrjy3ZlvDIKm2dSqJWDzJnCwk
TSjVKe9RBUjqzQt64z/tAm3uirtlm5BdZu3UPpYifONlKqD5oyULyh3ngao8fPVYYP/VHmTxmEsC
VLaT5fH31T/8P9wHVHpFnbbKX1Sq60PyW9JIk+9XJ3hhIP0Lv06u8VfdgbdvLn0R/7GZRrI8oZEm
XTLCH6lfui2lADzvbBuyzKp2Fjce4u1s6BKBByHvGSvNVAcAyA1Hgxisw2DUPecoL8cPWnb38Ht3
x97XUQF+YI6KxMFHj12iE915S4dPT0jfNU1D0LqwNjtyXww5KUGQSbIYHBxF2VAcktIWX8CrKzyh
3g/RgdM8aUNcXOpWIVI7I6EGjMJ6LDU+2GW3NgTk1pTvAIgZcP3isS3pKOos49SGWN5g+CSoU1J4
+7876VnrreBxb+GphKFKHZTw12gqdM7Lpbf2aOJEqb4SmueDw3BnERKGqCI6v+xbUch4jHgtusl4
rihxX+4PK7qnIKXXx7f+O7WXxohRswNT/5fiHcubXZj7VcwzhJwEbQm4ZncxIZ4CpERo6aRrs4fC
l9L201cmlKBJ49Cogn4QAW7/HeB21sIwkCbbBradiQlIDgTxkgS959zapKkd/aFernc6PtWf7KJS
vebUpp01razBTHggtiH9q3B8kr+dn7CFtkqOzLMbjnwG91tfmRHt2laeQDPoqZuGHQxL7RALq4db
ikspSdYMLf8XJBWrhv5Zkrmkl7m/QQ1/oGMKCiesTX400rzZ6CINCSJgXrUQvTA6lTLOi5KLBRvD
IXsLcGnp/4bHodqGHH8KwTKd4N9pW0zlYqVJ9oafBJVcaPD5hsolQKHrhg8CZE3TJKFs9Tpv108d
g7y2eYg4+hRrWgfGSsQ93HBw5wFcVq5SDxN0kwItYYMdY7RtZ4lrzARvDdVInwqElln07LpuGgZT
BRWFxMW9zntKt1xL2p1R2LFtSMLTuqFF9Z9WetqekTQIFmJCLSpUBqTFBK+ijtTOzoC47zuo6pwG
AHhPxOsTBsdlITDjILrHYyRRIPzgASjdfT7NoUnyQn9PXRecdFgTHUkYn70C5HM/UuIDzUIb7MHz
OmC204TuprB812kKgLFXdmkELO0TRm9u4ocdR2K31CJS+wTFh+juAJy6euYBLnw8gV8s3knkEmOi
gJkjF9qyI/9yhAmw+m2YvJVpnuz3BNJhclzrB4e4HwrZoG7brqbL1EeOAI+bFnuddlffxQKivgY7
j2J6PHC1LFEBMF0lmcAX5j1S5dRtvtwLfIYEFpFGJ6npWWDdDdr3m54b5FjpOXSAmObB0acRsjfd
a/nwbwGOobToEEUgVNtmwvPZgq/mC5OGtu7zVxK4rOwR/fin3ewsLcIsyzW3tRUQn5ayyc4yf/Ui
vfVL1C6nvJEFBJ4bgW4FZqqRm5aLUq+JOqhBmz0R9JLY28lH+9H6j5En5TUFlTyYzr8CT5/Z3Km7
/DNT+Q9wz49cxfG2kJe20/4h8bDox5xJlHbnhoHgQWhtCGzYBYvbNuhaL60LoiCwSAOunyjL//pm
5uyU3LPrfjap9bGDXtzDJ0Ke4Z66QjGD8KUpVRi+n0xhb2IWgTDI5j0W8If8+RWapZ0ruhgpE315
kxs+gU2upo4sTgW2JBmaH/tm0iJK550A90ZvOL5h47Sxmqxf4BHuvGtKDzjn+NEnOmrp9FjwIKyN
dBDrjSH6SAGUF2P8diknLBNCfGD+EdIhlciBMJfVVVs2jmfqT/ojlsuy7wDhFMh1dnWeRZ3TZ01o
zWZAfwUdzKsfwhJGZVHoWWbaaw6X5lhGFFBUEqOct40IDsg+GIZbSVvE6Y1daZU90xXnoHaa+VdT
0F29JrmLv+MV3JdEgMG1Pigu3DMr96JV4thmphkfqmUnc7h9FZSa0eH3YYErsyc2jkhbU9x9BGBw
YN8ZJjTLAPLhe8TChkZ67vxIOcrUVs2W9TLpfv0NaKQzW0A1HyEZgvRAY+gPJc5c7yDTWF6wfOLt
tbaw5bk8ersariTL1PlMvoOu5GYGEUXvPf3vofDx3MLhH56nLWL1z3duasjiKcV7sd9SWBCAg/Lw
xdxLxkHVbmNZSqC9jO+4GhQXSnjkDGi3GH3JwOLNqo3fTJYfiMv2opT21WdJ2UCoWCf5El/+nEvx
gF7p3YewArwc4RHogty9VGPiCHfpyQc0HzNwuE72Xr9QJLerJSYa4RoBNok8kev63GZivU87JWyl
DHmHmTn3a3MW8QdujFNCyM54vBw9zHo0mVuuO+7nzVAReYRktOU/urB3xMUI/TbgGz4jo173tDKT
GBbOAjfgqreVUY6XRYRQyL9pS/X1GJin26r55AIHMevZaX2J95oWjvdb8QpYgHNUv2d5JI2LXhsD
I3RN/Yz0J2QtB3X6Nxp64bR76fq+DjJBy3QLJxjYT1wTidUHPTromyziDccSCsoB2bB18rECK5kU
otVx2QP4s2BBv6wk+AhYMLOfMvPcMaAT9AP8uJxsy2BfbPsUin/6OiH7LeNHQk/7270HWYbfWq2J
p2F8Do+dQvmMuoirGRJdtC2ek54FPqQoY/D+HooGc5qfVc3fRXMbmMoKZch0EwrvppnekHyho+nV
Mv5iUtleupfZ65U9Pe4Sq4xX5CyaeJpNMVcDZP3zHMcjIhSKZ5rshZ/3bqfn+GdAt2Fl3lN3uuGN
IaJDMCCnkXKYIlxuADmFHALW87Ms8ypm3CB6IvjuMC3Ojzn1J+GS5ncfz7EWdYZCR4jKnzhDFugq
jJEINAwdqrJvPkq15Q6lG1bKAU/WCmsooG9ZkCjyTznxi2hsAi+zvfbFhOYuOtH0ksQZHuSWx+oI
kZcrO2uH23sylQIz69/hAZXRdH24+Nu70llocnH3GKa/Z/64HK5R/tmPLRQn0HmxrzKZ66kKZGlH
tTXGNwJ07uLw7tT4CpV2KM4aSy2FNfCuegrx/QSjNJUpg3CA8Wt+EKcP+EVPVDL6L5Zu9GviMihW
MuX8WueWsdWa3qwzI+EmXQeQEii0T9xMJMOtc/oC9QAC/sqKfw4Q/U1MCQyPCibsxtVXnq6mvoxE
UFVTkAUitVhk1EfP7s/zcu5hH7RAMVkvIMrf/kjcPJj6AY+DYM1Fb+cm0KwD9+adRkxeoQi8tecL
u+KcT58PAqxZlR5Lria+HubfQujVOB9pBwRP4BKeR4V3EAajyr+HnYRq1M7kF2xjz/ukWqiv1lPH
FIJYFCFkvAaIxK4ScBT4AIEiD2gLBNFRNSCi1k69QBr9smZ6ec0XxYqoGDdL7BZ95uER4uF/z8Lz
/LstsEO3f4PHjP+6W0vXYStCd+Ajd3IYqcgGAopaQmbTzDWGbutpedDsutPfqenxVcMbvkhcdING
4kCvKfy2mQwAoIXbCf7Ca7UyiTiHWM/0qLFXHVcN8EHbSXlgaxy8UKrqk0zrxrcfI9ycouMNQkPW
wbvMo6zuHOu5xHJo0tHIUOoYnR6pyfnnmfFuth/NHZJfSamoYCY4McxVH0ixyRr2Ff879gSkl4jr
9kmzKmJkO1vA23LSsz7JLfyOPzmtDgPabaVqBp9DApMlOqeECpJZuGPx6YqBLzpJwurIJk5gNp1c
7Zdl7DeuV7aeaE0bwTVq2tukjqPPzeLiIQTcXnona8T8iYGnLy7VvCZH7fWkWAmT5rrC4962Ja/8
sa1LYri4QH2LxqUSCBW2mfUi5XOOtgeRwYWIk8NFIo1S+E6YyKXXyc0E9Klr0ekLOqt1QaL+zRU9
LycgYb/3WenMd7XHUrZNixsOO+M9oHh3BERCqANGL1axArfVHSyxgQHW6a5UTUiEIShRnXRJ+Q4/
5sZW8FbXssaS6eZ2VzKcCCAqflPEju/VZETy/vzBQZnSYFMbFIM2Z207hqienz4vNAFF9fIjrub+
feluk3SM4JudylLy59whYuuEaajBl0jdL/zFe1+fN6h8mkZYLQyGbyf0JUC6M8SEctDQAtxhzmRZ
0mAEdaYJVqv8w8M8U7VDOa+HFKl7rLR4T8CgQh7K91MG8Lwd4bac+fGjG1PkLPFFJJRK+GGQQcf8
wcbapwW8D38S4WGIKinVSgPL54nfJVcwNh5+dQ8aHXFF3/qeiK85p8ckGZ8RagrwXDyZLEqP9ipO
2hhdxz9Im4FzykqxLSlBiRum+nYCccVh6rWchzQrtESa7BhPxaweFWFTnq38ccrfmp6a0z8ysG9a
qoYBnSvvePzMPpQS1ex9JrK/AkejTsu8YD52oYPrgo2QoW9VC/DVF3b5kLay9/NS4jO4ee9XHwyv
MWLtR2gGOFWWw7AHy+Z8HweHMaWsUiNXLXRuStkExS375Qm2ZvY0JCn7ONwC8Gyh6HUs1vqV1Tw8
+2vBV87N1ZN1eu+16NmmhhD5GWSZnL8Su0Kf7htBLl7vWawNeWYxWNOXZpHEOWAptqh+DkwCqmL2
1RE9U7Z6fG4tVmcQn94fKJQ7Jh2RMXzQom1QtreaH9KBN5JAHZW5ClguG6QfuGAks92LE+JKrZBS
lemhtowocVMvGcou2sLeJzHnQ4UB6BishSs1FGW14fi/nQxOD1DexmD5eZirtywPHbIicqKccQP1
OtzZwZA2icz2RRMVPxgQGJulNp4a4R/IaXro+s/UQgZ68YOYt/YsN2zM0i63N0wh7ihnZSuc/ilY
fpOIFYt71x/c8hMFCj212i5dA6igq0Gk/wAy3odyA3sgnxBvaZDbMUKyfg42a7dE7hjRFcR1rzYc
k4Y/Z/A5aBZAydfz/jGAUAGIXTWmdLDVmMDK0CGEVcCAcV7wdgH3MSBI/pU3IlbwEQOd9ixm3bRA
xwXJbvhh7MFCJQy1KAGAd+6tiTMbx3gWV9xC7pdsqXU/giQiF/FGbee4zA11PeLRz/sfpBLGQxQb
rWqAvnRGbLk5atf/7oNq8/BtTnTLuMiOqREqYYX3uwbUzwYM3744Am/t0jQ2DM9vjgEGUydMsuIL
mgi0vhue+RHFVXEPNy0vftX/M7MYfleuFltQqkRYksvAUuSv2A+vtlTCC0J4cyivv96c2cozVwmo
pyKKMvFxG3uTkyUJ3J3cV2lx7RUhzxkBAAot2J0AmiIz24020lbwOF7rF3vG5HLN6rkIcz8uHOek
0gjegNbh04lERzoN0vj15NFk7vUNGSuBm0ZTOLNXB6hmcY8Z22Vd3a52qdf458xSWNu9GpBK2CjZ
Bfe7qocHYgDdBPu4xAN2+4Ul9DjVPbvCKiCyQLPSEHTQYQKSkOZ5IF8Lu4ArQWCoQixinTtvvh06
IlyIpoMlBCXj8C6inqv3L3fQX5BS2FCF89aqEpCgc9Zvjz3NuRgUW3+2+D4c6t9XAMv2/JBrQGvc
yNPiEHINjeiYJtYHrhfStc9ZiP6Za1GEcwiV7Mcs3JPy756+wAIhdZmOlPkADBd21YXajO7RNijz
SkzCVuy29dG26lx4HOAJsBbnyvywPJl7HgBcBrhWa6OFbd2uTuzn6fp+0fUtUKVScu1YWB81ojYJ
js6X6oCsKrckg6qomE85T5xSDoMnohgb0Izn6H03S/X7VLMZ6BNSVRWLWU1qFlxeREsP1ITYbeXu
zJoVObLdKdKfrctMNRguumVT4TJ7pkcD0fkC+CJoNWvu5N+JiKnxK+A1tgLJ1GdwGGITUlSYroJB
sXlMqAcfiVWj4l9oxiHRlpJzlE/pCopRW1z24q8xFzou0E48bzsPcElGPYEyBxVegVBr5baBlN9u
JE5OTtpZJzNn9lxwm38HlicSRuOuRXeaD3VtE365QCRF1Y+CBMdCw9/x0JuKpbPpiNMEyFM7bDzo
FeKP9d3wIH1/8jfkdzi3LdEmBA61BXIeBMvz7akokT2PJpG0TLOeo7FXKdG4q+LzWIEqwySSqTZU
00qf7kEWZnpFnrPRhKZkA4bm484mr144Zor01G8L8DQ9lkwHq23sF/7oQJ7L1Qi0sTe5xRq6wvpR
c2e4V9O4vz9TrWJ4wN+nynNcRwL6z2ysCXkDgqIniISvIuoNVz8K5w6MRGKKsK+VjftwRAn0rqWU
kH2Xv1ECXDfp8oFch6ITOaSZK35rlpnrCtEKstCJ8kxg57legnTEUxVnPUCGPklUSsL7NAEaa7sg
DLMLWC4XMGbsh7GIE+wMUYIluZLOxvmi2rhqhX4S+9lptHD+jVQERoQz59oEd/6Yzuou5S5XfpIT
sOr5fXM9BuihVvRFgQrQ8MJ6LyGxffy+mvbGHIc96GdkdQ+8a8QbmSzOvJvanFHysZkOhEK2jndx
pSBqHFSfrR+zThhY5IqJuENKBKh/OG61xU74znNivuCKvKzAEuJxJMfOiUgZf6bnSiyQ8grWhjnC
ZvBuXV87IuWri+DJnqR852ub3+0F/OLqDa5YCjaNFNmgqisuxr1X9ellFrjFUfhAaYDJpvkv1QEC
1llXDR+N2GHUMy3zbRWzSk9oIznzV58M2dqGhLTicDJBogHQfCpOHRGfMEIN7lWUoX3WQKQePOtD
PgNbeQAxiJ+L+8gUpnv6YqJdufrrfSgY7boRnqbLPVqfa3X+kjnd1oLvwdqbeabktxD2BO3FC+dy
267aRrZuXvttz4D/219IZP+zat3Am5S6wtnVbBfIQ4ZAy+Z/VgObaNMH4rYfM0xwCTDlRNoxvXkC
LIvuRAls69smSAfDMdx+vBkApgef/NJbsyVJq3SigZxSIKsl82q3dOjODqNx6lkG4vuB348j/4w2
owrsTufputJ+aogKRi/S51ROhCjfU3RFgFKUX8wl7UWWY2eKA+30m6uL26TLMFnwWB2XHDUGMNUH
KXnZnwHMyXAAhv3sOkbi3jW7Q2oICYVasV9IGtxPfE6vwv0xqlNlVJ/WGYVzqbKBiQwcam2qhyl0
x7LZipSxgIaaCvZJ2qGRc1UMcnpa6fWTO3Jyo7Ol+pjwdVspMssP3dkLpl139vUNRxUO0Z38qNBp
KYRz47u3aR6LuIGUqlAmyuTzLsk3bvVQizqWTiB6noIx8bti3YpIEwR1PduVT0oegpTqFGMDUiiy
juvW6aTs33w9tQ7l83mghhSJweTZG8wKJFszFMtOnDCAd3oKWCUXG0hPaYJ6jkmzdzhC77rlK7LZ
kr7U8+ycPbGsfTYFwg0V/4uT1RuNGgqU6sAQZVrZF/m2Tg/qiOAJ4ZRO3C/Jo20fo8GtN49zeRR+
q+0kR6JGe7NgTPDJnfBNnOz+ftfGRk8hIQLYQSklLbsVgoLHchXcSKd9by+X5mAhUK0JI7yoCNsI
VzYtrQqblnUsndH9qDtiCUHPgnD62d4MM+YyavF7Ihl/7ksgr4Pxmg3vHUedQCEv+aKa78Oo7+2L
0qCiRGmrO/qVpg55XcGq03oPRL1Y5UJ0vEsVU3a8sztw0tf0BxlpiqWKFE7goEHeMHW4POMa9DJn
jCy55xmt1V5O/7blLBqZqnMEVC8ef1h+Sc9uYJoUoPUaa/SHdJS4xDcmOM8Nlb5zXmN6mZYDtbOA
3CVpezWEXl36DyAnVXC+PqNAGw+lCT8oW2rfNC/vqFe0y4Sd+rzFb+nL59qfFTct6shbHdsFagP3
mINJro2YdxDby9RuIt71BhqunZ0cF1TQVIVb3ktl1jxB++MXjB2iSZeipkHvHfJPdxvmo5iiq/xf
eoQ/cBkP4pnld+qPW45QHp8EwCuUnSkCAfzt9MTcCFvL6ovu8jiRs59ba2FBS1QdMvg9m7tOH3PA
/1UWjkVGbGeTP/TmNqd3PNAGvnWkzL18oZekslKOhsG7QyDIYXlOOm1fe4FgmC9Q6QVgrSGllOwP
iMIYKD0w2SzqLa2X0b1ACQ++UJGCFSkyL4SOsQF0repaLZinn7AVm1amKM4JKj2h60w/8+ZzW5PU
SY83YwvXWZEjWeBhi3rHHS3GM8YiZJBp5aaL0IsqMjbmLe0ThJcvKNZYHuZLYkPivv2hAxho68kx
8MYninuDg06d3XsFfuYbxQppaxWvqKJ+QabGVIOVuuZU1xRNx+LV7i+xZbPJ1esXYCbnLC06FNDl
x/IVpjM1xt8mBhESZJCB0jDeXKwy5pGxhSxAaK5YigLE5mReLS1UDWyxwovajH+HD2y20jE5skss
K8sFlm6TadX5xddRnO6KQwUqZI0u+e7rWhTmphd0VasnawtUn5XRiEVaSqNdx9yOT9X7xS2rWJ1B
u0Wm777+B1uSpySZPjkR5mvAWacnKgJgFg9jrdSDChgj+JmgKAWybhgY9ikDs9D4Y96hCyfQ1pys
KgKidmc3R3kZh3Y0/aLftkfVVIuG3tS4nNOmoZTJj0VAt1ESu2RaEF5714M4v9Z+czRqjvY2H9yo
Qdu7B1noJB7gs/JL9HRVdFpbHWmeEa3F22I0e8QtAR+cTBSsQ9gOeAhSV/CqLPNyEvB57nmMvmqP
I/MyN3vj2FVQWzlhFpgJB4O6J0zNXcx6TuSkoYzwmqblbZ1MQs0m8iZOb7sre2dJYNqEouDxt8z1
T/yTAFRUuJie6ryeiKkAWpLbYljXTdKEQhPx4PqnRFteBJIxxuXtSraQp2KnTecVfiY1SzP/33y8
hIQAKq/bI24oejo5VJcdgSjaZgi7qD47xgJhU1Gan9wvddlgdGglR98E7hc/knlUrPAnAi4buWOV
ScW4+kk6W8vY7HU6V33KymJxrowUd1B6t/5RdpHJiDxBg7Uu09aurNZVccNCIf20STcXfUDk97H9
3feHaQsT+MjOqDQOiLpZUXgp0LwO95ax0xHX4v77dL4UHBi3wj7WTS5nw6rCKW2fhZEyki6W3vi9
ABsvQwTsD3J4IW+bt17SaauGyzXeOex2TTfCQeL0gprG6GsFWEQoIok2QouD15fyF3FpjpHTaqJ0
xoMIPGI5/qyMEys0N+eJRJL9ZNe+wDHMOEJ71dXoI4l5cV/IaHYfmeB7gv5BVgikCNhWcdS63a8c
N7U+fqgxe+FS7+y95UAIg9JS/zbTe+L6YHOsPbliUKxF747iM+58UA/C9xrjF8dcG98kQ6en6lNK
RW+zc5Mgf+rP+jnq0SKQCxuatvQ35S7Oq5V0iUGZMnVJSOVTfKF/A73GXqdhKxX3jf2CLHSp0vxB
xSrvSQYvXItTHrt0rsLBxQFjDyVUNF948hZ2x8xk7B+xRALGz1k8xkGvmB5hn9G0SHDDDbZEUCVn
KaqbREeXVnnz8CGDwKGbMXq54fcR4uK0wHwuYgSknMv9xANA20t8Rl775Pnmdgn1MklaV+v0PcfR
zqfjl2eIZucseFWTaKS+zkaN+exdVBNlWZ2elvJmc/WdAeA6ju8zSF78WDcTkYSusbz4xP03Yj2/
WcyzW2ah9XxAf/8yLnNkLP8bvLiSlcfE1z2vUCHOEuQbVu/o3R8SWuISxksWIlbw4EayrO2YMeq4
pJTUUd1QG77qpgL9CP6RuhDORonmfZmYsAw6KMg/yXNcKDMrG3+4qmj2xb278cuH7FKdbMmiUpR2
2UNthkaXc4+xxgS6Ls0MhraWKj1darAOB9qOX3KyosaAKAR+dHJTX/RV8VGkYkwtPQxiLMvkrvw6
3YEaW50rRJGIZkdyu7+QuTxd1B+KhQVqv+eNWCnBykH0PR4mUDUCEBs6nI5KCLeHt0zpsD7MGZLb
HkngZUoUKjTPi+sj55/x/1wUR9FR2VEbwPhQ71s6RirkmQCKvgPBpA7tJoP4VVVhtcpxQHOrgMUg
iH1f9PFBxKW8+WSdboIj28rNSDIyptGlfWvKnxK89K5MIuwlYvZXEqIMC+mdAEf17A/nqfRhUdks
JtGPHc1NWay7TEzW2Gn4yW5CiV+TVwaLpe02cUJ/rtGqWZP2es+q2hbi85ZJdfY0sQVf6TeDEX8a
BDfsQvet9wP7KuALEPnAmoHUj1hACFSuwB8hqLMB5OQLFQO19nguB//+p5y1WwZ2EsTG39p4eo52
lWSIb9Kmi3E7uWH3NSVTitFBaReXWN/bLzoFpfvtaLMl9uLlEGkPN7LC2JWeOkxxvvN15BVMF7cr
4irjZSaZQfULltn2GnnQo4nsp0BdJLNPhu2Veb2HT0oS1Y0UXAi6D9WpfOsDR4yUXyn+tfhApQv3
4pAG2IW+2GDly6juMpShbBDsR5kp/oHVxGehJ0YzczixeKvlXs+0J+Qmu7MwmvKBhY6hJmAF6cLg
y7Lq+wcowwD7XBKRIK+6SnvP9wVb6iY1OmUu+8feGUw6VWlKdo1/e2e3e5Np4qnjneBrFhlkG68g
ZLeB6yoZcNKcIlturyyc4ptQ6Idw7qUNbMbLpHQKijWDxF6JR6pFdpI4+Q9X4Nd4iYU6Q8UkLIsz
GA5jSoiDLnPWkIwLGNSleT50J9w9uIBuxwOODuvNqY7vZElQ8dDnygOMfvxVCC3DaUg3m+otIXC4
Ra0cEhwWpyWuVKVXZK12aXXzhlUvbxPGVYGEpeFtTtcvnT6FuRHy+KAiE9tmGvXr3dmcwDZaLOeZ
AE5vgSZkCgdRItvKUM9qNLy7ZbS8dkQk+NS2YWhX2KSRdjxr9lE6fxuxHFNYl5oakMncSUpHefRf
gJflWjC0CTVfcD1OK+HT+qOqEWMHOPmMdGgGHjeGWIbqliS5KNvDjre+OG1CRmXcPuxD615pebB5
hoRJShMmDhGCWu1J9qmaoaygGg8vTxPFjV1W3ngz6dQZhMKQXUpuuwf7yrUYdrG2hYAwb747U+ee
rQRYUm3TmaAB11NdYQX+W2VDabsdjQZN3lpYe05jKLHnI+XA/RvAbMKpjAkfFI8H+nuzXwDyf0Xf
EfHrojG/9FYu07EImKAVhNW95LgB+8+qIUp5t7fcOmNu5JkXYI7vGwba6W46RQJVhPFBo10FCshv
hOBBxoOnkD7KMqkQqc+tc5/F8xQSm92LayxfKZIVGcBPt7h5fiPirPMt+SzhW+LMaTnz8l4BruKf
SNrXiUzshsYTOYsgfWy7Nihw0m8PmJSmFARZEqpasxPkvF2/qe2PYjZomYIzkQAT1qLhFwOXtd/u
dfZcsKYLyoxWxyIH/WsvsRIZvPzcx76T/39k5/Xxg4D5q3OVOuZyf0Yk2ma7qjV3gfat/MDdwWSK
KMUF8hv7S3i4lQzeC9ktcdbpJIwkKmjhoZjXmoQ9L9aayfpK/GEHZN38PPFMZjBdvH8N26EzPn4h
gVn9nAzHjPXnB6wNkoHon8xX9mEw4rGyrOPEzuKb1mA1ATiXKO+irDi0bpq+AEmmQBm80/17fasz
JMnIhRo9dKJuwafF2S6E7y+sCoxYa5Fc9LPkK5ahBRYflsrkhuW0N25PLEKgoQbT4omC0OViNMcs
vqAaR7EJlyVHEgsoKQ/jET5kHiJjRDoJMKr1TS7HBF7WM7s8KNsFZ6GApk8DvgUS4VGZKIZqZEcO
TF5q09bfNAfOslwCcC7otbGmuk8wcjrPWz5JBaPgx5+fLOWAzYpF20iqgYsFcxcOljPKQ1LH/vhS
qNtvt4of9c26GFBM7zlAfA23P88cpS3SV+l4+flC1rbtha9fwZ3TU/ufrxDaeq8jJzu4qsffrOGc
HTkTZfVxs3RwQqo1h2VqotKhMj2lalWlxMpaCaGJGcL4dKbIGbFY+uYvIMUy8EawTqLWpgiUMFKA
OvYWKF6wn5AJ4aF0t572umQk3UJF6LBKnm4UdZ5aiKW83yACbbTzdagvatmzE9X+oYKXnESgrpLV
71sjKTU4ql2d94aCQ7xNvqzIdO2L0yU24amvSKIQ9zHh3xrQDU+mZjT6bWrpj6QF+wKuHqtedATz
DqVAyer5oyHTkAL0Y7l4QR9vqw+FXA8HQCuRDxeBatmMp7uYVE05xcKVr+huj6xUnChd7gwUDCmr
1HxtH/daG8IZGKu9GtHuS0cy+A3o59t2C5+70Soe2bN7paOGWgG2juYsJaCpOvZUBBrp80iLbzB1
n9BmMCOhx6UF0cmsAr7HGVKKiKqXNYYrM3EzOkh++op7194XtCDpOGwmFl558nUknTdWJ1v3U8r4
yKs81s+/cN3JYzftTBn6vHiAJl7or2fg2nwW7DEMfONB8vmU/dxdy5VCyklu4XrKKdFkagSR1Qiw
CsFehY6lnLjNeEvREnf5BTEAGt1JkihpuE7bJqjfh5kNfxhQxEJKtk72cqbxjqskX/+hsGHJdWII
6f8NdTidZNvxbxXJomOLKkfPita7jk9fFg5lvt9RiNeuI1nvogLV1tvMD0KlA4T6CM0h+VQt7E1w
oh3uBeR3RRvey6UGhb+VnGmvagYmnt9aZTrwCNpCJrwBjXA9fyCZ5/a4oPdgnWf6IWuxR+BsUGh6
cO9bLfZTxmD82Gppy+f52I+k9yYxz7tvR8ika1UUZKeSCbxtyivCcX14fw0eZJtZfCwp9DEeEaiM
yZBmIjq1aUy9VW8d5xRI6Y5P5lF1+84mTy2cpf9lDm6VqoLy0GOMi2opnsh0gDgaUyRXtlW8vH0c
eoTutACqz5OuVx5DcI5u6tSp/UIM2igt7y5Miyp45+qG1vY2gPGKev+EjJNpl9sQ0XYEG8bY1dyw
/7qBNxGrhX4CPnIwUcOtno80JinViHKHEes3kDIjyBbpN4SwkxyRQdJ8f9MQipiM0XnPCPdV2xpn
9eKuDB1f1JxUmgrRJIqSrPZuvhEUmr6m1c+1XLDUw3i4MlnO+IqmZKM4Srq+gB4IS02bLp9yS1Gn
zQMuHVZBx1knTPo0XTJuzYRI+W/b2YZN7udIEQEgpyDAYPAoajcZ6GbeBx2MIRTH+ehYb2vVmCZN
S2YmnmH4Dq/kxDPNTeRcdUrhNcLuMfxNdjP14Lm5SVd2yVD8NBsVnPy5pzZsQw5N07wu0S+a8ouf
THXs3uVs5mg0mF2rYToQD3RhCgl7h0a2yga3eZ69t5jPEY6FPUy6Y6aTvmLVzzFCP0eAeKZ2q3Gu
0BshQpBTC6JcbaxVprDhvpTEkLeuaGY/P9nAN1O7RAdxanjalG+HfQX286QhrMIURJ/OBiki1Q2Z
CfFOhWptg0OrcPR/1Y8UcIxCdQN9eA5urggyFEM1IO/YgZNTmKuzuVvANdek1ov4+w13XhYBxV1/
ZxNUuKwa2Z4xhZtg4tfiSMhA6XC1Und3cEAsrjdRe3IXBjKSN6LgApI3DtYqybjyFamaE33yY4UA
MkviV2lpLsX9ziJK7xCb79/BB40u3/4Qhyf1VuM0eOZf4bxu9n4b/rzzCeqRJAXPHVkGRcmyhDoE
Phnb53C1JYHyNQM74aNYQZQlXXaEDJqtuHvbR7oB7WTlKL/ZxR93EvxkeEXMYt9PxFKCMXjK69FZ
LqVhPLVjPkj6YTbzH1RZtfnZ4ap7kFIwSC0YeZ2SzyO3o/E8YAX75qP4E3Meah7hHdCMLw9ZfKYe
ukuDTVhLJ0Nbd0NAEpT2xn5DCGJ6Wdy2jHayIbixaEWhkKpSOHkoEYaVWSCd1yUl+1hfWxNBTWCV
jGuPJyiKaqbt+YlaVW9oyIirXzPm02NGwrANe7IjRtlyMZDtb90Tq2efQte6zrFNawXWhZOrDScY
BKUC91XpAznLWI4G3cP1A05mteSn7dW+dbMvvtzn5HW6Dtn+M/KRGjPcjjZKNqrv9IKK2yRNd5LJ
9+f4kWpW4FYSTtIZh2KFONsF2sNRfxr8lLziUK+gen02qPGxuPVBUvtTi6BLFO239RVX7vrFYBKs
ou9E6wB5eZHIbYwje6t7bn7blEEf1z2ZIK5JKzSOwIPHOLC6DkB7MMFUzdg8bjm9bVtYEcEm9rN5
MO7CMu/aXCujCzL7mstxSZDqzebAxH1lDHvHVWSz4GOs7P5AV18NDDMC8uUbhXk+klvqKMct9iVl
zjd/I44AKJSZZbh9Z5/6qn5iYBcO9EtGT+4ddIzPSS9OPvmaLS/afSOfRxxHKLXbZ33pknLFci15
SZhioyvSjL9lV2RmA1GAbocaNogkrqXhH2DCJgBoSdIdxAeybslTQGhmJeNd/m/VtHch7wZIN6Wy
T6jJsnlzXuuLmVWFl9web3y9USlwbznbGYYwoR0amFJEEh3+6IdLuy7yCFFQt0vW9tBvjr8qwI5S
RrvNo+CdcwRlJQpxdco9h0xvznwJDSIOn60KNfZC6woU+eR1oEoCaJDuyWjh7CUU3kkb0o1XF5dm
LNtNqq4/Y5HxoqGfmz8NLCVrHcyaGIuKzwmxPEAmAQ3WI6DoTr0XHsFioo0lVQGiNQhvaaFccAUJ
8gcerk9zebFfNmk7JOBo+ShsTnl+cmiQ7Y2FQXtuhGPsuYHL35X69ZkFWik8/ijS7E98XIxK8j0c
BxZ5H8v8ya2IWCCrRaH9K+LeDVERRZaikH1o7ksppsI8zNNWq47M9YaQR8a0baV1c8GP1rBpnpKL
oB7gEvar8s3zIUQXpayUsvbAiq4fXq0J0HKuL+acZBhVFUPR6u0BAwo3lytsZn1Ga/rBlqwjJ6iu
Vdwm5p81HQ/KB4ppniJKX45it0QmCZa2qu+LHejJn3+dxsxtOIQ1Qj+DC36BH53DgV7uim/yn+Ai
NgJa/bFFCBGW9yqrETQVsuxsmx2ngN+JK8syFIEaKIbAbbiAejReBkmO63ZHf/TMf47w5kqkxQDD
CzWMR6HIODFUHjkF7qqZg8BD2myifZxSl3Cz/Spm78GOBp0CKZVMGvVNKX5TdfWy5pNUqFVMuNbz
UGROujykZqGbYxPgZXZz6ijY+E8se87d2Ra0OMKwAEMxJCsnK4lXx4IrpB/hqWHcufgea9jKaahG
PtpDonZR6FqGrxzsCcGSrBHkUlMMJxNZtPGv/PFP5SHvGemc5tcAiaY2Km+gYB71tL6WoBE4wRmm
udGlGq0F9e085duI3Im/ljXHZVC+RqITVMapu76QQpaVix+qaL9937XlNWzbQsBelVXFfjRgkh9z
iNhS5FCWg39TxwF/9LwoNqjjbGols9MQjjgEufcTxZo9f17m8y1ingsLXbnxod3gArRQVgN1G0Zv
m3ozxcz8ttZ0hlZB66NNrjKVO8hyY7aUenOyZRB6ih/echmswtg2j2dCFOUVnZx0HNuSjaKGVppW
gtbnSUtNyf0sFDpQlK42jzetZ3psw0NMnNA+LwyYxg7aCAsWj0Z3Pry/Ibd3td2SkDsjB7TM0YS1
wgEtzf7hjMQVHWpryHOvu9BZL6yRDSvKViiIAlIAzIb5CGma1EpiCaC9h7wQuC5G/IxkahQOQfqY
Kq+KJ8QDMmibo6WqqVEv3L3F8XfkwoP2Jkt+D0KGpz7iHOUot5hmdALwD/u0/QlC/PVCXfBx9uWx
l2OT1SLxkV0l4J419X/8UVjLFzMBtc57RvIoy0LOMlUkD4dWZJHGYPkbvRjFnfx8NjPB3nRaJEKa
Q6AGwWC7KOizfGf+3hHSit5/TngAubvPyP+1x23q/ejAjAjUF2W1mgaw7j5O955TXr375/kGRYIc
AHFrsBioZTEyylpTlOsKH5V61pLRiswrdh5cR59fkPeLpgDvin0zYA9U6UdsKb4so0+mdV11y/P9
CByrbXSL9uhzFfB0IlahKzxV7zSL747uqMFiyvHo0hpqfFGO+LPeqPAsDYIemkpI/hk9HHumojCc
w8bUDScUJvLBE1Oc1iHSgXrJba+9IfGJ8CygApD8MNrIjyv7xYMGIfOnQdMp4XwKdMG8/gDxVryH
TyEygqBcJO1Yd3Pwh9J+jRwlh5MTjwqEzvnBrz1AN24o29qjXO++cytuevUB5HQX/SnL1ziXgRYW
Vg2xIZZjO6+nVx88xeTaQ6hi43uWoPprH7Asnu8GVB0VCPsn0Zy1Lo/9aR5KNkC3OjF5XAuLyBfY
xFenypF9Ub1KQClrjKHlYYEbjBpWg+DIiNUO5dTXVcc681/6mVrdV1dtd7tWHEZMUn62Fmz3d7zA
k7t7TxQsV4ZDMUpGBBTgD8tUv10fCGuOMalTtfXn3txs2E06QHeSPDdL8d0eSe6h1duV1HTn2Lbb
rt5fqs1XD/BQ6XXTkw5rEf4nNQdu40pJ8iPAkWbxhm3RDh0c3Ban4yLm+Nueu7zqmKa+TpHVaaIO
jQDhjrzGpPsdPCcmtKU8sMcoJAKu36IVc0zRv7btiqt5cQyj1nNqbDhfSQ4Z5epqhGnBEBRRkFKQ
ZdBr+8CSzVngEf58QjA1lVtMtjOwohClgLAW/FZVeXanwPpQYz2HVc3juudjX9m57t7tKwWJfrAR
utQCDhIXCg+8qnUFO1TjheSCHP9/VpPt3QVWmeDmvHxyFCVkur0RZ74+ifnFACnwWGbzm1pkm0KP
h1e2H/PZ4Q2fKVM0ZeGBtWSVQQ6ZNmnTMez4sCrGeK8WzUGw3Bi6t020+sMixiJpnRzS+x5eYXwt
EnmZXjvw0vlaWLqVyc+qvdCCK6VJLM+D+cwsN9BlSk9mYxR8LgW2cPvkfkUEap7VIxTi/OMvIVOh
gy0KPxIUI49+gKXu9AaLDEdbKBCzDEoAoOr4S0/g8WQ95yY3wT/nguOEawbaklwe1EyzncnJfKko
oTQB/spdm4SMcFKa+oDjg31BSjg/z7S3wNbeDPVYqWYEOpD1CmRFuSy7cu5q+CGeNeVWJg/UsdjV
CFeFdCq5Va4by4dpxfinzLXOGgCdKoCcbZjUFxJ10ieTSfzpD4IdoTDxdJUvna/tzAAaTCZQCPFw
QXznvCi+ikGWVKDiwQW6u48fOEg2dM5IkYlfuJ6BJbO4xJZfMQwzLcqTGC2yyldS3XK+xw6XouJz
gV/Y2ud30914kr0IgnX7nN28mTnmppWotLqNoqNe7D1HZ1L9JHxdDDgJ8QrD2IZlRwZ8C5j8vtFi
0qC87TOoZ1lZXuaSAxhj7QAzeX6RRCHTV+dObMu8tg99ZYNuz0mGw/J4Nl1+9yjkMvnWjPEQ0jEs
tRO/ZisDVVLES1uPGSjCCnD9MSuofc6JokvMB6zWK2swb4TZMeog7kqv91pcdVuYqmc/+gr7R9BG
MiGU140bBN7szjZSN+Oqr8TCLPYwqztotBjt4e/eEeSm993IqRFvCBH10eXU4X/yTVFCGfxRzRNU
WmV6P2B/+b8GWaGNtqXUIPlctyXWyNAB6RPFg3Vf9ZBvQnctadbJtWaAdeWnv0SdWVcIX36fkrWk
Jf3PqCNPLmVtq/rpMJWgm8mE1udmeXZ1d7fp9aFzNsxuNjCsKzRXwMHh6nkKV1WklbbWSpDnW5WH
TFv0ifCUCenWe2kVwKWKSllF0KGKaLL3niCetvajWXw1xSx2Su/H4TULCd/Bf5RrSDct/8oPUoJR
Eq8nmf48Own4FVo2XckTHNOaGe1QDuEYY5Sd5UJkv1Z5+LIWvBscOV4d2kriIpsQ4t/T+taVKZFN
2QPU+BIq7bwRy+jYKFZNnaWN/CNY8Mu6QgxdBy6GvFIlYyQwmjWDPeo6yKs731HzCgLzSNAiqq8T
hB5LDD4uSGBinf1svfk0onSLOPi5V4YhyBo6hoEnTR81FozE8iYeHmO2ExC4yn3fq2CHTl/u36gf
vkAS1xEqPXJzIgChM43qyA4A6HwFLfpMp+qv8FZZA2VURuqtN/Y5YmKSEwaAg95V18NtR+esGKEv
r2xjvgKUes1anKPzXlGsbmtcyP088thfwGkMlc1uWRMIkYtleifgRxcZ0cd9GJQfuNuThCwBQQ1a
ulhAl2uq31BOimVmP9jviyqB9haUFbELlDL3EppbDs5MHYKo7dLMBJXgnZpwEPXjM5bTAXIMWX+/
rFWbzsuZ/qbXwaksxqFPClP2pNBrU9W6ZYRscF21V/sepsPxjdZvI1Zb6Pwqq+viqGe7rIicQjs7
eiQ3lJXgSDFQdhrPiGjFu0Y0DuITabPBgtG4rlZe5wMmxg7PXKxREHvT9/z2VMT1Ky4m5eoeYnkK
eGfOxmaXOQ7GOzIzk1IWwGAMyZmgxJxHmU8hRh2QsXq+73rS99E55CD4xlJiYghRcZqQUTxAnVd2
t8KMWjcyrAA7F55oWh/6gEfbnjEw0RzUcG7yKUNcDLJoJnMj70bxnU+wYhwonQRtsz8tQQGZ/3q+
BWb1qTzoKwXEZilGRtqpAPuQnNgPVKlwdr26UBv2JiiGtADz7ycy0KSJNB+n87ELo0mGiq2ClEPX
NKrnNOMTFpmVVMNGbk56h+T56eGq4QUFlxu5PY7+s2C6wC2E5JTajTlxTAKI90UR62iJDczNfoWF
RXwQjZxMvNbJHYJxPCtzTysGlta9kQP/wuJm/T6QqaevhK9pLsO8dBT3gUtYVYyHBKFYxn/jmyhs
XJfcre71qribQFbGdfpI5b1cxG8IbMlmmX23BeFZBWRIgGLncJd5ZCbFmLRwk3UCmrVAUs5/ZrLl
OSEyFhcBGSAskSNCdexp6x8DDRgi4Nn0l80zBp00eENDAr2jZGDzFRF3FEgTRO8WTvk+jETIdzn8
xpzmSvQr4mYRzvBcpGoSQsSUhlcFgAK5uvYFqgNruGkVuSOAKfDSmPTVj2H5GJIzKJIeqmNY3CrM
qjvmn/QL7pkqVsR6Gx6B64Tljb3KxfymZZ+GbjOBXIPDD976uquGxyJH3MqxS2yKRQIrzhfJaJFk
RHrk17tVU19QXBUfFbgknKWLq8T/WHLaW9aowYFHE7UdB3ytzyAlKAGi/3nCHK6Pl41Ute/wjsjN
oqDOmTzBKPrgUXslZ7Isstk4Kf6xZgKiuwQ+hrgLBlXgqvnRenApRJxHa3hboUq0H6v52zcxHtcj
GAMB4TEgiiL+PoGQ2MxMmXXP3tm1o65nOoxAO+TPrBzC+P96vbsMBQqB+I+dsBxbmwCBKrhLGqyb
6OEu1SFbKWeak8SzbkAkCsJ16+1L6pp89k0m49NbANWpbQE/kJt22m2oOqafpdF67Z7V1hFwcIw6
vYqdEECG20qtXpGahCdg7eu4nPOsawbFEa2mAacgoW1gkjiwP6rp+pSDGkgYRv9b5ndGOCA166Xh
hPoNZw+audtv1LF2nMFkA9GH/XzHLbEG1afwMr9D4kirZ4tYK9hFylpx/TyDHpBWqMRS9vRldXlX
1SDKWq1vxIfYk8Ih/8s/hOZVJBFRxxolIe0qfdSfbbAOieTyDtDzdGm4a7xp7oPljgXVH5BSRh2d
4sy2WDszEy4eQ7fIBk8Qm8T/aIG/wIojkxTnHRhiAlFHFxWK+8Z1cAVMIqvBYRs/IikqKEbZtFz/
yRa0tLN153ccLeU1lmRhSioDAAroLlSsYHunDVSv+Js/yvqPoCrRJz/wAukY1zgHMUND1gkAMD7n
/Clfa9PWWHd+4RFOd3L3k+aUj28vfhlVpoEJy/Ki1BezWXw4ok0Mt1g5ES9D2iYrEpO7bp8igC7s
9x/Nmzn/jb5dcZNWLOINmRgLph9bo+PD0NNoj3e0/xC6iWLycgDcg+kLp5LDfielJ5zJuIvaq2Mo
tSvdqi5x9UQSkdcPzLF3xrTEStAzb7s2W4IMUVOXvBYEewQZMb+VeOErCxvqvU/6M9tG+RDng1tp
7ipzTS70Fz+YvA6WP/4jFWNcDe5pqOrVLI8mFBws1P3RM+p85Wh35WcXj6jstfcomieH8ZniOTXY
9wnMoH/LuxRKTbUG4OBUO1IUA5qs4g8SpDzg4UJNyJvjiifz9iLn9KjXxx+FpYb5dv/65s61DR+J
WlK1bCHQgI4kPcdRSAxQxRyr8+XfT00UYbs3UWJ/yPi9evTAB3U6FkfYMpY7yu2MCQmxlX3jhWGA
om2ocltNLiIAggy6wgemi9gVPWncNDDdyeLlex/RpjEdsNyRpz73QXHC+bAIdkpbnLl3ns6ViW+T
kDKukvapmV5bAmuwKm/BHYVPMYuUVWV46wQn5q/7UzHOBBNNp4caG74pk/LYqewFM9f+adrsYudO
K+E3i0DsgyvYlL/S75qltZgjWIoeYvRlzyLa/L0fb7TZV10Xi5lSFMpVNUoqZ9e3A0AB9tEWeyzp
LqNjdrkjsi+ihhnE+nx0ElI4il4LHeG6m12cOn6jC2Hnhukp3iGjovGFSxuggKwagvV2QYq8MM1x
i1Ld1SuaJqxcvvAr3MEH0dbQDomhgTDbUoVGu1Ys0rFhaba1hH4yo29/OhIsbWe6h6L4Hq45KYW3
f9DFkRGvGAMHLPtCkpGRM49eOFJ5L+kTAZQ6jSQrFc4CLKoKCaR8WCOlqA3MjRRAGYONmWFwtK9B
QUXvXMS0OVSzWrESkZvHOmQX4AKuzcCQ4hq8zFEIZ7l0huBYb+4QgwW1GLK3dLtc069FiXncl3o8
kflfp0fyYLkNnbhN3JAnJ4iA6wYQOnARr6ocGbnpzAMt83PZ18an/hijUjK+Ue+/KHgZebdimz6s
aAtCIjiORIhsH/Bb4hkxzz02zuDVLkfhM2+neBodZD/+6qMpszE0spREHjCbrOwZIPjXLMrg6+Dk
Rmy5enP6/G/sQb3fOmL6Ki00b3d3UkEE15wmxL0HbBLeQmEQHBljTaZndQ7CfYSrcIYcKPTEAKBP
Vf9Kkges803V+nHCrp7RzqD8whQp1KBbNmR2lZPjDy6IZw/lMdC+zLsbBvkMyT5hDDKCqFadK4kb
PLHVX7OnGanhtVMIs06KNV6j3RIRxPpjf1o+rURkwF/IGfsNZ7wcVukrQSw583fopmf+derEYu3W
qWSYrHMG5lvEmED8GUB8gfHZtZt12zWLi+yVs0uVjsOKU5eSmJxzxEEn+Og50jP1mVKdHg5fw/hj
7nNXpvclQiNp23vmz4yTASO2ZgAed3IfofLhEA8tqHwwnoPxQPnk4+4UNURapUzka+oU2BNnjpxK
Zc9C7HfgSsm1n9ihSscVZ80R8GjWIl1iGVtfcr1IRz0geTu8gYNjhqUOD8BG24GTKzScN8gtr5JN
8wFg56TWndWVuG6qdQxwAZSPELXZsANyybQR7urg1FmCMHrYxxiKUkbiUOBYxkztqyyI3kbewqu4
F8fNx1UuYy6wh38O1tBef9T3HT46ho9O1wr4nT4vBqbtuZaHfln58j/YUOwm74s99v8YhSO35wYw
5faQX2gXCkQ4KWB7FNS2bV1EVdfVt3YqPI/ywMFYEcGf8YYSU8e74y9YLEFmONU4gW0OqWkhCn1a
VjG1xL1yd9e4/aXoto0+HdxY5evXUOfudnkvwM2OlWgrDkZFCkRrBtpi36mZ+ZRuHl1e3aVlu6Vs
ct/ymekWaViL8x00P1DpgDZvVrXmqPpb35cwtENFuyrYQWUy+2U7kwl4JsdVXNK3jM5uFnw4W9i3
CfLIkQLdyqmT5gKfCztT+05p+MDOkjsmMoxuhkGzrH/Q8/bTKUOfc/MfomycHzmzoo1yNPIECDQv
GoiTWEVolB0gMTqnYpv5hBTCXpAltk93FUiCVqrwklOXCk94dIEO4lGNGK3gXANAmACD4Pvb5SB9
QOTUJvX4dP2OtvPGnv2DHSAd2GSB0Yc8KsaXbprM1FT1VTNAGUdrTcErLYELPNKPxjwj1CBAuY2q
KhkW3S2kxcjydLoeEOXTBuPaWE2ARS1RcE/X2vu9WxRm+8fLahS6xB3kxeV9TwHV0T1GmCNhuBi3
9OEkwv3JJ2b7KN+Pljy9y7HsK5QOw1xf+JlJ9CSVog85ZjYfve8z/zXh4HUuR8qhO+CC5x4RIRXy
BBZxMiwTsgWDDK9XnY3tFAKRujXydVuNvTjj5l4vZEQ3og/xXaUOwH+YXr/AEocqtcijCJLwvj1+
K1xExrkYkWu/ah3JPhOJRQVoWMmZrC146G+3wGUhlsX+ukSOacUZR87cHyTnCNh6hTeKGxOvGteL
6+T9bBegIl6oEeRszqSLZJFNsK8BPuEUC2ga1Wbkk9AuPVzUCqDKbTR0ub9TpZT45iGAaEPar5+1
EClYw6h4N9y3kzow/qDvMgu52Et+bb9Nw8dI6y+XCNY7bu4I3MV6qaqf9ZcD/DofB58pfsIn/HrW
DcNz9vBmRmH1nP3+GZ30vtCKFfHGDEvfLeyzf9US1wmWI6a7JXlfkUXc7OwQ3wf+Wqk7sWYlaou8
UqzLc9vtokU8Nt7PMhCEsmj74pbkKXbM1O/hqWvkr8F1Bf6mMRJrcMoNtycVE9RjYE3WNy2F1Mh5
/u+gGC03Eo7fHD7G/x8cKCCrxLX4WuA4qWeVfuhcxS9rOUIEA+ayn7FsIMW2i3Pe/3kKHSz6Y3Ks
3oPAVbhkEliyMZutwur5jHhAmBnzUwtkqPU+9/wv3YBO1kKRDCmfY1D4BLH+qWpLujszalP8QzY8
dG30YZqsYFdg1nt8PUZ580d3B4aavugukDIqjwOVyjV8ZiNNY3zudwKMlsR+AmDik9J6FQUceIRL
aPQjyVAXsY6aRQwV/c4AQZnohdjyHGbHNMPGFcmqGjf13B2YJgAbKWshzbcOfJkNEALZiJ3Ts53A
Iv5IQDeNENhzKAv9iqV0U/j9WBzOrPCouyA2W+iTIeICpXKSUmJOUC8Uj6wyv6YY9bCChjvRfuZD
Hf3z5U4TjdugZVak1jOB8/iq0aAbVuFEiFvQPXqKlAkVBZW1fzOxXcaG6k5QHdHXNbY5qomPpizL
byBHsNMbiOVB0GqD7ORte5is0FS29BCKVAfoTD6gYe0BU8Tn+isvD85oAh2P+4Srtp/n5Hvy0rXq
+kJeWkdwrZA32mg0MV/lkFuQqNC1x1ymn7SLNr+GEo6r7aoUvZ90JlK+ccdXl6d8jPVAzzhZ1FNm
KOg2lhkZXfOoHJYRjiaHTrFCuYfs2q99yRipcRNrOOxOcY3aGZn32RbaulC/64yT+2X5owns90pi
tg7aTk4ZrJH6vmw7dePdDm4IrghYkvBQ6dlr3ECuA4h6ACQSOOHyASZT69hu/v0s5bYux7OsGpTC
urHkst6CpIxDoliKQ16Vd0YELiZaYvSoUltKxX5ntLVbQHzoYety4kPvKxLAcR3/tdU/nLFnZ59q
oiVYXHwr+mUkk+qfHMYLSr9tOmKZHOu7jwR/Az6YFSFgZBonWszwfjKmsf7qfwOP45Iu+JrujGaG
T1a52G0g/mfZzZYRgIHgICDUQBMzAgdAZZMRQBeT8mPfC0cEfFTMhwQhHAFnVkiCEZrGTEj6EL0r
KJnckDHhIso8uDx/xRfdXjum+ocydwr6ZHa/m4BZGmFmetF6SvbA2q3IL43kVmfe+aHmrgdbwCCP
2cnac4uuS6PyAQHqhoNo5HBJS6jDEk1yQT7vdE9htaGT+yOJ178fr7h5a8fVSP33HcV7M43yD8no
BR8+Jdf0+Bkd3FvTaPDs7qetBQY84Ah6ldKa7ZGLrSwbKZEmtNRbdquwpOpoCuLXr/RJby2VDvO3
JVTBqRmjDu4oQEu9ujJuxplKUc576U1Im5Ts6q/RW/0xn9UTnIplIeVZ9r6/LoW8JCEGAl3ksi9N
Vih0lbavAqF1rD/cxon5ocTM3lQpuJtLiN0sruwMxbZ5bX3Q+s4K6fLbPGacvKPaVp0Mv+HWgjI/
DdNOOfACN/6GQs/s0cy9KlffHiRLEVzBAGfBDOl6RclGsy+5tAfFkUAqvS91q6fE39VRrTIGHQHi
Y5Tr+iaG/jywkE4DlQMre1c5BytJKWbcN+OeCCOQBHYQzXEcssNwBm12IoKfKMxwZIZWlmfrXBuf
EAO8Sak/rfUPTqqIcnKjxeL880oYLnMh3TCihB9wQJafDH2koo7IyItkI+jMx6TSLTLTP1+1Fe35
VWrKqAwu8l030BtoSt7zma6jjHN/xg9ys2NfVSiw4WQ6llc1NYtZfOt76QPeuPcAV0wWb1kAxF/j
y2Zme1S0lfYODzKxFW510sWWos46RzRCPn7hhNwRUGaDZ2UCLud36yNtBzqHqoiU4S05X9o6Jyzw
UJR+qTkvtiBmIg30OLOgsgAIdgfjYJeUbiGw7FOJnQLl+bxi6pRaZBqbtUs7k2GOuwBxNWbyaFCf
PWCWyHFr5OrGm72UXBWKeoPndtQhZn3lNDdsHmcJOhZHqntsifMVELdwR3bl3LOtGZwB8ZeiXXQP
WV/V/PjjmvEmaopKiAhYUQl09croJjKn2L4jJS8tIAt6fAqaz0ZFKxKxOAD58UHLYA9uFtIu28en
SH5gHNaldlHhrbIiHxAu32RNu1OFgf+TAX053mUPVdxjuf7jTT7fH3cxWE+ADFMZ7pkrDf8Qq+yP
ALAz6/4YTdNV4DlapG42jJaOpL1Tfkl/cFh+krUAZSP4iaXeuAzZtCGRySEGkaRW/Ub9cSKSvk2K
rJdzMPVFaCbrCMHieotLJXdfGp7M7Eirht6GqkFhbjdejFgDiAIbdtfGls6FhUnxxBjXpL3Ch55C
jQWTZya3yJ1gp7csiXAe5K30tr8hioOKa7BAm3VH03JLg2ug7+P8S2pWPlrwDdbdGLRu7iEfBO7D
NBBnYCTWSnJUpYqVkMHNbgqnKt/VpFZAiD7XfgBp6no+dDNKnlPM0xfKJiSIqkG+TvsWzEBrj6mU
q9eRy3PS0JUSc6SBKRQwLbk57xbpL+/hyRbXOolbG5ZOFT0qz4bHKhrYDiAZi1/3J+GafOgwE0MT
cydhTHNN0wS+0rqxsKULMxaIg094aKVU0sFGfOUAzZZBOn8+VgKMRTK+kIv37Hcs+L0+3hbghq22
Im5BIAXlUpXr9+zOXQJqSvOSI1omJcV12uXN87XsSM3a1Nw6uV3V/5lFQpiYohAozs0wG8dShy/9
EvvW3Oe7f1fUPjfWylT7d/KP6WzjerhOTsCyDBOCyO8y/Wu501IxH4kQSpjB6EKbFD5z954ArWYC
ojPwMkgz1GZ7HrhXHl8txzqIH8W+/Dn4ykRIa+gYETPtULD+nHLAt8/LZXuwWOaIagLa6/G8yBEB
nocVvY5q0foBIIOHksWLJL4ALz3mSBhaNROzKW7R/NgymZx2wMBnNRzYlJI/J9+pE9lJU0hbpaNF
EfdaK79rYixChIuKIB0i+HkPVda4DzefibY43Wbbsf2S8V1zfm88dtcQL2nRT8KNAZLlmmc0MwAv
QAwTAEtb9Bmc4Nn6gslNissE9tDFUAS7qCKY82mDUgSLNo/dzAnMb3CUQmJwZkbxliC5hZdhBXKY
dnHrLzh2am6f4os07ek7H1WMzbmPyReGbx/OTAdl+u/G4gX2odhHJcRSL8qSj/EQk4OkfjPGSt2e
KkvLsv614U86KQ5Xb5FDlro76i/1Yku2OZs5p1Zd1+pX+Pe6rquIhsxqXm56gs5qjG6Tfw6447/m
f1WiYQYakdo/kbl15SeDRq2szqXxa7tbDZeRRTBlm5Nl8+zKwVBW4G+GFzAnbC2Iw/E3hjFFUoxT
yxFmCKeS1wqehOeJn6U/hqbS6L6BRurK4OnG7og2PCbEEInsUf/dRHzQPk+tIXNBSKtajEUQFwnz
KXI62QoLF/GTWWdC6XLQZJBjkmlKmBcU30BRljHXVf8QJhmjTsIsT8xKbJlnoMSdbLCD4VeJ8wZ1
7O+aL9M2Jv/N0tKdLnZag+jLSo1eiXeYyRXMVNKtW/6Clvg7LmB9xcimqJzFN+YamR2/nUqb/M2w
DF4ZwHnMGTAqcLOrSX11GbXQywCOEzUcjd0iUcMqo2Z5JRnsO5V9ROBfTF5DLsukGNy89pHpf/20
t0fU9w3qv3R0URSrsRa0kLgm3jfjtnG+qSnSMORIX0Ky5p5DL7nV68NH+4FonMIe9xIPyLvogN7U
uhM5TNKwHZorYMG6z7MoZwJFAB2NRThLy83xTQ5PERUH8CNYwFV5IPKW/DthfcK9H8iOHHv7MMq0
YTgUFEUZCG0e71DlvEAcwfDNy/EQS/fFP5glMofhuUwzIuLaLaNBJsiAE67Xo/jZFlwmb3Fm3VsP
wr2B93DSxqQrCmCwH5HjuBORn+O3z9+qFwNOy0FnnkU+LlpD+PJas9T76VLC82jXcL3TDdcB7XKB
e7K0fLlDQm+cnWXqy0t+sTWxfeAb4REt9kytWcxtjJMgoB+G2eZpW5Mu6rTvkAJ5huyBNs7a+A7p
hycoPWSGltMloOnIwD8qHZVFaXr+iDbP1rxGY9AEov48QWMMA6LVo2XF8MrpZ6uJ0Iil6ousZJu+
/cbwwySX5xOs0qnJSuGp0e/jJCoqKMB6AN2UXkQzFipMHpJxQVie1nDODCwa1F6Rwe4ML8zR8bJA
QXg4bHhXGDyby28G6TM/YyNvF08jcuaCi58Q2nSpwtOvKPPzKkaco0ZNFuuV/TXCyxcrgJvVWXRJ
j9vAiFDGWSwpExUKVnLAQ9oYvrh09cbgQdo0P06yB4T75537WkyMhC5+BAkbTJuz2ZSmgdoX88QQ
HDlC5P5z+U/d+d1iHhSoRvHaxv5Zrn7yYRHlutGLVzVnoOKPamSpmmb8oYNUsEqd14uPIsoj8uJE
+jLT++WwlJHNVa6PmIpfiVinT/wPwxl1Gn3gNo4fHVqb+DjycRcuKODXM5xJIgkNh3jeYZdIBfGG
499o4LWJ4J299G7HMTzj46mIXSS3y0O4aZGdRzcAikz5YLUuX4TAoCwJ45MqZGmGlu9o3A4RSu6C
RVSPXeTmJWIBNEa+yQyHk5x75l7vClOnS/iaGAVnc/RLKiRvJf4qjYgwt5WLQttZPgXuLI1l5/qd
fnbO0CgZTXy6QLpR2tw/tf8xFfxqAwow8o6wafDXSFvaaP2TcGmXB7P8Fs/tZFg7BncSaRBiJfgF
GSmU4tMM8bU+S61pjtNcytto503DTMMQw7H9IzdCLGkEyeo0l+sfjelFRHrrCjGDBl3Vzniu59ZK
8sbhMytaALBw1YLL3GX/0OCClHvpAQ+gAr8p9/87v1E6o+Yi4VdP0mxzrqSh41xPg4bt6ozVTxUT
g9BZuo/m8VnSzJbxaZb89bD+ZgL7t0BdpaSPTx4kR46mWzL9iLhZMqNWu0mWHDiorOjkcwdrkHyK
K03+YMKj1x0YUkQwAtJK+kBz/Y9ihV6BNPlEl3+ZVXhN/o1z8Ut6e/yTqSLAHFqNR+E5ldII2BPM
IT48oGeebfeCwHumkTuoEno+EupY86Rx31ZwV05KBxE46bo5Ppb/uggJc5t+bMVlXZFPV30dZY7m
i2+mAs+B01jQCBta0qwje/MTLRAJvc2vtHIrUE8NJs2Fh4lesVvvflWuCksA5vMvpRvAq/iGlRVG
61nSpNxs3UYz0Bgru4nej8zfc7TW3AiYcWF272PG7vtrOt2oV9CKOgRfUmAsnPAndomu+NBFhwsz
XNIIquIKEcftojvkVJ5WKDilhSjrK2xIvNQoiUqdwg7hegQMjY3xArpj3Wn+KjMVYukw9adrGpkl
rKW70WURiZcvzL0HMYJDoDEIqRW9CACbUFltKE5fR71ynUfy3rp/vBZvbOlqEnXX271sKOf6rZ6/
yCeZQhgpOhdJC46tTSjPLIOLtp8FLxmc/bwCY1UehEWXd4bNLQEwfbHOYx72cAkToYqSWq/wAOWP
cd6cy+40a2mdLcIbRGbinhhtEBqjV27bMTITblkcfMBbbetKg3DrphNLU4A4tk5DagOW0lZqqOdh
ZV8cE0hwtahaPcX30TIFAQFI6zNy3kMJNTOlbrIAqsK71H42TJ+U+atkXWtSK/7TwZMfFSPBBWSt
td4e6Ukj/z9GQSSw0zcHFq6gwl/Xuo1+OXbg1w9Y7zvd2l3te8HSfmOLsTIuLhYYpV1+EnbQBFry
6tynmiXyc+0Ha8MKgnpQLHymbMeOM6x975UN+KDhgx/YwRRZuGR+zOUyVVP+p/fm8e5qYSbD6lhh
Xe+hlaKmIER7vOhJYogLS7NzCpO9T8LqoJKbQduewbZrXkDJA3fzaZ+l92FUiV5dIekldUYdbI/J
r0EiRVbdS+eYwUhObLaWIH4qOyzMDUqB+sKaFxZfR3JYORu8S/7NBQw6Xkki8WCUj9TagUDQnmbi
cVEZRtLj/AgqoKsyNd8X5lNMTBFlVvhNUJyuFwHHM8RNd5b3qpm/P0XtVixmmymcsPx3VDWfZsYC
6q3gK55kOMNXfxNJx10GbPmv1dxOUC3qiAqh7/sKN3eNaTsQyajgbG5p3tOKhVJPdTyLDWnp01Qk
aBLfFjyFxjFqvzF2XjR2DaP025bvKWPcFQKdYaaCFUhpwWtfO42MteIUkc7ORcPDudHOPpSFihYg
HH6Vzx2TUJWgmb+oUXOexbewdPs/X4hrxRQ3+Riupsc8GjhCMEqls6NM76yFjGWT/ZNbPQtYqb14
j49r6aOnVCm3s4APVg9kukP2WVdx9Pts7Fpa8vLqXFH+W1QouU0lgvkUTVmUbNm9qm/onno8MUAu
pgVgW7LLhAPHmK/QSGade0jRWhRt4SLkqJq80P/qDgaJQ4lRP/4PKJqF0TPMXzHQDVdF+WbqOTfp
b5b11fiSkxd4YflDip28fPRyUGF8NV27/7t0Sj5CZyv+tZd436XXOeFNJ/NZi+8w6M04EukzG2FW
tgyaRgu2mYHcuDDJiv6SIjWxbEGC24lLuyehjbs6p2DsnzBQbPGkeUANjwnUmEdBBH3qfyAjCB3H
BkrGUp5gLo4zuosbaIRM8Pl+rEtA3z30T1P5TpO5MGoVJqTvDNjMof2lJUNa3Jl0OLVb7LsTYQxO
0JfdUgq3ims55haYa5zXzx1aLhkycCZpVD9re27k84F3qJwd9Xk0Y/6YP2L2JhzDUQVVZ/YMkGJa
Z7J/eAw6y3QYwykmJCys2/OEBSWY3P8OdutPaOCtWVH3QKAA2+/Fn4KdQoRs+NHGaYTcsYiVikEe
n9RJCTbyiysRHuYv4OnRxD6X63/JU8YAQD/KlvgOp9ptbvD5DdIX/c8SPhGPQOwoSQFifICyJc7t
U2Zxtg4M6T5QYUSJMZtRCCMnzE9mNBcpgfGZafgM4/sxFHdlDI9XFXgKhVGXfl7zJGmNv0gSThkT
VraZl+Qtz62qozvnFW0tmnO/fmKZlQZG8arFriNL2LZU1YvfnlwNW8vAcIB8QMvA/fTkYTtno3nN
LbkZ0BauckYILDqUO9JdkfSbbQrEbXjVcjcsic9VcLmpiFiiaV3/zoZONCClxOISuhejhNRjhm6a
mYMgTO8hiV9q9dMvKYW0gX1md8WPVjRvS3fDc5rYfY99M9yl9WgItSQMAEoy83MyhP5us9VVlDvz
SVrwlwEBTRnIHlNWkHutlZ9140yfUFLE9OCm8dnl/qH4lcToGjFTW0ZSiV10gQFgnFw5DkS/SLfm
dy0eNW1tWeebek0EFg9mQGIEmWKaYFFf5WTqvyLtKW5g38beJUAMaBCHq8IAmTinx0ltX2RhFU8v
F08voHscYS5/5KO+pZZkrczJsFmLTh/Hx+TDAEojpjsbfAmxzla/pXpVFewSSkxgUNeHGUrgUui4
2tz0FlCAb3nj/cXm72syZr+ncF7jgFJupg/pTDcythv0fJjkqgCC1Wn6SdpMakFfu0EtzZh13AUk
0M/Hw6V8dYRgdRt1oNYG1unRb6pEhmo4utbnNhRi1ZcOf/07TM9+bihL+sF5DXz7iiGNdlAUdCWr
YvVQDEn2l3F+B7ecupncRu6vyhEerf04M7AVtJUA3xKw//90WaKpssITcvDuPTQRXci/KjkM6dq5
q2wRlXZO46X2Onsv7Nd3j4NVKH47YfLJ+DWUriq+yrkiA4La7IbUrKBT8+MsTD/MFQl6OxSpM9Pd
tcGXZBn0QOYIkg6lG0t9QCYFeyisGpYiAf+z7ev7OUxXUIC2zxr8F1PnR6e91s/02xRtZT2duO5g
Vd5EBaS36BKSVUnpRUYeGDA1gD8G4OXR5DhXtyzIM+4S9Ao4wDpBUBQ2SG28GeInMI6JddY8oDkH
bBoKWvsv1ke6m9ZEOlfGk54pRX0yKALOOVqhzBw82QxbpAxuBGlrkUtienJrIu01jpS06WQvYOTM
eAHdhH5P2NpgKzVKVuKs0Qn3ZeUTdIwPvhffra4TA9m9CCmD6McbFLv+BE68nXLzg+2yU8dD/NUQ
nzdzM0Xo4+oqTY+9EYqDAD8CV1ewIacyW/0qFcBbi4Yh0uLrrMqE3RjtWh7d9kjqx2swmzqYwlnC
rcDk//preNXRBmmW++jj+J1SuB6aG5yLH9RyRsfqEzWN5FnaKiA4xK/UsmkG9HiYhbeHKiPEgT6f
cGMY7k8ZqLpeFAnJi286Rf5+5ACr0yz39596/c4RjzDYSOrZYY/I4pZ5PRi6PVomVCaHeTfcSi0N
Lx6AXY0qcBNW59oaebw90BCYq+vNr5KdwtAUJsxMBxCJjgSeIX6FdLyTJNoiN5sz+Lghf7aMHd3T
P7xY6YDYSqLsAD6uymHlC9Ro+BQkeaEKs56NHtNiJTa2kleulY0w9zL+vLykcqiuIFq9BXb+DGro
qV+r3REivGqvoPDUDiazC8ddUkuMbS68O4Gy5DabIm1CsErL0+QSiG/Kl3PxCXhzbSnRo0W+0y4F
BRZhKx9O3pASCdi5wslcwjr6s45T6NM+ZdoZlQhExevr8P8MZm0mdTW0sWIML7ukcdsMOLOV07bS
4WgNCm4SuraTKB2qufwjV/D37o9Fp4CHLs6s5kjDKp2f0rwaIkIt7Q5EPb2HucoayNZ5Xi/hyrhw
JtmRY7LSPgTkyb0oEUh+q9TYjyRyPgoSnZ8xLKdx3tgGP2wPxO4k4JTyDwdHnN5BTbWaVLNH7B2J
1cpU/nyzakKPXk8muJl4W84bOY+uRbQUmNwKTQnA4OKdm0KuHeZLBj5Mm6sGDaom0ryIIGImrIYf
ycHa4/rqalBtF/S/jIifUmlOSzesf9KuJ3qmGpG1g0jU4ZBfEXEVQjfezlqecOUDtkQ3Xnv/3IAb
mKQN91jr892MxxDNG2VkNWeELZnaclyaguR3pUhraG7pQyTIQVI0vqHc3nWbcAMQJoRMBDgYQtAQ
0zlMyb2n8jE23OeGBivePSkbXjZIe5mWJl7mQTg3jBo5/smWLpA0Yciq5reZhkWPZskabzbUBLge
AsN7J7ZnOe8QJevTThN5PpsZyfbC06HIJ0ifB3P84YaqMCO4MFyRwXaGRnSwO7UFyJVd2ZFopLAP
vwrRVrVt7B4UWgBXeoUxzHW1omNrTK0uBVhi8FBzkKWzNbRQ9hOX7Uj6SgPKjiMfmH5oau93av7o
FH2NSZ8zArigTlviFqgdOoq+gt6DbbSA2lCNyfQIMLIr7XWiNEpnHhUV5zCFuQJ6RKgUxbnv+qz/
actc8N1UjZwXylWfGfbBEypSuuZwxJ1xbOyVSYb2lU+l5MCwhUMqv/A1ojs0AKADtpoypOvQbem6
7ABLW0d+hFW9gfiX6MtKxrQi23MbijKi4AClD4N1pSsFGcwNUyp4Zb8hWvo8IfVTkTDkfzEn2+MP
cgjjjflie0Krd21FDDuIjlFhr3Rrw6XsvfcXPl5a5ncKN9JMFsHvxupYY5SU1dN2nwF5AYJKdj5Q
rPHdDWHrPpJgM9EPYXKRTSII4vokbVPLDMUCXEUeIcXIqY3QF5IVcDUtpgIPgLHvnPDjVkb/a9O0
kkIm1s3vmalZG2XC3I1ojotU57xQPyAMcs3OnAgp/FM42BaLR3j09p9sJnLwMB2sMA5OruB372oq
e1MpHYmkBDeLRTMGQFPGlJ/5RR8Sl/guRPKl2nIFoSGvWFQNBEewyqAa2op5lTeSNHTiJernlHH6
1DQfQZvkDm907McKxvjjlsY1VV2z5v9iyqH/pIw949zBKxsbXRH8BfW76LJD7R3CNFg3aYmiSlY4
NpeWEZY+kqi5A8FvnTWJMh3ZpNZjCOpswSZvGgFXwOOJ8k9C0nUBOPY+J9Fnkt1RsDxxiNH7FOKA
CwHshyOmqhNKoBjCUcN5xqTIDAhgjoOkBhG5f3OEWTfNH32byLX+oHkQjSvVxLfCwpNhr//YDUat
6G/8MfK8Fe7MmXI1R75ufKe1WzxQOuZQdaOdOG8ESHRL7qJB8msp/oLxwkOjDo0lfD6xo2v4aDxi
1nycEDIxaWQSXJIL/RmELUNJAP8485InikouLDUnsWosKdd6eQrAjCaEca3A0cE3Yud01pjxqG/G
T2nnxqxKCuvhypoHlaRpyaAtnMisa8pm+YJ3CKnS6BpV/5CYC6XswKS9hd0ShJFx6tk9VOVUxDfg
oUvhrDJml6A5hP+6uP+N2mvMlB5+XhVSfNzatKHPGno3tYddigO4+wQUiKH1muvaj9NtYc4xe3+u
VrgR1AgikQhrsggvLlhymB1SjgmJNyKz1KzjaQppjgr+u+xRR0wVhRJ8NkqrBh8PaFg/tssCOjYb
2RBXxwtXyZB2Do/+nleEAaOHfXfSbYdjg9DFFRmbiacJVVK3mP+rDF6acn6B8tW83mgNQrBh0mzV
VLkGywxmpNhSxelCCXjF+QlPf/qMXt8O6AaVRwfmIhuSG8DsnkROKqEXAW75AYc+nL3lLbuM2whL
NaUUMGYcpOyX1z6UMrhMjUTT0EOMk2crzHXVplzFE8Xq8L+mAqbe7BeFwVBVGXY01/45WHsVQeWh
L0U7qpWcFJIcsiD0HPdU68iD5R+1xpCi5k4qzcak7dRjWMmTJ5eFbT9MVfD3B2q9o4jbW/xfWMeS
SoNJ7rVbyNie/F0J7D9/OQ1RNuGJwTwa7d1x6nnO/c35zKjt62DteNzUQPYJQ57YS3lbtKW4PV+m
MdXOn3KNEWKjLXWs+c+KagfD+Tfg/7DrNGSvPTDJMGYs+p1EVsJatMb549lX2AekXC/VYEeP+onv
e/0PQT2MNoqtFIo6MpIRnB22tuztFyD6v8mWxUpE8E3QzYTXT1TJ1mxqWeZguMR0SE9gbspwngwM
LKK+TtE4wqkfAeO1K08fS4MORsEracmEWz0TcRQXne1IBYwaO8hePyxEwPFGI7RnHnrNiVvODFb2
QMbTTsb532kmt+oUP4ICszwtfHVKv465cT4ydGSlaKDDtxkehhcKbgWq7gd6Wca1zCZ/eDd0AyVO
OLiESPgJjYq5XUXD9nn3Mq7vEaIMf3aIGjRwYKq96zaVNOcyd1xkLqTOHbbFtrFXKVwenhHfN2yE
8s2yhan5XNwXebdcL2BdTh5AMmv662WnkxWRKjOKqebtkw94vrp7+PLa8ANzSo6RPzKJJS0BskbK
LNn8NjcXdUst8n7TegA0W7Y7bf/idFcD/ZhOdrzTti+GtCy+l1jaijNV3WvOFYz46xwvjxE8uxfu
1cjLFIPEVtUbfxkiFcFqhbXK3yz/2P3dvyuibrBw2wi6jzpxeTiw9oO/yD4vJj7+U+RATZzqxMCa
vU4ZKJIAYRkMSKL486gMdwds6P5Kz12KvtPqDb8w30WAAvlCLXPDQwv6T4YOeBsOdKK9nRDB25Fr
bQ9dfFxuUSETeFJ1nrWbB6l4WcwLPvOEWpy3y+Hawkih2av7AjM7lgUMLWw6I9taBdPAuYumtPCT
AG0FOc18pemRZgV9MNkrc/SYzYy/A+nv3NaZDDckimYQzCxohZdI5+ODZdf5iQZUz1jn197jbxiq
OnVjtxECCVw/x9N9hDdKlyTDy929wwEduYOM2XXnyyB/FpMTd3DSAiuwqg29dtLbbsdf7Odai763
9Te1hxwT+1sEBz9ZHvLTNB0PpxwTOPpRJA3wOleI/sXS6OFC15xoFfsQSMWnOTdKziq+2gg+FS4S
6GBgLUY1L7O7Og6Xo7Se0Dmu8290u3NogEbf11Yr0xRoDkQbYDTGuB7Ov0GpReAKUxlr7m3oD1oQ
QAqQpyCTi6jioba7zcfutryNAPyJw8AbkvIDVUf140wJqsnWkmAv0TGqclIo6WibmlfEQi/m9Gjx
Jk67AwleEmKB7o2sVJGf8J3oju3iE28gwcUbCGdN0gdC5s36cfSOc0x9gWDK/1mwkwc5W6+SNLS9
4E9PJDFy5YdkTrhO2rUi04brANZK3cdNu0yObIieFRNhPsjCE6IWhldE6644iD+POGQl2P4OrqT1
IwJ3Kq4I2AN1NKA67AHV4g+EzmS2XcnSSooLsXqgKvV61N95h2Rd5asqTaY8MAVN1RQvLp/Ov6i0
egJ4W2OvT8DqdReQsUQ/K6fua7z8BkvsgdEQtSoehIp5UwTYtm3Y9hYCXPVAAF1Kt/F3V01zNa4G
ru8d4H1ETWPV2E7w2W8zWODXHNzbItVQTHbp2OYcgBJa6pa/6g7UhIVPUu86SMkahW6F+DY+m2NQ
2Q2hE25xgjpL8KHjTwe/5mZ0L+9GsvF4uL5Dd5McpCKGKP0Gkz7o/QjU5JLByf+n6fitkICZ5Cu7
SChaZkeUBbthhI2NeMgMqD98LrD/5TuUearog+V2neqTIeQBYNBfwH7+lauzGGOC9hkJeGcD2VFR
rZIihft6TVIXyHs6SWi5qM9CppTwIJdwNTNKO6rubApV/w0JwpsOCZbdS8rEUacvUH37+737DKgq
seaZIQUmFugRFfmsfQ2LEnkILeH/my+uh03cAzxpIT04JAyoCYkOU4OioKRvxxvDsoJmj3Hh3NGE
sV9rRukOfC91Fl2FvtV9gjODNLJtVU9UmaWN+TLzdL6eqz5MnCQZJiORJcsJ+PTM+eLkLp0aYQ+b
T936O90Xk1ctn49ECP7GGlkHpwpFLyFlzc+98ov3fsv67+XZ91xMAklWd0G0PsDpUOYMMBiFRN3u
QcshtznjtcNMus3KAGcQWuGNvkhzvNQY2hNDg068ld0xy5bLSoY5hqftAoNJd74ucS32878pntBt
pj+G3NJTYFitNzeUKSryExiAT7GoJq84vvI8A+ZIteHw9c7xDt7Z9489UPDG44WDPd6Q6DETlv03
M/2eqCEPmb268EJQB8Dqqz1qKxNptpMdS48+s5oiOUKxTq1VWxtsBNewMw1xRovSQES7rLjTePWq
2fvWbMBm74J/E05IpyZ84cHmcSWwPB2KUaGG4WkKwqpdwoY41vmGvgUDbjJAYahFpCJZ4RZwmH7e
0mNiU4cBs7v6D86RkDmHYNSuOfcj7XFKfjjeZT5W4Cv0jEgbK/dNNLL7AqMcY44Vlf8ZiDJxHAo6
e95NKhEbjxYxRSUz/DyQ6Onva8PBi5tNbSufXRIps+wKZjcts7CnTNY/XTUmCnIdEm9n5Xj2Zb15
eQpgZTqfQJVlpfcd/aRLzHuOiIwEidPMyJ9wYSniT+rScvPmB/NGp6ZLLT5TJyL+R7/ZX/OPltT1
b5vQvdi0CPZw98+R+c45XUfDO9rByR31jnmqWmfIZm+tedWP5Cf+1WEoSbzn+z6lz+RAwDPsV02B
vN8OJ6bzOUpKfOkE1YTdUPLAe06ANyC6wCoOJBil7/1FaIRu782PLIC//RlyCPVBUdDn5C95wPtX
5/N82RZnm36+EBIO++wLisJReH4kDyuqRJ2jX/CTaj6lao9RC09lLMcZZkjK1KbJRET/mcreO7HP
EtNIUPeEloukPV72TecluVdPutGOgKmYgmQytCYNZrIWXCHlwU7TCG7nU4eG5fCAVmhBNGbYKiOs
tqxUksAb8L1Z3Xln/w0QH4a3XKwMt4yJeLp4dehfiASAfeDfPcchiPCEtPTO+87KIUUbxJSmiusd
fdczUTskPFqVrka7NwbIG8rD2RtoV8xyEwixJ0w+wdwVcfHFdGTpq+CnViCIH1BjBtDySrvM+YtU
wjx3zMTdaEJDRNQPAQ7tdiU+EIZzjLxHa7vcsXaT4lR/YNuzEf/KPQD3YG4BdiZQd5E5Eseeegvb
P8KB/xX+h40bL6339oE4gpVmdciy25zPYT9rAbJaDt6WYhoj6tZ3va7CxTFrJ2VDtu48Dlaop5zU
LPr5YPsTIEJdNpz1jt2rwcxxuPmbHXy1mK8xD59xryCfsySSXSd49vLEgPnlyU6NlLCXd8qFZPhg
jzeVIBnZ49LIKHg0SMsS64nHs8I5yUSczGIdXdGbgZble/oIQzFnLck68rUOVGVqGci0S9gz7ViB
8BgSrfvMNShrP3xO+9/99oa5PnWY28VOrxXy/0oI5lSKneCw4w051zd85P3pKVvoeRkhMjt4kkBa
YNCwnjuyWCLi/LLY+myBDSO/uT1TC19Dlz71f8bZydBc9vOpoErDPigyvZxQT+iDkk7ULP6pHqp0
VEHgakcP2mhfZwBvhc3FnEjioMAOppbYwmJfS8V3HrAMriXtyZZdqvfWA49e2nkApF33OKo4A4ly
OyvktVhGp/zE+1ayttMWB935EvrPT0W3Vn0llQQmx0nV9Kk58t/qqaQz/4DEpJa9OQ3BonLhvRnm
yOLZzeMUx4X/dHE2sgRQg6q7Ryjg22dOoSP44d4izXanhs8w6kAASpx2oYNUtgjw+9iRi8OnQGYs
mzIhggywmeuvA92kP3W2XkjGTkr9Y4L9jPguHWuzdBTWDCnfoWfqrVg8H6NNpBPT20yoRICChyQO
qhj5BFaTM/DycU8nuzvrrGzpeF8N5zs6b4MoijKX5xZSKYe5yjmJkIhp+PgL+XPeXS7ABBAZEyAQ
eul57IPgPFymKatogPETlP/HV/DHSPuL4CamSgKbJm50iuep/MYXY+pIqPnn6QXSJT+mCqXHGA1K
Z4hKc+yRc9M7DThrBzG++UHOOMI/u3qwxRZB6aa2E3M9U8G93IYNh8wdb0OpLlnVLVTLONB6g0AF
IGr2HZS64vyqkWJ7fipj4LIh8HvuyH14f8mk6r7E52XtpzX0D9gVWc5J+AHMJd0EiWjPKNoFnSB7
7tiz26oIvXZm6DwUtzOkbQrGs/ThypE/ka1t9+wSc7fMOGe4RFHZh4/hluUVe25+RcKw/1o8Uir0
WqBySTSlnaYijyRjLWsbFPn1xMiS8gMPN8HSIa2j/g+DSNEOvhJQJnEVOwsXVafeMJ4MnScbT3sd
XGQril11x9GyfNrVKv/L2YGt4cF30HlNqG2pggVtbjeCf99YHfRZQbjl1UreyQ4BVUXTOSbn+aVo
wjXD8i5aESxwts8Sl6w/eajU5xidOOpwtmh4u+OLI399drT6nif0BujY2soOy3252dE0JV3J9cFd
3CJESkECuHfR+II2qoric+jjIW1B4dXSVBAsVDH/5Rk3VqzO4nQgxH4LdhZMd33/G6VRgn1knXmB
wlgLOzmem4Gh3MbJaRw8fwQWHFgkkDPeZ63x4B1RtK1SJQWD2D8hHbh7PbnwbQQNDyHmPPdzITgf
6wMuzzwPH5LAjNX6XcXN4q3E1nwpBin3Zxc0+IF7IFmI6fhwKgbb5t5FTmIX49BSh5vtNtgK+HkG
FHB8qA+seLjFKOJ7+g++gYVY5yvZwTQM6nw66Dlc92PT5/+pWdvvYuGjFJPgc4JZ9d7gkePH2uDP
H+dWWE4XVX/i9WuZvc1lIE9doZS4TkLnsecyq4YBPA44+m9vJ50pRVEUdS3chi4SRqteTqPEAGSB
eeRaorfPtw+GjdyR5H+XkyvBY1X1IXrVEOXuwVSVJTeyf6KuPYyiviiLeggz+kRs1NG4NDm5jbxk
bEZZh63X0IiZMhYnjZU+w8kThvcNiGUFWmZBHsb8weiyqFFIQ77qj/V5tsQR6EK7Jx5w2rKKh6qC
yS/Ff54R+9fQIgwy5RqOIwnv2xD9BuyPMcCVoCjG+mi5q8T5GmO4cFkZun0OheopYZSJoDuNrwGZ
JDd+s7klGUxw9fJr6UqJF3OA5Ny800MRyQ5QflWpbyGKag97pqGo7K3L5+pXq7SVIvtERUFt0Qz+
6+8oqroII1P37bGt5RyxMsO4GjbaykN3uDpxzOu4n+r1Vceb6JxOI4jd1p9R+U7mLAlyM9xXIGDU
O8fKel9sQbhP7ChPJEjViiU4PLgPSgEhz3iKkojgOzAmWS0ra4YJC25e192SuISbTtEf6CDf2YAx
TfFTIWnM7o89qRWyE0dl1CTtr7ci3QvoarGpiP1guAu8po+oLcAxGPJyjS9vqfsFYNuw79hwy+Ui
7tU2NbKaoTS5hIJ8Uity1E4R3LmnY72jm89Uf8qvSXboi/vts/GrrtMu/+y02ipl+bZURXDKtsuP
ljazk+tFWOEbwhpLpxoUwh6ZugVfP7NBcvPfhUv0wNxO6Z52Pk4tuvIZuGDdPP9pJlmcWHUROUCa
XaBEoGWm4K3SIpcF1R7UUibCa/8tY+85MLmaFlc9ZA61Karn2Znv4y9dWkOnSmrfjtg5QSt4shtx
5y6knevkuYUWq1lktN05cCvSGroRgLbzbZziQnheJO+398jBuTWMa3xx8/pO8R4Lny+AYOJzFrno
rni/tlGQEYXzP+hUo2Ms5bapeEnqPeM4GaPZpOQC9azXTzUSa3D4GioE2ky08a9P15KwwT0sXXhK
lzuKfo516ltjJ6BO7kq3wyS+rp3pgMfuH4HCK0EBf0udHUTruC8IR4v7UhkocA4a0vxxx85uAqM3
63oXnA6Apc2JrOykXH/U/4luTy+0a/PRWzHEXCUqNBkORtu9iL8qltmu+v8RJiFjGySPrSLXmVdN
a0kgcIBOnPtvInciV9Q/CbgXSHDIMU6z6o/BpP+M/NatZXs73BqIHeFtp/7xcClIbE/1WR+Xi/uL
dkvrxqJjhPf0MdIBefiK9XWLxLucKJC9CWGKkS03Qrw0QAq2ULssC2SYsSoOTCdxSp8ODLnryHgf
2kDwC0fdOSIcvj5109YrTBaRlvrcG9JyrG+3QlpJUFFeJ8B+oCr25sjJTOnGxy+PeAuHzpIJmv4C
f4zgSrCZy6091gKNo1Swm47CE8JKT9SqB+nMRaD4cLgK28c3J+WLcVbViRgCSwmvREj8AsONQzwQ
RoheoR6H+jByqWIn250jY7I5QsrtVc0BLyo074P+M/MNvpAzf2LuhSLhj8SzM9N3woi+oMCV7V6b
y2Y9T1GfzsJy+/ro/bXS0fYgazKeLU9CcXzQiPZOZIvr45tRE+HWLY7CJRhNZOsr5UOtvQpr2kIS
OWDs2/iIfC/4U5DxmrYPz1++FJLC0tZGqpUreYHxUJWw+NnzJvw2+NmZKk06YUXZxEBMP+IbFIoK
yUUYnAUygJygRwxQAaCfAKrqs6ivgs6ty+iaxaDrdh1lO3WgzHvqB1H7mNFMn34sLP1XeqXidhuU
lJXpP66x8qtPoScTmST+LgLNhPMZBpBs7VkfIgOimruvnoiVh66myJwzAO4x60iJfXXpz7SdMne3
3wV+txCOMOboqsA1CTWtLXwu4M1+98ELhMG8H+sjYscfY94/yllDtPc+2l/qo94xgv5zAwaoZ1JP
CdRXkbpwlIw+vHzsUo2DSGieoORKapDbV6dEmNWx0q+lf/GidYT4CJFRI8uMTtxG/Wu5wpM2TRTY
brM9Ful08wbOtMYJIgH0DxZNP+bx5nO6uJlVIn1prtlnnbXdJbtr8TC8ooGipm14lkSyZeOXXQ6H
Qlc+X9jBK7gG0xDvOSjE3XNjq/3F6GXBtPmxXkMeaUjbxYPcgvtAbl8mGxZkHwMjmMl0qm8yL6QU
lDCMWPIUadEAE2l2DPlNroqqsmJNk1gbiI/Pez4JUodiBdS/je/wylCFHMeiEUpdn5J9m7OJygeg
nNlYePFLkES5L9mu9m3mCLnVh0+dMIZFXZm0FY5eQHe0WoWdgbANGOtax8754FH+lJLNbPpi95iV
RqKeuWhAcdmWYREz1yhjXicY5jAGJHg8a05mL8rbCIb8/Mbomfl2QMFq0evwIgjJ4/4k2j4zqwy8
Xl8OOClvQ3x4ZLRFGDYKHkrB19awr9hCtCSL6epWg68vQ8guGdWETKiaZXp9Z2RPfzRzPueUyfDb
K+P9slgSmcM1hPh3TUSaKiPDpjn8J79AY0okOfyAyFy1q+NFDYeQJ9RmwHrFRZIOrBcHLI8qkjIE
hRb66WLLXR3NuDWU1rieCaFYut9H127C+234jWvF5AViXod9mGEZdrfd/VrK1qb1UeUZ0VjqGkW9
bOSTPmyUO/HXtkDvHgy17eYfREVAKiRvG6WzK9668aN+T/LbZ+XJcGdVqyVGaTqXe67mHlQrm1bH
fB5jyMG3He6MATW9V50hHUlw/53BRfcZrgvJxu8iWp4XPKKPsnQbsouy1CbBo6Ocnt7BY2eTqXrH
A1/UBm0mNLrlY97KHTiZcIAChJ9NV9Jpa7vShrpOZRKeU9sCjTg9aeqQE99uOh3SpVMz67UZg/Rz
MhHAo85+m+jyfXx3kgwdjdCmAOV2hSs3EOfBRz6VEQvrwCZPELUTQIcKKZikv0CBUue2sA0sOyNl
k7s+mOTk+KCbSORT0U4HYbhByGNAMFrlH0lO2mnXT3Oe5YurjMOa9fGDrSNwm++OSW6RH3r9Rh8V
JoLoWYO8RA/pC23ANnCuqAdcugbYoBIm9n3vz/RRnJt7zr2MURavjjz4nplIRou52Y+BmfKCK4Hv
aFezmb8v7RzxOGLGxGKbbcz7l4f6dFDPYb0fMtdu/BJckY8mTtvnMerMzrtDAdQ8sfm9WvRfSY0H
xt9CDKsZc+QwRU4A3uwFnEmytyN5RRL1NW9Krtpx3NON7MUHVbM99rbRyKBCT28AYcWmwDG9YMYy
2cbWWHR7fX8kUxJkxugUBWDYxphrM/ibROrwZAKspvOdUHCAE5AGJXq0AM+MBauyoJT/h7WO/OyV
6RZza3Ofe6sP7qPLPwMCEf3ivLFShOUjL6GzevVMQAEC5L0ryGJ1bNKQhiUH8/Gybxe5PS1+h7e0
DKLaiIqYkmifIODmIcyOMz4xXgv/QvpsokupuWRO1/ffWrQcc1z6tKHRt9XXJB+9IwNORMhdEIeG
KFYccOj+OIUAk8ye1mFgi8Cq5tn2bvNivOx3byI3fJHaLd8XNnr2HoZ/f6cekfGklwqc84rS70Id
M2oxiSnTvHaNVuZIXAuWS3PTW62xDY5mNtV1VZ9i7axuqS3A7hu4QY8XRG4xsCtEdI76OD31rPRQ
z/Hn8TzeJBblrYIqQgBy29qB0DeINZ0jYK5GT3fg9BjIUCX2/wxfwSrz7ovbYroEi8ugJE/hs+tB
pl/CMF7ASm7KpvYdacM222SY6KGRFAbW0VgB+cmD2yhRS6/7oimQz8LWVf0cwhkb3WWhIydHA/AD
2SdKsxrJU8S4e8FdTmJwiXP6f6NbCP27VfGgiydPEi3u3YS3rouveopS+0nwpRArHxdPX5np72jU
uG02c57wCSVBr41+kS4jxV5lyNMIDaSAXX8ZU/8MrdvVvpCdbtUBW9x7Nm3TkJ/WpTY85rIdfYk0
akrUMlZwYlKTyMaddyHcxfnILV6MRDEKTkYG7IQX/Ed+y6z++EBOlZ1Y4g+28HJEcoBvAYqM3gDh
XXqPz0mBhsLkrmL8QPSN2crmnJhnmzuUJemPzJ7uZnQCmX4xTmRYf0YAJsf+9yjH/4Ioge3zw+KP
UBTUuS5+/ZuZzHO4wM5LfFmGkvEpE1exoPKGcEQWI6tJgFpNBC9tvXq3cfg9sIdHCWeu2SsxBQeO
JCYgo14RfzUsCVyTdZ7Lg9KMsE5VArc+dUl5E2cx3U1VdN15ToW3DDQlx9TUe0NKgsj4zTfhqYqn
jMkPp+APvyxcWPIa8a6SQFyhGRCP+Oe4p7x4KE5iGiPzg/0yVGMsquzbb5t+YMQR/yE8cNnPPjRZ
TpfUPOJIgDKTmPJJQAZXoCtHE5mTl6+Zu3wAVMNio3X0C0IOwd2SXsgb9RHK7TDik35NF7ZKkv9d
tctVcx/wtiVDiRZ/SkQ0Jre5PQci3p4DFkvorhwKHZHnf5nbG1/gjtX/vusY6LxJXVOCDq9Q32xh
MiunZjSFY+j+BTb6/k5xXsGcdZxS7ahMblpBW60B0fbupVW0o+YpmjXXdATWKJ59qtXvfjgIhXig
4D60EeBhTWCDKImnlXMnB7g0NirB/YH2pdZ9x9tNTp/6znNkMqtk4GysX5tTfbcVi4Ul/5y7hIpX
+dNwtR2rxSxADztjdx7/+baM2oTFDgpJQbGl5EeSzV09Hb2wFCwBhtDwKQQQYDf7IkWcZRwVO6MR
bWsqfieg7ExzKT36uS7pmltKVXJM5Dx8DOxqu5sKYFDZyJ/0G8ViDlatOJu+NGtchTIdchStPx3Q
7m2dFwuLR+WPhdQhzgZRgS1eSnLaVjyDU/KPboJBTmPBm7sPpwf/XpDZ6pmhi+zDPxtna02c0foj
0P2EwCm8fgAR8S5V/MpRTGRWCPXcy11K3DpcFmKiKZmd1krNyNPH1tpZGSEnW+EjS6TuWV5XJu2P
l/L38kPzDavjWvn3cMox4CSyStcHhPKV8j27dHPeVxo5vt2HEHBM0m8kwv2BcahH+S2NiyHbcMr7
PQNd58L9rxkwiwZs5VJEXWmmcey7H5gCqiAemyd/3eskxT6QU4VfcBC1xa5KBO1LQrpozSq7aNYj
/zckUuk5tXXQQCHWcHCgIvl/f9/V93IHYtbe4PpHXuccal3R+fGeFR70hl0FFy5jLKu/2y+oh2fO
ABIWkf/hnbRDMBMX5BPC2ddjG4uIdUBXx9GTwDWjDc8qKsZYMZxrEsLQSMEWbtFCHyI3DgzEXTyC
n5jux2YgsVZA/SPudqvh9Jkydd4PA8XUlNPxKgm7DfENb7cSRjdf5Gc5wERNqqEO+UPvdIoNGeAY
ZlD+XFawRbfi04utI8k2YJa/js2b44t+Q7Zzza2EHjjcCCirsZj9VN4v+XALeZjN/416ZX+B9BlZ
/wusyFlJOMPWQIQBDsW13JbhfbRWk2IoDkk6Ks7JqBFnXPL19Cg3Y50oauDTYb7pEPlIWxHirpIf
YrjtTfqk3hwnXbedlJ8d0Ak/25mBU2Q5jYjjbw9L8pbFy6l6Vr6hqbIds/grjJtyRNooML6yDa/+
2dnbGae+es/el6YuFg9B3KELLy55CgmR4cHDl6pGQcvOaNBwcqQpQS/wUjpb0VbCT7eddPOsRwCk
cqzpck1zyJwbAOctEahpslacx+E1O8OKN3ZUXrUHh/IgkFW3DAmfYHBHOFOyLXuI7XZ/SXO1KOqP
KKPmxzs/ocMQux17kLL32SIJpDPllfoNWqk8PK5PUy47rOhc4BFRgVBIH3m+IRKTKoVgqR8jdQ4V
1nAuf/UI7v0R3MTEa0+7ybyZiBMY0PXGpB6ZELLRUis3llfuBvpVR5zdtD/TeK5NavTEnESYFFPL
Q8in69eN+Ct58vlTwM3LWh/CIcPYWv+k/Rl4FoY1RQ4hgG3OvPAMLdF0RkJvL7QUqW89l2kde5qx
39CLHmTZl3CcS6vxkNzFDa6+nLfi3SkQSjNG+gR6G1OqMYhKs5Ara0YEmRCJGthaJhROzzxB1oNS
XDFEVkKLpuEryVeEviBfBU/OW6mDNgGzzInm90p/Jy9FTwrM47VvUMp5p1GHiO8RHCt1t9NbSw6X
jvV9VQ1/C6pFH+6fd52CSC7NFJqDIi0B6mSpIK7M6Haw/LTU/NmLTFPDlxSuB/AJBdnvIdrzu3bm
ZnUekuhkxX3ElFqlpVOpxXULj3INSLyk4NDJn5jPLCsHnIaPum20lD/IRDUG+jvPgg8bK2i2h71Q
S+FLeMRLKfNPljC4lkoJg4DKayS8UVmU0a3hmi/laDysGJiNawXB/Sspcwqzh7Jkm+i/fjKaSt6L
UrqwsZnFKB4gGxCdUj+iEBFv11ZbKDw2J2BxCCjd8zpFPAwsJ/Fn6MQg5L/zNWnjdbOM/M2mw7C/
CGEoHbJJcx9klSwoTjACoh/NAa4H9NNxkQnRsfpV0a7mOW5HT4r527p01VPvUiZCZzh7vuKfNsiG
CszKTZnB29WRZcwwvYObiwZI7yyEL497aRHX67b9Ij9V0fD6AzwDgGmw/pH84FkCsoNfJARvCgoa
I1X42CP6rLNgJbE37Io4WR8h2O+1PNreauj49WGHTgk9tX+lSthmsTm+tfbtknPpP0jVI5uD5Aoy
CDDkmCai0CuvaU4YBc3w3S8KYPqMtR0o7QL1+vxatN1xfTfbZj0i+ZoknuZq4k46B0roLySHlU3T
JMmKFiVmJ8BTwmISEcTppcuj5QBUKLXD1vSfbi0RoGnraQunlOQ+3HA6wR3kRH0Qh7e0HXKnS2eu
OmglWXUg2DkJ77jG0ZkLDgZz2/ZBINlQvmrt9aZxkcABFRZR3xzQ+1GssZmBTiLSAa16TVagoQbI
/Xf9jUNNVhX2KQ+kB9osyYUXp490efpmZFmDZHmmO6Z7xZx6lENwEv8oAt2c1vicB6iNFS7/Kcg9
N0CR8I+bPcJUR6Ha+ErDfiADHbKmKu2qOh10L9WvTxDw37hzyG2dfBiXB3IvS6N7mLD2ixQhMt/t
SvTKbAm5sJG/WzRJkrlJiqNzegStehowqVayaFW8GqYQDynJUZZ8TcCAzfyl8Ftl8oWHw5FfNQ1x
g23hgPE8msXjqgc69/Q7lWzAOKVa4G5/fX7WP/Y4CCdgTQccqfkPSSdX9RyPQbQVagt90itY78eq
aDgY9PoFyEDOBglc81hqVm1v7RQLaZ0zh249kjSGwpmF5Z23/JstPmKHTASswakh+1vwGCkzaFT1
9zRaCyZ1982EvvOQvxq1zUzUek7uY0hI9/7xXquN2tEpfBlGlCcuN+zSlmKfMeeiRL10jeG5m6/K
xW4XhO+gtIrfU0GVWgLq/gqAD6THKIaQ32tfGbsNnQnUzrkiOj5zHOQh10IYIJOW2+fMMPsINrQO
9GPde/knHQSW/OP/wRgePKUNAuMG+zcBOzzLsyXD71+BBBPi3gKhW9JYjnXDbCBxM1g+epW/fsVG
yICY6tS9Ck+OiflSP5jvM9t3p36QdUqdzsIWqo1y4CT5PJluyhbuYnhkddsjyppQk+bCOBnbsMfy
jL3DeAyXPF1vv5gSQ8ECWuKSisSAxWe7ncIgxr7BAcuGXD8Fmir8uuAaNca5P0TMAgAO9VYg7e73
CvAUglRtLGmpK2dIrYUik4/h1KSTw0Odc8fUxyXvGjRw+sAm/sdmkiHl8i+9Fl/ZOzVU7GK4WXhH
Mp5jKAW48dzix1ZqcozN1Dkwrk/8KGblnyMs0PaSsQnJXOg5ApgM1Gy7FwYjhlo2BgYGT6DUlxnR
gUaLvwirbKjPGrej6EhSZIBTDKwmqcxO6GJSC6wX2rdFinmhWjLUwaeG+UB3BsM41hQjXrO59dzS
/3YFDJZ9zvOYCge35u7AWumaVvcZicbymGeVfApvRVJxbuphFWtawryV30ikkh3lgz0FIAkTMg0a
j6SVomNg5mK0cgmSf1shCov68TXpfo7INOOSGB1p5T6icXYvV5UcfjUdJ5uQS3jC9B1LTDf30XYT
wt/klTqjAXY4PddZrzclDTC02x9YQcGvpfAjPqJOrOOLVuZCdXiF+tRmEpFH6QWDXr00gjJ+5W/8
BeiqVtBohTKU9ZGbRCZTudrS+kii8VORA9gc90DUZBetuJY/GonOcKGH5PSHbXiA4vq3Rl3lbjcu
sOB4H+3CGVZyC17srf2HKEbrJtPcQyabzpHkt0KYy3Z3rSaZhctEaE9rljmXZw5N8dl+6R7FqJ+V
X6asNlzUo94w7wbzZ+9+dHqYuViRBkl4tWyFsolCoQBOKR6ZSXXRnX7AsFww/XP9m1MiI9y4LuCh
FbonayDWbkfZnv5TLxNqvCTbFt1gZagMWxJMv/Hmb+pDmNSJrWqrMlUJj92zWdvovequ4fYZpmuQ
VKEFIBGUaBFAiRte3E5oCB1CjAvtaTfc8cwsaABAjeV7Vp643iLCnaxv3bEE8g4gB3cAMHzCmDE5
w/fRg+Db1GqAWldFa6tlzQTZmGzKq+4t8DXQf+ygbTImczWEy3wS/4qUwcoxOpMfPfrBHruU8XnD
JJXwytv+VBunhmmtrRrJQbVYMHWNxpsTRIrVBLNVt9M2Tkib/i4Y3afxqh2VjzPh7uiHh1kF7Gra
RHdEydgt/cBXD4PUe5RfPB2jGZimWC5AkLu4MKrYyRE9smwmldWMhuLI39Ybn2PVdZhK5hpyUyFe
eupQGUrR38w7fcm/V4BGnZ4aV3MW8DuaaFj9QS9VAK4japMvdXuhVxeI5DwIfIQGgIBeroKhceAu
uycRAa7QK6VWGUWpFsLwQqo4irjOHqzlnMHT2jrZDvyARV6EfA696rRAtVPBSeAnRE6db/GRq35/
K7uxXLh0hgHry2+QW3jiGK1cYr+rEvao0y7TGsZ/ISbiXWVNAyjLoY8NulydksEUCbhQ7tblWijj
UBo2Lv1kQN3PgespjmUM981nFWoq5/I533Kka/kybRuuFWnYt0AOU8yX63S8PXpmK6Nrdbp4pi84
tE2yCme7JqG+87SUkN9nhQ232p0QEQ/XuAJuiIDb1yQiUJLzz/vHdKAsb0Td/WCwbNG6rz7UVNkZ
aMh1HTMjoBCFFgX09DmoFNB7bkhY/67rDdFbKa9DoMW3Pz/1aCCAMLM2av6UJQDvqfH7hyuyLsFx
Oj7qqrLW3T71Zj1Hj8II1T/63QcdziFGgz0H/TTHetAdHL2zS8WiNb1QIUF0ygjr+I/JlZAwO1x7
S2yyBgP7D5RxPNWy++qAp3/uetwKJFEMiRVgUjuQ6JX/9mn+9Te71vtCvHw4Eipf37f0hbQ0WGPd
L/9oTlkg7k/tQ73SBrIeUd1tVx+tXHwBhhHzlgwbSjzGcYw1vwUOPm0me5KMfag7nOu38i/rKUtZ
oRY190sEWP6xxROUmYBBYw7h3fpCbebCWbfGOMuYDwf1O6H0OJIbUtul0Lq664P7wOT5OctA8Gjg
E8LEcBaPo6AQKrRtocXa8hWMPsR2Ik9VumUP1Pf3IjDsLn7dRGKbIEqMfK0Bdtan4uCobey3VMVE
jFihnEolkmJCSd19/iNRINYTiBsELkOHrzMbIDDQRAyRcjwLIhPQfGlMGUwV75DBKVdBcIO3OiI+
SaHN6bc7ou6ueUOroa6GBMuYKe7pRrzSJ8qoaquVf7sWiAm3y9+9PlicJLXqZdtNnnFrp1RBcAOF
XeP32tZ3ckUmNCULA9AwF3K5f+NbT6gGEVjuVwLYIfhggbVo689HOa+1iuDk1RjhZoGrh+SKrJNl
Z0oGTrTSHap0xjpK5kBTCcFZtFeEmV8xEsuBjQhrQV4VvoW4ICnDGfdp+Et1AHxAildacCJJZ2In
l1/IxWvBlLO5OQOKdyUkzIWAz8BKYs7zPFtATWa/Wo4bCf2ydaubLj88H4IE2uxclnfQqM+fXaiI
2GeUtVx9GIt6k/qO6oAWb6ve1qLwHDygzWkNh9EtjImY8fy8FfdJ/mmFg3yOcSWB5WYjlSRMltPE
60GpSgjnGmnUOsUxjv2FYBtICf1b742PpXOn0eJ1E3VwFX4v2tf1wY4wgiSThfPwJ7VpEo0KvKa1
PwzwymENp5cXrqMccmcwxhM6KqcUBRVP5boDS3KH1FVjXqpTzP45yYHTfr+1Scu1GSJXK/iqDXme
753O+o2AELMEOmOQCZhCOKaoai5nq8qQ1ZvMrXxDiQylVY0gVGHpe6Few1nP5m2INAMVHlSfFxN+
CrFbnwo8FywqYKeRV40UxeEFBRnhUT/IvI8MMpDBzz+JJTfWJBHizj48LvX0WayaehvnSzxTy1tE
0sf4L1zct8sCuDZ+r2OXCf55jzCrvYVuTrsYJsBPfxWfhYA4hG7iSYARjnFEBV4VmVCMeJHDX+VG
Qkhq3QLdwODUcS2y8OMYigL+VYcDbJUFELUARHdp16u0D7j2ib2VAqF/bVJfWUNk17pkSn2fxTIb
s/7PHH2p92PQjZ2G0GuuGIbTlfOH8XjX02GNtObDGlQkEj6PUTIHJAVHc4K/muENgw93X3/dkopf
sZ4nihJRqrJUEZ+AvPFv/eaisinGS2uB45MOmI8Wg6x9Wdm/vC8dBa6EHf05gICCfMd+yr4kt0FE
q4E6LNjXbfVZIHOl6JyrsEVAizC3kaoYsfymU+v6nDNLy9pgGVETXC1uPAD4zknpXw3YprZPRwml
xfVOUisGGmZ95PJQ6zdoDFsrRsXN4Kjs0tZp4yAYWhEqLQcb/XATZIUQ0RYjLEJLAkkH8M23ZLQy
eRGFwLU5AW+3LAh/nrUqHpAiFAlvrWnyhRbU+z7eG6z23Hf/5xDPd4p8MyKj9HjoBjKgehTOv4xp
+lbwe9DXAf3Vlbe2a268P9nvafZuqroar1h4Oe3uks+lChRmDnUQ83BWCPqHpOwAHP2RcDHYhjjd
CPJpJgOfX2TinqEAtH8PkcXrld5TGJIajIWKN5IXKxLwDC2Kt23u/frLcP3gM49kUE72bsbOXXGU
yjGVWyfi0hzPjrF+DIQq/1LsW6bSV2AIRkPlQYsCPJ6268J7HAIYu4kq54c+2o+KCAbXEC9ZWTJJ
q5LGsh2Nammrcn6xc1vSO8ZQnp4ov46f0ggINqghOUcJ5KXEx9fdYlTQTr81jnHw699MvHeJQGbU
aea+oQIPKRwFLDU7eUi9GXF6YhFmPeST125Dz/fyDLZHUEXIJy/HUCE3KSdD6k4psg36kw3SYi0P
vuO5BYpVVwqKBGmk0M7ZFKp6ggye+i3CfwAYDQDcMK7jIXS4tiZViPmHkgaraXRnf8PH/8lGqkAQ
C2NYyd3uny2wPDJLye/8/3bfwmcuImITmjBiOSEmXxkX4BT/SQAgkthi2PHELywqpN29Kxa17gUV
t1CSOZxZW//ZBTIEaOBL61zzBe4ws3nKcJcpbKVfHuGN0FPoS3ngjwOlbEmC2I0L2sp4NjIkQX9u
LJLxsGMD04/Zea7XHTCOXf/ipJZWzzRBGF2d/dvwhA6pjlXK6BDTMHZFVlVAoBw8PuVdkYdKpfFQ
mDzmNzNHkFXttNQqE08ZRSKAybUGyJ7CgVInvShiDx2yz5phQOMzNIuHg+ZV63pOOHBcPvyBzqFs
uK76FD/seay/Kaw5jlxOhXhZMDMYBy0sSRo1lqZ+alIVOQ88fx9KfnoDXz0emBYn8gX0b/msYj5u
hzmKIZnK2h87FtgZSUPE6/lWKLnJKNMS8UOqYIA5/5XoXfkaQJYhvgrmkn5CuhChGi/ud/1wOEbG
KnT/rjVYMf/f/a6UDDpRpJOe2k6oNMkw6U5l/iFLXsOEWjUN2glniBV7rAQyLoJ6/vjw4jy74BPf
1iqsaMbq2nhBgfEh5cZp50FdUei3cfGhgJ0mGVFz9XLZkPHe8RqUO8onIQ5Q0MXuTsXLQBCUzoBX
HxPnLkTo2R4O5aXDqFs2BlsRYIa8DbuY3jFfGbzfJ0BXna+RqUptatk2asLHnftLkDK1rIzcrFih
RvbvJUx19mTLyAlMkES+IeEcT1yl8eLIzX0phiXq94+4ERmaeDh4jAreU+XCI9JSXS+HGFDfvQgX
hy72FEKle5dJ/8qhY0+HXFBl/Y6ylEdSw9C27gur1QRu9JJQJhUI07dA6DRF+i+OpPBq8uoaKma0
9hAbzIPzshmNJLoSyuhqEgCZUWPaK1MIOUZN6XosdINnhUgMJzgq0cxFsDRvGzIqolB7weJGZ8yp
c64nHFzwf9GeyLX/udrvibvQDF+42v+89HkgeHVFeAokRgqPVKkWPzMOjAPmK0G1EDPUeSbE9jWS
xAftAz2mKVSqs4HhH5jjSGzu2r6Dw4ekzA837UiLltfeezsdLtIePdKqeZ8aUgTCdG4G0CBtCGj4
ixfDfprUf4axpkXVhw5yRP1fcpJj/J6DHjBOQsoYm0yog/1gU5R1hjFD/9ZLLKs2Sl9Yn2I6QwYT
3EWmWAJMJ8Kazw+P9ojay9cA6q7YK5HJSqqgSD5ix2+cyVedRRpws7JtPJhQNI59NhmuiOODq5Bw
8AHLIylcagP/oN7bH0OIbp5ZUJdMjwYiZqcpfwQl+02id7RlAJCrYeQNIrnYKtytD/+cW4JLIceT
kXTwLT7UnCqCWewuLmIhuuYxEi2MLfzbH8f39FaYE6b7/b/pa6tRIa+8JnTpP/THnQK1DP8cIx5h
CPfD7oRGrGLD0qAz5n/BjZyatM2AEQoLSOqu5gw01iRIo83WOpVaIexZqlCOF40e5zmOJ4qPqFyJ
HTIV7oJUp/9fbaTQrgVCKL4wwoVKFQZV3EYbS/ZYE6INfIuhUqpH2Cn+xiRkvm/Xc+RUVsQsts87
j5rLALGExVb4pjQt1/vzk3GbNmSXOrAUZbMabjMcEmCl6zETWwlj1Pf4IZas/mN+jhNg0T+uQUPx
XhvNH4VYKQMYwm7Tyf6TCSDpHia4aBL2NSV9Dn9phNe+OKCronpAMXSeK2tQnrkAcoYUvlZuXjF3
jR9+erWcBSE96JI90ti6bCie/ucgXLI+pNI9b+Y8Ixc0bcAko0JXChkUcm1tPx1rMqJ+A8yOl3ys
KKnVy0lVWqcpSx7Ov/R1z6GQxaAyXomz+YLw22QYK/UnCw+Khc15MCXB/big/qe9la5PhFVMO1ON
0YKYHtySZ3FvBM+KWcEk6FFskm+vF7arCXwCzXIH+OwKfQ362FYVnqzvDT18RBiVEDDjOVZPsF2n
QqCbAAHtBBLQbrZWjgxGuyFORXlA1C6iEK8keM0ITXxGqPZcCUVNAoWlwkk9lyKkDms5lNsIn+MT
QgeQDpKyBv9qGGSTWQFB3ZyKlJrXt3TEFlhCQ/fyC5suUQEkp8fuW+HKbdFzkzhf3yussiGMbCsX
DnxCTN86SEaAVC8Vlu3T5qg8Uvdh1/Fg4PU3Oo6Ld1svTLj7OLs0AyhJGGZOn7MX9Z+0VlsNzHVH
f2Voqqv02Qm8iO8fQSNB5IFufXdg/xHN/gJDKJivbwzt7vdP7Z1c5SXgTa3D2gmCjtbVyfb1CXOS
O82ZBB6jsF5EpUtxzAjAHFbMw11wGplSU/arH8KfSARijknH/rMIvDH1u5Hqdu3T3AqeyrBLgkTR
FWF7Ign9mzLFbYmhxjQzfQ7Uvoj6r9HzXkkJlpzmhSmg7icU29j2pNNIwxlT7796fDfzkBJgmdF3
YoPfZfO1HOgW/xNV0I1PtEG0n3TcTmoK4eKHDA/zDK+2NzhMvrBuQTWcmUTgIL87y0cReSZiy2yg
F982vNKuUZVbYHtC70dSsi7bvOxCW27CDrtpIVu6FKQPIo/I8CB9ZaP6petN5VOxVkfnv5FKDQat
JTv5G9Og9nrlLfn/k/SSjtmaZhjvULjeJfhpnVRZcu3nIECg7ZhUfWk/vzjJubvtIRAMLZznPdrK
3owpmiRoHBlHjhMDZ4ReegFuOJgjjoQX6Ocb7g9pLOLAp4hPDW8Z+ETcvoDufbLLd4QkXZFr/NVd
0uJ68hVVhwj29GZKuG6ULnoSK2dP+Q65uzK5LPdSXWYrgpwljq3YLZvox4V0pqj855LAivbPUwAP
bkhY/3QMHPepvAp8k2yN0DfG916suZSR/tPhHoQwOH2LQtcosilo8kxb4NLle5Oqjpv/4wp43p6H
IRxMOECm6yZ+MauVMZfsNgDv8acRGzKctFQVBTUt9q2Ebms8DHfKG07u/YCGaRq+ViA2XLim1Jv0
GkQQSImyNON1MsXojKPxj9MEa9HZOd3MnHbHqoS3jtKctRcrtRoBhw0CLvZh6cKoku9uB4OS5/23
vwAQYWALEvKEcGqPaUrvQz3PtqH06Z9am6ynA/VXFdCFSGJowRs0Iv4/ssmljjpuPTbo/d5gPRY/
+YTC+J6HgPuuUHr5Te7BsjypkY4Pd+zrbLJZN4ftl6r0ib7KjXQ8UgeveMBrwn1yn4xKt2/MZgYh
Nec+W1FHQuk13UgdwF8bx9/m/WhMbUek8jISrBe6nD7r86aW4b6CQ3xfItAR7YzHu7IsnFBqe0jc
lQaibJidRntdKdAmV1k8NchQUk0wIyEEKUdc5lOmlEanI2rw5rJtqBiADRCx6nfYVTVEuD42NAoz
gOWfYBV85CHxut/ktD6ayOZHb/CBzQ8PMrvEYJArwbwil0SfD+3tfsw+Kv4Njrf8MTvt4wFBLv37
dSF968GV5CdhM56taljsjjChAwVlAaWk4/q4lNmuQVcJUO5Lzg6Lt9iTo+sq534VjQEw84moR8T2
Fp0NA5cTtQD2JV/kXH7K9213TjQ+QAIeawgJqogHBi3RTyKfqaXp0lIKyW3yxF6lxF/OByIN+gU5
FJQGkLzdnb9z4r/h8fG56WYu3+SdSdn2dw0KQWVjC0XtxWTG4IP3VYzF13h7DqKmUBzJT7RwyKSb
5vcPl+aul6U/wrEwwB0acvslkR9ZDwjtPAhP7fRgSo++9c3KmGLpA0T9Q6/FO3xEcLUkA4tcDs1f
twLCxPTbv1EdE7iP+TZPjL1grdGqOezjpWrxlpBCO1tGsoRLxjy6cmFEa3wMlQYEEsdJd1nt60Px
Ur8kNgXe/mzzAk4NmZUiHmsHayW7iUlny7LC3+XgiDV6yxQTdMx3rLcOTweREGJtD3iYWGtJ086D
iQclWNDDhmlwUAn/mcN3Uw2iuHHJYzWvi3e2HLwAUvpLnDJr6pwJBRIJG0ep9fSwvnrh5ydrf2xL
2+4ISdWEJPlY11E3tgY7I5YzE5PI0bhPwKaYRsqvHXYhvvH7bRpTZOm3Z7N99c/JBhgg+8ySGC24
h04n0Hm/v7ni9VkoEyd/7zdJeeIiVbKhnSQRv3rdwD02DLQttGlNbL4jGa5VchaqN8XXdGBIXDWV
HDJnxiQKy6Rr3JtbZjhAuZSSJ/yvSQaTgU00lVgplXiOVMvvmXeHd08siqmwbKK6VxB3BG2LgdwB
6A6FMN1mtvEL2itpJp7HrN6gULg1EneLEmlcqXtfpA4gSQ4zJvT5iKaUgtyyZwyVnfHOKDuOmMlW
m+ox2TO5462B8X34J6Vya/UVzNn8ua4AsqNWA7NA/IwLYtCo6Rzje9J7M215Y+AtVr6MLAuHlzV5
ksVgAqVaxHof2JaiZia9O2Z3cEZgyJSbwe/nVNq5KhyE84VvCeeiUgxbBrBT9h25tEouPCeQ0/VT
VFejTmbxcCqOLeR1KTrr/q93F2R1fgvlpDe9oXQJ+6KiNgTEGhKOCnHBOptSD1Z2Z7rlVM8uUpn8
fAzcWPoRmoGqZztTiiZl6wM0MlFDKtf5OuJ6vNdgyTBsIyW0FRBJg8rkFC2KjlXDoM2TM1Um+kq4
sV1cZdo4E9KfjpGhH73bikyQGsnFtRkBrH9su1m8zwKOoh92GpPByzBS3j+hGAuODR4f4K7+A3px
XDtvtUXfXoOx62D0TpHbK9L/k08hYxKS5NQf3ONr3zRAp46BGuu+LWmjHMtTwA4xF14l7OoFU+bi
Q9DLrfPXJ/0APvtTGfjwBEUiEyNA9igu7OgJJuB0pJNy5b4xpBCIRcQZdaxs0aJPHPW4dVrkjtx+
U228Txr+F0VFWVoy3ZDTckpSf5QzZPN2eg288gQ/xlA9U3WeoZEZLNtRKKkxH2kWD0Fx434JTUZc
8rz3IyYVcOrNyJTMO0Z3f6i9dQ+GVtf7+ldqsk2cgIxR7lCxlMZjJHrmIWSeSI/8i+Zt5o13ri/I
2TosmAhLxIfph/cjcEGSxW5R6gwQHVMPDBYNkXLsGyjW02b1Wk1cgSfI+dmbrtSLV/UR7Fprq4Tb
lVV+Lhv0RnBgDS1hxXDVmDKsQYvyDFBqLgXccCfCzbGF1N+2T/Jc+vJ1Kbd6CS+S2e+/FbHAzOxW
u00DIVtI4935r7OfyZ69pZawQdFMPxn+fbuIW4VY1qZGJAWHkTfF/65nOh/nQ2qqOZVvx5QMqOdK
fnskgiF4XC5Pk1sjFsH1eHowvxTvAFtzb3hyGhNGV2DjBNqOLpDBzmwotfAe4x7fAQnLsfzr3URv
yvjRvn9ZYTOjn8CKaisn2F+/8JtZTLPJJSfXtlglbRlojyabZ1QBxNnUGGrUwral1TfAukaeFFN8
+NdSfL/uhXoKvOopbRrt6FeULC5/GOsYGAFG7y+UGPqtV6z3K15inDZ0XFCX1/X2AYIAUII6ZyyY
ZYaDqFtHmMLt8hhXkBAw37nCjJ3OKYhUTX3VvkytCzsp1YJh0U4/UdGykGWly6qntRocb0eyDLr9
9oX/YS7Blfj+ZB/81brXmnIMePwV7PWkUeBiLmmPbrnwcaStzn6fRjy/Cm96SkFJZCxDCZS1b6ct
qe9buxuy5pZh5QVai5m7elpdck2IIfy280XJZ7d99Fx0QD4x5tvgySYJx7HXnbw9PsWjuT2k8Mrv
NUhw4pCPCg1usB+1KRaCQp/feAiNgNfLTt5AQ0dRzpfL3d2KQ1ZXiGaUXekzgYPGSLj4ChJXEPaG
CYnnvX7BBz9YxEAPWNp3ItcR/7aa9kiMnKAR2n/R7N+otmY80vS0I70r627rGm6UyxoLZxLcO7uq
EmkgS8NwyeBcin8y6sMtwGgsQ8pSBDme3mqrLMw0mSa9H0GNjLkaxrsQPOQhGNroX3WKRRPBnaDu
Mkq2IH/ZCsdo2hUpOy45Mu/RHc2KEDmzca7RowPzZfM7tTGC5wteDdeVzPBfW+Mp7R08t6nqXqwM
1bq1qRGeSrEREA8Vv+xOENH89pmllkqaMi7dhnqpmLma6QXx3rJHnA7tjch8EpXsjEPjzxj68hPh
Q9OYk2CEPNwQAIRgkowZz3wbeV+Qd+VWYLZBc3winrpAaz7Db8VfqaqnIo93plsEdAfsycBwRQ8U
O278STXHWckso2aL9IXxMhHcYFeJ6BNDBTNKGaw8alswL/CuYUU5/OQn2LUNqozi30bZXIC7Sr/J
ZiVSVi5YsjNq6Fg2z1z588eS7NY/lAyyhb6lDSx430A5p7WKmSHmTibPmr25Bjf1JCtAh60unQTW
aetGEUFxmS+BL76+k9SPaiGZ0IADV0t8sssjQX37Moh2StaTMEB1xGA+PKREYC9TQUIPZZ9Lc1Ve
+ZE/7VK8Oq8T9mP2pktkB2lUYxlHdF2Y1iKe4ZIKMQg/4STBucGIhalt+Oiv+p1dL6q/Jri/kEaA
xeJ35IPsxCrOyD+fp5/i6aHyz7t3Si3etjFU4FoYqK4RaEXUBN3tJcaZqqSzT3wq/2eM7BP9ajta
Ja8skuTcVAItiRHFC4VolbRgmazaqsyk8LzIaIsGorDOq3YX8+Wq4CMuGVmgXhhWx9SzW2+fHmNc
C2sk88HdrMa7mqMsRqXQVw+EC9MrQSfozcf/wvPqYtowf9cAfLsoavfWvtOqbAFeJLm7iYVGOLNp
dWFrHx6wtmUKukt2nHO7gn842i0hiwslhiP4uKq2MLy9U/gdFLY1IVOt/nau/B2W/01NO7rDEHvI
x64VdjCYrybS1BjTgQufRoDdq5aPdSJOfZjnIZf0Ew+uhf6GxKPI6BBPpmPkfSl8p6jP/WHiuWLT
EBmPESzOZ0M6NbYYixvSMO8EqacCaur2WuslMH1iLCVzGHL1HZHiwHK3u2yZUGXUUmB1GRm4Pdo/
K3hcMffAqr3AcrGBFmTtD3kPA5bZw87WPQbp5wItZPTIuXjZYnj2frRnr5xpVNq/NUjMmlhZrjsa
tHcyzbW3rvRqUA6wGlDFCyOjLIEr8baOsQgVKj0OW4ECc6E5H2hpdM1lrSY2+qqoD/TQiY+A5uGd
eZGH3yVZlNHPrJvdbftfQJI8rZ9KiGRCn0HvfHWkYDErZedxEZyMrHnN6kH9bR+AJdFCrLYXSBvj
pHb7zpYHUpOPlqknFcVGs3lcp9hgQRTKQPOdPmEXVJUtQ5SR1IVF084POV6ynv8ijA2R2Fy2TZx6
sO7pAC8nWqpYVu2KY5bSa6gLUBvvzxEgthyVPFnLbNUspkOVnJLAU3acIYtw8gVAJGwgEfEFT81e
+IZsFoIumZb90vvQxnxT4sfORH6hEYFsOFB/CeVL+SHY98TPRJWHxZni1yjQ0Wzoab9E0kHFdUSX
FBwfedK2wy9z+J3HshD4O7iRIQOdoq369gUd48XQ55TGusL+RLcvib96kwIo6WEko/GHoWvObwe+
6AwtDhljsZ+4Eq25WKT3rBUV9zg9KPcg5ulJcRL9YtN/5RHRuQbTx7lhgjLjCWfXpSQpRxC3yZI5
tjUQnvK66yNuMiA7tNsCOgoc5zfX96z7LOPMdArGPkNejNd76oTVInT3xftRC+lJT/2lqjsmS1//
yQlHovQkvBmKP0/M6R4DqXlmtwt8ztZGccKXreP3zGyCpTMDnPZ0OiTB4U9qiXO4DoQdk9c9yOLw
w88ZCmRW6cfkx8coIbzJdizVtsrvWTN95UZLR5vAPEr8fcpp1ZnMD8fkz8MlEo44jd1XYpOLTzle
xsWJnifzia7X5a5WqT4IB5OCy+9LUpFVoODipqCpPFLpaU6+curzrd3sE7WY8O7utWmVy3QMtGMU
Lt4O0wPWTDyVS50lPuAfZrdNzdav2RvcojiwN6Hnf/+zoZLKMtw8k4LAo9c94pY/Ph1VCPYbrR0X
81gk/9sgkeEmyR0lerVlYwy5r92jz7Iv2rY19FInwvINxT4ojpqi0NgC0g8ANZ/wCkAs1Ei7xoiU
hK7O/mGxWfiLuyIz3vB2bCIWGVEAnGXtoSACK36bTdZrQXR0Mw9bLbK7LPCfkdm66tCxq5Lh4c8L
3r/U4kbBAJs1isgjL8FNYPWHDuvfQX4oCmsQ6Sl03AflN/mlCfiMr+7g7yc3hHrV5IsvTMTsPNPN
/XUB5Mb1q8dpL+kTS/B1Y55KHwk+uSCA+uT4rtllEGWjdZtoxykn1LXTVZ7qOD/V1FYU25ONJk7e
Oh3GGTWjd4H2AP9Vvtho8IyVa8ukvDrkByK3JMizprpDjxnB7kXdRniEKAuG9urb5r0kXn/Vfwlo
xYcffn5lWs+5gYJIfBD4pCj+Xb+vpbTuEI8LhMNMyUQiaRs85gpBXl0frgeKthxk0UZ6f4VAv68x
Gmz9W8q44xE6P6cyuslE1FuMtcO9o4cdWQqTU/ojC6DbhCGxq7uU+PXGUHM7vtS5q/2BvmfuLVlo
n8wuoG80H5FguinD9d722b2Zl+iK8UCXKfRHy6WVbMwNS4i2BhypKrK+uETncDVbc7wJgmUp4Ntv
3015/NzNF0Vxs0rkUyTzGQf7rb/B46ZORNy+4izXJIvSOq2kXtM3Bbcz8WgiGUCuxVdhIdSWUz5i
4ISFpF7zPpXuM9gZrV6Atvbqx23Zgcf41nf+HJPGO0swOFBDIFP6kHV6wRT3GMKcmBhEToezb63u
CM2nHnx3KRi01jwH+EG9gIQqTthCapJWBPLZxGj1AAOE46TeuoB2KL/vAqfL7Sl2RuqayOIVhAc8
7OFZ2eTGc4Ee2a+w0QmFpWhPa9qBJwo7Ko+25AxkMBOkDEV63fiinLsj5oJlt8N55VlcjDNLP8iA
nRsKGd/RHqWnE4Ftnf/DGian7YLe44uCjvW2D3BqpST898tzqTwwZHLNfVQoxN5zaL197+wKIr7C
2U2Nn+V9aalmZO3Ic0Dr15MEVYZnHuYwlQGmas83btevq9DJqJhWb1oXn64Iqt6W9HfxdyepsqGY
XoP7wlsiY1+0EQKBytxdjUIqdkpGJQRSlcCQRGaGWTDc9KhPXxZ0ZVt88tIjLgujdIeHzq1wxD/H
Jsd7elQ59K1RezjtDNYNfQKGI/BIyvRZ5qrBH4K1ZZIyxRkF+6uLPpL1jYw1NzGWxQZP8JngpFSA
CTgJ5UA68l6Jb74sBS8YET6RJwmgtVAUf4G9paR+w7gV+wb9KWXXE5OyuPtGzrPCOqjJ9YUkB1vT
LUdxlg69PcCF2T31eH7bc/qt/G83aP2BuN1FCeSKd7+pulRqCJUAUECzI/LJtioSyfpBvPiisAkD
0OM4RCZiqEoa6dkSaYkzEMf7EYSeu2deYfT1pj36vjh5rAM1zMx9d1A1ENK1lXDGEJAO6yPHKcQW
B4KDbnnzmdstwXca7qAJNOl9BtwDEbziVQzGjkwWvgPwv7oIJ3wqbFyMSHpqZI9JTHq4e9ptlxrJ
Td7LiJhwfE0Eti7vRYAjQwBh07+T3G+mxXkuqF1yzy1BV1q6Pcqab6070zdGa98776PBcmNq9O+d
uxRRRimRRDP7upiWZv4TB+k62sr7fGwMccbsFMdBQSYDzIBdPMvQCAaFcLF5aMppAZZ3jKLKyGHj
NRksHdpxhWnohQN+/z4lbMSMZG5YE20Afmz3VSNctvaxrza0k/7TVRpoiYy3TSCImXNxsmaJgtP+
YdgbdwNr1xvperz8Q36z142Mgia9e8QT6DXvYO30KE7tU7NhmzoLxUzP8xojNZ+eAZj5+K02yxV2
8+FPZHMM4H7VeRtBKQQ9IqTjSYFeH7K0A1uh3qfR59e6tldaltpTCvelNsNWM0FJScFr4mHbvzKI
VZTVOGWE+1xmt/HIMymoGhk6BIbVL2v9EAMq3QM5Kt4Zr7jK8UtdZeUuVnHm3qw7HRyVIioWSwOh
i1nWAsNS1B3NCuWdo6SiXXPhizTO/pfD9GPlGdmWQABcslqmn7ocY4vbpBv3A1TPTPCF35ojm0Q8
QbcsfSvYuSch4ZgWEtkVWrkKN5wgL4o+rwN/bd0WtVOJYCFK+xvjnmQUigFsdiuP65zM1Tei6JvT
tlZeWSsxZmdGpiYJyEq0Sx4M2YbK4N2vzdgPETdYyEhlQot5v71LJqiS9/ihVxmoVRKdl5av91oS
72v+RuxEJJmKmvoXRVuhOuEmdpYc752NJg/trP9aVudcDpRn2TSV7UG6+XDO5D54DRdItpYT0UGs
wEUjJhB8SaoOoziC3Euq6ZncealXP0GdgmKmbeNdoLOz9rFRo4rArG6pyQQwbk/AcS7gmQ+dWNyq
FNOyyJCxqtvqmOXKvEBrR9x824LNSEBkLsBaJVzbSJQ6Q2GTns3/LCznN4WxRgI3Q3AKPtByGGx6
4P+3n1Cxv9QadoSFnHHAs5C5V/j/1PwYD66irKpndJ4o59HWpv9j4wBt+r5J7lh4//FXITh258kb
PY3eOFjigfMVp5qSDcqS9/TFEzg9WtSM5dF+S8NM3x9OyXyUmbuHmKJIVzcmYyy65RZwEpe6V6gD
mbboq8xM4hp7IhZqaF0oXq+NIp7UnFlOvihXlrXE9/pZKoavBAk6y84J9vjqyqdRfwyg653jQi+r
aMy5Le6kVbuNp274ZnNYR3rKHVOHXIa/c1emgxXv4gvVdiPxoGO7YO4Fqbu6KeGteaDAtssos1wy
0m7IwSjxl6dtzdgO3PVvTXxVKLxv8kDVfGrTP0po5SdGJZHfvdaYaYmLlAjxl1t5pSRuQPBFA3fT
ZROpbrxozCM7CFC5GRPTD472geovHADwjCh0/sDooJSEI6jCrvhG0RDtvHGkMiwxf5GBkQELUw2+
7/ndXYfzcyGRUrvkgrJF5rEesEquibYjntDKcbKnHGclZ9EweoPD4qkFRAL2LHzozKYimM+PC5ze
1kti+I9WspdRcjmd+A4t6rFOmPd+9DKLigEQA7E/5/4P3mFvTVRb3QhBKH9g2JzMsuCm01ize4hv
v2QHaUnFreSSUr96RVxxmAJFoy0fJ9aeNARpssEWVZVuQOtJrugoE+EqeaYTduuMrhjIY2YeRSiN
w4XGOABZ9rid0V4wcECZm15H9c6DUW+iD2qU3fBcKEU28LZ6+UU1GA3PqMBSb9jYIqLJzJuwFTIR
4EXwxGOTYbvRyjCvzrkWzMcRGk6svJJhmBuT1Pas5MXCnn7ktqtwf+1Ey7eo1Sb1QKaAwC1IvM/D
VhZ8JHcGhy8uAHgBsDQiFKToi8UST15vMFqLVkHR4QupjLeISA5a4qcg7+jgwRZGbNQm8FE39g6W
mGLxqcATzK03tO1v9NGGcrwq3yJwlPv892u34VaBm/n+iyIatvAsJJElgjz5mn1KHhsssIzl/GDV
C65QkaVaiG6yZWJ1f3nUrJgXLSpHtDgDSmdjga+z3taqeqNxDW7x6ZOQeE/qxSpLX9UkxIuf1CyY
ciUUj7BAJfxfM+730/LzkiZgf4jBDAoDJaIIa1tAAgrHtKQqKwK+vjoYNmRn/dkyngILE3A1j/XV
sibOjl3aNh865jGBqqmrIzEcPaX2jTqCzcmTmpe+U8LXquVF/oRRF8Ae1X61vK/N9+DZZ4QcDX07
E/yfpoBjtbVcxb6q1Lup8rc8rzNuffXtDWiA8zIBE+eRR7YdYCKtr09fhIbWCuQGlvi7GWCn/u06
g4qFyT/bY+CVOPWtNieHMSrmryMqdKNA7vjjbp2zYLA5fgGCaClGFJRMJhxhiXnqvrFI4yU1zq5h
AKIIhfg4QZLApyTHIeOUoBJxFqs2NoKBes1w6EscZoWfa4U5ELwD38cBQFOIxMfnZyj4Suy+CR8d
KwlMY0EjKBYreLe9qw6NBJBWYxTB/Nxk0Y2Y9qbAktl/RaIebBprLrYeeqr37S2sR+n3m3bw30/Q
P3ONwg8+NX9dswTvGMfnZWwTEq6pCfny3ww2qI2PgsONBqeA6+hX0yYDP/AyP20Re53B5Biybcrq
3iJY4ApKCUAWh2+bmR4t/Lj1F445i+xBhpBBgM6+N/zacRrhhsBQwD/kUjDHOnL3y25MdCdVLyuN
xo6Dj6OqIQXNcirDkV4RslspdqeTF9fVy1X6FX1HoimFiHmQciHQNT2FntbSNs0aaomiF34N7gwL
sl0Iph9q2siFIOjTUdtRdD/2N7jgp2iO05EF2mons00oEgcnJc5gMs++CWpsU0QdEnZ9B1asnJ7A
cWXgdVMHMbtmlaBcM6NXGcczm3HFgH2E7YTOq5Pz+91JcMUg+g9NH3Xjsf06iw3dSBZgN5ZzlCpc
SB7o8RTe2FEjiahqSbe+SOWZh9oB8C8tu8/E7DTeZtZ0P5QnONTD67VKlOsbpvek9hgiW/tie2MJ
G47ay95bi3dg+iVCAr/Pd+UgBgNt59Q98EJDJk/3suhoo1zQj6EwRa0FVIaiQLkd9WHPFvqz4vvD
8c7gKWwvnb/UyFnwhrTAyXKkCTKLv3yS/ntRs4bv4LUgMeO8gaoQayLxkC1lq1y5Nivz8IjyuWHh
JY0nrn8BrPjTNBHTtvFChXmewYIxRE7OZ4+WR9pFDCcId8OHH5X5CDTDynp47g9Y5A9YeZncHonA
Sgq+kdw9X58BwtoQVQo30lAIqKQReNqXh2vbjeWueDOzaMElwsOms7D/+8nzLkX2MFIrXYe5+hGs
Xzq8y9w7giL6eFWMshXn46DvQsWgjk5oeBGomna/g02RozS+h0HLrL1RGyI4ESUSEsGLMIyWFfUI
1tlykXXcNJvgKP7xkW8gVuwxL9adkaicxIPzEmO5MFf4U93loof1QSrYW7YrT75wcrAD/SDYxQv2
V7vdrCmEvqfoHLuOoUoMrndp/3uxmL/kFDKw54yOotZpziNM+DSuVPCBZ5YHGpY9gUx2ZD2W5qM2
1y4+Xab7ToIR4XeYqryR6Qu4CKde6KKfvwGUF/Zz4K5zCqB/5UxhgY/LvoTMBM2SYCcvtfacHBSs
oZlozwBB44FbboePWSwd0KBnAjArrY3vtbI7q/aZizDfFcFuyueFwpgD5T4K8W/V/JXfXR+a/MT0
HGyO+Tzbrhjz9hqnj9hkhdfcDp0CSgOPcMex/nevBnoXOM2qHzKuMIyelhe0+jkiuceECVJsQxq8
AMEqCpBQ0t26AZrTi/botGXrDKFLshph4i5UyHQAcjOfIvrc9czlzOiZS9LA38m4D3ZWAJiuVu4c
wet9+fStFP86I0iX5syWqo4dkMdGrPAFo4ItikmejbnJ1c1QH4HJTH+qeGfP5daKo/WXZsVDPqQU
rjoMKwXUp3wwDRLBfTD1wsltDf88x6Dg+HxqsF3zB1sgGpwxbNEfuHWZKpwYg3aVG7hUuwMMM9aS
ebnJTgtq+g3hxzVYcaeaVBglrkMAa163JXT1AthxakhRN6QYckO1/6bcIHisI6/FFEBprbWVPvZL
wEbH/MpFLk/zTdH9YnKApYzHUgX/gdetyarQ77tcAm1365JRxBPWiPAOEFFsKkgzlsKcbOzrLBrD
oJWvRA6YCXoYAI9dyZMycJPGeLmugODp7Elktc2Z3a/5zfzdE1aZVxONXvjUgi4rrYFEwZreK75S
KwVXgls9MifI/4S3X3xW/3DH7yNcqe0wAt3q92cLWipgDUNUHj0IAlsKnAPa2jH9SUnAk1UMyQuf
3c5STqT5BWnOtLtk3ns15c1MXD1PzSFzur4FLXXbgzPcOD5xyQyXbC3+P+jITUQiosfUxiWVowYR
CJR7jeQzOK6O0c8W6amfTNqQhNwBAbQpvDUTX3uL9HbNOq4jLBjOKvuNuE84ZxMSmtBgSCGT8OVV
tW+8uUtApztrzjYl14k++WE6iXyVcrpBT/wfAHCxJMznttNPE/lMCLl011WFmdhwtSmunGwZUpgN
0pGrO+w+6umTS6lhwDGc8kM2ate39gARXFJL9nZkDqvdbK1Jb5BzhvmlLiSxZw8lh2psM5MTNveM
SgskCY0y37GN/0XAb63PkttpJe7Y6KaRYkKs3fsSfPye0WKEGl3RXcK6xvPAquPl/acSGdLOBijz
OpJ13Y2+rpUs5caUyZAGaOV+J8PaVczNnNlYGWFMpJBVZayHOfNQWQEYS1z0quQZcbAN0qbVjiCZ
cqO05eUkKxa67vN96rQXDOjj/EjXNYyMYw/tNGH+utnVIEY0bsn+C4lPbns9KKfPcfZB1dOzWrKy
5vKnPrluZDaBGkPkbJQF2B2peUt3JZaCbkLFqc0etjWKCrKBmC4KrtSQTTnRH30PFI3omVfxodq6
ZVJ46xVrbo83ht+91iOBcj4SQX6x++kx0EPLzMvT7oNe9LXi9rjbpD9Z1OBHB9gn1xWqhajzIaX1
b5ahDo304EMY9lipqdZli8SpDQmpdoePAFUbaYWOTlP1mm5tzoeHN65++efB87WRy/lVjqVDUbr4
Z2I1SJ7kp95sJHnE2R0ZQWrxo8KPMBIvCW0VY1kToHRnelGikHrMVGj+Q9q3nu6tVtg/6PRIZGwW
rtXq0eA2OQP8xRZ7ZJ29aCY1oD/2ILonobv+YH7Ej1u1zZsdiiRi9nl3tljKmDGTANZB0+O9bp4r
uDcjSMLdZnaNrdmYAShwhyuau34z15Mbhy9HGX3PKN21PaFh0ZNtagmkvW+kL6GAm29TezIA1blY
054uUemTOOUPtdRU2wX1/Q7AdQc3sF/GdvEigyXQmIYe18/gyh+ZZzI9dTL0seUU+Pn+7PAbUZBL
wBW8doZlZ9Y+6eJaQdmeeSjkfa+XKmtdFC6X6iCNOLRV1Ts0MOyXfZmiFcmtnM1BaO7ahfWN/Pba
5Rvn+sHRkr/LAom6QaOnMuTD+tMQ5oERD0CFTtbnijrB9idzwSkLfCUkWVBHClx0Su8weOkYcvoN
ipDLEeExCopa6UJUImBGDOXOzrGziPVvCpgua5ehDfu0JBdcEEdxQ4UKsYxnCLvINWH6Kjmc/1dE
6ZwEXiq4v6oI0mYKlamKfOKbNHQLcD6PX6wt5t/P1oRGNuK0e4YQVtqdS1nGB3T8N3+OuklD7OZb
/DzPQjpcFj3iwnkpoOtMOMqpasUDhaEPSA9nobYWbVoRI/UD73DB/KpjP7mNFB+VZ7fVTq94LM5Y
t3tZ20kfAymZusrmlt1VS+1yvihhwCVh9oh5kqaDw+JIzAXqntl57w5D2nENGb9p1BXudmbxXbFC
HuP4HbY44ZhzHHEg7Gr/hEGOdLnULtwHbVRkFw3C4mLXc/AK6dYR+Yw4K8qcvK1fhGsLzSIev2vM
0dN414baz4gUVqIUOW6ECesquZtd0w/jIOeqwvWOmHgCX+PuCXBVqHbtgSMZXrwkQLC7a4mPwNG4
BfIckoDPNICKinfWLTrj4e17tVYzkbrD3sDVRwvcBc+TSHbtBQqDrIeHZx6+4gwp+Zw9OUvS4zqB
DZ9REDA6+mhlESqsRppRfqwOdZDgU+Nnvq3lw37T8OQvZ2H0q4Ye0QmoSMylzfZbIFTO9kYqMQDk
JMfLd9iaROfFi91tOJbeuNN24ZMm427Z9nFBw3H8zbytyNFt4zgnDMb2S+9Un4NND5afvZYKQQWG
AJCynWpMBqR8DuQ0w9G4pABITNJQqjG5jgPwU+ppLvhs3OL3keMppNe6F7AWHhDrulPcP1VfGqX9
G8Ko9vx2XVBT1/hf1XUnguqcq7ybi4JFqP9cBbtR5GUAhwoL2BZ3NZiFbQGAtjT4awTIKIa66mB3
wEGXWoVYySwrFY8xjXXCDn2oWJtWrvnnMrKhp97OS9O7oKvcTmmWzGurCbf2jzbKoMzGi/ZEjPzB
V3ZtXaHlOd1M6RaCAVo/nQXJlTOzuRqO3ySKMg1d6jzltlRCtSVuVWA1g/j93Z+fATb00QY3eS93
GEXcnHVJjRyHZeVZc4Q82q2ZxkjFFXa9PAGH+vhf9PN/buFmIccxP+2Ezaf6nW+vpQ82cngrumWE
gnSF+PG2jO0g2TOSYotLiuG/wvUrlVYYDO/StLBrZk9ydLz0UNuO4FZ/PTD8Rlymau++kdiB3ko3
7RNRCD+uJZNRIaN5y6uOv84jq2APBJQq6PvEszt/Y36zFF+nETUfNcjEH+KLvfStZZnPk+h/bYGw
8TCh9KFhc5MwU1N2KWjAJ60wEG8aEe8GVM3wr6FhQ6F+MSm3KBhI35rmsYSealJeH82k/u/Lpjnx
yVdSpuEF5txbT8fFOxV/6amqgmJYg7BWR/TkMsK6dxNEXvFHcvuERChP94N+/+0v9q+PtB68CyS6
Ju/f74fNV2FDVohj2avTsKVtpPTQYmA8g3/PXdO2uz50gIaqARoL3Fi17FxvFEnl/aH9dQhsQopm
JuylLGLWXLycElmexDEbRD5rcXKBaAHrPc9sdDjexZS1EkYZmfDcT0iirgurDhw2TqtmwFA5O9Lt
QH/caX8D/nZUrEIAuJS/c62EwvAksFn0pyCUL9DwJKNCqDy947HXMFGC2Rkapdxcz3QLdPOE0iH/
XJgqUvBrXXsETTesvazWSLWHNb/TnK8n0VXNFwkITdFMUl+y7EZ/BFz8gtynGMGU4mCN4lg+5XZn
tVU7DPEzou37yW61usMu7Jx/T+61lCC3thmAy9xRsW1LpL0X55JG9nieAyJHDQ0DU/jjzVphnM05
C59p1/BUDRySb7i13k5c9gtKW0pd4yJ+0SIMzgtl8n8Ic+BdohyHZgeEBNg1AKiOylorsI2HO9w3
juhZ/wzhQpXb6u2rk+K+iQ+YNtVIGkbMbCSx0pSOLZapUbfE4ng43Wc0jIARuLAhvZkjutnB3/9c
jweT/Pt94PQpgyNofAneUI/wIUxSz3nnvLOUIYmpS+erZiST+tQA+wcexd4hnIPqlQTsKNCgYCMr
jVXmE1J1cgIWzeESgI1HQ9LRZuwUxXPQjm1cmQV10jTCbDe/C8TVomSf3iReoD/HLfMslE1H4mGr
txvCkXZleWyxkCpzeeZfmv5H9wKtzhxYFBWogqXx0WndwO2eMRRJSmdFdsUwAtywUtrYkbT1DsuF
GLvzvucoT94vHyQWi73YJimvGSZ3uips7oMwsSWy5/IfHHncEMHuTYsw2vWpaABcop6ay1H3Q9QT
KvM50QKVKujA0HrQ33Y640Mzf7bEvHo5mAMn+PkejtaVf7mXl9uFXYlr+m2XzigWcdFm8kOimb2i
mqo9/9AvQGxe4bQAiNxrOhqvkHvGF9JrO8l0zuzRXmo/cDcomUpSkI+jJ6GKhdltgl4NEyEv2hA0
ye8gO4ag4Qfsro8RPYvIQdFs7NIzHXy1egEaIFJYBdz/gCcOsqsj0HxiNWsFLsy/BhkQKCTWme4e
39a2BsmjVX39/LRuvJaX1PV3nv5Y8HrvoG/yg7bgSmhRgHIxsdcsodtxS9vF11SIOofBieIlrcNP
hM1uBWOsROQ2FIS/Hq//m8bz+iQoCWQ0p2lpUcOp0x9cmTcY9dRHBXen2CAyfG0MBPMlZVeKBPp0
u1JLm6B3C0PLPkGqS3LYxg/aPUwJa2iMR9ewtT3E+NJ1QZtiUDpiiEadtmkNgki9w3MhC+54dY0p
9WeqT+FJ93KHsPH0pb6OtRpH/mRp6cAxP8xtPcCsSkr8nE2kz7qFq5mj+TZAV9sg9wb51HVwAVns
3Jg3F71PW9GaBuBwKKa/oz75AILqPvhIIf/p6jb8gvcFTfnEl1myFZpzU2yC3P5cHVWh2ozz7whP
h5wQ0a/jxkCpSZO4Oi7MXQHKeuBBOZ6BKycSF3mMbBe0iCNB+CqzqbZRHkZFm8dkiD3GtpJ8rwE4
MkQf4JKDK82Xos0CpBupPOb+8/NAxJVqklYM+WCWDxUIqfO2zLcImu7RcPo9EDLjleg7vXufb7c0
GrGrNj5LifWgN68Icdnl4FRYiG14wOUIPaqlzcy2JSMr17gHPs4LUVHzefvSCv15QfOhPlUO4VgN
xGdsLWos5ajhN/jvJg00qlDXfoXBUNqBgXWvHGNNob68cdAkyJKcUv2g5BfN/crwUoHCXou18jqD
Z2X5LNSuo9B9nmaapFJLMBzzDREF08sM57omLOBPOiln4/ifAcOmrHTJ11nHST3mICtH8kpUuRUk
b0uQoF2VG52LvRuZ85fK2D3VBhNbSR7aN4kne4QQHDGbd20s+pWe/8M5QsTE5SU7zTQcNNvSEubK
M5mEotb71/tgEkC6zhaIj6vENpU803y0UlIaYBgJ1Uj/RaJ+FA3RyGIT4tkPiFC1f3hOe4J5lCjW
je8RIGZSJ5/pecAfZi5D7V5l2cWYt/CEAyVALGDyJUIUojhmZi62B1WP4gmqz/VUgqxyWiPtlLZW
zSvm3L1Axni3u6Kzta84ZW1yak/L9kaaFCTaRiTqU6keQaSpkQkVWyzxWOsC7yzxU79C22+kMugF
zs6ChwVPQ9a6OsfrTrnwAGhAWEtbTaEPAlR1Y7GPzQled7c4Y4E0cT0Z4+fNF7CVaVbMvq9krII0
+pq44l3PgxA0pGw+GWTzIbGaZdawO6IIAqLDb13JlS9mx7C1yGWHxrFREBo8oZsmIOljdDtU0Cf6
MJ1c7xWjrUZkXyvL63vADT62FTwIA9p7gjxiEvzHSAxGhJ2ipIoGJdDCazCPw/RCQQTq5xNSkXZs
uRRZSmxX5F3oEpIYy1lULBokmF1PpJMYCRF/ZsXdxqISAmu+s3UmnzLQTTPCFxhmuljpwhNZD/sj
WrJ+ZdwLaq11fB9KQHELDCV4J+XWdu3f3cPmWHEOwx5Uc+EvnuuHyuRX14hZLoXVwbPQ2KyWgVU/
9XgRePy65sChfS1eotqy5H9tqRvT7rJmqoDmD6oVG6G6CxpjRg03G0WBpciPo8mCLnFYxBE67xma
tkKfLw6CNK6U2KHTZT6mH70zBAWqYi3SF055XfsEcf5BmJAiHv6hDX8l4O8iOXW6o0J3q7YHHDSS
J3tU/HNlIFT127a60Ag4/1IqddX3O6UydRE+dAOYyJPIfo79870dn3xLvtD5ZGTokd/bb0j9lrGz
nSv0U0h2mSwgBAQnrW5dxG5FXS80Zd+42mEXDuTJrWSBKrt/heqNKqD6XtiIYVd9qP5AlP8j3TkO
eahPPECdjqxA7FMEs/dWefKqBzrNkrarQMg+wsXuHZKo0fOn7+fMzFmAU8zNauPk04BMVAlmZ9Fl
A4Mx+1kLsyJViKFBU6d6wn/fKt0CsBMWwXXoVYXhksJc1PZ/u2nijrs+6ZKWD5qGwYaCXzCHA68l
7l6haQf3JT/NUTulYk+Y+nD9ghfkVj6Y577K2NChMLFSMiIAy1OsLjnWtiGzJi07HTycDGejp1Md
bNwPuWnFtkdDqElpRY6qsv9oLV1lT3Umc1nAxuh1oZMm8/LmX6zkmiyFLKYUv2rTYeHwE9fwDjdS
5JogkrfjmPJoT7OYHX3gbmUlFSE2K2smXKSB56N7UMlSSGE6u9yPKWkBM3h+dtTB3DDldoBB5OHU
hyxlUyrbwjyO1JMYIrviSJZvSbcrbNhDHExHOgwrvg5tFYmRd5tzLH8oUDy2KAwKe855LU36hB/j
bxo+QqfiJVUDKE44e8eoJ7iORkewUxlTzfaSC7adctubXikMGNA7DJhkeUyKyGvavYdzVvwR4cUg
D5H8n0TLya2S8CYslTwNRcDZMIFrMp7BmzOXlT3O/5CN2u6xwkiisZNGFnmNDpY7LT7Q1BSTrmHC
zQwb9bBlrZosoGQeH32Fda9PvMk/vfpeqdfkSV5rTpb8+AoJaYqyycsk+SYWcwwF+0fQ58KtuOOU
9NJxR1LeURU8hFrsoMR/dmmIZluFKdGtpH+zTFP9mMAHcZC/cSv9Zwz8VyQu5Ldtf0KwmJleBOM5
qhp2LZhbkpw2QNT2SZaRvIrBMbluSfUZUVu3epezKUKGJm/S0/XtLm6RLVmFOTJwtYGkt4GD01WG
2PdekvQgH1uvhcITVON0WMh5qOQpQFST3D8OBJpEkUQM6nZ+zCvA5LBCQhSRaQmNQGUM622zEmfo
0oma/znPNx9J+QoGoNt7kWzkdWU6S+mEvYPAKe+b/Jo0icGadarqIOOufcPWCoZi2qq4nXdSHQBg
mBKUE6QU+mYWjemN1eEe0gLnSB0DWo9a6IURf02XD9GUW7I1hUINIL2RgFnoWIeEP9ZBCOD+2sxM
DqymKfCS+vDnvXx0x8HlENQI+aWd0jftsLLnJ3kp1pTYdqgmfPqdjv4HONnNEcMc+dx99KYCWf5U
9+lPHibRx9tGb8t2akpncLXOdFlBTKj9PZ93Jwa0R9ywK4DomCxG0gXBXWq7qVu3ct2SSNvdh3qm
Mk953TJxnBN1cJoWZbQQTGqm4JMCEz3HoMXCxfS6hr9hk1dqW3/CuVH+Nfh1hebjEh5OV2QhMud0
sn4LbV6Si6pbWviQrYUbw05zNsKt6Xh3Z368Aa1WRBm92mhsZy1IJmDr/BMaKTx1ofjaW4iDK/7a
FFnqzupQVaUgF46hPZmZ4dVefV0zzgV0/mK2OzNJZo8bhFcWpOaQ8DURXAtBV75zY/o7SVffaPSU
OqTGXg6hQp8yDIfNk75cele3U++PxQWpyJxx3YBD7KDiXwF6dR3Qk/e2Joc3b7CRVehwRDaLePD+
99MTdfNMDiBbazYQ/NfDEsJfD/c38ccd5Ge0ZJUFJBUoH3WicJFMDWdwt2GVL9Tp4BiqsqYIup14
I1ZlPwNikkRsUhO1JwpOp0+lxgxMf2MpM6GSRGiU0CNL8dhGH/Pqm6tBpKO+UTEA/V9GpDCg/+iD
P/g4oUaGjc7+EZ0H6BMsUNgfRQMbSMVotBa/Ob9uQwUFf7sQcLoLed5fu7Ucx1KcqFb1+fUa6HCK
98/w6KXTqsp9rbaceMmyVDOtSKpbaiHWoMzAK/5fmimL7PO6pcv+cVDnF8xwa39svsJdUolYPoqf
ScNGIdAJ1WYw/V5UwyZDivYDgvlQ8RZpb6nyp6fvLZ4eK4wmtDus/NxJO1zMJoScnaxNUjYzAYv5
bsIFGVQwzRXEN11UWo7i3PbwgnhFMFUdq+jgqR9vq+ZCPwJ4i1wzgMUg/6OVLFUojcdQGZpselV5
57ZMfVGgcozlVzb/Rwy3Bfx6bmR2iYOuu/0EcDFYJhtroExUC4PgY7QUoBep4UemaZ/9hem+/DsB
x3uUmDSFE+hlB/wn4gDtxXpb/UGeAOnPjvFblSWhCmJOAKH0uUJo5T3xLYTUT3tdIBPQG93c+jRi
oFnFnlrVx2wwUSGldNpsyOmTvxVd+Da1i8xJuxROkS64QMb5xxtWHDow75st1Y/pl0vd36CfI78N
wt00YdvAvz3NfDaOrFRLA7fhAaUJCBr+2hfXYsQ9u2YjYSnjpkprNwDpaGq742KZLZ/7EHVfiHPl
mdXrq8oZcR3YAnNa/xELcPWHw9qgbupdsGSO721K+pI9RPm8XnGGaC5wpcpcU5o9/h6QpWjx6WeZ
9R5X3QMN1eTMGflBoHPPltwxmZnxal7SrqBPv9FzN7xTLAgajKcv4Nr9drhaIwHk0OULpmQVdhGM
rD27WTwlbPyKlu5h9psDJ20kiSgRgCZVAQFQJAseQL2z5pCnsft34XsL6ndm+ck6Fs8/vFa/Ql1w
e5B1cgH77Kh/An0HRuI8lgjhFqIZx5CAxymWrld9CcTv3YtKCGmmzuuQgogdlcQX9U+vT29pvBVr
yfK4j/SalR19KpetX5S0xHAJrFay4TBWYD/KuE8iMVuYxnpjLJDWnTJ8o/COrmtyE1y4L2anVBVL
G/R2WfHpICv7hMr3ofiQPU2EoLsKTe0q0ATgVhk4oV3BDhPwI4dSAl1wjjl4taybt1JRKYDemn5f
mU+A46JQaf3tvuRP30ZZH5p1mKfGgXJrBK5KVmtK6vhVC9Wm7fXdGbFW6cUDQtZml+9jfuXN/+oS
MxZSHJCKId3LBcrZra1pZZK6TPPn1uUBxulePExpBVzXfH9/wjYm47xMA3+LrtqGYQkNxNLct6O/
0nPCotGFsg6d0FSIyWJvacVFVnjxx8Qh3cdpL726riZ9X8bLK048RHepZx9uVvdNiGKwqlTMNMb6
v4BpYBwmweg0UbmyN2/ZOe5m1t69G8KofLwL1UWQ/x7n5tiX0WsD5zikBFNYQh7HrKLesKjhg0X2
6BiJESKIPOEsX55KMrWh1izbrQPKRJd2dEMMasdsUHLXvredsrxOK5pYyuKYz8Eui7AlB6SynId9
DJtLctPTzaWbMJrM5CEWy9XVt5hwTpq6RoSrKzzSTlTV/hDAbodguTKh2SgByIMj1y9F/R0DiyIJ
egyff2JPD+wnwQt3i78OokTUeEN4rLm6Mg87kQSyK5KoZXdTy16nkImSgzCTbYkaXEGYMqcMcQ4v
Z8MVZZnzmMzcUSHVIm1tBn0cuIowujvi/0Mx+yPtVmZwPzbYI/Y0pPC4pyDATMa0hbLYdGL/k6cf
Azdz/s6zvB1RFUvSUiWZIpVp7h/GAEF6RMCahBS2VacCDvQ8keXDi+JDRhnCfZNX9i8fvDhfPGgz
maYbQ74GhbqIqXFJHXOid/+7a7iOwEjiyAHxO3cc6xq/wreiZW9VEBpyDMEEIu4YOwOTpXiVb7lV
Vy5imvxJNuzQ9hq2wWGvy9L3+fU+vl0HEenx7O/C4qXoApKD/dKUuFBJKYbUL/OblSEGAreqApgy
vbJExOkDHy0eDL5jEfHWyVbwohiyaw3nUPBl0bHVvDiUwwJyov+X9ga30I3GpZDli25cQ4OFgsf4
AqV68JNumzDYMrvhvsu5jGMfe6pAfB9gILBcFBwgRZgCzofYZuzZD9RD2xYLE0ojk7AwxQUJALMF
RW2A1+Y6L26R+7TRJIVO9eYncGhOaYsNVvIWljaFXtrPXclh7iPGTkn4AWsgXWcoPQAXnguXIUFN
rvpBV4FOsASgRuEZI2S+lvGesGhhq+jUoUz0co19desJqVzOxiRNczjUsg0HiakC49JdowHQaaRM
fkvAF6qiLrMte5G7rIH1WjtKm3awhlbMwnNsU7lCntbZBHdSapClsDbwJ80DuHJoijIE7xluahWG
Kc2ukrFBopS8o56iQ4IfBkHfDFBIdRCwcJmCMwAM6Uqxnd7VyYy/3/JWszXpKHHv4JQaPY9DOQb8
+FS4Pq81Ci0sJ5UF7CNqAwWDg0cDK+A9pxR3CM2W5UaxYz7kQnSqIEA/kohGjm/6wSHPlTeAezKq
1SaA0WBLF+NIHNX23wYdaB4G+K/V1xRIhjNB631qrpv8BhyRC5e5hoZaLPZH+nbYUNaZpTlij3px
YrwNGmWf3wPBNl3CqupaU8a3CmA4Rx3A0dijSCPk6QNK4IbP1w7mwBrCg78c0xsAmHPHr/Mzqlwm
6xzdtO6E7hjGRauO1UKeoC9G9JgfoYInvOyODQirXz4IUbuk5VDZblvPP4VZ5iInhcRM3hlUpefO
JExL1sF0VRHvolLYciOmPIra8po8/IdwzYTd3OgODkwyepoUo9LYCGLTQARK5l4E09totEgcPh8u
cgD8wD8rDCTaDJrx9lZqq3T3uho7FZ3WSN0wH2GtNbC7CjVBNpvMmxgHBU/gsUVRZvQXdZ/5lrVH
/vNXsaVwySQGIN3mISVyY7vQQjDW3fhIFz3gEsKYRARxtjxAhz5SSiWZNfO1aHfK2ApPwBbNbdmL
8COIFvM79/bo1wvymVJdIJTa+N1te0rBE1EHPVlGmbeV5hWzL6NzoznYXg/gG5/ds4fHWMM8QqSs
aUl/ZuhaE+V4zP7yeEoAURPjUFGDtX8dfHc3znqQG4/Xu7crqFfqFuUmeiSPCddit0LAi8Um8Dey
hiIm7Hx1+BvNEBgfsa/Ztw5/ypQvhZp+QBDrs0DokKsdR08tMQN+bzjeEEMkf9fWXL0i8QD2t4e9
awzhNbiA5stDEKZOUP4yOaFNUhBtukiSx1GN00yQ/J8Rszk/aIiexmClhn7ncKz0bUXUWB/8md83
5/YfuWfC7Wx20RM0yCM+Xv9+kzybBQx3MaLibGK+qM3x/LvL/W4daNi0YQaXbwkj9dGMDXrM5z60
wWQORZlPj9jMcwhV0bwcWKLL6U/ycBDuJK4lnuaxqn2Zk+kjAYIsQYSzNbUuestTX8XHrZeU5VaO
fuLGtewQpgL+F+w9rLNpnxW7hBnZbRKADWv1xvLkmZKDsvrudyYPZ/dzDmCkOifS8+qpqFozVl/b
veRtnC8cbBbl2RxTEG39yBAl/VumQIcn8DCbadWQl5/brYq1XXjiSCqqtSypV2zWQKc43jqdjI9i
Ws2w++XYJeyEzFxDz5wySO2ftV4yBCeKsuOLJFM9qsVt1zzimxRCpSAgtpf3AHfBV1odlMYP7GrT
ihNJHzCw7ZwMigvCm45A/BQRIjh/i0WwkTBUR+PJEvyiD0t/ULy04KCGW8kxxAAONmFLeuVJuCGo
UsXyzhGeP22ht+y9KnDUMAk2+rCQ5CB6A/zc/5F1KS3I7H6SXvQsRoeFFlPflPk5rtsrN/9r/CK1
dSBA1UhxcGeSN7ZZBUMNV9Elae+xbSJRRjEII30laSpftUlKkTc9rZmrOoAtTofWkvKc57St6w0V
1VQyO0XlsGWWLP0dkb69cangcj+CVjt9WzVPt1DBzxZcNtM63O+Xd64nPXk580OniH2pEWmya5XP
QexqS7BHvp6f1RSPFijLMFE5qiySSO0sVg+EaHdEOEr0l7MPPUuJRxkZ577xtuQlO0X+dw0b3VZY
cpvVF+IIQ2jBuUOo2zewdtY+cpCR4cIIdqE6KVvRFnttTg1euxXOad2ANlDjzdz0YvQgDYEp82Oo
RkMr6Y8Bbz/3/wf0m4VC+r4etkCpZEIWKysLbUjyl+f3U6e6x7H1Cn7xMN1mhRHIkesCRPy3v3K/
5ChjpLOP8nUH4naCMty8qnpiqQe425UK9WSdX54RzYmOvyE4eoh8hLQsT3pvu4pLNpuyq4vPuv/o
LCGHe4PzQk7lCfbIuhEWlw0TIoSnwS4JLmvbRG9mVZ9i+KWHbxLFi3qqzQqwEgzPCQMEFq8E/6XE
70NAB1hfMJej5s7lWhAD/hjfrDs6AOFjL8k8LRcadKeiegaX4fycTxzQJq8JX+aK4q6y8lBn4Og4
ypel1vOiI8FAH87/B5nhHyjwaQtIC7YoV/0CAkWkio2wc0dQcw2HM1HIPFpa5Y6nU6Z+vnG2awle
bHLaF8e2OHw8Zmhe5AoPdT0iOSa2LawIsYSfTPtPMcGbUuy7E8bR/Yy8L5VSVLpUbpLOU3UHRszp
SoIcnbz0tHdC7Ls8p3XTw7Sk/L+vzVwujDcd227E6eZ9d/n6eurVsmc95yYzSfz9wzUjCa/RANas
fRTXqhqyvvcRs1D7HJhutgaHLc7uLkGo/uz0kqJdCtBBScnfHVJ4vbuPFuh9yfsW/WFspytHbSx5
VzCUpgdu8DBZFID3HqCf04rou915TWdCel9kGMdjsShmD7bWGTdNZe2If9yFyR0IqCaK2hSL2ks/
e/mWVN8f6EOIpaEY84VoSqUF1PTJdOVV1u/QwGjBkwNI/fjZVlToiXq8ZZHgbEcqDEvtodk8OXq3
BZ8iSFFBYUK38pwUPAOjdr+rxXqRTe70JHh1u7BK29sPYosnIy6LgPlrk7yX4FGIK3bW/sxj5fiL
y9nJMdlQWeLfQ2vnHVaoP+8Rrk80mhXjByXSj7eOmwQmpHk9YwMdmiRCa2QfjZ6uIGuCFr4Qinph
pn5+80MwnA9GrFcvs/mEJkdf/XppEolDfDhOEbstCtUTAbrwUqoc+nuhQwzAt52ESK1mYPM3ROxZ
ZuWNuarHA/z9vf5Ad+91WY1VNaEZxTm9hLvscxK7fjeXoSX90OTDfpFFpPadoSLId3lbCJgIHIci
mCkbXLxPDua6cZeJRJXhJ7So1TzuCPN2JPc3e/V7wSx5iYwcLYy+ZXewojM2yMCcXJ3IaDpl6aEg
+NEyhl13nQOCg0uRi4jl27V+CnAupldIneTLjboHxDn+wf+ZpD/LUyQSwq4woNUUftYmQOiYaQZo
orD4FiTjcE/LGfZ9oR8lcbA9QJxRWXipA9QjK9jnn/qh0VoTRish24dotNdE3VUpCgPsYn8NC1dk
DGan8+9f2V9B51Vb3ElIO/65NFfie+36lU5ZuSXCnjGt6MgjxJJgKjX6ozChb9nIt5jgCXsbIAmG
LtVuDoWHj3sVDIFOEH5h+o0lTPEs7q2oBroqaMvRJTxvc2Sws0G9XCpWHmEGW3vjGhsW8bS+8VtM
TpwZbDNz76kt2UX0bfTQ+bYQWa00cVWlRuX+/RKWpjn4IdRj4WAffXxiNIwwTWq9299oGF8dV1Pr
blPpOJoIR6XbWRCtGgravYAxYpsQ+yCLHdYS0vB+2S2AlX348qbd4N3zireTcdw/nkJ+tN8fd7kP
N+W7ufwBBE/7uxMiOj1Yyk9j3IOXhGP2r5Z30eKsBJRoJ4leEJFwykkEJDMrMAZPch9GlXjCkJYM
p5PAsHhg5AXCayeByjChP+4VJeScF6WPlyQWlgiBf/fqNNVUJ6klezmqSpezRnYcsmojdZRH/f2b
kGxC6IFp9EIg8pRyKYmJ8tsm9Hf90O8DHGPEVVI3rak8d/YP6amZaGj/TwVT0I1LbSe37SGhVXhD
mXpepIWgNaxtLg7rbVoBVw885pC3dLFfWqx9Gy6hHbX7xfQ1e6saUWEozEHTSU5MNTYTkpWZqhHV
4u2MjwXK2LNiXXIoqiTCTYX6p8HRTr763A5/xc4Sp67dULOCIm3yRFX4EuP/F/LnjG51S2sQC5dQ
vsYKN5mHQFSdAKHy4fmf8HDTGO9OzP61HMQ9jEPbT55+rAeg4vjYzojwez8YD2E73iY684aiKZO9
VXyWWl7zifP9/cL2foIUMOcFzlm8xPwjLWJsBDiB20OPPNBk4qAn3HT4DMOzG0MXQZacaSh6yz/p
AvJYZysHKCUDdteD+CbQsZV3FadJUM+H8btWJXs/THIln/r7kyuczj2GkAZmqsKR3duUVEUmSsiG
FXhyTwOMVgJoVYp6UdUR/qPr+0weVHCiuid+l8iTvXm9y1i25cZVlZd/iCLao10fofA5k8bjtJFW
J5op4EV84w9p+JCHIxaypzGxT5L9+3fP00DqFjxnGQmcootf7aGtizR9ouCInyHwTFTCvONluHgt
517HDZz3GiGtyHwdsWF7/CsAoyIdbggqED/HEKI6LDubKl/mWbH48/ohim1b01+Cdpa8teYbgU0N
j8rbQCjnQlE0n7Eoqkrt3SmDbfIYwndY0P2eQ2xYVF2C87N6d62n5fK6uoXOrSILa/fpb0tc9ybd
x75e0DJC3IVLrnq9t/j9iFUkLz0SL4UKX+0ZoADqRwvw7dqYIXI4RyN08j5aDIgqE97nMSZpMPJ1
ckS7mCyukzccCYdscI5EaianrIL6BQvv1RfAwevDmDLnSuuNV0ecXoHyLqParwDMG2gobXRjPLnE
yT1G8ysNXwaEdOGQ00YWKEnfaGEwGKwbOrcilJ49YT4+bCTf/E1KnEaqauAy08jp/7ygCtMpr/xc
82SwsWgp+F7Nt6be+gDuTiXey2awBPMrIDIQ3O40quAlBiFYv8ktewIesRwHi54y6ObgX4JmUkUB
yyGvlkJnqGwnnyGeI7utxrdX301CLJdKbNXotu6t8mSp6s1q56xL2CK7319+TbPGqdDG9n4sWTnP
02TjVeiaGLNKz6lMYNEJ0Kl2vjRBiMyH9EZT15NxKr9R2AtnmK1Z+xKQ+chX02YqOHX11G80tWZq
dOGBe84/KEMB4d43gyigUg0oCjIC/UUU6aII6qJ26eZRJLiT0ybC6StrcF7Y8UteKy1eYGGkZqbj
mr5mUDXX4xluXWUBNyLY/wfnRnTJaiql11YOc7WZJxpNHURD2VPmEs9y/QqT6Arb1kUpJ3iXFJLj
CIoClvIPCUEPKl2tGyVx0g7FsK/oh6+zFbj2t7z2iTj9L1mbbf3buPbVIAwGgsOyPh5U/bEf9Rdw
qKNO/X43SJDYvli1ShVyloNd3X5wajF7IIZDelVldbr1Wen6BPXbw2OaCmnLUXvEMS4VXCq91cBu
uCZasEb2o0elhjKlW6ZG2isSzpf21CQ+YrGZ5readLz4sOiStQBXbQdHx4/QGVwq6h6rBYWKhBTs
/FbSrEmjnz137uTewg7yKYn5B5AG4FYjR/R5/jWKHhMY8E5UFleyH87jKYleYRkDOexQIucJN7ND
4PJjRJi6Yles4YXcBezReqlIsIsCrU27+vfzeIUvVAdvx6nWvQHm75M6azxWy3XLC7OxJJ37rh6Y
vKE8sgVZtx3o4V0uZepCsO02gxsXuC+OmPilv1IxbSjk17T3RMMaqZcZz13+glmKi1Sk+v0d75QB
rtlMuHxw4kiy7cbvrFtvWJMth758kvxeft6L8mVMOmv+B+ksEoRAG2IdvpZH+JbX+Bn/Q+JBRy3u
xa/ECWZfSZYtCTb9syhtn+XuUx8m/6g8obDrPpozcEXke+T6a6Pb1XYcm/p+4kanCASpEGqXYpcz
Jl1lzsVJFzP6MtOwvbj7nVXS34YQIT2JaEzgXbGyFlo+3BxpgSdVimkr1BHm1B4i1LFBrHRcoCvm
waLd98F77OB64c5TZ92HPm6TMQpwSR0w4tFkwjTxMGzYzs3ove6gmQT6iXhV2IlZ348Qv7SCHFZV
qwwH8BeLh+5IJl3ldpjxLIl75nTmxt73k8oDgIHi8o0d/sviX/m/KrQw787zEwyYpKE9r1RFMSV7
rJWBySstVzoDqNzv+MmozIt8jaF9H0SUuRqrg72YAM2EvFK8NfspnxesbCP2Qafvkn4vuUZuOTZQ
0Yo8MozH4wUQ/qBFCoz4lZrajE9BCgmu//nQw9DcoDk+j2q0Na0MclpK6HYZxTIBzgRVLarmEi4X
HyTJwasreSP9Q5nP4Pl3Lyy/K7VVcwHszUMrN8hKwtghBEmbK2EUws8xhYhqr/0v+rlbVuKj8Qw4
Hn1lGpVYV97qROZrPS2To2BhttlBoiAVgPfKDWLbng/3dxgejhgZkdAtR4VYdmuljdX+T7oXy9k+
+QgT20VR0p1LH3LrCIKRptDIptlbGYgCfeRjctTWRkXFEdlVUHpLw9fHeokEyK+LB2QTP2fNyZzV
CSsBuReWpdbme1gq1SE6NQph2E8WI6ZnAOAXfYsP4LHpVh+HFeW5gsBXisR7Yl7u3X40nVy1VZHj
VhlXi75FiGyTZRjgiPW4h8L7O2iSztN/zEglSs+QSAZqpFtUhur2V1tRxRw0MA1kW02V46MXwxgK
P1PLQMch5tyjlexZdwXhKVElBTUkMq2H55vNd1cm/XZINBskSe2yd9x2qcdcQmBvzOe54ClAa5ep
2tJfmGV9PhEg6FWa8g2fXQbQd8+dXcCFFbpIuY8m8qbdOAcjNVKatOgMdTSjDeJ01jsrfzShkpSk
r/X0zZeAjgZPbKPCnevOnh1Y/TR/ym7XrC43TkvYmMlcc5ByJw5t0UEtrb+jPIP2WpbMiuEbkO2x
Xc2o0upKLh6AwU55Mbcp9Og0TBbm4mpfzO9fAHye+YpYmOaog/AHecRSOr/RPy4PR8YKRp2xEI1u
sHIjVCkLrueHkXE4Sa2Fz3kP0aczyWiKbLNSBw+gDjs09g/DhAAGL+DkbXPgTiCQRMaa05WXXLPu
C+QOT2DxcpNfrEhei0+CdS/4WLxFyIE6+VI0F/0VTaOG7HCeAYk/vx1Gm0+3/QVsDRLTDmzC92sv
bSr/wPliM96+VwtAxW+7I0iRrtorLZ5Ni8xlJAtPGmYZVu8amlTK/iVEigXT7hY3cGuDLxnFz/LR
urONc7oh/L/J4TflROeDgod2Kq07lWXuq7wuRTzRlubcwCD80T9WgZ/d8+wZqaI0MJ+LfAMDB22C
7j56o8+aNGI+2KNnCexgit3RTYqT+tbv3ZJBSM/JusPlPe6bcP45/gEd/hBTx3VdCNc7tL6uJY+P
sB4yR2/iRU67dv+2s/0J9Nly0T25wRoB0tZHAU8nvFGruNghhHjy0ZSrPLgwcJ2AFUtFaE3H/dJn
TkETOgn7yRt5irgzneMbotqwhvUMXIEDgvkb3VAQKsrhA3sxWDC9TmSFAODx/M39XgRaaPBjuAwx
A6ar9qT63D8qBAtjfKUlsfC8vslWUV+bFjMFbm0Tz3Rd6wE6+BpbLV6CfrOo4oe0xqj63fQpUYc/
ZiT/lxFW7u0V8nxxrzv4w/MCwkFxHL6gZB6SJs3zDZrMJKnOQ0L0yzqVPLhUPDv5HoFs3G2Fal6J
dTEoni6szL0JpQW/v/qbp7LTAv9pmHVJjLwxAm+2Z2mFxpVX2iAVwNNavlYHebs4EuWHJou+ljPk
z4XgNUoDqawwzNzMZGgcb4XAE6EeAmNNHuxZHPGuptRyXWuAahL4t+x8fcpwWKiwGT+INQFjE7FV
I/l7G+su4i2LBdwB0iFi4Mmvlnn2wmMiQ8L0CaxuKc4xMxyBR4U6wB8qBEuqQjFLQ1h0sRikXvGK
ENRKiCIEo3UrlEF3LLz87O72k/EKaG6emAbUt09DhICd474SjYUhnR234Jg4R1T1tciseuHNVMk1
UA1xituMxAwB5ZcLlnUusmy93s4WLBxXQi04wlxpxFqkLp54+jX5NrZtPQJjq8/3tl6ZE4PVyiuI
KO5HoOhjwFWGMCC9aZjlVgCsqp+aLzazSj4ZdwNwbN7rvA1VUOc2BwEC6CzJqlp82akIfoNiewHx
RzybFjtOUrLq8OHdlZd4uv0Vp475IGRy+WwihDpGsulX7X5FjBaZOwzeNjFg2Gh3UdINs+YqhqM4
MvCczuPROn7b3sGXgIraqgYtKc3vUuKoCA/GxFn+TuflUYT+BoOUdamMy2IaDcPRmflKsw5im1ff
cAVM0AFuAJjaN2Pi4FnZdM9DZ3iZd3v3FPjotPIsLqOZUYom+IC2XSsSLt5Fvb3x/u9mphdVHJBl
ckvsX9C9ImfT7cd0rSEF7Pg2DWD8Efa5CBec01kJfhtkzMeylsOiimYVfwRBUlQtiDjTQEM2q3Oa
tygNu0y0dVvbtgZjSeq7X+LE3P2YOuhFgyG0Re39EbzYUWKuXFT8tI1Fpmn+IdcLXaFWx9xq5a+z
EIqsDaWTZiw5kAn8iqs3pOOVzSSkiye7578Zo3ktdxWgeNj28xCe+SURoIm5gz6GaH6dtsyzdsuw
Lq92c7r4Eh/4xedMYoqKOrfxIYEvbpkMDez5qlxnoc3tlpKYywS3KQPyLQYZgF/N5URQqe84BfPw
E62SgMByFvCQBBcYic4tP4pU1jP4vtPQR7Y9ejdxIqJ5LNX2T3q3UnQMEs6IwotR6x+50usvAzF0
n6/GjASOfwXTcGtBsrB5Ttzr+P5Rkh5SD/s08t/o+UC+UXg9Jelz4HOkQdSyWm7I02huYM61/L2c
+RMIgLR/Q9G0QBiq0e/IF1MDFHpt1qy+aIbIW4MEKQfF2FLni4UTh2/zYkI493xr1qh9TIXqJczZ
QprVMjg4kEZpZD2oU8xJ+QJH+EH3VX96y99F6T8ZRu6fKYOKU4eE7/1vc9pcK6KsXrgX2m1WzyK2
ImobxCyYcHbbMEfGXuDzQne7G3MsCrUroJDFGBYfNmnKynQQNPTmmZRFYNKSD9v5seBp6jHXaNhR
HXMaZZxkB23z5stQAMibhMc5eE9QnOhI3bbMOY18xlzkLwDFbPPtF4dOC0KMFPHL5eQMPWRKiHe2
nfmI51d5h2nMPJQA0gXI5mU313IO2b8OV939B8bBC1PhYRIlh4M7Y5pA9045yDk2b3yTcamWRvEL
RA6IIryn4JN1SlBvdnkQbpCavw5vDevPQ+nE0BZDesODZfC3ly0b7TH7tKh5u2ThtPsBAY2Dvubp
NKbwG/dHCh9mmD834IorSXYe9OUkD16TIIhWyaLn/jzGpnzX2P4venTf5fXDIi9b9TPo+hCOT9UD
kEnYK8FiTWw15R9WMcwSN1G79zEFQHTC85RE51/NbxrjjEPlKxjcF1JhU05H4DDxJwgZXU7av5Ub
fgJtCROLjJfaO6T2UOGDMEky1F8SV6oVWuQKy4UPEjeMHG3JWYHftho92DyfU06P6DZQ1WybFWir
uFeoTaY4Ggecbcg319+uapitCZZd2LuIGArRwNfpdOasCf1iU33etU2WD8/DHOWqgdYteY/6P5mK
4OJLkmsBMexmzGR4aKyCqtVUrXttcWOmUqFVKd5wFFNK8pfoH13aw1WO3ve1p6uIdtqIJ8xIzKLN
IHhMntfIgM1lBexzxap7CArwm56PqrCg2EDRlKs0lp9GiL2nzCxQTyZosTPLn2/a5m3UUYpnI6n9
jIDtwG8dV6y3UGZU5nktVb+apPSBc/pGJ11QFGSItVF9krmx4MhZmRL0wfmzJXj044BFak0ieJG7
g+hJA1IO2MMBBmkqSBkhs3i1sQdL8QQbve13v3Zt8AO2uowiV0c4/NncG81Z4gS9CY1BLXAmmDuq
xrjVlrD0EYdU7FVGkLPwGqnLraf3YZWWDzdGH7+VsflfigH4uuaPk/kiLVC1N0vHq/l5fx6N23Za
hBRgX2SXsqvYMhWHcwAnY2b6lxO/KDF5ExKsC6sAQBt13LJrBvYMkmztEOobVpu/QfiN2sUKAchF
NWEes7JguTv+xpBmh+PBaYxyb3pmACmPL9o1Lq4GLDXALINq/4Tqc6YWhd6tixdUmuIdgxd38Oc7
tfyfzRjWac3tx062BBpiidMy971USjwGyXF5Jyc+ptOUqQtRdp7KZFOERqtmz15B42zCKtZG5Ywh
CMv2noHrHBPEzrBvQr/Wdiw/MZbtLNUi0cwu15xH9NtM9NyXMgpkz9Ci7WUGOn+EbDGJW0KkmuPq
XDaQy/aWzKyNVUI90TVK1yqm49pp4rvw2Yt0akx2wvtD17WJaOE94zKXm4tFtzjIlxhPCvE4vi5g
h/yU4Tb7E1m38+0KItql0C+Qc8y9cgaUCPJM5+q884JJ3aY1BIoJJMEFgrE4HNpjOQSXy59GkfZ1
DVNusdSBuoxfW/osXsMA/ubn07OVDYYhQUPt9Fkr5rGyjB9PivXVOSEZPHG2N688wJLwNiCKyH1h
lPj6OqGYHJ7Om9+tpCH56BnT2wQB24TaFwDDvvYWPt61pqksHlS5cD1k8WKH4oYYTkaA1fOIAg3U
7jp/BFo/k+H7KwqKIGyljjZl6G5CF7WLBv4/cOjOyJJiNfZna8t34/C04f+AklLD+edlGh6RbUNR
3gLOnAU0sAS0YmJC1w3Wj1qbxJa4GqcBBBVZAJDJRzkU8IV9D9AppD9M5kQLPxjlb9IXbXPXLkye
HfZWMrlC4xqyEZeqOZQYDBOcn3X0gGpS6+2Kts4I5ktrUHp7CK4kibiXnmlcTvOsODWkhdpWQfSJ
bJg2vInDACxtn0W2RF+ib3ORVASO7VkCNXW+9Bb1GJDui9c4v9rRTvh8lt44Tr7RXlvCYqndhOb6
yjRFAQvKiYwjvQUyoRZavuhxxF9jHa4lN5HCvRSw8QB5B7EC/D5cUwuL3OwYHdVFvjW/bO6MOQYy
Yd3Qzynek6PaimLiqO0VoXikfXkJDVWhZKKCxdIWAGQvYmCrB+JIgg1dchzILTij6hywdrkrsAh+
W1zB6ffG6waAE47p1AtQa+tI3wnyQhkpWkyqVTRuUD42vDu8JRMYjQKXE8SO55ba9KRuVFRG2zjN
Fodew26WCJixtZ0IJtt+2kQQpPey6c3U7Azo0kX3VVoTfVR7wD7i+5UF480UcUgcN69KMNzUT5vd
5ZxpWNRmd13OwZjP/+Z28V5Ti+lBSPNpf3bAa/2iF8EIr3Y33H5mnOGa3gLIo/lI1npjwmnydfvZ
C+dEnqWnyPTyPvK7yiRVkHvyoAlMKqyuF+6RChRHxCQg4srY3RmPIl6+JgHslpumocUf673EGcS2
Js8lkHl9wC7YSf/nJo67Uh8jHcR++1r1AkhYaQDspwCcK1ndZK9qyyyVzgBO3/b8wt+s9JLqFOhN
1DUZC7MroJZSzOR2J7WhrHoB7amjMP7H0IHTbUbzsudk7vLxrsWhPTmHRw/i/vBJ0SeokffTqnob
uTXb1O6gwB3XBATyvZhrwfx4uV5ExJ1hvpeqvZjyn1Dm7Ap7L1Qwb/enjkjnV3ol3Db33T4MH684
hYa+4MDkJy3JDuCNWpagBnd19b7lMklD9SuM2JqY1+KBeO4yv+NKDnOR80wNfpP3u1jLA85cP5L0
P7i8iVjeBz4TrWP1N0C0uoYaqN9q7WibQv4MFAwJLp8VpreDoYxTL4YLW1wObFk39aL+odUWB5gL
lRvkusmI9JM1uzsJMleFjR4ONUIXBqNEq+plg3d1YEzn8v/x8sKFh5RXd2png4sz2qD0SnfJsoqi
dIE5fiswZGgTvews73qIEVB3Yqhm41dsbDu5jkS8Uq5PqtD0viEGnk6eiRBvYhX6rLPrekCWDcFQ
pY4zmSMX8G4PaRT62CqtY1/2oocqqbkaX16jUmfkwJSittJa94zWRyIROz4jEIELiBYsLfHn5UEK
vvevE+7yxzM7pf4OcD04Zh1ySVXQWEeWuu3tepgj4Ay2RznPxe7VFlg6BLByn8HbMQtgRZyKRL8v
Vi7PjqxqlPuNnDC4h283o1tRXgNqdmeuEfXTMLjy3A8S8nzYykYoRNc1xsDSmLNfDJ6XQM3M7ToZ
0u01GjxvIh+DVm7+DUzqdR87pjbx08HQWVrzcgUnNKbWJzH2vhV5SnwKYIWlDdn6V5c7gvzAdy/U
MruaB306M4/h0d3I59IqKOshbUHUYYtMerbPqBNnKDxyS2ADTW9scSYiUQzu9RBbbttUTw0q+j+w
2wf3a43R5UKRy8N5jPLWc7TmOWJ5Q4vxUNEQMfcq9ralPtuqmKzY/B2k5arEkIKUiE6nz76SwduF
+rjXSBrv0gYcoZqZrPgbBtXHyf7WSJgE73eLrDDeTEfjdzhPJGTuPl+6sqQuwV2z2z/mRMXrSenb
MKP+fBb5jaBYGyEpZShYP9oPP5v3we8vw35QGnxaF109WKR8KeZ0dPhJ/RFaLANHn9ubgcjRKRee
pVjdJOIVc0DU6QCEhJWOL7/h8We4q7XohlmLt3Lj1rGkpoMs4HWo3nZhqrhVyONIRaxpRCVP24ZO
eejZXpaeFfjv9qw6aGAUq9qUXX827QV9bhf65fN4bqfim2NKVXL9fg9hzSRZqnmsf7Q7sH4e/H6g
rbkHDTSSNDIb7EBnUR+L2L5yEmsgcipOFjMoL67DSY19+fccI/6uWd6sehVuUwW8DhaHK5NjKlSo
A3HXQmtBP1XLeL4B1gNB3ksKqaxC+AW5IWVKZ+LAdu88z1l14P8M006JUXEIl+dDB3+UfFMcxu/d
gIKB41lYkyaCXcmzIh6+W+eMNC7kdV3TnMMeBP2UgEF+Ug5Z+JFECF8bPz25FFxCZIQFZmvb43kD
BXG7uWy4kmflSXD7Su9ZbvWn2h00nZHWTkraK2tEIFnZBSjimK5nafwV0wYURsW5De8RnGIVkGM4
CE9ObB1aiV7iDVnyNQYzBFGJIEy025Vf20gEiq1md0FAjrT1qcfOOso1N3stN5Wk3fkOAH+Mp1MN
D6/XQ9pJAbMSjM301nZqbgUl78XCuempQT06rcy23Pig9XJAKcvhFAWXI89SX9l/6ryUU3j5nZUX
8eUZ5XkFHX9CJjfQqrMTeHUm60baaI9wOj8z33AsOv2XExGEgx/8DTToN2ZjRIH2lavKAMGXMA0R
2ULQ+kihLzep+vCFbHndsuvApcqGuY5fNfJAKP29yZhwB6Tgax9oAJkPR16kC/e1kWLsqtsxWaaq
PRBylb+KZk0yNiswa4LXD0ghHqeFssj5Dm6ss3cJmhxLz2RnHJ2cmLQnDDTonNvM5tbYK8bHJsDk
kZOloDg6ysJZUu0QzAlHnTXSvc4hIdkw9sjvYTGtcudPsSF5Nk3pL3ukstMog/9pcBlsuFX9AO91
FjlT9LT3i2aFoCpZ29bpvAIZgF1QkklGRjrUYguT03Kzb/lRPgl3vm+bmjFcrVYUz/hgPPAT0na0
dkptwbv4x62cTSRTTc35FV1p/1A52K6aAqvPmsVlhOs9cQl8FowzwLVAYQbKAbseaqN+C3anLIlg
5KiuI4oiO5Y4j2UHZSwUhRd/S6GlwKmWUvtetmL5lgV75OKFvIMVJyOX84oq/q7bYXjSsy9p/2QD
sVlt7m73j4ZRnyrR20lpMv+a49UC5dubq/+fDq2wEhGfXv9LMX/6LUlvlp7jgiefbmhPXbgdIOjS
MXDBaXsF0/1poePwptEyHMRRLq4kxOm5Hti1RcjCIIxhnBnK+PkqSeAom53fpLz+pcjK/+uedUi1
z7ciOjI/GMxMslTiZYDjR1zOcDvqFtzZgj56ZDoxf7w216QYO4CyFU0n0xzPethykUnfzpeXBdCZ
pYNbMqx2X08PZth9O2xX+nkObF2HujKlqNxA6hqPC9iH4R4zS/dHBKHq2LoTDfDG6qw3SuW0/xgX
gJpydrJeh4xfmEadW7zjAaCo1D1yvDzBceNNWCA4h0fMKRhtsLqMsWVZVxjSG+Y0wCTRVDpOZPFv
WJrR58vrf15E1oMnSggmyF88eHDhYH1MRvcBHwEh72gtsQuNh0+VzEvhhAfEMB3uS63cFzRK2jM1
8vPvFFE2Won1T9LUQdCxSKv+77q9gT7AavMQrtteX2lTlloKd+lpMD1c/g9xe1TPYaksfksXSUQS
3YS6hvBkksMqBPX3Hp5dnSWaVIcAMn4ld3vYE45tN8FKii2jKijxA2RhJ1VAibmwthnTQOwZlRjD
liUEppjQZWRGCRuxDA6E8X5cBFCnDUo9W7mGrr42kIau5h1qrIRyE7ZBHiiL1q1pYv42pF5UWy8q
YXfIDMnMshXYpuHlRPquaYqTUDazAVOc5cWrY/eDOY52IMA3TkrY19yCXNnpUtqOE92v4HmBEnOL
KOP9sZJOsByA9dVGFT3IlNZeRnr099IcLul+Ck3j+ke77QZzmy3UxRfMLWMXJs56iY37I1X0svPw
ZK7hrfcTfpV5P0EPvw/p3UytiAxSovOsFMwt9YdjH7MU6+QrBKdydPmHCxBFKFmPeqf0ghG2qiPl
TSWA2Mf254NgRhEBa2NSgzR9U+0jSrPQmyglCYMCjwQ3gIV23hIpFM3HBgvg1UsnIywbmbJ8coct
9FoCZSVAT7JpP34a0Hh7boJ6scSaXEkzPk9Du9p/wWU0pTSIAjmCJxzmtJrxgFYpYNjD3tdIyEBH
o+NWq4gOkG03D10Pc0KGiAXOWDGVoeJF876ikSThFi81qZRxrr5NRtW48c1J1ztEIXiAmHFy5Yc/
gq4IxXgqmleG7Cp2H4XqDOB6MIKkvcKaDSZXZn5+7hHHrvnjC+SUObroDkZbcQCqG4b2t1ndRPie
wwxNcenC9nQHTVWwVrRx9hN6GjXDdJOu/CNVXzG6O18XvaUnPYBLDAwB5wtkgelOsDuJstyZsBbU
JdoAVJj0iabrw/hlE7m8WoPv7T395bsnHKIHvAz9D0r59UCuMGvuUcra5gnZFWeWwoEpkFcwzhVo
AltytWb35pHdf9VViU7BVORP5NbD5eVxv1/YPxBo4TuQM9nvRprElRS5mPrYHxkGjX08CVaZDZqc
6WYwZeoxqXt3yhqb5inCzzVNSGQkFqk9qjdcnPX/xhKT8Knicc7n7hUZBgt3YQIFad8aHglqTDdX
jGx+c3r/cwyt5RmLn0ze/n2qsdrvpFMBKzERIYkDFaSvfS/2uq/UyBcMdkz6agVj9gXJF+II8SEJ
wcD/UanYKxakBc8mCWJfObCJNKet3yGxbFI27laqFDlB58ofR8fgkuQFM6mj/v8B+GWzZnjH95AH
z/1hwqzYMUMBOBlrZjsXnhvtqPrTzstDY2nScWdf0OVR6olTSU/qIG1wSlzpZlRVR3/bbJ3XUUZn
EfUdGmKr5D4Ro0CwF7rdb/qg/PI5fVatdzZx7i6uOPP9xHKN3WHM52QjA/lipdOmfbyFvPdxbW/R
nfHpSVJ/vAVmbFWsMe4hkCfZvNRLoCWQLzWmJ3NJSqC26ydIiMYL9NZmGwMSqpZW7ggG6VPZHn0k
K0N0nV97NrvzpT5SYNXmPd75I6V1NpkZQVdFzBvBENGFEFQuCK9h0LcO38Aycb2bw6bv5vZi3o6Z
nzEG6B5anlCWvCNF4+QwawZvjmVe1Y7KyaJ1/iNsg3nAv4FbQ30yi67U2z4kXDLvLNj2fWhIdKm5
WtvkC1umj+kLKvMI4tIBoNoZuVMVfH811HSSCmsazQHVf9cS1hsatrgdFUyPnJu9DHJkolIy80jb
osQLvOz3ORXT/WIN3AFcijIpTV4a9n5TZX98c0ziuvQFqVdc2ck8Hx9VyrW2Gq381AubWhDihZ50
f5Q2XB8UbL5dmkaYFVYvoLhiQI2Z/DDggXT/Wr6jQ5a2vu83TZcrYJgt6ROLG65Rr4htBO/yyLh1
z8ZTlCgMVhcVcZmkL9W8JYt/hFNXDp2KndVgE2v4rpQdnmRabLtSWb51bEzEahBp6pS26aQi8hBZ
s5UVXZykgeUI3Q+IVVQk6hMLW0zE7wHUTQKttejWNhOiUY0dqhILbk3ukVAXXFjj0/DMY7JgP0zd
SsvkYX6IrPrUtVL6hguAYEhUcGbenmQlcbHuEifZ2uZ5MY41ZVY17ekdxyOD4WNAhx9NXJNlKUCN
xG430FpYnkkb8tcewVTM5XICIZ/gxc3Ev3g8Qau+jJr1zB8P/UiYuyg6H7fq89M+qgG8n1zpcgmr
V6wRkrSvTc+6PpzxCUgQO67fplDVydrxOpne/813//BHWtJxUWBmTNWyJbzTSbGjuBp3t85nPE6/
bbUR2eYvWPe/M1dFEZE49vgdv4wclJ3mUolcRhR549UeChJdOkMvM2zKRROmgW+dvHegTLRAZMj3
4qUF/JmfXPmabrb2emdqj63P7VO+yRQbIjHlL3xFj98ShViDRbkB9hNAsxoTKzAD7ybO3jbx001n
nMuV+C8xb/AnFiM6ISPQuOLec0EITPZFkw2Ye9GM9PH48nt9yQHk7VxaEDSu55YhYx+Vr3YyvvLt
5/BA+/PH/azeNpYaaEWIHHhdnRFBfatY9uYqg/9nU1I7Z+qcrOinOFLe06TV57ao6EXPFz6wtRpc
jr6gL/bXySMAPy5J4mUyVs4YPVbQi/UfHVbcYNVoXI98xsfQTn00jeOX1QIO37kWYDTFaadby+fL
Kxu2i3aKhxWaI/vndIWBvtSxUptZyJ2NfH77dENHMMZmQeVxYDw2omeAG/GYq7wcdKzinbI5juO0
QjI/Vqf6OwTotF2HtOBCr07MO5vIfCY6fLST0BnESFDZAqvQRZ2t8zbq51SN7ft7KpOq1B9dIJ0+
rZogx2f5DtZmA2S43y/bMshtyC42Z+ph3H2Knj0CQM3EKAH2mrA9V4eScntXcCjOqTOKHIgRHP3R
+sKBrozlSy1QBnhif2LVRM9TDAegSjLYgdEo+yGFr+Vcx4gj/Oj63fYFdUphCUzQVeUTQkRzrSHj
0XbvYwIs9n/Ev9gr7OYYG58xsfY217N5LCAt0T2qI/o+uV6Bx/K4tlVXsSp1FWQoTIWv2VNUnor4
UOjCCikOmzNx6ueLFuhI5mCQpQw8Gz2o4u2kBNE3QDtDSv3iW2DfStvl4fINYbfzBY7uQwwMIHbD
r1thjZww8FtV4rAJnXWTqhEnOiQ6iIdm8eepCLRucexZwO2pZqdmph6DZADJJCvqyq+o2df+GTR9
z4QYwaD9hdF2G26zYuaqzgCfYLPWJ6EJFb+0VKl6hxz8IqhDHAOzUCOWZxPsmeb2pm1ZAnmHqD5p
9xIC3DMTEWUC1eSuPFYN5TOVv+ixKNK0txzG3v88c9zjkJdL+7QnKpe2mP1SkdVa0jQamZoBr8fO
G9FPiK6Y6OwsTl4Moq2lgrtmeZLsbzQQbLR0k6ez7beSwE4gXYSeZuIvN7VKIsGp23OOD+BldeDo
9k2hPpT6fNvPi5qKXAAr4kECcKQvYEkbP7kwXsPYrWo6Ppuh5s0tK9QDpxmF12HzSuMusa4KkbLA
PWsdQXMqFKB1MWCx4MptDngykRYh6T0NxndG9ICZyjkC7LhrqN/DjSJ44fSlNmUpeVY+2WtL/0G9
f88aE18Bt2HDcvbiQuUbXpXoLClku1BjuGJ/vK/CofN69RwocXUQxqO/YttFnv/QtebTWHPXM8cR
ZZVX1TqXmvZx2Sf4lqvK85UW639vF7DvMiF7uymUFMdZGOfE79fvfdUBIcSz/mr4Lj27qdxf+wWz
Ku+QtCN61/GK8+p4wRrz25wN0pWHML2YrjrAVSozK19NeiJqPoECQZCl2UU741/uhd0fmOh+uswp
zkLuveucShff1Dj+gfjQ8rttWP+k0lyV0Tv6tr7ogCx744jrmt8jL42NZ7WI8pXBVDgS9pAgVD4u
D4J5WTTL2h3dy/NOWV4Wzaf2DS92pk43eSaNbcLQWgE8jpw+2ES2cgQsfHlod7xMcXLaO+WyoB+f
MHNP9FJRTRQdaVvyaz5nTItqn/+tleMCnXFtn9RcDXdXxTVTnuFQnFPD75Qela0Iduem6p78nILN
VMeHqpE0kAXrVunxnf3JBV01Gl/79l0rumg5yKWVDX73/MY1J2PrMZj+8u124g8tzuWprsqmL6z/
2Eng10/tsKnq/S8X5+wW6AI1DQoEHzVu/idjqevZ1v1H+yuxz9KUsUQVOgUy2PvMOMaagx1/5jBr
Qwc4fX5CNaQUkab81QqWDe14xQ9wjKF7daAAy23OsYGKOAlFY9huSC4TjVTuemXqQce6FLh7gBtj
BDBFzmTVga0juy06rn1RMdcis+VyWVt3A3udhKy4tdwcTE1cHs35tyPFRucQDd1jP/GMl32H0s7t
uI6ogwMD9P43mUyfS2fp9Dl4ES9PeSn9lt9UG1XqeAE+jRlG8TWjMEd8vmxEq5LSaUFEs/RP/pB1
Kjlg7Nd+0ue4oSpGneXYgmrui9C9nbf1lGSNDLK3or7IBz+qyhnx5gDQUpdGDBFRyqMkgyZe3El2
IBrGCEAUYeBzqzs3bS2PypREnbV7bKct4S/t4tmhiw+nEx/tuGtuRdlGSyb+MOWZFEgLU1sU1enx
j8XV9+sAj6lxCSDNwFTNkZJet2e0krYhRW4SE2mmpbB/GNKpktgWQdHFZTJpZbJjnsLhD0s3GPau
tgAyo+Zpv1TFkzhbAk78ZDqOZEgNfGA1FdwDut2Zfm33OyJD+EDW2zGlzSYIP5f71XYgoXPfvh9U
62GMgDiQCMwPSfWPEwTlLFiv2K1lyMzfHwHPPTP69jm2TlxH2rln8yRHoM1sbBZ9GqUAkIiPbsD9
Nb5K2gwsKyHcx69SblJInABBhP3DyhsUSHtN40nBA67rfufrj6Eqhbk/eOy2Al6ARdtk4ykLnMRE
TqTXQzbRXh/575CAPPmf7Qba71cqjk1B/po0v3Z+BskovGrgcvPaTK/c+5i6B5tDHLa8TCMzBlIz
6H5mY/NllQaGDXOqZX8KKTjYyO7E/cpaeR6D3YD8QW+xKNEfFlLFE3I3Cvey38tXJr3mT5eDXUgt
ZqxeDdLvudHXKC7oXGq3cieezi3/DqVFF3RgjR6S9DcBPAGcrELqthvNluQYXrghuwgIwIKruqSe
4bBPUlnNn6bq1zsIKXTjm2KVmw5TNmtVovqNYX5jYedGyv57EQ93JwgFVfoUvGMgY4WYxCPlAd6H
kvlQWvPtQViE05uSFj6UZpYrrxqMYJZwp5A6iWziTFW408p9pXqpNDJNQKFfk0N/41QEtSmwzFhF
hpRkD8fC1QZqPuQfXzn1KRFK7un1gezR2EzVYRGiRXBt9kaJ7j5ZPtknxMgaTmjwZUjjRuQUm3Q7
LOXt7A57XnAOafsT2MrhuYLfZrGWBpLe9Q+cdk8TUfNf52AarA0j3AUC/YXMagor+fiMhbH5ovQL
lHh0jggacfwVzibE4o+snvRAI6rnkxENBxpCkOAAcoFGBNmalSQ+j/oWYIEmCKXGISnBw9GLKp+T
Le7whN75wt5EnS95ua1FSf4LDBR3BmSkPyb7s5IaS1Ko4lb0WRlbWqxqj4n5j4iOCW3X/gxnSvrG
Mg6l4KwdZSv/qLIH9wBYcKLieUkw4/CSnf/G+5FzhxP2+HzpERikZw0WdEM5mo2EXEkYD/6/iQ98
dETzevKagIPPDjdgeJi8rm490RRuVe0uX8YKGjKU2u/H4DTpZ1YD8+B7xHtt5SxvAsqAjZNnBDMT
7nyAlQ4sJuhOb15r0XV5frhm5b+UObyWVYitGgwxhflBwEcUr36Cq5Ej8RFO2w2/RkQ0G2mhSJU2
KlpuYzgXJ/iDqoa82ymz8c4IRclHxYSiqKz1xdH9kLpaFiGXSyuRb5aEF8LTi/Iy0qqkOZVJLjBo
uHqjCmZeQ6v7BVz0nYZi/SpArs8YRSvNuWLhGdvXDFusfaI8XR0QvyGdRv3tl/3ELz029INT95rW
XnEbDGx9PmyfyCEfSLQfDWK7mbLrjbyxqa/JViwIjD04FDBKNmr/aWn1BGdwZM/YwkOSdgqAaaCB
zlh+nc5ldWUgQvhw+jFxGC9zqDTyNKv1/0yl6volPFKjTujAlcNxCPAbrVSUU9qIgxLarfrS2QgA
SZsSM0qo7ScTw85GXl+oEeC7ExsCLtfsSEQCEcgNlt1I88nsX7vVeRH7dXo8l58jACcx9DUB0Gm9
Cdep95X5KGVP2nmrv/Qk+rnjcNQk9ixW5/ojyXptY8c36F8AMKxw+1l+dR1xIHxhSvm4cxJ6oYRI
igPoZLoGCa6m/7zAY0jRDF6cDzM8Vuxwdi5lWfwL70PheugfDNVYia0O+bSqdhSnDHFWnjf5XDqP
KwJMpzBgqW/3lPqVonim8niT/G8upBv2QyAXWlhPH/WuFr5aVI43cpyvwTP1fdC/AErKeB4JX64V
IFmBOhS/b80wJBOhzubP4oVL8azSEfBI5tSV5eWPjIhOWoY8dXsg55GlAZmDH2Pm/lVR7XTP36if
w3qCZ5AKu4lQHACHr91dWRGQjM7LLiQzSK82fAsot2I8KnfPB5BMEfZYuA92KWif/qyOZqWBV1Dw
TXa0nIxbEkFedgGX17Xe6jbuBPxgKZL9RJTuoVyVz6ZOsyqh+jsYvF8A339YV0G1mRzVciH68lC5
GHgC2N+SFBgfSjx0tJUv6HCBvcZbNShDZJgOehryT/Mdjn60b5z+pW0ieb4VhtPJF2uGWxmQaFKL
Tg2eR3RiDZ08QVgNLRHTXhXM93rvc5UaS1R3i2Ag+HXFOGeCHPd9xrGHpHBWnGSC+RO9n/y2CQ4Z
ZR90T1LvqgiO1ihgz7agF6HonIt84tMNhN2Wea3pCuA6+gQtMuUbhSh4LjQLnnXWwrs/BXsSpq+q
M58eOHzMpMr+5EFXykshNLDjVK7J+3QFEXmQ3RxHk/DyEPdUjj78Lzv/0WR9lQyxGpca9SaXLjlV
Df8qSJB9FnNjxvA+Q3t/542UD8UIwSgGz4Yj8V1MpwAfELXttvLzx3WoencAvP+/SuQ+VXEeNZH9
3uegW5uDzIuLZb7MrQuEbxXi/DB1tgVmYpMsu8Y95Z6gmv8l2T3Sy2RSsYaUBhmWm6C/IHMlsQCl
zqf42c+hRvdCZwSMOyBYHYvy4AqJReMtx0f/BsVRW+KhXG6bpp+5YRRA9mZW/fgoZQAEeN2lYWtp
vwXp4kI6WYV4rXJWIpDzozLmfYWUdsr6ed55RzkvuBkSPhrbgHNluK2/PpuMsr8xm/cgL3/It/nw
SRbSVbp5aPa3nFNplwNDUPh6YPfowy2ZQ/H5KUltzXiuat5YkNUAg2dKOA14N+jfAqfnnCd7cCTH
mmLtK5aLdKeWDw466DYkZenm0PsCU9pmyzHDocmaF1t2utKcIY1K2UnUGIyhETD0veFlWHUYuHNJ
mlLlQm4flR6QlYuCXip31EbZVjcSUwrOOJfR93A9Oobc69jWy9bHZSOkK8hHzCQh2CYMme7yKO8Y
g6wukrZRmXinOy1wfw/VNWDGrL3E7L7unDf13+k9vapF4QqU7R4ETxohpurW05ch99GJyGpVKpNi
L1klQ32D/BLeg+ywMK7r9BK6OtLou5gRkNmezEFXJJVWd0sLbm8gtmk+1YluTSzKCVba0ak1tTkW
y5L2hk7wWhQi0JsOcoVd7ptHewV5mXRcpQ8M1g3lWPs8UnrSGjh8lE3LwnlYz9j72at3H1VxZw1d
BgoBQs9vSg+91gdmSulxSny0E+o8UeS8Osnf96gCYnS0I5qdBuHawYraKLOLeNUtLbR3sA8aF9Ot
dVUBmhccK4OzyULzIktKNF7mUq9e8VCHO8RsgbWBpuUSTRUed8xJr66jNfGhK4xKXwgbrrF9J/r6
iUARRPXfLEZSXMWYixS4Ska6aQzx0vnpg9bbcbKFa9QNLIOri6jdDSIU2oBvV83C49pBheNqNNAm
xFwdljOFOxpbexphbZ1+mMAIa1n/NYZ7VzFytNdvoWbNdyi0cgPbVJC+Wl4WPhXZJxiEwDGSwpUz
jEMzZZHYeWVsOjV8y0Ic9S3+6QOOkVkbWhJ/p77VdydzBv7XYnC7H9ooBG3KOtiXzieZXtKEXLou
FMXHgkaW48a0SlRiuCE+Uzldod4JsOOyRVFvEOuoT6PBKvhoyqOw+814UUsO6Z/fAT0uceI7J2hk
tQ2gJcTH8GYObv9LOJ4C6oyCURs9UXePn2fZ77nVXzmNr2pc2Fb/T7cGrTpRv0ijEdNLlqAJdKWG
r56VKTp/Z1y9VAF+uxGYPMpnpqyid3RYt5OZs/cr0C7tVZyI5Tnz22HQK4d1PRiKHkyRF16zpS+V
MCWLgv/8bQ+OQ7TeU3T1l5JTkbT349wxAkWUW+qjPux5bX2iq9TW4LuZ4LPghw/c2MMut75kSed3
zdiVDGfbBHfqWxbBL8kyV/6u4OsTDCZoYdtopgvNR17m8gLvT4qy1GGtJRtQhtOyQfajckwELMw0
OtHkIgkvsmgPY+qM227ccU8wzxnqjrGHiZwAEbc/oEZ+jsrD2svkZbPro6NmGNCY0MPAYwPgkYHj
4KlGiFDil+rEpKPp6iGTVvkFjcCewru0VDGwDJ5Gyf1JAi19ZTtm5QhgvazExwMUcNqdFaph+eN4
AO6ErF3NZ0Mb2zRzaLcRL3g4OcTdhmXQjE6zoPjj3ppT0ch6ZnanOMMQF0FmkS6ieAKCRUel9ylf
lbpp3FQvHcDKCpC4Jh+mYPi2IRgE2tiQjTrhXU8WKQmbu7Zx0G/9hhOipZaH8Oapj0ML+qYY+o43
YoOrddutg/xLovEzEQ0TxiAUcNsi5ir1MTAFklMiy2BIk1Hg4oHBqh8cDH8qIXPPRYdQWqWCm8KQ
unkeqD6UhczhYw6GwCyPDPJJ+vSz6/uGtExX7rS4fB1pk0oRSNy7xy2NVoxuKmzwgSIAQBPXUlWA
BfnkPliKCRXxDnlhp7NnSSMwKDGhXsG93BVryVGjyPmrK19H8Vy9qstaDMZ3EglYE6+iFykhHR++
ZUyuaHF1mQmPXfO83DvjThOVjqySega4G3v4ZeCMzec/ZQygIQuCppu96I3lf16nhBM+SXQwCo86
4xP+4zPe2zhHaBD0kvktWebKi5nuy+sGNi2fSHjJyMVJAYsm1XXdNSrvv5zIqwMbdLZuUksuU9cK
rcQxNOJ9UOrMPjFMlLd31sUjZcamVMdjrfb0LC9zOqxUZmFTO/bGVWMgkzJ6kRjqFaPxrW+NwK2K
dlStWnd0Blq5Y0cBDOEYkbmSTCBMvrXs7099EycL38nk61AQeuUOAE7ao43KOpZ7NSrPp6mvqgrM
DlmDSXnpmIZXBpfPseWlAAEIwcJnNNEmnmE+rb3P/VlpbN2sXVVe8ftRAM4wn0+bkB6PmjT9VisJ
5f0vHnBPgVygDw8TpNDT/2XD7qbIF5AVoYjdyzZZm94DU6Dv87vTbKEBt9+n3L5mPFYQtBV23L5B
dsLfN7/UIpgR/ujwRVx1xCz4515qmYGBG0Fr0owZSVGBmQFS9vnLgBfbiqodmmLZfK9eOrFY8Pi6
u6+yMVr4iv018xqGfCDB3pb+7mEm45bXGLD2VE8cu2LdSCSPNgk+/UE0gcrWqfbla8GQmWv29dQr
eH3/Wz6+paOqkPkfFAWtS1K7dJ2lI5+QhPSwKuHP2GzcqCzmxHphXs6HQxkD8AUsrN6mcbkEvI6a
3KB1a6mUVUeQ/JiGnGSGJu8I/YGFsE+PLvgdjJDKrS/K7CP34tVk3uhx70AVCvUzVRJOJD+09Orh
2RmD+gv2WgVdXlPfNp4s2KD39HkbM5zUdImPd/kBtdPcMMVmrfzwT49tx9ZASZwEZ2zKFvE4MJi6
+8bLZ88AI8iYmbsNFXrrr5ph/RVF4ZBhbVVqV7pUAesTfWPcNluzVZ6Mm972ClN5004cgdIHnzb1
pkrrvPY52MEj6HithJc1IHD6FN6nJInhTpmlDtiZZVbZY4esUkViFWKeZOvHDTvjWIgOpYHIEdUv
jl1p+PdQXCMLm54X0e38pJ/BYnhXXMAUbJGL+r/N3KiSniD0Pdl/4NLXqcwOxlur26rBnjpmRG82
CdX2tkBNXJC7JAebNxIc8D7RAof7c9MVtUSEhlQCGyYi6/WulKoWxGGiHzKdgwOLtDVQY2/JdiGK
tsSpE4Aru4pCyitpzMVUanwgQ/CxjoQEATB3n9EArRCWAX5+hSq86jIvnC8/I5jXyuo0okTN5g82
4gjq/qythqy19rkeGqLSUj1V53PKeO5NHSMoknFMU/vaChRAnL4xmNbz9wlPwvCJAcOVoFUF+yA6
gd63lYyQu154vj5vGbpDXDzH1dei+DmPcOH3RjjVl3dMpl0YKoMy9kIfel+CEcqZiCrBl3yZoBGP
eV6Ap0/mLaGd5IZgRX6Map18TveBRycFiNHUyCYei62Z6jAH1eW6kK8S2g60oouYKVyXH9DJpUpB
Nf9HxIfUO9NTiYEyhn82Qz5ftsX+H8UrLF9bXof30i+Q7eReYQs5W7khYAiTW+/jhB9MGDOr6LoA
EOwLQwUbb9B1/CUQ5PRc9dnsysWPR6jND3cDfqhRrS3jqTbSLRdulky+RTEGoSnpCg9wK+02rVLS
SPyQqFsiJJtmk0QZytPLdGtpb/F+SiSpE+HNAkg5+r9XezFi9f2FhbBVDUdEcOZMBjNinOqaxBpu
IGDSA/9JeVzTUZx8LTY8pPUXn9ersPE8yh3/3941oltckK+ssN3G8bQC58nEER/fnWWfvUpG4N2X
FzkmfxeCzEEAdaKfApRebzI0JD6ygSWw/la6wwU+RdzwQOF8RPsvCwQC0ACDOEel7RZyNYCLMbby
oxK14LF8Zb3SdEDofBrB2SGQb3H9rAVTqJosZtjLWNhrdAwgMKNXDwFPBQABNM0s1BAMLXO9Ker+
srMaT99EhCdJ7fWHWNbO47vZBHwv3Z0vLbkBOebyw3CzXXRyHydP9Hgv/ND2ZqE2wVhWVKiZHRay
hWil+cMlMS1P885PHAQWvwilVWEiJvuw1D0r/V958/eNx28n82fmRSVOwUh+DfUj4VSWfwO+tbUI
MPpapgbPQLYlrUITJXaRtaB9hUL62YwqBnVbEbbN8ZWuwaQ56i+LNfXbmHyUv1P2gF1L4AZLOroN
zbRB0BCIJ29Qy6+nYcl+jUEo/qBqGRMaC/aJsn2PgbWDqlkwOR/8t+niNANuDWc0zpEnuJIQHxNT
kBsiVBuiiEzEd3RUaGynui1z+DYExz3wl4FPxCaUdMBERdWQf5W1ebx2xLeN7cf4MWlteTg34V+7
lqbQmZpnWHow5qeLuBVN/93kQSzwrtYZQpQZcoRKUY7gY8PKsEg8VjNNYS1VTjRl3A8kVsOZutLY
IJOhG9wLqvcaDgCzEHF+2htUOzZJ4jsE1nE5QZ55UsfLtdo+TtXd/ts8T3fRYJa/1mnXvxej6CRg
S4sJqgBdIpeSPpyMmPUDgMPcusnVYdEMXaZ0strnI4C4gOUXkEwL3oYYbIE6MpxGsZJeZGiUDiSL
QIclzx9o4+NUORwvLI/+NiV1H3yC9v7sx4/Gsttoor6BbQmf8USD6TtHlLvp+jJcNYnftMJfY2hp
zOz6tuydYQNBF9obIGhm1dUqVcAOz5kMQhcJSiEf1wx8HWHEPeDBt26NskGYVUyP5cVdBXX6hxlx
9gSylswAtKjOhXr4Rf6+k/IdjvBMtRp4EMtXZPKn71uM9yEtRBssyBH3Cl2KKu/LqiPxyopaEjOD
AOC3GeNF1CoT8wsm2eywYHbKDxbhShXStCQOBfWv8mwWvKnK7XhpH3gBmGvgWpSDpVgH13m5o1vq
Ll7eUkZ2gGib56ejkR6aOw7Evy0yHGfjvR9CmfJgNtV3JvBfAzoXGjn/aOCFOkDtbAeUVB7cwQnQ
pL33BVNk8mZEuASz1LtYt7cycAjnVqG74V/4tv2LHDVGBuEXQzmpgKEnHPBZgLL9k4w68TGbOQJK
Ol1I/RcUW0lrrYgZzbMMeuTNasXztHtMLPkpotY0ZP7BIBzaa9DNBKugPnrtDJlI6nWDvzuVkO+G
G//DvQNWGIDwBUseWaMHB7JHNzl156CRcjRbNJSoD7x7UTnwg0sz5ELbOPwO7mcKiwokBCSPHB/b
UN1KboxYyI5TNU22IIcF6ILiWZHhPcByQe27obFOfeyLcZ+/RRdvIf9IIpcSqVtxYD0/1pFvLQ2x
9yjwTB4eQxZSqH9IJ5YmNnGZYcscZV6wH5f5nFhEMWfBYSYdlc8JfDeYDNvafSPM2q8ZSXmo+GAd
2eedn0XiF+5kUPxR6W+HadHzz6srNlCSZobQEnaJ7YpLVfjAg8OkByVIAss34lGSyOlsKCceBFmC
Jj6E5dIcRiA7Q1OhYQx4YT92KvQZmN7iOdY3PkCk2vwcPzmNaTxtgNvjRKgbIL6ZbclG+/j1QA6y
afp+ELQWbSmk4jDLjFVXgclJ6iHbVzpxmusc/OWa0sDDS61ImXfHpAyuUCi0vp22X7GMZSZEzdiZ
W9SYedrpo+dY+lufwaiOcGNs/k6ainqO+nZITS+C/cXaXmbluakxhd2YLi1icPmbCO/oEj88oNTk
/oLTN+Y+zYFltRG6Z47LMzVNO76oY+dm1l+6fDJL36vXrmvwQzvVO2DiKh7z6c0Sftg1XBft+wxY
P1FSj95HgHz9F7XHKAaG+P+xgOjSxV+cFkd9cDP3c7Fh3q6NgPD4nA2lKN+igiZGWdgk2rrr3vMj
NNfCuXblulCmH2ocgwt9eiR1W3Nf2QoW9CRcu5DTC9Xe5g9/aSvGWxcmmX3NKgzLyShNPMdNolS4
VLgJiXFNGJ8qUNOkNFXp0vvfIg5Ol031Zx0pJPXKwI+IApq7r+6J0SNMXo45uzBFcP8h14WW8LGQ
C+tEbWDReEO2CK8A+x/FxSsGbPgXb6y0/szShDa8o33ERQNtLb440msIGMeGNwR0HiqcnyPkPiGg
Q7WCg5WX3Mg6pVXXUZE2qiPA0njXPfMEJqebFP2wQ/zgE8dgtYKXb+l+VWpYHboReK1Bh8T6bh+U
ovhUZslX+Dgwf5cgqXS2XGFn7AnsOTQVZINYOdcvxoM6o/fRFfkwJ3p6kmVrMMCE4j2VMeG+OR0u
dSyHasSPl+unp3ohd6x1ESxm5fg2Lmx16TLzGJaOOjOUq3mrx8dKVTSZMlPV7gGtv+AgBCM29hj5
KV1zZWZcFmNy1xZfzVABPGsAJLqVNeRiaNALoRAIz2Jhal0N31zADAKRBSzmnaKcvFBuTDolDlZv
gvqYuI4tb9HSb8nDmTFjvlOHPQok3xu9VbD1AQTUdPdJRsZszlWRF/3h7JwMSkMlPniFbqw4eKL9
Uu7oC/kv0JFeSAPes6Et/tAFf+F+TGsToWstFo5mI0GjeyMvqxsVqOUJok53Gye7BsEpdmsmIP6x
XRNa0OaU1K6JkuLS9keVLSToEl0kcMOVJNrfHlO31cXaYWZ83M4Zi/40IeTUIbrTGg2jsPIiP7HS
rWB8K9BeqRXIM2BTXy8qYSC3vXsdGNBuvsxpJ9T+ixJO7Ofn5EnLtDxs7Imhs5O83QLsZQ4tjrAN
61/N+O+weB/rcR1u4dahiaxN9wJnH8dJrZM/z/9QAXZccjmpZFkiEL9rDaPdfHfLRyQaNPD67xI1
v1s1ZQv2cSjdDPVbufwAO0NEU0A6GM4GGiIEy3huXMokxz/dw1DeQRP5JJYVnO6s1YfD+68EESYH
iGU/Oiw4KX8RrPCN6Ue9IgU0F62uxsrW/+TkH1/mNvDDlalJQnhfGBFl8qdIvywwYovl47xh8JKT
10E/lKIKZ7t6DuMGPk6iY601zx8ksnOWhj0s7bcSzKRE1S2lkN7+1rpAWzk+RkAQANaLtHpMDgW3
ZpViMnQVGQRx/iN8U6JhANraRfngLfIeyVZGhT/lMc2oqG64VfvLluxqvT/sLNh4L+/nNc/6jJLm
aLeN032vtbuPSehtkmhwxhv9oorTzKBwlkD8cwisRracV8nTI57hnT61Xf5Hi+qbrCS/nCnQxMgn
Go2LnVDIVQ2Y4+0FdxEMF4+BJP1la14MfQWa66Xu9W0gOaiFuyRTdeNxndXr73J2LDLQjC/9KF1d
n9cN6alV0CS/daGfhzhzVeYIWLHfmZyKppPwfcMn8bT2mX+gJdxB2KgEy8xoiwq7xJPGjnn8NLhl
FUdnLcgyBnVJwc9cNXuA8g9lSBhb0ahd00jzUfeHkHdUupQ/olmZaIJZXtkL2weCZCWEK+SYruPy
lcKkh6cEUEa5oVmwk5nx5WLgbBX2jXRVhyicJZvwXF+JMpAVA8Nyk7btc+wbu8hZyNcFqKzTN8FH
o/+0QDVjQ1FKL+wNEoBfeLieetFQecYRxYlmis+9H+zsRhSuTLO+uYgGTi9qiGFJtrvSZtao7cyc
ulES3/R8Jl3DmLMQem9pjD7a3yWQtxhm7Y5mKBdc1XLDNDUKVMqoG5YajAgo3h9A0IZGlHJ2PCdV
q590KjVj4hVIcQPPeMucBTNa39HdYNibexIJ/3CtEROkwagkqzHU7mJHcL72n2EXbocKGGwyTeUr
xIZ34i48W4y/eTw2ARDN4SqVqTFr0w6RXqrpr/wVRju60045Cv1JEe+xmtwJ9ooudVAxgADbpg+O
rxISKM2l6cR63wfgv4YnjapSuQO1Pa4o6atKrfr3uaSLzQi+7qgEQEFE2ejKS0eZi1zCWFKvxT/v
iN9+zzlY5vpoc4ByKicBmeTCLGh55ASdkdMjjIUHtxfQKkna78rfDTnHVIQRu5dSqd4jNWbZEOFA
U1qwG/K6vrVkBqZieeEOT9Ovj873kY1PEOgwq7ebQ+VGxUvz4ubSFAeHX48M8Uip/527oDHboytl
cQZeHTIOvAYSOnYSRiCO4yRMRE/ob0fRg4tH1MSXzvI5wJznKky9QkEaj7FGZDAGf/PIWwfzqe7S
6LumpGZ+P+Skdba4wqyIdnznHHHHOFkBzhz2omWqIIxp0901QDlxfUr7ISbzDTmo7b0Nc/bSZM/F
oroItss/S3FYdGPJByh9qc4v40CnqODp7oIj3SAtFCou2qRsi/zlXyql0LE73QSMBOEPVgiWUUOR
SJm3CeD81+R47uSNG2/YuizoC6QuVUeeV4i0MjiCEGwggg+zEthzgYZUtad0UaOYrH66w0miTgO6
2nMS4bsHxQIBIUFRdmMqYCx1XxTFIe7yM707CsGIxIdCn6pCV4Kco0gha3jBA4qvYaRQxTLVSJ5v
aSS104q4TQSppObVi3vYT/h4BrpaPknp6tgXqj4u3TID/raqthgqzvRR6uQbslFabzz1OprhUtOv
tCF2PUV3fGPd5IWoGWSrSlK6tcf+iwWwYYC3K+6vT0Mma6ICFSQ62Iy28N/+R2VJ10Zc9KMk+Cac
RglRh4VCV7pejBgT4wXUOAOyvFaTbrM5wvz3T0o3xlmhn4g3uZxZwJyT33/G6TND0otvYEdmsVL7
no0QNSxD10oMVWKIj8IoGAH1oZCJRvvCt1FMKkpnpmSQOQWaStgsFqxKPAPST9zKiqn0+4TZJMq7
/xVrIlTTEh2ovyazN5pvI0MUyQ9s09mm3r58uX3inbF/jczKFuxmcrJvkzD9pkWOXEXy+vXZdov3
YRuRUtoeaQ9g238ld6TEQtlU6L90FZqM4GaFeeWBze2MkD9iP8p3oyXTYPC2MzM3W3wWl+1W/ip8
JGxtT1iJ+Jo+4+qjeq8qtUKQF37b1FgYfJxHvylnwcRwCbr42vS+RFg5edPmn1TeP+or+zhIY1ey
YNYfdGHmSZ+341MP5ygTwjHc60LsaPF7WLpfqzY/DHcn89KUJLZP4/G01bv61QnEmVFWH81J1PSh
YENuKkJw8DEAZGVcMxEkk6E89JXellTAl24diDlPxGfmG0Nm+8hsUw/m5N9n6tP4RHF7nQdf34UG
ofutuD4aNIdlNzp5cNJsLnz0GLxQ9d0dx5x2Sc4lFhn8JxlUKOcQC6u2xzGBhLt5WYYaFUo7MKan
aGKTnePFx/rPDsBhDhVnphAw0gCJml8sjP41bvryJ8JLSSmu++uuL62o4lYhBvtTnrM+QYooeMV5
G7yj+bdrS8g56dAoUJ6B5AylHH5FwRmfcq1KCf2fa3XBrG3ret7aKZ7O6WjI82iN0g8bDmtOCjv0
BDFIhi8b2EIpumZyRxALDKyH/4y57RJd6zR7vOJG3z74zF+EBLUCELnt5GCooyTFtr8nmKupo2iL
bHStZ0N4XqP8dUqcLriduN/0CeDznTzDkV3LIm8GJDubyV9fPYKDM8LP4/NlGfSBevoxp0qvRdLu
4U4iqYygvHqSl9N4HtKTWXmknKD37Cnx4f5RBZy2TzcACh7tfuTMDOdxzMfk63lUFEg8CrnFGgQo
f+iwmRe4E+A11QN4Kfg5km/aYuYonZY4BFLhfFNdTshYoetcVLKJAFKAZQGTVY+NDVKAVNPD6064
YzcmdATtO0Y77/+rJPJxxtGLxqLi5OjLhB7YKrEyA21zAWwRu+YHZhS/9Q/QBbAAyvSz7hhwHVeO
8/6Puy0obAA5ZbrbbOhnVNx1GFWQH58n6+a36qmy+quujeX12LZeauSY4VNMEadBp0llRgz7HjEk
yoAT7nMpHooeaZIDpWe6zFmurXdQwrwnTWcOXDu9tODIayw7bQY0WyonYoAMCbwuzyNL86yCRLHG
THORuXr8MqhG+QxchrcZdnbIsYPJsfnWZtmRy44lMdKmcfos/34BX/S1jLiUMEvfgJqpr8LrSu4u
Rmhw2XNJ9Gno0Sv1IM+AtFLbMH5baEOYjYr66kSj2jwe4jsVYPQG+M1iBM/qss22lvAs+LLZATaf
LfaEGfJsh7W+PB3fGmRiZ0BxNaWb4WwGfNUcpM+8K/u02mCftMT3oK4debZsYQtqbo83TjnrBldg
aLyRSSReGXxcT2b7RT3T64JEp/6FGLpOr12j6m+M5F0YYBSjmos+LlcYw6HmZqFbAJj2Tz/L1UL7
1EUgi+MIDqY6rN5TyhGpSx9tohJbktmqQoHcdIL8ozZ8Xl+ECJNdswkXjIy1edvckfHnZJAVGTYQ
jJz6nOl+W6vBSbulg4ENn/6l0Ro08MXSeNdDPqxtTSLumPUx6z4smNsG4DKEFp8JoPxx3zucRUH6
XaHmdbzst48cuaU8+iAOcIS5NkyOexkk3NK0t++gaQALtA30wGB3VVLawwk4TGEKH1csR9vuVaih
1/j2/zISLX9cVu5Mezoq4sXqvhP6Z0YCGT/2Nx0LQsM8sbvxbwQ8ZljmNt5FDgbfAiVlMzC7k9Q0
Dmy1bqipqw+qvZunrHysB5yj0s5ZJTJ86oQ18bgEH5r88KBumd+pyjm8jtcNtu6IlE7BuKCUMWH9
ckJO9dgPTsavySx5CCbaTbVPtM/aQbanl83shvJ15BK+sE281UqvCF3ci+oNT5K0NThK+YBkVmrK
aMq1l3Gw05qduhrolpmiT8ZCr2R/8D9XPjgk8GpAHbFMO2FSFmass69XjzYpPYhaIuCts/83Hcx8
P51cGcTxhucx8Hz4J7YEh88YtmLmqAPin0TNmq2ht4NZeSfdds+fp9wT68TUk1RPHCJ0NJS07evO
upqz5CVcdudKBPnM4gHpbLzwcgAUR9r35C0gJkOkmIp0cvgO9GNDtQE1vm0oRVJhFrPzP5KkZlvy
ymo1Lg2rjPgO9vWwlWqCPEFz2dhdPnEB3dsiIJMhGHnP28PPZImP+7RX/Vp3hHLFxRM1KO0E732y
O8AH2G1odBzCoxViMTDOiSoO6G/I3lGwyOTW7w+NU9QP1ycUnGoaYa95wGnSoY5fJlvoET6kd0nW
Ktb6s0hGglzcXK9+85hNWOJ8QSYWl6kb5ILbgd12+Kfm30kPG+Tcc877J2to6uQIZ3e1RmhnvX0U
UITifTzgdvPAlFqwqF1MeJeocJ6RC/cTjMAS8MDmGed5FMeIyk9vlPT/ysGRafM30kv0uPEInoE3
m7BXDISNICL0x2PSJ1AojT6NJEtPq2wfWCrmrfTtkPkkt7djXz6VBVVQI5sDvwaQyU3IoIqdHJdb
d4EbTfe3Sz7jiJSuqFEAeW6Jx0YQSnELUcgjXYcLaUqEAAkTa1iWRBO8zPsgOg0+sSO2wOYdln18
xxvxetLIaygFDBzSNk18ZUUsNV564xbUCKJ37rk3Ra6zp1KxnEwBM7T1JLbZdea8IXXmrmtWKlHW
VQv8rV9ncvIGBlNj9URsjBF+vuler/TGe5IiOlzYrSROGRUMzHpS/SIBHQSYet/6zcI/uPvbhofq
4TS7G8tk+bB1s1f+eyxB4mwlgQuxN/x3y+sRYyD4upptnn6snllXsJ1js8PrPg9nc0Gbs2FXUYFc
gWxES5L+pU3P013xNtvHCKFaTCCy9qf1h8XX9cG/tCbR0iXMGPJ4i6kFZC5jxzzK+BDKiBf/CGck
tZP+ginj1Ho30g0/vKJ2ILU1NJ0iKaVmHLDqZtHaVcQyhQZ5G7usJ8WVfCtCv9/IDTAa69nS9ybu
P4JuH2Pfwta2Wq/7OyKTFeRJpKTWANc6npg0u4kHQfEIIY/rO7X4WVoERQ2YltI1e56dirL0pnm1
UOukb/PIbR7DiQbqj5hu10pkb2QcMz0g9ywyPY2s42mxUKsbM7aPTTd9q67gFAXnN+FqUqig8xMl
Y9liVKwjkBntlUKlenM5scpXbPIr7vHMyt+lX9ypYyVIimYDRt+IJiex6ajbgmCvq+bXuBaSKE73
d1QjG9C47j8tesLWmNywnjwAAn6fLSuCAbKXUhxF6Shk+ZPlXs1xMb7zt0S0GOv/J7uirS2I/T3i
qWh9acWCdxMGnPidbdcCZg893pt2teNIqOMN3LCVkAUemNXygxWQ+FZCHT1DoxA7P6xEAN2Irbx1
vMBXQ6E9jmdEx73Xtwv8Mk3EsBDrfFHCWfrALDoDJw5uVnwX6dVEaZRswx222tMFhSnG3V2ockmY
f/Xa4gpWI0Z7ysMtgGI0nPvbj+jkwewDpxItnRDCpXeVPovbMjTV4ndVz9dxa2H2svcChuUW///v
8G+2c6YHaQIdEGtPxzSorufMB8lXGzjOgjJX2BEiMweoYVShagvRXjIemodSUP6siG2zWSiIJ1Xc
neF09uM+VLpA5kpPseQwiebvz5AeMB+FosR2N9qV7YOdLSx5xuaR4rbwjexq4xug87oOD3kDlMW+
cz7aEgbZUgACi4gXSk6PZ2i+T2rNNx0dgacsRHtuJ1p7DMMFvDaGhG5z6ed9RlntlTWSxk4BDWT3
wD7NnaVE92ZqF/sAeITPay9KacBgtwUYnAaI/dxntDuDX0pqA7ZTDpZqTAPdSjOb7m7ChNLsEXXs
0qQOmIvhaZXrUaWOFy1kAxypHUzpFPA0wkUgpGNSkyQltTk1dTY3Lh0TOW8R1U2UP9qOKQ9zHvPO
Pe6kSFLaf/twv0FAnsLuFWHOPrW5OiRuCgCsTBZlFflA/ddUugnJa79o+xTrmrBla9wZaIoDNjTk
+0SHXgsEIEJWSQ6YB0pfBxvNUNDyfAjmoPnnhKAoRnftHx6CBp5XEtEVrYNytdPqh7rKa3EtsOOG
AEy+xIvv4iLteyob6VyrrsTsCUZBgZcj3lbWDPFP5ag5KhsBm5rmBbXqM8ZwGLHjiZYAiuc6QOV5
ep2RBXkZYRBX7OZuHlzkqtauORwKm8aVpceFq1claFkrg9okNgcgdHDVM5jIfFap/ZGeL4QOX26D
CBeap29G3XFcmlWOM0jKxEqFxbXdErZvFPj2vBwEpWOk63n9mhggaV6oBAsoWTqUUR0D3R9xt4iY
idNduRAsDmrDF1K95MT7i/vtN6KE3JmI2eg8iFshXKVoQmTNZ/zzjpltqJh58Svc9IbRyjq5rSWc
NQhyioCrk1m6CuCXyf9QZ57ljRpui6k0gxpMY+1U2tGT4uLoJhhyltUDg6/HirMgZASux0im62AV
7GaGF4+seoB27Xe6rFcaUdNZQkXakrG0YJA32wRVq27I91vbMCR/Z44Zukz5dMaEhVwpn93UROLW
AaoaA1D1if73e3SJel1d8sS7XIlivUP5Sve+AXm2lNM2nt+1MTnw0k4AP/NGVSLt8piUh9SDqj3f
buo86CIxLOCdCBSLwMeaTYOL+HuHjR2UOILtRitD+Zdz8ErlVcOgrBVMecf+ERZOJhrMSoXXaCVN
MpPAN8LWfk+oCHI+nokAr3rgb7GE6duVlJWCZuBKis3FO1EXoaNDIY9rGo+Y3qNzc5EzS8eMTeJB
x52MqOMWQIV55Kopv1/JYY8p2WBp0XD9P2TK3G/XDsAx9lOLFUDxjYUKAjAG5QgDnhidZNW5/APp
NeY3+21cV+ugviv53+CdlUzATGWTHrBaoZrq/GjP0POpU9ZrSC05p4HsToJ6bUXuGYRYwGRyorsd
DA94+HBl9YP8UGe9mAyTsdJqd2ImzfPHxGdrznq5Lxo3qJRrpODinATAvhHY3iVT/QHULAFsqkKv
IPhow2wCND9wpb0dN9UBtpVD8/hAGgvqZQafDBgRg5kxlUgaYWmNleLgb4OOg4LMJBM4rsqBXM7g
+kmZsekZpxVFaa6z/FWa9LLEToWTTF1M2WS/f7fcsK0govpDKdZ2h0C62UGfG7c1L+VFzJ5vlJwU
OVXByzqn4109ULeDb9YkY24Qr/0qefwYXN7Tr3Di6bs9dJ5l+RXzr/twRRh5PUI+VJL7lmLytDTG
YF/jnz9g7T2Pusf/sEXKR0HPq1BjTDUScrLQ9iZN0uw4NDw234pMIRmPVvrxRkNciJMNAMVwsX21
WhKSoZ/0rv42lCzjEpoXY79NHd2V/jizM/k7Mx7Rf13SyrwoarzrsA8EWvluNW/Yv4UZnr3/Lxz+
AZxc/Go3hUkBIxtgAgf6nKb/+1EucQdlcIGJONNDUvvY+C2gRakuRVtCID54WoR9gw2oG/MsZ2/H
9pQGlsGwS1eHaDN6uwFNq28PVlsEb39H4za9M3OQPTsjrmOw/XP2p9xxVX8Q0QKf3Y0K/XcwB+ww
PEGa94WAV6a1vcdFThCUolDWPYGGlYkkLUGdQ93oDAP64jrkF/nv6LfRA90y5c2kur1wbeVMTLA9
3zirHeb7xVIN2PDAyf3esW+Ra/GfWqXFyWOG25JLCBi+9LmaOTgoOT3bPloNhiX54xzv8Vhm6T1r
Iu5lmTQgWOaNgNmlTouK8Plni5csBRGcMXEDAVJDqFYWRnCWDiBRA3+7r9CX20Ny65SoQigUTdzw
7lRPwYn/c5rPs/pXFDFJcSKl7se0pXpI7ZfCSjaeFh+cBf9erIBm/YaWI3qfMU1A+2ltt8G5aL81
RLCSeD2XUbpaLBojpOXQVAn9upGwBxdhUw3F1ssJ/mSkubB2/17BE+Ln4VHOJLVf+6iAYrnwbPCs
igW9JT+eYEtkmPxbgNdHOiGsqrB9Db5zRrT8+Jdt/17YelcRc6TNDmZfjWpEROIGqelP31q9HNRr
YMtwLjk4lLrQyZ4c6YU2wZAoaCYbjdgtokk6H3SFIfkiuPQjn6Mx1PjR2BFC5Gtu24xq3zukGfNE
Fu7y+soDhTqLNplaw656fpxtGA6n8Sl5i9t8etoMCG6LOmJ7tPwizpqtcdF+SbaouN9f2brbQWgn
2VDiG8YDUKKv418R6FsNbsTn23IqBpwcclLfEEM0VpBFYvaGWi9E2k1PW5RyfKqk4Txp4H3toIYl
lCbW1K8Mk4PDy92vUrM/pqCkkj+FzpD3M3jcTzCsm9Ulr5EomgGfJAQ5sdMq8rvhs4qHzbF59G1D
xCZRQ4l+bUG6OFYfcZWeDv1iEYc8gvvOxvKvNTnw99MeZ7EVvp+om/0DjbwRfuSqI0Dmfl5bK46K
IIIfUFpmKJ75zAxfpT4gSZnQWUVrs4YJy85PidJ+UJgRyUKaFigijYw16LfnS6UV4xwdNIB6o8J7
uvpM8w8v4x8jL4M5LRV03uRu3NFQ7F7sKYL1VANAz6E7IeiV+cC/Vgw1HVhmky+homG97/1gcuCJ
KEc9W+gIGUKcizQfZjdnUwSq0wqFnHLy+gUJwYiLzI9fZgLVAccqDH5IvOe/BxdnpP/s49u+7Lgf
ydOdv/BrQveAPTxpGhVPCiHa/zAoS0oWfNHFZJ0WaQVTE4llI3DuqHiDdBq+n0RRzMj1X9u+yuD9
NB74AQdBJZ/yscEYkKunAoAuDkKFcrFBjK3h5bDMz6w5uZTtwnI4OdAclfUtriQ4LrNRqCl1C8IX
uCSbMdD8p3gh15YlAeCs+oyulLV8AQl2b47TfmmRhz5C7ggfjHDEKa4PzUWJXFqQARzuXrlp4o+R
es3COhldGY/3r91UShWsDnSzvQwaox64H1YRgeuQ7+qBf0mJKspNl0j+3OkV2UUnaQyuCWri3KSR
nKVjerjr1JSZfACi8i6o9cEUmqUOmKdsS9t8RCIHiheJjCeq+jjx2gzAgR9e44HxQD16EbddY5vz
FGFvuH2azRvnt5WrmhmbbzVnRWwo2JBu76mGhpJ0057xhZvDqlliYd4EtQQcS8MMz4nxjD7ipAS1
fj9611mNFHVKdJ1WjgcWSvxfacW4IzlejFdqT24x4TR25CiOc1EPNZ4DTTYGQCDMRDVXRFApNgqx
i8XUJi9P4aqe/a7ARBuPbeszWPJfHYxw2GDXZMja9buZnIXWpynP2tlg5T4jQGidR5tMjRLiLF7q
ExzQNxIsaz75Afa/p/D9MW/LKce9sv/mObroGlQucVCDfDmbK4QoQJ2ss+hwfb8s1IRR6SVi7ksh
Qre/ZP75mcQVS5ofCRLdYF7eSTWbi9H7AigZfSNfLVnY8dBm5NxBpb5h8c6pgQv2/0ba3lpPfWbC
3dCyXNd8vXKmFxAjA40WDDrARVlYuGfI3o+CrYzyQBIZ75gLM48zQkC094x1mN7OxrzYJxQ8TjpK
90hqjmnr5oSgtp8ZIU4eZIfmKmtthUdzVU2M4JVafYYTuaW+MgGnI+W5S/VRP0MoUI2wmxM9Rn3l
evT21Qr+ChCQEzszRGVjjgLYrrcjBb+mBy4e+tP2uIEmnMFC4lJ7eCYUueIyDlU5RCbAKpSuQA+V
4jFoT+OSEf19nxn88OQhvl82fCsuU1gPzQRUilu/+7TEZk+hKixghctZNGNQaoWEdQkXijkXl2vw
iNqH90UQiKN+qMsHfJaIJ4QweRAcmnfxc3wNZUn3yvG26tfrHHZjpxbct6tIuQOlrf/esjZTffYl
rqz1gwOIV7oN+4CE7xbvVgR0RMYUNkcwnWHC0l942YaNJiivXvMLhB1WqMCuT1tbm9Uy1DRenjFE
dJQQODZzN1FhYbpFOlLM+iknVDHMywnrrQH787YCGPq07X38K5yvriaXeNXN4Ibbgi4SmKVU7OOE
wSwvGQzvUVDc4fgQgxEWvtbevvMFcLrKVVBTKa8fEoKWMuB23qx+Tbw2fmndH32AjTZTmgNB2A3O
jT3rEHMXH8nBZxhoxaiDcb7/CmQ8nypBG1P8TKjzG/9tKoszWaikrst9pLckC6k9hjpWKa26JRm1
QW9s6QvpDMQqMzipPLmZsgGlZVTsVu+7wYc14q6bpo3kzKwGe35wJGm2a3IZjqAfM3LVFmwePVrH
zfjPDh+QP1iWm50HRPcAjNrrCDw10vKQ6Bj7Ur5YjWsOY1GITUbF2v/d1xrR4THLeTlqbC2Exz/d
yLSJvnJimSmRNrXzsefySPcpct2YhzStodskzdrCbv+6rJFJkb8YNSv8uLH362ZrOwyZSeVM6/Ok
psUDx4HjKGq4P9sLKEPqm0EJ8KjwDm6veTM+dwt/QW+/JENLZoddJECpB9tn9oUTLPvVctB7lWkb
Yz7+XRylESIh84JNSmpr5nsRigQISOBoUdZKv95QbiNIzMJI1wMYreBfvfcrIH5pwczaQFRsZJzr
3L/GeT70xc+dtFXVx5ameALHcdZ7I1ToqU6NYjuZCepL4itvrj+rECH74PFN+cnF2yBSZOIWyezj
WP3UGGgfy/RDSnD8OSp9Wlqy1APRfK0b70ipH2LpqtknM29/NX/Z6syoFwsKcY1hl38ahuNtzxhn
zgAMFmmLpsi/IzuDJVUfCcFJg7paqxA66VlEejlu9uZXvJrqtSBbu3QMM17IQqBsXYVEaK0Vy+f6
s0REO4BFW7TJWpT7KoqFxS6iHzqCgmG7s/DplRhWADk/Un3Lm2AnbdQSaFAwXJtOS53U0iTj2ROQ
Ja0rUB031Ra0L4LfA5YjjhjWKYTpmbu2OS0XsxuEZZg3AatM50sk8Ckfjuc3Ar9cfriNsz4EEZ9L
2wX9RswuFOv9WNpMw59n0KJTc36cpm0wtMMKkh7Lhqk4mNzYRVYOqWYA2TuYTE7ksP0kGO9XFcei
uvtn3kQ6+f0bUJH46rMzgk9hsgm9JzE95IOwoUHuhPF1TnJdV/3Buc5apg6zssh2K5/Ilx45ZwzK
b4HwD2UwptmEUjA3KJxRSvw2v17IabAPSuxo24e3d9n6WBgEccYyt27Ygg9pGlK5DAAdndzWIQHP
ZF6ZZT+JJRt+NJQ1qvveS822Nk+KtbNjnYcN+gYRoY2EgWrEB9nEMpeDLgBiFtl+laYhaPH4GyQG
VdcwPWWuU8YABuderCKIWKZfZg8SR2x1KSBvxBnhmqej37UmnAOGnyelTW9+7vtYq5ZFQ1GGRcmk
TtxCmNOYoMtUyRdsGyp8/DlB8aUpfnmprUV4k/OTAPrRxKAAKyBzYYw6zSdyMpk1W2tilM0xVVpM
SJdtyFvIPp5nu10CdEm3oiH1F2N+nTEGm05J/THyp60NsqbUa5bkoMq7J59xAPK6Ddk9f9Gw3Rtm
V+pLaiRVCVecCMbmiQK4M8VkylNdVzIDI8pHhoVEY7pitt2Z9ZRitMigDVAJOD50zX17CRi6vT6x
AWf27tVamlHrYFdxPjda1Tk//BFYAtF190cl17Pn50rdvkrmIafvAK/n4QndKTU/gZI4IWADdLxP
BTg9IDFb8gdbjCYO5+pREeMv/YKMOaiEIvesZmqLAwGw/VX+U79RaIMMBTeSV3j1S+zhIR1BQm60
Y05dgJuDyTxVCF7sjk0OxNkFPcB2ngzR4PlcVSzUtnauaOu21jUTwsI2o7NsfsY1bSolwaT7ZquM
cJ+AqKlxR5iIJ2mrBqIC0yx+81rtOvIkgOZajvKSkwSraReypwFYU2D9R5qGRCpUzxIpcMyOh/5o
NLwyCmjwv4KY4IyPZhHBt0Dve1tkOFsLaVcGzWb8tcm9LYxuw/C72fQriR1/TRnjnXNYqVcqaPoK
xSzTSffDIqoK3ZQ73hARFNkIAjW62f77KLYEq6/1IhPhmmKo7DNK5DMIjdULhMPAQciXjwkcaMhQ
1p8uPDo9jFdQi9aF2CWC9dsAwoto2xx6wGRpqFsZUkMhryf9edV1nwfcgrvBMqzizdCGcf1VHuXL
poJZ/tUGlmBnZ16tNTS54BVkNIYgur/F6wGYQsO7L2tQv5hCQOLCFIi5yrxS+OiaL0eb2Iehd8eB
395ANTGhSX1qJrSmt5HXvmV0ebYjkdJ7hkGW3FFWzRFENErHCi9Yz+3bNma4+hlb3yCtD+zQJN0B
Ecgw1gnHghPfVnn1c59zea5yvPeh36e2qqRngnLPhiXLhYkD3cYYww+s+3TUT0AEvUUhB6S4D+Xi
kHfRzxaTI0QLEFV6DAkQzA9NF7ehEVQbfOHTfsZpQZN0Iah0OhqVLyXrHTtSk1/JITQR/NSRhNKb
JO6t3A6qgzglDPM9OeVqB9io24uGu7nvYOgSZnfs9atJrJ4roObO+4cK5MczcMEPed2xPdNDcEwf
BFBbe5lkiOtViK7mDSOOClmIrqgVJBEubg6adDY5tMNXJeaJTSgxGd3QHQKpQ/8nevYUfW4qc5K1
undCZqzRoNadB7FvkMMZ3b/V1KK3Ww6JfouPMHioQ5M6U8AfeYzgKV/RiRIrSyBd4poTilTuPCxz
vV2tXjgydEB5BZcYDrtVhKGBWggSXNVWhZ68vwQgixCLowFx+DTNttT4fsaA1+pFmdTAAjkLCwB8
NHWuXmvcdHH9s9+iGyBrukFy2ay+oaFzIzR39XAHf/SqUa04UJLk+nlOBqRmwFUJKwhiLTRSKA7g
p6TJn/eXpOU3HkxDMBdBjNwJbVVgzgL4pJgTXChUOUQyJHvxmPYo2gSc9gF/09VwhSZSmU4KcxN8
DunUfAezmhIckejOh+9455R30FcSD/HXJNKa1v+vbT/mrfT8iLWId9rlZFavMcvAHj1d9G9ORUAI
1ePImDASL9RQZaj8SeEVWNxlt6uMFjy6fZLxzMrTgEqwK23BEASWcOEJ+nnjstTwBGbd1WhKS3fU
0q9xbCi+xuKQaCY7NfN9BKmTwEFFO5MAaPLYGkd4aRRnGD19Ptc1WhwLIWLDbNpcIhygouUyTNmA
mZV/VLVIiNfr3fZ7fO/xolSKonB3oqPsjjB5hAuCylgaEN3rtdAJpKuL6ZRuz1aigl7flDqBLpNe
AWo5yWI98xwV80kg0am5fWGFnv5yHnzLPaROnTi3JtdDVuzKTHe+s5IP9RAJqbWebou/BYtIk9IV
hyavk8mJifM+ysQUiDsg6Zq3cr7kP9oAeilgO3TovqVrgQUxKjCjdRJJYGhlseteraHzt5qWvmmv
WU13acytLjTbL4idPMpnhYV0ORjdQ6LkaO7c8kdMMGHdYK9jIaJILmpKv2Y52z2Zz2l0vXy0Iydi
3+nIwZExl7fPQy/BsTrsrbMsWw/stB2T3K8UkkP+szxD85NOYITSQPSJpo+1XdUnB6sjORr6RCub
s62x5KZAZx5oaIQqUioGrOZDqh288IbJmyM0i8X7eUpz5ekWGVUCUEaYo8qtVyZ0iNoKJPTrxXvb
PbYkvtKGUYbRHzgMRoi2TlNTxTMswIUFJeTaZLOrmhL69FyU7eAc7b6IGiG/PdWAaeDgKgE7WZcw
n8NnKHzIkXYQ+kvyxK3aZgItCKDfAGVKTgHzMarV5ZLzn/Xq9Pgodgd8gJMqOGbzBAX9uiDCWokS
j+oPOtkKcqu5OnKxqANW8Zuh3FXH2nuhGDuZbpzK+6nApAGUc1OI9yynAZEMaO7jtLrEJUwHEuhW
xX0r12nBtF9wR38jgJIkiu2dNphcwr+jgFQGbTke4161vWRIeJFeDG0Wv0RrnOwGTXip5ZMDw5QJ
iMajN2/s1dOvFisODaCj3J+ImIW7qfZWphjZVlk6ly6IgqRtEky2XKaL0hQ8QUZeHkBqtwH5biuQ
DMbDbZhjvPbn767rK33Zg//yUpLBduUGbw9q0zdxKC0OMZaZ7p0pig6lAv5mterNJrdvN0/Zgb3q
JEH5Pk0ThmZaE4CM0Hl/5DZUix9/eP6XgyzUvMSjsdnVSQggBtbWR6xReqfSwCGc2VK3IPR3nboA
XXEIN0ZRqmYXLJvBNbESO7JGr7MymRsZb58EIc/513ohP9ZP/y33B2+zF6SkF1LFz944atGVurHf
kW1FqXr/cpeK5/ScO3gmwN3akOlkKm3vFtyRA6zgj9RJ7Bz2aVIHXEhMbjA7cDPpyjF0m28I967V
Q6NX0+w/tUlylSruFDpsXKm4m0HvHOIDuqJaDbGnBCpoTrR8QhzYDBCUEUPmAdDu2O5Zx0GYXsUK
jf0r6YG76zJ7AyNUxnEC716d7TEPvFYxeG55QIQbxtA2e3gju4qbTm3kB4NH2+5J15Wh9uoqmonA
qfqd5873qdMn/zi8kqxrEp+5gM2ipRWVdlGSB5mHBzSQyxrXwBP3flEvS/nt1SCaPsNrq+8LTLdc
/yZIE4HvzeLZUETYhVNxpQ5sktlZIfCiKzQHffADoqG320mUPkgoW2wxBWigQ3TfwKpeExzfWvej
FkZ0ESkNHk6/lYfJ4/hpuLohTQ0b5luigArq1DLOWq0bX4UFvzWyrsXIhbkPoiw9eqCdaDUxYBkM
9lMBGQIiqVdRj8vLDFM2RMipLiM1Rvn8HECf5Be5pVBewFXIVEduFwiNf3VQFTTP5+2qFccHg03G
7Qc29kI+6XeiuNZPLJ3lLlgJa7PQ9Drksg6E6JERhnCVAZ85C+Ve0WF53jhjCCuqwgArTPPfp/CB
wnGgycaAfcsyS4hyQfqKd7lrBu67GQmeuFm0v5QIG2Xbid7jnQjd5FOgAY9/qbs01zs3BG0hchGC
bNsWJoufNaleyojiIMZpmdfza0p2qCn+tx9rP74OEzeGeqSaAkJxUQ/CZnSnuPo32B1HQR97z3yZ
1QplAaUw25EaHxy7yKWkQmU1QxZ2F8uluoy8Q0vYGRDZ5MoWplGqrqsIUmYq1jNKI7tjNBiYfnRE
hhFjF+H+Evuo3y/gMdKzGXZ0kKU/89+JIIuUg8BDmai+eMKZhKeF4GxL/lX0+I7FYqSPVToIGg1T
q8WRhL0Hzk3TFL8Fz91SJB210JMoC0MsaAK2E9QlHocGuNEUxz+2xVo3vpWsJkxjgD/03Ge2ofRr
Qd9hFCZ9UVXmBcktz8FXqwKYhyJbsJqOzXeWNSZm5hTCsi+Gz2ni7pRodUUtmXwFhu0cUFBtUX0w
WHebJbZe/jpweZf8+M6+RHfC1FsK9IPkNzhwL2P7fl7coI0LmI4dwIVduOX+1ndq2kxxY5RxTJT5
0yY57WvbnsMrZbeE0PZCiT+7ixCCc/n8nNCkCoQi8lylSSyrk1DE0JHIGtsF5jf0HHbwxtMdMo8m
ujJJuTOW1LpLPPStSGn+ENQrmmEhsNtUtigfGg2rum7rbbSutT0oYECO4T/jxYoWOfS0QTMIuy+R
dW6r4ltg/XN5C6VuWo/2iA1ttiDqFlJ0pyhWOUVe5uTybsH/m9CDZkxwl1VptB/uY2scpTGnfrcw
3JIsLNqVjFxDr8Bjh/oHovolpZIUuRvZU7Hpkbyor83WWIDnRreN3+0B7fx3r+A1UjL7CfmHb77W
gJTU+8YV0r6bqL+g+9eAc2sRGm+UCaryUw76snHIB3CcQl0KQC+5ZE86zLheUl2CZbJkRvMOjKs/
4b0zpcXpROEEwOLPDVaLkYmVUzUQCgUb32sUPiFwRbzXjKnxrBuJzk3rPM4Rom4iDpuyq10HS6Ip
ToVcU/XseXufhAFjevSmV0jpuBWK+4DzVk6Lfk1n84GH5Bo0h4J+Byodv3pllfx3NRlRhb4GniTS
DBo+i7AnTqkUIdQokoGqom5zxgHCgIMMiEqAKtEDn2zMT/6NB+xyhxrT8yV8b4CawLw6btYZUg3P
hD4YsIODEd/i/snkG0nsun3rGnc9me35oScqxJ4yZxiPKM5QBnYJKQoXYAgwHH47LNGKVsrcHMrk
053erWNOGoiIeK+yvXwH3BOje8kSz42Bh50qwPcYP2B4uEWN/M/ENa4XcmSraczm6XhjLr1Omh7X
af/OvJyHDbPQkX1CAlOfysQX+jCO8ptdpDlClkRP6wdGkwHv4tI0IOtwn17skfiXEdh3nKsouia+
aF1nw6EiyqhFhSNiHXklj3beZfIcbJ9lhSjqyWTIW4NzrmXV4d5zzh58240yI6mVgmYNXWOp7ZQi
0VEJDc7MsDpKxd9QQgpyx54LdMy4OptwjBYZpxhQYQIpxTx81FjuA91HgWsA5rgxAXB7d6LH6uk6
Oh3U40DDvhX5dk3HL/HnfG77b4rQPsrrCY7FIsu42gvYVbvXHw3/j2ACQ4uvZK8jg9d3f0+c/1HP
m+26re5TuYf7wrAfL91Q05TTkgLEci4NgeciYqKDLR5+A1ldCDRn8kL62oDp3e62qbYHTactlOW8
uJ3v2kk75T5KKhiouTd60FQ7N7vB9KwJ0ILui5k3qPa6aDLJWj8/mt0J8qFapX9vE4dKnCKkmMNM
Sk0Q+4STAmh3/e5ZU7gEE7w/BX/lmW7DsW7qsED0TMILt49ndBZmY79c4xwVgIuBHZbqO8aNoHTX
vKeQLZ7GU0Y97tf1M2XyKouXMk+wbjBqRRGKP0zMlkAMUgF3r0QOqDvzHXiMMEa+NDwPEukUEyUH
TtI45YJvaWAL/tvHcLETb92ryEHP06cxzhSqa58f3bRTDnBK+y6StNnux0kAw/Wn8YgQsbYsDPc2
usRCb0O0+L3Rn+o3UWQ6jJqY6Z/oRO4fAwnwmqbDvrcECNOsdc67ZqHPmR96e15uciKM/i7QM4XK
mftU3dYmzNzlXzOuAfyIC9WxfTt3vsbI8hkHSavEc5jba16+YUGMa1gSuis6Z/j5mMtBGcp5Hre3
4mPzzCdtp/LlftJAWvBWt1Ft3zy1/iYmAdnYXY/5mkAur4yFkR/rvlpzeHtcR+ASNTlnaemdP/5v
ZjLR8JtDpcITrKkqhOsN2Z2Mldj3H834NGyhGvtIFmAzic12gua42fcLOf8SnEWQ+iVGK45jGoB0
Fr1ZPqiwHizBXqMm5c091XkthLwsaBgXzhOD8pyO4kKUsQwdcdKXOy7HIIkUKFnOxE34fRa3ZIHm
qeY/7gC9zeqL4KX4Hg+v0VVqbF1gGp3Vtgib27iyihUePGbzl7GOcg+NJW6hWKlpurdVkRUatns1
+IfhezMEMhrpcp+IdfgReEkWaBsQh5raf0DA5Usc/x5N7L1xqtxBAG4zQ4U18QdpQKZUrk3d7jsw
NlwQZmecUvBk8XMqspxOyPcS0ajanxDnlFlJK5DAAq0WD52+weU5RPcT9eFY+54pfQekOtrvFlc6
0lLxd21tHHqOalUEkWkcCcMgG9sE+Q7RANEab1O7ylqIHQKjpkctUFXCm4os+8cvpJjaW0fwPwtt
H0P73VJlaJniwVJLjX4SLYeIYr9O6LTXrBwdBu2TeYIMvwpfjOgS6sdWIFwLr9342zwE4coIX19s
UA29UY80FS8DpfmbxqSolPzY391joSxNFt+VxqRmzJq8IiHaXch9MgDDiZ0OnyJJtSCF4PjRg0tO
Irl49OP7pQ11pgK3moGDDunLThAzdLYdFN0o7Xl/QZSp7HoKLtjtQXxTz6AtuXwQ4m4T6jSpuxvI
D9gkqqa+rE/SuIcSc9foUdaZpN3ywV8d822Hye5KbwQPlKwb35mDrpUs5t+4hRkJCKm1u45ufsoF
j2Rd/MnlDqc9xE1H83T/AYtAO8Zy12gVtWIawS7u1bmUeqpSnWbkPsgzhBhb18lYyok6ubNrb/24
OdlcTdbkthVaXToIoD37Gcpo9AqhXuD0x6A1bngXyTpWDBTYIcO01swLQLJTsSJv/IrQWvYN7FRU
G/qmBgTn0MF3rKSBKJUa9dInlhjU8cmiSRkKZ6MKUS+w318ck67OxAFbZpl1+ggq0VEjTjbXPY6h
lx3LO2qLFfhFq7z7mQ2g/O/a21ZLOeh0Ws3knkPtClomDIdmnUWBMcCLqhvQOcsiwFZba1gbNc8t
T4e2671ntlGt5rRr+kc99etPd/0+KTeqJs8ApD4a+OJ1o1eIRVUazv5nCj4drV8hTeJ1Co/L9H/K
XwY0saYXPZFVbYvPIhFMlwZCBG3Z33yTAYhHALBStw2MeLOpvIfEIc554tkalP8vyJa8aPnOuEZe
N3/q5ZjAhqjfpiYWhHKgPq+yX6McX9SYoL7+TyNHR86kdpQlSv4aD8WinGoatEM0UiN6rBdc7zV6
4F3XWU9JSZnarwZzt4VyCuH29kxflXlnzpSmU/gcjbl1i6Z2f7r317Qzra0bqtpKE+AeiCyjBzUi
8oJG7ItOZeLdGgvDYr+nD654U/z1izP3PzeY4jeRMjGOy4BShDx0sn5la8nUnZCZcU6Y3acxxlKg
nZAMQz+p90jXLnVcuARUdeaEHQSu7VV6vbqNbYkcxZ4HDdBcqJY30Gx+m9tmk6BHMO/t58l66ex1
pCWRIZkQTJS83bSSDSQP176N+D8C3Zim1uRABSiyw2YC8GjMW63ssfDIlwp/XmIWs2f6vzSX/4hW
zi1aZ/X0HSIxQPOQkuubm8vQuW9rThMgPcaLsh7hLJ/zAWT/R4oFRLSFgZ4+FcDH4H/50yBp6I/+
66/jfFxemZ5bpsG11qXstfCKNV56I74lOOiYtVkZ7YR4oPaReTyoYWeXj9kq75jgHy7WcFy/81Cq
WNnnjbjnkainrxduxyhEdvUDUsdT/lie07zUzlL7bpFgyaiUZrE0Ki/tUKObN3C+/+df9bBNB7ib
hDs2wyynWxN9AuXoyldh78ufCbo1/0e8oqPsIf22KblyCQ0rLofYxlCku489tJ3mDF3JR8NZhkLZ
+oYh2NJk9FPOliOiTFJ+DL7vEIKfP0uZ6cBh15pii9QU9zRYTyaeYM3NS6NgUE5dlH2xeuoLU5yr
VAb+EVH1fMrnUlW89SmhCFubpSumBpSLGUykAa4GywCEIWfL64KGybDZUxTsWt/BafW/6lK/iQkG
jSXNcrPIxYPi9/PC4WvajriHcvnoKrdE2iGgR9wh1G7uRJmwmfaFiMiIHjHwZOGf77WDjgdkSXGP
gQ0V6V9kv5kYtJoUxNi2rH8o7Ti8Dll88eNAiVhJE4NRi/P0h7AWzPZkNHXdlpdrzV83UvMuty46
CijRwmOFv+qS+hhuV5aDINtBdJdGLLU6+Oss5UIRuqVUc2+jhowEHUtokTPzz8EugtYo8hC+wQrk
dw5Rx+n6KRaoqcVP1qGrGRpoZs20Bhe6w+mOLly4UWo77JvFsOlXGeUuY3h7R3v12eHmSLiV9skL
K0mTtPfD/dYg6INiNQSnbhtVi+932loNJSgtCqd8Ch8mZHaD+TxKheNRYerg8MW+SOr2HSILdBwc
dVU8iBQY3EpfA0kD0mxJJuUqMLLuR11/E7w7dpfDsS3gnw9RS3918/lnGn3FKAic1VT5XKCmmn8Q
gyDSn94GcjPgcb40Jh0tRyY4RMSweXi6G/cMRYzGJXvBoWqraJLf8KT21rs3NN4WsthurPTmOn5J
W5E/5qdmpGa0/AZ0lK+3GZiQx5ccbcGFVd9Qqcqj3mjQpOXiqMgMBNJzcvzsZLVDvWpCiD83IKGf
XKfl2pPObAaFT9ByqxXApJ1qS52qBL6WE/I37cbXdbD/bEinGfswCK6OhWvrmC5RTOHz6xp7/Yp6
X/Me58TU0eF3X14yL8mdnV7evcSqLleurOI7qmGt5N6zlziWT5sndhPYoHBWqkRAZXDi4fI7uj6v
Yu7V/OiHJwX3aRRcK/drdXxem+MJTTwN1uq8gQfIhjtLxKe0TJ8TDpSYhCxIbv/cMGkS7zvn6Pep
ZRR/YEqhA+x+D4ssSejoQ0RnPTqHcg0Kpo68UzJXlx8JugVGY2Ta3bDJWGkaVFX5bRuzUrclqtyx
Rzy85Y6CJfdIjyDwKwq+ih/8ekWh4qEcGZ2qPCqIHMH0VGhoBuVAvGBNpPNjLlGfobWCbkXS+Mz8
fEJiHXdm+P1p+/lFeqpX4AjOIJK5hPAzAgV5Re+YrLCjZF3MN7gu6jA+QsIkgDJhEjOFQPc8p6hE
ijt7GozNMIO/zSy7uV8qpy7UFhCaVq5YbkUEgPx8psPwOPARs6fB6NGUlykliPtfXz9VX1HbqJgC
yRTSHSFZTAUsmNe/w4bGeQDM2WQw/Zjo5N2+gHROC20wY65saD/DknT/ns06cxi2IzUU/pne6eY1
GCwD6Qy0fzlBBUSmI5wIXtC2O9vmeNeBzpFYoydFG30UaexP1C8GpLEKwF++fctG3MwmRp1k6lER
ZO6g1E6SmxBtZDl67TqSoXEYlN8i7uFNom+PG7znYdYiUZGwXMeSQeqqm1K3OiM2DceP2gcT5dxM
jKZSN3whnPKPb/zoBcnkrWleRxajTU40OYRWsnBsCkXSXlTaGCifEyXjCE8dQtL1qG3UjdQWjPX6
wv914BHypVV1Bwml4OcP2pAeiiY+/qMAya8PvChybJA1yI450flJAKZM4b0aLLTi4tQauWcM8Hn1
5dZYDdhEt4OqMyN6UQPKz0CKyRhBZ7pDyUTwKUnkBQkbV4y/3w0f0j6VvShK2AKc+nmoWFzk0Vrf
7VHE0rdDtm4PPz2/aj5sXY+t127jO5SFk0mkPuRSdRrXfNDuxgHbRJumjWc+afjS5+sMfn3ox1WG
+D0T3t2gNBrcFSe75YrZXopf2BDhgTu/l/71BryskbTOipGIhLW0loxDpg7UvCte9yAhq9Rf4c5w
MigOHrAXMu9ZkgikHtAuIuJRauJNWGhPbHERvufpGNFaMRvqtCLy/Hp5F/9kTQ5b2ydgfV5OfvWF
D+bEYfPEBLLWHgHi1XkGnzI3D++F9Hyc4HuN1G6KOvZGZhv/iwJbxVdtjjWnSDJvrT9OAiO9LNaA
CbkzOlbrxl/nSUqG2hGsQcz2nhxKSIIiDTRKa4+pfpa+ewA5tfA9r1tgtTlWTesJM1UASjm2k61n
PMOSLV6v/i6i71j8uy+pd6NFdo+pk2PYaLBam0eyNuikvgTM2eiM6YaZi2abNbYQsmpp/GQvaIel
m9xJiGt5w6BGYsNNvfQMKvc18b8yPHODsg33UCWFOYhjrCVWQOFHZMMww+gHlMOf/JEkbfm6Um+T
txIO+3UcEf7ovOAa9nkEPswWwJrRubQkmhjBZKl4Y6C74dqOF5B3/etyt+HEAGsNghH7ssfvw5Dv
tAkSCbdCcciKd5cvOCUL+CtZH8gFVZMWqFbbqUgZ8cCoDCfZwSrB7dVsxTgf00YfLFEiL3ZZM2qe
mlTyccJj3+FOcs1XL93+MCyze68T8lDGDm84juRf7/tA5W3KxqTaS+LJRr5OBDn1MCziqYR0f+VL
Sa4KgjA31Cx08UXM5f6gouNV63n51f7Yv8Od8OmfQKc7Rjf/tmXsWQ8HCIM5XPycbqsW5YmTCJ2o
gviFYOvVijFlV00270GV90cVBVpbql287hr+9HuHbSWvGv9jsJsx9rMuSaymIUTO1oBDer4SMqWg
n8XdMm7C4gLFX8yRdx5JP/BCMtWPFxp2udEyaFibxSrZgyxH8zOIt9t+LLoE+Tz1XxAg5p+jpK40
coOG/g2t8cvQD0/oVr8XA7Aly28O8+OQerXN6Y4vwA0AJ7WhUz21HI2mEauxi25cZkIvXp/v48Kx
VC2vEJWHRXLAakJITmcQy3tjtttRUA7hhl6Ke57zE8ghoZGgeZKDYIekAgBLyRYoQvMbsXhiOXv1
2ZPcxTN+3iDzUVxl9QfwexJmNejhFw9QlY074IYd2KCPL4iIcv2WD4zObibWABsl72oDrMGoWJua
r1s3YVXenbABk7zwVRrtf9Nkxkq/xAQMzKZt3ek6wJshMmgX/v5SGgCz35LMVyJ5QmGYTX5oPuF4
p5rckSbRBucHnohv2dM047N0e6OS52g/q0VRCyUgxgnR8FE3IlB/LLJ0yJGwIJmz3EuQ1QUzIKyB
/FTbwlDOxNDYuiU9cONsAdryNesKPVB1Ixt3mfXHRso5a4zlRGAOoW8Ib4TtTe0bWBCOKPQcbLsZ
bt8dg806tWIgK4hzNtPAs8+uop2ZMyoj1xIEzTv5uLW2WY/tIL82hOgRz94ykyYI2kY+2jGsJjMp
XZZl9RYSj9zr2bMaQ6emooRyy1LfEYzcdfPWQPJhseTIMZz18tJF1SCcaABf4h17BtZxMT0zcW20
rAMZtqC0E6GnYWzXu3G3p98aUA+jVYgtoFO3Tv/5eVoK7ugJ3R8oLxW5Xr2dh3G6TBzjUGaBF3Ow
LtWZe224eM0CDA+rnHYKlr8+LjanOeigrcJrgaC8RjjRFswqdfnCJukoGU/IbosfJskoPVEz51ee
9dulcvdd2+KJ2D3S0cchWmzzsD51zFZKDU/2mgSIFtvH+7UTJgUVPJaJjnuadl9mGCtqiUUkUW9s
iONWK4L/W92qxwFyWU7/U8QaEKpRlhcsrxolXygSpqawVR7w626Lrn2ZjfuR37NBwht0bQUKCjeW
vYHtlGyHtck/ipnqWpkhyrTON1ogXzl8gkG8vQf8GmkPC0XQANc05/e6UtuFW9jSZ4EN2PR3BMTh
/gB7pOFXcPVAHEnYRMjli+UO/JTQcSjGr/9uv/i4/QY/WXTAop6Brx0QYQb9EVQVs2qUPnGY8/8M
OErk74Wr5aEBEpqD8uqgZ4z5hJxAb1K9SFG5E6feyotZpUnVuP3hmTO+Pa9r1a/65UjeUSvN9tT3
JMRd7SkI+/RTkuhN3C+UpYIUJlboAfshwiU4gT/nPYBOGI9BZx8Yt0iO1Fdn3M2FS0dmYtyEHzZd
CfhfKMIBwa79CDHZDpem43YmsV8ZXSlJfWz+Yz5RltVcoFRtCjMJa9l9GqRagCgRTsSv+ZGfaAZ/
6BtffpynKhgdIyI+AaZQ9U2tpqbESc2PHxJejYMHwHf629JrZNplisoRvjDa3mFmCQGy4FpL2M/U
BciIInNaufG5JfnyVbtXTaEUwpJCg5L4xHY2ZefuY6R+Fpn7zhUyojiKs1DnO9v0ibbJV6fa8SPT
yEqaUuWhqgzYfReXQjfeg66rHufxrTunyqjc/3aBMh2P2k++MLdATupUE6rSfAzIZtdIn91lgr5f
XVsGX9MZIO/CXRlM8U9/fQJlOZ+jkujDAPAQ12mDEd3Mhq5dOPSbJVV9V86hsjQv1NbFTWlI4jU5
NOvC4xaLoLWgQ5AtEfYutUd/ZOa8uxyTMBb3YHFftA+nB2RB+JVVzcp7BFs34zhEu5iq/OqD/KR9
vyOQJEBSQLgSfK+mqg5Ro+MHJdTHRVpEg2IMRUn7wpeMoEonrM6T3sICUQ+WhZwj/oYhNVjW7BDB
BttEpAlmYu19pUXmpJmTRbnl20lN8plXwyauPkjFXFxT/orBdKzNQNWNH2RdJnnwZvDlf6C4tBnc
DBK7zv1vWarfrk1/Mbv8W1HDwnQcs+vVf7jCgz8Kp3fqNr/L4GzS2Mjs4MfeOWrXjuO1rT4Vl1VM
xI81tlK8j+g32qh7qVz/rSjLlJFjCyi5Q0W61IBj8KqReaG1QX/pqIa6cRRvlp59i6OYwCritx1C
DQERKKBn4dgsfqmFdprHC8HkxXsoDcH2lHEOR9A7H8gvVpVh9j33iKle8FvcMGqS1RvXInKkGCrf
q7vNQrHGAd37XmHGryoaj0hJJUxJJNi6J6tH1i0J6/LRHHW1ivQbeI0Yk2fQ6GfHq3tMOwblz5fn
d/r1EXuKm72h0Waor5jm41PD3ga+YMslLB6I3ZThtHViw7iKGSnUwUsoWGaZftVFvQ7q+dMZZM80
LiH61xDvHPoY6kIz2+FIIbtKBWEm+nQpSD4GudfAy+5fPlHHUeDX4F4Iy6pv/Ij+szrNZIkejhws
8y+vfwzTMNEdXWs8DX+xx9MmlBVRgy5Wd8zgDEY8MuV3q0DZsNWC0WfcpW4izXCYsqFLb2/V3Df4
Z7ICeFskjowYf7AOiTHxh6eGRYCkjvD0dxNlhW41PeFp/ZtPq82rRRTfOk9KR9ab5TqjsIofQTlm
0ZHZtdkJSu06Cc8nn1rjgaOWzVf0fGG26ncFC1V4xTkoW+g+qaXAxNyfaooQCMUZMKOkMX9K9Dbo
7rKohjgcSPM/7p9V/G1HSN3pOsay8fC4h4uYUyGk2n7xBcBKp2pm0w2vFvw0QfcbyXaQizR8AOl7
pNedlObcMuZJE7OZ9WOLI/q5CBe4QhD7lWFTnQVIsCwRhHgY2HICrqQWonJsO82YzZFdUoL4uWN8
x4F/OI+9UFDJEnFthSZ+MuNEKhjk7eIiPauUWm03QuCymHoqo1oIZaF8JVRrmtsUDJXfAv1t4hC4
cTcmXUowFBVGiiswT+hWtFK4STuuO2OMuYBM95aFYwe3hpYZft747MxmDkeVQBd2q5aahz0CgRAU
00gtLo2nnJqFwxjLa/yxrEpWX9FSL/UwtnViIUrwkfyYXvYbxowDRvJv5S0iXa9eYIhhNITseqbp
andjP04Oke/uh5cg6x4T8e4lr7L1sndU5+oxu4wWPoaur/0QsDvr7OUsL/eUreB3X/9T830y/25A
5QMDOA7Vhbeorjq8POrzgANQz7V80ydCP4X47OYSFo0LFEv8X+QErQIOlFfv7BNGcBksGjkQZWyd
p+MSWJvDaJ1tvFA+oeICruBBhu7sACM1w0b/msBXfo8iPu+/75wrTxScol7YlijDRA21lQRWa6hF
xQX4wtJOaMR/q3ZBT+C38O9fqMNpmQ1qAXsL9PzYc2kWh/fYleBni93k9a2ipHL+1bEiAgNzotQ6
4lahGDuK7lciXvlgN6I4ZSUqyHS6Yfdl+DXgiFLbWNFmRPVFF2ZkB1wMX/NUgsyvISCA0iX+MGmB
JYnekge39q20W6Ipd+6c+V/nhEfYORo4yLaIBXEHnU4IukpC73ZiW5hAkiVJP6IKm0Q0QiSS+WNx
eejGlkA4NwG+rZfWVxpGX6ENvhLFIIfwi2ze+VG2Y6LILQ2BQvUtm5QE+sLqpj3JQNP6jwEQTfCK
mytCqM/b8lP2jzzNBbBA8SBvK3b/VfMfGFUVVgiT0bvKeCN+slgjGe9+J1J4cLAFytl9AkXltbGX
XYC4UeyGJsVSNaTzCYGpOHLDPsAqSR1JWD5yIUzLJ2HGh5EIInLl3h7pTYXK6cDiqNxOMK/BbzLk
AR1YiZUML8bqgl8wHG347Zq1GQKKA4OVx0eDSr8Xh+UVNSxzrIrevmn9C5gre60QLO0kS8VvO+Kd
LEWdNnqoKGVqT/r/fwAh3HwEo3sBdudkLhsAC8DWQREFLH9BPxblh9NIBQ3XmBq6dUC6aD+ZKHQy
cAWDFX+/1YakEd8BBIzj+idbD3rcYx4UqTbczUblSktW5sWBk/0hYfarbDXgmst3Ebiz/pojSIZr
9O7kL7KsGkHkT5AQwBZGEF/8xl0XMHOYsrhLBAfI+TrFOeBUrv+KYfsK7pr1yIu5N3pVf1wr7f40
Rqc6te9+tSOn27SLahyLkNhzR9TTbpLI0Fl4q7IniyHTJoicXM9jenna/YE9muF4t7bD+GWClwEO
MKNfwUp/jwWvKS237W9DsgD+tncKmT3A3SYSLdjAqDt5Nu0L46nA8EGx+E1ypg7z+C7xyu4fkACQ
Ml/YyPMf7E0g2/mYgyzL9sGKVqrAZfjv6heBQXdt3RZAgRG0998B2apSfB8xKc8nzAn1tC4eQJqY
N4Icur0DGsPMwUTsGPcPSW9gpwkr/uXvHxQPcK/0ly/+NTvFQCChzZLbhTo7Z70y31VpsTDudLKz
57GvVBPYnuc/nXKR8PAIQt6MESLIAW+kzgSlNB4xs7Rccm2emosl+jON11rLD4YOIhzmzzH1hyoe
svIvS6eBGp4MyVFcXC7zFw5S0nqCKgJwp0J5aef5JSYTMXPYlTzo6mZpcD9rH3+smVJzsYvC4BEA
ZPymXq7Tqj33sJygyd3AEtlvuwVkQPhwESJd6da544i2YNvoftoaNvJdkBNey0tfzjSM/eCHa6MC
0YE0Ky4z38KV++7GARmatp0MmL1xdii2b/r0jtdaoEnGCnMC/rMGrhhdLFVqSoTVFxdOFGu7U1/V
Z5gPDnqVTjmtz23L75b93tYkka/Fph9GHps+Y9xmMY4Uxu011PuGEs6Cz5i6DljmZ6L0xEQiZJPx
C8yHlpkrl92rZ8hL5Gb56UC5Cnb5eOZCE55RvG9+GOKBmIJu1kbNaCVRoKSz2J84CHywbjBT6qnJ
U1WJdsTDMIY5WTc3A+dVl5DX8xD/bWn+TZZHXOdOkgHuOhkqh/zPL8cuq+uObspaV8Asrf4OISQP
VywspyTVzbJ9rpjD3eOZTkqqaXYmf+P0E2w8O75nHOsHSMs5VrsIrslmv/rFud8KbKAoj//ycIqe
MmNt8Hi6BtvYHhEpaUJ9/RWXWTDTjwHtficsHke2o9YAsecVYHbKwdhNhobrbcVejxBJQZDn3orl
v0fSmRzTXtiA0va1A9SAUFHqgd8bprCTJyuneAjMFd62iOmIqHRIWWBugbuMBz1PL/7zDuNWWn2p
r3C2zgWHHuLOXt9ipiuuVAYSR5YsEcXbiDAgEYOZjcFlFLB6AWUwaI9MLsDQSV6xeHNzMH7vCcqW
shh0I02qFp3nwlRMHjJuT0Tced3k66+lxpGF6Wvc6phiY+DbmM+ezc1kAYRdvhypmTa9P5BX0DiH
IQrBtpirFJr0XxHW56BdwzRPAQUj8nwh8Rt3XLAoWvGjqQFHJwqdFk55omm88Lysbss2dxiUfPHe
Zk4bqJBxKKig/qDZvYbOCaEm897qyrjMZQ48u9A3oApP+c30toqd3wpu0GBwqcfw2kAAuejqyvEr
kaDG49LDWd3CAs7D/mtUPdaD0bTCJFy45soshNIbpQIIrndFmgVlMAfbTHwNg7ycxBYaEzrJK/Sz
2fP5GTlzWbuCTjuu0ltXWSIl81sSR0j3tFkferUwoYt7GI1HZhCHh5Q7dqZY3MBDcWOTjLwB8fAk
3gBCSp2t2c6W2EFZan0DK4vh6y4Muv80ilMOEuOmvVdpuD5RYWC67dXhxSA76OWc3LqjpxXLeS8+
0EefgckBHgUZwl7rZ9HJxsR28jS9nR2Yr4vb5YO+uhFQN+Vt8G3QFKW3oMWHMI8NdAaDIygXHFHT
ewVxbFpj9hs5z+vtvr7J4gHV27g1xbpFMHhk5taK3Bjro3tsiStmtHNL02cbjae/REshN8aW07yG
aWGXYkpdU9tuS62wDvFK/RM+PFjYi5FKJuIFybL4Bm32korpPtPmgdLYtn9ssGTnZ3NwpM1mw+YI
Yuja9UDBZ1ga+J/WUwwIO6vsmQleaES0K1c9FoX5f133DBYuhQSUH2XuhP/+8YDM7tFHsljJROkS
awIQW4VMqGy+yh7DNbI40dNMZNg4MdLGDmMSoVN5iLINnxUSgO3jzUdREtVL30XfRZe38ss5ob2Y
IWGbVPiw/P8n5ZaRwGZRsahfl70wAHl3fD2jCvzd+S/47SHJlckyjJHKXMX1DW3lDgdnwIW9hmDW
ue9wCcg0thFhB5Nt4RvsuHnHCSCs+U2EbAboQ8/XSfpe+aib05mxay0S8z0rOz1kYGsukwz1Z8JW
3YbQtHFnaGLZYEROdRhYZCGI1LqiVPRsmw1WDFqAFzNGHLBzR3HRk1mdU+TgQ5Akerq09op81tGJ
naxsmep1ktuDuRjFQZZ+wn99EsFDhqKZ7yQdRsW5ugNi2ubW1gpTEYHcYwaEq2BdpkJ+0rpwUSoZ
6JGF0YS4YD8Aos0sGoWXVVVPeD+VLUrMMBVZs2jaOXLi9E15VIs/wf9iPijFQeyS7UGaXOhv17vJ
TcHPs2XAgZphnbeIBwyxd7mFEqs5Kp9mTm30FozWMocofzeZro7ZpI3L/ApRXQV1R6ckN9Us4lts
qGPio6bz9Y6R89NACUbD5w17Co1tGJ9Zj/CiplWuGYL3p5TCdbA47CAzCZNhPmQNauOvYIMxrl8N
LJTvyTfSM8GcPltsjfIfND3c++9yxAbw8i6DPYPIOiB1q4PCoeUA7iIYpcszxbAv3UU0dGI/l6A6
lmqLa0ykRtfMWwEREab+kxAC0Du4Uvx00lRuKWQSEGi7DPa3po5a6tn6FQZRTMJMQNZCgOxlkcYQ
jNC4jNVFZ3x152sYLMdJTHhcOCRBvaK76e7kYTa6M+LeQTQnxhg0dIif5bHX2yBg3Yo5jp8Hoso+
KyMyS6xouW6yjMDqm2FJxgE7FaHAY7l7PJwBEuZRmwEEWHNmbs6iLJN7IjKd9Iza6mEAV2nrNy7Y
0T8AMikg5oxWpHLO2knvKWeNpBtLLopBfB08AqaP1NZCTSTsmpuCSjuKOvu8HUB8Gh5qxUJ7g273
fH72GH1arfMIiRqXjKu8MbYDe471iuV/E+2leZZj7zXp3M0SMShfJ3b+eEUZpP6NBPbbJkcKECIK
+y23x/ag0gMYLBCGZn81gBJDM3IxpYu7h9q7Re+BfUmj5+HXtGlxZCZupgGXzKMtcbkhlgHMc2Fz
ub5aixUmmRqN6Y5CIPeZBWSZrnDsNJu6AQG9hRoJnECUwowBkmB477cwoYRUY0VarB9+cDe2k25C
Qw4b7jxMSDV/9DkNXIgK1XPY3Ggc3QlMSSz50kt6aeVUl59bdI7zYgsGnaZhqIGOxELaOTB3KUqj
uuWJvgN5XOU0CTBsgofGqpRYKSKdG548mpSrFSG4r4cmxr/jGB1/EaCva+VVcKIuGf8rS4grXBpB
9WOYeyIsrKq32bK79He9WlhIfJ6krsHT20PbSfT+IHKf+lUme7S0De4dL+/D3gLhhPZ0hNbE1orS
4t+TsqUAHTac6cWH4L+pa1pE1/je/IkxTsXw/w8q2zaZm46Mc5ZT2UnF0bM738H4JSdag6idbPXd
aT9PZbFjKwzytD0BnhZnuTWwCzfdIuSazD76d3sobPxsV6HHBt7AoAuCdnbAYh3SlHxQYCcY8RKb
kUazlsWnjYYTw8nFTCNvuwMQFl9vI+4bFAQCXfo119Py6Y8JYiEnqMaGlSlYuEETLBP0EPZ7/TXr
UGUZAq1I4HPZBAKvNK/2dO3SaPAwkVTXna7s4OWmI4FK7QllQKEZcFppR/5ISb5tyQ7btlmZDrAG
XxC28NAQHn6ug2EQARVtgnuqzZQTiyLWmPSCzbvyNtEEs+gn1aD3+hK4c5pSPmA/J+EF8Vaxs6lZ
Ppm9wxHqClF6VOIOWu4JO/SkjEedjt+R3z1gI2S4y8FsWXF/WmOq/xUggffOCdb+vFDZVjjRfnpo
NexIBjUgyFBuDmG+CSbYd+xq6sUcJNIp1Z4xOcMdWiAJEdGztR8IUHjOLHRM8d9RM9+d9wWPTpnE
K0NM09cBOTHj86Drz4GigePpJXxmS+OtzXLxKYf2TV+xeSFxk4kvFJSS5qcdyVCnnDZz7A1iCQMR
f4pfHFS86cEpeYFUf7+aWA9JSYmx6jHbc3CnvwXV3t5cMS/UivzRug1Ohy45/DV5/EI2N2aCtErb
dCIigUaXSsAUHCwjJWsv0fEcMabaHEehoOZFiIveEABq1MCJTRh76cB5uZfUPGoOD3BBy1HiRxS+
mYndpXTmlUh2cFd9XUu8W6uOIpJAhoD9raEeS5/afjYgv04CMLNCaLThAT1RstlEzOOaAYeS6t5I
btx08+vTXOv/DTyRjn0XtIpU6eZXxZ4QQYLnIl6UbQ5tkHOZ8/5DRLowP20cNbaq98Sj30/vciDB
DjXkF/KqEpKhE5YSEAdi6jU84sJp4ZcaWhX1slwYM5SZzTW3ZmhPwFNoS/HDFlqG3C6Gm1QRh0hD
2v8bkN/LP9w+EgLkqtsWDqsFiwdnjj8qyBtNQvDOU/9dKqVZKF3aVoVmsckMjHg1cjHaStJHIr/d
mmR5bx8tPdTkBEpegrkH+ps4yOWfMrgupYibD4TyPsi4bvupu6PmTGLyl5VmhFCMN5cuSizaAeiD
cBVKbtku7Muoo+RWTe7R5xOeUjSaasR3v3M8pv3ZDJHnFZ3HtjlJ2EOggVCYL6M4IJFDsgQArHlb
eIj3j3Av+OdVRQgCPdYP8uJtoxNai7Nqxkzxp20/62WJPf8AH3pE77SzSPN0+ecDSej5diqhfPBj
1IOxDcGps1UvGBDxvV6zd0e48b928ppiFuGT41BXeXhM7F56gjvzEDJC9hru40BeMwfeHnBS2YRR
o4UxnwzrFrCdbwaiu0uyG+52HnspPcVPkejMgy44i7SOvANEFnhAnTIFm0/S1K0u1s0hqtXnJH+B
5+hKMxqwNqRdksv2JiXOPOMT6YKNpjT7Q9a9mMhp5P36j3EKhCINXHPXPhuAi0axlo64MOLObiLr
kaubUEG6R9yP46eAILTq0bwNObxTZ1xPwnsk5KQrPVTSyDwTgOFH08NYWQYpFSd0it00s3pLYMIW
vT25nxQsR+n8JmbAz3mAFNpFm4iCnCbTy3hWWkjpfz+45GSCnpS14CBtYFKNhgtGr9BSsUFxo7+2
xTjUuVxVApBELHeEI15xCNUy6Z813p6GJ+WCnAJ94i6cMjFb3mTyfUihLnlLR2KgXk5ncsesQqCF
ubkEeRKHq7YTwdNrGxo6tyyTOYAd0Z79t9YmVFO6rPDIvjGI0ZR4j7TkYckR+/6kRsjkkQ8t39B7
mbPpSqCDWfmiVgIpqVncL4xIUL4JDe/X+D4cp0YQIZGPr1J6FZUtbVenCZI1aEAjZGwqNyN0XL//
hcMLTO3BJPv/GGb9WUd4x9WSwWIDSjHLHfSTDUEhQ3nUU70pKSlfsUPqMj4MVY/6OKfZzGj1PqLg
u0cQNwppyz/wEzPiNQfBF2By9kix10CEJdNVs8bRM94y8YGUBfRbo6gjBv2scLb/glZ3AKqfgpBh
bBX44MqX6vjH5Dy0c1oSUYDFqKpgURQfV+Bi0DK4r9E+g4Cn1Vn3/LvEJ9xdA2ap+mWMCu3LGEcw
AJheSjbMqKS15I9wbvlEMqw6H/XHyq7SxlOUViHT48pkzpPJMzK4W/nRiJFTYQVLyerKlU4H53CM
8bPHXWnyn981NAW2HtvfOwcBWdzY1mwuRGcqPha5YeFAyxljDSJrJJ+8NV7ObDFZqBBODJrmneUS
85sP+pHbgIpZ5t4eHJr2v1oNYPutmctlmXU0cDiIbdIGdF9d6Rsviwpcy4nfbwt6mAEdk6Zr0oWe
O6rxZ5KoDpQ0G5agvXm3+rDqJD2E4f15jLQH0IWk01VHYkBrh2+0efuBW7Nz+WROEh7jriHjz19k
FUsvjvRhpavIyRZ2V5hzTcEt2GcNtzMZs3mzNglCuonbuuFI83H1wzR3TK2TDW/SOHnwMdogxRj8
tyWpNbmqsazQnN/P3Lh7+ok7+Wfa9cemEAIoK4fS/2KcLBuoVj2/spGFBv4AN9cG/EgX8bLN+ze1
68uxkc7/CSi5lPt1Y2KxuwoTeHSDbNoMK2pnCMhBMpbnAaB+W9dZYN+D6+jrPPKBBol6llinQqrm
6sFKEHH8f7HS4ZphQUzs5+K8MV3NouE+YqRD6xy7PALxrs9pAIaUvMx+GLNbBvIY0hXvQOkre/9G
lc4DiDG0lju40s7PJP0p/PRjpFxixJ4rh4i4nQ+Yd9OItzKFfnKym4jKYuPxzbTm7yySN+OOIu4U
+KB6CdCuL98ehU/1BaekVGLCnOrlD7SHaely2IiKlDFJGBPTEz8aM2H2+VhShCLVbMUvPqvAxBSj
H1gd64RkpXs/nBhINWrVgsgeN/PISXLlo2VE2agK1OxjwwB4+Y9M1om55RiNepLqsC/JInZx7FFe
zXr/hXIh6z0prp/X30pKx07235NaJRgr3ll1CYgLJJALl/52kDHhoCX4LHCIQMqyRNsqA9JRBci+
K+Tj5xSuvOLX7jdgfi9YdqdKT4q6AciOxi4tMRSF6Y32eqhm2NvG5ggS2G0jr2I27B9kg578OoDE
ZEcXFQBkTpv858/coc5qpQ9fKGtopoKWyU3lC8ZcgCD0lBta6nDuPCS7J1vBg7gZAMq7Qb3e/eDc
YFEkr6yY/KpvDicP+yLJKJgaz5tQuOpkb52Kt0v5+w45zrVaAYSW3nrZNfoM/NWCw6xX0Q3xOjDD
F3ZFdgJhERyCN2gM5r8UiLwXvg4LwIzPKJZgh0/dIs1xej6FvG92UDlZk/QMhG2Q4USpEODB/Sz5
n9Q3Hx536EtRsjmAZKf52KAihbDN2NaCJ7mg5Lpxj/lIC9zufYt4VIUS8Mc6pHfYwsfhTGs4hiv3
n6T/J0YDaaQqNWV13sorv57U/bfd/PnHUGD6rJosdJPyCy38Da8TIFfZGbvQ+m5eoP/i4FxAuhCO
tvHvoSdGncJuFXvle04VotsgxlMGUpJ6Sri7U8/QRVE3vhULUP8X+bkxcgE0XQh1IZPoxnOOKim9
XUjYLx3ARnrxBoPQpIhFq1BG6hWiZGnp69yDCoW3DHzwDNYW4Qmf2DdZo9qArzDappstTea0H46A
1FDAjFzRd7uW5Veu1+eSOSvnlbGMj/feRRWxhUdciQd0Nc6miZzYcNBUvoWZ+Q9+Izv8MEE+DUP1
8OqKk1nzPuMamtxWs7ug04tfr8Qw2k5ieEqjEe/awcmAHIaqmuiLbos8bl0SBWj0/PZhWLIi5if4
LO7s+yU5liIGAR0yg0PQTtoLnEq61Kq4gZsIbANuRXcpgCo1nhLSjMgwSQeIDFFHjoUD7Wp2lmD3
sKxiYfZG6WhCEj9FqSpiENAoAY+Rf1TO552Xe2HySu5W+ZyxwD6ljcY+koERWeh5focIUtbCxiit
wr/HsiRuCWPokBU7KDUaZAtqWk898Cy6q74K7oXab0CeIYLMMV775e0ZQ49UOqTnysfocw5A4X15
Ji7HNIGa5TDvYAcyBe87Ru7BuuzNuB1z0vsJ1Vq/J88NFe4X23d8XmBt/AbjhcMaB7aJLuN+uP5+
qC22oYtpb02lg6qQsvKGvxYEblOL/d5gZgIqx0MdA7GHobsgVdteB0GrlEVRzFTOvZhb26ODU71O
fnW8E/6YoW6jXW8fiaypWm8tpLvoeFC0ISW97uTc1BEqJAJ8/3YnzWU2um4Qeuqe17J1eQBiN4E9
SnBRnL2KCB/leZRNMxSeR6teqIBPfrWtljahNiaakgzhymi9UJ5CJrLPZzc4NNC6Ju6CDpceXhil
bQW62jcOCKrEOq6t2jK9GXnvS55oGOrVTpFN55MPXqEGpY8nJKE9W8UtSGYWa7AfjlexsFZ3yQk+
T4dq54d+oEeOSmoxG7Ahsynnhq4P4J3zYft7/enC/bxM9HMg6lolqfU9EYm09y2B0lEXHtRHiXdh
8r2c1W0zAh6gsyooZ/K1k88pycWVZaa1PJJNg+IGjjZzgcJ1Ii6D5196+tsCV7ranZmu8qL6TqUh
kUr5uuEjZYswbWsRV1FnICf+jpqfLBZezZppQfD/2djARp1NR122NQHdvXUWX6vkQlYGRIUSs6Vg
vZ2V1CM4HfUJYrlt/8hHcKm6YxTxp5t1KDhq+9WjtO+ObG6DR53Zqb3uZZ/H8Eaonno3FPXejft4
Jr9zOH74GU1IrtTkCHMl8rzGa9PyhubOAZY0qjtuQduUfGK1UTMYdhjIsg4jX+R2e1jlkcEcA9o+
FB5kP4CShbgww0BumYKpIj7rGV4Etpf1NkVYvhlmOvsPITmdk8Qy+vvQ0HPbNlVRDDXEXcL0eSws
f2zGnou8HMSdr4ZcGIlXOXzXtEVKTDuVjLjvz3FF06KWiw7Vv63B7QhMBoieDGszcfZXpqatOe/Z
Gocnsm+t/EfKqnlV+Y+eDp7Qyozia47QtxpH/U2hGs2goZmdqTalMxY/w3hjdxI6jAVpOBblpQBp
xClVv9C/5M2hm/luvkRxdml4e6+lukbx2C6QNFm3wwVWTTlAZyv5UOtLCwcQ0iA57u5Zs8AOlPOo
2SBJrYGAYFlahers7lx5Qx3cvyp/Azmv1R5JIOMJo0J4+up8hTJpet+tXdmKJZCadKto+hFDtBBN
66UGbVUqIudbmWZC5pAN3rAu0wWwYRxZhemKf87NUGfdq78o4pyM7A3Af90S/TURr1CMqpJ8h/J1
c0Bpc886Uol2qfOB+Ht1WI9iesq/NI7M69vanslPcAWaC/wfoXKMAT6MLXmm9FmT379hqJJI3pDW
bnEBzPJz2Up2Efb8cj2ShQE3eswnq3UGR6yhpxme4L6FLNDCvLOw6TY6jSk9dJszEccCDhtFCn4h
mPelKRpLwfeH/mSVmSu8fF4gwqLN4tJmBBBr3Crf8Z36oECREuESLXhYpCHBn8gb9kFgf8dLV3Dx
q2oddxUcHOYvOl1rjtGNPL9F2B/8V+6SMYvLk8YEKAV6YsdpZAqJ4i5uGj4vcq7KzlAibwoL+lIQ
NzvNx+KOhmZVcpiAnULiDNciyzhwryZO7g7E+tqWm/PaTLKb7KV25xPjwDS5PwSxtKu4t/eJAq++
P0BC0YxqLcGCT8bLd0xvNVLg2q1Fca7sp3Z1RbCuAmZXoliiNnT9JQjOc8/o8sS9PAbxzngkDwU4
BCuU8eyrh69u//mKez/52wm0ixVri1XxGgcIA5S22mWEg6tncLwZhnemzTFWOTC+WB2D1dyK+pYq
LjN6zmyEZC3mGle5INKZnwUU8jJus9JZQL9Iu0GLfQGJsX6Z0mYpSJ8K5sdkD8VXfIZBdkv1Ip6L
1kJYX2N+YzmqXONJ629dw2vfew/8qTiLkBNFY8FeGt89dxqp14SJLYfYijFoTkjWKZRcjNdWPESW
Sua524cgodJFi5pbLHfR6056nbUk7jG3/i88hoilTz+jZOwJYbP2ZWsDbxe1vdRm+5rb+Xsko9EQ
Ab1/xwlLpx54eDplrncNXlBar2uaMycZjGTI5orbB1J1DO0rYd7ZqbpYH1cqpA+cXW91lNmfRd/L
qNrcOAQ7RTpDc8kKhY+9ApPDX2QmGG+T1VVxujL76veu8MOXb/v0u42BE7Ile0tUuAoXq1pjF7Jc
/vxwvBZ/50HrCi1SpuMu6HKwIWmOWn52kizgPtyRROdkulUSkLPfU3x7QpsEPltBSnVaO34w2SWT
kxlfiKjB96XMjmd1gJgj1bwonsKANS1bx/04L3a0WJ43ha0XT712398iDGBBkfaicn9QXQcruT6C
78Y0wrujRy+B9niPfb3wpz3xyD+fzXW2j4WeDS4ynFWb6MyCFMAL5oJ5WLSly3DOn6brZ9/hkqwV
GpbwkBm6leF8HbR4oZuli0I+vf4flMtQ8tsIK4mU+/3+D/9Yx49hisJMQmmPY7rJCQdx7cjohXbt
Ys99gFMOUFKigoHP4yexcbXgWTYym/MdCEPzldiko3lrWq1AKsxcpIbHLnFONYWQQloYXmqMdaR3
4y4HkO/kBEZYHMPxQAuf7tRtcZqmIyTvcjxYGkQVdiH09DdDS9mgYyIZi1ELP1sIq7tipvXXD4+6
/hnynnfreLWn9k93bQI9sum2d5iEGDNZKYBEmBeyoA0l5VXk0z6IZ/azE9YFPJVjpo40unMLCcVN
zGdNR+DofsXfdVLNpHBsDwVYDGVd4fIUPRs0VYGNyaUdAwnhN3JEyE6SdZrHfmUIaLWbEEu3ymbv
Ark/lydUkxV2KySZeLES6cEiVdnLV95+DOFzNHjdMJkiXLdjWlgHpl9G7RuQVnUPR7R5VoyAtvA5
yNSJQosh4JMMqCiWbpFw7lo2TBVqHbI0JLLILA02IStrw7N3fVrwuDmcbEc1up6Xg06KnrtsvDAk
ZlCezsMK0KcGlEbuK9Kbdzw8XbFuTh3QiyUyPQSs/kRTU4GRV1gfKC/+zJsPStunvOPSmqVUneXZ
XJNvRWPX6YIE9v1n2O4xkjw2IUouFnw3BP5BFJlC3Ono9D90zTr+D8SBFVB3jnb9plI1zn8Rk9kc
ixY3vJuUfbY3E1txbXmgGR37Hs26tPjYyDmsmZhODJTSOHHVX7zSC5Z1qwIHqPHt5yg/bnxczfdi
LWdfpOWB7PWHJFITguDa8LCyKHV0Dnm/b0/G5d1Bu+bMlVOnuGoEIs93G2N4mtAB4LJUnWv7Rhim
2/8p+EQwpSWUQPmxqI/I3uhgQhz3IMtsct/iIzkKU1gYiXa++fFrnIKFEhfmX1mNWUUsdFScC5j5
w9CSE7qcWkP0JRgYMAcDid5gIzE2VhC8hZY3rILIfps6jxttrJ6Rl1r3bwrjd2aBHIdBBD7FKt23
4cGPGTa0PEHsceIcb2E3PaPEtEE15mhkOiJ3AbvhfBHQd8A9fFcwrdAhtPlOxztx+EYRdiNfufzy
l3HNhFfYLGnKjMPOHjbegR+7lThjHI1d4J1Ul/oLfqSbOkMKAjdYJ4pJpnYJ2dh1BDoNGU9nzmqf
vo0oPc1LPnVV81BU+obuyT8WyS9hlret1yvaNTAFpzzu026pP7ADRKU1XABz5qmNuF/S59lyBQG4
VlCekK/0JAaPFZ4o/SQA25fhiPzMQ19HMMikEtLhtrlnj2SQk0KjjJh1c6WwF3kjTYEcucxd2c6s
0MmzlNF21SfanuVssz5IdVADSUN1EhhHEEUHwb3yeNKQ72p6z+oZBnyNyUM3P0y3hF+Xb0UGMY+I
Lhzkm9WK4YIAv3h6+zkL9FASKlIAbPiIlSVi5Ix4omhcCrTQIKS+dMvAr3u855O1UoYswDn+paQU
sc2HdQ8WTa0Ywu82kWf2vwY5T2WbNWuR2im5xUuWnctLk7NGJtDG3Vlb6W456FEH8xliqX7HbvtT
luwkK1//DDUt8ZsAaOxBAws9fiXUgQt/w4lJv6kBon5xtQ96cFmMq1MChJFQiwaxV3ROqSD8V39N
xU4xPb8gYGQmtMLVKEDGawK6ueag4Pc71GUQCWE6oGmFJgXzdaXUZxkvQQ9VYAvNqPWfwaXgL0k4
8fWaKdqxumR1pU88z6vKv5cCp3APUTS+7OPxBVTD9xYLKDr9BV7FsaTI39lbf2JgwObW6f7xxPwk
/LfCkQiT+L/jtE6SyU3+cweWBrIpHvzpOwEkGd12jLYht03UZvO+314kijoyoXLqglpp96EUSI4l
ucEoueC0m7S8+uNhcLatfymoQ6oFCD57KMH0eoYYKYWnbEI7Kub0aeVfALC6ZdARozcl1woVx9yp
FT8oRqa+xYlnoiIl8HAIciCou8Q/EyggTBrez0nZRGIzABr8T1yvThFqZCB+8f+oqvlZAbieWPpF
mtTgrem4rDnTQbAOCYCNvPsTg3T5JZBlCdBwY4t6AZPHC7QB3OdEuuTHHhkAczIEzSf/xhM+v0Nu
8S7QIZ0umKdPGrf5py+oDgoLA3/i/dccZ6h5lzJyxKj1VwyH6yGv5cwj3UT9jL5Zqj3emAVW5Pxl
2cVrlFf7XYUTtmem767OI4gpXJSbDJYdg8dUS3RhSNi++2oJUp42smE9OLe+2HBlMeni1Z3oLDTf
Xt21yGuZc61FeF4mMgqrEk3f73n9fu8Q5K2bOVZTMFWRSKQIddQyBIxwUSOuln7a0+JnYW1x6tGD
FjdRnw3jWo9qX6BnVNuDxdVrH7f8WTG6RXSnTm/7Pz3ev0MZS+pQZZ4JEEJaZ4dCn1p9MdEhKtva
lkFdP1xIu9AyjMuzcmHuBVp+CBCIFQ9VffTbKHnk3zK7Xnes2oNg73NufE248f/JAKonNj826Tz5
bvvSH7RBE3WVM1ml7WRXyoDOuyZI/jFqnVzNQgvBC/EbMhSQm2ri93ynRcm8hppCJ6QUFCQDvcXs
73rCDijb6dD3zfjrvJLs2MUCfNIRBHX/mDk5tHDUrZxcph9LxC6QnWNHvEhvLP24y+X70tKxXzhh
n+SqFPLLFxojDO3KEv+hC8E1j37NJ8kvf+MWrGS9qKac9Zxtv4p/TwaRsIv29wFt8EcnluNvQlyX
QvWac+VW4I4yQBxNhwBkntgFV1g4zReJhy1EIsM5bmp+rBZ0wUhCpru0RAEdFCG4C57uqd1kYKNc
XCTCF6y0WIeuFMYwgfbty5x1YJx7+N3nYtJwvjKeduf0CBfnk0dzyP915i9Qvl8wMBWa75fSVf0I
SM/uWCQ2Pa0II14SlEu7NADL7oYEI2y0FQL5hTpUKlxDibol92eD7jrSQDwCdBpe0TR4ug66jBO4
p3+6QauQ3lzZKPIjJ/munIMBXNwC4nnlQ7EqwiAKy3WuM81L4TWj/ekt6Kh3dP8XU5t4N6FkYTTl
JX7zxPskahQCLO14AxNIqYvAY07dcNu1AovRHyHMlTgkrhdSzGDoymFZZ3dPw+i8rfL5SqI55cyD
fdxn8rvPHyLMoQFsaddk6WO8EHF6hnE7yeJEsuQQgc998pXsklS/8V0zQddkkLT39C1PygSmRgZo
3/icKMqi3h5tjx/Ta+Q7kW/e+32RVPSXxl+WgOkd5eOvyZbxuQ+FKYfOu3xL61ApFZ8QLjgGuiRQ
eXGaO2su9GhHIqjgHe2+JT+mr9Ba3nxdPpQH16wjOQ1as7BFVHVyWjeIZxJSzmIWeXm9N0JQdW5a
gQqDqllL/6+ApTQPXX93xuZY/5OIFnnRjSq/GeoqEig6JcigWAwR4tHK8WrYvf/1w+9NDEBqAqMa
Om0Vgv3479Mgr1C+zyFQDtjsuW0Gp29Fm4Bt8lN68sc6iiIMLHJZZYBTR1PO4I6oLpdB/3xYe5DY
NRaqxz8LYT5BDdj4uzApf/NRAyHDmXyQAUAgZItPuqYbO0vpeqImtd/mt1BN6skCioS/sZJQfXkK
qSkRrOMd7KtzzqtJBEVA0d/Kbtatkt1W7D4V7Qc8uw9wayh1PAQYcbn1bLVmXa3GiImaRpXD6219
7ttPjuBgWli2yMtj63/d432vowkpS86PUWIkT27lYn3pScXjEsh7IHzVGAMMunSqBZKQvFnGd6w3
kOLlqtz4TK/VPQuf1GGa9wf8mj8ghBznlZMD2DlTPRzLr391X58jSijdzf1K4AbglcsoULsclb/b
HwCmsY82Ibq0+bNlfCpSH3G8tVyDKurCURIXzlQOB53xXLxoC7G+shLuwRPY+EZ5DGj6vPIO3D3o
QRUgD8udkMoCS+UcYSfnU7Ro16E22Cmzj525MnNgawTAVZIl9JVnIt7HoOOoL4IqH0PedU/lVbwJ
x4D0BbXjVYfwSk85Zr0dI4TAyAXJ+5aMDNICIyo31ncv7L1BCM3KQ34+ebJjmdMZlImW4zjzFORT
QgZdL5YCS/r4o1E+jaJ7Wtm8UcmnKken5wnjRGdD1CidQXnF/uHXq57dUJf0EXJIzd3Z5XYWntP8
UVhYfkgNa3fezk5Yds72gixfRVIv2AU+ESjh4ewgBP12qpQOtZ8rSMPkt+2ytguyeHbCsJkXvWvj
+gBNRnTakNK6B1xVbHvf12yMWCBKAfO2Jcf9cm6Wo+StcTKtD5I3B/czY3F12l6PY0fXZwlN6ay0
cSgn+SefJnDlGnTrCXmqor2HAgZfK4bScxLcBCV0m7s15/SGm8v46XnwaqgtcseLxF555g4bfHFP
f+VeAsqT7Aet2dS0e9/udY//FoUVOx52yS9x2CcpcZd5BHdIl9zAt+9jX6J5XgW/3eg+rcfCsLHJ
yVeYwihwT2paJnOyTO5RDv2GNjt3l9ox2In0exb4Jy2cKaYkiZnRyjyfYdOBGCumQXSAclZJmtkL
F+q4J3q+UmJ3U8jlzDiuiykUX5hVntEYiIt6UHNeRvKqnJUEW7rAMaZlwnCtZTUFcK3Xm3HKF5WW
AoVWPk+0OQ0othH/JchiMVPiudsEV700b6ER8kPe/GM8/YwgK58N09Mh3r9VLCNNXZSxsNvrxTqY
Ra4N5BQ8qZX1+vUlBfK0tJJaMJ9OP/XZTfkfuA499UIWdkg21DUekZRdHB/FLSL/5J+3WEmd+ayY
CDHkyijmcGUvXmCvqzaP9MHnHoYQyLdZg5+W+Gp1Z/FaYpbA81uzQ1qwWwdC5lt+DmcFzDXSJKy2
E1uKFQt/hCOU7FMl7mMVPVh0s1aNqZtKLjEEGWszXTqKhzpp8VXfNm32ceGr/Ur6xTeAtY+Mw/Go
gryotWhckvRIcoWzgpB5fLHbhiPnpp0/gwQtx6kHNwwfokfzzXLSLmYFHGQAet3C2OcDp2tnNFLN
nHsERCYWTfiaPP/7rbxf4uqpxT70an1mIhpDURyjBWddI5EX1Ro1iBg4lMXkuDB7reHdtdnrrbWG
ymd1dYDzOGNctCbcSRc3T6WPSL3m6JPSoHKToicxL9yISCWnvRL+JdvkKK70AEt8DzWM3YaJTqhJ
dncq+ZypiLxdvZlkDs7+QFtNYupDy0oI0R5G5VMMse9hvdoW4YvmlxgbJr7U+++2AjgVg9K46viH
3N9uvVxKKELmb0zqq7ayI3NAlW4NJ2i1y+MnswJBW9SOdcDhkKWIlue6tcoOpBlgEIvePxC5Xqxf
25Ub84iCU+aMVC8R0I4aRkpSsxjuXE5wV4i8ALHp7G1tqHst0qk8gE+4zzYum8CK9o3THuafRve7
wZHIIxY9RpRCXMLZhGkj/htngF0Bcj2cmm6b7tXwWdzt9jZ6shOpwDXbiE+NX7BEtTEqQSukFf4Q
rgPZ21uSE6+wfLJSwsxHEGK6rKwAjxS+xi6Ylb+UbMS5NCN12J5egOl6cEMIE0gIV17eV1DkGnXi
mvu9qGcRxofRSPs1bSmqpdYvNn4okhotbWTNEWsCx/wO5BvaPAtwJB/O+Ye09CaHwns7D9Imotr2
AFsUQGljVkvpYzNCZNPOITBe9qxE6mXExnmXE+0SNAMNA6IpZjAC2uMg7zgm3K9YZtiqQ8EuVizy
ixQnumUPUA4jh+praKisGWZH5iEjX8E6PkCYXkPdOC86ZMv7HErNhdeLtAfm2JjKIXoGF6d0WxZB
v6ryRxozA4flEpe7PpSkyDeVxyZwrb6scggVQyCPdzTWegFHqDJltsAZYvI0NY93bfHan8TpCgsO
5quiLDqU1qzxv0unyHWwLRoPuAA1B7ry70J/jKc7lRdlhUHUnjE+hiJSK0CKmqPIob273kVl8/iB
+JHyb23P5q0in6zeCXCzoMLp3BDX0TTfpjK+k094e6aig1Y/S1n0p1TFahSuOkMJmEyzAXhSIMUq
PsH7NhZ3P7oo9yeqoba1gVwJF03e6mNpz8uaTV4oMcKX0Dk7UBgY7KsbWV980HMNRnAmKuAdhPBp
L9SjVeMB8tf60G56JEdu47rMWZLmvPzB/a0hj9rl6NI8o8t5Vad3oP0yEdxoGpePgTl+W8opgCQO
HZeQuzvVFux/PefX+qAE7yp/7IFCWY/QZo1hw6ignTq/6iFRerjuONvBrpTlH9Yi/JnJ90mD58kZ
o2x+UpXejqRKEH7CU5OozoirLyZW+JFxOXNxsKhtHhNiKCubvCNo3yVTh75O19BD2hDG4rQXS/Ps
VZvDJHj3u7ofCOCQBqpklZEpVvqxIGelWNHYzFQCUGfe6fHviWO16TYmxv20OJp0mt3JN17bn7Vh
KsW/libjscXfUGCb59gtGJfRTKq0mJuqrq0nGoZx17l/jZx2uTWv4q9WwLuLKjkRklgIjnPChCkm
dzo/mnY9INxn9TZYSQxaw0tfhZDAqrBk8d01gzNCkEEqga2WUgqKqH665d1LTeDbXaYJ+gLgoFLr
u6SltbDmh8w3t0lnoSjiRfFu3Eqy3gB/PVCDBi6l6RHLXG7vS6XgVEz2Gw+wxmCJiQA6SclzW4lW
m8eFvOdIGey+sCwJ2OcvzNfvGCQ0QhOsoKjD+CpYF7+DuLSv5zgAD9ZABPFX/uxnEpIa32brJMbB
05tY9dFSGDBuhpM+hm3fYJk890fryf06mCIsEpKcR8XDCjda84CqbrfdB7xhupJAlfPoQbOiXNIQ
6cZHEV5lpAWt7FrpNZ6LsPRzKsefllooR/1EGjFbCf0t1NWqJVKj+fNMAC1v1I43L79rR41UrYMx
W3CM+2e1R+3ENZJVnQ7IXSLSUBRwKaQlxCYN8la+mz+a6xOf3ATtvDn1Y8UdRFyUksUL9JEK5IGG
Cy3puTKW4TJhDZnyIn9pLLfUD7fzpc/2BncWykHijaRLwAdJYQwPpSYpp3Vdt3oozy4BPRS03oU0
aqJz6HiBJn3HfO7xn4+auaVg4u32oj0u9sigxvRAOlroQ+77TX2mEVuvpsClbUCkiU1kVHMXbpZW
PxyKWLXUz8CBqbfnFilDMR+t+7JD2MyPEJFTCdN1bdAjFxi3yzFtvmxsoHDGsEEeCONwE1yw5+8K
lRki29QCOAyDgMH5xDsNJzMlBM7bTner7f6wIqTsjOoiRt5JjV1f8uAofijVuA6kqpMf7aIrlZBl
m2piOwQ/BPLZgoZp3Xl2CW+u6Wtg4ljveLTYSmDNCWcofN53rQTdKpr6QVc6Xh71rSkuW1K9SHtR
euBUxeas2ObP2R25eeFl4UFQ5OazNxbryQQzRy/G9iZT2TFJTYdjNsO6dx+X5kbSCTFKaBiaP/Zl
Gr91ugURtUfN+KQHkgvl6C/iLZOwHaEK3Qo0pOayrQlsN0A80k+NbSe5GsAIby5knbjb5M1w23WS
j7wAyqpw4mos3UVCwJXKpe9dHUOmv1X7xT4xNCFeYFyAVSoOZJCXC2a/CIi5jiJSqmHpn8BUT+Da
2mBsp+8qVl9OeOzhMvlqmcR1E70YmvAT4S81zH5pkBBqV740mnQRHwfgkdSBh696CJAFwn2Qiw5P
4yL2k5vvF4ib5nfD/pAE1g/7koYhPhiq2a8hu+MpiZkt+ExCI+xwxBwOFL3qqWKC6z3QZJA2tt6z
ZAPHr58Iwkz9AsNSH8+KCqx3c6zMlAseegG7Xee1cga5QWH+/JdCDTz/XAXqg7kZUcZ+OS0a8PrF
igHQsrEbYwVB3Hzn5vQ1+rfge8Mqsnj3FCB2EI4yvvGt0IngnyfZFH4SxYuCMFD3z2XAMocjkgYW
zOCGlyn76W0C44gv5+RuA4zRoFRH1OGRX9W1YXbgbsjB71UesU6aaj1rxpe+QFCx7IFCIEeA1kzF
V9sgSJPxPbB5bGhWiMm4tf/cbpuGYJKu2XALaiWyP4Vtfj4GY+rN4K3ELfTfbXdSw1AHuH8phlRQ
TG/cI/97JlfAlNZsXASYp6Qrv/j6/tQegTWx5i+6vbwbo3ZC/O2Jzj656/ch30Beh42FezeaP1vv
l1ASN1d/2JBJMTdXCcV6iqjNI794hvRoyuO4xrkLufLO5GCnKEUEKxrM9098tzawDnQQ2FqJnH1c
GTMk6bIJXQ7JgKd7cmQC5rrud+r5Q6Mv6cYgENVjgVdQjbj0J2H19khV4NOjA/0U7Yn/KBH34JbB
Jtzumt31NXZ8eb7QA5tdO90s0nXIXWFxNEYdANR4LSjjY0Wnxvq6kMNPbfTldBJpEDTK05HD7r4b
WD4qYia9VCFWBitfZgM+5mGk1IU486iZ7BCqS7M+Jap90xJFcpTitpWqR2JORIg7lYZBEKMH/bT0
wIF/H+a7G7WhytwSvGaJhMNTLAWAxCuAni0wtCKDvlvQhRf35pR8NIsX/9bPszzERAVYVBukcMPg
uQUzyPT1+kWw8nyjS8SLk4RKaACn5hfoRnc4EBgZj9w3b/Bv1yc1cjUgoWprSk3Kes1OVCNoqskR
VwORF0j0ywwiiB6KLZdbGY5q1g0sWZbHDlWuHtVlI9Grs5egvXr5uWldcYlt1t0p8IHL4kHKPMzC
8LVZpnGTOgijCRbkS6Ju1MFG64EnTKl7hb756+S/KondO3Kf7iLCLmLHHD8Jgh6jWiurRPP/yBYD
J5pjUCWI7FGGWc9mebjEb/1Hga+S4b0ZTi5IvAqMTmnzR5l5yThSB5mD/ll9OD1+ibDfp73fcbPH
vODF0hFYGt6G0PbED/xUP32mEzx3E/5XOxkgJaekP1gL9GP/9z90g8iD5BMRTmLIbyubZf+4VweJ
9WdyAibxcpdr7rCKYyd4zwpTKOVNPZeo/epX8wqtSkAWmaI2hMkrpxgMQWDPndvulnEY37QRno7c
ZNelGC8C/DR82dDPANphBCCqJC3xhFr9Ry+JwPQnQWJJ6RAn0TI3ovh9rKTAFVFRT7FVRXt8Q1GR
9DOlLYp1JvZBqKh53CKr1QEMdMXwASGYVWBkBm4uOhh0y/+4ZRpUoKx3IS9JdT9LNuraHAgn0DlK
ewektB/aE34P0hwqXO3KrWi1CIsP36cnN15ozPYBttm7vS3sWKqCRy4cOR9FfeSv8eWTnNR2NG8M
eKIqbqNYf78Btvbt/MePPJMdxKIw1pfDmhIkeRwZLsFyBTAFJLTDl2J/HE+1hym/1usMILSmL26s
0x8kZEf827QzeTeFbvZx5DVGI6X/VOUKL3K62vBFl+9puUE85K+pTa6sXD81EpvftpqRsmmZjg66
Qn1/NMfiggXkg5/8ap9n1jHe9p5DvKoHq9J/+LgjDU6iytz9hyDU1mfm1GE7c1zl4v4E5WjhmKSU
Fkgbp/mjLm4FoT+tsdmh2fsJbKhjvNbTLstpuNEtn6gvNL3Ku7jJ2kKo9XucWY8E5uqI5IZaDzfs
2n2cgyNox40xrYduimrfVww7LCrX1sof7h0hOjkR/7d6NCsovnyMdiVUskY9TRqnXRk5sa21j38n
p0YkGVsOS3sgvaXYO0rvbt8O+s9OBs91yPibBsa7tmKiIhKBM6VD1VdtRImAt4gnca4vvq9rLmw3
WL1e0+6SyobERpO6dLyFlGWwQ6FnR9zzcy3Q0/1VZuCueOM5wJe6SyH+W7/ioUTeP2zgGh2l1eXj
MSN99T397k5aI36A+gKccU1w4IeVWckgvneQeH1+u3lzO0z1eMJ81pgnKDFL8r6WMbJoV1tyQm4D
6x1Wh+7+eeXePff8cHTnTxHqhx4pJIx+FQ31HIGQEpiw/L10vSMwNOsI4qM+Dulani7SFneACc1l
vyaq/OoA/JU3AgXqYl0QOdsOZVR7X4GLZ2y4Zwv4JLJUDoHy97oarEJ4KQMdlGfAuo1gxUIcwryw
VxIsB1AIYLslgb7e2eo71S63VnyNSNR6bm0La0N5KCi+JNcuHgWLDNhSxTpvRxn0Uoo2GUAD+N2f
RcdSkgTBCh8hz70ZXl9rVdnkyJ5SPCLrUe6noC6xn10+MTBhtLUIvlHIR+AzIMaMB8yRmteGq2v3
PzKbXuy64d95FD2c4/JJ+o0KPZPefjdIw2NKp4nt/WQo7DgCprVabgvxV3B5uSJgzuhWfMAYZbQY
pubJvEebZG6SdpZxs/RdWaiGs9VNt5UXAnklmsqbVYu7hQytqqRQTFsy8sUE0pnY5wFa0E8w6KNP
oNmLXhYgQcmV5QU4Wwdeh0mFaB+796Ybw808sr+Gsc6KSZ3nbgawrV7o/3+xPT2v2mr5cv2DFT6C
9AGlbUHB1Jy8kW1JvVP7tAJ14qiFJ7N1rzb/r366yhzccY44nDBY9RELVyVcBAuJVMAihSHVkYYT
Ln9rYflhik2TxiTD+gExDzjcZr4k1KXkH43pdkOL02en8WW9V4VbcZ/3GbRQWojY0Y2O3aC3LVO1
gqLHQealcX2Skg4T8/EKukwXdapAqXnYUzEgSYDkh3Q0nrq93FecB9jTDpD2yYKNtYCI61ISIgCv
5X1agCOppDloEJwf9kmCuwOvABANA8xHTLJ+5X8egAa5fuEuTlwMasxq/+kkkAusMd2YRDZidAuZ
+m82RwjJjrInLZ21Be2HfOdGD0AaxaqPrgJFhkBSfDCchky6OBytBNlNxRZMpJUb/o5M5q0CWQDQ
jP9I1N2oIj9ZfSiU7qzCF2bxdbdWyj8m8tdPCQyXHzmYDzPbdRtI3jRAbv4XNOXojTFPZF79sRdP
jeHCUr38Pt8e4xJl5CmdUwv6DFyoS6rAN9IzjRmDB19trkB01IEcJ2kVoTIeVi+rhZczNfHt0cZU
SgPPaVQz4+lc5bu9S4VA6RasprwfwE26Mm/guSLqJUIdzUmjVvc9THd4xtx+9U2QyrTQX8oGI6mm
uu+kJ4DD+ebfnsFtZJUXo0BExafZmAakJa515h3vMDlPmr6xujsvZTcT34Aghsb3FrTdgmqaG291
jD2rR7gHwwhYiHLjE/9NiFoDI21+zb5EYdmUNbTmDIBezns7owfHreWyQTj7NDb9qh3m9Et5wQXM
GIGxW05DokNvFF9pYnvbnW+n0y0/bp1yzcsDjUDzygdaYjq1siLYEPUEzPn1k02PRF7qfcNLJogd
yLTLpXBBI+Ufl2dQAnme52+QHVsCQ5pK3j2SX8rK579hW5LHqZaapQOJ/7MaXdFBwEQAIKC7RszV
JVJxMCm9gWS8P0Vh4r4o5iEKhYtd89O5aChPIQbVdqFejoYIGOStdWol/NDpFfYG0AsbKXs1Bt1A
QzPZGzeK4zsa7GdvkCtNG2MXL7RM8RJf/ZjjYyq/VrwdP+sPULU5vKIWYzYSnFBeyp6R8VQh35Qj
2csqfKZ/e7cOQcHiDdPxsm74KGGBoDl+UUvv6H/kD+pMaELssaoAIWfL3PjknM6YcwNLsZGd3Tpw
IFxowODLKQBF1dyJDIjaXlGs9f/2Vi5HwYI7FBD00Xo/Fynm5pZExT6vk/3ymZ/+1oz4kzdAiY9N
CG+n2FXmzKX1zhrMB3pdjnkuh66O1iRiEcdXcmSwTo7CYNRPXkRAovMYl4cAuvVRkliVGDUIAIG+
KIbupjfixVkHQ39K+BYHnoKFMBtwpr025GBWvRvR71UUu97OQTgHuwuzVfGXyh4prCwa/g/6dlla
45znU7BYbSlxLO8JhqYmhcA/M8YlkEj2ZFCHyT46VkBBxsPrmhHSlw1lDUN0jGwKu+5bvRj3pYk6
kqA3dQ8ZUH3/zhzfVYA9ZmdEDLG7OfTUot3xFQp6qOdsUeXggrW+l4pkaTicnjYWZSvwaLHE8AdS
dgw6WR4BEClxfiDR3FDmpY3zFABU4V3b9x7YFKnAnPVGvypyJ4z+e3vSGGrN2VuohnQNaxsXchIA
aqyDV+SIouoOGElzLSqHclaqOZ1EvJr/G0aMl7JHlx0ZV1v2eQ/86ASP6DyRKdqhGKt2Dk26Jxbn
Q/F3iBVb6SkmM8uhRI5ufM0dShiuubroHmWEyYtCtWvs7XSBpjgD3H5i6FRUN4jHqXiIH7BYmcLr
Nb41yfu7JAMeBPbUl0zvNH2HZsEKYpH+8bvKE9VqHfnyNMnSf6iUzRIJo4St4pwe0CNGBqHVMpFv
Cl4qUvArLTQLKJZFkyuFIMKSBwFtn3A/9gFHRVlE68Lm6mEIaUD2+sWduZTyTDKyaUDnKCbOmJLF
bjO8B7HfqxN6GYbWYwGJjdECgqKNe1Mbt9Q/zyoH7zIdlvK3pkIFymJlXDQm9b4tCE4SaFsS3C1f
80pMNhvbBxpVu/aH76hLyU9NH0h6oHT0wWsP7qGXMtDo5rIn+PTZI9I64ZsKldYzDbd+3E0jrI9t
Yby90UXgMS2PRaen2gFPTl2lbKkMHkZo+U7Wi9/+CB57twcoeWrUqAdk6xh+XaJyIjv081umR6/f
STbYWZ3WOqGL6ILf6JYZee1E8NjiTNS7Z0IBTUFymx6AOPY9F+H8A4BKHE+8ZO1sEhUOs65zD8D4
WYOi4OZD1pU8EILPRVD2TFB/ppFPZsauxgnc5znRwva5HFiWnFVbNdZHkSE1QnCDWAt+2jNU2Lsa
mTZQC99DGxPjfv5BYb21NrRHzL+hg/YAmuyVZjbjDPkUfhUKbvPZwb56FqLtsBIrBxq1ns7E/fVu
YxPAfiQkuUGBO2vyH3FEuEKa9MgwkjTb2AmtJXRw3yHnmxvK5bOqRUJNrGKkub6vVl6UkFsasPvk
491AK/Wg5Xt3cdfJBWrGYP58/yqcJjMGAd0+iY+cpq5VWbvAeH57dC0EwdY5wNAqwbRGPg5xi8lg
2OdYqPM3pnl0STeeC9z5Y4uF1xaoN787ANauXnvi1JJPl1z+/VHm3HQin6bsJi1yCuHuIxplOV66
ECbNtCzYih36IULpd29+9JtzYKgtGHhqLSG8d2r7iwiy+UTmFCWBfHLvf5EX4DRW6bmT6i6i0X6p
OUPOHpsexA00VsM9ZASRLmsf/Nrvl1erPDGSzVdNVJoxhelX9ejOQbwSvTHIu9Abe+69HgCuKGjA
+p4jyD/V9VHjnl9LnPla32FXamaIxFbGUZ18ym+epuguo+10HYcrI8ijLkwn5EOlBvVv7xyNzfQ7
GVXxX8J1yTgFJv5ivgt5/uiRJhyCVgvV6Fzvf3EAUKlJvR+hLq4QjhS93/MHZwMSQWcX3DAu1u91
ZdISN1dWZAZX+bdzt9UEzv7ykDFhZJ+hcjh5UmnRtOGVqxhb0ppKebeUYJJjzzNlFX8CCCtcg/4e
h7OCb4i8VqEhWtfBgbz8Y10deX6mqnmsEnV/znofI1wcxDEUuaaTh/rZDZHGPZZhHO91fHEMB/oD
sQH0/a1KeSuZ36GfWyDMC/bcWjH9J0bdTzIj8WcZ6bbIa4JLQrrncPu+6vvRsy5k848I7BT+sBXe
3mYhJxmRJtveVEEdhWq4L3oe7V7GRz+sD6+fVWT9tc+VuerR0DPpe1C8Aq8AvtM6pR3NSs0wpcCw
Ee6kiJLQgyHRyYvJFmd2qL7upQ9Mxyyt/glin/rFdJiIWatkqCUkWpdbJ/Ygg5pbUot3ZyTYI5Qw
xPbLjkZrI1/Kzv/5ZuxcGoEcCdO0cRF1utSg6ww4wD+Jk1YH5Kqh8d4b4YiyG0wSoqjZUO+LTF0a
fO8rYRc4WCPKuIhc7HHWyB3j2ydym94Y/zoDbmVrAPWdgGp1pbvr6cj+mz/IlZy7VOrTwrRcbE0S
X4D1IWvfEGqjyFyPFbLK0+7fYG5nMpcj9iz5Ey5uwYyAsTIR1iU/qmpIYysRLQuV/2v/HuULpYDY
/6xWaQrz96nKvF73zdtcrqqAY6mLJ2/uxMRxHZOFIfsyYYk6V13fE6o7+fHwKcUplwKik0+u0NjA
vaQbANJVfbq9wij3RNqQ90W/WHV7IzNkU+Mk7f1nY8tCt8mnbrCjpX6HTs2YaeVqr6bSNGogS57W
kLUqdkkPbLBjblHj0xVmiknXEGj9YfDb2vWP3RRXZSsIyo10OoCVHNUBYkrPK7xi9IlnVgnwmrpE
NsPYA2vw+fphjNSoVBSMN89iyNbci8i/8bCaTy1fi9gp4vu6bJjyqXJqyKOhl+mGi23BK+jhod7F
PPpYDJsBeWmvcAWfx9Id4GZQ2D52IwbuHnc1+8LJlB2ZOy1zWPDhqHudad6U7MbjnoWJilopkj8z
bZHbqOJogaOjtAbZuJpeWkpCSdTSDDC2TAVQpFCdQ7lrPdu4MY5V5+NdEwKhUC04Z3KUIW5lan7/
4duLXztB8iFFbOrliIVvNCtWJL2iMmJPpk2WeU+V3sr4KqGf25LoMegsNvVgcasdxaNFicctV9vP
jtx5gd/vu8Kc9hHoQT6Ni9x+zk7hKyCr/G1rJdha+7wu0+uhBZcne4sFWyf+ajzl8a72xDaAVq7H
JCw+PxLQz8Ytq4ZyXSMTpf786pVK1YYNDMMhMEVsLE3WU6lM+5dAqXIxufGu/sfVdEWKeq3l/fNp
6DE5jwhRjEpqEYnVQdeHfyC32uYjWkBPmCukX8i3wFg7V/6PkRSYKZT562PBpRkJHFOsNid2J9gz
3Ys0Two0fsqJIGPxQGE3nZTmFEXkB09DeEDPh+SWxV9u0TMvabEqOUFUJydWi8tKyTo9GsW/jDTp
FOR8+2UetdSC7ytpeOqyMGqCNE3GMgRoWqO23DEhcPe/E3PxQ5MHJmpNqidz9Ogqy+po1zXr0cZN
8SVYKmzRMd1WtFOE8XxvgQdMxQxqq8oN89VgC0WXZVXh06Gl0UKnBxEIzH+dSxa0wWQIxjMLcEvm
KGOGe1uCJ/YXQuyCMP5j47gU6jBPnf0K4Jl3JzP9BgHoT0ShYqsLTHJlKQ777tWV9dZNKXMIrLJk
Ym1YgvvueHnCLQUnPKxX83iuFiM9mDuZUXSXX/HQOZ5w2AZgaLT8RIVqi9FtJK6jDgPOUZsDVzXO
fG+gRPkzRA3QagecGxWaigDAZa/u9x218pazjSIODkdAI/6/6spIfWolMK2X+7cJI3Je2p/Ry3JQ
nDARJfuz6CJ+KQYdeE9g1GJxJbf5xrvkX8/o/3A4n43zEZYE4JLX01/WmVetPVso8MCaeuFwU1Ie
M7uqsT9o19saS1ozAlmFILRkVZ8EwYDSUbMho4BlSr8XE51Y3T1Cs00afqLALIt48GT0a9lxsLQx
TQmZFmkF4OvMm+alMiPAjY0jwYjRrqlAhxt9nM8TJczevOyD4Z8+eIXcooTl0hRQqrpP+Iem4GOO
k2/kXUQUYLchAHn26BriNNb0+/mq9zc4xRITKShqI6aX77cO8i/3L+pvkXJs51x8uMUhRGaJ4AH/
+Dhr6Pjqvt0PcbAc9Hi7/aenxX0agHJd01abFz1TSX3Y2eWaUE2QEK6Axa8P8Q651LqAsMIQMpHN
vIGmbPQxwpSg/mZJDS2o9YaM/Xy7SkKNSl3GCTPySXfF3oGCjYxC/UHWK14UfLCsNtxFcf9rG4rr
EWN2S+NqHxlUDSE2d1cpeN7L/RSJmDd+YDaionVl04/32KB8kI199s06mWtrjjDdC+B7WkM6yEX6
75TNxEpsMPRKTAvh2qNQv2FIiCkE5JR+UGpA1QI/nnsHxq37iEP4zbtoB4pWdM5MG1HeisSXgbAO
xJJvY4hIHZyZ+iXJ8Y9BX4GcfkQVTyiY5xbEOsT4KwmyYlK9Ef7lSdecW0KtIMTRBQITo/Twfsjy
he6rDLVR0ac5vQ/qEl1Ofk0k2ftoanGWB+sn0Vz+VnvGkeDQ5hm//8U3EolE3f/ti3l+HNxnlFlM
4/FNnv3oavDMYmx8BnfHmj4fz2MMROJDIopIolFPxD3S5PBXQvU/XwzP9qzBMmXCwbKnFYnFWxgO
c8PV2/ESBjkN3jdw7gsrYa8Q0Fnok6+9USql4CxdQC0RkMO/OVxYdWK/i2qPHbA/chO4eEd4UmUz
DqcLhPB5icsuFNzJxJu3T9HYXepEsDMx3YNGvtJGjZ+JOj2s4jYL9BLyrKZOfnfmdsz5Zkfih4z7
U534CsP3T9FRDr1B1pwKV2nlLeSTpcVIf4S8yKlSuZDQMubtbFIx3ZNLlbZvezNCXhxhN2aiTb4H
2duHtS5CfjAa3V9ygZ/roBeV51sBZ2UnIls6NsznUZjpvLA/9TL4oyq1EuUYxYGwpOMB0v1hwelL
RYBthi+btTLlHR6uganAsSDeqR4vshGMmvY6akiEthMLY/MGaoSgmZtBuXE9Cz5fyeO1a8gMC6Up
5Ad62EjXUoKzpr10bshISW9bEkB+rQdzaYB2zX6QnSNi6Y1RsJJ5D1oSh9hbpVLM6gb3kRqPqNOH
7dXRAvQuOhXtoPuInkze0GaTzs+30jtxSAu4S+5AUTzOsB6hW93brp+XSmuyaj8ANTk6m8pojhYU
+Zurgvg6xI3V33WNfgPhxRwhhnwfhzUMwWteRqxXsiwBhTVDNxP8Fe6Q5YiGuCg5Ky2CuEiETqJU
7i+zyueMxu7GV0SVMU62aXBnyIzl/e2kRqQ+LGiu/qT5o04CfS7FSR+DYDsjZUXuKRMr0tEUy9h3
SeLvKZnvotSxV/zWJfBgAOzJmUuewJgvf6RGUEQWxPb4zQMXeadYnbwGcVvMW106DIVrDTFNmIrF
/Jn/6Y8mY4JXn72bO7/Tlb/PGDTH/2DvQUgmpO4zX7lHah7RM2NwBGRmTOuQmsFkLGU2enV59PWF
YLai0woP4P336ACfbPobjKdfKjGCCQbWKgI6TzIyYZW9mUiiSw4HPwZ3Wi6wATarwEy3T9mTIP1X
1kGh5w+I+1iIylbOUMekE5YBzMFDD6WQdq1UbuqbsIRxe0xppuz5dfzllT/d1ZKWFie43vjeizCq
it9GeBMUP9eqynITxgjZF6sBA9uXrQq62zVnPxegFd4TD4vLFpUnydCLOUBETJKxYtYeEdXPWn/q
GwUyCm548aOWEwp1p8MJJpGG1uAIqLsmU2gjrjNGR63BqWNRBz4nj2n0v+OBM0Vhvb1fSrIr4JkO
O9Izl5X4swy0TTyRBxs22OAlQakzem2/2OwCBPE9LkaIqf2ZOQm5LHoGL68s6xef/FBKffWaSIfc
iH+tGfUExdvArHSLvE9PgXE1UEni5kFFFKRcsvQFXYTwbvm0P5zEdyceejn6AQgj8mg0SS8HWjCq
TrUEMjq4R921AW9KBe1lG6kI4rbhizaWcR9q0U8IJBmrtBm2chlBOUdm1NeqXw+Quxe75KncWr5K
0eo1rIuF4P4fr1F2Z3OM3y22LJ/Otf3ZWQXh1W/zlvYYgseOhBimP2RPrCcrfL9fJQZg7iVp6N8V
PawJb6hhIo8leuPkB9MUxObG8P8/5uqHETBMoM3yoN+Ca9d+nah57uauPfVUIieD5BHYVIeTYZ4n
KrfxmTzgj5KOF8oSYof1N0Py/UU/NUhEF3wnDSd0fkLRGc/ANW/WYdU13S9Aa0B8EodXzhNJTqQ2
7uWf2OV8gIG/jATXOUpdcWUkMkaTB/i7rHGnSxEUOjkyXFgVCmA5UjKNkr1SUXu1L5rtYJvFDBSv
vuDDdTiigQdvLx7v5MNZZW7gu84Uu06K91mCPg25jr1yAD7mt5VBLDILEoSpfljTbFxDvbIsGgml
hDg3HdkLf+ITsKjEHaXeWQOvPrqeoflF9VRCIcAO4x7LFSL+0Mv055/kJLmFsk36iNWTdh1VFrw/
jeX3skdRr/Sl7p7pXA08P7bDiSHrAXjbTCaPoG8KisXemafPodtd2FoQby1GvyOHmEKYWiUgQubG
yWjVDBq8wFYwbdfLW6oNhJt0aGcAsbQRFtrGo+yo5d7+lH7LyaK6nJTbjnkOcCfTfdT+kwk77hQU
26DkPLx5m2uFd1T8rkI83ijlbpplvP9c1CPSyh44C6tXSDUaUZeO06OL18pVzrRyhP/B30/92gSZ
5f8z9WUnlvtn6PNmpsiKHyHE/aq+aPNbyLiwh3bdlrztpulPgUDp4QJlZl+J4KGhPkDvnqqglgr9
+KC6WUSFGtAA15Cz3rvYkJzk43EUskcFdJ4Lt5v+kBOjhZHCro8OOUML1EkYT4OoNmkx2TzlcpJ1
dkI1zCF55fPN8gkJGUQyVWftN6as+NPhM67Nsp2pLahwV9R/cwQuyQmOruV03mZJ4zx0YPqyNQb1
zIlIHoC8RlMr7MQLT/7Xr5uITUBWI20wKxZLuyKa/ICFxPNUpGYFMTC4Mg9YlPpupfIfTzsdT8Iu
EyYXKG/m06tWcdl9GQyS+KWfsrzKMQfIiacSauMHbhnPkMCWlBdlAf/izjyMg7LiXr58SEnFwcJ0
qT1vHFoG7I2d7DCiG+9FbwBXfSMQUVq6V7qSgihGJpjDa6edYMmUcNqnilXBEuEwqY6d8EzeARxJ
ziJkW1xi0yqCKV//isU6jBR1CFwvl2JUseagPuqyp0/MInWMbujY/57yJeDl7OJed767qi9223QJ
Q4BdD2fK03al41OZB4EAlnr0hQ1o6lrGBLoA9aSWQqWPTW1kTXhVzO5eVI6/5THFUM0iBL2JYrCv
HZu65RUddpmqCSBq1C6OMioO0+nVrrXsC5UH8Y9JErkq6rIwWSVIHMYuMSIyfTeQw+RCOOcfpApT
PQJYxlaWkMzJ3CMwZ6nz39GRsiCDx9RqYi1EAUowIELmi3Eh4AIwaO1Y2nhSBTIJoztzxBcLkahp
irpx4TlyFuv7VW0UNTjXhkX5QKwkgkkzxAEDXdU11zeTr/FQUwBPQrx/xmrSiOeQLvQ7vvYGV6mG
46FNguSRWAmJUpzw0HehlsZBto6b+YiR+zIejewZLZqcOKCGNgja5bFmzS72NejHRN6iA3L1XbyE
Xqk2cHgy7YSFP19KwMJN1SvoK8q0DGDOZW/W+2du1LpJmWJ6qg3iYoGKdclxGr1Lrv30nwGt0JxG
0A4nJ+DSAAlLVN2p0KQlzzsp9qXTwru+VBUzMkDuUpmhZXkvwDngzhIkNZypxfKxyI8dPffQq+WU
OofqbMmhmxOYcecU8fMvh7bPjqyYkmphpYnj0z+vqJsgflawsqAYdY99y/Utj7YSU1GDMf7uiZoH
YhmDIXmkyKbBOUTOY0HUnwg5Nv8SqhbVOWuy58AGe95mwHxts4hJsM5u8II5/b9MyW5EtTmO8Z2U
MRYzRC08RySMaTicL1nIHj6NOsBj2DOXnz/JjOobEfupzT3KBzaHTU1WldteE51WWceex9ayEf3O
jumuSl/f+Eau5gRB45vTBMgTHDQLX5c+sV8JsD9mf3G8Nkz/16VoV8zW695qSRjDcMGmre5pYgAs
hm/Hx7lKCgXeccijSa3SBZ/kh3L1DISOXijiq4JovKEij0p5xDdn8+yAQu3+U/UolMp5x98uizgp
dE3CrFYKDZxVEMid8UmvLQ8xPIaGH3qQ3E2DmYJJLGmh2jtiyhsNALO8lGh+ilH2lBlP7sZtu4We
pvcPzj1RFjppEzbPLUtDRn3fbVEcgOGdYpWKf70hZTemTcr1RPlI9T2Soj2rGsxA+cvjZit2W+no
Gg3bhfv9Uf7zSIxtLfJeTxw1WT+BCzK/Q08eL/P0wxvXgXQkNcuS0LUUFhZJmJhMQ1YqOPGOePs9
ZAqN9K9oAp/VWrEfg1Wr1U0qLQHyw5wMWksDIkIQEVyss6VZpABPy8VVQxtV91Hu3y4MDci7gYW/
zLsBSJtjAZ8RGVCNgYtESNILoP9fLZVXjcDQAyVUPWjhg51VPSqj1HcYCPChFsO4cyGZFFco7feG
4rLi0mmEk5/Xq772wgMuDLa0pF4A3FcXstgWjDLwC84B2YWNlGLbp8pQrqocpCiQCTDQqcut8zld
17SOzYeyOxjlNerKOXVpJPyeWkygO71VUe+cggPCSmd5PG/uHDLpdtwuoHLGQ5a/28Br2vrZNzcD
aarLyYZOPBjEv1XopTjsiwXivqWJdYXs75+bhRldjuWp8M6bAzPLDLpcmXF2jiNTIlFGvoE4ciuw
WqPh+lBqJtjjLYUREMlDzVEQLZf1AWsmFIPO9LCBfelW+YOO7q/VnQxZGwT6Y7S+zXeZjXXgbRe/
494KekrivND2+L+nOf9lHzB7Tcfq23mrkOW7X0Y3MW8UsPO2ieqiuhUNNraq2UqeDMKPFQ5kukbi
jNvMoFNYLR5EGlMLy30KfG/GmvKKa4kDM46a7w9dzBM0ijdJi8Chwajhq0FLxydXGOv7DpferUMJ
hgUZhf2mfG9EI+Ywo2yw5Ph3rzNSvqr7btY82Ls1ZNNx2qmgreb2AIgmYCBT2JUsPUr4GlS1a9T1
bMQJdT1Rn7pYrzikV73v/7CgXaTuAD39SXUkV4hhnVhPQVMdrE936HDlIO+Wcu0XALc2ivE3x32m
RXq85O5sXKuq0yM/xa9uTJoyI925b8QRBd9gzjXQQzldh7W9ArRUosGn3iz711vDRxA83Vt3GU08
hLG2OYkwhPrD5Pv+aCcLskMwqiOzKKPm7VQ0LjVEQBjs3+PVpdD80uexbNvEHGn3rMHOlRi/H2vt
LeUAgPONFArOyHmqj85tgX1Sq9yHSUO7BOdB3O3CXp0HuJ38r65XiAE/7hOOliGbHpisqdtmPd7H
vwb9fIH/WqGRaXiObCJW3hQivi4P05rNVBsz32NOVzOfFcL4R25u1HxVsS2vrMl9E7zfLQewLWRm
dCJFDf7eN6cJWe48/YgkKaBDWqEnnF/IWDl4LYQIvlBlUIoyqqFCIqDOQGiye0bTkfPKgR74WH2s
aOo8zMELTZtCahNey80hjD+GU8eokbgFzjLVTVVMm4E4AMJ9Ou4Cr4/z5Z3Ag5A7AY4Eg6Nkf88Y
dp5vifY8syK7wdFbzNJYEyPopy+0HgerNCo0t9geSXCXp/Q3Tcn6JFUWdRSXDBe8FiMljXRrwC9u
vVsVNpdzUrhI2f6fQmWbTzSVXUy1EVwjr2Iof/mF7pUiD0UUsy83/HZvJy4My7gwC3qWKYN5GPVp
fIDp15Wq1u4u2F09i4aKWfVMQlLabPfikhE+6Nlq/4fuY4ep+qicPsdpq0Q5x9paGNjNmncEv66G
32r8Ek1inC2DL16yeijkUuvnyHT6x+5QJgGrQO1/BA0LerM+NcEF+ZcY24ldZxQK9LFQTJy3AkRp
V9XCyRetvO4sM7oUstiUNhgOYDRVAqTX4bHYFyLjtW+7V9wiX0YhJJQe88jDg7P5IVFM6x1US7UY
36epQ3e0t3t4uGPQ4GV0+DIy+tLYacZJMZmIvTxkM2H02PdofdL6t9tIigr1G9t+WlUUTLRR8LjP
xAkxtbngpAtlaTfezgINwACDrDXhl+C9asA8agNi3d0EsDsuGSrQ3TKHBU12wXfqrnyBmEixi/Xl
IjqG7DCviVODiutjLMXWG2VUXN9O+KtjgELBkg80zWFNbj8rfzhoUifQFrpMrnAe6tj8JBUtlKLf
jKCS+9ZKnjsZq1/FKX/DSYoGdhE/p9fM3Cc+AI1LFkMcHEeLjCiaqPLBhZBlunJmj3QYaaxQmlu9
KrUB5h4kH0Z4rs/OwhWmKE6jJEePxabPQCcSffx2b0XKkrDtA9ewMLBSCHnx2BCwRxA0Nf/hS4fE
RIhbUsiOCuihiaY33vyN9nkroy2UdtdOzEkSkkicJIVFAKWvpBtmUr6LFeBDsOM60irG/lZrsVQp
DUGldZqiFedzNH4dI617gLlskny9p5OonvCOSS83g2WzeCp/KY6QcYIOznZL0KNiWj3Ab1/py+ce
rb+OiyGZUiwMTQtHGKnf4+07P54jJmcgrsfW07OpIhrplwZshZzXjFcyCK60cLu9CcCQAUwbrNOh
SrK+le58ZWK4zN2RvD+t70WyF1QYrvf2Bt6fAWs9hKOaMu+YesgNIiAzg73mz29A9EjN9l7hSlJv
ePkP5+QgBqEsQy6HCt2638cRD158kTZcO02nLX6mH1f/ehnrwKH10GVzrAlqCe+1iL12hJMenDEz
fco6ZbqaUhZqRd6Bb0YaKfUXDrPW8zH5MMRN03GrPPOi3BVdT4gsuhjo3wQFQomwEhJLl/Rm9c6A
Z9LpF30Xefz9oevEcXxnDT5WZGCFCeEy6uSkvFJJvFFV0hChUfTDCc1bwJn0kcT7aJ6jf00ioXhj
aWOzKwhtwhKBp1zECkC7uIvYyVXY0QG0eKf4uPmNbcGT4etz3agboS6I+viKjjojaDpxlGw9TQ/u
fDJYqTpgi/O7Yy27N8TvADbIzQf4i5OZQkFgAwUwHYma2N89XcX1viIekOJarCMtEHgFqAylHvch
KHX/dvwcyF0HU7IcFXwjUsGlQ1ChqcxGB4eoAs0RfvIu4uduL3CTBf+YBt6u8dsZv6cdr43MZxwj
lJPJphzr+K4Pv0D77RWFqwXHChh/hn4JAYzOlV0aPYZ2NE7UddVxAPiHmB8WcqywvYcfRvxfWZJa
aFLM1i9J2WDe4Mi6Ydb0VfzJg/mNARNNibcb3biIEytLHsoZBgDQn2EpX+IOY6XEDs57s7s7Akia
CKFjkLUgAkzP871hS72ywMmK/xsLREULtXhjbg2sfGu902EKfe+EToYDjYQcp8NLNn4bSrzNLmqY
Kj8CgRCC+EsABLzZhOpFzbKqbtlJBTKruDWyc4Vt8jo5XRwVi6iPpP7CCfMIvnFkPqoeWFJjH53y
9E7fhRSsBjy1OxQ3nAvdfbpmTvEOMlzJ5LrzlnNonm2VBM6XRPMV2+oANl6Cs1Gdic8snJZtGGO1
tsLi2KMMjYPdxIOi79oSBqLZopE0t990JmtMeIj6y8jbjDXSL3e7iM2tziFETOI5NtxbDzzput8p
MMhtJ9uykIu7a3RqoUdzW2b1oHKvcE8ZkYHKXnq970Vno5uug30QHAiAKZTK6/Wk0KKyoVMLeMkG
zmH+Js10V53/bbD2JDa225nTOtHqdpapdJ9d9HsQXHdRMpY082NpeiB4fFqcVuoJA/35v+bCzAro
2jdCCkAXSn3MiuFPqtCfJM+uIs+eQ8oiHt4DB9Ea6rlGZd/XEUpVVjoTTUAd8eusqnBHV+kV69qG
3kry5TDC7VVVLGG/zMsm1uwKzPmlATSpqd2URSvnxMdW7fm7hslcFgbYtrtxJMHdgXb8jZCWMY8d
ujt6DxACCw/KHZGDmytWcCXNEn4e+YChRgHdGvZcyUjZMGIoPECnCQz4TX6PFZkQY1wcWfrd4CSb
O+ZzrnthSPMAwaeJ6XEcs7tGig9QJkc92YoFtRSqQLV2p/CM0VCb0Jw+zrbJmW7YAvH+g6Wb9N4B
gdfGDBepky0Jykjhupr3NUEUkXQQ5oLdD4t8BxRwgMsvIxS5t3ZVoIp/VCVE+R5dy71n0Q5YuhKv
k4bdzbAWcGX+xmVd0ov7CATMzQXttlY9SlKl1lAmZ6H3IbWf5zegKDvZQO9vIdWYmwKItcbO0nt8
JFuGS6c7AZR3un/zEcgoLh5X27MVGEDG43FGdVOOMd1+T3Ctbny5si6hbCO+EubSxkbn1o+EOHEN
ZLbSbr3MnAZYiKOmXCdcOuEYHVZrNt8K4N2sJjNO3On8f0ADkdof/lvtXOs28ZotjBrGvRAbMbnh
RTQ4jjt/u2WwPTcf94XQFGbfWk4Thl0QygHmOw+kjydfg5HRvZGzJn441sSAAxaJaM0W4seqkuOl
q0eIZVJo9veaIR03gSHk7MuQsC7u+5AGib2TRiX6OXmEVXtkaZO3tycaCeo0Fx9n5mNOrdvMD0UL
Llb9PhT0gDRo2rYrsnCJmU6M/M/XounKyHMTcw6NcV91u9u0d2Ol0keg2+GruHGk7NIaU2+YmVej
WCtVpBnQgJ6i433Rvm0yLZLN0cGGN1I95neWNKNY+RlcHCYtu7WEqvicR8Yh9x61el1fo6GXEAJy
jvOZSWY5ENlQvnoo0q8jeEBqKR4Jh3x0fbGVl6jFZdyhSozOnXAVSwjJcihlHhFSthRXjHfsRcW4
+QOnbI35z8msL4xaw6lZKZs+CCmuEXT6Y1+HtWYEs6j0PDTlOZvz+VvFWqaoT9Lf0NKGWkvvurTv
L3Rtf4Cc4xQ4oqv4CA6sDkHpR6AHrsjS/zLNFDvSesjEGUn1yVBo6rfD4JtXECWz66XzWQ3JH4RI
zrLvEXt5xknUs7ZoJU/XKwsjT1yrtk1wjQrfhqxZaCTgEW0ZXsk1wnKv8SqhPksx4thvu/w6mGn3
PVdC1aove0LixU/wDijr3hS16ig5Wfl4eP7FUSpfQ2JrkRUjq2Q2L995DkBrGeOLzqXMg1TFBDdb
8+TKj/Coyo6LxEhF9aO7kPPdw1gRCX7y41aQL+QEQTNUJ347h1w6PZo+tbI6AKCH0agYdPjdQdWr
zXhNOMm7pq6wOiFLNJtsjTCJ6hp3Pzrk+5c1E/YJAIc7FIB1eeyzQcM8IDAszGPfutbvrrqqjfu/
f5tvSXPyv2H0ZDqMHn/gLvnX7hnyeGFW9My/kcLTmty6y+cC4tLK93U8IIMGemwEuWnTYrkyXHoO
DJX9T6WYKwMmsCO6y+lA9cYx3zJ+YfCM3DU3ax/dSx3p76kWenfbrT6LeJ+CXEuol4nCLiGh+Bv4
BVSXfXH2yFtjKkWQm7/laZn9tebml3plZ4+Tl+0SKLfqi6zTKMJMzsHb5CxXWOB5TDTIrRPYBpP/
4jWhKRba5gZdjdIF665FZE0N9Y5PdorX+VfvE1OGilvhyyah8I8aYD0l75x/a5C80X4Fpq2NEHeL
9O4QIOMN9hsQAx8HNZ3S6IxTDkzFDoFtOzqOq4oTJ2RSKeAKww6vxKNa4WBjPthL9FCUdTloFdES
yfUJ1ivyT8vj6Ks/SbPXwXf3DYw9NThuPJwAhJPv4oPMEINZ2BWjscRp6wgrJDhub0Cx8ZDlQsDH
nz61OpiOLOyi1TUWPutTwFkRA/AX4rPOaeykzWPo61tLc9tvTE8vMP6qS9BrIRUlVZm8SGitQgn8
AnUUK2opp4amSAS0uZSwL6qYCHaYd11Z7dKKPw8TqLbNlo1zjn9h8LKOmsJObA+ZAzZdwvtOh4xD
66on4rt50+mY5qDhr4Uf56Blq4SrbzvSA+2rvuhiCOukaCEzXSD7HlAcDSfEAMsd9rIZRatBG5lY
5NBokyR13tuta1ydstyUhO2MZRcQNiImf5t0hnrswyP27yBicgM5Qt7j1az+KQyYKS/PbsRX2flq
bmUNtARpvxR+SrdnrOqdA9EvjvolyDSbBzx8PJ376kvFkx15Vu52hYCZtRkcrWNA5PAsofJz9OiP
q2SuD5gmeim4Il7+A4lH+6PKqVQ1P0JyAJvfy9yrYiErDbNlKX18VLaSM4hxCh1b6UJ3bRRZ7SsE
tEhQwZ+2rffUNC8UeKpKH9/mtwmEb0b+EmM/tlFyNHJVAGUW6aumSEDcVRs7MGjZN6XqEll+U/Rf
DQgJDoCOTTcpGRdq1Osc/N5kmh/K/gQtq+RVs5+2uwr1CQZgP4kb0Up1TYMW5XhNm529hurbkIWd
DRWI5ZxxLTJlY++jTjWuDyMRD7UomLLKE6qco8oyvY2tav4rnj/E0b5huOZ3Occ/1+F2QxSAEgyn
5QpYziwjjSSxRAnnR1RZ6P+YvUPC+NV+8bfsDuOhXb2hZ5vDJeRjbfU8Ws+Jxbc3xq1rr8pL5SO8
KFT/eubcIzJ7UdJ6WNdVFgetoAmfFhN50Mso9QYpozRIC/oqLC+ekd0ogcZowuOFo3VpdFrI7lQj
PFndDLUKnMpjeHhfy2wqkqL1a5ZXpRLhrEurZXDA+YCiSVv/m1MleIzVrf+oSjzJelDmt2Lf2EGJ
h8OBfbQOor3ZqkcnFCw4On6KspbBs04cUVVDu1m7fvXbSMHo7QE6Lp+QxuNP8Equ1lxSm2zQia4k
96Nud4uNM7cuaX+dmHAKmPMHDEC1sb8llmcwhoW1ReyhLkCxfkGK4zOYoJKqheCfGYLmEbM5nmvO
Gp41UZZ9Lt3UieCc/GUhuB8Gv3U2ZAPaonvVd58e8YHcEiHV5+jgUdRRn9soUVldH4y2/zKH0Zsr
JG9zdFMqeMbWklQzWEsjyEbQ+a/OOGdjMp7bOCgpVcBMkMWoQYTs6vlOhufYIijysLSsdiBx0vfp
sQGn+LjBkr2b1O0wEwTRGXnqI2d+HCoZg65A2nmCWA1cOV/25XwWULhbUd9/d6T6Egc3YcCUt+HS
G3iEGkhpQkuXbLYwCSCiPC0Kt2vnuWaj65qSya3sg1Dmc2c72Y21Cksj31kQjS0q6SZ+NLV5cDCH
ZG1cnBkS3vhqX+f82qdv8DNV5l05G4RGNQU/GiobrGyVBOzaG8wg0D+q+tY5akEe3zh1+QTvqg8g
fsuOeoMG2hJub5GpqRcDjrQvSBtlN967oiJUQWXcFij1pnYCB2bzIcub4nrF/neiJLWVoY3DnG+l
4hlCpujJovYtiHUGahKk1P20bFRa+CUAKIzFVIhT+lmINj6ta6fF6ch++vhVnX3sLOf8mYu+zEL4
aiFGupQIRuCa449WlNK9k7rm2braV/JvWhvWmmDn9KD5rO8aOuTs3BVjo849qZDtBKbGEj5Ye3T+
eFVP7JAtrMOiMiRnKdIFN5k94/ci2gGHAFg8gyjZryc7KaRsbQuCG/myLCwYbUKFJuBt0D7MGQIE
BSRuUhKulxndycS1sck3yVRYyD0YyIbYfzMTP649bjrjX0j9/9SnoP6dXOJgR/kHHCwSlLrdUw/D
1lYSRUaRWWnZx59oVJP9g0noyhO5gtEbiwPOBjy1hyjXN1shFb2WoCQUTpo0Gd7HC9rYfK5KUJKB
iqNsLjOIDpI/l7KvrDdzvh0Aad3iDLrjXog4bloDYH+bO7PZWp0dlP5/YfpXYdt6iPZA/WImYFQv
4NWzRHT9llQps0RR5sNSoyRb3b9nFU5qfCtrVjm3095kTKXT9iuBOKzHxEiFNh6qvTWGGLtw8IrR
QyHWhhIwUn/dKiFk1J4hfHrV6dKf/SIxBb9lhb28FobXoauQtKqNiDHgNgfAvzeA0m3pJK+pshHl
eQmfybJh29Tvby+DOOoBTLU5AVQpfOkoEVKRHmcu5Xg4t1O/f2eMvXMt0FikXczk3cOwBt+09r5C
vtQFqRSo2G+XgnEwScprAqVxxCZxjro/aStcdjzUREa3VAud+KmL8KjN2gwkhiVmUWNnwhLv8gHo
mFIVyAQv9hEEC5oIfwBBuWKsX7r8Qy+/+uOGQQZ6eXcr4dMr4KO+h2zO2mw7HbI33sIgrdYjNy6K
ewuWVmmNT4guI5mYztqq72pjQeX1BGbXlLOcLOT85xMaVn0yuprXjQEu02TKiq6WhZ4N9Elp43hP
WlHTixITynQhh5a/wO56qk/qBCI5kxdkLdX5BH/VuoFwxV/LPjv8s34KAPtylvxSWlApkG58XpSC
hOjVgeme74MQsKNHRQgZBX85etsORT8zcjPMGIE1OUCSNOMmxeIST2RKIbKhtF/eOSo2SqIkz84M
zwHM3we/EMuWvm5+wJSwy0foA3YPCwgSqJupu7SY28dW2E65mojwU5IC0UPPo0lmki1VQegeKsoa
I2DIjMxPUK8P1/id+tuXjxia1w87Dy9JO4bKDAvqU4tcq8rMf/qjRyoQ+XUlLwgwYUgD2t+yN3l6
5uDleCOwqwhfc8hjOGjrWr3ZjKLuh/nnf5u6UnURbQwv4C5zG4tFx+9VpOKJLoSJJ1DEBilcTAv/
r2RQxiHFpRR7/TZfCkCCFIkKFDrymLNrKvyphavJuFPvvYozDFO6oaTaufe7FAlLiHiqoJ+q4Bsu
E00b+T5vwMReNKFnuj/VErwfO+cxDI2dvrr0inu0NfbJNcQZZGTKcr5iHh8nApx+vRLPQNYOwNYq
cTb0IoCNcJvK1J31u8sGFu6mKQFCX1Szsl+dcjy5bEhkRQ9eQwkdhAZugSeJnAG6PYhlXRMUh74E
PdC3IeOXXszx0pQnpkw+c9xKtZR6ujnX6nDibADaqRC1UZ5X/6U6wa9AUJNKW+qqYFn3K4k18QKG
fV41xWkU6zUdeWPZKCDhun4dNVtvBQQmNmTB5f7b4GeGuimjpVeIK4Qrnb9kWTbnOBl8rFG+wtOg
uRkW/FdutccNFBymKXo6/7uGcxkD95nS2YG93FE174Mpj0S9Lr65RbTmRCInoAB2EBrgYY3cnnhQ
mIXM3yNSENTzBWgghDoyYGN4Es64d4uYEcayFc3wkjILWvGDVHIfZ9len8kcQJl2yNKXRU5C7qoS
V+i74rvK0YY/rWPjO/R7UCkNEMtwpelfbDL6OXERQMkwmCOpfbNX54mWFt9TXoxEel6t75dR7Vvt
/gJoWDro3yLg5ZXOs3uzGqHH0TsmePJJXpCaYOZJ/SKZ97Wd6nYDc70T670vnU3NEScQvbGLaL2/
MX4mXSZeRlVoUQk1JFobCvMTHe4v5DeC9+PxJYNH14husa0jMoSKO8VWAS9mm7+TyxjKxnuiwSp0
CWBAmgzb8JwOmDOjmKPksgf+sFv4DyJEEnYhSMAqgjpKx2Qw8VqMSipaFQmAou81IFjMrNLq41Af
Y8DoIXRene4HwnPicWXJEbnRNKPNbExYywllDTvHxFaq6WT9QV242ybBGYu3kUoHRi8GjJgpZ8Iv
qzcTKceRBMzNll/REgoT8pw5Xg5T223K2atuZWHLysIeLDlzVsw2hIeYmElg/Q05LFhy0RzhXger
AyFxyKl2NiYx7DAtWkDYTQJU4jcFe4SM7aYoNSofnVaycLQAIVtL8FHVZaVcWn/SiWxKO12TNmoq
Dwltw+6D5Ds8CaBu8ygTnKb84I70Fne7FMLtnW31IWNdkinQ+DuEqrwIJZKorBjnta/Ug1Wel9Om
aV9/v3I3r8KGhBm3iBcigvvNMoF1o8ngVrMl9GY5fJ1H/aSbife2SLC5zdWVKlHGP6CJXyu0T+YV
Xud2Gohnh5/uZF/JtCvz1ELlmFs4g7nL+FpHyUj7p5uqesLz6g8LIfbFnrkOBU0scstnU47eQtch
kGb9zGA5/MQ6e2CxWxs/2aPPu2CLdVGKLxpRY/qZXf/6RoY1DrahTjH+FKUZNe+JhplHkX8x0WuD
BhbzAWcE+xeNf+Ei2tT1uq6KEFtms8y/MmIgPc0BTZQ+nTRpRs6/3kCbjvMQ9hpNQ2yG0fGJkfWq
oT4wLK8o5ipqP7u2SSBJzQWQBpejqxAFqFztARykwmnBzzyXuxusoEIrnVDHIohAqrj3XsZ6+w7G
QvP29THN02as/1Km5keaDdvXvygIvKeeou6fQmjApKB4wWT4vFb/c8XYiS0UxZRyFgZwBY3bCLP0
ObPRstU709K8+AI3ElIKvCv+OP1U5MopzNkh4OCmcF7NDG/tkwuPtaLNSiJSKAh6FCSV1US7KKGN
yjPseLoM6O6wcmJRgrMIza/fmWJcsDYREFW+XN3CPKyGc6lEygVFxsAmtKODCHqtQi5KxV/bxZuA
oP7ublWylo55LY1H3C11X4DUd8fFWENtgOeZo1xwHE/DJAcmCY2CJg+HZb44EE/afJtlFa94v8dG
iJbW47n9J2QTAklSlYUHakD2jREKqzSFmU/qbS7o6DcQtGoYmRCpkLWXnIiXRWu8gvHOadNLzvcu
EfDm7AupI7gRzO+oy8HP84WEgfJ9lSCmolppaTUJj/JdeJlSYs1nyIK8SzappwBJ2rCyWDqN0JQ2
DrHpaCKdRphmyieN+Me22AY2v5qtH+ml81ZL+a1zbcLa7KK0TQtwImbkCeACZt885eBV/ac0dFGj
VM8XOiiCfXyEZGD/33nPcuxrIotDjoOojrfpNJddJy8sF4puoqsQemSsOObI3gGD2Uk++CHt7JTN
5t0eXoBAjX68oN97WNR5lXPeWjRdPt/IwNqmFoaprySO5aS2KQD1OF5XFENwLclQFcpKSzhxKuaz
S/OKVSLcGoU910kFapczILdng9sKwfpC6Dtr6q092X11yAoQttyekcz9R3Kr3NlZarohS+jg7NY+
vvToxyvvpBkSdQykf1ib5OXPHT1kmwKDsbKZyFV8Wi+u4cx49+S0JzSYyjJBwqiDLGGXOjqchoml
MunMSUB7V36KONlxpCcAYIwOWfCDJYBeAtp5XuVcB615hjYXdLZGbuUJM6CTMn3bHShXxdjWRiSz
BQ9Om5LCMV/1+HWV4OM9+DQyugHzGb+69Rex7obnJncN++dNtbraFA5xNQh8Z8/eQ/gIDCQOHOOu
JBX0gd95SDXgJ6Ujr+4lgYR9UQ6HLu6fgbmtBNftha0GGsYLi8s8Wgu/Ji3i9g5uwOAZ7+dXbH+G
UNLXB0FYGHGwISre/PSc7BPlDcQcm/SyGOSkysmXMRS9JunmPZg3Ix371LYWMyLTYdEZM7si13Lt
y1T0/gONGdOcfYcA8eKdutAOmXnw5RLG+UxSCCBiiDD/jdqYMNNhRrsYhkkPXt8WShRjTB/tcs0v
yTsfmyvWgG3u5AUm1EPSZmIxPxVdkvrlxty+wYzbg72A154a3zw1BhTzsBk9dO7LMUt4R+MZcUzS
osaxmsMTW0+ozNk7/PamchJ1qv3vN2wiapaV72XlTBfCcbx0sl1NZgLS7x3UJi/FsvWofSdWyIW8
gQ+Txohi1NhlKQXf0xFtYDJDk4xu/18iYLgmK9hPg1bWS1z/msx+9eC9irl4JhX+/pRNmlSBC55A
guB6FyJnEulE+Wp0q1T0HT62vnY+2hzN/x0qmpY9mVemDGaVFG59f8W2F1cai0CrsS7elMVL941K
zTKNc2A67/lSdo7Qa71dxEl9kTmelQqqMpJ4Hti3pMq0E7rNC7TteN0jiGSpzsTWTiHrGmJwHd0u
KEITd8LTZdTG2AgRn0NogLoQUItJY6ZR/FmH6bdkbe4bD6wRVYoSwzR57jWCLJ4B5kzNkZFGvDGG
ClGmYcw8veLHrPJOvwqPZqpl9wIqoZjNHWxFhzdo44mRYZM5vaiuRHR2hbUiDmm65tckqJzB93TT
behomrVzZRM7mdZtRybrbQY6+hxrq0CNgNRL2wmk14PVUNe4FlAPvZhlgp/gFqYU1gXIxzr8uhkP
o/3NkHAP1R40uxHNZjda9NTKL6IZOQJNHA90/uj5QYzo92fwmzrhtWNEuYHK2zMUZGDwITe44Io8
jmR5Re2LqnGac8AmUAwLTDm9jMv78yaeBMwsCH0W2DKzZMgWBy0MsRyXO5omMa4vLi58s9Gnmt9S
imdg99q3lXgku//d//UiyWi021ux8k6gYKBQ0fH22rcs2Golp7MqQ0noxK/VbPXQdMSVPP4a/fWE
oaxgVDUlwu1kbFR8xq5oITINuz8jV3ZtOdGoYXAE52SisJP9vRRHZPmy9l4T+NUl0YcIWUvzeBGm
RnfXg2GIbr92z0Cf3s+ZpWbrO7avsdH9sWCcXbFR2Jm8HTbOihZIU8zteUuBN+oK7RWdcVws/gcs
3CD3tEMIHZsxlStgPfy3f6Tc7X4tw6m/PgzZZVEabOwff+oY8gny21KOK1NTYkXGbRIFz71aVP1W
BPTzN/HABagSKrIdbYDYYBZoBDzpHIcLRoG+o9gH6nd9OFzohQxOCv5Wn92J0tjmAP3jfRKX5ndt
cBij6l4rZp8W+JbVaqWYrHUunI2SAwgaV64VgU5YepjM2N/NCQ5W5dgXp/VeBh778qCKHXcSn3O0
0AHfH60a8SLhupm76zWv0hSj3efWPhiEGG5dyT1BRHlW4MiIBzirY3TXy78AeqtRhSD+1Hh75rk9
27DRRdIANzZRivBMnwAa6+q3s2hVb7/zWilO9AxB+8g/3cGhks/Ec5ZhF0D4uHzNX5oMRk1lu80Q
HB9YGxf7vW/KNwaFihScdz0kRXrQUIju985paXuj5j+4uV9RZk39yez79gioXoyydv6lqyLHxqqL
PRd4wEynKE5+kJg52i4bmG3Z8sPBiNLLUFwzolyU/Qt1ov4cKnRDGH6ZYOsm1PV+FLnG0znQgJHC
ViL4ARki53Bx9s85q2JE+90E75V19Tgf+mCTmL1guFx7xvW99xN7CmlDixhGaoK98IFFv7xlExkm
kldcSJTsrGJC95VdpEjk+TWraFXnzM9mB6kshU1ac3Ol+8i+k2ZAWzIgZ0ZJuCMpmlTO59vjdtDU
RThQdzc2HB1ygG3LVfjZ/7KJs0qF6aOdezLDFdrrN1kqhby0BvywRYpv1tFGOHb1H6UkxVvD+nPt
h8mPCWSZ1SirnBFAcqewY5CbugtZmBVly4nwvdZSIALMJNkLXYARotB0a/3/Jhxgp0KXjfcx10P6
fAUazzGPsckwBIi4c3jwtaSBo3en0A8JDtfKOlIbuYL/0hKlagWEvi/vSorUU+cvH4zZsvMmNWJO
aEda+xBPq+aPbtmxcL0Y7Lqbge21hZ6DB8UKZ77SY4vg2Tw8lhI0iGbywJVAmBG43B7O2z1/gvm1
LQcvQIPALRNqXxai11OuHtpLxZk+2hGT0DhUoD6JF4sB+mRddAY21zjG7y0QMz62Wwr2zJfabldd
ZjW3swIPlE6YHszwmJs6Jqnqvq3v/2HYmzpRXbS/rUAtr8lJnlXN6bsksNHZev3pBnvlWEqW1+1O
OTPt2N5ruI5/4jelefjSHVLPJBwV1fPd9oQfvW4UmYeFfRwDPMCzOr8RyqW9U/XfemZfr+oaM/6h
eZ2v6OTlt4O6sHIUsViglr0u/o9PJUovr9IzzxvTp9o0nyP+znU7NgGoPFstEoVjYXBDb+RrRg7k
xEL3betG8caQrUFgMEDXKT5TaF2KUghV2iw8WVE3qc4G9bhPuwCQfofSfYiqTMMwgKqgsd6d1HI0
Q+1fxvw2D/8zzxUNjdew+Fs1L362TkossxfcxBEYOx9HuuUHDzFinesRNX5dP0uT2mH6HzDyF7AS
KakgIXj8V3GrtoM5rsxQIianJD8XEnbW3MqO3WWFaXtR4XOdDoTEzaZgKwMGtVAGIKEN/RF24KR2
3Y+QRvNJjdiXRMww5I5cDRjV7kkq+niAOuPiZ0eVB1/SX0wZUFuQHoVAuTLF/JTio/0OM7arnh2c
jYdm0SsjVdmu4lx0QEeQFIe78NREM82HNLJiKt16AsObO189fvhVEOcfUX2lYySSfpVr710Kz/+P
LZ/kLcUE1ovVWD1i8DtjDFHwfeZ6CQBfbrPNCAdF5+Rb8uALuRBX5bvcTIICGRbg5k1HjHf1WDOk
eUQ12qtE+MccZqmQVidNVd7UXtQjVcqfl+Z+rpw03jHR2Ce/64qnlS+uKu3a2taE7SR60TNMlTHa
+tQMleVSzIa48uJ05tctxQZlTIlb7SpnmZSmF1P3zXD5smJBU9VWtjzv+/kXDeV3qIn0bBvRErlr
pc0cL9fIsli4Uhm71XtYnDLgTNdP+Z+rWNbHh1Cl0AHD0KPOT+BcpcwwBKQ5rVxr2U5+22D0cDSQ
AltCMyI4KTA9hk3iCz4hJJofJAr+j3PYBTMXkfuo5nt0Wfjja+CUVAedTIaRcvdYBrUgstFUIp1F
kwWYH0BmsZGIcJckXYF3Ox1St0PgjWpmrBMgVA1FIbMzxBduGodFPgUCe36EQXZnvQopjBFy2GpI
bZWOL9oEGw/Mxo7UldLglXEOFV1P8tHzQ+BXOb8Q8G4EXdKmvowPgwy1ZjGyW7oLRUVb1B1i0OUS
F2iq/MyWJF49cmEBEE9o2qaqso2PXa9F/595Dxlm7jYpOMC0knlvFBrTpEq3A38kZVbMja9eHQsF
b3QUd6jQ+ygBafdOYL04c+LLHmwkJBBf2RopIrcFQiyUOpmB2vIxSweOKs32ssWVOuIvarjBQHTr
IbGiRLLOW92wqwa4Fty9xvy31TyhR9uiRa3FmH0rQHi50ZPLqMw67iGbBw4l6MsmtIj4AsEOFKPD
CqpE7arfGv7wSHZL5oHO25xPqmMe/DZyUk2g1vxE0JyXPixaBSGpNnN6TTMx4MGKm/M8dCDpfQXG
c4exsfK1VUIT6auGHG1IlBrfjrXrjTJw2mG/n3i0pcUKCuTOMvjLV4a4HWusXMD4ypJu7PH9Kzm8
R3RL35txLHJaFtSHdozxWb5a0pAPI/dEm6VcRU6Tn1yAUcRu/4LAmhKE7QKWDvb3R/scNvAXzQwq
vQHrl1T35ANUjABHAxlK/hhlzjKpUSG1JGfXszQjGyXUkdpXcKH98IN7IgRFbR+jEU2+sanwN9N9
rnrmv+Ixhy00ZN9BgcocBBWqq4JFpO+5w9FClC+q2gsbekZVeRzRPU5G0Vn5LAQ244U2UMo8ztmB
LSzkLZxWRA4t+RmooTmpKcU4Ts3Gqpmzh93uxfgiKu+r+0DBao7J7rg8xtJdnV2RY6Q8Kz9iwJ6h
Yk/iVb3RnnFJb85B1IAdEciqZOTAPLMexusZviyILIUZB3ZzwhlXkAAK8HtmROpuDQ1HH/DdCXMo
8QYQxob+ci48i5JPJTp/FjLYQ4wlNg/ZI4H7L9EBU58O7eb8DeF3hiukBd5pcRH0xZe+cA8ubvKY
IoISTpw0UzQqkYqNH2GZNw8Edz1+m9FwEB+8PtGrV1u1Lyr+mxtN+1kYVblxbEnJw+QFPBxgxC8K
LMEzMHDTWVl2DtT9rjlyP1wVufSS5OnpFRpzn4HP2UgCnspulDzWctytWhJal39ptI12bIX4ENkR
RLmJMo/M0UcFs2yUBugxfxo6y2m8xHh9n1+qRRWYj6qXohg4OrhVQ7tbhZkwHSigUwr6WSJCURz9
VJj+WqQ5gd+cTZmJBZoOpuYeXGoMqfkKlMGb00dK46RE1SeIShpI0aVwUjnSr5/nNPZwXgD6EYpq
jhI2LdHM0GCnpwqsO8VYbrqgS7koPPYOpp9Uv5kKmF3wSsw5Od3neaz9sOhmqu+SZQPsQSIHiDQ4
IsePEQIjG+jlbesxU0uVdPnFKVLM+jugpO+422ACHKl57E+XuVzyYaKUId5fmBrtuxiH2xQUPoZ3
po4IslYESEg8GwNW++FC/v5lpcrzPonFZjbJFGhePQpI7BM94UTt5phZQH8YhaJeikGRfxo3baCh
O24tw5EUfoYg2K2MjIWDaFuwcrze1z8IoviV4pdxF3ABjUCZjvXt5uSxzuIjb7gbLfh3E9rQnIUI
0ctiUcV7ofv8UWu631HCDzyCcDSzqDdIrq+vWBhHPYAMyCfjUthF8hTs/8IKWApvQo90/HPAN9AU
y1KkvGBbX5ywf3ml10e1kP4QuQj2qgwH2LvPipDrJSydygj8WoS2kzpceeC4Zp1NonDlE9PMpDyf
w7a61rzyXNmpQ1l2d5fmPH4VLzvzCaNLv1G/mWLcxd1t30eIclt1/Q8ku5B9b4aVA30kY8ahQazs
rL9cp9I4LTAVWLyyayzHBTXeykEPc7lONdKNSggECIOWPTYljZj05W19XNnt74wPkSN0xSx51lFO
0paPwK1Qy7YX2iDyCU5pcQ30rRkdrIyQIBoP2WBl64Ak+nlZn2qiZE0T6lB71RTQ+5jicWm8PUFL
2LWxiySKJaAxfs4H332QwUmW205Qfgb3LHfT7PgesQELZ9P7bBGBONre1psWnNFHZK7qw5m8h6pk
z1/zS5bJxUTvMs8TP47r8fbtOATM+RZg9PkHQQdGuTAiX85ztswfvtqR57I483ISBMWE0FCuDqKx
xtkYTjMCamPJnrMg5lc3wOtwE4bCbAvV++HAIg2xE/7da5mS4nk5N/1blvkUm6o+/UXlWqczxF4w
phm/MRzu6HpAZIEy0Wk8KqLFpkZWvjfeGqyya3Mi7kgYHQQYRnxfzIB05A9KTTznFffMLBpNemmZ
kl1fc8KeYyTh4KkxaoSpYPz4f5Myu0woTOoS4+LkKMVF686s/eGD/CdgOlL0yXwVtIl4jH0QEsIj
HIz8DqdztCQbIqbvn2AMSDCY82fMEOZS3UKWWSIwqKXqSf9Zl5DBzSjjHoDRN5xmQDcqs+2jVPeC
afLA1fqqJ/6Ki3XWZAoN1nRLXrvfp8evDI1t0hbXcpg6FZ+lzEmJ19nCJA/ItM6MfVwjQnSmahPN
rKpea+v31+5jF4akb9vXFhEMzUbmbOrVo37Lt2UTbpVXngRTSf6YM6+FwPWfLvbBMco3sk2bcggK
zACO/cuESEM575+63j5L4QJkJFClsfje9V9w046Au8XinjygO2u+dRSLthJJibJdCpZ83zwd8Pkc
F3JYtCNhUGf6y/jQJB+gwXuTeW5KLssg+koLKIYfzGiYJn4o58iuQXA3/2M803bZA/brD8/aairy
DIVQXSvNFNFaFGZL2BGUVniM8wepAsJeCLKvkj7Z9PkoGpnDEM39OTKBtuRL3wHYZvTxQ5ZFKBch
4pm3O2HGVsXaUCgesRSWFA51UVvLswvIVp7DHUwzKtqVUVYEQKBOZ9YQwNo5bMZZsx3g15SuANxQ
x6ZjD9j4PmTn/ghnwZdVGpHcgVoifoO6NO13w+o2nI+EEZCi3eFn4T8uA24nQKOFP10qwegpOGp/
MHltj3wVL5Aie7P1zwCT9CsFWNqJgRE0IwwoUXB3T6P2ihL9vY1Oppb6ES7uJ79TqGnuPgoAxMz+
0Aj53gGj2LN/4rJcwCZNZZBHxcyRPHtMJFTmBsA4BQHZj8uOJpkj2FkPiIClumjS2oaAi3SzdmWa
bVxRwX3gXDhbW0NZwfFuy1AXSjBu1idz9EF68FwE8s5uSaV+jMxYDXL6davPj9bXyh2psH16jbsI
QIYoDpGAk5Lao0ME1vi4tE6cCQ4zhQ1f8iZ+cPApx4eyukCgSZi81d2/kV8G9Os5Vr2BEpG0SsBw
IlX0XAjTR7ODWQMk7JvTs1+n/IV0gQDL0fRTMVbMWFA0dPeBoisy8F1ScbkxyOI1EaDkBe4+4SEN
3A/oHqehrSsLMIUS0PlYJvgDbR6FxTPXFkf9q80SGRGbtOp3gDw7wul0W9NbxrAUyBKge/p82+z+
v2sABNM+ClvVIy40z22vNQw8qDvGVPogDI0FGLOwAEFLboRNMbygoMrY+wLk+Wke0Sf5h1vEWZ2l
yBTumzaySpF30Ci6FZVYvLvkTUxSejMqUG6duyGL60ii1U+77ab0QIKGGYF39UTR91qpxtoFdaO5
Z5WfdYzUdLvh1OePtkd0yPP071r+qpBmEwHRDyB1BdAf/1FJMPR5/YvkPQBDxoYg6CEACNrjehyH
OqKfAtFDOVlLuzzEoi7qtIOe55Ft5jsPimYiDWuGIKl1aN2ZdF8dqAa/9uE42T86Io0HSDolYvIY
oHEz058uT81RaEO9D8Ges9V4DqttPTEj/M9VTT5NlDM3wU7HQRBp1DOH506ZGVVIVejzShz0KFAI
T3fZKLmOZGst09BGGRj/9AtK0uEHdNYLsLZYsjR289bdzXpjY3+v7r/4/zvbkQ99XVqWuApgjZ/3
DE5zfU7AD6RYO3KUzQ26MabOFF/xpJNuxr7FGewgF8LEGkfw2Kg546VoWROo11xi78XJyQ8dHIey
8+0n7JyyH9tgonXntUHwBn+5BzhkU2gwFxRxfrIJ1Pn2AwU6RdeYTUTXalvvviQhqAnuZFoGifmw
Foaq/wAju+fD1+ogdSJ/y6aaUUz/CoyG0k3uGRFRw5ZUntATN4JPKukUZvGrIb4dj0ohj0cI6qo9
2SDzKCowgG22v8mc8P1FwZXCqM5cpdV9Yh9brfihhR1DTLOnFKr6hPT00ehmlECzRljG2Ap9P2/O
W8GUJp/YuK2irrcNOUA922/keukrhf7WDwgkjvCA+AuHsc4/kZ2LImTNdu5ONTNh47NkVhFXI2di
abDVd0iHT32YDuSvhuB4qK8/QdxC5nU5wzeOZHuHBq+UOQPe5n61vWcotbad1qWnJl0W1jh0jZfq
iSMxFq2BOEdsONBFeaCL4FYEf8fRt4eEeI7/NbxnRF7nK/fnqjo8acBZs106znSslNFv5qHS5FgG
LtgP9RNiCJWJMcnFrD6r2lNFsC1YQmWpS0K+EZlduOIpbXWmb0LWeyWXDdLdk4khlK5jcbl+nJvo
vpxiUx0kJtZONBO+3/rUwCORumtUg3VL8oUrG4bioShhdyugNOwA2XgonpZ5LbgfNN/HRI5KIE1K
O1wAPCKmPpILGzjXNKWFm3tiy47ozBJfOog1wDy5i7VOLJT73mCXOaIuc6Kq7+O8i7Sjxz88wCNa
8/bRJskha5BkHcF2X/7PiYetjxwIJs0F5R0NNL0lMetYKPNcXbJBdjT6cblkglxkkvOfxfwbmNjS
sL+L6dtSEdFKfSLxgUAX8F87e2KE5e1tHm9E7PCBFrXlaLgg/Su+uxbaZWKJ1wTjFjaoBpK8hlvq
Mdvj1KGNcBfKtdqJe1fmFgh3QBldi+cDs14AYRYkQePBYx8ecViT95aaoPHiVjkU3CR7a/Yf0ytO
HNHa4p1rwZT/AXJmiDBFOfC8giNQOWfpsUzA3PZ5JNbuLIJxEKAd+H1QkNz39bHCLg5qB2K+s+hm
pu57PI38k46Q23AqL5NnYyulrPRQdOHW+vAtXJjEZXj7SqPzFFF4ZcjPC9pa8F09dufauydYm6jT
29VpODjoGVbt5Z2J3FBZBX7Qrt/BoHozgZa7hSEB41/1tLupLGIAZ5BK3QksBNxliblhWpmkGwsB
3vTlGb0ErvkgJnpRS/dLB2ylk1gFQjR0hDebJLd1BZoYRU/cbxqMVuqX+BsF068TPtE0ppmN++rQ
WCNwp8BuKDcVnFlQkDjaCgadlTNXcV1chX8yiYOqzYK+S7BLkMkMLNhzdkp1A+FTLvO4RV80PVSN
jPxLANZIg4fovpe5KKK/7WT+bKodlhj1+7BZYBcA3WN0oCccFm3QgjcKWycx6HRdsuFoUuD9g6xl
pWfQCRgYuqgvH5nYU3ewD+SQd3hEyXVm63n4WgZV+eN1uLJbW4QNiXpMPyC67A/Hpl0eTVI2vgDV
BRdMpLx71Tnx3U2Ppq1ZF6Z0PVQyz1ePYScaIY2yGQsC/sShWRctsV1J3B2SgoK2nVxViFvEkA//
SdJ+2wdfVy3JM8sEOqTT56gDUyw9ICS7cRuDE/GzbBHfAIUE+6jttQ/zSlnMGhMZvtY6/MZcP92K
Gc0lOjgrKUV3mgKY1uE/6me0FtKiyB5QXq2GCf1ubRtKxBgtbVGQkEKz+a1I0pqfKTKINEHcyxkj
ZlHxJmvacsvtrepQUQBA31ZG7wqrQjqNIEKbZHGsf11GwJ+AmgNpsg0F4hGttbrJBgEueHQRt3cB
1rsfEkuKq6nY9fxzbloTRGf0ewBzzPJwgySZjCBKKyoM4zRGFggl1QvK/iZCvu/OCgI7XOcQCNxn
OLsXyECfiIuzWWL0I/F6hzh23TPQ6J7YD0EnX24IJNi+OCylRgRX9SqAMzBw/2idtiD1zKmcXxeh
IFk6Sw8Q9J19vyBTvoTpFagjhx0BY5qfXO7iDpthUKRdr77fZpDSk6aaa7JJ0Inc0hnWs8GISgLh
Dkkf7DvMx7mvvwdZ0unle2cWlrwQI+KqRMBnetMVFMdSZpvgB0pyLpNca3hwkc/J8O2T565rYhvi
MgPDT/IGUtkSPU5ADfByoozF/5eIOorwXNLh3C5V7u35nO5ksp8CyqXDmQ5OIQ1DtwI4q3ydEVO5
O9AayD1YJAK5I4wXRprMng7g/eaYV3Bef/X2ja8CDo5ZE/WDbIrpYVmVBW0ykM6VjgYXPhalxP30
FowcqdNKPheTL4ygNH09BlUZDobE3vvHVEdJ89g0EoMt8umlqduws0XmdRczBv0qUH9vnIUYPkR1
S1QchvS/5NbcPXnkpnQeZ+Kfww1cohS5r+//AdVwLITNMFSssiiWcwupSjxBsO9zfE5kzBf8SyVU
JXLm+YOsqhYgw5IGp0Zy64ZINdkV5ymTlI+tXOKusm9Ru2I4l3sU6POcnwM+j637hl5wqg0DYYUo
Bbr6VyBMTpWBxYaamHs61ZXvf4T8xeXVJEMy6d1H5DAt94h3Qe0NyG8AYAmU4RbVu26IF/Hru6hc
dUoREHe30FGYcdy9neoqybFNrgPtMfzYKomINU8Mt0uJVaH581TyNAahNCiJfc176XG5Vr8B+LlR
IqVvOR6BaBULYBCyvaNbCAOvBw1eLQuIiaJezoq+LDufztWBY7pYYix78X2fdQAv7qaG9MdZIMRG
TB6bI1gmRiulnD9RM0/abwN3RnC+H58tahsJ3BxMQpId34eqZxiJLHRQgIGm3b1EtnUpmWEx1PdX
Qhqar+K0dulLjxbfY6ZKKka6+YIX6ZiFcR5sM0mvj0gv3ycV+NSh5GBpxudj0+Y2E5H/KZINHmUF
qzcAHgZGP4neyY72rnTdxSChYoi6KvcwCyIVKKw4vr23xEXRmEZLtOY9oMl76RZw1FewOHIp2eYm
oGGyfp6s+IvLCuKAhifBk8eA7yekmfm79lVi/3KWXwni6+eHt/0ZIn/mWzbpLXrmfZ7GQiS0gaaY
Awg9vI655yElS9ibK0Pfmir2c3DxMCdIqXrwP2o9zlxjbL45qF2MBNJCbjkKwd7OIrVKmLPIQ5oG
FnLR6aoUibFkcbwoR/g0dY9oSHuvZJhX/aYpdp8PcAio1fLaZFK8OAYcyhAHpG15OLPpUVgH5CpD
o1m1o2cv444XFZLRaCaMMtpl0jF240w9ISarFH6tRLofLiNNLih/7rLFjuNDFsdpp1kfYN/fk8ei
jd+6ZOevyBdKVcwGTL3LCYgGxXQiSFtHB7ERLfdFne/CT/QwsHXEgGymeoD1IayH+wHEZqZdJhU+
EkUNfTG0wFXkokJjQHAf2h62SFYSrpJLKi3XIZdus7tv/yIdFnsYQYqWmgwlGSHImz5lPFZoms+x
6YpAq86674bcUjCKAaDy/dOPqKxTpMZcbA6KaWcEXjZC+QAqStGtzsCzAfYfRbSYHTGCeLR4P4SY
IJ6xJxk2yxby4mh3LseMq9QAjSCDYwU6uDPZEr516Y4gAHoNxcvSiKX5lY5hq0od0tRw5FQACF/x
u3Z1M0l30ZdKYOjkdfeIrUi+hhsM+/btJdTaxt0x9H87p6iy9s8vnlpqTLE5HS6DIxZFdGp/b65F
VHd19hICEu9cxDQreHOfsn9x9/iBQPwU5A/7XmLgMrUk35L9z7go2BZUg47Mim3nWnqMZ/xqqlKS
+q1JMhpGvR7Pbs0Dk/k/WzGgi3/9MHM/HQPVcXjpYYJasZj8xrSP02DvIH/vsZ2ETzf2G6fYkSol
knrabc9rH+jqtIqVjsnsnz2biJgfmoDZObdqvj5Y5Hs611YwR88PaJt+deWsr4IsWV0ohVzIsz+p
Yl44LvC1mtZWm+3SyUDSUPc1kQK1UBVlmGQUW8y45dyB+ObG7k+QuLhKtuiyBUFLJYxi8/Py2ecc
QYWBmMRuetcBQHU9nfl/Os/eczoCFfO3nDvrefSrcsKKbgV0e7qdtegUQ/DFDj7SbOTbuCEBgRAD
Xi0g9xytJ6URWeJkSZjfO4BHMwUXdvVPZc4j58JKGmw3TrIHMB4yp/g1aJq2tiMbEN7YgdIo4nEM
AHKueNLHaBm8bhmvuu7O7qCHmsETsQjLom4b2QWCKh7ZvlVUTx+JbXeWNJw7jP52/zEDYMCCiOnG
izVnAC7GnDjCJYCKocjHxgihB06xSvzhpUv/3xUa1FfGcZuVbs6ESbymjVf1PrlzXtHI2RSZoupf
83jq+PV8kL3YebZgwg1blUUkhS0iNYDctHWK6EmDQLSryM7tvoLQmMVkVrNeRKVJgSDoKB8bV5ZB
QF313sWSd6nPCCNjq6+wqzQ+NIMRYJYwi3v+4MKXNfIrqS7BKoNLcrf804CPtIwIOTYmwnyhBz15
JlnfLaNlmtO2ttQk024SZ6CGfzoyZ4/yNtAAXi/4RahRPi7GLJMaT/oXnlO18G0UChXuMvx7Bp3Q
/eRXnV0yrPnD70b6Vdq/py7sZHfpP1R4YYLSMuYtKZBD90DF2h05l5S1YicTFGIqj4LRpbIPmsyZ
LrIG9kzFNNxFDbAMQ5crSuBddG2r5g+0dmWzEAcP8NWG5zyCshrlpYwkt6u7/SvWr6FzANQ1BkpQ
zv4fUQWhJlTNFQJBLSTomAP8NJeAMsGV+YpMwvGnHq/pFbPjHBZFuujVN2dHp4/cQGboh8pgRT6+
/oUw6dI0f5I9w3TIhOvPWLY/Y2BFyAVmybzFqq5Oj68su9P4F1KgqLOCIkU1n3QP9TU2e//0NYYN
9Seg0jyN7YF1KZYQ3RSpn7avjTcAblE37MX1At6Qd4qXB6l1yb+O2AP3hOUPX4YtL+zpLwz7Y+Ul
xiPuSjGs0IR7xI+8PlPMcHWmeSsyy02fL4okLNJekb/K86vQRv5JX0QsoQYGpsxxc0AGspztGu9i
sYIQdehvjcdUDbfeovaMrlogifs9Brx3cEWo9nLQ+9fwIAM+oKcqWs7K6x1v0kzYcRIQcv2QPooq
Cv3ZFWfaaOTjSS6SnJHel+b1qaqKderRYJlIZ+JR6VYA3uwK1GOxaNe+l0GpyU+l/t2x20EVf4EB
5lbSBpC0CM9e5pDZo3LBWlh2jG3oYGnrXu5c45PXDsMUdplNRrpFk+K9zgJxPjQ0xVEOWOuBUuRd
0EO6YGGDm5A8t/YE7zl4OyQVDuX/EdAswAWrObUNk8eDOGzo1y2hqENtCBYayRW7c/n/1Ixf9fKI
ElBby2CGJc007uY+q59TtdDOhGHl0N+jawBfHAEMjwZ94tE8KVp6ye9GczR8NBnEMDTA6/0jPgAH
ePRubCjA2ZjWsOkE27lXjSnuG9Bzk9xs2+5GBksrbl2/ziymO68zSP7oWOmUu8wy+TBcmE5X3QeJ
YMp6RtZFyo2BhMy1xoNTeJ2ucw/l0DajZz+Trd+prkHGzTnaZO67VrJ8dMXRdpI1ooVZRXy3bR/n
R6DgG6lrQu96vIOzCfFMhBKIozdiw+d2/BZuMupt45vodKjyFaf1FFBsgrS4kZ70etwuyAsazC4F
7SJlbfYbCbpspbPAkGs2KU3bIGsXtDj5AMtHQ/ohavD/UcN3aP2VwuqKfut5h8+pPRPjqnc7UV0D
J2/KaatUnq8JD0Epo+nlOsfLa8f7uJ0KU0aF3UwiYqHXJaoSQPKMUmvAeVjzIBS1uOd0u3fFvUs9
nsUjrrlsLXFaBiS14iCkKnZfhwhnjT66Y5qO3XKNvzBMOBdjn4CxSqxPLLz1BRKfHpx3Mhb4Sexv
bLJfbC+o8Xdky8sa7sCeJ5ZjiS3DiCUQLj8fAklL9kIYGYHuJg09d1wr6SqQwhs36Jb+1s0XAA2L
X9fbt/+423nsK4HtMedNE/0Whn8jR4JyzEppaWrnk4prIz4OYJ+iWHomyJfQZhhHdla8r0jIvc2E
p9UCvM/N4yySByhtl70SdmrNnuX9B7kI4gfYe/0nKhJTQPBZyjlruVfi/37S9iSkzmoXkbiHzpyJ
i11WkHhjiLMS3hRjwdHxjQ7xEtborrxrWb8sPhB+xjuwmPB7huzLspjexEzAI3HBvZf1kHV+wy83
WlS55iCjoO9Oj/1Zhdl3zcE6vMERvU2cdr7dlSeQAMrGOchXKZHA+28B9E8UJJxEB2E/2t5aAMVo
ILvlvq2iQtzUkA3fj7cOyc04wE7IEEECW/kgUPy3IsVbV9xLkYOnrA4oJwd3zAPQG1Rjk+PXABgG
/8K7X7lMvV2I8Adoi35GKeg9X/BEB2M/1zj18SbDGX9I3a4XOoHwJZi72YbI1wn+BufyvG3QuE05
0iAhPhKMtJbSTZkfa/3Gpdiy/W6HafmZHziTeaNpkMBy8YPZugCaDH7sSbE5TR4ESFHBa1Oat10O
609PXQosn3/KfwTh3gBmGvIscdHUUR+7RDzrjoBoPSy/htDcnO4WdZxMcT8AuK9VC2BwwFEi4TCi
45tj5BiIRaS4yb/yf5oNChg8otkd8F7OILE7W9kTmCR8NGmcS3H/0MK3t3onvRZchKlKJHOaui8z
D8bEQyWqAvDUPsHfaE6X+YnyVow7Cuk0Zkl99YkSghgEUIPIR5tiX17PmAkMwNJx18I4N0uzWvpL
xvlIXitxHN+j0rLFINO2y35PzZrmJ8TxER+/C+pBfGXdGFFN50BT4+AgbBgPBEZXumjUtzD+9JPE
C8ptih7xGsDq118Qwv9Dz6byDRPAiXmARDl4Ab0PEVBF3tmMzCzfLSBu3z/qu9D/EjuQsM5sFNOL
ZtZj7gp6hlOC1ICM5xI56GFq4lCO6+vMFV49rVqSZhFmyrQjdIXtIGS8OUqoTdpT1Vm9gTBb83qH
6wCaKbpl3Ru0tOvXCv7prszw4jRsnNVs74jodFc+jqWyxxD5257RHGDfzX20SXITeXBdH5PWUZii
OXdEvabIZmNxAM+PnyekGHjdH1S70f3IMCDpbxN5h3yRuiLQF4o0mYc/bF9gTvo+dWFvfVlukoqM
KrjS9jAd6VQUKMR6Tuqe67VWsgpCC7AsZzMuv9prdNTMqOuhU+IF7LhlQzdaCQE0ZTlPeb83mE6O
RCSpFU8YT5QY26KfjQXyUbJrTT3Dp2YUfbN2BzWnvD49ZaroaZCGu6MqXee6RpnX+yY8+tW/p6tg
B2w318likAlluKsviQ0YWt1FlHIWZqcmGI+BSVKg+IRAF6IGu2lqiY261KrjW8Hi+AuDBq5VRG5g
67Q/SpptD+y3MGW152j7i+n+gRg3vQVWKbyeBJWsx+GNINhgznlgGoJl9ycDzrrD5ZYNMFrK2Bf+
G52JXtkcivGERCAxbh07rCR6gUEZ0QNp6mj/Q9+SJtZ8Zxml1EVdfTcCRIm9Ix+53sfmUuCnbAGp
og/UGGMMqRuJJt+06HfUN+Ay0OAKrB1ht2aiaMq1mqahuWroRln1/JvA7KxXifts+HIHohrDRxq9
hcjDMzSAqz3bjWaCBxACU1MQkYyVrmy6X80JK+tobLMf9MBEN9MfdDsUAXudvW6vUCaOnrJVFNyz
5KCQi993PbOtiCib6VxLNMr0pywwSnCqYmeKE/kRGymovrEBbjCxzLdxLyA/WFDuvj2JeEXtCUg1
EF1aMByxvAiv6j/0cj7o6H+Gpav/M2UwISsuP5OJNdPB0dkLUTORrRiQbJVdksSI+TR03pw+3nU+
SXBwNcYTkrHMFF34IVKAgHrzPb72zphMnmlJLGBeNFMPFwFXsYEbI4IowOOMhfG0grFZtG5mPUnn
hdiSQfBpQvzlVaszkDKfFj4FAKulBAI87HXdH8MWfv1mydPoxl/GL9pznHayGJ8NIAWPMSBIX2P5
cW7G4dI4iEdMFt2Qx55QOR7+dMbiCvdbpKHp8SbjJmv86qX+vqiy6GQvNNRjZPeE/06p7YjYYt0B
BZ+OCfxvrbiUX6jk1x01lKNNi5Zz/oc3IYGKIsKF9R59aHK+bIyYnMKQ3AxxHyb9GrAK7+aGzDhO
qZTb91P5o87fhpijupzxdkY2bZRJ159gfFHuzYKcm0WdLvP0HZhEh6AytUQhf2CmeNP/NrAzJX73
uTkgJzGIKMrxfiGeC6m2Z1md7pPysefLzxXRo7Vlr/CVj1o428F/fLAZhNM0ZQylbS26IAQbVTXZ
7CLSYbbsU5bNoFopbubgl4cQqP4bSNpDfmDyHCHka7q+d0aE0YnfIcJLscXA20wWbVLaVutiLLgu
Y3JHJFtCihJIhKtSVbi5jfQPe897B5hYI9lv3KRQCgx6TEtaJTjNrnp/88j4QYIWqAbiRcKz32x1
ohDpUudy0LTTJ3lAjXn0yYET/KG/vrDCpNnZGhBjBgCYDf3p5b1Dctyp5fgS/E/R6f89+SvmIeLl
75ZbeXs5fxX10lClrlZa/wzKDyLu3uuMUoEnZZMw+CDPWu1ZJWNBOq4vw7VhziyIVdm7HS/odU0j
uGqrubC+7ATVqHEnZJNTkaTDB+U+zjVqgwAKEXix6RZDoVogYInDA7QKzuLncK9/XMwAOzsHVihy
KxsbDkDPNbtxYz7p1jxUkW7m3z3qUUr0UcAnsQRYX+ax22OU8BIIavQZFF63VDBEIkyeEReReQl+
nHnzfe0sy9Q3hIVzjJjcWpTVigolMOrI9HBTdWbJuuktYTfkgBoODJvBghBZ9JVxpzUVLth8rBtn
8prqAiqOy3rb/tsw1Cx2LNLpPyNuUR5+cqBMKGYRuo/Ov8jVv2pmlLEOGR/QC26HnWHY+Csk0hiN
M3Gq3lA+PfmXy12ueqamlfHHnZr3a4t+UegusGzkHIBMJTlKczSWLsfikRDC0uzTLX1pyswAMark
Sn6rVfbYTzSt32+f8fGX+6HygaerXpmr/u9fVT2w7SAiMq2e4eFIbVRxPiceto3BM4/JiaKwInfG
55nBB/BKMNyLoszCECbLcenrgSh803ZX6Whp+61LqAidbtEWwue24kmsU5LGRiJtAbgk2CKSN8Hw
YTpSk9EjQFK7W1wqTZgYMjVUDADRd76f9Cc7YxnPZMyF/uP+P91D5p+7ZsuKXbhqqHv/2wxVOM8v
C04PyC1N9odAcVgQmspc6fFfn3HP6SmSo7T79ThtqFOO5gI1Yw/mJ/as3u4QpUpj7/BrZk0geJac
spAveHYgo6zDAulhcbsSQcpxQ5dYkkIuGPOfaeU6GVDkm/Rzaqxo91yiLh0DfHwjaBrcgsUqub2W
MDLgsLsXOlfgyfWEa26hoqVHA0CwNxydfOLgnKIxjnSZHhXkC5iL/nqmUiGYi56YlHaGloBlBOy1
pKVKWFOuMzIoRldGclwGpsg+JqBMY49v37LDmiA6dkqRWxPkUQmF4ByecOWrP4Cedlec8HQJhD0I
XvqpDylgd9MrDSANi1DQi/1O6+n79/VCSoLz4NPYf2zUCJnb/x+96hxJ6cIAIRpXQcrSQ+9dppnn
gw0baWFN5pnNa81yrDBrA57CabYqV2uQOZKhL8Rq+Oo5G76aKWKDPIjMdv1zrUtTSOE4zv8fWxF4
kxlGr6gtUTyK227PWAsqBItbHv32DB+TQUzUflVy7LERMmtP/pgUvAVbnph/gtGTb+p6cKdp1lXU
1RsaLFCCxvlMfnaCxb9yBBjrkSE/uHAJ9iVMensKB9VzFH6JokU5/fA+HUEoTLoAvqX89u3nGxic
+Pk4zM0gsnvFDDiZhpqpWqBi7o6qqqvJLBCtrrqesuprZLUyO9o8S1oVdD5pltF60Xj0eb942yRj
MAYCRGk3MQzWPukcPSC9Jkhw2nIVJp0JQqs5wSS7cIqf5GbdDnonQjxF8hDgfIE6RDUWa4CrJUhn
vnMsxZW/xHW6VArEV70V9M2YotoTWwQChAZaw0QmmLKhJUKdEEmCvFLfG7SmsmBXYp/Vl19zyi/R
f2snRG2sUyJq8MnzSy+p79o86VMll6h7y9L1QdbRDU5DFsZgVqN5HzIN1+F0Y4dLxpPcmoiwjK0D
F0PqEMQWEioswkxxIinV9WVkxZxm7adJvHRXdY+A1BVU0xuNpb6fQ0M0zzLD8qT2oMJ4EXuJdt1F
2oSaNnKPx2b9cmv+AyznlnQ4zezF/syviQUrbkTMyx945y0v8W28s0qJGIVJgKxLiSKKDf4+0NNB
kyIWrryAGwXiDZNrFFj7jGZbF9rN65vC0naVky30ZQtw57PZs4oWpzx9BACyjlzpBpjgfHgJwYt0
mZh2TOtqsYbOi8lmUHVqY+jh26FERPaYp92jRaX9HtShNyZ8erU03/NUB7qGJIlGfPr571rD0HPL
+H1PSFVHRpdtbpauLR/jX28kjH9hVJUyF8JJG8OhGb4WLWpQbZa2fM5VkJLpEuqywrT7FoUwmYkC
9dVvePSHTqP5xoFwM+zGihKpX2I5LInXMcKPtwzxKSXr/vD/2hqJT2rq4paVHnTIHcT23dY/bWYN
VBMNA2quLEoi0zdWK/+PeYiJ/QG9q1RNX9NyATUrUaR2bk/sEkGTlYh3WwDnI1622UEHDlgEMJtd
HTJKvG7Bn3ijfFR5pOSIUgvK1aI/ScWAFzmpJ6Af1T3FrFYa4vx/iHRpxRZFbKhtYbdYhTVAS75n
cn+2J4G+isR35LT/OMUzWMQicJEPg7U/TH7+dYxZOP1e6IwCbPBZxUR33NYaytHYvjoBxZRwXgKE
si98gHIbtut/W4D/kWW3UiLRJr/Ho+nzH66gZIHj1W18olGpALRL17QfictyGtjNf1k0Uf3xb0qq
0h7pyWsOuTQJc5hntxgUeb36YQNDD229YuhdiHPn2eGYW36XROx+0gOi0+/qD65MCJ+bgGnAOqi0
s4cCB+ZYHoIuDje12aZJq+T2cWCzcihxApyt0zB+MsDl+48VuGYwHpJcenV7hkvJvheW+Lsn37PC
EdQaEmW5ZRGVdoYCRqtHfhBzSBOvtDDp5vevd1F7rrPRqfYGvewt+/8yVRFp4WdKjYXVS3ZSF1QW
hO2vYzcc2zBRa0Bmey2a0Le5fwg9Y1PCLiqOF8yKaFndEPrnBDQFQbudnOyV5HdcvWPK8qhiW0yG
KzxFcwvPiXts8Mmpz6VRE8ZI3a7MdH4cHzB+4WGSd+VUfPv0mU9zk+d7s6m9/0CgZ+TBHC2PX33M
kulL1GJx6zjckD8/UFXInAqSnSDMyPGKNyrkgBpV0VomsAvZEXTvFG1SNkkkX4Xg76iVxFYX3Vee
vxWZ4UdZtNZGvetfOcaOtbx1xJz3XWgXDMNPVSNJoz/RoQgL83CYOoY6tSnH6dm4a22Ui1XofiC+
+1vbrmcW4ImpM/YfC1xYI2ovYeInHV1QMvtiLtAWGX7YJcVDHQ3StRZQfcIRqVuQeeiqQ96otOab
hxqTXVrMTxXaPKLdkzkP85PPmwVxtQlR9u+obG+6iuRgaRMYt/mvyf+l7EUNogutx2R2TcUzZRCD
jA1zOi9INspLQvNKafcQUk+kPhWdPr33DbusglzfhYahLrKuQKDipg7+kK2K6edQzXbEMs3sadlC
v20IMfkUGGEjcTaZnQTz/p/Xg63U6Tj28h3TcfIK+dopObAI/iYQGLwhrmIKQdB2bQqZZhUST7Gg
yXRtchQ0uZfTidrI93VNKxMo9tRcS45z2Ktiph+eYOwDg5BkfOolnys6A/IGC295HGTtr9Ne0EVF
0wfO0412RCmvweX3q+5q8XeG8wIhPWjNmeFsMm1c3aZjzUX+IrLMCJPmlTJcWT8/cWriJujKnqke
olcOj5phQ5ELr1dJrgIUzKjTlV7IP9OxnD+vizcoO9RbKhgQtcYUfDAOpKJOAnUeUSUwB1qIANAy
jhQ0MA8an7/r5bGwqlLAH6ZlVcuP9NsTwbbfPXH2zvnwC/f7W4T2v32m1tkRa+TKaYQZCm69CATJ
DXZz2gM+A6XeaE97a2dFw7hcs8E4k4Z2gVWOQM4PAqFZUMZW44PNAt2CRa7gQlB8yqwSlSBWQ3l9
9nyj4pO79mQJII1JfV/SDtmTkUqnvPeAOAqOmnAjLUd3SEp5eVWG4rmL49XDRrQYufR9KNXpIMY1
h1onZPJoNim3gOq9lp+HukPzdYxKTzOEyVJwJauoyDFM9DNo5ANuv1G5J+8yCcbk5BQVamBTt1XD
c9ciFIuA7vX1bEQAuNqH/EkOy53x1I4Q7Boh0tSpmPFzaUM4Avvi8bVwDnCv0ct4DIIjEorL77Za
hjZ2WPxpUplNWWK09s6ldu/IIaulllFIN5ZaYGCfamNFhWRlDKYMuZfaYdhSyrYEPEtTeD1Ma/As
ME/iktA97YsQZ8jrn/v3Sksh37fEHHmYNi60rqUz6Gk41sIOfYl7IW0w8mYL7B1hN5mJERv/J/MN
NjIU4JiLz+wOoaYLe/JR2Go4mUkjQDIWAegTIUNpbFdLh3ajPIJrfKx7ZT1UvFadeb4ZRt0wvgTS
4sRLyliBZuj/aj8H2B/0eh04sQorNJxjzZtOCabMVSWYkxdLNSRxInR28jQbOloVPR5rMnQzszcV
ZrhqFNiYgeWJs77pq09HXFWGRV8B6suAZfd1vkRSuxkKA4ZsMVqbh6WsAcLYodORyhNjV+8cKG0F
6jv5ZOHLutt2vhg5wB+tDPQ655nvTziIM3XuqlL3hLyB1/S4X7ev+QtB9YJyOqwf8ulq85Kfuqly
t2EqdUfVTLoXIOlsaV2x1VCoJj/PS5+IG0p+WlyQIFoAlKgSAkA8PavNQT8zKUOzDauntRiPyNmr
vS8wYSxrJUw+wCjnriDptyYNQpCSfdIajVBR+vNq71NvaVr2NrbJLE8ilPdvVcTqRihAULrdMc2L
5LlGetUm7l5ieskIAG3Kr0MWB72Zq/i9xDg2D8LxS/CXkIBK5pgTai67sqbAetDA+gIVjxJddV02
k1HypnrCNvh5SFeAMhB2/dumBnx6R8vtD+jLKk1YbMV5G+4zk/r1exflkgyct/dl++Iu2oc2E8XE
OjVkvCBuaK0jmBoi3WRg3VhVGFHe0O5UbJvkIem5dJD6tuwhHZndRUp2fb2a8G0VuiKyGbXtUyWr
0EC9V5PIReeS8Ogu+oAQil450YN858gwycsLJ5F748RCbnYLHTUcYR836xZGfdmjuyd1jlRTU3j4
RoB6UUZD4fPSo4/tvHMfHNEL0UkIvdaxpEHM+3AxmNsSlbLgNNNylMjEr+nykQTzIw/4x6eT/hwg
/quW6JOj7sxWIYz3KpuH6EpuiwqKWS4QKdA1m5TMv+GGuBHpivCFb5UM0fUbTGiWs7A3W0ogGZZb
wJYiVRP1Uioe7XdNAhAuN9Z++6HJ+obU5Ie/joFJ3pgeeVC4Nm0ur3z0RuBuT60dvgKSEcylbgax
gLYxo/J3sHEatNn97ZQ2ohAKKQfCirJ6+UkboLU0+rKqHob0zvobCxWp2Hfp6UFIqESYJDdMwsFk
8slrLZla51KWVyNuL/1o5Hnr/guupbkI24mFxxftvFQnweXqbhv5VTLCddRy8r32S72qLEWg2/Cd
5mQct+mfc5gv7rLIqeuu7JHgo+iJYCYNVLtvKZQtC9kysoV69CPBlvWwzl317IOwCMfNzFMqTQF+
lJSLAxijrg/blrj2qFfW3JiqB6byjDMfsBnM2/O8ChBTO4c+gwvVCj6DpFOP4MNNZblzf+wk55jq
vPa5XZ5mVUn5e63FRfTSTc/OIThE2beJVBb/g4tLVxFBAhv3FnCu0VnFyC7lFTrlK6pJiVjVZyyA
rG4VOjsgRDMA5C4moqOf3RNtNvgFcNvaNisAiYfDTEYL1Zg5nEkGirgng9H/JN80SU9Ozt86K/zc
JqrVPh4bhCpu6/HnsQFZFlXj0KOhpG5IvoMa6ByCfhX3x3T3uHONJfQkdLEUVfXi0EFAwX0GeqtI
+jnpOIPt/JpkbAwbj0NEVJkBSVLH8xANqexVxJnwsDKhXyfXXNkfiUkuczA8tXUulN43q/sMbWhy
1MjK2XD0u+1KmFYhSFSHheJnBx41ODYkkzRdluDsslGQGmLgEbLp/AS/lLdJ5OsnO7XNuqn8eZai
bdT0+xL2WGS+dvG23stlTd5FnSQGRauWVIBwIHGzgikDqQzK2+a0G7KHwKE7+1RPK9ekkQJe3H+2
cRQKgyhK+pavsSEeBIOb33k9N6VnFzfva31DcVBkVCIbC1PJ7TD8NtRPlUBuZkinpXfgjj+hfZFh
OCnen3p1FKQrvRN1IQww1w3TarS8LPGTIN2WayO4u+Y4csywdG99Kj5CWPaHi4X9eIpP2AOxuWh3
gX6RK0HWot7YkdoXjeFsYbJUh5BcAScK7/hWd4mqtVcos7so/3qdRvl/Tcja4cY0zb0O3Faf2Wop
v9okJaEjMoLYUod2FOgIU/CAtnEaOg0raKl0hldjP90aAPuBBBIABIEYB/SB+kc/HjM3hy95ucw/
AAGivt8f64YRkLDBQCtJPayUkxC3sovn1VyqvUhNPqoZU29CU+TcjxJutshk9Cn0XKEFLkfTSjBy
q0JSVc1/bAnoPS3K95gLOAEGUYGlKThjXY88dahheuUOyHrIpc7eu9X+PYQkg4GNnjWC/J9zISfY
zAXo7wjD0WolynR1IjRXxPSskGbWsKj9U9nOx5s6mm5d3cWnGQ/0xlo66/G3s+DD/ipgpyJQXzM0
znj9kYbHzjUviOkOLedIw7t/dkHK/lAQurn0Pxl+wue/cdApfWYlyX8VkX3a5uQ25nv1YqqWqHVa
8CiBmJZEBtR8OX3lfuYCzy3AcQWfIRuc4TgwVU1NH8TGpTe5mTp8vJ8nk5BlpBBiWtvDgfE9NLWI
ClQDE0FZYU0qsr9owaw9d2qP5reFxcJcrjXWyu1Aqa43MDpIyFKBCMzhVQBrkAqCdFRHcq9xWrXq
pMdJ2VWlajbb7N6/9xO1y2TN3NGf7aYMOZuW2JN3nNzXq687ugSQVeOXHUkjkZPUkIiUbArGNRhm
GhlbRQ9yKOiWCPARb1NwaOZOILE+Isp181l7MDqObNbgJxMJvN84h4fwusgA/XlBGQtNdbLkwrOz
6CaX5Sxpt3UKiVyThiq9mA8gUmJmdkxmsJ+TCeL7348FQSXQ1H4fK8uSCT4zuWmQ666W9BSWCgcC
JG8JwyXznMEs2dy4HO8gKBaXd6jtW6d8Y5x2QNE5for3GL2NZJHRFBSCBFNQonwkFCKMCCvN8sDC
aRVmwBvy/DZSH9HHYkA24bUBKLgcTJxk2AbMUnfqj+srZJVXKW+RJdlZf5M6lnKPWJlEEdLM7l2q
kdlXI5pwcBCa20P8FQ0TWlXNa//0iKenYM+2wVP3Nz/QDdDfLI120Zln/wbvzdVIoUAP3phgEzRi
ggwwP70i7cxGQ4/sqRxrrZGDNRDuYBqTyRcJdJEzSoFVv/FrmsScSoDG4IC67AfrtbqF91Oy2JQW
qgWFu/nKC7zaxCrRPTUfaMcNy6O6XUZQ2cCD8tQjrrqbK888YzI15fwM+kZppgMLLoavoU1qOQa9
dDxsSRD3AXVTf9aUdl/UJxfchwP4PXZeDC8E1eVK6rQiMLVzCNOQODmWfnCIYkMwU5MQXG1gt03D
E9pTKAXFTmD9Qs3hq+CAFSvSetQiZbbu6NnOLoIPZ1n/+XWjgIkYw8qYHd6x8lm9TLcY2zhY0VPF
pkMrgHh4E8fDvFP8FjCQETD7RaOvy0lrrUlMRuqdFsNNDcZXYvBmghaXgEAds0RIjckIsvLewzI5
frehaIABGR5McO2igO++m7xzZ6ZpVM6VeE197F4vye6ujIx8O9JNb0yaiX0Cmi+3Q3MGwEnv4NIf
L7vdEHHZbS6byou80ptXzGLBmvbHR8AFLEVYssyelD4UneQhmrPyFBttY2s3uXTVej9U3kRNSu4x
9TtRF4In4wiBIFbIDeGhG01uUAULAFSUnCZ2RH+HHxH09iLZatnTG1vGG2XPc1NTcaCatt3amFaD
yor/spOoT2gb41hselwRJttwSy3YOeI7z3E0NUaj2cH+Gobbhvbr7n1Eyp8lFyYiNx95+CYNWlvz
Ge7zlVwEP1BvQ1SN4gFC34vh6QeEHkKwTs2j8CkS0RrE4dp8+Qvik12J2H9tHdYsy0JC9lKZJTJS
KvvMvNeuwsIKNOt36vNZvLMptug9+pUJkIdilTeD3L1CE3Ftn/orCssAaIVVodW9GBA3P2oMlaWQ
HqpxcDjhYlY29EQLiDecUBbBHSFnVwMcml1i8avU1vfSgpBIHB9uvWVxO1Ak9/9enGAWPp2rBDUQ
J2+m3rQ9VhkU4D1GVeRlSCkEK7V22zNtHr1hW7Lvw8qJfMdtx39hMy+Fuz6SLAud+uBm78c0Ogjs
i2aSBzgcCC2zJmItGZ7hiWSskVpb36S3vnBrqJYBBc+Tln3TtodpVnqleEKUVmG819dapedS8Y96
akIGaEHb33XrT2BSTrzv/BsRSBg/P7Q+3AksGeU1uFYxiwEn8ihJ4wVy5zwx8v8SfKYxvurTFZeO
zCJNiKTUrMo8lwY0gJdpdtMR8UqQavx77ss7+Kh3NIALYqK1gfDOgZW5e/JBOSlzOu6j+5NMawqR
BQcN0+ylZoGhJjb54OKR0tSn6rzlf7CL7H5uZVKBkOyyBPWU/TAnvXdDX1dZA3E0WIR8i6w5rz8h
OvFYGoDyZ5nO0OliQUwCJ4PCyOH7YxOuFgVI1IXmMyO/uTvG2lZm8/L9HGb4Ppbd6/FYIfhGTU2w
UqFOj+esILxCFQhW7/pZ35p6GFnqcvdA3tBfOx1RqHsD5YyCeEDOsGept5P90ftKbVYPEv7whRmo
NyEFZjPY5dZms+ME6qDnLmrNn3H48m9h3eaO6Es78pcE88ScqEHJiLvLSrYq5GvKevy5RDy9PHEc
yFvzMgc3+XaD7q5FYGp3ZKjtnBiLFOhN3+Iok9uRgYx+O+UD3jcicdDL8Q1NPaBVcnXjpEfg5msX
K0zBiK/z8/gsEIxX4awAxdGX74V3GhFCiotpZuuJhENTr7Py2jUVqUAfYVXq8EAN37xC6D+qainN
MERljZHpqAKOOrCPECq61rd7h+wFxd0UGh8vuyaQH5rCwyd5PDE4yJU1Nkq+BOs7Fj6qYaQPSxzf
UrDDeZboLWj7wuuxWpXT8GGqR+xQAlHQ5BZbMandq+98Ss7sLDjzs3blyD3Z4Bhw+cbCw9Ib/noE
UP7MEwgp6m+drQe+XtYNPZsCCOR79hQxXTqGRkcED68j5OciWynOAxJM01ZYYDDGBydhWt1u5Xtk
XlmmIsmDFfeyZCcZHqd+WN+33qa5+uF1OBoHfdCH4i91Zir8hUx4u3a0maQ5TburIJypLAE+MJHf
nBgqNcpZr3fK+oL4NP4yd6iDla5s9BUjgkSj1zt2JfZqwfX3Vrr3mX2aJTnhp6mPipb9+YJF/Heu
yCQ4lzMj3bvFu3NboKVuXAvBtrWqcuSC+k7u+1B7gxTBeaCwTGmvZ7TFjRxje4qg3Im4ZqakYRkI
wBCLYBafvQ1r9c/Exns5BpIlrP4PYxdWtXD6DSNTOS1c6sCKA0xOlCL7a7yvGHVPYy5BsKelx0t6
wO+QyLhnmSORPjD+pZmtn4LPaK0HQd7nbf31fpFPPixVQ1du/sJygQv7z6kZVmb29JUvUueRNo2g
HwmmutmEICAYCUYCqUr9Z6tR5Boi2j/t67xSICAnazm4QQSc2t3ogkJxQEGuGmuoBkgRPNsOA9hQ
GhIAml7ZnGqRVgelBFOSq81/FyMLl4c24IH2iFrJ+MKeX7/4dUWNjzYqFgFmtNlLqN75Mke68uVs
pqBAqdgX8Dgi7BvNZ+V978yjoiKYfiotIg900555XML2rrB9AibCei4Dw5jCbg9fldMjsM8eblts
+IBCoTlTgyRJ5IFuCehjvpkN6x3FszW0Ywg4s4+cp4edOQ33bwzS6JvHidBgcS4F/PQhBEdWwRDT
gBAhgOw7XPyCQo1hXDrOWf5gPRLBtECyWuffWYGcRcsmXULTjLRP2eAMnsKjvzBuirJIczxpLP3K
+asoCG9YsnPGTcKXyHwKRwbq9jYcWkj4vGl4qC/Y5kDSELZyGbaQe6NkDF7HtMX0UEgGlYlGvPGo
1PxUrSbqKS5spgaQKD3PGeCXmP9BU7nvenwrGoFo/9CSW4QvphdumNs3GpAKqAps6oSp+gpkycJW
Kw+L5wn7SjkcXrOytm87pwkCbwhmJdrOYU5E1lnQkHpQvX7Q1OdDxOwX178jjr2yi7i4Tl7SxkzU
jdNS7BkQ+8r15zPtZ2XjVuIP2oZiQi+CvGkdMaX7KOh09Lz+tr60bdluKxIhmw4C6HLgx4qrKLFF
2zBB61rDvt30PGiAvEx5XO2PSjSkno/pP9QWCkWFYCJFUZDLXW9gcwoXN8R8J1jKtOOGZTLXYy+M
vdto7Q6fj4Svnp+N2ojEQFEt9YhCz7MyQiulToqH7wCgO1Fyfl6aNuhvhv5v8mciyAEENr/VTye0
u4iFeu2NxWJsLG7KQ2Cni/tg90QyxHhgLSkD3vgbXlMMaoz1fmvHK0U4Y82X+wS6bUdkhFRB8bPl
6SQePVMTBTT332pCR/4ZeOxlJdodAfW6Vx6ZwlPapctz8WF9N22lSQda9qLakpyicSIxAB85FAE5
aqBC/ha7BFXViduF0Hk3h19RGQ4T/MyYXOaZnN2RkB7eVpNxPXrQu1y17rOPvWeho1WNuN4uKjf+
Ujghn3Ah/Ljzpr6rj4FopXaIp4Pn+RG9klrUJajmRckRyzcpxm8MLYjTSbeZeremUzNR9wvceBX2
21Se9svlPbQl9RNRTdU+fK67gpdOK/zw3F4HePphh0Uxl+r6ZYw4s2i2/kIxys8RTB0/GdDOPS12
E8jgJAdoe+g2Ew2/Ntpqdi30M5BkO8XRO7Pqu7tiSyzsGzyPUu9rwy19a/ZLuCE9wEWXkkuLls4Y
Ip8hd/iDiLRcDu66Td8IWE+XWEy4Hokg5GRJWtG+V7ytR7Z5SdPxXFDekdYyW2YcCRmstxR8umbR
itFGCRNXK1UxzQNqPK3gaoqvGRuGow4dSyqaUJf9trycoYG1zh5fS1O/iUGmykZlr1JXRE8RWZxt
+7cU43kQ7Vyy5g0RJN/hibiOVV0siP+vrJLQQg9WW1VJHeLhwAUzTCaZRf+T2Ch8/mP4ZZBH/Hjt
MqLq5cc/J6rf3KWB5P1qJA9Om7GXAGCp+dbRtnlb5OBxW1TeVRmrG/l1XxX+a7b0RgQVRNI7TYWC
Oks/wpZHeO57rxNfaUTRBBFB+rVmqmrpA8F4OSuSY/Ai5dOTRK0a0C1GMSQvcSOXfZupYa+RyzO/
ldAZBuby40vxSlZcoSIBox1IC3FaU9LAk1mCMo2xH/vMqMBg+mXfYIiV4AaI4NdvytxXULE37uoE
D/ajBaRkuATnqtQT2lKKpzVYjsT9gCWxi/zmgDUlRiYLlLsvSuF+WhBtRGGoa+0TqnrXZglZ45mf
WpE1mTTgQv3kUQS1+2QwnF+63+/Uamb2XdW0kfHnNPQ3DUqI/8+AJeAGQsxlqv356YS5eqxwcNMF
L6CFpWIW/yyyqy9KfK38x0p0NO3qZLyUmukmxQ8sDqgfJWT2yAa0qMqv5c9gt9qAsHctq16CT3T0
crZnz7UW/MbcGVVNSO2sfzkgL6COb5100GTAUbnAnUxFXk7mYFkhjH7jEk4di+kYQRTzDgWT0cIP
V0mvP7Lc9y0ZyqxNHdPRLps+aWqAJZ0qrR357VJY8Q7UPLVd5pNIolU7TWrR5rFFRk+WInDQ94E0
xcctbzV8izjwkKLlAd0V2wUyjHfmTaM6a4+CRZBf/U+tAP6BH7UVwyZoqhfQCtiocFOTNZJrOB0Y
eoHfSn5KTKoHCNBHqXEXbXJlW4eYQVJJFbaRi6Y9ea9TmyJvNQ0lkOLMsAIaf6es6js8OsjFmoS5
EiNIq1pPLKWylUOxwirFzrajrTqQ8/GIRKIIwme21V1AtSZYxEzpmzcOk+zzC6kNEJc8z/HwLpdY
7At9KFt/YtbYWl/ZmGkMS/bK14GHnG4xwp6FMUGah/xLTsftr/HLgWrOagqEjgdfemOZy3a4n5Jt
et4YZOnoTp2JPdq2zPYU4XDpPWYG+MFSDqVm5quBxCDld2hO/efuoes9TzYbu+E79s9u+AKxyqzI
MC7kVU0n/uajk3ay2GWyQg77c0oKxrRP/EwxViEVr9eyRSNI4TEgimC0XsnkjFZKBpssKIWFuB+E
bZB0G6oOKF7kmWkEyvUeHueeubEV1+6PElsnsiXwvaMC9WqOsczbRjm0xRjpL3Rd0JDlQSnXP8Fg
zhGQiTusyTsh7FtpmYPGN/EL5gxQbfVncEPxQOxWOsqDaTS6INggXRNwsKITbT5dSGsA3xxT0b4h
l7UrG3gbHOxlFmSDWCCZW6cBTF/iYPUXM4K3keS+fGeY46nv0UERopuv9ewbHz6AhQTPqoKe7l6z
niiSZFRk3LmrVNhcnqD8pSFqOthQc5z8QuEpiLfbVbFVbLcai+/k9b22YB9WSb2UYVUgLX6NlP0k
KLmTQKCpSDsxf8tDdK8jIb1eAFjwDglVODq9oklWdyqrNCbJwj8jHif5znLkOkCjP4acTGzPzA8S
vbvNe3K9fuA6DK8cWUxqp54gwng+cNZxJdG2oUQi26DKUnhCYq0u0Klpa3TQQb9D5YQfSkWkFQf/
j1Hdb/ZduWvrnYC2JmrFgVlIefOtsWKOubuTJz3+6qPlBf6f80DsHr6zm3yKj9Ir3cW84w8tNkld
9c+o/WwLEHCpKPfM+djgmgko7DP54FpuhYvL+bpvuG+rWY6kUG5bjEG8PLXJrhkt83hgjyacZpki
veu5cCKUfc2VImMK0+P7g4XGzh1mjO0MEjFAM1eq3ACQF+FchB6hiruO0q0g1oE1l3UVzhCO8CIY
cAd+BpNbbhsMAA7GURW+g/cytPOo9XWZXMdbX9k5/JQRMgAprt2ScTurGok2S/BDQea9wjbl36AT
OmkHj18jB8dP4BG2R3Nsrnh3e+DJ9F7TozQtKqFzGLW7lCLpizXZmzhIVpUTnynnN2k1FTybPGAI
8NZRk8mmDwIabchDvlPMQPI5njQMuVcCDfwH41wu2i0DN3I+AHk6ntyUGnLP32ffQCYw58cl6x2G
pWR/qrN7gjCslDygS87e/b4e0xCmHH67eJz0yyuZXSqHQQqai11JBNOeloUyzwvU/1Ro6i6ktkNk
Vm2tgfCPgf3hnMaqPL68wrJZIcrUslCxKuJzkUYyOyZwx0ogRjWbfTy2LWX+5LjdnIUrqrDSa/lv
edv5oveGgHh0cgxO28LIYgvs/geWChzg9PYuVJYKMe5ULH2ING4L0yos0QH+MQIxc2Px8kRVPkc2
FTtZJ+hNzY5t06T3RxKiYVVwB6vx7SkjVKlMv668ZsVXvghyGWP7m11DtNY8maOppSVIU5ieTnOm
c4E2i8iDCEXd2KCaVxAcsJ09P1DAeSBkdOSZyHosX78tfQDk0PGlMZ7OFLNMPbti6YWANYrzBgJO
j4pAo74vAEeiBCU77CVkdqsJpV3PD8q7wBRfyoNtEUOslJ6xMITddfzPqtZ667+ijtFlIPhRkL2C
EVOAZjG559t1OZBAROSf3N/SS7TQFEkyrdpQnhcSl2lAkXlkDOAmOS93h17NB5SDUF3iXqAUW+aj
GwFcWxmVuC5dqK+tBLI1T/KtAGQirj9TWi4IKP8tQKs7ALJoAhxaJ3gp4aPDhwZP0lUxrOZMclbF
pZDuIiOmtqX3ZF3etayvQ5Z7+qOqjMsX/zeR+wwIDaE1r+H+rhmQygIg8rP0ZRTitDWIwKWJg8Q/
DQjj9v8XFuRDC9U66JOCW8bjkptSJbCLNcIc/BstIUa5odU2fsArf+P5TzfTZaLUEvfhDFMyOiKz
0Q+dHsuWEdVXprFHJezrHaJnt415LSsz9p/JMMkUE2w4cgbpTD7p2v+qf2h2NvaazrMIonNYm8S6
mwKVXPtuxWA7tXHrVP9OuZQe7oeXWyOZ+6XgcY7P9ijqywjiSTlkI7DCEGlvPz5fu2TG+AHXJjC8
A8FH7ldM1lbhzxbXnLljn+RS7gPXoum9Euizp4FJxwTqBgU7Dmd2ioQr2D2Oi5TpPsUPaokUGjqA
1m9QSHuo6bHAkw65bOPgVSwfo9o+jbSC7DkbGestV2mrxs7ZDqnXX6ZObW++Bp4KSJtFEE30dfCh
8bbOVToovT+5ctM1qK8qxu5XuYRWVvR4zoruylUX4Dc3VbvjpmMJP01hjZjttezcCeiz1LQkfnUd
R4EpHTn7NGpOpDN6arDB323s6Ps7w8sFqLU6uuwxzoa9TBQMI0aXqJQLkE6WazZObjqXNr1nMCoS
tqjZwc3dIv30IRCf4s2ZtGTYQv+hFV7Bm7h2hk//yx6F5x5Y5uvG7TGUagztzCVjm1jHFOFJAO6C
Pv1qDth9ThRvnR+/ZYBeEA4teZGemHJnHGBJL6bundqUn8Hgs5MQXIBMg72In2d91YN25uNg+W2y
GYq6gaP/r7OYPUvhwlK2M7ZnhvP3+SNet4eCNHqRhC0l6BSD73KR6ZpNeN9nrqzsraKSf2DfkUnP
N+SeVkGCWzaZYqhHKS3JmTE0hpT8jbmFmSJCp87KPJvfDsk9lLS8/jxPlTkd+MkXOL2AQpvlwhOb
8ZD8VM3PSdlsB+OaO+d74vo8ZypaTqDJHH6AGyFMTsxk1yDtck/z52D2UHaZhJRwuLVRTQmbpWqR
qXTgJlu31N9bs/R1bLX684oYVUYZZwK5u+rw+C/yJLCObdQf05B18ZlJORzQqsDd5LaiGzzSaI8g
HT7KqPm2KLk8TLD6Q0s0COe1aIZCdPsyyaJZ36z9Ia+28XHLBGwirTsZ30gN/PtYcqbBH49kpj3m
L4rexrZwvrImRqf5PPAsw3IvFref0gPK9vlqmAAZhjcVwKwnFiURxA2Nua7mHPr6aa2FG88rBcSo
yELWUgjRo4GVw6AkKIQbX5b9wPaXu/wqHeBhliV/4DZyjbd+EUsmQ1toUXXr/LH8goRJwVhfR06R
BJr2OFIR45nFxg+UBVWptWV+sB/Defm579brS+qLopgnoGbQTw+Bq4drjYSRCIcgQ3kOlkLS1BsX
W5WH0mXUFAUsGmCfbB4lnWWb66HJ75iSq+S3LmMSD3XlUxbLdpLmA4Qe7al5nDDwNBikNXaU4F8u
RQd0Am0dUgBlkaTH4f4QyVQr2BU+0xl2twVgqi4iNUSzYDqJ8IrsxEpYj1fNwJ2SYGChzNRWpxDY
suiJJxDPCCCNPeAZeV3d2qbsZ5xVwrr47K44Dnw9F7GB7xvy0YUtIfanQjzRCL6zZLa6UEcs/nsn
Jv0CEOCHE2Wv3CyUB5v3O4sbbAha6lNc5rQvP3diwGFSbZV+jR9la+rRI1rbF2F7Ezv81ndoKQEQ
yn+zFElJyVu2RmTMn1gpD3jrRcxAL7DUaYuDoZXMNqAXMRnFlkITmdumrsPwi2zYNAG79PSZKTTC
myS+V16ssaJrDZKc+HDFqZ50yeEmp3WwcYLUgOQbO43ALBy1vQ2d3apvsYAqUA29zq9q2VswC7hv
SE2GrwGorcwBduES8pR84grtmajQU3FGkRFdgoXJdg/6BvX+kFPPglqDzJ9L4pfx7Q1Czfs7tXL+
EHu+6UhB+euIx9I2Qg7mQZNeYVt/FdU0r9+f9mUPQ5l7MRclNr/tchd2GyACKKAoR+XjFMUcKEZY
nlhRvn+d/o1TDCFFZ1yh5enqPCLeDvlTutTLEmKLrpYGxszNiKA2u4uR7t4Xbjh+gwGfQ6oIEFWK
wf7qKVB1TfmLD/9IXjvU3DkZ1aYWieNPnC6+LnzQfw8nW1BWxgSRguDZhgpHkvuBithRmFU75TC9
RaLVOIALIq+oES127OOR1kVBALy0Rk7fCmrrHyyA5srRKsS2MIlk63Y51oafduLL4befBYJmCIaG
gO5FCEv4jPxHTtX46do0QhvaDnNJgXeGqMefL3/GVVLjUkdeOdqP5F0aVtApeovoQum2iXBE2ktH
5tOGdk9nfVcsLuHWT0lOlx8oOy1gmYZYpXXmOPU5dhctUAWkdc666UyYa58Cra09cZy1gcNkDUAQ
bO/i/QnyqY15hxZsoWanNJUoCRPxJbMCwWnaecopI4AiVNbsNc80GL+WK64YxTOw7aMCa7ZlzzN4
9t2U6p2BjIKmm16HlTsqwCa9gyp2Y4/dEsle96ZdAYAs+HgLPdu9/xiv35fNwntnJUjYHELJe8KS
3CY+xvLc1kZspWGYzKlvn8arKZp+gqmc3WfNhwHteJ3MpRATVs0LMSeTzbUKCfgb2HSvAaaUyO4T
rOYKZa8e3vkuJCO7/ZRsyt1c1gt9dGkijyojdc3Z7Q8t6Wtn6+viDkKaDSwbJYijLcyEFKvJ8eGZ
B5cDrGAhIUBsKJgvz0xHmd4T8EW0qCMSuEJBiU2Mlf6m16X9/zZA/8FOPB5Z1QMjLkk2g07akNg3
PSG/wg+ALAjiFG0O9Qq5xk36vVxOfgL0v2Hj8oWqjsM9wtFx5GHtXhuy9OHTdWPidUKYY7XOCP3X
y69ZV0xmFF5dd1OeVUvyW4m3StIb5AwKVTkjN9tI6olkT7Jekrx4jY4WP6XKrxXgusVLMwBIo7it
QkZi1aKwXTV4AChUBpOzU9xHzepMmhLI9r8qQ6CoPNP5nmuJR0dQYLNySWyr9txd/ttB359jwNf4
PKjMRZGFUYxo3zGBsD/1Cs7ePAP8O00MrljvXMPjoWqQQ2LjS8JqXJkHUdP6LJxybNCyjBtsVadX
sje+F/VJyf4wsnQBKhumAtOvdQS+HGVnDH1CzJSEEk77Ootkh4VrZ74j+e7b1r3pDJVOuLBwXXz6
NMiUDldmq7Mr700a5wuTWPYff7mHKk5OyG6SvLk6kGPxycjXibl35UIHgnrdhwS/Rlzew3bs9Knx
g25f2dOZsozTnnYRqxdgy+C/M6WoaTp3kUF/yGdfs/k52uQe3TUMSroKXNA3H/+e0gQIsn0049bf
E249EGvctUrI7vGd34yfEMwB2LNmUTfJGQq4dM2tpS+v5oR63rLuMtDr4+8mp5VSZ7wC2ly8l8pB
YNfP8gqqRB/mlzLNhU5+t9HP53ZSRhFH6hPFQic1nZhlK8vhT1fCoL1qBPmuWi371QfuYOVeYosd
mmeh7sDavp0T1zetDnKRLL0WxfF0zDMLbuZEU7+hsOnHGznQInd54orISc2jX+MdBUF7IKfgttcl
tFq/9sYKHePfyMG0NJ755/meuPKWyXRFLSM/acxuJwuE1C+WikQyDLpMua7VaSBW059fGwCfBkBH
PrzpLfwbm/JD8VnKcoOR4yTtAYdZoFCGkXnWwD4h3p2oy1lXJ4alGAJdq825v9TCOlxs4CXNo6Vz
8WbsBPsvTBhTdFO+6MSqI3DeG038nrmjJTtjrxTr3VGTemzOLa0RQ1A2vmI77n9sHoo/0NHJqGxL
7OJ4wtT6pd3x+wjveZZI/U7RXaJYtXs+N2zRm1Y/+Y4GTf/ka+sYTutOdKL6pkOMye6KmYJpjn1t
ZPUjwK2zdI7YcMjSP2UCiwUS2bD0Hln3D2D4Tbt5cScdsrL1g5Z8Uq87mBBW3lLDJVbZh96463Az
71IwQ5ThUiqxTL6QiGFoxj05vYRaWVaZtgmrq58NWQQGeJ/BQAVwN8LdsPQgA8W+4cYN4AZ3gHBv
zaqkp7jCnyPFe/uPOMu2u8cQ8AK3fl7llCTqdAU3wBltO8UY6FeljO7+gywB6evDIfJfxIHKPTxY
dTf77H7lM/GktbGeLekq9SYKLg0H/aJh8BEREX1FjYdwrtLTWsU1WntFxc8rnbAleysgA2q2Jfi6
JOLwxOmOHmfwykWMoLHuNBfXXPqPC3w2o87nKCYq2vAKeN+NwmP/5Epim2vPPVYJ7BlnALLovr4b
Zshs4JEu1zVZRLS4jbrQ9cL4XM1NZepf11/BBTszZ3leo7meWDvfDyFkkjdV3eVpic3iDl0n6ruC
NXOxGiGQ6HVvyMUEhQLxUaZsSGFlg+1kWIxAhB4/AvC4ckZha9t4/eV3AqQFuA8+FP5gjvI/Oj21
YOtd+UkBD8Ic6TkEzvoff0iGJfN02Xrle/U31BYFhaty4ppA3baUvKNo4TtVqLo+On8pcSGb6nD8
qruAze2clB11B9Wmd9iiLCeaVAagiv7Vjoh0Xgmoin6ncJ8MDoL4SJ/ss9VagJ8ZZi5EXXnKVurn
aUQK3WJAyKHAykVBf0PGpr7FgqTQY/1AxCjs+snwnF8f5kYoLU37Qi96YLDJIPF11I/pag3w4zWo
jXdFGJPnhrUdnxSKdgnUhAO3jLZLE3zCt4rVmec9RoCtdyB0xHoLjyqyRUDB3EQw4BDZRZSZvSMb
rnEMUs9Ux/aDFVlmUTD2HYaIlP2tAf6RSa5N7xYF7pmOqnx4qDIC7XvJUsShLKLE5pIO7ao5Qvep
IA5NqyTCSovD0eicJRM3eSbLe8L0UyMUzNyNeBhJoRKV+qcb4aAIVCPrIdAnPU3rmHmvR2lQTzDm
8jzakbEmG0v5ep//IouR7pzfqMoENbghVPc4a6bUm4+alwZRqGgFwosPLwdNPbKzLD4ZYi0e/CUi
8qsD86npOQjpSXiLDxtQ1grh8mLgCB8M6vtQpr4wqvPVZ7r4BJfAKwTCD/cX0A9Mtuvdo5KXGsnh
i/XlHmexw69M8fBeBYSvbx3Bof1BsMgkPBperhsYBK+nRtjtLRtjLZ20lyzZcbMw+alt8BuiFhHF
YmeiJ1Zb84rk2ztQ9h7sKd0NyQZZkNBRl44MIIfjdkeBzJKL/oFP7WUkcl+JmO0cAJ2xqUn2cM4r
CLl0fFzR3ElnF3+cBxDFUlaKYDm04Xow42BQH/wZbtapJnHcgztOcUwQRk+oQIGgGzkckuJJy/Er
4XdN3f1OmCONzkrZZRNL8Cl+dCrj1CLCYTsMWJlyTxbej1fYR+BnmAonxGpHS381GUteYmFuKBQh
s/pol/+TEEK7MO/mMk4TiecVawMbns7EPyjsEWQrfFdtUsNMhq9WQjQ53DiXBOqQuPECzTmfkj19
LDesqBCn53Su30tZMvVD9TCiZKd1sJGGw1jlkTZSqCLod6py3H/48dAvbweLxhHutzMYheRpTjGO
5YatXiIb9UjjTt7BuXOS4cM4DoiZX/XNN9BcIiHx0GWR2Q85XiM/AQRNw/NRZy0bFSqED91o0req
8Na086SeqYZKtIYOMcJrXIemj/CVo6SnujtKo9Dq3MpDb4i6MpJthYp9WPqVBjtDxVUzS7R+lDRK
jk497gLc9DhnPyCnIaeRgY7EXSfHBXpvTWNI6UxsXpKJT4j9gCCCtyrXDrFiI/nTZoVrDY96KIIR
+m6a4uD44E4I++kWG3O6GCOxc6P+hItdW1RxbFNkBc2zdxB2XaJGQENJS+ijCtk0yt0PhjT9onGv
rUaikl4j+6ujhY66IBzpF9vxvs7R0XVfJwYzARK5Z3eU8FhiTcJfuGxissl86fPtO0s8rQBaNowK
m61lTaER66fAkKN01bP3dFbZTDqjp4lVgS9ezdNydfFzOMI0Q4SawupCqnrpTLlopktuEIbLNLOi
5Ci2Blv7NHaJ9HhY+ZYS4VZzsYan2r2c7agnerJH1da4z16gEEh77iuzDzD2VZi94gjl8vWcOygv
vPHv27un9OfLgWP/Yt3RZ4EsKPRJoZReAIvovsSvEMexeN80s9Y/meJgcqDRpq/6frziXI+1vukG
cEGmkBYXr9Gkgq08K+EmDw6IGrLee2RSH9vrwBulfQTqgHMKXrgxIjyTy4BBzJddes2ATE8gXNz0
bz9Hr133phGsgtFm+pJ7lfq2ah+UFk5RGfuLYn20TwtI+UGwRE66fKxD0Iml1/skY5CbJPgdcaX2
RYsqixOpSAFudo5pARmNdS9/Z5fOtksUwCzaQTehN4ZvsaeiM9b/9dUp+xF+m1fmxtaD5f/aNuu9
yCZ1moaVUk+IoZEH5kvoLMaAMxvYWF5eeG9fhZCTN9TaHBzh+x05STefkSyri5Fx5CreOlwDYB91
Ottzo7JF6HNRbgK3RUQcr8ZJ0V37bQTrWJUKtGQYHRmIItNCsqrD9VFfpQnO6Jgr+hsnxOI6obfe
O/4bYZA+l5CiOCEp2wnHtMh4KDCeWsKItq1tsYv62yDib2Bmj26RaxRiWt5C0exFOsyLm/lmaVk/
Kbyv2Gqt8dxttRkyYkcjswzYZGPNxIlF1Y0vh51mLMvJD/A+mP4WU7/3YxAPFBpGTQEtbGwksAE5
f8ZZU/YpkQ6giUnH3KHETXqNkyH9kkWwwo9nGiZY/qyJaR3D3W0neMslEOyOQey3IL5hRVjO88Oo
xUpG/b8ukyAW9/Ao9/bNU+y5r/8XclhUjzyUhgG6SiUjH9j5MiDpPt/HJjtMG9G69eBWkNKUNj8W
daSqwZPhbK9z1jHjQ6LpdsVCvgfx9GOBuSs0rwI7IgGOkOwhqy9koHv+iYQMQorB5EEOQl9SofA1
bKtS2mFuVgCc9FK/nC9qEB42qMV1mTYvPBfsub7PEm4mdCMEBNmU8mf7JEdQzT7ojWkfMuslVCih
eBd4MZKgGAcwVb/6TOQr5IJfBMhsX7x/cWwmINFemRzjSPIKpDKH9vAHbsgGsHn3TxiXrEGy7jwf
JNr764GWRNX3OMmZwxHnx7XbG85TVBpBHPJnJCQtqZ7rp+qvChvROU7poDTZTFBXBKHlt7jyqJAp
bgZFaTKHROVsZym11NwSl8e1UJks3+g98xnBzh7zZLZ09V7miPxANCDTGAKwI5Wi3qZYT+4m+MFb
TLHMQigKdxR4987q47UGdTYAhVi6D/SaozY+7iTpR9b0GHGGsfgB/7VUnu3yj6NMtlqA+hmXwZBO
IvtRdJpTe7I6rraZbP2Vcv6Xd+XPrpv8P4Pj+K40GeW/16mk/k/JMr0slFQZPNloFOqHCLskEWpr
eJhqEDUtH/y7DgksEpHFdNdnM4BOS2nHAlj4CUocRmFZECRYpIF+ew8nczpVbzDNzqQFLOpBZkTn
MlRFmvYeG8ZiB55h9tTPF3kxrYmL3eSgLvAAK0JWT9pucEY7Yu+V3r2mDSzNKfKPmnezyHin+0YK
ay4QEEZoHNtZ/j3tNn1VeHg+QWjhjkR5tLy/9UlMzQ0T0Mu8BgjAHD6fxUwT6rmFZTZG0C2tDgHC
xIkUJzePovMVv/D62/zCLzjz5cjys4GtemtVxPyq8pPd9iDJjm5Wqj7PB7QBEqZvpGL+anpEaBdU
71FDPl0st7YzQwonbS1S6h2AOV8qhwZIkY5sWEyCoV1HfGFXcH6qeI8sgLryCeOOdhuer7S4/c8O
z3Ll7MxkEPRC4/pHvGwl9xLXnJa4zLbD6ubgkKNSYbfq43gaJfcq/WINXlAu+CYe3pzvVEwc5TD7
ocbgj6h6CrGZ2jpjr0JiTc9SnDsIADIxLa5wty+KD0gHGdj/5fxbJd+jurWDzJS2Dl4yWJnmxcH+
InWEaju8N4EFXFjJoWw5YaNn5HRxmBhbS1kSXHmMm4bKuswmrycrgniP9UWqcdYtRstJRjK0L3Yi
sz5vQpcBznMbSaTUGHfJsS9jJTG+E1c8Zw7FsGjGfdhjNYJ4xL+WoM2YG2lDkuNquX1kEfk1yHWH
Bs03ql2ZSIfxR+34X7VpDrrCUh3ATjKj8i+fO7Ihe/FlhH0FCWgx4kjW0OZLtEEA5/3/Z+sip2PR
820ZInUulCP9n9Yl3rTDLGpPn8BVNQb/hbMv5rOoSI0fxA52WRJbpsJztDgP7wQOKDtEx+IpTn6q
BGMrHUdMFhkuRL1wD0udwiKtaaBUZt2sIds/FIJAn4676WNGkqtMJtgeJogHTvapw0J7UoGiZDVS
X5tTks+CDaBp7OligWsH8fGlPFQ+AGIpF/YEvCfMNsrn8GWzoftu9CKQTrdKKvAo5gzEF49n9ufr
acuiKNpLrDJbAwzitNv1+/4aNod2xrd18w7WWJfJQwqGDj4+e2lF09IO6iDTEc1dBSUsSXtFePjV
rYLC6sYGv8z5NgWZv9iSDHPH42z4WBMb5QlvShaJacM48zlHQgpl4wcjHDKHb4CCFup1TDsKuRVr
ljWo4ftcazVtRFZadw4F6wErAFA+KhkaajBVRUC5l4CKYjxC9vLZQ7/ml0jFAKYhCHQqGvB05tDR
9cMkwXfwNlPUbIHvi1kkMGQ60beDVVs1Rj7uVeGo5pG5v8Lv0ApdGHoJ3iJA8G1VC8uI3XGGojGH
rPEtzJH5IjH1DNh8zRNz9TsQoY4boSfF7oXfp46/QkCv9DmjQTyQxijjEkkdH/MzllQlD36Ttm/f
TGY//REcWEdHvslQ5yUQXxrqTJDdzfHqnFOcwI51hLRe2373JgiW2UFsLVRK03scArZiquQRXa46
yEO9brkXNlPCfRik+HUtyDuQrN1OcyZ4cOPZjYGqmWxXmljl3XWwtb4EOmVU7tuETfZ1Pe3s8ocq
FzUKOUoETbleptW22Yit7AgOCbDvIrcoEqQjDlC2/gB55+mqMEx6DiqPetTmW3srtWrtvSk8bXQS
vWJtzrwJK8hqXe1SHPZClhmcL9stqtS4qA4w0Ftueqeu8F8iFbjoKN/aUWgmEt+VeAPkcVDFCZBJ
JLj88OhlhG5XmxAnbgM7L2kbWVV23fyro6Wytm5/1N1SUwLKFC/+KazsbRIEVhn8zgzJhWxCLKfn
AjCKzMv1amVJpSzN3lRnzvndVoe09vvfm2mVBaQnytNKP3zCXILittO4kXKZeEF7mwRsJVSNvxoN
6Y9hPtwm0ZJ8OVpLHTxDM68bqRZbLTHSZJPs/bFNLvYfsik11+okWZbJOxZUBGL4IUgw3Ju8Dvuo
94FBaI6EQk4xnUX3Sw3gT5tR1FhTGZhB8EkXQVnsHlFV6gXAg64+hntDq3gYaGNloqKHkUbq7JMK
6ny2GsvrwbvhkUQpd8Ggw66skK4MfUVp0FtUTPYP/OFV707HzA0CaohbLMP5sJxlWacxeZ72E4wq
ZrZCOXMsAWPBs7RAX5q6y3OHVu6VIV5mnzlGxi4YrBIX5bonyuwSBGYkiX5PqFbUi/DZxnV0fRd5
cGf/kcaxZW3QLNq4MWpySTpX/aiJegaDnD6x2o/C2uEWbKo2g+VJgXX4evAiRd6WkNAyJt5S4DvL
S6J8bWD48b4ANOj4BjKg0TTgjUIjjcAY4clr06UtMHYXs0TxgJSplvI/QpTEtgIf/NH1+6euWMJ1
3c4Es9q8KkwSvn6NwCv41P8HsWu+FKPFycawoO1gDFf595TdvUeodJJxGzhK8on6xpdM076MloRe
xYVQipDqFawYdsyYHhp2aUKRM1la/q0L+PnpVQWFwlL4UCFRthjNqwt19E2uQFSWVZ5QJa1eMaSd
teP/7gNtQlJsng4EhS8KFeu690wzUoD3QCQPPLrJaOA8xwBJeE6rHASS3j8m1fdqV8V1y04KvVS6
W6zXvAylGkjv/KJQXuinMt1JRMTM9VtjvrXqb6Eml0ehhCOhZ5gbfOKZE8Fxa6Pqd6MSryb3cFBa
mDE3Meyu1XpnCIcVLMM5PfvHhcGc958y/R9BKptShOMOp5w9nCtA/6vIdawnGPGsRdiSw5EjWsMP
wVzDR0AgzqYiTjuW6+zp0mulgbiGFLpJXuUxNX32TxGtlFiCKbU71kk/1XELWDxv7GbQTHujIbJi
iqThT+9+Gjzn/+6ZhzSXLKQM2F2Fe1hqI/XaeFpDA56BUVoXMtwoOVCavoH+ca4vte/F2mDg/6OG
+mjzdjxiDi8P19QyyA3kdEcBZc2XzctctHz6Fj53uass5SbYeSKDGW9GcXz0nK94ptusKNoArroL
lESBFwWrowIVYNqQiz5lNwa2U5W7lcxtwHNfC44u9SOWgvCrsPMFiNa9nWMknriRtrER7zB3rw+C
jFLKfKcOESrqRWEPFJUjtWD6SsKYd0utQRixOHVKQo5t3ROyZzrb/lPvMpZZ2AuqdMKIioQxpvW8
KE4TwkwD6Ep9VqIv77POZ8R2DF1SdrWOdp3HrdLsg/U7O/p4JFfbUFj9DMVERQbDltPGNoTLpAgi
psN9K07HnHuj0pHjBZtN2Ws0ZbKSnILCKCw9tLZotSCHFtkLiePyRMqGyponwfL0XHjqsm1l1Rsj
5MmLYLe3YrpYy3DFmIIa4Z5m9KypYpEjqly+POJzJ/t4dcTN2diGfrLfmnPKNf0i9y1gv3EHavo/
MmLBpf6d1bcnPBD0m6K3pJmhQKIPm5uXX2JY6bmIqtzr+zU7wEep+6Sd/y/BeqA9r+kR4vVJtvIE
W+yDpw2Y7h8ogfPYrsPrdXYWuPNOgx7SY+fjpyBQ4m+cJfcfeE4fdMoueUIiBK2mIosWXM2LATGS
lSERiZeWwMq2CUPGzEszu8MrkePuQrf7r6SNZRaBaNT3fC7ibcksy8/wrrv+wuPzQxvYOijeXynf
q11GcTVJ4mrx7jJe0ePXSHSrJHUumqSvtHFkmQ6vi0u4arn2Q7hbmXwZ0WOXE8imO+We2YcsCzou
Djdaz7lW/JOp4KZLdx3ZshLghEqm/O28ututEWOJefcbPkk+otT5j2+7WyS1fw9pOKyKRU2UXQrk
UOQxk8zN+7hRDtcZd9sT5/txokof/fO8sxM7PSZz5Djhl4RtndWP6U1NN7ub5WpVmTAnTTQoJ2rt
BgzZJCyP+x2pjbfUHyPOkzDeROyacBSrP5vjKle4gCeQNAZcsdwkjmQt6qZvjXTVSvBpGqwf+EKa
S6DzdkDX1zM4ZHoUM0G+/sgneHQDu2Avd5lJlfPRr/TNuOFAZe7H/5b2Q+TDs2+Y7TJ3g80LZQPt
qiBKgZ0etAA1FhJ/wU74O7mS4bGsSRZeG0+90+/Wa4uTsrLIurdw5g2WbCo1TxOVMY+BqBAObE45
UmdHUnfWM3TopBg6fAFZHhZkhyPUXgkohUWjNd4q0iN2GD2FZ0KH0t/Yngnauvz8zaZuasaN/BZF
CXlyBCywYqRqo/gNTaUBHULtJJ+x+1H8BDcCzVg27yxmmbtPg9n+QMBxY7PsnsQr+vtwlUWbuCD3
acT9K5FoD5PNQ/yn+J3vXxgC+goU+9PajVWPEQ1d55RUdjxmIEKgLnY3Kja/r9ZGYMfFG5Pus8WZ
z0OA/pAeStMt8DN0hNqZ3V+QOvsd7tWkOvnNOVFhCD1TNgOJjZq5gPWN4vTmw6EYj/3Kew9GTYZp
i0J536VXNpPpmBuhvsuepacqBIWbK2b+6HYiegHCJm9I/0hYmayuR9cQNuyRQejmXUDNtVOyNEYv
6QB3ZOYO2p1FtHdRh52Ei9IdW+o1NWCTevyDlTozQeRrg+wyR+5sUkS0sP26wdrTtkyWIgMu8Di3
5c1Qo5GBjQchmBn7vghpvkDe6jNYP2zKZm+VsCWmEFWxcRPl7gJRkpPGAFQwS/2luFRPHgA8lCSM
x8Gk+ZbAfg8V13c78i9fivir6cZeGpZewKEVv6XmURU9XOxizq7ULujsqtB6a0KfO0N61+2130gn
Dbl3C4mcnaA7hMJezfaF3jo/4xP30ww48XbgGN/FUPpkm8ydOY/W05Lv0YzQl5W8caIf5WaZtEzo
gbA+2J9v6mjLrtBbHlQoEH7Vxf5BiSSkJRMqk2xrRKnIOTCoPjDl9e8C8B++HnKxd4Ohf1Z99+bU
CYUPGspqUJmmMJ5JVsA2e7uft5QyTZurVht17kipfXxCJ1U/kMkx8bnWUchaJ4IR0ZdaYxeNtrbb
KNC14EyCRCnPrv/666f8uMUKgAWSarLi4y9pNvLEoAfjW7A/RLGBTtwipZVMND5Z4Q6nAvgK/FqH
Cc8Zc3JKigcXnA9tNx69KTIPHLMoadhX7zs+KurOyaSJ5vivVHQqyef6lBcbwwuBr0fG+OG0qnKV
ptg9M/VlgpH6y+DKOeymOuWv/0VwUgfASQ5hU+pIdJfsZEsWwTAOdTi3+V5Wqmg1rJiOCdE0jYhf
vH6tbWrlGdnIoAYXFb2/wU2xbB1U9KQvasZhkYv/s+somOvhYu71aOVdE1rvafRaOEqrVTDywSHx
1U1Gx8Cfb5/LIWG2HtDzCP3/pQdON9nybULA4/zfvOBc2Ez9dx2bx+YQbAgZ4vXwAvalfyWVTgfv
YK6wNGP1uP6O9pzKD8WoVF7GXr+PZIJM295Lx0XJ80nBlX5zGUwulgLJ7XfZHM7/M+FRUem4tPmh
1QfwnacQCqpztChM/XG6sO6a+aNR+I6AN/pp1mnauQbMJY8SK57/9hXiGE/Dxb953We2jkzXk1BH
gGa5/Hz+YTAnaygWti6dtLZmJ1z5SJ8wxTFTCqGPA4V/oKWLEFUIU236WnJJSfv/RhVHcZsJuwpC
f0qwIP2sMEe9sYNfR3fRkhrlAOGSAb/y+hwp9106YbYlyFdGXhgkbUp4QgyYD/IcbALPGVJ1HCY2
NELwvqT6LThGh+ncDEGFnlWrNX0UrmpnLlL8LJfq2pXK3/OGxsHHlBnHpxTmuhzoY4JcoJl5tkTh
fjPGuJbFW+WRErsgN7/EcqoAwvzVL5EF0bZdXBawrBcyqJsP5uQSom9K366qr2rEe3+fuTxY7wZL
9isFX0Kw1rx1uH0nIyTLmzbdkyzekiB/ZACIH9DnVhZxQlR0Y2Vnx+HYX5Y228SVOSkerUYjgDqZ
v3PG6kRSG1VQISQlF33KJ3qg0B/boDlIIfP4tSMN0Ucw35mhLssDSR/B3Y4Cv43ozwKKu7MoQLJ5
jhw7iZ6rvp3ASVxNuxZTVNyIZznhZHf5mEfumovcMnRcEm4mGUV3oIC1Xr0D03JVatMBmCYgL8iQ
OTtq3v1vBarpqi4vxjs6n0P2joXipexZVagQitN7goRPqvm8XfkbTguWCEc7F7wCGTb8HA7HNzyG
+NgSBwwfzH3HZrxCLIq3hqLWUfFtQ0mb7W3NAnRVMgaC6zkvITfnVQ9HJEnXK2fso4U0okZzFm4r
0J8JC6pQHgbZkeONpVHfzXwjcWoYWqLQ7J3Z1OBKfwhhcA0gzvn445GnArK+ad4ir3pS9TfAV8kH
BcT1sPazs71F2hmmWxJquAzyVB6pzgisFXsvqnZtdZwlnYYmMkFyRKgJ358ZZUuMcHSoXdGKLGKX
4wdDrOYTMXr5dVbqib749GClJUr2tIgHvrexX6kcv/rbQ66relcqU+hDjON43V+jP/NmnoYd6JdU
5ip7NHa8/ulQzUKC0LfMhY5pz+nzSG1xn5p+MAHy9MJ6Ztw2iIw7ZqBFfA7jg94+GZC6NBMMYBoM
UFzFXy63Nf9Fi69LuqXXxCguVEZp9nGBPvWC+aXxH6okl/G/ppU+ekSgIHQszvM8Zjgkg0kn+ZVt
0stdu+Hzef3iZ+XleyVlQo2S/iekk+Uws/wuBNZh/qDLK1AGdel0tON2B0Apex+oS5x5DBdNg+v6
c9XioD2z0ggte2847UPD7SnjPrMUrKMWOLvpK4/w4LmraaoSsUhJpJlrie+Bbqry3hYICg+4VNIx
9mmAtzKleJvDkGyUXvBQprlwnTPt4lM3bR65acfy8BsJP8IhtKQB8en4fGtZwZYE8wPHw9gxIDO5
enMOdZXIQ/zUV/bwZogeTf0HZ6W7IQ+mwEkFE4m+iUDEskQDw1zvFL6MpcFnDcuwqSEdHTS9bxBF
EvzzAgDlDq3Usr/qCc6GQ3Lkm8CYUT0/kXPB8N7cc9RER3qNWqmNl9CFDVjuTSz+6kcYsElyXC1u
quZ6bJ513wEoLquiaykSyaLHuaiqdzMwF5FPLCMxKCN1GUqwpNHYyEnm+clHbh6npstrUrfL9x4j
2o9a0l5FZWsMH+rNsjf8HJCm4cRSmEF8mfANH2UvmNA/OOCTstl4UzqC7XFhPcOGkOqcgEsESOc1
xJlbzNqT4q3GpR4tT73e/HpnGd/Zvx6MQmjXTpiL/LFNkLsko3lFwjSAQdd0ALZNPuHgMWEcXIyo
JvgLLpKNWzcC8L3XzKpAz17bu8n8VRs0sy62LZIcwFGW3yzXpYCHbg0GPWnJRndtpDk4PUuAobOa
oBpG6X5YntSaLOpbl/30tMWLHvwfrSmwnGBZJvWcfMHuMqItqcPbZrnqNsBC9pSTNGTLD/BJOKhs
vB15ej3tZCSGJpCiXbn95E7lRua+bi2JuBi/0zqD4sf2WX14R02eePWcCi+lv+blDGlXzgyiOIhR
iG42oAa3BqeeuDeWXpCjZ+2z9MHYGHYresmk4cWCBXMHZTFkPq9/K/Mx3ikjFbAvasrmZNavqqaQ
zKTgVInUa+gcMrRFzplkvEuB1BSCdh+XDTIiN9seed6RfaAy23ZDuhS5SgD+o2iwCJxZs4q6tKXI
KgPJbAlm63oDYRpL7c4qaGMrq+9Zcs8Cd5iFUA0PMM/DqKrmHqInZAi4jyO6oSv5X7PFZdBuBURJ
taGtAZYx2Ur6lW1DO9dYPPNT0c8OlsDYiLjGi1zM0qTjXX/ECzZcYa4Fkiju8XoBllcNOS/E0Ekr
iQI/8lIiQXSbwFtmaSlhkzi969Yf6XycVfh6yNa6309h4SzcSRZ3wHwxHS0puIrsp+46bucatmSq
t0dHkFQJWyBWwrIJ2bqEuOQ9sJ8HxeqHGTzBF+eanNXFKCcDh1spmg8DsMKFdNZIkXA191R18/id
tSFDyNSB+OzZgG+Kw4Ae1afBdFFuEC+Fo/xssBUpS4+lD74CZL7QBckM1VIT/LZXnYBxaCnsQrAt
zbs481rtrpDLlo2FMPwq6FB8tpKs0Q5q4xUCOIcej1r9YWzL3GN9sbmrqcHowCaCWnnN07smK+pq
ksbt5Z3m2Eo7JbTdk7Zl2YWH5G7k2m8osUDEuSw1+DnO5wXJOXt0fHaUubj9bKwqSfFsMd5ba4ko
D3qmB1CjcaONTByrXs+U8zScsT/vgkurDXOjpNCXq3r1sZ95jAWKnlJtL7tO3/w7JT1zYjGtFnjT
q2/GrNYkdFn1VGGNuJeneJzaKwU+OdQup5ClmCfbMMkwu1FMDxpnrgnPh38OJ5wtJ7KnoIiWsNta
qs5tANDtdpEuumpjEN/xbJhegjcaotdRheJuGF+RJnERkBF08sCLwHwWpGj6qUK4ma+y22sPXqFZ
1TaeSALNyf/Rey1Rp/DXACT9TDK4o/IU1fGkffc0US4EGRPQnjDBQ1bXSZ7hbLdtP+PAg65/HMcV
Th7x3lRSzRJ1GvHaLcTiJHC1vj7yLcG+7pUsbhr6vB/Cma8IuX9bIUY/jD8D6SYAG+GwRhUzZGFh
D48cInkolfdHplFrgXV3Tu/ztJYB5WhYOrNx/1wo6ix6+eHAz7DWleVScKjcZ+oQhWYEw5H7jr20
CvUJnjlNjNtjxlkWwh923Fkec07ZnNq5xsD7Yi12lBExtO5RYkdf0q22B3Ox+mJmEEWtOAW5JEEx
PCNPUIQfX8FdQwGANgYOAU5tYtpyOyOaTkKddCBmc9RQHBp6nF66XrmEc263wI/t2Da4SAXv1JDG
Cg5LnqNeOKuLF8VOlZj16KBmgY3fs70H/bdbDgywzRtr1V6k8/SmN3hMQ6+yDZrUs2N33wgbbzJ9
//KenRs3CcgJXOwwO/rpVFBt8Dqo8bLijm+VhWmpC4aiU1u03go4mY1w2EKt+jEHYjGJRzenkKAn
klpAzbqwpolZ6KPZ2qCArvaIFZY+O9efhoxp3YuJe5lPUMP+0NxIuQQZQ67cWzqfoBKrc9U/X5cC
j8A1v4UjEdkLbBnvENfoxn1GXhWFbkeieKsFwmrGQtDNF5XcgYDgUAVfPUA3EdndShAadseQtKUR
sgchoFg2tG3XnT1MG+K8S6GIIJFH+UH/n4GFlfQ5xB1CZRME8sY7SvEOBWcVX0QsPnHu+ofwod2N
lOa3i4d0vr7AABGQNiEtkwcNLe+Novwwr3jRuyCVTIXT6TgejVkh763BwAvD/KFFYSWfMDBTCpGp
RsrN3/P6FZUCtNLwvBCAQ5Cm4s5fghfLcIvqiINzrGjFKwA59nqkHajy13Svb+a0W4YQmo7XlWy9
29rbNU3pWPzIKnlr8R45fS9aB0dL3n8u4mVjBpgQE/v1cZkHI6IzS+gqJNA18d/OvXNsOjq97Stk
n6029AusCwmYvH08eiLOxA9uZuqUslaEEepgUVOMgJ4Xhs/aOhUwpWSeJZBGEnnxKPAW1NLFM33i
Y/rWNmRiPVvEWU7K1lsBcnOvh9KKo8JV1S/xn5KXu/2IhblA8IzggzLRb0sAFusdsqDxe43jD17v
I6mp3aFLIwa/XBRN9MjRVkPSUcltcxa95xXcILpKDqOalVEZRCOVZQkoJh0NZ4Jy40J9+D1DQYwS
7JUuBdxMhMq5h8DxRYPq+YG44GUql5oCl0igdpE7n9aDRX7TA79mRvozN7tNNWCMZCKVnJOapLPM
HtJBujTUpJknmVDT+overAbH4ZuvqU3nl3JY+yrlPM8Vvh4+SOEx1Ig6jLOBrmqAdcJz7GdKnlHt
dQnpsFJIy2O5blLx6HMqzLUwlSwY1wuq57O6XQFOd2gfJM/Hb3rShvyaX8EQ/iD5h/Hn0BFXVRgH
NNa6kr2Yhp3SHUCyeg5dOjf56ZQyjz4qz0JkSW5Z0CWiViMOGEHYn0p2lIZK+jRPavR38trxnhn3
PYPiUoiWympN3EKJlYpK4lnEWGrBMHUH2jLKta8HfFe6WgHZjxnNIbkEmsLmrSmLBjDmyO9lVmgz
shHwRBqRfhn2JEDyXJk+6NBIRa1S6JKTeTZuievNnpyyZPjdXkbBkGF1vbrZqn0z6vvg4WDgw/x+
OL+wt0YLNh0rqhmmvYvLKMyIPOLEVFNzHaACnAH9yrNeRMc9S204jwJmOQr0HLNuGBrZ2eVRNYge
zB6MtPZ01u0lgvi9O6ysFhIhYLt7wUsIM9Z/qXMERRZQ4Y4h9oxSIrjz+vLcFGVK7y9F7f9MkNIN
kYVaf0UAVd2xGO5y0fmhJASemPmIl+RnCaFIeqoLO646lzK5e8+PAD7/GefJGKSjQWh9MMsGw2VS
bBlj/ei+A99243WvtKEPXOO2GwpxE0sF9lJEEpHEgrMjDiyZZhTFVDc57n5k7nFqrYKKSDDRs8Tu
NRPJATYhiK8Bbg9CWWtyuLEPY87KN08dfG8uYLTZb1uIMH1yZZ9LEHbAftZAfenpMIO0tMyVqpkU
AzXKkoxjv0scD+Iu/OEpH7gpj8KDW83FkpMXYjJrddJ3IRDBf+51ZAQzwk9KVjMrRVIXGLZQRikg
QSNkM3AdYyvVil6w9u7tfE7eDXOAR/1x7a+rYMxowLzEISmDli8Q2NkVIG5tps4Zpw3OvxdOLADf
+z+5Kp0CWUYHQdaGAjaNuGn8w+ITy85qxufzPXFZ9+NUJQTLcqUZzznPpNvRrKXnXRk14KFgIUYI
Q+ojZxYrsMhmKqqUvIFFEqrZMEIV4jz6mLBKUf4EBVmjVgZYwRyb+PPH1qzU/VcA1a1n5sh7LZj3
RtXuXjf0mIowc1FX3v190fuYFl/VXefYiuxVne/Z2DBArpUdZtZNVciF7FT06dR6Tw6PbpW4AUaE
kWZP+FW4UXBdTEJKP8gOWiFi66Dcc50HHEryEH4uPuTzGG/I36mnbWedDIzhp4bsEWhEIQUe+T+6
Bwxy/iNPact+8mR6JIRrGP4pW+1qIyPO/2BGIdnYL6Gp0lltcItfo/fuAJ7IqAhO9gxsp0VXfHLj
34rDTMl5WNVHic8Cmj+Nn4k7W2aR3XI1n8hPX+5DOgSpbU15Miad130Cq/N410RgaRpnMGAc2Iu3
yndrChhlWX5gQHcei7GtacDZi8ocIyhJA4ln9cBxV9AnlktsIaK36ai+07UJFliVzqpQKoPx8Gjx
rAe8AYZwGgnX7EHgoNNMc9uwexa9LDSt6/eayauWEUvYFn1iSK6yhuRYUUDywijb8reKZGBiBLdD
zmCdXb0zK6y4uM+6sT94XMsZJteHdhPg5eDAx/8wv8PATR1M7xk8dop13CSLLKXkcxKekRI4lbFA
wVrE07R3UkH5Za5PIC9CGYTm2weAQZA1jr/ONmwMq0Klka7Y7lsn84sZc5w5qlLPXHmEoBXc3zku
SG8h/xh4doc6aTT2pUmv/oRHsUVr4SoIPceA+cp8r47QdGL9gsSMhWZMwu/8fCgG6eC9jbX7Z1cY
Uqe4mups1SpuoTv8KleychVQyAz9Up7zyLkq1RSaPCGCbrJusV8WMJsSIIJX8IfdF4Wl/rky8PB7
N2b9iTGqh9q0QnBktJAR58fCsC6t1jHM/4Za9Aj19GIBt4Bl0WbtVq7fARldKI5E/hxw53Jrnbs6
sEKbkkSmjeHTHN/i3BY6mTn7tf63qyd7cWgMVAzO/xUG9/snTgcOnYQPyrkY4KNDn+azhH6/aRVy
h3tHhquYbYBz+yXW6TWZbnuqJL+zugwDD7gddSXexTll5YnhTT1fpf3EkupeFcPuMF5lE+P9wtPc
zoLTorcVCNolgw66zRqAuNYLPdEp55N3KiRQRbkYW2P4M3teI/xQQNLTc0ZJ1EQLC9h7lWqRJU+X
bhn0lKFoWkCFhI6RVpyghCuqs17BcED7feIzkHuWYWWtUXRjwGUGwEGavV8tOwye8ZVqdkozlyTA
1oD8BCp1oHHd/aWTmT3pQDyDfIkWhI6QD0AuUmY0uFhhikDDfjEGs9iNVF/TFU20Dkten6DLB6PQ
L4H49UYZfMuZYrUKwjqWuejXdsZ2JYFf+hBkEV93wDjMZskOju2EQ8xrKVUJ5jjBK5NV+AN6GgZl
38hYzpKylexKe1QeeZZuP1MkM0lZI3LC/ZLysJLBYkPUnoK6LV0N5LSUP8aidRByGHnFqsfor9of
9cidDk0T5yD/ybSrlJ6UzJfgmbVdeDS1Oo3aMC5Byk016c3uKRmb05cYbEbPyAhseNlBIOEwzjwM
IIs/iNh3qLwLcIyeRu6nhYl9bCoTHyod+UjW4s2z4IU+IQI3aXWqZ7K6ipZmyp/tufucgEEP92BD
Ek9bvJsZ/JODk5kG9CJzdPAkGLbUGVNWRWAIhqed7xdfLqU02WZci0VFZKfCB2e1ieXC8UGQiBmw
gmgFFog4QAyiZdTKK5MeRDw1SolwhTk2bcPgWYf4VZBoBB10+QTPaI1FrDaPNglJPUObiw8glY79
pSDFUOQTMbvMCKC7vK43XfNbw/EjSTzdcXWZqXtdIrkUY75eoEyLXcdymoDDEBwwrdno3dS7Pg/l
Xc9AT25m46bBBegxf8T/C++QvROzz/RiFXM4wRiee7z/ZIGikqrfldO7x6LwP0+1lKpLVXp8160/
A7bLEQLvcs+vxUo+cHjcJrdT0IMe2Jr4IEbLoi1+XHEJb/t3rt9jjEx2V1bHEQkQmeRAXqJMYbfR
Q/+ZPRN2wpjA8/N3xUi7YRE4CbhtGUCc/YJm8rwMyV7vkLSYfTVzEWH2VxKNoxl7o/BeI0W91Gk8
nkrd8uX62o+jcN8lWcaNKdQOXF226pl1oM/wckTdAupaxqOsd82VGndPZyHChEOKcqLl7fGX8XsD
i9rUuEK6wgC4EbqniLIeR+ikOQI/EfbZuy6mUw4w/SiE/6ZX/uCaEpRi7ryIs/iMWb5wGCqgYTMM
TiaaEq6q3AgPvSEPtpfTA1LkTgNywUJZSrMxBtXTMezguWLD/wUgRya2HZtfTOOF+dN/k/kbc90O
OB5J2vCR2mcYxWLCnVxvUx9jlHdOTHSG8JaO73HknPV7eig2fNGouqtPGtH1Z5ug9fO4oPrgy/eg
TVhPUfgHxkdkBEKRBqlgFsP3E1Yxp+ehKMD1FFSGyafZ6CQSZ8HoKz3CBdbINqAXCQjt2suU0RAv
z0BqIF8oxthxWUwmf4Ba5p5ciDIE2OhZrnhWS/dI9Vu8Fr68PakY5yMJFGnfhIb+ML6wXkPTnlOC
mBl6NRk/uuVRISw6URGtlqAek1vdL+h4JB1r8PcL091E3pfbNXpXvvh4OqIY/E8lDJmcsZEBlK8x
ornpyEGZN36umuHzAKZh0LGKfF4UJ7XpApmuLP0QBLym+/I1EcyHv1yaXPh2Xkoh/zDoQOW5S8rX
XcCbKImCUI2nbdfa+xa6v0PjXHGnK5v1ldD7e1f2/9pS7GSTxrIfgoao1biAldyC39zjoOxKNIhz
YxIp4xqgu1ZWS/YsnY+C5r1d8rVucmMpgf6Oxk8XYh6DpOn4PfNoSPgpVlk8Rl/qAIjCoOTy0scf
80hsTNhXKc2DDsKpyGyWfTYLOpmnSVAzcK6wLcwFDM1KKMliUockKeQl61eMXyw+6SEE+vbrERku
tPZpJJgzfa/dzjXLjlh1YnptSxD4Z8smRf+bEwDBm5oEQqEmeSr4RURXR7koFmRJHleh27NwVkdU
cIUggfVayc8/Httjc6NbY8JH0kA8xJBjuiWYqdO1VGWbnmhZ+QtZFa49gRmqvdL11UBUrVINK5py
Kt1nkUnXS30gB1BasNfwoqR1QL8X7S/lGHlstgrfaUdboMY0rXqEqkKVlRrXzjwGhonoDZZEHTBl
Xv+L27pHmb9q7+Q8LMNqVU865NhngddlT+1bXcka3A0Z+nEE4wsO56deSddGYjucYDRIYaC8zSQX
sH43gSUrENmnlFhHnp+yfrSj8pizgX9EOqH6Wcneb4gl+4rhVmuh6K8q208MQk6/ePJ/VS3rYlWY
7VnHlpmc4dTcla9eBvCvYG7RIjGrKc+vlp3shUp+yB+57pO3hPYTPfbyDErqPX4R+DeGbkCS09OI
n8Ucj+muXUBRI+QALDntJV1iYCjI1Q2wF3iPtK62U9YVL6oqFPvYnrERoPyjaxLjqiKC+Mr2FMmT
z/+sMRcfmnAeMxxxusAgaV1eWQlYs15UFJmL46fwQMn8ZMCccxH7xMa7cknJm8eAnFhNsvF6F6Ys
tKWBq0XFd3T2ijxhpgxHKzfCPmAUB7HWga3EPvg1GESIKbUgt4YRMKJ2FjRQO2r1P1Lxjjl9fJEq
A3sBiuwCvz/qX65/TXInNRuUcp1fqGHk1zMa7xGCYNq18hbOsaCdoWPhYBPzEjZqoFg/ISJUTK0Q
JU0P24JVK9wBn0lCqXm+s/imDLP39KICkb3T6EnTOOduuC/R7JvYo+gYEOzhHs4nED4yXrX6NAIe
HBo0xQCotYprCIK1MCdywitO/ByrM7iXrE78Xvf1JEhJh+fnOmDneZVM6CYr7c/UfjsuYeOOZPne
X7ECGxmXVNa6c17492JK/ys/sDe4foS4cj8SR89jewt4nzUBlNJ0goHoPDsn9qrCD2LLlSMiibWF
dYHRogYIaC0OtGA57sx9EjixO9jW0FIvQMEHDIbBKtlAe3CKFGHuOIkhk1rkyzUooiMDZo8d39J9
Cs1NYyoBm32rdQOU6apZse0awNw7HRtBBGsesRYVrBVW3KDcxWOqGYMe9KOsDz8SZTsomAaaylkY
Y/AeEWKSNZmn8A5JPg8C/DXkVukQBTbk99q3wPSVhgwmbTkN1rgOrRSFeiwQpuwxC2W1zGrwuAAh
3r8oO/tyEVF7ZXKx4ge9NUnfSZQaPea2PX5WhCrRlM8jXiyA70cEl6T9AOjhlTlsmjYlI6i8RbCe
xHmcLoZo61MYKxwz6xAAJIXYkqxE/CwP3UxYUL3o42EMS+2keSxrH3FArMNqeIu+eQkXK2HmuMrA
ylNKOv1wkAbBBBLyQqKGvfFUg8DIRpk4NcjZiJ3W/tihZ3glvJ5vRwGAsTf6J6fTP5iuXDSqi0/V
GTZbMoYv8rVmwFHQS/x2xtp2ZX09m0WBHBAzjCldANDQkSpuGTZCAa1HHlEtb40VEN+YxSfgVKdE
fG5qGzsEtT39ruJAlDsxssSO48KpfyhfU7/sSJeJSgg7h4df0qqVi4eOQd0+LWZjEeW7OBqzbM+f
HzR+3KEFouG6+wM+4D06kgZ7TuhWbuegpb2jstCUiLZemjrqU0ZcdwQlOA/xnLa//ct3Urb+gi6s
9sjePsz6soRV4niiQVl/DJ+fg/cbOhSCaedC6uEOJqAYwOKy1Q93ALbVmzcMcIImusmgo1itqMVI
sUocZ9xF5oPQkcEwhnVgZDqrw+Gpm7jRxBg9DbybHbN7tnIwWfGlT7D3kFb66EhssCM3ol8H4kXM
ytlfEyJVrwP8/Wysw0H+ixtHFgiKQr4I//6girS8Si0tMT8w+Uydsfo1upBMqyzhrgmVtj4pSpTi
B2l4lRDiH9+FsF8nMjjOsVIhA9PSZ7TJdDFk7gPvgDXb638FDGDM8KknfN5T3/+33D6YMVy/LltC
MPLiCS07dJ0DKXasK+Ro5OUYwGDNcFjMPWaX87DZJgc6/0TjLFfbwwK9iOmR7/umFnuXd58RXuwY
xxRJrn4q/mag+1q8bOXzb5cHrAGQGBBtO+xKPE9dq3+7gMxKsIl0PIJ6tsKQEUIXBdiGBij2J9Jt
VGd71a3Ke0pIERQAkUvdaTvi/gczlHfamVTnNxyvnF4OMSOqro2MXpBZrNG1Tw1Pi8KB3S+OoSbk
4C7eSFLwdu6roN+sfJr8LcldW1YhfujBIL9Vd2axH5WjEVjtqJg+uFGDw/2QEnG7x9XHTa3exqKd
H8A1bJEPsufi/jz5sTdJ355tTNCf9Rg/I6o1NbzxsIW1WL77YsfZ1MU8H5Boz+xI6WDuIhaJ1KmW
TkfiyEJe/Mzl+Oje03sqCmm7WhCJkC2leHWR5OUKabuVDyFtGKj1yz1fphgrr5GaKE/obecQCS6i
sR7hzCKelMuoAK1RNBtO1woei99wJ9zR+F6aHirg//CdomA9jhAI/nQG+ctfrZgPCiaRT3Xarr4s
n9AEciPlDdbGKIeGLboDV2o+DLfRYC9s4sX+tbZQ/el0lE9MAYK+y2f/cdMIpkSaMWAUWDXJ6rwY
ZuAeYQvmV5YkOt1OL8Sv8S1nNR5jKCFyMfC0U7uEgK7wvi5eXLEt0O3gFCOsPmUhewn1ZRTvd6DK
IkcUWeBL/j9Ey32p7aLN3YvNgQNJh8SLFODwUZUA/cFky24Pb24uEzA6xXyZ/8M7StJYbvCxDnCo
YrOdjuuSYU+1QC4XlNWIaHk9TVwnfHuEfvIDp7Zcy2ZyUQc3lwmu6s65y8+aAMn0wtmQU97oTBtH
0Cz52Vvwfqx/TTBRpdJI4IOvGXewSGV72bw4NPQ5wGcaeLCh6rawKQbgYB6O+adXabFVjFWiLlwV
Fii5EQHB4DSd0PSlujZ3equs/YePTPOqExz/uJ+x5YQpe8fkmT7buZIbmCuXOCKMrffzRo80CwWE
vLek6fjIHtODujxf7L3v8FIBrgY6MPkTchKHX2QuoUkghGvlP5CpRmFRRcasPAU8A6awLnj0RMbE
rSCGPkg2Qw/16/LxDbz5SbVvkzV3fIqEFzLCWXMc8MZZnctYYWswzx6eVUWk1KCObL5kVwDsnKm7
XawiVcF2XOTwhsAKQGzynB0Rr925g6i/y/Ygorz+bUNkWqkNb1jZEhBANcGS4xskz83yweM+CqI1
JOTB2rX3lnic0HguVDWWOe5qZQwNiOUUIAMcz79+9xYekU3duyvIxtcMqy+Lognta9cp7p8iQg5y
V3Q45nvB2y+P1EQQHVxBxZFUC3DJKHv5OpqVN8VKMcbqnSUyon4j9Zhf6HZXkNrg+5kbbJxxV3hS
TeLNbJzpYrVYJ0A4gKLXKNRP6uEMqHoWqhmCmtG//kWQPa6L+RCCf+yGVgWeMQPdDz2gvQd+ziAJ
MQinh8fZwLAahU6a6KcuuOVYsBkba3fz6XtcwloISpyQ0EEIMtfDVuVptWoXg5gKNYB6mP5C/M59
obLAftsLVncj2BnxgLYkq424ToGIAqFKNGnQgp5Joy3Z4p/6WH4ZB9/IElO+9zFaa7FjOyh+QNih
BTw5Yq6LUUj3F4RdTdrjr+FGSnBBT09XrXK0RCYpEjYoakf7fSolGaH2o5Q/+yayhOVlwBRDuSyw
kmArbImJx/qoq1drsQMj4kWTLtYxBbKSYPKnKNZhXKeF9daqNZPl+YJ+Dzgl0o5Xs4E4mBGVHzpw
CcoDK8/kyuKdWQQ2L4hdCye/WMuJxN3T/n9yBNagynxpHtUWujot/DOg58HzwSsH16B+Av5ENWjG
uo6J5tS0i/2W5wt5RevmL7ETDxoh7JJC03c+Z2fP+sMzmPMrewMyCKj2Mb4cZBi1z61ZOWPMXLj2
xcyyX4BUDL102a+OW3bLavnelZcgmJgQdRU1Fz3jJsnwg93nG2JommLiQpglIaZd6119DIRv0Y42
wwVQapix0jtjv2/FnBJgmaDFTTFFEQ416/1QfT5CyLyYXZ0Slk+t6rpXBkmWKR2KpLKuyaJrE9Uv
PgRT5Z4BrikyEtGZKTBvvtyaT/0iLsoPU32WB+VcksGn4AHfcdhC0dmixDum4KIkw8hBEzxUDuqj
Lf77C91ADimKn5iYCmDl56bfFerBpnjwHNpT6dbPh1Coh+gpBChWk7jmApoiWCQ/Xmlg0xhXzkpI
PcD5VWCu5p7hu9DUmleU/bxwahd4LY+HDgDn7IVmF+XhNRTreYHz5npY+Tcwpl+SEBPgvXiSnwut
EblOzUfNWWhkXvchJJvKmVFt5xswvT2nU1FsZuK/5t8RCjSLmWnf68evady8xJboIoKaFw/lpLqL
06V/5nXcvjGkEA5cQYeiST2ayaRjKpv1LrtquaIYiQeYp+wHQy6/aXAL+GEoUG6VQur8F06pBGao
iNh/1E+8U7IZtgBAnpikUzs10+PgIouVpulxQq7WB7QpkixP1ce+QoFkrCbbhBTR9Rfa+enp3MRh
o5eGaJXD8YcMOe2U7HgDMkZIzFACNvhcM/oNpA4vYqNoYIsUOJpgTXMJFD/kJAzmyEJ7VY5/kfLG
OC/70yZW8mS3o6geq77D8ffIwGa+iRCbLJQL0i3mBqySDyEag5j+TIzXKKZLuflj4yPCHdcQqntx
+OebnMW7EPkejN55hHhOuvNhUXIomArX1+wH286tU4s9cOP06YgjtByu+++dn7QwrJ0zGNCa5E8S
e3pxDaCyVJyTfJUMTtNpYGIjeATLzzaWNov8wxXsFANWbObpFEFt01ygyovHgGuNCqY6y8f/WwD6
wHv0ENogxk98Z1yD3p6H5xQ2TCz3RSY/40VLDdlAbiV6Zf6cvQE+oQwJBoTXSqxGFqNcF/m+KywZ
UgCHW69CTCUNJmW3zWecIEVE5B7NhLRhimWAuh5hopc6TuxcSPsE/XVzcEC5vapM20yAKcmL5pc5
3ZjvaKuLyq2PAXI8iTWRAXEGQygwb4P7nPOHzc2+HznOl9jKzfUQUTepwQPlvVGfO/0dVZJTcNX8
qY4eCHqDylutp9IuxI50cMotfgLkUyQtRYU/sQfmLtZFrXUlmMMggyWpRe+V9i/idqEFhRfjVWEJ
1T9+3kFrzsKVLqmtK51Ec/ND2unlA1umVALVGGX8pOsH6iwuV5xR08Qw+jr3/gdb4QOZLcOV+Ihh
UmXsmruW+HNUHbWk6lCSa7Ynx28PzVA1takCbi6C8ECeeKSxUdtEB8eH1ZHsXFF+FWTXGquEnnAh
vZiH6G2P5ozxuCV+bPIORBQimLGt/HIfJGjYEOheqPZh5UoyOAUWf/2eCOO4X0PfpdLifC8005ig
k2SyGhAPwK6P+nFCIQaZCM9Jg/SzWDNGUnbM8aoNRBELvSLcOK3RkFTw3PEUkGY5dU6px7o5sy4Q
QO1JmrCVhLSc+2VQ4Q1C7ykttxdgd54UWrwrHm9kssTyc+9CP5bKWm5DZj/mL0wYebP1r5y/OiwN
Ve9W/kegbiWPswciLc2svx2UnLBf/8hvsh2WuRpW38lxKCTvaFqOzN2WkmUhRKK9krKpxASx8vhh
uY4vQ0B/8E7rwIApZd7wRGu44IteMneTbHMfRlrhhF4sd3vToM45bkhYz2uf98tULDubEmTJS/Tc
KYWtLqK1oQatJlbkP/YnvPvYs91+p+x7s3Iy0ZNHhoyMuJlWqysKP7kH1T6wVejq5Syj7EV86Wr7
/iB2xQ0daZAQVn/fKQh5LbSIDATjh8beOrd0KxgbklJbK31ZvgKWhLlGqKFZCRNSnJdgYvGU+CQW
4XHHhPGPeyjXl4C/Lh4NueGNeYyF/w+amiZOMIxfkd79jzGpyIH99HJklv97d6sSKpTLbiGQfK6r
jZ29lxObiRjLBf+csVABEtnjTm9cGejcrLw88ElEMCTqYoLQbfvcLsWYXp8InJOdFczS2ZG+PrQn
V75nES8wTbgfDGToW1laG9x9F3Y7ymmFWwbKjabvjZMbXXZFPMiZEz2kOnjT8uhONTa0aCTCFSO3
8RbIpMdB/fKlaHhRdcxE/3zy5TTsspRTaRXdLYv7Pq96x/RSzSh4gbsmj2/641X4eNnBQ5kcPBCl
HbpODG4KBF4Ll9uYQI09RE3/4WUmaBWcflvCDNZGeJY+y5DibdlrescCrSMSWn1/0ZAhfZ2l4Hyd
2rT99nXgcIWTCUXHgxC5dk3BQGn13lpBhlm4OGH+oafvDEG0TajdJupQFTbQsVCVlZFH++BSx0Rm
tz/4CW2KG4/zcwBqBCHBaaz8S+RRihNJZNCayjvSFz05Rqx4PiymCLKmEkIXNnKv5MwSyWlgxWTv
FMXxBHk2MKCjMf7LbnIfFql/KxGVEgY+Ql1QZwHl5gGtHN/cv2tYEhzSfjLi/uSXziTsT/fEM0Wp
83mld3Xhw4boLac1mFEj4mT6NfDWa+tU6nUI6kxEVFXbUNtXXe1pcAyQkdEmwM56w77lB8IxPE0e
yIm1Igyp4EvS0hrAH/ZzYGtNy9EVK/6K+RbeXykAwVnZ9DRrdmbePL8Kw7TYj+sFzXD4ISgGFkhk
A3HV6/ulHmvUtGAl3X4Xv4M0X46cbq1ygXkeKYxk4s+Wjx5QUf6cma+jUSKkaKkyxtc+PwRO7C5S
SWVeT76xHkq0MExz0BW8PXjAdwAvAOSNApNwvbu19OgxSTT4XvQ1GAttcDHlM++YO4UcPwZ18uf8
UGtYszcC4z8PU4aYo9Yf2hseQFDuQeSwOwH2Ljvze1NbXAOKuwS8BozlrP/SuDRE4U06pUu1ttzo
KV0Lvl31g8/Mu0fGdn+0um4hkDk6t3WA+faWBJUtQ9eDT7hzTXJQ67KhtpW0pvAO0qSrIYOVa/kw
3hf92xUlFJIFPHefSHSQMKTWAVUKvQQLb9g0pgnIXg7p7Ib9x5lNRD3lml43wW7B7YAYhh8r7wBz
IlBE5Uz+J8Hp/T1Dd+FDndIqLnjRSNeyJsT4YXS/EZVZBTCxZsbnKA8zXTaCFOBcI1gpzpCloMNN
O3iOxbIzKoJDw7iVDl83C6LPfezFN9FcS58enE/F0bAAdT7n3PJn4UXqrjCovJG05argndz1j3jR
bcA/OcCch7lhwe38qvcTrxzqHjAAPwX1NsZ5Rsl43lwmmkDb6pglNFhwjhdxyEpbvT55zTQ9ayDy
r3cTp+zXG4A80MzhYEvoJgWrK69J/uTKE79oN3WPMXyqydur84Zq2qK+v1B/8ofrnZxGuSADmliy
rfTnX5ijjM/ilYHhwY8wWhi4ve5w9jcUS0+9O7V7ebrCl+VspnMOcJwtd65SPA9TAIwYZ2hP7ZDw
pywWdufhE/CvID7GD+NFCOJkGjf5bRt2UoepRGvQC+wcpm3vWuYu0ybIlj2CSeJ/UElw9cDJ0WZM
Z1gjf2pCKBD534lcHHyd93XWfvy7KSH6IAKj52MB4bnIjZrfGDkL25GR1g1RW1mxPY6V60uAu6yL
g3vC7MPlMEF8tYVvIagBXW7N7dXh5Up+LQ6NT7LRzVjFROcbdZz5TSICWMKYZs0ZkDVKxAy//xty
M37kXlcq3j6AN0sl9RpNR9a+klaKsCOOtpHXQ8f25aiefn1+Mpqabov0c/4xbrGRRTOtwDAG9XUT
OjoEKqC7SKp+zabBmyzVHYpdTNNPU6b/KQrwX7xl2IkNkXK5BuNt4ULicmsPJGZ1B2XQX0px/gJ9
pe4vGR93jzp97yde45j/ecRCOUEHXjGsTMpCjcAz8Zk3fIiMT7P5PkTD99tZaHM2udnnCvZVpyht
uZwuuwBhjaoWGjSr9LzZgQT+oEd5FS9rvkn02qPB+CNnFAoT5MS2JFt7nyufWkUFkqLahWeb/S95
sM9oJiob+mdDZ8ayJwDRlR5udiH6mlZazYRB/I/y+P3U1i2y6iV8IVViI4NO9twGjXlI6z7b7bXl
JzyJibwuKVz8sTfKTNQW0MIo+qQak9YRA68ULKnS3iONR6g9e2WynC+54g8PtDj9c8Ac935OCQNk
cgIcHUHNVt9a2vwiPi69QnS+GOPHI1dC3AcTkwpgGrDbhwIchEKzd52fRXfR16z8KX9V3alfXZNg
pA3dUhcwXIkeDYcJJcP10fV/jxD6vhiUlzGnZIP5bju2On6pYHUGHrsfTcRhjqQjy1B5rW+jYg6F
MOSdHmmRPgX1g5pxriqZm8ERHzJ3wu+AsOpqmcede6Hc8Y0W8d3XhDd3e7NIxEwvFtH/h8ImsoYL
Gb5E9lLSrK3DBaY982y8BhnDabHVbmu0EGkZ01x3X0LI8KIAqK6AXAhtqlOKBTanuqc67mbnNBHL
LXNahKRsO3ZCezV7EgKRShJCzu7xeyyip7jUK2aZ8ibXZ+BmCZpsiw3TUANSdPnZdr7Q/TOIXA5z
NbeSNoaPzpnPgTqlTpqiIWIO9J9mu54rLaC929HQjiXY5lJkKcm2hQ7hZg0mAIQRYIn0x2xUzp7J
Hh1F3lUXr4vYgjzVRcDOqYXEo6lAa4KGODhKTJ6w3ml/Ci2m89j97UoQvkycEDkpZNk96qRIAG6k
/fvt10u6QlHEuPgm15x1FDgmc6hCbYCxvI8oZAoWmOoajmDnuezjqxQE0tBbTmyedrV21mE+HNVt
FoJBpX7AhZeK/mTfsOrS4xcu/OaeiCYVADd4OjVw+v+h2YCkmG1qGuKxgSUmDzJfLIMZK0qYKljv
l4W+58mynK5GebJ2nUoKyjxCwDjwrXB7/2quirbn7zJMP0uw9iQNkwEudCIhjuaayRPQdQ62HZx7
L11bB2PxqIwB10Bdve9g+veXZrxs4a9QU5o1L0OK7CIc/om9j0j5C84zT21dVjukLpJosDWpb5V4
JfpYKqG0Q1vHgPEB0YsQMtqFePeRPeuBNAYbodpTDwGPzpSaNIk/rYHJVZHrXYc4YNj+ANyZJCgm
yJjSCa5rCFQPQc8FKunuXiAM+zpM9iFPcYoafe0+W5rka+rRQlqaTKTIpZPmgpbmjB9kgotYmoQs
DRzoCCxxrJoJH//6qm6bIRYBac4E05kzqYqoXV3cWSfBwQXnk5b4QNCjK6UaiApy3xlevgF58sQx
bd3HbUMU0sdA/gcjX5KXZcuWBkPkvOOPSEevT/YzJEvT4NK8pHrPl1xna8om3oX7WhRs59zP5d/D
T++fu4U6QaDW55UehHsjbjSHlDgtBG+Js+nGaQ2K13X375/G82sPCDsTq5jk+zqMQSEhfcpo2YJ0
VCea9gF8h4V8Ly6KP8VEKGpp5swxC6Jrr1sZR4lF0T+MwTNmE/Z9lRjWTSdV49sd+scpLY31JK17
zOl1q7pGC5Hy2MZ6KPDrGo7eL1pDgFr5oneoRPKChJiDrjDTE0Uc0gG7Y8Wm87+OwOPePmDOYOLe
wLB9w+URYXVybynet1CZ68FeFB829yoymwvNio2/ekKQvkUZTwYeOeHwH4vzVYoFi2O5EluYI4pS
YfTxGFfxfj8avZKusYXvAzez2vsf1QvTFcZFSHMVvRvDLiRiM3yBvBt2Zjb15W10EcmeTHTXmjA7
NqYRr9gGGXJ2/AC6AkFdOS20/FKzR1mI+jqsGzUHsZdV/zKiwRI0CGbGQL6PVjeSE9HMFxXhX83M
8kGtWagwHbX5jJDb3n7jgPpqDlFrBs0NZqyAqY/mjlD/7LT8z+FBymznxazGTtdxbAYE/A/s4lXV
XVbKlPqriNzp62v7ILuiPam7YrA0N3SyXLW714dbTYtfvMwJjz7uPuB/H4SvbPAmmfYiSlQ3ocqo
SzHXWT/4WiRtaHAiGGMY2egaEZGpOcR1QtiuvVjdqLDo+QV9Z4yI5n5QfCfay/pM6CC5IdJ/zup4
j73TCs0Pre2TT9tOlO00YWIQ6mwO0PNKE36r5Jh6O3dxpm8Ymz8vPlBXTU7h9U0eE5gZLKr0h5bz
oSg1tC/IioKGe9gOJc03C86iBGdta3lstE6qp4bExdPYL480Q1w0AbHyCIXxSQcrIxncU/TwKdHs
+DPPzzt/qVHelWjQ4Y2vanKuWYdktiNOIefvYcjNMXbtVjaPpcH9wFvv07rzCBBrIY2DXjv8ZnXV
PuE9VFNxnJdTwnfYYGTv5IfS3X5kbT1DJ7Vyhdlta8qjLTQqULslUxyhAgiRKj9gWOrRoCMPGCZN
wUtQYkm7Doe1qQHV/NX9wqyka92tbsioKW2rVDcFO+V+Xa1T3XpTkfQjCTS61o8G2eO+uujQx2dk
YXDFI052yQmUVzvAr2eda1C/OaNLjN+DMSA/a403Tojn34SP091J9udoXeesqIzDKlh0xau/MEkw
PmkQN5JL2QOhuJUd25E0gugeNMVyr8LG8K7ZMoywPJBvzNDccqX03P7Dq/S7UekSYHN20nUs0L6L
JLMbKyCI+HTeqEnSKmFCIrndnN5rXG6YIVskOKqpPqitUPua+hCveXJvx2tqKpfRktUXB2yMXbcD
HJxkRkTjMXYWo8rVZbVSt9hJAhyXpG4I/K3nquy8SW16SkC3yT761nmVSlRDvk4NgqZ21lK1ptoC
tXM7ARPrq6qxouchQ4WpqP05st8szinVxJ2Oe9ckLMKiyCc9TSdMMQvzbtITNei0qUflrRuJ1gko
E7rwI2Lp7h4tIUCNwtv4zE+bC3e8NdpFnOFkNOnXBGtmPwU8jkgdrWyEDdQxwZWax+k0sCxUe2ud
M5afv+Caec+n5Y6uo3dTtZ+vZO3G6gOcLcbjIZeEtOXCcWdwXQtxL7veFbo1OPMMVyHvlXyQRMSX
s6dvC9myXSzytonmfK34SwgtvIcsnoix2PNd6DT/7MaiEX+Dsf3ew/BLQXtvHmLS++nvZcBMwkHp
Ir8vFKUI12+C7kpxvi60LshpwWj5NHlvFNce8TzovYtB/QDw+30RUAz5nBSigk1t17TC4ZSbfILT
PehKiOsDPdaC5tllWcrK5XRjG49lHG7d/NEd0nQpLCR38iK+xj4t9pXgdUBRpz9pFA1sIBY9j9hi
4LWntItuZyS60EBd9UX/2h73T4WMBgT8M1ewBv6JLBG2HwS4OKXR2Fp9Pf6MS/ns2i0iKGHyPsov
lr5EdscZXpSRyrir5B+QtOfTYo2zGgXi8EY9RiauYfv5dhp8j628j5cHXpapLq+iPm0F7sEFzIZm
2eAeyUc3jq51WhtQ7wgRTlnESviyrHxCGJOtwr1gyosltoH10TCdThq/aDyRLRzirLmfLPT+/AvH
lDDhdBB+H9GTd8ID/ME9wv2VItc9LmOfx06/LYZlsD5dwSffur3SeFlH6OafSW1/eMIcdmiWDhYu
eDG4Z6Avb6AVbFT3lskyt/aD4VcnhmlNFmz1x0kNN8V8M88KqrqbKJjzAKUhkZuUiW0J+7YZwZMU
2HdXc40D1cy2WBTobb6Tan2d2mrwUczVq0LL4CUUgJe5UDKzOXTou+/FniMNBaJ/sEWc7z56J2QL
JEjNJydVbUJnh7zYO/i62FjSI2VpYe/PrvQxbd7mp8GQUNlwavrMj4/K9Z3lJwaLn5lh8D/NE6QX
6pBD3yAVnsxHBLZBYTqsa8O/7pzfQoNi+RK/TQ3B+v8j+cz1SB2Vl0NPuS757ND8HRKVO9pd4b/Y
it6680cDN02HhIZk/nE0+hwyuIEAFL8AJv7BzcKEWAz0YBjUgAAvsOs65k1wu+aTC4+Ejqn1CUc5
gkaxVMjjwqMFShsFSKkMZeHQvnddWLG23nezPYU5SJyPE5vc9e+qsADL+LpVpJTMtmv0HPWjPNxf
cmvYswMgzaBF05BWxtLDSXjMn8EToQm+1qh5bNQrzw5sAJkec7rEiRLJMeVNXWMM8Z/5QFsCiJkK
glqtseAshW8QrsO3tk2pzXnlKO/b7v3FN7VTdi8SibasOPOJzbdQ4MbArVTSkHsg0Cq8Cn2Hf1NT
FHziJ0xJQ0/uhe52Q5GF9+jbEH2w3YqUHa80hxd7lxTDWS2OHUJ5Utf96T1vyvfWwNZOldI1XHiV
0m17gkT0jMsHzitlZvpuRQwS0MUDVOZVg5aUMcJRrZgE9h2LzWgHfWFvAy416rRpDz8H4rV0xK9o
dbz0J4ZHbjj0MRVY+IRCsXBqy3aUZtIct7aAXRtDsHZS+bQwj4dfHfq7aGAuTqRw1SPMXqW6u4u1
8l23d5j45XNx+WUATbBZKnJIs1EwYHlBW1ouqA1wFEK3W9OVSOLrL4K/zedKILMYvqSvq1hWz7/t
/pbbkBrc6B8KAJyRKGyPYDSsARo7XWHZPJ/a62Cv5mHV7e8LW2vK8mN0mP1BKr5W9Pa1SPOhnBvo
G0TXBS1HIDL35qsgrfjYXEUZq4oYQjo/EQClS5K+5BIvxy9RUgGCypmdYmz03GARXa6sdtdaGGB7
MRwTSdj7eCmPntDa442CVb9AAILnjq5WvCW/Px15r8kAzTUsyw8QsM6kttcvSX7dJFDb7Dx7MzVJ
iOduWu0FzJ3XTJrRLSe9kfYpKQm531QMw9K6+ojiuevCwSmnYeSB5RXA7Xn0Q9t+faQrILjanJKH
RhiYmOFs22r7Gy1m15a/WhmRKcBDvORBYfDCUXe5YCmHCuH4E6t+Ma0ZqNL/vEsDtQfauF+IFsgS
Pr7LUq50/LPwOFOS5Uukx+zfftpNIJVkmgGCOCmOLBM6eEOs8mL/CgSZL2a+SuvV/Rtfmfdj9xk/
/rN8m4iaDYgKPwqTrNgbBjihmmmWnBFzG/jI8u+cQ8C+eFbGTcuPsRfCWIuk3nimIDK2+bhfS/Q7
naKbDkln57jgwHCN/BY9fAR1RJ1sHEmJwmO/xZKRzzitmPxioi/ktTObxkxSFvHrNB3/jqpFVuwg
G151yI8UiltsvWdrEnrlQhxiYAVgPFBpG1/TIILl8lsydfXzQazrHvP3Cbm0HNfHYMncnPUdH4EH
r9Yy4R4CUCHWJzzi8qZJVkhwYRrUMi5/SPNTcMEyOTwFPW2Gsru6MLvKreRjVkf1paYI3I4rmRi7
wqL/fbMInxg9aflEh07NJ1av89UJZuTncgXtY+KnFnKUbiujF8q8SVz0EqtudR0MkKiXIJyxLG4s
D93LM+Uuu6bU8yn1KdEVNAgr2/rwhIqGhe/6V0no0HHfOwoKEY8HRHnyv8m0infHARfpXtyajMR1
aDkV6jDQQW2g1WnOjBB1mqXuAvwK8FIxwDoiBkkEZWutyTbTJOvEMr0X7jGeLjslcD3wsA2hBrXv
OiKlYf6FyPiSld/am68jLOkPX6df9YfCoqx1Fl0yiHa+YbJj8pnXMsyk5oL+f1TKLnO8yUdLaIfu
DgniVLZJ3s2FOMvX609kvFpvIoQ5hg1q5/F5RsKE0d94QPppW0eNPD7omzFi1rFnc6Nlgm0usIKq
WWPEaqmLaI7vtUfcikANvNUtusBVG0pIQ/u1cxuyfniO7azBev/+fPLS0VC9Bz/mFkhg4VVeI49n
jGMWtNfAFkc3zabDjkZaZTllwR3mQnWjue3WT5qNTEcMieZHFkBf9Q0G+oZ7fCCAW+q6zbNufKeW
dzfbmUCmtHFH9DvHCChFwvQ+4mwAddcObDfQTt0TBhEfptcZHZ7/isCgyD6Rqlv3i+rVo9H0kPd1
dFcHbWWfchkRKMS0vlE//OL9Wn0cQ+jbfnFV/B6RbHZXiuYhOBbiNlNm7vX8uGnnKUKktNpePrnE
zuiGAouVpcml2/DjUAyTYDoZW26P+5NeoAJMJWaRZYaO3F8vpJTGAo4MA3a7mtqnwVnGLnCg0+yw
MxzdIr9CpySJWmXzBGObEt9zdUIl0xA3wrJQteSWGxWrYRLrh76PaguryHxd6WZQVwJ3qloVC5DA
Qo+U03j4CjcMSPE5u3GjzowgqGXYkRTDdzYbwhTuuXpicUs7eSiZlbXylddLFPBPtnRYV661fOmI
5RRA2JoWSbBmIX/VrEyrc//Gw3qI0Vh2XcM2Z9IPOK7JpXSxuBO+sAaAB/OQqjs5fMtn+5aUSRAU
2J69URttqLKn1zGPQIuoVJlw2i7QvnCQh58P0Xy1ulZe3JnZU9eS6AxpGvuhfypQQ/J1+0CQdCd1
uH9p+/q/fCKsi7imRlysulAWSF7XpATTNtzd9s8KRGMf/T5EWJSV74SotzWImzM1fMcWpCn+vxOP
RS5qSu1AMSBsGro8kaLZsuFutP4jIU+CUc46HkKsvRDkt6XEXjmrTeN+a47qvlRgoTz7/SjSLU+7
d4FIsXNOVMzXwIKVCMKrN3AdnnkzoFMwt8Uo1Y2eRCf4dFKPtF6VPPw/LmgeolRUc7gIwmQoRF6B
t/Xx8bHv4cIt9zlTPcT7CyYr9GGQhrAozkG4VD/NOXkkaCU2SGBDZvpiOWw+lheXhMaD8pf42rgK
NI+IK5uWEWe9spA0j17DA4G+xCLC1X/XC2K03vMpK9/RS+MKdQTIeEqfpzgC6LQTV4tTSM4DEMq2
HkbSWmOooxhMAQFHQOFqwcRgiloYz8ZERpkoMyev1iKOUbkYKBOIuyMKAgyVzvt7uid1SS5XoFxY
06zInxzZfaBNneXath28aouwpQFQqzPVhUIiLQyas7Fx6bTb00J896JFNAwIrLdNV8NCdyCZ4ZiS
QosbrYxCgTaDRRfsS1ClNIUW0A3IdfW84IDGsHwynjWTJ2x8kzU0TNL8fRkHgJbCGdnfBLER8CJo
/RY0+/1PCbg/I1wfE7EZFMqkqheqz261s7tJs15dF67eneVW5ImfVavZgmWhDQdF3ZImzRrCI4d6
4knWxao39VU0SkQPCye3Nlue++u1MMNofJM34V1kw6kA1476Rrq5WxUWGVoVe0IcLERyt7KldgC5
3D/Ot51dEQMfmquUlhVm1/B+/3my8/46iUpE+FDnLj5Zn1T+0oJy28M9zl6tefpohu4j199f3KU3
moNzKn3yfLpjZJIeDeWL7O5jvFRgq7yK5AaHd5tHf7IaZU84yWltXtDl51LzgUNsEmAOIaG+jtuD
ISp4qF05A/rYTi3nhpsvs/OuHEO3Fx9iidqJJKAfWTuXbmbhfSLEQQH1NDHtQLVZG/b7SaTeskNZ
xBmseCHmeaWsk+D8yGZ8bqxHXQTnKzvSesafjeenxHdK30FaGGYdstX45KCu4th+kPVYLXLPHyix
q9snDepfYFJIzLAsSC4egxLeFfxeUDSfnTFQyUNK4o0CjWPBg5xGvfA9ucAe/6cPZJoawgPB1tqj
OYjaathbYQq+SA/Oeqmrja3uET9ZTaD533yxY9JfXiWOB1btzNLIJuQo1GIWhoMyycwhJ8bxvJfZ
V5C+WQ61s9AFDqeJryH+nwFdJI6SxtakJ1hcG/n/VR6+ydVZ4vqMG+YVipUi8EQlD145IGIYgsDc
SOpc7vrw3tm+XK87P87zv4Z+5lwSCfMNN4WSI6mg7jHT+YRbYpWlUrpXl8/M7iQQfUuB4GGE3Vzk
IYrZ/oLGUnqcdWRiTYlKsPYsqhXND8oHFCjxtqfpoIS+jDJJaid1IhnIDAmlgGwnCdisuQJQQEzH
iCb7Yd8bhLH838OzYxnLaynj0g/SNyjyNlSyh6PUIG527DL3vPdQ3HkNPM2cA+b5DVBJlvvu4wFH
THIDsEcbs3ys92Iv9rwCPz+iUqIPTyBjVEMttX7Im78OLYl/5d2r6wBbWsf88KFKJqxkWu1g+HRz
WOg3cpMVIjT7ZOCJ7p61DvP2fSSoG7JoD6kkLRzXeX0n/kCgD7Vyy0sPKUoKfOpl0+bkgGqvVY70
MX5f06s7o9S8/6mVcrAJeBM5J+ZwjjiJauEbOqMVTiADro8jJh/m4lD/KoPXUOyFdtBQEEWrVnVk
2q67/EhBghIsvFpKLFio5pKwPjSaP2GKVWOx6UyKPqOI8/D2Zd6xVblkdOZNXvBBgs2rMpZCDSAR
8dNE/77VbsunlutcGdTlNWX1U7ylnrqUiFt9eeZ0xlvEietsBcC54dQ9ROw8c95QSmLTHdknLgiY
Q7uEDSZYWFV3qmUcVmNYP/yIoY5G4K+7RRqIIWr3F9yDRzAbV0AeOXcSQx74/8xGFtR4sVbMOd1Y
1jZLqpYuYHQxXoRp9w3HJqMeRX5Ec+9/R9ZmpexrmJsHgdxRmKDyVg1225FZfmY9O4Cw7aFCYJDD
r7VU2p08DB7bsc14TKy36/2/msWc5lZr4EeDH20ySGbekCYrI0mvyCWuAdDSy2yEN9sI39sODHVb
PgGCG70MoOmPJkKAXbn1h/KM2/ZZPMY3W6jD+sACulsN8HYn4QeEP79Y5SKkD25SFUpGZmH4vNog
ut1Ngc8dfTBLqsMq43u8UZDIbL3gSyBocboc2f6UbcVxsSsJBY9v2KSpVFwM4glH3JELDcFqaNQb
pFVzsDpuAk0wUOf9UIWf5dmqDAsPx86McmxdxYfs9ZGVOr6N+3n+Zf3ZRo8Hqcbhd8Atl7/VHAkA
cA2/lHUSgoa1L8C/j/5tcvy7cozrTxtUY6Sf+//P33qrRAuRtb0nWRggbuNFvBcWs5ncn5tOfsMg
FyPS81u1HXVlMjzC7KuqEBVbLPxrhkFyYe4LmSX1yyP6X7KYUG15ac43J1oGoACOdN7DDHz4+9uo
gLjT3g0HWR+xkgcmtVcItHggz974aJpXxzmeCvd2WpyCDePTEDm0gRagLE5A9Fii7PKWf0SK0wZ0
TX82CiyzE9j3F4aAF93I4yWMjCfEAwIn4sdfLm5gAmyu1xdxVYn3sXKvQP384MdkbRDYes2HVyPX
qnY4oxWy0sGeaeBsFm4j6HR4UFsmmze3VgK9CXpCFbnfHDaVPr1wOaLO55N2ZiG2d3O3SxNVZOA+
75qhqwaCaxiCy3KavuMlOoNh4lRJYEHFigAJD1+qyNhGY6golLSBFYDa8qKIpb4gRDSoGXDeHjUL
mD8PdW4Ev/tFpIV5tRmR3o+FlM9mXt/wWscwTJy8GdHogucWo1A1nhMaUOFBoXL/h9C+q+FzuJs7
AA6JiRqu/tf3FnJ1OCi+XAj6fGicYDGt6V5zMUlwDnaw1tqAg6S6U2xtuCgtsq3VuqehWQXtNNQA
nqunv8amG3jQb4dmOJG2wbtWCMJPU6fyG0fApk2H584Dabn0iXiKXEr7ws4PB1xm5N6pxVxdT0fi
nLSZCtk1kPBTLAV0pdK9UD4T4f5xE/kJ8yFrwG21pWss+/+JAQx29rPeTTRPdB+K2Vc3HN0fWZOU
ymiWfzgZkyLxYzTRdR4d9hrTtVIbx29whFI/1k+At0DCGt/YCAvo/+PVNgUhbQaAAXYYAdY8O0Xk
DETINR6tsqonQ+jWwAzya2mTks+Y7UTPqWn6J7jdja3S8EAQ8gz7khBQHmR8wepeWiTNeZzsVe8r
+nPuTWd35azTUU0LdGfHOqKkFxdNsH5M5Tz5fHMgoJVAKRzT5HdPlMn8FiqsMPN+Le2zBlvEZFk8
CHhHsbeAWEUmVLa4P8FKnQt3AqpdVZhAi9VNSeuEac0Y+9fTu77l2eVCJ4qepdD+PasY3Z5xXF65
KxH5Brl3AC//5jP7ONm+GGO6cYQQcE1f9Dao9JkWJuGe765Yv/P73fw1PjvYVu8leWUXQ+gc37PY
oh2RF1DMGb5ScocfD2bOlnRjAlH+xlVD0TizClDOQ7jjazyLlrQYX2quXzHMXRm7cgsjDJBPD7IU
P+8F0AbI06O7PWo32lDpPQHh7x9iuo/jpxDSYMQVfIlrcLCnOhXgawnjXzLkxS6wVwnOzCFsMbrp
HZbetfx/ZOOQcVo5UtfKhKdPvagLbGSC1moNagkWzMG3pxia46q/g03NTjGp2VAqEWbBsz9yiT/A
OC06zXu5tCYvfjZTT8AOt7bInPYWOOyGrkUf4byGKZHfBUIUUi/PKw+DYHCpEmC+KzSH4ovjsb9j
6VpC4QalhGnhOBgqHFYOtKVuHfK5Qr9T36uRDcQLhlGh18+q+R8d+7D2s72TNdZujJNXlmehn1q1
jlM6qzZDBu5JJfvpg/H0/P9EmoBGQleOai9e37xVuP0TctyP5JvAOyj9aA28TgMl2fjYuYK24pr7
8q0W3L2gyuprrBcFKYisAaqQCcSXKKJp35Ia1QZz7y0ZYks9yeEL86JDmEuwFMZrXWLHEm5EG7UG
KXbs/+g0WoEDz5V/cp6BV/Jgob+GbyTf5EYcbXgRXhUt5DckZo6B24BN72OGA/6kiQUDXMrkVCy6
EEfAioiij6l/cpA2YDEP9xlc3mzGNbHZxjh7ZEShOB2r27ry338WHEqdfy4UkjrEEp+fr++nUKuq
OfJGX/4Yc4RmhT93YpLqY2cgTB/mGOOn7j6lEL+veaQFaqgGIrb7HOWuNFVLdktMIKzXPdtW389x
QJNESU8UIfchSIi7wYKh2AEZ6nGAPmG5vClFIUyChU668UHDIfSeNtzBEuL+M7xG5m7/SZcD1JYY
NhXMXMQjgU4ZqrUeWV6OLr3GJt5/I2RKo4TM8D9HvW1y/XIG4k4WDXHZ4ufrtSYH5ZfsXnnzMZhk
HrhOMKsBMtgS+jmj+CJfffMWh89ICmEpSmpOj1Ktr1IdMkdIwr57hKTUHcz3qXuI/TcOoj0dF1mW
+Ck2mg7TP2UPwqONqfZR6+l9j80OYL5r539k4G1CH9rMRq0ElbgpCu+mKd5osXbMCOryQT7tDWyt
6OGXp1nplH1hKT125iu+yZ0qAu9BZt7q9+0y3Jle8der5gwzKXb5GadrnwNM0yjwGercxTAFJViN
9UZzNqo8y8hpqRyhjYX//l4RmMsmcvWSQ8fSYY0HFlVG0Y7AS8qjP2WhkNcoFwyQFN/B/ApMMiJT
JyHEyNPwpvQ/fa/2JE2hWo78c5dLLRPZAyKOhEON1u04BCKOPXvD3H6OLX5ndcaj0EnMmSxmyL+r
LpudYUgo1KU9WWYpSgLPFK6LoE3gpJQXoJl5wcsKsaYwML/C8UYvGGCX6iMOB24a2MaegDPSuj6U
O9bW7zTjR34K5RO77HsitQKab522Ezzr93aWaxM8Qa2HDbJZPLrXctJnuupFy8ouJHi7eg5fyTUe
4Y8j6jrrwilrxAmAuazF7p/Nq3f7RqxSj5UTyu/k64t6Xj0eBfIjFajYgzPIUZ0mRPQ2yfssuE3B
sx4q3+95UkU1vX2icKjyQRtkoO8hsZb+7UfRXdN1c4edPa9OljCHVzL3k9LeVBJk82EvYrV7mJVD
KgEnKWP0DOUFaeGmbt/UUzQmi9jNk2Yd0j/b/9gAyHBglz+wWogbshHBGJIUXua5ZqfTVyexj3SQ
XWRyQna0enevCO14SGTQft+w3dE0xLnjhvh1OncBkG2M+XsWNEVjs54yWAanrC7K7ePqErWXKRnv
T1NQXhDE6qwU/GIeEyGdWitqv5X3WSAfYbj6u0RCisIx3B5ny/R8OiQXVBaI0NY2EqHku59Zb9Q4
4pv8m3Sghbq7SyTBtL6A/5tK0ZTk9MgUoTAI0uBC3TLmCuh4safHjUenwsx9Mneu4gEqV+RA1deK
+b2XCGeDP9utN5nR1ElHPyiDS0B8qEWWZc0vRVizvl6AFnLZICSaGnqith9MvNC4nuXqQtX0gHjC
92FD5S2N+11Xm4Xc9sZ7ho/ZYhElnCEyLDNQcaLVStsYS+7S2bVDQ60DCppfROLpIHbiZTdJCAhT
nJZIwPbUVY7M/xogJZB04WObYDTZIjOcsviPH2XMj9xu+UQzX0yvgCBrs7+hfmb/VLmfrhIBvqip
Lqa6AWJ/fH1EtMAow/wcroWIkTahbe1MB8ctuX3Q6BnOwSvLfEuPOPQncmt6fAa5jAkLgs3F5EZo
17478RKWJKF9g3tNbmlR5xV/6EcfNRewGotzjOt9DIPAh+CuUpktnI9dLVws/2lkpUtDnhLsQM56
GLxTQIaD8Nuqdn4doU9RpBbsEl36sTJbPNLQLpL4j8J/lI9FurMnTzt2+rOBJhpZMK6DD6vx1zJm
AjZqefj+om0tmP0E7ZX12IARsTjJydCdbFxJBL9K9y4YB0k3NYad8NTILLWJDEVDDoyBdSpmznVY
0qFyd28QLlYKU7z9avJZ05Z3lcZ3pmwoJv72jWJ68Y+rUL0OayzfVNmK3zbloCW+mSI/NS5zzpFk
7+P9j7cIzceFNktE60lQYHkjXb1t+FugPdqeWKhpexZdmq7lDul1gwfS5JTXW0bip/vYPUvipEbi
CZbnh9I4zt8+tSbHU/xFFc8h/Rdu124RocTsbvwUTwc4wJSej6MdZhsyo/q1rxuQaGXATxjTq57Z
jZPBHgsQvKlWHLiSmGia0PvbcjH7pBnp5kMSNhL3GO2v5clt91P9J/CslMlt+AdhCRgnUQg4SkLw
Ec2aazTFfnAgpabCkUUxpi0VXVjgzsJPVkMwrZMVjEtUlOJ/TEwo8oL4CGbNydfCYpz+wB7o1/uk
ZSgfY9eUDykeTNVUrq/yIAH+lFfDDZM2cHTZoi/5iQ+8R9JIrb/fjyBrSrLI0t7FhwIOi9zKO9ar
my8CuuO0IcD5b/C7m/AN8Yvss82RNiSalKNUHh9nIQnEcOH28znj2a4+Y8Myt0Q38LgXdtzsXO2P
qs0iH1pBlbixY//i+ocgUWts1t6kXW7vbPtBnshGImTEgi1PKUVJ0Zy/GIUP+4RMiRmyh4RxsGvl
wHNY3tEnUVb/ONeN3gkPPRNmGW/FoQQDjnVONvAh3iYwI8efVditz31DQGzXq6AM6SqLue6mo6cN
C6N6VwVoDKpIQ3gfMypV0zUA6zuahYnuznWto2VzxPxMg3FZ+Eyy4Jl6RnTjXYyrcWzocKvSoojS
7ZH9REkQxoPHt7nL149JLMOV+7WP9hSCqG/ZIhzbJiurnsvRH5GntEVh7HWxPcVm18bPyBQSFZhY
a5DSO5ABnNQPf4mYK+iIKU4JGz2a1Eg864lU7+s9YUdgzjAM5+64Z7j+ODT1NquXDmfIUE1Gb1GY
7K9vfPmNPxWcLc/wAoIhICUUy+FJlMGJgZawzR0BSmluVcITeiwXgubXiOYK1ww7EUg7GXSL7S3i
MGryfvmxee8Ouc4Izq4nvRqnujCic7PUHgulQ8r7N7yKWb5sSC+q3CDLzgOHfS+Vr8uUC+2THQoe
WvtlMCFyyJ/wCpZfV4tDL5vrVzsBo8kNBDzHItYYryOJP4pvZ89Mye8MefryttQ3Wjc/RadG1m4b
ddQy1Ak+XspSESaV0paQvKeqiPNePG5yEFyPX7Vhyh4HSa+PybytsnrV8OWbhyiGZ27Fe9PsZkzh
zuj2xFowB+dkd33vjCAK7pIajf14R5SMk0ImDFVx42KPHLxYd9zVg5f09uJj+vczw5VL/KnKnXLZ
xxoZxqSMhcMJZC0O6YeiL7ZHo+ZKA9P9IgRGxejKtpZsA0AaHAqECtQeRlduw+7nz76QeuTwf0AQ
OUiPDYBfaawP8yvZhMn4faYR5bR+vK79AZewpNjBxWDNDC9eHS2HglOgYT05NOyftE+2Px0cDVGe
W1Dm7byJMYQ0xrN5fnNWe7FFRk9nKj3BrYgE3+vaDLjAvebqOAcUqTSW5Cf4Xmorqg9VtQNmxqx0
ldgkQEMpWn9HcDAMExRM9xvEaS2NohqQZkmvNkel4k3mB2E4rR27aUue5v3fuzxrH4oSkD5xH16q
M1cdWwJB1x5q0yHMpDe44GC2XYozxvf/LmKhkYnFHjgmmm73U+tta7i9pIV5mlwz8Sidk4/LuzvC
/jIXh20fVJT9euOUHF4BzrDE/euzRcOK459MeZ9mBk0oMlb7Hf9mi/+iNGoPyg7xr1zJ2USHkdlv
ikQLETAC88EZOk3Xs82A6JSbszdbRN6ZD51fKyIPMZw+md4J9xfTgFWjv3Fn/UDJveueLoHcvlqU
Q3s8xXyuM7X50TS/vgJXKWwcOnjg9oBKCJoQY3S3kqJugt7HBcE7kG+rNpm9qw0VLw7jpgI34izt
yC2BotjOwF87aXQkeyi37NPSwXVOu3XGoxpaEIMJb9+Wclz2ZR1lU1qct0L3JV8OyTeugEz1zOj3
mFvQ9lZgeLJFW2Cr/Fp49RGyZGd4haC4jH2AS/KVTiBrx1KgcRxM+rQyJwoTVUSKWGsj6vLslpTG
xDU3Qh8y1JorC0FgK1EKWEHhaelLtK4t/RXJrjVh6l5V3m4FXrUdYMT25x+KTKDCE3ginVx+7Jwh
D+QagpeM7izGud1vHEnVRQpUfB9e7e1RB2QUnHVmENQMwvoGgphl3VgdAGTmpS7LPeiJ1awYql5Z
8gr3sc0eglFpsb6Duu5ERJ545Il5jyS0YHfrkqwkeywFcdzQpaI9cFafJy4QmYT6Q69l9QoqI0NZ
CTHzNUB1378wkS7lMbORq5pKcwTtjMzrbcAdlMezCaM72/wn6pVFewEHehGU/mWuBPhCs7DPXyHJ
Fipf3p8jJo3Sty8PhStlzB45zRjaeUuezNKga2RWj/pdcekgVWONDfel+Yvd4HlvkyaBzh1lpFM7
mdZpmkGmEZDQG05ZvIHghl3UcN3lrjULoxcDNFRpdlXlip1ybFoKQpm2ijlUNOm9iBAtMYcoGJAw
eacJhifoG7ZawEw81UnrD7M3FjYoVyb4tT3g7zBELDT6GK2ewAUVQfvipQyjnQTrBR8a5d8+oXJq
kKTK7tdItNV6UmjyQWHLLV160DioF5h0/9PQOOL7ebrXT1K0JR0XxVAoX6hiPcq9lDQ9IWUaoI0X
0uJMHejOLHE6dppCkH0qZyLb4yLKHMEWv9bIfeA8JuxwPd6nszV3w/r1pZr+PmKWNGsBd88XQTty
KeeagcooZfcvj3l9fWKqnswYHiM8TKreaLxI+Zpq5VxqdYpU6ee1aMSRti3OUJYSDh7c+YsDN2yL
gIApe89OS85iXHI6VzbLnyLXPj4xJ5ApkXesYy3LzJlDi6LWTDGM8/2GnDHEohPlD8vcxYFENa4m
z2OvyY7z9//jNrWrXKk0aRa2sRzuE17JYhzGsNM0oanNzrIP+u32Gy/M5aOTOli1JWDPjhB2qsFk
WsFw7IspGSIgFN5z0qvstCZKaM5WHyeF6suyyxn9dojQ9+GXTcK3YbpCWHhfRMtTeBoSklFhBCR3
c+pDDkJX+X8Mmb8vnczvJfUzrNjVUnZZa6LBAx/886HqCHlnhxGLbvYHTAGJIP50w/ys+MaBIDry
YAReFUf+Unn8KKycBvIU4nLPYpraV/A4LAIro83EVDvFWoXQH4qpM5NdmxYj6sI8b8Gg4NxufIRG
4bL6bniSJ42S1Bcn6/32kuCOZZVzLVycS7syulcW305iS0NQiJl/ZbKpxetKGPlhFv2+emb2olp5
jbPECST4dcjrHVTiqjrs6oaKy4hrBHysRkpooSvza8nFBoEsLcGd/CJ14vv6zZ/il2QBi9zCgXcL
gvAeZlhhPkWMHGcFhbcI07V3Cau9U8AaDB11EJukq/YAFh5EpDIyepJoSC2+g5RieTL3nV2Qk0vb
d6uFfC9rVWFLPB+NiTJRdA97mSaecQzXHa6oTK1ejAX87b7u85AH7vETZ3ksFfG5BPX9fJQDhllg
UccdYVrCMyYWPZDlxNfvB/yKIXSPba9AltwnHkxVuVaM6GEdt0hceO8a0lXaPdBp02nwZ5IFZaOy
mDf0vexCxbxgBTzhMu/xaaKZnPzoXH5GuHbI1xSvvicVuVlhB+4Qj3TvtP3jFyo8wxB9qmOJRnv/
93ePRAJvZaJgwDa7WQFcD85tr+D8DrK1cwm0k0ukUyw6rwvB5KSj8/CTd9Z5UO+clKPtQIOMcNQN
QJS7nVL8w9e45k39BVK5wfsNLzQoOXvcbEgQhjc3/XpdmIj16It0L7AvtXP0aehbXS4wEgaqOlua
flJn7BT1hvY6yEb9uap9KttQ6xj7O+0L+wPlrMgL9nMBJZsyX1ObRX6QcBNH2eEJWmi4BzuVal4L
G6aK2/uKrcl8wDyFNzgADMce/6ikUupmgEb9Kc4RTQBEZMNVxmRo0xXsBh6vjLOUAfvaAh8o5mEK
C6Ef019gnQkjpaQdg5yeHiIDNWJOM7bjR9+cwRjhHcPHeC8gI7txgGrzrQaBs+92swKUWCVROV9K
MTuvQS7Xurym2c1xiX87Aya4no8r0FVypm79SWA/5yPSYQy4b3rUeuIutG7Pw0wx8k/fT21r4W2H
ReMZkxL2YRlK5eyPISpzf8KReEZEfnrwcC78joSyUgCMKSIXk7GQoxxLV6Pas2OBGdZl+BDIdkxr
/IxOiohUO/Z9RkUpkA+pIPRbUrGTbE3R+C3ZkT8z9sPVTPMCqSwzIRTdcL9eLLD+FYxLz+Pxpf9S
lRtMqOgmkevqh5iKz67HPXhQUYNQ0iB6y2dWZJpnE7kN8xy+mvynt0lolAmEr3n2RP77HfvZENcD
wPCPGiHNHwi3syJLTAxV4PVKelv8sO5qiD6ZAO3ABLEwcOQ/YDYHxHjo0VfmKNwDHqlpXw1BMVe+
tDGrDuUeG8f/CSv0SYbJGLp+8HVA6flFtbQGVeCEcovM/NzFAW93tVwVCuKJsI8CAZluI3cV1U02
CUbbLI/yODWe+5QvynGRJUBkClBMpPuyOiIkLFyJFIfQZwd8fjy1tqRT5BDW6Pbk31JfETMrL6M6
mB0ekD3ph1k6DEbLOD+qmmuE1aIWXGJwH1X5P0TMIGgyYWo/JDGxn1b4UjOgwOmrI2AWyMJmel3x
Xnq+BJo20lxgStYIjHk+xayQqRpek1j/rp+D/CF5ssY9sJGeQr+3sPJRxUqhYcJSOVV2rEl+SfGq
a/wx9Z4lfsf3mX7zDFYv3BymzhxDlnkH/CI3Ja68DH12hLVlufnlvK4wAhZIENT+QH15jicoMBOl
N8iSBPVPQWxZQxgJitfrvvnOTebufWjy1Tns4SlBbkeJZkEZH3C0Que9d6okRYqcW8884ei5UOp4
z79PoWyLEni04YNzNP+x1NWQ5Ei5hig8vehT341Vc0vnF5Epetwpyiq18ffmJjaEgPCUZvgP6M6K
KdXkW3sp9QesX47MQ98r5z7AXJlP0+xP8XfcEkzmCBJSo1yvf/gbY4MKb75Xn087MfcQejeMieR9
Ef3YCSOGKu0xen2jvKd94tHvRih/qUGYDbOnGdZf13chwb1gOnOsHY798YyJQU3vpBzbct7ohliG
xu950pv+WEbZ7ad86GpaCnFGxNGT6ypRG1feR7d8uIXs/4ReZ7LapVeWJP+lhJPU0MO1PedwQI2z
d53lIdnlZx82O7/MFiQ3F+iMpsRwSnpX84O+hI2wDviEoihp80UgEueShAc5W/XGh5JQ/443jX7O
6JXcLchkRmNamkF4rFSlNxqmi1MNrcrcCI6gifBskfXGdrmfHmJ0PNeTO66NzvfiOtc68tzgEroM
ZcNxw3ziqagFDJDbSP5Hr/1dbVoWKvUdrhe4TItXqqWdf5CDVfmI5n/AcG1heJYk32LpRE/QoOwS
DwdV5NX3Aojf5BRIBEWd9unwjdF9kbWbV6jSC2w7UEIVtBlqn/+Y1+WleFb+Urcd2F78ALCRkLWG
h90amwgoqJZw9Tlb+Hzgs5IrGr9YwQRTPY3107cB9YHkoVINOE2Io3D610mxxIdhG4QrApM+B3/h
ZjN3XQaHv5NcKYr+jRavOSl9DNlYQEeoAUv4J5Ufv2ehaoLvNVtskf7qFtGqOKVyE0e4n2hgl0uV
Cf2pqzl63W2hwjurvhCAhiwYgs7HYoWmzChftj/FI4Cby5lBedjVNS4rSx78uvJxdjanljE0HHIV
G09CJyqnEB2TKpKSJQFZHR3g9Wg1X18txuE9t1fEsZHUFfcFATBg0kArGAOWYhHqzwxJewMKg0A1
9lspdOx+kGYYI0Hd2W3to9OPFkZZ8fVGXsuh/WzCrQMqMMWrAOIhSAKsO1wJEWSnA8dRA9Fyl9Vp
+z/uhcN6gAKKGLyWiq8IiKNrV3mbf6aoFc8uCh4mbdUoNDl5pXDbP6rkc58bgklg3/WmUbMKnxPA
ehaEqVxt3nRvbaiTAUVabTr11rXvwvxiXZqwXrYC4lgwhKED1FOBKV2mOIOmdSwo4xnRNORhundc
WGGymw9v2A6Cr3/JJ/3L7UbaCyal0ClFdRkSZ+JqypFDV3+CUOlgwBDAneAAP3XURYqstXgAlw7M
FodTGMWt8f26Z0rDHzzzn4Yuj75XYG9txVbO8s6/7Kd3Op4Cu8YNvOD+hDfwqXf1/S0tIxZZ+e7t
Fz7VlfM9SriOn07CwThaPE1FPIkqbxz2NUKvMbOlbCV2i7RxABCcshZubOsSpUEk+8dR0pY5NMeW
8tSDMAUPdXJSGdaqXOo7bv7AGvBKEaJZDtB9XLfGDGYRSluJ0Yv7hh7jr2nEnT1R8gGy6kV+YYn4
tOg4Y3GyQU/5eeknRLiY5PjyUXrFrMmqAbu3HEud2/fx5sO068fxAtUrioXwMYlSZTixu7zoOGoP
Nc6r0aJEocuKADrvgu93TDwNP8f9ZyL3nREW3HKz+ZyX2vgZQPDk9SCmx6zbbe4YQiplGvdek5n+
cX6tUURXCgwzOX1Dj7KbcWfHnsb/pkexsuJhZFn470uyGUR22hqLuTzlLJ88rW3TfnYL45cFmcBC
vXLDKQzr1+rSchf2Uq2AQaMhQ8gXe+xDRHjnJzX4BaHkxdk2olBxZFwSRAKD2z+m5gG0/Bwc+NNg
zEL+4TUuGkQIfJXfhDaga01VN7JVJFbLjT0dn+Ksz/3xYZ5jdNrC/dSlwcJHcHD2KwHeLVAhtz1h
18QnM1p6dl/ubhhdmeIK6i1Ufk3SYZkeGQQgh96XzdeqZ/zhIy4DH6+VxOJbk5EElVfjZ2rx7fOK
No/nCIY+5qHCp3c0ZNvRXgvc8z9DVGeGFsfByfLnSw00ss4LIMLFL3tXuvYskIY13tQuaKnDUWZA
B5Qo81EJQb8nm6hpZr33cmxeHocBpH33wMwUHbaDN1J2nNpwqeZ5VIXvLO+aFdqkoUjhGlREwnkm
5CGwPD/8UxKej2s3bKPKAimlNbUqvB2p/+2v84MibupRP11kfMX0kKlQrafxqbWxGG67M+94eMpv
pmhY5p3+zH2gXZlU9tTebusIXsRVaOosUen9nx+U/5AX5ZiY8WStdMJol4I0iaTnVZ1Zu39x4nGu
YIw+b3EiMiKNG75zzr7LwGmnZjJUT3L5S7rvTtiHBsh0Wvr8GAgfoX37aMo8H+NniGiHdsJPZfUe
ieou1LOmJp3aVHEvH0WYf6O3TSlPNUt+z8JObgLNzBMRM3Q3+bDUsFjhfu8BRauPuuOauSw9V1qj
agnszIMq1MUB4MUkxTIfdUCPvxRO8Zw71rnbC9dnNns0nDbbu2l8RBjvmnDHnkpvPFEVqmTWpUhv
2jyO3tiaUzOCg2gVVrNx+T6cYhJUaPs1fo6XKtk2wSg5EstPnrCDDYRqQsGXr95/+vW82Y5S6db6
r9ruOPNar3xE7cbrvyE3c4pcpIW48XKBbOE5zkGY4jfGaPWghiPyXUDQNxm3ooGLlIS7r9mlZX8x
Udmx6XsT8khyVsL3H+aggcSL7Y6OYDmQkLoW7nSrn4zwptEe8Q4QcM0n6EOJ9T3paBnJEoO+9meA
LNabRTEnM1RjNsPVqkTKJO9yO8donHULW1duK7Qx9XOK+HD47NzCzDNP60W5a4fBvhzvx17UOS5g
4juQP7co0/vXcq2Mp+5FVo1FQLFjsYIPeZCyVcgPI8LiwdxZE5WCScq9wsDZ/xFevjv8H5uwpqAw
mWMruiD61XBIT6mMCMJ/KH926YIPfXiu+/IaZFYIeZt0ZZ8xBNkzPUCyVlDIBEhcoBsCCNZOzeZk
lugZdPGJcJ/N3IiLMAbgIAPiFyL6uY/uesfeaVufyiYzMZSuCluykJdies+5RPZYITIIhbaYbLjK
xMN2Q5VwRFbWb1NfZz0pfduw436wGD+oTJSaA5EwloXV+bOXep/URq9dn1ONJJuqpKwV5JSgrswa
cSLOXnreXyf6UuGLQJYKEemi5gofQALo4/wuuozakAmKYY010KMjD/ePa2AqWmuZ0JGklTvKUFdy
3uOhO+1Le1Bwuf52r3XxT28uRIYeH77Wq4ixNeClqOtzyEQsj8/NX9In95HmEyKl+do5AxJKc56b
aNd+2xSuFSB/fA79VxypR8TCaEL9lMYyTkywsw7j1kj/4nQQGv0EvopIhVZJsF+TmbMzS0tc99rB
ao7xIJjSR+17RoIXNFK/Et5E+z5Z5L4kx9PqbqcxWQmpvh5YlSNfsPvJy3twDxbw3E0X6HZpF8N9
Yav84i7hBOOmjsk0nQmcXABb9A48MEEmHWm3/mVt91G+N60Hlb8wzx14TS0hzRV0yPu6d660QbcP
E7WRKbtsmR6LeGRlBsHfyZHKsyHBC8RNRTob43Y+fW+iSDedgKG+S/6NJP5e79QV7eX4Azmzf2b8
0haZt39NX9SeTNv5LpwJ42nOFulNihncy0W09Irin3FiNlSEjhaXdKaPaDRAcDTo7ZwiTTs9OlzP
K4gQPwg3o63hEeNX2OdcDDAUHpP5TVzmvsTHjJi6BNGeDxvMAxPdzqmPL/YHZbR3ApsDnKP6Q9uy
GdCR70rBKI84Dz31g1CqVg4JuXNd9pbtUxGsBCJP++A80ohtBilQzFsUsg2SXKpeVcPfUAajWmzg
sZ3o8YZjLupMpzdtI+mAsNQVVAxtemB64O26ykHrf8I7+9bv+X07Zx4uf93WBn0OhVEzqH+ZMfMX
yM/CYgcEbO0V0C/q0wQlG82VnmdgMsZ1Mp0sY5hpCic5JJsANlSrYlSHBNbpMp7p7w2GD4gti8Q1
UPlu3O4J0wAzQLtYqmFXdfguLpbwThC/yhc6uVhog+yybNIdBb3Oxc8AmaUUM7BVRNaazQ0P7hal
YtGYhLOjETxKyjQDketjx1ugwnLavg+H4l+s9QyM3joWeNcgmMewaXHedNmcXKizLPwe273A11LF
lOYj1ThXjzfVxQ17A9pe4wCGAulsnEgHNt2vdyNmu6jWmJVY7n2QV9HK4XdqEeshSzhDLFwFXG5a
joUR28ZjbmxPhmJYgQ5aLMwGS/TinFjKEhfdLAxni8V0MiuEMW8W0n2PI0eBQG2P32bf8kWX/TC8
SJK0OvgOO4Xwsl+iqL9NdYvIegnG+7zdb36R7tyDxSqoUru+QKHlMRFt5IlXZKEJy3VUxlUcO9c4
iTuCjj9+gZSjEPx8wKgmwOPTPviDSBmwV5mZigd77GftUfaaa/QzOpVwfQ12cMbbvXja8Rd/C/7z
slQDeMmOQ6AcosE9nXAfUvpVNDe5aiY2xez6gq7eTFgx/4hFZ2c8S3ThHTCPW//ISyCeq3RRq1Gv
IRZlSgxIzu2dYs2wvsWawnTyraUHHlPRZ5D7cGWvvv7fmpUD3lSfqVaf1/e3MaMC+yC4Hnoqy4J+
cX+YL16d7lUokAv5KEpDfc7Lz78PhWw4Sbmw9wBsE8d/r07wpIgRgx7z4TJ/A0wRVUb6IchVZasv
VJF0UgxSa3QPVAUpjm804bHcCSu0oT3XjfPi2ViVzDG2It43tBw3bzfH3Bmkhd4ZBrB/SMv/A4+2
RvZcy2sMhcdyToqNCQnlx9BMxVPSpV4r1nJsMCPcpfE3ulzk8ZyZnaytPNEzkiW7T3UJIoWgDoE8
wTbhRw9ZrFZWBka8ISbj3C49HggLF1GwxeEUvOh1vchqeUxiskDA7FtOaLDyT6uV8bERERvKm6sQ
rJ6c2an6OPo7iIHH/937+HvnTPry/4TrMsg2OnaID1lziGpAcXUmee73l2rNdfLGZjnNogdIpb+t
jiD5aN15M5XRH1USWS9Z3KfTuIoZm8K1EKx5Yg/295vLx100PimL1e7CaG4DVmlEfl5cPLBSjsUW
KvoLIA4WB5iHig6rL/sB1Bpb8ttXhQtCMWzxRXhcYLGfHf+9htlX5YkEDgsNHoWoBj3Q/7HlL03i
3KDmxA0o5e0PpQ/t86zQ+lXguvO5uUWLnjzVZOrdEhfuq3FewAC0EAA4qcqRKLXBFwXuMSSrNraq
DDfKw2dSBVCX3jAekLV+vchyo8u6U7QQyaPeVfpLKUTGtruVSnPh/DjpRfNaSkHanQenVsT0e7+F
BoCttDRN4kPU96fWVBlge5l9HwpC3Y0hnZBB4Q72fIaQZBRzbq4Tna9OEwmT5nU3kq7C3L87sWN1
UWV2jxYhJdfZWepvj7yUmCEyytnGquNoHdVk1o3jSquHKQm1k9BK8/j2HF0XDGOeQS/OdA2cWEKe
3LuPICbuQEvbg18vzx1oXVgYqfY6Gois9bU1bDiCthJbkAKr0ISihTY6qVaQRKME0WnJRuojgRan
iU3izSv5OPUaP90r6IEGU1j8tGGPApY+VKGUyFPpErt0e1fzYTcYkFoJ7lhzN0+QfTaWtD5A7KGj
cSLoMVVuwfxNXDkTmmmlgjRd9B/4MoEdGy2fdzaZGzdacd908NcFxGCOx7WErfXFQJdFrpcOfmZM
8JH6PJmRz/EZTfpdavEL3slmvBsaJOqsmGRgnoPLulkfivH3Lyq8lvTLnMHblEGDo4jv4J8WP7P2
l2viiYS6u9cO6mwfnyvyE0Px/cteayA8+fAotmTQ1m/OKZCCSaTVb+aNQLrpD+rykAiYisRMNIZG
7CwRZgIxxSJ/rqu72e4Kbr9dw0Ju53V9MJbAnDLZ5RIfK54npKNFp2UgaNuFIshd5sqRV0ERp7B/
M0BqUnoLZt5IgMCWuKykdv+JF2lQMpfOsR8Kn6VEWlNDgPl8rV7SX6Vz8Ac4Bkih1B7CEoZypSIv
Ha14K6NlWgS0tKxb0eL+NQS0WNtHByV1ePlQBxEUBUAhW8Dec4klM7ToBRfpYnnrgsqLxxBn0CWq
OPMMEdmUYOv2BsWMT7zt5kUBiV1L9sb+OGBOuuqwTfdf5QS649GqyekRV1fptYeGWhc1K5qr6SqE
wYCetiq5kJyJf/XI/lN1bZgp/IY5Nb+vs0X9QHA5GbZrYRwdK7c+FOL4YP33UbJr0Mp3Jpm/p/Pw
FX9Ptl3hF+oM9nifD8JyOFY5SiY2OH6GHJo9naCtHURuvdXaixz4Wwa0SZEmjXELYPdAF7J3f8ao
7yAoYZzgO09r9TFxJqgDskyyyaJdrtw0hWl8Y0vkTujOb5wtPLZ7wrDQn58WlrzlgXlCIDL/QPPV
w9/5mVchzGwZf57CV12SQ2X4vTb97KjSxkA6C10FJnOToBh0CmyjhpkHosw11jGsoouXpmmos4sq
VsBKL8VdeEIDh6qMVXrYRnci0rPVKXYulu4IptzzmreT8kBCYdA6Wq+E7jDPzpNAmZD5Nop+iKnv
Lmi9OZk3yoevmWvWMMrbp0sONCTkRPIitWjqcccoMKguQ60Fztk7J9G30nWFt28FRQzdWBR7FKwH
FMSEWiNSVaSuu+kG5StvaIrk4dI+xO37HXI8KmPxFVVhBFVWGcGMXMGEe4SYODoTl5mxZET4/n02
I+kigFTHIKpsFbLn/aYxLBeQg8AYhu2C0qHriSBCsteMZ/s0Y/AwMyt7TITlMHajKi2a7FLn1+Mc
4gfunD8e2GrDhSNjUBrGnRTJ6iKc9BYLj76Tw8+RSKu8KRFY0PQc1bb8jt91ab9mlwEAYmbNfmBL
JQrv/njgXsjvj2PwewUcwxklDuIoB0JQN9cg0jrkrr2vvAs57vAi68JLi8cUs8VaHasZRpySWlHj
FELw5+gm5w/TX2rfq3VJMY0vQ3QEYo0DYiU4CbYnXSMGGn7c0GY6ALCc0jwYUaH9n7ggVBWb61Un
ndQHd9C2/OLxPd9zS8hbEbExCG0nxq/dtMwhESTRVfFcSGX45bmMMgJp/QL5VdSP/e4ojYkL9XH3
Lkl7JLzsY5rjvBVDR8/uoAFpeSW1cr/5C4NalLGwtngx6ryxnuMLm2dY9JCxLQemtAuS9cBilqmN
q3Iq7yyoX+0/B4xXCsxT4eTaozMEmA0fWRfINEghmbt28Lb74E0YY70QIgdLrwt7jiOx5X3tZegJ
3X7c8o8AVEbz0JUVsheKQp5AHgrC6chAM5eXV/ryNHa9VmaH2e7Q6NolZkbp6vIwFSSKsSpOKS6G
9T6K61oaazT3XWgVxlRCK7aK2j3muQeVh4OwMN1eVIwUxbu9Rj6LBeyAIooTkyriE5m4GEF4RVr4
AV5k6G1XAfnLQ8jOWuBq8PJ+/OdhAeSbfuAe+bdTOdZP/24gw+dKfiV6o+dXoTjiE2nPXN4tOx3n
4cU2ssvf50ZWh9jd4ZpfvbpH+DfMgfviOYBC2mz2igflz0G5drNVBijB2bGhxIMbSiPEv+NB5SEt
P2kxVw2AuO6cU8V5vJgho/6wtGkB8+x2v8IjwR6+s1dMC49cCb+cm+22akerVkqpOe/wAb0n3nR1
rMeBMzDEGH3OVkMAHpw2h0CujFdJ/MgybZqgZCWTpzuG+TWzsb2wralpUSTqIsGvymaKmF1OEv0L
ZzSreWX2siyF/IpW9/iFvnqvApDuUMO8icQCD9aYr9LUP7J8ql+sOSa7Chy8OdUJ+t6NwzLVjXdf
v66bFCLm9AI3I3au8TWBQF2bTZrnZ0DUWNFVvsQjqehoC8Fwpt3M4rPja9TvcCRkqEQfUDtravfp
2dDCvLCpX43urTHIvp484h+XHwh97YhxXTVqJJH9xWKmsqL8aJYUjE3iLfoxc03lN86VFxldh4uv
zFPMfmBMu12FCHLQ7TkJs/fC8nw72UhBPtrHISKuH+5pFitMjYyg8mKedU05zBfrBvF4y660wBJu
6F+yVMRT8OgbZRU5vcV2pZ0thNuPQhul8Q+hLi/XQdkUBVKNyNvSYGciRwz7to//Tr9dL11BO77j
uhwhBvX9MjF7SzcP4whw35tm7D99qLqXPoxWzFUxv+outEzo+z0Gp6A50Dzs+A6KoH6Pd7JsfVMU
r/hMX7axDswTiKp+OjMcFZM/lnGCbbcch9zZoaFAXuxTISwQMAml9Tfa0e4X/U1Q76W67vBwwbQc
gUEpASFvkQsiO1noQPqQC0lEGRfqPeh53Dfw12VDL7irClKYg6gqi3Nle79C+Y7DsaxNraaoDO8k
kcrpAVhTLp4A3EXv39vnJYhMuy9k2ydedNkGnoDaqIYKBOE+z1ChXDIaer5os9Y/9vI1bzzIJT6v
KROAhkiSCsX0E45LnzzWWWdQZG6dVo32F4Lz4hByb/0Dp2gcVYtaWCK3e3ZP9BxypmyQS4UBkzqa
q8t0SlE8cw/t61Skb+AGSrjvVf7oJ/CM/6zVEBJSTEtqJyzNooWRTEX+6ovPjzr+jsHFM2TtdpUD
Rq5eIW2m7D7u0d8M5kMcyUI3rg5ZvIrd/gKC4wGXqUkelU+hWsFMtU4Wo8Elzv1qWLBv1cnJySA7
pwKoZWcyNuiAEqjrglvKAXc6gpqG55ElU/anOMRtkbjEoLWnh9laZQ22yWYfVttgHFbvJfgwyvWP
foXHs1ftjr6TdrSVaFfFGIIyNaUy5aXJNhD/OLuYSDpVy45wZRg4isrMbpxTTBuhiGG0H/pIEOqr
mToj6WfPs5xNsAUxZWbiq3Gcuov2utywaYkXRGrwkUBfjRe6VWK4/EsXlZeYnQ23W5FpKxOJjm7W
LzFue+BN0wOIUJb3Xjyj/BuBGuxg9cva9uCubKrWvcXS5okBuRYgxrKq/H0+QZcPkpXMUQ6xz+OU
uSuY5QGXkz/4lDFN1JsfJPx+/ACzPYTM4mSPcj0yqZkNJnJLFFvHyzosYzfmvRKH7hqoZLFmzVRL
HMHdfa30ocCTZin97c17QBhhPdni5XuYWYEPuy7M04x6tjj8EZRYA7UuZkbs6liE0BO2FMdgAkr+
sl4itKCRiWO4VfIqXnKNiFPTfNVBAfcKBnF2Bt0vKu3Jf5qQx41zxT4vbcFRs900RlLxtJ4X3gEz
DZP/PPzNvY1t7TSK5Nqx47XB0u42MynCCpx9cYoMjGa84MDmAAN8YQVFCMcLOo8zeSHK7n1co6uV
YoxhCvme6VV7jnCMfZc1z0kRl0XGAc//BlhHxzylwZoEjr49MU0bkx4Kue7Si/30JIb0b25OymZ7
enpfrC7mTew+wuFLduoGdjCHSHmViEGn2F6mZNokpTkbromUHemTYFIlH3Tb7NeaRSMJP5jux/Br
wTyrpslY+bajEzHy57xMugtDywBEbDdqF8vWu8KE44nqzCFmnzYpM1GEP+t3mwwO/tvMasEnsE2P
HABqeh75cfY+RCO/jEq7gBI+RGlcnaLcDQLm8B9aGOiFtSDCjL6UVFaLHDlI4hgEv8sMSaoB5sCa
4LqsqsWOSnOowH2OPWDjC418ofYrc7GE77Q8Xu8EW/jIlnfhUYiNOEAbc6bKPbhDAieu5RSyCjXh
Railv5ut092ojOgmYNYWzaMZrM1JPK17v/Op628aOYHlXcGX7iYUWuOGn1qYF6xSsxbvLCVITkMi
cPnJVieH6gf3soqk1dv5rjzId5TnGxkTLNevJKFYy9S1jhIQFDBOaV3L3d9efTgvqbloL2f4HB4I
pIfQ6dIM4v5mnCSDffrk075K4AYdO2Us9X7D56dsV6mSxIWbvkfwfdTKo+KJgXfagv/jK5Ror/zC
FGThWZ0ed7p4LEuBTtwlhZAbQdhSC9bi0ZXk9IR9pV+nkFBtOds6eL+bV2Zn5IhPkUhtDUGs18Fx
n3q5v7VHC2yM1iTW0LZWLL5/sU/WoJhvPLpo9W0wMvFRrw4DDxWGQiiSTXbCJzfBuA5aRBTVM00j
QwZorKuvHbxJ+UItrwWM16U5pkJE6d9olnlF7nHRDcq7RwkHiRtXozUgn1YQEZr+hLRZVcgqwghC
d8N4DjpiJDJpF4v8/N5+dI+qSHJXWKwq46fCzV4nN7Vl8nyHfChK6JzHIAoXbMopmjkRfFuttrfN
kRIFUPE3gwxLvO7uQmj5f1NtIObfetCw8PfUQvpy5Pvlv7pabe3V9aZzxA8WD02+msVEEegtBL1C
EwpgveToRetIjfHlTTn1Yt6YaHtBIm9v5FCyMIqvWZxkN2kayMHAiWn60iF745AAAR7C3ZwapZYA
rlfCi0JW3VHxHBRmj2hbdBAPtGBVuMaF6WVs6BS6yDxhb5D87sbJZg4hO0EhwFJV4pi7x2QIpSw5
TbrqeZUIQC6ktmTvpXU0K6Osf+nHAMQIiAhQCrWDlBt9r5RzwPqq2EhQiCbH1Y3Sm1LUZWo0wxml
K42HQPneEznd1fd51H8OnmZj2BlWAXov1vAAGn2uuX8POtk87tP02R9UICxA3qzjjavi5CAzCnt+
2Xguf5LxCfQoUJTn4aEGVt5lesq+Nb3QFlj51Nxtfa2qpiWisqWQsnwxmKBob4IA+4CnL221Tvmx
26OoyZvL4ZZX8tr2zhEWHfvV79hyULKnsDqfi+VOvstSZAqyqQvwh+WY6kKPTr87DNinRyrNWYXy
76UrvsmVsc2N6//2U2TrKEp5ADgOYbOWtFx5zFKKZPmNdIeJKQFGUl9vtpwg30N7RsiXoFa5x54p
qRNVsVJ0sBkcqhoQpulbIXUkFEgko4a+J/tiu4/N0nh//BLPGRPsGEPDQ0yInbN/3Qki2JAOHLmg
HJzyQU72ZEFdjUWsrNjEevsiFRmj7EHL/IuExLBScMWUA5skFvCCv5FBewHraFrseIIvvFA9mUOK
RkqdVOKzOw9xRgRWV/6gJ4R75XTb8cfIBU+3CvmY+l+sVf088xVBefUFdwi7ca063HQnd5zKFqSz
fWFR6ioDRCIt4t3Q2eULU3wQ6PaBhs6XS8pFbUefz/NgQUeOLqWDiW7SZpBH0IFfhUp+NypVafiS
Wf8zXAP6Tg2QyedRPR7xbwcjLUXAw09Z+8qtBGWHEzeUM7kmcFCD0iRJ4seP9VhuPWK+V6hAmPQX
GUvN7w9DsoK+efwaXoZJ2EFOc9FOSMIfQaV9qFffVPDJSTGmSkqKUVIfrd64vlAtsv4r+CruSnGd
CYxVm7t3eGv4vBB4K7z02I07nTFhs+vBIsNVYyfuaj5FlowTrGPLY+G1JqTS/v/QVi9aX7ceSKlw
jCcSP9sYxPYzEWdSAU4wPOsOcQpgoFYBAc9ijQAoCdOU9FcIQcf6ZH052ln8jxgKpAy542buahq4
FhX4CE7JWxxV5wjLbByYdv7ThROznrNVomIgfG7BJwiS25uEG5Nx31v2qwnffvVmzPA1GCmX4PJ4
MiQsVkvuZymZv3Jisbc8pHii3LgKEUMzN8xYPMMVvpl2nZ0vkAw3BRn1eTk/i4+yO2gv4V1EPX/8
bq24YqWEDxFFHZkBqMprpkYZOlmZPatRCZzxb8ffi80gk3yUjIIItN4T6lIeH0p4KXC8Ud3f1rZW
DPYl4FGjYcaJHiXBGlUrpeaFeddUoYPDYwdtxjtF5+dlCN0kLTtEFUsCQL3rw2/8f2pmvRpajspP
Up5x5mp2UbI2+GB5yzTIR8ohDuV18shLiNLNMIQjwBwQOhV1c+4M3HqLzxwCES8VqDV0AQoSzVo3
p0o4Z2SlbRRrRDqE8rlYCvxXwvak5btcMZtH/wfhTDZs8QtpC8KNC9m2ra877FYUC79dxthcpf1I
gt5O577FgKDljKR5u1kMmclfzTTOv5pq1EuAOByVIi0u9K3NraAN1ls3ssE3j1PiE/SHLFGTDeHI
51JzyxMArtcyoEJ7xwV5dX+S8shbQ+eDFBrqDXT38V6qtIkSQqkaQ4jfDP5KbE74GKg92EfcYNz7
bCi4cwOMX1Lf9B3vONN8W8CTK+Wv1rPQ0pPIm5yXanM14DDyOixAed7zIwdzGsvXVbr+hDlwtHH/
GzzEDWkfB/pLn1tIVBFW/pGWMPAMxh3eHfyO7imTSYtK+cVVci/zSzHZnahj5JvhsJ8V05DS9bTm
ddXSDWsStY61M/oCMPCUxoSMRbFAYpx+1ozI2UbY+Jfo4vneS3LErNJQ6phabbO60yM63Xj3F2tr
cRWK4MvqnO9UcjgHSVl1iNIUsp07+AXEKI3lAwimnqDauWuoPBUdqelxrmEKbB+g5taLSrd6A38P
TwLXQsYJc8ssGpnf1K9wgejFvm5CLvkceaGKgJIZVhoun2KOCoNJ2i7rnoLE4N6G7rAJqNLNsYON
Rvdiz3a4fqRX4654OJ6JoDyACXYIIiE+YiCa+MLYOagbtnIKwPUhlPP4I8z1g+WuFTUjHOikhVKS
izZpJAjeMuF9cj+ipxNJ3AumqReLxaMQGmmS5aisr2aR8I/FUNppRQ6SUHcps2QVBS7PqSuTINhx
1f4SPSq1AUfk5d2erjh4zPfG549MVp2vBjLm/ln3N7ObqAE7SQt6sWttlA72R+ICcgsEU0ufKOU3
sOFZm+tl/NvccXFpRVpqaZqy9mOs6eV442PUBT6YxQ7VUokT7scTsSSdhQYnJS6Mtezaq0ZrxjhG
TlHSomO+4+EyRexJmGeoaPGDUVKVoE+xcdBKDwWyx3wxaBDVtX5lKwR5Hv4kzpxAqPEJ0QCNOaaF
BztsEDGlSVlo9lGJ8gp1XkCjHDW2QKmfaCCQ5SFUz/Q/RZYySOIjQf0e13Ky437zG4Od0UY22d6U
gJHmW2WwVGBNYRiXJ0DvNjJdUxDaQiNYt6N7EAXoC85lSYPeT2eZKayG/BlsWHb02rj4BBRzBHOA
A5LcNvWzR1l5OmBhlH3NWobSHnxMEt6vNvZgV4OB8Rn/GZIEgkge1qCTcMitMcn2eRVCFRAW/PUk
x3W8JvGz60OxXLoogxnaRmsmoO72DaVoP3n74A7ZbdSi7M37VCoTS83gccYT6kw2tjNQuwtwPIQN
BRxi8DmnbVke69eHDG6QeruPrTvGYt84gQRVQNst6HxGmIMixx/abByI0u/I+XqsV3QBZsLWCyDt
ZNHkTyvaKkN3OoF14x/OGZ8PoOywXccSusq5Ve7artg0j4lfCGn587HChPB8zYFOE2hcE9lFwYR3
l0JzSZj4eiwke4UW2ktR9fKq7Q7TzxH/Mo4kUn8oTSN8q4kszhROZ4Vet3Kjvq6Khsl18uEr6bJ/
tFeYq6vkqwYhpFiDM16Xs5tv3FG5FB3ZuUfPCRsQZMc5m151xw5CFMwtEjQ/ykC+5390G9IQdcp6
X5M9fDguufjB1NVPkrjzPV5JbVmH3wIBLTfUfzxI6BJlRHPi0VvvWOxVF0KfDoh6vO7fuSVl9/lk
MHSGY/HLSpxh28x26wcNNrvDKZBzo4wsM7rOCSq6f38miWPDEPKqLCA+k7Vs1QcSi5SUhTJUnC/7
pS/YSY9joluyOQBxWcK7AkXw0WtVsnh39g+FV0VzcaoWaXYX4TVArYRBEbYv5Ztw99JJz2ThlDZB
wbFemdSiJq1pUdBxNCIisNNnegKs9gTz0gR8GTunFcAKCn8/vuzvEhW2NnYhC4ln5nzAZLZGQTCF
mDYFC17t7UN8GbnO4PLP0xzlc1tGsNQL/ySy1eFpmzn5+6+opzX7NLJ3OiDs8UL5ELFkAN0EKZVa
34WHZRkEv20QyiutoiPMDJFgmkJTD40EiARRYLCmU4JngcOr5wf7ayH+Umgq7q7CAWixjAENbQWi
qDEeHM+CPTpc2U+KrggNccHSg6BvpKYQf/XA7dQZ0iuYAelzGib1ua7XhG93duGjx27cRHh+kef7
rJYRhqUHgeUhq/E5iJcZu0L8RHwWQ68UywEacCOT4I2KYwbinJQMMssgB8+GxAGcNYRqtQGzo81/
UcB8Ybggf6iuBVm0dEzBcN9raHt5rkJ5b4uUBEn37U0j4r7+mJqP2xKaCk+8/yHBnYlXKQmNYNQB
scogYESTLNsXCJ8ALuJadUOhIXJb/8qVZbbyeXSR44sfZPE5mlmIjySlIhKPs+tkizPrydeF0MMV
IPtNuMvDx+8ZIWchzFYgRE/o2CzqnnApgTJBQbApLLkaCDwVLEfPH6QxZ0YeP5iXSgpZUtSzWmBx
64JzpcW1+QAZ54n/2kfRNEiIwzw9vJQiWlJyJN1jaL5tKSYAf2z3ZyJ4mSX082Sx4p+6mxyvSrDC
Qe7jBOKC+08uS3VtTsZ6hfzI3SdrXrTGd0VtraxgCFyqPdwiRPeUbsVkuk+XU6lC7rlRYh4Tr7Bz
EUoVGuZgQz89RV9YIZkj+vQ0g3vTNnqnFUxvb3rss4RLevRgH3P/c336Jdq5sIt+5CSWN7Gsg4Qc
AmkjSNd7Kp/kGhWyFBK5PRGu6/b8xKovQ77EX307+e29Le4lxlg+ocJIlXMm59A5CgumGEfz6oOW
b/jIclzZzQobN7nIiL4e8W9g15JMqI8dYGaJZ1fUnfHgpnJEDnX9lc7QtjFCelr41iMOvKSdeQ9+
SZhqzYXygXHvWAhcKaYYyQjapQ52K+w4VtLBs+ezSfSYC2OINuNSjETGNejPNZ+IEUwVrhgfMOJ4
+tfPlIsxjjVndx063OzSltu5+BWo+oTaGMuPCJCx0CZg20nFsRZ/zmGhrVj8iskmvM8APKN8eNbE
z1BzTeiAhFATd1pUNEZkG26X7WBsX8UupLh/O10yHRBS5UWXBJtVCQDZjQzq/wy5MozlFi5NgQGi
9xqT+Fko5p/LyhbsKC0MrCJ8aky+JU9eym3JJaGt1kGMPdsLAtKzKn5KSjESphDOSr8OgX5By1cG
UusFhuKoTfZ/xzXsbuVooqSVmbWHaKOSVxvrQopiM1Y4FapuabWQJKm0urcRD96yosfOrkiEkGGC
hSnXU0NKTM+dMPajChPegFkUpFh3mTiFNLamGWhAHGpdP3o75bcdtM16atDFJhXOtQ41i5hVJXgu
pP/lvMCGnV/ARq4AFatlZzL3kw5EHQBBKrgdHC2pB/imuoRUdtXNqTVW2drabZY6iZysfnIh02RO
nN+O5KdbXFkJA8G40mahqZQUqSPoZ+LxR019FUw3tzB0zdYoYPettwB31ya4OE46gcomb8A5Zm2k
MxLKyW6DsmSOYcpau88K40Ct/GWHdlIpXWAz8LEfC85hvBbR9YjancIrGzwQ+aTu3b1ZimWtAQZQ
9kXrAkeBnPZ+C9uovesffnFNhddJQT0vLn/d7mDdjHtbTzf6A9P2TkOxOnHTugHk970hMGGnc/xX
22xom2gAAI5dB14k1ALWuEWYQqk07R8KdffLHQZfldATGpW42rWQ9Y6xlZJ+g0X6DvCKSrAfgCJZ
DyeXlIMz9fQ5E8zKrZMTOZydU4PsEmVD+Y4vyIddGJXhMhzmc6V2a4sLG1+MmLNwpQJJHZFVL9Gm
tVMGMYYP7PeXXIMPVEIOGWVdYfrJ5dul57VnK06d/sFHBqNsbmR8tWz9ZBv0Mrg9Ag8zV8gVfYsc
W60ZO5WXss31HaZeSR7GyT7ZGsZnvnfcRQ34t8Xdq24PB5VcphnrXN6iRgsLbSR+sTQuHz9nTvjL
lvprmv2dkZ0x/So4nFXrFMopnE3sEyAe4TAg3voGrgx3z5Egijl6YGy9plPzHccsktbfVPpLRWkS
0z4SMMVjRc7ZJGzflgCdG8FjX/Uz3c3Vft0JZvUfRkapX/5Z+M8iJmmY1HfcSzAuFC5IhqQIu7TJ
IdWOWDlQc+Je41k/qMAXmLDtnUcou32W5UvyjOfYr+qtCj/6QtpLFgLex54op+U2SbsJM0rtaCSx
LIdwjacvhvgJJtwijACUcyb3sBaJCpzzjiDV0ttuIIS5fAj/1lum3cFJbofqRcq7lK1Up9vhstkz
ryFtjjPZw4OKle1zAtW9g4guv/wWecOcqslMkfWBJDkxUh6PJXIF4YjUEVZBqxNmmPxjjvIPwcuJ
kODM4X+FYZLeV6Kgv6W0CgLe1cVNhOQ/KJFxtRtyyHgQx1m4ugb4NrDWZeu7yEPwf3IoTtwdpJ7M
pnnezvGND4yPAUQ+8KcSQzU9xn9zadb9B8PXm9PtbTOAqwFTSY7d3yoemAMAeWo44V3RFju+uvu2
P5HgBksxhkqW4d8Pa2W/vvtb//K9Zn4ltJLDbiJP2SgGthhZk+1xwLk7Mw0oOvn0rL2Ykr+0577r
arT7Ui7cmOFAbGN6hq8Noku5y1GA/zZwBm0GX9xYacOxxfna3vbhSCO0p9qyuq1mwow+kt4k5HJ4
unWDiuaeQ4awKxfYlcOe33z4zufTz1d4yzDwT1hZrYQIEDs7Y3SQppt0z+qQ+EWQvpmTpOtWgFc5
7+Z97RRJNkiVGWcLhpuDTSeqgV8OV5p9IEuv5/nwTcrdR/LExvKI+43swegpIkpHpU8ZJywHqGEH
NgaksTPMzeCCxo/qYe5kCo5QJUtBCV4+iY9pK/JfjvzzHMAJNUSCw8q8f5D5CSX8wbuRLQnLWsij
OjiblwdzVehiu5+xRQox5C5/HhZb6BKq2Sob1vaqLFLy0hge0f+jDNWuDZ4HoXURh68/CMInWjAp
f5A/+qvaID53vBSJOeT7P54X/Hrnvflc/tnQzIqU9vxi1Akozz78WFPV7B3BpyQMThnM5B7SbK4D
KZbw1DviDHhG0h/acHwNdne3i6pYrPypcSg+KlimgpPieXp3DjtADdzM45MVBXRLCsMpT5XCczox
eJDPFd3UV64tIxsCa0pcPaqCLpY1HoTncNF2U4UDPej3bppV4QawUkS/VBKvtmLoTCPDCWDUpCn3
VPlclan/e28kfNI3Ny59HPWdCTcUkQj0NC5K9oVRjkBPppGqen0nHzeg48tNG1F88A+pSvqzPmn/
Ycg8IqSqLQZFYaT1MVeZb9THfqQ56ie5dXNZlJdAYDDGMj/0nw0u6Ijk/Y9oLUUMDVZobEXVG1RF
Dazf/096M5Yh6COHiRzsddxvyoby/Kj1PjfacUbDy89hzN5Kyf1q0Q5ATEkxSbBF8FIsatWuOvJ2
GBxjEpTjpTXMtqGg8Y7Sg7nvhqxQbxZSDj3ZiAp8p99ywH2MbV2Zz4/HEPr1fDlsfxRk1z9WlNIb
PpXuMUQXuln+/KEPgwXJG96KDXrkP0bpvgBZPV931VUmV9EQWxFpRIQIy1JI8KRpI/xR3n62uTCp
UhKo6XZYHQlN/NhBlXKhvbMztHi8oNaaYoWW5m9XN1noC1nOaN6AwCjc3/e4XVP7QtojbF0ZUWvQ
ysm1CKZlFQtoi/9WyKvi8JsOD61VGRwccunp/NNLSmaeXXdDO68axGjanPeA1kDK6ggE6VzUiytG
Xl6sifqEnCEslZOq5JVsrjNZhXOTgD/vxjJ/FbLjotL2c571tk/jkoRSi/Rhtib+VV/Uo2diBdnT
oYGkvY4Kpxo/gOxSHjKpHtEYL7GHJbyfXQ6Og1gxDNdLUWw1c2beWJ0uZqH2q6VBkDjr9Pkv/a83
+MtTGTGPPRsvNx3cmvMECPv1VJO2MmR4YMCLEFdOTr0+1vVgu4BeIdJDDMhzcwKCqQfS4UA5Y/cx
ObelRpjKdCkRrhecK5jlgh7tiEAMaBwwfPj0pFauLQxkCXtsb2Rhb7t70SyCIDW3Cpqxk3W34Iw9
ezOubEdu2zZzPkWj0uT5WhiMuVshgkdHEf+R2eViJWgYEp+8YUn1VB4ZPShqArR2gt41azopyu74
HFS/IWpevJXoyLeAw7NzSOSbNvP7UCd75/mJTDqt959qk/FYhv7NKc5FYmXvGHCaS7QuU649GB6A
ko5oh3ln5aeRIuz3+2TGjOtACTC1ZlMkAWHHHzcUz+e8IY/2/OJ6uH5BZKzlGT79/t1lNAsYPTku
5gWbEkPFLJzkUX/2qmdKyhbUK3h+WiV/GCHnphxR0EVbnbLS81ku0FjMPwUOqWpFEnHLnD2aL5WW
M56gvrchaFie7QWEKXzy+LmjasinGQHFs4fcNG6QFeRPsyeiujUPc2ayzvsaWB0zpUfkjnoVpnjg
0qfpSBfoCZe1ogpDUEpAk/5PF2SguBvLTvQIqA/RoKeOJAMSZcyo3wOL7o6JUSJAZsCfzfOqVzDK
5p/ShOzQgHpiTESvSoLjNl2pXWe3gdKld2BkiK4s5BUxr6D2yYjX4XKvK6aMQFYWkqmhraj8momw
fVcfaTh2g1HPJIutCDYRONX2/4RtmAaw+KOIvtg1JaLfuL9SDiyc8vdVSG3k0TX4uVSYZkLlNJzR
xv5CJjzK3s+1BnQQPMBxI4cWfx1Isv9ftIRMOV6EU6uCKeFeF93X5sWofavWni3SRbgdzVK0Fmvu
X02zP4ofJx7ZgXEBN8Ej/pwitMagLjBv8vO7DhsHGBECb+kFRtP5dl9gaQFKNCBULQPU7dKtEFbP
NsyRpXN3rmRdBrQIlXVWHs/PxG8uXfltht2me6BlTgY6XTUWEBMjablUbdgdiTj1B37lNITIOGTx
cNNafJ7RmV8r+Dl7eH3GF1qrrl+Fn1mc42S5ub1rQEpEKySMs/I27GJWchHgns3rloiSsnqQ5fAk
3rKEcGHzdAJei4De2lfif8jAxt02w8tKwD25JKV9j4gysCyODnSvgZkbV7XKazSTfBXSgybFR2+C
Ji0mbfD61sWnvVnLslB6I4dRgYfX+T2xpAhXA6tJzyJfYM5bHv1Pdc0F7LL7kcqdGJ0t/nyopYzs
szTUAVJzsN1qsixWogPvzsiNsSf/DdZC9QgRE/nqjv7gmV5Vrb4/oFIs5qdArHV8cEJiuhoJFQpg
+pR4BJMA7Lpfce+SwRN1DlhOrRuO+muRLT5DBD3wcahxsWwAiJZer7doULtsDQxjYSSTU2utPnK4
XDiiq8seeQt44/hoXxQ4ZSM51oo1DljOZj0k6KqWA8ZdyzENTyXYKL+BUzhg1NRvT1lr9ZrEm8lW
UMZL85OX2YjXk0+NeWHhpdmj2oywZX3JsJOWxLgADonBeqfdpin4ESfI4CBvzu1odSdC7jKmDtF+
Ug3zVowaCng7SPf2BPHYY8WmVjOCPKAd0D5h9F46bXL916Gfb4PKloQZhDkrTD7raXkczYLm/xPn
HyrdsyuDGdKTOWPBSxmVTuat324mpvHWspPtvAWVSR3NOl3rzRgYZywYD2KljkWX1BbjXCrQVcTh
upKMT0W5QkwNZnAQOswGKJeEGgSx9YbjOHzhKYjbOjGq2/wS66BaCugcrx+UuuDI218Pr63V7bD4
P1M3R7SaAFsBhECw1b/UjCNcM0ZNmF7L9eUjN5JgrtdNymzQCXwVuc3FxVqR29ronOAkoq/VivPy
KAz1VABYyh9EMDpEv5g+duDgpwryWmsU41dzcBdBNJENqfnLOM8IN49NqSnAyRNOKXhONx/WmXxr
gXX5aKK3vIYLuGv11eKNnypIE13e+X/IaiNR7rks3vlMYUCI/ls263l1JlpUZZLhprlT2mG0PZts
/MKk/kv6SVNgFyQ/Y2npjKNFtV7WlnDiIHuGf6j1N0b5EHEmxBporJCgHJ+0W6ViC/oumeFz/1Xw
BBd4EqWP8c/PQ21Bw+BYQe0Ws39srbTkubUuBT3NckM0lcISVd/9SQr6wb1k/NPk0gy8sy+yS53n
d3mi/mCy4lIDQVFoGRkOT6THQ5U0Da5kMULhMAI2HxoShkttPGL6rZGCtGGsGDC3tFhiuJRa0nOy
uHihC3SllpQaZ8dLKmzjxXWFLcIFO6Q+KS/3sVh8Vtks+NSJTrkRw6AezvE4RSifz5x0HO8vjqsa
KTLWvhp1VuDor+8LlcXOUB+3y9DTbcbnPSM5FdM8WfHTt7gwqURheMgRXjm15IckLhDt90zIEjSp
aCiIL0sy11t/LOsW8kEjOMTirU7mwX7UlzJ17vkx8Ss7D2cbyQn8GKH1T/Gtyn0Dz3l97DaAIkq2
heeJMfNr0TcLa+/xzN3E9JnUPtzwNhFfkTvB8DYxU1ogpyXfJsgwVxAB2W9E8xAdg+ByIUp2uwTu
rz+1io/tYrHzoktpy20kTcZ2OLtBlVhNmi8cdpHUJLe3z87R0zdQxToGgAOhC4jhDt6aUlbYTViC
hpsFYGuFR5wwoRZCp3H32eS6fIWsJeHn1ka4fm9NcIEb3HTFaTXCCNM10yB/TooF2ixMp1TIk+c6
BVCjbFrUNEj/65TnIUGNwTJMht4qfR9ybGLnrQg8Eo2AP47uWV73bV/jChVJ6JsW/KJ8QyAXK762
lFNN2OiPZeiOaB/Yf7ITnzinCmbZCvCFHV4ow5G9QK+kFO9Gg6k0auKCbh4kqFaAs1QcMcs/m2f9
zEMzQo//EhtmfKJpFjKYpbumPzqaCJ5e5GtmbTEtljXPuZeef5knzkpDucFJ2UVMN9RNaIvLBz3o
BlUqKo92pPsRHV7p6CuPVMAfVU5OyVEFoqrYm249+580RIz5bPYTUieCbNtrO3n64ulRZOFGtXgF
abK9LwK9CGVc13wJ0klJaSlIDapTBCsFf8Euyhj7RoIVKyzgZtoZP2nvMHmCXQx+e3O9WdV6g1nF
4hZy+fYlxPclDtLnpxlh8NHaeirURwTjDE+4/tCDknUfPSrXBaI7p6YCSafRHG5+Nua3ZwVd/vxv
QCouELuZShPmeFjRFD48LP3+A4Qdw050975cu3q+o1vOY0oAY8ccMEcHBg/N+Q/kjOQEwOVHL8kk
begE82rDafygL69R4y2jnmXylvSeT1qlTUgVuKGc5w6UZunLvgmaKDO+yWNGd57y6Q3M76aaLQKc
c7wNxux8vxmOwX9qeSVhfoVoWQVFNHnNHqiqUdN45NgaxI6pbrUn3vXDf6cl4nnmHhHKUZZiw/NF
uZO0QI/x3+N3rT5L2Y9xEM6SUb40u4vmFXoBK0ja8Aj1dZhv+IkoTxksv7OpIXjfVXOmXmOVRgl3
Ff1xTU6PCwmX7De1h1sWI61x735SMM0G2lXhPsdgxlsBnbXnbLbl0jUGZ/CYhWWGKnvo5+C7ZQuZ
JzD8BfyIga2DmRVBhQ1Li6FUkyxy85vpF4Mct1BEPE9UqlfHj5zrTVC7VkTM5pl5/DpFLSLXg26y
Tor/KdumLP89IB3ubaX2fAOnI/6ceqFhjVB+L8QIdcUiHbpHlmXqJSDV5lFq5zpf2LHGO90Tcvpz
sXiYSoesTDk5S5xwZXgQ5Jm0xZErpeJtCQmaE/cxR8Jqj+nZzV0Q9ojmRlVAyRAvFGKMw2lR2PxO
zvcHR1jnj1DnWynzu284tk5H3uuBU7cR7whj/Am42pM7QYhmA1Pak+n8SMDvwjL532pweehQx01x
775rPhbpHvTLs+3HwZTXAXBfREACz5GcWRxJV8sFdN5lriUFNwZRC5/aUqebO/ThZIv5bf3SOTuz
tfAlA/Zm6p6CMQ89dPNx1UL2wfOJqCH3bba8VMuipiEoTHK6i1sqxHvMt3JV08+KqTD/rP7XoVhy
pGSavFafu7h7bXo6e29XxWBFDAzWHkc1ZOaOiv/VvVSbMK/ogiOUB8NbPNOH/EeeYGECEL/jZhr9
H16Hk/q/6JR5njKFGnzfGdaNAqhcJ+JzzAn7tN9tLuaOdecucGbaGC6/O4Wcgl4JQXB7hWIPBxsp
MAu2cmD92z0+0e2PnRenRNRGw30aNebyy0HqhyGuxJGZ9dES8pidzzkHU3D6zo5NPikichVfM8JO
d+rxjoXIYWWGw0CpMVFRf1Y2zviDu6JKOks1Ne7UUTAjnwOTJTI3TNNqdDKh5M/NRH5EaiXmCGGP
BWRgaERdvbPW8J3xGsDJ1VXKk1csSQci0eR/+vsSt43Pf3hPkN7WjEVvIuSYDwOCE+bPANysoXOB
qd/aAwfyOLtMb9qdVE2nrKAw5Vgyu+m93OiG9yvlW9TD7me5RePOt0/XRH37kNKN6n0fD7P0GaaF
Q/YCF1iqTOuoHDOUCbhiu9P0+8f4spyZkzKISO1/OFIWEEScM677rlvhkeG2eRxyjBVn8MalI1lZ
jAKd7wtMQHQlVofaGUPh2nNO1LmuOrkrQoBcnPC/rtm2SgTMrQovGLSdITuU2+v/lHAxx8XJZfG1
E9rjVS/jYmIDSu7Xl5Q56eFASihoB+NYZrXlIWx1z5Ru19tJ8CltR+tH92ml7S46S9jx0NdkUq18
Hr6O8j2gqYE53YUUotDkDyi4noDpmnzz+YsiIbhtQwk800FUZKMn9oKychiYP7xX72Qx5p4k+70X
SYLdI9A+LcD0CLu6OiuN82jHbwe0cMQgaWCMD8mzYP63p2zBRVtCnnDLbO9Xeb2bWvCn7k5H5lWf
JDRL6TMlHRDxz9xzpxktfuxtDcDQbuXfGI+C2OmrFdGNQOqiQ56IFwDMBr3qT6UmE+axEJBBXovL
IXkCePdUdRM245kR1ADSbfR4gVUABQ5R4hgHk/eXppZYQrwf+NpZLwTvWJ8QK0hTIqgPTR0y5/yD
jWrW8pTAioSY1S8KNckx14XxvB0Wi5b9JBb+FejHvlZvHUkQXwttMe2uayZhn1hcNUgO4o8a2vTZ
XhpW1VPCFEmmaB6/XuYczTTOHx6e1FmjIgZ+KX5MSKXqSEUn3BGRjfRrjaandsBRBD/QYycdvXLs
ILhBrKaGi400Zfp9BTFM+PpbySIYjRJ7FmSSXGNLtusVvtDH8lN69apGaLI3C7T4ZS7CSRGhK1we
zEEhEWE7XJ5oUdbKtkqg41WDqG8JDLAE97Lg3GUBXIq0bTzzsiGt7S1dMS3EvqCsd2LTPadxMS5C
2TjFV8IL28PuREjoaj8j9VyZJXwMMx1lkYs0j/xv9EjJosrE9A4jENSor/CDH7+CYt4idwYgGZ9A
AF7ghtKI7lNxJjFpoDDK/rRiXkipD6JEervzTg3H2G02W9eNHPFj8pamu0g+cPlVUUETKsUd2c6N
jji0Z3j5pMNbQVW8qcQy40g6bNwQGPLqL8c77fVqiYJBXfAge96Q981cnhwAxuFT/oIfVQ8QO9UK
vVZt7qjcOL2OM9abCjzEpFvgQo7w5keOYrOKn9EelYUtO/OrTzjFgK+Wp3asx2KWKrvUHlsatTvk
mL/ECns3Y1SZGhkDJLKoWAecpBxinzA0l0/7Ui7GNtPrhKQVF6HV+PyL8X/qa0YKEHshXW66omaT
tRddSGFfn7VKI825Mimf44slwVoHINwFCha+zUN9t5qz5xG7EgSe80+tW9ZiTkixAtjSToCKafWm
1lRv62jYj3yYBNDtboUdq7IAz0ZZRMzX2/5PGF2peaWNWVP0XQfxXTCDItaSDetOi4tIGHuLxwVh
EGzKyjSUB2JSMV2V98R41RWjpmYFCfMcKUSs7Atew0cr3UAQcdXKf33SOmsD5VnZg8SvEE70JuuG
0AKp+TqGLV8vUXKvtF0hVQE8Ghm1b0gsmM77Tc/m0y5od228eFMYh20tuH8iGA5BoWzSPmzs95jF
StixUohY5m+APz/drHqteSUJ4/QC0XVXeW4jGPutty0TnXELBwTRMk1spZPndoippmNcmUYKiTiq
nSeF56pb1D0yT36qSxv57TzjEoMvDirqKDjtJdAEovrAMmO/+CIjV/fG8tVaCst/ceWYynbfTVJa
BIMtjZcHmb4GuVUYi6E4w9/Rrxt5JmIwge/1+/KVEoM0p8E1cR7SwsDN8iz20Zuw46ZLkPRE19/c
jtDY62PXJUu9ONyOOdgtzjBWasXg3ORcQSNTTa8cf8X0mrSw6z+BkX2/cSPb66gzeqVtbLS+yM51
AAA/73t7VXkG78ieMhyRFdKMcZe6n/D5Jk4Z7Rlb/xULt/0O8tfaKOyNqEMcQrTm5gYATlw0EMd3
CCsvx+/E9sypDQjrb+L2+rmYQnH3wnGq6lrKpO7kTPebpQA6nev7vfZ7Y/TUS+iI1JDdrgSeHRJC
k/rY7AzuRW1y6Tetv4ubLhzKbZ0AAqRWLZNZTWBmHZ1uGi0AhePjo3Ul/M8GFAFPsPQiU+jssHaU
ON4KvQ1dsbiLwbn/+YQHjNMS4FYZGPqp9cllwK2vmIjBIfTBa4nwc6ffEAYaAQkoOtP2Ed9e+dVM
T7LokwNYRVvY1l2NVCqoEfH8EXOEf9pEoOpy1ye4WM6/RBcJLVXecFdcQmiKNzRuHUF3BnnhG85c
4+43Rw8+tmTVF4T2e/2udFg5rMZqA2TSfbrkjp0CpKYXGXzd57siNcw6ZBw3RkiW27UAR+GYxe4m
QtYVdoDabHVmM5YiA9ImfvFb/P24YVG2666U55WlFOlmgEZsIrXwrYQvE3iXz731l9khTxVDsXuW
FOZLXPFmP42k09zAe8V2NGN5tKJX03t9EUQuLZmX2AFLqurSgAbhGD+iRxsCM6QvA3hVqKVH+Od+
nJamBURyexdvHnncHtOfqxE5kuUxxHNNeQNrHdBAOev/1Zo7I4ocViaYNVKgpcuo7oQWrg3i4g3m
m70TnnJFzJlUNUIu3c9fTp3p3fDtJNrK7E044at3ah1SGlHsD2MoRXdOxdAQ/PzZFj+fdbqQk6id
W4Aisj/AdUQlID+TnMNzPeDHCmQwl+0SMhr1NhQ918gdcrB77L+CEq6reCTWV/SidKjTon8bc9is
L4q9y5C23YPo92TFbb5ZDsaD3cUbRvn+XbdgjNaMOmzVAymAWky2A/hYJ+JqdG2xDiROEsAe4/M/
aw/+Antx/Nw771/vYHfFpVAVCzQRZF4owXiV2vWzZOvnjRw7ku4Kv2nYpy+YW8GQV6nClfObvFl+
KMgKoUPzkmY2/s/Z60v3dFEIO+ZQ5jFIGyxTSjd35O3l+ZG/TP2RbfHFEZ8oBHTZtSkq17AdKBQj
TVzEPVabSzUxSxUjczy6KKo3yaud0UL5ESkCFv8QwZ9YB1UfV2jKEg3owC4cQfdqIcOn+0V3P43T
v7kNUXAz5NX/T99Zm0jTOeurIvMdPognVS5hlNTmQAtWcVbuYY5+YLPwDcMSPlFK6sXEZcXod91w
bHttJUhU1qlf3qZop9sisUn8Jl7xZdZNqBMbrTWMx4PCr63TOE//LYYmFfI680Z4NeSBXDhs1EN0
7HcDLPlY/n4uLjMPF97zWafy6RZ3xmTT1+/ddkT06+Y5m5Za9aXRvJcLn0k0C8kPyI2xVovbib/D
6kDI64FLPNUk4DYcnFrgpth7Ntwcn/hnkrqm/HCqfvP8kzmg2EvsF3/HedfLSkWnTWgvn55X9dSE
rE9O9o2dkLVQZkW3Rw0N+GsVwD/d1EoKfZ+j6ztAMCPjnygi3HE8SJpnIolbhDsMiPRe/1NZmED1
4e4KuOa+/MenNqCxJ9VZzt5Z9Ve9jlZnPxAWizimvoGQ7gUHSGd0BVyKZNBYsEAaQEpu5fwhvNmq
D8XhX6+MU++Vmug8ZL/trAvuY+9bYTF1TrovGnsJ4WQiIo3vi8noil36AtRMlNrDxe4G5oBuT1D0
rJWdpFGpXdXYJ3Ty09fINtvuZjeV96d7SfmnfKK27ZyLMii5qVzUZAqObNrIXCQo4xVbkP52ObEU
1XifDXLuCpNvUJ1UWWn+B6kuKuVrvSpnCk4al+fkbfm7o8WRaMiyCoao4L7PuodapwgcsR2/34rj
HNhssJviMOCy6yRnr21x3WB5xbvHrTocqWXxbuDth7L5olMcO7z7hP8S+0XHr+g0Ts1X7MLiL2rz
IWxnD7pQ8jln8epDLLYY+XDbtq5SNuQaRjvvyEffF7YiRGw0Ll/avdcDR/dzN9Y8u+w7zuV2a3rh
HwUPYlT7m/XoR/EeqWi7vB9oc/OLLJjHqnlwsqVt1KudcIeGSgL+OSkT9wcfZWxHj73PWaXhifO/
+Tg7IEoGBwRuBqQMlfBUEYloOVrSu8udcw3ouipfWa2PNfKQs43XC5hd/y4I/FnQomRI1cOWdWGz
5kU0pDU8BDbU3vo9CjDERCVOrhuZwoR2M73DszwL0ChLnGQoNU2H+0ma6c8zU6cprBRaAajVdT3M
1mSV804JtWwY0naRPigsXmmk3thttu9vkDBS8+fTHZkc3a0WrHGbxL/FSG4hNDACA0ORe55gci/c
qs1woCrI//L7wYW4cK/7XwgsI9Y2B2Tq0drp6+/4WWJFET7RKJALHwmD61D8dNf+PhXn3rHiLDZX
d6hkXo3IvPCGSI51rW41HiwmBdOseaqaP2vbhM2yZGcphe/ZrRxT8WTXVovIkNi2bhwXW+/78P9w
V6swAupK4w6ABuZF7o1BOLnP9IYoShROyYa5/33B4jxj3e5ihh5hiZoy2qlB0mZciKEdYJJqnOBk
xrkK4scwo9rin8v3T8Mbs/XQXOs2loynDWiyOyPNQ/OKRz9BBw/isQSQCujeMTmqUVwC+11bfciD
eyuVJ26C2mS7G40hoEmj5thDV8ycnqFOL9B3LkTXqcpUtO3/e2d7xGAvNcQ+RbaZBas15JsrlJVn
fFZdDIUAdKyCRFJ6CPBg1ORXLLW1Ree7hEYZNlqtHuBm+ydf2UC8F4doUfl3byAoXDRx+rC+udNA
tW+GOtcQ9gk/zlQ316k6xIRfNhVXjvDFN12vxoYcDGw9Xd4bqYLzOP7e7tAiAvQ2yM+rE5DFPU9I
J/a4j2SLUUwGSyI6pZvqRFflIIuEC2sjfIM3g7RGEMuapftY7SVuhC263WY1FZxtBGvAItjlqKMO
uzvBOoi5twB4g/qUN75udWSY18CJ1ON48pRbBe+mguHwBBb9S0r0o0VDwxbrdoy12CeZRGffP4Z1
IO/XmiJ+WuLGyCRCK6MchLKAsJ2ptkFxJKPyx2ZK/8KKi4HyXOYQFqYG5j0hgamszlErZwKfoa0e
KQyNjjje15oXhW5px1QE1cjzNOo7dR8ltPmmFrWZiMDpIhKdf8WA/DZryAhTTsOUEAdhOx2Il3yy
5bIgljlTnhkhilzImeztMM+C/86PmEe32ZwgVduc1Jv9gyT1z8zRYyM7W9G77Sk3/Y1dVgKI0djX
0Sb4Os4k+VFtXeDRrxpHJHphveFVIY4LNxVRXAf6aK9HmtP8j1N7PYWzvvyMpNVaPBnNnorddTAm
EQh7AIvuSJdg5D8evIAwWSKEMpLRVLIiHGklZbOWA8i0T7OxXaOUi4IymEdORHJEERLBdaXVtaEb
1PPJirAI6X1wcQS94EdQEv/MO533bdWfFfOxsqnLEx6WmjocKlWACHUSkcdFCynETISGX7RyGzpv
n29nHcNXTrvTBy0+7z2+XwVsagXjLDYopO26Lcgb2V/AFOVWvwleb8Z21JgWUm/BXvm5586hZVvO
JeiIiQ+GdjvdDtfkZGBjsaI2ylzNdgD8V11SEx5E4cZYZbVJAW4TW0dal9fPgoJ3Xsm1Ta2D6KKL
iunrDCh0tZgnrxnPHEAb3/HEh8hIGVekEmvodesvWcg20+vENqxzfsQSl2OcqK9klr/aeGKO8DyV
PQkCRbc6+wUuu0cK72ESWdnvNUpJIMEHzldT1B7ie4Nv1CriRQyuFy1M8Qmgz1osjMahL2cfTfGl
smEN29dJqj078bg0Vvw0I5m7+qudMBW1iOkqhE6v++aWlFlKFhf5X3L1th/ma+m1O+NNzpauT7GH
+YsDGA55gYDkw9yLzh7iC7Zk8Ff2PMT0taI+tuuKh5S4uYZH3Z+Jl2Z7ycB5sxUgk9QDpwLUDUV0
ARPVH6wEY2IIJuO2aI0eOfrtHx+SyQDZ6+BQZ63WpIF/4Hai2FTm1AEtPX6AkBF/EANcYxqUZmSx
CnEgKvQDmW4EZm6zodDRFKY4Z+zB5OdejF8XTjcx3KmUXT1Mxt8+oOYXpFwDCTV/BkQJKjcxV6GZ
ezHnY9KpbcqrmLChiLQJgRiHPrlnGbQWaD1jhWMzXYnM6A3iRWbs1JEGzeaNMbJljz0DB3H65L4o
tdYBI00WL+ow5rEsZj2PvnPgEtGThkPplJX3rAklR4yQCgozTBEUcOa/nqqSLsKYdeD0Z+j7BDAb
Nflg19x2OhEgpdkPSHfkerOpLU6tWtxMwIfhy0mtefU6hevcYm1GT9EuRYzG0fG9jtXdWrkyBPhk
hTqz50WUPFipc9A/pwbaggK88qB+6n19UuAbt3JKatJxy/CC3NbisS1Ml/9yL/6oE4ugnEqnhGjS
xgn2HP70N7LVsglJfEav5dRDt7caIunj7oRb2R2sHyehCkmCiAG2VmvIdszJNdCQb2Cu9B5dLChz
DOIxTNKNcNQeXethcyKV6EtBQnzwzcN7t8cmvQpYuK79z3uQcrnYsCjy0oYpirAT0/4xNGyphIFy
qyOiLxLff4Bpi5bLUlbJtIw5v0zrXLjVvLPSiTM1BHvJ9jJWHGTiGtdZ7MvhptRipwQ95Oc7dgSX
Uw4iZ9m/tr0tYq9+3uXQwg0dtyF451zb2bz/iuEcVFv5eWmO9ANGD2tLbdI14GXwBSOrdh2moz+F
HGX7e7BsRvY4Hcq9mEAxv50zOnI+w2QnyoN5m3l3tE/Pfh7Z3C9T3UN1tEvbxeK21N1kIIX1QvtB
qTIq9vDTUg3IxNkD4rZWJx9J5y9/Q910FsxIVHniAlNMLWGxHOQZemOllKPfZly1E1+ycC1spZeE
tAHFy0z3LYw5R9foLdp88vbCPLhEaktjDzppeKcynhf1gQhQ4DOY416u0TX3KXipo6EmBiGBfcUL
diZiPVyMOuAZJAe+uOf7e5m5fV19dd5lbPC0z7IybqAAzH1pFRzigOX9spuMm9a0ARsIp+6bdmP1
s3RqOMXxJuTURod4rSGSpIH+E9ysOJp9/NZOU1T6X5UpGlE5eQWDHGDgPafIvpyiYIe8k+yLWYBi
3EFdxPASkpeynk4FQUXKUYuUlVFMC3oUkPPxJzRWEEDf+K1lFI8ehFSgHyzipad3pRCBmEgu2xT6
3uwt5F2NE2++9KY5uk3HN6+F+5E+rhUbNI8WoDn3bgV0goxPCsXxaominslCH6A72vAltFAWzjip
JsT4Drgkph9Rx24tWr9XWJTZOg/cZTDCpu9TluVJl+80CVgHa/CCUwDSWowheGLg5PD9gRLZ+yha
CnbV3wk4VF1rPpSvtGGfGhRbnv3sMKGOwpJhSR5HQ+gXkT9PQg5q6L5qB+8LwWChIRiLoepwg51o
x4W3Fy2oVVYCKlTOa6UADwwa1ZEewq4G+77GG1ntzrGBhadHoOawsUNZUzQUs7xU8ga2fKTew59s
Ud6s+hZTK+G51obG0ySXEQ91iljdLgeSUS2R9m/2qp3ZNmUBkGzya2FUETVfydVwyfIQXbUEb/V1
OVH1OU50H5aApcu8hoZFF3uMS6mDpY7ih6X/uBCDlivfWtn5+l96W9ooYwfCWPR9fAbTNVoDvFNr
NeSfsEMnfXZhX7MbuTS/DYKeTZXsQK4T0EVOKC4N3H9R6vsEeN4YJ6qW9WIjBe4xAGgiI594aPf7
zu8tGA3to0eYOapzT7upLHsF+bheIMEDlAgz0LJ+K2fhZ8JN6w41x0ufgTCFrZl6B21/DO/bfeKm
q8hw79uR6ej1CTni/Fq1YoqukSdtB4lkiAjHxQXMZ8OPaG/UVdPT2TqjCo9c+srbiA60WBU74erW
6DGEbyuC7Mgh2HvjCNwDXhF1CMoKzqw7KB8pgcF/6BNSI6KkesYAkWvIfBUNLsWs5nfcWGYJzrOp
/nJw3Cu5wHWyLAD/bfZ/UeDr3xd/LJjUPn7yJwD96y4FBLH9lj9kcn/FK9RK6hdd2hbZVZSo5cGy
oT9DmHKyo72N+BrW4EZxD5EzKOJH+o3G5Yr3P6r7r+gvImdckxaQMYvcL3JYkzRp1DhJBh0f+wNA
pToC6jP9uJzUMdUfwPLfIf20dXcEsD4xybo457EH9e/kgV24+d2N4YttzIg8P0iBAYNbABc4X8rZ
Jhxh681rkRVhgOEfCk5snihpQrCIv61KxRqMow3typxmmHAI2IYlXFTn2aUTZqZU6ZGyXA51C7Af
UHkzkrb+TwsebfitdvkWEZ/G/kNHmD0FZ6I5xTMyhZWOo32N/fQki+LxcdgWF4vqQRPVmefvvvn5
8/y8LrhzZBej772orWyyeYirzzTAp9nHbHtKB9JbU+DWpQ8VTiBGrINsgaqqhIZ5wMLSXvmUcjGm
nIoLXHcnpsqPIPntceMVnwc8ToCX8MeI6Y8LddActPH6CMILVx01i717SSbtYMKfVgfojwPbd37D
pHomRUYMXNN7eGRzBNYUAYnec1syxJEUcOVqXg2xW1AGrKhBsnncTOCLP/OR0xFbuam7iPDjsiHc
87i56hHlSWM+ooeuEVVOouzbZOD5UO8fHE4Hqed5dXndzxu/9xtehzs7bFQeJhsyAHb1vW+7/QNE
M1CizkVgJMxeMl2+8lK2fF6BGIdE1DfeLLbROhIv0Dpp0GWaSH03jMF70PRyNA4sBkqnYm+jwa3P
lgnRTmnCq8EZAIhmJtOnR8qI7nczgTyN255fnX25mGg80Psj64RTWh+JB87JI5/ZBresMZS3mgK8
VxOpwiVxaPUX69LSnqvKJj6cevpigEdHK34A5fy0OrxOd8VPH36svxp/C7waJrH1Ge1Hw1uYMo33
djGO4DflJYOMoyhO0hRByatpjjBJQGi3SAzBFPw8JFTypUbrxoxwYioKv7QUvAULAsBDsfIVXCJy
6qenbEBfmBIpD7ux3J1pnn25k+LxIqIKLDSVpFlKOzeJcG0mT++tJcyeZmBeve2fiVfPQ9DKR6UY
OA2CuumH/u3dV84ggjQ7eJ1pq28hCoh4KXpTbSu2nsVOCsaVkANSMfB381SnvHx4/J4fIz+4Avr/
Q/n/PlD9eoLPA6b/E/NMdI39q6YZKFltJvGNoYkU6w1fJ9+93Kz6hAmSoVJ6LaLiDtC5aHgP9aK3
9hnZVLsIj7tjFSrn7DL7oNTkeOuD31QA+K3BSwjnt/lbfxLWDc23ydWfOX4h2MkjshQP1JMCUbNa
f1Eowq0VvgcRjO+KfJLO4va5qKsfEIXvBrMsWz04yS0jNgwHIogDmc6PdTAJUQJzjX9n3i9LM+1V
Zg9WWIRYJVqkrNBQcFGbm5ew8FlHR3b85pFeEM7y7rnl7cU/Nb3d28+VAVCB23MI/IO3YjKKjgIz
PJql3nZRGjp4X2xiQl64UdJWmAF1Y0+de80YPRnJsjwLcF4rG2ukIDKjyIi8vTGKcCfGcQOuDKC1
wPzTJmgKeZhqpHLY+UqP974aV4SoeqqM9HBiTxesYr/Sp8vktPaXAuqjMB2GTXXCz3O3w0dY+TYp
2dF0BStHjb8hWY2XqXp3pGyrgnwiFnuljYXPqLzN+KKg5Fu6+c1cZv0nKPwZI1EQ7b5vAHgWTSbz
W58LU+WXD37C6FqPjhM7OUs7TCViK3v/zXqg2AGoFfTDnfQRsg38uj0AjBkiaogjHgWnYaEI2f1/
bgMoebxsYOGLAu+L3b+1uUwcazWVrPhpE0LPMNxsWgXYsHibcVji840n2eilpgraPR4QZOgVhUEz
ksb+Wr0K/xe21cZR+I7zXBHK3p5uct6AA5n+uRtnvAokw2O6aSSF3nN+7LQtE0u5ieykcCe2oL6h
GSh9oCOmLfXWuadBan6ma9GfEhtBxnQQ/gjiT2cK+DAzatHxCpj367R0Lz0dmE46FIyLimA4ulsM
6uqkJUWwA/d1m3kVdIdYLyezz5ym0ffoCkSDqEyqdOJWhSw6VwnVt3Dbdu8ueRcZU1OR8cLf3lMT
EvQdVqfHE1MTSuncMhWRZS+8P1JggVHN2IwLwkwZer+zGDcF8Z0yb6kj6cVmwc7G2XpSmtcl0Icz
M1ygnORxZDyEauhaa9vqebnkuxvOqpo7gUF6R+GMo94LLpooIeu/hQd2IUbdcB/cLzGofNSw6PlG
RpX5qx0Q3WnnLVONOXeIFCazktJXkc+x8B5Fzp8RC07XEGnWlvsB4hLbtlcxBW38Z7RfyBIGouFs
XQCH6z5WGEaxN8uIrPm4fVzBHImhO+T1vLFdzw+KEDvtFGn1XbauwjU9SyNqkbh3KtzPnp1VrFJX
AqQOIamA8JsQRQplXfdtwPxt9UCsVOvHqMZ4riz5MRvTfUDCu0acoQDn/Pf7tH/mNfv5RQO8xv8W
tXNhKnB5z+C6YfSDhyBQN8MZvdCNViB3s+2Q9gUDzPq7WYyR2Ye62PvSYZLlCF5l8YGM7jIRtH8S
LoRVAPv8zJmja0CGGRLpPBSQuOG26AmSwWHYItOkAUZULI/oGjeGd7L9krRlLqPbGy1/kojLFCuL
if/MA6yKtPQ8gcPsNStgszUQT4Pw5cOOou8Cwyowcf6AhCAAZMncpN3uLsSGjGgvJoOURS6Ip0ZV
NdUxnm8JLVyOhoQQQ/QfQMFqacBKZ3rQJ0bb3lj4Xf6e82LiLaDnli/imUi/yBQ4V7jnLFtUtpnw
bKHnlpaVBOKSq49sGa6qKyrAZmbVH6M44SMGncvoVE1WRzuGHIcRkMg+rei83wWXmvecQFlpXAYQ
5Jbv07bTpVIaBb8OVY6izTCiHjZ8Ll79uOG1Uc1Chkt3JbD0WT2WwLuDipZUr0mDYi0MRZakBcBT
HgGCyLvnnRmEcsDX6ytwEDXkeaRhbSVQp2XMQyYQzQVVDWoRnuwUaEng9fbhl/jBOCVndXPymijG
ejAmku6Cj5SSeOOmFyCnRuSsSzdpI/d6uJzy4bOGvLWG/b2q1cZ9+CktcSZXfcqsYS34JS13EU5R
BLmhot6b9OG8GZi+HXnvQn5sdPtJn4pXaGdh7tfV4L4EcRd6ARBAkXAHbZc7ZoGyGnP8qA27juBv
gZ6Tw6M2vEBfaen1XoWqyW5cVvH3STpG2CLgPGkhiOaEq3sAsw+FL8gZ4s5Nr/wCE4/QSqxsni1J
X0Rv9qIUKIHKsdSSWdnc7lAVfbzWyvz09e2kYOQKHgxd+Y17ZNDbP8OLKrI85f1mx7MWPg/0eTyf
QTPOI0HTut09UbMcmjbEwAbzYx0KAXSUXP7SYOI1LfLshemQf0OSt9RcmB6VD58vqmAJV7viENiq
4r55lRPk2W5QdKGBM5r0gbQ0nujOqAkVyKDy8BMqeThgjIdhCFoEabFWs6JaZsMMefbxjBJlQEhj
/TX+8Q7IDckMgCtt/fiNyPgDfypXtNg/eKINGULgokD8U45wsedl4pWPCykF9HBk/5tPqL2IFrUc
SepYPVB76LLoyYY1u3F5r8KNbu4Ch5p4mvCL0tgZrYMj6BqxkpKU8QcSsQTlzDp7NrWyJyhBj4tY
JJKycfgkqwtidn4KHWTNJgcx6ouNHc+qPSS+stF4e89mGbPOPr07gF0mEQG2tpXqG3LS0xwFyME3
QcOwsCKiA7krtsUt5vDuviiULC0p0cNeDgrSIsrZK9ZkcRv2BlDKdMb1tApfG4prL/fe0W9/AqQZ
D/QETOGxiONF8vMno9jLaaez2AOoTdAWKP3cbF9i1Anlw3IUNqiRxDt9k+QuD/tNfqX2FCiKbDP2
5Xtk8Z98vC8M1XZaiWMPMD5g1aUs+TQG0uDcvOW23vNvhcdMp0FoE+Mmxw5F30Wrz04sfok0xmm8
HA5VcPEfBqg64HLs4DyQkG+M7OfD1iRK1vgyVIAozmXsMF+riipjPu37JZEDUIHcRrmPeULo5D4D
ozEf9C/9yxOt/nJC84M845XzB0O0d3lPvPi+Zi6AMWc0UaEL0GqwUGGgf9s1Pi6UdWSFYDgFrG1k
tqZXsMnzFnb2d0A/DXS4zkb4I0+0KPU7o9PfqFO6mperiDAiNpYft63XlA2HJ0TUPNNY+AvydKDv
eaS5EK8sFZ6xZuvyJdlqGy4fF/4YbFYOPv0P9tnEfnL4iglgEhCrCWf3E1yPDB2+Jz58ulLIWlBT
6HxtO9qaFTNl2V8t+vrAcq5bjFHY+B/eNzPSNbGVLj5KMYHiE9YMmO02JDmPaWx+U5dDaf8gLPXK
wKhUZ9eA2EiaDeKwDl5E0yiRtvNkiwhRMTCUhwStdZ7a77slS549UE3JRoONLgsCRXfxJc1yENfB
D+P/3hy9ne0FfYQMUJSaVBWQdAze8s3R8oLk7BHxlhqdU6U6+XK0LMiYjFAVNIWqbuwTbq3mkZ8X
5p5RBRg5hYbq0Jf6qU5Uc/sqx2FfjnoWHBOtIATsyMhSXlw31SsvTLpMxzwAaalW/L3R5YidlxiQ
oZvcOIqcFn1EETkQa5Y14IzUF9HB+51m3t/n55P0VsPL+guTkihKtsJjc60spCmDcXantE5UoQMH
+Ie/KktHVMp19HiuB2f2HvLxdZz3Wef8/9vvWa+80uZlMVKr9eN0b2jNDMwSqaBX4+AwhWGQVmsx
3UtVZQwqN7wOn4+divENSsaWqYe/XIC41/OaZ4Qyf6hcA0hO/r53HJd98n7pERWGWfS3/3S04cJr
D7JT4Ifg4HfPu3IwiTNnbtFo18oZy8n3WXbHFhnMlx8mwg2e+zRFNcf+TN6JIy3l5PIza67fGz4J
EecxAF5WRVUeGmagiB2pO6tW+R0gNO7YmKXdMheVp9/hoDBxQF1sSMStfFyqncejSyalQnFK2r8v
KuG5m+3I4vBloUUPXEg1nK85X7DGMTsbmNa8h8eCLGS2vW8zcq/piepVlKWMmMMVWvndMB+LqQG9
DEY59ZSv0ewXiA0fLc8b/i9pAqv24eFuRJ0z7jCi+2HAZRWWyWEIkXpXnyGp23KA7ffM5KcAJyQj
bGHYR6/9KxdDgyJsBum1PEntES6U33gr0sRKxzZS6q/coVAcw/P89iFZFPbvYfqbBfHdBYwCRy6T
2no3zRrlk+HkQX50aPH/LqkE3rHzdx9aDmAVDItDqJhSdvhYi2fQ/ys2jjfNR92lWhgkjRRXlFvs
MDbXELVA1BoClXMTnOr0an7oeb5QsNoYOR+exCUF8CbY8bl6fT6h1MNlH/VXEWF5Nw2ypykjsY7b
J8oTqADaQzF226WI6GrLR7lk/FY9VG0brR1BbcZ1t9WBtrfwxzQqBTOTCamydu5gECOk0b0iGGgk
nZLlHZIPK2Uq7TI3h8Kd9hBki+EzJOZ/oLgqSB1xEvXj1hAE7d+ne0IzrzEa7yEqERdshn+fI0Yc
f4EgdB9+QqELTxm2pDqL01w1GMVGjg0KeXyRwQmdzkMx67vGHhpF77LPWxOMAuj3TE0qVYMMiIl6
pKw1JTVCYunn53xBITxTC9HwYBa9eLNwgxLkxzQWWpGZbJalEK9KW4b/O4LssuDAYWseaE8QDhH+
ByEpRbA7q0xHHma4STT7ee8W3usBjjsPlaY9L1DwRGZVFLQevMpDM7IzbwgUrB1dMXRS09zD4gfi
iQQiM7+6RonY6fj/BLIDvgdZ3JIczrzSdmg7zvXdC9fyS2fiWgY5g1ID5vUFX7aoVDhYGANG817N
WC13DTICYkvEm16vrYK3/A6GIzAUWzpqefPlhcsw7cxUpZqewS3EKAfzFQto235QeAVc79tewZoM
SJtBfiIOOD5BBNwtqWONTR3YWYlxS17g38A2q+EGBdySojJZsk3pHDLwwOTcPcQxSSFpAFHwMUkS
/cmdick7kyOH6lYmEVnlhvF7rVEaGnXUhW8U0LQh8GAZMeJG9RY583ZpglY04rP4VieCwrximH3x
HmTEDb3ryBs2bQQsSZ+RJCXRGrCCr6YSDDAIIoj5F0z7q8/x4VBl652G+WfS+AB65ONNI/ci22rj
tmJndj/WtveITEY/ATRv7buG7NhSEiURp3tAob6tv0kuwwlx7qZSskSPAIPmyWMwDzRN5ZBPaRm7
s9XBaVpsnhW/PDsf3dMce79BoHgTShtag2uLvqVUXVvTKojmLU0rXwuDhyXCYapuDHUgHrn5ldPR
iomrzDoECf2ax+st1SWiD17ejxeEi8cQdzsIAUZSz3RTT+c5ebcbjcYwgJCt4H/kdN3EcJqKkwP1
QnQQy5g5IT+Tdzq082hYVc0fW5nMpxy2GGYw4YmH4ac5wBkZsjnhVyYvX76csXKdhA7FtyWWGe+I
jn2/Zfp33U6B7vAe3WZSYfbZihclHfUwGFmuTwx0RrSIRBg7zFe2UOjRMXew6Bu+MnTXaNU3HOo+
ejb98nMCi88QHgp61ObebqN0PmDXWLSyz2KzrF1M0PfpB9SF0W9DVFW9YFzDb+Twvx0qUVXIRb4x
+sWwAzyqEGj0Hsv01RQ28GziGvYgdLMKL6PLIUTi1I/Dd+VzR2NF68LSX6DECCU/VBQwWurqVX4A
L60+xnQlw7F9IsseZMXtL3ItbqH6DOL0fujDUkvOwxetF0JsDJycO8ShWi467P9MfYbg02UjrZ72
Vf4BQq3Ceng/+bw4MGwBWiAulv2h1AEe04M52CoAJaiNHcFr1TsGNKW74bGuMU1gknOtW3mZhl60
DvYycyEtL0JLWc2XXNK/NiJq7N6mJ/xYTetjsHc24pDPRA7boDSdr/STCrFb8JkP0imYkpk3FzkW
sM1dAOrAHq7gJWPSgHfrX7pua5CZduQCFPFGs0MRlP5A7JJjvkVULr8n3gHprJ38Bkw+A+ABTcGq
f6skQHH1Qo7Xk01FjhTPLrSFmgn3vNCV29pePjMHJpsWil0YLc2gs46WgImJJhMAJJZtLOYZ0fBm
kTYW3ADmEhr1HhoeBTT2CWl7jgwLyxkuxmOSG22UNVM9hyz3K6CQNtqCNCDchWeKAPmxp0TPxTU4
HvYcGEKfgbnTAj2NSDW1Kon6hvVIrtxG0C8v07ipDB3SWHbGI/n6J+UJ8Rsk1WmWpT6eSjIeXLn+
y0B/zO9sPqcGb4Hwxd2t9dS6rVifitAVuA+QfwOWNwJEAIaM1W1iBXld11G1qOdzQzyhhUbBpa7b
Q7THNCWHDW+tXq1J2ebjqg3+9VlgwLAL0qexcSJV7F558FQdgKwgMdQXTwmOHJSYFKUlxaRButTY
DBp0moFAbEH9eoiHEpIr1mh7bRBVqno3BtTfA3PqrG70F7/LR/g35C8T64WlhXNLAp3rpgJdJ9td
+xCTWhXjryLiQMCT45lxHrJ0Efd9p5IByH0FoyzzronhAmheqd5xjzjQtn76wVc8m6P4qWrO7j3P
pw+V58meCKscDeXYap+6LYTYvCfTC31UQmg9+a0ou0S6iDJYe6laAXQD+M0DSKy37O1MRANMx6xb
JBIV9DzMKJc37Aj1knbwjxtQtfiBgyJobbFilGW9S7kzX9l5ayI0jwZLJJoqnwrRDtLKbPaaT5Sg
I45KETwPgR2jjn673nDBlthrn94fso0F82GNlereRx8ojZNtMpsfm47LestlCppS8xg2NkacPkbn
sFfv38gpyRA6BWrEuQcUe4AT6WlnjfSCyUuFwkaR0D4lSirXNNQ88tTjRtXNAFr0YbJMhhK7tBDy
2MHVDUitAUSbvyRZL8s8cTz6AwIu7+YlCViMYBka2RLh5hiZsXDZsa3kgLBPGvuKZ88PgAD3/gYm
8za7/2Z1UMlPKUVHw8rXGu5zSEB0nNwfzuV/JZXrdS5S7esf5SlW3yKVf3Cu6I/kCIyA0Q2dr3qn
D2QLFgEATQaAYX4Mhkve4M1ul9oD9VIawsF4N8gHlC5S6GumKqVZ/AzUpjQgxin2WHqZFcI4pk6C
q79DlVtoSyMzMwOnTTI13GV1Yl0K95yaZT43kY1jxgIbKVgIjniJQPQHBtJZ+lx8hC9Abi59yBH8
BZvh6TLx1n6Vx9pLKStQUQ/MmYdE+9JXIiCC79vOcgSi0uID2spaj4g0yYGVsteugDKBAjs/WKHE
ly5CXAgpEGelZB7uoMyz6acZR+6XeGK6bSjuooJkrmMJYZkYIh2lgTIGkrgHVcMUlk2XrH5XJUtF
DwoMPzWN/IQ4TMawHBpeBlstve9sS8PU4vpBva1bfPhlKeqN14cZJA2NIyKwEBhjmQz12cT70buD
LACG2pqz3rWf8iQb49BhvPcbqovyKuH8LYLijszNjvW0VDYeN2X3epmlqcRu/cA4S0lm79MLeqTU
amxT1Yk73sNV0vsxk0yR+E5SWfJF5HfbpxTr3n3BQGx8dgBE8k3vOx+ZIKPm8w0zXcNMBYly2uKP
XBvGQJm2ltHqFj5fo1ozbPuu2K/Rdb5TqGntGGioGO/s6gGw4O+VTrDjNUqkEaR99yAoDYEEZy7e
G0OFcdpISHLO4BspCOyJ69SNtUEh6RznK5y3wTHYnIaDZ0fP3Qr5MFrwJz/zrlXp1UfhCBMiVFlH
VIrmopWpoQ7O5GDeqFpTx0IUokEwxXOL0rGPAaQqnwsyGZ6LZiIrEwrQ2sCosml8piLBn4B3eeWu
Ok/h1ak7MM45Wv6HPtz4aTYOzVJ60t9ttATZmkx1rAdq0urjqqcDk+yB23vdnyi5PjhheelFrsuG
iD/pIgylNyqbgSyr9/e6raBWPksLrop+zdpmjycOlIBh4BYXEFEk1W11uGwB9ZzN6v1spVYdQBpw
TXX957kRPNN6BN5XcjLdT0SMQLjKiCV+k7JZNpokCmh5bPtqaSDH5gUO9E/N1LHU5NxIKxL5a2Oy
V0Oz7Mz8oY8s+EuIkee2hd80H13GkJWMEl4tSZDDwLp/8l8FJZgKzj+0/VG+7zFYl4CFKXcucHJS
hQLLq1AtNQ9QfFPUjpBfDrn9vjUQqnG/pJmJ6A+RmFbgEPvIfmjtOhcZYxmFCdU04oOTXl2s8PQF
FXU1oLjTPdlSy7K1Q3UcSWeeBEp3qPqaAD4h9eRqbyXqizBqEsHpiz91L1o/i+NcVF4DVMF7j1Jg
uTli3uGwyV+zv+hUJLmNGb+OHFw0jX3ipAtNLczAmVl8FK+ZCdaC0k8MGLDkz5pCYrufgjGMarAT
+MytGtijCDJ3WCZDubTgye6QO5vJVBv3oGaNjO7OvYxINh6qnskB3T/UcOlSv0ph3fsGlPlgcMvt
1L6EopO/8XNFlND0DL/icRmcx3FAUA3CTseqzyYh0zgSTHPnvjmppaypeZiIpqd+0DFI8qtJBw2G
/21teJLOUY97/8Z5RWmFwc1haMr7H+jy8HoT1lsg7eAdmLXKm3iTGD1KOgHtEW6HC2N4uHSD55op
UhUlA9WJD/pozqQOcRDECHaV3Z4gnxF6lXb+N934VF9gYTQfHILJrFQUpgm3D3BqMQnIj61/2WC3
SkHkEMhyTZlx8q5b5q38ca4J085MLutUZel10MungW4wBmACSW1hjbz3j9M/fAbNRYMUxZ6D/jgx
1nIeH5SGghHUL77sVL3w94idu0XiibKfJBTB3bH1MLfc+zyspb7GmUD1YyEuiU0YzljoizEhpXQx
4ULT8OvKQ1K1vMZlnMulU2Fy8aKMOzQj2p3gK4vyBUW9djOhKDVVcMJeBTWpkUaKfiVNcRY9rUY4
FRlmS+vx8j/NArWX3AywCzxFXC3PWoX1ED5dbSeizBNxsk8PRmJiLFoYYztKViV63YxDfHxtD/gP
nFpcm0WbF4/3Vv1hQecqp5Cll3tGIv0bPNFEJZoQW3kHh6/gtGUxo+JCC0wH7glUi9Oqh++jszMS
lBVqJIN2oDTLt3Pm9PI+XROHOCyGYQkIurw/eIT37NuF0MHnu7WsjOB5ddFJnIS6Aojr38xUfg4Q
qNcMdFAF74fLInzRB7CzsPUwadSe/gMtOLgD/Fv/TQbwG9dBYsJAwhLCG2dDQw36h852jYsjjX2+
acA3LPSc5fXdnqrr95tz5OzvPq7htV9w5daBB+rQ4tPvF8ipdmqRnFGT3saQ7m6pLfGMmcS6hSbO
DnZ8xbTjrY9x4+oES/U36KE66iFw3kcx0sVpJ5JC/9H+UuOjzIsdzkL1dpJyjPGj0xI7kFOKxJFm
Q2RcoeVbCUlHms7gSPYW/dkM8KTevquVyELCpQlu3edlFyi3Fgc05LP6hOQaaYugtxvj7KY3yuBp
a6wLkqNwFuBylgZcbIshlX2mqPSUiyXLqlRGv9NIRCZPF/wBf5ptzZoBPXOt8pkSfi/dIUHTvgOu
pRVuCMoJfx1rY1QN7+2PbESaS3ILJvXlC6GJB3s/yKFG/3wA79VgaKwuOj3WgLywcCXpWtaxZgGq
78aWKW1rCsZx7kuuQcPC7eT30Eu/t54ruxm66sEQa0HOG6WhurHnHX/XPVqxPhKO+nfdlDi1TghS
rWOqYnBHRtOeoERU7pRjgBSl7lUEFMFGnJMSI4FeIQRVuGMlTUWWpet2q7sqyO1T4NyTm1Ualo1H
2XNSUkixpzD6tumsDXi4Yhfn/fj2pvv5Ze3nu4XavAMTMDTuQb2I7vpXmkeTDbdzPXH4LNbizGBc
Wj6u+JDsSnRVlXkzlc5FFRlQ1RkNqjGTifXwlkx5l+5Tu8mtRNsPdg/VD2/PwNgO2Jk/jmtr5HGQ
bOHampHfNCM3gE0kBy4h/zSLh7i+4YW12bgYaKTsHJdGsfTsj3HKRi60VRdRplzi1Mm7sndhRdPf
qx4RoiFhD+cnneFtjwqWThWuMkC+KYfD+0RmHYKVkh3YiqkQkOE1vvEdzx44UfnPjCmPU6iHhq7R
7NPhPJsVpphfpqkAYMntElOV2H2SqgDP2Cbe2srHKGOkijJH3NhYxhLcMd7musPDEe4jS4vTVm7y
j771vyYDUpUsin2ornANBBlTzatfmXLwlxjXt+wGBHKm7pZNT3ZKZb+j+z+uyMPMHuQKmNkcNp1G
UlLYwy1zcJCG9OWkx9KfJ2dpvizAM2kk2KSvXL0Emcav7hpVxGU0rq96hlBdN7kELzUOOKKmd1Vr
3JRZ/DHe89CUFPb8jO/ZwS8QmfkbAKiFBkSz2vzb6BorWduM55FtAZa5NbiaXSclfZaO0NGW7X6r
+CHYtqVIB617/uosm7s9T7Rku5SiwfV4mhWUiaLBeW6lEFG/ybzXIzwQKLcW6qrMqWIjiUaMBCU4
h1J+dSn6GadSLScKCq3ER2u7R85SkbP+05I9iFcE69p+94HMduXfgB6Qde5Gd3nPTjWYTTjv1h1N
cppYjs37E5qTooL0T5g4zxtxwtkUFKp7TEKCW0mnogD0xeYK/OSx/lJAEV0bgvn2BuhEC7BJAMy2
0y3TQ0q4zp8DE5++06Dqg8RPaDaMzrXE7tnIUX6FgXrpEAjSEGXyxY96nqvUHETZg+P5CDFdQDUv
PIf/PXdO0AnExY8CZx/5eFxmWmoJDbOBldLXa2I4oAS4/36fyOwmYh7WrMqVkCxrU8r4sl5EhFas
m8mttwERLbi/7LqSYXxUUUXObci6Gk8S/3HlBf6+oEZcBrSaGcr5KPHoneHVjhk5HAGALyFunFIQ
l1tuR9l3UTrknZpY5b3Jy4UnE+Hbd9QdECzHvpbBEstjiTSVxtE1Aoi5Cz2HXkny9pljA4M0AD6m
5KeFOtrqrk9cc9auCKU64NKnxd1ZrJfBZT+/0AO4YNL7JjY1uYrVL2p2Z+3wN8ud+gA6N0mLDMi/
VA8DO90E6Nf06NI01+SS0KTVkWIZG7jEe+lWaCOyHyzrtkQPfZeppGIKXiLm4WSzyHcGp591FJtd
uNOptMpnAXdolOUf6rDIYxwasiJQZ80Kbwr0kq07iELIXpgTOPFt22HLStvxZQpvMZDA17sOpFu1
NRe2hE/Mongw/vfP3NG8E9kAaZNhFxT5dosIgTv/I/IIyqPD+6Ff42r50d1A66VB4Cuofvao5SN4
TIX1J+QDo6U+NfDoyOJujL+yYJPzBELNinXhTjNiQNN/jzVkV3oPk/ssABvvGRUtS848BFEOSjQG
S5SFHphmoTgKQKXNppEPs4YR4Qt9okRWsg+dlBrInPhBkQA+yWY+1cmAGcjXSF17KjB3ol433ez5
D3ZanIwWSMzb4b7CdHm5lWZTzT2ZY/SR68duKk4L+rYxd6vieOguGxxvtCySVC95pypM//SHzY9j
pCKBUzYgynSPydtqxZRU3+uryCiNo5hokL0SRLF0oyof0/j29lq7WW7PpxvCrYN1Dv6svCykBvCk
WUM9kp5tRB5cp+uEfw2flSkxx1PTEQeiGBk4IM8K0xuA9UUMRgSQc2O/V21WD1WqWtmDH/aBIUia
W63heppCGwtLiukIwGw8mJTKqoLr8UJ9pw3ymO7cRiNbHDFCdoW/Ztf9YiAyqYySjRaqtqBhzvxI
G9W7qE8PhAmEXkgDhl/9uYCtW4LuD/dg9NZZH/iw/XecpAkGtl/v/zpkfogAr/V+aDTGQvzCMqMj
10P4FOe820foGDpjEAzc17XeyDZx6TgCghOprz/EZfS0INEw/WJf/ZwZ/ozNpNHizelH2/wUlOV5
G1EpOZEC3cto806pTfS37bycGgYIp8J4zbIfK191EC7op/tKurp/gIWHGo5JG0ieQbfm16G3X7bO
z0P4CNNqCQQwhwoRK2ARkNaPw21wraKPQ8dP/Fd/jfawfE0DPS4vAyzBbMW4PkwcTbO4J7xVcm+z
turf1h1vhDcdwSudO3htzVZmIOf7+QrJp0GJDCpIjeUgsJdsu9Rboqwd6TSihTcd/RxHh0BECBXh
3Iry557FQ5Dl4bWw7v1S/uDW1MQnKMRoYkqquFYNG96tUPKlW2RMLKi+Au00zh+PiOmQtPtGYAJt
BwWlNWF8aYVSWCni2Jf8/SrhKVTQmU5isGnQ+BAECdlOsqwgmNx2H05CBzd7p/4AAZO/NYrrnCCu
NYd1tijxnkDG4eVhUi1CF9gPK0iJgCEwzy+E4m18gfZAfWB65cqON2IrYb1zjPc134Pakh+ix7PC
HwEQTktG6w3H5ZfZQiouMbb8+j7DqdnWKJoDHIAodFItwFgj5RYlBdAQBxFg4bx9pQs9I3O8bksl
j3wKljPrcYTD/ihUjDTpFx9qX/NrW+rri4Jg5yo/I5wwSZwHLswJNCVTyF0xWKt5h+w671nPAXlB
ZXQ+cddE/6hrQ9fjLGqftYCZpCESo8JKod1IlZ8D1omJaFpEzJtOex4DIRoSp79AxJHpdiGFjNqQ
KOEWNq2I+WPP+1Qh3FCgHIbHu97pQYg2z6m7j905uzFMpgWqjS62+EP7FjyoRFvV7eoqfOuZ31AZ
5WO5KduTRuKxrYKPNfxumps/Ng3Xinx5Eq7cq0iQLXU4c5tzdUD0Z7Z3be6kafwuuD/Y66qMNPSi
p+10nTII64AFSQiYiYn37dbw59T6WXTy2swkJaEppuH0u1aExduH+B32OWPnud0K4X8EzVVHL46p
NEvFJRGu7FRF4cdkhfgQ3IUvVqPWguqLuVNrXSRazsJDz2BwDEl+L+R44qUMYU5vp+4F/k4147Sa
LwgsZpoy/QTU3ffKmc3Xepg24HRDW/2PynYhjJcomscarfOpEf3UYpiEEv9qb/qO+Ya8NZsquQko
JZ4KOR4iEVqURUyAjUVNN+js76cTYEj14VZK+6kK0MIhbc8Uga2E4NA2Ruk5kB9QF2YMN/y7Iya1
38t5l9FDg9LrLkn+sC9R+CTFhGpGwLomrt5kt7jtwk4MOTXYaQDLc4HLAxMxC7+Ky42fJzPW84Lh
XOHVV98WsCcBiAE6imMT+Wr7Rx/9KCiHj0dp9Ot8Aws4EzGgN3S3lMEojx9H5fYElwy3g9Dlw6fn
RuIDF84YuKma+27svE/9rsso9W9zlUlYT0xGALJQwfkIfWqM/stqqyvR2LkL9+MRGcaoKPKEd6Iy
Y+3SNB3lRwr5UndBvpeEr0Z5rhYSk6aFL/ZrkWP8vK/1Of3K4LBciDhrR2/CJx9GqMx3aRaKcKl4
zk3nO3z30R3PUQxDma9gpj2IWXq2uvnfxv8DB952+nmUZTHPbL6CxGuvbvB/Hj0AeXo30fT0aF8C
UTFhttmnMEzg+FW4vaLZkmeE39TWn9OV4X2IODJ67HyW0D53GFaTcGIurAwFFZozFyZsswj4CMQ6
wITyfRH5eNMZXZQPxYablpOZPmGKXxjhvGSj+Z1K0qeVoyIKBzsqm70xOFvutJu6k9E1Z2+bxQCD
9wR5rUUUEZWK/5VkovKdnyAkiyfqDpHI4hJ49BrB5YnVfnkGD8U3k3opRN3o3x8sApvGSq6fRnCx
xZQw4Ffpft/4ohL/vbSXaXFeaeEAThZGKA0SURvNnJseM7778XJpMNt8avkcEVxYQVOsuGoPxmG7
YYAz0+X/SiOl34/s4rQVzWwCFc3ixwqhBH2U3g8Xr+8xJ0f/9Q37FxDhh/X0AaMbvBMgykNEurB0
22r1moI+Br+mZGYaYnziqDbHyXyRtjj2GB7wK6Th+vrWsAUo6EEjBWELbvGvhD8DacHmic2uEgsn
mHmK4x3a7gGoTH08JO15GlURzVOq04BUC1pvz6r0MGjriJ22grbsq/Vvjfr68TnvPg/fqFqQMLQK
WYOg09Ryp5mQ93+3S6rQETu8PP1C0X100tCHiZ6pk42GSHbml3qku97x3SdIe/R0QAo99CkkObiN
f7tPXduTboCFLA+iqNcvN1KEUZf08zb2LClmFC6oHZgNOZelpuTz1Ir1GVqqXBdlWt5x81AXq8Re
p8Fq5krcf6X+FFNPyzpd4pfkXDBzj6GAAKQYUeZQhyD3h+nEym4oXeOu9ZwcQr7uo0Hw0CySX2yz
6ecufxqd0qPJ0K4B1UbU+Wp7uyi6qxkdMm3Zkk/g6SNfJT5FhypQsOQaT9i2iCdss1wx56qZA4rK
JW9Vmih04733kQxGHtD/P3m4JA/JsT8J+hCzXHnTkTzymFkVNnYP4408uEdDZvYttVHPiNVzNXj5
1//pBuZUXdt3YEbWtYQ/lBR9x8A579FREmd5zpcRf5KxwUtgpdK58ei8bsLq3JK9h93AdvXBhO2k
s/C3ktHpdG0xuRIPGY+8ybj0VpVFTR4MOQ91wceoL2LXDWZGck2L8K/cpyLsotDIdoi4OL3P9jwx
g/zAzhL5FbiU6+TNcmiTjxgSrlothSOhVLNsazE1lESNUiDcah/DH//JtdcWbZ8eT4Xzspmwol3A
1NXOwJKF5uUzh93/urVEP00/wBdSyNFEM57vclMd/+37tbHAk1Goi797e+6xQF/n3wWeNJDaEsrY
eGajHah2vC/p1EZhjZVu4sH4BpFw5rQ2/EyzbbSvvXbgNc5n7hTJysfo58T+uGkDan1a+ku4oapQ
AFq1lk34GvIjaMKKBENzgtqOy4QC6bmrc647tiYGi1UUnPgG81Tco6vynARxA0UHt968KSBfwzi6
CfmKgcwex7+jSo8d0nnLRHWb3t2KWttqlty60WGV8AwE77i7UqqLW0/I+ksDw0M0bP0qg5xRxZjT
FR5bDC6blcGrB2NZEpviQg0oDs7kSq4D6D77LhOCqAlT8Ln7TmEe+aC/k4eHbaaGXjb4LC6KqxAN
UVpRgPBDkODBxa60Jo2JFcwsVbpzLawUeiPkapRKaa57bl3hYAxivilZ/kWEs75l/MD5XWps8oaD
grwt1kFQiSeyPOhKzApHBnBOoFj7LQE9YQZyq6gqMWC+aafiPcbD1GNfZ9ITw8vWoBv4mQ4SXOsJ
XKUhZYDiqitfbqXtNZrCqPKujrs1V1oLO3u3BQXvcpbU3MMTSmUfAIEoqXN3CD/1/stXe01jLmwr
9O5IzsfxlQKhVBPXMt6amn6jGG8FoaV81Fcl6ryGrY2niuo6/9rWgC8uoHarYq3kkYq6dCxJQfJZ
vtGaLwMl5XQ1dnw2Zhee7pt2YJ5+7FP7Xam2OuMTYhQMAJUEx236yKq5dUwKzIVDX93Lb6RQIPXI
tbS53yOGngxRl3ybkdbGw7Nrk8InZGl6E5ydnmCnzWgY9fnboXzc8RbS0ltTpHht2E3ut4vzZaRg
t5QV/U8qQ6/O98Y2zp7COXuLHK1rH/QdUjvQdAWkbE1mFTDzI3xafn4Lq0kDQa8mkrWsJPUhxEHU
xNQQUjOqIjG3fcUaatEdxUWX0z1qaq16WyvieWSMYzYplLpPeGmGoemBiJX+sp5lYVzjNa/YWXXW
DrYyLOVOViIvDHS9dPb6BhDFHIWCKqU/n8jdTp6su+amfQEnVxlKbGRjOIS63xH2m4jbwjm9YnaU
xrT/xLT8Gwf8LXBYYJY8sTk5gF0fL5yu5swap94OXrQGte/i0v9tTMjxZIXYfHk4DqCNqNLwsALn
SskKEXA/RtyZq+pkfY9bwt4DyowxlDyTN0LLIx+d4GdbsPUdooXf3aOsHzH0qE62a2WaQVKmB8oE
y+MuLy+fOzhzpL5DSnzQpEBmXBbP4JXkeUogslBf6Ce+0/LNronTYGFcF878WMdgBKVIU+fZd3EP
1hXhBeSchttjhlSHN6is9uT+h15FDgPRzfsPUc+FvljObcv8hdO3qFWboYfI8IgpBHYHQC4CnEE2
ay6k5905VgkFXiY2h9TtBQ+QDqEcKe96QJJ/ObV4++nZphXwzI552pk4o9+XiH1L8JizLBpKxC9Q
a++4/GhSfQmfg10DEmhGGpNr1tGWDvIeKm94ORnhzelPXwtCVF4y4xjkQaLhEd1shr4Nz9qOLX5I
r8vZB4hQcKOKJJrfa9Qmp8Yqfv6gVw0ikJZI0z6z+OHCzFIDw4Uk4uAoQ08vAC0fzlxpYMuTmxI5
eqA/TOQECYqSqlm1b7UJZiofZZ2oAsqhFILiIfe6i3AqK0hzoVvb2AoX3ZMgGkbiQqTc+RZETc3c
VmpPPLNnKLVNu1R317weJulCucvMuGkuWuV0dfb9pEmqx0E5yQnS+tLIqC5qE4ARo5AeI25IHuao
bLjaBkvjB5BG8LWCpiZtV92VuVgO/UEKdLSGCaWo6I1eTeNPi/Dn/YHZAFp4LKNE5rtQLSaSR1D5
ioCoQa5rxaU5ain9jS089R0mULCr+l/U+0UtQFSrkvTpxgI1wFZt4Ceq5Coakl2Zwy6jL/J1CpMb
SAG3cqe/3exoCO2KJ47NWaOSneUQ93KoZDy5RiDU4zY97Qq/DFpTQM+mFocek9dKHz+KhXboZ7Fr
zKVWF67JLYBgR2KU9WIZ0/R+Q6uIvYRvWhIv/cRtFGxIzdl01IH3lqt6r9XYO5FI3Q4W+7EDW/Oe
srxYOTsDDwR6oqU1z6U20UBZX8nZc0+HxXWT5qxgE3zmfkMTHWJ7rMBu5VOb2dW8wE+AGuVQp1MS
QNeJ9MdSbcWmn2XLIQk7kWD+/BfSwxlt2IxKp02qSA/ZPD3C79eRFPFygmERwhi7ZPY9IjsLobij
GO0LSut/TQjCx9mVhI9fUQ7UP+o200gjqjVVFtrlVQOIM4KLaJ1e0YzD0NypEtxIwdcJKx6eobAd
Hc3Xp6rxgVQvGtZ++T/ejcBRgko2axWqKb8BJbSMI+BOTlScto/iBknPo6Z9e8WlqgO+aOZm17/O
esmIo3FcLIQeNTqxRFeXR13oIiTYaKFtCUiAXgKSjjk/9+HSH7AeYgXYRZ+ZkHviiE+g+pTkXmUf
Em6wD0Yl++4vyyNXkLmywT8RAcEB39wUCr3lgLN3gNxEj+TcsKuYHYQLlGHPgl30A3PDxsGizN8g
W4kGHB/QEEfXrjRFpJfQ4hrkauV/bmdGma2JOTmE7j+UhJufkAK2l0kXYa3TDPeQhV+H4DhxIJUs
I4NyzKCpaoxkdpHuo0HAMtHfi76lk3Eek8J48LCGG/OiDqtD77EYDFg9foh5hZEcZAZjrdwvJvIN
LLT0H+0fO0v7aLD9lnTkNvqqL+t5AFs8EmjRHKmMkBhpXovI0EQOx4i7yvh3aR9cCpPNR9WR44r8
mx0ffv8twUZkeeG31dsBGiP5IMJddkX6opM3+ywK7mDkXz5EETPdc//+TsbIT8ajRDO853fCLYbt
LO22OdzV95fVgGON3lN9fuqbazKySgHMeiWkqhU5qHx98giVdQPCjN5cEsbzrOGQ0Sx3daVZSBxK
HervGQPuFM50AfBO9dIjydGLsq1bJ68F8lVuaO87ex+YtMZDRR/ghDfKC2kuLqdaL3BfJJIZOOY9
+Bx3vDZNtt+k9XLICmPVJHgNUTzcsBPgiXSQmaqrzBFJ2U8vShYADaSzOBMVYgTQOUqqPY9TzM+a
EKym8pxpIFwfpzOL9S3OCMmXSRTt6H1ty8V5oRjUqYlFWtp9vzUS1YlYzNYMhEfioPjca3D5cU+Q
4xRE723zUtovsD8xiZPWiQXr8MarTWlx9hE9jfo8kKyWY4d/O9UKH2q3+SQ2cA5x5/0iSWOIU4kC
HunTHjvn0G+A/DMhQ4uVBrVbCKRpQC3sK/VsY5lJFm8hksasKY5yR2KRYx0pBCqRXvSqKp6Siux9
wLRWaZuTY2z+nWwUgn+zQ7D0T/3jH48NWIxfDt9i2/XvmrJCIgqyUUoorwCkkFIL2p1t6ZfYzSGD
a1QIkc2ynHsdhlwFPgPe/zh5lFi00YKXmGrqxMH1qDt/tdc3HKDNkqPlKY6wPx33xvtJwioFzXAj
M1oI9OfxQTS+t7KVSaX56R42cE54WMKN9C8Go6/xgiaaGrcAoXV8ANY/whlUH5Hduc8lqbX4nbHw
9UF9Rv2+u7EjpwcfMdbRJrI7UORnaKZWbLqEoKWuZ4GiLgX5upCUX8UrWtRN9fD7OHgIuMOlvlEb
Q+ib4RO8SVJPXNzRgXFNLboC0xVK0UCRq6BajI9zDlJiuwp0Bi1paUtpW9vdY2edrMQM3qBmKBQn
NzZnuGp/pe4FNzjjVMK0Fi9SvBzzz02QrvYkW4FOiKPjgbhBbvDSjnBVulXc1M71syA/16bC8mSn
D0LK7gnlgPxwFETb0acZes9QIEfWafASREKDPYPwYej8Yu29WbuI2S0o3PnE9IgjY4lpAs0SWI/t
wI9ot6kw7qfibpGWia4aNZ4vJml6qXHyoK039YoCzxP4pUfkan1W6cWrxbDLfHRQFlImZLrYXMJE
4WmgWYgAqmkKFmQUI6KoyM2iB6oUkQ7l3IYLRJ9bIDdOVqIWc/1BNApwXyzaDyKvp55akBHB6HvJ
xtjBZgwudWuFahyK7e/LqPqCJhPb3+Kz/DE0UvjwGlb1UM/r67s2Mbk1FjqVYTb9ERsMQptl6PKY
Zw2DzddckY3NA6r9cDKiDNRQlV6YMpBE8Am0HJvht3CUzUqawswXFPFAPu32/wfFcthd8ZX++48W
4dazTZVl/k8dBViQ6bfuW9j4xOE/VdpxYMF9K0x7/Za43h/iPKgwG7QVVULy9gyTYAerUDxMdkob
G+/vatgo2SBEhJPILAf52cZ/Rl9txGHRFdolpkv6YvK/spl8YqPaaFbdlHj4Ty2141rr3a/jtc67
z16i21PP4CbtvdteMyaQp59ac2XaEAC/DA0rdDHbSkqpmodqPrS+HkrqB8y3Qrwj6EebyhMAZQ9/
ULjStF0GWXdzRpf8GK3m4oIb6dkSPPYouXk5Q99ZUi6r2z+MkG/mhhwgUTY7TS9zBXhDhQ2WJehL
JWYw7N/zKE9KtMvcaxBnyGsKuprTWu2EbSc7fRrKTzTYhLasMLCkF3zb/+VkD+hEkzBxHNmUtaO0
xLNRHcr1cPqhVrYvaTPExKkGScKJn6IZ8QMyn/kAFRaZ0ue1FIxzrkbofLhNdyKPZlahrLszJuTu
kud/1iQmlHJMIEDhcmyKx91G6USpw5isQVaIzcuDSFM3De26roXw3xcC+XUIbFfL1ndj8UdG419G
EKzcrYHsWIT3dKDAUaqwPapZlk8+9A8QzWbLZK7e4mmOCMXwOM7veQItsGjQpbUcQy8/PcT9a3Vv
czj6MitlMBsCeVsuPETy47Ad4O4YiolKFmL3ylL5zz2jy+IQ6GuhqHc+3DsLSXUCrOtXMgNk6PKt
iYf/tiLXTBDlM1UM4u04x56JVRIoLlPI6QKk+DJLuisttOvyaOBYn6/35KrlnMoj7uukY2LqPfkC
sooed2YcUBieBmHCPwKE9sPDtALGyfak5X1L95/cqkXgr84n1+SakZn1x6xh2i2F8n0WzMZXO24W
9wmf9i7UyrCNenBURP7/mlNE1IDoIt9/pgm/78rqRD2JdWWawtmczAA6n2HAoKKb/RgAnXwGsomn
KG5JGLb4NUBGbnVc9inxAx8FaUewSI/3HRa8uB5u8IEpcbwzm90xzNfWYoSV2MYb2keHaWe8Y3HW
T9K/kQhVCe7skjNqdLvB0sEjNr9ENlFj5BX4YUjRHaGOKZipj/xjcKYvUOikKrxgIb7FUuupCm25
LMtctulU+6cQyklcujNSRBtrCJAmODxAv30J/nwXklE4aF9DSjZUYOE9Nvvk99BY43D/ScWmpz1q
WaElRk8lo1vdRGAj5UHb7BTvARU3hItov3VA7LemjC/OsvNX9EqVZqPQRz4OblD9PF46ZW3sT8zp
DR42rgen7wi0cRD1SUONSs4mBGd/86eZNnusu5ZFmkcd4Ok/CxLEVl1G2jK0Cn0arocmEfBmRpHa
d1axCV9Osh82JIn36+iXKc9Yl06JEt0zUBKS2yom3dhULaAvrRALnXdwGNlVA0Db9rPFSymi3gCj
XQUOltvLFdkcuH1NXHuVY5XqNEqD+4NoJhg5vxPrOOA9VgZ824Cer5sFHDCmdqEMSr7tbDwuN5IG
vdZCNFanifLDUs2wuUlbekgIBFjN5AYSqqdt/vACXTherrRzKK/nC+YWW0NrCGkbt7tv3s5xX4FW
PqkMrZ7KEOWWWMIGULDeGoMm0icd2fXTacXcdd3PlhSZcOIQdCs06wkc2+U8IaZv11vPanPecaNT
He6Hk5ShROWojM8te6acCofq+W6tmgXK0UoRqsZ6yfz/AREdJj0K5uJwVPlXQfFJWIdlmj98aXwu
QW8hpsJUxG0fgl80PQ6NsoIz5LnPcUH7zNU5ecJKGsAt9066p/ey0upW2Yx67xdGfAZObR7WUvg5
fkptUF7Nx8DyMMqEI9Q+MS6xOpLxN+AT/OlKE6GLVWRIxQZ+l5KTzEWCKKPPAizLl26ypHGXR9Q0
AnHJn5NfGBiSVEMWiFgkY+upnXLfbfdJtLuyvZXJiYEtpGbV8Brj5CBFgE6utAv7FuTxkf5HZY8m
blm/RV4HhrLTXHJ2r8mRDgIyKYb8msGLWRVsSnwEP8LVjykwPtlGzE1aWtWOQgALiljHYh5Y0uJA
8uGnIVa8brmLd76Ks4xvTpe0lboNsnpXRdKjpUCsOVVARAQZ2LbKSRnn2OqUd7KBGUrbBKASfXvg
5f2YPv5EqovCIUVKN5W3QZ6uUSUT9dz5UwUCF/xyoI1U0sAbuOKKjSaYJ1YETpxd9pTV9DUL/91t
a4MbmeI6NKnSwU5/uSAON91aCrZh3cfItK6mvpiVqBqSbVfN+Gnct3PRVKu0EM6y1cjk88xf6XPt
DEjyb7O9EXgPqK8xxOkyvV/1gbzJoIk9r1HxIXvkAMWIwSlW2o/rxRK3CuYe++FX3q/pOlKigabL
aFM/SW8PeCN6X96LYNHAyYc13hwmLyk5DWJNGM1183tK+sLhEmdbsM+dDL/So2APaVEo1uGbjKK4
XkA6PZbTvUxDw7zI33K/XXOUNmF9o8zO8OJFFAlvNQRPmZv6RmttP+TU/aVV1ayXNRynlyJLNXmv
SKK7zf+XMCOig0V8TpTBAJ/krU9espodz2Zemg15Vty8eJtpoWrvZwhmS2ciRKLl89F2qvx7Kx2i
/BYB6yfxwoZ+zjBGgRrkpyqkYiniHXDMRPkM/AShQK6/rNR3Wg0573lN8bBzCOdkqvkkwNGwD29A
xk3uyRYLEO11Y4RoRIVRaITYjpS/FZ4Ki5kKe3o+msIHZrYJ6HEWgo1Kzg5HOiz7NXhBhrXptubD
S2f9abHO3bM11txhHKbsRPSN/WBpivcPfKzPo2JweFtunFxvvL2WvebSOcW46e2j0InZEt4jKJh5
m54k3u8D7IsYUWb+DUB1p0J2mqnIInYjuQIFYyBGpJTqF91d6YM/sq1Yjokimg2yscIt3REK/Bcw
cOxwFwCLGubp760yP6s3KvDMivODIyfAR1h8g6Z31KdLFBy161cve7JI3+fsdsjm7vKYcufLLTY5
mYHknAkK4cce7Lvl3PZn+yNQhj9MTGMW7yeJJu4PEzdRIHpVYg6eLROYpS7NdFgvnaLNnnwvQ2DV
7AUi67Vw2Hkj3D5GsDfS37mieUfOCTqg1+tqSuJAxoxz0Mf973FPoIFO5hbGEtfaSz7u5droDRFR
dkBzmSaNdXMdGmG5aGGFaP0CzoFkEbbJIRfw15VL776dRYC77nIGkUbb0g0ncOlb4XJIIaSQzBCF
QVNmsd0wVKQ8TbJ/O5M1Lctn4kdYZ9osIjcSIC8Fzcvp+DQWXDTU2CmBvoa37dljVlz28WpuMqx9
+JQtJEVJzxzrhK3Qp5gpzJ2VyYsyX+fs8zGT0HRQ7pTXCrEiJI+iqreQ9CO/bWtBNDCLU8YMvnmM
ETFVumj+mnjlMZORGj/JXVTOhBQNkfgcIKLG25GpQHo1g4im4f9v+jvJZr73uqgvW3mOZauevg3W
b6RxivVNufoJReOyGGCOInfPBJ1rUBaBZ60BVvvaWg5pCtzIQhhUbPX70ViD3zPh1mqtwZ1yQqN/
b63qSXF/n5Nw3r7tSjo/cmpMa7f9qvT1rg4d5BGGwI46q8G4WjyKDCYnCpU5+Oaxs2JEX4oe6UM2
xdsJy8ZN1SeTZS+WcUrDEHNqhHfkGmxhtw2WqCIYmU3KC1iAFhMdXRVTeQR4mhbIKp1nsrLLYgTO
s3l8MjtKou8MyyHap4jkMX3z2l8p7QRv5yq2QoKV8tovsCY3uvgRX/0oGE+sCfYCBNVurNq2BNcL
hS9qGtO3ouJhK7gN498r5j/lFH84mbnPjNYnQlKTEAnJxbgjOpgPHKSKBbjk87SqSmrx3+C7eejc
0jK9S4LwALKTnougNVs6g0v+EdUwKbM1wNZDZPitIxvtyfYhHtzkTOYhSj7Eo90g32Wfxq76aDuK
ZoRoTtoVHSC9GnSW2M4zSOiS9si9tzNIfJJyaTwUnwyJfqsDgtX3SmUwIG9t2V5n1nPMhBKvriZy
xCsaCWp7byk8O5cjTxCYGWQoHF2mrfl9P5LU2BZw5dAuMM1wKaYtv4QIMuux9yuz0EwF/z+MOQy6
/7A2yC1vLjJJqxvpr9fw9JZ7mEmtxyFhB60GO8D5acWEhPYtCmDh2REdvzThyA+520FrYtc5WITe
c0C01ohlFSJ7FlycXI8ZuGaEK28Eay7f8w9kXN+o6aey/MyVubJwRyhPXqm0YO/Pc3Pz0SaNfzbt
uv+/VWBBaIYJ2Yi1E8OKwmywT5OtFFS0mO0Qme60TfWTZZoSM+rqN0PwALOvirQEBBmsPZb0Ycjz
1ijz9jp+xPDdcm0Q39HDOHYpglEOUwkscC3H585HucckE6rzcDz1Y+QtB9yMDrS8MFLQCGJylG7n
yBD9FspFC5MJXWn46TjkRDBYlz1YCx5ujCNiD9dye5mmshFEsXPB8gdMkbo76EgA/JJJZPUDrnJR
GpBXVKTqH914UOwIFobzm8f+BJG+ifuIc1J6xNKOeRFZ+gyMKnhLHaOEh9ultKx+IAO+7sBAlKqM
SscRLAiY/C5erqtbY6d7Zhxtmj2i1WMqKg91N3b1qqVuxmJqPGcjfU9ox+MYbHVVFVxgt8lPXstI
tT2d/i2zki5mTBhotM4dMPGONNQEkzySA9jJ6bX5qNchHwmFnwdIeo3JKtATo+iK/1IiES85Ah9E
jGCQzTGvWBdcw7oy/ceXiLSzM5HecW/QncaETtbgiJx9bPgCa6Y0HS21GU45T6uUEfYCZf+7xHLA
/WVQMbS0tL0MkEeU6Gjpdp5AFpZA9Sp1KcyMa3KsawDfFUmzdsBEN2W3HG3OMXqO2AwOSqhQbtGx
2jzbXhxclexzvTxE7wEEoBbRfUAwMXEOtpQJFBjXRYQrAjT9iieie4KG9lIvWsj9lV635ivM7Z/F
EVUCyqVrGlAwio0nHwEGGNaA2EXMAE+IAqXgUW8NtgB1GECulK5ypwTfJ5oOXk3k+qIWzFHvG5hg
19VmJxPDBXK8ooC/aF4bxLfxRVm0tBwb0/3AIpKvmWxvE4/Bm5EAeX9sDcLtdc3VBcbyqaDDAXVC
YX7jP8fP6Q4twdzbsIPIO4tWk40dj5w8rrbnXvTxeB1qV5EqNL9UglYhLD2y0phzFBJusV7JZKj7
bLwJLYnn+QV8kJd5JdZB+GosDqy5IA6eIrZL+KdV1GMQ9r9hkhbj8xtlRduX3MRa8vO3E8LfPZVZ
uO1adQrKXfc96hHlVekqhEDkLDr84ckDpmXf08hjFXVIfuIeEe5EVisRPqihAXtjLkODfIQNqrX3
DFel+aWoncykK6zYfLYa6jJbgQgDCuitTFq9h/sUolpj0W9VuPPN5Ppv5u4I51V72LgPBGZQjK83
qX5l5/7q/15fcfOVBb7I643xyzdntc47l0VMNgPJwqvRtL3oj1+Y2sec8iSb0NGBrjM5ankHoBEQ
mTBIvlbelP6kqNsqH5CxnaYRAtrE0qKz/OoUs7B7ugINzzwfYxszrYvtJTMP6iDpvZ+YHEzqs3Bx
/wmZJPUXz5rEK32imBYLU3G7iIFr7cQUUPfTGHLZz4rSRp8cEbFpUNuHNEq3nZtfmxe0iTsZZUPu
rcfLgfXcjvtDRBO6M9VezddXCZnCDOyqLrGIY/nmEHCWK0U1xV/8YbNDeYUqoSwDDmKqSkfCN4oL
wPouNSRm3LxTHoflcsTdy9e4sT38cyfyGc7AtZ++/hR3jUwDe3ovuMcVQClCvBkGAKN6YVvP5AJJ
FnHc6vyx15IKQYcUhNlWr/Qc2hF8zdanrAe5x82KIQvx1TocuKfkPTr8nxpioNSoUUV40KPWSFw9
gpN/99tVSWu/7D/ZU51XYU1wHRuz+hRBf0uNeYgT22VigBeJ6Vx9BhC7e6TdIb0ONjIlSkOSKngt
zt0Na3FLZgBRKZ7Wnzfi39yGVDbtJpz5hgjlGxO4nnnphxpl22ambWmh9tAHo1SoJyXmXMcw5z0x
zOsktFJA7DH65leYRF/LX6kOLKuMPJbkjRimFQtt64Odes3drnAYFcXeQrEAT62sCNDa630MXFYa
5GnHK0VHgMjNyp/JuPpZ/EQOQZiAM5/ce8maJdPw0ODqvPX6JWyXJm878LkOPb5QXzZW8+b1L0+m
nHPHBn4aG5YC2+QNn9o66ErOnpIHk7KM/4VsU3bco1OQggowBqZJ63Xm7oqv+pbtJSaAHgh7lugh
lTREjBasIKbmfV7+34PbolRrJmwuebHWWxfNe6miT2gsTyXSlMJ7aSpn06yGh15cF+EZOm0Nh4Da
mtOQL7P7pXPyzeto0J516u+DqFjBUPnqRzlf78VfCHZieiiSkrb8ir3SETNGnB5L1DLGa8sqfGtq
au9887IL3nXr0tbyTZgBCB9tlc4tPW/nVVkzV3FJbFvkZFogeBB9pVSlpygkjAvZZFYWItO/LcLm
bpeOzLE4vxtD6ynrmMPxLWFsg9dzrA3vgWR9mHurbEcxTxbHJPZRJw8AkNUMlOwZ5I6of3Qghvvm
H849BJ6KnLCqQU6xJKq1Dm4jqHNwUejILMwajcjpLl0eYtpmT3XS6CVatem9MvWGjwI+al/GAjjP
8SlklFpVPJ+9SOFN2RdvLyadd5hkROLhkyyc6C+t9BCWFca0GmA8l5QyZJaBev7bdpCncWPsHHkK
zWeyJNFmkiaETejRnJJj8bZGKzcFqtNE++g3PqR3ZdlQHjbPFe/21MAj/FWt4GsdWp3UNfTlHQre
PpANR3fqA8FPC/e1RW8tB4uglzMFpKtVcELy/XfHlm14fANBllMudxGkAoiN1IBQSVEVnD4yl5jB
Fv/DWFcCFp0LpSjcyUi85uWpxDXDK85mvMkprfaxx1ZXJrdtw9FomPn6wZVBM5pf3Q7xZ5HSjrqu
+IqNwwrJwsPdoQ+hLa5gnITb9VV5k6Gp5722coIsJi84h3zVJjO6ur4TwhO8j5r4u3k+mhmOfoYq
RbS4/bppITfus4quMdZWZfi/c6GXZbyaDRJapertMfTFxm6h8OwcXM8d6/raBVqMfleWqq+yHB4j
iLZScuFDGb3B8pJhAiYxSdLn18IYmMDmoMb3Vb5demwEGaG7gwBkKnzrP0YXfAj0AE3OtKMM+4OU
X8C5cRqQaD4F0oUt1j2J7YHVJtO4Q/DpJDfq9qSGMoUOVF0Witgun1Nv2FayH/l1ao0Q+VrhCaKZ
KeSwGHcIBiaKoAURxJPlsTmsdU0aE4kIft9rpbxgT0wYqAqG22rh0G9ajLArVfJ7AaW3J+YkZtLF
fGppQGEvnb4uUqVrox7TkCy95ctArU/Y3ddaOuvItRYGIOcsAcQDqtYv5tlrcWh3l19AoP0/Qvwt
8TUShSFURkgoGyG3pp+4ka+4nALiH0gLC9BCnYpd0OuHgFosGzjMDxe2El9JRErpwP5+Th+OdB3d
nfm46S3OWyBgT0KP0o7WJvZ954h1PWTRYm1CDqYCa4byV0f8F24cE3WDTmp111ONI8KCx34vbq4C
mSQk0IqvIRYrpOzosfkgWc/TEAwpbJC3GhKnXo89y9SxaxQQ/R+XTgFe2PwlIhdP6Ah0iRhMbuVk
1PY1IZlviFodKqT4cHhfNeuAfGY03P0IDi5+g5geLlXQooLPZTYQxatQJc+Xj0g7UJoiN5wOR38C
/8KVIQyOl3uosFp+nzvEzfl1SXVmJjA4q6k8xP3GG8trdMFqpvWI5/GnQTMOerX2zumyfG/Wclee
e2TU34QtDbatT62PmmlPBIaIxPdabziFtOpWxJbtC7z0Lb2GHJcZ/Uszfe23aCvjqCzqEmEgtB24
mL+OQIFZAOavUzx/Q3yrOo/+l/CxQw6MTu/SUEU5fbjDHWM4c9dnvqXTUkUpBHg+M/WcITGnJ02S
mGdKzNuKz6hwCIl9wOBbiP16Dz42GtYJc6zpYL4e9ZI8tVH/kZFVYBwjJ8p3tZhpJyb6U+9lHoZL
uXiHAHHYEBaeiz34aGVKn5BvFwBWx4s26y88yrA/XsrqmYBMOAORPDBbJrD7324rIhZ+Zs12Oe1Q
SmfMQs3E92HJ8+KyUIM9C59WLymedsOVErJ5wsCFeug1NuCJ7DXl4XHfXF/uJEvyN1QjOjVPN1fY
0yfhf7u/ZkV8r81tFZQYo9TzVRK9H86XatKXL3gp+3S8YmoT3tOugs043T1mBevSrD8zMGJbLWWq
ysOFCSwtH7Rs5V89gIlS+kRAWazUxf6jEfDIX/qHOSA8ooatM/W+azjq5ODvAjOvcp/jLZnv8efv
Hjhjzbf2NFJSDyD8e4r0/ybbIub1cC/qFBer5yVZWoJhyTqHwQMAoR2dmkJZz5p2r/8Km8P61j+b
Zz+QrZkaOm/ldaiyzTCsA6PLpl/m/fHJfSUPLGpLCN3FpOsf5RaJfbRzv/9cfQGh6gVTIlddBCBx
u+QzLG1DvGb+C8lLsnfj4gEsNwE6dc8kM7eeyao0qzGJ8nt8AucJJNJn20S150PwbMbfvaJp/b8m
74RcuMr72QexxyNQcrcaIQhywR129LNs4IoVLmeOpV3j6pUqUFiZnITSyrVtPO8YMWjiOszY78V3
LVPQ+WPXtC7CQ6Cbp+7Sf+N87EmRpOZ0WTJvSSya6R5zrAhmlQ2YbbE1qPPOkvhKsVjjTx0s1wr8
RelPTV7jyv1178PT3XUgYd9L1W7GITXTsOm5noQarhYAxREHgDG+LmAAYp2pWaELHvY4v2woS9Lh
O2I+PnBHD3PPK3JpTlTJD91i+xEYbWvdwomFTLj2/J/Ay83vt7aDjzJTzddSK10uLzLCf8MQdp38
UpqQWNR3wFB1TFQ1GAPCcgoWJFTtXT8weQ/HuXxirzi06Mg9OlF/DPV7hFoPfJJ7XK/eSaVQ4l4c
RGd6/ezM16FSKS6pl+wG1NpCIzmKlKIhotvdh9KSQBnS9GzHWVeGfVykDG+aOoNaAueDTo3kwEVj
fDDCHC5qpaesvorVclw9P0hMTNL6cywYTgUNucTwzJXRdCs1dq+TG8vk/ydOe7m9i9CxH48UcrR1
xYsnMzr4DnTruGogabgv00YIsTX7o2aka6F9FwxcTheG0yTHJ2a68Oiq2Qx05cRNA2huCrU0rJJn
UMT5N9xmJgJoWHUBRad7RcFdHGNQzEQe+ckyKz8SwtF9FkeRng8Nk0eo4lRxmACoEtOVBr1IDyMY
fGu+YropOpZ2xNLeGF3BObAG/zTxksxdIgee/fuzRhRI4RzbqhZgNRz8swJiUjuhH7bN5hQ08GFZ
Ag9XMF5c97QDwit59ZCWSGrU2M44ryH+llQU+H+ummXi6cgDMO7h4qPhgXCGTFFKlnf1LxuVS6l/
RbhtY6JJRYt15Mf3kwrF2kLDp+oAbQPkIUJtozx3vhE6UPOjQirZuDiz2Iqfcuhq4WweJ/DzE7ef
5wbIAJKkjQ8AaWcY6bIf8xNHEzvAOUhjwC8gHLjwhAfKUmu8auOHH7pn9vecCYypO5muG+NzupO4
FHkll89qfGo45Y88bmHm8XjXplZy3cZQFYRhYcB1SMWjb6XTx180fZEGVTFAkq/WdipQN50tjzUU
YkyLs1418QT/gUp/sGgevd+kfnwTVcUgGKrMGrrvBjxfN7DP/h9tEHAnW+2msb9oOotuc//1sNwz
wQyCCAgtPv8FkMQ0JXtz4jlh5Iic6W/l41LOwdWP+ifKvwDhvfWkeyCxGsEeBQBCBKAxCGYjkR8h
WB2z2/gFyYJiUSHllU2QHGbR4+XklQEa5Nm+taqiT7+v4/GV5lsxI8HxNJFNqRvLxygGDjsNlfSP
9p+n3yRPQPFD8alL6DfRJnSrgkFkCZcu14YoKnBV9RLqPz4kUQbDTJvfIi6BggQXW3HBVjGCtrIA
Efy1MzvSGLYSnzbyqibB5rAhWdV9Nox0gFBJM7cXGtJCAlpsN+Yf4oI4RMnOZWAi5CBFUqMfGyDr
t/djpYkOcqHpAkGH0d+PDQoh6KAbfDPHp6SBudhAik/AK2efV6BGfclmjAm8mMsuTnBqjd7DY+DO
GqmsRiDkH7RJI7j2/ntngEMqh0nXrT29Yz4pW4LBgBmvbih0dnGTNiET+GkB3zH3wOZF9UAvn2nL
8ijdd1tGUPBVYwmI0zIcxYGfBPSpdp4Ym/sXeGHvZaw3qeWg/NKo2nyMO5V0UBGVTJ0QrMdnsogY
9vaNZPvxtmGc9u7yQONjvWGAe3wzwbnzYGZ0B6UlQfkf8sFUC5j5UBQJ6zNzY/fNqZQKV20U1ON4
tHrem8cVv+3coMRYDZ+mLqtBlW5hxCAIMhl/9JRn8umBB9lWQyEMFSRSfqSY5rx2/wUWGnMAdntD
WDywsUQcOmb+P03XakKB76UzsjMDhcuEEo+82obEpEIHt0LVMXPfrpZE5eMELwPu180pg46qrf63
8gWAmYrsT6W+ZWKxNKu93vDmqT/GWkY+iQ9LpZpMTDP7O0hL60Qo11bMajJKwMbWTlKe4Oc1GcIY
fahWdThZ+OFdLt+EFGwE5II61U+vuC/i4DlnJmTAsvKT/KuPHUGca4iLr3Z5HlZVK7PtY5F6CisO
uMDv1mu8eT14fVi5SyeOZpsux0gVBYwfx8Lvm3VAjIeXvAhGn1HIF0Mz/gBbSMzo/JEwM9ftVpbJ
iWQGBa4wUQc7KH1CdB37NsprZdM9SrcTXZX8Ko8ojLsAUkB99rNpDTxrSeVHwD3n1Vj9/jW1VkbJ
LkCB0wtDmnBRl1QszHUR5fgtzCFl3oV4BQ4d6zgTDKAcCevC4M6JoxcXR+mHdszclBy53ZVloWaa
knQfAXpQxAluLfpJkv2PEFsivIF+3w53SBFYHW2v9D35crr7m+9kEDWjWzNlgh3JCawG0GhFHu3l
jEjF1DTZkZmHON8hhKA6b8Vx4zMbnBnKwEtpke7YUdmtWgQOXMH3n51kmKEgzAawbE7+yozxSGdw
hf2Z406aDUXDPZDe+NfkDSXLabmenujkQQYHinIRjCkMFtpRmTggMzIgrIbnPrmuRMV5DI8IaBew
M2WklF+3tWSauwst+gkhde2isI65NpAMdHgGvXNBT156KwzjV8AOUmp8QSbrCHMporZgE6xeVqmb
LeCWsLaB3w+luLXc0EE3j23SQuElxEqnKYgjMOfIRw2RzqYqQC77VBQWbbE93lY4GMhtOvLBB/Js
5Nz+VZfJ+DTyPTUDcbfTpSIzjU2HbZMYeuFRw3Um7UOQCPvGwxl+G0e+zx3IjVsJ4C5Qtw/8V/7t
LCu3UvRPgr9acznE6rL3mXYcCxLagTHUnx9MionMW4hQ344DLNaSiyp0VuBICb8sz36jHp7eGYYj
cIVbcXQFFgB3csOLWK+keijvQswlJ4FU5B2YuunnXb7jZpBHUa53G3xbM6zeDcLix3bXaS1ABS8w
u9y+0pj3leuSvuaF63Tu3g5mxrm4rZNlfOud49hiu+DJxfKq+U6a7mBZr5XkSC2OEQb63PEbVqos
2TQ+KvkzMMSvc/70dM8u0QCg532yGhnkQEw0x9hoLmyESkPpa6a3kQ1qamROmtz9WbtBCfYK2Uk1
hoKt5wpUkK0WgADkJku7Eqa8cbUrq35DrgOIwsqAUzo1dOK/xAogoe7XPA3tNLoMXMCkLsRjuD/v
sBX5ImQPCH/Pu+DhgOtiBe1pUfe5DwzDxpqF6OCyNdnWHGrkX+MtKGYyWiVs1qcS3rwrruyT4ES8
AGdiz6yQQnMDFEuc9fsNK4+itOGQ/ZS+Clm6i/EpWgPEQa3eYO/sovynVTKQ2oMfm2VVS8ILTe/s
Hqgq2cNBExyW6Kc0TJQkRi3Q/77usBBINfqc7yvnQyzW9sGjslcTUHfIo0RKwOIMKwiePAHr5O+z
I9fV89LUUhkS9Qd2+6V4LcDWMenarVi3qeikGf/nt/HK8QgJCUNaVozIhoVlCLLbfke9GHL/agQA
zNUPrLvIapBl1tQERMyZ/0nG5/AENP75VeJp7fQu1WI4RIChzGRicq2pIxv/tH5rcHe2yBCZMjv3
e30Wnf0P7QKI/3fCRRiz+h/94ksSjQNHhHTEfLgeNJfcpMI//8YOxGgPhj6nHihPaNS0qTLXC/Wk
GOtTnFLgKWLbnisRfxDGzyimPaTQbBCHvLIzyS0R5KQimbkw89B7qGyPDET+bJvpeuefRSnSDAqQ
hfnBLOVNrimlQCK5O5peSW+JUFdlbVnUCi1O8sD8IkaaMnnMJ5CP8fEMISuoRacTy2YKikAyFBT2
uZXcUiuQw9MnGzksmkH0urFn8+USp2YxAv2bXCoW+fUHbZEHurbPyQpYIfM3MzoopIM4J0G4yJq6
MRnn5tZf7YFSJp/PyjzOlJ85RWKp7vrw8gNa1lG4O85kY6FiOaQpK+siAx8gp1CQ+oXcNS8ceIeU
ZhfGtdUwB0CIZ/AkkMHY0U0sr2fgBZpeSK0/Wr9iJvFSPRPpZIgvj9wSyIgD1RYloVVOtTA/b5w+
0hvqwxU00jqxR22c0GSk2eUALSo8slZu0PTzqI2eFj9oE9cXCWw7/tiR3k6RuyBjHD3atLT97hIb
GZg00sufYfHrMrIJlUg8UfaV87jpJzF9hOVkRI6ahmSbAT4wIpaLo4EWdkjjRGLIq4dDiB/f+o9w
LyauTYRQqEmviW1LMG9ka+2MeDQT+hYwhECfXIO8VZL4548M4QIoVCoARSK4EcCU/2yBGNQWIuEM
q+k1o+0xjYxCgpEe496kJgLIrMJHPXSOiBwGsUA6rhc44XS8oZT4Fzg2yF76o/CASPxSD5BQtVh3
zNlhjPhOezRXMK+yN/pw02Z7i0otXM5U8ix1e19yY1v5Pl5OCdJnm7Zmkhzb+3+4e7QJoYnZf0BT
082PeiP+4b/Ds4U0SsTn9tGNolCDTwhbu5BBNVC2eRwt0DOwIAQgk6xsiyLD0YchJ7SqAHEoxqdI
JO5fju4DnkFOXY0teF4YL7FQiygC7+U5SJHWu5osudPzY4mli6MGcGSwuK3le1Wij76bRx0aUdu1
pSkcZUI8khif9gYZUq/3ivh2iWlXZDPB/L/ODGzv2X9dVk/3rUbefmdV3L22zAIrML/HyCMHszVS
m3Gn/lmrBik4FGiw+Jv03B9OmlE6jAsq7rNoXnvJF5fs2SN4Xd7kUCmnbhS2pVf52zmVRaDEohN8
KnyIPw1Tgvejiq8W29yRDgfbXWiIE3Djc7UVdi78U5WNxxB7dawAggf8O0O1Ns1BhNWrEkd+cfdj
763UIQ/6exjce5EN1CsbTO9NnOl4g0iTwcZFSy7AarZC7qWBTf6bRpTtBcYbIcdtbUo3BbfnGITO
A3iY8NShdQolfaZ7VPTyVLYYtvsbUJKMNSwVsp5IvIoYaaEXrtjFVmEta2THrqpMQQdPuDoZoXYO
Z3Ny5WXxd0PX4DPM0Z3+ZG+z7FBom3iWQX9iwrbIrC0d2O3HuNy2cOALTYWlbdcUCEpVjQUg0b5Q
SvmmfdpcbQHRpz4o0Gwe0hIoBDiOXbaAMLo0W02r9cl8h4STcD7Y3zb5o9wwzPCc1ck5akNzrNwg
reKn3EiagyLQw9/D8eNOoRh9aAcvs4YjuGaA/TOXTCgWumXJ977Vz51vqQXkR61Wlrqgwb12IkG/
timGWHfbpyf5J2NufJZ988daBZfFZx5O47VcLk5znlTJv6x5QLRHUtzhchRyMJ8J3ILxSSpesNa9
9b14PP/QnOIqiIS0s53iC+1Hm0UmUBdaE+Jz42xmLm+tjFthcDgzDAYmHk/pT58H+fFG92PAdc1S
jH7eUPiTJOsvOBugASY8a1oTQe48TPYCOvDqn+K2mIEbYfHBw1ywdYBuzY+cJXZnAckM7N7NEtYw
kW6pA+XGeD3ohn/KytqydVBD01qV8F5DJpszNNZxC2AYxc5CO4c2bF1UbGL6yAWmED2kXrxH32de
rvdqx72ipMMuD2uFnf+2jGuRh5GdcD7wnpT0FrVe7jiy5E2PrX819OJTnC8smMTMRoMRg2G7fYTn
AUsiKeckDcL7hT8+jHWJC7aFcZmMHiokA/T0MTAFwFD4yv/9b+zn+n4boZN8eIO+c6/cEiuzqMEP
Nqc1Ku9nPn+KMPsfSKHNfqSRwi4FQB2Qdibtf9N9+asvAknzKGDW45WB3k+hsAtZTsNicN4xWlKV
sRruDAu+6OpIFVJ63G9Usk6k7FyTTrHjxaykawHb7JBpiXDbzr0zP9q303VBxb9MpBUZ5YWpi+Ab
dPs76Tq/TqglRuxXeHqrjF5Rs5yjJUTaNrRpCCEoruI7h911vkt/OsvNUkmGR6m3dcGxQyyvxYzD
XbtiHRnC+YfdJIHROp/+AVwbglYTa06dgUojZVI/lPo307ets0qRPJTII73OedKMSlSeVdkZ8DB0
3TWASZIofjl0wKRP/SJqjskUvdDWzV+zvAzOMYAx6sETGKR3m/PmOPfVnJhImko+fk9HyHYVlVWH
7N/fp1CLTekrIoAHXFnPgpjV56L0VODxBSTYyllF/qgqNOBi0U7zDqfC7Z/fzkBsqCHv/VXByBur
2G16tBYNvicPi5Zcz+g352GsGkZc1ikXyq2QkN9fVclrbTTgdj94r89/4QqMqGOnfDSYHMuRUwOk
MUNjrW6m1z7BXloT5iZgjOmFeOJYjRmC01T+qYygmqq9PWKB+jx/fm85JdhsUAbtgQcK5gHwRO9u
cAR0f11FsOthI9kxXk87YjyYN/lQ3YdxGhPzhwe1r0zZQNueqNq6l1yeM795tAHIJiEdHQl5eM2i
Jv2SoF0qOqQu8CYe/v3xHdcSAiCJL9mJ1Wk3V6jfNedYeYMBY0NGeAfCQ/udxC5n1O5yZujQMpn/
+T4gfOyEYOeiUvsie9IxI8gpfd99H/WDfg+l/HEP6NLTz9YoLXINR4WkHpZoD/MtFoplkD/17DwJ
XYbwUvAARHDKteWH5prZCGjL4P/X0ituUuN7Hef+17viIoycZ+ogEDVd/D9zKmEX+ICqxDz4RD9e
r0h62YNXeG8lIq+xcIr4LsSfowJqq/COoqQtlii20APJZXcMLHjE0OEKAPgRShoqXE6QR6IdU8vE
b64kY1JwJFq8Fdqm4HEqQ801AlTtyEDlgCWIT+W22ZQjEoJwJPdpKWZSmUXnjXMjOCkLV1q09dK8
Q8+LfTQf+UjgXlsuWpNmria8YqkjQWJZgA2MhHUQTa90ymV7hT6q1RpQ6wK5ADIFQhBx6wWlw2m9
mx3vNsu2G1dMA2BSGvCt4EbxBG2mfkUcVqdY98qMfMY2jOFJ99QufSX5TRExw259Z1WOzWv56zIS
pT3yp4ogTxJc4fnrP++VGsaocjkh9KnaWftKCAPHeEVd14Osow3x49t/oCb18DqiZzZsZfiNwvCm
YBzsACTgIxE4O8+TdOn+H/eGA/5H9r95B1miCl+rbXVM08W64fLVBMzyyMNKMR3fDTwy9S2VexJ7
7XHuVwpUdAKdqN8ArPx4la9iFJKglRgEJhVzdjxsehSvBkEbkmV+mq9Ku8U9xywVFuLOr/7RopPq
32lpxuhaxMRNxvmGXLEof5as9q0U9V7DcUoKmrcjBBaDyGU4+kCfbAGNVuMl+xLb3/BYhzyUrxE2
tqFD3gX3ovGhD91cB4wjTbO9ySdYsXT/E1CP2KMheCexs/mylE1fisvdOvbECGrBK8AzG8inCy6X
TB7d4lqkZ55f4i/aMLLFr5dOn/WY6c5os37DAEE55/QF2ZzSNu03JXWP3mOzXyt5imtUm6AolAnu
RLjA+AQMSSb7VH7HzAl9fB9dWdQAgfCkmvw9qQn3QUBXS7tahV6nVTrM9FhWW2NJQFppvqQcAjFV
vcVmFPfSektRkMPdIBdzvkjpBFNfXp3PdsmK3xE/hMvLvUBsh/6WfitUiLKHxIC0sZPMSNj1v7Oj
hYhYY1+E8HujG7WjcUx0abIWh+4kLB9e39hL4P7BXhcolBsLj3MVqoDMXXxKkWWqaxsZvVuW5HvH
HNFcHx3DcA75BIB0UnGjVwkQ4UFbf41Txy3o0W8di9kAGWaJahHHsBp+FsK7sd7qyDq5OyVOnJdr
mg9vy7PVc594tt2iMIw55unSoQ/hMBvsZm7WpXT1p5YmPTwZ/vqnOflOER4cDfv4TyGtLFLmGMG3
UQ3N409+pUnAOUCQah0XNWZjRtFA4g47OqgvxVFDaBk9D8TMwFLjH+cA3NB/HrYDLF/MV+N8i2Ok
Vi632lbY9rZ0TWMFktUW+BtoruU+5GYUp1i/X5bgDuR9Sda/qWeJ3Bl0VQVPomreV6wVJrnZ5lD0
hRcVq+LXAIj2cESsvfFU5qQ49TNieUTKn8Rt4jVe6wGusW+aGIoIFK8VEPmjiStvd7J+nRQGCPsh
ZtgN8td72QTrxe81yAEogmoSpLafxKNZXJnW4bwLtgcXr9syDjiWW7c37XC+LTSO/aVsanq+Lh8t
lNVH1H2UKAiNPEzbQmK0BnIEPDjPorhU8dO/zdo50EjXYa/4yhGQofzrNccECDJu6EVUtK5k/fXZ
IJ5TsQnnFHnu/1YBIEtzsbVIIb4UqnOxruSarK6ZGYIUKjITs5SmN8/eBwiqOLS0YVPYddi2ww/0
WRNU3YXMTz2uGldH9kbC7NVK/y12pLN1rD1NfGO2gsOP+2gDsoKZeKxQ2DF5IM12OB4UwPSK2LB/
2P5o2/vhpN/VM96g1urWhli9EZ9gb/HauWJYqvZDp9ngFCleuy8UDIQHLK/tgf6P6ig2Y/ON0csk
FxPd2MUl4rOxUjtnlNXaH/ZsKyelrgNBEYlpktHWFEt7cC9YrPrBL93f9xGNMycxFawPMIsd8YXN
vDKy0bSR6e3bkPtb2M2dy/MBnms/ly3wsZd4Dc0XBsGHlLnTYEAHr7uwMta4PNLDPiv6WfgLiXeI
6oMEGnKfArqlC7abPllZY6+eCoHBIEX/LpUmvYuzb3sDqF4rtN4jTybKaMrXduhnDnZ8KEupEUWl
GaPRW/dkVhWOAcZZLFOBkIatWFzk+QZ5+vDJlJE9t900Z0nrQhMN4/j/4cZimKB6Om8nTinN1A+I
KfmGljjGUSmRh1qSkEy5rECongjw3H9/tDCYzWWzWLz+u/NFGp3uMhyskhVGZUTqEQxEwBuD0Pgz
WiyV/OaQzP3WiqX85NQS4iHoovreHcTHTIKVcfYSAWOYaHIWrIR3SUzBOaX6/LiZFcQDMoaDE6yJ
Zb+VTDnL9EbItQecw1fXA3OOTFIWXdNiOjs5ptAy+TSQ+XTsJy7BA4byT6K9+E9VR7lxRmuQ4P14
KqEua9u3szmG/Xb3Cp0HA7I1F1D6RlOjbHTFTkSQZp0iHsqaQn+TugyZ6gGWFTAdo4qrivVKIklb
bGMDHeRvqZEu0Cj5t1Zu/Eo/DicEZ2puypWDFXWNCi5eWrmL1yJ0ZZOIvGM/DRHzuh+5l7qaRPWy
OWU8ygTLjO8qpWwo13jqoPTEzs1rozzOzTepzg+XE0X8kj7RIWKPIBGtq6GAuoCvPr7ghtnzxZs5
YPjmC9ftrxGpqjt8UbOUJbYAXkAUxFbftgoa4Tn8VOdRnZpHTh7ptmqE7kTyEFf5Kt0MifA/toaz
dMdE5rOZ2bwK15lkykcsbky44W9hdFepZvOBVmoCDZV1hex5/ye3c6N2IFrXW2tD5rGFzRT4v/TM
LPcnC2kAycWHCZ50H1xSKj91zRY62FW7qgch7lZST+AK/uc3nJfZuNT6EIysawpkNs9dkWM+1bso
TloLTdJ5e9etUT4sE53+AXSe8qE3/UoRSdKML2U7bqxrL9uTtRwN3dcmnc4MYupjq67YLWmQfs5P
tB2B4ej/JQ1YxYli8OcXXi8XpP99rfj9qrcTgg7vbt5rNIdY+VBdTaxy9c9M2uWzC85TiMTs4sTJ
avU9E6bI3dJYsp0i+v9R9bz9ghJaI38ZZI+mWVTK4oY3Ei0S1Juxkajunjj3AbqjQB2wtrK7rh3q
ASQecAYkt508Tdm6NRGw8Wo7N6BtzEkSXQ9/fmcQdukvIOa1IOKY1MFbMrLTEYQuwuAF60wByTwr
3X/J87jDjuAM5oq0y/sbLBdFxViBlkEmv0T+E3eg4IIRLdEnycngSa6eWcF4UQOIa2ZJqphurgx/
zduO9slsQMy2RZG2UBbCLhy+rkYAd15p8+9Do7GstrryeFb5rpBoLsl4DnkVvYycC4KR/wVHuVOa
0mMrl47ufBORsj6Jtq7vw29Ke8Tcv71CT0RqThWTOeYfOMjuhymiIX7nRMPMu+/QRUVr47p8ie7k
SrcyT47vesks8BhMT2n8c73+GkHodOI7yaRty1aEpbs4w7ChNfu6kNnRUxDRGkGX/fxa1C+sQuOt
ePwEuCUx8yxUMllsKaP4Pa+rp5JgRvcrk0jkxaAnw7ljQVAJLkN4zvaNhR0/bvbYlnkWxK8SxwlB
NrmJWuEPPb+Qmz3DjKC8ObjmMjI8czkWcNSNgqWqoNbv6O9pWe7VyFW7xaXWYSmHnrdFoPg0PpG+
En8JtDv46iHdPgFh5RY7MkFRpdrvwQ4V+uv/b+eEKL6LZLTg0inoitrFxV2icP4ty6DBx7fpy3fy
li5y5i6VWsrnrtKPfNegF4wBwxatjlkqmBOrRxeUsaJsTnFYfYhmO90YZr9ncpMaZkgtCh5PM/ly
KeN57Mgju0ntx2cZ04A186BKdFTHadQcYPZqXcD+/NzUhPKPQ6gygGURm73s489+9wAV0QKhApej
NQATy4dR53ua1kWSl2SD9lvesIDKXSRR9wTfMTyVOBNVFJL1Q8RIBtAlEwdHvkXDBPhmsF5IYEU8
LqgR90IWBg9+hX87dM6iSWto3QE7BW9CqYzBKjUyuVHzvfLCuKtv6BpNrY56Y/jzNrC/tWNTTIxU
42rpc8Uq/GDxxtiVMPdOrCIO4p+9cpbBbDdKUBk6joDzKEbuD55zOf8Dwadr8e+u6HoBlO4FjKH1
CuqcDrJVKtclTZb7SYSlnzY4nJGtzabc+Efu3dckR5LMxor1M5mv1Un5qK69SeFU/+++7Uhz2jEn
5g5SbB71cIGX+oolCph6AH5FW62QyTwQVUsJNWKNlDDe5XarSX7w9nFZTEPnxzHoWT9csxWtu3yf
ynnXEOyfjNVQFHrM1pjA9wI93wDWDs3Fw0/RVMULVrNYhZ2GJwDwHrv9a+IYA37Z7xtVV6zpoYyZ
PsERoRW7BXOIklv9wxDs4V8KfNkJl1SnIC9vLzKvKgjFK9LeFZhktCCnGliBkjAmZgo46ljdIukJ
N2WTg8Pwu2Nyht503fQUQxEYSn4oNim5ZEQmp+Y3HR/7HeijriHAbCYNsSJCgRcZnFppSy0ykrGs
8A6r/rsX73vC4bIPhCIlL3gU+2IEZHnCnpLCMmIhanAc/XoqqXHYhODCj+BW9x0Ucrfdm1+fLFqD
IGPpAEYG2UHN7WbcniB7ASohlc/9UjOZy8wpliD3PqsPC7ghf14UOCeuv5ysBdX1lK/ZN/4Pk+T5
saKWb4M3s3lKIrgZFq+BpEyFKUT8I5DYgo9FpntKjGPb3ioLukuZ4w/K5CcP3EGG0DKada2G7iwf
UQRrIVyhuhOVUELZ+rqRM5TcrIACmOOKX3vuGKkUijG4nc/8J/6WlPB+FDw6ljdmwCsVwCXDycSb
z9CFc7McdWTPYvdexF2Vbk2HE8oId1YSTLJmORZYTYeIQhsZ94sTNtcA+jnat02FskQYV/25ICtK
Ybdw+IBqjp1D2CF8oYex2e/D7QOi+YIfzp6IaxsovBxkrGyk6r6V3s/hUVYO5lEYluwiLHQWtST6
saXtIKZx6XquhLTXI/KkeS16B5PptGuGaMjfxCtAcyeEXxb9fLBaBxT+HD8BX2zcVlkj5nkte2sP
gN8H7IY/Rs05hP4E+T2TFl6QvyyAEUVkeEFinKBgsKIAEzgknPrjrDKzPOnSa6gcKKK1WeqoPoS3
IwftdUFFkvUTYf1juIN+t4GfsjMaUusxIxcupihsg2WqxlKztQo/7v149X2gbvCkF7BmvpRoDMo1
uBVYOuKWuVVHPCT5xmu8ReSqqdiTYlijQ+HgMaQD3omzJ2AV+YIvKOsUcT6DizVVPwUXga9gYRso
TOpt5Xn1fcc9fPDvwCyH1gFdFm96L9ffB7aUh7t59wmeF6uC5qUO6vjPPdri3nmTMzVwIRkPN73s
t6LwH3KZv9BC9j53pXBEJnpsp22NAgI/0oeOE0trj/LWnW1AE/e3PtBttU4U2AltbXipxauN4UCT
vHvlMynI4MyYR6qofWnKYTz42SoBP0P/FCLypoKrY7kWQMd0QHHI/SiNcLyKJ+z2beoE1I3joU4l
xnO4TA7HpQ9XbBI9W8qRJOGzBt9HbjBZo4THuQWkKbCDRGszw9W4DW2V7OnGrE+uuoi2mbuA1z9M
JWXnhpYbTZkkajTeQCLgbNcdLJJ1bVY8D8roM16R+xrQZmxa33rwITDRn9wBYJlr53j8RgW0mjhw
k+Dn7sYid0WFVvAQGJvPDIaC0vM0XnJcsKJuF4VsOYdKRMUweeN3kY5QvHgH0m64QBpsyoLXn4Dr
ms5gY6n8hxQS+SCYP4qOaqExNebFgy/RD0CnnF2aKtVr9T57MVTmraZ6xPSauHBZK4pFpC8bnaWl
7yi/UWTd8TR0h1lc+gS2nIOTJ2kk4pa4AxaUX0co2ONIuXLotfbo/NX5bAJAuKyZ9swUitieAF94
gp4sEoEqqcsfPLlJld+y6LRTCdWxVFhHFkV4pHNi3VLZ5LVgD3MSX+2PBk/jRWm+JI/9dCz1ZOBI
jMFajKbWFMqf65pd1BKICnVo+G+A+vqho1AsBgVOgBwJFMrW8LyOAHr3ptDG1vfZyqVf82V3Fveb
M6qc3OHDzEI41rOWj8VLkD5DzZld4dVJZFKuuRQyCZW63V+ONdruX2rXE/KHy4N4BdZACCVH+zMD
TUwsY7whgZQZr6zp2VAz6Lfcp+wPJB++/4LTZqg/lYoJp33dsjihb8Lv7URyRu9yCehBYsTxvwdG
aKfLWqj18FG5Tm7oasdlphLxSE8vDmcip/0SCrxMMtQvshGgxUt8vnY2ORlbQxgmnuJOoJAl1h5p
vtxs+pWzOPt8vO0A8es0T4tB5gOUIn17lmeSP49KQUToRTutkuMfe275HFp/sNVpyX18FXrZ2/ob
Q5xvbbY5rzRiZXxeqBf/L6eFeShjmTaNZL3uOUieSrllMZSbhvj27TeHXtYIrb3SuGITRYydLPlJ
gmC1ZFjoOmnsfVkDSNSM+mFPx5BAGXi/OVbLuWGamWifkM9RCv5jnb/hr7xdbajYOhvOXyHEz1ma
ao7mWmPSN63qCb2cOvINyVLewja5n1Yuk4hYyB24bGpE6h+J1MbI6VHU6peUZpeqrhi4qnAjWBBd
FJgX79szhq2svVcD+Smw6lFYy1jLXAY8yLpEFGbSfEdgVQlAn5GR5MVkcK+DBTwMJ19PV/pqZhW/
w3Iegvocf8ZknDpiLYx7qlwXJFbypHbjM0IPGnv3pxvEO/RA4GtH28tO81vGTqfLBb+cUAO947rt
F4NOwHVo1p8ksKKIGzdraqaIpWwGVQJ4N5hL2lp8c9UINKSD/4xh7WPjKMxConaSthdr0/Xks4Iq
SvwNJtZl3/oypGeAtZ++CjOL+xZ7iU6ObvQbOXUmjEF5RhHyZeLSSwW85voHesOJ9nEsS/1q7uFg
sTe+QmYnbdDYoCW9Z0Sv5HmdPohnmwGzDPW50h6rxy+7hugXCQEp4UF6VLCFdiq7Wd1upXqMzihH
qrj5mBLnU+2AgwWkmDTdbtgb377BSD0fMw38lNNm1ImGWxZhmPRx+evvZ9v8aYzOf5xTxXFeRlAJ
XmedPICTtjCxft7V+KWITH5ynyOIRQfZzG9xUWs3QoYuQln9kwsq12iBwKEJJ5VPcVdJj2f+BZM7
XcGOWMLXv83RvGZeYYxVqeEB4k1p14XjaNyTbBaXjeR1yGPf82T4DxNPQcdPfgrrner5jkXOTqVm
je51rjOyb6EyvycLqVkvZdNmWfqcCbb+zv/Ghabp+mO4/DLOzK6W1WfV98FvT1KgrP5GbZ423Nor
NgCJ2VHup/CYsesY9+yBQ3DM5NllmJebH4YwWcB8rbYt0rTGXDGPLxtTr+p7yHytExqR2mEe5jVR
U1ukeNYBFD4aWXzOOUHmVqE8OGguTrUUAcSAtWvY8/AvLQioeGgPrfBBNkzLcLYm2ui9c/TU1X0F
+cXXJVoVyRmfZMcXARLRZtwcO6VABFp4XIUJYjt/2l7fR5supVp6MjUBwXX6IyrTL7i6Q0dsMeal
rfR27KOZDDik9WzSuUwpNxD21EHKX1X5Kl/AKc7I8nA7Y5idB8FyQr2/tJ8jl7vn+usfwMzrEsd5
e9eqvw4ixY7LsA5C7HItaKFzlTEGs/FCX3rU8ADEktIaJSRGFdu2p27aMhukNOShqe70NHt9yq9U
T1TOQo5mRfc4uuOqEhLMwtWLifW+9FEb7oiSNglpTlvobpmKOcoS733w4iva9IUPQN00zlx7uKvQ
Y2RJT3H9ZgiWhqornPANzvrVcHnXF261iMY/q27A8EIgoHMUz5WVWh4sJBeshMc3Hx3c76naiYlK
A/LXpIEQXY8rsWXid3HnoLBoRNC4GgNDv+kxyXJ6OSZIYcvUGY2oAy81MZz6GzK5D65uOtTEZ1Iq
KVH5FM1Qi08OguYMF5c2XjkaSo+buPMez8QaZynK2tjyd90dj50yjwLamGPgL2ntadtUKaORp8mg
+EapkScj42iGbdPXRVkPaQp8Wx5nKcCrVivW/QjI6imnWUDFnfhYB0aJuQgPkv7t7u19tu9sksuE
75fs2pGrdyS6ncIRtbZsEF7j72JwJKEv8RqEJQLOXvvHv1tsJVmO1rc5/f3ktMT9kp7GNH3YUbmq
L5F841zxQnSGCJm44Ih/wThXHBPu3Rp4Rw6dtZbp82OHQxr01K9Jj75GfodX4c19Dlv0YkqHXsWS
uS695cKmn0TNoq50pNoieTmW4MTN/E+fDyBTO6Ldem5B5OZ/JIQn6rVvYIlfaxOzUusy3AsVajMr
Y7w43ly2FCk5gLomUpHyOXTdZVsV5FH3X48VHX5jx08NjgJvICEJouknRHWotb5jugeb4yd1tExB
Q+Wz/t2FouvPIQGDHIrcLjBT5462bfyJlo7tgKo3G9tYOup8zmWOB5Jx9XpFZ32ooBFmQg3Ut+A/
dz5JEOJccSNVc1w19D1QK46Ye4HjAzcBTfrNa5sjxomg4hKr3Ei6rVDa4fVT3kJbcp98va+QHvcZ
DALbK7y0EcJc0OzPTicrhzpYKUy//ZzEdI5fo9xeTnWTXQIcU+3hUsInoUM33I/nOtsElc43EIAT
m9MeUHelal/FJd5uaoDmQ9wqJRWoCM92es37Ci2iEI53dO1lG9V9MFm+aWlqriP25O+XPbA1vI9k
oPhEye0CsjwQlYzLx3CBRgk6Sh2dcZJVG3CaOeCsuqTIn3LHBy502wdi3766bxKFTpxYmG9bo4Xd
jnJaQ4IIjw2TfiU/zaqRsc0rhCTLDpsFQyKEmMVZCobkY8CbdRHM7Q/czEfO7LLY8AEoChzxQPCj
Tv84uQXo7EGLLAzsu5eZRQeYRq0C2/jhPcduE489FB2wZryPnDrDxazEUgEfews+0LuVclXwpgOX
Liy1IbHyQ1GwYEwi42IZGYxsK/wlTGJ0rjpnUnCAVTMsO+7a3J4SeBdmpm8amh1mtq4+1srVV+3h
GAFH/HcseJaiK0FeVJ1wwNzYS5/qGhb4WlHO6QxyGXxSz2XG9LdzAiGQrz0HtqErX9LCHnVRKwfn
mNXgmkfm+3Z1MMPpKbbu9VB9o05ED9x0HkPB8YStqCl2xeCk43IBzXz2QkGcgqt+Rt296WuBbRWa
oDiVlKb0JkNvDSlmt27t0jKbIFnflXqcV6EhrXY/71TsijyIrEuGr0NEInlUc2itACeHtYt6/bfl
QhX1fTyCwgP5RQnx1B4qApLmxS1iIXjjNadm2N5eO/+AjGeIh4bYRK6NAvU7uOx4ePY1svbkxY1e
n3vGZUpw4BbUMxbQuswau2yVpc38FB7mLNKJXLa9ZGhElnjN5m9mP56LZPEhL05Qf2HjYC2moLt2
UOqg5uGK0oKi5clXhHxP3Mz5rwsgjrDMtN1IUbrxk+4SyWiAHNQL4BN9xMCYngyptZLsUWr9xyrc
gY7hg4PBShwfGlcQMcV4FmW643SJPsDpaRm8yeQpftnBoFdoacufjYy+GC1jcfuEy+7gO9nb1Ehp
B5dPPUuB7KgWcm5bMCSR/BijTHAamN262KSjzeFX4d7c2zrBBAo1YN9nkqfKACRfFDQU5WQqB+uH
+PGa8oCcujKvq6wbfBwq5mVHo6nAq7aemtzX4bTnWUYurNj47GLywaFD6Y04AUe5p6IDfdSuDeaX
EzovaD0ysFMrruQ7cm7swk0LejbLGxM1T5mBIo6AezHGd/iuWA+ERJptFlc13l9mcDsOxS0hd2CJ
og+JacgEsSVTgZQ4kE3FMSq+GSnDe1FBXbRMg8imPo62BswFG5NOA1p7SI+mPuuqvPjOPpDP6gyt
tToQXK20cAFAZlUBcN1NE2kJtTxEuTVp+IrtPNBoZw44luSYVQfgt9Oc1wwAaQIt+w73v0iVbclG
iKtRoGy6Eibp3l0lVXLr624Z6xERuYKpHj20gcAyOeeoFVSBe0+seHR1pJmSll7DIJvGnGan74mW
xy+xX0QuZpxdfIxgW4rEoDssxnsbsewfT7ciSsEh2N+FLCBdEDLCvXMktqSvSiTCqf4hp5A3g1w/
nXjbYn4rPWVhrkH3l7AK1eU/Hu9J5B3yRtGv3FJcvhauXsdozEZ6Nj7vJt2QjoKldylh+uo65It7
KSHMQe4RKIWgz9/HsQTkru1afyL4BX6S3U/i3a9K6wpO3BsO8QuFgXHjLwe3kJ8WV9qOZ1EFX+cg
pRpt78Dbf6Icxmc6FQD2kTqlEe5jknQDXT8W8ZXMf8yTcdbr3befORfHnYVcMKuq+YJJEnHUPDKt
y0ko8U6esKp7EPDesIMoNhMLEHVzp/qQuCh6rdWWxN99J94ZwhY+gBMC7oiiCUZnUxHFEtdPZ2rX
+8Fl4jOrTCfQAFEHZzCzjzO5Zg27B61GDv2cxIF+yiWzb2dyo/DBQODIEfW7/Nc43nLVPeQOFmZ4
uPBRAE7odwBMWNYthAtMerXDBG4yJxCoGmR9hdCZdU6r3GsRQCQcwHCQg+/qSp2h3asgxz/hda7n
5slp7kAz0RgTkSerkHXRWkqmk3xf/JAmnewbISH4oa6LSCBtGh8286AFXxlZjik//4nC6Sg2QUwt
Kg71gdS3vTBMYMwuwCgHJEKqNo37wXysUq1jMBOWttxZOVOIH5TTGWfhqz+d2Mdn1XzhbEaO34ZE
Y1kLzDED9T5uaroRwoBHgMQeQsVIZaCpfOw79yx77acOxEoYfSUoBrruf4ijiWvqSOPZ+7a/mf3n
0LLu32W4T79Xkr+OGcI9sRa1Gsggf+cIyjFPQvAcmpRbVEN7/2v2GApWC1brFD+JPDvKh3QJkDca
wau3BJqRU3ygSZGtKRG9NTSsjYti4541SXscy6TmrIn33olet2YQUe9mOBOCdZadNiMcFr5/Dhdb
SJNSdHg2wz4jNGQ0hvfLRaRONvCiUuexi11aXbjHbstZwcW7ysOVFcVU7pRsHQ6MYatPc8K1uFhu
t0/2ZAnH1Xy118utAQSorlF1AAoF4/RX54+DLcmEcAaqq2NYbjMjm9v5mcmPsFPNvGZVoWfAyrSp
Z9JZpWvv7C4Y3CqgZr+F1NsNYhbWsOk04nJT1zslolK6FMUoD48/9K24Uy+ozr9tMcLur0KwJkz4
nWc7bfhvANxbXt5sRS+XDJTGM+9yR2Fv9sFl0o0fcNbdEFX9xeYs4i7LJQZTV3RrCrMGmMdXWNko
oKvFQEL8oABga9OwGSC18U2tl6a353Sm+v8q4r+KNzv8994NOqB2nT07mBGV+2ewyspe3JyYIUgU
qkeNSWKBJR2qBYCZtNZs/kOoSaPlbuiT32X4LyhKKur8y9MVuC2ABeeruoVygundnBiU5DKMNANy
LGlniDDJl3xLkCJ65Ay5p73YjQCsZKe7iw2p02n/LThQavT6otFU/CqCSS7rjquf7DNpaqLqRVFG
jkcQ7qnOdOi2yITJcjGpFBMkuIxCuQNpvR+4BfBMtbSB25lYXR+6em5t5WmVz52dFTBtMpXaEaW6
KrMVaHWLnvPBIWFA3+WfjnIbTbW4pSPBK193suqG2A1TEU376KoX/auSeiXVKEr9B8p6S/HbbtZZ
SdmyClA1yjj5tGgo3N/8h+kzSdgi6uhBOWYbyC/QbCLckHy2XoIVDgWX8pjLVPJfrCftAQK/eCEB
ZxhnYkcyZ849+z63w1HGsA0VdinvJnOlkmEG2HGI51VzvgvvmCPcuvhiODsk0iRhsonL335BGdOK
S354pBFvXt7BmPkPV196YaoxaugBTJlT+qU2p5uI1rSueGnoxYK7jIjwGMJhHTgPipXBtJ2IEuX9
806KMmoxSTBU/HOMkJaJ0oCj+n0Z/PYD4oUW2N6MNAyd5oNgzWiZ32QJWbyoyd02whQ7FMEjx95k
C11yVLNfWi7rycRqjL8z3Yv1jzy/yLo7WG3N2UKcjVq6SNlbyTkg2FXkcDacDJoLDGiHlGmij3ew
Zo7WY0FDikmd5jHLFLJIzAhWl/FHmJ/KmontRA9e+fsYd0PgsnRI0XSWOjG/C4OigqXJyml3lYML
BL0UNhbENtmENmJS8vXR2LX3W14sQ0GsiOTijpy59LseqpHefq60K9y3J5yolYTZe9cmCC0UtzkL
tugKfdZEfQ2UMEMaYgA1ql4CdXOeAIdl9Bf3w2XkI/oVQ0TlWQHa/Kv5r4m7l+iBfPPAgHBl993J
zYCsCQ4/UJIV9QtzfNa2lqN9sMHWHgF4922tcsghtd/b8oaM81o1t7QStnlB9SI11TqrwMEfoiz/
R0lQlMP+qrSg+rjrxpbsaRz4LrsIY3wlyrBhazuS9Bsw2mKybZwPGvRXsbIh/JmqPB2pXE71yOzk
Ae+WGK+39otMYQZmEjuPyMrrxibeS8WcotlwickfRXWqJL6qIAdb4XsUXMq4VWBOMoSku+wx700x
ZInZWObahj9ODDdWiOfF3gqVdagTI9Ba9ExzP7wn/e/iEUqdyCpPyb4eXKFq66Iex/6WE3f9b3Eo
EDv+B6XzjAKxDb+PVHJgVucfY9SRieEHxLXdlX4fSkh2ZGzzHBhaLIEiMRK3hFtXvv6X4y4wF+dc
XtWgV6oUdkMkJJ3HwDBRCmL0fU1ZOb3adA5rIuzqjM3Upc2/LH+7IYUHivBBZuBKtFCxuMPhHSI0
PlOmSRdY+Lpsy19Ct5z+djk2Jsb2Ffv104aSbEbca0CfNsHK6Ssj7DB6NDQNlT2LLmVYxz2g6YIH
uHJNxI74gjzPio9HoMb5UEFJOn7xuFjjXei9vVkyoz2DHpDT9VmJ7aPvtgjlSf0QTlWn2FD1jvQE
WWW3OCTa5oKn81v9me0syvpb3OjcXlPu01rBPfc6VERCE+SmlTMQ5gz+oW/LoO/ivasu9zQdy3Hm
KpHHRdQZBxA8tIknQ8X8PrZl5A8yGFUUvRiSJkbEPJa+TTkiImICleQIgLz9Y0ImEvGxYs5gwy0K
Ub+IUsOBxeGWqBypIm9Anu7sHFr1hgQU8SlST162lZcQDdlKQSUOIp1WIQTuHtEggbnSXUqkFIKm
5cFq01Wkw31JloEtFKP4j4XfwH9LkFQGiAFWMlrhCU2Jsx83XIbSbgFdG2WCEfk8jrHJqqUCOin1
SHrQ+He+EyL8pORKKuNaZpVw5+fHvPLBzMDUZKSPUt2zGZeHKCr6GQVZwZkfLhxTkMrV3myC6rnx
+3YNqpQg4jAIziexX7OdMybWb22NVOV7swBApErNQcHj2sBZ6Od5sKcBOn6vUQA/Lc1XHwYQ4X8f
k49ihBgD1wrRaKBIdenCZY3DUcGMZ8ed6QINNchIkE2u5GMTaZ5bIEQiKPeDzXt3mhhe47Ne//qE
o5gOSxesyISnOkvV1l+y7VJtmzH1A2XjNIrwAMAQUXYBDr9ogMgwwvMxg0IURVya8e9sy5/4I88L
DPo1dJ+mcEGC+B0VNsJOCvx4yuqYxfYxVHpoI/Qv+/SDi0gTqHIa+pRtRjXZeoOQE6k+XA3+SpYx
ZFK9sSqxZrXv7ThNLDpEnODcFUAH9k0iMyrX1++JKGoAw604cQTTqnRQtbKGB7Xkjgei4GEbl01l
JaLLb2tgxv/9Y349+0j0SfpbsLEdDxnW3s8oY0Nub8kDqbGLyUlLcLa1QlEk1UMmsZjQNgTI/JRE
Q6+d9hIK7vO2SmB10EwW9aqVVvDvXSF9tN1WFBT9GXOmX1o9CO/irC3BNLk7D3YIW3s0Hetmk9r8
zYwexmu697xE6VyUs5BDLmQbksownJyAMZy4rTOvWW7ZSvXXxU0dxCAcFmv57+FChinAYl5FFZ0k
qJdtp2y20pKg8oScvppBY7bMIjQsfdizLuhcIzY6HIhrvG2LmC+JUFxx1LLTCoDFsWBTHMDMWzFH
OU6wjLpHQQjkp8HGSN7RpCZpz7njT/dLURRFm2txXzhpQt5U7z43UnC939bNSA/PqoLPeRSK1vHq
UvYpA3A1e25nU4DtkcfiyT6fAWHkP1APydvmC9sCNcMopHvtNYgs9ybskvKtawVW8ISCi6mNS8pJ
sykAA0hhMAhgEexs65fopYPCvV54JEhTW0uD2QPUOtWWXc/bGMUTGOaxlubyeB5M3UYBFEe3h/jr
k5ZGGscYVVyN5LZ3lDWlL4HzHayKFQ5Gd3ny6a6nmqaLTCaXKLVdRdHdQtyx5nH9V1DMHweOzK3o
VfiQMHFlMTSpcaX6AaKucCymwO762mSZfOE//i5/bwL2NgGZnnbCadF5/e7WNXD0FVq2g8MNPKTV
VeiBBpTjt7GjQH47mek/HFJpe/G0IUDLCzwrt0A17EcKNfrwkaBDn8aismXPb3GsLVwmzKjIBmym
z7EH4ZvPwHAZmOic42TGVka+KWipSi979NDE7hhadObqet22/TVZ4010Sl+HCH600OlODl4LaoYa
YVYBG5EI6FB5lIJ0L/VElSLP8yoBM21Q1BBMdZbJ5nq3KDZ2AiG9Y1qWchL+L8SMc+9lVRc1yj+H
Zmpx6p9NCVK0k1D89jpshMGYAyaA+iRPrVhWs78T+SF+2I0pRqTInCHHFZuSMvps5BjDiG17SZNy
awcNPpzLJN3BY30p/HzDnY2j+bW+xBxlUIdbM8Fe6M3h5CADAJMwVM/yWI8/lo8bZF/OYZomvQUu
q1cFJPGAW8h22NRnN2Cfg6efIYimaEuKkldKTS426h+/hmiCFlUcw9iLCL49czyjxXR8SnHoPHB4
Q8vNeoTedJYtbK98nV1Fg1QGz0U7t2jjfdB6g4xIegALOmj9TxPCYiky8MTncR83o7EFMqtleEBe
KHN2HvvMythO4Ofz2pJHwovSE4yUwfUTdqiP07Jp2IRNpTubPfwd4adTwggkoMwwkXyz28BE1ore
7EWySfGTirLw1OJN07DvzEVa7lH7yzr1wwxkwh1e3Y/bAKuGPGEVQ2ATXvUBDhmrUof7hInAPAPm
hqlMTAlBK+gXXtDWHLSLdctK/fPaoLXz2nYWEBhSwNUxUCzUA08U6WqEIp5+F6pv4OHcvb7XJLYu
Kn1ADRxDt3k19sL5c3CPu9zsHnXm3LGHZSjYdavIuwnodXC/hNI/tRzrzhgf7FAxoT9egJ6NGpkN
KeWhMLU6uuKFJP1qt5voU/4njJzxl7VJ44yqA/4Kc7P0UEj/8yUG0AAdazKxvnXrTFsVZes8/fw1
5N80cqRB80YeuXLCJpiiAWNiPIchgmIZ0FbRYibP0qduzqae6QjV+N4weTTvFrt1VfiV8Tvc+lie
5g+ImkiV5Wf8FhhnMIdBcyksTBSBttaS5jLzgiqMBpzOxxMIWocU12xTxQyKV1FtXVLr7xIvd6KL
qjxoBYD+qmyXwV7gGt+K3FB/nbis5hAlmHb/pecKwXPLU0ebrV07vi+ouasMXtL6dSx9b96P+QdQ
SkAMV/m4WxLxXFLCm/bvKxQYQ+NAc7BvQZweAkomP1DvjBoVpSBq2BsMzf3b/FcPqSNqjcDIlw4G
wihqKN13ilmWMWJ+I0ze7qyYXY2yFJtgRm9o95wiyQXCVblQIkxNj/sCCHgfR+sBo+a93GdDF4ce
7fnAgHNf0bbiwjZ1s2Roqn61hptrZLzxIUnDqfoekC2DQh39W78AHnSKA3WhYSOh6jbWi6cbxoLy
kw9zvqHEp69+oHOyyLCMFU2rsQpDL6FjVv7Aab9cUhkkSwHF0zly8/QhP48Csns5l98G1ybgnqWK
tQ+ahoRu6dR7G0QJXloAENLW9N2UE70NU4876wfp1/496ZLvVYhYULVlYKx9AtAY2X+UAbnxOjzz
FM01EeUzvHrOe4Q24EmWRSY4e5njOlLachPdZ+lP5n/DNG+419wrH9AULg7TIJPsSeuxXqP3/8En
vGRlAtT0FrHtOMAoohIp0uI0xdUd31s8hJkTA9vo1mpfJMsto9GBVeu6ALR/PoUMtFw3tqIAx1sy
U9AXlxGY/zB15sjSzzcraujGGUHjKy5eFqlaN3FXFNMTc0kxMtrvuBC3yi4tC1TiBC4QaNTVgKlE
IHNn43jJglHNV5iZH0aAMTyxwhkQrPhlSYzoJqRVigmqFX40lBYWBPlPV8NYmCM3/SdLotIph7Te
FJVUdWTl7VhM+Huj0RiVhg6YX8UBw2TrdAfkFHgxKekxYCMaQETCBz/mKTsayS80bPsY6gNoIuXs
oBmm39T+t63QXkT2xuhD5wsaFUVPWV0zOhlqREAp5oZmxMCwPenPjkS4EultFS8LwwkUS9+8GWVd
EbbWtiYGmswWbN3HS8U0Yy3ifRWih2rrbHyA4m4b5bEvtgho9qOrrpMb/o8YitUTATERUoa++pI3
OlBm9yi4u5DSZB4DxUwwnXD+j2dqLFwEm7ifkTzK345XN7a2OXP2Udpn84jlRjCEYuwQ8ewjVBZL
V5Cfz4+r8SpVwjafLlaUmzDgkbNPV7Z9qjWfnt7TZbeRB/Ks54bcJPsSu/7cVE0WP3LbTBuXwqNu
efWlV+3X7KWFvZDkUPfbAl9b8IkBkIhKzJy/lbG5NKvwMJZJLYBYVv+LeAPV7EYqTfhVRMQ42f4W
cXLvdXFjuh50mJtMPYqSFFTHZTJZnzwbAWYaeAsx5kPXOmBvlaI8KCEwVc2PTtevfSShpgaXeoVy
1XW+o56HQy3eN214sHCs8JB/7zrPjByFJ89g/Zo/rw6tdqA4V+mcU8Sd80vefqXBl9SO7QJvk0KY
kNBBVM+3gO8WuMTHxrfDhM6M4s7lZqTIO9/VWtJH2JddAUckBtFuZCjvJNR6IITG9pFlwT3JfVMO
lf/7BVarjbbYRpyyZ90BblNB5aBznQgCaMGXklg+Z0iJR9z4YnDeME+3NYdHXLqPItgVyKNY8j6b
K1yULXk4RGCTkOhjaEgYgPmMeOjJrEoFMtczIAc09CnKOdlGEluR6jXgPUSJlQgQMI+kj73+SpXG
EQKrsx02ndGujCIdx9bqWHS6x3La/UbTEY1/u2fJjm588zkIXKMWSMDMKcvhc/UXw7eBvyizHJnX
bxY+IWICi6iigmB/LzpxhFl3UzyFw+A3HhToxiKd1fwz7IcjTty90ZFnKeoovvkwJ8FUmDggP2fA
DP04DcTpCKonpmovQ8Trq85alMJmBuU9Ha0iZuPuCNQY7tMsZ68fVtiMm2c1i4zeDmJj5cXdEuNZ
gT6ycGRkBfbBqLqRZCPFoVVz4jNVHI0g2mTqyFob8FUitC53Ro4yozOpYlBLzKwucEfxhs/BpIm9
DnYYUTJ4AnjZRAnxByWiKoX2+hC1wm+LAyMOK6Z5MucQmWtJ6BxuM1hsOogtChov3Wr8a3PDV5Cs
ig1NcKp68+YPYLUFoXpQ0LGeXwPtkeNCMCbbr9jeJdXLnhIsPRrttRppXQaxmIeOwkYIe4NdbzwE
jeKNu+MAwU19oodpydeWionjoxkNmnDztfHWnYw7H8qCj6SlTGBdoRaiju+dOSXrJzIfHvVZozJ0
1ekm54xE+lj/ymbynyq5nh/KkgReI4YK3aVpgzgwMAHH/l+0+3YAC9xRQ7AfEt3EBxda0pLQuien
SJE2F+nB79qiHj/8v6NfcgvuIAHNN8HrIeyVSjxTYo4oeedyOcYF3SjYA012OZsBISW7yNmvYJTA
c4hUoapbKrbWnbbQ2W8rWfuKFJhAAj3V5e/MHCRG796SVLiJD5zTSi+h0owtRIFJutSn3ARfKGXK
kxrrRhYe89ipfKMNHs22ZcnPm3wrS97rztnOtxuFLgvMvaK01Jvr1bLbnq9yHware5F9FAc4p0Qq
1s2GRVsoCZDQqoX1zs9Ss8rsw5s7E9Lk72KbOU3mgODwd0voua/xJiyBnX2P7SvvagPvLUZA4ypO
CPT2scRz66i9l3H/CxspxI7/x3OcXolN4VSUaS0Dz91JacaLqpwJ77Ooy5JZzCTjrvEWwvUNUmpB
LZcrEtDOb1TkyZYJuaFuBeaBjg+z3l4WS3Ajk2e9KN8H5Vb7Fs4cHxJFPNz3UXEuxd7u2fJIhsoH
JnFrjBPmGIMre1njf2INjJtYwnK/IExow9zj1CbgVLDkhncxotOPCCf9FJlk8OBGTyqZi231oEDo
FobR+sO0uPq2jd+41dNgnHfwfCti59LkclcXdqWg2CR6SkH63baalebm9dEKoVFP/UvFBXdvwrdf
roE/kKwxu1F0TOj3pMHlR0KZF4oGzPphBYB+T6NpJGl4mxvVZaD6r8rLc4eH9cTpULrD5nSuL1cg
Q1hKdF9fnr6HIridcJqdgFyhf7jxJ4XEujsVtWEOw3VMQkypHbN+IPYunO6F3QmJr0Hkb8MV3cGq
d59Lzz2Wxtv0nOqq+ZAWNhPy3UrswaUdSRHZ5IbVHnHmv/Iq+CETo+mYPl4KhcdwAJvMuycX0ujC
U28kvtAROk5myygBpcNv5DbWfmvdH87HDJDRGBdPNiQsQLsGQratuyjwIH6PZmhfB3AyMm4KcinX
q7fbsWBr2HRYOGResKLjPQ5mdEnfAIuwr54ij21zJat3PcwOB70EiidRZXL6ZxY6qUuBXVhosyfO
EB6GZ2cYQllZ3nz/fCPEa3p8mJgUyvmmab/2d0uvVqeqixPXiGnVFoKezwB+zSlT580AU/w7z7Yv
J5jP4DQVVnNtn7gSoVNjY3zq0jVD1AQmz7eaGvig6W9ktacApAV1lCIKp5PYq4DD2YPUQFOwiy+x
TILPhRtkFZd5xCYaMFfVtkbkLJCJ2t8AbSQorFwZKi6En2CKkuxQVV8GvhmurQJl4sWKBNF3HVUH
ivvRvkm4UUWDhPsvceoAzQV9/RB3pySVaTPFgPdnoEMfXAhL6Sw3IXZOONj1b6SQ3hbHmZX0rR/k
1+YYa97nFl6JuS3J3T4KDlxfa50/a40ZrqArUk+Df74AdvR6juH6yRgaKfoa9Wax6E5/nUCGT32W
tVHpOI3i2owTR8nErACky4U/17nryWX+TpoKFN8O3hoByzyAqdMSIHG0P6zfoLp8Kcog205Uus4j
rI/iKMsJrekC69xyNxC1YRRgCtGc9bxsUmmgmuSU6ZtuD6ibX6wwU0B+XWrEDPWC/vcpSw/iu4+O
T6kE1NrvPiGZlNqd6+CkZNGpPH63a/OyCxEIJt5auK6Sgo5fJ2TvMzpkEZxTdfY288A4N00/6EJM
Wphzg4ntYMUSZjt29w84ylpVSHcPDnhl2zGCG+IUEUGMdrHfFksOQ8e8xkp89AwiFtFtybPHNd1G
vxEqLJmLFVQSaIEdfTiKhsxf5j3qPFZVTb0Lqn0S0kzBa/b1z23lZkEG7SeDGgQPhW3oMC3Ptdlm
zopPDPw3AIrYm7c0ObJiWQESTJcGeIOvjmQVmkYH4RdMA56o+4ifWo2WxZfFWULcynMyUlUU4oXz
AxA9yO5/XoPi6DxJY3p/PVwVIc7RhPNQRM+MHu/nBsdChsISPwnbNUxWp3dEXY2lEfmm34ZGwto+
vNrm9ogZyEfLiVB7jCdNFV6Gcye9xczqcnwZTYERGlF9EMnq33I67u+0XZui85gdA7GdqclNIl7V
+5JtNMqfs/1+Fm1oa2/Npx7XA5LC5SAeCTJqdjTWLfovxNWZEbkUTsJqr4BTGZvba9qeACNHKxsu
w4cKRQg3FndOyyjzPTytofoz9S6L2cjlNnxhJi2ESd4RtJJx5ApJEzeo3HK27/C9h2dgfC3Y1YOw
qFpiFITyiOtzU8ZG7e7D8hrfjoapKysxnXwdH4mqTUdP5F/N2EAi4T3QZU+FlVhJfPx2soWVWBUO
hRcaHzEBB32i/sjjldyoaGOhHGJqyrqo2khp6RggC1eQ1RMtXeIbkQChMMQwNzPWjWlzDo+KZLO9
vd78zlIitLBcs6s862mL+2rb61zbcwfSkpwtHsQAbVtONUG0gMkwuED+eHQVuXato1jePTiEq3QT
vBDzU52gVNw8CqAFq4pv7qaRfvpHPDCScimv4UQI9Jx8UvpJG6R7aHb8voJo68z/3dUR+FT7z8Mc
LTwXPhShDgRqOD+HfboS4pW4wmls6a7vE+hYtrrNqVwIcyN6c1s7N5+ql8vMvYt5sGo//RP9dmsX
LTo6wKDDlYuz9MAKnca7iyGldCrwfNdSlg6EreN1JatRE7kBSt+Kxx/tJOgRH61kOmcfP1jVRuqt
cMNhEf6zrIrTbUhkydOoPtJuYxl/CiqKdCe/skqe2h6z4tyQrLFbBs8ltTxSvawbMj/0T2LpymEP
WUDj56QvgURhuHpsEzKqBgBGKwyN7/hZLlAq3bfzHTP11J+T5jbDC6B9J15O8urPnkXYJwJdT1PL
51rCmBL/ugPKqjh/p9aDNZBVb8SGEvYnXLRQPyOPfNa/jFhZTO5tJF4i64mxl1Ey5eslZ8bRNQ8N
EesOVdr6kGGts++gUB7s8lOl2kNNYC2nxsucYqbCcl2xIzBjRu162hN4PzDWrFo/0xl/BMmX5XlG
a23hGlb1jllaeTM5Qg1fvKWQ+XDnDAhBKjgcB97an20SpRqy3WJQUc6wcNmgSMPHoacEsRtxo0f1
BtCFHnZa16Wn9GX6XIzqNIRywaYc353Ku9XB1O01d5DMaCVlHEGS59t1Q7JfgyjJhvB0BV/TNcrY
5VM+XVyIO22qciRz57NW7ELDH9RLxmq0PA7PsFv0Woamt371Xov11jLagc9jM+oZi2Y30LO2Ogq/
V7HBFNt04XZS1DSaL4Tv9nUDPHWpQPZXZQErAcsHQtUbs/zLsLGCVSsSmcwveROumR7Dsx/S71OV
Ua1bVI/LPMCjjRtfcSPySrUBBQWENZGERchbDfG62QgBtSavRQH0n7+BNQyzz7jGpsF8hUqrEXTA
pzCs+U56HxXJPfwb2JYmVsckLx6Nqo5b6T7i9BlWh6IAkClSnEWgW0+cbnNs80bYt7bq7wiOJ+Q6
xFH+FAQ7L/voNNOjGcuE3lazG9oAAOuUftmWrkE3uJK3Z59YFveUEOjGHAGt+ym//e4qHkWAlav3
PCDSn2LG7AvYeXJrAG0DJYvPJ+nSvk/WQvx4fVEzDIGyB/9z/9a6JS4+R0fUuG47nUewSYm7YIEJ
tW7tFSGJPm7LdQfOCuMX4QcxYcVrztTQw650wMbPEd0PNDVbLUd9k/mOmZXfE/nUno4m+y/dyxD1
Q6KjJH2VXl9sAFOCqYMWRzld/DMHUyXSRMcqCGyXhA0j/t/3BfRhwj26fH8WVUgjsrOV/bvp/gHu
/nA0uyjUAb2+R67oBni04Di6Qgz4+oSibt/bB0kmh+m9viOsj/FOVVPRnS2PqoNVB1Q/WJPVwIgb
2faAl2nEIEXlHQXU8lmfb20sdthXorBGQ307KBbvzXpPulMhErGAkkMrX0nPb53fI1p8/hONfqZi
YBUlyU38QKHcv9AzrpMqWhtICXz8AxKPLDXVy3HZAkCZtW2BpscwYjT/PUtx0pF3OTjqj2wL+KlJ
Z1zk1zGAkrRpFa+r5UeRpWsSt4oPx/BwcxMaiAg39Q0mUWROFIna7xcSmWR6Ly2Kt55arGjdSmkO
1/rnUHv5Ph3dMg2zvVpLs92YTVIBHqowUhLvE7nsmk9muylpyLbYIKVi0wPhiCFGjI0YEWW9TPOV
AepnSWhW4Z0rbJ4+eB03uXCdLne2cBtWNf7jKFRAhQK5Ks+fZtLRGHtgGwIIjHqa/OAJRQWQvMO4
IGHa1D2k/bhsb6FZrenwqQfI6kXEVZoziiGxNBhdhb8Lokfn4DvgmwQJS0NRbM0HGq85lTYj8mkT
RtTmUej5WV/gLncRVG3mN8rLCeAdwDjvthc5EdxNo54xGumUmz+k+mVNlKjhBm/eqtrxTGLu3K0a
LFT/vhid/Nr+ri14Ekq/ksZjt0jBBacRrFz9qrFDQWd/v17GxGwhhTdC6+nXqdAwTu4gF3+ZGWAp
EQk0rGlpWDxFz2nJC7oni0AGvpd4XvaQgvjcaORH/M37fsQf7hXvGurPuQQmICTV4a3ygIAlIKmR
Mt4JDJ2i3MewtEOvwdO7bxCmyZi7vaafdBc0u0Ia1dqzmAeIKe0VeYipq5FSdDJjJnfaSvhfqW9O
q7IgZ5H6z1M9hYasVqHZqIlkLCm87PcQlft+R+GD6gXblhd1Ix17SihB9DI7sBpFCrLX34lDARUv
Dv9PAyUWaEO3i09wv8e5TYsRZ8+pEH4WsePZXs+zCKji1P6S9dhJPwgMegyWz6TMECVHLBGWGMVP
dMEVYOp9e2JfqOwW4IB8zz9FAiPY7yXShK+rpa7yLzcEFBJjm7KX/ccbB0PiZoLhIl6zbaZaArut
Br4Bzysl/tZOW1AiO/GthfkF+OFxPRB0ilm6lY8ZHjzX/HDXqx7dzfNP/mDqJA2lIu7XiN7z5ug0
VQR51m2DH23J9fH3+WV6NhpGi3yg05ixGJYP7JEagIZQkjEswDH0CXjCEnu5OhgfXCjW4h7SQf/v
lqgRQf+Y0qFcxB5fSLTAFftN7ZOxiH3+xTeZ9C+wppwiF82gHbBe7PrYmJpwToeFlv4fARxhtwH+
I05pWQHiW9fGJlVHt2CYxChKJovdo3IeddjIHd6J/biqjewkPsV+LyE24CTJf+wpMJ/nKW4okgrS
xv/XlgZWN/NyYnohquQuMo7S5199ergxsBtL7EXcEb4a/sDje5ZQAGbJlbpiaDpXfBvMty1709Iq
Etx+qc3DgYbY0f0uQau0Ow+vi2eijdeRBusKU9SnqSW6gITtxVhaNXVzkpZEm3udRb2ZbdsITyzj
XtYh8vGZHY1pRyKR2n+rMJ4TfzvJ4ac9FcH++bZ4nkeQx1BUPpVazVwfIv3g+XGCu4qmzQfniF4u
f34U+EJsv0cFaaEm83pSOcuoeqIzo75TUsGNTA0YO8apAb4mwv8mXhWqeNuqCAZ8d/vayWQTjkbN
btKFmoX6uGS7+7KK7FUO031wen48p3mrK4PgIkZhAc/if40IXw9Z+6NFI8w/+6zczN5IXgHLwgje
6LPxva2P1f+M0cTzZ+yuHq5DusUOZXBta0awlGTxu8p800V/1u8YRqp7fFRifQc7J+ev7SQFS1qu
IGBFO9BcqQGUWcnNmiXOWdWpky4BaVHwQ8s2N6fHk7tvXJDLj4cte77EgdIk01kJklmESRja15zY
evuNjWJLOGj0pMwM7uhuSe5UYVIiX81Azq8WhjY5mMur+ndMSVa4oESoINbPA+ADcubk/c8g9e+F
rfeZucRJ/6uKGu20pKjAcise5Vod6f2IBXxas26laSGZjSZmj3LxU3jajFAKeocWyMt67HofPhAv
3+TdZF+je33Tphe5cExOK/OB4/Qrl7NIr/C8oeZwTt21SPHBXmOyeJTnlJqUIYdKn8WYmEVG4Pjt
AWMHsvJzsAgAuDAB2B/yXoMz/cF5kSFKGsugQVeK36U4X83nem6tza0m+FIW+v2thvVipEAA1ZH1
yPmIXPzwQ+F7fCE+J+7YqqBtqjm7aVVHexAQKBFeLtzS3dqCagp/oE4dtclciE703Qm33tQSrC67
M4cPdvkWBvaux7fNzqTxc8CpDjf0zIo/zXfzYA22Eubd9maH28mX1VtNJR8HriMiswpfQ2BGB/Iw
oa/fqrd3HiBxBHm8DS8tBl3O53Ddlsm36TcXUw+aSLSdNT+l93DjyriyDiDgeT5jM/IVal9BeodO
wrXQz8F7eMYSBuHD07ZgAiM9vKpg8Yodas/IWDIueBaW+x+OADYsO7Aqlad+aIF+hGV0EfMSiUxF
hhGecI4UR2XjOTOgRy4oa6qAulBOekvKmbB61p4Mn032mEthBASoIrKog3Oozepwv5elo3Ly26AR
EQrKWGibWVe6X90LncFtUprsIDyhyYPg6jcJ3zzmmd38h58Ywcnfk1e3z8UIAoyQkeL0P/1rZcdl
v35MgBF9TMCvqF1Tr+TDFVYr/rKPPhCDBGnugPatZ2+SFUGXO7zG+vE8inHfTvLTmbtY4gPIGoDW
P/s/Ocn6/8cFUO9X9EjYb1tmPjhZVIWRFlKWLWzfSSPuzxyO0Joqoor/fXyVaHdsO7fh4PId3+WI
rHFPrV2q/EABTntgV0tfJu9y77tQ+TXBA0j5bMVGQyVfCGyHoPymT8FQ/ev57eS1bWbca9sPoOuS
hADNHTUKFAK3S01NX/JgeecHBDuHbRfBQbVtxnBFuDqcX2lRO/2M1NAbJ537qqP4Qpore6yxmqbC
3cplRTuvbgyxOGcgHD7eW7hTCaAhqyw/W0Jo/jP3VYciWTnpSdCd9cBMgSiox4VJoNV5cl7d7g6Z
iMdoliiU5lRJe6NbPwnSRZp6ay1s1yFPgOByMPPIq0r+eNItdx8riJhK0/gpUmFO5WlbvSQk9WY5
8g4gC9xMR02XzDJ1rNWhZ18s9rn9dzeJXeZQGHiddwEa2/ATakwxAm3ndehJkt+gfQzvF9uwA1+N
6fNIaFIDx01r4MGJEXTThb699uf0AdFmGIgHPr4279s8OGu2ft/BGib7nwh7tRbcF9r1nXh5qu7l
Zh2RXYBTUoQy8GE+BLevPSJT6Z/of3QNTNKtK5tDHj0idRnmVYTH/muVTv3leFvC2mR46414lHib
wA6vB8Kas/cC2TzN6JKSvf7yQqDyuxf6GaRNpCa5AXEVgamivUARSN+pZ5ApfpHweukUuX98NOcF
4J45Buw6qu+f5nlu+1WW2xFAm+D1KAp2Mf0Q6XVV5zf7Xe4VV4uDn5aar+iKUhrRmi9P7dWGTsYy
Xel8yVIKurwh6FnriXx6m6tHegaMEJuv5S3eizitZq7hSAWGD22PvGdqnadY6CbJi1Anc1uMt3Ne
cAj2GgF5wd6oyQKs42gbVt6MqNzUvsZW6APz8CdQSg9tub8t9n0SZcPH4JVsSuzFfJQetrsNQMf4
0WpqKXoqXVJaMOOCEB7E6PnhI31CQw6fSorCJc28Fmu8Zr/aEpjyiAD0FGbV9LIRLqiLdaixgqEz
CPD+1smYdn0Pfce2OxS4cPleNMLUZS0GAHofRDX5O6L3IxzZM3px7Raijvg3sS4wcgX9sYTJpnXU
QixDDzyv4nLgziwm1/ny/VwkusJe1jZlsOJKRzt3vYMXcTjLwg8jvbHIedS9r/Eih1+hGf90VhOi
hup+nbTA8Hgm5H9QY4FZ5/wJtYKB5z/WW0las7WpMrdVmOT/8I0+qmlhV0XGfpwWaJOeCDd7ssbN
kXvdon1twpf3rX/HNRLu760KJ0L/5VHoF6CCRete1EcmH/zvArJ7D67stuDGq4DBaM7x5jcnUTsl
V88/x0iwo+tOcegvg6dbg7cmkU6rDkpyvDyXp/Uw4Fqyk33/+vtZw9wCIb2NJpIOXNHvHyPw42cT
KkU94YTcDLSouxTkVaNcplgxvRZjDPDgrekNjbAzRMjn5FkibcE53t9xbEpCLrPylqqa8k/q5ncP
5JGDbgod8g0JxD4JXJ/O4uMM+Zi+ucNk/T8F28rABKOtFaU6YoJxnK0qja8VH3lqZzuJcOxBac8D
r4BETJc74VCzI22hirQXHz3cIajp/qFtC+YwMzW/+lMzEe+jJUKovZNeMdPKrhXwETGrHo5D/pIS
Aq9G2A5+dU63QBz/lnF6AtoC44BXQb+Mpqgy8RjZpkH5fiKQaGmDMGR3mN4VgviOyhxi3C7E5a5U
rtopIn2k0zG7mrN/HEesKY9SO51nTjwxUVgN6YxNMDfKtWVMpBNdtInksAgUV96YxNusEt0/XfeS
6pbNWZYvHLJ3Lx6GuDcRARLMp5c88py6bnA/VGldfnGAAYbyqG/WDNoF7lTGk2rc6vE/f/rVEbXO
W8CGM8KmxtA+NusJ/kP8tF0J9Y39+c3StAS5e/ZnJ+p3B1rPBDfok0M5D6Yc2iY7o1EDDkPUjk5O
go7bUzA6/bC+JRw6O7v5W0WDlePj98GtP4aqtjuzYN/w+EteTa3ewIg/GMpJm7i/fZJeBjzZdBfW
Tc+teXeikTdXcIhxORlGGyUH08c4fyWjJ2lxg6ClpR3W5cmD9UrRhIt/tf8pzmoBGNmaXuT5kq6n
sTGfJbCHW0xvy4G760MqprG3/DkVTJAJnTrQdIAdH/xtWnTXzKSwJXV35Ina2jOg7m1VmtI2RTRy
K+KkF1R0xgBSZXSY4MWnUFaN4sYIMG0W6GvcM94QtSY3fhrLKvmgqgAuW00GsqMm3wwmStFhfylg
GuFcHcqcoOe+0OAVkV3GP2bbQV2RJONCAkKkTyRfxai7U76cfMIfS8GUO3aPGe+fRIIKTPEp4LOc
tqPF56wzXZFQh9+2K1DXE26exC9hUj587bG55s7PNpTNwiJxp61wYzsCboC9lLpLbAAnBaIAoMXE
srqlFAPnWGTPys5WIsoqhkU7uDm0dlaHev+biGcSDFNvgvuI3WbOJ+spuLP3LliggeDyJhkB/SlP
CiyBktINhixbr1/iZcIDU1IG3lC54rYzykKBpvLRCYhciQJ2ZRZy70brFYFRkjn/s9p2+yU92O5A
e1tjHXBHPI6txqgsJWVao6wld865RwOlehGnSX2CCuD6iPqoVYsTnhJlD7Pmk//rBoUButr56XTv
1ikxbgXrlbx/YV023k71VsQw679D+u3fYqegkVATSbD6FDGQnzVvJlItzGI0UbbyU4wOHI8VBZc1
+8s75poC1DDDHfRLO6OrRG+gElLO2AZAPskKkHKvsJ+FmcH71lSWWyi2q6oGyKkcy78XoM7Cx1vO
yMZerRpWsVgdSzfWN17fAxd0iDRQrn3doWFYGXOja/X05Ayf2E5k4fqckWSzJxRL4YNV7p/WeMXn
ueXWSwp3lFv6Yo92F39ekJ2vZj6EpPfU/jcoMaAuBS+GoV0hUjdXMoHXac3F2GjRoqq51BPvh5Ud
Zq8JuzD+Qbh9QjfQCW/EAn3xatPlGe/4dOqTTPUbqMSMUkremgeESczZ0I1rLsN7/pzM2+I/vaWh
k9ZIdFej7OvAM6BNsGqEff9ZvV2q6FYu8ObrXIH1o0v7nh8c/ZoNQY5S0iRtzkl5BZnFB0H+ljLd
PSx/UXvJ3BkIJrCROGYIz//9Qx/3j2RNea+/LdqwetDbsjTFVA+BcSwHl5e1PR0O0RocW5mhXTqF
2RjiOveXeNeYwcUKiEnMwxEjnVAEbdMMg4e02H11fpmyiNGtW9Ot/OPwxv8gOoCf4nV7/UR0QF4o
KzPIaYMBwKlnJSXAooaeQPANRPjCoe6NfidIyZk1b0WAXQ9274XJCdZV0ewhayyyX48+BSO77M6J
YvtlQ2VVKCDnhhVmJ2RevHU61EVb3RazQW71hieVdnlilEl6oXkARUqFDVVS0aR5X4om7mdZPB2G
q2IpwbzOJi3/TltWiws30ReCHWbEZuRid6mJwSjHScSnwecEdZUR3iCW0fuBJkuU72mWPg/2yWNv
vjwfhH2TbYmaztgu6yOV5wL6zlfQCYrIPkGOfI3qaePubot+zcioVx0KSKn+KCBgfKLsT9iko7Ep
wQHwwnUl50gqiY9yhwFOwW8/MG0TWxFqupAJ2CnR+MdAOwImtS0npwUj+ZfLxr13XbhCtWnm/DQt
BDpK6t4ooHmv025Ysjer4VSD3tLcWp0VmqWSKqEDueLgUAllkQnPm45gH1ZDXEBjKWN8YmfxP4k9
1Wp5gWgQyHtNfvKzJTLOWSAk1xcZDzx+tMAtUR8SfirO2x/BZ9A5pHLsWuw+1+JbPHbatSbo5LhV
uQ0fFyZXvFgZ2AW7nHIf0VebJCZQkdgR7TioZnPctwGO3LdRbgi3ihgTNhiOXO7PQfnaESaRf3ZU
hUogCgkLU6R9zd5HwtDGjJF5KN7x6ol0YLjvX29uv9gaP4o3SWvK9QE+c9WcY6z6g/+xqvIensKo
v2TJ43GYBmJcKJjMAZVFe3DZ1anC9Yt2eEPNybSpLUbcviN9jRYCdgGlysbKsPp38bVMVqq8TGu+
U1LE28eEEF9FPggQ2ZSHGb9JrbwsmI3XNkPhnt3/0hAsvPFJ43kUXMAFlKS+1YzlcU8PamjCKQ7a
0pO+GGZa2NeuDacL6Si9mbNY/m0SPduaoxLZ7LvCgJ25dzo8jtSTYsDcXy9NfqdFm0dP9En9urSI
yXN62CTHwM/wz5pGi8ucuGH99E4BSKTdiwY0JR7pi4qYwIm0ixJbO241NEYjLsLinjQv/gYHxu0O
fCQlcMR3/eoHe820wdLHfQAHDiNdxg+DlAuiifk6vSGTD0Zmux1YixECgNubk++dTt80bDu8joCm
cypi8rWeH3VQF4O/JW8Bo3boOFDY58SNdbDTKqcn2++QD7NmhtzVKQH7zC/eSXjW0SmTVIQ8lRL+
RpZBiGCGoU0NP1h7KOBqYDgDDecfPyMD49Z2xTo74PpKT4FgSU5nNJvYuTHc26FFGY4NvVlthvKY
Vdj5VOJxv2xwiIWLojas89QmQS1NG1T6Bmd3mYNaeiWoSfildY86p1ISQh7z+j3bMyHl3DMqq9Sc
MkTha8gzkFy+U7m7+i2hDjz1x+mI4ydLG6mBzWKHonh9qYzVrMqbxgMTQTsvRx9lUHhcsmRfRICz
qPiOhhv7eUOPbwn2Ois31u5D7eLlsktHQ8hlPW3Fz61vpWw8eCZVmen1nocydZxOHnCdMePgm1Dj
6/FwNOlvwdvUhygjOQYLngJat9zZ/1s1pPGzIgzvNLzIRy9KeSvN0gC0VShJYjwEUkNbr865RpsU
tlh4IrLpNCnthlV+cZ0SF1gij9024hFSJ/2FDtZsSQPHrnrwqL59JNVR5a5KKUCvfsKJOBDPjImS
FrGMWr9dDM8AciP4+PkCHtnKEb39GX72rlWkq8YQMVNKzFBPWSbUL1L79sN0x/21MjGmf1WNZdwg
e4fnTlRSLx4YrygtZoD8wIL4PrbcZKLl7Tq9UemxHT0jNMNjKw5hHZc+JJQn/S/AascasKu4mc+T
1u78Xi5Hrr3mQ90hTgdqP3fokwwFTUXqrGRBaSCNRIjsodnqQFeW1Z38fJNbAMD2/i1kTuux/Gto
alPlVEkq/1n5CPVPtFiPnTIB/2oaiG1usDAb1vTkvU7bweuGJMevhHt45kdnoLcQjlvcuqqKeMwo
N3/26ovEnG6lflOEyTieZD6EN/scYhl8NMRxuJgjXLJkucM//vgHejTeRj7ULQv+K4RMWt98O6un
dHWVAmjEEUOLhIs5j7y6rvsLrGmGcy1fmNifVbg+LkAC19I8GGApbFvDLBIO4hWTyQg7D+dfwaOi
mGF/zxqbaT0fI1h3f/gM1ye1DDwyZ4/BJPeTkYnSo7hgiN/T43xrQ2qA8Nx10LjVir3giVt7QQXR
tQQPzIKkAGLqp5022WKeasgG4CQCftFWM22+oaDHToX5n2KgY18MTnGR/ebqc6fieXTcwHHae6cr
vMWUUtx4GwhkbQi1e9JS3dqyIXRw1X8HuNz7fMtLmZ5bovDAIHOz4IiRB4x2FuAOEEduOGN8OzTR
m3DqIZl2kG9HWRINdSVMqdFJSdX1lq8jGAFBJHJPcnZW4WL80dv8QDUVL2yOZsFcnZscO2feRCU0
7NzYVFadLaS7qyQgV1XNfe4JAarOa6ho5ii4Mrdre32PYM1voqOMdwK4qBEDqZs932Yxk9QwmdGy
xeX2E8Htd9Mo3/t0S9qLV4FJCyTK+Hm0Ms+kObTnxkzTqO/frVhfgbUrWizkge8SZj++IMk2lVVP
dPo76h0Qsc7OfL2OsKFQqcJ4iLKJZkQl151GYLYm0icCDHPPsue88hqxh/6YCRGbMn8xdDBJ5jqi
v6oOuZrn5zJ9ktIyqOa6AMvNFrkJyKFoYTHDNMQ/YRxlPaqzf6EYg7L3kIMD6zcxaJtzwIHP3S9O
UmmtAySOAT18xiMfrZmVURNPL/YstjbGpUo5eAi1oZMGk9zGQj+03LmO7upbPJNMNqP4l8vbXooE
02nUvyG6cKU+QKTtDBIM3hPKu3EE/I8lzkGBnMtoxi9ajLkHvKP+e2QU6N/LiZaDlonjH4kSipdD
dU7uDvGKRQuWt8hxx950CiH6ywt5AJ8g/doR6R22yTkHM9g/rQpgK4SNY+ABPrWBF53gDSLeNc0z
8pgYpkCKMq66jiyYZUsFHHkeEyDSLHHvo/dEzbLTNbl/7H3bPgr4gnWpMIcAkC6WqnoHdVFAGErA
tnoWJw/pmveWMKrMaVtPLsmDF6D71BC44af0Nucqor9nBX6kYukuIwPwEJ/+qf/gS12oLWkqy4cp
j8yS8MxpbW4VOdO3SmMoCNLFKPLRM+kGVY6T/opMyO8VuoqkTUglfqKOEcrZlp8xTZuUxK4fPS6F
NReczr4MplqqEoiETkiIxEXvBRl9EEs1iT/ApKfTFNZlnGs203qMX22QM1HCefK1AfkROCaYObU7
VhzblnSXYoa8OpGQQ5vaZdbUYIIIWfCa6BInkWySqpXGlHED1zhVCJ+pQQ1LJbEoU2R342ooSPfg
FhUDcxxdGun/J4UDeG3a7UPp4jCdgECnpNyEeD4RVxglatmlQwY7hWGetRF9jY30s3gDIzZzwsbr
HmBQ9aUOvBGGfZz2N6u/INRavMHFWZ7anapSbMVUNq/1DHo0lgHD1Kj4h1qMyrYGUQfF/brKMMvb
fkUe1whHhbVl0wzPf/YRTa6YtH3WclrNaj+z1TYIuH9yb2x0PGowdom83qzOzSe+YcpTJFWVgjUl
yU09lhOTSwSmt5f5yFrBBjhGmYnI+BCIf+5pbZGxfdXtquMFFXjvy11jHvP2N7y411mn9xKacVmx
C1PUT4gosO9hmayERwM23sGbM0q6o+Rw80r5FeDwXcQGPUc9QbDZifSRwkp6fL+h1xctKqJ832ww
5Yew2toXojGJLIxZmHs0oYF4h235Zv7Vww4rRVyN+5b9L/YWkK9tH+9jNWwnA5ne847YsfKB3J1i
WqO6ZSTt6ta4Z8TrwckgkvpCmDzWbqcNlfuXpCfvVxgwhoGgyK7tpAYXLiKt5qf2TuTfN49s6ND9
Ymc0kDg75o6QVaZO3aviGilYkAI8tGQCxzrKr4H9xUoKkVhq5LzsI2KpABihzhM+/jXDEwVyJSJg
YDdXmUnEHlAUAuzVo01iwhcLjsbAffncumdhizQ3E0ZKOlu9VSgNi9qOwUmOcyj+df0Umat88too
HYqsjClQ700PTHp2uOOgcf1Qdp8tjYj2qoy4UTsD/4I7bsxc+NkgfdbeX5AhgaWnhFpH1Ukbfr6P
St8PGEFfyUuOHcNIRHf9WyKxHGTAaq99/jVXuGm2sEL5JpOPXmLOzuymNAbqsrEPHkJQjhF82kBi
lOPWAAZYJ5NvZjE2unyZk9Zh9ek72TL1dRaQ1iCFENqJ6rfxFxpuk2AEuEzmH0iR8Irf1y4eR9Ie
C2uSyO7QJyXvfew7aRL2tYF1lXahHb66TXp1jtfsD3CcN+ndCY6SoyOEKPfvOz4djK+CvC6N3QGt
gHxPTHbLn/1m6gR9Gg1COiQ16mGJyK01GsJoYbmI5t7TMrI54n42KDn2zJlK1dEI/joN9gqh141R
ILVPrFCLIbFLkgvDNb0WS51u2L8CxBZrovnrXVzTb9PfWILc1/RRLUBf1TUcokbgWYOGgnrDmF7b
+A9Vcm/o/Co76sTh+5Ldw9DFGIx77s5Dh7jZ2I0nLnAIh8Ry8dyXJQDaMVR+Y/V/hXP3GVGCQ5nb
9f3cU/LMHtpnaEPuNhLgek4EaBvFdtUWduVV43cA0bMM2JmUtvePw8y2r0BNom5LbDbfe4I00rZY
JadRDlkvP5jzx/Mo1mQ8O47bOonGdeKyEZgEYjXivpBwWwvNAMWBggP/eNFwoSi1ysBOvk72kl6o
QC2jSZkmeg67JkJXOcBffSrm1pT+XI5NMdb2rSu3SeiI2dYq6FpXNyJgYAzv/300oGFIkUAoCQiE
RB3jFHrpjnAlza70F2rB720eL0LGk+Ow7CEflMUdYCBqNrzGMz5RQCfKTEnxytdIsbgZ8igzGnzx
s9mcucRt2yjClHF8NrhPH3LYBVMyvjVZh8RsPYp/lz73ukKAAh/4rWcIN/3yI6Isjzvykg1xS6Be
usWEc+fqaL+deTYnb/8Qzqo+1eF5W3HAjkyQkSvsUjrAAi9/1vW9XVH5aONrx38QDt7EYB/XsBe5
JNXLAhSbXLVJK9XDPst7VvXk0fwWnS6UKM4YLlkC0ZWvtI9PLx04UTzrMbXiCnNXmT25+q7Q1g8J
eGnZtDccTiI0q1Qy6lBnIoWze1U4I+XFEb8uChdKm2TQo9VViTcaDjOTAX/wGTwfKAFzDzDcAGpJ
hpL1fqbB7IKi0kHFQNuRHSwhRUJh7JX54y/NLoT61rdzfKET+uHoQPAE0T7k+v2+9zBgqsD/q6u+
EaO0g6Kp2RhLXFrNySLpv6iyyX48c173xghvzF7AaH5ExIPdYHkbsweZJGtHKWLmB4Ze1r8YeC49
r+z5cVr+GZqXfC5c4wFq3/HtE1KLfw+N3OZSmH78ksWI+2Kno195YCufL638BCIFXIZ7pb0/ioM8
GI7CAqgXhA4sXutkxYk/nSU99z6a8d4n6ro6h7ApQTlwEUdgeSvhesnEfSTkAXg7liUDxTsIMHk2
4AgzWMiiE5+aULhQTsjIEStdgB2PHLueKe8/2i1ZjOBT95V2Gcw8iXAJqSczePH2CcTlrukc2XHT
QBVSlLe3A+rbKfAS70DHJSrQOG6L9bD3+eLyOOZZE5Shgr8SSZY9j8tDEA6ZTvAb+9btn2Z1fxpn
oBB7mJNvvjPtjY65f/CWOD+KG3NPGFcsZ3FKou5QOx7/qpEUctkBi778mL+vAW0DOkfq33cDdU0Q
4sTkzI0U+zTMbyB62r6IoT+ZwCIBWg5vYjCZJLf2reTV4QcR056YcNX+pbKSYP3/s4Qoj0sZij1i
1WW+aEMVacEbwxuhymgBhLNqd0Vfta5GZbP+icWLEA4VnWMk1MxH7mUa7jZJIM5u7v8xE7NY8Clk
S9a8ss/nPw7JG0DUvd8i1lcrgisKsr+GE89zAhb2GLIR3hn4/nVO8q9JvZ1OEeECk5vW2nf9JObN
MpUjpAwwhRpbfq/AIrcUyQMqoIDs9lnVOKCXYWqR9f/p28tWiihJ1IootSrqWwnO/vrOB18PxIHG
0GGu3bEr5Tf83tAO9eGEQnAQSinAAiGjt1RroquNAglLgLQXVdCdVz5RdBU7mMFjty7phq93LOz8
yHUXjvksGcyWwaA73NQ6+wrAbWbxWH/zxV4XH/XLvI8N2jWaQcmX2YTZvGEzLYkCHb/tBWmuVRSL
wsP9Nf6KapGBFPt1iFO4nodJKmxroqlK9tQoKrPknG2rAl6ROYABfZ7uKgWnB6fbZdAULR/pkSv9
omBbZB4g2JOdU//Vz/k05J/pD9X4GChpHEDyPROirGFJPDSi6oR4YjbZD7HYHTyTmCSqv6ugL/wy
klkiY5kLjgpBqpTxhgIOmPjeDn/Q0EzxcDEUuukh+sM91nGXG+Br3j6/8lYuU9TJ7f4s9LKzX+fZ
r2W4Z13X0D9cTToqiXewfs/4jRIm3zW3j3s6D5Yt/Zm0R6fnCmsMKm1jUHMTyhOnKF6HW2DPwfn7
R6JmtpP6EC981h0vsfvvAupmhCn+R7s20bsrUOCEYtWgOOHewiza9VO5E+KoqMpi/gJYK6AY7gsC
OGwcSMSSVHypwvcgod43hdDUFHqOsrloydRfpywv7rcbtT6lwnwtjjlwJtj27b/5XvIIDyoK1jvY
D6Z5tbtkJeKelxPu6sEzIMHbCwcweEbDSQB42Z2ede9Ze70l6241qpuLhGLoRPfK1TGfoTq6ua0b
0T0gLW+IcGLcQ+faWqsQkQOGe4uYQo82x3cwaQ65LPBJg0DGHgM5emSibPCuS0RH+OM2I2FNQM5p
TxurwWdFAHXDRrLOID5NBSbWvqWm0Ds+BrZJ+lbqh1G7APovS6tcPdzYNZYxN9+94+q1y2Deius7
jI0H+HXIM3Hp7O4IwblpdRX4jvkx6kN01fSk3grrPgHDQ6Js6YWC8muQNm2GFEjchDVTkaQgDhm8
Oxrpl4f2Tf8yIW+FUaBMXgR0hKflscAHBwXI+VRAXjM36V+jfP/qmknb7yE4/iUU017YZAH3M4bP
nUOnkkBIsAvXJUmagCytn3E6b1TTye8w/fVs6e5AzsCYb62vd488YMcOVmMoO02SC5wFJk4aeYLj
5pI81+7Yw6rBKuHVRUPdGJgLeMYwDIDZflUXLJNQrL3k+IuSUXkP2yOCuYTxsEjufG6L5/WD/Gkw
M4r3Zlu9cKfYssH7mzIalIRL7lJAqiFaMujIkJzbOfErW9gC6qBQJNOxNBeb8gA3JmaAzt/8w2go
c5swGnTSN4wJGzvIe2C8BBSaxVJRpacJAVBkb66xn8JFZN6fkH/sRJ5TdaZF52+WP534ST73lbgW
NzxlfGUkHJ7Gd3ls6YUKphAgUZVgj9YyCixF7hGybmR0U6ivQlKoE0qrxWh7iGx1dV3DnLQL/20E
692AREPOZsRWUkkpZpz+sFvZbuHC/8BJzfZt2Csy0MpleErE+AkvczCAzHNc3dCM73LSAmY1e3Y+
Fe5teWV3wW0V3BglxdVA9teP9zj3ArZwXGw0hR4TRg1bJGi7RUfHHshfISheuiKp2FVLzu5B1B6r
GO6l32ejzqYy+o+6aW+tICcB5T+rRt/IKCPS3GW1xjf9bywB9324u0e/c4I0KoUIoEKNu2GKAZs2
18uRNgcDW96xFOHoIpw639/deseRHPYZnYRwY3LCal7Bg1rc5LWRXXVIDk9cL0TlDqg/AUZWlK1h
4U3RrBS7MjQAKHoml1vR/2ltH8G+KbB67IBNYBhtcS7uJyNtZgxTES6/6zYEMizeHS6UUIbmKOjh
zo07RU/v0O2j2Cw+3MXcrrIK7lhiMx0ExBEp0UDykGxeQYgs89+u7e1P6jcTcdkR20JO/uc6tOC3
7wHcIaTUFVKm63OF3ujx9CTZLSYOz8tko5xMDrpQZVYhIpWtSzZAot1OPnAjpqB75Nj4vCkl9Yn4
9zeYYpmM/uZtOagBDzqsJSCSuF3sxp6AJn6aO9vazk3ZzOQb4im1Rg/n2qJc1eIAOUTf7HAQ1+nP
svCMqvYzPJjvF1Qs8VDjBwQhK3zi8GbVAfm4HnIRimBlBH0eDXZo6y7krhPCbG/0+eZHqCoZbm1y
o/0SZP2+s5O9eeRvaaOCdqNaCnv+Gw7TrS6BgMCT4fHt6Z/H39unRAfWinojWu0hg0BXAc/S6M5x
/erH7Xw5olziuncYi0P9g7QERrnS46SoBFiopdYaEK+rA8Lo1KOcdIZvjQOpnHutdL4LO3GI4fGM
HiT3yRuW0XaN7VNJgO0qY3ymS7enoFPgze7M/FeLLznZPAw0mlwqfdsNpCFZYp7h1hJy7nJ2xEdl
hD5Du0wd4tnIg+odtsvQfAGZc5rMpSGo4lxsH4hJ09mAuxXp7WR8SH5jYjUPgciTwxa/Zw9BLZ5W
eX+y+EPn3tP5iVuBBqDIDZyx95cQ6J8xWYOeAEb1eGBgbKK3JlZja1+CA+O77W4KOWSaM+Flj6rT
hkr68FDQPI18bwIYL4zR51MnKXdszLMyvNF1a9cQDthAh3CG/U4Qog/mjljjis6Z9P1KfiEXT+pZ
Q4Z5Zoip0MPwFk0jATYnv5EQNQzvJApAihdIujVjCU1CyxTb9q59ud5kKApuRFLB7DTZCqQh+5gY
cHZW1tBtHOE8aTarSExQs3UesAbCYf/dKMBZniXYFtx/caZLK7VK0iT+j2tLBLQ3iueR/suKBm+m
HmiE/YeTFISSdvmvvF3dw+nzuxZwSl57TmReycD1z9BaKnYTMsxBo4t4VIFXAi696UeARJ86TZR/
Az9qVp+L7JCZLnjS04ATMhMYACoQ4hgaIS/zO+gNOu+va6e5z07e6aF0xJm5KxCk7IF3R+ldktH2
0jX6R/2WaXR4TEE0NaIAR/d+2DP4ApFdYSGDvQm+7rezcFP9cKcYmGo0P6SiJGn9XA1fRM0UfBEh
YjEQnv6W+P4+LjNIvDGR/pwNswCyb+df6MfHgJwwxE7bIzxRAwEC/opfmuPOu2DhVfTewa2WHpeI
MuQH8YPAo5x0+QCZhxFsdAaBmnbO86qksq8upOtLn8BcusixLepzUKJBmo88kKy+SeHv8PH7stLT
IXKf6D53Pk0Yszp6Of3e4rBFmpxHCc99WDIshIk90SlN8dVKA2cdYrXoLGV9ul/nfZGBo1JJZDvd
6VECq8WwPsrsjbb26DkhFrEvIIsGhwcQnIwweq4/Q9VmkE5fO7Mi2Ync0fz3hOpv5enifjWvL7m2
AE2+D0/3RMSLApO01EmKgIreldL0QojbY8ceY4FmkamoBz4Vhxm/gTI5r8n27zkkD58VKZ1lCTxP
RleMjiSRG1oI3zZEy9rjlbzz3lrzuaUy+at2Sm6lYRVEQsMmNLCVRvEHK6wb5Ondosi2q3jOIxVO
Cw0wU8fA1ZCmjBF3i8dM3GbrKwl3dLTnPpTnOvvAO4wPcqP3P7t//WgxGz4ITiO4+h+geXVGtJ1z
nE30JALABgxtEYz1aUo21mR7m6Z6Btq592Sh+LPWpt7fKrh8HNBq12TMOHraJ60SzQeIzNx18/W6
9wqK2sHSw+uQIoWQTU1aS0u4x28xg7don3vhVHoqeyeJiTrfk+0wpqybiP46vtRxd+kpSnacUzMv
wBbPs95j8AP9KvRecO+6jybFH5q3WUffviBpsLny/xiP5773MKKFeyoKuUi38VZuJZTdreB4JFzr
0/o1rAFmULXtfRm4vDBgfO67zZ/sdZ9/J8Puv9q2K/5yaQLYmce4ETEQORjWSuRSsJ/m3Gg7dcp6
8Zxj0j5YpBQe5aOJOaxzf2+D4V9mlF2+FmuDT0pCLSkxRWXIVlHoxAnSA2POGFPp1b8aM4W9d1KT
BzuiA9IpYKV5PuGqiBVnDk3STyNS5Kt3xptdcTVY/daHV5nztnSc14Kdn83kWl5fHNhVIdTx6zWx
WvBP2lI8NF8d4U8VJd2g7/QRujqIbru2mlD0+Xvgf2juOzqxgeApN4CgkclSPajLSQCqPpwTGa19
zJinMEr/yBlBFR0lsG8pMuazmsDilHbf7OTXh+p6RmRj0caEuxegg67L5VIqloKRHwVY8IkXXNt8
MAxyXctr9WCZajp2d163z4XuSBf0VcbWWp4tSw9b+6/6jPy4swp51KHKiw51sDacKoT/ksKkauoV
nT6N3JsaLGCdJ8q/5reLWM3y5BUduPLfpaJnY8yLSy37AsRHedVh+L9dswNNB6wMNEYBGYMD2g23
nyirOqncVCscVQjS8wgyjVnDload1Ga/LEP9/Xj5sZqrq+/8emoldhF2hgmO31Lmg6GyOiyuGYPG
UWxKudyvzGxRzzGGeYoyzLlUK7xa+IcDOG2yWVvEVe0r4BzwzTmOTfWqQEEEFBagBWQkpdngrWWc
3OcICZIR8NRsffh3+YxiBooueKeFBr2QtzlVicQ8TbuSA/uULTgINTH6hB+MR0Mfl2ZZXmLVpW8g
IOxO4Sdybe8XD18lkOxlUN+8m+U9RJVJLePVBGslGjEW9wzTTKwh0e6q46A9yg9j0HQEgF5yhor2
ZBMIX4CBm50N1UzUtQBCE7fSn3XYnbx5PFipTVgLmuimsRDYfZqutOu59YGuGxztlxrylGDw8MzR
OcSJ5Qt4IZz76AlKKW1K09rqnIEnmzzdVw7ve2kjxFegRUI4eLNAsoFtIR2k6nsdCbyrQg34QOzp
I+XAI3z2CTtaDFbIlgGmxCmuKTXG6oVhGpM0sqnyA/2ydSuY1YbscN7Hfr5zyeLQ5U0xQ6FuJjff
qL1zZsOJpD13iIPddz8gUxdZYig08w2ajO/nx49wQ62iQx4YfiR/XDmwtLLTB/PSq/XvTmeHrDLZ
VazMXFUKeWjp89l5fkGmmaxZcfxZb0jgDiI4ElSxqyv5BpNTXnbw5N9RoKjxxZSuB3gOPTJkooxi
l640QFT+CttQvN81KsbK+sVaDqyzDhYXDzVy20a+c/Ja6yZWsw5aX6dIZ5jdFpIEE3yOVuQGzuK5
WIEg8sezh/jraThuaidnZgV4FLxVh224v80LxrQhMeKW36EYuAedimX/KEHswDBe4TJx3Bb63WqZ
IxWYHRo7SMZtdksBlhgWJ/6mU9gW5yqTzRgUuIqAwlZHviwCIiJ/i1dscokmYngx7KufWKFPUmaC
htafq+pLswo+mKJDqfXIXNiDaoVRLGBPcXol0Ju5b+0np7LH9GG7+7rJbGJCOCKsKFxWkXQMouv0
p98LRU+1vkLwoQFgjkAH2zVHw0MUegQWZluUV4PPnBROzIinFxrcP7yx8BBHDFB0YSZDClD0giYA
Ke4HLAGFMrhyRMe7hkSJ3i8tcuhyKOEuFwK6tDcRZ7bRf3ecmPCKWmsXqhJehDZte9tvkhBHP8LP
IQLbtzGUAudyY4cCuKdMBqKSh0ObUovj4aGPUGKOSnnSdClrRZiXXRvXqx4Lest5xheSVKi7oKdi
35PjG8leFcIxholZvYwSQCWxPz3M2jDvXgm6No+Vrc5lp1tTW8CX0R3yKbu2lapKXTsBUMc9Ml/X
xJyj/1i6eL56Sf4GYro/3vTQ3uCltp8IhhYQB6YdUmDjoyhiA9KY0Q+PNTXKH+2q20vs6cnGrnZs
8vA4qtZn+4+K5XiE1hSA2p3L8YW4JkcvyJ1yh1ZqdM265AUeg4Dsm7Ctb7qs6/y7aykyqvuKbAmw
7RrmbSnT8+CsAYWL64KA7+kq7HzwB6NsssE0c6ua7Qtn/HFBK2mrhnnC/IR/0OPow2y4OgHa5bFb
kQV8qKcbI8bocJJ3RV/PWwdJc5Vwa3KT9IMobPSki8CiacSp0aC8PWYxHqGORt37sp3YgAi/5SoK
jCtRXTZiHnchd3zPSCK0f27nsHaVs6Fxakq9KM6GxrBZ1IT4g3aPcU5uK2Yp2T9rtx22yv9b75XN
b4s2ZZMgJ0klbIuiY2DTZYCfcVmD4I2e/oNdp0zYMyYMp3tSF1im2NvPQQYjrZZobFSar/LPWnb4
+g1lc2ctInLr8v6l4y7j7+xmwlEIcl6HVB5yh38i+iTcVOvTprY8QYBvHy5q7oWhgjxt5mtAPovK
BpX+Edh7gXCUA0mZW85AA1jrvMHEYX3x2oo/ZsKjTjRh04yMyQT5mSWSJc8mG5v96JyVPxbZaGds
zsGtoMgsTmHg3M5HCAQ81DF2WdKpMgxvrjAh1bkEC4sSFTjiU1HXAIMQ4QQRDcpux7bh7stNzgfE
5jvFci39axkJf7pGApR02bOyhNIfbIyNaZBCNgbBplGj8JcBWuNtnw6LJ63oXXScAOBRk1Arm6a0
pbjG4MKqKAV6vm0Xbg+IiVMqzszGRPl1vVS8XgxLS5uNlPgPq96xkfqbR4dE9qAR9syuJwgr2z45
J3t6agkjy6rl+dkZPHVyjCmNzyv0ZQ1TUq8fVoJKc8dnU5g7j7YpNFo207SsVrlpo56IPhRL990t
fxnfJ63QvMtnR/wtFymheqW8TrMZt0VfFebSL+SHzaf4kr4030qBHMzWiHijL1kHGqwrJ/pBi0mF
GUUHSLcGxz36wsAiypQwrfG4/fBpqEbDjrIopbw4/2vh8hss+G9jqXgkvvg+Wc9K6DS1IzYtX6LO
howBV9GRKMslzQLETyGdte5WO/O4cpnyixLztdZ++vgfvD5vgTm/uO3K+VbStiuex+0iFQXDxi0v
s3hsADQVwsZq7/tMwE4Z3OAJZ4efpy8k2rB0qHC4uWWp+hJc//QJI6s2A9rdTK1fKpZj/mwhLwto
cvfavEr3GLw9/wMqmjhiAaOB5YSr2BSmg/jXbVQXHiU7IZ4HlPW7dbE7cmlOmheNbjfHg3fUi0CB
Hlnz1Grs0+YFc50XypFkyUWSk5+Hd7uhq4ytAMPbc6+dch5+md5YTuA9YoxZZVlHCtoLe1zReMUZ
wMLJAB/dt7NRW1EkS3hoqZJjinXK+L8N4h5/VP48hlriAoyX+/Fl4lpJyCUyxO8Wqvqu9Mu6mx6O
Myugu4DI+2Owaxx8aAsvLJ5Cf0iEzuUKHZTu8vIB9DPf+GYXMHFCTe3BpBDSm+4UUspexktDyQ5T
tM2D1voRCnTHCkiei+xJhjywrHHTOIVkmtDFoiZqHqmI+Uvv3NFVN0pORKTC3BbnhMim/JUpX4Na
ebOOKPWnzW9tV00dni0vfhv40Wp1U38/4Lj6xJb/f0Ebn8XymeYBI+rT7u5HGLEqwPkEcBD+TSTu
PE6FCgr13/N7ORgjukXj0zw5vtuKIB40pJ/iPyGbSFC4kt7tJ+FgsCT0+KU3X3kAVjfTuq8dsJ1B
xNFnzhDaokKhk3kio9ffXrQtnLn3yZBf4Xheki23705m+NXiaaCCrPR0jS55OWd+Ki9eumKxXHLR
tzsYWY5Q1hrr3FoUFaOLYCBxmFS/YfHe4KNHoC/PSm+x9sF0ZkdN0S3jbB0vT9sjKujQBD+bAntQ
wgupUOkIGMoCoKu48EVjpelT8FrE+PMsrP5fNYZmyGm7d3v5tqZrkIA/Z0lpScnZIV/CY1RUt4cm
htalyMJLKF/mWLqLAHZ0sgifcVgjSrg3Pi5580Z+tPzJWdkTIeWrNBIPOicX3ToYe0ZoVE84SEQY
DpILCcQlU0clSJe2RvNrAeG0jlH73l1ibewYrlV9ZJgi6MiB/+TKkbHBvplSnsrbAZ5W5wSuyIcq
Nre8j2aFOigY//aMvSrOlcHpYRGyU4Q5paKRKFj3u/Yzy34XTFz0ByoNoB7PL6/gtGCBdcyIU8Pt
adNujNze7TGGImIrG4Eprzipz43ys9ZHfsqxBmHABuMd5cQKr1jAkm6ayFSU2EXKZmKllfieYa1X
oCPIWcUR2XjvCqfvLduXo79RS5DY2UavDInyyA1Vow9TGzZDA8JfjhkDcKwM9LLIbBmRhhn98Pw4
J3ql941kbqjNemb2lEcM2SBjskBr8JoRhVk53gr69qyDE/ey3rHEdillK8Wwnphqo5DM8GBxlS49
ahT93e5nTxP4c764bqY7ODuCn5g3GAC8WrL95LaqswHzfJ7vH+m8kJSuJoEqawQUFUV6B8EhbctC
wrhmyP4s25RxX80c9AIC/5U6QJz4OUWZotIRwO4qTfce3FWXDj4bFSuSGWAdhtNVOQvnY4tjrhaY
pdLOkve4BRRTiDc/A6jtRkRARSJpgYKSDAW87U4aC8CutLAtT9qTWfVqM5gusPis5HHU1Mj+1NC1
D+QgiiGYRZcVkPgTshvVdT45ArTdgm2bKWu9bW6+N3O2mep4q0AT4YHYBsVHr8+GXRnu3oB2OAUe
HbgUlnMEbHBWjPWjOsuvNWn9nSnc0GTh7kok0a35oYxyc/dsy2FWBl0OamRe5F9Yu1bkLqSQcprf
3DTWvPFobBhzSTbuFwLw5/VLbRZEbV+dAkRaNG7yTGcJGLM5w0oQWa5FhllNW/aqOpc+MJfxIVaO
HGCmSDkbp37XkoLJTp8xWfuLmblYZhdvUsE73PyuLQqxtlDOC/4srHLoe0lip3Iw8udmWM9DNTJj
r1Lla4/NovxFA3r3CdTV5+bjcZnJTx1LcoNNEJSNPmsXNUNAxcFZJfxzffKiehAa2JZ5wtFNXhu4
0kqLsXt1wb9+KKeSYmRWhZsbFfonherqzLiaHlEBfkQwY6kgbXatoiW328zkqqB87q3qmreRhs2d
h557r8Gz8xwffXTg3baSMoyH292z/41aPb+SB8DMm81GorpUhGQMBQoffxaIkwO4qZivUK1z5km5
2+1DQWVpUHWGpcXA90uJAkg8d19YJ+23pzcuWexCXWyUIZ3yqAirb8IyDM5aJo7/FRIAAWi34lIv
c+M2akbvncC/TgaE2UYgsIHmYtW9wfSVT6bd1qn4PRG77PLsNuc3lDU/yO8JbqeOzCzJGg+TbGOp
O+4CxFZpfTAqD2C6HLUtE6WuIQFezJ48z6H4zbl5GVZIzy8IeJW+X2RoGy1Ozyilb8oGqtVXF5yP
yA69TW+g17htvMv2fywb8kiTzjl4jg17/kkipzG+PMtE8AB2yM9AntDyPn8ETuEqfT5sDXEb00kV
/5Jvb7lnsRAepqxT+D+MKXfiMc/NSi1hWr1fmPz4hY6MtrzkXpQpqUPqClG9y+ad44BvjUDBZ2WK
PTx5gW2DXmSNHQkm8+Evq2EPLEHp+oU4iI3SWWo0lmfUndqgaIAm5Z2Jl03EpY57JJbaXAkIYBF8
xCer8cdyt7172Wb8G38Si4vIdUGOD5IQRChpqMeJsoRwgZMm9dZiOGfFzjGt+eOQvrNqAJnB9q+d
r2uRTzPkKbrRgVn7qCG5Jue06X+sx2YXGUzuf2dyKyS86mSCf5DdFsCbzgus5kqUiGzBLUMoIynq
yXqhpbt+yZouO+rAFkDTXqav63GsGgr1EMwbFlm964onAF6fg9xgsscV8yPMx6uIZJ+BEivGjxdj
Ru+Gq0ZOX2EpQqj7qY5Gwt3eQ7JqRr8u99y8hCj2V/sDJkB+69R5xzWpyWVAcR3deZ3YchCgUy6P
LANMe6DZyG81FUFHSDZMVSWlUMmwspn9MlmLlN23IzdbjcEyXbL6ZmtE5wJz6cHyXi99XT1AFYL9
UQhQREpGl/nhMQ+nJFC4xd5aSh3ExGLvHCmi1MptsGVZ9FpAnpDnWu3eBNgm/MAu2o4LgSXPAtmJ
SyfcFsluNE1yV8AO5LlPTb9gOfBHBVZuUViZTB0hVmyiSfgLAq35jMoDebvkOLDbTyXZMxIJjuvh
eqp+nyGsxgNs9IPnvhZD4Zb5O/b8RcjTlla4K+roLQN38kwhhADluO9YQF5vz+TjYXfH63T6Pi03
MMBqjjUGHlA8W5dqMs9nsPrbexBi2UCofngTStQrmxWJ86b3thPqbsWOK27eHv2C3aCFJgTMNC2k
p8e2ybSsJLm0a8/jBr3Vd15InAHXaoksw7S3SkTQfaZDfsNgfumM3oHQgdvgVxooi7u31UI0BXQX
K6aNSTyTZbf6UVrAzqcD2CWtXTAraNYaGdlDbY/xb71DVot6zHYo8+wy4BZH7qjLXqhBRCnBmaZN
kZDnVzW48TooYbyC5kVo7T3LxBchzvJSr1gOm+yCy/6U18nsBH+Z3pX4FRoTRHQy0fc6j7Z15vd3
JUy1vCCNoLXqVLIj02tTUX3N2G70+YYsQU1tE4303JcIJEB123gu9Ov58DbqxaMAwRfgukrN7Smh
Dt7qtPLEJAp/9vhUr7Is2oyIJzUeD67hpcfATtx2HsLc3w2e9GWYy98Q8Rk4e0CoqIlFP42UExC7
gjU2kRppTC1RyqpmXS/MS+SMThFRtghUdALC2erc9iHJCKRcRM4TJti9Sjq6EtIVO0ZjY/PSj5YN
NOzDmyIReCgH7ZT748pMen+c/uAg/SFk/XsiI/y1rBup8kdnXet7ABwuRxEYM7rhuja91sWh8nu7
8cBNNhBf+hc1UxtACDVPkfOkxIWYzjO5B/cURpRqjlAMWlrG+kPnD9VT7bKWFSLqgcemNRpNJ2V6
o1m5eAUTGUzNo3irP7q/4wg4YD3tYZG1Msj5MyhMTRKEq195cB3ODF5JlxZIgQIkdNz0Tc3NHw3/
jwqVEWv1ndX69CGcbOkT2F0DjP8b6C5jM656RAwx9HdLQKOQH0hAzgP3GdYDy2JEt+yQD4ju1KcP
CzumY009HdxtoiEpvceaah57DnUJdHHfCcCI+4pi+mUc258Ik6E9ivgWHQcGmEZmFqNDth11Iszl
rzrcRHVWLXD4KiQqIvWyE4olOL4BACICO5/qPF+9m2Klfkm/kMLMHgbwHLfXch84uSPUZ47Eii30
gLee7utW4gkGeWneMx9wwm1gwlEVcL9DyoYdeFSn91Fi2Sc/i09qPCGn2vkBlkr97pG2MGTn4hsu
A2jOcHSZeWBFK+LyaQ7J+TAxwiZ2jWaxygLbZtYuoHhWRuMhmNLC1jVLPRaLNdZI2BLdFrc8NHVz
EGV0pMz3wL9uyiiubyQCySGR3J0ohlV0+FrcFNFx9GJWVDPRA7TJ/OnpBVDtz1T61Xo9qu4TWgr/
c0zcQHq6Zrdls5xvIbAxhd4BUHUdXaXzDMFuUqthy3nSNZirV2Y+uMfsOR46vEIMtg79aILSZd38
8DhniE/I0p7PK75wmpLz5/xzBFY4sO/oKUK+vfAFxa6d81RPHCjKempfE5PJzBFZZ0Jbv6FfWDhf
E8Ul++bA76CxXvRgNfv98Gf8Wl3j8fABp5g9j61pQvi5MLkxWi1ZUZQrcigxtyQlrpo2WDIocjE6
trkXe8sW2uP3Rl+zVYLgRZfXo/J+qf0vfUyWsAimF5aaiIK50DJDDL8Bi7PSdbr+aNv0IS10iy1k
w64X+AA3TVuBe2RXTzU+1qnDdrxVFbMC019eGyPaGYf1fsG/hpGR2gLkaKeyZimHVBpfaflu8jGV
aUr75fVM2rSvpUkyMcryOzeCxPCem9gdRS9lSrTmI4cQU3X+Bg7iHl+8aai0r4CZf4kmkh2p+Ty6
kIX/VOpPN46UiBRhvt0GaqNQ6fM8u822aFQDkguDOtzTGf+DMxPvf2CHEl61kTNZ5A6JYH0WeWM6
u+FcOBDC9nTbVTnN/RghV2TxYuJVCMUUAarMoWaIrUxQPCyGhdM9VIUYHrZrXzmBQcjR0NoIWksu
2G7C4N4psnRuUqTamxf3fQt8KUY8ZbloBr33tzM7bnTCpXQZwrZQb5naE59bXqtwVt8ikJwZOo7s
QWHrrwYbTIJWsZFqisrIC4spTY3PW33U1WDfQfDEpyB9Zx7KbvfFS4esHcRyAfmr0CZTKPpB6iTa
tcKEr97h0yfESuZpxdq1eBVtT/WlQ9MCR16SaYP10UdM+nUVTj+DTGAAf/QK4mTAzmZhGGdSck2a
+czDJlcDZoSRJ8es7y2PtOmHs6AuZtQcWZAcHMelpMsq0JeW0h2WysLlXk3V8WRN9VM72hVspSUU
Lb6IdP4lXP0mDGDmRi0vuOlmb74lmSQC+JV6yVdR5ONmn7sLNxs/igUCorFDw/rmEtTHw/ooDcJT
X1b6zcE+a6fgCF2wwLEJYkBAsh9PkNff21Ecgrq/4VHwa33/HUm0LGnzzehU/+FvWTvlWbuFWrMF
Q3ANZadImyM7D6EZgUdtJNOTh1RcIqqQnYvFuIKi4F1uePwTHTcpzgTv5qeexCq+M8lxT/cQGK41
He603+GEB1Ng8uuV84dHrloFMx2TCJEg5CQyijULtCzxAAfgVbPk6x0aWO4licVswlaxATjEXSb4
NFDp6ID8mkE3jLAd2fE6+DJPZPdKTU4ZQId+0pOokTEq462qhMxq6ClPHxrNtb+GdMR6I6sMBzcc
0AvTP/gh1Bn0538zfF3QQI6yUGHxGL9I4HvYBmStaU3G6cyEFj69K17nHFn8UcWxZ9eU1pyFqjmL
AOz7Tq2uMscFtUKUNWrwZnemwqJlLrIrZdWl8NFsGL5Gt7Yui71H1anzNL5MAg926OHrI7oHgduU
sebtJSEI/1T72Y5k9lyMdgF/TFl9C0HyfxzN4qLtQ1j7CF40iNnOO1Z/4IknahiYVtynlRtyz6pL
73/UxkDrkYu9D8Y9E9M9SZwMUvMSxoGkU/V6cZetWIWDe8IAste6q89g4++ys7YhhaomeHNLvjiQ
bv8mlr41UZezevq/3nUCkW1o32MLPEex04yA+QkPEiGdHgxCvKr6l+OiS3PJYtR+abaJ11KZdq2w
rouw+nOsbvsQ+bfihpRcFiJEc1FeidUsIcyNlD5ymodtCXMKbN3M0DQnZj6HvOgi/RM7IeTcLn6r
XrXWl5mqb7QqPrUpjdzCcvRBJsjRVNGdeu9R9swQIRYWb4VzV9wnJ6vCcQfBtc6dzLpbDjp8BdaQ
7FJ4Wtdn7pHZx+4Er2pVSMoRTIvlWucvu4/g58sToBNf9bZUqvZhIZvxkL6NBqEm0n5+b4ANH7TB
ESVmmmolrFWDH6axXssTPttiIc5ngKcTDVD0h7nXra4PUsiwW1FKCukvK0mi8MEHJcuztOLquRNu
QPq5aDphkfmy73QSYkS013qZQxQlIft9v9Tje4xN9YmrKdlIQIOBYazvc39Cv84gUmrBWVqnp/N4
Ua8XMXt2twsTXC0lrcGG8el7a/GCSFer1cuNpA6llBte5s2nNdGC+wltXIOq2dP+DF+SDTrWvqrA
lzUF6Q09HXuZTQTTt+Df1q/D1rUU/Gal0ze2/4Zxk6KVkbhAxN1AyZSUxKD9LX/P2c7AYclv+0O7
/G9iYB7jQ3QO2R3FpQSSW3jbpcphgAaRnzq/iXCQ6SN8rrtPlmZT9kmA1I2UDVf3zNd0JowUf6V8
ysabQ4Cnf57keSy33kVtpeXKBdHS8I8ir2qhudIJjeS6OuFQXIEYQo3q4cf8LmR6tYJlUn3SWlO0
Etdq3qnPErVLGMrRMbjpuy2caJ6D0qC63UaCVGfGjVVS8Hl76Eo2TdCuhKrEJ4O1WCaFZAMQMxGB
UUp5xrxyGZeSsxo6fY1ZZNiykPnBF7UCFvs9E07gj8Bttwswpf/TaPo7YeJf6q803WaDSvEH74il
eLfg8Jhqljkd1/KJot6/MIHzZjbvwgWRpbACAAGVotsV/JY1FqpDlr6QfjeCUt1Bv6Is2VNjufaD
Mi26gzdqIyCniNdoM3ILFRzBElYz6w9UyHlLMsdHdnYBuYz/wfv4Al2eaySHVGcGaKyVF40TFClA
tASgmj8eUo2TlMBDDD6FJfU5cF+J4mVoze0naog7zumMuQhP9qvOu4Q+PmIydNoau3F/JqwVAjj7
cm0IjD8KnULxBv7Co3aejvaTyf+jIMmznHZm4XmB/soa5qVEypyviZAi329w6tvQbo9rtJPN19sn
LvWrtb26aztRaeNizJrA/TZ44imfG2/G8A8Ja6LJ+vSdP2fHHuHSBJyAC6thA1FUBkpnmjwoNfq+
Ak/+CbvsSA0It4GTgexm/EE6w1rr3hbdydrL/G180FqePAgqD6OyjFA3PtXXAKg8yssdA7LxbSyR
GbhlLhG9amVxQlUtAELitOXZuNILL9cZhXxKSxH+lgEqTT3KRFdG8xXqxf05u+YZES9NCA5c0hq/
KO0iIugr781al5+MdBbHqYvxKCt2EtBMGvT36kSKGqe8zxq3PenTrMcbEyRIQ/PqBVj+r2rdHRsc
vBJytwfMJ7FYo8wXBC9sc1L1DFs9m0zAfJU3xhpVgeimqpqO7l6BsguAXB2Ng1dosWh5RRx17j3D
ID2pQS6xlH5Z4xvT8q9bPQJkDCdEZUBnZORGZnaqdyEDfd9NPYPnbWLi8aoknJEe06yATOjQW+NZ
Fp4HXYY/Wzi+QOXuKw90nfDiw9iWHPRkHhEfzL2aJnDsYuBY7isd/Ir+2FUagRC5l/4CtGIFfVUS
5/H+WOjiSOkrRyoAaMpdsfW6Lt8nYg2QZWGXAkIb/SQQm3GE8D+AZJy5E2D/U02Par/DwJDpkLdn
VZVl3XgtF8OmvQSAkeWEp2DlgSubXA5duxJsQ/hDVcPDgk7LBMT1F+r3MgY+z9mawK0PaoaKKcqC
cWEZDX5bL9hNQHSRarAoEgWoqxDmD9OD+Jad3vtZutljmukgDrPSNGd/PsxIO65XUe2X+6Zonpfs
bB+hGme79SfDgSHpjqyCsuEtU96+j7hWhdip2PQiJVED/ORPK1D3oayF3e5dPQ/S5AvNvGhc56jm
KcEvdvximHkZHlLwdhxDqq1tB7e9Kb7g+nq7y1k9zHwuBI80hbFcz11iJcA5aTbljUc8GxxSIV/f
ofLgLAasH1brg8OQAsnx6/HwnxL90Lo28eBcJE8flB6leW4qrjrr3xsxWsozfBGgqDUJNyav2Htq
PJWUaLCN8+WasCAvxNmiKbQlFUawzRQzKH825y3NrejAKfdJ5vP7vqlqlQfOWberiBobwDz+99Pv
e32q+l6brUXFSF92j+MqfSJRLks0bA0dX0XxLUjAfNE5wfS72hdjyxfeEGRQB48WUSo8Pa0rl0do
lBS/+0iT4fZxdMuyJ/RgGnuGzk84UFmzqVhmCzIl3oab7LJn26mq/1sY2JjQNMOGl9koMCyGLHTn
J1gvj3w4E3KuuU03deeDE3XO9O5uya7D4m7bRrrUATZH7LW1X2o8HHqQIOsilkLpYEHNrj5qRW3m
W98i6Ul1tmwwSoufPimmk1uwMJwpwyqoBqiS6eQYmFVXIsw0E1i1hXQIgvqsGNGsWYEomWK8PM8S
hg8TAW+3/m/fBSv9JvxL2PNs/Vz2jtCvDoVANyuj41qfbYA2QgI3oFoycW7ZWLqyDLzmSSBKEFt6
uwBXRKBjiooZJzlz1EgKnWqvsZAc0pdWS+PVQRf9xvrtdKdpOm+Hl9zuvfcS/jPRygMYFwr+IZ+b
U7TqTumhyss7khixV6+9z7RBpKGwfA3zy4KwHtqkxeh1LmKS1Z0u5SIJAQIIjkrX/NxMCFKvL+v9
sdSm67OHPJH0FiBmn+xLCqhiZDLxrQovGgOuDRo3zB03rraNWpI/M5Mbt1p47luZ/CGHS3PAh37d
FpiY7G4NG1IVwkK9edLW7rHQoufYuNI0YUZdC+LZoLSGSTHTD4pS4lkOTLUbbWF8X6gOKzzhAxzt
cp0ZhnRyz9lf9ewJky3jsDY+J1mINPjJLB3fxUBITQfCbarFzL1u5h0xPoIW74aZgXG/d+2JhaDD
TQHBD4V2UBMhl2nrJjry+8k11nSdMje4Fta32eVB49AmlgToUHDxEZQE9YInFdjxiNBUucZ1yDtA
7XVGFJ9pVg9hmHsxj/j84ukq+QVth3ncfINtaert65RGe5rNS0mCIxMwEudfFmKB4yW3KBZI+pju
5xZN5pJajumuS68nO2qx32fvGtj6RMKZa/ulAuzLMMp4GQQ4ILYVETirLHOEZTZNDOHxMkVwDjBU
0p2+vdjqt8nLCgww73Ovutuht3NJjI9XOpUMbiEFDDwGxwEhcxQE9Bay1VMJYp4EAg0tOzEDxppu
c+bjb9vJ13lOZNkP4NJsjKvvMg+THSQXmtJCleIBfDOfpQ2N27qOtuIlX5IlkL79HScbqFiSGuaE
JLV4/KxgSIeyGYLUbyu/FA8siGfyh7MqWfq2S1rcO++nTzZEDAhXHR3KFC8hC6ZVzbHjECbU4GnT
aOIGdKLvqMiOSrtqCTVyV8r5kcEBTUYWzaP6ZnH1UFJJPWWlckEHH4eYTDw3naCYYINK87xHYyFU
RPZSP2/FOWNO7SUs+klfV3PZSYdnxTL5TQf8Oc2qesEn0mjKaIy5RWZOnYg+tf7F72y7FIKRulqA
oxppydtSR1cS/RU/qPQVwKSagzGfbDn0p/yt57+364mK3epsLyGmu1F9f+yc2qyDxfj0rko37Zbd
M9h/NRFTYNE+IaCG4y7nqiVIS4x0pBPe7JXSiG1t0uR+bX5U3mW5tTfKoJLsylkM03OIxInDanA0
SNZR9Qe79rGQyzxBj1oFZdbjPJvke6MOLRXdGM813zBwCHnnVFLTEMxSe0raGKVuwE4x1lQMmUB1
7GIoZWCza3xRyQ5dC4vBtOHVYaTyb5XWZusL9O/S4yoRtGoYFe807kkr4B844wuj3UdBk+nAL5LG
hl7gBy9d0mgDypwQKnwliDmBAWWsjP60KJBWcJsgJ/QWujZ+84L4+FDMHX6yOjQ86J/+fenW2t+a
qVp+IwCTmWUO/qg/dVYCkgBrXo3E2oty9xp9pSrf2EY4MsZITK1cb/LpLzKZVbF9U8PR6jotEJS1
LaakZs6KDD4QG5o4+tFHN+wpnm14cCFND3j7nJEeyMYRmoXdistMjGtFXdbTj06htT0OdhBstCCV
43sNW5XZKBfakpEktOCNqHY/HZY1tLZlkKSgofuiAflqegbEJlGqTdLYuWzvLQ+KMwMvrR78T7wH
LSiGfSszYx/RJdc0842hmh44s3L/XkbXnuYviv6Rj6oxvppRo3gkbLGhI3amCbg/viHjtCywioIc
BxH6pK8V+G1KJakDndOOpvJ10JaIWCyRrmepqkj2rURaghHaRmVHuPQ4uLf4IvaDUCq+SWd+lVWa
Wtj6Adbre2zNKMchbz9WNR36fcJNbKkuqWrb0zzU+Q0JQ51YaurJQpok+q9i6xph2hfIyqMJ6EAl
JYwTs1gGZhwZJVZXjSxHfzV5HgKhK07YG0AS7vdANPfj7N93rVIC7jiA82kEJRuYKzEporalJ6Ag
nDwVtcMYB3mJPOyNaWSFS2ZebOmIYr3KwhGf2MKYkP9K1xGZuVVHsYKbF4a7K6qnybnlyFKvRHYW
ch9f6iE+C5OVuXyutEXB4L8TRVRZE9AKhZz3TCYpgf6TRJ4nbL6iqTeghfNGDtEq+vNrc3K3Inp4
hp/rnX4hsbL7PwPUS0MWve2hvRdY9DBi8os0/hXUJDz7b1b10/bCsS4fczvJYZwCb44hwXhPleEb
OphEMKHC1Z0uG54gp6v7D8Oq46c3Xq8+lklV/rFPJNuHguvP68+0IfpBVVMGTmHyna5XLG+1yQ9N
sVbEJH0/aa1ILeJc3RqsXiaj8c9L9gJCkf2dJWbxk8cTNSJpLJ3gt+SCbNKo+2RtadCgYbuDsKZr
P+0ugv5VadyOyOBNxC+iwXGwMFBFHzOphlyChqJJ5ALqLBUItROY6dwgeB3LVg8cMIW7P/WpbsoH
inO4h7GTKeTL3S7e8Q41E2CeFnTrk1tSNMzWnHqdQBk4OTXvzSrIkZLCeQ+VmWbfH/2eTfN46/F0
iuLlZsoncO3PEy6+HGOfSoAYmcxE4F2+YinWC9m7JLHURB+Pxz2nlmGQTPcFP+Rd1BklhHR2JLUR
sWHy+CN+7PWV4HkOCOkLJI3rAZcbu2MAKL61x/JQrA+tYOTk/lhtylUo0wyJJ6gRK03+lT1gZMPd
Rum9Rpuw7xggrKvuJJD5OB8eF89V51oDuAhWw0UDd3mZdW/dFUXjzkxTFyHQIEH819Tn4XWtaXtM
MZzX4mI+ijUM7anyCv0WNztNMpmhju5vv7Jf9nGwYChAd2OULfB1LnaI07ejnjZ9QjdN7yt/PgtM
suwTXGgCr7NNnopwtfL07+VFHDMn7MHSfs1nlkwJi2KsnRToKqHV7+GFsoMHm502BrG1nOWbzl1k
oEwHJSVVE9MXysE5ywLs60TPUKoGd3NXjk2niKvwRiQDRaCl+bbHGLcZmTWK4SITypYIPyrDfkcu
0CVXWkbpLM+I76YBzZIPBF9WPyV34RQeEw2NGYo6va6YM+LJLW8K6eYspeQ8qV/7Um2THAg23kYK
vZ+o5PHuVl7JrXKLlzg1Msl4oZj5zElzCM4+W7254CPVC2qxLUpAb/fmL2tqiVNe7gQ/ZoV0YyVe
qg/HahN5ovaNJJ08NbOQzjwG5W96/aSTQvKJLIIUDyGkz+1lIe3t7NNykQP5RqhihMqHhpV+YcFU
aBmNIIaTb3gtF24UxIApCZttkwgSngltAO++KqnXB/Q/SKLn9Hm2FiwDRKjNJoVQy8XVBTqxyZRe
snitEos7tGZ4LPqRR+5aKFuh6JnA+6cl2Vjnf4ymM39KuJhRGltO0nZCz98GcPPlhuEBL/oV0nfx
3WL95HvjELLwI9fT7ymuUhKLXZXUcDtFhVGVk/0FbjqmnjF/9b5qU7mCf58VDOxz9onJSsyjckXU
lTmXAbBnlS4eYnLe+zm1ifhcaM9dEvbUQy7H0NDt+RqID+2RzcyJuGtp8lD9Yh3vUHa0DHAAwjf1
/6ntgYTIHf62u+f/l74YHtar+1ohebSOojSOXI945jEeYii67MYTUwm09nH/Rp6B2NMeyLju1mRN
YSpaNe4AzN0GD/04CeoD+iIYHhkeCyWTh7xlJVHL23d67PjcwsuCNwnvBcZB5dHdI9GtDCFyr03+
z8qydhXaxu5AaDEa10KaOTEyt2ikrKfD/bC6CR9Jxag73/LDffNVBtEFQo/x2qtBliJQY7we0uuu
8w6sugJkZlgyKdHK7lkJavFGS5pDGwTRtC/MppMR6nrkqKC+lUlwEZMUTKSYKv8+irPs07IXUGLI
JmqWe1yjPrUHmMW05WmxZJmI/c1xsGJL3qHhFFMDZVT1sZPJxI5bKqn06JIrkMIdWEgofERK5X8a
Ec9gAn0bvBN8kS6sjVeYKc6VtHgkRFXwEQ7Rj1B7NxBav5Q5/MpxwB+i5tV4yjojMTnUnekcFDDJ
BhYmZq5m2xjeOOvxEY+MzakPyalo43vVqcKaGhf+Ny1teM9Fh9L4eG50fhdlhZ/dn+5CxF+ObzjM
IhnuuVfYKZ367IJ4QmeUCyaDVvC01Bycw1JtQEHv64TXeOQCyRFSRmltvmFOiN6luLsPnZPwO8do
qXV0XjwCM9sEXU3mz4q8kH6IVHS3xT47az0uztEG01RifTWpXQaF4GhkEo/csC9x1oTPJ/BkNsw1
6t2WnKLlL4j3mYpjMYW/9aufmXezZDmxNd8cFsdT6lx0JkSrIfHL+VLDUehNwM433NZAmwsmjM5T
9Iw/JNmHGgKiILplEgaXL54ACiwrG1WioeukY6CGMon6Z2hyodBCF3L1SRPz45e3kfV8tgNe/bXt
hwJR86BPUojfkWnhW4d3nr5eFizzGUesLuXDuXk8YmBaPo9CTd2jUUDHi5qiA91Hl8voB2gp4ACD
J6d8C9VeVkcCEE0CLRztw1VplrUcF8RCjehvSINSTzpa/6yp64YLfLYYnFGLsDy9cvlZF+INNzCC
D2ylLCafrwXtEd2CcVNBuWkYXENzJ2ft/ABfgTzfom22/zxp8PpBxBDTXwAGtWZmCrbOtJ7IboAg
Ias4KTwyFl/REDcC/DpbUWhQraxp1JxrbNi9MDgpvp9vV5yDuuMQh4L5Py2cJX3fzhS8YMOk8YP0
xOEcXTDMRfFWx+3WdX4sY1cGusjISS+cB2jX/2g4bh71XGjqP7zpQw6M2oWx9nj8q8ZF7tIqk6sr
QWfnK5qMF1wEpA81bG5rfRsnY8qtqKZNPvynz4dB0cOVRbG/tbdy4GJzFmivEFsg3BiraZho8LaN
eFkbT/q14jcVBDeMEau+CqCOXYAS0LLc2GOLfMHaZYQcMl+gBmI1o90Hav7YjYF/Gg5wpqKd3mNO
UCNA9igiVkrju+UvewUy7o0KpuAIrCvzNSDMDE/k/Seh1LlA/wGSH21Om5af9ZWWixRHOMF+zP2M
SdCTrUn5jCt6EFFVjObaNTGtcyJWo8djjUHHRa3wwz2COHFKbOqMMmfKh7/KQd45InH4195ieRok
wqRyMdiGVL1y6FGSgMBsTxJbnlCSaPRZFjh0jbzF/3njkDmFXkQadljkbTcOYhYaFzbLgeqsFIY8
cOcA4cjt00ZlOQ8vjqvexODOrJAPaYxrv8DEXrEToYKlNfHrDbWk4Z8a/SBYuQ3+Wo+w+bLHJIuV
QKbL4zy83HNEZSgA7NfehS920iaA6Tvhg9eW9kbBOetXgSoRFuFE6Orl1ucLZKfzZ5s+XJUHVBrS
mlpGLG62bvwb0ShoRwPydlFreepnhoQCWn6AAxb82FrgGZwzUYpcjHl5ycE2ogcoO716doKhqozY
eT7dCY4Q0U5AdFdZvud/ur6lIw5djVhJadFBDPg1ANWWUkMqS5SfjFgfN9W/mp3197Mf8lwnn/F8
JpNsB00xKScnDG3WRkAd2k66rC7MdQ1+JtLFrjcc55ltQla0QF3B5zKARVaZbxl/sANWSoVkKOFm
FBhQoxmylNXrrY5EjYzej9d8zvZUSZnWmDRqTPEDDCXqkoRpmVc1gx/pDgeBsnAu7K4Zd4qRLTcf
mTb3gfBhoA9T7OvSkOpvUe5fILH78PVOSTt2WFPfvMGmtzb3YVWjrfM2QMbZ35BVWV5mSRHabN9p
c61di5pkmqu0DcxJIS4zBW1SmtBdCZcvMzvaWFyZyQ7SmQdySHlxhQ6RKTPnsEh4apay0OnqjjD2
YNCOsqbVPTw+DA22qogiQImpt7HSUx6jxGkD40v7qsd8cF4vS8thJ+NWwrBImNPbIH/ODs80z5Tv
hBeHRb21jUnzVdxFQmen53Tom1k7kgQDR/rEloJ+YW08sy7HFe3o75I+cPkPvKOgCYpiq+5yNljy
l6Wb1KrAf7UxbsGEENJBtVQUTjAs/2tbbw9AVRzzs7TIopzNCrMiGEF46V5lrFCRo0ilBbRFlv9u
ThonnA22/ldrnNiSnBR2qq5idrKBIJl8AFGJeM+9TMOYb9E/KM5wgcg4DWJzGW4GkA47j+QSKDit
2VxpWQL6F8NC+ZzEhclyBjg3Op33nxCcI0Wn5kareWJpPSznOXQZrzSYicn8568b0zkBORtKFLfs
/Hnjq+U/H6lu/8n6q1Zi2Ge/WQUCAhR4q5peUZk+df+pbt8VIiUEudWVoF4KeCvkuxaTRh59fCWR
tjE+BceadVwacUgMiwXEEbL/AZru3dp42DpmxBwL+G341BZiSCcQB+6gHgosFeUsjWyAmvoLPExl
3yGS2syt+FoTC2478OtXnW7kvfRXn/hWoNTub4Mr+WyGz+4/znRebXowezmGNNjKIdf6LGtkC7c5
tQ/aOHXdqqLItQO3xI/FM+dy82UwzelSevqFGxFd9xtOrJjwQcmgjDMXj7bO46s5g+/YwZJLoqvt
MXPl7EFrxl+lsVnOCVu0cN0OdPAKjcv07r9mzIrbTu/cVcXOgPIws3YVfq8mnPc4HSo8zit99qWO
Z4xW/JQbrFFNMqMbpuGdfxfFISMg/luLO+yUmIbkOKg2T42eZan2glNYkBTUHXncXGidikonYuGo
M49+QSo1AdxVpAkmQCfb2G419emLMrempjim1iY0DGkPccoT+4KN6qit6xZjeEYE8Od9RvALcJ5w
FikQtPFufNhD4gg38e+y2Z1amh8kJZojpIDW08tzT7MVGfleXDiS7LR9UgLMfFeKVO5MJgLTZ8y9
G1Q7MdHWWcDuMVCRyRqBiH/LCSMtp+p2HXEeHq+y49lBIUVfVp8i6CusTxMe8WJb9SbmXrWAVeA8
l9n8QNMYyDbcgUbMT+mAYw7QDt8viBNSoveQtcLTHkE69ZLLCHakmBODns2KQj5mMsBZPa5K5IiU
hgkTw+ac0/CXa8FlTLihBro7oXyjeqWQJUztDX8FncXtjDFTs8UG4rgtO5bJ9NiZk05EG4lYW2j8
BTd9CXzlS1aE/aiRbPo2wMlmFzQuv35yREZYwwyg6FEDUjRraW5cyBTFmSDvhrSav+RK1yHD5DYI
5I/smTNkaOG9OhCU3e9JXQcSN+uho+cgGMFhzUiTiJFGR0KmUoZ0IsKMTdiNpaU8BIiEgU64ZIcW
Bp0ZAGbOTUiJgF1gkcpkkRwlCevLo8oFOb9CZD696ZTdi6k3wf6ldvap6sf/ls1HSFnmAvZtqqWJ
Dj87hOm3xj+8BrwatBES5zQOKAHUQm+HSTTtpeJJeN4PRYxTPfvFQtnvJRT2dstRvLtq5DOolx13
qgBjbFfGBUSplMdFg54941U8QJx1enV5NI55KqeQQH1GBBxQ2A5vSXzRf0jWG4rg2keQFxdE9TwR
YnZTuxiTj8I4AUIwP8iA8i0wQVh8X0ECJbTMQ4k5/qci05feBx/B+QwLX+uo6e/2Xk4ZtndoFAkH
TX+SHkcp8ykyBku9F3uQYyM/ipsHnHjFQ10O5kmRt0BbJYYTOOtrG2qYh8xSn0zUIjL/r5qoW3B+
VzVo7C3dZEY63Yz1VyKJR1TvLQCD3GmM/k2reKJmwQA8bOKnn1Y2s6+wNxqtTsOTeOlbV2Ct3+oo
aFSxFcRgIP/4cf60EckY1ExX9/ulUFrApnmHCOcSQoq9QwJk2/I38Lm0DY5jROoJLi4LGLFNcB7B
coQqH/fLBYKUvaZqwFJ5NLzgreUFnNZxA7bQXIlyqcDbKWBaUORX3APiaiMLvwwYhRZQn7+iuQv0
OTVxDcyJyxgEKJxKOeU6Wijr734qb+qNHfhw2nxfwfuSHRDXVNaz2HiHqdxtid0e7z0M1w3nXXOF
0XLi3/MjggkCE5bY49l17AHrpikwXrlu+FPMcNmUcHRPx6F+ww8jkBurL25GRr3sD6DmAT60Q7fM
tO4O7Wxg03DVIsaxdB1y/JRJ9ZAOwd3xtlOEGDkVRtsztmJVVYD0Ayv1mound3fmyrxbCMeuMBU5
Gz4jL/6jGU50Y6Yg5yoptM8o8TBxeg+MGHj5teH1653Zyf12IVMwsiNgYWy9EYipifZWB06HCFeS
PozdyLlP2I6rnU6QY8b4T0JH5N4UPjnP+wQ3Bjzja43OPqPmtGeBd4qnPvM2w6td6qcZXZH64rC7
h4oE+qMksInezdiVwILFXad8T145koXRFd2cwOP6Xd7RhXvA3/bw2lL5guUcn49GyydmHDklIimc
7np+PAm5t7e9zMdGIGJNuJM+KT8KTQjszRb20mNlMzR1DuWfF99vxhw3ftKB0vsXeanxuDQcYvAD
7TJoqO6maWQIBOkRqMhnDyM8PBv1iLCkkBiLb89wy79AfB+KQIOWuSwmVHPiws2dDo+UOPFr8nhU
fT5cO5mxdiPq2qkKSc9obnb4LIKqX/5lJWcQ5cvLIZsnTyDqqwO0zhVrwciuEg6z47alM6c6wW+D
6pinZSFRuaEDaSZH68iTIGtkTH3CNkrqht/NXwxUsFFLViU/9rgPYw+LdW0dpTH+lnq4GAGDbFJt
+072udnDGRrp839Uj2f7F+pa4JCNBEx6fSmRbjlXiXojXewJ8LAUVH9h29yJ7qKHoEVOstCJGP+D
zsMij3YF8C3Yb3c+3DJ41WANRODytDyKbysESndQX39P8vfzh2BvCw0Ij+rawp4+akzKZxQ+fcRa
62XsfYeuKbWXC6M9ivoAFEV1GoAT+tqWk843Y5uSYvNpWBZFtNfowJRuaVz1WrcE7vvYnjMEMy4C
Y0tFQrVJ0LAoaOx3EH1WsQm4asBTB1AE/Whq7RFQmq2rOUbIUADuMH30V0SwZIJ9IfMM6XKL+m3r
uBxRwwqLr3uTWXsU9SSVe6ERpDqJlFzQNlJ6mjTTrfLQd3zT53VUnUjCnXRyN/ho5Sb3ASbdUcN2
D2ZXJzFUJ4hj3KlYC1vls0FdoDQLhKvfEnlxknkjVKiT8lizeM8fB6dY1lYrxSv5ImicreZk9i46
pPfSMhEE0Ml/3Js6Tm9k9LJnL0n+AAq0cda0zaFO/Asm6jyVFC5AWGG1V817jldEii3meQGznnzl
JIYaH2aJPokd4VonhQqcTIIdaAQ9kFiIeUzFZ+LfhUW/SLttUE6w0/inKTOrrhlT/0fHS7yhKZoF
4EYk1M9YvYGWTh2LfCJdKCLztziNv/F8SNObwgo4pWuxlkXyycVFuGeJ8p6UxmHlnnVch3VUQp+N
4mMluxqV7s6BMHw4b54/RLljHgrEKHJ4ycOFL/NmvP+HYZbFAgGMPF3XOaKAXqhX20yD9wDoviIJ
+bHyZVCtXHJlcUkDDi/YSzMhUTSFxXDep4Gxi14VQhTqgYUMYa/WJM7mJs6QTXxtMo6e7sdE9N5r
2yDzQ0ZjYvwldcCDjNpsUrp0UwqabfG3DCZHPfaM3i8woDKYCSI0d7pU6hGq2Vx/ePwT8N6jcMtZ
RmlwUDjLuKHbkfGwuyEm+fwSBrAewB22Zr7trIA1yJ7ZpBevTGyOdp5seFdLRqieE2N63pU8sueX
XpwkInxgTmb7nVPXzVCdv46PfVdm8AzL/8jAIE1U6lBOa/EOyKrvZMwbpYKWQvzkpxAUgYDJM5j0
TK00dmScnCC5dzmbe/x7J+o3lgJUcbjDFQv2+tQ1Hy/6UxwQGoGKjstiGOWzZEU+bn+51TgHGVQm
WHxEMvMWBlwrKve7JegzgGbHS3aaZaXoKInBu6udN7dxpz9g1pc0kIdsTcy/3jElTKO88ck7PaDE
4CFwhCCVilzfzJALHFKQ7doSbmu+1NlaZY70hnUyEk/Rei+KPQwV5lOH33sY65G5C1Kqg0oyq1j4
TtVgRZePPug4GnvlxNKeGGrKczI9kRMLwfHvHzGDpQswiHN5m8d6ah9pup1VXcV9XCeF3VZ9rEdf
yqGlnsO+iDVIrUq9DLS4INzGE1OnPm45QPOUELtDxR3mtBe0SFxLdmY8FzSQD6bppLApA7/ccknD
G8f1tJSSAa1CwfCFc46nud5hgjMikbd1ktGTU0EEN/tJ+hTLPPamHkrW4yvMNtQdP9agTVMk8DI+
xRIEkCKEnZ/81dWHcRX6EUUD4tA5nHcjWUNP0pCyrOHREl5PhYUO1AI8rMCDNWqD3gjXhmfUmYfr
RPNM6SwTl4DSsvSTeA9NSy1IspG9/1FRnHmpG5zZVGmdfz1bg9E00SghQZ45RSCQsXUBovEc4pxJ
iFMbJTKoSDc94IJZmVW6tdy9RnVSWVXQWeNxVQXD1bV2vcwKbm7z+dRAkZLMaMAxk2MtEb8OwkCT
PQEGFLvMOQibGNTo2qdHcTBiDv1CTJr79bq+IpSABf8QkEUPVo9cF/DLeuoVHN9snwrlEpHzMsDq
g5GsEKpkPOmkk7yzKRf3ZK5ZTQw3qoG7MdD+G4Z6RPzSYWvQye4l+2BUS4Ja4x2ZdVmMcFcVtDN1
DAI5DpsNocYQYYgnr2RUQuuUBCCGKdGgT4W/Z2Fj+Z2rUUPRexXPyvxz1lxYXbKPMneFn1Ctk82H
fU/4PXDy1/fijsrgSWYuQ0pWKqJeuKPyVYaUk49dtyFQBWVHPKKwWYTTvtjzhDQmr4HAgnlRrmWQ
kUeOrwOABqABcgMi4nW2nKUHMFH30KJIQtf2eC3nOYfuvkGx1/FIS2PA6eesA7oXTid4B5dSGez+
8Av11TaDs9iLAjFqmA3Lnv6hQzLxORd0NiOFRsweNCOBR42QTj70jRMCIRUlAxHQ1LNlvgLroPGI
6tbNq3Axx/ai+C2xLUXW7ZVCJxUdN91pemhi3HRs2VKtYJqR2TxjOfA3YFpeBc/Vsj3aCb8CcNOu
1FIzQU/7W1+ezqiob4vGSqVQCIGhp+NK4TqykrcNyKgsf/+AnxEOZRyrkkbAMtLaIzC+Q8raCKZu
/+glXSPlUGUxbHQiQhJSr/uk3SIjMYtffW2lNH/f51VF9ykUpYOaOM+EjD36uctO9WD0Mp5qbNM3
hUbY0XQLiNtOh8aJGVgKAH5ci/S7NgLtWHJwp1glWg3U618La8SkhAjYX48iobBwYd3+KsPAtXNz
WEvqXM5dBkLdhGetUDn5WENawmTKogq4nZgCueu21JCCjnhPu3Q/JiD2cjDPNgjPlWbruFSXkTIS
AAL6d3/7guDblvJuZRrctepqJdBQ8VT0F3YJ2exdEM5xhErEyWmymxQFkHLHIpj/PUwkDYvpaQyh
G9ZbKSrTNmp3RRmqY69If7RwgCkraLK4TLWuPLgJ1+B3MU/FkqDd82FG0z6BRaiid+lI5gJsr+VY
WzQgObhGVOhJ2ypvKOXzb9bwfg1ouw/uEk6FvDfmA7Qjp/xbZH4Wm9kcNCycAUC4Uasef/XxCgu1
5L6sm9Dih7ngUVrkr/z6mkU6YSGBc7M8u01/h/SeOj6hau26kTsExV4WN9MnQxxWXicTtVbgHq7k
MYeYh2TLJ789QDRYuLSZ6Az5R5/cGYBmL+D92MvjW8goC2ykIvzWesbtVlhHJKZcTBdTghfuK8iS
makfqGbpAQoNQYpESK484DZSQL1o6xB5vF7lt2Qvoyvl9sjzwTDFfTYSRv0X81UvM2NB4ch0g/cZ
k/Lkq2UiFifuxY4DTnSf48WeFJ77j56p7xmu3lJr/zbPn9QugfwaaHQYVwR3FKasx0v0a5XZ7KXb
uvYmiqCj3igejRB18q/9lm4I2Ia+xWzLKqG9NaFKLyC/5RGc1E51HOD2Dw8dEfU8ZocREqtJs4+l
8OV/wEQG8K/opxGOF8kS6Q+orDk/LuRNsWH08Fcj144IMcIH3w6BrGlVXM13j66WOkYdS5Lyv/e4
vsnhV/WBZw3YHM1iqE4SM9E/D5DUCYag5+STHnQSTRqIj37ZBhEQxKKQn+7O4Dp0Nn9FolwxPZHB
nONnOhYf9xy4cY5TiK+tL7FCVODh6qoqPPiTcRwFecn6Eg6BVk9GTSsQxN9vWhzQ3goWn8RU/imd
ctNj5Qxx8cmJTJBIYhjTdCeFVZfzl2zmiSBhCtxxopnPxbd0sJSG1dq3idXwJVje31S251aI8mak
d+tw7cAngRNLH/cn1XI97n9YAIOIycnZVSPeE/3reNH8aT+IvfXkEI/NB2XvBRDvy+d2JuQWIfK/
ZPyub8QZkth6jGe/9yWMVDDJE9QHEI18DevnOhOeToL1AeC9akmGiV+Irp/knH1V1XsOvs5Yb/Ii
k7r4TWoNqrTWDUYGAjQ/kQVQeyge7Hkus2oSNf89lP0uVNA4cVJHLJgClK7ckcZPFvKAOFZwI4Ct
E0Xg/1KDg/kWgLLyk7v3SpjlDnaFpNih/DTqE17chSCmtKUkgLQhSvrN9SmRhNTvswIFMhVe5QCS
4RMXSp5c/ByPNylTIOtEB+mioPcPWyMOrU+6YLBqPF8PJAo7gVVNXSo/H2NRys6cSsdwy0PtfhUZ
/mgqGLhURCq29pGYSPzFNtQiSpgL6q2DoSNpLJG00L366hSsQL96fKrVmtKgya1CQu4NPalTaAum
31D2IgSyjuDveMMvXx5I0nQMiyJpMPrkXvGxBaVANqM7pjRvP21x566vNqpVwOAj32J8gtSWX4aT
j5OA9BAsQYhkLVnbe5v6fUHCBNiDa+phdvpnJa7hAoIEuzQ+2t6fnjvIJUN4c65rVC5hWEkMfWa0
7OCJ+z3Xv39f1EF1CMdwLqtXcAQpv6Sin/BBOGN3xdqU4ptXo5dBVv/UpY8ltnkebQm8zgT6ragv
uy6hAnzidBU6DFSZaZct4Y9WrFpDR3Yv+UmJVPePfXyQa0dfeS8i8OMSHUpnvFwGpAtEJazRBwTj
00ofV2akncrCsz8A/rNdr/b9C4/lAjq2XbbWjIeiDizdjeyUWDPyzRNdQOFCX/c+9BOD3nY/tI4F
upmTUEh9qXIxj/ICkdGzUKqJLpP3fQZp/Shc15W8gBo8kh9bFNpDQNyqFY80oe90pAZczVMDYw+z
tgrpCiE6v1DovlsHTJ4Uvn+cDJ+9Rq3u2Y2qUiJ5AlB87L+5L7iI+zSOtRtl6SzYLBoBrHZTAARC
SWncBwJU48Gm/ePgcBSELNy6mlRtsH7uWr/uy8bc2Szmt+8UhlowIR99Toin1ZHqDIA78CTEz0Pm
JQotsH/EQLrXbVBuiBIdO+WnIIvE8nAFxPhLiuo5t5K4Wy9YoefiGSWxCKGEt0IFjQ27BAVJFbSS
1A1NrffMWY+yAbmvx2SrtcKBNLRdDEwyRENKkcSlFMrvwraCbOvHcTKlGLDxtp9kgRf8Vrdx3oG/
16ndwIJjxzdRjvOa7svqU835VN6NTqdcTND+8bzjdgesSHPhRQ89bo8G5nMBYxf543/4fHUWyKYF
6LFEFVb04l4oHkezkOuWyNDwkqsCsA1xkxRztXrm01Wu5hFuVHGTFMpS8PmgnIBGz4eIsIpfs9Gw
V6vP1fI+PO5Bafs4IsTPbNj2AxLBq2vjU1pATUjUBwEULNvuo8Hm0NX85RsmIAPsQO+asFgK0fl/
bgbIk6lyO5Eul1H/g2avltlrRZN4Xwz5VZ+hML5QGLXTmA86yl0l3irKnPaonWxVaitQ8b4/jM9F
e0lZSqFt19svHGv5xlsiunwjUMKWcJO6D4NGANoW0L3J/ZEZH/3Wc0Sv7oSE1VVosw3GP/lNtNNI
rg/A9cUKzoxE5AojceefKDFLgDCNU+lrHmEcWBWduXawtDmejyhT3YrgNl5FKAt8wSs0ggNCuJq5
ZGdUPC0nYbxl83D+uGZcls7JpGxRKqw1BKg3LgUacAgygyGcrQYWLhyQUldsjGRzUY72kIh//XiT
mi8EmCkJF/OPl0JdMO7cVQjhjGFU14IZJ6yoJlpfOpam9TP4Yru2XdR88SZbAH9hpCSfR7DJ9xPG
UUnJXG0jHl8L5C8y83fdxpP5l4k89+vObVH9sOqkDDX48Xh93BV6ptQa7LPI3EYOu6Fqc7nMb18b
ZOQSwnN5ftaf8QYG3u+RAMVbwaDJ3mAOpgE4F11hE/MpjIK+2Dj49qKM66LjYcEyqXoBheo1yQ8t
IamE0O8V2NJcq5ddsiv+t0cPoFehtBSjedMHUT81p3ZlqQLvWQmDzTWIS3nMB61JeX8FOWsXSc8R
WN6AceaBMnyErM3AC5GEWsE0YpXJBwQAOp31pfvOAu3Zlw8RC6lkj3q4OaWnuKNS5ZZkYfZAu8NB
yZ0TZ6rCJSSX5xcr3ASCo9eMAW7uclNJFPFSjrh8ni7GUGdEAz6EQH19HM93HeKEGTWcjZjtX1Sp
ZLo2GSfV9/uYS2pqeaMv1JpSu9CpKkGSJF/rZOV0dtfw5tV27hhufkyTPHJRzaEe5TVt3zOS7/Au
uaXf+xsvGFEBQHRRFq7X9GJOcJyJ+DCKcrGgh9j5da+NIoBWUpluyp3wwh+9GDBxKVxd5XkPG1Ki
Mnj4StvcJG5iEEkMiackC2RXz/2ue0BUDw4kTzEaL3/1nIFiJL+Uz2IHZ9Wr95Eku9MswG0vTND+
S58kmBvlauAcAVXf51bOJDlXT3ttQWqRvAvYkWY5rx2hhWnR17T77HZxMsMPepD8Eslsa42k2SYV
WU+NMI5fH6ejMy+ju9NxVbrlTsLK6+C/dFb26chcNkYQIEjEFMkMQJl37Bt7+HjM1AVtAUTS01je
Vs/Oi7hp4LmawS3RoM0PQZ+AdlftcaC+KYLXE8SrtsFu6PSAH3xBDTbLG8aTS8BI7RB8d7mOvyOb
s00WipctTt4tuVicAchZoKbWWRxN8dJQH+IaMn69hZZMybBS0QgqUKS3+UTvu+aqqb6hPfsUy9h4
cPwNR6jg18S84RUaPgN/lSNvI5iqs/BdCkp8gGpM6MxVI7VgYJiCTwyGZLeDPXMu/AfwM7qxztsE
iYwP6+Ioh1cBtbF7vJhZB5KrTd38ofs7m68ISYh8kI/eDbENcLt2XCI9PpQMu4SZtj9ULVDvDQQD
iY7lk8w7Rtz0k24nP7uPfZ78w5kBFPR6f1YEEiudVsujsuhH1WIV80vAQH5qWwbzvLR28EWh821F
bDFA4ErpzcGK8sbzhFN/yna8XhWGCq6XiNYh2iyX3lmuPL5HpCi8Y2hXtKdSWgFFi7c7PZuOeRic
U/iHP1qEo5aJprZoBZkqJv+ezPORDHHaJvmParaFLB5/mwDwxCa2EqfdoerK5wbPEs4TNGkylSEM
q54HphmQZrlWQfNbmVDRnD5TKFX5OslrOiELZ4XYGKZOm9m7BEniSlervuBezRpIiUphvPGsM9Yg
WGdiDPo+AiRh7snAmT6zzCi9kJs7bVf3c1EPCR5N5IIfUgygBkA0uAHI+OGLyEIrunz1krEevFg9
yQc8oZndB0AHetXfr1e9GztQMNb3Mw2IhxniZoRjxTWod4pQjtLdmSWGs29aI1KmpszjAxX099QK
Px9K8UZGDkZzKzUTURscgc3D8wujyJ0DOipSCRS2bJ/aRkROD9yYUu07LbEHirdupQ0CbiSWCtYP
cbr+PyfQ4grnkNb0WnvJrqp4K24+F67XUZldwkNcl3qfJZ7WfszryMsCxET1roLNgf2HkRE6T9e4
rCwwUzYORKJEHMwxKNXjuN8DndCFnAJOhvgWuXdVqTayFwDlbugZVybbvzqqV6IarmcyDKfkJSbc
C4WbvBh4mLQRfcPjBhJw8MzZZym0abL+XfYyRohKiXvXQ6dyH1bO38PyOYVo1KIQBXiDNh/Kxn0m
E07ksOZQLWWsRRXa8+jc2JJUcYg6sXhuU6RswbyMo+TZ9Wjo0PJtupGQPnZPd+eJfMRdg3EyYLF1
GHYWMeQnR53TSDAOWTvFB7Yi+AT4g5YH+ceB0tGEHXmowYBXQpsStDRy9NTy3ZYjQzY5qoEnf9WO
t+G+VwhMSwQwQPwBxTurEfLOQcZTvsV+uoX8GwRJ3gcFohZs9mw1pZCsUcr7HQkSGukqOSrNSXlp
4a2vg+spQQ/kw+arZ9SfHlfGzAUBV3nBmV1L6JYL6qc7bir+Nxs30LAk2wSSyni507Uhbvx+2A4J
64+G2OxYmZOu7xNk5DoO+M6+fwSXjxt5WgH5BTGiFlQLXrsi1FzMFjDYsAbcXCFyA/7YW8Ffa8Gt
0p5gHlPImOqvbJtUg5rbkUYcaDTmNrpIOXFhPq7YYCtO8d3sSd4uWQTluYFkOEqvrfaaBaEz3or4
H2g7YErfZBmLJ3J5y9y4Q34KRgAEaX4LVnAKHSkBe5S1ZvS94CwaQuFgkiCN3FV5JPkNFAuwXJ64
mfS8i1eZ1Q9WYRBZtmk3kbHevZGjHkkqnGfIf7oH1PjhV0mTelrw9WToX36nGiq9Uaiq1r3yrbXp
GHPDW2aZ23tPCdhad0ImZXFUhqfwbN7R3e8aszgbkm461c89koJhSEu672GnS9nSHtB8bpGeMy6z
sjc22FT2Bfh2p+jVzCIez1GPfIZDmD8lco8X68X4oYmqireRn1Ih5FULTeOK/AqbGJoTYQn3qugm
cuOm8YgZ9ZFrv/7QdwumA/g037W/dK8ydtjkwX+02XGoHtmWvCxw8BxQbDewtK+vC5QHBwdP1tZk
iLMgZw7OG2+HTYSi100Bj4W0i0oHJGHf+aZvHKn2o0Gyi9DlL+bMGweguBffIrBTo4Eh+hBNS3LB
vkyZ4Crsn1wS8DOi5T4/ZGVijRAVSAowPhlDYvJHiDMd3Ro+yUyd3QCbMnkUtFSVBOpcv61toIzj
JEbVnmAVk/VX6NO0HPHjsae55EBTV3I9DPJBI7U+FHrJGkBUuv3JdqZw5d7Q4a0xF4mydKYAxkFL
1K2H9VDIFw/DIIQ/SX7kb7tHPjBfavL3ukJN3u5TuKnXgReGJaHzXsn2qiEJ16Jpk1jGbQ9yHCGk
Yi7pHlTCBVP/XA66CSjB8uV0Gg1XN1C3Y6i/KRH5TzihntMey0Bn01vHT8SMAKUyrXo6NTLeQNZY
gcoz7KEFBPEBhumehkRmQtyY/908H4yBH/TwtT2Be/SItFGikKyY+pigcnGIiCPmAdS+UlQPaoVh
8++v71HffxM1+aIJS9Rr1B/WO4znxOOq7BzG6Jbz/Nbq5lGgLKC23TVd44lFED3NaY3jj3U4dQFN
/08wbtJwLut01NVpjNzla0vtcFu0BDqbRKqUHE2ccxcuiBdL2P/v4/Uc04aVbEzjJdQnwU+05Bww
BGgTS9VduHwELRxRJKU1xDgGLZ8Gx9oIbPtg6WOys735QG622q4cobqhdKjHQCDGATVjzwcZwZ32
xzxXqJd1iX6byQqAvBrdEMqKlHLlc5ePgh9KBx8u8dT7vYHVlCZtNxNcqM81t/i05yO7OVPwMoHr
V16E/F3I1nY3n6vv66OAiltTpcHvjqF9P23rd7AeRt2ciwq5sLMfe9NxXb+qkE58ANoEhYEyC61s
cLkGc5qDa2AkxORnDBPKx0VyBSJ9dwTkFuiy/nNZQX4FaupJO6086xdMw++2/7rmcFVNgEKItThq
BhS82OAX+tSFT5te2niKXcIVy/1YSDTweGg+aY2ZCE4vKwoXeM98iMSvQgRzAHPKW+i12AHG8oH8
+Iwpt6OMca6hYNmPFB5c1ih/bLq3NGVFca1iHF+A2FQqZzzkE0LLtoI82elVgMGF7eI1DV30aF5o
aMziqc6pR0VXS/43cCoYEcq1uaTTeQ7AckXA0uGSSaddJZFIQ1hylhWLfFKbtDZtHmdIO3CQX6wE
bkXJh5rkhyuKgzx4Wmdn/7tOTWdkwSyTxZB7fTXA3QQIZcvWLbybGWsgxwHZnyBuqoD1e2/ShvW+
8JBe4ERZ9bzzkNoUXmcyKhO/ZSiSOXP/20GGMfM/BY99U7MZ0kgF5s+yo6fhVg5TAIuNRViOaG/y
Ju87KFqRFy/PvvpVob1tl0GvSxoXUrI3cQ+rVmMYTOUDM1v5DK4j9+6KrfR4ATZadTh5geHrkjYc
02h+NhnXBrz18NpK2AO4exiTxrYXHj5t8ztcot6mJFNBu9smpwyQkh85w7aa0VrXN/r3rYlFQBRU
1Eczy3aKbM+WGoN2/LnIHVfU2XAvYh5qFL3Ot+j513JAaWYz0IfsoIWA6iu+0OybsHgenj0WDYj5
/0ea6s0PVgSMbehT/P52pJfNQChxmyl/RawrCf+jpQQHg6MBnY1uxBujglVk9YRTtl1TWm07aXzO
jSDPLqTbCdp5/+PHAIvMtBlxCdYy+d+S0cyt89GyKeYt/q/BwffjrKjzLWsFAJPTYuUeZqZg7Vfp
SUZLFeA5ZbilfNlU/lv+AijU0isa5WNp9vShACXuA+h0jx6tkC34jx8IKtro3EmYsiHxuVCfFGS9
U0REGQanEZOJRFhVLQ8i+a88SrwrtzxIquQSwgh72Nj45XMpCEl6i0Jh/2VB6ajPPAU6CT3LAn/x
VlaAhQQTylXmOQC/V65l6pNftFDxOnklqvLNUtVi5DvjQ897zDKKWZM9PR5CAP03SOkHLQBHJUKY
PfW+hE2SlwBFqztxKWCCqqIJAFSqs9Vw7QKnuQBWLPo0TyRo/Au2uNN35on9maqZr375bdO1PX+v
hNo04ePJresNE8681NkIPaCDHXy/10w5XOt/UcVY2LuHmWW6zk7kEeXZdJoXIsggCcaR0rBjoLm9
prwyskVYsnxs33r7tRgyGsX16cjAlLXptfoFyijPJ2gv+Rj++faQ4gi0bEf1CLN7t1jvu0f4+iC7
vx6EimRqpUbpmZ2hz1T9pkmYtBQW0kPC/pMK4ha/k41jBrJx4fcbRk2+7Mc/3ZiyBnTqgcxIfAEB
1V4ZZS560BetUFhQtZql+awDG0gdDt7TxGNuS2omctjb+gvXWRy0LO+2IBtQ+ZDoynwYw4RrCvhG
KUqpaz/5Dw6ftQcG2tdTESsByORd1PfPJbco1yUkUP0yE+CXGAPRkgLZ8Tqf+xWl83WBUGTtnP74
3ELsZ5oZVLTEP2db3AU/E/Kxaa5nly77LPbj6TlL6/L7eoHlejrvvMZH54HCbV3SPq+SF9RaE0V/
qpJKrX814v+WpjV9K8B3et0FMmnmehiR7LcrOVVo1oGNI1/GIx/hAVvQmjPLIWvz7OGrK/Vy6dsZ
sxWdksDBdr3mAb0IHWKcqnDDcp2JoA2W5BZpAo8sdldRPDHce+0LPOIS1bohWF2GEeTR7tz2t644
0sLA4SbuuWz9Fk8dlzRKOFwAU2UfMCQU861o1p99SruP5KUMc9IYqd86iogfMvj8Ku+zi1UP+RTX
Y3YaTA4VDXBUjsuYlTsR6ag4ZOGpBTNEx/2mB0yH1g2iMsd9PM78ZrxfLeiWJ8bQNvArfdE0wAz+
0qoOGjPZrg9Q1BlpOA1pUyxTwyfINf/RmhHvNtn3tpzOQ1jEvi+H2ioiWdEybiB9F+/vc0XK1U6h
LQ6hbglnW7YzF3BD4n6GPsvLWynp7adWsbWcSF66RP02SalJaOJOHOGMIQ9HGlk12wq4gbSX8BbA
rnOa31KqGv1IvRrPWL2FMpVqHrSLVpsxc92w7gMfBAoYwBE7lJDaKMipr04abjjmLHjcUqskeR8a
40V7agueW4Vodh9/3o3okVbJa3Z7b+bDnSa/qw6958KWAUVIMcNbx+a6jew49pUCsca4J9Ycq3F1
JipYM9u8XjbLfzBzonEvAh4kKdzWziHIt7QCtA5DDX+NTRLW/zSH+Nfu7FbDIRKGrcJdwJ3I+gze
QZEIAiS/MkCO6cdHRxmITmu5gIMIk1Nml6EGI7UnSdchAWNhULvQbrV0qpwGO3ILMZaHTU6XLhpB
fWJcQRM8BjaXPSO7UWGTmsuLIGtEboQ64fMeRtYo9szl5MKcawlj/80LrXwvHpk02taceaTphim/
IvGJWk0JEj0yCL/Mn4GjzVmkz7ZTOPKyXCbm5MZbZVdqpkxChydemFhFAojo6Jd+xyEtB7jlQlFo
LIMiQYC/mXrAxD9LNDdAsZ/eWGqq2ZxvSoDrWPOTWFCLngasnz90HEAefY76kWd/w8KQOR+xZzGf
vh7bpDXT7EUjxY3tBb0Uz7C1axUkseAA5O2bkpBq3J++XgC9W7ok0FaCCQFQerRMTKxOz6H9LAYk
pjuTna0UNI7EAP3klTbr7VGm2Mp0HbdAiUUv+gqe2qs/gnoJYe+S2trVz++cRFKmDydT8f3/w62r
OGZLn9/WJAioXHCG55VhrPQ2BTf+7bs+ZbOLiIl+P87htOUZAP+wIccOW/hlLz5mcGXKo9nu37y2
HEGbkwI1Vg8Ol+a9yE+vqIqp1GuK80Hu69a/wtOo3+xwByeJ15etioOEJwleo27SftMa63x80xgV
JdEVTrVol1zLvRcTvymw/DIrTALx9vR6tMHwlioUzzZ4/eOxXMkI2EL9rWH6kMCR0SZFOrKlfNlx
1XhX3cX1tXrQsIQTVwnCjUDHw5FYzLLe6lZQmmE0miSRnboIei4CCgkPkuiY7HrE8M5HZm71FK9r
CEMjPERQMf3fbYYNvCnkuwJNY/TQcYIu7LgO7tySJHnrfnn3Ul0E3h39oXO6jWWQa3etG80k/3/i
epNspWkmOy4cpr6LqgCmmvmV5aB02VUCanP8EHIncyw7pWZ/ajEo7BTD65RBt15DZBbAkkn3IgvO
BzkUUATIUR1hs0sEXpJmt4UM/aZLY21JGGhKVVf1yLt/wUFJsexDR0Cxfr2sBBJXy+MIOVYlGeNv
jGeVmkVFMYMzg5iIMTuydigu7koLo3JMMei78lFBq+mCtMwJx8ozK76995RVS7szTofWHS7/MSUW
Y13J6mLyWoUXA4yA7g705Tedo5I62j1ggsBSoX7gPCzT9JOo51Ry/vnHbUI5ClA5zcNbrsoLMBn5
V+NCoAVA+vqui7c+Asb2xVVHvD9cygdEb4s4bppH5zrHCYxVH6xmLvrXNS78Q03dHvfGrV1JPQva
KHX/r0Lt2d4Ma/lEaPLJH6UtLStqFDZiU4XM61eKnbgxUy2gmMk+X7qPiK1qOR2wNUEBGjHCZ3AG
hHPh72x/HkAiN0OawvSHr295aztL3GltcddyR9STa39LIWurfmaW3qNARXSFeU+MoqKf0/uaOapI
851Xl9eUN/xCUh0ahmb/dcm8Ft5lBXwb4UG3sUKnliWx6wo75O1u9Q9aihCzzUCAQS4tSbSrBVu9
8CnFtO4RFyhT09gpCuroLpicHcgwG285bX6IeT0GE+opYAgePc9p44ZsF0+U3h1iYa0PVEnPPM3N
+YhyKZ8SUzczsZ8DNYG60H91SPTf/8926s880aqwSPNnWlGCDZzQEKpyqGQuRmzCHPycKLq2kV0g
MvoasVtkSgpAXqs97soN2bKSUmhxCUbtSB6EMBe4Y9x2curk2UrS6B4eMp7B8e01Bm17iLjtPVmD
xVg/o9La9RaeHDXV+ef68/mgYLsdlXPLLiXQ5p3ZISmPGIPoTLzqGQVlDSykSUKK3IIlYChpDohz
TT8QFTAc36/D2S48RqdgVD6bDOWP8D+65M5g3m5YnCgtuBMIJr5Tdw0k5bgBuDwsY0ntE9LAXT39
3TEWN4pfzgb2Xtr2waPmtQ34rTVlVA0dwNA1VV9VP7vPf4RLq8z5X35Ft4CwIB8LO5xTfDuNTTR/
OQkzV4mIgZYaHJhkKf/ACAUjcanBvzIFVsx4vzTZxOfvWJ8jh8iMw7klphZ2YotUI5uysbf/ngV/
HC0jsOKH19SzN0F15yfFSofW89rfVRvtpqHMdoeQJ6v6kWpqVKrWSeaCGbhRZYSnVCg5maDwwhOc
If3VoL+rZSNV///fRamxPuUq29WQQ+UydUNDAjY0B/WZns9gM3R+7e5BUQEUATfhbh3qOxDToHaJ
y5ZPPe2BmY1yIr0NdveiPRx7P2PDsvCw1Sdl3tsbT3nOBlziJ5UDAenPg4pdqEdKpyI7xImfDr82
wePY1VVIfxYFsT6QuSxh7N53cZePU6/TAJWquD8RY/pNSXEfwbh8onlzT5IvDXHgQNvPh68PD8Lu
sNHU1O655rGhKJZ9ytrrOky8icTit2EomHgg351haDwOwrvOA7UREYA70oZHw+PzBOiTxz+L3uFM
xI1AwItgxbQSfCKnVR/PGIku6DQQewI/fsRR+DOnnKmhVmy7RwZKNJtEQNLCtG/ErUYXai/g3qf7
ZdlwJtUR6+UmRyaTSzYQ/g2FK/rSiW1HdQA1Rga/KKFqHqABsyeT5DpVsBdR9JwK4hGgFtXV5x5m
n378zOR17tCe4rz6lXlM+KUBDnsA+fSzHXfB/l3Y0jl+NVyvmxfk3CXkg2GFXt/gFW+ndaWCC2Wd
AkPdF5APjiE1eAM2g3V0ZbQEO2CY5iKo2PGw6yI13to1sm3/Sdt3iOwu+LfiP3/1gT96gTTKwRWO
mRB1SnCLs1xcwvVUotJ1htM7gHMK3+X/mfZok5U1m2CVCV+2U83uClDpMa19TNzuiWQJJ+VbbJ4h
YEAxjd2PICocITk/PgjQJmtTo7dsIugc80UeQZUooGIiUTILFvjyFdwuiXkbaaJz3+VxmBFS6mWt
nyS2Snns+Un5nnzxHI/ZDwU97iklfwq9e+MAXNyJTNej3gAciK+l0SrluLKL+fcHOySJ9YAH/gon
H/qbXh0LC+e0APDx6tOMtk0l6Tv5ieQXrmObf0/fshqY1RyfkERH3nCCjGkC2c7P4TIo2z3GcX5h
ixAj30a0L2PVxVJQ9QwriKbyodqhC7WTCv10LJxCLtUvh+LnjOeZX5yWSuvXe8IPIaEfjae89eqW
pkBGQvpfwfgOSz2waf9QG3QKhQf4f1Xw8Apo+9CxX3YS3tmL6nJqVy6q9G5PVsEklODFdIdTUkzr
QJncuDkWE1FgdZFkyzaXSWDsDmB4fdJ1gy5bhdKJtezjgbmFZRY++prcNu7Lo6Phvxnn34o0XBg1
OAyU48M9FZG7DUcN5Bc3D4HHaHF22tREE8DEtMPARzehhtqj1OOdBi9CdU27Rz659n6CvnfVe8Z2
udrYv/FFDFMhpYhnin7yH58X72qUyCn7S3BY3tg6l/rPMWa4mHO/VZG8g8Vi77s7caU8RAYobDkq
MKLxyynI7oUiF6OL3mOE+IwYSCxEuhUEJc1WyHz5mnt3lja0nSnpSL92kKWMVwl3elsrsVDQ8i93
eekKJ3W8wh8XjHY3KRiLA1z/9TKYYvsE1vp1uRaHF/sqO/Tq1PxwKOLboqR6jxdurtomheL2Wgp5
HmmjTlgDCteGDtOGD1yWnZCYDoRpdAXEM8kiIE5Cp7s+feeXyawx4rr6uW/Vwmybr0Ihlxs1eFdx
mvt+NAbujMVLIUWnHVsiWfpHtS2hUJNiGzF/7IWAzKDcaoJ3k+N51F2Mg31LtbBRNp9qOpqerrjG
UnBZ8TRkCSpxtvjCQGS7boR9RVXxSl9msUyF/rpCrG9oJdRMeWvNvjzczfzOA6zkJT5KY7qWeNTf
np1MEUWzATvgv3hDpDRw3ua7MJKWp2sM3JneNFqlqCtXwcRmwjRaJ78iTGP7oagxps23ydyYjVwA
t4Y/21Xl+NXgcanuF1d94VwnslEdvGi5Bd0mAjsp591kihOgy9E/mpzlcOf/CJe0w4JF4LYFnrZ7
rG0fU+/59sZiwV6bQAkvYE6hUCtt7IWnePQZCVoRDF/HHyR6MBwX19fRnnxe2A4emLbswu9ypFwG
RwVtrJ4iWoCgZIhjeSIL4QoLzRPWDhokOIhZFxnkvMoxn4xhNM4/BhBSJ2EfUpNaFZspROvAb5Dt
zun2jOFMPqLmeyr8O4vqBjcXegkApvNJot9Q9ztn68fDmQm3vXItkRaOOZ8wnirJedfbaDjD6cAM
nezVau6G69EVM783B3aupbVf+kjkqCA2ls0Vj54QhVjzXCi6gjPLz9wOKoXrIbEfi/k3eYBZ9ZS3
qUzupdQBdOC346ctFDQwWJFVYLnmsrGAj1VgYHtG9AJvXTx1amGYw+N9FiAzPbnJh6b/+yqIs97G
3pY19l3caa6EMXatmhFT+ZK6wIv+OXYyBBmjtiLPfdTZII1fBefHB+mRfGs9zHKbNePNI52BpXMk
AQE95fuuCwkOwKFD93vREqdPo9Z2lp5XoprpeQ6xt13j+1W6L1RAp39Yl/L0d0ghjZJQWIsXRHeu
aIdxjfSTV79B7HHA86kU6fyhk068xGm1WA3CE+v839qK7NaYlXnEqCVsLh7zdecqqJRVLNJvCcNW
fa75Bl8nOcFBiwVNR8s4CgWIzHRx+ipznASr9GSBsxoy+66M4f2XJ3+YzIVeZ7M6pPVwzyfaqtf6
x/qo3gmLbRKwN7d3Gj9C7ni3ns1+piLsFtmZnYW+4zSZdEDQR3DhP1zfHs+wo+RL1ptXa/Raxalj
ouT10YGojzrKziwrPoJzlzhvm3Zim5Y9Zq8MvPhkJyoSiPZZiZ5TZVl5G6s7tIUGjIHMx5QGQoVt
Wsl5H+pAlbh4MSYfG8TjmPEkA3ExccQpZuyDWQDiMes/d5IYlZ6NkxnJivjHvrecYkTTD0VFTQz5
JtQqi5fNmDpEd3m5IttuG+MoYC2WpgZ0YD8iT7VINoITUt1qZYBSOZQP5vuXwVzL7f036hbjbwYM
O558jxxFFaZNK3oG5+XtwKh4i7ECnQkWM4a3mOI1B6g++rI3pilL9eI/DtxNXDfbodHYagMM70Nb
D7gMSn1l2DwnJSXiw+Psy85VtpDrGGOC3ER6dgKRCfFgI26g7bZcIQGlTg5iUB8dK4JiVTtcxgQ7
QC+qak9AoV1e0ElaBrhxVZ1mxe16AYkDZCPP8alf3LqvUFFaPsaNUR9XoXHWZEEinVYis1825BUn
AQqh96tUB+aAS4TCU4nYmWzr6rDwpajW6lkVyhk8KFvkdzOGSSCZiLQc6h+fMEkk3lnM3gwkqWyT
0HGVfy7EWEW8qtxZNTpN5a69eDgJ+KOPncuQsbozgbUDkG2rlc1gxXmAP6TcYvze72hz/jikoEqy
YfFxZtLlnYQaRc68H0Hw/8VRBMx9KUqtgzGrgcOHQv3Um/ke0kMmWc+ast374VAuMNAiBC6GTeRp
sxPYlwCxVgMTv7XziJlrTGf9Fb7UW1U802jYmvrDcKqy3gQTKuH7Xi0bvYAZ9RTwbomY5g50yj2M
VUF8mx01CJkJXJ0sIHMWX/aPRVq7fpeQJnkDAhYaQUT2GIbJR2O1KBPHKIsEk+fr937E+lPXsEBK
NaUDngOrGHtrYZcvEJcqlo0gf8ONtqYydxnS+vQYhssSGNv9fcnTHGoaNY2tw0O9EO7DsDEycu7h
GR06sXoHcR0arrcGbEzAK1LWQUTX97/NOOkM94gp8TEysoLleUbwgeeCtBcSlVjul8hgeF7EBikT
eThheoJF2Oc0PIgpez9erBahb1wXnTFDWUanLSrawRo/+YbowBmdE5EBlYmk5quznpiEALkoZakJ
oHjRRngRPm8ho7CWCuxMqFf/awb3/ew6JAN4UotPrtYyAIqMYnJ+1ckTCYfak+49mCFA+AnPheXL
GA5SmCynMr1VJFPgghGDAVw3lqGZl65ghidWJDTpMgA2PiZhLVO5QfoH5Alg28MIROhLyoypDdo5
IMh4XTcWy8N3ACDyJz6KlHKkC3SA/kDcUTxuwUZQQvABupGd/JLbqyZAby3mf7myQ0ON68Mqehyl
LyKWEs6RNdwsrMosRlOSyatdIV2cn40U1mz1wfORS0eBTO0zqyCoJpOomz8+/tLD8mBD4F9dWlSW
HG8KBsSitkiFpFZomdrzzWHTFhqwhPQ81n6ZfkYZODZ0XNUmqa3DbbHOobsg+cnCoLZM6yLq80hY
YF7J60+QDScDJTgBbdzZF8eKNoHFCUceUbvjr3keqpczU0IbvXR9NlznjOz6Fxgp9vL5d2dQvkLE
bKuKHJAFAJjWqByyoVbfOy+NwiXJMXmNHkCZOnTiC2/PMnahllv0+bJar7atZUWFmwRQG8esEaKM
kBXngC1M4kn96UXm9xeSZOk7KPIgvHExtGkp9TuZ1HhDsqgZ4oUOBqUop3vc7632FKwGpDKUABBq
lK8qf2qmWWqD31gXpxJNvVhXbnbtOLlLcxG1lN4aYiov5URXrsL9HNP5hFWwXl0hQhwPbfqMhgQW
Y6bqE+KclGBEmrRTiR3m3EyOh3xXo0sS7Jnh/DfpfBinR8Wj5HpTrto6wgGGPt/uN+2Ssi1Z/gbV
3MaIMBPodl7fb1Y4Y6oDOanz+h0v4I51P/w3jHaVD+ndxde53Y4xg9X0HzVsEw6Bx4yIwfiJJB4+
J1bzs2z2X4iFMCPpo1nyh1dhlbNS72BFjTRqLtUKQAVqYDuqQXa7jWXYPJBlJJ3bDs5/vPWGu9N5
rAQnWQHV/WOfulWx++1hAP5f+PvDV+oLiP3dCKeDkOTexObOTuMexaImdPa7m8NzVZ0KIL99PbpO
FeZtXR73XR7sy/DcQjRMHvQZUcv31hsgQy4LCofp9UC1GgSo3XF+Ul78hCL2LFz/AUgYlT0rHjcl
vRFM62PP4cKLU2ENequjZF05++tVSUUkJ0VQnyMB+R3nR/KoL+1bDh7kuEaMlAxdg9n/ZLZfGS99
vu9ttsX+9eYTUY1RgG3MPA95p2WUMVjWxU0QQ71Vrr2Wroti1Ot7hQ9e0y9W8WAfHCVeFh8qZDcu
ozwP4fo6g0Ni08b8t4LXs1MI7E+km6gpBhJryeTiINp3qD/lZNwyuvFT3u3K+B3xo4sEWaV5kc8T
fuk3W1lh033ACvK7WAiq7CzpST5TLmg6IG2cFfDvIrkcEWYccbkxeTHr+QD9B2sJgNTmSSyC/bcw
STGoYk+qRovHTx6atTjG522Z6SP0WUp/2H5KTvk9GH7LEyTqdRy6JxOxmT8FnKQwXGbTEPURc1Ig
m4KUnf2LPrVsm0kTLO26zK8ue58nNzMUG9mYYXTT+LK1i2pM2p76TprKfVd9HYsRQyD5ZYlQ1aft
C91IdrPuhEJ2S/tl9mv3OeP7tGl29cydnRkov09lckxQcFP3Pb1ASyISbmbDQU07kGv9AJzd+pxr
wLXrFwnf6Uc93LYmRtO+ztEUJOQdyckZVVU97bOmyQ8esgcSyW/aveBUGusklYQ4+r0AtypFMQwU
G4R0yvjKoScmdtikz6IRE99i/CIiGLu4OHJ552aavJjnAeV2efMlJLZuSF7LMi9PsmWjSdaWQugQ
2tY/irFqpvBhIuuGZUMmeyhGA94vfEZ8Ujs5chWokxxPOScwo8uTvVmaPqrI8hy7zqKf6aAYbp6q
zL0x09OajDphxf4cv0ZQpOocFWUnjdI1uH+h6vGikt6M+61LqHp+BS+6d6S1mKWmT9Bjs5HSMPxi
V+KUoc6Y/HoBUX6uKlpCRaD0nxcjyuGvGD09+LUuconS0R+na4UZRaU/lGjN0dYZnCQpBbG/nYzk
tKftOjkEBUgb+UYfH7wTgmdDPdB2Mhof+sfvhjkobRNdewT1htAMdaVgz23/dFK6az5URbAqSzAg
aM90rTpDegHyGnuO9pBpyGPmU82GMMxRLFrYx3a933NOSmXaUOKOeoErV/Mllj0S/+brpgwb1INm
ocl6QzF4zo0b/nJhr4DS35Z1vjAa+Sg15h7RSKrX27dZ6e2OmPl/EGE7YZaq0nYmO2FpnD+Q6PFq
NRd3ZpLziCS26Zo+zdBqKkKA0TrbzjGaehbVXIRO5TSK3GuH69CGOPEySfpxnx0iUnAsZWiYKyfc
tFI1wF1oRwU7f2tIIMPqx8GVwEN1qI3TfTtfZBNh/FuorUCFP4UMoVbDjiZioIbkJ+ShKA32qOGY
Er2rnAYvHQricpeJ9vhg2/o9EvydfaxUKIrr/K+3ZXqi8/pGjbOOdeMXbzjxChZGiDTlWWVuyJqz
RNFal7s33DK5L5n6prFqG073i/C0rK7vcq7/AOCxGDoIbHk84NStuUkmnBCMwSsxeayBTK20WuSJ
BkjS3tb53iXlOKTnoj3SRSB+n9SbW/inPPaAFr3DK6BbZZkx5OoU7AVNrhEEaYcCLYlHJDs4Fu1E
i+v3rAlSSjKe+Fq1zo1c2Logq3+rhkb84yQU7/WuhOOA65cemapoGAhXU8ipc0HuYblFxO6K3nGu
RuhYRP98zmNHDX5P/u3xDEAuxU07e6HZDsgBFKnTz9ILe/shfpvQlmliU4/Oo0IAvLW2S3I4PLbA
DrD7cCTG11zg4bdBhSp5E+XkeM+TkEVFs6yectah+G0oR1D4u0ULFjRwSLN4oJ1P2lVdUwJUSGZ6
eENIh1D/jKKaSypqGaqNINnCpoQsLnkJ2UZcW4YvD3iQzuT8K6SW5EGxDWJ709oZj16uErFSjiuE
/ip00steJmbel3LROlSW4EEaKAKfC/+DBZnT9KLRoYTbqJQWrPwatemfxZtmUby2oxpo+rwehEuE
FGEI4nlK5kODgIb9VGHccdnmGLbkDfwVh9BzvWNQsVJs2Ejci6e4wUb+CL36zLCSm0Ak1KN2hTA9
IRodTd9RDCoo5BYZarDo+ora9wb8K593qnSyQCu5KlnqFGM+uE3mLuKSFU6oYcL/1oPEqxp7XVhK
unGfONyhF4K6Gc7F0fmHk9QaFwiagc/FdDHQ7WLImAFMK8t6aOAZ9lhJyvRnI693k9BrVwWxhLdr
560Hbb7dXNezi64czdU3RlvfM2GxOfdWhVedFyeIv+OBu07Tjp4/lt4dfyYl4tWZcBBQ8kxKY58S
yJG98sP5cdPoZ/O319G/YTRXa5h0mCh9P0h/aUiRYN4LXycJ3VOahcj55qGz0itp1z4mFr4F0T0h
uERQlA0jBZFf2Z1tKT44UsNYqrwY6NUPc/AmU5i/T8qHJecspIMD+4YPTPplrsgXbB1CYlSW1/cg
KGKNGbHUYpebTd5E5M11cGnhttJOuseiylyjzdyzlZbgo0Sfdln5bwPIVNCziK7/j3CoZJzLg5Hk
j9EN5pdFknESvQK1KRdvTlMjqKNvcVP2IQYmqn/4ZVB0f376eejG7bCktDMRHoHG1bVhz+Kqd0vP
rUwwByUKU+f1gLcq3gWV/BfggE0c4jZygV1G3Ui5sr9IEMdN0b3xeOEafWpRQtWndvb2gGnGrlfT
K/fzVJ3it5eA1UJDGVkP9QiR0hWwyBcK7l92Sq+mjg6bYZXz6ydeq7plF+bKusC9bhjyNMZezKzw
FIHp24OtVuCOYNW5I+a7DIVjzij67MdzyrgGNVYrBsfkHJAfL5vegpCuHCUurSFA5GJgQnPnEkQe
ZODsceP7I5e9vnCTALtQ2l1pFDoUNEV6Pxxtql+WaCDohB48YMVDd9LXUXONfsD5PelaUKPGq/mJ
W4Szp0xAE+6V+Y4B97reEqADi5IkrfZXI1KF/cTKyqIV0f8TgkLsCFnuqUXcwgSh6ESoAv0vTh2Y
dSsO7yu1HMpwry7aK+bBiM5mXUDXekxjrjnYLXBQ+sFSfqEAqqKlXEYM11NpDiDCtko4s3Ur4B9R
VHPo6xB/YwQBYNHUAhynuS/FivOGI+/E7GKS7Zr3HqrKsCoQEoBv0QeHnYNzz2Gb3nsEFjUQaMqk
bH4gEnxZeVVpXGD/IofUR7POujC4FexS3XxM+7hbxCA+CX7PAbgZe6tytDbHNu3CgLotpJgEXqMH
68f0vxaLs7bwtA/p8UkhJ9YJKyWA7Fi87IEnDwWDHn7sKSB2MsDbg0zsozCGCE+5QvuYIO78Vw5G
YmlbG8o991pFP2nW5zSGRYiqBwt+tI1lo9ThThHn9Z8hNhjOA2gMKf5HcIbxtI5aL2DG2KseDqDW
sn5oyPHcpBdxchG/zv0fS66heuUi//8iLdHJg4c97Z22DMk/swuOE9ceBTjndntBqDdOFxosx2Mk
y41USGpyryTr5kXvIin61c+lCzqQvql4A1sn116C5gdv9w+smw8rflBAGc/I7HnWs+wFpTK+Xhm6
/dr0GnucMMF6ZhuQlnKy7YwK2NC+EijZAOVQvBOLFc6TQ/jOKl4w8kEgFuMJ+5G+6UL6m9ExyDvU
H5bERMn3ADYw4IzlNESq9UMGJgliIOCTXZfoTz23algPnNayPWzmDsNaqijkha3T9IkEXSA60XEg
nPskQ5UF6JYJFtkJB9zeL27xeFteJm2860NOAr6uTVZJ4W+I76fBmW1qebAY0XejNoU248PPGVHN
jnPiNtdaruD/xJis8TU3R4sO6UWcPb6MS4GmOCP92cz+WIHkcSA/kzb+Zj3NhLgFrttcJyr5hG0i
KXT+YLkQH/nNiY39D1gSdwHCq8vNj15SH9eXt/4d6i3BlDyeUfpIuVaGJu98waxoaud2ViP6rCFJ
OpRWnROzkgmCOjKRZrOHfVevsiurHbAkorue2Elmqh7yaHbuvWOQBeRVk1CZPc+pz55Azr+moXbA
iM8J6t9F1/O2SVdQDKGnWQ0mE6V2rylGVNFwvmEYX9XhV/Id3qGhS2avZ8TcQAWc0ELEndvMdyK3
1EGRpJK3iY8EMX62osgkfSBlSv3yOgPGVMBIZUU7gwOA+XuqzJzU+CYbQu+64JLEr7/zownND52A
J90OCMHbR93/tZjBU/qXhatuRmCZtgNeje3qRaBWczFzdZ8KBYczltz1pnGYRfY1ZdPaIuVdpMB1
FPgvakDlitJcgXca0ZGdcWWFcQC51pwDmZsaKpPAlrPQmHdXkpPiIBOhqpBXWI1SGGqW8pFme4Ap
7FiePQTTaFxU7iYVOAMmoZvn/W2fjdyM3Ks9bLOuUn51Ka/OAli27v2B31P72EjCjxZ9I5byC3HI
BouLSvOV2lgemYUt9tvF1QJD70MwM3DZ7OJ/AaAzlk2OIfFHIRkkt/yGlakJVbb4/qzn1dqix48f
C1KooBav/XLrSEs+aj9s/zc4aKxwAxijpliImG0Buf9d+deJv13+nc5/7xbOJR6ix/6rGY5I/bGj
Z22+ZZswMSvzbFTsCx3DkJWmFq9+NMHizsTaPg4CW3j0/SnEyS0SfV35JjPQJcVSvPZNcQ+Ogxio
1EhyMQTkJERhZnXxoXvtym1y0CVbq4SNY28vdtRQwrp/pjuR/aZ8Jz+pMX8b0LcZTH552fhl+YwK
kElmz955T4yYBwM0h881bfM75CNq1qJJDfK6es/L7b2qbtU7hGHGxY3bO3Olf33NK9+mh1idtj19
DOzYJyJY0ztmVb57Q/zgY5pA1du4V16Z8Kwlmx4X2h1mT7w5p8lC+3bwjvsjxTT47pQhH1Ztf3Zh
4pF1F+phiLs7+V9u6J7DPFYJU3XQr8CZKHpNtDRyU3asJq8yQYzpJ8Qm0lPYn2CM+95s0fauB7dw
vUyDiwwKIG5+0fg6+izo4qDF1BDNv1ojBffMXOyAVvwrvvqKl7FLqgWBs3WZPEMQOEZ95urX1/sf
Kn3zs/xazVXfliqi2S+uV9n3JdpgQu4qELkHDltlrgPur9gVNTJcinHZM1taKhF2kzoajbtLZ0oY
OrXsatFbhNlUpFUL47fCZAUCSB0frkGelvsdl24aTguGIaIbrIyAcfpPe/+GNSAhp3bLOv+sBjJ1
AIcsvUdBCWq6DsE9N1vZf9j+l1wNufKmp493Uj7y2l+RQvRLrhIdsXcNd8EQ1L9RBHuRiOxGy8gV
KBpU9r3BqyLEA8DpZlOf59ZtBUy1hjV+HNDcG+Mshlpfcz8nnlTIhHlnQOKZ5mZzkfYfEsQuqNTZ
2dUph5LpVe58PPWZDPZ4s3Bj6+C+KKpYLmV23/FUOJWzMEthddQ2SJP2l3Np4a/2SUYO98SfHpfO
tdAipwrDkpVpxeFW8D29LsLXQU+eE1547/4ZiVlypvlgm+3AVIwRDjnz+ooRwcucNZabtWoODtWa
7RU+zNuzRAOerk+m4rv8FcUJCYG7oQJXBJtg+YkNQ8JDlb90n97m0bpjCHPW5ZNsf7HXRtFubdqA
qTo3P6WLJfhmqxNZncaZaGl0Q8+rGEdaKqbhaN+YNYnK13c840+7SNmTQ33VAJMA8E3LTEWIX8ue
8kxUlB9zGR1yrE644PdlsefCoQsvzd+pje+zrepGRgirr0VYI/1W5VHRmr5fTJVfEQ6sCuZSEoqs
10pSJHD0PeHHPkhz1WIuqwXgEBDhUfM7dsvaQ/m0I8vkliyC/77t/Ex1WCm92E0sl+09GWm7KHlI
OOdE7fg9HkyR4alCJCw/CWdMkYoNx49CftoBNuKx8hp1xZn9JWZSjPYcBSIFUY+tiJJAAG8Wm3HM
HF0YA2XsC/QbIzyInVEgHy6pxmGjLTRs+1byj2Nk1sc7ZA7blHC/Xpu5j0DRJrXEQ2disk4mEZA4
xSiFz9YWAC0OU6fOPP90eRNsKcfAGjwY11BZqRwlnt3ddgn25omW3oysYPHsrvEecY5RzLoxxZw1
g2G68shdVjZORJqCZ/XDTBpw65YG7KWAaF7qrmctgNnO9919j+jDdccI0G0CqqS7G1HyABXGh644
5AzuEUuU7lbcKjj0pqqYDnY5242IEKQyeI3Ly+WeSxYJFf4NZ7pBDtl9S+HUSfTAFCVy3zArqlab
I3J1c5qcZRxZNI2IKLBnRzgVrmW5zHAAgfsINezG46SYc5P9QZPCvW9hhne9nGGZdeuJ3nMtVrId
Lfv6f/qwyRfwC7ASLrvjQDM5MxpZwl7iLq9RzKi7qA+pKqlrBx27dnk6DeZeMnHJ7pbeU8/TSDjo
8hakgh0RNw95mwlvrQFIIRsgx3vJvrG+vRcJiu6NV26bN2IWrcP2YjiWSU7iuXYZHE0ydrMtFIyW
iDoP1sDMQcCBN3G1T6GiSjP+qdDG+gD2jWTpdC7T5byh0nult7HPM0YylTdcgKAHcR5Hm4KX6Zjg
KRQPnCVCHMSV/3j+Xd9zz+3O8vCva2IW97Te+FMlzXCbjQtc3mAM+iLBxDEUQlPGpG8LqqA5WLPp
z/4Y/tbjhovwgntBHejfEgxIT1/5LS63WRoWufzf12j2aab+vjVftiLbhCoyPEC4G/7Ao7wYChlV
ibScA0zXSleGv6tHjqUqA3YA+kX1A0N523osmWKMGx/nhO9cMdvC0vQD51D4He+wm1sfGq1QLeiX
fhCc4CyuAdcWfnCRrMLvLQaFBgetcUOPxoa+kcn772RL6VYlj8lKoIEDbsfBKsu4bl7QQX643O0H
O6Q5Y2vGTMej1t/1W6rSRSg+fTNBqSXpCSndqdeWvuq8ZiAceuyufgkMPNvWfK+enSyDiZ0rfAxu
aKSgBCVjnJWXJo0nPPNgxZ1f35JY5OUFjlGNHSzUCRbfuz1HvhWwlMDbxB0d/SZUcaXLRmBp00uE
bPvxiN4/FYrKMh9LIPzmil91YxqBEr6FkptvR7VvOGUsjPb2OjVExRJTDvwspHoAFsJ0hmjKCENh
30zX/wjBFuzDTkzu0rwSjcNCeLCTrUmiDIDLRAecc6d8Dds4TIckPX6q0275pSRRW69hxEHRWLgq
Qz07qhq0mpBIg9EAAiFQTJYGPz0Sx+QQsjLo0QAizwCWubZP5H7wTAXTA139RUnYyuiKboedvmTP
vcAZyDu/l03c47hvRvUApq+O/8gjE/iwbr5AnJM2cr8LK3I3CpmBkWFSZfUKQ4TW4ZNeJV9mshgg
19Swc8ENjYQ89By38piVwcwMfGMKm90GvqonirxJHC73W8Y/t96WxNpduVPkTlhDfVghJbh9RNgr
SI0ErUSSL3SSHYFya2QR1m2uOshKOGI0/0DBPQATYbmAK2g43V+xENLBufmvs6uTzTVF5qSFQAaf
imCRT8tuiPMaIVEubqMmxCD5USvwP7yzN8B7kCwy1T8Njr6S2nPnQ4+Zfz1d72p1y80Jdbkoj1Dg
Tj3wm4AzLCovBeUc4yvk5X9FyX7e6IjxprcgUFxM5JQPVWk78x312ZDvm9czOyvlJSi+wwXF780i
W47od9GSUzZhkIodIvLQY4L3qacvONp3huHAIkZOSHOPf/BeEJOVrcXNGFiLpmNZxfkquTqawgCv
NjS0+glGYzTwJWcpXmKbntEPcztkCBlZnnuERV0nhu04db+QKnychyV0NKXbNvnG5ITnfIhcoENc
+J7ldj9pWClCbjhhG7aU1/6vwGt0ZvRHvh21qbKtq5RyZeB6kXmFk0PtojqFjtQSF2U8wiWO81mt
xGPAnZmUNNriSNT3kYpMZ1/NmPkbUbnBiI6ztKI/9kYpuqgvFLosjEmUmO1nRBi/JVZ98T/yfBGx
c9PmHv+xGuKjM9K0FRsvclqdZQmh19SoGos/Xd4dMkqlUUFG1Us9/pGCW4rDPxARaLIM9OJL4ZCq
It2c9pnOwh2r/zEEyWp8cmiecpFXKsWM2KmnB/+e73pSOj8huHnqZsH0cYEbvOb08dDHeyle5LWV
4Eqidz5Gd0pEWnI0XtOYVEqKQKqxn/BYhSvPxCsy3VduRLH+sP4G8cGwcM3ICxbOp427YG7JlVje
1QgNLB7iUpZbFV0rm3IZ2pyluRaBsgGWe2q8mm5bI0Szz/WP14Zuwj9iUxdaIXjXiUb72RjOiO5F
mIvVQi2M0+8rAW0C4ENH51PN7+W+n6VjxgP7rHHCa7PNxUXej0F8/FBts5jyHgcksEnYdzlLAfqi
7p3PFSqL76QQE7znfJg+A8jpQ3LmbPI70eZY4/H0kA2LZ1zusOhh9d9+oV+79WDKhdnBbca2soSM
I7lMR8uA8gZ4czatf2no1aMLstLjTQuPzjIp9aTYfVCkJjK/ELOOUTc0qnveC7mjk7s0m2HOgN2C
+bzAxmzq78sHizMp45OlUmalpzQfq9VTZVUKjHfrSsJhbM0nKx9PaV8TZX1VxMQ4YksVtcZivxW4
Y9PYGMTahFGXBOSLmfMjdl5jOp5+E0Ck3jOreSnH31sIcYLrS9XUGAKAN6MOy9Su8U33/WQ4/6Fo
oCX6OMRbExQt3BqjCCmCHD+J6N6DVcczz4XF9ECsdy7kXZ4PEb82Uc77hJEkneyBUxtSAIT94ylA
zjTTwSquvj+lNEBin//z5716y4tZnisnBpzOujZL3wEN5TD+oQSz7FAASsjXedxd3010eIJRwil1
7GtFhoGFDfQVyGUa1Nsv3c9qOnbqUonDnHtQpg0s0Nrxl5N6a55EMq3VOMJddLGER8KN/+L9iYDS
zZkIM093ZzFYHjslIZhpMfdpNF+Ba4E/eE+/PLzKj364nhkqhHiluG5sOfE2uU1AbwmZ0bf9kcij
sbHKyW733duNdtVTq3O9xFixjPWZx7MrESpOjEgrdJgBrbTzuj7vqPKvaUtbWxgv03aQUp2xefag
F4x/AmPxdEaYfXwoMvYRTYG96H+BxHvwxjKZvVwWnCZlHtHHGS6yVC9lfVvSegzKwiT9L3mCvtA0
I4w31+f5PA08n7OyiN1Htdx09sKy43+g5glj6kD1vrQVmxJ2ymgZOGBf3XC/r3zkiOPPa/z2a7lt
Mnq0VCBpQ5NZd/rpy109vkCrMUmTwAr4crUdyQkBbQuRv0lmHz6NXQ4g5STbTcilGncHoKxYMsiV
qQjGY3SyreMZvY7hABePwKWtiL5+c8QBHAgthX0gsAirXS9xCEKw7yyHAA4M8jKOaIBfTh5u85pA
DPLti9VUEHWzzADTyZuQjfFFjnXMshtEZauwDxrk+DXyVHovzLJUVOmm9bG8KVgIrs2uYx+9ufzT
t5ZDGz835SP1hkLqmDUMeySf/uBPeeFjodX18Z/1XcXw8Rw+dvFEJEb0PAN6DI8QpYjBfJPZ74R5
C1T6yDOzIqFnKNnX6fD0GVsfqmRkJ9poIBkSsRrhKESAWz59z0qkZQRwn8e+gDLpPaagKbbtXozJ
xxGmOsZpF1dawizHxygo0NBgNgl0rqLLhnbbXAyV2HUV+WacUHYZbzDW0yNJ8lttYqeyDTJ1+hjq
47aPCSvmgYuTvyAtIHIKNvGs42lpW+lvga8h/4KmXZ8hCo1HL90P0eWIyP+Y+6lMzz1Qays93U1N
lJWTgfKSnGOiLTkP7EDJgrW+B7E/LA9gkoGKLz9l6tNXHsdI+O4ZC3PJbrpdEJx/oZ988ZfpQa1F
GmxKyS9ma0rmZPdCqG0x5xyJil/+19VTKaDR3EdKkbWu73V2gdSu0fknKI0xz+5Oj03mQ9RAOqdz
LCeUFPoJDdQQo3ohjntUM8r43ovw3RO+KYd9H/zCkDsnpcO/W1K2YaTAj7aoRuryWEfw0vhkrxoI
DwvYlJhgQwfm/9sh0WYp86Uyob3uls+rBQHjP+TQQAPwEPeaIK6HQpD/Z6wHq+Vo4PLw4jqAGTMq
Z1KKtKGtNHs79oUZpFRjP6g0xRZN62VH0xhWLRS59d4+SjSwItPrV3gaWjqtt++sVboVpD6B1BJz
D8tpZtgTFwQVwJdzGiepumFLT7HQCWfaPKLrv1l2ElKhOOGUUIc1cwFHj/vDAid+gOvBGGb8I24G
dw/N+10+XZFDyOYjVnXXm2BUHVfmLxoN2FUtyGiR+eqN9pr7ifp/BKi/qKt0Wt27qJoLiNRvWUKf
tz2IhffhoCkGSH+V/J1kK99UNIPC0jxmViBUp7yFUiZGDZ9HHmlQdIj0P/bPTC9nOjjUfNFKSEm/
1ei+Fii8XucwaoCr8XoqQeNIgQT8aCoVa6MgTJ0ZkNXN78EivmaDa9ZBJDj/fgC9+Q8N5nMTW1rb
Y3d/IFFASiOJ+/zyj/pTH2f3PIdkBSnfS5EqfNy4nRHkK6H3dW/PoEuVcboM59TD5msD0eR9pVZd
/DYBo3vqkV32NRo7ofR1ARrvtjtIm1LdhJzGprbX9yOOJMN5mw7uNHGitM6vxmowperugxGe4SSZ
OlgCNIC/uhlznxpl3o1exMXqbhM3bQi5Gi0pGXkz7edIx6OalPLUgaRcoqJObzNqbOA0rAgzu2Pg
/WxdPpu/OxsxFRi3dlRGk6S+4Z2RH/7IdYJ1ncNNwvBEbvlyE1j+wF7Fq313nREDCm9+/taZaoUj
o6QIZPMqIjplhRTWvFaPLvUx/5aIrnnxQLXm3jtpb7bpMi6vJIl+ionQ/uwFJ6GSrIkD4W6eZJdl
zTJPdLQJyCh9c21Xc/Aylf0QRiduNk7bYZjlJY9vkQzVC2FvEMCJi+Kd6yfeWtMFQl2dIw+HYr+J
7IQ1blXCm2263egDtcZCG1LYP5cQ8FxUQhFRGrf2ddei81wOLBIMQJc5xFUIpLsZQIA4WHIudt66
mssvXKZW+mr7PxmXBxVkI+9rFle6BwPHuyX0hogmmbbtK1kK7+mFUe44CrzWVTB0EQ011/ymL4S8
D6+pjUd51zS9k5o768d9sb4gyDazsQEG0Vmh//uinlG8qIDXCGLm5HV9zx0fmGkOMqxJwlZrCxoq
qgQgYeKuNZpNzasIAbSFlL1fXM0+NXlZEM3tW9XMdnW0yxnmu55F0wClS1X74XUxVYjSrUMmi8yu
qPTgsZjjD8vgyKoabyNWDm2keTUtx9hUPl6MtG27nXpoIWYW2daRZJ8DjzMym/hPCvsCPUO/9kvD
UnhqnyluisOltQiLo2njFRi9Yq10OQHhMCcIx3iun5EOhsLB6CYN17Neem4kCVbSSRGG3FqR7EoL
mrr/EtBH6tVyHg7eIgIDq2DZqBA1U/KgZpwbHkOQKeP13Mj2gpca6MMrkHpRBKd8QVF9LMtLbMPv
EzUFYUpBHOVSMlvJBAoklrEsUffoHSx7Slco87IflHxRcmCWQJQh+QkrlguzkmzDrhM65mkCK82V
xhEsOp7BDoAzLvNK/FA57oMa0fG2AO/bgwjycBIFoNkXvX8XJo3r8H5kOxf+lvwGdX+/fzhkbkbs
O5Jtp3Bgd9f066eVGWvuzbDAxsIotAksZQGKU8vlbd0jUf5EEUqYdXneB3vljtPEX1b1WfLdjd39
uI7Bq+QGfFd6x2h04n9mJjQL9rdKNfc3hDodCskJs++PjYhBVEtfGIFrqtI17TZZmufMjehJ5T8i
RnrK+KAf6k9LjzgG6XqFmvBylGuMQPdfflhQjB10xRvJg5XWEoTixa1ozm+zr02Q6D16OEgm+1wz
vAlhYW9MEKkwQIQ9Sgw7+RuVvri0hDyMyZhOnjMXawYk6RakuxofGM0taIhGILUehhbih27aYBpA
BsnYPv67AVY9/3aBBP9o4dckCnN62AbqUnD4EY27pQfgoigL93myVs3OiBpsDr9gYrH5TXxevt7H
rsEGNZ0b9H+uQ+SZViBLlRrPELYX3b+AoBWnucYCcAefmIp2v3NW/2Y/3cavuzS6z6uhKgqBCq1Q
JFjbCEK8yv3B2fdfMga6usyBH5lEWtVZfol4metn7gFFJYRwL5vkrQzbKFndiCbf24Qs0dack0Lk
uXy0iZk1z6ZD6m6hDywD2amYDVaFguU/Xog9S54tsytfis/7BPVHML0ZSidmso0+tvU2pIrEPg5a
a0ds6sCGWnvnf8YrmlPnfNodfVyzRbVRxp5xVyrDEDzvOHqiY8vZhzd4L5TzOzoY0TPoQWvHxyCf
tBJJLk+QurWC95bQW/LlyfPACZSH72a2wmE/TFRCnW8Oq4qTrkIwt0Tp6Zln0I6wDPw4/YS8ToOp
YCp0Y7994JvBFwtq8BKLJSn4QxW8m8pBRDtWRAFR+dJP18SjEHsR2ha1H2u67TgNv/Vm2HyaM0TX
Bm+qxowzQo9QxMXBUdGihhvGr2DTYGkYOvvZT5O/d6uEU8lTNRY+uMLqw7WSLKd3ixJ7So30BjyV
YUeXbZMYqNM1DfI+4MDOFKOOyAtgWKMFjh610xtPporpRvyesHJAVK4SkLdMpDbrMxe7Exl1des9
KLtrTM3MhG7UBM+M+YufCle6RZ6L54hKDDoXW/HCwg02ja8cq6dwdH8BfDoDRv2yDPWnTWhwfPwE
R16jVFEfgr08wuR8WbXECIefE1qoE9q/kAgxnfw5p0Vti1206ylEakoV8QBVCP/a4v03nGvkG8Z6
NBgITO+2KysOMDNskkpXg1Ux4P71AmWmr5ZmiYuaC++qhS2hcq5SQYJVEa7kgi2cHVd+XGiNAux4
N/Zg8bT+1XGJMrm5I8UgJqq9HHMSZIrXFxb9YI5Tn7q/T5G6HLvAzsnQJ5yINUQ5llkmtlNvAwLC
jjV6zlvcX1aT2CnfntDrpBgirrfDlsYH2N7FUxCElLl7Sk/TgsXSUtu2aHTS4ZA4wKx2INlNBBHa
QCmBHJ/EFwj0cAg3O0z/ICPXdIYNTkHrTvdLlUf3fSwnMAUv60qJV85LN9fW27E4aTyhiti3Fd8T
2dNblpzGO51M6UFkU5ZGcm4FoGqqX5V/ep3THJ7AIl6tWETKGSaogXqcD/AVm0LclkTpEP3le1Az
UKDoqUJtdrYsmyW7CmSR/KMz6MvNdOgasI2bqHSiJo9LY0Z79vifxNO/qkDda63ww56Cv6zUO9nU
qHel0Juq5CPpp/4yLFSRw4WS5evzmrSmjbur05lVwz5huFY+1asgkhKlZazkr2210UeIVd4dAELc
fPKmBBOm5tTnWIXio3HNus2pGKitdaJYV4b3RrmgWxmMUpdr58CAMF/cEv1dKHZqGI6tbxdyCVRm
SKLYAaZKdQxQ+MnMJVHyvmqm2vGqM+rUWK7As473dF5SLUMWPVpSh3FvS9liMIgoB4c5ihj9MJBq
jL9bTgek0FweXo/E6srncRZmZoi3jlkFr/rQgjxRVh526mPRI6TDaoUMVRqx0fXodqjnS8VgtViO
p72b/Y/WPLtDolS2bM4rvQG1yeMLrwtpq05xM21hZL+QIJmOlCqq0pGw3Iaa+EhlUBm0ATZ/VCEA
UbUlBvOP4o6AH5h+V7wuL1Ivw504w7GS7+JVAIW8/Acc1/EgHju6C+gI6JcDWV6qlMODqP7XnuEY
UKeacBBuXhrlDPnv8AKSnAdsu06hwrk+AFIE5iXAIeZH9qCg8YpNsty+r15K6ybFSLdjfZddvrS2
NZ3q8G54cjwk+mvddp1KaKA3ifMxiZ/E/dBD0c8y1wlYWa77XqBmgv5h9YM9R5NdJKbwxSGwZ/2L
7hROyOAQmnyqb9Kmluo2AiEHQymCuAABfd3EBu2tcRXoE0Y68tDWrhIkbpEfg3zY9AGsfP8BDWIU
+FFHnHKZ04kabIelsFBGAnZD/i74V4djO1Qke4f2BHO51P8RN0E1eJlZMYV4f1YV60CRnr7cUyzC
tSCJGwZBmmTpBFsO+YJDEBECwLpmPKaioTuM+7WM9G4Tp6ee822Q49d6VgxvM+K8WoqWEYQWZzQ3
4HH4w/GjjpFhn1KRb5ML6NkRXKWfvCQwTmJxviL8ZQsKEa3vE8GQ21KGevAtbol/sZhEeUVYL3N2
XWHGsDrSiax2MUloRivmoD43Knw6kihF10T2XxJPbqerEnzqt5AWAhvkvN1uw+vY65TLB6aa0CRq
ZD9tYQ+HMTnBIsgflLeshOaUNzczMY4+TwyVFGVo2AQzGZRIpeYMK29PH2quPiRiVmOedqPsZnj/
oWAFMzQFy7zPXRo+EYAJtgLRIA+3x7k+D9GJC9Lauf6L6YV8BV/TF07H/BKxWxzKeZrmuWdfsnTq
xvnZymD/oW8cUCpZJZVCvPekA2xhIA0Mb5d7tQq3/fUN9mJLQxefKKfYg5a2UVRPDWSLmFZ4eNNp
JDlUc7FYokwU2PqFdzOa9oRoGx6iSTVVxIitIgyacwE0iN0WqqEc2eVNOkeMoLBGYRfxueYipEZS
n6yVcAsWB0SIYKhrDbvC0uEpKW6I0tLAch0uVsPDISXsv7uk9l6xf4lhxvL0/1DkCWmeVblw0m65
+NC01N2YPo8y0VYGu+t9uHkjXiWiRXld8jdmAD4+9nwdR7B2EJBjmaDnczbbaFfwZJuXgIVglcWQ
odioHIvwzAFADr3u06PjF5jnUJaBMj6ayV6V69CM83mD4IR3DcFy9YjZVFgZBHShBcb3iFC/j9Jv
cK7jCPQIJPwwyu8xsDjT/+UHkIJ/PUCJGdMJnT2clBQ96LL4b6z+5Dwv72e8caM+rVR/I3zg50lr
l5nb3xicbeE9h8lBBDGyGO4VcbW1uK490Ns+BTroI7UkqaSqHgsSfU20B+a2KbzSJBnQ/EL/K7Io
J5oWiZBvZnE8m8pbG4bVFgS/Ikj0H+0VL/1v42mUbYJ9PcM3TqZ+Nkdat8jihF1dd5cPiZ672moV
hwLh/aV1LTdecYwpNHFJ6wxe+bUBKu0kHAn3MOi8uFwzv7bBCEINEosOCprK3VTFEfIuWK0+gmNe
ISGuPx+HX003hDmk+SZLydoV3bR8C4gfNtSnOOhOfWb92gc/jXHg0pRfPiJmKJ6lFZE0bVcHhuCK
RypXemc92rBT6AmX+LxTUJygGZb2AfSxj5qck9O6edMrmdJiNpLCF8RxkDT4aWda8yI96i49Ibyh
M7JrFMlQSn7UQdjAOFXnetdIE0XUCRDm2571b6HhjKc65zTR40ACUkgISSDr+7V+C23Cwy/MJr38
uyr6rT/dJ8tPp4KQms3AOcnakTMhlXrOvN6MP5HHV0ocV1hMDhdmNisZvvlYmjQEt5b9Db5TKFXy
x5qrXiUUtHPMnZOtO2jYhtBModWqubajazssSOZSiUZTImP0Z+lkVNvlVPcvREM1yxchCzKXz2ZK
PB41xbH323kgYeWQgIKalomVLw6Q/XPzPAXAlrKz77zWb2DVQV4200Zcg4TXN7tukx1dzuMyMKa3
SQboJHRXPkfZ4MHUUcVAqia2oQ7HJ5va6BoAZ6n4z0+qZpR2+Ayy1HSzWMwV+C0JjXa9dB41ZWIR
ctQtTol8X+JTKRjhM02yuRU4x+W2pNjU7Ko6mudtFFKSp1gSaHd3BFo75E1pCNBYIgyr4Zi8PkvM
jWaoi57VchovXUecN4K9Cvziq5oGK/WZPJanN7hIUlWaI5FsLfgIyTPpaxDe62h4RE6Ru9Zd4Rv1
j210B5AEDhHdBiWTiyGrdpEK35akdiv805KeYPkk769Dg01fygicaBpsCc7dvxat0NvS3D+8lFFK
DphGQJS7AjhWMBtKiz3w+5UcEYlIMvCOD/G9DizwVwjnVAMmSaajSMepue8gdAwq7mMzBgTZaVWY
K3gIBQDLMT87aBcM1qwBXr7U4g9+GHhFwmtDkB1UeVFDa6fXFUN9z+cTPq3lkqmH7+vRdpefo3Na
tUbvbmq1cMRBKHwHG6fvZhQ3lbCJYzdhLF3xRobD4jrXmGoXIEEg+sHoYDpX2+/QQS6LwwyG3Tbo
22+hP0pN6RcNtP+LhsUpvZhr6ATzD3tb5nGWBOFNQTQYutZd0mktHTyLR+qehMNwAQKEO+diXxK1
t+uaY1gBRgdgw3zWJs9OsTbXe8DZ95jGbw/IgekhEn+Q28itNI/3FCsdVcuCk+wAWRrMQ3WN5OLe
8dy1zYCuxrk8ch0e2NAIfnD3lB+Lh/YMW45eJP7Fv2kppjpCji+N3BSLY/VnbfwKqwuG8Ow8a9RD
iyMjed79RXRwDhUAuyaqPQXow/WvMHOus3dlFlHSFTSx2H0dE/OdnxQ+1aJr2GgrweDWwMCchWQ2
fWfuRie5HfaOg7I0SObrT3Q1yt8vGbtMlNJly82UUko1388VbcQwSCmOsSFqVLi3anW7jfAjijvd
JceTp3QNSRUktxR8hVBKswltshVToeA5Vtj1uKGaj/uxTDz8d1B8wc+Ve0tdotRAiUOcdWTbF6FZ
fjs7ttn7aYXW5OJ/veALQiTLmZp3oToYZWX0aobYySpL/v3pArn8BloMk/hif37fXopBAPEYHQjW
fIK+ER1KHEKoN79grDgmagE9KBNI53O8LvrTbEzBbIIQ22FHy5SFQbPXVRn4bo9kKRn9/aifr2nz
zay7vkN3H5Zj8JSkDhBl+kLLqalnSkOV+WdwTJn0I1clmURa9EMROULigB8mK7/R9O/gkeFMv+/q
M4JQFSQ6Hkl2TkUMI4WSFHhHyYmETH1Aj6jidIv+8T1qSGw6vtqDnhy+6yK8DJB6y4nmehGgbVTK
qDK8sJ4pmTKQ/hkANA27nQrO6BOZ9yznqpkk3QxSS6uvPI61IWTCXyzKEn0srXoIECwV3RWkOkL5
vVifMh56pg24v/KPNOvOSo+iTvTmV3Tn72qf8ZyYaY17eToCtmpkn194Z3gWR+UJUpI/BP8jzjnv
L1C0kAeRt+dr0tgTPmDul079doFweys266GwhlzlFTjGvsOhBdZXvrmtOKPdf57d4kTwNKgm3MSx
BD/x5CtrqRW81TLxoQBM/nddJMwYfothjQxhLvHWhqe2xsX0NgceaI0lYbMTsBFQTr096/GgIdSY
JSKctIol+EPAMAQzobb4iekbQsuEGcmPnVJxyPSM6jTg+P1rn/xbeMtdig0jbxyKtMC7GbiNZNP0
wVhjre9tT8a1o4c+Gug/8SqNgLs1LmBURzl3wiPl4nb9nqAanPJHxOl1Wg3Nz80NZZfrYp1aZLQV
5nPeQkzWRfJReu+5MSBZE90fNz3749Wy9bf+yZMbWa80JNeakDBa0RK+nUBGyjkC/71hzSJts7an
MpHUqq76Vc3Ggr2sOK7qIZbA79cYxYe9e6B//EyUxPq10h1zt9Cms8EaxKxNAYEqujlTUuhi+chU
2XlrgOxaVe5dISIhSOp0uxyxPE9QdpjZmYHkk5z+PA38szDpwfzEv3NIWzCYf9nsclpGGBAwICgf
lKQyuJ0c5e+aQv3uzAC0lYRHkdmUAsSTwCkkqgdxiC/0fRJSXMG5LJQH8faxKXIGEbpPZAwqCEKN
Yg9Tdcqaz6k0VePnPwnLlf8dokyaVrxqYyuuyuH1ud2HwXSZdlR0C1+s3OaDGrR9uAp6gurj7o8L
grlT6zUgZiCCI8ns3nulwRbaegqWH10N6Uhf1lmsuR0M/isAnITNGK3oq7MizDVZVDCVTHs51DR9
HKXz7BVD3Yva7m2xxp6xXX183NRgZ1z/qT0cvnU56iP/P5Jh/quRIgqN5MU5VqlF9I3h3kXM6N4J
71b7xug71/h7f60OkTOnWb6slUFhvD+O51J2S844Azu9B6Lz0urs4Gi5+VErUQGnW5U/PGzIWWXw
Blsyum3JfP+ipOKRWEqUvpqTEX8HAbc36hJWtOupuQ70a1ikhKr+SHNTlMdOaYRlmEiN34wGxvxk
FHxqKlf/pJ2INk4xTAzKuxcuqpsdgp4Mnqq1UGMpxfkh//8Ung2ihgQGhAIGtA2I9787x4+cqZqG
DCgdbw+x/qPWwRfPh1f0tfrSR4Av6dID5S1/cQenMQsezHON1g44gvnkRv2f44jM4V2L5lS21R9u
Qztf5A15ORwhvnHfPeqf+4ewguNNnzg0J4NkIf+J/4sDEsA9bCYVfcImwn+eE9yqcPmT25xwtSUj
NA9FaKdFjHhei/8IcaXaBbHBJUIqrbAHmRb7+7As321rxhMaXs3AhWx4w0ZQqJA4XhwlNiWypnMU
xkC74ljgdmItOKWCsUOpcJnCJI7f8uRUZzDsxAPgigC0ED8yVKLuF+j0rXXD2ZmAScl6IMH7w2D+
jRfRB3gQOS0amKmykqHgteFh6KFIis/G6ny84QgWY+UdaOSFgnAdYNKNQssYRLloYFYta7dwNJuQ
jAI9mAekT4q+aMRmBC8eAfzcxfueqhl2AZuhgahjSndDannp1m9fmcclsTyYiLoi1JCEk96IOIKB
oD8/EjIZR481f1ogbF/r8mDTov65vlXtMl/t/l1c9gTcScz4cQPvped4YpEPd2UOQxoY1qcQMt4M
IybtxDM0+fvgICnelefjIlTJ7Fmj+ix018IN5u14B+uxJrErIzUmc2g4bMKL7ue2xtZgkqZ2wsne
OAisixAnmENdhA/RovC9OsD2vZXMEkxREiB0aqFXhIxxqmVIyy+M0AbTDpoZP2cI8tx04mKUAUaf
LymiQt1kXP/MQ3cdtXR+/EGg3CAjfkscAjXtL2cQ525g4hrM9iUEHW+/MV2WzkqMiVbpj3yerZVE
nwFCVYvBuUUWG2ExqedQ2BayrUIJGwEVbH4m/j5dVd6L6TFs9/aDMrq1xukCcSDF7fyh+51glq1+
NYgaDKK9LHJp+0JBcEznxOU9DczHhxsPg9SVL3OW+qxRBQKBVxOd8Y6CHv+dwIirD6uc2zK2oUUX
1rbosA91lXR3qsemORrzXuQ5TOfXIExNG7uKSJ2vow4r9jFwudTSLC761dKcSRy15Xf9McHMw7PH
Cwi81ksCcsnjFqZKp5L870xbvKH3hrOk6bsJ1ry/rP6IpZWw2E6pdH07LxhbhRoxRwC3laI63nbi
7s03oOWdTLJwd2+3ydRzarvKeDsCAafKQHiKV01AYY3pMZ5zmA7P2C2sz730X2H7xXBSHFw0ky17
adc1AI1RQ4ZU2TVxHaN5rKecs533/pdaXFw8ph3q3e9Vc2lSTHhz1ZGOakE3BFNUAuG4g46Zpi6E
Qf+Hqik4f4w7TaE8ISYcmj/ZymltDtkCuE+0EI4/VzY7OG1TsmrW2DB+i7CZulWBrqY3wUaOfNzH
d/uLgzdVGnoIKMuyDPhT14dQLPoFomoHT0pvHno+KAy8C/iVuPsD60pUo/3Ij3c1CSioWNw8gX3e
p4h/j6U1YoXsM/pc7qEsYU9nERbOlEhl8p/lEmSYYekNl0VF2FSfNQ1Drg8eEU4OY9u5fWqa+UdL
SVYBAReFQE8zhxBu3H9ppQBkMJsbtT3L9t5Vpf0CDhV4b1RH90MKx8J0wHvFGVogG90HKNvyFuw9
vXG0xwiYy/gQzR/a+ilnjU9qU5oP86cmP98xrsz81Cwt4jSNUUwVpcPdPjS5DnXdjdAqi2ErjPCU
VTDqvsWJUH7Y/KaGVE/vFFKl/IvFIbITwRiycbg2EK1qXbrZuAB55QR9xaMTcMDOCOuU41C/nNQQ
SAX3o9e5Zclw4pTDCZbEfrd69OMW6ECR9HS5jBytkDyXIyC68QurxjKujhj+DVsBgB0repRz5qy7
7+BlxsD9TkdtdVQuJbR4JTgoe/VOZcBbpZJJrq3bh7213pp4Nl4qu4yfixFJ6rkGUPSgxlSLTzdG
7xUBzQvy/meaPb+Qlx1YPc81Cbc5sbRlnd3hobszInquFU2F4i2Lx9/hWh9nABT8OZOQQJMn5uDO
B9vqVcZceuXBK7FqmTEyD8ig43LDXDQv80zlFpLtRPrWQGpTRVzMhC7MPdcKVu9s3iba730yGXte
rHj7P3yMDRDDKniOetdbf7TY3qdbT336AZxG6drYYczrSpk8Qlk+fL8DgbFcXcn0gOOhBx0SHdoD
9E8O2GyDjiY6LdTP93yAt+veodAutI4iSNExPNr0tpoPhFs35Js0mOkDak7TxCJVNcNbX2MsfMIz
GPmRAyQfMYh2fsYoKr7UpLLOvl359nLsQ/6gPj917lOfRm2s32qsbtRRtZYD2y1EJjFUb/8hEy1w
UMj9SAAh8VP7w+ytM4TGceAx7dgxoeZrkg4apSVLdob7DAhnnL5w+fbraWxwLmdy7qgD9jo+SW6X
Sw/p2i3VAwGOyS83p7y+w4zkdY4zqO0wpmBO00J333RBzNjMAetz/vjAdKBISXEg7eVDALADWwJK
y9rYGCfKJdK1UrsT+ZuOzSwGvsJ/u7UthgVP77sLOxWKq6bMWWtKo0ROM8F1U8Jy0YvSgboytrX8
jo7MZE5aekgt58C6CSmqBFG3NubK9lqx47UHFbbykAZ9PYgFEAfIC0gqgDLs5DeM8xSbER0Iuoaf
wKn2PqpbpvqXwYozMRwJyRQTDINpBkId8BqnlTqmBuz8BPBs2j5XJyban6rsZ2AlugZ7RHqz6yGZ
okcD+a/8wYZxHjiCSd5OLmHudYjixMeQaq79yeciJf+8mMZE5N5bozKx7+PN4rCKC4a20cac3QzL
zOR3PLRR8WsDL3VbO94BfU3RjyjWbOEPmJKyeaPYv67HBtReBnIXSFt8TtEz0vugSyUDH5OJAEJw
0i5J90vZBjId0GV5XqlhZCSYPnu6QAEW9njQhG6N9Ffkf93H44DVXb9x7o3Vb8XOP5b1ko3Hy+8t
92/+M7GVrzjUShgn0/DmQXTxp0uWlqJmRd3Y2AbPNoy5icYLzMlU5R5i1+d70Xi0cGRkM4oAmJKQ
qe96WUMl4rKNhXJJTdvRKk2PSKx6eUSkTlhPjv2Hr7OYEMr8eKXT5Ksbed1cNL1yXmhhOVs4HBVz
apjYGQQDL9+QI0uwL/ULdrsYnNS6NB9pKM59qNBOXrNRVYTlKSzxth0YwPqBQDIyhh4hpd1Q0A9s
utG70au9FcDe7hggeYmIoScc/2a8TuzSlnhIn+kjuHfsJjYhWsrI9LSQTqJVGD9++4V/w245d4Aj
49AHXY+a20VbpX0DPvbriXeLBElyynYqmEIGwNERhm6zZe8nK0e0wv5HpmqdJV/BzMyfHxmvMY/A
zbnsMc/gYCDh8J5zMDctUcXvobXqPQV+21t82Q2q8/vAghbMqUvSnCYQMt+6Afkw64fxp4nk5WMR
AKvMqe6hfPywo2h+LvyZCLLwVaN6GQrR8klWuirr29VOeYE32TCLXOQ9e9zs16taqakKoiA7e9yL
kEi1ngO2gQPaX2QhvwEvunU8bcRUJWEGZcjB2k0PTiEgsxgo78xl/XCfeGu5pynb6t+nsLGjkA5O
UY8ScMhVOgUFlGGVrJAqKNZEvVSK3QweTnjwa8oj2cONrCwarKMroQ+3O8a3akADJ/3pQjYbZIOO
WzdKKo+DzT0V83YzKqdb87wlCW/3giUkJEhX6bdfpisdJSiNSbZ2wVghZ9TLXjbRZzMKpXEBO8zj
hi6aQoGyT3U5oOTWgLJFSyOnJVD3GAnD+nitZrWrBZTjQi5b9rLt/6s5SCtIYycmKF5OAQg4TXad
jGGuG60JUWhappo9TT4vfuteNxlYBsK21sXR5hyMvpOjte2Ufqg+K62HpNjcj7arLeXrahjgjkha
lFz3I8xCyiHUC2Z41cFmWx5+V5+bWq3vusALbryrDpnBLu71zRLH/V3Z5HoBl55FMD53cdp9iu2N
nBaeq+THvVdrgX41qL25u9ue/BgfhdpRHUXZWeoif9TnwmJkKckKq4sFYuLQUPaTSmWLnLfTXvz0
e9FMPrP5CWMNcYJ87Tu8KNPErjrDngRPw3FICNGNKEM9ZH5qbdpxjsC2qzCdoID4ugZQKkP1AOMm
ddBtOhoGLhA+kFdvAoAUq4B6HuI+prCz99Sh7mawHV25kT6YKUeX/9MhJ1JltjOQoGwlkWr8rEmR
RH0iRf6ysXQMlhSbvaKH326Fpk3u72+WEtvWqYCGZw7ACkQbEzdLapV2Ug2LImzf/WTPoFk1Rpyt
KKOBWTE9KmiDsfpseODIeJf0U2bgwiQZvXre1QNW9tVmmjG7FoNk3k9vIXyyibG5hFciavEpT0kP
yyEnFLfryvRAxqUEerCLys12IUZVVXijSnK9ec9m09GltMb2n4ZHljBIvIPXt7xz16Rx8gYpDXk0
Bsb1pemgOvTyw3bPTZ05CiDdhaJ3GClXYMlrLI2WUjQ5c94tTzlyMGLn7wZgTCoQToeMq0J63l1v
VphBbclxzXbawteVr3IS2NbWqq1SdinQpZpid2vxK54wow8sKgjFO/jy5KAyyOCbxZ0dni5tfmAk
SFHP3QElOtbMFb8QowA/HhWIl/4hrFjHcJpEp7jthFxAoOlra5VhYscyjosCvN0dVRHhmtIH5cIV
H00NTokM73QBrTcs3rRgNzGov5QcPwF3CNltIbnVIFePLA3UIDLch00ZeqSudj4mMbbsZPDJhXCu
1E0cQBIGwXnebjXWheihUrX1bYz5La9FUo+uHt0Kj9q0pgf2Cl79dIFsgV+g69PtW+JiYdK4XL0C
n3A+ofW3KC6TL8kRFAMRjdwTHdBf1OIsPHZJY8UEeglZnpHYrMYpKeOtHKSodpkhQYxu4e5NVQFK
+z/zm/CbTKI5nHP3Z5lprh2JaUnTEZJH1LJlzoCuMsvoFfuUsV6LX/9SofhXuNrhkSD5SSrRwDw/
eIzTzmgrl3gUFz/KAf/yA8tvM2RrUojfzAD58hnycMqjWkv7o5JGNOH1kncGGQ+DACwonySECbmH
xrMPyzMqThsLYBAPcSNf0tYaIIu98skbSv02wRCphI+TACv+YCkKWcBvcQPoh/o9L+Hcyqev7FuB
htdoB45K662xCP6ZNWGMo3HMYc8mVVs2s/ZOlYBwFYJeHk8lMG1gVDdUu6GIBXBUnP4w1UNbJhLZ
WqZZhvfZhd6e/ybkYqe/dwjpaw0Vx+dgLrGg9eEz0zKytAXOVQJ5dv/+XuzcEFJSg03mEpBcksIw
QSTqzEtNgsi++5VIdT2/vORJbpAdRRThE0nGjhljBM9oX61iMnfYn4cdLTE7Le3xPMeEQpT9BXFv
+PuS7vkE+QojR4pa6GmIJr8RBAAq0WoCL09NqwEXAxcQdcBqewtAUkGhELyWl1j+jpbCJDznzke9
qeVgAUrHZgMGfETcxZyW3KB504U24pY53l+ZNCGBpCIaWYPJJ7HBcg7Uzw7sh1qrJPt85ch9leei
86Vbx7a3cFLaJM33Jppw0C8qJkIf6B6pzn+77ip7YA5QPpJ23ttkdvzBgoQbNE9PX1fF73IQNCg4
oeukRnhdp5+XfcxRyheimvCweyPXYMk6oeT5pXLOT/qwwsESME0fVtK4AxFhZeyY36bkV6p0QjU8
MrVa/OIquHcS7Xc8pvTcA9h1SKudA58CfJ5zSJsRsExk4Gd5NIVEaotGOWWLoxfvM2F/9OJUMv2Q
GFoG/wD+HMtPhnmDe/4xoheM6EE0Rup034zVSLLK7NB2OJwMb4BDA/+gA+b/sIRQeRQZmnLhWHmq
G3vHa5H9JNFCJu4XpUwYkxp80YCVjtdJT6eXUQj1AYNlwnZdnXEM2XB0ALiHXe0RIiDZ4nAEA5AU
b6gzEylCA+wXPks8CZOFqGZLX4TxcLFw0vKlEKfKIlgvbPRWIvHYEWedPcDbZ02xgJUivWHY0mPw
OXKU5JuODZJVr50pJqBFseJ+kh8C+fMcXt2fhQtV960eGnbQnL9ZkZYFC32QELTgpD79NrEj4n7I
l7Mhwb9s6fCDWlt+iVhFbv8eAJJ6RyaI7zxXjL3zzuBP+489Bhme1PuvgJNbwwFwTpyvx96Xp+f4
h9/CzlIQc03DtJ+yCjQk/qKiXZRdLfurWogqXRMCw+4Kbdtzsq79VoAWH9O6C+sttSiIDF0hmBKQ
72ZcP/5H1QIkNLVxq8+RJIMsBR4xYxebtsgCvDZTYpwHRBf/bGBy9zsmF1OfIwIvmREEDSmtP/p9
sBSYvAvTUJz05Lnik99mOJfY0CK2rvi8fQ8HLiWCBipVNC4RCMNg5aXndS30M/fYS2LoTfQgJHVO
PnRPZWZmXkJbCL+KpCsr2/W/67jcWNc4ZVxB8VqhyrFftQkntqct3UY73UdUd1T3kUsTLJMqu3Ij
n8HCPO9LpWu1PJa1lNPy5OPlo2k5W2UUlfLaniV3kH7ptPG2zR5AVp/53lxjiXwhi0iblQmDiTEA
R4bakTHfqk6X8SzO95MnPrpC+BXBivGObmlMav8Syq+0OTpv46kJcL2BErky8cpXU4OEa+c01ZAH
Qm8rmgUT5nORsfCt0muAJJH9zIjp2iZwh0JWN0zEd3WDqXhgJAzyz6Vnof0j6/y4WK4eh8lDcg/Q
kbpBWO0PYiJTm/I8NUsT+6msy/wV9GeObOfJRBgGWQkwbtyWLN4H0LvvILg6ee2OIWYsycjBx68L
i7f2FtsImWlzUChc0QMC4OrgfYviqmqNRNmCv8qypZaV1QBlvCH2KiZITz6oKT1MdnnhKNgyVZk6
uGyzzpzSTWAWEjU9mLPjB4OP67Q81uJofdlCldcsTdiCl4gHALPPHpcZvNBTNl+pevzkqAeR2thn
T5ZY6fP4Pexxx43EO+x1jdkD3K/eIOBuIBFgI988Q7F920x6WaHp821VxSnzpHQcpb1C/FcPA0sw
ldKawhq7aYYVajHUm0Xlgef/uilLqpLZyCNZlPakCSXsfaVnxcV2d08mlZC+Y0wmGDI5vkDehEzF
nr7yPGpgbQ+m/B74+CADoud/IVq5mrzZHeZDb7I0+mzzdKLkkm67ums/Ra7K1Ykpo+rNGjdeBx5n
2WB5Jw7ZqZWiGCdVENCRfO8LP3MyiWjcx7+iImBZp7tGp/WOxTWWvtcKfIZfSZcL6LzVnrboxADc
CK4rN82NdeoP4zQgIVW0+VuytafKV4nzY1IOvQOHGDrdcR2pSd4rKT5blkbJyUs+9Hn6GtyxCvxp
UAepe6Tf2MeYXgBGRZ6CPjq6Je0fBbnJY7V4bI0Ekzr7Ibtnepax/TvYczFhOackFGzteevTLZRN
wgWT4NN2GYkR5mowvquAneoUlDz2Aj88QSTdMkNH2870g3qaVVX3GMIn/EodPM04KBJOwIa0wLim
04BjrwBl/gaNt1DmpCExmBV22ijPluyE3SoCQLs9K1KiGT1cIa6p6Z5ujOaYBZenTgP3C3Gpyuxa
G7S8kwW4YUKoPhwfJTclFf2YI+O5xM/q0q2mhfqPnQDMPhzwQdSms6Yb583+e4O939R30ulPpXlP
8LXj6WKCuInt8p72J7roKEo7Ueqzles6OWWpVJLEe6F0FtkQmbrBXiWs5yern8uLeNT0vt7yRCcC
Qc83r8GT5SL3n1ZGuc7u1YbZstVS9kcvQT7d21XtoUb93hO7iBqL9+XNt8sGOyjbScH9lAPay2Oz
UoumwDxCncIk93Ad/Yxo23bLWXKYF4c9nVwCGb4Q32azEx2mPsv0x5jpYRux+6HBWl+UMDvDHj6T
dDn0GGmwjceTIPn6Eol8ptTQ/Mgcpb0BHB3ulrdT7IjAzXnqzxIhqeD5JE2l85gjlDLeKbS1U6UB
1yvBmgy7bNrS3PW9YYuw1xcErkIbdV9/m0872Xko51tV9oIeTClyOm2Cy/Skl7UVIo7x2tzB8NAW
Zzja/e7Msb62c1LP/DEfiUrCTdMgVQiPE+qZsAksyqC/xO2Kapjbx5ZQTi6ER6UQRMHYblfkiGtV
4pHUFey7QRVlWx5pj9TPp7I3Z5ML5j3x/8Vn6CGvmx8LgIH046ilrAEpxplZJs1JhC4N48JxFYu0
kFx07F2I9m5mEexizsRbEHR2K6052PZobjU6mJjSLTP5VkWwgu2Rok2ozTwQxR6v8VTwcY06JrNU
5iJSfDRJ3CKR7dEHW37Uo2TzGVZ3XRiTwjfNMEfg+qJ2zbDOXVECunnxs1M2hi3CXPe54EbPIgfV
IxxQoUc6dTtYBduHIVlPyNzYY55jDcsnm1t4r6rT0WEeIjOD+lnf3x308WiGKkSdkCTCXAgfQT4u
kQsOxCFSsnp24VsITLbZsUZC5RwrczBzAo9VBZq0N6ZD9ESeu6yETetAGuMTUG8A4kpggeX8nyq+
bmNdzYAIpNlKDsTYfqGJcAq6knqhd+kmiggfdZlNGyf+e+aKrhJ0eHBp8xhxkSwRWQtAK4gS5HFL
0IwaPq1ZzoXwwVQi56Jy4s7ICWBcnDRs4uM3l7qg92X4bcrvlfiEc2dR8tk2DC9QXK0lLO3fqo7T
7G8nTMs6ps9klyph+RRNctehm/yX0jnV/DubFDQXHwE5HE0Kt9NmI9W71VZaVSqKdAAUcutTXFA4
4c/D5VmQJgyYGfB49vWvRsi5fL4/RdQw75m5sKc7QluB29IATxZU+6GE+ZWtDPbH61RjJ5I9kfkU
H+F4692Ha1g3bCGhfVeTkaGtL/uF/r64GZW/mAhfBSjpF9+wRDjIE+rd76hQfMAn34GOjkafPw/D
xnf9Vf8OF5ChE7sA+JWGlxJoR9eNTqsEfLZl7EWOgZvU4jiFNQuw1Xz2wwrZ5jgmp0gUzFUqqEln
zX/ED/wNMtkBq3Oak5A8idM2f7B/l2ggwJFCYL3eH3pWlU+7x2whhaqzvKtKCWTgo0vv8qU4K83q
PohI3Lh3VCVgy90ilEwCyWC3gYoFEb3KfeftF2VA1obD39o2qzIWK1Muh0dKXcaPH2HK5XLmd1Nb
YzkHAiaoLa7M4I0JmDlEgjU28BNEdSGwLyi0JW7pOje1h+zurXw3mO+/syBwF9aOp/8iGiBLzQS0
pCARRTNAPWUPshVB6107+CI4tz/J8iLshodCz/WeTdztNWEHST58KJ7orB2Pmow8HUIIeeet+4AK
UUG0mlH6r+EqKZg/o+e6YoqfaZGl+yndZNojKkWW5g59E8/GGBRTT/arJsBypiLpKWhFke16rPbx
aFBDYNdTtNWZtd3QNnogVO+x5KYyFG8VvJau+pzWw1maaYFUF0Psaa21vVQiooslMnFmMew31ugo
jPqGnyxPR/43hU6fJmVQ+14cZcYrAbVQTmFbCJ51HVcgqvN0zRO0mldp7q1h68GDDXOQOuve7bzi
j2jFdL1qAza8myK+UIOVg/q5EhfugB+7hTNF6d3Qjr5V33ZVfrl9vaSgwz7zywrBamBtMnaxajmJ
PLx7dKuQKDefeZZ5JQ3uzTH+VG10iKCkYIhK/L9wQGbveDVcm6h/Ok4yojZc4G5TH+Vv2/lrFdiC
V7wEZ+Gek+HuSDYs56BiS1JhgGjFFrIOdZcuNK8KsboYEUaIdADE9Jegn5Y30O3H5KThRI4l8L9t
qqo1U2KhH6Wt9kdYIUZWd04wMlUQo65gTkIW/fHmp/6FN0HQRF4RJEohHgMFY/HqFIEQwPA5x0QX
vBM0hvBvIyG9/oxdwF7Sa3XvboFVanJNnX/Xmj/AvYudw61hrPsZ9/d0Cc1p27L2AEBYU2QA01dJ
l8Pmmhpt44VYeXtbCMJMtRe0tQChA+ThJuim8lLLAJntZlTe8HZTlanBjgHChRwCUyE/ins1hp3e
PBeVY28XF1e8nuROURZUlp+iQC4sb9uum3UEuqi/57lAGt3Wjfl8/TP1P6I/Nu87tx2WDU4bBSyl
KdNpdRMHWhNX6tb3wcfroKTYG8eFZT1IVuCYbBoAzWMJ3esQ2ZDLQeC+HpISOXNZBpcNrNVKQKVG
sUgjmNeQo0P4dscJ1LUXHqbrINP1q4+zoaovqw5zpeA3C0S+KKxup6vVBDHmsakhdxCxzXoYR+AA
TH9ldVAODmNQ94Viy/vAHkvW6RNAo4E9ygofLP+t3217Y2i3UCQPfsZr8nALrDXF4/7vn7yxwN40
U0D1zt4MrCwgLi503SZKMr81yFSDvGIbT20epP27EP6D/E459tfDLdFwnkvb+HV4AK/70MRHS3Ph
16FliK2FO7QPTT8ytH3RfdBOZ3Pu3nZ3foTg3rTHRlKjXckGGLRlWY7tYarZ/TAM2idbPK5ajTbY
X+EIC2t1N2Rln8TGFQL5eC5eknyHx19rQ8UyphXxnsiHvM1LaLjh8YTjSeKETvjVCmxUot35d73w
KjulJB7hvRlKUCuRBLndP0QO/pmcFEOHIHJb3dVu7oQ8YYzaUTiconJWuQ1whmt+P3P+cW7UTN8h
QPasjyil1Co1Nl7wQrhxsVD6fg1hjhvQMMSpeUAh/av0LdfX8tNFHZCw3XI+RnfLV7sO4J5RYSF3
nE/acjRCsb22kaGvokZXGIVC4ETsrBAzYHxtXp5PsiD5mGqdIO3cpBY5uuo5dE+Yo+XLRME0a6h7
6paLeU4adFS+shztERDB37CWSJrZSK6nsJ9IeyZmf89tmpceUL4x/Dz926Y85HT8nSreX1lbPlWA
0I4/2VXUa7+ecD4zr754dTmn3W33v6AQvbnZv8I2NLA+yjBiQGFaxzGo3g2LrGp9idcOYuKHO03O
npphV5TUrr3A56mZOeJ1YiWsxDq4PGJy6l0H38vxpZU8UjUpJ6YMgrbniJLyHO634ra0r18lc+xK
cSsaWUXojz34wBKu9DnKIY6ZkcdPEfhY5JnqNaSpRNYogJW6txCAIxl4hxpHYtltwlGh06s2BiGi
8VFmFvIkV6MPKvqNQm9w3Afh6D3cNbdO/BTp70dJOzqt/C8TVp4ik2S401abFSJ+dJhrDqKcB+UI
6oH7u6Cd75fWn7EPGzr98ZrZCEmtVEBpQ31PE/ryQygYiIna6BILqeU8aZ2etUYMFc1ClePCO1sf
moqWaB67zHQdLMaXetVR2cLacsdhgfLEb8hEU314QgRdPsmFgKp06Amkj/iuK3qmyWl/3/PiM5Ol
9Bd6qCJvgAJMaKndDtnogNHvTsbxI+wVnlEvIVkClM55a9uSZUlbbLEkCqEbr03LxXisN/tumrqH
n03ycPDcUQC4H+0ka9Y1J2uCbo2i3X1OE6E5S2w3FjqLDcd//boSFaFTw4VmEz6tw45JDXyeTp6a
SGepyFbJDV73dTy5eTXDniB6S7NgOn1Dg8EScZa6TE5SJUN8RuqpgbXYjv+LQ+6WuQL4M4GUAgc/
0MHHeM6dkwisoq12Atd8QdotztkpOrNdn9yH3s01W+sYA1ZtlWVuJTPzNBgYViBFqm3uIK2JVcvk
mPL68doyboI0IjMm7OMpduDL7OXbnDabrVbllSLfnOr7nEyj8Oe6ReNENA7ksIQi8vXcsbUnkaLj
qb1EV1FluoA24ppzvW0DRkc4UNJeL/vMPxIbXFuDD9xnK4t4BoIdUkND5PQfaYuE7o/+XWzULj+6
A5WUmaBXkTTpsmLYfv8zrLFUqC+uOMUXuo3xdd+QUryz5+qYDO5PG9Th4lJpmJCrTlfk58JY+eSM
6gcLGCWaq+XpBtM3A+tdQoOvZtk8Q98a/plRIyIAtaxpBOgn1wznLzr+lDXheLbhPOsig9cMI0mw
5tlzzpX/XQ8nzKy/VvbF+9AGog5hA074L+RWM5Ixc/qPIwQcT057yXNfzb5FCCJjACZJhpOtqDQ8
gsHoV89Lg1Yx2siuQIC3iPIFbPzp4n35YxextK25k+ioSwbp8DldvcAlNLEpGSoXIYskhigYtkQK
28fzOdl3NXRuo2pjsbvJW5ma5ETk3ZwqMVeYVNaM/1KtZ82yty9XnYAGslyg6Knsl/U3OUb2LS54
mw5bSegBIm4my2R6sf46h528ZWBgCqGYEBpxT5rOndSPGO7cJ5a0J/+jv7Y7cHvTPkFUJ/igbSWa
mrfEUCGcisIhGMI8nHsF758ifothkueP31xD+UmOQhSN+LZYBwTm1WK31+ajNfXR/8l+9SLH+sO/
92UzwA1gzhnxjlNRBkLlpusu5lNarXoCDhUsYyXtPVzqhIvr1S5cRyEzPmn0AE0C9U1pUNT+HjCH
+5Du1Ms1oOuemdfVEUabtjGRXm3zSE4l2OmLFaJiNabFcuDLBB2xcEkKHottNIiB4WEYXMcXSuJ2
7TirqlOWgvq1h3SSjBBbRqY4tG0LO70LQjZUy+5ZcR6YPcW55RO0BY39SXH5lAb6COJ26uZDiaXr
o1PQxan3WaBSIjIXPrQEDDQoSbYoG15EG1aNIUysyTeqeuLwNDk8y1bJjuyu5oBFf9afFxZ2jrsg
Wyvd21IU0xLN0pffbdYq5qN+hwgWKkRgEGaV5QTjgwWZbTwIZj1xFLZDTEa0hh4wTgUdNKdvKHZC
GBFzlywtUujh3eMpeidPRZSB3mCDsAlWRcWzAvL3PGzvpdEWfTvxJsjfBZUIQMzvULsJPfI/tDwk
tjzWVXo98ohM/7QttgO8Kk/O+RmPl0cbhPLhYXM12LReskWvRHgdGUCvEYCJIJ1uY6TL8iOSyikN
XifXMPewIHh5Xls369yvC18SGPdH9DxeH+tRbiDEMQqowIgBSWRGqazkA6tS1qXI9EVrXBUmqw4S
VKz0KPEfSD2Wdr+4V9fm/mg7MXhRMEb/Za2M+Pkz/VmeGlnzIVTFnLs75YWYwmTYlAYgVBK02oqR
uv+BCphU1ALohSMlvzyh4ijyLT7i+1P61NtJtP5wh5BvtEEgbnllPA3yRXoHLYP5B5yHK52UGvE0
sxX+Biw9RswQJmcrUE+Ut3vD6dC/ODKmYaPeig9qWwSTasDW1XKxY2JIVLCKndhM40YsEbDkA7J+
sHEzja/CWsrqgtPl1NonIoFIyZGpvHWjMEaVndYJRPrjVJYqEKmgb4Hz2TXdUe3wwqP+oc2H5xoj
W+JOxzmVQb7co4hW7Sci+aVd69yIRL2DfKNbuJNNvqt8u3hJKmWv9dZOs0X3vClWcWQjTsWj0YCV
l4rRKIeNrBpeG6uYYvIJ1hsGgeoxyP0ylzqKFspdlJXnlhZ8pd34eVvuKwCH56VFtIRr6SNy3Nbh
xy56R8DUzAxXnKoe5cHU8LaeMenuuU6sN1qsebegcZtyYIxeV2SwpnWaZ70MkxpCpaK3JpHdrtjt
2y7ARwtL5HeDRPo1XXNR5uehnB79Ld+c72r3JtPLZCl984fw8PWK/TqIxlco0Yi6eeikoK1ZbQgF
cNHj0tnNH8eQ9uXiOBPt7+tQd3xYsnqTnMKco+YjfsN4tQhUb1weEMyj7kUxA78ZPVxPvmPhNcz3
S5AebWGm4fxAwZ/S0E7DQRf6LJamleqnW83jMHhpG/suNeyFLr010vssNrYI1VQZU38whLee55nP
Bxl2C7FcrB6+K7oVr6iGsSTHTql0w6FqbDSD3OjQPcRpDKoU4xEu15HRCKEdLbzu0ppFWOwQoQX2
UAXmaxFxyJiQdPbGpr94EjKgQtKf7n3DDE3JCAX0JaeyJDBcELq/jXP7Zg1DkQMhGtcriOExqBIm
aIwkIlzK9FkOXtTPCuIhWvC/QEVkJjR1OmpJbP89CSCeaRzgdjNHwjMq2OlUDON6i7+b3/SGkGnt
1dy8Ho9WPA/s90+fq5LbvYGEEqbz8tlAzQiNE03cN92HwevVfgh7b+SIpkgz41GyqyfNEI77t0A0
6QuKEP/tsdXXwGvP2tpJDogT1jDNcMAZR23ajcgetE/z6vrN/rwFAvXRkBvMrrSjMKH9Z0FvKOzH
qKikdVNyhqvV3rcDVSinnUKEldZfmX+FUSaHhHUerkBzb9ewimxGKlypTs4EIAjwBymBNtIm6wcK
sAv3mVoyA4smeIycgXFYt5APlkrJMPYr5/jIrWekH6d9oIaUP3wXfkqAG4VnZLGP9QWBlYQMfVtN
gsUFvV2erIi8Wn/bMxhLO8XMaSREwYHTW71QGELl+n3uNnlSJzDDkwnpLGJ3VM/xJZhrmjwRc+wf
H0yNelFmXSk55kpa/HOo5ygrMpcoJke3yb3PcMUzLVRvpJ/4F3pZxXBhI7ZiEXWoXd7EL6Z8vXxu
yZsKX2N+5yecA/7G3Gd5hrEi6vdH+8/4E2n6c0wr2otaHoT6rGIn25ZQtzQg0msjNbmJlnbANHaf
g5Urcl2Q0Hnheck9K1phGs49LX+gEUfyR31LdQeS6gXHdQ7yN67ULLlTqtEOLRQGs2UO8gqXFmFV
XZmxBIrO+4ulLsuoXbHCOR57B5Nl1+zGnG2Dp7TBVoHVOSQBZALG/CXIBvta9+iUJVYnqs9jEU74
pJlqg0MBWLmixJMVje20xzlNkG0IN5QISzXoaya3nnR+rmVCLZXQqoCWU8dEIxyhhQXM+mlhJyjW
7v1NjE9o706pMbLfW7p+j5DPEplJFvhRCG9ykjFMhjdqajXTC4UxFcyGqj7JHF98yeR0JZbRNRLn
HW6CIbnwzmCH0oWYhHPAZ+C8AsAr9+4I5SbGfwP/58QFybvUwq6e2A3FPDNhKIHDQBGTQJLCnKYf
2z7PGqmp2jXu91JmmKrQMb2yiTPfpYO5XITxBAkmQnVGZbTEa1nKFSl2RTl1JJ98q7bDJYZcE1Ft
NFZiFDxt7BQ/loJ1QfiUSZAi/Scyy0d5yehRjXuS2RbovcvIIBdXQt9CwlIyYGkeIStf2T7ndac6
9QE7J3Ega5/H1qF1IVsVRBYejY6owe8rG09AxDT5tvZ2Txv5j0BTvdaKrqoTsKNPE1Mf9sWWQOhZ
KGOepeo+jpQyjkzdXer2olKNE5NBGsRMR9js+s2vi36S1SHzjQw4tROL+ESZhsL7JnCVm4FV6AQ/
MXMMhWZ4JXXn1muKcaF8Ct1kKZb9zkke3xyWzz1Dx5EkAp3caViOKzSEwcskEtL1KazT1eCwESca
sNpifV9EVnmWxmrVeRPvGT/aLI9m9lJUA0uFXRrZxAjnvDCOuIGYgE7OwdwegWJz7T02vK0St27c
JGK0rImYyTI6yrXlb89cq7MlVVpF+34WxTn47rjD3cFqmKiznlI04820ATQQiHrUqnYfwGOnNUF8
YjRCW+HYMLgPLKpm2kSz6iBCWmgu60G/YGcrU8peEj+AsOzjWbEagqY/rQT4yrLKciiwqLTRn/0S
sF2awBlLlxY3UQqA8Hwq0okQcHuy9fibZF+7Wjtd3RLA3k7V+Rb3XheB+HM6LRPXKNii77LmhK4k
1TRqxZ5+8RXtSUiJy+JdWxwfD/wHONZczVifKcvSGVeeTQ18ahmCG/6gD7mOpt6SlVeWqsvUToRE
QzzJIJDUdCPKbgECSPvurGRKS/mK5+zm7YiAPdLSVLDdxsjcJ1K0lFmcxx0Wnun03em4jd5LXQRL
XW81SWp1kbai5SbADc9gZiWsvlH3wcgvBY6bEOvQMNdofZBd+Ug/T3ZLzb9qZOtmPelxlK/7FGo+
kAP3n7/5i5i6hddi4qgRkE8aq2WiSHi6EQWZrNk3FvPY+14dbP3NHsutwSmRY60Vj/iQdlUp6b5c
C7lHj9Zlxcsl5t0UIhZgDTXa1F0iqivgnAm2XjaEWUHIKbzILxAPyAeUTpoOZzoejT453ryu8Of2
TicE4mjOF+VDbuJkTV9+smpZb1qsepyLqMO2w6FFzleKp3/RbXIL5w15RWvAyComcLMHU79YFP/a
6xRfv0PxDxajkcLT+eKjJ84K5jseohcDLL0BY1D8DCqTfhnh4cjpFMtqLABFPXKyTZ3rDBNoKOqR
/S/N33Ok9MSQj1ISCuiJO3lHOTtFn9Xp2EAlOhjhQyeEOx+5+Hi/iwTaE9NeDaYPuimxy7wQ0/Td
zt67RwzzGG/w6/EPHLSoGmhTtQpoB7l5vWn65F8wP3cl51ZKHuifa+pnvXn1d5PQ8+TmajcftnHX
HBzKbLEm3prjW7DKZAx5nRRdv60nvd8eGZL43IUgL67YgsrnSi2AMqVuxuBddaTc2mRc1XK68+ig
TRg/bfBRek98u70M4YWwM5KeB4mL44sVJax3sPUv1L/ZrP0XAVUIFdeOB3C/y6g9+mmqr946mLXJ
o47veoPEU/ifRBidEwm7nZklu1H73HLaiM0JUe5TiTxxKH8yUDE03/4P50Q5PXeCyEk70qkx96re
Y3uhIfhYsMLHHCmPadwp4O0rR6GMuaBBitegj8swq3Yd3kp0md+89QNDxvCvJET+oEFq9wRLn2v8
1leLHNQVvphIeKKPGlhMaTv9vw00yF2io/fUNQM0vbk2jXiu731+ddFQ5tYgI5MC+BztckNeXeq/
+vcrRNQCuZGLUPAkALnJe/XtTL9RgRRp3gkTFaJ/esKaAkbwoCF3J5kb1W8nzqZt9crND0hn4dBu
SRh3i+JSL1JhLNWnBENxsMa3jOqVsMFUlNzAzhI4cpROsJyfNVoAXTkIlM4MYYj0Yo7YzG1yCwOR
6owTwNER+7s1raQ5iZn8s1wILqlTysSJd9DV/h3kGJD5okjN3adoqpUx+7qaAsonYXQSFpMGmp2V
3n8a7IGJqyrxvA7U6vIaEhU0D29+hhw6mM1Bvt36pGrOIK/paB9eJpmnGua37jM/Ib5lo/AUPaPX
bBy7mIO+jPXZkleIxPZK6poF4a9ikmuXPVI0iEQmCm2HD5aR8JnaTp6xhex2F9KfFRRmOxHAuOBM
KEkJhVO9pK03toYzgJdnZMjhHkGjO6UucCRrBqwhyuDApJrcOLsDpi9TgjRx11wDsjqIVrMa6Fi8
V346K6pGdjZ+XoX4c6ErAd3yzr+SI1Ps/aEoOpNfQIG4PfeMcZHlZyJGODPxa2bx/KEJWSl/nMZq
y2infzi5Qj63/i3sG+JBeDjeGW9Z+Ci0ti/OPNQra3x0Z89AQUVVbtRdstBfsJEGS3RRNwaesE3a
GZhfiwBPVrVLx0gGhDOygFnBEFUYGxQuqA+Te0OXo1OjYkARADP0+oVRdh2e+N4zdQ1kMrYxblx4
6JcIk39z9vq35KZcYGsI1hSSBOODIT6jvEL5nVJs6HyndZzQtAVg9PO5j6ed/Ju6okKpFm9CZPYo
kAYv7twSS/jec9IuOBPpCCkX1mJbe9EkT2zpPSz42elR1JDKO+trfLHf01tgwi+RTMi0UIkR3J72
Sfvj/UhW4NHJtlY+KzEANzY/AO+lDevJKvnz7eREGmL8gzs8Yu4OElm5rT/5Os6xxD/b3lSFcZn6
jk+GXgNJaeToqYSq8AqSqG0qWTycZzXr2SNsOMFd1ILOEh7FJ8luY4fQQcrRCiPu7LlRaJxooML9
K/bvFMfnxULAOk6F66hYgfdoxD6HU6LUiQWDKtTSQZ2AynCEVqFJ+PS22FbpXJOaiL5fAxcNUqs5
lDErrh2V9vusplYzNc7KFeySkn1DmMSzsQwEiNU9Ns/vPZraNary5b6k1sz+OTY0cOEB0qyJTAZo
dLMs3puC6ntued4Ql9ILavrV3PayBSBT3w9W19/baERaKLFOu511nI4af361XDVX9DI9duwPh0Uo
ItAzvWTYddSVlULGYjnzguD120gW1DpIARJvRZXIwi9YXr2PavcXdt30EGMCo8a5NAc/TwwKhHsI
CenwODqLSmBm3Es3RLuYqwJi5HqVYddmImRgmd82a6glxjjnNgfj53finGftx5RnKMDSgqj8ZSUR
tjWeHEW4iVuLGt+/a0QJgwhDTc/lKUJ3I9kicsWeGEDphgah8o1I8WnFOQeJBmVi18xznfJFAAyR
KMkH4aj0zg67OCPHQBzU7m36Vfb/ge1DxBEfSC0uqtc4eemSgtaw8B+fcRIZ0/E4LPQnPG9wxYlH
Ytd4HZy7q1TtcnUBW5ZDUEyWJ5ao70tRWP9gDzGnxYuTVYrSs4hpjIjLyY2hLtX7Odi6CLZs3H2u
FKTV0ZHpHt7FTQtjPz6DXdo/ZzOV9so1f9ctjJcRtebfpAGYgkK+e2Y9mQgGH45SkhPQy/VU7SB1
RsV+KoULAAtu10J0clVNzNx7spNR0EVraW4E1OfbyMtemhi8BeZdE0dgkCSY9ekD280T62Scsppb
F4Rg2ITHp0RwvO7Dl2vBqhJW+1fsh+gAcnaGy/5bW/ZR43heXFN1J34i77vEyF7QfPwm6jdzI+KZ
VaZUtF4X8zj3cZDEfzoChb2Kq2/CqnajIwDl3+EDMlcCwsGj9tBOC491seei7Cl5kWPDP4GkP/HJ
maScK4Uch4FdSxNGOFuJ2lEXnsG+SaCTj/V/tTt5MZ2tOzKREfD/iUjeIpFaueGmA5itEyHUKRL3
yd1aX/XYbIOYIKEjTTtr0vGJo2qkStr0ftQ2NH6EqGOiED4Z/God2qYEVc2hLShQEBiTfYG4LMc6
Qw9LYxjMY6TROjhXlhWgWwC+cxVkiAcruGw/4kmh0i2hoo9f6L5xTBv1vbhFwNOdzaD4H4ci72uJ
sOZAFuMzMVHl53iLehaGaXbPKkC7cMgnYQs+/Wan05dgJ/rUvFcTUOEEPn96GttdGN0Ks1KOByzz
4aPj0DL/vwcbRdYs72uw4OE0X8RNiP2yPN1jZdq9/9qij71toMOLM+jJuScMO1XkO7fFPDNU5ssy
9voad5ryThV68f+gHXgUjGp9HG0vk4c1yOMHoUs2hdPRY2V1VL4rAa9PvdrrvxMtZszuLvwuH9dq
gbYeeLYNdUgLxdrI4p+8PmSkmcyH8hyknyc/LRardjVNgbd87Srdgmpd4Jx5Vf7ui2IslO+7Waso
w3I6I29xqe51ERjLEuThsKq4FAyFZJMgZz5rF2SDkoktjoxHxsjAUiD82ifACjdz0h9/ixkCHpjB
bzQ/JbcLP/P1nMRQFeGrThywtU7/C/Ch1VmCQmu2aCzbYdkEDU64iqW+aTytsdK9jc1oKmxjG0Ji
sSYi4agwBy4HbmabL6VG69x5Wb29QA/PjS/mypZ6rxOkTWL+FgDdi6JpmNO5H6mRV4o12UBkKQ6K
wNg7zIu+yiVFAkXuXiIqSZwXMvblwkDlaVbXOuAFPP5QQ0/TrNXYdtAOLlRxUvQEm7YEZMb9UnhV
NJ+PgM2DaoI8KHrw5TrlxtenG58PVYXkF5IzPHyz4Awp5k+9ON5VZdWojQR4f1rG4FfGZarPYzpL
mqQzNNoEbPNRNVTk6e+/eI6lG+NgiS45p603cSlCQrD1haCiNfKv60gvmUTrIGy8Qd2542C+o94y
qrGAnQig0r6Qa9K3fDBZFS2jmxNyjV66vTYNMyLSx7HWwrPZNiuMa+/E49vApmsINi3vdIzNOwII
vpo5Cu3aIl4PCY+xg8fXliVBqc6bzO2XA1r1NSnvpcPwqU+ZLa8gpOn9J4RDZMkLd27enbxmhwgp
zlKt2vXK+J9EBlwQpHyPPGTKBWREVbufh4d4GR3qzA5Oj7tZ1zR6lnk0tgTljPDckuaSmhrHKBPN
VwRY36GEFnN65ka3QRCOc/EPT2bZqdQwO3dEmXZAhPC/l6qJy5cWjtyupWhGfp9fwbMpibmoNY8M
eQO/R7x41NE1p9duHdyEUotwUINvjTvmY4B37fRbHT9ju25eFwHo8qn2vYi98onBGbBN4EMdZMVU
8FLXVd3ssFye2cnkfFA4Lk0IdCICcVPNyZng817kvxgIBG+PwtMwlPapQtfVgYkYJIW1oqNtMNgV
J2Lh7pkNXuU025pyieFTUKSGqPpQoL8Q0psJIS4zpFLpVJXbXB/yOPgpkocAsP+RmpcZHszfRIy8
JeCfw9LIlK2u3hyGZYkHhHaNa/pBYFBkJPXNDvckMDo5qD9GWvonzGfVqWoHGhis9BwKHDm5RBPh
5BBylvOoFxcANCSIg46YVUeVlL52KNMN79NhHA4bkQBMMkmCIi5Mtej0bUsatI1EQzrVHs2lOvES
D5gYu5XE/sKBx9OuZeFLG/uDUoTfL5kjcRPJoztNTbwBSTvXxZ/PnXHVXJ+BRf0Aiw/7Yo716DCD
XXVGWYySh8O6+kdsr/H7Hwtvv5LUxOr/ICynaVAi7rz5w+mYW4zdzc+qFggFeoaq0LweBr3rp0Mf
Gk6J66qj+4uRXUeQk7/9CPwEzyUuOnfsRVN8YhMLBpS/98pI1D3Ff+gclaFNJEWDb61cVRtL6WZp
Ctt1Sx7sv0YjSsTcQXkOlMlsMxVpMAKiH1Sre+v6tjaMws8QLPNm8Y9IgNk23vnBii4Hgisc4OC8
O7jnO2ZI2vXWKS0PbNwzdRzPNQq/Pghp2JrA+yFNJepk+Nqk2pGrTHC0LNP8ZSgb9nfo9bA2WQ11
AeU1LytCUK/aVKX0dCj/UcoEUQ6DoHXkgCkHUUQ6gumIUt5G5r2HJoonaVNbf5lWNgC15lgKamAA
pBKsuITzNVqIeEuBNDfjFeAYz3u3GHtBso9xb5kKyiRei5grZDOqbTtpoKCvKlyKEVyTQmFgyAIX
rNhFsT0A0kXrCLTw/52V9ZGs9Yyriuec+cbwuyF4t3MMQpVeQOkDlOq1BvYPfoEJk0bFeB1Rs/81
BPZywRy/MdSItrT+DGHWG/hlHB2PGiKLZ9xRWZ4VoXlm4FXJQMArrrbzzbyMOK7dVH95yDheiin5
8D+wRUdH6KcME1BS8+jhlE9rVh53pcwbRZXTweA7kBxiUM+jikiLdnZ+fm6VP1iMtI1aKGiu9dbR
6n68Gn9I5HlGEr0Ga+Rk6RXbZ2SeTFZ1ONcwt49Pm87coHo1iSX1bgJ6xQc2aWAmZNjoJxQK8YRH
hVhwkdcvqxe9sBsrUf25gguDyOfTD865YiVjNwbkCpzUFkWyNP33mrixAGGergokazCVt8FTZtAV
au/wWoAxkLaPTRv2zzY/FzhY6CdH00yg/ACb2plM0Vo5ZFPEVpjt/F2Dekx1Xxpb0M0WAihGiqpF
91bFcHAQbSy4YfPfHBNApV2v5DRriAKzQiXGZZvqFQMv3MeDDwEBiTuLFskXF6q1AJlnxMm0/hwr
YS4Ma32ClVGebYoWab3t3+8O/GVyKcUNew/U0NRo8JODrF8ekqoM72WbtQbKkICpIJpbOFQ2mWhk
d3vBj51sW+vavs0EextonSUmi6bQIMmp3K5sqW+nogfc6IXadKqFA8CKV2de03j95mR8G4YQoiRo
1X6Cn406vWqR4P1yLQn3aSVBbTPCaDHX1IBOCfMvJpnwRthxX7kDYTjjCMBJSD7e+FsCtP9tVpgt
FMkZmE8pWFEiLOjGfou1Akabpe4Wzd1yJOQdPLyy0mNvXP7OUt6AnqMfZX6QyXObZWUPauY2q+KW
WGLWshGXYsMeEhWM5llzUOIg9ChYx/zoXTrb28LJD9SY1myZ/5lwcrF0eVpZNO3NZmaKEfTZ1gLk
FNO4GKC3FPRR52TyIr3OvVMwgz2XL47Nbz1wIS4F150Z5kmARoRP7WBKlWDFJ1RFpME3W1Zjl33D
atIlzEU+Z51qBWKWW8UC4cWgJV5Df9zlM8izEVPFqc8vVTweucE+cDeiaFci6OXdU8ABq+xvji2x
4gwX6lIbXoCxM+N+hlsmjLadnV/luTtpCiFKHhBNVw/JCphNISwDMrfiX3x/YuzWB25B0FhH9VM7
mRq2iGfPE7mYIJ6NiSQDvq2XVT7laITMLSsH82x4CBgNtz6/uCkrbsGLlmZFXC4sEe0aEHNCBcLS
U4C3P0ZD7LGKZAWV3/p0t0I/oPBNv5iYrX6qF1ukOgqc0WpiJ1zKAW12FJh4vq4GZiFgCUbUMQ8Y
+VYuCFUx9mvlDAPn9drxa5jD8aYb7ZD6mx4cXfTXLhPEDrZLhpoqAonz5S0ZZdG2wdjY7wJ4wUlt
3OymSPmSVkXsokfXmX+8T99lhE9slGI/ahOS+DV7ABZ8a5wACXt9IMzGp5tV8ieaZ3pqzbTcUtke
GMrhyXwjaUA/2r1OdLUZdZ3/tMm1gDjO176UPdobhtLgFBliexhYG9I7J15PAL0e19LUXqW4lsLy
4Deuak4VBl6qAIXPuGSjGaT9L7JiRVl5gVAT0I3tB9Ln7ZjFoCjK8ev0h89iIRYJWq2wNAHv9Q/U
/OJZ4Qg3GYwj8zYfNdBWfLWoPDFkC5gzfDrDU95kytRWU0HLuKH9iUz5zde56sThYkLXMHClS3Ng
ngAyOSV62XRBCmJQt66hi2PrRlTO/7of4AHNOWSFYiXNXpq29HXbLCx1FwMmueRbAYYQhVoCac/u
Ov9o7lMPDMhemUiE56ao1yunPmKs1in/ORi1z4rq5eDA9zxXWCidsAHIwJLMZVsBrLKGZCTyzwZw
S/g3SNRfpow1XqYyFMxmYEoExm0K6t6iUYDQ9GG6hqqK9o73BdymrLiCRS0ju6K2CEia7TY1irEV
bQJ6ixLhzhju1BDOm1QYqAk1fYRVzuw+oHuV19nXRQLlGQLAcd50unMEKmaMt8z8yCJo6hEmPXTG
TLSi6pTw4KSScqdj8IumrZq1wsoIaqjIrlNQeZGI4kv6FL11R8syJHUqXqK/c09GMNrbSJUhDfnm
rQjWYYRDy5Qc/yCOntSbWFoHfzDE1F3oDa4ArsREHVQmFJxZZwNKgxurifoWeuv7G88lGUTjD2Cp
0h9UNZGjrryLMwKh2s9DI3qs6nk0msoEoBHCoQCPLA0ZIBUcNyb9t2lK9v9GW6uJU/YFcuIb53TL
e5n8jx4TTQnk+9IdDnb5Xgn4QSB+oh6moF1lU/echY8g3qFXusMNiGEhaOoOjvgtj1m1L9jHR8gi
ZITPZUswHgR3SInxfE80i8osIijDZpyl35OhWLlRHSsxACpPloc9Q/mnW1x+rhY+c552NcJ0sawg
mORDaDfjr/UZFpmj6St1yZPeJQp+fBCKC1nOVP5t72ifE1QI9Xkqx/FhC0tg/BWsVXebSEnSQUtw
Zq+vyWGwhKQEtWK7dyW75LRlCFuyAesqeI1xwQB8KyOj8iIDhnwSyXxiNFrC003mQAYFEZBQ49RO
CsYvsAvDV1ksMsHU0o70OaLdDAcz2mRAHYslYq5Gh4EoXIBIiXu/gQ2d9shYQcnpZ9bsF4OiuguH
P5QbPCO4Q8xaj1kOjMjUHrXlc+b6R4GmiRyKOaP0uFrAJ0GRZl6+n2HKV4kIvJavgE65m17JAGGE
k82rck/poGNx1yFHQr5rscSHDu1YzE2bwBZs8tym+a9Fax7zJ8T5eUqr8Jw3gwMjBByd5QNvsTEf
WjruHbD9o2Z1NTqmr0tmH1tWywxQqZgKVVRvUc/KQIiDB56aXY5vD/BRYHa6VpgkFMVSdD/+7jgx
NLazV+RBZ+GcQr6ax+y6Mq9evM+QvaS7DUJFBGmSJ260nH6gevfEXuiV/Tl+o7l+3D00KMMy+ZKD
ySIZs3TVri/odRblv0mra9X6kzCmw0ciIDrxTt5KoNH+PNPzyV8bmjMWWF1yqtDMhJNUNniEgXul
yb+o8Ng0NTQ9vuwM28nFaK+B/QhQuB2wv87powom5+qKO+EOaZfgF/VTYhTA62bvBbYkRASnOJl3
o6b6i4zQKQ26uckg3AFU+1caETHKPF+eXPoWPx7gC6SuRTOSmSmJfZUIWwcTUtGZ3Io0m85sRdBy
6RjKn64q/tIfCf9yJ1K+lG3cY++PbB4Fh0O/cdZC/pdEKeRhy2Vcpi3rqmK3NLRsTcXOBYhEDXSv
X4dJvmJ3xwNFmX9aoWelH9QDP8SStNrYKfiYyRHt657IaoZhsZSPdIkL6iMWz+4arhXro3ZjZByU
8L/SbRtMnczafHzrjPSidMNKt3L3Kz7I4n1QiFWwX78qJb9cG3gjbxWbYm4eSZkLupAYZgnLQ8ZC
WZjkYDrDRoHydrM3pOH0wS4kgOnuyQSGhotcElF6oJqZClWtkgRAh1zdPKY4E3EMdtOG5XQGG9j0
raAg0jIVQ+NdLElVvVyVu1e9W+1mWkW63QQqWgvkNcJHzIZMct6n8OTBl2Uf1np63ol1d2NVpOg6
DYfyAMHRqdvwGmWCr8ykMkHZV+QIvnN7oFwoCVu5KAqeLXwGHXOJNslehvIBd/UKBBgDVy0UoyEk
9P2DK5w9DoC4jsb++V3yR2PhSZ198kDj8sJ4cyuF+eRL3+IRfiFWzkhOeWabCZD3fetHC2HwyFkV
USPipc/2Wbjze6FSnXSTvE4xKEdEGzGV67L97UDus5T6hMH/3jPMjSuW9m7iovUs4RAMgb3PS00R
XZy/hfkUd2H+RNbzbCZcge/OGht/qbn9/fL6491wSa37+wLo+7UTwZQAWjhBewG9C+C79gjv5u8E
MzUodqbeMLLcddf6BjjoqYqNEOj0Rb97Yz2xBJ6aUNWiWVwjSNx7tVr98S4IdiuvyVhBQ8xmTHud
GM7S5N3eoXFlkFbruZjvdqMPpeISDK8oujtngvxAUpZXpbdDIQ2ZcAF0mfNjbqwZI0H+Bu9z7nR8
nWTuC+Qs4pL/2iS5SslIKlYlglDvINNwq4aNAeACdGjjqAvm+bhJG/wUw830C+wRkelammL5DWtO
k5xNvkMRgyW5wjhEmwelc3tRe/k6rzhSTUVwqSWE067pel3m8ciuv2vfuX8W2nE50GROGB+yR5vw
oyVOP0X26JZvUTlSW0Z5hkyYiXnyXvwfaklerCXrhd+t952E+be9zmh+ingKhp1+t7h2D9D6Ho00
x3DOs/TrwwkCHWfoPvCQ3p8FnZU9ZiDgfurRWk8zIOcj546ll6m1M6rlEkHBHWDVI2LVGe71gGQb
GuDPu9dFF3KH0jF9WqZE69e4yyT1JFkTobu2CEPB+wP3ivIV5bnoTozLkpJK468TwcFFvF12wSMS
OJ9wvlQ7MPSpfMY0yJ1MuDY8VHVMKg/xvIK5GaWo7dlI6QpUbEGwSYGrwFKrVfNCCgvRnKuXBEL/
Q0vvbF3YATCKYeLanlmX6mZp5Vvy3mGlJZPECs4BIfW1/fQLbf7kicPs2yq5qwngwPaUdCpFN4b/
GS2nJPy0mmLQeEpTUmshUzb00ZSok1r3QLTmo9FGUQH1pg1PBntvWnMH0EWXedxF+D836I43GplI
e7xHG2K9HFPD19oOkiazhIgkX5SD5tS6dN8nxOgMSM4OQ67XIalG6gyV3q5BLn7t5bJ80jw7UICC
egj42vNxeNzLXcR7PITjxRNeQrES/TE2DiXfl+jhPajuqV5jFgUz9ZQmr0Hrkt5bkeVC4sbMrJyz
UlvrIRsJN4FuVJxAYp8Jo2pUr6WACOqfAe6AUoz2l/LSCLpCQMJGwMAExx2Fsdt6rBhR4IRWN6Pa
gOvqCUnAB/PoZp617OUwMho1+cZdE3bDh8V1qnPzZDQbst968zTPHuw8vcqm2Kx8ILDej/b5HBGv
PdbhMzLAKHuUB7/WlvFVvlDUCcZfD9AwX7DuFS+zHgAq4Xu60TJMZpFiJKjgCnXqybpkmjDRZCPV
J8HvSoUgZa7c1v8ToOKV+FdVQvooRwLQcaRP44C0kRqJGTWH7lSWgi1m8lEoLYHpNtBPOqKHRmsi
hnh2Xq8KGeZVp3b2NVaVipKiwgi1AsMm3opy9yqvLQvNaCfCmXLPJnTF39avh51gWLDNq/JCSBEp
7KmE4J7wSHYUKvQVMuU3EJZho9POX5gEYCD5oQ84f/RV9VGDLpJlHWXrWa5GEsvnKO1ALne03jyt
k4FMe0CW76Nyn74eTPAF0Cr6WOfV7ZBM9z6Q+cvMERA1GmbBiRFVDLAXFa5Vb1JozrOHDlegaiUM
Nx45+2wWDNhuv/BhD1ebv5Fgy2SAHQqdCs652WTl6LdZdHhyPC3oU6uasKlKXbXYZxWkaFpTm+mf
1j1Dcg4bz8ipNLMBKV9jzQjJWZAs/yLFj52sZOFtSrGv3nEq2VDa4/++/GSooTeS3OPiOeaTQBtP
7nl8DTZ6g0My/EJ73L9Il5z2ts0MWxZmIJ1NxPNJ2PK9ARGB+xXw4nUYjUJ20qr+TEjzI7RozNqI
UGSPfXEUTFmoGuAabtAqG0dFKYWj7IfUtsgrMu7mHyhBKzM7AX4Y5z1zBCJcrx9Ag+6KWeK/WYre
dRR/dnSXxw/eHu4AaFSpheEO6phG+uU26C9KnRif7ub3ET4KQ1LeTgXPLSDWHI4CNi29gVEPPEoE
q+CLBYWQcBWJFBGAmD2Nvrmzgwab1l3PH1m2Uc01mFZQeGWwUq0Fs9XCVj8CE5gBDu/27trVYoKc
5hglIEXSmeew5Cjr+jjf+e1nMjANAlDugjtr9171QuaSU7/eaBEO0ioiEZ0fDDSMvTkTPDC17ugu
AWVdW6g/Igc00AWqYZ6bbbDc47+wX8nL9yYSl3s/phbny6oe1r8YoIFvHyTf+TSh2xId/5o+TZhx
AW6VF+YhBWo2bvnhxmfWkHewYKUCfWmW/Zmks6NS7NJnRAaMxrd/t+iTnUIMJlLGYAOje/Lt+2XR
e9AL0gJTnzpOjgiKZLOSBvP0ay+D7H27G7ZLwZ5a7Ashdi0kBrdtMJcEkp7P+HK8Cd9GpaHW6d/Q
RkwYc1w+WRVZ/tzuAB2Fh4xiyNVAXPHQdFTDwN850sP18Zxmxj2JiOIX/ynmZtIk4qOSd/bh8WSn
m1eYuZ0926y/FIBRGiftCXo8s/NJJMTcwWpGRouqJA1Pq/hnVotVAtHLkw5FVwQc58yK94yh2DKp
sO4WbdsdInuNv4ubTIxR2/fA2+rokN8s6FnQ2uPajo1/zPS+lohwPlRWh2w846KabpnQ+DGCO8Ot
CgxwNIIf+kOJObFkutyYTyrDyAL3gwDEJjic9lihA4ewb+6ERnIEHcMChGqO0DX63kubcd4Gh5Ry
2/aORRGbEzWe7WTLWjeSWOKcI3K58K8e7AZSi8qUZ1qRYuH3ksXCGlLvc6XkqBNvg6q0o8n7C1Dk
D4DY8J3TUkq1v+ys+AOh4IlN0kYiMCEovWujhxcA9I1PKBd+FUVFl2tQcfHPZ8IcVNBcojrTQZ6s
+rOJ++5o4birn0NzBKcOxd3n8LSpWlEPEMg/qPe30dGCprYR2N5dFi2LR6QBOvUCCqjXj+0y6gux
MnqNqPKscDY2A1K0m1imNUX625mQuieEq1Os1uR5gW9SxVy0vr8/y+JgpjJw/PNOiY38KCq306Zx
XvPRyWTisBKwvIDO5c/a5gqwvqktXu1ockBcPeMKwBFJBrEajdoB/3K3Tn1ApQzaPQU64Hrvz08K
tDZRkvh5QJREBFNOBVbXNhaXT+mObArqpP6xgW57fZ5GGGogg8HS15rw/IUvXCFqwH5MLvnvR9eN
kA6ZqpIhN0iH8awCkadk+m5UkO6qy5cseFHwQFuaSL5qHPN/aOXN4HdmSTxm9fmyygSic+tP47SR
DgRDO6ANF8w8SKGZrao7gbrVA9488LMG6XyspjDB+YS2VD7UEz6+MuuRnRowRtS0AvtVC4JxejYd
0zDNw5n/H8R6rrw5N91ru6tQWBTiYn6eaf4AYGMYnbqfE0WqcLecbtav2i+N6Edi2hzhtutIjM4f
JjFgoK1Ugg6aosH7rNJWbYUAKE6iwIbxLSRbV7dLnq0U2xmRIDFeRrOqGQEJLmRRzck3/PxzgGAt
0RUIsPhEteJXeU1nkumf5xBkthB2ED7RQTWxq44Bavn4BQ5PXjXUfrVVrXmdNp9xcsg2vHHqdF1V
zfb6dEZzGf9o3UvgmM5bAPNWSAufIiHEJ1s/N2casstJ8PE460TU19zRtWGOJAnaitiRNTrylhOV
Z96H/WpCkMMN8kTESr2n/syUz/eGWeGAUE+EOuLohwcSKnUbRJayJIGvoCWeuBxwKUR3lrAWXEOJ
mV/0TVR8r9Pg2bUCyEKgcJuHobKBVcbJnCRXoT7unG16XeFaZdFZe9KpITPzqas/P1b3s0Z7vvHB
xmvZJ3HQGiDvenuD0AOIwBUhCvlsVSq7ga4yAHHM1V37rnEOyP0y8KSmvuypDiUqdQFxBI07KC/b
MtUWwvB6W7j4zb6WhLsPm8XPEpCwzPVQKoTOeYLKbhIed4vGcS5q4M3FaQ9dlDAYeyABtKL8dUxV
cqwhrTGgj8vld4NXNpS5LydQdZPSNLBmZL61LpfeTulJ9H5CPOuhXqGf1EOxixLTPvdMEIdN/KOc
VPP6uVwTdrFb+gaoYHV/dV7G8LSLH3k/oDJ8cJCAAppcpKAbJH2w6jOQq3IZu8L3tsD3AU2+Fgig
mGcglocIhGi+IF73/ZL33v3YnDarKGKicrMfGcxzv2Qj01d//hRu9n+iJdhAuukntAa7/QSm32ou
wYBoOZS2WgD6gWVPxqwLX+/ig5mxEVSvGhy/lOcCMnbnQiqPmag8YIYQ58NfkiGOXNlNxS5DZeek
IqzXrDyhwGsTmjJv87GxBSQB/CbL7QVhjwlDV49pIqrZMO/5GUPhTqJD85oHa4Q0xU6VyXtZA6z1
Rct26LaOnUcPCu+wG/cpmGbBZq3FTR1UzAVAp0pSo2paHA7fKjDivyFVM9cuoSk8VVwExN97qq/t
ITh4+IMK3R0fjTgELQp+GWCZJ0VysuSD47eEvAQ/niP108LOby0yWftfvgHVMhhb/YN10FrlsVY8
bwVHCo00lCqQsGhF3/Qd5EWsUOVO5o/U8TBgZYPx+p0jflRZpOpk1zFTBhxiVUdNjyaqE8BCYDF2
eE6+nSw7NhlzXk+XDiWdIlYXPI2qGk34iDvIR5wcihGxCmjbCjcnmc19eB3xvZCbQrOcFFaKQYFp
GvvvDG/vJK47nPS7AYzwnZXgC7SeXAI+yT6ATK726nMWARmQIUgj6rENj4QII+n1yap6QELJ4BWf
MO/EvcjyGC6k6+i0aKPsZDq130UbMqy1AHetIUvQD2uNLyHO2E8senCZ4c36kaLZJsxO6LbvbG50
KdIq48YpNZsiNWfrZi1LxojpF0BrI2iKICp0BVSvAIXSadbyVwfqkX+FYyeLZTEVz3R0oOKo7tJN
ZZHQQrNAy3BZeRUKg7Tfb0S8ATIUPlMRnpFEvhHLKdnWftK6poVadmwvhe4uMyhcpeGgx3bYhChl
+p+pCeHTMc3tw9P0ts+/r9ll1ukLcLpTbYgajQbXLb6NJQT+2hy9Xf5GvXaUkdjohQYLA0haGLad
IAZ2WTm80gsnZD8Qf7/KJIIjkBU27xyRqAqeRWffoDxwX863z2zDjM/S4JRQUv2XJZIq++zxEaqr
gYQl4ieMJKdTmuyy4CdAtKK9sq8Qk1Si6950LUF0y3k6vDMHwZm8lWZtqS0LWrbxpJMXf4wMlwD8
DP6vSfLPBUA3PG5BBCPBWOLif8+NOxOcmJ4tPU/sY+jL6QmObZoEir9SBjOTFi0TZDalRuqe2Hna
co7glnc/AgTIxGYTVAV8FtbRdti4EvZr1xA6ZNJP/9+2juw6Aj5YCZY/aMqF8JxeY6RiSWqeMet9
WH7L0nHWsCxTBtl7SBfS8TVOp7Thm0R6tk6uq1oh/9YpRIhIBJWTQ+WBiJJiA1s9bJ07hKrFuD+m
yIjEmu7BkB1/lxrDCFG/92K/3GX6ylIdzsESCVcJUgsZ9igzk6PDcIDNBMvlBRSf7KI3nv/5FtVk
lU6MQ58hHYS7LgdLcUyF+utbIQPuKIxz4PcY4FRJF25TbPEC2QLbWivVYKXP0CevTrjeqjsXzKDJ
52WiDo34UUxXESYC0OxUfLO3zeObdBuYi4DQ/CjALOPHbIeuRD3mDYs2hAwpiXkq2pCCD9uLS+1T
g1TiyXPtYMAM8w+hMTlO9a0dLLDUO0P242OXpTCEnMPZ7NPBgmw0tVlIl17oNwCYKaoj00X8fgzI
3boA4k+8G5kKEnWq6ZX0MFK0Q0donRZ3o/l4vD3GzQHluNHPwAtmWadd5JbmCh1FmjrHH3vPqNXv
xEzYllVzPZ1Vwt9ri445jIs/qlh2kToH6WAcz6bzUM8O36+66xUCkCBFrSz1DdDh4VqSdh13fbaQ
jsgXIHUq3m9BYRJji5sJsD4zqkyeO2BUZXIkG7Q3J8XGKjrFSfCppLsvkLvxF3jeh7+NlyBRRut1
A6iYnKcF0bHjZWZmOiAcxj9gRLWHwgo6WH+aH6bp5pZ+fB+mfSTPmR8eUepBS85MXKj6kKxpnMLQ
YgQFxNByFaHnSo66932xL8GrvYXOKYFVz8t2M78jQx9awRRELRCDeEPevHvS6QNQ53kRWjKdu0pD
ujc7GPi9zdqjKxcYcS/sxS64a5o+EI7Et4YNsYh4fzVtBMTs653OjzzQ3R8JT+i875Vg6oBZP8bi
5ZYBrOu82YrY7jR53eYCY8xmGwJI7ucBtMsUHvZWg6TLjM/HiAI08VsZwvSWFdjJ7OLXKtaB51cf
EK/e1aGyp54rdfZOd+WQMjIEtfm+XdXuOl1ikemZv3Pw0oEOQ8xjwGSn5ps6NUwsWa5MYE+oX5LM
qgqp8X+q0w7bKOFuxIeKf4imETw88jcWtbuw6qClCObSJg0le7a/yGtTnXSnKhuKUKdC8dZ8ojz6
amH8865fz6GJxj1fAc7xzEhyuJ2fXZOkpOFqIf9y5TUeDCj7Grm4wU2Cg5RRkWUstZdlY/3Ry5GG
xyGNqFMbwnwtFyh7oiazF8za29z97VEq/pfR3OEaXqPDmEipwBnCUJtmiBTgj7eG7qPoejebOhup
FPkP3hfFDlse4HexucuJmtPpXwAeOPoHwiCLx6seyquG6QWXimZEd4CoL0SC8juzT6K8NBZypB3L
A3aoml2Sak2k25qcPAKxxImP97WSju41Qfyh65mhhAPDci9I4//mIDbJYX+RK8eBk095QLcQJZO9
NZLFVnwnUKgMl+xw/JiNiYF7294S0T+IeOAEjDLQ2IkQg6fD0muu0tYaHgwO6olGaqfGdlBbo9CK
xRgCAtCjBJzzv3m9ud9rxc3sadcRJJDHEr/NVeC5jqt1QrmfRzWpdcEEynLidUA+RvelTGlnnNJg
aVO/gHKwEoQvbAUs24L6VdsFAarkrwSNR4Xh9BSq69d/eOTaytF5Pdws0vNHdHLmh+USKiO5fiG6
K0CKoJo2ew+gOui+RGTaZyPH3dDkMQYxf89hXlkWncqIuYCmvuyuO8bztu03zkwbhLV8VTi/CwtK
YLp/MCMdR1M6VLJg2srsR3A+mx+pZuO55kY7cICwyyzAg2ZCh/wY0Yi5zwq40odsD/FWNL4LNSo6
Yo5BdZpQjZNTBb1o08JBPRdiiHFg1TCCy6sqs6+2l9bvBbNy9t0jaGAARGJOttZb12sWIovl0K12
X3hgZNQFtsqxb1iSlDbtU4KUWJAIVnW4xwDpKzfGN/yL1n6oHjE/O/r/CMjWnZGtiXlJTJBpc4+q
w0aMBShIEo63LP0KU1JTlMN6mf/RBlDPCcty+pEp5/juAR8HPzd5ng3MdlzbMEDHiZjIrNHollvS
wbqgkUhWMkHBgSOa05DXn07pk02HM89JhYekdv2EezF0EnnTHBsNHT3FGcVIjmXWtBa5Yj1HmkvA
ty7mROJOQ9DhgcwcxTCkOdImhYniZM49hKHheeYNt82rPAdyjrouM+C/6W6i5n3SBk2+sKqz7Jbx
SW3Z5QPkZb7nQGuhzCto8nbRIdMkY6vvE0u0s7FHkI09QSPBcwTzdzKI0lMSQkuxFagtEKB/K3CP
Zvj0L+c6w1jKuR/gQTjYLSdLpMHZeY/8dUoa4u+TGD3UuIDqIpGzqW2pTjRv6z+j0ER8MIVHyNrE
UdyX5hrjaZw6/2Sanb4dJptu3+XLkCSlIO56PAnhx3njyIj/tMTXSnqScbJbAw1NhRr79hYFr3Jo
KFiqnsC4Q1w51x3kEOUUivM+FADSjm7gYHKfK3GtdAIeC0zs+ln1EoTyOD4WBVtRWdT5KAhU4eU2
Cf6TmWHVO8/sWw02iprqKLInBEX/8jsGbjVe8bmCSEgsRJtd+cA3Z0HWmYXdwf0GM3YKWbe6nUQl
yWJIm0dGkyUW3kRGIb+C2ffBPH49dx8pa2cECJ+cf9+PDtnKmMvNK27JjZbKuscZwLZCRZBhPPa2
4uebb+lZeKhtAPRcbL/6Ym5L9dXz/1N3awqP1KuDZqNA3KN09+B5n1VBOUcjktP5rMMEnaC4uoLx
4lPbHNgHO8K8CqtjRXJPqcI+vpTVn+l7SL24w5d/Qa/hsXQ2ZzdRcKH4hcDoeBePO3dEfs4aNGOE
OtbOTsAK9db3Q44OFF53dCqe6QQJetO1IlTv0SL2qd9zAq08jPQaNtia7NfQFHqRQLBgYN2zDPxg
xIOU9dKoLn4SJXOmWjuAILvefEh8r7CjJEg2QiSpFD1sVp0aUWR/hUpurI4CYiBaNRB28km3/0X0
1X+7NvSoVyiukvxLJ02VtZH6oCHBUWjCj4dANrnIqaLHPs7BeMrtzQP5ElCBYl8iYEUoGkiPF/GV
ZbMptyTft44cLM2Xt+7Y3je1HOPX7GEmV4bZwJ0bUfAssSUjzwh2FFKKmBL7Y/hY5MN9LzbHgT+h
NmWRY2drqTHZ33gD1ScjsP0dwZ8jDwFe4Z6d84edc9Mo6LcxjTTk9jDm2JGmYP9hvxs1M47aKwsr
H44k37EONfaxrXMp8+3CKS5uASRF+31xCkPYeY8l4SilNq8Is6AUvRXn72HGzbOBUs1CZvK+H0Uq
LE6oRCWEWIpPudkyYQi96DE35urXRB3kIjJM+/c2NGXP5BIzNeyIH5ryZainFLQLKeJ+vr0jTXiy
q4rFqss6pN6LAp9zz2O2gd+iMbpwh2ErqxIgKpMv8TMtBAJ14bcNMhJuXhC0Ja0RITfEj8iQqdPu
dyKkvRflanfuG+uwNw+kkfwHDz3sy4seLdlblgpUgacm9HbGGvn3z35a5N7fzU46FZG1CMpQou8V
zB8hP+KmaPx2/AVwSgArjhAh3nI/YmUKcpmrt/PlxHBngUDBxUMw5IlkKAoQGVT2HEy3VnPGVVe3
Fx0nUD7OrRYIsa3vWxxHpjIIbAG9/u24AJejGoCzkqIZ0S1uPLg/hbGYkT+HsRfNkqyWXbcOFhPl
5qKw/n831Pq1g3cJmA4YMRZtwnUe0PPQLZ6aEzaWV9Q6QaesFuWL9ggt1PQrVAUtZEQWMCH9KU+K
HJaM1CQiTd0AfFcyJYj4q92z1e1zy7ju3Wxyp/I1FEDzkhiUX3PX3EOiAbyciAx1b7qCvMbae/20
iqWkICVmX8LYkXkEY3BjwKbRaU0qil5l9NoPvANYSYDOFqu5hcxZaJQnOHneTvtFYGCAW+eRQlr3
Exlu+iXUXha0x9nHfYNZ9FvYSiE62trqyQwiMKfeG2htwtIav79E+NMRC4/UmGwHEB/uZ0iIocGo
12UazQkumwAEeFb4XDRIdiNAtE4K6tqqQKWl4bhQhmkOPLXJ4YrPQu5ENctEQcPMVYgQDmlOJOVa
x/NBCTMVNB7D6pUQ6XufXSQiNnmmAZamjswJGByCp0QDcH1LsMGuHUr8a1rT3PHUP1tedZChJGWz
wWukU+0PIMASHl1gzpkgOfZn+78BenM/QDxtiMFh8RD0cOcFAtxB/1KcSnttF0VVNemaLRb6fRUp
t/GTUObfymcaCDPBXcbQrjO/t1pTUyg0gFN04kbxpbEqTQobFQCCxQwTebjMF1WF7Xy3dqYGoodx
dSt6UcLdxnXpP2Pqhsu9gt/RQhC31sTySa2ph75W3LAL3cnepMUeKiD2d/NO2dbQSwZM4+Yzaw49
Kzjjwa9Kra5P3lZsZQA6LujPALw5qBmTiaYsipxYZjp90QEbS7WoBtHQrM9QibDiB6Oh7II1CFc6
s1y+tfBKS7VLZ1sAFe6nm8ItZjENXOa0UhW60MNjJ50JnKteVFBi/xFzkHcxau5HuESR6M9h1npB
+vASCL6uoifNB500ROSqXpu2BWZ9oUUNhBTO0GgMSDUwR5p9YhbIn1WsWpUFdIHHlgOoSiIvgmkV
w+W0SME/BXWPRgJhoNz2FILM33SDWmrRd3pqFFtrovH5yH/Y7MpyVtzkEq1QqJAJBtaPL+3QRAKx
6voCbcq8hXsaKaRkOgudD6LOEE9xgGXcNqPebYy283EqXTWsE1S6p5rsek0y/LBu2YXyIO5TEfNG
ApwVQv31tb1YhjlZrcgF8MA40ne2LuG/wTD108hs7//M9XEWvgDwKqETODszEdLnbYEnfNTSHQOb
JvLDVsWMhanJKD4ux8y87kN6mSR3Lo3cPn21k4U1YAEvOxgo+zhs/zMyXWqb28ZOY722IyEeCxiC
rKxdh7pXC345XS9nV/9MuItlWcfOsJpMO6+pwbuNGRZj0Zbc17unIKn4tMYmX3SkroTZ+VLtuj48
La2whCHncaT9K8MJd1MQJyy+lELLmn8Us10t6YEYkqQ4b/3G1i67m5TWLjyC4tMyKR7W+z65AZcp
yjSwJMyR9azLYVnm7XrQ/mMe/LzlXKnxyx2mKy+fKCYi3KdrSW4RoaZYSCW0wLQK95COk2DtNssn
GPaO23F1c1mkuRFZegOoAdmEnRyEAdvSMhn+q+VdPdJxALt7XhM5V5MRXbGjXnSjDXODEUAqQbCh
TLyWe+ZRXJK9yjAGWs0dVw/8jLefFpDKSPwE8f1/zT2RzpBOTszNZ1HNFmDpUHc3LV/jMcwKUYpu
KN82eziXaqD2rSj87ZLf5562/rvw7yVwCucdPaKGExmAKx+YesPP+c+FXHbhg0ZDxrLL5IfWXCns
Dy7p/1Y26St8hwIMulEkabHJ63ErG2w2ZGMMWSKJnxB/rA83azwbWav35M9a0DoRl5boq6401/E4
Tn+xjW22hBUCyoJWbdzgCcMQ2buvkyQiqBZQvPWxEbzYSVLUIutGlNVU8UXRAj2snAuHghHVW9KM
qUW3LLR4iIlt6Ak6rNtowZecqGhw5AzkA5U8oFfjy/sExOXa1n8LLt62T4k7hxrxXvVwxN4CuY9o
RHFtIBlDS3bs2fF5XJQMHwl3ErpMBNUACH0V2d5GflwOodBU31IgL69apcNlJl+1Uo24yX6DAnev
aUN0KbD+CIH+Oat2u1VQIfccsVM0K3YbEAeDJ973qkRD83YuxS18JydbF1ze6JdzaXqjRMuoTTKV
IAIS5wWWA/CqBNPRgg79hhW3GAa7aKajhQGq/V2v8ptJCs5bisiaMICclos6PhOEIQpwZVqx3t00
bioDvqmrQVk+apI+fykc1OhACv322YRnq03uBXuMq0bq/eLHcb0WbFZXIqfH5R4+Wuzba2oaidvf
qsPQwR2HHbyANQbIB4yropd5D7CKdyuforherlz3usFOgZxs3KaJI6C71KpOhMYzMfwQxKT1Aw2G
WTvQI25jsgyh+AKeXqTPiM2sxqwTusjAi9Ijzo2Oc3rPDn2JeSHcvLjQbXICYutEYD2jnNgK7TYJ
7Nb/5QBqQtWm5Jd61cGxmZbF8ygPIl3h/1ykgnaApUtpreUg9/yZe0KI8wxv0bx2QcPQfTdKosDz
WnUVs4/j3s5NUtx5qiOr27n7mc5McRDss27k4NUW14w+pqn7pk0vD/HlomHDO+P94+9kzBgpq19+
8dwRMw8oosFwBWYB9+265YoJmBeFK3CAWzak0HyGHxxgM8wDZK3RjEy0CGtwOisadctt3kiKb8vw
PE5GLFxdJe4TzPSAgjuXXlasmV7NXiwxvc/YHYZPhta5DW5I76gT6TrnPrWwxglCUwB4aAYjcHJK
40vQU/y8bAOp2MuQmiprr+iiVv6wjwTQWSTUYNBrZZOHQiRVF1NFMZ8Otijan300cdTDkvenlse/
Xx9lbTDA70OsEPbeIDLNbk7YOv6wHjOIDjFXGk+CLaQwbimp4vXLLDFJjNykPbLuPsIRZBIPY2Xf
Q8LhPDk+Woo1SXwYR4yQf28IYqqVVTZAkJPxB/98V8WoWijC9fuKFZhs2/r3ss7iuTy4sC9Dk7hF
oug+dMSYBAJy4W+4hM88fcVffiCF3Q3GLlCpREKavMMPqVSUFJ8XY0TXb5/nn+qECs+23kbUod6j
o71Dwuc6bUMq4B9tAZQ17YSDzzXVjvxZzgQuenMbWoYsC7rEiJwz1lBR1MWsq6xhSP4Jxd5XU2KQ
xoLP4Z4Jx55W176di9ceGloRCrDVhvTnd6k5z0izlwjSHwcKVsSYT5heMV4VX7x5TRXJ8yVM4k8M
e9mI40UDcnqP0hqjmXNfRVdGB3VwK3OXJUtHbeznMkxp23pzkshIHVdQUntLs6OZPgRrU9R1OEnj
azIPLA1+qJOk/9tDC38vu1XDzH7yukjK7lTeg72abriAa98PK2uy8k7loRyR9wk2RIr12CbsudrO
ptueR97SfOndyvk46zwaWc9Mc1dq25P9UshxaaVaUrdEY7AdxsrxXFSzjkMrfdrb3qO8wPptCSdW
XYn65WRvsPVvKTr6jJFI5UXMEEpSmiDQ0hP2aeUHmYQbKZt6sANyK8GiRQmlFogwxpRwPR713pQi
MY1NULwVrfPv6YFmDphbBPaRe1ApUcR/1VmQra6Zo0Byx7jSRhP3sjhqwlxQgbSk9JyRw1781d7x
Qo+cLr8MsEzMtCSME0UTzZTqbP/oEUMzjjo4yuGN4Ab1RK1g+TT4LE+y6flwX3+xB+T+eVUMvJIy
ncseO7i5U3fHajK5hQgUw98vWvbQXDNfSgIUijECrwcVbujNQA+MTpk+JgG+XVFwL1HcURWYPFtX
cbAXhymt6Cv/7AoJAdVBGJgqOpu+5MXvBjMjvBa86EOt4DUGlfXehIhcKH/2s3EmiTf3vphVD1vH
21sb55tCj+vIIkGPOtqQ6Gx2BsuYr6mdJLmYHt77YUX4XcbHZpc1MzoFrv3Th9EqDeC8YFkYwXlX
xLW9G/OZcGj1ptikTO0zX+Sduy8ZJHcY9t7GHOro9H0SbrIqafYkZGQYNRsK+P+HzN2PRYbO7U02
z1FDAF9dqqj7Sn8LL4Leg9QaJpVIPQvB459IWuFS82mIyc/4yplDfCuFoeczgHl+qsMtBiNtjui+
YIRr9sB8/CIXDAtL9I/hsWbETwQF4OAP4Zbp+71gtT2R5nXim2NHbFgTOu+5RGSX0Q9d6rJjgrq2
gtJ4fxyc8O49cMR7b4gAXQUUPy0DjFpKUz/A//1Hd77TsOKMdvaXWtgGSBTu2BKaMaFVgmY7VgC1
s4jpy/jWUoIuzF84Og8p8Nq/Kd9YI/DEutl2XZgKyj8QAlO2SrtKISBMdNNaXHVe1E7TgwV9t1KC
Sb334XoxIu3pedO8k2MpYdPNRFqlPqXyw6iuzgWJC0JKNUQIFREecWcxTCQzyR1c2LXidozpqrOX
SBsveQ4x7fWv6/YteyYpawcKG78fbpAP3z6aM5NtQgUkykKG6nM61H5w2giv2epB6epS8AK8dRpf
OCGwJd6iVAPqdy6+h1HBJSkF4gztoA0qfkFEcsgSH9ImTcZmavXJZQvbB1/Xswp4K9UO6aPFuT/f
BMJIj1uhpqVfjJVWXLHuzsPAwccNplcpg29rv1dQg6mQ1injxJzOI69pJv5PmtH/9kpY+VZg6YbQ
iiefdNf6W1L9KVGZ41TkImzvxamrcUFOyqPoeM85ZxhwnR5Ffw5HNaY4UNNGIkBxYqEGrLsnnn3Y
xuGaaKSYbfPTbw9XsuPYg9/nn4EdO0dY1O66FUmpGJGa2BVT3gKoNlVOb2YmfK5djCJTe1oXOhfw
XulXuQfP7AiAp6+6RUAxa0uwfz5na2s717BIgyyYkmZXTE/VzQ+hZE80EJasVrcQx8RUBgzmP6sm
t3tfuKbQ0NiWPz580+IaEqNZ4bz/2mzgHDk2cNtiMp5BsneIqKoMrvq1X1GCYgwuG+ePZ7wQWswK
2H5jQPJ+ijlBN2yPxTsDFs4eZVvSc+bKvkbRu2Dc6cgsBCzff/2IQlYlnMesWN42pfXaVgykxFXw
Dcc2gRixJRz2PNtEut+p9YSwV1F7t23fHA5e918mNUw5zGbXbEwHf06ndRo/C2PlFH3vMqdda+kq
vsE9wQV/JItxTGWa7l4cFm+UBq9jY+zLdXPxB3qQUH5224WhfdVyQY1Wb6uGBWTO4F4UvBltamVZ
ep87nNEZc9dzhFyNm4y+ZKHWglsj+wS3FU24w/+KWfH+775SPGdLbYa1myFXF6oVccr6wWOF8lqM
z0/lVayda71z89Qd4kaPwshpHef2MBthD5KcbhzCIzZu/6HH5y5gfwZXPgISo173kx8PDTrtlNSe
/n5GQ0JWFovFQ7eQEPfxTgJwJPolit78PGyhLN+lXx0bSG6mVV3eZ+M3/4l+iFiKaxfpaIGkvcdO
1hfCXLKR2e/GaUS23yon60C00L9Fesgjjbn/7p6bjpbIHOUqo7A9awnsoyA3L5ayiWcPjlKxleNx
peLXThrTDqh7gkFbypQIhCq6S6QVTTtLlHtT24z9rtBF1jo6NlwZS++E92aPA1vhzP0EleZq3/kL
wouieWR4Io/Zd90e3Sc8SO+DHj3JyoLh2pLoBVfzmPxwfZ+XOsjZL1e3CygxEc8LRCJEWYA6kEBo
GtiG7xvOjhwQtCHLTniBdEHT8gCjV4Iqgrt+oMgCKD+Ph9eRUCNjnpeUjmSf2Z7D1T9xAUFWYUyH
K5C9rsZxr6I1YTvwRbEMUSC17bEU23t0iDnZ84l8LWoH1VMl3zs74d/GsindlRIRiSluuLLWvvb6
YAe5Bxt+jEHtJ1YETsyj1XbqzMiDXRh/uF3Vio4xSOaizww7J3d3+ANM6r/+96z1g7+d8gGVAnuR
d7ma+vTRo03EuGeLSMC42l9/nF2LGWpiA4MtTu5J+pp2Vl8fO9kwpHg8IsJIy3RCNSAha+8iFd3R
DqOhHoQoDnX1Sc+Uqccv4yaPh9IskUNkNHgDFAp2efcKjMX+DbIFpTw2b/vULLZ33Sf6Xq6l8Bqd
Ol+4Sr9RjpAJ4iHX0JioUBplixpYiyDMXtLzMOxJRMi902wDUCZooLZT4n+f6UWWoGAU6u6pfSZh
5giz/gCUtEqAaB34IIvGoQ5ZoQu8qz3FTf/BO7kEEgFkgVurCTq5FKTBqIlirL/LYUhrv9904/Bq
AGwllOQcS9b2yersdYR1yvyimDXSpbrVMlrUCCf/Jf+osCSnaRKsjiHvE355GDY27fhaXgHpNhnS
lDOGjb0vd53kbytvKKzz0HM/eHVGI9fy1qa/jKIXIU1/R0jNu/UYfa2Sk6ssyw+h8UCaS9aZyX/4
2Qh6+Dx7TF5Jf0DaL2WDPOD+r37wx1Uws4lRkX5YOdjvwTTPFL1IJwCUZDMAltxLIZfy5aQYjoa8
NLTDmbJ2mebHkqeAyBekGvH7QD4/ETEdFgkrTpeqjKC7bgfGfP0mZdtidkXIGzbZpaAEp/lScbL+
o7QgBNmYMavJnToD1DfC2OB5xJgT6bAigvDwypYYAHEvdN9EcNzk7GzZmOjqCgQsESovgGRjkgvG
3tMewi9aiz0DDiME4qLn4js4w0e7Q9ahZwA1bD8Ntqpxluv/GdyZtnW3UcjOlVdsqj/+N10PCJgq
CUJBVOKpUyaQtumahWG8PmcDAzjMPBACpA7pGjFA+C8BlnUuwTucL/GPqBYjEWM2Kf8MxytrmrRa
i+FcQpcfNgXMv7702Kk3M+YJoub7HYuuUA79+hic9Izzxh5xkpvcCut3MUfqCU3fDiKkjUVxhJWt
3AzzgfEpPGpqRAbNfULTW2lvRIN3cthecmZo9wK5nIvs81XrRzKaLDVUMhIJ/1iqm+pt8lzsRLUu
/tSZ4KjPAwW240TrjFLtZX6KzB6YM/VkfguDbnib4GcXwSOV3LddTLnsRvHFpwUcArrtqCl9v3mJ
qaJqdVNp02mcWhHUSHohVl0Fw80Md2NXxyFdqkjWjGd2AGS6+VwdTd++XR9EaZm5KUCnaaW+NLEW
iuHCfmtQCJ4f3nEtF/mAKWgW5uiJc4FwDde/mh2NEFUuP+lA8l801Pgp2iWF0EBFwOMF8rldlMIt
5xQfQ6RrduX7iNPgT5OeawiYIB19/EmykcMc8BIES66wZg1pftOShYoXqjKfU/rJJiKkqBRGfJ2A
v3Lt3HCmteqrU5ABKP6tMAy9gTzWXEWwB/TUMgkEJddKUKImYS4peIKJM4dKFzdn7ppINq7wrWuZ
tchWwsUi9sGfDGdn9LpE25TOVyMLMBiHnJvjaN/Q+9xmzSCnq/3vBC5YnBQym54BoUXav6lxjdQq
0fSnCwycwIFIOXIzI90ePXBq+MgHxlSbb0vvLPgf4sivKAYi3BPtVbLk51drsrV2S1Hd8zpWDsbf
SwGWzJHQJZabKeje3KdKr2a4njn5kD0HuZYE12BG7Qy98GgEd5ohU+vpCuDOyTK2Y9mg0ZUgEIeH
phWXWQTcvpGe12m4vhQkzwaPUAg2cLNGJ8NS9EmDZMn1iZa9g0Z+z5iBdvu6dl02scKQ/5LSmiey
Tb/glW4v+I2Ifx2krSzCDM8AA8anOlaZZ10iOoweOEXrPNknTrAvk7El137+fcXJaX8evon0rp9Z
2i4CdkJefMSAFqClNHtCIbxtZDPB+4Ow+iSLbIKDpuKjyj0+yLIcBcSKIixGuovqMlu7lSCBYWOt
2NGjzVdFejRFGF7YHZrhmbx3tSvu1N/pGHq8jwKjTywLglMFrQT2UBLgsK5amIZXWHsMhjMRgSs0
en3UoQ34a4LX3NrSfqAgOEOD32bGetx5sjfsZkzHj1voroD0z4jJ2zxj+bxYRUj9N1/k7AQjh8pK
xH5hAPJsZMc2WXC6CnQO+ToKXZdcGGQxVq1AYb1H0lfovz10peSFr8HPnsn5DGZnCGJGkswuxkCU
19rwoMgpIBOJjvDmUIPFv3HhhrG0Ubicnm6elonkgIRI82uDz8A/cQUzW8C47l71IhEI4p6cnMng
vMkU1kmBaHiPovyIfFXTN8LrwguiLZGfiRHJh/SuWEEDcC2bufER9wD14mMTsHqvn91q5Iidj5yN
gJuMAin1t0MA8jOCKBrJUfsSrraoNHBS5GFCb70myiSS0ocu0zqVDP/7p+kKOdIAoBAaTXBKhC9V
co6DCNi5IRzA5HT0o9574uvwwjQpk6MYVWWJr94vXYhx6BSJdbky+mFji9g4vsFO62xMQtD08/GE
MITLjoWthFgctb2OUex19mLP/ImEhw1ACbnO4Q3XHkV1NeWrPfJIAavtboMpV4zTiY1Ce9tJ2lOI
sUgbxcwhWKmaCj0jgQ24uJRkJm/Cmvf7CU8QzZrWaY7iAY9UZIm3yNAVaeh2Ax874VBETN2YlzYo
21YS0LdNy+xvI3rjGTvKK7JVphfvwItBg//Xj68/LcT4ZtO55qh9Ffl7rC+FPcg2KfaxhxaIL9AF
F64MBPfkSFxgkOiI9ybzrE8BroE7+pTB/GEWFgc8OVD82nxIvyaAlyrDDJkiWk/EutdHMJOVTjrr
F5LLokoF86+WRbSRM3vJUm/eepkwkj+kWQQGOQ32TaLCwmBtzNK0CaNmcjj3iWp1hsqYdAqrzXWB
ohGafH/M6KGeB8O3V6ER74DdJFO7wx6wkUW04Wupf8XtAlGQyPNM+Qb8i/I/ocbv4uDFFsgdC8UY
LDaE5xa6RkmB6U6sw5OwFDqFlke+/8M7FBAMYelMGnv74EcgxeJVBVj3jxO3XYO46/mPkLG+9i6r
Sl+ZPeoAZZlun0BO8FevtyLLQ64LhSITW63wWmrEopBjYVlWuG+Vxev/jX3kjoyA1LcaU4bm1NSR
5CXTO798GuFdkw5TQOyOsT7z+Xowb/q85grhuv78Kyiy/8o/MdhIJME+SmqAGNJd4W/rAr+lxOZ7
Ylqb1K6wJhxV+HKinNhJRr5B2RspB2/YUgIPj6jlZu39ugGiYiz3wTOuDEEZ7MLZhncaobaOKUpx
9RWjOrXjnMoGjTFceN4Su9JbiPMdRfW3zYFWH+MJBj+CVY7PfH60b6DoJG5yG1OPhw54Jf037auk
aVjTHh3k67JXLQJn2zt9yLIYym97pruLZMkGo0gkBOoTEfEKQQRcGCs3ykbog534Vn/Ir1UBvtkY
ZDtKQJbGqO63r8XIrPe52562YlkCeyxRsIw5Y74P8niuI8RQZXFL2kxhfmSIZw15dP6jqVESCD8G
ACe+VDGG7tVqPhR9OcZ6WdCayDausnxOMuuO7p1l7+pA2LmZvmRVzIshzHYp7POVY+t0jCvTDFG/
dJnB5AZHFR9YRvT1DWc9dx+1WVRdpf1/TIxRkO7EIAQOvIQU7FKczRXT75OCQ4n5hklndHyQaGeY
KqdI3/Tkn2OWv8WEbXcD1gTEDaViuxqVWxnVT2HrS+UlCEJKGR+bOTZ3kuJc/PbYHO9dSlWxNM0p
ahh/1EsWAI22eiutcdaxjGDvQ6t2v3E3IbVHngyuZCVlb8M5eC8joJztyL8frwQdVqfUSh2KuqTU
2TDjmc5Y+MStpyfak06Mue/ASZKfvWZ+KOFYhwb41b3WL2TpYAAZd0vf5tbQWmw8H4rMmjXbh9W9
Yv48UM2HPBdq50bVdPBvqYc1mhjRrPJZB4ldGm+qQsqvyrdEnI0vZQayqgBC6TnnOfW8gJGxtWyR
Qt20p6IVIX/1LJdKFNr9ZIfDBRaqWa09NsQV6LhU1waX0YV2/zlxXG6PjPp8jkav4CN6kOIuVDgW
+vEi5sgq127CnmMtF1cHKD/iGzMLPCE0s+kyGfi5apatih0AaPI8Y4vjobSqybwCgKpMw/n6X3n2
6mYN+JWaQsFyXQdAB2rt3eQetPT+mUvr8FurTIyzRybWNQG7VM7geGFozJJKyOH499ZcUyAzWqii
n+TCurqOfD6Yq848JC9p4QXtx8qQyllQwkJxZRY/IUOtJPuPFEWaFnspEAxmaq3WL14e/Mb9w6+K
2tSME7+/Rw3Ew7gCKAzFwtXQq2Geey6m2S4afzD3trR5kOuS1XcJ5wg6WaGeoJooScyUZfhBPxWq
eFu7qddazmfUBO7IXerJC+oD6zs8ZuMjubJTUsZ1Vskw7jJIkvOKW96m23aZJKz9NmqR5HjFLEvd
GxSN+dtpPHlfm5v2oy7Y+GF9/hRwi0CR0JfAWllfUByoTOTAF4Voo2j/KrCTUvZrBbo9HKK935/1
/2snMMLJZ86SPsyg7BqK47jz0jJ3BlgCAoReh/NM6dB5q3vbkr6D3rKrZGnhiJofUVvDkzv7CZSD
v0GwKe4nWQzLMn78uCYmRYnVKqj/NTMc2gRN5Iln3+fSfPsSwaLmzWy2fF8KEV0Vf+i2W8T+sbyW
VBX9tZm4SgimjTyciZKyJLN3waHUU/rqNMDIiJtzWjNk2mA0/JylncKSffCT0aSDaS4JuDZrlDYG
/6dZmx+UczrPnytHOa5UC7WsYCSvHJ8VcbKQkVJEaLHCE/9Pd2B5/JCTxQFFc7cUwnlVrPVog+AJ
h+SPjRbHVhbZkwPAfAS5HzOWWglK/I/herTFhC5a2w4UxzPtqT3IpRZ2qv8n0hRrqAr3GtgspUT0
QjJQepm4EajJCLqSbcJ3mZN1eV+IZexzS6ZejK4NANvqX32T9yXbDewWw0oGKSjcp9fyhzJZuuQA
AIc4IhvtntjmpZ+5a4L1PFtfUfbrQeOTt72mwlMVaYhOxm82azkIxzcCU37TwUDRjQMktt7BJyDZ
Qm/Xp8Xs8CuESxJNv7tezYdE2t9o9D/Wgm0NwOxkxpTrQjZEH8Xp0HRtoWKMLQXPe4IADrH1nvHx
D+Q1LVk6RR9v3aPjJz4//spIoVRKUyHiYxGjkwNAz/32+2l3ZSsGQwoEGD1vwYeN9sNEAIZRRCKt
Iz/J/FrT8tBSK/zV5eBBqatMcdSkpPFq8P2ZdCu7pG6CA7ZIg0k5LGbelZ+Lk5WP6PYkvGNyBlYC
QMVFl7OQ/CmDEWbgHUYHPzGnmQLV0rSaLoIIZH8rdiv81ige0AsEQH8Z7bmMAo2Eqc8U+bzYycaW
svbeqyDOroZw6GtAKHBpZJG/ddXQeD/iVe6uKdabXEBTjyv2ghnRz7PL4VuZcrRPbvNEhko9iKZd
ozP0g0uucUEmj2rs+GB9iE1E4yUYOVkVHUXl59aat7KH8CHRILSCqV4vH4vIELJO6Vioj1JSnEh6
xydH9HYYJnUtFZir5rOVsl8Jzwyhq9JIzkW0EC0H9UN73iS9TJRS9sFdUdB0k8EaB1VygTV7Yuh0
gSVpRDpm+IHIFhHv5cgh0gkrmBSMDs/TfhkMRPlvEwJN13yD3fQ56MsO4RTr7uAKK88BlDXa6ygK
R+wp8cNfT0f9i0l4ksTEnZg1vKoUiyKEwfYyhGQ4272/vGUDrsK9oTHdzx1YweFoUJHnX9Ax4tHP
qRVhldrProvtsymcSXlw+FT8+grXTcQfB0wkVElRbISUTvLSRrAtfaioYd4z7G/FI7EZq6oqg1Mk
eeYmzyP9RwYEcePaP0Bu1wayUQWF9tICbUaopmkgNUQScBza4+8DNkCGZJpH9l3KL0Hha/OBF6w4
VmUPDu7mzfzElC14WYqBxFs4RMtqBTiMefSAzTw5k7SCmjyovfNucJcMDRf4bEtvtZ5gBsbraCRk
T0XXwz5UxuX8Bv9r8r2twmS0RIazJ9sChmb2z3Ui7MPTc3bM4AsmADJvO3FXGucr1J8guB04tPrk
U37VhNk/qxr4IT6hIa2EeYfHiRe0W6JrdWD4RvOuwr7Y/yqe7J/LcMsS9gP2sjE+tXpEfGf1H+j9
8kzxrqMuu0A9pzThnoJpv3wf2yGC2wwxbo30fSS+8lJhiFETwiqXGAY/99SAhDITwdY4hGYasmrA
AFIpM9kK+HNirnFCFSJg500VxYsURD5SVkbS50j5GwKx32Gn8jNmX1O8onUv74hY3Q+Pz1njhfMj
yv3yCQHkUihZjdm5h8HfMGzO9zPnrh3f94XFH66ElWXUpPOXmfImAvdN9VY3ibzU0zwbHoSCkwgH
90MALHKYWBwFRTbAkBf+0m8fQSj0tvCOAoDbIwV2tvHmTHlv2M/1GgLAGUnE5r5tqv8cmdgvZZkF
x5eB3KhbEl5E5bJnLB96wjTwUqFNWewdNGtkIhKUyx2hG3OuiKL44Q91J4u4/i+HmJFQK++nTXYK
OLhM3OcW/rnf6tBLG3TM+crQFUknzyr6uXFB8RqePdnzNbnrLOglssgH0OhXmadqgTI+zONXxHTX
i3cZYUeMOs1NIt71M53fRPOw26iyoQf6Hb5rWwqyP1ZR01lYkTV0MhzClH8UuQqDwRkUKKXCfu91
69tsr5mLzm4AtgYqk/6qUQgtNcWSWfySMtac/fyvBB5QJOuU5MfV732sdUhkCdIRUBkH1XTcKnHc
0cu5e081Cb1VclOTkRFRsHG0SN+toulwayjk1+ACtGMCv2H62m4i2J8DgD/5ganxIYmL9BGnIA6p
qHXwJEX3ZaPX/E9wNnvZGcMrGzP3CSOYPy2D5XAA+kjU0zCU7gw5mAHuBlVGBkIbLuOQo+Xy/ZeK
QcPihFSomiPe7MyGcj51GQLYPqIJxjGwvbrI91oH+DkrNrg3Uo+LCg3T/G7wxrTHkDD4rbQNeiMk
t7Is2GyzIryoPTnDxdfLBsyUwOlEazI+VSog9rUpuzssF8vcSEia9i+jDEAAti9GVGsAsh/l33fe
BAicJPjUgaNsLpIOJK3FWodhuaoGifZqvBgYf7moxxwV4MgmOQjxcYKyaY58t117+yyjDzVO9/lU
4yQXsJhA7h5SU05Nz17CQcHpakE7Krd+qhye7IB/7vBUnCXHqFVngcIGSS+dbuZ58A78HDRfyGRi
hVtpAMkiBeYNbSe1cBMkz0ULDZzSzdFyO6+cI4wb1iks9vKkUkDVHj6ry0XuK5MdP0MdK5Gg15YC
NQYHoZr4siSNWzCj7rSiyMYH6Usz3keG7jrx1a9O4ivyGpLwQ6wNo25cixhwO/llLB6JQtHbWPT0
6Ckz5zl5LYR6vCfG8o1MtL7JnNINC7SGoz8GtlLnTTd14RpdToXMT5p4n+6nIIXL3AsxGDmQE2q3
a4635sNzkrpIgqE/Q9mGQzIbWoz0mnF124ZSzQiaCFWC8+bI5EMdRblWK4pGqbSJje6lvtxwUUiS
krCbfnjVExpf05sjysMxLyznrfi4N261Hyp/KhN2sgrDMopayn6oDPL68WbdLWskEiKFxlXqw7cr
KjWgt/XIIgxgsVNi/ylDtDk3c0Ec49OdQfPdRmDZULo7hnocT5gMqBpGXN6KaJV8EecfrtOU/9lt
0Uw2BCDMBsqfXC5taF7vC/yB91twNvQ9n9fyF5cuFWXG4FYylxMbCq6NjfWhTjb6MYK5k6UlQ8Mt
UdQLe1gOAhvyd7lyy9ehEZvr8mgdPSQW0cUARBAMxmsFbteUGPMsWjILRIJl0hXmSkWUy/HmwCHp
2Fa8+t0t+fos8EFjSwGoYDYOd+xfTzm2X6tc8qNFOxbIegGcsOXNR1UoEJk5i43itZEBh40Y4rNG
5lV3sflfFDaFRx0DDcnDXXeU6fXaJRb1rfQFhWqyIdC8s5DZUGlVBbfTCHeaxGspT599II8verXA
+w/Gbbpz0nqKV5Za8B1tRiIy5OaX09bre2MqZuvTasjwNbCHcSZDKN+j0227T6cWbvUuJW8tqNNR
JsbPl15b/WriIi1aSjxv4oZK5JbV7fKm4XRqUQ3pD06VcFCCb4nAO6rzQpPRu1zzK6CtLypJJQ7V
HoBPYVrkh/6mwnCvUtjH5Vx+nmRTkWYf2AuAYAM8BbQgDcF5mOAQZNhnMVphYI6glvK8+1j9wYyW
RgufexXTW8vYzyMnr6mDf21SZH5ytsHsdq35kaZNZvYjmvD24PksQGWEgA12AavBa81wu9gQmj5x
e8iiSVGAi6OMrBPWUf7VegdmMok583+2C5v1DvImN6er7m88ua0BPj0arHTVHMuD3x8kp2zHziN2
5JwmMrnWGxljMqkKJtkltpudWksrTH3MEVZdsnWb3REYuHstp9R5cN9LI/WXiXRBBRU9x4NAEMU5
7RY+PYpFyTDQ4DJIcZUIW5sqzJFBN9Ut/D2e8j+sXf9vAdRLYLt9KIflGjTtelo9VqIFfLgTaFfy
dA5Yp2F+5N529snpkaupGN1BjK4ra1O7QHEwoMXNPdWyTm0DPFmCHk4hWVZnJqk5AhsVapeisraY
hBg+7q6mZRn1Y+PRmHa1M8h+vSbfvOel5d7ofpnq8jvbAdJy7JJYGdkm2gHisCY6udcxRmsGvsXI
RASb/t08h2MMiQZWtOum1XPVfOPe5dmZCANHjvCRPEmcjOvjmHqR2jF88PA/2eIShprVXVWAboeC
uE4evMD6vb20FgwNrhL10w4JjE9MksoK+TRD4TBCWL4KSxRYCV7l+6RGO0UV2Gw5r7GurilMVfBB
Br/bGjXAuBkoWPysiBQn3MfNNh9C0aucrdI3Bg0Un8ZRieBSGVNtLw2X8Q4k1Vd552K2JE/hmWqp
g9PJmc0G8Cqd9CzPgvWut/Wp1i5qe8TyB5XFZCKMdIl4qzU0uDEWlSxe52+3r9sF8OdjANuMOh4+
GdHOZeN4qBR5NwOwKkZSDYNF1Awohjmj/Gn0AnjgVLNFRWUNhDn7wTwh+FzPaxyTq5tHpx6yLbOC
UKGMFAMT46CBQWk/xXQ2E3GyCwWfqr6z/dcoaZYboq+WVRPr5079EpY7+EZXcpakQGviBOyEM9Nh
JmxDoyMtk0dvkJYymklwuZH1T6pG8CPk3smWK+FUBmF34BPZN3IWJosf2bqMylYDZiizv81rVxOg
5554n7pvZe5U2YPjTSDn2uVawW3dgQJSRtwXpk77dMo7lxx6XCiI35Ziz8UVMTu4FvLiW5nfZFeB
pmhA27yFIfxfNaCpwetP1WK45NNbkaXd9syYejO1V/F8b7GekaB/gBCPShwmGrD2T4tahdSAFCLu
IL56ws68rWYmrlOn6lbQgpPD9jy+IBEowrFC0QbBq6/SEFiSo0WF6CmQNaBmFi5FnxdYs+wOoqdb
JER7P2xpPo7uMJR8VT9YXFZbaoMdRKi+whcDWGo9PdggsTliaKSRfYtjcrKi3kUmlKfyFEJBfOE4
CNlbaBzskuhIXh6sISZPSwN67JVj9e27sWlDsxQRDAwD0RoEtC8NEfyKxuyhlKcCw+F9DIYDjEM7
STsv1qJRvtEV1X71LhIv+7Al9D5t0Kiiy3XskT7Ppnc/Jjhq84tbf7PF5C+53wqi2UqrgFj1/eGf
qcQ2EYq0nD6GiqKWiRqHohwoCHCh3mb25uqlonskQ26dw8yKinOoN6zht+VTE6e9W4WHKV1fJQ9n
79lG4gKmFJeIoJn1g38c7QO7tvPzYk4TvY6ydV8WKKSVamJx9RUeo9t5Epz4ALpqkKqVMuy4UGfh
WCB0mwC1GEYtuSX40prJ8iahS81VatHNYdBz8aEppUINeLCuKEK5XsDBWbRQ8J1kPoW/xTJeAXaq
pfZPLUT8fzYV5pffLiyJf8gUeLFmCE0d1z1aCZ2rIlwMiaeQIzKcIu41hQTWzhM1LTi28mtH/EC4
bn2ynHHWHUIL5HXmMvg95YMJ3UGzvUFXRlBOuxaRgYCMp3+hZc7E8xGZEs7+ov7V0uhhazeElUPP
US9qP0jfNcdEPiT7vgfTkCUxlH1sYilBEwqNZvhI5Ao7S00KrNoCPog5243oXWIC7COIw7+WUkKq
jtes/vWAmbbjjVrHJ5gpA3mS+EkZMgcYSAbf40B5YO02jmGKCK//xi0N2jlzzLMoBJUcKOA9ZX4F
r4SOeUAzsk8F8CpQTRplfxOv36YDDmg373yY6uYGfX2UjsgvciyUvVar1hNzZa1beLWJJ3RMImuo
7f7V015WlnStH17AAjNDzyTFkV24kQdkwhinvd+ASbL5HORqVDA2DoU+xWdwSvSPpnjSwKkPu22b
TPzOuAsr7MGgavzTEww0v4m5Z/CAIdlT8nD7zrW+rE90alwminM4+XcVu4pJE5Q0gVCmbUgz2jq/
mkoI/LUsu+ndiRkuktmo9IA0oF0a5ZkAOadj+QVSJTjwtCafCuHtSMhiGFKtrAQJvyJ6/BWUszkM
iChXutOPvESqzbQx1ABrczQrGTMI2736yLHQuU4vTU2vco7WC1tBDi6XCUp7AhExWqFYdWwc9pHy
GNT6HsiPUBmvUTzaVsmoxQ7X9QOKNozG086YuMxRNT/kP9h3xK1h+UKZpQgOYWwxgyjR3zWgHZjh
BJ2PlbTCOuPnD/GzcDyAwpZ5zeox/FWSdRPQdl5YrSkkei8obIs27hWrzKoqD7KFpOo/QO0YWvCr
bT71MmpCQfrM/PMkXbogAJu3VLjmFdilGNNNzwJBCa64a8pvW1+ebpY1mwa0lHZxO64f8uwMaw7L
Ip3BWC7Bj0zhKW7ZkT0O/ByyDKZkHr5a0fh6kTcGtyh9bz0aF8EMGf4E0bdpEo+ibtsJaGc8ppaa
yfPu+fAdDLSTo3fWrKjxZIZ+DiZAlfRo/F3Q5NmdUruTNI5Y8TyO31eG0siSrdcrfwy2sy2ZXOcV
Ney7Jv26Eq9qebm1Cal+A+YN4m+BUmbCHELp4TNHf+KFP6MwBFA2asCjk1du0f6l+hE5ZyCxDP3l
aTDIdbO1x2/xK+OsyJ2jlRvyCn/xE4XVE9JylpJl7loJ/cUEGpK7tNUMNHTqa4JOGs5zTsqB8trZ
vO/9TNAwiB73ALw4sa78hoXcnKNA4nH19HqyLk85fv00v548fz40S16My6Bp/9gSbxe6/gSePneJ
+PGHfrDAhPQ2bBc4fp8gaobpy87nktly/9IUvONsYjMtuVmc9XsbtrXxzP5k77sqAwsEIUITcCLC
SvysWO6AwJ4XvBlpnQMdUJ7ictEqXbCSNqYHvrVqQlIw3x6YsHPRP2tGj74tQSWntmK6uoEGISwF
jjxNILPNg47chV3da8xxlHCEAbMOd1b+LzlCCU7r895pSIDk8hxkpXZ8rhT0IgVRORgXCuNiumXA
9mZMvWNij+FsicUFlPFswtVCaPc0cmvHgKfu0ZhoYpDM0aJ1PxYVIk0vxfnikMmNfVxY1Edn2jZP
umYIfau0e9lRJf6dUM87Xt4pKC/qKl1rTwVuGMfUHPNnTqXRRHjdUiUzncjGEdcwKRDdnBvfDSK4
ZfucJWusDx61J1V1Rtc/HnX3+gZAAOBM9S7TFOeCT5gw/AqLzxcRw7xKFTMMFKtl5SD3vX+YZ5Ms
DEbRWyGqjd5z1mGDmyk5YZXwi6eriQxSw5WkcUVZlxSi1x9SXtCPdhijfxxF3PbUpqpBEtsXnvE4
gEg7XeL2mrR+BnEYMKyMuo8Gd7pZM2rbFJU/52R8ObSZ0QyihhwgUC0KHaih4iF75XIvVEUlnB1U
6OdkE1XEQGThIiCPiY3+clGiIo88jGTsuGnvBwtnU+j+L1y2U7d1J7SdPfF+Xge1WaC53LNyr6o2
pwDep6yF6vAxhDi5tnjDTBS3900rAxLRY5GB5KVSb+JYv5YnLLwjUBzBHwFlSybVj6s+D5l6+qb6
hhnb/plY/Xzme7xs2wLKvy29X4f14JOpybzatJpFANuFBh6XF2q/598X77M2ONekxTUIyeZG0IMC
xhE1Npyfp5mlbdAYRMhfNbc4tLysmBYN/VY/ivzD1HqB5cNJJIoPtn+wn6lxdgvvu8stRcSK2c30
xrj/wTnuxXo4GsQc/IZ2Izh+1n1bYZ6YoDT4oOz6zcanNqJo7y2VVc5GbQYlU34ILzT3wxtl1+aZ
7f0k/1+G1O+eOrVE0DydzTUpeUYPNZcNitj+wzUU89+jeAVvQg04Yi4Y2yQyQVH4bz77QdlYCaxV
sf+ibEiCOsaJ62vp+t/h21l6OLG5JH4k2uP6CirqOrGAYUR0SlJoKi7dgFxF0fD8bK/aL6h5Lwze
t23iMrLrOeBxYkMpzFedZbBNIBLoi1lGFgQQiRKo3kaThNyHIoopyfhcfAguEfrE1diW1n5xkk7o
BwHy+jU9UBTDogWMFF7Rsof3/U7GN2TBWA3/yYb9OGDbEAt07v46MFNOGmtI5UrdLS5xvMjDWxYD
lGRH5f5gYK7cnLZf1PZ4oIqz5kRZHMvpsfNfJTg63d+CS7Yh9g/T2Jv7ccau5oQxjOS8wm4rnDAn
/bqmS1yJ++S9+GMC6arzYzNVYQnfXyIxFnN2CS3prpQNkhOA2YWs7uNaxppvPFRIdCWEnbGh26dp
0plvOPnXSBpG8HiBydXA8MGmMTmVyGnvUnWV+7BNfZQoN5Ck7Kdk25d2SvSGAS/zhRid63dJO1qt
99gXDaxpyD9Ts4G1MvRh4NKW6ZTUM8Y21lUwLMPZDPG61YMLzFuzfUG74YngStgZswDVb/SYHPBf
qeK8D2EuGP5sI1AusuMcUWjMlea1ZKXSgUDlfA1M9SxCpVP0AuCdQn0JNtGZRojhTKQeIgkZrSNQ
ZFJjo4CA2oBv93DQqadTqxaX06fI44Pe1SUKIYq8eTz6meiWMef+R4MSCSE+c/wV2ojat/2mg8Lf
JOXlltwGRuZRr9VrnyUDGFrH1uhLe0KQvmAjss6U3otx6aT45otLiy7Ey0xGUexEQIfa595/LmpU
IJ/UGj+pSC36NW+eNdrzsGG2QL5XdkHahMzMuoAofssNcTx9aP8uae9a0i9gbyKuZacCjIjaNjAO
0ahQPRs8IUWzFI59LlJhZcWlrNavfMC/9BoHtWzvpIUAetcbqrar/kfmtW/a2VqX4hXD3gEN68oK
Q+Gb0DoZMzfhj5Qz+E960bCBWq7ddMd8dl+MMF+Vl7QNBYllRoZE4BebG+AP7ZwX5s6j8gD8vvFk
UiCkcJa8dA1xy9yKYiviyv7YXeORWDhmf6Ebi0tK4bap+EPALOIWR/KSWabIBeGCaxj7UwDD46R9
aIFM2sEV63tmUnY6MOrm9TdBwgZonNWA18OQWQT+Kyp/YI/OggEFsBgLjdDogBQ1G4AOtre4pzQy
WRMjahur4Q3n4CmE3JO9PeEjK4cjnVUGx4mj1gXAulg7omQqzok3SwVOmNRWsS0SWq24p45KXYbo
7QdZGeH966MPiubj9s+a42b+M6lnDVsV055FLRUsA/5hvlYcZGKPcMQK0l5m2gImi0mMfBC9eObN
YAlYsz9AOfawx91PxM30U2KoIK5QHu1BKnHqmJDwib9+HWwDchmCeqhkkVsiIt9jhDkzdruU6XeQ
MUb6I+LJzNa7W9E3PX7sf4/xRWpoAS9hyeOLGkZi3fSHAV0Iyduiw8qE7KTNaSjmtEzVwXNosr0o
PFy2n+lbTfyPLa45ou13PlbdZ2Wo94SN1M6pVScsDdO63ahf8mPFCvMRrByJzTqN8wN3dK0v7aNU
65oJ3QsC0HnezkyI+ZwTpJLuB282occizEoDGkrxMLzA5DQCtwgOIGXo48SKcEsJFWdY7loV9tGZ
G7RrxS/ogY2G8mCpGchpTVLLGsRnDlQUPBdrO7MKPQbv6UWWCWYlrU3nb97VvknX5MPZ/3D9cq9V
UMdKgGMadzz9HID15FvePoVcwTthpbY1gnIQzk8cRo50xy+LCRzyPdmP9U3PhTG8QC+SC+I1gmbo
MGUIiDRKYpUSOEPJzLerfQefi0fxMxc+ZPQwACoKBDi8ttlysY8Pl5iz+nSnLnti+k7oMw/h83hW
yG5Uo0+9XwNPNA3xH2tVoB9M8BllO7bX7zl2CnTlNCQEKjkpfis+Rkq6P5l09q6AwEgAeBM0Yk6g
XXvFZpc/D5UW0IFfyS/5nAEPnEz7sSnA4JmrDdwgXMhAbnFz9h9kVOnFTRU+cBfSrrX10SEDYJUQ
bRmi6f9GxiGGKoT7+lEkhiJ8cbo3es1H3q83J3F109oKxDQz690YjdC3PRbf/lppl/OkgsM20fe4
yezxWDfpyDtQk9ilV3dbXqBHwMpQVCVXB+JXESnyDRcF974yjbfRCh2dtA5+MAXhtmhd64Slxvcj
r6eo8aRKfTH0BskoYxfMFbrDUolhG937kmh9ORpGyD+cXAaB6j1C43oy0If+pfzUiWzu3qHmaAPL
YzNIliXKIaP/y+5GeKMvHbUzPONy17OPyBI6JH0KTQXxGcq1JULoqm+9DcyzEUWIdozJiO2wgq2G
iffClo3rxAq64Xk+gsOTeUIxCDlyrHgel0RV2PTn6BoVJ4XLcLE9K7y5AIGB24MqlWuedbpKKbMG
5ix+MEkwklbInasRKZZwox1Jvh5JOOeqAVAjeL8Zo9KHYlNIP27ceFdtKpjVnZ6RUBhgYkmqJLjb
h26/W7zHmbvYzUMikDo7rEkbuO+XpqccAQaNqgmkkYY+uyf2Ev8uBfVUzmND5WBF68KnoUR/2gDm
CxXk/gXmCClrnq9XTRQQ1UfiH1KGQjWH2zpKZBJThGgKNeUjkj/xYeso7si0g2kCbnn7srpf+Zcn
mJ2qcwR5nCfn7KSjuxIL2Pcx1k5UMdzkLYIpGJukQWo9fd2SmPX0pMTYdxgkHqpy2p0DydHeZEF2
UWL81Of3ccjghpIjTZlvWlVrRni/12urM7ayYs2yxIzYb6ioGXch4uhVzyqhcQw3LYs9gwgs3Z4f
o6WpGAjgFDpmQuUqZJspSyb3IyjnvhoF4Fru8Xu8uu+BB2VJjRBaSpjrr9ic26FmhK3PQ3s+KKZ5
g5nftkryjPHZiNWtcFUZvqQ86U4UQskaoiX36Zni/gRGurP+BXOeVmTt31MOGNRv4Vxep8HkhHkT
SG6IFc4wZHkzre/G4Wl6GSfZWbU2n8Lsn16OJ3fu2qogBREsWlSnwThNfBABW/3PCTxr8U0zAnLC
OlFdQYznXKOzOLhkrgsqAqVTiloQ+7Ut+dcYhbwBscfjkpddcGvhvkPHOCQcNNBuOrMe0lu8tD8l
F8ueLHludCLzyGHyeZmLgCW6EO0T6ywUhDZRf6umLL9CTPHssh7ezJIJAFDfl9ZPZSml0JS6pWih
Tg6X4isB0xozOgXx76dE1IBfw2EVqcZBXUs2f8eNSPEfewWimfxJ2sZFXdRu1xVdaFufScDZo9uN
SVBTRF+UqqEzRIYyYcuVD6DAPkUt2zmFPQCD8qIUi3SFqt36a61WQricl2PCsyzPGD+eVQxa9H0m
NEBQt/27ZYbQBbyMKnvSyTF/tLnArP4DjxpNOimWcGCW5iF5ameUuunDXDI7ea1Hmj3cyRKq7DH9
q5MzKioOQabeTNxGW1+TSLUKknz8nvUfKZ48DuAxRMCeFeuRg2s6r+Umtv6fp6D+Wer2L2SfXAK2
gch0DbmJvtoU9P+6eS2ztfSNx0/hF6Hcc0jxpqtl4obkq33gDiQj8KpN7RB/3BS6ey0Z9XATsYtB
sxJMDqqdDCNbXgP0AlchpLqiJImvplHHv8jV3srWkNNNNDAqfWHuZfh0eNkbmocw7odr81TgITcK
8okr8uGQEDBlqy1tdh+ea0AOLBIfzToGOdm2gSB3zDqM8EPVsyKMoWvmQggeU34Dchvu5B0kqyHn
4msNCakKqvYcum3OOzwsLUHXc4bjV9KWFRPtlgORp9mG0SlQhTKp67LOdpYk5iW0GXA72lVCSAyJ
81w61qpIkXP18DJrwtb3jy71in+vra+PemGRIqQdgxLj5WsxiAiFuP1DdQUMabK77mEhS/CoTGkS
LHSPvFkS/bjGGOM/NXtKqpdDiixf8zGelJzNCNWcVIDE6bDI4mbrUGJ5iJiY+xeqmlb/HMTzT1cQ
fI05cmRqSWHp4iUcQKWezknUYYzUOmHKCrHH0/BPE1RBQEQqJ9RdhS3RV4O3+4zaUYNC53Gu2grM
6YhzeusVBouiQVe2xB15w4tOqZYUxcKn7X0m6ZOQTBsk5AcJCA04q2crRypQfHR0fm3IdsG/wHO3
wKHXEVY+PFloCvrUkoKDa8kX3lUyvH8DzGFDNrDfVHbG0B0L/YAk8zFUHIFis2no/d0SJI41xLI3
+7x68ZQwiC+WYaySZDUNuKv2bXtKEfm9AORZwY6ea4ohdNFvUBCO26NMTFn3wDP5hMy1yUg+JKaf
hqWGz8cUgunDBBO3/1EaonRBTQM3cmxlpMq7NYDDp0Ix+cAjTTk2ZEsk1qtDrtTd/jn6VxGtUAKs
sSaRCsCesz8rVg9bagEtLgQFIUxAWbk6DfgsT2azsjKX4AITqHWgf+9YqocVrMYYNoZxZiv0uyZG
sWmwONTstlFaapgI82+loVINaZ3Xk6FcRTEu8HrYEz45kN9N9VSdIuzTg4UngoVZ5tfKzgnGLsUz
gQ7rEPTTHsDNa6kQ6qbvQu1iOR7ygeGG1NuqQB4xcTevfX6+lQPz/ij1Z3md3YEtQckQAu0fZxPl
GdicPL8QRSgj8Md6sM3naqwFIApCa3BnJRd/hHK5IKIrLau+5WGiBsG7wr94gCcjJbm3wqOMTUBN
AYGAfAgzd9SWwhCs0a5SzBbkUGunqBP4koGOLrwSpmtLucmj+/WUHbn7OKFz99+X/ODzHCABfQd8
anttwTQ9WsmT6gZoNfLvfIzmLkB1U0OdAArMDuNIv0taFDjpfYbbPfbIkKkiSTQP+8WmfdIM1tzX
PpgdXL3bH/W+A9o+UxKssVVGz2iG7M4GGlcWhy8EstxpVcRCGvJc1/aTb9w3FuwgoFsM+EqCDvVu
9NTtCWvP7/XhFbzTdUcgUFm+OezAu64HDJtyXp2a0bwC/XW8jNTE7UXbEEjkGZ58Uf+TFqjbJ0cf
QdkRhLDWN37Fm2rQlvQn67htFp7uz/GBI8bgrD1Gdj8d/M2T3Za/UOvKwlEgodckH/qQJt4dRGZR
IvEdbjyFQuyXgoiB7lNgQnjJwcBwZqwRiSUeluneaF8r1RCxxzk0m5JFXzM9xLqjA35Ss0eNLKKC
cgjYDCA+NU67+U9W+yip/33u8t51OjTJk6Y7tURPf/WobpXtITiH66QnUTMvRnA+fuW+4OKKGM3k
l167/49FQi+KPVSUOfEXW2TiGR+c9lAiQ0Tc7DfrWFlXOVO1ji9RKSXP+NpEKAlsuWM3HVeYDYEA
rvyZ5fjXeH5GX6UYzJrM/+zPMyXH9Ht4I6tRf7Wo9RyEuwmTgKNEzmRQC0ObA1yD1J5rkUQG5GUN
t8syup540mYVy3Ge7o745FP3pRE53HV288JeW/KVYuQU14PUfUc2Y4NrdnuL7k7FPreJVXKIwuCn
ZxYUEQOAGFqqpBqcrV64ufCw1odcHLwQ8tKduKhdbUSwwO4Gs6TtWIqvJDSuMEvjDu1y1skkKb+8
ZLrbxDK7AEdgyZZeT28gBXaoqAY4fzrw5pN3g6pczlIwtugWV/NVRwmdVeACQywDDYdt5snLwZNd
s5VNok0Se07JxmZY4EgsyR8BADGWuiyBLMux2oLxoaWPhfRTJDI3236g1RzarlQXCCgOC22BCnZ+
ECrkI0zbZzFfiVUrJ1ADAC+DPnYwXIOp/QDZzyE96xJlZ6LE2pHyWJN7+UiW6HOXtWtH7tFiZ2nc
B8nmFmn9HWvufQsE7VF1AuOOHTXUSK3aInQrfskQHMbMTkSwMb8Wa+8ZHYKH0DL6JFz0wgWHNdxb
hnDjgut9yGlr2jc86Jpa6rE0BzKYR6AJ9NhwU6arY87opTPYqnz9YfmplPMgne7KLPYp8WUSQ9Mf
zN2RoeyB8R+JXsaRq6r7AVyTP70913bRZpMcr5TVpK1pjp6KfLJcsUijmTXgtk4r/oUEAyNo3ZsJ
XO/8EOwFHHaEP/hm/a9GhYA6Qg7e802jfy5MNZfLAZXdouGrWI//HtXZftihFy5Yzrodq4nse4Pn
bHrSVeO2L3sZ7J7b3RnminQwLGeMTf9kA51X/oMqy+iv39YFxdC7i0Upzi4cOJj6txY1QdpIM8+/
2qvjB8dtf4+md+p2HdB2ZO2zJJceSfodEzhbkBin9npnrKD+Ou3fGwpaUogqXIyzIu5xZh0Mn1js
O8zGORbtf0uzcMpaqejyc7qfHu+bRWaRL6wddPCAuAZcdq9LGiONGzaQS2fPOoXWaeO+MMOUa+9N
189DYdKhNixB/P0+bItBpd0yFZqshVon8YImB0S9La4r+fYmEsaetdBRKhoeNNt5/GqkzEYnxO8f
aACmo04fzgYyRnEh1p8vr8zjZulGNxwAGtJcnga2rrEcM4b5CjlAzw4k1lKxnYduRpoqKDUO0F14
MTnKClNS/TftcxtwYcsGQvOZMAQWcNPkZmneFL01NY/e2RdL/0qPjWM4YRtyc5GBekebDVQs3oIM
OHW4LZHXUzC1Xmp1EDn0Dr7eSnfkYAzVGsn5//dbypdxMGvL4D9BSbJ3UpkMlTye5mLNtppINF3L
MQow8R/JSuAL/RWzRRsMb17mTV8zXK7qIzYyv7jqLxyc3G9YniLOqDC7whc+MKrcOnVhYHvYl021
Kk1dwNPLC13csEc2BgOKpShXw5B2f9PmvhuURonPcwCoSXVdAx33hDJtTIB473N5GotG2HXCvLfy
74Ggd91HM1V9S9IpKABphVtc1gVNq5rncno1/G0IFDYpCFtyAoeNGwL8WJyX74Vomr7LfdQ4MU5C
QiRNlQhYYSNw4DRNOjGe2+3wJv07i8+g14njKljcT5/l2yZy5BR0CSbnLQF+xA81j5YU8htlls7J
psfJVCyFu0mopW9uAJhzXqfe6zlWVe8eck3pt0MzxdlFf5fxNFAy+4b2wzetq1L0QYRfjbR0KL71
LhIrAt9Xkeesl/Kt0TYNj699N6jvr1SXBy1fzwYQDaPdyZZbSf5H8no6FrIbyNBlt38RbUSZ5w9R
lEDkQh6zN2DxzATCYCydpVRxxwluMGmdu2Y2P7MGR8XPgYnG+jt8ARZGLxFfli0WehId3qddi/AM
msfY3Ni+K7GV8OW/LbLhEM1fx4phk6n3AE0nb4C/VeBj62iUYC1O4t6CvmxDvEsFPqeSukbkzuEu
lINyxPWlfbCKlXAjcmo5APBkKJVhhBMRlOsSAvEXgUlOj/b2Eah9alH9w587TIaLFzy9eTUUEmxl
dnPgdvXXnKodsXDdeTP2Xp9dttLjBFfUgyaMOqo26hES1R39khCw6llqiubGbDZ//Dvtanll0okC
k88l1r/vi2jHlXRFwowH9h2nl/a/3IcUwlodtVInEWTtWz5ywiZeGjfqLfMpZyEIrQQfWm7isuAZ
AnQTllQTFgLGe8Vvy78lgfKoEw0knNxMjKjIlS6hBigJdI1uxs0hWGkQ71khkpyaXfqKoH32tRVi
ZMzwAVtj+j78joQ4XeTmBBUjhx8GH4AcjBDBGDCPpWe3AoHO39vBFTe/IDd5LcTe1s9sPGqaO3sC
RHCPVka0E2qoEQM7U/4fxLn3RDS3OZQrxD3jQFMhpuU2/leFgKkF0bpGky7qjCDqPqhlWrtNjHup
x8L9BxBdxCAKlhvKzB1GX07IykwG5K9HAIsQ9MWT9vtyI3NnTr42yQqTMKCcH4qIFll0cfmLIG5X
NqU6Q9sZLT9AsFbUzk9eq3ktJw1wPOKUkPH14AHShqXhxFoqgNuQ4CW7fWljkKfuq2HaueYamqPe
oj+WEh92paAZ9GR0o5PJmCmFiJ0pZQ4p08hoSYQ3wG2ltI5FjEWvmAxXbl+uhuFWF3J26AEDQ2+y
+og3C76zJl+DMnWEgXrGlRmGiGLC08jcl9dcMz9SrgxdbCwYY7NcEs/X/SAojLN7xyV7g9yTGPNM
fNo/0d4vBGwPiFAlTc+MM6eQoDDl3Q8i+IkjzTn+41wVoHrDvDbrEZCiVLPVUDBL9ovI/PZ/MC2T
iLXHIfPoFkbhzqC163gQrF5UjiHTDCtZ8AKHT5cCPzfHdZ6dgN3AiKROdbA2YVjEo63btnvckaL7
wjQX/feusxTd6aSvJVG7z5s0koD09Tranz3fzoxWptGVg7HTMhuUndT9KCIjzcULT9AJdTsLncLA
cxzAzH4LAu7WDcvg/Ag3fdd9Gs/QMacvh7wahp1fRKl/D6O6rauzL+rrKo3COdsbGfYpBOwN2GN6
pETEqSmbIOQtHBQ/DOW+NqUAyo13R2z7ELlrhGudnsodEdXxSqV/3aPsnIubr6Krjum2sYxQ+0nX
2ayOAre+JF9ZcVyHAnytVDOW/DYGVg+yF/MuvuVSmCnKjLTsDQ1ZDocrSY3L8nLgRQ+q+Do4JdS9
TK2r2PE0XX9oSYaOCMmuuVOwKQTwtcOthyRqkkUqwxyABOl+7Dt3HxEOWZHK90VDy2cic2t2qJzw
nChdr8NrTkTsM987ID8m9xlN4Ameepsn29KEIpJK+az9Pwy6Dc79UKeg+jfQtuUQKHq+b+SoNF+U
eREGGDYa4o0Wr5vXRakAsrGiRLPFYn0Z8iP+SV3g0d5G6bBMbLzXaIYGMlOddSxIXZt4yJayr9U6
xJrxSTgiPN0sXq4NTe28rhfnpXDRWisqtMCZluTEj6Am8vhWNj8QnV67HE22BJ64iCKGdLajHvm5
cZWWo+lKaaSOudJU6y22nIV6JMztUWYlG2nYpSl0GdaIpZx1xvqONIZfNUeHzZi+x+tuAF55O5KH
IabjbWeJbLnTvzpqQJ246BpVXU/lmCOfyfUssv8gCyxt3Dyh2QMdxTLW/fcx7rJ28gXW+sTSBjnB
X3JIfMWfkzuVNcNi8+ZbAWENpQFkspyfLqlMMht6RiGew6HylgYpSgkT5A6yZfT4Y7k0nBR7NmB5
gAgewN68SbGet+7ndKL1xWvbNp34wzjeO8owemdYiFsQqikWJyDYp18PgyMbq/o4yKAqaGwETfWf
APCw8T4DP1vMjcQwIMCCs00kRfwDc+yeZTd7IitqbWZY1ccwWfs3WI0AowoUr13kEsNQqDyeC2H7
e0aoMTzzRa8AD8d3TlMvggiMpY8GXcJvggdBVHetX5wq/X+n51qc06UQkHLcPZqcsWxwQupWe4ak
2sKb5T0CK5MD8QWnEspqcjdkiyFbCUrLBY6wipDvrlUEMbJxBs47gMx1yqEeiccwGfN4EOTWbqF7
4NLHGf/Fgyw6icmLz9QlWYFGMQ2+Oc9ukblhAZL0bKXtSo2DP1BgE8Xxk8ocdfCSs+hAvuEfTrI2
QOwv99es+cnMH+gyRdESM8zeItlGaVonaq1SHciwGiHyQDODkGAQJO8hxujX8r6JKP6JRz5ivgk9
jsdPsmwig072ZEJcMmMddVLSYZdTDClP2HKmJj1QtoeQRQZrkDmp1ahkpWwRdsUShkjcGgOylssT
IofLybmGpkY+Shu/6jJGqY1iPhVmuQmmQux3S9BFztsIyZP58ZBmXf08zaDKv55vtCP6lnyDshlG
nrJkRtEm5E45Zq6shZbf8GmoT4O8xmqOwuWShsl/iOV+6tSc//23tjwKI9Chln+y8olzhseno39Q
HXdlD6CpIR3RnNHTVA5fl+Cwuo6zcu52MxuMspU4ZGjXuMILT5m2bMKhDBDx2jkUmTNAOp4tCEGP
41bJ6CJui/kKQauVNwnG+TiV+KC6KvPwkqFsnFIyCXBWOzplMwgKcwvsbv37iXzue9G9llp187kN
Y4FWoSKet2M153imtSu3UGKsdVr9U3VJhqcBvqiKclrm9zwaHzf7+FlAVHU1tXW2iMvmXpwIpbMz
cyx+xdQ/nTHcoyvLgCsXIXTm+ceEAN4Zfu/i3L1r8iKD/oBKCcCFJ1VB1x3Sg5vj7nARrpVIhhy3
jKRUIKSJLVnJxK/JA4CZultFKTqpY+7pmB7+VnXNcWtyrqjxKhpUMG7+fBVlQkpe6i1RC1AikW3F
vYDd6Yu4g3EkU0IRi46wZ09fXn+ciKUuODtlbGWaPIRrKRdhkqTs0Dwmcs7AJKCudv4SysoIGj0N
jSZfFkjrVW95iO+20SMflhuueHVf77QgSC9ebJ7i31+DVVF911Ow8pNp0zBvSwNLZygkj+P8Zsj9
quzhguaZMvimnO6LqLgMv3vxepjY1qTVKRSBIOBfVY5VrVo0OI320cXZnWBHpHe2JXwyE8YiqwEG
CxNV71oQ4RoSLLqdGg7/sAqulVn5SnyPJaDN74apSKoT7D+iGSQhqvQoigVRrdy2pPizKBVOTTpO
ca8/yhxWN4dOclMXRvEuenDE4gyoiVZRA77gAejgfqzyG/mIDXMchgvqHwEzC071MGppidq7ytJp
5TYMVE4i6KCbbJJ/h6+ywTDqlIxTIopLeEc7cUOyP6+0zqlM3iRS5UDT7eaQMPLZMi8VEosS8Pq/
d4RuEvQ9+Wxzo9h/mWldHQUnmiqu0p8alPKJuJuNQYrxtIZx0qcNOtXF4SEPirc27NzcQcJ8680H
dTQJlD+wfC+aMd5EaK/7p4bMb8K6fFV1e7HP8W4KkDTBtBHgj+WYz0e1W/EeP04oGayRRAFTuuLA
QdtE4V7xdWFhQaqIc/t6+9A9PZAmdTYk/LyfogCMEv89NpErEbZ68s2f4DaOoRtK4NocIcUXZZJ1
iPvAzgYSqOvUchFc9r9UOjmpTRdFeGWi160P7YbyJq5hgPkNi5rau2jZQmpY7U3gwDvuf9pTlPlX
sX7qv42L/FwvIiGWZkiPrvTQgy0lklcaXIh2G/kbV2S1ibUKsc19YB0nTJQ6/emBLqUc3ybkh/m5
/dv9IaZ6NoPI5TE1c7sOVpcfNwsQWN+fSG2HEoW0kgcLLGDvbJwG5n3INyMcOGrgpOKWjH5PfNLh
5orCFuteFVYS8XDMVIRpX3dFyFuLUy75zRvv4AeHA9npXYvVZ9h36FCI4qQ91VHmmog7nRq0Y9da
YMI8NmI+ZzM2AlGOZW47REtyLqn4fJRJ1aPD+Qmd/uWr3Oaj/2VxoRMwx6pSrh8PS1hHdzgAVTe5
muKM1WsYAQKJ/h4HqCXC3ZNMGXkIacHvPUri/1+VPuhsbLiHSmiMmxVmG7uiUDPT4/PHk57bBjLQ
b2XMeqnc2VGICby/r8M4mUyf8wSgzwY/HPptYMkAWyEbTrk/JVzzfrKTtDFzRpsQmZh5K/Q1xAZc
OxUWrSNVrZY4R15YHskAVhh5hgamvQ88717HxPjaqMDeTQa/770mIbK8rodk41GqdO72Z8XQ99Kn
sxSTycioFCqpkLz0FIZlzv/z4Q1oN73s7gRnUvSaePT1SCaIDk0kmjmPDDhy7u7AgflTJUE+anUQ
EBPR4s4HBJWY7jKFQtnISZ1T8Mwt9xC/wFNSICB96wlUK11fsTvNHv4H7/Bf34aEs6hKMpezMesV
pbDAI9JX21ShCiCOn0LzQjt2Rm3yh1VoCQHopdpPL67hoaFnLt17+ja2v66CAujnboSwqeB/FnTe
MX11ySrYVibOGZKxZmBJUqd7ug5FlMXAO4E852DiQtTRKyurb93pnHSWVrFQdWtPtYm9+Wfio/+Z
dPG36n5ErX9OdA3Xjp3C/QfZIkYwJ3SPwWZpyMr08jMPOTZmSqklrtzh6FJpQXsrNxqlu2tKa0rs
3t7Xg+9KB8FltNoU1MmQnu/UcxrZXwqDCGrNXLE8QdFe9KLdKdZ6uDwT2tu0JBrhYM77+3sN7sbZ
yGcO9lnDrI5/pEPOXMvWlsfhHrDubHZP2kCftPwrh9CxDQFgdC4sr3H+LfPLKhLcruf2MEY33jW5
G1QxPRCFzzccvsb2w4bLChibMumfX5M9uL+X5jd/VIrdH8kNkzecrPJ3tmJBRKWLQq7CUbRhGW9/
sysDGSZ9KyQMzJVkFCaGKTMN0LYsu0wSOVgdRj+eulUFiv47ZD1MBY5G47fqHrLsLWd5+y2H8Kht
EQDRHk4qFkiML8N9Cm7Drji5P01lxBPwiNL44wbHQ7exWW9s5SiOoo/pVXohnYxJuIb/My7UlQaq
DrP6zbCYyy97320pjs2SZeJsumsCUR2SmQW7JAvmjCJIiD00fDX/wzX+EdCjukrFsQj+u3oqax8R
DgArCxbKtsruf0LZfRUwg2QjKBddRTaIstxW6948BEVyn8Xx0lYJhmFhQwNKteFnsu7M/ld3CPw4
gVAnVPikbfCxZyZ8k10X1k9BXpXBjTPvm0PiuvaI1GmdyqDpv5fSETdHL3xAMwpvRfTUX3DB5Z90
34wAJMfx80zL5DjYKJHm88tYE1ekPwWGUkCPbKaTmk4RcroXydlNjRJx3sPtlAWJ/Vwtk1CqSSvQ
FsO4LirLi7D6jUNeYCUajhAuM5iT9bUWCHEIkQ8KEvloRg7X/oJer/4p3ij7klYnIRbUW1jV0R8i
D4MmqpcNy6eaMz46DgJBRA7Mtm655hYcG6iDme7ACFC0nc9FGoIC3JJO4Tb3OCdFfHhthbmUbBZX
gmD7gS44APzLfI5eyMgKTaIJiKgmncZgxPfL1liPIvwlTJ/6/W0mMhMO1xaAQjtTeK1ZDhu0MWiF
tRpmd72NSYcNZp34nLAknzW5Spe+Hx1+glUDR8twELBzYAxNHH3YjGAHptUCze0SaWV/ijjkqm8m
5M4z0OAL5XJBNImAmy87svdEsbRQ6RSDBVEIa6WQZY7viDK68J8Ssp+Y09iNv9PhXMAyWU2XFvSR
bdu8NJ9yFGqwAJ1fJeHEOmU62JaOoiZ2bEFFUBfoXHTDWrSDhSJbiF1/rKh/0M1UA2HwXsSsl9Zr
+rK9Z0TXGMbbI4D4kWQNRnwkGaICWJARgAs79/oIvH/ZST/zSCEE07AMa2vqbEYzpHLZG62r39Ua
Q9ryE9ggQmE2u4erYS5RyW7zRvvM/u2gXYpAEuE3MFah5Bz5LZC/ObET/rosshA++NZBEr/oh+TC
1NflMedIh4QaOjR15Cbm+9NcOohcO/nOsgT88fK9IB1xCaaDaIdIn7a0wU9DeqbAozNlLyWbB5Od
couTIbKwXKj4cvcpL80znpt69uv4KrPD2+I0INF942RpXsJEL3TJIZoOG9AHTvC1AXEuzBkcEBsd
03EjBtyzw+I8Zb2IHG5UVn0BZ0WLFuGBHlOLphGrB+YHKpByw9YbjPTdVCsA+U+2ULAV9exgaeEX
vckx9OXj8vhNEicaUcNtrxZ/uTFAdAQMS5U+PJOqhb3Ec0bIQvVCHRwFppzYA0h44uHl/NbTkjZB
UHHUkbF56DW6wZP+vLJPE9JCm7nakbXT09VXvVxCDf0tgUcGEFEWPEmWJYk6fMw8w1JkADw7kPQg
NPyHlAfi/yj2unflAckmFoTD/XSmNeL9YK4gncRXjlhukxYnQcuTLOO4eT5gSwrjiuPicexG73gm
7pNDjpyoE6HDUtd5BuxNZzIU0KzkrLbIGX2lSK1+s+UOXwjz68IUGFih1Zk983xNlL9dJ79IopiX
DHd7V/eEIiVt7OuyMsVmsEArd4Jb4AkCZwFre8uyauLFxm/FmCSzEvOUlJtwkp09LkvWG1KeiCKc
xgvf4dWZDr7wuTmU3DWuOkp/Nn/Oz3/jwvJiR1rKvlxh5BEmUOHAJK2Xss68pP1/CmSUmE+ifo/N
aJfg02hjK2hPdcwRtoeqUAHiGPWGIRuTNWbXQe1cJ4JjE0D7kkuPPt/jj0upS1CMNkVMiUD8ysK7
/gyztEGOiKTqkSYgyAqNt7+3+j5sSp4bWyd2agj4mVg2ypzlMGEWfIcqh8iFKvtK8o7EBwzO56X7
Ck4I7n8gpCNfkueJ2HVoELcdtkroZfYi72zH5TXBTwRE/UThm6sL5AZ8ayoVRRafdEsGKFu8u6ly
dkvY9lu1sKxeX6qNJOIZ1xeZG+LBeAz7lFPtX043HToKYtMOppfhLC1rFAWdt0x56MeLn/qa6Yio
wL27XGMIWdgB+r3jprkaDtFkbgRA3aEVbaGlyuUP3zqgX92C6mK/as5MaECTSJsi49zyErZeKz+x
a75hqdXo25A+Tx5faxWgxQF10sLjnNJ08iay7yoGcuetc2uTSVNyHOrMErWk0hu5td/+LxaApYoW
of0WdoHPVqVCZ5dmwrUjMW/QG8KMlJriwsEnpsaQyXTAiFHvyzGmjppUpry8F7sbmTLXKQgIhjdx
c5WoQRGuuehk90cOJqikswTwmq9kUxPtx6ZCko2bkUIdyHTXnP2MnV5eA9dHnxweT5NV9EmXbFQQ
vl1IQs9JDWx4L2IoO6QVXtNlbcbyeqisy09fM3R63yhtOqb3YAddhj/pUx35z9PgSwbKnQ8Tt2Di
CExMBNze+YnWOUnwMhVUa/rfd0J0ptMnXm2yZIVf9XxS9bEUDbPJdHvJFcDeF+jNsysHKEhYlAhm
T6Z5nlLxvdxa55ldIbFvCjqjfnDslGtIDMclMBEQjeLAHzEckAngrGorEoTyswubBZOFStVgyQQ8
PPyuhYU7z/GMdXHIvoc326qUmYcDFTDo3m/JXIjNNTHbWCPz0SM140iHtWEZ1ut9P3rmCXkbgUCg
PZLDF3Pba35/I2qSH14gBMm9u9h5vgNQPHd5V0RBBuXcrJRe9b3hDJWmWk0ZXQviq1EWHLDCwwc6
Rcx5OK0MZevce6V67mkz1FoUSKhSrqoXJ+BJb5XWPNfoXyNnzsPhJ0XxjN2Uo2bG/09utAwIIERq
l1B4saH+capZoppns6hoGf0UK5w5HBSiW0xtW3xXe52TFahw09z8zzNiKAhzIAK6PiPMhyU8QsJi
mRz+KMLIgz2VTzhwuHpLN20daqAI9PuRncJmVlDQqW4Wh//mNR/ATEa8fuOCsIUrR3KxmXBcjrTo
/sPYDl0iPc6xf0CkC0FQywjf9/q3hoe64o7EeM5eC0xuLC3zk/5PLX2L7Olxf5XIwrYcr89733B7
iPp2+5+7z+/kDtLjdmFCur5doIHe+mxYDZ1wLVJ743SCvsz+35UTgwF/FHwNjp64Op/tWHIvWymn
dhdxa4uNlzGvF5Wri4nILWJjoLrL4mILA4JpfXiH37jS3judaU7VdT/4k1TefzTGh0WF90tcrIHT
vSHjPVj7/URQwQMSOqzqZMPO6MXNF688r0vg+BC+OLWzBel6Tm+hQKpTY/tOp7FMCe+HctkBnbj3
l/3NNX6sKLoj9/kCaGPC/tO3UdCQNuTvEEniQAWfHbwjGq0AUCjwzRGbb31xbSJwZGcgnD1XEBF4
dutt+SFRPAYBWD7dSh3VEwkx8byKenHe6K3eSgYMzd5/fdMvk//XOMr/L96Iwwq2uKJypdguVA7L
7keMRraJyC6sij9DupmFrEsg/hn0A3MTC21k1Z7MuBokOB9ujDgGkABUYGqGNAXgQ3G/GIELtDoA
1xRwNnOMD2HEqGNX1zMAg29giMlZU4qvGefZEgUa1Fk0291IqxpDd8+62njCMTwTQgI8Z0PJrV9j
dKiFi6eIHjOb36/E+jZiGlhrs6/c2iKOCU91H0ZbDxSf/gXjxo4ZFG5s+evUF06SzLqN5xMd+LAf
NIjAKaiKBTUg+3UAFMXjQ/dVmRIF/cSUPvLi39AfiW0qUs3WVWOfb1etW43Ww5Hx+waKxBB1v5Ht
yeezLs4ISyl0hFjZhXsd/AJpQuOhpB/LkVr2ThkoeUM17eLUYdQPpmL7KWXNvtVn+N8wtX1xn+H8
3NQv4QroDSIY9fKpT4I/H1B9jfSsM/RB10ig+HzDRbXK6kPW60CqWMnb6atsF608AKbIpg+3yoTi
j41LFWiAMQ3tk9hwIm8DmkQgd0Wj3xK8rwqRVUr5n00g7nErQaEgrP6iln26YDxMrow8lIRpCM7+
LI9x5bDySuw0oW+R/DQyAfG23y5Z3YdHAp06oOIDmQ/AC418iR+F9dM48tZkZcYchK9Sq5exq/dv
HyyccO7dkzDhfWipMlc9EqwKTYvr3MNDuyjHoMvbUSrt0wF0IIaUE8hlUyP+POna55dtCFGHjOSz
yGuy8Nk1caZkZNCxFg5ympfOJZWiwk+n7h472V7vEWYVfsey2EqyI3kHBUMOPVPGLa1KFJqZTYXD
xg+o/ptplhKdObQdMVPU9oxuW7CKVSvQk2Zwj69JjbbUKHvnKkQwNdLnPP782jTyYGhUDBzkZ4Bv
O4uZqKNK4Cb/qsQMkxT2s2pIPxfIUzjrTeSHg/M9AyzMq+2Oood4Ez0k7/MSppaQD3qoYndAlg1p
1/l6wYZUHXd8XqFkc1o7mRNQrGHUi66eF3menKr3hQ2jd4l4naesCcZtMR91K9uwfT7J9knvckn1
wGfYbugb5vye/siriYljYeXDwY+c7sLdZevFWzgBMdWEewNLzu7AjxfH4IvYGwt1FZtXLpm1lknn
sZzy2BRgiNmzYeWQvmLUhHt53HE5xNzmU6qr4LGb7KZtLTSsDVWZ4OZUMRa2LBFv7H3MsBLSgBOd
p4ZhS1+JgNRS4pU2ozflizI7QiCNpLcQ4zX65N8DYy+TALo4WA8+GU99R2V2V2WXHn7kYe787Jdy
tlt70zy2ca/1ER9RnvYS7iOofgR9wG/yZNAv0BbTJ0kwd+4PIDOYhNxvJateLzlVK2i5rmP5YvRH
UBQrlMqnRi5BqjeZY+6nFPw7sKoGAwHnaothjoFpWIve+ey7Mui1j8+qf3A4F8LTkb9/RsHtLECD
oJAfwuuUKMceYzvMYWufOFEMwTntDWangoG1Zxj5Fs90N9BkxKKWB+RsWsK693UedxXn7udCIDyO
PqIr5PEVzRESukfJdhWw07kyoEm3zDa0143dPxRxhio5hPvMm9Hvzw2c35Dmebm4PxO37S2mIEKX
4brOxNY/1RyfY6eGIt+69vwE3soF9yRN7tvkO9dBWp0eN+OuWa6hc8YZmQz9gCyc2V8PLvzar1Du
r/P/A7YiIzBAe0SyFuPR7Dl4XGjURPIu4DShWP9xwm6U1Ld2JM7132QHM98Q+TVtK5JBgJ4A3zEz
bYAJw912IV/wri3rGwfT9b4Djyncnuj94iEXczi3aV7OxAAWXb+jU8R6ChRDIcMzfKnvbTm1p95y
6IS/0k+95fC7ds6jsoVPIdAQVI0euXTCklXVRRxKzjlklcQPWUju7Q2W9/ZO+EzMYpBQlYIbpEf9
qo+GURfQkthrHYw+laBquHJ80mUqPcucWWUCzy8CcdUGZtWA7dBc6NxaWwSbbbhOD4oEGVMZNvvc
6012okMdkrPy3ypNhN7fJIk2/jpi/res2Ha8Hp5LSTiQG+NzV5VKRWKpGm6T5EIJj1Dn48xGOGpr
mCB1X8lUDxwcUAXcfpQtgcmw9rCHmkKmRmoIdPYVy6FCpG0LOB7ys7HsU5XxBO28Rz5XRvvi+aO6
VtYud35h40tU74ov4idphUUl0CN3A80wSmRm1uGTs+uQwwln3BRhLjGPHCuUP35WsH7KSoCyigwF
8qSBv7RhTyxuJ+whbA5SsObk3BXA1JReAxvnrDlBXHAph/naTq6nU+0h75RMrr8QHDX3bw8vfIwz
baC6TwrzxqH6ZPr3J9VUe3UCALL1Nf/DegfCZuqved/Q63Prrho0q8lnjtaBS5rEcx0dJZltsf5s
SOv2KLANkQO0F1wXpDvNrc5XphrbMmMhxgkc3sJa4X/46S+m7w96rGIeen1IncKyxIvRJ738Nw/6
uXvuqxZAo054hgAhOYnMPO9xordD/XxaCjnPdrnZf9NKaqJ592/2vvptuzNQRaLGfyfZC0TsauQB
+8qDgJmtvBdHQvqr10ppM1A7W1MR2rYTpkkVJVNa96RmjjdnAjqKfRnYS6R/1U6/QAC6VXH/3p/S
G9yDKe7FtBGwxRb/66b/9AyjWm86tM6AaS6Fxwa+2WR7DAuUbpBbAoN9FCXdz+GJsnmgtgadxC+K
MkgqY2bJGi2zNFMqEgp9hmva7i9sG7tkTF7WsQYm/FanrW8maEmIynGotq6KNgS4aPySxsH6mrgu
l7b2tlJgEnKmqJub0Qtk211lXnGDeqegsyeDt2VLy664yfTf97Q8DZt+ccz9lksSCDyOgHR7/jEB
TmPXW1x+tjpxlpIgV7uGex0H/FyuRl88uR0IdWVl5v12BfsdJCKy8Q5p4VjhH1lgCuOPmmJGjevx
rxV3bh7ULcnStMWMbmDKkIsMzn8Tv6cN72QcdKYrSU3uHXcPLg6ICKaQBYM53uMLNP5g+9JF5Efe
yir9aSB+8Tx8WobzWJ8WF0E6uV5X1MGvRCVXEPdsHGYk4CO+94ywHld+Yyzwx5ItO/apEZ3mkMhf
blKB6pi+Az6rH+eSWSqsXlJGDFaF6Z53Jm1RyKcTg5sjof1Cg3vKP3nOYv2t7SKbi5uvBeg3ltCa
rN9DnEsEwcw8YaTKWDM/ZoCwFSDicx/QG+AJu9Ke3OkeYlc8/jCvjVxBu1+vMySPMUiA5SEaUm8j
fOQzZc6X++eXVXbn8myAPtmeNZG2ZinuR1KeHshmdwoTkS2J3H4imnC0Hj8vqaSWsvtjOipwVQfg
UxdMObaIV0MrNXE4VZYF7AGMQBUJlrEugut40REUyYtSNu+8i55idzfqZFB7fHT3mxdqFPWlgm12
uxKnt5S6k3Rh26SkTAgaTA8H9dEgmsbOKiCZHHTtJa+EdjzNYCkY0CW6NPM9c7oosHSZDjgnzIcs
DUuVlxldHQofh/Skzw3boR6wdSYKW/SaRo/fT88tgceibUdPa1a7SLvP/Ay5l0BmBRA52uyDv9TV
kyWuixrmSezUTZwwd37xeZVlzYDZPRI2EVuseP4iG/iKR5dmklQtr+Jc+oDHv5S2JKpi72JZtbPa
c7m46UlpGAaKTfIEjMeFkBF3L/twHfppI8/ijmO9vPyOBpS/CloMMG0/bz9u1oVkXofeLtODOExB
q7Pr7GBmsH9DWCiwAkSI+vzgHYGea+caH2wsY+ZZ678XDn7yPuihhvCrdV+tfuzWQSrBLCsTteqG
kBXLuMjGrVcQbk+DSCcccMXyswQugJeF3Fkrwzvl/Zalp82+kwdhiw4+g1meHiz5cQ/VEMGZWl4h
Rcb5s3SkvDYvmeEN1zQql3+r7bejKgrSpJTvPQn8C+As58BBq7riuyBayx4CH1X0e7EQ+fzVr+WJ
FW+dItr2tZbE72tY/X3/RWkDSZ8aWnGDqp7rdq/fNAFrCwypah73ZRnvXc2CiUPhcTLaXGOBacK6
LL1ncZBHdVfQZQGKCJrQL7blWQCFIBETSO1EbwnGLBKormj8Ev6Ib9d1SQ/0CgEZmHncnglQBiOy
7icAu1PXJLeRz6shZJ/9L+IZDGDVjl29E/XBG1SIaQOw1WSrtEFlw+NCsGwS3nsC1yUvnHyGS3IU
GhvVQn5jKWV55OvcbZR/dsliR/jVxzGLX37hn0qRK/j9d07ft+ULJ6gR4ing8q0GXVabcH1NqpGD
Q7PyZZMuHS5zJyZ+h+pGYyE4XDYqJv0KS9QUlMSOuj46+sQdd6Kp7nNidWhXLTHGyOthe31To9Io
Cg6VwAFgHiBxFVUgxLT8w+0uLmYCgP05ofFtwzivahufjIfp+sBNB0hLoZ/vfe1KyhMd/xAxBD0E
OsyYfR/cZ6vp5ebog0DvPKfI++4ljzYbvtogMkXJ08r49vbh7A55qCu3vkxD3cBqcNndDMu2iKX4
+FfgK4XFSG1ERvAwqPW2u1pAE4sE82mMD7UrdqNKx9iteyBVfsosif5wbmQubguf8s1COirrsnqe
/yI6zQkRFoDpkTVnWO3I6wpEeWKHOzSsu5PA2FWxEB77iBKGN0hjdljZUi1Abny9FHFjrrPwvZbv
XpaJ0bxSbLeC8U6S5sG+OmVEbjASvtk3zoSWHgp79p4Iwus0PaEkwaYsCFJVyV48vFhZV2/CDlXr
jRLlHYA9eII3/iTgGzviNjIm+EAV0dGMqeUEtxqdtI88nTalRYx81d1rN4bclNdX0qZgeqMz6Vds
BXpIIzzvsXj+B2usZehzGZt52X0IKjIc+nlpJ0Rs6OeIn+zujNiVls8Ln7fn96L6GDHxMWf8a5Vd
GmqzH/Zlycq0ZvJKW5jClsjfwm+oHKZ3h/wKgJkK90l1to+DnqLDFet6Uh6EkmGW1b8JGdMkB9Zs
xtPdcj9KySZ6DBDeBsdl75E97MB7kfOFNOHCxZJNK8UvJnokSNLNBpwZJR9BzwBCKPzhdw6/1J1N
+SqjAJ3ToIR67eoKevAen0EwYQbavsh0D8RverxwfBoPzmVjYPG9IsqMw/aSWdfDJxvY8f7aFs1S
3AMNjoh3hVFzlHrskWFRv0UHbZMaio+19WCCHBsndBUwKj8Uhyh2lIaDj02fwRRcD2XuPTLrYm5W
evIqnC0JP38ewcpnUWDEz+7yfqKd7X9/Tgd4I9bYco9wmU9l1ZWyID3G0mQYdU2v080UgJx018XD
SQzSM1aEKf3nUGtp8Nj18nmuclLIC/d1/aPenb7UJK8mef9XsQuq2Jay9DTIkgWpbLURWhjvHuR+
E1492VIE1r7KnlG57oLVyNZG+SrSQzkbnIAXxlgqiXS2kp9GFi2GANkWl2rlpyBQAGvRRS8tJXyA
uyBZYHgEjvttwPdcCvdYAp2ioa3Wrs73X10HMaJy2zwfgwfIp6uJ4r32XJ3nMRdiVFQn0p/2e1qg
2x3ciCDO9liYjypzJQunc2y9Q26fZTEqJwvKE3V9f77cpJzNkQpTJlaRL/gvO9dfG0iId5WRLzlH
OycpJ8r/R2ZmhTtOcd7Lx4i/mDeTTYTHks/gTB0o2urnIdS7Tj0oiUvgP2DQrXosHRIc4yRuN1Gg
fk/0P+XbSLnE1eeZj2iSvgMwFZ14YXzRqE6pfmmtf0sNqmuf73bCKEc4pugBWfbEYwdzhiZpns5v
ZQe7Qgmgwygj8U24C4klq1XykXuSQLCqi37/vfqVZ8ibPTtRw0J1VRSTvjYHe+tr1wmLP79CXAFM
zMUYF5kn2CvwxKPcvGM9F06BWc8pr7ZX4fk7NSQgT0SikwY8IhG54YmP0yN+/oKyoNmCP9cgK7nP
cgHTrtbQ6cLu8IOZjVXSUEBr+tMLYp4yLpeJ2zEEgLeZ/DKYcNbWe+AshToQ5mkQn8XSETyO9OxO
bpl/yBO/BXCgZ8LQa/Au23QvzZKALCg9tu7oCureLNBiak7PlmdVOzIj4SWRn8QSrRLg8tOvZvWZ
7XcmjqWuI3D8fnVz/svRAkRXB2xK6lkGRJ4jSdxvI/6bfvsmXuFNowTiYq+4+kJJHcCqQ3zBlT71
GcE8ZHCXKIgj90gYOIrb7XQTGB6yNS+L6fxVF1WhDuwCVqo1xCPOlXidufCp3jIt4o+Z0z7r4UX3
dJoEJaY+E6Um1BEQuOy4EY3JOVGM9WeUklrg62NMgG+R12lhALu1or4cevMz4qJUs9r3pVDCGesl
eZGvuePzaerBWgDRfXgTg2DLwqd562DP08FX2bhkKNiK/I8cRLLkyaZbQnomeo/MQbhiHMf15uEg
uhv+uk1SYTTEeITDSihzhGB1AXjt1BNmjvMLNoJbYgRYKesXxtBs+0mmrF1bdarx/PC8EyPe6Zty
dSNiy2WALVhwquwaaQvvEq0pA3WuneY2XGlwCSAip8PjB6w3yKOMyRf3m42R4+UlnfoJeFKN8s6w
McxyhIIbkBzD9Jtk7SZqvERY2ydryhXnq6PZZI7Q0QBz2DkYv6fti7nhVBLfym7Jgd60cdwKDgR7
ycRNFd2wBSm8Fp+PMeYn0Is7Oy6bxLk6G8gQqLgad4CnPLLxaJnQUQQiUYcvWf2TITpFINFA2odg
Vm6AMyyEEypV9yy18Xpq46K1UHYQS5wYBu1DZshmqEUXqm9bUpdSLgSY7+yibGACnI7KAUsYCORM
EUBXftRKjeVzP0Ed4spJdQlrKhs1SN1yAC3N2W2GWsjNSp0oaksXlhOLt/Jor+Z0t5qP2TmvRyVD
818C+Bnn9WZFE6DmFZWHasKK2Ws9hPBePBt3OUZTal8BcaLJIS+0IT1CovP7gnTHuqcS1DUd8oSE
prsJRLznj8T938QByi7SPFAKU8Qr33ef8VIaZV6UjdIFuyuM469n6CfYzM00i/Aor+KJFIpS1j/m
MVIIkXQ4c3ZForl5XILLd6imClsGtTEBgKg6iGq3ZgrJY2feAGKP56WDdBVB5wa/zfXSpgaCVpcd
nsiE5iQIdmC8QqDE6IsHcQ7SY5boi0951hPPy6jgzZ3sOibTxRxLHZQUkIHhwYpaY9QU428PUHmC
yBHp4cClCZp5qTQIy1X/MXVN2OqPedTLCZR8c97iKLD+SFliQ8oIhGS6v+DyoTHSz7MLYdUQaFHr
YG697sO9FUHJv7lmDCKO2TDhffUWUyDd9dZJZzjeWv0zEG8ljSGLkFzIj6o7hc6QKFg3tuqzrHXx
5NrWgW2s57Ls3a3efVB1NYT5CfOLHrWf2pbQjg8e0CLvo/RuPYXEBB3bUeCS84AJLFGBShK+qe3D
b6OkJd7v38Lwiu8ToY8q4M/OYHxqMNUN99UUtlKKaweJ1alJ+V91IvSsFZqpS9sNBiBynl3IWPI7
cjliqjd4viNbx/dELnn/4uMcRsEA68RrkAr8MYOEQ5FEKLtcqwIDti2ZRkrZ1Ut+Px+d+a0R9jlD
18EvAXkiCIxU2gfaZ64qT93bS9Y50e3pVpcBHHSQSaLwAen6XSythY3e7/vseeQY+KFj/hoKIta0
mW/6WPzw02nA0hbfB9dtx8akFC8z0mON9k9YoTykV9uOabV5UHMQ/lc7l/cPQzs9Pu/Ovt78eRQE
pk37yCg6cdPYC+0YtoRxK3H2OmJFmk2QUuUVy3FiLEjOp6FTKWVVa3SOEqGnu+ZdeGYeVJhe2v8b
oc/cxybnzNrqp5RL4VaOHfczZVlBD2+GBlRTw7MSJWQIMDTEaDbZD95efLweTqEKcDHAB2/ClUrj
opcIyrMKjvNlpwyUdpBU9hxa8TDOcGNyMCXN7LbJBiKYnl6VxD+ucqj4LN0aMlnEmYtOqJqRgDDK
rO5rFZoi8NOH8ti/iOQKlceC0mzkiJexFe/+gALNMHE3uWoncAHJYepIHbTlnZmWsZqVfSjQte16
2V4jticA+JgBwM3YUwDDOGnKYZOyAwazUTcp42i1AoFaHiJ/PS6b3spmG70YVXyLRo4vn+rrvuWe
c/xyUT9ncOFUo9ftcmlSXnvb1bkiI5j/EptUhnzI3VuDrupcfFStkMFBxWVaM3FvxddJzVv7dlet
WoT3O7HRSOhmKWKE/eUN1QQ5BYlkogfExEdJYUsHby5JpN4Ls3sRaSAa1vLKpg7kiomEf4BBcKow
dF0Nn7K95Yx8BG4n7QxFAuD+z7jXnKjvcL6FDO74nAB3HyDmILlxPeIsvgNAu7UgBWAAUtCEbvwL
+NJoLKNdTVBcpe4DyVTPXODzfBB1fnfNAc/pTy49GOTCw8umjfrTxJnDKYZ9CYhjAVohTR/K1vYv
46Ks9NlVEPc8djx6Vg8gMDLuIrqLkSH+DualL9eyt49uUQHwPRlvMtvhgd9MDok7fM1VT9Yh0ZZ7
bhCKnB/LBos5UzPjSfena8NSzEaJ7/4By2sANP/ih5WfCdX0BZYMO3aX7dX4PAf6Rb3bssenmQAF
M7KAD+Z5kTTg0qvfLCWpnY1Dw5t3uGhPz9wgpXrTFhINk8VFhcg1Qz2NLRKalzJE7YCRwsoKOMWw
ovYCmmvtdMp47oo+cuE1a+Rn2ndU/v+WlPy50mGrGqSxZQqTRe1r82spTcW6VjCNMyRyCDzc2EzL
05Vq9Mn+wInLDLtxHd2PTUIq1QeUZjZLxEoAoXVIXTQJDdxfzQpmsP3DW1UWdsbyQjXA1DTvW83v
I7NJlgEcftlYZ481hNbE8xSWX9L9pBb0/EVZQGd1cSQ9v07ZOTTZIJq5bWXTFdMFYL2lmqBWb2hd
iDNPQKSTG24F8e2jJ+s37n72TgEwGjF4x0kE64NhvCQnwniWl/CGZNiBIN3frAV/oz4xPmIX0Iqi
klRIV8bgf875MIbegfjHoarh3bzF7Ehz2+SlzxuUvcFZmRuqkMxy+FIqwGLY5gGT/n2TOvoUNBNC
6JQBS1MG5X5u2DhEnk6nBxGGVw9CR73WMkR+sw79W+N2Q4MPSDH8THWYrEQcW7UEeUBHd5GnD6Jn
uUwlLgVUlnGqWS8AkpZG/8xaA6RvJ/dfP+bSsVew28tTihX5Fq/v0xbwEXgBFohIFRPu5rgpy8AG
R6auk+IDUSZ4IejKQ71y2W0s08FkJo3Hmsf+vM/1WOF4JiAjCVfLjauMUs0l8ZGGkI7BO83uDQB/
+MxzUVGntxruCyPzfd91p7eKyAkMRsLalhL4l7nc3xDNe4diouRc8Xpy6HuoLc9Hv982BKn1TpQh
g6sXiq9fGp/kZFItj6XhiNUC2cfTuscIUgis57cO0e6fVBz3H4pxaK4s53w2YVtEr/bM1cpwbzUD
+6pyyaOmG3Evwdd0QJc2jsj1Mvk8M9lSm+R6sFhTbzqXvmO/sAknDP3TK5GhlZ6FBDLoWVe8q21i
szqtEuRRqIBvTy7bhVIkDSaCuSWyYt+woY3mh7p7FB8RZJn3rH7rSF+Yku8jJ99daJ65S7AYtUlH
TbhRuFUuoQgnnRh4WER2i0xnpBsDZ1AYp8DwqrJFGVYhGFhION12DctKrtmA3WhcQIl4Xs4Fuu0h
ocKxjNhb0O9tcV+b0ntUHLzgRZk1bf8tpYFaMZ5ZHnGR8g2qS9a1n8b2jpKjRrmt71mHrkjsisHX
u1/Jt/w1TjD/lLANCa/gZiUnAGvOLeTUXpayn/PXyLWrvvd48DghPZnsN98OgygPBjmCqcA1m6nU
/TlVXatlwKGU86iJL6gV4GT+qjUNE504Vydw4vrjrUQfPraZPU+cw6trKLep/HoZ8+jkVkiJyj3o
uPaEZ7m7S/9/BdX0jZiFDFys8iOGTE/Kk0RphZECZIfdaDwLxIAjHrGFaF9jaffQyWRWi1VyhWXy
61hSZW3Zft5y2V/p9Vd38LlgrMvz5BYV62V12Bn4CF3FPEc2k6XMUEjRc/T9GScXBf+vAZs+Jdms
3weQlh1HrIYFMTFpzJkZW2yiA3E91QKxk68RKhesHN3q2SwxtnHu1s1PPztocm27B7Ned69GaKiP
h+IwrjnMfPCt7hgDoz1m8urdrt3LbpOKZWo+qoNz0wJn9er/B73Qb5LKT3Vgyw/qLQ3sU28l0ZSk
tp9r23ZAwLjhWjLY7cXD1HjxCNrbaolxWMjobGoBJe3lif9cicqm0s3savD/CqGsR5hLepWMKNXc
fsa3V6S5tY3bfSza41Qk/vz4Z/rVvNZhixf/NpZtiGH9yMp4AoCN6LIJIMko3P25Y/x3oQfDgj3O
EvPav4sBw8fUqMgb4wGmzLeoYIOKYQZ8r5/fdfPEjPtRj6GAbJ6W16xUCtEPVNLhqyQWX2Cr+nbG
ZExYw3kVwf6Y+tnTwTRsFQh0SnFNRkasIqi9WauIT++oa/cV1eplrfQ6e04XB7KL4yx+6KrxuqkT
7sRp6HfWsnneZPDkIMf7KnOSn9Vnfnngx85JEpEAE3IYdWNkI5zpWSbZ5vWumEs1MTeTlod9NpaQ
x/lvi9s6QYPZoYXtsGYv+FVFDrU1Q626+XwiqFxNNtULJHeYWIw/im4VddmvTXDYlKfTIj0UXiFB
+K6jnmehqyC1dgCgalNfwuxqiSmzOPDItUhH6U8pcswn7qkjyAVwxG809yv6S66CZMuFvJntWf9y
33uDVZmBNis/QBDFhbb54S6hSiOd63/1gdze91BSBRI61jArH6+ORIxU188Pwc9GkCIQz0P6IS3P
LLgGvFWyFZZJxMO7DAn6AkdkDHM92deLfDg2Fmr38hoWtNnFncHnaitmXbyDJrfIaI0+Qg5M4cMA
kOBhltLQdVSP5eKgPJ+EPAyEDAIhZhWCwouY4ptijmE3VjXGCqOVz0xPv2C952VbFvo5Kwz+Okyt
KNqnvJMkMiLL2aOU0IXDwp56PH2L8dyhkbPqBbPUp/OssBJDRckl2xeAvj1FF7FVwnQ01vrTBlCi
sgu85vHK5QRrQmXdCdUFVJJ8f4ytjYH1JEqbD/4gJ+8+MjR330taJ0YsE9i7wEPKF7cNdLtFBxW5
t7KMNU/b9SHGT7LB6LjtpjQi7rmY8alug6MVkdyISRAZZ+5s6nOFsKJJ3SHcct4tTqCZ331EnMFX
SIcWDq0Wvj4OVoz9+KtNkntFjpNtTZfGXqb9ZsFQk3V7UcjZKgcm28CJeyNCtIzVirfxI29rtu7e
mDRopo6TlBcLMSsp1rNIHguLw9jeMTwV8+urg4drXYU/jKq73IoqWXYGM+pZPn+Uqj3zkCuyi6v1
0ocYktbGikesY/MOywf/1yG1eP7gmAsLOV5islzRrDORGYF58JR4g3Moc8U+GmX+7bsKDcjMRJb0
dRysh/Ke7L1S8gkfZxbLcbaI/rmm6ZskNWT9HIXXK0FLHT28N5D/qu1glrF0ZPiL4dCgwI2UOnUq
DHbHzgmGxhHXaGUeGlQGvCmai50agnyiwjmOOJlF78E5eIpVFuyI7gh86GA3iN3r5+R55fmHn9Eb
bbQfpjekEXRKpdNn7/jJDDe07zbURRuS3N2hM1cuVTUay8qoAUR/RgAy8RVDDEQ2LYKQpWFaE0Y0
E828e8pxv/674pHuQRDmNsU87GWzm7fqKYoJy42SXXB8xtYzpkCztZZC6Eyp/YOnB7M+q+oUtOkp
GCf+WCFQbjGc8UEJoHuQ3zdnoCJ8xVGhV/ihvcaxaXkqY4WLsRLdl/uXUWintaU/9mb81eM6waoG
BCAZy78hbsTHmM1EbtdB+IRhvHtk/Q0jQMzfPfJOK03cHNjT9BmX9AqTjZSSYSs8QF+4r8WGTUrW
rBqEYl3aG2nEepKmq4ag+A+T2vhVRlJaC5x31VqV6vnSsFOTG8uaFHRv5ovGeS8bAdpLOywqrBqu
h1Si1izQIXZWq6aIfNfxHCRvgG+RJjRSOsq8oHofh2m188MqD9/mC6fmORkMZ/KU8Id1bd2lwCeu
LRxYq06RkM1z0Pc30zKrOUvh8HD0+ONt1Jugk03FCWh7/xHAdZC6kR763HmbOk5uT/HtX14/x0vR
bY7Clsx/WmfxPumDBQskokthjAhyTw67X8N9bnK3derPtO7D1CAx+kHW65R7AUnzv/az6A62iIF2
wPN7xTEfRvqD1oIXeJu8V1TRMijrN2Of/OlGb/32kGU7piwr26sufYnA1gbpm0dZEo3cKCsiWCfR
VTJNf++F0Yg2IrSST1E+xrxMl5JQJZoBWOdnzTPDcxJNsrJQibeHQXgRBxZoDvCar5ibN4UHgfl4
tj0UVx/rXctv9Mas1r0aFCw0O38T/Nc6EsmkMdv69A2wvc0jzJSZ1vUGHP3c2/BNcQFDoL3Gr9WC
xYdFj98SqsQAdNbFsJUE096PrHVG3X5LVrXUfjwmU9gRjyiyiJm4mEbphhc36K1tyXqOg3sK5/AM
QRILFf0qwwDLwW5Y5RFVV5nBNjpPNu0xoDtR7Z4UzbntZmFFZhTxfrkl+zxvfSCwcLYdq5QT7q8P
82TfcytnhDmiOS/+4C/kYUz6eTOTMgP//+TM5Wpx/JKzLKgeXPR5HV1mWF13ZKeN8UhZzTSabVmu
jQDkzZa0F8x2Dztou/Q2Y0LD5bf6lsjra60iYhnWLu6QqVycQylG1Si2wXfnKhE2B5QYg2Yi85JC
65s9R/T5GyzfJtQ9b4TY2gbP8qw0Xgbo7ADuDOUbsAODPiEiQdflwLjDLO4cQUDCl7bRf9vfLLHN
d49pR19vCvDlGw57IsWdXMj3M/Y4omYWPpoCj7Z4Sl3F1oQYMlcMXbaZjYY+XFVVr6i6aK08yq3R
AS0RRAw5J743mkf6uJBu9HNu6eygk8gNxnCjWdrMFpTrznl8C/hv6Azr6yfT1AA62cLH7BQXMMNS
ujkQRTqMPdwiGa0EKD9QRPfwTcBgdWxdkZ/5Wu4XnBijU84HUMPOCXs+Ny/lrJz0UWmeL6623AL0
RuqkDLo9+dwRnKBgQrriuHdio07g/5nZzcvfYP3elMcBI/Qk6tSsnTMj45qrpvCK/8RkF+tqGK3Y
5JM5d9RfsbHX/kuzmYrIXBLXHCgEyf+2yCo897RT6Q37F1zzbfKEUhn2Y0Gsn1yrDyY9RPRrxhHq
VZR9n7Ck0ptBJrURZyRf/ghrV1GEN7WAo372LHIzALyTLT9o3eFYp0A1L+uXpNKP+a6QGH54rm1b
XVBp2ADGiEHDwB4Dv/cOpYYEa0S2/OeiAZrbt3FV/NCRjy/bt958CUnQlw1tb4ge8E6pPN0iDTpe
ZWU+tOlNXKkAtJwMcMoNUMCELvcCzPuvihZARuCi0rqyHa5XKcb+SEoCrXeM4rQE9wy3/qCqz3tA
gsba3RRxOBykO76Mcr2NLwUSPKKBrFIXRBZvQvJkHGBt15Bf98CfimJxJbWjpOdgrTJnXoQra7m9
qOqIbsw08d1gfBGJIYmfsRcIClKhX7iISKKEpYhYe1x6bd9XsVnGGPfYgd4c0lcwgRmAVmhTvEf4
NdM1e/vS8f0Q5unVYy1TOgv+TugE0AkR+rVSEROEDz/AOQMNA2LO/BszIXY4qJ7mBy4H6a2Xtejn
qNmlISjfy6gqoc2ZmsyqfpoK0nzW2qj79vVMOqhZ/QZF+F/hCiXwhd/O2gvYXWu9WhtuIS9q2SLF
VlbdRJEIj48o+l/CRTQ+AsmcUy8B49wFx0dzqmLKAWmI3OEg3R6Yt+PVcdXis0CAdGwS9pcWApiQ
OFzqfzSABVMP9e/uICh4RROhTT6kRcYDVIhE9nRU1tB0BHm+i7IzjembG9PeTOLWlrTmGMWGqdQH
BbWxtcoQ8pQ5R/xvsIgXi0YeFv4U7ky5Nfj0Xh0jhW9RVPeMd3marYRohSMMw+0yTRXyvxQCe+cg
c2Y+dVosbH+jvmSltGtWh3P7Wg9MX0Nr2+AKIGL06OkfUdfUzBEG+Y8J2kkDBTkfxyz4qiaYdqd8
MsgiATe9Th7BhUA4n02t2qikSz88MYnJqY73awxKCuz4vf1PoHiA6AnqZAixvxtE435cgncXDhNH
J1FeZH4ALBRQecqPFZY8epSPtd+/Q+04ZGCphT8D4CFT0cWtIiDP3zJqNzLqGG2mbMUwpfr+ZCuo
KYS2YeRaKvoGX/LJ2fcKpSkfjXJlEcIpjtns/ZNDLqkAIhOKCt+uz8bVIzAozdO47S2UJVPdVGxp
40mbCiIzhlkgx4vHOoAILMs6H0yRHDYtQMVwPlbqg0balf9qgG4d+d6AaFjIUKztIraVzH+9abvj
RYwE74IoOlETe8nfITD9xDV2Xk96o0Q1rZKqf4PA3/UcU0cIiVBJiMdR/R06JtoBCQpZb64kmOAv
2BXfW97pfRNHEygNeSlsox7GZCoDHP77JkzD6B/s9wQCCwMRcF/PKOobyqatOUBG1hfj/XFzE72n
jFbQ8Gn50sCYOSfM8ZeZ6SuBSH9zsMudIb20HXXpSMZdzjFaIp0oTM5DIVsc8ZarQC8l6Mx1u5BT
Gn6M9yYPMXV2utlhnTIS7EPEbADqHfW3rxbNJkYpvIPMYfM4S/WmQuO6Xa3r3zrcMCbm6IQtAUbQ
Oba7vfkKQWSPHOsuA8B5gzM99AqUPS59/ZtlAOPaTp5Zo0ZK2ggizC1eb1tXK4AIn2zja7Ao9ROS
LbOSGibQ5co8hZ0EeJnlXRkBx7uK7YYkH95XdeUUJKPFaC9BUdbplBp7Vw1MrH15ECM3erO2SCWd
gh54z8E4dhnAhfd0ep2bEeOhXMMkskKqxevbP4c9saCfLHolEHZfVoWsLmd7PDcFaxHJE9nu9PUr
5nDrUsbOGFLnFRgj/USxD48ruu81qz21sMF6MEjFBKxSgz3gaNBWwE4XnV+wMamrcSnx0th+dIkq
S+kZGknAgXrdB/kqoeOCEUnZMnmIT54l3IGvCdsNnJmhxLUkOuYHSowiQPReLdws1XTFkblqQLzN
tQHbL4KEfvuA5BkTMe44rg1YUn6H7PeLb9dOJZngb5nAxtiLUjRW6revHerg0u6Nl9I0/Lw4Qm89
R7MU5ZK0IZStd4WkKFlJ0apXIe3dABBpeIZQnHOQ+1oJuOdnmD5ejCHc6+NinsfxEEL6QQMrQxss
O5rbZdmm5iZd4WVT5M4rSTX2eMJcTZ0GLadrilwvdduOBaPrvOcyKAhtAfk8ayjesZPf4b7pP4AS
VTz/ipC+ZAcoufznaLVByBib21ihSspieyzr2x9zgLEzVbllPXph1i3bf9vGGbAArXQl/DY/HYmA
1aEzMqvZ1ajY5jfwBxXhK3zH2MzXZHwYsYD594o3WoHgLwBFZGUdiRCCc4jX+NZRT+KOzOaSLvWL
1ZBrZnrfEinSx43IeBUqrSaKpSxwTFOwM1Dcbfl0AVlu7zzJZiCvI31BVQJvwQrIOg/OwHhLFf2v
OfTfe2f9+QLb5GEJuOwKPa+JIcseDe91apRncR6N7xLpUOqYj8v8Jpr6eAGSmFBOcql4WusbRTuM
iV4Oa+qpZ1ntYtXGYdgZUZbQMovKn4cqlWzuZpeiZY14cI4H+WaLzLEc7mdVm9dtBJC0vT9Rxw/L
LhxOYlxcHuPJEDLj+rr+j5Ex7FyPhsTmB21536Q+usFwAg2iKWCqh566SNJB8WfpZqarqyQ7CHVL
8XiLfn0lMpTUIVZhiS4uuK52umti4LqPqPG/KwQYkPvQJnzYMqM8+/PrIot7sZ4TzyvlD5IJH07O
SwgfzA5qtFFrRWtt4pXxltruHvTwLMxxB8KYB0fEZZLuKsOZjWMxsFO+TfyLDcI2ELQTBFwFc5XM
TErAbbEi0PnMdXdaDsJvwafj7UqrgmGeeamcXGgql66x8YMY2yUPNqshXmjmJBlf0hGts7sqouGv
bDEHVI6mdGC74+9NToVVrD7LwVV1Z8mwImHzf6+XxT4M2+cV/BKDRxqTnQAkz1tNLNAtfFpNqih8
i2jnwz04E+OT22kqvZetheLKQSGNbNL2W5kXQa8YZ5rlj7T99FB//4VtcGJxN3K3afEMDO9fFGLB
uuHMPWLoTAQWOXEKtAJd6Lhs/dNxq0qDzJNOo7Lx5yAbVw5vacIQgtaWm2s4fuQj9IaYBbtfvUw8
BtnDGp87Ff866xuqAxdl6MOSK+lI1w8eZKsYcSqF9nDY+6C/nIWBySinrejRx0kVHtJmJ4dBKsVi
czEaWC2gEecm252rzrR0og+00Rq0V5Xtypon55Nzjx4iJmvYHKDswQwLYM7LmdSeep9NL7yUVsWI
0ZP/axa9RWqRRGiJhW2oWXpMPE497yE92n3jQn7wvDY58+7MrFBsExslKC6UHgnasGLJyJsKXaOc
GyJX3EfiJm6BN4qg0Ww/vQaQ5VMVar8H8ONxSD/+qbyCr5S+d3xLUdMi3ROzN7HYK7n0AnUxFXRh
X19/YtyvEt9sy7hrhuV0q1DHCkNUnwi3Gcv/YC95oKDt3k3wU5kd3uXXv4T77e8aJtbuDcDupPBn
IzVygonXqqlcLekFBUO9LZwUIXBKgTiy29vHDTUYEKoN31YpsJ4Rp9GzEr6x1gw8CHSrgXNqfd/w
EeerRHj82thAIOnKWlCKoXRYJKpqBQA60CxtDAIV8w6/zewpDrBBuVtQt4E4mutnRuYNWPMy/opF
fyzOgO6TjtARDYQMhvMtqG2X4XC/4VliIrhqsUpsfNZ2GAuSQsCSY50CK3SXWesrj43zf+k1tnYi
LS9hkMzop77oWZRETDSy0APmNbsT+geNaO5cvhifjHKKyAYrPPxgdQewPfBQE5vVGn7lULg9VjfQ
0inBdpk4fw2YYac7A+/xqd2CLiwmVigLXIH2sfGGHtbYZ51AbUxfGY3cUVBEzcfDsT+GfzLMtmSB
SIPCOgaCzvMqPlNanLalmv3MD1WXMRn9GT86Rdo3VHD0F0/V+yseJh7AuIJa0Ak3yxHvqh/F5du2
nohxu2WrK4TfBYIrZS9jfxQO/HoD2H+78cwEdZQ+chd5BvK58g9cXryaf00RYJnHAstbPwxI2gEB
jmhs648AhEcFPSq5wi4oXOAqMkDkn9KqQRWN0+lsOM3k2Lncc0lGSJh14qMLwSuXY2J3KgHbhOo/
ElasYNWSkeTYy2WJ0LlD7NYvjze/MlGppjhuh1eCmpSOWudwaKxq7ES83quGQyh9eEWPhpvcRDhv
qDU2gLftxyiXcMrtfE4vENOxxNIy5PgsKh0qzmsyXyBJJrEpQXWzjshIrzHHwqMdWw78lKA+RqoP
AewIYhY0Wk6oqu09TB8tckm3PlDbJ4yUEbWVowtQ6DxaQk12NiVLq2c30nlcXpH7DuRuCcn2eWi2
U5Oh0hFWYUI2CDNplYUAsvOb6L8kKCGu9nJ+tVi1PQNAlTzhHmprgwQRaO0FpeoBpD6RCMOwzmVr
/0kkhkj+d9OkrWMHOtXXBA9N+wpdZU+38AgGVRMVMNe5izSVmZHBi93kmEcKvwutlAUgc+JtsU07
Fx5pV2nAD4QhltQWIg5ngBzzmq5Egjs+obhqtaY5KNTRB7Vp6n0vWUEeky8rKxCmZuDDfl14kTaP
GCeYByIrvK+W+eAYesJCcg+W/yzk9uTH/hmvkZKUktAyj9yai1RSbekQwIJtf9orARYXZtY9jkEJ
xjySX412/7i2RjxjXYYcwaZ/hKEMVYzkkdzXgwPtvP0Dw9h7XjYv3C5tjc40WbfEj3IGYameRDC4
nwCpNn0rrmbusj35Gof2fy6/JSym4YdnJ2689dT1Jphc3shBW1oE7JsffchHymUqVhCRcr65566X
v5jqp1gCo9j67JE49DRtArYZqVZlEeViT2C4DiPKh5JR7ebcZMQs50sexJBM9p7AwsebtFlm47Gy
pBCCXdwIGTHLBhgweq7MT/RAoR+b+1atvjWvkmYH7yfruHgb94hEDomoIBHZlZTqt7Dg6MKXeAOp
vqONLxXEHhkyDkNNTTV2uof/gXJ1N/1URFCirDfb0y0ql2x+stIcDQ+Xx0DOXh79rMIWDQAY8sv9
kMA2wToiF8Paeufkkz4QkAwrPthlB5XXir34KNPumd+el7mmK/zDHP4y/ALPNC2vv9mU+BOJHuJV
p6jKhDAAYoKNZ0Yt+f7ncqlsFBT+175nkCsleARiVodVzN0hbrg9NcAgqXjzr0CR2o1/zG90qMcz
0/2xLOnIfIvS54KQCKsd2/m0AMrvJvtO+9LsGBbnZUO5uIGzVkiviK750iiY445iu/sGmLQXn+wo
mTV44Jcc/IduY5SunnzGEUGVrxiw/GR/slQaA8CeDuIs8KS0qagyd8mNCi4sioHthRq+x4XsDhrL
re0JEd2nA1WpeLYC6kbOmaezWnlhkLM8BNEe9XBp8jHNlU1AZfxXkkMWaik50UGvTkkOfgfvyKgX
4T8GDT3B1Z8Zrj8n8VvCBaRvfuNBKFFLZjXobmnHleKDODczeh4N3ofaugpLD8n8nq1Ipy9BRTSd
GNxkuhGXIA7dbf9++jtw54JZHW1qvovpifV4TJ/Lu2fbrN5vo+ilQc/AvnyCJiELynUllZCcNiYn
QQ/u09lKobnrXFqxS9tUboHgyOE+qSdVOw9+WRHuuaF7qW4sqXS3ehk4x/Mii0fPNFgry1JPRpva
5Zi5GCkV9H5XqPckFpvM03lKAzQ7aacOlyyfCfI5UudLNi6HMA5sNYV2aCi1oFtQOCRHgVY7q1OV
bHG79t4nfG7QTK50fgDs75KDBPSNjN4CXDR7SJIP/4TrgWIGQLKHWzWLX+6nrbqOqRoz1/GML/R/
Bxm+5Wuv7MKHY0C+2ie8SQVnheTHxIhe//Tmv0ikN8GwfQ8Tk5XX9+iiprQEeGY7n9QyrXZeHYv8
8J0EyVEpSBLWh49RZFU4coxAYho9GlTPfwHvGQMncE7ERJRmkzqpaGQyUyYZV/aCnewsPsK4R1zm
pip/m7/iQCxKOSQCPobQ25ee7hlaIvWDLcRsLS+93ryw8cW5WT+50c096Y438rzgmypjd3ptndxA
oPbFQ82sEBqHZSdrzxbUJszdVzkKM+HyjXdAcXahUcM9xQOc0eDrNa7YhocXOagmPvDyHtIoP+U2
y8SnMNZIcvuTV2Xky7EoEX5i7zgxrVTbKgiKXlsEd5myD4qUkQwpkMndje3yzpVOEwOMzWV/7nBl
4LANOkXKgx/d19b8hwjClfHoTgWPh8lG+8AOKoWU7mQhrzeVnlXJu2AsXGqjteMLoZyL8r+Lbzrs
sbeNLMYTEB5Jb2eIVy+HY9e44HrxHnzew1U//iYH2kn+OnYBiSmkF5gy3Mv1VWyugTrnqfcBoe68
Yz6kwhPkf/G5/xBe/WD0V2rFSxHTSqSL7H/pSEtxY1AmXqgjpgnrIT1VTKYBMkCX0BUngb8qykkK
C8FLjMyNBHvaEeVzKJb61wer3WR/Z/yVQ3wMJN55zxlGoMbh5Zo9K/gbUwIkdvnY9XJ82mxnZVB3
TmF3OnYK261ycMI+ltfdzhSr9xq0ptzz/rRmY+FUW37oSE3n37Gt0NBHlNQsq+9naaYJIi7LLtui
IfpYr97BWijEsGVhzP98CIzeTHxlu/pIbtNeRJrMhVNOYN2ULS++ateslt39hQ5KlnBFV954EVvx
nj0KifYHg9X9yaBJwaZ64ePgrSZSnfALKLFo4aj1vUcEnwdacmeS9JEITe339kbKLZTj5IWITC4i
x0QWvZXdR5bxTxtCKUZ72ZX+YAcVJCXGwLCRenPm9tqAiFIfl1TYoqDRPZqvFPKIr8FXvxX4IrQO
u0IkpV11NOr+vmcn7kqWm8hW8Iejv1y3giF6Oz7uu9/6X8lBsKNeFNjvK+VWXbWLWFwL9Mnwo867
z9QIT71c/dyL7MXdG8gBHCPyKNAiYuIc5j64khnijCZonYFCMPsEoiIkiEqRCLg3m9xjPGXshsVI
1dKr4qEosI6PHF8dZGk1V9C9vQp09UMpMOdAcpPs0RgMBiIKtOaus3IqlDzL1N6hTHNP/TFknlje
bPqlHT6na9eBBHNV94HqUL9VJnPp5gpt57x+6DFi0dzkVUkQwX8v2WwQxk5sUW7FuO/r0VzARcdE
WqOwnqPHntbL6XD9PyJl6Z5R7IkRXnw7/OQdA8SVdfTkdOvrZYcwVJl81V1SVOoVuak54vkxRzJR
OPB9Pzx31UWN4oXFXdvsByZDErzbGryeAbrlYgj1xCQglrWglifRv1kzL7vYj7x61sFQOmOA4aZ3
aUhKLz/kEXjX6j0OFRjD4Hw+47uIA/QctoKLBn2UStWTUEfrISdqBCrtFiOqWnP/OX21p6WgYURx
u3JlC3hLjXyyypSMqzAwLCiBKs/5oed48raCOjsgEywfj+0PopCXU/k6q37N4RPretqEAWcfaRox
oTlSmD0sLq/kfVZRD4KqC/lDTfk8VsZ/XoBOm1OuuWSv4CGEpvG6+dZ8QL4RrMa1mWjLlqy3vux4
5xeCafA6ceZFi1FV+7EKvI0uAtV6g4hU2KAw2/WSYSOQd0TSxgFp48GU3SIhcYDLeVE8hMXpExex
Siv+jJ7S4SX2fw4sHnLlEI0McR+7BxVudyqvRfJfCOpcHGufoG9ER5MHVP6xSBI0K8mp+1PZgdKq
drV7gYlJo1eqCoqP7FyDuMZSFkXmGo+Qx15BIXwBeARL6UbBk36F0Xv6IjK7739Ww4+B97k8k6Zn
bZMCBehw9a2IZ2mmZvG+J+/bzoOIdslpHxBTum9gnYPOIzEydFVKQSYuL5cBZI+57l5hLngGQ7L6
J71NqFJGPV7kMxpFVvoA66pE7N87tYvj94V74mSgFJzuV+yb7RKVbP91XaiErRgkGbxlqb9RE+4x
gVZr7A5rGEgIqT3Xbde9tWXBTKXICDwwCEHOd7nra7DkNwX4UqbxnrA2lRjdOfupk5HXBES64Nf9
WZl/rfLlM5Tl9K2jDsskx3S42UlGykg6ZStn7enpXNfeStOK81/vhJ2g5ydomXDcA+KaH5nTnaLq
J+5zr0lnFJok9PjOFldXLWDqOOuZkSBYRC1IzMNOxDDxdG/MdA+tSYiJVUdf8yLgknvyD8nWj0AA
0iKnIRFtATlb1AyG/GED7yaVN+v/rCBBQFhFX5UTuh60EvRcTmu2PrsCNnWuxtQOs8u0pQG02BFD
7dtkZ0Oq3lNZMpVbVvE577HNkeWfHFKxNb6gCpIT26EkPUEeNK6o1pbDHvqfbnIZGFl16mF8oS9e
9wTMbi2KMJ7iFV2uYGVxZB5TxNe/J0hFECGWxpGXO5+Qm+vwvlV6wf6HjpZN8bRcJGP5afsAveN6
fZNQX+zZeUrDJXGZda8bFHksfgYjPTM5r6frGWho5HabzYuCnfxSh52oYSFmtnP1kIz5db8iaxlH
3qnTJHUw81cWeu1P7QbbycOtO2TSxM1Ji+brttMINwPC9LhgMWsrviPhlAhlMMKuTdcqICklLB5k
pltYoIivJlDN8XGnj0MyQN5YfcBeE/pyfJHs0Ts1VOO88kD/e7eueKK84akECqGMaUqqDW5BlQSk
cTj2ht9RsG9LN/sKr/1P5RBBnSb0QKFI6DLoxPB7mkvYfSATRVW7DFN32If87bdB0rsLXTsuQpI2
9BkbTiKjsZRNIY55tF2q88U8RCo+Fm4AVC+B+fs8AXeSCauOMmBmMv+QgUoA47oatS4Tq9FMmVNJ
LcDzM+nfK08jiF82SAmK7W3Y/jG2Miuo4EgnPj798c1iBkQTRcq3XYKRfYw2WN6smCQsrcw3NfsC
TTbNTr3Dq6rao7MueeBd4fEVdYCR/2/6YIQidKSqr/3Km30QYcnWs9pYCHqkyuqOyuisevhhxSsW
+5BF12dDaXZHjTA2EtzdPMKXwX3qbI6xJXQzdV5kUreZiweqrP35paUUKof5qtdHlVp8ULuXLwbF
mpZE9yZA7xRDUKc9uAF6vYJuQHuR1caQJRhM+vulnjqjPz40y5pBOBlh3EjDghUanXGgslnIjp4V
za+v4Si7BALmOaMWJu4fHcAg++xrV/3gKaCiKYyq7vHsR4k2nccg78zj625ldX9DXvEhJPn0030U
MhwDvxsmF58ImYjkXUd0x+ATzwNqzSGGV1uUdRaeaPoiLsxHc/T8SuQjuvNZrNZR3FPnRxDfGX6p
uMzSPXLB9KFmN9oZiYSdlPxF7R1jeNZO+MXYFH4m4/XndVaY7Iq50VCgQF+AD1YeX8BnyI0LIP+X
TEurKy23o3ILU/Sn3z59AGgU8Ge3MDYN0pqucXndx59bStDEwY534ROFCTCfgGvoDAGOcDMW8q4F
EUXEjuysMy13VUif6TQs/yx9NCV4gMamizy439nVyBmifHr0SHPgcPXYQC8QvFoqDvncf92vH9dj
2T5isheAcfolrdufsEir7fwkRyp08GZ+nU24AnF38Os0T33+MxJQWE3wevuwNXUvRysq329opc85
wKVKafX7HALd0+pjYpoclErIEGVHCUZJXvqRIDBDrN4xeRiC1SJb8jsV4j1dH08glfSP+vqAcATS
BAgQWYR9LcO2yOVWLkirXYfVl647I8Jdcd01RWXLbOd8lR+mkM54q6yMkds6H2+yyEEFouB4AeXg
12NEJFFNCzAo+494QDOzUtCaapQoTihknh9YcqtLBjxMbQC6P8SnPPcG7NmCub13k9dq6Ap05kq/
hYoKGbBUmBAP0iPPoj0qrnPiBFyMo+DZT/FeUdihh9R5LpOsLkM2YYjF4bTuRSsJdtzZH9oH9QbF
hZUzWiE8aGjiugLK3NhfLlx5HdPLLIYjf/Z+UDdbqQljdnRBEpfJlHn2s1IbF0nQ2gf9dsRTM0+0
6JIOyaPSe3OgvbyEbfrsT5J4clRgFYuSMuWGrzjzfXLUCvYxPvvGameXwhMlGSAQkkwcZSThow3b
+ikIWJv0bxvTDZchPiPboAQFIgvuyawYgPqXUMj0+IU38lWk+qAFXmyXgNVAZqykExedvQ/QkIDj
u98uk/S3dnYhb3BCGu3rHc+RiIg9spas3JNAylamLaZNWrpjCFfY+QWxnxIGmegKSjwS2uLFEMPg
Bg2jiarR9UZETw7XCEY6P5gm7eu6gQb6XnFQkDjxu5bSSEvjpu7OD61c49AvKRPibifY/ThLwDJM
g8O4DT/eDc1pouZRJQk3v47M3XLhELYtRN20HNFQ0HSrlas4bzcFXSqplsMt3WxD/t39TKCURKmJ
Zdvnb+bc/bqq4LVXuq3y3g5gnq/8GRC7xGBQl46ypCf4QCkRTHYjjgVmpPF3TMFW5bCOydqx18Hw
nWV4NJYjfHGB5YzDG9wlgim0y60VMfqV4zpwsRQKKdFLmuN1bClHv/SGCwSDEGpcL/TnQygVG87Q
mMm9ULdIvgdLFjB3b+iYaI+DuXgBkrAh0BWtQKfqQbJY8UndyfSbUEQo614X2JF7IsjzXAN7nl3v
wEiOFafv9WRmm/bVNeHUd/pV5Mg78RuA3bWgugLshq/7T07AbgrDJWBc+uW2PAcKGV0Na9Hw8csR
KFpeSUEF1H+uHllEX5AI4nW6X6xUARgrjVs/JMWf587y/VQUc3fGkfXzx6bKOtqG2Rk/Ul6FBfcV
lgqSyZWgeEuv/VW0S0P/+sUSJcc53dzDf+FNvbcW6gxYz1h3vOQDOtG2XfxNC6KzobJwuCiYUQsW
XeeYFS6BKqmVFBeyLEeTeoUpUDXG0S7UligHb7we291riyyfxLiuDkcPLrfp1o9K6mn+MkUDzpjj
FI1lK40a53BzSxr9f8kZ5+T53WmZ/lCJky2tamdhq4CvgzoBnJekkX5zuonjugtlLyqhsbEsju6u
5xYEXFRxX0A10Vgb9ZLtW2msy2oPH8mjeQqXs2di5Lxcs6aSaFUy3vsGAFePyWAmImfueiBemqSd
sqBSKxCG1HE7JGbFoNrKjW+SPAq2fDHTh9fnCprpyxoERTqhL9N1Shsyh5iPtN7UAdbzP/mPAaQV
5JMRqgm5LC9xVOcqRTVP+Y/0hVZWLwJnuBi4C6yGLlQiex+g/K4Ovwd95FGcDZk5P2IDLJM1nrwV
S0gSuXQcI4JgydanNp4OdpzmRjSLJ1IAEXrVLjbAon7bmo0Nv1JvhoSCfyPwXQcP0F0nog6jO3/i
o9z629kylYMHjYaRrfeUFfNsl82x2PY+NYHOF/DPmXNKx0OvFjDkRlAiVvSrnIj8/S4Nc/6eVsOP
0H4QHMOrqABMqCBHb9mEZL+aSCvDnhR84czOhZAr9jDnH1t52cX1cFvHX+o1uBFBJFd5d9XzdrOF
rRp3n6e4ZE/mEieKJhS44ELPVgwqAyeawlVfd5+f+L2Jyk1gIgSqqCUCxBMIAiz8QfCm0muRcUV6
kBwm0gc3/HU/NvwQwVl4gOQW1ZKAuRhZp6jg+2Hu4fZ9DuTTPG+dCnKdpKk0nXgiM+Ux8W9uZ4nt
KSVNkiiB8ltMNRz6E3Eg0QnzRPrvPWiaJbjuUskPzjoW3DiFZlApRZ04zE/74jBcqexKHu7+UfIB
EIQULr60OfhF18FWm/qpjJlfEwMtG3hdYEhzoY0O22CvT3Whod/+CiF60xIB5Vcqn/aTYQWT5AvU
drm/po5wuV5EePuHU4QGaKab0pHECSvOtVWz6llU4w0FmWKazIaEz/1zTP1YfJzWRxTmTzGdsBI+
tzxwhiEWKXpQoy7D1YYW5OEUOwpBmXcjP+iZF0UIFrXUa4hq35dIF7p3aUJ6NBJ0apcfgtwu8i5Z
TGnYu/gsfXzFSR7K3KXK6TLTgnUTM22P7xDysKLrmBd2m5FC26PRVnvVA1KAW5NEYf2eD/frMdZp
GwO4g3ruCt1TTYyvd6qZ8K5UKCTu1CnyHV7uSA+B/ZW6AiHoK9R5j98dOD/P3vrLjm6Z52tR+moH
03OKhPhDHrBWeJj8IeZ/Ee3lIA0EcY3i/J+XH/7qWePVI24CGP5iSGDpf1rc1mntcErG0PyhJpnY
lfe93Z3ommRT4rR1UTnZ0LR3s77pVSQ23v83ISJaRvVnWwCjU/QIFum/6F2n7+sqlqooWz/ijBST
KV9pLU/3Ywz0JxB/4jxL7cHwy9/gsjuew6JFIhZpKcLQUQndZc0D4LcF3zMv1OWibRxi1G0AgBIs
mUPq26S3tucSM80CTf03CnVEhFFIo2xSky6v6qhihscxFKYexSbemY5YYaAP+wSe48ZYVZubbhAT
+00rPBanX70+yPeCsbRyB22sAsHl88lHqboySuVkI1H8vkehrcBvPSS5ymYeUZEunaLdczAsGzTh
p60jzF/7EpM+eY86iIximMUQ7VUEWEKVFdsSkoOvkO8m92zGwKPwCSUED4xNvoi48jXsphFcdogH
KsJ7igpKlW81nIkcQASsBWPLZK5pNMuKuDT44MWXmwsQE50sHZ5+jvy9zt1JrIfjwJZF3PPwthtv
QPUrGbzUmry4tQAerH3XxFtHVGDUZ8dPDSQA7HYoB+2Ygi3LauT6rQKXtc+ZDH2L2H551n+Tkzzw
xMv+W3u28RoUg1KWuQrpHlt+GdMPXwopCFGkJuU5DLD9aYmow6oDXfF0pRRGZT+y7QGtkYwkSV32
vnUVPeHdSKewUURL4sprtveE3YeHJlc8TtV8I36w+4AwNLE1f/eKxafhOQvY9N/LtiZlYr9x4pLI
iqwePd+PDpgczmIiBw4ZJQkxztmc1DoSpe2v3Gp1CfuNOwA4IWqjYreuKBGt9lYHW2NiZfE45hV8
smbsIMD+Uy08phW+XidxXvvA8NyLSiOlIw3CHRtZhaQuAiOD9RlMoho+xdfg8yKm2EkcP6Y2AJY3
nF6vmuc0CBFJziHhcCXb0vvp3PywvUIxvNeocfPiD2J7dCA3pkNS8vXTTqvf+dbelvmkivn3FwSZ
vl/3mwfM7/Q14gtL9lwRsFQhQjxhC6/enIHXuXuNmhQZyjXf6z3T+zAJx8CUk2AWk04RJvqazUeh
1Igab15SCk/rI5tM6K0Agh4cF+JSo8mfT1CuK22vHSzxrL+MAMfsWMn5s0f0Vu6HGz0pnNch2tjK
EFnjd8s6JNmHYiibFI5x7VEo35ODDySH5+W9FzPVvxFjk1/R7brPDmoWnftu0iA18sWvOzQUR8Q8
CT5RkYzPW7lempZOj/djAaoYdM6KdHgLDTOvcnx7iemuk6KmZ80kEmF+UY2DtkmySYGmEH4Ljnsl
yn6DeIecX/Ejw4TEeBf4W+/uWP9vZhsqLuY7AccyHAnxs/EoSRmlfZc4dFahjmpknlHS+lrxaGIU
S4SDpXGdLaZ4AQmoOYsyyeBzuFW6ywjXYZuAw59oG1NpjfyXcIjUeDzDFNckmK/A1UFSNIlaSZ8e
BSEi1xnOS18rhH5YC7T71IHIFTE8LkhriP6D2np37DLpBhY960SLkZREZ7yjqn8tsrN18vGdEXQZ
wklAlICIULmOHc8NAJ213qve23zB8DFMr05ssisX1oRhHUj76cXAmlQEi8ZSw5ISNr7XF/UV/6hC
c5T+dPqrZNMk0CfoGbK46c6S35tdnzflH7k/s8gm5Ox2ZUfFnJ3OdNBO0BZ8wjmErRFXB/+uAj1S
+FXTBwYh/ivrq0Db7ssj2KiCyEvU9ywM6q4jnnZtOyhxLGUMQ06UwisgB9k/Enxdam/B62kySnXK
TsorfIPWLjsma1IbgmNYYTAjMwp+B6lYejxvbkQGkYyx2iddoicIOog46zLLHFnaCGJB9d2/EJA1
26vug3han042R0mC3QcKo1GqZcrHyVgWGssJSqM/+2p+H72x85t82gr7qpv+rL0Rc9CVs+L2tkyV
vgYCr3a9INRnVLO/1x04BInp16wlRiKvFs2S3DCefaPIsMEZOoAf6ZuDNiSSMBJlS06QS9Y6vyAH
D6lGHOjE0+s8iAYnMFpcjqFjEllMCO8oRbn6AoLqmvgJNMfG5goPEH9J7QHCoQebBD9Mu9Mt8dsu
w06PGyDa2ZrMUh8AKbS9cHi0An0vGfNS30NYABKM+M9McLeXrQzp5Wbh34SyuibfXQ0UZ1hSTxe9
b7wBeUcMRL4ChcRgwQ+OU1VwvoIy+KM1OiJG11B3zQ7WZwCLI4MYBcV08deaKw0Gg8/kSvBgPOHJ
hvxOjm5utJK2udAjRXpueeM3+XXtetjwO5bbGpK9PPf3RrGnRZEOuOBGZ/m3RRx6lYrzh7i+LeQ1
bNLbsK3m+gpOrzovKah1vGV0En83CHpSiKbv40snpfbd5R1JT8QKBF8IqXXD8yEFPevLZ+OA/6N8
7PMLJ9OWZD0BGxkwz0wb9eWmNqjpswUh3ublUK2+lgQNqaTBgRXtfEotVLfEM2QIBTkObkA2CwXg
0hggh1alVLePDo1o6K/5SxuC8lw9PRi5K3EVew9zIQuSb/4PmUGABMelqN6d3STCV9JkbgRCgQgS
eDRSj35GWtYzd2o44UQNP9onkCiOV1ucfgk+8jS0MHCo4Tf1Tc328jxxwNfV6l4e4V9fKcZTMrdZ
mqRVoMSjiaHVCIVfeYETMu+OIheYZ4Sm+T2ePj+mwIiXka7eqr/J6F5GHxeOO76Jz7igrkRJaCs3
FoaRR1UXQfN7HLcjKG5jUOsw/SiQh0ZC8cLZepKukYlJYpopzyeorWomG8qyPqsyTbAhGDk3Iv/e
hUTek96vBHcdDBCc42QJib48KONsWLivz9nGlgf+l5aKWSjzqlBlbFaNuQ6Rw8Q5fg3Szhsvya/3
krsZn2IalIFSatPZ1ugLM6Kvgr9Hm2PxvRY8FNeAwUthkoRO3rOBrLjPe6MejazMGxalATxBIEtK
VCEFcl0zKJ0hPlSJ2mdUCK1kau7y6aFHTWsJwTms4k6wocf9itU9paN72rP2VJTwPCQzHRAcPpT3
42fnBBpjV65g0v1n+Epio8bxqY2GIDlX+Lcek9hdM2VyeJSxS/Ltz0/889ZlG1syPEGJ0if0uvv6
HhhUMUEOmFPEvPUVeoKnl2UzbJj79Y8F3CiQTFJ7OhS307Sg9+/LliF9T2waaA5/V9LB3rFcnPp4
WXG4d4v4Xao6aQ2qiWtawWejS2zH85fDt8eFOllHULbEXC2oNrLRrp0ka6MVO+bafdEFOx8Paj8f
cehegWZmXUJK+VylraW8fyq3Jk0TxS8ziMXQTSnYaDcApJr11sb+RC1ZclI/e1APHa8NsjeUvFwH
VxqLJLzL0IiwiQOhUfxdrGh4yVbx2o9VwgGtZ9ohzyttszmLIRrBNlyIq7Bw58YBQ1tWbVA4p/tz
ITQUE8dkx8p4kHz0PYZ4OkTS/r9LtK2cYADZgLc3/bLhA/CSNCn7gesFUz1IyZnN/ERM6FqYcBsg
W9AaCCzd8TaDOKS9EUrR8yoEOhVNr4+DTjJV9zUVDMW483lwcGHKWAdDvfDM+v9h+pLvOmozCspC
TgrmLwR095hPupSQycZsx2lhKCOTpSJAKM3NXxkik4B00nlMMY/qnctfm2XSDp0/vtQGok7rxMj4
b415Rwzmw9R2miLJRguBnIGideDr6C0M2VUPIepmxjr5/J3KZWCsmioast44+qHxE3tvQWH9E7cP
f2D/VDLA22mmZRpEC1q9MzsT8Hp90avnBUCVCCVwfsozFhaZ/UfnhiHArRnZEtzZ5/CM9dxi1NH+
qNJtlcNAwT2wjN/K9/5CpHi3Tph7e4lizmpxrvrQC2v58ThznTU7V6HstdebNKKmkyBM/zztfJcW
OHoPkV1+X8HA4uNNe9ASY+z+t+syipXH6HYLNDsyfybigcZ9mK7kAxqRz2PoV4JQYuz4t7bq5lJS
RkwHk1zIwY3pz9xq6q/5KFtZsc3EL9/b2kH8nAPU2ZSfYzkMwwsRDyWT8GbadWBQLufqmnKFZrJj
BPR4uzjdKeo8j0YuGdP8SBhvEsiaKfCb5YEIlJzWhvHkUXRVnlI7Ks7uJvG3Ay65XDjhbxV1bFOe
C6rNEQjvmEcrpgKoBa0lZwG1Cacy4BZAkXvF3deqsfrPEls6GM1QVCQ4BvuqQ3KL4wg1qUaXaqtn
oqI++CS0nMPbRKnJiMSQtDdGNvzt/PDSB3jGTJRbQ3SuuYOkaeeelu8CnAjrz2LaF6O6WkRtbXyE
aUc1cKFXsbqrWP9aUClvwEBli9OIB7dHv0H5iP83TRaVPAfmFkmqAYV08hxhBafe4k1RbYf3qZKr
11UGqEsYFo/Bg8Z2dntxpRPEbRymp8c+hUh/VM7FM1bIkZ2sLSclaQdXMN/10IPoNtBhYevF94ru
9huPtRZG4MnLs7yAwAJZ5eDJA+/DTzpTf82PEmeMRQGcDUpw2iJZ67Jfv7Pkyx5efRqpuuUG2Obv
X8oaxchUygOJdatlZJhBhoUpLVJcuCBLnvsk71HWkGucYebujBlhSt6h4u2DD/BvyF13tTOtiCtT
JRsTqiGSQqKGmBNBA4BC5pQsM4Z150C/Fqeh400DQOMWv4or6gZc9fmm+9FDPgztfZ1nZXR28wuv
KmWniagtBK52VwazCNO7uV214ZbTzXXTA4VEbCi2zdTZaMN8n1QNmlq9+CtqG9PimhsHZx+ha4sp
En6zUCfrpqZ1Q2rl7mAWzxw+mgPCCnB9mV0So/ToI4Vx0ur5lU+Z8uUvh2Sr9DDXYScK8T1wlqts
5mRffSincUJmINK95frl8J9KMjLqyDT0B45vVKiRAYXwSOk4i/VtMEaDueAK72NQVfN5sPb7NPMX
MXtKJw+zsZrNzD5FCXai7yvxQZosK4B477XKgBRk09heWcG72QPyeyeFya757chOOm6msrGnKxih
rl09JHbK8kN87M3fuY6SxKqzQgmryWHIqcGDr5fE7ERAY6F4VeozT6NpLXkAoy2zeOCMrkrHItDJ
FMn99d3iJVm53Nk+K+g8u+mE3+ICo8cWuu0RsZZDeRlAB1OzCvCiaE34YuTb8bRQBEO8uYtQPqEi
E3Dc2HUM84o80qexi+pvjvTZDSuCEkkIZUFoKUipn8o0gxcn1gSDJtcN4qQyeUxJwqBpM/jx3GJa
68A8N4KH80+wRBZecPgCmaqJdnljoXwWL/571Itq8/vMSBBTSror1ydcirwQxfFk8TcevjPdZ7Rb
gc/tvUkXlXDgew9Cwu4IDn2f0D8Yqkgp1tg3OAt9+3piTY+smui/0XPqvjsxwxOxejkX/xWTxGei
09atZ8GI7mwDBtp/L8HgYaQwz2wa8O7eteXIqEmNM+RuQUY5tjByFGQiFGQkmQsSSo3Djtgv+E6r
KEUBc2jPeLq4MB5wjpAFyFXve7a1WjWLt3RbSd4J7IxJn/B9S1NyM4HyVDkik8ueS/QRcx/QtJGh
WrbEFAlfAE7wQjkXOKNY4srY7DlEp1sEAf5g4gc06WMVRDwzgWcVHgZk5VBt7QvCUv4T8akBtHmg
Qoh4LgN0VZBRGMPvgNEBXbwp3jmbGym5IMCYUOwZZC0BMPZYG/06dnbOoxtzrPMxmMln0LML2lC0
R0eK87URX+zY8iBMQfxqsmxthZHz6ZwVZChob8zXtDVhQAAH5xAjIkNEW7m8ifuYPUpg42koqCeg
hPRP+4iTb7Cp7a/vWR6e++YBfd2ShXZIHBM9PxLvdPgbrw2nzkdKfVWxgSU8dniCXzKaCILIaULx
PprCllPOxb9mac4BWEhmknvjvVqZhPAsUbRB2KnvYUg0CroTsgVtM+A06ymF8JS9fNnZtZ+bXcOa
+3rMZMMxnni8pPM+R0oF8sVmfmZmYVaZug1dmlTonnJSD5ENSMBGVL2hjnRtCDT7GrSrWHI539Tr
BuT75IVhHcIyjaDqRTwEXaId+Ec6WaNY70gMf/GI2RmVuEHAX5V4hkG4XQI2nNlpXa3q/qANIoM8
+0absZ1UbwHvpGGfq2BWVt/el33IZz7mYzA2VtO4FzUKkGr+TqHbZme4ak9e9BZp97KjnP3ses5B
pggoDQNOqdmbxUEfes8DDvJd42mr3675qdYMQXuk2AZLv1EvimxwULXYCiAR60tg8rjb+K76wJ95
7rwB/J3n7cd9pYJh/MovGvsZAesOrEWf/VtwRYzLrOv7XOOGhdegcDBQzzjTXZcFc849rVGVKujl
zL4KNVbp3NKdd4IVxhlhMYXTn4V6+ThJqmXWrgy/IWDsZeceqCcIrLouuS87gkclr/XE6wqGn+/E
+5xsQRHtSMfLn8h+K9VGgb/zAKn0vBl0x/kAYSmwC2VL7eblI+nyjQArDg9P76O0ieQvgenOlFfB
4wjB1VIR9SGoo0SY8h0Vd1IgwqKHTgAGt1atZNWnZEMHD6o+Nxp3RQpegQ7T4vxLVjr4OXoXD2K6
vZVEmhBWU3yU32Bgpcq30q6+m9EzywprPvTbM00oRxE0pTag9fpFN60+xBqWM/Dmr2vIxNuoPk+r
T8CK2sx+oiPn6FeYOqyMW7C/UdQzfMCJsOTB5x0CpEvLVTpeZuT6bA8DFy7LNn/FWOCDUdyd39Uf
AfNTVQDbGcQmE84X/auiabro9HNL/Qlwq1FrfNrXA2qymvKcgTATJrvkv6HrucRwyawvmKKEpf7T
QhBm7Lfxmk1Ltn2IEl4Sp00hRBM55s7UCSu47xhu+r0wkhUHIeYzOOE8gz6r0Wu9fUFsV8JZBXI+
k9RwCplff8gq96KGrOAUX7y8rLJhK2n2CWujxI0xUOkEnpOeTPbtjli8n6z6k1Lfz8unwHksHKG2
R3593nt7yYUSs4Sd/SlE71SSJa7zK1DJZRZ+Fks4u554ETbvIX5BgPorZPAShfQ8/zaeN1l0rCGH
T9EBM6I2ljVUb2b9bC7qoB12R0c3cKihOFHUNn8CYxiAEzeGEtKv4CcFZd/6rcdUjJAEFHYofrus
ZdPc4hzUaj6A6QHBK4Z5bUfXGidkL7VvwgId6SCPY1SQ+YVWzyM2UP+eXFT7mwcYxbt6xa2S74St
4gTMvI3FSyj7yMoFFulLutuGBF2WudprUjuua7xHxQBrFoHLhxhVsJ19ugvbaf3iLGhobSo0xxrx
4MCQK9cahc+9JMwCSNfcjJRIQ4AQms6cpor0tB5H+oIpsxoEecV0DIUeRZN0aBVgGJbsakZAdnNw
PF6i5DB5KJHcC95t/iQozURCBnOlYuZ5hm6R+pczFNTouRrMvXp1EOYOlhCOMD0inlK3SI36LtcA
US723Vq2RL1T0I132EyXZOn1BK7+XwUC1EpkTV/V9xQXQitIl0XtjlbOETAoybDGMh1UPyFBW0wF
yPN5JxGaJ5aNwuMX6ERmdQAZyz91LMnJ/4CWcfrBmcS9fIfCAc7xbdDvBiWVsK+LTnLOYCemtyFH
iwfzmK/1JHJmcVOUv9fX6UJrq1CdDGB6i6vNeQnp4W41IUNplzqk6dC90FffPyq0DlQTTJoJPGx7
cW5re1TxAj37U6kObdGfQc6/pVmMhxm1hqukp9h30Emlw92dHL5rstH6kLQu7pjL063L0Dyicb2x
dMAPhTbTSsmTzUnOn1Ziw+MR3XrK5lUwWwxX8HpfD+sB7QddBFWtbuzSY3XknqDNRTiOzOgxvovY
ChOYxNpGJR5PAXPZM5RPcm8XCI7eWzzCLHM74+8Q75VFs72bs4X/hHeSNYaUJSPhrC9EAwVnWQDO
gsHyc5KvfaYLAUk0aVJTA6UlPGiDO5QPQx7RAVQ2y9OE6235yqzuLiqHA9LGzVrbljbcjJhz8ZZR
g/vqm4Xr6U9dQs/5cG066O+TmAAybywpJTzxZuYEhQQWcKlyOYG4mfu60AXa1CeLTszD1nxJc0mH
oOuAn4dPAgyiNaR1tfKfYih/mBQX6e+2OMW+2hveG3oTBI/5ZcnoPGh5DlKrPOogjXzg1X+Xo9TI
umIshYrbsKTtuKGtif4P2bUk44FE99+c1bZqvV4TcAlG5LlL0iyOwZ5vD6cQNkt2Zxy/7o4LA3CL
mf284YWR+JQ0gBtmgxXQf228EJr9j143muNYTaY2QpAD+1bw35twPMTOJ3btQq9suXpTINcEB0Pa
rs/aA6zV7+ZQOCTyPDo/pqsPLpolgckTXLXAqP5MMPwENXLWR76mg5kp7ZvbA/ox6eUM9/FbiwNd
hWfIteebJWldLpWP/zUGKevE1lT88FE9+EaIXfV6kjwNz9ItSjFfbicO1AfXyz61hKCv74wQLlbe
nS/7XbykbL5Z/4DX0Zm9qplqh4zBVQNUjK+uPwMpaWSd+32bWjznwlYP5x9xFDpdAPu8/NPRuuh6
Z2SoxOPMsUQuRIyjuRUwQDBPoWtIw/6464QlH136V5GV2JVtQK76kIVbzRQT7LvjJ7gKaI7MT7gE
Q+IZzYN/vfUTQl9MlK3I8bQlT0IFzDArcE26aYHzB2Zj5r+u7086utWhhpolXWjFWHkYM1KsROjO
Zie+cRWA5Z3bFhzd6hIvvxePOrHgRQQuEKtqKDY2qpj8C3UlP8NXBsxDLdb2rh4VYDYiaZ+OFKL+
Nn1akn4LHqJ2uws5bZfZdXEjrxY4R8KNaIh7ddkZX5jNOGm7mnDtnR6hYrLpjcHz9UbW+0nKor4M
Cc56sNXXqAaCC9CzDhX7kcTcn76lqzl4nUiMQFhE7lUwpdE+HXhppxsePGlWaMmBa9pJdHWuj58H
nrwvTFYgcmmLAFR1vuAC960z0lfY5vJQbUnXAfE4IL+uupEihU9+vnaADGN3vVWelT1AuOeww0IU
GkVRGGmX4/NvHjCSZ0+nRhZrK1p4DTRsr64MvbKgj2vlLhznBROlRT8A25oVHWhIimhse2DHb55A
wLikpjmnKSxdjyEjoiGl3Rg01iSUWNMDjA34zM7xh31pKa/e9yjIH6MiLDcDocle7ry73S30YXce
qViiozxe770uNt5p2yYJIUBwWWD1gVnhuUzF8wNZ8TSKVbiUiz2YNgnt43uqARDpkf4ldlwk1/kJ
dBfIDbv6O0f7ZmRUjfsiW2U7PVfWTVCUILvjwieG1MlbxpG9shodEE2bd4qClUViAc+dn8qdlxPm
Ph8DSA9oDLP3oGUZzPenLjuiIiGQj7legsGVhDMBZQWHGoTN9Uj9wavNudyB+y/XIYNM2ILZqLQo
4Ko2+ZJqFuQWcEOQTzl/Eh4Hhzn0Nq6VlW9BcXqDqcVDHFZtflVx4alhZyDopt72rlBSdXmqA+SR
Sw0nK6uD74TKyJ0I2oI8+ht4sQ1ACdTIH2M65TZR21fR+TDMto+/KRXBawIjnsOJXAnRVjrRxW0K
uzP2ZW8dgEXWhF94fLJ2bMZRQGmOXg8o3YS1dz0JQrHBFbsZkhLHLOAQLFxuK/67KnRQ7dDxyHpw
XJI60uuWhr/qEnLMBnNkefLVxEXBjJwMekuopq56oo9zpx5iZqC4S8fveRfLZgI54UkKcZXuixNl
5OANEs7X4/gmCTN6x0m6V5BZohZBgeGiVzih+VUEmHGeUBBcQjpJksllUltJVt/saWiHSB7eKZId
IC+WnLRGrLyLMZszMYZzk+/aPBdUOUo8zLchYsfnYqQ+cG2j/zwdj0CjGiv+xMVM0vKcwBS1uSVB
9ALTV/Agu6aFVuTxKG/2Ez9Tn4RfwC/maBcAhNnxC4xZ1uwJPUH0JrSbxp5CoA72mhk4P+gotd9P
KcGFm44h2gb4od1iX6Lu5+1eQMDGkWnqBXa3bLCr9CwKo+L6DAxUBwfBIr4i/nOFYB5poqdVahuh
eJ6S48MZlGswvGAQvtsV9dnfBOEqWFOdiAdLZ8CPnBsTF42NP4VkQBj8+9MwhWu5ckPpGFQXDcnd
X8Hfw4cLTobUUoZXc7dpzzRhC3ik//HJeNlCgASBvDrGXGhB0rkYHVFdaQ+ika/Gycl9Owe2Hy++
CYAwl0OXJJiS5ZDoaLDRe7U4ARTx6YYwoKcDNsjvgO/oH3bab1fH1K/nxtWBYvo8KNUFOTTeN1kF
8m4n+EsPnnRGu1eM9ZKWImMwSXOHEs92R1pQyVYuoJrduvGzUpN5/yCGN1nlw1p7uPt4/JRc82ef
5yMSimoYFKeBDVfg6oM/WS0pSzeyoV17mdUGoqlMWm8tmaGH4hDX37BjZUQb4tH8JLaliocmTghZ
wxelIXs2wD3BdPV8QGLnJryjxh4TNk9WaxHKbcHA8bGhC4Dds8nfDbZfIvK1dwmNrXvoq0ovBxYv
pLBmN8m0OUukzprBqOvZb5paQzgNfg2wjNA0P8KwOvRu3a6d/r3l7nep+8dCR8JTwBevzHl2N3jI
gx4XLgGIb85J48N98mNNbOE1HFlCMoIwIx1e/eIe3N3zE2O3YNDRfudFAePj7DbgCrN108+UcBRJ
UrJpQak/pLpbKHh46YdxPyGWNoXJiwlfyGgGvQraK/MCUxcym7zsZkErXNnTLDpBMJrb7TpXOkdj
0KKAdh64IPJZ8CKDYbAGXF2701dTDsfMELXDXg0CFJ/6CEceQQyq0phxDZ0ttm5vdmNMHtmsCgeo
Wkq+Ikqr5jOSy2AJMecmYBm+K2byZr8kvQV5NH2cGgZfZCeHp3C7sghJXT9AG1iyKOfqTvRbrdBt
03JvDNvtgC45KhyAHQ78pRJ0ka/GCJx8CCnxOztJYtvRLeOfCQokPJeJuxWrFK08TKgXJ6XpENq9
S2yOGBAz+iUXws7a0TbIyZLM+v7Aks/aeZq6TLobfwgNtamltLbzagTa9LV1w7Lo3mp84paCqdx9
fSXZ8Zhq3jSXOuxTKKIYAehzrO/qwQ2IBzj72/PRpciwpTLHHFI/ABOud/BwSU56etn8z/0MU9po
Q1HqoNTGJF+icK/gqOR+6tiwy4wGGUeFFr8R+Y5KnEW3oJQ07awn4rO3P6OWiSBWzba4wE5TKaaV
vLh6yCCALN7W0FG0+MHh6FHog1nbBHfx2WRrmm9kyBMH0SnkXoeBUYG3A7cu4c8BYwfedXWxCrBA
/+804vCN9MUFv1JLbkGJvdhtKJwUFQ57CdnS44sgbsPRXGZxhLHyraGUHh8JiAF/U05WfW9jzJqf
6QiBPMoNjx/5WYq2au0Us2ZzY6Mzeimvo1LrvIIsjKluudhdaqunvDA++xBW6yJxbqDUUKZBH2EG
/9jzAD+AB/Zo4GlFVW55QBLNfr4DRmrDixRWPnlAHQxkl5dWlu3rECaExG1UFSzRa9hf2bKd6DAp
xJ1bhGl64WWYa2E6M+pZm8q01UFeoVjII5Js+kkxN5ZpO+xU4l3KSuHvUEliOwMXpoBxyp+PO7sm
epzr2CFzrIIuy+LK4v5KwE56BHp5pDsLOkA8MuHyDMlDLaOOMEWoHI8F/YG9npJfiRPFK4BlRuGM
fRwCc01CVQ2/GFRO6+h/9snIhpOzPpGcU1My4YkmcxFw7BOIKhW1mVRmeKR5R41SwGCXGNW6Z/FT
gIUPVvqSuaf76R3USrsyo5WzLixxfe3VKUxZqcXXd9nhA2qJgLNPyMfWwtcjYgJHPv7TdZkkiNzo
prWw7k3qQmpyvDy+aQaKfsAaj9uwGoJPSwDXznFGzQYksJsaDdTsCU0zjwmJ4UYGNNVnEpxaZWx/
hfF7wiq+1yMyaM4oQDaA2tKU15pOc+HEnqQsG0yqOvg3xn88FzPVTdiCTH1BX5Zpjo7jC9jHOF7o
BmQ7F15TVBvjpqQPlCMF+4NL6RLEGeZEOn373wl/M8kCRgzaXWDbkKmSN2wm22nfxs0hpX7KlASv
j2UviivRt5CAmdKpXdLkTjgSrQuuHsjokO+vCghvfaUwip4hKBIIA4iyKDkJZiq6uRSFgVEblgEb
6T44iHuufZPV6Ump9iexT7AqMGrwrvLkTfqlfirNxwdLVt6Sx0oPqm59eiUPSni9jTJG7uTrTh2w
i3hxdgROfT6pPh5/+Btt5VpP9kz5cX0T5hZqcE3WSlvZ+5/Jl0XKPSlFZr0tbDR/FwrITH+Zfa+e
HtnBJvDckklDHRgAlZUMeOF2+hk5ygVUmIBTWK+Nsl/dIfDMczGmiMCD8QHAaWRbw43fgDuTf/Pt
Y3K6DGO9cpAckcwDiPM2+4EG6Z6l3oqE7pW2EWsDvMpzSTO2kuc4xY8B/+psdMRQk7qWuPhC/9Hi
/YRDH7jPbfoNUUqbdxp9oxGpt8OM9dhTh0qfcttPHTWVZrZnG+ubVn6YQqCbwGm9yD7qaPA8nE4w
/WlxuewYsIe7+6+n/VkhgI+UZYPTek2PmO6ISCzWuxE4XnAUbH4c0m9UNWVNO0/BaxkvUcxXrd5F
7MI5pGGfzzTjcpMGFd9xUhRzBGaL6OSLDlMt4bevlSx0sVal7O51HIJUM1GbuSC0NVE+jfgkYtTl
oZ5AVE2EEEm0ygy/cRDYNoVGwnboWxK/4q03irm/26OAMtslx/kjUYuyKGWxYHt+RDMIWMTux9SQ
dOiLXB+AmVyr911F88aYI0rZg9lbKf7j5gJrDcevlMAS+QxGj5YEGJnMk7bX2VU+tJ3rzIgYntO4
bgkqAbhHeFWZP71DGYxv5PtBNbf+XIZIt6mu+W8rLVExX2jyWprR6nDgdSWqcKwnuvCjdeJJx3AO
AyZ8DDFfxkTiKnImIWj8bMi6Kp90JWLXi8fOw5m+8A7a/ufvw0DQupbK1VxK5Xhz8mCek7Uq3gYa
G8AwmafWBrK0vOrsSfM+pZ4yuAzR5Vosuk9LRP8snm4FrYM/1w7ohw0P24PNxaxc2lD9KlJWmbf6
C8g3FSqOzx6Zng5TbNbmbAEwvmvxdz0o6BU1G+7UhQ4T/iMsY773YUKyXgiawGOExuip2fNuU/yM
b3FXmO4v/z+xqwgC/fcMOcTAjaZTy36P9z6E5Dk8t0NK+hjCd7bhmdAgPTyGXBZfReUdq7/hv8Hz
gwepavXzKv5xyTrvNZ4BpXMY4tWtX3Vkg7nv1ix6yj7C/RwHP/6r6dLbph3Fed7aiGJXtJzM4vUe
8aLUcVPg/EJPYIPjLSDIApCn28d0ynLdkfLslnFO9/uwEj4sDx8XwWm5YPCogHAnjMd+SFSI4Oi2
mBX5GVLy51eL5vt8oiJFm1buGSIK8vemnpSJlbaZOjDZ7CVDUfDNyYsQwFy2JqfKGN963S7ml1Da
UcwcqEJc4HYXRzQ8lUbsumBTB2KwpC3gTcx2+TN//GBbIjfrSk9RZ07aMUKkPEodbVoQfyfY8+E2
A3Iv9BkzDS+y5JLsZgKrEUVJZcAYClZoCupQ4beoyNl4DDD2EHj9mNenURd02X/CUUavsztxVN2d
SJ3qjI3pibfOZAHi+XDOri/DalZqyEiQHYDNSaorU/jaB79wDepgY7x+CVIHTcMauTOc9LBlTz//
2fkQtg3bBIAoWVP7GKR7ZgQ/QAodx010HT2XzxJkmAqqC2bdneVhJmlT/NXsfO2OeUhVAR+SsWlE
j/JoTMDzbodzgRhDuXAtDeKu9FZb/O/o5YJp19216KuQ77wgHSu90t2UnmH1y7Mt0wRTjbjIb7Td
2cQh3dsMeXrbkW30h5CXMRU8BSYH/KArGmPNwFhWBnd40tiJIzJf7EbB+ZVZzR+FHCZDiIhv79p4
QfqgGYO0acl3afyQ7ikgMc6NNGvvF7xLZGPp1sjj5kJrAVYQltwZEsf1e+1p2NHYES65+21wHTVf
jkqNWQGEmEbcQrKvys7r2ozMPKYTPDXpqvSK6fAmjchfDmIgTDWhBx0RCK9E7O/Y+0sp4cx+oBqQ
cqhTOaeuEpdJn0OnUkD+qBtickA0bjv+5/RUEYuT1fGp+Ez1pUHb3E7UQeZVMT8uUrOrP16hO0Vd
zn7xNtCdgSxS8hI8/USxYfv2c4FTZQpEK/QRC4tsmwZJBlys505r4qHCj+b8BIkFXb/QgGowOT5k
gH6VpN8XiVCl9gTEkIIEsRtLDgjnUXqDD3uJvh2HlHtf/lB8vT8iFYOg+m7RjvuL71s6Nniq9NTd
/6Z4ho4I4X7xuDQ4v/GlxYIpypiIDNbEEv/i+tYN0AeNCqt8/c9KtYDbwOw4l3/Xb/HTgrvPdaXC
9N97swXFyILtyt4QuMARfuA2f5od6XpeP2rPN1TYmvipb47vWglAVs4SkbOmjlHDrJlQ3Aizs9AP
C3tnT4bzHwRYYe/VCebZ/tpEK5jA853hMvbQ2IDZSHoq6YyEB+gxBFHAQYlt1IhDgktYUkx/R12R
aGlom0Tw11bc8LSODaDS9C0F83JkNzceAsbrSBxTbw4li27L2Xq0dNEt+T88UNbqrpXofUYaLcRN
I9lfE5rknT4x2xVFpPCaPg9JDSlV58LwjBzG+T4jRhlyRwBHr7SvzOunRg0djhnd3c/rvFzjwzRz
tkTZ5AtpiMxN0AgYxnngIYqJJb5vZKmpsz7RzD1x8gCcS6qytIxV91UaWFIyLcL9EcSkxYRlg5wL
+p5xuBYJFVczFM/RFQknBhRe8Sxq34rGvlyUySYnQfi7KRagk5sTDWRC+ZucZJB/5z0d5zQjKyJR
3okG9Ihxcfm6vSoRzdZDPZLnVL6A/9odxnf9nzpvgy31AA9sxqXLAEZ9L/cvWKHZdt3G3MGkX3Ou
MInuHUQH5fP1rQAFOmt60/dBwsMtqYXrBMgygmhr9dsptM0Kz1CtGOeUGCl1m3XZEsSJVm+ee2FR
9oti+iMQrmSjeizAYQdgqb4bRd61jI4AmNItc0xkLgrbqQe9UUIqfj8jQkhAowWTL3o5waNcGEKw
twnVJyvUrN6LdAHGgEer2DUx6Fcezqh6SDgeUgQwPd0m4gDMhe1mbdIA0GkUEHdJ5V5/vVpj0iw4
UhbtCFn4pSyfUOB9L1Q95W/6tA2QUjGv+Ay8ruUkqYweuowBZQtKiTIeL1DuWW6eXyoyR9LsE5tm
dZ/iPEhInfAh4zOFdtv1U3niZwqitEOK+Jku5Ll4SnOHq/9Z22RHcgnJQp2KlwRdP1L/7rPWRkP/
uyl2Qhix00PLG0yjMeWP0jQDX1jTWh7MXGGHyE7e7PfM8OSTt0pNYicIU6Lp+SUvx4+oEKJzMbmA
DnpcflMJVnlcRXKUHRLwKEY+gaD5py3zpsH/8qVnW/8AVrFm+xLRYDvKn5JwdKUCclnI+ACHEJgY
tifi9cjQu2dGx7d4TagnxDA3slLjwgwqs9gGKPBn+xwsNwvlQWxGOKcCE13Jt096MwMBvHBeXyZr
fQTpDO9hM9eBbafoBaYWQPpOL7pEs8i4M4aUXVPCGR9dOgLmvSLoA1NOb1PCjYz+dyR8JieDY3ye
LbmUzCoMeMgS2Whbg+y6nC4nk5XQ6VfxmAqknlyR7J3VTSeLbJdkd5KYtqNbWdCEgx4J8rX8dy/O
UcBPQTVUKfCQpVgNh3p4GK+c5kU5jeTnPo9mvo4NvFx8a7m+/kTRsgeyRROnQzKTzTUl7RJJ56cf
2vKb3Ds5R3tNxL712FE3CZ4PoR/BA8nktLbsJRqaUrcEelG1MJIFK/++BD9xB5/vjbCBGI/HlkRk
yZi3crLYJRmcb8RxyfVmOO+sl71dAKYB+9IjXM6O3CiZnb75oLi3hHfSGgN33+2v1ICXOpD9R+cj
Qm2mhHurLOuMSXRxvoO4/tRN3o0HxWXMGunO5vtrzbCkDikSOK5sW6sEFhgEuU5imUp+nAjxuuKW
Xriqc0tqMxvd7ubIZAmJ17ZYD+/BODEuD9Q/oNIEqKWM6Oe+/DJtUvZLQ9zX9EYI/8TFvZyxheQy
r4JUvZL4DofT8u6wacsh8eZUjAQfxVHr05RglG4oXR1J+5gZrlM1r1WUX7/aJJ+weKqeQ0D1ZGMB
1qdW/oDnddZLCA3XAo1ket40AddAKog5+SbPMd1hcICaFTUko/+I/Dbn3CirmAD6QpcwXR/hC58f
EUNt1wzNBa7NxTEI28CWt0/936vNc5A41imcqq+K9tt5eVGy5ivZwYrzvP9dMUo9ntplGeFPFAF7
zN34sZM1Vbt/p22HkqXc4xmGF50gW3Q11lFDmEOvSmh9lWoGTh4gSEToM0yxGQJQVeZLptlUN4SQ
YU03ZvM5gASf5vYFLPi1GolHEjfU6aa3B9+vqtCP/0lvvGNb9hpiAnNPmvfyJYTRXONJzMUJzTAk
ny+R+S10YfPmhpA37LdniuTX/eCIfIkPlwsiu4taCduSpSSz71SDvBqPjKU5+CRKTymjrzSe5WMN
m90jTdMPUkBzBDfeypOEf0iSM4x0aNzYW20DfiUb/oKc4a458yxIOKWCP+2wB/60pKkoP4JgHcrP
CTrdKRXBslM4y/ItNoBUzTPK1mltqu+AOauQo+Mpq0PE7wBZzYmO1bhPxJClw/sYJHHtd9yrFHvi
e2gPWj/C9pv4rNVl/+8oWcrqaZJwAQ17C7VdX/cyn4L+qcqJqMNaW0+zu7uI0+PLmGKlDc1qb/3P
jTOEzPgkFsoUOmjUVdSVq5doGgRdbRxv9iQ8dcAlU5CxpCOwt5yoPQgYTWYcu6EPRL1sLBw+xj8S
cfQsL+iLX7KzxJJOnwLEffmj4VxJc1SqE9O68EYW4nfj3Yt9/vCsianGxx1SwWR2E5p+16tWHhZ5
zViDcI9G84fNqhFkq07tl2zErMetAhwbMexPuQ53+N9ry6Z5ZW5SX0fotyfgMeDhvrkEYEv/iI8+
QB0tnKFpbY0yFQhPRqomPmbF8FfpewT02bAphGMuNi8wZmplkeAQ5ew558q0IRXy9hoQjRQtir3W
9Tt3F+rTflSLU8DzKNb5cg4/Ik3xQW3UoQqqUWcbzuWmaRq2vKXCnAjKwVSidgKT5qQCBiVxjUFU
7zq/hu2MoP4icKW0BjV0f2tryWcrJjZ1GViqGfSYHcSjZAa4mD8ti1T9BYLCiOaY3qIhPup12xq5
t9m9IVvtb6B3DrqD+cFZjLbI4HcxJcVuLR7wGTumDyBg6HNAVtXBsMHVP/jGD3Ne3Mp/SAWMCwZx
2KA5B404mH8HBtC12By1pkz1oga06uFdYsy5X7evYzuTmiKXOu7DEKwjz6NAZXUVe9K1Kh6koQfZ
nw0ufnSeJEJKD0daXmntfPhHzSNQVidNipe/G+eu8/zJZhtLyX3ODsPVdVSMR2mmCWXn4kInb4LE
wTW3kNj8EXMIR1DOa1QPNpdtyf7s25x7ovCZmg6e2folbBe5H2BonRqQbdKSR0/oqZKDsZBWcdJT
KrmB2lxWh4FlhbZF6J4iAGHDR96rQmrTwL7IEMQdsJyzsQJW/BiHNaLEgZbY5C87XCK3K3tWbMMM
QUwoJEZ3gqdbc6JThfQsfwNhezAB5VWlCLj5G5v0tpoWo0hDSBP/sszO0iFqYl1uF+Ua2Oi/OLAG
uP6+ZTE9y13eeLrlmwMldhsMTtOoUeMebkYvDB5/evqdm8q1CEV4zLoT5Iy46iFyH3IS/JIXumXM
Xd7dL6qd2Jdw/g/a8FcWwqm6ux6GPUoA3YVAPeioyxV54pea/ZAaJccz5rArf404xcM31JLeZlwN
32VRr7xWc6tg9W0znFgos+YLLN6059h5CJzcumcrXTquoCdgFccxTXncWLyeG+8ocdjZGlzYmRN5
AWd4ESc6/HKAxTP0nmq/ay/7/IEbYjD0sXAgcVUYZHq5kpvv4yvDo3shqd4OSs8rDEpt5yE/2oma
3u+e0LBdyHuWTiN7iJXVqOSQltopakgUL4pEJDn554GJKr7EYg2PqeMPtMEkb9oBL0VxisQlml3A
QA8dNy+v/nB0hW/ze/yfwphEfb8moBBguXR6XemE+YbZ8oI2KLWLm6WhPWzWmIDmfMqWFuiv/DXj
DMoxOZnKJPxU0tJwb2sUErx3qozQ/NkjN90ddxmyhrlRMtsrFYCcSpVRVW645YdfBcg6u3DBbpLg
EHe0gBvth0sKuL5kwNSPD55vO449arBoFUCSajSgohddVtncp4oBA80BccMN+7yVMsLjNqpwbMEP
IPT7F72/a1SmMz88vHQsSMoNrZ7q70vMWUTBaSRJughtzgNDLfcr3QtNysTtRw51K/xqzqFtadM3
QyxQiz+RfWPVjSL2936GkJjKw0CFrpuVJUnCRGv6myZE/JsaucTty2S170tFk6MrGlve10kD9OWd
panNg1C2qm4H53GuReW1ToEhxlNhNhar5ZbcvXOyjsd651Rz2Xf3e6SVojzQG1U3nhbhXYrPEV46
xcAnARMLi5DWlpbIiBxgtvS2kR9JjXt7/46lKEbbXC1M8BzgRZNp19nRTXDYwvBO1E5WIsDra3XV
02pi41LOkvenWUKsF+3rphCMn7uwQqVbt+p9wHSiglsVB3r5qMhDwqqc1Jfs4n74V7kmfkGDGxFA
436VetE+cEBRoEZVXOWmnDkF5ggYeJGdbgKwSgxSrK+DlI/pUOes8XvUuZNxOK7B6Vchpio1uGMw
TTls5liXy3CdPKmO44zFmBKfV/IXBLSwswFOjGDk0fk/8hE5CQlbYErvNXdvpa899kLrHgYknYRv
CHKS0HFDxTRM4nsJwqj4nNpuPbFr2luBjNd6xyaaiOnPYBVf7hkeAGEHdFuM3640FZpujGLCY81b
QKAFzgAEl2p89VAPLrJ3moiaLn6N8qkJKOeoWLjF/oNSmJOoA5ctXc1ajcrYecSRSgtM7auKOki3
9d1qiyIJ6sEl7Xqk4JuV1bwYBIt7S7aQEeSo+aYBPk9KM2kOpweAe53snwFHZ+1M+L/ai2yWy1l3
hojoOheJUuJob7gsz6n7vSAHcgkyFKoFYm158QxZj2/naO720qu3PakojqHR1fvZeEMCdVt3ebDK
7pZIAhsiWS48Km0qQE2+9kYj/oz21gDCqsjH1k2gPUkZfIPvqCejMxeWs/f2a07Etx1vm8F2YIUd
zNNKwS4bd3lPa/sEwNHd3HRzBx0gGPl+17H4lZ/88McQhrV26E5/DGcIHj2SUILaeIPwSneXrcO5
amFHapSHlDmFvngtJki031eZgdK48IBYHgncF2sQHvSUwd1C85Ep0TW8y6fWSSW4PqzoLE8mRBvc
Re4AhFa6Vbk4yaJ0tB1sGg7q+gfPyOWieNC8Let0ZVd6wR7/bTJW7KySMzgkMaQbUVsM79yOR3Ye
dSmCLJD7qf2vtf4EZ2nRltvNM5V+3zyXswJXuogB1cMIk2IVQdHgztbRPVPQ59mqFO2B2seh3CWh
2FJ3xoZsGobdpbZOaVnurSgIAdzLMOCLskVFJh0WeyHqe44DhLs30ucnE5/7g6FQ7jvxXwdRySXB
yH5wkZ5pyMW4PRBrL0FKV2AuDCK8Vv0PN2OVWwArzNi6+M9WMs7/ScdHaWNwOAc26jGmIABszgip
wJWmf8g+mCHE0mCszTPhIvodj4i51vvSJ1P0D/fyq8BvLQF2174vRoAB80LtB7LRXxIXht7H3zOh
ufaH1FDi6/D0lCn6lFGZ02xd/fYDSVsbh7kpAz206K34u5fnWzm8cYnIAIegCN/67LTXZMcBLvyF
BwnO+XmcfljeJ9i+84Z4UN5h72JB2GgyxCtl8TuzyZmjVQScta4BR+g+2tIINVhQKp3glIsFlt8W
e7FMIBL1Ns9QpD9y+YcilsVR1+SWyjImsvM0I9SrA5NpFI+NRZ7+dDVkwHMlNdy7PvnNZKIt5grR
hJh637TPH4LfZgWHZrZRU6T/8tGyWfPinSNR/UVKWxcG4haaRIVHlcZmMrX1n2xmEBfWYZ5cNjp1
tqHA5c3aupHHK0GN/Eq+eIvBttPd975fnRBcpRc7dilfIYgx+pIhZdx9C/VXadAhWFBm2NA1ALdH
+kTd0Pm27vXrYgI+sf2OSTE4/vNHlNkv0Ept3zIIWkMvsPdAsLOsuWiSJMccMyKO01aNhWsigkYP
6mnIoqPa51Mrc81r8BQEWP2cpygNCZXx6cXnXnDNfnE1NknOCxFKdAtFi5WFqItujsc5GIipmhht
LTkE0L2DFqcV7zqEDZ78/GGAaepNAF+uHUs7pWvXtcsrsNM/RdfIkW/Uac4AG5cQMw4Y3/UK6HwZ
TI2JhViEovOsSbvC+1d/68+rRJ31Lb3DpQtp0V+RGUiDpu/y2sZ8Uv6MNGEP1k0bhdu/pI6XCrul
90qZh5AngaloGkyVPe0dCW5pk93VnDUTNuCmbUkLm4GqaogHT7d8aaKrcomP/yYhzfdQAqYM9tZ9
LKLOrl9ZvMaACgjCnL0wp3sB2mOrMldQXsliH8F52McdRHFRU89thvDY2IHpyWgWFaff9wVyIz/X
QAIqfJNKSlfd+aCz60a3LtNv+FLrQ6xbxaKN4HxGQRmzkUR2Bf11h2fpbAohlBzdwAjeE48POeIJ
/4ObCFSX1yiK0EUq9ZZd3VwINUqEqVl7wvEymihGiSKmrPAAYAEc731jMQlT2UOzlVTd7GuVf2dO
3Sh7tGDZZunqh+bwqbtQ35p9WVGyQDJ7Q1Ovnxesdeq6blJA31bldsLGydcf6lr8mn8S/1LiKfKU
ww068oAc8ZCnq5+JBOnyefo5eMLZYvqPQVekdwPy2bdoS3oKHJheHf/HsOHQVvHkWoAesiqlseXN
Hm/+Y4mmnBMX7zh71taSNiPsEk6mj7iEdhAGaJLJ+5WuA8zv/jyNhc2jAmFt9urLoMkmt1akJXj5
gdeK8n89vGUwWppb5OJeR2IHsXvr1XbXBOBbQycICs+856H2wqsAqYBCWoR+2Hyf+WqBf3XrvU3U
JY0sd674GLstg0QGhtBMxkiXEQtP8aasZHW26bMCsAqIiDZIzTjov3RwWKJhXuA+ueKH3HpETpHA
+AATx8QeGM2w4WwWYM5tad34As5AAQ+Ft3Hvy3YcZ+ozF3KeonPcOvqXymZ3m9VfW79Jq4GyiTyq
uERfW8mhESL1O9Zev/R24J51Cim+GfjJx9B7sS96jDGqDVkjEgz14iKueD6FLJj1+xrJ8vkMmdUI
qmPz5Ayd9eKYwKPf4UPk80M+E1OgloRCTZVzPtxDOiCakrPxTyB14zbhswwVQMX1RAWkCJg+CU+i
2QsZxxvb9ZNmpctQpsaD9tmbmgT0J70ah+4VVxmzoIHN0XSjrwgey5POMnvKB1ho8Zp9kbMSevby
7gtr6XEts8he7xRsXZgvikhdov8QH7aVJQX0ltCHr4gxxrCYRcBkjYLHyqmlXIzfvXdmLvJXif16
anNfsh670O5M7ZWFxDW1SloeZic+ICkh9hioajeIVPo9fgrnLcYZXcwUycAOEI40Lgtm8nypm8/A
OkJaSK5aznA+vvccOaHdiKCc1v+nC1Mris4rMC0F9dky4YnRhRnvCnPE0qdOXKUQ95mJYChWyQu4
yLubfVb3tVlNFRtsjxQG6qO3zoKK93v5bpznla/gTaDYZzSecWe8x7cchZdnWNZ+olY+Aoq/ILA1
eOVxM7BDibivUyYZK8dnLozbpOuxTVrkLMG5QIemLjQlWp8hjMGUY/oYWEC0cRusMpA86aQ8WQ/g
rWAxlbdPosb7xv1GyZkrp7NJpEmfp3vOG1kMthefZ+oX8Xhk7NpLvRs2AX1/OaF7cyb9BAg/Prf7
XP156BLrT8R+ExD+iFejkAQRImwRB+cx+STF23TxICCzTbVsZLbPsGXHL5iKyxRA6Lk7Q/Fpn+4p
0uGuSbZbJ7Z2YvbOS3XWHhEeNiMtvNYrY3trobdfnoNh3pYxQtPlCuRpjVr+j12r7URYOqA6m3X/
8wAf7S8A+yjjiyj6sDin78Xt4GZNAWo1DzPUHJyEvlZV8QQXQfCtevruvJoA8glevU7sdGzE5ysN
l0ByvQ7GkgAPbEw+gzTtPu0kmeJ2BBxlEmzKt3mwRdUGYMAszSifh7+2nORatXMsv9YwylXKjcy5
rTspQr/VfrQwGEskaluNiQA8AjYM2KlM06ffHmSmItcJSpPQwCHAPDTIqYTkKUBQSQe5xwX7KY1j
7ZKZoeq3uUcAqwEGF8hxJaX64rigA5ulrPbMvGUFtVpXamI94kKgplfPzmi75Yf5yBk8xk4BnXBl
B++D19YF9CxZx6TRLOTRK0hgQ3kNKl6BpAo2fUKsPfdMud2i18gC+HNcnqhUOJ2cHVhqx/PHOXRf
Rwb8/X9lqgiw0k5zP5INjC5KWr4iAZQZgDHZ++o82CSHgbKw+J5oXhLrT/z2vRNQLF0EZ/hcHk8z
75sKpwnfD/jCNrKNUvFtcjIVF/u7+Tut191e211y9pZxb7pyfre4bY+FnIlIPAku+/YLFg7v/rok
Lg7xevG3XXmhhABr7TOiQERvKX5takNzvhko+NpHIloRw/WATBlxbihiwOwrH1/fPL537apYsGkU
0vIn6/BkSiJ/srYubEXjvjEsLLKLmzYyqzmGhfgcJ43/hkxtSQ9j+kFbf8I8wMivT6MWOJ+h1n0T
F4G/BYk8IXkKhgkt691WhIKEGrQ2lNEbI/BpXnovXmNafJJE47Cm1ZrtfLMqO5B7Adv8T9mgJFcR
SpXmFMSLDKhJMUjijmUz+HOvpuRwlhmo5ZBi4KZIALAHqWQvB3ipYcZIdyX1eK+CCqscw3T2btfh
0QxWTcX+upaTxr1gOvFrUjFZ0+HMYey4Q2xJ4NtVnXKkQMMhmjkLFI05CkWrKGXtZ/nKSh2JL1MM
8jRWqXiRlVUBC+aFJipTbIZErGVQvm12pgboGVuiULVeIIZrRAe1CGx+OlWu1XgAwWzVRmgvRF/T
g7iHsHgvuvFvZSfSfU8XlKdrmLBpWKW5wPI8nR+NwGuqjoVwQpHOgTmOz32vBrO1xomBvBzPJTrl
caHzCsMcYUq5vxkVH5rOVbB5r0NkdLUv8VBOu+d9/uv17T79SseUtzueGkOVylDftwzIEP/bhow0
E0gHJ7G08q+1zV2h72xVHGxSbuvps22hKbDtljo0ZqvBsbq1CTsBL3EvQP/6iJnpQSK0MGLrnRVS
yGG8+ljv3GyIXGBMDluahIHMTzjYmSnXjvd4+0NATvpFA3cBTYhSbQV1k/lKRJwl/hkLCjh+Q9Ka
WE3xZCMz/bh/KVwqEnhHU/KlpzBR+1z544jFWAcef49boOuYYfO4SyU5os5XuOLcl/LtLOVTK0jE
BLtKaNL2ylmAp6p//1nercyUCFwCgzBdixi9wchuoweCAmPFgLecEzAQFEW7V+FJZMweyXhvMyNH
04RVPhO5DTap3cDQ38TAOx/R0JRzlS3ExqtusWevmQRm+0QOe9XpfOUTX7C6HzUXBCYUBn3SjjUD
kmg6S2dgxVjPEBHY3X5IVRiLWBfFvb+SrOXlrvYFfmLBmMe4c/JnVPYi3YD/eF4V850Xt9yASVMK
OsWxL5Hn081DHojTudpmsaHe6cvOPbZEv6zBtO5A/E1Y4QGbThuNG+LQwW+Q1eTF9kqd4Nh6uy1f
rI81d8ALKd2+ORESThBVVrJQVIgqa0x/KEoacnS6QljfZtysPEVPriiMPRgvIKYCTRuGCzda71Di
gs0cRhEjTgyPifuOaGgnbmQVOFijMUSsMdq4LVm5gN6i0/A6YBIEKgsb3wwbgiAup+DWzPEo4GFq
Sbbdfjy2Xihup352sx2OaNH+Df7lAKvaJrxVux6P2a5Cqn/VEb4AU4Fore22N2Bfwhllth25+4r7
uoybrk4ywcFnsLxckgs14pc5UT1WlsNFLMkkz8RXasJb5pRWl0JqmbobR2RDJ0jV4IjIynwniRGo
TVHQwcXiHKAMYwIm0Zu/88mdA6y8AbGWANdYAlmfR8dIk1OxdOjRNJ9lCGSzdeeuSd3EjM2zaaw/
CB5LuZvTLgyAbZ4mK/5rLWxbB/FcuJfJJ2OddvZ5Rn7uz4DbpgxIgsjMItMslw4jhPaZLxL1eksJ
CacNZycG5mVGN68OgWBrb9AkQ4U1B54Qep4ckbJnUGgotB1+xhpCq4SscjWCuPsYBGml4IHz3Km0
CHZ35mGLnal8HipdfV1+XsTsW2e4ttMp6jXg4hx38egfqDBeOBxWoIy+6JUDvAVJCckA7tV/JXYo
AcY1kM6aMcejMcPxvp/Yx5GihmrJFsz0/I3G9MwK7hxkHkDLsTgQJK5ktlww2u7NhoYMmhwFUxXn
17yctC8HuYjeBv5kOfydZFkMOeNkfSKgqqm4O1Pv8qAD1mC30h7GvSN3uZzNwQamY1DaeZHLvBec
Dd9jC+4qEuWjTUoGECnsR4x86/S5nufw4Kqk5HgjFljmhl+IinNnM8yif3adR5xYLLp22RKr+OCP
DEaKmq7JhgUc9SfIKthqBJx6eKWnhkA5AW9BfAj64fQMQEsMLbAqvbCI4SksCfDBioWMzEf7O03s
OG8rFILRzT4IB7IawP9jFN0UwsXzYG/vdOlk3tdw8oJrPkxB3NM5iPKTCtFhTjrBM+4ZYHXY8dVM
1Oc6lh8f4bk4QRtrH1H1Ov/gXDjnx/oL3sg1Ro3y1Y/7q+rjYTfrP6AVpigoid45N5Jf8hljr8qB
hNJLAu2I8aYAx52ngBT1kGjxgO38enZ9uQ2O96fp7ACsN4AiCQd9e+PxFggj2Hhl7/NmvyYj/CSK
qq88yqH9IZOhO5TkTC4zns53Ag1Mx2qMa9vyBgFt/gaZuV56EMIY7kkqXZHGNKUiuQpKPRnqQey7
IfRgJszVB/snls/JvzDuNv+u9XdgKbUsZErQ/wIHgHvxbRIxQh86qc9h2qdL1PPGCYJBbct5azwC
ErCEEyeEByOm/Ord970KJwPQj5moebsIm4xfeUx5NV4zMz1mCwC3b7wV+Ot+OYrv8/Qg9DegBUC4
ey4tbfwoazLfCr/t+AHsaZDGbV1zFha6OI3HJwDwgY35kLr+JVoA+In+2sK6e/JQFB5Pq29lmAF9
EoCMCOXAAmJrcK+Rc1Tvl/7DTph5lnxQFI6ob7mkXUvL6Pl4e7tC1vf4f/C5UkkbYvjwLTx28x8+
ixi61058Hprwa/nA+ITf0n0eXTVYc3Gv5fT3hmFhjb1lHDyyaIpXMfoigr2r+t/R9qaVi+U40y8m
DbtEB83eBjGxZwr/O6xs5bTbhK/XZOLIDoem4VoYgz71t5Jd+GFGUEhJ4FR6C/4nu82/a4G3M9m9
TXubJHLAP1e+6iPTZH1JkqggET56VnjKncgjZyf8G/pIsBUIb7ZnkABz0jrBrTNjt/srspwcyLRI
5I7Rjo2ofcyRKuw+VkdMzt8GgdjAXwizLCpGS5/BopcxRH4xYhJcufc1dCDwJkaRJSV0MxyNKDKO
OMnVH2HNhrAC/19AazfO5xqKjJg+E0OyVncl/VuZE4STRa9h6HxIxFaKHb18gJNKw/nljZ8DGvBD
6xnWUSQD8Fkv1M7cECNn79Na/5kO5vVosL9gRSr+bAeF71GHg2KOzB5gS91vmVpVaAhLEFwQ8fsW
7N+l9Dbk/jlBEsaLkXSIXUYabFkSAsqujTA94EtHnhkPJ8nA5g8qsRA8+LZwhoRsMCB2R+jgcyoh
2Gx8X5M5+xQCrvzgDF+LtsJClwan7s7X132RSCrWWylYAbwNRFuT7Uz0kOzd9wNWG4Adk6e0NZTG
/eHwY6JvA6wrdd2MQs1l3d5kj1VGHP7WmLVCzh3c3Fg2LHgCEyXOt1qVlGHm5e+7sILRgrUHiMFK
SuBf8pkciVPDkE9xYxKOP1Yjc4sj7yeL/mkJ3RWBvRXQQO9k0jNjpgm9uNx6yehqdLu8/dybyg9Y
nUfA5Lr25BXkCcNNRovRLiLgHClgPOmVGIxwgbqs50rN1vTBVs6+oEulFhbV6eRDdemYbUvRUWTv
AKkAxViNbnkF06AySanRZhyHDaONU1sOYyCgJAtci2UF8xMBqr+MaLp5/9M2iOYvnDIt/iDn0/E6
+YJHzoFIEDXvhQrKW5BB/KJHBIoi8IPyYjWDrPULZ7YEq4XTcRpZQoXRDpaOhaJyx92USX+T/Dlx
L5ZkPek9yby7L/DAHbt8PLABG13eRqd2rOTKoP9R5Mc8MR7FAvszuglZRXiQPDUBpw0pReZkuL+y
thKDOtRys3b1HmoI50hgIIHDP+zLUE+oMoqOFP8EI1Hh4sNlVWQ2GIX22v021vbRBp2PCXjnwSSd
3rJ+rZEjCpC9raiVwZRUX9t/+ARppSZYLWrzgEQ35c4ieEM1ijCmC+Mjmzk8RP92Ng6a6BkBjxWh
s1fQxR2xNwxraA8ygeSnVzI0Wzm02nS9mRD+X2WcvJ/gJg/DcaUjFW3UPdOemxzs2vcriBTXYvAE
oOvMe5SDt839uAEcw5OvSYWftUhrP8fu7If9LnDbwOZsPHON/554H2x3UccUcAeKWF9ZkpeCIqGs
rSP4iKC/Sr+ks90dVHXc80NCWbiTPeeDNSzzSNtgscuYvwMWS8gy8Uwu4IsJy4hF06m7mFR6iShB
8ld9ie0WSX8r4Grv3Q90yVnPpu2MzmoLfLiUhthPzhc8J7mvDuSrx9emYY9OIrPTAEeD9jCUvLUI
ffhLy/KO086zHexbqFDrWTAbhLqoYFcIBHE2cIjGawq1uW5MWBYiRJEUSZghNoh95XUVHHHQt8rv
S2lwqyuLRHlYWJN48CcoceRaRxjp5q07POuqUiTPaKmw4HnWMSB+xYEwHi7OAtEviLZGD0rfcDhq
/ZBDDD3v/OTZGeEfj70k3ZZsNhGntYbQ9cWxOhbF7wVo8tA4NrQHXYTZpbVEd+hv8EwPxJ7g2cU1
8OZ3i+tD0M3jTIbeeu1sn6GCwt+tmkV2i//IzTqJaOqZC/I8qaLwwmtBlY8OpIiRvA7u2Y9RE7HR
22ILJkOJZUkh/EXWeiJx74Tkzkf0xhTm/msTOTl/4nFQiaThUtDKftOeV2XVOErmz4YVBiXT2SZA
VllMhty8I5Y0u8oPyGwjmsqVC/acJKq8lZCZd+chTsHM6jea+qhaHwCGRmPF0bpcGA7g6rjqbP/6
3/tIhgl0vYzM4pa4sqy8OAfdhtxjaPMxcdmim+PXFHeCsh3aP8tP6pU+y9a8ttsfo0mzPSw9J3W/
4KiDkE6AOddh13pTcLrN3ZV9vrcHbe3z11E7gmv4/Zl/I73YmikhJpiG8X0FClx+08GxgrYZWg84
wwjfTWGFmsyzW4F2Mc5j9qafxPvZx50/F165KuhxlbSopEezRREskEaX8Bkf0VLxRELeVfc4WA3T
TKykF5wFBtfwcgxV8boH17uZpOVZczi/Gcx6M/lHcUmUPc3rzKconcRCeLshYsBTF0/bOw7qd/4h
I54iy/dFqsXQ2Uj8XIrprOQGQkcOqGlSryXW4Y/a8WKwmIDFtmTNfbToqt5f6vmApmRoyfnW8Iv4
M59O6TgDpFU+NXx577hLaPD7HLdOG+DAVwX4Qul/qreuGWWGSOpKC7Vr86nkbajZEO05DurTK6O7
LqVx+uY5BPsB3PWfD1R9YIxr9D7dyV0JEkrDUP9tZdRiqXj4l1fN+zawZ7081MbvhQNMwW3ELFe/
XwsD5L8966SGubOzlbpCfzkGg0WVVynf1p4mOWxqX31kRgWD8Hi6diWiujqyZ38sC6K9p2A2ZFdF
p0nTGr2h9SUPkfoy/LmutPB7Johq+xC1DojJwOtrkxl1rkciwEs7zBMy5Viaj5m4WqYXxqYH2SZq
IoaWhJWSWo8qQebtfdWOFRfFotZk63j7gW9uPBRyOvpaoa/xXDo+eWjRmyW0vGlaeoEv4gcDv0iQ
R8aSTywUBFFx/oNL0oyqJ4Emhqj2TEPdjDqTIkb09kcGWKRv4BhMdiBG4ZqOjnvRNfm90/CgNsUs
+lZjHDsDNyZP4nvBXYjOW8WCWVvNU8xzVgnB4+Y7HbH9L5OTZWnFsxYqoFf+pFQkuAelaxBNLF8c
cVfbRHcJ82v0+IDSnFxdjCXV69w/YdZVq5Tgcu60JJhM/kjFYcMd+8Uj8UqNMpk4ExF9ChLdecIy
DQx6ko6oMfQ1PYKpXNffORmf+R+Rtf/XcPXPuuh6fsG8HF5ZFF9dZD3FzVJWdLk6+t5CVZDMWcI3
rrz0HyMoZkNXlar01ZrUN95482vjdiHpJicbztHmub7be7jfHNx3bEYhnF2HBoMLUgq/WEG+ZmPO
MY55+ntpPg2hZQ/8IjClPYqG8CQVZOcnDk6eZQfZBFvDlJjlKMlJicv5LIlkSZ5vywBCbiSRoq17
IPIXubFNo+YTt7+0gfF1UPdgp3pWnz4DHQ2t0BmQEMIEOsUEeoLT4bwkFvANdQSr9nt7sLzWCUhz
MwfYrJH3quPByE4YIVfI/H0cI2vUgynffK1FTYDkgo7uuPeEVOyw5DRrZgdzpKnj+g9fgWbGFPcz
axWfCtuYZGMJOO4P/BfW95kd2nDORldknfCx9uy/ipMudMA+EJDy21jnI2k2MWNStiKI3dOsawgl
7fTo/7PvGPuz9aOC7JWg+wpxFPLAnneY3qe7I/t9v9NAFa1ECQcjjSvDiQgMKOIDGL7Ex/T3XlOQ
7pJ73GP4mEQpJempDcol9rrr4CXdfQEN3W8hC91MSOQ3gPHORwQuUEUsNPVlaMh72bnj7ChbbMw5
0A7NUX3hjwvbEwHQiu6f9iNPbgU8BkObB5CpoOYBYr1pD0lzUKiYll3RGoL8ERT7nzSZsrNgrxNR
80qNfr9S3A7BlCKOl6FPoHFBdIUX3epfa8f1uaYjJvl2AinHCqnme/UYPkHFtzGXz4hLSR8wxNQ5
2I3NVixaC/4WJEYeaP0/IYP33Prr5h2bAmM5W1lj3MtZoUx1DH4dAkdUOdCe9RCQUTGLuXD1zlxu
ZhPNkF41YyZE28kKMZ+/vXiez/XwR4EbB3iWZhCY5oDl7z6NoWVARpIadC/nwN2nUGfmdqTlCzgx
0RXd7mKNPTGS5HeXiqOTv5esixEfRkACq9TbTmQ7kQyxQA7r+0qjDiIcy4zVU7nYH9gVKO+2+UXn
N6W44Fl1ifhVwN9iPP+nKzKHT7Zck5xUVSEwak8MNSN8B2o2mXxMeEDiJJKbx92lKlSQm95HR5BO
0RaSoa+qU/Zi6m7zd4nH21O1tp5Beniha5LUBR+KZgYfSg+acM5LEh1NGejud081xCsUYVgY8LT0
WR52Tyj+zZjPqtAVR+Le+Ar7Cf4iPdFkTNAIMRTa8m6aZ4rbcbwsfkVFP72qxIWqZMFrPubFvCHT
LKziHpAb+IZo8dQLF+AFP12v7tchBWtqi1h+FlqPiH4vG+RIYnOta+gi21p0pQL1F6hTPVxwqwKt
opQJiNDx7igZs0DMModC+sAik784RG6Z/tnliavz+XlxoKHHodn5VkKhIcqrfJk24eh88Xq8gjPR
p9LqnnhVdM2p68fQZAl1CmhaYNJwxu8/Wn47binYdiOY0aN5VCkk3OJVS8Rb6Fhd41mVQpuo0/7W
mHUkwRDS2rzjhh3MA2jj2NHubiNJM0fdL9WUYYPqsu0aYk9PWEYlMWZbPAfi8ms69KZv8sJg+l2L
8jiNdwv/eVVAm7k8B20ok5M4B76F5co6YshZbRoKKkMTq8/wuyLIxYP/Z3eL5+3oQk+YqKCJca3W
o/XqoJWGFvkB9lRSzK1u1gP2eR839UU+NejDUQEyi6tTfK26ybUwFFH/6OXBtKh3fBnsMzPydji5
tZI4XNwt0pGZfuJNYgM6Y4JRsdaWJAct1EfkdM2G24Sdl7oC10RGRWvvtUouBdPU2QbU+KDrL4jS
C5zqjRlHynlq9Ife6b67jVdC4RYOLeLkMdJAQ5OhskvHEW2YBe8MH85vjqtPMa2/vkSgp1ROYiNG
cB4NljnR1rNobJWc4stNA6R7CbgWfEM+NLYURDPZYN6vNC1v3Yw+m/Q8xmpKUUSm+UUQa858tzaQ
1PvOsReBArpR52hpEYz/P5r+md4dEIyInpck6Nj7nlx95B77ZOX7JJRMhWBVGtyDfkKRErFR9NrG
qCJGnPl1zmMp8N1QrMC8kGc2ekMqk8xY9lOAUkb5u9eZAe/AbTf4vDKm6J6ttwmNy2k6w4+t4pT/
fKMWthySmCoZxoGhL2kISvQ9spG6LNznCj6blPI8R4iC7oUDatXqlrI78mWfHlRKjMniVK8fU7gS
I9LuCtTQqfXAMLc5Iopw+1lUVUI75NdLqVe5YG5FLifVjsahmnc0qBsTt9ufcfhxycL/HzcHNUut
NV65Cx6vYavjw+G7GmqS2cpNSNAiRUuSoDtruUTKCuLhO6R9CKWfbi8/OhmobzACy/aDEjs+EOua
Nbu9w1Tl/7FCVouGhrIx2N6ZPlNCPnYkZwFY4eYBXQgbGRE31FrBfpDIMvfkGdKucc63CvK/6mZX
brSWpxJNN+K20wT7WPprQoy9bJGp47tVMlzAEl1cIvjFfFSRHNn4yNXmucb86Ga6wQCwjKnQ02Ei
lgGZzjBBw/0Erey15VOcnT+vbPZiB78zw7f/+nWU2/EOvuDxh2swvanyoJKlP1g6PtjQyfQpB4IO
Xmi7m+25bGhWesnZZcx3GRsONR4BnwRk8wXO5CP3ga3HaI5Z8SKF0x7cF1a3MV5WNJcu/liWSkle
XDGBw6rtjtXv5aNdWjMA1E822T+qcUuBZAz1ap6NjiKt0IuogQRiHVxEbQDcoBbT8JmVCq5QGNWX
dYic5IS3A2p7VzkyQKLm21JfEyx9llABJdsTV2Z6en+zEvn5FkhpgXTx24W5fZsZxdbFQFYwPH8x
G2srSKFRxTQa2TwvW4n2WHnfgf1BPrUsmVug72BAUID8iBE8dS+0fV6jEt68YiBexi+f+6Xl9QNP
TJH2TqUrQLI5XN/3IWyPsr2CFGa2D9Z4VClWDSrG8xbQ2pZ78aWtjTuDA1UTqN3yy4biBhfA4tJI
nWMYu/ovJwnkxvF7JhgVENxr+bsFi7sQFjGHNU+foKT3DUux7eZxYQIF0UvqS3lLeQUYfL/ERcmg
JFvOzCkm3Lv5UMoZE6naEhBhVRuwUvDPF1A1EcXFDVXQgPVECl5L70Xw8rDU17zMzo9JZL96AieM
nYzEoJKw9e7z7RY7Of6pQ8paVK05YD7WubnErkvba/KJhO+fy45IQrE9iyd+UO1iXdyrngCnsPcX
w0ll1biUMOhOZKRW0JFWVTEpWXJ50GySA8FHOMya+aDehy5ExeBskyxm08NfxlarPmWs2y5y2or8
xpcfJn1dhfvHbJHFFfCulLzavdsp2XD025Dmdy2HIpyQ3+iskCyfpECBRHu7Mk/GaG5wCXa+Si9+
XM/n4O0kzKjV/pGXRWg/702J1nCOR6wlEIdbunO3sOvOUIXxPYh73CsnDT2x2V2PLfF1MMR18cEG
EH/JB9MFvilfkcAzjSfG0ENVPUSSujYZf4pYZEFKrCMgZlWldyE/ZXIp1EFtFGkFtIrlnEEMFuge
rjVzGKmsfhUWa82uuzC+vVI+rV6J+D/1RWjGYPWMvKCrxcI4cWy4GB+v+p28R/WQ2bQUOx/QEyqM
2EubFDDZUBCbrHfwra9rnO2qvw85fHqsd/t1L1TAuXad9zIoiKUSFoKJGXC3tMYmudC7CiudRFSG
+irlIaIgnY2xOUwd0OXI/UkVeRLhGK21gNsR7tvzYxaDTeUH9SnYhXaw6JHQ20dX6C534cobMu2w
L8nyf5QIYkQwgKy/6d6ZziPujh+SNTJO4Yuefp56vwtDgKMxvbTej2zV9sDymtFV5ReygBL/MYyP
Z+TQgjgvpSwa4EIIrNcAxwLq0QoDR+1V8ktX4dc0k7hHousxOdlA72ouu/jLxYAIDFkOjF0URr5O
gxLy1XtxzxST1tgLoDxaeQIFOjlLBqcxBjy04NI7VwVvWc5EqLpCKNLh4/K1Hh04tAqY7a6/ziwc
TFT80BI8SRmAjIx1wrE6JD3XD3/GMPnZdW6I1IbvP+YsIMC/CfGiGlGW69VnwqemyH/5gxZMnqn0
s5wuiWl0gr61a4QW59wR8PXY3z2cKMwjt5PsFRKGJ+/dGe/bifAtBUs53BribXO7WA0HuEz/VbHY
XTkSJcIigZRybxDdjK4z/kbQScTta6yKc2OljqYyZohAhjuaZC6p5+PcoXHHe9Pe3Ext04ZkBATm
9ZYRvtvq7qcKHOZObrEyjJj8u6psmly76twqnFlvGkgu/CYrRWZ6UmG4NnVXw0IXkuvl28Iwy8R3
KYDiEjTEMAm1PrC/wwiCK2YKGHTzXnWZq+Nsq22bI3i5snZD381/nkD/bgF0112ESLAyV1jMRfN7
v0wcidmU/8GFfLDCnS1VfjEcRg26hwPdYfPZPNV93pF2sl8pn45qppAvwXU1/YVwkZyRDhbnMDIk
tlEO1VQqwTlOeSUhT/hf6muNlZALXabBIAchugvSOZPOjlhLyW3aE4qXxV7UpHvRvkvhlPAlgJnU
YsZTrwGk9kRKpK7oiU8rJFGfH6CyKI1tTnJQtCtRX/omFH0MVmTgPykEBGft7d35s5OhWdhnHNGN
pDhsV8ShmzAI6p29pjlQmwFLUVyLrp1zVkN74ODL9c7LN7slvENJH90tcAeWnV8Jkg6vnyZqG9rg
aS+2OrhOllky3oN0ltxKauIAd84xVO6I/Be37ijBpvOOhU/oxedYSF2Z4Y3HAjZHgYL/Vl4D1dmf
SgYsRfDZCKNReTIGcLJMhPBXAqRLqUmZ7fPshtbqsmBRLZ5TJaE+A/CtIRoyiCwhGMBblQ04B9J7
1JAcuXkOJMsFQv9HIew86ayuEb4ziCQ2QgvY0LaK5tLtPHiNsdLMfwQI1pwpg0KNWDVSUCV2EXPs
LkVagbueSqGdGjyR2zhF4PQ8KDZii8trKpR4lwueZE3qyY+x+yt8SDKZo+/mnMvCz3tbpJNIj/ej
hec7J+xqmYAo6kHKPDhZGrvLJSCusOTNSQc5rgfyQrNtaognZqaESNyzuZnTzqVWS+4w9l74/6At
IbUETukRY8CfaE491pr61foDEKA0oBVQIdhOrJBaGz61UaM25hKPhKplIL0c8xwE5xEAplO5joDA
LEFaCrrf3Ij68mjQo9Mt5uEh2+U+UlcNYLVviu3a9gowDxNCKkgegh26oUoLlqBufuB2jhSj8a6X
aVYVfMaY+c+BYipUn6CJ/eHCYfkACBoDPeUROmDyfo7TgYSL7/nLPntWCmPUN0Y4YmBM1YQSwLLt
jEAG1lgDtTIqCP61X9L98g3UL0JoHrpTZIVihIUXtMgwl3nzpfaIBRhpyfXAbEyGsFAFjGnKCW0p
9O/j4kKo/RwyBeOtnbGAQ4Yy8N7wJjv8yWQOIimPWGlGgZGB79B2z75nNwTJW23RkBhpv+/kwrg2
iFdtCePDLiwTyirRsro/sDnNJHZf08gmgRM7B+7sZLQ44htBqTuru+e3zRPnDZluMDz4XeymApwW
64OYdNArdVTPw78l6uOz1jFaozescSjE1HYGQdHSAm7sVSR/A0RT7gDhNR4qZ3r1iTnKIomCIU8w
3LORWwNPVjtAFnEkdQvF5R/80eyxQtGronrEFoII46mKEWxzYGyzwJDt2IEv6n1CkbZDJ+seCZ22
qtMdPHAYYZmYyTg4ejEbUWuqI+0GzbsIBO/lR5zpKqP2f+UNaZ3/FKh0a3CLmQdILQihvyYnf7bu
z6uB2BfN0ksvJNjQs6wzsxb7OcJA33gVXvhsXe8gJL0jcucdhAfEWB75UsN7uMKgjO17EngQQUxD
eLKYh01cgqnqEAQk6E2m9YVrYjtqiOXh94bkFra0V1+THKtdzF2S7RAlVy2aXVujTxfuvE6/Ylcf
qfeMCmawc+VPsYvzsSwgH2NxjcetOhVP4Ood8LDPisRH5HgIWUianVMxMgY1vlYL+Ywj5yc7/wAK
N+KkXX9Lr3AczKgslRwv2fh08dxiXbWJ1SPpOwtF6KKhLTduscPo719IRKnyp2wdu5OJm0BMHFC8
y6+XNBpNxKNRK8IyyYY1cCWgk2+dC6m+y94FCZoOIA7/GNni5U+lyijKgM/i8q0lHNgblkZhbR/e
f/jDK/yK2jaKhqBfMPj+lbOYFyya4eL+UeUWBykhXixfsxbgFktcL8/zkn+RfAb9gnG8fssoMT/8
4sjTMi4h1rl/pqN2cQOaI5IJWVd20uAHNq0UQzN1Z/jnnkRlNSacCxrOn4gJORkOczbQ7EW7JeqI
QotNd2+hr3f+uSVVQYnQbZUEMz34iN5P6gfaH6kOdRqj4m3xOGINmfbM/4G0VPBf4wEwpOvM5ilM
27SkHv+RTkgIJgaNSUsrLiPJXw9Id5+HWFZQ1kZ7rOc9O4TAXJFG+aQF1SoOKBeTm45sQwpXv9n8
z9e9BN5Ir79LIvvK6mf6RT69YvRmgTZ3+QMFoQBVFFNy59UKE7gMQxkLJwPAZz6+irDvqEPdjQmP
6BsOeslG9BVksbweKX9L+F7PTdOTc4GhBFcvsLqw6FFZgtaQ3/6PWnRpeegLtVUdLLC1B3f3CMWP
O76p4wDM4emF9B34L47pc2k7D3FuB0WrUPMMpNbws9PTXViPL60ixl+IXI1JoziFJ6G7t8L4QKTp
8kTV4XTjX4igLWpwcXoTFj4lBa9yW5fRpY33exQYNzfqbP3SUZ44hFGAKrzmS3NB0tvfSEki4uqL
9ogg5h4rXpe9e/in1JlTCByjDZwLlXIzryf7TFZgULXf+1jN89RNwrud89hENr7p1C4Qdb36xlp2
Mom/6c8uwZAU8/O1e1AEPNDUAmxCro0YIhM57NKmVzHP+yZqobMbEZnr5P7LWJUwNgs666ZpTthP
SPZrYHYkpM5QOwPUGAwh7ZHBHT7C5omZaHDzciA3FEc0FmNWWzIULn3HhrYowYOsRFwSc6KbAxbP
tKQxDl/n6c9WZKO+Htyi5Yvb5aQj6V8g+Sa0FK0xqQHBk+DgM/fSDReaOmQG74jwH+/bZwwA/t0R
WaBN5OIOk19aJgOX6cqMBDyaFsf3G/808KBmTN3GLu8sLqlG2kgKh7kYiuOPasUlMxuTL395a3U8
NEd1pBPOo2NUcUD3+y9AQDai5zvlJS9pI3tMU/UALRsu1JB1c46qotEDE7eSeAsHjW19N0q55SFG
1Wr5hrLSxNX53e5/2MGykTCT5V3gjIX50TkJ4oLqeTch/mMrrUgn3WIxlToDq5Z11rs/gnEk0np/
xGq8Kjjr6Z3f9oLR0cIeaxHa+F/CnOBgTPcVb3I3rPof7E5IGQqvPmu9Iqo/60pYwMBjyUS6yoOx
n7y/zSLBL0gC5gcWgoxWfFmm9XWJRdtwkCAhDZrL5FaowiUYvfKiN6r9gU0bSrkk+YsF8ZxMWEQZ
WAUYCi8cP2GdLNYhaKRY+o0DEAf9l4HMZdWsMpGNZ83viFzWopEjHs6wq84Cb4CudpXd1sNsygL0
obj7LGTFukOrdE+YrbIkhXxo5lPFv3Uh4GBc4InQKT0YqkuMa3mqZn60Vxlwqv+eKOWPsgXaMTXS
tAC7GQSnh7I75C4TciT8nSKjQlFHjbG4kjUDETpI62rMFC6q7qVQ69c5jLXXL0MYMHWW8dyO7szn
cOMGtFUMrIBqSGqZYPHFSfSe9GPqt/4cWgx5n6U3vGz7RzHqUjRPhaecVOe6nu2vFjfZN/nmBIgd
YIrpX7qe3ATMmIakU2AgNHY4+nDcT+Dk7rY4HHPDih+dwoLt4qPswA79O+WzFr0SlVgLnSjLqzQr
Hk7gfHAJQvqCX46GqkKxFjd+nO09FKm1LYlEQqVGz+xxO60U4JyTlk6Vi9HN2jbK+DXFh2hnKvnT
NAGBwdZ1Yfzwif3KTB51jpj/ck7E85gfoS77ReCx8Zgmo9rlMn2084zQRb68qMz0nD/aOcFnIuFq
tEQcwYkn+iNRBQ6GJkpa8jEwFfd1rikeBVkQVpocapDoMGcMeftpM67VGz369sxLEukYWcXNWB2/
op7hS9VN+Nj2+nP1QGNdU7uuSonB04JPMJM5E/MHXxbNC25he9fAFfe7yA4RLvtrnQElBsfspwdX
7+UxAbS7fEGSrLPw4fCPWOkphji124DQULGYvlfgAyr0LUa5hDFTGIsTX2gxaIBPGxaDzU5vxqL0
jdDtimkk3NDqnp0sr8eev+d8z3t+lHxrMxp7+0D45zKhtjol6jeHBLsghc3kDOhoJjioPFopfc6R
JCmBexkXFpqAWy/hOR5Yc54CzQAj728TYJhS4cX7OdLZGd37gMsKVC/cNJKf3v1l+e1rnZ3SXGPO
qqAnAk8clysdzeeW3AWAwsbduGeilwCisNuoJI1tIbS72PjqwGtxozI4D8kvBilYqpqDYfpekzGa
0T+uPHotGYgsYuJhWPPUzfgrb86+TUl/qdN6wDSChKnH8OTLLF0nGz/zszmr9DGP9lg0xZtUHAp2
o875ZujjSl7jhfIiGFFHKgRjLYrw4LUnFSvHHa90EbUw704Nsut05/LB7b1mbkHiLgo/I3adXtcY
rfNBy3t6sBQsXsRTMEXBloUKMtgAM4v+kdXc2gGycoIOP7DH2SJAnXPah0BxJKysw4wu7++hdSM0
goFOCTWFH8bAXnct4FtmaB1+EnjhSCfOQB8QjtT5eko+cd0WG/Ic+WJnnCIqm9htdi5ehDAQYfoN
LwUv/NjAgoMTfHLuex7B5ZJM7CpKpc88qFvhdK04QxG9Z/IkpHStgznBZ1HgUG2FZnsryVJb7x/e
/TBewnG8OrNeYSWHbjxFw44P6Jw/1bSjqD8RI2L5DUmjg60W27cwIjxgzlAue05q6dOJzuE8st4k
kKzJS7h555+nDxqWuaz+576R1dxOPn9+Unp9n6aTKwT/2hP1iwA55X8xeQsVO8IO8niINwaMUuid
14i2pWhrnsiCzWZb3OMQAj7I0pwEnIXUr7vcgHELadXWIReU/olQBKw4WYq4rFPGe3kwlxKWS3O5
mA5TUAZm+6FD7oxRfwYaknIxj8vHWuc3p01nGiVhv/C8ij/iFu33c7Vc3jmpCiCN8is0BW2Nd008
GCnKbaBwqjN4GVq+MvB5oVzJYNHGqFBKG40GNMHhBVX1N5yTVTPZsyFZlxjphLtZos01PbMRqXGU
a35bmJahQN0o3EF9hJ7Duq5+AwnIDtSAXRkSyjyBFEzMIr5XQuJm+qeRh5NVieRraE8G4QQtDD1T
H4S+WsQC9HChRbgqx6tGdIYYpa5/t6+blvP25mrV6oef+iN70CC2pHcwMekyZgUxnmmahfXqUxBG
G24A4ETqsNdc8hrCuWpbfFzuZjDtFSQKyuqGPScycUIpOKF9zsPVrwWqkcltZt85EbY2XOBPcXNW
SnB3vAO3yYpncLHSXYLq55rUQIam5BLIFKfZ2eX1tMy8RtbpfKoFkVXu+XzwJ7HDX+yesU2F/fnf
hPwZjsyVeEP08/yESJauJu/d3XFAQIhuazr+2a+wrVsPpBwtNqkK5O/0PDpJvwqHOCYCM4apCVO3
oNH0az1LSIrCUit82zfOHqlqS2iFVAiLc0gxzij3C6S+4hD/JCGdO7xPioos9gzviKUeNe623TBU
MCcLA6c/22T8i9Sp2U7SSVNVZJTP6OvDprjE7sPUFAL1FuxBEs2ah14hLC3LUAP1HxbjnavqCUbu
x5r31wpBJ/8qrRqk0b4eernLXY7+F3r5AO1neSM+AQzRK7shpcSyOqON/t0UwQsqo22sacBBJ8zX
yOYcO2BXuNH8jxgR4np3teXG2ESeEi90mzrCKtER+eZkz/UymmRS6QKlCPwIGdD+XjXQzdECeY8a
jw6GHe3KabPbzF90mO7rtoXIsuZ9WYTIPY0J02atJx7bj91JPl3Y7L3yOrCtqetboNcL00ga9iKY
CZYJKfsaasNNeH3+eUQ//6Xr5SckwBqgRQIXEhi8VoQOWBI/UcXBFVQFlCrh5bb14qAmzUbl350g
uZq4Kn2E8oIBRhXnL+5I2FZ4RPGtbM75GOYW8yEcKA2f3JIl8tAxjNenlqiqSB+dLQKFTHPeRIcR
JyHd4nzUzAGvvH5GoZRpvrnEa3es4xoEUY2eoZgjGAoPW8Gl4e6qJwVovoFMfVVM1arlsZSfPcid
4EPcECv+UhqnG+4xuKsQHnmfgqmZDwqqgrKeCQf2M3jUyjqeG2mImOhR+D5Rs/iJaqJh2v4C/Ey7
2UX9t8eguxXsbjShsL6sfBnwYxXdkCPMxQ+bBD/Ma82/PYvLY+XmI+iksO4a0j2GgXdTZFDPyX6H
6M2ngZGeWmjBVOcul86plz1DNW+W4oUUm3mL+0h1SGaVLTuX3HP5/puKr5kWzilAl93zjD73imhV
XklF1IyeDnAbKkGa8z7Ou1XVYLcW1EF7YMUY3moTNtx0YVa07JgCRfUv75EKTQCGxoIbd5U4iP39
W4+EgY5xs6wE8ls20IPBkpFhDQZW0J2vArdwFJrjj/UmB5ghaKK/24N4PsJrnuM1eTgnNHbPplla
LPuxak+qjyVxHvNlcf+4Yd/3AJMXy8QpcJ4EeFYPSSZwBOe1816KRB0hyE1Rkm+rE1QeO2SxDmwN
OQ6rVtjjqOb27q66UZuwceIZZjXZOSbq+TGA9MqRb1MZ2I6kAY02DBfM0UJR/EBw+PMFeQqT0OMP
H6isehad7W3+0vNz313EfM3uzJLlipBhSvMkGcLEtEOOhTsqiYQ50euF4/zzf8d/SqhQRdN7UKBr
P3UrjHdn/+M8IILGaRB046i0XK8LdSwMY2QcjvW6xeS4h69SzXsEwUKEYSKT46ISF4xIA92JyrCK
khY+fNj4EMJw4O/TtUevpfj/Q/BDH3PAOhoLpmgTxTs9vYGU9cFcjsiiLgrBL9ov4tSGZBLnOSbM
SoTIpAqudbvAYFB8lw8hkJcclF92swRLnISOMyiqIPDS5J0aamcmozneglnu1lx3gkTiPap+Nsvl
TFdzMLaLjq6RjZc1FoX0YZVBobi46+Ut14GufCWY/EOjAKWiYQ1y7NsYh03OpduNd5ujPcR+nhAu
svXe86CA3r+SsxhFjU7w0VfjDKpgvKgpRxw1Qwx+GEaXi4pPasGWbJ6I8H4FCc6F/IMgf4KSZM+Z
Vy41TJC4lXXPPM3zZW53ZD6khu0kOLkaM2uDficJDn3kXwunNYgtcaZTYP8GKabKC8qZvpUUbrxl
zPlldy6FLLiyw4cI01RKZCOloKXQylA0aqa5ScykOV8B32JRZ1HPTwn2Mu99Xn3umEUY8ljgVv1a
9XblJ/1t1zOorg0hoP8GAb5PGU8rsEFaMFQbQOroUPp58j6pt7I7i63JmazSyuLB+46d0mfkxdpK
3bmjjGpF4kSoggk9As0+jBOkerDcsYFgTlitYff9vdnJTQoGITzGCcCU4tPOsEt2Xj1Makb9fDDD
JqqE9V3aR6pXSFR0+c/SW+X3LuHbzGX07YN0XkCqP104+TrtxDN9SPCSg1OQBk+mpFXEliC0Gsf+
vvgKX1GT6XalZ+MYaGIygGgresL9woSSyeq2ML/leoDfUXC4gEl/sCzOCcBiXVc5BB3IECB1RcqT
Am14/0EvR8sMDZoWNVjW6CFjgR1A2SkZct6EHbODl7ct2YUZ/MtYzqwSR+5uspiQzMWFROMNRfcJ
XpmNlADeaF+Uq3dMalda1hfCMzHSK2b91dB+UHCCpLyIPjTVZtxvNiL6iKaa9hDyozWjAmF8e8Pl
M4ZsnF1OmuscKuvS011THniwzA54D0UlvYtrHu1GCE6M2qqkumvW6Klhk1MHHpAeZM3LZJshCQQV
YyWu42Gr0i8DeXKoUxhBeEmF2YoWiwUt1b/j8qSqrMXqSfP66fIP20DKGCF+Ej1aab39HQul43iC
mviF04eNb6KXnrdS7BLEcuXEv/uDRe0bgL9WeIvr+Ypxsne3O4CGHUZAbIwaRYpHBpgO7NueIc86
mNJjJlsP4YdRQXrr6CdKTelaN93Oo/iZlVMJvgQcOxclZuadn3X9AHDM7137q25iDSJSCWY44a6j
qWavGBJq6Vnf4Ok4o2rS+cVMXUZpR6dMYJa9FHq1zgW4Z7h1/+XldJ4sITBGsYKka0MSTFnGwrYu
5m95F8JSI5txcMv3qbUZLo4mFxudfJhoQWDBqvhQ24oYc+i8Mqvb0JlS12VfHCLMM5OwykEHgN2l
f7bjb6IBfrm029GVruwSfY1gXWvUBy7jepCUNZzEEVOtAgIbIcLvPLyW2qDT9sodKiMaIb+Rl4WP
j8HOVZbxOKDP6AWP4OKNPz8WjRjRKRlneiYiK0ZuXoudGmuqZsoHrAjWA3Ln2YrjuCtnXTCvS4pj
wffY9hSGttj0tXYX5fq/cnWopA9ZLSo2eBcaNc1CoKePeO43hhwpLkBQjv7rAJZ7gZMHRuM2mdf/
0ADgasKuwgDpaseIARuJO44UkjXiNaS9diTTCafDj1Z+vs7zjjQfgcF8eQF6VUcxmAdhb3mp+B2Y
/SO6Jf9leYbI7vFkdoHXZCHQIkOdDWyl8DLnglFW71ReUJqYVEQQkVgUHHIdJI7fuw1lpeQlgvry
Q0FIShb07tOVqLG3vI5RWPjhJYLzbzeFhAvFTcLyvqTppEwU48DIVBCWaPNOabZeDuzRPrTDcdwo
Qn8Hv102PFgXTJX9ZI7lvYEI1TOj/Im5NkY2Gq5PMsRLsXK0yJvnaazGsQRkkit3Vu7ptGqiE+jJ
8MJXCNimOvAGMvfEU4RnoxgYvVGiUQVOGyICmoH+p4x+h62XGeX21pqDUKs2CG8Xn9YQwIeW+VA3
y+H1wxLaOHPae6kRcm9UtjInazfCQElFTEEq87LK10O8uFpGCqR/hj5bSOSfRIOxH/iOcph0eJQX
ETtpv3YQzPqvx9260A7uXPO6TM9ueMc7jMZw3vkQ44+SKgWl19kbINfCilETgU5YzZe5hu05Cw5w
13muoQkEt55b50IGD3TFM8JM0G2sG4lZkJADJLNW4cpK3Cc4nYElcEqTgF86sMrVEANH9XVIHLh0
yBsvKVvzmG8Td3rDKSgLKVzIwO5XfVdJIIkq7abfCZG+7MRba82RQnpfzvRNgLDD1BkeIb+uchIn
qk289/lozCC3zrkfTi+e3VBA78UGaDZ/V6Y+9n1UMQe0N/NruLTAfbcMy7ClmxCeOHF8E9wS5ry9
qvKOE5Qb3v8HIq0UhniuDB6BD2dCbrvH7yZTQDsIb7lkGs8mk9R+IMkDHAHbis8dJH5pb+zGtFBX
SHS0Y0MslaJD5PSPy2aRv9lEV0V/xzUwU4CE1AjYwcr2v/4ErbJYA09PxYHlKydyWBN7kH4m+yBB
TSL+2BAhThWuK4S/qONx0CHhLO890H7OinVNZRZuwJPT+o+XaVlfRBtsOyYDnh09AqG+6o6kFupw
P1fljkuscMdl5lkzUu7Pmu+Q8q0qY4p0giMXsM8ts73uKRnBg93e7fHSWHlS37rqUVB0hnyTRO4O
iTQ+8OBZWKRi6kfxGTgm/c+YRwSuxcmFpXx6RlH2w+eprVnwAfFoYaUAoN+tEqxzWoB88EC37KsP
S/V632QLvCCvMKKF62kBzZD2GILd0h06O4KXi9ryKFSfX2m1TrLp60u+Sd5U9Wlqdkbss/Zd2Ror
4Dgm1gCq338iY1zaAMiQcxALsxAFz0YTmf5vG3/eD5fuONawtEkFPE7aTQD12gqfSJAAh/EzGLr7
3DU2OkoaSosINlMBVHNLDrRU/zumfOOGLX9mToPTXYhZlU6JU3psGYUyaBtJvQTvpEIL5R2uvF90
EDFQVN0JPftGdL1curJevdu2URVCKOFdbHr8jJemj7yiMZISKpFiLiQiccILETYz+XCLaa4BXexO
TvRFyEzhwVRWBtL73ZNKIYOxhG9ufkFrshlFXqtE0TXLzXmdn/X7RtoB1E29/oEbMvl6e3cVPGyQ
YsJjN1OfedrUZYeRIU1M2DtotSClXvxXvyiUu5D4CPwssxL/Jl4tEqd1ITmhG4K7xXX6Cz9nulap
f9845O2Qc6uswniRQS1j3mW2M1B+OAqR3SXpPH0W9J60UIQiFl70uiYwzaV2PbfmBXdDVhuGmfVA
/dyOABAOF/jIh9acLRI4kv5k+WNSv0dd0Ob2XZQ8+IGFv6bXqK83Hp4zvpnUMWhyfrzIV4khE9Jj
fbCeiQam5YcjHogamm7fEiTH0IotjnfrnDIiIV6PhBDgS95FfvonK0vz4p4pRKJIrdQZ8CRvPOIR
l8mHIZG8Oh3aLELkmTbxZ9c53DIGtl0k255wJUgPpSWLzWbeWbLSuSOpIZI4KUUWt/J2dI8BJMem
4dQmzwZaGOWbGpaFyORTxIYk9dnSd0MDQ9NrkGVl/YQ0WodOmSy+QVL79vz3MyhXPjYFaUusJQbg
OD0OCCMhEx0dyPYuHZL4fZoT3bw4/vUOsSgGlE5mFoKmXEAfMZqepzr3YQJ+2Slhr6QhNUnVuV0H
7XPXBWQOCbKHR/gMd9aHMW4hVvUxnC4edBu4xRFh6yrsy2pYssF/r42BctxSpgbWdxfPDVbmue6a
TluT+3UJhf3gBzdZU7/PJl6z3Mmp6ubpah2pp4Ahm0lZayGmMRVLtj4WBT4JhGx123zjG04gYwYG
YRedMh3GILT4bfONWjDpv9bNrfuXb6ow7mQSDNsiyXXTBuFmbe7hMvUWvw8KXxjm8+V6YYW+Kfki
09qeVeX7sAzg4sKSbZT8d/wOmqqudnmI6DsP+X+u65NHWpd9xYtaUdzsRWnH2TjAqxmSwDpD3uk2
TJJE6qLfZ3J94soU9FtZFSspfK4KUp8GC/XJGRRVY6uHejH4wcG7V8zJcKNMrdH4Mg3SP+q96tU9
df6Oswiuqp9pIXtM73BVlQ3cfRAJrf9ACMMUQtY1ImpUo2YAmIoeD99EA67oc8GuUJxeK/MoZkTX
netCO24mLD+BYzbIeiakxLvB7wTQw15MMF8Prwrztrx7s8Ojlx5fUtVNA2KMkzgHeXOffcIfVkkh
L7BttVAvjKDdEE4SkQDq3+NA+2NXpo7xmDWbDSOBBVHRqFBi76fqMWjHrDSlGcXU5d+s5eeA0FaI
jOe7Fnl6SJlk9VyJGhfuVvOWgqPGjDIyZGMy9ho/k+kv44uOhwxdolEuR3/UX4jWqfBXv/JUpeV2
Zb3YH0TzRU8Am4j0TS44gwqMxhXy+flkL6eOcqW/8oX6SWxjqBkJl54sLegIhlkun7/8Go8fQYk5
WnFxLbIX9vw3uzgkYmDwkO3aTe9QwIXBO/TvtNPTuzalY4TfjQfVjJMtKn8Gf/NU9UDD+QB2GLvS
whmkKmTeKoEns21LO5aiuWyN2P3zU/CIXp4RztCtEW+u9X3oTGrTQR9gVTZ+5+KKftnBmFoPwSxs
mzv8uQvjAP8YPzyuuWXybYDKutUMusymucjfjdttNkOSJYLp3t9d7oTKNLky0I/t6EMx41m46H1T
4TiqsTcCmiSkln+gkXfXP6VyzgEvOTueJBa+p8VQX9/oaVUfkWiGR6Ruz+Tnwn9ajTfYyPZbVsjs
M3FPvkAGd6NLspMz5Kkw9ySXV/3DaFW9SnjIqcDmxxnm+CptECp8M5StzrCkHq9H+FMjnxJ8bTZq
EeKRTKb2Wt8cArG7v3WygwRaANiJiusMxKqrf/yCswlAocg1vR7T+QU9XXWC08kQS45E4raR5Alu
A1WWqSAjHCc2MtoDObpe5VYAD08uZdhRjBoiEjMtyxrkHeQi/dOEO2SLQYDjIR/1ZGDYOnALMpxv
GXb95rdGZd7wmFe+H7taia5sLKYtRPszksU44CdY8TuDVprqrpM9VO5WcuRPekfoWE35Gf4XkAWg
pNpgzrxhsJCD07lebkhURcvYaDNfcsVhl4fQ5toaznqEaOVc2cRvDoWITgunlVVb60gp9nbfE91P
A2sv355arorTH5DOj0xMbmw+1KWPjUC4RaLDu3ZHkyZLYBJCroI45OrxYef+J73yLwoQ3E/oTi8Z
8w/VUwB+uPrRLY8eLVNZsv4xhlJh/8M8rTDlna1HRshUaS9McNt0npkcTfNdYanrFJ8nidFMor4U
ERS0mYEV63+wWpX/SFgDBdd9IFszyt2vAtltyn4NVqCBRX977gzq2aSPbvPxjmUlo67WXL1PKesh
Mok3ighd7ZEsBZ1ajNlpFYKhDroq9Zj/QCWu7tQ/lAG3BBKfytnahCUCA5xivh20Gdf0yJrhIeIf
9fUHTagAuzim1llCGxD8vDxmL2j42U/XSm4xBNvUorO/jQ7o0tE9gSN2Q9lptCHMaT7O2NpHS8G+
iO/PwWlkv6mqOda0Rmk/ZpM18vIDdXbyyjzvx16cQiy2Jhmw0CxkRQSZmxQrvtZQ+0bTfG0QoRSk
bhhiNgZA2GvLQY6szh16PH2sUl0IzkttRP+t1sBpqhdhKdrjFSXxpnbKMlPvpx/kaZJgv7ZUT4UV
Vls6ZJhrQY8HZyHYoqbqM3LRrR7PohF6Urnn1Pls24e55bg+xXAA2jYGPq3NxYHqoS+TfLMHZh2k
Rsj2l77Wq35E5tncNfEKw8H0n3b5BEcrBpBSybn+jvOj3b2IMeey1INkzabHKhWURRqmtLxrYbKH
+AP2z2622OEw/GVILfhCsrigl1t6scRGgGiUvVNZHK/s/vMOrJJwddd7kChyRw6GpFYfuKx5hW/p
WsFEADFVUrF5vTz822GWmS36o3j1oVqkTQsYQV1GgtYJYwmQIt/PtdQdIGDvAYF/xYFU/UJePG5A
yzEtHJrPiqIlTe4u2nm+I9wQqAgZYALwPW34TC04tljnMWSSDDhFtQW+DVTykkVHxuCgeYLSJTo5
oaptTOIGmjX0Hjdoned0iugKPXx0EJCP/lRfgCNIHGfw5myA8Nu8OuVgxN96CIQ//7spnJ5BJoRA
m9jk2OXQMMypF3+zCvoJohFgEjasg51GHviuWTnOff2zZDohciYgsS9BFKWhNfq7SN3wzhPy/pHb
+T2wYOpvb3uT7WJNpbecKWv9eLI+i2h1ujaxFwCChXhn2zctlOYI5ZJN9P3WA76Dmj4ZoZegxNdT
tvjv7EXEafRaPWqdz7h2mGHBbbmUOjIuUBAP0d4nfGNIACa1TGGztqxOblXyxO4DCI+T4BXozRZB
tTBF6KvU5p2IOOQF1f2TJZAI2YJahsF6KIIl4CJNq7QxlupKkBOXoohUScVL5ts2J/g9z2faFikb
JYvinyaT16qsSoBuW3eLC3Sp4w/E/1TwWhTE3cnXjWISROrGod2FCp8RVS7HZtcDA8ISAy/SP+eV
C8t7VIBMvwGJV2qdyEQCHlRYBRAfha9qcJHTHoIoGtgKvc/bz+8a84D/Gbx9Hz1XPineX4EZo5Js
a3J/1MC7XkJlHsZHtFUs/f5lBWHDtm6191cbF5XbyK6vOeJWVh2wCi8bzhC4Ndjv3XnADgXB4UxK
fRSGgTeZOaZ2HkmctxeUkQqWI+b7vxAHSTVO/etAmVVo0/Ytzg+Dgs8lTlwHl/Twx306sCKV31lK
HHnVIaPeNOSHv55H8cB+G0fJAoTYGqrWrDEQuVe0ZAsc7vmF865EkscsMEC4OZjkRTRqN+51tfBj
fO3sEyjQD1oDngBEzjNtz6GrLT2I73J7/I19YaZ8Lkfxn8EDpSr3Thgqcv5Cyk0yZoWPZwiy7ibc
+3gz13ova6UbwyRjn6VkStV8rvneqdeyBlQM02BNQtmNWw98mOrWVXybK+PVCG2bpGMhYuE6LrES
2bIGXt9/IQiJnfdpoNamX20FMBZMymP+39GXP6zzTBBb6FQO5j5WjwCenNw5RnYgGYpf2/9XPYdI
Lb3HNvwB1mryUs0hSQx6jsUbpEjrum5jVOqDm//WZHGhPTVo8i5+AUaegQgFNhMGaEAbs12u2Uym
qYc9JApOeI1l/wgcRyxjbvxhgYBHGnM91ylukXkSiASeK+mUpo7kSpsH8tutQmtaBqwqet3cL9AV
+hbKfVuiSo3Uf3jVH0YsvGJczxSIxmiwBiBqy9Td/miUAKpwHTUL4uPFCX3Q0Hnmi51VEE/WmyfK
w1R66MlK5nRDYl4Nwiqn8Q122QuDHnzeYMcm7G4r7uJ6lA+1vzgD5xCw77hCPAKZz6/5sPXol64a
Djglrf3IO7BqJpkfqUbAA0GXgepPhHvlVDeW+MbJTPFj63pUyu8pgJ1NVCt/Z7cPJxWDkceJSsn5
TSdVX8tTY4Q9DOtrDnILiyezt6omHp7EDdYlCrVD+8WqZ480MZNQqa44KDz63fZIqgb25UcuVqTX
zEsOpaK6mSNBJGt3AD8ucMHtT+Vl1LjMV3exOERK3Z1LjvlL1kT3Edr7MtoBJ4mOZcx/JsU3SKr+
EiU/JEhgfk/eu8tybsAy8vou8DUzGKVegUY55eY/Vrg2sBIpVXNh3cYfmxcbRZNeG9/N6pTKoly2
bI/yHajDNlXhSBR1P4nuetfpL3VKckVypOTndPOt8FbOt6Ef8ZwwWQpPyZ+eNipHyJ4jlf5OfPN5
Cwr8HaS2ViVVGRhq9V4LKyXQjujZmQfuapsXTXrO3ZPnhIv6Wr264T0/RTLRNr1588R0Rf/J5ILg
COSOiWLGhEjikP86wq3FGZcbvVJVjoUBAhflMnNpvQrnJfxkVV/AaBfJGyYdb4vDF+qTULLZMq4q
MI/1OSWvRcTRNRX4t8qOtsMw23Am4qJpaZNK0NjDerb/kdN7cmUK5kHOvIbk62OdGYvOkv7Gfl8M
EMbw/hzJyYFrbXUqvsH3/wud8p3biTwkdn6t/QUmUlRxc1SbXBG/+Otx7dBuMaGtfmKN8ctzE+S2
bvuD+nmFLARVco78vbGE/Z31EZ+VJfteqKMSRaoWjkBdUj+j9iA2hagwtraXj5XGGFvSsHzpiOQ0
z4FHAGW3YBGR30dHpkTsdMYBhCwNo76ECcGNtHGoQLvHU5NFtie9yLY5tl+SNo75+nH9paih1TT0
LF+S+/69WkthxU73wemM2YyCJL3xprbI/zaaChJz+WOPZ6kQ/OoTn0MIz4ClV67Im7aAKAlYJbPG
PvAHxE6SEsCNwR1BwcsxRFNTuqlxNJrc2PrzJ8qP4Wgib1T1Tjvk3HEwUc2J10DHpxB8caJEUPXW
LWNl20Jejxmg303KTWolqpRto9KIGVjC9gxAQBhpT9kA4yeOBju0UTNY+E7A822K91KMiw2f73dP
g8ck60kjydnYSxk4iKLKlKtnGFTGrOuBCcu2+bqBrf0NAtOBXAUfhK9REySn3eGXkuO+a0uEkdy2
Cgs4lmJ79xU+Mwn00tOyKaV1EgIQbjcKNrFXsXVeeuiU2IsRyR/P5ZFPKTZnA5JFfvBo/OKmlzfs
syy3OFLjnDUomBQbI8dworseLT7GLtYJtL/WhmOrqyRDNvkFpjUyQCHTn2FAJ8NDdURN1/VBwK6G
U7+vg11tZvXfTVnnrqdfeEWNYYwlXTumEDPvqWZjLwdCuyNtQwHUHo3SQnBd80+/TaLXrXKyopjm
ju/XnIQETl/e0QR9puDos29vYoy5KWe/Okh0lhPz0q0WM1JnrFW14pGq2MQHl1OL9MCtb3JLWmEC
y2jXd8/iko6Pfq8fdSdzSrGBb6fK9LQgsNmVHYL6z4UXX/od2YUU2e2aBs4wpldeG+Ph8yDrfFhT
+fcMTDEW2VDWl8trahpbuxylNjEEVAdr+xU8o1okfkuZGskXNKulfkf2BcBTuO0vMWOSWw6TVV/X
5Y5mN4lRSayu4Dngv2YoovRL3JG8LHbRZk94z/B6X1uOCZYqH/0wDa+BsCiu+amer1IJNiYRN6e+
HonC+cQ4GVbwEVzEIWKqp0MY7iNprx8yWpxJahLUXRfIWkhlGJFZ4J6znhD5rpJCikjsXk+60vJL
oKGb+89SmoAQiJGlEKDJdymaOivo1X08MBykD/Mu7oaXDaLQ0QKjDniZOE0iHaHTyGtD0cxamUCh
HKhUiPf7spvsRKwZSly8Gl3AZoyoROE00W5CE09bS9e+b7CpXlfC7TUoip/lQaEd8Z+DS/YouQjV
K2Xub/0orpx/tt4SS8AIvjKmsM6CGxwId1XKW7hTLrGBCzAeGrH9HukHArTuvE7YoEL7PJPkpyWE
HTlTWH7ZKmVnMXph5EJ5KdQZSLwYSV9IiE8J+YMI7cUqTLtts8xbVtxpH5Mjua9Ma8REY8OiE84H
qDviww5wACa/dKpGP4EYAwM9ES7PqCfjE8CbqrMtirL3MTeIIAUyfpNzxQwAinXF0t1kTn+xTYTx
PTo7WUyG7mEvA/TosBxlGOOlexLckx0frRwwZysmpb81l8yb2XuC30qOMRIbHZknrZPKPAb9rKNm
kXoxJQUVCtP09zCBqgRoNazFEcCjNgDdeMGeNlqK5z/Z9b87MJNqxbnAR/57wl6MZPk2VghU8hFw
rpAvXJXtx8esLQfDy64ORssdxMn+Xla45IrmBbcOvJ2Up70za8K3YLil/miRbo/vKSgxO6Dpk8KY
0N4sLoidqFp4lz5IK5GIRTZ4PhsVuQyOE3nOzWpRT2zVyFhVmREWtlR9HQxwC59GndiOD+t2DCnQ
8mxwLyVqGoS/msLBsLYKe2FsYLMGPJ6GG4+aVOz16Is0r7SNQTSzEWep+/BS+R/pnTx2x8LyUEis
vLj3u+Xdo7xvjmvhNTWcogG7CftparXmZ6X74FiyRkS/9rQHh71MTndBB8E8m2yvtLT6R1LmJQ0X
9OEWQI8igqwDEiOYTCirb0FaH32xx0UoAEscxFGyU8axYtr0ec17YvcZQLBtYbgGDmvN5Jf0GXEO
WF6+poHgMNmeqadOV7CARGrjvDC6cTMCMYBHOQxfgGaFzX9pW3rGxc0c/nl0ix9lgXID5xF3F1y4
45VZ0b3NiQJp9EvKDQfWJ9IkdATUFIpd8BZBUoePctoGwisVF+LWhrcZITHVekmChHtI0x/xj0ic
1Yp6TGoUy3Y+N+CEKZiIMThDFFZma2pgDZdrJ4Q6nCnwuFxHHhHP/XTfEfSe2yTmGbGkzZQW8x3T
xlH51HcV+mI8hvJipfB+n8mRp32Hr/D3Z2gxGiGo09sYlNwKepdH/wNP3kaVBo+7W7Bf1J4wK9Q1
S+f8y/EJ8HAg8+fvd7f/7ciJ0vrKzPrYoB8egEO2pFJ9dHzyJTZnc2tNJ/mfSSCGy2aGwBj3F3vq
xD0JlJddz2gvPv3ftexFC1JVt3iF/HmuFwy3C1QXbLbJd5rAliB+ISvGf/pITvzlPkoB83KvMyBW
3dEEK4afTEwMJuqwF0dQj8qc9RSHg3TK5Xb1bCS2PKLyJ4u5b2rVxewbOwBee5IK4eMuKzVTS/pP
8LQOwEdFnIYhy8xZhWJV+q5fX+pf2LlhnduQISff96iFaMMuaQW8uY0CXXpCincoSVmykRv09rP8
ZkJdpk1GnPs3rTsbIjNYRKTIJUI5KWpgIvw7hn0xHIPrffWEMGt4APHjfDmMxKgunhbdnxOc9wmg
9Uv4VEMGw2vymZc3OvwvQ2GEM54lkyCxw5rM7iSJduHxcxdcd0HWQI7ORB7UZefxLWeky/Fgtob9
kL6QdoqyGuelb50qMDoR8P2SWKBQ8Lf/N37Qwlpuxr9Jz26sjCbx66HxnG3Ntdehh8yIo09QxTra
Fqu9BpEX72ZtYKRJ34qHkF5mXEmYbL7zMJuKz3wh3A8Tr/nsCvCtxD09+dvGpjqA6yIRbsVFBRmw
dyjyveHjtTcI+CS2dob5VyLr3dCOV0d3KJuKhAJtifnwh2PMxDLyzfENU6buVUocYCc5TmeFA09Q
A6okygkigFbIB0UQIn9cmypH4qDBQ4RciV7Xq2TYBQLLOxflfukF274xpcbKgK0UwNLtw5AGbdl8
sQvSm1poaEqCGr8Ved+nWbxiVneLI6fbe16TklrnwrJmR7/In0VlP4YmH6D0Apwx9/a/5JxK7O5P
3BmH+/dB9Lb5pZ42RADeuxVjlNuLyxlYQQQVYvfjn1HUX1UOO7Cew+vjMNfkt/NJkRYOYmaLllCG
ATSXmPukogHVoYx8NfAOp6A7ZZ5+z82KHklwBh7xgICxhhtNeovuzibBPhySWFY5kBlyrHQ7Iv7d
EKwXxh+q/smNvdByF2h//9QZ2UTAIXHsRAVF2QIuVZEeKeH+7x9oNMRh8xs2xJJF8+chxhUgoVku
01SJFDQdomDKnl+8HjqpG7nfqfPVUHLNOIYHOzrM+v/OugNmI2S3yesVorAooajDn3lQi4fS6mPQ
NC4Ukla4PWhwaxcpcLCH6QVX+kpJWCORO9a0AJr0Z2WVI2/37HlomtugDysLHaCrRa6fnip/CdNV
5LIeO4qE75HCYVe/4ez9d8cr7GtmJ+6BYU7AQ+zPxpQxrPOwFhuggXgXrWP/GMrQu3BYD5l7l0dW
TM4SXSi7KHH0ksA1QEJhr4oz2eCXAVlck3KupdJ5i42TwJaUUJJQ0Joj0Z2CMK4s96dKWXMNbrbB
HysEOjS+uVJjDdHUUbCdvu1EPyNg+zjnFyGnKpln0XYZKZWrTU+OAaGrApmIl/6ENlXrFZ1CCUcr
EnHIsYHoWdDNASpnXWpMDPEHr8u4eEZy5JtSP5JZhMegYYoT44UjuJfUsIMRsTL1MV8VLWHKs2MF
lcEFu4hBZJn1tq/ldZj+N2oLTk4AAD/ruTeaB2aBkxgNuGsbM+2wbkS1WrqR8dlDFLz3OYEZKdK5
Q76Y3sU8OyvpsM+6MHGzantBJEOOKqzcMJD+Q6Bc5Vu48wtjX54tDr04P/qtWDenmnpWC7YdV3sH
8pMUjk46xaDEXm79qCJNg5yOPn5rPWprHPpEJjLOu2Lps9DDbHBamID6ZCQQ8jSEZGFkFNRM0LRJ
rmkGOx4vSZ1MoOK7qOnCYmPlVj47Qef/XDCtxZ3RwBavHe/9SsluOx0WotZl2RKpqets81i66+bv
83+r3rzsjT7HkgZxd+BSaNE1uCaruCocO2cZ4o3SnAQnhUbHn6gEojhaX3CfDXgfRaBQnnRnnl5z
6/fLErZODqJAt+KP5gV2MNQqLM5kimMLIUr82L3JwG2X3rJnqjxPwTWns3BPmX9q8y3a4/uXfSby
OqD/oT2fbrEbyAlEJK7SIV2IXnCTtiW4HPu/XxhIrf5khJrZa7mZ0OFvTH3T8NztoSsaOMPCuaoM
lS5pDPh6NjRhmpStF04RV/X453wtB+2ptoFL5ItzHN+9esVQwOXRPCKDzEuuGpJdDZ5/eeo7NFDX
kwJ+n6nrNlVhfQTnBAcdaMhNfZ05w64jIkncaVpY7PZBunPcNPoTrHq31MikHB5hUVw/tmmXH9IZ
hFJfXs1EPj9/gp9ULXZQ5RqsBu+FFaOXA6bIZR8bNd/Ncjo0f2FGujTwGYCNZ2EVqXLMJwkbI/iC
AK+xl3/Hnqh48pyetPJD29BOq6Gaa1LUFxB5Ik3JrD6fwPSwGevMPAiU52zH1nWD6SDVQgpS96s7
0rgYYrtcJWG15AjmkVriBt07YePw/vkL30LmB0THIS/6wTPw9zudf5tJIkFGZYZEMSY7GfSDuki/
iYwk/zpM+SRwBJgv//kHCJWuqHdiMJdPuLo6w5hf4VEsuNlm7VqRiayvXvF9s4ys9uGbZwD83Hd7
q8EM18Hp5sW3yNhPJug6T+vtWqffp62kdN+heZKJQGd3SlvmIjwIOoc9sOI+s9ZzAsR0Nmxq7dL7
XyBTbjemZb3TlvZ507tSgWPJnVJUKMVsFlGRZQigHXsUW4la3hmmjNcT18CQE/vEFkIDL8HiSgvF
GGMC48IQy4lYxKj9F+S/wRXPGI2cVw5IRQ84rwZ0ikmH8Pt6booq3ohUVky3sxUF4AFKiFQW9EAn
E1zvzBuAXUJS+Jx75wjEAQKlT6z9d3JNBge6Li0duwxo2WbyQliqN0cYjn51my7EoblzShhOZzFK
jL+Ur26mXHGjFfdc2FHR7GsPE14+1JoKiojmRlIxZqdXBqjL5vHaBUsOi9MaQxYuKaPJC5BNdAFo
moaj+/WxuXJQWIg100SeQcNvIQH2R7cdkREq1a8pKN4WeHN5q+fOsDvzMfS2v4R5et0jATh5v+zk
FrkjTUvhBFLvZbWnqhJ69P6yRc81UN6w6sP7HEsiKNVngQ7X/y83aRZ4CJ9F5dhku2Re+BloRRvU
w2REIA74sBEQ4+Bi0U6vV5Z8gvKb+uRqPgsEqkHJKoDBylzGHChUH4mAE0ZX0PcCfwqPAmMSDRqK
3CbNXRKj4JRNoLFtQHkAgkFp1ztLAFBHG6I8h66KRRh/7WYOaEHjhxNKLg/DLRiABCi0+v71MlGZ
itlBkL51pIRtblTisMEliI7LpxZoW9FdJ9NDDdsN1b2SBVCKNg+A1fblefKpgTU77UlwvGEWrknA
OQIWfEQt7mLnYVxDcNwtrsN3jl2MXIeExlex3IzJAo2Rhg2nsB56lr8pKlFzUHY/LIrR7sK/7kMT
5hIv1Y6HYCdvO0wBvHb4OAewB/APHJ7BPKt8D5pFV2Kx2KJqPgUp6XR18j4uSE+BqZycB/IiVrzY
wP1V3g/bv+eVm+Msw5nYA91Gj+lfKwaMfS5nCHVnEL5E024WAsp+kLXeMcggQ09okVMubI1fyHDk
w4e3jjrpfAL9Jhi4j3gSCn407ZAnS+57L5yXfkFaM+q2PwDRxxAa9uvT4FzJB4sUtZWHaRwEl8fq
0SYQHo4qJIiIQ+OUE/ArqqoojSIlyOtzd3qs+Ts20ftYUr4by2Fe1YlLDDTMcPJbf/zVCv6jo8RE
+Q8Dmk7xDV1fzSC1M3pB5fjR/OUZTZiPV8H3DQBAbYYDxW+pcEk5GDyeSXUvY1xByOQi2x86Fu90
36QjADuhrA3YroboERWn+kpGeMus7ViwhiM/wd+k1Yu0UX5zDgLuLjsDjZ/ifIyqVzYWYkxO+xAI
w8SJvgtgloYrncqH5hu0h4cCzeOB/e6HZmlvKzaRRuR0jm2GhzgFj8qQaafYcU2G9QOjOVYgN6O8
J4AYyg+Us9Vx9qDA8EF97ESCJ1Gaw0UuAqHNcnSzZTV8DHFKmuqJyitpOieuJGntzLVvhWAgUFR5
jlO1S6PPZgW5vGVt+25tsWrRn5dWSviqUPy8nBq7NMXmEQjT9oDF1h04I9yXQ0Lqctej7St8Do44
aR0xA9FEos/WM2NZTUlnesKSRIdPQV0MzEgI70h1Ce02LmeH+WV4SQ5I17qzKl25WissasOSzy4F
KbGa6UD3GIAAiPL6od62ZzsPGW4LeHUfKHRHL+/DarO+0U1u9G3TERzHMeUN6RNHfUkvYdiDJFsM
3wgnyTjp7Ngq0D84yLM6NtQyqHzb4PgkpWZYyPWZsmkUxIIDr+7FVG7MAIrUxc/RBDJUHbmIHx0O
OcYT6nX2NPe0e5I8sMzJhqAEtG3+NyMDutDdmzxtxvht4tLHjbWGjVNLu7oK9bncE7kBSwD22qXg
PfE2qeXg7wPrN2QrFz45rBoi/sDNA6tlgmG0aK6uPu4hkAxG2oEPI9OQ7SmHEuXLN2rTAXcRlPua
nOoHvgI7OTrugxwC0G1wc0Vv4m06QNaMuQkDsyUe5ICmd+jHPFk0sj5th1sfdG4QsAZDdVcIM4ED
EOWSw69ZaGEZzOeg1SE7Dm0+jjk8F1lgg+NEmA9OKM25/tAmWEmosGW+4I9OMzOohUsNrefgIVEX
jGd0BdJ9EugmVjaLTjyl8QL7TX2vG5AXjtpHtxRWn4DO/9/J/FvczXlaUGAKtqMAgo9QxWfPEXxg
kKZIIEt5a+VsXJPDUdS+0tDLhYOcd0jixoy2nLvsBLvVqylp3xyIiy/0C/WiX2QYClXm1H5yz7rx
o+GNOjwmqtNQ08ffh+jH6WF90I0LY/SjVninjK2Bakbju3z9LIYdpl2ihDUKrBb5VzIntuLaLXta
2iUUtdS0Gd4b84rCX4Gy7I8cVycz2Hq36MlMhlchbyGhVEkrwqlD9bhg9DLJTG/sgSgt3Q2rHqD/
qGmVrgUjqiZlPH5gTksZLP11tqPq1pF6oKsVi6LxKPmtHV+FYf68hwPH00oma6dfCW/3ua3iDwtO
5DiizYqhhjM8nQYrHFaKXQS4Dj4rT0wFk2MWIpk2lz7EqXkIGCinh3p+lWGDKQ5pjthNJuHkPdDc
HTrKOdoEy+SgTfXLC62FZk4Bo4x01db9XT1mDqEsiJgrT+66FB4VfMhJOULWvxJ57aw26UvEzBGw
E+MmXF6USAbYSbAG98x2JLs2GwwZQYr7YLDOVxpI8I6Uqlwct5c4vYnO61Yxd5z1SgSXdz1aW8oM
s0tL6cnCd9eAo+r3VbeOPyoSQPqp/KCd85owVbFhBM39wUenN318HhuE5Iuu4IcYlS9g/P1KmW1y
wR5ty5NU34UZHCRA7CiFXhXTbjehzHktMrpETUw4jLRdlrd8pwosp92+5loemr6h4sWfi769Gm+A
sD+F3VVPRCHcy2oI5yIIVrA/sZCTVWKSJEiZQfQjgh9HgMwrVYhnSmwRRiQT8uJ4SWvg7v3WJ+s6
fhVombfVTWb/FPRWJk68KLO4f7H87P6uWHRrYzpn0UsQ8WvQIX24UwWdlIjn0Aeu96jPVMKGw8NJ
4CB9u1nzdViFBerr3qlzHISxX5i/nmiGCUTsUQ9lS7PVnQ/Dwd/iUFUALiXvmSnnZeO5zFnnXxEx
I+smxVsQgBPpjMVF6Mu3fbA23+BnUVxBxTnOiRU3hEFnmp79JICYkomagyTDSkRPKuSDS2MOg9o0
aG2M9WD3yi5S5AvHSdkv+12kpsaNLUNfR+7n9RJPFztt9JoTysCdRTkQeRhCq/y/I7NjO/GELZxc
kJCLEtcPqQTy7+3nGVBssQ3KJviB4em2aUSBXs8C0B1ZW39NUf7NHMSNiEhIWsutpGQz4JJJvy9d
TamYBuvsDWzeI+RxEDX21zj5LqTrnCN2nW04sO0MlwKd/M84+KRs5jDPnmNVw/RI9CdZ7g3BdJDN
iGezlSPtyTpBgKdyEdPJcc5GqjlY2GaL9w2xvWub/GZUTfyOxHhy+TY69z2JeC5alENBU3boDvyf
k0eMFHnNXu7fnoqcxPs/UAOk16o77J7onME8eDBbDrWK1d1sZCFylQqp54l3w+KcmjuXpjGQs4Ho
G5UZpNy+J1zpKY0ls2o2wFhL9O1V7DV1FkP4W4UW7hw2cPHBTyOizlXLOCGJLBV8xEQjMBk4sm3f
bzZxnTNH/I5WHuSvzC0Hi2RqXdgCGijMM++CCoe9O02yPgdoT+b7/aaTZd4WZfCFeXDzJ7A2shGv
Z9+mRpR7Atwjaxz3GOKiB04sh6UJ23+2voIHWAAuFytvEpasPF25NSc31FPlJsSTxWEfpwrlwugC
rvOF4oJScy56UhT9q8qiFLeoIksL+CQsHrHnOkiKufAi5KO0yiCbNih0TTlNOfKr10Yeq4ghwVk/
z1SywhDhuZIWXKs7/vmfsI4RPklsZsUo9dqitSfjxcN/Ecwtz4hPO/JwBRB8pep4mxYqauG/d7NP
hJO6XG0SMUfqhoruDrjtv4ED03Zt92n/iMQijWWKcByU7Z2gYX2SB9iACScXZAvE8W/DM1cVpAuk
fhxI51utSRZTMJhUwODWESAUINndkZf5LaXgsIsTIk7DnSgx7QdqtGmiOWu1QopWmJjiByK8aait
sF1jrkwLX7dP3khKI6TROv+5WM0iNyVcHrnOnuD87+DY5UILeWqI6Ajh3+1hZAIEGfnqKrE0RQNl
m0LaWd98aR4PdMdqiTa1Z0FG8yW9j5aXN0VVt+S77Xdrs+4w0Q3yW4OzHx11luvEz3PZCJm97KOl
kHxsjSul8wQeTZAg9khLgOVkirDlaRJStKNjvXruNxQNJCXsRduTqIX2qhQiTw9FYfeC1H/M5ww0
SZOKCjjaX6J2lk13HAxTMaFijNug4BtzdKxSb8cbSaI/eYciGRI95BHHUP2XgNV/l1ynvA7QV/Fl
rFPsbEXPsWKgxtTrObIReyHX79DffGLxkUTjdZBXbJXMHTgGSQK2/WgZZ9gvsTetBNUx+oBIZ3vd
T+VmVZ65ZG9fSb1C7dmmAmi8Z6tGTS4Aqyjr+n2OBdIe5yAG76ULjxZpvjKpmQuGaPytjnd8F4iU
lqVDsqwzEBy5ADKTRoWPg4rleAB7TgJuBNzvwrafz5OAD+6HHYTdRsNrMNQ5rEwBZf9Xd5Sa7OeB
y4H4BVA9sTNpyHjn//ZNIvAL2vGz4qVbO39Otv0lzUUh0QsBGeQ8j3VHNMg24pRQTNVe/IjB31Y7
cxB9a4OQstnR0Zzm+kiaZUx4xUAZyuV6J/gv+TQYC3LUVekwOQQ73h+p4a7vRXL6dStZk+FEjwaD
ivlDvMVJMrxTjs6GsTkhIKsBlx8y/VVde3SnLG8YqwnBbvWu4n9azyKyhd6HP+Y5fQGetEkOqb/T
puC5OG76TAGDLSCrDjLZN9swgHWyzNNHCH0izFc9jwloUohf0OVZjI6qtlu9OHLxljHE5My2iGE4
j9VdfLaS+URfUfQrdepmaqCg3Ii8JL78JBDU9h0Ka7I24915FKuK/PRTldNJlrCI+U+lGosd1dd4
SUHZKoCAC2pCWLHEbK6guv258uUlJcoBJsn9M1ByuIn3nbh2lpHYnZcYgzxZwzZnB0GNsHMbX7kr
xKdXVY7g4CZNUXogVY7BVTCeeOoK3+KNIpdpeu9vhoCufqay8mi1YmuvfUUO2B7lCDBOmMuONukl
RczRPyiRDJaQZw5B0Mt6MpTUzCy8tKBCuxMJFUoyK9mv42O4qmVGfR60g+ghR4ljJSKzUuv6Typq
MwtFi9IzSVYFhl5DQu9jUB4f4jiY9tOAjbG+kcqTm93Y10uGTblh/mwxeqP5mSbm2NyklGNubIUJ
ZQRUsQcnXPrF5JfoAQPWt6Fbd+xJvaykfzLSbUQ7MSEh6m0dbDMU1D1qnlTbSUQa5SbuRqdd0xbz
SPYO8/0fSZCnskxkVt22PTrSthe9tas1eMADLR3W8tKjBD4nNsBmZUyi3VgAwIpAK7zzqsiMkUWP
3u71nnANMQmR8aszObLlYPGbh5UNV9TeuwnBZuUkzqBMX6ikVdSy8qORADjxXchSJojfdpHAtV2i
0K1lgZk1VbGla21XuztCFhkyR1VArn9NbKjl9VTFw6UYZDW4KXEwkmpzA6+En0JQ0z3Wj3FPKNTH
ySfRSmZL1BwVPtLq7t4GcYh3lU8+IfGSpgQstVK9a+5Zvodz7L8x9tsqR+CIe5BaIckqOYOfTikf
HsEaUkbh0EXdzHAvXXAabcIbkuRcrZfkrTGk7SxxUAUOR4ROu0ZhP50EhpeM07Tdq/mZWNUqoXLs
qyuh7rNpL+eb8maar80VOCr6M1VvY6JvH/twA/+GNCZI8CXHfCnlZX/j3FTSTyvd3jjfzLs/lFZo
pmOu7Mnc8VrB07D2BpMS+59eYQ9k/QxKb5rVmCeTpOK/LYvlrBFVEAPxShHdq+Dx1D6Ou4pgIoMO
DvAFiIkB5/TIbWmsyzxZcHtEqqdqEjVvP9VOVAHtbM6XOobSw3z+WzfqDL19LnFLJ8R9p9SxG/Vd
U/3VNCK0RbIKm9RdFI7uzHugf2l4Zc/4xUxMXcBWal75upG1tHwpkSdyhKuehZNfDLZoJb48XBe+
UTK7TkvQqGdgPV0N7LKzuIzktwQPnfy+3K7DTsfuRC5CcmQWhyUZ76KqgnvX33Ze5x3Sbj/FQsMm
sz7N1NoZIwSMi+9LpdcVi5FtWzB4cdLUti+SwNdPETarNETMbMg5pbcdc+vyhd+v9mO4pbk6gFpP
kehyEIU4wHBdt2JmJtIZaeGSEJV6zUUfvu1x1A79nKM0RxxYhspy4T3tdyws5SevF2EnhRTVkbs4
uR33hT520gg6VIWvZK0MPojB2gWlQY9JSzarSiwArc4forLRBXXHyQqSF/zPi513UfRTlB0+AN3e
DG9yXgBoKnVV1+PLZdy2eu9UAgAca2jtiXrH444EjbY2WGSrQ1rVvuLfSHamv6/A7hc40v4UHlDw
bhx+/NH+gCuuShOuEYLDMFOEBY+TppPPZWaY3KhXQtIEgXnhrILlQ88I435U6rVEUOpP4E50u7Jc
oG9dhFsKdi/6VrWdlqwiQ4ZhasEPSB1orhv/9QbzPN1PMOu2Gy+qzCOR79Rjmdf/tAJpzQE8EEP+
DnattL18QOjlS0Vok0tBfL0bVjO3F+cd5Sqsu9HtyZ1Al2jwEKXtMWwAtwCiUe1mDYrFamaM9z+l
nLGEnN+O5NFvH4BMumdWtcsJLJDA9KtTuNDPXoCliL7RJCP1PTmiIXBfjO+Ir0I5Bggkrw03dtxi
yhQbFhWzfge2jS3XNs00mN9ulflgZllPMTQPiXDdnYBGCfXK30hM++ipaajqaqT/3hsFgMfCeYyw
U2sTHRUoHqyNFABWvPrPlPmAtP4irohs+gG8HWz6a4CswYSND616E+/gkICkbfClywjzlk4ccPUG
T7fdeLuBwL6ZMKGKcaSmNd3eUCWu6DnHt6oPg8wkN3uM1WoJldyLRALAnU1MjMKyq8A73M/IOZxc
y26TBnJMmFswxRmQuTOQKxlOAWZnR7dvGg87o6BzULPZ5200dYUSyYS8LT4JP4ITabfjLf9LYiNg
QnvVbcaIbus/T74gz7Xd8D2bWpIgB+kUOPv2aGXPme4AOvc7Sl7Akh8koNzfHeJARG29KTrQxOVj
2T6oiQmhMVxBTFEENbE6mBs0ai4TwJe0SG10k1TbJHgOmbM+H5CfrjTZ/3X/y7ZmGqTc7jZ3Uu9n
+53zAQi5AKtRgSb5t1ZUmw4ZUUsyTXzQhrQbSvm3wk1ThCcrIHeZNi1OPHTYIQ2IDIP7xctw8DSY
AUQi0gbwsNyQXm6NS04ZRI1aVp6EG/FNXULc4lKUgXHgJS/uC4up5v+KBpWjIFoPcqKxWAXrNols
sYBQEacL/l3OSeSRF7P0aovvHxQNFoSDywvDtfUepbjyfGQS/lausqL2bUaVaAjDiukS3uj2dElb
nVNklANqlar3o01g1o+yB6bu6zc4IKiPQGn4NAF6y2v32ofoC1X35TIAopbHVT/P8aXr+7sB18GK
5DgxLDFRCp8ZtjfwTFqRZYXTcIC4PxVjeFxXtP1HbvB9KCBvch78x3liDa/f07sSX9CvgI5745fQ
Gaxqf0inBxY6Oeo2GEZd5I9WA4mRix7hoRpEMPnLmF+9enCmq3ctgtXYssAEpkGxfDahP6CD6Gmf
Saa4O0iCzXn/Ps0lymCX/0lR6jcwskcmnHz5cWXuz5P71GtYAwfLcJ4Z4dehgormVhatYELoTNvS
sWZwNUb0hoemT16+9anVOc1t/t08mG1en1HUNt2Zz9hqWNr2jz5lym8sgTAdINp747OOpkrSJjAK
bVMdW+6n+IEFn2P1CHUnY88ZgfjMpALc9wHEzLCZSX+wsFPQbvIf96fLfSm6pAWntcdPLgbs4GWu
uKQxhaqWnS0UKfqyEfcNLW+w8JxOd3d6ZiYXAqlaldp6sKFDrE3T8HVaFD6vapS4Rsfu7Peqtjgd
n9ByhEx3s5Z3csBCFDcgee/XhmJN3nLZbRdwiuhZj9pDM6shkPQ1KVrs7oC1g58Yal1mDRTBah86
M9W/T8zIqLSfybqJP1UOChYK4DiIKXGKnJllVnaAyqSpC2rWxCvDyDt5gVJ//Jb+3U8OdpSoLAA+
+YIz/zrdU4NIuHabUpo9WnYyBKyyda3/MxrIXbiOHrOTM0ZR4/2Vq7hIDnrILUDRDOu9hySOqxTu
yMGD1myFdyQ+AMqMYmGEmtG8YQwom20e+8MRhsefcGTKLDn63C8tPCxBXoOq6N/FVPGI7a8Rgb1b
AT7wcaoUeP50a6xtpxA1LlkMQ3E9ps5t0pVx84GawRgc2rmHIsNkNUY8AG9JvHEDAPAOL+qKk+wW
4j/lZoZBrIICuJd8y4oUtdzMhgkqv7AkLzTEHRdpMkIVDrePDErTl191KFNn09vpL7EY6laci6vY
nMKyp9diWmNV5R/y8yriwZpE2Tclmh/+7vWg+VAtFREhonmYtsbMKmeDGNa/HVFD/ES6aUBN/MBf
cYWdJt5E2ZUejtBrBiZb4yB+iqx94NA0lLUkalCxdkaI8an+5R6nQlXzYSnTQH7TLh5nvvfGpejR
1Y5nBXNu6e18bhkyW6wHQ0V+rKLjHvooeiAs9AcOr4Zn5eTEPqSmoa1NjYMRIDe+4w97s4MJgtqA
AyFnUR1UgHHfG+Tq5u3SHIr9BYc/nnPtLs4ykAAWMJQKgYiApBCzGY8KxRSXHaLm2omMYN2p/b2r
fYf7kgFOzn9+cjTu5FcEJmA4x0BRco2DmgO2k7RaGdTRn96ajmlVE9Y0Gl8ncLGuz90Mf3CzA/qi
ZUC3yZEuxXysj5dGEW8VQ1UEK4fJMMTZ2JgNzDUF1UncCRE0fX0iitjrGvz0/EdFIBr8fnweTvUN
eQS1CLekHmh/ZU0oY0+eyUeoj26JdUtiX4emmCz4g/OMjcVwo7iZyOZiAjiGE4S9RjgImCYzeTwh
BtqORDlCGdfqpYNLTnyF65+62DeDmlHodja/WO05no6Sv1zhIywOPnNchGNQG3nBB2hxlmTJg2P0
htPmneov24CrbkBPTDpjw0tENbwGXeHUN8jnhihwzg4Bhs7NGL5pAqEXBQfr/de881/zoFM4goaz
KsKgB7OSVrSPg0sByiy/m5YZFeKIt0dG/p298fCK32rDYFqizOPUxrGVFBaflujLzdER4fZZV0oV
XmLTcjEAQk0G5+fLQTi0T4Bttjil39+6IxSh2PFpPa0zFo3WbEyoLEQPgC7jjmDRfQRfYvLerL4s
zFTdpwtMEMqaJKDSE32ypq3pGNjKCFcjmXcMfEdMO3Tl1mL/I3KrmBNf2pOtNTD9WoE2XXr75yDX
B4MtlB5RRVIAg761l1DG2zLF8WXFTMY/HMV0L4GbjJscAlQuUBunvhhY+C9/rcH8XuXlZdhYaJ1U
6hAdn7JhmE43yZhXUj3nr7D6i9z1zJZjXmyOBV2qMwQcH4dMs91PZdEQ+fURUWCzhInLV3+HzEd+
wpzJBA3ATmjhmaX2xF7k2QwDm46zxvRXKlJjy/ZPcmWo/dxStVyxhLnNEfEHn98DRGuHoB+Y+hgw
nTWBI/OSrOzB/egsI6wGXIUAIGmZ50GxyF8A47biacLGozYFF7/M97X/9LC7P4B4ToZIKqNe8ate
uLs2E9xzLpz81CH61Vn4C1GwhVieJElYSxlxhzfnnX7uOvDarXLcBWJfL/inhGvHxl89MnPI8hgk
2hnIvjuuKbhnghoYA+Y6xwvaSBDKdwQI5HyUFSYYtmI+ZTQKNV29JZBsoMl4xrb/138apJOXuJ4K
UeGD4Z1k2eNqAfOAVM9htZrKbTqgyTrpY6aQOYMLNkQMpaR/FEg+Rpn2hNvZn5zBvhRPEjwNTK8E
5oOO1o6BZuI1SSacPKg+LBDuqKzOKJA9xUifaokpCBBWbwUZ5dxJxF1I+K18w8K3Yel1A4lGix5+
mVye3PovfpvlEpyjfWO7Dcgz+LKiJIovQz6FbiLOJgKdVUClcCwkaxst8xozolBRJtRJkMM2K0/7
+oG5i0iSu7mXot/mGkzXSCOU8e8GvDjDl966MVYMW3rGqNAIGQouBLahJf20Tej5QY/SoN2ED83l
6l9neqpCRMtW4WhOhOL5tTZmPpJfYEwoB/Au9TalRek2Q0InTIeq6jJPKa1oeoVdYj4dp7PEUlCK
8j+ignzWaCXLVtUaGxLLIZSab8WGC3NnB5QTIDTiSR8QkZle889nwEwlTQiet+2+VPDNVfy7LmvJ
maSBpQDMGz/kLko0TZlw2wYgoW8XMr9qvyHv61u93fjaG2IKuWT+okrZYSq5y4E4aDE/VeLr3ySH
5yF5X90UZWS0mTrm19pVf8jYpMdYPSpNBlpP6QAAW1bw2xRqqS2leq5qIIGogb4RpkPE1ONz0yMV
IoGZCAis0+dQ0XGad0C3oY/wTUusDygViuw8qmWtThtxTEL+HpbswXs3wIJS0rr/Ed4t/oWKp1mG
wFgkwDuN9t03dhMIYslkU6NqjT1llMzr5isS6VE/EAial/GZxtNbJil2N6kKmJsEOs9o7eokGvrJ
eMgd8B4C+0lXBjyOOiJGPz2B0OF+O3TZDDmyfivK1s8Ch0UfQG5k8iNF0uVl9Ao1vLadpI8G8f1B
8AKli8kZwsH4+rcOp8RcH99CYTtIffr1ubExewBd76iBkkTQB/ALNCGIl0MmRRZ3RA0Vf8plLBSJ
G8PN/EnHR72PvNn24FrJ/yAWgVDpZqdrzzQSJsnZrfPoESwwPVyUwwiPs5u28BWbmuQ3SNh5rrqc
NfM+iapCi6m7+3W0CAHT6pCK/BzZVFkLwq5RlbtZUnrAt8Xp1IErGCOUre5ltjXZbokFvzawCFC4
Z6zMPGbV3/mylR375o3ElRmZtNrw2baVDsZHUANM3vtP4WXyYVfdbtpc82SdE8Ux574+2GgdSrkd
6R1Zo5eyg61g9ezAoO6YgvprZeei9pg3pgzZYfMLJrTiGPbH6JvEeYus1tZSg6MMezyNirVodDjG
M/mQXeIIeUKQhq60mSPXMjJEB1wZWK91ptuE4ADcl+nao14u7NxYTOF2DsU1/zqpYxdnpbqb/sqW
e4NJUPQUAuL2jSS+7Vk1oDOmikl2klZKvcgDdzihxV1TxDp2k63b+Bwk5W5WN5L5CdFY0BouYwFP
KA29mS5JMDG7EimSNtS0S+L4Gsd0hW+DSLTOJ25TQdujhgnzO3/eqxmNWZaTO1duub9rcqQ9NMmf
PuDBoebTKhvil+aAV8YkkeHCigMF9GtVqL2TBVOPnpAtQvqW+w6fylNYM6RJrZIttnC7bCxh9NH1
W2epOs4C4TGv2esYbW9QjsD5xWMOB0VRh43KYeZ2Xyj+ERmgGhPmhLo0i1TYl5kKgoQxM8qnGxjI
LxnlNUYs8/NlGE7L8q3P1n5ikROe4HcOSJeZAtRgvgBgmxhQw4TaovGRq++R12O2IoGrpKCJaMUc
Sj6yUzvL8jlbR+LrEKJpdKlAa/5ysfPE0MwbsV1iZptd/jFJ8KFRXVgMLjfmhzS29Sq0H1slJfxQ
QXuAup1J2LeRr9Y6lyYW7liTp5W1jsKbQoDA93ffPEPVmdoQUiHdcCJRlJYCLEiuYTkWN21JEjnj
QtS/DlaQfDHf8tFWoLtZCE24FZBIFuir1fV5++hKRZYtmP0c2z5A5qgh6jcY4xX81jUL1j5UaNoL
QPx45aJYA2m6CFAyRY+6W1FhoB86APSrw322CkDm9FJa6vNAv++esFly63LR+p4A2F6QTzvpAx82
6einfE34p0hGZLSfodPElRLBErWeVS1TkPLwSdz2Ko/c3gAxbKFbrhNNWeqMYgKpzIvS3k3/TFKZ
q5oyO0zfP0+XHyAwAns5knebV1GP/iIhHetTVQ5I3e51p5+Prib1RejqJnY1OjZXKt3kvQ/N5chP
gM2HuunzdDDEB7VXBCyLVrcjjUaO/3JBBpSIgnDt/0n8lE+IDpXeCB4jjdyEHY2hl36uddzLuMI2
ieenIwiiPbg/ZY7D5Rs3t0z8Hkh92sQYgCGaMfaVy1r/mc3BnyToWR38Kwi/tIyvqBiVm+ac5mTZ
KAO5uNoGVZ+M9KnZ1vWxfhfhZducLTCRHcATyagF75OP1OcaLPi5V0cAKcLJO3kDJM81xOh0y/qN
qTC4E64kRgN6jjfZaOdG/72yCX/L7sy0DYpwnODV6pUvTLyIbZ1SX+mxZVZ9KwEIClh6PBHJE9+Y
YTkvhgQeQavfqpwLNnGF5Ed0XTpfC1YnGMSS5ULpeHmwjhCEC+xKPXd/hej9cPLbZiMy6y5Rezn5
egNVQVeuX8N2PFShD1rMKKFk/PgQEJdf5pDNo1DzZUEp5uTyCgX/xXmU9xs3iNEDO4KZ8cPH9ECd
vF0/5S1GDDFQyX0SY7ChDJ19l1fxa3JjMvSjSkdOTsYGCHqeR26lQOMGcdFuGfJv/zuzWxES+5/J
XVlNmwztyDueKn7fQIdk6UQTfgqOB3KqLawlt7OFCayzbgHkMPLKckdRWq5Q64gyYWd8eHIRcu/i
ZpWrbgz4d5P0MLx5wlh0tb8/Ug9ErWb63aQpwCV+2xerAM+bz5Qtf71K2vAXmpEqMn4+qWbUD1nb
oXxaO99vSZx5bS5YsE01af8Nmo1Goh4Az2oDVE7dFYfjOdK/sDUc1ADci9XjvzbIlzQELmJr/XDe
eWBwy6L6hqDMuj6Ta0WEtZI0VeRXR3G4BpKuQC8Fa1Ug0sn9hktiZcGVQ0OGsQ2Z/7PncnWmDnk3
P348Ii8TAl1Q9+dcyzw8QzQj7YO9k6yHV55jGWDD+4+vHhZcOpiV4Bhhttjbp5N9YXZoK9u74AtH
Cxo9nzyqbxhWlkmDhmufNWps6HG2j8MdjluX9HK9cPGDz9NEg8sd6jG5E5pcKgNYSa+O5uEJt2+K
/9m7bkZIbYiAxWTmIqKVir3fzMKcsba1vZjxzHF0rYyFCSA8269JluxzfucBP5vFmNI2ejhbJCLu
6vn5CBVHB/Ysq3NOp4ivNFAyFp4lCwWykbO3El6bjbeFtUzyJ+U9LR8Ljlx0LTcrCAvmLJiWmOXQ
0LOoEYIwGmBHdDTXgPZ9cY31a4HTWmEQfHXZ2fMVMfJbbGfXKpK5xHfWE+LShnWShnqNeURzmaSR
MsGc6UNNd8LnmvVF4/TXRV3O+ntW4UXh+UFizKeDCwTNaHZTvdQ2yL83DyOpbfSyd4gpZ8K+9ZkO
2hMiktsxkuJf7u/+wFsLhLpdAgUkQGVoJJ+7qR6BN9Qe9T2E1LdW7jY76+nS9vlEU7RNJdGinRUr
Ks3V+2bjVBf6aG6d7UrPHKfm6+AjSSDSnIp/5y8Ew5zYxTvtTLSOD3QnkiemUYAjCVhaYqXck0G7
2KtiiZO0yOvGgE83dqHKQKuUuSY6MSLoDtCAlfofOy8pLi+rBxsp8b7fqddxkWnRg2W05J0L1wQ8
yo9ufBGXm+GgMWhlmnkAphWwNycj6qcaLPzobPFS6MZNx5eFmGKuG8c4NzPY3d92Y6oM22GU/QhJ
wqn14QUjkMqFvfUpIl8OC2qurd2nacHjnU2fMpSr2VKFidab24t11pDfV99s0pz4cywy9n0rNw9F
yrp59W5X4xs1/HxWw1Kq3SEGnBzO6qoMvoxN0bT8r4grn1BfjnJq1+3b87VbX0MizxMsFe9uX0ez
5MZ8lvqVYF4rhWSSm7YWibS+j+fQn8KcEU7eApK756dnssZ2/7iHjTOwogQlS2crDb8QFcfHsbtf
VAnzeEyhwujHIweVaYuDqmfHQBWTu96Vqs+OA5xM6oDMAInOzCnL7KEU/duM+7PqjfhEpktIBm0P
eJ3ozqxIb9lD6R9wPazWIltGsdo9O3GxSSw8bSzp+0I1HY6C/nV1gK02TZuLWD1NHat+WFyngf2J
S+yraScVcJE2NNGZ7jNFKJkQdv1uUhXYzAoaKtSFGZQtgoaDjrHATCWWs3RX5hjMgP1WgCZT5eCT
vqKe8V2MmmVzI2JQcB/GoHJIdUAPlRuJcP5G4+5QJVzXM99z4XaJDmZK6Z1+BshBW+xTlET8Bt6K
IhlcWkdgegd21D6z+vWVBJ1HhCpzmxTkqG3l/iLOt9sBEHfzRwQQM+lB8I2EdwEgYiKlsK7lvmRY
L3sB27awhabM3YmjBbWK+CxhOs49Z4SutoGOGdVO9udVa0ay1xrfshs6DzQYaCIxqfqDKiHlIAzw
UGGCn+3s9XVKVknQMmCIC0MjeeD1WjkPzXwbYDSsPna55cD+6c9PvC5BmXzdpNrvP9tcyV81ObqS
9ynwAXlXnC8WFeZ5n0LA5V2JvfY61bUzC28CwvL7GqWb98qJKpTrn3gbUlkoDdLvTAdmpL+Ceabe
Ulhs46dmp1FSWWtmivw3hzTwx3ULVwpYEgr3c1wzn/RWm3OFbFrAXJEBUmF90hl+96EHL4WmDG5E
Kh9ROCcQqr1m9jdnAhYz75bo+1Fgp+e4jmfWZsvEulxSIEIH4OBkN0T1eCdpMgMkQhPh/l0rFWGS
G+YtvTLI3S3joC28QCtz1roZRMm9iNk5TutQNAyrjqyu72jEGMeoJzwQ20dfXEvWfRRX9x4eM1MJ
mRVpAK8BCYcShAx5usWrqp0mtWdkZ6jZKE6vjVCOBCesYNmn6sxgwYgbqwUUoFX9Va2Z4a9lC9j9
J8CtkeKIY+BWeKZeRe3LXgF1pzZ0eu4XetS85yP5R9KR+UWXo/m2FEyMDPaQ/6yWAdsCS7zGvZBO
4AGFBr6oyYL3aryfyla814PkPPOOD7+kvC0+4tlUfILR6oLezuXFA6EN1YnFZ8MiO+10PbUbOi8S
JIgkiP23IQRTm+HbwxGPy+8pvkGyYNLfABSu+PHN76NM7R7fusxOkVvHY/ZYfMd1k5fb2AL+1ju4
CduDZULJ7rWdMayOL3hWEXuW7H2n/My6lNXFfzvGiwsGOKcLfqwoJXfYtzV3LlQh0om63mdCTLhj
3tZR05uSlbQdp8aQsinyQLiEOsvlMMbjWWkGXML2u0eFyPdJHIhthqO/HfbNaVRwpcr57UlXD8mW
s579MyNJ4ZHqGuUGFi3JUldHtyQA3MAe3lAHsAhFV4wAqyU7nzCqLhWvnj2mTLqm71JQAbYdLxc+
o9ESpFrEHu8TIfmpP+R8cYwlowBrbhVq5odEF37IsGxnlpVD+0uJwlolu8km/CozZe/UnVBbhtWw
dX80fnzBjmANjQ89aSwhAsZZzpuhCydc6Cb/KYEAMW7X1O3D7Z5rpKVz1MhOVHoqVKV82DJc1WkA
Uyb3hKvSXXBxHk6t8LGUWNT606bZbH4BTcTc5e+7shAklB7eQR4PfLNc/qlsod/1noLHH7T01yhb
s1Uj1xixcy+a5mlO7fs6SMVuj4H7JwEQBHrC8HRrUdQV6+wOIl+0hXCJ+9w0mDl8lsvTbZe3zIdO
KP8MBWYp5xee8pybdDBOaN8oXzjRAYsCHR1Elk0yc83RojbHs0l8H7bRI3NnoPcSQxokriA1s1Q/
Kg3XN2x8lafiDdgY7mtsjjvzpucEG+2IA9rlchDF4j+93ZXL2HnjwC+Kf0FlncCxCGljwjsxyfsH
H4EmHc4d9yZy325xjG9i8fPjU0TELt5uhuOgu/WYtggDc9HKE+4UiOR1i0iPs7+a5ZlZ5PikI3Wc
P7jK+1zEW206n5Vd8ozrhGOmnIY3sQ5PpYuAc+tVU0bns69Mr6YP94E1zLhGfg95XxC+Nma9DIQI
AA9qTZvdQdGAcKo2hnbM02rzmtocKuceUM/4k84/sc8QA5Iaam8S0eesFlFMLX0RzVM73l3UskqC
45cRTYACTp8NVxciEh3HODYmHSpgEdzfNBzxe09OnRVbWrOzWLi6AaxNbzp/yv1e7pnlEz61tPiP
RmejIm73nSzu5WCcztN4rNrJr7WSRtKpzrhHASRajvG+M23kR42+TkMGF8nmq56g2zDuMXljORkR
WtzoiIlGPRGEgeRVrDwt7tOO2u9MbOZ4hJAZA1KX+cmmWvw2Ly9bTOJKy/rkvW4lMD44IOQm59ZH
SMfEu2boJK8cJUodaZl52BAcrsFJbUhQfVjIwK2qpFZlM14AsWoVdysmo0VyMbTKyyaUGBVC6yae
nrkUzI14uXhdEscJ5UnM+l0G2VokcTFWEFcZzWXFxKdqaJjspbjH95mM6CrsY9hyuXDixPwLK4cM
urOAMlZ0m7Vy8rdduEZtYgd7ltEPlWwjQiOOAwzxEWDMWbdPLpfwP+THeYIJi2ioLm5/aju8Gck3
1uuzTGOBD626FUU8muhf6ROw8zzNmCg/0XXi9IH45UuGo3Vz8CPHT1jJiLBtLdQ2DzkPJau3X+iX
mizFOSfT56fKmD43RLXOVoWky9J738Y+5jNGWtV+Y4qKhI8TkKOKANHmp4fiH/UCq39HYBmSzZPh
TT56ld8QP8p9zr0y/W7qHmJl2WVQuyDugB5Fc/CgtUdMegrkWKhEzBeEQIr/bTw1asB0sf4ndZFW
mGhxGXBkSLjrhyKkzC8WE1+kUXTkjfATr9aZkKhlUlv9dIlJam9xruddDrhgRg23bqt+KViYt0Lu
xWHjub2KDGojn4Sw5Z+MMTlJYHuLm3XGMTqhaC9Pr4UXMPgdca01pCrYJiQ8WSBwz9gR9CfpNDp+
+bE9fTHuLgwZacH/82ixKaKEipXHgNX4B43TW+fP0p0ybofPSuO1PmcqHGsUg6JscSy2GGy/7xcJ
uM23Hbd9JJL5sSWy9lV+fM7uqnnjWhCvlWfb7j4bbKfBt3iILkt211dm/t7Cx8D7xFtULZSgUacV
G5TXE7cbo3wiYL78SBG+i/iW8xnxC0NXtCo/c4Yz5Xw9QwjLCUTa22rJS+Hwk3hSTql3OAr089uo
o9c1OqO/U8mM90NGac32flSbGUhwcaY7YBA/RJa/pfbBPJiqLdOzIfjR/xgs28rXfnBOE1+fwZxR
UGrbSIIsYi8qPT5P9ictceZh+tQGH2NdaF6ITFplLMv1kg7+96TZrhE1XX9mqV4HDfVr37vxrEl8
HcPjeZ85MBnIO/v0K0sgukIAS+Ed6sNVSKR39t/Q7S379ppNodZ3Yl1rDe665+AhitZ3d6GooZmP
j4ZRovuLGw5od7OiEXLPFBEWn/RPPHO7lGmvVMffvvf4fdqR+AuWw0aM87qA0JO89DorkUcSpTNb
JkJMUVzEh9IB0pYrjIIa8ND4PV3a+DLmvNT4XS4JQxZDbIrTHyY3Wwcayv0kyDbsVf447347hltC
+g/KHDP0tmAOi8w0uF2ElkIktGoNBO7ZriMST9lecSRilLA+ptPOgOgWtfs7nwDnPt0jx8jkre2K
UCNwTFoZL78dr1N5jGDJ2vU6JFjWTpOY4Z2KS7D80hPEz2RxDxSx84ksiJf5wGI5fyZD4YKZjB7d
GBWdES0EvrebNxHMm9BsH9MDEPDk7fuYInAFrriKAsSPfdKFJWKLTIMA+8ERW/cz3EkTOSTgH5dR
zy6poaYYyHIWoEPedtYMPI5saQFwandT047xOYAA4o1Pu918h6ruZDjvnScq6+r1s4fBojDZlu/v
Jo7oJpXUuhhtNKqAbSaFGSADWmu78aFssv0amq4WoieE8AHkDLI2xPQDA8GeQqRdw9B/e6cuqQcJ
u44IXs+5qA0KLhq7vwZElUANRZNhSmdxjxDlVRQmgg4zO5Q8ji32gq2+b039en637ycOao6yDh/i
IA5Rmql7fQRqSgTfqN5tQ+aw1hzA2+282q1A7RMgwS4cgCOlIp20WdGhFVXiSZkqSzTjnqWwBdnW
1he3ug59TjlhtesRWyy05oGxkPoD1+CvRTHlBKVKFuaFNb+c623dyORQNk5LsaE0SRLmRAFf8MYM
ysqOiQQprRzIWREKYGUYzBIkwT7WGRiP13zyDUzSMMx9r3gU0knpQ1nBE9QvgZpYlimPwWjZgkmC
JQjp/RIvdXxkCdfay8H1+FvdSZJYkSrKhw/p03qkm9kjUc3qPfSH28xi3XtBoUVgdix/sG4K3t8E
fGGtPL5OtxIC9ZVupagcNz5RsWh9xNI02Huj8Hayud+dUv42gdZ60wR1/R8yizcjV5zwpsRBe6Z0
t2iv3SDpMu0BMoFpfP1e7SxTJOJQ+3zB0GMb1ncPY1fjIv/Qa25ETvmNfwYXJwlaoUc8ZOQGr3Ky
JFu61J/mKFADyuvuxuhs9JHjPG/ytE1K9lz0rpzLvGeTwT5ydHzytv4YWxD/nyDhB6/ezZKsdogZ
BF4ZuCyzes+0fNWfvGVqcFwBCGwvkZ2i4G7VKMYqOz1lzsPFIJ6lUBki8mBsCx3VIOW0UmpjmCiu
aspYE0EZpPX043bWvjIiT71rQpV9lR0LfZrkmL1NA77VMolEv1tYvo75BUEaN/ge/9SNGIO2eh/w
KJ14C0uD3f53c/bQxc9vAL6yjykWWXkDKaRhzwAgZk7nE6X0zGNfdBUWF3IQYUGbTPUPKn7KG7eu
kl44N7Hdaw0ELFdGiUceYGSGzM3z8xgg6HPOpUuDvEzo3OymAuRzvq2m59a8EmLDhtfY3FuKLY/d
n/r7adQHFdVBFocYp4hg3yfCnE0aTGJuYgdm/4LVY3qgH52LRU/8F6uQdQBeZgg4Tu5c9jVuco6Y
qh+8+Wy18JsUItE1zvlQMOHYQ0i3AFFUWfg4MD+wPK83i75qI6dULSoBbThXg0pPWDF/5oCYq7m1
mzT/53y36/Xbhedv1zMx6gTHCDkbKN6EonvzMMS52Vmq6C9h7Asc4re9Yc0LoQ27qLUQR7mjELrA
5OBEwhpK2RBcks55PZLP4n0fzzbuFccYUlUuZokk29nKXjAYstNXsr3MpFvPd2uPOsa0ov9wcNe/
5QQpkPKqfKwi7ej/81I+MPufrewhF6G9OEPSsw0Snelqt7Y54l1CleiF5lLxJ73N+boG5bOKMiV1
xn9MJ1GmDX6Gk68/6FBIdfSC5UvPC6GIwCk9tb4EtToy1VSw9zK2ELEmMXgrWDUn8RIZzG58DNgW
JwY/he0I2Wg2IOv+FeZ7mJMOFpdDhp8PRnTX7mu1bzVpFqdk+X6EjrBSBZZjBE2SFYgGZxIvGmmO
wGVry40j9uOZYQLLflqAHQbrQ8llIDJ9ro4KgE3eDb4QxYwWl6D0A26h0C5cijjJP7WhvzFwEKZh
wl//z6v7xH2HO0pfwI1EGhkHG24kGBaMuwqViOvIoQHLQdVN9fPP/I2LLx7qla6/5DQfykrS2hm9
FiwrgGyYYP5VHTI5cEqsKOqNQrsxGz+xzrkazt2X2OoZAk0SYME/FgORV9XdRdIqOfSLZ/UY1bxq
nl32w3lXywpx5XWv5P3WfsvVU0gINfq4Mu80cFwxNOomirXpIQzn8tvEQSJ+IPQdDOuVN/KLY1hX
McxQG0jcbNcPfWM7JLOu0Pzwkhs3Gg8WIGfCxfzR6iUCs2C8rkjk3Re33oOs98CGFFDkr2dcIxwq
IHa+ddvqfdrdZ4757s1Pwu/RiCyWBCcYlZLab7NlSzxqkG15a8Del9KbhxOiF74I7dve5myHSSbc
nOBL4ZqhbO5QgQ943wHWQDiNvtvvmTqpIaSUNhgpV4MJsmV+epNzTRIuZmZc81XhpLVj226d6tWC
qkVdfa81Z0TJCkeazJFteFnMEZDapIa3imVk3OPZ4q2bjCypAyO7TSdhkT4FtdX92VBFMA8LY1cN
hqybvSKVh1aOjxS2ufoMdgu8edogcOTII+YcNbVo6MwoT9rhq8TqyqSWLJsgIbZzczfMHMv/juHy
Ki7mZyHeC2eBA7sPSvWqv4G+hT/4Khre2CirzF2wHguWrTweJ3LdJfJfWEqbec6ztr5rikjFTIG1
v/Xb6vIlKKAbwXvdLeBEJjFnVFHWrcdWafbEo+c0jyAVgKtiV0JmMNBxM8saT2s+Goy5dABxek2L
a5Nqs8W1zBKB0mEUQH2Z7xb1zb5l1Eo2vB1dH5Jnz8jTp9TuFeulfHAlJwo31AqoED0mkIUXu7HX
vUuEGJ+m2pj0vEuWadld/8sGhoeKhuoHVgSTurh93WGs50M6jkUSoEH1pFglGkyBWCAb+V0zbPBY
jePS84f5VQWbJfCa9i79nvAX7hEtuVsvD/Pr0hRmIK7cCvFQS/365/hJLj/1HoAUPAO6VW1Kr2c6
6vS3G5ZiRn4xOHfUmQgBdnYsTyA5qB3K8VoUqbpe7MZSNbI8WVA8vDoAi67ziGAkK+mJTrv8LI54
bYjaCfe/scURliCFBHM3yS4bFSlr5IljS86bOoO136HJ/Y/aoaLYT9xnOaKcyjgz5n6GFBz1qsdF
ALv8RXIwrY5/JWxDjV+PuLMBipsYVAuZfq+r3fSaqgP8dgv2IYTOlu0epLQPA3l/ffhcvd0PnvEd
uQ7OlBuZh7OSEJjqTUT7XkNWHhmfiBX0y27oKfpf3G0p6Qx4a+lX9baTkUgTqTFJgginntzAu6TO
Zs75IyEh7n/CrXau/LQsB7wLlN5h21XPFbmqFaafRhjp+8o7HtqmJO176C08IKKsUPtMZtEArHWv
TEXtQzDsRQnaW8COG8kd1BircZVN9ssDmrzwg7ZekbmSRxSAulqj58YhsraX97+m3KckPAurpyYd
kZELtmsU2UL+WlDAZ+Yc/rYYlEgIKPJmEgaEfgKpzv3SM1JNLfUA67HmJS8RvzP+Sa+XrSe/I5Tj
ZBQ/Oqukuk3trcZ+CQPE3/Da0sGAeaZ/qshh4F76meQHPHIGq0d/qkxgxov3SLBun6jVDZRvaP9U
Thmyp/7Y3bNdLMfcZcb0ynBCXcVg3UfYtVy2BykW/Mqdt6nPOue8xHTwbbxRrlM9hLTzkQPIcBZc
TC6acU76KzlGhvSNWyM1jA8eH8FWULDe7EM7e5n4qs8vKErZRN/4r42TCEL+e5BUornEWH+Y0TGW
+LGO4Dn0FSLpKHi0AAQJJ3hCx1su/0GFHNyhvfHJf+s7H+JFpaFlDB8ybaD6OnDtB7fZqRvaeW6j
RpV5vo1v6mQR3aBL6i0UuNLCI47A2zWP9hfkmKqejsu9k+XMKDaveKK3yGyRhohFWhnapSVNDLbS
nhwYI+laTzApv3xovBaey929tMSeGMtRX8Jt9CyreuSOqG+J8XbeHUcqPQZooOP3KBBK+u0keNcN
n5p385UZBj/9XuzBIkwtCteyq+FHpSvxaIaAMB30Nx63j/gs7LwDUaFwMUPv4DHEX0ovYfxaN6lg
M9vRxktFDEWm6Pu7Go6nP35r8HoNxkXf+rM3uSUIzNGfsczslTh+q1mkphMFmzUyjWHaOajogXWa
VFOGNcsFOX+AuuM/HIEeBt05oVlzMOeUkPacaFmM/lH/5h178BDDQfIMHEvLXiXPIxDY50kOqL6O
aKWx+0TYFZHjIs9fDnTAQxOlw5Y5OpKvzUQDZBxs9MHaB/mE7Ken8vhuqEoiGIG6JhTLTA4MYL+Q
vvs8Nk3uoyoM0xcTE3Oq7Xfy4Za00uo/MlOlBMrzEy2WiGLxxgyKO4eA5Id8kjHcU98G0ubogApm
hfrHxDNOHipuKcbMd0riQ5MlUKnjUS/z6QPvNA8sQ8cUqm680CwYGSn81AYEpS5K1/ihqfBSFMAs
7TFvVBR/qK8N27feFvGhz2btlZYyTIxSR8NdHghQ3/hFT/7ZIAwCUou1ROk+DBjCFQHd0gUwlpRu
BdNB2nBUxszLEH3l+J1c3bOtI6V/ZYdQ5f/SnEdrJLoAAhQq19fWfFc3UJI0bMqh6j4ctWVEPbwk
PN/iq+GVlMaKqIwfjeJ3I7/TNj35z/KeZR2oSuV6qJHBxRgED05KYiCGJqVuyRhL7UDKifFJNQ4I
Ozt9CfTMVVdeFpeG6vbHzTNW3DPTgRCRr0U3LB4kZRn9HHpIAiyGn0Hzurtwv0TlTVbVR/7kPSTc
ZI10Fr1zxbIbnK6CG2pVbPe9tzlul3OBfZ1BKNNnbUaJq8g3gjyaokzN3TR5V36Ceh+KtiviOrIf
LUFr5+qrkzNsc3JlL60niMRzVjXYcDqot5SAsnCoAqmh9mTj6tAeQO9U6P6iuf3dEgVmj1FSvPWk
Qi7HSz2zRN6cC0TkgKm6NTKOaRU0zXJMncECcR4yf1UIjJFePtVkkh24VLOH5PL9+mI4JYTENTrO
oIUj8X8ZzSXjLyL61NkkdWqZlktFD5kM32JMsPwbL61DW8qRORVihZ4HQ52z1Lm/IibUulk/DPoY
MG7yBjk1LjAKPz+efmWi7YYxh1xCxez5U1UvEPee1DGkKhyog9qK0BxvbcQVfuS91D62pPnubQgu
W4HcUggYiHvgXs1uG+XqN+DcLsanUbW2R3d5z425DjbqYut3He8O9AARlclQRvDtWlMM8jTXhT0K
IZlJW3iybRrcGbSNUin4RRMkNFJ0ReySJIMUWonn3+9f3nXpLpKMC1o3wE8aosBq3juwvgr1JIX2
YlpnvMw8ZeBVTBWEa7wJgz/n9QtrFFCXMgTafDNy7LGWOBgiDMkLhE/zUzCJ/ApfilLpOzKfYj3v
616onnvQzDlyBz1cOc/4oZ0Fzu+OXOEDU3fHlqL6k7PDtRJrD9vDiO/SdixxDBLU2LylYKfcXpNM
LwhasJQ9T2uYN0JfweOSP3q1p8GMwG8QXh9xIbptFZD1FEnZBir8Llt4fvSIeFl9ce0R9vGOgRrH
hsZcfnvveFmK4XtTNhwG12YRPr4VLiuh33OLldtEy3/F5VezhIK+o7ifIVNIlWskoM7NXtz+BX7O
9ElK+kiU8xLeNWftQah/L+m1kgKeOcwD2Qka0L/EATqfalPQmA9IwSeCD//FovE3FDUOxqcNoXzx
iCQ28ZPbB8o96MwWvVg7HZaSzAPy3cP8LRnyrg6hOPI8wcc+sySiBiJ/hwMc5M/fXYEodRfRB/0q
VCa8TU1uWdeUaCwGYE/MucI6h+xFOj/tQG6MgBzIQl+nX1Q/PR7bi908QHiKhURLXe1s7np9RRHg
8SP+G3Fl+YXjkLwGp+0sJx5iTVjQ5yK/0NcOVYmZ7MzuFMpgHMVSt3bDyq1sCiiLauHkmChbh4W8
00sGnHb2bF6GYD4Ja6LetYxyImqdzR9JoGNgoQtttDc7w1O6+W9rzPIjdqKSYjGfegxRQ1USE/78
xp9Jp1pXUo6fbMhTYYMNOq0ssJPlEpMJAaMCmK6q1W0TVIB2FEnNHdIVxOqGLEsagtFQQkz8QVlQ
RBXiqesUJtJqCkBGkjFqRgDITfO5G7GfgOnXXtvF1Xc/CdYtD6SGcxs+lLNiYb0ezOm23Fy7tWfL
3NKTk9MIcWUMqT3za1aUxRUSFxvjkfjz6lEzF6q0VwpONiRVOYQ4dr2C4YKXlOORWgfU70DK0+AF
Wr0mAVpWxDH8mEYIB8Ynb/fviRakwKj/ABlYlz77q46kOMeMx1GzU601DevnjCq4Z0Ma60dx+dZV
ikQp/SOivyES5TMoTgexezdFuA3x6F8Ovsk3mn/wC2iGoqyvauWa64j2wQ89qx37uwhdfiUG5RJI
wWbFo+fdlvMInnCWrLdswXEIdQbJfudGrd6QFDdYb7SxoJEOUO0fK+C6PBpjjjGcNjr1nwrEhXqn
E+cm0wft4rwQVu2wgLHy454SnSFqJdLrLSLu459y3WByprySRecAc5oK8BAjLDXoGl3Uq1233LWO
Uliep/vtU6Htf0ghkFutXHez7MjzYd83nqWrmWdE0qynjuAHJYdrUjrWkEAmpUi1Q9zurwkKbmgB
1akTZWa8bpyH4Sn8aRRu6U8jT36bDoqq9LdswUe6Mbp0B+4wQMhL2Bg4WaUIwSIyn2hzKMbqetNF
y84utLQ/dLzkB2ijuoB8dxV3mUD1cgGp1odvRLPTB7Lc6ihCmaqGbZi2kIR/TTNr1mG++wA3Ke0R
1+ACkaKFYK4Qzqa2mGiIn7ubVMHN6Uw0s3qDP7TId7EZmBqolr+CCpSfZPdUch8elWZNwEHXxz5Q
QCTdO/S4a0NyBiZmho705V7ajGZnd23zpIDG4o/32aZrKcC2Bo+4EXji4MJa3JGZ2OokSeg+yl4t
AbLSq0d4QlbTOI0UeimQ4JQewBxp5viCZd9S2Sis4td8uFUxIb7c2fyQT/nLP0y+fF533JZl3GK4
958W+uyHbMbLVmual0LmPYFOv/+kxUrGI6SvJrkK7Z5mKOUsjGhwJNe1RVeVddUMhzo/+Mq0JVWk
bZa4MdR5671nvywt4o24nw9K39dhMHan7S0Aky/N00cc7WEArvBzM2YR6I/L3gJ/P3KYm6vKtqIA
oN4Nc7u7ma0L83+JYsYRBGclXkcNM8jzYd2NNKSV7si/CuXUq98KT8wStn7NVXczx7KV70RnKj3p
eYFnjdkkH2mcfORoJ0guIU13v9Xcjx7c2C+wT2aGU0MxbTb4mzWzK6eq9sMwKYjk7hbEePHsEMaU
RBS0IHXaxXTxQd7rCcJxXTPsFd3WgHNu3tZ9UaBuiG3l4HYTaqer4Nxf0XUGF+eRj5cIpkfDW6Ki
SqDO7bQoChM2iBuK1xgHeMpC4krsXMHeBPu2MChyPpDQyMsDK1tSHhoWHpIT6geP8LFw8c4/34nX
I3OPqXzyfibtqGc+ZuYrE0GWYerMrboPfjTzhi2+EacPPJjeP6Y+ZLDkoXt07zh/C1BjfycEI8uP
FQIo0c/iX83drqsaRPN6N2S25Nh/9a+oZsv6RlnxYTYaHggzlxHv8QimFL4g3HPQ2fzazcXjRVlJ
MMzVYNnudsckMbmWkRuIdjh1f3+Qi3txJyobEo/sXiB2Np6kUcpI0A/QoV2Ne0KCeri/EoNVzIEG
BW4/ufT+WuPKcjcFeKd9g2k5+WXQMjIej6g5SdGQ//KNm7ONXYj+KwlF6bkfnmvnuX81F5exvSvY
S29We/3lEPSgJOAWmcekpzCeWgtcUG1JCJc3g20kFPdKyKNBORMSruEhDO0qgnyZXrrWU+pnuD78
POpy2C2yGRFjfAgqstD5l4zmKWYVP/CcrJNEYKPb1yEt1QWYEon/cYnytRfhufLhg08GdjjzDSwn
1YW7WlH1q8hipZLB1lzudCgBQjKEZTGQbNN0r0fGomsnrQ6Rq+bog5mcqRW+neGtT9AJW7ANieTN
Q75mbLKc+0MRAXX6f5RnQGfaPlsXyZojnLo7eripCQ9z5T2+cLT6v4HS0YvRdO0gy3+T0zHvouSF
OdW0qk1YG89y1XVwpbRY1LHMB3B09ZUBUdUa0CmtgKmDfBJdBCXcQGwlwevBRGtU5/ciszpZtt9j
ihq0981t1io4+NPlP+FPsrnMyrfdRtsYcdwJJxb5uCT9z70G9n1EdNQ0Kg+CHXtd0GVHYxQD1zOF
deHOHH5D7CjyGHek48llfDC34Y9bRmFVyHrOU+piJZuTWyYgWjUF9deKGFPPVTqRGAjBAEDuc8xG
uebqZXQ4L7OZg3JkaCB6t6EFjDFguAR8tF4TtYrZl5S6j/I18bu4jwq2MJK40aQq9SrTYvzS/miT
61UM4XKGWpxLAXavLef1EHyfhn4JkE7iw/wG8Mtow5QQ7IIUjDxDWwMwm0qgnw9SCnxW4BaZLS/Q
ePnvmoTVAuon33fGqh5wlcBhuGU/AwPO7lXM2NMXEg+iH/+mosWdOnhXqpBAUzdLbPoIC7dGRRgg
SWJE1n8Zb3vvtPLYU32wHhMAgbNKqYoPOWu6Vgt8StCdUR44JhfZLVQGyx0+YkCPKvNpUfS7hRzA
vONNEorkjGix0q5SmosX4tNv0zVU6vZy7qh2KnpKHjh1XNsEht0AdKSBbUHOYKs2ilkCORk3xVgr
yBD46goVNdnzd09JQHKeKNeuKpnXG1hWfCEV0Rm2EIeyaZ7rBOcrcZ/ydirLWyvim4MafNL2EbWU
3JttTG4I82aa7ORg2gK4F/EPtosxw55pUgfQS76mhK1Yxgi/1ltnHFp1kOZlE/bcGfc/FnSHEHQy
/E2YeaJ7xVWmOefT7QR6jk/j/paSxcKoxYMrESn4O8jF05IMXFBTorDicFF+1wlQgk4mDP5YUHxi
02OrIMQ/iyJ4AsK4Om7VNn7g5Bcp0lEAgvV6dfyAqNW2j9k1KGiUTj02fv9mAgw+wsABf2uRcf52
qi2Lv/PtDr/sMGHC1H9hCB1hPOUjnvXrWKpcQa4+QAWYxrBg8XU/ycv/56WQZqCZLi/AN2peGFR7
JqCXA9ULSUQ5k/dYB5a9Yd5Z+0FlDECtLzPp9+/cB398HQ1zh3Gxr9XVk7wqecA3cSSBoLm2n1Yn
mUG5XiQ03EpLC1fKn3JohKd3enhphS2OFDyJka18OFL/HPLUyHKzTvV4N/0iHsUlULxwsAyWds8I
kkAU9jqY1JZ3MeYhuaSdPjqTKVIGw3WDYj169cfXwgynjP85PEin6dRT81DpJfhq8sHTTQI9kbGr
r9ls3TcHLgSWey1xdsOhbdwoWx5dtI535vqFQJT/vYDZMYl7FYmw38zCrYYnPB+h4ZpyuR+d0au1
3Fd5CRwx5H7051djeh/bMUm3QAd6bL2Y7TsQSgJwhNUbHDNg7wy/CU2XzafDAFOR7mYuM5R/D4mV
XK0n5rfD3CkpyR1Kxmm6bVeij9pF+UO3VXM9eFgUejR0cdlp8dqGCLYyvzRzs3IWWRnEM8FAeqyV
SoA3d401nb960TBRfvD4dfTeBD/w7L3qL/S7bWRTxHOsx95W78p0DlLhJFdXxz7BvUgCngwusyrB
uCA4klPsjxs+NNCIoy9Hr8epGnGu1hJkV+41VXtNiN0aZX8/zSusATScKvSLP3dU9TSivVxraDsz
uLYZLdRFL3WfSWOPnX2PKfq+MGijMeccTqt8NIdEDeeqwsLZ1unCHlUreDVHBPWLYxXd3aleznax
1RtjA1Itw+GStKCE8TjgkzFsM3qYQWfE/bEOconAAlMw/kpj662kaj26328uVQM2Yh0ATD4lrXid
jco001HmBakEbQrKQsPUpa6cL1S+XOAKqtF+KLJw1Pr60XCbRuw5vfCvRHBfXrH9ipPf9YLeWnO+
vNBKk1QZ9KFuZhRq3tNlbQr3Avp3y+3v2h5WqSsme7wr3sOE2pilBYje5RVJ8efhV4Q+09qAMcPR
zxvC/+UpIw501i4SALC6iV9N4TTf5xSulPLdmgLe/4bT+5ScWm0aAObHmk1a2jzDEMapSVkOGBWz
G37WgWsIwks25anFZxYRm7TkpX7HQ0Qq5nDMowIZvJi9VwX61s6vL/yfR+pTJJKcdHdaQpXGuA7o
2BE8xbiyM6amHiyYNRSUMUjK45TLs6uwF4AQT/YhZHLya8RicOkFJTmQHH1xOgTPD90HU2s/KMuE
VGG+sINI4u2DM70Xl4IQiD8igqSWOQxvtaTFORka1b2R4ksQdNdPS2trICswaSEL4dzPB5CqnyPg
KJBapumoN5c2KtBw1vh44G1hhWK7hVQ0tm4r1E7Vzd0oFOFVkBJgTEgqyW1rPwjtFYn2AK8SUvg+
KThNW5nP77JNpWddB4Y/6yvTpP1nZHlNf7o1MQn8dcQtpU2Df0RtyGkAjoKL5RQV/HlkKnzRB4Lv
BNYLgdgDeWDxCJhEgFVh2Y4i4OnS45O61epWIDSJ1ywmtL9bdyYq+WXefeyGTJSaq6v0iARcKGAd
QvAMWbQw1X2wNsGOWWRA4AWcRA1thVUXuP6/96hYVJzd4bAogFFqffYPplvdsWRRYbMmakFXFbsI
xpUuCO7/qjyOWF7HAfcQBR1HeP+GTq66Zy3jMNwlH1NPd/Eno0FB3Qu6v3zdl1QvFV40K0VmaUY8
YDcBMDKfrceKqQC0VufR8warC5NifZ3Tj8F4k+WDlGfmHL3yrElS9RZOFPPU2aN7OBnT5gYb1Mvm
3WIRziOLCPgbrqXq4sWFNvXfzPLohqwPC2EpRjrUjDsUJqHEZAdto0dPjX/+2oa5GFsStWqy606a
di6IKu373oKH9aCNJhgLEP92fQlBgoa8pSNfreIH4Tf4GciLZJzZYG5BsOAg8lSfwGwV2hpEDa8B
aDThVamLNxjVdDBW3Gz13UjKSAzWW+2WHC5T288qup4OOI7g4oMkM9EJIhP3+r968ASw/G8fKZW+
lg7nIKtS4jkIC5wGWokg3LgEISWims+EXXlUsrzFjNzqvqensJ1ty74XW8IankcLUUNHt9DMXW0J
EyUmvuRZM9FbAtE0h6NH+CwEDaAr0y4D/IOZf9yw+wK7cKm33QL+ZHJjCkDFaNvt44yRbam7eHWG
oDQvSsFdl3UjrxRiqjJ+BJlMv+htUNC2fBbbMhviC2zysJVeucQknjTyKrnT6wQ5WaVBq/51ZCJH
rYOGt9SJzXD+YvIn1yH4lceI1wakyUeYYY+HJFaBZLMvMjOkYRSM4JjN0Cqo1p3oBeo3k4wSJz6r
MCCCNwltk+enVxmzvK9AoSgykHVxsxg3JTz9VHCm0KQHnIUMTQZH7EoFBhNV3PpeHtYUeUIrvPPG
IkZsmQBdJkZDfB3/MHcOSZmGw7W/UfC49TgKdtir4/J4cr8MZKtl9sayYm/JakYBvx2p+9Jq9GZq
ZacEH9E+JXJJlhm/6HL1VDW88FM7YLyEyauWlCbCO0f2BxvGC3UKjBby41lLn0CZYVA95+T3z8MA
ixaViVj4ymhNqF4TZ/dswbuG1e4W42w0o2TKU2yXrM3bUB3a/yjnTj2woc0LS99tk0+qby5jQepL
uk3MWkS0kAJe/+HwfCdlW/9rdJXZpOMxbW+1sD2PrQqNq9eYYKegC10ilxbqW4/jp1nD4j+q5ifT
pTfFoo82TF27KqV/WmNELWzda5+pUZEVFKVW7XJJCfDXXtAAy/x3LfKE2H5vLwYC358PtlrxQz9T
FKBH2U1X5aTGL8rMlSM2uqcewPvC00VIosUDLiqgAqNbTlPvbOJGr5r2ElULLHv+GZR1npaUws3z
XXeKx3aKRG5sBHy2/ocACayLV1eX11F0msA6RQ/rJY/+OMrno7puGKjJGodcSsCWH7+6isVUkW/8
Ykqzd0uUtvDChwEMzH4k7wyXP4/S1wv6SrsuNjm6g8t5jrjh7teMTljwvq4oMu1kyImTLB22nMNg
6uqQRUtRIZLdXbSg+Vz0tfsrlz2jYion9VcYetBTr6lDH4JSvwv5ukOYxLkZhkZDZAqPwtsOi2b5
Q9o/ta/AH2Tac4kTSodgG7boOEkodFto+OfZgHr06l9nGQd19wESAhB/Pquc6+SkxgzGS8TDhZ1H
1T+Skd6hdl9mbJR70VkLFYtcTHdIXPSCy9E1ViiEEBrp7Q3cwbpO8sW0qft8l752H3ixa8F391X6
L3DbcIke2gnQR6Hm2bXCft7t4kVGBxjvYxxCnklR/KDg5GIM6KR2ez8XTAgKJcd+/dCvx9P+dV7S
UdISG5sftWpa1Zs3AIIHmbrWKtZUMW8ukHKgMrn4+xOxkrGKQ1t1viFCjjc/CBUjtQhgGITp+fdI
JOiiJQeylbSchQWvtXQOQAYTNw07Nh8J6+QEub9dv/nlsxnIHRBrJ39YvKUNJDFiBqQf3GMy2lp6
LTOfSOXq+Sq9YMwYo/3kKbO0BqbG5e6PHNLsj/fIKrTmfzPhB7vv8Pm3IcoCGhJg7bMZS/Q4XVZE
LGQRGHetjn6BGcuuJOY9r/+LxMgez/mjvfTN6nWx/RpVHZfcK9DvzeoNhfNSV4T5zCS3ddZCLTxZ
R2s9/MTQHpPBvK8uBcYaG3WjBha0XRGCU2w2EATBlGN9VthTgJl4itKbgo6SZ+lt8uSXOORT6jJq
fPwYuQUaNytO+6H9TwuAmjsKOZgdpbk6aVDjxFJlIiNeEa2s4AAHvYih6gqNONfYnw5X4f9wGGP9
PrDaTATgHA6GrMP7XgoATkWBxPVKe+hN2wdlLwRmK6co+HiOWGceAm6lnIDwjgCSq06tqnj0hh6C
Rt/kbV5v+R5KIcR1DDGD2glLH3MlbI871hQFbM8DROIUIrXmkqkiE8VqMtcj4vBFm9EuKsfP7sQ1
NFpfOkhNGBe5E4S6xG6MTBJK+WfIF9v4sEDUPJAl9Y7ngc2O37iFoehOtPZQNpWeZM4HD42c3MIN
Beaxmq9u7oUmBirULwIyYbmMuJzJA3X/wBKcIRMur1Ub30doQPWsqKWfnfbLrufr21xXgSSEEGEU
l/J1IlQRtxMZq4NZiAdvDBb1lH67T5hqd/XkK6JZgweUNsyXLECEpAPhaxxuhTTBciJbfQUsZ4pk
N9I2WcD638Pi+WUbeXwzJlKB9Y96rLKRY8RkST96aZ2Kge2yO0BdG+uvKCpGDZeAsjXGxvqvR3Qc
oQ0dIqprq/LMBHZw5bzVSr6kqzVpZEU6eUS4Bn9gdp2zLNa4O/5q6Ohw/F7pBi7nYfPNIAN72iSA
eOwac7xSY1RDWjq1Q4vz9PP3I4lwMJXC8/RDNYQHu/WL+2heveyF/ImQ9i89VYl/GgvPOC60n4eK
98B6YedzHDXW+R5OSHj0u/ya9KDl7EOVIkvcw2cTWoyZMqnsajdUK5wzuYFcCY7zclE/YiVnZsNk
OyPKFda/J682Nfs0yzGiEFPvUSO+muv2TzFGPB/OvdPdw1gy3W8fabJerjZMZrhSnOuRII1PAMOB
UiGoFXxAnzSANmbx6UF8MMh9MsGiXC2jy3wMbaHI0TLylJk5dZxH45rywMYBMEV17jznedwaKNC2
l6vWP1n2QWV2y2frv+vBlZrUdKH7g/Z8ze4RJb+I2+bhZ1CjpxB0Gt9USRLJhhnkU7mwqOx8YuJY
fyJrIMy9/RQNGDP4/Q/a3QNYOZLAboEFC7Yf2H7BjAj9WdiOiEb4ci+oz/txzmPcwZWXN7kMMyjc
1xqCrB/gh7TYMkeONFtKYi8dh6/qMxG9ZesBf8sGfsCWvWlQ6V5QmxEEmtNdllb4Uj+W5Bh0MWCC
3EzYCAqp6Nq4IZljqW0vNBHHtYS7M4mghciu2lBSP1BGNdB2fFlb8o4I4kCq0JYV/3Dohf3gPzvt
mlmxizu1dOtifTJgzspyCcE3NNsJtsz09HqmfJmluSHwt2crT5Eo6AxTCntqQXJM7NtEresWR+jd
Te0KLzEM1WbPmNsRXTerLKjfogsKm47Q9oS0/zvUIv0D9f0r+Ooxg+YfGN97/NNaGJoOjdv6/pj6
jpNXoe17oKTuB05qwgm3L9jGcA5C3eJCemZM4eo72sv2VDtMawc5NQnKQrZVD3EzoO0U7a9wXDcz
OdaVKWN/RAtAnzveRdSb8aWGYE/hvinXpA/dVnK41rSfmejpxiGCZkQD0yBgyl2ytPN/iWDXMY9m
zzYcP8fm3S6/3ie1DbPH9g1pFvvIg+kt8nzCt/qT46E3xtIqNaZ3SJHV3tHSIB0KHSnbtZIQblw3
mp9DuCyUso7jwVutJp9AbxgdCP2ilV47DBMRryJ9kVMfexQtjknPUcvKRHi/f2Pk0ipmoSe+AtpO
Ze8g1fVxkuLXRyhei0SiYbecAC/hej6PyG74FVdah7/s7ulq9f9J0dTAwnHMstviLhbE8wOiLWVe
z7euyERSfL6N5KkDOeLLAVugj+qHdOa8lC9LU+xQ8k/78l9C9qNRpZtq4uWf3LMPOfCPT77kjQZH
YvmNnTvXrMU2vrSi3Sk5W0Foxn8Xfb3S6o69z7MExaZSLFRP6+yCHeIahxXz5JzAZTCAhD3ZJnPE
xOwmO81n1ULK6Q+I9cJh9azUrQHG2zEzoUiHL0Jch7FhyxfeyJFlfcA8l5MJE94NSbbLflK/VFgm
nCTy3dRD7bKwf/qz7PLe75c3YOPGRa29g3n5rhBTKq6RfqbAKTykEdt7QOFknzDV0dc4btbHBbHH
rShOuRXROMzh1C+laFAyL3MvFDVF4CKAK9v/3QLFjB+zHk7EIa7t0QlqiyTNl5jt33aO+b1RTLjx
YQPMjrlB1i6BKXDuQferGNoVZp4ItUPnLw6TPXvV+RpskupOeuNl7IR/uQCrNx5aNSrW35iVQv0A
WXoxUYVIAVYx1v5GNPx8YXx8HtfWVUq8JNMkH9u700D23L2SdKQ/VGACavCLL5RpRLwG70WRBTfS
rByQtIyE3cedGA/ywkAXFJAvEH2Jkiy+dHRwkQB9Z31RDcww42wiVIqj6oI1393FfoBfKXOFrxy7
RFqb9mM3StgJM5sTmensxeshPibQTbIG9cdJRVs4yFkogHUMdHo4ah788echam0hj4oShTKIg5M6
aYPDI/vYldRyVS2X/FOvAr/ZLBg1OEWZjPWAwvTsxAg/ZRVxb09Ky4NJrb+VN4HCa+uNsJkgdYe9
vsko8SvBVHkryKNwILLQrYT2ONyI4x3wyUkpVqbaYMCZk5u/gi1v3m8CInMjRFEl5ukNrykM63AV
t7CsXh1I8qE99NIi+HRD7oM7UIwh1Sc3Mhzcji/VNy20T3iYDoUXPuDorFBE5QDEQmBzz/Thi6sA
qTGICvao6Nu5zjWfJS+6kfuiDEdePuz/HC/fVkOSE8XFbj+TO6A5s3RwH6X0T8aap3zhOYPImV17
emIt6/0byXgrQxNzmwlkofrwh92+jiZdpeIz644MA7ZEQcnJYVfzQ7n0Jof/J2Yto4XQWB0EKpZ5
RhgJ9bUoLYwu+nSMRFmlPpedcHVfAKMAtOg/15Yp/a59anrFb9E9O3mcB73k8GkGKEMqBBPjZqyk
o/smSoyEuGtb6SD5qCagycmzQhzWd73hBYbZsjMNchdS2XvlAJ4S7PfHxC2VnFHoqZuBAeU7P0DI
z8RluQumLa9UFRugksfH0b3mtKlb3cMRfJTO2eHqfSqUDFmavV3O4+vjA/kqnp455OlT1b+8M2nV
xl7T6LojUWvOHTUcAHpLyS7a3wN+atDFntj9kzaJoaDl/LmYTcg+ITbApdqu2z+Lqx7sdBzHxLv4
i7s5H9PJOl9af3AuvpM0Nh1jUeZh1L5svsekmmT0cFPZoqqI/4biHmUEfBU9tUwPHhvTXQRoNF/y
ckcy1cWgUtK3Fjas7litCUUfMUzBcAH4xQYvRdMPkpWs41qqMCeeK2NmHW+9o7FgSkpNwXY/bglW
Dq0WVw0TAmdS2TEhbNMeFizdklAhczpXbay6da6myxttlkA8RzrLCXhFMiNTtoyi6CSo3wUkQyqg
Ziitf+ynZHI/zog9nZ4Da0xESxzaKAnPHfYRGf8EqPH9+LEwuc2hOHIG/LKNdsqmM+Hmy4CTuIxQ
PlJJ9Jqqd1kXG6sXm16NaNKKITu/k2XfIkf6F09T5geFazioh5SvxG3gvQUiJA0RRo7pTkiarJR/
F7+bb1psZHjBZfRbwkX3JIWYknPou8bPd7sFRAcqaaCXQPwzCYw6sUbmsbZGi+I5wBWpbJeCLTGt
44SMgbAeJM1ijO4qb/guVq4pEQuFhjtfKw1ilG6q2HhbOhAVC36ZLJ2yrCVsbx7zI33g4uH0QIuP
UhnG3a2ZQXj+9qeZv3Qq9c1w4WT0veagjQZpOMeYYoz7ci+HP8HEA3tdpX+3/u+/GI/1+PE8oT0L
TdiZUMFb3ES6uHtrsB2HBWZ5vrUmBh/u8u0dCa+qpY3IiPZqKgLfbizDVFjulhNVqTqS9Pjm8Z+5
guU1fQUBlfQ4IWAYH74WKCkiMXjVEKAchMUCCLZz8O9ilPCdSBAwzGcnVBs6DkZ4D7tplkmZ4saI
p/BZpy/TxnmouxMZExo/5UZBaUFBQ/GXgqWSLoHhWFb5Ppk0yqydaN/8+csT3Ji1O5lbnKrxVEde
gUe7o9kODXqyIaXkmlenUgLtucqBmxidSxfyrSgoX4GeMx6MphwpATaliG//tma9vlle+iT7BRaQ
3FMM8Yyhr3B8qYj6DgoKHo7etNmkRtteh0FPriBK94IOplW+e6Ny29comr1RxnLYvpNWjL/1GN6T
o2CKh3YBDHCMGycScxYOITvmaFdo8I1WCyZD0aziBERahIlV7e03wes2RN5o4O7ohXNtG2bbs+lu
1KDXqgLF5mFIFU1sC1yvMsXE/gh0zVMxBKqilrR1rPrWk4/LxiJc59QzLDqHG0ZbSvbLPrUi9yME
Fy3KfDGCwjD/v/KvJl7V2hfjcRn8GnIt03e8dPhRb2tsMcsx1S6Qf/Odj2i5AuKGEtkcDw7g6sjr
GJ/N7sJZj5JwgfoDU1KFT4PDzAbe4vfk1xTvp86JhfpllRNejIHngLiIrwv9MgZ5+Qq/v/Ay1Tay
b4xmO4Dsq3nE3sdwy4rVzCbpB2UNsJZwjRMYDTTDipNNYditlYmprji3Xv9K11ceaS8DcK7RrqXd
qtvKNisoyWb0PiGZ4x1WufqudputG7ltIUhV4eP7lMeavMKBssqb5DQnHD6ib8Tozi8XBl662b9C
Sayuqqdm0dGjpqPkXB8oL6rryG7eD5FCFVvwWp8XKlCoAV0pB6ApIM7TpKoHF3AWMSBNTL+GEUzQ
sA3EfP7jAB5fERPUVQEG47//yaMxaRUbJiqYkElW4r4LkO5ewJDuIUFysH0yfpaYYOuCYjJvtI07
nH6jT+PktK14+96HU7hhUfBk87TGmUnNPDAcGHenKUGk4y2Qb1nOIxMAPw9nmhLHUnwaBpF22JUU
9tGu8Rn/qXVfHixvMNDjevvkiNVc9kqIiCmhg5OLU1nVj/O6/I9cgLCmG9/U8cFg69TVYDfiQKq8
GnVEy6+tONixrrNclbmCrznwSydbJBz9yzmmt2sQzHKDrhhyHw64qDpJmon/apEWry+kVVwj9bsT
+JoBKGXuBvknwuE5yeMLffWJ8eQnpu3yFDpgRO39RYzPuOQZKcfVfL4iGdh/7t9NNnGPn4iNKcT8
/0j+KtyVlcRUEB38pcrHDhFcZrSIDq3sgEr6IJ+ADPSN/VTGt7fW5zSZlwrsKg7qxYF38NlesjfN
Yf2fjpzNJA9uO3/fGu1en2fJFHZQyPuvK/XIZOjl16OroloawFF1QaU1vnD/4yf/r5UinqT1iEC9
liYfUeREdMHeZW92hckAcWkkY6XlUSYjyW8UDaVUaO9EgTTRwOFvOD0nvqWvdAvpeZyi+LS7apCI
LOcmvf+CBQWLfsGnbTEmRR+5wNaZR+r6UzhzPukpFpg6cOYohivzAKK6uy0Uy+bAwD9F/W9NSehG
lsceVpeiUy1tmgL7ozsE7GcU3KQoBXbmAZf3O9R8c187dYl2GYEROoOl+kTkbxa8bGoWsdYe+UYT
YgKxN5ha8++Pe+RGGssNeKSb2hzcnWG1U67gDWR2NMb5jzuqP7Cwj+txcMRRVQjxbFpz+Rr7my0V
lBFZAnwi/7NJj0htH9dtGPArrHoA3pku2aqr3ErNFYpSYVN/PrrNbH+LLz2tGR6FBp4LFTnX4ioG
yCOLuAuN58bG5tVvcusIkzeLDqFp/EBgU8yJU9G/g2mpqHyz7Bnxue61QL2DkavsVE02mHtbY7+2
AkXe4WzigJFxP2DgxXsWhyqxyPDeRqb0tbeTyf/U3BNPo91EKi0ex05qTLSMPY7MU5BGf98uvSA6
SYdQdJl5UG/qvKqnFIfWawMS8UTrscM3KcRynAbgapXYw0fN9ZDDsztoVfETusn08aLbIqG4ga+a
6fBz3qL9QWvilOO2fv/hC6qrJJJh4/fLd1ButJUafwmu6D1EiCkBHRVkVSTVTh7xKmLR1C40N6fk
ntqDbUUmiiR/LLVLCYg3yK+GSssITHIpxM3vq/0UbIeB+1UXx1Yr5FBjZOmOiSZMGFaG+KPjo7LT
y24dTxUJ65y21JQbWfvlF4I1KszyfvWmjw4bWAmgVCsvu9Gm66slXRP3PgOtqmTBe0mTnP58Zn5C
Cp8b+uTYA7yMqrkp7qDaAZH+/WaRw3PMvZzubQCQGH3BdFOM2G5huFZxJUw/IH49eQRz6ek2LVcV
PjBIuu/mi3JgZpwCw32+XQ/zmhIeBvYVSTLnibwoRUuTDCkzzIeZuC+wV9Nqy+26vz2xnQAzuoQV
Jp6sPV9NpJFfdK/cvkA6Oqueq/R1Rz8EQNDiLJ4GEIGcVbKRh/SqHH0kIq/pFqF7jArPeBsB/BCF
rYpLDqoUJTVixqcBHKP7jjMRo1pdMwvYeTsOOixi3e7ZhChye24reURloLmxFhOSrofL0Sv4V8OM
wPLjsBObZbS07GSEbpy6rBiCSTtJ2FRACF99SNWrYhfWfD/wT+aUD9Cuaeh7IN+DQi7dz+JLNASE
dzL2UbIl2zP5PiXnO8qXZ1DNuN0lh2kRIWUNsX7V3LJHtPEEdxKsXeiHAQ8rlUNwj2uajymF+qfv
rbyHs5va7Ye2IBt9JmgVv3Kq3vPIVhg9pWayijAMcLlixOBQb2+3G2kaeLMpBDJtBlaRVdO5D6bc
bFa7/hufR8NECjCu8FeveC7uWMsw5HkZ2U9bBdLOYD2wxennDJiLV7rCOzwVNKPPxDO7mSs+tpsW
eDMDODW8uBK5O2nHUq+5rocFcZK3wYGIeqzb2uAI9HHrMFCoZ3Z59cJ/mMo3z3nWcdoHCh588BOs
L9bjNLl9ACSv7FEZbSzt/kaky79b30+xPOAHLwgcASZhRh/smhxTkq2UBkzMp52Ylsd0RAaHxXys
tHxwLzDzLBti3cL9DDDlvaaQirr/pRxxtMS90ls38LBvCRYcJlnVCDMMIlQsxBk2RIIAX3F8Mooo
PSKXoT0epXsvph/bKKmJJlQgbt3E+YTfE0vm64of/zR4aY5JkYITBP2k1taxRIWmaLcYu1MFShhx
ZZtBIVJBdccgcZ9yPe3ogYEDnxvn+vVSbET7p8VHbjYR4BqE3vSsmgLf1ENh04gGrqGuc85KdD7t
zjdDy1nK0b1DAsMJ5JqX4bkTsmjGDpdSeBDlc/AU30U+FqPdDeJb0uNHjBw+kpC52SLTo07bEF5B
QluVxFVWheC/3ll1bPrmK3zkLfJEfAGCIRK5pqloteRR+W4nZW4sUk9Tk+g5qX4uzHPBfYYueFkS
3pTiIheGBAD766DAezV2z0ysc+X0JESWiB/OqrphhMfngaPxdzAS9Yqvww4iMcxcQQxTmkAG3y8K
ADaNUa/4w6OGUJr6xFjG6bzXfjq3KdgdwrTe02H5cjRXoAfkf9ls30vqWJ7ZcQF0HgRDebxUiLz/
wNuj/3D4oTq6epN79PlOCQucKBxayxhYaxiRoQo9u9iH2DUsktZdJyBDim1Cc5l/TS6qIHUnHWYC
6x9Ogob6aSEaZiW0xuUpMuX+sQISJ6N3X8/EcDJA8KtMTVb67lpCRvxFBgwd1g0h0uZ5ImXqWwWi
kEAl7ky9q2JwTa05PijE2qrQkygYCK2ZQbZsShLpjwcRu5ZEIEWpcv9smNlGOO/jk88g0604RAM6
M5J5fg8RJRIdMAz0WmFoN+g7gLhqmpEP+5j9jHJYKqw0NXm32Jpkw/JFEfUyHG9g+d3ADs51wNY0
AnqGjzJviHMNnGxCrMmYQ9RhLVRSzt7x9vplHpOVVeTyypNQYoTt3FwSupWBoGeCwTpZPG6WKcSA
Ww3fMjFD8vEEncdJbpKZdS36UEy4w1M6QT5m04eUOMycovLHFQIsJgoZUO0BuAYOHJcX0KKSalpK
JSf54YMNDTyNEjiQGNuTtdG/m0w7Epr3d6nQbs7WUIGOQZ/Dwt4q3tpPaYVjR9IrGTvdfwVtIjtZ
dm6AqoM4NjgFDpez41VKE358amdwhsYjWlIPQRGfLslQuQG61FbJAU8NoV9wp0EBPN+3WTJBEAd5
7M4AnSpXRTs8icsd+DllsgUSclsPqPXDLX7hhnQ/qYGyIiWqBEZxYlh1JhFiltqHgmVc+UNOc/1k
BK1alwthiwQC2hE18+h2M/ArcG9Wr4GQo1EGv1eBIc/gJYZwbDmhSrYeheSZLtFD+SIpPconVNt1
X0huSohtxl+BWRAMMFxhUREBCh8YDaYdp3dAPQBa/nrUIWsJrXOARN/Urg9y2vXBRyduAZTLtPYc
WDHVWe+0xZjQDEGFLvJvKi4IWDGBtiOxkbG4vlqwINny6QW6A7guIDOk4wd2NQzFScD+a9JnDR/U
gTz0PEF/jSCC+33GbySSKJGNuTiQD6u2SsUw6VGtihbYfXtk4dlLB470kAZsd7QBUwYlAFrJK8sk
cYrcyLSmbFw9M14xtr+3Y0eNbY63skmoyggdRD5Mm7X6dA8TqKnH+YiWjH7A9UCRBxlrubVy+af8
TjZKnTFkLAqkhMgT6dqH6D804oZfzn5beVAu1X/d2g2UbeVfszSHUih27nzGa1kw9L7HKkA5Pglc
o3Zh6Lr8pE6mrpgiA0hg6LVm4Gn0fezAJZmR3l09LUv1Yu4lUbUDk+gdW75H0C0FgqeF5rL/WCoY
gtrN2zW6E8JUicMB20wFjptOdjyNkaMg/Dww02dNAZZLBEBYDBW2QG1kCL2AegOXbtZiKITWwMBh
hb9uvIrzUuUIn/73yWdCjr4ApK4FLwUDUM+4uz3MK4pi7FCmsaDpghSPre0LcZZF0EEJ0JALDpkK
r4vuc0bHzs1AstjUamkR1QnMxiOrpkaWrhNuJ+b8YEpKcynUta0mHheJFNfGm2HCpwdtIsmrQeHI
G3z+2+Uex4bQNY0HjkY6ChIbU4fXKhYv8xtnjWoPX/mBLGwNHv8Qv0HAPglZJ8/PjmzxFqDEkzDe
8mA6SikZQg0wSwEB4oTbl8ZDenTLfEK30/ADfrlZUj4CinfuF9YITG1Sc/vBhWK/9N8cVUsXc+t1
y8IMtkVdIeYCm9WD/vghkce/qd+rQB9jottJ58sfsS3COhXqQGx7Kt6Xvesx8VTWeEMzZ8nI2vrD
dfvzvBYFnLuBsUArz4XzVap+RByAHfyleZ+V4amzzzFIR7vfPRu0pvfhVH8scfHUI7h6Aibr95AS
fGTDrW+TcZFVwgXVLojERekFKwFcs1EFGwL3gR5Qfdmml3y5xiSwoBMQvoo2epWKp3iunLZtWcuD
48wUuDDWLaE4sMr2J4iO3JMK7gDFzXalCeE44eLphj5hrjKVwwWEx24UgWDSICXRTQlorZ++hPX+
K4k/lXL9rbpz9N/AOM6FmRglj6TiLjemnpcBBFKVrdFzViHqoKAShtC30lplVOvAPu3P+o1z848D
w6mG3z1BomPzIB4o+jis3mswg0tfXdiZXjZUks/3MnzxphlYB1233AnQVA2w9pAnqDLy41hZsuk+
YujRI9H0gmottye/9b8uyO1YP0iw1pmdRYhahg3AqnqnDWgzR4p2m2iDfov60ImVJK6xspGzMuBY
5YHvltz/2vQR0MTJMbgWXOJqhO1/MrtmvXdJMetgsD8cj3HS1x15We1GdRlRsP8va4eui9Dfgeiw
2tF65PQwbm21N29e7DhFPdtR/c9+80xEFOls4RRaIiP4Ai7d2dKxzDPeQHHtm+yYtcO4PyrBT3A5
K+lO5RrDkPzZGflnMGx+tlN3j1s14xj+mk9Nq6fa3rkzhffgo1CJh42u2V/zxlIslkMrz+3QWzTi
O/Kovddr/+jyPCVTDCCYiPdH/u5PITQRPHQZsx6xXeYKR0TDw7pGLqgvxiIu+mmw5s+R9hLvqIic
Qq1wjjMaJmHw3pNC4MWh59iXHYW0NhHORx9GUBzJFEFHX1OlpYyX9o3KhEgNsKivjM2VWRWFmo2+
DZW434tZF7CHK9RXjKz1RQuUZj1ewkoOvma+3bPaCNUpjdMvxiqZnqOtg0rYM6cs3BEE/0fR3bIm
3RDi4V3GKji0xio7BfmSQyWbVMHH63kVrfALnBgoYZg62LaT0dnOe4+4+m/KNlJZQNYqMTT1AMlS
gf6M0B/tjZwJGELdOHV1hsbONTkYw7cOtveDft+I74HoD2zu5q5IZH3QS5Mu8ioIZFtZ7M+9k1LS
+Ck4p69thqnfDtHehMp/oKZz9q8U2mFB/D7awaJNMAy7X916I9GjVAKGbOYDupdkSUV8uEUKvlKv
jZkFjFqXw0rsoL84gXxE1uzQNsfADXB70SYvAMhi1QCRJGsH12WTWD2SJ4cc84yRDCgu6vmi30Ce
1s/x8Iwkgp8Ojo+gWabmpiJArQmNAPXmzd1zzx3HLjXrtbtzrLfqc6GORTeOz5bSPjpcP10mRQS8
AmqV3PT6v1qmVkKMhhLoBfwjHeFtTDCWUkeSvunzH9Y2717VWXNcFau8RQHfc8bIYmvTutMC4EKr
jfsf0wKTUWqxI/l1qls4pdD+Kf/uRu/4UZDePsMnGLWj4BbNeW7N/6n9RWTvPs3eBIfwYqgnDVpv
qubQmhX2h0xwYN2X22hABpykM5CzNjtw10V3hACPfND9k7CpmACst3Xnvil5bakJEvEgx52Y2n1P
NIQeSb+g/HlF83Etk7wJArTJhlD2H9fzItEwriji/MuCaECiQLjYJ4YixviVTlkJyvkHChyvFLJR
Sdsdc1Yf55YBLE7vfuXTlaAixAfjCvIzmvU9CoFd2Hasl1x9rOtxne9e3JrFlLPY62y9puqXoYnE
6RM7Owtb2ebRfYVIndltL6Aa/Z8oxTlodwy41yPqExyKjCg0vPyYL/H5dJR3vCe5s96NbL5S0eCA
x6gPgaODEorm1nXIO883RUmDo5F9QbAWFB7W/bONXZ/0xnP2Q6uWqP7RIuU8Jl7O6jsBjo2RJPpc
y11UDW4q9ORHg4IA/XkbjholhA4vyjvTacAwd6Y5VhZzncA+T7wNJORODJtL7LjKTfeaeySdTTT9
b94/nFKo0MOhpkUNTs5qImi0ddiSvd3vb+ksjrZk63IxS8C/KMACo65P/5VnPx1KF9bOw1UCNjPG
hAaidCGGAJTTb8rxm2vnbywrxcDd5X2fp0vStrF8Sf4mPzHmooC7oHjhMXLQ9vN5nF7P34TzMDdA
TL16XBagQr4KhOfnEalXCxFhisOBICQxNs/JjryhR1Sum2/zP4S4AR3pt4dmlQzXAd6ZOJ/38Ya+
qvSx8WhphOpvo2Z0ww2iYe8128o15kSO6EFmqzx5LZg+ta94ZPz9A3jwTL0GOAjpCk6er4leb+5R
GUe2lqp/ec1H2m2EAXJzHwM1aBCmo8HZaD8RQFaJA3QpJh5oFG5Kdh+deugJlcs5tdlhqiHSFRB9
YeFORIu3TPokDY1+wvSDUqLWiLSByJPJpyHOPYMISwn7gx0O7UhFXcMQwDtc5JdhV9Wp0Jh8sEa0
48EM5wuSBaZdahSQlv0ADIxxYnEDMSNVyKL6GGgHbki8NvhVeFS/CkF0XTwQCsxYWNMVjoPX9pMj
FvXlM273ExEPSeUsgWRME1019fmiej7nDNlG6fh5J1Q37C+WBknZRVhEeBvBN4hnzgbCaUInctdo
JUVXYb5F2HG3uQzNnmp6jcCZGuakx5KL0mLS93xoiMUSuvQw9ME1GhUq9XhPZdOzVmh+7v6n2yXE
ITGRJ1NZL0qdiLOTDgbRaXTEuBqbJih9KckBSF471JseMiVR/IH0gBFKzdqc72dHaT2Xqh/7zfNp
euQ5eor5wGASfcS4Nz1Ay2Oq2FF4bQKC70C/5TOyyffuIo4e/VxP4dPo9NWs49C9iUTwO0j5+Lsn
nEG1D0huDW9J38sOOUxlblGQa3sDdqWHn7EG89q/7cF5pwBdcs78+j4SmES1HU+sDxXjGZ4UooCF
pECG8bxL6Zn2BTQY7veiX7cjyINZJMS9wOcjRElCu7QUNIo6lKUzCLoknzJe9v9v5JXoM6Ib1Ccz
RfWUs3qbls6Py79nTwyfIyL5hyvYX4WqEI1P6OFzGN5s1b3ERPdOMa7OJ4c9WDxxF4bal9uqulFS
u7q2+d9RGiRI8LcLfPLGRGsO82z7UJLRW7oegWwAuW+9gE4tsK6IiwlDhMBo9444oPVGkiK64xW2
TTWxj7NDv1ulvCRP7N298zAoyAmFN0FAwxq8bpI47wNLr+gavRihSCD2tQwNPRMHc4+Puyyylzl+
Me/iDG/rMKCnlHVwgrY88bmzDXRbNexnSQcJkO0nhWdH4ie2Vq0k9KKygsycibNTG5E1aOGIs/gB
AlzHlYudo6DwKGu5Fxv+EbagMOtMtalFtuAaQvn6jJA5SbY8qmii8giTvrhybXMXlD7g+z5DH04/
SxvNc3beqF69iDR3rvfuFu5o4y5dnQ1RkWC3uaMi01hXMWh8UeYpr2t37JLxNVAOo50sLA1GtljJ
2uIzEFp6HiPFeuB6v4+IoRU9q6dNgMOjSRaERoyb8cwaiUcGaHyq7K9TgEYnhagQdd25wlnQfVXB
tyCq+RJvyeSzvvFj2nD7uOhsuOIKbda8FiorD5FrrpWhOT6iCkeNTGF1rJgzwnAhEJjZZGLnJ2Dy
tzG0X/Q9ZlpIpTm3/xY9sIUL1k+e7KKCTB68KqH+Him74uQdrWLK2t0kc9NEGo4GGbSU8WL5AW8B
PGD4UB3IY2BlQwSHhmNZvHtemrlNx2GdQhwR8d7lRzKFJ50aszyuLZ1Yf3x3Zu5bE1baMRYwkEAl
Sl6Zez9Y76zbNeIwK6bZszvCJ4DUPiB1a/lku3MBBTakGmzspsiG2TrvUhmgDPAsIOcNHUY3zqDR
rdWXlw38k2pE36Ig8cEz7KO9n2Dzewc/z8E0XxAhtaPTtYO8TONXciuGDVI4DSnHfWZgNf4Boqdd
BmeSInJxNukYH0KkArqgiE3oTlAPgjTAntgRl15BDTY+xqatnaQnhaPaMs3k+hUlZAFLT8qaK2dZ
yCYjKxgCHFPFeaFWyCxyZDWJmd1vG2YDjwpHgLXWqUtz8KVqB3RdKGwt3tR0yVGgLiOFb+LDBlxm
qMSOiCv2HRyqQlnBCpMuucIcH7xdBHaW8Qky+Kkh1JUuxG6MSrzB8NO5mEI5csbCBDu8wPUCeceb
wA4DM7LYq0+rhQ+UTasQt8TaTcYwDIVIP1wG98mW5i48MiYSS20FLvpyooFNYVlNYACMwWbqXjzY
XlqiQA6ouloTN/KwHKVWL3HLYg7OvPRbyyk3pQaCtrkB8x8vLzx0HhvyYW6v1X5tP42H6eQxrkKi
H+o/rdCff/SUwPZcStwc3KCk9cYl7MxcSpOEgBMI7kFtsaLQDQGKf1TVFlnSP6/xQTg7HLmwKYQ4
Le/OVINb+aiAOWxWBgzyMAsUG/QDf7G1BgioMYizWDCsMMgp0aFCFGJkmM4+CDpPioHPEL/dcxDJ
Mbe2Z4MQryQppIh/SvgXHt6Azq3upxj1UXeU3ruZqSInaB9wXcVDDkXER/xt/nN33dR4R7JIc4eX
VYMM8QGJhCLbMikkz9oqkzpUINKbBnnm+eYYF/svekEBYmN1KoJNZJVsbihQJ5fDjPIKIyt6gmqB
tNQKpRdnlBEPNtAC/RD69gGX4T2Nof8K6C1Vnq6/KfE8fAW8MzlfPzfYlMpfY0Arz34uLcmov1Ua
6ot9AksClRpZSWeK1EzV/DKiXN4+Ojq+57OBTWkoBj0+/G6TgPN+eWgkYd9/DmY7gnohfL4V2YpC
Z80EcJjdeoswYHZPiIzv+N8H3gw1evoG6LrDzEuHvmOCveybH9xwdKa+jrsz231LaBRFxUIIBZJY
+Vn5k2IGVaqOyiPSdEoWhjSdtHnTwny3GNyJjfKPPkmeTVDF/XNkiz/eZ2+9DlsEthbGXStiUo3Q
kKTaF6BN0VN7hWzZbv+Bx97Jy7tmr1P6f3Ue6SEjnj5syaAdi0fmf4v/gutBjlNO1sW2ykkOnyfo
PkuAxmCQw8eAslJap4l0rApPxEdqQZB2tDJslkVq/3zEf+lSDdQtpIbKZonsO2X/5Sa/TpdA45n3
06fYzyTbSzmx3vNyEhRkY7HB1inqHIUN8tLaTL8O3FtpXuV5+oBFsVjhaDgYJua44ePeOBdFCMMM
RIYbe6lF0B+sH14Yb2luxiPC6qwifv9pjD2vYFPo6C7ewkY9oN1C03mYW26QdmjIAwBeH3DFhse6
Mx7DCCEq5+Ml2rQ5RDbsePyMEGR4AeqKpggm7v1HSr77WFuU5+O2Evh8JSnbYfR/Yr2Id2qZ2P/5
O5VwrXDvD5yU9rSlHNNRRr1hXHIk4zAIp/ENHESy9SzoopODR4QTGmAxiNTrOmV0dTpVcDffMcR6
rMnTBRG1dMXpt0r66dWaJscGV0Z+A6jJwhqED7QU9t0BgC87kbjYMWEuDiTOxNIlmYnh7Ki6YE4X
dbyxmpp1qUstkSbwTzjC69vw7vpk5qk9SQFNw/m+PUexa0XwHudrBIRjDQJqDj7cf0PW8B0pvPFb
cFKK9i5XnbX8NmlVdQgQNKY+w6c2c08SCIhixqQNw1585Lv5lV5MRYOdr5WFyLeTR0iFiKH1tXom
/81ydIUIQ8YtZeP78ixCcw+rjI8k4C62xbm5Kr+winH6TnFMzmD8hCPOtfNh2e2UhPitEGr6qNdp
H0BEjRkcWXQEU035Vmz13SSHo7KCh8I1L+PLS55pEPF1d6DyA+cJ5CeNlN1Bng7o90HOU17XMEiJ
juRDnzaPPPzp//HsCUrNHff6ojfT9Utgcug0NJf0edhd0U7G7bJJZUCLth9ii+S0rIZqIrXceFd/
IATob0nbN8THJdpUyeXWg9GwK0yUXyKyWI8SX1PjGnjG1QMA+nr/B7AslelG6u/Y9qJE3+vrvgJ/
3QVtZbHfwj2efk6BsMvBAYCORM6dILzvrJTsKc21eVia1oycPYB1DzZdxm7MFhrBwkju4JRCkP2E
isbzYEu5JmIvot8YRaagiNsPokJmBdtnC+J3Q9OEVmBwe03UgBpsn51QCpwaVfSJ/ORwa9AH+pgi
BTFPL+WUfPZQhOf6N0ZiVjS/yFjOJgiLLyyHcLCOHeOY/h8VPh7IsC1Ez4kx4H5ROQ7XfFog8Exc
0uFH3RJBuOpeLFcl9tbC109zM/Bf3tbMMF9ae6WZUcvxjhFebvgjof39o3H8KXr5HR+KTabt2eJj
E2D8S8k39VNLpa/qSEMPDBlpFDT+PuLgU3IH54j0eAHxQOqtwqE+zdjizzY8y5+MniM7GLrafwD5
lpGG2OLsQkmYr5m2qkVmepLxcYSe/FMgl1R5ZjSq+jQyuJkUNs/knbAWdP7/okSFQPsVDnwGs4ji
0+HT/h3CMxnbgeBExtUGxZnMRoMSirXRSf1PRicK903jZGXExrPdj62bjh68nNbwBlSyOvJEOJhE
uCvH0W+aerb+fo5vRuuNmF9+Jd1IPYanGRmZzi2IfMr8yURCSlaoBHacN81QjuzLzwdeW2/QQzuR
yfmn0Y+W1DNhrZPIjxsugiD8ukIHfFsZGpnzqgmDO5QsWK9MK56cIaJ9Brll8AwOCLAq/Uxar20g
AeDGX/tM5SaF4tyNadJzcQPzicluXpMrU3tcn9w1sSuG4eDw0iNHIf1aYQ6H75o7rhj8cNK2S4RS
mXjxgrSE/0sOKQE2IRFiQv5PQKc+nI41qADn/Pi2cCiGzS0CkKTH2ZTdzfEwGDV7pnBSXSkqb5EO
ScXvto3XDUR69JiYyWOC6yZMDSTNLQRlEOyIp9hogqivP4hFMLVhVk0AVkJ1PhFQM5DwPQEfLVRE
/F6npQCxy5vza+ZPuUdSNsnZE0eSc1MKZMmqqMM4LK8WFy4XUc5fX6opSprZOkrmLb/PTrM9Pgd6
fB9A8nahnaQDi2BRDreZU3nLR0vTqfZNHAoVBa6nZxLTVrAvlEe7WblsTP0maI0Sgq4vTT1laGRV
EPy8MX2vbKPWjuoKKTvsvdcYLo7qw0QjWymDwEV1QlmyyBfFyndm4nqlseNsf5Q6d/xHUFzdNymX
M5n4dGmwyUOhfeiT4OfSuU0AGj/Lu/CIRdYoVz1hUqBD0H6/gzkYqAJ8ZBvjR76nH4jJN02ci+Sm
ULx6tfeaRfGv03cjo/mmVwLuHFl45agU7TTMxb5Eq6tz/R8fWhBagNbx+2I9pq+y/3J7OmqxILnX
Lg4MB09s8qWK7qaYQwxx8p5aU3sRTH9c6SX/2grLkRHTuJ8vobAR27mtHMvsHvQhXkaitLUj7DNq
2sYtKPMc65A7wh/t1vihvRmLVp46JmbeYFxcLiF/mQnm3ThRwtsTwaXBiTYwm9h//lH8v7g5Ir+G
Mix800CPf1qHcy+6aMlLDZQrr2hIn4Q+pZX+fgyWrawTgk2u4W9CDJm19F9JVa+zLNyKZ072wztj
ZtWt3YCaTryHWFlni5BHBIO4MwvqRO3UWRHTMKzl64tXNsxnJWCpkAdrZsANkgMfw61K3c2bj3n8
82/mq+7n4dTueASEgL35i4sInMtC5WYDGFF4MN2oF2OSXHv/5wK36gkEnBTr2zinlgeIzGP2+vJq
V80wjFGxda8M9tfsQ62N6FZn0GNil1D2wIOP8xubTMsA39wSzd8dF6FgIXZupmNwJM/Z0yaFfaik
YeYRUMDsi2jV5PA5OUfPAl0Or371vyijy92skmUoOZ/P6b2Dx5U5LyH1BHeN5jAbuKgqv1FsYotA
Kp6+URY+sENX2txBCH0X4/UWpQbT6kpT8AYqiCt/oO0DQ9a8vBktILn2boAC3kfDRauUGQp2AHXc
ddn7SrqmV/GreB71q1BFSaq+FiPK3dhiX8Qog+icXaw3In8EVZhzytKngtkdTnGG0DfQ6cwjViEl
kbtnolxqZ/c5NA2HDbBAJNrPH9vOckk7k6XGyM9iJbZuAq6wWL+CM7IpYqafY0p3wp8Eylx8Vf+I
79bTl//UDBbu9IK/w8gbtwlK9Du9OdrYgHfCwMjjJGfZKUD74mqD3dXtMZxqDTXoiYZ8YAzrkfj0
Z3SwaZuNSlFKbepId084MWu21ujtW9bUr7od1Cv77U3B0uf8XbmvGOZuwq4ORLgsbHqDYjLFVAAC
xmJBbH2WkN8/mVeHm4AaOoPznoE0TEUVCY+qc34vc9aCIs81rI0L/caZNlEQjiR008/uxOHbRzzl
Xf0EW5JTpDzHNYyupA8oTfSqfiIMx7tHRVoi4SurF45JNLd2W4axyHYEcXVa5uJZIMKSRZK4WAcH
RGRoHhG3zH8YlePM9GTIdWkXLEV6IXFgzJmBCTVF1QzxTspS201me7g3+hkaruByk+NTcmwfCK0t
1ld7jJHmPuuPS1NrwFtSjBegJPJv0O8YvTLDWMuV5zlSo0mb9rdNeoS2gXrJ5jY3G5Ohmlz1fL91
ltbAXgPtxFbDLxtLc3ZRTANg9HTGMxujs6yEP+n2gVAQTaNxoeQMlXarWmgNdNxzykY4DgNcgQux
ZbfAZEARs8Rf3qABc9/i101ScgXFs4j8mDzwoWcA79xoT7TwZ1vEkNr/I1r3l8gwKMDATTa5OK1i
smnnzJV0PdXhIanQRSxc/cPsm/oUbCkmgMgjBg58v6y9pBCGqxgyH5s0k60xrUFK98Uvu6QNgdZ5
/Zhu/pikV4NF0RoxNtj9rngO4xlvmR3dMDRYjn/hjmVMkqcmXZB+CEJxoHm1xIpMIQ42/UtmydI1
eliirWXrx5AjQgmA9YtFI4GEy12rX57nn+kS318Azk3/xMpaM3snOBIKzE5ShaCIXfmqoApkrl/4
o0mH9/DPRlwA+k35mBxXSO0m8mjzF7I/82PHtHRcb95c/2gsA5TYhC3jhhUGXlF6mc05v9YsYlBT
HZqeQ6TIeKcebvOOQ8bVYXq7kr7ahEgKOGF9BsnNG9k3RXs5424ZDt8LTbf27/5tlabO4ab5Aqc6
oRIJ/cEsTbZlhL2Ac8Uf7LzF90EId9f1s07nLiQPXhl+7qKnYX04vsxIRfxnntjI+P4nAOy8L/zr
ZLYt9A+sseT5FabwxdQBbnkMBq3HJUztxbosYwl9d5DsmIqCWCVnYYnJhDr5Pv4EZ80dK4FtIpkD
TDLRyq1NCJmQ8qaC4sugtbgnxCauXlCVGpwWmobSrzoUV8MIZNwwBhKKyL/fBpnoWzEcpBCbw70x
a64y1FOhI+Ku6vn7rYRyFw5uFHyG8r+MIuIX2a8wSXgcXd7UVz/875GWYX4Pje+tw1M6Uk6WzjSB
2+Qf7DNLzx/Kc4VoQW5e6G2NPcDy/cqibaNSgCnvu8JOXC7wgrMjDAPrBhYoMBdAn33S2mCZGlw6
MGymjgQqBvqw+JWsDqSimbqp3t4qoR5l0kR3wsUVfj5LxelA5gSLzWgufj74EQANW90DRjUAG4fy
5uncWeL+ECy6ZL3OYoBVu9pj19QiESqNg3U/fcIb/hS/Mp3ZlgoiKYhPVpto9VE/L5tDTqeSWLBU
X1akrd6WcqEtIu+u5XkGSkdL32N3MmB3WO+yz8ZXzSSE+SFTTjqGKdGpHG4PeTzAIyVMEH3Bcg9b
35w8SEd1fKH67h3u3BKcMI6+lnWRScIUUaywliRG3mdoHv5/9raxXqn/nH7CgKRnJh1mexUbke3c
QhyFU2Q+3IdR/SOqu8PUU228Ak5uUswGweKSm4Zs/Fsz0cM0Q8GNwhKQLqryYlcMzq5YPqikQxQP
czaHs3rvWLLcQ3WfxRk+/+vINg8OH2jV0Xxyt3V2GhlRpcd3LoeNhQvZ7xs4EZhV/ptzRe7YvbWu
KJj06nPrI4KMZypAe9uAe2u9pibnDYFqU+utVJPZTZkXdbP1rqoTFH4OyttqSQDWNd/iykKQ4Lky
2rH8o9fh0/CT/WhNJjqHmwZhJsyMCJl5/j1idWobFE2RTgTzd6ioJV6ukmflXJy4Dd18sctivq6S
o/WrGDiPMcqKCvalYFKNysECEiI14Cc0rdzFIGUEC+WLc/bM7lWvzey3SMK71auUA7SnjlycQpk5
ZPHLJAfITnLfTCh2LlO9SS6OEyDRMB4niXQu/SEpyi4thq8g+7w8eAIlWah/kTkVkU7u8mTOMpYj
/HKkMF7YZM+8U46jTEsC0bC+Fab7ECrtmRVVHs5q38izJgfWPgBYq5Ln/EGxcS4/957NfuHPTBJ2
6CyxbAJzg8JDZWA+HnXtie26shPLkBCGO46OF3QYvdxzvSiimCsRucSCpG62U1pW7kO+jG2y8/T+
i9Gal6Q+wtKfKpPoO68wBL3vSYamWiPlbcVs4Q0atIT9PExCuBbGFu+YTD6qUi+idSR2EQjeh9EP
4ouszIXifQe7QO6TLjYxj1lNY4/t0WEtBPzwo/NrqX2UlVTwQpAiJOQpBmA4yNCYp5FLDO0Uuoex
0kOi7RSFhFMb0OE64xoJhPyhMVD5ILRtfstSgW/sPoF7wZE/afwx1qs1w5v2WQ2YCdrYxPVBrrz2
2MZzLMvo2SaybeLGQT18DHG4jazcHXotrjnhYgPdmDmd/0pIb28Exp8WOT7fjHraSfhqBV2RMK1e
oY14iKNlNrMgXhu5wd1HbjPS/FOy05MP/EtKsK+RhlbvvXtG7RL6zqQmnJKt+0eScfs7XTvbNyzP
tmjtWpwjw71bg1E2Y1s9qHdMyg5obYtBd00AVm+DSsmaQqSpPtswpuVNfIgZptSR+UEwh5Y3Cxxm
VIHbkPMz61YBq77oMORpOLV1u/x6iF2p8ltqE79/IfjmUpC2xfzgI/oYVGMTId9gOtWM2j30AMew
xRimM8cBkMAt9m/Ib/EGSh/kW7lehO9jH62Y+3KWuoynD/7Y4zPxm5fiqXvtIgoL/43NSWbk/erH
4qhuUCATD1UNPFYcKzpROzl0bJ9xjEqfIuptSTnPJ1r2HifmrHkJ5w4l0Ph5Xeh3aT1LkpGKAcS3
o2rhsovbZd2DUJzWNYAhHHzWBq1YXf+WvfUYUyRF6IkKrNiEcDgzzsl1zextDOXley8JFbMND14t
LhbxBTRxJ+CTCVE+rGtEqaIiQg44jeL7Ga2vgc8Ih6t0OkFtavqknxYZZ6kpeWjDwQx2L5mRCJpd
JU59km//lcYrf8ugS7RQJE5VpR9tNfhlyrul2352arEwFp4fr1IKtq25OSrjRiuCTZH+wBDoVNuO
IjefgHNUBNMhOCwOptITJU/kfdngozwKPRM5q/K9YbPc/U6HbeLUvSy74bT5TR/gR7ELAJdLPB7T
O6aYSaXr6P1c802iegHc74pi6xqBBp3zW4xAgL6a5JYER4/WxWprXrEwcbD4XVhJciIsC0IKc9qD
MQZV2gA9FRR5/Y7/q5yx7O0vtAaFwtsw4QwhTBbJveKOkDyO+0duvCkhoh1rAvbsqu1L41kOpyIv
C8uM7OYpm8BMRMHbLnMy4tuQJaZfd+H3f2eyvRw/RnavhRAm36bTfwe0x43SrXYba2oR/JsDY2no
pXo3E8ghh1AG6x9nEbz2WnMNbjmV6PjzPBrq6cLZHCymQcprEssR7Z8pQYbxhXE4Fb2mEo5RDZFK
/gQasfb0cRdJKLnM7JpyKBU2nlGe19Yau6q8MLX1GrbX6BzgDmUCfPOg4Z+7rGS01zYMJgiocESQ
aAn5TEOwdiAgmtZQld08hCUZwlf22rPDrS0JckZq9dV/woEjHcmQzHynuOWQgbx3J2ltCxOzjeGB
/JswXDqZn/RSZc1tEhsBCORPp1hHG8l4opdIf5F9IaOOp9Fq/txBlxmHXqgV2fNJx4jWr0zvOfTz
cfow1sYMUPqm6bO9gk8mwLLDuMKqd80J52/ZCTsmV6czRNVJVgHWJU8t9i/3lhkW7/dZkW5JtjJY
Vo0ZyOq3im5MKuFMpw4I0Ug+KdqhAdfytnMA38gSOZJRhUJBefDHIkNfNdn5we0FY3/Twhl8WreD
SG8jx6mAHcJ1Rrn1duUxLkHibZ+HbvRDVnuZZlv7F2RKShXxgb0l4JHdoZDo8wn8FU3NcLXY+qcM
VMCnO+94g08jWgvd1ma8sSYjpJ/Nas95vpxMr0op0cyFyzx/cgD/cHLqN+nKqlFu0WCqLT4f9tUu
YISuFA9KgNxV5GhiTv7Lg/5AK1HvntmV6tlVnSUuVXzoOp4VZnOpHlaME03JmrpeTFrzR+nkwxKp
qLKz3L/zeTL1Fl+m7qoQygN+XRJ177z9TYQfZdKbMvg+N2K/XUXpMOdUPUpON8HT7mcmFIR9MqjZ
2e6IogOvkpRZ6LM1/PkNvmp54OzMOThlnfw/mpZc3fjHRN4xZO/aQBaGw8hnsaLTkh/OPF23colY
wH/NLVcnUJ/883TuLHz2InfSjR/raVOWVGGFcd0pyXZA7ljAXcMqLFG8cKhWzYPHLUGcgIBM8Ug/
VfPwWw5TVlgvCiZDRZrZ+FDVTeaVk1zEhsJh/JQn7vABJgd8d7Fi0OwZAKxH4dyk+PQ5/Tg1/Up5
Yk2MJtZM2JYDw/a0UiDXijOQGkRZWh0R6hCOeOr8G/kRzuqLwR3oMCbDXhOU3yXJB6TJT/mfZsrS
Q/Py47HAgrxi4olJShyh49qkjBndGOpCTa57asApMFlhF3V8v1m3f+SruhdDd81ec7B9f7L/O545
+KTapH1i6uWHs7R9l+/y2NStBjX9jRSVVoXbNEmHrq2t4oXMKPdxGSA8SrzkePQlbSNKpaFu7JNn
3P2R5IdQGHN13MjBIT+Fx4b/UCZUrKxehekabI1O3OsnOFst960z9INxcHqXFg/D2S1FealLAHlI
HMVrLi73dlF1cVV8owys7WxbnPzwHqFVhZ1cFvHELCDwiPc1v5Laz5i7WRzZ62aZMA51j3hrHDik
Ip4nvPoiUObtNo0DidZ3YQe35dj0Nl5+XUz9gc8YK6zIp+OeHPvK+rtzvF+POIQrXhQR6YU5MiIE
rBbdcnVw3J2KNAq1HAL6Bjzxwo5S2dSg4wkO8cz1oOI15Kvs/V75ZTWnJrksIU61VH4ED29rlu/u
QvzGmjQxYNqVfC3Gi/OUjNugOiebrbN5USHpS9zzuwl3Tz1oCSDIx/BrJ6Z1FIvXR6bK3khxlUNb
yicU6lCMIlV7aPHhRfe+dhFJQ6KlmZ5c8oc0znzvneJb1Vn5+4ErfihZrSkVBmMM8iJdnkjI7zBq
A9MlPgXMIZqPukWJZa+MogMcjdMYmWht3uHwJ6xhMQrQ16JeXZ7syghKoxNeDiAmWtniYii94+Tc
QppAQ69804A2DXCLTQtmTGrpHFtt71s+oZt0H01+SacsOWoibaXPj2HNEK6Ff79IZPcZbMMS7Pih
oPg+rrU2qBrU4Ipa7x38Cy9lgcUUsu5ksDCxhK19d+Fyfhek4exenaIdTGpKvA/xBN4fqHxk4Oi1
KUaZlbDfsEgOPFot8kOiCT2cuK8Gu6XwTYlelce3K+16Siurld5iyUP1Ryjcn7qerTq95stDz4Qz
SDszzsofb5yIVLQ3v3eFt4FFmvphZVoop6vKW1oi/vGG3vp2+vwdE1lgbe+TZv4BopFyv+A8GR+M
yc9LZG61bIf1PND2eLJ1BHhOyuxX14n27vUDLIEEIMntH9SGTvOil3ZRtax5jE8dr2q5WFy3XlYD
hFciQOmRRoeXzay2DwGChZkjsggtLLsggNo2uP/Rq78NLxU9I/vNlY0ccpmlLHRCqEfXswFyO9jL
yUlir2hnsEbfeJkvocjEF34UhMJO9AIZ11AbEm1z4TkS+ApDkxAW5pG2m6m3jF0dlqJt3JSH+cvC
NWWE2qK1uK/mrj1slOMCi7hUbVv4dbWP3tngRmQpUwRSPaG6IsytddlxKW99mP5mCMgEJLXT4jot
h7fMM1Aj3Vm5llSvRpwfzl540Qr8aC9hs7EziuczyHWPlBX63QHW28mTUaIQhyEWJvb32yb63NgJ
jxmiu9daypPC5/jBmEGrKwkwUqWJI1jAYicBhB95e6vSTMXvJWFKCYg7ehOy6Pygafzh1sU+1QjD
mlJeCbkjL4i0Nbidvuf3WTnIyg38+8zqXLTBbCBDUdco8A4xMaGOCrOybQpFH0R6hxlRzPxrajoM
NOYfmkBQoOsKDAlOIBeHlNkFuf9cSTYF4nj9lu0CbKqE1XAht/9OnvEZmhOAMTXkLoCZRwD834kx
7eIjj3HXNNu+Q9QxUiyeJBaZw/8JWeoTP0uqbT32aN9fU9gwWhwT0+N2kQGyzivCk5tk/nvsa7Yp
oZPHfSj7TDG9AX5AkeZEUo0ZF4aTZ2JlPKuO/mRnc9vbbKrihwpTLia4vWKn20jGanbgIH6eGBUl
7JMGCNAYJITDocvjiWUmco4hc4j4tnGQkh4JYsrQn5NtRhmaIqmlyDWKaXzyKXVkWJpHbdodyULV
CC/U3QRdZuvJNZEbklS0aZWVDGPUaYVbd9kb/BsuUQ5ZbzDFk3ZCHpvzoh4TPQas9NE1yZYNZnDf
WfzBXlejvNF9sTbiFaReIM/gtQmZAUokruRb9kdyKn2ctul2dN03GE9WlKxr3yIbbylARaWjnhDa
t+yAPGubcPS7bNSA8vaoVBLh6wJ47I9CiDgm5+rR/USVVH6mf4AwPKdRS91woLJIe5he7a4Y9N2r
Po+VxZxx740cLCBl0b0RGjpwjZeUdrB5TlyK5XHX2gwSHtKmN3a2kNjpM3fMb5WMSFEgSguGPWBq
9gf4bXdlSgoNLahIGTDsKwldGcGm1JYsx4QwdEdtMaMrO1pvVaECTfSzoH+maC1S0FPunjflXUsu
IKLjS+1yeRjiBHulw9dbCdz7udmwtz9PQdX77BmIG/V4W2tvzmobW0epzBdHJs17o93NxBPdsTM6
uns8zdbolOWgTZMrZrklBPQrVIkAzJRoFYbZ7+prajqF2uw/xj0m7INsl1G0lHcOh3Jg1hzW3vlj
qFptsdeo5Dz2wQCR+50kdLrmSFnLSCO77fDiEg5oLtmYTfr9AYEA5mQTEQEUv959027D53obYWAY
LEbFN7nYYKjaiHYfpf42kzVm9FaO3SbRBpxjFXNbL6LDUmoru76qaI6ed/F9v/tl5suDe5ykEAZn
gD37o1UdwbUVWT5jJXhnQAqKn+9qXzakzKbfqKki+gpAHrGD18v9GRe7g6r/9AsZRWkjDBP0CFRA
u2FRu02vnz5VbvQNqpCyBHG9uc4dSXJQFL/xnMdlHPrJ7DhnEjz9awOKj/FFHBwU+LTIS+v+RZiC
m//DMTDa9+tbILtuh4wolxAryOxkldQVgI45gpzQmGnxX5xAz+umqRqt6QhpjIryMDGuoxx2LKeu
zEZlw/+3w6AOhRGbdLzepO3bHIieYrCF6U0BxfDSaYugsek+j2KWM+Rl+yzBY3Lp4OAsYMadOOfN
uqYLYdzUWVHGEi5ZxRKbmveAE1PewRpaKrQKOhORkGTtWqcZ6BYiaQ4XiYzvBLctgKDTKprs8MEJ
jEBs2Z0Y6WspDyCPI2d1vbSVjp9y0b64A9rMvB223vwCarAl453woyviLnENNKoxJMZIZoCB/HPQ
rOFmiFh7TNnZQR18Eetk7eG+b5YTilbVOUuiOOpbs4Yiv864zamZw9sy+b0n4gjbSk3EG/2KBqZC
kOu4e46/yyQCMvIWJD10WPJBQRkNVD9Gk1lxDTexn+rlvU6ahzNPNSMTnJA17XH44KhbIZXJYPRT
zjM8MyNZmCK2kanmhC6h9g6pSF3fYhC/kpuPMl94BJ1DGE/9wKzOhUbr1eh1Zdd6wrRSoYlXUK3N
zjPzNGSbhTe9ftyvigjFJtMvWy1vCPHXCZgckBNkT9cdcg7hiuuOU+rqBVH7YDRtF59u2zbrdRbX
/VRVZ//HKfLpbMP+i5K43JdV1Wk8dWIAB5bdEa3SRzRLqvsBgMwZ8SG/IrO4O71bVHcp8fESAzPp
DIWmZWnnNJeLJ2UwCugPCg8tBQmkwJxMSyV5ZsPG9SlNJXqavdQ7G1Y1AVSBR85yBuQ+NbVYbyks
vBIJG1R7m3Ukmmu/wWmWVs25Rc6YYyzfWKtscB+vhfq/bMcv8gO3Od/qLJQCEhxiQha0S8AqSn+g
VgDD0VkqhNYF/51Eu9iicb/xyxN9bR+WkjJodzBAnmDelwks52DQKhucHi/D1iEY8BrMX1PhPGvx
taJly0o+/3KioRPADK0v3Xj0gZMgikTBnVX/8iQZZPwfcg1mitHzyJ4EwtWZcgE6FOA0IDhRfIcs
GXR0gc2PW1pG9hdEUYZ01RJ+7/txzo4xZtb3J4Nl63KgQc/qCa0DSPKOSoa5fJwAfqNry0tGm7a2
m5fakjW1+x2RZZIk7vxpqLjuiQyR9P/G71PQvg4w3+QOUZry3q/K7WjoY5uwC8D9M8VJNvu3v1KO
lBgheFzupibDeyaftHB+9mqcjQEQPeu5G4EEmrxQLdrfpI810y2Oki5jjILj9lQea2MGy7I1Sm1s
/Tn7gqXNozdCEQlWUZEtV4grgNQIccYVRPgXzx5+JIRsU7PhMvNROX0XR4HXF+Kejapd4A3Detbd
qjqt/pkNyqwKDl0q4bb4n5AweFcW/yAHFECvZ3RVTJbB1qAF2CeD+bXko7SUJskgpprCtqMKJ7AX
aSkReZnmBcOC6zZrq7zudtOPF+MRxXPDyLdVx3sp04dGD1XbEr1Fc5pPp/IlRA2gocl0KlGHZY+G
jaS3FNlSJ0CWY1CIJGssuePmCwJfOxUDZZmOTo9N6Jv9+ura76Gc8VfCYIAe/Y5X3gUnIQyx2sl6
vXFLXsU06A0eCzX8CEjc8hJK5SqUt6LTTahPF5rNECoStdPEzxKUpct153vnJPRyv3kcDtcZ8nCH
Ghx5n5RLztj/KI/QwIVd6i6csYiQiSz+uzjscnqhiNbrta1Tyyn7ubMZfjnASYWoFK2KPEpCgwg7
xC1IIiDMWyjYlhBkKD3hARkbz60545lnlkCWSOYtHnMAdLDTL09Q2Qh+Jf9CgN2PyP1b02NUVyGa
DGu3PQESqI37TMqWoCbw5rs8O1TLp4tev2ebiNOpbTSPHYcPSZGgL0Sp/Qiea8byLvVrKj3cLgeC
7ot1nEw7577KLYuu1w6HqEigz34bYlEk4iPz/z+f3UtW3whnlF9j0RhXC71TmeV6ubZtqXDNN94A
3ExFKpefejZwgtckM6EZq5JwxFB7kP5Dq7P1QsOFv7r5gQQBdfNvg7t0SIXfJ+Hidy5T0VZdMJnz
bUcQlMtQ0qCqb15ZV76tFZJtUWON3tNvuJYaAYQZ/4m5513/0GRh3JN/F3T1Ucv3wt7SugvUtbsj
zcpGnsi0H0ZYFVktmcY6jZ1XGBkzoR1OZcrz9GA5Q72rSOs6li2MLwLbE7LeQwZIZ/kQi/6qLzRU
SyXL/xnB5cVdciTg/gh9W4aFeYew8KgUHjLQWC3+ix5jh64JFPAWSz/gt3JJDbVjRtt6/uYosXmY
GA40mDXRVUia14FfBlH2tuMQtot7qJfr02MxVaLZkOSyIv/PfAm6gntCZmNnmGh6dYPQVctORVXA
vwMir2hiYID9bq06QfgOxIDo6TKauhaY79s5PdfdGHqy+ogd3BK1lxJnJ4mkIvs6KYRgIReIgqir
gOqik6WqcEK0Jv4YIzziUX5FgEwooafamDDqp4WFZEcET4ioRTOXGIhbE/h5vOlWJfy8B8PwprFO
zfqwN1axbxPwy2s2ehr2GETPa+i9jnrtwWfB1ncdQt5G/aRPPnD+Z9BcsNe6IAel6VjdMh6a6FCA
TceZ8zoBMJdsJ9XTLi1If936Iwd7V72Q64f3vc9PPoZXwkm36+S+zFJemLxbUJMFsT5Ap0qTisj4
ziPMeekC5e3H1SY76qna/YB+2gIT8mZxhQOh1UE7iRpGK4ASYYB8G2FJoEOTuUDnRpDcO4j5Uxe7
svU7yBs2b6gScEYDBF+hv074t/N0kAdq7vjY/80TaOTkFzJkIB1MLiM/p8lHBGiywBn6A+X9KLfG
HzfggXQ11Jv0nqlUF8NplZs0WebGGRg92UfD4/4IUWwe36+gi0WutDxck8Pplffsk87/wenYzmsT
uRLWH8VCmIW1UOlPhmBAIc0ylWgc3f9YHjUovrdwewZTw+3KWDJDLS9rJUaMSM3lo1YnImEvQwFy
uIZlrPd6pVVfp986lA1ZBEV8aofcXJd+PoHb1iCi2aX8Us1fombgFLitPsI+93Dd5Pmu13/uG0Qw
yC3y/JG0xaW1r+lzAE8TKbEww5wMGoJkNVDlbl8n8heMFg+Ib40+QAw6ecG/2bOgFkeyA2Irk5PC
SyAku7lHvHvJ2/HoU927O9aDAbhN9BWvs+fXbxWjZLza3ByeMcGM5NvGHzfwuorrEC39ofUNdjwx
0MNKVrL15xgUGmXv9qRqcJ/0n0WsrXowtoFmSJQ2Hlk2AG9+VeKDPCZa5fyt25p+tHidJkoj7CgZ
K9LT5lXr/Xxnb1pygrPjNOPp5xopaRI7wjG9Xxyu/zc0NloX7Jy5PTMBFORkMt4P9QQoOKHAY89w
YAIFF80QN/ChcuWDZyxirpM4RzNgSGOH/KMFDufga7Ap12ZBaVS0+6gPJmAH7ZdqwgdLeykiyYV5
1LcT9XlMTlTPI7AIQfEnkea7BIWYgoP2wnxGxZUfaJQsfFikylv9h55v9an82AxrmNV3iNki0fEO
x49+sm0cXkHypdNECqngItSyQlhuqWcgOTA7vfj6iRBzq6qo7arfY33/mzckZn2KEeJASqrFqZUb
M07fH4gVf+zB6c9SDdb6heiEMuZNYiD30EQFzfFRYI+jmEKL0EfDn3jX/Iy6xV3eLod4qCSID0/X
MPrgBTfLov/f0/kIiKhOPMerA5KiiELeCY4mnNvcBub73J/gBEhiOZxs0rJejRFX/jdjiTmC8qHp
Bl9rjQh62QT7sg6N9gbHhc3QKusT47d31wk4yRkCNcJnaVycl9Cn9LGwVoH/FmWMaVAFy6oPLTCd
DeGVWPKwidUXD617gF9vStYrMzgryOdD+YdKjvIEG1Hdk5SErIwJqoQ6/hssCtVmjPDgiL27woav
aJIjkexbMp4GvAjurPOiZEPidaBkUwZppiP4T7YGakZbfQ16DIhUICRHwy1VbiwSKbKPtbWfQw+j
cf9G5/l0d+Fchkc3/1/7VrI0RxxDA0EUg5DX4nHi9Vt87jr9beYN2sQSov64++UPpGLIcsGwex4D
1XcZcfDd1sADBLT5i6tgp4i26tDo+eUskajHCnLO1HhR961/vx91jBZ8Rt/5z29A94dtYYTSuKlA
/OKW5CQDMM65yzdsTKG7a1Y04qhqioVxPpYHbxADIXAtwkEvAWjpUlW+AQKOxCQ+A6obQ0p+69Pz
s3AXBqfygfMorLuzkxBV/ixDnfutav+GS6/pjNQ9MVXDQ/B28zQxHejlMFKDCAQJHHhmah5/HRaV
du5cfx1YhVwwvDIrWFVFyLX9/gs1jM6+dhgn1wgcgW0JedmbWsMNRiqJk0Di4uU0jc4B7mjOmUax
XTH9KyznWuCrydQFUTho7qAkQ/K30Un5DVmeUFFIDq7rLppBT5VW/eoXp0oBYma0B9fcocAToQnL
XjCtX50lzlOQ3n4pDm+zcucabYovKt/Vi/mz6QzGD9/qZLuZXv1QDRZR6CS3/ErUhC1XEq3F2wx2
KsG0aMjZ8iKoyWKu6+BybgaDB1X3Iok9hg9KgJrYIUaZ3wn8eKRyFk22lDvNjxu0vqgsZR4GBz+v
sZlHaa75oSSnv2FqmUCjHtSxvu0mY2QZehwpAki/9bSuqVHL6FMAhZqBunRdedGfAadEuZyHrZYB
TGQQ2SuiCNGfZZnak2kRORBfb+7zJleIiZ3P3b+xuwh4mDI5O0ONhPjTu7QVMfJ7GwsJp1jAprQM
SR7Z+Ml9o2dHRhHVhURf31QKS6t/rWzJ2naZjTD6CoUjsf0ETJj0JfkaUXGesi1RF/ojDzdlRDzO
O99cNRWSLkULtHTohTaa4EY41MVIIGoLGMRTcgmCCOi9s5o/motkTEq723x2ENsgoBcL5Mo9Loec
QdWn4wAqxaEWxeUvAtYT4NKV+3H/58IR
`protect end_protected

