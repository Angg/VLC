

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
cQDd3XIPPlgRDhqULvYHvwCty2ZrVwzfefmANvx1dZIylIMC/SlAcj88wfYJOEUSOPC1U3p3rRJH
cF/G+RPdfg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
hcwXqOGXIKp1yMXglvtwKNDD2csTguI/218BbAfP1Qe5YaY7t7J14bh3PN4/sY8v5SUfs5PPhYYF
AVoQ7+Y8KyIAkFOjVjl8Q3cizlaMAyaX6UCc4wmflvCCOjy7mkT0VJKPELyiFH5OE1gTiKu4NfqY
cLpas2QiSAVn/xZw83g=


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JJiSVarYWytdLFzHp3wkrD5+jxEb6zxCxwIxMuHES7X4vO/81ppoMZmSB67P59pBX5Chyu0EswKT
bCRha6XDZljqkcBWrrqj3cLRE57UCaEr1RVpDNBMw7hjNrwCb9eTELEwb3X0mZPKBqVrRNroBMN5
Mb9o7SPJ2GKhIDEDF5Q=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
x9rjekK3vn0E248BFQkRU8rm2REs1XV6NiMfscimCVnt3moe1QOgVJzTLPCcPYvThLcZJXwVyFUX
J1k2lVxuHKaC3FNNToKLX7girUcVANbS6jS2AjaAfdpYmQXF6epSjXy+KOWM7AfrGv2r7XNIcV6T
P4He3ZDDIABlWanBaDiVD6NYtB9SspFXaifjJ2faT9Et8gWmYJogYQ4BjXl960BUcxWS5faBudWm
MidcfsfVFpzH5bJ9L+thBkdIh/P3Rjr9ssCSzEagp+1l0DsZGX583KqMaKiaZiIsR+KyQ8Hrld0H
vh5k+kh3k9z7ewkJNwM0LCpa2Y0qGSJOxIauzg==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bMGW+/GNxe7XIGxZQsPwYg9NhBUySelE4d3DawPwcsMkcAefxMJ1JdlslSvSp+VjxIobQhkauqfs
plGQEEjRkhr+3m8iz7uiwT6s+TtBZQ509t+m12KAHsziCshi0m7JEPgqnpkYUxS5ZbKQCRgudms0
J1TIIpIIdBJiHjiJWPFKhl2FSk46olekE0MQ/LvS36IE6UC8sP+H2MLZpAxpzqHuZ9TNFvVcyr9C
pc7viw1i7pElJF0USsLWRjDFrkLdXdznJwKPhjmDvq2WWhH0UZss4B7FZEDrUrjB/HO8EjVy2Hj1
fpw3eQ84VC/StEBHWhh2/ovbE1xsoAsXeBE8Tw==


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pp8HZNaXt/evJqKzoiOa8A1cmkUh/1mQf/2Vkpam3N+hCoX7wAAqGU/zZVMPYP16RpMjeC5zeSin
YvUeVcdgv5x+e+joKUcjexTi2LwQorDqPIl0bCwYx4LccUexnWG6I9/pSM85Q6QNP03F3dTfZ+nY
q8I48HLVTNxhG5xD9+JTBp8D7rjXe9TJGi+hVikOsYhuY2PrwtvuAWhuicAfJnsIE23LJrp0i1cL
6oyVsfKsx+68L6qOWniySUGZ5yDe5zDF3WoQ1oHIZl8/tfnTJcGPsIRyeo3fpk/6/w5zWnz1pHuZ
HvGPaU9zIF3KNoE/3qKTDNhAcVbvP4+ohJfKxw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4784)
`protect data_block
wUfRnjv38VcmBjA968UBahqkltWRmbPeTWWTSlt72sLelnW3V7xV4xzVgbiB2fyVeyAwmrmJSUob
FnTUT56dF4p+TVJggSRyz3qqQucsokZAD8woKxyqNQ3yKKBkIQaEJDPKeOEzd4w9aFlLal0xOxj/
i3KIV1rUZWeZESqGTzH3iM/Am5BBPgLqzRD15LNsMdrJJ00gm5IPbTYEDnmr0wmDvbs7QHdbaIKm
9Y5hU+/mvyICvEViLIbFjHP1arz/pQ9ip8WwnbxpME5+TwBDs9gRBtqVH/p5QZSscmD2P1UVp1if
xYxAO0hOcQlRfB3tNodA7vSNFk4g+ZyCa7mQVmb5FnpUUW9ZyvxHLyncDtm8UsMN1bCtBaOww+dc
CrSA3VnW30/7qDanKUGR5kljdWUPKSCXzRnlPn9o/1dDOpk2JFUGAfgWczKsPP5v2XEsWzfjhZmu
xRT+02ksFTgNJlPBYfiXhH75WaiyHPHYfMpNC8jhc92633bNxC36vpTGCG7oARP/p4m7XJzj+4l9
LVNwfcXJ82VW45NH8SIj4Ed1KqeLTh78zxpFTBydM7UohNaQOG243mNBZ0vwt3R5WXs2NN6KnXH/
xIMVgIk5+qgEt1CErD5WwTNNgMaXt9EvOKc9wYIyoQETNq28OoVphxnpsOcKrqqUCPtfcepwImY1
vhtfrpA2zFysjZXlTruyM1IyBFQvTSI2QqfWBYTo9SCZLF4mGCI7DmuKjemZlY4dqslxyFw0BW3L
n7qhXJWXKVsK1FyZNnxURy6nh0Sm/mDrsJZzIL4cPRzDUvhkWRZ2VQU94P7cJIe2aM9SkgavQw9s
ddjGcRAUNoneqKytBK91JKiGlxG4Oe1x3Ef4zmswRii9ZjTmsIcJaY0Vxc2vjKLPxbmoABVFqUB0
jEIUjJ5eUwOYR5MvplIr1owrxg72dVCNX+MzZjJtb9nksgWbzynEjjnv1R0HsAAHjQLsEK8piag3
wHGu0ER3KEooZTBEH1efEb2tGixC61sIL+vb5g19ZK5FsJisjYBUhgNT/Pq/VUwJdoQyiE54BMRt
uUikaaLGsDDbL6wd+aow4XSRcGrk921MzgHyPp58FgHYxay4F+pYjSyZ1/qjNMbfNU/WrRVnsvjh
grtejDKazbufnypxJC07yMIxn+h+BtuIG1IaczHJLJRUliQmzozBwoPIKm//0NNOxlVYSWDqYMJJ
UPKDIYpa6WIK6yWI3VGXbQh5dwIYK4CbOXcgY77tG95FRLFfJgRCgyTxUXBpS+bD46DcI+q84YJR
pmQ8M0g7Qo8QdBTfoEAQheUERV/fXKw2nl7g7rbhp8T5BjLBizbNMdvWV05zT01vq/cRRnPQ6czm
E3j61DbGBH50ottIC/WYP0yOgME0mY/cJurzWv8NWvJIHkhqdD2sBj/L/hhmaJCqygD4XSKC+YOj
OYOJ5xonCh4NMN8fKOzdc6VfsEQq/4jLfdfFarvcSVxT2EVzdTt99CFdd23B21YDvK+Wm/+lfUSX
XLaCN/3NGZvNiPNP4W/CkSu3tmTIHsOsrfKRxUm4VNgJFvwVySH6AbftfB2GL6mt26nyc4SuMz5K
xgIkyPYpuCv0KZp+kBjhbPPcSk1aoiwinl5pr1VigR2mjxjL+BwWKJpCh99fYdLCwAsix2mWxux9
SueMWLYB6tlFc3kfdin2EoZw6t1kQos5BJ52dsTv7UFkJiGYVteM9gmLOLXPwRydtWs3iAB04BIn
rfbApxHx7ut0A3Y95LsH4GhTLauipPrya9nc3sEZZ5OfVZ5dhWy4xMU1cxPnJK232VarYh1bLeaj
e1nrCEbuEu9kloE2+ZE6eJQ6imgAaZU3ReXq7t+OgkkP218PSEyZdFUaqVtKDBnjJ0j+X0rJhz/u
ShWrLguJ2hnoakPFZgMEM6+PiJ8KY1t5XyoOWQZIX/flnc6gEx2ZQw79WFWFEBWLUv6b/FNkqgxy
8hkEjBOQus7jdsWwdZLUfcYNU+IcRQbQGbTprz62/ENlBdtEehWFx0D90YOXIIm3d0qYWRyqaP0M
9SYwmE4LdIbFs3vj8s/7AjJP/JlurwxJAKjfOA8bVKLvPrfdTixnCL/O73kOpI9LbYZ/+Gvv3Qvp
GUDQ322bVDaYdrYm6LcI7wvuyYOO65NSXAnAkXo1q5Bc/0yuipcNsGITQwmZY6LSsuAhs0naJObS
TZW0Lyr9X5V11aLI5GtOjKmyqC7KZysayCHrr8yFgkCUfVgq+JNLO5D8jciXsUmXvHxftmZ4GEuY
sdSEJAB6sCerAel2if9SzXsI2aGufMIwUTAck6nqB+ufOu8ih204oLZustjeWyzFnPSxR7km19oM
MEATYPPJ4B0RQJ1c89Hgf8TKPmLZc4Gs+TkBglR/QXXPCwxJ/Tum8NZhCHuBv1vrxgmznBA2fUEd
RjhGTpvF70X3DB1+ufzI7Fl9ZizJ0UDfhKBXCb2Vu3g6QQh6aT0TBVnQkqaUWMbuJFbO9y1b6GwW
ewvCr6dVYSe03+tAa3YavYNuKV2MPyvaeVrlbVY+zbISYzyUYcOKtUZwSZvtq22L16CYRNEol+uF
du5MqU1RBw3goRhI64GaaNNm30fnFlh4oizdjpgbiBZ13QMvv+RWeTkFCkFuAmGJlYUxQmxaUbkF
e61lYsQT21Qx7BI0E/4RyNPKfqw+GYNYNmjqdYfchhitoWYxNuP73d5v5g9Udb9Ei1uYVsAd54Pl
8HMBOHH3ldhVeOmfyqfuS0pYfnSo4YqUVFKo60wyA+8g+XuPFSaMC61Z7XR7Dp5U4u8vG15PVK9L
IoTU9izaSAxOahQRG1wiCW+5OvtwAv5DVPKRDt5K5QNDfjsimngt0lCky7iB9TTOKNjPvlgkHRtK
kZssL2N30R8MZX61Cr2fjeAvf/REQobAtdeVDxfwd54px7BW02vUScXJA1sV6v4RZPn1hzYQ1nAw
uJ+m5T9l5QDAI7s3LKHgBNJdpf85UpRNnTdw3jKKYvY/SMH09JbtQzI1GZLBpjPGFdU1Qryut9Bm
O0TE9QajpERxPoM0fRwdkfM3fOhAnSUgH1Q7JguxmudrBHcUGGJ5QBs7zLZjTgqxRxcSoavVC8q7
AZGN9TaPSbIONHuvqR9QKuM/OZ9lwrAcjYRXQ9RFGoPCHDrnDTGlFZ0a3rzxZZD1X7SgkURQaspB
LhDmT/WFMUxGM2BdoUs3qsf284aquzY4z4jfRasihklpJSHezYj5e9ouvR7CCYJl1a8GhSNG9elK
YiE1/VdFsqkL5cgTArGTqNvk6qJHFN+99WFx1gYK3AtcQ1VYfVgeEfnWVFosOVa0VedFFrhjCT1H
F0LnN5o9g0QaHvPyUtI+GQcD74MwwygaI1HmKwLgIWJJEbByeAM+l1S2rLIs4CPNhsf/RIJWqbcY
wUG9zCFgUIxMQ8JpVCtBwP/HgTbtvZjmYlhU+lVYb/3++LrZnF/i9TRO8AykkRqAlkDLC28XWnbh
/Q3ru/0xuTqhtdHwi/0wlMKHPjGYEPA4dPtc7SeIt3cb39PvSmTiiEjabCq9icUEbIurE1GRQ5A1
72pEhgB7/WJGXKhCf1Dzg2m8TPXq27yAWIha3ipW5mcTozwJwpNa1R34KSzIv8DWzuSm0C1Z+0ff
D7pZ+Tqy3rr3d+ykPB8IsntbJ1CYcDNeIGZgZmhjbLR/gkEwmD7x8E3JySunzCo8UFShtObcxU9a
5M0omFo2ES1Nxdfo62ABCvVNpdfKhIGG7hQCH/Zs3s4sYyPQbmveQYVcVBeg60kS80A23kS496xT
gv3YEwA751i2RNyd77hhgKjM1HZYxvSJAhMEz2F7Sl3TkWnMe+4atcjM8QPZYlU27r1L23Huqo24
JbpTR2TWhxcRtlOLEbj5YRVuv9/xfj31I0oRTRKl7NM/iO4OQVRBL630TI+rxuqKnmHgSuNuCLLx
BTwPQ9DxD/KJcq5maPDnWhpzAOXtrunQEewfiqaZVwUJR1bX6DgFfiCiucta1j8/zUrC2qL+YOaM
j26GALwL3NwRmnhNjh0v6RPoqURATkZR4XW8vMd1aS4X6zkiJAQ9YYlqc9tRhovfB9nP6r4FSqzd
/S3eSnDRW5DJBTb/LXjsbpN1XVbCIWDphLv+4/I9ftOEbu6EDCZU0bUXW9c5fmBs+PjoOrYZo7V1
veRNsXalzuFU4Crc9S5se201L0w9CMDDZhODOYRbRXhKZGyWjgKlXMD2HFrsafGQ18Ln+774eJWF
X3DAUxxv94inM+CyI8YX3PcWWJVlL2x50Nucmx28jtA1wKvneJopIZIyXxpWL9nm8+Nss0KK4JcI
6z9ZGG4L+RSAw+qsmzEltJNhdiMmAf1590DloHi5zEjGqChSNaiDjzN9CNZnuzGTrSjmTiOHQ6M+
SVVLVOHQeTJQxRwjuZwY4Q3fBb7dO/aHk+8ae/SyXAXO3VAHyuQx8annzbpV3CoGj8ublx55aRoN
vRxRJ1hB4ieToH4MKZhJrLgol7v3rDsFH/QI83/wau0ZoEdvtdERr2orubsO4gKcjWCZJi1TNr9N
TncCIt4NJUa7irOrHSo/CmXiGpy7HoirWUD8dCicQqnQYV8UtxLXo4dIwM6y9ttl1zp8a2MWemrE
IAcKUC51nhw9CrEfdPCurGhR8Crk3nG6KVC7OJFNXPqgn2Fe8YVawh2JMN4eyisTW6DVwbDg18dr
AI6Le9FYNZbrtZIgqOGRLUY6ywDGj6eftAypyCYqE+OX/qqpm/Z26zSQC2bcGDi7dFz2vj85l3AN
c8U6tl54QrvWhOmo73HMhQoFM11L0qFpRDlPqHul9Jij1cIcY6jM4w5TX1NSXjJlSbs8e6BGbe2W
IOWVEK3q3W4+hJ5vBViC1RFqopEW031ka726r6wdnxTJM+Wfj8y6wz2BuFTcibK/KCLZekGeVEm0
Di4c40dHqozCmZTvOr8NX8AVtQ9XWr/P4mO0u2gir1sr3bHEME4WT70txkFKo1LMSOcbXa1IAPXc
JJD/+DliGB6UvXB+pllxv5sMAvhVOl6op7rszaxO3ijL9ddpjr2JVemSA4HsxtsdLLOJjYTihRA6
fsXYzzON9J8C8VtB20FBd4nLplOyOWg7iDudVC/4hc0EHF37hzWyeRCyxDj9Y2MpM4LBT/noSpEv
5J5/yC/gG22HpX+EL8EVSbx4BpXLgva1eedoCAwmxnHuZhnuvxGV2FYbURJpLvtyb1XVmESlcM/4
nkTixwTrH93bcF99NGWgU1xZortNP6j68DJXh8DeWJiOnpnV/s1VTvMCoscuPNNERlhzw+LoNxEq
W9AeWb8K0tv+nIgMYGizuSMoMTkwkJyv/Hravqk3F81neEF2GzIDLiBDE57BkHQpKCf9CWIUrTUh
ml071BO1h2/Hd4T2sdSDujjP0bPI+E6e8bWMo2QXS3A3NH+QZPy8bWH6pZHcTUl24wQUrgjRpYzU
6H2ymPaVQ4oY64Y83+6Wxk0M+VQFOGndrXCpR5ig1+B1v0YOImYfEmbBdkSE+jGP/yZph6qDXYZg
J5DFaKoqMfXRkhHohSyxZOs47j+/zghe27X6TjFso328vJplzdIIbROeljSTqGmSEN7UehxWSQO+
mPL4EETh8fIiP6/BwP+gLAq6ap/06iIdBDeBfjPi+K8tGmG0BxMUIyPyM4sUUApj8az4eR72EGrv
533w4hcdbyLZhDtD988jKnHXlSDQ02AxDzIG1J0lDX5aqONtFSqlNi9+hBvZpi2r6RuucKz8AKN0
u4mI6ozfQfNP7TF/7UZyDXiI3HQ/csfS6/8KRIeitWCU8OomI7dluOTCfV9vT4MJdvHUDqhrE8Lh
Ov5n/jTVtxDxhW0VtcDcRtVgJ6QXpekReagHrO8OKSIUlPZSHNmdTV9w9v0lE30EFKrEN2rpo3wW
XHZBcwdn+c0aSiqKRU3eGVMkAldUz++9FwcOxlFO3yjoM429WQfJkHW274hZmDQNoSTMJ7C06W8b
ESF5CwUNkDgzuiHdnpJT33ueFJfav7nBz5c8GPmIy0CoFJ6fToAHhjB7JRRGxOG2OLJLF9otJbtb
kPScipCIusvruoOnFUh8aPMZjO54sFdsUse6Tf2pL+nfiVdZ1DRPAG94rYTLMxKCLZep1IkdAAaX
aS/oLm8AU/xZ6jl+hLyaELsnm+0zb2TVmsK7THityuWzQNAHVySERp/lbqnTy1TxMb/Sc7Vr0qDu
1mYobMHtctiyRRTtD8KghwPgwWkoLat4t2Gev1P3m4SD9EEVfXwWwtf7J+JJ/k881NiQrTGeKpmG
pw8Ljl0wDralPThjcdin77mqk3GkC63McC89RA4d8iCIDoZeT4CNcRGoDY+N29QXIUP7Sew=
`protect end_protected

