

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
gD7l84kB+WAh1ATog3H36h0/cMgn9QL5jGe9p9PjvP7N+FJAVvGVlrxcgBw6dZaWDNZqNANQuRFv
ZSE8fsSCFg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
YQUcxim/tlzHeVlJ7otHN7u41KO3Yg5DFb1yF4GCsbXGLtUvWNlkFjY+UPIlgYImR4Zo4dTHJQ+j
3BaUNSUOqAVzT9CfyUelv2YD2ZTfAtzIe1Mboyb3+StKnuzxnZmIhVPiZlowdW5lQ1r7BjDPOsge
ztxOfUTbvYcTUE1ABIE=


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
eu4MFD/NMz3pssr62VCh1XDd9mthYydX9VaOq3lWUwHi5/7e5dl2SAWHtYwTnBgGPY+jCcMycJhy
WSlkhQxVj5BsMm2aAItwXFvH2mSbjlPggtI0/+DNGQ4x8LQSFLTDYnnQbBrHlJymsS+/asMkXACD
SJ2tF8LF5tMhAlMPZZ0=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rNAzbNlIFUMjdhvgzZ2FokzvR4AuFtV+1AHGDKa9QgeBsZ1e0Fom48uKbJ9iakvqUoUcKKAvRzeY
OBkbx9P7Imx0gvIgzFsgiVw23cBYWOhbhSqVb7mef9aKx8yeF8T48n7gKldUkwBHIPeqaayRI9/Q
HCZO+k2+HCjRZE6L/Gzd+IOdEVUFOg3NtWFPk2JFkfZkxs8X7Vg/xxtvH7uvp+/EbVyiMbnwDT/p
NSqOyA+rJwBJYD3xRIPTFDI83XJLCF+1i4E8hyu7Y0F9MtjKugqEHwAG+JK3jde00nzNNaeLVUQ1
OfFMZJpkk0Cg66d2cvJY/G11oPkmvTq/JZ4+5g==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
apuTRT8aJu0TR7Ciy6ONiGK4AT7TUEiokS4gFf1g+kDg6PdKk9VRun4HKszIadRtahjPQo0of9uS
yvu3GS4EQo+Y+T116wnAIXnZSa8EQaEsDkziOI+rCvXv8IgaPYN8Cq0aRlASFL7IHOWNI49V0c0A
FIG/+5U7ZyNQFCVwuE4gCgK/pA6apm5kY4FGJft/EdZ5YAbR/nCTzK4P53+XsKHrtGfw+/MthFWz
tI0OtloKqc7laKZWKOVFqWq8Qmq7UL6utFODtxEQqzczH+q+Gw4rkUyOosIY+cbB67hX+GlmXXEF
jMwvUcen9t6c+wiH6rmBDcUIiuUHHz6q+jCwJQ==


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dfDj35aI8y6zqcW/IHFxmCDw2mpyex25qQAUnsL+tIRxivv/85PqpCOrf3b7NWnwUKMrsxtw+JBY
mtlPsVxQKR1gn6VkaHwbEgwxXXxFe71Z+1nWQhfF8Nt55jGvq1joWKMrurSV7Mo+HkvHMSszXj3v
8ElD0S6sN91oml0nObejOhxzHf0ybK+sGag+CFA7aBr4k4rYglf7AzOYrPl3nNoCkyrFDQFa46/w
SXJm/os7zUHbsDI5GGUH3BU+NktHZV6GK3iyhtHTwrMgDtpGk6vKHMKULM1Gjv9g1/jp9Ao4cUhr
bCVOXM1v2e8A3564rmh3if78zTzCKamPRAB5Ig==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5312)
`protect data_block
8aYWzANd6lzwkn5rzdbEEv/7IoVdR+5Ka6Hknc2V48xH+1U0v4A8e1bOMpS4qv1+n+oEEj48RCmf
MO0sTHGqk2MV9a4MA8Ts/EnkQqMA9WffvqC8LTVF84zGo0tXv6jpIAZZsyyv9Re8K+qdh4SjkYdh
Icvjpc4EyxazqgWmnpe5ZHzepMFNsXITyjLltDnIJV44arG1D0sa2X0LwYsVqfoHMNNzmVQ/wtT5
ZEFYhHS+HlVkbWdvO54Zj+trKwBbqvxmymCctvD5URUVup2RCU+lNNmJTRnGB+Soz1aRumpeaJAx
PYOwqPb2yeEWAH/9W/TCB00tnl0OKb6gR82Nmk5S+FwM/Nv5KgmmkNXg2+ZWSiw4brOR9eQ4fSih
DDn7FXXvvmgXsf4/TrnLpbJ/XPCK+uKJLiYRZIhLVFgKHbDXM7iwfOwMTQAhuNNbBEM40XSVLJvp
N0PSdtn5607h9qgEWuw8hffVBO9TbSO/Y11p0kb4J71obYk+m2CGz6lGSeRE6ijJnSZcCKncKA22
3XAoh/sw8atzmr2UCRCFmF5H7PMacGEwDpvcwrQhbcGoIv6DYP/wjr8e1BnRuo3mAf6Wx0If9cHX
EEWGC5uw5cujxKMMqRrWlBRIG+kFkYAO+2FPPq3sIFRVqDC6desAI5TP6474fivp5R7kWSmYRtyQ
z0LAfXrGqKtRHttQdu6k2h+F0CQrmW3YUy+aLuu1FgB9YikhqbP+yKZsm8c6KhruJcf6kHkW9YB8
E7px8lNmzhJaCb9Zn2T9fJLQ/33FmM5J9hhyjh+LluWJaNRMoxmEYNXe8s5Auv4aH5I4tFhdFq/b
cftca6u0vECiQakWN0v/qnPZKMxMuAINZSEjV+S8X124zFU2tAtYyGjqgPp+UCC35RsqhYV3UyG7
xHh0JSmjbR12o9L/TrS1fuBi9ED+M9b/R7g/IzXXHGHcSH7oWtKQYHMMRDt3TOVsybLVyZsLlFKM
7oNvcrCcjlhMB3NtnEMjW4V58CnEKqA4gWkn4Mxxws5e7MJBLo71qeSbMWahmpxnuxxPUjlhMR8r
CN2oE8Ck5/sFhlylQvKSGW58hLdiGkfCaNrHFOKy7YiPFg+bclgVw3fytT4c9EVVhOx6To/8TsIB
y/kSKq+GUiRChY/08dwrEQ9sOPbC3gIGxevvjbgELjR/H06cRaeADS97UB6ZUWUdyFxjbr1bToAr
+XPltmMrgARWIE6/wl0fwSl+Tl4kQ2g7WZIRxCa+GfVG8me3cmvszoTF9S3C/8+kbmrw8iOmPTA9
Dg37TpZYF9VYdUqRs41vIIMCNShWmc2hRLXNtAb1/KyWuhBicxex7zw4FY4bxVUyWzr0hAH4FaWY
Hl4HjHlQAZ4BuPN15hz77pFH8TDAtWMnRKXulzTDDh+evYlBs5mUWQxN5sXtEsLmHfSRJgJFEUrv
FB344kZbOdwNEFyxqEm7hjwIvh4P5KuXDz/Lu2//YbY63vAJowRKeMGJEomjgQksK0J+uWo3Y5Ch
KUElJQj2IocEJE9FkWgw4UNTV8CaVsIprNrZQ/l2Huuoc5WnUGKO5TLe7xAIGLDxV2BKO1nrw9+3
bjiIdOmrbDMtSvDjbyr3vB88rMhERi/MbuhfFqd2jfVMrYd0thvkKiCFwguDjIsv7cDs5eO2OJK8
5KdJBnxwMphkFY8nDrPpwN9rQI5ND0NpZWtQaCsx5cF9MADUZ708q1ZGKPgsI79/gTL5o7NGIHPp
OdbT07ADWasHcPGNpbLBJ7B/KoRulmOKWWYEFQf8TN+dbmgD/Akeqzy2xFWIWs/IMgKGp8gI7mVu
EvW66+1AhxR3Gutdgk3NgSTYQlcakunFCf7H91dDgST+ddIn+AlU4L6zDuza7LhNpoYyIaSN4neB
CBSopekrkTrWRXDnrT/G90ZssQEpfvamYXkcNHNfM4Qca3uLKrGjK5HQZ1SdfIUf58sd+Jkk8wZH
Dkc6TGZ2nWjgM8sils6EaYruv3msELQNraclhibAElDKeO3+rOrUXHVkZF0V6Je9J7EY8bDum+PX
SHgFXy1x0DFJV7J+e8QSI/gwmDEcDgVkBI1d+uJc0SP50vkAu2QOxBcyvaUzX8u7Pr1nCdMchX0V
okwajltvPyNldNFmzDi/AXANusjG7z/+D/Cml9tvG6WpjHM/pHBa3bIOiS6g7umG3RGWFLFeOUyv
ZEDpymCPHXn4wTV/azZpIyKR5vTQj194K9yv2kC8hZtL9roKqOORMrFYb2s9iSOp76WsZr2bKT6u
8o04HqoSSWCznB4EP70XjRrwaHLzBWBgT178RIlrxa6Rx4bOitfK//O/o8Q4x6wmbo5vWWCOjiFR
lncZufFOTTMHqvJ5/y14Sf1q3XpT1w5MyS10wV+RzeU8Qjzwwl6mFyIIURYmFqSD+DkS0cjJDZ8r
nVybhv4ESRs+t8yy6mloOqh7bBMGSWxtQCdEYQWm/Pwxen/dte1D3pewS2j75ia9CV/Ta42YAW1S
QfGimVsOQxuRK797mrL2kmesN7M0GMRV0U1jkOPQFBC2TMBTq5ZE2rGu01Eg9EUVrIxzKf526eaz
0p8X0OFffNTztnZNb3Yespu+mPR6T+we1Sbk2USfwjs0L6+/2iVYeZJUmuBnljB8J6CAM8JrUhI5
bpt5S49F+uY7a4hhSy67d9KX+IuDv5C2BAfag9oTlEFuU2JRamjXR7umUe00fq4dlzcjzlUj4eIv
wjku85qFGZKuKOxTItGcb4q3la+kgC93X0zN/+rbx+cTgtENXQkSRU4dhEU/k1E4G5PXChY44nLA
UXR8UXRfh6Y09MnR1XoitRcEWTooq+MGqJTA8WPMViFYQK/kwMbohCIUyIn2jaIppSccQsz3RHWp
IxXPgXbPw2IATPa87KQ1nSBhhr2MCEAGHfC2AQIZoJHly9sopI3NKvfgHZbF7gn+Q+UtXjWSz+9k
lbuWdjjpKC787zofZra+aQNGIVqb9HPbNVQsOvexmoCstQKzPbm0CP5eSJ6w5xcHm2kZTy3lP/h9
n4MVzP8Muw7w37hjPZlphkgaNLsSpU06ObuHTEhgQshq1/bgWn7BYyra3RnAtwtcg8WaT80AgI53
xCqkwUl61TNK7KpLfMijbh05J4EuoDJv8MzVuo69ircTIggl52UsrpRi7CFmQ6nJVJwi3WEk8IbK
SMdDKa8Mg7aSVIn2NwWRj9tMKTXd0LGamy0kNoKVJdEvKcK0jcBvPRG3V/Yyb9MyLXctu2Z/HowB
93O/1X6j4lxoTw6/Hp6HHvegjZtkXfCNa0rr/IWaSARmqLWtgzwBAfSqGP8bo3pSLBARPj1d/vpf
yTI8gEQ3BQWUKIJ/D7DNfFYGdhiXMKrMadcE3NpuWiHrBmB4VnR66POsNA/LvfCv+gTHpocXreWy
fZ4MeePIorRgqCkRsnNdSfIeseZsxZyZ/7JCD5o1Z8IhR703d9PVbjVLYVIPK8AClR3fdqfh+OuE
9xzaJJUYCCfF++n1xL5YJfEr46ZZKL2VEMwf6H5LnElPmtMEMHK05Lb8/bSgglBvr4nDrgXBPaI8
80Ea4nhq+n3MwIhueaUZUHi6vsiAs9bwt7LNobgCcx3eXG0MD/uvY8jRvgi4NA0FimRFLJoh0z8V
9jxmnYVtMRHrFcCY5QMgl6hLoahqmQljO2HpLLnCP7YJGKDCSw5BmBqHenrYjPySOMOovn/HTzoo
OhJ3HGFIeYmzO2b09LhMtHkBKCMnSC7FMwMj2XaTe+Wun7niN/c4TVmE7Q6rN/MoStQlsUFELUsz
fc119QOQQr1aHR5A0655EvC4i8QOdxZUCRsT1/yuSjp8v+V2CPf4AiJYULYnc4JilkY0L63Re86q
rt6nsev+nxE9vtpPPSjy2fDuCnk1lvn+EFNT748ZC3TDfjry82jNs3VwXaiuyic8F5r+56zaI0tG
9OZcoNX9B27Nw9VD8isll2mKO819/+0vrkwXT97FL5TSB576lm1BhA+NF9hzdmt6cqyhTe+PNSpL
FaUYU5mdp9gbhspGXBCA688eS01XFY7LFEDkwq+lA8mcr4GwllcAaQkYTZaa4wzwmgnIhEH+b45c
JsMkY5eMgWpK3FuiJoJNh/opmSysqgzrJX+dg+silQH3pOcLqjzHjK8OTsb4wZTIutuQLJQ4+PwY
VxlxAFhvHQ/KveIZg3naZiG9begejHiP0CTdO2Zf2milZhNNXwmnP+Gz/4WqVAYIyeTxGvHxyqFW
OPouoc2rZpuBYXm8iYLi6jFatWu7foZdCn+H2LNA5ycGDJe9v+1WzbMvS+5hj47/ovNYmd4e7tYX
CuwSNuM7YiUPFkF1AZTX8NUsQFupZBBJffrToSVZw+5vbyexFlLdncqBpHibUrH0CJLQfeFZbouR
drSvJ1Tk02acGGazERhB7QW0MiulN3WoUCGV+aMhjdk13m2XQZMEgzXRadC93xoI8WB4Zt/8hX6w
O439hGcJuSKrBD57efXF2mUfKelql0txQZkQz+7rkAYosMhZFpgpKWO2yjQskmksPak7Fpj9Z7jh
TRXHwWaSlsKSqnw89LCXXmN49y6FAuXdardhPa3xa+2BpC/dCjuiQjuhejUgpOSuVNdy53QyYrZo
kzQSh9NJ31rN1BbbOTNjamrSIuz1/C+RwGhexHhRBVfA/yAtdjZiJPE1hXnHIx+H3OTB/9gSdz0c
IoTMixIY9KnDpQepLfRoyl9lh5FkRdUe638gPSyqku/fwSnKal2xxR9ksLe5bKDkeUNpnqLe6QcO
rWCQ8udf3PjdVkUQXcS/oFQyngCa4+O5l1bbbNmdkCxpjaSR3dyPuZS1xSbrVq0bVzBvPuhoWagK
HUzfRWSLWbmi0Kdx3iZTMK0BrxK1R1IYf6qAQeMF3rLKntWIfBPFAT8/pMsc3c6whF7BklwGLws5
BxL3jPhReUY4RP8Dwgr2IkN5nSPpx64NNpkXmsworCxA2thIQ7Kxmgs45iJs94hTiDSduzx6/OmD
FydfHjun/0D6fD/Kx6/kkVUlvTP3K0sla+4OFoRGrF/JAziGmyC8Ru54rU8rseEoniN8kYiUWctt
6f8nbMSbpgf71ivf7fyWCBeLjpvN8+VLWQKYhfSHmkKJhjY5N0VpCJiIdo3+K7uKqAk4pE6RCNVd
xmpv0yBNNvoPMW1cIJ77Lyl1RTDx0Dz/NTfTHM8O/bLVIpuxiZ0EtQt9M+yoY4h4qfk+L+c7MGTb
P9YVVWp3hE3/aYR4all6xXyGBi8DxB8rlNQGhzMJx85eeXpximRm3gyiFWb5Yb71XjJ92eXDNzfb
6YEI6tXHj+oMASYtOx6/utsCUaU31a7KXodHSSadS45Jz0FUb0I1U+VIxexlwZa0wPGfWrFzWcHs
2+yep/DBEBo3wIW5hgGsTbZpppEq0Z6prbhgC4kMr+VejU8kTzchoumEWk5vvEgqxuUhV4ma/F+Q
KuvTO+9IBcVV4UGRfJhMY4WoUVoNBg41eVJuq+RpFiBJTdtq1uKMrkB/fmqKIbx2DeBmHDTWISec
gPmFFECwnBSpTJEy28goDZRwViBeWr9P+mYYf3cKdW3tqfLm8XDE91cXAjHrFr2Y7SvO17Vns/r/
E7T/s99eKDc0osr0fo6dznBIDMSV4BT6RLZriRK5HGc2b1oa6ixLQNOv/+/ikkBiVBAbY5azTDCh
x+BaNInW4ddFfEQspjCqlwXitQmEQK4yLt/9ixtyZGy3aeHvV+JjSI2mDp/cFIjql6+ON6MxqSWu
GcdTi+A5C3v8RRlXaptcjySw3YdrOKaKfw4iNZpJ7PQWEAh79JDAYm0ukEhL5scvJMRLyxOjhEWZ
vT5IEDkE6493elHRPJhWhbrAkMfK6J9KmXYkdBYUxu6PSUPZObGsBw6HTlNkrjQcNP14kzERzxu4
sSXF4DH7TttefxjAFZD9t/0Tp6ghjRQOpg8AGhybcgnYT0YBKEP4o6u/BI4Ve/HDfSl7nlWlJljn
DaSgn2eAr06JpQmRe8ulepFbyM9skHIAAjDPlHehL7Cgfzy/3IPP3uM5SmKBZCkTv/umeEFD3UyV
WbTWsDqGlkzJHFrvk4VCvsphIN/mp8rozfHRyn4QUUqxeOj34gp7OJ9VfD5X0WttgLfuWEHrrJQw
+k3xWNzjY1EB+m+dhr9DNTYkCQ44WZfhA5TTYr/xUPqIVI0gKrQvIUVQ3mNJ370xq/PqR0Sbf1jg
RkMSBUHq1bkBRsubkgEwT7rCknGbWsFjWJgLzoo5vyh5X7m/M+ALmiaIUZO+5DRkcruoGyNs6uQ0
KopLxpdWKJBo1l+G55QV6wBGKbqFez2556YHQpwRaCwzIxBddhCRusIPDT9Dmu5F1VpT/6Xx1ZkH
sGNKRB/bEsAKBzU4B7zhKqBzyCWF+69Vf3MmvDPvKD+2P6iALsOx1CEddAcDn2mSa+Do0I+sW7J/
NEoaHufYjw9eEpeef2N5flvG9w6tOky8SqpyGcVVB6NTwvtApvE7RMhIgSCvAK7dEiZDzfT+JRGj
W8/j0fDzZTur13ZaRlAU2y6jcLSObUuYij3Bns0XTSigMF9CaHzN3FumMzezmPVV5B+fCwZrMzUE
iTGZqqUr9ZTHmkSgzGqMNSLnLJF7708imrg9YT4cwhx5pW4YbNjA8ouJJ559aMgEf91NKCc7YF6R
e9tdUThJ2JaYtxTw82V+reDJCBvKzahYGxX/hI2H3Jy/uE38EM3qZwB10ozB+2G7cjoAeVTC3O+I
Ji5LcVKreWqeMOY9mLuiimcCSdvzC/OeEoFWa95/edpHhgxB9dmrenn5vtZSY6WEWgIPwYoBjXbT
0HCW42CPpSdnXWO04iMR5Snlq6JLYYnr9ZlRBKDWjk3wNYL83klP+ly2YKt3+i1mCHSelL7svgk3
V9MUamFZVwzpFBxL15arDD4k8m95tighHRHSzsuCnchasHDfLWXaZMZMV4qBR1vcr3iS63kh84wq
W618Rib2C7GNeqz0Jvn96PUL3/I6a6C8CywDtPBBKd0cnGT6GnQAXel+ZgK4px8+tbM47B8Enxb/
SqfGozBx2cW9TDQ=
`protect end_protected

