

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
DNkSCrKrSZZGZ7V5MEC0Sa+FIa8Gkzj+o/6NpxIyEzT1r0pebmEX5gzn4ZglnkddvJ8/1f149Df6
ndMlnzvmbA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
W3TEk2OoVAEcY9sACr8qvdTXcz4KMrr0wBUYfTJiYRXEKj2r9L+Frj5vlPoRfXyR8BXMuNIvntP/
hRtRCfRyewmxrXe1oHJIEkJM8D6eCjNM+zuIptS0mt/AsnOv+MMQLDkTVqLaJNUJXubQtL+dhzzd
RD9SIj/ZMKv/oOZJjHU=


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
2wWKJdgoqz3pSafJq9a67M/dd2FxPncTZHCUPF6InCTgFQ7MOQlzLhplRl102JxCos5KzhVt25al
HkjLSxu9PHw1ru871OGKgua1sS3EafdVjGCdT5iL+6+M9XT4bQzC8cVlky4YWr6qOy3G0Bl3zGGA
4U8j4LRDtMi3U1kOYa0=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Kxq1/5UngNEJdxzilglpkl2MQX9t6W7lRQYEeATFLTlsFzdBmcbPaM4E6/H6jb3hTjltHCzXXzJL
yu68g88g81H7vk+zIgG9p+bAH5mVTWnGpTcQ9Nq3V+BFNfatOquArwL5wvfxgYh4qmnz5LLzO8Vn
ZipCR6RyJHvmX3LECK4ZGhdOjgqLTbHPcqhN/bNhl+BKCVrOY8qTWY6WSJt2I/pR5hbR+Gxpp0v1
fzycz6IA1AnyF4dzdl4sorgs97DN/Rwyy5DX+iGMZoJWJSj+jKc0DU3coqqjuApwjmgaPZEOIkHt
fmd8I93zHpUVO+LU0o2VXdLy/rhhX4k5zyqLIQ==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
MMro34sbMT/dSBUUDKeWGj+AS/ioQgVbGWAXG3XMUY+tNHQekxt+oKRBWcwquBl3sw3SJLbR1Rnx
TjJ2MDDzEH5uCz1vX7jZaQbMCFAU3K7MBn40b87mRKYgK2nBkQ63tKhSjfklMsYEEkc5/qUdspSU
GIdrS3bVjN2jI60HeE4r8Ae7725zNCxoNO7hmmiicY8i9qwR3Jx3RLeEISc/SwYIBg0patrQcspa
o2nUblqCyHtuSc/DkaBV68tb1S3LDYROKbnkmBVtPajoK0FwTW/5ES6DuetOb0ujYKX5ZJWNoJr0
DsAiVxbKY23jSFr7uskYGQGx1K/crFks1SMEuQ==


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
DXzksdzpRyBvPJAO8RW4ZhlhoWO1yMLSwz3BzpxXSQKUFJz2DfYgIojvnKP+h4SEWOeOMQNr+agZ
sZh5CyJzK3n38AYVr+qSmIrSxy//25NZBDMRWM06jl3lxtySkqX1u9lRJvnZzDG3hVY4BI+zv+3m
Uys3/UlD6y6GV0iCZqSqOjNMRk77t+OnDh3CxzRxxv1qIqIA3AkY4LV1fP5qMWjFIYo2yfPwXZ31
leLLHOibckzEYHfpK61VUGsfYsK/Omf6e+sJIk4DfwW7z+qr59Fv/xjUYitqPxa99lpT0eMUcAbZ
NbV6OJqwWXo35ZdTdYOXEUb32x+tBF6ayvy+zg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 909824)
`protect data_block
6+ZT5N3qKm2jjMRLDB8m3BfdAMBEEytgnZZR8O4mtdLSJxKisxz/uWtrRzYFuTZrhAkzHhFmqeP8
EEh+jOHE05d9FFNjp5bLgNx3sqj5znEN8dyKaonNowzk0xVdxVFhUFucrn1Ud5yAa6lPxsEyp4iM
6ZChDwK+VnDc521U7AwWey4NaOJVXEdptnT+hQ74HnrFpaYv95sbjy9Ops1eeFaB+GHLdrOY8Ake
2+kJMZh0yyZxFc1gLKUyWD4R2Jg/dymA6W1vbBaeYSr7QZA/lumoyyLncbFI5tu6U+SgJ/cc77dD
rLFn8XrCUSVHqSAaeUadvJr5Dff4q/QtHdGjNX4pzZUPa3z6bSLAQm81JGwh0iE6reY0dV2goQIA
h6V+OrTAAxVY5SfkHOilxcvQ4mWJQG7xu99FMYC4ZSc+oSDGd9esowVJaenKkJFRZwYI3Dye2Rm1
GoDWpvLyeb2EzaRhExMHPgGhC3WRYkIzJ5AFxGQgYAe6upxm1j1uGwmx2RaqOw0t79Y7ZTBtmYLy
1JYkPxjUGZGkiOAMJOZhUy9Y24+tA3WSrDkHqwmsmzH/n0uM1luBhBnrT+1gFAEMlsZCsapbZdZY
LRScUYh18uPy31KmOM9eVvYkV6kWuRXWs2uKlgnDWygULzFABMX7V6S3s9e1E2ZloDeRLQQ0/ASG
HS2Lu6h/eRCN/Mc/SWic8AxBTnohzi/C9ohatPTZBvE/wmgxoiIIy7Tr+7efquQ7Go94cqAX5ZhN
vdIV8OR4E3PL/4Jwzc7SPj0v19d1PMxt6Xxv7490tm/FI3yIEN30PXAIcSCqSMZ6a033nG0s7VqX
Bqjo3nMGCRpfMq69r4pey+j49fYnEz5RyguIIc1UImH8WKya+8KQM54b4yhrGzr3aXQl2o5ImSuN
/AdYfSsbi4zBdX1qWif0xfOyCuT6nOJ7SA+uijDgSfmxo0wOKF4/0YYGt6fDz8DVIxaO9jmrCDvQ
C8vZUE3xrBxWwCE+WE3ZjuYdHLNpVAWwlU62B83UUAjwnWtC0vM+s7j9JekceW9o+/UJzE7ynZJD
6InjTzrsaCxHCVpQ9o9mICLzgTMIrFvYOT8mQQo/t70XG5+MvQVtkLUZKXksd+SjXo3Mp6x1GGrx
DnhPtDRVVp1Tii/qCJhI1vROLXJNHfz/LRWKHIs9vIb1nbz4SeHuF9RfT5xhvy3EpyM+Hf5Rb9e6
71BRWJzFdb3//i6heASoFoxYHkix7lp//Q1/5ove7y0PY4ZCgA59jAPzlvYSE5/4Taf1mmSXlkyM
zCzIzFO1bRWKWOzFZNWG+Dv7RYH2ei//bs33cK7FqFRi+5b/qKJz7cYj9THOqx8S7SLEufH6gxyM
aFBhl+thv5AO2ymyLcUt/FDK8OrKoY7B2bRnN9jN2CL4ApcdqKh2PA1Yz0/Sltg0VzBPOTA+oV8k
MOwA2FoLrNy/OP5oPE4WkTs3+cZ0u/v3jbAJn4PXFZHYqe5VQ3kuyELv8Uqf8eYmv6bCHtn8PxRu
ih8qWA7a4cuTBkPfcmIGCgFYqtqqr8uir0A0NZAaUYIYqmwtZVeNhS42puXzPBQEUhy17/jeX/Cr
m+irfrCgVkgpA0wwsS0d4qqfOLvCMBfqb41GXlMzxscEBhVFb9ZBwBMw6/1Vbf/3Xtkk+YMUOEgg
SOJ4swapgaayiq+hWfV5s29amXE2SXR6tEcs4fu/0ZLe/SnQyb8hhE2WwB6okIgyIuLzG7PKP0l3
wCVKRKgk67lwW6Dqu2QNvcjegSJy+CGXykMt7NE4IurdBA0zz3eMoZ7NFuFHbJygIbHb4fM/rLDX
4LM9s1RZ5NWfJzmgliOolY3IdOvupsASOhxJ1HVU5KcvrsEoA1ufzi8t6dK70KpnTfB7fdG2r87d
jy2Y/0qnoKAht11dOHSlFNFjDiOe0J+cmuwICxzPk75/+8k/UTAl7ocW6cpWWjz5e4ieQTjft1Wl
fgiWbMNyOtyiUYE/0/1n8buDO4RQDxcLflSmwiF3FsJraHy/NIWWtn31nGZUzO1ve1sIPrmusQAk
CX1H08xqJkZPMyivlvrUn2OrpRfkh/J5G1kqokWHqfyzjTQ44Opxzf+g0HyTIvD34JoHqf3E8cTV
bumR6YtaHEXicCFcYycXOXWOhcPUUGP2ESXRc9sVhLt4+x9BMmBQcV9kiVVYSgaqJmrmIxN6Wlzv
p97LR/JHfuzKMsweUTk7jw5P9X6c2nTVL0G5z6VVMNGwB5Zm7/VLy7d1h1gD6lEg+wS4Hjmh6cX1
wiwN6x4XP7SIfTkhJTIwEyi3Loodrrm7CVH/7QkVToNkmfsO014EkUKrz31pz0c0tc+RwDRiAOMm
+/mkTJ3hdURlvyUWS3RmUpFRXonxC+AjxRJ2EUYOpH8vgFaJMHdyhqyiuOfvxWHs9+hfkClyWkQE
n9MODdL/qYHhGBlcoe/enU4rgrFW3QvzoThTbJtGNZPSZxHZKYiDfFNhuNefwPUY7uNUm9ZeIBug
4dcwUAqfB0FCm3sB51E+YJOBNOq9phNHxBy5YFvLWcEgYBcBz2UGTCaT4imZlad+ZdOv8CRw0k+8
XCtfPsWPR0E7WACbJMqY7cZyZCqmZS2JYvMQXGEG0F4PCABc290PLUIwS06cmAluOr+KrDR7mre5
ULsCZsrex9utscCMr2UuZT8LHhQe5BWr11k0dO5rvoJbegYp1GIBtBuePKtsGKGG/fkm6boAFM62
wWr8CjeGLHY9zdjkr4oT/AzI6bmABk/HwIOACztZT/Lta6OTNP70tcvZgKzO2o8WN44Y3OXjDKlC
lfyb2qC0Umz5pAXlqwvtW0VhF0NaPXb3mGKiaq5ol9/bja4Y7QfpAQml/BUaPilpFxq/Ez6rZw28
U/Tivm+ISdt/BqbUy6RuYtnF6NKG0WM2tmblCffTAabs6M8w9q4aKWLZWwR4Rds1PbSvoxLradVO
DlWsLouMxRFpz47ob0Il9mWBGZ5wCxWU2Q7iZt941R9FDFoZGYd81hPyxXisaGNSwSJrqew0gNII
kkrP4kzbDSirZqQUPPlVn1d7XVg1X/ucOMVC5hYU/tvEy5xXzN+h1mq47iCj6uxaesYStiTniPp7
lMOXjh6+ml6iK9++s9uxxi7PAG/LYeqwM+pEGhjVL0GYi7i5+HUc3xjBY0YrSwa5WN222hy2uWrf
ayixSFYeTfZMvCSk0cRcOMzNB6gmRZgnbAkeKgot3hW49Hq9NwxbsBP0X2PsHc+SOZxgqI6hqWqe
LRouJtDIMLXAiCUvs45HvpJD+/uqswwr6h+s576y4lhULHv9Si5qeorjFTv9IB1KGMZxBQosjYQ8
HNT1SmWWFAzzTy/F5Kc1ZxlljQDCcEpnds4j9uIXLmaUTK7MMQSXZqWbna3uyaHGzQ0/1YSKKJd1
pi7XaOhtVLCLn+S+4Yckqk+aEvX2vO1ZaGi5dnVSLJrGPJ+k/3EhralFpEW3rKzlG8zOi33EKy3m
Nc0FwvyPLYaETDODVOm3rrYnUH63KeMo2puwqD9l0J81Ixma99fAveIXF8M6wnFj+NiXjfx+HBfd
X+CUn0hhdZmridILem+I75X+BJV1wKESDH6X+FE4FC3MWO5hBmQlBLhOZC/bJKP3zMXGgnAsCnCA
7m6ukmmjVL9PnGm97K3Dclmns2ms7tGZqLnWyKzoqkqY9oGpoG5aSggs3VVwZCYmM/5PSBw7wtEb
WnGo5uiuspWEJ+7ZXMIUR1hogtZYx1rkiocpTtU+lUZ3uAgHLd2TLx7vbXPUJzZnYAUz/yHvylhI
MNz4mf9S1i793tmzPG0qrQUE/ime98Sx+l2JNxZkoVBvv9u8zw2YjXyI7cLG1DANkHG/LW0Qhywy
7AuSB6AfDdb4GAWwJsuPP65MFsb1YXIDzOM7nGXL8AseoxWBn+AlT02oGhjgi3dzNKRnho0IVaV9
Tyq6t4/8eH+E1JMq/xt1xBC4xBp5P5UJjuKUqaw73oObsHb6sYbr1p4eFuAd3r8k8J0EvC+D2Ewt
AJS9+dH0X5wtqX0ssKxUB+MWA1qYxrQwyc3K/mkpwFnUL+YUaiUWtzNiTDXjif09I44qcKwPPOvp
CujTgZrifrVVwTOYKEbInP+5TS3bdllX+9R3CdDXqYIJg9WeGvxdeiFAsKpvyOkGP11eerWgggZA
eDT//4Pb+g1euEbMRzIi8v9JfP3gE2VmOCrBoGK4gs7cKnsoeq0PVKMiwaXz4Ew1bFA2/DOLSiXq
sayP+AOn7Cgp6GaVmKmHumuFuxBnwKTHNcDKpmSmLEfTu8mx5yi2i5YyLXA+sNVpi3Z+uL4xOMLB
/NPdrcRaznYCZ7DPrXT43aBJAWnllrcF1b2GhyVc8Mi4u5c95iVXvU7kG2kBAlEWXDLI8r28S933
OjCSf+4Lh88djymWZhMPQJIHP+zExPhPupGdELcrmjmOQH6R6kixpVm/5IKJ5HvwZyrDfuaSUQQs
5lI9On4QqJWT7h3j87N9+7e+a9viaoL1DZWX91lQH3TJMwMW4/ByGFcP55kVK0cML2ZmLpkysDNj
kYav/0wgkmJeB/PXbdBpkT3qSmaL2GunnyW5df7iYdtyVE5SbM1scuRIsLNOPrf8bc4Ufa+drVKd
Wn7i9dOXaJCWSltLlElc0KCMyfPqOFXRmO44PxrBWSya1z+B6sSU15kcRemfFA3LVwasTxEF03zS
6wRW10hVia7nWV4C+9h5yknia+LVmzHpSYgt9UNbew8sangLXu7rWrqzJvF3nsXhDLg3w97QGh35
V6Z1arXnP610k5jwEORVQT1lJUsY/3MC5NlMIP5fWqjFKiwwMpOMGxTYYMmj8IFbZ3BjHv2Jq8S2
fJ0JM8hjSp6RocnmSncuYce18OQf+rsSUFH/v0U6mQs/QIxc7LAKT00iUEsYkcnAck6wI5SdnjUU
qDxClI2OiZ0LW3ZqktKxxmwXCd8cdgKb8lhHCFI+r61PNHvCw19PoecBKtqziZPLMGbQO7ha6na+
6Pz1pNLPMr0gocRWh3qAii6m1Mt9bQbuo3XE4jrjtpBgiTElZgFSmt1fYfekmRXvmsQVeM1++1FQ
grsvy8Z9sujxIrBAqrZtIqetXghIw5MwTxszfZE38CXtYBE+Ay55Sc6QDTyADPS2PYL6UqieiSMO
3Z+CiNocZwTusjrOZOuN/BQyMGMcmkOO0q7G9E/SWHyeKHt6llikrd8Ny8tCShCE1VFFF5Lvhrj5
qtFdOiXnwSWIINgORvxpGwQ1bap8tqLbsuhshvBUQBaItjWLV3YEqn0fy91t9ejCYoG8+LTJ3Cw4
JfFirjBjI4Wgnd+mYQP3cDEHUaRdqvBHkn0QlheX6rPcFI83+JQ3RRxjcrRaBbO8qSK4QjKuMddT
jaN4OGGf6reYbSkvTJkyRpIuYx2Wz6hHKyMqBSVo7BXUiGQZWQ9o0Re+QLFwf1T5tRmjs4gH4G3I
zbiz/jg4QI99JbbFVyQh47eDzf9/aeEp4hf2FxC+5B/qpcJDs3ISHHx2amG3571f32/Q0VO4mMoh
bo8QkxghJizjMMR3UOA/1NLwVuOW4qFnIm8gVwOG6l8oGGZNYFlyjxrA1ZiI1142VtwQXbGiGcEa
9CZjWC1PKjIbrDweutFWXeFBDTyLpfGGfA9IHffTKZ1S9+86s8DVrp+DbLBAvqSgEr7UpUahth/5
uxC/YfdKu3NiWC3YyliVSnKNqVMhGf1Uiu20Z/0GVcRnscAb2+uaQOPbtrMznN64QJeRiy+SirvI
F8Y+gESBKv9eTP/NvsUwPeQoU22Bkx9srXrDIicqpUMErgD2XIXdtLNQ4QOMpdlx6WKziDgFjW4s
8kaCrwkEA1jd802IOtFAJAmlwnRmSFqiybWQWjYTqKPif4rk/SbjAPYbHBTPpkbO5lzecn0lGi6U
06Sjg4+aOAITF8IFNb3pe3eMea1U+WEycwffnUhmpO4Xzcqydc6yTt+OC6geZ7DmBLndG9Fyi4PX
ag4V0AXCulhZiK7flqk4Jjuq76dCwDwd9EM1dMtTluXoeo1Tlwhs0icmXxStasw0OYpN+uRJwpGt
RAgPo1SSieXNtfsOtsFH8OMNgx3au7PgOiFYG4kpcblkXSrjTCac1yMBdMGnaUgZ3aC3rq7MMqZr
rElie6d2Xl6h8YMsiQGQHzW1S1v4mEhlGBQHe4MIcUNflK9oaKmGRmahO0q/kFqSQJDRQcjb2LEz
8VTKSCQxbyvH1/CTXcaEqzbPNILVsf2kVvmDCtxqzSXFCDBdq30AbpHdxX94fGq1m9TPn/jsDhN/
wsF8sxXFX5nw2oDomzXBN3wnmE6/iUo8k2M17X/5roGmQDuuZu1EKRkb+5qaNnkiuUjYUHeBg3gh
Yq9t1GSFvbex8yaI9ILdXSfn26NjvP6NiRv8amvWqtQuKu1kaLWarOMh9nqq8waGvlgCxMiERSjL
xwTVyzaAEpxFwQCcak4kslk2lOyEVoKI5VyU+18tt9bqtbzvDGxGOpci7H+1+i5qqG6TZjyHlfLi
cRndI8yROw4V8Vc9Nh9bXxn+dhHIZN0LN6eWWW0C68AeibfvzbWjnjRK6Z11IDJUfhhpmJ9CwYKR
0ROkuZTIHKS/FDvzMuoGiTZ5SAJd+p8eBc8FlM5Ozbk8uBIph8gXEpBFKdbsXTbJoXOqPYqwbWqc
Dsy15YGEyHz/G9eZpMS8zMW7d0NDmrCc9w+Q0SyOAS9VdAcWc4eRSsPKFTVagF6ZD5JHXQy3aUOt
ukm4ocQsFNF8hk33GwiBl/mevbjJVGauO9CiPiEa4nNN4/tNeQJ1V+mzkEltbnRnJsNZhhph+vP/
YqA4aHjBrPOvdK4n9NPoRvdYThn2Qz3xNtPpuGn4vpXgxM8BWvs6ewU9wMbWklJjY5B6gvWM72hn
qd3woEd2puoT02c2lP3045sov0CyLSTfHc9qRMRVJA7HPV9ehhi7reCArR1XTTgQatCgU56zYfoc
iZ8X3/fJvq0dnSGSYJ42mIVgzrBu7S1IDiTaqSQXeCCqj/FvOC+plL2uXNJZ/RvIBBR4ngZrewiH
AasFIiPcKnf+pWJ1GVToHYnmNgPna981qvO3zdBMlHA0UZuqaJMSXVfqUN4B4dig0PxCseTfdyxa
7SgQp0CTQqoW9/QVqmqq5fNR/8IB+gI68iVGdKATt6wjaVcDm+k2TAtFBQT+0JVkI90jDhC0qVJQ
kYGX2mVOCT3czBRDBe0ojaDv0vNHTil2ThAM9WGn+lm/RW647g0YNhn0p2P0Q11ZraV7hIl2qLJC
GnBzYU87/mNPYwvo4EZur6Q5MthidKQWQjKuk/+08ay+PEFX/Q4P4PYk7gewbOhASZ2DA1iGeIRW
s+b88ubSw1HG9t0VUHL5TVt7a7YNWl4ZYK3/e1dIK2evFHCnWDcHe+Oe77zJPlkpUqSn/MrIG7gD
msOl7dDCyzENs3buEnHYkSghc9O7m96E/ryepiT7gw14zn3fYqq5dUHe1idPuPr2AR9VaqMOIPod
z+2aRV6Ye+YqswNC+cA1Va5ssStiXIjyQerzdK+5WIPcipn5E+np3YUEebLnRRK1mztD+daHuYAv
4DFp7KHAr9AKaN1ZbS6bsNZihc824iXc1fsuwP/t7KNwQkPQOTX/rpQZQTstXogmBjxl7Pzdjo9G
VjywomTzCVzhNufQdTrkSmLTWYGjumE3W7KAO4IG0Fa0iyWpdDRGEeYcBa15P8KfL9DJQI5L1IPu
/XTfkts73uudnQqEL0fb6vqv2njusOs3K06fRCqM9Is8PxHMERasuWWG0CQgRb/U7YwPr9DWC+Dl
geDRYG1z0yskhdQ5Vl3j+GRHizD66liF9MeroqLgspLlaUOlfZnYvjqrwjNBD9zXL4R4eL0YPQjA
zs+GaWkeOMOOBeUdSOub9n7holCPZ/pPpGc54MqVCLZfIMvKyTvPOK0R7C83R7EjbG6/dU/vhQvm
s55P/Rn4SF5zFUsIHO3RTe5sjBLHtlyRM8K+2ZePe2riI0oEnC/bw77E6k5X4zVkpTo09dI3g1om
YfHy1sz92PvfS8PU51iwpEQZ8OqjcKIA7q5FjGh7GTeCTpLFSjzQo1BTvBluUUaz+DdwjiVuP9z7
taC2T/PjbmWhLO/MNQ2XEPbUeeqAZSbdw4cOzLX4RBJfbwoiLB3Qr0Qik31zvmJXd2ZsZj83qPRF
d/FTcL37wXAoVx4O7SBDgy4h1FK151NmV9q9RiwgznY4LKKma142mYyrPzyW9CYRWo9cHM7bIBjH
6l7y6gJE4Gna+3zPTA+tgAl74oUUqMqAhzONkAXQJn6jbtA4YWkSVLhXbrsBPL7DIX33OfqPPtrk
BsU4vCJ6xJ9zrvy07Q7lnDCSYQkMS7lRWj+oOIvPMWi7i3bE5FUz/1tOXLc/itmWPhJG56zWLFhi
di20AYS1BPHSA/+AZqqvFicQpmpyxfR+d6LEUC/b2lycPsCrHc3C3WVZio6qROY5OA4VKgXnvVEG
kKcvoU7pTt+eyFHFKw8vqBawteHvx9DZRTYSQM02f8kU/daKXO9LayydoSRy7PuqqRybcwhcZctC
39VEJ0fypDt5VZJXRU5ZpBDz/GmzAcW164jseKDHeXKaahcYCROFmXwdBNdgLNIj7ANmfa+j/EMv
W9d2uGQy7Gx8301+ENgBWdDtZRnSc6uG/fiHjgLV5cagCgK+cYR8KeQahguREkKdo/KF8dfA9Q8f
b+fE2M+2sX0N4hebgKCn+9Jyy8ajmuikmmiqz61NjwsPl000NYdKd76JxxHB7Eqw50keeao87G6z
tcBz83wmSNo27M59ZiSjwD6Wm0GTxOOZnpeNutQm1DKTyNx3Va4fXTPOENdnJFhkI3vIt50r6w17
z2yIVvr0S8anzcmzuvTxKotFFszVgKTXX8uOJsT0NIRH/NAnveMxl7Vu2je7XRbuESOh/OGkigLl
7bng/mnmnuKyzdWZ2/VpojiS9/S7/6mK+LDrOVbZW3xJejo4uIMwslKP6s8bcJayMTraR730hN8Q
TDKVUrFoAOzaNAli97UUc33kxkgCHGK1i1XfvUFIyX0tMEjoJ2qU1EJCitTUOg1+PheTLLzTPZpR
uJulzB5Z/W85SC6FqrFaJ9KcBMpuIBGo8Xk14VH2ixT7+LpFWpJA/KEtOZM65jCYlriwhNZfc0q3
OyCYjPIRNrzWB/v4NnLz+okeaQdGsBcQOZf4EJd/hfxcTKTpGcaaoVszzg9+N7u7iWBAEMY9RUu5
g5dqKQgFiKT59SfWNXT4b1UqZA19Kik71YDVDD+cJAKQ9IWqmi4FTv5bbE4w7Z7nXLOXzCFq6uts
xRkosigED0uJd/4j8IZwPgET9FjZpq1kWzZ5nwVXigEO7xznWOPcdaQGg4akaS/8ND/vmTLQ04WA
mQiOrMFgIouQJsVzJgvE6w+cFQhgtXTZ1HJJqvvEh9tkpU8s6C967fy3esKHWOI7n/j93e7ypePx
3s/9woL38GlZ0vRU/hucgVH+VXLwN6CW4Lu9Q+RJib0o1G4cD/Eoi+tjSc+oJ42JgDFTsIPyAVBt
M5J9K4hLoTsawDVZTfCpPqq5JrooEyicKJI02m3xsN5kbDv/SwohnIiGNgOBD5BTQi6VMGwnK3WZ
aO924A1fGlmRrNQa+HU8nB3XrqvFW3SbXlXofvV19Dvbozw46Yd0aI3gDX/vrlz/RPzJnrqrCGVI
P+gcVmzckfv7GKE5RwWyZ1Sngk3wKaS9+muYvXs8/nQwtNoCELWFC5UKyUYOFti6UnQAwhQy8MAX
Zppkj72hDV7k3z1zIKyjxhzjApkZEnG05yVHIRa3q4Pe4IpX5bHJ6blTt3jvTejcot0nFILFd98R
RFi/g4OLnHLAws7juWi/FUo9yCQsxC30TqigH0gugrzQEhARA5kMO8xbQCMqctQbUFcCIAmPjc0M
Rq2/rLmADfcIMjYZP7va95nk7jezu4H/rHf/8axmEL1VuU6xFjCJb07iaAIs5Rli+JmBSN9tZKQL
sspmKejKEliNc8sobbOHAN1LV8OADoH+5Ermotbvd86tOKrIgZmdJzqF5AS2wCMyfLn6b2qSS0UK
yI2VNOT//hH1ArnlJ/fOEgN27GKE173iXzmOYzh9fDcQgPohvwly6FuMGgL4Pbwdq8WvmFfbOXIG
CRaqYQp0Ex3qUrYNEPQBOigaobmsukQwFFs8dkUtosM/fLfx9eVWckgzT6T2snU1mYb/4MqHgh3S
EF7QIFmljsynmRSvQ+cLa0gL49blM5JZmgBZhHyXTq8QrzOQmEBTZO0M8q8GzwOM3PX44pGHTX/n
i25YjMnLoWd5u6RGYWgpAaYn3nl7OXK/m8jAeHw7Ec8/8Utq3pdtcVMJRRdXigrzfjzgSWiqaFng
h1zECM/Mf50ZTuEhxiz6bHk7TjmIc1Rdc0iEgW/au+d8d+EwCq/rdM75pYK35/FKM4Y1gIoP42X3
P5tsSr5oI9oIOIOcTKgVoDpxhc+LwIdbLiwDCodwhYFageJuyrzhTrd9dqKKYLhGhuDQ15+GdC5X
JyDP6Ec2RIJzpIrG1A6RY3EVTAJoaiscZb/vKhKiX0bApH0Npg9Lo1ulBMI/BQQj/nDqeqig2f6b
WJ5f7dvUO2FSDlI6a+PpGXItNQlr9yLOdqZrQryA08yVFWjCPcbsDaZ/7VSihJuCPzgZ8+y39nvw
CdrKpBPWIuQ4XlnmmIuTu1nXhFrARgyGTpckqrZGE4qrCaHySweF3gZ/YPgrLlgEbAq4qEctI2VT
46Kygm5+vVJA5bX4DJVnir2zuEUnafMBgJ59Ku3eyesgzW9cTJEaE09BsXW8MVdS2WSiHnZnLatv
HHPhhwreYw9uM+smJUf8NsCp4DVJpw/QsB2kqXOScrUJu/MgX+oUVwLoRzB7X5fw2HSNSsFP2igR
g6IvPm9DKV9dhnMclOjj3jH+4j7Sx5m3xlhe9VYmppTCK4wB3d/gCCArioTSsET2Hqiz+mlWxAS8
FY58tnzDmkqcjLAruToOxQcr7ScTp6AWHKVpR/pGXvc2WyxKDdyqfBqwd3UEGxNBmVE+oVNzSDIV
DwtrA3kuJ2l2UYnB0aDjpMMiqjxOXNKjJvZvKFZz5j6xEoD+KLPiosYFudrQUfQ1ezTKUyVlbTsC
h36/FwCWgw+D5X8M0brlnEddymv06DlE7s40fKZ8OTDKPc7e7I/KDT7MVlURM5Gw5+Bxkg4NjBUB
4u+GbusJVp77vChdXs5WZFavp2kqm/AKWnEXMYfOksp9mIAj9r/FZo8ZJaaCDiKIf/7UDz2KN50J
7WOnV6UhW2kHmZ8PL8NufUIaHE87KbqB7qYqWh/YVNzXGSsmCrnghbbEf2XUffSASJBImxXfcMh0
6JR1GxtWyC5IYZ+oQSUn4mzItpUD9J/kJzwcKtTbNgSInButcT6/7xCFWpHxcP3ygNH8ZUNx27Yo
i+3/Dvg8OXX6PN2mcwnWyhdde4VazZVPd5qw7EhtQmbkUGRriVvvhUeDnaoEdZIHU+1GEzJgzpEW
BRGZfIGAW3imPug0LOgrc4rk6U0NzGohdkb43wkqGH1JD4N5QgZ2+zyX1ybHOxiFu4g24R7hoPFv
hEg8IbOJtLm7wPWO1+3pup2lDgKnDo7KnNuKA+C5SEN0do3M5n+p9YI67fIkDX8t4TRGK06eV/BW
I8GRgZdQZ2FPrPJI57DuqsIoGP1cuMo26kcZ+06EnJBWK79/qPme9j/EEI+aQj8W7+JeWcSlUkp+
VqFcvfhUTCdJ4Usi4nkQLELJpA+HOocfMuktSFG2a9zcAseQUhBs0L9HXBdNMdh6qmAz2BEVWbop
x5XQvHj6EHf+Oe774D4xQP1Ezb/hkFt4rgrXQ0oNNKtWOsW2zBO9IofUksLWgpsN8DaNNrbJKWQS
hfm9P2PpKmq0DdTVjRi74ko8+xrFqP5+kqlDWlRmTb+CTFD7tOVFDGjYijv6nhTnktCsUHhWHFcY
9REeHcEa82XMaHWBUUKeNJEmg+Zse/LYitk4GswtRyl0mEO+oU2ZMFslfS1FANp3aBa8G5EDwx4C
RXwP3EVkLyZDz3niEruegVo9sLpFWZ/rHP4g7+oaa9L6NY6THgionX5QuC2zCJhh49XXNzUawbVL
VJyGoN+KypWuGl/lFk+iXg3YYj9B2DAjL97jA4e4Gxm7UMhwm08w7Cwm4JWTbT57ev6BqIaR90dT
y9EDpmbqFVZksgHmVvhMa5+ofkkSaCcbgoyI20X1gVMQ25PPjUZNG4RvKptdcYIsQSZiWTjwlHF/
T6yZq1komL6rOD2sNXNcqj/j0gGMNT1btrhxQI2ejmQIDjBoX/FrQoWYuyg6hhSTLt8WzEmVQO0c
L/trRluc8px4ucEuVMQMiQSXYQOOO988Vcu9f9hfRwUDpTTH2/bck4rRHHnlFRPCR//Fwdh2Hd5J
bzo023v22ft8J1BD6og+ztB/kNlT4d8+84JxnTfr/cNM1D1qax9/Zmcs1lHjZxCnaApYknIG5YlD
eKgGKMaRpx7WTQwxWFaB7gnpb14xVZMhalnQbkmRGUPmjYuaeK4YXDUaoUuEEirmIxKxP5zIr3op
cUSkk+O7YJbnafiuMq17LyC7YtG7Pz30Wr/Ib5jkD7P0v/TbJLhg4I4gCUuPa/aCeWc/9od0AB6u
kmBOgKT8hfLyeGie4/3+O94ZZUToCwrTLGKRJPjleZPaEQJoQcfIPgzsQzmG6Z4mSfvPRozlFt/t
zJjr6D8kHvBM3SwTLyI1Wd29//zMV9+LsmXE0u1efPDzHwk2ZwV/o11WYp7j9gY5WmOIceklNqAb
4R5QxjD8PSdkoCRTLeAYebhB/OT8H0PpNSFvxi150d+oulTyUHcDOEO2A7m7VHbiV+pGiaBajgLX
tKTCecZ5eQCZdspw3Ht7sXK58nQsyjvDP0aIBONLA8RWcItcO5yrOneR3vi60GK/Cgea/cS80Mnj
Ww1KtqlXTNg4wvPgpWMPO0Wo2Q3kK8uQhC75Vo2QO7NFzak2QOsI9tBSeg26KVi6AYHASAAe0nWn
irkJLQxQXpxP/k1w2S+v9kAkxKRFXpVXH9oHm8JQpCPO70ML4O5EFF5vL0qGTIz2+w5FEGdiOhbM
KdRyQhU8N4q+O8PyGB+E2SrebOEVhL9VIqWV+ARUcSoitDBEGLP4nWSLSS1bRurJH07fqe/VSTKb
vOJvkhxkRz5j6aZv9/CqooiqPuY2ruMK6bQ5zdFWxNZYljsfQtE3vJSqtFPCexYE3LufydlBg2li
vGaorUcUlr3bwao2ILvFeuP3phTt3m/dTby/Fu/p3Cnqh54bz7XKKF5mJN2o0aogD1eI0x6MNRXK
dBIIilwNC5G1+GDnooFRGYhTDZ+td9qZXh0vwYgkLx1CPZXH173KBsBUCf8bYzYpxwG5OC3JvBWd
eLV4vfi5yqNvGX3Rzp/Quf555jVe/eGp5Dukdx14FP8e4oYERCMfIUdOFarPTCOSW42lKlLV0HGA
tPFv4HHe/HIlY+ZfeHvyi8ihB0x/yYuWnX3W7r9Vu0hSCdKZai6RfQ93m3td7FhMuW8XAgn/9aeP
068jMwkIXGcXRmuKOqdiEJ4w9ikXodUHn7weJsR48CxwRY4lZJMfBDEjEQ3L74U0C3m3a+YlkuES
p0An0/nUKZX4Bs/5hKWB6yXEXvK0YGTbpRQQL9lwoPNV5CUncrUSr6DxR9D42IoneEPOVV73YWd/
nvxpMuu7L+NSStXyjozZDU2q4LWcfWikEcb8OM+lrqATKCzeUAwOD/IYBASnh0WACDrPsZZ2AV9A
vi+a93jlGpbjX0If9jBxZlQB1syvnUmoqs4PBHxJ1CYauboYx3azmXjuIK8EzoMOOlI2gO94c8u1
Bkcf47I5DLubEQB+fLFtt59BWWYVkTaqUd/+E6OXAGAfmriu4eireqNN0Z4sd3Z9Ft9U2vs/2t9w
70FHxgLcwG3smr+syELU/mEoEzZybMyTjxKc1h8ZiYyXuxkaZV4H6erSWctIU3R4YnEYaJTrPVQx
lPAjYabmR9Mu3tLC4acXDl8X0rnU2B++FPnVSMHheL1qYLIaBVrvuP/1hT2yinGBvvtDb6g2ErgR
oXCy6iM76LITjZq0zYn+mylVRGDdDxdrEFXzv37XdVNLf15jtSmWnNZeAeCdtMgcqxStCzbCJ6dS
m29vZ5DzucrlnxyUTfgqUJCHV5kalf/CQla3cmcN19NhIbdUvZvtM1fQBCnbdOB47QlePp6Hfd/b
ChsCs1sG3mEQ3TykPe0UWIcqbJd9//Xt63NjvdeXx4t4IPXLT6qOOSigz/X2EkTcVsoSw8msQVcv
i5Dvmbdy3lSTqYALJz7oCH+Qly52OFRgMe6yRpB/chfiUkrI7CAUL+vnca/OPLGRiWeDCAycfnNh
dXzLLq02RCgrC54/UQteweZFVPstoa82Uaf0fbyLCiy3IshAkJWguiSQXB5wgHwOVwXod/20UHqg
LQxWpT0r3KKb7gifkWtWkhrwUckffk0Tu90DjaX4tx1A2NZ+kGQsJpUbK+xsQdh+E6warydokSqO
VreW7ULx/EUqx7ENtElywfCC8xPSFIcSJyRR2upfHktpM8G4Ct9eaG51QFuA+Mds2JE1+kjaQxzU
coDVSXTva5Zh9gdvqEB26AaYmPOkHQ3iiQC39nSZh2shB8vKdb3coUmkxn642x0Dxw+/yGVbtXhW
1mWC3gaGQXX89kp8aMtKT0LoxFLVawjlhUYiBBzWXPi6cVywO0gV8LJa6m6gPgoO2X/mHutRggZs
fj/ayOP1Z21HjhSSnWciz9rZmF+iplijHvjXiiiGSoU0R0zSmBJJEbxs9rpZxEAfSb0goVJFOxlj
+gP35c/Qi/RakvtHgb9Giy4hFelAEr8JS9MC6Y6capyaNvxh9QUBLRF1GHUj4AJ2fHJIhnB3UDDZ
9PodyY5hOyvnAllf6Rl/EnHim6ewwCm+NxL55WjU4kdhGY9Es1n8M93Zge+NgBVbbNYTx3EVjaK8
GHzsLKQM7LmGekgcO8BBzo4af6jHueWgBYdfRsFugrdfONmCeuwL0ULOWzZSHZXo/SwGjf73LqlX
as6nRqmvJsyLG7vsrF/l46gCA/lDS7VdODaApJUiGkv7eWd09dHwsKVEob8rp1Ra4XzbYTjFt3Og
o6LQQDYh8CSNLOb8B47tZPd24FabQm6ifV46j/DIA+C7wPsxiVUpoUx8t+8/F218snlQp6Ap4dkC
eJpdXq8SYSniFMvMdcyi1VF9GQ3XwouvWm/1KC3O8kv3IT6MtR1MH2Nn7o+rkzEh68z3da7bsAzU
YTIsxWTUv0dafAbIU0WOKLOUoJFg1+FKu8pjDXkk0yYAue4f0ALbMz/gxW73Bu/8zA6h4oHJ1xDp
0ZszhiXuUNbT0pHfFTrv7syIiCEwQKYlTkGd8y44WwKrUZeIlj6zNT7SLKtUlstLBx5BfquRR24v
L/BK0ug7xGKu/TjcDly3NccPTueuWIZqKDF2PFm1zB6QOg4d3lcveSZehmiaapLn9+dmHDx3zSJF
o603uQK1kL/0ra6/eQCYhu8xnKubdmYL44BWXXlRGEVYtikgb/uLWPDEoYZeSgsZr3huOfgL8OnI
dhSjdrch4XPMbpcQryARfC3fn65UdFmWEnz2Ig4ixceHwQJYtlPImgXbXdJFLpsMhrDnKQ/vVhxZ
ZVEdnCogUrq5eAK64dcmS6FNI+qZPqZrAArPTi1HGzo1xceTqiY7wYvd/VCNw0+crn6IhTKgff/I
o4K4OtZ+5uMEd18VMhvEFGn4DgUX0pmTH9mf+DOZ/LSCfPjoea1M29PBdqtZ2B8oc6ZxCJOsfZCk
U4GR7oZrdXeKIGTXR1I2tV73asVLtqhvcMJ/T4KQ713hoFLaIsA+lztWE6wMixeEyZbEFy1mU4ME
mqinITQSlyGHkG8q9MyHKIhqjQcojxsz9m1oWTYr+0Kzajodmcjnuc6k9U05qU2AD7NKbs4ZJM0q
LDfghblu03e851JrFmS849uexNjZfryHtwCChYfNbudCyMEARFEb6x74lBa0V50d9RbJqulGVk2G
rY2atl30nTHQvFRfsgwNh+vciZsVXSBIzctzJJaLsGM8xLnrgPOqw0578bXKoi3LToE5AQaPxC1q
lbd/huc0yAVPw1HpCFMDGotpKIIv7lwJnBN2wuIbfIl3TpMQqofmChfCm9ig8SKJo5/OFSOzsB+r
u+fQ1cp8qSA/RSfnPFKV28dDePRvJBluz5WswxJsE0TCuqvbNJpCfT0XTVfvKbbOUw5LRzwlqRiG
el3pnWCcN5ludPPN/HBVA02rUDTSglVthem50wKwHPmERRiCZb+GPPvrx7dKPPEYARu0yL1FCYqs
Qgm6lyk+S26XXi84Jp8V9Gb+7MQdpLylBykOHSXGX1z74i1Iz2VGh07ryzEzJCPzrulY2cSya3/5
XIuAyejW6ktThnDZAXmm3LrfGBfadyl+vpb4GbYO53jGNKtJ9M6U7LLRabYk5aaCacOjav9hu86t
aw8OQBsSlbeyDLOa5Z2ULphgZ0pXwmtqcpEd3yld/yPoXQMLOGou6aQNwjATRLXxxJrDYzTPT2WQ
YMiLNbQvN78t/kEH3aTzHkE5vtPeIZjhJBOgXybXys5poFbZyQ06Y64QmpuY86gVdp//orCbRHSF
guvG+afaWCCgrZoQ4AJnFG0FyMPXJmfgnFYV6NzxOgTWJ2fON6Q76MLlIb28oVoKCNyOk25thMl+
UwVp3dA8xDCkUZXaIvgCoccE6bBur3AGxT/HRXBr7naSxEY+BcdKxuQr0WSk7/W/7AHEzdBuhZxQ
TAeYJFtmsISbhaYcRgTRJ+uG9x57QI67mj0ydPpHBY5W+hiwj6qqIG9SpwHal82+esl7QLbh1vmi
kDtAIjhmE4MhhMT56N8hj+OTUtkjxG546CVWUPNVBTaohyWXuKK/jgehG+KjAX5ddX09j3G1w9V4
LElwKi8nyoUsm56kP/+8QFdNiBe6Jcu/vFOIY7wnTzCqTgqnsyqo4bPbpKcdpyx9jis3YJFhy2Bo
q9fA4JR16lQFiULwyXmVfVDo9osUFoZp0QGMWi4muFGTgrExdR9uvZj3x33FIkApjC5FVIdnq5ks
yaPXTjYe9ugxCAireMi6CLowjofJwsaD+qmSzhmRfbVE5w9OcHFGMN+C8vMzOjtTi83ACdfTNu02
fOHBmzvwSpTQHIzc1FkWHZP7ERDVycTo7GBmlATO/MSqcanpM2oRoMfCP1NVdyZnzuAeE7XBwUXO
6Is3KKmDwZ5t48GBGjZcQWvDE0wpPf6/5M5OH76Xbxo8U8e31gizqzZx01yKO1ARWHxMeoWX0kFK
KZQ4jaELvJU296o0BGtYBFQwsVaOPqeUfbjostv8Qqff+RNiWZQDKLlvx6Th04HmuqYlttif5GrW
MqQxERCARCbE9p+3XKgW+05OGiTjrF5sr3xUo5uAPKNmlsqcE6t0ikpfcHfOS9irEaizZ4Ak3X2c
ew1ZAaWa8S1NycU5RJx6+XDp4nm3HBVTFgf0z0obLp2oMl9uYivOaS6/CrX8XSAWDx9PdZdKTLYC
yVdTeiuBiuV47l+JRI7UJdT7CYPplFBVS4ZHLbiAjUZRVBJWGqCzu3LrqY/PLhswHY34VupYjrbP
Tahs3o+F8WBEcitNS0KhaodIdA90JmTTtiEYfElQ6BPXXWDJ+8pZh9k8rA8iGBbXFO833Ws5snZi
mH817zNzOjVedSLtyKao6viQgjh8MXFU3vvPo7lUVBlVJAP/WAGQRakQTwubnQ+dCsZ6+reMhIey
doeceG9R0RUgxsHVN1vXQDla5V8zlkBA2GalDtDfOV6N+7UXX7uZPGggNkBgE3zpcy6SsRzMNWk9
ohcPx8F9Fj+OGQyk2KkAQkRbpWlpQCv+9kxKBQkJo4ebbkVlVZVWfzlbsy+8VTyQquZnZs75RZw0
0S04QCIvI19m5AIv9DHQsjELPvBFRh//JcW2NL88201S9o7GZ8bi0D984ADNnoRRcb2HO5uFX+7F
MKlQOS15gWD1rLxnrbKKFSPf7Ldri5tYPSy0n3nizAklo5IxOH6kCO4ACQDiDd+GjFlyzuJhqiW0
66H2YnTzXSxZ1xm0QpmDimlyU0ybyWPBsTtwRp15H7MqsH/Dpv/H0ZlguKyot1HHBQNKv8+pHIc0
Z83S/Bs6DfY+ysoql85bU/p2JqYQaWGlrm4Ux/KCU6cxV7ePuISY+b8kUtX4wgi2DXUl2c88sANV
Lxx2iNYYmFfTakhOYocPJ+FSXoW5P6mAKFhSOp1V59X8hgW6kztXPywXYT3d8gyqOwFjLRwRG1EL
cuiSWAekUWAR+zLQ+pG8EJg3Jut7X7Rjlb4tnqMupmy2279HWteGO65ajcd/neo78KCy0Uwp3XDQ
TTuy2wl0dpa3S1lMHjwdqzBQR2tWzYRh/wYeHyuM4YBRvfBSn1YX6sPAAogNNj+LPB2V/8xse9fz
KuAAfCOxADbtM12AlGWXUvEk16duKHAcXFYC6A8jbSBeRRdbG88uuV2zE9CLxeru6s0SGW7G0gIQ
9jHpQkUTbt37qe3WXQ+YnzoF6YR3k/gb6o8VINTxGRJIT/4xBmtM2WXKVam+Pm8NZSHmYHu1L+6Z
csm+oQiU059v/2KiWwHCqsEK2YPHhOPEUea6L1SeW40+MHUdX7tF4ClogQ/xznCKf5BGXuTrGf1r
U/6E/7DB+cAl5vyKayEhjuSHgdj9ObWI8ETqGmdmveTOvvuXc8MHaBAfu1baiyObhXXKNMvZ1H/L
gHAIHlzdcImsHbdhLGdYCTZEgqzfrh9aKH+LA2Dv5DXUlunOPEERIG2YCo/oBNfcQ+oxNu1x+hC+
mDmZkdWZpPGio40eYatMfIxklPhqXxGrkUfcpHA8Fu/2X2lql/QE4dDxWYu5xwVUE+kgcA59udYQ
cPlKO+MUW3h4KPIoIZQ4y+l6z0XRJlL1WQ+gFt8DmF4V17sIg6lHjglt/sd1nAhA/mTQ/zhP9eC+
8KNiJ0D8JVzD6Tdw7f6lQTUa7X3Vei6pX+QtR3Kj8lOL5eMgu62G0CuM1+1qFd4YJ/WfBGKJjRo9
cifpfGt4xckVA29kTDGh3uNPtg1Yp5grOGRI2JvjXrQnK9ip+y++9p+uUa8SzhWftTQ2245rYlwj
7GQ52Y5hMDDdg4uciDaEniI6RlIl/aDbe1OhpNS02gmH4hlixlqmuJgN4lSEcPU4SZReLPFTKMOk
VJ/hxT/FO7z7jLHiC8vKdast3v4hTk3t2pXYXttaQ3B3QLY6UBmTUqOTCMpcsaWhlLJBFZP8a2TC
AXmm2K041x5k++itMAV75JG0RKxV/dLhC/vTvHi7hMAHRPDctugqJyVBr90QXi96lnk6bClbxJuD
ykjv7bMV/uTt52e9CzN/GJwL0g+rxiDB3sXnF0B1cP3XnrFis773PlzWfNkr+DRFs1eCHisxAC3C
3i5nkC6cK7AluW/mYoprey2C7zA76DVrFots7LC9cz8YOKAKnpXwGtPsES39Y+eZpieKkfV/f3RY
MW/vU4FydsXCYAwMq2OIvsqWuVA5kojOnN6UJsp1pPe4oB9ZZyLCYRQOPEcsCrR+dFf6SeWIDT7n
Wj4UQTTgx8fdOz4ZggCiQVXaOnGkUhwhKUIb4CTb5JEbct/+PsYF6d9k7SwA8D5baGRCuHMEfzys
qtN/aN2v+p/bhyLd+SiujPKjMe4K+etn2+FV6M3KDB6hxqVZUJrFfK7McJrlIp2tghyexkOCOREg
1K7ltMvnuEHP6M5TeWvypLsUzDhoCemhKAzUgbs9QxQvzJb6/QwwzgUhipONj8Llj/v1H7PxJ7Ns
fF2M/CWu1eIbwa/WSAhFAbovaUEdosl3VSKZnDCtCUnHCMhFuhioArs/uJwmvbTI+ygKR3xrSZEE
+xZ+Jbprft1DFrK0A7IGjfKswY9kxTqatIwnW2/FJpBGd9xLukFyB94OcP3XWlyHRG4j8JsVLAVC
ROb8T8B9EGccgQy1xEBSnEoWqHETjrFVQBltX7QMTJWtkCmqNlgr6H9DeNaTh8VlEx7cUGDhvh8Y
OBR82J9T6ApqXiwFi/OW57qc+xIVRJuq5by2JD6AlptEV+fMnIFpbGYyFkILU/tAFqgfEcri3vbh
D1XxgHuT/Sus0OF9vjjhtaqgBtvQPwa+2LjSbEn24P9p9Xk7vU5xEfpxANxGP8donwQtXlpeCJ2p
cJAQ2IneieHM8qAHdUk9KlC/SXbp0yAYYn+L7qQD2jNLTer3otdUB/hZzN61h83oFuKjkBhiehkM
6Ul1B/27HW/YzaCxm7zcl2jkN0z28wWV35ZujPhIvWcXYQreV1wEMMrJxfUmpNFNsCWVsHqQSOaP
cFnLAZy5hxPWfJAoZ/ReE41XHHrEDUr7uZvF4P9t/ye4Zm+auO7hvPbgGSfgpThgcZiCSCuRnpIY
Spvf7c3UlZJGV84lUQBCbvkRbddXHHuWWFns2xHEAF8WdWFQ2tBVBfQGFTq5/he9hbnPeQ3H0pxT
7oAP/OUHvjbZv7EPyctc0wBLVSn9jP1VX6gALFhE+s8fIpvzA1qNG1qkoxyk0Uk3Y2nwq+inYYT5
EPryOQn+GupraezXX4WdDO8v37FqhrmSNM6pgFYSsp4Zi6YlE/9ZAYs2lhml0qQRyDQmfZJyfJqT
0wG+jonpRlyqh6qDU6HvpWD1HQaEBb5wf0GmQC1rHlbrKYAy4KPJmc5wx5/W4cVtsTxxET9gVnfy
fO8eK0nqXaiI3fF19fXgE4q5c/7KrgjQojbDQcCsCF4FDSXj6qT8g+FP5r2TlAuDoyjMgNS2k8Ik
JUlPxFopH1lnmzhs1ZpTqx86w9luTwVrr9/lh7gAog6UUVOFCdRD+br9c5/E0gGTejrG17x2QYwq
B9yBk2j5IHPLRJYJdmIkVooW2sKEn9dQYGS+8R2ODxSw277eUSzsrPnZtFj+hTgolWxJ56hdte0s
DBzNM9N3t1EvYDpGKOmqj8r0oek/hr+gtxbPinaYZJiuMpv4SxXrFJ/yN7MB4T91pjb0tQM9Kx1K
QFu9yxxVAMrgjys0Xt0581/CItFro+/x6x1IiMBEffKIoTzQIhsgBf2Ipf3it0GAkDSCaYeiqCYc
VadW6Ff1rk/yOUlZ50AwEUKQ+iniaPNrhlfQVI0Xx20/s73o3zjW71I0omRgxaQEyBETq+bSwGji
t39koSt4sGyBisEK48ZpMzZi3buWbDBoFmG5M50E8oaYZANGDEHhfNQtGzkj+mH/Wd6lPs1N51M1
BnMlicdlkUKx2hY5EyFGKzcDMzWHxn3BAhLHIGURjPPSaljNggvghEodO7G4rqM0aO0Op+aEuZQ7
8W6DDb6lbv3WEC4vIPKEK3GmETEySptxFJw7Y9N3sIYnDMOOIu8yKNK4eOt56GiVn0lUvEUIfClP
442vmzR8sYxb5c6qQfpovmFkt8JC1MIF4H7YpJWM2ne1HEg98yYhL4PE/OTTQ6jOOnCRIOXC9/Do
gVzZEu4Dkoe2G1hx5ki/8YMQ38B//U9sbjYyb0VDE7laN9LEd0PgGbT6s9wJURV4F2Mj8mUYLtko
3zcm5XXNTelBegqYn7N7qPK/tOhZMFK538yKgwcPQVJqjctdTyrGAtqbcmwbuNLLMeMfR8RVeuxZ
alGl+i1LzelUkytrRzle29emJKtTETz70RVz0tygmsfSyQnptdfo0D0SRvNX6k44c4o3/kjSzdz4
+Exfqq4tv45sIpWBFpqofN2KyXIJxUVe9znuUhdPGo8XEHgIYR2v2FNw5h8nfZrJIWvUa8kyuxcE
GFBBFwrwzQBiT/9KEPkC/sPtWG6/iew4p3ZMIpRw/BodmLReTbhthg2tUGwdinz7tvqf2dgyKl1L
eCZZrxrrhpOw+M02L9VS7aUnI33u3BgY2d9oPnYN9NjLHs5cx3ZiWxnPBFVItful3HTTOVXUo02i
yq1FSlJhuzadmqgLRl+5Cg+yoDWRKws+IK6gycsSj8k7PIoEcxyHXMRvl8gefsNpykiVQnGIviZ9
ZnhXE7KfJlYzxDh7vqKdePoKY9xZuZwMPQjfHuoyQMgyPs7h7s3kUvF2kfMoyt+QH8IjUYzN1CyC
hySmgi7iFXdaXFQEJU1o3AfkZ2Ie0bCC69wF1b31DpFhLGMqpSnbKdsKUgjC01G3Zw7XusyxeSG9
v1o6gtKSh1F+p5iTY0UlCM2VC0VB2fj7ZDqTxdpMYa52N6UNx3AZqnddKu9Bxwe2uF/IN34p+ef5
pXahqW+nWtaKj6ylIrql3Bq9qbQZLm5xtrJmcTbHg8yRdcufEShZeBoH4omaFu9P02lUiRTrB+O9
4XI+GbHrbxrQDj508S6srqjKSbzLCSBLw1y8RE9F/f8spdtjfdPnm5qwhfYbtsBgsuH4tNDbotTQ
iv+2tC6P5U/Ss2O+td3UCJWuqcuDlatlCjO5/oMxLFW9gVPI9+Tgy8Z+AuEzb89Mv6xwo9r1WR01
j7IIX0XCpuCXZPbw3FsZ+0vsQYPYw/CYch0LKBhBy3/ZmwGK03kiRImIfE+EsyuS1qznH5cjckyq
dLk8vHDWSKnsMQj7MIvKmKfuQg/ugJuSc/3jkndX02Dp+aXzbcGm8Nkv988fIMxCcmy/Yf95Q+D8
R2bmhO8oPRCIt0XrOZK2Wl4WWwP7tTD9gDzuEc/rbUJFea1ojccHB9YZYSRemRam2OCReKgvoaab
Eqwtk3kZv8L4Be5qBWh2Z62juFAfhTjiDzMttQKZq4mU9G+l+RKpO83qXztL3lekcv/MnsZv3NHn
RBWCM6lehECkKtikyLGF9ikjZdv8rPUgZpa4tb+/AQcv7L4DLqDOeIuQmKkG30DzYjaW0jC9+p7b
E1IfjUKPrBrBO45VXHyH3TsGPEtULMKU/8el+mgP7JyOMr+RDz/ceELzu6qyc9xND/5opItcDaW9
ELq37JdqbTNKC0hQxtL7vEdRNt0OjGXRQghvcpqevDs7WzPjh0hEvxFNmviScuAb9dznSxOMUTHX
LW8oNN+oZrwq62csY95ZCze2rBy1VWuViYXEkWd3KTTniUc3MIVBncax5lwqKTWEhMluLaSDTvCi
UNNEb+AWvK+Y7hEDqNJR4H5hLZWhlZ8qhQMVK4Hee+T1DCWgVcBXp/DYmOh7pfLFL5iwyg9erBIo
fdN5HSulaObKLSyqqyjYuUwW+fOICcZ9bg/29owtsDfvMAFZ75DT9On0K/8ut5riU9441EhhaVTA
lInPyqcf2P63i+Gzd0TDEn+4AKrmVURfV8X2aZtkg4BDKYKQwDI6uErHAUlVeB34Ny3rYtOhzDhi
LIwD8TDU8tPFa4wHFiySvgAllCcjOAnatGbdSFuxhPNCsh6hZ5Zjv5odMpkHaKNW6evese+dgJSX
mjnM0XnIIMDSxMKIlnlno7dXvxSl3m/KD4TVhS9tmWK7bBSPoukjM4hmPSWLYMY2QMWNb61ACWdw
khBZ3EvKmEKSqRMMDP2005d+IeCqiupozQsZ0ucCAFZXIZhOrT3/jmsZDbERMoXLnU9/3G18LZoE
OJ2oz3eRinqdwL1LdeEfZu+nELpDvR5PKGnORVCIh7gYKzEH7t+o1WtcOd1jIlkGgVZfe5IFbIdJ
NDyZB9TUHBQR9p/iZAD1P6EM9FI4ZzIS8Smi8W1kxBM6/+mGI3O0U7UTdrfGkFlvAwaD2ZWdgVc7
6eiyZsvAAfyN3tvRexhAkd5PsGzbZGyBvIz+6qdr4XtvAPsou3r5EpUfAeygLIosGqT0LF7jlFiY
jKHkdd5x/MqtZIIvMm3QJtzv/x4sR/6EyP+sJW7LbN0DJ1QX3H/Yv6Jy71Z7IyzpTdxyIaW6WDaj
YZfAfJ6xjMQa2aMqyPGUbDJI87IioOKeVpY946bCwOIozF9nYNSX1AN90Y/8Ou+EJc8ke77Iukq7
tAB4y9ke1J7cDxl0pEws0qT4xyrPP8OtiLKU1ONOl6IGru/AGgzp/uMQxIeWJ0AC1Q4bEQsMKC8B
J4azJb50RLayobcTACKQdk28MDXs2x4Ux00wqQvm6yiXCrdg6n0otsDdcknm1oDFIAMc7N2k8k7S
6AX28gahBI/f4r89grM/VDuQYdODZ4Z0yywROnlOim15z9gs1mRQlffIQFSzlrMGkmiaSp5qNp4N
V1WsrqG85Xj8DQDKBjE3otoFw/irxUtHfzGR/kbjbPKqgPa7X87QEKoMWJ7JdJztsRu/S6UHdAJy
ilDuKjbsycuyUZgPg+XYADA1PIU4GXjNFJ/P2tPgmRcT1FAJbKSitnWVMfhar0yUMiJiQiPi2o8W
rQiQwwK9mXC7Gi74bSVJ5uhntrFhAAsP9ufqqey74mR3bOsu+80SK0X5dNLbch9Q6AG3uOtH6np1
MEK4+Rs3Sbj7nw/J4W8wZGDYzyy+DFGZM/pFscXROsRpDOXGo2E2kI9Ntcv5GtcrZlLleZ9R3ip1
UtBi6nrVDhReXtSiQO7EzfvSXiu6B+ZcFM8zO4hTzxS6wrIqMCU1KToHH3BAwyBlB3+Tds7Sxhki
+2aCY+2iNmueuzLDlmRwFfCEK2KWJodxsdbyKiRFFhIuPZdPjCUuc0LkQKx8xSlWA5JMoN32uS0H
NsW/f7IUrMmFzYK+KCa6gnr9GTnqWpoLsonrvMyt49qNQd3MLoycC9HZIXkHLoh9CLkmt9umUmdg
cXMy4FG4vNk5iaFX1HR7mfQLdijXPIa1EFFocgsPYM4OzB8q4ounME0dcbATYMZ1I72ZVWsf6mWe
wC36J1pRbhl3nDNYjUe7XbRSCDIvwrWMpJVzBZQbYRTKHCjhgAjQ+rxhDEaiyGas4tYeDTZwovh6
EOy+AXYRvr8ribkfIJ0RrBq/4obPc4In3F5IwMcV1+ax0IBQfb+2PgLeQf/R+YrRf2IoQ0xTelWX
CfaE5TwgW8KMLr4UYXJ9e/akDDdYotqq4tFTWJ8qeeRvp/MA+6jrw2eyCCCfpWOUd+7/qMnMY0Bv
r3BkK49jJ6o81M+H2MWVRJ/KB5IYNHcXAm+YuGoC7HNxzc+KOooFa6q0wm213fSYl0BBYcy3BkHx
vDOrgZpzkY1GJQ5bmkzfgr869LoioxCzUxFCY+F9sMKI5S3VMbzVMpNuSsL2j3O/dPeMLFj6n4aP
31WAPXxn37lWHKvIGsYrzfGGpA69BxpnP5d0UiMEyJIv6dIOcRKyFhU+746yO8HgZszF+b89J0RN
dga2/cfa0tHbB7uwgAZGyuH1M9b/PaRJsCZ/zPWrx48MaO1Dfi46wV3WlXIiI94PZFX7qx4Zi8no
Qtct6Z8tj4khyGT4rrCpYVfYaqT9BkBHWEN3c37a6dA1FsZD7W8o+iicpG0JHIXzq70YlE7Ia7FJ
oxJk51MF9tlaLl+0+Rs5qSGRx/Xun08HF6h0RXhy/IcP8nwY7DwmGlRY4coA10bmnvvd/GT8HTvd
OF/09A7d15FlEp13R2/fisk++uW20k4WNuazTvjNTAuCIlbu1R1yWXRHFI41YYUEZimYsfayWE/1
9a2X6sjrwqzEl+Ks3lH5muTq9A06t3b4Lz56XL4u7dMkr0RSUN/+db49av4o6nohhpD9oLWrGVgk
xvYPDQ7TqNHm2sHBs3st4FQC4Rl/wUX5lgtUXra9bRUJrR4xAZdfGCHQRBUkD+eIgExd072zDFyS
e0uS/SI0Rv1Kmk93Zqu9qeXcI/NJyiqvWG3WYiudp7wVcNHtfq8zBXONcvbmYqy6VBZinKO0gwut
xpniyxWzXD3MQ5Rqa+7jqBSeEpSwuaOVvaWcJ0Mw7D/PN4u1egBIfx6BneF4xXS7V2Yjc2UA4Bw4
2bTWj7QJpNrYbnwkDLZ9pzmKUyU0qzq2q0t8+T25Pp4ZxMQ0Ohs0bgKc3e+QZ1C5a3oR1WsAMvOu
Zw6CT4WsP7nWj813D9sBABHcxbzMBb/pRFIEGpTZbN8q9/ct6ySXD1gQi30Ck13HQVLz/fHYJnfh
4T5C2RGkCyrCAXMrLGX6OCBy+Vb3qlz4Ng1TVPMr30O4bGxg5bYpVYHM+8ay3WYfJClny23jkxDK
M0sm2BzE0sDvqZYtIW0yIweBv/h0KslnNaJUOr1Z+m9OmGXTWmKcth/WLIDp2iaE4yNk5Bxcye4Z
rKG/prvFQelYtl7LGCVOIhD8mnztrQQuyXgJK6g8kPQLFCLS6h8VcmWwAzfsWtQOrLv7I+qmugfB
gZu35hP23JPSL2BFk8pUjXgXy8RTghvNrTtsiSV8FsgvfI3SWLNAH9hL+YLkFPAungR2I2UaK7y5
DajyWsNC5e6znyVad4GDD7fQ66byeyvTxwDNAI6rdz2WTf1tirje7s7bOlJR2lVyc/eGIszna+yJ
xkwli+GqneHGjzXv8Wg4jubrOSV8jVsRDqzXwvZjMaoTXOUWcg07T2gtA6u4UtWMZx/z+2IGnSTu
pZuaQA1P8fYAxIlferTeTcg+bVE2a8QdyYKdi6jao/DrJ57zcleXrnvhKJog91vj8ZGs28R+30YM
4Desadld4L5ikBRv8kzWrhRc4vO/XxjYc0cZPDv/gzoX7VHsqi6VUpdw3a7VmD2eLZNj4uCEvzsS
3Vi5/HurJv0wLZNQAxz5+vA18tt+GPwm6ZDDdMzDnME7jDB8T1y1R/ou8/pEQOFr+O3DA2CyMobq
ZhFhCLOwfYqSvOnkotp04fudbh85T39fW03SJNALjxPMiMZnxxRhXyRtmaI40vkYiLMGTpgVtrll
TcCceogj0Lof9x/Zsd6FCnDO5C0Rnn2pWGzSBi056In6j4pPWJI92mA3ShYarTPmzQJakASlMOdq
2j2tEUvM9SNPNEed13CM9NIJC04c6zmy3LbnSVKVhggQHumcfb0sArCdF92ivpTvNEreKRPP3cBK
eGOmcKIrmjZ6IeoZctRHtVzz7WH4Tw6ih95VpDVgHcdm4teaZpDY/XpPpejboCu3KftJ+ZE7ihwu
/DbOhBVHDZD+aGmwaXCgPBghGxrAMbSpL4LVB/BS9mx9vK++HB3XsZX6Aw6nz9px7LJI/555hWza
xHPZ++3kF3LMhQdDUkyI4wL/LdF9GyjVjvksWcOYTUC+u/66xIeOTe7NnWVHa2kyNqfkzsRgl0Ay
7WEPkNHpimBaHEEuO6H2udwg9a4ngybTVbVpXTe4Vosh/mbZfkPg23S/xGmDG7wlyKqrTJuxw1R8
gteP/jEyZDzebZfszpfOORvwZhPICycmqyqNFHmbg+vX1FieYKV+P2DHYTAlpQsjsU6uhrOW/mCe
OZZ9GgJ5CnwUgtVavvhAyXWmjViYZmdHg+hocMXp7t8abrRFJpBdv9vDZcRRyzr2k4Lkbw61lO6Q
WACHY+PFHyWfu708r68XSbhpW5as5kA8pITocnJHSyed3UdAV4by8193OBabOeiypHILpF03fVxu
LZ0vE4BrFDRv6Gol7n4DgfwV4PbRlTqI1hcdHRB/thT2pRX7R0udNP3MuplVLBMKJ/PIijfvtFdc
LooVNWOiJB7x2kv8G4RjrUD6RAmcYF+LUmoRqoKzkl/gT0xfNJjhvrqhlIWGldrPDnmdN3ZrJKHF
p22w8Q/XjJXkGky5mLbJnzF2bxUuqYVR+bY55Uge8DJi6rhhXt0cHndsevdk8whEqFbKp/h9QIlZ
e/9Zhq+aDj02Mv8whnGbt3vUk8orfREGMp5ZMEOYoVEd9A6TgeJ41GHnA99z7KBHQLJrY2+BAHR0
tXnEXguZBG6fqoIckDrB8rQeIBQOtBp0cWs5d76wZ47jRY3LVlJYFJUJwD0qY96zn9zqbGQk9C5M
MRNrNnNJRxw8Bxs8gfWHPvZGXQ91FnbNpRNL8l4+xefqvlzyg+XW+cwEFzSfpFGBlYymKX9Gon4s
Ot0LbrTDAp89VZXB1jTGmzGXf6lfiAFK4NmbhCz/803QQ5keO6l4VWDugaOaRfU6FgGwMsNCanB6
FxR1ao0sZ4PrRAexui1E6ignc3B8lpliDl0sypOxMm1VzElxj4WvXhnABK1bzp9lk2bJ2pQ1RGCJ
o7iuuqaN275Kq1i2RM2Qv8LmW1N0x0Yqo+zBnM6Bk1mZSgrvUTz6hZeEzpZ+qMqrDRwMTzDHOJj4
KT48sG3MpIZr6M/vb7QXgpc6Lp1DvJUiRoSHadBJiVLeKeYANW1ra2ESnQyCZb+m5TIAPNpynz9T
tte5div2z6kOILaHRnqwFVEiJYNBB5YdSZLkfEx0uKPgjuL9STosO5BH1vpzhJofRZEx8Y0kNZ1c
MlRfzyxT+dcONQ78IFI6VR01I99rS1X0lPrdJ3WpIQiS2fAMrQHph7fzzJa7YdfQpO7Ca0Bp4PZw
4BAi7aCWKyQGC1S71dDU6H515PdiW4KzApAroDOqUZfgRKq3UoqmD/X3n18mjBVPgs7BKuIIUU4k
if0ep2O8GPxPIJGGINgev6bWrLi7AEf8Y+aieftsuLkZUmKCHEFkT3xCW5ssY+D9P06vVATFjqdU
gAtvchX4EMowESnAcuMv+ejUyLCpu44dLNHwOhQW8NF6NYvjB9dppzQOsc62Zf+1KWykf8osqhjC
yRR+ShbiZJO7SiPz8P27KVt9tg2F6+aFnTMY7KLRd/irLXa9QMkVPV+iG5PgEDsiECNpGgz/ktnK
/OnkfNlGgvS2Ko4SOxobxNIcQ0vO77lVe4DBj9DM26D0L6tCf/UnzAQy31SzkP2uf+rCQCaIhjpX
1+AxV7+5H861G3/QJM+FJQ69I4x3tIz4WGTJdnnuC1ixcHJhzUyng02aodp0ks6MxZtL/BnOpAUN
AoJ5FQMkptH1xBBB+27ogn00r+fLTaJ2tmjuajxUntXQcnAXRCx5l4rWrb+MfNQ+/fB4jDGJDoOw
8QWBfm2ogvFqOGRfIRbZxeFWozmb7yg9ZRthiDgGxBdJOVzTQfYQtfoB04r5iG6BCLamYv6Vnzau
fCiOEbrSxUEdZJC7ZagqSzl9V25RrtfAxW0Vt9jtfopkv9Lu1Josl5BIGQGZbqobXlGxl/e7Aord
1GUB2fTgMX7JQFpPECnRtdsUKWjQP3ErL7FJ4WUXi8kFnkrjOo+dNChheWbq8jPuUWCFBsCJ9ec9
gr8j2irjl9Il5wUgCQu2wZPQTsNgg9ezfFiPfd4Ex7OxxY7CizAjteC+G5c9dTMcxXs4poNmpjlf
bayKbmgOpsjPoklYMzgni3/cMMxnhoSwVj74eNFYNKVoe/vFaMWA+qhX6u0KuZh/6dcMv2j5mc8a
luYXtC+sM55OdeQU55x0hgWtbBlZzTijZxVgQn8YOl0vk5+qn5TttAWVA8KosN4+Y/iJMrQud81I
+Q9qgVP+PFzQoy2DmB1lpmYwEiyp5A753ann6g5uEqaIZhbKXj/69bQdyDnJhq1PeJfofk7Op5DM
gjgIy/Gxa5wcEYQNm83/8aJHDyvLUO97lRcXSFSVcbicNU9/DMu3HP2g70yWIB80jwSwFriIzYAL
nhy5ipa6w411QKXuybGcQinkKELNVSV/OvCjMcMzeKzW/cTv7lGBw5mKhM8/arE/95LUppnyb1kV
HG9dOzKhkgYp8A08o7mvznA/c9ZZGW0S0lY210EOSbk+XDLrPD8MIV7EK+2/xvIbsJ7UlrPT1WK/
DklT+Ndg6934LG0JJ/PwUYtB1n3RClOmZKklfXihoagOyorrqthLgexMadOGhF3ax/eLL7S5FjwO
EB/X4PwawvGG5oOgiJw8QgGx0itZESNyNcbddmxe86BMkP6L+KPUaaB58pWL9f8ZrzbiJMMDuyh/
f6zAkaZJpn/TihSAq5ORWFjTXxYBaMeAiLrufd4sDZw6gMf0iSfB0YtTVmGKfgwdFWuVY06uf3vj
p2PANqpjqqtT8mofiWR44cmTYjJR1sf5BIRWwP3dDQru0RSuAyjl6dp3Qtc/Yl4YM77+v7XCNaYm
2JFqK5CwRryGliLf2b4JqvJRkkLj1kuLo7szV163KfpRnzh0YI9fEsUSH1zmLkBVfwNi/JlN2XG6
sZvZxXF92YN+Aunpw87VxJIQQaIwPjpFZ3vl5S4DUE15eoLx8hwwMRWLW80VUJFVbMw55+jjKG0/
sUkcAqSbex3d5v3AqvVrY2qNIvb+TnZOMgP9xPCqiZiHW5nzIXlZJv8G/M3zaPNLqC7ZutVwnoKv
kNwGtieckB9K0zqXxni481usi8UoFoInQGYeTKCbBnbPptGKwKf+Cr2XFjYvRoxTizZNwwscFhQO
ghYVs8cSLGYFIsopv5e/epWBckHS58SWtxvx5JqPohOZtsQMzu2AeoZwnOD5ph39lqnpH5Ik033T
psTXTLkGv+5i+cruI8HtE/1bMU6Bs4w19QGxAcY65/PSuvTYDRD+r6bfAN0/K53z63X4kjSOBbLx
ks0hX4gdaZj4HPEqvn57PRPR8lNeUl5/2sgaRZLJbkO5jc2cgmqW6y/mnMrNfokImfkuAZ91bfJY
f6Afm7c5PUQqKN1+5xo5X8xZDS1w6FKttHQumGPlp22rKtBX6t82oB2BXRy3k+tzWy/US1s7nnkV
ATadwNnq/Z3yjl5BVIuEoLWqMc8LR8QNBDjXW16LgpPtu95+T0zizykR2NeHuJeGrEteH7dvY3bG
3nwVTA5eWIExwDUiYUjAcB6y5/Y8iGbRAURlxJ8nyoWZiAUrG+LTWff+YEnIST9WXhoMnZpnDpVo
x5s2wRf4HAUgLMZZpe95dQlw2G9DDr5I4LPJRGUklht9jSxWWEb+7VTjdHX2yh+/yG9X9GFnAMDH
bMb45HWRIzPawmW9BSxXDbtvsd5TKptr7B6+ynGSONn/KRJuUnEts7iOudn1W7/1nxVIRqgplaih
sIEjB/Bj2cXjpmjN43E1yhDXQBzPemnpG3hbyWxU2zSMncytMQYlT6iKgyRhW0xxjFggu7uSrICR
LGw3bS++nZP6tWlOQH03LYtdPL2LqwI8zFUaPHPoHJfD5mUPZmnS/9g92q3LSnQWQV7+4QwmhJtj
0J8pHmRNvQXeSgO2dfbo29oUmqS95bmfNAcEbJUUIqdqJV4Iv8VOo57+MgKkhk4RqXyE0CF13yN5
UFE1tCzlEAdb8b289EqDuZDXmO2L63DLGHabqF+JiCQtJ96anmy/UGJuZF2nqNZmf7LMHvpytIao
IPBkTKx6xme/CyNhspzveqTufJ0c3EYzvsQs1MUMhyKFGjTRLhYpXaifFj/B5nzmG53KKDi/VUnG
QJNS+zwTpQvgqMNYOenw3l/s8Zs1FPLd9fr2VAekk3cUyhOFdrw2/XaN3izagTwsXt6UrWiny2Q7
2bxFsHJQbepAW3VC9rfZwMuPLasHcF5XRX3cjdS+cvgZ6jHFWqaLvY1thCGBw8agJ6cQGRr4FeAz
GQl0huOUln2gvB2igEOE87XC5GDOeWkKDHXNc22ZxfKPJjxXIqg0W9VW5n46wa9x7N90NhC0HXKt
i9Kfn5UccwPBbbsrD+xIpX/ZPRjMTIDMvUnp3vxhKcMLWPsO0lHwVV5cP9Kv3Qg2NxGlVpaFzIV8
/n/GemtTSMjqfhftYEUx5fMLlYrHaI4ISx3q+o7FV/aMnSnnoGthOAdgc25RvBk5uGuRyAXL8la8
cmYKxN5q6tVauXUibhqB4aaDxh1pZUNGo8VcwZrITGNNnjIu5k+ALYlC07rnZtBx4RffDp4DpgpH
r3A3bPE5VHhcchuYqYMwG2MQgQsr21Q2canf3PV3yf7ZWdrVf6uhTtKlP1fANSAS1gw3l8OJ6ZHM
tOIkQvG17XblC+FJdnT5aVhxb0gTUsSUa5nA4CmgkqTFG8yVUdc+4ZqBCsnGXwPlcXi566zsXP/n
FJyABwF/expP/fc3Ky+fFx5ayD8/DTL6sDTmPFKPP9/uoXpSFhMLx7Jxg+WIjj9PWE/CJXDl5icQ
JKu056PDDsjOwoJrkJhJCms0QPnd+nQgdcNZ6h4jVwYidTElPeYwJ2ZGT2E1UO5MC/HAhW9VN1mN
JgLRp0PJc5XiWjFEgKks4CxBnQ8n3rYDxkFxoXLR5oYteOMyzN+ljG8yevlKxgcSLMJ7UWg6PdS4
0w1E4/CvC+aDbtZWx7olk2tESWPPIW13iBTMWp373+NMgI/nIS2z9xwmrla6FcJC7IeP9BATHYtp
hxSKec2qG2IZ9s4fEbsFQ1UpyKW9TElTGY95/HL3q/RaX2AjoTsn05HIFf6kPQvsvS7SKRYNC4u7
2HMQ8kcjz6NQb9Yfnynj8tp3/k7Nfc6afMNh0nuqHsJxXYzb9lATTe5iXwk4KxYGT6w56lqTYrPA
xculKGtipIYSrnkGZSFqf4yxIcmM4HEqrlK16c5iixYMgqcoca7ISdZb/UUNMSpmyx7+wdkiaVVP
26l/nLTasfcAKgamcTywt3HTTgB2u0Aita8xRxyLJR0ri0p+Glvqaa0zQ0WZHQbo79FjhO5fv+r5
1BPwHDGlitKPHNr0B0lGF25XfPMliTSnfA75QcQ5Yd6bc3Ed4Mz32ec6ddFnLalTlnFT9AiRJuU0
/G2gh09fDr2iygtGb7xShZ6t83WeZmh6TSWSNjcOb+y0ESDQJ7j8w2aKT1KW9366AlTgEFOW6HP+
/KTDovwzGFWnZGTMjpdP5zXANz0IZCId9jm06ut+9mkgqoLCNIPm88/Pb2vT/YytTroS2+uftLcB
DPRTWx4FJ5EOsMW7CqYdzgS9wbyzBs/ZvbDUjzrL53yQqHXl9V6ra4ft3RRBMD9oqQhVRtSFHL9R
rBo8DD3RQxurJcIRh4lVuthIsnYnRITJyYYv0OuDUUv0+aihu/+0VNLyRdoHN+2iSfC591aZ4K3h
QeDWriR6PWefsLu8I7ktGocgqfZ2D3AtuR22ChfaGEhNoi5JLKqAVieyC2QG48DJFfp0uM+q2vNh
JgFiFBS3CyHeK5/7LNcHj31OyKgPoqChuMIhKUs6lCjj/XKpia6wnnXb1YNuN9RiaEslcCTEkYOg
3+szjzbf9yz7p40YK8kCyDIhiOmZumYLdYasUs1mBCHkK1x5BFIcmg6LCjSpqygqVKXIdH2LOuqK
9p7W5/gYzJ0KclGe5RUBVFxwn7ZMAxe72NlUVyk4NSENCD6bdyvARgfYcDdo86JIcvkIxHT+iP4r
iN759dnVT3RbagxsCCi38KuMd0fUyfC9wrIfule9Z3U6/IyFtsbXUIFUxwDrOkc1HKWksh4EAhgf
JOvOj2QC7mS6Qaf5wlFcgwdHoiCNB67RseS5hmqRytf3o9egmo+EL2TpNEPlujfqbMNUaFLB+PD1
Mvdg3cdz9lKrxS3x36wQvjXl/Vo9/cgTlDDAvKFkUyZkCrR0WmSmFmHSNqu/6m/68eGzWWSAbbAl
plNopqVNTqnKS/mxJOHTsL49/FHQFBhr0fD5mrtWotWd7u5UOTBJx80fYVJA6e+QYJqw3vDqYGXP
KILUQcV9WgxctBCZoMpusAXhJ9wRgdplQwlOz1cnXyC/e4obiibow4ZpsPNhG8C1PMkVqAm8aeWy
COpsvh0TvTDg74DH0AugXtBJVqX+bnCqj12CZszbyAhidYUeKMRYWW6APzSIkTskQSv1wgu4zpXG
1jzRQFSX+/qtSNDgRwW7dyYfa1ZOHuvprthdweh+16dQ2wHh3P7JB7t6XsJrXwoWu72vqCkQMb6v
jWGnP6Ea+79mg5OHJqnDtxMNaiOxHdkLfF43E+Vre+YSs2NuYUE+m6TUHm7ZG/Dq3MyAO4VNdX+g
99BGgdxDmHPvpqpPhuuLfbv1Q6ehO7zMqye9Hn+UqLOY4JkRxh0L8PErpEjidpo1OYwKOXUgkz5d
8RmAUl9em10sQ1ZXDu5r1EBhI3L077tClMXCf/2Eai3KlleAMCPM6gegHg3a9OYwFWcZddL3mkuS
e9J4rVkyzFnA1/d2XRe7gLtVA1GQcVolIJxsxlNvuxXNc1iHB4p6knJexDxZIcJoUTvLHT5sKHT1
xgZm6LAOKLasZfaSfQebhnjYjP2jKqueFc2J14QbvPcqVxpW29M21buYjRWGkNhAhIFzLO4QbGa7
QYDwNE6tgYd6KFtco6C4X1MmrERT0WHTvnn44bea/9FQw7twgAL0PYMg2K6UWams64oMpwJF7vZK
QJzGddOrH/CyDjVRx0x5+niaeq0tDAwv7NKZ21bG4SQwvalS2crOQQ8LULygUvo4HDjxHjtCaB5Y
020r+z49QnlQafeW2EDU8SGdYvuzyepZNRhL+pAuivCUPAl+aiQ6AWGrWJzYKZz8BdUgyAf5JhvK
YwnNVV6NE4y7yyZMStR3A+2K3HQnldc6n3ZpCoVE+H6IwFRrMD89x6YbN3hAz8dc9iaEn1+Z76Nu
wQ1dgdDmYj10QCnx/I5G4dTNGsFRowNTW8yzFn/S5JlNJoU0Ifr8EmMOxw48kGmnXEI8ojqcYTDc
aZZmGXGKy7yahm7NAMGKKsdjAWXjLz04F1rwyDixF5JiQbQvX7ffGBkHjemvuzHn5fUsZfprfSxl
j893QxvVDbTWky9va6Q5HaYczD/9N8jiJZg8oEr5y4VyaSXLWkqsCZvIwDm610iVSfakdV7EG/Fw
nSNVQ2fstUwWzJPtQkSYf0om+Erwgapa0XqNe97DDKlGLHM4+iCNAo9ohNmvBpESZQhgNqHV3MAy
7GhFQHnv/TeigeCh1pfygEW8yJWqAG9WClMQVfFLUmW1iadi8D5T7U0325WABgCbOfc9gDrgW/8h
t6SU+cPYReHsuv71D2fYr5lHppDLVnTJAg3C3lze21YHn2eEc28exextrz3QQ3T8RBv5mYMjvK5e
HgRt3p4vM7c9scYhTLF9Muy6xCVXSUwyMOOVfoi8bc+pt7XsU/msjg8MwUsYSsRsbGo7YIxaxESV
5xfQGxuUO2jwgcRlcWnPUn1x1zK7wzvgtAtoVJJberhKtczHKSGPANHaeZW4YHdxmj4wHVOnFxqp
a+BuY6Mrs2XKtQTlFvqBpKvWcY6L662Y/Bc4EB36ZmKnslObh1/8lKQY+pXoF4vj8KMqB6y3teB2
JjRbsjjXUT/SlTb4Ju1mLveRcH/UwbxgFOVZqumCG7xqVvn8GU/s1pwDgK5yuDBwwnygsEiJ21yk
61PBG5W5NiDvx8LBKu7AQM9SRBSGRR+g2dWmbtPC+KGQSWylE7hgbHhbi5tE55wvHovKDQ+vSpmB
x/p3z1jo8j6f4iagqx1fvpA6nTHz2Md6Oax2uyZBqJO0a/2Zo3W+fo/Hne0zIlEEzH0zG45LBNJF
UPIWIKeaH3asMhsE4OqNJLzgk/mhCRKRIpzXCzezNiGrc9ULZ8XboCf3PJ7UkL5M8HfcegYNdzZK
I8ZxonXZRQlaJRzAKXbiDrePU/vkAk2RsaSgJJ7IERpKm40xw5dC9KIbxZMRgSLJ+1OJC58AgvlM
lJpqo6n9eg1YszB3TLYWQI1fbvGe1dj0ZBcyLIIpdnO1O9x+JvqSpktBIEB9wbIQuUBlSB9u2XLI
MqxDZTiY3yQ8Tx5AsKyQ2j73YqWb/T9GtNxz7m/RW9ImXCzCe8sz1MwGNfsxp5EA34EZ1kBOP3TT
vlefJTiuKIbJNkRBKg+xS8gEgtSAHJ63moBOEa/9B4RAjCfxU0o+O2ya93ZoMEhh1fn+S/oI9JeP
o5We2n4/XaM5R44jllfvKui3sfNPqoPhBYkBEwbgsAuEGbvJ+Vv0Zl2cqzaVzGp4VqDW1ZoHHiYX
7GYvGBAuUuXMF025LW3dXTMJKWvxjdV+4BIg+3rO1kVdjVs1Qi8HiVW8vdD94eBzwjUzaEEOXgqp
tkts05qX4gYXO4goL6sfwT2/k/0fnI58urnjW+3kfl9vKA79rB1Q+YIYtH77Ci4Ux9smqUr6FsZ6
ohICh5/s3wDW9fG+yR8/JshR9IUFcdbxoPO1pAPz47OBOzKIvt6oXYpaBcI6ypqe9FvlnO8xrz3f
WHHiuaa8BV8lPsuPlTWeWAfI7Wau4blwd3xJ/bZIEZK9oWVRi72eWl6yUD3br2BQKImtrb2A9cpj
Xog5CYxGmUxhDIsr2SvJ4m/SawrKRCihdMXBFu0e4ii3D29ArKA6EjJqQtggsY4eJ1fUIPqaWD9z
6TPbf6u6GVSsUdxcGw9SHFdqVw5FPZjSZ/I3r+WdW/ckdg3gLSd/RIOL8UWwHeHVd7mMjA64b4rc
6/bkc3AVcicIUfKWK9hJj7tIrwq6WarWHfLTAHPcgXGlmmhC7R7uXkvGwKm4CfCtXVpK29awpYHR
W8YJwq9FV+PGsAP2dYvNzYiPwD5BjARxjIOUEmBh8AihADE1Oiu0acaHmtTKfHzcjy57Zzr1eAPW
37F/6MfsCxwpCmRI7gFdVVX4L14NTLvkI0eAn77+eVfS4VurGYm5jyb755PQAuo7lGwEbtSGxlUS
N1+LYJiihljBYl97mQtKQB/L7/wbd0N9vSUB54tkzq6sVrcFdIKRTq5KqxA9Hh3oZGuU+ZHQJLkG
pn+zIIJQk0dgu3p7jkHMk6gdt7DV4u/ACfT+gm7mJdozXJhIVYZMmECyr+W20elAkEKmFZoOTsAb
A+L7wL5XC7/uXgT2P5geH/9ostZC7Gm5tKD9S88yJtKTknhChK3WSeDL6nXomoUlbzVP2xE1xSK5
gdTyYgw52braMYlrKAcsx9QPtgdMncrjVYPo8wfy2AiFTsKsHIeiaHK69otxFhX7wsQpSTVTaJpN
YrKAsiRCp5BMxsTYmeoPw0e+4HdC1UxjS3K4X3h3OC50WDdw7duyn+mnDb7bpMtT0F7aTOul/mBs
Ecu/QCoNlYOhutMgptXEwlyRnYO6sxbW6wM+EDywxxo79WjqnzotjByPiTou5rijVZLhZ8+K3K9t
j4soKwQslCFnx7fyY89AQvD2HxInmeg8qdLWJc+MLyWM3Wb+jBjJhd9gzGFzpKwAg+G15CAnyGG1
l2LiK+WQZjuC6SdfFdhwj41QUl1ZP13rIyW8pVSjQzpKEmjX4Ubx2LpaCD9WZcARbRYHTkr22Xck
J8tKAlcRc4uMKqrtkWUFYGloB/8+zNTiM4RZiYM/xeikRuOfDKUt+cxDMjWcyrMw0mBPROWeeAe9
ZF/py+7ouW/fHMbL8l4ElMQPYkch6B7gW5FmCUFTCNCt4gMvXPV1BBWXTZ2xistGvt2LLqrYFqk+
Jaon9EX7Y3+Nam+A/zuKFcOD6sI3D4d57qGv9hJqANOt67+1snBny9GrMgr8a0hq0AK5oaWu1TwP
ZVtpbcYAKhEPQh7RXZCjZvf/t9u++gwB29TSqffQc1tdS5Wzao84Qhd8bS+XHZOCWPjsYLM61Az0
Ue5OEGkQvga5+TkvL4S6ak/vLe+BsPMkA7/1kAp2MhE5cFtsE0/rbBhZgpb+J2yNSW+MjVCZvHok
1BBPmbJfxbUpEvNjwE70dO9JX7FT+xPtE1RIwlItN1SMGlDWB/qR5Eay15BovdnKU9ZrgPjiFKuI
n0PE20r08Ic8txqGi1VKyV+UDTBJIwuTfHiEQjkyrQ2ycc46SyNIvCEdOWQgt1U28qDcjrhHFIFS
+EuUk8SkiPB7wJYQUtle+PxB5aidnxwD4KVmS3Q1wNiOtevF028Ad9xH7Zry/gchSo6wviwFLFaW
EZ0BRgINYud5Cqhs3SoMEEm35QeDMQXZdUFrmFyW1pXeAooWRRllHCY5STTa2ERnxqh9wnRAihww
eXMDrge3v5YTHK0APajLVuc6b/PtIaODl1yEtlUcjr9ejnsPp9oOLQEnWEUdttzIXpr88xAQTKHO
HT9BGSpOudM1k860WaMrkrue4k8Bf9Offf7dmz2SKOPo0X/yay+z+lfcVI/le9dMxTelV0SLEPPe
RnbQJY/h4IYSthS0LVmiDgWU5IVP1i519BkCkaIcHhfUVLv+Di1D6YCYogT5afGsfl702fJPrcNh
8XdfzYTYIhPOhWbVYAc0JR1TcROHTCuAD2IOF7DewpccmTp8z7k41E/OpjcRHE4H05/dWS8Jrp9X
XrsOn16VBo6RLKlXaxhWnuExRl4Cppe0g3kYm+cHgDy9q7AzxE0G47+4kbbcF7wX3txqWID4JOL2
gkjI+OlubR6tIta98ZfD9aLrd6Ib1FkMBYIraviaTS6+urfiqQfdUV31ZgIZyHDFaA5t1k74a1YC
RQoI0kDKqZHElTcve4QMpLlNdsWvPSkQ6XzPVv14J4jue5KbYrO3oLv3QZGbFC4dUpwOhmgKAuRL
gi2c2ghSYZbv578kQzIVQtrABZk0x1vjtk/1My13479nrsiEYwPeCRYpAblb78SBqn7UXWCNCHwi
B6WIl/B8mGsia3BehAIASmu56+8K+eiofpvC78/xpH3QZiIgeXz9Mzp0U+mxZBWfA4WSQigxqy29
nMXIeSdL44szOlVoKc1ww2lsuhgae88bBaUTNGJze7Icqu1XIik3BIJKZO3gxe7jONlwkh64iCRF
gWVoBb6wTwEPnuVGFChvgHXWRO1fPYh2b/K+croMNrUHWS/ksGXkVAwGU0naMKUktgT/9cJYwfVB
q3FgseH4jx2ZAeviqCcZ1fEXarCIOuQ1dguBqTBekJn7phCU6FP9lJojn0e1O+z07Uel7EJVQ5in
aGkwZJYziQG576jjZXoETq8Q0+5sLUpF9qiL2WVjNYs/9rnmnpBcTzEXut7P/LMbgR/94WXk4n8M
15yFLJ5mOQbFkiTGkvcN2eRzIY7ugEZkJyDUosbsMh3C2m38zdjfvrl1mg1vDkJWJuXpuXQtmm1x
VAR41/h97g5dN0+dgGJr2S3tAwICEVPcTFAT5ir/bP3JRaPjJYLglvqJMSMiaSsDN70MGP6oJtvh
CatNj5OftTfbM5go6ATlBZzsc39Ro5gQPv5QIR3vd94qDEty+Kc34p/UqI8mX+jSUKvruToNApZb
us2oeWPQRj4PnetXcGjvjUZYEPkW6l2ksQfmBuNn1znc7TTpFR8CRkzd5yOw/TngekdLEAEktNbS
doQHvzVzvkdkNxkXOZqw+gSl2iym49//4lzVcFUmxP7NvMBz/VwfWQsa8r3Ce+xGckNWuaYQVdsJ
7IoZnWgcO40QXpksmNprqms+yq0OH4mJuRCVsUy2UFMxZpZJlF66vyZ5rJfrCFk85GzJsOzJ6fSy
BNKx/TOGHAdCoGKH3FMwMP6vwbVuoBkJRDFRQWpZnXp/skx4gtz7UAzaSSr2avJCcnaGsZH2Yl23
as/60rtoGIEyu4kQ/mHfsDLNDredlJZuQWw+Bg3dsvGm77T9p6pkEtgJ7UBuK4VfVBB8miJ4/dcU
gyjjfEDnOikJqhHCW7iGCFRxy51VqXI3GS2m5iFKgyIjaZfvlmaFHiYjlq814va25uva4yV3iVkX
ZRlY5jYZom3H2vlyrx4sA23Lje2MtcRDq0vVwU3MHdPQhxX768RFrUxKg3a5CDHNBnEv4Gm2z79v
JYyuihQjCJpIaSBcxuWcIrBp8BrBYWjung2rnXV9U2vpHAI9h7ljZNMUzLlYpqyt0CbTzo0q+Vea
TWOwy1ezWI80plmZeNBG1mMdaM9NUwwZwYPZ8fH/hdSRQd8nSs7RzQr8fbiNYkAVta/AnbZCZnv8
TNfIC6UfDe9hqaGDWWi0ivMfevZstaB0nFylwEaGz9GOiyqA16D9aac6dSnJi681aNrX0cADKcfJ
0V8EHSgARRfJyNThNj0syHwO4l1pWBVAc8S4kHDJjFWYwnK9sajML07qi5763GrU0Wdw/bI+VZPr
Sfz1/nPj1JwJm6SWPgUXla68W17vV2qTuUX0HrqFbUgzkmVQIU6XsSc40XKrsK5Q+XLGqJ2f3KTt
ftDZoUYCh4p34OOyB++F028ARvl3N9qkb+mCi3+d40T3tEE7lq4XYdXdh5drH71I2ZgqFL7fTAmX
Wd3AgLGRtOBaKnP7btQX+oAkYWg/NCfMVZC98YU8UTrRcvQDuS/61XTeUjZIFK7Fha1PowY1yX2b
DUhdZcuvzm79EDEsrga+f7qgB4mRlec3NzMhUQSrFd4ffxhOtehtZ287OTKQ+DwG/fyy4beD0fXs
y6Qn3IfExn46cdfFBCkjqcEaXVPyOY6YvjHkk9UUD2o8Rm50FrdSU8kRMWXolbAPSA3o0++fwboC
H/psJAcpkEQ0bAxC1Oi7d/TAjJKJyxXzSAp3IGxTQWSFDAYdDtFvP0+YiNC+irV72lfIMVmCLJHF
HY6ZjZE5tmhDlom4p4dl+6LP7mnwS4q68BZ9ZNJJ885JFcGBjAT/GbWuHFg2tQszbZzsLaE8d+X6
KOdNEro/o8jLZO/9U+J79S5PUQ0le2pI6Mq+5KpGtaQH775YzYvcqi0HSSrsV6oYMaMPu9wjUDff
ScXQH3Vg8B9mMlioGMd/Q5eWJQvvBAWv9TBbMnC3SAS1y5Zm7yZYuzyXN1BJ3lthz4E7zYvGbxpb
EUh86IbjKZXufQNbuQdZMt5/H4n3JfecRdQlYpz8Rv3RNk/BaYyV6kCV8rQHLDKkJkbf7w9VxrxQ
lNsGbz1jk8vMfeo5xmgYhnhtNtfcdy/83hE2gwTwXr3FxWeytWeHsRw6s+00H31mbyZqUsYeLvxb
rk22wfIFijn9m9Z8tX+DX+toA62AbNwvz+8OSYwZvahRZzCgOgGu1jT/veOxKn9WHLTAslMnneOj
uH6RX6RMHiW9VuZ1JeohwV3zNr6EkzDOAMATZM9X4NQKgVovd2F4X/ME3NXrUVCtOGDfuKLBMoMt
w7QejLVzfRe/zWcejZwT+/kyD+MYdZLTriILgW/PAzIVvidhtAEPxVTRG0jOBh0eivt7vD065EPf
TGtEC+e45sM5QgO8z6Is7Puj3owLknDB73U8ToWeRpENSVL8rJo6c6iJEoakZ1GvZU0gNc2MC/WR
ldG26GRcdzvkZnU383dJw8/hE090Qtbh7KFJTAblDos1lZH6AJgDQ12UlTlKGNHafOkvlz+zwz0v
B4UKwavbxkf3eKZE7VrtK70pW+5Ibxzd3vvFReBy0++e3APuvx1S0z+okuZKzTZySK5joOBeGBqr
+qmOTMdMIhl2Tug5oE0gc4jst6l4jF154Qo+JjBtD0ENjK5Wme0pHlMENrEhhgVVnzPgESjsNB/o
GwBGOomFCMuRJs1UPtyMZlPJ+t3PnH8RLCKlyF+aEDv1kkgxFX18d8H2C6MrEO0d/Sw5QL5vzmt7
v5XebCQTG7OLphPfZ7EWLKYdAR/++uIxaZLoz0i++jcwkILmsblqwzW5TbMQNLPaz4wA9BsNt9tB
KyqqAvbAr1PDF1DH586C7xJT41BZ7Oc8E0C5e/kZm8/H2xlH+8dsrbj/OYVKPYTh58CaF0P/3yLv
2OxxXJvHo/2ius0KNoMo1k8GY/rPSpkpKNdG0yVmr+WxwNX0eO2T2ihPj6iQyG+lmANxhyMEGwI9
/DYu3Cg/mf06UPmHOb2CnJZR/ezko+c1xWL1zQn/PR77kLRnEHVyanpI2vrZQoHPD7qxoxCr3Ezi
XcyVGU5ghICR8Br3+ejXuZzUnCiSGfIM4GPEJViudRVaoSKF2N6MQAyBsym2jyy4KEDeI3mnVE5+
bRaLFWXDe0xaUEUWluiWmFmGGpJ3AFlocDv0eW4kaQhJyMrqn/PKMKhrrfmLYKtKBnLd7HAXXVbC
DgYj6mN6vEpTaixXb7rFql52tBBnOhf83Wxu/jWlPlAawldKvg7oWcYxDgX4IH0ua6CbH5r615O3
X5oDtkI/KxnBdbcS6i2y0cjViOWk65kr5EvvFJ6I+q8pqbPPskmoqqoYE8yQYy1fu4UamoZwC8vX
Pg+13Ukc1wQlOWQ5mtrX32jSx8ArjpbvoYoz1HZsE1po95DBQQYYQVgjQ0zgf3WZ304kS7nRlxjP
fGW3lJX8OkAPBNS0TISB0LMu+JEL1uYrjaWphzE6WB/FRGOYafr55dpycHWt4rhwOBGHiS7joGfd
exZeTgtKLj2q3BiPDhPkbz9AyfdWkE+UIq/FvakO4CCq0TgLh6qhMdLd67uGneCVNrbrO6224pEX
Q5XFotzn4kUXzsRQdfb3a0OdXWAAwWbd7BN6AXK5U2ofOE5diw9qhheGHeG7m3jwZTdxkvL5K19F
SG+ykccoL+emBhX2o+Rny+5ufzJ1VqO5hFpJp1LqeLhwwv0btZKIYKRLHO0glv4IxtQngnsPN/h3
v64RXd8mNe6AFjcpWX4q36i7AZZK7FaES3LeU18AOMyOIj1GD7NHdQP1WTHodMYf5kXe7/3/ANfM
S79+k9Ey9oqzRFHUjiaBRd3rFOiHdTUqDSVapFQrzemQQFe2wNHmhwCI6+ePdwKQbe1/mVLcRcfN
sWlhq1G3yC4/iSHWf37EAIOOFswqTcGG+YoacvlfAcMfuvEHlBDZjUZs4P68DfxxlRL1GH2+wsSu
Xz59Diz+5EFvaqKaOFcQp9RkFqA/Bq0dsYZKC/kDq59nJq/9GSqFgqoxi4BNz/T0G2bh3EV4Xs2z
xemxaLwtHZkKB1ct6mmJLX7/+pGWEE4ICMQgu6IjYzvqg0FwwItWzJ8jifWKfySTdZwwVrjaJcvq
0jPzbtyhLVMv3eZV+GcHf5kWdQLfQoKG95xSxN+nM/rJn1p1YVktNquTaxzaCNrCyaIbhD0nDXst
HmyjBVclOChmsOAA/WwkpXVsi3pZ5ao3FggjM8Fv6JmK+ndnqYN2QbWhCxnut5wPr8wAz5QWLIBZ
MlIREo/TbODiVpyTKjxqS7pDcDjC81g6+PH8xzVh6rdS6Wqi+2XZUiZgaQ+hzP1cTETPpVluSN1q
0KcxfN97xh2Ce7Ery5iwHV4a7E4dnLskLgYXU/gxgpBDmpGLZA9Z+m8AzcRYq4/7UVYomFJMZHl8
lOMhuZDxljIkPI/NWxEy3Zso7uGx9t831ZmSykE6hWNXQBbHl/o9x9vJzqxj49xb0ib6zLpCcoRe
/jtXf470JDemxzQyHMy0LJ+eXrbal8KWCq/BA4yJRlLuHZeguxxFzVEdn6VxHuoKf4IfGuYEWoI6
EPJubrr3xoVOTtoqwF11O8qotZ9o1Dz+oXHhq5e9twrjH721p+2AuY1nJ03MEjouqct0Sp765nAz
AhfCobImBixgdRDpouV6oUWgPEx5GZL06ilCjMwpWQHoRd86mOBOqticwRm+3EfOZAy86cgnIFQn
3QtMorLTIo0RdOfqVEmVX30Pl/isbfclBIWQbIEzPzbadO/kSO6IwWBRQUOu9EVKujQeIh+zXzh5
+N6Pml0Hr9dM3Co5A/eE9zelZZ7QF8V2e/sb9kHAXAXPJ6f94KXXtANNGZlvrksaTc2jU814iZ3z
J2E2ADq/ZnlnkDCPRGmTZT3sMCA+YQI7WTM3dUslIqncECBnge17Kao6hsMDWaDqt4qVuKILp8w1
6auD2B+HhgU4pfG1lmLJHkD3W+cbKz+zvgf7dUXWad+PqPLw5bomCW7RGW5L+dpgLdgnv6Vcoo2q
V0efS+JZSdOEmDVZlXrYdNnIDarcW3LvVnUFr5GtVSoApgapsqdaLHOnDR5mvjrkNgS04c5hNsBB
7rhkWGdONG/wYLGTAGegmaNJU0wKIWHci7V9gVP/fIkukorJA24HM3VXPcHRfW1ytihqAnLrKK3X
WwvKnjl1KJGXupDrDs0Cvgx/s4HxyEMxH0BVG9HdyPyAFPbeMgtCtJoju33SCpsqsqcA9kx9RCmq
peEmTSeeztodI86oSf91WDsbEy0zfI9mYQ+4tOjUA97XHhCkMptGXR5MzDgLpXaCd/SR5hPxCSnN
AjslX2JP9o1Fz9WkWQv377UoGMh+tpoGH9YjrFrqJIVsZ+li3Vpm6cBk/SqXC1VweZcVVqAi0Yfu
O9LWaTG1n15c1D+5aEdtqMY8FrVALVsTRq1hVXFnCVvWShr4sc8vJCzC8rp1ALeVOaFmv64ZxbaP
w5hEOKPYr4CO6JIyJRKqkH0WFEG7LrB3ccMt7HPV/B6hST5GAQWTj7DBI9DWcUotyMQlJ08gsIMn
Y6uPfNzcd07UKH0H6vf55qGXs6QWGyONa413HNMenEztVcu9/TY8F4xPeLgj7J6f48l7bg0ngSG/
JRytJZzR7/OUF8+JRiGS/IHcWinZhT8qxZhArxrXfgLI+biVrfjNkjNMN3f2w3baEwSMQJ74pmwz
jU+lgdImDuX90aGmP4SynrHaGRMUolB6j3As2BCFag+CEbup/0vBkwDw60SFMJP5UvsiMCUKY0An
RDGXTqf4xZ4MpsUb77WrUKKqXbtcCfb3ptyecOW81yzSROf5MmsgwxWVZ9H8p6ISRD5ShLVagdTi
yWxf9U+wzxnrcqJwwjcDgI7ZJpHNKc3lubH780zgWhCkafwSQANlIpGmq9Ya3iE/I5REwu37mK/m
G3kWbbdUsqRgw7Vmz8q4bTYeDZeyHSzyJpMUINAS/cgRLJj7t2LmzlZgbdTd0jfnXMx2JeYLkZkZ
i97MdHbOlv30iqWMCiW2VTdABUza8b2uedIjQkU3qNOQqDFdCS6lo8pN7bdELrBAj8HWcDw9xjLv
gA2OyGvPHB+TEFIfAq8NrUL2tr4Wv+TLwGPDhbjGV5wzhCaW5qeXdNuM4MqdAfT8DSZX70Sie/1p
5JY4jVgAM59v/eZ0bsLyJufkFmvS5JFZIVO3NYKepcBqFsWfbd0Qh5A7cWghxBjNSXp4MoawJiGZ
cAP6G0MhGkMiZjZN/TZl15nmfICvJqFbFY1a5W/bXShwxTdJPDkL7X8kryncJdTnSXiXLS98Nc1x
MROF+NfwBflwmGUBHW3DBcGMYdnwCpE/tvfI1w6aAAQ1l73WvnFUysyqDa1QGOTG2nb06qN+NJlH
WUzBwrleppV/3zupZzclRid1dHOh12xwSGb6SquD8MgW1/e3Q4y3PMaq9Nm6jWBJC//LYf7CjxEj
w/qt2UO/1ayMnl27mDs5e51FrNlLTtdmJX9Y+WCCJChkq8FDKWADHgPCzyY7dVxpPI38GlTcORL7
3f0qhWRCiEkKCfUVx217p1QTW4xS422qPrEIU8Udc4neDP9w7DrVGU7JBTn61no1fE7hXZyRApS+
1oUp4P0bWuSBkt3UuGZdDn1UE5KFxRmUt+82TSXdvCoy4tROTyZ5iw4LkW/3kue8GMBMP0ymP4fd
o32THp+DONbxa7jc+8nRiWSu2ywQH2Wt1Kp9ZaCwIObnxtbFrITwfUBTcBbawD78+ly3Ah8YDaFE
2b2WOvMPYt1B/ctnnF4sxTluPXEU9a7CjaO2lk6dXzB7pdk5YW45b5awAMqwqwZpTp07WRKEBbp+
dyeC3rE9CP5qdJLYEaCNxLRuBs5SNMRvA2TCRm+/K+DeQU6frwOoyqhtBUT6pAe1agnwG2uYiZUW
JCqtnrElfaZbjLYnYiuEopZVQb+WTYFMZET7ZPv2DKxnc1WuoP8wYHQCHEBlFd7qi8r8fH5/URbN
J+PAqMNt0BY7heYXjVCFZYAU4n6ytkortI7IGM1yraYlkZl6YDr+Bc7sXlWkNlTGFmIiI2XkeLFL
CBFR7c7WFNsNsyY8aRVgcnZ18L5XyHbKwjgSqX4Tgh6cf+OXwaVCkEnrZd7qA8pZGR7bN7hUvrOA
fpW7gJBS0ioDU1KQOCj8UY3Chdg5NC+gvbHVIVXjW/EaJNojPHGfi4Qtd7EGEi5GzI0Zn85xfbip
PdcWI0HjiRljdb16uPVnBFdOkQYs63JEwADZncfz15LVjRuq28dqfWPk+pTxgytrQr/anSoqv0XH
e0i1Zhh2+w3itBYa5pcGL4cVvfvXBk0gAoaM9yq+Ry4UL+kmnUjKupvg9gqIrWunzPzXN6fG/L9E
o8i1kYq4eUXTsCtyN4pZ+api1ONS9QaZSI6fgZwCm145uNju+3qjxqlH8blt6qL1LUaXLjgYDIKd
iVlz6g2yrXHqDuxA8XJo4YQ3vQtsWAftYPRk3+UtzAYAU3911PJ2AzkK6Q3WMCpmRRaNdXLIQPve
D41ptpZYvcCxDgsq+UEDoVp7AYrhxsICqGXH3dj9h6OG4s6GCWjpNv1S7iN9hgCbN50Qp27mPIsg
LEI7CA03cfg1NuFpeYFYOZiGit9eYAYAKNaePHsVaqDVNapZkA1+PDh+5CSsqm6wpeVVtlcssK5I
ewTm8S466rqpqJM/tIu7xgW/6AhQYvretsQEcVQRv49kJ/nNaz0V/gJtWsa4vmOacCUFKgKcskv4
VehZZ5ls69nH+UJrq+foD3ZsCub9ufrYdUF1RvpAwa7mTbI2u/jvkNVzyNU0/LvkuoQUSk8P5lrA
nrPEQbBSRXCrutWKQpp42v4qHLN/9plaPYngai0076s0nFi/1eqj0Kmc9SaexSh0faaUVbuA/Lqb
F12PVJ9gLjBvixneOvLGDeZQqfT8Hi7qGMMpuRgRXprrTR57B6H3TLkcvpuVAafWMF09NOEGtHBv
xfekp+dQJf3W2bWWsE1nD4rst0CRldA2A+W1E4Lb0dJHOGxbxvwWwy+r/0OHtMH/WO4sxUF8GKOy
uM1W/IuEquirGJmi8WWOdBYJn+AtDoe0uf+RA6ZPbBXYgwXDyHmg7IXbUptwgQ7gYr1LVZDzEAQ1
yLmASV9NxRT4R97ortrClDJxQuFRAdtXWiEUZKRJ/uW2poYzgoU5IPfZrMqX+iyFU4NiVmqDEG7D
F6VEQKK1VpGkXxgtTGQr4GT7q/13UrmWmr3R0WkE45xPoh8LFPMtc+u4wFOPzX8mN4/l1z09fY8F
s3NeiyyTXytgwXmmUZmyX1mhsEt0LEElv76XJ074J5miMmkbRt8eom5UOd07PitZMSgX5ZWG7+0u
Od78TFbejQ3WKlAFCgBYA1FrkjXm6GBbtKhPdwFFD2o/U4jQgxfuL/I0f0daZGdmtwakBGnAAbiF
KWmVa0OXzA7Mslqa4rIcFZJbHL/HSC9AS2WD6g54gQU8huYbExhIlmIeB/DCIDFRHSUybuYoHi7h
vYJ8lsjmTQukrnVYxIiwbW9dxRA6IcWhUFIzFbMVVSI6QW3oRF6NptOpbhMbuj8d3xV5/JlVc0jj
GYLSSvX2jEjPOpIjg85I8UWNVm2p9JDdAu9BP9f4vycoUMmAytxrzNnekQ52SiFxWTluSiJO+adW
1q2wcVDQCYSX7QL8xQX8WID9UFnE5sXlByuFHVSvKCx6xg/oGKPmMy/EXsJz6wz+jI1udA+bbPCl
WCkNxbf+/tg2N24K4qh6Lj5q88p8Ca/Ow2O5uQh/DT55oxtGaUZZOsbUCwmNk1GbZjWflZNc4mNb
8HAKh9oMnffecmXLkvx+qzo3WPS8dOzSASTQ+qVq+l1cogwa/dBFJlqlxavofwvJAyFgQSEA5Gj8
F45blbmOG1FPQ89dZpnLyl+DAm6L88PSeDVhS6Z0YcGsiYba/sIz5KUmmZH4NV+I+Mic7eXIJz1V
3vDUIin41PmxjdXIxSzZ+M00cwwhtOkwQCRjQf5caxamejngePyhx98ArhmmoL1puXTGl4cgwvgU
Hfx1HI95Z+qpzxfT/lo3EzKsI+rSaBmXJKA313p5XrR3umYtP4rl5oy7sGrlNSglCHyZxHN8ZazV
bMfCE6ebLLM8+xDSOV/wDcYo20vRzgsdeYzkzub4WrgS7EYC/mHHymNWKjdn5WfUZe9E2x8HoxOf
Sip0423NIsUhqypAKZfn6gfWq9dlNSGQ0V3+T2ftOaPlL9dUz4dZNAC5RLpNEkRPcAmOPjk7UREu
wb59cqB7Mg3h/4pt7ZRKNi002fYSYgfcpCDCVHjq/ufULkDUlIZPDaIJM1ybM3MBKn1tEGhawMYW
zCmEbeqF+z8YEykbQP6XRF2169fH+rxI7ih4FQWs3aQUfLvXeTPgNsTTBQnTs28VVei7f54FS/In
zEiEySUMXSU8VpYI76kRhKxHz3aFQFDO4mwJeDYf3TX/aq83U7HAbBD75a/nvFG1LEjPT8BuNrYk
x4N7uFBfyQatyk4Yrh3DflkvdNH67K9fg5MuBW2/hovXkqw1Aj3vC7cKLB1MAoCL4aBwLnahChrj
Aczfr9hyLY5yyaB4DvYgoOKS8XY6u4bafNqtATWHDlq/0MByuX/pdUOCn7l4BCkpd6PemD/fkpz/
ChSp0vgN9ZxfNNvor2RcylUwPRtg4x2uQllgjKPD5OXTR2tD+0HOIZZk/vGB/EE+lxgH6e72OIsa
DlpmgfXnsKjnEyW+2yr/5CJiJx3EDqoJBV8F9beIMrALwk79oBvxWdc4zJt+X8JkLfSBSuSNguND
KUk26ANTFdxrYd/q1ZbxQ6Vc/jZDEnwX+GX9M8KAHd6Ea/Lv98CyyfIRLVgnIyumDOdV5J2sdoNP
g3X25ZIO5R9sR9rYftCPMP13mutnBzdWVTfl4FWwbN4ePDN4UcEw1OFiqwYV82FwFd3stQEPlpk7
U0wm5Ey259rqXpu/+QQXNOXfn5ILO5ZM+M7XSS0HnAbGHPB1GQx7EJ+UDJJwbxHbOEEN8yFpKRnl
bQ0Ske/AWdA4MhAMN+VJ4XzD+h29ugN9aXQjDQO73BqHYGDrEJ8yvUDtthno2T47lMe/1N/kCjt4
92b0nkxB725KB0KZAt48VEKTqNg5qcR8hLpjQxN+virvxhnCVuCppATU9P6h+IfqYNrQOzil9dWZ
3a2EYz81YGgI+h3+wZWRDCNXWc4tSgi0pAp/hVBPa5VjYDkDXOGqs4Fj3VeVchnFE9VoHsrnJzIJ
M0k9nu8ns77lXcMsVqm0ramrS4jEBFy2wPohICdVMuYp+oLgRB/jD2QVUfHUxQ5xlyKr301M6vtt
UV/vJ4GeEk0Zuogh2dd9y6Tu2FwR2BIbhBSWt82MyjWeAl/O7BS/fRhB55IfXLhG78QtZ5rOmvSQ
o89u2d/1O3b/ZLM0r9izsq7SesHU9AJJ6ZheEtfC7WuNvaic8J0p97WYOaOzh6sb7SpcLLkCt0Cb
7EKl1nlGmj3KCM46g+XdEnCMcNtYk8YJQ6qxKztbEhRZaSSW3jzqvjYiSuZzY0k3J+ey21dYV6B1
W79nwOhd2YhbysoK2lzCtgCS4HMh92p4jns1+W/B8U7J4orBsnV1fzDW3KK03jG4QPNgRpw5bEGz
j8YW6pg2OF+2byyrjN4w10aytxmWwbX1OO9Bs5Hx1HCkgUZVKtkr+uAZFyjsACdcVz2/LMh893lD
BadJZgKsHdtltQYEiNVfoCAsEpereTGTOpz6x/mUkDJMS1HAvyc0DTtrMHShtX3Xge5h574Xv8xf
8DS1tTeyFj3D+9JWOXHBKHKvsNc08pkWzde45wlNWS+UnFs9/fs6GJpccW+QFhSbQVT6r1MHKM3z
ILXoqotCxtPRDTv4Ww/AY45nKM7VjNqWqxEDzkNN4javQ6z2Qe4e9sWHDLnsY48HFQbH5MOmdxtE
pNPxys4H7y/AMe1uT/EkCr6qc/JOjsM0uD2hC+WWknrZxzBQAMh6kLIqjOcmbVHW9Sl4P7C4TPGo
/MsMJyjoB9oNCpCyENM/NU83wE2FQDQRYLZtTQifnmon1SRQNzCeHPHkYsMrj02CRo+YcbdEakwe
JSdUPSJ2Zdj2nzgtGDDNi0t08M6AN4npL2N+KaeOVgp1J3CC+Lskz9M0zpdvwkRPnbozG4WfqS8c
Tk++ooiyGIDkUXTjScluHjr0jVs0wlc5/L5mExavQPLlpnW10MiztsXCitTEhnKQ2Jn3JfCgUl1G
W4tSXqAzi2E3LbGXxy2mpxvKq7gHC/bKNGCbMmx1T39yIyi0BEqY6Ycv+OaRf8ZMpH7yMpwqyBPm
y0I2xW4J/IgbRGzWxOiXWNljvaJab06UJI/Rrrtd4wTbsCvCwrOkk4J7fCpAI5hphevEGhBnSAzK
BtWczERs8JTv8bRiuPP2w38uzuwmuEjMrn/ZvmhMIQAjCrd8VaHvFDRicisjr/5fxs22AgrItrxP
Ij6RB8bLRuz46KXMAa+vN/j/d2JWdeqMffKpyYOGD9WqTXItafn+R25887qNbTsbDV6zvLItjVVr
fAnEssueZEuRpTNokOiVPXP+3V0egrsDe9ptu78SI2hfwS97LrrFOEFvivNcb/4kkeoL3wgLlRgW
BjexzK6q1xhO+F4zguqjJapj6+nH80S9OOj5M7rhxBFfo9Ush4Y4yAGD8sUa+xbGd3bnPUisr+jv
XwOY5aNSPZj0lmB5GaGl9d1G6GjH364XIsdUoFxWxEYdnU1ooctYU8OtKhUA28crht6xEcXLcktr
bikHQqFbVx3dXArZtGNqZSnmDDx8YtiNzas0V0FvCdt6sJ4l0VmbtD8ezOefb9hElx3l7AYa0dT3
0mEEI8pqKh4mH/6ClVpNjGyYwfbd5snLfbK/fRDfUQC1DFhpLulgrEm33kirDMs5bcyXaqnhnxXu
o6SNVnYrlbmdet8qPMg2trc7oKU7QNfDWb93b/bYGc3Z6COXRJLD3jCYongF6SZPZPRzthmXQJ1u
2qZx2hZWs7C5Dpkv7nRQDPIVHmcxLjz/PGm9Mx+ZMESuk7D7OHKQ1vaKY6LMaylTaos/gF3pM/rC
80bG3LN/kyJ8mZ89rNIyTF2SH3fjmupRP+lspHocGbM4w+8iu2IGMdZ3meu47ACjAtr5pUt1MLgb
n32pGMcv+h1fmFGM62r1QizZ7XUMvgQ2w6zXzplVEBG4/tZe16GVAsznpiQyHqYnTXtBpqqxlrmT
zmmQ2jNpkeo7Xgx2rRMyKIy4koPW0ft+qrrxMscTqi4cUKdl2bAyjsIqiicdjWuTrlB5PLqDRmBe
fd95x8fWEOo8qEYI0cP/I8N1HdDhmcmAnJ4d1TY9YcrF5CXxaQxtz/IRXytuQmMEuIozZO5SUEEg
XbLbunWywReSNpP6yPLRtlovRIzdRqeovaB3+F0hV5MIcNbdEoGWrsPG4WJGF5Yc56Me419e0wfa
E92gOgHsik02UY4b2+A4+BOlLiOmilo1SAYBeAW5SaazjtHsXCfx6NaReVbYxWYnaFME6Bn41gm8
Sr51OYQmF/53nhravHIMpYN/G0NxtESN+oK+xa2b16z9c4gx03pk7EYwJyDOUjLzlwXRRvh/6aq5
v+DOCqKStgh4kj+iY0jd4xb7ZhMUTryCvKGidMk7dZ4jqXihHuFdZJwv2KkY7UcoIImLCJz4Oehc
Vmb+zQ90wxIBYFAObJEnnqkDpU7GP9hSH1ZIJjc6YXlqYQgWPNmHPYElxMN3ieJmFW9zkSFP2zlH
sE/5npJmTh8Gv6MElfwmZtMS2XX6R06spdqfHrjyPRqXtRS6W3inE/ab4ivPJRGOE+j4ggMOh4oT
rQUK4DrtKJAlFsKxocy3/+yt6E1Fn3mESBDKXMO74oxNOZGk2sxoMV6GFkypJuPvzrbAmelp4sBn
xbgvZf3pbGjNt7hhsEOjgPoFZUxMhMc9YrymEXneg7fyCu6IXrFn3XjjMCzXI9B4Uak1hAbDyXf+
0uRChI5fIffczYNthaJ9kstywPN1gwk97DbgwWINBd2RdMEmD+Idyga+sUAiGHKVFD8UE5ePGb70
EH+oTtq4xkIHm5a97YuhCGLQ6ymIKiooO160Rr1VjR5hnUonSHv77Gfn0wMtWYqG7nB1t4F9XgVO
y2NWha7dxrWnMD/0BBqoy0RxPpb0ns9pfln0ZztNEPbe6qwDswfE8yreYpTK2BUQwQnatHwvU6kR
Kx+C3D1Sz7wLZ4G4o5KOjgsYE5UZB1TiKEtmkxZYqLidrZL7UrUdFmwsoBuiApbOq8tOsghq8jsM
cCingNUAy6Lljp7HTH26GNomjib/T9e1v3AemZpVybl524jAQrDQr9L5+SZzEyldTlRB41M4Nwxd
oHOZU0Mc5zlMMPE6P4QK4jODmy2O4rVcQUeKa9Pyk+TIiKwnWwdacMpxBXTrSzyBrqqVWCny6DrT
tSqOFRL/HizLQDKM1vQnIxVTuEstklqHcHbJfzCWyExh9xyxc9L/UoTz/dZ8FKfBDIbNom335cel
YN553ytC5msI/WScbpFw+ob2A9jonz8VofHTn37SyF7imkKE47JR0y360KB8gcbBWyiJUidmH7fO
LhPGfBAQXcj7roSz2HFc9b1tD5wEefoBsS8cWN7qROGgTVOpuRZThLQnDe1/fR0M6nJaeuoXT+cj
CCr22mSJT0wNOigzMm22L+tNl8qr/Qjtb2GfWwK/e1JF++7Y2SPrgWmBBgwzcLz26q6BmbsQl6Lv
aADqzqumbsMn0XyhXVupazIIq2klo7ElrfMsMip4XHcDtF6HWON/wXhSt3yp0puHuSop5D+GoO2d
Mdr+jL/9CNC3PmFUWJgD+MbcQ1Sg3/osazzEYMeQ08BuuRfZTPMOjOfZFihiPuGFlwybkBEZOGpa
jHPQIOHlJymU4/vTCnuNSx1OiC8IhsqGngXyzoYez7rUyhfK/Gt07IUuVr/Djc/GQod4z91BL5fL
giYBtRKjRSETMYKmYMrvzt2Icw+wUGsSK0tVywgNkqerPM49aHszu6Xitock7zWjrOl2/6eFFhCc
9cwF08nN+JMiHIj5xVEDYChfsz3/g1EqbtAFEC8N/BVk8YAy4v7HJsRWYmwcWCmDaVI1G3JVaZXf
8+1MY3Z4dMLsfeT1VC2U12HTU/MDMHLi52cIpQemWrmipgBfBpQ3M6lYhcjDtBTXBx8aINN4JKpL
ZANpi0VAO/xSDgpyUieIIQfqhGhMGUGA/WZsBxtNNAU2B1B40xTeKfwDtjs0b9W9wHup4/XdE4/a
hikKRaSMxOL8FMZJt64yfidCCozqMUE5iHrwlp8RV+76jtCHF6dJ1iodYLbZJVD3q4oN/Lgwcey5
IF4bgx7fH/cqkeYWKTt5RHdCY6OxGRL26M2oLKlwU6lp5S7q+evvfa036zqrmJqUcCsUs0SjyjQH
Pgeo/MTpP++7nGcw+o33Lip1efgX6v078LXLRZHBc+jafaQoi/hWeROEQ2zSoXpxggCisiBUnD09
AMRhhJCy7lXg93LJ329y2S7nkxS3gbG3nZMXGffu13ihLc/bt0C+jpFoPyVnknmgcvoGtORh8r2s
Ja9MDBRHNDQxYVJM3oGzvraPF2Pr0DBK1QYZpMbHOcVL6uKubTdfHKNgphZPfTgvvgS0uwkyP6ET
MUAcYvyDLO0iZWXgqS2b6Izis4+uTZ3lVVeY1mdpbpJEYpAwMsg/OhDhyGXoEmEkiIVvOJxY7TbZ
J/4J7J3ELrFGDm7U+1W4olH0La3FaYPZpjp5fF9fsDjHDEWJb+XPH6N2vVRw21duhGRiCKrdFWFO
oDgiyN/sSFAyoJpLdkKv35pyKEbpX4zzFCzyRzlFUDuSHZOSxuAA02MYMg10SpF5lRGFLbQVVut4
RBhGBssu7VHxWsoHufJwftafKV6CfY8y05a9YtvwT0zgKwSRdGTHdbffiaoTjn7B9UfgKyMEttuu
KZm62OoSBZrIB0UOMNiF6WHC2wWUzAamWmtvV0flhEjHVQUw6a9lfOoJXVOUD5BkFy5YBprhVY08
1V9+K9Qfr69Zw5cr9okdjiWmNSDfb9D2mkbFqhjzzsOZFyrlC+Lpc1lVjHQDGQqvcVBwiSJDM+nI
F14LWEPS2Gn2Rba2fcdySvJ87drkgrwNCbdanemtca81xDCX8r637kd/tvK6deQ93iuRwhrYVyn5
DqU0/EkbZ0KJB6lCGW7h77t+FdmGqeVVyA6iyLD7IK3GBzjOhg+GXhk4yuA2ixK7s3oYHgyoNuzs
A0x6ay3mj1WVrVOc85q9UY7rj6+VhIKYBm2EeRGPO+ZV0jwE1cwKMv0McZBmHPTuvy8xC6yeTY+t
kokRmTuNGkmT14QtgQn1aUJNeQBeDfDpz49Eo4fycj2GUa+oVTv+mAUrrCkg1BiWPfsG+jxIEvCa
ZDVJa5nwmmrViuLgXi6JeyA8ZdNzaH39G1xq8RpE7eO98ggZtTxcc97opdRlGg2VO5m2zsbDxt5v
ONfVanej1YeJZd+V40Viq/TpAxR/1L49SYfW00W5mL5X5fdS4s3oBqghcUPUZG+dZE0NesZgbZjo
SOVVq/e5Jz3rUxoakGPmVfQ49j2brIJ8D/8EsyhS7WPj863RauTAUTcGVIVasS5trzu2nPbOhpps
gIZZBbZjxTyOuFaq8kS1GwvbgENRyDTNdRnkupCQTGzt4Uom56viszMHKt3K1mUvpMYx7CYtvj8s
BLV9cxgh9g4b+1V3tx8cYz8++blYBrZyjkBRh67CGF5rtm6gb8pkOHLCspt9eR9UhCsXZPPJVwow
dilg1kFGvsPJe2h1hwCPm2R2Q2rm4SAfu//gFIkOMbJ8Jezjndg+9DABEMqlWb4W40xhZIZZMsKl
6EeM2g1sZ/oVehFOt7XgQoS36MLzdKh7HRwnuWxJ1JCdTOFh3ks8FqM+UYz+G/ns7Cx8Gfj6rcWZ
PpuCGRtpLznZwl5UPrGmP8qF0cuhXjcpnWG6/3HPh+GpG+cRwyiP26whqdT4TzGPJQuGIpna7V1a
96d6UqslVP8l8xK8JzMZqKAafuY6mgTrx1E54g+uEq3zBDncIekm9GxkMuDh9XpANVqbP4eC6MCq
1Ee4CiuYaRw3MkNKDaG+MM33TBM6Kxho8RBWzYHHg/MH6YOo0Bv/sRhsLvBf9eHGxlOh2r52Ho96
x0cBqjqoK2sFcXTC7iBOsd9uml2cbmZMExjYGP3B+5bQzrOQxqoiUS1EAvxU0Om0EgcRTP2pmflm
8izgsY28RRz5xqmhHYP5Q21enEixc91yGkDiv8IH4U6AVxjfUlG8t3SDox2N7OuIfN4tcgpDYdC2
5XTF1Z9lEPET8ZH+CBke97fiJnqW+taktro13Yt6Rp5+kztct7FeiCa5gk6eH4UFDHDB2qf4sIvU
DgYmdEi1+HgVnMLi1d40VVToYwTCdOM7la3sAX1YNmhCM0tMwaY+UfKIawbt4taZ/XT7kLuJzRD+
Ul3UmPzkOOzuWNQNlMaEKAJa/3saMpeOD/XAUuOPYddPYcIiOgxPBPgU/WwJK/IWZdNy4ST+XnMr
HELqqZCAtkvHkGMpNYq3tNcIIBL+9GphRr0/4rBJJD//2THvYJ2CKlPxUf41QgY9MV5y9LI+OJGO
WKgOBhLEs+HAr/qugpJExWaNbJdhj1+9juP3H2JRIVE0vLd6SkEwvkwsEzuh6TRetGLPPPAHlABb
QOiWmbj2dWmUoD6UIplAcpGg3kj5s69m+gfZRMUjfk4ih0i+c+o/5TxcYGBZMIzT1fF0tC6W0p8k
fY+swlv/9ex3ft/ibzPBMXMWKdWhnHMNdQuumNOdW0k2302uHeggylj8r0dy0IbOVn1q1ITsTj0g
bVikgh4Grmuz8fpSVFj7oBXDjiDRmN51e6XVPC0PvbxuUA7oYCT5KhSSVEvJ+i2ILtd8oUDJ/T1q
4Bz8cf5YOFXjhJ8WAfqwZp/TDRbpOdwbKSdQsfE3uVqyvYLOR1Troiz+4mTWOXwfiM1lpAfQUWWg
xDiNTDFRWwxLG79LLpiWl8EauOszG8UARdKCoLufhsuLRtFev+fE1T/7Mo0DANxmthdCYHMF8O2N
obhbd5ze0SvuAbZDMgLzTa/cxrxLsQzG12ujDTADaWK+bilUUUG8tr0Rtmf66TlNRL2kon7t3kcp
47Cqy6U0vzZw87MN7euUw3il87KTrzMkvoMcvF8yKLOiXIa1aeylBUxldwFmYMWjoj46uQ6frGcd
PKp0M2U8mqiAZtCjCD7hhD9tddlOIWnjUHZ1JObLbXlV89wUKZhEUnCsS9+na7XOqLWs1p9kZSbE
sbBHGzJL/WbVgyuA2m79yo4qnLL5FyeQT0wZWOCyEcNets/k04QocG7qbCB9etsn0Esy1l5Kfb69
AlIbrEYDED3SxllXNovKo2n0WAod/qGJOJ6ngoyoJzolLIJ6lsbDhe268Jhox6GGCa0Guc3whDwp
YJSvr3fKjy9iRdHNwCPU2MZ3QC2xiYzWb4REmCmZHis6KvqX6iaGF61jyPZ7YIM9EtGmIuVMB/WH
KefmZziFpLmVDRYdm4HwexzZUVTdUiaBjhKZtK69JyGlpEV2fcCQmGlY3rVuWHwPTSJG9I3UXZmp
vN8SCFFR22PS872Rat/+56W6/dYfws+yfdDBTMVAo5qmXxUJIx2vVfN/HxuuSxyoaUD3mfNQEmL/
amgeFNS4UQd4Guv72M7yrVDq43/0+ktu+lUSTCr+fznj8GbXbMVYJGmk+6w8vRWWza36j2pfOUEY
yqTaLnlUErYne31+MFN0T/D3D3BCe6BcJ3C9lo53FrKiIeB25+7sa6bHLEMQcYa42tAWgNhq9MCy
Vr4xe92JIUInlgZAdyELiIINRJV3RdpA5ZDaam3emDZhxL4816j1VdaLBNpg5p75sSIhzbIBUrL+
swrqmofJPchy+Za2rBya2A37v5B2gHjiOiEQTWdzMXBKXpyKxuw1FFTxtcqfHC2IPACeVcxSYuq8
tJCKDzk6Xs9h1xGvr2yBI0kjAdFlNHiilV07ESq+4kv7d2G5yfJjJp43TaJhXoKD7VV7XDLjs+ba
MnO2iyw6lGmnTG4eCZd0kX6WmsPlVw2apmvcBL2B/k/B8clnZ2kTBltJFRCuQ3ilEjWcKX9Oj7j9
6P2evNT7SLSPfPYs4cqBB+Rl3CP6/2dXAeaf9+jKF8ijwaUJortHUoHkgU5V3VyjrMp4UE9sxG+M
H0hPkBGQTH6oDUrIllP7jOUkjUPBG9sM6LkJ1WVNz5f/9ud1KREbh2Ro4mDXZX0sRKUg/S9oSvR5
q8j/9/CjLQxdgtc8COvS9yhAbzuuMb41/IG43WQ1B2uBsPrGM2n8RboSboZIbJFurknfWcxHwSex
GeIwAfe5VM+60UWjNMO7fqlEisGCK+2wdo4b7afRMHbbcaciSXFu78YWQ6YDW5ocJSbZO2UVhnw9
VCLDBnK6S6y8LfMuuXiQE61PUydEgtryeUW0rEm3HqzEEBY+Mu6e3uhctLZ+p/xCJSEk9gsTpQs8
/eC+6dw4HLk74UNvJBCM/I7ObGu/9LE3cECQhaAIMWoDA/EtPVQy/tYkQNwxA7QZIbLdcIdPkyTW
7c4IfhY5biR+EADT88ut+OFvadC49iTUoDWA8sS236ezrM5+q5CztAKLEQw5ZqAjSVtEK+f5Sree
dfJrRJ/2+qI0Bqwxfy+QqSs7O4DaoehHWJrgivHQrh6aGB/9q3EADAzFOBFxLCJ4133sIagtWXbx
r4XDFWYxdKoAM/4QtQfDoGIRcIDqWKnq+FXWbgx5PsZMwuUjjbAbhAJ4BmKGGQ1fNB/M1xuJ4j7f
jz1t0jJeEf6+FdtY4Rr0558YJZDxqh63nGH/gXRRkgu+s30eWVCbsgKzOBy6ATTWDyxEIzLscjHb
QYtXh/ttnBcjPiGt2oUZcQyt+5/UqwbF45j+hVurdhoWloB8mo6c9cWsOgNr7//moxEly3XAzQnt
+jpE3PULvFHEZBariDUGuG/AY4xMQ+WJIeOGfvqegKc84inaHa1jwV/ZlCY+MYdboYdxl3hzsI0S
/kXRHgDIJT8irtccn+6pkHzQpQYb/PDmGVn64UW/KwKcTn+Ba7nx8GHuVTgYopBryotVxsOUrFkw
bcbLPrn43o8XNhElhiBruNb2FNsuWhXRWsRCSOItcCSY39aVpeyGC/Xr7/NcZd/+608A7I+UBUTi
iMSYZ5ipIZ57B1tJHvxpwy+pD2LRj7euqoOdcZHOGrDr64ZNyljOjEPkBiWAxLHCxY9lecHgO0sD
RSt+duMTn3mn2cfDIdc/y58ljKIKVGrDHGVkpJLxOd+U5P6CylKQXp9r4uRT5JpDm36xqZoT/fiN
UVYgMqkZIGxku/V01zR+ddcz4+ZTrLNL3TNTmnLiDl3bRSc9T3L+oeb3UfCEII3vHAvWnZcZ9G54
IakSjObRTGgeBbG4a6R+5IKE/brjIycVriR3qt9g7XK8fN1vu94k3mVDgH1EPxXv89O8bAfgBIHI
UA6ihj9Il30aa3ocL2mGX76+DrAr3D7UhPgKktsVJuIcFPlczqyGXSIlYXg3OtXAjmz8f21lFMJ1
dAnt8u5j++K4BxIobFI51Tax8ab2PggkHoWNV9dlnWaDQ227PuMVTIctD4Va6HBI0op0m+MecMCc
yw3CVHdI8I0K+tVhKP4ZlQQmGb3OLHp4LxBJGPIVUk5UFdfoweypG/p9X9vn7h3gZJSn8pak7DZs
d1B9sUOaL/N7hWchulmQQSH9ZrC/kBsmMIVxSprqccPBqmFO529Ob3UM95Piwg3KCDNhv48fkKEa
A2r9oT6NAZcts4YMGYv+qlOmEtyKGYNoBh8Z51jo+75L4dJnCdymtzTINJ5z+V2LsT5pTmLhpuis
UXLv+MkIlkpT2QwJJltF9+6xoiuGPvQw+vCCSOatzk7fW2/uD+GqhEiQ5ECK4VI9qQB2icys65B6
G9Uy4MKJgHWPexhXkAavFbSVm/HED+Ha8kBxqdbMbVZT1gQzHtkepZoCmybq6oMqOnNU+RHaJYBW
x02uFfKH1LUMv5awQZFZEPjtxRNSAknf0Oe0CVWGc8FKIXgd2Rjm7snKorYuTQq9jXIsv351s83W
WK0iMgh4gEVebBbWyzxcUL6xvQUy7FjkovPY6mOKW/OrnIBJbBM9WiTmFn8t83765hET7oihH25S
SN0HjqSxYRpqOXbrkWgSb2h0k8giBoYYT6k7TwNldwluzWlBEGybsDmBZb30h7HgyRM+6fXjhxeh
lWKObe6GsljjrgKUu7CcdraV1fUO/uCpyGoIWV80T8IdwrDVPURXzev2+Hy2vBKrPNt8jTGMWBTE
yU7uJ+Iy1zA7AVrc90p4pLvhVuYOLlXXi55g9aOf5Bl+R4qWSPfWZa2IACGmUtgD9I0KTuvDiNBY
LI0bNX5ovSnJf4t2l6WREVwP1AKazHYM192ZllbrausJ5qoEp+sTbeWDeOcJhb2L1r2gql2EeRvg
MonDXQe84tby0ofxyX0sPqCaQNdrFjtLslHrH4CsQ7vV7si9C86MbmNVCEZZrJ46/fEfHueEr4+S
MnhTsAp3N1GuUbZ8n9aARDcwz0+j1+0fmzeTDAZ2Tdx4rn1Z+x0EjEBwINjqLXjpVJagzhILdVZb
w6oD34SRuLtTn8YlrEh84T7kwvDgic5kBDAzMn+HBW/4gwThIUVF+FFm0+9ylg32KEff0O70KNz0
O4oJaBME/NoH/oNpfexrQTRidiB8C6pWu6aKINbmpB3QS49kDCe9U6adp8ZAbdmVQ7cx9794Enkf
YeijMX/m7g2DocRxARSyUSS8Re5fAWDCtlYwxSiDh2GzjKaaFeWwL+tGXmWA36iKgJvXK9A2F+E3
hllr0RaneNl9o1Fylomgb+x2+98/XQre8nqgiH+nTf5HwVF3m+tFfQeWBndvw/oAVPB6JL2uAPVv
RUYDvUjrhibgGrhNtM0WuRzUJdVNKWM1+HK4K7oiQWwMihSnp1/PxVbIG3wyWv/oyHGmN7P3Osqm
84UDpW3s3xfNRgP6NXMpFqaRWdOAXTnzNwOgWzTuMYpJopF0ykgMvZ2GHCkcJeas16WxHxzhL36W
bd3cxLRJmNKb41S2dyquf5RPgPPXSEyLTp2HzOeqo2yVH5KANyys+EnDgoDoOivHCP2FGCY5T7/X
I9Bl5T2C3nF3QeOFzI5DLdCMFvY8U6xpb1X1zBItf7Ub85smEkzO6farJtE0LYlKWoGJr8mEjZn/
Tz2tuq8YtuXhznCrM+d92mnHvNo2piqPkMOCU0BfEeOJ5ICpbccigCbFO0HQ6Q6tQH3vbEmJ6WrM
igL9HvDFg6Ye3i0xs1r3lr1HNFSQg1uXEPpj1PqryJb8egahPYiz5ABhJ/rNIvaRkMx2ZU8dNaet
QaJnAm08qOmDOTZpbgHxrCNxBywwGJSZiLhyOxCq1ideMvc3sRbiMA6oCV8HDJy+YlPrOg59FLdY
3HFuQ0drlWjEzuiCVTgNaQmVd1buokQHAeoO12w3Ttu4GTlNjr1C2p4Es6w7C3H4PbakHyp9m9jo
gRHmVb/ykMyR4pm3YqMxKUgSPVgjle7DuJMCrZ1fDPrvxwLniBN6UTaXX3SCFuqPArIfQvhVSyj1
4Yj/A9Ohw5qfxl5ZKGHEV/t/iLDqZAkNUjBWjNMuZNz21v9irsq/DxW3FmHDOuLX81X9DciRS0t0
iNv8+fRWMVDQvjP4EljhSotsDxIQnlLmEFZ96/Rnyc0J1sYNEnR+ASS1Lbo/CQyfdHvipKD8ZO6T
KRwMMP4DQ6UJvFxeNLVjQEEQYBQ+f2keorUiTu8DoCJRRLkQMurj2FfSOOrdu8lAGVnNT9T9ex2v
zP66v9vTk9kgsHUrjcJ7bRcX/mo9gy/xvJTDq+0ixzglLW/VVVZE3PIev2GOSgn7DNXI918ODpCP
qy9eK1K/EQG7c/VKSijPj1IpmYWDd2ar60JezKpmtT/XVJTVLDzwSqNV9kXLTF+xWsGiFiQHu6+h
kvHP6Ht31XfV6z2GClKnWTHweRmL4ylSaNYQz3jaiaad8eFNyQsREPsxBpn1cUnTrvJKnnlUTTzt
wfKj7DVLipZtg5REFrHHjZwYT7kh/s9JBqVFwiJcMz23nax1jhq90DDQ7AUqpviJOnhtOGVfxGhN
KoMEB2PTgZB0QzFsnBrEyUHUmznL4/SjZ3XKvAslJg7ABW4VbrQjrCvai4qFFfGtqcSCHDLUjrHE
oU/ix4ltVI+EO5ay//ZOIGl9puv/T2oJ/QQPkfSxohPPWKRtcsAirQfoDzB+NvIM/al+bgJOG6Ae
BtIDhD9nsHJhZz88OmhPtxgtofv2ygRHLpl12Xsw0R+ldX17NusQy3oA7S96R5Yt2nE6jjnCzzlc
SmOORDFWOIMms+tHiNkIuiK+4At16KYf8dzSqulzMP4oybP0MQFCtiTVFJtB40MOQT9fUR3NcQW9
12XU0Nf5yJqdroNdiNFdoyJCLzUQvoe3W1AoSeos6nNR27ii4Nz0auZtq9lPZtqmJyH4uTThvy+u
ygR59a/N+V9OpvhZ5qVNnGjn03DCwrWfOJ5559cPE3EIfeyH3vxn0QDIvATYtKLGXiBVZWo3nPu8
o/hTMk4ShNMH2v78hLXjhBAwDVLqagMW+tFyhPie5tAq5OyITWyjq0t67S8hNZJm0WvSjcbu/wUT
R9j9cA8kjF8i3U2XJZJk9b2cd1tp2ZFqCysKrEG4bde8LRvVuk7miOcN0fsrPj2nOxdLrvPFrq7g
/FkwZ2FlDd3RsmuBXS21aMuxBfwALvMvE0LCe9eN3aFFrBJTmCufGXqXXZPUNxuErymmX0wwpdqK
4iJvDSVomr4DcQyCazezhA0v3Krzf5jAybcFzHSNvs8YXkij1MTJVoI4It0OlcWWqEu1PmpS/DO5
3xCBCSRt1nbBHKWVCrpLyHbtvWM/UNU7ng6aPkWpNSHv1+IULB2hcO5Z2m3AnSUQwBAlpEP37GQM
Uq5B7HLfK1SWj3FCzp9Q9Fh0j5awRP9I4W9slsgmU2JyG7Ysw/ieO07W6XO1F5mMqKrdHj64dvbN
BXx7hJSFqvDOCBqczVOKB5wZMGKNUXkYtsUe7FSwUZfjS/18GwMppdbgLAEF2ssn7q618VLgz91j
2/5DJZglpVQNZIIGNHcA3cYnvkwyJI0bEJPA+0PSBI0SjfsgUPJHQV2w/uALbuwlZrg47vuWldVp
fQG7tVRqxP4eXJnSwUuGO3y9NCmEbw7MQxH4R9gSjFKnK+TgK6ITkTe3IW5aSXDvc8ADEfR/Kgtt
AhLb14huHzcPAo+Sd+bj/25O0epiXxrlHb3dAC9qr7ITe1w1hvJC+nuQs9ebn4FxJxT/ZRCivbox
KanFR8Y5MOMayhoDg37ThweLPw56HpeRr8L5ckcSrLYo7OHNe3l5XNfLW+MiUzgpE+x9oZd1dJ0x
ZPtlLyo1wqxzpM0bYsCWxOo41gjfl1xsJQKNj8AfseGyqmOT5Qxg5bYI7s1FEaVToKs3jUsHc954
YOUbDddpVcc8vae7jcE6YKzQRDafcNcM4HOcwSu5kCl6kh4h8WpHNokeCOCZYlZz62dm94IQPR5M
VTKdfElDlJ/1vBmoTkqr8VjYDunucUQajGiTxjH1vDINZeCFqc4kymPmaLWMGEZTVE0XLgES+bVp
HHmzcxkcumZn+vMlAVrXa+NQfStx/MKLkwg6WuQfNg4oOKSdlbYleTiIzl4/FQtc1bVEh0fWu2bS
jvrN10T1jFKbyLoxbpToyLTMewjtZXb1l66kcoXu+ZPQgJGdEnUTilyu4uNr1KT0YpiPYT7Xf3fJ
jgtrIKKDeb88B/xG4FiZC1ScDuqj/KWoVICUG17WDXMi1fr7biMe8bRyZ1KJ8ElIlFmoznI71Von
rGez8s0OgyM+doolzNRMoVtX2sEtBxC7XOZjyXJC5s9fDcEHLy0cYSqBF4LOBskb0JUL8Dm/239B
7izlpU1WGiRhcdoDpiSGcHwAnjtHzNv9URQoEsvAhzOePVJncK2jRCNrTXcl9gda0SNCv4CYf2XY
FmLe/rQdzd/Vgc4xiOudKX2YPgkbn/VmSP7fhvCzPEJmOpOaxJj3OFre9yvwPwRaDln3tQcAJHrX
4YmyGCELbyV31kgcuu6axAeiMlrW1iUMy5RHRCP6aNdb8tR8pYKUWAHFwj6fPg519ZIjJ2+9sEMA
8f6iNOmI3l85LSXLLgNwL1l7xegUbaGLyj2bjBLGdDXDkjASSjkzUGy7hI5cIiHyVeuJLbEiguFx
GsO7wbawaNmOI20dttHfGmeY9iBzj7hualwXok58LI7aulrye3CuD6Y0NNQ91mbjgbtxxj0FH2iu
tYCPXUUi/bRU+K1tGJTlGeZ0DqgHTkRqaDwxZbjTBXhYbTL9FDsldIXJKqhRWma6lXt+f3YxDAeA
dA2+LZxrEH1gFvTnsTtiEI28J/grL6b+RagsZhRkZ5CuprWVxqrPs7F59OjIkgsGJmP8L1bXaD7j
nyxE6K8GuekZvIsGZNLR5LUIw09ndVhaQn5YdvivoNqnRBehFvxpiIIka8vwBoASJyuxv3EkzxsI
o20L9rpM0XOpK8pUqWVoVayfy+yArmGQlhwv4/ozLQhSLuGSlNcZ1jt+GCAN09pFcv9rRkdPDyAT
qYyCFrZlcrUTwqJOv6gYIf5oXSLYfwgInJpkDIxtqmv6ffeUY3Osr4K2aZmP6THv23ONIW3ZWqEh
NxgVgxPu8zwlAWXA5w2c9CIKGOsspjZyUpm4L19rxqCv/tv4In0ZQmaSv9NyPVjt582DNOR1aXy3
y6V45S6gWHcyohaOlmSHuVavQ5odUpriBD1eXmqWYa0dCzNZRWzlZu3vOnnabzpMTiUnzUn7Df4k
4NTJRFr6Ye+6hwcRFxfm+9Wt9ZtxbV26ppH9US2/t6bW/phXxOR0e5zWqYcNPYKcNrVrX3p3bsaR
7sqlb10Q9OfjF7K+PiNi5Mf6eOqkRDzw+D4hUixRXDuj3tAfGAo3e3Q7+bAJX0pTI5QIWTZnBw8L
E1u/7L05gHiwjdmTmXTl/tDyZb+RYWtzcOUrketxDKcTBytK2xLb4P1A9EwkyZ/N3aUQNF+qp/qW
hEIemn5SDEVnNBSCWgt27RupQGQU7N7W4Ib5zy4wf3wXE7sr3J+UWvjCFxuFoPahrTeg1pHvyQWj
4LbcUOtKl7neeU+gXoYzq1TLIk0FbF7Xn7lRauiOFDFKXRaIAOrvVcKelcDnnFH+hG9LpIZT6eWs
Vje+Fr9PjDMPyb19F4EV454YApGOZ13STH27yoV6G4GPxquL+F893AhpW9fYU3TMAiNSiha+BY5J
N1ihD+i/RjuZ8k/KMFH/0aD8HGNjOVLaMfZfJzX4ruPywlKkVQ34aVtcoE1GONBrE3Nkdbscrwa0
c7OW9WLLMlxHiTy1cCj2aehIzN5Z12xAn09iEZfTM/BOWubBqyc2Wjg0cfxDEKbB9f5/Xjy57Ve/
vNLB6dGCx/hojdmbboMLzuh54hdlkFZCyGHk66gTYsHlAjIHGNapo49fFBv3W1olRFukOgqcd66s
z5Eu0xJ1kGBVD3UR08m28LDXRFEAA7mIoBLUSyawVCykYi09GuUBRdziY0LUbJgIpWFvfcPTjENZ
pg6NCoRg1BYoUO2az+0XVtQxz8wA5EDc+yOM0E+nqcS6gH12x9PrjOzFdFkK5n6iGw97Ko8ecoki
2ASR3l52O2cUxY5PGASHL5BruppXnZDltMHdNgztMARcyJ+FYW9WeUYwWihLkadGDttpBvOT6nzZ
lQVOibImLacxWSmrF+K8BALxIEIrZQs8FVC4xTpaACwuonQKZQBvx7GDT33NKHipjMTNcyuciKlb
Pa9HtqwZ3U99H6AiZAe6R7a9WDF78n77BliMe0Ayx+fxLDkNypMUzK5hMABw4gce/gxHGM2MsR6e
Iq75WT2wK6l3nIcifpc9O5Ak51MNF/IXfvjht0Dk2aVHYhgc4c+R/XMGb9dwfXii9vC62wtle4ds
8ZTAdvktMnnBCHSFw3+p3O10WBfyxBPSfHaM2HPA3bvTv/SFrMyzel08oVwp+79t6Rkys64JDUk7
+nRNlv7TyRlT0uaNcKVfjwioK91vLZJshGYgRcO1Jjdd4SAemQqvqhjm2yDhVVVeGLxudujnUYU9
6tOC1RIPRh7UoQ05o25kOkKXVQI4e4X8n1nq1kprxC7iqg0t7SeMQpQDy4MLGpTqrm8mIRcuRENt
VFSVRni/PseYzC+zuejNzCAa3AJfYHaoBNwasmbXes6DbK50bGyuk3Hg4HPkQZbEM+A8sRof4cjN
1uqdNlG+Y4SdpNRIxZJZF/r0CHjutJq60Yu31bHDbcuMBZ1NvX+Ryj598SuYVbcLRqpL+08/z/8W
Kk1su3azzTz557iPtdg80/tFfV2uthv9CnPJFyp3fdVPjRq5k5siEBEcPbqMiCjhmgfyBNlkh5uk
KLlsU1mZegiSSRgbALC4rCsckw+xxwOl/RDPrcJP4WFLOxBP7Hp33zrbdslA5qVcYi+umGBc2sKy
yUUGSWk3exZ/c5AqKilQnAFdlaCRKR77qd+tSezjldc55RvpgKMqieu6WL1KJxqFjxU1bYAdKPUO
eeABUSiEzbiYRRIDtSDc1YOMy8aokKLzqJxN2SI3jyhGi3feK4tb2xWw5ZyFdFHWo7uT5bTP8zFj
AviPd+Edc5F230g1sXNyFHe9mlXYqiI9iyjAdPN59yc56BcqL9ItkLwi7nIkKh2Tw7lEisSpRdxl
5j0dRGwuU8kERBuh0bS41eZStoNpoL1GgxsKl8p5cERwp7Y5BJluQkkMIbcddIgYkGLJOmz9juN5
5Wi1KzLGlsxEB/HbISNQvtbY2625n/OdT1yeZmKM8hORCelZRuA5q3II0g37t8kZ3W0BkFNqHffn
ducA/xfIhYzacpovtr8om+rjbXh33QtWlsrsSGxd/1fUJr5S9HEX2XoGCf4Xygaf1cRdw6li8HOq
WBs5Oix0rZiJvWdOMxmriW0G+Pz5Shmg09KWLduzBKuWQXH8eI0MwNYWb0krsTN6eA4Q0KGozGdM
Bdq17rOITNFCliJezfOlfAmBwlDRdVb+zlV/ONw9+UW3AaeKwG80q4vXTf2SIKGWay9f+WMKATjI
/q/sH76KDIz8RWjYdncPLcBO3ei/iG5Ke6IdRxuhIPIUFs7laG0RvpLGBrTtLYnKHH2TT+Mc8nVK
6VYwm7cRWcitIStanPpVa/wyWmN2nDjX4s2tAo9RXMvROh9fyMND2meShJiXGiFV/2ZzOwn2CFYn
xGQ2Tjg8tSJoE2OsHDHl0MkX4SYIKa3XktMJ4UgxAONh3AbvZ2ofnZAXwdhbmvS0B4t+mgFcdU1N
3j3uB3oFPQma/rinHLd5kufaIs8GYm1rwUFfaMlMfHRxR4XdrdjeZB18WlFkHZjve/vKML8tbCDd
KY8JEy3SBEmjIiueQTZxs83LIe9oaQPIOUoUwDcprfJmo2r7rMLtnvgs56bMQ6n8kzoTKH7LBUWl
bzSHhoZEpVZEDky/90N6oveRTeZ0QlD9fXziyNUCnk2m+Rx1eOZJs+sdYzQQdVpINCWLUrHNWMZm
2DWn85SGUcWdogmyPGePnKY3fU0JW3EPC1rOKfWvaQ78HS656smkpq7Eoh4kxmM3XASuBm9ToDkQ
wXxWe+nx64lPx7YQcejgrP+jAm1Xl/K3/oo4sgwvBwurUf+CW73vgzhEQXPVquGqBuPGjqfjHgWI
tpTbnJ86DZ/0LJf6wO7czX4DDZGFfLJK3ri7gndjDhNZlMX6TPFOztXJAkzBJLfUikjnVV5QGkW1
ApuxPvqXy+IElKznTi4Qqds4jcuhsaG3hQsMzBt9TV0Pq/f70L9kP7ajNory2BBn/HEeTxcLgMVD
flaiIFG/MIrtOjV4vfFl6oqQxFfK+V3txy6VOap+K0ukP1wBq2SykX71N6NzPYCN5ycdNWhjin4X
2QoR2RK6pUDpvDnuSyrDJqKDHHO5mcPTYyL4xHtYXirN1wnyv1LsZKBFBnQVZmAt+Rmx9k6QEcLX
DOYXvzo+xWn9sE/9L5iUpwB6mnIbQe27EpZ+WMSLMbUaAleiSIxI9TRx0QRIjsZpveFh6uozR30Q
RuIKrEsS62eud1LuBKpIErnl4bPO8IOKKyhQOrr5qsI2OHXkSUAUuWjDHV1Hn0jtR0fNjRyhXGVX
+SJPWhRRi7jf4gY+F+GgDJN/JLtHT8S9l7dFmm/17ZiHjw/KmyNL92JsI3Il4uvlwZS+kmL+WW8k
Gnd3KCK/qp5DVq4zpe2MyQDT0Adjc4wDp2B5pLbmKKmzWl1AMiLZ3Bo/U0kUlpbl7ra9Fp9mPaCp
TRBHMZut6TnD3xVZakAOF35KlO4ZGlsnwgWXme4kFbouN/cMn61wQlNOoVbsupvlQvEV6aXd/X//
yzqYXptzUAxuxRbhAcMyvlsvVh4SuhpKExw2iJNAHbMN/C67eRIldKGHJjqJ5QMbN0qQcR2dKhH2
L/nx7K49Vipbr3ITeVxrI2NR9rgunieBfELDih+Tnp34Du8qwwh3lgmEWHpGr9CA5nw7/cVWbFBz
oaBa6Nny8JMeu8au9v5l9vTvZ2ST0p6CtrrvNLIZi5HLGltVlvYrxVTiv2+h9dUTmpb1Rc9duk3n
J9dcGMsNfF01Ad3p+tT2RTJ0QZT62nidorntQjrgl3S5uCEkHjlixG1gaCZE6FpyhPO/MlOxE7ok
H7Slo8lnqO5t2c2JVQ3Vvomv3Djx0eAnqk0vcnxszH7B1GRQbSBs66UrxqJ/J7Fs8U7r9XviqiS1
73UypFJ+c2CGHDqbDdkJPsByFojOT3lM3G7e3Pg6bilItJ29P58VKsBbI4zpJMnzgqq+iAAGSPGV
Yr0Rg0RFoAjl28o+km+CrnTAABaeu347nVeqVIK3dCDYDEI3abGawbG6QFG7YzOjqxM6MuYetfM8
aEWsMpOfUtfl2LR0sWQkbBPWyb5lygseiT+ZLJweVCMEC9leaXDOhz3Jrv7wMQhAfQpvAJc3mD2i
kGoXASV7rFWP0NptEY3btD01qcqGBwy9SJlOUwuJiIgExN66SHWjMVRkNq7bso7woCesC79SWz2p
1PjBKWrTDkzkc0ozVG59BX1WVjoagBEF/VAnzV0niu9znsRb02IfnwL5AI45+yNXTgkeEGljwm65
v2JE7Py8UNPlfT6zpRnCFiIn76dSHVEz7Hm86v/aTvRTT1FaF3RWnDpnq2jKrmEed6JK9gzah1u2
tTgxduyQmcFCSlP4SpRBp7ZR61uxh9dgzu/rqzo04IsSBg7Jfdr94UD66I0CcGBL3GRYld97Rq6w
zSIglGfhLscDZcvmACYnM/c3XE+0gKldq2n5zta2ikHN2MuqY2Mjt6N5+PCm2k/lFSfZpetvfFGY
Yz4JPyNQKbLIGWvSK2G5OUBm3ASJET1O0TT1h07gFYblYJdPGEfFoYEDzTTcNElXyVFv1x5bv4rZ
Jqkis/sLoZr/cEh0kLq0yt7oL5YcReeFUrukcNISoVF5tDCFuBAJ3HwS1CSSon30ig8ffgnrqG2h
lH0jYdurg7GYHVeUX/ocMyVH221z4iuc+mqRhbrvWf3c7kf8rKRHFDl59O+SBhdkuomtqQ6VQh63
HWLBn6uEZjSFuCYJ7tGfUNwiPbxChIZMmQeo7sAPMAGnTj1czA6+8UkwUU70wGVhqe9uEp+bLar1
o9mg9ONXFPsIv1a1C4N1ANDmI71DbGSOO39SRITAmLJiVlfkn7JHRjkOs3kkKp1FqqWgNcRVcEoc
+iYj1KVH9Y5S0n5mFbNCAAP713BzqxJbuSGVeXJkhxwywDwiO/2MzKOAMHXaZCPoyLWkokGcUugq
AkKt0PC3o6FRViBGX0xHAK2JDUqqUqMOLTGZ1KR2dpqoEl8syoiF+Mhliu4lyKchgMtsP0aRUhdm
pmk1KJM9paFTx/3wM+QRbDn3AQuTSQSTYXcJEnjf/21QoBfAy7IgYmVkwDFFGBjIlHz2GT2udFOr
YBHzxiPQSrhHKbeZJl2T19rPomDBHa+aB39yxbHA68BOS1ZmrXgnb0qvMVceyYpa9G9lPqVmM6Kz
618LHz4dL/AeXOWxU8yRlO+p6iM8MbA+mgeF1mm1iN74hMArkbEZa48LxWX02YgwDCDsbfAQeJ3N
OWWhUvof+zWWGV5rVLou2w+xNFeaOkRyhXJmHHghLpJDKZXlsGloTSJjjy2+9FnKUXngNH4zahJe
rBcbhEYNi9G3aVq/1uiQzYC7Lb9fajEFgbzD2V9QAll5ErPsGhs+MLL+5ExJEah+z/2bu5UV6bd5
WWBiiP1WqkbBBSFkosAblQBYMqpiRzBs4/HdD5uIHNCNZSRrHd/d5JRcSYZfW6h3gai34wnbd3nD
pa+NdjMrarJkYxAhpGZedg6/viIYUAAUNwuA7YlGQ7DTmhmE5H005WjeRFFVEFKsoyeRxOAyqMmT
V62xlbnC7id7I/pUgOIt1YAZF6PyuMzjD7A+9Jm2gRQiMJu65iTaQb3sRP3rFrbejUzp0iE4N56v
4r/0m6AMZ7Pz/523J6/9mZYIfGSWGBsYyGEA3bUyJGvhopOx5NcZ6SYWvod66U70xx12qqVfVBHN
aOpJ33LKH5gF2l5i7vNgfQ4OCrOvC304mVvz24Z9YdhQLs0Pmchd0bVnoChcMjpMpsRqgrl/4FeC
wHwHiGbBADrFMEJzIGmIrszE6KlZx1dcUetNVJH1WngNrR267asyEpMdy8YT+SJK01CvdqlUUVrS
gcKWDSpFl99EGjj6/rRLEFDGhqufsEE3mLS6XL2iUAsz6P+ZDc0o+k2VNfj78L9F1jxpbqJILyqg
ZynaR5etEYt4ugNu2qTURxkJSY1HusJv0P+Cw0bWR+1pQsUc4dRcvYD12SIRT5GfokcjPT552l3g
d9XAON0jkpFfH7q8AM8eh13uMHkGIFRISIqtDKPM1c9MNuYU4ECYdfBQZdvE3p3ri+2oM9hbJ2HU
8hATrxPul7kdg5A8R1g6FDGpqZqPSbSmjgn2wY0DjCqPUmRgb/34zPf9Revt3nZuJBZt3DOo0pjV
Fs63hsOD16RzTzodkChM0jTjhnkkv4T28i481Eq9Bb0D3cle8UNGF1/dZh/uAEwY+9okoFkiAPOt
6rboONgu/dK8n1tx1MCG4NsnfonC+S51OfbOTUlup6acG5TRATnFr/NppoBsnqjGxSN1mu5XZsuf
mJvrOuOLRynqNTOf/LqCutkEAK4uXaPdtjDNqnqJ1Xe1ivjTOxW7P5ieXpEIIsmq933fRuPhZiqR
7KJPMY5kiBrM+291itL5SBngfy+oZLCT4uI84A8ZMyV/fDffOsXiXnAJ2xwAlud2Egdn5oW6nue1
Zhle6f+cT4SC4r8XfpQMdH+lm/DdplonokyHXYcJqCNiEuH23WY6wg84zFhLHxB7POw1Lb9YqyGn
bFyYtKpLIQpxYHT65BGpPAlbz+MUMjR64TK+jH/VE9CUGwWif/miMpvx0kWzAoyeI7SrUsk/bXib
9USZQ0wOD5oxtr7Ts71VHtPmM7qZjcMoqz1hUJdErxZi6jiiAD5pjSU0dvjnQqkEyAYO/YkKe7q6
G22RKQLlbA+i7bpIeRSymJno437xWkrT93hLhpNK0rqplHewQ3zei3a53GoY4unbz7Rd9TQVSNLg
bu9CDcrHWAws8OkiF+o7bmtz/8cGY0ykVt1To+wQ0kYpB7JyGmFhP0ZyYIeQC62yWBDMX4IyX6Ow
LhWek5h+3pnNyPcbA0Rt1s/NyTq2wQSfs0dARFqUetN7SBiNTmUEPAfOYisMeJ7RTMujM6P0V3WY
V47I3c48tx/R5XxKHjUsea/+YeSUpFtcduD0Oqufv+gQQZfJKs6NvPo2imUilrlE9ojjMgI1pAwZ
kH8m3smfedBuxfECJUosGF3kG1bz7pLpzFeYhkXpbYGHTNqxT5FJVvby+AZh526YuVfIvvQcaC8j
tLd8IdUVgUU7fqJYw/NGp4n73vJMkisUGFV55Z4Wq/s4FiX12CHvzU9ArUk6jprWHdGUD3id5xlP
CdcymTOIsiXz2T76ilsS2sYyIkKFtqMxXuCKg/ZEF7XustxFzPQSbqXDp9YjIDv2MtkxlLAN9ar5
fSvTPSXwc0H0Oq4e/t643x9KbKKIlZ2ylLEmV18+ZBm6sFnVDzvXr1IK5agt1NXfjCN1gxvPdumd
sf+HSMDdKixtBx7ac6h+lk94qrcyDV261l7rRF4JI1Oo4IlAokPgdPDggBXtOlwli5B0FBQmd+wl
MOt7QtsBiL+rtAQ87V+Gk8bjlhK8+YHDTzrk/0qO1IZBRH+slqvki+SdVWOZk/wGaJibbL9DbQ5E
aNelHaFwsFHMWAZdP+AifwE/nD2VhC5xnVtiIBKckHzmg4tNMkxQsvgzDprjGXo+M7BqTjijcHne
zZj+qoFdtlsrze1qiHpXCHZMPbErbVwpbT3GwN8r0xnxFp+sn8kGSCao/h+b4700/UDcZnKx25Wg
NyW2qOlOczAKCMz0muxXxoh79ILMG7zeIdAmrBX5bwtcShvN+xEiSqZRZ9C+SGd9mgKL2isPAUw+
XNRLC9pN3TgwGuN4/gmk48m+/N7GUaLUKV/I5I0GrOaalgIV/7ttN4oLBgSMtd20gs+43Ox4SH+Z
EDbdkWsBAuU024mfPeSx0vcuxLlIptSennfym7r0kD7qDP6J+kWsLGHTg3e5m8vlfSYFwHkgGTrl
LHtM+iBUx3rp3bTCHLY0eMDjffLGarj5VbG2FiL0BdUvJVopj6FzlTTTybJc0L+2oxNQwM97k2jr
hI2cJLgj0oz3hDTwCY8Hi6XOwIM5aYLXAGM8LDZtgNp913T/dYUpH++AVI+QP0JjV698iM+rqy1H
74Dxz7SIkZ1rMeTDahUBbdFliPifdQqFOG4eReAsImSybkE4ObXeYLquHlcwEiYurU3+lDAqpwQK
SYhqbVwWi8B8XHkorLXeVKpDP7zawgMJcc0JH51ADCnmpxbL4yvgLUNeGajg9wxnJ/yNIOj25J41
sDpWUszLzDwLXCECq7/4YA/oKqRCpMLze7+7uQHLWK+6+U+niaLC4HjRVNJ20d2iNLPRKh+xcDIl
GeknTOaz5ohgjShenwcFw5H2eSAkYl8qWPznd1BbB7ISPGpbWZmHqGwT8jhpgX70YC9g5WkLhXsn
WKcEk9fWUhlfovmVFT8Q9Poa9A8zeopwvM3XeMPp8/xmYPm10rILGqxW02A6srgpC2o4V/hQR39t
2snKvRM4qXrlqkFfWvLjlpSl8A/JwiLr9PJ5FilAktBn7bvFWt/jye/SPFXLovX1lgR+kQE//PU4
WPvLCBFAj3qK/F8k4hJLt797DIHtfEPpv1cv/E6/9ooXoCydF0Az+HIqJR/C1FkPZOp7VBSwVaUQ
Mp+VGklvg0HqKAJ/LJ+6B8uosKoaxCY2j4sZ/QDyxKPkuU0wQwtmyxnKNmKHzrFLC+lHQ4MwCH+Q
G+r0GscFJ+kfL+UjMGxD8ccNWDNVmNMHJFkjAoY0O+nW76pIi6aXBMf0b51JyI0KDxGz82Z+Oh+i
RlT6Se6yqBZLfJ3Np9dB2G5pxpAKK8deQJOlJsEb1Khtydj9zhL/4vFmmZdTbKCJBvAhSRVmcrxW
qmZOz/yLuSKaFWGyhq9riqDLlphYTD+RhX5kpmud8aEP+WgxhdS5vHqtB7Dit64uv6qE59NaqeKY
ZExhUXfpoIBVpjiuR4IY3QVYozipjeH9Mxv7AXpuwqlao9Rwn17ZaP6Fuz4wIdMwxFQO3bLLOGgo
QIOVuFHNwGXuAipGgXToZRROH2OSp/vawPsKh/XMYd07OOFDNgHyx3VP+6sfTQxSY/E+0D0EtEO3
1ExmBSn9Rj9HfwP0AnqCNKLNbaysfZ+PsiZjaqmJ/7zz1KwZsIQevfHfOwkPqb0pf9SQvd+UCmQf
GFxC6MRSv5gRmEWqC3HLfnj8XqWsrtCVd9awjUiXhNn2hoAJk7W5wjZv8q1GbqvNeRQzMqzBgslQ
RpY0Z3MC0raPvul+h92b8UHY6YLlv+0J7Om8V/AO3+eTLWPcKdAPDDIEJTs9z19QBhVF7jSLxuA2
PQ2CR+2D0J6Zni4ce8kcdHwZ5l4OZXCLqghGj3GIVJXc/oXfF3B2gudTVoSpde+Hm9ZxuvguASgN
qJqCiVJJwPFNjfYr01WqAOI3BhVydYhiC9elwgtF5u+PE367+OSHE4v9P+7Ood7yBi5q6jrQKXVm
SSLTovQ2ufNw6CZ13J55pMqu0/i2GZO8roDU73SdkU2q4o1v1c6/5yJzcrd00SOMvurFwDQRcP2a
gMn8XefNYo+gjoFielnSh63lZ+7gBI+zLrtR6279RtdBA5kA/OUSQSA3a03eh320mYChHDNIt4Y2
f4Zn+c1oD8zhNMDC/ybOb9mZa4FYJCtGADVTU2109pcATFm1nocN4GVJTLycqAXB0x2TAs1Hdi1w
zqKLV7AqJCOibgjSq3L0YVvFPRWIvSwAFgp13GisZHeiz+499Q5pRUgBIk0CYayM+F6KTHbD/tBI
Rd52dicR4c46Usufj1ivebj23SBkkBSCoWAsZ/RdnyGdxQFSKTfp4sN8RZuCtnlLFu6de6alEhN5
kuwq1wQXdEIAJfiT1Jd59bxS+EdJxVTQfkmXmGb/YO75Gt3uHN4O5Cm95yAHuFywm1bFuozlil/7
YoHp9sNExLVoKyEj9MkvaO6Wtpwzci7k6qWyfZ62v+dowemMNo/L61qlfNm/9WM5QP7UCnzDYCrw
r1TU7p+SREeyaxTJB4nqCbANe0sfwADqpL8QmlRGIicx9sB4OPRu5iNxdkK3kNEDXMwvxXgDdIkq
9MhX05u1LHjyVe9MQ/Nwe2VD72DHT1+LKllATGI/r6Z1y7BSRXfrZlvP9lWV6crUyhCQ50ykjQwU
ZN1RvUHfq5pSehjyO6RDsGWyqomfOnb8UDnAySKD2uJy7CQNxM6CmjsZyBb1JxZTeZHBjeBy++SD
5rjOd0FTz9aB5GOyreYuZsdBFDaxkbLIe6xnWpFt1uvi7fqgLD7AWWYClZZgPaHAPuSptSncEjGt
/7U/vIfikSQXPy1fj07eaDUFCuuKGbu0KFs3lHLLNPAm/bopXE1rSF0+hIcAhEE7tLetc2C7UB/A
T8WMxuNVA+i+Uu8aBJ3a+rjahrWtKscSnUFuTDiUUlC0lN8P/WgQ6HcVxfn8rDtX49V6YxFldF91
v2/XuJl1gziPwvVVGwP/4r+wEUpM9hOYgJqaRELzK2a5gwmpl/aFU57L/83LqKDss1Tf7UnoyQ3v
eui3PQyRfSDK6GludijqmKG6n6XJ32ZraHYN5ysowCEOvck+RyrZ0fbYxi2HluLJrOAcBYGhVRRq
0vX2gHwUydCzCLhj3hLrKy9eHYlpqxZiDMwPNhN9xAp9N9KIkfyGYp+I2eVDE+zP9sduFht+IfEE
R8q+XxxqfiCa1hxlJ1g9aDYEtUiZmODwC7IOiW621SoF4rz7dWTkHC8trhaMU30HQm9fS1CL2hSj
0P0vgzn+yGrWa+oVaDp8x9i+X8CkYnsXVz88z7kpe4EkqFuyDKrpg1jHGFX4E3uGEamHG7+3/aFV
vqh6EVQp43bRo5zJvklx1oYUvETG6PQhn2EBRE8MudP4DJb+sH7Bv0qAmY7zSj4+6uTJd7PmFKKx
+Pq57msfV+GkEONtZlWHSPhjt04+5pYQJc/t3bGyAT8zE1vyU2yXo3mXWYJEym8E4yQpsKGJlG2R
9imIycxfekSJdRXBlNP3CoJZ2C+HzaPvfr87dsVWlDerFn3gs9v79bwMnZB3FejU81a+Yn8y9Sj6
LPy5Fpu0+AHnfkvURlUu0nx6XrtLYWCRAZVwCSQrNuNgCOD4zsth+eZzV4WoJnDD/6dMJ7vd6C4Z
ktgRvkTOLPYX19THSpvmFX6NFUkLS7zYPish35tfvAMCQziNF1fSiptBsIm4qAKCabTPlCjYU0Dq
63PQLnodetHwyG/pubVyk5NI892foHqKOjXX0y98Kz7Iu/XmULRjq0e2Z1/ElYI3yC0O2arLEhHS
JIHa7a+lHKoF1F56vrBhKPCCra8VCuqfRGIbHNbaEh+gd1Kn2wi08SF69o2TmTMN/xtn0mvDLnJ2
UYZ/BobIgVruFWxJdOJqQjOw8Q0GWdSYYhZ4ZE4xVbVTeGNPVK9+LhGLFKaDLOpYvSuX+hd9+/HW
x/jtt3XrczvJSwCvjIBGlN5LjB3IhZNQM04kZtNIS6ZloBlQ5k0BN0cxEi/Fv8/M5I8PsrXBxrL5
zLkG1psyHRSUve81LKciqeKtFCXGst2gRWtaDwAy5zT2FW6Pp+gsSkMDelXVgk3hxiP6Jb2fqu9N
IuDggzB2aEshBs6pYI8HDzfZdwv/r3gPz4IWVx5fvQrSOcmET4WM4RfUIMJASH1lSSjgdL1q8fe6
DKpltH8lrwdxYBzoXpTAktTc3LSHYY8zf97cg274uvJfqnCRBaizWkGs98JosUy4UCvbe0lsysvB
Dmi5PwYjG+o/Ux891KFUEJxorih7qmTJO37vtIfKlkXICqzS047m6BFrpNxk0B19Esv0XGpGj4gC
QEZrRebRJNbVu0Z7uqhrlpFaRY0bZ+ZM30j8jGUQw6nWVFnB6ZbRg7veFi4LitpQTFHttUxWDys9
EBhUplk7Ko0E7nGTum6iholKhBUiBJFzgez5gePvCqEYcjVgNeDntbJx1Jj/LDGS01hswLhqb/yz
HQGlfvt4LNWfS87xzgD+A/Vgatvj/LdMfYLjksRZ6ZGdRJHzzka6aYadVkemjX+IM/lCzWF/bce2
0/DmCKHj6LvsXgggG6OScY03levhv0JE7brShce8srgKCNHeADod9DqWl2FuIdE3KB+/l9a90Dkz
ZJIbGWM5wuyN7kmxsCsJbOepJG5+sxHGtPwn3ZEWKer6Q6BfDEVtFgNRWxyUTnWukpaG9Ifn6s+E
h88dqVeLX12M4s6iuXnHS77ZEBE009qbLQpzMPm8kS2D0jJ2hMLgnFdQbH2w049Ad2q5LQiYBWrj
3KsVHLDnD8JcFeW5OvmD6R/fZK87aPEnGlvGnzZRGcjaPDXHLoBkK8RyJqYWwoywnvhk8KNA9gm7
iyv/UzPBkXlNfqgh2JZQ1lNacFMRPAtwJHxDMCeNxQEWB7w/p7s10S92Af+LxqHx85ft7rxzqKgz
P90/ZDoT76aHZ1smH+MTtUVjw1YyuowP+hjBt856E8w1YtiHQrilIT3S/bIHeb/1Ob4yxbjy1MeY
l0iLkIZpAAnkHRhSZ3pAMLV45aPn6SgigqusUnVPf1+4q8e9jga4JX9qbnJI5RLI7adSaIgCNTPm
bToGDtT8WBx+aBJYrfWKL2mXbUpzk5DPf1SbaVIW4GPNME3CxmTRHk9jDKqaA4/Z2CGcsem0FbLH
rvX8ryc9updnCP/4h4R6bV8tMlVF9QqK3ud5NXvr0T9Qc5wwol+mcu/JokQwZ1laMQEv7ry3Fla2
vrRoAgd6AeXtzDWxMwuWjV8ZcSYk83KMzCTz+7CYVs5GJjoM9R8KYJRGZ3RPvJ0Trf2vrMbJA0Nb
duxLBWvBksrE0erWXImUv0QNXTgOhBjPQbibahOkkimFedUP4yr0yfce/FF9jSnJ6ucLMlKEueES
FWgGecsudAIACvwacZIlfkH+bJV/zPdKyJyuNP8lOfWpUDe2goeA9dj7hW+h5/DIFHBemtXpRAhh
wh76+xSf1wH2oewdvRVw5++1u7uj2UefR65wb52pDULNK2XAGWY2UHI+OT9iXm6CiUckt83B8gTI
SvBxV32Z4rO56cfCgRYufmvKTB16R9Y76EXRDAPGzhos4pERrljtsc35NShIbW9jqT2lfeFRYW2A
gY6o1P2R5oq1i47/QhCV1l5+0VODNOV+gV0EBlLlHz2EDgAykAbBJ+PourON5KENdUUk5FvAnCyy
idUORNolgBT4VIYpXPZxwF8+bZhc/VcHFJc6Dwh/Sae2SrJqmGvL0f1/V4Pp+uyiGZaDzVNviiH3
NeobyYqG7ZcYnxUtjbc0KvWXCJtZNy9TYztLY1BRX2GuSOiZVShe/ktzpu2B00vzNuiONTl2t2E8
Ur/BaJp3SCI/t/dNJQgC3e0GL6EfkwfN+OHb+/iNTZ6Rlk31GOb8E4xZb593eUiHsyIzuBWp2uuB
2aY8ox6VShkWEMwDI9uYsPjlwr4/b5wSCf0PFNwjAC/n51DfbnvfrXqxqvV22Cq4Ut4MMNO+qDnD
m01CLa5k56fV6y7tkv8Rc8A6aQ7wEeCKiaYV0u5RUS6VwWlO7Q0iRM58xry4PSgnHPdE4Grvg3YM
pIqPDD/EuZXxxZfYkyHB4GBCBvXoo2OJ/uHJLN3kerqu4amLvws+8IBE+1eFB25CXrS/paQayOQR
Jx6vzaKzRgCJZdfArlGgNsOdiL/TtTPeRFzRUiNymxWG7keHUgy8pxoqNTzU4TlJ4Kd+6KUOQ1xB
xLP9c2OWJ8ZyT5nEiBftkzQCJR/sECXRy06FgKRy00BpGXzkNXE6vMLQsu8Gt3Pl/ZuRPFSHRTp2
FwaougcNLWoY0FTPx5eHk7AstZ6poZMDepztqJlu3iSOPMiBwC5vjB2VcmjGv/CMhbsutesIejg4
ac4w8tvP791GyFJxCocAndvByI+20HFRkQVfJ+sD+uiMntLez4ZqbTDuyXXUljZNcsEak2x30sCs
QXZ3HmEIRhzSaCoH2VtW6CxDHDtHVtYIw9qGPyHj23gI5orCDU6dhJyJLjVuD+52BEPt9qeT8KFT
YFS2+tF3GL8cVs7RHV0Ovp7cc3/d1delbWGfkkAxDRcREMR/INFoY8Gaz46bFG0v9VUK5aisDU24
+Fp4JIhaG3BzTMdhWzqxf93sKgBsPbBzhyaRPDfhgPauI394s3fuHcGLinG689pOdHVmPUBwVPbX
0bC4unvnuFS21W8cQdIAUSc5rEtcS6Rewhnn9EmohSMphf4YEaPoLQ0hXMkB/mmMsFqPOxDT4bJt
jwmc6BxhOMrb0RqeUKxLfg/nyT4KMYXvcteUdW30sP3XQyZ9wlCrPYRedgyq+w5JFiv5HCq1Ejwx
sFcG41PcB2j+soLXJE7iLmQcc8bjojtSCNqaQJ6SPjSMrW2/G7prFMJ9ozzutgmXAa5GXsbjwine
4pM4aL6dnT5EgFmjJBJcdF1PRlOaZgNIIqbJRNQ4HK5gyByS9/0BLfkvg7jmKOowP3UW/fSvsrt7
JpKe3wRs7SD2iCGgC2zSjUTZhItWRi/55DjNePeAQKuIAu5mscG3VWWSWNubCz4KiEnghiBRqwM9
HBAeKwjg382EOwa95lbmpPCquWdFtRsCRLxJ5s1L5e3JCKm0c0jto/8n0YgvjGl7yJfJnWg3Rijm
CiMcJUO2512pOlxIWEmQ2i7YsX7tJS7t7NT35eVSWNqkripuO069hlG3kUw3+QfKwahxOkZIbc8T
VehLUQna/3kOJ6dfBXpvIhf13v9XAi5hrI81fxZX6MYJUp71ibad/wyYLUlLE7d5GP2wxxo9eEU6
EDJ6yLj4mUcAxPl40QOHCQyweDkof6DjnRSeRb5Ih0LoyYbXs4475Z3wIpp9+nI1GJEFCr9/fBpx
UpmZ9HFUjyigK+j7h+jjqZ5RrfwE7YT0pmV7H/1ydPIMzespN44zQH6Gyv53wPsLd0ONSgP3HSCK
9CxykQJpvo0f6h/53yiRQT4IXNdEL3/PaTZgdWKTrU539eOfmE8OUMueDJXXza1IkEsXgnO3JRad
8Chgi+3dTzvzbvo3o6EZ/1uXsNBje1AnI08WitB/fT6cnWGeISLYqXhCVgWtYLALupR1I0j+B7BM
JW5zPdgrzc9v6FL9qH0bhiIPho7zIDPn23vkVSucSXYD+7rt4mCrwPmgUHxjvEIjjZfJKQPLFosI
S72pN668CS3ASzrudTxX/IufU6dcxbShsLe7gSD1gkBmxzVM/inkbqXA20Ek8LsfCP7JZPV7ZV0X
ABLO+BImLNufvoRVigUtml8zyiJA1orGB2Mfm9pzjhUFhg7iFwLF81iQqvDfyjI+pAxkExI1qEsn
1lwhaFDHRv3eaKXzFai2mhbN1evJQqXARKh6+owYAD+cwdZu7zPTxdMGezoqK+Ye9rO6Q+fLYGlX
PWPj2Pkh6i7TsJMMZ81IJZpeDxhyYhei4c2JKKmI2elW920pfpUFH/OMzlMoNJi3s+V1k9PYhbOR
v7bpnL+UvvzXmKFqiQun6XQwLXUydbp7CgN9QF3tRLeWR9WawXVT8Q6KHhXVNRgsRLuCuF7YaaZc
RV0D64VtOg7hhMPxpoomUcMBoyzXFnGcE83Hhk95Q7b5paGaAvf6me36TEF+Hzw+h1MDloBkVr16
OLi4NbvXn0xM6YacU3w/Tu3SUlUP3FI9dRmF1oG64QcpjtvCdcfyLUDm+hn1it2iVx7pAgwRA+dC
FoPhzjWUqqdxITvEbLVonB5EXPOXDoVAUCqK8dcHLqU2yOMd+wZSAErPIU4Oiix/vTn8q3+yyX1t
x7hMNvZmhnf+IKJoQ8+HtOkGRert/JEYn0Jwg8CtXgnUYeHqqJj461JUAJRHDIATrzyzvp3BdJQS
xO71DSPQIjQaBqMo+31iK70CvFHL8icVzp/JHu8jliJtAhLtPJI4wl4wrjGV5YGmdEBQxlE6gxZn
cmJem+nPntIGZO40o9F23yVN67OYB0xO0DHFGmwaYIasBMCigYkX6NNw3x3oDTzNNaUKnzU96pBc
TDBMqPlyzrhPOr6puKdO2ogqb+o+2+3tquXW91NSie9tRR8onKNUxuCjy0zPavDsUqLDM9KqtT2B
Dqwct/PJumwOFQ9Qs8C9FWY/G5NMGwU87X9qR52fssVjFrODpAGg5qtjvUed3b2pxgRJmNjb3E77
lNn8K4Ms14B9X5a0Y0zGe2XZNuGSF2lgCGBfdX+CWLnx4qoH6Y79yFlZLcrFUWO2ukqlJ+2/9nUz
7OSin/lX6+FtmkBaA1ZTjUqRFoBvflVd41faH0W/+zF+60rHoegSeRKS3s3jITvKNyaK8WkEnwgH
RVWcSGpIwgf2fuYUS2lPYZWR4Y4w3w+jt0F5v976eeDWmvc8FZKckmvSWrRq2wwi6yQt91esR/jE
ySbN3HZnIdRvpZG2LSY5lP3Pj1T0naLqclrVzfHhSwc2TZGWsR6My5pxcFxRsM1LS8dxACSc0ZOg
6Cvn9SrzY8QVYd8p8V8Un/8mxYqtSctklQ9iuNUE8HTa83DqXcof4DxzqtLKPKBFRF+HuPjK5c1U
qbXbIDnOkwzP2g56w0yBkj1sdjo2cUa+T8JqNpCtjH0TaTyZaeI6vwFx32O3Om2wiR/hosAcdTt2
o+dPs175nHJIJkPwNSkIGMdWHpZzFkwMLREH4nYyUt+tzevfsHVdzsxTuG733NCPjlN7AiQA1bSX
WV6BHTT5I8PhJ6VtAnPZckakBMLYmDolHIVUkBVwIDKEzLyAD09V2Plx3LiRPVGSa+27x30G+NHu
bfYpKBIeIJpyYmD5f1TrNSZzu7uOS1dBP6oUsekcK0GnuwjFu0hL667Cm9cFPugIRMwSrzCGo+SH
DlBPwUEKHGGyzLTygsEkbft72r46oi/hhjQI/8Kmk4GdjCco4r6SBt89V6O3QbiumMF7N6M3nLMm
T905guPcChSsJP8ZcY5CbHBOQ++lv8q4j09+XjQqADxiFULN+dhgmu+AIXEcPifs4Qy5w9EXkwkN
o//v8jDINmti4pqSY8hGT5wdScYvBvLRoxmBLyNkRAQt17Nn5cuToavxoXbXOgh5j/kDVRoYIBZh
OcUxwhlfRpMiH1x/xB/8eeZqmdtWrgcJuISafCWi02JyIAWBn5ByBvPHEZbHugNs/q7vVokFyVuy
D3bGIy23vuoIy6AjoU9K+CqBpETIHqR8xuXMVZRGoUJ6BDzkU4ZulN75YhRHcClKiWztRVLUx6aP
kGWGE64JLp1zmCnlL8cHlN+OdjXHUwiUqCQbAJAKtbxIAtOVRSp0CpQeGTrRBljs7LIkV7kUdq1h
LwjGjUL8RMXc2JT4Uy+KvyFmMhF6qhrTM7kvelAVGzchiCJDp12PFCK0pq7WCJXdI/KzZLQDrX2U
N8or2qwp1W1fxqTaRnMWl0jr1XeiwfvB3Jwva05wL/N3xqTqv3FjlPjkq+sHpnXLvQl1F5KUBZhp
JastIx4rRIMNNl7IxcXHj59ZQyFdbjR6+UqJ6F8nOiYjVN8YXdjgqic0H1Cx8/WLMD4CgWXFAtMR
pShk4HTv50ZoV0jHHSelJLzAnlj8J+EOjzqSCJDmK7OURPwkkbnY89+wRBC1fhChplM7iyNSWiDf
GXGtRab2m6sU86DopR+LfCcDDbbIy0nVc75n8tg1sBlcOM26I3OpvO0GWwC5rtOeYAIHl/fSSE4u
peYWWKKZQ/XunFAHcl07efqb5+N8iyCGNmkijMrxk5R0WMlz1/bK7GzimKLYtAEiFNSkGss3EJ7B
G/4NiF78caXpMpYdIeKg3TiAnBh1y5slPk0uuRrJjjMHBjXG/V7zSbWNZZUvBjg9V6iORkJb5VA8
oUIVNg81Cg32FKYemj5IcJSYQGJJCIXmUapn1xG02imXaxhf7y7pmR+tG5/oAbhCGQ7X24BuzIpf
QxBDBRHB2FzJt3qlDFqHqa5V7BBupFfxs+j6PPI/WZmWNXDFToRpcW7sdd43HS0EERAYj52BSclT
UcHt2qcIzPZjRVDdO9Ofr1hkVWj7W04ahWRiA4oFYzDGzJ0nKOy9RwZiFIX9YEZ7prXccJLwNZHX
3jcV4GD+dXH+FAh50IzykXxpBd6nkK+hSB5DZi4KDxYeAREiXdSEkMpz3fQy07ulwH5+jfV7q7de
rtoJrV5miL2bnYQEySY7WX50k1/y6SbEN+SamwcysiaQ98QqS/nC6r41FxJObNKrDNG1rV3Y8+AS
othRwiEOS+1KVQLGfOmA7+kLBmDANFeIJrlbQNIsn9YGY5kiEpMLFRUU3JTB0zZnsv5mtfUGwZzM
nF33zF1tzaYjkWGRpcWeahvOBTPXSVX42apgUm9/DOrlxVk5ZFHm9o1BkMyYdNkuz71wQPCpGyTa
Io6JPcpmMIL5GDbzop+MM2hMvilAPHC5a+E5GgDHl1CHR7JEiA4b+cTzYgMlFjeuu67Upst0SwKZ
z86x3wYIjki5sIMNruXVS2S80sMjQGJ1LoIgmfFZT1+jHIwg6e5gNRk4mgXHyd0woC+us+njjcAZ
BkzKLn25MtX8Ytzj537kNK+X3dud03C91aMhmUkdqQmHrAHdHvQ9rxV3CgYjhkjD3O+iM8r9z5Vo
m0Srr71NKfw/dQO8N+tmKR2oZut+IU2U1rDtbiH0/Vt2C+ZRa/FGVmzo4gZ5ePqx3vYlAcODEysv
81aAgZMfHo+dG25Su6hF1VlTVvbORZ8ayIWYFBSiQp5PNtvhoRh+YNEz+kL1QRkkLFjf6lBCPVBg
N2iFsp4nF62bavqyIcLUZ6ETNEEooYgVTdKOv0Im6fazKh3VVIGXfPoSgGFQvTA1jeyCiXGfI5uL
9/8dJ7GZK4oOo2PyZI29he6Td/2MUNwJTUzQ3SdDLhYrEKyeYAo2Sp6ruJmhxarvHoKgxDh/JjFg
YGjWODfv/G4hICmwbWAWpVsho2qMMi+9wT2xbewzrqGIK7uJbOqQ3fJwzjswDv5TxoYh/zYJ0I+B
m0jO8szeBYcu5PJQSgVIQp0q1uChzYXXg2w9Cq2Uz6arK1tZobvpyBQlhEQoW1ipPAO8+yx+Nm7e
q+scgx8uh2lBv7vogMqAI6BpmefV2zXO7xLJqWh++vh///KgTBbYJs/ZGUS1xl2nuFEIPc3QTU/p
11JtvKCPD54lapb1zMUuUvuudgw9KU7BRQ0Nf/NBDBACzM2Dcj+8KwCiKPtLvZJR9ZvRBiXvLBfo
aEIssfUbYGuUmBm2DzF3iIpLVihhsbUzreWA9H/Lolt0yScwz6wSKdCmeVJQ36YN34dr1BZvAjru
TeSF17t7knPEN2ERoG2zKAt4OdBkg+lEaV+H8ev8EbD4Jrm4SG7Y1u7mheeXkLDnVcX/YLATQgBn
SNyWm+zvYKPTHTH1bdHjiK3rkPbxvnnLeV5MZKb+GR2NmD7LBVVAxdjXqhBTtDuzMlCsty6RCYdI
SmoZHODY3mRghAFkpdzSyJNbDl5GrtMm9UnrdO77FgkDuV/PLDdAA5KIQhHz15Ddf13BgDfLDmrE
ask1cv0Ydy5UaytR9ErFu+9RK5IDW10NJYMbLCqcPNmLjwNG2SoclID1lIO6ffBsrtdm33hImeFM
tThFv5eApoj8K/o9iVhfxKqBHn60aHCn9kM1OajBSWIWFJ4FItPDE16KCuutc8Un/PJ4hc7fB8iX
C40dyayyRgWR0L8XH0KdUshkehoYhD13x3p8TFwfOvGC4Pd1eJxfmMzYM2Mv53J6dfN06+oMaQZb
zTSmCagw8nN3lV7PluMJIzPyyGBuktNqmgeBvlb3ZjOeLnLS6bNih8GrLnEumugkB4IVdOgiLR3G
j4sQbtuHfkLdgQkMB5xho95WYIGIbH7OEHexWWlT029T3jjV3BB5Y/4IERPLcPuBhv6C7PMghdT+
jCgbOFXllqH4hrvt8klqyLdgDasdF/b3EedljVfz695JHt3rfzfbmjQkd5dMOmVWaezlIrrDoJs6
CQyugCU4FkuGpS3ZgmTllUuJJAZZ5miso9xHp7+OuTxexTmg2KPlbIOf5UvBdOfxBvRYa/QQdRl9
XKIW9IemMQwEoG/yLJvM/4owYs98FetDB9KZGHsNtSXlEX9H32vWJZw6GkVQc+2gN1aEi1HbFV38
JrkytLs+/RZg2lWJVocOPTS0pSintTxpzvMTvJUFk+N854X2sb5Y09b3+f1ouwgkyyGFLHKbvzXq
TbSCS1xxP3fVtI8lGJsyU9Yz+z13XX7tjhY/KXJK1qofcBp9kM8Mz5ScQc1XXmV5cyq60c5b/6vz
Xw/8q+3ofgWrxbxnX/nvVgE0He1f+Qq2TtJG9bs4VzvNW5/l2BxGIIZxvUEx8WHCiMfTOvuYmxHo
7cyogdT9zPuuCcu472zGB6aKd7eIBlGCm24LCwCOjHQ2HGq/UE94dOxIjBk0JfJCulRDdRA2HGR4
xfTNZyWciCJqN+L4fxoKCc7pGBwVF+JgzZMT19FsvOCawFm3IvI8zPe/ObMtyWJ/T3cgKYKE+8eu
nbSpwdH/UfuZvVqTG+M0GdFf09fS/7jQRmxWfuWg8uXxE2ZwBsJ65dUOlE7fn3RC62QDe3GWi9Bp
lcpvyaMxZoexWi4lXdAuDA6ufEea+74DnfXeJ+W1uLGHpdnMi1bqOOwwb03QEqfRT9Cn70gtxnDg
MRA7kqyghgv5VC1aqMGi/dIpTtzdeIFn9iuR2uJ65Cu8rKAiSpFwvqTrE8ckyiHDNloZ3RQlMIxo
5kaRzDbpmJKPFjfif2LZHQ4nqxf6LHm/1W64kA5AwYre+aEB27bSz7VIWol+F6H/9Q8a85CbS4Jf
93zU/WNn/D34uZrISoUARESm0z8R3pGBiL2phn+NOWS7AVubpuYSfdxpKE5lwJIdXbqHZddBExsT
4u8vs9hr57Zq2DKgyc+je42sl/n+LnTaSC9lV1EXgkO8oJCfBqXKKQrGIEuP3PFB7cW2Ayf1zC1i
Jon7IdRTnzEYw0B9GTX+w4ibuxZ+G9EH0bb72b5kOE26vs+q32XhTL4e4ROo7DtUw1aRJHIo58PZ
IwXu8cuk46CjjcWzNdKynxcR2jTm/2TBqE5PmVTAIYYdq8teTG8jb1IC46tizTwaX1VA65ldjpzT
Mp/d8UJBQYUBfkYvYZsaTgCJIn1SN74182QbvBh4FuT0J3++8G9udrRF17OherV1IgAVmllz9WYH
z6/gPYKaGBs2meDQrG4UCTSwY/lL7/pWzvTMoTHHhXgZOOZUGHuMz/QlAI7d6NhWwIDnI5lWodP+
rs3pJ2aY2C3Y4ZuKXqaBjSeiFr3H5WXDqAXxakwPEZQ0qncHYPup51aCB4H+WBAECRCQOPwh5z93
sOCUS1qQFGkukt0bQ4Dabj7/+6B7u+4WSYjRDr9Y2fTH2BjXR0AG9lS2EqziRRYvkujfWdno1ao1
geqqpdDAChMREkwSVN52qQktVqX5Q4YuGpZUfewZxPR5yE2QvIe0HbboPf31pW2OlHfPTibLtZ9X
WsScqFEjblrGdFZZA19LWLp1lJW7v2ziYm8zyicTPyJ/nANsyfTvBGSIPQYkNeiSqZST3guUKKdu
KFWhStLF1wJMxuz9LtDmgMNtdS3rsO2oVWIMoRrrANSpqc3gL2E1Y2XzLG4JBoTjHsp+R6P7yoyP
fPkWceG41MKN2uw2FCCniam7jbJgynM/lf4Z5pReMUzc3vJ4O4/bnBzUuq2c6XZmw24M9cmeIS4f
iTygINThxFp5M8nJV6tVk5/ibTfe8G39YfR9cQpZmcz8GGlseV0ZsaJDv4cKvSH13S45cRJiPns9
dv9fuUZtpbpkks24f91ePIUFRovRvi1PT06beUuR097Y+Sq827fCwyrL/WckYhZKiwN90QTikcAY
taputNpp9ioPeyhccY1xwTMNjxWr3arzpkT2xYqV6J0o/p6JxhU7P+AGPmLzqBcYHWDA+NbR4Jgp
0tBoPWBlsQf8hXz0GyzVzEJz6/IW0FuIHAl+AfAqqRD+cjIEZTSutP/veNW+cLNAoc6swRmS9K2Q
7ho1GrfyOXNSMpCFQsc47s/XmOjo5tm+BhwlDgY+X8lE/aZHS5W4FCEAowU/VWDwAPGEktDAod8o
KnUCl0cu6CLGgoEgcV5UtrJgJzzj+1lUgu5F04d3kOIhmr5UwS/JPtu9hDMJ6ynk7vl5X55BdAer
FqHmDp1k3etOJqwe80NI96vYeeQX6zFjklv5lSc+vceCQwfDCh7yjwqIBtDWsYw0BjxsfjLu6rKE
JE9kaBhAM9DjXdgIzRM9CT4W2e1h51C1Lv6m7h69QhVQM2EqysDMf/PG/7IT3SeIkxdO1w5dn/cw
S8d4BheydmzhU55ZmbGhzJfOQ0OTjzwZYbluYF2CEJSRZVPKbyOLslHzTGz7OI9GQ36hY9F7+50v
AmaufRgQUzjwpCVcEULyzM5L887twPrLxbFCq1D4XA97xme5fUYl2ouh3AQntZmb9veuZFYRJhXi
LmlP7T2X+JQFiNygXvKChd0TDKs1HYs2Uw2rIJC74ETi8m4/UfR6D/EkHP8pJAzKTaeOVkIzJBeV
If166llzb12sOUkIy/AwqzzXn/tQIglg5ADOdgikCOTkU67TDalkxkdfeOxWMOaULHwB3RSWL+jP
Kwl21VNiPyCdDipWy2JGxmk+z3Ed9FR5h49AKrdQlHL4dOVyg+HUt3DT9HEQEjs6jCurR6Em1/Qy
M7HcnXTvM6Hv9c33iI0jPvEri8K4XwqRGaKo5ulSfBfWmJJBF4Q7z4bSDQZKsO0vy9WNEUQyMyo2
EBoCFkL8/RzUwjHWs0N471oGDNyjJj5p/JkSaei0HGLpB3o2I6K5lPmMNB54fbvrVOmHZYtVH0pR
V3LJSGyDEAXFko2fZXzDeKUdiG4jSDDk8p1dc0AHTYwnW1bgbIia94YZF4pdO3aWfmIsfgygySgF
hik4KEWhsi6WafCUuGNpJCcT+/PtqCnnxfiBKicEKNta79FllsgfEc5pJsTonHwvQ2nOH+8ZRIk3
7eoBgMIx1nQwuwTLuBeqMecPxxsycWgY9iVehpXOYUE+SGKqM5XqG1ajelRIy1ANZoDRhqMK/rmc
kcq1RcdrFw4+qahzUFjXFZhgiLLntVOEeY+szoFZagDzJpj/TGjRrkLOQyvamQw3SfeNuioJMayv
YRe15eltS9qSnoSC1ytIzJe6YxFae4A5M6u1nXse7ARCrb2p0W/FczIFW2iuXfdF+bcdf09oLNCF
xb0dE6aF/fNGNwRDxFVwaHrW5bRB7Wi8UZB3nE8bxBFMuwRrFP5h1rJ9qJuStX8DxdStrnC0XYMq
WYOwnpG2v3GXcJHlrpmtb2+TFnYcgmiMxcYriLVjpaYmUmHE2l+LIh+hTQmymmXXn6QFiOHVIgPJ
aq/JDH117gWxOwN0B5EOUvwmvmK5g4UJEpnWTOsybGnP+NGSIsoMF/dl2HDuypban3HkKVN7kblI
3yjqnC3w2CrnAC9fyR4CCo8/q0kJsjPStlFVCGTSMXgf6ujHlzfUSQQKtBD2dQG+ABWQnNIxaUmS
FdbOWLbyKLp2xVzr460x2MGdsC0PwLS6QQjLNdPkEApsVJA4GgIAyuX2Ovvq4Kj33Qbpo918/O0p
sZyH/keAWuE07Fdp2RdARMDUv5yDGGcqLrZnYGHKIbxYZm5ppw4phZJw6k8kipnzAL9V8vSYPQ4/
nppC9oDLZJYLLUNMW3a1yrFmn0AOFZXtbGBrC/FeMzk53Jv0/UwNX/Z9I5+kZvLEzJ2Rr/Rq3KpU
GINSE+IDIsiLHg8yYedZqv77cJbSVN1heBjy1lKLR9SkXpMLFCtv193juQXW02r/PMV9f3N+iD4e
Qtc0lK/6sRpqMWlndAqvyexW4ziejB9+d0a6/0cQr+db6Qqn9HD115juU1kcCZ7Uf+bA7Q56pvFJ
GR+/qQDyqN+Cozjjy5J1wasEmkdFau+Qlm5raOmrM4hqTjVPzmT8DR1ct329dSIuPVrZ4MeEeObh
/DVjCh1sNOlL/ggbc0ENsXH7IeFlCFHNpYJh14MauuhXmRTHXPLWd4q10DD5FQC72IRcrRHrEr/A
3d957WyzWjrjNHGGNhgdm1SZ5NcaG0tASCWovc+MUKPsGzFmjIGoGkzoxFb8CKWyteYglRh5vszt
si/6X4qZZLyUfb70AQob5x5EHuv9lyi3tbu92jSskUWyDDbRXdbt+UTqC7/kTYqplR40Bfi1qrCF
py5RRjlLIVU52Ol3fwATo0kk7Dgbq9Mi7xU9A5M80M13bKCEwv0D3S+Wtox4ub1em083CUjlahqk
AkmUwOzwCOpCH7hva1vmGnhVKXUGUSM5zmWuLJlcXezLeYZIL34JH1qDwlu4FFAouWh7EgzPOSBZ
M2yJX90Pdb1r4YkP4nfOOKeufXEUk1gQziRSBO35wcV7zF4w+BY6cV1FX1lY4T/EgYKHq/iygxAR
nFCRgilgnYENCCnfqWmlNSm4lvkcJbjnOP2JxozIXgB6vqkhisosIRB3HVlfVKpU5oHjQ3BRDu6D
ieWnxzT8gvyc0MwL+RaAxqMW6mb3bvHGiAECqDvATH9AQeaBXMSIqFwXMZvcTBhcZw+93dNVZxWz
HnFja3p62hFipqyVV7YTve2+tNkQuqxNdnb8renr5sXCizt3E3Pf4Ow6uuee6OhdVf9uGqFt7eI2
iDjVFXp6dsTp5or8HUIu9Tq8VWeX4aHthTsiijp5X8EEgZP5l2MhuNuKqYtMCeGKjE4vKSr62fVt
txHHQKVEwQ3H8fOSwCpTH6Cg1/bXqBoJ0u274RA7o3Fhli8xVCH0zP9TLK5FOIo1MUDU5JGcvEw0
+4ApYiPXvj2Rcsjm6Z4U9jNX7pHdugJmi2ysYLYH3Ff+ukzGN2zbVclblp64gRgPNfDAlpgnZyl6
H0JKvjnME3IOORC5Jy8AxB9rujSaAK2ahvENNmBRfLZ1Kh0Turd3lvwZijXAfsWUKf6ENkbipqAG
H1fepLdDv25knOxSRpD3fxKMWxRmnRkFVvkBNJ9iH/YpfCu92AsHea6nXyEYSfRId7vqP5ltyuz+
21ymh5IU/GLw6nSif2iL1SooevIqWX9DImy5QpBjLuPLSn+znOTO4S7nRTckPRLzQw0tbLZS2eLW
RyHumUdm2at70F8D7ACnJbtyKWZ0Qks71OCCnZK+6Mmtj0zdK9+wVh4aDlkyjVlmP4TZKvZhOS+H
S0fVXaol36ZTsDFpZ5qZQMKeHcldt65pQrA0c/uabmQSduUxTGkfZA4+9LlyBTCrSZoBG2eUmZ3W
qWPvJ+OBUEdRwKd0RWjZ4ljxOXq3hHvnCPc8DFk1A32EjGJfcsCQ35KWX1hLDq43t9fckHiIp4iY
c1Hsoluh6haxDGSnBDxzLvYpy3isIus8FnonDVuk2T6BB5DKcfJzAzA/ChxhVJh4VnI/uvzsZuWR
KmVqDMcc/qt4kEZhFPV8T8DdVOa8okdzPrtAJkSCSwKlji1VW5Pt7Q/hNrbJJ3HiGVxpDDRWF8oD
0l/I/ZLEhY2uta2VcHPk/3N4HQW3mIBeX3rVs8/1pnHT5UWrREhMBaaXnuEwDEFs9KQvKD+OneGH
Seg0466BQHeihjjnsarBjzAtFVCzn2FNGRcS26HnIZk0A0thLE7w1fh6YGWLj3C4peqCMX4xUKXu
RT4xQXgCchw9qK6ywUwZfeVTMQBFz5RFr4UEYZcBvBDuFOJM1M/MDIe8S7PoPTwhWClANSeLagfQ
woPW2lQVpw1+wqOWAhJQyZyZBp2tUmBBlPIBwumcyNhEHyvwLtSOTgJ/vS4wa5zluwLklihAfEvg
KxaVmkReFelB6wWOH4KSWUn1E3i8pAs+JUp6Z4BEsjOfu4Jd0j1275f9VATfvXRf+ZmDAxMrOlLl
SRYKKnZhDzj76GnfXnheX4tMNUP2SXPBGyTdh1nzOIoNLEnTtuT7BCq7CtF07hy9BHLenOlR9Q8g
b0UAoQtVSi2bNTq1Qn6L4cjdfWLTRaSwjj+fOhG9hW29fCYMa5nrbx9zgP0lDdaF57Vem6f3CQ3f
Mruq+XPX91C51SI/BMNKuxm1/o5YvDj5RDws68m9LrZBM+4Nh7GkcnIJuE6VPwQqBlfq3cSf4qIs
5PWND9ZaxkkKN8muIezrpfm/Q5R37vJm+/KxDxSmxfZrc57nE+rIdp9Qtwbc/QryHCWzdzD/e12y
nKfHKoQ+KEF2wCfRXefiI548kHqcohhi/Pb6z5q3zZrJwDI6c/jc0XyHkDsSr0WTSPFr0nJBJY92
0AsQna7Ig1wjtr/uSP76U1ScLu4WvxWni0dRfOLFOlQrZHD8OD92u7M91wMuXBq0Wy4th56UA4sB
FqAkGbnRVn7f21ehAKArMNZu8aCQUAwkWIU6DoAN+rRoBGl7PaDPkbTzYflju7Z/F+iF6CJb7Pv4
djNhMuGPnV4Lwljf6tO+WdsOOydqRlGaAv4gvVEhwnB1uhI90tqtEYcSCPQw3/AZFnklLsnrbk1X
8dMYPbeQ6bxVu4yNFCTz08pMtU7RDice0z2gOIv5xxqpRCwxrSqKtYl1ynTE8SDeY/TLqFwr/EAn
sH2oolQfUuu71Yv7vR2yzS1YdALWnmgWrKBDncTnGWcEDc4GTqIYfk2K+5kCOzLu5pFlQu5Zm5UK
gzd7g+C6WYl0Yh6GhoQfI2o9A9nSXT2kWDGqTYrv0mhrSvQGj5SR+NaoMn/4ihu4IpJ6vN9t77Sl
amoW8l+5F0mxkMrioIFQEJQVbpwKx1ANC2TaKp0WKRuQoGzNh60AeFGRnRPT3sgZRevduxgVC7nJ
H2vpYYPbdY5FT/65hQWJobUbjBs/XRtZgQAup+1eNWLjmlXOBcCg4KFxAd0jHrLz/F1cxkWnsJAg
5J8g+H7ai9yZxrxq1UzSRFTRJgtxJ8F9+Qjo/gKavVrhlXHjZG7k6XGQA/z5/W+U/MsQMJade9hk
VU2Bbw4cubryxjJkpNcbZQyzoKPDFYhDONImUMMlt4qfosrAm19FNMj28+BHkXRVJI41Ssj3j8If
2NXqjAviZv/h97IyppGU/7UlMM425o6jANeI1kMIIHheXZ4zypkwvP0hmFoHiMUB9ix7SWcMG4Ms
QU4zDERthyfc26KT7HxNCD6d87mRl/6BKB0BTr203qrcv33blblAa8hCaNgjdJ96/k8BRjbGu33/
gdluHP7IwGBIqiePNjUy0FHzuUZFu5QtX5Ty6KV/8U84TYmsaKwoa2jDyz5hPjcoxPRGi/pGnrG3
1u/3BqxBtWjfSBDhWk6SIMYMbFhxcCDP1wonR5Aw9Ipl7SGgVoUdlS+qHbDIkAVUwCaS/drSqVal
Cp1lSLFO+cz0YSPfCaqKvm1uAMTrTLZPRnTXNoqNSqtfpCp9O8C+zov4qRlhkTwLDG305T56dsjq
Yq54K6hpdwXUNffWo8eQQ8ckibM795A/gy6mm80ENRVB3hdhF0bBBTwb7m5QFdpG1+DdaK2bAY1C
XzrOBv8zE2ezSC2aEphi/lGqdKcEItoNcmgixISLbV0WH/6uaOvWZTKFpyn0diXNe/ZNMgaM/RHe
L8898fPeNcP+SqmUs+IlD6Zd727xgk8MGezZtgcZyYgxPcnSWnzROXs8DlFkPgFsTRd/K0TZ3MX1
E2DUn0+qqvgfDhyUkSZyF+WkR8ZjM1HBQYSYHlWPIlOH67Sp5gie5jQFNkonPKH26NjZzHOgnqZE
y7Is+FWdCozC7CTeriR7t86Wlqr1vV4vv5hkSWYupKA1RLjU8deAjvw8pQb3PcIH9aN2oAE5/O56
oCkSLjU6t3b1J2tymr/GqxGWtScH/HOPookuJ0XVFhwozLcaWt1fT3GR3/FkHsCJQ9a+Ghay1KM5
FDh/XD/wAVRJV9V/UpM0yskl3sMrfEc2TyI6r4Dca9DDXkvWqpihEQphSnvYdcDXpX/IMnj4mCbu
FpsHSZZbkYBgyN2TtGS++iKioNLzCoimTd+qG4/xDG+ovx1AljOo68uNj9IdPgEQflD66l+Sbspk
fzsfO7qdJ2bQRpLE/h2vH3Th4NutVtrOPThCoJ2M3Y3naAZ/OIXXozaqnFZT7ypaxnXbq59M3opE
pnp2XzP/IzFeGVomXntpRuyrR96rZgs37nBQnA1/HfiZBvlvdDwZMNBTAV5UMxC8f1l2nL1RaI2W
NcEDgVYKCf7tseA8D1HgvPcuS7IikqoDUu2orFuudrPPYKyaiMqB51echSsXZjUVgeqwgzR2R0Qp
q8sxNxNbg4v+GyBwqXqtLrz3tJgr3SnMaeJh3QRQd7LjXPiQVflk+Bzi29Pza4FZdaw/0Xc4Rp5C
FFxfWZvpVxmiUDzcKeY5uM7bYhwNC1biJF0iQZZQz/RSORZxtyFu7/PgpgkxoGdlsAYCI/LK0C9p
CDm84QGCH/occ7tEdKv3xrgvP6ugarxfmbMKAnRr3Z6L1r9zcMXAeNSdtIAe/3QFJYgdA48O3Rem
0Hs/Ecb0JZBs2xrXSByPw2SzN1odHm0d+oCYxQCIu+Z6WcolD/TqkLz0zpvCTNj+embbQuIseFBD
IR3p8+BiGjD79yKX4WDbpcP+xj/JqNG5iiLvQjic5/1Z+B1JciN1T00g8tNu1z4AqwNUNLzhjYnr
BlAvRJIPD1/cMFc+r0k62jITfVGKFMBHLP3BemR5kqNU6Yjw1luutx4RELzHe8xOdY7Iaf374fe4
HvIguZ3Otm7rpfpu3VBrw9UN+al8OvT3jyG18rkRQq5DUVVl2WO3U1WAn1Ht29YS0mREVVq5RqQl
CYJDsn6DKpTh2WQh5Js22OZqssb923uH88byOARz8o0C9pjpDJ+uMG8dM3+hrMQLDdfQgPd3EuLR
76wb1CbSzABHDfLKJl/sdlAHLpj6WL3rAUo84v8sRQs5UmyzjA1g68Zqq2eDbXu3GBZw1NPONAfN
X//lH9TRyD92cuVOPRx0KtnbHOVw0we6tBHbODOS5xGXtOAcOrOA9b4HJaDkjdQ9QJOqtM2ffquM
NLFwZO00fMPYXAslM76Ryquq7ugSOOWBCPpfdmjeIzGgEoeZoFPwsZ9JUA1K32yMe44CQTcArOJt
w6cCG9zXFaVDXW6EBzrp6vik7VMtch/sfYiiQIZCv8/mRscy+NXKVDkecLJmhQVCGxIHNdc0PPn8
tVwih4uXzFZzEWiBLsUG4Zwurp3ShqGXk7UXp2AW1YPS+o4axdeL62gkeDY+bTSIusMz8arcGgNM
QtbyV9fW6jDhG/wuzx/5qEoQE6ZqzThPRqZhaTrzpCNTDCjNAZJvkxzllz1Y6upV7wgCxPngzKlN
g0fYQNMpqDz62T2tmBs0A6vjYKskYNm1qu+lBF3oFRhTL9OS/pmZNyPElDw0qRUhhjwgJ5MU2a+0
FMsPeZ5Wk+q4/uTerFrvHpq5t2FNt8iZyOr3T5cfox7pz5Xw13TCBvc43B7TsOsPrLB11fGgoK6t
heWTsuY7VcQhd0fMmrhagCxol6qXawbya4TZMPbh2e2bZlBlol55Sbigf2FECh+vpZOCXN8qP17e
ZBDpVRSQjCn3iMCjzO5XBkQ61q5fPuHRnlqO/or3t3E1hcfQ3BCOUFSxsLDmgpEslo1ojaWwJ3Ho
a7DI5q4Ml8dCkfEWuJ8rd7F/sNQaVPIxIdhdAvo08ONg4ZfRcJg8tSHemsnhB2LGVqDV1giy8+Gg
JAfqQFrbTXMGWtD9/187ceNNcMfcM9gEglIP7mTgII398XmCRP7d57Hiq5rvkLazW04lfr1D8ajA
XXqi8L5MjOrDrp3OBInaAF8ti2RAWS1MfWs9vwDiC1BSXMcTuzwQX6aDpN+yByAcRtlgJ6SRU77s
1u/aP1NoYMqh4ip1eKPuGi6LdfhApZgrMv9h7mgEr0uEVUyYfKUAlzaIhCM2An6uYjeXB+Zuc/GU
63cNXw/TAkfe1Fn0m7w5eFPdDGzNtquxs8h+ATV6UFW/KkOVNEJFiPBt1D0V9R/7o5NVNL0BofOi
u1JVJNfJ1+mcT2+udOlDqmwXbL3qg3IBbMk1sI6wmSg0SOxH6R7EPvYtaB6MRb3manfYwHCZWtIM
yuKrcO08q6Wq3FG0ZqXqNoqWRvcZ6XJXL/j5atsTwzsmX0txaGLdN5a6efD2D1mousL7qZ8xNQMD
4melGsXAEpl9wH57B7KSk/F/YkV/jxhCTDYbXDlZksht0CBNZh7bmElmEN9bksfQ4M6xY/oLDlvh
gJbO1W8QwSPHNFIJlw80CKpRYV6EIOIL6+tWUxwN9PWmbRh9u089cZIj2MWCY2HIKYeI2bbhDBdu
YL9rxe1g+aLlzQrO/H1Yu3aEDBrqYVzX6TPzsPetKe9kKvldMmeuH2sXjnANRN7phaIRNCJXiRcd
MsP6btjjcHXUXWJf3i8uVDpxQ0SiZE0VU+wG/lvMMBeh2a7CzTQsZcH1pliTzfPsZvEuj8ZIgqLW
h7gSfpSQ5nMAZWkviPprYNfI0D0+JOVaqJY54p4CENfP83mJyyZisknVb1JoiMUPPpOD6q6SfIQo
LHyIDAtD2C3WrR42OtzdkiUVNvzFUxTX+MuAZDXz7y/U67FlAs6nUq4ee1AQXiotXTGTC9HhLxEU
wwitRt5fOoDHcLKuqYQXyAakWrGlzxUVGpSJ3wnkzE4J6+x1l3TPwVa9Q4s8xGsNzbB+brwVgzIQ
4M6IEVBhS5Rznssx1SHn/ghDz0snBkt7WpyoYQJjI+9WAgfMxCQV+ofLPnumbAnt28hZHU3QWWfa
ScenTuOKqPNn92/KK2Jne+6kVOuZWrcBdkwl8LUI3fATt+8pew+FS8HffBWdCFMgd6IPJZIoEYfC
77LrrYG7EKd9oXtmLvrKSYY9Zdu6pn19PWQmXl4SnnyqDtYWMiidrkjam6cWTw3lKpUBWE6gmJ71
k9Xf8AF/3kBxO7UKnQmS+SkS0ATrXSGcWUrmqXgYyNp3l9D5aSfVpQYwT6UQciqEtBg6TY/gN0fE
P0iqDrzPoBc5Pss6fYL5v2OSNGThGXKTqGpK2ZlJ5s+4q//Fwd3XOqD3fXGrhgq2HhUqekTJgRjs
dfgGw2apz/8flUx9SORgLD3mz065ogW8vvHuapVk2LtJPoW5oqdk+RGdWCOUbDrUh8JIShHtTXMw
wWir83SaNd4QmIfBDh2zK3EQ+TJdhho9em9w1NMoUS50wJtXDMaasDvSAjvr2nYBG1dJHzRBlz/C
ea/nTMBJyMn6WOimmqpghBUdvNeg2ZZLITX9dVWNoF389SAsZHb0B8p3ogQkumb4g43Ny9JtiHTt
KASYZAUBrW8BgZORBvwPoLigpOXL8PncQPyCnzWxy9U86537btYZuWP7BWqf1oZzs0wY89sU/+YX
Fh956/cXyzKjQRSLeVlfiK8hcRXT5oUhVRw/NsCrLWO5Atuxe/lqEWALTXQjzvC21ZxnZ3ZXF7hc
xvzdpNTvubvbzw9nzFEiMYgH3qsTanAyo5Yt0l3/XoITz2qKu7CQI7YATl5i8R8p1keWDS9TlWh5
BmkcRb9IxxYbzHBpSzdwY/Zm24uoOsP0GxP4l0jIVzUeB3uqxOvaN8COKqP2twOfCeP7FujVtfzx
+dnXvg0/zCShBn/OuScFhg41O1ggkSAfeJYm/4RZfAoDrgQ8ehA9rjxFDwlshXTKo4B1oSIKasaZ
IrYlnJD9OmU2AVrcmhGJYRkxZlsqzoMJIDKnDdMqf5f4avXT4M61qkGdCwOhimcwA/Yvs0BMBEAz
i9AW0F4hCMfcJQdPm2MJIfhSiLFb1RS9MQYyunhQA0eRtBUoYxVY5udDcRzPmw2+aT5Tj/DJC4jw
cwapbrDg1g2e2957iKtubmC+Gpp73TkYqcoGiB6cD89sE4IPOO6QPAfb2WDp0LJNRkwJqiDZw5Cy
xXXtFYzWeEhB+80nCobYtaQLffL4ai+ZHWSvE2STSVWWBeSfQRdO1Fds59NP14v2a9gxm311+AmU
qcu2u2rtskovkC/cF7kO7Fo8jqCF9nHWpiqdtKhEEByemdsRPAUnoq7qGKMV1LnRTypgsC8WAgc2
SdhG0CZ/GtGrJrnU+9VDzQt9vRFxtAfruVx86NdSd4hqSyAoilZyMqHUBUq18cbJpD+70OgmVs7h
R+/Qc02m6IXD0UWMgRGwuMSDJPvdAezUx2yRh+cEwXvOpgWPWzAr0DYob61cqZxvj8sjp0SMLs8m
5P1ztwnbE1oKtovPLbBxSJUBUAsKkS9wiOxk/cig6GdmIoqwjH1qOhihoD9/DKynjjw7ZJcuLps9
ovh/3AwbuErd90uMPpuLxQLBXyOHXJ0JY+lpteOAL/Gk0Fvbp2Umb6f8ORDo7gg3ccA/yIRaD2Yj
KNn8I/cpzS6tZKRRAiITex6/pfmI8jw3XdgQSUNnzsG+f7qmDVTxwjrFN94/ryXTJhpf1ksRP7L2
0xcGj7Eku74E7/zpTx1bDPIkObQHXX0LmeHq86HdKjyQbMkMcYSD7+RHUfZ3uxGT4/QIS1y9m64O
bdIfKAGM/6ibordbJc8CY58JuxCPrIrzATl0c2tbkDUXoR92BvexB3oczKovYM4vpilgPLVHl1tH
+egUkbDXHIZcZmQrxBCaEcqVZNCPyYa1IkC9aVyXtZXl6vi2X8cL5GfumpOR3NxYNkMIFNYIs4SY
eeF3v58eAStsxeYysotDOtFg3l6SBjswr9ndXKWdOZofyMcnUCWkPEoKAOEqaO2jjQsav70NE3Kh
CUNu/4OMgqI+vAMMRc/30orWBt7qfHZNA9BpabTYi2UEML+HtWN1aJtPjqOJkxuaH9ZREXecZGK6
XUfNk8QQDx/5QoW8qEAslhZ6GiqxMU1GEq/DsT155DixR2JaR3gt1biCwQ2tT2gkHCCVznnV8Rt6
h4yvXMK4FHpuZftivSIHxzu59IwGTtTmNWbxcgcTjc54dJcnvFsXn56GQWNirieOt50P8p06yOhR
VoKbXDxjbTSLlBsNNKoJYoU52SP/s+U0yLDKmkCjdsQ4GosXBNvmqXfEmq5BljOMVrf8GzhjF5+2
ZXk9ZJyEolDhYQKEFwt0icfZ4Lsozt06OvTF1eqJtXpk5ew+pm79CzeEXcZbPI5c+36qkyEn7lpG
uiZYkJeDdUS+OTgfEtoNXy1c+ng6lO/tIKEHvXmV+Is4bK8xIIhmMFDywruoXMj5v9dp+DBlzi1V
QKAjRbiRU9f+2XJSej3d0NwHjiZ+bMGY6MYR7Tm04frgLeBdA+yQSw92rUZNupqeMmvjvo6xEFYb
CJ3laMbAQE+ROVfxheEGZ19Vb2bpPFuY1reBiVQdv316wEbzFyTD2fmysaKh0HXI4KLFWOldYO41
DBdsFesJuSu4SvtYjcMacEwz6MM3d16hC4FKl9Cg5gQc1CLoB7anhOOaVtAhZKCqNqBdHT4Ybgrw
pFSVu/kwFJRe75NaQX6DP97mbhQpABKL+S9SuWlxM2xy1ASurWhG+3x6ChCmcjuhwl2c5y2cPYyb
zy8jfhXbgWVr3qTktM3Zx87CrLHK3e7owmHCvky0vNHH551JOj2kEL84Il2ntKB4jilS5I2kkoM/
ZQopMr2Q0Osw/mx77Uf4ZTajCuRb9w/bVFqvPbbHzLrC7GjYcsLOOnlvkgLNcwITG79Zr2XKcQdl
ovaeCf5+VIkXQvTRCaU3euATjPk0UtsSkYjo2cqm1FDHwFtkr2ULh9FeaanoyPO/PJjuySP89RNC
wB0WsxhVh3vw3K6qUxqw+PS6kPtYPGZ9D79bB+yes6v6Cdh5zsCiCF0GyauwKxFcLUKEnIK8PS4g
D5VupJcv4nVpf9hqMpyFOszhlCxA1kMElmoE5Ey1e+eo7v+w50iD+YV4tCAVz0Kln4NcgtXK3D7v
5/1wMNccitla+XUJnvSPhRrD6UNNFvvPKck4J2iS3M7gXHZwYVdvOFU8E+6Y1RuGzX7YVletnHg4
V7zL6FymrBLAIOOuidajFT6QyQmpMFIqgYp8ohaov7DElWoGA+A1fXUWVabJE5sq7yBw4mvJlPOs
MV+RLgClz0vSUvl3tU1ft0wpAQZh2UJFhfhz5xN0wzYK5CpHaQEbuKgZIzbMeinY6gKO/aP8wCq4
6lLC2eFHqx5C8xNaa8BFmC+6uP/frTw463Fsg+C/E+qBm/TLrRclUYmuyFrPPPORRwVRDBot18+U
rnZf2kUKq4f6QAyUsW2qE6Lf+Rhjiz3+bOFy3cn8Neo2y7RxmNyFjrtg1fICCL34R64L5L7rCYQf
TqlQlkCSjU3MwBT/SPy2zrDSbJTkctYdZIVtW9X0ExSR7AwPbCmqU3Ux10v6SR01QY4aTb9kjm4h
VK7dXOMacSUWcRNU4BCJtOuCLsVxom8ldU5i72GCFpqujU01xtY+xbmmKaSY9sjkqG0sC+5eDMKD
JvXAMcb1GyNnyWIpOPI6K8Vfsaygef8wf8fVH1KGs/UBg1TejPfrUxiMLwm1XUlhDwpCQ0BIlCNz
jXYzmEuERn61HJdT1aORvcn82pYRgCKSQhuxmEzxMaeymlF8sT3EKN9NM/YgIbBtCIAdHUNfm3Zu
px0Ig8xP4hvvdOBzTk10TIPYx1ImomSsy4ka3WxDIvbairYJLZ/nplWSSxs86+IltTONX6P1eDLd
lwtLqfzy2x1tC7YiExCP4YC9pVImHOwgnMyR2mn63hY77RCybD0SuUEsmVlj4Vr6M2q0h47SxRyp
OHbN6ylnN/BQ0mf6+Ik/zbynkyYuXXlHaw67lrUoSqeeDzsGlxJm9APPDCLKbAHK73OamnufJQHm
WOCfDYm5PMKOpukls4m2bvW88+QKp15SkraVEhTI4k94yHiHnGyEUHUNmctFC5Pvikq9QZwzUsd9
goMi3fCyJGtbHijAW+ni6anVT8TKZyEXfddnD3bcbW82olEqNlnhz93hcQs9DTbY2xQ3Qm25/OQs
INcOSQkuB39EkQHg0irOzWb1PdbzqoMwod/kA8oNm/urawjMfWF8ixsqAhIaWniypRCb/SOvtY1y
r+kJmjHVFhWXBxE9/Zuz0A+Y5gztGgw0e6Rs6mCUy/Bq6ztclpDws/R8RioF8mj8m74KlOLBaArv
OR7SvISy5okkrp4H+LdUdFvdbmOm3rKOpk0Z+nxKa9wWjuRuQV/uQy4+ZlOcPbVaR9aKKqjFabOc
NVdfnv9kVCpyebkihM5SR7YKmm7EHx6xgVXNcga8wUX3+1PoDphu8SgeMNPIuSdORcPe2+JyBXva
7PfVyszR7U2SLZKeTEm1RhY6CB6KKBE/ZL/c13lKH9Pvh2LaWpfCm2jQ5w+Yzybilt8ERSksmpZc
OX1fGVA0IUJ+ULd8gWi8/6jA8ZEyQFaYICHiJh5s3n4ougm28dBLZVEcceFTc5mJNA00GjP3mpAF
nzdaP9/8bl6q4+sJmRXqem7+HvBDtdOX/Q3FOIxv7OnfDrD1x6RR5YfVo2YQt0+ml+/y58Ap/W5q
zqqXr409gA/epiPoHJ+P7B/kUzcJYoKBFwrAUBU6DzBTvHn14Hcw9TwaGSWGi93CraayOdcWLsq/
lPmtQwVwaBZsl6V1LxilbNDGeduDCUKcFzrCfIwkN07T2HS3lM0xJsTJOP/cMwBlAJo1Zrto4etf
/2OkgFf8FvMCMgvBaMSb0rxXk1ag7tErKgAtsSG5xlXMIBt9WG+6DN+nQqeebcNs40xlguwIpuk+
uwqxjTvVzZlGbj7rltktELX8ZYfogqZX2a0FPXJJaLzP9GOrbNNrP5ebbU97c/Y9VZQApDabDohm
o10UgsVcNme7dahBycXPI+9K7RK8Ca6ilxUPAp5zKVjUcIrnTFkrVs//YC1AnTrdJqNaMwNVEeMt
9+/oxhH10ec6ALWqB3gg1UOFKMjK6eNRtf/bxs5OOG48iIOkBNaXXmmYwHKEibQOP2BC+dW5NCap
WC505YiTBI3nFUe6n/yDcjcnOOu+C3zSag/2Fe++/OJXbxB/4BVTzDQyvD4U6PX+sQNzy6dTEVVK
r4VdLv7/qxFOwHYyzaOSKf4UkHZosEg3381YN5crwkDzBdqRKHZryTLdzRWdccYCsgUOFJ7fCLXJ
WWM7MiPHrFwXjNDCjWirVJ9+7UfCQANr1b5EZBbkWocWPVh0Cu/nmpqahHdL36Bha7ItSVVMPWAU
XS2qjyHXvpmnU+p24XCxuSxJ42VQs3CMPXGhLNN8L+XKRfCjS2tyIzUljcvUuWrYl6DfFq0H2nxH
YwFs/0vpTSayPyzNU84lwuMF5h7Vxj/8N/sJRWLlbAM2SaEJa4bjH0ttvxhmTBq6MYi4NZqtXhZZ
L4eC1Sgg1mObqcNMV1QMpIoHYB9/6t49ILjPLis+qd/xeJ+FubGhaeWtaV+ZNaIRd+DKa2DHFlvL
MtYsYFaYQnYcvxgSU2OYC0q2duAYZKS31ICxWzvnnTnaDTgjze/aKCzVVooSosKEjpN88JBKodSJ
dAJz8xtrTeKID61GO8kLt2suxPJQv+EfbXj+DN0/iEpkIYtBYHah1oDZlHR2vpThAGwTjMuyzl+V
akmOcYYuSEJ5ZdLw/BBNVb2rOnHlzNIZIn116L8Ba6+QqXH0uYkMSTR4RNkGsqYNMUE9SlyKwmXN
X4hjHrsGK9hId88Oe0LcSxAzLi2BFfaGEzv2hMdoCbclaQgcbbpJgpu9l55lmKwsQffbLTjCzrcT
kpiUG3xAN/+DW5+UakIsg4X2chbMERcti8c6D+OCzKLp/abaRwAbpLF/nDsEH0DqbMkxeKAEUasU
BW4Xyv45NRTy0g4h35HqtBBR2qdHbKXpYqdkjT9sy4twAOxm2RZIjIG7VtFvg3cVOxJfY9u0h6LN
FzMy5O3S4cM1G5ihvnFXkOOZlDChrT8iWYEJdO0UC/YSzsEF/IyLMgw4HN3y+UxTfIUCQhjN14gl
CsSiYgngzow9CuI8Wd+mwGCPfB5V1Gf0TUx+vzfv9qWmFxXDRY+gBvxKYoX/DzO0zbggvAUUKN1O
OYy4Nf0KcxNZuNxAOdq/lInDiyjs5uq5Y2EBW/tYLsJXrfpqA1zziqoRuuMi0P+XTTYStnq9vpbA
lxCVthpw8bbkpvJunwZ02bDFhgEejkrkEWuAFrRlA47qxauqCtw5J0CFWhu4g4kth3QMyKDl2Wlj
fEyaIckmAGGk6Q9EGTIO+6msfa8nrXBdtH7wY3kbPBC1E7YqS+JnPvjXPo8BEen3qINtTsVGz5ru
uENONWjkYyk9fGQ8FM6YKbLs2TPstiOqn4ro5U2aihSFIa7q76uaWRMsqsCXNrk/vGGgFFx0HhMi
jYo13jajzb6WbUyEpKqtbrs3rKuh/ipekFhJZt+/ApQAw2G7PBxNkaYt7gPyXyJodBFowza/WNOb
RqElhjDnoWTQFcbmI2ooxU4SKEU3wDFUExY1ZKksE1iWKTuXO23EAZ30y6e/uGIHVk4LExks5vlz
k7JQd0hxJpJsQzYqr58p11rqtKeshztX9DjLoU88VIWcLGo0gaogSuKx7qFRHtpaiB645Z5LCwNS
x/X7ihWczSO4nxa3rsLGhwxGqjrRHw6v1hZ0e3LhYnK+xsEv7vVCDng5J4oi/tIgSWejbPrHpAcX
bAem/sCz95mLibGEgmdVrPK/a1dZ863nG8w96xuEApd6cRXMOt+GOJvdivruQSXVA8y86YaPFFPY
Y8YqwyDF/OQTmL/StsOb4MkoxLaHl0F02J/n1/hehao3G0RclDhMLqDLamX6Bj8vyMpIVgLO8hc+
XsfCWC5ILYpdrm8ZwYiGS3o3bs9jMXXXfgBlIv9gpro2PCxqHCl70y8ZArb+VvFI4o9FvJr1KBL2
x/cRb/tgeWQKTcwx78TCDLhtyWczvqPP/TxDOCzN5UXgn5MVMKVpVzUouf5tdRTN42+yrMVIjoao
z/03WK0+tY+0kX6+ftXONsl38BmIRpeKQ4XzyiKiDV1XSD+w01x6kvDBsr+vSUMSVAZu02l458mv
yUyfSzFxX/qdNRF0fE6r6+wv+mTPgZeQSY6ZNCC7VcvvLMOKwqflgY8Mf4yG13aMNZciLhpHDy68
IJOFbpLogeSOsfG1VfTcmwTBhbpBnRiWY3dGhxIWR/HzD6ZkwaQbDutnEsOOhnsFuHEHDbVltJnL
mD0e9pIPf9TpIGIE0Ar97ToqgwDqweL0Mcw5QsECAvwx/d3iDeuaRMZn7qa5/EuzQuPiQDJLr4AQ
sG1UTXEe+a1JtQ4AlCwCMgS6zIMI0BClVWTISe3IYkdjNKU8AOLrP+lwHNtGRyVSpyNk22R1HVoQ
ku+dHPE0KGjpfaw9DbM6yd5XmhH3sHzobqksTUhr4YwFVG1kDbOBOmsMY0LGsYG0wD/tjbAhfWQ9
T/QDP8vRG659CEm4uxDrGabAW1FP0iF1mJeaiIeFjGzxNIcBf/C6jNqHBavfcRMFh6MkqcFBCP5N
RKTPhB0kOBj4/CtcpJjq5cyehf/3n56s81gYWgEmLhbTdRFyX6tlOoCHLh14amGYJJ8tbpmULnML
3nCS/OzlZyV9m59JbFHuwSGFVKDoKiz68g4bt9kjFHqVCpdmFgLXNKMkdw48iirLvqOojpaigVPP
mfcBG/KPWvgJrHNgdtsQXVBkdH6S9HlIzaErSwY0Vu5VICA+R5afYnFWb6elmKAw2cDYWgjCojcR
b/NDQTuDo06o5evCVK6KbP7g+fn5hfrzMxTnBz4gAoqKvfExkp/0IcHTO7rlynMJdHXwIl1cOA+w
W1UMmiE/PUsajZLo5a7KVFVpWavS79CtK3eLlvFJ9C58a0+SSejU+rk7Jt2yXo58n7J+mpS9WhGC
yXBqK/M9HqVFkeeA4yzb77aIgFOak47Pe1VfE1011qoy6uggpg+myqD7k0vrqgCoF178dBkLth+L
DWdFYq5YJNDHlWXOUJ7Cl88pJ7l/hg6Z6R42iIDWs4RIGmhinItU8fIEBrEFOd+xm9lagjazQTd7
5KKAqHvdIDJoWIF/JPt2aDqRYA1VMjSPbV9RgUn8rWhOHHIXPGyrmiplKhqadZV0sNvzj6pSOk8N
f+qRxBbeHMzJTv+Hhnv+qNc47KFMTh0FHE7OxsL8xDv0QL/kgrfVNaFWMoX1jLMdvrvnCGjQsbH5
f3RotPBi/fvjHc8jWyBa7hdYTCDFvtUl0rezJyyFLDjtUu2vI5QouuoaZg2JM+9wsh0nxHG/ff7p
dPYQJdlc/GaRcYilfoMI20jrwfJWlS48exFzdHFFFEPsqGVAZaIGsmAdZ7c/5OGOJxlKBowuJPDf
3pp3J0Ub9ZgkpKUjssMimaeoMZNVH2kZfX1o5y4RTUlySRCuj+vJn53PaMzPURn7u5n3lXpsA0o1
CLoB9PVkX4Eto3cgzT9uWjEr+HJ/StEg769Y26O56/07fXkuAWVyKnm4EaoEST0vF378eQFEgTt5
Ba+eZH/GXVDXgHeBk1LLM+EX4xpxJ8vJFgLrGiZKQJulU748sWuMUGU0A1xv+SP0ju9aEwAx1i0z
9xBNKR0kQS4YKighVStfwdlD+AH3cLH25UPT1m0EWOy7FNSa62aE3CkIfO00lGE2FZLAbY5PK4Kf
Zu+jHA6lFRb+qM3TwPiCT4LSqMsq89WogYJJ+UGcnQ15jPBuJZ5JyVbMQ8tQVoNXtiQ5WX2Pggj/
Sw36nEVeIM+O0kqHyMA7vltCZzgOYG45nD/EP+VrYx8vS4CInP1InHPs/KQlPg1YpK/KyqW+nNSc
4qEAPabT2wMZZu8NNGRYbTl4VeCeqEzCc+u61PTGTiGZ15kKARhDcfu4j39ON+tnd+0KAdc32edz
KkXiNVRHYrqYCqVhX65rSCk8naPeaKid8vTPcIvpWX+Y+goMWjXTnEWR3Lr4YIdDM6WuTDttMhaJ
/kFsow9eUuPEVfARdAygzknblP/nz7h4t+9nLo7Cqem8DKRcUbFOSj22YfjCjzC6jCzjiP86MUzO
gybaguEAndLEHpxFJ9saihzz2RIY2iVXIKfB4FnyNHMtn8vFSJdx9h9/vllsUerTg5pmaa6254mR
TpCGvkFvz8w8+cpRFMlSbfLtU4PS4frFhVAlYl1dtNelDy2hRpigVsA+k+vZfl4Wc+VJAMtjnUrC
WCjkQ02l5YGvk0dfnIVl+o6eY4eP5SmJ1LIfZKP9ddwjctqeutpKk2lqv9Zh+ZprbjBDr3cTuED6
rZH/ezEUorus6kER0UvQ90n03/p9lLLDC1oQOkmsDTeDJUkeHus9138KKmZAK1HyFH3pAMzxCn0E
1qT9WLatkdj4NvwIaY5u1Qvx4zY7a9m+kk1pMKSKjR1JLXPhWkX6sFqceFdfOco7t447CUD3gJuA
gYRRdi/ErYEc3cGMJ+ZfDCJbDWKJS53FVJJMUx3aqakc5W495tJF4i2JHMYx/uG9HxZq6Er2PSsb
J2Eo5MIIaiRfOZwNN2P+nwA0PnDqN3n71B9gcwBhxaLQE0OmOtWjkbcBXYI7QwSZ3mBpM+Mio2WA
ou37GAIDRJACut0m2IDRPPW9N6icdysWDNQqKuZoy5hL9ZD2dlESGqUUvK8womm1EYxtmrORCc8U
nrHi/zxrF9PsKPveZeS4Won0utVqPDyol+RlENSVNdYNT6DAR/TJD9z5jrmyXd/uTMahxNpTzjMo
1dKPIbXOOA7vOR1zDSr9CI7CsTPJ2jETFVcqAFVZeAyCLiryk+YzqLGOCF4VXBNccKGlD+OS++qs
UKbqRlYPXMtKUMYAeLHCc5PgDXEh0QUtfhWEOnHEUmBAJWYmy5+M4fj2dPd1tHZYNikVhj8SiyUO
TXki7bB/bCKIaC6uvOE2dhEZihf68b0DyDsC3uqakmgG7JpC/VAkaLx3ssWTZVIbpNyK9mHfjf25
D4v3rQy8rp8g545ZaYiZlT6X88k5WFfWaoksw7Ts4qpjhd/6W3tq/Ke1qsHxh9Y+Cusc/1vgQIA5
JcEKD4A4BNxEyMzq5l9FT86QpBvT2VaS4CmLsivKgS5w9LwNGOMo2ShPYQYwfUJPtmBg3p3dr6ox
rSu6HXEsOv6RWvinRnz530L3vRVsW0AQ1t4KNhA0otOhtN2Grv6zwCwc87slBI5nbJ73iSp4iY5y
bCPbvvUKiNr8FCAg9ENuh9qQ8OenC0bytEsC96TZFow0JOROmshUybigg5akeQItNhfMHPRIl/ZW
v4DnzcC+0At/rYTXufOXBcYuSsFipqCLYQ1quaqZPZKLDxqdhXZFVuRmF4CqdnV+QlJbaMl4WhvL
V4p5BK6k9WzSx2DUO0opp5l5KdcMAJai+Evpk+x+7CAGA+lhElId4pc2HbCkRTFaobCDBWmiWW0l
q+5zGMJhByqOIwvm2Z6Rg+WhXENVw5Q2s8cHPm5ugZu7+hp7kkbo4XfjaGwu16YyidvqPZl/bQxR
+lf0ldlbFNcZoCry4Xua/gbzfJ+S8/H2CdU3Ve+UZewHUhPv16BvZxaxxYZw5fq6fVhxjQUkugFg
WfjzSTnPT2rUA9c6aLVpCgTKK4z8FKsOKrB24SnNX6tgidwhRnb7ad5te8CaWyHfVkxQQkWJ3992
RSNX3hCfK3PcRCZ+5l/ZSBuyTbFcx3QHcjPiRHTnzUoLxKojg+en9sOnwMgzRybtQsBaRWf8fd3v
bBynrxpxYh4Fk6JRydfTshwrDu19159GMNnLt09HOf9UaTFqbAzT2qe4z0/Tr7Iej7VZfEatDo+a
b2YVuZ6KIfwIQ/J3cAKbqzR1lF2l1yNWwHrbcg4S7eNF4vF1D2oRnn4pJ39xwgYZc/cTcf6oWA6b
L9D4Wa29bfEL/Woqx1Vxl3ihHD7IQekCxZfovfOZ66VPUSirvI3bEydd81y5tNoxHyBu+DDQQL21
giFygFa/r0ChRv7iCR0InV4qD3nyOfWGqV/hF2nZ/VpfXZOJ/qbrTgLj6zSMSatjV1oc42fyp6oB
2aNYccJl3S0dK53Ca4DEGTMlqAk27MAO8V/1ZVxxMLhYj1y5QB2JEkLhRNoddtHR4n46NcUg0Ltb
TFU+N0mjh2R4BQGaA4Y4osZeqxJbowJXumbrI7JghH4iE74Bw5BakNzQZBOKRabgo8q2qWM52ba9
5LQ/y9rn7JIoJnuImFHxyj1XHxqcofGk7n9UeyX1AYpKVffU6tjPMXTUJllpuUUfHlHl/vSo9lnk
q7ZT+QfIKknae1WXGjU5kR9848PhUiYxiUIpma192zAYyMaM1A9MB8TDbpSQ/BZ/8boOLEmw1uwD
Fa6xZBsCRkznYvN+Su8frhB18NPC+Q3dBcrdY4fOcqkZo5fpn2C2s2y2AFof74W0NXC4fdV7ZtJE
E5KuTgoTW5zDtI9JLVYynfGXolHJN5ZPxbMxOnaGanR9YJoAaw+/I1kcOjAT9vkxAiiT8fcFwtt5
l1/N3Ey0gXDkpZUzFGP6roDXLgOhbq1nketgLbp+qdWXsrJJHUPhWh+Gqz+yBl1EPU3ooHkTvD9e
4bJNSqNElAOBV4DJcFVi43f/JmGHZfqj9paVgE/ekOi7brukrL6SIf9w6YEQVKDoiVXEIenK9Pbr
/zfbvw28960dbIHuE9NhUVQ1KagCLJrwIv6mOj9nllU68c9YmXpnOXgUvq+a8X6UURmXa35+UbKY
oxvP12mnoqHT3hPjbdhiE9qija/yVKMYkVUHkftB1ZEVbadMyyOFOpM+vw+UNxRqudnOZCT+I0L9
WIzgX0ey01UGE9uXxbv3AwmGGPV7aU7H9Oyqu4iS7umoYG5AD7dSE8GHrnSl09bhAHXaC7AV6J9U
Ejw2VZ+oYlIHCUNIP4SzQw9wsgjMJdRZi4RZqGAjjGHYM0dyXwfl2B6AXKTEG7mGTkKyfSpl5X4Y
cQI5odu2GRXlbzbf8qe/pS7INrY/LX5cCsj5lBzIBMzDSBtduRT/PoPXEJ7/1LkBbnYjeTI6jlGx
J2QPEnNsqn+oHYKryZdDWTqGYxin387jU17ZehwDabZfAxj4ExImL9awRO5Ub1+iba/ljCpU0N9a
sUe2E2Gdcnj4maB12tH9sCOzfaauk52fNq/NTF0s4W6djYwKB0V/GWWuacsdAJD7xKkirKpIqHVc
i5cYcxQZJR6vZ1hBh34hF0BXi9ypnMfxMXCsnpGX9+eaGNQbJKARnfrfjYllLC32bcasV4yUhAt/
jUXisPaFlDw5/lvzewVjTx0KIB744moOQWp3i4K8a1UZAactdj/48hqFh8dAiYC6uI99FyewyVqY
I2o8NN531pGAAZ144h3x76vsESVc4BdNNNvowhj9ZlJcCGRRENsyUsfhF/ZCkqcM4ykCGDJXqy2a
7HpyCJCD2IBEbf/AcGslIHxXAIz4JSjnlFuzqe4nMdm1w3xUFQK0IFzQIs7typh+U8xeq3iZXt+w
9PbQ0JapMkhgdCGdz4i4guykLaUTzNFdF+NGT0qU7XjdGrE23cQt32x+IevKaI7YZrYF/631O2gD
lJwAMqJ5TXeE+0GFZXCs30b1btxw290/cdjBqPcFfGVhDD4YK0MczNC1+PtvR6ey9D+3eUHAU6uw
oO5i355xKtg0eUqPH9g9IiCLlDJ8ciuJLl/Z0qjv4u7OIy/sQEbulJmk21IstP2JSS8oiuW3Dcv6
CmsurnVKJrO3ckSkXA9f1Qnn4FraXzfKfjATo6lRL+tZ5hUgGG1rjSkY7Sj47u1jIWH5uQCPt3kW
ltktddki+C2Qhz3zy7ODTYiNlQb/eN1h3NeJfJR89UKCyKUSu8QTCgM1APJRwbdVy9+ZmvupirRl
slm3l5FIc0iZOlaWl+wmlrvC+LXDPiyOuPTwxWZuDZPVqL53D/6ZQbjJAMnEX913krKtfuifuahU
to5cRTvbTruf1PcgphbO0v3qTDXucOThVKjRTSXmBAGOSky9XdS8ux9WaJCRozIRn30dfPNSCOVg
4kfPDogRYUx5RhC9WXN7EKkd2ijvGeic/UXAcIjKMxgcG4+dO9pukrD0R9reVxrU9fw2Ve7eVIlh
aYeKoNm4DgyZDN5iy7RmDTgNghPZ9q1Ji6GArACjqMyY6ZAP3A1rWMND48eHwRfcIbHp/znc6Rc2
h8sWdmIfmoXPdVr7X5wUsxioGHkinuI+kvuei3LuBVR2KJG7/GHRkLq9PHWwb4rLILsM9QZOHXB6
S0e9YKfGZF6eEKelctse/aFyPMb6ymnqnPF8umSg0AwPaY6y6gLQoOej4Iv50UZ9/qrTy8vC8M9V
y1j/GCrcE1Du1pBONUDcngMJ3nCeb631hYftMsiz4D3mnQW0qYfKt935mMfaZGi/h+obyNriRgjJ
m6nAjhpgIL1UnJBqVe/OTWjS2FzNRRCyHxTUarGI3xbIN4OOGS902L8+5emTzbtKdxyzb99hTKZP
JAN6KzSIWaX5rPy1u3UlgDNK4GKKEN5dFniqd9Yvo+KinpA4CY4Uqm1LFaJ8rpIVTt13beMYQLy1
8j4Zg5cUMmt28BZU8mkNhx57+hznRQj3InuK1p/D/CFkyya/BTETlYQ2Xl4qk5qFaKDvqHCsfNU0
9ktLOuyunD6AHzmvoqw5N17jRkPM4Nh6WuR/5ql0+vGRE81Vu2XRsa1IHpmUsxLsugii9yhKDR4t
U8ExX3yvrs8WOjGqO4ED5YPh3cX8KMbOimsgEzARrg0OapaGotcwqgabGy9Cx+WnyE92Baj+3iVX
v63aDhzHheJWdFRuG2zBe3QkZmopX8FyDOlN6WhDMgaVpepo6UZ3am1glF7Ga1Ngrb6OMi5pyjM1
QpJW8uV5Br0UvQFMOBncbdL5cR2VzAlag3sFWGvAs0urX70YP3Ycd6g51lf174Na4wG5ObIgjlLg
TG/YWOTy6IGWGkj9LCMXKfX6rXYfN8KpOTV6pnCPU1lU4kJJoaUntbmwLGl52viIzXVMP3zzuHiS
EAydbBuRE5nzTUb2YyGZWqGvDfxvLTVUAh1+QIFuFQAqnf/ZzUAmPXUsy6Euhdi2ic/yh5qekKUu
Kh6Z2RV+TYgWzuR4+ZtheGL1Y9Y+yyUJxfFbXvdkEhnQIZYzk7WT9F7psVcbPe8lzv81U9zTUFL8
l6vn4zPhbH8d0Gp52/BFdex37e5/j/HoIkvcMAIWVgPGWKrKWmKKnenY6IIDfY1V8539ComCQwsK
y/07GJH0BuMo+H2VCFU9Y83G2qy66mUGBz97w5Dlh6X9506nzTNLKDNVWvyhoo9qP2K+ndzjZ2Uz
UMgQL1AJ8QmqkfS1i9E3c1HN+DtuSPvTMM4g6iln4Zk5Afwr+OgDE2OAUKKwqiwmsQytHgTjG9LU
SitlzyzvTPAFd0Z8MZsq8ekKAWa8e5oqKsQ9ZobJLQSNk1NlDjuQ0+4JoaTgxl6mpxr1mqqeMuOk
V2HJcdIrLzLLXnp1mlQob8kseg4+gM9iSCI24z8aJB67GLXrQFEjmQLbDiUwkO/4ZOxjHkXg9XdY
tp23IaaxZCRKy1844w1jFVd4rHBGLue+/W1E5tYkAsTF2a9R3KKZzOevyB+St8hHUL6E/VIPCwZE
xCEqWcTAWwJATgf4J/0Z+efwowkuCFk/crqbbWbKhARfzbSSrhCK6nTPsMLuYNo3QC3DkZe2urh9
rhBVxDN4P0IbuEsAUKfTls+hmdA8uyTViDfZxiIducYp9XZhkb7gQt/66o3CnixKGkNHm8LGTg63
4njbZzHn0LFhPMJgSPpFoqfSNmUKqQTAvkdF49Xqwm2aZToDz9MzOIrTN/sKLZG+SQr6aPa8iS5f
FeyrkfpTymhPej6XWrmj3CReHwIaDLPtEX64Ei90LbGumBjAkT4R9CCCf9PiJfFgjrEh2NhYMN/b
my0qiovd1RhNnbFEMzHe5LVxien+9msywi5I4n6mbm58wd+cF0kjeVlAp+e2RMykN5z7mBMjv8Px
xPLs/J4ou7I7Bnvr7Al0Kxa3IJ1eRAPMBVH1fMTz3ZgHOH+2n6rEBEaqeeTIvXMbq9zh1cwrVxkb
Q4nWf+GjNENw9CZw7PAgh7R/WStsID/6R+m0joWGSFRL4vclNg3OKPN1mA2MAzhjPBDIXPXOnIRZ
Qo/ZRWuRpOlHAiOns0odQTxQRsMOVKojg9hwfkwPunZodtsO3Dml3XdpqzrIjVF/z0E9OUnAVIcs
nfkRknvPjTA7J3yerr+s1cfSupEzqVkDuiG5cMArG3bC/IOslR8Ied3PkQ/J2tOBA93A1qppKApL
mysKqG0lITxpiWUHGZB+S2RMe6zRm0U5vUE4xAPScpr+HYj59zkm8nDy68x9KfZ1nQttuubRo19F
F1nVmnsGLel8M+zNyeyHV77eWSTaFlfBZNIG4NbyXVR08u7T1xDdfeGuJJ7sx/oMP/hXnuFlgq0L
gGHxQ46gWEEd4jQK/h8M8vvod2TFizYmoq8Rrh1k4ng2+RbVrsYSfX71yvIQTY4Ihjc4VrGFt//4
RzzJgY5b6XKjSnynnBp1yo3weSWVzSwB5ldTwonTjokr67Fa6vH37rUjPC4u9I9PjKvgyaMnBu8F
79F7Gjl6Vfr9OJBftYkOMxeO+26qOH1JGZEd9t19B9E5617/SBrTMJPEJJy1H0ku5cVYlJFMf1x+
QRQZc9/JlYj9rzQEc37i+LIZsavwqnriSUAdb7JVeqSV9L4ucxSmIrF8+gg5n6gBA7Hcuk92iCeQ
8KlVWYzr0XCx9rSh3UrUCWG2s0HSqF7CSqaR+tvECsq3vrdeWGt8harHXGYNJFAZIh8GPG8WIjO9
Wq7gKGBDaCXT9hM5GwFXN8THE0JBotp6Xf4fxN3gP9ousV2jiKR0GmfBS+EDajMnU2sC4D74d5PK
D2ywlzNjIu1d/0n8JjgR3dItqMHtrfRVoa2/nNY796zMPipWKYuD5w7is1aJuQldDo6RgOlBN/cX
o8OyOLyMlXYSSF5/wpWxFLQ7tEqMEpBkcRsmTidaMmBf8IYkj/VD3vq0AKu8ek67s31PQ2OHyBnu
NCABAyTcgzRaCtNvFoi42RVVtklzuFq3lgKFsz71GfyaKeC0Dngbs9tLvUiGR7TuS6/PBx9hFzxp
qpghIcwsdsjV8kJBz2kNrs9vD6YO+LAzpNNr6MCD0E8jv84K+vgxgWR+qUt8uhYLKT+0IIInZp+e
6M0IIEEEBajWeKhH6T52OJ6VXcOzivtPGV6ioGm7F60Ji5N0Ja56Jm8YL9OoI/YJOu8Prla1fqfE
WEdwxYHyAqV0DdBadTdkYO1mj1NeHRfnM5fPlEUDZ5d4tk66gnq1LgfVhoGfrKWnwo1PGh7iOFWc
b7xdG1WhA6a+9kMn0n1WfbukDEbcQuHtRXDzdf6c5MwUcWV3sxpUdP3LfG2Hq5GaLMTKo3OCCQ17
O3ZeBtyqQK18lLPjs8Hnghy6GWBEI9vbvABb+SZyE7JlnRF8mXeMerPiTCkcp2lHvYDgcHUGaAmE
AAOcYkOJzwNHMwB1/0LI+T5iV+ZlNYxxf4X3TSQQ+IpyPj7F+IPW+WAsSQAzyD0eOJzlHemh6uck
sded6M+kVs9RI9iZv1QXbjUn5pJDsg90U3OgbtdqoMNrXBgBr/Dw1LXILaJZdTF2A6EGWT44X+5M
Y0ZhYbyViU2WKefszA9UYAtizV93MZH0Z1qREBgdP2jIzW7xTWQ4TqiIvI10ypgFWOHAv+wW3TyV
LEFrV+Rc5e6c7RlgUEoZ2ap6nUcT4egfBajog5J1yeeEbXBnQpdA0Nb34CDFLnYtKe/zPVUpJayx
HwI0XHhqT7iE7wG/MgevTxFIrwF4VzIgx+WF6l5Oe93XPYST79koog9EJFZlQe2XlcYDnyBmAHKP
pZJjsmjVznkyxM/r/Iu7zTFOUGhKYozy+Oe85oo1o8IygY+q4vLmGam4CUZbVzlRFppauVx2dQ+E
lglHzrvy2sJ21+/iaz9KF0hZlvedrpRBQnBPqKa/4LBeLH1PZvJPbXxNB4yjng4M8DgDEsOf+Jkm
l/5lTKJteT/5zIBkuEfEflSvgR/apIF+o4m0dG6wthIbX96pHN2vAZbFZE8v8vP8GLz8u5Hw+LM8
dDfGsuVRjyoWSts0chwfUVM8Zkyd1fYIpi20VfP/lWbU5ALC2WjktOInnnBlpUh61jOBCqhnTCW5
aCkpCrgm9rTL3zR9v4boaHwEjH1Aw1l+bZ1gRfNb85M6TKd0UaV8v5fKG/hsPFpKOUUH2P6t+HIw
eUSZ8R7F+e3D5Uro/+Yi/VyoFKk/DYnj9d9a0PvzVbvYuqprUDMTqchDhh4v3AP4gPWsCP5LDqLH
ie+jTWeVKeetlynaE6LSGYQN+uAtKPXx46UD2IX6Wtg/BAbsy2eAIi+edmJGL6jPaFUV+7QXDSeo
RbLhFjuyn53tl+lIIZkFW+93PTvSrW5zpIDEW/j0F64aqE7llFlRJmZZiI0GKR1d6Qy/tp9lZB+x
l9/5WXTvCYE8M2RKy+lGoMgU//X4maG3WTBZZwaYOWpM7feLz06B58oZvnBuLbyIxABAfF4eLGNs
0nt0R5/RtEf2tcaADqCMVrmahHtqx7oNGINLo90UGCAv6IG3Q1grkW4FmShaxY3p8tWTXI/3ouik
y4Q6ism0Wm2UvBp+p/bcSV8R7Q1s/0mIPPBe5tGRgp+LBXEONj6wmP1Rv5I3tSe+zsekQlBfeu6n
CYhwKKRK5QMOhAnJmpgdUwdTjmuEEwXxbnR5Z+dyf5az2p/CJ0AdWIGB5Tsqna1uiOQmCcyKfq0X
SPXSdWnG6MK3XAY5D0PCXvbzF8vDP73FwcgTvQeD/v+6gGmcrKFjifV7NfIEFLXEG1/yyBmPF1/T
KyG5Mq3kH8RNLgnmaROwQWCUs6DAJHvPqAfWzs7IXugd6M1U8eQNIilFMfxmQ0z0M3IAbZQe84ap
ysznNBuKj/inomR9FQKhCaglNhoW/KkTSOFUbB63N7EbfoLdja8/SdakdWifrQBGDPmNrVYQMcLA
tAICRbfJ6KwLW8IJ1NhGGvb8U2EyP1YpHBzEb7eXWf3CQASrWWMknXESSv5o1h89zPaUWtBBEysD
43XZcGL+3D8+3pskradXCgm0n+8Q2vjCBZrbQmg/NlqvVP4nBgEvH/uEmvDz4E9ReI148jdVhNyb
K1F4emePs1d3RI9UZ1dY2zv0QlioOZYz0qiGe4CLLxeqRv8pnMK35cKledySlelppnwPh1MJdUZ7
tRnOwsCHDClyblq6OHW6mQlPY0FfhVLiPFLgY/NY4UQxa6kEVkuhpNZOH5oBW5KA2OdcoDa4BYOZ
7vwV6hzYSNKqdUS0W1/7XDqMwIF9mpzzB4H7A2vqVJ/Kficpps7rSD+7KpRJbzASkinBZibYtqIe
HUQyGFUeIXgimTp85o2zFGG5s48TTBQ4TJgqbl1h+xMahzWB/md7bvyRvJhOZL6v91YIn07VOI/Q
WJq6fy7ej2QFLrntCtSmtdMET2NzDeWB4NGkAZ3A2exNgn1/vVSZw8ftA16cod1Mb/zgHahtkYqG
ElHu47rp8zlRPCPot5FkoNg4lyzfVGwKY4wdrz5a7Hu/GkH6JVeZSnx164l1qxRWyMt1CSVhJ+W/
sLLexQqATTgI+ZI5W3+WCdtKCi77nHGLzoHA0kYj94AUKmjmlkleUPmr57tWkEobjeoZ6MfVYfzy
/t/D6AVEbh5vnMjwK4rdhZfHUYnn6jKe830mALcLQWmIiqqh6z5kXtVZW4KW7n7zI2o4q/5kGNPu
uapliyS06aw8cpqBgEa9Uf8JI1idxkhvdoY8FcVKZUEHz7K6WxB/xqeAG11ZelGB3zpinmt/oYNI
mONL2TgVNMQiDZZTSYq0itsQtxT8C57p25pYs6FKmw9B1Dls+7LP3xepveYLBpAxl3XaJY3UwMh7
swq4HKiH/UBIRPodvcoaRblyP8C3MN5G79OVXHYVvcIY/kI71pizpTOQpX17XrTRrQMXqsJYhJ4F
aVhIiJ2WOCskhgSdIfQJpIU5ywINmaKZMjv54wQQsh0AM/+us0R9FDVF3DUk7J6UarwiYgMvSk/Z
7FGVwpPl7+XNkOL6va1e2FjgYYrrJilf826XuxjLXZJdepJmdvg6FgbuclerQ8XFTlmKfn1gvjCI
pqi9jwD5GSYqoQTvwam0YrWZwdzwzJ1J1u5+WujRJ996MN/WdRhGTQrs7KilmcaBhjZp3I3xSjRk
kQHpzUYbZ7c/EerMcPdwsIRGhSNzeb25JuJkq7TdCWeqshPhpZj5hcH3SE1BaRom+HfwNimPwfSX
grqqqG9JEnA+g9wEu+OZMMqfX9usOhvxbrkejEDpvBXM0+Qa0biS+XMn6KJWpP3rDacyzetw2JTE
qPNMO3lKk5uXQ6EkVVPmnO4atvEe3T1ePO1Tk1ZTi410RrHtudjRrx8wiUXg+fAgsPXI630n/nbO
Tie5mwz/aauq6x5HSGsZAfWjN5VlQ6+dsHCM96MH2z9tqEh73/JbV9fkAue1Ug8ANXrOx31/pc6+
iq5JYOQvMGWf4j8ffoR1XhT01R7+rQrz7vjqZ3Wo4TVjh7gPe/2h5ylhOxpWrpLUWODLl5ZZnBtd
zmnWwRmizwZMFtK8vQJ+7+K3GFVIyv2FakjUE4s4tN5VUm3RPMJDsSU3r4ejMJUydfegOrUyI/KM
MsAbU2aREHijyRzBc5AGlMEZkoZknPGUr5LsmX1fTy9J3I1zZNxv9R+Y8l+jXGovhkRdhIIWCLev
iCciWEsVCmmXRYPpqtEN5VWtMt8Zmyafm8L30pFiqRveP8OA5ABgWI6l0crfPWcUzC7Cir4nX9ZG
ODb1aZoiaQLD2sSC1ocJDNOrEnMz03KKU4tDU1QX8+BU2yHs8ZMdCHdGOff9gEZBhMKj4YqGU22x
/EBZjg+d1jBAneOKJhOicHvS5n2rNzXzErZcqtLk6Go5EWrsxp8FcYxpyHPkUOUN2Xb8Sg1QY1D5
Y4lrNK1ieGqY3pLT8FSjawsS5M2AR3zncs6iGc8UgnauD8drI4rR3z4zYNTubEYv35Y0as76Z7Om
sMvQZtq+hAwmF57BQaS+G2Fquy8aymXUGqoybwQYobxxgUx0+HWZIHB+8nqn5x6rCtDnsC3c6Anq
n/ABk7rwdU/x7CB3jvXxeYI9Y1Qacg3FlyJ0B7Y1X6LFnH8N1g0XHfr4L0AVXX9Nq2r+A08oehR8
WkVTJ+98Nt5tPQ/cUm1/IVDukg7npyp417UxZ7xrGagEjg9vNe0YqHWtN45FJoBVXgyrmfoFY2Yp
hyvHJV1C4/OXwMwB4CGw8F3lgaVZWXNNzyhJyfJbmaYqf8BktqKOOSN8VlYWf9uuzloZWw2KoLKP
jKkle9PdQaA1lXSNhbOirYysY3zQlYfawxthCA7f6UL0hseteOC/D4ipHSzd+v+mItmVydltH4KJ
4a2B0BWs1zmc/EtU+t8UpOGs9tJJkqMpWgAtoz3IdjsxX89Q0JOpfWeJV60AKUbhcDnZWEdDzRnR
LoWNszsCRLYgGJc/11LLj8FgDP/YV9LLLyQu+UrhhmpZDzVv1b5vi6tmZXbwmtJ/Bhv7V3r0u3z8
NNvYXJOWVpxquNInzjAiPnepe6PrEPIEOeGQ3Q9P9RuUQ0R/2Bw3mAYB1GAQsiNxZrELtgIaDwFu
Vf8EiQDGnXBK4K/iqS/tfK9iiI6XY/REZtpnjKs8rbY1oVc57xx5H7w+hK/4cI9qtv4SerYkzEbh
/u0fE3LTZ4vPZH5E6KzyNKMwsVUpXVGlKAk3lXLGUFOA+P9XSIF4tkGoV6HIzuyP/GOViOjZqAz2
Jll2juhGNav0B6FwRl6RxBriauUvll+IcdQ0pcj+myEjOsfk2iYYdx6tqT+fiiJdyyX5a9MUX/e/
nnyOPwGjEwmmhZUjwzY4OinXJQQBE0KUSGDHHuUMgmt+f6AZwxQ02e1URVnYk4S+8llfgeHzIQL3
a7CcIZBw6ULsXFoTcs2fPuJ8vEcp20LLqv535cRwNV8G/A14TkE8pdSRDzGguMPwPa/ntmTGL6SR
C7eT27hT1xkM4bicipdD1BJ6p1V/f8XrShmMghjZqLY03F5ZEpDjsawbhVZSMb2R0OvtQ+vuqssB
bpfMcETcXQ0PjWDoIcGIS3szTWCqvIOfIff3JoN6m8WEzM82vKH2LCWwtyvsSJScK99OzopBm2DQ
xlR9Z49xAYPhFiHJzSxIGRzqto3h7v7co+2wdtpDZxBSTWaHEASOQXwz6gIP11myDZyyZYQFYdtt
X+J6CiOww9Us/i40nQhjBANo/AmdkjGBtFcKHyBDPMq9IE24iOxopFDYaIsuXtYEdYeB3tvE7r7d
1MhaePqQXTzDmse55wcBzAhALGaZN9c7MWUmuLXEWEK0r3LOVOVuJWZ8RV+725gnWjWS09B2Cxei
mf+taUjLVBEANRwkR4la7xMbzMhqEcJ2xbfnoz28O5JK1vPsqSjKcTh/RV42Oh/GQL0ptwpJQWTe
0kMHftoNk8Oesb736XdCCZ5xrHBXY2vpYBUCeFHe0TxnRUqqUA1rzgNU28Mc+tV4csEcc1B5ssH2
830JTl4mV2IM7kNsIPJdwU7o9mjeQRBrAMto/0W9tsycaQs4YZCkyag3M/TK4oMY7BBKybkx6V10
XP8IkVTPhpcYWgSpFZkXgw7zgs9M+lMT/Sl9pLUF3KxfyN3do80MXQHAZBxPWP1ccKfncdmBHqRN
ewuvorSKeViEQ9d/B1erfrt1oCohDUVAccJRbfOr27ocBl4hJ9UzXfBVH55s9uFehMzBaBKSFFR+
U2MR700G/m98dFWXqi5iMmVQXPzUpYgJ/FuGhAZDNcKQMfcC7ZoONpL7kRxfn7fdctzZaJt+KPQX
/0jIISd2EPetBgqP5NSxioHzhnkk25HfHWj1lH/pnT3URl7fDSrrKPIi+UELQIbr1C8Afl+3Ju8W
bVpv67unTriKr0zNls/GikB6ka9fHRlL1EGL3RRP7B1dh92xE7gmZFavdJmFdTyA1N7EKNH5UHoR
O4lXC87DNVZSLpys8apUOxQM2NV6pxI/55VmfDeb2yQZT9J4FL9Qp2Js9WKRKvm7TLhw4F5YTTC1
3JyfMV3/hpK0obWu5UYwKGKijBVMozbTe5sAH2qsTLLlreDCAFE4a1Odhm57mC+XxSJ4uAGAq0MN
Ybanv7v9dkw3K2kF2iBF84G81D/K87jGNw7iWJ0HzbCcYVITbceXdLfGGkAgZE461jAIv2goNzut
16Ksw1u+sIddObGQ/ubYT0fx+Xv3EpjWD+IQ0DWt377nIMajc0gUer13pRneMcIgHYsh49XdyEvE
eWebBF2VXRU/tmn/eiHI/W/XnYhJkPCRp/ymmYgf0lluZRKEqPDNSf2RhaLHks/nL65dGoWXHGxL
FSHr3KUw/XwCJ4hsQ6FpaNmcd/EGBndMHhga8IrS0Tslxcjo389YOlsyzKvgdWEUe5twhK5wNlaq
rltiye7gKevOxqAEvxo+FYdTCD9RR76BS51fwG1l7RNiyxn7RL1vlZgNbNNE9xQ2efTazVN3nuy8
83BpJurHNMp1PtlVo/amPmSLAkXPxvSHP44HOvogkmRnU0K6KdgKjEmUCPwtHu6tysEuLErDkZok
17oaFGQUkhztVLarEQRVWJ089vbDOWiS9dYyr/wkiXz2A8b9Pw3hCZfltw9zy7eFBauxF1rMkMnM
XYE5OSIg8zb7+ibExotND2TbnX2J26NwTBQaBXSl8YfEEudVr/DyFfISGCJD4XV1mdhfXLbv+Sdn
Qz39tT9X3hllZCq7buf2G5tAWcH+MaqOf4mlBzhx3Bdjq+s1Ua1zl5MI1A6U5LdZuvgWwzcgLver
UdLkja5JPvU+PDzdFpPHW/Xs8wFBhDlDMRyVCv6pWf70V1heNsKN0D6VY71d+M06FByuGrsn+tUl
NZds3j0OcN1iAM0MWp+kSr1cy81bjEmHAiicH/qdTF/535UqQhkrrcGV0/nUAHqKGK4PddtU1toP
jfH532FlxXwLKqiVKr9MjXLJ/VUDNeFaG/CfoO7F9lOGGOrk3FDJxrMVFGSuaJ6gVeZqxgOQV/c/
EgGhgqd2RPvZdS4pMIe5X2L9Flj1GLVflN/6LbOOySHZvYxn8f/rmDIWR/FAYD+NYg3LNRh7jg7E
WaYLOC53syCBpBc5BGMNmAIOckxtmulCw2qZ5JNyQsOhdoEiW+tMmfRjnNQoqHj7qCdIQv4D51M+
8sh1NC6wQ9tZwOGi8cNphMe5TeY6F+olF9hKwj9LGezQs09xw6Oe5pLTKFjddNyFsu1+PMRoTJ5H
47OSs4cZBMNUpaflFgI/k63KmrnwgRa/7B+vylFV26aw69aTWjlAkCAKnaeuU+GTAuKQKGkSUuF4
Zp2EjfTiludS/Tyi6VG++kUke1nB2GWrlXfOyReLMscONhZiZaT7Jd1qpRTJ59roDvDdFZR6LJ3B
q+3aohGDSAy5F7tlb6m40mAxU6uixwLodID61trpCs/HXJswpGtIuMMu3uxdyX5qY8EUc9WugQrH
Sywn8A1vySq+Kqp6J8ccNeQvkBi9hlVHr7D8Sx4d7tzf0P+dclSudmTSejVodTZPcebEt2AybJdk
J4k56THEtYXh3Jmu9Nsn+APLY0f0dvchTUhr9/cKd9ZzUM6CI/rpqnZp8HdbqtmljXEWpUgkyRNz
TmCD7epymTw8vSmDJohf+cNt6qVJ9FePH17qk9z/7cmrkelQuhi5UK8MHFJ1mvYQAsXJlAc5CC3Z
GrQjjCoF+QKVXXSIcLhqqQpijmIi+7ylBmhfK+I8zoZmDdcXD19ODt+HO6KXCpFMSkMHquqqkD02
KeyvL9+Ze3q10ul5s5d8fFre/sCHMy77mjtky7+qVuMYZwlf/su/uI+ub6YZC42rxzeZxs6/dfHq
DsFI08vwt6C/kqGeojZ8Y4Tct8dmZ9qkmNOOqD3EWjaby5ZJOiTx4ioPtcYs/JZ9+e18qCpPuvOp
Pn+/kxpc/63UgsNqkLVU0B/2x6ICDIPfRPEFeQKr9LX3gDf6BhEDZ89NPHowhurn4NTgpxzn/Lx2
UDn1cDxSZDDvPwK11rMbvW0NZxdBTe16v4GcOPh1jajaABm4Wgw/38cJU0E2rrkf0W5RlZTnFoDG
4hzyaYkaFX4MORDhgNY/eOZNP7UOMSTD6KsIry+9RAHQsaGPoXHaEy70foYd4Qfd90tZX3Vd4Ky9
IFkh9PkAsYIP4JXakqtDwVhx4lcJMJOpiwzJJB96qb+vyqkjAIxs3ad3nm6LSIOGGvBkYA7vy9kX
T9m98s399vyXCCY69cPRdsxkav5sAGdllW76UkKyZlJChe4o3ZQuK/kgjuf4E+XDxGo4tcwdgFrg
fD2P8LCJtm1eTH00pdkopPS2dSgsiMcm+Fj2cHNz5GG86pst3pZtt2PI46Ac/Z8gA7okU4wsRnhx
NR0LjBz9H4/A9KLRowCndlij6BoPcuO0+VisWQfjQZKYxfHsm2ZC0UdVM1uRMQ7+ueNeIXP/NcP4
QELfqrEfQ8sFeBb8rC9/6fMGKb0xvIBl0FWeuYHtQgIGQsVgRUiPIFGwc54z9034553bCymlNQUU
8qPbzX+83Dd4+/Fy7Bd0Xam5oE6OykrD9Z60oLK6brDylfIvmFGjnkgqLGwT/fz5PbXPCrBi0wSj
x0Bh+w4DGBAwJWSGGa9E11Z26nkkw39PK1Lfb5gNctUXPVKN2/0QdthtPNmaIHAwo15YKlTg6eLk
J20y11tpngZrWMovBEXuWni/DI7xFZ5FtGaI7WvSuyOnbVuo6YU9s9U9yt3c0xm8qIb2lG3ThYiK
4DyOs4vyFr91vLZj0lXtKVWBXBAOq/73ewVHNRFXW+O7wKIKb/DVEGXt3grkqePJ2WFhUlsgU3Uq
h4jWgxll2Q7Lq7oGR8OSVSn1kGcntYh4MU5B6zz+9Po5fgEbj/rEGhKFfrsBtxoaboiTETf8gmAV
/SWq7hVQqTaSGAkMTXKAnc/qnrjNsu887XyDQ88lDsBZH8UMiE4Kz3molZijiWywCQKwFDwNQeLo
Nj7j3m8gsBGFE583B7UDYe3UUGV2zHsroFQ0wdwSsJ99S/tKpi3XXPVXT5vpUsFxWhRet9cnpeXb
NisaNeBSh+hxlBJXzUOmdpOmeqR90W0UxQvtAHO1ArCPbln2/J0I0CVIXrsnMMBIBx0qlyicslbT
oChKjjhZUyMK4YOTEr+BUMAV6//Y6fq9X8yLEYhX+BXLjOwnTf4/RMohtouTSEb9YVbcknpLxSVc
Lx97RLMx8p419hW/SScPJj/Xsh90HbhIb1E2jDj8oUtGARLTek+gr1+J3ujlpNmFFEPFBCHpnnfY
x4+jEgJGJMtU3O1TmKPR4wl13uF3zKbVwZciPAa+zoeCSfCzPzu7E+Pe+z4RpJ8abN7WnmWnxXN5
RallmHy0rTzJo46Oh9xpHg4IczV0EDzuSuUEzGApFjX5CFqxUfzfSvHgUw7eF+UEiz5GcXD6YRhV
BDPHYORYMGTj8uDk2bzUQffpe5PPovloyWtSTyCyVYHmAyBMQ+lxeNLTeXFNgS6ypFLNkpauEHI0
ane61EckvL/wxN95B+fRaaY2CixnU1xbcH/Zg1b5N3EpV/mhS+uwOcFxARFXHYqhB8YNMZg/HGUN
LePz9qnE1+nABSum+UEhcAqTOWnpZLYn5yNOEOHvoiVssWTMGeqT672EMtXN6cq+JXIOty6530yr
n4k+j9SVPq+A+eUJ0cuNwQqgV/DARNZZXD32zS6zB7mVh9LoHCWJhVOtcRi4F225Fusya5JVdUqS
HtGopMjqqOXiBBVL85eM+TGiTGpmZPF+SnR6JRofNdzCWR3Vcrfy0MJ3377dEDU0kHl5/VCTVZL5
MzG3hfW7OhLKtzqlKFyal99RFWwyTNIdhDwgCridZBGlc+4Nl+GBqR5pJQASejojfMdmFyOLG/ni
Yithmzyof5Kn7bRSzb6erNx2F5mYUBILRxZ5AiRdaXcGRKy95tkEcnFX0vNzRs+rm+QEGJ26Lkx4
PUAOZOxdiFVwwZjHgsyXOY8LFJ4XolM/lnxmWn2K3Rxo4jNRddvG9D7XzuXfM3my/4/Kw51r1/I1
vQBGkumXlQLxOpNlt4Ugcdn/U5273ozPgL0q7y66Iw/WBHcNXZvh/SJ4mxJFjk9VrRJ5+MAmPuK4
iOESpHgiOTmfj/5SQUTaD/3oXpCfhWty8E/Vx6YjepRwGdZoYzVTI48qYqZzVAIG4VhIKkpsakcV
ImJi0/AEDuICOtmgBXtqlOf2Qh9/15bvIRSQM0UvSO0nP279S0CNyRBd8ilxMazyC50ugxqNFoAB
YvUj1VmZC5PM0Qvkdu/4x+/Rb4B+9glB5OT8Wl2i3hGV/g4uLShpSO4Ab9uVOlTz4LnuKbUV0gvd
hahYO1SMzsZEpBR/UmHWA4nIv/R7OlZl1KnybgUwr82R502qIv/JTxG86hFtY2bCVnVMmApAmQnc
6ZD5/uka7EM3L2X4O+HxHGVYncd3g+dmmjhcM/Vek0J9uusYdHQV6PKi9Uu7LJWVBKu96+3PK6/Y
VLJexjfD/UcISjDGUIvuLdre3uRuYxZ92lg2Ej9LGRJyfVzWNrhUkofTZ4sq3DMlrE3qrYezG2OY
JPFYiNJq0fo33ITBRX+Wqi0u9chzThXdCLbaLDLLgOHHHy4QUpzmsGkFCu3ky6qXGmSVf/vCn4Zj
PBT/QKOW7zdudztcNI71ymYqwXzPTbwaAp6SfMZC8c5FdSLV4cv3FGdADC9ZT6L+nz1mIwxGOs4T
qiq7M+fBv9IF5Jj001ly2BXEVJ2jTZ2somx4WIfwKCKakuOR2TVvg8Dyc1xTqSoBN7jy0JpzcSwH
q+97YriY2h8MhTs102er5MWhWJ7RFQ9ycKRJpqTcpTRaHN7l6VBqYkleSDBhBxmnO1tqIZ0YJb0r
7JXdmQGdqCAbeCPulnqXzmflv7NDLtNTkUhFohTCk+mipgt0ezMgEiJww/lJypDoEKt0dkN/9Dtt
FBid1YMngUZBa4qJU1WiR1xi3WCwy/7U1u2K1Acjb6A390gY6SHr+CJAma+3HNzam07zYeOd85vC
lnhhmHnW2YUVDHWmx0SwZjwuZVPtDyPvCRbHAP6E92VSg1rz/jC6if9npkF2oupa7Uh6HdMVxPs8
d/RwJn0tk9lxIw0xByZ59t23ylFcTuT+CaH5AK5cfBIenc3u1iAwFv91p44mDs/6SZhmPwpYRwIj
MCgLWaYNrwnfZ5t/tbRmH5iJ4DaHM+SpOh560+2sBEQAIDIL0GZrd54AR9/DKBbx+NnQR0e8xAB7
VkmjfF26HmKLWyyyHRxkgOQSE9XDTS9aIiRSIjEf80i5EDMYyzQuLiERCs7RuzLetHpI+oocP+Eh
gv9bIHHtUTO4VwhM39nCdSAhqKLwYV5FTe7meHeoeRCMPuKT9MgH0VBKY+SiLQWbwU0r7ntm8fr+
da29EGnPrbsS6uiTvo15cQ+mh339yYx0GjU0CSVx720NzIEjdOmVkEHVQanavI1BGbtNTfs4kxgX
W8vV33jz0IylXJRi1JEm+FphZAiWObFGBsdJ8BSr3jfcqlnxlw1szIKh9OMPq33d6QDNF3wbn8uB
3+oklDogE/Cmo73wO8y7nrtclFc5f1dUnnCzsCIETQCQLlZH1H0QrvP2rQ5w5DGasmHzNHh+B1kV
t6BfI3FNw6dn1CTdc23Ixj1wdKsm6EAZ8yl2zOIUCM2E8QvccqZRcwJTXg/0yaOQXf3pmpe1t1SM
5bX+FREx+RYw9nErjVt86LE42sNOlTnVjNygb0PCVItlFc+IyGZwDVF+bCXWReLZVzsH39Lz7KM1
5G3J85y8SO0Q/N2O5gcHRoOCx9gOzZW9YD+qiEYv3s5n2If/wIJTudDqXPisI7QA1fsAJaZu9epv
w2c4B8j4fmIiKG5/+RNbpsoFG9MF0Ujyqd4FSkr2FRP8Mn7HvYyLoeua6PWZq0cRlZ1iiNq0lftc
QlRrZ2g3/agRAprKiUluelxlHITNxs2DIIMup/v7+99zK/BdlsgkzzexC05/TyF7zQft1A2TMz5W
DtiPLFeNy6qm7utLR6BIaf4hNow4dT+OWn+UlmI1LjjZb1zyM2/Rk51zcVkjz7z1762EcjeZ5jUu
5mhDDliNXk/AFPLue3JllRb3rC82ECXwqPA+03QAN0M8MdK6W8zem0jvBbCffN7YvKOIXthOFqCg
KV2FezEJAgLs2gfYnifAyM+Zjx+ZqQIeyGm30x9Ty8erSKkGymxl5wzxY82i/7pp5P5J21Q/1ldn
nsIAbv+oNzEHxx31J0rBsINYqCJLlQdq2KLNbuRF/QEO8Vo0CedrGYkd7V16yJZVeroYnG1djgk1
WvAZ7RDfqwfkJisBQqZoeExTiZmwgUOowwFSLjo0oGHtncM2AVbsnNLfQBeDJa+gNrgakRkG38Ig
6ju5FWyeCXSlWpYEtvzDnbvd329SRIh3yWyKSFaryc1a6eINcAFwkkOXqLfD1AZDvFCRitpsR8Xh
uPhmD4c3/G7dKWVzt00/VRHmI/uiWrsV0Qliu7eccp8P5gcfAZaGkRpe9wMY+1EXrX8OTJ1aSi45
xYeEGTo0WMw1hjcPBZ6bj+KXnNZf4sfsYluBmSy8mCygpBIUvl7MLTLoHYOlz9KaeIHP/bdRxBJL
E8vbEz/fWqb29b8lzurKDKknbSrQaBwKgbs+StKo9TmHT5YTgWlOzXa0OGs6bOekvIwe7qsliRpB
1H2Z/TZU2xhJqBq2z8wS4SvcPY/Z6qMR++NIT3XcblSeiDBwOO513SyaOzcuebuJjIAsCd6Qak07
q0NdD7dKE47r+ooyOLxXfP5rIkCuGvslnTPG8pB1bEYFwsZHiMSsXIPUdSnyihncuOpR5yKAlpyW
/O/7+jcAfr5QH47UC/nzLe86wRfkYm/oW4UXZmdV7RN3D8LEfMmfltJtSNQpOEWtPDjJ13E2LQ6r
11P/GXm/x/QJbOhH+dpdbTDasd9RcLDAVQp3lcvQNgbR1BLKIv9vN734GsI5CdxZRlsj/4V40nGc
QS3WzePYKM7beYh1029xNErITBP+VomAmwbXUjPe14vWkR67tdrkUpAayGMXQh7rVBBoFxGvsOsb
XMEWLExxw0rfBJDTVFB+Ks+cRrAg9Vn4GEQ1DZSERKiusTSUiUFpQUpnkK9GEtQAVcEQWVQBYFjW
uXj0pcO9RH7oti8Vo+2JxtfnDhmOGhgYF52bSQ1bOBYe2qWfgDFQ4wXGIxoSqc5zTYHX9VMu3Zd5
395gAKVUfuQ9XT78DY2w3bs42ShiwDyNrBCUfhnWfQXsujJA8AuCIvpayXM3B5o1RwrmlO5+8atm
QToDGJlEGE3aIphyH21LkVxW6u60iW12Iy+4lBQv9nu5FBdKFU3GelLmzIjNEm81/lUR/nU5+ndg
EWpMnzzfeqUkbq7XqSaUMgMuV+MtXndmHwEPrSMhH8FcdxTAKdb3eFaEEBZGJ5Q1Emh9117O6TyR
DM7Rlt3nmkbRsx/MtAiFb8SiXuxw6uHbnr7fUEBi1xJ60jfvZjQ2gFnxuHR+gXO7WXgqsu3YlKBe
v2Gq1P0h5BvEvJxarV1zeAPIPChTeGqgjMWVze2bCObeq0st6k73xBsqQMem+6vshnqcW4R1JXwm
5wYUygj6DK367AFxOMjMsnPegbqZJtdOjB7ysQR+m/hDbMT+BI0gunN1IGeyBEb3baPBrkGVvs9f
YFE8YxijSmj4KslUdAEyLSmNOQNFhShhIFP7kgNFECVc42BCz1Nh4NWB4QBboPLIINwaQTEnzyt/
+zZQ7Py/1wfuSKF4+hxoVzgdmaURe7/3zYx7odeTac1YZcZsEX3LALqXxJmm8rmfEA3R417g5EZm
eZC6Lfb8bnhrEW2hWE3LDwxxWpQh2CAY5CSBcNbA98qz5Fq1mOgqMm3Oo1XsScsR7slexXJLWukl
31J0NvAxXs+V3ngJVs3NqXb21WI/N68VCiYTs6ugdKh7F08C5KErkeLB8g0cDiVSEO04TPkkyuvs
Fus4Wp5jZ1UQ2Xp7JutjOCIB21TN6/qzciWsnH2hgCoNTqUx7oELRiFT+RvjaSw9dMWFHClA1Oe+
dmAGg+YroZm04NmTwexXlOtYzzMZCRTUGeqUleuEjRmoaitEVKIgQqzub58KbKSKDPZBqEkWIVZp
RgvpMZJtR/DGNfnF1W5mKA78JmptD5ycmFcXVyId0c2DzUwULmLCWTwur6DyZyRYKfQ076zVJZCu
FAeLDNXKI78IO9T2/2e/4D3GTkKI4WPRwHWXgbY5Fnq62kXEOvKSBEgoOOlMshQAqaCWy9cvrgbY
nsaEDHw9kwyJYrPzupaoendchh3sgXLdH1DgMIq/abSmzsuFEeFuHxxwU9OeCgf9wZGbzu63i+6J
pYneRTMSMjEe1ch866Bee3PUYtth453iO2qN8KFW+7/lVWGw/kkfPX+7/b8S8/Abf606aIgJKZyY
UVt3zAo2ADS4Hsj29in6GJKG6PY05zJ/GaiJnzxNGqsntQ57ckJozDGMWRbZBMh4YvxeCsHR1fw+
vN8rrv0Dcw9zCwvUsFaNxkzdqEprQz/mxeh/DtPdylJNLQ4QJVVOEmOmqq5vz7ycx8vj3eqatwBF
TNkm8p/un7e/pS6aRerl7uD09Y2mF9xLb1lErf+Asv5hjQ0fC8WtFTg8eM/zkJJphIRVqcpX4pd8
7qPEhIJ8ntiBf6u95RdEIEOXgDqQ3Ul7AIYRyA3dziL8LO5/HlMlYXXy3FOT0aZX7a82FR3Yf/yB
gkQbmxB9YtCtsN8Hnrydl2ebLx++Z5xUhzhhDAWSqVDJFC7isSeMpILjwgeDrIv5MaRkVqEtaMdu
FNEWoLhnOmcfXGWVtEX6eHV/+zXnR6/f1FVUAqgAAD7cdtkh6mZG+KaZdZ4ptdQ2tpc2sKgP9B7n
ca67QioH9g0LX5KF/qyMjsIIApKF1eEYQWy8RBpYy5RHqwi5cur73LSPxzHYR5ya+z7tmvN9CcYG
EfeWul0rcdDDO5vZ0WqwQYbEZSnN/Xos1+S4CQGvO1P+t/UkYBuVuOHmHTCqvWmMqlaT/wnr4EwZ
V6U5tRYfeGKSkdVWKyqCO2PJh27xGWX9gxwFeyqMfMSoCbY8qwWlbkEGm0Fufu2OdTuwKnM0FkfD
S+RXGhRt95QTLTYYg/H3TneqOCmvCDGExXpoL0CfbFrxpqO4nEaVTgTTbEsDZIpDfjysU8qtMyfo
Ih200uupAZSNR2gh+gb33wZTq3ASXpGzPnOR/NViSLQZ6ha+qiar0M3knJMldlReJ8cReT1ZaAnZ
lexdceNvnc91QJZUIIrohyeaqymUs0HrNXUBsNxBxZysQar+cYbcjzhp7jyqHzFuEtdK3tthWPex
iooZT4CiNxxNxBRLvgeRqcpk9Rr2I2I2Tv7SnWK48mpAYzjumH8Xv/n2wll1mG9XR96pPooCJZt4
HsyTQlefP5liJyqGCzHGHAytx+FW8hIfnc9+07iwftbqW00Cm5BDS6H3OJlCkfEEeTQy6+hKanVc
Z8bxoyAe52MGxiARkOB5LxQb3btgMOEYQN//cXgLU+fnCtSlrW0rainYlW+7a2Jk4fQ3wC2ps3I8
pAJbkxsxIBWgaa6btEqJiG8YXKVm/xci48dBeItArbQJt2A3iVUUaqnBeX1MlEwtZb9tpW3X55iJ
aS1apNS2iPEk+TovzvmJRGJnQwkHPVRXoVEsE18ljbTNg7QTTSQ95+3DAbrdMBHOL5e6vwmZ/3gC
9IS0PL6Hf6v7RZQmjgBb9PhXeU4PPVSemf5WXXekhvyQL1nL7lzsBvpLcZ61MvQmDV6a+bFE+NLa
pVtU9AeBTSQjierbfiV62UoYUBOI1Uoy7QAb/CEc6p2JOreLNQGbqGfrm+K6H32smJKrybTb1ZMq
znim8w+hrg87xn70ZGv9fWsXVBQJiPgTl13A4GW3jgNQb13meTTzYJ4OHMToc9R05qy78XD22Yg3
6ob2d6vW8jFDxTYcBnaZCThZQKCVD9OiZBkqzuYqZnCkEgUpkaQiCSZhFqCRQCV0XALrBF1dmCl1
KZDcbh6FvYl2mbFTzUHfICevsciB99VRJUI0szLK6pZpj1aEwNGXBg8bB+gPx0t7Sn8OD+uzV3XB
B6hsDb/AwLE+H3l0B7VW1qdmFFhsuUyYYGSeZsGSJxpLFsxmG2dOK5osNn+oq6Qn+VQjmV+6lEUN
PJVpOxjtZWZB9JLd3QvDewfby2SaFEibz1IalRfKu6YF7IoWM3J9o8GeFnL8oDI8haVq+1wNTPK4
XFrpJSm/pux2Kbr4ktsoWlsRiv7OeBllxvcN5TeciuinBkZKN122nRrNO7JYIDkq7rTJsHWqi5x5
k6KuPVDn/95B+98tQYh2BY0cUn/BoFbS7nm8n2m3Ra5Z8JmAW1hCsXkwLY7IMDCm6K40e6ou7C28
A3QuHjA/A/JfX7KY5apgDffkyqGweyG+3y4NpFYt6Pe6HvKnhBaZtt97sSdtwN2eAo5/D8mAGQVK
AzTTx5n4549dEdSzeRAMAc3e7he7b/EqXzBijMvvBhRj5TU/5ZF6dRYGFailXmWFeQY/EKVQhh2p
9wokIWw2VZv/mQSkq3Jzht+XwUkzKf/tsL5dIcSnW/g4lRf5xzfw5CcAJJRTG7GpoyB5CcuSLSYa
iTNKvzvb2ejZ5GQf2pmdwT7oYBkfTbyHZ9oGBNGvXYNBF5iPEp5ZGv7QsmNWo6T+V//MQmKUCy2h
LLc1yEWjSrAkedmifJGChU0yC33kJk+dxwpzGMQiYlJ8Prg5wGa+BNLgmGm2W/21/hiYP0fdf/+/
pft5WDZvEUYn/OZUkL+2BajSqungPYtu0A2RO+pyJUW6g65tyOJMrYsM3zmFFEnroU0QJDAMwa3x
NxYiHYHm0dc261Q5olg6V9fAivH6Ii5EJsjmW9ME94SdPqaO+SdzfNJpQFlwkpWJppzD/6WXETFc
Bcv2zaPU+J5kWYvzW9peYkVekiEK/GJpshIT1yVwvMcbR2gt3Hmjmsrs54s+BY/98+CRu2dnCAiP
rzalhueYFvxaf0kp8IM3HH/G2C9TBNwtvUzVDE9Wr570O3dvgKgdqIlXNxVvnGzQt6dDPcEX462J
CKw12lsV0Wrkl5Y+gbyiVuXFLzxLKTP99JYrPCyXs03En1ePd8iAFizmc4iB3pbBWuPxnRVbEjRZ
YryGmTbL9iHm6qQvN/CKimLD5LoKVkbgN8dvCETnChLscsRnTkjFuIJ4fte04ssPtDuwdjMvjEon
RF33hsgSOmbdMGEk1EzshbeThC+24j5ntN5Nh8F8CtZoHvGvxhl7Gs9CYnpE8OLlaE5+HFAAL7EB
u0Ru51FeDaY0WH7n3h4cJ6itW0yJFfWxBRZutjvTqZDcLZac4dtK8MtN8Npd3z1QC3B3zYFuRXA+
wqVSVdcpNKEUjbN9/sMpq88ZaUmVi+lEeYsvNeP+sTZHX4XZgjp9v0hgYrKXAlIDS95wT4RuHI41
ztHoL/wSdJwhtlGvGaQJYKqmevzRt0KRWafMNEraM8NNZA/p3oZ8MTliTLmGiticvInNTO/+U98a
IbTdnNA/2dKxTCz7WgRBMAap2t4a6tJCVj45FBIQvoIXWlgpUYplxfB+PJth1Sy+jGEIXphObFHu
A5nAEV/dyhOdvwCJe6YuHQsM1KXDJOyD9VKSybT8bRZOwow4wtbt3mboJ9Mi09KwuDA3tE9zNYA6
rOQtmBFblyErbleWePPMYViMvFAndrZ6+75K8s1OXgbBzOfgF7/QHEdfhe6+ZheyjDmFQ8wXw9z4
vB7aqAtup4F9vrU4CkHGip7AESouzvnkCj9/10Qi+oL4rBL2+jW6M+gnvCgB3zNUFxcaZ9Blwt9w
H5xirqT9KA5i0HSJDupY7hRfGzpnrxKsD38kHfUsZIeEyz70fK+eG4qB0x6CY3mgcDYR/7iulDyv
PMlvyGOrbs3fNEl/UWgp9EDCIZY1uHDNwl5eqBFnDWND7Nhz4BU4X7ej+sg0GBL7p43fwdfMHZKX
cYNay2T1wQU62BK9HOTKIHZ9hI+q9OOiMUBxo3IONGn9+mlPEKi+yEX2WAXsRluIrEigVTNkhggT
c45N/C3JejOGYeSh5ekFYrAIOuHCGiikfAWxdQGhdmd7sPsFLmTJ1ttsWjmQ+26CKBYeeac3cKrA
4ZiG1ayM1fu7z0MzGPdDQtAWC+6L0lW7cy2Km3X10O+rUAKflWScPqMc2+EFgDmh8kiLaTNTxzf1
Hj6rdEChVvVA4I+AAK3oPOb7cIZp2obuLYq4aOdjsNJSbDiJ7RIawC4xZg3NyZ03wQQyozwoxLdE
E0pGmxyTqQhQ2zX681Ak6Lu/Wej2YevwieWcbYboWSgdV3w4Fl6v261khaP6iMCMrS3gh2mfP4jV
dJ1t+QDh5HPgsXZzjXz0+pWo8Y2b1DY+EF/thgkBU1xbxrUkJLZ/f78yr0xd62OXkGoKfHhfcEhf
RNUT7hmgQkMHSZORGTXtva9U1TWH6+SXI7D95bsogka7nCg8JfLUsL5rtjqdwnKjRvWa4XiOzoRI
FPFJlpcORR7TZln4OR3L5xG3YFaULrzFTeXn74GdEfPz1bUtYXvMXuxqjjCcwLmy2Kvzmc9UnlGj
Z01RdIWn9Pr+b5lcKkSMjFcPz/loxR7Yh5QwpYuZ94Og3KEtY67bNwfnItw9vUN+ObvmYQznm4t3
dIZQwy3O9h1iMxigJFcj3U3KubjoOLVtZxsO2kzXn6OnaAIT5JPHe+gWBKe/bFsvDF3AUNl3BTO4
bvku6dqZ+MjytL2W5gg9xDc2pnF0qAqE/pQvmKZrSIGG2BEfyJYkS8fCxOCSWRdsgfxSNytIitcN
m7QDW0bTDpguVfMsaHSR2vuoE3DQPJBZhjMP2jy0ip3CvxgZ4I450bgU0d9Z7B0T61r1Va88X3iv
E3LUQjU4BB7SQXBUWJBOWDHfTLvLegxZhMgMtSRu/hMaJgA1O57t+MPIrC2A2Acijf2ws5ODK7xC
E8fYNl7npmZ30scZjnkwzVgt16Fs8EPJVVfifSun/TLekXbzK7w/89LAZRcYuNlK5jsM/VeBA1SS
QtWrSSC6UGWTwZqANm8rEW7B3I11R417qsxLfK7HS5k/BrSXRxvagZg1r+rR5Mk2uFsXi171p0zC
ifa3+biW0DJOQh93qR5KSk+4cv4vHKFgTjsWj8b/FGufCS7ZVRJPY4ONhEJNqBFVv9pXBJZCeTJN
j11HzAgn7SZlmmsJz5TIFGi/xExnCQuowurZ/LoG1GG7T8/+u+DSPnLfe8bfu2M7J2FkiQSiJu4K
RjxBChljJ3Lg8YLFpYbQtGlb3mPJTMcjNI8q6P7OdDfCH1upKAHjHpi52qUurvdCgL2dEBGE5q74
1222Bq+jvvihetswBR55v15+7Hkp5sM8cQdZ7bqYIScCpYgO2pD1G76t7WHo6rundaFU0/TixIPf
j+cwszfGCJiKfK0c2X9tijIa7FY/khzjeT7RmxmpGwL/1GXAAUM4IZdxSmjCT5mwsBVRGBux0B+k
zlhSEVKgRoPsB5vSspyt3tDVjsw7h8rg4q7Ap3UwqaeZxplv+EEgFKeRQnwPr7UYgtKejGjiUfbB
AJ+9FfmjxL1+MwEgEkmlD6j60ATEJTvNFBd3RdoMGMHgCcN48SJuVvyvIbKeO2KbY3gBxAImAUON
3FqnSygvbt8CUXHGn4PkxG4XZN0fruxqVATvj0kJuZgs/B+uCKBvlZZj/gWQ0abBasu9zWDpiLNv
0QMZj+YhGgU6FFL/zW5NxF3SUpBO5L9jkWANOdMvLXSxhbcO2X6SUYLSHYqmqqGeWIrILoY6K5WS
rqXoGkw+uqM1RG3QWk4tj3s2O9EjiyaJJjfRIz4oF+pAOhsZKqnI8Pea8IB+0otkPq2rtD7aS9UG
90ChyBYVWncWTgOHsXn/3DppXYvbB095I6nnayiZBd0AWWWFHaaKc28TwMlFOkRgzXeeiC90a4bK
HfksnBW3H55Vd8Ii2flDLV32/xVktr9tVL75NwoNQ857y21VH9PkkMLizGA7xDG1z9XUa1NMfDoP
WVxBsPCb+s6U6QiY7FDAJhHVVsOC9t4EheEAnn93p7WxB7Ksvkdno7Q9zNDiDEVs1GsL9RIXuzPS
J5Op3C5RwZZK1piq329r5ABuEk2DBXGayAVsxX+HY589mIv5v5o2opwQYnxJ1xiOkx4cYDcX4Oys
UrL7JY9DDeVJnEfNC5YaVWxSh87E8aIpVeUcHKQFjwfdXFZq38CykcM0PGb1zLMo+Th60aVfFzkZ
klZVge3rmjyoMRMUcpqa42cmI4BghPMz9YAO7hjAiEwJ6NEK5jbc8uxyro3Vy+WP26nmPd8fM7fk
IEh187Qhdfs/k9DNyPU4qPVTKEcsMZm/vc6nkUgvp0d0drDllNyIWUZqPKo7DybyvyLsAjMWNJO1
jzpIw16s8uGtsSu4M0PjYK9+8R/i6HYcU6UWdBKZ7ONShFQTnqr/SFO22+vHHZb7n2T1V+I/hkkP
IpfWyJ089wuHQGRTQOyIBFHGFhQbGXikxV69jsd0RbMx6OfdGLl1x29DaGpIlVJ/nIBF9kL525pS
xTWsvGQtLTLbiDSrlLYUJq0SjlNjs6otBojRJjsNhewtP+R7FZqje8+0lSrGGItqUaYDhF93dRkI
JuadxwWYZnOj2fvfWNef0tCD/xiF4Co2C+NbSfFlWa0/DRbt1mwCiqY+HH5KObOHUkHRCO5uUBKe
o2b6E+koLdPWM9XvgIxbznhTAOCGPf48/tx3D5UBhSEZdfBby5jWObL5kzqz6EHccQ2DVzIbxFTj
wRwqEuRhgEv63NBC4WGZrSfIATHMkVQY09tygQRjUStTPs1vfEmbcfEC8CBDq8pPl9+pQXsLJEH0
YqoY+rN7/mLZffSibpg/Pj65qkv4mlmewZRWsjmpjFSUnUUxatquDZk5Um4S5H6G0mooH5ghVmSR
p8DEVYmq2Xzlrz5AmXxRFiA/YfbNrl+LxN1qNJjrosBZcqBbSsu7GV3gC8PVKGoNHhkjY1xPWvFh
CpVtw+VnTsLcpz2oDj8XqC5Ei8NRkpEf/jzQ9+LPeSHkafO3XkAlCBg5bxNp8VbxBpMBbGwdg4kZ
RXNnsyBLlehigcbiVHAjP2N9j6JdVzRYLIEJsebu6X6e+OcrnhkjywT+ZgwhqN+sqmZBL8FkTmYy
/AWTLAOiH94B5Y051b8O9xtquuMB0XyexTTSG1hxfhuKSbcmH23tAAGOEVyl5JpUJy9SqBHK2J4R
v7/ZDpUIpPhka2ajSo1jzU8xaE8PtamWZ1PSHZVnDuu2zPJGGb6CyHQGt+wMew64hShyxAWcR7A6
NL9ixm8SnrY4mirzDVINsEpGznV7OL1DSvYxTE+EYWk/KCXSe7jZUGmP7xjOq4XYyGMLLIJrlu81
QhCE6l9rukig5Lm/YVeGcJiUK4XB04L0OgtI/xeEnZKhzmnDb+K6eazG3DMfu7yOwdgexMFLxFRU
fnffMsFF6Z9+zPJ68lTnc9c3ok7xfFE1mPvCJR23sYtXmPXIYwdFL+duRKjqFjePFoZad5NfyoMX
xQmAO7Zn/ZtYOVVkgIDWoVYj2hIMbiWpcsdtEts/BGB80vF7xURvhfCqQH8Z3LZIk/eQ+lnHBDA4
0EZeziW56glj8LLY40NKuHJScp9EDrbc1Ad37lVpvDlVZblRQ1FwHDtQ0pUG7a+0360Id8dcj0XR
4fUkfr3Xod/wNrC4LYjRqxLx5/2g51gyjVk5g18elPjePh6ypUH3WXJZKXVT3PT6xaZOCOOzzFxZ
/h9VGw7cVjGR9FXJEf1NGeUDzY8Tv0PJ8dp5UAGrVhN4xW59P89v5Mhl97XbHOIc27aaS5/mZEAf
D9OUVBT+vKu0xnmI92+YXl8VxkcVcN4CqUsC94lZ9cY5HunzyJLAT7S7XGaF/+ry6xFH8yRoN056
KzXWJVMQzFUOjZ7w92lAfB1reor6vqBBfCkUafdfIYXBgbUfVm/o6ICJuOH885ntNUp2Nspo7b81
DR7/mPpq8rzJQ+74OCn1uO8Rx1mInInTK6bEFDEzHgHynbDWiocgvW0V8b6b+4IsMAankEwxALyo
iqtMaa8JEx56yMyXMulEuDABD8EQOaFX5JYskfOyNnozGKwTy2d3xJjjO65w3lb0J+k+EjIOUcfb
p560kCSuOYfkto9Q5STWCCMxtVYMcRc32KNTB4L9oEoHI/IMJX5YJhjOtT+y+lyc49Zi8VBMlL0E
WJLPz4bRmuS4DD9d2dPdWt18hSEUt03c8sYSZcjuSMEAJMb4nyFWYpupHZSZVHnJ2Icu5pDiKACN
Z096gtRYouZoUBbqCVrV4Oym2i7VZKMYYcwYEpFpwU0Hil0OBtwPocDPmy3UsxsYsvoS5jA61BDy
Wh62zoPP0c7WKtuVe20auk/XfYqfiQHb4LcN283Im9iuJ9+Wc29T7mshQDMZC/Olyz2TKpdCmZm8
GUMFZZn5djHEI3M1BZ2SQiQiHKpRRzv/mad4D8I9TJLNerZ8UUZALna+a4aoMPSvBHGftgEl39LC
Lx0MRXDr4ujK2KZ0PxWMiue7yuBlNDfBbUW2F8q+blD0grGpvgnfRMuSs6XjeNDmqUWRed2CJ+K7
g1yCvQxnBFxIg4UyxUVFG8+CYseIIcLLqxhpW/0XiVXKicwdhkf8PUm67uc4aPtBFfdxl5V2BnbW
EMHsUcZFuuA1nTzrXNjJK7LpY5xgYpBvGJkrFHf1dPtEXMSt49Us8qPhr/BX2S5tqwwfHlgPnMXD
4eNJhwR5GFzNQzc4tumMR0nKc9JIa0NsTR27Mp5bZqvtWNnA0Cqqg5OSWvwPk1wsZbiJahqpx1Rf
o71xbXiFjX4K3hnkYgJUYDVUzP7ra66h/2HysjsUGYyGEadTwR7sAFjsfUM0/qgMo2lJrzw8+pTo
SM1gIyl7WvBQwxACJ4wA8OGAVELITpaibodENZboLIG/yflRpMdI+if0jf50AQbcDaqNCjAZF3Gi
V2ZimlXOSSLVl3YTD+5wvPdEzHD4G6foDp7w0L/rI6YLf9Fdye9sAdwLTN7xcIbJeYBxIk6xYhQH
qs+0QVjwShG7ujUF5kb3RJnZ6/r2c+PUiP49d9E/ZlhUdZ6cOxy9+dBZdAr4rNGhco8/hOFwrxwv
W9B7xw8KsHp5iCuLsf0nrXg1B4Wz+3N7j0nNEZ35XxST3pWaOi+Sf4u/NIuVO8VLvjSnufFj3TsK
yr3aSrxxW0j5wEuesNFJLVYAhFvDLRF9fQiYouTDsZvJMMsTUXjzNscMtlFm/F0VrkYYxk5g0xeL
iOkzAvuo9Wuj4KR9yR3kqRnaOt3rO0E+cbL0AFtZ7HGjJzG2w/oTj0fwKkX3Oj6ITQFVcGCIXlNQ
8CM6iKl1D0UHAOD6kH2r0fZbnbbr0O+S8erkCmFF+EPl6HGOfWesEhALJcZT7/jIT6foU0Bie0hY
0kXWKQ/ISbIKdij8w85NDaB9ixZT4RX+yvTyOn8oQxG9UacWC+tLzGvuPwj6i1MbPvP5pckb1iHT
gadCb4DnpFtUiu97Y/QRV7/MGOdk+/2l7iZM7xUdmI5z20uxr9ZqfPILW06S2PXcbrJvdXn5B7QH
W8RArOb1e6+S8Pel9BKtHL4OXqSbimbePsCxuPHXnGtD86fQ9GYASVS76y5yp5pERbp5AleMDUPJ
ML/1cfXfzvVjee/SJIZZNYmvyxXec+eZbgaBPAnLxB7vH7ByP54nqc2y9CJdKOLDbgV/dSg6t2C3
FDLH2LuXoiS8xQsThYBZT3foCZDJNMH6zC79p6iyTO11bYBbeRAjZv6KfqPz5VVfb/Lu3DMDuua9
ijMgf9yTDKK7YCPGswIMZPhOzTPucDm7wl1mwOJ+qzbzquhQ3oCb4Hny+Xs/b6glG+IeFu37h8B4
bVKZI2b5gH48EwijOcqyIVf8hX23eNARGKjUhqTRcOMBici72HbFRWEiw0QPi9EtavVpWbtlibdF
MiYRZFOXEz9t+HjsFI39Mr4kqk+axcfJMGqhiih/l7y4hoH8ZsNmeN4NxuyqXPO51jDtjwc91V5e
BW6KZEv9h2jP/OxbV44h1ns7y4CTJG+qGhRkr5DEe7xsQxVRcCTQ13268GDht4SLne3Ews1Agwvt
uy/uHKTb8VcMzgOHFZrGFyqJHMkIgon0nEKvnhNY3klfon/2+99drH8TM4uaAMEp8F/6DOQZuhB2
Urn3JAJcqAFukA3BFa7dqQooy0UPHN8GHJbLLQ1bOdl9o5CGRBRkRwX5O80Ee1L6veAC4PUqGUCT
jWZD9Xz+raL2zRsSKEbBZKlr7FrfwnD1u+Lck5dlb6YKcSWh/6S8e2LBDVkZMUMYGX/nuIAQYdDX
3vLaHvj6Mp5z2Q+gZSiSr1SLLwuOcMoJHf6IcQEIAUCg3OgHiCFJ/IYRzw5WafIXTn8Bc1otJzl0
/wm+sZ5qVZfgdodBy0zxfmHkxwgY2skqYY3IZRCa2cnY6lJMJ9PQQg02R31kx2G61HwryTkmG2vJ
6XGVUca1aV6OBWRa3iEpAIW9zXHjXAK+gkcwSDCChl4oQlTlmx47fb5HT7RAiuFAYbdlidfKgKMi
reGqo1Nn27DhEN5eNnWiCDJJJoX9SFYPsunMrFUpilc+LqpBsTF8oEIRrTACxZr29fh22A1D6N4q
Jd4z1Ev2g2TnTl/Rz5GDO12y4vDsUxwxfU7PapMq6Vg5de7attsGWzLbsr6TTuUE2awx+j73aY1J
8OVw3ueAj+SkmGIhE5K+2Kvi/a89YAnfAFOPHzisQ+t56Y5/q1UbVcGgeMsnKKS5Kd3doHj8JiCF
gmDa8Yc6CkR2Hd/xKBIRe7ZSt39znS1O/7tA7O8JIb6dIXFLQDywWRTzGD6HopGpVfJBiuAjNDE1
ZovfvEnhrJOZ/ntB/4qewaoW525npEZfdu+qHn5gRVv+NtNIxfnBX1304Er5Gx3BpOJtElHP4yz8
2Zw3rorPuwd78yr2FOp57tcWkRHkh5gjLYMjchbqDEuVf3XTpnNGK3+iEFp7hldfxJfSluLyhsK8
QHa29DChWkoI362FVF0FSePRx89cOk31rSvww8ByMJAEjVoGyy8CRC3TnQbY6IsuAr/n0B2K1LR6
5Oj1G6jhAWZtw+FfKi/kyBqIW2Q6nFFo9sFrTveyItJZ8AQUYyp5cGMwlZhsI4zqjzbjXyrPmu0P
LHOFPNgh0OfFH3PNT56qt7+hQ7/qWgmU7t7SimjK/R9KNVnj6hSmSAJGVrzxek5gIvkTd/qbYP07
tLSv/I54WVNWhLyUuWEjf83hBLZIiTeC3qJ5sUgn+addRlfC9a8dR6VHC4vT9g5KUykrhtD9QeXg
2xjRnOqp/V0GeTmOsCy0JJO14pJ87VCBDM3bwlrh6D0usOOT7isIFwHtgBbUyjO1DgAw38LnYrhe
nVaQwlZfDZncMNxP3H7W+A8Pqbfp1NHiI5r0PB+OsrUJD+13QMEGPauVhSieOJyAYICkL7+fQpu8
eLB4yh4sLvfVv0bNPXQaRwZ7NxmWUCo4SBMzfv8acw8KDbhxh+syWd3Py+eUc8Glv8UiuCuD4zVO
+xDAEvlJXeSK22Gi/MGM79JkcdXf3UB3VCf0reb7eI8ISd89nd8GT94PMRvVTMYujkYQjkaYW2mI
bN88g0qpHpMXyh7C6t6HN3IxwhvF7VRRIpHnYNVa9jOyfQ5G+M3OkoCnOb3itT27xYRat/opNyX3
uRTIw6X0lEQO3i24n/j2wgb2Kex933jXvtuzAvhLkEBWdszXyAdpOjydicMavSBkqHcyiWKNZ58w
VMy3cqrtpkJzqVZZ4PWL8O9sQm1tHW1g1RgNtllv0Mo+eabexl/AAIHs8Qcb/bzo32Wdn8uco7tR
twx/0y9yL6Ypz/JgOCJRasfooM2EuhJFd6p6Z8xQ/uJReQ/EJ1prx2KitF4xXYpDxLcTxhm7sAbN
3GxuOwfiu+PzpSXLi/7LiNWgQoyrPoBosRjNmMhRBMqijg2XoFQw2YWUmWgiWG7pKSKoKPRrcGa/
TDEzkHZ9BtNnqphE0u2eQHfx/0cecK8uEPpoTBS+K8pvdOAvvn5/Gtx4qu+ypwGrPqhKLx2Plhg2
q59aW/yEGkfF1A5nEDh45GNTFadiQiLvtKWQ4ZxZxhb9sLEZ0c3+Bg89iCEbmV1p0HFzkJRjAJgK
1bvR/8w7znIYOSHz87LDMhmZqk4eeygYSeIxWSh3Igzi7l7/VhV8I/pfjyQVooqRekejQl0pJOmN
GSqJBxLNMo43VoxA12BvSFGeEuaQPWi5XjstnP1I1PjwnMaz72c2A2ol9mYpCUewG/VE9dRMe6uU
n9kYtvmu/KP+LT91xPN+ubHo6dgYZ/dhvopnMgqNkJfBG++XbaSRLrho1+a/A9JcRvsl7DwF+ZYY
2sycfpz6UiBQ/RbOHbNE52RPYofTSRL8WxUNy10aJoNBSseCQsxTve5v7GZOKXjj9OuihmU21dKn
V4QtFo/BsiVzNOKepzWDPeMt3qAIBW8Z+2l200omQ5PfEPMcWmcXJhdkXksExrWJwh/t0H30Vo1/
6HYb05xghIs7XGIhYkbR36ysaZQqrcyEXTb3J2Y9lTFdcFrXw8WPLLtbH6Ts+FYgF7QAmBhUJnlH
w2F8QuGGQzVWS1/gJfdxbaOWHlDOgPZBF6KVyK8q2GX9PovzWq3n8OXAg+1lQ8Ep10oHr4P8J5vs
IDnwmLUpdFjrEHa4Mw6rtBg1/4iSrPwMDxfsqmIYHjbx1qIvN/YDUAqgdduZhciS8WxoN6W7ADFr
m6id6DBoQ34IV8pZo19w3eIJMO631wAY/4H47TfjXZQketXa9KDMtQ2o4mlBK11vcwOFdnC00qPs
SJQzAbCwrNqhGctA1uU9HRgImdtkhcewXbQJzKM1B5njMhfRQQy45mzkd/lVbn8y6qUxjIqkd+Jf
E93lNDUS20+Kh2qMRz79ZUhagHUb6m29voVT0/bcBot1O+NJMPSOfZ04oSjvXr5PY2hGHUwjxeU2
P6ii2O57U4BPPcmr+RGZXv9VwqJq7TWn3BrQyqsc2zcw3JwAbnitw1rOWdw1kS82tj1BPJ7Vgv+a
cVWLoUaZjo4To4eF1FLAHyspZfEmnr9KaIAtjCcHCrbWYWpbANHMllEApItRbI8JCjdjtOpTF4RF
ntOWEZmuseiedYKYQwUnyD+udnlVsNF1oblwsFvHsaeFpj6JDNGsWeCOXwvX4qEv2eNgRpSk0Acs
/m8569/FjchmgVOrZpL9f+x71WAUqwJ4TENG7kvTMHli9mWdvT80UnqBbX/+wcH2qKdTo3fDHS/d
JvXkqDH5Z0FmgNsMvMsIcDvB7U48VN0CBBLaQ5c01p7vJkvGsgnYmTzjqqQdcUPBd4JzCSnkPiTM
fMa0bm/61aoMtLjSwYV7AI/5dYnbTkSHUpZttGLTta+7y2ImIcvKGpIHkBd9Pj5kpFU9UoUNEysu
/YVF2bpNzWyzpzCOX4Rhvj9c4iDIqtgLZ03vm8IMouAb1XBjDFRoGAU/gKZItC26R1Q5YRbqG3m6
eFa2LGkBpBQUum5Gn6z/McrsC8Q7ISRszh1aoGrehxOMyKGesfaN+ifrU7+ZpTxb6gcFx7OLyu1S
GWzMcaO7IcUF3IBrR8QIuo03hnkkG1EJhWtkahs+Lve4no6I+1HclkRxSsuOwpweQbFpXKqfpclT
ckyyEFov4puCybzkruYgsD+bzbTXDWf3VnePD0lUjQFv75JcWSmooy3kVLZFHUTPRMG4MmguX8Tw
mG6NfGUK4FcsMtB45txZjFTAS3RfipSZZOfG9CwPZocMY4WudIc3EUVcl3IwQcrdBTR3060OZILK
yoTJK9GDzUBGYWLj5OK6kRpxq/e+7qVos3/fWKLTsyhwyDyt57fhs/Fp4ekS2+cRFaBcGl6GlPyJ
uobYxhyXRhCXx639aezbCfAbfZw639xPm2vev/tnlS+q2VKpUdQQYEvpywKAV7q8gD4EIMVtpG0J
p0eYhUjNGvyl2znEv81F+Cdulkhfr9SHO3SPWsIOUpBI2hrXaB4pYegmB9DOl2gQrd5OcHJpqF0D
2clQgE2ob83HJXLgzBGmjQU4kqc7awWpxc5eu9uji27CgWbaRdI1dkNTqa8rQj3F499ybYLA/wdI
jjaceqUonHxe4iB9eBKCyHyzs45q0ZHA/QX59MIg7qjFMZNXoZbT/7JfK48fatHzsnWiABkB+b2s
cx0eXr7R54GRLKYryFaj6JnKUMz3Bh5emy52tzs55FG2VQiBb36wTIdjZ5vkmRiyw3hj3nDSrAVc
AUZWD67RzB8uYqc2oPLixva0Q27w4zllmLISVy9V2rzp9AuQiBYwo+kjt6tqYd10xJ8BoXQqfBvB
xKOOB+z156m5OMeXfR0+G3BxIiEDqSEf1MZjObdk9mz16BcuwKf89CaJUtFcggMaCPPgHg0Nv1JH
M0eOTnWCQx/8ePq97FP82aMp5rXs+59P4RG9i1UJdsiNyIt3LhtSqVANfOK4hSPrpS2tkFWEHVwd
RzERCJnctSO634n0DXGv+zKdJiQzWlILvUdr4lSO/jzVKbiD29mqw0/fZLBAGZS4NnxhQ8e6XJsi
pGQOPyKi6Em7Lee2BWbXH9gUnfvU05tOvfU0VcQoiXVWk+nhQHYmNpZTfUroV+nUyd66IB5mKnPQ
KcMoLNIlUy6gIc0xv8DUyYlWGJK3UbtyfLQk80dxJ1rs0ZT2lfHK0A5FXK86/o8gV6ch9D2rgHmL
uCa7LzLMot9XXrUF69HqJ4cDS5y/+RTIJ8xu1Z/NEVp/SiR2ZTbvxzObIbRzDs+XVlUUchi0GXbV
W1Ccmn+UIaxeolmVa2AzSYujEXwCUyLzBXvElpcSRwSnAzV8DtRllx0TZxyRQ+it/5No22+/GjUi
wjMAXECi3r6pNUbrdiaxT2VIKmkY3NzNoc6/UaaPdgJmsaB6e15pZ2p3cESUbU0Py+tPz8zojwv7
gKGkivOB1U4OGVzwkflzJ/LXaPQ8UTZMBA346dcJ+oWNoE9rw4dFG8dFY0cD/FljCfvaO4Xk5N9W
wqZJW/AGQyYXOkyC+JvXh4K5vvyz7uJQhK8yjIk2xsiN/C5R8qZXam/aJQjBh0fLzXWB0/UzXtn8
L4kiWIrlx14CMQjSN2Pxj1fcMzhh7IuarNoPHbX43qkK5SQBsfJYy/FGYsg7DGWhms1+nP+S2PY8
e3jzbd09EA+U2mv+I+vjuGed0PBjoDPOPszKkbi+578S4mEzRVgBKQHgoyPiaD0SANxFzq0+oAtV
UkKY9e4hu0H1+Pj9m1qWGSUO0QvCIvro2zm9n0vTwdmu6ZmewoNW7raUloGKsnVN0qg/q46p9SvZ
0V2tWbgUjf/c51Q9SJ0IiSSRnvOF4H8Nt9LKUAN9G4dk5FLRQXODmTL8T6jCzga+1KFPWO+7WNoL
yOYRFvuPVKmH4CAXDOkOH3HT5EXLbCUFho3X38G/XsFbZgJXdMFO673WY17NPEOQsWTnvDFQ47Ee
j29H+1n84bDNSGui9AAfRX1B2+7Vldfkt3UBmjWW7MirRVriusQHwgzA24DzL58CpM5gQe25o1Q1
nQ9ITXrldRBCRQnJlcUlmzUdDeJaXHGj01+nKdRDBJyAHNd477c1AXqm6DdqxX6hVLWK8phUDgAG
/U9NmFphkUTL5WzsAG7sHq9v+YD1fRZHrFVnmwgDdAlEZS6x8I9yCbgFOxqZK9IQuDSWfgDYfaqP
YFwOoNOdEzQUK2hdNBMT870h9SFkIt79/X0L3kyW8BdQl5Azu80f4cnhX7c8sZnIKtM4mBe+6iH/
U+xyTz83kqshtZJ+P+J/gBb3A5CNQN4IterorHtEzjCDUuyfb4r/BgsIJl0ZR2DNS386yT1C2z6U
Es/CsfmbELk61x1OPU/9yjQuEx+Xfqa/qJQQ39xsBU2Hy1sHT7H7ApduARqBpFN28iX50ckPZpYQ
YKkEIG1BqKa62W8agBZ9gjKBcDdEDq2zUA4DPfwgyftImHw7So7B2o7ka+EJtcQz3TlI6px26/nK
Ln0CYTsSJEujDTgNuwZXFUDpMl8bQkfm/LAGJ7cPxCb6Cu+d3c90nCqA+3EBoXH5806HMUsaoRVu
vJmzNeCthXuWJukHmUpFWCYN6p6+4f5DVsZu3Rig7lO8UG2KV5yUVIravmevA+ML975Eo3hKYGId
UGRjZlugUCoHpzc4Fd0vRl45IfNq/C/8Yk4mZtQCQU3ZOiC4uRjVZP5L4/ImDDzzg2u9h8Ay2bOr
9g0Aa/E6pO/H4H1uCu1/IM+vuvf6MaI9eaUXsi3YI+QUrilOBmR+LI+8A8R3QmEFss6vqnpFsLy+
ACezZr74gpfyD34aXClIr1u5ww/TdcoK72NQWgNUSexmyzP/bLwg/czdKR0GWugtkfYtctDdWeKY
tY1/4hjXSvlN3YQigrfpaozpjeadZYFt+OIZ9t5i1gIs7ow/eYczYAk6vfqFJCH1t/ztbWLzOgVo
FuZ0FfZzd+OmI4SFf98Tt2epzb9WVeabRv7GcVZgCAkPPnGV/6jlGD8V2TEIvFRRJBwYAVvkg2CY
+gapIxMknKkw9P09rBrpRlmvQmoShLoodt67vChJY79VDDuj3p1LFnj35C+e2/4stt6N17GjxJ9f
0AIRoqJ4znCXAgNcAJAHrenLfjhrdwAiZ0av6nEoghMVbh05GEkqVLq0wBNLuMWhFjfizw1qgD0j
SJhvdh1RSkf7pA6bQDrnvrkTXlDMNIyFTplzaMhMOMI+C4sSyh5yIn+/JWSfNuu/S4OBcAdRo5Iz
lEWAaG3XaBaqXJdODg4597jFLGG8Vjv6iVbv1nDHkXWQpQkayUa1BcZTqUB7WgqqU2kfPM4VUEKy
D69o4+aLch0NPIDZ5dZBOmnh/OyzxPfmTCtLRFF7U7VXBAU09pStjKgPYVdendv/OIG2Yohqll6S
Yte5JxZA1Y9YUR9NciuoUnEYt0rYm00DpMjoO1Lb5V15jC+YF7uiOmUkwOcrflv1WkTNvtfMHcNK
jJ4fFkW5MdwJkH6MnC5sPMwqHTxf2DKyNEpu5c+cHoo6otdpiLBhWjEN37bJP9fBQQm8Kq3ieAqG
RZC2gCZ1/gfthJCOheFeKXdnaMwq4V5zWP+3+ICSq0eRMxSW8Hogjh4yt+5Qy1nfTD1D/igvU2E3
sMaDSnGhzljnUMMwfnG0Dfh4VKrxzUC6aJ6yD9tgBryI6Ci+YZ54IC14nSL76OseGUf+lVj8Vavm
5T3pUcvuVtQ/3mCUaqg8hNmvw9p4+tRLyn96mI621n2mIqWLysa0kmgV4kcCJlzL4kWRatTSss7d
dkZOx91FfTdUT8aD6zWawij2J3tdgZgxHIxu92xfYkV1GBzZavHpj03o+WBsY8oYSrvAuYTLpuzx
NupGcZ/GiYSTB/3ryX5fnAxCRYJasXdjzuffhws8GCbV9+NcWq4J6PIH88p507JMAsAEF6QTf1G3
qrQ/U9EKpUyszNUYzRZtPmDVj+kBb0uMAZ/ZJSr1lqczSdbQWfTSbSRqgoLzLND7BKGXWvIJQuYr
JD0kXwKogB02hbvFMGky97AyhMYpk7HCGvY9ZVu91CdFWrGYglgaJam28OGXsJXuTwgBlzmmtwmi
JVVXKPrvGcag0b7vySEEGyRco7pEWFa/ijBwomS81SY+sQ0snbRz/+qkOeoXemcFcblrWxWOuVo2
sG9Ez14/jQpTqEydAtmU+dwPtwXB53OGNqBe3siHORmk0WhO5PLnAUg4dEvrRg8F+6CWKKUcnfKH
rLLRDXvDsI45pVJztpkgdGfaDPfUyO/BuzLpPr/HTuETHu9Hm+TBwwONKuho9q0jbBO0850vj5n3
b0m9EweVkVRD3L7YGPiz3ihvJrPDqqQgLwTTuk7CC+PI+X6Und13SEri3DGgYpJoL2uJkM/kv1UC
SmTPDIcjhaAH6E5IZ+8ExNG8b8GkzN79+fuczrLIFEfqR55TPJwfhiV4867m/uV89pUKNU0QpRGH
MYTnaNjuKqhMMzP7i/pZKscfKm/fEeVt6dhSSChbu8oMX6OgsoqAQloLA90arrMKxgXqSxBG4ooh
EMrTPjKjmp+bOC+15Skk/nE/4KIa6ASxRk7gGQzGuGs7x+9KrvolBAfhkihApN7P/npS0aRr2Lio
syxUYs8gTsPcOozOATRxKN9Dkqf/qZrpvAe992JeMgx48Zrna/moDxFL45WYk56o6Sfh6r2TJCCj
eWnH9CNqKiYNDEs+WghhFMabqKJhLm33JjYMski/G13Hn0hgxX/uM1L+q9AAOyLXAVfx4/htzoDy
LEIGpdSdV0neuspglqkXWNaOViAkkaur15WgpcL4moNp3te9I/6Pi5bjVRPqI89ZekSGffYx+rII
8GTE3Dxc81tIbIXtfqcuyBV4E1vF2JmHTvOr84iomZyXEqBS5i2AoCI6zNR4prFplo+Ra+TTKbYh
aGhKiFgAsdcVjI2vmO9nPsKwJX7kGxrz1uwWZ4nE5OKaRJhIZrFwL9g7Bpgk9+TwXgoQYDphFiBH
KZJwjvRCx7+xg99fpA/GuWWPwyjqULGZZj5x4jObrTZiGT0DA7kTc7kvOdhvFe71KZPUPSrPHY6+
iPkjgitpTUPq1Be3YY/tIFbxEwinAsNKJ/Ne1rjmPKA6QEwEH12HI6PGhDbaeqQhN25Skh3iBK/V
CmbTTLc7CO/RA+l1L1VmkwHft/NF1W77UlNF30vyoqC/1d1OYL63byDj45iA+SNWWfiPYBt7ufR4
ghzC4AgTOXkSFEWWxgNx0e0hg0W0gh8gYaMR4Y4C76w+9ORGrg5x3ycAGflQ2sgZlWz6dDvr9aQm
F3wkcB3v4SFLxRsLkj3a9mf3mqIQg+hd5qV3CGSm3ah1rW5rWm4+o++tnI54L4mSsM0UKPlMX2Zi
2t6BI8H3RXyIwRvbKj8yEBxDAS9/YTU2ZomKP9E+tKxKNikfk0o4nJmKJauY8zzc2rSeopjo8QUn
+N+tiA3jjpqRApqrJ3tcgnSGPR0k8qV/+qlYk6UKZ2Nh9jFfWXxeGLfR8sT+4abQ06aYYGritVZ8
BKPDU+LubNpPZRFiJ3EtktMMExNkYzD8SMG7+m4DczbRK2fMEMSBMbPJ4uAm4vhqdJj7D5XCM0Cl
MpHgIwYIO+xYcBw9HBSqHZcF6mhDcd9PorhFKDoO+pJ8F386y8JgT+PHZKjpVEFvpqO8HnGglTLB
5k0W7EvNP1fdlrxcppMBLU+vV/cD7RVe4eHsj2pge8faix4EPoK2Z++NkF9VTeRBm9qtvTu8C7sG
ZVbtZrNQhJjNyvPReLHlzbYC78xHqgEGZpkIurvcr3qm3OFr/cD8eNP+FzYgnf6nKKb2hmTHe20q
FqMmAgpSMEPQL5lRwFWUno4QCz7nlgykZAFEIWvRpFSh73jNt9tNvFxQlP7fxrOR7lVfhCbm4zUU
k0eG+59ir4vw/zz2+HTd2rqlebuz/Q1IXjtrls469c7664wCpc/HwRwcgAVDNmxTsV8EKUllYdla
8VufrjroMvqqHZ6hIXkSdWWi0FPWbYu9qKBJNvkt2XCbi2iIeK71OT8vLifIObolPQ2hC/tkpqGh
RIeiGEYK9+AHXgmiVL0tXFyDWNK1XQ3Dx7ZMOFG/vOktjsRCwn3hdabenh49fLpK5EENrKAXicxG
uC+1S4TEoD/ngxOWMNMwP0ZQTZ4Es+++OrdLCNP9GQeIal5/CO/tb2aOL3z9qzyNB/2trGW2vwJy
ihjTz7Y5l/XuEOlpAOoFq84BQgPP7MxN5SiWk6BqOPOiQvlrOkDrSVYm9umpousRF6rLPGMMCda+
8lCsGu/OUSKYwXz82rUyzhJP7pcYEO8yi7LYZt9dLFO1xFpCPxbHWXkkc7ChlPCxgy6RZJ+Vimrt
JVOt73UassBO7Kzf7x9faWuakfxCLQGQ+CMQ8xnQ4cZqv9MBv3pdO+WWtuW8ZOOO+JeQZIt/zLyB
cJ+FQWcYPxhAmxUet2vD5vqNBsSC0W5mwPGi+HHqjFQVj+VCJO+TTvGhec8wbmdzwuLJqOPSwslZ
/xlkCkRvZylU6uSEc6EhRFbudvVxwCLOM6wQGoj/PB7RramPcr0j7T905WfJEypSwAQKGnoHKlFq
o8aa/c70ipG7EvuWPwdhSVe28/IcD/WmrSjcQv+j0yfLMfe3LXZtn2YLhNoSJVoVaryE84350I0g
Z6eXwPQlZIi6rDoCLPEQGi8PdMAklDtDMiZ8yLFrAmTuHvQE+7Pp3Ub9srFfphCiYtlgexdM+lUa
Ll+HjgFkyzfUDD1kiHpVlz17vw75HKEAU/prktG2qGVc9feQ2+Ci7d6ZmVtbhpRSPp6wvbawYJq0
v3QW/xaaKTYDpUX48w4bRWJ6WB8Eh7equq/lneq7wKmk8vzHVdmatXpVE3GjEyV3232co9A33HRQ
2oQOHs78LP4eRygFzVZBgVAdyAIRx/gA8KKclDZOMGg9Vc4D4rbucB6AoWvmxrlsR5+HR5Tyg9wn
PC9akeY3yGtB3gG8YxycdN6MhioHFU7D1j1u01BJfmrPBzDUiyfPVwauQn21XlYzt0DVd9zodhm/
5oCEf5oQpDFRP1n8azST5Od51f/t8Ciu9iVa0H/RLWoJvgEJP+FnvBO4p4SXHX4kNcOB2ZYr0NMR
22xQXdvtMNev+ygoVTY2dzXtaxTUdoSlOFeRfCaOC/NtjYZ0gpvFS9QhSrhy3pUgksF4yejBsTiz
RiD0HYgLL/ODZyPCN203aHkmIT1MZoS0ZhuRmbarae6A8OfA1LSB8QWX8U0AR2mrKjKuful9VMt2
O8Kx53YHgK6+ZSgrTcoCod9VfYw5/tvX8YOL0fWJRz+HyTuVXv9/Kx8YS6nk8wdstrRUAo7/gMKA
E9OGbvLDLHXsQJqc7MOri8TxCpNpmtTClvyOkyX8dSrXSYRrI8pgEIFivlzYj4HofhPtqTrFWiMA
PTwnsdf8tXr2THds8WADhsuU9hztZFBrM+7hgevXmCmjV2CIgZtKBmg6P+K9e0azA20hwkFReUSB
IRyosAWz/qpQHbWl9VIe+B0yaNvULuhLIwjQgimh6+ZlL5VP88rI/1Mh9Jne/vqTjZ+nIXnhCKiC
hk/mHh+LsPwY/IV3xXIw9MCP4ZlPV2tsn1lDR4PKSPvVGLJthkkn6/mSkcQpaIctvryLI1dTkfKY
iyf9TwQ5sFYarPMnJNUGHT05NybzrHx4mLjlRL6HoFBSiU+cKAYgp6EF0/0RQgW+2PmkDPcJ1W4i
zM3cjM/osW8l9ppfpun/WiItwbpp2z/mY9MUgVYxb6IDl6NHoXpAmWr5BrS8A8EV3lh2E/X6rTNl
I7Vr1cw/eneueDGaqCDilHh5fRESNJd6D8HdHBsAzKhbk01hxqzywsYHHzBYHvVq4ncooJ/8TQ3I
NI6pZvwd+AIxwH9lwP3MccC7CNc76Oxq5wMcP/R5VuglJs5s05TZ+jV5d06tWaHmjytlA0WN11+t
za2l28XucX4VjdV/crRlHhiyzsdt9i32iG+zjcc1gnoj4BreiQM0tdFkd06yGi1YCizbbJr4z5uj
drfngtjUOKW8dkUbGIfJKsQv6fFHKCUfZ9chmtB03iON9M8ps6QY4ogCug8tq29DmXbrHmiLb2SX
mvP9pQmHV69PB/AIhSxVHcgIiAJ9SORgmnTqRflm7AjLVFDF7Ue8ZwrNzcoOoRtgPuo7cKe9BS99
Kd11dNlf9nHyt7oacKeV/AxXcNiGHqnLbwHxDqBXVngdcXbLwfwjRRpB7nXur30UwejGHXzQ+SZX
bBKfAIaERy6kUeClNO5yi2yG3pnpLM1jx55jiG1Unt0SgbyXJJXKcmiudj+pBs1tRO6WCDEZxzj7
gGlnRQHqAg7DnVilDSeUy+oqIeSFt/W5kZmFO/UgUBj+BUTZEZZKlNhWk9wvz57qzIEd9SysyDqn
P8wuh4nUir+bmc7MwodfDMeKQYUB+pfcSprqWGyVj07jyU/J2pwxJFho5TOEwC3aiYiBmMCzQns2
vIL59BSe8j6moU8/hK633dFaPSoLHS29gnfUyyrWGe4Pa4SE2DktaWQX3RZcn9JSdIcmKU8nFFdz
ruKx00SWDpI12WpvlmRq6jOETAmB4mXaO0lz2VSoavKov1A1XAl9L5MRdgW70JaVR2v3Do5MqHZz
f0et0D/+mkgdjLcj3oeTx6xV0xbmom8nsLBxqDhys14oPM05/QyefegSFH/4bos+8pksRscfoxj2
9pSQlLakvm5dps5qgYODMXaQMnc3PMFD+nWNrOV2wuI4S+HCuM64NOJmIjWppxuHTUBmjzud1TlS
OcApvU7uewUZb+cUr05R+UYMCG3Ncdpsoxl2I9YIBsPYvvNB3opReDTrkogumnSWm6gmF8tU5VUn
hpTaVgXf8vs8+mmfL6ZwBqSPcRcJ+9xrADOweU5sJKLiLEq2eqwPmgwGagSeBPFJwTeIK2VMCYTS
Bt7KMIdKiT9lCainPR+BCHZjARxs2AkyMmcnVUZyx24r0UrPs3ws87IyM7dxPYSoAmAVD7D2x3mv
jR1sngebi4eKKjh2/r7G+kH6bH3D+7v2IuTgfSMYhhIUJp0LBcaL0lOkoB+UuI5E5crQ+yTUrqdQ
hTpbcF4IJJCSq4rY9/8kHoeSXrYUrLZ5o0T6BB1VF8MlGGj4RRuRJYdXNVMmKzBGO5MN9fq+BrJQ
ezRudMlVQJLPMhdE6dP3jBLnNjyVZVZNwULReZ2UnUHbERIr99ROO5veFsZzApkkK0QsCqpqdO19
Mm/kIv4hYAFrvt4vQbXmqyuMxR6P/1zV0m++R1B6Y98dKWjCXzXeotN/RbOq9nSgRJwwT5GwzeA+
u0HdvyD7jeWlveSPsuMBF2kl/6iPHYKn1oC802E+fWaaxLwL7ba1JfvtpHupTcmZ3QpP9wYPGhlK
NBHJRgZhld2YkRIPndcrQv7A1iE6CkiH7w5t+xD+4MzXYkBMJiv8m8KJodr+LzFRIO/le9p9x7+d
jtNUqLrBqnFAx5yAtaW2VLrNXhxfzsKw9rrC57spJHXqpCUC08O+qiwMxao+5pBzmsC18Oi69Zpq
flL94sh+poLMelbmdD9HC1EfgMN17rBjlOaJxwkE1M7+aSymR8avytBEdPxCes3MJSZZW5cTBF0K
aWqueeNMYNaioosTnNmezh7AXdbkbFXEzwBV15pxC5p08qbNLKTyY8cMLEPgfYBEka/TGQHtwBnL
GKRStcs/HALP75puw5DZ45tBRX9CsDHH73o7ZbfDjrkg97QIp2sfuLQYnn53lj34ld0zv8/vLg/5
TaMedKp2GpOivM9YATvTBl97KdAAN4EZm9SxSqwPTP6r/c7bVRhokuMkAtmUu3/Q+yji/0tvLzbN
29ZNUHPh2g33POCte4/snWZAoMJ8huUxV8Y1Z2uxrtLn3LvxdI/7l4iXv/YDigl1RbGa8i04Fcce
BYgwcpxKD6t3jHcJ5GWymiRe1493G9Y+y7dcv3UG4Nvjz0IyJCJIY7lwIObjajkWmBXPTIB2mWoP
i44NwVBZ2Oxdk4rX3Uvddet2pjHdntDSH/OMNnU8VtrZ4McF/vQ29i9t56U1I+es+fOM7oqCwzsB
jWreWbfnntMzSOB4XdwaFuRsn1VsnSM1GqKQvyTsEHF3dpJ7i/ljrgmcj6/x9ubjlef0lC1xSGKK
NrikRvqGwwDNx3u//QsDqy8Z+5wp+UOYR0JF+9cUlMJHLPUaYCgYr2oeZu0fKO7+2YXc2jee+tyZ
kvHa9FjfpzclPFGm+MgsCOFctPttIiRgH+AQe2avEd0WAy1tQBv6km916oD7JXU+8cgVVQNMjnM+
oLM6ANDvqFbNnDipKK2L/cvmRMgMIHNgjAziOLEwZWtVnBhCGLOVB3cYGkNRndP+EzbPnKIsg4Oc
97J+yq2Y+dhQD+ObKX3PR2Y2j7w8ntU/9d8X0mGg/uSixQ/a5MCnlB33LccEzonCIJaAtVyVyQTR
rjHeV/75xFZcVuncax6w5Gv5LrqSwrf28b8l0O/ePNXRj86fw4ksSO6IRg54PtIU41HLr+qo7eYY
ZkbHf2NMVpTBppeAu0F3Xh380NB1pQUKYcfcTuuG3pxSvY133TbvN0O6HkVRDxX5FapMXfJBTCR1
ZjojDkbbn7pM7qBt6um8N2AJlO/uH15lPUxcpyShenlcNLXfQFme7Nt7pqoCT95eq2UecfxcBILO
5nD0bfnVzxjjgQxzwrtpG5a5SldBxVbOeNmtxOetFByTlTmwxGETSIhOuvvb7uA9lp8vk+ZOn977
CpEogVxV8IkxRT5hEN9X3Uu/iMwHi0d/2SSrKPjHxSTr6vFtHHed8l3YIOLuvDHXbTTlxzCjfieD
H0ZDjhGS8CRj6UpM68Vm7xbfnWDtJLx+x8jo3/c/qeXny2SGyV8QKEf0+58DS9m/3S8nhWCU8qnN
cpXF8dMcZ0lB2TkJXvcO5xpQiy5K+yKluHquaYsjwp+PhcJ/XEGvxKl/z3s3JAVs8rveYnA/99YN
rzkrNvaiJ2tPYh3FlfXzXReVCyrd5zg8RvEv3Ky9dFIGplneKCPwA/CowimJ9jWhIz5mrZI1g9gK
YhH2Du23yblvnxETe0z6Sjvu+c92UXruWxbeBqglMxpeG2/x9k8uVHQkjjG0c7/OuaMGzwvd5L1d
gr13H7ipXCCLAlyfNBTu49NHG1FkOD5644HP0Xolqvq85MPNQYnh01ccuDJOb2s2hSiUxrPS6ixC
tySxAhZfpqE2Bq/KpuCDLdrHERr/rypwofYuVx5+VC3lYGEgxj9SMa/Nwa0laBys6cNHqtixQodQ
fKlaCxjPezgUGq3AMU/q3y+K+lrAHMqS+F22Pm3XWzpup4sL+cFCPsWEo2gF0YFMENPL6QyQWPMU
tE2EphS7gM3rxb8ujPJnGgdk84TNaUe56s/q9IVfROrUHOsENxIiz7PwXQg2TVB0Lw5gO4rFGzas
hxL76GPRy2xrs5DWvISeZxM5wdoT1cRwGPKQA+3ZxyVGApfoszes1ed3YTQ2+PjRP+rcO6aHeUm5
mdltdEcuLDMUY+EF6zOZFB9Z/895JZ1FA8AMNpJzec54fcmaKnusnoiHRMtzoh0sLtFPZkh8ZKzX
yhJVZibRex0S4R4j9OGj/ARYJZZ3obaa/u0IvCH9+13z2b5lrAEVgrVn04vopq/ccfWKiqwMF0dg
kmT67vdkrpnthy81xd3KwW4DTxrdBRwSVfjNnvrnvbBWcwzX/y7z2ILTc4xSYTT3pv13cGe5Amzs
pdJSYitDxczUsxXYopR902Z/xEEtJziGr+DLqE5qZ1NmC0oviztiZhQBx7toHCpiUqmaYiSiTsUb
GwY7/NWImscEobJAvWWbgP7yPFKGV4tRQinEtD/S7PeO+NNKOxVYLD4JoFkuTJSNIBSl18Hu0yK5
elFtneDy5SbxR62oR8BPv0xooBcQRsxC9zAMR8ZLlNS5LEhf6LzFXHX+ejzElRVr444fuiSCjNa4
S3kOaRlP6wkDaoS+fT6KFCo7gf/hVCOWull06EXUNHM80S++KmNXHMoRnrKzZVmJ4i0HQVSoCQi3
HplfQ+EZpC+5XV3l0gRauyWKE3wGqFWCp3ogRr7bo/fB/DniYdYK3HFcatd5T/FVjJnfxvWcLzvV
ed3CEXu/CMddNX3jSA91zgM3cdMG5ws3zfmR6S8oMKJyIqtX7JdkXsTd8qSkzZU3sxRjToRp9gfh
wGMM6ggjUBQIB5wyFftQVkMo40ulpjcBSUA5DG0kxxpfGpE44dgshUINddhxse+bJm05u+1lLMED
rYJWBnp2HD8AcW6qRvrf/12rthH2UU1wRpExQUuewLB3HwR3k2HrnnDJ49clG8Hh48mzqD8s907I
hGxej6oz3pYL7ze829Od0BEUieotcovmElMFH1LHXnSIRRcXCKoflluSg3tb39uBS19YgXQsnQRh
IDhInk2YoO+Rlbz9U4XKEULVgGP+u06XxZmge26KePUSeV8dnAIK+zx++71HTbFZX8Om/v1eetMF
9/I65ljitvlyyoOac6iVcnPUZHzks3KUyVKtAE4uQBE+DpEgPAbyP3i0wC9oGaQAjnYpM3sBbYak
7gbFCRHdydgRQ75SxeSiNghfSX7vYXuW3Nhu36S9obD+gawaV4n0AKSJrXHzTIcXjIvs5iI6jPql
nH7VegEWA/J2lzqHelxULTRAfWQacZ7nKLB9Wq/eu2+M5HlUV/RtmOR64DDajfguOCjzMFx+7X2X
IWUFnR8HeW1Am45BSLFUQUr2SpJb+g3W92RT671Pj5M+WBRK+kHczkhC6ofx4VP7Wdn3JzCCOxH3
eokoWWoANQHIFixtqVlFAveEQiulFqTiVMPE2ju+Iwi1iA4OZeszCeAQS4k9y5HJP6T5j9PbR+2k
8O1NGPWXMbTNjBE8dOYNCxWP4ueDB7XnbDYouNQLJxxOOn7OMGPjNmRDDPni2dGhd6j+i23T0Jnh
nchrgvb4RlpQ8f3A3hf57T+vAiyH/YEFXrK+75OTx0b7dTFwEEz+hPRDi9e+UoB1/S/HS3cyyNyK
GThCaYz6SrlesLiaUAcDKHL5ioWbrNtZSBZoFT47EATissg5FCBntOlw/vZYSgNjPPJn/dyu1lyN
f6Vx+TqlF+HOGpNXJ99Rlgwn/5+RZJ/xgzacp9XrZc9BT21PacgF93B97IqRasa1JTrLCSlN1Sr/
G72tVXqjHzEyErsA9AXRLaDBpiou2Yocvtw9W3ZcFG7UrItI/MdTdbPqptQlQ0f4HvMk48to8/U+
kGUCrz6TJYJSpdQDi74ZOFUKlQA3xfMyaH/MDcocZdcmrz1484JZ0XpkOfbe8TsVvaaiDsnqpwEd
tE+7+JTSaItIF9B/mlPaa+XixVmzr9dadsjCxDtDA/CkmMwiAEgLwVS0GGLM61Fxw7aUThxC8Bfj
489/E4ZgzZSH2gpE7JVmTGBfL53+s3JTovDSA/WJOyK6hiGMrhvewLyw7cbhNoWMq/NXB2dPGahT
4GaaSoAYm6f9C+4YzRIZIq2XqSeZJx3Y/uvx+oQJ5eCGK2wHJQydlnqzlIRDJHZdoahEmhc8qIjm
GL51gUkEBANKZ24nK8hs5WXKcJvaFRTqLZCZd3P8f7XEMkQKmHg7sD+e22yH4ParvMgTEV5hjVx+
Rxc9vSsfTRDRb9nSdg6nHbFTlpE99gdK4hOXIIIOjOIPULDReojWRcYYClIorA8mtLWdT5XEauXB
W+KGoPGiZerSkft7+atCCLGtPhPEVVSOrdaj1ZAuFRzy9F/SPDVuVX8Lx5J00zL8d/Osa2CtXQE9
eJ+oLEet4RrImFm9ONzV9FZMEAk/y4TnNWEHTeE/xx/DAqqpDoHD3mYqoPol7yHdoJe/W8Pf77Ms
yEbUrr9k5mkaMCD/JoOQ5a7bnKW6YYowBJMOyumRScMNFEZQ9pBEa8YbTf4am/YQaiOVa+u9LKJJ
qZJ7xor3wvoe/5F/VKSOKD91J41B8f8SlWm+1b9JUFMlcfbJV0o/V0SmE4eDxEqxLNlj97D/uFbh
uLOftw5vgw4THiEbHkTdPAGKklIKAv9blMHwEobJ/XELs+Y+w/7yvfNRWBuireme+T/Rz+QdJ/4z
sBqjzxG4N4s7aCAMdqVSnd7E1A1UTyDMAXy8N2GPoM5AEXCdz8JawxxCfIIIFl+A0pKA6CmxBHS7
hIonH651Hyd+XoKpiu0iR6sShCjGeceCQuLgnGcFHK96A0U7+ZHdY8M2SaD11qBTSy1fgxTw54x/
ABvkEShE7zkO0sA3P/WhWwi1228ZRVxXBUh77/aHNmZKAO/BcWHsYMEpNFKMInptzqcebSlJ2uE4
iM/4mHbhhTHjR4sL/pzIDhZNP+DPHim1o7+eS5g9cLiJn4+90tp7xNikZvtn8x4zTJ8Cn5OjupH5
JlWSEgz+5hKI6JI1CVvTDSeNOIKSko8wP4jWupeaDz/4UZNGSJJfTkhMdeunqT3yrOoMulzPItbY
gn1HtDHyRkJL0M5NUlMnKRZRzJ2vMhOsCLFU5Oxbo3GjaFEZ7C4P3HFbIkJ7dpGl4XdB61TSd1hH
aTm0mDahtisab3Z2cA1uHdpSFxLgWUTCKKKmMy/iv+nHkT5s22MGzvBe8Qdu1qrgUD63C5GZHgUX
9DwTpRX5rEFJsBYJx6LlPc0gzuEWZaKllTM1YXadHVnsfsW5Ri+OIvdi5wVTuK2hvSloAxSpchtw
14AcTXYLpLLqolv0A9c4HGXJCv1UfZGzG32Z4IXOcLf4QoIPpGtYI2tYN8r5R9mnuSyW8balrt3T
Qd1iJNEdU6cKELweDoQc1g51gQytLFpNy+VMD8CkfAs1Zyw5+qwQ33y8OMHDewzfrl14EQGivHfH
S8Wo1oER/gLDsN0Ufnb0AOi04hRz/m/b4QXajLDKnBFi/4UEougdZsymOVm9f+b37W1q/s8dnGFm
tYQmjyKfuWGlNdVCAkz5ATCCPmTB7bIQsEROvcBXEHf0MhJwmQ14920RR92EudSVI12ANHS3jhKD
1/BGgGeMJkoGR2ypMtPJFWOywyVGUlyPQD42pTFz18fjbStz6ZT86gWTbxsCsColVr/zIy7A8+tE
R/ywBd7e8RDnfTG0ngi2NYQFfjBBM+Y4o4dTyoEDtaei8aTQ+gEa9MAwOMcO+gZVj2244e0fABEt
7RbgOmTd3zJy1GtRu4/XAss2Ib0SnU44WSq75UM9e9zEXdYr6ctDL7XSrHQdrEe1wjRytJEoFASr
VnGVbT8Kdq6M7jlmuWkz8QSzjrW/cFE3x8YjnKCW/5ZyE5vhIOYv7KT/MTg/7bPlFavmF9hb1uVF
zERT9N4QtAeXFtOrSocGpmcM6OE3ci+hbnSooWEXG3sdYkG7GrKwW709RJG+zyB1mEnMtAxw+4tc
cKY18UIesQAYUXIKZV9aWRFSM7H2W3ckwwitu6czcvx/w/34caQXgftYj2UxAfMYNtf/rkP0wFTG
ledPK/SUMDCYPc5CqJYBXVfLcqCZkSnkJvhg7INtbJnUC7blepwcpLziR79lel8QULiljshIGcLp
MxBBx6GXzeWD9H+ny0lZXHQwCOP5FoSsw2CF8Odm6HS+Zaf1TO11BD9OOqu1kaNOuRjcNkRvEIyU
11E2U0mAi21TR4WwCQbOwN783jQS4NpMz1bVANtwEZSsnuSsFsBQ4eyo+Oxl4VrcWOuPS0WkrpMI
dfiNxxYufRWIIq08nvk+FbxTrcFUuWR1ZKPYGqFrYebkxQM3NrSgo9CJf/b7nR7GqDCKxj3T0+f1
y2MVS31O9kCYcjl/ACyovkVryv07/8sZGf1ApzSBj4I3zt7FWbeO/tF+QOE1WJVDtkrbtSWonGeF
ef3lvfOh1RJJDcKxv1XV5ALN2c04F4xTwPJdRUmSbe2uFZsgRHgrJWbZGikqvIOaJyiZ6iQsx6LN
RGLyascz7wbEi4EVBvfNTiXT4gHnpzz7rsk1u2z/NVaNWEwb7RJdWzW8vYFyF8+beUFhIPAnrG+r
p3vkyjbRU6wbhPyT0OGcAcFDRUWxiNHZtGFTfBVNadh5fAccbtlfk4l0zmQrhzfcXqH8fe3NVbth
ik0Evu902aZanWqU0DfFLmWI0ecSKrzD13eooyahigmrzFSYoKE5uS9oW6t//iSNBXA6RNvTHZ0L
kCvjV5UFIjVoQm+Y8bf0QFffJVITVXY/PnHYh3/KO5h/qYxW1R8L82IiQOM2A7ffa6TbfsIxgklB
LXOSRkKgXVnlVVCPXrCyhW/o/kzX7W2akKEQYs13XP7+5lm2qaFoSi2D8wtmQ/Yjcie5iu4aN+3F
iASBZHuSLfuF/TiJ00bLRREyFlmEqe2QGJI2mqhAVStCX0JZVLHZfOfbU7BJSng/ixUogByFfbTn
q2SO4u2N8xuntpn9JbYdxldzwYpGHJmqGfSnVmN1qXu/XL7fqr7Vgqw2falRq9c33GKYQXDqH7Ax
SSdkqwpaQAbaAHwDlByvzedrhgvvGuFMO0MCQZhcrJWz8w3mbaDYsQXUy6LVrnwGcP5OdW1U67Lq
Mumu9sXRhZrf50vx1TPntHRgWCcL3eh8UjgJaVl2LkJ07qBPruWSr7k72OvQW5g8ca6D/1YymwNN
46tkFx2bQZujKMPF4Fx5FhRZI/P7D7m088olRC3Fw2DLvjqb0Y395YKmKDTkil1lEPUEKHfcWv1i
PD8mH06J1jSBP1DWotBvgO/bRBQ3HOWgbiVWo0GY4VYDFYiWMVF5yH2QcBpfAxn4b+FZcdFse65M
2vLM8ebJRYpr2TBD0JVJR7qLIwzYegEgTybe+UfQ/WeHwVq4DAkd2XBPjjGAzDekaC/8s2PIizPf
CKUEIgS1/ka3acnCMPhApU5W5herm944XSo7kdwH7qbdJDUAJ8iluclxXX9DtzpAcr3DI75iYuAv
xwH/Ue2B2aLirmYgtA9Z2THFFZgM0GGOjq1Z+JBA666pv2o05kgYY8R78ou2eVzX7GFUHBahkzVj
kvkXEZuiu9LvOgw2t7eyp0NOjIs/zieP4UG5vGa04lccApHVv1mBGEWUqNG3v2nJeUzLpa2ElIVN
JPS9yIR0Ti0jGKcb//fy0PXbUleXa3/qdyxFVtauXUkr5tee4STzMH3wHG4CSfJcx20+jSTYSeYq
XsCibYBOrPsxbJx02ezz1Aa4EtalV9tYNu1UikHpvPAWVZ+YbuZHCjtLTWjXkJBEYOJe+S+ybw6a
8IG3SFQWFggE6jHCS2oLq698mi9jk8z0oGyXx3IdBf6kjy3djqqZ3DgvyWGd2Xt6mlejTZlhlvpe
dHek6D0waPKRZHp3ZzyfGdRaP41cDmwcMQ8AH+fxsbOvqGL+kKNGCjdY2RQs8WNTXU7tiZa4sSyj
cbWyR7ZrPlh9O2ZyNNwjdzzkwVazrKfZFjCl9Urnl0+P/CmTfdyJva6hfsuTw6BaiVLqvTFkXjsL
hnIwVxhmZyfirTOfU8/CnC79dgckam4GNvSN+XCtZZ5/eqsRvQpx5YSWIGO+8Za5909UaKyI0+M5
ehHCRrhtz2871TitU/4AGJ73ROjSN5AVLpN9BnswGI2zE8w7zsEoqRtCsHG2gsfNVQ7liCG1hzIB
h/8VJZVcF+Lr3SWbhu8YDdmbad/MMqrzC2iA1GhsxYnE1V28OHfD+llk96fTCbgYPcBf2Eqk9uRv
YCTNXuYbLvNwUAgTcSwm0W+/pR9g5sdc9Dn1TW+1Mz0a4OKzeiGSfoU/G2OE3G48t338mk6dTwhj
LNfrH56iFuh2Ix5MBep6J9R1L6dlvYSyNmqhe1/70GeyPTX5ud+aU0efd5yvGd7ighOWnJrSDUiM
sIFygzaJPO7mufS9VQUIwo2ZVZKH8sF2p0isMIKknh/LUKTNWN7Fnm/gFfIu3IDCv2BFLNaa1rXn
TPICm7Ojuf0Di+1a/Mg9n9shC8aTVFgfaELlBeH3Kfqs4i7/lSyvjJMS3vHyh9ITsP4rqjXEoCll
XxoK52Kc0SQPWSIiNUjNANNL6zAWZqRAzaHgKgAK40O4UJSqMlTELDflYe9nT4EnA8jyL5Q272rl
I8JQI/ZikeB0tGrQkCIz5Fw7ZVE63HhoBy9qGU8WEB1DEGylv8pE60h5ZvVVIHR0YpH3BwBTh9V8
8yWGElG5kt0uGBHkfDyRWW86RjvEgyu3+VAs3Z0fAWb2F5pK0zmAe1TaXeP5dMrWzwt5LXT18qos
H3YiYE/ZU7DZ8sQV1UKIUdJ491tDKPGQS+wPqEa6YHGws9gg/0uKEynmCsbhyUpJ4V8BgbxTdTJn
3HcACy19H4J34PF7bSv38DyV8tK8vLcOa2anNdAzfGL6TvEIRvPqmqhWtgQBYUhaGX50xerKDGUx
g+a9su3TsfHoOuyQkhii7rnsdAoL6R8vQt4QltGUSTqV27eSsYEueBcd3BHP4XvxmgXJjg2zNRj2
Gzl9xyyKesz+FyVhUSczXf5qAKrbyrXBPCxXmH0ym4QUQWMabKxu35N+1QvtXcV62uuWWHQjpKH0
1qsZyxlRV+jxlbj4LEHNuQAl5EN0akUR6AL+DMFK99MfPhtqkECl047Oom6EEuhFD7z0R4/IXPpw
i0Yp8ShGLRb/K3kQT6mDFH55mbchvnoaAwfchikkyERshV/tejywfVwQq5vVlhq3LGacrLQcgvvt
cWxxnWGK13gy0JoQ+CaHO2rclurI4aflym0hSD8aFodFsqIQrSZ1Ap5zfi/KmtQNAawzgR4x1nHY
tYE6jovAwPhqH8Ctr7TkRd7QaN+MRjAv1eqvV8LUdrONUF6IJKAy6RGcOLp7IfdJn/WuBhPRl9Oq
wHZ+Sh7gTdEFC5xyVNqhseE2PKBFvxMiIYpyzP9UaQ5QooIvOY33SQBYFrbVWUhnGqIEfBjqdORR
To0fFK1QT9f+wb+G45oa/3f/gDLdl7bWanHGMsmpJc56Njp1TTOOv6hec+aMcr95nAvxiBohhnlW
cCjnQBH5iyYZQJM6HF3/tP4w1uNaeH1yqpnl0VVmc60du/xCXMaYdHILLJqQBDdgZ+12aXpnS4Sw
sj0DhHgpUyhE8ZbmG5Cyd5SIY62wy+Q6c3mTfquTNfnAkXNPUtkvsZUTKB2VQ5z4UuXKKEAFrK7u
hrxM7mvHK8/Vnd/gJQzbX2YBZbkfZCvbXvKdDcfZvnGeBmY52YGqR5W+vZiFEfQk0XQBfp/DvGnc
OUEiGqWM3on0/9nvRvfq4Mc9HMmCeZKcJselUherOW4ypvPTAfkZD1mbd7GKXmt7wxqU8077E7Y5
otboPsBAZClPvoBEYJMG3/5PxcnN5TFpMpqzcadWrep8e2VH9Iz3UYZBRQA99jM8Pe5D3aCHL785
XW+0REzakI0Vyd5Bjzsw8X8JDCd1S0hjZVV+v/0znoni2CF01veYMq8EisiSEHFbp+wBFyRivouU
FL968Xz3Tslgppnkvwaj03WTvYrftTu6Z8Dz3fm/mVpubAJUdDg1lqhrEMSPaT1dR+OL+U27a5Li
Aim3mNzHBWtx0xjqiCCmLMIf6fNTxAgS0+mjyyEXhNk8we7MWak9mFeglUJwEg7s1Ps+7RCdmCy1
VbM1tfT9OQZnyrYqTS5SQWPKoQxmpS7fC1pTeY3iRMVLA/nsWI+7HhO3uSNBSVON6+WMk7sVrekD
s458NJhFivLuLkqj9GAIgjvUndokiQeejC5+YOS0BzZYRCmJhGpJoEtIahO/MtFMxHHslLQ1brMP
qz3dTxCkuQKNVvtF82ns1suErTf+cl/uCZ5EauS/wep9Q3KJWIFjXmViuHFhl3o2sbmswiz1JiR7
ZBm8Mv98c2Jrj11snZXqzDmvLJ/okS+sgcIkDMkipnNCl4azUB0LY4I21ezaRICY9EqQ5zquY2gc
Pg9LyhW4/Y+9YUsuvg1mq7/Nq1kecqv9P9kemqlfnB+OSpTzWxNY22lq+gcSozCbtBmaQKMLR+pI
wUXHi1fLDVOdXtHsoiAx9yY+WhvZkT+GjBSjsXyOVSL4B2g+RufzDHJyRekWFBVXFtJz6Bs4y+7f
NTBuj57wDCyXVtcm/Zow/dQiq0vAK/jVVtGakGKI8nhonCqQUpcBQX2nClUv+kaJGabmJqDtuhho
vhT75tsARjEVikwxaXYMces5EmPs8/olsh+Fwv2F8exIVfatlv0PEqSGOmj7lBJdMQV5NivWvFpn
9cEgKsexJ+N1FWB69v7b2M0Cm2tJIUudFmd+cXuVPGxHgZfrdn4CGjkcTKYOJbxD9UsXXzUpXECe
NILm+l5Q4HTRNap7Po+pchBIUI98aqHdXj6qUYQLe4fKml9dgHy9aPOSZl2b7yPrK27mKSfaVDtb
cVXg7j41ict1Msb5IPwLiEHdfwQFZfAWRfS/8V5sNS8DTyfOrX9vHivHjwKZbmWOeUjyYtXlJeAO
Z3pydbI8bDPB5L5ecBCI+xI3+42DaMkbHunmDxY1NfjpNe6M0t7ZklQl5y1xiNRrBaBc1UA6lD24
5Xxx+KDBeKD4/9F4FdUt2p/SVOWf7DV/bf7De8LD3A/ZtnHGybEeTdWI9hipzBES6XNqF53nXKeR
lz93lc07lVebSgcXchukv3j4VIRdjq+pkT0iO6K4Gntg29K6sLax53hDJMhG0cxRJJgFWpJ56fTL
rurPQSryjuvZZwHZ6+oMV3hXaDTnlD9guwYZDez6FyvYdyLIZOrJdAJRD81NtJRPpelyXJ2MKSlI
Xr10VVXrSeoZGlB2lzMV9fufwWUcwg2MTgqC3OmvQ00S6tMd3Cizf0C4+99tniOOePkPfYbZtsFJ
eV3NNcLNy+S4A60VF+VzNNZpCNhfGTQiouVob9L0R2Nbp5LyyzSs/lbTSrw+9y9B/aQ0vK+Dsvor
B/EYeaOYlz1O9GxaA7UyymJHxXNcMUxs1juJTqit9IY9It2P7szXDFBgX06RLXEC6U2YF677wVPI
d4uoqdrggUw6FH8zRpPrwvlarCpLucgUE7z8vhaHgilzcTudbMFB0kikf35OZ/IcuShqWGRp9qnN
veb/AUNWNDPRvumMNGyyBDIKFPG/Su8pyzNMtmQJ6d452bcGaaZkltxl2fNIcLKQQTZ5UasSENpK
GL9cjILeEHvmyz5s3iKL2muZ4x2R91IaPlnagVLDjCB44FyR19vk3Xpp18ZK8/Cqh7sqQBElm125
BMUM7KAj0+WdVnBh1qUxYtOikGyfRDEBjClHN5GClJMcfIIppu8xpy7lOALLDyAh8Xcv0JTi9UTU
3bdonXrRtEXv/13rXL1Bm9Wlt85oyu805OXcmHKCs9F5orCOd3YjssxBK0trbXr/jaGhCjPvmJrd
J8qShd0nO7wU3UCEpdqU/udBcaQKsR5+DnBNXp3554LO8/GT0k3JQj45/WV964XRBbqCaz9CtKmP
WrWMcjiYhp/dhCLt67nn4mDWYvbqZVTxEfvYhGPNMMS5V5RjyXJWlf2MVTCsm+0MTK4DohvmIZfG
7kwWHOBucrpx2CrB62QDLlukDzoDWuCoa5yApYc9YM6PVGDszAPFGIxz+oiHklJrMrNGfIuxzUj6
lZzwo95/4UAe4My7ZxYD5AYZncCTmFcCzgl/2PdjqpL8vKnz9LZfYmduXA10BubdyvcDuY2vJ9H5
M+bYHQRK5UmLEzIbSwPOLt4iiN/Bn+whXu8XOLs3z21fngtdbaO2yscR29O5XIe6XfjwxJBiC3NP
16lklebEsliaw29/zV02d7MRTiW4Z7WpyhcwjYgbDLnn5MO3oHS1JQ+H3jc1FW8jLIbRh51KROS1
si+7LYGQFsGOevaRxEAU3UOoWOzCYW7vAMBHO2Yws7iLrAvldKym3/P9FN78qrTD68fvUULbcncy
pPIVYSG29BV9J/RQud0VtU/Cp1bcGLcJD7w3DvJK1hROEIXhcyGIS70/5qoXWq7B0W2h4cb2Jhrd
TPFRGVUiI+/5/OWus7tchaPnrUMNiF7HMgqV4j6K1+lAWuJTYNeBamRMpBaB6EWP9UIu6UdnSbFF
z3+o1obUn4bnjbIWdSWAA5OpVyOioCBFz9ouvmJ0O7aVN9i8mSB5ShZYePqRTwNPg+m7LNdv1r6x
K9bkOEKW+3pTovlzyXaki8aVtlCy9nDMCd68aF/QGn4CTVSyoKjNL6QF1SvdLO43kQnnwcX1jkDc
I83C1XgiT3aTDKAlrWso1QNrIIYx5LCfHwWI3maA2K74YdMeIXvmB5t8RIxmXntz9m5GUEmMO9Hr
gaXyqFpL1slYIrDb/sSWLF9hgvCc8gsSuXt6+5qQtHP8wGmdWgvpjfHP+g+S5i4voCH0C04GiAvi
zkf0/OC3nH4wrYqIxO0lrr6FKd3P9cbVhSIbWeLz0gaLn4Z+jpTmLyc6zs4CUxj19aamUI+lrC2E
DSO4+o2DwMT6eR2p2eqbijhOLDKhZ2NoUfbN+QSDRDYa/5FyBHK/ff8plJCMjnWn3XTZA9LBXkfg
aJcAoLZwmruS9NyTrzpoZzYGSmuuxcN80brIdiI/wWaVfHvIsxfFwh7HRkze7NGWfIF1wU5vYk9x
VSZ+MtQzpCYZzssNEr2hvXmC24d60jqLgpLE4KQuA4mHwQph0PI2qMCVI+jYod5X60YGjkTuonHD
1psjPgvMsij+OLNkYAjfe6WI7EFMLJLzATeDMcAAFn7gGgECNPLZfmNXjoBEREDSvtog8qKFiin/
n1Ihl6W68vFScB+kzX3mfXhIXWBg7ZW9oDUwxsK27hBoWsWUhkjX7PJMRDEoPcFaj2saOSrWNpZv
HnjvYEQDXaGmimT8RFd66Nsxzbyq33qLl4qwK3a2ffIfzmSkOPN6qLnaEkJ/4khTcLBRPvznA7Kx
uEwXguy/VjTpKreWLsq4fRfOG9lSi3+zgtQUFO06rBjLFucRmP4yxhTy1IAlD83pg7R2TiDmbeeN
v+iD+ZWJsoqp4cP7B0hl4pRWxqByWpKjwWO55/3QaIbHDb3jrnT7thWZK3McdToOSrsePsQmrJYi
CWiUE9cXRgyeFtgqmPxboN/YOVR2/hw7UmARhBRIZ8C0eG8p7iPudZxdj2M8HzdoGGhP7AqUNhIS
CQTIQQgaFQDgcQgE+uh2/L3WEW/Y27KoJED+48L11DJXJpZGA0RH7D3yigmQzPFpVfkNMHaH39vm
ZjpJa5PKSrpfqlwsdJhLCzvO90LIxRPb3ImgRARh0woFxbbjKrLbhY6QATzrm+J5kTJeSCUt+L5Y
KXPQbUhw426dd0Hqhs/v58KNWvIDNWZg/WdzHtPpzHMbZKbzEy0DKrElXsBi7INui26eeug61U8C
m95oTQJQA77c1+oTAlqOs/FGP8kVQhrva+x0qhU0SdzaxvcKe0aoAQVq4Lc3eCxWu/l1dOsz0jXl
kAcbcpMufSAMGHHyuvI6bYbs8u/I32BfO1YWXg00vlz4d5Bi8z6ZcgZhbLCBfTIOKu1uCvQUkQk0
nVVuQNEDlhtyQrVy4bt/zkYuJ97VB5msuihD0EiexiJQp1Jl2CbprJWRcSWQP+AL8Lfne1bJSNIB
UzCnQ1Jof9Agw7CpcL/OHXv/s0U/X18cc8GOF1xUNhHIeJiVahtKwVn5URP316bxARQOvDisD+tt
YUXLN/6oZi5fAXkFD8IWIFbP2UZXuUzhZ0XOzB1tYySV9YID9JoAb/ZFTH9TvtvohxsESRmUDjox
Q0eea4BPuDx0CjoOPb37f4hIJ2nC/tuaRFQEiHtKObUyBy31cCeVatsa4szXodHQ2iIxkrLozzjD
9/4TFungMDhipTqqKp3sY2hMgJoi7YvrWadwatofgzvFVTKDrpHO/RnJRKnwrYhuLJT3aDG8zwxU
x7PUds0x3S47zeu7Y7reTJnPd9/2Q4KXdoHdoG+SocgbRMpga4Mzo0JZiZwGNlXcwAMpTvGzkNr/
Q0TUyHiE6/9iYcXVaFVja3OsGscXLVAvExm3XMufTn6RUIdZtW355TO2LewvysxTs+RollJBpnKM
WfVImf1oEZFECqgjAD5MmcNNfT/Zgx1ZDB+FWwDSV4wcuzsp/LlVu7A4/t8L20c0znhrqcQij9R+
CEL+U4l6fi/D5EPjRoXzFpDFK3d0BZHueia1jhCHNNI7M+7VVWOBvHH7fjm3ZVGVQK8kZZOYT5H5
UOHl9iDsTpydHXbVrViPb5/08B3yH9m7exmZB0gQX/mUYNb3RLlCQ6SbLjfuWm5L8NuTScySMzyl
7IJ15uohSq1ZCRghGTUawwRPWBzrAQ7RyXVRNOOGuBzi1WbmSa2amsy1kXeKjnlqowwBgU2dtU8y
38PR22DTRvPSXNUSk3cEObNO8mtvDiP6VE9aj0dyr6GhQXIicT8XnFahmrjWrfhUAHI87ZRAFyEc
SKGIbmlXN0qEkfHHJOBLil93qhk3jZFPXTRcWm+/kP5TGtq9js7+AQSd3rlqQtxRlKP96RI/Z4gL
vOsCuRjYYrZ2pg/xBVOZtdF1o7hxD/f/f5VNwl4IZBUfqFFwe+2B2mph09/gNukpEgC7UuBlS/OM
lbOgcuwKk9n2dddaOZIyiI+IgCfEMgBXg7EElZPi5V7s302lcnEdd5gTJcYDsibJzW5EDD465rBf
fgzFxnj9JLuozSGOX9YdgDfqZz6qxVwRVBaOZGDLN6xUAFXWXJV+JM1r1yppK6ekzFy10fn2dOeC
pxYBtz4a+PDC3OzepIRv3eRqkfAlOsytHzI6xGDM0H9dg/+Ee6NaqKTtHk3dAuuuuUnqO3wsGZ6n
UnP3bDklbOnSj7HhuTTBRlKwICM235kT7GvjZfTsNExse5bx/uXMC8KCVtzIDIpKgnK+YGunE2+1
OWwO0sW//Xfm3NydU1pbyzA6beOEYeE7F00GBBQRqyP7xE+6fA3ZeO2zkQRZCFLMNEin54Y0Mzyq
wRivGd6ljzP6enI3h/wjDptbDGn4Omn2LHWR02f9gAAWv/fDie/vXDOJ4xrbQRKQQlEL+TPOZ7B+
CUjuSUlD/E5m20nXbIffCaVBIreXu29WkTUQDYqgs6tGQYgpT+tnLLPoA0LasHDz4a+FrcmtD/Ix
tXXZOumgcB7IXUlOwomRRVQEmoYEPfCnzcfDIOUHs82qtgktmT/bnALuzyjIvNqMZdNz0xapj1VS
Cx4vhmqvrw3WOqC+gRxw0pG4q115AZdo+E++ioTLrUpas9hqDbQeUXiZHuQUtwypSvIkPSm8PtwR
L7tj2pi09hXSq9UWaw71duvmEvn7d/m6W+Vxr4nLLI8W5UAxLjZ/aoBb74fbIlrvvqyHysAdIzyc
Xxop5dDVTUaNWzlnKoqi8/wVjoQYgV8MucsFM85vrVx0wKKQYqlomc8aoanaDv8RnVGgOLmc5+vb
hVj0p/dbdZ9C/JPQspXI3Hu6OIMNuWOyFfTp5Wxin0KMTF4WSAV+VgMyKka2uSdkhhG4mcgBheyK
8bGxqOHdshDpAGq3dPfIS7+5Y9S0XSFtKgxGfx2XAFXYY4tGT8A0lAPH7xgpwZVYVG74OscXTSw9
e6ga57xE0Vwj/5pv3QhVisqc4yqegjlfjxozXyUs8Hg+kCzSI80Y8dI8ySzXRNNJ50yh4DKAIlHV
xBcAZKyCb2l1ssA4pA2dxnrBRoIIbBYBX7grYcQR1XuVdqqpH3cPBKVRPHoCh6BOfiN5krea6PC6
RuIuhPyIVbFimDhLoLFplC/WPA1aZk3N61l2Xk5PUdSY0hGZFMEF2QlM6lndCnYQGqhWRIiAIm1M
TLPHfiYYOs5C/JD8vFYnX+5tLKQfQZBrIFuLdzcNVDMqIGYlH24lpQAd7oN7DEH4TawVMzAdHEe0
Ns1V7QvYG1lHOE2k4rTxKbGJ5Cm4DOwChWW3koNbuJR+RhSL0NhMgG4VyF0pSybr0UE9gmeNTJ0s
NxSo5uR2MurRX78F3s/jgGrCiSWwBhYTS0LRjY8/cgOTMOrdmBBXdnJUKf2gbD+fkEmW71tlh9jY
aYY9RLXmJZTLNukVacEJm0C5zaZrkyWC4KAomcDq528KTrf2KywUcu3J0oBF2VwPxHSBBIUcHjbG
AmDo8ziRxWKPGyhZOAUzrxMOVcJ3eSAENbV0lg3Amx0R7u/pM+mrkUHeV8b8nkLQeq2DphLRwWYP
t/WTUOSwuBwYwufxjOxSFYFWEn9Kh+sUldzWu+3Uq7EACu58s0DkxtR2QxTHLxLkebdGsjbaBTFI
y4RYnCycU1jnWkFWTDN+JNj8WyexaELca8BXGvfnb9HmUVm2NO1GI2ACi1j8fnTmzMN4N4rRr135
GiGJlfe7xl8XhSQViLsIRdF3GLGz5rff+aIL1Ocum4+mM8XIs+HqOU303YNTsCyzRW/l0f+vuH3R
VwjYo+tBzQZe8GE+1VJ+QWDWBXYkkg4+a0bQWlNmgf4Nxb0ZNwBNvj1aKVdjO9f/MdozSSZdy+CQ
DDt5MZaemIMGC5CTIN2CASRfXSvNeOUaTFsdSGfQzT87ZLPkEBbs6LUHEZj+4Z3p2QutV3d2jbD0
EbMhRhONi6I+shgU+G6Qekvk+swfToHi6Zh0bRUai3hNipzlEyw/uDeaYmtlX2a1Wk/tZmlg6nHW
JIODTRTuHjrUX2qk1FcL+9K8XfDgRRCX6OoLL1Th+oMCxEYSVjDAMutAsWQ3ejgL9QzuQrSok/9v
GNldhgiMGnDOsI5zcoDpOfc3F+hHteOL2r2Bny2g1ODLDAG+i5ZqcosLsuZL1ycrWdLY58QeXz8h
xhIhlYW7KDoQRyl3OTcryMQmDevnm/KUQJIx68/WVSrCFZxHW64r1ddzHNG2zTOG6U/XB19cz2LX
y4CQhtVD3dvNaE6CLgdabnRzVRFxwHX/HkTVymKclivG0hNt8gdie1X2Dxug2Q7ZwpwyW5GmWb61
4raFDF3tMoHgOtJdMGmKjv0ZDRbt8suGLdsiLVRWS/mf12ZPOd8D8nRch7z68n2G6zXWA29pK5iH
rpTe/3cOT4RMQgJAdd1hALzANUVzGHC7kxWra3wkjACAAgLQNbRsAdFIRCBP+TNPCabB3SDb1FcE
b8Y4vjZWvasCwTpQoW803C0A3Dj19u/9gyPgPzyNyjraO4qBhEDruRO0VTl6SdpTwZI74P0cCHy4
s7uBST6au8laUyU7CceNBXcQ/hXiEVPIjMqZtpDbWx2ALepwRUlbxvUFbm7f7+ZoX9y7K4tSciQc
MH43g1i/lIVXRfrUBf9UgYt/eaCEu4+2ZT2gBkyUUJ4kkBYzmLfrZBETdzVTZw2zVVBHePhXtJIc
CWt0AoO4k2B7s+TJHE+1jmNEZ/og734JThiWlx70vDfq5xSwAx5cvdq5PBRuG+egV2Bctt3DYkH1
K9KZU72KUMFpyLUKjh64rKPQ1Mtfr/4OOAtZhjNs3eFgfXjxFWIonatw2w1nQJBanVxjtgpMFf+f
XLmK7McJUSDm7+tc8cKILk1iL6xeBteF/P0mSpo9zVqcBxwiORgj/56Gf6KDd+qTIJ9ktOZQiLg4
+g8uXVFcy2dWyRT9PTTQHZLGvyKDyxi+ENWLM5tDzZ/jqZAs1GWHwdnfxcx87Y0upioiP/HqxV8d
4anzm6HBJn6Z9TAGp6jynsea9TOkHGh2P3NClGlTdQWNXJtdR5sUV/XkhGSei/NJjfRBVGRCDRe1
/QmYsDOeYhl65TcG+m2Xgz8UDC/5zF+bwC99a6NGHC+IEW+BQqWL79rBGIEiJFeIp9MuhL6COg8l
85vMHcpx4V/8kAih5fe67WXiBwrgzwUXooYFr5f8Ym/nC2FKtdDrx21//zHOQ8QUUrvD+r3HboMU
IvSFHN9ENzYdQ46BNKvqPWrbh5kgXPp5bVHFeQAWgcrOxUPVxNnpU9XjkqEII95M3FJUBkoFZayn
epXDmYdxtcZH5gWEymDPBTQNopiy1Rx5mHwguxhReq1Z1mUdnceiML0iwkl0hqBaq6cTbfwIgfnE
PuftMPaDh6rgo9A7FBYiaBd01mlS/KDPkhhI9DMhxQpA6lXVZPfb0anEkIVHvPg9zZPvrbnPaWB4
Wuj2WGAWfOMqyQCMytpdYcLLvwK2y0yx78kBRNf+svAxfPUCA095oyomtJwJhEZv/LKyvJ+O2oGN
sJe9L7Y4vIxcsrJIsFmepJKZI2FQEw1V6WCo7bdxTW+m1QrqxbHTi2adukWqfY0ae9F/iAXncp+B
8XXIYW+1PpZpWSywQH89HZNWmPF8iY2KwtHsugwXdYyUrnUa/0WzEradOVT44tjhP8h6Fp6Akp5Q
l/lnEFcVadEgEsDWb1r48fxYXAb6r/8rDGjeSvx/Jm5qVZxXP8yNZPVkE4RpFxylMcYDxsZX/2BN
oILarfL2VBJOzfpXfU/gOjek+nKUwlBxt1ciYpUYMRSq+DU+hmrv6PcaBEBK8xTqvsi2paNYVM+Z
e+9qDbdiFVaICpfEJ87BlK470EcuLp4yJpsbyZpMkLrR0eLnh7avjm0tFDF5i/XYixZdwVn8yMwy
/R345P6OdWusHhWIB3oq/QSOMtNSwV9Tyc+A0RX4Rw2sfvd2gc3IwO3B+VHsfSyZwYxVdgpiYFp8
CyDeo0wpi/LVGiiGpJEGDiu+8/SdCsX+EyLwRfJCqiHYF9I4nDsDY6dxvmrr7+VlOKFtv6x5RByQ
ELifLwyFV9T1pHkSIK2pJ/OMF/aRJJK8IaXRvRhNUKZziuNiYvb/HwMvpVfW64UCLiQu7Gt+XNoB
nT3wFw4ppn0iRURrfkPA9VwIE2LowdT1vznphaumSXP/6cuVVirjknY3HQDzjihz74/3fT7IlasV
VZmILl4HHDG0xcud31Yqv8RAjIWRjLs4Jcdnd/BP3bIM4G3AIJOaM4qnJXwwAkfJVGlq07m13VY4
2XPMUDefqLxzSPD5C6xAV7BZU9neZxMXtN5nd1AlkvCct54qBL/baidwpM0U9rhiqKWUBpkW2sCJ
Za5RKuWTv3sjBocjutfWcUs5Mw4AJdzPmWjAxNPQK8I0mcGrsGqVLWyxFhS6Y75r31uAfbHipHq+
5yB2lHywV9NedSiQzGXlJ6Gp2+a5+Dg9V3XwCzxoroYnSJ33J+kUJWI+1kRZwR1hsSYEAvNaVHOh
ERnh1H6MoIgFGBFBNUUq42FMoByRVwh+2GCTTuRYKQj6NwH7KF6GIUnNWL0tFSKNAM4U6bvPNB22
ykKX3JhjWjQHFnueluM4KIuLR0WtTQuyHZXEtxQTEErWKp5S5qZqoHvcUhTX1bvkT0j+WwO0sGrd
cum6WlmzEw3I7qdlpCfReIkV+nIzFhk1jPynX5yTOJd6nppe0KfIWhFMxyXUM6TkIhHiPII9rhA1
zBAA70FwcR1lfsRawEjePQ+vyoxazlix6bnCnj4LNjwvpY89p2VxAtF1UXVjaBQBPzrzqsFb332s
bO7y3mu/DuMd2/3BWDSC8p5VsVfX3Th4cd7O5/0Knmlr6uFzGb+OdkWRfKvch2QPotQ6cKJv2Ook
e1Lp7PuBtxBythJ4cmbORHEyLbbNHAIg5uYTiUo+Q6GVqBYNy6160awCAgMLyuqV/f6ZqBXHfY6a
hn2msKSTdcbgzRQp/i3k7caYAxZ9y4Og3URPmQuRIR+USmTFQ241x0fekRVulbikForliye2YE7r
OYjvtonwETHTEJ8TZ2JTxZ1Noct4fm7/t3rZOYyb3pJfe0ZqDEMcRmTxipBtIAUWY4OuLtpEYDrH
boSRSeitps18x+Kh6em2azE2u3ao1lo2VvJXL8Mt4PuklRSQYqxeJnv6ytSI8LLffntxC/04vm/H
os8ejNf2lBbeljFSsBg9UNBAGHKNKWhtR7A1UJsW5GW2iCsFwdMBB0tQX47K0BrsL2/nZDqA9G7R
45hs6Xz04z/rem1Qs2eCO9YKHGIwFKz67+1HjTyItn8GDESWsZdwMjFmCEFZDqov7c/gf/Jamk5v
AobWnvRd89KpWDen5zLkMNr/p30t2woJD/IZMS7jPembiTmIYP4feM9tEgX77qSa+XKxTx8xTZht
KB/klKWzNkziqMk7vKJuxakf7xPLNjhoFV1LmoBAYwrOukFO7GWKJzoJq8m1yV1J674X675m+g3u
08ftg3/Wv6TNrj+EA+PJ6RIofdj6R53QCKk9t3JkmJgtEJq2wxPxGw5lqhGr1GvWILybrz1JQVUb
LmDqUVNfMH1eA0P7qrrB2AzqjAwAaBemuiNt1HbE+8BwrHhqQ5ojq8lzItts6pHtO0wTSvpaD6X6
+0dRkkCNsEWP6381tXNOQq/n1BbC2zWbV81amdQO7w9ptwZwDVKrWxHrhCX5brGaqbZmhM21cFHL
QA7eBlefJACuJT8gR9GUvFnk4b3KbkfiZNhMZqrVqPV9x/a8nTJ+UTvakpaeUVZ8OQ6wLvg2c96r
oMtpfagHYNH2dL6a3IWiZQPh30PMMcJSHvQjPlp6gCv92snhmlljbP43rXUtG+5y6nbdoYwRKBJ+
WGzDDOjHNab2I+mkY9GCmmPVaKzjfqR7nFrywKodj8wk2RW4MpXE881LSjp5RGUGiLgpExo/Os+A
nEvJa7ztYBxDjdk7RrohHsVgu9P9/ykVMJ5Q1l2fG6dlyVy+aI9lVb1hpIAzSHbZhHiNznqdLDuT
7XQbu739GNXLthreZxIgPVD+MD9da4XUoVCvdxBum1w4AghMZZ1VlByaVU/DRDi3ATnZ98Ev+Um7
qrRwu5EwplKe339hWI480MwQ/qA8CjGPOTizkdUoot8qU4skrq2pQ6XRLciEEFhF4odQYXRM2f1B
q/h6CSVMEmBCqw+CGB9il5azGIYa/vF0JwJ44ed9ZXlor8f47v2tgwjiTfmC+4gHt6lskLMTHq7J
QzZoC/qdGiYMNnxYqV83soADGSQh0f7ICRr7ix7y7CjpqRgMcfrxbGHRGeSCvF8vd6HW7aBuZXGL
Yaj1m4NHlmTFyo7gM9NWmlPrrRPpLO7Dlc7tBAZli48qKvw3m6Vr8DeFYOq3AcWrIo/7OiQt6mo2
mRiNY73I+fA/6UQo/NHp8Dw9NocBk4e9B4lQ3xGgg+uSWbT4ufvc+7Y2wjoYT61Pgrb9K2xtzswb
ScGSj8t8CkVWZbQ72QWg8HwK9MDl792nldhxjzLqSJ+isWI6pG0GDxMBSu41xbTHhN65kDUopTiF
GaLFGGgzWs3ZosIlkDw8ekYeK8l+HqRxz7PwDIh7iI4KB86Kd5+Culk9OejLFMrkax2ZTx/5qtBS
nA/VvRrfXspZ+XUyUiIRbmk5xQ6vdszSWsq0lAzDtpItPYqNZHMTCutM+vJbcLb2XlLO3sMom2qs
8XFJNc9olw58bCaz1FVUHgRzOJfNmcKLVfBBf5uUxXmIaCp0oRDxYYY3yioNyXld8mJQiaTceT5+
HbU2RmHin9dGRrJCDS7Ru9U4Kpo05bJ24/xqe70yeIWv2CSd77c+13ZPm3MsdEGV4fIIdkaDAiih
pKS/CYxlOpK3z7NJjYaQJ/oAIddP2CHlQ9lgY0apsz05Tyx/v0sdckOzTRVTLnRBZn64rbt6rwBQ
h/FmPK96zhE6Vm4YxksTB8eG3zOURwcqKDo9DC+qV0xoRi3ApnmyzgUHbDBteLwG/6DqaIYWCMt0
l8Y89JFIQOW5j3l5Qu/TFOQKxNypsBzJoJ4wnMxuAehvtSjjEP4LwNdLaJdr1qFTHfDIGpv8Wpv/
mXJWJKvwA4wn2YGt4CjVpPVkoCgbYcZqi49R6gNv+MyzIjUeREtxi1P+67ZNwgB/dQoKhyYk6smr
jxXA2xbSdJCwwH0/zLyc5UHigUqZbPVk9JqNy5Ls+mQcKVoORuk1ONpFT/aMkXTu0av4qldaRGv1
B0rysdHD+ak7P2wGAT30clXqKXXHVLmW7Oo74L5Yf9wV4MCudSa4ieAYnEoHsGPzLBogi7LbIgBU
CxXyAlzeH+LFspGNpj7oJha5rNv09xlrTYT15KYw59lym+VZeQPRzVo2s2L/QDpz1/pADb9Ophc5
0NPTWjyPttDrbel1VmAAGeuszIG3ajZ+3+hWEKeHcTYpVuq83oxsOnH89GWBI6AlArEE01pQ4BsT
e6vtxiNAh2ypD8KCXLYtpUGO6NRN4GlPJ8IQ4LuI13XfyaRp4/zn0knFTKhD4jxUAx8A8tTTvSkP
BWHQNJH8GV1/afu76xTXJIzt83frQryIeN3fr2APSoESChiS0kQ1h7lbD4ikQ0tzL2ARH/1iGLWG
XcswdsbSXqvUn8D6RNesP4k2/2qOvGZL8zwMQKf+BCjnxH+boLBEoLPhGloL3uCIR83RFhOp3GTd
UzOpfJ8bhThWahCbJaUQRjTt7LujNBcgyEx6/8Lm75PDRWX9H+a0dsOIaeb8iAZjrP4t+4jEANo5
qJbj45nRNsht7zld8By9QF8C9eH0XPwGrQO7HEDt9Qy99+JrZ5QsW3qe9Z0duz3X6H08JzSCKSo5
GEIueOZFC+4dczMil269tWr+EnTnWa4GDfDs2td6esig0PyifCKFIiKJQCKigHsowTJE+qAqZUyl
T92+6AKEESJwq29qEX8l9tozI1VFJxpdMcaU9NuD4Rio6zJfkKQmuseCduvq4pIDhHea3QnHeLPa
VGNmYP/8Iht1/61CbWLV+Wf+0UNCDsEglYEFf7AHNSkTfOqzBrNsnucRi8HHp2yo2/d5jGsjw3/0
zyKgcUamF9193yRWoT7ojBvE8csScpzBnuqE8vwqwWxnCK/ouS5PVak7DlzIDwbqYSKk6TllZALO
HLEE9qkoj4/QMTVjXsFtahOojYlUNAiKQTgaX8l9r8FO1dk6F2q1UfKsdWbSpPtUU/IojYM7qPsZ
x/VE2KCWbpSi/SsWoJ2mmzTTRktB0Fsciq0zLmLoUrgFfC1oymp4bDWNgxi/4KpFtObt03OTfSuD
AW7aODL93fmniaSyqhCwiEWnRaz0EHQyxrKjtXxDC8lkSqxzcl8VGPOZAl2elj3ojQ6876j7xc+V
xXHl7cwXy/BHpoTFbqGfwiOQTPXYDsuI4SJLKtkuiz0h+Ff83bgz4TuC4uDLqRk8MjwlCpGC1Hz8
9NbIIWZnq7li6arCCjSsfPBiFoZpTEQzX0SY5AbkyUQrhQgNWwMET7fKVh3jh0LTg16j2qkuHL50
Wfnj7VVz8VQuvJLdv5fIOwSS+L4mi8Se8WxB/2BUZNnSofm8W7e4zXKowsqjmEIahKX1/JK1V1m/
aqwb5WOevu+GnKvHrHnDDrsIXpSEft/FbV/mlFmvJIfDK25L/u4LXeJ7y6iw2TeKVwiqsfAOev4N
4uvC28YjA5rJrdTDrDgnCKJLpHcdSW04WXs2vc0hlVGPakaAJFDoaKHVCDw66AjMJSNK/Uhjwjki
muRrjgRI3O2A9w3aTwETAfHA6b/zJe4UuLPsOywjRPbvvDcXNT9P+4l3FTMOlbKu4d23SRik62ke
TAr3DKm2QBk576/sH1ATv/SWH82knWBTV4PrdovbkaLyf1aK+XZcNAo0XCn/QW3/znqeDey+JsoT
bT6g5H/wZPPnSElJ9pPQtH/rbvVxjm+3loflriqPXxXZhEd+FEUb0MjANlxnJ8gooB8BnLqcxyAg
lGWNh/RSf4ufcEWxJ5oWqVlPLe4peQntcsnF+4e8z+GZU7zCaRMMqj2auDWf/pxw+YHHbQH+BoZt
2+s1kk4nQQDPL7UkTIFHX2HgFD+YAARSaQCcOQraLkbi83XKeZT74Zyfm0bJjs2thFAGr4VW955D
7H+b9FY54AlboarO3zkIn61eURtSsfBQCZmEV1znQSaUX93gZLg2pIWjgScqBjamChQMJ99b0o8S
jL+J0G3RFoody16pk7aLZlf2FsQlupWmGZ3irEM8wbBa1Yte9KBnVRb/vZwbS870g1HHYfXGupIk
yZVoSh4iJG+c+zWTapJ9si69ecnMWAPoYff7KzryIsOBoVJWFV56VFNrtHszwumAiNlbaUzAmMWH
6mco8zhR77rufXcJQ60QvvY5tsjcQqMRjUa/t7XUfsOtyBd7qeal+uxyc4uOK1bcX5X2RqekISOI
Cy+vdZyuWEj9F/x3YNk2CuCJxG3x+DCtA90+PkXU5dhjODs/vT34unvE0uYclPF4/KqqdvLpOAw3
7z/9yXI+Lkl/gux0E+n96IN/MvE10Y/exu1bDn/2ks3oblcFk2hxhCh4MQH976oD86yvU1vDUcR1
g8D8nKfgVtbDww9Z3fTZlQqABq9F/ptPEj6Gd0bmGfSHo3h3axK74HfBb1AUvb1tt2FsWYSv+zjf
Qd1vnAMIV6kqjCnCAfDk6wFWO08Pazqm4T+hIZ7oI+cDAni5UZgPdIeMGSEbkO62pIVIhhjhMYRf
EGZ+0w/WPdmNVbHPf3DpqRN+94wa3YkzZyxQMJvtIT3mhZW2LlQROz61UAiSkb0yI1gb6uXhEMVQ
/Ux62s3cwoEHXsOEF9eL0gNrP7pO6WzdYGpd3nsfgJEOar3G2Vso1P0rL1Pc03/2nxuLPrVhiuLT
vD+ZtX7AWiAwq4s01YDkRE/M1QPip2DIfQNKXlUukgWP6wmQgoOiSLw9q9HfH0Y1E6z4fQkp28Qi
DlsMMldFg+XHkvC35ZaBbVMCOpsfRpuhSmWwFHbFSoegM312AR2tkrPy2F2cqjj6DPHtlTyYMTZZ
zkRY15LJeA2zb91iv4kcm4HgWYmVYS1IrZA69D0JInPXdxx6EgL7biZkYMU+fKLRq9vbgPtN2FZk
E7rgF5MSxsamAGm395CBkCxr7hO4TAG9z+xfblokJOABfiqIrUaSf8Zg5FaG6NQezMfJpfjrt3s8
k4aB9oUpkiaXaFBFmvOEMbi89ojzNvkkjKIAlLtaulKgEr48zvae4L6XgnAZRCVi9nv6Ce4N3E1/
9rdlmBffBpeRyoJyG+keyOcTrld8Edxj0Bux9UBiYCzH5Hh7n/RCOWT0wFYIb51A5GijHDzaA23x
AFpFxc2v2AV2di9CE5+QiY8JnApq2ibJa24anj47O2/f/mOMcqy9KFulW+WZYVK8001oET727OGd
Ho4qN5hqj3YzLUz3AagQLUH6t9JJf2UQ8T5Ed+veGxa3asMW3oqKkbRTVZTAGwGGiXsTFCY0jFKL
P3Gx0xI3ITVx1THXqkwADqsrWaneDNpCflJiemqYIIPzhCcLgo0zj0UXD1VkqtOIsR33iXebs/R1
EnZlHRjRgCAjk9l/dvsI3gmyHb4y8X4V3nviI02SAQGDKjwTt3NUgEW5dO+FetXbuyaJcNbOJaBc
NHq29619kXDQRQAZHE4NzoHaU32AdtGf9GY+9L8Oj2NBjW/h1tM5/WfqxUp5aPq9jPQJ9mgRJuV1
++7UZrWW1iASwNSWXlLS3tZMjL0CPIvlk2+0bTjhhQC1hLLFB3S2+v4k4ZPngtG4omg+PZqRDSwy
9+/9nrQVlWDPhAdo/4N5NkxpteHp+gb5cJ6yBXr3G5VQaj3iXQtLsmibZxVjjDVaOFwL0RxVBT2L
wZ7Fdi8sYmKeYUWhvjkvM5xHd0Xq5WCC0fhKLJc7nXuA2ssIWAZY6yPvl3GowBdFCUuW7EfPCwSN
czQAmhAQ+hCynvZwfJchEorWNHPyHHcmE5ppcsVnBLRYwJCe7azaOC6FkzJauYlUoKGOsuXzyGLE
xElt381VHDVja9hCPYzqQKHxNbiVvaxeorPcv6eZWbb680q0dSoTrBVRGAlPwKRv81MFJb/Aly4e
SgISuu9QmkKLu5Q5aCQ46OUHC1isWeLLvGpOoHaXR0r471VM+OQgYIQ1aXBuknaGBpaGJOxS/in1
CSs19iqwMkxIm61gjupMHadHYoIjLx8sRsd0Z/OC47d4qdUdLOSA39i0jxt5GfylbtuQCkoPGeZV
gSL+Xjyod870tM1vBigR3Q3oN1VuQpvEV7J9E9hmJIYr9X+yX3/YIGgF9ttNZsQTLgpg5QcBhZ4j
ghUqeDSRtJyOH1yCuVt3/dVTYXZV7jL1/1g/u+OsR21XC4kGP/7Q5oiikhWnsnzOvMaj1VOfPB/i
zOzoV6qTvA3wwQg0N3/0nGoimhh4iB/gSgYD/Fg1jQH6x8drX4fBBnB3bUVjMhy+ncwKTWlqKV7e
mnfEvkm4qYmNEffjOlqY8z1TBKaJkVKgxePEow+YXRQkZ3xxPv8+MrnxtXJhzABW+cRR3L/4qlBL
+17+H/qiliy9cOtcFFf1+EElvUbNlRrM2HGJctiChuHzEugNO3Rek6crApcC96OQBzEREYgKZjjL
x1qpN2yhM3K0PuEBBtQFaz6WXSRsEHr1/rOKlKal+GTgoH51dW2E3+Xioa+NlyqNOKxUyifAEfvH
KZFkQt0id4dw/kLTNXJfD2OIgl/CdT9cPeFa94NzI/M4e+e0c0NnaybeI85GNwFzeCbCBwVcHyZE
Tn2ctzpnwn7lqJeorSLI5Vqly9C5vRyqlNUd9aDsNjBJEeKqyXxI6qYA9fHhap7YB11jqdB3YHMI
DuHm5CgpCR9zgsMEiAEDZmBm91xELUmeVIn8BmhfwSlGQgBszRkbSAp66gfevmfaVHE6yMjiZ7VE
Qe8nSyWHVwpOj+HhxbaP0+GHRTVQVr6EfUszCe0vQ1RbAE54gpwu+pQRQARBtCcHpkWqjnRO61dG
85/nwuVHroCW9iAGw4Z9GDqvXElFPSeX0jMOuMK48XTSJRta5N1RcvZfgxxxHQxUnQdftZf3Ow03
eUJR+ggfGqZYtIeq6m26dhEKTEfAe73BEp4zSDBcFfCMzFjZlzUMN23ZJAkE0x2LJF7kzipT5LEI
gTdolakKnN2AtfkOgr4xrP/tGkfy6KSQsPsNmzUlr9U8f4JGcT8LKmOPYBR/syaki/wYmiUjsuj6
tD7dIMZCLzKPq26x1FcTqHnnQsqWayBS0mXmmh4SRDXAJjFY/gwwVZnhhp+B0MC6sZQHlcdjQuZb
KQ7hr2jqVieo4g5B4jeTrc2IeBPURbhjCqu0o3AKsFaRxmhCiOZVqYmvcxq6eJphEKo+CYqNdaKs
YYL2VIN5NQrRW4K5V2BW0F20N5yQjVr2MdjQ7927Ckpfvvp/U1cos8Eirr5gmcBqNrCqLXqNU5J6
1cE/dZco+EPmJQZS4u7n7OJaKYIlxt/NpbHdTshOOtbCPkbT6EJUn+8Ooe1zgRearz+EC+poYcqc
L7KOKe6dTrsmky8o4T3r2t/xmPP+STRfQLsaACWMMh5wHPjqInolLsHKExlMHCGKG55ZKjmc1Ve8
xe0l7ctOKZXw0D2lE+Py8cmSxeESo1ik9TaAUQ0+IvPFrCJ8SLfwl5IVBHvJstZ6ckBhlWEx7X5y
x8+AxMlp23N7D8MdmY2rIEMBB89Y7Tr41kW3HmVV769JsKmfAgIyjHyqhC7jnvbf/h2tKVTPtBCw
2xh2Nz074p6exJJjURbIo4oDc4k7VnB2eO+XmNoMYpnGfCecIx3at5yYSoE2xHZk3tT2MPx/5iaG
XD9cxlnPY20vwmxUh6488+L6DsNop+EvJsXOCEdY6qtWVQFV/cQWRwv3+dm+qWLz7a4ez6Dk9Iph
i/3FH7T3YbkPJKlHziGNUqBeh2YqW7L1ZPrSIiT5hlJG1EWC8+B95xdKMLSKuwzbCNuwVyr2zMPB
ZGV07Hv6EvwHz0cxGo3RErWh0lzeDLQEpUhOCkD+8HLWOBNjCcP+mGpakf8KqNa7JD1VwcejLN5u
BAJoopyMrSLjbMYVV9dxYRQOIvpQeFU0ch3xs+tmCGh3cidelvO2Pxuh26rvbqtpMi3wuoWGQF8b
upUyQazIhlYeC+jZj9rpWvgyyYsZ8vXyOZULlWHSOm8KecWIsp3sPGiFMtnIIg0zZWQluWOlZEnM
PtZKrXlkwTE22rkCSeIWyMn4n1E/zRzSgC/bDNzaL/K5+BpRUqXuwurf8c0ph4tzEujOgzT3N8oX
BsSShxtuBbuccUO4xBWyd6e8m5k4f+heY2AYHBHt08u7xt1cFdyPRHb8EiC44JeV/6Cfaw9Z++pj
PX0xjuMMl2hzL6SGvqOtp46KKckNpDy+Y0PDQaYL3bbB1w/m0bXncTzaR5vsivrCqLo+G60d8gU3
lPItk5f5DkpriN4xPDjT/bURmg/KCf2sEXA27LhjZ03+nw0LOlKTOJIm8cLS+UWpHmSRoipcHtFh
T5hQ6sMqVLASqqvq+tm4aONKGQASrL1orNlwCfoWCCWBoJWa7jvMJFhVVG7ztU0fkxmRUa20Gd2W
3+Fc+dGrmbvHONHDjOfc6MKjQpigZcupJylb0TS5qugYzPypPggWRh2pAqs5U9e6IgG5lRrBFw09
HiZwiXaf6EBZd7WlXxqWILxfrNyS7HIufLTeZk3/oNQO8TnFZf0uVMkrty8AwLvpvk9p555RpGDp
I1UjKZia89bFzJAjzoRG3U6WM4BzAUZNQQMgp9hTitmbY+pklnR7mwCQNxpiwrRiZkWEXjxb5+/C
osZ7j55wJdPFdMbAdlshE4+nMU90K/Gn/2YyQoIGyYu1AJReGbuZdqpAn/ZCKA4jXEQQ4mKs54Hb
t0bHm20AtHAmK5d5cIKHvoDxySF6MCIMb2bE40NDhGiHlM0tEO5rMwixqqzh4+stjCtWt3mC6cOK
K9Z2QTCb5pWMaoGBjnTudcD6Xajr4UH51WesURekImCT/OyEjjoU16n3h1NTfWf8TyQNyBXaIe3j
uDcoVpx89i4KzvpBfrnPKIiG91nd5Ph1e+YauFLu1JpThZGeTbIxx+GOngjtcsdsa4ZRlRBzM3Up
9DeQOaVTrihhGb8Jtv+O6ZnPm52gC34eQcXrqZjIUcAPWzRk9ikZbssYxVeCBAWsZTky5/5OS1P2
0FVEhbQx738wa8tWTrkn2mMac1/8x+q/WB8c7G6LJ8VijQLpPbOH/nl/iW8D8YD4zMQG8FqvTevh
JaspgL3hTxqB5zhfnzuujx456BUiYNcMV9klPkjYBym9l2Ic3R8GJ65QtS4TXFkgWPqIuRywLyi/
Y3JIGD8Sg8Xuw7sVsDsDRCxi4z1GIXNFI1O49Yr6MYRq8Yi8Eb1OjBu4Lr4uM/DJFcd0oliysjAg
jXBMeLSEkZzSDRipcSsqsnG+OZ1/17UXrwBws4FOM7W/Acp2w97iu3e6arHaNn6FmVUAYnwEohnm
kftd/4+QwDlMjq6UbcWvgSqhX/67z45tGkDzWQk7a0ClQRrXDTL4dYxAaaHKANcsoow2zKxz0KN4
j3wx097tIpKaBfMIUcFP+ZW5vHO4LJzL7HNJEZ5SBirA3DRA2itB4kU5FBF0oUU7aYx/4HDJUqfT
GkWFaEylqWppqEXH71z3LAX7SJHCFQXRg/NuC3DwQ/jfZu94WJZfvsggQIZT9UUhSmeKiukZGSFC
Atu4WgCd2mvZlO8p5uE3M15+LJCXJgElKSLlJKLW7dggbO41eON9gAGVn+wofZ+uh4/71qIRJOwM
kMxMp9Uhx7xcHRv66u094KMUQrgY3l0Sl4QQ6ogZldFCC6syPwwDh6agZsrHVK6RRCcabYN4pqtm
u/OTnoSR8XF+yzJbjw7Kmo8/3WIiLKhn7DwcJ/ZGpiWk4qwcchH32vmyk7GhB+D3pdKAxTnP77kf
BcVbJQ5upV8WidkReBurdSnZql/0YqYqGMOiNDIkjS0Mk/eO6KtA5xNGz/ARFSS2oj9Dilt5gold
fxKhduenVkOPirRufxQug+S/8qWJHlfrQIeRJR1PbKUelIRbZHjdY9ybcbqp74tj2Z5jc54VKjhW
fXdc1voDmfmLFwfdsRM1YQmqby4dN636eliojl4CUMZQLZF0Hm94sD4KryXvsuSiETxNp6SNerk2
nvL8rQ4VDeZBa+Thg3DhBG/ccP2uK2NHwouQfxwUEnTSI18707MxZh/SjRuBPVRxz4qwhQWdym3A
NezaHlNcolEOmdkB/vQ+BF86d3JJVolaEcAXLOIMJiWDlLUqkRpoKi6YkRt1zMrpKNTDP4RP40vg
EaOTJ9Qi2uem/eqjCAHCD+YgT33VvJbWc2348CERsweo1pnd2hl6olUmlj0U9vny4DfZJjTR6tPE
fO3pgyyvMqUWd5Y06f6u1YJ2oL7h2QjUvqvKv3upiK3d0+r1yp7WwIKB1N6R53VXG3+BQjJgOyH+
qPNRD4Whg/O7jKtxaevQ2qOW9NZULd2tU+NrmyUq7yzZK393kUBPia2Uc0g7M8K4I4uxOZUKCiPW
NO2oVMug97crqstUzmtYRjjv0wXikaLlvZb2gSSTjbg4ImOrYD+YRtz4Kc1iv7m7/F5I04JJXJD9
E2hnOmdb/TNc2ho+9h5B786glbPsfX+/xA79BuEdWSDaai8T17UQBvX462mKSDgxfjw+JndCUbop
G82JCHbLDxyAqvim006clN8RNtFX9tW84IAARIn9aP/SFUVmIGuT3ID/sqMoSW4mbGFNh/E4NJHL
m35NEL9bQtgm9fRlRJ8EOvuq4TQHhhQD6tCDuDjeTmkRSiJ40lGwA15f53Urz2YC/jtShWURv6BD
bGu2tKFnupcBZnlTVxp/rZqZBu0hoyOzqJ5XzfABkobvxjBb27fSc3oaeWe5sAO8jO2nn3TG+g+q
8ScBeAjygKQgeoU4kbz89DzKkn4XTUneZ637fzWwnp/6hMMHf+eNjBXpFaMjJK9IxKV8CWue3rgi
uLeCHJ0a9ETDsHTf2UNxkJySMtyeon2Q4E4Wiqbr4gSaoxQK/oQ0Ln/+28rL8VNY5QrOhIuGft16
pmFcYUHwHyMXZjLMsfbRN01bGWZS6sM5E5bvgbFA4K1iy3+dHjm9B2ZYAEzQY/+YZiJBv6K/VHJD
G8qiRkCXwKYm3oOGDaPH31k1ELQztcCe2UNQZKCohk1UCfuW1w13HBUsEQq3LRVLj1wH1FAsIdNB
YgrMt4wynS/BLP/hXoSX/oRlg4tevtu9uL3OH0RXBtOW8AU7c763+DLmhh4vGPSjGtFRdQFe6bna
kh6uduKIttC/lnbx1LAlGvPVIiCaoSJhKe/OLVGwV9IS9QZggN8Dj9KNQZKRJfY+WYjM/RliqDYJ
JwBVVixEGJhzXg2BLBr3FUl9X2cvgpYJBr30PWLqq9SYEMQ1trb+Eekg3ABFTiU+MLbohxRh6hSa
RpsYtLP553dyT4jfZNOaOUUBasfTWgmkxU6Q6lLRiQRlMM7ineu7StqfcPaiJu0rFNuvhXJ9X+GB
bewSTi1efLbihqC/eO/nroOoxWTnJmswB0ASbu9SX/NbapUaDmlhLqAP20YEKFLL7sm8k/+R/hqX
V4kLiAkWaKl0OYmAc/7dzWNu1AqT2jMglzp2J4j/i653BP26XK+Oya+E810jMywre3LCDK8qGkHF
WnDNmeDFvsdjopB3JRHKcclAZ6opWB6NZA+8VliVcbk3s+KZgxr6tyg9ggCdb256vFfGeWF5T/dz
l4gUuJcjApoIUqiNK/UZZmzDz/tgk4JEGe1+qFQIvnJjrUiJSd2Y1KxnzxB0cPPE5183bA1DgU/Z
h7uNdovhUlxESdkYGaBrGNotXrjy8XnK5xylH5hun6smmFbaBBVLeg1lz5v/XtntvcCFh26v1+5j
M+s1FpQyCl2t2UrRRbYHwe/AgNS1n2KMUBOMRWEcHIRVRCQe5OLmUf0IOgmH+Fho8g3UTPVSTo7l
LsuwHcw0ZEMPMwsy6GsJCJXHMCEJ59DQEjRoNuxkCOVAfCTbh2f0azYAIfcCqby3K7XhHUIWRP0l
bICHUtgvHE22vAn6h7Nqoow+DlxFDFIy7qp/4dl8Y+KW/FvcRAJOG7ULraLzeoW4LZCD2p9cxqtK
IfM1EuNP8yobFZAm+nTl1GmXKkLPMpdlhmnxm4bhNjcjZDLfJZYFabczWzQgcaUv9MN2a7RwKw/t
neuduMHQaZrSbkQ5444d9fUq04qqdjFSHjtHasizJHfnyWdiA2eeIj4eWBKYwfSksGE8dDNwvU3a
Cuu+OAru0TtPbriMAPPJOtUGdJFrhFI1KE50HIz3YQluOmh/UAN8d0Sho7FaCQRnqzqens8xVjje
nYP5jp6nE6ANs6uO2rnckOVI3VDCCDE0NTNSIq66tsImK67J87Wy+k83bhWTY1h82Rhwlmo/6TYf
8NRn13SB8ik1JIE3188OxfCWNvXIeH6cYZ+fJi5fiSNRLXDGIXexHdnWIBj52xMmIP4tXEHs3XfN
DmTjRecrwUYQnw3SINMMpjiS6mcziRsy8hSu4iQINdkhrO+54CB5BcTQ9hjtBgkm8+Rdd0GKrc/I
M5UUguRRDJBLGr55OLzT9Xho0mLj5GG4PnMPdtweysPWKqj7wEbQzCTM5cLyPSwOL9GZTU7VJMU9
7Mj0VLZTBn/ACwWJOBbuYGoTsuz6wfKGnYp3RdKA1kGD1s93r51BcO4LZBXPd9SG0Wrf3rfrzHgU
T/aIddsc5iExAUUrK8Ky7OUa9FVOlSMU5TnUznDquQnqCdvYkBrG4hMt45p0/chZ3xfnLYeIYiLQ
OMaKl0gtVbnh2Vp8a53rpGyrzk3pAzBszaCR/8GfE4gIj3tuP5fJRMEnjGM8u4yWJlfGtep/yO7Q
NAtFF4zSaH8B9N4j/MiGba+dnXMN2BBWlNFKs8rVFnSns6AI40Wcm7LsN8aWIoA1+KiSFoRO4i29
YfD/wDCjkmaBJPJAFcl747H1xx7bQPrhlxWPhuB61Zyp09uQlj63/mLXcHeOFE7I5aDnN15acIhQ
VOgQX6V248LSTtxesGs9F1PWsMSmaDOvn04NGUGz/Igbft/IyCBnhONdwi26uuCdMi1x3c7UEv10
QR7YZNsLR/lOGuk7TJZmtYFKUG7n3EHdipsoaLfdmG12GjZqwd+ZCgYK7K+INwcwQErWL76yJhyz
hP9yBY6kjWZtY2nJCNsSp0/MF5vgFBbtpet/JEtalMSz+XOAe8C3IRWs+ryFaoaiKvu17YfygTr0
U2XO1ZRpgK//NmlJfHx+5zdmFZRWnTUaMbyuXP6PgjAMHBfgTWwi1QXXV5NXBE1JJly+3CStCjR4
0cFn6CkcxOP3MvunMvY4wNtB3JcMQHxDq8AS03ZeMb47l9u2leX5iSHBBCzuaTF54DuSmsVnR4Ww
JDxxHJ6vcFPAllaz0cx9LmI/eTPilDPMw0IzJo/a9Q/bBSmssgUmNRBTKMFvRnMZ419sjYL7C2I/
Z1KP6RmF0orobvjfdGpdgs/7jzAUMI9AaWGOkDXqO9Vz32n5YoADQ703JStqpWTDiZQ7s0suiW8b
iQkCDaX9gWXVQewj6fzjulkV75ED05XBeHFqTgNuShrgL//2Xyk4U+D4OjCls9lP+0DU8IBnVIdq
Ss7OVWSInYuXkIXiFgIBTH6YgdkzH5vtyGtT+78dDjZhz/dfXa4Atc3NNWN1J9qSNK01qvOr0B2V
vB+3B6cfQH1U3KOUYwBzbvNg6K4MdmBulUklfLr2RKTF8xDFVRd4SGCUyVx2FFgLaBdO04yuuiNp
2OOuJ19R83DU0nqqDv5LwGR/k9LEY1/SXaA2NZi1PysbV+9MOewXbwGxPAcVassdJiLIQIwHCdtn
bpWpTC9WsLzKE6nxa7dOyAc88eMmiFgQLJK1DQ0RkxkUKQSGCRcGWRJ8OngLWPfI3wJh4C7W1OAz
SUyoMEeA7NI7TwtDCqQDgYWGKeUQimWWRthi5c4UXrEdgCzbqZsmVrPsDwQt7eFovQkJ+/UaAedg
gYw5t4961zWH6ENYc//7+AwrpFxNr5gfl/GpA/oUty50RPb57VSs7NXV4mHLeQe5WF5F0QjYBZSy
R/OAcnSJORhXKgx8N7HmhXQaoQUCxGwgoR0OhuYvoJrwG0fnY7Z9RkRNoK4fgNiiIuqUoc0Dj0pk
SjU/Q4f8ctwu/iwwCFc2RfVasut2ECkZnyvMM6nhh1reagVYq+Xd9tkKcGm+ZNUgnyEi3bJ8RJI4
x2i/4A1U+yqR+wG1613MlVPXeDbWox3szKwcWA9hAdfIHp1s6ws8G+n/NEcczIeMWoiRZ5p6ZFe1
5XEC5X+G6IkhQp+UbzwMKkge+hTNi3PGP2zir4bOWGz26n2pYjXQiVnpVMLYUXMHnVzntL4gSPtl
gK1PidC2D3aOxtAWvmaNbPLVNa8P44JQodI7tf0VXk8Q38ygQ7wFhtlTiInPFFbvnvRmzdmX0F07
D3ysgwcv40PhA1PjCmIIWJV6p+PZX2EgGUpBxgXCH8TWxoSKH7GnqFTdq0MPQsMyLa8KoeKq5LqF
kQJ4ymKQyC6gfowSyXgeITauZaQov6zfihr5PR9nOlJAi1SPoJctGGbX+st2Yq/6x3UMtWLHo5We
v+t7xlB11+0vptDi0toNPc6P9NPtv4KUBneujvqh+9BZwCMAP79CNKQV1scHSkpDej3BVjsGbL+K
lSeVOl3zi8heP0ANRw3NICo4aNL5Kty8EevG1YSwGHxvHttw0mO4Gyou8iXFSnW5mrYZddczEjL8
5NMGXtytzQxHkOaP6l9sgvg5NOidAibRbpeHABnJmsE/2y9TyAhQMwFhgi1T2130jc27XxyCkVjm
NYVEEKmiWumVCm2vsS3jzIOCBZSUODBircf2P66cgT5UX5jOZRYJ+WzlJ6uZkw5bruQt9mk8qrzR
APiMI+jAsmsUKI3uyp8ndBYeLpRKU6KbP/tNlYgm+Yn0CRfZQyqIWf4qLRl8prJrnBxL/zEzorTR
wnWUUKmT/m8dJgMSrfJhKTBDodC8KoqSNimec/hcUiYRqdPzi2L4Zh0zc8vjCxfVZDJC5RaDj4/x
Kzc9y98PUeqRz2tcRlg/3gmQYvif48SMQVxigkNN/DAzJLa/1Z47jbDJ+YOSmaQFqV3ebVrbHZqv
l9ugCL49jlFbSPJQtONOY0JAT0Z85SGnRHFTGbeQt5v4mkpwyOpruAB2sGg4T5GyO8U5mniTqK81
y5ccwElYEqGllxbSBaA53n4LprCNAoym0tstPD2lIhTJSnAt66aPW5pmZuQ15yw+Svf3fU9vpon2
P56jSjBzFS+pQewRJvQFrpR7e2d/lAnhecaDz+FvV82T3GrJfjMhc3AXZHFBzVkbXvgWWOuAVzjj
dlvMJijQUxChR2o/jXoKTZcyafvhL497P73gh7t7rUjqY9kyoN0TFaJHydJKnBXuOnayKZgcD9AR
n6OhBnUM+FeB8eVrse/JCSZdiksWBQy1DdGSSIsMI+jSlouGg9FgC/tsEsAIa1NkXZIhnx7/A9of
2nrLovcItlJKAVI9THT7WhivUABpg9W5VUrf6Ld+Y89zRcltQmIuwi2J7yawXKfYYBfoZHjfEdmE
iP9x0ijKyRkMTURZ99PclLGJnXCZT5HORYYtaeCdtlM565QViWGwQaTJgB7oXLeVe56x6abxr319
tpF+uXMXSoDySdZxByotvANw4CioEjRzc8ENWcDsCQQWIAp1mHhn2skbY+GiwwG60s8Olb4uruFp
qEmVglO8XCBEMS0DPUH57QNFc6YC7T7FdkriXNE0M5vKJFMzcaP/boKGcVfg9+XJtHn4MaGQE2ir
ok2s3qfe7XHxuZ+/wxly9yrOy5EA42iCYogLzcS2N5xmYskH9I5RRbMpIj65m7lQy8gCR6Zq/d/9
0ur3N0z6pH7dEaQOw9z4N5f86sAkdvAb/vSH7WvyhxhgYQa/duV8RrJxNrBNs9wXEr+PGUEHpMH+
vUnf9DCYpxC+ajwXRQiKbQ7La5cGR10NMjbqzI4L0TSBiN4RKwI7Ez2tlhuIzlI98bBTLX3xQ+EH
c91yXDVAxE9fCkAY26xQq/geoWrBhR3LeYXSlLOIYR4lZQqwB9e5+tphCMuRbkQ2Jmr1JXc2J1ib
CcoBwSx2/8zsBj7dHW6qT0u8Pib9sfnK+v5IojvdU4ZWfMue5sf3U23N3NoL+hbQJWOAsZ1bTsja
Rcn57kEVxtMR1SzmBmwaTm0Ymu5BwilbOlCkdkKluQpLVxmW3OiAsIg8WhPYy1EAynXkBeUzXanA
bR9ppKaIe4avfJ5B3YpPIqYCbMrD6Jk7rG4QUAzHm4xFrFNJ0nQat6m0taNMFLb3UhekrISMCH7P
/7rImihAy7Nfha0ctfw5M1c7+eN5u0vUHiPA4kNzDpbT22O6k1YJsYTeeVYG3Sx3uGszu8aNk8lP
AxVKnmt3Bzkj++Z3Kpy5YMB7QXeQBCZjaq/zXeh/r0H0VES1YRooILIi8OuPowzk6jGlqWlUmz0n
Cb3J7rslSj5xboWkY08nzWm16brQ56hZtdvxpsLl3rRyHxBuVDOWKRiYKh8k+DM+Rvi2En1O/V4x
o6ycpicHFwZgThqggPB+1ekmwzRg/+zKpvfdHo5orsAPICp9zKDddlEx9JR225ZEoN9aae3S3JCV
kJGF9mtsmIk4+NySqhogn//0u5welKQxV6pSapiCE/8YveVMSrYuko15q5GkDuqnJIMAoDTmfoKu
km8QdZzxwcGYMhObxkNN1INRRjYYqYff3mAdyHVd21WdxxIx5Hs6N8V1kmVrwiBOypKDSndzYoeK
kiMussniJXcVdzHL3dkgiY+3UHnyU7tHJgQI0rAUBLt2I0VGNyV+/7w1l6vodwhKeBmnjKOxMGR0
hu6lSIAqhSE9s8HxiNKH6zw9EmWhW2cbosxCkuG8rNTNO2FHmtpozXyYut5sNVAlsSdwRkGgyTe/
H5orsLvdjxPL3+wGPtDpxcNukP2aV3rVtWtw75weqfNbE5292xYbXSLDce66PV7Y4uocnnj9WaRE
19C0KiuOxnMpDF5HRjJ7CWldC7Su30PNf274Nm7801Wslr6OW1bRdTcZB88AyiLQ2gMtYjyszO6q
GiHfB3+k4YuMtRMiLtY8JF4oufUncBZdU8F78YEBDMOgG0VqfieTkDSbjv/2mas00JIKEbN+l6A9
KvKivabuKa8Gn1unIrZh2cT37SDLCc1W/sJFB/WcG2SUV/St3d/QmKN6nRFOM160meFx0a9vaxMi
Gw3dNoAJW52LHylwmdUNivtaNhM3dECSVyKk6+T9mhuMyVQhpa3izeKL3gpoFc3r5eMwAcsrMoza
4ksMxbqO7N4fzlylSs2xDhiCEcwyv5KDSsdLRfSXuKOC1Pc2ioYhc/LfljO4VX9+C0sRHRIsX2ku
rYPY6shEKvuxHy4WqaEDW0TFXurKX2kKmWiWX7GQ7PuDnHfQT/TNpKBz6qcJS7EY3Z6Id3T9KbEt
w3T7IrRjZuRo6zul7hhRuKGi5WY9exe3UJRrPc/oGpqCiAdLD3OlWxp23q43DJaWN4rRxyNhdfMo
aqHPfkXGK6C3rU101qPhXXt84rKddfgHjkQ6QH2z9u2XV8X2ayY57D/v69zLN476HRUDicvFlIIh
/rbFZRHOhV+eaE7R/saB+IqUkSA4hcRXCu23u/0gpoGzKbPF35Zw5cpHmiNExMAOQpk31DqQ8RpZ
2xrDTw82LaRaI3U+cU75f9Vy+peobbrAtXIw5dHrEUd+/okdcdYQuKlH8eYtS3XTCnapBQVF/pRR
2IphL0TBQJOFBdBusBWUTOYTTmq1zRctPJPwAZ0t9nw84Tr5mxJPXqS/NwQ3wMnOI41Qxh17QhBn
7zE26Bu+WBcWVkYlYohT3nzcaVWBZUj7BfUnmtXcWam1lEm6aePqE0h4fr/nimyEQ1i6i9iAKcKP
jUBVLetWmVxWPwNBhT8EcPVhMPhECyet98DRbdoqrVOtR5Ltsk2ckMVONmsvbhTxO5aSkcVgyN8v
Kl8BCi0XoYtaeBgArxWep1+hUMYjF5ksr/SCboVlW4wJVZGQaYUkokVU+Usyk3muxDqfuhwMBIdq
erR27+b5O87O5j8PXpxSzsCLDYi4jw1PX5ZaP24vhRFsimSaZOw3rWryMe/A+7wTuApjZB/8N6sW
+dLvhw3JA2GWGC/s3xBP5fyuB7BOAwbdYZ5fIJPN4lL5iOqfpTYT1knMHC7R7pxD+nploYn8c/s0
AEkSOl2Ff+MHHJL9Kbglinnx8BhV0QJ+GdetukogyH+D67ybNcDmzqk/8MsYzH2bHKfq8dEp43JE
ZpH8XujgrIur2mllTjIsq7pdwvnOIxP5rUNNfCTnitYkCFKiZ0rQAYPLGEqOrcyCZoePS+S2k6CC
SxWWPpEaTLIRY4OZk0PHGoLIYPF6+3TcnUCx41FubA8l+f1LwktNwK9rq4H/1s8rPppGVMQfY1yb
BRk7ru33f1KbDmD4EI+Uoy44OWhlmr+yZcdq7UtgUySAYRJ3+Hdo4EEAjFUpLkRJ3rlC2ufEwKzR
dK3iAdIfSWeg6cDnOOYnC/nTTRfXHMzCC1qz0oJ0z6xgZfN3IiMJi1cnlRjZjYjbqCRoJhsfTGWn
dCjJwdcqOnqiFCo19xDAo4p7yr4ekxj28KfnI2v8tFyFboeeURs7Xz3Dpcj5po3Vvc6XIAcgk5i0
56E5nqe9uZ29KlFsKlpkvdwCEsvNSKcxPyvC7bR3fRLE9wFOuAfWaFgNjyi5QlF95OPmPz/M+vqH
3w0j5MDeT2ToX05dDi8MXFHaG6fkNQUzTezF4+8l49qMeolBVENDCacA/+yXCiAT9yGyUp6tvkMH
PQmNSCPRFTwoQy1IcmAHHaeduYvLIw2kwwbjp64643L1F59uwiufALKHaKMdvLCXN5pzD7KSbcwL
leGZLiPPfuXgYO6bGCgc2+kuMbVpGlyvBNMtWiXxYPfvHeTBnJJ9uyPvgSorjrK6v7/Gns6enVpO
9WFxgNfMwGmD7AcZPoxV1ncuV0FybmccGHbViihgjvZJwn38wI8UdU1pfctukJEsKOSf9m346qAT
h/IENFTSyKyYqR/CdDwDsvom3+vA4cT1WM3+btpMywwbIAiwFBkBdXDBZ2bwyfTgNecwUnNiqPF2
ODaR4vwvm5+IGeK8e0A4CzvxTOGyS3geAye1sa/LE2cC7AoNVMWOHe6yeGHSEDoqElEuDvcuEXc2
FuXnGV3Rna/pigltKiK6Wmkh/nbW59Uw4XMYhg/c9wB5euw/74sg57Fnf3NofCathVvbMOm1s5k3
88A6BS+apm3LcjMpF9IKRnxMGNT/OAjBuD4oSuLchK/lHcdVeXMvN0/IbNx5z7qViPgRRfA10WnU
Ui/7+rOxIoc+CKCGejO5Le2LXqFWVwxCLKcWLzLqvWb/KmCNLOVsWxh/XpwHn4cxARPVEn8QJo7V
b1wwKyrh819bYfzLhX71SaPZmCBL34ArMyjU+nqFhgqkzBjO4xox7pRZsFxwmXGVwlPbXiHOSlsQ
1e7xdevitDY7eAttF12XyWgYy12uUcHLkHqibWgFfTZ7FsU1t8GdGJ8BntrtGD/ZWbLUlUkAZVBq
TSR50KqrLD/NYfF0BqDnb8SWXIqefeARvBeqzfmLGou6oULiiqAWofgxJG6xLyYIDt07nL9BhbX6
Vd+0c64XwihwwW1RjTH0mxJHcPYqGu7GL42iIEe7r1/MXmBYZsUu63xctmCXm+hsWxBV1nXNXh0P
7JEVGOO8SgJloE/o1tjJz8jZjevii9fK3XDglGl80k4DucXHrrXawH8sW8AIdFmGpfIy0W0eNq2K
ZpbI0ijmwYd8jqUowgweEuUBuF2p9RbS9J083AO1auZIRYMyqqqs/FpfwhLt8BGuOz8KCABMNyfD
oI9W57CW7Nul5H9K/ZWmlU/6Ug7LC1Jm1L/gDC4CAa6AF6a3OU5KVOmvZ90CCy0BtF5bNgegbA+z
afrttVHNSGqn3XVBBop+GWaNBM+I8Hny+7pulw0WOz5sCJLWNSA3JpunD0xRm7xTjr8vgU7Nm5Oy
Mtw5y1aEyaaQWKNyRXd2mXDLdRrM90aCta8StRqPC1Hnndho7vvwerurwN7oyOED4OJJ5OBmfjCB
v2jyBatVCJYah6iuRV5dSNRmx68UF7zdOxrpogp8l9nZPX8fwrkQQovW+PKdE39UK93QJO7zSXpD
trjdP72pS8qLVu6kQLhLZppwQh1H/cn0LTjkimbJllotCETPLKnAv+tFidaF2OwhowR4zM+VbKXN
vSph88yiKPV5mBtPwpphwv79CsyPY4167w6OsZO3rGSm8Ox99G6zqjJECOu+VhFYkUmBBnbjFRxN
A8bb1nSWine5eFbSV54G+Gj0oXSeZrmdWMyu/nlFLYQrrNHEvvjEnJNCZQGi2/KNYBmen03RbS7X
48ky/wth6ck71qNQSqydLIXZ03kjKX7Uv0f80Pr5ca7I8V4vGDNeE1UCBX/KfpVvesnnBIh/bXCy
xYQZwye87vVVaUtKEF9qC9ozxK54w0njQ2+qcj8H39oZXpKlHksLsQQcEhU7ZMDAwTjJdmNv6FYC
GxTdS25RZCufXDUZOR8JsJeT1nlEDJDp9w/NDcjlf9BE+P2f8e9dD0sNDmJ/amHnP/dIOGMFhMvS
0Upjy4Kp6D/dNqkHzvH4/2UX9YmI5tHWLOpO37H1Qi1khkDMfOCZGM/psH78geNGQXkZhhizC282
i6WXGRhfCGDtJKdf4ruGhA0W+36bIEts7Sc9rzUaxhy5o+kaYwc/7KLrBBWznYPwGRB4Xkr1Upd3
quZjDByhrNczmJAycO9ofc0O3rleuZvrtzvHyMv3DMnovyMN8uXOGC3pcOJBlnorVi68aIdN61rl
dZLyno+l1Ujxm38mAy2U5lPB/0XYYW2/8MYi/ebQB0n74l22Au/Hp7ipZHeJx2VKpoVukWJDb+7R
YpH8Ovmesec3k5+7eZmzgclmwvG/qXTLlvd9/RAiJVkDLSniElATKBivX871uOMPGwL/Xzjt7B0+
gtUF4XN6iIZsipHR2erLLxUjTbtdikmPsB9NwOUhpVY4MHGCqvZ9vlxu9N/q/Ifo6fbHcFog1WCd
ePYPyPXELVredB1gaQQtVNL9MKg2NZcbTdU3X0aX8f3AbJZOrrKh/UY+a7uUtAHRIEVPE/K4K+Ig
Lo+fv7+FR/ePymS/7Iee51APkmN7/041WpqJPAwKUqUGvz9sSre1maYJ6KaP0e/+KLyEvj8kRhbH
1vgWqXIwWX+svrvfiLYfLvoqaDONJ1dkc51ciW0tp6uS8UzVw5UtiQOFhzwgZhzbZn7BuvmZjryI
ZP32d9bLvp6WPL8cbLi2SNsKr6T0z+bApXZ9l/pKfwkGjnaBt3XIjE2KICy07Hk5+IkByKBADETs
H/e3CcScxtc0qQjILCinalyMAX5gbHxZ5NjcRPX5JccoRE1dn2/yoG6L7f2STEVYOS37XxAC9hIi
ug3oZamVADyCxi6WNq1b1Qn6+7ySVEd68BnlvANzeXYgxnlLK4QqtJRLEJYKiaziM8AZwcks31KD
R2d2a81hpMO0C10jlvslll/CjHERnDf/PIrGB16N0Nd0rCD2OEGKAjNqzbRjhUxkrgvZuSg0sdtX
t0nm5l3s900oEuBNF+wRs5pV49w4wmozbIuaY4dn1r0X8lzFFmsWpQntmRTvb1dqi3blTFKT/A+7
O/1P1k6u8EMtfQDN5dxN1CiAbFZROblwpdEoEQ7eit5f/ohHEH4Tr3RPoEswRbimhrjhqi7LZZX2
S8IBqVAv9T7XDc/UxAm5Nn3aeli9wCCzlbqDyVVClFZ+l+GKaWrrfbABfu7i9fkNQYz3pLSowNt/
Rm5vByUin6Mvhc8Kn+4bMWYQELPyOngiV+EXkhDS3y29s25VJcZbv+CBV1tKed5oKggb5NTGEuid
Co6mVToN62FiRKeQ0kBYFddWOXpz1y9IeMzxdpJVkUGEsGIUwgC090kDXYdzTB8eVjJCbC5K5Y8L
Q5kNJSQTfifwIo55o0RaSBOXPSRacjqjxyxRZ6p4UGW0kTnXCh2m6Ml+CW1DMFBFe0bf+wgKbT/5
K7tjyxkrb5iMOWj5hT52D6SsW75bXBM5+MyfjcCAEB6PwJBe2R4DVzpPlgzV/Gemnqd2657fAsmh
vs8rrrU+Ig/hHW82q7vkE7pHJoybIPhk6jZ4jGe/wAYjyqF7Z7qftNJBg1TGgYVaQlGPtnoDTbO7
aI84GSNAtVlrXwikVPeyWMUj270ykHTDfB1yVF5UHSMCxW4llaAY7dPsi6mAOSYnapxztR8tjzxk
zgBkeGTqglHx8wAdgh3DM5EK010LzXkU0iPa9uE7cUe7DPsZRtVIgQlaXX9ZRfwA4wPSq7sydVFQ
IJCB1xLGebDldCsZObLeQmgB1XXUoguQRJ1LGYZSrxECwf1H0uLXyIJlCEUDd51M5QJLys6fM0mB
sqciN2apB+peugOuxaCW9gfB1RwtsrnVROT7T6u462FvCytx8Tmo/aAITdteof+110ihzftzsIAy
LnDn13SQQKO3oZGosv3+8G8hMhFF+TdNpQfYnAGOsgUW/WUpP4RdAj4enTtvXBP/WPRgta1ZxNgQ
COJxVZ5C0up0cq4FVYmjougc0sllPhJvvQtgtmk89BtxzF/qodagAOeUT5LL3bEmrP2KZjYPdeSl
jZSyXy04sr/nLBcvy57ER3kXDGjieSQtD8eEsLLiYcCx8rhE7gtSKTOIhALK0lHfx60vNyi4QJ3t
GB+ISF7UuOTKprrD30+LgeJTcL3dW0/X1i9ms7CJNJ7TJd0di+rpOoPqVRX/pdfzNV5HlhJD4NX+
JPAlkrUry9ZV5fz8PWApq1D/PAvuRg14y2jOC3vjs4ZjAz8csbNlMCB19v1xRLom3Afkpl3AImjf
J8fixNqGVOK/TPLs8QilF9/xSO6tnm4LB1ovjvN+FIBYT44rOq9gig7Yen0sYZRZG0npXtENGCtW
FVI5Lqhbp76zgAyAbBDHSgHvqczH1E84TpZflSgOwXQdDetKsyOLoq1CEtJmWveY/2bRr8c2wNUg
NcaedCxsnhN9nrEQ0BACa1XaM/YY0YNg+uNqctuKHfirb8Ub5fw9gJf/2lVHVlSeDL7TzspoTiqB
squ8RdjbWTeOE4ZRIQTCQcJmEd9sr9vig/+lm8Oyt6h+BKu2hqir/pie/sqDahsqlNAi+iVFuEKA
1yadbx53hjAeMGpmS5FYUreF68FiktgfyUh2YBTeISnJ1qOewvg+E95QkYwSAHAh3xqmEJdsO5pO
RegrtkdcV9ObJLT09/UZpMvmMtiGWbPKttonUSlIficGAR/enkCs2y4hsWoF2BBfxOp1t50u4B3K
8AzADr1Qv5WSjaEAPkpQODN5tAcn+0CQutSUCHiACGY6vij2gE7PRAlqNC0zlV+PKv7h85onWWQz
CXbxZnStz2J2cQ49y4VXS/sTngx+gTT+NrdRGfikahNAkEP8FS1bd05rLbio2ug1ApNStiXBFjko
nNOuIs3fE8mmoK/+MzzymYJNjCmZhVci3l9cZ35IwCdJr2zt1M7LRIVb0pCBnT2FptI84x57YsmY
LkYSXDItRlQrkMwIvAYj6wdsPLaGBHZrWW9qCsova/IyVCkvkKWtr/oLE04pq/xF8cOC5dUScNOm
G8KuOnKUJekpd9pf5q1U+nN8HTjSM2NLAKSzI7JHdz/OMdXcTw+DGnjDMnA6FxVOkon6RGL1K/Jj
h2OOzxEAZySGVEZPE5dgkmDTAgQIuJKBqUaBkNPmTt1YSkt+vicMKQMAnRtp0TcrDYbn/5+rsskT
rZA9nsi4ETcHz41oc0IqUPJdHqTAG6tChfxvHg1yitwjBCkXJf5QKGR66XApeWiVqLK5+PHYksUV
4egfnID6isCANYP4LHr/PBUUJe/gf313+sX7J2LIk1GAZfzf5maxn0oOPPVxT4v+1mFUIu1MOH65
PMXjUrSCJuCCGHpYpzmxwEpBAoS3A3yAFiVtF4LYlSaxOu/HU6CgyptTbaEI+LNPtAE4KSyvS9Qe
Wv11sD0JmxLA511A2lsdQGeLpIqZG7mbxpmfxn32OaFHaYv0v64cedn2J/zz/y6M7nRaUyE5Gosp
5BmcZJSeJASei74eY4ZEYijv2O9tCBGzwnZ3gWFzECeRaWh6gnywlb8zc024K2g2DWeqtoI6kd4X
3qMO7qVQB4H8RMvaYAC4EUI3K2wJrABALe/CoBF7ZRegtgrS7veWkqqLQqxqTq0A3w25TkLjMDaH
d6/By/zScsE6/yRnHf0azOhxe1W4zYP9svSsee7T/uO16Vt6ljqer0lDIYlLH7CgbVAFwvV0sYuG
W+r71FM0JLilsw1kWKfXwPbYpG3kSTk2qVPBnHiO5i1b5gqcDt3FnMVCxYwbgKZQFpPQn8c39hRe
BGzc7o6oHyMx/u/Th5jaOw0LPlnYdBgxB0C7N6pUQfRd4a8wwnRmm9eaSzX9Y0ybrGqgVvMTe7FL
GEvdgk7EGIF4tiu+k47tZjzwbjYgA5epRzSXtfJDh0nJIEOFMr+/xnH4gfWNUcXul+FCnyfpkVVQ
kDDO7ze9c7Hn+f+fikrP0MVFWf7bDUq9eNRiljuB2hED/wjfuH8UvzVWdIq4He712br30o8nfOBi
okSM6FBBc5C2qgAculhzndfhZ2DQpm2H2WVP75RdDzmSwUF00eftFpIkSnKwVc+Q8S07ViB/zCly
uOeNVM1OJ07+rs558/2khy8RuDLErDOhv+UPX74kyPGN8rrPClW9efgN9uF++RbYs+/a1MWE7rbQ
MRmDwFucIcL/8Ci1+lhoA1Mlj4Sg0SS1qJ4Mb6x7OOUWRrGL7VwE11FwnHA+izlK4R3tuVz2aFdg
l5HixApkQVB+cCp0PUejXNl8NRKOqNZrTib2EiMn7FEieFj5RyPHrodcZVFW1YucwySecju0lL+k
ftYXny7WVSpsueqMeoxy909l2rhW9YAqOeI5Knvl2ShLrWFxNr0nYsnUUqZZZhwQYXYvxWcCcwxj
/hN9GSFjHIf1qp3EwAAc2iREFkI1G3qqzrNJjjGry03tagIsTgsX2LwpPnaLdBg/dfVQJSwmfLVa
8W77lcNBBZzYJ2W3EEjMonjY16xxOy0P2FJja+Ite4ZUgu1YdL3BTWDRQGNhuf1V3cy4S52qYTUV
un8TEE5mqn94TKoty6m3eszMbdMLghOySwj83OjqH1Xt4JKALsOTzjzlgEmVWmYc0TWZX1kS3QTz
RHASG/AzEqWiltmV1UweOzEMOJAkcIcY0ccVlyllFpWW2pr6grBuyEy0JwfKDkkrV0/Oyx7QtDb3
gWaJYwoiZ5vxxmSse+AAyWoQNahdV9OTXSuLsOAWik9ciGS9lJkAGW89rbuC/qfS8m8YEpGDnu7v
N54rg5fqJTuXjxbfNkjihYQ03e5xEPDrrvhe3LhBLOA/+kuNgCmzWE8F9Y6Q9FBE5kTOh2s4yZAH
A6s/1ZESt1oJyGn5d54u14s65munzUfYii6hEP7zfsx4s4EV+PJDatqxAFmP/ZNP6shJ1DnINcB5
eNwmXuPvPgG4Eg8aNBjPfGsCodOzScEPWtWlSkbQj6+J+8W0fvO1WAaQTdBaCyj4nPNzG8607UxA
vC4FiTEJo+S9HO7bhcGsAvAn+vtcsxBKLmWFh3OdD+ddiRZEjtbZzEIp+HcyMOIJax1uKmQ9s8Z0
GL/Ajy6fZb1wMTU+i84dJIlOBzD15EfVtwmu8IlaQFJ3MZfMDntA/1sh0YZAC1/StUjwsuiYwztG
3v7AawQgEXyHHuSa2QmmQZ2BlDvQCzb4hj9G3WW1WDc2Zb6wnvVFFPAY8ygzmTrH+0LoITwWh28m
Agby0gooDz4U2FWMn3xjC66OOgoIWXsInQE2xrI5kg+uG3dEB+snfRJbgq2seHzom0Q4utSMHf7U
JDQegY3lnRl1NG01CsTRoyZRhk3G+mH/YkkmMhXclMLYEn959ZGp+L66EgZ8JyqOXJPucTvfDaVZ
RnTmKPEybovwGBeDLN1xSFJga0BSu/m8izZrwrBnn2mvvz2Ek7bbflxE9+a7eD6+aaCmGXGbwJOT
SgUz4hLQomPMU0o366J7Sx7+mSOAmqcFhqd0D4rjUnSlULiNlXn3vkMmAnd3O7eSc6OSBQ2Rhp/i
Zc7PRoy2L7lzk6gmvOfbV6Fvg/DC2cne6tHLVI+itWZTCZgFHv0K8Bn5if+mph+G+Mb5GizttCmK
6a4CW3RlxNL+B/TL3dx9hQDluq6rtMLI4Snqgh6zjumE3I+0LdqcsyJH1eGffgzwVE3+EKPr14jX
OK52tj8tepavgVB42au9PTCL7Bl0sR8mYu0OXwkpLMnvZbTfbYfjKtbJO2B1yG9fcvYKTIIQZ73Q
HEguMHWWgga0ctqsU9nRvU0xzhppFeeiDOXPJFSRW2ZmUcXtE7EscFFrACo40cpitN4m3LWG2kqo
t8rYPs0KP09lP372NNeXppCR/dpnW4hc7JoG/F9nJhMpP7yIfX/uyMsQKFhvnwVDH3yDsFZe44ju
eUFi24rLvLcStyMxwrcrs7X5cB8KmAjowpXLrh36Dge5WWxvXFb+p8PWcs+GGxqoe3+dXaX8J+aR
tBZCm74Yx4HyU+x4VZaOoFhZpjhb34OUNs61jgBZintVuDTJ71jOE5B34zU7RghRgJ5C1Fmmc/de
uvo9KU55nDIkJKHfpXyx80YdSL3W43v/uWfWeT1JzYi3XkxmNEzespQVYlKy+xj1AoiaAcbC3Di7
EYNIfW13fYvandUhq30Etv0c7Zt3los36Hoda8oHd3C+WR9ovhfwuAWc4xnYNc93NuOPKh9n1Y0i
FMxuyMywri0WBG0ZwYf2Uy/L26OTbupMNx1TtnOzv51zx6dZa6AAcN/yFZCkG8PW6q2slBVzcBwT
gAB/TbYJshyhMK6hhh5n/HCCpx0cvBm9/fihby5cIEjEO92Xk0Fhre078bc7Dt4yTG/NLQDL1PM2
mIKj6jHhiPkYVJVx2YG4tTcRJfbClgACvFCmjBonerCN8CYMBwhhyp0o7H/Y+OtsQVWxkPoGOBRf
DPlNKTrANUUGacGNKU9+vtFw4xZd+AkAuW2Cv5ZwieaOlBnao8L30y6SMQ9eP76F4HWwc7r/dHoq
nQHdf1E3su2rOqFbVhDY6JqtOfXjfgmamdBL9ECB4smJtqpOs+Oo7TMl4TOzwt4y7ts72cnZoxTI
trADHUuxxJvShgnSXHMwojj4B5QKkDm0t8cgqEaXtf8ZNzlX5mSXAg4B82bfnqEw5Vl5Glx3iUJ7
XS+dd8JjCvt8USyUVFT90XtmhVI0kG0uX0Jm3OWeaHB2LGrcJ//rsD3ylD5oKZrBTcz2dI3wKxxY
F3Sst6RDWzIH4CdpOvBqTGPBmmF8tktM7Ce/qb7/Ge8oQOyAed4CNO0SNsijRp92zcRRj/c6Qgcu
yvpavMnYn6oYY/qO96kJjfb1OUW+LaGUBuqD2zzoKS9G/Q1KcRFNeQIV0xBvHIcmyvJr0ME0YBBQ
55IdsBLrddfCqCDLQc4kjfo/wQVRk6ePGgnbSG1FzOdb/aNHu9asAy1VOHri25kvtOksog467AXm
vNUNhNfyOoFWEnDBKYDtgWxR1+5NJXbbCgMNO61bG1idZ3zyl+v93amhPMT8B5ZowQ/rHABdtYRy
vnvelFi/SCPwX0h9qNBxZ8th5z/4il1FTE5eCiHPSSSlJYVZK0hHqC3MEn48jcjgum940ng/7scW
7kzoFjsKiea8zOCyWloYWsUDs0+lWrNfeq9/4FnO3r7rN0jZtiNOWTc/fyrcJ4h/eqa0qSs/9E63
0O2yaGXB/WHrs/rtibKNXZrJYFYXkTxgWMCTPcVHUb4R4e9wSK5MLtpc+DMTXWz/v2n26a6zIOZT
Q9zs5tsz2TSgkI2HjQuxU6FgcepN8Oxor+FOyuSebZbDUrMtMK5JTSxKZzAliCWKJp4DOLp3q0Zq
FdtiUrdJwhQq8qAjq2QdecxDFrFiCxevSI3bHoqu5xh3PHgyhnGQlpPT0bo8abYz8NAz0AsOO7N7
xE3KqO5aPLvv8I8n4A2r4rb4ZBqoLns4f5oC+k5I0RziuGq2DBZmdkpKvyL9u1/nngJGvpiHMwsP
B+f9KncfhcIG8tDYDI9sjjEJa4BCocA23WD0/u9c5eGUzKyEbsDTXEG5Oz5QIOvl2c94DXhvaeAS
D9VkJ+UQTknvhKi6RbuoJcIsaOLjutCx1cEfrjTB3Ydpi6WSpStDI6uHN86w5wfDu8lW6cyXBxMa
YQvsr8SrQn1J9KtOoffAC1PQeD0YzNJL9jYhPXnQckSaOzk3sSWFI82BWWBlaqOcg/mM3p99KYL1
rjcrsWe15DwQjkznMUJ6WDGglYluD3vpj/+qK92f8RHrmB3Oindhe/sI5Hz62X9msB2igfO+Owxp
mwX0Xzqw791g6n0Og4ESvdB23iJBO3xTodFxFEi6B7wM5uxcGjwBqFK3mJ/JoJCc93DtNthkkWXt
B8umZ53hNm9sWK7cG/S0w0ihwfNpAH48P7VmSzGUAPh+wR0eQmm4i1Ty1Hn2tcef3pL3xnQHjxtH
t2/BycLMBRibfcviqyMRgAQlxtrXWLcd8bIU7hyoPAYNztUpj0L7wqk9nrxZfe9MNDkpy4gP+1Wh
j3P0aH60dsIgbEqtg3OIE+hz6aJGERllp3MZUIofGYXZ7LVe6mXu/Rj1J3fWnjQmZQyiFqa1I0vu
IBOqK3e9SxVL34fb/JHHh5oc0DDXAeeLltBOeZi6p7l4sw9xTbm70fYTcopd+WGeaqWDoZ/vklMD
mhxPOlC5cBuvWKsCdvJij1KHY9J3hknjcfRlxW04oT3qLfirrEA7w8j1C+ZRKZ576vHreazB8tW3
ctXjLIsOG+J0IEfld/oiF7Ds9Bxja9GSVVVauxL9N748FA/uiq6mcuCTiXlcxTIHN7ZrDcat5kIu
SSVU6yWIH6gXsBaOCO4z64rACGY6FYZggqnNLgeeKgQNwozTLbKIzkji/fHh/o9LUp0YpNO5EsKp
sX2mbpz7YratIq7bSJWEBwd04Vg8t+mKxf69mQ8yDLg0oBOY8mOlgd9xi89i75RMRN3PGKDExY/Z
dL8Ni3R4g1f7REuh5Hjkt83w7W0MXgZsUgQu1QrGLrAXYoe0IyFmeIYIgIsOmwAYoorXyFLD8rD7
G3wKeLwuVUErwGranfUp/Z3NwE2C7prL/DN0isXTnMrAsjFJwcJG2u23DhgqjMohxyQOT4pJU6T1
nS7tj5jQuZe9zGUnFDY5WyMZmokpFsYXCtmj3LFX0X9Uz5php+6PlAI+xQtiIp/FT0KmY0mJlKax
fbyO0qBKOAionPr6Xm4RSZPCNtGhWIbNjGaZtcuQ6KGwKvp9zOgeC6FO11mTemnJrSnTGZTZZMHn
NwBOldEs93tqX6oEE7GKe7Wyi2kM6DvVvmzwr+PRNhJnwosUJwtWwtYyt1IkegU7VVn993Pbhygc
LR/BbgndCvbt9NBTLjorkfexzbHjA+sTyT/gAjsM+Pf/MRGUWwAVVwP4Y1S4yrBgJBLLLVQIzuuR
ieS8CfU+8+ikmXQyaMlFwbfonCwMjfHeQGnCSRYccUA7C9fcT1LydshZD9Mx8Xr3C3kKaCTUbfBV
SsR4wyDr51Z3ploKtMo1amsWLDZ/Qg0mHXY5dfUq981ybv3+drB2cdmRA41NfDewe4wGMoBdk52h
Awmw9ZVAEh4PIcfd6VTBXYvppcL/TsuS1RH1DoS27atkEvaylOsDUJKKgPSYviIr8Sy6XCl3nyx2
vzlVysmBzkjN4G2z1m7u5kePik1/hLf3E7ToBex4wE1HPtuWf32dkzMPA8Y563IUr5+uJAqJygGI
zItGbP7tP1hxOzJuAagBKNJT/EsniY+D+P8du0dCkeNOfIUIPZND01Tvj64uOCIr69EpN/SAvrIq
lny5LFQAAxTJ93wFbKLeK+faJ3G/3WdZLUxAC4Ua8C12DtlBN1E9QYyFwjPXDtZzwz6cA34+hszR
3MuvV3uF7A6buTk5lEQZ+K8PSQI9zu+Alf6MsRnk2Zkui+HpiF7cw811RDG9zPBTAK9sluL9VoFs
g2/f9f8E1hsl9GnqKYv2VdTXfxSW2P9eoEX4LxkgPT2yx5Fwq9sOOXiqEJbJT9yrxZUQzHzkMeQB
TnvDFQgU5vYwg6EgUi2SP2dwgLP6MAuaHpxwj2o8t2PJs3z/dpTo//GKUaNPPXpFDM8al0mNBeVQ
h/4GoSOIqitF6UYv9+qvPZO7yYA3kL5CUqsNJ0cEZNME9grKTLBSN4LqwAZUfwBkzo3ifh0Y+jgy
/DT23irq0HZQMlqHsJLJAQY8n6lU1Fs9paJABbglum+xemVh/tBF0LA6NAgQn5yrrAVlXG3oR00G
3dNHEYmlZyRWSSOgeba7B9Q2XVrkUzNGLUaMDmdYfyAJgG/4SoHPbCy/KzkhYFAdGx8DmsfwiHXe
QsNB0vtidWvynKVAp5kWm4VQiuik39+GNNNPUKNRBv0c367E7E07qtIhs1ksDkRtO2EqOTuU3DCO
E7CRhueV4s+2/5yKmPrIK6w9Joe+HOVQu6jmIr4aH0CzTYK2ltCuAdcSoRGtB1jmc408a2I//iE6
XTH8BUGvxvn1mNRz2+4dKm4LRsojgm6TnXeKS2nnLgrHY9ufGoBjWkRd902uBosFEHei6kPgkhnA
8858EiWOuFllqKYL5CLccQyKJq4lkJNbTBfpea2/18Y0ELRYczMXCmoofb/+XmMqBsdeJ4DNDMjp
eaThxzEoaLS6UG2mkmkFX21zC5ZJ19V4HjGTYNFnw07BScpK9Ay9rdQE+UWHYn4NC6PCPRD9WVzH
6eDD4xYzmhg0Kh/uSqN7rLru6T667bKxY5xT5SMrowojz9p/4Wa4YH0F0xyZCzm6Eh54fTLz4rcG
LBwcYQ1AJZeYn8zBt4HfWvBfPVSrN8Z2BGk1mKWCFcc6zSoweivp8zZy/EdOoB3sx/6aGiJlixV9
Qhdqxt9Gx72l9PPiQ853k8JlxOCBmhtBMyOdaFnocrzUw5r2Ybohl8Py85psN+K0CFUev13bM9Ao
+bg1oRb+G5tWyeJM1mgFZmBhw0HLani71VfpFKX+l5TOQtVEyfWCSmPdhSVvdcM/AMgnXNXmHlHq
cmWhrgSdCPRpHq+cpZGYL/a75EE1Te1LpQC6RCbZSPG1OIEIdttAAQd73b7oXFGbYXxt4bNYYjug
7ApEx3ozhAbTkeWPetfNHpPYed3dWcLt9vi4l7+5YWY6h61753pHdWwAiKrlUzeP+Y6xLFP8xsbF
RzOxNJZIeDocJvM1JPpbGEanJY1daL5ragEOPHbt6OWuYgqqWe4IaW6TrhA7MvsseY5/sUy2c7WB
jF8j4FwvbCioKmmlcyB5+7yzyr4fM7yASzotymL+31pljciJqZqd+vpfCt17AiSm2q437i4qjMbu
kz0rOTY95F+DSeZ3W7jogBf+bEk2brYG2uGcnDL/ZbsEyJJJq43KaFfLBtBqjNy3TXofCdj4FKj5
8h9h0sGVfd3EeLLGx8NVYt5hprjJZh69jJP3gxcCWJqTtZBl5jrbvl46OU+VyjLQLW1RloZHxkL0
WFOq1V56aVljasTVICtoFP8wnYsAV73WMpH/uqhtMOFf3FsM6kE9joBhE5QVTsgIfpofs7D72bBG
PkiFVXkw/OV2ueysE95HEa8cVmGcV8IPQbCT9xXo16ZcyZkhIkdzXJR6G0iTC0WGiitYBmeqnjhv
qLy81VI35MwJFJr3m+IM72/3ECoi/ooUFM76o5tjhLD3xtKoBW14L6Fkw/tvZr433ENNJJquWPqP
J4lT3TqisRXqJxDJOpQD3qB6arZknFLoHNOnzOWyGQpF1cmR73448hiW/Evq1FjgzVf3++1eE4rF
hFqLVOCUfM2x1CixYdQeQC7a/GUNX/QG2ntmffHDagFBlWp3Ak0nU6xdPuMAUAeDkk/L0svguuD1
X4s65Yz8pNQBygG230B5QMWwWkFRwiIaknG0jok6jU5MPXg6dx9JHbcKoCMlttNfaDl6kA5ggkWY
Z0ZLMOyus0V47s5mWs9LW+6UWfsNERLAxdpmtuIcIxosHhMn9p9iCjJsUdjYvmFTbeY+P9ydGTgN
Tt/0s39chqJCvp2h7vG9RZZKf6IjmYidvlAyto1w1K23XJQxSKUM3hG904kcUM3WxC/r1TpwsX1/
exynd5znX0y90Oac9xi6OToZrCaee6JLrIRXk2+fwCFG6UzFZSHSsCctwOtsFDW/lSzxATkM+iBK
nE1WXGXX3zxgTtsA42d3QlN4Vnb/k88UaH/i2LdxJR/lbau0RKLvgbO5tcXav06GT+TdWCi63cBg
b5rxEiHMdVvLwPDtjh7lssUtmYXW8LzuM0M4mIhlIjNSxL7naIANuktUuRWKy8IL+qQpogJ9MpLN
aj+f9LRCkSUv0hgWvRpvp8rAZrK7Jn30kB+atgRh4luM1ARoiJy5upT+fwrOyiguRh2VW9Eo6ekt
wCrXTFMVSaGgiBjaarG5/+lMC//VhB/lFV/5z5HjgytCD1yqZEHNJHVfhGg/gbFtEN2+jihDi9yk
w+ANuP4i587d92pz5nd3sjz6YYDgWxkLweXwtEvd2csgZs4hd1O2/oUtApQHRUYxK3t9R94ivtPg
zerW6WzeN87G6a1NNewq0IqR2LiXJ3EeAhSlrb07qsgQ5enyt13mycnkuZ/m1u+6d78AZKS+PDf5
W+LOgwDrZpnkvuHn4JpZ9FYybBSaXH/Bu8MNExMjn2FVGulMwYTSWhJebX053bemE+DUoSBbl/Xu
dqtWGFWVYHkL7+ZmmXYtOxe/5RGEvToo8v8ywX/VZw91YCtUQO/L+1EdMal/jvo407VLWYhyWCkd
u0xhm9yEQZ5rDqbU+614cygu4vO+AWwCk4BIooXS9aMKAguUXAcuVJ3tTvzrdc/xMAzs3BfGlP96
7IJAgyru3Wd2gepkHvhIIJLcrR1IgnMlGFELdR6+m6bc0TU1Zsd5yz6mBSFc1xtUtg1C1dS4jXiX
KmqMa/iIANqxjllYQ63j+VdkwPfsgMRNoMCR9aOKboI7mZaiafPCtfDeO+OGqj1HcdnaxRMJopdZ
zlMIgr3OenFpNcJ184Zo9EWaVov0P/0Y9gMQXFNVjBODc0Y9R+cjg1+hqFw0C+RrOyQ7EBbfUKRe
SF8sube3UyT17Ql+inw2UI5VBr0AxCrlJfaVQizT+RVdX45MRu4f0TSX3Asi9KtViEr1reRfW3QZ
aIslQhQxt7lvovL/fv2q9pLErBYtW79ZtsRxAu0mvFEWqqHFFpaHRF+SjYMvJnlACqXEV6lNCIYe
90wVKf0l6NVnJsy5gI26ZPw1Z48dhUKS3g0aCIn6v008DV5LYFhQvkUuOCwtCLJSr6Vihpjt20dM
frnQ4n82wqw1FKRLX+M5vJhcpxXwCiPxAoVcg+vsV7JWgt0L3CACEw30T5zJ8DOuM7frRg8/Iufj
64Cc3ALOGkVlwICDIHjEVk9ZXF+tzDJBGMCsGYQVZ7IXwahRd0NsecpGRqcmHOzWENkvEtQGpCIc
4I2YAajTHzl6GiPlonJe4wuPICEY3DZvr7ude35F0CCAe+KphT/2grU+1gzBsFUypPKTL5mBU2or
YmRAGgBjYVAf5GiFvX4GAzYlcVXFfpUCy+lXI77jcnpWwlC29ksRYfo+SHOC0jsqN30UG9zQJEvo
Vbh3yiy68jrBbYBYTt1sSNwxawI3LdzXyll91RkaEGgGGgPVjQkYZuB5dYPM7KBOYJmwdk+XpIdR
WHDQ5qOVuoY3otKOb362tf1vcTPf044C6nSte2maxLG7Bb3SSXStCbo0/D0mQkVp11eIK9a6704R
omX+cLYvtzLaZuNURGcahQUw30biHFCGeOnljUC3cmisCmckMiQIui68/yiqCdMlJP6kvU40qqAW
9eEdatLnZjnKGlIBAFj3/V6PQxYEjA3JcTvn0ul3KbvDQPNtUwXSkptm24O+cP6HtIBsvQe03CxV
1s1DPe/eO/3O5dZojNFKGRsxKzxJJ5gH4czYvMvov37ViKFWguZPF3j7b8Zy3LdJMIhuO60e1fi0
F9dWUcF43y1TVNxd7A6yp9FYJpL6rbmn0yTvWyPRLswskvv66BYot+H8xo1vqfwkG4MBxIvQALIm
XAEWmqQ3TlAKePfvKobjtHJkE73W3l4nArCTJrO9gzelDCgJ2XaEI7mIHs3o+ljqYMN9oBkQb2+0
BNYXEWEaPoehPr1fyQ+ADHSA6jaAvRMqyhcdQ2wEt40Lbdvp/3P1wWoS9PXNSCYSuyuBKn6X07CT
JcggmGiTgQYoqyL7qK/Nm1sGTpSSALhbKgYVgUjbDM9oGzrcQil2m/G6ILmP7s5e6PeDpIjUyTLP
RrwNTl6LkLFXFMy7EP9MqyL7quGD6Ly1kKfuLC8Dho869IwVp5z6shQZrptMb+JxerQjVoMqUWGn
sp30c+M74OhNSDTQJDZGp+BuUizFkZsXo1pUo4xvfOMSzbbOlWLS1ocsHkzyS3j1pxA59O3h9o7W
OLqizGSGIY4PaTFMgqCtfkEEyZIZkuOqwQmc4wRdATPyfFP3Kkrs1OC9BSARVsZfYyPIhZwNw5c6
fpn57sdqL5c8mXvs4uPUTZVkbBdR18kdxRT1k39xTqzNmUZorRSu2h6p2k7GJ9L/60VYKymScarp
goCjPBLhAAOUc3U3JHdsW7QpG04yk1uZUR3WEuFNdqyZ2TMrt8PimjpePTYPDdntOokGZoaTyKcU
pmATWsXXOTfYz4vIg30ekHnElLhPGyYaMqNfg6RAFOZNKfareEnvD5kw0jEROh6bIJb11BQMZj3l
gp8RJvj2ccaFq7Gd+8kBfS5Fl8RYnDRYZz0qtIWibHZWg8RXOpKpCs/8BRR7GwoGa6lw+8Ap5/Ml
+Xgyw65rGG8D7k6c2tZhua2bgWBI8OAhX7mcZjVXGB3Xcd7OSyzVaseBBUIyd5q0pVxQdUjhUkM7
ag0tIQcyRk6tMh5GQljfNoJ7lv3XnUvqJsvyCLA+2iCK/foGRRWZfeGzPF/5gFQDd/GtIJN2QkQB
amu9mZ5rHudrXkznyaPU3AjJ4E4nztR9ub4Y2sfhtam2bg8VRpaiWGhpdXyGoBeekY07eBpV22Xj
QDR1SjGkYVmPoPC2PH01NPKTteM3SmLJGijJ8RK9CHXWZwMPzgrQAaqLfI5rk1+VodioLzXWtZAg
29Tt490f/IocPeEb/Vf7UTX/Bls7fLbV33K1q62gUf2LtnI3RA1DHUcIuVfuO3d0WNnGq2vmrdj9
xIR+0YPVeYHTdF6OL+nVVSmQpCTfGK8pj9QJqh0NmMxHozFHQ/WtcAXPVa/e6dRi3QGWBSvtLVNW
A0g73RSLcXPexM0mwaPBuUh12vv+yx4q8pkZg2mbwTnJAXb8zYS9zCKrDIDOAptc/QtFswT/3x85
ctFjErQFniTO5wb7Gy5a40pVvkggyCo2M7sl1TDz6OZYS+38ARFQMfFY1HlBMckqLIUa702ParR0
b9YcQCbMge9o0b/29ZYWh7FpKI79HV3rzQYI+Pdso2UETotSyfxUu5QYXMOTZr5IhtfJovfxJ9aw
yu3CSXblGBwbApvkB1Ff2cl/YQTgdOyKXp1jOtDe0yjUtF+pKPlMBBaNAgOCwaHaOZaQR5ifxwQT
3LrbI8gt1Uoy/Q/qLjAi9Qyq37/NR91WIsAIzeKFSoyK+TUk5q120sFiWxu/NlgluBTvHsWhJRqA
EZOusKyDYj03TCQ+2B2smX1YrA24zI/GmzHo52Ix/mQn7BxDw5xJqScg3zEq/Q3zJ1MTYlt+dMiO
cUnsZ8f+AsfpbasYV2a5M8+drh3veg5Gz7Tzmex8QWpsUo0/XWckf3RQh2Y+3yr8r8e1yFLn8keF
QL3hDtsDJB6KqqlGkh6P1u7JcHiqJ9/rhJtpdDGDthbOtUzBPIB9IKKWBmxKHqRnA25Qadx+rqSR
RW+GoEW6azT5qoileXL17TuvcUqRiqG5JeHFsQF+ppxy67ifQIHQU7t5yZy72Fb8L0ZMgUtsB/zi
/6DAfYeJfG8RU+C75vVxac/azeWzTcfFj/BFUUlqJu1qdZBqKU/d8PTUD+a6vRwPitJRjbordxqk
LFJnDtY2Exf3i49M4TWpr95YePgg04yQlm+qkvM6OMi9xTK/vXjlGFNYgB2BF3L29E+/KKSTXpIA
aiwKS/VPiGimd4ZSrFBMBZOr9IG3WxNFvn9VhmVsVNkAGWMHG+3Q35mJR4y0lGcOtqzb8uAlTnU1
81122AakGm0KNpF6We11Ggeolqrkzi/UfjRXkH2Ng2ym7AM2oeiNqMcqiIeu2eezYamaL3UirP1l
dDR49eXIFdrhomv1+CNBM2+PbVX2dDr/QGrhj3R1OgJukSJ+NpLbzv9+hqJCOFOvF6/uzLPVpglN
EWXy1BT6fqGpPlvfi67TJa0UOnqz89z06gHCnPmJP29+4DU8/T7fqgmMuKfncqTPXqG0+pEn6DfB
LNgTW+KQW6HQ59nHuCbncNdEAy+QqFdYrLUfGcHKjdSuQqTH0yP5Wo7N1RH72nnj7nbX+L4U65w4
Ku8lkAyZwDTZxN5l/yOoFp7w6Rus2c853vzZjZGERXFDOleKTBpJvfRue0p9S5q8bYc6W4dUACEj
Brhbd9LaWHKxovRVVn0RdmTlJb//HZLXNlkFGvJY63EdlrYLTo8ICIFpFUGxtht/U7Pg3t2ENwLu
KEP/5h7qbiPxz3Uo2zNWtDEaLSU5474PL8omGBJIaqc0rTFacJsKa+hDQP0NlOfwUyrx/3hhgTsH
dH9RrizyetG9AaOomYpovKYVficsiUxZzP1ogb6RONgVzQ/pXTfOHST55mCwHmo3Dh2hAg0mX0IU
gtcZj9s0BvcAKvTslsfbQIkc/11LRHuC9WNDzgNyjvMRUVX3pK+dj25JhTcaa+7EbFPRumomMyAd
bu+f35YQCNRMxl1o0GArcZh21IMmEUH4UR1sbZJX3ew/5gn0eBX6WYos4r8pCYgqTenifZT0M7B0
uVpUhUaOO7r4H5BCYS4y7t0AAjccrUA31srEsZfqdb0JcqLobvAQ37YDCgKq8i3I+TGl5YYLHzBX
YiCa8NnO6twGEntDPBCTeS0UIiB7X+dpDa5PBGSKHZ/Zs89brCr+IeqSSaHFlhXjmjmjfJalzEpM
geAtRDaHrja7OrA/Hlon+bXs+ipxy5eQAUYsYltRuyIvD1RNO//MZmz4ilC47HXLTuC2NP271gTs
5cAuZIJYn27vfvPv3mC/ZZsS/gztaA5FGeZYm4JAkbuqH2AOGm5UNl7IhU10aNXATRF66Rj7Guup
m6bEoS4ME2BDHWj65uu5Rf0I8QlE8mzbviKYsTNdobCQyQd9E69MvyVg0rkQcbLOZ3Uk/WUJVNf2
7VNygFFvmcmH/sB2oY5bw3mRkG4jggJGgagaVyLU1Ek4BC4YNJgPwrmi0xb37LfFtaQelOIf1s6G
BoY3H0lW5CQQQEQxCUEKh9+8NvVf8c2kKaot7WhALLce1VAyFJbOOxXNgIRyIArydPF1TjlNcBbO
uwBIUjlI7ZQl5NqAKyRL+80z7MQLtfHtnAy1jB6bhwEutTJdCoqGSuTF0AaOLPkm2XfY/d/o126y
c6FUq3eK3tyq4vGp6c/oScVzQ5Yidm/J1rrWf9bY0pk957FULuygTvvmOAB+CRueEqWj1r2u41EM
mewa0DQR16xfC/Xl/57GqaAvcPKidSnfG+A3GfFaWaJU0Rvr5+2Gyny9PzN60rxc9YxGQBBqzDGk
8glXeaBWAjayzoKoeRxmAMhn159nD00SkkbNUSToMKzbf4pmKh/daizWGC9N8louCun7I6kPa+07
1coRkTslE4kMDGXBbVqUytpby354scsOSoxt0o24kn9rh3EkNlA9Hp+jBT5geo0OC+fFwbpp1Tnn
FO6DV0kzWszaJg2QXFrWoUQ3H6fw2QiDkp80yXDhhdFTCApRwHxUt78KmArvhLWfvpomz74xI8+e
VKLXlncFwT1MPr7tFBiPpPutSL1AACJuswM21N0h6SHBmolspdBmWEwBANCamVlfV5utCUpAdFfY
n1TxkwOKDrJ88GKouNTvwNBi4DhVdREO+vAaClkUQ1pBf+GJqDWRdCaYRpznzI36MZXM8y+PJ8sr
rn8O05m4KQj9dxvE7YuLhG6c//8Rbyve2kEdfIRV4QwULXeXjwmxQDRtLKk4b+82k42HIGJo78uj
YkdS6tsNr2yCO3Xhz7/om+rYv9/iAlLwbA6dGzIyxMbsB7uQhLpYd4n6szXYdJpummzlSJ6h+c05
1bJpC9qHwaQMk4zoCJk6BzvBQerbDE0kiX6ES7B7O2D0zi6sIzYoIWUPzMKXvpbGFtc779UM8rAJ
eiEZQfI9gcN9Hd31kj4E9wabTSlMJvijgYaWbe2RCmNl6m27VXsU3BAk8QrTq3E5qL/m+1ezoc4y
eSGHVg/G53AmxWJXOzKUcwzOMMBLGRb5wOM5FFd81kjrm81xWNCJ86g5Y0Z69AvypH9ewlaqolZI
nSPyzOk/Es+ZZjDlqmz8wmxoKITx8JJwWKyhDNyFfS7go9ImvOO7Ff4vyJ9QwX4pEqBE8pxHDeXM
8ujW0pBLiBm8xyli00+SviYvgcWg1B1msya6c/KavUG2Wn1iPPlVAy4on/Ts/XamK7Dghyhg1V2Q
+ldPiZ34H3q+qRZWe8kLcy1L0v+ItKeLdyaKsyXkcbzxxYJTb5KKHMV7HtLEd+nNyVgX0akApGR4
GrSqnYcArbUsUlod8wSYU8/CxI6MNLFmmK4fHAE8NxWZggykJcpA7+q6qxgBAk+efsWQewiWJLYn
ooPe6gbeNoyCI0maDEUcKeRdpgVdO6BRvwqGVR56zRgfL2JobhUbawMVr9eAEWY0lGdPKWvyp3vc
BcHX7ScfDAaSiCRdPfVqguMeFFap4uBjlflnpVDhgEn+zduFezvSOhX3H9gbVkBhT1l1FY1kUhMb
9BYYhCxrWiPPAPHeHwo0jid6+i3KMpEzng/oYW7HTxQoFdTEVD2zi2ond7DVEpCH83tAyFPjablc
zOQTU1+BOz69FrNzh3v6c1PBB5f7grkvW0f43fW9AhdmFUf8Wy5HjjK5IdmYmYvvx/ITt+I2mQc1
c/eXPfJiEq+dFUWbQ2gvkEkVMO2Xmqlj6ZR7QaL3RBREC/sUPy/+/yGnU3Zghg6yOcWd3NB3n4yr
D57fmB61oBeUsqAQIyF59cU0JAUnyjFeKO8/BfQ8jRLeEcFW3yonPCbgPEaJ1mhslJ8Ka8ps13i+
0AIbjiJIjp5gQwOe2sa2SxiJFREILKIrAiBbb7GkL+MlhpmXw9NjszUtRaVoNqkBrygUc/vcPzYu
t3RNo1ieyYQcLX4G0vWQrytF9J8zrvcbdbcD8JIkwSHfGlmifYR+ZcQRd/07hV5iHI9pR0tF78OG
stHXiPXIWmOjWjJ86OAsGXl3wmiF8N+J16rQq+9XYIC2Lbwl1G6UV9CHGmogynVa1nqvm7zXQwTW
Swla/uBVA38l98byX6aFZoY22oh61Tpwgc9a/oyYkduF9qUm7ZrswXaHe4ZBN/5sk+WXJmYhGMrW
Bm7ebOSAa01Cluzfwa+HCyYN1YvBzg4YT725Nt8DD9RRuJdpjMSc9a1sJDd1EAKphqVDPWvfAiAs
dgr74K2JD+cg/mlHl01YKvvKLY7SIK8vQINRGIQeRk2gA5jwrAYnEMhwX8i3enPcanD4o2CeeY6M
+rVWWHsoXsi/4M37wvwlaBg6L0iQrB6qjESqDZcjsJMbODR86+9OUNF7EjSb5Dbw4Hg9z1Mks4g/
sKSSyswEJZmHo7kohNRhmOz9mvd6lzQnvaiY0a/f9mW48A3AGr6T3Nqp63UK+B3StUJ0as43k/v4
0jbAL57lWXAwtI/1h73AqPYAsmHEQk757MlW74mPGOXaQnLmO30OY0ys6t4R/Yqghm5Rpi2wwILa
Vky+mTs/WI11FA5lD+Bq735+Yvejl0PyjPUyohKiI4orlhNYHkl4YyK4XsS6FNnX4c89WQ87OK02
UQnrteCgg4VFkTQOKYl1qvvIGWaSQAaRTdpcgz5X6VE3wcBQtGiya6O46v0o+ATrhhO6d4YTfFhh
dfDB/OUjQpNY7DcZ14yVwTCfdLJUsAU3JhiSibkCeaZMHjK5dsboVr5QQW6DlUOW9fKiFAqAIy+i
sD/sv9EL/AhmGqvXEM1DgzNMiigVuX9nZnZaXSWYUqbt0Cfct58jkHC7QMsYVeCaRcVkpb+Ci85M
JBAGvIsOSM+GIYEqJK5TKE7jH4RpdkrX8jQaBxdyxoG1DjAoRDwXE/6H3ly1MNnKwfsW2Ta+QYIe
PYC7jZhnQFRM1Ern4MtAYk3rSRivQyt3JlOAvpM4KW7Ojzm2ic6ZkQXNOgHxC78zeL/p+uBfLTee
Gu4vQiLttssAlw1D52ORrbvPNQoN4ZtIxeY/3UIK58a3XV8Zbi577Rz3oXVtdi2Rbe+yHBsEiwcH
yqiXl0bH19MEq0BUqz2AqDI7Ad+M7XvS4kadaX1LqGTlbUCqF8vaR51emW+9J8Fd0roAeGR+rB9C
O2ELZUYQP59IZ18kXHRSnRMDM6f4+/IDbaQp2GSPSNRBP/GikaPizTMNFyJnpx6zE3xmFl74xahF
yoSqxK7+N/iICQe7/fsAimJAOoqmdMqAZAblXFDCaPhPx84gcFUC9LBjveOLwPnZTc6IXRtVqLag
6IrhI3IKIUIV6x5SMemVcdRUsA0owiU3jhGh7Rh2fU3vxoBIlwtuoYp0+Ck8ziqf/M/AWN5OgVCn
n7WwDQTRCG9wkH+hU0VzFrHTk1JsEbx5sGEWDu4Wwj24QtY3jTZvzuKioLjQZx8SG9RnA7ueTRS9
tthuGr/ChY/H61Odb7D2qaB2l54EKVbfTkwSpMUqxGRt0EXJIFgAhtXRP3sCiTpucdgzeQr6Sf4b
/Gns2D1DA7nRrwTCWdytbbWba7ghPEO8QqSdb+iSR16sqlvu4NqqfHVefonIfVacONe8CJYY/ABT
AcEdOyYTVOzDnUMnGRwRv58O9A/F1kid4UbweniUJvDK2hYdCFH1uWgYd/2sJFmnHpSTpJaFIyxq
bKXy85QTB/+ZbyaARfJn94YLimA0l17k80ob9kYQzqOxVtYCcm05ipgmfkCTzn9RqMLgoToatRN2
+yUofL7mbXJ4JEzrv0ZdW3V0Y8Xs2S5WzUsaTXqG+CIEimg4Qp/eBDsmNs1d9ZpX4kr0jKNgVDm5
y7BJAImPjAPy5oUFz0PrzXDH949FvmxOItm6oztoC+JvcCfvFFVOzPB8Wcwnm9W+NYFaWGuyBXrm
A+ankKGUTSKM1mxE9w5s/DHMjyp5GyNDRDyIvGCZ5EF7o5mF3FfakVb2kuQ810hoB5rIEiugxOo7
6AITsFvHeRvnwW+tPTbBAQ4LPoRgFnUcwk0oCP/9rRPsr6wAElMzo5fu7qtgoP0/RzstBhNg2NZz
UpwMUQMW5MfUTCInFds+pOJ0SCiYd5iuGPMNhFKqP0rOOiIBAyJWDTzu0jN6tK2s6AF+76qePDjK
/0NOb+ydW3g6FlrS8wEYUCxMAb0iCrdLhnhVnND80+Enc/e5rHcLBm2VR+REvGmbEiZWbDXDRzC8
pZcYBTEFgcMYcEYjDQwtr+/5hTYcwc27fR3f7GPmo2t6h1BbnfOvURPI6UO/hVg8cay2843QCZvN
A5W9ZEt/hxifp6nrsMK1uKq/0hCPiXXXzpZhrm6l4oPmjJNZhkm8utOYmu4iEDdY2cYsUO+KVdbr
RA9ZR44NR32qoojSwtfgE9K6rsrvFHSRa5m8I4wMPBmTvHnF8M4GGKP0ukJ1CQVbgKEtaUVaaNy+
W4At3AVuvdGcd2yONKGTx4OED5iscP40VuCwbK7tJGYWDG6YaT35Fxa328gwZKma8HWJk+HKFVip
21yJg3sRqj6waFWhM2Zft7sA3e+ZtuyAAiJJppfvWjgYuf+pUEeRjSD2k/oeKaxyzm9OqZkkcxFG
+H/zjttYVX+JgRyYHugvqKlQm5ttdLwALYFwybv2TlNOQVd+Psi9/60pj37a9W9m6RJlBWRpw9z1
AlcM4kbyTB/qN2LZsXTrRbF9H8NqaaIBEP5l1lQsdkP8SA/ys68iifSU1QMwFMEtBAENE0RuLmpE
XafaE0NUuCHTj/OB3i7ggxabjckjBu6ui0EjjY/kNN16SuZjuRBJdow9p1q3LvdADVei+yZRXUKO
lo3tjirbyEm/ih2NtqGcQl/rrQ2uGy5SXFfe2Mi+URJZi0iMbWWKE50Ze2yn/ubmssoQH7UXfFwt
eOdXopGN1C64LczeKzzFTJPY8Zo2TD9Vqg8beQjMZUfpRchmmFfnnu4oBA61RhohG+IFLoryqwd0
8HTNvRPUaTQMq4KN0Tn4NDO+aK/F2TUSKfMCy5q/YNRBFpIcawyIWkIsa4TdIKdDR1yTZxa4R2AI
SoP7ZhZqqqKBfuZgoPY8lXOUtuQEhxpA6sJhp/f1+vzkKxBs0jWdYUSu/+TwNpXUrrs40x6rdXXz
bsYVHti/m4SFJCljTOo+yiF6ElciAN5TGf28P8VmoxjFVMFddRf44dQRwR0YQ4CyJgPUn9HWpBak
XuHXOr3IZtyFYba7FvttbpuRN09XnPt5OeB9mRGte7Bf6uA563M1PA5/wb/V1UHypt4V2yz7T59L
pOOBI75+EEyJRz/gE9W+vAq/PHpvNCwzxMi5s8REdQe/LFTsKiaTbBggRLty5m+ZoQSrqT/9VdXL
3/wMlWqPTSIpAxAa/zATm0XxMSFZjKW20z//T3/13HamzD0Ho0LY5jqg8i0DbbfMphTOFmtPyXih
dLk/oOWepXL76gFpSFXargl4HPUGrPzknzGlLxFpneK52uAlATKVppMBQ1H8gzWpOM37zuNXj6/d
k62IQjJTI71hyhlqD7Eta7y4t8MesMGxnXTfdv4zP6ayU2H97skd+WBtJjc5RDCMcxciiuSsq2qh
Wo54HnChKtUfiU15hQ7n1jPzKxblV61BjLlMKiyskR9rr0KsLyY/M0IJu2OZ16ieLB5BL1yjItLE
aA11YemL+28axtHyqib3VJd0Au27FrokhQdVVy1KBhA8hhyrfAvlQAwpOrOa9aDnUkjSlQ7/AQZ/
uyHxIEeo7BQvAtGa6brCvRe5jqG5+rSEQ7e9+LOrEKMWpU6Q7K0gac238fQDjEjdQBBn8GGhIgfY
shCw7ZgrQAqBtYRxMdmtznwpAqpnRalkfvIa4O8suflxOM+eX0IMltTouqC90/qAy/4VaZEz0kSD
nz5Ggxy8FsLcCLeCF+0AnuwtQ/0xwVTgRT9NKEoso/MMhpzJ2ICUbOYcwUOJhRrW/tJNRkL3oeJt
9AyyLrU0ZvMD1NZDGsQRStrXRL3Xevs4bh+U2fgedktfbqe/e9llbVz8ATvn/eJbqSTi1/tXIxym
1ORe9rx5WKKDWXVmMe18FvFZWobuROfq3Lt6YLjEq1hLORjQmfjdcUzi7prO6oSvCWVP0ZipnSIq
lVvlgGtjgKdRW0lQYNTBLi4GVbw+ygo118eExztJiDRRrPsaq+7/ImIlB9fpwtH4GiamOEgH5Dep
FXJ4aLWmtJAw4L747aBxyljEIpbPyadj6eX5KqcvxKDmM0x2rAIkMfVI6xkXPXw7Fzjx0kMI8gv6
fO0UKdRPbkJ0dYohQtB5YTXWU0XsmJVgEVZa/1GZYwxvjgM/JQcZ3/xjhYcJ05bu+kpQtkczb5qa
H5o+PIGv9l5fyoOlsYo9r+oqagK4BqPoGut/i6jjFSPEDD5HGncLnJkUyZTG1jr2s3aig3U1no2+
ZKwZcgwES5SXIHHgNgCLX+5pHsJmnzg3Dz6vWq/gW+LI0rkR9B4F12qCEPJnMtzc+lfb1NDyEpAk
uNaGAduDdrWiTwJ9iUXfOVPqyJ0WuV64OPAwvbajBL1odEulA7uHhxP1cdtQfAuCJeb1/PdNHeAg
AuYLU0WKW3+mUVNHRs9jXi/39OFBkgytGYK1DSLhLm/Xy18nb+RwQqWG+6RfG3MiHVLPND0JyMAS
Ui3ECyRlMjp/IQ4rTUpByBRcm1JJuPS41ftyM8d/EKbGFVyDgvULCwBnLIq7znR+onjZIgYNUefm
ZJr2K+jwnT46Ydnj0pL+hZke8OcJFbxVfQlIzLOA/YfsskSabLkA0XKkUmUQUslbQe9W8uMRg5Eh
AxNHIZx+fxdWay6gkW5mmDNie23R5eNvBoSwgFlvGaNoyrguo6I7dupdeYZFj+L6NdWoXDbiBAEY
raxaTnSZ1H95NgyzPX0XMA5hdA/5vaJw4/IT8ABJ09t1TdKlB+BSpFnvI6fm3hRsx7hrZql8v1zm
QI1wvOeobo+HV9syiZSk0O7eVey+Pskd0NQXx6P8Yo/VOq2BCZyJiHDUifxBwwDAbtjz2843habh
8DVkQSgqDg7LDx7si1InGt7sHpsEGbILa91J0clSmpnfsL2CueUebDAFvua63yWvcGsVPSFESPZE
kgZs0e1+ICZSHk1u79iHhuW8B2mPJatSktdqWx9YjoOO6tXDfj2UOFpRUHIJoc81YrhchfYiWcxL
jgBntsAxi6Eka3kXE+PCeQL/Oba+bOltWLpV+hFvlAGWrHfV40lT3QSVSxLfVzxJ+nWzBmEs/HfD
BjSgAiZpxcg7Eourhm+WI5H2s6YoRGiPsDcU82+BcQqiBmfbgatXwdwVa2RRJDKATEVG/xip/ZLx
kBurhVeakImwdWRxYsK47crQZzxsOVZ/eGlzpfgi8+uIgsd0poYPJjiAeS2D/ve+4WtBxhSxrC99
unbwkcXXsglKl4uFvACs8oo8K5UL96/aAin+G058xmsuQxYAEKFozZN+NZz02wmwChsKwDE654Ky
daKNKentFPyzRvYswU4rOQBMGXrkBH6pf+1W8bzbsDowlPuClrlHNje72/Atlxwuo3aNbbPRWW7F
y6C3qbBQ9riFm2iiQ4IPJ+lcw4/q1pD0E8252UC9tyMjZ97ekQGN1f17zzrJdk9EvPGdc8EsoXOp
5cbc1TlQuV9mHCZ9GSeB5PDaSv2/GQXyXQdjRp7I6o4oiJSAerxORoiMy7jb+VVf/BhooVLQbzJ8
IA3tNY0g8jKxcLmJLdEgl6WcjQxUvHKlsFUVssaNRm8Zr5ahh21KlWd9xVwejfW37DLztAse4xUV
D7nyDPHH8O4hu2n4DCAuaV+wWZbCY4ntTGvPIR0OZblIhomj7EaWD7JftQqFTduJ7ZZibozD617p
bj4u6nYII/dy+C6hjr46vEt+UcaNvXJJYDLCNJcdkxH3ROz8pz2gu9P9qqDzlHuo5EUlumxu7VIu
IiyWO97tHEyxud6hhbGLW8dpCtfJesu3SpkH1hrh/gVeveAmqD9GC/9v+lZb89MmiWMwpL22oglA
9G366sYEQoIMSWL9U1/I6YF2a0oIfILhhY4a76SE3j3D/YJQZzIK/ybBGuJgVilVRXzAswHUE4xq
PxyqwI8vFO+KpNkgyLabZdbakj9bvlGm1HuUC95c20QU7Gkv05D+wx6Ilhsccm757netuB92ZBqi
O5ZIt7QrrQma9fqOAbOjRvo1N4yzneU3Y67WxA4h2Hf4czF9JLV3fLNIAx35UnKQcVdgDI2xk86C
Vn7gt84cTxlPtzQA+St62d/dbPAawLLoKM9xDrKfUneAor2KiP7WuOppoXJyl7AxR8CYLtaR/RsW
Dle43uq1HZd9ICucMcVwRyA7vVQYyHSAXtM58DeTFvwBOXjcKg5EmnVfaktouXxHpPNdxVdAtri/
bSDceointDRWRN17DqD6DoCEJdNP3p0X3IyO0X67jgUikCphX3iiQhKO2zD+RrlfxOmNxEfHRRmi
TNQXcPCOzZBdFj+op6UlJeCuLfzs5MbIF5fdgkI1QWhXnXDBLOiOdJYWMeXKvJBlLxy2OqPi67Eb
zPpG15MLSCBCpyc90A1+0bIk1Ja4Wb6Thno9q6pguOSyMdOLJVGj9VD4uvRRZi6yP+dROAjC/PQN
gaDGtXNP+HVPch9vSTOZ5VdqrWvvml059CHhTQZkQ6pZ6ozz6qicIABgXgXD+fL2v9p25Wgx3hCI
69QivsLK3ycV5EsVzcbqpFhELCPHyPIHOQsHgAMYdCPI2qrY1vMCJJgrFLullqTtcA13cOokCV6T
rxqQkslT8ELMmoh4xUi8vf8QBfYbt6Xqx9yKs3GwVF2su048riP2q9ikLhDmCqCM2CYg+5tyL0Q4
fouRZgzQNqBwppbaUBGhXTapxiHqgYINg3kFTxsv4q2Ka5n/h8iS0FutaDnaw9VQ8R7aeIhhNr/X
RB5KiF2CQ+2xLp2VfJVPHURb8pNU1VUNdILA0J64BbvdeDv9ygkPBy5gbGu6lzXJwXmM8oKZzEVr
NNhT+4cYcbmt5C1kjFu9aAos/jIKSVwT7snEP0UMZeKJEyC9+WoNoz2BDru+mhbwT+A1XXnHopH1
wfIdbf8GHdoy06rtBJ2Xy9rVdZASLBRtgS8jHApp5IXrLfA6aXg5f5T3MJzyf4OuT/hTbGD08uI1
zMp21BwFvyIsKVyJ1yHTX5hk176OEs5Uy8OB+JxoF1bKA34BgwKVpU44iAf43iev/JyeD4mk3/3I
JaJZxpSryCB/9mXAcivFCImdUZK80g87FQRlRn2+GaP1yLVgaQodZYyu8hMZq6Vnae4zcOOfs/Bl
Ak5ibFW6aFy7DxrsUQ+avIB/oJ5mEpGifivHyL7fL6uXLUW4qf+6thJzpn+wPM7CsnESpIDLhGuB
HbeQno2v/0hyZ6339a4+zz+o24bF/YlBzzkMLc90pYx7avB5WY4c28Ho3Sgks1yrws+tRLOmy31K
pzHzsxEDTz/8Y9EywMe+I7XqG15OyQV+lb6YslcSyUTrp7d81Y3b4lgSb+KLQAm3nHhuTxa25E30
09Bkx7faD1npG/zx+SN6Zo2lMxf49TTkHhI5IR8W+EGFy+8FWO9tOrQwyz922rVyDCAYazXTP24v
sLU8NUpSTMcUEDwu6RpA7BOLy8uL5AUNMqr/sIb0apY1h1xQETwpu50Q5SGhvGcJVpSkygErjUx6
hkD4tjSpK0e7kyuhssRLIubRUzLoqvZYHF8VqMxmfbE3OuqxRVVDcEY4Wy7flCVXLOB35wEJXvT1
+92cHhjxQ54gpa4DNFa61S861Xqpr75g50Ja3PijPEy9X9yHM1DS34nWj/Ha8CDkmcrhmlllkkZQ
hpb5bg6gdgkWdBDxVt+G/t4GFuICzE4wBGmUwfY/ezWB0OathR0pW0ZBFZTs2AcZP2JETiLkSzS5
REQvWkLGe8mtnP5GkELz5I2ezi14bSt2b7odFpgxR68KU3jpCw/ZeblOlvtkxsU1mtybnpcppi0D
Q4fr+vLXpxzdMAVC1ON/4UaTmNw5EjYnNpNABPtjFNvs8ayhelyvR+YIoKdOScgC5Ust44eb2nqf
GwrodzZmTYHpArM+IsCUORoXbQokDQr7QI+2DlQvbXQdll1+P7P1hq8uGdzavyf6V+umasWXig5q
NUKtdVsbJUeKBuV5kdiH8EPiJiSZqkEsJOoi54Aki2DyqJga34iB59l7Bfu2eB1E19hjvHKLivL3
GdNWEtdi1z6mvwlklpbBxzZOstdOKILOliyPMK76loAnDT4vwZvLAN3q6EtluGw4uG1x0dVFw3Jo
bMZWFZ/FaeC3OUUlg0bq7CGDwJufJHYoMFN6JAZJWt1MBNWTLR1/NUEHhoXP4xjBjpI3Rd9FArcx
/RoAGLkcZYUcODplpgfkQWg+qyb2QC7nmZHuBvJxJkbogafT7zO960UQMwu9OkGlEAdM5VOl629m
FsD7v+kaLDAu0wJ8GlXiGRE8twTKBvIZFJHDtpBfto6hGmHjI7HmuH9PytwzmjhjJ0/SP98BYn/K
7MDLymadZ6ItltSMTFCsNpzwJLkD50x4W3n6xeITZQFse89cjhmPq7Vpji//CrjbL80JIpbifurk
zEZbdQP6iNAGXjk6yB6KwYBsgDIf7b/LDEffzppu563nOV8ptuoD09+46hx4/EmEJil90ya34Ifc
LFIjOfECnIuONteVBU3+OR3q0qKQrY0f6qfEnvYb31u5QjhssKkS2SxF5bYs2YlkcLY3h3kq4ZnO
DLrs3k+6AJKN2zMLLBTtANIzPGHw02GIyB/SFeugnU1uEQcxzxs3xBoEfeTeO1K1cHx29+dkOpVl
MuVYjvueYA5PT5WuYNr9eRI+hJeC7Tbsluqb2C26opi/4N4yNCg1R1EqjrlB8F2cscn3/+xKvMCW
FR0QOlZdtCO0QQHQ0UCo6B+pvtsFvaIx41rPNz60TRJxX4F2VjiG/kCKqYP8WFzuP+WCxu7EuaJa
YAT/KPU3a08cyW9tZ3O70kNTbaviFvdh8SlMdmy4OJK006NiZ3y1jFEUM4usQTbVTLOF4r6y0xft
gQosTa5AnNjaqsL9Qa87AXAi++s7iHvwaK6n8ghQu2Q08b6vuzIO1cBThgSOls61KQLLU9xwQOqJ
RFmvyJPMr2DDjfBlFHZCD8nTDq+Oox1CFjferoSP1145h4U8aUmn/ZGYlWQ7yoc1RmlAKBHpKTxE
I6i1YzOTBAUBXeRKMRCybpvipCUTZMPilli/noOKKXn+1z/1s+GkTkZ1x+STEWf9tONDu3rXYFqj
QJ97NpxOaE3mEUzIIuXTFygzjSAuzcEyJR4TL3sReHcu4gtWg7+NLG3ZFwUU+aWf6bI9p6vvHrsP
BsMyo5r+80pUHXk38T5UaUFOUNRqvi6ha2vCxFniCd72DFSsq3A8eEjdkM/HQhjbeCLqsZpbulZ1
kYKACKND2ypfV5qPGER1YOMIYMHjPGms/KMK7C5RYmPtvLsEzdDIThJf4L6/A+KhV+TbPt8SmpQH
GSCAa7oK58ekb2/5zzC1efXnNHXmEiGwY+lelyYt7xVra/sML3orqlLnl5rBO3hw956tPXKREv+w
B3QvZGIJ6sgpH/kytTvfVQ/w1+gmjGCgiqpajVIZk7ilaIGQm/abd6xREoA0w+pd1I1F/fbrP1sJ
IryxbR16RWv6FcFJmZHdkFHCoEjBIIIBG+Clb5JQFT00z76zO70GX1CJ7YVvBg5ZX4ftDlYAUxTM
QylvR93+wHDHaTopFfz7uUrwhpqG9fhhjJdZdLfLEK3QwPM1aqhjimoEMo1V3I/b8Hd0u81PXgLo
oTBjc7VTgjFXu5dqmAEJpi3k4TnAC9eL/eytoOeuVBSdKpxFS3Va88akrNsVlIIeum3im+HHEZ+h
dSUf1ggaz8KC5k0Osj6lpQL8E5Em/hVbw8sSxxsBv7D6n2UnS99sFS7aKcYTKN1TuV3T0pNryzl2
UR/64gvrrDfTkKgH/M9kgU1MzNcWR2+mV7GPIe1gfDfAYS5F/2D7MEkmt3TlPU23Rx7CPl2/Y2kx
qV87oONfhi9nP+S+jqSC+OvZ8A82xmopbDXqGIOTz+tv6Aq/N38Fsm57PQDH3HIRJGjTJrn3J4cH
03veuzWpx2hPfuYKGEpncvamBHCxLnR+iWPmvHO3A1iU26BP/crniaC80wK6QyJjxXqxabMGb06g
G1SHoS+mZplsT8nIlNaMqk3pqb5PUbPORD3fiKwlMv0jUvlklqBi36PVCF0bNCkDHyCtPYNkCvY0
T+DPkAGU3hCgcyGvjf9capLuA8xnOcfjrEoiemmtwmACv7N0EoOrkijuRzYJ1PYONMhzwmZqKuGT
g/HCgmF9HsjGpBsdHydfCU+lItBiGncteodwqFMyPALFdeMQpa+ZXuw4v+7osr3TUr31/3SibGj0
cZBayHzloSehXsXHDS/GUZQg3AbmhapqeYQIr1+raHsSJFiY0VsSIEv8xvIknzXrsOvzGdOnAEJs
bgFlFMtzoT6qAG6ej3DOk+ZjLeRMfPvhYFsxQjAYAKKsc5o86oDYY1xbDfvtQkhIwAk2jV1HrdIt
NrKM7dwUMQBGaL1RQiB0tEQt9WJXHnQLddBef98mhWQ+mZcdr9ikqJ9p2vGKbOMq+FL0YJ1Uup/R
l2rCnhuS2Ver4Q3xMIuaIy9wi6F+xGj4zCpb9ZByPFThixHmNpNTUCxeplCzxumQ8WgjoWsletWP
3IIVIF8n49w8gtKvP0G3aro1viBNj6avWPhEkVcMQnJQUMh+8YBy1ng3Y1xBvJMjEf07SDZrj+kT
iG3Ue3wjjYwos9jtIQiN217M5XwN8k/NZgzYJPdn2rVCxjLOtYccHwKLSiYZ3i7n1ayy7zmqam3z
pnW8ayq24PBjX4rX99a12xmEzpfQZuiR9UnTbiRipcIK57ZHbXbtRA4Dp4924taZMJvP17QB4+c5
QCkBL9cpaKVLZPTpvexCtSEspjViqPaFZYg/4bGxtIKohRk4OPC6h3EJfEFatYFZtBmXdU4xOyn8
FvYbG3sEvg14ePikkFpIzqnH6UdfdhlORNodKi5nICjibBb105Bu8v5wORtsRKkVAXzU4Oq8A/jf
ky97BHh0QmP1LdmqN+a0DFGc1kAEZo7XmF4L2JH4HW1qNi5ErUwfxRkXiwiYJKbN4HEB9QUMxZN7
SnkLkVxbRupc5uERrVTFhogumvRn3JzgivC3IplGPyjDHyQ8Zlrzt+9pukBHuClZkRDd3ndAkKDO
kZN5er6Vr2lwkLK4Cy0nLDJhZDOaiCxRL/r6B/qfyYPk3E5udraPe++J0uLFQOOW8pR3LoOi+lG9
5hOTZ1GIWrC60XYoEvmOwEAmNfl50vs+LIbIiL7xrQr67+fM8uOkZbfjcSLD1HRFqAxZViKtEi1X
K2SF/djpX/wyzUTMBe/8kIvMpOwKAF2kZKKPE2KomTrF6xfBMA0TN5wBfnYzX0Sh4r6hqFJh79Kx
8D53YtorHgTOAgcg8Eh/N9rqYyG1kOapuOICh5WzYxMOCyAT4O/Dfs+F9zeMn/8ArwZALvdvDHL9
2vHcUcZ11u54L5EIWD/ARanPLVKoyDEKjQl5klQ+oNKEMuzQwWn+HBfJK0ia2u6lLrmqxNhs5gEg
RHa1akfx6LvNfR11bAwCZeUTyjNodIXOspyl82Ox7FQfAqPSXLnxDf2taRy+mUxZaZT1DgWT6LPv
KsaIPCN1euDcSeR/Q/0GiFXNzMS8Zz+bNpzAEKRqiKVpGcya5bbx0UhW9Or+S+JO1196qZ6KPyz3
Eh5EhVgv1DcvQmH4QQ3M1jN71r9yKL48KomjoXCo7G+17N5vjdt40rljy1lVnrZ6keqo71gnM/8J
tEPzOY0OK3/su6lnLqXG4m18tM4J2jGH+DhPwyT1WWlSUrfcnMvv108e01c2h6xoDJLX7FxUyh1R
jchbHLXZv60asHdiNMEQc/5dbK/g6AVSM9EnzApqHKYFRqqUFp15TMYP14nPyrOKw4JMiWQVI05z
Zy70JjIssbnfMC2AfkAqOG9VW/fskmz7FakH/4CG779yHBPaTSEPIbId7pxLGfugUJMypYMfDmzG
OKd+zJkkGuQiyFnx50FI7xVh1z9BVko64l+yM2tzNVzqCjkQ+8RijoZangiY6oyP9NRwDTi94o67
x823JKus+gk1/5NxW83aDwsUDRlVvqEFUO3Epl1eTKnUBPitjwqjiziWiu8Rio4oJCSODvMHJkdY
3mz+CvgFHwtR13Mxf3gcaz0NHTxkQ3VLEq0mDXPcFSNqb/EGUxcsiUO8Tu5Q9cZMqRMN6Y2Trqrk
QFSNu4x183sKJXM5UoH7wlsKh3iWdcbLspPhqGGcOQsnpMUCWFQHT4TQDsNPt0uO2B0z3H8B3hun
W9liCjEcxo2OX9zSMsE8vYZo46TvXPnLAg+kc9/ZN+lBhCAziTGe5fuxYl0EPXj7kNViYlaOf6VJ
w+IFKHXAgtxUfmpkAZBK0/kyhehfF/hwB9w86AVxoTa6e/9dGj0qmAAlkzP3OJ8QICtmgy9qTviN
/Uv7Egd0FXy/q1AAaGXiES19aI0YfQXdp/P3dzmHw15s5DbSs3iOHtCA3nD44HKoQQMSWz5GbbO5
HxD9y3hdgd0am5jOM2V+Y/X5anXqwmxE8D6yBrAioFga1Z6pgzq2eaEPSAIPdbAz4bYjk8xBEE3f
UwYlJh12FdpChamGVFJgn3RCwOnzxpTCDfDGPiZJzIWbhEctVD3fQlqN1C/gTkO6RxGBsYApHV9b
PN2Hpv6nA96zqPUG7JMGqO2+6vb/XEWo+bGdfExqGkK5iqSA4tifhdl7+oHmYcDrTYOvnLZ/H6+P
q6vVH33C8bo1L/Zpub1s0r1bCeseh0w1rpi47B4uU2fkkgmrCJEJSa8Zg75AtBL5su0/I7mGJG42
hSNKdFQVGYlyC9zc5iuJD/EvjxE0RzMLQUFpp1WlmVFDFpRBnvdGraWc4S6wm58EhC3F/o9zjRvY
LEXMJOB5tguUJTNQj6WFKrJIPRYOUdFXbxRVL58qmYHoaTB3IVjAxe1nklc4TVfZUwD0uXjTpSEu
cfbNzkItj8icZl5rOj1oTBriyxGczObNTGWIsUkdMJ+uFxy/AGZyAAqszWgXEZpwV4mifMZ690oH
ZER2CQp68DgmDogBJfmGIowxtjXcgKHsT7STCCZtLhLBaRZw23Vy8+OkHQyUCjzVhCoVg18vSeVe
NCiYInh1venIN8Sm/gU7UcP/D+uYquYyUbxQZ9iJW2c6S1X+9tBy8DJLRUGMNIKpLQMnRG4rMxnu
92qWPWdmvXpMiswkZGNXfmA3JEnjmpWI9W3d3DEHR31KMhLxdOP/dxcKZoBrAZ3aSEqj4wS6fK/c
OciAMR3Lia01dC5nw7DMr+j1eA5GReRvFlkRCSld/i6c0iDceayiv++r6A062XrYZ8R1jxU07IJp
8rIG3ENTJMk9p8vw1YSQR+HqSLA3iLx/U8nAax6w91gm7qWk11UlybM2pGA3Kxl0wrUd8JStCyAV
eSvVdT26TlfWPRX4Br9auycO9khw5LfBG7BZj3iO5lGwnVL3L83AjFdPuhXgHxv4oJdQZbGOvTFY
q+HgxCAo8lWM4tX8L+Yq68/07QsULGjjBwaZWA9dIhjSpiyLVRwjeuAYf/rZIem2DXC26KCKdgom
VBXGgJs5sGLMqMHKocWDNDICeVjmsv/mI/7HwFm0RLNphwZimKkEuvt6FWs1e2Gd8bOXxQDkZkiF
xsBlPYEM7yrwvBlIzuK07qqlmXj23KQP0LCkJ/JVMobOu8aYIJW7wexUvotbVcJrEumYhXNpCMhT
wMW3RnfoZi/ce3tcXUmgaFTKHC2gx5pj2Y8omKM84c2qVvqaP/dpr3v0VSAUQaXjgl9Kx1nIMSV+
RvcZ45dgnBqQqDzoeH2rt2ehjrt/PjSsPFDHQk5gIozlk8JWHLKrhiCD367nyKst/2yrtt2Zeafg
EC+hD3jX67nhgdj0Q/v8uZrWTuT9ltWs2+bvVh8xjb3Q3pGjbya4vMYdx+nFx28aPlhKWgJuzqyn
QzRPCGqNYVbzX/Gqrie1ejgQ4ag8I4X+ISRwBFC7yBVPCCVQzbMjv3pE4VQzilsyw7Ll0chXfviA
UlcNojWNU8tecq7KA98HWCEcvM94+FxdLHif0pyRfWhoE/c2sugo3vkxGhjwItEEUcCOiC37XRZo
LP8s6ekvRA/5pugt8qKm5uqWb17Igz5VvSoXiNevWzqi8b/SmWuAMdPZbhBRJGq8/aCdsg9Pyndf
N14OfMIPcMyUsaPHAdH+DFS+Z6rE4/Q+qiMPZlMj8gU+ag3oj1aFzzqJix+wYzz24nlewDhvVn+t
MCWVqE7mJmurySlK7GlhnFWhB6bNNplgF2B0/SfidAcS8IrrLfdMkzwTBd2Ge9Px5kBfDin+rR0v
dHLcAL6qpMhTZy+UYFptz2hboXy9dTPLSRu9NgcAB/guhwPzq5k+1lzcsmmPOxuNJRBdj3pzmmsA
41LShi+HNOF/w+AT2m1aVvMdiTyzSaVwkOdNu3KZgmh1ChLW2ipYbiWUKz3mQpo2YqG3RJrqBqfN
4cIEc9OiZIfibClDXa+BizMO4vQtzSohmsxMgISEvqiGYxSpFoTMR1W7PGV4WgwYZjv9f6jLPBzn
1DIpwfHMqPY+9PZiVDe6Mgipdm269iaYevVQqM9PPquhyv+VSdiXX5mpVZIQOfQrNjJZ7PalAU40
gR2plqARtxIAFLKsvNEJJSEl3Zh/rAC6Fv/Hk5Lb+3zcM82muCNqEqZ97gEgrgolN8yZ1U6jBcOl
4dgkFyrMWOIXXZwVC4sOMXuoAf4Nl6BuxaqEGkYpo/PubpDmje8O4t0fR0H+bIJXRMRWZgPcRMlD
dEOfS7viq3QXRlZ14ViXI6ery5bxVw91pE8j7vHNCRpycv2oH/wOJ14wjkjtp+AgRl2fO6h70PpO
PkOcfa5Px/7oDBGy3kKQpqJ1j1wFCzyWUtajMKmgWst9w729nGsa+ETpDXKYQhfVwFWvHaiuBTvr
9A498uSfOTgZJBVO90xMLlQ5e9YVxPQA1e4llxABOgg0sO1Cmc3j/p0/9PpSMxEIOMOYCvSNmZbT
cgRioS/0UaraPY5ahzaKQTTNGkXvuuKdULNXW6iSPOzq9FqwXc5VZRF/J1Q+/ftDEghHyC5wlv8F
YezIjk05W11oqFE6lm2Gb+Py5Ue5zaUYL9UXhtZkT1OR5spk0FvJf0jbUCex191gwNT/jN8XbRTv
KwoKUObM7E7KJLEeYx8S1IVhJbx6AtWWVXVtZT8DrpVnlLYlW/e+2YYdoLMENflJDBhaUts701IT
ZwhsZGSjBjv5kmfb7PVRIAXWBl7oZQ5jvxs5Ybv9iKrBJeXk3miKo/sG3h6U0FXtMTLk/imGvQk1
ynmxsu/IKgZrqoJIZmS9nDuBJBVtjLaQO5yyF0zBQ8VHclkOVayUsCUMYo7CRG23rwzuzCaVpbrf
f18+KR+J2ulrfuENIzWmhVas4o0iWn3Q534azBl3XErEb6FFtaQhstmU2PqDMSkjPbw2cSCUJBk0
IYv/312yOX0qAIxxdmnFuCLFREu+G6awAjezVfc+wh+RqGBowJV3VQSFRcn45Kzwk2/9Wn4688zR
JqFr1Pnt1UehuV1tPjtHGiSJl55cjKLtuFbwhvi1R8y57C5CoCF/Y8x8THezBG763nk8ykQYboSc
Vuw0H2g8nztMX2zzoZyzFYfr0KabiFvq8f3VcpxaVPetoUfS8K/QbD05qCsS2OprP62wyIMabaI7
Y6UzZvR+NPr9vvqDneaivPL4VJhvtdnDC+Xs7bsX8MCijHAHwoeljfU36bgT8iowvd1c5YYm8o1f
/U9Q/pnbZ8ZWXXjyg0GPhYgxg/iIXpUric7AN1+6VhId83ZYZ5Mv5K5J+xrrxqySWVSgAhhP3KDp
dP3dHUsy6in6GDtfSC6zGSa/YwaNYCxEUtAHJmAzhMFn0CuRG/euh9066WzFX0+7eAwSUIt1yvxz
0KM/3OonQ33brVh4pGf7sEG3v3DZS+c+KRyRNWo/yWLwNBQJC/MNI41AFJZmUfDKcwBUxQzUZFmJ
WFuxU8UipwiADBTBMdrJqs54AmZfy5hwHp+4w9ZXx5CUQd7slmQkbnCxUT2CVbIZYCI4m2ABRZll
p4PLsv6fZx9+RdIUR9ZfkvmIS2DnUzljgJeGfvn1mNgroqq4OvAJwgMzmIAIlRls/vtS+RpkcGJD
PjWfPbZtns99d/aHdf+/BKAQE9DUWv25ozZBMZPtrYIPPUlUTYkmlmWIe7rREp1ieLc64jsjDywI
OxCeONx+B5ZEt+ovNhmwVgZly1Kg8QQSvCaI2r6JezBb8gKUhDW3JDphackW/dTC+qKiJk64mt3p
OuiNZZLsFY98j5N+awUR3VMp2KKxdNSUN1evL8rwNFAiXCxHmSW4hWx5TVuyasXE2FcOskH/d0+k
qJYXrD1Fyeocj83SMZLNnUEKF6OuEh3LUFji0oCmxxvPHzWDHgoBNqSf33J5+Pbt0peTyZ7TvmTh
1ulMF1PwDbIFcbPMe5cGJwr2MF8jfqepqS4SbeTXTyFcgX6tsifOxBUcWcbdmEi8EIZbI6kWfRU4
0OPTkprPhISg6vftIHLa5drRkLAbdvqNw05PfpivXnHdgLh9pZH/ghrHpzb4ysj9RDff+hnID0Bk
DP7tUMVm2GViTERtIBbiMybW3kt3XtN25MqDGMoZhbGpexxPvh1VB3kovidWTWCqvBN4mufdJ18v
/9NNntTrDS0nSEJ6Rj3CldgF/fMNCziujb2nxHk57mYHUdOm9OeZjrFFERkKZfiIHZzYg0nbUgcB
GZyfb2ajJc968i1/xFJ9IaHz1U44KE102ouQvwsI85D8l52AB5vpjVAPhAPTXA7HYllkyAjlnItn
TlJT1o3mCPI7AsswWZ226eZfJ3IvY9neM12aNaLsFSzwG3hnQp64X/Yl0ho9sq+DT9hPaL1M3eyr
HkMVEKE12GuP7ottfQZhsPtvaPdmfp5uns3QRZHRMHqE7S4PFIzbVcrGtoAT7xk7uXf1YlANUXZr
q5XhutO2rwxahXHNzgKQlIfAXRggDJ0tuF3Sk1IzcI046Jenhs6OxrD6fLo3Fb6+NGj++rz/2bPL
dyK3jsiIqrKx4k6uU8JSJ1y2kCZGe22gnyAigKAYrOZwpwGg9hUJVZLzbx9Xfw85Yes2cWlEqnGL
MiQeuLGITOQ1I5tBgswuJC0v3RWAKcUhSRnYXkIRHEdwBKLxOk/Qy7jLaTcS5Y0wpAvKG1/by9CU
FAfDEphPl0ovQ0MSV9Jg7UW9O1p7khJoRJ3fRsEUs+x2GyDLUxIHvKfww3enlKVQj/Yg1/JZzVvE
5fIo8bR7iKBAQp1FiJPtfz1oDv24kIl9ghRBc7VXhG9fEF0yD7yJ87WbfRdH2Ca5ZeUdK6pRD/wD
DiGNnwGcWl5o6a6c7i5GkrOy05QcFfS5TQTupW0xlHyYIHXDzZxYNm0a3Beo8WsaaWh5/U8Su5eO
3elZdknKMDCKA3dUVPti6qHm+i84U1h7ihQM4AanX49V+t0sbmhrQwpN3I7fzX0Z+Ke7uPVwdBP4
xz9WWtq7AzrjAJmMqGeW8mLVzKAcGSNJQouPR6YVZblnUDMXflvMlpNu70rmXIXjoW42hSgmqGAC
WHOq7nmTB/3nsS6O9UlecwTmrBAE1JfWvIW7aTy1wJVQvyh5Z09ChqfcQmU6Qy2xVOsWDvIFcqGz
ZQpm0aF+YTGOZTV6qQFJ4sWlOfYsBlClbnVK4wwXBc/AUB8LEcBtF34rsHUjyi3GxhQqiWPrTOi/
rzRDNiso72lVHHRa7PUp8i/3fj9UUZXy1IpBJN7Iuwflrroewe75eWxlrTqIsrOS+tQSHVly9W5Z
W52X5DZYV942Fr31sHbSmgulF8VWHgFsD81yKRPh7yt2oHawI3cjK/UfaZ4Gd9U3iX5OzpK2ICuI
nYqnVX6vqRD8VygK+4V4AJH9AG2kG74nZjORtM2qY8OaWhP4sy6KoLd6luLaD3NUzqomrjj5nenx
WISW3/7Q7YE2g/1MJco7cF8dOOxnlsW8sdRltqznMSnOM2EZpxmQqew/bKId8n8fFQYs40lPPBxG
qs3hBEIlBYsyjws6wjAYE+Muarzl3fYGNFjysOEXg4z0IUapp1CRbR4DuH2QnzYO/6+Bea8nIslu
1hn2Q3HR0unksUMSo/3ubNupmF55ee3Bk2JArDdIdYUXZrs7TpqJ65NiPhxm6Z0Tke1m5kAdUSNt
L8YgKHDsYIfWGzLX1pq1gVaJ+yRgGGXkIGmUzH115fx76wz5ex0W+XUQRaC7iM2138/gGDu9WkZO
ar2/l+iklozqDDome/LasMqUxC+mKB+Yk9SXQQCS3v3kPGvKIToIyJKcitEZ+oZe7VyZ8x6k2/n/
ISmkNAspJUMJ2NXF5rJQyk67qyAW8InOBnp6EjWgx2AD574DktWr4DgUtbGlsdKV+rL9akVCKs73
1jJmjtFdAqzng0yTwlifl5Zaw7NIjXsQcoepikd3b0FwGb4iKogZzFS2Z8fk2aG6EWcAWezNVStl
K/A0lyOY1s/1qzmoSF9R2UC9iLgVyidIVelHLyjdhMCt957J4Hhtb5z7uJjSHfkdCzTS37KYyusH
cBO0LVB8G/9HB5iB99gyAGBfuKe5X0v2Kux8OnJxvd1cizBCpDBLsIun7YiUW1n+d3CCVOrkX550
74ZPi3Pzx8dOub2T67WbG0YTGGJ+yIFXgnfQ+4M6D/m9v3GlkrpChdSZX4AZzrb1vYKTXOJV7DTP
JeKEfQHQuD4u0kCnF6iyTfBUqGEd0unEeo1BIDPcPRFfN52i9LfWfgWZ+klc+3pShrm2IKx31fLl
NqXThtsfmtrfOzrlanSnMdtv3QkDTYqeij7qXMtPu7XSTXQQY2Lc76+AqTHhYe1yI1biilqrxq1q
JsxSK1eGv2AOMQMj1NexR7iujNGp/Tz2+xVwNl7Kpx4zj9yvhIUQC4+3fFjM5u0fU/Of2UHQa6iw
T/eLaBO+6x2lZsnZFnb/0Cbx55w1K4aakfyouPVHdI4RZIWXzG5rpMfIu75qzIYUTdzW4g01GKhV
B+/Id+LBqXxCycH0GRl6NsYttX+3KhND9yJYqX8EMl+NYApxto2CnjocnndUsg9EEFVShk1vGvZ9
o4frHm43dirRpbAFFXv/V+yEcBOOOp8vwyvvlSUTiHoyleiXm9GqMsWtyoY/mggUSjPagH2weF3Z
WWlsyXJn7RTwkiVZPVJkNZnw3aRFqc7TMx6EJeL5Y/eQsmyaiZ4C1YWFxlYoVXEGT52wsIC/kM0e
Z1KrZN64Wc6M3txL9Bh6Oqs2hzo+oP5GAPeZb+WxGi/5KkUx81hbpYC1GCrMSYbDzs6+PWI+ztEP
utlecB5RqfmHpKbcuGffuvdpEZglyr08IIbWXE8nTExwSCCqLrIAS5F/gKve0VCIUwOp1x+df1b7
t30Vwz7AAvZf2oOZolQF2U9b0cHkSgvpGhI8cJYmWX/WMA4NiDNQE/I2+Xn3LN/vb4S5+JNN6WpA
Nw0JvoalewJxR9vybf1KrU8Bh7mXlHXv7WVufXY1ALtbvBGJCXMOWCOVMlV8yV7BsxBs/sHE/5T0
834u2zIqQG974Anp7/C9YR7eVHYeJz4AWdc0A40rmAEpn0XdE1sm3LkBl3sA9Wws1QgYSkdVhgLO
fXcsZs2jnnK3gGXJ/00Jdg9E7P9YmivmxT5moywqakdza+av6Mh6OWhvsLL2Kv6fRxwvKMM8vagS
0GXDAOJiAX0ry6A64KKcDv5NYnAaaW50RmQfMXjnFxRkpbl59YHqWtTCJSaFCt9F4/sO2KPBDt3q
7FB1oEuM/L9N8HknHse32XWDOwQ9wOZBBSTjCLA115ulWQhGQPwVoukd045uL8OgVKqOdgq4uFv1
j6Xw5F/WwIj1MtfYi6oyuMkIWcI7dS7lBn8ziGQJnC+0oFx7yTvGTse68djEg2FyNH4SjXWv4s7Q
Zd7eIpo6swffPnaBzrOOJVkfCbkqRdhpkbsyKtfplmeNGivUejmTHdLTvF6Q2/4Fjik+n48wdAhx
D2PxVpdIhtnA5pPY8nwuz3XCTg2QHuhWHgjVWMB0nC5NH2BAgjLcJ5ec6+1Vv88qhiq2uKt9M7mG
bJOv+gwwQQdZ2Vy3gsYWwlMvlsiCoBkW85YNSooQuYDzS/ADyW/Nor2ZKiimIvOTJd1yToomNo3p
eGsMP//JiTLkpgprw+qdkSBZO4i8GN80D2PDqyqsklGbSR48kIQB+liVUXzU5mjSPQ1S/CBypltu
Wv58x3PBxh05IDtT/kJd4aZzoZzZcVsBgUS3js/Jp9qkrwD+fa8mN2/bmQQhLvo/FfI6wKzwZH6Z
Xj3w09SJusPi1x8zNMlogNBDDTzEjWBflCRyvNVODIHoPkG2x7JDCXt/0m9jCMRPBO/PEaf6lAm/
hmvMjGDw6AJaznAWVX6/jlZlSgw8nM8tnJql2oYJCGioGq9yfLAyZ0LVof/uxf5GJndQmsO73MUp
pdRi3FnMSzi62Q/6bDZAMX7ybnLVBaU/3twU+PT1SZ3YBg83nt0E/FtGmzRE/F91sHI4dcBkGLMt
idbQvLc+xp+dcIfTqu+ThAvd4xJ5gZh4ywwcL/Yq2MGbT+qtosIfdRNYPZ/MKhOiRs0sM7bqxqC4
9GAwzwe9EcGdsaO0OpqFWOnubdKE8/FFrRvts6O28rNqsMMV34mUcNmOACwmxAHRchH4us5m68tP
sOeGkHG3pMLgwy4JyL6TN3vJtHzX6X8fl3Q+DwOXmuSu5zlpUCknPolqutY8VapEeVJarf/0EMch
awJvJ8ffV5saFtaBBA+Jj6Qcy06mF+gyoYmZm+x17/trJ7b26R5QZFGI5UPGl+aq9+fSh1Y+kcv0
tx4ZBgKte1W/puveNrSXfsfWVsdIClidyo+YONQSYisBgHxYxCe8ETGgyE0norADIUBW/majAKfG
tuttqFH5DbbpV5uYEK4HQfWNgE1M3e/IuP72o8MZuPDMMKP4iRYzSLGZMKDPDWCKproe7lr6nJsl
Y2yx3bb/NKkJhdRU0UYZkUApKuP5sicnRIt3/SYUwy+wl+9n+ZLr9AqFORaW3oarIZv5zq+SMkgV
TrUUdAK8qPIztkzjA1FV+7b+wGQQLK/TPg5e0USHGs/4WkTMZ1dhgqpl0Nq2qAG5rpH2e1N5utzn
irnSS49EUlbmjBlg1trCx88sAzXt8uwN8WB5xaIgIyZJ16f2qQtwmsw49zeBPMHPcqEVjWO7aH9j
yLCS+hqQ60FlquRJhug+B2bApus/cuyadut1BnTP7wl2UvVxhadR9h2u1XIoSB/kh2S2A6k+Bv6v
a841KKe9O/YwQ/yu8qc0+BNfz8eHK+kyyQiexDMJh6nVvB0VdkipdYZRKLONUFM+QhTDDdAcyDju
lcJCdvZSpQR/HCoe4N2csS9Q1EhopxT5j/CmtAZQhVh4o3fBC4ETFqlqAPrlXAuoQJ5RCHwykfms
fgEpS5CIKQHt0Lb1U3NTJWc6DwDTVwk0j0DPM1mDmgMHVR3r5yQe6DnYdQ8ZTJYt/L+XraJtPr6n
7eHGtDH5yMiUCBTS5M3B2v9n47wF8h+lMw3BATmKTqVB16pGZey0ZNHtBO0n5Ad1jU4B7slWU2fh
3YCNjyTEY2OPYzU8ICoW5I3Upx3YBMc4JlAxFz9RXNORc064clIBBFssarBkAZ1teoq7xkvncFs0
rtxClSFBWCsM9GU/1jvxjXMXlbOf8RhLrItk0tXjnJG7Et4ZKktVesiXZ+VKyu78aPjnd8yhBXTZ
JQLa+LkAu0e2W5MscW+rNkNf7pu2mmGoYIGNe5CEuWFVStAQA6KwCC45eaiDUKrA9a4py7VCdsHE
LBZDEYle4bnUYumqzSFtwvyhAuEDiXDyUlPqZ4TFVox6BjGkr2DgmkMUpXZCsldfGiBkJTT+dQJ3
Y6E59ZypXylldj24lgVi/5mk4jCxn+9cdMO6my3gKVAhOX41OPpnF5oe5EwEkIwa+vB7BhHkN+Be
dlFMGvF7YBhVC6fPabqTLKdseyr+O+Wn5Q6FF7BbMVos4wpp3CyqQdVHVq+yc8LC6IBmjZZIQ5a5
91ygwOAooODVMkCCf3lJCVbIoPWdUX8CD0+Q76r3pFEuJoLjqsZh0QCdgckHWb4B6GUfGPZvN0is
J6z9GByl1n0oC/+aSGqU1R3FvX2IXSo6MrO0S49lDwLWOhYGXDRxV34MGPAoBE+C0/bi3hgykVaR
xbfR7kbhsqufHt6xlhiNpBFAtsf9ESFbRBlCtex68rUPh38cQeXJVfxHHWfVN7RV8yI4WSk9+/Qc
O3nVXbdcDEBEu903WIgPMio/BCSxthNkuvBVCrpu2wJdThm7I/abcqhJXfEZUO1QoE3PxfQi/jwV
jQQ2v5/QrNSkp2XXqMUAcynDAXvL2W51+Yj38lrXvSG+EpkrhpghYZwaveWNcPeYLlStInZL6g+3
BhT+O0CzrctMquCZtKNZoEDsqu2xB7vzUqiazBSOx3tQEWuUg2z5JH1V2E1puvgrMcRYY7jUBW4M
NULi38WsYONbo6SMT8gH81ahzyl65NA3wLcNGzcnF9aZtA6wMUJGeliUAho613t/2gYvWnab/idT
aI1tCTudC5xSqBoXew+5BPJRzyT9qn+KkDlq4VQnkqi3F8Tlupe8db67YchWI9IjplZJn3zT+XQg
jJsZ+quAeXeG92DVXh0lU4YDd6oe9l2Wu3VE2ywsyUzuA6+IW+DB0wLLDsHhg8AzYVCdZWyEkJRh
G+fngqS3Q7crSj3qbPSaZJNam+j4fSKxTjIr1OBBl4whycPgSzC5NG1pGu3Rwb4I3Oc2OoySlrdr
lRRjPoiBhVSlLO27zM6UOpIJNTS1ZQCc6woZZuY6XFdX8/6Ux9WTtlDOuvzFF+9TatVgE/YL7UtP
EcSKMmRuXOBuBi7t3kednhhOot5hgfpEkC9BOiy4YdMvf5bksApou8thi2fw+E27gUhr3bX/6ocd
pIb6u0OCidS8R9nXxOI+/UwpI/QIhsH/8Qp/UznSj+YIHMWqHoYSafbnbke2YUso5MZPwdRzAdg8
qIJJFst14Ir6yb0EONAFB3rlZzB2dH3hwTyPw5zwswNwGTnwvCQyZRE47F/lXqcoLDBEUcBIxrj2
EidDJlYYq0Whw9wXMqM98/Cn4fh5Ce4cbUpXBdjxPzY0XFkjk5SFIcZw0qCZUulOJ0VtmspETwkb
/dlp9QJBd3M+b/zDTftXQtBj77R2B0RVDDeuElQKpatlCmgD7ZAr9ycELcpFLxbXb3miRUyOs+jC
Lgt7vRMsb38EnlviiUwJuyEQ8GMnHQrYLLB8quiarWkdmCYi/bifFPKjf9yCU60Xyjn/CkX8hA2o
GSSgX0jToryeJma25vxBHZ2tTuXHIDfwTX8VmZM2Ym5vAdZMMSKPkXcOioCL/JkQdAJe167fm8+S
tzbHwiVRF7a3RfFIUzuaxVlLqwYdmfzVqptf4sOd8l02/8NGWwuPRWDB8nQSievClj8nBFhWrFDP
mLJZXJkol8mPAhgbfumzlY1q35hbAHvsul2SQ6ZtfssQlILOvk1s8CUVBSnS1cR9ETFIfpb2sTKJ
pubKXq5lBsptKNGlPqTIpLuR1bHH/s4gPkcE1mL1FD0Ea4YYEprQ2Jw5CElRP7EMgRtE0fBhg2hp
FQChjJcgfgiq8HLCq2XqedELsD51H+Ux5W2cj92jtFzHLA1icH7a5ZsFLdDut7xYSet1dpYVCec0
6IH1ZcVPlj71p8GQQcjCfFej1H+ejq+P65MsjiB4fEAeA+auqnyF/a1yhuiQjR6g2+hgsVfs1jgf
2SOYvProflrjbPmrpPE5Bra6BV6M/rZify6LwOWvhbD2tGcpx3TGs8CgL6M9quJ8GI5v8Rua5ILz
VeyL1Fpvni2M+AHifmQ9AgnIZgpWhReiJF+0knvSSp9O3hx2i0AX5rh2mJnSGIqVYoOQVzLnfSPX
wfUf1nvbSfTRb9D/giLjZu2DO+aTMG9nmnkNIX41NBpU4vyqFH8uW8EolArOnalG7ZCrizRmmpJX
Xq8qNCQlwDvJGseLPcc+orqlR8LSD7t1VCMJPwB9S4uxG1A2aXQpFqAb2TAPJUJzLD2j9rdgH9hg
YkZbRqKC1IIsXkNVbwE3Uf6lRmidCf4HyPDJpPtpzvulhX+O+SfY+lpvVzQdXKDl5fnHvG5M4ouQ
dW5cC1S5Dy8vvVH9/GO2mRhAMHZnUJ7eHQw55Ss25T2xcimp4u+C3AOeVZqz+vSudPcL/3Y8W7CO
GzvogYkojChFT/xf48NfT3wMUneH0fY0I2YkIcT8zcjUoVyZLfuZrZiA8la3nE7LQVCXSRRo20rw
OZ3la7uXa9AdlJDd2t8/bEMQWVi/zZb6EcAz81xWmKfDXrG21DnPKGlUWTP75MzHQFFfsFr3KxFm
rIoT2oBAsi8i4abAcnfWwrUCA8DqK/JJA0sU/+SqBbAgDcaHeJRtpV4LUReLp+CoA7fQfYULKEDp
B+hllyohDlrrsKeaX4bfpfb8BDErcmj36F5rktlDZXy13sUivFNrrE02ZGE5ZiwjOom/L7PUrA9B
60jWC4wXC5s0BsT2WNjKF1svdCp+ajmpXPL4s27PxHEPIYBveOZs04PWwGWAWqZYijCmM023Yx11
lAUH1c1iqG3JfA2tpua4DZRmKSB190+zrZp/IkbuAnZnfUuMqydSooA2wG27gjWWU9tXsFsxlr9S
RBJUYK+d7TxViC+74uE7npGNdi8tjKFMVp8NDQHQty9wG+moZyFmcYypR/x7VxkzOj8l+E9gr9nC
qRY64R/sCRnm8b6q8BoCFd813rnMtQ6tb4MPvb1zUmFfeSRsYP98WuDVtl1c/MvSflljOjJcDDzS
QEk0+FxNMb393LstWzeSi/tnhZACy80FjNUEFccTPspocpiXzEjMOBmJksSE91R9ivPfi41BTQLm
cGQPCd6bbViG0iG6t99Jw8HA2BKj/YUOlGD/wuW8oZCs3Yir64NS0UaQPKFn9JgBBSrMaDulAvp3
A5D3GTUm/rP9DxtN+s8PAHa3eMBZJEehsnBF+eCEUJWigZI5jj59ZvpaK0cetcRc87rBKLBf3LoB
LAX9WnpuC/20xYJM/PKnA5xKTogQstJJQebtNkwKmbjFCaUs9dxxeDN9Sm5cxbP/JsvVKzwxYajx
Cg49w9Jz/d60oOaYxth9LXm5WDf82Qmh8ClnkWBTnL7PyzbKNkuArLi8f3TjkllDPl9dM29ZFU6W
w2p90tLvN12srbLb/T++CIon89srqHNuzTcA2wR4WydV9hsPB1US1R5CCKTmax3B3GKhcsVUwc08
qIys8Gl/n51OkmXaQsaIYwMs0JlW+H7Nov18Is/JEW/f1O/PxiRYLCIb64v9/ckj3s0HOU09QPmO
fIlX4G9lpQEfFfhfmeUASNv5xuBbzETgdHWePjtvaY2lPGrU+whDsDZweglNq/TOVySl9yyFxKlp
mT3PwUE8uJLgSJmRcxp5gcichoEGjIJhpRIN9Y8+3inrUILj/uV/kZmC+wfKPK0f80y+7PJHgDmK
NS6CVx9SNPb9FRG8jg1Rdnr4c9IKD+97flDIwZrClKwzFpsdoSN+GNsUECakQSRDPkibbNDZhoDD
d8nIowypGc89kDaeIC9OsF/2MZb7UxUtwrcT8jXJuIu9BaUIpz2wab/AjTi4sQnaazi5lNUUtabT
5A3ZoftHs1fIe0W4EuGYw/pDKHjG3DOB9HoPlXyz7wU+faJ7VeRp1A+9X7+SGrEHOV7KaFvxWfuq
qNG+xMD2/zpp81a/fwX2a6qVwIw+34VnldmnGevbfCTQ8lOSTv7TyU2vrC0fqc6jt/zb3gPfRPsq
XoTsUHxiA81cG/5TXswExkqABeIIJKAMuQ+tug64pl0z99jdTFf4FR8GCd5qQIgwyqix+wNxVof1
AVGd/L4udDWLutSQ1xKiK3EsgZTULfHL7GCovgerFimi87WQajQPs3VbW3E6CXybz+6CuknaqBVJ
Y3UF2dzGwwnImczIJjynD+/gQs7F+YkqQMt7z1WUIR2Q7LftjvoJXJwG1sc5YDakfDskZwN5TjpU
kiUcJMsO2B47m3F9nrCscNHUxnVapt9cs9+dC8TwpNPKz/RP1Mmf3CZVC7EuscAnVPzUG8KjiRrf
HUtErqoxSUxCdlOkOjcOqIk7H6+SgHn1wk2hCxoDo4xvVPOcgXqcMMUsxHWmoVu07i7C+u7Z6zzX
VpJIz+GhDUCbTU0CN2CY88oJkLVrQ/xL0WFkInCFdAHJbl1Xz0NxfDKEHPSaLlktbcuR1ibyERhZ
EGmMmEYPdRYXQ/zSx/PcVpVEiKV2GJKkbdDpSf4GBcM0hNxT3bYZJwQcZIWns0IGEkbTLvzbh6l0
4lidPIKPrf2MDScHGTX2nh0PYYYib+Dfe3rJuWKfQdFNJOy6jN4qYiBIb4rPZnH0H+jgVGTRy4HJ
IETdHJsPPdPbxDYOr8O7W197axHnVPr2jYFirPq/dyftVBuLFaLKdhxGkaEvr9o8eurCq9mDPyeU
rl4NgceKBZo1z1RCoROUxX2PqUCVuAWNxk4elwHJkwocMyVe+ArMNSvd832Qa0xqqsCseSnVixSW
pUiWgrLnRUWm7Vaf0i6GqoamsOZMaiRJfLJAEmi46ANDEa73P+/NGgwQGxvBwZ1RjQLRWk/LEZVs
U0yBGGTRARyT8BiNfrEbAVu4UfiZI43HczoAXSmSIyzL72ZW9eh6Gr6c8r8VgD8XKltb39S++4rl
ZQqC2VJk/eV4SQTNYmNQVHGRAFNLzn8+Meaml1bISXKFZk1SoAAnT5oBPaOk9MHw0LsLRQIFHsDe
ZzbX2ujwK7epWKkcK+YDcN5WP/39DfmjFJuTH4/4GPswiiBNjY5WXraKtUuTwFdpyqldtf/X48Hn
IUpNWAWmzcbBsjxHJ4wZS+jqsbi3h7ExXFsQV2fJs8SDQVVg3/WU6fV+yMKFx6hE7xp9KwKEOEbO
SyZ0k/XN+suyjoqcGu5hlxavwFO5aFXB++v9+2muU8R0uzytv/KfJNaHZ+sJDrp4ZKgYxn8MfHjU
xN9BZqGRYZpRBO782jCZB4HOFBYTkusTECaA6tM9vG1F1D4gev9nZWJxhSHlZgY4pqHTK3g5/TxL
nkVnPrp8Mc4y8bX+GwFvjmVca9RmPyih4FE+SIiW9Rm+SJ5q0GhrqSgSM2AVBE37fXlVoFFtDjfs
Yh2etU9d5M9j2qgL/YwtWzpER8zvwMi2YLaDTF+DxKvrxSZvVet+0QNOwpbGm70qady9gdbZ0BDd
LPUBrfV5/lHcB01o/MDdfkL2WuMOiPlFjrVfBvz1MyvoRDIizS3qzGPNdyxotWDjpGt2gEwP1EG1
HeFyCC7p5FKB4UMzDifzbCgdeVWoNb5i+hSygippdNNeynvXqeDEzKE0x+Ab7OzULX5XvGsv9KFS
PjhrTsSTtFRbChC6kA0ujM6lfkpwG9yXyVDCvzH09pljKY+T9jTV2Gb9VjeEFs5bZ0HFahyE0239
MPWK/VK3r3Q0nLLSZNTOETdtB5DDRTnP1HxMGSMduF1LJNV5SsPHLxWawjk9f+RHYBQ48Bqh338d
D/5Athkc+DTB7rQ+J0BImJtB+/QBDeIZ98OhtwlIqXGd5uBHTFhCDbN7mLj6XFaabSmtgXSHCI0Z
dZi0WpMjJtZl4m7xBMDYAAFaLtnbl2smuRshHcXj0KG2Txv941b+uYCKlhNZFrPkuAJ0WLlo66uM
MGVJbX9EjSgre/jNEzuDn6rVy16qSqTJ1N0rc8ZIfnRu6k1iTeQANfIt6jgwUv79EeJfjogRM+3E
ZLcyMd3jV+0f1pHE7+3dN/7WKEXa0hK1ruHt10UnkY4/iVjOEIqDrOC1G+DtERaYF/ZGxi2Tejzu
GIm7LeMmGWp/d/ShkiGpPOBtOcRF6qjPpscKvGfbdg1G7QPNIh3gcH+Zv54Vkimt9n59D4r1V8TQ
N5nhKrY2urL3+GFnCwPs8SjEPjU9fc5U+Z5d4GjrcbrlvvEqHh2gkMZEDhthBP2cIcFHcrzIaKQr
lGvN+YoeFC5Sm4NHOvpuJdzU2Z9LAPBfYY5u1RaXI7XHWQzhLY2z6PO0VqbnJxlv3Rz4ke8Hbg4Z
18fwqt3Zjq++1IKsE1T+qqcjaiaNjcKBhhtAqXx4fOAJadY74XP9kq10aP8rZSNkTw3VcNiO6ZRB
EJIfRo/qTKPBhCf0ZsXxSiyYrwIck+JovNry4wo6KczkVRAn7vxc3ZRvd5CGFe0JiZ5NiPdfsaYB
N6+llKj1C/l81/AbNuSG7jfx0P7PHx3fZSO50O/df6gIrwJ0JMjJM+Lr1H186EaAoGIp+KlUY1YP
KxiyqZssDPTNkgtehWC51pGBPC8iAPE3uey9QZkyQjwr3e96pu3+0BIUczk+fbU4V0VDA5VGut1r
pWOXDk32bbVkvj4ABjzLzJFHtiBRVxnsIM4gxtwR8RcOt0t4wmXhLIqGJEA0OJXiTkFUJqD0KkKC
KusmE+wVLiteUgia3+ZMwCx4qpzMwgX2E9QKo3wTHxnAlNhNw0O0vwJTC0C/be7ZYtHFijIpPZP1
FsJ17SUSA8+0HniAk4k2QbrmRiQLJPiZlHl7q3y+jLkF6yRaWtihhT3MFvvAYkeL1c5tTq42Gz1r
PReSDC73SkSj+rEUmmFU5b5zb4oNB17yZW2AyVamMHrc0u98+Uqm74o/IhXl/64M+1c9hBOf7dAX
8aTD3gr0y/h8JcDtiqoiQDBXLP7l3m1deHN5/NQ6bF5utWVJbYTljeVZmzPNIqARi34MBlZfUxOD
35yTYSQBioR7sBq+KFuoUfqfrVAE6gS6U7LJ5VxrCzuCZvtxLkjKYvhIMYNMCkHbncNNv4DjRbcU
jbB3LRk/UfawhV4OPe+Afl7CWi4rSKxlH+wcEpwkMNe1QRqTNlEkfyRtTFtRl0L8BeCeknF1PuIy
qx1mZvcMrmXI+fbGRROJ/9rPitmMS0o2IBDfo67/UXHcMBRVcFfPif1JmcY4UwENsWvcAYxF/M1L
uNDAmzPt3G4YsS8m3Cry7kK5/XG3UyswqXs7k14SLBbrcJwkz0lsLk9pobyzFAQJsbHEAF9LAYXw
zD3an0lzAHs2cFS20/lsotffajCxOQSpDKsoevDTF0/vztAiaN50BhSiVBaZ0noaOg92FcNpPkYf
78ABnPBE1EsRK1675ogRQJ/tOi6EiVgztZuQieFIzKjk8F5tNp4V730vt7i4hP04yiBM8l0U5RWI
GiLcGG0VP0rFRvklpf3zypTw3XyRfx0VQP+WqXIwTLznGX8MIgdIykuZocHoNFqfrXJnpOBdGOX8
RO5OwcQ6VfsDOh5g1Tuq4b0fHCT4tV3Ub6tjSUmFNax+7zwrr4lf5ik+vefqU2A8Blv4wMTPObgt
EnguPhc1dBFBUVjxKYK3qlce1y1KmMyOCltz9niZ9msLgbii56NYvucFnJp5G974tBTzYd3WG4oR
gMT6X2n6F6SFSoaZiqlDcfElBA0uGpXlOeb5uB+sq+JLjee847ryVBxsOZvADxRsMIS/MukSi8o8
ETaNfJKcR7El8C4VvLNFX1Ki9fxjkPaA8FbIfDhj3e0aBeQIAKVrFvTXzccbcex89vq7g8sQF39K
kah4FlRsAbHZ2uPp40V/30DobYVou7xya5KHwR57hVhz8TIU8NvZBBXepBrchju68lZAAyn10Vr9
A3nls/TJ8Jk+4eZWfYyUzwDcMQ1rogoYVitjjZXQQO7ZNHiVAdZsYEkKglBIW8orLKlxXEFPprKD
U0/7CYpCyJAp9AiU2UBYyRrkut5Ri0pNnFYPHhPwymgNamBF9TT2+r4CwwniguQvevj1Q5hCP585
OBYac8FhuRs/i3q4H25GRstkXcY2LKPLAj1QPBERUd8VD37CIc3+BdHIqoEjOTwoMgDYctMMeL/a
Zo+I9gHlm5fxb/BLFgOJsTAGA2/Mze2xZd9twPcmH+YqDd0DRjjhmQW7XB+CWA1bPUUm+451F1A2
wl1oxY8Ibf8kMMNScVUrsf7yMiELFI9jDZ4vdadQ4ADqMo4jTPStnlQD0aD0cfbwH0Zc+QLIafwI
lj1wKDrU4Sszzfqyw8C0Y7LAH1C+5pF2/7jDO15ZQjEmMonx3lYU+DEcbnFYOPrOryE3ANJsjuRn
6nTavTp+e1ke4/vL5xqh51HLiuAdJD8HHYIKNTLlAMrts/o2OUrvdfpLYDa2trlioRrBZWfNcpgo
4VrKjPCKy0Q3SlJHHVjhqMAUam/3tO7Sqn84WK7F54PypFNBywIsGp1wODFG7axqayDZKp/G2Xo3
s3MwginBk4T/Q35QX6fATdhziNtemqYP6fkD69Ru69a85JLOz5kKyeqE3OpR9N1qgEUng6XQWfWe
1M/ha0NOszwfpn4SlNHrMNwLWDm7TqnoiD8T9eTs5xQhIg388T/8dqsyjYrnGCJBmxU0UyPIpW5s
LAaul3Fgo52vz0y1b3uVRU8Vl4SgyUDrhHU67IXlgLfAUSRP66g9KTgyDGpPcPDCkwde5mxI4hjK
Z7aVrlcJuYA/t+HsupxC7Pyr5foYflkN3yaRIck5w2WJkFIfBhlIK93gTOdctc5gLb3mcsLaN9RG
6ai+3KvPhvuaqIsWt7CuVwtA3JukYqzdyNBjfruEJv/++BtWkhtKH0+T5xLkucibvydzi7WV7HFo
5oLRpAFHgDW6j5c+JDYZOukatoIn3MU8VQz5ulAwNMwJjhFh6lt9qli1fHGKpxp26xF/jq040LU7
Mw7x4S13po0798iqXTWi/JYaJMDQzNGvV+Nhq/n2qzS+K6kUAWBHKkrSLrd504SLTzLw4xeZjNRB
ARCn/73RmMIbJEf8ntwqSQb+orIGMdZX0z3gyFtgHIGVkxMjoH0nbUTPXqLbGsUHPm+YBzWJuuCi
CShYZRcSx7yHsqCSaosDhWnMYsQKoQyVTjh5UAu5BNm60rRqtqEM1D/Tm6BmzeImfIJ8Bim3sJKH
kBPev2g0NJJgRGAqb2fbYYWWuO92EkZhsSF5eMstXihxLdHfQYc3xK4+U9JAuLCybfql6ffIoXGN
GARu/ZnqZgUyGIFpjso+Ic268mUetOinVtZ1dv+i63p1bh7lhKtO/7s0mOT7xdzsoTb5PNWb8JPu
UT+7WORdPOlV+jPBL2Qpoo04Hh5pmKLXxHjRAzSfP2hS/ebU1PWv9qvqe4THt/8WUq1g1Zp/Fmwd
IWNpdMj1OpYOIYdxejiTFpWH7PDsKdDlzirOhKJAPOgjSqU2fC4thul6qKqqNX4O+j028ODRdyFB
luuYg2RPOp9jdkX8+EJq0hcBPyaAoHlDg9LmeuWRj8wApDKqy5dJBO9wsSIeTgAEwiZ3RI+Rr1Yx
5fesTqa2cI7u2KrTBRC5xhbI9+X1azaTk7jOe8LoP3Zjs+ld5Xe8PsZ1QpnUXd7cpl9mm8JtxAa9
kerMrje5F5dU6XU+perokjwuicJ04Sj9ofSKYNaHQZrFSJEx+6vRIxFMDNSPAkbmiWGiz95Hhnt/
F67KqlGYOrPHsjBVAzUF07BvcjSViBZKWTJbdRiS96Ixt09/TWdVPkN4ou8oVyk+F0FMGADKE2v1
18RCgpuNBhyJ0MWH9oz1HjYtUxBjXPoonbpzeRog1dB7rYGeviuPABrh4CWfAanIXa8IuUYD2CJB
eImaKzwIdvESQzdmpVJOhwg7NZ1swWe/bGv//8kHAduB8C3e3Lo784U4IVUqrsEeCuqhQmzKoDVw
c3MnqvMFl/S9ZKmR1ykA7Nz9/6fw4zV0BOLof7IrdyTHDFURfJ1adZ89zDRJmkbcx+WS0C6rvVSo
1qK/YGcusdx3FIjEPfwmFXBz3FAJlnJZ+MbLXZHU8b9OAmixyijvqv4NtRfuiq2crwSBRLxbheqY
kcXCG+1Oyb3MV/39yqEGqoaSRxGFt52Rflok3OJ4HH2IoAM5/u9ZzWdbfTksSsUziCP5mMUI+UsB
YMBKx9WfzfahBeVNNRfFuDLfBOzj6XNLFZuM0pTvY6osC4wVdfJoAqf+t4Y2QBp7apm11QMXAVX1
HKsU781l4QaODBbuPaul3SVDseGwE6x1+W+n11sBmQAR3e6UPT1U1pIckIaEzMBt+d9wsRko44oJ
LIpGkLxi/Ih6bJ5izH+Ogp9wyd63sGDbPE7hyxyNoVZWTV8dzfC3EDfRl/0ix18qVWau9SLINLqS
5rCO+nRnaYLTJ6EugkVuSonOk52oI7f3Un/hSje32R903p8vgQlT97Opfe35ToWQUj8+Nbl8bMfb
6NF6nP9ITQK7f6gC/O8rn0hbDK1oHeoq+C2/EfRHhXB81UTWoZeyVDkiHRgYy3TG/ELPVAK/DjQy
hckfuCV/W3eRHOZ8Iqmc5gzykylUMvqyKR9L9YeOd5OGogLL0CfAb+i+arj/5QZgGgqiO4drya75
75bqBqSHJCy6PIlBPCREMX0aLSTCsv3o3Iz8vcPDzDBFQnOPP5YVGq77iZ3bQPWSu2/hUQZYer6j
T1xmEiltom835yU+o+Nqj0BwcilguE960LbH0hF7zaZBaNjxSSVm7dAq2ZPQSurQ9TYaOUP25mOZ
cdmtL+EZa1dYk6l96mB+LBK67jS50dEysC/lqlHEWt+wfFvp9NITf01vqHUBmkJ5VWyCTtAZiSrn
gMeoAOEvB4SNgbfrfboEXRqFsh4UobqQ67lEFlQ5E1xpzmVOnefwqfiCAAz30VzTnZyGe9OUz1OI
+Py887lJmylKCbIJ6V/cRQACKVSd376RGWoSp3E8nYfGXisYdgrAyoSBQB7mCqpgY9DSXK703V3t
TCmW5v/QcrANijLVlboX5e7qP5gKdT/h28TbWJzieL8mT4MRbx93hW8mNLYL+33/5zvWfR0LglWg
pqyNe8q0ErXI4L+taZ/03Ltz3QxTssiy+7rER6xmOSI2yU9a+S7LxV+gphqHKHM0kbghQe/3w3Re
pIVda08ZrtmijZDvo2CZJEojQ5DVXN7BVGa5S8548TMoftA9xJxz7KeF5hpfM/tssbCsOCKejewK
a+eGy7fMTzS2ZsytQwFgsrT5svNXssItImbSx0Eo9WKDJ+kZCxVsv8lCQQsVQU+KvGBqoDLLnb70
tdZoIs0STn6iKTTaTrRJUtBIJoFRPWtd8KSbMN7wF7H5F2G/oXs90DuYZpc9Zd/BNMlY6aN5vIWN
pWii6wDIHfsU8uOwXoQwpbUKlEqEvAH+ZHVsxu25KsetqMdgrM1+M6MXbMfvXTvKl1YLkEm4ty0E
PSsbKr995zxloz34GkuL37Y+o7BIHtfbJo7ePFeSOmuhP0gYXjNp4NN3ULN04AvGaGwUyTiZNecj
djnw7B1pipucdeoIyqYdLscgznfg4qSdu+itJmeMfOQJ9BZQclqnlz99KrOL2/u5Dde8SgcLpmg5
frj/VsRZgT0mBDB1AL5b9Nm6C5g40BH21fLoz84dHvp1a8H+Q4Agwows51oO9JXUjC8AfFj9TObT
rYYDWFZkOkRgEpcAVI0z8rfODWgD/LQTjZA3SbrEYdkpFcJRG803Zxzl9cKq2cxGxldF7VVACiBc
lo+5rEtPZhtvXHAgQSF1djPArbJdhc9z/dZ/cQemF5eKonU3sDHvWMkYWn4M71zWO917/PmiHM4D
cA+yDsTA1Qjh0UFDb4mla4nTTTBf2Y8koIpMBePMKvB80W2jHzuC0hGHqUol1l/1UzwEYABdPAZg
2w2wfwJbLwTc2kLWP8QNqlvsNjpHhUolIGV19j5ZPdQgk3Syw1hKcYDVgkzsZvWU6n3LHBLGTdVe
M4tdDP+1t42MvgVsEOIitv9UycMq1skwLijrQqIuH83+tj/sHxRK0xE4hcXxL2V7mttk9WTI6tr2
64nIBL+Mhs7+CtEV+k1cusIBspXhpoRflgWxrpxZWDBl6pBjwEAOLaoisq6/S/tvb0WwfYCNWVOC
QWzjUEaxi2lGANSLuOTXRQXrCoIZ+BL3TuODhX/5K/TjArb8yYgimICmXrtMRBHhhtpM8iRIEBWE
Moy6/9lTz55pO42G833VubqZ2y6okilFqZ62igLLe4HAEn0h8L5igEoGQPL57e6iQMJPFN8cSD/c
2GJFa7IRK9GqKQlMFe1418tgsNLIvkjUjYlmt5GQXPBQMxbr2fT5uAJW63WZWlJXsrb8trIcy9uV
f6R6sBEk6ejJJy9d/WbsiJ0Vv88OQYjYo6CDYsj/0tIsyIYh48GNwWLIGwQPtSaB+ADkC+g9fccQ
usiu/Mra3cX2D90FsE4JRvv9lKry9/4e40ypt7vHvCw6qqzZHtNmAQ/I/NqpMxMWQc1pleT7zX8H
3IP4vKZaEBRtRdQfnriTVS/TRLsQLNfp+TCBX6SHkV1X2jTW+Y4FRPZCEv3B2HYEZJ11caqReA9f
58hpcdUMeT6ynCWACJq9Mki/swfm3eQCiq/MMq3OaghPipl7szC0e02Y0WWBLTfdM4L7KAmZZ0SS
K6DqLzUVr7qb8OgYr6hWb5BpC0GS6dRufdwgxq7ArBx9d3ZLQlO9Roa1HR28Y1joNOGtoQ4uDaJ4
/uYQix5PbGfe8aHyeyVcNQh4k/MmvMzztd9xNpemTJ+XJ9AkFYI0c4k42ofOquaGvZwdhzHnEnnv
PlKSVT5PKcCKVVR5EgiACeY7XBsNwNVylAXDuUeZnMqRk4V5NGhXBUZu11DTJmARLFJTVjNY6bzn
jMqcJFRf3K23G0g4jDAXnM/28USJWHTwL/DfcTxknn+pBKfLkSGHFGzWUy/14r6JRQ12BaWSt8B9
ILW5TZhYaPodm6CL0YTnpuP+QuTrCx5tflpZRI1QDiTLrObVAUIvsRUxWFgpqPaoFsrxF8SbQDbA
Oo0dEAbteTTF5tHHXzwg6z7a11rhdx7hMgfPFWkx+HhXNg4hUnbZ3Cht4qiLCIoAABXXSNl9SAHL
wfIwUeGMzuErXvfnNI4fpjxLYnRJ6st6zKG5116IXcX4mfxINSOXHKRNLZ+OkJnMLKfOeDyA0UJx
HG6DcIhsOhQHvRtz8qefQQ84ofCdHYQBv2duWT7vo6RYnKPM0zT+IcI3tvPRVqGi3uBUb5me3IB7
6bMZbFcEWfwxRmUy6joIKd8H1NqhRfXAz/UcP/V4AYHzKqkjS2BfuzlSRrvBtkErYGi0vCxvs9dW
Uy8O+A/dmvdpnu5Dvb2I8dvn6vsAM1szyIvD4TfOoB2uTjjyid/w2u84dUn1d08v0cyT/vpfD2GA
YTVjdd+aPPq847VGXWteS8/t1Zx+I+roz5XgiK5l6YuK1OsvasSiaoRqfDlAH1lApXBweIAdSbuo
kIjTG+DSxgAsr6QmhGjcNd0bSJo3eNNznZ46BTELJbVpSe8lGfWqAIB80nyFwh8LaRojPT4VYoDq
MCwumc7x3N3K5IUIR66XN3Ev5sOvaZR7lN8XpAgWMPvyw+ydOajNoEy38cTqIUZZrVNHPNpdw4/G
UscMmUtugaWV+vO0VtirLIEI8L5Ms8Mv1HB/OJbuYB13/C2Ghh1tzvSPF1ZxdaA9e64Iw7oX2QVV
oeTGbW8F4xB/f9GgJYoCc8rKasMzC6xXfJlP9AY2GU2e7DDpAOspOiYUeoEWmrhNV0B2LYKYJa0j
dD8hWAH+SxrAH4U/Dr+raRTL3ziKJZs4+7RyjhxxCz8Bm6dhyG8zqvii6VKjQ0YReAZM6dE4WsT4
ze/kch+UvjQhugGt8CxrXQuBpx6SjQuV1KN5Cq3b63C0719vsHc7ZhZu4ZbsGyydsBnew71tEBIJ
U8UKKZVYmk1K21Min5SF9nkNohN/OWDdIpXj6Yn83cC+VvF4zeh9TI7oUWX1S/fH6ONOAemQwFir
EirnM4T3YHlRxTzcPPZG23sxl7Azeac+7DH5ZojkhmohacuBAXZOU+SpUK6we4t4Mfj6yRXlBVOE
wrZSY/MfBKYNSALJ7QyM2fW/tED+L17AMHUEQSi5kwcqWgGtKqjI6EPhnkS8950o77tgYrh8Nx/y
Ws55AFoTnzrbII0Lvxq3tn7H4t/jojbdvrtZVDVYVuNjlf86nJTm5g1E5gpkIVVs2MixnJfEC+Ty
wHXQ6x0728QCuHqazUQ1DavQaETJIvxeJM2nR9+XqhbgiwLZCk8qzq57sWMNfvibxorUkCuhz8w0
4yJENLeB6tooZOVjN2UqA58DEXVZbDS9zP8lwMpM0Qxv9kIvWOp7fJK+T/praMLT7t66COvDamux
aR2XFdxGzJRVhFQBYD9nNrRUp08Lf517osl32f0HAEHl31dNew6jff7xDY9JqlHm31sD/QrsDBux
9k640zht9CcNRgbR++MLNI9/ZtrsuPt1ud5ztxnHwzWREgMXJ+CwM/bEl7U5bblAsAyWtctC4aKV
uScHheNU96fX/okbtRQkCNoG7/SFX4bYAIcz99BCEhkBNQJ2trvgKKfpyk4XUcwEf3yW2pRgK1wu
2vcdB/nRBUOONqp5xhgwGtH/AWR7OUXWovfGlK4WSqBMPEzxB5O4Xrz+i/iQCBPI718EXu9Gvwry
ETx8793Czhsf5wBir1v/JWiGiYuX0oAgO3hPHcuDX4A+twx/t4ACGezTIZptr8g8/CAHqlu6rrHi
QdyVYqLj7IE/aWpljfHp0GhnQnj3ofdHN03LHlO7hj8pgO3UyZUrS/9qoDwUUAe5x1htBm/OFEWz
e3FR3n9NhLYuI9qwE3eNs/sIxZ3VT5mHZEQsusHCMPz2pJexOY5GMDEC+/+KxvxMmApgBZGCYxv0
YR2paXowYV3vDnhGMjj04h6NnzLguh1mpvmreDL4h7Y0NufhFFC0F5Uov05iDWp8jCUwPjZ9io+U
9mbpZ1OjtuugVaT77Dimqo52mCCrO9D4I0r/L7d84NR/fI/+lROktLE37fsGktVDx+cymgoRlpSx
KzUHdj4z6UgtLEJdeLgYA1WfYE193WwFMvmVHNfixjgAIWZuwFyuArmIAxEHLInnMVAQ3Ronod1Y
+tt36zapIJD3O9joBEGnua+ouT+ypg1dipVfa9DqkZGhrAWpaK8n3Pd38YTBQz5mfJHNHLroD/6X
dABkHwLtLefyTP2V2cNHRG+Zu1AX0c8mvVDPfySXFZyGJ44Wr0RNfyKpSvw5GorO/vucKDpI2m5M
G2LE/fp+C8eH5duE+OL2GCQsTpMplC61O7Hir6EZrfjTo7LJTGgXZihvyGJe4y71ouWlsDtJe2XQ
me7UkEEnzlkFEXDF9DYtvlG9n9N7mXHKQuI162LD9aVyxi/4bH8wqWHTfthZgRTnGSFWBchUlA97
nEcqp1/+GvB9uWal+AACLy4Bylhrh/ifnBHP/IBECx08hrHFuthTwWQIlNY4SQmPk3tUVa5KXAn0
C8OW6MWKj2ciU29/pX6/iufPnjLo86MpawjZdWp8nBIhE3YTBf3CCKQy/t0TZFC0njim90i+qSex
DSrEfN/sE2JvX3fL7pxctSBHy83BzyrmUpzkQZqMV4qlyZIrmCLO3GDugG+HhlsJjT+n1oHtQW+7
tpEb2GRvPZo+yvBQLFknhlCZanLu6p3LFfHmMFm8Jz6Gk7pXx7klG6xl4MnYRmecJbd2GP1UFeup
m+HT7RHWVEk47U888B7wjxZ/q/iQAeUS+kjdg86YynaXvLXfGTaxiGcGmL2on8mNoyqG1VHi7+t2
1bCZtpmPEbXw3SFq8uYuXRq0y/Dv0VzVgBdbfSygkkHHVQYs935Q6aUQAdQjxaXawk4m/ntzRwJP
bEbUdH/M1OALtVaEyRYo/z3OAbhv+kV/NZFfwDD+LZZ53EevOwElwzRkFQM3uVWu4kx7qx9Jhzjt
KcSgDf8KVW23nqVlAicn4ES6QtjUMToPVvd+uIfQIlU2iH6XwuyUqKHGb0WhchP+1DQwNkC9Wb7w
KqjPiXrpg+nNw7dk1Z+OjQ0g1cXyd9yoPVqBXth+GVcH/qMvyobvaOa5rvbdQ1b1CzchrgVZYiFS
kK+iSKLHUVb6i1xiPfJoL9IaXawYZf4V4OxG+uQB6j8TPy737DY6fK24Dc8zzQ9YaYpvpVMA2XMB
wyyPC73uBysJk2I+5AVNWxT94EeUJHCWnVtXELdwCiOykIudHkq1eTQDgx+bntfDFsmH25KLwK7t
jkQpo5Aqf+41B6j/vb4hFD2eoGTF+DxQ+cxOl1NbzzYGeFU59WkIh8Blbd/Cot0Au9MgziqFG5P8
2wz2WymvDxfPlCHi0tTcfQD2qhVRpWSKRN1OzYoWDpopFFgYI1Cb4z2jAQJhfvP3Xz3kI3qv3sBg
6lx63OHF1Tx1XYR1g22BeLntrpSXEuIupqTUyOyxfRqPISf6n4OBxn2ZxgPgxNYpgtI5eBuLJ14E
HHL8f0O/7ymlWXaHgMKpp3phKwXsUmWlHYl/vaEYNWeK+v34J5WaQJuiHNAi6eKf0gfbVAV+ix/P
s8poeWKSmuZGDppowOw1ySVpoP5O4h5+NIlt5nawJoqnSpIxmefxdDk1tIOzDcWnENSEO9bpc9oT
/np9hFSf8mMLQzNkNPBlU7OL4PiPni8CuiqRTLw2WdTM61h/z7VkDIPNSSA8+JVWXCvbF21r3Zn3
b7mRsqnHjYjjU8uevmOCm3woptmq2FYiqDzfJTD82e1ScCJwRh9//hVFPMUXpZXxg6sUnItW6LcP
3R2OUldRRN0t3zKulMw4gwy0JKAHl3vSEObNm7BUw7KQk174y0p73FJXy/BOuIAIVshkcGk1N+Ai
rI1guoNcJS2CT8Zh3Q/CpQKHLpY8hDGGRYdEsCYLoypEEXgEPTqK72twDEqU41occVn8hd276vwU
Q+QDb7tojm+Kj2EM/X8sQfHQY9j/268ev+vz2H7h5NAaWn0c2is4MKIlEWzvVLkLxAdiKO+9/r31
yZlIqXLkjUBjT9LIAXkbtab+IXzjsCT8sYRy8vi7IdAaEv1IDxlW5ySVjiyIizFTbrAbCJf5a1vT
C7CoWou/+QXXjgKkY11q2wXgXpxG1aKaul6TO+g3LQCxuvJrLOAJdrGHSTQlrsa3iXWD/yw9qiE2
CPP0MBqBEBSlpqz0SEa32Fc2+4Ivo0po2h1G4lXCY+tyKwNVgKELfUViMDCLMiDEnjm8ftyRfGic
FJ3dXMGoRq0Qto2IgyQKqeFYTTsAYEealyh5MtT9ba4VYcsQ57nTtiCDnL5mSA+j+mxsrPHmByxu
+k6cd+0Mc2xQBNeYvxtKFTzJMRHxLKhToXObCHhH1TalQOMNBs++rlKlf7cQD+8DMl2FeBL+Uveh
pE2bCmk5ylKxmx7CPPHznHkXygptyKV2qJG8X0JOrXuRleycmH3hcMDjgJYflyGeXW1pU6P8uwNz
pd/raKNgkVSXFdYS95YXPUuR+swnKsKun+0/Lnjn+ZAzQ5l/AzJKgnfX1u5NR31OfeLHnKQSLUN/
gCzcD89Ixo0Sz+ntHYUu+sWVpmEs1G3TgNPtjIM7cLbuOcN6lQqRM7jhRJW6g1GdwP0WEBkf66hX
E0kELNEvnmy+m+/TsS3D4BRDlghlUEQQPBlvuLUrj1Be9m0VU+JYRV5r3KoVTwD9C0wY9d93sYdr
79LVw14Uwa88qDhilml1tBeArWhN2ktsNBYV9erz/13XMD8xKg0BjgLevRaE4pFH2JRFa1XRZgW5
Q7NUaKuKKH5+DNyHKroe7tjyO3bOpCNJ0aRhSTuRyXMEAxHrIpwwo10hPDOHDLW14Hmfg4KK+6WV
5cyPn6jwpAVZEXSd/hZ4AvznaLgfreMVRFbUZspXlVyq8sA/tF5C/+YjChqFHWXEupHi+UU6OUyW
kMskwdwBLtay7DgAk2nVEA8F5a8VH3Pr7u/4WOakGaEC3e9Oltwf2SwLcNrcl4qOYdzs8PWmqYhN
jt9Yp+ZRMAf88uNL3Pkkq8rRqrILo/CK+bdunVP2f4QszCiumsxpZy1f8Xu2cdH84aAxYheBXlVv
cCNa3ZEecO190stouo3chyOiSnItswUf7Nbj3n/XWc54ysPEZZkmLxzSbFpNbuqG1nH2CcUDlJ/3
pLZe1ToQgj9Dor2jyamW069fdEJu8GBevDg4RQLI24qBbAj7Xff+9ySqlpDBwRtaYT/InadXgzMl
zNCt7m/nehDS9fK8YVFGxQwf7zCO31wflKz6j6hpqg5s8Rre9WJo/QjnVTHg5IxfidHEP21QvZTG
a55BCc1mN4GmhYAnjF/8+5Dl+defQml6t4QqW5B2AKwAHL295IS4DE0SOwUEOTTOjaYNAI25QocR
geoPjSDLpQo7FPXnQTVcPuaLK/PSYga9+9r1IPG7Zlqqs0/qNr3XLotDmvODs2PiMEl4unxAf2pL
xr2r0njvniRytobCWFZT0uIIXb3Nk+KC+NV7czfQprQjGlRAkfsFUwrcrX7LFo7li5HxqYdCCh9J
SHN6/KXs23Mp33CWhCCbguxbMuihgERVg7UiSwXR6E5bpyW86xF+DwkAQJJmbNvsOJgOyhD3v1X+
yCuW54w0ReKs5DCftvycvYtuMaNywjIwdW7/7V9eMJHdrC67OG3z4Gtn20vD0QiG0vLFPaGhgD9Q
UfF8gvam3vRreJ6llEVNIs1G5li26hU5Oa+nem4gvBHCG32uc7rcDe5KraWlhdr23Y2JmmJrf3Q0
BOZkwRh0iyVAnCEyjmdOjNrbAQutlHZbI3R5K7nuwLSedhUv70A8ZW1HCLKRFYv9J2gyzDR/G43t
yncFEU4rBRd4w4AwdM1zj4dPhMHIsnDpbs5DEhsz3gSrvdNfS7t8Tt4ZnbY33dY8aUXW9d6NzB+W
Dl3TenGYOy6b9mNmzTxqu6zZ0U2RG12te/Mz0WxgAdA4xBr4r+lkI4Q/wd5xSoJ8dZkKvaoOhrQo
bgpY+/lOJsTq9vqcu5QRTewaFZ8ews+bx8vSrxfMffgUt8NOOFkinYqJyAjombXNHAnu9S2PHudv
9/2Hj+tx8mnVcV/s20dCrvOosuASEPhbxfyqf6kzHF7/iZo2E+9txMnS82GP5Inajb02G5fSDcHV
0tE3MRc7uE1Qyc3kvqmdoHchy46kva2NUATBhHmZGdPiy3ndRZvF7B0OTsItPqO1l/L+VBpX1pXD
jJYxhbcJHdKvlJSiPXVANyCbYc1EvXvUJPmMX4H3KxxawBxscXKrbxUc1m54d/eVfI/AmhjMvTZ5
tbZDe4ZAMyH4fFXvezjLkNYnTQS/uA9rp8Kqw9V6RLc9XKAi+RVeHcAqbcwadYNgkcHazqIvr/VU
o313VOzsuWY37c3csnzAWIyCqp45Lgs2p5Dc4reJrAnCAZjV9CvUwBzdXid90if8pvyR8hEyzBHc
SF/j4XRf667vxD7FAyxzYeGVwfBxm6nsxCgrlgn416HcSlum9oLlqxKom0SQYG752wx9VDsne5kw
/5teyy28loH13M+v1/0kvSOWAdTZEjeRt4XObmvmme3MuWoWJDDyAtNmJwY4b1Hi8/KpNbr8j+eW
TIUZPK4Vg1ddL/6e4AwlbC1tP8HKgrofqcTc0+gurwwm3vQ5XbWojGVQSr17JilkN9YGU9SB65k+
yfNrZpMXJrSO0tME5u74qwED/2/bi3LqB3Z3ZS1hmkL1tdQWkOZIzo7FgOThFYzYmoXlM3fPt6A5
NL7mJtJwmqXK7+hTz/bC9xzt5IvfLZsxvIE8NUbEv7m74lXJJUlSBS/PhfFBHFUQgHfTQfw8nrZn
EyAYog3XJWmxKsyQtXfU8/6DqukdeVfELN2rDjaxtfZpWW99KoPhOMOK5o62dHTD4OhH7W68SFuw
8kntA0n7aUUvnMwfnmzJBZs9Vugjt2mgfHpA5tX/Xi8RvpGGX6TwOifbYvGTU4RTkmr1DN56D7Wa
nbQX50wPbX1A0VEYtbzKFOj/Qg2uj/VKWBpiJ7QO8kP2Nx5YL/zF1LHuhvUwPu5LbN/Kke6blbPE
QHiYLTnhWFYf3cOanlZuUp7pGspbhUxsbBVWSE185UJdeHxUf/CVI3MHfNHx6itf+7p7lz18X24E
CPATBF7ZoqMOpGag74CROTYOZ5TAf82uXaqBPa9RZi21ShFFEUhH5i+uLwUyO26gq6YNstSlJe21
VAHDtg0fkxNVtTbfQf7+I2nqWjJTPZKn/pCS8B9qrJgyv/CWhZB8LJ5Tk/cdW4cgm5OiEukxpQBD
wwmVXIBLrpSF2OYqR+oazY33WBAzqvxZewFFfqzcdFKAp40TqW1vJgYY8hdAIXNsTn9QbXS0o3bF
2DgMrLcl6TjOIkH/+xYIHCBTpcSsh2dTatthuWo1FwmG59/hakyvbsnlOw84GlLf0rHQAMWb0hyc
Mzjohngn8HJm/QraPFb1RaDmnQ+UlrKvaL07oXdslfoxjgePG4EYgpdYANzbi99mg1jgCTKZJtaP
jcMdrHPeCu8ib+iYl1KFUjKiD5f01gCuKfC+Pv57AbFku1UxC/JfSP37l0SHw/BatpBK0CxnEPi9
40jBL7WJJ7/GCJRvaUyg1cb3SXGlxZIi/VceEKGxdryf+YUSyb7Bhp104hOBYS+0ylwQEjK62qMx
6Owqm9zv+9VCeZqVLHA862EXzTnnxR/FMoOlZkGin0n2KTSssRdseKBrHVEePqKkTaiIJ38Pm1fv
9oOpPVPdWmqnxzoq+LDbDfa3ssQujSTDKGJOZGwjs2oCLwremM4JxI1FzCjRxyls5D5X2ej9h4su
6/uAwnZoxaXfu6Gy6IO44qfC2Pyk72bIuHXqBhnO2jWDGoBg7/yYDzRj0n49hC/BC8w3tr2/Mwpa
wdNyc6bUXVgf/rG+PPAR3qLbnP0Gx+aAGlwU/8RljR3scCMShI/T3J6OXt8Umq29pGkC3bE4fC/2
JrPQ8Q7f0jQlp7ZBMwIShimTmarKAO9mTQ2qoThfB4160/MyVgFMhXZIdOXN6Z7vRE0dI4cOpXQH
VZVM1khgBlfl12JucDK+oYvw2d+QdCI3+TJ83JXUgrkrv/veEwa0dAGhmpNsFt6av7NtQ6iJjXnE
SyEvcSf0RdmoeFySeC+xGBLnqQBMeOJwkJApoLbQZ+3jRkroQoT1HTle4fvmymeNrr0TwV6tTAvh
i6Y97uXZyWcFB/5S48nuqXb54uCl5AcGPQ5GpgPSSWfJwyHKu1gT/YnPp0ZRbqT5gdPcILcYnuZs
/x1B51P1GtapC52p9TJsBGVr3dIfmTsXqXe4R5jjumGZ29WGcy0ooK9WVG1SlXWb5gMaWnhLPsiq
gqa357fZvWW+tIP5BBi+WrwCU7wamxwjJKQtU0w98vgUAjiNPujFa3+1M0P39OvEzw4Eww5/bq5E
9tFFdj4bYxtvhH0NAWacvdgPttHY789qFxxwcUD8Xq5cTg4hv060sH7uu45yKBPz7uvaCb6F732x
srCe3MixUEqFcJAU9OqKzR+ulUNcQPVHFGeA0Ke2Li3l+/1P074TdhGmAqK0lRr64mjjoWtMI1em
Cyv+8xF6mr9OoKJgOq32LAJwQ3svU+Y/MiZUEgByJCLWaeNCSlqLJeNe+Lp5F1HFNu/Mzc6ozNzA
K9O7tgsmwR6pVagHC+qVEaE/MKc7nxmC8wD7LNyuci5HH2iiFtCanIEq0ht0Viz8pUpSKZ45VpvX
oEGUOP6gz8b6CuItHD7OYIo3hBrCTRnLWU+zg1WVcsisXu948xp+LNCQcBRNAAUuvTLYBsMcedle
1xQb1DPJR8z10723kVNoPforzoRDLbXRy2Cr3tH6e3YHt2l/XbXLvqHOQyLUMKadZla+3i72GnU4
olpTfEwM/kROxL1qHvjsAR+JjnmNjLiqklRRPchDEZuns4BcXwRLvL/aFnJJnRp7Ksgc66KBGVnA
I1w/NcBlO109K+OYQz7Xw/RSPgOcO6ZaKpa+e9a2o2VquPGo2iThf20ju9RJsw1Dk8TQGFAd9gEV
Ibyo2rL5KqECGkm0871nH4PoDFJd8McnXaEWeYwLbRQTF3tkr5xdD/uLqVv2/3223ILnb5DOaISg
9TN+p3RQW0s55YjnT20BZFBxu6P5EnMHf/1WR0gJnQGfRdk9vEtpfmDXtMd+qqz587kWDIUAb7w/
gY7U2Fd2OciHxZ/4kfgA4wVPdJkxNZ80NabPc1CYYfndZexr8gb2Y9moBPJ+PNhbtpKAaHlE9k9h
LIqi7yZacTyEBsp7EdcsrZgopk8oDHk3i+czqPKuPgGUDgKXSf1qlnkxjCqBN5gRoyZSA1L3TaEb
dywdGQ1ej9Pqnq5eCE91BeSP5S0rjhQqpsMHye29wIf9tShh7cZ1JxWKtvQDtKyVkehekqhXYFjN
SKDN9o8POxWUVOOWaV6RbaG9nZyCqzmCpvwQ3wpqhZqrmGSl2ZVILSBn1qm6JWv7xxA0ejp0lFwY
J3mK8aSuGvIEmSBG1NiLK0onDU2brQc5sF/BQCYS8dl+eP7Lr3ObAuJiqLQX1hDnNa4hUIREb3HQ
0Qf1hJCIt+JFhYEn78P7XUgGAIvghyJ9OLLq4iqFnTXGL8ZdtN3s02ZKWK/StfS21oPjHcrBGoRY
cEN/WdAECQpGvekfc/6fMHahr2wawlTP0WNUG2+aqDDUDtUALkwc3PKfe2OPMUixwLSSRZd37DCc
66gV9djny0NQVI300J9AkzY68yeSifWhVmT9yLvT5XaFqrcgEP3J5xvW7X4UJh3Y433+yTGCxfGO
E0z+3oOAe8BSmarCgiR/Nojh6TKsH0u0i4zP91SEeE7Amzcyvad4jXtBB7gcHqHx9JeDuskRvdHw
LFlQd4N099mIAi3PGMJTaJOQwEnMRZ3n/Rqwgpl+sSajEZ1+tV6iyBflu82MGtvAjqoZ6XJeXwSR
JDsoUMd+AXyfHbuq/xPCStXwNW7V42VOGBPQaRUjtHwYR403WVhqGkRWxTBSIti9b1M2vANa33vK
dN10EpYb0HZX/SZZ1zk/EhEbre39f+SV2KD1vcS4MFSkoX+2SbxhKKXx+11uuaE4yB7oUmnYquNH
I/gmJKOduymwEP8PWy32+Ifih/XNfdtaXatplJhUjblkYA1KlHMdIVxuh9U5P1EUY8CgU4oV4whz
GTGCoGCmDdWffLAR2p9+QORZoTyO+WXvHRCCDj6dA6SHaZNAPws0EC5naweQgnrYPHUhVLezdfhs
uvWOzw0woNg5cUShLJEkq0APJdzXvs4llWvlVFyEaPOTxziuH4rFRAldIlH+r1FhsbFd5Ct9NBKd
u2F6nnz4yvjHcDJx83SuKuw+Ycg8zrkDTnUCRLcU7kXmA7nafcpM/96NCR/UGFI+Q6Ow96m1DB+V
IQPzVxBWiKeDyGHF7ZdUngTy9haSfEHL17rN51cxF0sSAa9bDWWsqyesHFnpJLmctxh+dyzi0QF2
0U+qsPgJ8ruev58bZk9vQNbBC31v4EL0jFefwoVx5DSkSkaZjPsh/k6sxA5mnYk7uNCFix9KuDsl
37QK+p7SPCZTxKP+Rhv+Hx5E9vGXx3fCxC3UM1//Hek5fnZ4zK/S2AGlE7EFQ7+yjxyOzf0eozOX
MrNbkCLQP3TdZJhdYuVHXS17nM2GaTSAQY9uUjyXk67KBBnwbWBQF2HWKGQQtqw+zUyzjfafaHB3
RqzzWlGNHviwJ647r4LlJr+ELa1zcRFRp8om4KdVLGV0AyIIfq4V7t3dhBaj59BA2YFzOmPN6qlv
QAA4orpSQcz4IY3qy06xYGRN4i79d56pwOspPmFdVtdAxVCONYULHN42VZWCp5Gba+2s0hVmW72/
prWRyhEQU0WZCMPfQ8jj/pzesD4Plyg/ybiEuKseAb65gEaCLKCPYDdSEy1EVNoUcVUO6cniTr4b
r3VwFfeLDILMGOybNgM5AeIS+KwIpKrcUcWZADxazh8PekhEwzMdR+Wx/IvE3jLFyMEOnohIVkMd
iEWl3r0hVFbwRzrf1f9VYJQROeKDZD1cqlt6FTwcLt8uboKs2r3ABITb3b2KpUSYqwyMQ19vphZe
b08yaoD9QO+SH/2P37U9aibJzBUTSHCkkQqDFzkTllrtecczuDx8HQIzO6PEKFUXysCkddytpXpf
y3P6OhIQOmv7y4ay1lDu22gBXH4mosUP+XhuizL+YeVeEjtsMca7sJoHR8mhR+IMsEfMNcwhjzsO
uMwTv/sydFAH3dEfFCiIQzgIBcri2vIIs769c+L6zYpS81NXuqm6QkgdBTioZ61rukh2GAP+2ZF5
2ZzhlZ5szGMjW0p046Qvf9OInXKF/huEhHf3I0KmvsnEbsisyhFTH4gWnOUv0nbkmyttxUNT8+yr
HdXM8Y8S00pRLsmPn88iPKbXv0aQBuK8Tv9tpnOQ/r/d/Iw3RSJnMSmuZtW5T/Bp41SQTyQzqykP
t0l1Q243SkwZiXU/9hlZJFq/TGuTYjVJfDw7rXnqPcq0y4tqh8a47j/pW+2rafBp8eUssT331lmE
IyN5JfCz85y6Ci0TSza2hbRU0mXeWu+TPrWozMHDTzVrF4rB6alH8VnVo9x5kPE3xETHFWEdkdxh
lBMQrhJzHOjJEvALsY0Gx+CPA0mddU1tYQCedWCuYyk9Wi1rIwqa2+0TTcFxLkuEnPulPn2AQ0Ig
iCVrXK9WkN6WHFasjXmhhuHBW6r+uvH04sde7OOilly9ux1Bq1YLxU5en1hXJbbqpvxpiJrkIsDZ
3CBbZRH1U4XLquchH3VMuwMS6QjNw9OZq15c/VwJI7+8t/ViZd8ttj9c/4IC0n2CQl90caKyIARz
YrttYRSOwOppKC9Q8RxlZizBH7Ynmm9/T6Cy5BgMFkNuMA17RBXCijEP+o/CjUniAb4jzfmWrHBl
TaHV/kC7WBSzuNvfkwN9F1ColZmXWJio4LU8I+PcNGbeiMS6xO/ddebji7c4vw3gzaabKn6jUsG+
7yAWYfdIrnZuctYzYMsyfS7yHxmV0O8SZpzsldZZj2wEzoc6TXFTqeGkUs6iZprWSRpNoAWw6uKu
AudzPUlXcn0cVRODWnQiF2qWN7WsTN5+mkdPVxYZDefb7+l9ujT+rEIZ1GmJUUjKVdnL21KOGAuI
xxBcRC6bLvNTw5olEsAmtWDA7+ptGnQ8YTe/qhSMJKphoRBxvUJJSbwMeaVT+eXaYjS4L+RV3Y+g
SMx+IiklE/3qHjEQqWYS4Gr6pEPU31ONCtWLeLzRzFOvKnyitlKpxpmTO6Ca4ESqF+qxeouy/Z3j
STU0yln9THZkKjDaRyvj2MIG6VhGe85A38ddoEYmd1iUlUGAYC09nwUVIk7GD0m7gYauPO5iY/xs
Y4PGAOtG/2h6uwhJ9wsBQDyMvX7fvWfypmPEWrlhDud19yQxNYN4en5hEGJjJksL3N3oqGoZtoml
YMSFnRF4IhOjv/xzBj1U3czMtMWZzPWqXEt7nTz0W49+91RI5GNdXS7mkceHx2BOUhLB4xUAfCbJ
bCMI7cMkThouquxRUVXG1NorXXf6aDNGD9xVqfSqTAOy/T9rj5azDLXRcnqmOU/KtrLEn5YbmuLL
hao9XiOQiXqRKE+zAB5bx1kAXHD4kLSB03G4H3M+74u0QIIqAp0oBdlWzoTJgEoHGAZoQxPEsAqy
7hdDD/UcIQHCwnfk8vM9wCo3q4dq5Cqq/vycbiOmAGJligkv4oP6eUS2Ybl2KC3/muFJoU0IeGe9
Q/HByVaVZlSH4aGSwqV86n45wWJLzbdF18P+Kowvyig3EFYWXBMRzZT3c2T1nGDZle4ml4t8yiiB
VB3AATwdJEGC9Pec1b2rwawzc8edwfO5FBLmRsJEcgGY18fCbBsf7ghbJebI0vo8vGYaQ4Iqv/KD
mm3AmvfFOt2s+SwhyfQg84WbzCdRyosJpJ23jSC9eDxnvCEP4+/UU9XF1Ub0odzxnQRJnKqzqcQI
y1RT5CyS1PXXti1aTJ4OWkU/qFWkG0j5eewW2pME92YWxB+kFK9R3wRqvjsSiuMxmY0bF/Qdvxiz
sv6gUmnZWi1bcJ30l8VkFJNonzO+our3vPFsBMZ59mlVK24B09N5bt49mt5bWSdjy7DUsUgskDl9
EvGny8A0zoclthXiObzXs70h+3f5KYkWiO16UNk4hNPAMCGZE/u+w+7V5rmHsms4RyTDc72EQnxb
fA8qlhARtFdbQj5f3obx7gUIxaa5AEy8ZKyoQRwQsJ19RpC3f6UN+shTM3sEh9QSdMrXU/T/6hgl
vjQuwmUw1UWMVqX0wm+DL13+R3uRMnmU8pvLe8Q5uESHdwR6fcWj21KR5NQYgFMiVvZJsot6Jhzw
9MsMXtBOvAN64FMiJCc/PN1BWCcajtlowEU4CLFBXUitYlWT6wW3H6Bv1oE5THbnfKsktrl4mKsP
OTnrUl1nr1QQyDyasnBmY+Xkp1/IYUSJ7FEx6UbVLxYvgUt4gRr3vBq4axU2I2oSmZnfPGy6rGNf
HsCmuW55NJ1p1jPWDXnjio+PbXEv3s8Dcpp53jRLlqCucQ5ZgWdSwfZKb9REoMa8hycV73FAUR21
tSlDJU9WWoUEp4MRl15lo8EOJPyTtTyxG6ZMk/d5exMDKnv/VhKKP4JNU1eGNpggdEfVR9evpT/v
hOus87eIXDyUU0Sm3zsun2ambVAj5Vcawk+qCNiQKvR6UauTlAt0RT+N1MH3PB26Vupugr5l0BqD
K+8R4YbAGHidoBF1tXi5oe5uzStjoPufFarqSl7mu5lN9ADwDRCxubxKCjfe+EITewclq1I5hMjG
MggsY2/kG72Qp/lOUdHB56vvXp0BcG+Nd2ItZuLxHGXhHbQas6FL8bIJdTgUTXpL0J+StfAan8gO
VYqVVdCFOLA9o0dkC/qNy7jrUhg+d1W3IFLuFVBX+urZ/mt00UTYcII0zWBdghhhdodJ0qqGYERp
5nwJgmsqYcgcfDkTVKudDYKz9RkYTGyVEGwJJzvqrDDNC+yzi79U6TYMNQ/eQynoIT9kivbXOXZh
CyIbUkGPipXNHTqcFs1E/qENf6pAFGsn7FMPrn0L3XRxgrKcYqif2mCtg/4Zlj1Q0/dav/0yJE0f
y3oXp2GBqzXE0VNWO1AwJIb6mvW8CBdRhkyGpqDLF3HE66N5TgGSv59HR0ivQ9zkmDv4deovbXsQ
Jhs+zRoisjW20k3kZDT+gsiz5nNjIE9j6qs2sLlN67IitAnXf54QgK4HSQZdFCHgGtfi7cYmETe4
A11LeOGoX8Svc32OUMpZzT/bfreNERHIsUdCJzCB88kpej4tW+3Za6d2V+2ugq86bI+SEEz/wp2M
CmNfHoegofHGOb3vcQC4u7apBHTSQ0uAnUpigxXF5tMbXDcXfnbh6yu4YRyk3XK3zxCNd6GXXTX9
n8X3SyO1cFxwFMCvZYHcGNn1FrQdDvshwJdviUvG4mo0DPLPWLpurPFWmtpt5VwVyxT2Bp1lVIoy
PmPUFOrF1jlaxamwHTzfpe1WUAJkzpF01xmAx/BW/Yxd4MCMXBS4VgfJPn2lo4+/hN9tmgpiOCQG
jPbirera5PjmQ2PjETLjg+Ot857GEMVao5yeGu0TBnMnfWa1lw+gmqgbcnvf0zneCP23arJxgmIr
IGrJrlESXIISZ1rKG7A0t1cMTI1prwFN8RvDnxJWPeDmIL6NA+Jzegp1dBn+uS5zehFivDxo2qfA
xGo0Xsa+5CsHGfVYLoP+04Fgb/PB4KVRG5Vl3ybpl4XGeccok5K3UZmqaqfIWV6418ZaIGu/nLtw
nAcTuh5qKY1jXAG3kny9xDfhZbQ3m6eq6kkwBUW4+OdWQ/d7kuba0Re/yJLwQWCCVp+M16AqZHB7
eAqtNVtB8b+soMT3PFsVaL8ItY8FQTSFkKhoNWX9bwvBugcf+8LpiYIHPtGNjsRAnrdtLnWu/t1Y
Irfwnx+muw5x7Tubashfpb3r0/m7CNS2SUPCK3vsyRATNyDxFqdam46XwUV0+gaEqeOH+mFRevwy
n/4Ik0dx38UlHtD3hFSJitIq3iMZPIN6aq2z/YjoDBI6OLKdy0gJ5KaXwzkJIVsOcbGOYVxGymRC
0b+DyViBQ3wD0gBsB2exyYFHti5GkfdSIyizLh+UajLTEz1X9gY66bYUnfcBIjNTyCkF3DR3Z62v
SvFDqmjFDXforzK/f2SXqLvWO/iqPwk+jWSjQstfu84ABYAQ1XHxq7RfiaLpg/l+MNLh6+Gccdly
aGjUh+sXiu1gnqyy0xa9/Z5QWS4/KQN6Ewihd75CymltMi3HH+GxDvAfmSf2RxxMyet5sJOSNRvO
SRmVdR5AoAP9nHkA65pG/XLWgk+q/AGZAfDMh+FFIyVm+9SvcIcpWJ2aiG+FAhFKSMfgHe33hxyu
EcaW9ydKw0eeDblsYmN1wm7voWNIZw5HtkYIFqhlu+bZ1mXNJmlu1X2YvBKUfrkU4uBEuJAGR7ti
2+6Q7B4SAi7F6J63QVdlpkobiWVavNlgePzdGtnLZgvgT+7MS9eKJDEvMbOBuWVVjyw0QKBMVxTA
MozI3Sgca1G/Q/JXzu9U0mCmtzm0BR25KRiO4c3XeUEIsehe65P/gNO+nGcsiF5DnhMIhSLVmtbQ
i6a5c0idbyj+JNr7r3ZSey0e+gebJWY76DbcFSNAPXI18xY9NFJyd/1SekFp2HIQpcPfYTsc41qq
u3ZuisOQIMK7zM949zmRKe1DMdUlraj9DHiZIwkWbN8sX3yvUIsDn3QYHUEScghTh/kZL2lRkinD
pD6PfkzwXgihR/4NdmaFxTNFaSORYKU8wk4qLSekEJ6RDeWWURTOiRwzUUKtCYPFv3HfM2taq0zN
Yl04l+msjWlgxOiNbFpdTE+2BnuyZ4MbM2nvYYASSXF+EqIC8Y5s2FdbIjqPhclHDGeOgJsFJPQx
0LXP0AQgh1MeUK59wmWpqvY85vWgclR3cXIJg5BxQgO9SXBM9ShZEti7MHMW2B8AnkS4qxMcxsRP
AysZzLRpVvFIsBz9L7YSUgo+uJMRsHXAFw066rRHtdGWri93cVu2gYjp+/XsjsGWCJ8ydq6830bw
Y+wXbaYE0led8XkfFtg3gN0LNRNVCNQrXogW8nSr5bojhon9NPBQGVTlqgSc3yE7KYJMc9DOZmOj
j5AAdkUxfCnAITuJigZw1el51TVtNJbjDM4qk1fkmltIEwW4YZ7Icr5vdW6i1Thl5ftjhg+YCgjs
S2S+FhthAN5AptuErBT2Qt4wIKS9FOILLjQQd3dpbPJ37zvWE4uI+Im98Nl39R3rv0GPKJepy86r
lh6tpSvpano9KpWlwG0F57XchFXyHrctQMpybYWW7cjtWdhfClol1cOncCQsHsoPNVh08wJtc332
ii7ZIpHWdZr5dmbd4pnN7KqIom4prRjPRNG4O6FXK/oLp5u1C+jrS4auxEwRYhcTesCSQff2jBt4
GqAjCdJyXB9xIIJShh6zbZyP1YMAe8EZbNNKPWkJv+h6BsR5XHdns99GpgRgexZyqdvxkNYg9SMD
mk9vfl8visxlysJXDSces4IWqXuAcrqu3U0cNQwfOt7XLkHwv/mWpx8u7npI40TTCx6ORUfcOhPL
DUCe9qwCzoy0Mg56Ya6h4bBaQdQ0K3E0Ru+MQnY8hpPph27PFvn0J6B27txI8wfcFteiQS8ZFAki
LeEJvyJSNHDnU+zAACkCkxh3FiD4gCEjgZGN5eLiHi11JD4eKeQYDBLwKg51UU6AMnr2PSbmF3CT
xxcSkGO7JiZqBjVnBBD0oWo/buv6LefaH2al1CxFBXWy/Inwe9gUk2IPOo82rXaxkFBqeppg2h8b
DGK9YU43kdZquGTKjgcmmv0NwDr28Y7fRl287/Np9IpABmWTooDmiPBjI0gRGf1azZTuvwyTAZsE
tZlOPQQjsUCFhxZGocRfX3OmbciTOBKm4sRR9UnLzM8H3moiM8X56eIh2/70Ui9e3/gAFoinDtc5
RVl6vDHf0dB71f05asj/ydN1Cmd/gUs/nqbtmqTITMmp/jJtgfIDG/rF9nvg9zCLzuUcGV7la6FH
Ii15MuaL6xLCWBMdUgMg6CwCQL2JaoYunnQsZ13nMSXZ12PHkVY8sRwvBweXzhgh3TASIMCjr1Cm
ViMjaIMLA7LvAY8cRW5FdvRtgaWP+RRJcuYk0BjEt3K7a6SY66hFzjzhZcw9IUdxikh0B7clmrLr
Kc43NOol3XIFDpsk4uzWOIh5TIBks1+r/ExeZhcqItKm1PPquD6jlu/uN31jmp6bjCeYVjSjocUL
/ttx2A5dFuJXF9EgLDYkULwaVm615KAx5gXA9043OEPf/KP4Yk48R4xR0uIC2mWFEITXzfG813yt
YRH8bJ5eTZSLcd9XHu9Ba98iR0AZ/WwGx+uDpZRzDyD1u1NN03zyQiI1IoSvY4l5xi78ga1/+Xxa
KHj2In/hFeEw0VTxleXw0aDnO9c9jxNydWrfNurjad2djJWFny9+yf6cKChJFPmvnPFJnOmhIXEQ
/7/yTg07wEEO/hXZkfWvR133IgaE/wv+YHVwDkM8uPydlTOlgw3LiZWrP/RtTxqfoXHLJvm+OU1z
bDebTFzrPLITeVMhmchYXSzm2cfiPUkm5DY3GwrN+b0l0dOlKiT9h4hU2xdqyawO6p9vQ8krCzLX
M8JJORslKeprq+xIXIIPLwiG7jrYe+dH8HBEQTthJaSUNtqnQYhiosHAc6He4XNEaa0+FDtIdaxM
SSMAfnwlrJbTVNdSq9HAqtN/kQjZ3ae69VkoEd5SH/eCUezC/A7xfeBnoyw8l7Xb28JquxsdCiA/
3RI7GV0K7gGsJn9M3bRJ6Kredj6xhaByMkmIH9w57WY2CrUc69TQxyFhg9d3zyRAT2cMEmYuXM6c
b07KmBzP2+1gsVSFYnrGDvWosYDEh8tVJqoKMJ7egq4UgqBVULj4slRf4HdKYlbExYQEvmXLmgku
2rRB8QK528Mxs4ubWFMIpKUYT3lyFbH+v3A908G8H2OWqRgIneXK1He/y/IHWwI0LQ5L6h/n0MbU
F1RwpMysE05Gq4VI8saD6bdiAHKzlO+HVhq1sNvCRDLAL9YaTojlNfbiTx6HMbm4fTUyL73FYfC2
vZva9QhWgUBWwgnsIt/nbyPbCE28QLplfQ8xA14YV30h1YLBypMm6GLr0CcjlZaz3P0vDaARweV4
pduyWRVQ51kxNLQiBGnGqxzseNJ/L0bc4SSq5sNDExNPy9/8B20Ch/VcMITEhc0xUA8U87A6Yqw0
k93EfOORfNc/lY2IwSm1lK9/PKyZ4Xum5QvOqQMrIDwMae2TAQjx1TgZQIq3iknM2UymM7N0FIng
YPkORub9PV4Sjo2ir4ETibKWi853cysH+JSm4EUN811PlN2KbJWZmj2n/X/THY0rz/0k35V3HXc+
d11hSTH2ViBjCQE5ibsWtwLUnrqh5SnKuPNg3ED6T1QJW2KhM0Vg3p7NOOWbItoD8Cf0ISxqJFE3
OS5RuLxEovk7Sje6xnWtrSj8p+1/qYgFPhjLf9KPoCUrfCDCwD4gcn4NjGCS9Ln6dc0t3uyaGIO0
3IWAycLj0OKG6C5DC9OlX8EqWmC0NRr33kHKiNpslPv+ds6W7UDEz3fZUCWHsau419Vbgs63A0UL
S5A0/wC5iI5GkQCN+NE4+WWcmvDKN7B98OGGVtoiW3g/ki29OL1SSHxIy07n8jj2KSI+8nBB7+HW
Ll4M4MHaqIzbx0J0ekXjmAS5Rh2EEP8v22P1pIKYk4YInpnoIMJZ8mo7gNg/jklsRUtMZwVudn3J
//OcM1kgzvZToidy6P/077+45F/Vhq/wzFkkStyrVkQKzEzSfWxDaYWRQZIW+JoLoLi8nsuiBGAe
7D0QGcJ4gJrgy5VZb4+LyjPEarJ7Ylk4sgsdM/45hzI3ytTNcNQxA7vQccwluNx6YIploQN50S2t
nrY2yhcmwkAkZE7vcwCnoFpjwSYziXBRKC6M2W+Qiv3Axc90c6p2HHj8g9Sr1xcoDj9ZZMq933eP
fog87ok/koy7bIREk/k3nzxOCjFF1AuGisnwIpZlY0rotyiWi5uTjD28weJ/dldpWF62hcRi0Qlq
weINE2B/73IFMzUIsVEMnoSPJlYAR2N1grLd7dfX4+7tO8xodv3+FhHE/IPeABNGHfVsl4LjzCx+
3hksdYAJTh2V4fUF6jsxBDp/p8R+Kt+TUtvLBFxMg47TcaYi/dlauZz4rIUJa63CARF7TwHW0nUg
kOelehTsyDXIaZ5x3DfGogBRBGg9+3KaJ3y1wHh3VgulXJUxKavRpr9bzuO4O1Rqetrwq1aEIkJ3
kQlUWqU9mHjfvaaBbsB/VgufhJBIuASy4eZJDo8AzfLpKPoF4EtRH1unMNIuL6W71oI+e308i1xd
NRcBOIRrB2eMe3VM+emJ+3J3V2OBENGpMYcQHbllPjIl7rXrRsa13Oup77W+uW5RFZAuuc89b/mB
g5XHiEpo5LRFT15yU3PWYCZCiw9kwZDdt4aknZr9F3BCQFCewP21ixjM2PQ1hqNSD9KS0EV3S/T8
VoiIdNVhrcc7pYd0MWsXmaLDsx3iTaFZcynA0YIFNR4bL5OpSam6pUwy4z1nsfld8VQbE6b9THcl
sgQa44gEyOKYnLemzjFhAp/e7GTwyRmuc+W1QovX6HPN4BfGpBSyCzxel4ZB27OMSWjpl7Qz3jqZ
tY+RlVTinmLNVC+PR5Jg6kMAXd1jIgMgaPshfXU0wsPHgejJqX/1Sf7oZGjBvIb+BJxiCbjC1ao9
freu7Bl7NNuydMWAZ7ZIhcULTj4QIw6Ciu/dKp2FdUoN1S4p+xiNfZaKlddyjnAaQX5IcBTUfVpH
KXKXPn65GJihDi3ttNE2ivGQNv1k0uH7vfaJ++cp2V0DQb49FwRn6kdUhMxk630Mn3dU9rCnZIU4
kZd8EAtJ1ObOPj0VdJF3PjSCO2ccqnFAkkHc3hP99eEagd+XRRRzRxPxzTXHckXQd05awHxt/ZaU
tZ4qvYTLfgC/OnlUWzAEO8W2yhyDv/0e0iLJBIxtTTjpS+sNSqWVrd73QwaBLHltrK3+By/AksYp
/9x6i4mMMuZHzMczHeIR6L59AgmciEwplcNkbn+wdkTSga0SQl7hOag3Y4Ti1qeEFgdmJpp5iXG3
9itfJxhslQQiw4j0xpsp7VLRRKA7bdrq1CJVMq6VaoqXw1n1k1oTvGKE12VSLJ+3HDK7t/YQWQ/L
qS0KRMcMLtvsx5XR0MLlfvW0lDBg/SFPhvxdYcXGlYvBmOSyq/KrXdXj3WyLHXcoNqMtDNmN/KdG
ozeLgPctm9y+iMSq0D2a4r1B8/faQQOIo483cTckDZCDt/uia0vK5G5KvdIOQHeg8VPCrYR22oah
IJpLoRlgg7HNJkHhQY3EIwiIk2kZuJ6yce6RuDmeEWorP+Jg7AIz3edsy1cMDV8x4iP61bG7KC6I
2io3LZbg+GlfTH/KxNIksm6YKxMFoYwB/tPHQsZr8m8Km0EhPTqcfUNvEZ0wSrPpbhAi+GQ2FUTH
viLLBhhiOiYwrVJP751kqyshD9cdepMWZVemjItTb8/77jM0Js7PYevdZcCLbvLi6lry1D2VS5tF
1kKCEBLAQXDDYGGahfLG0yW2nCIq6v5M8fybQFWAUY/M22IQis7NTwEIrSt+JPhnxH9UgT3IhUDU
p3cjRSJZaXVDCJ4M97xzkqL6cqFbpc5Wxm/wDgMS1UHzxcriT40s7p7CyJmeiSUdUnBBp6JQBLcJ
4uPpabNKOXMXF9y5AEP52Pg8wHlpskwAwEfXqULJPxhaepHF6YbB6xnIWI41OnCUat2ojwt3byr3
fEmjTF0vFHp5i0aQ88sSkOa14P/QqPPGRLOq+D1sd250GDwnRKukW0CN/jyBE5H06BiivpQPV0yo
bYQo9y9dvtxmilWYuRFw/seKijX+7bgpdcthDbhaYkKf8r2xWbYogdQ6oxRpoKJeI0dhg/WuqxD8
pKmTSJfISuyGTpViMZm5hup1TJloTiO/Gqx2CUqhh4ZDKy2eh2K53/6+iga8WNv8ucymBed7+A6t
eW1kRKK+cB9QiKTns9DNi08sHqNJjFhGwNAH/1yJTR04cqruQfUhiBOFE+PCkmP/spe6SSC+JnJe
dxw18fCaeczsOGP3YIwHiWSyT2GXlMcwGYMwDomIxsxFAeHJsdw4w7GMvqC258dkX5LB1vAH1AkW
WhkjaHEpOvi6mtO8oGf7s4z8mKxavWYHh5++rOJNMzEKJWq8Ra/O4lutZd+U/hvYTZ2NQnm+xxk3
ygCLDqDnUGosei5rny7FyL5F79XxFnPXtnDN42cQ/aWtoqjtD2bYQC9OfEiuCOi8wM3lRIAF1QCW
JACo48y1jARA5yGjdPKLvAc2oPEn3MQvUMRDUzFB76EjGGRAEchp9BotdKnlu8r6+921z0rO/m8N
brnK3R4+sngqI3TWRzEDGvzXS5CsoRjaEsKG+lDYxlwjl6jmdtNCT9/g5gLW1EL0F60AvbJ+bFT9
qAqhPE3SZ3wE5g9c07reixP3zQeaw4hB/h6HuXHV0fndPGwmZSWOExoQNQtD0pzABdnu7fCFlWRj
zwf2jfbO/jtcJr5xoo9gvIgvVWkDwRwOWAV1N44ROawi/HkANm/BU6J1XVlXpUTyaAC33yAH+Ctj
gGCL315m5UdO/Go11ttic6mTgTL9mmIwFvL6Ke0G9AOJA4noH6D4d48PD0P/gncKghP2dt97uCwr
lwFx/8c01htuWMgSt5/pkPDigjq1yhno7h9GcsVyW2GgwfgW5yrTsUf1Z9TdrHNREGhJqOy97Hxw
4hGAtWrGcN5ZTjibbxCXKnTjlpC+bswQjlGVEkZ2AV2N2LHXnu/8nC22tXc+cGVAxypwsYFrAbA3
BXCDYGYzEgOYjw4gNS5JWBZZDR4G0nrvh1x7O7tl1/YMK2vQ4770gdbQng7izNJctgR+1faXuQ/2
5MfzOKryFWg/pKlvE28XGC2/aqHMIy/md6FOs7Bqg+9/rnpjJOurW4ENC2QRmVjCX64zLPyTFgE8
IA1rjqtlQKhSUS+KsvCWQ5Yt+rYx+Sc4Nf5x3Fe9cOT9IXuAMCYEM0GGClb9Ywvok8fSfm6h4U0t
2d4fKQzZhs/b5CTMf6l5+n/AtUoAW52p65GTe25VRlm51P9P7/nmZx5wu3g7Zq80ZjcldG9rT2dt
mWrLmrrHH6EyKQfKH4nzrHeMPkKSTDpzzayq++6BEW2U7+YGJ15N+Zg+PWF0FFfnOAKdlCCE74rb
KD8szrlMU89+ZTmsDkXGVJy8w8lJy60kB+Pw2tyK9g7muT4OQ38Reuq2NEyBoy0FKw7QM9rkbdPz
ZVvkul8itM55nge4ss8z+kUZF99tFLQa3RnMuznokq19I374t2VY9SBoKXI69jiLJA/g+j+a0pkG
jED9YBiPCNvTelzDl1Drk6yjsRw+KQZL76f9qaDYWsAvoS8pL9Z91rAWt2owr8DR5zTnWUD3MAay
uHuIpvomS87ku1gzjcwuiqZLpo4RGcAZJ3RAHgq87JrfzxItLBfGpOX164NIk8oYhp3IfIlzuo4c
B1bzZ1ct1lU+GYXQq0J9o+IARwLauObyvuA+t1SMeGurP8uwkLH4HQO0bda4kXVzWPxrTk8P+NNp
e0dho+0G+1d1yloI6waWC2EBiNaizxBCeiaufqE6jxwPVRR939JvjQ+MDKoJNQ+4WfRzHaTsP1JL
nnhiztG2V6EJCLM0YvFW5+HCHUXLSHRMoXbaFdDD4FSRFCHa68L5q/OvkYEaq+ZgB4QyyeayZNCn
Sr1oTlVAkEG/PoXjXThFGxALuEX2I4tK/7sfHtJYcpdAu+JsilX0WKy0p6QLdZtiVWxXdtHKojH5
LRLV37yzJRbRPYuLQFNkdJNveJjYLdQz7fYc5yudOY+H3/Vlhq4W8lO+2as8olzHBLfBKB/sVc9J
hFVO8W4uYNVHdADgrYiJjeunn9ujGBG5nmcqEjGcC/Fm+qxzs1YKPjW8XADTEpQ+Ezu2/3npOkN9
cawnU6ncoh4luZwOPz2mbaUQzsLH1epLNInB7rpYzo1WpvI7WUW086ne7b/faQQgKabIIfi66FXA
2i8eMOxY+gc8JhIqNOe4SXbCQpJxT32p3BTgOGEiBLN8vpiLnkbL4DUcVslCYkSELzjoZPCLBMnZ
lL38bPT/zGdUEvRAc3aUYfXIXGuAvhVpd+fDX3vDPaeU2gPaMsdyYHZsjtXdY6quHRmcTsAp2hg8
am+EyoZt7i6tDJxDEGVsoS3nFR+mABYnh1fcnVugRGnv4ID45FLU10VHHGL6B9IyTZqVK3Hl6Jnx
IjpVfJ2vA+BEyiuXqThiE8GrNUoRHz6I5TN2e3diWiNd6lbkXYJfH/tXgJ8EquUDtzQvf/UVQCbA
ZsaOFgUP0OJQ11Xfs9S5dp7m9RkAK/VJtVI/PyuUx3VAMmvKNLjnYohlUMKWFav89pt7359s9ALF
3FXK/usTkXbpQXPRffPufb1i+CGtKYA7I8N0FV9oYJqKhH/dPWmBzn7IJ3kGQOtR9Gm/vkvl9xME
a+7AakPjiUDERUdLmWrb8fLU3ZRoRqvVvBlmL2YDgqdwJI9CwBr9K32q6IWkoPBNh+iJtKKV1Je/
VU4cGWEDuhCuneZ8fio56k7BaQnj0rNOwmzqDbDoWPlxnTJOM4pq/O4pcrj56X+hzwf5sc+K6xIu
2DrcRAArgo3HAUR41vqsZrtARooT89mNCK2B4lBCbcYovNkjoGLOvBHsUcjJGFTRWqUSOjyuJrz/
S50NnLEX0lcFN+CE7WVdUuAvGkgaQCFGEYys55tT/RCThcGFrkjtZUuzHnhiAHI4mTkcrSrIw+Sb
EC0R0zS4ZJTbEsPbTtI5xcZQZNC6AenJqgDCwrTea+fwZ7K7EgEIImoERoMhMU6GSfO1/Ywql64f
DhTYlRDb+e8OGDg9v3JDJfDB/0+Gv1dn6W6qbFExmDcujHQUvsl2SNbmWbesEN1qetm29R7O0hln
8ypOBWyncdM153IiOV1yHWUDp+41k1IOd2UzMLYBOA8gRVcF9gdD0CNI+NNZR/8ZkgMX2CwxJYYU
SLVP2pV5YqH9VDq3KpzOBtqq87I4fMaqHn4VLlEoCGEBPUI0Gqmp7CLpn9Ng89f1uvpiMo08hF9m
ix3XX4qHSJNo2d2UHgN+E1HOAs0gPsyFbPh+25zcKmP2G+Z3tw6cIS+yVYkE61zRyfH14DLKY+ie
6QL54zapQMaJjWEKjGEdnDfmmoGC3HxXy93qMjCMMNpnyhqboqkYdSg96hY0eOWSPr/c72ETHIo/
Bqc8OwGXxN6C1+FCRDz7P+YdX94f8NY0JdGcQW+a68b/+jSktOzopZmL2hhDDLS13xBBoln+zqll
Gd9IzEU7rVE5C1PEdgPGM84kpv2owBPOgcxChS2rtNnAjM3ffUZUKXS8/c2Sj8uIiCw22H8ZsLI+
qQrgvvDpeEGtT3RgrXttjWTZyRmz2ZC0z/tF53T1AAk+1Mo2hXj196HUjRURh7MnMcYE8ZIymJmb
SsgOwv30e8an8+lMXYuj47RZsm04IZP6yb7yLO1LE6wYMr5SV55CXsG8amVOTAzULB2EgM8iENBy
AU19k7HLmekdxEzVGIkH0PkHGHZ7mDAjhrvgFxZmlPnssnCtv0VlCLYur6Gibd3U7OoarTxP/irZ
MOHUq9weC1m1FTro8dR0dGoyw1hTNG9AA5KTH3+1ta92CmBXCTy/CHDNYPdo0TKlyARYRS6R4xZE
5+UA02gCvXdXBRts1za0KORarmeGZelijtuctDbbAyB8H6C8eq3et5/kvPSbSHqOKIdPE/UyPVu4
96WwTY+8kSDHUL6f+5vETL2y4Lh4MImHuDPD+eCFK0WX11tzj6DzO4REiLQQdPoxoYFUe2fYWGD3
dZuU54u7HjeIfExC3OWcWc8qOERTBZ+FrhD4cGa+OgHMXJACPAzPIFyfqM9d2hHQcMwnyK8H2BN1
wUSfWUsMAPVYvNzHScY9yXm8szxGyhquiYp6KDECKzfA01Epywer/ocb+/d2bFAoQSZIJXSQ+/kJ
tyQ2jdcee7g6syZevARRkePYxLUO14k4NEQ2IqMDCVUr8jpk7IurSSRVNlc/CoaW7qDExqrE2Pv+
VzUTCafD4DDRz0eTHb30+gs70fkoywAs/HkOq4puRfyuqpd4WBRSsLI9mYEmFxJhp/T4jWqYklRZ
mkxpDwY8v4LrJW2WXYIVxOF4U5L96mXJiQV7pnO06yy7O4UxE2mPO47Yl6QinD97at7B4YhdDkXk
CoV5DXEa83KI3imcyAT2UNwajyv/cPUSspc43aHPm7EfAGAVTV5loNXmGvwcafuObzRr/fzv1pHY
Y0JY/awdVfzDSm9xkCS0T+BRcXHQZFQkiAJm/MbtpWUj1wSyF3C7Nrc0aknH5cL44DM/gQOhKNon
R8PKiGdcYsYBOa4+xjuQSYmM5sZcpCFYyNMERQ8rBW1InyveKm2Uh533J31STBSMVlhX7zpViLIo
zFazix7t+bbtov+NAQX29dTH2QKpUSxrS+0GMW+EZHOmd36nG0MfVZlUHtYkaIZ9JzoO0F22vexE
zoqIKDAh5YupPQGyI59vW3h4i361gTT2/WPIsfr6AfhAh2Q3IRyy9uQgkV1HTebX2YQJWRY4lx2+
Q3smo0cHLsbuW4EaOMNg3CecTXn9tt5U1geTcVVnnH2AtfYPH2LtzevO+G8/Yu6dzlSH2o5/W8eU
mpJojRf3N6pTqfhsyy7AzagPrBqwFiO6jAHCeT8Gtnz9qlWrsWP8KZed25igybziMRlBmWHrJT5E
BQxZNCqxFrVMYZBGkMmZsMcJbckBOXqShtd7XJdSDx944KSVcsUMZo8vf7zAkQo6yPFsPpMec2il
Ih7stLbVwMdZkMX7/7G/kG4R2/xDJker7KtL08yApTZGwvMuRzr46j0iH1QclGrdu9bclOKCS71m
VUlVYc+Q4uthhAHgaH02JMJ5LSfCvvlk1l//Sf4aQz8ZEGuM7iSHMvjPJ8EXZkJhhJoaXZPNomqp
NxSCoTBNHBeG6lUw5PeOE6Kj9VqYDAksJqbtoa7ADk/2CFSuhr29/1S4zqwjOdxVdObHggWYh9Zp
emPzNnYPMtnm1g/XRgbVHYIh21wkPF7/8SE5hptwA6+esilYm7ADvaVZ4J6QnNL59KStekvCQ2ZQ
1y6LYOtO8qRN8lGLgGZuv2YWBV8betY77K0vAr9ITi4eZcJGwlugM26s+epR9xg1NMeG5Aw+neJV
gQDBxcrKwUfbqphkfXnmtViHss8WZt1sYTVcLJmoVdudzxMwsPfwtnZD2yO9xAdLTQMYnDn8fe7O
ELJW0untKUl9xSVIxECn7m3NI6NF31DuiRV6SSoTOXPZNudoyfDP4t71qxSDP/o8nxclBs/9rOo9
JO9oa1Ibr66G9A/CCpVwc//Bbl907GqU+y1WGDRQDyGTmuTN8RZOyAEYAohjn5K9ZVvrTkPIRfAO
50iwouu8TFkcAS9+zb3fuXyokKl34m+CTyfaWRXYbOt4sMU2EJtrjbSgLZOhI0j9Cz2APly83w34
rZO6PUO1lKdAEKmNal7xcLufQOFN0q/0m1Uwjko65kkuXpBFBNCKYrQ6FgWa3mEfiftPhskNcjOx
dPeV2Xs8N++7Ou05m2dyn8cTW9VA8hmgsR+3a5jE/U7KzxL6hmwI01cdvRCqpD771E1Yx+KTcee4
Gr9ksZ6VNguH9BKwTrWc2pCmbSaxcRNqUMiLPiJvy5PPvIK/SGgD2AuWBhBSPtFAu+eEPCJXO4Lt
6cxwmEytSZYz1BTlbg8azc7tJsdIydrFQJzqkz4PoJSMlrQbwGrmcb7waMzAAVyCfnNT0+7EMLeK
nHpNxiZL75ypOm58RSzMC+J5KZI8BkjDI+zsb5aR/O4FLmJhesGxNmYVnEAi/jCZIwfVJMcPqfWx
fQmvZsQWj1R85SsDQYAsNb6krubNVb+E7biQFDUxf2YIxkkiE0h35jEuOSRPRTuI6CQb2HPEQjEm
4mC0WdOhtWo2S/aFLN5osqyP848beSbX5QuS2s5rgXYECNzfnG86b5JlGrzgWgemYZ3QjhnEJYVX
AhoIhIqKL9e4HYnDSwVpbIp3K0WxfLjb30NaP+1VoZU3pKAF1XIkP3ZDPBmexo2wmtv0g96bzJA6
uEufXGYbdxeycARss7uKCT2bG5hhkvh3hf0o0xlzwcLWbJoFTMkTkGHtBrIpJt/5FIm1KR9kkgsL
sbg+k19d4JAYMopM9xAESCORqO8qEEJY+uQoQ9Hl64lOY1C8+sp5bu1//1YxhK1KMqJu9DtjBCnn
n+cpOaCPuAx97o56vzS6kbzlYyq1VfGqav7B9G6EvNplCGaGr6WmYExp7gpvRD1Vgw53dv56DZ5r
FdlTN7yfo8AUEBh1RaaOn6GRf+YWfbh2t/5xm5KbDSw++GTOommuO5IfcCbNaK3rpN2XKOiaG/S8
1gxhmYsWMWmBnQT4k5sHsi8JmKpcFFFZZFKBZ0pUBU0Bhw0CXMbnA2gY/C8t/LlfKYTFE6/RfgTi
MmRIocGg8m2iSfJyY3MkmTuZTGrLHFb8sMpns8+XnG6ftldfqFSDaUP3kHrgr+21ay9UdEK/xoi6
TYTh5uVfoso/mHf8YX4XhuPW/FrHyOSQiCMGB24/KleYJNfIJD6Yhi0wnFQEnigo0NctgSxz7Foy
80vwze6kUQC6vgnmDeYmr/JBadyvbaUBHbI+HC2O3f2jnZgbKqOYAvBh06mCjWXlcVE6kCe2RyDJ
jSeNDUTkWHdUMXNWrY7bxV9gALGP9WTIm3vpXv/iLNVEfFtKUnIhzf7xhbuzEeSGObrm5lcmUDss
E/QMLDX4Pj/+ad0u0cEW1NsZ4lVDSH4JdPC9aeHJrAd8+q+b/0M8MwMDLucom2emhyVQBndMZv2k
Wmy09YEhMqKugPXJAgAujNN66af1W8s2lp2EqRn+8BkE1KqLe9kp/jVU6L6SMLajZuo1sL4D+W37
uR3sERYXg39gJdmkutbq0zzW2wozullR+4mLvHyZn6K7hmVn7dNIKMJLQROjQpfImSzdAApd617v
G3nhDfrkbiMDgad74i8bYxYRsWZzaEVk+ocbOC31iM0mONqK7VuZ2vb5NInA1tImA9BOZdNSmXJi
LROWqM7Mh/sDTwc9x61tunhH3J+c9DRURTZpmEqCfsk6vTEZTZ+9swkXDJcHOW+wFDbA61YdxJJy
1ZCNvr24eUlLIfWSgC4LIkaLQDtCykjw1olX2lECd7kFwkQGWdotktsJv+QemVGEi5xs/Fsdd/gv
YkX12hbAR4OPxTMlP5vVIdaof0tbMRmkmYKHIf8ARMdRwRky4WQVxPxfN4Jjr1E1aOF6U9VNzoz7
LMZI+vmGyxIdpRBMDaG0+63Vas7Z37bqs/iY/SXws83BzoQf+jsMFCBeOlHK1W9MJrZe/qzqsJbO
RSPHegb6eIPy5AnK7GC4LHXcPTCCWRxgeDXRCNo7HgQ83d2yFt7jc5auweIuCX1YZrmwiL/QFB3p
YteUu6cK+IiOIzQIXsHJ4zuubjjQ4BXNIRRCgH59WAUsv2EhxFqoKEd6rVQ++Q+IbBj16UIZ6fQR
+JA/CpsZfiCtBtSQyY4Ep46daHf17eEo0Rl/AgQWKYHZ2mdDAqESoloFY7tMIiJeA6T2AJnBNsi+
fJukN8SHVIN8nre7nnIrhfxk/YQUVu1X9a6s6cBDePOFwSgOlqN0vdY0IpUwfLGm3dxbxBM+vNGY
PQVyslDEl0wqskh7kAOpDFo5mMXAbOtI2mSvzQJYASvteGFL/h+Cwjqc8QhZHq7ZdkhgtNazH3xw
1mEJScm7Hd8KZOu28rX3xanYDS4B6xbqvSpk3UiJoQrCPVog5RmPO2alSf27oFhFiVES74iKvgjv
GpJ/A2FoIPVo/yNyTdrQ9kT9MytRLIowl0u06cDdRxbHAAkl24Esrt8r6erIdCqU/QqMFQ9zRjMH
AmYWzyB7V1oAXIpIYhTKU5S6fAScWC4UmqAGnt7YTQKgO6MW4xbpeXXyUSSO0QfzUG4r3ic1s2us
gL8qXC6tPSda1iOYO7VEfwrUcBu7IZ92KXgDtzgaJoURmZAAlutRq6+XnhlzGqpeW/rrUbbb9Cvn
gDBc3tesdfeChzOPnSlZHdy2eprN/AZ5ewnv+tk6tGkUeFU4IW+8JEfM5fr8C1f9LdtomjVXKGZ/
jJwiO571/aJ04lIUdyjrunuAxny55jnKNjZQ1tTs7LZUdkcZfjyl0KzGpm32d56Ju5asO03R1ifG
WYAwyrnyzOVaPL8pVIMNP7PqzCDSYY637/lMzQHq62KdzQj0rkqr82GBFhtrni+2lWn04C/hkGyI
YCFmiVZSg6JHS2Z8wIDe/XOZAnRx72/nNhN9WB4nEl7LpDA/KpRh1EiJAclX4xZ7yOCoNaguS8MK
q5uagR6d83DK3d5oTwlebmHBtpx1fqzIz4148Fv15soaYmjFsFfD+OcIOHfWF4jEs/WwryGKniRh
+S3GddBZof6fwB86/6LAtK/rBIDqNfXKa4dWPkEfI/+E6dlQOepOU0iNqPZi+hgDsEgNN9rCg2yM
MPM0m0G2NO95m6GiAbpylh49RvN8LjHj9BogppzYY0OhCttZ1DNQnY54yvcSuDio8/j/9i2lTZN0
HgiSUYAUQzDq5wDXGtjOUfPvosuOkolP1bpNOvUbFaTcIvPeAAd+BH6NRHz2fVFwweP+FAz/Ulwc
tU85BERDaTpi4C+OzvJ3JCpDErzsIxrOTHsbDrvLErFux5/Va8r1f5VKU+mAzth/ptyOEy01cYPb
RAwHmWMciPG999nrZYmM4kxFICvTk00gK7pdtIIN/91tbsYxIsAKgSHlXDCRaFZu6u41KKbva8+B
MhStE3NbuFGkAcdpIeFHjpLUpcUpL/i5YlZ+3qlcux9sJ6d0VY17Gqduvtnl50wUrEptBO6BaIHl
npiiCAG8erSTvAsQjbsSjzz0Y9haPFUEzELspQo/rbaFRyyisG0Q437F2h30N+1u1jgbGbPjkl/p
cb3tz3o+f0HPAzFPk+JGIBsIFZcqAKcK9SXLXKkXCrhLjF/PgAZbVNgJP6b0Bqz00NNiPrYb7VsD
Bxf1Mgb5Mec6fyAxlZMfBxmwdZDhFswyRAzrOM68efuhh75lNZFN3l2RpfSepBDCNMDmEkL3DXGW
1XrTxk6epm0erQQhCXTCuYxHRuML6YcabcmPwKlzh5NzK4zKsNlqYViXOaDgxZEiPXdf9tl5WTuF
YI8CSNU3pS3J3DSHYzN+BilXCLsnl5WFcKW3WSeBzhQ2q0ciztkM7tW8MWWchOyzcm1ezo/3SUJJ
/hi6F5/aJh3rb83LdyOBqFukPTyAYGwA7HfrNnTN/+tbiB19aM1OTNmSZf3nyRIXmKE1K0soUh0N
hiFZ1fx3OvElvuC8hFK8qcgkFTru4Mo9NPcRzbznIT+2w7nWvmKNKV/9oCTUmEV0j5su3R2qcm/b
ayVRGY30L53Vvp27F3A6cye9v5AN3t2NqbU6UGLN8nQyGlvga6M2fybtBV5wpYClbiFygayx7H2y
rB49xgExjYMPKmtVbNYvFHLlQIXRAYbrHn7SkbNY0A8QyJoIDshqTZr3iJL4KYG7dSexuZ1974uU
r6RMk0v5QjQCgVhBY7FmPxiXn02mcrfbrCDmm58zJrtHd7T8wDNPFyERa0dCAT83kJP1NCU5ERdf
6YqZthDlsgafFgaRiPo+zhOv/6aqryEj1H3MhdETamk3sQ3UPsK0G9jr9RTj0VBu0ItO/3FL4jRP
8iNUk6FBFyMd1Vs9dBSiVS+dvNc/nQxyPJ13A5iLE2hX0jDJDhGX6s1PKnAXeXyY2WcW3Xb3KSf3
wj1//wJQDEIn0ioUutJBiztv3fkXwAhjDGMvZIQlOx9uuvHOZ5Tai8O07VdzBYaQ++QBEpMtZZX0
3PBkHRWsKOj7YWIBBOrQtIUUfGq5fQuQqI8jwYdZyWiEGP3c1jbyUxBbGPP+tf0kJ3v5yEvWUOog
VIB2mXQ02a77HiTaufDIdSG3rwo1Hc2h4mnS5RPKfrjjXanXB3CU0B+kB0j/70iQ+JehDiViZCwZ
C+kunO5NAxeoTkbmAukzziQxFnT/oA4n3AGZDmE9qkOOAd5vI9DCUPz644KPhjkWvs6QKSiDGzX5
9RgLMYpptUmL40ClZX2YEKjf9umk5LN9ffrYJ+ZqCzrzqxoDVaNka0f97Zee71x/6BW3TNIBXvBn
QGzgCrkaMSERt6WWPpA0Z9PSg8YhAfJU3pN6bJkSO41CXQ+eIqsVHEtVHCaScGcZH2Ti5FMokZGl
AuHxx/pdVFYEwZS+NG4AlsZGDYlssoPzBvjhBDKNBmpbtN/M41U3gVcBKVmUEjS0809js8lGaITX
yDa5S9CpeX0iQalQIlWrYGNDSFs6Ico6zNmRkrlEqesf1QX2opnZBpNQOdFXSzeFFasTjCi2ENeE
cUiEZrHmT4SzrlWAW23xqw6K6V0v/Hn1gaaEnbQ9Zy64+rOpPYSj+IMGnJ9L5tC6zTcnS1VKhdwU
O0ZfeY+Ndw+XHCBXtcm9AKueAxUsSg93iWwfFmbTr8dH3aO4BL1YuZLKKtMoywuXbEWLYCvHGa0y
IeyJOqOjA72LjyyQxCp4naiEf1oBbPIyAB/mGtj9KcSmEN1ifgyktWPCEfYKKuiij/rv49fxxw1v
xu3MeriHRaOrepuItnBqQsxqemYSketsAauMyCFqQ2sGkTekMItH+gRl8BqKc06IRqGpAUXOQcfY
4h2WDr9p8c65nJVlZV26Xx3Fn2aeEeKYX9//6s2/i3TNo+OAgfaH/PemEPLswHfD8Zcf2DGWMwFf
5GvviFIGDg77kdPFmCRFFlhFBPzEdE4TjJCYMMBCGXfZ+64geWsweGk4TE9xqisIGWy50NxQhA8Y
FKguvxD8YYl2mxnQab13AdTMGvCdUh3wmWARVydn2e/QEZzVjzasPb5OM+RO4TIGi+RABb6Jbnbg
ICp/L8VIiSays4MEXFR1WQWJiNhlT0P/8K6DDhoIKrdcWL/5DmqU7fPkrHPLivTEBH33VxejgGrc
klyPqON5mRhytPdw+AYmakKsRZMydXizCJiuh4/Dh33DMss6AfAZ0EyAaKJZpkKw6ygTvwXvSQAj
ZRxhaaXOus5SHWBHIHm6GR9vJAwn9iLYrTrKBwKqraOVcNpUIe7ZoK7QPFV4m6nWnxJVw7vgpnHE
hx2t31+4TxqxNT/0e6l3M8VPGygUQu9CK4UHXf9t2oqx+9rFCayR652if8h7q/wjVTIpuenEiyo/
lI58lGKU2ravcsyVpbRyYdM4XGbHf9VdBjUrqvX2x4rdHS5zx1uX/4slF8DAfJ59H+98tJDw6iw2
s6kU1weATJ/+veL5uR9zYfXxmjs67PHe7K1EZuwvOD86GV/fIH8erNRSx7Gl7W7DHUu86EOFMckI
svoqjb0+oj7k0PCMrOs/qMMbeuqesUvQGjqW/jobDCAENcj17583+v/17mJHZbi35finsvLvzXQF
i/PhNPVGaucr1BQAyjNgpbz1Y/wHtxp/ehcDmbR1H3Eib55eJ38WM3RsldHdNUO4z0JVdtXImIKV
i/HgKwZj33T2Vn8rZIf4zqW47m9nqHGh5mp6Rl6Bu/F8QlfCA4e52jhj9FrRy05xprFLPBn5wuCn
NFHlk2Yeb4mUxwbLh7ZGPD9jE17P10UFMg/tlSOJ1L3lpJV0tIM/lLfKpNPgJKkWbJ5zi0ZT+m1Q
7iR6R080ypwG9WOS3DaZ0v7ScwBZ5mDKhu2cigvPd+jYBLyNhWf9+ofV6F0Y1tz60DyRvQVDxqAw
GDT46exkKj4mWjHZypmEF71WexGwyKbZ3/OkSTqWNERTl3f73Vr0nPyKjbdZUlYKIZYWJiq7nHIQ
Uw1moU7j2+CB+VV3Il7/uel7ZlcFoEqIXSHo8UOTXp/iURghIUMTMZnHIIsHgTbWRXhnNNaVx7lN
3rw74ze3EHlzldjg6jzQtpbdoTlLCE7mk9wGQoo0qmtbbiqNLTlmYqsrXlNPEqeqDyjkYujzxgMi
YtJWyWJV23UGBonmIk+gtngj03MfnF7jjJQoxYuoRrlPo8+UJDRZR0A8t5cCRaclvoAqGOtVX/zd
IUqfSS+YZbj4DWVEFsHCjIN3WM/eC6OtOf/jptAJ5+zieJEDYJOKjFkgedlnTfpVg0rXJ3BanipU
KSCCmxe7d84D0EDPrFKO+cXC2iADshl2a+WC1ISPBGvoBgXPy1YMw7Carbe8qq0LS5W8cHwCJ+HY
rFM9WDvGT34naOCDskZPjTlymX0MsEv1dyb2+9U4FRC+IRlycTp2KOFx/TqwcxR9iYAEnNbR4/kd
eZ6KQbwbLjQjg21tEdvP2/TIjpZ4zcyqRhl5qWkZop1FaFV5qdQPPaZ5l0wxiZsAQKt+4HCvXg3A
l2BTS8WER1DHk+/VGZgdekkFBOYa1+DyoyPFdVqihCnImf/VPA1JPYJ9rjxnTHsWgbGlxQi/nwlM
d+yMaj92HWuaCx4z0OKIrTRNRhAtVh0xMHEa+vL/JN7bwzMn/vD5ExGIwBnlBFZc3MNkoo7vnRIv
sxQzzFb8qrIPHFfGOka5+aLgcHjS5TROeZ3HSG0LiSKhmW9sjZrn43ygnXjBFvKTOPYQmdPIsHUW
jcj6/ZNfdZh2kQNR7Mj9Flu/j/eKCS8P9t+vFg+yIygTmK51thK3NaundyBMZ5mXOJVAU8RhHRyD
eNjNeQC8+l59MBY1tyh7Ltlw+EafzDOV0Xoky5UihPJ4BYq4RtG1zuO+fEs5kN20nPZEK1fW4/5V
NYMvIWnmBm9xhYQ6y/kpwqPxF3oXZ/146CYVVDfg1ZJG3MOBKdGHh0+BQWR0eZor23XSNe0I9T/x
8hMvtwzk5vgPFKxRTQiJno6+1p8ji73MGPJ5sMJVKCSA9+hAV3TGzo0j86MSwNgqBSUbh3a/G+Nq
iedelfIcmQsI/50oTF/0epYf7LifY0VMwvPKmZEis+IP2cSU4bdWH3JhKFgZ64DrwL1Q45Hlowm/
OnSU/VRmM3WK7GBLQOcntqtVUq41f8QcdzeHa5PELN3lQXDc+/M3PqYNR7XnTeo5DXqwtVcobIuR
nFarQrMp6N52GR3Ldte4aqJwyWneyje8lKhxkdxT8jBCFNK7c4tI+2zmdj2y+qZiSB/g5fPmyqId
UbQcTU2W3Q2ZPPhIJ5kwVPs1MTFwKCvvFS5VrO+5dhe3MWNDefMb0x644zOsRS2E38GJGJVpeQZF
wNXnsWCpBK9s7MULBB1LJx3ePudbMOtTWnNDWjVbS8nyCXLucLHEPcueayl2tlVDJhsGAJDwjtAZ
ghMfnL/JJch6vdafsmfwDSqO+UgPiH7CY4VH5nPDmJHYG8hXfZnnWTnrxwIWkf/ddCqCBbgTc3eQ
J2UaATqcqpaQZShA1dq7/4CVeGAx7gnPlNts7Cq8ppgt0pKrmtSZb9gvCbDZwIViF8xLb5odKCfN
Ar1Ia3OEcmGrH5jJqLebQYdqNtqiy6jU9qeZycJFCZWDP+d8pPioPXmwGnND4OUsbtBWb6Hzpucl
JC3SytP3qpWcbwieoDlNV0HcWlDe3Y9BjxOJhW7AVPxkt/d2zhjV52pncaH0RyvVGrUEzZZTFWDj
+ZXfOhgWRqzE9dEHb9sxLdTgJ9xpz4v8NHExRBbUCcSuDkrBQdM7VeT8J7AXFryo6XVnROwLUfjy
npBZJ9Egq7VCaZ942Mpm8uZg3kLf+QGBGsxl5Mjy1GJAnqZduzv9MEV+li1cAqRGaNIhQd5IXdpM
9xNdLzCkbLUAY7Vei+8lBbjEF9HxmSxAQI6eZwsQ2yzMf77bMAJcFyD7j+2p8rFgneCNvcjQUnEv
RWQ5jPTxQ/nTtqiGaKy3ibCdOmdJdG4oVUxiNT+N9ElwOMR9ZPyIbFEFSW48yq5SlkSApiZ9fMdi
XvqCDgQ+q0SSODJiWjQ3j5s6rQX3m20ONlBtfxRVCLBUnHkKmLFyKZusFy8U2px4LthQ1QxhshlC
WcyjVjfGIZebPNTMzu8QiuJdP2gEIyhGIh4ELNJMNh2qBUtg5c3B9/O/okCLWuluo/7MXV89DXZ5
y/2HTcvFWBcy8gB1nWAKrZVVIrKmmF+4ObofvHwugz/0fc0YBZ+1Z72qyZUm8hh4adYkQD3mmAV3
7Cu1j1ev4k8kv9dL7765XxvIV7TXlLgtSN63S2kITMoSs3NhjZeH27XoMhZkilB7FLlaJsNv5jjZ
pfXqE729eqzGVc/lh+hRlz7gYkQFhkSArAwDpiOu/W1rylgTbEeMevMm/RdpQeWk+aISu8rOLf3u
oDAVLNIUFuoGta+gWA0/o/Hvd1f4FnrAZk2rHVfnLBB+KnzdRX0wZLlLjSAw+YOiEsJLma3MrMqj
8QQU6FLHe/wOy6ZDDVNk/CkzEQxOWkXAw5gPsPQvWvuFBJafIN6c8/mv38gtizyrJyBrp6SjtlbO
mgU3bPnH8RWNAw4vSlzba82U5/4+JWpdK050/Vo4uyk6P9PIcY6G6BaeYJuyZzssNj2DC8QoEWmo
Si32yURoK8WKoZAQA4Q7iLJ7xngdP7DxVkv4dpQLBljSN7TIVOo+5HTqVTCTLxpN4ZVloPbd8fEB
SMG/0Wf2T6FVKdA6EfSjAa0EdkL/Hr3/rDlNWUE62eUs8W+5upB8Qd6DBvgvk/bLkkGvlrZ1DTWA
tcEIk2kr44+fKZb9XdGV8tcRmBk37LhLRJ7xn//qvvzfAfyNQ5LCgUZF+Z+3llpVOhXas4jOa3aj
ZXNfLruG0z0+fCaXAtUkQtLsp5IrVekr8rhlb4WEmvQssEQhvIgNHVveWx0xo8mk6kzCTMOFNOMT
RiGywTWbyrKb/ZT7yNx+RGtHeA3K3/B7SY8fOfycboS4mQrUUNvxP7DYiO4MnPxnq3I5B7GD0Ukt
NbJFgXbZJ18DLOsXihglUNEhn+GS3tfHd+4zlJDGfqJC3hbehv5MByz7VTJLNskeIxYqI2cgxWmA
677LrmG/1gJ/xWNkhyWXdjniZJM8LQjSNzFrmXe+QDqdlyIm28ZJhYC18WQHnf5IuzcQtCbW6LFO
wZnPp9fE4iaVCPyvZDD7JknOf7PRQrJpXEsA4P5+RSu7J7SNgB5U9lHtTnEykDI0QYp2uroYlfa6
6aa/44a0Ic3gOrXBeMp+BNG4laUdjUsRrVwQOcVKyfvVUxjDG9sjhXhICTrbdvyRqo5JSImY9XOC
G9o+wFUWuT7OdJQjFNePsEe72fguUkleE8nbRtkH1FAXU30751ngvFmochx1Sk13zX5M7fy4ya0W
I2t925pfjObWxafw4XVEYW20G/bswbcWrtLEoOClZnGhUQJU0RXVv+aND01r3XTfMzVm+6DydyQq
P+p8BMWLCupLfQoY1UtUhWd8QXmGu+sMmRUbV7foKy1SK/5EA5Mzq6wvRiScV+LlStGHp/VFuC8O
osGkwtH5hUlqyAQ2Q5mOEUmHLzoghY32Kglhj6oUWopkYozYfXubV0eWMmkAxC9PwZ2ndQCGxRaT
T5ellvo55GQOf4N+zWI93hpPWtan4Tlp97kZ+FFF/Uf+Od04S8wv7WvVJivCdD9s6Ujjbmzd4+n8
eTcnKd+Nfj3yHZpilL9FQ3ieBcwibv+bcxSIZWdmHpDhkfZyGHqsZAhjYvbxtEvT3aDEmzA8ss9a
YnT6KcfkZIV/DfbDyPbniKgq7Q25CDpbwQCoVzDgVhFL4g32vYfq6lKXYp5YsvOZCX4BenCNWjyM
Q6I90owcPMjYbSd51qzi3XAQeLCUOwF7iZxDR2z1XH2tBlJ3Ee241A98cqjlRm+/n2+BSN1WFY0w
6rHL/9p3VdPKBFyj4+iXx+alMW6QfppYF5LRAQDcWFLekrE7H1Zu8epj6Jd4qYOYtd3I0tnm/tQS
x65F8nD23RGl4uOqW1fmk7ugTraflX3kzC+YvjjAg/F1vUI1WwQpW0T+w5jQYwZfGw8qysb+dGkF
gAUyCjSRt0cBKm2L/+EKYAu20SzTy+squO1YD+dAGVirNQrJ8IgeqOZe/vROMoHj8R/5GYs3j2/2
IZve4uVtXgs1ndKBfVHZM6lkQtYH0wmWmh1+nWhIld5Elxx9du4paGMBdyjHbuuRHOgncGFW5TNk
0pIk11LNBz3VaLW9Lzm0+nkMhAlNmpBnuDmOlijhgbEdnmHBmNTc9Cc19P1LJ/XGs0Y7rdpAFRwb
o8irg70VerPBGlgMwajjFcf8eyexDoZv7hcajG8hAoSXs0gMy0S7zNi3bCdJZvzCcBZLMIq2Epzx
VROoKJ+bdAY7mRe/qSUJ7C007WbVF4Y6E8L2Swhg9QPOVksLcZtMN8I2QmEfUjNAvRYCn/3J4qra
xmga/ELBGxdfz1D+DJ1fy/5+HXms9fNNf6xx9euvOvchvNaoKahsUM/AFbbj4fKSKZD483PB8gEP
O9+J9uH94gdqusHAiUInFyaxWOABnYMdn2FadLF0nSrpGpcd/O/M/wJ/u08xfEPN7IhrJNVyta2g
+En92AlierFVgwP8s97YNavy/qGN85F2hZffQFlnHrRg8N8rn8St/oSnRORfVZkAgXCPWhicfKK8
mq3UVp5cFv3QBMbznNXJ4i3uWG6BF5Y7FOxlxEz3iwEdIopk8cd0iVOccRi568THE9/iKmozMPUP
2D5v6D0biEmVMIDKAM7Ex8SO8QKI5NDpBMsZb+CNYnfgavGg/xaNf+1NLtEZg7F3aSiGHbX2m6qC
cfFi2op9suyTlCbnPjU53s12xELH0TVRT/JH3rd/stawKIcY59jpLL9BqhrShZmAYccu8jZiaAnY
30jwkzr8mpWAGrTLFjojz6QHtBDQNbfVtLVisj9XKGnLZ8dzllZRZck9Wt3zaXiRq4iI2uAOkuXX
wf/lto10lAjosVaE1J4hBbIbZhNEdbRXRVAR4YRiMzPQU3z2xlBH9xd9LQ43WG7RZFdC5Fn/HyvQ
kecQUhJUQguHUvNxFTFIxtQedojOylHo6eI/lPeMxcrcpgacBhgHNawXX2JD2xos2mlSo4XZcWcf
Zl3yplflFwL/06EWROl14wYfBmA/5vfaezzCGSsgObzBXo+xIb1jTGC1WZ8ggS0v+5E4jc7bIyI3
XLqJIhLDHKFeH35K1lGu7DwbzJu/HeR28e9iL8DnWir4mMwdU9j2Tf+oNrwqCBvZGHRviW/lPoPn
SkKEjUqSJRVGotDOF6pd8zIcEKurnYYQe4G0IuGzJezMvvR5IlZTP5m/Wd8CKSCBQX0YE0p7yPql
HWsjyBfJmcRUU6yKV603PeflkUAR28XLjDlV6/qlwZu8+K5oQWEyAF7eyCk79FM76Boa/kY2Wvfh
GMFcg0oAJJiJQoL0aiw23CcCvsJRblAzQf2/x4Dhic4gwi4+WtiI6N5b4yqSFEg1UC5WKNpvabu9
uEaaTtSvmiQHQFIC9YlGcDCEkaMfgsLaXShTpleZP12Moy6qCjTgMlF6oIl++lsIvwwiNK7tijeS
0NF3exbeqebr9A0jT8DxOMBv4hLjQxguVJnCKxOsatLG/IXC4ncRQo3AuDNUV6b6dJbKqw8e3AMs
wWrMT+Um76tHmI6vOiZ6zsSbq5MMOA2FmelChPquoJXGoFjbK4TXjUQYyZC2wyyEVGX1xjXw84ab
hoXnbokhYI9rBlzCdsx9gNBgL8hxPWiGznZYZhGKWq/k1fiEktaPlf6kGbl3nqmzpTzIkOL1Za2M
4lJp/74v5n3s3+fMykMqQdby/6weNYPmY6PNO8j1y6RlS0pAr9az+z6HbArMcUG533uKQLmfF1eb
r+dVsmCYG5fMIfci4vZnzassrK2W6ooCT3bE6CsYJbcUD6ZmT/uCtmnppUhG0BpfMJsDP04Osqm1
oRbzdGKb8va0hpH0xYF6DFH03/WVBe1LaYSEQLQxdlcb/9cvfEGgLReaQaKjnkD+EJlhFyADA09L
H48yVpqlhfB8zGfdp8Illpj6FLaK7m+8weuoDf+Gf0G+iyTJGaHxB1KFNocrZoi3/HpNkoqV24hn
qZHg51HFlQAGv/2qvvqF2w2s28yv+S2wH33EPUMN9938NQgRRijuq718rz64w16+Qd6+d+hJDEwX
sQTQX+ffuPoOpHXvSY/MEiLNsnehg+o+6GeheuGxDWTPSWgxwmmod+w+Kjd2oyB/wH78BLj4agyJ
T3w4XnJRreiAeo4tpB+SI1dYFGsfe8AIj+/LQyJbs5/hMC7hPycUz8C1TKktPbnlWPpAJKnRdK1x
SRSkGWzuGbYOr8Iw/RUyM9y2a7EGkiWapcGuQhucOKKKl9TeOb46OC3LkyF8kanNsxPHld5Byaw2
CY47+gjeMBEHt8YUX2MaCqIRtXw9w9qYFW2M5HXK8I2DxMp0E8O3XDDDEakH6v6qPF6RVjbTizNO
5XhydYhrHz/DO9RFz9YOhDbQqyUT8CObOBXpLFySk5ZPEplH8w1haI72Y0slDo1r/tDePu0uyfkn
bLHYnjcVLSxwQ+fXF1VffpAZbw/w8w8szchvmoo9TnjwJoht2ziG4CBAetcX2KTL/db8l94yuTDj
nYG6DeMKycpMB+zauXYHyFgs25ZSu3XoP4VTnzKrxMB6cmpYt1qiEv9ZuQw5+f9IaWewELK7fLDo
siadNe1LF8g/PtSJdEv3qU9Up50uAMtJSNXuxzN3x5PSMzvFSyYorNKQ0Z4NQLQ3t7f08sKcp5pW
5mDTlhfOGb/r7CHatgGJnuOSgNoH3mBwI0pMUCD1/Z6wUim+BbGfjr62IZN6iSaCupa6derWb8cW
A5UbjbsrYn8oN00GJLOI6m3PIH4GJnFGSZYaXTdbgw4WDzwn94ZaVXNjpH2hjpaz/A7VVLRey8s3
5I+z9il+S80D664spjIfBGmWHN6+s4IXI5I3Y3tCIquQj0pdIO4XnnY8zLXlEwa1aapHzbckrArp
MonGefitQNk52sI4HbLKRiVKo6yK/PomxCELwVYnGqw/VBpJA2/oQxRT/fZ7qf4piwl7ZVHK3RZs
7cG0Ll9vKv96KLuS8fX+pAohcsaXHOz/qN8KesXh6+rdxOnAbhQ4pL45UvtZnFROfPPJ/qD6Vljr
QNktK1d+W5trEXFMcFVTV+8acbszZxb4tyXI45LiHs233Y363ougPJLQmpRVbvkb8kSmJ5Q3GaqD
9J5XfX0SGdnFaXfZlRrLRjfTwUn8DdGkintRJcmAL5Quja+5LP3qgBAIqXWMU7YPFGL+65VXJ9Zs
anvSJFKv7fmI+ASn4EVP8SI94a4BBexAYzTO5LuoJ3aD4hsNdaneS2pLPLDxUbibbUJEtN2gH0NB
Ma4UaB+BEnbaZ395IvlUXOGYypvYIV1WkipV2Y1T+a6ekY4IFlCWss730gOk7T0IQBRtNxrd+ADi
3myg2dLGEPIsLtZntn9SkitYPwOk2pHtteP1fNffdotsm/1uMb/Yupj5GxLzh3tYQyow13paMSs9
2BzTX1r0hDtwbG0ZqDSIWq0B1jJkkO98huITlGPsB+Vf1k0BR7nE3L3NB4ENSkQ8rQcakOM1lDw5
VYWMfIF7byKSy2Ws++o8rBmZLm/5Lb6JvtLgk/xanT5f2Eu7SB+g3OJto8vDCw77q/UxgU2kf3HF
xJPyg0QAKK8tg97nHKLcSxvhRV3A4Vug7NDJOwoywn2F0SqgZEG8hHXvwOw28ZQGjM5SB5A1KAYU
sLeGVaaVAPQ/EULxpTqKo4OSw/JkUw1ZOzebWlu/LesHV/5qS7xN6BdjdoBs+MKbB1uKL63I0OF5
g34DgFxH1gRhn5VP+OzSrbA6KrcrfZbuS8urmALxY0RdmWDUOW0hJfeHNfPpkPI43N5U+0hFrRcL
/UfCoQp9ZGE7W8C1nGvgD2gsslBw0lTPbsLeCuhmG8xDP2Vr6qjnJavka6hW81ig4i2xg/j18g/D
VUvt8DUFPDhld9pRmA7Bl0U2/GG1K+4Fe0EUmzb0Liz83TSectWoNRt7HQwFG7Ohn4R2Fq3u5i3/
u3iBdZ1L73fGpiqbjSgCjjcNgvjr/DWHzRB/E5B0w3f5lHBd7Qxrsy4coJvanq6anNlG1piens/n
tXxxKRCWWLT9x5jwmc0y9bH4q+1aTkm9qI8xc0H3ErTEOyZ2O46noGwnKoHGnQLoUFW843VEVWsN
IrZ5pXsuOsmu386IBA6mWy+uZSJglObrp96bEG/Hl/UuLy5Z+ZUj4Jik+EjjuYiCf5dpeQDc8sXa
OmIUv+Pb9ngnve1Ocsb388DAQ/YEkY4InARm6yjpx3Kkr4iom04K1GwfkN3N289qaRm8ygcaQMIm
IB0qdrJnZTcNSfdtLmeCYySpV7nWoWTmjuAN3EQvink/MKfbiEUt1lVItor88jwIWw0ynhfY2WF4
3YQ3RWXXWOR6zrmYggKxOp19Gcs8ak0y1Id2dWmtbpQrPS9oljVaIrO5Yfvse/dpig6a3Da1XrBC
RBaUBB4YIM/3U1oHUOaAXWSo2HtO5tEEi9M8BCXWW1Nu6+tTgZst+rAWar54L1SBBJSomtgni6gE
D67QuaE7iFP+6eU9/n7egSG+Z/KWnKcEAFd7GzRZ2zn7ay1LISfWrUGXt/ccYtcFRIEw5vCaSiX5
WShIQmPlr5sqiSOiErIIMgXHpY1GP9GRyQXEQSo8chxUZ+Ba3hGHh7gaXVLO0IXFl8YtxJ3IuAIP
EwxgAUMlcdTQUo4D5XZIkumgGMhPpTtXDkzLNGkEqfWDU+CAykcowR7bgSBrt0xxkHl2qD1dTVIV
/gexy+5JTEmADiuZpH6WB+wXQYgzt1zuaqQ4o/ic1coGRggm/2NosqkQjT1NksO5WgbERqTGWrS9
7/a0+JHdQ1X8jczlflzjbvoze1vTq4/FvzJxcopHWsOjQynG2yTqy6bVWsuQQc+fIcPx1861Kopd
+4ejrA1BIm6C6CdvdSTUdqGHok72pX15CC9bWv7mIaFAfBFkb8OAau1vmAvDxSsI+iriiylZzC8g
DYZmeUX1dNlHTq2VJZXOBBiMyi9uoImRu0INY80hX4J3DRwGPMP34wQ5Rst4EJzyduVzBNCRMSUP
DgIQlXJeTyDnIv+2tH+VyMHO4hWYoNV6tyhtiOZVuxVZhuS+ic5CpTOhgVWHAihgB/vCCRyQgrc+
SehtHQS8hvWc1x+NZH0CM4BPVOQ6CitWpMJyKj1KhG5mHQt//K5rgYEhPEdiO7MjkglqDgPTKuCb
m1RoeE8P+7KiVKj8aAJXGx6yznI4j2VsohHvXwoedeo77CZns5Ji9Fq0wF3QKalASepc6KO+tTYU
Le84ENMw9lP0H4v0uFMXyCPcNgaSzwytnfUenwKFSDH677y0TDb1tm3/amHvHS6Fxnhr8z/JBRRJ
2mPGMrLtLzdPB+AZRgoSne3136CaSw5DNr5kcPzSaf8Dq4MxirE6SsnAS0hcYqeSNsSk87ImWUcb
TYyTgwN4813D9kCwln/aPrPlpPflrX6qGMqROBtPGgQaCqcw3bIR3IwoM0bWx2R7Cz8jcQyBIBcA
QlVMO5OvIiWuR+C1TTvKTuu5wUtUl0MObdNhKDlq4bqY79dv73fivotieGPcKEOKZNQMSAIP7KgB
x23Pi/aq+dg58WUrWK+smlZEmUv0xDNzxVp+FmQL14gNtz3U84lXhU8mndFuePcXfKQhQe9dHyg9
LqJ0s0FS8c60cgUkZUD+WxXGs8H/HXcPNcgQmxzwPIgE4xYq1CnXn8Ahn5m5Z+bZ7+Iyz989KdjL
G77//bsCfbkLyfHEYXS8+6QGogdjqYNItCguRG/RACypSySBnyXzDbYNr9A8QxDZRxXJXYUTqgHx
WiHPwrw+taD16D8DrybTYomFRnhh5cMAXsR4+LnRXjP0uaagDqbzk37yaNGE0kOPkpqyCmhaA3ee
wYZ19i5bFXhIv7+yeEwnLnzvkYVKKCNKMtu2nUkF5SQkAJ+LlFrwCVvWMv8JA0MC/6Vel2W4zIgq
1WCSY+r/laSGDVyWgQFfosc7iOjsKzdBxFoX8ABaAbp+zlI2vmY5Nv2xD/gxYq7KdO+LVbCiVn+D
Vk4CQCtyWhS85cspZi4bIoEDiulq3g9dnM8u5vm661oYO0CoYGXGED1vfD1mNiQnO4QNMYcAtMS8
P5gRDsuq73GTAg1mdz57/vycRnABXwTxUHUM5TBwCfSItC6VapN2s21et9ndfSVLlOG8TsI+RRFm
NyLNEQYhbwJtz1VXniBopiiqrBE0pVZ/6p6E3bh2Dkplhl0RQ17n5MY7HAK5SnCqXCyupU3h9xuj
JQKpYZ1aEldT3Wgv1dwNOofGbv8Dlgb3I+unTtXa2T/y0ZbwXJX58y8d3zYFhBubbGZrkpj77kBZ
ECMX1MzwLnP7EiIUsHIs/s2peP/BeTNB1sOVzd9+DHMOvgESd29/Da75cZs8fHUu7nnE5ltUNWMy
2gSAZX1mLbfaf3+hEvD1JBvZ0ZVzUmIRbGIy6GphMtDJybteuCPdg43uarIMIGr4UqNofZtEv+Cw
yypk3PtuJL0bTBwID4Vybk65MGyIlJHFQu6b7v9Tx66cCeV2r06DmT2LyYTLU8uCzDickqOEXrjd
0sKgiMhXl57jM6wOHMLspQJ0ykixoclwToIxAh96ArZmEPEbkfxumoAl5pOYBPdYa4BZq4K3L7eZ
pbaEb7IxTK9SOngAFyM9QtM1jliWdCFDhOBID9YlbxOsPyOu6jR3tIg4M88YqKsyQ84q1NeqX+9s
ozqH8d9Su6B/au8OJU3bk4KcMq9686PbjNc/vg+sYwXnctigF2YWt0B2dMReeAjLgfKoOtmIwSSz
ODLiZPO00SSEcxnOad26hLUSJzqJTYc1KL1EZGpexig/ypxQjtWiUo56qCZ/Ym2B4TOaui+kNbyq
Kqt19jOcvNggBsDnz180uYhirw1g16HQPPdPu9UYFtNHWhh/B2If/QFP8IsCL7NW8vThc6Q44cdD
3DY2SBpHPw5IbAh6FKr6wPMGlWDjvFli8O/XjgmGYC9upSAuHXmENzF2eCh32ELCQtnXumcb/fhK
OnliNdL4fSABe2FoPosKnKquX/xADGZ5Ig+HKsXDCmZCVZzQf59IUnzALZmb0e/idyvuF34GVNNb
r3Gxdk2G+A0rBdU540kWFwxrWCddxDgwKOpexUtisKSGun0M9KZOGvheVWD2qYLcKwV4Nb+hk85T
MV+oMTadYnSkBRwOjR1jqzUmMVGZMlemWjygFSHIlyFT7PNY8BKCbOmnh/fi8G4OQrI3sHXfxVjL
t6lGtbs6h2aDdsAOgFGxbWa4S5moWfz+kNw3dRlhJeR+U+tSaXUmaFhYm2WqTV2rlqJqEee20G3e
6FDUnYBL5NiNSyNVlYK1bNmJE3MdkG0FV2M0/uyHBUYgizX4cXYoXLb7H2uMEAsHUQtDcOAnBlcX
xKBDlYvBGPKFSQ3l9AHDf2i5Q1K6pEpRh8HvB9SJRrzaWLaHuXP6ZZY/1xP2xO7rN83ZZQVgPoVs
LKOD0n2lCC3WE5g0LUwvRPtnIuJPiuOg3nUwivuKn+hsEHogHd3fhRpwhTyTleJ4/qDYT7PKKYQv
mgaDdGK4o5NnTsE/46tru4z/+1FB5GlFpwtQVeSJSEir93wI2jimQA+NH4qScA8+VBdAubzoZIGV
cSUFZpcj4wsnxPUXE+aGzUYv/QPGAAiWQ5t5XX9Q3hY/0oTU/KD6k/fbCOh1HQ2agLD8hSkOfwPY
XTY4nhpMdF3tbYVokeueiTmabCN4rMRXZ4/opfcAAsHSkRt9npg/AwKuYa6lnsdLxMaNXSc9ktac
X0iW+TWUddadcyhDZJP8fzOqp/YTNClGqtgmiB+vyvqknR4A8EtCoaJ/5JjI6r5X302YrDIQggf6
WfZuk9MOyVwvvmM5TQHpqAg3fefJ9whJE0HcMFwel30/82g3aCbRfVIue8VWff8tZ00e4pcIVA4R
qdRSnFr5rUM9Ng+E8DeXpGHSRLwujQGL8edHC34r9dsWfIYe+g6ycaAIk1cug7stGWoyVBrPcSdh
dLILB9bdq9rTyTAGTU25ikAbS9NXV4T1zkZLspo2XCdhqx2mtLGdh/pxgFtB06GGQo5uIs0LS05L
S47KRQ8fGp5hrpjXUlpr97CQ7sKxwuH//S4tZC7ExAhSngSb4w5LAtAPw11OpwW5dd6rdgmWLviu
IR7zB5k1arzIj40YQvWPzb0bjHqF0ZXyDUp6j66PHsLpBwgxLVuqikYmj631B7buuq5Wv0K+ApFJ
UqBIoFbJQxBE8fcarC6T6NK7PmzNdM/8yIzCmWlDgQKnFx8qILX1PQU+8evWKCvYalYJm7tN5zTA
5dXMpuR1zgw4w8l1hlQNtVRC8475zHWL9NsQ/VMpT1L9lKsDyzLZ29lMWmVB707V4xAPZ0vhGvEl
5tksBvqanJRg3OMdqqViNgUej4TwUiZJGJhzVwAItEgA6KDay8Zam2QVnNDdUG+9cWRG1oC19Hyv
ILscL8NbxQe8el+33a9ebKIilDaAmDZNlyIH8RxNDz0Vlvq7s8J6Ht/CHtzWuokJDqJNKuzS/0BZ
044C+yA1aOV2ft5Y6ul1euEHIcoCEwYL5m2WVtGv5EYkqPeLXvXlMwqM3xnAz8xNKuND9mk6sXSq
AefQwwwc2Z5JUSqAcOX2fZeDuKsFmq9Q/zt7BhJxTH1WrwNM3hloddMKaEwFH9LN0mHbHS4cONkJ
/TKFWWEG52pfbrT/yC/1xFkQxF3ycDBnmPCYwt3w4ddW65/0aYVr7FiIe6yybTSglGUzU/H73tko
dwp2uRqgFR2/pyFsiAxloI0yNhp1IaUEtQZxJX9J4n3NZYkNRmvvL70qGuM1J4PwrzA/BX3vF63q
V9mSsnGeDid/6gWyk85E8pV96P4K6G1NXChbSHVUOkrkX4+YiMTzY0RcaB+zBkxB27x5ych85ZkE
wl+ycc127Lm9UVjS4HinyLFGhIXA+cgZ5dkGC/IGSrgg/qcoWJAMsYlLnPoxU7lX9GBmfjvektuQ
O72hKfwggq9zjUL2R6J3MgHVv4KZhANOGStf3RN4mgWO9jOfjwh0vJ9gbKo0rzZCzi4TKqzPiIGm
CI7WqxfHbHmKG5eh1vBNopf6hDo4DhK26qubkvK9js9EvxS5ux8x54K6sAQzDcGAsKJtK89srQm/
YoneV/kV2n2cANkXISdNFEC3hMLXPzLprMnzqSLR4MeHX7RAb/TM4i3wEJrX5rNwP+dbvykz2sbM
DdzoD0AsBmJJiIB261MPXwRU92loJy3VW8uWBmhPyckTO504RBd1fS1c7m3SYP+vxfkJPyCKtxfX
kK/+5ro8F/FtOzIC1q8WxsMVZTJnpwcGTUHzqw6gCPF3i2Oxe4hruXWk/jcEsib9B5opcMqOyLZR
e+q/9cZYLBsDPZ6WPFcbHIUJIoKgZbc712ZkPb5EhcNiUYwRfH5GJ0xAOzRzoXs/WgcU2gZ9DvwN
f/BmxqiD7gLCQGGD0aoaVa/RS7Jq3wrIfuPRsb/8x3RGUGp1RVYM3XViHSJev2IJy2RAUvicg3t2
lVWOgl3ZpPwM8u76lZ8UecJTaiwkluuIKTY6StjKZRsKv/RfKrb7tSUlGXaBdXpACQ/wjLXdtRJo
fgKaJ2mTLCepe5ntv+2l14aBnzycIrZHNfIgDOzACz5CB9C4RVEWT3Lb2HWpffwU/HIUod20ms7i
MZjbjdBx35qSFmSvFmGHCqP0/qucIBdyPTeGOVG1D+qv+my7sSYx7cL5XGJxqAAiYsZuAH8NUoVQ
8ve3kQdymCzLRsFVg7TEyBd7bm486s+pGoXUoZ42mWqPInN5wfTPwNv25NUgTooqq88ujXyGcTqU
Xs1VLv1It8HY7r8PMG8S2tzGdeVpeDa3Ul9BwGrTL8oKPOwK0gXmiQgfce8FZyddLTuo9VsHaNx8
zqHVklJ28RSezx0As1TJ+QlgIqdFh0lpNEVaBEi7IJck4b76j3H+YdA2yAX79B5sWEXolrXrDq5r
/f2lXBnYj853r5iSWivI0aPU4xPA9wI+b9IbX8v6iIpjl5BWw5oHYlU4GF3OI2nFlHQbXRepv5aU
l0XpupOD3jDS3hSstSVjXAza+ZXc6J2hoYclO8M9AleNpKJsTTe6m9ftnXxaYsY9jE/SqE9MKvUs
B6s6ERGI57ubU/TEWlUo2svLxVi0d7hreVUkRDz2e2Bw/PDg+P1dTnh9kvye7tBKdyajnUbEU5Q9
NLTU60qBIytFKrT3AQq1WiNQcu7M7jlEAzXFq3q2eS6tH+EkrK8p814P3NwCix3CxtV6mQqqL3wI
l6mggnLS/n/RYpf+MmJG7msp3brxeBpMGWG5biqA/JIuswd/ItUclPdDM9UBK90jL6/ouiGE3eEC
hbk0uS7z7VpHax0Ko3DkfbzPDYzdZEzkHG67KAzJRBpEofYq6iPFFh50ZlTv9g5TBGGcRrSZLd1x
gcRG7ggvwVvfMbdZIGGZT7PXUQY7Eog+oHY7H+/jMyX/f5An+hE1EVYIW8mgqiheBEQx+m2iaNdS
/SLtd8ySHvylxEqp6BNuJmLuc1fvYRdLgzOQ5ccI2fwvRHztQ/jg2uiOZBJ6GSA+7MQbLcj7RNzt
4LGU/NTqS8K/AtrTqpAJxpf3Nz3P0v5kXxW8seK5uKwO63kHl3YtZeOpochc8/xJgovoMCKrlGIk
PXXNMSKLMCuL0RbNK2U9MgzFW0dv23GapZhAHmaDVQtm0h0CaG7SHZw6q8ZANOu9NrBMulbng+P3
3cdRB5TFqZxIA38yK6rc0zlD2rbpM9S2r+AWwpjc++/01xfP1lhnPpowQROBXIZYqwfj1b32hx6O
dIeiQoMf8U97nUmkhX/VtKYnbAHiFisWlMR6E1SUyrv6dvMnQ9vcIssLoxXtbmQy1eId/UP9EsSA
GIrc7eYmjFaz4Xa/XEKfVvalu8Dn6EMXhf/cgAQXeMeqblNB4ZlXA6wkPPJstYKU4oCYtE4z6KrP
0S2Ql/tVVDr5SI1J/edXbc78xwQ7aPjcgj1sgYm9OznlyGggJs3tQ8AXOz0N5uz3LiZxCRMHNyBi
vdC9jIw6TL83ZTp+DRJ6icM+ocpGmM4V0MgKzh70UgPkCnLaAVfRvlrDzb+yYzX5MqYM2LCqfBcy
lSwr3kPIN+kCC66yQGxwhi0lllT1UqDjiNnX0Pr0OQxLio8wXMkwcIKkxp2Pej5IId+OqP7G9Pfc
/YBlmg5OENuDaR62afLY7ncx9SnCYCl0gTx0f05GJXeNxyTrQMi+3GUZCpL+Zz8hoPq1tzwzb69h
SJ0LN35NGY2QptcKZjr83xPUmeaCKGpWmRfmXWde88btw/loJGyBvJi4PjWFd8rMWXJ1OnaZ9Psr
q1cKuf7j3KPN1u5eGC97YIlSK9MYTD9tj1YyPw7+otbUMukpww3AYbSCa4uoxXg/lMFI4/4Y7DaH
zsrH4QPU7lUEXV3HSSkGi/Q14ICRh/Px6DejzZPwYTQW+yvTEBrijrs4AaXyDYOWaMINaSsA2LSZ
OuoGq1ODyWtqP1mgXIlRe/J1PjHMP5hkly1w/62JZCCuTSEXM4F13DIVip8CiUtHjbXrcuPDzToe
smcMN79n7kfpBDCmUm+lxzR2qywumRJEgZcxBJ5zMZ1jWQQ2wOXSR/FqqAD40gxUAjjsCVRIw4Oe
Y5Cjz2VKX/XFh4FhZOFNj+HNHbbDc7XCmNSULgMKDfsjY5ZMn8xhu6tKfSA5UvCZU1HhrZ0aDMyf
89IZVhX1abmhD9amiBWy4RHTqmx8gu66Cj4G48xNfBBR0GAREN9Kp/dh4an4L5CkJiGDCia73yNN
OPXXJKBnVKSOoOlQNzMoeBBO8uMOTSfOMGYD8KobXWIGzop/1kicZSppYzIFbkq7iUdzmNUqXAPb
KGVCtjNqg+KFFWY4DVvnsinfQKLrKPKLiIQsAlbVJsjSRAKpUUQ0YXeHQLMYHok0S+9zIjsdlCQd
DUs0JvVyS8JHC+wlA/GVwc4uO1g8UqH11/DkF32jyrK+pa/PKDXZ5eSnJkfYPMypT0SSq0XXfzOl
w8u1rtridpQIo3XnLAfWaStrlFmcFCP/ZcYpl8sucCtAVlLaL5bIyKFQDSwrTwW96b0O3hBe7ORM
67CrKtZXMw2zc/b6bxyXdW1O6nozZ4Ovni+802o6g06bIQUyzUDh80hRe6uwAufzBx4SHJk0FkVb
SzMV9/5LMOXK3jOQFTcz0QvWZsKvOia5rYUGzBoEyob6YypFy5dWJThvIZBWpjmodEZV+yVEvVwP
8/NsRtuTObx8tH2PsnaQxXHq70bpk1LBAP6UepLaPOrceVz/qRlW1CvqB4I1sKlsogn5xRM6vM96
dMCYLQQqP3kVNGWa7J8/YD7BVtZ7IGwZaJlWt9xlRbBExKWnJj6k67kYlyMlH9XLf/ZtYoc7exND
J3T2PuQLxJsb/ou3I4p8pzEtwhsgl1EkR/hv5FFEq/mEoTLtkOYVmB9WpJX9xmeGFf2BTXOJaCoj
FjhgL34Whnpw+HddhTHbwG40ZNk/Z4jNa0NYnHgR4Av68Y52KDqO0kiD2l+8IKLdjHZWC+kjA5IM
EwA3fovZ9ZDjpPgzgcV0hxt2mxZ/+2xqDPL+xQmIAWWIEb0YLn/oNkflw8TwZrM6MnEygbhszGTI
DftUpFIgADoduBQnuhF0QBCC5KdM5Blvn8wTOH0/Wrh/I5of4aV9LtnoBJUU8uwuHDSDlU0TYsFQ
vin6AA13exdVuUk+qHMP8wPQ4ZMkiPCW3yMgqYp/EeHD2LHt6uvjQt1FG0o/KTyp1ypBYNblm8xm
TmKvvfZt2RU5vQneXPjTjDndgNnrVusgxXs8F+sjMvhzx3JF9cN2sO7yPHoq4oT7rnTblIkzI1T3
YK1eB4zPHlRendFalHKqbU2y8K0lajZjx9NFlqBmA6J9ODePiX1Abgr9GJ2VK2GB2TcdYVMAzCYG
4vX7tkhA4GONiciQ1/8cVz91Z7C/Q7ZYzzavLAiWDyA6Bur0bvIzg5oMmOKTYUX+KlXTe4RJzcmC
arMbiq98bHjhMm5qNo+/jznIo8g+H1PYTA0qpDttfnFPzeqvkSGkEkUCHgwblIQtOh7/PjbT3hCu
/2S/HR4TwaF9oaPckdgr2tmYII7C5OinRQOMUGbiIYX8Qclf/NCvtCA1ApnaZ8X121bPC7qCjX8+
+GfKO+VeMySqWdKAwwLMCew2q/j68Myz/e+Wt0twdvGro1Qq+vogRr4Q2x1LpVAw3irsyBAxVL8y
RGp4EkCq2RWvz3AlwNNJVwhQjoMxNrBlUfYV0mHWOEjzW2V3sG1K1xPxTAVz9VdCPIV2D4QS+ndP
NcBy+x8qQT5TV/pjilgkxY1/SdWiZQQcgiBgbkfz1hmFYXaeO/ge5Mie6fGpoUguZ8SzOUqNFkH3
Yoj9KED3PlFgqxVc/fEWobPYRCf0FDcq7zlZKieHZgq3TVKY4pFHdeQNTPdv04/dWq858C3+qfu3
mBQErcyIoV1zRNRsB32X5Z/Wo/tE0QKOrqEwDMwiJwuZJv9S/VQCNw5IY9+0Cxe0RzvTw9hPkU2T
hMBPcConmfCbrYchNDMKcWqcMOCBNDCXLhHjd6QlhmJct4wCnQOZKM/2VpEHGqBc4JNuW9BtaRsQ
JGP4mt4DEhEza9YeNiP5rz/Upj2ererEv+J7R+0/wpSAqdTqMxDbLhiaLlmbTCU5qdqncHFdMCrE
BfmzFbTWQSxFGp2sMD53FwJVIzSa/b3zhTVyDzyDC7pOEZNdCJSCCBESK1cEJG4dxaOFBDdT3o40
Bv7TguTe+XPHH2DLJpKeN5GVsxIG4h31YecuYN6RFTaWtePY/PisawEWMME9HrnUs3Spf4UUw1eP
nS0v4xQNZ5u/keQ0HdHDNYt+efGgXaMulT7p+vEPLrgvGyFLcA/vz4UHjdECKZUfqGXux1GTtLnA
b5exL/uh5tlbPGj00HY6VZ2rbnKb+swASLgGu+81trKGxedSzc9vHE2YMsZrkM7vC/LUswcS9Rch
/7rl0pPMKxTI0d/sXkkwxYINKAFBhdeZ/eaGsJS76a1aE1ZnA4YQnJwAS6YqeUgKaQypfnSdhIpi
Q5SRCh+D4SIDAPaHfhoth/RnrdePN12r96VMDd6KIs6jBFRX1IGPkAx/t2AT4+438BBmJHcWRRh9
U8GkaB2cgV4dS7vZo268b9eozGSq5MQEtU62mWU/1qqHfJVtY4MgNxrH32VflQJFD2lv7/ThNCMv
p1uXi0Yv4ByeOLsKWBE0WxD2OqLgxUzWAIUHCVVaPEpYm+4e+NElRjcVuvZxP+TSkywH9LTjvjEc
gy7YC9qApOYwkMkRXqcwCntPOoc5Bi5Thnewx3agYJMaFdq0Ess0sGWrfgxATk84JOD1kjn1F3Pm
EqLhxic9alz0E7+rshF0sC3U8aCc2mc8i9VmPSnxyKnXwD0zu/N+sYzWlGI7hyaBXeksH4a8m/Xx
DwHuYh/vfbtijkmwgInonZUqw3sIsv1VoQXonTgiGNexAYzQB5buVwJJzOv4x7UZLkN2oJqXHhd7
y9xoNF9e8iGRjrmIzB22On72zyfDSMRBsDsPbzOSDYP8HYbqQij+xwYyzI3TvyykreBQiAqPeAwQ
l/LgHTuT+ZVFbL8EgsN2w4OuU6z3Mg1YNq/KztF+R83l7uzqmF76MVoMTPrbZUVqIyMRbA4GfgWP
YJfmzOgGocVNuwcWZwCubbx4dBJAvbqm1BJtdqmIoNWu0jq4jmXxweUTSjX3jbAW+WMx3xDKtmyo
j1bvDW9FndVXd49AmiTEA9ngnBtPF6g4eANeTSY/I1x14tmcdKQPlgB4l54TG3xAWHgPNhlkMWMe
tFH8WzZ5Xi857o8NRf8LVWorm1oDIrU/Z2tBgEqsP51zBi/sC4kR+pmj9TDaVUzKQLKojxIIMFPD
a+uP0VKN+uW14YfMt2Uj6UQiPHg7uyrNkOFw4A7GBTuPiGcaDwVKcVQ9isH9w49ha6SC7WCHT68M
JEYW7YAF6UbFg89Jqrqm3ynvxvM/k2UAOeHC3J2JJBH1anzW728/todFBn7AaMnhpg/Lje0wxJHF
f9mXuNXgOJO9scpZJgBzPwNB6A5xjT9Upp8klKj+N2oTgWi9XULX72aurYXCywjdr4acLcPsHQ8z
Ak6kWMWq8ISMgaX/uhVNHJVQSZ51mskAT3XoiOE2anBAZAi06QYtwYKQU4AMxXyh1JcEfcym/kbX
JNFn0Sde9kYTlxkwMjRRXGN4KdICRwEiWejh6cBxvIVhWr4ukUFNa6uXltBIkPj7+/T32gqsisnJ
fVeNajFyXiCtS2rLYh0YM9TSKOBlrj3fEOnI/pc0cPfIh57/N8uz7mWVEQsJpmd5PwrBAniz0jcH
6c6L7PIrwnFpjo9PgvwxnfLw4G1QvelvweeUfEC9OWddTECVarmkFMut6aKLrJmkvFL4pkt2W8Ne
8KZEU33pzlAVSYoSP108OcSe6cx8QI6ZfzbOCW6EP8aM3YgeCM9ENzlmjANpmDLBPEwn4Aw7J9m/
9EAtub0GgzoocGtDMFFzNIe15ejWOBXqddnfPVyA5F2pxdt36CMC2zQu9O1vfnOb7if2ZmdsuZfn
7uaYnWL3+v3VwoH6o5dD4Sa6SQM04QHYjJ/XZNWLpGOztHUk+1bYxYA/aMedn6DaBXVvohwjS3az
grnBbswNItVUQ37XTT/STqLV/HMs0CpkRUUNpdCUmxazXEtgHZo5G5EZPNUAtdycc1B+z3E2LIvr
absWWs6RMTRK0D26wurBllewnR9XZ6AzP1uZGw/TMEYPB4SaKn9fGnE6qeLjiCLVIMCVlzSB+UlW
tt/IEV1Onxi0qU0gs/8EzCC3l33nuwgHjm2THTNzyiIHE/kwJ/kFmVIb2u/lyJ8L+EJwXE62YBxr
idOMh3hbZ7o0J+uxGGU7DFX5ILo+3+DA0ZhRTlaQkiO4HlaMY2JXg23c7HfxTJAt/0iCeYYXrm9K
5L1p6VDUBoCbvefmlvMX8QWUJvBgN7fk/KcwY284tcwCP5q/Jud/vgfFR2fzcnXsnbV8xGGTaLbq
9/bmbKNe6m5jzz2FxdmcuJQDbfTb+w5jfbEpQyXtkDxDnzvOlR1QuEeNR0j/4XCx8HHVpgQJdQx/
8WD7KmSIdG9WJON4XOxOx+4nqbrTapDbvjgkr5TSko5JNr/6rw9H+97MhX4hmbPwRIWcGC1R14CW
xnbu8ZPHyZxTZ64odbZR/6TM4Hmzm+V1Maw/d8pezmRwzp65yY2znSltHFYvO/hStJlkvK7aVgVx
CFGf3wllKAmhpMArbueRc4/qexOzQLwzjF0u3i4kiSTrZpVSNZoAVloYj7OzuNjWBRxkXcn0Y1xp
P/uKpACobT3b8bD4g1cwQMov6fLAG7C66Qas+LJbGZCvz7XzddS1wUNFuj0aEVRx6FiAFZ6JJoB+
YJ4WTo+GpoqEJ7xlqdXIy93CHmKP+8Z34OGHBXTpH00kLJtr8RHO6/7BCj4X0BQHuqGjryP5HDyq
JmcCUeocLqJc3PiTgHvusg5VMkrIaq0aYolYfTWy5S6nw7TejN3NvC6SY1JXQSG8L4tVvXxnuVw0
HjDJiE4v0t+Ei9/2mxciNCJqHrYLevlkAq1n04b3+XNwVO3O2y4r+JTNMTyJa7Pc8S34aUppxJvr
e21WGA7e9+rdbc6IGlP/lTKzoIm1hLCcUrf7GcFpp6x9Jgrl1Da7IRDT3thyRwgEyVWnzRVElhly
PMGkfpcqJMelH/rfhUEXt14RGTrINd4Ci8ubGF3/TPuJcGLRd99dEB02cI2kDwHjnOt73cWawvV/
crQL/xeOEfVT4ZrLg8tmAxkxeg3Afuq02HSIIKYpHKgLbJD2IIpTt7SfJhLGHXm4MruY0td+5u9k
PUy+UQddO9EZRYyd7MQ7LTv0J9HO7alxfdWC8J3JW54G7UUua/9swDFC/oMnBPVxNA4fR2kc3NRu
gD5sk1N3zW+qsF1k6Td5EJdH7geiPGEE5+i4cE3c/pNKqH3A0Wlc/sZqtHGPpyFCYn9xbaI0y3Xe
nWtgD4WDf5HkWwDiFUoJDHtMuIs90e4U85xlMCV80t/DAHk8rvPCe7K9wVrm3PiP9w19fNBf46t+
mUFkuM6XJNu0QWAnRVFtjr9GEBCiszFbBlY04XVu3GY03vCu6QlgEj/Xj+qqE9JOdHxzYkDaOLp0
1Lvhf+QE7mUXpImeRfvgKT+6h1sr8uOFv9BYxdUOs9CTzGnP9gA52PXnOpmYIu+5u9Z4fI62uEqj
lZGFX79UrFD7hwQWMlwbofearCHcpVZBcLeLB6e53Jdvqr82bJxjMAysJ3cifErfwulK32SFSsvW
OiiUwPVcXloqai5DyR7e+h1SbvCSD0SXqQghxQ7Ao+9+Uae7PwpDWYAFfhtPeP+d0ExyC4QuQYs6
WdRufr17V63M8x0l204i+vSovjYTRLpy06ybXEFngHvLH5rKl2mjBQGZ9goYG/OUx9N8Gisz2FYI
Oucd4dCJk8WDlohCVUfCyy4hjCiDIHRd27zSioDUnrvxGdNNgRleRxknkKWZ7G9K3P+SAcdQfZ+/
xEpg/lnjzDgSkZcLkroTtN3ruyWstuoTCOkp11PHJMzmJujGojmMfO7UJzc4viishMJAIla65fR7
om8IDKQlnCpalDTqPK1i9YP/e9C2uTZK6VpcyGRwTZvyr9/31JalePvceeJ4FETB2+EwYKTh5O1R
P2+UvopKM2H3PajRDzZl+YBf9d68jrJYoBu9H02aRN7HTljgs3kPP7b2+uWvjM7Cuo8NTCj+dDDf
Q3s3M2cst5RODJSH+QLQLs5WJA7pU2d8wPENc4IzLj6bevyi5L/HG/tUG82ZhZI3hTTw8JK+mUt1
NKPkgV3SdG+ZdmyMBqQSqckEhFyB9K2ewMTQOtPVa590guw3uJL+EWil7jpUwKGtSaOTSSUH6SEw
74AWoOF7UGE8P+TvX3/+jm4tMalAEjOuaOSKdBo7XbLpr3ZGV91tk5BokxBSbo/eAqJKElHe9HX1
Gd5c9oLgNoN/hrGULNEuCCMmThaupNbSsz3tEf9pPSYaZc3EjQw5Lx2nHjmXSSokqIK1nrmFXb5l
J551cXrIIeIIgzvxYcHhZDVvwarynpi0EoBcogfXR0RBziHnuoN0mnToCpwTnszawHADwKU4UR6E
ABv12jeoyljf2UDy8Mvdrn3ketDGxfNZceXcfgmUhkpeNO1Cc2RraKubtH0DGhaTapYyoWZdOOLj
qPtwf6sQHFlv1BbBEh3FI/6MROEZHY1kNoI7P0GCQTg9H4M21y9CUd1o/nnFerq7qZ9pwPf3uj49
36JzdKHxK0fAG03T4AmM1zstLt4i+7+T+N5vehY6jD1qoveVw0rfB7cckiNGNAC4zbqH/HPAyEac
ywod6nx+m6n4rE0+PFP3Vm6SJIlJxrKJlSKQaBbsnKRGDNW2HPZdqAim2t31PvNx0satKBGlY2xt
5fNzDR1A4cfPdfPYFjhmKSSaY12/oh7r9Kko34vxJ3cecwJc/+B6/ncpChhSGEW+ZXThruDgA9Gw
1s6XtdrQEp9KSQmS9F5c13q/mdeNLRJEwIfuXPHiS1X5a9R0x9dYSAWIiC+xl5czborSetzEjhzD
4Mn5qypeO121f6/Jb5qnxOwUKiuEDZlwzR83N2MLOLf95ES3ZxoMNYWygt+bL+5Ye4Xslw52INgR
jnvAKDz+rtppTahH4B3jtbksduI5vROnHNfrZilW1R5ZurpgEjta/u1snVb9KYvUdPX3ZMBS2N+E
LwNe1LdjxmqsFZeY1NR/AZxYy72S5FX6hPnnXL4f91J/6D7xZ8N901iC+uEHoHyK4+I4DHvVdRL6
vAmLMdjXlX6LxfocZwVZBBKT/eHl+NT8HeS0XE6kTB+23w2zBexDbpTeglRSApwURmTJr6y/ihmr
YGqUgY9aeQSUvbBDhfVYxsS7vgwuV6b1zZJfKdWlFmPeny+Aq01DrF0wXj9vlNxBFwBzZMbDaS4U
TOgiFTwxUxOQ3asIvEco/BzwZCf8KUIrs9BPGbzbdEtAExHE5mclyvxtdkJ6J2VsTgWFyp3w2hRm
G4QLQS3gnY5q0o1SYdOHAfJH7uSZwpWCZocPhFXYF3eT3TY7ePdC1JheZ+Q3ruxfSBNkOu1DL1CD
Ps8B2sh6ciKgublQTfzFQIn6p+PPnTR4fGdsXwGPtD1hNABydmrYQsrtIzSz6AxP/krwwwOakjrk
A+yh7kKbW+gARrxhoVr/SoVDxfVnskPyFcjXZVqjdw1E6pfdzU4uuTZ18CczJFlifRs+nfmr2g4U
cy5GlCZjLga8IZ3PJsnDrcUqee2jLlZpcaVFLQpjNpHr5ZngX3bJ5RyF+VQF47kUArEMhzBcuSuG
qOEtQ2en1aeVxrcVSd6N3r65YfUZ3Hd13+e9wArB8OYcnysbLkiIVoP9g8AU/QUPGaHpWpJU0smM
QwBnK50/f+NMIWhy4JkKfIW+E4vMXF/YfUjntTRtKIaNjq1Y8zZbm/N0clswdTMYTTBX0K2EkPN/
wXkDavw4bGnyZPGESmwUUhMqKavUkRoqfW7p0Z9maTya63vCFkJZ9diCE2+I/y15PLN2Nbzhy9Aq
yK7B+0u+F9BFrYZNs+GSb8xT2k57NAyBq1cop+p1FeFH9vDvaWQxKYz7d7d5kFaN/iRPRvyzRTYc
v+l35ilyrOeq30C2q602NAX7lvjrO98QflPHfBS02ilSLx+B4rL2w0sGZEvuOTTo5U0YqTk0ldvz
WJMafckqz98MIgMo4D9T/VC+LhK9CePk1TCB86jlNMUNh3g4/qme2CipjT+vx143cY6/00LyHdqM
TRWDnHehThg6421i2e4okkKZ1Fs1lM0AZpZXsduJK4KJTPOLTsjL6vSDbSbvHMJTCuyERtwK/eIC
Sz706vob+gbfAkFqsUYA0QlMDApoZf9pz9SuLd2t36HMLBrkW0KP4ex+J3ztM0O796bIpmDkioaZ
Xe1r5r0kPdsd06mxooaPQukTiUrQodGTcG0bT+zkLkMnF0fcIqBUllt3EeCfYOR6TVsTwBG7VA3a
eiC08p/doeP/6JQ8JXvZXBylowpM8X0AEpAQcfErY8D2NZirKSI+JKApx+2iSpBD9+GM+wsoO9Jv
dvaNnTLjxmLB45cjgjRgyeG5PwKvmBpAyrdYmytHmIS2zCZIluCm1SAeub/YEyx26UMUgLc/oCLm
3w/b5HtxdBUC6fGUczTwd4xsc+37fwit0jx6017FyfBeFpK8hXVu+uC8d+oahD/nLhgATKRSWhEL
tmAlUjBYCjJVkZICKENsEmjaWaZsVw4HtpW1COmNJ6k1/XegK3vRrskiJqP7xyTC6M2nuduiAXoJ
jIoj6pu9Aolpwluczmhjvomt9GIOLVumXVP3rfX34KxreRx9sOuUfyMSZ9Hjw/RPkz9IFUY4FF6v
IFnjkv58EGmATw3e3gm0xwYe7oyXhEcRh2RwKlWK1MG7AiExt3olS4R/IrffNdRC3wn8Fqlwp440
Rg1d/Jn/m1g953sddSIFGKK0yXIoXVy28KTqM7VT+IyHIlpcz1mhgLcW8R+xNNdlq7NV5BUbSZsp
cEboZ4z5rPsWZIoxDBwEjWQ1qkvDK7vGvGKUwZ8/Fz8a3MhGz8gGuqghadq68O8Yi1W816+S7nJG
02DaWC/+nGOYluwIdkOmYQDtJIB5hl0Y0qTeKJhOVuR7kEq/20J2m3xBEzojFEUjPMzGaVGxWFjo
6eIct9BnxWuwCRf0kV8i8rmvWja7P1GOk1QDOjSs+Mp0wMTzlq8FhF3KG6BqJBtVPklhpZl3+GTL
Ws+7xLnmC3K4sbhqrjUqe8yKWHbmPRu0Zk1XyxECAqQRVlfsEcX1UWkKY47NuPkjqIFYLQLC2wIj
IHm3KLyGdhiHlHiH3+hthkvx0Ku7PHvXhf+g1ZOvVz7bpFcoakBFmsQ7zhVTPOHYANutfMqQuQDD
4gVL+8ANNO9L/5w184P4nBWfszDWFZ5sUQfMRs2cTzXcoS5GFwQpnnPf2wLW+Bb48vWsGs6pIIAD
w32yyLDY3ynyQxniqdqhbCCvbUUnXPSkPKLITCpIFf6X1gUJvnGBe1tQA/EbyQpU7lGfk+JMaM4q
Gq3P+b7hfAJiec0rDw4m2GE45tRD0qIacQZZQ5Al9Cc+NUj9xa2BjAS5C2Wnmu9vY78ldBOXPp2F
BijEUMA8Gz2B2pCjas24wXAf5dsx/P1V7FtvXuKdU2OuXlCXoefe5RW4gTCyPsQ8eE7GPaOKpeVh
YfM7O46RuKqTMNhZ971yAarvJaebwSIWzm87CaQZhcrbbonVaU9m5jymXlchJkop68yeLvpZOsHB
VWgqJ3aYUPIHMWTIVmLTzbj4r+8d5zqZIXn+cXAl1MFmOavmSZyc8IEUWv4rV6TwwFLUiGNI5koM
Mp8AQMIZIFwCWHgpewvIEzlkT5x08F3QNus3t9ZPIdZnvRnZFvz3CSCnzI5lpj1LGACJ4006gJA/
5V4brE+xIy04TDavDj9HEy7VSnOvCXzxUruC38N3UczTKSCpB43ZtZFKPSvtoMy3v2gdbluCdSWX
5ubBFKbTOo2boAwk9z6IjPMYYwHHkrj5FE5xd+gf3UJByLOVMQXMiR/MhSQ9zIZPo5TTgU1YNktW
+mCbYd2Z3rhT4fLxxvaqRBkqTXG7EvrL++qr9tzqfGAkzVw1G83xYiGHhH4/AfF0kzxT4MIAdXlw
1kGza8rz+AgrOXhN4Jfwhlh9JKPwtl+70dQVFk3pY5O+SjfYFZLBhkO+yNhz6UILCEmqAlusklHz
M39IxMmTPmm318T2SzFkr2eglAI7L0XjsRih4wM6wM41cGGuHTnVJwdql2K3kB5zYMvewPo0+kYX
44pHAt91SFNAoMKYFSsLCJUkrxfdsZ4brl406STnc6VVdkLJoL0tgkrobqO1/+Oy3BJk06rNYwuO
9WUEEUlcJ2lFB2iXW8rlYrKLOrzvVqG04DY42gAF7CTauDPfSg5AMD14zfgTdG6XGcsKnJzpZfMv
5M6XbVpOh5Tq7HE+jHbXSSnzr3AJ2LegAGsh2OM/YVQPH9JfVEeLHAY8gjUKkkDelgPfCWdb02V4
mYsFjz2aRNoE9u1fdcVjjqPBgGg2PvcAX86MYvfdPdYg91uf0HP/710KX1JSqTJxqNTiVf7n8lja
Tno1w+LpujD143LlYzb/XCLQXOKSpS4cja7SKD2Jk4ecVOYLV1/G2x+L/YoXE4FJXv7CBw8Ms73x
aJF6K3qvveUP9B0b/Emt/sCYKzURg8OHKMUVlWKS8b4fOVq0kwBwni3YjHVaWxA2vKyGtGKo8Ejl
HAG77cHp7Q1sKp2yxLV3Z0xWQQD90g3Qbjjo/3yiy/UhUE8IdxuIAKCcJ7e5nkj2PGfRzoOVn4Nm
YHeBuwmCr5G99/ptGBuJt9QRjllysiNMO4uYl8pfaMxR3Yin/deBdCrEzD8beE1dkAYbN/MFTpPT
N9VllkrN4ITmhn6MoRW+HYXM2urwsBls1wzdkv25xvjsdWseUoMxKIUV3qbGfhsyyU3H2sNIMYXI
uPXQ3Jmt/S9dOduc1NSJb0s1A92PZ5uZwZO1adNSThlyWDFfEYe3Uhx0WvIfbSIASIOCOceQ7vBx
blUP7va3Fxydazla+mi9LjlZsd+sDDEpW2YyaUkBB/ZZNkMP1gz+ukx8+KyOBxMbQpNL9VB4QkGp
/x8B+gfeI21G+eAB/X/Z7K34teo0VZ3C0ccWo7YeJB+D9upigc2Tb19rl+HyYGShHiQoPAtuk6bG
Dk/YIJmUdX1jwdXpr98rV8Ni77sQzZaIZnGJKK1O5BsojnBrWrA41c7p/qIoz2rA7RWBL0DvCU6O
Z4oMR0XeOstiaZgTyLZuncoHw+VyktEMh+3A/aUsDMrNC92p51s0qpSHiZzmE/V1ePv8W7OzeGnZ
V2f7SJ2A8aCSCBR/z1mSap5Ji4gR5fwEbwtw01xUlfskYtKMB4wxb/ch1AYC/OUxs3KX2nXv5C+/
Vno1vi4cn5CPn5NiiHn2BN/H+DBEoA6ldjXbSOql7BhdS/R/hKquMG1sR+IzuHSa5GLfe2nsgRGT
Egkr+pxZuHV/QGhVz3iQfmefJ3OuTp0CtTv5pz16q7z4qPxakC7gBX1mGsQeImMwn7Qwe641MTBN
9WZ2zf8wAvafmKc6dc20X4uKm4lZN8d2d5V/aWJzaZTXVOZ1ynW53YnOuPH9VTpdJy1EIDUkvFzH
Ry53NZ6lC3/1oPUqMYf2RwYOB+1L2GwVmQWfze+8mkH9K63IhTqGs3ntIBYiDX0SUUdAETmnMXcJ
hlOr5Cjde+XEcFGEurdVtHtDttvfWBv6hvgJ4yrjKlfgT4BDClJ3XPS0Y/FwNNX3F7AwmXtMUCEJ
I/OOe1QTpwZsNdY+uLC/b8P2vg/6S/oWwpvqK5hvKm9fpjoouBAbX/DhN0C74AjsU66u6Wpct7IC
0IUZmDOZpjRATwNfy3OGHGst/jyFfnsqtYtM7507be/+xmPd2N5e3aEHKroyMgjg2tYSXiCYqzI5
OG/Vlg6TQ+JfXMX8YKldF1bfD7109MDnJHW0ueLRhN+X6gWVCkJIKxlwCVOMCv0hTYa2i+MF0j/S
c5R+p9ojmPSJZHg8kMqzg7NHPAM195p37Gvzzok26Xcm50Cuxx5GgKs8eHGSRcaN81Rs6KNBctx8
5DirZ0ZOQHCRmtuQM6olnhTMzfHxu6BoC2pFA2ZbXXFJKRttmRvQhZe3Z1X/xAo7MkbF8pOmjeWV
7Rg4+DDh+hN/xOXnrsP677Xr0m5Zu62K+z1EEJQ9Yx9vcJwMHGllTkVXaVy82Ctq05pweMotBIbu
1CtRdXxBy30zMx62IqtDVsn3fXabtW7uapXJRODLZO8kKTFhgZPjWoxjza/rEkuwUpptdgiN5KcM
VBOpegBBk0TPvkCGh7s+QwMEu6IrNPmWwPYOH9nMsuKd2ds4spXFLHDuVWrvjVcRYq2tjnbt536W
Iu8urz7hC976vladpAL2WK9CMIXSvempD34J8qoHUQrlrjIJ/COa0udE2kddUoE2hdGOnKSwdB4X
f0TAivcOLYFzi1gOIJjJeWIMnJIVkzpqjtwqJAIDJY0xhx7mpWQRfu90zkrER1sYeIsmu++dbjpj
8E0gwaPhhoecQZUVGtB8Mat3SpeivR6I29GhUv+yD5uNKa0659KKmNzWc5bBTklC8DZMEN1JCXma
iRUdolgjDHMNqYuFx5RqyIF+/P5LL5HDf55yHSJD5d5fe2cRClMQ+3YUABSqvvGZSGu1QVYrZzz7
ab426c64GkTSUEcz2pDA8RSVQJGmNlWiTGaFeU1cZaPUFCJU+P+UQBFVu7Ogb00R/G8z+V84Bsgz
m/p5hiUyAvOxNKLyefiRliorhgwdL8PY+BoX05TPsFIJ8qW+rnPBnKU5cRWAYshlnM8X0NffBdfn
u5DRzhjCFS6vWexMYGWnLqLIZQ4U+dWtWtIIrF5+s2pqHDUioDFZn4Ey8bsBlvPnKE3slZ6YypZq
CXxT2IE2Q/9jnld+OC2Kq4GGgNOrD/fw1b8gEWARQX8DW1tXBcExu2n0byHmHloTzX9hpQ/AYX/N
t+gJTMI709eQRE/ArzwXpyJS7MAEeVCx8vrfrZ7B6euZp6Zs1jxBBto7VQFRYOeXCk6GS3TtSBYa
+qvrEVa+HBa/eRvvsazqA7kN7iICcSC44QYWIpVKMsWPlLoAqOPthVMZkRi0pbV8oiUbvqxTAu1I
ETPoi760DCwskQTdy7if8vZ21rgF6LlFOH79j2v3FI6E7jno30E+0Ncs6xIS/PzBRz9EgVB/TgLA
sXFVsFp6uSRPAtgF3YwlHsbFZGs8dtN1CZOP2Doyd5jr+UwU1Sspu5NbEnLHu8pEAczJg4tCw3KD
YF9COOLETh0J6YyYrcROK0x9gWYBwxP9CFOd+M5yGblaAnfXQImM9GibfNHJ6CCeO6QKgYdcsiLy
2vi4+gWA8ap3O2UCvw84YCfyqWyLYseKk3K9Q/saABsr96ebHHEMc4E/UDsOqddQgepHnTOCUKmL
8DZDqf2iR+SeIdf68pZjW8Y9hcWXiIKEABVcp9ERTSvJDUqnMoINjH13QIf00M5CIBqg9HvaYPEI
1iNKpRXgVTsg1sZjb7/VaWEcwyJ8HF0QJxFsszapqQfNllNztslg2nJQgK/LFYwyP1I7iLFIg+ql
ySFxjooLp0OxWlnHGPb4U3L17Wsqpr5uIj0F5pxqy7fn51otCFez5XxjLqZT7C/9Fkev70DTN8Lo
l4m0nJJZNj05CVisz3tIJ/W8PLsm8RaA1GeF5i45I7PTM3rWSfbKTvADhGyrr4bhKIVc6incQIBJ
xNWyh9+vReaWyeUhtNImXrCK/wJ77XgFE31vLKsO83NCllBSPO7cWqkVTQ0AsBwxToHhYqffyv+Z
QCNQ75r8rsZW9zLRPZblT73TOswuc3xDuBeNBEHQLEQyI+lgOGc0lX8X8cmr3jYTTrvjpYdZZqZP
2n/djPs/0UirnOhpqvsPFs65L0Bqxbt8BRDeas32aD8znFoSix59/C9mw3Kkg2O+4T2RLNsHlj43
kmNOWWbJvKfl19lWB9ufhW89iVnxrPRuv5RjhUBrerCHTZIyhxYNhM7eckjaHr+n2bph8NpS5WeT
iRdypkXVBT97o6iAqQGyGS0NVoCW/DalCbSemI+ocVfl4+/qcuNgDETmEDzYGLMFRtp4I/dP37E6
F8U323NV1QauPwBbs+DKP3QAkTKXDUZtzSormEMaS3klqcK70pW39ZzNEOTF1h360NNyHsmqkIG8
0Vj2+xJtB2POtO4f4FKcWVJNeT34lxC8PvQHzFxsO0IHkRiRc+o5Q/St0xMWSIJB1jNomB2yw4Cr
K/youN0hycNEUTF8ieBSHEfDKQ8caG4C1D+tcMzbe/YXzb6VxdhmMiMvvdolrGP9Wv+IRRJpYhwC
DhHFjPjwlvFPJPHRgop7KsMU0wxEA+YtSjKPkKKlcHoIuTKFEBFBBxCN+Z15+BUlSv3ZPNwkAf40
2C8oppjmZB2m7Cdj2eC6tCS/tmRjUImeVQ2uhiDMk2OUtkWPAEcNxM/gat5hMphrC7tBBirOzEqW
tDd4LmfqEe3kLUCYXvgLK5d0wVKyPvXwAtekBHJl3A2p8crXs+7R30nGHbPMKeXeeGFhsnM7w/Hf
PDoqj7dk/VfBZJnzGmmFhuuuDWl8yYrvgeejqQE0jPKB1Y6F2vMSo31stvMyAqRc5EHa/V/zJWIc
ybHFzuOQ//KVUVWZlqXGllbseg93Ef+fhs1MBPNUOtWXK8lDkR3ARNEssJyfxIIulXBXwQUYZZJg
p2dAshnsuo16uzvfCVE/CSa9FTk4U+2rB/TEpJZCuEIcZL4gfvgodP0TiNogL46t1Ydyc84zV4+f
Ql6NlKKmG8/j07gHW01FIaobjM0jAxRjd8pL/xPChoQ2ZcAewg6K5YAIUBrLfhx4nEIIWFQr8Rdu
mSI/nSAfg27Wr/Bi8YzE0B3IY9aHmps/bC+DQZAZcN8AjJGiGemWEIZ/D09vqTOur18gca9/u7zA
nnFK1r4Oei/lTlRujJ1cL6Yg2kgakeQx/lHl7Aed3KEd307MGUH20LLH3ymYbE0fQz8g5I0MJc0s
wxS9/S6a+iJujSA1DoTe+NkEryTu6Xm9BMwlTlXg/Y/X89g7Uc10OAo+s+A2KneAZ4aYZ/JGEo+V
liuzF4Sv+wcHYtpSyYpu0PbqTRfSPxX/e5a0h8fGyzlaXgT+jQX9cH7sOhs0cLbNkpmmaT0o9LoC
QWyqOhUpsBvYjm2RQrXpCWaXHhijT8RyXeysHGNha4q6YIjt5MxOnsRIxIVIqOaY094xW4HpZP3s
zQkrdEekVUT2xZlN0moiYMxK/25t56uA0/0Lil7zH09vgBmspXZkyrtYuRzqSz4ASUmjZCiTdOnH
HOgO+R1vBOhvKmqQwCTSRQBs0Nr11UBM7A4e17XhJPtr/98izAbZC03igIsOVH3ueAJmhoM+0N3s
PNrammDogMCia9o8sDwVccjwYbccdrWv2jRfKcdmbxCzlBeZO3uGzvYClp24lwwgUpL0nCqJHT/D
j2ot+qcSmvB0sbAOgfr5hnafr3tgjhKUdJbs7DYRYavPSisWOYv9PWWAFHNRn/KNSLfAvXmAUx+N
nXuKj5+Sd4xQG6PvDFHDkdfQU6b1tK9+LmpImk/32T+VhXpCUf4bvlRrRI4BgHlsCYL+UVTZFuPC
Cs6w0juZ4TRQXllDKfv2vgldmlktLx3i01bR3r01E6nKIjhzjyT348M+BKmYr7m7yMngSvjh2sHp
Nap7RDwjVr2Q93tMa7MMkI9FKG3tKeMU2vExidk8YgAIFT2NrXNuH+muX+A/Uc4COXjzTIOQtOSZ
tEa1hvQvewq+ZwFtE6aT2YLJp/iPrwGrmluamiGfrIO5xSbh9qx4umhwFUOxbQmiyPSRWNfcsCDu
mxrqtpL2fMpEOjEHWKMkM/OhsaSKBRRUS0NYxfYRdGX/MitktvPuhud01KRib92xiRWuT4ZxppqB
Q2VHqLCgqB8NOg5nnoLUgwjVd3AOMx86tseyfmYbQHTTBg/UKWKJoWsHV6Ld8tHFsSkwLiO4kpH+
kuiJBPkg4FQ45IEN82jtVabjp1+fTVsHUblvbyypwGaPYF+r/MYh1mj7pdlJAJfC7ibUavDsP+eI
7wjliLS/tr88xg7rRPJ8Bc9eydXbd9it9YivYiAXkFu6+fe1ex9o4nCKJz600QRKz5fomrnLnPBA
CWHnMD94LmuZU5+OPJP5e1+AfiMMyFO6h489W+K8Cs9InE7V+MrZ7Wy7B5UEY1Bhq/wUGyLOUl5T
GQTcYGSeBzvvW6V5UclFsyqTJlK3N+u9VGp6x7NSMqiZWDUaBLKsKZb6JwGtjRSqLwhm2LYXj/0h
L1Ki0jlVAJ8bLwyQpvhldj9vTAcOE0HTlRA4W6BSGfOPlMt3nmxXr5v4POHXa2pikKn7OtHNAWRi
gBP8XHvXkQMq8VPkYNfnajQLY8YBZs3CbYnX2CVT5W/owvYLCtecOtlXN+yagME8W4ueSasIdz/n
ACkPNeS64fkNe0PjDWCz0zyC9CK1oaWh7ZOMWKFI54zUwGMzBmlnws4IDkPWg847pRqPl6no1j8t
uk3/BZ2FrC69Ka7+1RJ2BSwFxgyNKiMNkBENsUbc0mMc8pp+Mb+jv5ipEgiV+0cbqG7YldeFsRy4
Hrj37ghQ3FWDAKiRVZFVIWasU7a/qzTW6/0bLI4a4CcNb3xmCzy7I7sKvEWVvAUmvqxUUFgdpXPO
lMY4xpY2ANal9ezUVqsCIsuDHfh/vAiIrer3eGvkxiszFPiDRIu1nbVN4g2prevGgrcyKUf6Kuuj
tN1SR5S2ld4tcKtuRojThyyXsEVf/92hUusMncO9iIlNdfq6n1b2ODKflCuU3LXcYL0DwmLQ4d9y
OfwkWcXwGDdVMZMEcZj2lz57Q8diAXH+y8siRpPID4yRq0DzxDdoBkfbUHXhPMzYcRtZbtU3Rfvv
mBxgNj5bgyGMOKKz3nHJ8gzchmPm5Py98BrEL0nEnhQ3B6s+Skdcjzb8vjRS3mUqiDUpMs1Z6s0r
wMARWQ2zHBICSbrdtHTYZ0RUQaGAja8r9fserEq9tmJbKSHarxbyYdxhpvUhcur1qqSahy5fBdte
d12NvquATtikqR9xyt2QHwBA6FD5OLfjcUuw76R8k6o12p+zZd8LeRlAH9rGXs1rpsbST7xgk0Xy
H9B4PQqa+KQkyxvzi0BdVCWoY2yvxo4EnoMzVxuFr8o8Bx5rRIQxR8MYb54+u3atdYFFZk3aTKhu
k7poiKJ5YPpcfllQPUjNmxlHmpIy78dgpiQrF5gkacmGLOBMg0A5nUL/txP0WpeJzBTbopac/zX0
QPpQLUB9X5S/OttlSDgv6+CoG4ZL/GQMx3Rl5I3eDYNIPk1fowWbGE7E7XMZaEV3ZZ/DSxZ99/pS
6QMRj3wt315GIOD6+Se1v9QFNkcYcouMiYmAGNQ6RdRZ/+upQUX6LF1hNAl+lhdLoNGJ3ZlInMVU
99Y5F9Hrc/Au2SHKsK2xESE1iZI/2Wi7mrmkpJs7f/XggUXDzObzAsFcHLx78WkOmVWSwsoQvYjY
l3ojxDDqsTgmNYu+N2UI4lbrBdzvkmMBSZ5Z2kCM8tBajbEXtQGUFszy6ivqM06XdB8RDthVPHKX
iq2XQi2K+PV7MJQDWXzUQYl5r01XT/CfG0E5XG0GHzJgaZzLTD3jJUI49ETovHWDZ6rEm9anJMXf
YoSKyZgyPsosfW63To1m05L39TtvyumZSR4vvXUagMDP3UHA8gzLG9aiKy841DSYoh7/3i8UUZM8
DCq4/rN4RJx04sTqecp4GqufxuRd+0PC/rCiTUzYdPVO43tA7XJjoaMfJqJoCCDLtkyVdQiiNy9j
HHphwutFGWk6xyqTlbagAsBc7LPv4fjH8wJswJPDJwN2PGukhZqsuRiQjvK75Mcg4S56DPzDyd5Q
pnOA2ivBPeFmSuczDM3UCdQTWlpc6GmBQtsPV3kYe77dCIKNlPN5F9MVKJ3mcir686VU05OiZznO
Ylhy8R5Bdjy4BB5//r9OFCv1GlM5kqwkL9Bjv54mZjZF2YVey7JxYHCrLUxvMm9V+er02YtNz/R7
ENgNnmECo70U5EztXNHvPF7yHNGROJAs4ZOKba3LvmPKjG13qd3nvBOLg23QnhZ1/iz6jz/svlji
psDo+uhF1wEqjoyC3NMjK5XXzYubC5q/jJN344DXPjGCuPnw12cvkFmBwvnEbSYET1wzySsIhUmB
S906D9UE7jp2g6xMEI4UZdryu6w8GXIxNbUt+5fc1C7F7DB9A6ZQLGygI7SAc0DV/XwAZphDSJDe
yDyTwzZU30gqTvGjb2n4GjxyKgcGolTryA86fDHxb358xm2dnabg/W7cP2Kmk6E3ohKnMJ+FwSdR
x6BRfB3VnC2zruUH1km9TwKPQ0oI7jslTm9+IrGL26g6F9INlPTzV+ee1TemZVPUjv+YVqDutSvl
rL+A+1tOILAp5qWrfm/a/RpJEP8s+XZog1+6kIan7tYmlPDOduV3Xw86/pdcqchGsZSQMVPEsSnt
E8NsmgHNXqeMCPTYrA/+qDN9M8Fae+LUAzyzvrN+YBL3pzZqJQexqbhG4I6ethKJtprkjgfNGivY
hpsztDkiFxWALr5l0Sd1B2TwBpX9bcQTrfuoI4QsbbHU7eMCnWvutx4eiE8b1jMFBD3N8s2FeklI
QP2IVmXn1z1dLYzzi1DBFiBbxpEoqwj2mPst5891PANgoHmHjenttW4ios5EFhILoqT7c8A8zsC/
tSVfWHn1LbFzwNrDmLOr08i5jXgd9uoRiXyUsIMqQjkHzJDIaBJJEa9FOhIOI5nSVlhu9jsbA0OY
LdQubzw2qpRflAd1O6QItH2mOrMxBRjW88akGNVApzHRn0Nd/zMCWuXdvf93INkRF4aJUlWVR6Uw
Eb9Q6UxPORnW/OrXQBWWEMaHnh7c4MPhbo/nPxQ4pT4v7s1f/hY74ZdG0BPCOnaUEjBUw+mHBnOC
cXSys4mgfxovu9gIPruQ/CiF/nUAkWybET/phaEitT7oyg2dao3CLi/22270X176ihun15xoepbh
9YI0QO1q8ozIa6DIeztydTlQxKbWKOgkRiLuYTIbJ3YiGdR0H6sVOyZwD/P9ywmclOhx/NzbxHvF
ZPQpdlndtsbB9x/TDBlMRZhjZ2HwiroU81nY22O15BxMRTzeYDbBc1cJ9L4vmTYrLg/z0I/RxipG
nSnjKXwkmV9i+4c1dOcNItyzuF5BeipqSceyKKSWK4mPdQTpS4wX+3m0QJ2MUf9RBWQ1y327489A
wMln99fPmlaOdtTD3wGn3o9edHKVCIcVu55hDVC4FjLHg0qn1gmpgDW3IPGCbYB9ZTpxO41lOEH4
OVvSfE3AiCNDXF7NPqSJma8tsUG/CCoTWrs5Ioiy3mtRinUrZB4W8qt1xjttkL+QIdaiWWCs6341
M8xR1DEw+lrCUjmjqz56M0jh5ozSucMzJPXMuYS98/E4qCtEjpRmbiXlu7tn20+iFTBXhFdeLWMh
dKysBtm+VDSr9dy5FEKjvkOtjdTiBXtW9dBVKYRnkXnmFVWzIggvw+5fJB/xEIV5J1oyMoWq7CzX
qlKhj0Lb/3wMDXbh4cNDOp35NQz4TSY2gObWek8hyo4BZniM99x/AB1byetDNQ6BDwTQiEBWh3WT
PbXHuSldssSUpvrToOpv716zWnUo5ns47ocxjxYMM2AdtaPpv+rqkaVoTvguX14yWJ89b3IMYOLE
75poBoYZgQ0qVuvM1aPyucbtnuY6is2G81VhpIhwXOHaeNFuUV3A1QuLTRU2K99WlmCT9unwe4Ib
eLc0NdsLDWUbMrWwF+YPfiS2mTrmiqLzSFGJ7hCJXMr9AFGyi2o21z/2IJ6NvymL/peH3Ldf9g1V
QRsNT0n6N66M8/P8J9wnPod6a5h5wnhEofpt9JVmZJzgz3KKxlSDgSAhiwRHDi/zmp7v5gxe499C
M5kcYAiITcL2HKFv0h+kYLR5ZSXYVBV+tKaCrcE5RNlXlSmJqvfiMyR0CiifsSQFfN16ZwaX/Nfb
rEtuPJBqBEJ2riPjcCBLbF4dmJDdt1ViX863Y5UfsSxH4RbOVBJQsqCOyi2YHvyyUr1zWMiQNAVv
btoxO8IWJKCH+672imuYxU62ned/3MIQTBBJ+87UCUeFTss+6YNZ83NKmYuoIw144aXnmpSXrQdd
muq5/UkRlA6NJxm1orpAaUMLXFhlm7EVeMaPR2ugFVN+oGIPHWodl5w8GdnrXB00I8chu3EZE3Kd
evtVA1hCaxOo2/pBsVgwjAtYuzSsuDMgbahyJ0C9QflHSO4O/gE0bPTQpSp4gaeP4+h1Ehanyihr
IE1hJOxvpnvfqZPEXLzRzOqfc1Sxg4OOdRSHa6JAlcYh6JJ1cdUV/yuVmdeoGx9tsvrZYcgjrtQG
MrMeYrwLqY81CdMCZ4YqI10/tdmhDq+Gg4tSAku0AzA1LzDAI7Wi7CqTpgf9slUM25U2EdBG8heT
VXmiInCkHFqtJ6b2YqyihJhqn+skWOmdazz4yfW82KE88wU1tfXiEURWCsL8RixWieGl/+0QCpqF
t22Okd1fpQ50ICtDC80LMURTVnXKdPGOT31vgUcR073vJ3sxoVHExxxOA3j8GT4MtM8HF7BnTikG
Sfe/MjFIuAVRBLNyRVHrjoGSQqCLjcIxYFouB1/WruSDiKz3Wls06crMllRtQ8jbsHsOiN7rU9lD
aYUrRwVEq9H21POW9KKAM7rSMhxY0nWQhxJ1GZjm7n3gfAPy+dUZSWknj2LhOPWhkdBYCvq3zL0o
83n4wyrWL+X4E6PqGdqT4v17krepvHj2yhqE657ANkH/qjR8GORIu7MIP1A5njXrKUDrdR7De1bc
xgN8pyviSiuMYuonEJbCpgakgNitBwTm4KqTIZCE6fex3liZV0mn67uzk3Fkfj7b9n/ofN73Xl/o
Wf8HiXJgfe4wH3OXjv0jkbagw4AEdreqaYyFVXGjC3OczcpdoP2rFVEtby8JYmCANL1hM4pGy3aw
O7ZJw+8ycy4Q92InxpfQTIaEVD78noq/UwXkdbcj1huKBFM8npKNyTmK6R2O1qBLbgM/wSN6nvDf
xpkLeRnzNR+jks2TGpY0Vr5xhVq3PEDDlyrIHkZK85OwQA9KgCd1OjUja0MJR50zc5yNpRb3UZGo
yY++t7ALr51bzNYnvlakRc1/UIVnJ7/saN/WIQ9HRXaTDrTzZpAxks7OIRp8xmEN+Nv0NvXZxA7K
n2dP6Hz2v4m5LZ8Gcp8lIwd6f/JCTtwTIUoQdIIzkd3D6GIChxptPtcXPU/uMj0WVlGqLKFc3lSJ
INm+IeDweWANcviKoyNiePzosL/JisnFw/1HPIKksIhfcRYYo7MyI73ojPJxjgO4FvJqnNiwoy8h
Ws08SPSnpGOAcKZlyZYf+PMlJp55/GjsrLL79o3ljpXLf3YVUYc8noaM0tujPZjqh9qNiIKsUh4w
TJMVRNRKhCYv9aGt0lzOKt0eBYqNflfA18oDmDmGhWzUqE1fhAi7+hiS0WBunBLQD18Dl0S3Dx/X
E9KZfEoVg+s/waKwghcfIhpwKdBTY6Nwz8XWPj6xfiF6MXOc5lXnHb6rRHVXstHL/dG6fNSDRn9r
NIrngjjfXTA7rQD8YC6MUoHWsuXvEYKajwlWHXxNbZVu13eJMQtKopUsUMbcZWp3B3/4mnNvQ1OZ
FdwW3FVVAo/O/OmMK7CSsDnH+SP0tMM6JWOvKLCO7ZetOKDPupmv36UPYWJk6UCRSSifA0PXQhSH
UgWWwtDHv8ZpsK34HHLJpfh3sa42Aeced4lHlrSxYt27EnapQ0em2dDziURctb95CEO3rLvuh7RQ
vl61DvtoCG56LA+LJ0cBQ7olRQbqFRX859C8SMliJZSG9MpNqT+MUPDDIYwZj7yQIW4UGvegGbXX
bMpIZbJmYQvB7xfO1nop3ZC7nGby78fWVJwmsz6x0j67boBuzSkdnfGkXwDGhfbDwC1AOBZ+3+34
XjixE3e3K0mFUbv3acSX5xOTB/6MRH3Cc/scoc1+lRMXo+zti4m+99f0kt7ngijbE0mdj7pGc3OI
OZ5WNPnakggcVv6LsN5IryCLQnRuPV6OVNjaZdpg59OiCjeKoRiI2HnrICQbukJT4AOAchMPie8h
PEqzcplEwgaK6rySClxHgJvBnpjLb2nqdNX5ONC9Gns75ltXL5FI2VDu/Zq59iLgBqSIFnCCFeh1
gR3NRa3nQb1ae/6nGSvD1fimQxyswklI96phOfT81WBXHxuS1QKEIyfeUOESE/PX6jtJlyLhlF6t
xu8aLlwrHNKuAPhuyBffD+Q2EL20YUzDEjmVBgh0Ste8BnGmRy2LDhCgTOGx4IBN2iggmpMa5fPZ
DJ9eXaaqhh86Y0TMs0QFjDu2Ff0eFiH8ipdf/l2iXi4WX8FRmu+rCR/8LCfZ+hkehf6fRe0F+YE0
63yDpC3/0HVTtGD+yTQ7qoypbJ5VfS82LDbAhiUF3MGmUCLb9VSBGyKQJwMKj6tqpGBh45wfAkhF
M8L8u872iOFZ1Lc6YGCbaJmNBRSwx8a0tUq5esoyzugvgJks5xy3z7Mek1EUOdgTl2Bg6MG5gYKY
rNwgJ2svyuJX7Qg8CEooFPhv3pN7H5S4SQpiVm8aTZ7Kw8lRrXKuUtVAXnZn2FtSCzw13zp1ewBn
mITH7IsCvIawsMbJCdTxvAsfiBy3m+XuUtuP9DJ5XHMPsfZ/L/MdfxVr5oaL9dY2y+WLqbTiPHsW
9izFdkSlg2vNYOm2MunzbdEHyOcQQdbQvWWawhTKVdZ3A18bSyETrK8PSQeQRga2D7vXPq8pIv+G
nHuOhayehkBnfSyZkDmGkYUEhfeOMAszwdBXWc70nN5dsdsPfCOiresolt94MGw1fvhYYgMBY3lS
zUgb54atPTK6CUKBJkuO1uSVhZUe/AauMqLUZ0zDaPiCQTZXFu+MTM/hdifdcih0+X+87s8TJSmM
bYHeYUGhnKkqmJqIZvvUs6NJ8Nuoey0baNSCWyqtJXg034IOueL5kOY2VOKLdbmGjXSOU1AAmN22
dcrr/Ww+N9KiSEn0S2ZQoq01S6AbmS83bi4I5ofx/5vrI07XKc5fI7SI8sfvNeGffYS34fUiHL4g
z7yVMPDPN/6IOAzHlj/FbibBX0RUPSRoxR1ty79GgJ+XwnBCHsZxAn+E9aMOrFBOBKp/h5aL1pKC
lHhozL6QtZ3HKnQnZXH0h4xEehyZXwF3mxOWJgin0H4giLp+GB7KDIgsYcro42ajv/GEVhYOrOlG
/fb8/bSwGZ15iLa7ZGLEg173TD+S1CqGR3E+ZwzCuYmw47zMirk9s4rPElEiSvjbCv1wFVNlP/7f
2UvMk8eeQB3srqPpovtreexCyoVePWl2+yWvO6hL2z6LhcVT00mWiog23nNdicHw3tzmdEpdOB9e
o9MhMzsIjcLId54NuDFJcXsz3GuK8a+buFmgWQGmqTd7rTH8XvWTdoqzxL9HZQzixvSgRFG/gFkk
Yu0nh0F7FpeYi+m2KTb1vbOlxAszj4AGHKA05LCYjZ7++ZaRk0j51I3SgxDxOIcDhKESrrJTcf6f
N/MyvmRNMNM+j8OVUWx+EEEQru+A+ZwVOIeHOeqcn+QOTIzYv1h/3pEUf22Rthed9krbJGUTNvOX
S7zaO7WcOIe3etP68ysLQ0kQNjKzvdNTX+HHqWCFfGl0wMJdFBPOzhe5MBOGd2WZWzQh/ipDnMbt
qxU0HclGgXywlzrb2pvSXXPpcBl/KBp1I54yGgq/Qe47c7SmcTw3RDEgjtTL9qmLw/0G52bOF4xT
FKoJd4omocOGUR95jrE1qWM5YrAF9w3zZhU7O1hjafkmC6gZrMcQTFb5ONdcvKkLySbD1uzHkN06
eqM8Tv66sK3PlXPMYZBs/HJf8X9bkVnKObNfKoKuT8WzBQvi9nrh+saHIPloAF9uCxGD+sYrUtnY
D1S8AracbRGo++p3fvaAQ5V1Cnr5W32sP+fx4Ro+W54MtKtE5c9I4lBzHZdOcgXVIgbiBqciP9gR
MzECX4XzFLBLhiCipce8LvrTnchaOtTQDMxHhiQqmc/iEtrK31msEkKqAX7G4rE86rNQ/fsrJTn3
6Pum4wTS1iKMUVpP/r6bmhbgdSI8KZilQa+MI34Z4DkaeNba0oUhLSaw4hiuJBpvWVAYMBP8/0HH
MbV8oSBJN9s925WP2yLzf13suXNFQqxNBmGoNtH+dt0J/yQTm4xv9ngsfi4CpQCpwVTcrqRioHCy
NnPZz0093bYXf17OrRuX1AZ0iQoAvbMZlwfAfuXFfL4CoBmvYvWO3IjKnmmfCMYnbhsObmq/k5GK
7lSzc5e90nfb5L5w5C+V2ri4MwRFCMOOQ1LtB8kvG/sGLEoWQpYdWmrnyIUY6JL9kPlvfmdL7Xpa
3f/PRV9P8yKOHmLBERaJ7cwi7EFFjOK2WC7fB+dORO1UZv5y9tbX3rvo7AckCAKtxlv0+aaj79xU
6CDh/P7CPG51L5lNnG7x2pZKBGlL9dL81HfTcAQKbKs+hk1kZbufvKRtsLyHRQx/SodRkyx+PEdB
iZGK/ZEjvo5VU0CD6sTjnq6pqt9bIrzi4ImwN6neT4wcpHkTxJJBTqf5B8fiD1TFMreBTRkD0j6r
R/sxGrCVTuYS0g4CXDWHTZyc5Ams0jlDCtvPNIY990IEDzU4AnY2r25+km4b5wSvNM/BEnlvueuy
yEk5/1C1BybD8p99Ffax18e7AiduCn8/FaMO5JYBnSadRnob4Rr15w3ugOYcYrdepfs27q1cHUn7
uy4BNqsI7VD75I5NAXXuBbwDCPGcs/OIXTIeeC24SpvYm+ZMaX+IF6QrT/Hps8ackhaddSdb405H
Nc7lv/q3EbsO6nJxuK4AgJm5lufaykz86udeCZkNNt2w0q/fRDnT3OCZzmXPVG1Hn4TV/1MWvdON
c2e6im0nZxM0kExcvnPaVt8z7bZn6kkaD4rMn5f85q6k/lavE0OOT26h1RbXIev/GmzN6KWIeAuF
45n3FON7joIJFfnebV+5LuJ2VU5qcHM2RMHt5qfP0GHwzmrEhSFRzDakJSrOQjOc8+MGWa3EqRCm
foql7XAmEitk13Qf/EQiz7FnH1dmKNd3J4szXWEqG1Gi6V330Rx7qMP2KCxit+Xt2ehAkl963BHo
m8IeNd8T8ysWmjen7xtglncbm54ftdhAPRMIGAQbpLXHtkWLfja0T2XTAJt+tr4c+VbpNj2xMKlq
jiva6/ou8NnurITVMtpq136ZL/KH+P/zQ5FUAArRuv/fRPuWF/vxz2bRPwjuwbFJ/TqLebdN+yI/
I4gb1zSC/GsF4SrMa9kadv+FDg9+MGNP2sbyVaeoJ7NFrh1Qpw9HPus5uhsZ80EPTDcvLbcy41FD
h5oS2lLh23GW0WhiukTAKmNlH+sK+rYwWYTNzSGIxZuGsh/8fhwoY7Gu7+jqS3Kg0iricoxpaS/2
kzJQgLn/Z7ZZRI4vsuqbazsHHyDJdwNJ1RK1u2zkN43fyumCNVA0y7GKuTd7QRl1rxXxJ83LO5gO
25GSjNlBJq5e8lEsL4D86xvx0MM3boMYeHTLp372q19h092yFuOKbgJ7fuU2DeOQhMuRRHpLvDxI
RfV5H61fQg437cvJ0MOBXc7t2fv85esrx9fONGzTM+hyeUX/rm6IPaV8lGYxA3MVxKQ4OvsU7EV7
ESDTyjvEVgPMP0TTfETkw8Im3hC9VvGAY/jWIW3RHaURkoMPSKxVO9Zcv2KrPbRMPl5nhL79NZRx
gQ+eZCyIxEGKFRerEw8zP7reR/8oZpsz6BBD/vIJrX8i0JEbcF6m2l15+J0zgqOH+tzvqop3U0wr
1i8JlPIIElOgsRRhEsEkteQqJ3Q6XizUXKKRSo6Nfvn4ZWrITSX7n2JryJ510sZsCxndVdksDpQ8
Dg2v07+Qkvk8OWO22B/f8STsKbxc9J3IhxfFBkOGMR0kfHbibIIwlHegEbRBIYpmfklkKcWzuh6F
/UBIEwqBlolYzg0T0CJIoU+YmExL1xvE7R5OU4GZ3O9wsm+4P88YWpN/9wxlWzAhyDZo3TcjZarq
pdEYyq2e8Sa7opuYmkP/lXP2fLKsJ46SZL4/eHVjbeEm/H7uwSnuOKSEmqgui8HWD6mcf2RR9v0r
Xd5KQrhrsXqMgAkR/NchbwoFTTSN12mKrG+ds1eVJTy7L/XqaVvgKb6+s0TnIfbqczPvcoYGfLs1
byDiKjIOmBKH5EFmFlGIgioyW8KYeafvvBPVbKZoM9gRyt74bntJVMqHNcGA/v9LsRXhX+s2Hdbn
o59IYAZFwZvGtlo/KZdBNNfSRx86keM3mXrlX0mBSQ8K5t9UlnXOIOcb27nCuywCG1YYw3Fng8fZ
nB9NAnQsXxksTnyUPs1RAPrURFRNZnNLRihz9bZDSM7opTfGed5BGq4tCYbcTqaIC5bL3w9icMtB
ajEO+HfCsw/GIFxDau2OXlCS64BGbnLXowi45CU1f9hULov7E33wwIioMY+72VYizTUY7RLXxJPI
C98XlKze0ClQmAGWyNLTyRrvJMGwKmAbEGS79Tub112w3Mx1OaXupfJs2rUY0qDaapV0wA4DWzEf
7eTKHazPqhDhABl4HrSBkMJ8SpknSg6xY+8WqK4UXuCW/OqZScfXMxNFfVhBDOuUNvuvDBaOuhEY
dwodmzmiXbw6ffvyZZqgSYpPG9D9XoSHbphyuORFcV84oPGuNRSq12w6zf9fO9qiv74dzmnXZhPs
QWEbKcNG+oKezDzbIygw6BIlGpuqUSgapr7etnHWeYmQRu343PTSxN38IQUq5sLR2z41MB/QUKZj
6WqQM3pNNcbWeRzPu4ZEVIhIEMNN/cgwUCBfiDcWVncSMKRhQU4qBeC+KB8m6cK3AIIBl2yAsjGs
SL2T39TmPLY8Uyjszw2F1x5pgH3RYwvB7U00whNue1svlK4nPCB+EElMqPDM1g+1D3rX3nnX0eP3
XH75CgRqvNAoJXcO4QCmTEZh+nQdQ75xXMCVTfyPtb5lodnAaCCAVoNp836y/GT1yvEyDtkf64rR
e72siko4r9Mci6wpWZ8uxWBzMJDJG0w0D8HjWdgADT6TBEcdaY/vlLCFNCiH9rgpj9SYkxRCzoVm
YCA+uySW5iABim1mJLsYjA+HAC8bClzVIVfQjkmusmULP2bYkf746nCIvxqJOqpMlo9CSR1D0wm8
N9JhUtEvlrUpKFH6XcnE1XJRxk8GDcY8zHw2v6w9wyQX/8gZWLH2S72nQtvzpoThZbUpbsku01iv
8tnRq6pac7HZknoPX6Nz5YITvFiJmPga8agK9Q2bDHg4JepIz9ttd/3BAaYC4lCrUciwgirNb151
ydLKjC46G3uBn1CMCzaoAPJDjvk3EeXTY8XNtrNJf2r0G1O+XpSTdcABoPkfTx0A0SbsoDtT6n7Z
ufEQtZtcKh1LXQZUMH1gWIXdVjxI9HaFnSDf77m1clxEeFZGCJbV79ehqNBwr85GE9cbTSfb5Hd7
M6gB6RuILqO1nloN4uAQr0Sv9OOJ/x6IEAzqmaPue6tptD9npnMUWXPpiqTAK7LO/spcZKjS5dVz
+MJWJeXfMmr/2r1Sy1cb8P3Ha/A/jYV2febUmxN+q7RMV1LLM/7+LqJVTMHIT99QW9M6LaAGNkL6
2k4rjjj5jcyYo7oFVfzM3g7PHu3EMofB6KdPCOx76c5dTdpnTaFXmFwbfECjyViwcIII0jg4gIP0
eD69hpoVQCCQwq5pI3TiMdJv2fNz4BMkDorh1hWuj/T8KDuxNT1I6tfFR1b8e13HbU7rP3npHNwK
pB6hcxNw8lKaz7Jx/zgzm6Z6HGzA+aqLqOo1rJXX9ILfczUFw5gEvwlviPddIi8o2/y5j38sltCD
GB0AoWRj21/ScisjrRC/uKraGfRUBF1Hfe6tV19CLs0DDZMV3MopXOxqUda7ewKAb4XTXUw02eI3
TJPJyZBHFBlFep1G9G0mZ4lRQZdFAFelzlKt7v5RZMxdJkNsutmvvanX0hSj8e/ydk2jcOsgN1of
a3w5c0ojagijEX4/VDkgAGZJ43DYxu1o6SGv3a/K2NwQBVjFSHE9w2zZg669xb2UXPyudmYm4Ab9
u0JHFF4dSM0JiiNiErYAeXYJqXRI+NOL7ofTlotJgTn5tTSlg4eIKv1ClaZ7Jr4RB/e6C7FyWLwB
IIgIDyvVlSaF0W45cfbRg5RNm9SMrmKnlIwMbN6T4QEb1aWaxGlWiB2230DTWczkfNN/z4xZsNBo
0UBWsOTDsb6zT6561+Mveo11NOo0P9v/QvFkTV1QGwNYIqV8FfFpRJwbbk3BDqWDLiL6qWpQ97Ru
ZvG8kbXpy8HrXhesMIwfTf/vcgjLRcZJs0QYZMtlDVYMDy2g6x6Rt+72oW9O4q8xIUxzGDK1lTBa
HJj9m2FsH9SFxtdozaoqq+b5BGr1vn5/Ij3iP5LGhoq04Edrp7FXOFZOmlbatC8P24HrsP2kEbmJ
l4ikIeMQ8CcdB6sRVfmm35yooZH9+GJY24qsmdg+BM+hPM6WvnZ3R0+wJszTQxYvYl2lQfzrGAA0
4u46Epir+OuYxQqX6lZ1y6971Q4+9U5uunRo5Z3mWHoxZjFiJO23OVHbputnNIte8grvALA5TWvP
Y6KsnfXnjhF3BpzY+J4ambeTyH460QDaA6f3yl6xxXgXYRyXxOhTZez/n3V3KAHyAUYlrRFA6xo/
+hznInCAMJH1puuwu6lUTDjznZyphjAbE4p0Z4Gx2yU85YuMkfwAkaSwy/DvSGq8IxO3SnQjJ80y
mLAEXBUbSrPDbK7nSH1YEM4AMz3tOmMXKB2UXyAD59GgYwvHivww05pU6vnp/H7J9h6OVlrnNU/j
33lvOqx/H0x25aPcy/3/mWSwmnSQyUb80WWac67t1IX6tKJH4+So7C5S7hjUb87vkSpuPleVQAC2
GNySUstx6u9NsUkKPXfLIs7ucO9nLFhHVF8r8LW93dr9uvbZWJGYUsemgiBqFMAx1g8QAhPBpZIi
6ZVWYmXLvHIHyqRlcilTHhQ/oLHn81HgsTuHaZm5Y3PUAHeZwR8ida/x/fOh67HmdiRUMjIiGRNu
3z0cBHQOYXOoEJQjZN7149qQ8A49fWy/da+Z38doYsMB1Ss+beF16iOc5YVGSf/8rqGxq5pOd3PA
vAKC1FB7lb58En4t9fIIZ6aAiqR1KRmE6TT1FzELfT0Zt5Nmo8KPX0C806zc4C+hB1/5EbfIHcXN
tDI30NEZTscm71pxXGzN7ZncLx8getfZr3PAuntCCg8ZcbdKx5cb35r07b6CVbQmEzoGhuqcKfnL
L5TiYfDKdk1CefQ3v9RaSgz29vEBNUG09J2I/1ykbvVpsxTnXp9jhdu1V/9ci9auUQK6ckJLOLU/
mALQ0KMiFQMXIZUhunVkK9XGPXKAbknKZ1lTb7w/HbzvHF80BnWLTZ3ZTLPmjapLrO6WBgEVLwJH
gTjZjAE9EZzlsdgd/ur6AysZ6aylo/a51/Gi2im6bcOW91JEI0gteF2IptpeHXfgGAYEvO/ioEAR
narTlXASDn4y7p5Ir14KZOPeAM72jaOwtpThTPnnr1n7bqzmwnVNTh+1Xcm+dRydVt6fNLhWRH2g
jm2lvNy2HGXMhGo1FOggLfm3mldMnd4VPMaPc8HZmDR08AKE2QVqGypkAiicrSWYCIq67ZiUGtV1
DXCvqiBbozk1hTf/c4AMLPaYZzOBfME+ei7IOOOLtNaffWJ2qaS1bxsVldhXADamQCKDFxV6aNpB
mSGC3vpVhQB6xNESxrNaKq08vkso/9qtILvacL9mrx0q1PDGMHmTsZI8zS9ov3zZkkmFp0OI3IKV
3/MJf9N57Mt6bqR2usRWtRVdacAksLGF5a6mijZ611xzgw7wNg1Q8dMIvx/Z8cuu7dbwd+1ob9mB
fj0VUBMQu+UwOZqpNqy9aGRkMfUyvsU73LE6DJY/nTA0UEomXlEqDYqGNuyCXraaMCorGGOOZZbE
ualUSgVULd8D+3AAv88X7615lMCPQjfLSNJDtf2+KkB9i0VHpYJqInU4X96JPhqWq9cVhCuOzFMi
75KZZCeshLhRI4NHj+1zxdoqU7bNXo/NuD4aUkAPDxvyhxFUKwXSfIL+vmLQnK/0cex8hkDJuBrb
p3uo6NgSrNuJ74O6J2dpUo07bo3RWgtK3UfJywhwy9AOI5ibeIcPuQP9JQjvjBeI/7wDucvJMn1N
5KKucsMyFlsFhMVwAjPDGm2RgWOp9+FRuSbbFsSU8YF70HjosZalqL6ir61xdYGbeytU0Hh0irrV
qMX4k7lTUMK2g40COuzWm0+3v0hUSE6MIVIdxsHPeYkX1/54xXu+R0vUFslxBOnHuDFNbSehGtWp
uMGdeLCALe4OQ2rb1nMtxmTGWUI3Sppw3Uzl+1+8Ts55QLfspwRpKk9JwQIRCes8dLEhF7qwrgie
BI4evaDntEaGWsJNDR67/t3DSP5pJ8rCxEo7jRTtNqc1hTh3mWcl3uh8elBr3TG/49gpAMmbAnf7
D+sSI7yypSEZ29yOsIn3/ZXTE8o4EP7fjoqI9imDmJkmFBnjpWerC675TdYm7tMDWiY4slgho6Dt
p7gMgETUccJemgsSzZVtAC75shxEPuREUyj8+d044+k3kjGFXayiL9x4LS4iLLM92tfuzBn5kdaA
VSF+KpL3d0LarvUsre/1vA4BARXHa2KjrsFnS95JiiX7ykqXi0ISLQ1bhHZ14aHc5qBP2rzJqdgd
GF13YzcBpNfi5bq0GQB4z8xsjAdtMkaDisB34EAQ4GolNGGzfvT367YofuM6nBv6iypTaeAZ3Oog
+9ydSp88pCgTHNtfD4rIlgUBbdlkfGQsKED+MhqeX67kGL7OzVC9mveK3mipJDpOW8qaJyKiZj+/
u6nKiSMzPXQLkHDkoUnsr015FuMYFJh8dzxRF+s5o+9FO2TI8CTGa5v3qPx9ZB808FUtruWAJtQ3
GG3huoIg4S3GAEHlYZD7GQ8vJAHB8JremK4n9SRlyGKqBvfVXBKD/Iqg02yjLnUIlwHIqQ0cFXhG
bTyGgPo36vzN0kFNsaO6NjpYonRbesNMlDy6TdG5Kg12n8lwDqEhXldL+69sI5QUl9P53qGzziEY
Y7elC+1kLinT3/QFIK5BhnH8WpXxUYTHApZuS8gh4g3jw2eJTEB5++3ccpsyGF9uOYuKTfmM0yYK
DYQ769+FMrLhxCJSXuNip4rRRbpXGdRa1S2tsUUDiHbyF2kDdHs4kMlFAT2ZA1UeWEN5ymRm73uk
qDvM78KTD80A1eT7j3wKKMpDwY0oslMI3q8U8AnkAWCI9f3ngmP5uvabFHmif58g+IC3tqSGR+AP
lbd/XGHgTQyCQAVQ8BAmmx5ECWncSMnjhTqw16ID79sdckJhG3n4dCUaY+xEulJVbameCpRxxYOc
QcuzIu4ZWff9OQ+ubtlUGsYwkN9FBxJNxxCN4AgoC+8tLm91S3/qHVxRSpDPHpViuqi4f5JgS6O/
DQCWwYGr8z0xvUuNY1DtB2mTdo+uiteUNKqMKeEv7QXVTemxlG8jPA9/pbDJv5A8pJwxIYvO3xD6
5xSQygkb4YpRo91RObgD/am2UPOnGvs762O9aA55XBnmrYsilj2T/UPD+NEPueD90dDfVWxwLh5S
fJeHaStts/cE4nkpLz1+302wiSe0tdclEJCL7SDFDs4Dl2x2FZkQNDVL1zmS79IUCMbFVYIERpHc
Kj7PuPp+q2fW6JN7lR8Y0hO6xFZ7qllcSs+zdIgvHzXTHG0cxBuod+r48+XM7R1pFlI+Tv9TRSAr
JwUZi/g7WOqmJQhZoSg5JiUndUeM/X4fR9Mpy4QPxuLBV9QRKDy8i8h47t/cyxH7WHQrGflhONJM
ZEbwd4eQFI4h7fjOKWIqB0riWICTS5XPxiwpPFdBpaQq88tsqBciXYjvUwL8Zv7232In0FOkzv3Y
Eh+GK1QJ18kv2qAyqvYFjSmW5sRfgtmNpBPzmwt862Y3ljUSy15Xaj2vVPXLNmILzoj3l8K9NKEV
x+1pSMeG6WtKaRkrBExavbgiOzSP1vJVs72/5T0rN/7Da2MCJU0uHjl0ReqFi9fNfOpQ8nXEOqAm
fLvIiPY5psMa1H5HuzEnWlQdHaZJb5cQwcSc3hUhIWt8TypYI/xKgXtv9CC6rlOR+tT7DPbASMup
UN0lBj9x37Anxm8tGWmnP55zBDNkMM3Qvzhw1Dj3mCDj9GT7m5GsQjgZLm3wLucb1wlJw3TKsPpb
+bo8zCUShAD8A5IB8qd+feRCLlEK7jsmkDOEudwWgEUABDCmIQ9K/3a7VDENyDoJiaLZ6JKsrYPr
FSChT5skrMQX4aaQiM96n/c+iSs0rXYDs6K03gdL0WRO6ogI9oNSUi9KeUR/lzj6O0IY/cSJuxEj
Cc30TTBVBNJ8/F0DvvOMoc6wgZYT+fTp8M/P5G61RY/i6EJxYWWFtAEKyO6zPxehVr3zvh3mazv6
Twebg7vEZ49pRcFEIlSpFXFo1bOb4hBD0VgT3pMODAgQrhK5vMIVK/Mt8QSbSfW2yYLX8NU2wysy
y54HbsLZwnx0ccAgsXCoUWB9aeymJz25xfkWr40TEmb8JKimmdIF09AwxVrhy1vFg8Ba1OlO1poJ
/5Z596U5MlYXf903Fo2ZKOzyhxfIWsRhNdP/P/sfr94IMGqz0Y09u7/YN2OlfKjUcTNbAHrYtatw
++/Idz06uiexCxKNW9YiD1yAM5ftwtxv5XN++FnmHQvawoCM5a1TKSTGy7J9hn0hZVhWCyF66CgV
spzpiN6GG4AgyOur7Wbw4USLoRKGwmST6f8a+6Pgsnuyie5C08tRnWRg3HvgmCWOSe3J4CHrIk9+
UuhSshwmaeC+XPRAi2g4MHdt682tyRLUQNLK5l++kECryoOG/W2k3Y9ChExieddu/nR0XWoKpOzb
WjCCQWQG9JJNK2RmnwW66P00mWXfG47aSC2ZHhtspMoIQW/KTSpW+7J+0ipq5QzGJczudlbkjIwj
pbqgqNDz68mfM8w+T4ltBsVTtKasElLK4EYKHuomifoq38pSVC0O0ug2Gz05D+IJc9/V2lvUrHPr
d0H7Q4X339iZe0MKKc9fq9pYQEM2NGMYjeH/L7O5pul4UYwm24RgVxt/N2Vop0Epji2R1vAg2DIP
pi+oOlBsM3/VgRUQ9GySSJcOGu2c1yqD3Sa2SbTFTfzkA2lqlCqHQloIiKwK8yEAWo9lvnRT+1GO
BS2WYBv12RUDfGGPCB379IdsVeV5ScjVyXhG8bJBlrYPnurfHZE5Xg64/aM2NGKTpb+KtYc42IDE
asE8zMIuJHZ00afFYoiPMYj7D0FUPPoYx4M1dEJOOQKx0UgrZhlVQxeUxySNdc74ODOZ9ZQ3B+bk
300J1aBmxVB6gNOUCKIDqSFMZNkLnVyiJivh93xBfwnaA26QQxOjZmLXYyjgnjouapZmR2EJJEKJ
CidwAs8tO6lNG20hoi77YRnFBKmA0p7odUxBdLL72I6SPaRxcifD4Dag2u9SZEYTuKnORCbgIqFr
si/DLg6TdY2OvAPJrIiIV0iszrarI827TDwFOeTX435cPDVUhSv7ItLv+qb8Na6nOhumEI8pBuAj
kgeUmeoAnoVwjL6d4cPctKcjNSBvcdhWNvvmrIkgkItt4o1bf0+KgC9ijAcbo5KdS/s5NrUAyvm+
YYvEQgi++V7mPI3l63/UPrvzL4MsU3xW9Np65Ol86HN1YbRJuyCmdDfI2gIQ7+pPvCdgt5GrHXdq
Df8AT5tCgYVqBFLhs/4ce+SCgWcFO1AQh4Ef3UnfPDJrnCHuf1gUYnOWDnW1lCBEUspw2A4AIEyW
YzTQQQUH7bEvP8TpLM/kMHyZGs4qW+dqiPl3lzwt28xIdY6F3jRhl8tHuynZLnh//7LwbQj61Pp2
yq4cWUCJpQ3r9sQat+TNBKdwF/d0EEclOpwS1ab3IzaND6ZtvmBss3xcO/kvF8iTibA2mQ1htyln
v3IqblzdW7TGVtS0aOXE7aAtcKEB1/P9klNFib5Eeydm7eU/LrAYt0iFNKKcr7OeNK/0LcOk0QXh
+DjwQ6cPB8b3278I6rwOK+Xrxi1KMG0aEYzdHBE1YFXiU5dhUKrxwE8hFtRyblr4VNcaptG3cpq9
mx4XEMRTo8WVEytPpRk9Mvj+2myiu7dSXLTGIoXJ0IsEfN0Rdx4xyiBZMs0w1NbRiPhojuQsmj0H
YBrqTXg0rO7rS2+BQgr+E1OTQ6YTkH5NxbwfjEM1qu/g4DvWp7oS7qMQ9dKD9vWCIdDVjNKlXZC9
+RiwOtkyuzx8/Rsd6IvjF/eR1PM+Mr+DZFR7vtzivLCFXO0jZlvW55+nKmKM/n8Y4m2xdI5T+hFu
0rVI3LXC3pBrsHiVfJwb/huTsd1CrwjXOsadtOoQdNvEAQZhxjT4ZxBeENHA39ihg2sU8X3gT/nR
7WAZCd4Ht1RJ7kzhd39j+xjvKUpwzeBgGJIMPNiLsvi6adH/TK6ti7SKLgtMOV8Ulj3n1ywI0AN7
yKq3h9sBZKidceFjOyLKRkCDeUBWF0p5ARD/sf31HP5Wk0NJq5Vrjb3SoTlIXUYEXdIZGokls49w
EEkz3yde7fbRLOzOcy6GRCXWr+s72VutCea5QzjVtTjdtzh3+1BKkDIFgSsZ1VkFJM7NzH53h7NU
ZEz7PfRsE547cukOweYVJK9heoaItCN0m0ArM4w7FhdQEfxrTA0jvwXY83jdrM5bJFRR7Yj7+jkV
46fh8AyyROzBDqDCFnwiMDoZowYDGmOhzSpaD/h6LYHZ1CcRKvjDfWQRueCyiUsRXEaBI7vGZ7p1
FLveUzpzMA0MXvXI5ztTFWbCArpyud6KSk9GFcezkH588NW2MRkg+59/ZAPG/VaElFyjE0alwZb7
M+e6IBqgEjXDfaFdTLVbAr9hKmZ/zwdy3cNjL20c5cpGRNs2tePehCW/dKwqFih8iZyFw09R6Ngz
CLum+C3tIQD/pK5kfTfT6v6rNJQqsXA4PZiF1NV6+fu1my/4ZAqEsIqNz17lcxQbjC6yqKEyfP0L
e8VOPNWskypKYUu1kecLjoUfugMS9s9hAzL7PXWaQggu0KxR/3+ztlH+6IjLatpOB1nfNW6xmnPa
aDEP6+K+PcWPlC/J75BMlKMautpYiwXkD6kVuMuGOWuOrfbIN9WZPpEoF2Z6p7dCBDho+Lae16la
VQMfo4bh/YPFk5RM+u5+xA3bidDwlq5/zVrT1I28TweYSM79TAUm12S0CRpUbBeKJB0XXB+UL+b7
0qCKTKhlRSQFCUecQPPhCx0WQ59LBPdIjroH/cEATVb/cw4B5OTzTu5pVZopIBhh3nTEv1+FXDh4
YE/EcPqegFWLKd4Hotxs6DGb1QMM5VRS+lq/DKhbraaxgaEJ1i2z5yVLUdrDNMsvE+jnd9h3stIz
c9j/qvzPV0acandFX3ue7OmrHFYWoHUtuVxJJ3+Ph2HC0zXP6F8eHFXzT3gNtKxhdnC2+tNtIvvN
wsNu/iYbgkqaZjD2hiIS9PicFMMKaJiDdkk0PQu0f8Frr3BU860EeZ0o4SSOcNfGJAMic9/Bqa7T
wcoLJh8d7WgKRdhoR0G67/ve9cbShBzngO3e9nnt7JM2NLv94bOQYUHBHbdcFoKOjI1TqhH8YXlR
p1zWn1vOGHf+5zRYkW8pYryFmiGDNoIEYGlyjQH65hvrSp/PK/XMaxuk50lcEhGUwvL0/JG4ZlvQ
t+nc9csGJ4oU2ty6O8yEXY6HjutwVjJShy9BVaaw0VWpd8K2YvZW4r2NGU/IbsE+JaQLNSb5xxMv
fUzhtbhdDHc1U1eCERFecG7L8xsBjMQhW9hKVwlY5uaS+J2UKrkoXjYYoHXCoPLoXd6m/Ez3sow/
3MOm31FwpkdLU97qBCb+I+GlHi1sFta9YDpYeunBBjqVh79Q+7dbgPDVxTcP0cl37mbC3M47UqJo
N9nHLjv8/nt3MPb1xlY7LvbWW03cJmi6nrFU4ZYcA8d5/OWyXaqLvkHXed5MyOcPzNH567u/Y/O5
OEHU/jgA8S/+r3DwNaR0/Uuwpk4ekW4yCAfAbQgB6q/nJ8LbTV/MeKkPxXEqZt8ct0+95g3IhHgu
IRFnIcTEfHdXbMaSjkbnXiImkYljMsEynihueCeK/oQBZwKj1adrd2cwQI4XgSOaWFnytjSWXltW
Emhv50XJDK2EmbbaEIy7iOZrUA+d729cPkmgxtnv1qRmZQi58y+6W2urVnEqpAd9grALJNBIebiv
/5s3vgJWCAaJETfVSDxTtFOpsdy4aBoK7iq2VaT7vJKPvfC9dCwmP+yEJAIvTLbaYH97aUV38rhA
AcoqtZpE1A9zxUZC5EesvizHha0mTiiyMYOFI/MGdO5mUBrJSFQ5d06YiWx6gsreg81hB+lkfqvI
J5DiaKxrEgnOAOlv+zc0WlgcXCT+uukCwcP3UEcZBN8rT0+wUOzQlKjXjs4QId0yLKK05U3AYoPu
yGX5z3cmjrLsxh4x1qHXmgSf+ocS17342pf/biNeuphIXx0Lej5v1lNiWL/HgI2lAI543xCIl0eT
BfoC1QYcxReEWf8QkrQ1TzQ4iMY2sxhzf0P12E/uUoIeVhqgYBSDNkvUGS1hLKc8nhtbZs0YZTy7
TVGnGYhqVD4gPPEgxsZTr8P6vQ7B5LNY1ygTnVR3izm/DPcyQLjt9fqhtFhf4l8gaew1BPy060Nr
ix2uZlMa961TS2BLKRUBgcct4p0ptvmvdV/Ulei2vkc/+ImdExgD3kiwNfX9NZljJu71mK/rDHip
JqcBoC6agbAz1hB3VVUOCKCURu2lwXfJp44hUHdAq0cPny0mJOJLxrT3J+exytMZclYN/bBhH1AP
D8BvHOHXXjC2V2Bpb1OCdeRhifgmHa6u1RT8YRMdZtX5i7lNXoX2OZRZ74yGFcefnfEU/W9DLalP
vkfpuMUebOVcc9ZkIUn/dF1Pa8kkbkg70xUe7gkyaSYdYF6rm6EOQMnBRThSyDpImxqmikChZUv/
CQu95/s8zbekrKFsoxneACKh/LZW1kkUdd5pzno1UH9vJqB2Uz7NB+qk2V/1oLPEmeenPQJq07gN
qCJ+tdkCN5NTCHcJyz/pFRUYskjFbVfGUFmJ3ehGvDiuDUyYDyN9fOWHexILJjemI7pA4I8CYfQn
pPUJM6dEYkHLnxTbKfQQe85J2/76+LK+Sz4Ft4tcIMvl9MgijOeWjioDckxpED8VdCXsvPHJEVgq
fsdn3Am+AO9ZQ3z0uOV4wEkYv9nwD0/TtYUWrsBgdGqcT9emSocGccRKEi0ncn4fsvyoUxtUkJlE
RSFT+RHzK871imTHIW51L3XKOD7Uz6M46Ro1pP5XO8z0OgGmBWnGsIZXDX/gRw4WjvNOoT1DMMPV
tNbhpk8KWlKd+hqJF6CBKG+eoZ+GKHFj7i3i7Sl/0da9BDrhCAecsxrckEuz3A74Z7xzS0dsOvVo
fkgThTa3O8cobZzhfHL7AqOJQ2jpW/Ioq2EnF/slmPRJF1iNkwmYyXQPtgtwUoGJrEwIa1zVAI+F
3QgS0sUmI0SjWgCYRbuIcvCEx5cpm4bkLvPTSZQabrCltUdQGl2ThizRztWeylnr4YEbwJs60yWH
LagWfLlSbA2IozQcyFRSYamLElWaWl44p5VgaKzswloTiYysy04BToL6XIDfvHchfvs8D7kkLqbn
u2hhd3HCGMgHp2H+sZcdBDnF7s4tuJUYVAkS4EPQ54QrzFAmmOt12Jq/Q3YUfETEognZbyK5NYX+
KbWBGYeo/VanTdyDy446KGcuKtvpSAoZerilM5dpaqFOQcv61ac2pbPsHIhnVWgSa1Oo1nmgUjfQ
l2NryHM6lquf49i+dTDDP+VAYa0D2sB7AHpWk3ifEpyClrTFTEoUZeWJuSS82J1QK0A/6VP1bIEJ
k3wB60131h6d7/Vt4bm47waNup2BDHQEENQ6ljrGUbWHL0Z0cNaJVYiZDe2lKjYO9f5kFbOKzKiY
zriSg4vwE6C9K31tGtS6lEgyR8oXjHoprpoT+EMkd6sIPlv3kOStxTfK6hDugCj9XjpgrC/FMgg9
y989pllQcVmQtp+qE/FLj4GBuhRgVYXAEZK7HwSRUC52WRVFNhpiX/ATPxm1/3hJyoEy2tjA+n/h
mVUgYj5RylKNc9FBjYQwg/BMZBWGAgzGjN1u6NZYTTjWTPwRO/Lqrm6k1swOLMgsYwa5XMNyy2aj
FKoCm1dSXUqioXlR704nEMG25co6oys12ExpzrRlHTVjq7kaUf3J7TZcI35AHHSq54LS86PIRdTX
bVjFmXj3Gaj17Vu5rcpaY64b5KRq725DE135fQJ0C5PDOagUbCSUpl6MLqVaqRXC3oqCwMD0IIDQ
92q/j0ScwokRluK1ECj3LFPBB1PKfPPoho1rWI8108ORhjnTp2318K9cATUlxS7BGUiDb28BNlJC
RrL+T/uEaDB/NnShDWpYyV6Ikxr1EMtVmUE2/fA4Jyma3y4Ialnlyy4BXHRpffCjYXbbKEXkFmiM
PNFsXPMB6xWwepk3kGcweHqah+EkwkjeArgKzG26XZ+qjiVe0UyOA5cQfmWrolEEdwZpH3M0xLVb
KIP8JnWLZ5jzKBoMxiuj3XK0k4+GqvH1NPjfYBxweZIdICfX0g1bgdJrXfYtk3jfazRJWPqsLGci
TNhQamPBZa8hMRRytgoxmiqYGU0/5UTLF2pI3bVXsPJmyTBStkN24pDmptvDi7CHx3VYaHdKuc6m
KssBNNLnmpsDMVQSYQmoSPIQF+U6q2/8BJY0svwGVbrfAkh8jTohdezXw8ep4Op+/TvjQwr/YWpj
2E6Q/CxUK5e4wQ6r58AhX+bY1STOLOROyzmm/Se+6S8xy/3p7cQw/99elN3s0q0HjVj3e2ORXbnV
oRlpAE5PgMHM1SR6swJj28k12Q7Q8xEOz5m8g5LfaYHdImEIDduVYGDhGwzbwEPCvLwNyVFWnDP8
s8My+ZgLQdnJAOse/dGMEXrovEMCMHC5NzidPA21p1fA1kQlN7Jg/p4DTjdRXYU4xmqNdBArL3sm
cSYHK7om6cFdDajjn9kqHZNB//zskeJaf1l3QGlAUtWVod3zuit/xsWQYQiTFowTawAYKuowD8JM
ezKb+a+BrBfHXZvtP6xa1OyOGUjuJt/Dy8E9ezWblrmuBi/HSr6RszoKiwW0kFFltQbsVGJ8DDXM
/ApsMkABkj6n3FzaYm+o7Gn73lbtSHn233aomzW41UtSP22CCjevcjsViWF6axtw8wz5I7BzUvbc
Rdmx83Vo0WLIys8MAzNdsfEkptF4ykpPr+5MKdH9xbidNvnct6AKrLn6BNGyd9o1/e9S9Zd+yrKo
U3LTHDsbKBrII4ZVizV5zzUBIiCwx9aeqgqmY/adn3Pd+k2uQ9XIYX/K6cII4hEdPCgvF+E93WEu
AkWufeRPUmD17eKhOfdD98tTDXQKRGHhAvudZFV3JKLHJy/I9WpY4ERITwNMUZTOXgcgdrfHmsE/
LzzhXzoPMH1OE64GI7GuGBKg8EgCxfaEQyygS5BhwSrRNkAFwq1yy1J1fWSPiD7VSGlowt0dpXmQ
yWzFEpBl4IHDAs6Tu0G3uHymsSLl50QT0VnWVK7ufKQxcwvM0UlhwKXqs2sqOffLAtjh+XjIokY7
YxbbLRH1h5fTmdR2ukIv7LQbzc2LEU3j88w1WIZ064GMYT+mH9wgfS7i2YrR3V9nr2LlVFI8bqDP
Wks5OP8JgoLUubO81xHiiEKx64yaNSiUMuJNpuGvR0JdANH9yzdKovgiXSTMf9dz9snrQMo31wvJ
Ky45nAw5hS7PUWHlUqi+rsCKLRfD76k/0niy4i0CubPDZxZ9cdLXaFrZ2zRr8xbNBgBmwHljwzFn
nFA4gBa/qJJiqFlB5gj9E8fycxGhqVeAp0cALw/7/Zlm/QHZIHzTUPu/59DtwsGCmM7zBbskNvIn
2+9zK+BnSo+nQLen+erC3RcyKyBlIw11+QzVr2cWyxgEcOdsWqwrlrqzpHgnRrIZMkuPIdO4OZkj
7nhSvyaifEoH4yei8mPdLKhZC9NVYYAx1pNMDbADhobBgFFyhfMpPyVRB2ZSuMqirbYxpLggWXrM
U3mB1RRwqOK7KygFlI1iPDHoDDWnUI2VozaBOk/gI8yeAt5hKIF35Drr8DnNF9vpOocZ71I0iYYL
LBdZMJb9GEuwR0b+Ha2mebpnN/EM4NhLzjsjOenrqk7OUftAn0mhQ8DXU+oWr8foD2j4hGnRGWwU
1W8dFfZnpjFbGZJZGaxZEtFg3h1OoFSJ++3t9n2iyJcRwWlH2BUAUvwp1WtcY7Ww1R0zWR0Mq/vJ
ZekRXJu0XQyawxmuZQwkVeCPv5/LmjeaM0LfhmbiuXCSD8faGVKjWgRBsluj3LYiBUOArxaI5jIw
orft6PQcIRTg/v6E/MKJ52FwDWLov+bY54vOXqeO/aH2q9KkYnPOxqOaEZtPwQk3Fila9tuqiAVY
qkeq8TT7Hzkf7SGepWxsnrdCHmMFz0y++7WjFuXig76b53E+TbhHdHsYODeKc4+nnA/7SQ+3LkR8
YW24FoQkxCezgJsVzmBCW4LTboQpQ89GT5MQzis3Bdx4MUjr9xmvHrSykxJIIlZcS1/ILhBpIZ9L
5iCRCi0VX99IO9Gafd0uHN7yQNtT4Y04S3iuJhwdys6QwJwkAFHJOS9ngXv+1XPmkmcEkhVxaNwY
qKjNSWHCF3gCcPKj4gq9Yhz92i7KyUj2Ay71drgmMIgqDZFivqRl03OnWeGY13qr3uvf+/V7MZVN
zphKgK+cQECY9++e6f4p3KrVDB/xSFwd8BPCAAhZQQXtoq0x8dbueKZqbdSo9bqjh/b8R6cG3x5G
Tdygubn9YmamaFuV/9QHQ3FIoGWQ/2jgUnb0Det7jBOkTXh1aUVUzhWJM1V1qDDJ9LhJ+Ng0q1Bp
Lm5OOqRhE2EE3dgx6ttvLS04kvECSTt5z9U55Pg5hr0D3ukXO65zcIDAFLaMiEXPaUZsxJoFsCDZ
WprcS379TZRf00cGvRx32gGKs5EfvsqgCNSXWYoT/GgJ5ylN9whMXFCB7TFdomIqvkNHtowRyufw
T2Lm8FLkYivdUyLcJUq1cVuomgPTVvyKOfLqCdQMmoXZUSbEbfJJGjiHT38NCvPZsOq3HtNRPLtU
b7hakR/JHUsE1Jva+dZYLGUXjYBMtHT9zmVygpTKEZq7XXXyp3pByluzWT4Z3yJO7Zm9E7E6lR0V
dx/NI0BgphdNJsx9CsZjIGOQbpGoNKCyo+74xhIsLHqBhRD2FmetoPVfuszHf2dHapgawVj54uzw
6woV1GyGiIMsgcgFn+HI39bLz23fA10CldZUYPAqbs5YxXFpN/UmDKOp5vagR9iewo77v1AMkdEE
NlEf1Xp1iPU3eT4U1dAC2KPrvl2m+FFiXAF87X+vsXOhyjaVJnGy63AaOfxVMaboe/rO5ilyArFi
sEFvSKNwrgfHg9YmQw0h3Ure8WSnc9wA0TCynC400Kvwc8Dkt1rnKlDh1IP3kVJ/Lm1aQrjxydFZ
6KPSzKDRhg9FzvQvmvmVjK/YdOI4d0DEPAj0FE7suY0eidLg6OnWjQ5BI1Amlw+YSGYesv6TRlGW
BNLkRFLGlW33fKQ40y+XbhG+gEEq1REwuD/IZ+ofNrUAWBX6IdEWoMO4qnethj6fpkXAyQshTeUM
T1Xzw/AkVtfDI1qQiZHQh9aHO+jNsE88Xik5SQMc/GnPtN155BLQe035zoI32horVK1Xm8XI5tTF
8wdEs0gR0XBkDl28glQ6SaYrUZMiQ2a2vn7pobe0q/lKlPAMjOmPudGFpjjRRiuMJkJDjQ8WvGIU
zo8iEVf0Xml933Re4huoC0XI3+I7eN7S3PO2Db3AgxqG+8Gmn2H6W5q8GJpRr/YcpfnUsq6gnzRH
Dr7OPJ8Um1F2pnS+iLzy9XqvG0J/X5KaoGJoStEFgTETE4lafsN6pANUDwN0wK7Je1VVAx3gkNtt
6KC57qzyDHQlsOPww1L/qov4n4Nm/ZiQKa4XNmSLr/RSCiVQDf45OVCZLr4fqI3DwM+aCo7mnVoD
GwCFavvFqIWSLaesnmsbcGDkL/ttNk7PCP4mF0mKzpHyYlZ1OxYDARb6leA+bMq+5baFFf/Z7wR2
KjOiACISZzXMlsxRXUQWYT9IQXoeqaMbAZ+dEDMhnJ0Lo1t8J1HeGq9wbOX3ktjz1IHlqpc8ZZiG
L3jFj36iMfcNDZkLzMaECBqG6kpSHuZN16ByRgpoy3c+0NKqaBZftDSvlTr2FiAXJVrqnFsyPKpq
oqwmoek8gvM63z3voUkbdPhEePJGOpeAlFsq/NtpMy+WJB1ZWLaal/QzamqNqWmUK9csvECf3+qg
uduJKwB82vRllS3RV146urgl7suPk4Me+pxf2wZ1Gs7M6FeGJ/BpLVk1OT6vZENEOFLvKqfLL1yD
wKpOVCU/qD/p4sWvwWh+z0QDULZmj0PITfICZDz+bqvHCdCSIOjS//ahXkJf85L3+DwC4XNJA8G3
HN2hO4bds0dj4wZvbXBo7+6YsdVdIMcQjmaZ+wQtm4QPPVmlQg3Q404vNuUXWfGAIpMDv6KnAo93
gBekvgLmUh/TfPSM3GxCmXJuZcRtVbEmTB2lPNrIXflDY7VUK3qitrmr7pvCgjVmfj7dKiYb2Pro
wyclZfaiIZPN9IQ2+mo3xzSpsJFgpe2nwY5Q+aBvAqI4rTkV8xCQfx7tWHlfe50sn8288PULa6Pg
CSzdlpziWqwAicUsbuPrp5bJJ+FaGGDTsCghyLwtvbWdn5cVbYWvW6sdWUadWMeIhjesdio6ON1Q
5r3q5XJxBCetCz7SktgN8d0uOw80jMySMFalSJeqsPEjR1g1sjk2mVSr/gPgYC8lBUJ+a80zuYYb
6T8sMd5xVsBAH+n31asN2PfH1vDRVf6JgMJ1I13Lbl/O1W2nIqLYbSSws1SnMG4beRGz6q3hZosZ
sLcsrC266/pfOLc5Aqf10h3DzO7Ja3MtE6K7QvPOwn5Aq52mSYlAFBbwx53XLCRP2j8ogf9k8zcR
e0q5nxLKqFpclHiTUZ5QzItMvQQXgGT7uR9KarJiXUhU+pUnPkscyWqpiAEKMgeEBK7GkmKHRZ8I
qB2rX7bKQ+vYhe8Y5/ewXDbBiKINNCzxPPV1foPxnQbI7WpunelW5Euov+pC6QdVNckK8xUuuJDb
LqPqxhVAZUfPFVNv7tfapLt/ZCEpzl2wgo3ehZpHjeDf+6hki3HjYPD9+VwQAKeFlGqhgr0fp+tw
sox/ObmF+y/m7k7ibjsfJ0ES5e9Sv0LdcmS7Kf2kZ9nVi5c8+dn1jtbGx761tdcdH8Xq6xESlgTI
XOfH43gYVgu9HtBjwH8ZjS0fOoPjYNjsGcO8ISk/DqfHHk6pTLujnzLwgqxreRij63+FdmhE2djO
cpZHwq4MvUAI0sOLj3m1SnbRVE0BaP29GQgkg4kpnQDxGl0KqLOohkazLLG8+c0pLjPaMT0sUzKp
w0L7r5VTzxEw+V3cPaX3gNPT7zBCg3ISTLSL27Ptrwh3PrM9yuENLGakc+S2PYV7Eex7yuSxiIKX
RD1K0ijg1AZM44A8awE10LBWNOykhgA8DCuwGpyAJsqcW3szLVnPET+SLLtPqQbtNJaUadmbHEhT
xdk5z70PEUgh56uxsmGln5z9jEha7VHiAsIHEcM28Klb6nQDr6t90XIQh3X2qpIXjrtDWj3UKT63
5qpDs2tYyb1B4m1H1n96uqgwDgDtnA7tKOu/WTAjIhED/65zkiNoF/2BNy9fqIJpEVPavioK3iLt
OJslht1H303DnjSrI8icxWWHHdfkeaLYiRKyBgfQxBchMWDxk+r2thLLeEkcmh0h1xSt08t2rmEL
jcIUCWea5LzPCYPQ5dnYkq8hSMCYt7z4LjoCtn0tF4TUMI3QquUdTygeaOaA377WeGyDY7+/wc5j
8hPAZLAMjJgZubiVNdHd/4Hm+3xrbNESUX3ffdJjE60NeZuqcApflt6DV8moxiAhBKxKwwY3pfRw
5JbgVNmLYxRhKBTwzjKDPRLaZvIrtNqqdec4WoRr1GU94ejcn+bM+7k2gCSnboTY3s9J/q7bmdjE
MTIYXJtd9/asZI+2s0Cp2BHfE9jWPfbcYrId4pHv08N2oQP2y2EEX1mV5FT6DsUR1xhJuHa5eSer
lwvRXpdNGvMps5EZqWHmzKGtPVSD3W96un3ueXZJrjVZ6M9dKE/tUnY8W+nshQBhE2YVuzlMIio+
pzXzxzaDClKeExoJ5ruvKSmAsLC5JyPRlcBsHCtGKRPvXJ7pHcu7UmEOU4YSw5RmWbuR32txEIfA
rAWwwqkiAC3qZZMEWYRNjqLOa/nxpwEXQKxFEg/hTOUEa5bTYpfXjqlspqHQLXhkiDjx+HVPr/RG
c6x85k1AKLqrgOIRnxZ3VtCKKOiZIBlFXLHjL2w3XDWfbGeG57uCOnlmrr0M8CnpomiTnBW8mOU+
/aRRVyU3IGQ4il4iwBbbMCiyRulujfhrV6OapB+ywtgHzRuGB67LMjKTT5EuV558L05pV2K5YkDB
tvd+EPFwOYBKYtNeftzUjVhRtthy9jsR2/Bln58n2BP+CXlG4Jq90i/CPBkwmKw9Ii9QIfcuKQle
c/plLXSxmpzBhmi8zdlfsbLjcnU6wndWtF5ICelfVsDE5dsgpsZf+udUfUaELcn6RojrEVmEsOs0
GiPLb5NYD/jXrB2ZvTfZSXg9rW/QvW+59GWVLFinTJHb53nRcevBTNih6rRDsmokPJ+7JpFQK9Mm
0PY811vNVPe8Jeh8+YlIiYF2yEnaP3rb6XJbeo69XaxxoDqlSPOFD7Mex82KqlWCIjAXbHLNfglu
phK6FU7p9zLT+3RTdewO7/l04pRW2lPJ99ZDfytTxZc5231s9lEeVH3/0Cvhj6boIsPk7HfICXIJ
y0UZOZ0U1MjJYwqsFHJuk+EfVqYvQRmOYKnJrzPpZuA51bz15FzBunpDchca+WOj0DLkRu0fDu6v
ftoOMAXEUiaD9DDHHqeKML9Hk6ERki5slVb7rC8eQaVk+CgAMuKRZq/FyU+PuYCPzQeOpK3Lb4zL
xLX/SkbgNDAUg02sQcxrKLb/gXq3wk8zi1nV432CjAvxjByHO+gffvJNg0MvpX/fVjpZHdX6nUJu
+NFfCzGceKJUhN6rMt50zuuMpIbD0qrsBzmlaDHumYIPb1pxGPqAECIMhcY/WgJBGdtaZTZzbGdv
dByCpcoYOtNUyUB5rHfdIKqpeCwrRpQLj7KRnijcQtnuq2wzoz2EsrUN6YGjYMovB/6La8oS9TdV
NDkDZXGhoqa0JZGTHj3KxWS4FmXSGVKgbli9kM2ID9j/nXc2gWk5e9S7SO174zVPpb4So0rBxK9L
t/HRRq+VCP4QNngIZKxWBao4qtYXe6/Y2eIbSfyRJrvELV9Spvoe/OTRYxWGWoZ3zCDseuLShjVm
WZlv+WegpZqgEfB0l8AYWoJcAYdv9IYPePM1EqWTDkoYWTmigls7TaFzussxu0uY3o/eRqqtJAAV
uMPtab5ZaIgXhj8eXxniCH3gyuJmcUSdmSlYYZ7Cs2s9zXA5WwrCV2Kfz2oXR6eX/g/02TSm7vrb
i0TNeqs2R1zsgIkhdmNavTV7nkUCedXG7KzML87HfCFNzD+AoNwbEHGfIXVZ7Vnpo9gUdZb9LU0g
oqoxiCyONRnnyv5vdxLDKmdADzc9zRClJ8128jamPTrq3QXCje4DziKsJK2gREVg+FAq9sK73Kx5
GAhMLulQZnS+uxQBo76f5afF+9V3I3ewpOIEbu0Ex2F6GgV95zK8UeBrz0EabooWzckdVCt+Vm0C
axeRodu10BvdaEJEWTozoZBUhK9GUC4wb0S7BPbZOKJy2yz5rC77DSgqG40AUDFJJ0FA0jwJ870N
f62ekGvWP0HSUDi/OqMMZQ1y+ACnaMbONd1wr4EGhNumTFc2m+DmkjEEEph+Z1eMIMODeMM4RfjR
yowIfaZS4/48CRuZH6ge3zVC0B1MZiuuvfSnpIrhoKtW4ID6ZwEZfHVQXio8MDMgqjXZo7aS2Hmp
oqnSeQvTASTEXDnEX/UWeO4S5AZZSBTIIWX9junKoBc4J4FQO/Sry8H4okAAZmmRlBo6x2zyY0eP
0iwRxJhhnu8UonJm1uOsBMQN9491JL2cAH/1DLDqC4rhXKyeJ0KKzKtx1GuLbRTlUzEHgpk4Ub9y
cc/nSepBq7tgPkieyPsy0zUG8qr2HSn2N5WYEHe70MsaHYbTfmjhvrhjPUH9bZB3/R8J1F1JTPTW
62FI7QKxOzjK6656BfVF1lKlaN3icRsKJ6ZCFf6aX9CxJy6a0frixJv7I3sCg+K339PR6Jc/rn1t
2GNHjBSp9N7eMVWNAgwVub+fTMNWtctYU8yu0C7PUYZXT3I6DcDZuQLixTpaZg3ssPhUyI8TTBUh
VzUNbJBu+bRYSsFNuYYbbuXK8sXYkvS/uVjb+A8+5Bs240PCUxJvhAPLG1Ip/WEVy8MGnao0Z2Nn
jplKgJ6Vt4ystbwWW8iLTPeFv8oPwoytIgguS1PmCYm4CvXYvZ+wynfISLTUdz48B7rohDOtx9gd
wwCbYQZ3aapYJfjGyZ1qMc8Xa/7zmKG1pi1JjMgrmKxUGTSE6JivWXM/E0B34eVeud1CD6RCsdEW
2DeGsmedoAEsDc4U2M+8qa9b5EjfbCcmTrVe5iAS/yC1A9tzjgNIe3aUMpUbGb09HXdysXN78VV6
k8cNQYfIQsbpjx4BBmUOCNEZm66W+Y1JRPmgYqcosuIKu3dEjf3ZstnLsRWR3QqHw5UQ91SxdtUy
JOjdOx4B0ChZfWBCYUD5C/uhRYnYqn0aCIyDSt32kSB6uC1tklBBNQhQbDtekYjqIrqfdJ05lbu1
CwsabXo/VGa04QOXjAH+93qUsglulSI2ch7YhX+GtpPxGnLKlefNUrTe5P7eZYgadMT8fe4uj0fV
CqFwW9FTwT1EtXe4PHIL7/v3JkCTVxTNWIB52njSSaXX+Kaq3MyyHgxRtr9nf51RDfijEYnXntFT
5WV9X2sgazr5c/q1uz3GH7n2+C1j8SXCN1kALBB/xZ68HWpvw4DnE7d1tzeOLcMMwrzf0DAcs0gw
SS+GOi3B3cWkpB9C1DjYIjhblQPIM4LQhTltxkR+9xKCE973wuIJpwd73mPWErKQekiHl82Iw5WM
ddmviJCd4TEknHqnPWECL9cxs7IKiLDcJcMdMKCgnmmHKX3bUY4uFn1ndEA4hvuBZIrgVGhnPJ0v
KIqcj0bQSDgbdv+h2tQok/SejCh6ZR8iT7RRNthDvjnO/hzAshqzBOj84FCUPMAL/WfhJae1cFkr
4jVDI+J6ifgnU/H6t1paB4XgEIcdxO8Nl8Yibvd6CUKKtD19DrFbkiwKtrs98EPyd1xMY4CNZ3mw
fuw8Z0y4o37Bdgrwip6hFGj4HadO+BGlhVaPOjsnL/FKjSG+pPBqj7KHFCVNWEuoP3ygdRoZdoCU
McQTRiqSoYmAuhZSFahlcZKv7CghZpTTBguCR3/lASPpSfyLcceNiQBpewhoeeH668MXfMTvxJqF
GeOkVCirXdGBkFVNUm+1mcQ6bWKuJKe9229gj7tz0DC+bmgKRxDspL9Xa/oNCJtn1Fuyx9iVnABD
vxIu5Tty473ED4ypIVcX4ef+H+E/ApPEgrHdl15WiSZ3/3cS49Bl5qZLneoEH3LQnagtg2zd1iu+
sCZwmXKmO+OxANfQQXaTLLydn9rmTk1MuptJooKXnExUd/rQZD1PfpnCiYUjtqgpGr0H9kkDMQ5f
SJjvG1ChZ7kPgS9bc8lPpEp+Ad6eVwKf/WD4lR3BMZhmH3+sLLnIaTOW2w+n98OqnBZoN167tHaD
PvpjVdHB3VYWd9NcKTmNoK2phRCP91CD/DnDFY2KiZVL6n08oRE/Ls7UWF1c9yTweH4n0IzXJRsj
Uaive4jeFGEd0qCu0Niw7b/QQm8jwZL/aEl5WD5t6WpzOO2+iolFPEivqeyy3D2Cq4hKKHvh3XO/
Iq48j2k7s1xET0e57zxd9u/a4KvL6bXtrdQrt67HiMDcUZM2vG7tgbJm/lleu9/Wm9W0UZkbvKrW
FodLafgu1H+56TCo4ByxxtFqwf/CJgfnvZM5fZuO/nC/U+5SfG+0GCv2wSJCsjJrxFfxbiWJqzBY
Aoyn+dei9+tviKfC0tJISzaI6WPubnP1QFY8ffB7NtI3XMpjfnR7jOF5lhlNyG4C63irEkb8Bu91
jpy5yqpTmDjTOqvd7YhuZ44wAVXkAcZwK1vSlx5gwM6AxUGWNqNegZcw6q4MQLTDed/Hw8w+uxdA
vP0+co4Us+1SyOeKtS5o8X22tzT9m0YtEchK1XDiY+MjsiRDZaUK2yhdxHVgw7CXmlbq15or3E8/
oo0RI0exuFjzJS0ZVTEpo0ws+sXO5nFjSDphLy7IV0mdY9YRVvVGCdYW0gBywgtMvdJ36QFHV/TL
g65Hl1cud8ic2tTkHSZqx8cmHgHu1i/jn+GZXfaIChFVGmFgcXiF2i0xUVMYiOqZGmZ5XUakekaG
NPGCh/rDArNclKgdAzfIAPXU9NxPSjjLzYendzH67OkwOTRak9PvqoDS0RBvQJIgrWvFg2zv98Y1
FyU4g1NlNew7J8UpFU6U5AyB/9MisGaqhkyOV1F8jxP8eiSEw1OMdSi05QPbUYubrtEigjHhgJDv
RWLM1tlUgZJqKyDIAwWgrR4pvPAq/e8h2fg/mu8biobigQeaJCE9qwUigVM2LLcgSseldrgo9qYf
KUyIRqbTsCAkwSNtSP4VopKUdKhxkjCN7vROgIW/2/augl6T8XgJcrVVKfGXbXVhdCmGwSxkZmMx
Zb73nxcjMJ13TsLyBtUFcP6VKBdhljTfxyaCqSZALfkhFwYKJNUtXKLE+vENvpkorwMEUBOIr/OG
nPAkESii3SJvvHE4R1vQNVfH0W9ogEX8wDExHcO4k9W8spAmstNJge0vrx+6fbfEnqAEaowKrX34
8ilZVa6RC+k4nDIz7QDQwYuUbqCscdTlM7EO02Bdu0JZHcdCNeNwlgxvTO8BO+dUH0pWIiUghKvC
l8e5Pc29cibCqQXcIsVJ3k4tdLzcZfJXQpJmLQnlUArvYPJytCejwHCcSS72MOkcaEGEDN8IJ+vn
uU8dBUeXYqF0sJNt3athQPOJGbRTg3hCGRbltE5pNUR0f5B9CtpY1Czgj/cNis8x7Orn1PI39eGQ
JchXl6zLER3F/Zq24Ph9bPglGoraCbc0LZ2dS2SgOYciiCA/uMquDOI1+KPx2//vLlGRTDbYf/IH
5SMncx99fGiW0lcEPkAo0G+QTEwEwu9r2AKD0+EU+7LY9481VxBtFAXlEoVhFkt7Qu3YebSDWlSD
X6c5ihZdOYkmPzfEsZujFU9E2qT9mEUpGjYZnJM+5NszD5hq7tZeKi4yU42kfnDDlqwHl0w/f7wG
zK+mKAD62O3iR2p7Wcv/AIvUDI+XfgTKAt9bcRW/dB+fynw8ZvPHohzd3CgCx9Fd0iQTGNNbyXHL
ssRqoJX9gFvYxari+Y3uwGHf2nHpWSY2HxmdRs0h7GjvNggA5JVRkQtEjIrTJQaR1AZHgs0bRs73
StOZUDBKCmvB92FwWwsqwidQ+akQhY6k59xXqqPjG/LuSObK5wC5Kc0TqPmtRgPeCTsDjsDehmlz
fribOtH3B01cr9iK3fNh6b1N6Y7Auq4Pozj+eiqdBLLDV5e/O4wwf3BZSTE/Rjn0pmeSmoe5u/2f
MG9MyjU5M0p7BgGnh9fNH+HovrdFdvH5PjUcu6gAY3wQqJTRAf8T1ATQJ4Mv7DX2fMnp6mVn0JEH
biZzGcVuqlmd/ONvs9Z0orSZdbJWVjJVcjvzwv9MXLTnXgj/c9gav4uZpjHP3VH0pyl9LR/IQnIp
NPZ4h7DtmNiYw3+y8tL2sW+dAz+JA7WeANPpoiF+FGi+0GSH/GoNkMD6AvTLGrBcA7fs4o0hcWAb
qCkIWVnDj5GjCjt8CQh+fWPpJ75TP/TiAJM32dz0aEBUCIG2JxKDEz/KyiPJ2zlIJIms4k5mkUMa
PanV6Upy/+ss2ZQDQL7cED9Ru4KzMH/u/XPomOB2/WfG2R1ZBIUudhOYBQ3jiYTude1R1M0f7OG1
PGprsyXFgoZyxki/6nsgX45F8NoCwEz9SkkY1CHiuuxS9YQc/7N02OHT6C4e7S4sSXd2BMnKed8P
kfqZbtTt9GIN2Fv6w5VBPbV28zlgdsxMCK5AAXlVPy7rCZ2yfOUkL8evba5G3mlhDsY1emz5IQFd
9B/nYoevBj5N/aVVuEOjkWEghytiS5od7aWutBAOyqnjYKk0KebducMTCC69pSCk8mPPhsLPqqNY
6JTzrjq2kOSTyOCAZxM+eMb09dLjwo5xbcGDhgB7QXK0Qh5RubfIQ7+D0im8y1SwfVEePBVMVe0D
lWPFreBWjzRBT8j3BOwYSiPLzdmIt6TwwcmZzkzQaGwFJnEp+sPqzTZswJDX/SSH/kqL//qPICCp
bHSy6fafpsaq+cJem2SeG02E7XgGzpR2LBkxfr7qstQrjmJs1TP87f3vMQVbpFXaLSV+NhlAVv5x
OmT2yE1szfQQ2LPQ0vs2D06hyQXr4nC+d1rGqiB6eC0WWYV+8yBkcTsHu4GhpOnCUSPRtImLaugE
8TD0JQFpkKA/a6MG3cNQc5QXwRRnNmwoMCyJtX9Bo0EWcJFFHQQvCD4bb4nlV9qNB0RcCzXg5ElW
fI6fZzkJec/y+nxl9ckkTJlDdjzTLD2kGTgvbCAv+xizdi6H0febfFZCjzWhqJJH2XmG/gI+p6lJ
v8KSuiT/tVu/dbfWYRSWYKCU93W1x827BDOREfnMEepKYLX5ujjphIJj085NYLVAgEZPmr+ZrunZ
ZmL1r+cqpKeVcvxfaVN7/dP9mS2OiqB7toNWi72nizTAiLj+CT9z+aFizVWLN7OwKxSlPHeddT5m
guOymqTWgPijY/VkE66NkclKIwDviRXDV+RZ/X7usqpHKl3vxlU9/D7k/MOjl0hbC8q+4JK7jByW
Y2eyun+zkSZroifw1B8PnLDIsPbK1oqr035pP9MLZTElzXSblCgUaLu3WQADjm05qt9VOuGdF7AB
HFWbyfuby/eaJVS1VMYDgTlKWpqhW6HJ+sVBKBASYnQuATGADYgrIIYnU4qYWvjfqu3SmJYYJibD
yV5gUxQ22iUO4DYQM4cSw9w14Nw0Y00Z4giVduxntawb8Qwq8x0ChsRc46+xy1Wfyy/s+sh6UBbE
NmY77gsMx16o6UdaBAujoUr80OPfQ+obhLYKanLd4DY9pRcihhVj1Rr13w+JVYAVywrq7iGdkFjO
r4h8oxCWDlgDDX06v8RvQy8Qqsw2sMSZrW8WsGRRUxhssITjjV0QgVf5G1O8BRVSd0CnDqBq8ZQ9
V9TboOFVpVMLkfkoa6PT3CONGw0yfkjVdoFkmFu2nN317FKsBeHY5OT+evEjpvfwf2iixCWoRYcB
tFPmQcTSWaykbaUrw7Xjy4YE0Jdyu25Zli09pXePP+r3ev4LI+ZN0UOQHiQX6o2BIaZKSnNTLaGW
p7a+/idyeSB7v70QJ8a8xee+eYRA93QGLyrN7sNnIKa6JDfSs5jMEpCpKAwLMGHE0eM0MoiL0l2o
zt2t8skzBTbUPmUIyHQDWPBSVxF0CXnhdEUOrwSPTL3SSUhwi+47yPQqUgkILnVRVY4IraEFzOzN
4GUqCYtKnV2I4BpnYJgdO4X4ihbT4k3WKP1u0UH+F5u/I/vvb4uDM3QW4eupyruyJzpdoTnnDfH2
IDOdRW2PgD8rQBzMHaIyR7ozY2kC41lPfBcRkftbd50pcfhFRZ6MaCfiOfczZuBl3hw7cPbcPby4
pUUSatQ04zVxAFBoiwHUn2Mhtdp8GbvN9+NHXGH700wxPX17YkQjuhY5tQGUBNM3gmu/VbrO7ToN
Nhja+jUI9Rxli5LVLZb2850JKVPzVnKH2iEmuUSBv1gOH5qQbJ6ycfq+fdf4PoZ04c62nzYGDxJ+
iOqX8MDBj0D6sRxzLXZLTpAm+sCmhUq0720ckbAdCv08WNclCVbLGXIH6V5sA3qMrM4XFX2F8MFj
P9ecRkcvEcHqzGOfortkHmIEx7VqB6FwnPESfy/uPk9esqz04lHvo9S57xf7lCmPFQiJYIvwEb5A
zGq5j46fRcfXjcYY0Dis0n94HLwuEQU+cUkL/oh2nIo4vqRJt035pNYb5Ev6+fXnWFyxwghTEk7n
d34Y5bGhwseyfQ9j75b7ogjVpDuSdIfIlcpASAOWFi5X31lp1otT0UccmRCs2DNq7oO6Rdv27Aav
gh7a+OuAkQzYkomFoei1UtRPZznsSEKWQuOMs/SfezPAk91K8OuWgYOsvBS3z949sU3H82pzi4wM
nwX+Z0lB7OAHoXuv92lwIrExsr1snuLfUj3QtTnWEnRX4Bs7R8rWzILJMwRwvZToup/FDL8+UTWx
Ge2PgSDVi7rvy6f0LHwJaL+58wcggFWXaRBtYcFQvDv6RKzdkKfUXNnqYZCfIkqoO/N/r/dqem6m
oBD03tslprnR/ARRZhtmsPsKC25L4SftqUoZriP51Xv1D+J5t5YoYkiO8cX+0gP+OQRaIW/bNyzT
HnnAVlpXWi1exif8qFE+oh9M1uOaGsUyfK622mbZiVf185Ms0MNbuY+uTJZqfuaWKovl1tLaBKjj
/cDJKTZURdaTgSCesEUwrGGA2Q1Zh6QwhYiZWXmiQmpkLZgOjbbhb6rqWRVbqRA7bk5zckamAVQ3
ckLngh/P8v4kyT+QgmXTk+t3NvDT3V+208lUB8NYAoIj6iyV5Y2FHyYypYCXoGe/goehA8FOecrQ
DTKq9naZTej0fu8eKFlmDeSfzoxHBhhIDMXbLiVLW22MjFlJZSh8tIU1jCZjI4GAT+bDRoGlwdxE
0L6G9cK1P9OAO1E171kkKcO/4LyQxlfxjQv2PCeW0NC8T4m8KAbbxg8xPejOL/XYF4QIcgrtFeYd
TPzzIJUgx6nLtyq2EPfmlv+5n6APyqLWFmrpyfV2f6F8RaaIx8n0LaG3A3FKr2XJwYELfcU77aoJ
g5C8aAejemUjlpZlugk4LEZnvApT4IM0BWiWxqLOYSDLXpmxVejwd3GyzQNYCm2/0WWT83tF4qNL
5/c7eNVbU3yNhSyTJmWWLgjhE0OGWmszBvkHlR73gQBoA6Wwpu/b2DJ9UqOmOEh1C1KIZQ15CkIQ
rPWX2Zu9k0EwCE/0QbL7iWcBnAfdhuSeChJf28oBTKjyZXMXbu2fbplX+nZbSYAWORpulnHAWUnA
yDay1AJfjum2eqchqvL5yfdA+Ky8TBapy+NJHcw4gqirMRdsl6UiM8MyAH5e5kwu/J3sWnSpSxpM
If5YrH80hKq/UmclTERhFAtU1vEwHzvZACvvHq9i5Jb7MDCm7qsJ7zR50QT8TXqwCPyaye1OXz1Z
LINaRscXGBoeXzYrcs6jC9NfSGZ4tAXNcXrWJIpS24Uy20OcngCHquE41n1RghqLDsOQkqkInQ8/
nWnBopUvMinOhGa35mxfzms1OrqE4IRY+BN31rohz8afAX+abjJoCUP1aEJK+cky4+4KubbtJElD
XoHSvNsCD/nNLIIqQabVyDLiAJCHkeVY5DrS860z/waVMjlCWcgHPJ11x0q9CB3VvFoXjdpNG4uu
RRGzhzs6Z3/sJTzGTvTilmJOitXr7FMmPm3c2wq9Grc0oOfR4Z2jTOUzuMIxPUt6VHZOCr3kC72z
GWDqGopms5yGF1f8Ljr4H2ywNHDAFctmbGU8g/FOWX32kE+4VBVnXC5y5gndcFVsBnryvbmr0cps
vs4lugOWiJXI0vpb874zfvi1+IOeBOLOE70n/cBPyqSF36lSZxdf+65UzSp56r0c/taOIoFHLciD
i+w3mtIwHMElnm8w7vghsbXEkxtxZHxxC9BYRYD2kBKQxazk7n5njP3mHo69CRO6zy/EmXXPp5BL
9+7pJzQ+hDogn6KYlKovmqpDnFHWM8lai1QgL9bl/gaVpoEhF3cUqA52AgvmB/LfovwLnORdimhp
zJjhcwLZFA3RCVrWhgVeX8wsVLpXMRt7ti7t+Yl4kkQv0lJcWcznHjiLLNG+sxH+oRqO1uMyLDNC
RFdI3QlyZ0PuocPvauD+RZ3wWabcX5wgdrzkDuAubmdT7cE1uBkWGXgg5Tc/FarlfzTlaVQVhSZo
Xoo3p75dguAbgidHw5tDgDF9DWCYEJapd2Fe/k0cdhttSdqv520mZNkdPOLG4/oNrogiOpnENsGg
pQRrx1jj+y9Gn5b+Z0BOdsYOZk/YWbIaDXRzU22tsiL8+Z2EJrfgwFPFtzC9qOB4B4MaxhRxkaVy
HUZ4ylJscudW3URmtPWuecYOyoTQYoMmvC9C7JaPF3WB993I90IlRgCubfhZczJAqSrrCxOo9CHc
Q8OF1uyRIecbYgoE6bMrKj9E9cjDNuLrl3UGJDfpgY4u6giiw5250+w+efClGQiPSY6cgswhA6RE
jUwZgIxkja15yYSGnLAVh4DhkED/J8MakqpivwKIhQmtCfftnYeX+DSIMbzgj4rDeJ4fZaMZIqdC
OWjom5vwYNOkpTglWXNcK5jTOdx7oXPhVWRKt+dpQDscHOFRvAOdD7IFnrCv3sOr92NVceyDAAzM
108a579HDOnm6NVLhFMYaHSbdhF9+3zMiSoObay8kvMor96mOuXIbWXgeMWGvPLHwWxwFjpGci/I
1+B++E+jJWaffJtbbyBSqXoNmiFnb3J71+o1DCcyk3Ywxhq+T/dThq7CjbvL4/VxPukoeUNpPCkF
tCzXlRTqpnAi83GpWjcEtMLZhTh9+avdeJKZ0NCNzCmV1BxaaovzBtyhQzyxb6YpTyQAbGni8jOP
2lyO4iBG86jovyxpvxWS4TG0uKT75rkOw2YuOe7QctyT0L///3NihLUlL2TrhANSbkrNuCLF1Dsp
sEth7Kb0J7KXvjjFLCEqRYeGM+IovQfyz/ShULLNiD1SSGujIVrrrrUCBwTecNKchhPmfN6kX19h
CsSJ0ruyQiAsp/uPz35niJDYVw2yglQGGbklc4Vtis1e4r6hSBK4LpOuCPC3GqPUvbRvDIpcKISV
OvkR9Z8gSTl06fZBjq3BHtuzbXADhuSo54UvxPzLhtpsS7oaB4p48CPxKKFP4+HkYvNb3o0w+vXE
C4EmPW3aCffrWGURZNN2Oh+iFjtnut6RL+JDkiUDj2uM3Q0Bifw5nJOqJ6KwvUVOqO5r/JR0pmHv
I47EzqGTAeDJkZNzkAF18kYQ796HZ6njtj+AdKtm6TnPi6wIcaqGF4w/obCN8/RrvJaiJv7hWBHW
UO9SsP5VLgYeSq/wyWJhTJHSovkrTZe/9z51x6DVyN6Yr16yqIcq89ZNI+lg02f94PPaKuUkaaDP
7N4vc5PaBfQxx7VsrNmsBdBcu1dP57JNORUdlmrYSs6jpIMS/wsvooaCCOatoZ3TWBc3IQ+i1B8a
BtoB++FkU8vXBpw11Fwkb/+/W0EwmRmY66yPleQQgXpUfOxYe3hT7OCfohU9R5Hz0dj7K/4ShO/e
79eh9aDLrUl7VMB3hhgvTzDh12O5IyJDp44jS0yTHwFgri6DqXmWqSoRHwfi/QD5++yANKMiLA4O
8Urz1+dElcY201GB9aQGn4RBQB7SEv2Gxd1uHZcMpM4KjKQNgH3TYPkA2qcjYJjjsvRPGmibEh9b
QrnCJv9qlZr8zAz+M1tXBMZIJXihn88Kgmq6JB6xMaKD7gh9EE+8uyBAjQNgA6kSBVsS5aYYMQ4n
hk9VmH8Inn5junrqqZF7QVi/fT+A0V3b9WkHfcfdkoIB9LPVc3UgRT0SpnH+r31BHS8CT1IIVRAN
mS3KiLgNoBtkDnSRbPu322lzwRjZeJjuNn8tydG7whuPMotJwVeAcR6mCYw9hetEpVTHbVqrxiD3
uqSySYpIcWhLORtMdap9TdsBAjb6uKK1W+sJkpgn7XeAEduYK4Al2rsRbXFLDqNcqM+OOlnfxr7Z
RrYXjEaCa9hpC07L4nr6LJQtD6KLNKeVvcPC7WD4S9SbBqHw0P61xuzYiWYs8iIM13XvwTHSvOi7
2FZNHA4EsxV5fPiVQy5PIIy5RR7PTtgCYyY6oi8qosgu5Dn56fVY93FPDo4Vl7i19CN3KUyhx/co
36oBZXg4sGkx5DVPK5T4qEXJ8/RDteFvKGArJ82oZsJw+pVtJipgTmE3QrBJod7UYZoSM60zuFPv
RQzk2ldPZjCe7/uzkC5fceZ8pSaRsHf/YZM+VpiQy1DPFe86VnCK0QaQFFZ5re5QWC5yIge9JEcw
/KcZ8eq0n6Juv8NwjO8sIwXKY23lAytPlsmnU3ILdypwlyHL1efdOwWPS5vKOu7n0OzBi6oGv6WV
Y9QotiEPnMLSm/NCOBQIETLOextIZ92jlQmv3SMrI+VZLC4BJYiyXGh7f4UB/A+m2hZDlaLKszId
7O4nwA3s9W++QTcxrDB3IHFI2Gd3EFNRYleeDB6m/ctLGeQL19tsBRvQAAUumENxsOTHibBpQ9lo
oj8MB/hcExjZLISFSGFY6MNR17MtGrb2CCqVELLCLsZsOuQ4edp2ye8Dyp0hNhq0Hp28y8gDNV2T
u7KPAk6W6RoWnouXluGuFH0TvH0DjGWl0uP3h3qrLjKjX+eIPWtGT3M/w/gea8BPmiSsisZsODkt
BKyJsvk8BIH4xwEAdqNx/lR7ELQcKT5PZ5VxxvDszY865KbVL0fqLYe5EivE/D4XX8QI3vXIArIQ
/+lntDi6ehuCiUPMfpjxpzUEA23pT4mFR2M8KbbbiPyOMn3ge0wjBTO2vI2m2xjc2g5HieiZtf2Y
BxbYuiUXMw9AkgPova9ODVap9vwXouHTc3rJz9qPQRA0GKRzC1qC7cM3Joii9JXOHRCD4m57QhiI
n3EgKzGQgRCH5A6Ze501SacYOQEXZEolcIW2d9JWMhE179pDkMD8AllNh8WLKMmm+snYUiKq4DnC
j/UcQCj92/5oc7vwovlf10sa07f3wQC/lyhfMnvWMpMfvEh61vlYGUp1n4jtpw3fDlozncIRvS+K
BRCOeP9KDaUAp4gpzNQZ/Cs7c/P2pi6Dqw7fgDWlZvJhC+9N0uDx5GpTEQEB+2zXWKPOeNFHM4K5
KVXdMOuY+Oj//tKVOhD4nM42Z+ZeQEK+02NiCIH7XmffxVgIL4fIWH/SUodsH0qa6Tw+5hgkS3bc
Bvt0+lmzc3/CVCHepu5NBq8vtUzYMPzBCC/Zra7mnBQ928Rzca6sGGpUUPEmNAj++Aj+/xBxnckW
19cJzBl2KIBuHBcNWp9k9G8OScY+aSoq2/UdGumx2aNhrxOOwgntMVA2EBvgPBuZiq073rToojEx
3shuIzWPWTsPKilVjLzBX08t5K729Rg7ks1/WqIjrtXSeTCl5fkA7drqFkHH7OteZm5JtXzJD597
yH5bq27RDwso7B+XOWOGaacSBFOgvyH/lz5qZUh3i9P+eSFJx47k/Z/GmFONEglAIE8cupqHjDqS
pPS6iP8nSkbXLKL55vqNN7a+Zfn6Q02LD0/bm6O0c4LUd36+fLN4Q6SY1c+EVUN2T4OjjreXH+a8
VlTnQVlI1q/E26+N/iwOIBnHdVjLSmW9/QoudF03eMhfe+DMFMLco9UCmS9nnCMYKol+r1lHFeca
1ed3ndfIfr1Cm9Rn6F4O9DZmCQPAUnxbnDbGLDo/+xFNVSQ2gJHXKkWTxjaJu/sVdiONICZXvnUP
qgN2zmVdKVlrFyZB0ZEBfNpOGIb8Ju8pFAQwaV2gnMRjGpiOJx56zgOT4T5dhCWgk2csuFydBIF1
PuYkauZhq5uSboUDrcQAh+2M6oUbTx2m/badCmU9NWl2A5xjkNWhDBUHaoVIdVKLLzCX+Gk5pUpQ
BwSrWGurXgmtuIEiXX8ACVZReVQhbmb7v9uigFCHVNokG2W7iazTUrTb1thdGj/D6S76Ma0I628j
exvERqSdoFaB6kZsvZSlf7xHUJt4RPxU817WM3f2zutsxU2/qu9XN5C+YuS9NyYQM6fWlwiU2huz
aqlYKFNirIwfQgSYUSG/zyy1G2tsyFbFaoFu6DNv9/z491pc2JSz5+7CS+3SLNYMyHMs9Y8KUrw/
mNDUk+tCubmJ3irTnHlGgn84ojXBH7HITGkgPSns/Ez4CUkPa/8OKejEh1bb8p+QrRSkhugX1aMm
ELNcofEOlDF/Y/4xGLGEC2jFqZUXp4lEglM6rCT8uYItXWJSj9lsG5+zPGHPlAkoVx+2F1UhFovN
KykoIXVeYx9XnsyNVT9yCs2B1XY/b/Cab06GQIFYPDwNhppVXOK1Dl0fj7eCLk2NxNZbhqZNr2Sh
nt49wnpVhd2+nqJOZ5YtMgYa3aQ4rySusdBXFoiwx7/YF/maSBg7c61kOTV93hRz/6d14eEg3X14
cKWjsSxSnSCfHzl2/C7kONuFIFpDiwvqTSic8Z8BbFGFt0dAPepKA+i+FJ9klfJMlwzONxOtCEpc
6DYexP7XqBfJKQTNDvpSSOZaQ2fyCIqjt2wVP20qxcJ7svoc5fc8VRj3BXfHE3krN10GZ/SafAF/
Domrs9NPM63I/gpKhYxaw1RGcZdC3mZE/dx5KKAWwYPIb7e/3Q24tJ9HqY3TUmptwFhgrDG5+e8D
beUOpnEcftRST3Cem85tO/e/pp66t4IfMedd2/NQ4P3zNlmdIXK3DD2l2A0eA6y7lSkTkJloTAIM
EeqWC1e08t3/+13tiWxGLygM17mpOK7HyMG7FMUOycUFIit5NDLtA/vuRWuTZnE/LthhXlRG03dc
2OycEZoKeqi4Z24AKAiKtlVGyQDhn8r/u8RS1kb++w5JKm0HMLwrIDVSO5qW+iVZES77vD8BXgGD
M6rvtf/uy0SubzjZ6naBB6+AZOAu1LXJGD2N8uoyDWKX/mxFnCCPh449wFoU7o8HJsl8DCtf9OFN
+OjsOgM5GGvORD0teqpjlDGVKk2RQOjMjhlnyHRs6TZNIdFSFH/QhaaUp9ef+ne05NyTZJj+7sVO
ts3oFyaxbBsEfzvsEfWQgUPnIesCB7Cm55XxxcXqs9XmXbTGyX0twJXOrxQwaPC09U6xXLQ5yOB6
NBLQMbsoysIsP8cLILDdkoY5NoLXiPnyqdBU02OikQccpAOgA5+lM4k8swS4LwG5OsdxR1Kj3MD3
6UVi+D9KAxxurXTXfxCA8oMvRLyLVj6QljqxMHn7mVW9jImuPYcw3oggUTF+nXlAVQhQfjpl9fJ3
5uGWy0zgN0dD8fZR2G6dELs1dIP6U1I83c9OItaw83eGgrth5mcbumoQZKdFc23DvbaNiwUDNzu+
X+mEdPtyIgq+Y6CUkN0DrlIEotrtYjqZfoKTbg7bkVmt2/lzt4lXUCdjL7ZCKn3+q+DJPK/6bPxv
KDsGGd+FC/HsSRUaOpFVfAcs6AHybUghlhyZNZ0XDDABYlFwaw+gXgagOlF1XEM2JxDDR4aEn72i
p9ZU7uFcqwTNpHYdRZ/uLkjmhyZzOu7ICzNsEx+kDRjpUPOnlPCRxdmLPyigLdsFk7lzKBBhohMs
ftmvDCAD5LuE5m4+lAIeZJcExgGEMW2QPeJFkdI2ykUvCNsWlPKBx0Owdx5hkX2n0Ioji7y+vHl1
MM6RGVmxJx8NROpp3vA/zYK7K68QpckgVKQ9gZsAgFpndFHftq60Z3+irgnZMQhARuby5n3J0DXx
UaOB03WQebGVTlEkl50DJibWtGjofuzRd1MwONhuvfUJWE1+I61HIF+mTm08aj8cAO6YzbqmfhVp
GcIQCL4OvvJeyZopdJIk7Qc3ry+u9Qs3nQDAf7cjCR+XZqqyKbpJRwLIvYMr/+1GjAv9+xA3yekZ
edVlJIuCWk/6GOdRATbCxu1JJconD/XDRxPphAvH99cdSTmyxdMhz4G5EqZg5rPEhWFeo3EG8O89
XK6swt4Sgszj09IhPHqZjr9mOA9JG+2tfGYc7Wh/Ds0CBqVNMmTlaguKkuwbSG3WTDuyeCTjmAkC
TvhQitg9JGN11KPpaxNiXpBl1onhbetGWP8GNxCzU+C4dNK4cLp14J0CicwHf+1Sen8hkCFQ6b/R
JZQVKh5KCK4ZlIh2ZuYgxWs5bplwKvyvRwnM8/x2ce5rDXhiRTkfptjV/WAP3PR3M/DO5w7eA7AO
EeAbW3PxPB4/YPmx5fTg54e+8fi4ITW0i6t5jBgKahm48KVBxu//TV2ZDpkCcSgvXpCOKcK94DEi
7YXihqFsR82RETH5aO85ifTlKqC7SN3ogtSt9WZT1pcHg7h1/MPK+0wH1inpWPps2RfLx/xFkBU4
XbUqQ+UG6zIIS2y91Wu+21clZvbUxkedtZtNdoNDT3927L37zLNZf7bWuXEU/Q2aBnO0D0W1YtVw
qIlRnsc5U8q3ZcL73XP364HXUpUr/+hJz6o8y9O0kwldYqe090uDa5fPXL+uT5VEzxI8hMsrvqlJ
sQ+LP91oHmwswBfcSq0YbdjFQO8mH2+32Wa/u0u7/2rYxq7xbZ9gOknMclMh9qoM+RediCebLyPh
4Kw4xBPvEuubGP+Akz1g0U/AUVsbg/ZaiyVRXqRithkGRUmdG/ahIF0wX3JQXlobptNQEZuafdWr
9+kSNSS7x6zSMK4P5yi4BTjKXfJsQ1qOYvrlJ1quT3Ik/W1+8ByeYmkp5vh/J2ZMF3Yq0oP/AbLc
/HQyykwwr1hgryKyikYGZXF8/0twnoUx7VGmD8EKl28UMfbf2aXiaAys1oWKkIrOGn09rUholl5R
JYvDHq5tlEKfEvKvjHRY0O3BpFYrdZsdkplmhaNjIrYe8QbTHnx/CAAPZ3tvhb7roZfeh5HcNI/+
OuH78dzahA9PS3nXsJTB1xTeY0Wh/0RDdw66zTDtJz0gSvgzkEwdPYechNaXqTW/iItLX/3Sa0cZ
bRBuiXPGFXmKzDbljNYkvAm0Fddp2ZMX8YNeVuhWAirBvin7UYElgOkD487mTdNkfS2cRhPrabb7
aPE3DYPmVdzLJ2YyJN/jmRRgx1g0h1Md1+OpBUPdMX4hmWApwXI4j+uSHZVcioM8S7Aw9ArVNsXz
cvIX+cD+ty8jZ15HxNatc4REIgMbuQ3hba7SjW51tN6xSikVCeCj9GfwjscAhDCWtxtJwH1NX5Kr
Gi8JXPJNvQGJ3jUNh+XMl8t6/DqJF2jNDyADg5kyCLLVgvW8KoghmNk1lbfqgQUrr4TJOX33kB76
8pVrMlBPe8rXqn18AK/ZfZ9Y717lMdLoNkwOn3W0LF1sTU3dvkqwD7+5WHk88guDzDLO18s6LV3G
pelCNkxwG8mV5UmswY27WCaEYvxKTEZzbxpj6qoVhcP4bm9IIJ6LBRQYNSglVQ5Le60lCjA05RN2
rAIA07Kn9w3zgLw6hXpFX2pGxf0yzfXTSFWvcD3IcGEmO4Ra58N4lCAJOITgcROlTWRn3y5GGEvv
jCYJjVS0frUJfEuLJs64d/dTthRE2EysE1mIezMGzo2S8HDFi9HFKuzLQkR9yA1GGha7xJmWO2x/
HRWHtVfiFcN2BrTGNxpfJlUR2Oam03Z6ZwmzBzy08Kb4eX5x4bbZrLKZa0/knDXGfSChhoUTYQwa
k+G5zktCQNmK5eolae4EFkMu7vPT7WSyqsbmgieBuufmqOzTpaKgB5/zpt5mFh7v/fOIjm3UDi/g
PkcqOVT/bvwzMBKDvyHA5tZXIIxavJpy4dBFDuHvoEH7Uzxd5NeA3D2/I/uMSJplLQ/D90U+x1Fy
MtckSNJd9DXXGx0hOze/tR97d8NsIGVoOpILO5rg1X22LWaDYI1qUQrAJWzLril0gv53j51Rzfl2
t1KFN+7Tp+XP7+Zs5Fst1qr822XJIpY5AExY0Kl1SkkG91zfKOkfetbQLuiO2mtkQNS/gpaoFp/Q
ysvDBdDGlYqxlAs4+bEpeHfhjxpdbXl9vKXQHuYFiPT3vK4kB8upZSpIASosss5Lc67WmXB6pmMn
fu1ooCEB0X8Ci5yoW+4zgc8ecc18Eu738fhgyA4/jK/xePYRlvq615rEiLf7/k4yfWZQK7uoQn6v
/mQXwUPCmQD4ij1wrLnRGVUF+UQjnyIR94zjYJda/eq5xYnKT3W5phtx9aRb6v4wsH8V+IkMm5QY
zm+1l+7fhrHNUcK6BXyOj8gqPewKuEwQdsudC9/X0hG0xvyshaJIzotJwSxEcJm6aPFZ0IiMdyvV
+rrF+/ZauPRrqhHLaSjqo6k3bTb6roq3Pfcwmu6HnzWHoxumenem81oxLD2+DJ/jpQmGlnDZLaYc
lQw+RHL4ygyI9ezB0WnypiP3T37I+0kG/HakQg/0bxEAaGrKd8P0Wjv5hvID2oNsoa5bb4yvWqtn
GWhQSr6jlVwkqCjheA/V7oFItMYzp6Boz4zr/2IPmBMYizle8M8Dan14StTv9/3an1Yk2HHoVHvp
Nhcjq8hZp8PBj8W4iyTxkyAlPkw6skg5jaUSd6ppveibnAwJcnBlibzRrpdOs8Z2o3skFk/ChjHG
7Yldh0ge9QNOl4KP4uv0QwREZu1LuyIRNeMCv3RAqk7V3/fyBZSzwG9eoa1muIVkkv3MzAjH9DoM
XhBtn0QCrHg+UwqLWSn+XrHck3zmjL1ZGNATb2xHu2wCpAHI0ZgrNmZhbnDQrz6h+dli/PcLMgax
NQgixpXREmO3rqSNylP1bKpfAV71ZQIWYeW3yOrcANvTyXdIazFe3mPhVUKHYtPgQup7f6ZinJRd
SVqj7Epq5dXT4eEjy4w4vc6tdZS9tHqmzZjCHnsKUl9VU6amdGcX2LvVgQQVUOnx0QI7tCNmQJyA
mJ29G9H4ZBRuDjnauQ+qQwblLiak1+0dN8UIqR9wMCYwqvirFa1NoRLvaUoaCbnkwTGjsljb2t4C
u+ot7jdNtxikI0FoVrluo5ZRGYe2h//KxD0amdHqE0FmWFPpj5nvKCfYOrLZWPyKb+CREl0oyOL6
azvafZP81ze+VwINrWtZOeA0e2Q4HBTh7y/hX6U8HJB8GfBUAwuT5h6mYrDjZJTBZblweqFJyATL
Cv6oGKu00No5jIXz658AJTeekzPtVdxJf3/MhCyXe0kcFZdN5VUeBfQn1qYIy3aSlaRV6ARSP3ZD
oZEie+xbeldLRWmbtztTfONRA8IVD6esdk92ZKS2/47KHr2/1Bl85nR7u4+naVmEPo1zXlou5EzD
Nt6CA+Ul+gdLixpGBjtQGKEisga/XMZ55guwsx3x9u6Pa58joF74E2G7rzChiXqo4hiYRALNrdIK
rD4qL1bSWgToU8dYwr1l5j6cRahbs9O/qHC6Pido+0MMCyaKqOaoLdB+CREdK/Uu5ZMQzE0cxpQg
pWFJ/5luRctwaN2w4pkljJ5tVEQxVIDuBBqwO0UZTFZAa7A3c3goK2RcW+KpgFlBPQ4M1hQg9uiW
tFNIWkQO4drD/zkzObGt/CvWdvAtXA/7waGpMnVAlMkgw7SSB0N5qjoPGtwayWJPGhPQsZSoavfn
a6rdCXyFbHaX9iKgm2j5emhEPtYhdzwoFKBgwBFAMfJ40zg8se5t/Xe3twnKuQoaIRbt+pLGBcbv
hV1IJ3jsRsMoxOUi85ACvB4upNDuCIqj4Xpzkwi7Ly8hfu28qBeSPwSR4pJW2TrUuhY0ipPYDr3b
pijlRYiR0WVKIwZ3nbSUqvVtdc/+rHEiicr2T2bGj2qFnEHs2GmLjnSIWo56EiRpz0vw2CcSCXhk
ITw7mBCeYk5TBDagF+u/cbp2k9S6HwvDZoPBbpD+Ly87XOZ2AtXdEm1XaGE6kN7sj5POYUhLrBzq
ILUCGro/TQ07E2uthWQG6FbsXQPvN2SRyLcGV8hBRTcBp7HEQ9L+MPdQR8SC3gofsa74a99XgYsx
IctG9ph9GTFmkdCf+90CZETN8tepg8++zKdgt+1ONDt+uyJz8Eb8u7EPM6L/VXRhOhqX70+OcFuN
pfoPqh6E7K6qkGOCPbBmItDBa5u3e90NJY00mUzL64wVjLamPlXRfup8C8+fWuu4DRJSTZ86uJ7C
/UOjf137F6GSyb6OrvcKgQDMXVM2RELtEyuXtfAB/T0tPxnEmo+5Hmoyv+g+zQXj0bK2rO0Um/6+
TVC2l7xCvqKLTKJ5rtRldtu44E09LSsKrWcTTW4q3FCr8gts8tWQgQ3CLC3FDCj+N8RMAougbSqc
WI7YyiBLmBA8VBpeTDwzJYFPfGxWORixGSaYcf0K3KENHgDgK1dUugXpKozkw3evJw6vppRWc3Yh
qphhiKMRs1uLsMiKdFz4W6MY+dThcShtTsNeNSof0R4zuX1N2j/WdHqFEG5y/FQQQf5pER0XTwKM
l/La9l4Ozowfzkcgcn3zr9fDfsbZH/L1CD/iyhCLbVUQLOUJ+jYAVIUk8z8IIUhNA2AWbos7bW9+
s0jFepUXfRRbJRSnZg0Ikq0bIp2W0td6EmtlGeqBdwTtIdWZM964+UC4GSM3gRMZRx7GxUg0nv/U
bNmzINAz3rwe3KByK2YsPPW03xRMY4sWXTQBniZRDdlo9ANruuowCWie4i8CVL5Wwe1u3FqYHtlh
TraMBkf6ammQQFC0pf0+V+ev0YriLUE4K5Zwu/zaZWdbGC73zorjeEPAMBpAQuIfdNVqKfHGNvma
vhwp+Wt0wzeccyJe5nyr9WubQbKN1utfqgj2bspOLdIXQ6RBCaZKUAqiMmb9EcLwVCSWcCOaNwXh
vxV6UZvQiPnFSTdeIQyj/8W4if1krl4t0sAvQeeRKJSOMVEQCNFVAzlkXA5kr6f01TkFhK+ZGCKF
x4KKQa/j4V8XIMsRTHWC5mbvVzt608fdgjAe6nB8dFn0AcCemoHq0LgvN9+nxUGuFJXpeGnzxm8l
Odnp9f/7GRnbKVjXIU/8USbzWvgIWBR31ZlDayVT9+1ai8JEl07s+9OOqGhIFCNg1kLAPYqwTJVC
6f91mHPgOPbHxy2LiWCeHdWCjCqm4zEE645yLzqRomJL6AhvCdYjtW+Jbk90dTuIojFB+l7GQU6H
SJWnFD++p1tf+8sHcgi4P0uimC2vncNHQPRe7U49FGtALntz8JU46myyOP3GqS/7QZCDuYuBoXod
n4CdiIfAygI2tJbIAyM1ATdwpgKkvbmQgbc8u/7awS47sTbq4+GLYLfWWJhj/qufwUltTSr13ICn
ILu2c2iEbOSUlXbpoGW4JF6JhUwlmPCvPfRUg/VUFgIo9i/mtGsozDbSN7quTC4AZRIA2PNXCCO5
kfeqyRu3sD+euO16PvklniFSggV0aXkTCK1nNaY02XJd1VP2XyqDH2Ve6VG6w3HqWWdzhSZhn0lG
O7HDn8ktwFvDNWTnLYFrSiYJpNX6FEWpcpZqaOyDACTVXeKJt/N5pX0Vu+UHiQRjXGq/UXniVv/O
Jg6CKzElCFY4vriCkJEHMik4tLhKkT8qeDZ9tZPG3dNpeqXPorIpbnxDnQ3Udyl2CdJwaoJ84saW
g30qEbRYAi31qOdEI7Dt43Wdk/JrXaRYa5DhJ4BBZ3VrezMjpeCvMKlS98r+tNjrwVOgz1YeI1Cm
Tr8jiKgITi/16FyYwhjUel3FtRYIlfI5RQIIlI8ZUfBcQGtsIAdU7sjDKt7G4hRvLTRgjS1H5iur
15kxb3oZk8c7KxpYgsfN/d6TPwca6PLcpN/PETpjBWw7n/4y1URQiDg7Eq32r0zFQNWBEBqSqzsl
rS2Jpw72geiqODyZ2/s1GFjllGDGeSsuXvKmKB9ND6hLCVEVD/jGRCR1wwH2rI922ZCKmnTFtLwZ
XQiRrlmwQwu53sgngvzM3s98Xh1T+LzmB8tkSJPEJtWqFuECfyiG7NCJzhOwiktFG53f3T4R3bNE
rL5H8RDoaJYG7tpVWekbHw92nHCW9xeKPeHQzQfykK3tZMTJxMM6M6UFlzL90XnF6z4MUOdHXicD
hJ9UqPum9Bp17EBHw9RyAQJgP/59bXomTwU2WT7nnpecV4/3ZcjFvVBeUVUiOKXuA2RrFd9L+RrU
FfnHg41Cgbcx2kvZKZjgSVwtsP+WfhL6tV7uFimtgeyaCBMPOnKhDoOe394MUdMC/AflpZOlbUX9
fqYymF6XNbLDJ8mGkVxGXM4mMRjbv5ldpTohMeyjrxTxfzLb0lelz03mZjYln7r/BeoKLc3lUn6K
OeOnpE6tSy/eLjLi1rhv6t5n72xGt7rv1n+ywzp6phauAgVkpW0UipIkI7I0l0AB8Re0r2oMmGzd
hH5eRd1IcYS9FNcqvv4TngReu3F1ss3l3nlRjp9kwCk4fNyAo4fyN4un/NTvhSK3K8b+lPLVysR0
tsv2jQIWSsUqZMh9STO9OFGxkU9RX10nAR2Sr84dkEBMDa6k/flrCXRF3N0AfJcIM/ZDNa3cXV57
PfxOeBtZgmGhwQByqtmVT3zP7747nd7/AQBkhL9ypqrGPefjFOkyZimSeLjjgEeZ3iQTiw8n4fCB
iGT6VRv58kxl2sg83VIRJgfDXFa4cUQOxT5bVcEw04rCER0ESvyQWblPi/o7ULh2PTgCQ18KXiBM
BIBR5KqyRJ5fOc9spU+4BMNNDz3yXtYGOtERTU/zU3Rb2dGZPdR0xOMo2MwUKOdZj/3gTXRE8Hoq
PqTYz9e8bZLbhHVLuLGG1uLVgyKMaM3I6uJOjIPXUNMhg+Z6rbYfaPjSzYyIW2AkYfCCtXRtFbDX
otFB3XtPhSinVcAmFvdDP6s67AuxYnrD4+YUYHCP/gT3i2WL4ACSaMwC2uXF3/i3fUCix7Pa4Bdj
1vOB/cxGIzGSbqfhNXTPJ4AgWP6rgn4J4VqOB/dVm2SBEtR20OeHu7dxk2KrOh52G4mlbuvoyBaX
Bg7ACllj3eu0gxykPhXOFUFlMlSZHoU7yt8kyMj8rbulGr5nqCLpg3hBHcHTau9AtYUtP9NO9P6i
0sA9UO8vUwyfpUvsCkWjcNAqsruXqU/NDN3yqcOOcyCJmFMHYpaZ1tk4lShx6K0Lzhi267sY67Cz
kn94xV21yerxSTQogmNtxdSAF7LTO2zgGeB160pdzU7udn4KoWBkSPQIYFw1iWfg7WwGeVtZV4jz
6yq6wKVfSlbvJ8gwIZJWgYKpwRP1uUP/cnJ93oAxSFVCo4ket3AOGRiSahZOTJx0ozyoI8nE0VRs
4HklRzyBT87rGRELrJoyJ4NOwwc6qwUGw1eRX/vp8FX7U+BFD+tlXpP0JuhNF1/gt7vYA8gYafUn
ifedjkVAJtK4l/bpkEtzGrz5Zvdhx6DULe/biH/6NoLufUe1yu5g+1HwDnL2tosAbjM5Seks6qBn
NHySl1k7/BZ9rau1EbAX7GUXuL1GU1cTK1J2CDrEJsZzVY/tmR9WZJHPSVmpg6RqWRViG8ubs5Hb
DKYtuBxd00XHHxdxAKiySQ7O2SFLDfHA48m8mmqKrqzINArG9vMCVZ3uSdzvt1EEY/bR19IPtHa+
xC02ck7e31is0Z3+BBmdF7aI7dssDDPy/m/fL78ayS1hUAkByQn/au2CDxho2wjtuYQJWs/LKNEZ
C0saFJDZfMpOscjBHWNA7qApsT+NSFZ213++e/JrcOYy1gX/KWfKh4aigbhcXPtFTTj0U6MsLfSM
mVFyjFACA9BZpyx9bRGy5ShtkX6Kky/9/ZIx4QqVz0u9WwZ3AuqF0Q4lnOU2keWkOaXvSbvjsDYx
xsLTFpk6bpNpFMWI9J/P+FNtu9wy1SuE0rwMeqqjrrGvq8aSo0cYOwWQk5QaDyJRlRaPmGgVgvwf
/3x0JEdsTcQZSed68ujfSpQ5PVlSfY2mIX0oOnQVI/mocUQbICbFByWft4goeGo+ZjfVAeX5XAvD
yrNmm9eVQptPq66ovIzniedLueHhfDMSRbSbUy4jgzzHcrXyjtCkPb6eZ4/e7hJPXnrT/gqbRMde
RwL3AnxOqeAjFOQiG2K6dG5oVsI2ksn2YcfkZf6Wkw+JkzsVGGLpGQPQ3PMvpOfwdffl4TPavuQP
2AqqR20GK2tq0Q0lcnZXM+udhV4/4aExAgNz6ed1Y8NRrVAMfvPzT7w/xf+UeHfMp/yYOySfe4GU
Bo8a8gBY5FbvrgMctKuf7uEU/nBk2MZReou4MST5oamNgNfHlnPLBZ0jj6ruqxycMIAfdI4sVI2m
hEhKBhTF+46jgZca+euRxV9VX+ILkkUiF/26zxbxU3FbuzMwtUia4HLcBw1kO50pjXaMYzXos8F5
TDCDvVQUFjKg3/pLAUCNgxpijAY+mMXR8Z3I+12BFZGnjnrfdYDvDGZMhhkSkOsVvPFwPK6FZA+J
fguNuDxzBdJThB9NXSXw/fRcZVBtY/+uF2S7q4iZTkDmHnrlRRFV6VqWGjogD6s0emXlv+WKxBM/
Bm6kfVjJjoiBZ0f6TB6wHvyAhou5ofoAd0ZDhYQBFB8exP0tSQ8pe0hbke6qopIRWvifkK+9nQ+f
Qh+GdTveHabJDcRsCJHzkZyftOFFNuDsCcWAyWGkcqKAKwEv/Xw5AXn9MnXoe2umGl4SirdRMD/2
3v23ax5IFUFO5YrWtSF70QOoZ4wa0rUCf142SiiRL5bhheGw0RL77VtZpBLyEkCFbEYw5fVNfdtw
dpOqhDaz06S/Mujy1H8kEIEB5UU+EJ+/2MU1gJXlS3GaCoo9W9L/LlT07plWD0OOiUE2c141rANS
k85mJH8VOYYqaOABOogxVTxaweMGAV9SCOi1nyX9Swy5QLsmzYoFm7fEiMIpI5xnbKKjemwkd/BB
9O/lm8bCJn9SLQR2cIdsV9GgRzEeLcGgEValqah3re/661WMYTcV3MrcBcrKztfX0Rls1Gtzb0Xq
9/xrzf2ugs+/fxg3iJGgYcpmWsts36w4M3/NePxOqFcYKlRUJPA4H1q8lFsWX+aMLMQZPh9UIu40
1T6OdwZRr3I40W7D/azmj7GGUmNjckDevBdQ9j1GdogQrn9i2qFMgaSyXkp0/a9XFJ15e1LcxRiw
/GJaaRBcFYkyY9VEZxwxaj9e34MC8qzDvrOgf5i+ZoNGSJb4WEJb/qBBjurkJKomxv6GoslwWRoG
/dcA1tQFNSWWrzRoPFN8vyC91EYrAZ80MHehMYbqsEBQ4wp1YXcTv6av1TyLl6DYcKjp2Fccrz8O
4+c3od+hMkIOYKCAlgCT0QbKejyadmSvc/lV324nyGhE22WEwRBdEYtP+5+zazLBeDw3V+hAne5P
GETgi9CF/qveQr+8kkisMTL7ZGMiUpOPIYv7nV4XrN3CqUgoTE/YRS1q708zhoFSC2G7tKImNE01
OhnIh5m5RzRokwTiUEQINhfri8cPVIHzqygv4tyGoh+MBlunqoRQE1f8UhxV6wLjtFisDdbH1Ztp
oUYAgUKNlx8QYm7/OTGFrGVLNZR6RDsJtc2ND8N/kMpBauHCXb4vvmcNIcjXVcBdK65jRr3I90uf
3L3hBUV9dBhX0KrHxF/rCoZ3S8mlEfAG7SWCuj8yUqmv5cSrX712yUpk5OrGwzHoGU8UCTQ8rUXj
jTvZwUE6kL/7pGG/bKvtdRyl69VF1+/kCfY8uUVFb4Vgh1oBdoYrMjI77I28zFP81R+AGHr33cpb
FQ901sqjB5UmL+8yrq37/oHhRkNKJ33p98AwGxTZ7b0917FR8BuP+jloWQi8rpCo6BRLDaBHl+wH
xJnuvZ7iDd4HjsYIw3lBvzPdSDz6GtNXuGFomfCtOUmiEGet85d387GLKB5YdFktqWk7vUASEp09
DXpV5fAyIvlQXO0qSGux3+Wv83i453KyF2gcmIB7JIJawbXpDk8P72hh4M+Ghg6bTaISOfsEaNxc
Zxuiy7n9UCyABQjgTtAlZ3f38OvA0U9eNyBKFTT8VL+ueCFpGSiwHRHiLoodDsS0AKttLLw8zfoK
GzuOpxkpDecunqlRy/XS39BGcJeRx5xeWQJdSs+ffFu33zlbzixtr8tLfr4rVO/+6HUPZ2RtoJtx
bk4iZVTaz1qGjG+ZV2pq7K0MSUeIxl5UEj7BvHwBKZFtLxqB0DdBXHMjuqfp+hcQwGPZ0uYNYTs1
2COHAmEaDSmKKCAdCvoPC33shaqRRcWwWEBz1g+A40yuWTtoZhU9SxCcjBY8PL1WC84V0Q/8AVxv
mJYHVrtnC4H0sMUeAgUWGlM1aCXeF5Dj0N3itD7byW8YpWwyLFgFsmPa7Rk+pd3anq5eyFxRfESR
HJ57bfmq7au7xfhPlxeiFMbRM/qg9b58nRrc1M7plPpEshi02ZFJb3yerfjy/kuT8f1gUjdCdKvR
TRRit8GBwF4rkEB/LNzvENqwD6m4MMe8WuBCZKXOUIdhoqFufZDTCPT4z0TerQqViFv9gXOK6iOc
2zJhnB0f3eZGYEzNB8yw/cTba6ynhw3HDWXNsw0R46y2mmnEawIhL4anIILlZCtR5c01lMYyYFOM
Zcf6Hn8D04BMNXSX5ncwdzuPSUIfxhaqJehyGDDQmXX5mTiMA5O15oTy+P30ncw1583Nm3XaBu4c
O2nvYYaWbzTWfmxTsUUTLnzxDVRTHlwCExNjHiPv3LSeSuwcLeCGdNf0IMuTuVCp43mgH68DzQhS
D/vrCd9paEGKbU7Fioca1v1yw7+iZKnS0aCWLOVR5xvSuo1qpczAlerE9dlNworQHGhokddPfFQ/
GT+gFpBriboikBtTjfRl6NmgUAu4LwMUTz/piPO9V7k56jJLrqYD4BeN46bKP0UMIt3N2kpIK/8D
cnvnEhkb4lrUGNW2sD8EXoiXxJdaMra4o7bCp/cb0H6cCFCK9U4fUcS9LqoQZlCHHbCRBCKD68ya
ZAzutgBOo51pS/Q6Q4/XaiKXi16JbSqHrwPN1iUrfnKE0ibDANMgbd1shozo7LQZxYhmVwDi4CtE
zT7cDjwLIdmDyZvik/ZOcxdPN3Qy9O7JFZp2t+oN9kh789YQ6dZ7jgWIr594Ny51YJX677b605/4
hEL2EJeJhJoZKks2QrbhJPUgAcVCknJb0SfbxdJRcEfMK/FVx1A6rAELrv0Tc3Hh+MMzMOqVtBj9
ou/HqDC7l3HS4Idf0cXVCS0VxVj7YFIU3R1k25matOclIbiu+v+8vafhQbrm8o88Fq/Q1CqGfU5a
B60ZkhbR4gnA/frxIZcC6vamUj1FbiNhcD57TkySugF7lgnMgXqTUOQ29+HSkRxpqaJDOLB5J/Ku
qX5W2u4ceRIEx1y7McCRgqENAWBFkklEjLdOK2IG8NyETfjuEkZKa8pZ5F5hmCaLPT049G94Tddo
uyrZCE6sMiCBOacWzgP+wT3pMur8zmlGygDgY36+XyyCbTLvHSSiJydudfTHPvtdi+gs8Ldlqzux
ZJjW9cOwwkdBHcgyEZtItYn4OxMSIm3uhfWAC0oYJJlKWIuUlKwU0G2kWqtqYZq3pOHa8ezGEjVI
zw3OWxBwbMnjNbgb0lXpCjSlrk907nmrCTQSvqoOpXxzaZnYno4RGtTJHQ6Vzg9nAiNMExu8vOlB
/wB5ESAk9bD3W71vLN6IKtKOkQy80on8A1G3yfo5XAbux0lLrbd5Kivek3+VoGXo+4hTbVNIkxId
0VlOP4vYXK/t9CmvS2hIVDnanpcu/UgqMKrIVP8ur54n5YSaxYGalz+NDZ7+CPwsL6m4GCRRKrcU
U7PlIJRIUbyg/zTNB1qSIU+qgwvrBsHGuXxISNGL/mV1eq7WOTHDfbsL7k35ibio0sxfonnvJcUY
RanXN8rWXvHZih+ZUh8yEB2ZJSlNPHyLwopbqz5kW42UV/8WfLgUCTF/MiwEovANPKVAIkr6pH4L
v+5l+r+m1LJnhFRKeWR4Egcf0WI2z6vH5hxdf7NfPfs26dq7XHHLlq1DcowU/Qfo4ISLk7B3xGhi
zHZKoQB4lOliMK2ZD7uDqQt1Qkip0oNOXvEhBR3dsdxnIUlPsrs5CzdP0hczTR8bl298NxXLddlm
pe+ulKwro51PDxezRoRdMJnHkN4z5g2gbDWotBt+LEUYU3wod81222kvLwSz8e9gtZq/kQCxXkni
F5QaaLVslA/qDEkOsgbgflJCi3+5bRxN35jK+O3IVLAdOSvFYG360TJyCqY+Rso+H9x8ndpHXNVS
pD/oyaGMQEEW8z98/YgGDoMEF1HhxoM2hAUUS8JVuClOqJUTpYBc9WPsyd2UI5yIurmHhWUIxEmk
GDfV0LlXHRQ1yl+/+wSGaODq+7SEuf1kzHz6PV7pDp61MqvBm+Bse7Bkvhs1Sf+r0LZWMRyZpI3M
1zqb6F4CsB+FL/j9jbZCyUZ7YCwrUtKB/dpSU48E+3aHnvhS4Uu2oLCsbopNwbZ0yyjWm++zjn4V
KlwQpDP6Y/hf1a8iZZG//wtQt6X1jp2kQXEna/aHewrfLTwOcsQiw1ywf1SEYi0iUob0ISNmqTPc
MTAgHbff1mPLMKx1ZgywrFXkJA1T9s5U5AUCpyqm6QGBQLhs7K4rUshJp6vNcV7Sca6U9zDN+sO4
DvwBw4OmDhVHT1eG4vflubbS1tQZv1L41p3B8kKPP2nMP5GbC2in9tqW1hyB5y908U3XQKPc8nTN
Mh2fnJBbylA4ZQszm/oH35OMv35EwMVFFvJIHYelBzrv51Z5UapvoqRUtA/Qcw1ESbra+4eDGuSv
bu0+QXIvhAeAVpXcDyU2+rwCNa8Xpu9Kp8o3xTUH4ux+9qyPZUUOdpv4wSF4CyPp4OhYaS9faFhC
1/u0aERFYuCTfwoYd2jPr4Uqil2SrZZCPDWQCT9xz4M/HTKQVxFAb7s0ozThg/S8WRF6poKtwC2g
yHeuRg+Qvcmw3auybCZThMZt50xixAzd2ffp+hKJY8EEZW0z1Txv3yuRC/qhvgCHPhQci88oio70
cUOhJ/zscIH6iOamRNz+KUitE7EJe1fbklgfDT8/ngDoBSjZrJaR7T6EwFVn9NaQFkn9cwogFYgb
ENpBm4gHJzoBbuK9j+GoQ6xMLLIiRmB7HNEFaySQ3LRNv/1o4EKDpuarZ+upkZzib0ROSL8sFy5h
CaiCkXBeWEGTZ0K27BTLSGsszpU7Q5Y3JFOHoIr6ZTK4ShyZEqVM6nb15oonknQE3f0KOGGwDxK8
jQm2nahBOZUavQJ2oauvrtrPZdBSvAjB4/6dwTq8t4CaUbwMJ8l4A022U0jeZPhmNweZ81IeonVT
uZuqYeZcWOnc9jtzmDIBvb3y3+LuLt/A3fv4zrYKpavwGUrFWqICs5Oj4X6XY9Tn+3hO49O0ACoD
tLIqi6HdWSs5FMblugmtqaMwXKnk896r9rptvSUbDM3PKSZ+TRLyfo9OSTRnAJTcnui+aMqs3yuE
/a/Ddpostb5eDFhdRXK5tajTlXQzxynC06tXRNXi6/GPxIORxTA1BoZ85cDNPPA7FtoBh3oHzdv5
6hiAcYh4xOQs5sdwmQv6QeTP+sfpD7ScdLuynLIkTYaVQo5m2BL4ATxdgKpteJMiw7PmukG1DpnS
zulsiP2xXdvoPyzA3wvdYfgHbsU1vrfnbo9bTAnSs5MjtkbDlNht1N3me74pPWXq5JnH//shyw3+
J4O/Vk53apTjtEJ73rYba4ZTrSQrQBviDuWeQRRj7zLc8ZmwgQGZ2ajYJd2mmZgoc2o58NJMsCqt
RxcehNdEzslCe1xFIdQolzKgXwBWxAdj5MFv9Q5OuxFxTHLFtJWxDQIMMy99vBl9iSF7/pew8lnD
JlhHtsAyKyKnuInuCjDgTrPvWJTJbXqKa9F+NwJQ3o9oTw+cTmDxfg6AEceVoU3x93j2arX3tRi5
0/Zgf0Uw3ll5PSKtGn/piYNXDL2REkE67pd7FIZTih/e9YR2Ql/3rh+dtTcloCKgIRPLSidAz1/m
PuMQrWWLTEYZaDsPJJrI2pVLHhuxf+siChQCSIWa5wSPzSUVN/2g6s4vQ2H0DwlVW/ZtBtqP6YQx
Xw5IosQoNGv4GSxywhjW/BC8zzHtakqJCRwMhhSn70+kHERYR4R5E5WZ1+RHNC/3P+VT8xfOiLsc
spCQNTKjzSJEu+xGPzMtXV+3TJYpqG/b6qee1uMXkRTWaC2dqFYUqlq2EwtgdR8+mnC80y6SBTz1
YDEU/W5+n39Z3OuzbujtpRh2/dylVTMcWM1fr9P5FAYqGlfOJVfOoRsNSqkrNxF+wn2y4ym4XeEd
1F1usdvP5BehjcrbVtxvnh1uyUppby5DCLtgmVxTg9LmAXDKtl3t28em7JEv7XI1C+oI5a35bPvV
s9C2RswCX/a67oNRU53qQ2LaXcS+NlSMVzMF17slKIuAqGctWkQkVaUgJSNTcTMEPXwJJfNQcML3
pgV5nOS9+0oc6q/Pd9RsiQSK1Q4TmN6+CtfqboL5tNH5IWAfZp6bHA/fjuhId0GRTFnibSYd6ecF
MvhjP8kcyA5UlpFEvYAN3tu4tmfDME17On/41C3lNk3ccD7QSlSuk90bqHXncdTLCqGEkl4V2vQN
pSSqGpihnxlbKyZJVL1A0kgPR1AP04khIrIjRbNBUgNVagnSMPwhYMqpcyk+xxPu6iJmgrOzV5Vo
ij7uI47kQophihbbxl8CeZ9LA9MCSdugQTltwGPIfJoX1XzvkESn1W2wW+aK512z2erw8cLKB9UC
tpi2RhhXVcbraSTatYN5cML66NOV/74x7CgSJgz499d4Hnc2eHmFdQqX95dim4G4DpKUXE9Xz8Ek
OYL17DgLOjXV8MZajbeJHVKc63znf/zKdgscL4PSh/nCvqy8GqB739njxXVkCjnEM2/eknP/xHhC
hPi6a5hDR1Tgl+bAsOhUuhEVgliSr+zbLwAD+k9OAJ+i5VTYIhbXQtcZrMDmUwL+5LbgJKD7j/05
Rm/zO+talRtvKwq4h0PjRg4+4utHsAt82qk+T5Jhts8N+StlvJYF6+vagdg8+hlG7XJnQi7D7q/0
84ruWJyvYsS73JBLa8rpQTfHzN85xm0kzqW/LqQOXcuexEz58CzBgKQJfLEDajY4bo3eUWypEzry
HJtHSDeTTnmIwZu82rpVifbfVJp7GFaFxNNZY5Cb+gog9ykfCNaHzPjJdheR4cnUNNw3tg8lpMUF
/JsDrGJaZOde4hYp5YDpmwcIR8Ze4Vhfvm+mYGF2Jo7HHSDFsKModkcIryi1G6zgM9K2Fj4JRNQF
gYRAV9Rv5FYhvVM87e7qf4n4SNh08R8fRqw+6YtYxAbAWRUh2gU0rXvesvNsJ2uDCUY8BG5BJkyi
UwO+AzUyhUxm7cBc0nlQOI/KHP9ltmlp4rBOcwTM2Kp+WIvhvmvCh5wz+cBT5qAdYyS8YIiX/AAm
71MH/ag3qAEtrcDHkn7Mnr0Hs4DSmIuRU1LFjvA0OC+dqObRy212Y7Fu/Vp/9ceDdC/iAOGm8zTG
uv8gomlcc7iLWAl/Fffd9mSw4B9mG2erfaKodO2amjum+LiSSIQcWoY6H4O/pIQzeNLjtWpP5Q6K
3YibO7X4nqVJe5fZ02DlqV0w0AtrnRbsctSE2aKZwS2vmXsDECtDF+7oLSxkFVIyfhJKZscapg6L
pGgIydJgqHvV93r56RbfsR2SbvfWOCZDuN6Yz1qmwbTeiQUJ+G/RAL/WdcA+Uog8m1P3IZRkzNMs
afahsUk3+3SA2bH3KkOqbaZjT73UQya8GCtRjeQuKdqjFvwf91KqypFC/um6CoEvCfspfv2cNUQn
X44qc31UVRNPNgQTB27i8mkd9s79BZiVFGqYiJXtcYtqQOHvhHtPOikBPkuwJ6eeuJHQJwP2SPsG
jXXP1z7VHI2yBfyKrh9VREvwFq7CFA5gmL/3isUa+fyaNNKKg11SBc2gc9fe7dn59FcX8/iJfSyA
XZaYrZpMsIjRxjh9nxax9tgJnY57DdybN3nno/Ac30ECa0QZsTjpC22VHs0rU5DMKtidJmoh2Ziv
zL++JhW0LUSpaZDWfgxveSQZJJFxSs2YCCmFTsaB5RLcYCv+9GFjfBv8MvEl58PP8AiTe9fVl+UB
/dAHZP7681fHb5i1WZzdHJY3DO2hmpkqWivhXEnzCs0h5bCZGccVdGYqRtDdL8+gZER9iZ9LpZzS
qQK2fRwu7IUILlSZs1hmIr4IMaZuBMqiR7QIu/YSloZC+/jGv4AC9mHtNG+r74ucAt7rDxyzR7cL
WHred9uwv0YtvxWrQ8CW07laiBRC4d6jQwouQiF+vl+e5/u+O/mcxe6+PdTccYNjfsoPXDATdpbP
g+aqXwgPJ9nnlERAoo9QqfEhAWBX13YGoie07HjtvoQUSLIjg1dioA08KCMq29XVUi1rxqVD6Lag
pzotI8ONYYFaHmx6LJjV7CkTtJB2HwX1wBUZ+tZOq20Vqy//7HiW6Xe8IGcxWzhjzDw9bnlmn2qn
cxQTBPJuNMttrqhETirDqOHLtb2Kvh1QdkeOZDPs9ld/3uY/oBizCiJaeQvh2JxmHImMUIWvzl+L
zB7oPEygV8OZ0i5AZH2OUUQ3kXlJpmFhYsSzFCJDPXRj+e+B2RFyRN6+UdDB6woKeat4sQCAIJ1u
LkvLR0WYEUdGPBOd+cALzw2qZs5zvptJBG1/IqdgWp9zHBwkoaWpOBo49aW/NOdolUvuiFiWLFLA
nOJkdma2NkImT1UJEJVeWt9/9SjKWCSCIb3UB8mSP0q5rMGNuReewHR5xTGnAR9W+pzz6WVIW2VL
aQKbmwkbrDj35Ek1aPOjLeCX1OyRRrFa8uwhnhIx6GJNzF+5CcQ8CdPcERw3tKOoajn0wa0nRKdX
3Aj8wK+7HgIcILXsTw9O46zCx+9OOdY4+p2e8E8m9hKNmYhqpiRHEoffIIf38dLmhr96qeHr1RNP
05us8wxWdGsApZuDPC6ru63QmSG89nt/z85P20jE+UU6q5Sn2aOxPR4MiUjStrTC6vYWm5ckoOSf
3aiaww3nOFAmIOP1qrotyiii+9V0Eu7K1piIu3BlaOLKl7T5ireEDPINVPHJ0xf05Kn0A7Eao9hw
A8UAaFGltCejBEoiU8dBa/INBuywweWVxOfvIZ4OB47TeneCyAF6GsoWE985hYk5k7F30mRRNb7f
NI3ZJH5JT/b/c2Sd0gS2qmZu4K+YlaFSApOEwiyuYorpweHP1XVJ1/2v1f+tfhy1Oqdmf+YFE/rR
O/JAFIaNn5n20p14pwLznwE/YtBahkkq6ROVuWhjhmOOH8subgu8A8URCVyofqJnGcQFdS1KIa2A
wHMG3iJPl9CY/DURkWa/ZQsq4OKqOmZcECxhHaNKWks8qIhoAZFNTeY31eigb/YIAQJPJuj4Er2S
K1Hx6iqnuRWKv9Qy+4jkODJmoXq1QntgXap/p6vRyxUWcrVgejPBY+mbao/Un77et8eByfBBl+Ao
PaF1xvFnkqFycmbV8Yp2icJDFS4IyTswuhLuo8JwiMVbqiHB0S0fDA2pSFsmCZisDb9oRPGek0rN
FaFlhhfzPKWVg/OxqEGDKHi9b9obvSCgpxJMOrj+MaYQxnnig9LVMc/L/YC5vQ3NkqWa/HB7PFy6
Cb6izZuC1OVTUaYQ/7y9sqhN2B7ixq0ubNinuhO5rKJMmw+7TlbvC+tFq4wc2awnGn1gaomR6esW
RnQVYUWgphF6rW7q7Rn4GAA9E+cAOIydXtEgEhPvT3n9Z0R+G14CY4AztMqltYu0AUuWGHKcxdN8
MLtSdA70/DPQwYaalUGttPUwvwgk3pl77nvK2LAuwaGJ/JOV4khpT3b15aNtsZZF/sogHioPWiK9
mTniGY4adVOs1TEnn6JpTdf02z/F/qXCYO0KubaetZKR1G8KMZ6TxYFXHxl+0O8HVrjeQMG/2J7/
UuvXg4CBCGkV3GPEbMjxydClCA+vr8025y/DV4QzQVeTacXuqE4arxFUdhfKvpWSYnP2/YlVEjiC
G/d4hXK2QQX//L4U1H43b7vN3ot0NFXvYeKhWUpIiC1KpbXxzL9zdK0nC3x1CO76QHFXOR1npKlr
lBf1uq0ZuCEJH0YFAzgVnY5tiqLQpbmz1LtLNmhRpAj8lV9EGgGvRC4ZyewXQBkCMiUQa+pXYnv9
WsrJWilXFUnmsMjLkbUsc3FHM8LZV+9F+uR6j1Ytm7pyTkjtieP+dPkxNBnpxQFL6+Hf/iBTBEyb
gsP7sdC/6lV1kaxOYMsf/GS/gzJL3rlnOQ21/dz3Oi5tK/3daZ5gFpsZhZRypxfRxQI/oSgR90ve
jKdHrdCU7dPkcj4YAlAVn7b1AUWWwJoZNujFZzXsr1XA+8ZbPM7OGQjY8SigOiLdyaG6w0tZ95lL
i6ctfYQuNaKBtsWXvFc8X0aoCRjq/bz8eIk1Os0+dSPtCXmZX0IjQ8nNr08DqmMxY5QXgE9Fwr9q
NRTXpqroK4rMG2Fjpz5QEjfFeSVEpdz7UxCa04VFjfylL3R22y26mfhPTlymK9ETESZajzBLutFz
B4wOaSUJyt5Q/NAHEXlCp4uhYZBcN7lM9GU4mPF/E49Uo8shXRMt9FJrUWNsB97ncpND8UwDvnbZ
8OnERn5hZBDHHjq0J8i1aPjbGSHWvUYSNj2VHbACO/uuJM6ucDX9e1h2D8UnodgknBJpMSRXuJQ3
PbYOvD4E2lZFOe8y15hAeY20r/soF5/MPrxqZquimwC5QKwGWwQCFE9+mFbJcRfZPxLrN9nlG9dA
jBlzn99tv19N0PqX4XgkY4enLo2woeW5YSSTXbRed4rublGDOvMNa/dlnmb4ho5Xf1YWCuszabNd
1tO54hqK9J4XX3tAvoVPhIF4ekKtmT8yZjoIE13HrPVVuWdl1jnxg0pjtmXZddHxncIssekoUjSr
acfoLZdLumMcnxH5jYRUlE+cLH6Y1nDbr3TuDBU3pr6mbGfkwQP2tyxIunIBtyRJypVpW2LC0x7F
2XXNg7ZU9MFuzu5QzgKe6Nh8Owu2qZfTBkJdTXTkM9TSukOR8U+nFo0y3wSnlrWwngRXSn0C8/iO
/RdPj8/mcA/kldveUVGuMYe848bnSPQtXj2BqPMqoPRjG4MndswL39YY4myLj0ch4SMigvl9w9Qi
s84DGmuBHaOQygwdIri2bXhE86auh5ORg2C9fG2cxTWWoZCHKq2bwbAAW0nkHik28j7Uo/JjmtsZ
w23z19WOo6VsoTG6e167sonRX4PC+302PqQiCFT1JkOtAcv/IR2n9HfN+8Dn3andsFBJ2vxibD86
SVK+tfBS/OIC5czlq4LNqBsYzhQAyJKHXO0L2QxMZaeJjoJiQxzC/sycFRKcbhZiK13nMCAzkuzr
qgE+YMjO7rPRgvtdcvskCBdl6DKHSfzIbckrUBn4sLktruWuni5MMokEitwtiMoJ7ccE3bas35aU
VdjFJ2PnbQ/kCx6dDS3hLXnEmKiX+kqLwfmdvkoppeXyuIpyA+ELUjGVOstdKLBVsMUg8ros/eqE
xT1LMCSeRPke2S1z43a4i0HoTlD0ICUqQaotfQXR2nAMHx9DXTMqkfOgMclJzr/PRmMNguZ+oWJr
h4oEQlbErRZs06ITsgYfUSUR5tchymdFYJyoBYz9T69nlSmAVKqHXlvHqIWZdMauSbk+LAHvfsZr
FXcmCjgYmXC0ZZSFgE3M9krH1GDrVEVx19VbQrdx1pFjx2GKhnj3Ym88aQ9BI81mQKccLl6i+t93
xgBCl4mnZcCR4Slfp5+/SjNaWP8yDLNDluVJaKbSkPlg515ypur4AHyQcGaW9Q0z6NMJFmTrk2aV
DQGkhACOCKjAS0Dukgvg475q5oDTQUDxD03HfHA1c4FlozSoewbrO7cVblks8PzzfYKtEiZLWNQs
OK4nazNxtM1B2HL6uH4TCn1cyzEaalhPmEfm78OcHW5qVUDi8vYCjq3d/A+svq2DiYQ8abufPR5G
r3rnrdNdYDw5vtd/dRLnGgjlEIKA1GwwIailI6jgspqTLnNucfjMYrDSRsDmjBUMTkbMBH7rwBJw
4FL29pu6+5kv5Bjy7mMKviJPLgJZbQX8zCsaRT+wS2t9i1h94e6cmTH2+IeZvS7JVKRw9Zzu+Mjq
cfNyVxNEA0OXOc8QxEmQAjv8hlqhUQ0rs+C4aGzyn/cjTDFKSgSCaG0bpMfiTk3hnquSBB8NqI2F
ScPgsRe8mMiavM9l75DQ9qb2/T9nuBF4xY4dE4tN8qn2mBjfwNhSocb6JW34B92VZfcjwL7KRkXn
5BAN21lVyzeIppIERZlSquhS0RqrUJpyynVXPRh3to4wSXkuIYw6ozUZZHBNkuiqSdCc1XyTTNPu
7/EkvM+tDIYdEgoqZWDqggNz7W2VbmWzm0DqpIYWgMTwn71MLwf3UVAAKh3xZ9HK3ghUHWXEMEsA
kfDD9JJQ8P0LtiKBUxKVX4S7ssqkmy+8qBGCkka5jvXHan7YuHoSAmuQfUMLuhMGgD+mw58YuLou
jr25+ivtWXxsEKnBxpzHvEntBxxmth96k5f4Ms8hgw3FipzRX9mCAJvGBiLYFw+ee1VcLB4d5VIH
cOs1gP8xkvdxqDW9QW5PYwPizB3cKawrDu3UZryxCcT+mqUZKeHGAuX7ZkFGsHuWzBqgyQibN55L
gxX/FfPsbb7qImkPCTUiPcoIcXihycf+LZrTQvRrgBZL6JQeI6jqboJOYEplz5vn0dnPZMCQ4MNQ
/b8yC/4mawofDO4xmHhOjuEey0e4Oxittt5++0HveXIRE1ZARFrmqtWfgrosfA+TLPOmIBAPtn/g
A17/5IBfuxDHVCWf2bqSl2TgDR2NUTG2L1d+Jd5IiR6INGN2Ux5WQdieOjQZiruLMe2HoMUhk18p
0JWXD0o/Tb/LAISFBvtwoGqY3NDAVkDU6ZBBcfpwAzk0HPifVPz5V1ud26OkxAvwWyxi8SNDoYAI
6lY4KJUNCQy4muDAeiilgcF4/hlNqTzv/WJio0x6fkjfKrxI5s79d4DDXNmayIlbaOEsJwmBZZsX
OJgJSGk9mwJDCUgGzvD3wG/UsGansuK/3beSsXu0Fopk5EUc39r5uR8ZPpmkcTRUsMi4hyx9nZwA
xSQfw4YrK5EBHEEaJHw6GqEqxKbsHRzd+B3ipYjr/x1hz4CKb49upL9yd/tjbig803RgxAWBzf1W
hH6gDJOLFNH0Gl0NKvVTq2LBxbVB7uyX0lt8e/a6boKIEU9ZZpmanSELJZlhF8lcD7Rz21vdAH3X
NUl8j3envf4oQcJjOnqw4OJM1Vuu+OII7paiFltGWobhoFXsyti6A8u+d5UM5Vw7OCals5j4Ks/a
RHtcCMWVTciHZMgNUqiJ4nbWniMWZu2WJlTkVyLDdtwtLAQaA6EL4/XhxRytDU0q0PXHlH2HiBKv
HmPd1Rod2BkrtOROOBuiEvdtxIeDhh7RIkYIWxgAFb2m/sKHSa+h9lk7ctFR0Hy60BR6YYCFirws
UfAuRbj24wjCSJEyOKdnhROq43iy19S7yAfAF5kt7StY1gkyVEl6YiCyaLC58s8q+BdcEkVx6JaU
wH+KDIWtxFjNs09NiLMD8rvgJkfuWhGIatrMrrKRO1GfdzPYL4TFzXXn6Zbwn25wB+WMr3hrhPGo
K0cp81dQCo+hi6OITC2cnv5gnbk/2ObRfgGznmE+G2HFFMj5EeUtXHPaPfuSm4v6/z2Plu2QQXyY
PJEA3g1iE0zio99tNgeeIFJ2788h1j8vGWlvVWJDR6HKPstjI7I04cwL+D+bKHQphZuJr5T41Pp7
EUqA6CYBygtNdIFvB9zq17Fd69wtu2dxmy3zn5gZ6u6+33i95TSsthQZlW66YPJW/wcshgn7dVR5
sVuQu7CInF3T42IssPDawz483DAQsXBw0dh5BH236fh+wLYSDrIHKPWnbpBtZRFYIA6NVYCLEtac
XYbvdwGMgE87Wea0zL3QzoOV38ESN/BV4B1lF3VOcusuiI6tfObh1M+pyx7B3L/qHK1sfV8CAcG8
/Qln3Eo7Hr2zvkkECtAp0VNzkGAWReC98fRbzhOP+Sn4TrK11N+yOrczJg9LBkHgekHj+cMJ+zNc
gkv9l7ELp3RfYH/YHWAycd2F1YWUfFKfjmLH+uDkosbIWPhXm2QLqpfnAJKg4kmEebgSgYcQxeM5
9osjMUk1gI4ME0lKnCNipZSd4L6lR0Ixo6ETvzy4IwesXvyDRudXLfF3O/VpKkoxAU6lOvoXLbbV
CuEdT+4wwt45jCApDtig4EFuCHHxkkxdBuiwn2f/NcVGsUZeTCCt79e+qrR/rfW6HcFJuQ4MHn8a
jDQ4Mn46F3Ow7Gc+IPM5TMv3RECs9W5qTe+KZc/NiF5cg5078ertDH4KmMtlrZwmJPoybG0Ms/Np
TJHPDx4lKGR9JHoI1hamGLNfhp5rIeLtnTy1DnSy49+YaXPvmyna8dM7d0KIdR5+oOdlF/wFxVgJ
ynYboZeFvSuA+uq6oEPl1vskVt43JLAMgyqu4ozDUA0cz2fvd5RAcih3YQ93nVK47TDSf0tUe8XA
s1GOcwaKGbDC9TJBFdP6fGzzNrqTvcHxzjXuiXx9mF93SCY3olA+gfFLSeT2MmJ3KSc5J8skcDSj
TgMip4a026b9TuItWOBNU13yI/MBE+u/5mtAWE51VBDl4MjGh4Jy/7D9QPgR4fVijCZkjlmKLYDn
xGuDFkYfGN/WrnKQiqkUi5H9Vekb1y8GNXefPCaNXZyibgzJLRWTzow38l94EEGk9hAawGn075sX
Cpp1y1JQZPMYN1d2y5TT5ordgh9rEvUPbhLZAzSTLEwVuhO+tiKP3hgtLDhdmKr4o0U2xfOSTLUt
U0QJc1svOppuVhACi3TlwigX0j9f7hLfEFTB5cCWi6nrYdkYfuOTQMpa/1SLj8oIPF7vTfQ6pHCn
NejFhFyFwMDZj5sapCG0dJ+xl/6chEzcrEdlaiUrAcT01O2mJIGxKUisMPUEVjI9O6EoOGiN8OKH
lBKIp+87mgssdG0lbG+OIEYscFjGPDUjJPJPn7uXRmhapPhxB4GDWuDZyqOM3tIf+uExqkETpErj
p4T4vAtsA9tox0JvUsfCc/T2lhbQX78VyYWAL2Oc8/fUbbIhc46BDSngSt/MaP7sv4zYrDZkqKs4
NlArVWkz89uyF58aNASem9mqAMG2fiisCWQrFVMsBF/WaeVPaAfyZAAaydZDrPQzJ9UODS8iyBZQ
4dx8QbgZYY6+3neuv0OuQ3x4K0SfojLECyuV+YmQykOGibFDmfBCaC78gHW9lzygpm4sIo6HbYww
6GZ7f+opVXV3JoP6odSq6kG9x+PZuJu/14lkdL+wM6msgBzbvT8rnd/E2OKq7AOAI6sVg86++Nhb
uLaNa5XnmBJeEfh/pyWN0S1AUj0S9wHGXbmbVNzcvBp7A1CKUxiUNURglKDYSx+rOn+ChncewL/a
+XwBK5C2YpcLThlDFrVCp7FmE0vkAHq9xu4MxVcu3CPWZR13QiIefgJR9tlxe77QAmiEud8WTjbO
tqj6oYHRvCdifPjN6A2iEplInZhmlHs28Bgv8XbKF8MjwH+pVeeHNKX8Kr4oPAgIHI7ED8ljeG5k
R5+e3NXfAuyg6bmYqggXq2SnVpnBHDCNwKO6mqoYkUnIKb8QVi7K6HiAumDqSEGW7c/pPTxCa2zS
gAGqy5gat+EP0fcA/FN4z7ZewGLLDdRfq4brQWp8SNGJtjpZbF23rC4JdCdTkGmFl7d1IloKdvvo
t1IYLJwx1mTCU4n/9GrklpgoU6zexhEByCfLutHxxDltfJ57lC+VSdvEdTvJSCDLaH3z6lzUlGRp
w+xyBeoUrFSPxV3rjWFdkH53F5G8AT1Mu8x34qs0pLzvxGt4cALe221yYChA9qiQrJLYWJ4T0Zp9
vR9SZkZi34rfll6xfBqXtP56fvruixyjavEbuOxElFl+lE/2Rp3UbNiA6wsG3pG2y3Go+QNwADPb
LR/mE/Ko4wUPV8rAg5O8Zxd67mXMqtbFcmlksxoOrt6GGcq3ken/zbm6xkiFdvNIe8Y9du4MKNtU
WABQUVdOWZ6OH84XbDd03uTe5rHsTvQzZQBb9lEZjomlZ7Leq5yUkusbO3uZ3B/+yTbHGdtafjAh
j6Q0ecR2cBXQ9whRoQpH3mVu58qPLxbLjQcHlCgJrdFwJcN6UPFBOnXEZOZQPrynala80LuIONgb
3hBQ2ZK97E8B7Nw5PoB39sxnulMQ/2PqiU4qSsJE/KG/dcZw+5i4Il6wVffTrnOzyzbOAN+SIp6R
IQwnz3zEjOKRsBHyTJ6bJiaNtHnBaOgp+0B7+y9B8dtnD6xCI2I9eYsJl250dchiPmSWU1btkxMP
jkordNOcwVqD20jFwAxIBfEcyO6fn70AiAmYZLODsdT6echeqyXOo8A0fcGzDX31gtCzsdRr1SfB
gqdwMdctKyAeNs9o6JC0by+FUDXhCq0lEBeZD2vFHW7GoR0wwNyfRgGp7glnGzV6zAVRu7hw7rP1
4DJk7+SnKmeLEg98VUvhvhQUXIkaoYfEDrByHDysnJs7W3vsRhSfm+ghsbSpTDpRQussmBJ4QHnd
n+p0l13dn9AnD34UppjZOCHBNT9KlZm4cEMUlDimwohM9e0W66y33oevJRll8NoUdTut7Uc/NcEi
nehj/ZYCFqeyuWAmoMkQ/hTJJVlAZDTlhli8nA81ARxakE7JlqkACSisgaiTi05E945+XPwrNOZ3
avp7FTySAhiSIZTPrfngnmfo6wdMQZyn+EhVdEmTU1PVJk8mYci8wcZYxa8XJc4u80UrBF9UB7JR
1E3bgsC7+Z0lLzzyooVM4N/45dLK5oW2UjTbeNUR9pqyQnpEy44b1Ptw6AEkMzPCUyekTXR3wU9P
+AMWmMt8ILLqia8G+O0h1iKfKB/qJVwYgswvWm72QoFSp0lujw/UihrwcN0+sTJdFDF0OyDBMOBU
0hW+a5FhyznBglNmfVPAN7EOhiEgXWpZBr4b9vl+ZHoNx/um8rgFNuGR4C86WcKhpPpxC+w3Mn1o
waou05Scg6OMlPC5uixD3T+R9hxEv/Db/TjuVq97BLcgZzYdNgRixf6rovYs2Q3rmWJcKvmuPDKl
9LfSb3nZlFbfaW7mB+42gsmu/rP0AzUACoy5hNnyX3C+D1R4qP/oWAkkoABcPZsSpc8PjKNH5iO5
LOQp+VdLdHAmkjfBnOpJeCPewQBWkPYMz8q1UeHIYEtffShayex9I0hk3asouzlZzAMwRVbClnr+
iEORrj5Cz+DDkIaVobEAfHryzzhNsZ0rHhkTqhXWd9KFb2ZEveHYCO+Hpx7odwsBqOxceP0RXUNP
eF8euBg6u3aEh5ntQZ6Jf/zPI4q0l8/pdHN9Y2ZAMx6lTcemMyxNqMkJDrvCUvhkybzmlxdw4771
6biRmUJ3gVC7ctuFDr0LhNchwE6E77gXjllV0YfECGhh/KJZ1qXl1RWr7MVcGp4GXEPcrD91ofIS
cGEp19oboN6NJbrv9+g2sh4StE40z235IH+SzT4haOk3yKdtZndxVyQjXzVH18Or5FQsROOMtDQ4
HJtxxZZQeT357h4LJbRGGeu/65LS23qgq/IQ8wi9IdsomM601FV9fQ2mZ85TcVggoHZOLZ1Lmruf
5R+rz+93ICARvuXX7dUK1JIKQMzGnplMcDZn6wICfhVGGXrA793tfAN3vcDxM7QIFleUIgY2qak1
onIms26L/TqY73RR9B5/LqtvCZtjdq0wa4xRkYQbrtF02RDIkrVax8x9d2KytooHO9j57YSkfvdn
nye8Ol/+OxqjIaJvHAf8U1k4+VnYmVcXUhTHti8Tq1uOcwr5OBfYY3zv/LPID7kLkdGPLtDVrONd
ajiKpWzOz2Ql1HXWQtpor0xaZGXwICsn1Ldm/cFqpi4HDdVuzqJEvDKvdSYHO4LLaXxUblIX9tfB
Kvhf9CEQA2h0cga20PsuhTHKvSQQGwkgRvvLF5+HbNmhXgTXJikRv7LwyU6CVG241y8Pseu+gJNk
sSivCCXrubpPCm+L5IGAOvdADFnkIf3/xLUZF78f/uHhFTefIK9ibKkct7ZCvYj/ZIcwnqZlRSa3
5AmJlDsmN8mVtC6xvy4iR3Ay6lPaR6yB3IATQAPeilH0zfOOqYcXVdFC4+UWXyOHxF3Kro3xs0QQ
fneuMUH28Wk1Wkf4NNDn3+MhBggTcGZCkJlXIhnrG9+CM8uMrPdeuKK7MbJHbUBgN6lSfARqwFbM
MsIHvsBrtE5Znm1GHbpibbHc5fL8LDtrefb1k42esWqsxFpKkTCEJ+xBC97yUreM1jdbEX18RmVq
vkMnbpSj7CjFpPE3x89jQtPF1ywE3SOq5Gn6x4KkiDamwmYL2QxHh3uCRQV9BKd/lJhyGz3gX402
rWd3hinzVv9RgGhM+WBRuB11vC82PSE5pNcFxN54bw4JVXfl+TViZxUQpUeQwaCcK9f3/ctlXEYx
OTLLoAumrASSJqSPqVB1Lko0EKtZ/sY8/0uM1F8NjO35t2KyhlEBaSvHv94rS4b9HjFCXE+HbOVJ
Q1SheBH8vcGKcuzyq6W9A7G7oWdQ4WyPbmqtjyr7ekhSEIPl9aWfwl4oyx3McDBlHuNlipabPbFN
lrvDUZNB/6IOPNswcXeAURuynFKwbcUNjp76+ARwAOz/7QOzrTSiCon9npSi0CBzJ/GAXgGghtS/
Y214Y85hi3dv6h8A+hwMtbElRAB3Xhq2CpflynRdx3EH9GWwhtGIjgznb8tZyg9Q8yDpHTYiqOoV
vY5fq5jz1jo2UMvaQRAAoB8KctIP0CbDbOaUdiclwfKeeTVSZNWSANud4s3iASaBEkWGuy7B8zKb
0o8t0PfS/FUsJfXoMGaU7EAYPAcnSusf9raLTB/z28n3DXHEbOLomeoUelC7VX7ZYUVfyww/Z1r6
n9LPAbktuPkc4GFPyGHvZfr2lr3NoJAZpX7dnnsDrdXvh47AXQGtBOYaZyt5jweF2ytwakdFgfjH
b0BvMObO1TDP6vT1/f1TFoO8qbAEopnig+E9Dp3WJ0Ycbpyv16denJuvV/XAo/dUKIhbiqvHA5h3
sKk2YSnQqFutxoNhyCsW6tSfbCIMr2xL0GHDHkP8GFwz0vwhlnaomKSUFj41ChKiyxONBrKdY6Yz
00QolqsD56eY9FSW+TAMIqoQy0YtVY+NMUBMHgD7DyGTnIc7qOg6hiUpnQ0KANULgK+8UCqzO74I
GwxkNwcrBBojGyjHZWxHoK6kUhcqhCPxoRwBPYhbY6xkmopzeD+Uf/baQwwJ3LVgYwNgNqHhC64h
kdZI6EXPUiZY4yILO+X/6yBcH7MBerOv1cIyWRqN9paQPY4WGeWrXn0UIVlo4xqEIO9U9PXTbCcA
vOH8whwXvKwpAT0YlXbE4/HNRCpebQvuf3zWCTKzK1NSWVwlVzwuu6Kz1iX4tE6z4r8GADmC44Xs
x6u8ZOxrM6tW7OUBsdTjQdGoL/OGhrPSL5DCv4xmHkaYdWWouj+inpCeCHa2VZ3Gg13lv/GFcwHl
V9aSR/MvDxKZUXDtIDPmuwLFmsOsDyZ9wTJxCN9hrqMKI1J2LxFyLaqXQqb2SuebHrqsuX+w7gSQ
65RYqsOAr1BxMRKMHXRYNZ1OdNzkreGukxJa1zfrw+7gNb0oHfvYV8zgqoq39j6XW9V159tvqel/
sGkNEtvwTBlAMMJv2wnXYixKv8ZeP+2GK0hfDgrTH/qdtLTSrTdgEAbnNHCZSrTylA2x8LLENq96
ED+eRlIlyjA2s1aENXsJbtJG7E/9JjOtJ7DtfIdMEBLzlbgmGqVBSDRAj9gqBxPx5SC10dJSVNoy
gvb6WM+BRtNLWnEaO88b3WMjKUqegUST+Rv2VceQjgrA3INxn2PuiV4TsUjB+sM0iRvOVk2BXe3n
z8f+0KMC1v+kAeaEZYMI4to8W488RAN7+HJ6QLUEQGm8jnjLty+arVnVrd3yOPQa1z9vxmJxP9Z7
L746bJWsG+6Kvb3RlO4t2N0FtF76quZBpMgpQrInI5ezkPkt8cIYr1RTM/lXJAololS3vTtrb0SO
VmUZR0u2E/mMV/JNDmbBzOE+E0kIqO83rjGPLddXUBE8vXPzhVQOqDjHdMji6l6C6rYeZ67NLayz
cmEAe7Rj9kKuaPKQeBTD0B/ajie3tYEC+HsJ8NWvRevz9ZSw8UCNv5DxrgEZ04mMdbYZntjPhOgy
z9hEfWQD9kTZ9cE8n8Hca/A9bD3iGb95VcNZkRiYojrXXSNM7bDUybrsLdkoAFCIsqGWl9X5XlLS
XA7Yr6gZWpp68bSsm5N6HuG+LWy3s6bQa/lDW/MGy/a+gw88uwWC0tCr+QoMvuWPJj8m+QRnmxMR
rDSX995tbK2J0w5YlTHop/7fJpcodcy0ERWuvZ6miVhdnKL0pg+4kKhUiy6POXHaIl5rHypi36qJ
R6EoBA6x6ozNLv+Om/RrDqFyOvUN366PzM3ifRPkeJ1LX1xB4RfWW9HHoomqCD6vNOMHSdmIY9nk
A4cNbLt+Qu/ijfISphgoHdSuCsMUZFT7Y82onMCfrdXO17vFpifrlSVNxAg7P/S99FNdNSw368IS
HkG7NzyUb8OhEG2fe0t16gr3zD53oKnLNf/PxsWD4dfIfOCSDQXHIeinWodweFXmAG3owlYxB+pO
hHLZ2OHUJsfbZcGHbKDTKyHO03d5/Q4e0oFgO4vQQyStF4ao7P/OLxreD0R7asvy+8wtugjcOo+H
IM0ZGy7mPP2B/7AjDJAaVY3UNQyzp59YtDdH8v5jV+oJahV3FHTcXqhgJHco1pX1jNfIdFpahutw
5zYrPouKtR+qVG9jyq/eQsHh+AYzdnJKWR7mMcsPXNHySUGcRQTGZseu9Ok0mUcIarCGMX9A1Mpl
P9eM3pHru5NaCe2q/0L2C64OaIgdr/2yskxIDxPJeHDWColY3hnGuUMPygHKxdoMLnhjw4Gp+13y
lLyS5mIQZ3tKaemdUapg/k4LiGDShCiJjD2eX6Lj8WGbhEVgCCXypJ7lbUOKPr1KUpsPVJgikXga
mq/lkyw14EhRFzhGnf1Fu6nxtZ9K4XRuBhuqdw37MMzx/y72VrhB2kGRcZBIx/CD0rsEdUM/lgnk
nUHWTLEoccCWAV37vTdC3a62E9SQ/lUJtfLAhBrC9w59Zn+x3okcB2eCarHHE+3wv+gVc3xwTFOD
lbfhYlHrHGxgQnu0Ino+BmfbvfdZzgFnNE9y/uryIYHdRQnkUOyP5n76e7F8DeRnvKMGthPeiHq/
lFlQN35Zq9aDO19jwT+KsjzRH96kb27HKwMLfia2uMPmy+msGwnzYI0Cbu1emFm7YtHyLcY3IpvY
RJOa5OUFl2sHJcY9k0LTPpXnlRLI11DlnpUJK490L9mQ7t18IdNcNCKwychAueEGvatvncT6AEJf
V2iS3LkzVZzeAoscUGezbBem6V4W3xwix7UsYxakApmxtHsV7oYVmm0rSRBeGtXWoJneEr8H2iRZ
UoG3K3i3mkq+GzqqgV/ZIaY/WNc4nx8c48O32zYUmY5IyZBOfWwZyjwW+OM2CcYQvHLAWNOMs/JI
JAHMT3PVkHHY+LcDWHg6baHvW2CQ2fE5hNrVCpKQM5TModAQrOEAiTdS6aWOsTXZ0RrWZO6F/n+w
CgDEsvdaZ+obcDO4qJ9imutwSUqMFqjXQZegiKN+zPLLE4PlctI6idOkgQPY1framTXVXLxLg090
QvH09H7kEG+Ajd0cvMWrnSKGnTCJ94k+E0mwsBhSRRZxYEcM+IzhfK7L1KFTzR7GmnfH6vbkZol7
11S3OPFP2AY9D37c1GkScH0yBCcywJc1sFRscCA+ojRmHJhG2np+bKwwtaVekvyPONQU2TUfJj+q
jqKZjPdSeqS/jJFznwww/l9W4h+IBKZsG2WsB3PoScSocCCVoWSOZuTj+klR3dsUcnsB+7S9P7Mk
EoCC2rbIzPk0o+eltOzdsbphtFPpGu+CYUimrXSgNQddbNLfQOafn17va6fcVhF2VkClakaNTkh3
tJYp4lxX1MqZCxNHRo/Yx5EA3zoUcjSJ/FuEGPcP/psA3XmgrDtAxmlBorj9dfgwSXi6JmQ/w48p
Sdo9WnHUTqhMV3TEXeVABw5LXlkFfq7v6bNmlu8O8QdfPEWjPT/l0UYPY81SUkHU+raYqKxC/fFK
WfvMvqd3z/UOwFQbOjPfgxiVyBUq8Mr79Vr6qVuJOSG45Sb+GLb+j7Gzug6bNRtbva+7OUCsqqVA
Oqf9fk6ph1Z/Yb/ZvaaBnxsnHc19QAnOXwFf/Wzf7k+pbgdYP1Ix1UScoWyBtV9qwK3TiHDRIVwq
Mvi15GMm+bRDBJbzQT9WrhAhmJBZ4BW53qGfJm+Li7sUkESMUS+tZiygdEAMOHucA9vnMZWQV9Dy
6ZjNQUe3aQAaak2y50h/aPWuXTWjLz5lvqptsqFkMLWtIPfhVXZREdS/fQDf/rrzczjW8axy51UD
NSzOdiUZZjLlg4qC6lBhEtsnMLvMMynw2pS4znsLwZUZxDJIgN5mMoW2mQmIZ7mkz34Huq0Bxcfx
uJjVocpIx1jp12/P19MTxSCVyVt2pV1Vb9yo1ciYUEhhxmyXNoAjrPXzdBIuaG4qxtOVGjLOHcgc
jzHfkLE7UAq1qwNIU7e+/SRhXE7vKHilTY4JbW9kwt8grOe7TXWAMIJE9TuXX1P7TsnXom+r6yDz
mpe3fRsf5xfxazer/hg9KWD9r3mRjfot/V3AWpPza5MK0IK4S9wMTCi0DRnk8tcyGQfo6IYX4h4K
Vd6mMgjkEjo6X18+82RMLaAv9uw8BHergs3HQ8bQw8Dud+LWZKJdmbNu5+ZWO8PGZyR8/cOT3JOk
Nf8efWQJZr84kmCfxGF/kVveFMwYgmyAIB2X1fUoI6hVygyCPqI2n1FZX91Jpy0+y17FScpEauFt
Cm+AnvYTb3t+DnpcWMZGkrrjAOytWGl3NXq4Z3hVPtLDbWQyILLgLuUVROCMjuQspWuDhXzXsIpU
NrJvTa/5JQQEHx8st0AHNesxuDISq2lOk/U89Ti8TVRP3Oc+lKKmA+pe5u0CY4zOEnsY9qxwjEOD
x0fNVwcw3iFqyDCcb0RgkdS7MzsjuZsSo52DIZozEnz+dtGLMqMNlQOutNIhXitPX6NrTlLKjWrb
/xVFHynxZ92EMjOHesCIShzDOxXEyw2vGDpCCkdZRW/woOBcIScZwx+EfA8sShVnTnxjG0VZF43z
184wBSl79F60mBepAfuHLkfzBuV562551W/rd4Hbx6YQnVqfe30heKgeJPcjmH4tKkIOp/RYys8J
VIsLemuQt1ZyQOTu9kW9YFfbU9l+dZHGID7kHZfrI77biDZ1oFpm9NUNgt2L049g06SEU3noYX/f
Sq+d2tjD/TynkrnNrPRrH7Eu4wQuFVX1nNumJaL9ejSXZzp3cjBssre8EzvXsOtPpX09ipGodJDf
8B1nYQNaqMUcg3I5KqSzFuryIxY+sd8D1JoN+9EICpM4E9v059xYJtVdy0ke99zxUmRPAVpHaSiT
i7+uJ3TA6QjeJOrVwZxtoqpmhhfy1W0kwGtMitOay8Eyv/x49hIDeaLGx6fkbsWJuIDintSENSiq
dw7Bnycn57E3jgTFtb6vL2XQDWN0PcZHkrcFHjQniofhABz3CQakf7bJOHmFFWSRyvBhS626ekh5
1qn/oMwvZJwPsiEw3oLicqeQslRdP4VPyWpoKhy+Atwux5k+FEowSV2pLUTJxwY23Spa5iZysgcQ
09kMC0cUgURq77RoBfP40mf1reXAphef+Fo+PcmsT08bXRXgMClFZiUk8TK7oPvwJKIewbal7BA+
w2mwQf2EpN1uhHLU8js0BvLjePQumo9EBUAfcjflu5nPdwmFTYQSc+LvbgOS3XKM+LnpRNiPN/Es
tjSLLdMaWXb29T1BAl0TxkS+2hb4C0Ks1kATlnxn+HlIaixTbTKpqG6S3ljYk84i0JRv8QjKQfQR
xIAaOmDc5/CevyTz+1hQyWZ8t6OnRtZTVlQ37VXXPyjIarpbeDQVYQb9q671U5N5fVioXAfdiHP4
gsceS5y++ZRMf1rn21KM1QV7CzjF/cr1FuAORh8JVQmx4mUcqqLn09cSKfgvFx2cjSpaGaZhe5DK
SVG4nAWrPYFqmFpnrcMk0el+TH2PjBREkKurrU0wHDOlTrO9l5osXbuo8M7Q7nAJGXbNozWImC6o
fScyja/bUhrEU5jAXii7ThZcfahT8LIg2GT2g6d9PiJh4EI1dOgsS9okrCwxMw4LsolpItblUn1h
m1vdgFmDVJGI19dfuVnufeKj2Idr0+9FRxk/f+SUSNTMAu1k5Dgaiapu9zE0ojCYcMD/BA0OoXdV
fNqI9MBGoIXI0Oqz+0k3275ogtmFRiCtgfYxaREn0CuIRqbcXegsVHZnT71OmKTrqJ2yUCXNrbFk
PGIqyE3wkFN0MkxTkTbWj9flwaxFitznwVubpcTT6ZjHV37mBZ4romcvGeXjNe/BZfNQYdwDixeN
/slGH1XTCj1PGDQyOk5AGqwX44szjPAF2FvNnfy1LMt4QuVppAqAmXUij3AjVGxe61JoFYOfENby
O65A+3c/YTofQ/XoaYtFvMuT1NoAIKbY68TtNaxOEWkCGMdsbxccEhvBeM22dEfF7fPZOl5aQ7yJ
VWsnpbUeSm15hGMb8Ui1ATk3yRFb/6YhGJEs0EpPkjwo29/bgBHYnFnE4lBfwXN1aECFUrNdCGgO
Fg2pNsPfkNHK1cSry8/x/QbBNxr8nU0loEvjk9mPoeXLcbYPZWhatIgyao+tonZGlhqq24RPQk+h
29XM1lhO3OP/BUoYIDVS9/73WJe3E8cF4tc79x85tCSTRWzTpZ+7mzR6U2KcjT8WwqFP0ZHFCism
vQOKXHFGAsAj1EE8bgNsgVgheZJTABeNWqjOR+FzQMJHEdcp2rOXyHKaQUBvVbUhjxbKUT6CC6Fh
mwe1FgQUZwEGN4wXkbXuZL7GH5IybwUGpqhZkd/nrHBN5CRwgKDkvvC/jnXYFjUxRmAcHbOy9lw2
8WXFdFgVcNa/P8i2PKeT++afqsmkgGta+mox5b2ivgljmDKVCjBTStFgWIIlANGT0TiS/tRGlgnY
DrikgybekFBWMPYtCXRPW4aL/BLqIVvToele4f/6QqV+7HvAcO2Ryd5+diMIfFjIf2LER6HlsHYv
ZAsQxAfeequniQnpZ5mZ5tGg6v45bb7lBvfe/2wO3UIwXfFfA9/2Fmqw1ggi6pdFeE0rqruSdEOB
Hr0Ymj5pX0bw9eHvhh5uxem+nHeTpwyHCtNO1ACqSqaSV01qZGuOaONwiroGP+3B6HEM4IvSE2Ay
jEkeYMwqbxwbq+sxt2w2iu5wNud+kL6UOUjLA+m+RwUAWLnTutud7Ate5GZgfN4D8HS4wY6JwI4m
IyqrSq/OKhiHdLFdcVa9SbEQCTvOSrbSwkX9wCv/mhDKF2ZrKD+b8MDbHntqina560qGM3IP5Tlz
Pc7exQiBwYg+g+fYlkhnSNjJpy0nn/OxLs17tGxm6ZUq7V7SHBs+MQPUfo9cnDrhLfVREeMHWFEt
bgXPrPE4UUMZEWEKiEGgJ0t5BjU77cve1XAsW268pwNWAIGmGQY0FtteJ2bBBAidI9Q/zKjXCP5m
lVpUG/cStuqgEMv9/SAaGwbLZmJ6mjJhUswdiUGErIsylr0QZ8Zps4YCQKqi+fFenLFrovFAiByA
Y6c2zsoNvQFcUDSDEQQxayBjHZ5batC8Ii4E7A38dTbT+fanM+0hh8pH3uiEWZZCaRMxZ5U9JI1U
sHCexE6l75QonwaoEYTNqtgxbkhRz4AtyU8UGQeOzKMz6cpa54tSrYH5Z6+lGqfX7hgpSOBFadtp
Xg9hB3MdQl7EJY5LUzMtXerRCRpt32bPR0La0q04Rc+pjaAe/buxU7phGpoJFxI/UU1QRbN3TH7u
OI/J8QQHVqasiVEsLg/9FvKlf9iRZrIfoPzodemXrVapfHuz/3rt+grAMtrnjqlrlyYhoDEkZjRV
B22lLJGpZxn5qC2PHWH3o/TvRf74P9+kSTaPwMM1hb1NgfeKDfxBDTqzq0RpFW/RPAgFd/80Af+B
FBY110EWG2N3Wv+N12jaaMZ4HlS5qkvLuXZBSM9Vh5Z0/jUvkpebf9Az4jqQKkL9a6QDRcrDeKSY
AV3uw7jZ082VLUu0FrtAxrZTXqsAx9j8MaDnZ5sbqHdm+wZLTBJeEhmhylqZx7QkrQPlzNdzlKra
pUgKCdP8GizhuG99LrGD+XIS/9UlJZT3rgzVxn9Y/V2PaVt3SM9dj4338XaEzFa4+RVbvTAK9l5Y
Tw8Wa/wk7xbEM6rWSjMfdlt5PW+AUTxLHKNrgovo8+xJyqce+2Ii0buufIA6fBNskUj+pVpHtIsJ
2o1A5zlCpeaQVm4NiA0x9QF77NH2giaKdYY/3DK5c67MB/knWySOyiit8n1hYh3CUy39DR4y2Uyl
3uS4TeIHEQB65Lp1r/ktDFoamkUxdC4bqP0eKErygW/sfTi+kdBiScHQMFqOrK+KP/ETZEEoRwQl
c3gqAWH9pcHAteRmMnAxPpGKLSJLVCpkPWyN8Rdft2gxv1CALuhYTKlYVgCmvxw8P05UbGm78bEm
xEl/GXw6BVGoZi/R+NkjL1HfFCbvT2+M2BEcCsunrXwFPS5xgAk9bz8rNV13laB17BQxNlsmAF2U
FNzu2XXp7am1GbqgQySKUkwU6WLP1SdLcn3vsGkTUi9qKAH6X0eOhweOP7q81fYjXBkHRhpvjMJ8
0z75L3Xedg8+cdDCi5NNT2SYeRpw/wTUiHWjjwqwSFpM5Ke25DIdyx3hqnIpzYOHu4Y9Hr4B1rs5
Jt8GV8YZC/suG6fx2WWffxbNxz+x0gva1nIvfD3sjemMEDPKtTbE4VMNJ0DWKLui6/wdh5YqJQFO
vNhxvaK3AZiV/9IeSxL5XMm3lqbnWP00oJHE1TQDi/37t6YnzLN3iiY6aCvDSDc2BVzoBaKJ04nM
XN37R8Ct454OZJRRdI5qmlDkHyfXKgD+7ccf3HW2VCdFa202hp+rf8DC4mL/g49Or9/yrbIP9amU
VGRb/Ndt720XKOCgkFuoCGjRaTyY95Vqp+xxJtjJDLRdQt8eEFbwUmXIQG8bs1Ls/GSasQwU1qoe
JjqYPAI4WNZrkV+BV/nLH9kKNm37CASrThEBQF/K3Oo67IYyqpgIRNj02VxQisxeQMK2iAT+vTwm
l4AOmsBD/w+DwZ23zFh4Yqx4b2PdC+gBIZ7ZyudEHKOOcuLVVNjTk1PwqqgTQwdmbxqU5KLCM57w
P17AdSnE9lK62n8txYkqunADF4dqS6ej+miMnQMk8PmX3EivSVJsaH1kisbKuTYxLXAipx1ubGa0
GGWQrMiUt5As7+/ymRgLjVBU6d/sJu+JfrwKa3OMrlp/0AY8faPdgXmUZVBn+cIM8o8QgWYWKj3/
gga9/AwxQ/nelaBtB2lYby7BJ4fRa04HlzCk5RbdiZgkhtv+En5sB4/OJDj2w8G8cP79XTnd+a84
kQDGLZqX4bdtHrvpem1zludflf8rXKNhkFGSEL4XKVnFjamrFU2qC99Zwg7HRS4CouQ+uysOQI7S
LPvd8EpCkn1CIL1shT1x99K6EXWBxyadK2p0P6nBQaTqi6fpzgzoxj6xJuYBqYInw4TyHv4QPn4Z
AtHy/7exCTdFJtXB5pFtg6H0xi32zE3SWtJLbH+9sfPb0k0Z+nWHSU+g0GgFh7eWw8baKKtJw4w7
vyQCMcquehYY1hD+KEH+4qu4y9MPCODCRb7kvyHzytcR7dXB5+k6JigOrzR6e0OUaQHJek4aJzlF
hmZt4y2rSanzykObLPKINaocjVg9yxdSqHuhag3AljER+KIQdwjk9IL3mWri5oveqggJUY1izXun
lCw2wtDNOzOT0H1AwyTd53NA3hzcVtF2evARyx3GQ+rGpJA+A34synh7JFP6QhoP3KJ3PAM7PNsa
Ms8hL1PVPyVj33Ar0LN0NO+KcVm7FWAQsgdMpjc8q6Xczu0BpT7S/kwvYIgVBVNgTb1l0DZsNMVe
aqwJ7EatNpN86acWmi606hWSjQBuLfXfJjwGxEHFcjApuOgBaOurthLS3OU6aA4RwE3BKuudd8gi
dBZSJvlH0Wj/A9QT9Ufc+feLWXdpuczoF1E00loCQsd9oNab3pxQeIGk4TR7SWcLWLdxItKn8tWj
hngkpNaphBiwn0EA69MpCK7jJKDW0AU+fEj9YniuF58VoSlWIMOaILmZT5IToCCFTfFf30lxDY9X
8+HeHTtc6YLWymBOHlIqaETt5iWpJ4x/Wn1bhSJeX6mJkQBWx9QL8EQE8ymAJYgNSY/81BKRopGf
frVcxxZ5I1DiJQIktesx/uttYCYf1seLSJQriXk6HyVjGHOOkyE5cvVGoWqgIVarZXv7lLx9Qdcz
mJDuDO9R3CN3bqQuKNcScjhbH7DWPEI9MdhKRknLXU0H/drZ2XDPVZYCzRKdEOe9lKO4AdrCl8AH
BYyPQObXCXnr+haYxt8CMBdMzm2NZfnzaBGLMrRAXFyN0Tw8NckjqkUgC1nwVeaxBWfi7u2JRir3
kl0UnU+a1ynKwfu/lv7wNr7SBacJt/5F2g2G8DBom5GoLIstSMb1f8jaYZosoPjgnom/ZQek8LqL
uSzeu3M3GNZaau02HPfaOYn5HeFXnAvQJLak0bp1uBHp79YZWX8+0xYw7ChvzLoVHp7AUmafryYu
RdJZnfg2sgf2nEdC74V3aFvdxhRQmsvwDPoz3ThcQnh9qgluNMFc4iumS5Egli9bCZ7UTApI0h37
+oS3RVu7qnGFPqg20pRoATtuQzxqNxXUOL4Oyv+D9pEphRh5u6XBwhfodmXUG2B9XYhOzEWJfScU
XYD0RRS8cs/yGHDYRXN+CjcmUfAvPFWh5CZSN10yZme+xgpEv2khmS9+K8oi8oLZXPA2iytX/RmR
ylID5/q8B/cig7U14IsESyKjOozRw0SDchE0/6+7iNrM5N3iNiqXVj7o+oEm0l00ct9wr8BtzXBK
7PbmPoH4kmhCRh0oGxFTRBpiHmV8ej+5q0Q0kvuEP02Uio393ePmpofbRXoLK3xQxIm+cBhz3y26
96fG0TGSWJmbNs0l9ej0ofvpHAZqQcOjbNL9u0cfTyjsNgTg+57PTkKtJGE481T5gST5rS9rqd/Y
8X851Kra3q8bA41dWcZL1bGKoT8b1NunO6sV7Y1CULMl9THKRPA335byupvrlzMWLUt8cd5AT9sw
v2Jg1ZSBcPwSYAoSJE3lGzTJwxT8xqqJkD+nFveUbRXiz6BXxFeLp+YOZTfJIdODtqgm91Bz5JT9
f5pp7F4CFJNBirkD61Jd80evTW6PnC/dV1xDnYiwibB8zlvUPXZ58kzees2GxuB9MT5NtaSCyLQX
3Hci8HUikbqaflFnliGxkN23dS9RH6ueTNIGWEBexorD/UTAaXtLM+moavmPSEQPSB5TiM/jB0Ea
14Cs4JuGtG8tTVCY67pyVc3b84BiJGzVs5og0LPAxorr3yz+ZAJjC25sW2plSnMpJ87EHgidrBtW
vl21RtVbRh9tzTzra+NiULl6H9LH7GLiBTe8eAkuzCp1N7MkqQa0oB4yq1cM2FwEw3+RLYuy1IvF
mWnxUQypFSqoXnLzPW1IdAPxO2NJhS2hjxlBgEV664Skrm8j7APTcMvIIA1rygLgbf4hzn4WIwiQ
7fML12Gv91VDuBPyl4nYh0tvSTJIsAa85G1p/9v+rXM2Ml02tDh7u1kjTxZ3OTgrUyoVVfLCCsh9
MP/DU0hdnJenZwrN4RFqAu015EXnrUVVrFYctaVJeBbrizcxIo3h9NsgEEds69y7QG1lJYNRo6Dw
jGaOcv8FvsW7yAnqaIqSbcl4HYU2mg/J5B15bqLiCHSafgo95HqBCqFqAHv8PGYDVasp6HKVWD3J
qW2nTiW+DHz6yCWE99dX4fMX0mPDJDygxcdTF9bHAZIQI+HkopL5NJDzb32bcAaCi2UNJHu6O3FC
QQVarqJChPG9lP5Q2TXdeo/Vd4NjJvWVvTMtz9QhAMc7nmQbQDB0s/tTshZLLXizgXUH9PYG0FLP
y8gLZ+msAMuAVQ6xHn8FFELW2z/ChdYMy9opppyzKtngtF2e1n1OqA8BeQ76j8Zk4Af3WgH4013O
AbhIyCFJbKihR/zsCGy+AuM3dk/bqwtyqrxcOzzUXq/g2kyy+K6X5SbvRFFGD1VIIg39J6MAPaYi
IrL5D/IfM0V2zvTSyd1/oIiAQhL+UYPqIhkYgwuF2HpwE+Vizn1y3MQcLNukmeFBMkT62Pt4JIBC
BeM46IZf39pfGK72qhAv71IafrFfp65E7wlDvtdSRsDgfremAWFNwszMDzzo6MSPoKawFvWBH1zh
fKYDwetCuTV1eEGq6sulcUfK08WA68BPDKM7lOzZa8zl5OmqDHMvYCmE+b07KqoVX54BQfak6ybM
ysM+ExIhF1R1b+uzkj/La9EMRWa2qk/uWe6ukpZ/t0N6pi3opCT1mvx+7ezXgvZNqSbV0Wh2S7yd
FN3ynwmQcMKS0FuCBGGZHQ0Pwd7LvGjKAxRkp6Hui0bxYcx8kBQ/FowpaLXQnFsIfjj8ccYlICZN
QqdJhrQQoB0V/E0TAOQ4WTFqtSvuqwAlJfJ2Jfk8OUqFc1Ikr8V2qLkpcSngE4Il0HnpsABly2rF
MCtixJIRHeCnVXymuDFNP3ahyfeq582lDy/6RP4/rBsGiw4pG90k4LzqhNPveIBiWSxjThYyfThm
uh02UD9xkSX/Vs2yO9xPte4CMghcp0SOaqNeeT6fVNdyJLu+IFhDGK6xwgyRwCkT5L/rZB8zPInb
8o90fh6/3BxlWoFOkk+IpLOtBGfZcsEHllwwOuxtYSok3EgRepZyBahEGrr2bfTpQGyiDTa+R5g2
45Mwo86yZ9eLhqI+Y2/TLIgcqFkO6mxq7m0C1/eo7f+bxCkr3QvW3vYb5sDV1PPHr5+BI3AOF7r+
EhO9IgLQQvhLfndjP2dh5vh55JGNcbeMJiKqwEG+D6wvwywqTUJ7O2C/LYdRBBKP8lpcFPPCXnZH
lkO0j4QqfA08hU2AXv2h6hIjNjd9aAm+h1SF8idDHHdhbhSmTX14Er8Wx1V+eYPNHWRbXAUVKKDW
nkYGKnUIfRtDLLT9CB4n+qW5lmPNFZZ8BwAmDbsKy2qaGKQsluFQOaCQiJyL1ZVX0P9q4vuTxqUT
4eZpgflCQKE64qFNUJ7TjwNfFV5R243xhXfSL1GRreVLb4t2fKhx3c3Mv8AUTSfmqfmZJsr2CNS9
liDrX6g6udcXQkelo2Xd+SKQGf4IeyS60Jpx87EF1DgRdiWPbEMtAfaU8U+n3jEv/2tEnvbc0PeU
IjcGRQVTCEXOoGOlYXVarHrCf56UsJN5oqdX84zEscUGg2FWrYFC95WIkLH8AziBmtuBcRu8gTMg
jxw2XIuoGgKMPzRWkplX5K2yIcw6k05mVKENY6nHVo2uAJj7t+DJAAWhii1/pfqUdlh/kAPycubz
d3htfmp/MipCPhX7w21WZeywkA808UCXKNODXKeKAVybw4tCE7iAp8gT3SnXJsBIbxVkXQPebxnw
wkCBi63inCPYQwO0Ae0OuSZTjLB2w/aPuUoDP9Uf0BYBDu990AmebmXngUw4KtvT/zSWJv/zWcgO
KzL2nxYKVvJAeslw8TE5Lc81DzvZ8aHHu2P6va5YrtkjrGyM9raTAqmowq/cG8dDVFzq4LN550g4
zGWg32XK9/jeKbLs0Pw8OhZkT59Bq+SbX/dNfH0lNVjqqQGiSGHxsoT41ORNKadw4UK6XhzHeof+
I+IhIUHjAqagnjhpBe4PUPMtz6uEgHwl+P3Up3J5FNIwlggnViUpdRO6PcMgUOX4pSyvAN6F7LsK
DQjzSNl26Jtf2DM+iFCGUdYjz/62TR10FbeLwPDA+v2UZ01UKs+JgIIWoie/K9MHcdiAf78szPLc
NW8qKE0bzIzVxRfH+2Bh1mMvHRQWuLkvhLW0OpyPSkOfeFx4D5zYhko5INgq9bROv9aIfbm7wja1
+CMW/jjMouZMPfaINIaxpYHaIFqiZAj2Su8/jhJMplvl+vVTrZ8mPeENjaEZt52vD1yXb5T7jEGB
TRo0OBW1T7egH1sm3alzaPlkAR/yXuhVK+5pfFILloOAaXwu64kkyWOrPQ7P/xKMY9ZauasaaXod
r1Z6XqhTnH6o8StU8FUlHR1WCKYutMkyJPY+JPXojmjdI6mwlA3EoO0fANqJ+3G2MigSiHVOSVUk
Edq6MaItvDWw/+POyc6KFQ4Fn1aMAkziW30mZaKSDaLL5/5sBEt0DBzpdjxwkpmMt4TZFACmBM48
++hpSlzq4x3DQIQTylXTRlJUzWwRdJOmFWFRcOsk7rgUGrkYKimbx8XjWJLAhGgeF6gh/HL7dMRO
X8re/S5RvE5+s2kC05DuaR4kADcgaW8vBunmwImm4i5s7ee9t2HZiFN1Sl5o/9jsh/fcM+b5RdgR
IiagKC4SuYjs/1wK6tWuiPexAvziREF9FvPdwFIwhLYfn+tvvXZVXltURAtc0M74lgWuAy8PTF12
e2+rXMeA1YNlCC0jROE8R+IpXRfsekq1PczK04BVUETFfTXhdcUauotK0RpW3k2xvmPU3zXfcVtU
ifCRYHMiUQnkFqQMsGNkKt1mgmbAy7xp6J/LGcHlZRvzTA6ZznH494HpeUvHfx8uduMGPu7u1Rao
8NyAO+z2EfuNZfGOc7mCAy57aE6kUT0FUJCvkGi2ZODD4jydmTte0oTKNOwJ9XoKZ07D2Y/0cdcO
p0TbKvB5BnRv1F0WsIq3omr5t5qT4uCZ/dThZngnfR++wCUOTKYFj9fM7naUgkBQvtik1hRujQu0
JmxE6+A+LJb0F+aXDx5LzfAbV3Eh9Jn52UA83sZg7BnxUiRtPiobPS4A+Es8qwPtJOb5eybouEvo
cBEN+80sviuMrU9MbQku9eTpc78am2jk/Ls9SVmsx/5IhhXeI6iKx01tzV0V/pADe+OYfFc5Ngfy
NmY7hWeZrVHc+OYWt3KnaViGxkrXQgDbU2oUNCY8lU/Ieev8lxqCVaBmkoWhSKsUZrtHUmdndWE1
EhWtvIwC10v/sni6ndQz4ExFuA/d4LThT1wIb3czMSXrK6rymwGT9EIYgLI/aLF8Czos3FZbopjX
qDnwYNRQZ01m0ksknOjPFwANjRu9X1asGxJPHpaaU7jXyyGMQweYHUbZXd78KmsFUqfZhTo2rFH7
GVhpM1/a+4HkI8tyZu5Y/SA4I8BYLRO+NRgY6ggBWlBH2QDsin2MenqYmhvU6oi7u5IXKei4gAYW
Iig2UoTCc25gS8y67Uw6RZSMDz6yuD/JI+pGWNjo2Lxx7eOI3DgJBsjFFAnujxygZfgzBYRSEspN
PieXXbWJT0RaMzfc+E2KtiRRWjhe/o0dxfP7X58FZjxksb8A3Ye2rG8cA3IkDz037oEKlAnva1XY
PRH27Tm8pAoYv/jfjC+CWOLXku6LN3/UR2lHB9RjBf5JkENG5IeMg3maRwP6t/Cd7R+2K6162O3p
kdk/soYoMQs08XXCY10511boBWFiuM3s0NbUoqi02lGLJDZCHw01DvT7t/xXL1APPcPCycG97Llc
HPpB4hKEeZEcnsZ2LgpMXB51bA2WSnCfDD0ZulOoT4OJ3bCNDUiSpYREI8C7VoFPJAh8EWBeU/hQ
4SgL6fxa2KkA8tWRQzrzzwgB8/zzU1Io5tWcewwoq2KFj4b5r4paA1bVnWcB9kslM3usbUrBIDSW
hiyTY6a/2i3/4XrQ0KQMTNCSi+va2tw+b3mv7UiZHXVpKKn/b2R0Rj4r0jiZ/lhNUy+KM3LcDW+U
YO+tttBz0F0bKAsZ05oQr54Bk2ElnV45zfwl9jc6xqWKwDncY8QCa44C7p9jVk6CpYPXcBoJ8iKo
UrHUWRUTXO/oCXCdX4BkvyA+pxcquB4vwP+CgjmdwpJ9tdSp7Y9jz5BEFNypoudaPs4I1TYcDk3X
NUtYYZKWirebOeTE3bckuBFS03b5O/JJmMf15QG0Yf4KUUCKJKRmJUayeZstxo1BBnnWUgbs+Ugm
rhqy1ZA8B/shIvtN1tDec1NrceqnIDJHH2P8c7WigX1I/hT0y3ge/fvBKVTqez3k6VOh+oAtbTfP
b4VqXNUi+a8EwIKcWSYXbl3JbDbSo86bIXOrGBzVm/HpFMF2Yasn6q2G026AIIgAN5Rw23F/g5CC
ZUs2qf6fAfW7LI41qlX09DBvRe6YW0o2dYpkoWq9ngtvK8YKU8fuq1BD0xGWeSD6MNOJhk6v9Fb7
zhMBVhdBxoe0IyCV/O8Ia4rA2Snaa6TwmQmmJuVpECh+D6eaE5NUG/aGAAY4TcILRBDT5cE3M3Ke
MTl1706PwtNF014smvKWSoXU3p7qECtv7ZLtCCJnE+gvnms15W1QbjjU0/3+AajNc7x8XwjxBO2Y
XLm6iOuto/NkagjZuIizj5vU2FC6hYGOCJDR/x3627XUJeH/WAXl8tPNgmkpRq5lwpDIymX9EC+0
pqgg0Q8sLQD9opxERFF0wyue4qE8Q4yabKtNl21KTTldOLaAkT1ll93yQm0E7wJZ+3fFG8ncL59l
YS50sIpkJCfQWwstgRbN6KLUU8fxGiUq8XPpEyiiiJYF5QhXcsmdrWArURcH65omG1IZvWaAYz+w
EeySa3w4Nazp13zA6esGGEsdLmRDIVGasxlQiN3jmQzKZ0Gxuxq/gQ+40qxzGoPPE9c8BZfjX7W1
crr4xuqSIaduKauTc2/lrk6QASXUfbpom38sjuQbgGus6+sNIjlX6Cf8gFgBUVwYlhnkLurz28O/
JKPm4OywCMjunOj3MqlvfI7icCGh5qRC+4G/g2MzOzs64CFBqNQqAQYcnw8we5zLzbKifIGGYJq8
DqyIS8Fgn7wXmaWLHlHb5aBZWztHcND3j3UM4qrdL2c0xB1bCAyemb3cVQu7WVj+JZ3WMZpBonGz
qL1X7QPg4ri77bWaYTqBrRLH7l59SJGYvpTdznMSgqAJjAgOnY1JZsgXGuBnMSQxdVM87M0m8U7w
k7/q4WXBkol1Jo8zd7PRPnR8EAm8WSPLIGnHo06qj5hfXx1PDWQ6yCcjxB0eWdsD2PCAKqt+3ZE3
SPWbIX7Q/K6x2xHXZAR80ReAtfsOF2c8C3HAel0x/xsdxP63j9emY6Tsrl7mAJKT0a4fTLSFTqnc
ZqL49KLViA/WtVVjuRhKVoGMAmxeOz0OEgpMbc+CiQhXN4Nb77u184wcvmL/e4GDyJvl4z7wyUNI
KKcQLnX32X5CMsgpKtmsChc8M1QCVhEhJBimsEltzmtws4ASW+E0oLS0+LWTYG7WwBm7uTxXW+QL
qIEkzb6zjMIcrR6Wu1GqkJEshqh5qgyoy3NhdE6wEH1GHkrkGHD+yF2tbv3ap5xHqPyUy4SdHWzb
obcDelWamjPsMe+XVtjjYsqkV4yh/Qu1LBXAL58/ACcRvdqIM0aQ2sI8J+NRZLKFfKftIfvI6qKJ
gHK2zSSp5fHk+1ZMZiMQv9PeFKXTwxxYOwDmA+Gt7qrTeLsZByZdbjSwriGSFKAuNKsqmzy9abWT
4ro8iQ5qjtATvQ3rrjkoQxCDYQBbIh4OWz1FEPbk0jaokf3wA6F1EyT8fSx6aChVdXJ/uSl7c+Se
Bd9zmiCsPKTRvE+6iU0jIOjXVrVjSoF6AbGs2HS4Cxf57nMYGB7GqqjHLNfw62o44n82eVgfSB3z
O2a8JYTXnELwTYNhckUs4PYJQpodxd1AoP5VJIVYJVXSsKSO/eXokVJnkUr8/i/8p10R68Y4CNkS
sr1eaI4SJ+b4uzuRSPkKFCJHrwv2E+GNHXUR9kzADUQ/dBmH0X7tSi7S6Lu3Erb84CmIXzYLrBPP
2lAx8YGBX3wRpa9EwJRDsH2lTTCuXndPWA1l8oMrsMfiYa8lLNw113++WQyGsg1CNmmQSQJoMiWi
ubp4z0RR4e37bSQzLkD+z59nT/93BRKMLa0OqscfRnJ67lFdZFO0djdm+jaW667sPWPvCKIwIhUB
B1q5BEDcKalHrhT1RsjPfpxhWBPZ3ngy+Ph/wMU96o2fBsE5pcaFomQ1za7ex+yMIiWkQZaz1nOf
BiU3r51HYOSC2+WvuSxcXt/N/iTAu67vKfwRUZzAlDI68gcNR+sl+H9xUFvYWBHGrc7tlaRoYANM
kMVzES9kphjgHJRUuE94wxUgkxIZhhdX4hFfXDK+5dzX5j6TnOn1rkuw1LK1Rb7hBAH2CQnNiTgw
yX6HwKw8FwcG1+A2Ur5YklsPZdpKubbEx7xDeAW4oHPX8OZRe7Cb5cZ5gEYG6kc47aSpug2m2f4l
mEaANYyWMb5gbY6o2fkzlcjlRVHhYeM9YTOTCeQ6Mv9ebJ91xNMiZOsYr0Ncmk5f38roKw5c+zGW
tundo1+uQIZHLMfNLGbw4mLvn+yx/GBSa6lw5ofmdCkLB5kBe7r9UVT2klA/imgxNO+AdUsWTe6c
4MB9Pg62VA04aWyT9QpqJQOkToq17VXGCAALgAV3yOhwCZPuKdlL2yIuhCQseRzXZZf8sgOeq0cb
SjLeW2+IuG3sSJ1qPqL7SPzg+NuXIg81TxrKydZYBpeWoNjdUZXJ+KOUrqeNbhHqzmKdsZMcgk44
/axSEt3+9KwK9R4UcOJpcYrX6zeLtvOPlaT/PmMjHThxtiPZNN8fHYfLk5kNsLHv7Ckmr9SLDjiv
bogOhuZ8h5Z6n0D0X+e2tP4viit4Fl3enJArp/4B4LRvkseo/1a0AYCVJcJQEEASVls5R3wA3+2S
Gl8Lg48Z4tjS0boepB+YV4wFZjTJks6Phon/PV9YjJiMeplke0/w4EKHPq4iOsMQ4OxosPPoVs1P
LxhIPJGCzPHjj4fu6NMZU9m5I5wkbctOyux20CwJ7Ywo3LeC2aV+OIAtHAA9NGiVrcL8jpYbybp6
B9eZR2EUqqVTyOZr7z23s8uyvYXTuBQMqiabJSiEYQnahgtGzsGbM+ZH1cNUP+BsQsajmt93kOAr
u15GlXmgQd/yWtFr6Bj1j0zjlbDMAd2CdOzIGIliLFj+80v6oM3ovip8Ju0qKnf5T69qaMAHTRE/
8dEDJbCwdBvqZiKpFxdsUeSKNLEXyB5Lp0Zs7/XV948BL3rkV0g0ETg6E7iA9zsJQjJMrSKG4OwP
308d7xOQn1BrId4MHW173eIHpQeD6sZSeu15UVeLcpKr4+uT3+6puQh4dd/sCsqzOPvu4Q1NUpjc
sEtNRXfCYHaqNLgDMUlCKcUeKDD/8E/moNPJrjtEYuJVHrdEOGHhbLtFPntUWpLCaANjYgPxhLJh
CM4DUTvmBxXhoSn31okmVbUIJayxidYPRqbSTGeqbgZI1ucP+dudX7iBjL+ozFMPRGXuGYqz2Xyl
wLrT0OjcATWUuvlqM2n8QFmg7dC1sqYx0MhxNo6PdLpSKTSwABjdWNAQImDXh0UKPUsRmoHnV3l+
9AFbvXBKo/hY+fk9MbTrGooySf1nB0uZJ88T7VT+K/WXHrMy2gUxszlaB881yPL5ikQ4tc5XV0Qs
nsm7LOJSvczSwm+xp6r/9KOfbrP/rd0clqHx813BEpJpXgR3AT1owEJCFA/0FSb1fTrL697YNrNw
5DAj2gnjruMcId2mkkpI7HYv6gOHne648cssKKXZXu3NoDqedGnSoqEOJoms76e8QrCuZsR6YH+F
5CXo5kpkf3zTsq8ugaD0We7LiliUCkczZBcEDCgPpiAIFhKlvi20tDf4HAqr72YF6ikDgMedfaQ8
VXg4ORn6VDpoJqDKPG6fK6pKn2mvMlqeGAZFQABSJE5CcEGz439dCgHqbj5USonKqx2qRwD1UWOP
Cb5rXIhBl8f2UWO9LhZMRO2NPghrIUkhG68qrpFotzlXj3zFK8+2TyLhpJLL813k+UkC9hACXRJT
9x6IxH6qZmYHM+JzGASHyRHmiEQa3ac0Wp6LQYCttF50RDjwK6vfGKQX/qw/4y2kvotW//XFu05X
delUvhmtMD1q+yPgJqU2ufH0vY3gDv81gAJojINunUQ604PnXedofRtrvl+3rPgWY8Ee5p8ZVKeD
R5VifbZFoaUCpiG2ooY9Fqg1Ls6S2KCwdEnT6MbPMbYXRVffD87MUtlVg68cWGSPOtnV8GX1dxNa
OaRUoTcHc0NWewZ/Ur5oeZg/wNH6qG5KDhlqzqFBZr3SNKu8Uti38PbVFYJsXKMf4ADeSS/6mf+I
3FxC3fQ2O3zdAhOmbI2ytTRB/+knAjIoKkZSCzDGlDd0yappdukKBC1niQiGl5hiP/VAHwxl3sSn
9pS3P/H6PWnHgSr31aCoDp+PcgkfSlcvumcwIW4iMpsc5NQA4weOW1t6NYtUc50+B8zHioXLtp5w
kZN6XzvCoR1uO+srBh3IU+nbV5enip1I+dqTnQWywc3h6nflFr6TQmODxtuq7CSftJE0MYlIol/9
xp79DH8NrGydPkbrft8LdxMCnhhwBJSHDbEe0Xzjf3dZ59JTgTLqbtR5dkr4OAiilXjgS7pEL64c
ye0nn/zsyvW9uVm5UP1a2OYjsc0cYAXEmUWNZqPkBgn+ZZr1v1y3neTeQdMOSaCTwYIsoLBGdBnc
+RVoarPaeGIInXQ6U2v93MNmOL824Cl55dmmM9QLbWNgdUa8SNDbQB3tkH7Fg4EA2RfBzq4THg3p
uGJeRpp0mVakUSKXKsgBdpzYeGbsnLBce0J/13Zrvro/y7cNcdqjWeFfYlqmrzorqD0f/wOWmjg3
99ICW9/1m5aHx5HEFI3KEhpuHf7yTCd9n8kN8A7+lM8CSlnVc2FSvjH+EoZZe5nDxRYtnjfDx0TC
v01QWbUQxIm2uicrlxFvTNMYPwPpvU5SQ+oLsI+JOsfsWOOqz2U1WECskwIJbpo4T+sMwotKxK5Z
83XEm4J6bR5LzeCWJFYGUMujViHIOa1aZWnZsCNyIsJlx6WdrPYiQUSVUONNZB16J2KylkZnge48
fIbGLtmu+NPu3/hL5JD5zlN28e+C+AaDgcfVl6l0MeToXWBCJ1SwmS5ENX9fR4vcPQrJFE1CnnPD
7++AvAZK6VEVrgUpkM0jJsN+xJ8TUFCp0ICu/3iHYaGYXmTW1ySW2mB9A37bPS/e8hcLJNr5vC5t
PLD0VpFRbNZgx2bBGYvadUWIr1V1d0hyCb4ZI0N/bvveCOmP2krGcQ5+FMRvRtRcpST+wCkiErIH
xueXkNg8H78xld6UtaHKNowksjg1V6OnQfQnxNGn82d5/m2hh1Ho7ZVI3xA3zJvyAjvPnfNAzD/s
LUBkJJxSWYVnWpisHMPEs///MaskHNTcdUc0cQYVDTVaOqBRPdKB2IYEXTztHfARDObz7aV6qEh6
txZD38iOkLL5odX4UDtX8Yxir+vEDg6+OjZ9d/iL8Q3UQWi3BbdVMM6Zes/UL+SiPv/1U0PUrvNW
9pY8wsjB8Kq8ocr1AZrEoWlN1Jnn1rcxVzmitY7Xb0QffSavhU97+rFlF//w2IAaFstVam/9TIcH
1b2E3+GTZYVSFzQGIfoFstMySxWTsfRqyQxcmjE6uxfoar7Vinp28TwiTP88buZ+6yZ3FxDzf5Np
5UgBy4A8xNJVwcLQ37xeJFk/mNDJ7evEetIYevECSOOD85VzFzcZrTIrOdX+OZVENa15CGj9BKPI
OfTY+8RCWFQ5nkpycp0LW8ZeenbsqVWv6h+buq0Og4eUlta2K0D9BJBJ/zly1tdPUux0xwf5Mk1u
9aUYDzMD49+bhfW4u6rsF7Fefn4qqwYYDB9GGc6VnmGLNMUu5QC9Gtj16c3dvjAJF3hCI/hTIk+/
wOQiRaDD7/hrsVjZdpTKD4knaUunSAqSWsiJC5Wg9um/rOxEufHTxra6Qvb0qTsTUa9/hjnrpcBT
RCx6Vke+0OY4nasXXPt27KJYhbgrBblnOBcKWTMW3iEvnw/MnQcZt+7NUB87OJKD1Fjr0M0Pat8Q
IaXkKdJzRREcp2J9wKeTi8/x73Fhuv9AQZxoshORcwsL1nBpIg92pUc77R+ADNGOhxR4WAAy69Vq
J0s8TiCDJZGSCF1OeiJZ/vJA2jyFVmDdzHvA+69kIggu3u9XWWTYYMUkFUqVB8NJTy157TNLayhS
myR0hv2af82CzqZt46cMaVTLk1ZDijsNfEty7AHJIscdah44FU6bvhjGkxNpT72NZtuE+gw6IeOj
77fBi3DXuxY+I9ddSnEMQwus0oYnDkqHgGzsBHsx5guo1E2YeJrsWsYLZHwTJ+7Kh5hrYk/1ZMDL
qw0maAMbytGxp3IOcZhQwwIVlLYI4sU+yPk1Un2CICcWtLs97vaWpR8sKSH6Vu+aU21XrgDbtCzq
7Ph9AP8kWoB4okF5tWBcoc7cJQvZlJ4tXQMkN94s+D9ysF7pzXXn6lk/K0D/trvNk5E+iH9nV3EN
DCWi4zjPQS8Jg3Ig/WUGenHcSJvVmrO/RTDQuYIjU5k+z0lS9ndFCLyP6Qw2OOEtQIxNTVHCmQZl
jI+Y2AkLhTq1nSzgD2N5BTf+q5nr4o6SprpnoCJNAvT7ltD1cX4q0fB5HdXFAWt5/PuTC0ZLXK/C
77aUmoHIog5wlXV5fUKPpbvYPZPbW/n++scJkIa0tYtg7D1ijZENvQVWWj1SxWtC6MeEUKV/cear
Mgd1Tguvk4PCq6G86NrFnZWefbAjrAGWHskrcZljLDrFDqg8juFGwGGtyPHiFuqEmkbMCfL4wxUE
JD7rms6UXznpfXYJGI43ybOxsdeDzM5Cb+xc8t10KgLVtG7W44HsKuezmuIY3wMHg9cacYy3BSaB
D0k4mKjVYT701qm2Zc3hmrZjiCZditYaJiGWJSoUkMAgUlB7eZrLgHANrM2W4o2MLrUxTimrDzk+
ExK9wCg0+aEc8BWhhFiRTcSk2AT0XdCQ86NFVOAPbortiFjMsR4fwEElvb/W2DHJCNvRIIgh/y56
3h9iKORksaa//B3qqVuVerK8LjyWWAaTRTKxBIkrEe5WK4AwlNG/HPxZbr8xSGm0QEeyaDesEiC2
MQ6ReFFI4Fm2qw5T1DWBbgrSdY6cb+Xd8GgQCBiiUYH9ufKmmOlCWd+FmJqBgPA2SO6TeRkPKxIZ
4A1Zg6pqPZYgvFcWbHDN/k2SewekS8wUy7615wU5MlotVjsxCV+LMpV3fOOR/pTqR/r5GLJ9wwJd
gD8Pi9wHyuX8boUEYzACzG/Jsfby2t+erTpYNayFne+dWVv1Zdo+MCZyU5JzSEvKFrRs9Ku64u+D
sLaTTSjnGUYWoBP2sTSoP35iwpg8b0W7c/HyMunjPc80IDbSqcF83cSu7xOFaYx755mw4s4ZRua5
vuHrhHG6MfyQTFPemJHx5frIa2kOmGsJr0mWU2FJdoaMG3K5nA4FUs6D1rbvtvxT4iy5XwADqTuk
D6GosrXjSOjRf4TshFdXnNq6oPFwZsSWsxGYSnzVCZH6BYTMONTqpQzcrvZR4RjlO+QlR6syaNBg
8uc4w8BBdL4FUOzM8O4TemtRGnefU6Mwtfs4NFC+NrA38Xr4VpS4RRAqS5WK3hBT8yqkYz3g7UQQ
y1GMU8eTPhKnHGhjBa2Hn3/ViNg8ck9k2tBUw8Z1IAnJIi5ZycuziuZ4PdZHQjsMV68uJjSfW2iF
e7Vb5nSxwBothd7m7TlKsL4878x+nnzHvxiGrakGmmkrBaGP/OUq7qFxKlXY1AKu0vSLWlhgesAl
R8E+P3HNsg77Bgm7QaSzOp8iwaWR3pl5379cCWg0z9Poxykdh0OB+cXoJZU3qht7EejVhLzGBLJx
Djm+rONmrkOEvs9wA8mVgK1YyiyE38CZsoVCIJlqMjHWBKuCwVq8a1nW4O2sYrzFTouT/ruMRuv6
lj7xBZnRxpADJs/nuolLRvQU7XerjkvMuEM1c134YTGQ0hodjieqRNqTpBrMGXJKL0S27yiUz7jW
dUYpR9qto3E8NIVd3noLDcQhzKrHWtz+I+dPBuX9V02p5hzOFzoqX7hhe9F0+Tyym+Ilg/IRKJxl
V+ft9ElBQa194Hf4AHyolmW7vqcGNKJJ/XJOsBClWvZMI/kGnQxJ/swohpbfso00DH2kQwhVyjCa
GFrYXcets2yrGLNQMMycvlXdnJAd9ZI59DfpG6RQkBAVrZNgseXCzHLqzIdvqsji/2nJy/M4SqjZ
B0tXUJFkc8DhJEfvmGbPRyKIfJTD2waCihEltKAuzRyXC1UoPsrPDABkOUmCpqHfk4CiwVgVWiF+
z+5mCE9MB8nNKc2J9R+CUpnsVh+ZxTMrL+wCE/KqgUxKUR/ki7pLjhOTL2GHYOBtCe8VVaeCAXL8
BrT5AIN3wTR0Popn1TqW0RAtBTey3j7tDbP869QMagiAn9IVQV4daMIlrpvwGHfKB6z3KDegiS8u
dTs9z/qMBMErKuP/HUd4LXnDn1QuwVUVCc+BIAuxN0aZs7G4DzGhPr6ye0GkIWoDwsSUSv8Nh0hS
rzaLDR6Kn7tpji1iEqG6I0jQ+KNVxJMx/GKgGeRuAX3KqzF4ydcq3G20D8aubHwybyX1g+hYOSAA
a4OTf5+MSJjrwfEjBcJd/gnvvR1a/XQeM4+C7LinFlYukw2cJwuCmVKXkFsBq/M0plf0Fx0p+p2n
t61jSiih7kp0eSd6o/cuI0O8dHAka7QvUDsT4si6JhoalLJ4A/Bz5xDz5ofeRR2l2OOFzMGnpxxe
BvKLwFgAaAn4g2cyO4iDgH11MMHJG4M0qSq2Hc0kxE1yCJ9OGBp4kxLqWXQT/X4jNYQxe+YhoaSp
Lv2DwhwhCIAk3OerGYJVgSSt1c5z/C6QknqW1SHfewVg225YF3jiMv0BpGntujxu8LW3StFo3zHM
y+7Tq5g/p5AVCuwuECNeB3kEQVWVgGXTPJwLMHz5aeQ5yu0N3UWWpIAognQr+KfclvoPU5bcJWH3
aE7vdkYfMxSmh22H4gaXtxCuykri4CcbEi/FmVGM8eKH2PLu3AnrlGuoNPBKLocBjCx+yJyc6gm9
Yv4b4f6OYEbOGhFHwPmf4YgZX+Hg2rY5X0es6mU0MfSuKjVfYQp2Zc1rlyF5yy1UkcK3unDq2JLR
T6aeGx+72i7fiqzZ/5xFCuNQ1sbBvvRbTq8KQt1XXrq8/sszVdZSA/wiG2PVEUnk7oLMPNMmWxxD
GjkMIeDV/acjy1gx1QqsRcZRzZ8aMOgiFEbyaQ+cOOHq2omblUczJ07r+IB6V3tgqTINHZbD7oVW
MVACIOgrcL3DVH7jttdmCoD3+T29OV4fEP4k8VZSotz5FcklqUBV940D8whdYiQTo5M3AMVxJeW+
REPwFG2VbelkTOU7oQzLgkxjnQBO5YHutmri+x3UnYLzWERjprUClU/UKr+eIjlCXSi209EkV+eR
Qeg7aFqVrCUAH1xQv+vgQ/MsCZaBnlF9R8bUns7kDR/ur2U4cEwm1zXyDzUiPhbpH+5Gm0oykHhd
DenlrTxLOUFU9K+/CuZpiLy4a5JwrgKQgzhyR94DJ8qSYYAGyAF0QUyiuhZdNbeGlxovoGXDwZK3
HsPDB46tr/Q7axWJqUO8gWO+Jj8mwIsB9pr7LT2Hab1bRRzPB5ARKnBAbXwkCIIgdfsv6mPsELGj
hJ3QWE71BpUFrMf2wYKOF859bW2DhUz7tx5GVbWjLJlyvlf3mixteawdTnqkQ3+RTLnV7/sjusqr
1sw0hmP+rJDaLuY1qHtLsZofuuIqtX4fDdWY/yxjIMKgWBz7ckUUNaAHkKbhEK9gqd891KJKrBQp
KXq+tnxuFYgEQMqXNZe/wtmUF3eadmEF5ze04/G3djyXvD2pf5h7TjWzLchsSCo28uuUJSc6m7dn
4E+Qp6kcNtPWCT8T4ubkDJX+Mt/oCNrn1RZa6mb87isVw8qC+gJBSga427h69f6+gqjvmnmQqoZP
vm7w+XLrzDXo2Dh6lOa36ksMFN0Kzo6rh9YGd2afpQk4JeqF8r0qbgftOVMqh1vqs6pKdsJds77H
xdTGE/xSHBPGtH6pyevk3fwkVie/80qjXtQZs+qIBcDZ7s10BMtS/mkpa19zix/VoPIxUztRaP5r
yPjyhlFt4Ujsk26WllPrAK8zVzWqCbPWluVnkSIZFmSAzF6f+krvK1lJIaegVKFvBeXdvgnwkeId
X2WQv425ZzyJ6O4ZyAB0STrdqmYM5594xbbmR98cifPEfv4ejKDZYbC1OHTflOWrHM43SdKKtZJo
g9z3NjLYqoC19CtVWDJUBMQP8bgt0Deh/BNGmRTLp04YvbXnLq/u9x7Qr0hrMRkdYGcN8Eli3lni
C33miR4cYwhUYgGtSS/9d3g+R3hgx6HuT0wLqsorq42Z/HO4VLiQ+mUKoo1yigcXMyUwqjXHiXCY
vdM6iZH/Aqd4/+5b+QD7ouxgeH8GRtWJ/Aps5FUw2ZNliscNV5zWSoaT2sGd5a5jK8Km0jRxJvTc
Jjc77t4PlhWjzBX2hx8CFmzjoC4yqonUrve0EVocfUziUpTJlhTvbDKN874SsOIi2i+iIvjC/I32
gr+sRH4P4GEjdol9y/x0Woyr/mol88Iak4kEQ3wdfA/nEXxG/Z5ZFliXVgQlC0QAUpoIhM127cTI
vch9LptQ4ZGdNeSLotMHcY2p0uaVciPJv49x79W1zqTqopmrLDZjRmBLxTiAwCqKHtruG2/t3b2C
jz/6KKp0fXKckcdLZICnRlvmGxSvQCMDWw1mRnyuLFhf5QaTfoejvt6GOf5ZXAE3VaUDNphFgCEJ
uX+UzbDj844OOvULrW+14bHcpECjVKQ09VwlOlyw7WtChJa9nSxpLlZbh5waY0n+U0z9Pd2NbP5L
Xmhf2MGSdNMsJ/lAf5Yf6hIng7he0+lk7PKPx3kiNmkKqlS2CzqU2WUL2fgB5RKyUSAL8gQ6eNrc
8f3naaCqhYUFMeLfFB+xo25eZ7VqoFCxJZlD2cR3GxdvuOzM/YSKL9jY2riij2m0B90yi0+gtAx4
IqeZUII1wa0lMgnGaqek8SDdWd4aWcmWnznHilIjcKHUwD5Sj8XIbgvdT1DexHQiXwEvkI5bQfvb
KLtZ3GNVkci7y+PFyUpiLBAf6UcdxCHtRrqbvlr5Eq1MXUNbrTJqVyTmjVjNgAXbqRr+aheAeWvL
5/vl9nX3FWD7bbxB10pxWbnDaPBxl864XTqZLtEKowAKHQf4SWDlQlq2RIYq7auOAHhL33eIR1li
hA3KsLzc8RYCe0pYrmGMBd1q2MHNyT4HcZNlA8tyMFQ7/P3AkUNwPhFCGCpY+RVy+qG0htn0xYnl
sQCjvJjHQMUs03teYhTnupnzCJEe9tRssxVdMLHWjb1Sw4WWpcCPZiq17rnKaUovS2pPRqnAV8ST
QuyH582q8LXvViVM436Z4fZbRQ7EogF2m+BTkVuUImBo9raSD6WQtck/hxqsjQ2sk5j7EQvENhW2
5ELH8+Dxlz1ftUxKhaQAQgQkwbhyMtOJbndYvYhCCZrWaXqGlVt/OAqRQGHkAip9vthKtlCwnzdp
mDnfOaKWwu1LuWpwpUqwF/VqtvugpCsrj567Jr4ECaRWNXnuvS/hXYCIQTzf66K94EXo8T8VDSNK
4YVCG/VnbAaCilf33089cJFYlvaQID6ZgOpZYgO7lFUMtdoRZVfI8+7d8iDXRQRv0IZpPnBUm/wv
90QaDA0e+4KqRCqBd2YTfJikyKYHiEaMDuhUCYg64oEZlGDv1cKGdgCsvhkrir9Hwc+UW+TxrNHb
Am9uFgumIIapP/WQJIHLInXXGM7x+wXKSDSKfq6DbzINaV2Xjo4EDuAB0s/yQKW5nCBgZaN4MAxx
txAEIoaijBWhXb13gAnomjAMrk6i//g4ytEhrDXebVb46Nz3dK7JVVEedvVYUnlgI0UpbNV2av53
N3K4UbeyGFhnjfbx+1oVlUdD7C36+ha/S8rQeCBXTs92Ml2b0f/uLlryPAYfqEOzVxGcKPfpobka
5zfuhuUiqMOHO177L9ZqeWn3KcZQpmFv2Jetc084z6ZnXhY7gjtepLJDvoHWewAlbkXGVSh+3+4F
qdej+CZSNN3XmpWhDEnsthYL/iARgB4HK/X3L5Kt/lHbQLy24xP3As934cs7XciN8s2Ac5daG44W
Kiwruv7yXqA9mg1ukpeKTw6M75NWnvTqWALLDcKBUrhAzjiydoyFL/Zzg2FdE9tSmXSNW95vtv/V
1UVXFDZ/i84VYlCUcnkU2+R1H44BcYu7C7CbD+d3rmheBFjsAA+7dwnR9HFJ0yXJdYJqaepwfcPb
hLOZShX/EgouWadJfxbU83vC6LoAZGvlGXLHKMgBOlNNf41VitAxj3SnuTF7Xll0rN4xNBWpG/8+
ldUaCZitlLqfQQO6tZ633wqS7aZ6JTNebkEtySnUR3CTpYFTimDmI65IuKTthm/h+8w4Q43E18W7
VmOrRfOBQCAuEVp0vTsaiI7aQVEGhhYN2NKO5gR1L6NSU+4mqnM3yEdo/kJqFQkogdwoDGCkuk6p
GWoxva5ESPE6wZJoXLdLUIE4W6eUVHK52V07lndk8k9b4ogjBZcxCgt+MKtkmprA4p0iMvC4Bzbb
FmHqIg0XUbtEfwV6Qa8qdnEpycXWQA2DPgOdY+MSL1dbbHIflJKqN1ojLsQf+aimskgjE6TIzN14
F7WcC1PG9LXmlXRQZvGKkW6YHY9GC0c349L7f5c73BGd2TLZTX9SO/tfWz3loED35FrHXk4BuMnD
bJSnrcF9dRHdj8W8qkSnkiZqvJubf670/X+/nzoqBhY8yePk7Yxl2Ph7ROBuQTBNym/id5waisNY
mO2n4sSo/l5UlLi3VNmco+wOaAFeVDeAiNzjDBrtX+MVsexLCsV0qtyxrJQqohw3juz90bkg2sYi
7UT8FG+jz0Au6wl9rzNAcgrV8jPVFx5Y3Nr1i+DV6fc1/qsI79ohkhH63Yi7tQuGzUhLaqvmkOTr
0Nf8505syhkL59dLy3XGkwjMkGzoV6HIP6RM2VnpASXNPyUWw1ALqVnX4E7hXVHPgpRj1ttTvWUE
WlKORLfkdfaJQ6vJMdcmqF72QVOsVN4CVGQWdxEX3TJd6XpV9NG1bC8wvUJ8uK5mtN7j/OYaAf7m
UMaI6hrHpy+wjhpAxKnT7dyB67XFEWHwh0IbCyr9pDEmSjGH13aqIg62yHlffdRYtV6xARwUaNDs
z6Mw+YQQv3h7x7U+83Ck7IC1v7Kg8EzEw0x7JQT0fAtdoNA/2zbh/4gTG8/Zq9D3VzBbAEfTY9F8
uQPnmS8tSNykLN7rAwbBVFabLIajA94Xh1y0j3snVfjSN3QGGmzBkJfxyrQBgABr8kLI9loReCD9
8E+4hDQeuW/AY6UiHKvvgP4s62vePrGiyIidV8dNDHwVw4ijByiRyCmzFnoSP+jm4TA9bchAjYLq
Wvuy0TVJ9EYT9KNBkEm+HTDNiSUUb6yQazURrw4O4r3aRJ1Tn41Ocqd8ijP52FCfAUY2FIXTi2ar
shL7bZgcTUxBnvyyhHs2Uuv7ZGebim3H/1e0/GLV3M+lRuURyssC6xvt+8uL+HtAzeFIAyJByQGX
dSudTj0w7k1ba3r+GKrxvkNMXZypIaHsVaWdNrrq4MhFKJkNDkdMLcXHG7LpgXFov1eoxK4dsPAK
wrddokVf2LOY7cZuxOc7it494p0g7M1XJCeVkgbBj/GcnKYxJRS6NjNZ8FJUitCOMg3v1uaaIZb8
LO9CoDjn7hszZJliWOvBLWmTPXk9aQ7/2V731xly7cfLM+so0TeyLe8tpmmaDT4iV6RBIGpiTDmD
iQPfRzEhOBCfbhm/rdjRNV0QYflo68U2eaRL6xM21n6QbEwHB/aoC8w5IU5xoi+zw4M6JArUBVOB
4wiZNttSAcy16hfr3GOcVvibrq5gfM8GQPUX+/BrAMxjFCNnLLMzOcMToU7rPPq2+WOiW9l5KlpX
+FQPXN5077NBgAy3nTqQsI40K6w+kp6T5yVBsb8swNcbwf63cIzWtFs3UfAyCsxfvcbGwxfr6PFu
MsrFvyzg1/uuoIw3RNaCNXbqT7lJMVsbZYE5fI/Q6w/p4oq1NNrUpVWXTNlYwD+hXlezEmhO8qpS
fGIcHKEVTIs1LeY7aoloduzT+W+Obbn4RVjDM6W1fgGLTVjlsuFtxbiaJKb6/My86gIFNG7pY+S6
XqaontUs5D+tWZNSrluLy+Rtkfz3L0knO6wZfRYprsTzQ3hPI5p3mJJkYwhwXhcMH+TQTYcutFAk
ROIDcLxg5NvZ6F2SPYZ8ZwL/dvdPFN+CHrfKH+9Sr284lBIDiA5ptREMJLdZTMo8wBd04r+IEGvZ
8Z3bidsK7XEeLGmWL72dX81ZCWyLdPheL3KFRxhjpL23birhQdU8QI28k4hgWSUnBd9JfHsTRZZG
/zOgQCmBijYutOu0c/II5TgkUJX3XuN0yC4BnWHy22qwqej3noYFTqNIgrwAU7yHZaG46TF8G2Lj
TVsdslNwWdsP+CtqDtcSRnHjRj6si3BVvnbeH7Gjj9NYlNUq9BhcZrVeYQ1QE4z47keQIwsap8Xl
8oww6Wk4DgO62XWNUOH8YM2JB7uysCFbNxih8XCSBOGMuXkM8SSoKX2Wva90Jx7FplRS/IeVcWx4
fZBUwU9wj6BSyXjOv83pz+k4wcN4SuvRoAb1qU7OBNKpRYQQe6D0EsYb82MuUJ885VkUJNNUb4HJ
JzMQ1yIEPSDbpn+ywyt0p+KSFpBxK0ZjJz0mL3+rp+xYdPQNEt56irF/lFcyrs6SakUEb3uspTxz
JcKnTlrc5ztoSDcvx4SBvXhgschUw6YMsrIvgVg3Ji+LsEPEh11tY/DBnnxwpI0Rgt+p+hC9Hs/w
5bKIn4jYuS8pLMW9hwAuiSA1pGdDrCiIP9ft6CG9A3QtfRAaDJW0i6ARTuxn86Em1m1ij8mo7VIa
xu5ACPuw1YNAFRJ0JMBPTFaQ+pLtkxYI49n1Rs0e9Y+YspHiNR7YScqZk9R7W/RBUABDJCCegCB0
Ah6bZOVlh05obXOIP4dOtdG6LnKhMgQmNxczpaXinSUV/8ZfXFC49aXAE9Lql9IO5U7npbXq8AvO
JVtGB3kJc6cs1u6h1vMBypnTHyDDDQQMOe/6A09u9jQJAGM6kMWQNoe5/vL/hViN2vvZ0FypmQdw
/8iXhtaYH+BdlPHOMJnGGRq5V8ing7vqrZ+LajYGs0RR4W21oB2VxP+ShKyx522suhFf1q4SAI5f
ercOAGCFYOBAhHf0/BNZiYdTChlV1TBQAhQzO/D50KdaMxpHus4UdPXYvrTL5SeNgCuDZJ4I+wL3
LuAq7xdSjOCGoSARn1KK2rEH5ncK1hzTvKzD0PBcv5lmrTz3R1AVX0dOSXm/7H2h8RxTtPJd/gjf
/Pd2OxKi0s/ZENRmHk6PsTMTYVIjDiCixOyf9vfMKquIfD53GjPCmoi4lwB3dfLMRIQ7JeJ/gFD7
fCgAAqygd7Fg+02Ga9OvQj0PDe/fUdY/svyYd+6nAjRTQHTSj7uapVARGdK9YHOnEeND4AsZ4AYv
sGDfbL1GKWxrXfre3Dq6a3sL7crFT10YPx2q1LWoa6TMc/f6OR7m8Tbhy//E9Os3OoenSJ7Y3Na5
zEWGxZ65AYlPm9ehI25XtXYpft1mYMdWTVDcavGFGnXrPohyRyy9GhSUqg+b7wvKUI0td6WS8Du7
ZPWEeYeZcS2sLpcI1uwxar6Z7ymjS1VEv3e5UJ73j/QxLZr3nBtCipkNtGrz9mn945wzRyzjhSph
SmQv68rrjWhDc855CMQreVQIHJ11TUQuAoalUHre3Mj9Tl05eYP0OcO9/6SsD9SgY64xA2er5tne
P7EFNZ+/JuX7Qj40A6N225w+Yi3TAmn7J+HkAroxS17wdKARRDkNiGjNTetfb8eU2SsDqerF7uFu
SW/zFMw2N1hkGj+a/62vmApJvuP/DSSa1fVv4TzwNpZ+vuYc7GJIrCXHxt9mwwxCmiM7dt9NylBx
utBQy0aQpRgcY8OBI0VEq9Y2XtgZ/K4PZDs8PVlkFOSlqHtsKYCxR/8GzpqvmmF7gA7yUhbWH0n2
a2WTilNpgN/nfN81LgcukyJA/QdJcGtl7OKIqxntZqTFxKtJtV0yz6uvR5R2Z3GAwzXtgSPnMEmF
Bz3pOBVUe4cYnwYT1TuodlGUNSyyLdGuLO/tRL4dvkuDXV/+dD7XQfatIId1ck8DhSO3wqJm8HFO
qt0fe8PSkuU0uQeBZ/JGorjdAp69SU0Y4vEVW6EJnQijIc3CMFKI/8xogh82JUzcWhlU4Z9M0DXL
YR4eBggYOc5fiQPIoborDxt1MMMFxTBeH5zWIXhSfLSIpygozkZjJuGx3eEz1ZUqcRdHvtx0Yv8E
3KD6qkC8prJyYNyaVF3r3T85256N7LwW9hWe5/ddKEdCRj08Ep5Ql4x9qcZ+YHIc+nKn5ILaVL1p
zeQmmjJ+43OqXXf9ZXLOXKy8Qyea8p0Mp6TD+h5cfav82HVOV4bQ0G0sQ1K5YeXe8VIDWg4pFJeM
bT8/RCaSXtamxJCcJ9EXoUfYHzP+MZLPlQn7VzGAfQ578GL1tJMW3Vu9QhJyc7zAaqZxN4LdKwT7
CuVoxO94x95Ok1oEoNBIR7ze7YfafXAnrBMzPpau0qvT6a2q2JzngadSzrggu8wzgfeyy1xw3GWZ
nT5cEAZlfCjFi9hB43T+fvLrMoOSh29OucAhqqc3FmdNKF98soO4maoNxP6rIXvogGADlXDNyQwU
62Ll22egzMmYbLGBvKmkpmHAeyBhuAXBkbXQT4auZdq9RFqAzeKmZ6u3/XBpOHAkkAhxDuc6mYiN
HsYzAWVRMMGN2iA2F77bfVBclf+xRjVrOOCqGUgn1NpiQUg9p3Fsp65vzBc7ImWBRYl98SHYtjuX
tTP9ncv/hU7OoFLkO1HgkHFJKwB6hgFjQQkAZs5kfeXA7G+5JrIafLgYDUTf/EyVvhgAFc5VIdZL
5nFew+/+n18ZwQm0SiQ0I0JhHluAu02QEttFDPTLudPBaql5OjEUNFzXYt915oHjzOwaMKFDlm3v
s0b7csjAPQV4BSbLYsiCX1yn0vGZSk+iNObAVHBcul+a/fCYGLldra8WlTmhOCxZ+pyXT49ckDMN
WRUTFZJFpSt2+XxlZp9hqw7vBskC1jwxmPS7QPi67MdugiKt5mQvikCvViD9LQ3hN4sLubc5cn4h
gqCaMVGdexRLZmMHK4CiZqWng+G1lIl1iwy5mFkZphM0Ydsy3gr328JjZUosvCE1+4ivMXtQG5l/
VkcPbs2om5AFUJCFx6/aXIGaUtbn0Maoxw1d7txXOThbMjKMRiCFQaPLJIcFkdhX3Eh9KEGHO885
a2hUj3kWTq9/qzaiSv00r3FJ600Fl7Q7er6oG0PygpK57w77EwOCu+4+XDC+nZ7TsA9naB7SGoV5
xkj4w1jWD0BilMwo7asTiB5aHUziMiaicxLODbJ4ejvDJQH8LKOpdEZ02zrc0cZKe9RhOYMueOB7
uN+gmG+p73mLQtAtjXseZ4RrhAhJrCBpszo7sA7w+/TlzgTfkHbE/jxfHicHIyQwAnYrXkVKIjYJ
I/Nod7KNF6iQm9gM7fwkpbAKr5GwxJisXr9hawDkRiIjNn9ByYKKTMn/EhkNi8096YIASqNqHoWI
a0Xfj7FrbuCqnjkSf+Vc2TvEPXTtoiPsSAc+h82G2/m2WxIe9KqK/wF/8ege3HKIdMiwRM76dJH5
wZjakYceSqTEkyD3aiAHxn4692lFKUyiqRKz5pvZeBvgIlyxvmsO1/JWlG7Jsk2V/Un9bGCMXU6X
Pe++F3J15gAmSYFnak2HFi0xS8Cgsm4UbC7kP14Gcuobol85svwHAuUPM9gKy3WWUcNg2ks5iJlt
HPmY7EMzURHq+swHyPKsT18Nro9o0toCh2e5P+KxhXgvDFrHuloRy/mbX/XKcRFTNGzbMCXeXLuB
GDKzZMU0TewJSiL1e+OgTZ6q04Dtt97Nu/oj4dX5YasBKMqkwnVqvq3M2GUoXCSyOqJkqxI1qdCf
X9DqO06F3D0sGHtUtc/X3xlNwcgKnnL8jdPM67xDzDsywd+w3YnOvhB3XHwZddUOa1vbsTiuFG7k
P7csJmTVd3f23wXV7kFIuI0vJ9F24qga6qxWrSEd8zKFfcOtCfZa1tcaf6TrFXmCYUhAc27W0b1j
/C9t8kWaapC4oc/76TPug1YyembYGys4OC8LrcgYHvEgjINxVxbbftdLEGuk8OKwxO6K/AQS+RAr
QdPOBezWDsEYBZ+e++NoERcNvGlkJy1QdSvOLP0qwoWOxN2QaZ5/iHPZ7IQH+7fjlWAII092uoOY
sgf1GGyW/yma5LJY9tMQPY3X/E0dvC+n4F20xg8Hr6PhHUdNrBrQnZvEHCx+Hr0PEyB5CQSO1e0q
P8Wutom8QDeplw6XoTrdjlP4Lh1dCpLttAd142qD/ZJGCZpa0sq4iNWYtpsaSQ+MidlhDt5pfJ/O
nSOvJwiuRC1KIhg9tL2X1DniXCtBCd37g0zjCse0J2Ugi9dktGLUj98laYKGYpocl5h2VYkiWsMK
kqSaV9QHEdHLJy9hIGDuaV7raz7kdZygr/V5NVzvpCVGI3PJc9cu22jd6Mcvj6HXUL9k0ZAQvmtc
fLfiGaY8+ORrzhgG2fR8fxU6IXUhElmD89qistNKZdjdhq93n0c6xs7HSPm9u+oByecde9OEZoAh
m4Be3jlWVpoZAxG4O77eMyJVEKD8yhoyPcdIsd9WokMKVrWdt0E81QDYwtbZdr0sLNr58EbIHRSl
zZhrhA/GyIJja989ptE2YCFStaJn1Vbvl0FmuJYWaCKWjmefcqrfVs6AjHL/mW8wjDUzFw/fbCaa
7UxBJxCQeeRTSxq6Vq8etYEm3nExDug9acmMTvsx3y/ilVcUu1SriC1VbM/Z1Cqi2izZx22cPw+O
gi6QIlCJ1cBTyT2pp3QaeIdk1ZZhhwawIiRe2aN2vWFdloZBqKewWetDw6UypGTcb36EuWRs2EmP
v63kq52JZ7VSSTwg7Dk9Tr4JQdjIBduNoiD1j1Dwu+PedHIfbMyzeGWAYWF15qAHnzXcwPmQADhV
rX0Zr1wX5zwC7uHH3VukhbAzHLNylYkQoH2T6NHHjz6iBDAJGlr36KMLSbTzntERy2mDYJWHEDYf
PuP92P3iA8folsUyCQ0FwKenOn+luxNYlh7DFQo6bePT5ZX+oqUXa+HcMFyL8IhWfPC336nqMk26
qYREfCHI/COwK1+x3M1ivBi/rCaWzd+Sw2ZUG6Bw+uvo43a7l2k2lB6LPew0kMbe8mnt2mvZmyPk
gFtKyDzQoK9ly0ADP2lwsKJnoZaHaJI4tQbM8JfEH3CkUADC9p+ec+Ck9efsJdGbggQ1xXGikMRu
9q0X/K26knsHndgg7monkk81Xkiud7vptJ51u2Q4t0YwtjNSNTI7LcJuZ11cLfUI+OtLc+VEqjuO
p9VoPvcv7vd4h6lHMhrH83uhLoplBw6xxL9l34w9d0Ncqdp7AmOOu44Gs3qgM7hg38cGCQKDdGzg
3ZF35m6+29KCcVnhpFv42BGDxeH4fdRRUVQN2OlceC5FJZxOdCM6aJ9PGY3IeJ4cRsKMsnmwZIlq
6fYPG6QEvwkDdKQJDGDokTI1wjqZU0tTYloQdpd2raewAqvJYA+7H2UviVElAG2ouPicT/1T1Lno
wa/ugOlFmvHX6TCOHqVoI3Zuo/fN9mewdsgLyeifWU8V3JqND7AEbCeKXMhq6Btc494hV+KoqIhu
7maEISaGmR5bvSJLII6KbHPx//xCOoXoFpT07FI0Ae9CjilCefGfoUHvyafSMibU2b/8H21zSsZ1
eUFy46ReyILHuk9sqDTKC66yOCtPPjEd91RSP3ff3/bNEFpcU841TGFbuMyKJyHKCppGHCdmkKex
xbwymBwgoIqz80TEW+R074TdLGrVbFHnKjJ/yKtHhNST4+eA2s0tIUn5Kj6TP6UguQmAhXX95Rii
kh41TD6l1f7UmNt0ur9T3VH6oDetm/8ztvzMAg+KPkSsECzdrC/j4+ejlEAwWWRVKp/oujsszLwO
iV5IBYxY9aNTCbmeb0MO3kF4RoGIK80A5mg7vdxDgrybO+6HBb2+OUQOfh3QNdHEf307wmLds9CJ
aEiD9UrZ2ZxIa/4UcVkPu4SxQgU2rnH7iewe+YFiD6kFzdmP2qVtWZUcoKeUVsXgfwaddaLfhcZt
txvPkVstvhwITsR3+rMTF8ZEc9wc9WMph6LKUJnKOAEd6urgj0AytO2uEa2SqYsUwuXVpyt2nG2v
ewc2+N6kTel48rs8RgWc7KhfHiI3N6vG+LMkBerUU44CuTb7gCLk5IxYL8Ij7yiNjhy1m6uApgbc
Fg2UhhV3Gd9Ib6JO1DQSChrGyT2CRu3ewPCOw/yWOPor7fz5PP6l84yYrY9R9Wm+6n4rpZavHBc1
3+PP8vV2+AW1H85rP/QX0pvpsJJMqDskqzAJwUDE0gZPL1MbN2Ah6xnT8/oSE8GIgYeXtTTt1eXp
cbqTis44XYYmAeVenN95spho0H5Ncz/qGI98D9MmNve6GS0bkl+2WVj8UrV+4vT1twPMraRwG5EG
LrAAlVD57XX+H5kzYDTcvNPXVftYSSDzhHkrK0aHOsEPmJ9/9Tn6ylj7pw7DAAjpyz76r5YEJPoI
LF6kOd3DaKtUKktxP1Fg6t9ORIiMHsVVFvbXGcVjIZGNAQ+MNsra/jbNflQ40dOH/q0mb9ZlLGsc
7KUMqQS3eUI+h/pOi/iNK1RpIhdKmiqStUm5RRTls27vWU+lAuVjPLasqfA2Jg47Qibm+TdoSfVo
HL74guls88IbCvJSYmxpm/N5LHqKAn8BUTET7lWlJvLwV+sox4KrKLpQ7RBdbhLduOe5B4Wyh82T
x9VYv7ZB2zE/h6XvErcyyLsHh6uqE5NTMVqOK/hUYoDhRW0CshwQ9jAPLY6sG2NXS6KvTjFzu932
SWdVgBIiRoKyn8ZjJHKe1BI9tv92mdiTp3sgbWAqEybN39ewjJsjLkZvI74b5KRfV0JKgVlbT9a9
l9TUZfi67hRVgi/hg5V0FkDTUGFj7I/sAls+6rfVr2SlMGF02j54eaYjTBRZp1DCsCe4V5yarGT6
VRo+q2uxKo8O7TD0XNbAkU0DbxI1rLPA2ZWYtzB/0BFGJOwVc+UYp+cWPE3ByN4GUVcEcSXe1610
PW0pZOakQt4wPlh1CougnQqw2GZXGu2OCUZMVaDSOF/AUNVVAQ2tqGPBQgbE8YyfNmlSrJBpqWov
GzBRopKCml791X4FBE20XlzEGjRC28xGN9qwTxHXHCpnYRpHjQzRAU9OrV9DkW6JSJqBMJFVXYFx
ygvEcSJOt1GljjxGWEMSMd2lkED7jOqzy5VmVMUZC6GicMFm0lWCwspoEhdSAowMIWeoeI34upT5
7aKRhQn/lVrh76cyhzJu88zyCfVIFqoGR9J3KJ3ds0VBW4BBeCEDb2kPkWFSZK2ErJ3DABnYwRwa
nscgUqMtR10YsWYmzKLTjP+2IYQJdCBw1YjtC6AML1NXEAcqFh6cM/oVh32+fk75vrVwGJG+td8M
RyqKa85ejbsE9H7+P+Yc5+UaHYpJ8uSy/jFzoFQMRrTM333XeGdbDW/qqbKddP7uobUVpJ4XqNVn
DhlFRzjRHbP5Ctv8lTL4FdnyQBpHALXPVGTvl3gtyImxTmALPbxGcahiB0gQCVKXwKimqAGO6fDj
tJBywqsuG+5GOHsegoOfOujmCyFcpEFJUWXMZmKw1ihv/5fxxNryCSwZrywivxfpY9iySsIIdyqe
uoF5ywVFbn6stZmXW3xzb1YqUrXkkgqDmHxJtKZFK2sg1Y3HQWOMMNG8eXjaUKlF2Ztnsq+j34mz
mcx8ZV+JWcsPOnOPZrLu73qgVe3JCYe0gDNLVOxz3lzYQIHjpbbFAriR+0Zh3F266itsTiM8oFQF
ZwiUBcrQV1vnYkmGSfatZU43lVLYs7gcpXQA2VFGeMT7MoYVRxOH4vvmmasBhcTPYxA/PPLA3AOY
eZXT77JAYavl4km5AVL+TWHkzoWCIit1kz6Y1iIzOXJNGOY29iinIQfAqFzWuJGc2wTUCXn+WioS
jVkI8sylFsWnVsCrESZC0je8r4MtzIjJWg5I0erE3sp3D1qKtVifgnC/FNuoU4JjKqxg9PEb+2v4
mf74MAW5p9pLwayMBLrD/DKaLt8lj88RqFnaaJD3MeaKlaZTtA4qv9s7fkQMt3g3K2becPeZds54
2nGBp6lxe6h2wq4KMJflLo46GWvtMAnN7pX+Q/mPbBMY7W5EFbj3SWZ5x/OtJFysgb8rqAAy8UK4
1LsEH8xXdoVt1oumpZaBwUUDUxJ/6osuQ5o7zotk0kVw3dqh3tQAz06JyYJ1vHnOdmXAWFkeEpmP
qfmPGJ/z/z2CbtL+KyIeRTg/h6KfP6whUp2TkzQZFnLfra3VF0P8Dj7Kp9ZUSHqTJIq4dG/E08j2
josH78elSVzDlof6Geqv0xesJfxzNV0GjDXXGCD5viontZGVcmvYb21W3Rr4Nk7P4sCAg6MF5z1U
VkvmCgRYhrkwa86wI3ehtqu1qY8hZTvlgIJ21+frjJCNL2RoCHrFxQWNNgkfSvbaUYtoQDx5SyaN
E1ru/031k/uX8bMF4kEkcAVtiz/FHNT7Yeh41dLJVVjAZa4wfnd5l+Rmq3NL+NT7BVO7s7J2BUeV
CgWEguG5LKQK3x7xix2rRK4j80atEwxPezsmoTlGIem3ZESV8iw45kCrrmDAkOTMz0e12leuzqOg
cUEFBr6RrbJuRalCYdcJd5CPJ+Wto0rN5HsSBtYfgfJQZcYczkIkNZDngF3PlkFsdk+CXxRcPgmb
dbKwXsUaNw5EivRcVvkutYqNgYPZPZ6swkuKvjAWKAL7bxQhCFwxC+LbyS+siyNTCPIGFt8I07FQ
pn7W3eQ55+h6JRbbc8dkMcPaK2vBANJ5rq7l+Vu2VJqY3LZrTKbscjahQFMm8SoTk6WrT0svbUCw
1MGExpuDu3wWBDo70+CSVy+0tWsW0LLuCVQYVq4bfbNpyCoTG5QKXuegX14F+wJv4j9yaP0bv+Mf
8nXN0IS5xY0ehntHXKYtOmAdtvBmKIe9xLUjCREdu4SK6EF/2zezlSIvIUsh7aqLOJ4omeBy2N27
5AUNJ9G3cNBIr8PeZt7DNtrxD/4QOU4XJO1bYFbyGSC7Qjgu/zv5S7TtGYph+rUWZzpnpctLwmrn
UJAq5dv6cvvQ0cdHRZcEpPxei5o22xjEzYvRHMmaG4I2AJTvGe+PgwYpWBQXmraXvu5ZooeiwCu8
y/zBS9uvp4REISZ3C5XLt0hv0rIL+62y/DjBobKZe/WldxavarULUC9ndew22A2FwaFZOVVIkEjQ
GwXYGn64gQ02OeC8BF2AJN8fgQp4Y4KZuZ9SqmaGsnxZxhq0qVLaH4CiCwhCZqs+6UlaSeCzkrcc
rwCIS3JQGHrPKKlUHzjfHugOnRUlXcAkm81fLAxEDtKlA3+V7buZVYoE3jAaK9hrHwDNo2JeV6er
VBv2+sf/HGpC4UshhewzWTYoM9RLRoaUXFgg1Jok9oEHsX8mOK2nbQa6O1SAceGMMHxqk45bsWdQ
GiNHB/pHYVM/pyF6kOANtqGigFZ3t/NIejHA5ss17K951PGa614qK9qg3zRwIPDsQU8G7Es449f3
Fr9xrP2fi4yExUY8nL8f2sZu29ZO16Z70jalULVxs1di948Ecc8WO4Tn6hHgnzHFGEb7e2AhyTcL
dvotTyBdEyuYgEtHa+i+YDRchE4mlm4F33ms5Jcewhox6wljKtO04xShd5FBIxrJ3mP0MVyNDhnm
Ju7kgXTlFiGmxMx4YjCljbgN/GT8wtGVNiaA0zENZxL4KGPbL8h1ozVXMKJXiSO4D3nCJYcewo4Z
sfQp2xqlcJqYHVSSmXMx0m8b8FXDDiCivs9Fji8JLqEqtCeEeoQSzlfSdwDTokbLERVb45RPGRxN
42xFU0vqD8+wf+tJoDettraoxep6qe86Whx4dMlI6AuUaLJs7S9eMYN/eAwUEVVgtVZyzjOBZrKz
oneJ5uESV5UxpysGkxf5fVyjr2syPlRIEBiLCEep9I+mtXxifx93mkf45u28IxwazQD/EN/KcX0w
9/PLg5Yj2vqxU0i6l5ogirBKfXPo3hFtdN7lQ99reTjAPwK6lBWvaWqu2J9JzpX3APiYhs+f6CwO
iM7HvaflwLx4zbDQdGJZ1lufOqvRM4/B0PbND0J6IG55QBviZFngnyzaeOycy/j200sX+Rb37Uk8
QHMPKiaIclitY4RUim/XhLXx5TgSVrx4yncgxC3bpyjytQkkwMDvSWPNzgoCvZZK7tgnHfQxdjlC
rlVX+ILiUGfx78xaDezXgD5XJhwsT/uickDHPXqYk9s8W6Dy0TeIx7OQ4Q0ve4U7JydT0NSyP/hd
H5HCOJj7UMs0L/CaU4UkWlYsmNeTQRnmht+k7NAup3OqOBGRWhWIVGvGEseu0arlBBr2OZYowm/d
j0zS9z8Z8eleyru7cyQ73N+Tuv1jNcXPaZMMI+TaErUwgkAM/khvw94AxAEhtfwh6V1mLwcEB+18
BTl26/2lO8GsxBWAWpjQ/1vON7KWC8JT/AmbOUo4LacNdmSVuNtEDu5ODddlTvYdsl8k7TuS+wkG
dQhlLtuluM4GsGw0n7jFX6CrhSXatKk16+/Qa83neUK+nzWOFvCkn3uGIvtfKSjjUA/PHXK/1D4X
Bmj0ogbu13gZFI/IrDEGDaYcfcBwb40K3IHxhEAj1OgpQ6olNox2M1FeIdA0xo60oi1qhYJNbeee
orNbEDgpOmcLEjBcJAis38FGoxy4NKihsi5MnoRBj6k9wWELaTnd9IKXxyAzEmZzWFqiA3Ze57iB
cx8U/PKie8sxO8AEJJoL0LStmbEPWNx3A3UNjtbMrA1RHOCEdbtVmlXdT704ox/ql4THQ1Fkm1PV
5WutB1RO8UoO71QAVZfwieTXXP6GaGQXhcBaS0sw76HpvUvzjWjlCPi7GHrbKOZTtSant4S9q8y3
XEthh+b5kr868Yg+38LIMkhJpW5kuCEEsTxIUKwfDEPfbnbcmGLVi+brzo2rhc9KunqW19MsOWsM
9yyI9Od3oj5FApQM4fK5cKt4H3li3rsFwJXYW+GAyvYu8Q0NiXbSuXikk/YU/HXyvFLjOdBiY3vc
09MDlE/0mIxSQ593C2OSdNoKC1xRBSobQlt9jAniJIIsgLu1JNtEp9uK8X97B+/LUJAB70VKQpVw
aoxHFzwrRndFGUp6t8mCqAf+lChk66C/axXI8hhkQ/HH6u3VRkG7PmMh2JEKhDT9iNAXI8woJUWG
ArVgWtQOTtp/ZOHzjhonURdo+9Vf79+PCBS+Prv2B3+U+nOcduBVM6w5c0Pk4DdWOPACHD5yHjU/
jyiTeRRo6qWlb8Rqe34fWMNyRiNP+7vC/LKh7DSWJfPdyXfonVpFGYaijU43iDYME5KCf1Diiwhx
r3UqeaGTaUif+BbLbvFpPKt4vM9Z5hBaOrmWulEWX5TyWlYV4R5ewfCMyfUGV9t+Tw2iATG6MV/Y
7YyCU/t/X0NUExSfA3OUxyUBJQQ3Pajtm0o2YfYKk7a+GNKmTNkmyXiblApItjTNASuQuXJk3uh/
jjeR8QTXinRwfdkxt9rYZJIEK6CnT9fPX83rTTTFtuof5Fc1nLWiKKtdZjuWETzkUu9EckdALMWn
B7UPxZiNVnQMnMvckeOfOmyV0zZwg0Nw2tW6ULto2skBbTtZVE6afRPQoXMnnj2kLmFLVYaPVoAE
vlq2bpgtpaeRwyPd2gdatULirhOA0eP/3cI7tDmLpP+Qv/iPebWH2IFYi8nGGtCYoOZI2qX4vXnZ
BpS4LwJ0e3ADceafHXVAbd6odBH/fRC/XbMaOD/AUbjYXtPzvvx/jJpyEWm3ryZaL/Yl5PMkBbFg
M2aRkrTMEyC+AO8szFndD7G+CTo0crxYYXMrnt+xP6kivkQplUsQVaplPTRFQtwKo+UyHM/rgBJ9
XKdnAVA5PvwLi3K3h8tFvdZ2xHqDOmIxMFLet+/EFd1AQjcztg2xEV/rqY91wadpFjuViLDNrDTg
yp6L9ALtKHKA4LzAbyXXJZFBs3UhUx1dajWYuJ7TifIEKpyaW9nTqjZ+S7IGpU8DobZJ6l+3owlA
swum/OApyLRgn3wMJgpRpYry5ZWXRq4GvOzHZLWCITgeTRxE6y8XGLfLjcUgHYkLttGgpftKOVe1
rwJ/HGJVKOzUkB61yNPrDsrCkzsAhbvgnYXgem8OdbA9+Fm2lPoT3aX7rxQv56oGpz9QmFGMGjky
vi51PiDnUOsFHjoYXbm0c+Vr1do0+7BHee3bXvwmV8vKg9L/HxJKPK+9VSHrcTo64XFmnLZwngAf
MV8GuDiyifWE+SXPs1prXFRqHLuV605VOWV97p4gVRaTqwOwfgSmHCZWLhqCTa0NLPEnlFCwrT+x
t88S3iQa3zc2RZzdNx8ADdGKFIYFLuZQU9dvkF2FSwxH/3J+7l7KC7t2AURQzb8rWMJz8FDhaxpK
oReZ1AwidBDw0vVVk31fdAZ59c31Ilil70qjqifYu3gx8D9EAodQsuJPED9QtJvleP6DRP2GP0IL
glVgqFT6hxxPbz3V6Yy8ebNJt6YFqRb3oKkn8pV0BNuzdK6dqVTZTHTKv+ca9m0g2Qo2VeYBzAZp
Yqy6rsxo0kUKktIR3+roAC0Ew5evBna6SrStoizFwvUmAFE6yeOrODxh+pFeNE0+jmh7JojiYtzC
euLNEmePrBjTnsV834HNTwfTEOHfswf14l3/sTlD0Z1Nks4bFWrJYl8mZdAPKeiFb4wDnY5dwUfN
K7Xmn9lHWCl2/jjLtFtaiZDtKEIU50v5k37ok28bs0n8EQKHXHZP1ehfpakaQWiVDxJZUhPWTznp
SFVeIrV6flT1QgF6uIsgIkAkzK1CMlt5e4PLfEpRhKy8khGsFJqoLwiOFCSaj9W6iEH09Q9mt1CC
kmwB5B98BMORxv/W6aCLK61lPynbdnmc/intFIKB3fzHRtOoADlafKe6pbfcxmzRMD8rIB8gj54i
jfjGa8jN7ZmEMQPim6T6SVqF1CBCJIdt7SPrCORgiQ3doak6WOHKaKEqw4NDccjeCAKALoEhxs7i
pPQlSpdqwCdJbrP2BsSN8q6J2bxy+XbM/ST21ksrpJsTA8UK0NiqhSxuhk3jZ5usWuwvSPf+PUPQ
womZtgck8txPFxSkiha7QrWB7V5CwP639ypxypkeaUfWl1w601ZZViWg4fDNyh/DBYlBUQUmNh7F
+lCCIJCe0L//kkRqLSGISGm8zTX8umBkHdX0P+U9yURlTB29lvl/hGf/ksH0mHPfX2fy1riq+HJF
xvFxQsqJIjgYhnJQuO8V/qKDBT3v/TVc6hrF/Up/ATgDjHKwhEmFn6OcVj1s/JHmHdqGz8cnUL7F
txd4vgHE65u6qh5Sg257hsEl03iUYSat1ZIyjzbdUXDyVFk7c8G1rOkViOoiWyhC0pn9q4QDiV3+
NWP5wGBh1LXyAZfY0F/klA7bmXStcsAzEKi63Tm/JcPYXZXO8iSEVr+bDKw8/oQ03ZdhAi+tTzNg
aFrqGmHfvarmb4CsrulJPicYqrEEf7unqYWsz0YgKgDj/pVWlraFDl+7mbTIkEfBXBE0c+LMLRpO
CinsWGw8gg+HI0X5MqIVkZLzyWnCiblliabliXn/yrZhBqPcD5t9pZ5EwaLnAY8Zok6q4htie5L6
N0EJOq4ekcnxPQeu3y3v4b9FPmiEvo91EkW9ime5VBHbgEKgIYr7JqOxrJFKtwhnBJZtb45FY0X2
BxG0WiMMw9BXWEvR+whrN6wzAr5e8TPrLlSRTc14jpagsf6b2AGhEMRUcmZy6liIPY5PAuVXY42V
ZZapT6QTXmeU6KRGc/zY//j7WSlKkkNq+JL1Er8yXtAGiJIJv5FrpdQkJ2AwyFN2hz1nm+OK/76g
E7rVezbiErd2UQDt59PLHffleDLuX4cnhzkXlP+jGhTu8E47CsfGs2okMDyNvPNtS4cz9xgimAaP
IAbmcWZJADVXT32htFi65KUJvVeq0dU8StyrwLVHh87BkM57qZRXAGHXWZpiPHW3G0h2hHthF17h
dbBBKCachwuYedK0nHW3yAltNuMQ8w57iF8zl9QFBsJDKiZN6Ir6uozlaXyVIdX0DGjkN5kSCAmB
CGeewuyMibmD6rZIyZKIePegc0vlOAwFjbNeAgA3XCqi7B4jcLqx4/VYgd9Jq0z/gsa+H+cMz2bh
kaz4T60t8dxl53Sfm3Jn4PlCN5P0X3qz7+HVj1CR5cNivDi+kN+8HeWkaxXVhaV8pMRRGkUFC/EB
Ln430aRi1Vb1zBRsCciCQsZ4YVi1gl8ujcdawLh1vEZWgxLT5nvn9mJ2BNZau3HPeBD28HyFUY4H
LA6Za09A9mSjjNFh5Ndp5CdhZci1bRQRwJhsDULKO8cRHrmIaYajjWOuLF5T9wrLguSrsZ7GXjH+
OUFNn93aFwtf4tt5I1E08f0Jdrs/Z4w3SJF2M/4Qjxh1z1O3k+zhodHtdBHU97UBDt507eJ92aPS
uuZ/fDAbspZQYWLEWnnO/lsktHwvg0aw0lVARcT0o+aqsC6kZV3zX/kiZaZJWG/S5xSYPzamlMVM
x86MvA6fCxEPauIziadSr3RqsJKPZ81Fupe2w6Yjp9gkHRo5I9Ww7ZHoCASjDz1yYd1lxmYGwmWU
9kpuEIxPjYOXShb9zShTBDSZsTQjxkYxDXJCH9yFS8xEMCZgeHlxrRG+d8GPrYrlFRmg+qSr+2/n
bcnAwKdkD6EDKzBnoJk9VvB2XjN7ZYmK/S/IrzaFVXMeEye8lH8q/FAi1zGAynTazZZg7JpUP8Ye
W6C2/AFFPx4O4lKrZ1a0GetOvUxDgBU6oOB9m7EMrH27myR8HyeUN+Wpl5h7cdxWRhWYNYL8QQ2i
GTFvFhJ/ZRhihq1krdWLPrRYaMvvjjxf0DYkQ3vGyIR+dBL5Uj7gYYER7O8DBM303bMobiOGVLct
0JrwDGdfegwfiHzp83JU06y8KvBfdNO8EA70Qs7nV/mpwFSwyG270/tGrGC7OTvg51jnF37F3W8S
4gHTHvRbv7KRDx+uQ8YxxgEIEubnDmJBbf5NzWArkmVUDbGYQIFVjW5N+doYyDsrQdoRPK0dEoSj
rfsBnxMft6b98mhLUW2/gjAnvMgneOzSWBsBUc67+lR5iypuJZ5pdPexI0Ax3Im4lDuVeScr7OpF
ZW9gCDoxWTdtLfB/VYrhGNHeTMZHiuAiDcWahLHiLXAFjbyEpWEkd2b8CZa8cLXrn0WXSCgT82cX
AsbE7Gb0kSTGu6qUFtkAUfRQk55IcxQvlUOd8loayi2rF0clNToTw6XFJ0L7lQ5qIm0NcYa7wq1S
lLqwlefrOqfBC+WCJ35v23o4fLJgRJFNS3mH+Ow5kK9luD4HxKd6cjiKPJx8PFFeBDBZ4gk1qeAa
Y7gsAJonwuk/rqY8vqS90sby97AyH2cDQaetaWn6LmjWiEWkk7Nx3I0MQbEr/4rnaHmMhuHExm71
uxsylrBLi7YBps5a4rMA7469IsPi53CoenBNL6/lZr5Am1Rw5R9Pz0YGfL4LBhTuogtXkQCvb5KH
r/aHAiL+eZvLLyHrHBpclA8J+wQwOMMpt7srRujaJFNtovFZcn+agWRUXRYi4vz432vE+tAD8Yqg
EaSeVnx/L0KY0D6h0t5ux3nsGG+AkA5fBxXiTaB9OItBG9/SlP+1twK4UpSein0IZhU/m3No0C2W
3uoOfJ56q8ca3B1mFhJ0UoQdBQILwd87gqVZiyIJrij/+c2PtAoOwt/E6MPWgvtJ9M3jNqxMoLgZ
P4wpWbptuwU4LuGkrr6H4UV0xeLIXgaLTMn6k/aRIuj5Yj3/6U8VInTcvr9hremQvF+42OFkrf/i
DRnjmM+rc05YVuVACi0sDT7HPTplsh5XEUm8Ud8WzkFAqtPVEBE+8Zo83Pb4boKQiYbRj21ai94G
qE3vN3HVm7oI2qO6A7OH7OzboVFH+60ZoA5PvDZN3yG2giUyWQVMsxr5zd7Sg/v37EIWd8NUdTQL
rHCGstOhjIMoDeAwSc4rGROtFX7iz6MZffsJn3a2cblqdaNqfwR99O6cWyxdxdRBXvCwXGam0CPg
YOqHife6WU4xHUVQw6yWNuWrX4rvU5y4yNG8pnYIfcU3zb/vIPaHWsMb8sf0Nl6WeEjQn5c7cIlv
FVhlsKXado+LsyCYli7J7CSZClDkpXwEwH8C94Rz2+2EF6uj4OtyFPUok1/TyXWHHFSz0W2FO2Jn
qKEJ7/1eMfYQ5eOwgekUwa1ppG2xl7xsfl5DDNsA8BN2+wzDVWZUvrgXahxC/jWaGb1lzZa0GD1H
RWIUuhclM0RS2xOLvG0Jj9zlgh3fsMjJQdGeKeptcrPhIM9aNl65W4vNuwEwXeME/CFdcybUW9XC
sg66Wyv8h9Wjl+EvBolWMQLgl0PvQQ/zV9ya/QljZeRy5qgfv19z1Y+LJOrdd/3KOI7VtqKddeA+
Qdf5LYs93jvIP94xNNxqsbDDPmJIRWZmCsLp3w5WYuMwquGq9beEkgILkOEctPSQkFo6PWLa/IeA
x1GtZu2qEVo4JDo7vESS0qvJndZDulDAZGwWM2zQ3h9a09Stgf2029k8hkgM9MzQVnxZummySJzE
P3mAUPl4gJhb6Twlgn99fT25SUK2/qTRcGFe/9U1N3w2gsyRhgzXeSSuP46pGlYpQ8u/eaz80lAb
5707NVC8qjpkAfX8p8DWvoqjjMSkvuyoxHk/X424d0GV01muWUZc/aYESwscdbnTyjDEUUs0YjUU
Ga0hrd7+UyWCLPtntuvzRZV9CXJ1cEMM2zMzAqwO+Kbg92alMkAtJZuteG08X2Ts6tmz2CD2M+be
wFaDDAJYjk37LgLCNpFK2+2IvgOIjBO9vBbli7lLHvIbFpLToUOLfyH9vLB4+igA3hlI9R7LWafu
OtRoboWaZoJ7N3/aJEavRwcYXVq/h3gQ5Pxtkn6JdeXveVIxhOuxUG0rSO+peFgPDolP5yLRXjl/
fL84R+wkfxtHpVvnZ7K5acTViomIZkbGsF07IVM2RibQMuRwjnZipsXVinfwPOZEWDoBzMiIr/M4
+kaEc7zoYf4mpr3Ymo2l+e8iaBlb2dr2UJ6O6bdXSthqC/YQM5t6Yf0X2UOCuuzUqU/UhjjhlMqo
GDTmZNknt2xl7Ot6ZGTpb3S7+Yw1EeXhFZ/DpuEYFfMYyccO76inO6Wz16anKGuEaY1/wAirGHw6
AsBn7XgFxlr1P9TYJIti13IGLbQeZh7+X/fcrtBtrLErE0g9Xop4QjvXL+pqNW4J8JMo+HFQCx1c
hmpO1vYk0/Chdnz9L6O28qRhhqGSfMIyz9e88g7u0+IUPsJaxxySxQkvBUnmCtRbnd9OOio+lBXS
yi6wkQ4jAAsAXO0xLOUt4m8edzMMMdsz80zkuM8YWi4UkT3z3p76XO4GQABiu0f/MYnVg7yLt3mX
Gw1d0SZ6u1Z54VmwSvqFurUBDfskrxPAenqpHgMbn/StTfDbgFiMAUGqP/Ae5gaiaBbLiEGOeFqa
0B6nGWvHuE3dd3rxUfuQN1HSXTTJWj8hBuKLchTh6qCmgOLl7OyDpDgknWqXPpaZuyNZIVmYn+pc
6BH2QfsWpEmN6CCeN0XrO9qbBNPLHQKvZUTPHVs+B2QRxVmXYtmmsvL9LYNnMSBW46kFV/SKScxT
MSjZ1odmm14NPUyYp9Iue8flTQWrmafrPB2LjOZn//Lvjr4SgGiVL3qp9kXK3GK4WWA5jJoZEmMR
V378xIEWdV0u4iSyNNbpE+7s9/oiYVKoKA2J4ROMkweJgLWggwHlDs8/iuqcQRfL3/SAeNuXrUTO
YrfnJTOJPVX4m/J0hpc2arnZlpQKIWgxwGPEKmGaEWzVpCRPJSLNHTXa7Zm+qSBCc5yX8+RKFCVt
dzko8mUQZwjzfGHb6/SRlbv8zSzeSbA2FrWy8jVenExiHFV+2CFI5ReeC+7FvPgAnBkE+QmW3tYU
Tn14hcw4mhI8HfLgZWR+xviynsX+XuBlKrAhBn01t0sHqv+bQ9d8WWFNcT7VCj5IThdfL9sLzVdL
4vCiyIiF7ycspZMDKk5qm9EH+wRQFDMvqHY7uE1D5KKdrRbS+X4e0OlhRldbOArxDGVP6PRfZZ4e
SMBGqR1F6zx88yj2cvgIMf3ubj/5MI6G/Ve/FHCsAVcX/bgv6SpFmLbcAW/XbDDhVhudaH/y2J/8
r2ctN/gOD6iYaPST2/HctP9tPbyIxo3vWIpnq1TQUGDDi9fQ0/4awz0tdJ2AvSdAqyonQPidJVWa
l3grIHEOf5bMxiVwSEkFyPNguiYROluvE3J4qQ4bISAKGsQbdNO/NgqJhRakFzqiGmpEfNW1//5V
02yBtQdNFHC1N4R/ok7NCM8+rCUWeBnJKzbpbkHrWo017oLq6aSsf9BlauzhQBFYETZzY9DK0PVx
PN4V/3UwnrGBPjO6lt3Uu0MhOGjvJqTZIUE7AwewxbWKOLKNRWX5q+T+M9g2Rm/VkCs9WbJESn9h
fy+ai27yxpYMJo9MuL8xb2JYw7XRIeDmREJv9iCAsQN4ZuUlIP9nmPY6uk6yYZB9ASzEaiH1zkGQ
FpgPvcFJW4+Z2/P+xG4vpR0MQ4/5FfHGFsJQKguzXVHD4Jd3Nr2qI0BXd6yWOa/wxZjCspOGJhDb
+byK5fC3NTxT/DzHn9XrmEoDyBMFlk93TwZtmNy43edILbf1mVpMGMIrNDrx8NwgdKne6FNvNIDS
pSlk6ZtaoZX6VnMJY1CYV4qhZLH612O0vPTUnv9vy3xO9J0CGG3EaBM8EOxmuWtd5kFzV4VZd4RG
ay+RaKYyVTD3SnQcvDvUEGKvUFIVcaQk3VO9FrAjgq0xSE3fuY2RPFirZ9Cvk+/lXM+QCnjvHBFU
CbHQNBHG3zCnujTNF3HowY2psCcS03zbF1UQMcwQHgo88CaXhJs0PSl/dGZXDqE4CAClxRiIryyu
WtnKXa/KwtN1amztt928/9pUGZyBkb+7LlswcsOIiK3H1+vys4M2o9Xei6qlwvwiCvD+RuLy47IU
h1EDpmN/YsmFdk3d1fmN++wpfYDydeNApi6orjZiphE18Ay/somyMFqr6GQtXtHMmEpCv6Z/sHNY
tG4Y7IhA9x39fPIZPw+phcyvfryclrtZV526Teh9s/f0G02c5YccLEws7rcYzwUti2nFf/aYlq9j
Ku5GnM6/txvOYybAwEM1LLjzuGHEEPuJ0IdUMVp85Va4xftbroiOKKRDSO7q5M9+3P0YBzL+J82t
94qejgHPfimEBMTEYR1tcG6Fbt5FuDdeG9r82M7ovGCfaxHvz5t7KMlozmBNWP/w+tSe0mj8zX3p
EQmr8Mmwj6cQqHhoa3tbFK/FHEDjGqwJx87c/0Ig2fJFuOfqlUik1v2n4x5SK4HAlU4JyHpKl/iD
MlYaCd/LBPUSI0athiNWbMPdihyHg8BMvjKxXPRE4Wuii5/bYU+rk48sZ0I3qtru1h9chhS9Ge3v
yrz+NdxzKn2GdR/sW7pELUvqCWmoexQMm73eQoYwkyTD7r7ud7XleIO+KS8tYB3IuvdKAoC4ZywU
e7gGBQ0t67f3TY9w14lqJJsJJ46yT6trIzTfO+8VAE3uz9c61nzSagpVOA5rtCAlNFm2zhAplRna
6Y6QFqrJa5PU4Ppj0c/7dx+onE3DWJ4fuCpbZCfapBPSJwdNgr0wwkbpPezBOkGj3GAxBhOoSMuD
astQBTkfxBh+5FyT04y2amhTWvw/wVecdSxFNl++SpQSxTJVPa5ahKl27FhAsB/BeUmx6R6l7jIB
OVwAkbIR0CLaTHk5nLM+7LdLv9mx1oAWq1uo/tG7xmpatLBHyOn7PWedPr72BKmxqx0OYpm6VHeB
0mJwCn6ylbHcwGF60vpyFmffB6hpySQ/ElLsBrGD7OH6rKDZIdo80y0AYBnvg0ah0WokJGu7ifAp
edj78Pg5ZbiRWnxF/D102g47OlN+mA6/LN1L9VhAhdrPlKpNKcM9LKyRkZQGSaM2jF323payO18+
FpH1vIJVcSOkBQYlwc3ZQCp+RpU2zGv19RHvfhKH8xNAuA0fgmEZBmWlHLEpi75odkpzxw73pUUX
hhf6H7NY0wY9vIn5UoVYSe/UXS6TxF7FgV07FQq2I2Od4NwRUrOuiYPJ8LPaUb65JlClMFhNiZZ8
5icsd+JJZMPF0XXIZnfi9C8nZGmTJBG+KpoRhrDAcMQrJ+hi2WHzZvAjA2slLcAkzYS1nxAGqPBq
BFP6uUxjWOZ9D1GtgCnAsxIwDfzslcm6hqOnEu+SfyKfoSiAVKJIRk1ntvErHckHXaf9rRs1t2o8
ObCFXK5ZTgORgYuzkSbtP6Wrc+gjA4qAIcj4MIWENBEp8Ujq9fYOqrOF/us0N3hzWOaUJ78HVZEr
K1PiNh/euO15om9vN9akuYyTLUTtCVqrvHTNpx1gXMgOtr7DMwVWgLJhr40g68Ox2opEHE5pO1p/
9B2hHPjFQ7fyvrtCTFA+swPaqgCQndiJnvop1gwB3kjkggbJ15WI8R30wz3otJEM/bUlx8UPRqin
bGvaUdZporq0Vtt+VbZaWaSUgqTDKkQu386hSYi4pbaNQWZka9+M4Im/UKdGN5Sqq0my9YayArAa
OF3sQ4WPSnwwWtbC7pGBqDmQOYtjkmUgu9bkQPTmYBAsgeVdfNeFPEd9R7UXZHqVC9OPvLqM4xTD
xPqper/36IH5292GQgqAkZvnF2TUD/Q5DCjDWWKfbNTP/l4JscqI9Tkd1wfKAx17XlPpdz+had2K
PKP23lzqVfMx8lvbx/7ZwruJRaIjyHbCf4C2IdmsLija4+eLDCHaj/knXSJFjsaZiTXzwxfOpAXb
hgzPRdLA95GWGNBexUC7LNZhHITy87RedR+3gSkp+LWUbCDU2iGlm9Wd3jHWr7CVPEkEfbulEZoE
oJTHOJwJv7VU9aNjggZ6HrzHgWYMiZ9+WUFRbuyY7sqaPmQpIRNnu0QUTTxk7ezOhxNcrAgPtXlw
JlYfgB9S8J79qLagyVnsJ2vL4SkZ8ugLkVRLdPAAYqZFZeWEQpdOQCkN2onhEsJ2WaIzPe8e5g1k
gWlf1QaEivPkICFFSyGCFXuEzT03fsZ9P4Xv0yezvFdq4gaLZn/7d1PSuYX0Kst3N0xekNoFUKXT
9i40Y7LKQWLxmAkU2LE+fqWJ1R2aPr/vbqMMVKHoLUkTtKLa6UBDBYekeYudcuvozkaLHbn1RUx/
PLlpuslyFgAXppk6RUDJuTgSl7nDyTaZSrAvUkDORJMC9ruD3Zy5BP35XaRY7VmXzYEaGO8r47U6
/BeWnBci1Za8my+lOrVvy4RVFuzSwCR95d4UScREt01cWjXEVodaS6M8sL11AMxRgeBYJRVoSWx3
ytSd3JeJTuATvnMeCU3J/aOrC6+605gfT/6XZc9yaerXbivF9ILIO53KM43V4ubpx6a7RBaR9vwT
z5kx41L0vr6eDoPwdGF8Kvf4ncfI7jwA9mvEmSSGzfSZqpYYvZ5NKW+5hp8DY+wMdCOwzikz4HTs
IS8vaEqbIit6JYi5AVAum+fFMgHxS9u998511ugBu/uzprmeGYNZkXle/3MS+VI32/vQEZQ3JBm5
eK4l1lNJtpeBFyMJnSvhzumr0RfZ4GESYh1cqNl1AL9+iscMfZkfsk6BPeSfdMUsnRsZGt7UHVPP
rnv8alT2QQvDOgLQnONgmBtXOp+0eFLn6E3bo6vu8WSgNiO1c4p0rJBfaOxwunA63oXk9NbbNXdM
4WEboxqiF4DCfWlhZLcRapJEvdtfBA5vXzjopDZgUerMgflh1Z/3vERM0nvx7XIoSXwT9EiVDVvR
CBw9Y48EL33mI/yhgUR8O2MF0EahdtxlIs/1yUXiv/gvtdbStlbSZoVw+55ZscoMwYn16fH2Au2/
CWhdZCRMGU+rNSQwRbBEWVZ87DnTrEMVDNrGNFCflFnKQohEgIrsiW0+K8Hs1iFinwRwvwqVkjEd
eWeccSSCcsAKWvEAGfZ8y3Ib5IujrWgy0ySVmdlkkX3TtoJU6h3wh5b6opK6Nm1mWU6ryDFVEp6r
FwJ0Iqy/ckiAFzu4hXrbQvSMwj0ctp2i7eTS5qs/8i3tRAylzss2iXlUs/bmTJskOdePzZ3ob5KI
ZKPHvOenTxCK03yFknM55CTdsSCtBfrihOp71Dzj0OtblFVLV6c04rrRQXAUucZgpakzKENHJL/+
ebNuVOcfFW1uGo4G7AdlfO6JCFMxpeTvrCnYS9qdIp18u2K54o82qTtkyE7pWgWb0RxLDLa+Qjfi
qU3GuwmeBR6Uk08Fnwr89tH2VNiMNnfaIWvaG24Kou5SUeXtL9qScpBOtlO+O0bbi7BmZ92wuhZq
qga/ySTlddmF37t5Gbk4dByyIC1/o40HY7zO5Osj4NNYzk5PuKPjmuc6xwagKo+en4f74HEkeRTt
gCqKwfszxDnd6BDShYRMAygU7ql7U0yu3wTj4BH2xXr4h0hjMUe876O6bacbvymiIPS+q0N6u6pZ
qG681UY63TVM4DqppZXMOY64WD/tWfilMNztJwFygS6sfe8l4lHeiVRDMcWoepPoQMPKXTR5rZAj
UJZKiGioXkox0R0Fknr7P7BwC7tKpOAp0/K7oT7ascUar80dbzoY9n5wK7Fr2kn077UZPcy02CME
fUYm3h1qu/jAf40l8IgANGzz4H+QKUhuBOyfUVtoERU756h2Hl18Yqob+JXjEjprvmAO+/Sqi8K1
FC/h9Zpdz2UQjM411lrKdggQjFXmF0RlJruL8mDQp9EaU+sg/fFdfXpwt4/EEX4yypvir5Pf3Df7
goBmcreP3pusMSA84MHCsoP1xh0Zf2m9UXLfAX7VBeMaglC9Iwmy1IHNQ/uLP0QyW2tyZncXdD7S
IM8P4ZFAAnRVoysA3C/9HeGIivq/ZyTQm1tbbsW4FvvMVLrAuxrUFrJsEP4iCC5PoT0dhaEdfodH
CQ5U3bEkl12qJFKKUlBr5jQP6w0xuTVK2EaYet2JC56W8OX4H0iRjxBbOUVOcF3fF/qwdslL5p7I
i+iOvMEvtDHVgma+0H3iZUmNj+PyK7APUFTAwLiDEWZWgVUIYzmL0ICtXyVsAqVVr8/hpTOB9zNj
u4NLFdkfogB0KyC8dZ4g/epO17gX5YNrvhwcS8n8bfFlXNws42/nrCKkoTk1gxgII+UvzdlgCL1T
nXZEB3Vvp54Go2bTfR8XfqtDR363QcZQ18EFv7Gt6WcvPbuNVO9YpccUKB6VHoYsYAVMLXRKuon4
zLCUiYMCEnnkHBjvLHqc6xA+5UwcrvrlFYvciyWMCQkeWcTLeBwmAFrr8ztZRUxj4tlYU1/0iDOC
Ztb5K5PmrPUG9N/6e2DdutNsxjZP/HSI0oHxWiKvi6ukVsRzrbJQ/2mtKTYnDjPms1boMevy+2+c
aFNteLbsLfSuQ+sA+rcdLm1P2QgYXxqrLzBfO8D4z+ZlgJQj/yC9MB5oJBY9GCSQ/p/hsoVw6d7c
n674YqMjfOmfFK//LZ2Jt2yK0Vvc/Z1AK1Nq8ACvgJNvbFFE9hE9qcxCKnewjUPHMKdAZu2+G/i0
88HMzxqqwkgAAwtXPYMcZ3FWJ6YhqlJFBun0+uYEszayTxqPwibdKNmoBuv2oRgOINgVR6CZljpX
G0gGqVEeG0Jz4yJ4HRlSBt6xB1eCc4VJK6OuyXo97kXhoqI6gY5afQx9Cxx0WlBUTVwgHLSGSuqU
MlmvAuBGkxK8SwkNpsPFoQDzitP2kwutuNGInJUe9ZLiEsZ5hcNEVJnC8X1i4OvHXfWck9uRXBB9
bTMtHGna13wprj8ooMtuoA2sC2LZZJpfZf750ezhdW72HVgs44LU1Id23CQQxsaDwB0NF+JBRWzT
1x/xzpt0boEDSERL12PMz09QC6QEwjgq3xyMGFdpp8Yfd0FauloOmyVnA2xORyVr/n11tr7nU8lr
SAlYIOfQSLlwWuRHCF25lvCI90JDXKoY69N3ngg/3ebg1yahmoqF/I3eOVqbNEKsRsvREJAv75DN
BH0v0WnKNYxnOIMNh41Y0xnw5tKFoyL8JIKAP4B/RL85kbBd0/3lCyXBHkoyCmtH0/aVIlwHdwW1
FVnVEd3ZqRKSnSn+iP/bKlUefcGMrLEbiop3RUgBGKa/aMyl7I5Nm+SiPdbge1D4BFUUsjNNzffc
bAn+dkoAOXGDi7GwgxB+yJPKv+DbMcxAYuaX/TD1veaQVfsEoidRQUoNBhwZJkm94+cqDBDUe7Vw
M4e/L2VqtpdYad6N17SVENTLUDUix74gL2v4ZJqW6HAUrI/2gSC1xVxkclamropE3J49WCMkE2Gg
FLa/9HQiqO1JvsPrh/8RMf/w/dI5maUT5H7rujEulDHwarmUWIemp2emrnXgpOoM3u4zDBUsijjs
Nq68fTQWpsBYI/e6AZc89zyL5+21n4A61Bg7zFwbJG7b7GWMnDj9Ebss+5Q17vjKSu/2G3tii1vY
VHc05giORozhgzg7/n9xLSJFjP9ZLIDCLwOdWFhsnB9LVuVU4vKw6Kea73Q/dHVoqk0rTjzBx1so
/lhcBwrOJXF7bXvmj5ohdH/6rxt0ULhKlkusRjzKPMEjtzCZLeFEM6S3CRR4OHM4EqmT9Thm49An
gOZvktFoXXAKrqATnnJ2nZF2/irzxBjFjxnaZ/+wO3pgQQBeQWcmWiR2HquAjzWce/33vMjogVk8
By+7O+lsui+p4T7wmsG+c8BYMs4L/TzKCKmUa5aXnmXuv3IaJKjfIsS9mAFzRyQuaQkBYPF0xMgf
ug4RY3mg5/n+/PWab+lNgybgD4TVldjBQZ+bwEWG6aDVpZSwDGs5u6V4H3y1j5yJM1dsd2C+A6fb
oGZY51ngLuFVB2S5NO2Sh15oW1GySkGFh3+z1gvvZVjA7d629wagRDDrknX4paVyTmIucYA3egQT
y1X+tUNe8Ht6EIj/vOFcaC/8DtMn/GLXrEXKjryGiNr6l5jPubqQZlUgpCHZR0L6XXROVsgMXmAs
wkUrxTUTyGVKf4PaNCEKorOKVSOzrWTwck8X46vR9SNN+1NHATPLe6ZPYmHHU/XaTt+5idjrhX0F
HINwEpkDS6Ap8bs5C0LgqiVtv49t18g2nhaRV0AGESA2TKy9mxDfqE6tNRh7W0UJuzxy7usGWMCl
2vI28zAlJ5g0IhcK2lv255XFukLqDrN/OiLLG9lrCHSzOx+NVC1QZj/yaEA62f7FqxaK8XS6L4eZ
etiPaRrDrTeYi1RCyZuXZ49xSKqBLqYwudhCZed6DAUFWwHAW64GODZXmj+8YVYHYOUpevrENWBE
1JL5Oe6QAS1ORUEbB/cQPWxDC+7j4uv3ocXFwxdyezSxf1p5L/ohHlHc3hjEcOo7exLDegiVE0rc
YpnIgdGupfN57RUt6nlLkSgCETQrvU2o2kbpatJ4/eaTd0JrhmdLYqsVfoi27UPj8wUrTYbhNfs3
QFMNduzR4YniVQX1Lp4xMW2pKob3cZhRJ35EEAzXbS7OTduXOwBc9NUTeq1ngdhf0QKqpiBL2nUu
XwzZuiaQc7DLSDI9bAidBDlW3rmKWcA4TPHXN1SdJMaTo9lzNmjzhr2B0fc3ejY3sUbweN8IgA3i
owyTX8WmiYG5sh1VsH7A8H5lHyv1S/nGAU3ZpAs6KERsSPdlAp4nnjts0IcmwJ+FvDYL1XjBkrQs
VOYM30TnfOf+Vu3YItgqseSfEsPbOKJCnFC0OYmiH0pc9TX6cqAzpGUK8OQ8wLMG7PwcCT+/atjI
tPlob6h3spiZyP+eUQtgWIVSu0Bcqp68+aRckfJLVnlhgj8It3pq/vKFlxwQm2Mc3lmhUX0VM2Xp
ZOg61pirsrI5eL4bWLCPfDz8H8VEHFWEJMiXw+rt9/0GzPcGy/3qpsXkZ3XuS2NQj59hRjCTJcG4
lXysbBHp79rPPq9xjy/WnPs2Lo3DCd+V/konx+qm6XW3w6/mpY4EiFxxvn9Ej4N6NQ8a6ewGRroM
aSgr0uT+ImHQ6f9S2XMX5PZndFTXV8EnwYNr6kMADZue5jzZNp0zCuYIU1nkGhwSFSPfqW1ls6lz
OZOyQaBQo67LGoJB1TcNdm55bpNnJkROxnXp17X8idxspdfZJpIXI+R8DqN4W79VZ0C6XSVXaLLR
eJqXJDBZmjAH7hTOL9K4u0Tpwb33ZNlhcdyqOXcgQZB6Cranutz6QidG/x6Eozl2GVnLYEcq/Apd
TqEaSEXBFmNXPK1Ihq53QPiPg7KCAOv5GTiFG1dqJtirUfdlTeP75P4Wuf8Nl9Afhvhot38BEL6c
pHbKFWMScx30aiSCkXbUmCLQmly4H7Pm74wHBW25ejP/bXNCJ65gHMES0afVlnd/PlB8VKZq2GiP
nfFmUn0hxyEx0KF4FedbO+76m7YVMjDwsUCA1BugC4FB4Gu1Rm434wWi53g4opIgfacSgGTOwoIs
n5PoL6laQsC/KqHgM5VtMf7/dxV/RHMf+8qClXrH0/N+PQn9RBTaf1+j/hGJ9b6QOhfvadDl8E+W
EFBC0iwSxxPatFSirc4/TxqEU7goPCBnYjq3nSid/ZP6ZKgFTr+j8MJ+OnYxmVFvlZH95E3nelpt
eRU5lOJvle6hE/r2ZXSeimLwTGzlYTdotwUGyw9JJGciaOCd371zSXoecXJEVwAtTt1RbXDcge0Z
5sRXFIYSTTyZwww2U4WuLFOmXxZ9WWH7NK+xBe2IupH1FPQjERE5VYP+g60aAhRDzU08i+q5QI1j
kX8Q5WC4jjVG2mEWoteAJizOSRW0FJf6YEnF47h13msZQyn3JFBP9RzxMNZPcjFpFgtc0/Fkn1da
syx+bdispCmTNsHQMtRdLHOgvhKZW/jYF5LBTsCIVdJFU+VQ0oCMRRRyc3QIoB48AcmNl269Vvse
krVBQi28pGrqm0jdHDU5ObpWKTO1J4o08OfqvcWOW2b4AYV01xvczQchVXBrt7pbOx+KZZTbpndM
8AVleJ1UMDo3bB4yYKd0G4uTW3o4900E88+8hKZLlFp0HRI0QCduu6oYkQ1JmUmS0jntQbc4K/uC
XFbsDjB3tkX9xx+ib72+CdhngJNDNJuiJYI4WEbcvv1aYzAiJaqtr+Zrx29QyRYvhvccTdQ8g3M6
0yLIECLF3L3vscAqjA1BYEy4Vr44ll/hL3XWm3y42MapTYOO7cn9LqRaoNOLvTyF6cle4ps0YEoe
KSijy7HFcPDquIsf7SiQFEnHWJtzTsT/TNePWfdk6NSKdVBWazs2h9FDIvAzKwRIS1RisPyRRLGr
YeWDGz9r4cqTlIMAwIsIqyidh1Bo/KtmStoa7ip+LWGw4wpbT+o61DDM0eVxym6gX4L5sT/v28uU
HMKkWq+lZhBP5kSTIfwklJUfJTPgsXLTVLVhmV+pC0A9LcTmoYkkiwV94qXYa2s60lWoPmglQtVX
CfbLx+4pDi/KM/PyOXKHm3cUfXHReqJ7vPT+sbXwpQ8V7yhe0KYEQVtiwM1Xu/KQbg6zdGeYDF2c
ESU4WBOR4Fk3Tu3IogWcHVxMeIADx6VC8nGvJWpah5q0B0na4ACFRqCrryvseWK4PnYLP5NSiWL3
WEjA89i0i3GPEAXm80fhHSs0T/mf1Kwc/fPeZrjDIOEzgnK1mqoKHIb1SpEBJtZPexvF6vvH3uSQ
bPtb2pgSDay95JW07WFYZSxzROoU83zm6+RIeD3UCviMzuit8nh1/9QHD2eHdrnYi8T+k0miWrKe
Qwr7GXKm/zzwPI2SBSnKmjva6i6JUZB+mnyTHWdra1cx2Iyxp/rG2krua6wQX9DP/UQb6xCv1OVQ
uxazdXVd4185wWXJPwMxrN+ehw9tqTA9E1VpwZUvYHHUSGEK51H0zOyi3bLu9vGAlIY+dfVyUqk2
hd8OO2D6p0I7eDjkZU55YHFQl/FUboSY5lLoi212EqosmbOrJo/9JZBGrNrtQ5p7NpFvHaZLY+Dy
qh38S3FF8g5c0uYHtQ9evMAEIzcFGS0qg5/C+7I4PH6VsvpZTvsTeOfELreNBN7MUV8KgKsgUf4j
5e9uP/oEIn/T9ZpTV7ckqcy1YTgvApc7MUttvGWmXq0VyCk4UEtJi4/smX2dE4+cB2uv/j3Wa+Ja
lnIFTgZt6mPfbRMiNzr7/8szyZCFtkbb/11HVRnuCES2JmaFaDG9FH+TBQ8eupf6oakwe6bhYaXg
iEm6ogavIrHT3PRznCpAphQttSRaJLVU0sIxegNCl8r7dsIkgzmTDZMlrpBvG6cj1XEHo59Abdpf
/6TBgOSD2ceuveVyF8EQknnoTKOOs2mUQRJvChiTIMvp5lJ84qisJAy7LYQrxy8c2DhEEoccX7aD
NiPes+ei3qYmP3DTi4nfiG2USTZHeL3RnZXBz6gt2zx34FPC2h1O41Duwjuu2X/bvgiTbS3bz+a3
5ucuSXGp3OmFByx9+1eoZglgoD2s6ZgdN2+c2syiWtpeIrl5Sh6aI235+wfOSO3SlQMx92WdVhr4
C55r9zeIGL8Jp/Xy5sdvqLnZUZ737rrH6I1OO8ZJEU7jn72nSfvZTnc99z+t45dGaOu+9jNW6WrU
mn9oSwub2iGBLxJmSbTyHgoyUyJUqebhp+zXSYR/MMGfOIls7eSg8aLlszfVyF4PsY/2UI8+olDc
CJeyLnwRjSqW8QRb8MmqZEmLr/e7MLFerDABItyZruUcYEKJTBRDumBMMchZCsmW/8dwUJhUB1cU
oLiVXg42lr+cvij1SvE7KQg8bbbLjB3O7YtoOFTFS+xxmsfG5hdTOpf+gzsQcjZMp8DqcYg1MnbU
lYSsSt7W+gxvoEGlDkrKaP4Ezjlv0EawBOCYvb6kGOKk2Aq/jOezvhDfQPxiX5fJtpWdsodd5+kl
G4KjVh4Fkkanv6Jn2Plwzop/sYg0HiJ2DV9DZBXjtGg5sPRRAxVlXAtgIC8xeEQxuMukNOEItAOe
8O/Uw16YomiahI0TOleEuaunOSUgCpYeuzbHArojfjXpWWlLWObNPb4dZ78wA9fW4JA65EocIPzA
xRNaGo5f0xXoCqH5WMmQD4s66Me+54ga/RrcVF+rj9UQo5iAQadJxLEHi8PxzgIpmKeYPqEtkSLK
b8WlbR9hRahx7keurufCo4WAqEZcvwSdQE/IKgQ0ofzc4giqOw0jjljXoqT/KNFQrAHww8X153Dk
+mfS6Pv0jopGDSEyxlG9XyifyJJpBqujVt9/Y1bHSV3/AumcJ6f6rgzwhH/bWtQ17UN36gQJSE2l
qp6AzfKbJseQTRaukkH4daswhVnp4yXDFeDq3a+pC4OkR+iuualvHP3m7Zy1UYHeRQFXrmakxNcP
bXjKBTUi58CxXs2YLkCl8VLWKRXhgHFORlZl7GOt1lzxl4hvwD1loFx8rzKv0N7e2liY0dkot+c1
I1BwmtHdHKky1BxdreZ7CpGvTpKwR7zYPtFnONBrTUFy4AjIfZn3PpXfEFqnPQXKonAfJwpzpoFy
q6o+SbxAhnU8xDMkqWKhbhq1eGmufAO1ZxfC3xTLPVN6wFP2+NUT/stbXJ8ZtQQ+35rA6jyUUTo0
Q58BqcOam9UaxNoWgZArzVXk5qFMq9kO9oOAydNoLUT179BEg4lNP0M/XbjcAgkKT0qNQJS1nCDg
130zcnIUdLbn6iP4eBfOwhpXmi1C+j5ldkvCkcCbv/WJF/cKkIsKkXApN7kOR2sQQXC6cQlwd7qd
juPLh6u+p8qrWsqW8iJQgqYBJecGXj1Mt8EFeNaDvnFmgjHQc68+DQkS6tJcJL2Wg4UQMc8oHgTL
kOVSR+xayqVCxZYzMnIzgY6C/EJ7aqHtgqpEFUNk/sU3wT0TptopRfdrUTsOvmYWjzPtOS8tsocQ
dznBa5AtVTjJRQp1abfe2b08xGISAzP5tHuI4PUwngHkYV6w6cdtKRj3R/N/5xQeZDedFQyskECC
KurcxLvya5+GQ4iqfHTOAeLUMto2yKDp09UsfHzXsa+30HyyNaARrlZ4SiQ9jwyI0KvzxV+x3GsM
ct8PwR5iJ2jYs08qYWpQYrUczQ2gTAiLe4XHrO4O37KtbPIlj0H9he20PDGkCgDGO48twadwC7Sl
tVPNMHy9taD2EcM4uPAhDfCAH8Y1c346ucMCDcqnGbBc7orIQjAVsGistoCMUUiB+AE64GBsQ8o6
QnC7utim1TDV56GVJf20ciUE3msC0KMU1haYpjUVgwcJ4zxaCNERuQZ/QwcK9p+0AzdqN+v7rfWK
EjYiWTxnSWwwWEcudoqsxRYBUoRI18m6dRL9n0E8dDmGaTLju6kY11joYIdO5zzd/9QroGJxB5oW
5So5iSRkvp3NqQKzPAU7F8KhQnNZAoHf4S3EeFuf2wkkZefAjgXqwGTl39DL0z6QBKMZ9PZEMcC5
lI2GfApwj/bpDWRzsFrBI3afaZBzxWi1DD1pfOwNvpMTlwhnqo62yq65TydR1oNtzbwKqAOmDbNB
/lE0z6x79GNHPbpC3sP//FRNF9VLAFuPdS2mm7MlxQgh3gocFuyBh1yl4vqrpfsfgGT654Lx1Anr
u7Dt48u9q8gqo4KJ8kY8Qzd+raTa7LMDKqbBRhPvY7agjP9KjDjpMwW2O77HvXoapJUrouH+027y
QrUZ0LzGDnd3XDvI1Hxk/5JHbsVVPeHx2Fe+zI8Z0JfOfeHS7d6l1aA03aotWqB7gWjYIb/uLaIb
aTjjoQQaYLPv/LndF6GjNEXMIgddKiYr5BC8loYnntYSHVOlVrZM9zBvfw61thNzqRxMc+N3FDjo
AcDxfGHBH/F77VARo9Cz0TXnfRSRVZklFEFlN2HvwCswBA7r87EPf26mb09iMuzdwx2oD6hCOccs
Vh9z3yPCffLp5AVjgKv/NCAhPXZNtQoYOwLn28Z+bPBZmVnLlbMVTuETeZhjY/G+TxOQhM8rWpBZ
NfOzxw6xO6WkreY0KrU723aNecT1F8a8MxVmacgtupWN0w2Ulhdtq3QzKqUz8AwQ5WK/tLfC7ovr
9TzOEYs0CaxCnAcUOOCZqZGzEq9xECxMRH0VTWkzGlS2PADTJwxILn8Nbi6XzHYUGdHG0I3wsygo
YRYHvvTxkmE0j6lsGbItXYCixXPJFrVdpuGNTmc/vrHCvGwcDhoWJeopsYONgo2cqX1LOYQsDC9w
cafo5aWmOMLwLj4XF/U4cFwBsUfKLan3U71u8iSagfvo+TeB0hP7Xp3EwBil6kJSNGOHGwQ1M0mm
DJYBVqpjsopj4p3Bs8NmcVpQZBDInlNsymIdRMCBEZcQGYUmgIgpLyA0dbRzEXUz6cq4rPWRMWTc
EIKezBL/CW0XjZnurdrfGO+GsuxZMPkhVz2oKbCV7y5nFwtlaK7hBQeu/ac3gR8d06R4dDVSKsvT
hKBj1sdNv4sgWHnQtvmskVeW02gCGu5nMCphL5ItHtsMgkumrgmqiPjjDv32YyvIESgcypoq8Fyv
lSSlUzBVhMVCYvGls5wzeXakMTXVwWPeemY9SBvTLkmCRVzxUT5mZaQ1tsNohEwEhSAMm47xm0n+
YEWzj5KKDR5NcSFxwGnBX42WYoJctYtoI/hcEgyAF/e/lrtC34C5purH7hHlJZyHIaqYRecRsv3O
JJe1763qHSmE2bol7u6ovUzAMhMUHW9o1rX+fqEUWJCZiNTyQkjmimvYJtLq9/+1zO5cc5TgzdQJ
/elECXbAKqif1Lcth4xX+8ONAlTjFrqT/bhFOJuYR9fm9J+Id3QdCIpQt5fDkUee0tq6a8DbG8B6
P3ast1DS9S0zEAUij+0CmZI6BmnA6VnZFg4Jw07NXcpLeVpMX3rlRhGY+r5bC470TsZDmSabLmue
sXZx+EmM8anbrGaX9sZUgkvJahv4Qau3Vg+hwvyXoqhASFHRDai73CPwSTgru9D2GJrti+a4LoaE
r0TVm1rJ7tPPVRLldHdABhqMICZwbtgORAizVwzaY4R6RYHx9rhViunHYl1Bcm1IDxZzn9nwcvqy
LxwWkIond7N0fHXZCCMyvWEEu+yxgYZTKgcdw69g8WBFh9cLTY4wZiifQCMjUdMlMhG8Sh7KpikT
3DMJ6R1Cho00oSV0FTcfWz6SeQdVHrWeQwxpqc8eOqI9ar+dsyzCuK0oV8vPWkW0e97onKOoJ7b2
pQQHD30qHTsehmG5GQP3jTV1uZReyCPX8VxPB76AJ+7WlJGdumOCgAKQUthGj2sCKzryXJSe088n
S6hsORSCsfzJDumq1SHuQheVgu9SJDhe1HPDv0LMX1YdIpob2gEKvgRfLIlmlvrU+/IaTPRD+c+z
/Rgi+XIrXQYJHU82Jp4wPe7pGkR9MYwCJAwdQVjW04E8a5X/1zTuEU+y8hgl2dlEVLX2/txZxnpT
AalmqmmPzVUNKOhPJU77irLmKDWpPB07ygnPogHqDTlDYi1CO5y/JtEwDQCUjpJYBkZo8GdCvv1r
V+YpeXUmtNnKMj5trwd2TA9+hOmlOWtaWpJCIPVm7Ughg9wVzgYg9hgPQ4kIffzKzxQc+rSohCHR
KBnht/f48cXRZIk0TFOMyI8lnv+peA42NZKBWQt90icZacb0icy9gy3lGsAz5JXuN/9kHF3lPRjt
i4IKivRF/LJzsX5uGGWNZ6aE/s7YehcZu9iejFEumlZ5oQt5NzsscZg6I8QzUmmMDR6B4lVn5ns7
AcE/oHGS2DyStTYKH5WljW1EEh3sEOMeKLOUcpZAzDNg/NIJ2dt3V+zRjMoHn94jJrquHK5+ZPt0
EEKr9kYdq9xqbm+SVnyyQEmouv6zzs0bMtkcxB6sWkWknaq6j5DZlTtYW7QyFZHAjl1mBZC+HZqX
tFZ/Y87rH8LtS/2sAvLhllGZDJedlkHiqIuCHRdRm0wvSXVue7p/+wVU1lw5qttjt4CaXZMqbrLW
NZkMOa8q4z8F7VMotxYi/1Z6KQbzN8UFUDVlzWs4zXL0m58wgd86vtX/oVyYYtGpysZXCTQHQNEu
07IleVPDRxH7kZwaeaqG0++5vj6TGdXtKob2+2d2BwB1LbPISP1lDc5wMapYdbg5C72T1py6UGKE
STNXYGL4g4OqWYpZ2RzcGFv3Rr0PioY069pu5VMl6SA6GBowojNFwMc9PWW1utn4jW3bRR8Ci4kM
CjT6hp7LrMxefWRbhWsMAT2mXwqYcNNnbFiq4xqcWM0BgJXND+bMYjxe6QM4pbvlCCyJsrOFxNpR
6QsrNdD50RCOigig6R5xlYV8KOjfhBIu4zz05M6GcojyG/V4VrCEJL716xMcaf/uA0b4rhb0Jyrl
1sjMVv5IyjxXgxbSmSCuhG7sa2LmZiQzL6MwPGcDRr00BC/HTT09M4+ztAKyo56Xd/4LIxbrZ7s+
+5RVf4h33GCPaRy9GXL6GwkZUAsz86VVVlMn4B4+Uj5sZTZ2QjnmYEcWkdjCUo/c+UoSKZ0D4Px+
ecjf4BYufQWi3gRfNSdemtBh2RxNl9mocF6UdVvTlvxlLjE/PJREfmHP7E8WZdM/H3cBK6n5LfrN
J/kMEdTn7DSQjDhR2TpUj7/ndmJ2SZOoWFppvSjMTKWoeJ0QrlHkktu8hu/AFbbhprV1AZfZxcFu
sv+2QIDOkXTiDTpIh+9ThtkP8YgljoLpMu1BMiAjwKQCEYmsdmEQdPJIA+yWhLsFIklLY4akKHxp
DRiQWZYKC7wSpGUDJuZ3aK3E6s+r2xBKuzd/oXYLjkIeb8AAByF4S8vZ78yJaI3r8ic4sWZqhwm7
o6rElt7zm5QOpAZCuyA3IU/L+nGWzD0u07+QLHAXCON9KI0QN8VpTyWoDbFcDGJI//i+jUgIMUnP
IvulFWsGzTn3P9x4qIYubo3cmgqWkz2wQ01bosf9iFhFz/CFsrutex4JY8yuRzC6pWn7/ei9Gu81
4QDPC+RXqavCqdAdkQRsZ2kfZrcnrDezmMN08LnHR8twnxujlqbIZou5+qnndHtRY1xzQQVfpi+J
1m2fDbB8888ltttC8L1ICLCuRena8TErEzyvm2ZLj9Rv9dHQZvdOsIvfyxDmnXXbY7h98bFBcqDs
WtMD9chDSmlVTKJkZBKM5rS4NqBy72fJR/T6BAVl9WJn/aDAIwM5o5nRm+g2mQanwHAelUaXWJI7
FFN6Vq3bu+AEPBIGk6ellkDlk7hMCmAwUDKZxXYzvQmF7PfsqxxYzhF3Ju3KdVgMqdJ1FYKILE/K
QA+gb2JAO8NnLjU1jeFMBxe6BMC7dL3/7NWNRn7n1F2v4ucXEHdvn4zQwylWphwno8I02kf3uNDC
TnVVAzlFBOtRU/gRgsYJAZ/Gh2OayvnrDFiflTRvzCTsJzFiixIAzY6An/LQ5o/0tX9l4EEEEg5Y
ZM8Wg5FWVEeXDKIvcRuoO65+1YRo6Cvos9bMAW99HEaR0tX99z90as4XIEiqzJHzVWUvJVVpyd0k
rFT40Bysgb4pwg1Llb2VI7csbNDWmYGJhsHePgZY8JNOkVegOrYmZ1Un3yEbq0a1fot/Nh9O7Lvt
+XcqQReGOV7AOwOUX1+y4FVi5fEGX7dr8fRKGp5+IYVfYPx2T6W6q8CzhXcD2meAIJZVSkFEDZqy
KPZ1cKtsrrAB5KIbJuoYKljm4Y4EGSfaLGK78KiwS1DoBnBRRAZEVD46d6Vy5Yh4vBo4LccDg/R5
G9fBN/3INkdI/SCt07zBJibKWf/tJZXidXH7YPZQhf4nGeWI0uHHxTytgRV+DNcwlq4QzK3+pOtR
ZM5r1iBFDD+tGDq6ZLjidcySSTrVsVAOrDpsvMnOIL8boANqWKbPXgYAA1RwMSdU7mnjDkaq4aT8
s5xFIqmIQ6lo9yyRzpHJGJE3C/LQw00sUirCuipAQtHOthINuVeviZRKwUPLuWnv0CuWvnxtLGba
q9/HkGjOunaNy0xseblYCVAK3KaJs4BqzfAAbNDTLZnhkaq6FDSHreRgRDeaHHd4nde/ksUvJnM4
WStsXYbopfknj07frWBM/XwhKkAaPj9ZgzgQ6EHCu/F0tPzr1yjB+HGt6yRv5wSyQgIhfnAwVU8e
gj4kFN+rirCZCuhDCZ3mbCWCkH6LB/FlGrQ2D6AXnyhJFoVZ1UTFxEiySu9qTPgT5DULGJvwJE0p
9ypAhY646rcqEndgERMeajJTOrwu4/zWf/zoCB3aIUuUGVQ/PMVXvq8N8H0+jIrrBYinUgaN+0/0
eHYML7nTmXH/1f24qOX8Uk7r9dYQId0OYGau+BZqr6NfVdT9AQExffwmpU2gpQ/kRhkxovYlqI40
51Ii/mPC5gDI6fS2ny1f5gqkrtLkTQNhgeRomnWb0Q29iYa0TTiIsGA6VPCyvifDkfGo8cDLxME7
BpGXZLCdblBg+m5oMnWuvMC5OMAJKjGGGdn98VKkdzYfdTxXhoTjwr0bbo4/DLAZ6yUz5Vw4V+Ww
JNYc7uOVYp249kg/P4CYcOhhHIlpDRbM/CdWL/kuFFbfvopZCDMyFXYPWXXlPUl9LPHMOGUFOPmJ
s6HG7csfIVUx6zSGZANHDbv6KpSq37zICVxBbQN1qIYDcFr4MMmKfnCK8YboGmg12kRYkW+ShNen
2pba5V9NIhOMwzPbpJHla2fh4gMRBaKqEQ9qWcjUBCfm/CEWaf7FCctmLEBt7p6iPR13061Ms17X
Fe2SH/s2Smd+AptyIa2EHIyESCq8FLEUoyc2BZsBlgtzntujzp5onA2P0ZW8e4ki6v5S5hctovwm
uOkvNJlvoC8nMZC/mZPPaLnaOy3VTgVdqK79vHWspxq8fqFFKc3T0QxNXw1NJbIw2nIw5Ju6Jnxi
SqKLbdmwfG8w0WYTrybUbk1vYS2DKl5R1JYi+biPXMWvPFL2TWI8Ii1thg25dHcydVP07vwYHvCQ
q4fKtfk3QNY8qi37p/S+gWTsxN0T26fAi3xOvtnRcuIVYwCaZjk2A65oArHsqGUa+5kLtRQgVuIm
1xEGHQoAgQ+MQVA9Ca3IzMRYrv7ah0le6ZXCsr15jdmg4aa7K8kmtZNhpc4AjBx9sRpkw3HKT0Au
XuBPWF4PkX6IjFj3ORjFrU6A71jqsk6BYTfxzeJirQzI7+1qv5KLSzt1fyL+widxDZW5fcoFVCU5
SxS58VGRwSp/DVirCvVIgNfdupfODmvnncchLsSfxAdpwlTasZ7lsZmWPXLmt+U+OBUP43ezEIOM
3a0sgxfDHIN8YiV6B5wPxoXnKfUcepRIl+AHAIGeNt/Px4m7SAkKCmwrcRsiwqPW9qZaebpGZLqS
PVIXmxRoVsQkRss9on9AM9tRwah5/FhJQZeaUXZorWjDzIpooPe0UojJQPZPWCkF6j0WR7RLoyAd
u6J0fIRxB+J6jVOHsHFgGoQX+mNb09XTk5jK7oDVIsgxSLPB98qraVJCgnDhHbeJiMfw++HElXr/
7r7hFGaK1A2IzVfLH5oE1gS3fkiRN/fSB1QwX6O/1GfYXWX1gPPq36nvB1OkQ8iC2LB/kgtOfVGK
4xJnbvwVrgfBw/ryrvT8eqzLSuGQI5uimLVc1VWMJN+TDZPqTdyRQjLwoWlWmIEs4yLr29bHdELk
wAn41bfdCgykmN5KkHK6+sgc6Ry4qD4kJvC1JgJxd4CW7JWjy36tCnLHkuxwcvPsV9CLBZSXI1/x
Q9Ewx3I9JDfJYjlhOgEVvnhfiP3FmXAITp3PriweT8WDV2xRLAyuoWGyBjJEnzKpdPbgz99Sxvjj
u9rRw0I4w7ys9DOVc8dw0hiBW7ByCka5yJEzIysJVA4fBbS24W0d1st0hOJhxicq30kPufFTNnky
UgyvL3X6FzlP9DhfTUzvF/6E4BwoTqM07yqr7VXfQzL80+GPVv/lTIfKtcRzaFVunRCvjOVPqlgE
vvFmapyhpwIHj/wmOGr8HiN01pUSHNLTtejsQBSEawuVx8LFDrcRWET5aXgHE7PVrLNISwSIF6IH
LgL4EnEqCNWqCp1TbNQ3SK++AdkjPre5WNPys1r9dj6DcZF44bU3Nxnjt4CAhJlXgdeu4QWt9Ycb
R9vgZjxDvBqRJvyWFrpurr/E8rmyVW8n2O5sZpB0KsQGTWzJp9dI0ILIGKfav+jsGQ+4hGJ5tRNP
FnbGpB0ADhvzVa/C8bV1eMlzTY58w0PAagmpEo1N+oqrxjyfCt5y/sYqikFef7JT3bLD+mp8iCTG
Tzv/FbbXNCetsfvoO/icC25hAKdqJkRiGqfzd6PK3pv4aJxYQdSWe0N1C/xGpfz976xLJOjef4GR
B6H4f3Z7ryFE7zn6pY/+I5CzeOnF4KDL1Vcmr1A2sAS4dsQgSWNc/DGz6F/Ieq1DcTJdiujjT4mn
ayCVAn05j2o2VSo4tDheqI53FIQ7zQVAvsTQ0/d/kQpbwssCNDp91HWw3m1BpsvJsNQYsHVX+/ye
gnEI27clrivRcrKuvPTWmpGxvNcJcupihjNr4BHLF15GUx0l6IWyPNMqIAsEyD5gd2p4S/vv3ZT8
eBgUI1nrTBeFQjopMIJGOowiB4eKw5lcyJAuvJZ+ycRo9HS0VZ/AF8Gvie5F5Evu7jCOoPYUoKUt
xnwTJLbn/eeJE9/4lzxtsJRoqVIiBoXXJeMs51ZgVWIwTDeQZFsUC7WPshHpwjEfXYHITSNGSgzG
gSBro+kh+Yg6/4SaAkmwtWGuBPOHAiQhsdSgg1P/71kEwJx53QIOcyYkXE5u3H1kA47WZUjidM2S
aWRbWVECUaU9GsASOpbx9MuPoHp8vvZV97XkTuVMsDJz9fkBfPDtMTbbd86au4m6iEEHKyN79nW9
r0srO0t2I6XodIqCgeYTZAINRSdgVBBxrJ70udKLk6AJqd4y177hcsXVpgmfwj+EOtycv41GMYJO
PoH2+8RykDgGY+Szpr6LC755wuVGTbrokFnqdEIB+wgTw/5gDBh381ROPLq9qmTkW1GFdxsiapmc
+2UsbOmBq7XHdsQnFHzYdqW7ACUrcJqueOmdY3GGjAIF1KCJce3L2jPHhfJJ30NRXRx34YLf+6Ga
iwXvNwV+dQi/P9WspoGE6iEnbSIa+HdVD7qEiOPfOeGvBYshQSoeulxA7Li6sijbnvCc+C6EcAAs
3nrfAnAIwFHF1HCdbAx+SK4hbNQvJNVlzpj3CCzWeFXJTQ/n7+VhKXzgYhhVAJ6f/HQeEAbwa16L
kbZsFme4AcmV783Wee2VVP8eveHGuoxJ1pKo49SkLIu98rXkPEVMkqbqJNyyoOt4YKcO7NVI4stz
2aZ0ccvPdwLoS+UvzBfF4kTZymyG2B+AoAqa/dT4555msl/GUXdiiuFIVco+3+FH6FFdjCoE1Bk3
Wy/e+mvFwmO2wkktS8qAGCEFQCf4u34IaUwqzsd++hY3BUSXjuO7whOTaqklMymbBep+HIHR/y8x
3Ux6WsgO1ijqUBiNReDAMVmNop1rvhWnCj/vZU9bFWWbtC0A1nhY/zIdY9UbIJjW1K1WBIQDTUo6
3MRF7+XcSH33CVX6P9uSp9ONDRzJ+9yQ26UEk6az6Z8D3dMmnrWCkYynuG0wgt6gUri+SqYZAUKP
pDBZJ2Zi05Hho6LOBhrym3Y1zTLcF2/qeiRlOtE+qEEgpKJydVhSyx4qmu2s143NGL7TYaq4llI9
CcWH51PidJz6j2jH4feOT5FLFQqKIFYuMzwjXH5dMa5hZ+/d6WLa69MI9MPNV733c7f+0gXc1VeF
92np3eVhvcC4g+YEK5k2UqqBr9NireeL8xQJ8PGM6cgFgpT+H4ghbMsxGxtFg33dSX4+g1rLI7ub
pZItGDGHgE9fPsDatJgcvrox2O9oDW12dnmOvZiqsJLQ3+esAMYGlItRtLJFClVgGaHiJAu8ioWf
1CbmuzIHIGotOB9C874L35oG6b+CgdFhgpOulbM7tb5HDd9QbTKO/GT/wwF3T4UDtUAb6TqH3sa3
uzuS9xcDDtEd2kUrkap/kBXA4nVluOHdtn8Jd6Q3Fs1KjCXrM4iDZ3uqbhrS2P0y/PiScabvEW53
yDm+1dYq48YCz0AouFdShJqoanBeBXyzHU4ioMBXcFApbPcrykJ39XSuEnvH+AzgcJtmUkeL8iUW
ccqWOzvTR7MdyJAbo6pahEjNcSFfVT3IfJId5GtF1FSKy4A1lD7kvBZ8rrAoqQ6vXwkkanb8k5HG
g2tnqlF27mZC1n07yj9wzuynhPPIEUCWUEe//MCYrP8h6vmwIfkY4+ZTXUiO35wgd4QB2mbzs5Zy
a0ca5seTBFkQFRNgVZgzc0YOgl4aqZT4HB81rdpqJZFOalOHv9Sov4z0vP/iolFAlXhUsEurOaov
hqaMWVKJMlvQNT+2LD3RLVUP1v8ASQ2J43S6f4P9TKuur/AEmHPyrZ8ijFW0/lsIOpJ54wU9/3RN
3gGYkjvs9nkeb9e1sa14tXyiXgYK9PWjt94JsGbg/2anoYoV5EI0i3euJNrZg9sSUDsCe9FB7lYG
YhOsOxfw+XZHqcxPfkAGIZ6C670MVyKHRr0Eyh7dolT1nfGja1xkFHEwz+YDxsJc7kHEUImK36HR
5PHvM9KgFtcVA9iOdKw0xLkzRxBwMNmqplCnjvVIFQ2Kt660gBmm+cifrGg1Qx06e+QmASiWeQ94
ed9yJv3lqyuAjlLkc1NLQ1J+F5OPUG39D/TJqFW7aBqElPXR/eFyCSoYJW6W8KjeHkSjx/uqb6Zw
iEZzmL4ffRN3Fy7v4k+CyZVcSTor+gWSEm2dUEksbU6cT5dmtIKofZd6datWQGt8NhK3l+RPyj7G
5Ql8CEbkvyPH7apH4PGkaDDPfwY1VT4R/S9vbG2TUSidrncDo8OUVQWUFkpzGiC8rWdh8X+NbEhf
BVundo8uE4/sMf2/0qJetsulCmP0ogxWcZWsaOtPoGVSfM12GzhETFI2+V1fo/rNHCUU/Y1oJpWk
BKOUXHsZt3YSFgoPL+Ifx+nWOuTPEdRuWzsvzNEu8N/VZRh1j8HhkRvC9pV/sQ1evAWGFExppWbB
mhK+jubs0KPDeYH5YMIGYEUcLlNgV34ThWRGCXi5PghpjIa3/9GK+6hfQY7eaizsHyfHC76XfoSz
v3IumoOLE4CFDnT8QeBWayJxAfHky5rFHkMXP7aGbM4zvGYHSG5VJeYsPWxtK+LmOwJ6qQhr/QmM
W+Z3N/RsaJ2h+SE+GQ/iNUTUdDcIW5JTpHUKsnLm71eHMjAkNiL1lH/7OMONcu2zJVrKgYJ222Y7
aGSiYY7AviFeTj1eDRMdyKLsQ68SZ1earW9b2nW6XsrjCSFmNmnMjndWsnng2dIUNFYCzVH4BEj+
nZ12KDdDvxTIL0Jtjr7W3i2rWSyBq0Z4OfRJEi+oerrUHo0fTomFqO99R9VzeC9qysxR72ZikrHC
GStyNQbVuC8aUoEvrX7c82JzYuDcMEpbYflVPvX3ZpDvPpi86eWSOq6b+EBc/27Lc7Y+B546d/PW
Ae8EtaDjzEi3/kjsZOwuUzPxJbssz01Kd9xgPNOOvoMfD9bpPrN0U88rK1n7M+4ZNcwW7GgYK84p
zdg1uWXVVCimpLodbSJsWMfwYgFCQCtufNRl1MLRbrIw8GHlpaYqmxTZOf7EFQEh/Rc/FCKeQgmz
6mBsZ6EDgqbaYjcXeTNXEdBQXviPP928jXL462g+7SLy9dKNwr5IR+/lEOtWTClz05jBaJKn0dSn
QHo3tEKukZ3ZVDdDLy72MDWcZTak7llSwSyFOSi4cbKOkezH3isyji+lHkdmn3DVAVTXLrUFRgSs
o7ppdZOXAQkOb8fAHTiimncwHCDju5u0Keybn0uRoo3hyrXAlYaL3LVzlxO1ZRNOwX3iOmZB6gvU
xoTWhGBBfMjLOY66njgnZ7s0hONcwZj1ysjXnI1rs8R4zG8AY0Y8QiaNPYkOGB1GjWoNjzWAUTw/
n9gIUMEMH/XEqbgX/FIgfYfD/LCO++/gi5X1eSttBz8fEaTSaY4DTqCyiWQ2+t3fc3fez10v6iw3
yoPGHkhnqlDUASC7v/YZa4B8h4xIJk66ToVqGUzIrH6krkiRv/sk+8Ltz93Jn6iIkm9ARZZSHD+Q
crqYDdUjHO51myrsbkQO/4Wy2iya1I7NhSC3cVz9Br/gx2gS6ThuP+/ufs2oyaormOlXGkI8UJtT
zRuNTfdBEhuIz6xQrpnHQWme54qR0+V1zBsdLr3uB+0aJai9WmqQCUZT4pYLMi6jyKs6WGIDSFk1
VlGgyvAXxXY0p19dM74QNFYE0CPUpfrLCek3+IXy8RiYDytvWWt1mJukdVJw5vplvY5DDkImjGy5
LA36gd46kkoIwD+Jc97x1EqbV+gdpIdMzo0596o6Vk82F8vp5yxPTVALwgoVkaYluJO/UrSZsJsu
6OW9C53ol1D3lTnmf51ZNZAZN6x4RG3088Ib0Co2/sXhwjnHSykQrg9HclvotEmpCdHw7aaWEeDk
4sVkU/6RiM7TNAWY0SNO1KH5um+olWSXWpelN2GnHWg/T+kfxfmUasSrMKvYe4+t6q56M8RQnvXx
GZiZ6RjwLpXdlRP0C71Rj39r5te81um9CaTEwb6IQz+LBpYu66GUKsyftz4jVtFt3gZfVVfyPyoV
t+K6VJUQ8vjGP4Q4ZyP9QSqdEacdrvRBWsct3M2aG+XYMCd2mbgNa5ZXI5J5Gz6nslCHA74/44Uc
0vTwhOiqwQojVtbXBls0Z58G76CMJN9blnGYVRMWTrR0/z/VGMdJ2Tlk7A6kNo+CcS2oExjZyG3r
67JNZYM+9yc5jrRZHF/KX7SGgg9itJkQCpDZQhel63ORke16qRMGgxveu0vmBQj6LvtAb8FZM+aB
ap64ovL4EU6OIgq1ud/pJ14z72FZfrjjcEyYxXmP/FpAgMLtY0q9EfCoMSXG7X6IaSyINbiB+d8i
j8TKVFp9z2ouWUuUf759Bg/u6tCC+IUjSKizIjQZe57TpJiFS4GkEL2NW25MDaMiV3QORD/iyqk6
z5bIB8oFt7hEHMKu2JnkaONT5rhfbgdoV+p9738g6w4XuxQqxuQNJW17fv4vzkDe+nM3KgKznyuG
/1biIvvHilDGocNyYLpA990u3gHOc6VpsS6hGTFUjP39At3JQ/GZg8bwYKpjfK1PsFsmi4S+WuiV
J8N2JJIHU7kqscJxktJdUjpcaAan35ge+qhvB4Pww63kdceq8z9Mp0e629iFh2dapbZYruD4XrdY
K3yCjEvLkh2GG84p8qqUXdcZYIF9GXN6vAA7ZrdMWNq1t6c7v/vK66412eryZFiQf1Wdm+alv5Wi
IukbitzGnglgCGLvj9AUG/YvXobwd/RrJmh2XzLbtBmGUN0Jr04n8Jsjl7baSdlyvw6FQcT65kjt
kUM344ptuUv4spuo3va+szG+gPM3NOqtkEjgoAqXpz4p+vY9AwLaVNYYW9OvNLnLcOrw7Q+jf3hf
HAG5UU7ev9y3Ss/A5R2AoOnMYjk0/hmPc3tUytizdXO9wwatlz/9vR8iTzwdaIbmnQlcEwCYR4AN
qj+QRziAjzIXBniIKJQq5eHcoSOMiSQDG9veNbNu3H1LP/DF/kc5VQcpGMaZr5yD+q1zGFhvze3W
BYfflxHyqmkPF7ofSGckveUekBW5SuFba8QiKxLfO33nveY6s1yjL4gVwcI06+SL/62GQO/hB5n5
7me6qwZp6EJKpQGkdOY8mYFPk3+PCwtkqZ93wiyebiVIMFNEPKdXzwIycPoMD8QV5KiUyy5CFqiC
iiFxAQC8hUjLJ+WALTWZR3++OTQ1Jae9VMyFIUv2QrQvjieq+rG5nJWr2ZfYFUer0O7TuMD2yrmD
JHDbAPs4i+vAkJCSnhwTszS4hPg1+uy1fP6/ZnsAamhKcm0W1pdcwu4mnP5QxTobuNLsFpCqY3rS
zSSmM2PS+h6KFpZIE1VGXzGQSCEiX7EUcm6p3z7+GmWhGJaGMen7+nRAWFcw3+QWDbMTATJ6YFZA
ez5TzfEtDRDZ8N+O6aNAjtaqILxFJtPDuiUvpxEzFaFZSvH/w105T9FxoSU3C/1CKOrQjEJlOKUX
4LEzjEFeJdnNi73eKbzsotzOMN++Te1V3DOjmJkXKrwqwtKzs+iaxkzFUw/Tf6WH5DTIVmc5BE/H
Yi5Q7Su8hf1gxzzZbuRVUDr+XnONDtu3vvOjGbKWy0F0a4x3Bt+vbD8H6v28XurTTFBctjznsc9c
gXTRvXHVmLv6nZPuWCftUc4xip4ZNgPFrktmVVBRxHy9txfYuxmxutrmXkJTKfiIq/jMAAjrzMd/
ga7dRok4saQYYOJ3cNoGY9K1PzJlAdx/KQABuXIpoBF/1cKzIYxNBh+7fyvF2Tf/CYA3lP47I8fb
EtFrRyXjqYZRvHtlV+6mNHnSnFSml54UBqtXQ3+hUkKNtYc4WC/uOk3Nn80u6xnBh2UIpWdKXHWf
xmkme397FZ4L66NCAfr9EAWi43AkEdWGRra4bZEheisFoHl3QLp+nRlrEM6yhDReUBF/lXfi2leC
fvwofYGt/tpW5zrak2IKcLUVARalw7cYbsgMMq2oiHm0RTT9vo+DfYmPGv4btgNs4GwuLW7RHMDl
CgXA+rxwWZhkuFKJ/9YmZ29SMTsUtIqYORNPt4xMFY0UeTRDO7bbq2IC3dxIRFB3wvXmIXDprav4
6QHMJ0AItYG/so6D4d0Pa5rwKMiij+t5EXWRNJQzv0zaas8JY7IYYq5ts+fiTXBvQAafKNeO7fcz
p+P0/4S22Oewe2Km1++kVOkmCqC2gLIzJzhONazvBBZBUCnCvR1BJQp40FqJaAy3Gi5qjBcoOoHF
QI2N2GoMtj4FX9lhb6BDJ+i3mVT/v2QSUwwQjarZ6hg+FenJmplo12YCiJ9Z4V5FtBN3KmOfowpg
hhPJkjZI926sA56rSofrFdwzumzjNRlNc8+9PuzMWUEdoaBD2zm00CW6lCrKpfpDo9jLgbHBNIpF
pQhyiCGyGbcadvAde43YvNTBljbS3NOlKhkG165KjA/W+EJR3cI2Na3U8j5cQRdVrsOIMuKVDD7v
lDDgr/aPQQjcfUGPCWRN0aQjLSozaaxi7JUi7F9IXLLujoY140oRVGMcJlNTus81Pnzme+TYt/BO
vjFgd5wQ/oOBxqYXN0e3TihCFS7beHQzcLi+ZG9uJqkUpj8I9uLNct7kRBH9qtMfRZDoFz4vIElt
muQJJ3D/L+SInBPasAI+ulN7KZlTzDKAGCz/tiinVVSL0n4omGV0GQ6dNKmV7BThWxfY4nP0o+RP
7fxjfztaz+tX2H4yMrliRd3WHo/gU9XW3y59mC4puqiQs8qzk7Rd5gbHbOYHU7847415OXsTIYte
/p+bn10Wwd+qHIyquICpy/SaSRSE99NeiyxPOYATOLZ3M5acRrvMosEEXs17flLMDdIqFdHXjDI/
5f7n7CBnpnOb/swT5Jo9jFkTrukFhMdpAnd1vNyTPXDyGyZm3v8/WT9RXAPUHBK0JYWc+dUHZfps
xPBEnamBsLbB1OddgSdOnZthcTyDIr19wCVQC7bFMqUJY3v4ylg9SDrzJ23Dvvnil/NCUYML2220
gdsxbL4q+/mquwJiO3Z4Lr9WfEuR6DSjBwixHf77uOCWfS4Vax3vt8qxXEw9snL8pD4/x1ehT71z
DsnYVnpcqhPtnsm7n3YSbjclHXBbOYjXjbu8qSEeHaqhWMJa6HieeUBFlGGe6cFywoXQi9HmPa1j
9gOmUQ6o3JjeDOKoCUw0azR+l8YXwNxbjIpsuSojV4u36dVS+w+gOi6arQeWgBL7qD5b8FPVKIEI
gdnnokouYkzPGlIwOXnrwEp83a/LmU+LeyXyJ+fFsjFDLbSTJgRCNHOklbr/QkiX8UaEHP+wgnQN
plO5BYopEdtCwzpkF93b2zbs49UFwsV9hWAzzn5q+60WPCtF1vegP96FCvUkj0ripePSPJOW/RXf
2eYeZb0eRJBj3p5hqenZKn0fXCB+7c3gh55BUYWg3tfGj7Qucdb2Y7t5Y0EgCrU7fh++Vwu/Y20U
NrCQSKETh7B9n7mhzohr5m/XApwMqZ6LvtHA1RvIqC7ORmvVjgl+TnRUWFhU+gx1QZ08CDiu/ijh
5soEGhnf9GoiVkRUCsczVgXpbiSSnAk9A4YOyGnoMNXYJRSINvehAySjZtse31ujhXff5Cphk3d5
1szyuGI9U+3ImoS2gkw/TVOYlceBrbdikChPdbBL7y4bpEkuW/azzrSqX1M2zk+HSpJ6Fa+n1FbQ
bBXz5zk7/q6t5kfL+dhJhgmTg3TcY8UQRPBJDEmA9lr4P/A948KOLSBo5tK1MXN0djpwkV9hiupP
/5wOoFIny7mSVjikr0k2qvVXhE1Uf40RB58d+fz2r42UGoHHwLNh1FdXTnA+ZalguRuFZatXhyR1
uLvKckUxw5UoHRVHQK2iJYUC9lOgT/H4c2PE567FyPyNV+nSLZzDZyEPy0wKc54+h+lgB5iIjyLq
AtLbgw8V4t8I2ZkmOqHFQjw7S17JauEOx4AbIVIwhFFTfF5kRDL9dMXKWlskCkNodFgYT8k5fpuy
BYnYxAqAh5su2HQwYGAetlWFLXM/6OBvB29HAo2aZw+6ul+wSeKa8OrW+5dBM84CLKtjqkzi0tYh
99imYw0D8sk4ZKI5tuADnhD3dWYoDyK4efiKG2SuFn04R2ygk3O67T7DW9bd3I3eSjdxBKwWnPjW
gEJIWeCbAoDxCTYqqQjeru3CLWmKTX0oSMJTT4SJ2VmhBhY8qz9Y+/ZHyZIEyUw4mbrErNgGCQdm
0qqa8D0BtZ82i8a3xk75il2B3wZuI5Yf8OWwXZo0CCzRYFbkhizawrxkOw7dm2af51YIPYxZKSf3
MSaKE5ClZk5/SD5MD0swINAQsYLH6ktdYzbLvn+9YNR4KH83rylirqJnPdE6RxpiYAoJHO6wvT7F
Wk3WtjedR4LRENGteFNfWtr5qsbYWc3JtItlqwJlBCLjAYLSUXGx6lKGAfrk2nZEJr2vU6gIS2Dw
c5YuPLIzjeyD8GgZcRm2CZ+pJHs/s227HrEkXwq98pHWU9Q3TWuJdTr74FyUKduX3LZWwycqw58I
uw5gt+23Wd6DY5EJJg7FVLefe4wQHO69PG5bgkJx3vvrb3zMx/yeDFyvTr+J/Q6nwt6CD1t/aJN2
yZm/nPy/7VqCcZY5UUpHke6M+3xJk3aUBLYezw4+QqyGj4M8kFehB7+gA8f/cQo06z4IKsBbKDif
L0QabJH2/lFnxwBhAGarNaFbNq01Lb/jqSw4t3FuXZagOPJx7ECOzX/ZqUhuKMWlwzO/02DsYuNo
zByC+aBWm3n1AYJXiepcx90MLWCq06MvWmaen/35ksM2NGm0Jd+kfHUE7I5LKtzKQ7WCjVROQ0jf
DG2gdZDyv9T9AV2CzThXe573Lj/KbimcsahnYp3NU47F+Yz+9H0wJW4Kzm2KlPeEJENkFrir7MIu
Z6r/KZw6WtFc9b1AyrHu8NnVekkZFFXUg1vPBILv2pCBSK/9JknevgkDL9b+X9/QxS1VyLSxriXQ
zFNymR2LA5p60X16k1hpfYZQo1RCucaWLdZ3YsptH8DQSDW9wg7OeJ7q/2QCvGOickcnGSFf1mCi
XDFW2qJDc5/cC/EZmplBqCL3ili0A6/UCWPsQ9raZ9tn9VVFI4u9BBBjHqOyhZmP97HeuAhDoMjO
1ij+SQrAwH2LQ9JwqB/9r1boF4x7lPH2AD2xX0AETxW4rpNlbkOmLXEzQ002a9S8w9oIdgsLyhld
+PiWdT1oupUq7BffpA+LBNL0w9WoE3zoieQa6mF3W7ntX1bsACb6DYoMsY0C0NAXv6fU/qDOIwrn
gbZK+bfZ/YOlyRx7UsBPbJEnr3+fyyQfWqzy6maacZXI2ZVAEWWbKCFplJV8V2KfLGUdILiI+iw2
tr51N6kMWUphLxxew8O48kPbqpaUxl9wcM8ymttmF7vIq4t4ROSjIRA7xymefy1glcoSBWiHcwrU
oQ5CHfZNpBilMiBjaXeyLnUgDQQzU+rkTTHbYmJ8hcWB9Brs6ALptG/ai7H3OerZxYIpEVPgMZoU
4kqBtsSVjlK1yEwEH7r1wBQ4EoQcfxQttsqpzB72VaMmM2yOt+Ma5PoNZIdyvj9y2f95VU/3VqiY
+iopsz3jfe8tbTZyxCT0pqmHJs1L27OwMeam7DMj/21b3cjkWeGfShlENOV9+sP7s7Jjz+iYwEYX
okbwv54trJZWHfQO3YPqH/odUdMjqIfeEQujYFrsNwLpRaYkqv449FzDe3hCTOkEDUb+cXgJUqVH
3P4xViNyL15NJX4aqkoRl0Kt63AHiHPukS+pvMWKJJ1nkcj/2gqv/rKT8XwztyWMzFKHhr8eJ8NL
h3pwHfQRN6xE5aXfm9k7D/BKtcSCRHWCLzgKmNgb4Xk12+IS1ToBq8jq7GbtubiIyngDFWTfj0z1
+v7rK/U71h+HRvN1pXxPlUlQtdSUbejcZtA2CbTviNq+2KB0ecPQHYlErWsadE3va8KbEQQgi+E9
ZoKtnZ0wan6w9N0elLK55EYkWQZayAGA0w2qVZk2ifqWUCIg2rfybbZXTmGcR0PY1ouxbBizi1Ao
O2uh+uQcyYAAqX9PeKPoIB82lbjSlzmuaDfZHsevsOM60Ty+7JaFiy6Min4hUt9ikt3fUHPSv6r3
JxO/xwEMJs9OSKJYIEidFl8654n/r+Nvm6zrlmAKHoGvPFlbem0kVnodJ2WZxeShdP70gD/SDD2P
PhDEz2Ru8OcDMKQsLu8gl8R9LGY6VFBH6K5nIjuSpOZdMCSC7Q714I8T626J4FNHfIzWzkAwinn0
Wg0YSakPWr8cHKDpYEWpiCxR7P+r0eimQk1SsIUk4EWqv6BH1tivyEznicVtUSeFuqrkzW6/h5Rm
6TLQpLyT8W3bCimgSclAzNjJ3YjDdcGRtgiXVxsWJXQf83gKE+9vAd4fIK0eDp5E48K0PPD8SxmQ
Wah262I391VnTHXcRrPaD0O/LRKrg6NLr+JPodrJEH8URwWHZJlwlRizIrNxey6Abih8T0/l/ZNs
TAT06LoyMZB2ubL4RQzue62AI9zYphYxIDnLJQnW7+P/K9Nz51zcrHeSEjDC4AeMuRXSaP/W2Fj5
/XTOFHGhIsd4ir2VvA44SHFcWwtEZkXYh+VaUX9YJNK+sjgtit1qjB/kRedGojmafsk+ZTLInVK7
gzOLFmztJNCQeFC0HzBOt7Klr2RmcJ+VirGOmtGbwiVa9KZ5CVGKiLiNoQSeyydC90aEypBnzng7
IviIMdCuKsWnZgHjgrB3FDSteSwvqwyi/tUG2JJaTp5tF2JhPe1UgKiXrOdh711pDE2XfBhwqSh/
/fYJ6OQOONfY7j+bUsUeF/mP027vDiwLzj6qx4B158/nKBC4+o0s/+wlLTmOjK8veIlWqmikJ8uH
Y6KbSzozO8kiCcjN8+KpWw6howznDBz3/ityo0JTdD0eOSpjJiPcSpUJodgp7ocNez86RflThMIP
x354rRhWLaOLPq9XjZYgSV2gWMkwkRoBLfZWYf9UdB/KfUulN5nG9dGE12z9pKZEa/GyFp0K4Cnf
yr+zkHFS8FDTnzPzMlamqYlXloKcJFT1D6/ZpMktsJ3cgzatg9S1Ke9bTpT/SwGq/XVfxSJTX8iO
+Ny4uVXAuGB0PKqxfwEfIpLuqfsHKCJH5Mzq5MWgoQCrwi7F45PBaOZ/OF+Fz4/GX3tIx3Y2NZ46
2thbQKQfNEYXnNHu4iwCkm0fosg7m4STuzbkrzzvliMPLJL0hduEw5tMCmoan60rwLclDNuUnb7C
JAEx4PEvpo4I/Cx5LLr7vq80p7IAy0FwsGBdeA4/Wee3HThZX/2O4I6b1jnUqBS6IKzIZXftdhBC
OyLsN9lfPixQma56MYlMSFM6o0F5p75W7/Cb551VyAk2bk93SDHueBWF1vJuiJFSlG/i3mWDR93e
zhvKccIxy28pHctPJsW033Wmq1ZtU3Uc6uqtqEZnoVOtd2+5UtagXgUkph2rb9FGdrt1DO5cOj38
hEpOFrWOBdY8BqKkfi8kQVXZazoxF7alM0+7toreSVKsn7BkEs2EoOhkFDk+/6W0XXGehHyCBxcj
0zIJFzOWNbDhXM7Ua7shfrGAnPNepzSd2gxBuoFmVg4bkmC00LV+KtB0gUGIUjDMKUHg9HhYvngH
Cr8gEFmGxTo5IVIEAxQo56Ef3ARaOgucu7PMrcAKgUbrTeEE2010Va+1BU5OF2+xWGBlzNtYPdEM
iDwmwp7KEHM59PWPUAVu43fXhn6uOa3AGTrATXrQV9N2uGH/8ggJk9fkW2dq18RJaqlfJCSLQr//
zi+qDE858GgmXmdMzGJKbF/l/nZJ2Iy76TICcqrTm0AYSDdeirdr4kU1/VuNNovE6QCRRw8CO6QK
hZJUh5xJ6JRsF515VTpTcnAfoK+aByTlUjaZDzqowFaRtr8N8PuRI1FzWikT/6sUZ+Qm5eQ/Mnr/
gQeB1AGo4vdRfZIak0oZln/7Y9Z0KaSkMJHc6GHoHaTk1pX31ZAjB5FTfUvQbK0R+WdJk858pwEZ
WZ1t4+ov7So8fzD07OB4RN2WsjSFl4jYIiIlbGhctarGLVBki2oBh7IcdqCzbwhCRubgs1xgJb9l
P830m2gcEg9vgghliqlEcNwfixh9ElSAVO4VNIPBA6C8uH82DW79blu5JwW73d8d7fjCUmiVKgT7
2qKkyhWpggAT+uqWByGB04WaUmwtUWWEFQ0BC0eoYEp/2ZxtyFUeQVPHIEXI5kd4O7e/fiXb5u+R
0yagXApwPoU9adiThkxDZTZ79PxmV89RCEMlsZWRIrbWbP9th9FE0VO95+xFTB449QST8eE3i7Oq
38i0hFPaqtpXgM7BaHfKZdfKszK7BucvelibAWW8fin5JnobScgCe4xCLfEucGGhJACkz0qZLG2i
asI2sMb9o9IpLftzRtnkpSpilYMHE1bVxSkaxuNVdsHBBCfF+MK3KcZMOv3n4BH6SOT305NyIkhy
+g3s7fY4cWQK3fnNG+Z5zR/GnraTnD/GDboBunlW3608InETAkd5dsEuMw26Hqf3206VZvETOYdw
hRywFwhrm5yxks/UQZv+tDDC9CDCxdb7kr6yyUkKKJ4zNDVEDmsb2/39FBTJsBg2KrBaKl0NYd3T
2N6iwsKNelD975Be07oYIym/kvClXc3mVWBQy6uP1oaXrSjujYs3leyG+9pZ1b8mAAM92U4sgsJc
/vt/omqSzfJ1HgdAbunDHueSLwDIWomOf0VuFICs6wua0lEoi/2kQ3ux4xMrqcrPCU7I/t6bBh2D
JXJ3BclGgx0RnOse6Lis1MMZt+fyYUpi4NiTwVeYOC0sTsqvKYf5JuNMm87iF6WNwA3aBuTZM29c
45nphVMONcwv+L1lSoDtwrDDJvLi8cObDT2ivx3pMPN4HvLTnwq9Vq6GQPqYV95ncW9Ggi18yU2f
trkJCC+3cpJjXWZ0aMf/S5p8tShVBdWmWE3LWwkzQRHRnC3uwveWB/ax7BvqS7fdClU6xswIDVZ5
2TcAJi6WrPlAsioRP4kgLoAnQQ6CgvlkhIfOafJeDydWNTqgHciVGzJ3WkRzbR2ffCe6Uo9ZQ0GM
g/lgmJZ+YYNaL+KB8zyhqms3/7vV+6BGxFpMAduk4FxicQliNF+rP24n6MmEqhoqwT77xAwd8VCo
+0SV5mFnYU2fAPr0qc0rv7sYBS/InXD7irxztzq6GVw6tbdFEPpSfkuIEI5UHzv4d0TqmrKQ2CjU
rAwMEHrivMBz//DAoebICUchb2fIgKC81+Amg22iXf7E6NTyLZhg+LkaTgbcn00fDtAb0enq1ZEz
fk0YKjpTu0x94usPElnwH0Xp8elQRblxDO/KWoLA3kjEWEq0l1laSDUjnNj9wvBwZcomcJ7fZmyY
62N6ZIQ7rqocMWDBqTWN+rZslXUoKu5CYGLH/5lwqDfH0JPzrBpq28xcScOoejCL65dhjcDJ43Or
gO/llXQIjs9gGWAK9r4BxUUoS35cEaBolMPoo8u/0MwTr/NC1CyWDhBOzmz56Y1UVpqLfZMphRdR
JrehGYTIJO/3Cp3iypzeIXZD26aA1mDmt0SZ69b80takLlPpACBXaukg2Ylgg2TEa3f1C082S06m
hn8e44akjn8M7Ta7iGyWMdEHEL1WdsjWVYpX/5ULEMr2lITNb6sK/g3GxbUUbABYDh3F21wH+4W7
vebf40JA6HG0jngC3NMtSztVNxxmJyzcGSVBOmXRXwbe0EBBqXoPVrBOMU0LPKGXz1RjQ6/fQTDw
y1RcU/cd63LLSiIbdHCbagoGwM+jtwtcqSf/s9FaE3w6XgyiZfHrNs6PYifNWodtnSSEooAj6pKA
YJAehhba+R2k0pakvzNe+FJH+ISK2tpkxtmpkQIWTlAu9RrT5zD9cljxD9e9yk4iP2VlKA1PTDHi
YlzUc4raLbrwRpATLnGMesCoLGg4RDZEsEpgBjE9wAaHEOdNZMT1ZeTQg2FASu5DhwFAmec7Z6FV
KGPmX24MgDRoEGLMvCdpAtD75fW0t/DR5So+1a4yORdet2l4RB73N98P9TaJ5xEieOWCTaNz+epd
MGER52Mq2FytHgQ8VvHqFAJe9E8oE5yFgpZ9xbiT/yzLOeNA4YvCQhbqJpd8f469UGiUemvyYy2G
IGs6leibiHn5W6Xft9myZ26oOpKTpcKIYi+8heARYmMGQllp9ezlFfxSJHj1YQJsbghP/axOhSjA
xJXnX0BIIxV9yCYo4MnQoh1TJPcRKMreL8LkVrF/FHlTREC4NAq2/o1A8W673IzHh+9MZP09YsYn
F+PL2KDb3FHRr7f6UIYfwGO+tG+DW755BRYyRD1IOUBXp+StQbjGCv0i10xYj0JFDNI/+Cg417vc
MWikXggt5v1gPf8W3aD1nmqEdgAoLIg4U12n/fJPADy989oXtl+VMFMDNCovi55x27Jn6i5G3T2I
ySYW2W3oDRrMp9eaP8O6DQKxT0tb66hfcPr2FITKLBUCNgxScD8K29KGgnESqUHMkLmlRpbMy18V
qFXbj8oSOr3x1Tb/+ABBfKx17nqmCYN9JtXAlLLGBsvKiiIBKQN/HOG8IGBXVGcF/7qJDS//qal3
Wgyy55DdUHExe0FAZ5PSHbSo8675Lcu5QKHFL0sGt0mxkF3Xgdfk8W1+vU61Csfiu7Mmkw8p+nUH
nPQvPmhvOUgun8lpeMaoivw2RBts6CjwGI8u8SHQsGnZOsRV4BJ25KFXJbOFtE/l2WHqyOEGSGbv
+mUnE9/4NP7oT21sGjvER7xvewG+WNs3ikFZ+OrRVXIRzzssFKFhgBX+BiUHAXQ9hcUQelDELvjz
EonINcY6oRX3M0twhOZhAUv7TKTAPG3DZyghcIPlG8eXxgWrLlgVj3Hn8NxoSbF4GOwF2WxzDYAI
ZU5HcJqXho4oKaQShGMmlf6cwjqEUTr0xDACJrBm2pbhvWZtYsxO63qlA7jlhxBeIwyG+gGFQmrh
UVm4gnZDcBVC7gXYfz18huFmFCaTpxnwfKF3Yol9SbDvAmZFMzqSanLvurDfPMNkOLvS44fMATS1
6nVeoWvyMPpsUPewc3c5sUZJ0iTT9DUa2T1VxU6raTIU0789hJxJDOUTWYrDUbU89UTbZHJABGmy
99VjqSxa4SmQw2kU2rghhnQNKN0Nf09S3EIdIDokhij+FDYtV04z4Kms9xBfArBtXtp5CSfwIoWP
fE4gJT38wCTQkU+vwERX8cDhkvo8uvNk5VntNYIKdH6v2pV51VLKFdlMyxXdb9bXO4CT1X8Pgj7Z
ybGJqDAaeKqXJuw6+O02DY4BCgj4xlF1acJeXN2fb0F9RZ5PWNVQ/PZUNm1mwo50cOUJh9FO1nqI
Lus9imIf04Fxx8wcLz+yC09/SSa0eyEsjs86LZm8OuG42Vw4/6Z4HaytliNPC0qLcmXYBwwKz+ru
mR+D+EN61j+j4v7EqAXfVPBvU9yGD3BGKmIxcx1ctmAcZEw/I2LGUrJoQmhaNbi+JaOypGs0djNd
gTvMUzvjkbzuxSqWCsZUa/dTozenxr4SBh6SV7LOe808Mo8RmCxMyRpU0hChnXWRWe+UtFohwiLH
htP8Ju2m7ZWUSCIVmd2L6+aPhwSe/8GxHGYeqpDodCs7cCACMwyzFi7tu453g7+WOtePjfZUiz3A
Rj6n6FQIgsWP0hUl767sO9Y245Ymh94yWNVeAUIdywK8xkIeWwM3pu73hckvUSBghEVe2JYcDVSx
jDisg+4MHqY1VdwIkCf1mPQsv2ewlaU+D/2eq0kC17vGIhrxjfwcWNC+IRJhFHSkdD6LSXHXJ2uL
Vi2ET5jqUwJYPRGbHjqSpMmiZ6QWPmTf2MaE5wefHttfcGxzl347jQRQ5EUq0uVlzvoMJa514d7q
L5eKCmzyolkDcsycXu7t04MOV4fwpzrAR6tyywuxlKMFX3DXzYfbR4x+8f0aKMBCzylDt+tU1OLd
wrGe3nj/wiRkq5ZQVlMjuOSpFt8yeLf5enW+mLk1HredWkX9R1UaTXbVc4HeGQPwuiV06MKDqUmH
mWgZsDLZnjxCtYT60dH3VNBOHeBecnoLseD6nYyFqjDNUQPZctd9Eqb2YMytCBQbNtVHjVciiMFS
lP62wSU5zbjYNQNnPISFH+8ehUCAPsjWP5nOi6V4zZdD6Rx/ZB8BNqnImCCrwbXfx3XiqDHsqq7c
WnBQ4jxDQcs6V+mCE81mYB9n+l1WCv11p7aZs/1Yn5eU+qwETKK8vC8yaJMg4Jzh08a8fgfl9xxf
EKtYYamtioD63AIvzaPb4PplFK71jlgEQPq8TLsE6QNaAitqWVriCTMq1wBOgU05K6pbp7+DwaLr
YpV1u1tOXKXoVFPZgRVaN2m+fRfHOf3Ae6BdyJnGRJgCnWStSyTRce8co9nPNWdbWftoHc+oh1l4
Evh53EPwPtBTIUxrnIGmdqjQXeClOAqWtsgxwSfuhXPVkV7PWhqOVuZ4ejtzUFY5KDCOeCbzOfOx
Hmlyvz1h9gJNuEwMKO6srx4PWAroAt093MC/akzEdv/RrY3yKro5JKVgZI6sxT1RPpU4cHCOQrlu
2mgG50RjG4zTeR0Xm/IAri5uC2Q6eaTqLmI39FrNu1+vho44DMy8oSSDFxdUkx6oZsORT9bQ5k4E
2Hq3BTU+gUtV6O2DfYoFTjXxvDNO0rKKo15ffisTpIuVYaZw9Xlfc5+PtEuqL3BfraA8ricEGqll
ZlIFxOT9ghDMLANBNSTXAHCOIZo6etWa+tNFWZjR2Q3Ks5t9kWSsnpekya+4bK/K2VJ+OppUATLk
EJjkM8ZootrSDYJ4g3s1D3MYa/35YH2UiaDBjARp2SZI1T5hB09qgtjCL9jM4F/+Jc692EdLc3Pr
jodU5pMMBRm1CxeIkzxaDI7M8sONQXswmSWKCAu//zi1OTkCBF7R8dFYpFehS7u+2lhnvqOBw8xA
7+sDwChe9mR2mg7oFcSN9EkAjEiPWCO9FP89RQHnpA+8LEeoLLLZiAqgNEwUjWgWCkNLqdNrTngc
7sq+PLa3dQOVQL6Gj1+93GR3Mtb7gA3M8SOKhgMEEkLaUZJZemYlwDZbt5XFwGnJ9O+OK5gxR22R
F8CyqeEItz3CH8sj9CTPpNn48I/4E509oZRW+WKOMNZ3hbE9NtxsYflgUvzSsqj2hklylt2m3dMf
012Ut78/I7/vlgqC3uubhcyPzR73I0tRD8wg9Io424Hf3QMREvUwYiG++QGPIUSJ/AbiaLlEsz9m
cnBNnMd1CEPGBjmer2kWxe662GJVUEIe+dgOBMLDouGanyspJwLtTPq/tQBjc0UOPp3KRH1fT047
7YdR7y/+9tYGsgyRntBMOOg/Z2lEW7rK7hlSIhMlbwI2Hkasb/BQFLtv4YnfvRdMxvi6J8mqturp
cbZn6+5NBz41uiNGQOy2zzZsKQSwWgAdyIkNzBidbhO5ZdWN9lKPPgh/3+/7m080vXq8NxVX2jpF
8oQcz7a4PWY1SeS8LLcpevCTvQ1+ZgcljHwak/MGhAqKantr6YQTtE9+zoXfiXEt6ODvjPhmFxxK
uYJTek+l7qE7Xih/19JAj34jvsPEJA4ZdUdlPptYzryvDuNS0ZOpU4iF578+NEMRDhB9luofD8qI
PNczo0czDxANjv6y83grg7hy7Y/1hjgVqzTZlTnNQ5MVUuu2h+8ChRr1PYElSDxn+KUgIVGG2JoS
XQ/7QAZy/XogUuOWiTwrZMAQZ2ejwECFsiNt0DxZvKlhsnIrh2HXQiTWQsv5PzHfT+1n1x7iNQ9m
o2ge092c7/LEx6w/I1hwdNz2AbSR/s8SkZyhM+9vt07kfyzt9DNYAmTvo/XsGkGpeKaX0/Tmhmhe
dphOa2Izg5KHh/sK9KFXwt+oQggoJ9BHU3AuJzC7YpuGWpvl/8BAu+ocmIh7iKrJ0bkq7K7QRteu
6dGnc93CpG5XYMKhT/G2e799PrDCPHDcdXjATb69Bzv6iizLLg+nWk3CKXSmPPpEBV4sFdTlB4W0
YnLtg5ch+/HfyAoLaCOPHkWVDKAa/vkrhI3GZXzP0Lb3BwauXvhhBiejiQDDBPAsnWJLPwuKgeoz
IvPsUCrCR7nx8sZ27ZAmUtmWnMBm+4EsWe+kjbMuRtNbdipOs/KiF1bh+OkhaF7zKMezpyu3afsr
s1qSmNbmFQeernPj1ndZvK5esIJTHNVhn2R9CKreXDteacPWAi6DLC95m6FSz3KRg9ZeRtxBI3Gu
vu5gbeoXhDemZIblmmpM6ySFsuc6VCUj+78WdyFkxCLqdlnvgXrPI6cbeuneRqbnbh9TnWWPGtGl
EoKk2sKwYsJqe/H7yA4qTiG6UzVhmCkUxz9N6in9hd9fM7kTvWT2xIp4ZGpOrviWjK9T8exPExNB
ntz7mBbLve8hY1GrWMYk3IGVxnMtVUSRJ58SVRtHIlx3c5RxycZP5oBAZCu1IERC0LNYJSb1GmhG
9ucYUOyetHJJoEDWPVbTaAFBJhNR+06EgbR/ZUg7kgGmQ3yqVg4tdFiTW/FIQtc/4FBRGhBZTaIS
AO39V0Wts1oE1f9bGvJPhBsnkErmUwc2RiWI9TLhwRMUYQkRgY3jDbSfpTxaoNlBE7F1X4zHygXk
PPJUrUSs6hqWOxx7AL81HFG3vPD/mloDSTn0Du5ZZ3k+uNSjCyIG0sTw8Sglw5ockR38YD1tuz9s
E13QugEOigDL8RBAcjv4w0S45PvOADUMei4F7NStIvR4Ghg4RLQ5XAN1YE/lRE7BoATEKhyvzofd
/VCxmVEfFwreZdtrTeBCdpB7gOTSamE9scL4+7r9reic69E42fl4+Vy3TiceYysmt7Rtx8tQxDyN
tA0Jv5tzNuqKrqcU1KRbNj6BcffcUzQgKs7YseiaqDQieTobW0CBLucejaFVTjMC6Mx4tVjCu/G2
bV3ZH4tMKWXSfA6i08g+H7PAvdawYlyUNL9iK78wwkvgpWGXqCs0hiEq8AVbTfYlXIw1+UrnRAPX
4ZB1wcFLb8EkYDB4ftw5uEZD9HM8iaeq4uuW4+AQ5IJrypkqQvILmrRp58CqyqT734rID+sMQQau
BdVn2qZOotTnXLJQxPlc5DcLW6NroKd7MlTLyNDVc7CQTgFtxIwdCR6bgVjN04pBtTLoXznoJ+py
fIRt2m3Ry+72Q103lljBbx7KlAUWyF2cTSpu28TO7BVCq2m0657oisDrMzEKEs7yJGqxvL4cs9qA
EGJ6MNkYBxMYhGtMHnIjRc7MXzFGuoD5njCs6hK7/R/UM/OviT7BM8D5+k1yl+JlC4NiXaWFvgA+
iGlH0ZcmWbqi6a+7Po+9EBdtxCB8JkFb4l9ZmQa7eEcwWqyFGaeefgzKAJLWbUWHhtZUmfN9AtyR
zvbE8imnffKiTrPevyhJPNxOxUpMf5/aSnZnGd7+/cfLqIZNdNAwHDVvgnGoDGwQg3Eu5bdEgFI+
yMXdNKIIpk9RUcx2aJ37sWUYIoT0cLUyCX9UTdhcmwSm+bRxEsgffvSM24t3mQCr8rS9+xppMzpV
Ir/AqbDJuEdGi/FsVBtNDE/M9uzZTc1FRv+gCBC5M4cz+/wmftkcezMKICT3nCpIg0911iOXtlrK
pSkfJ8iiqggbWR+ljTZu5/ZL4+qwV+RZRUgU81th7pHSgn5wXxoHR/S+YVoOUmAaJ+/3eKZhVE/R
kWPfsSi732u90ldH/fpq5/a5uUBxlrujqr1QILRlKGRfwCwHuCxen+IpbiOFqo0Q8vJmWiWkycI/
a7Dmqq9mqPTHvsz3LVIgQtjfwBgmH2r2E8Hv7CDjnvIp+TzTkVZuZeluOTpRFLWdTi8NEnvdlzK5
ZIg5Brt9KurdqAoBgUBrTm5Iu+8fvYW7vJNiIq0E78EELHHFk+ewySrCiBMQhVTFO4TMxQ1MFYP3
I+P+pYQSgl015blfjNrxdZaevrSyjmPFw+WrCUoIFUhPGOhZ3Owp538YSPh66aO6BuuA2t3u71xe
w53zqGofd3SNPNHwwwAT95XR8Vah20Wh2jpmgLScwmBt9LL69Y+U1S7TY4owzv6gwuphhO3iUDyb
4RVp/2Gg4MECyFivaj7whhHFMgrzuOVnBqJfudfk7DBn+HdbVIx+Kj0q8J3kRaqMOC5bdZb3MJew
dd3amjWrzfBqdFj42uf9LD2dXJZWRzbXj5rELKjCWZ3Vn6rBwaMxJGy2vmupRTEba5qhT6DHtCch
EFtKrvCw/JPmnjjh9UWk9FG9ie9Yw7Qklbn8ts7P0aDyUBA2gSnAeA0eQIau5mnu/Tx4e6MiLotH
NG1fN3L8tjd8Wgmm7ORA/SrSOiLVEnwa5fyH4LM8R5mAiovKN3hWq2Rg4GR4rmF94mdJcr1tTz5J
0Wce/GI19VYF6AjuMN+6bpkU7M5iJOMlGtIPYPe86twoS+m0T0s0sB2xTStfP5fkZfflbA9vUOWL
G43GjAjcVyqfX3vvGTDg2Zoa67lfINqvKqY+l1lOc7suD1iAA2AK1Agd1twUzdpgzWnxskYPpwPu
EeB8kR7GlRDssbMY3rLCktEBUh5sh98NbRK7OAf8XVWmgl01Q0h48F05lbJXVC7CjAjmwlii7g1X
evxyMNzdZFWaYyprfl7BEzvBf8I5pChymRHbto/2xtk9LMKOUvLh43CtTDrDjTJktlfJg6aXKOqY
8ZYi4ngBl5XonSLYgORFSqMto+qNZRvJ4eks3d99vb0s7TZC6/HXyxgRoC+Rzpr66IU17DocE49a
S/NvML5YlL9XJyYC6uBPVQjH/cmd3HxpHJDFJXM5VD+y+qtOKjuGY5PO4fcdMdAKZRAc8SBIyHLa
gjBQBcjENym2C4h7UarlDFsiMQtj+29xuZPC+EbHZL2LUKJ2kz+KieWEkCE+6U5i9c2rooFZPtty
p3Jv0fcjBlXlbKnoDeudRW/XWd1nnsem5IiOx2xpUOJzo/h0fU8VNlxMB5whYiFVmn0Cm+6TF2wq
PVgpkMCdIwBm8Iov7ptnIm/9JSzpG4g5CHEbab2NYb0iiPI3MNvitNfqib+25CemNQAl3AqUHWGK
2VJQOJT2dhdDtxZkXR5RhqGpRRVCqdh23xrQ9OnodoxTo6vPJcwQBq3R7onORYpzm5grlHBpcpO1
VujqK1kEWrLCdPE8C6T+sPQCG2i16EXC+rNZevyxBkz7kZXXFwq+PtHmCT9tuvGeCFPPtFE2dZPO
UspNovO5FgdSFm/Gu8u5vNUazEWkO5++qH0BZ4QFUbTQPPZefWyayJz8Jt1Nsz80KazOV3sosVBM
e1tvLvU+f8+bJb0QPfjU1721dq0GqM4/zpr7Qrlhw4JsbCnWZwZWdOSRAxD+rkdnLgbqTCbu60Db
90plX6oXXyOFh0j56rYlARAS8Di2Q0swT41/5RsBf1AQoBC+ZFukGiAcz3+VBenVNMBLReyZUeTE
z6DdtKJZXHgszsCy4SjUzQcc/oTlDeK+gosR6atFWI1Rr0ZGp5KCPbYUe79FR+tM1mMNpQkS2Va8
O8Ke7OH68WvDmN3ub1/uBAil+1tNubSojiA92JS8ikfoTGu20R18w4pREI1NilKNbPFtgCnzVRFS
p5c+SVyJGywIbyBE5BXW285J5yZLsyUhkxILRWxB+pnsg6T5uiPL3RxP/C94KliJMZ7Hws3a9ebN
/dm0Z6ybpn9ncJlRpzhBA+a0yNlPHawOUzOw1JdjkUowQWDECF69TPJAfsN7tsCqLrRsCEFncKi4
QtT/8wLpSEaDd6FzbZWTNSt2x00zrX89bfGog0YRz1nsRomyp/PiO4Cca6XuJDP2D7pAsWbP6TKu
Mo5yMFINyPA//TnfkYS/+HoYkAzRZeNS3fnYeXW0wEPcIOub25szkoGThCfQMS5zmkb+alEtM6DG
zxDb1ucJ8dPzABgde46GqRNPVqQXPiyXR2/ltOxK/Q0loG6/VEQxSZRL8Zn+1hKVW04xpAM8Q9SG
aGS7O/FGLluirygKJIzIlz2k0CMtlQtAto2fgIhgb0pE83r60hYGOv60eQGNhpUgSt1drVhlneMj
uAgOmG4i6zYZ4y0CyZ97WFGauDso++4B8r0KE81MBBvgXZ7yGgMVtnE1vmg25waei+PTyxm0aslF
tnyhqMjRmm7brydTDWsim93/9a27OqAfX6miTKtkPdZcbcfYoGkS03j99BgJEiFxxQhMNX2Srf5+
nGI1KBTDTS2ow2MEcrSqTcfMmo8gy5yZL/T6tja5rU6CjT+mpQkV9/V2v01zq0/WIB1ABXWztCTK
QZupeIsuQzRazZfeaLyvD/sGAwkHWYn6YlW8V8Q1NQM64PaXGQPb596qO/7X9uAmkSgdfsdJ5UeF
wIX6q9bXRgualhg4kBgcQhiHkmZ5ivMV5hIjPgox/54z0wFE/gmuUGGslvS6+xYMm5jgzlqnwKBq
KS9oIe8dSZSIv33xpE7qJd6E+K+ukM1V2fVGGlPwethtFFz3raWRJR52XOh47NZCYj1Nggk5bulj
UPyYGW9w/9gaoxtUopR95FrepD8LbvxtNRl/We+OTD8vm2PkcUWX5OC3fbafmy+vWi/WKsKa1wH9
vvSUIwxvlD97coAJtEIDeuzhllCTtgPCaHG3kJk/XNDu3uvQpvis4MFUr3m6rqzaAXWPgOoLS9VO
ZmJj3H6OYT23H5+/JpNpo94mvc5MErztGxmleVssCZp7vDUhWvIiayGTYBjTfrzYZavdlbLufcyl
QFD3yaIA97CpGOkL1af4DAdHcbm0YsQZx9XAu4JepJIpoZlgKCYrFECB9CV1wVYPCXo20CT6k34+
2lNfNuBue6GA8Y4+XmWE0VKItmvRMdtSL8tRVFlw7pX2aqwBUZd0jF8/NNCrk1VjSErU6sh80v3b
GIhzJx4MUkr3R/pRjNmwWxL63kqF9K75NWHZVg5t5BoY291T36z91RKy2HUqzTAFIjbCH1jWoimj
WZgpmpiS1ho9chSTuxDP4BzdNXTQTVtqwkpzrAuibJmJmXYhrEE6Uol13zjurqyoU2BBuxyH8+pv
Qpegm733uq6cIQilc/QhQYYLxawShTqhCkB23VjIIvkY+oEwpX/udXbPI3Msr25vJmb1G3+Xq4EH
hrp0TkRrFTHbpDOM1wZbL3620fUv6lf8uYEB7uBamoJbjPoaa8SbmypE8Vv0NKBVzwLuGL16K2Lk
p+uXh63AsGvC9oY550IuF8TpP62UmRSgJ8mD5IdxgP7/TJA1TR6EcKJ7e7EDSLtqDcXplayKclNy
r71B6HUaZOb9OQm4cX6CSTaXR17XQsiW6SKUHsWxz2IZaijGM3jRz3jYHTDOa8my/9IChHsHVc6l
7SEK9Gq6iEJpe2hejPY/+irbgF06WgoHC7QHHLFXhWsDhIqXhcaHpzjtylr+WoS9rVKSiWbAFDVr
kN6yzrrJT8XU965y+0d38hPPsOZshr33eLpIWsOZhLzS9A2ikvMRAN/AMnB4L3KM3Vb/06QtSb+b
LYWGhnARfF73UWhRyiSsoKdV2xzUYTRLqyZdjKqm1ZAtCVtKlh/rbAjA2n+XbJllyOkbtshnnQqY
29krdAykJE0lOtnpJahHZ2uudzfkxHN7rnYnjnVWXf5LN0N5KAcM0tD9xX9chVDRvR6ZWcCDobJq
LNywYZjs40bvPsU8d44JQYjgO0ix2rBvKkcn2pFz9p56PgUec0GcAz8+WMFXD7KjQi5e8boJ5Wkp
Dz1Wr0nOev+ZkwbnNJLVFGxx4gRXudzKxwlc99k+NuReNVl2wcu/uksRvC9KSxmqdxAorO0n0bAc
w4bj5NGNB7zyCJ8kmsSGtV34btxBN8X/0+UmSEcvsZ8rRnKkN3U9yoCVFIryJyClbNuKd3Y5BkKg
LBO/hDEYlDhhVwltWyktXrzWXtf5l+NXmlFKF/LzW5ddmHhCRL8nvaM14JnzXNSCyrmTSxfeg/a8
gIbNM9nnE9D8A7hZO02JUGbAKUKwbh6NaSLg/brXQwVxgnwjBt6JuGO2a0gzzALN1plHe3IdIodo
o/PScrATND947Clip8TnaXB13eC116TPwH5Rp16f/h6zy1QLZLgtJVCPC9ZjSbcKhJcsI+7rAxvK
Iv+GRQVCTcNNsDml8uGLsmnJnqqGvCQ87FVwlngvrMa174RaCpE+dG+9E1geD+kGLeW01ssu73Ab
PTKvXQNQP+0Bsa6Uz0Vy7UXltbd9lmxmG0Iq91m9pVImimGQu++O50N0oOudboMHmpH4dTwUFK+P
PEAYzQi4U7XHd0XBlGWdhI1K5YMoGp6civ8f0woYurv9oo0VQCxWt146MJcwhFe9JIQDaigJnBk8
mfdsK5BtCF+AplCR03t/68X8NP3g/wR/e+GkvFGH7Jxf788E4ZiSYgp7S/cCma/yjvG6OpH8j5Yv
NZhZs7qvINBFpk8ndHLzaVHC0Rd81bm4hsiDff1cNT8fJyjl79CXBjQRgMerwo5Zp4/gzykS+vG2
85u2NgjrO79DaGVPFUbmG5FiBlpodZZ7E067Uvj3CgKvtNhpsydNEXeqz5HpIzrI70ubZvRcBZVn
p2WmrQLBu1H46jteiiXWBiwawyBp8zY9F7gEICwXys05byVYHi3X5kQ1aeef3TM9JakgFYYuYKRj
olind1ZcSPHWA2euDXJHRPqQAq/xz3WtIxEsyM0zhC8gqTT9AQd9bQAhiNn5Fo8bRjtAwuIXOUMG
2CJuXxury3f/Q0n0u5DKmu6Qblgq2Ypuykk+GSVVTIGxAP/XAWN+O2Y8UH9RSzx1SZRBQGigL/Fi
MX40dTPy5wz31kD1MWRwIO/a0EURqsJvhq4FZReK6xo/JoF06qO7MTRf88yV5W1EgaIoBdDmuAAW
GtgPpQYGo6lVB0dXj/8X6aoH2HXejP0l2ub1KMMw3f7j817NZrgITNtJ1vOe3sAUskGM+Ri1LnmL
LCrS4jso7xiSFXU7UkTo5fpu7Ct2A2T7fEHigPL0hOxJhO3qmtA6nSeU2xc72cp/Q22S/TeJEUFO
Wi2sOe+ShYVgpypGWm4cU7PnRWCAaXP312DqiWzRSWOfBybhEnQUUx0z0LGdTksw581WEYtzcAY7
IeiywFN7igDGyahncIhAvNnQC/mP5sAFoy9/Spoq9kitxAjTdtpjbzrGA5j0oWS7+nbyv7O4BcqF
LNgp1CjsUeqqGoR+pFIyD+MMvKCCqa64JbvsV3YDFCuj7owYXFC46+G5edjWoMQZF81DK17ukKQ0
8nXS4qSeBxvBN/Svm9sF2XiAJgr9hp92sndNuIpC+5Di4E3dLelHdupZvAMpkplotioRyXVyvilV
/fEyfqtNJ3mSIqB/a/OsUpmC7uc6jX9aJuMZ6YbmoyqpFIOVKfTNAL09GjgLQ/xykCXzWQhe8o86
IYMeSBuX234Vj2xYwCgsVU3i1G7rfOJejziP/YLPzdwgqMj4Qu5VlP2xTns0Y5BufI55wQ3uUVHA
ZLs1wau5pVaQIimtF7xAC81Y+s68A8Q314xN2uMRr6SSZ2GzHAfmX95jQ9inCQe9rudpZSjTk290
q9vQhg0OF2/lKlAyK01LGgRBJ07/j0h3mP6c8mj/LRCqciEnT3KZxXal0ImrSJblumO/wW9k4/2e
9xt3imE/jsBRzfpMmo8j7fI9bMzTdXDkU4E/0vM4xdGdmKY0969UWfh8F0jsAZPmL+G7G1ysBgv+
i/a7p+UObFTA6h6X63SeIsOAvVyySQFaRAq22kxWNlMjTdVv2OpuFbsduU5YYYlukJUwNr2cFquX
TbDi8MzQoTJaWQ9mMRF7zFY9MchDetVokPalZwpiwADO86hoPDZpM5NZilZUCkPosU5EVciz5MQ4
1p4dmBxjmvwaadnCrJgqynbKnOAMkLpi8kMGg+uBM6zISHJ8e3f0pdP2pnN1a1tWVHgJOTApOUjK
affK6XSF2f+0dKleM649hIOzwOhKjdB2b/69Flih1lwEVj/99h0cVrZbHJXkKgfQjkhwbRl54sDA
UyD7mXc7G8uRFLIa4316tEnDXti8Iem3CZNohYts8I25go1kNlDzQQBaCQWK8VeNjAVhzeAbWBaD
bIpWuL6gABvO3wXzvZpSMEJAl7WB5Ts3mOhIeEEBPwkPhRqWn9S0VzDcqqNwIhhTdXTVHWMuvNkI
V9aA4dwv8nStjXoRtzPA2+chseIFSxG3RbnuCc3nHgMjjNBOOrYmsU+B/RAnZQJGKsJeDZXnuch3
zMux3fOg0PQi4BdFGnVp31ft60R3MNyINz/VVWW4xe3Nj/tCKIyjXX4M1waB4AodhE+ER8JotKrz
WQxoo1CfEpch27E8nq/pJRG2yoB0LcLFxv+pidSYHz5tniDRqwkBWfLw/pGJxRLM/vF6XgAUpSYj
1oQjq+Lm8Vw5ecsIFMcdSg+zf4iK95wTtS0z+DWcZkKYq3Xpjc5Awm4SyWxfcr5vFLSvCGWXdHqE
X9gVHLvTeGenwcKPvGK76d2pFquLyQrWln0R18UV/EuCcbKODvMu8y7xeoAc67w1WNi0cy91CEN8
VeQZFpfsuPkqg0lNC6hSCKViZUUj9q9wlHZWQ0OqICBTSJmQx+xHRJKnMVU66m2ndm4I3Tct2pvl
N2aQ19wVi6gbiRM0QiWpbMG7SWUkikKogPfUIB/0d3aG8hgzAc8iWH26i+saHnfmjjC7HUKTucXx
BgjFXkcphf/C0VYTZWJPxuF+AsKc/OPuN5BahKY3t8RvNx7aGX/9UWE3YlLj8lgPUVoIWqp6jZt5
WS3BVQ1WDyAgYLe35rur8JHiI+D7iuT74oi+zxwjVqvZlAYcWpfVY+J3uu8kPmKb2s8U2LCFYcdI
jn4fowvxMGXqaMJ5/U4CBLv2HoUa9zlbJZuHgGgUdVmgXJ65qEpag651TyT/SwmYxhrOQXq/BacO
TMlwK+dFhB1rDUTSaSGMsQUxauVwmH1ytYicv+lG3FAX8dHlvh5IOfR04g8V/36sotcVurDUO3Bp
r/Ex0+QsDhqk5n38QlGwz/iqmDRA2/RA6GwibMQPIvXhAhS6heddsr5876kUdvFQJo0ESkUQVnnn
HXiOpPzjeKeDrfLaMmaoOFxLZGlrtL30mOltVHTN2bjYzZNerfkHcnFVqx7eClACf3sU5Z83bVFw
LizK/p0ZjggxAS3fn0pG6ZcB4OSC8RXniq8PmEHl+HSLZzGKx5up94+EAoFznMPRO0YilSa7SAy7
WvkB/IuDwlQ8LPn4fZIOfdfJBmRu70odi8eb60Cw9dQeUcpJ4WR+B4ro4UoZm0YREjGqvfPrsOyt
3WVu1q7gVzChC/28WcbyEadklKMdPrDfGHnsnGjON/x9CH9jNnrWm7HnIPeKJv5Mxc0/qLrYjYMm
CmyYZHbccGCxhw2EK5Xm2rPsoSBq17cMSky1TA5tTKrx0OlcVvmvJvkLwIWqzOMFywf2DCiHBDYo
7ApeCLGrAy7ZT0IYFTVFZSHblG8bOV00pZpHWUQfru9EOq1h3oDFtsyOKWtQmtcsIB3T91QQRq9U
2igHzz4zEjkjSf/RGdFEZknZyZWC9OWaD2m656T6VQzUOvZvDfq+/UBz2TcMzb1KXUAblfpgdkCm
pwKw8gYrITWiYgcRls2grdingWTp4rqp563HjvD780C1PaN90ApyCm/sviRG/LqfJLOJAIE2tIYW
wN2NoulUJQMxZpmDioWtzwyJzmmhUCfEsQKPPiiKuV1huPd5a6KyaclHi8K4KxrUBCNUUerX2jch
YdLtVQAQN/tVLmjiCFAsj5ahpDThWA6jKh8hw0IqmstGsW8TJm6BJULW9bQwvXFb4GxPR8yGIeNR
d84uYZHhnLICFAtjwqg2+49Sew2IKpJPFuL8WCx79jB8lHeeJKJ4z8YIj2UD7mXVjwjPT6bRAJV5
LcwdonaGVwEaOsHL7Fv3SznL0hQ8+DiQR2xJt/IAQgp/yNRmbmiMPVnyCqoSGNJbWEf3TfrpakDq
MqfNmCW3fIbltzGIc0M2NDtmASO74Rd0ZW8wqg8h9/DuB8H667d1tX328IyIJTxQTiqzr2Gcl9Kz
SoryfMe+0zRgwniwNJA398zn3DARiFPtVr0Jn8mDwDieA8DIdy80i5LOzj4tkS7gM/JiT9h1c1UF
X+dlvHaDTLdSyNEfPIfeLkhRvsi3hs8vx+Jn4CCpbkW8206c6W+KIC7kJ9O5H5XGJ8xKzamJ2I8Q
XsyUx8JD2MTBBzVm3tjQN5cMUIQshFdpeqIJ3ZcQAhuDJvYB4A7rCppTEQbj8l+OuKK65jv9h8Ts
AqahbFCOQd0Zg47mDx3y3eRMdnbUQqLZehdpDy32mJmWZ6b3QR7E5g/jrLdeKAxHt9XPRhBrXbY6
XE1ikJlupoFFj81QUDgpV55jLDSgjl4mY35atTdrwnaGB/fZKsIxr02ujwqyEDvI6Gg7tFgijPfm
XOy7JxvqAHuiJ7IdkzrGxrSZ/nl+XryJXIUSUEjWCdhnhJl8Q3ex7kIn6dYy+ZvkhoC1+5F1OvDp
bWZj9wNQspWprjEGc0s2NqMvk3LP6VduK0yrYT+TJadOySbETxxiyyUddM/cpcy2va4HDxzEjgRh
w3/oCNcmA4OBG71DmtgmqqspkyCDY1vy2QFO/Sh8mCd+TnJd1FKbX/rqUj4uZj/ry9Py4Vn7RdrD
gz5aODT7sLzGzKH9rsXEekVRPwEW0OIG05WqLiVmT9XuAs5rbk+51MhbW42BPUlEfrp94t/gn16A
Yb/Ma8IHx2Dov4TIuyTn5eue5uF/fZFyNQZ62Mgg9jD5+XHoK4hGpcZ++iGXki8kDjVJu/crYX5A
yejnDZx/SwzdKruaiAeZe1hdjY2USJ4931H/x0RgFWvkioGQE1Ki8es8gs8pHG3wNJR+r5VJTRPc
cnyitXhLBTGapEvrQcn9FzYT6G/x/rbY2Oj1uy7NPBSf2PBuulABJOjIBY1PNPB3cyblXTHmax3I
PkGO+mBWUx4prGM2QHM92o047mtDCIoGB7+2Lpr2cAbpByfDwtsVL9plCkf+XoUFqqmt4OlrepA2
Mftitp8pXumE5XLFZVeLjXSIBnuaYSHljQUfTlVqdjd3cM2OjAmwIRKb+IFODDD7uGCCHmav61rj
F8TzYH6L6UWpwmdWqFeE8dYO/CEY+kymFLjRF6tM1SuMVlBx8IlZ+y9QfsdeDwZeDoNn625fhBZZ
t4SUxHoPOZiW2O5oHtx4JhAz1mj9yzYMNuFP2SPUtnhjQ/d4fNp5H/ktjvOwzg3TiESov7wYD9VN
O1MslfqcaCIbvHvclqUiJjlvBufawds5tyTKsxDlb9w1vGzgzWHq8Tg6t304QLmDV9cCFlAanV9d
/RwqbguwgliD9OIqcFl4Fg7iitCUtOhIZFfCYW4saFNbdeUjRk3OT4OBGjOoEVltKm1OamNCGbqm
VC+6VxaQibM92rYSZWVGCkOQ/i/CRrhscqvwUYKfAMp5cRWHmgQPGIiWIdPckxLCPIaG4qgzLh3d
Itf+sX9aarYk+fhtAOpcYz/T1zWXIytliVtgEG+kWiiMTTikH8Vfa7v8HelDYCTzwZ0m2dP7jhh1
GZZeqzT0Zpm05BpDeiDZ42VCSBjeyLqVyTfy4sbUsRQm1J8rdUsBj895ZclAEb/MnbbcrW1nqLUw
0lWiJY7RwhXp+P99g9BM4H7mvmKYZwErw/cY7epmM5+Xn4EN2XJicZKh7M6MOTNPLiQYAM4bTtPO
1zsurALxVequs0jGhOgE+hCPRg0E0yQ5CIs+YsfXE9l+QJ9P/urfkhVVC/5cP+mjVauoO0WWd4wG
hxtImeqsbhe93npvb1PhXMEIg3GKsfEGHRDuT6nR+9F2NzMDvbueDz/aiwLOGQUlLi80iMJ2cnlw
thiUOpFOYIPT3xTdJFjx7zADDSQtQdwCZ1lB3UGpGoh3Yo0aew9PiTFuE2hxB4LJ9QudR0qJxLY1
Ozhe3rFVx03Q+pe0CbajO/1Td62XCrKIFvBorJFAtBdrHR4KFkSVWvpYYENwpSfZRuGVxKcCqKhN
W0lrI+73ZbBSnE42I6jD6mP/Q/75ppXeR3fcdEkL2rXQ7DeBUO6qbXqlpyfOFJ1u13QmnGif2i8B
DKKNP/GpcNNgh6ZbMvq7ivnq0t479GiCckNrO1VJ5C+Vm6nzZWPq913bZGB2X6OoKK1ePbybJs2q
UvwstxjlbDY700yjBxMgGZZlC4pkP81lpx23K3PVlJg3M+2SQ+F8frUSzkKPWwPwd/dtEEG+3iUC
1dmFQzhWZAUDXAsQRuI1y+dRFpah513sg50+DFFTvxQnLEA6RtO+8pIUmdOh4DlRs7Iz9j9ziyqt
2WAqgtnOdjwbYZ+IsFE5fgPTToT/mt0Whr2FhZIbSAIuEZd/r2N/+yxFPN8P1OEIzns9pZeI3oVq
WTbmsxkj+ZakSByKmCYtp6tiqU+eKBAXI/lnsylXsI2PNAEogoLea0kZHFW2jj6S3x5xoVYtOolb
7tS1DhI+i32/ka/NaYuk7qJESWsbU4oo1p8aLSMWTzSrPqqUQF6loNTh8cBGdrSlS+wnJp+ySO5k
zXL9XkxURtY8bZeHbgaTepTotl9jRJybT8/xp8TWWnbtenK45DleQtUjbq9RBUFZzmTF5ZRvlz6S
7BgH+UoujqcbA5kYvgATfj9zmtXHNBXZQjSOPJWY1EFAqXbQilD5qqZ2kJxOixidJYW9lv93BRWc
4dDBn34M810PSKLjcwDBfDt14s3hYyRvL7MxA5LA9oMNY7K6kfmhOABCXPbS5DErpsiwzpvnq+YX
cjyJeYpVcF212iWhYNdsdUvRgCs9zsJxTK+RYPBu5qJiHo9C4yNsrNybtjv23/CG8EZopPc0ImhN
QDp4y2xaRYTDTb7i3VwApX4w9PD6top9bXAib/yLjN9BD4b5xag1fSe5X0uOk3vEwpluOVOM6yQ8
tTxl8BycpkCbTq5ropZMoDZiUIA2sI8ACbjuiMP/5SltLhy7gmuwdWuUrgUnB+czB1gRmWwzpanu
YWUsgv0109bjZlRRmtW8/+zss88ZTMvUnTs4WaGzqrbm8KrZvw5PQxwQW9Yq3Fq8DAc6W57z3qLV
KfDQS6IKmPii5C+YCMZnsJ62G5qLtY46ksNe7UPQeR1X+MHx4v/trnpAQzA/2pjQJ3e06CCcTiOv
godxcn394cCDVAnAOcO7RP3YCURAjW2qYCma4yKr2ivm+xEy9kLeoqT3+VlZ3VU+Vg0FlK3g+zNB
OE5dQToK9NKdhGJgY1yJBJ7JQo7mvbCfBPVRLlhNNjSFGinjut44X0ilyYbQ2VsvB7zFdyZAMXLb
+3Kzu1nHgfofiK7ynTwoqzJM3U/j7zbr+sxrgL0RT0aaR2Uc071P1QzJ+8Vmlr2NnsUFKEpjorU/
BMXjKYprbsCLv4WCHP41BP/KMk7YDgoUc2crplBmKXn2niu+iOSk5fg7IwpMqLTSEgtd8IbAmz1D
6XliShNYjEpk1pp66qyeVAWI8r0Wifaehz6iaWzYritlIK5pce3uBSJR+lQgku+aGclZ4f4e63eQ
QbM6id7shszw0RHSDNETYoqkf874fs3kdWFulVadktPUP69sIuYT1JP3djinwO67ezrWWgw2F7Wf
OaCVcxUIxpdxu429AZhQ/i1fCAhCY9AELjrsUCGmhe9NAmbpmOP9CieHaU4VmPjL6lbofJUKkAcr
XvT+PESgJDvE8BODwJkp575OhXI3JTEu7Yf30cYN+bWIgRpdU174gQ5Z5Zr7h1HLvM+4wsP7H1Uo
1r65xyQUMAX0h7chWDgzsl3sv9PrSI9j4+OVEe+BTWEYoti/lUhzXsaHoeqpru/+JM6zA2BQInUs
H9xrVVNc/xhGRr2Y8M2Jv6cAS3qoQ/x8LDuSGUYq6nezK5skzpFXzF11YGsF7eXVvfqZqgrrh+BN
EjFhyGB4FYbwyvrrV4SwoLoCBVWiHQde/EVJRbQJq1NtfSrUSOt+hb9dGPWYUoelduPNfj91q5Kd
cc/+xXUCz2lamlppUy879y1TxKF/EMYnBVNCUBWTM1qnQFbHCPMzZoU+6TwATRRG0midM5RiCfgM
wt5O4PdOsejzPL6tCtbEIEDY0jUH0XjmmyrlnMVE9pRdIQFfLyIhd/Ytps/HnfnD4ZrlfcNnFgoB
Utg2pjfIHOd8RZTSuJUojoTGF3ICWWwRRoCrZxAuTnPApGVpRv7w0ceADeX6RBDrwfv2SvzhQzJ4
UWaCcurFjJm2j+lnA8AvF2IS91IX4iAowld1mAy2Nf2IVyHSjnVBt78BzChPx4c0ZThwRTGlHjpi
/CX5qc+t54F1l3G3bi5dhiBfRyirmrEG/MeqOfOOxW4QRK+wdLWj9nc18x3AGv+CI3YKiE8qsKL2
X4s3Voo0LPWpnXBcNkJwtFkr1MT9jERciz8TUppLDGvcmT/xZ2gtkzjVxEFObakerJhOWvyPh54M
szF1lXqF3+rnxwNJGRHrARxIh9OB7+nVpQt1m8r8XVO6/r5oTz9jV1SIPu3p6t53+5aMp43Qe3ai
0zOGMssYYojyA0HxQPg7ghSpv3o4bPplVE/D1A6cupNKbe4gQsH+pSVvgPpwUr4yitFZELbzNS/s
Kw4Ld9neVpwZiJRzLyy/6UT2oJGfyzPUbbRFodiGn+LrG9OYJ8GDhpRkNcbUU+5UFrnYeLwyLTVa
L3gmIPsDloBoxZb92+/dxxPtbIlqbShQ2LfFzY4NKwIbgQDZEkgUoi9Tmt/N61ersNSYgXcIkWH4
23Q/RY7w3Yg4fHBGwN54GKvkOhyRNBGq0Q5xA3sMcHrXD9B/J5NdTcfIdWHfKW8N6coEpUj3Vw4c
84dGO57Zr+3rtghzvJhgqGakZfaubKFpll6zbWxIjRELubw90FxKvqMOqZEAwrDqJcuQ75WW2GiO
VhDrjuyPUzrqxr1gUmngCnL5qLGtuKbOpDYqbhnTYDjBPkJmr1A89ZLm86JQjMXJqJyv52vhpGYG
3lLBuZkMuRIpl2IkH1U7j+0vqv6zxbywp9YJxh8EeCCS9dR/HbcO3W12MZzif2GnKiTEjbuq7NQi
o/9ERHGESA/G4P7+mKUfcTLwZk4S1Te3MTZs3MOqHBc1O/woBsHDUNCtqZ+ff4TZ080OKfdvOOFq
IJCzi62WE1ORCJ2ygy/DgvluJWWpNPu/g2/bk01TaKQ0YNI/MSlfdFGVpSeafV4wlnSyKUFyCDy2
iWvwH6XOW1+14iyBkpj4r/EGpHS3xttSTzWuPbqr2fKuTFHddW5Z/3p1Ntk+WqHTlyvZTKpRJJXm
FnrRnuIDN+PKgpA2DZWa9z+P4vYHxUl435POEb+Z2eCY0Bamc1Sn+rRMLbGuS1x2L71ANoJHBODd
CdDWDLrMSZgyYYr7JFW22LGhd0vvW4QyrTlr6+kuRto518U3Ibhu66DY6n147VPm2yCjDwkDHDPj
yQ2s4CoqdI9NoRdQV1p/g4S0Fp4w+/E4a8bLjYzAKtULZ1VfcJl4nDmUVuO7flEzqFO1dFMVF2zz
w8zT89s9/WfvX1OqPvSoPFAC1yYnCHqCzXrM0FIW8/jAg+yQ5X7nh9R37PJeueiZ/wxBKLwOW0My
2sswP6SqEs216W/LllIYPmOmrGLPfuZsRD+p0cYbJIcQRatSRAHw3Yw/ZQS27Queiv4wob+Ofd2x
bYnRACil1LN4P8UU22SIQZhc9CPrHeA2JwO6U7imw1GtzpsevboQRbycjnHiTfbDnoqV3zgHZmDJ
EvkVbviQF7lpVKZuujX2hCeYXVsU8DSy0QNFDkC9HOA6iqOi/GiAA6XXV9T9ByEVStkAFiUkQwDz
UNxvXmA2AZGj1q5oMmmVou2pIiRQMLE0BvXihvv1ZIt7nn4Nfr3HpsTvnv0rxWMWtLNtl74aeMZP
sLt1cmvbDxq76+mLc5grKMqPgpPzSdEA0uL89noYPHqFidujRzTjw92eW8gfTr1oTGtsdv9sNhOJ
th2tfQhKgF0ACZSCwcNFzYi1Sqw5j40WAXYUsuk7VF2Jjk12/WpoD0FzE0wHsb8J9vc8PbuxDwOL
AxEMPBNxs7zkXCcL3tfBdvhMLDsxRsTR6U6bbIWP7JN+CtTPwPytEwQt3Cdg+ZPAZukgdkiZYZ10
4PhBp0QW48Kt3VHbJJQOa8sVZI5UqG3iA+X4QfuNngSkqe+ZbfYY2Sx0Pdyq7azpsP4UvMyaUNjV
Ad8VgB/oOI01/rKS5iahlZjD7V76riCM7yoyon4yk0rMzEbNcM636BucW0eafdZKomoIg0jIrPZc
yw+PI+uCtS1dcIDiroZF7Rx/fdFoamdhSb/MeeQqjmv99zTCQq9/jQgAKSH6xtd/yCj8V42XlDM+
rhZNKvK1VvvnH2kcCcvIUp/9lxPzFJD4mCXHFY3Rw7v7fLLBH34F6vtAkLXR6D5rGoAjQcU4wIcd
UtRbJcMalPodAOcxGBQ63XdfgHwKrDhuY6bMkZLS5FOkTDB3V2T+RCIOEG3PUwLuZGs9nSQSltn2
G7dn4QtjWKmmIpGyw+j2mNUys8YeQtJBAgGf+Dba5NJSWb6o5qYe6OkUrVr20ycOtSjrcCkHgXmX
zJ0E+Lesm+6fdSC73dsfjMaWbKKxLnUabpF+ZW78wtFpQHYbr0y7eDU0DQZgekwyTHpIymw0BJCv
+MpbvUxcQcF++6apH0dOq1fqXCWgZBYxXVcWBlSLC8ZE+XWXvlQE1eXU0EldWP0ETHHOTfk5h3un
ELPZSRvQcyPuMAG3qnGY9P8kvGRj2ZwtFFVGIsViQfdjykdFeCCpPQJV4HoEuuwidh92VvK4+Sr2
6gqHOHlWO2EGXN2RwuNuiHWHP7D9wm2MRSfBwAcXQwnHIcG0I0PlZrSN0mUfiHKaN52NocSrIJYK
q8G97yU1LuPT2bQSkHqSu6GIc2vvqJIC1T1YzUQtCeQqtHqb4IuArnovTa4lT1cJvSyBzE1YNmYd
BdAojsUaSc9fh8mHpQqjgSt1yuxlp8JuYU4ATg6TrlrZcIiw35fmTnCc05z1ZvYDCReQokRBQ7NB
XkPyYxJp5jm1gPdxwgg2VGOVd0vdIsqg6FUAf2e5SGRhFHrhHRd/jZKYVcfn583Rj4DvSmCCS3mv
j6AWcJPH88wMn46Rwq68HjxxsPx3Hp3z4+KjO1GhqMvrp7D5GUC1RVZ/KIwBLmJx9YgcdtbkcdM3
19r0aWB5VMSN/hY2r4Em+aBukDbD8P1RGb4XMsw0K5qLnxx5NlhO2fd02wWNzejJ5Za/99pruUoD
XyDi9j0UMa5JCU2GtZsGGCYbiJ6cRbbHNOeLSEsikSZlfVgdgKzArYxgsUZgd8aPYT/YuHBj4WrW
yRdb6bAU04wT5hAatZpGsBc5MI88ZXsSGTGuPLsUV0CmYxSlsZC7iK59ohSP5ehjo8BVu7jCGThZ
/ENvhou9u3BFtmIVRXmFsyW8/8sKPnQ356SdckkanqA79ASIk8mgCM5vXU0YeLQOK7i7JVMXkz20
Nxx3HKe1kro6BR4T7rTmuLDo69M1wtC2k65iL3EcSTEO1/ajatfWd57gIrb/941eJ1hTlaQiHPtG
0AuwrQ6Fq+i0YaiF3ajmnJrwmsCIe3z5Hjh4HB5xdVWwXTQLD26oIZ/SeZtHtuo9CKHmR5aVKn+/
xsNeTv12Nl9ihwX3HkCIF5mRECFkvQlfQWkC7urt7kGJMP6EHMaz5gydoiVG6CdQihRIFP49GUYE
YigZjoKFnrp4fOzyC3ZsYXPbE6ZFvpc63W3opTtAS0MjQFxy3vcNNQbVEynW30zMfEmLrn0dcIqU
MTHg3Nx21S+3ERocFJhzRC10ohJeDpxWtY/59jgL+LPFB3gEgcVkVgvItkc9Db2ZD8wZDM0dsIyp
NpWtUJWmITnNrULZiFKpRSk88GJ4s0Mc9clUdPpPsstcAYO+x9cJnjtyTie1HwDkztx6WuIssVUz
BFsxoUhoZ64kYoW7SAS7zIAwaL/+g9yl2bK7AxQrXOIft9GqOm3LcLeytlLyQVybqxcvaM1hk8Ed
o2WpU+PYQRwkvX9ZH9pCyo1qHGek4JshZOmSafBbAcrDJu7A8XS9uBkQtuij1AYZXY98Qy/Z1W4I
3zSIELAEa2Mpv8kLLEiqr07wX1lvMr7dKCtzs3+IQoZfa89NcDsYbD7MYk6d5JO9BlrKKCELC+KE
o6oqh4xw99NMq63SxvmMOXNVeHO8fmd26U9vTC9OWZhlYBIwsEJ51PQi6+BFIWUUCgfBTzwohv/w
Itv3oCXQPp+RkoRd+HbeDrRabttTwWapG8yqM3LZO0fuvkIc4acqNWhTWBPHg6i9nXV0NXmnzjL3
5jwIA1P1zqj/YUT6Q9LMwtMOz4upfPGRR4/lDct9ujhx0P4/MnT8C5p5idM5P27rMvmmm7wvrZwj
7GZjB4dAYFnWkSWljOZ+7jlQ0J5NSe3nRRnIEkAuJXF/t9X7Z7AGhX4HFFmcUZjgw6leyWw+3FiA
5U05OT2FtoUocvyRaoaqJOn8H5b62bbE05hSG4pGL9+0/i9lXQhSieMopvb8nJhtXae/pv/DN4Lr
e1ouuHyFGlCfEKLtlNyxcfAyopICv/onn3XdDZ85gY+dhnfCIO60IRiJHP3ikeG+vnnPctE37nxK
1NmN8Y3BKhphW7c8HM723Ldrb2P78yzp9uvT+l/AueRTdtZOxLEDBKBtMsjIa8zD8yHZXjSSilD2
z55Hk1qp/3Yps1xjb7dAABj9mKBmpegt13cXI1R/UU+3Yc4nTmbbv48i9vP9iCtwMmROL6y+XTH/
Y2d09IubmVJAM2gEH6LsNY0ekih/btNL1Uq9dYEvNhfOu2FfZMya8KmDSW/8cSTK9R+y/7UUYrE5
WDR3iDw495/rCPCEar5zj0oyolCmDLPur7E62S8wUX9hkoYovDxOlgkfFhLX4vznryUgztRlovLl
rFxFaPletlN4DTABCxLNwwOr8Dk/vzjIjRWuhI1NgDc5cylJslET/cJTkk7f0zdF0Dta9XGtkklB
M+T/UQh9+hM4HotgaMkDMOnq/PhMiAA1nqt3MoAKaaNkqOjYatmXxQVaAwy8FXdhQ4D4xfY0fiUK
nzp3YdStBT0+r/34Vk/BtazljE48CHLFn5GZU4rCz+ZVgiG0lpHE7DyCpwqyHEPLh8xGyw/na07a
dY/329kmS1MZ9EySLlhOnM55CRAga6KV0m7wJOCHXIsuSMdtYls6iY6NGtBm2fygnz4l/tDcyIB4
cWUR+rrJdRMEQqyGLQmSokA4sk92CFwQM93oSRL6DjO5D7eRfrJ6ev+F49IandP+tBE7ueE/1jA2
ggT93gtBNjiHwcBiVG5EodbCerqg3GgQsBMxjE6PYoob2zNnDLg5NRbSVw22aJo77T1NEG8cK2bk
86IQX0OrXOlJS8KOIrqL5lV5VLm+ENWZ3zlHroEqYtrZKL94IPD2J0dnA4jN2uEf0hyumU2JZ1lv
sciqODG+D/rnNdb0Sgg5k4JJtoKsWfa7c9pu3VDqgkZXDb1hK4G+Fs9GXJaozLZyA18cVpGLGDVi
64s5Ahmx3aZn7tvty2EH1t54gpSq59vUgVCUddjXDA73ki/+1nh2ZaurKAderiTfs8NAUWSR+NfE
nXsP36Uibfh9KPZr2+oJsaMWWggCOSyG2n3o2rdzoAG/7yywE2yYWF+GRrxNZ3I7pFkwvaalzp/l
O0gni2EFyMNdU1a5g/2gfw6cGpaPGBq/mwoDv1RYc6t46Ig3RwcbmikoLL4yyYfMAMtIeP47hpEA
eglEbh5iIiwTFi4Fp0vN7H83MYqy/1h5EZKqC/hUPllcsRYj8r/z1mk4mJgrL/vDWt0Qs99sFn7q
C8UmhvfOD0Z51szaT9+Jw2xZUT1I3Sp7nktNxAO2gvVAWEo5f+p99jBSa0STc9BBKirrrXQMgHSw
ibf2LNJbV2fbr82ClOFgYI0Dp8XmYPC98Msp02/dd4hHdG/49nPY0Ba2pei9C10TIqM1zDyIi4/1
rL8MoP8KqbhziNW+wn21wqv8N48vBAuSVYb1kOJXQE/nExxd/6yYvXS8I2vd7qGulzDQTBQqJWwl
1Wsvvjp2/68aWt/FxQ0wivdNE6AYE9ta5l+a4eHadJ0FuLI6Le0moCGoPyXWARLVb0R0eT+NJdS9
kcT/m0NdWLKA6KX4ufQ0DRNddQ7GUKu8kHznQWvMd84oQu4OClwiiidGlXCpSNFosq+P6IDalTaI
ygZX2D0m7oU4F7hPd79Aq9OJGbBlPFnTVEZrNXIH+J39FK8Tlp3FksqexxxZgKsZPEacVlggt90J
CbS4hzsu96OFMcNE46pNYw29cM1AczZnHAKmyfrkBTmdclAfUcLe7KgQ1G6NHRTH/0lRaCPcU3/0
wlntFOjtCBaotLHuAa4PDUNfFpuL35KQ3ihlOsawdqlEuSWF0uZyCB/4HR+oYH19cYCcIOOb9Ecs
PiQMAeNLHfnBJ6QTsQKPkO7hjpCQEMHdzvjVcvAiJJqkuva9UB1OxieNIPtjwKY40DyqOMla+Tbc
aMnRgU+wm8TX3dA14qHyRAKxIidhVvytbl4nM3eYBZpbH3JEx9pbW53iRsrIJkVmQVK+EQKzIR9H
dGKvgLs8ZMOaBClN6bml1tmRB/lmpTQSp+RNleDRzjHDwuzOCkODQKK5d0Fzia+bogltGwBL+K5H
OlOI0iuEwJ6q75UmjY3RopfosA/3qPHVDYLeh/SWd2wxUBcQruyly9klyL9j9hjvU6yRrmuhrouE
i4u45cTE5M0fuh+Kwgo7P7pHRoALyu7A1lHZy7yGGwEDM3Zl1YalZI/sinDQBko2tJaZ4eJU8Uwk
HBXC8PICS62eW0JaKkXglgNmCbcYl9OVlF5Mm6effAsDkPp3aIbY31bfwPyFRmTQVEAVT1KvDYoK
BYV4nU6FWqLdxxDGZTEzWQX7IKXOfP3EXBSBZoL45ksbvzhs4eU4cQQ8huWFplbkskEo57CpHNr6
7bhWTPk95tgDoYBHXGoBynnevA6cX7EZ7Xaqo0Iqsk/WPvHfDLu64OLTzGXMawTrWhmcVSldqHc8
/cj94GJ1fvyqkL0a5NrIWKzlIIP1EMobIBq6fiBkN0IZEcvNaFJnm2TWY57TCms/M4WnWrOi9NMv
8iPS/l3RsBoaS0qP3sE3qumnVBCNjFKbAfilU9EYM7jFm3q18ES+8uitzOjUsFsYWK9qWgVdrRxl
8jBbSYNUcDNca4+CZkXdUWtybF96RTjAIagdIqb10E+5BinlYcX6WhFl2rmMpd1d6cNLY7lO5N0X
/PvOCREcDL99fc+HWA+Gcwu+wYy73nQrHRUN9TSDQumAvLxM+f5dorW5CVi00AgGRJaraJ2pppXz
Hfq4i5OvGpCwmWcXM6hKpzTft0ZtVM3yI2VgnKMzAKbx1zUAjBCKBK9Z5S2kWhFumNJcQ9LNCAX6
TwY9kx1bL/84wFFFvbh6SSNUL53MFoDOGuJVr56BphZj1NLL/aBnSFCeZJTGhOqizicpzMPBfFks
B2sAlFxZw+noqpotgynB54C3GH12i40UYYKnUlfwKpHZFUWqUQzzNOcN2+xG3o5qUpV8VsVQTqfi
00DlkH+Qf6FNs+pwM9x9+g6UjWAiR7HNp+nJWYRvdFyhIc2d8IKLKxmk7Pd74uc3WVhwN0vA29Fd
ozBQoYtF7oR8b4ArdiTOxOW2B5hXcuNj3q33s3b9LZfOOotPPNtYx7jJNeWP8B+WoldFfVxnoKV8
JIT1bbYRE9IagmUgOGHrv9ns/gJqFpfa2UCvAJiLEM6zNjHpIbnoK/004lIcp9MDEDvF/Hqu7WYr
fKjPVfTAZlL3TO7mBq/12DgnSjbjpEroGbwOdhWeM0lNqAmkc/EeFZ0JGt66gmgfIoWiNPMZRyc0
HBmVDLiGivzHUU+FRF95Dhdg2wjNoA5TWseOgaZJGB0i/LaZ8ecCSmjnCEam2b4WldWmyjWzBY4m
PtrbbKNrz23Mz7JKTfOVlHZs+Bxn09Noh4LuXr0iyR/Mqt9/VTbDxkBB76oUXkwgAh6gPpQgO56y
/TfrQd9KHRonsWE9dYQPIQy4rSZZVtoPUqFiQbVmTVZA4TXbnE13QRGVp6Y1W384z1GZRwpY0cK7
WGW7w1v1pq6q9e0HnfSNCG6kgT+IJyziSH9G2dCNB2Ja7MzRuyYFyzZ8RQNm8ev05Yh6lRbfhBqJ
/TCIFNiieypbdsQhyIBjwkiYZhY7VkhCDCCvp3miGIuvCLF7MV1fVp+AAQoTGd04EQnuv9kJus67
TyzwkVbnNAnQQW4eRz/swKg/7GJo/ghJKKKByabpHVxJV9lvfp79a/oWKmwpuBZdSaBZoWXQxvv/
98s7nZOmxl7cZCOpV6K1MriWvGMefmSe45R5RnRg5c+dfG8Hl/suiKiqSlFSmtrT/pF93J9ENfhO
nU5JafrCn2q0zQlxdfc+1dXRM5GRSHoEadnFqrwG2TtC/SEN0u8S5ROqkv1gPM+DtmXIRItqnr5H
WAWWS0sMmyc8cl2cf4DqUt81iueC+Qa7pNVijhmLQS5dUoQOiVivO0Oh/s9w1guKTvrNXuhrpd6r
3y8xzmeX44k1bEc9iyql2rCYR0tVkDjVWsdaicB6apHUzShQ2lnZt4+QTdWkwy4C8kT2vNsZ4S72
G9eZuicdkOXH351P/m6BCw5Mk1kPue0Uu9qSPLEox+zhGJBAMVC1JZhCnXX1oxAwOiJIVmZ8gqVu
pmqXQJ3F569pnJlksm7faL/zK415G99sEAAR6L8hgu3dqQtC8l+qhfE4HEQNXftNajOR/j/BFYDJ
dsQCx2oeG4NYS8YRM0ONi0Ce392i9zOCL/ST9cZElWaf5/sD4d/osQOW+lPGqdKw8KCCEQkBgSEt
CQVKos2NkrTRmxRA/SgrNu1uy5HGPjXZE5vWuTaQ6bBZLXTGg7/bcy+3lWxdo7iK1laQurRo89QJ
oQbWGqafFkHXFNLbUeOAAjCGrvC+W6dFSsE5G3NIkn8EpmV050Lb6r70y8GUwxhN9JG+g9Leeybd
e0Jv6knL1xyeuMAMyBXmb56b170eLiis74O8AJvbiCmT55k0wyCeDFhu6A9qjbYG2HL4bbBxuYoN
WuTntybSaD/t1apulBneY9nRxIPImuB8A+C9Ae9Zr8bDq+CGAXN0KlMEv+hNRrnAqK4FoJjYglWL
rNOQhCMs+jBjlntpyMkuyPwZvvAoqUC8GH5clWZXhIxjuic7z6qdA7TORlrBnIjz+b58JSXwmgUn
Pcf/So3BZJAeHyBQhnfW8R5/1f0zeHzyMLCF+7i2n1/rwxtYcTG31sfbuDhE6+wz63XbLoXsoA7c
KBPbU8g0WN5dbBzzNPaSk25FkvY7E4hD0iXFHLvGRrnGean2VzMd72v2ZyDi02aVHV5XreI72Gnc
3mqccvdT0f3tAu0X5ZKNlQKDBO7S5BlZg6Y33t9wyj4UuDnAReafvQ6Z0+jnvuovMceaH/aNlxK3
GSHH73YMA2L+KXXUsIm7Yn318qDvItEBU3txLan1sdjJ4rdQYZ29QNVD96zOo8mDFHRfCdqE2eWK
BcMJKbmTWgIUbK2IdXNggEHXmbtHyypg7/S+M9gtCM3yaldssU9i5HE4oGiau4kKtyGcKU+dD8bn
b54lROu2RfzUcRGA/0qS+GxBLqk5/qlIBu9N3GmD+xZHM55dmUDZhyXQdrpiOKSRdzvOBZuKYUjE
UPtkkinFeQIaUlW4ABgTFbo/N2y1rwyl4R9qRbDZuXL5JPblfcbJDrlZMcXcNO9YCzqfTl9ds2O7
wtPIS6TFL4BI4L4wMpzLdEm6e6/77MAldsnwvrhj2+MLUU1Evq7Sk6bgUEsQjpc8ONz9/GY2wgyG
gLe5Te4FrkvLR20n+o8ON4h5kAGasx4tc4rkGB++BdoltbDB/iJwyc3NRs/Kop1I4nlHjZffwWYH
SiT2PZuOfvuKCf/p2oiPGLCbRgNBISPdxDYndiFBZ9FksAjhjY2E6/OipfzZG6V8brWShjrOGRQl
4Mu9X4Ex902aEbFaE2k1AUnRqtyqE66JHvTiansvyLCsPJAeyj7qBoIBM8rDW3ljcr+4ktlYwlvL
cUXN8PBfVB1lXgwjr2f8rCD3T2fHhHP0p9Wvwbz+uKSG5T2QexBQsGvv5yfRKXMWOeHTuBxxbK/P
ZkQ9jOg1IpzLRbkU0EP8eXE1Cru+jfciejVjB3sjDQEN12wAacqQYZVavDK4oCapKJzGYTsQAiU1
gQtnOZtwUMoTLbPlT9tT+qOKVflkIpN+WppQ4HQq2JdwZXElDC9pBe+KjG5PmXDwrI+uF8w2QAVM
yPJxQ18l+q0S0kpDxfafYize8GCJ/utyBRxFc+VZtY3PS7xI5HvHzBhiR38VRPjWV8rFMEbSj21k
R9mP4AYFEBvyAuS0FuCRRTRmIT75RQZzDD9S+NUFnLMKL4FKiUDtOHOH5tl++/8g4eelVztZR5hQ
RAD/r3O+lm8aLnu3ixQLq7we6aXwVJVsjbC9RajZ/EhU20PM+m3ljeKjfYKlpbFhzkyqKG1TBDS4
JjmmurxVDsNEJeXDFLaN/2hsopD+7Yc0ruq3wyft3KxUv3ye9QtbJcAPOGX1DZpXmlLECgABrwdb
Q0o5dYOvCB7RyrBhdVFywRp4Z1ibTq6IaDrQSLpXPLcT/weg7T4rod1X6oG/4B04+A//bHYblhMk
dN2w90UAFnNcIHo/+IRBSjkbKjJe/EicRlP+0LBZjSnva6QrwhbRuHeyR1jpXyPxxed7EmAvSQPi
N5Ls8ctkUGF0rG7KnDPimt9Si/rLZxUwGs7ZdAvYUXix6kCOh+9WSMmPCJpQpvoFYgB2wSzCtqGz
qKLPUFZiml7ya8/33qmYDbO5UkAFQF2aVyR1eB5+YOHHf05EatRtv1zLEaf37FlRRPXsGHPQuT/p
KTD5B/xcAC9M2luou/bZoqK7RTCNj1yR8srJp+EExPbdQ/CoP+fR2IVHL7fUOcPNB9QpFLCV/1j0
BN4dfssHNFMsHEXR6bHc/6493QQV2u4WX+d46hDgQ5dr5Fgb8IkjdXrFLsqaS74p1a+2ESVfHgn9
p7BIdwBuJhxR9/fav/yz6G2gOdDi86VpzAOt8F4rcLhqbyA39lZiLqKg5SVFLnnM/xiG/VMza4Nl
Mg1eWENQfRgU+HzQ7Jhk52FWjRgStvGUqKyHiFMTi7EkZJ8SCFgWcqtYDIMnTG1lgcCAWzBSOKU4
9PvE1AhA4hsdtNZLlW8lzsiCvtgsQoKuOMfKGfSbTM3IRrcAAb1fI1iiM9Hvu6k/M+0oUod5z6Hb
t77CTFB9f+WEuK9IC8X/yXgzWrImDmpOhGYMoHTxUqq/xr6iBHTIIfW4tHqJBVKKFSrMo4b3k+g0
THnPwV7YHbYVRX2Trsdt0Tbr6ipXFQvCpZ09wtIAvpJkknEHyGfCJ0J2ELeMfhUwjK2AJp+mFvFA
XlwHpZAuE7Hr5I2Z14v+GYo0BT6nASRImfJ3YIz3xZY1LU74yeHP0DFqNoEEeG1zQoPOnLK1tGMU
kDgh8ewStGVOq9OZ6gfzGwfDtTxatA5tI7o17t0v9Bw9INjHsgmUIGwzNPzhKElMWGlTKXz1BGPd
l0ocBe39VuARMzh3BcOO/zM8pfuRBF6/ZqfCO+43hRuvvr8vYUp9aKadeGVED69E1CE36i3qbFIe
rcT9n0oU4r7qQYm8wOmCiEZKKdaEJu1Yuwnpf5ORe3LDXcZqNEcfAHuHDl0ZFZOHoL544ncsyubv
SNtS+SZHWuogIVk5uJTQ7XPXh8h0Qz0pI603+tVD4Lwv7906dnpBHW25ArveFbxWP45tdegsM0D2
Is/gw5XvXExJikYjoCejR4IPw358a3d1t0bDBR+W4S/rs2VErFsONfWv0Kpck+mpeujRrXXKVLbe
U+SFTthBX6X0ocyZW9D+m8n7RiYrtSclcYunNJgGFW9nSu8qhl8XG90pzMETPfVymMaZNUNGPwgr
bQJ7sptdIRMauRXTt4YU/a+GLOkxc2EKcusxA123TZn2D9aT6EPBgSblnpZ2ZLDJ9OFXG9+v6KTW
sUrVJk2ZX6mEfp2YwM1DACgcUMD8TShU9Xv+vgfWh9PiL6C4Kjtf7SdAki8vT6Pgqsbv+/zpQCdA
sm8+ihu6+gdKRGa7Zg0BKnXTQrHKPMXchUptqkTd8BI3rDT9CBhvBlnp7bY8UWZSGedDf0ubUtx5
oQdS0zT+30ctAPImnq4OouHfs83W2LpLbErYtwaRhKaNg/OrRrILFBraLffsHVDnQU9nfNu7CUvj
88RnSxQadhn1xYgWAJs0ExuJtr22mZBktYUxTp2hmvKIRP/oIOdIDoYawfnpVBUC1bJxkvu5CPNR
EDoiH+blvmOTapZ/wzrlYE7k/UKHv+HYWnh3Szbh75XWScEZVM1QShxbIvM7ASLF2Yr4cMYrPrxH
7q5t7Mp7YtjxSPS3MfCExwZEQEiOBIna216Ou3TXcpkzF97YqC6zNuIAGhzf6ns99NJFcMCHPoJP
4OkaGxJO9vo1oeH+JW03A/gJMq1g/5DRdf6m3AaRb5/YUSOYqyRbHJAkpxOyfLtoc0WeVvOztOp5
AoxpQwhpo+/BNXotAPG0qK/b8Hnlsf9f9GA7Y1v+xUdV/tihBPFMO5KT1IsfPksbaFW0+MHhONQZ
CkuO37W+SoiOTM1OG7m+qYdnmLpUxkG6/pOsAVCXNd+PNMVGuDSv8vGQDfyKWk8+Dm+66JyxquUv
p3V++5jsEAGY5TnskyaxKYCTReYziTGqCDgBl+/o/8cKOZ2Ft9Cv/OkGJ789VyCech0cAUxpV2rP
+yEIlVg8KtONZ1QtvUzFVNpkgctF8jg1k0/wdxbfazVBUGJH7rDwVSZa3TrU7XKwmoJh9YMglKwC
yV5H6EX+UY0tJNkGwlUktDPHZM3hRloy1qqbcfDuz3cM6cBKdoRnZ9TDhBajhRJ1tbdAsA6ghOpW
XppsgTOSRw/dz0RjYZ3uZPs6P4wxXtehzpY8d7/I9HroIFgDt5KX2bADLxnpGkUiBOEHpUBGxzgt
zHx+Vr9nAAS0ieRh9uuuhIGSmqC4vyP90RrYgRtr2YpGQPAPj1tynjRgT1M9WtRT7kPCoRSBbXHS
QmBfeAZEAVof0mVaoXgtFcaUAymzD0jONYrNXm7zsR8jwRXmoUWpxmHax6lQgaGDItvOd3ZHxMqL
gC4MWKELjYIU+zhrerhGd98FGEP0MhXBCBsfftJHKO97bR7Z8vlcEJdySrcwrP+KyxzhksTvtZPk
zb1j/LgvDJ0sukaUBgYTlg0A0c2Whsj8KrtYkc5Rm5s1Hwn2nByHRjKYA5md1/yHBmX7ccWMT0yL
IDd84DkfT+MP9if0XUW4tMY1O68eQeKPPGLW613G+/6Kyeyv2769tkM9i4odhXewmbHa2wy1bxo0
YmQpAUMNK6Ss1Rwa6o41RtNJmC1h3KPAn8khuTmZR5SA2QnSGK27Qm67bEmFZb1HlSUjg5Bw+ofo
eX2421ASEWJ5earAYQJWFsm6IRTTVM65wlBQ796jJMCPVmmbih8dMJdxugTnBQ2/VslOWpeTCm2o
TkawFSztGnOVb8BZY+o0d/yOPvBthH+fAYZf9TSPA9Kboj3ivuZlKcTSzNJdFvM5TcrHzBf7lqvT
vIuNtNk8B58SljIpKfAeBWrsgfz9RDfqheNdbpXiKxmYVbj9f5Q9Kc4KFTmY6NKPtVQn/57ixZcD
6LUjwoIpDN0rVtJdlV0Oyta/farY053Zqyv+LnH7YxKXpu+5FSKQQR4O1K+vBmW93lVAt+NtcmJX
4z/m1vikL/Ae6rhZzkRjVxCpPbBxptz5tPyJN+NxfiU8cJQ/0d6xKvc7aFxIJp5iNp5sn+ZstTsZ
vGp3XXCY0Cy66tiE1rJdX+w2sl+areIx3EG53Rqtpo0nfWckiAhrAIegpeIKRoNvjBB8OT7wAqFR
i9ibH5dK+ixa174gNPX+X2jM4yq7gwSed29RWIFTexv3QMuCSpqYn1OhfZZd/TvwFgfkw1rj1YZA
RQG2vQOcFY/AntuPG9S4aWqRhEgrOvPSecZoCxuGho5OW/7EnBvAdUfhHGonl/j7LWemxOhuk1K+
OiH1MH2NwfHxb0/Cc5Tz8GeexNvVKvzbnbKD8HGHq4NKOhzioia1PzkLseGM+SxqQ8R8HoSUeWkv
lVHODfA6AVcy2eb/kQzhTFxtz7Hi/Us8BzaYpTEl0IPa7xRhaAJW8cPSngsp25GWXpvoekCLZ8lx
n2P8XG1B4smKP7V3mmz+D0NrjBey8kme9Icz0Nwo96bRx8wGCBbLth24WxvzH9WcOvIMkdZL6bGe
xfLHG/23mf9znm3LxavrmbHj4Q10f4DiCkIa/7oyqjKSy36/zZzl4sqd4IXbFVmRzeNJ3BtPCTqS
w/opQMvp7rB1yQGGnRFSkEkLMdBqvhwvCmMwn/wHB2Fsa9SHq0lbaAGYSFElbzQUGXYMhRNEKPQN
KXxdPcsB3PHjfsZTlg0AnwiizI+eAM9H60O2QiYE8VeGay9ErXHEt0vu0/jaB16DB1rA7Nj7Vumy
T2kdOm8ygbZ6jluV3J3GCHDd5KbsXHfioe3DlkDA7xBjZEEWGe+iQUoywgbffXJDwBwGVxFlp6+u
go1jrX8aGYjsoXwoIuwblxIxhMKREU1kT2UBTi8O2Qcbd6LPUu3+1P0iKFHDILg76lgm8rU13Teh
8b6iEwqXskfnJljF+2r2VV6LlglUAXXvAzQcanF36ftbIa46puIjW/6cCDo88fgVfV5DN/W1D+bP
TbL/MrV6cPqE0T2y6rJIe53N5ddulFwjxLQUxpxBLwFPGKN202ISV1W0QCr1pUBE3a1b36QMJbOs
y+W2NMdRLvPXmSIJZbuFSexTWlu5Du0ESVbnN8EOjipotAVb5RwQuPgvkkjcNmadvmkBfA1mOPEH
i84d5UPPC/eCtRtWPUR+KOCp/GQ5wt5FBuJvly++qek+aWGU7e6hQ5I6ujfLw0peBqwjngP0tRnu
emZeJ7qDh5sSO1l8SCxvUe8+QBRr5xU1FljRfFHgPGagmz7286IfgQhB0O3/tpLYw6Ph8JLWerIb
Wtzef2WuXRIprGFsmc3RR0lETwakqSKhJ5pu9Dy12X6tmg1rKfVj2AqV4FegUtF/DJ47fvM+u4Vc
R/ZE8TG+FYY2jq4iykJEO8w2kNVaWJjXMQWk4Zo5ZHLzoUGm3hSRlnkLy2M8veFEYtEltMDgLPF+
6imsjYr/j1sDJYZCL27IYQMz+EUpNwbjtkC5eS0OG/rm+0edgubvn0ukzD6W0lsysNYGILLIKlFm
Q4SG6G9VFyZW9BGNT8X+BjwF2+o78IT/o9cN2ZtWXyd4wKrCoAnEcaCE9ITyJeMkghSMQLGrzETq
ldVYSc92/TfLmBE2D+ksEaOcIcSs1+JfpFGWxzz9xpyLqytebYyA7XM4IBv/p0Thz/fJbV9sHxD+
c7BePdOLSPcetv+LeRVn26ynRcXC6xq6xndRKY2THUf80v6cdy1xXw5ja4EgsW+lZbTbGCB6vuNw
mkGOVuqAty0lldXQvPEuO4yXXnMswqPJaIgKkjhdBgOaMc5om1L60DCxcuXCMlk6kIgiVy1FvoCA
oM5rL42HR1c/hOfl6Di0aLWJVTwwzEiAGDW87am7l9fM/pDGjP9owfztXylpqRNfoDHSnrocEkT3
7K1tjiu/gl1B5rDYvJqypOiiIXlicBl9oc5jNvYFtFQhIsWWL8vSeYTuaDYAmrRi1JkyA9JKgh+7
sPNw9pW2TU6Oe5npcNA/SuVmDR6walwfwxXH9B6tbY3QzF0M7R5WwVPsoBkW6UpFW4diiGTjh4+J
T0ofyJ3TwUjSVtqzaWnWBmVcvyUZ7cpudY9VFRJxaLKUxLHeLZLKL+MYnqq586nB/HcY/pZ7kM89
t+aJHQZ10hctFboMYcQKdBS8XonYNcT20tCBYpH11iPZU9yYBbcotAinm1i8FfAFR2hl0B63pK9I
Nu14UY1f8dkpNponQYg3S+8gTYGEX9nQozoY9xyFcknoBHC/30SVpe6yvDKpj5wRA6ip6TyaiEtM
pZPhmo0t6sdjIk/PTIwBpuH3XrZFc0WIpVdKhOBPyelpA1UoE1oq0x9USOgluPSEncgfjw9wMSCg
cENqSlGoQft6zrLWxrADq7UmC1JlJmtz+zHIUXtI3j8V5VcBLtc1WpxOgWgiHfJ2cwQ5rraLiUwY
7DV62nGp35Y7jv1ZONvyFjA4E481kD8LNT8S4CjKFr9FOBmKlZAGigtMA79uVaDSWBl/GK3SGowE
YxnuVf7/a3K+0EChQ7W+bibx2kKopaAbUCzwLJn4LM3cQxQQtsvvAu21zi8/EpHLIVJrJgDulk3Q
2HYx8ukvVr6K+kQx8OJW6Ri4MB1HCaG7zY7Rxb1rzJn0XnpG14Rz8Gar1yTM8ECkNASKNpPMOE8r
QxHuJWklzoQOPi/DxWpWtECnd94Mbr/HrgHYkMB1fT8fmf+UuMmb2GSasphWikBSFeCqKWSRr7g0
vkSI1jNlQ7YF6sMN2SLyLImgNXJVfw5cU4fz8d+gyE7+fZxY8SHp7G29e7O31jo5bk+/J1hENF1J
fSERFghNS1C7GMcC5xve2ZyB+OHMr/1GAYoxd6yUnMldnZuMCKE0FU6y8/AKsqfGJO5jhzHbx2Ye
MfKY2bZE+Fp199oV9sBVRfZRPUOAu+Ltw8+cu8JMSP017cjtzdWxDTissHK+1sZ1TzU0u4VdACDa
9AgUgon/rrapfOKdDS0L62wYWRy54yNHncDtuQtI3mmtWwx7hRsXxZNBI2mzpfF9xRCJFrq3r5y5
hgXJfO0ppDyBijfyc7alSNmBgqq/NCRqahWzhUnPmYk/MuTcE38Hje2W5JKde7/6cqBc49MAyBHv
k9D6UHzOWMqJDH3lQf6Lkp4gzalkNUv2MDxQjLxZOuZXuJTMwXmJkowULOPbMGsPaeIis0GCEToC
jX7HhWypP1Wof9JyQO2Pqb0CCpoXAtjl0TeBy47hVFzx+G4L29tyiNY6KhVtisr1ZWk1YD3ILBL3
7pquG6UuPQySlWeT9N3vNNjdK2BlJHwPj8yLEDbJ/WDoAKx5u2S+NBRMh+47XMPZqXPzATLEmPDl
L5+gPpC/VjpfCQsc99apa30HSPUBRB8nYL7Afdosubxmo9ONtjFNStC1X3QQ+GAFLsNlDHCxqhm4
G/bwALXSCWSjCOU153E5QXcgy/WfnxecsVvx7cAqHQaxMsvAUkX3klP/eZ2opMEB74d9MWLOF6MT
+0sBteyqDex0hTJ/xJGpZlFsj3wQZIZJkLFXePKKUq+zATzsIGQoaSEwWRQzVfKH7o2uBPSVoMfV
/zOZcWvs94G6wsCSMW7vrFkufg4JoGLjkIt9XokfPxSJcpf9WW0bfALQPynHwmrZxrETjNcA/uqI
5uYVyhbY4WCSblRLNdwpdd/H6lmMLe5CL1DGvkUfEaki9uNVEddOQw+36TiUaxtze9jpyGvFwnxr
/8gF5SeCf/uIldPn7khWmVC3WgVWcW9oaDywb7C/6Wd7/GPnt638LZRVQ7SWx4ilfuFKLU9xFpb6
s1iSWXdGhz57jcdhfNYojZB9aVT9gSSuPq9L/unbDb3Cy2A4/E5fAEUCoPTaNWhkQpQ7AxEa34e1
+sKsJS2zm80CxFE/GB/JdqXg32jD/XO430Nu5RuKOP2/dzc2amzKbhs7YIOepvBB1eI6bQD7efLv
0PwEiHaye7ifVKlcpAmByhNgVvVMcM/HkJbZBDj4qP4JXXwKYdQ+2oUIdnEmCa2O+uUE7W9Y3dyt
DHTLSE6utNki6KoTQ+aleDlkFh1u5gaUq1Go6y4WB7Et73aC7JpXf1RhZqafIOF2kgkkDLpciyPf
w0Exgm7brMV8OAj49Z1mIDUn53vFwlOZo5i4jUdAp+5rY6V3jCLHSiAD5mhU5GtKH1xyNuqtLo9+
8FcZdHH2sD5Ck0I8m0yndqm53McKJGJwvFqZbX1evhblFCinDk56GdqGJTus11dcdmVPThq03kqM
wn6jdQLdbua3I7daWeU2cNgSAji7dC7mNQgjQwF2wfHZmkxJHmLHW2oNJzFSeos8zJME+tQthhrL
SBbvkj/LTnwCVBStkOrkj09JPlTHq6I+LF/NLGkIgRh+tBAQ3QNCqxSaKTmtc7RptQooh5tZ6yB9
oPxk6r+4dMvjimLY/Tsuk0wXWPmHdhewWXPpAZy/jZhUDMbQsDyrIYObQv4jOqwtcURulEoeATKD
74LIFHDzFlBcv76rTyfYVxV/ysBBnOTcguqCcTZ3DDZir9XNRmZ09ppj6dF66g5Q3AF7YkRXPto7
qdEOstalpFav9VwKifRQtjecLKCR1ZcuZ+9uULqMag7nVGCa9iRIf4jnnufx4A6XC/bzJmRtAEnD
67H7Eqp2RCjLCytM3yTrEnDGtwK/Z/UEVB0PPl/ONQsp0ZbOAqHCkGs/kWc0WRPEAifAGPqBP5OM
NRkvSHqewMfxLkHFdyxS+zqgFmZMp2tIeS1YVh0dJ75iG7DzV7vcvAMcLXWyxlSfyYB0b45wodyK
R5F6FFDmPxD3za0Wz75AMUGHq3eVOd34+nq2ygfbtU9dsGgyQ2yL6jxDvkhrbGRgzMVbCdesI3TK
5HmedKVPey/yw0uY/28kE5el/z4qvd/cmVVGY+ZdF2yRbKjfQzqNupXD6wD1w9JoWkzTXukGJzkf
pk5DSXwWXk3H+kgn/xtcn7Zq/qaMgM0Nox13L1lhVjN9eMlxiI21mTjWcK+LHXYokALqO2om3RNx
ybFCC1F8+M3SMngZxomgHqtcdTs1einbqXxM8XrjxbMn10S42XdMitzqPElyntsoNU/uiKI4Svs1
Cnx+T+/oArVl0oeqjMw4DXuHCuqRZHNAJJJrCFU9HMoUV/YXFGSILcvVEyvtz220lEFvCWf9o3fo
ovirDMtqPYjDOcwnrzfR8LcKsf3RqGb6cq4gR3efCruIUDNtQ+MhTYSrXKy1PBusorsGgtRT5+k2
63dEl9xvEipBrK1UDsuU0MTl68FggDFJLDm/Q1uF6lWEj5Tx66nRLjhMRX/Sz1eiFH7asT3S5ydU
EF2+zntx8LTATdc/hOa52oq5MTPrBoRval/Xr2wTCJHEVdysRMt/j1spXTXhwseAQHtzN/0fiW15
zZIpN7TgSI18O5PLMY8NGqEMlFo5st3uuF0KX39FF4lVbW/c6dRqJU4LSifEXJh4sHg8cl43oNe9
DFjI+W3HsNIEeDZcTEzfQmIcjK25KmDsXPJ7XOy9XbhL/g2SYeJrcJ6mFdWn0CNZjVYdpUfxjeaQ
J3SaRKK2D8PCNYFyrJanA1bHasJNsnXZ/ACAbiP52KNjeDdf1cM+qZjwZmH4Bun+xeOjYY6aY7DW
zLOYuyQLCe+Bop02rxAOBiwAuVE63mfoBRzDtq2TIsZ2QoG9HUsMTZUpMy1MsP14nONxG00RDJzn
TzbyfzxguYQG0o20HJd3+Q/ulw4hF/ZoW+ZNloE9fX22Q/41Pmd0JVHJwuTgr3szPCOrt0zBCMd5
Wc4b1PupUUyu9xroku4Q+JR/uf2sY3n5U3VGFqEtvpFYd6JKnpG5LyU3N5j0Lqvrf5u2uXabdLJx
n4cUOoE2RESxNYFj6IzROH9KbMQeVm7UFaxBAGJ1x5QBqVilkecR9JZ8/cwvNRn7pnoU1HxEDKD3
6LMc4NwwG7os82jETyGa7LbHNbGMfsoTyFfHTx9BXVooERhxxKuXwHeQWcS63dCqVyL/H1xF2nsn
biTpMF+9A82lPFxBIdr/5BfzH59+A+gawN/5vMSFUVqKw0sTx9MJQpzg3m4nNJ+0QNK2Ue7LHU+Q
LJPFY5icbyi7l8VC0bzCMEi/C7sn7ecReXKpJjqtfCZldf7k9YyqHhnsHpTTGubtkeQqyCBbauSK
54ljmt3eV6Z/fRFx5QGkhjUu9re/AvrRPrTym/KQsYW0mQ/Pr2LQ+O+FJrIzQ/Ouv5VDRvJzhoSg
4cvguSrDAZQJk4GtQ6WVQU1kQdSU0RZUk++mLrDUSqNZaeUbaKX3nC8ZcDS+QxU3nG1jvkVOmJUv
WwpOQCFTk4zmx/dkFd0Z2ZJI5h3usYZCcElLWK9UZHUUI54t9EnhhkhMVzhxQHQWZJv7Eh/3IY4+
xnBcmsT1l/PZ83z16NHESfCzmIqmchxdwBmjd+7VSoox+PYpDzyQPbU/pRxziKmzIDmXSias5xYV
FxN1CN4NXo2IIaE2LbRetbrqvgwmZvBkQhqep49WVTqXFlIn6RymJqcEa5W9si8S061XXhW1b40T
mKNxqqYRvXH+GNt/d1oH6EY2KiRVf0xWwVVYsqErp+jX/4gLukqbiM5TTpk6NPkWbGv+O6qXHHvt
KThnn/KCK6+7BItyytG7ZDZH6UxMWWKrFtAv7cv1R0nCQchIMPbrIIYUwKz+FdimD7MVVWqAdrtX
uRMwxCq639lO2tDKuFpDmPRbuVxXkvJfug+T6Lhq/s6Nr1S+ach5VxWNJBs+MFuyQO/jp2q5hb+o
aBK0BzPjk4HZJHunfh7Gl9z5Om5Q6dNF1YxTS5LjSqMASdLktUi2Kt4b5WaNKYjMlqd4HNSUPk1v
DOWyYz8r1XzEhV30gVJ6IXW4fMx5CC9MHvRB/wAbxFOdTqYmHqw1wq4P0LM/9qoyI1n+6Kvn+ZN1
+sF/33/HhHNF1MPYEIi7lCmw9WavBXhmu31WrQ7VRz6Ou9B0yLp224W3BXURIbh/WHXXv1rI14UY
qqPIdL732KR5tBgGBsNYGf6aI1ba6kmOkfx8yJitwRqzFvIOt/iQnMJG+QdtSCgA+Zd/0G+tnjnD
3ztzFj1/CWLTSmdHSe5JUe1bedH/wUEr4bUVT+Cx0+Y45SaDHSZVq6lpzkqH2aVPwmf9HKa5m8jf
8irCNJR/QwBAVhBCmyIuatIDXCmjWNx/yVpSMrYqBIlxasjf3W12snEktQZ9hLzCPOGU0Ta+ihSg
4c6duwa/+tzXDT5Wx9v2gzcoY113xRbeohrGkeVhq7Wfz7NbbrVGlU/Ay0Am/zyjYd+6JSe7tbRB
JSLRbMyPwwgCTJ4AboKvxaVZad6ARme9jvQ66dP8zwe5suYkkWOsjlJONjUwxUhc/VIVc/qBkc1J
5A+eQWzvywXawfa5Fhs6J5Ngn7Xo7r0znGcTC0BLJwH6lj8h/6b1dWtvoC+lLzO04TysGFQ/pmLa
fgxylt+FPuv9COurTwZSi52BZ3aB+xMUq1CJs6AV99rcpnd0X5cLaUotAXXzBWLygE/XeTdr5PO5
tyTTBbwSzlqr/UYOIqqHZNlBiNZPAM7aHdgXEfzXlKrsl1hek339xRflN3nx+AFY6TQ6UV9jgngz
sFhjWIWXrugqaJRrUjNuqDPivYcZQAtVFKyEn55AFLgyqNZBbLQV34k1Qv/+6U6me6M4bXMPe5mD
pBl1jwRKqmjZ30jTSXuAWbCZ2xpkLo9OZxrTV6wdnQxFPabsjLDmOOpIwwXvwYWGB3MaLsDm3sT9
LGB9g9/NoAGMg6WsK5Ay6c6zsNIoAl3rWTecJJFNbDyNj6zqEZW1nj8SDvoc7AgYMelXlcFUh2mz
a6XDY9Q1I6R5ez9J8hMTfuUDMAcmuHK1ggxQd81r6hnv9K8lBqsKol9XrQUlKSelpCfXbczbB9xD
gF+md6iRC7laWSXIDbFcQcW7OlrdUGGn9E2g69gfrup3PpavqxfK6t3EfNK8I/ngBiL+45kI2URB
mLt41Q0VmsG3OpkTtdOwgYizCmFm7GjqafSou4oZJtz9eL7ITTwZdVNVLAit6yWZ26vFd0CfRBsb
UsfjeKrB8ZKBVyHU2CvgcEoc9Wowd8RCl4VknOGXfrhuYY2h8B4FV/cyRpM0SFLx6M1FaQpaegMx
fPHuBxaVUD7xGqMSylbFJZsktKu9rPIuNXdkrALLqwZwwIhTGIbcWO5OV/wcccJYwmkV3n/9FhrW
U02YaXn1DiS+wNrpoqXxYK11ZLt4WOGy9wh8xdYIeQj5rX/+lF6QVCz5cUKOhZMxGkHgj625xFqX
fIBrWV7E6SXnLQfYWsTabSCaEfUKta7Gx86JIHA06XOW/wIy2vepMrSK2aZPL3812e+QKRDAAWcc
kSmcddGoDsks1ORcjjHWP76UvLWSe7evP2E0hqsTTq/SL/37+sqSin4n9KULqUlxZJDceo6U7c3v
jy3jYlfBOFX8WJohaip9qRBtmwY1Ds/mI3MoZqZm0ybyq8TA0eu/c6anElc6rH8d8oU9vlMV299d
kcAXtHxb3PKQ25gaMbC4INxVi7fYcJfF/9PfhBnYiRA7AVqi88Z1m5t/h2VAicYg7b5OyTqlNCMw
AAvQ8bCCGd8OovVSYg6PXRdjCcxz+tWf1V51nFd15xgVP1B4SP+4HQY+vzfTc5xOwY6FRicZTuWQ
Q59D4He2ZLiLXHFoYxL76oYk2IkTNPXqztiid56PJIIilMriG7Am8M8DTOm35XVm/+jhv9+3XpUs
lo/lXpEgtbMfGJhuM7JOlQ5/MVip+8h8QSH+J0j1LtUihBOWXx4Pv2xBLUVwbChIfFsQp2kOjLhK
fyjDhZjFFuutQbL5Bx5HUih++1LNLUSCVGmk6QuzTtkLoMYznm0TWZqa9pLPfq/SKPJJ9TNq4mV6
zRJlkKBtpb1/YgIxhray1K3gSL8Wbu8WSWtBDQxTWlYPo0kA2eYfNnOum6j7/TihLTCz2I6dCdmz
7LpJAmfmY42zoFwJ1RpFin4SrOvVCSkdYNecNFC3yLVORNDwxONJboAoVwf7IArR6aeDJvAiDevK
yx/olO6nCB19JlzweUk6V8klgpjUzPadsdW06YB1ob9FHH8xk9Nz8nnSTCeYtfQ9VwEZ7x1mmdYL
/9B50vF25WbYGbvX/afUPMa1uDwb8k3+nH32Yn3Lb8RFvSprGxNF0IosG564o1AhUCY98lyxM4kk
MywZKFrhH8Zs+7YGBvMCFTMsUAXrXpiMGG3RheFi79krOBDEG949CNPYq+yUcuO7aPP7JfOsoMjJ
hQDRY4vOSJYZKBRclf3VDaYl96fx9FPHsecix58GwS2tRGVt/8cU1PXSHpuf1XdN2yZwD3omOJKL
oKsQWW5lCm+LjrPilZgZbCaso9YlAyFSrbFN9C9i396xS8DcX2zhL2zCAy7NkDZH6RKuW+Mp5rTR
w6A9LHlCke65t36/+7iK6Jjw7zkArYTuuuflb7SUGIJsc5E+SSO0TIzsOpHmJL+4RWEjvH3VR/DO
HI1No8XvYwCyvKTLAKWt40ZlOvoVWIM72iihUWGy61l3ItDU2cKpvPb3V4iuAWb2I7aHbrjKHvEx
FU4OLZlGQA0n0sRJpLefcl8H3T06Q8h5GM75F0HrPSsr06EhWPM9TNCMv3TOkbVk1+yEvzQkgIJs
4CHAXJPeFYki1BONGdOq98N0KyPIy3Xp/996BPyTLKT2h8s4RJtz3HP8SsITfSriJl6bwcopzCN7
t/hMi2RbAn0Efk3YeQk6qD4cff8hOD3O4EpTtdGa/XVB6DR2ZX6f3woA7LbH704+rGU448RDyGGG
gj9z+wOU57ita28N9GQfzSd1QNTb9wLb4UvBq4OhwaPWrrDWNyKfliXT45J6jUQc+ZVMRF4jFpjt
ogb3TUbVySVwO8bIauCaOAs2vJqG2EEUOC5dntZiGVeE2ceji1D0j3HjfmolxEI6zwKyFGvqt72s
3yKH79MUqbYnB/pNnfCywGFf7IDjC8P0aBiOQRV49+pynQ2nvgKjfTsPqrjCQGnnoxkQjZjCc1RI
3sqX0lcPct6OgoPaNXwnxmvbxSiKodWJAT1mfhtXCn+9hhgYuY2I0h9DObK5Orai0vSlp0c3OaLB
NcbgSPsCvUNsXD2+/p72kl5fAcTwuuvHcyeG77c2Ga12QJPhrbu7rF1VlSJjKMU5W2FM7A4Uwww5
ZQrSySN7YjwVryjATt5L39535ngNBxsh3ypauLls0MWkz9o48kVlegcg2+XTFGXx2DtSRqYIO0n6
SKLR1rY6WP0vJPA3sbGCNa2k7dCqh/u72jqGtsJWemrb6G5E0DBmnmUbPPvtcYLZcc+1w5lMPDUW
Q8k/xdczzK4O+vMlvNUakWipG/P+W5nvEqh987DWvEeLDkN0DUDbjPtje6omDR+d5ZWkUEbNsYJ5
p1LEwgIxTu0ioK6XprFJkfrgtCGoIhlgfeBs10cpYhV9GNw5L1Z0t9da2TYB96nV2uXQoFl4KeuA
JVlDZFPZm+mU1knccXV5oEFoTSazxBZQ60KZjfjz+90UkWffMERlOKUOFJ5NrhTaZDcDGJlKNojF
T1Rdb6zvwpyoInqBR+Gc4bINjPHD1cLsgdyCbKBVHihxXtTwcR8bNN23Q9LxKpBvTSTJ6l/mCqO3
rl47Lu1QgEc5ka0QYv9ZuxDk8xfVF6hQnG6ubEwn/kroJ7Cr3l0WoJ1fYS9UM6iAhMVL4PoNA90Y
z34DtWXj/4P51ws1Y1Ug4UXYDHm0jIkOW+C0zy5OK0VoxlIWz9o7m0aTwLUvvuKWH8klpYDVSkRB
KHcyy9DPc9IP5XWDEAle5TuDx63F56SEXuqw+i+LYERULEOZM9u2kyYuyMDCFQzKPB7ZXGRhOeXd
t+Df1270g3olNWqFpVVc6r1leavf6xhh702Kk5hkolqRkCJ7OvshU9GZruOlUdLfy23Jd1a7s6QU
gMCAtVzYl/sqLhdKHzCL+4EE0y6CnuUlt726Vbd1S0bEZnpQA7Fsc67hwgeb1LLRjxHwx5XM9cci
K6mKlygsSzXljs9lrKP5qjOGr6rkZJUROS8/3SFIZikaBPcIFQapQgcuGWNmuspEy1zjwZHfuhV7
klMOMq9DFddSuMX6T2n/slr5oO/J8C9EFrwSLoa+4tKDrWZSAJNr/wVXWEuPzryhPHzhcQM7+1gq
Yxau+dZXIoiwQ9xAOaYMORmR8yZHOK2txuUGZ2ccUswf+BRumxC2hkFCzmIpsGqdm1B/Hmfy8RZy
85+ixJ+1qbGwW/h8l39KqV6OUb3TL+AGTZ7tDGlQLQEzELFKzp90bbNbUm6jKA/PBqiW3aCxMxlR
PEPXk5qGDQ9a4/7Tz26Mzclp3o0e0ez+jLUUGFWAJMjXxuuA5VybhBZxQEaTpYebLEUCKsvDxKwg
nLMxCbbsiY6csE/0E9QFxb8LtmwpTjXxnpnt9tmoWgTwXzha4cvk0EzuGXTPlmEE1tCMe1qqn6/I
WYSZMxFrTfJp6Shd5ZE44VGNQKSX90b5hjDNG7dhtOlE98PA6XSsupJWPafW3Tf6nz4ehLZiR7V3
PEO7ceaGeJtd+odNCM3TSAj3bV4w0ksx4wrWfFjct27+L9yA7vJ+325/7PAKfNRTN8zcWy/vLIN5
y/J32P1mgL/YzuhAb6RXJNAOyBdNLB1PYRDX5+CWX1Qb/ZtNwcQgfqX3j+kO9cdtO4adMJdWuHXa
4KnuqnDYXxMbD6YmuhHNIeIJ0RO1isLdcuyUcHxrwkdwpNxVHDraHJRaOf4pR+9No9+dkroUNmCU
hCwIDDfSmVytZrnUmtLa1n5S+THCi/WHXfrzs96fQ3NNBPxywiUIv/9eafsE3HpTeoAjbK1w4seL
JuHeqNoy28QEshecnAuTBKHFF4Frb1iBFOsJPed+vlK/wSV+OVEQY6aeHQHgq+X/HkdKMLDW/lOu
ePS4vsPXopB3eHiPjfqo2DmpVX+DtGZYdcWhrXtaWrSzpVNcUU8W4/SAR9qnr9esW5YxKt5tz0d6
X7HBMeyXYjLGCPAMgA258rc23U0Srqz3GlBeUhJePfhPygY8xaF4yy74dSZ1zbJkOAPLAM7Hqf9D
Yt9SCKN0Lh4Ndn5a524rWunQ6v640Efu+c/wBOtFzl2fhqSdiQ9I45GjqQA4MtP5RSoL/EtIbTmo
EocJbcVWq6Uc9GOIBERPYpKclZpZ+11Ot8X9Xj98NFaOhAhkbI/EYZok5G+8A+GqDzbhqtqW4979
7poGEMenArDBv8AKxqb1qMFn3GxerH4cA/va7SsuWmBTWyxMJf0WezpxAFbUGp+JP2VpjfZiQ6vU
xuIDTMFxmlYeMg4HLxUjFxTSNmAhScWvNLWTOK7U+Xd1nJ7/EzAfLpF1VqHKYMxyqkJTk4dCIfVn
wEEI6auR6IVNlqp1Xs6TMhy4tWAmyUPFACrv/FlJT8mB5bH+VgAegNxxvxiGd6YxD4oNnqDovBTr
fFV57I9z57yx6aQIC5cLq5Ve29UVZvI+0R6uMOmiTJeqc4p9mKKIUvDugg03UcoXy+P9r6PySYPP
X4TwLH0j60UsL2a+TfhxgneW2cuFt3alZFlhtP+mAY12vlj/zz9UMlcKsyKzqdQHndPr7oura3RL
cozgtiA9gppgUKoWaz5gDH49uid1bZsuGdp3457aHfW3cvFf02FQmIrVpLqxhivmI7IRKM74GpeE
hCwFDcmUnMt9+FCPAwVvmq0yHP8/dTETCtRltVtfE4ngWhVVg4C0Zu2JQpheBPpxdvpv7t708sZG
oydQjnZ5wNpHyalQDXIaDclQ/3AHz7NoHzgKsdBRgm4AMyVDThFJ+Ft8p+7rhZC29V03WbV70TR1
ccQ4gvee/quyUFf95FHcYMlrpGp2LePYF9J5q7IgKdnTd9OruGMQIFI88gtyxAT4JnrQ/V0mERZg
aHmxOfL1cGP3d7LE+AgRnVTKz1Rjx7xMhh/TIOTUEuhOq7CvzuDQri1/ZV4s+Ql0J3AOu93Bq5Bt
CBOIJ6bwC0DwHo5CLrOv3OoxVgueGfEZ48jLlEZ5CTYjN438SnhFbKK3DnK/Ahg1CTXV1ZR3USTs
3CdGjP0X2tN39By+niEfCQktEnwps9X7iHxx+V8yFMjl4FkAOFItkjRh4BXMBGohDdufNn/6KIQ+
08l55T5wuB8jTM/sKigYT5GUdklMha8KOLLJKssFJM2q8fhiXwG0EmBDU8aZ9+mR7yHzw+UGiH91
zz5/crHAhxiru0qr9NHgVYrBR2mhqlaUN8nqZbf5YUiMsCXSaURCa52PlnaEhEQCMor8RbT5PrIS
Dcqej6hAsqMCl2FcBIIpPmj7ac9Pf2R2lNc30XXsSvCJ7GBL7JfeWyKz1IMhKFmH8N+P/7xhzu7y
zDbjO/3qWI1mAHimBHnaKpT+Fik1Xv/FtVmP9kbE6K+EhOTvbn1DHFgO77r+A5i4pJnd9c305Dmk
v5p5zO7VpEv22ijx1S+zTQ/BnEWMNAo0P8pipl+xnvym0QnwkenK+qKueioevYjmja48Q9v0ih9s
rN8wJyVLukbfm0l5cr+18cUUW24S2PIfc/96RM7h7iEXtGjN6ONZxYZJbVfMXbinVniqb3aB4bC7
+Iyc4ONbmOx6VUbGviAJXvWj8kcWBY4Ktw7JvQFS8oAf5Gxfx0BgelMnWhlIvEmxb5o+JIq5T/7l
xWBBwcUB5/3J6Vza5lUfrOeaC+CZvl/rjkMGhCYcMPBV0ziJ+H21o3MkIcS9SS09DHUvinlFNBjL
mrRFD9mrc5xQjuwxDtBpCm0pI2Ch7j7Xd/1XmJCL9rdMav71LWhBx9Y8kV25d+0CRWIS9M9ua6GK
kiR3mAZL54JzeXCLUYIr1JdBxthMf+YSFUBwlSk+5o6KDvgdk3d6bBQxL4NE61ch8IGJaiXAjl3k
iffzbAdkt94w9g8bsSN7APzTiBPLb6+f122N+bb0DYvKz9fAbi/BX6knhF3qnanvtq4W7iZpYrOh
SVhzAItnbD1KAL8eyUzRNsNvPz8kLrEVeCTF1Gp2SNjHOGQSHcomvgM0LMvKSyuNhTC73SSxSFWG
R0tdZODrpcvhSd0AKhTYVQ4TjFT0mKJnOLTEuHqIN/+p9gc4p5Zkf0YCEih56cKvUA/51/yfYD5N
37TqPY+tVFnJh3mpeNZNCzzemYJZIBkciMnyVKb+0A0CLMZL7zUrRyBo8NCvLO/s63ijOhJNNcl2
77UgB7z2fXS1/J8Lw5bocbRlh+akboMm6/xMxd1HbvhI4g6Y4mVRtQYVgFpRqutW21kwCfSmxp6U
72hDepRnpc9txpm/ZZNuOthUjaDwUw2+QxFKNcGg8ckGxz8ZaaegfbZ83qCdMZ/eOcCZZaG/zOZl
SpPHCvVIPN/5UDTggrlGsb8UY2MGc16w96zZwKDg7QIouujXBZhqXVPtSvsMCHxAaapKLI2pGJ39
BdcBBadUXN9WR3FpXC1429mNS55n2ccfjzYbCf8naNO5YAPE+xOxPybkVwty5L//YTjrQafuUYtz
2iVOb2Oe1NXml/lRWCS9W4121+EQ5/N/yN4x5cb5/jtmVhcB1VZaym837fSjl7zmFqPMIBF6EtJA
9KhEoakk7OoJkJ86dW013YVkv7PrQwRjTHbMkosdNgFDUu24WibkKTSsY4YqzMEtw1ZgyDVy8Jpe
vxUpa9uGxIOu1Iw/4fH94JmOiwy/F3opxK30MAJFkkafXfTalhYJfq5m/aTMwTN92kw2Ns+2KSIN
ccW2fnCY6IhoZxQri3d3fkprVcas/9OvYMw8MHG5XUiFKXGSu7DC5BZSbq0pd4Yd1EEhJ2MGe1XE
uLpfE4R86KWWZH2vHj1zhq1ucxbTFyMEpPvfyXHAG+ZiEa24ubp0wthMeK1ekf2ou9gyMCynz1Jo
0M3nprV3OZZQYcKdveIoBMqjGcg+IZQbzs2TrUGTthW3zg7ioSanbDivtGAOdJ47fgQctPT6hDba
aG9XZ/IK7eaoK52seU1hk4l7TdqhcF4n4YOFlkHdLFJ80WUeB99X/xZJFmLTiQZBhA3Ubbm0h+fm
GDrLjKw0v0vNWVSmS8vweD2cFyzN9LE2cr9T6ojIZl1OFeGTvaHYRzocg9bh9DRMlKf8TPbu2+K2
yuWdQdgMt22BE9kCcgS/isPPWn6lbICCuGzf5jLA5lL326p8pzPqeM647EdRpyuNfmJRG1dyi5OG
TUHpbOuG1GGcNp8uoWWzy0ttc/q9jwxm/hYtciBIZyjRMsxqohlj053IJILdqFhLsfG6FjW6+mHn
Hh8iBe1B1OW8LzruYXN+fZMxB+g1LCSORDxaMdt1d9ePLopiSFe3DBtYNRIirXDfU3HcG7KOhBF7
5QbMES+ttlo+uPWuQQ4IoLM9RXuQkFBG5QdjdKkSXcTBrlFE9AmEkWWZAn6Oob9rqdh1WRdLS+/+
SrLIMIouFl4q300RzFsTKiFWUtaikXWqsSCjYkLA5Mar+FqDuhjnP7wNO7WDgKRGDoOfgqszyIHX
Jd4RVR53AaTiwDETD1vb8Skzi447otQS4ArorKVsp/35DyKXAzCyVBAvewVsn9Ff/Ho7FpsyaUL2
20+l7wiFPylGp3lGfX27qUCqduJ0tH0/eRo52/ELm7f05uY8wqSoGQIDF5NdkLzSN+0mEwASRTiO
lIzX4zmq5a+8Gs0ckYQnk5gufMY+KDPsph/PT/5m7ztn1nSJBoa+ll54DxHgUJSVe2riSryVXDSK
1GL/qylHyfFCjfTPgxk9zH/zcLsMdzj8mRoDNKt9lJhxsf+5lxQG8mItJgwNzMNxzV8qQIsVN34s
B/IBv4PJwxOug30QUtN2+DwEX5h0Z+NG7v8wb/CHcBk8Bool7QiSb1pVX/XLBUuVA76IoHH0piok
jfMkoVTKR2wz6exIGMaCI9mfW31rPC8BxVQ2/QkZtbSzonwj8kp+6CRsouwtEjJE+4YJDZ5mODwn
Aqp5Wyb9kv1WNmeU88Kt/BhQ1UrUzROmbqXr8dy8TsKZgc1/OXCh+wKgoLIXzVCQ+5Ogkhk8aSMj
JsnrSpQhS85DW3QF8sAY+ept9zbsfhw0Hy301BBlmTOGUXpt1RvXlRgaQeViaKxPatrW2DTcUChe
gSG1Zqv7iE5Nf68aT9vLMWQj3BMHtod0/SI7BfZhlxHbcUhCGJHJN/G9GpUmd8/ezFHFWaFj1LeP
+aLvcdr9xsW2TNFP2ZmP/RkQhLvP851/PDYbtWaHa7YZKwAWz9Q1PiAlhrxUTerZdisvyJKVOESS
I/6PlFkcKgXo7vGo+iCnznIxtshowFA3s4bs+uG6QJbxwBhDnpnou/mnqhSWQjrgOYqCwSTo8G/X
FadGr92YIs3KA3qHa6XHBi/NjrcjEihMndrFtxxbBNeba8o5xY0HbqQY/HclhRCT4ASJpCytEVjV
3ahQEIcdg7hoPWRy1u62dykm3o1g6fwtLt/sTg14PEi3s+CoKNT5POBp29ZyEsOZ0iHFeRynmFQi
Cy9RylA7BdorMQp8HWIpCzuZrG1PkYiEAmm65tIQENzwIqYlGD0XsQN8k9PrYtfFg3e9d94AIxPh
hL20kLEbYo3lPhLixup3YkVY7rQeVwyZnjSDr013nJiRVuIa91U/TdRVsVENbBfzkASxVXQ93+Tm
N5bJuyR9yi5ra9PFzReTqqnFrsD5DfhUq2Y848mcEO0oKjy/XR9hPJ8yJthb8wgoiHVR6CFVDu4S
n5iYxKpPGKN64yZ2q+H6MnBCW/sAEMZRCHq3YtpTI7/DGPefCb0JVmUdZYr1X/mSUaZT+Raod2kp
9FzCkQ58HqFgF/zkUqk6MZJFexoEdBiDMyjXNT+1pkXsueXs6QpF1lGfOQSqXVvLt86a486DHlQ8
ecvFelI11jmjXA7WjfvkfXv47i4rx4gE8HOEnOqykdmFKbMkr21M2NNyPzQXBHVgR4qBT1iyvr+q
v6on4xqpFciBgy/xafH/kX0X/QWmDaOX3qsDUx2G2FLS+d9/UGSYGh7xqgdWrQNKYvmlJVR/rh+q
dUknMLBiRJYW5PxNFRcvOP8qwCiDvmov9cn2zW3GjJNNTUWxmG3BNEE32YGmKxBJnrgNlZjnG5u3
pvKiJzGaGs0leLpGcuOJwSGojYpTWOVqthU+/6rtIqPyHPIMTH+mh1VjJ1fjk4ShEHHqSa3yNaJq
w9Afda0UR0JbbsO4hbsn/ijV88SuroKJI2gM2xZSsPb3NK4bfxCnJ+B/WlfFQRmWYuh/EnpgMqvp
Yh8NDvL5v52/klqPxoJYL2VvKWZTnXZmEMDHvuj1WWDqysW21p84l46ZKET1dO1a9P90HPVO71kK
HAB0uH/aRsFFvF68+AnON00RKEQGEb2UF5rJID8/oSKNIHMBF4gH3ckRP4gZkBNcFsVJxm/9YAUY
XiIE4JmcrJGRDtuGeGMDdPOXZ2bJWiKBMBHs2ah5FI1hMCIN3blFUikxpQiETGYarIXmSGtekWja
J1fuBcNYuvvPBExywKNrhQYelwd58C4dYlo6/3xbkmSQYtxjMY4wbxYCNYQ3Tw4ETg9xzkHuZZRN
gWK4exj22EbK6DzdGU6rwJhtiMhrea2GzD/B5AgT17Tk49g0XJc7zi8QhVg7BIJSJHamFPA+jt9c
HFpxmtv2wm0fEXGUe3fcwaAr3cbZuP23EDqmMwfvfWII/gs48yzB37gTi/7/+c4HucNvzU7miwLX
+rUVzFtqGuqF66pWakgbCaqVJyH0v63B8C09nTqBxKQRJOUDPNbQiF5HloW4RWBokPqwCCaW/W4x
ETET4w/ApFmXHWJZbJcJZ4ybOAPUIdxeFAwmrXzKHBAAvCi4a5msEFmvfUmAxWNPsVNqha6jNeyb
6Bd4XxEz2ZGIQZBjQaAqpVbIW06E0PaauJ0261YGTnDe67FKk1uYuTcbINJpf00//4HXJdZS739X
d/bWLa8QQUacxG1RzHbOHFnINGNlrTnavx/PKrs9xfAloHY18mKnW4pENhtyN+xVOceVvTVBqp4D
NyG1wM/IS08tpaTE6YlCDOW8/PgFv7W4G8JXXDud4da94suuDe/c4KCWWAU2GSRnxZ+1P66rvtBZ
qM/+BdmQvAa98U4mb7DbUASt2CpgHeEyB+zZVuuDkAyF/VSRtRGcbC/81M5oOdEvlhKD4Kavs1J3
Zmw+nM3GY9Y0fCqLuvsI56FkCH/kVAxzGicSkOQT0Sx61ZrFY2pi6PAcIYxPCQeaq62Xv4loo2Ur
xsTXJw1M3rKjEm2IZE3nqPtnJtBv8Q0Rsb33lM3L4lyZhh1znNyf4/3cRqEA0PjsORvwQ+8OJpzu
Fr9IumzGp5KalrXnpkq5d2ChMAhGDJl0EY0KsP/KMvrtG8xLOZzBF1VI1+Z/Bvysu3BPApnPp1sy
YY+XAxF6aFa72tDQMWq4BicB96VT0scD3TLaa3SD6wFG+vZZXwAAxz+wMoLdSEzNp9CtrutHzjpe
mpGqM+cKHQf7x9ivezw3M70pZm14sni89t8zWOATQqz2zVX1tqwpBSXYZ7EedtSeSV00B5BO/dE6
mxJbH+9QNMj1KdP6Kn09qei8iKqEh3FrNJtGp4F2WZZjiFZdUVtynp+vJqkNZ0xc0zbB33GhLEBt
GBCiTBRB72W+Db9REbz0KL0MiR/BYrlnUzGd5JB1xCVG3XUAgBiDIk4m4AFyM9mDbeFgK36mY4Et
b2gg3H6dcuSeA5pxJ7m+WxnJpihDM8DeMoMFMVwLq4Q15KVDQX6i6xVgj0s16BKwkiSOlptuAcOZ
UhxUl7p720RcVaR72ilAqZB2DNJME9NWW2EvREZIRO9O5eswy0qqANGlFvuoBV0lud0bhHaOgf2F
9Z5B7Oxf08+8ALBru6l5px7vseMof1AOOxPL8huyMV5IFWiANpZ2UvdKUsTvC2ak3z/va57WwH/Q
NcYjAIYEA9X+iA6NrZKx/HYh4bdhwUYZFAJoz8xQRQovPwg1UvojqLGhaT/Uv+QO54DYJV4QpEsY
ZbVfBZELiU1qDhnGhQ3ptnpHUDRWYqwJh6L36feZYaMgNoF3vCxHgWpgLyILt6SYW2pudJWy8YrA
LdnEF4P+tjTETFSrCikXpBv356JtQ8SWuUZwTRi7SElO1IQcsbqQ/BRlGAJbo9NTjSN1RvGQn6sp
fT7HbmsQ5TXp7CnFmEs1CzAQXDLSZABNWFTI0f+Ykn3yP4skS2GXW6bL96+MJfFvUW7ftk3sWcKn
0O6xG3QKRiOpuY23vfhD8Pg8ImVL8XMmdf6ezrfzhbpA2167LlBjgmJLe4lWMV1GuAudFK4EZY/T
P3IpW7CQHSDpi68OIu/WZLuPc7wGXud5LeWw3pRo3aHDFKLRiMI/dqpE/9/+2F8VTO9a0FZ8kpDY
JDCtPZOA29Pu8Rdo8jpHicpDLlT+WNy4ZasrTfBH5zezqzYfxR4fb5WLkecL3HLISj3d963GOmvF
zv7f/W64JBUq4/rTR0usuWGkasmUO6dhlxg6JOBCh795n9b5U277ol5zwscbdbCdbf7gBpKeYifn
TQD+CCtvzWR59/qgPfi6JkFMdFV5sx4yPwitf/72LM2DMoBr/MiZmN1bDJCJMb8BOJxSl0NY19XR
3gMjzrYDRujn08u7bH3ddqZy8u0n9APLLefXXfhrQ9oqYJSHXJXnVGuMtjllJeBKE3Qz59r5Ngbx
1fwvtRXBtiBbrINJrHkpAd/l4RfsqGBLvDcNAhAl6N+20pbTQMqh7JatcEIRlfPwnTAqu4ldUU7O
dpKWZ837W27BwbTNSLTiovFr0Q+zeHnVq1JfHA2SfG18HDZbFpRhOKOyAfd+akwpL8ong/lNNq+Y
YoIZ5e/qMBk2Cbxl449dyDlN0JITfCRXHQBF+qtTEUaWThnSSN5C91nI/CwQ5zOAZrbFPeG2sUh4
PajkAL6VdbieSqXRzVbkk7cbpnOaDvNWFOKP3Sq/0NhnaAhyGj1LN3AyHCM5xPCSCXPTVTvuWyIZ
tcXJYa+n0j8CSLL8bp8Se9PMyIUp9F9LsNPIgO+0Q6xOtpUkoAV9IaXqpKotWYMKSEJmUUmZv9Ag
3uJTC66Alm5pGpFEVKmGPDd+yH+RplCG70eG2AYvldWdYagj7rlzyR3SdnVS33ytrp7NFWZidcK5
PxNmNZyeYLzEPWr+FczwSaSjTVG0et86F5hTBchN8xyVA4JDb+hEEHEHR0y/HryBpgAaRFfQxDC4
tDR87Pm1+gEjaQq3Zv9VouS4Z7MvZ7x8g6fLkfjHBPuV1qG4bw2YZ619JHgbQPfxG/V5JV1qjtbK
eK1aq7JtCyxKYvUsD5DP1ZPmv0wY3APas6hIsxysasmwTBtZn4WdefwH7Kecf8dBPpvW1zAbME3/
AiX/cEIH/dmRfnoA/H8Gal7LnX6GYVmewGFtrScFRju/tVtKcvapjtFS8KrlI/aC6YXqUG173gMf
bWy61RFyhnvWVC/pJGJkwmzd6buQVJQqfo9dRiQ/OyxSKscLGHytKUscBVq7+HKCUv8Ml0yR0W66
EfvT5IK+BoZs4eDPVH0R4BVAvAlTpQuEXQbMIWWnlDDAVWihNpoHhwM7l8oANmdLsv07SMc3lgiN
ZpZECd/4nmiDcOzkqGz/b6Uc7Zg9Tbp0rlu4/dOR0uFEf5zFXDVDX7SImbIUA5U0+yhZ+hb9X5fL
/2k07k/6XtiA9UslpQTqxKM3azJHACIPaSwdtOMyXt3a1u72SNTGQXZItn7lyz6LG59Qz6ri1TZL
QXPApuUgdON0SIYREvzg8dHvMwy2Ook5JZdvByXWT+cqpONWrhgU5KuJX5NoMDiCWYe4L4iK9BY1
/gEbldi4DXV+vV/nhB63tfxuMGhi/xHFkH24oj9aMAap6WqUQia2BLposicVqhUOdRz+WSK83lUf
nAads8XlXFQCwly25tuN02VdIgcLkDQwALtQlxEaIgU6InZAl80TE0knXO5Stnqj57Ee1Iww/c7q
SHKbaieszVnjzpwt3KIcAj7vLgMrNZct8+Q8mezcHWLcgwyGBH7+88cVKGYUYEdkZgRlBmxAQxmT
M2EnaAeOTO4Fze7coD07kPVB5Pj6im7t5TvvYWKJ7HmShMZki1wkbv9Zri4qBw6oPTDk0cOQ4eqY
p+VwadHfqOwWiPqsMqfg9VGnputMfwzQioUQg0JLteX826wh1CfS3tag1+GUHymXvBh4yqmTFZ75
HYZr0D/t4T7Kyiu/cczXLJ5rA8EMrrwdhi3A3Z36HPNSP1s52DbzBJDfRbYyx5PRShe7k4RGxrlX
noVvS0ubkq8YQwWgOcX8mlHR5W5Bzji3ngJuMt+VIlBTMpvz9eUw2wYC8jQCIheGJCYNJzzZrT8+
cWApvnjUkhgCflrPILYULJKTev/dO88Vqd+vgiU2lT5nw+1AkCIV5Wo/oKAvZU8Dm0OQwereHVaw
qUT/ohjlNHVA4B02NT5Sxz8y2FJ3qHrvyDap8j+r0bgYNx8UeigckSCVEePVaxwEp5HDTd+YAzQi
OQCy2pPL+aqy/Q33YqNCS+H8vAKLbgDX5ossq46PcUArdTmlR16cN39YqHR02MN5gax1XfX48fiN
mCOWo4i/1LnA9Sj4NeloGZ4LP7nvOld1qqrBqqFzFFZSClxImKcx6tYTcRLdRcOA9ZdgC+aVwcAw
8Hm9dCp4xVzsw0UIN6221hDUyDpG3jB1/yXpiA8Zz/zdLdozX0xozv0Or4f8MqzRTcy8+/lKhggm
qKcWty1hu3SoMC0AVtgo8odyb8jR8Az6RXgdccmbE/GigLkvr46N5u98LuA6qOit0SdwLROCKFlh
bkqxdzpkOj+VKWLIoV2R74tsMsuhrKFaxSMjm35OZ9dSO9JezqlpDT/1+TfqTL3pUFKPHB41UP7k
tewYfbMKsjcCMf8xuos0GR7qKCgTDfp9HgaDnx00meInbGwZ1LeDcytEe8a7MUEwCEnTQlfDdooO
iy5YsX5GeSwAFTqEeHGyykAuNFmPpDA+7fflcAmBmWvVv8ScGVD0YnGgRp83ioMfqEvctZsukFWT
RYgw56z6GpeH/g4PvmPEl014fRdYNHDPpBHb/9FbErWck38chkvMnzGTvMMa3VKzOoKtqX9qYFj6
lOZp4qIHI5EFaygqZ99qsld2g7lcUt9RlZsUqIqj0kgBNA4YNmvPc7YeSgwXkt2RDskq72QxWwya
CwuvkHLUeKAcTTlagYkpneSDEBLFRKtt274HtWEeAOZQRZ8foi0LB6vYgtI40m0YD6kGpdw/47Eh
JbDAcAsI1P5DLPWHspqSm7baqfAJVPpNksCJmr6+ARQKZXdaDWCHasPGbC53Iy9+amgchYUG4g6v
rsEZci/948SAbn4hKeheIMvnEh/dMv1As6VAO220TscNHo3aABQBfiL3d5PbTNZvUzFq9JRzv854
eRmDK1PqMa/QkQb14DKIohS6ThYo++6CAERCAhnDLjDz8MrbWOWzRbpkllgLecka5ZJ4FggTQ3/x
UKKydw+QP0hmZvgZDD2LVx/Mn9HN3bVLEMD3BSRtkdhjghuNBrGUlbYgYy+ng1h0d/dqsNHcXjNl
lk0BBFuq7Rl1sVZHp/26ge6Fmpl+FaxBf23jG/0cGXVtU0rZyf4Bdf0isFkdxY0L6v4FD61LnIxT
EEMhKzNj0fSvfLZjkM5vKgF4kjPr2KewfIECqUADtDrL8G0KmhSzwuvAYiWC+3r8WefH336mGFdf
Mhw3kqdGFVlUWZyT6g6c+uQ1p2ntj43+6QKZWyNTjLeN/cIXZ/eJXKxKaV2JvgzE9XVtgMjDRQGe
27VPG4oSmwoRuRS2qU0Oh7SDPyNVi8mG4nglOsQ5qesCqQqdFNy4q3v7Hq/c95e11LYGUvA2bJt0
K8Ec4KUH46IY+jmlh3CBxjGbzsmu6YBlB3/wLjSaRUjmiMapHdvKcblIQCWV2cI22LCn8Fz85/MC
R6r41EbnWgX+E/30Q4ElcOVxPruOHlH78WSdkpBiRHOjrCgi6aG4O8Dg6xyx/dz6eP6+PUrsV6hT
Debhp+KAdcq4UEdOyeDHmKWhvq5E6P8S3s8oC1OTVvHqy0B1Ihoe0e8TLzRk7F4wROgbtAbttB3A
/klBcCjcHbPQgDvnySdqy+Rh4sGsEFYwZW0QBnNSZhIqGVmW1l/9gBuxYtygBfqtCYJdGezfByaB
ZntBSiyS3PgH9GlHHMa0mzCB5+vcdvJMZduNv/InQRm4D9sdRzvYmxMb1qPpb15AmwJ5xfyu3jhq
nGgIOY09I6ZwhL9yJem+QRy/Staw0GQTfw89E9Cocv2HssdBZvQjyd5QLPEY6YKXWhlmdlOPBRij
OncSmkjGuEYFhWxKfAmSLAK5s874P1Fg16+ND3YSLFU17HDOtSkLRpN405Fv59qa9grGrDx9kHE7
FNFgLQk2g/of6rfy7besQwY4OhNIVMsR8NRGUcYWcCLU4X7qwwBKV7gUUn2Et0o9I3hq72UD6qTg
+m3/jwyih35dfOLFcZ23PRkhMzwU5T27OtPQ+YUSn0DCk1avE5UslEbVDLY3S5o2wqC6GUODaKCk
Dr2mWee3rvmJq9hObS2ArJeSGCbFpctCYDzxN5oc9NnldQYuwksKBaaeQ61gb6HDbIbLdnQ5+S2W
jf15loUPN1z98Xfc4FhaddVmn3XXFD/n1ns3m2zkL+k/3DQcdLW0IIILk9d64PqeJzmFxL5Ghz1R
f/OribYB5rhWW1E3tTUPWWMOH20RrmV3r7DCWdTYUQyqaVGOJZTBvsbAxzXPqMGLHhxXG5I+4Vch
mT4HEqiFzZH0YJxCVxJnDiSIODCc1R5nCSw91AxanyKVk4NT6txEr7h9R2detQRZW5Yv3do1RQk2
7tYWrrVdoCmeFLekGcr03fVKDDvrra4w4P5XXicT0HkaWstMLqiKavsujfJAgOFPLszs0tGVxN3l
fk0rEBSsKsBF1t6WIF3cdSxHmJQlcDGd8jztSZAIejboQ5D4Kc515BEZe4pr8HxhrbpfG9DjgRJe
+QWqD/z8Ymfr+lSf2HVTRGwCxcbBaP98sCW7fuoQv95busvdw4DFFj0ZrcK0SaVRffVBa30xnPyY
QO6/gfILBMMHDTS7mmMiE2FJ0lY6B+5Agzi9sK1PTXNXMWWTOOfGACKZxHyJEPWihKz/XFCll85/
P0acV6YBfP2Q9ZsGGrfPnNoUtQVAC7xJhH1yXn8ur/9ea8jAOu10mj5wMUlv01p8nAvXHmCTPVBW
qG3Q9FnWCboDFcyj+VdKDL1Hazqnnr+zc4g6H16zISa2hOB4bcE/IHIJN7nDOCtUUMjx7x2mG0Ol
OToJCrRqUTdQNGG/KXdC5eOerulXmpiYRn6NEUzwzL3Owp10NPTUV3k07LmRk3w71Ce5uiAwHff7
5d9lITSdXxYOm1uXny0ws+l2zToXEV4WqReW5aSsK5fsfsVaKj6BVqHwyO35A5/cRjP4tDM/jJq0
VV6N/Ma3SK8eha1+HtXJNNkXH7vAQsAVm/jWITXP69Et+UnyWUkU8czlIOpMmcqEZU628ZYaQkR+
6tQw4RDsEwsvYdkUWgx81qMmex3wFwzYjpUFDW0lctqi/j6xHQz0vYrAg9kF9EUHRnJwhkvxcaJw
TH33C54jaT6QsYcV5CIxiRKOBNRLXduUIXMVXN3lXLqUYaUYkiNTlouIW8CjtxeqU6DwwTEqdahz
Puh573rqpM9NlNM2g4Jkp+QEX09i4aiI6cSTTWxXH2LgpVUbuzUh+y+mML7nW0FjWjRJdi9NEChO
uFlD2OWAQYFX+qMEU20koUpANDhzuO66f1upTVDE2Wu/9JTJlnJp1iPjYxBdy3fL3jq8EgY1aExO
I1s/Vs8+/XGl8R6FRYeswzyK0eK9TR21FUkriOoRDZeLcMDDJ7pQy+jnvcjZjluFTSNpsC0t1lqk
Qi2DAWeHGJTtPXQMHXbzQsqeUsIS9Hapk5VKPhN2piqRLFjvwVrkAxq1H7vEkKY6eyWd5JFZ0AfG
deIUQrmwZvPaXr20wKHS70fyTvGN1aShhh+X0jkJ2OIt2g48blTXNAo62KguYpD1tn8PTgyjxs0D
cvHSn0XqCElqAmSfQ0RdO+yy1sLCyHAT70oJbWnXfBZA5XGAsHUZSWxIy1r+le99y38KH/f6kht+
+u+RsEPXTc07tTUgQ0kXDYRTveTzzv7d7jgvpF7DBigNdKCiAxrN3V91MKtF1DEccipYaI0JfifT
Jpnz2fr0tfg0/SDkJqYQQxAu3Y2stujndHEsGFNq8YtpNo3D9/KTbWGkL5ZBZIrgEByt0iYjYDoK
jnZAplB3FSxFLYgRj1D2gBXzRGlVEGL2MYQniOkMXqEFcH0Q2qg5pmK4N2uDcDvvw6OHHFNAwjk/
NDnWPBacmQk1bjFEF6/6H0ivhBVv5wOkDWWqND+GtAZcJhLc9k3KVGYETzlFhpJv+cUL6YIROh4Z
v+SPxuhhhdRZUccub2UkMuxCSdpGpEx5xRXn4lCjgGRfBJdVJWmCnwCGmRg6bVf3C4bbrqu9Bc1q
vpFYDSQGD9DPMSAAUjdVT+UKmWIWxdocK7pQx5+0OXmsZmXL2lcopHX3rLaRaSNLWu6Y0ygUf5A1
ld6GP+Z/juThLAbkpmyfkG939COxqUKEOnhQgFSQNmSOc7mRID+6zr0k1sgIEJzQ14H5PYA3HxTN
6j6e/f+QudcPnfA2WnlQ+OOtksKCdqc3HSRRQgBgfCZXufmdb/CvGS87o0oExkSG7UEFKO44FWP3
1L9XosJ8OZnerfS3v9d1Y/D586cQhXWt7W03d25gZ+D2+u17oitSurun4oe4+MN/5bbIZN0s24U8
Wf0PvEzMtXpg5iVhfHMoyGd9HN1PlmmFXkIvzm4FcD3i8jKKmB/FqQOWR7GW7bx6wD5D4oK+Ff5z
jekGmuZECIkydYzQUP0MxZOhN0bWzeVR3gFkDgrzrafoh0aiAvSfDPl6vo0caK6SFIheY9vtnRbr
lJliDnzN3GMKxBRl/xhyFdT46edhxoqRTp1XkKSXRsjhBk6MrVwirhgKneldlXdVuKPb2SSWRlJs
HKcHK+ErYO+G7gIU8NnAXtUt0fNkkAXIg2he3Sn0fZ+tNgnt3WDeRIhmOTOKBdtz02q+TAJdHeuK
usXox0MgJzfQxqDPqkJB/tLfOI+52FjdXoD//pvMZTq169HhtV47CgfF9oPrt9TQGk0sTmviDdsb
Fyskqs+XrIDl5sV1H7WEjPJebBI3xkf2pgmwY4R5Uv0tUBcE3GFy3Fi6p4IORBSZKD6aqgJGxGCn
smdHjGEquUzZkCpPAnUFaOgV6E+x2BWLARMMTlZyLrvZvtsiSyLEBQvG8iSQ8UQYaZX7Yk/hTbHy
1qkSQdHBQ13b5UbromwGZLY0a1SZ4blefohpbwQd9XeZkQRO9Ug6L/zZPThR8uKf2E9JaThdOZKk
RLzS4J3YFayNiPaY4bi/QaB7vC3AAvbRBl0hzcrb1+zJIROZRdntECRSenHmK1kxeWxkXX4irM0C
SAmhv+vV/KXptYI7Uc+3oA1EuBNMkKJrgyKyucJRwQv5tVddUbs87kIn4wjKy4LDUMg6zwcycaI3
dieSOvXp/oN3IoB1JYObsDyYpi80i8fHOtksJghQ7gRIex1aRELA159oiYvIsSnNbzbfHz7NzxoT
dTKMu8bQkUXATO5vi/eOGCIK9KV4adQVcS5LlyQ/TrwM8Q277ejFXZDeP6TBpejTQUHAB1yCZFPX
i9h5c1QNpyVFr6gmW01Ri6t0VzgFDLsraOG/6Ft68b+8fECt9LXqahif0BR/9a+PuQ9sr3hWvOaY
t+6kr9hu5ukIUgwALwqW27cty7pWEExdrYCR8dFsRk7fxC2970V48acfb/LHeUHTwcai5P5sRDZO
6byG1kp2CB8Louezm3bVWspG9d93+Tl6I3sP75DZTRXvXDpzBMtfeolecGGowXFTgG7hLMTsivid
F8tzNrBpnSkKzJkDCOc0v2p280uxbfJC5TVb6h5qB353Qn00l0ny7PFVhJVLp7t55pYUnoFXdSrT
A//q/qWPeeo8LwpIKjw8wmG4SjvM5KNItW8g9hiLybfCTckfU6BPx2aLF/kyHViWd4urC6+MvqK1
ia2UV5vglljWvIrk/6RqbPdExsWptp8HcI8Y+TrqJ6fOFdasN3DlV9s1YbW9p9tNFnLn/OhWgyWj
xLMjjCk4HXLKcAOIjbflrdt4ymSxzuihxpLxD61AB0nIql/VEebTqTW2xC3L97hBXNOruOZ5vARR
zUcIj3nC/zPVGSEoZPBAcEQ31QMv5w9+O+guxEfReaASwYXvSqK48t9tkpNudWT/fOG0bQdMq3M6
Adf+yZf4vu8YIdOw8CG+6ezllj32ayCIiq2WhWJmFsZmIdyJEKPcejr/ubFO9W3bXMluOT93IrSW
NB1RtabpwQHrbRRttBLXXj6dQu+vJ88c95y6S9tn90N7A4gMnJyqYqJQPUZ1GoDrtPUoRvxy0X9c
AGipX6p4275PkpHcb8GdlsYG2T87SrQo0/Ctf+D/iebus70jBjoQOEN0fRlTVr+Q7Uf6O14yfbPz
NoFsttNDcCSaC6CkUZnSiCaNPmPA9ehcRhIt/+vN3U4c8enD9/4bQwC7CuUrl1IAv5zV1cIMHerX
EW+h/A3uAzVyIQZZrB64RPiWtp2vkvVvV5YEFt/CeihgVYpPK/gF8Q40CnfIbTRSkJP8Wmsqnc2k
DkC4LUhGT0w0VONVLRO4i0mizB2QTK+1eSXnO9X+1OBD4aWgDcX5XTWAoLdW0uhhm1kZn76CK9B2
dUuiwTUZ3rwzwya9jOtcMoSkRdlRn1qRFBOerEx78gqC6ZxP63gSUsyut4kHRPY1gdpKl6sIDZEw
VC/+nVgzadLCs7i9gol8JcHX2Y2WYKcKU6qGQW4e8BvzNK44rA7oGKt3vPZ6C/Fz/LdAoqFBb7lJ
kXLT2Ea3oemkzIQEh2+N7E3tLNh0apTgiT6ASgtgoWoDuuFuUkWQBsTptWfH/AIuNbINrwNpgneQ
egIJmvnILnkpO0cO2G6ZpLYFkGCEl0Let0rSC3T8js+ORJMEpZmhwAZA8dTmlf60Qey9uoSJF03t
afo1Bryu6fGpK6wl0qWPNyEeVjnSkVq6ireQMzWzj88cetMrYZJPG69K5OBEPBbixE/ZXFn+gVlP
Mc+70Qpxpm/sHjR0Q++ZTbKse2Kq/y5neqV6zLWLP87MnNVme9TO6uSKlrTy4fwgcytJvn20VjYi
lw1spk5LQHhowucWqs+WpPHQ96iO7ai1CWK5Lks551msWT+t4KxpWEVhwxpH+bHrvIlxdfwOzJ5I
j8AiUF5w+ye7DAisTR2VKXjUCrGQLN4ZTxgMZbzsrKP2Zq/EScx1iuwVihuhG8lh3OUbA7it6gUK
GYJ6LIVXT/Y19+KYj5CRp/Gnct7h6ndvKdsnGL62YOAVcdzawaPQY9WjxiHihv/zqFKUEbqbfkT8
IXRaK++BQQ0ofgOGzF4SHfHAA34GcrPusEX3J/EiRc4NcHCxSnW0glJng703l7+bsn6BYlph8gjJ
+iNl+O2WES4jdcr7e+gOqzaDD1PsyYhEUQqj6N8khSQ6x4cDhtJ3mq45xk6ZQhtajXH0v/lpB/sR
Nvm2iOiRo9FZOubUWf+qofhoUD4FJXzw7r82HDuYaqmvR/O4qz/VZCgY8Wz3Nc7k9sIWmKV63xMO
Rj1iX7Z51tkoYTsixtFLWzy6mBYH8QOOjwSGuC7b9HZDCGx9FHg1oEKvS3poHTlP99g/gdMRhtDv
MhUMLY0KHVj9fvFazfrYzZsPJ1P+Ex2blGhaAXXiI1T4cCjaoqhERtqLtRIRowVR+5WpRQmOvURH
eVnj0MAhpQYcKVIleGngNAYSbz+2bsrzDiYdSycCHYHMg16JCZUqlHu3ppQWatVu6wDeX+dGOx66
mlRBFTFL0eSaTAICUxuC19k/JJ87CWYZHwXm95MYHo9Df3Cnm4FTbePfvq8KnmrS9tD0xZVhI71k
VocStACMsiiIkvlSm7qmg9rgz8hiuFmdJifrAT4o39/D+1Dqpi5ya4xbobBd7JirnepFGDAzRWrg
wELC168FvvfYUi0P6anDKQeytZmh6mzbP/AlchhT6ygvvXYD2xbB0l6WFb8HVcqrG5B0arjHcIqM
6K8zl3SZLLbyg4WGJEzgvmAYn4JvAy8nBREZc9Cb4DCjX+VlJWb+HskaFicHaeaySDQcBxZPgCfR
zqDZZsK4AGsYdG7fmdGbfyKkMocC7P4SA4ww+5YKOVaXvL64b3wef/apaLnzHf9+QCdRXOgTE/K8
T5I3YiU1ObO++EFm6LEilBENpByRC/jwjb23Ebw21j1ca89Jj+a5kcXUChxiZIm/nqZ+OnNUotRG
NTg2Cqc+lq0tV02/EKH+ngVrRZYAcUX9gQDvQoRdVQ6q52NkzWuNQNZwUdAK9HTBWXwrsK2Fc6kh
hz5q1Sep0uxD/iah1jc1eTrrn1U+TwkUfkNqZv5ZBYe11izOT/oR5olhA8+sJ8HQ7oQ2+EtU1wDL
ZhLTgy+yk/wJYfGkH1Cv1hoNflKNohE/MGsjcGowiqFlXI2beKyipkwaXo8RavCSdoQNfrQYPemn
7PvvPO/yjKxsPsj/LugPerSbmW9PufQX7XkIVBYWiAFrO0efFAbhLcX6RP2XUrH4JocYsCRSy2vj
36CtYve2v1Ymr8Uk8mBsAyYYGcwyJ0hEjGyC1dkGbQvt+Uu9PwwC+29WTa1t1zmk64Aj+Uqkxn2J
lZ913gegO9LCZtOl9K+7ZdH5thOPTThXpg6IH5g038pkS1US+x/pb8oY/sD7JRsWxHTl6qwAcK3x
wG1XHzGX0dffignjw1DsgocyLs07reLajdeupXwpVoCWlq+wXJOwHJbhRo9WdLUHaSAnh/UxsxPR
7GIlPlAjvpR2+oLqbW9sdEKNMvLDXamgbbZjycGM9VLFM3qvdS09sginQ+BJnnb1PATU+1RoXGYD
WihRKCpdtUjmTU8VWTcY0Wdrvn3Ah2d4iZx57vyg+vsU5JW4HrPi9AtxKVuOX31+6cWWN2hP4n/A
EN7SPrB4SGLYs6NM6lhJZzrS9yldNYdJFhNCEp0dVy8Gdlu2pbPCUoMCca9LMUkGjVDeMr5BEAfp
1hvBQBOqdtyhEtwxSLvHnuqOtNamZbRDKHTBKT8G/cDZUOHCH5czfggtsLHnAzng4wsSNPcHdNUJ
FbdeohHajYUIA4tZOCfjZfOlYDjy0rAoncJB5tbuNlmxmo96aYUlBpZoItxU4XHX8OJEH/EVjhbg
io8Xg8OO9d5hd7f3mca3eR0tC2vEeFDXMByTpiOhms8gv4zllX8l1Spay4NpsYochCtixK5gYZGy
RuCGMtYD/AZlUZpyJmV5nv9DlwNYKOVQ8tovU84fyxvJmWuo+IrEecRwF2pGDM1pht+ckhAexNUp
Wox5rEUWXuGHpYG2sCalS2wWiK4bWh8mc0OiPR3edyhHEmm5APRPCu5JvcDVH+Ol/eIHURnfos2z
TTH2ninhDqepzPzIQ7BFWVxvG945w1Ld6YmHAIdNxZtkwp+5N4bYVfs9EZ6Piiz/L0/sFBDG4SjI
KBcd8wO8lGPE23ngTQqDUrwCHpB1r8eVDOX9ygaggRke7/RUv1CQYtjSaHLVRo1bl8R1s5aRt5HG
DO/rNafO5De34MJaJT+4S6giZ0EgWQ7A45m1c1hL95oTrceXdWfKRVRv4tzsnDBtYj4Zxvct9IPU
+0DsYdNdymrfRzwiREAGi/T5lrnlp2y6M4NUEHOgpktjbmgtXc2ZjNl/wKp/m7kk7m/Gz+uqk27p
qVn7T6+iHpVCR5OBs4iSflNDDu7H3APQ5WQvJYC6DCDYgKeQ0H0aP8LRaqyQPI1V84SdCNm/TSCj
khiZ1JaIUPsWOZ9ovoz2wtsrTwrSenBRw2Or9qD4wp83lYoALnHkR7io6ysqqvc64cf4WZSFN6LE
B6aulPL1uZwPvjFMj66DqvdzaJrQFND9U+ngJdshBNzVmFI9aSkifar2fq6EWsUHQzyII5TFTUju
8UQFRc4aHoaK8UB6n8TktEfqWn8LzVedLXYeJ6BSFplsX3YfR4RSNLnDkUzLzOodgTtsjGOyA7G3
3zG1WtXVJgO2QjvSOHd+VUQQBMwA5QaPAv35D3qM7OzaEVH+UIHzio0WsXZN7DpzA65NbuIAUNeD
tf6iZSRtGd8JAGWj96VXDgFS4iklRkxz3SYkz7h00hU/Q5HDqw971Pa15BL9CxnN4J/eUzKhtC60
H8y1Rf/pWFRi/YF4FXae9WYCfb5m0SdTEOfuzdPmON1QW0D/W1Cb7qLaa/5NBHb8ostXSoy3tK7T
s1JpifT8Ak9rIrh/kJ75dI59kvyovkHQDIzt3MgWCO4F+6Kkmgip2OIZArgTTA0Az1mGnpyfcQjm
6GzoxOGhHE4221ef8NbKFtN9IrP41u/s/gz4xo7iSxc3OByYLHEo5lDMNl9KoMoTxVH2jcpjbWiO
3hGdhoQ7tLQ7BMGFGzDQ0B6uzMYHboK5olrQOwzseT2Sv6sTiVEgj3JQds6+pzLNDq1KiNPCmVYn
bJWEkHEumx3PLTi7jMoFXzOOtczJ6XMvIa5+FaX/CjX1uIbVTuHVN/KgK/2Uwn9IgHvi5NrUKgQP
LDhDNNnsFpvlF8fhnWokmItUpG7DX6O/BGqpPmu1gVm+obnOFjH2iJvPWzIqwh5Xkq9jnnoY2LV0
i+Sl4iRFeRpSxmfbpTr2++WSwhaeM+odgpxR55JyeXrigAo40SX0b3VKDDuRtgqtCEJ17291I5pn
VbkNJZEggzPZqkdV8W9DHfmsfM+KuaI5rWev9YhoaaHpWnFftl/fBUIqu4gqIDYTV2OhOq551FoC
WhWuKp4KfBXQE4I6DAipbNW8LZfLrAHJB0DY2Ww8Qzj5GGbbZS3Xv+SotdAgsuHmXNwzdK0vGR+p
EaCit+SVKsWr/vXktzH5grN0lns3Z0C9UHR6CAzcexJrljmukgY96zf47DkDbvEdi2l4OKeMVVMA
KTzgIh1G66qx70i51Y5JQIjWw6Bn2xUPYx53hrGpihPH8fjo5rLwyKjwjRSSVwUG6dBOfAdRTZd8
k9b4O6fblGntwBq/njcti/ztCQU1A1+5J70Nn9xmr0oRXoT8HGSzoo0hoQWUQhtrSunw9C5SXcHZ
lBV1n9Sutv9niecM7BXAHXyUWuBT/w1vfCEFNinT7EDRDhIGJCwgTwBJHXZTRt4NLgKrws5G2Krj
kzN1Pudmz6WGm34wPfxwSUk+vdpoHUU1vUqOzHB/P65EPDdWnGyoqMommXf/GUF8kuG3laLG4MWK
WOhh/dpXzyL7mqO1Ul0/O7yUYT+oys9/ImruJ4Ej9f3wbiGR3VjSempGuKeBP82jmz8v4cXG2n4B
6e9NnJ7S73GGd8A30ajpyt/ShOqVo7CvZDuTsDupeh36tBh/BmCYVRXyaVcQNGmkOnfmfwm6Axwh
L5E1pgbC9dex+94JxXZxYg4jX53GT+vyhTOcG96aBNJhNriGcbR4sm6RrycrpeuBD3bSJAKRPEOZ
XoAMQN6IQBRNlQShKAh1nqA91pbEoP4XMWG2/2hmAygC0L9z1Z9jSzL/2aP8zQiYoqSSnXR+xTRk
IJJXjuPWqwEK98D/j0OVbk6kEagJffP8NrQvYSKzlshltKGkiIY7LNOkOAUy+oFs2vRW5Jhot7lO
KGSvzIqoSnPFous8JZcNV/dslVhXFEPpkAsLpH8Sk+wY+GdErFWUaAA72fAMaOCqZJo6BpSnBPXD
6NN/XPZHSw3aQR3Uyax0aftQ33hdFLEZDRU5ij+bHUmbYu0IteS+0btJzitWHhvnywHEauBPXLK2
E47lo/PTTAtbfaVNKI90UJAWM4k0n6kMzHtsxTBrTWzA/3yyGjIKjdhY1KCgPEycLPzfBAOlJFcu
WzfxjIBbFXernUZ2q7cHY0ZtxUKHyE5zE+CQ9a+e0m0hY3ROsa+noqO9z39nAj9uVs47qX+eCIVg
wol2Qb8epUT3sqi99JHKyUz2R63PeLwCw+Y6E3171WGXDphGgxJEFWWxtIQKFRzQhsN5J3si2SFG
K0atOdaxqxj05HFr4Mf1KYQXipDlURA8ZC74bylNA0QSCRuhdU8Nu+zsjmbjQJAd/qPmspoiV9Kw
7B4ZaBioeF64GK2u+580fNtAdaLmz5NwMwPEecMI7TPOp+MjoCGE9vCps9QBbd5A79Zua23r+SJc
3CsKJKHCNGxGTRLjnYvg9pXVgmV5diBzaWWcT/V5A9eenKorvd73OjCK/Olnp5ycHDhHRY0PR6oK
q2dGlTS8nzAA49dox3X0eMW1K7gxXum7AJGYFidRfjOA2703elZVk1fEvByP1mI00d5VcPDmyqE0
9pyk+2kIN9OlwTMkFCMzh6zhlw0V1YmZKoYRfItp2IBOCJIsZVHZdxj2ZrwNHoMzDBIPhlRcjV1C
z4jfXPiTGzAoi1ny8fkDxqPkoh07WzW2BkA8TKV8BwLYkvgYhPAdFvX54zLW4Es7628+d0/Faxi5
rx4hh4yesstTxgAEqq0umcSOiC1nn2MpAn+GqNRvQcviY+bOFrgKVEHLa6t1ZhFN3+fUQZlLMCCV
YKB70Kn06RzewuI2mnHVJL3YxbZIYw6c/KRxH5i6bi+vaFpEDHuCnAewVbL8T7Z1lGBT62hPMgBA
rDK0RUgoZt+ARDqgU3Ztk9w8MIB8HtxNGvgugQChkDlvME9e9Ps+Qz4JNPSs77JCAqcwsbp+yvO8
tOpqptMqXNBSYguykERjrIK/9xQZu7OE1Z/uTaHHXbVmaqo36BDgDijEiV609p0sINE1qaAigM0i
ay+amn3VCP22fYBjPgRj7U2+JiWCPhcQ6ESNmQK76anDvbOK8fbrmNnnk9p8bpAgJ3BHSjAEJKYJ
g7sOg0avNyo/iScPQZEBQGtA/lyKFFvhJU/VzPYOvOq6nJ7rgrA9++q3rA2xJn0Qo/OXYjutgVQY
7b8AF6hDftrxmw8e54Cj00kH/7PcGFFlKWM+e3hr+LmZCA4tQ6v7/WvfVidrHgJd93hcj0YbS4qj
kMwjTLxi7KBNNq8bJ2JAKVMz3+lWuKWze7a0rJXSekBS3gt8wOTS8WoTyk0A00HSI+4C/MQ/7AS4
nozVJcFbwD3xhQXAC1Ime2lvyGkNw3ICP+FZQzvcCayblMG2TPzzT11hsgCrJktRmG17bJCu3lWe
afTOVvAkM3DU90QkenyvDMTKn+nqz9dxXbDz5wtVaOQCmAZLxnNrmokc+giEefgPNldbGDhBqhox
nsg/Ir6OsT95kvORB5qyFc/DPW7IJaxP/WifcyJAzWo1pO+yXI9DyoMxsio2AsSLIRpAk6uxKty1
HP2moTpOLYOYC55BnyWuAHlH0kbMflrMD4SOQ6bqVi+ONM54IUMkPE9L+2GoTsQmmkDu8DfK9+Ot
YH2mTwPObOGt47fcN33Cyd1ZEdVzZQSvmyvQobsz3OqY2vvFy+rfuCNL1u9OhDi5IwuJSNmpZ6WN
5GP69O3w3USmSg67FDVtfd0Vu2IGh94FdAwaf4dS944yAgYE9JrwGqDwsu5hXwKGTqlzZhzlpbrW
uodjs3URJ/8uNa4jSQA8p0qlxEOUNpnBPRKy/ewD11lteRNmZZv771aIQWshzwgevMTXHaAbP5wh
dlz+DxE+32GsgKfg4ONoj2i5NCBEUG+fN88sxHh1pPKIPP8o8qcXdm1VusnY18+VCaeNQk/ADCnZ
J4+Yb5wZsz5Y1Y7456D5fveUZrFIZ936WPuFn/uLy34R9vjdQrZVQD57epPVl2G/lGgetBp7xAw+
utPisVr7CB0OYoPJAouAmAM9X/h9dGCjWmKiHKuejbD/63J9tR0NwXIRRe12B/tlp7t/1RdXpsHY
fcSqMKtZYAwon1c2BNINiDJEPSbEAtT1d46ZsUlfUJTyHaek/8IqAcamWwy4ctACBAVGqCSLFGmQ
8YnW+9jeJy0e0DzsE3rYzTaDNqz336T5fiaKkt7g4Ld99tdQ8B8CxebKK/GM3bOWFp+goVvt/r28
ITIIv42Y+Ctw6pREbiI+rrNr9MCqWpACU6K0uwI2m62U0oG176vllQ97dNXUzFmtAU3CDpqUuqZo
b9MwQam0lIWLPd/VVcjAb+YX1FM+7u75yzQLFqPf5QiuvrMO9ws8Cw8BCyRUdhJ8C0rwfO3o20du
EX7tumBhMcMW1mCwhHT8kKbrbx9wTix0hHep3NCSUgXhJnJxDXFp1T+CZocXhZii8ZArizEz456R
sQeZ7lvYzmPSSx8hp5nJbkZ7Tt5dxCs92lfaRwH8lxGq+CIc7p5ZghqyBV3fZ2nRpHi9ekoyBfiS
+YZooOTZYGW8YvIpw2ro6COTA2VxqsN5gKdCBp9VeUFw3C3l+ytdZ2DqyiR3dctTzM5icE0oHzgy
avFFmo/KTjSMfo4uEWmQB5MLZBSHVP6i40Mpld4yOYUNSjeT23QSXXUiON3/sH/V5U1OasSuq5T7
E1+Mx+X3kVsF0E/OpSMqXg1BNA+VCu0QpJDb5HT/ZqA1IHg6lAkVymq7IFn93Cl46vVnp5EL1pJW
1tcblyhdU9K/RprBY7vbq7jiOGZ1R175VggwRmQNOgQLks/ho80mn4Zi45UBlLhT4Jifcu3jMpc3
eA/GKMgJfrWr55sZPkuT03jf++scGdACxmE/LMxAbmrpqZ29uiRbruVExFob7JulzVFvNHg16RbO
oT8sesBzBSYTNFb7rj6UO6cyTXoLeJmis7B9w9E0ByIphdZCLRvSd0kUwLPvwhTfbu2xF4ecvFzN
1z50jtYCUDAzDgdygsN0Shdr1EN6TaWK5DlB1YtRwM2s69WdSBt36Km/u2IUaR9jAvAoa7JTFKOB
RGig7bvIGQrpRJWib5ONwqxh8otBVZNmkzKPGj+/N88zbBNWASRtNb7yUFPZYBDMPFjt8QRG40gz
yGV3owmDaGeM3JEWplFD5lBro4azRaZePnWh0fonZ2vGdme9iBaTaxVV4vKdjOeFUgM/2tjufMt2
Zm1SVzpw97vmEwxUXzG1Ypao8vOqixa1kL+g33aeyAb5abkmGFGfOMxXXV0NZknmAbKTKF9MDTMX
Edc90flNK7ow5Ved86q26ago+atxxcuDP6pdO0C9+TcXMovCM427AuWZIVHtu2jjVKeJjdZ4pCnb
EPSppr2I0LLvw52Cu4qts9Aoz4m4aj1rruBdKilqSaWBz9KDNl4a3Kfy+5mxA3ETQlfgHFvk6tyq
y2ie6qhDj+bfdR55+Yj0C4qUlXSxbDHCckh+deCwlbfoN8oxEc6R5OQcaw2JdjqJmfbjICIJZSjA
1/7hS1E0OT+DvSMi9kO7aRp8kwwKS9EqkEToMp+3fub2v7opKcTYqS3jAcc9BvU+p3leL8Iy4Zjf
H7iloXIRN2baBts+wdPpVfLIB3CL8xzzIHWISBgLuU6qXpuExJlXNdGCn23RM+5JnubFy3CPt4rE
QxJtgQcy5VmpD9OLFiVpJcr2n1L7p6RLf++F7n5qvf2qlhA28K80md6xtVpc8zpmwuheqXlv9a6b
JPsbPgtTodUSgTcXAap1p8V8QJvOIcl2uTST6h2gTUYsXdnmwCE6EV+RwrTGVodKIZ1IQjBBIB4H
/3fTk8UhQHDabnF2l19sVms2OrQrcDZepFwdK2A2TEnQvQirMgxGXImzb5Xwqzw7ip1ed0F83uhB
SvcPvHhx53mdnw6wTL8W8kgqQEOTy4Q+JJu7XUe09wNBvQPMF9SEJ8Gr8tqFIHuoEOiEdvjdknRU
1yOQXblcPtr2t5b35dstNmyG0W6kB1zTqYKuQN9eYRSIDWFF3B8iv3OXMML2OrDzDLHNv/aOUmhe
JyJUuIcg+jFYLxn1cbqnQRok1hitjgKKwzLm0rbfeZfGYQW8Eu8N1n1CgKMg2q/dWZRt2WuBiyNw
yCMx7lv6Sy6xJW3X9iL+wXLVHIaTrXaZbcchguRFEU3QkbLOLA6HRLMtPkUv+NMdWPtAJqrQpQBR
ZdVFdzuxbPO8L/d/EkKn/Oim9Qjiy+K01FxkQmnNgb3QoUbSioNM5Ir82TZTX26tQHpXdzmhnBMb
qWR/Oi4fIoaGEdqYO4q7JNgZZYh9lcgz0VW9EVWamIebjcEBFK7HW4234ui1+95v9QGmBQfiWAe5
uBOC6CqR8CIrfnmNH1/YoDj+nRlCho6WvCUT0C/MZ8mjJlh5z41oGwpeXFIUaAznziU+QW5DJUAj
QPnGpTGhyNYAa9jVUy2fvc+qitp2PvvV2zza2Wp+q0opk3fiqptko7+pP17b9Y1Jj0cEThgzef/J
NJy8w9PYjGv9KtmPIxmUvVwywOEIqQnpkozZYKn9tCAiB7WEBbn5yEgvMIDMRMEFzsvFrBSzj1do
jZGFmasQZ53XPnalByvAfRE/26ai/d8gx0rqpRLpUJuARVFPmGl75I8VHnMidWC1EVXGuCZmJz8k
m7jx8FYHN0i1ZXLDxjBOiIRuvy0cXio6ksBRdtkZKYKmuVvUG2+DDibVIk65jHTF18AC7MWA0slU
wcwAAo8/BJRCf7iG2v/7c7b+siwHHBNWZ3U2YPYQC0NcT0CyXVBw/nnVi6UG+WLmEsQoFEQgRSEu
2eABd+Ku5Q8CSCdae4aD2SsS+a04/aBR298/Fnq87oYUsAxHzmbtGC/Lg5PcHA4x7XnPV9LH3q4u
tXEG9mqy+MD5zlVony471VQ1uqJ3gzdEPEpKV/zAERCpCYQfPmx4tvVFxyoURJXmaE8WrOUerCsc
K4moh7mJYUlizQyguHY9duo9tFBG7QaDaV92orDLW2llKeo9q260p4kj9ZdUBVVjK7UNoS9yZmjv
JuX+25DFtzCTxsEmtAIiX+LnD4ks3kCTqdlcZ7WWfbleQ70xl1DyuQCvOQ3H5ibpU8DKv2BLRKdo
GqApQ3rDzA+STH8hRy2X5HxCOOW4FODHcg0QSOgvpxrIj8SbRdrc9zzo/dMnDNcEfPPuU15uvykG
hyO32IIAKftSIrRgemJRgrhGrOO/AqMcMaJp0rdqhW7QTNUQXIRIDawR0umRQN1bAZg1bAM5QBlv
HaTAz50peGI3aPSCs6vAyd4TQk9K3N3VxOxYwWiQS6nTn5Y0JWNf+aABvxFvEPuF49LBDi8PIwbz
9bz+/r5GijY8ic0AQT0zDDMrZ0BcgUBMdDcdKlij3CexSmfrnrj/xac3PMZaM7dK8v+6LYW1yein
6XYoGJjMxpSflf84o3yTucQdfPft3HhOR3YmOUVkg/KDkZLrFd+2ef2GNbUGOnLSr+s8FGasOaJQ
SHgfzw9PKtcZJieIM+tIzE6m+c3CCXmPcMlBUzY+S//EH+M0zY1LC9XWYlklU/JhbzAGkhjWDzTn
xceSGQLMVhNweytScGGKizGDfFlpl/Tk6UsAstap4LlgK3684GHlRSiBO+Pb74ZLup/OYEkrGO3U
T8hqdwbeS8J6s7eJdkS3O3Wb4vrLOi0spwxo+PloJmbHNN4YOhqoRY1DBhqq6ETid7UVHOjYtAuL
/OZqDDRTPYkBSMvNGmUuP3ayGHMEavEmR8CEYK3Y7UhlyKHHHSNUbXIFyIsfhMaVUTJCqiAKv4gH
K+ZP3BOm8MeAAwX4SC4MQX2YBI+2l8/gFUblE7cIgu7GrOpTdSwlqeKaUg8Ogaspo3H5vucJSeeK
LzQ1vtMzy67igOKwM8yc++9gvmRZW4fOWBwKCsHwPmE3d1hpFuRqaoO1ZaTH9CHiVruMHgnLhdai
jdjnbPQMF3MaLKts89h8xGpygAcPeUGjShcyioYZurdJ7i8RMQUjqEVtOJ4gvsyY/wYTghImK1nI
FNf/GS8gtr6u2CewmqLm1Icjp7bpd1W7W0uDp1sm8ebGQ7vMkKHx0nuFZsnV9zviRupuO+O4Zj9I
LsdNyoKFRSex+zbbM/CAO6HAHyJPfcatexVpEgmngNqMmEJHnspE/jzXAqfJ/MsB3iGHgOxR8Y47
ZIYcODHRW5pB7rpoAKk0uolwzYeyZIMgthHDNiOwWuepMNeko+FeJ9BI3pk0reKrdEhfNFs/SRQ7
yw55feQ8FDRFQW5EirLE8nWtXaNK/qdDcjWz4w5meLPhiL+IsXAvdnK8jMXXwIlY792fxmebuJuP
oz6AxR3ZF1wpN2FFX2hxy1VJJ8ycUpYfCiZLKtBXHNyFyOQ0HzKxme+nWk3p49HGvfWiAAXV8Iy4
FdF0qXnCAOS7t8J3hPzNAX7QeK78ktmmGr/IfnVfnobZZxVHlE1/pmRIzQCdbQBK1RL/tiVI2j5v
7YEppD6aOlkAscbGzkReP0Ot44XL3enjzaRwutWOsqDzxs1yWv5GUPx0AnnWViQYsUtXBuCOyElP
naY0Z9bc7gGVM1LbVvALfUO23uxI7j7DRKvSQLAlF1ooQr1Z8knk+DKUimzXrUQHVkE00N3wGqge
hNDxe+ibXC2YSeFXzJWIHJNro2eZ/rZNUV7YpGhFpaaCTC+Yca9xyoGa7HlGKfB69XkaBa/oNDFU
Oc5sTpvJsEloAQ8b+fAFWGM/h3oMYAnbmlRkRCBDhl9Jl4fMGTT5xsbC6WttORZ42UFowNCaHTiP
tz/WZBCfgGmqLf6nBol/ljpkmUpv8NpfhlySXhSAuHxFhi8jJOy+bNq9vVbh8mU2eQFv6CSkbRZu
75Hj0EuaQIiEqcJFgSa0wfgnSeR16M3JR+WR59q62ENhznV6wWmaLEcfcz11a80E/N+UsRXmiK5u
x3OGr+tmo1CYOGXbjsIJoum78kc3HzIAhbt05KxBDqiu63Lo+QvMcouiY0cNcdDZ2JauBqzBV+A+
tU4oqRWx5/fOo0l5Q6WhTSYh04T8uOyU/DLWrlSKrwjtnPWEVccgkKEwkpNZYjRUikIWgZxKwbaw
f9BM06WLGu//jb6ayV6oK2BoWPmptz+EQm6tvcwRwQiCEITi4SyPj3wMrlA4tR5BF3s4Bw0rLY6E
ETiIb5NeMMKaxqIYa5Om0Tv0L0BU8QDtJVMAHWk5JS287bkIy+TqjyqflEvvk2HlvgHtwK9u3G3C
Lwt6tZf1fCaaJbl4XSW5Y5mPJgHhUNh0KzWSKTQ42gZ+XeNCBorAd3diD/DSzQT7KS3VGLZd2y0b
n3Z2tC0vr8Whw692ZCNSQZT3Gf0JHyLnkCvJNYLWVC61QU8ka5HJL0wd3PckHYr94mfDj9QmCKfw
JLc0YMRwseZKsHiWuAFB5cL5sgoiauo+GFOXFYrB+uTo4uo/xDcIO98TWt8i/PgLJGsPP+PVk1q4
S38S1VxbsRapTxfYgmdgfAtG2b8sup7SDZRYUPitEKstOI2DIGQZfcyIWz1aXBjGverzectXtgLk
hkE2AybBJRFbJSaDW1kYoUd7r6W3WL26gDCkU6qMykQAf/oTAYwcfN+/UmdqvtJwkrdLWf3TC/vS
RU9cgbdHqTFj5X431hePKllX/ecgomifHVIfjVOqOmfRrnhSwlpxByipBgIvt8gf8gh/ic2oAonm
HFBXQEQ7U3D5iJRhJPHgJjKneXoA3MAqEc2RlQ1Wy0QdQu6H3TXZokDSAdawR2638fy5w6tNhQq2
u3w7BuSSHrRZfTdtPz0xEMr0HwoaDOHD1H4YC13XDlOEGFa4kkhesSZAnwLFx9g5WWiTtJRJUIaS
Bg+lg/HZpSzafokDuErkKDfgJ3IJgzitrNGl9tjcHYWZGQyKBMHjCMZmQLh+R+wxOTBfzTjtfnVC
hc3FDup+FA82WknbvKL6NAFy2vHf63uCI2xYrPxCP8gHddfuyqRrWa80vpc31gvGnhML79TfyhvA
0TwoeDJdaJ3TrBw5Fd1cGyfADwwtvbWbvMuA4WGKbgWUoT3nAMHaWim7SnUbfYTWcIA+vxgqW/2L
dtnLLDiIbxAACGk75soxJx1igXXit9i5Z831PIEerpKm6gb4dvK8cOjqpW7IExxNtlwcHVhBRfV1
Lip1xGBo6aPZfZZsIVC5XZbznlaI73T5JBFQDg1drB2tLfMI1uH3UkjclXhwkm95WmaT3GsrZFqB
AdWk8IkemgqiPsl8mr+O9hkm0qrRATpHjzw0JNcqJAERgYG2dzqofkz+I4zPaCfbgrXSF2H7lC0K
ykHEbc/BlTaZ+EztfXUAMvpxPTt5Am6j8iF5u4P9E/0rg5UO6bj3Kbb0bWXxVvcxcFdePvUSxFbD
k3lisczdK6Ha4A5ODZMG4ioJcu/t1WQyCkGJZ6ku8UFNNwc+qJ28kZMM2p5G4gBkyP1HzFDfuQtR
0H+Lb6Hmv51E94UbD4qlcQHSlDhfBd9+5w7o+tytnT2R7GijF263+MpKr7+lsHsOcksSZ6woy6vE
yB8djuZC6bVpEEeorQ1r8PPRwiQod+oBJFsane/2bvetdnKVIpPS0B39jayLusWXd+twSB9ez0qW
x3Pu7ogLoFfTzHaqgGk0Mxbq/7FAZQVkE7FDoAe4ShHIQUtOiuQtWz0CjGIEqiUTjq7RZk/R4QeQ
ZkLaRZAPHV9WNu7vp8TdUwFWc2TbAAvvmDcQWinvwj/L052ryAjVI3fxC/pFBa4ngiYlcYJndSlT
6jGmnOBHY6zRzSTs6IE4psRyk5ipqq/Q6MincAs+arFxuKXXpu+iqbXPi5bQzdbmowuYstSBDmc1
dD4FHQTD3v/2K0tCLkR6TO3+AC3xYQUFY+rJtcVUn/IU9tmesJ63IuDDxafTmBGkUM8oSxAtNcjG
ZQhlUhsRAlw6BDHJaTz2u3jraaAnoi6ZxzJPM2zQ0L3t7B7gBYXwr4hgKwsq6+s7fZ9g4JHZrI5L
6zn5cri2nMdpc+6ErpUuqcJ3W3ympD5qgDu2/uhqqodhkQ25sP7YuVE4RPxu/Y13O8J/Rof6UcaE
98RXW4rgrF6Hz06R3a64y54nacvE37Z+PuLT37Pkxty4FAI0DiIBYAu0OF9tZsS0eID5LhuPreBH
qjE4mG1bwIvMcHR5dezgnnaQkCOoifSLpxs670ovzIB+mCprL5gYhnJVrR20oXT5p5XWM/+4fFeU
mPkEEnJL6vslXEr75kJffPKvrkgfo0H2kN8+4NoKelRebU6E5cQ55EmLLs+vJ5WJce3NyeyhEfbE
TNt87PxzfJs9RDZEodt5/0ZmttJ+5xlkgTXHZ/PMOKSYhhCbZ2mfCrMAnEQSQEiNQDS4qp8Hs5xZ
BR5Xx21opu12oDYLHvYpSzqyHNvJ17xiVmd6DziMwJ4wN38g4j6XzJsxHyeKsuJMZ9FJDZYv78eN
xZF8vD1zfeFA1t6n+CLWvXxdusau5Tt3+pfwCEX6a8jnDSoUZDhFhtBy/UlrWseSnF9zcm6es4YB
kAlP/VcRrIuPgR4glwDXkB6g+WBaLMzN7I+8jpd4oZBbH7a0j/iadlkaEDbIJQNcUcSE8hHlX6At
9o6jQ5JTN1h38BNTR/I3Qi+kib2sCgO21OfRQHtU/psRJ81EiLOj9h+tg8vVcVcCE+Qrw2s7APcH
OrandyZBoccoMbuioDs6bAkp9/2ngKYdpOvpljvbKfGUYy3KQRtl6DtvvhulY84UnZP9RD+GnL4j
ZL2oZWYeBmu/H8fwqUXOGis4WbJnvKaTpboCiVfD7gyh/RwaXtZ9jz36NQadMXkBVTAT3xUJGBy0
vpQd1PP/AakDyBlfCUo1YcjTI3zYVu9nTt+unAMqjuUQXdrhm21Ep+KXVG3+Zxb65aplOoIZAS71
o3qBtDH/PbesrOWHIt1w/jjm9QGvaxD4xP6HquYzHahnMOvZrYFXGyUa7+QfThJQdUDTJREXcpNx
u6fKAntqYu4dyhpwDYtQdjyOaIMrM3Ou+vfl4V8uUM43uRsT29+bHUPeE7oWtAlzYoy+PeAB8+Y4
s2/hZ7Tj36HB91ETyyEUwARqpGGZOK9fxpyX2nhUnBaZL33mFucUvQTUb9H8ldcR7XPA6GijKGh0
4GdVCjn7ja6B6g9NGSjaBwhaJu3Iz92ru8imRqUWrfTCQCXLHVrjR55mztCYIfvF0beUiZPqlqsG
jQxj2Mb6P9c8M0wMG0R2EF/KzAXIxh17z2DLs8kJ8MXNMDxgcDrDUDdUGWG4VXwds7YNE2cn6f6B
ysxtSMCHrHzOVP/Vl5Z4V5EOhgk8ickExZPuBhO0iETLPgSs42HJ1son+QAchA8z52Ui63b/egi0
SU2Zo2RK233zPGE4tWrdjeynzYk615pEnfO5BEyV2rdil78UYx5Lzit93J+oF+nneG3zxqRB/Aof
dPXWKghqlzyV6AgDbo7LasbqDJnUe5tw28YNIDnMcMwBsyUWEYd+nXRyDbpRSVxgRr/q2AS4ri4A
kVpP8hJWYjocCyEAlg9B3I5FwzB76a+Wv+tfNA7/Q8Uox/NOiui1vbQSiGFNNwcHzjqEoqtu2TZN
6/DLrnlVfrw7OI/xeBGiLOU8NIY+79sQLPzS/br46OpCtIhj9WaiSeJXP2BxtXKUn2EXc4qFAoFN
QIceLTWMmbeS90PS0EOfYCvRg2fEDvVYzP1uM8YvwgiRxhJT8T3WLzWK833y+Otai1d80KHzIS9I
LSoF5X4qRCYRYNKo1rjb7BVGVBfoNNIBArSWxKB0GqRxwokB0sP9K4qD4GrbQh3IULCF+WYOk1uu
g4n/iRQwBKxKC89ogACSg1r7bQXbCpFRlJ+t77XH5MfseJ8yGI9Ks0ifA+jm16AJUp7a3P76Uzy6
M/Wwg+i9whIFcc96hH9w/s2YPdmPLl2lTRRHk5xuv82SM6i1DkGwg/8QqM1x/rsGWuLDmNrIiBD5
qb6hszjCMPpEMFBpw3Si7UoZgCDYlJeLLZgBbv0rZZ3VPUGDY0WLgTwkU+VwvTWD/gPIeXP2X5cO
O2oIZEsL9cq5c6do/nvt5OIsxvwda4G2A/4yLzA8c1yayDkLDWCxq64om2Kh/AQ5Bfz1cdnNj1Ar
mGUN/j+ph36FjmMcfb4i6K3otGFu5fCDZJdeCkjV7eMAxCjN2mpTYxay8E0k8cLV7rwSXrs+cccC
Gn+jmg2CMODDIanp1sK6irUs3zKTyZ+x7JUlsWUhqzXWR4W45foGGZE74mvcna9Z6HDN1le9rmw4
yppCFGcNiTE/7VE4hclnT3NeaTyCljtmG28s1LMy0xNIeZlLKNPJxSg9grA+q221Aj69vzKsgv1q
qrkxo8zKno/FXR3rFYFWB+b4oHegd1+5dT2jKrP57Pq44Ykr1jfRZBvU1AgwwBgNK2zP//BW6EAg
8Ph3/dc3pRVCUt4rP5zEYkjG1IlQJV8zcjNyt45O9LklUfBsw/cpLXJhTv+d+XIqUa+37xuU3/zm
aRk0JhaaU/Liqm0KOx49Vsz3V67BRksohciVTqyvX+ae3+Dd7RG+oezRKY1Xng6g1Ywn8zKl6TBA
RzYxQocejQ4qT+yY5ZcKM8QejndWpS1Ja95uOdPY2cMSvELiXQFeElts2/1ayP+cSPQ+NGP26sww
FRt8CD6wuMfT7GqNr5EBN6yWbe3QVjANHI2hwjMK/uPQsiyvK+JgsEfEndrjr/cIoVIGUqVhATqS
fwOTXxYC8lnxShZ2JzhzifB293geZrYkW++Q8KY4TxqBuGb0HDS0YL3UX4MJ49p4VIS4ytgGoNH/
0IjaIoINuT9D8E4aW2129UahRrb6w5K4eQ6raZP5XNjqbcZA363n4az/85sSmnwsUIsCyLQv9dAo
I9fuUDf22qBDwF/u0ONmlCsljeBz9gQA2EA8M6QegkEn4rPh6368LXPbUmp9pZ+zFisTjJ5uciUY
BFqTw7cF6/Kj9YA7eaisEn1JAMXbjt5arRn9tCaeLKcg5777e9Ejc8efkyQNWMkbriVjYQ+0ojHu
ZITH0e50Tncklf53p23AM2sf6mqOPMMgnEMOMkzXtBykDHcU5jLYxjh4KM4RmHhFXy2W0ZznzlZv
MYGe7UVeLCjfYAinjmtdtzKx0VwCtnzSdwM7FhgfRftD+XyNV+N15zFOpnFcMRU5K4LxG5QFwiB3
TkeKutSkRTL5kN/8vP+NAfC2VsStP7Clyp+TA+kse1tg+44EFz8XZkaDDsUzNgmTnfxqD25Yxwjv
7b0/5+tO0cTMBr/tm441zv6ar+Dtp1mbghByHDyE5XHqgyxF+XHI6Kz8a4QJOPTZ0ps1pSxvVBK9
dueh2l0bVN48IltEpKkvs/QFsC1vIktEkwNcu2tx5kdjqVDeXKjthxFPNHwi4aGkq2Xx/KxJobw8
7PLa7xcc9q/gP5aIuVAT60y1uqrrNjspHWYXpdOq/XHKn8rU493zeX+ElUjxIR1h9/8Z0/eD3zuL
qUaF3xeQVRAGbJZtqvzcwA4t10mKhMx2wuDifhK/v68Upk+XSuBpR7NLmOF8sXZcvdMbcbFjinjH
SmqvA4WN27uDgxVsiDDH4xHnEImWallYn1ZHN8oBnxGrNWq89v5/bS8mC6kP0RrlDor6W/NU/1Tf
Y0Xb/kzjNH+1gE4nClO8vxaBk/4Wui4b5zc+gIeBH7Vl9sUq8Mp2Q34xxCoAFzrJlsf2DLoqfFbV
nOprUNvy3gd8T50RpGdpomHoOvLkmMxsh0E9jxjE5Uphkikok7ceirHEsrEAOYcdtuMXKBPdUZz7
7PrYfdjFHSfT2PdH8Qlb5nSap5xPK3/fvLS8KeFsSwbdorI3xAj3hssqliAHR2wFAv7JYUNQqdIq
0yumr/7oCGSCy0ot8ZKiZhPFomVLPM7SRCYXIVQfI1RPnPlnp/+0QlCEzuFTUMmB4DW1ahrMX6K5
7jzOyzFMG51Ju/gIfFwuEDCbfGktBZJBFsls2T5g1W2YeuHW5EyMHvwpaAW5zrUNqT1QZiJ6fKh8
nwF43+y6FalfnAHZNtl/Tqi0ygaUwFQS39JuKYrQqDqEDFTzW83G/sxdRRSE7Jso/l6T4MGGghTs
8vhN7sTq67/wP0harJN6WL33k4TOwr2SU9sR3F02ZukkV+NIS+3OLzFK35iPmida012Fy43eO2sy
qgvKHQdqLYCpMGTYObaBedSsyabTQWUXwcj1mKMfcYDo+LET18p/f4Yx5XczjlL6defBgHoopg85
7U3W5qP+9YWOi61IthjbPwMhjE0pUxvzT23Pbfxy3m0dVYAPV+ztr48d3LSjnZ/lkV3dTmD33U4M
1QgOzqId1c1lF11ZEHiJR5wW7rDNJ51Jejr0R7osfS16G4fE9kA3ut55Ba1xBYN/4KBicQ0EzVvy
17RUreWNVM4wkKYCJ9ZOY599KiFJDztJ6LZZ4rTkA8ddRVIrvgnSbsVaQmyo+HeVH4zHnsijsrf3
cp9ScGHwNMRXGK4Ilw9rY3vxKjqiWLIM3Z+IbBYFIteqZ61uy1UGvCsyVoBqgsb1+2Xu0W4BgGNX
CV8CFWi0PKRxLLjSVf5KImM7T2PJTmrf+bXXLQheDZnnHx158Qn/LG3UgKuPId7Ma4OzHz3qDeEC
Oa8KiiFQwl8SaX/ZffIAvzYHIXqGlFkNOLBnUUUcUicJoZY7vwE5X+4ML0E/LZ3yaKUXg9ik/h6C
PduMZcmkoxLYNtxpusnk1pJ1+hvoZfuk4aOgR802dVObJrvrPBeIJuVKDz1BvJPPZqx/GkQ1oQnP
S2f8tOjQTS7RbYVFl0Pqv2xjdPeySzs8RcmAX/S9JWgH124a0HwfqT11OkeOj8dF8xXu/l0PV+wy
sDJDI6PuOEl3hiAgjGS84ZwNXDLPZ6gPLGqezYsPir7tVPolxm1KozmIu1yY/3j2+NXgQFEzMe+N
5VyBw0szEH3vLeGW/EgfXckOlp9Z5O8hNwsBLagd4+cb50481gOMADM+SX/Jwu06mQMdRrYai/88
Jr6sq9tQh+UhBxalRPXjcWOcqa6K0ocZJLPtzLwSUvjCnSYPcaFd0gtqdLu67GX7EGTt8gQnWepu
MIzzohN7+N+ya7ntmf7JcdDXuou7AGfkm0N32/U4j0t0KrSUgNCx4VOGpqwls/cyXJ5lydj3e0RW
/EXLGOsADBpWftc1zTBpx7m61DgmCSyULahFgmiq39mmfDPxUbI4cQjd8emw74ajbVIxqMolGP8J
OARmKvLnDSaurxPP63oX87HSpj27S1jHzTi84f6RoxtwgXj5eTfEyzb6OOu9cm17pz0PzQk9NiHC
Z50DZmslI4hhcCKTOtLvABKmTQiCAMegrTWFyRy6vzSQRyCIZNcDP3LOSWJDPYhyJa2rZWexuUmG
aHd0fma8ArujryqCP6GF5RuMsq+z5f9TAj80rym19QPaQL/zDvkoHJggC/Ml/3m01O6g0IR1SJTU
kaLS47aExg+dbU5kZQ6uCM4WuywedObVm/jhwdHX7mTnQdL+/Lfff7gJ9bZUChaarjQJN9pD35uo
h7GZ4+gNwQ6CO3AAFgmdEhDQX7o3/1+4NX3cBdWG6gVCbWT209mc7VKdp0Ra1DLb6Q2u1KrlkF40
qtQxs/X7SPpc2YX4aDP2kCHbWC6o6V6gp0Jse3yqq/yyGuAXLbb6dpSafSeTzCEcUNRJMskx80yM
znDnSrzlB7oSvrrdsOy0AWc4WW7UhO6+ROegLTrNd9TQtXBTS/1q0M+IbGdVdnDlw8AMmLL8gGI4
vFDCHadGN2pCxB8fjNJidaDzjEX6dw6Sr9K95uFKsG2k9XXfSrEoSvv3FLVar3QvAn1Aiz2nuwd7
HA/GOdZk2497JZzhMZhpx84WVcHfP/p7zchYO8Kp2SEf93pe48Jzl4t51oFQLHSfFdABipxaarcr
1U7WPJj5Ap2kc5C9HE0d9kmjeap5TPjlUNd+swGKXJrBrY7NtWnao7OLcNjBiaTmNdaznR7G+dA8
Ellb3glaWWX8astJ0p83aisdzwqiMfxXrjeIVmCOQSpYn5U4nWarMIFtyip5ZkPSAsdZlXAEwYju
ktZR/b1fhLQqn+38SIG5ZrVKasvutsdHAXaRBIC0Sf52ODJ6yZ5y9ypUgLJPXoV7MmlWLiBdpwd/
/HgISSHK96egvv2pdfl1s1fP2sRbPzLWZ14vC2eW5pV3hpgZkuLe8hsnL/AHDBngXIFGv6l7Xo8C
/9mOyFCerGok6BxK3HCWEEWeODPgJ+o30bqb9vwaAhfCdpJkxWYAosdG2MbiY+VqtCXmHy/+SPrj
FlcRXI4gOEPIFFExG+JZc2gvYhNX1cGydvaNDUvAwzOunOlqLaflGehi1+5rSi/Qaby5D0VhxnPN
DgJSe+iSFJhBQzCsEYTTRjhdFKJM7DnkXwsX0U73vi1ZeMMZ6/57tbnv14Fzz76qvFzKH/3uKHM5
V63gnDLOxM2ujoYorrtDbFy/IUt5rJFO03cfF44nuBQTSITuFPk3vMsYXijMOdMm98nQzr+SjAM2
0MMua753r4aocq5XPmNSJMxWIhhD6L3O0wnlQrYMRi3Z1fOydNvK5wvfFYfgR4VOwtesqmmXtvH/
fZcz3vmiHbkw/iWq0xuOqnLpAK4rv9VXgWxnRieZZXEvGzen06nBpMFYUu2DZKauUTR0GfTckn99
P8Pd9OCqEOujI0LLHE3t/RXovnJnWdgYh9j722he2E6utgkKhPLyfgpSfwAwuwuv1j6SVj7BD8k3
ig7elAqVSzfJI2It/qplbdq3v9s07t0TG9NI5+vTZu8KbcqKG60sULJM7yJ/8/q8Rm0k7LYnjjMX
Jrh6scTZE9YRJJThPvnGfrmDOITXirOY92jbnoSfunm/6B1DiZqY4MSnRg6EVDb7M0wAKBAxtdQo
O5lfyAkQKTMLwRxIfrzVfu6nPOHRGY6EAJTCQ08D4ZJXnvjUzJC1oGSQkV8o9wd6EDZ8Zf7y97Ya
+EfmIC8rJ8GFiG5icd0+d08OO+s0AqCrFJElqTEmfBXfOkKBjUNuYEylZvE2TvqAmPaFqqDkrVvn
AEJTGkkqO5sM/Z9IozhnX5fd5R4bjHWvR2Cbf5eB5zIKCHPkK66y/MJasjwZz5snS36hR7Rvg00G
1T3cu/Yhw2Fgu87Ffw6C3HLe5M0sTEx2ypkxsHgzJHV595MrA229wcZYPmDYHqBrLFImHStYk8IT
nb8dee2JazUVQhlvhQXnzrr2fdfdYMDUTNaJQomMj3FV2N5UvVbA6jawd+ncGqKATMXd+v2N5gN5
VRtZHOE+weXNiL4GOle3vWhqoX1MdHYp9nR1uo3ZAUJ/z5DZ7dYrZxc3f5cmnpq+CGJWI71GPjrA
FSQxmrq8SHQrovd+rTlqXwaPjpPEwjG/doZrwNAj90F0QFktneEItv+9EmNbDIuT/FRA6ofjUENG
YTCZ2GsoZ4AQBHr6i4RE+27NQoBOByFxYiosxZp98MHuOpGF5jPiMLPGJ/wkQcap2NEuTjrRuZMF
WwmhUQnhoN9/4aFuV3lnWYxIpEwqBNbuRcyYFDSjnBARugXDIVP1b0MEXgqyFh3ymlVsgZweAA/Z
xz0cbHh/AoqcbAYhj6+OZlN9vugsS1bJgwJxrcWeUBtCJ676zyw5OGDZcNxuIOP164s3tOlOk/G/
YxOJ+eGjzMlYSmyeouNNJxJOpIxNgoUfm6UaFDEYeMvixo1y6OVvvs+5EiMm/wHq35CkxMDdJIdc
0UsZI3BFPcx9OvU7//4EWMxg50WZL0mmbJnU13u8Rdsxg8KJzFhBU4KAU8A5ntDjorueoLCeiTfA
4LQeHJNMpV2j6oLU8cxUnNg59j+tajvjKxXI+RV1K4uxw3P5I/vslFY+qWnrfD8EKkKH2GHWfuNw
OSb3s6volwgByYQ+0euGvfh7JwSGwjhU2rBAzLXu/y5yTtOpYRGaH3guyWh+H4I9k3elO8+Nxh9D
j2Bou3c5CNlQJKBKJZOFsQswZQkBTZZ/Rw+1JclGIz9SiCMQf/Z8FAnXzke0+Af1O8F14Fj219+p
+i+XsqNH4uADRgXLmrc1WhllKF0jwTWnajMnFO1idas6vJZqfq1R4EVGxGyvNv0Jbe1YPH9y4HLV
YM1B9YPLrcysZumTSEbBUMZrUHZqi1rAFt+6LrvrmluzzdXtoePsMZjNx2qffIBEbOo5Hd7+iC3B
rzXKyd+Aa1WbV0c2+W3U+uhDe3MPFR8ScSD/8f1jzRwE1fl3wbCl/MN8YfuIwpDQ9z++A1d0wRtH
gc08B/HmAqQwqIRDr1Ch2eXdyFJ69nt4/asITnELqafDWx1v7K0P4wVoyQi9ywm9rud+Y08f/IxN
Qt/KAWv41V6NOo0Czy20roPXoL6Dz93xmOUfo7zK8FFst6m7vfZY+XZbI5EzWADrR31qQw2hE+IJ
1EiD9S0KuFXBcdv29lWcKkB/XqJLqwFgDmzcKS1EwR/IIq1v6Pj3C4KTlm3dPZvBEgzhCC9uZedA
yoy6TDBuFn45DUc0ouQy9BcJad7+f2JApfvXFve8c7csE8eEWCf+pGqXI8HwHYkCfK3jRiAu7cod
0J5do13G2SBg9yb8dSFFNb9DGIdkwcFBQjMev/qYjmqsDKcybAVnjQfXPek5IZvMbY2yp4pk25zG
kEqFK944VjWuFPgu49i9XWRAKGRoNNZZQkkh7R5Xu1epZMHrvmQ+xuX7BUTlUeybuFSIiI75SyqW
86lWjfacMCOtAyEqI5A9mG5CpnSF2WtmRzdArKggSD5TXDqpijGdC8bzeAYhyDXempUCKueqyB7l
sBHoUPZlMBQcmV1fxhkOfYiz8N09neCgG4NpC1elhGd4X50EPkEdu/t27SxdyZRaODIdLSvugzT4
s5RQEMMj4kWDRZh4gNe5mJD8hrVXOoSmEyJBexWAc9mPDnLD/PZmLE+EKNNY3ozOK8nXAIxscFlG
13NwvYHKYz3pjOvDe9SDdC+yLnPtqsde6hQlUs0tkOUBCpoDO6mvmPZ6DquBjrGLOlkv9xm6T9ax
cT1nl/0HMSCI6KLBiYm+mVJGVxp1CsNYAAyQoHTXx+/xFGvYZ+kw2P5kNTm/4dskW98u3BSEdW+d
sO8DGpvs7zywJSyBWonW5Cml2dFDsHRPeRxjocX4A3H2xinAQEswf0wttd5riu0CiyJZt1KAlLeW
5pBhmrU0mhC9UzecnUnzJKDWCVe7gv5qyEKGHixc4VzFOfVcLO4QJbp9AGiHybr58YyFI/HlKrH6
j5aOEanwJNRnwq1CrLp3XHv8uQ5N9SqXSE+6rjyM1ChWxKj9zPjmghdDYjteb8H9+VoEWY4s9/oA
t5E3krsMUdaWTs2sj1H3QOJDBS4QO7zqHjHzJE/JprD+Bbf/jtOUAVKZ6N9HqXa/jY8Vq+9e60BL
wP0+Cv5Zb2UFOeF8atTj+XjIldmxogQv/L40zMuNG+s1jM9vY26n2YhhxbkiHVDnJJ09FmjZ11jw
rDQAynsEuQGPpGdlvUbWfyFQCwRaklX8CL1bEK6wxZ+UqWzxtpzD1wxloEGiq8ORrdXFpIOjuugL
TsE3CUJF+E07ZEiYYmdiJJcK4+PCEplxf1khn90boNLU5925+bvHbnLmp6s7aPhqi6gyJnnsPnB/
mZQBjiCc8NG5WYpKsy8jf71iiZeqDY9752Vjpsx4L/idYPnspOqk7Zfzm3cV+Tl9CFLwgqnEssO/
7A/2nFfDQXaLik71st9fhGnEMs1DRtpVUX1/b2d9adk8bqrCdR2CxC7rpsyF5ZzGu8pR6eCGTh4h
CBwvxHAuxouutvlyUDNsTx1LZnnS9Si5Zeg9Vz1798w5NY0dKX0Y8rScEMPWYP6gWqiJglN/wwpv
Nc3i85f11Wj0WJVgr8dsJix9r4EpvQFwz6MqzwT8Eeon+w32tvJWzHaqCtd+8p+50i4x/f4Bi+yC
8nsvdV5DGv4HZlvob4lVaj/tAsEvPy4m5o8Zk0CXn44mUGOdAYQpBbCgtAxEiXE4CI2Fhc7JFIes
59YT6pGFr0geA/+k3eJ+ZgKaYFOWcV06nXBc34Ap5peCyoiq9lpOvxjTp+oqqQ3djXJkLfElxc/4
gnCpjez02pL/G6+VCFeCgGVXR4cxQmLVFXUgEazyN0JiYHjR7c5pPESlAk8aEG2dB1hEIg/vCFhi
8h1g//tsCdrBizXLSomtgkXVPfK7jrqimG0HU0MtbJELSlKEXyWKWt2sTecx/6RRMJbvRzGpWg2c
2afXmymKCFR04fPWmosu2SrKonfLMWZcEbeMgmcQc+AwZYm6sYb38wXf1Yax0XUGCwqUbu4lOjWj
3lAg7/fXhu9YWD+yBIB0KnifutzmacEavTpPmZGGjJU5msrFtPssifK5TJb56P+8HvO1VTdIziFK
K9J/HyL0Nak9W9BEnXNaSfO47fMhcFF8JuKdsEnRaXxLzyb9z0+5LfURZlOAoNLwR5QVxc+efOp3
r8SrDk1TWwbn80L7tKLOs0m4YrquspVdtOjccercBy/OpK2Kf87g9oR3/0WwClrmGTTUeSl4d8tx
wlMU+Gy4Er7ifTY3Q+ilx+rSGd8yPTU8s2UnZ84JaCi08Y4b2JaQFISO8PU+jsTR0uLK84j8cHbB
JHh9k8lX2t4yJUIw2xjtyg6/XdthGk0wHnQnIQDS0CUEmP8w9o/qp9MjHQ5UnoPjnfuQVnIr1GdL
QBRbsxFFRdgnni2DNXKwVV4goWZ0cgXndzHItX+G14CWA6Iw4SrpmxHQIkIdw8ml4zEAlLB6P6qg
sxoL4+5KM6YnXMJRHd9mBx/NvUoOLIggxQl7aKpRtmnjkcwoeJ4+aALBYHBz1ExIWzm7KD2uGKxr
RXMJuwqGrnSI9D5X8y1XRNt97TMp6n1BYCw+A0NQ/0sz3uSS1uGlkEtnixrAle3XgRDLOMKLu2Wc
s720WNlE4X8UdHsa53IIZbJsaT62v2+E38YKbfLWzDH8APdJii1+zRaW0cOyfrLMRDJtUD45NQVs
5eufBN0H4H/F3aCWAeEwEAc/G2D6J8ida5ztUTltrkK6V3tlWgM2xx5xhebkk66dXruvmlva9B9k
rU1mZJxe81l22Mnm0qlcyhcalQ7Rn2kZ9L40p2aG0KJoHoCU3iBXF/x6XW738X72HTH7JkT4SOmG
6TFfeo3ZoyDr65k1ezR+PzgFqHJpTqxYrebCcTBCYTykqNCQmKpIv2wQBONIekSN69yfGpXpo5PF
UWYfnYq6HN57Yi0jWxVfq2QRLNKUYpy+8US5HfXwEYZgpX+7CdumlIRNPztJPZKWRIiMFcI29gKP
/hxuII4KlbGDB8d9qn0FhxtLuIsnC1Q0BYV2ZWkFYXm4tiV+etUN/NG0/YKTDx0o81JflZv7XrvO
Xc6smYP647fFux8IfDM5HxjXAaU1+HCItWBC6koYdsyk861Vk8f4Ta44xqX+uRbWExOeMUCJ0fb6
uW9ThOk/6KLWR9x/5mHAnFJ/YvmxzIqU7CxfrIJ+F36kJCtzf3SCCUJIfsWKWImiz05E6y6xcMcc
NHIBtvRdLKc42dLFLFNS2IfB9k477W+gOkEzHGgkjYaNTOeukBfvrFLuM17NQwfMTS2ctOA02Z92
niXv0wiwxZy7rFHQOxBIM3lf8t+XPOTKmaxZ0SUE05Me9ZXdoTe7QvHxGutc31tTAAocBpx8p/rU
dxShkgFKLi25GkwI5wCv2Xq3b6i1xF52vucFTVucJSdvsWWvhPGD+P1sBr6Z2vVmJJT4RQ22h7X5
LxyziH8K7h7TWzM3FSyEveB/CEAI18TOlep1lxmP3lVq1WcD/TXRJo+PU1lNpuJWFELtPJ1JJHE7
vBipDV1up90YYaWRKkIoJvI3gLvqTMVt5oUzl6mvgOR963AxsTSl5gsWONmUAjGXurDLGkThwQbg
Nb6Rkbofpo2Rxz5SMA5oRGXSiUsraARWyewgv/AZm/ZV3IzYLJjw8ZrjoQHDV6/O9tvj8cOJrl3j
cKF4ej5PIZ2BSYeQhjj+VA25ti+s/C7Y4OGi6qEv1ZGEYK5kog11Oil4+VmLCDJvfzo7+xg+vgen
i3MA0bN+oToqK0DRb1S5Npgn7PBHjhehhZFR0+sLvk3qHnz2OkeNoeDNoysM4fUI2M5iXEy11Xqu
EhsTtd9sazG4O3PSTzaPvVAvsQ1dwPPernbpT4riGmeOAll+QmeYZB/kIPwQyGO4wINCk55hs2Dy
SaTrDd8AJpRczTgZJ6YN+B9GdJbHOq7vehC5pO75/ZXGlX2E/nFE8uE3L3YW7uCz2t3oHTgQ4CGe
v9/toxxwbcR1PX3lHHLFqel0iOd0Qq5naayXNw0f9U+XZze8CV3dv7x3PDYzdklfqbKV+jtugwpn
eYrEQLIhdDrJuKEP2yPupuN7fQmtqNSXuVfDr5P8ok9mRnBrhbHad4onIJRfC9kejzO+W2n2cf6l
Rl+v4KnCAbrFZKusxy5j8jf9bUlCFxgqps6CTukFRQGUUI24tKJMmm2bBKY/hhRjB87UQq6H1zG8
aeAtnMcs5+kobE68qef2wbHfRJ3oK5wloOaVb0l6qQo+BJBt2dkVI3rw0UyOa+7fv20Q4HPYI2Rp
t5vxkjKp1vSlepGlJS8wWnyHUsEFZIQKU2SsroFHRAdk6drpsEZcSJdT2zdLdYMNpKJatsOrphEO
/MopvDZ4z1MXmizv9UEYX5hellMTFu7vLB0WocXOGQVwsRGrFjrtY8U2MyRRsC4vQBnu9PEtAIVI
R4qEtlilqBwCF+MKcT3rasjXSahCz0fKchCCOM7RPkaq0+Bf+o1FtiR72HHqwmdvXW+Y9ZmgmBes
LKSek3KJdOPJc/JmzhSAdFxrYzoeddXkpf3Q86aooVermoPuGudlrC5cNQ5BligHx9ozUx3hbvdK
5Nkfi0AzbYVnFDAfjWOYhhGMUZtJU8GlcZMesEv8t1AWfblSMAwm4yjN76DGpktTuA+I5BPCw+Zw
xDE+w1V4XeoEjwcLnigJwHXwd7AcgZZtAZG/2Kf2YDs05X6cFXnxYhqzmJTwZDrziBvQeTCJ0LN6
OoRczI6fSswAAxCujqUWCp00Ke0ACM4q0Vl0LxxCBKiqHl77e4zsQFJjFz3LGVnHXW5JgnMmGK8H
97LrMqU983mQceSVYqYw4Z750sWoZfXiUtnSTrfug7wKalTkBMeI02orXz+FzZzAVnUFg0bHWkc/
n0uP8u7jFKo8IioCZYG4/9H652YWD1+I0vIGWcvKUC7jThDHd2S0rs7hSjCqW+S7/12iNb+l+cCh
YG+/qxH9Szso2sNP/g2gFcj3aXlHh1LUR2nbDBYISVJdMSb3CudWllybjwBNQLzszMS08n3iTtLz
SoF7KVui7TbyHZJahf3OwTohsk1FehhJval3612yrRUwLn1KECj7cdRchQXudUgVGT1ZysAhDXhl
o82xZFOsKkHYNbyVNavgEjEC1FZWCwH6BZRMTc7iKvang4e2HxmnK8XZ1bvwqybxqMEGG1E1ZFPv
UARq+XxZMmewJsdkGN7EDGJJsNohu7STVecsRLGRvK67gALINwm206MWQ/gt5BiUpH2Ff9bpClCH
Yd1Ls6amGVFLmcxiWPYXiqtLywHtsGvxCv3OFzQk5w7PxZpLRtchQ1flBxO3IIyHpcQNRzI+kXv6
yUtSK0qGJ99eAiEZE/xES8x2it+1EoWhsV8liCeCD5FrK19IefdQXYA4hP/NfzC6Uy4pSznM6Aer
frKn240W4f1s+lmiTr+EjTnMywwOL2eOAY5wIGWkax9gLqC/i+3r2I7/bqIrc8MtjNDo6PS7nP1/
AQzrURxzXmKtfmzxfLNgQ0pqihqRBOWUzusLOVwaBD66hYeAYi7i33jvC+TtcT+L2VlhEv8SkFUa
+VYO2UefuKnp2v48M5Sx+QY9Gwgx5oyetI7o3Kv8ekeBfh1T3Cx4cYL8aywi75pOpgkx8LvOmNkO
dpzFuANi/nfribIMjUmAetAAJa+9exCqrBPWHFsdsX1GU9sfVKSM4AVyjZiCVOL3tAlav6eD1Qvj
q95PK7/mSEOyxevHRAzXJKyVxNEqed51tIzOnse6UBG0GNQiuIApcwsO9Ym6lGLgQHuRh7jwc7O0
BQIB7+JlMK3c9Ud7osa26Aul0RI+2vhugm5XVnMFz4QxXmHwYCCFngjCO3aTvk3Q1uSonRBu/HUV
WCDCNNXJW2YIZyn2TVOLcemOnWoPO3hNR5ATxSWpmOweHKZO2IH5yKZ3AcpvYDOWPk6dNQkoV4o2
pakAUJb/rNI1PlHbeioiKA/zLyD+Ll1qJDr0K0U3QI9nUzSgmqYb42kG8Q7mfpb2U0JxPnmfJAI0
p4ixqSBJGUih+uMLKmZTLYoXpXTDIUAk1O9oVc7gxAECtb2X4IS6lso3qLqRlcLbKamwwHLf/eR6
OcUM4e7guq7CvArVBvYVdbSMhP8rSE8DkPWgcmf8OKRMlfYVNKVtFXarl9GqpBOnsNBXQJ5xQ5bU
s7yOTzfsrjvhxCwfb0Hb+LA/6yrrZxIhUsLowstxW3+EPMqiQsITJY1MLFTA+SYMhytCLAxHb0Yq
vdTp2j/HejMBrDrRbIxQBXR4y5wBgz7l2lc6u3YBkAZbrCQnv4s+mvi88w8k829whh1mL+pexLUK
M9ab9iXxUtcbuiNH7ERjEAIJTPOacXu8tnnd7iGdVsDBImrjHjgKLI7CBD3plTodHHBws6+hiIE9
N4OfgKqrVHi29p5edoAkPJuPfP+pLIN7taTO8od2ztpcLE/Pxf2shi/vXwAxBUl0KO2JFlq0wh+g
rqpNoHxADG0XoqXuaKKeMo09OxOKRMNKBg/HzzJVW2rs3CbS5s/iHiSF0QC2w/CkWBhSe4NiwHdt
nmc1HRW633iUntQczaQK2Zuga0tIt3YiRVvp7xFrJocif+0/x5pr+fcvHb/91c/w0rs2H3njVANv
E45mSXBpabmkhtNrT6e8VhagkWfAH/BD71CuoSksoOKrQRJVIbOTUJCKux8n87Dl2PSXhqL3PvNY
apFLuooaZgwc+cztw/qFuCFSCqcMPQnCzmZElCmJJP0SPpGeCq1ZoRosYFJGDK9leJueUSkRKmPC
1lbEfq6FGoT+5LFbD0aukkUw4cNhcegOm7cgIcLtNaRvpr1S0Gs8Fg52NoqQtRaLpypJ645ADm1G
OQb3bELZ9FHsCZ1TsprKTCV+Rth3hYsx33JnZdAKuh9kGGWyFAPbEsN/u/XqHgcqoVQOdHBUFCJr
X7FAMW9rU6OIZ6cWOK1KRF5+y51dX5kw3mrDAI65j1dMb6Txo0rQrQ7Hl6yB7fzjeKBeZ4D51BMc
Xxf537NrzlL6XIxz3iUmkZ/+MbZcvnX3gz9wcYhax1VG5807RqsTSSbGcxEL/og9TfLV1UxZ9MiV
bXEB6CsT8LqaQ3P886s0cMlEkhH2hmudreAC2yRFr6ZuuXQcRHIZ8hPmBkAzpXB347s/A3VhWNTX
uBDYYcXtj/ZqCKnav+b7vgbTSM4Tz2PuIjTwhig7shiPN868P/8Zqb6DigGleTixtEuHqTHg8zOI
4bUzGDkxE7Ra+AWjyKK3RgDsx2ejP7lPOGxFr/CmlS7iurx367/8SIpmu+rSY9dbX+IpmzMOtuVc
LSaFcsmtnTkcjX4ZCP1BEzDqMrkFi6qCYgpVz+5k+cwZWHmUtAWoidIoUQkszpaYYW8yCVYUeewH
6HClNay13gEtinF/YGmzFf91w/Wn2ddraeE5KXMvIPAXHydCnI2QsLUIf9XfZx16WfWem/oMMOwM
L6b3fjs8H3kGsUAlHg1BxcrQ4thxIGuuiU/azMpppTz0O4ADfjXkUKfA610g2xZ+aVYyJO42VtUJ
X/3K4S6gpppahM8vryKGIIp1bcjcsZXgnQM0HQTOCso1qQH5c5fke9BgOWM0w1sdwS/Yjfv2x01w
NSnpuPbJh314a0dDdN2ONDUyabBJbZC3fkk+0+gpxdV0rZWLMo1H1o6XsYiAxzNtG6taWkCqNo5K
0ZFKIJcTVp13bW9HzNlEeE9W3ikfL8iSMLE77a+LIuP9S4OO6T3G5II1L6i9qtCqyJOMtpApW+M5
a7bXITTXomDHbsY9N3rKzk8DAWBj/oMb3Nzs6Ctrm2yQ/B+OaQhPWyNb0dfW62ff/SkTrYrg9C3c
0j9L47ly5NmBFdvZC9XZrXfARb8hVHsSHmdZAzxwzv21b65prgKiBCQJyuiB5JT2Os4l8edLSY0g
MUEJGm+iaClJV/4eRq8PdUg3HSVlV8zhzMQdeUoX1Y9V69mzcZ2krVZimLdqgNYgaSqjmgJEmi78
TuawL4RpbKnRIfK8thbuPf+/h33UUcBjQ5tuW+qWSSOC0yJiaaYWUHvVieCFX7fpsZjfYjaNg77d
THKDET+rVn7JGjD8c0J6PnHWrt/qjsIq6M4asEJ7ULKU+eOS+512EEQyxwdzNIQ0OXZynitxJZBd
fWV2dTLakkIFhg4ANyucR/8VJQK080A8DR9qWwQ9GQcWwvYKpvzi8DjTX6csW1tLFZd4ztUJpP/p
vqxoBrPfY1CeFPCfmZpTLt3vZXSqCW5+cyqJJKdyrH4W1by15QRmqmHYXwuudYzuLF/SAmUPpIKG
qsXqjakpDO8Q1ZfLBDcAHnTIssmzfwSyJZBPJhZuiPViOzTCP8C6piwuAYgnJI8A766ljHLa7Nps
lzulXRSjrXH2P3SXXhX6/LeCP0QjCZH/YZ46K8LZUtdQPdpwvXZaTx/zPdVgruLdBRO2ul2F95pa
qBREaOI6PAnfdf/xF2O22SWmVBQDL8V/umLxPXhngkWBXHplh+ki1hOehvPq1ylIYOmDmyJiTqk3
rmiGuZrz3GfFQJsS7/gsvqBp+FgH/oEFHMfvWVJmBb9VyuDWAprpNLAn/ZVd5MaCamEy0ikJMSbi
4VM51OZlnWe6iGDR0x1d0LzopK6NV5Yu7GUGmEpcOKW12+OIJfEa8wpBJI9ABSxNvpHlDlK4oboC
nugZTP2dP4rMzgUvU1aMSZIMNoMgQeT8S0QUT8bZxr3Rd7EykW1LY06AyxeM6L17d8p8WoEy1oAk
fpW4VagUz6fauDZ5EM4x+lWmK117LJ/c+dW+hSEQ+hjOMqYNPolm9I+TbQrdX2CnVT5I3eJJLsD6
FUJ9gB9+lumbDe4VgZYf4X0f1fZewLH23CW8Zd5TXO79XQe0EmprnuK8zujJzRD89+l/d0+ngwBA
SgrrkfwEge88NK9QHGp/62zvgF3k+G/H2H/3aEGE+YMmulVxwIQyA1EiiNpzCwCiE5jGA4v7zH1Y
C/wfa+aE+b47KjNnYr+7hr2sTpfbCUefrB8dhKdLUCdZDlJyfkj3I5cDu+aqKvAZwjAlN13SgBNO
DfAs0H4TfpkXEkhRRNTWSbGXhmca45GExEBNGPP0Fye/sZdjtUzpgEBuCXxk1lN9R/QsoEfOvAGj
P14U+geeJySFzGgJI6Yo53tzu7z377Rn0NqcZExfls/9Bl24wTKBP/unmvDfqQFY9KsW6eiZ5lyG
rnRRhbh0wR61CXvoMSJ9GTs4+Gq+fd/C7bgeCt8l6FQq0P+m84uapNQYnaEYFB8+IHpwAo5wycTk
AiP+QPzTwhGgEi1+cymvLKMNtA3NScTPSaJ7SWGgHmG2oyPKu3di8g/QpyPxZCAGVMcv8+Be13kR
lIVJLum6MLFK16+rV+5A1yh7o5jMR4tAizOajjY/sHErfR2haBMfr9z5k8J13x9Em/3xPL8jxcIe
q0O2SI/Q5Be6KZnt8XK5kxS9Jq0gG0IozI0kf/ZuxUrUy84mOsLqx8y56x7aDQPqK2y+94VMM+np
VmHafBYR8KScpWCq0Qqz6JaYDzhC8fmEF4VKgjY1HVsHIrP94QhtKyXZFmL/BWq7GPSFwGJqfbDF
F/Tw9A0s50XLh10EG6Ao+EweNTBKkV71mtjn7oN297gCP+z93gSsfPpX5ftGgzhUOXSRcCg8BhrN
HUmY8lpXCmf0VeaHhvE2RwJJKWO4HcOWk+Z8lr519NijlNbzI0BGgJi54Y30XFpsJbAfzpXw2pjq
hODVP+uZY3IpCYPvy115cM79gnYH9w+ZX1xVE/K46FlCUXTQoF+8y3Ek3csG4NXtM8bbRw86n6D2
4CI1zXoAP6hyYZFpZEvUDN0+boayhCetul0gzFpfHNn9IKtGfRAl8szFXwBYP5xHReF0ImYXUbA5
lS2nvn30DxBBYzgXfxEg45B4xkViqjNjyGF6W6s6+gDVBidD6G3gWTL69uMgUnZzKss3yZEiSscU
vYeARQ0H/xf4qHsct78zZ3YaqowQcU7gOjiuxWZLL/Drh39cJZIyRxXzuJ9NHh2VDEYZRx+5F7DQ
l/mpH4KXe+nm5v6wGeNnMu0ACS/AGY362548kvPFlCxdqg/rWKtEuLK5pDKMxeik6LnYsQV1WaJg
7oHGub2nfmgsfqnWtdmFyRBU4fwuKT4sMJiHdt/7S1o/MGc+I+LneXRc6alZyX5xfC6zGl4pZFGN
ehUvX3xsvc1y///wxcy2inUxjHXILzScF3Mza8lLEGRVAa3DfLlhtrWgBt9e+PlVvfv3C2PIfDuQ
3bkUyRFaB3KKeCpLaiwk+0xYfC88+7tBL07NfAMG9jMfd+ai9UvHeTJitVsfXlptXdZhszSkNiiz
MN40PYY4FysK53TiYJEykCCW3v4q8n1YQoxKAlwjFcdzJ7lut0EWufKaoZ4vB0so6GSS05rTfbzw
rakCRcRLdgTD9lKvHGofHpexspn463uV6GeJSgHWGE6sB8aPnQu6sgIj3Q1VZ1mkQZGU/PgIdF91
QxTAhWAmzSkfAbRQOY/JYmjN5mAgeM07e5ypV4WUopmrO8HbybUxEYhM9VSBDmC4Elg4zxAjFCJ4
QCHFHSbPBMdBRv5hxq4cOFk+YemcgAJDFKs3/79c1WrhPlRnoKW8LpKYVbkKuBXUU4IWhy1noi5O
BajHZ5dTdTHHqtzoOe6jGOM5uW/4VOIJTLYK/obqrvgPDwODml0+SD4UOKYGzaZ0Hq82QdZ2/1eq
Sz19+qi43qdRl2ZNbf2VZ6xJpxIZUoUdd0rQ/zPwTewnkLQjuSfDKbuB+CY93QVXW1/iiE4P59yu
CLy+jsK6gJ6EnTdnehccReP5yeLJRrmPlcjnHWC6TttGtU7ElJbXnIt8yg3wsiSVTZs57KPY8Kmz
RcU3nsG52kj6h2Xayvv0TwWVOvzmr06rfZw5sMg/eiYpmBh8Hguksj2SHmSDAuam8dL5Xjkq7YdH
siQ+U+NJVe6OPOQ88/flOjskI+tIStfajLaR26uiMld39joLjRxN44Wr1CrcWNFW0fRjQMipe7Dh
GoRmx+adNnBRmUr9YCM0g50D171G9BkS90Ad8cezj669AX8mFOFlNQmLkGPY+aRlmG6fawBezKEM
QxVwEhlFo9K+JC/Fb348jiUTmxDRPXA3QYeXZIRCxC/cNFnCYrBYKGRuJOC/QeSv1WMir4FVQldQ
pH4JahuMq/ypGKU7joh4+XLNtFNhvrBnmfOcvhz4Fz8hHzEM3ypeQIGAv7KxMHQHJ33s2DgPXCKZ
oHJoahbChq2cLZJHhZiVynbzCKYVzoyriEXH+SSr9/WmA2x/i5DKcmQ2EA7Uew+6MEOU3yxJF35T
8VCfsqxEclwQmW0SakLg368anribs9SvLiYB73ar/BWxGWtluQ1KtgFHpzu5k6wPqnygx9m/XFZU
0tjwnG2N/orxhv6FC5ICnoXRnv5vQ8STlfO5/+KSdB+tXqUz5elrzfKadnZddyLEc36a0b8YRwd+
FdpE4OlnNqBXVV3vK1D6NZ3p5lunwYEDuzpDeak6vnYOVA3+Fw/8BGjEu36iazEp/9MATPHC88Qj
uf1Tiy0cUvn1Je1EmGGdQUWdNGTKeDsPZfiuQaGojMTkL1ZImNiauNveYwkMt+1YUkqn0Aja5QnS
8KGqNLDil9i7KxA2v7uqIss4lRmBlUvoqCKqS/KxiqHcUOftmmFpI7TTel392jzH//qf3Jt/SOQb
0UU/zPrzPgI6y+43NoZmTolEWaAnJ+Jz4oJDfjvVWiu7mj2VF1aFk1bYWZW9r4nKRGf1O+bG6fC6
uRllYvnh4FD0Wp1SRLzjioFrO34OkGxMtIqXDIe//kMY7hSnhneejA4izf0ALPYQUSMheYZc5t4g
no71+ROsTGkJLT3Q9Ly2DuF4+2fsw1wKLfAB6scvMIXTp0IvDVWjMWKtmmmSJhRT7hJ89ugc4Uqt
njKmgH6YBCFSRu1ZCjbl2brlrrYrXL8aKCzhhyVL2ccbnCAJIT4u2tzA7PUvNaVacA5vlGu4HBk4
N47wIkmVJ6fZVlTCM1wGLUkF4Azzxicqw5EVbz+6QXrHoE4bIjbkIJFP9kyPWJtnqJuiT867ls7E
tdb9k3gty57PEEqibdM68fLj7buEJzY2eCBOnMRRrb7R18tXsnmk7wH6zHkiYcFLdNkD7VQ+YMbq
Hwk1ghGW6eeL2c3n80zEDUWXxQo0uR3F+uDwNuXcGJSOwV9r/vJ2h0KX/Ewg4SsR+AW+zvhNpAYM
iKdA1yXOQL1jgq5+oeIBXFMIxIv8xgd/yIkxYJPf6qIrHFX6MVq8cskIyFOUDRwdjubwIPf7FgtJ
e5VyH9UsN/nhRGVpf6YyMhbf1PB29wk7J/chvkGcRBwKQh4bcvNkWKdHTwC6APC6q7Jn4L8aj7/E
hoIhh2T+Pss8VE0+Jwt3r3CcApdArA3SheXdOPoMOu2lOc96L1ZkpeHEA8/OfwS1o1yNzGHavMF4
JmuGa4P0GdrqEOHEIzNzjmSbj8dMJ53g8ixBdWLuLSeLVKIakkW0a5OrZ3gBmoYKjEEbJ8rHKltG
0Yg66qwmZFS4hhQoL+d70EwaeYzgdBITEakb3GeVwQ8Q03mpAvCedLU5Tm0Br8tmhMjLsTVtGnKf
vsLBGl/z4v9QYOpJCr7dEA3f2KVGBBn5UJNzIYMqsgQkUgs/2+Ogl4/7vPssKOY9Mhse+owKIxTV
K7c4w61cVJGQAF5+R0hnMdUO/bV362RjVdiuUf3c2CPrC96jVbgGj8u1Lj7d3pFMEvA/S/I2TBrp
GG9JA4Wu6BbFjkRb/FHo5ZhgMtunh/kTICUwwB2LJ2ANzNUkMyuQVw/tmOLdpv5AvODsW9Wg5oe/
SBFRxlzTixKNLTpwPEozl+c0QJ185ZxCFfu85j8IpmUrTMO63o6rSmaj25fOWM8apWeEOEWyIItm
1z3Hs1jEtPoJ4saLZWjRKY/XMK9g5cB0zHWhjxJgqRsHwIxADjdKD2LXN7qRojEuZOYEohhX0I1T
2JP3VSg5tacVe7sXfrbvB+EBSeAj/+xL7pxk9ZL6RSOdV6KjuPACU+k2mYtL82UaHsHUkmQnRF+0
CupthXTm82E7nVjMtqI4wyXXfqcw9WrxnZY/GvdGtiQFMwgj5RlNnUGf5c527WmLy8ViHnQepgov
kV3V534xPnhjgIEfm6N97m93oeUmvNnZLJNQuOo4yGJIo8iC882V2CGqtEKCZmKYDx6ymjDfnuoL
X9oZSJiztHVfheQDtw2jZ5kniGgOwEQYFFO7ZuHKnW0atZLtdd/4Ck228HM+8gUE+8GiQZeOSGqn
xQn8OhLuh4ExywqRnTPCZvzpOqNiNQ0GSSdvuSJs+1Ly5X97QaM2Pf6aG2A/q6BZaZ44jyh4W+ms
Cw2DXFglbj+7oqA9kE5URiJPSnKn/zO777e0Sgaz/b8vPuPfGOYEqT0ocBCQptGkOl8XYL6/Ib6T
bnSgSaXkjgTSaUTTvnEuaTSOorXqvmccArcc0gElgbPEykGjiLPD7wDdL7v2uMfWKW3Vlfv8hgLW
VZJ8vnwKP0cw8fVIizbilcv//nDD9dAOU7x0cEA/NLBmoktLrkEpinOX/2J0CWYOy3rEhPZoKV3f
EvD7I+/VCMeTLRAWRRKc9767rloGj1OsyMV9BbXB1ZNcdag4cLBkrefPiTgNEEGyTtp/QWUoJzWa
jrLfpZnkF9eC3uBe3a8vxg0lHZeM3leURyf67H9zWSLiTXXbnqV45nLQBy+M9LMyKKIQNH7gVbpW
OtHB46cZw8boSZdOFjfv37/WS7EdvGJvrghiCucLM/wbrEsDyMJOLiVwf5yZ+rb2yMfEezJLb3P6
9gg0RQBcP7gaiMNBzMO/2SCEzR/uCRHK4Hom8W0ASYeKMMx1fhBH/AdgLKgtTMcZv1bVp1k6vzo5
WTXexTYCdRUpo/CeqtpIzso7pPAKzGEhGRqaUkMp40aBvcXYvf3xSc8iqRrfHDLCdMdwJl0nL8d/
ZFwVazkcxETDYRUmRG2E9u3jDYLQVi65VNBajbPivKjy1eqURLU0wwD0rLNIY9Bycd1Q81pSjq9j
QIxApQZtfNBXFSYZoztayOd70nbUajgvc/R1weYCF4Sm3JZDI/D8HC/ECspevvQi+DbdKx533ucN
kS4M4nncnyaL3mWE53l2hI+pdnjAMzbclkeUD5OdceyeedgI1hmxONn7FIY0NB7M0xkj1aBKPsVe
zY01Ysot7r6PFz+gWRO2SOI/Y74eIHCpxuqz7UTE82xKbRfUK2h5LWIUaWH+NFe9xlbbb9VGw5En
vwMtnVnwqOP0JZ6xfbkiW3+F9m3F4XtrDHR6BVPw7gZTO39I+fuAicm6lZVLVX/ketHCMKeN9+AK
juMDM6yVtXhun38UFlETb+gfwkoVhtK2fxno+1EFEnETwPnLa4zl5vtZCVX9kqoWvG7H9+hJ8Dt8
yRD5H3fP+tqd7HHOYJf87n+9gSnkyHel+dxNGx+lrdtrPIIMlo850tT/ITTxGxcBAChG2iobWF7u
2EBeTBtBNHLLn7cWJLRLrVpYx14fL7H3I7bhqQd46SSlmUSBrzuZ4XkETfmdOL4iScdr+F7irsDi
N3COjaL4LzgLGFJ3UE6JwlvsAhJr3gwFa76nS9/6AIQc6kuoLwIcO2WPddnGDFdDOaL01GOsgbEt
OYF1rtZKqqasVXvibNWkDUZDvygoPEjB578fwzYhfcNObWG06bSexgnzHrQRCyzQ4GeFBch9lH+n
4aDZrdYIcT/YCLEcN8fuToVtzdH5O161Hdz51fbNjfZRKTG29wxypSUj3YdQkPjAiyImK9rrLZfg
1M4RsShnqeEOiltqaU+Yh9xGtrgouICZGgBjq9xB2JGqu2BR05CrSEPMvglgen3itlSSTiedryel
CsbJHDhK5+7H5X/SEnzUqj4z+Jz1lKTb1CqilI4kOSw9VmdsNydd8Uvb2cTX7bC/SfpQr8p9v8Za
n6inSeU0IqaItyeaT0nvmgeW4co8UhC/MzWqTX1ADOYO9pA4tMNh0UXFpypb4p5kwv5t2FLxlDaw
Th7bhCO6/etQQx/9sc7ulNTqTXdltyh3UC31ZElIYbp+SpndGd+n6zvqYvEG3tUppjtL7Ox11qco
Sr8lGUHjLy+D1OSCSBJ32SxN/Imj/rluoXOEFI/dO9GAh8BRl2ZuWDY2g3WHHSp8eqtuWB7X8EP+
8X5FJO2wdbSwsYHAr4Fu3rXaEkbNu5NlOPt3kVRc3dsmpscI8kPc8IxxpgfXzfwmLYsJ51GDPaUa
BFIgMmmXgdLRocAIG6Gtr3lEPYg4lrIDQhhq4D5OyEAWjRAXvac7qn9fdERnyjlvVPHnd0qgl/ph
o1tn7B/gTYuQP15G/iTcri0iEobpcDR+hWdzNJzD/Vwo9VAyv5c5FoLgPqQBI+bogPQutG0tx5Aa
0OLp0A30Lj3GIS0h+pnTOVq6F5t72fv8WUo57tJfV4ZJbzoLeI/Y7mk0QpQDwCyzBdzsJ/warHU9
YJ3NZn1JFwMC7RgKE879HvpPcUU+M0H5j4IgOCx29RZnfxlFnBmc973AOLQ8IWgJwfQiHWZ5ionG
+/t19rx4ZQf1WJqfyPU6IX+xu3LefqUxwNHEl7AbovhWvpdhHe4nrP2ubMXwUfzEPNnuwxJlTBzj
RR6+cve4r7iirl94q5g2ArJKdZTQQWQEx8RUqX+k8UgGIhoeA8K8EG1giKkUM3EnzKPwWdpz+4aw
cuSpJ4q+wFqoZ0EmbTgY+EOBdSpiKUIsR3P3r+CRjq6dJ7AzSozhRDi8FhxO1rFj0Dju7JEjRvXZ
ymePGEjwvp3DMxZZv8FCGrmIZ5BMJNbDXo08L9fcQNmT6nOO6kmjkC1Z/kwX2+fkOeT6orf6NeUv
IDVbnEwY1YsVl3Xuppleg7cboaQ2U3F3M8wZvHgbfDSXE6FqIUdwqIthtqPLStZsxGvMd67F5akp
tDRbGx8TOxh6EAFkaxcdGybaI+InR9t6JxaKg6tVYdCZDrIE79TrtXqLGBwf1a31c/10Y07KIMey
DfENZmvwB9au1T5Fu9/VzLqlh2gP2P8WGL1xDmrSPr3uoQgquyZm/wDcO5D2lBhue0m5z4DDlJKK
CcNMqkgr0GdaUQz0TxXiaTfrwhnYDCuIxg46Gmlp2fd+LkI7sixSF/WP4W7SIsT2vtOAsQWHx5kO
JG6M6Yjz93xU0G1riKdxrCXcKE8t3ARK1bFZlAu4x675qL4KWuBvHbI/QFJ0bsXsFzwqDjd2n//6
M+/KdiE7cfKzU++DRArn/Wc+CQMTVi01XD+qkB1B96eoHzvcRHznUnqf1Iz4NlRb2M/Ss6vzmGck
KnQw540mYGFEmL0sVBw5jiO49udNXCbch3MBBcHZn+c83eNL5Ot6kWa3TvhUSoVzM73QczRnxZKH
aSmXSf8PAcFXoKCFMY7asCr6wOyy/nyQH2haQ+ttDRYb+WNTJGpCqxz+f2yHnRLmJUiE+2t0Rypa
84smx4G9IRJ2/cX8wLU08YSAs7Q2idTfWwjCd3llIlScsYZRxTsWvaEWbM0GdBAzwvBAOkRdfQhe
9hqpeJBfH3SYtr6MX2oXuZCYnJALQD4NNtZQeHsUpjIoolFzLPeCG5q04meJMVsZNF55vp5lt8pu
lEg5HLa1zx+fXAmo5qu3L3jWb8+LqIRwqrq0IzrXrXcWu0uGkji/eOOy6/x5UMX+jV7JZfu8Npi/
TU/23GLWuVBCIXzGycPMEDyTVYupOt/rNLKUTuRDRFd2wgla1qe3qpOMdq9mBAeW8GOQNttcZkmT
R2LFG7NA6XBx3sx6GIxLomOeU47N6NEAJGjPFR75xXtBmYEbhtd5uAlcUgoSzEml6nhWiPA/CL6U
nI9PkluA7eyOEqDkiXXE+KY7ycZL4I/SzJfsRkR+6RjtoqbQ92zV05iXRuVSGrc6S1mcDP0XS+Im
5pc6c4niP705R18mPfo2uQboQS97ybFtYdl4m5QjbZG/MK5Av+MatmhpZ+vID9c4k1wbU/YTatxr
Y+r/sV2Q8l50UaRKmN8wHhe91YGqYRZCQAbqUqjMz9dYXlRw5/OcnFMhnWYPj/mibTZicWeHi0Yx
4OMQaQmEtpyA4e0Y+7uZMhahjuK8klSN5xfKPRHV2+jrhQ9BO/uPFF4BFKfNxA/QN4ItOCisL0Kp
5sXPxTzY9tQn1e5gPuRdBSYNvcgJmlhNhPuoa3GKC+T+usg+i0oA2iP2hy2tuHkIWPnd8raDoFu6
lkAimOeUwGpQ35lFUXRTSAqDxzhT2AmzZlLB9e5D4Gl2MaI+quxuZLiFyxCGwz167w3mWzpqr/p3
3LZCiwTLx/5ykfdDL2Lhj28LcRiguKWWPCxbvAh9tMsMse8f5U3/helpcSYficp42oVucBDIcaHQ
WEvESPoPdR5tvFKsWfCU8gLRq43Ughun2sGHndbyfuLKWIi0RhEU00SoNtYJ6t78R2hJTl2fwqDf
CQnZi4npyQ+vroVkaacXtM2sidIclINzQ+JLaek6dNFLcFTu+oegvKGTc4l2786j1c9SI+hf7E6N
25GGT7FxOU9t0ZsXk+AKt0gXcd8zGnuwSpsWzzFzGnTzUGJYbmaPQlZGHuYU+CIWyGFOOUlm+o0X
+KQiiiMh4fBpHONSYosg8QX1QCzrvqYODrR0XjVcoB28IdPRKPJiBhCxwD/dPQODjjU8tU9Qs9WK
ftVAYkfp94Xf8sqy53KKR5GcqMizvsDwu5QiCgN2f+/rg2nG1HScCo8CQrw6m6Ap3B/XtuHWbf6V
nKPVToNgo7Qv+1o46vvUe4n6Cf23SkjeNxrv1ZI9XPRjjJOpOxTPQ8P4R1wJRO+/dlv6Wn7MTbkh
6orgREKR+dAyc9fIC2kl088sfdEZao79RTVTySNqR6v03E9XvC8dXwy2644XD8Gsnix8wHUdmRfw
4w/br5C2vf7o9iu63bIAdBpSpbkZrPjDaoHt5er7jK4Z9IFf4NI1L1ox7uSV6+vZejTG9i3Jg6+b
/ZzOnXAPjGBTS9Roo01LfpJojP+GrAMRS/L5h9HemtBuZIFmsuHiHfhQVy47bI58qp4T2KIRe4/c
c3Td5GnxM6s5dy2wBwNCuIALmBCjcY+oFan9+dmdCyvM+JXfU2LGE8PWRDmGkHLf0Kw94VSTtFM1
hle9tUzL7TuaEBzEPtCG8SeGGHAcNV7BWrzAFfV25znvBot+Xo/3e6pu54nvkNz2liwTxd7E7WrQ
NQJwrurw7BE+ZwJuS5KRiocb0ax/p2gCWonwAg1V2lfZeMYEjDQaVBtJOBjGRmGKafk+aHx3ERh3
XA6s3CDPqpnLDPhx54L/WNJ1kjOOULWguOmnOQwuG2LTdpUvrymHnvqmzf7lnMfGlsj4kRpkMEV6
bFXRqqWe1QhBTi6PQUYbipfrt2vE1gSSJ8sIlAahQmodZOeRxQKYXpaeRqYXzMmluNTiVLZfBw6k
eGmFHkNmMLi9H6jYiEPq8RyjoFHC9HX5vPdYx7Nn/CJT1+fM+eMocP21AX0RDdS4ZfGzvd0wUqkL
+k077NaSMwWr2rAme2oqZUHZLT7wiykxTT92vRC3pfFeDi61eR5IEqt/3dDMPb5JLS+501y6o7nB
QLe7VTUDzTXnm+CIfhO+2WIjRV904px0LuxIPRx1g0rTVCKTROID0J8tqFlYpXXLlS/dwvfRiLcH
X2a1vPjQ8DcjBC69YLcbdUqpjZ+cfUq+Rpw4Q5aoM6xoZOcqb6NfkW/WZcDXyI+PZKkOfFo0g5zO
MSPsEA+0JC3CRTdV2NAo9huRDjDeZ4FZpvLOvIW1DalecqmyMfdg5R+7uzOLz5OHOgrBMlKcKyaI
TnHRd1+4uN7uEiflQrIPALup0d7fqYlM3jJnX8G6NkimD92/rAAGvhjCPeBSaL1lCsoYSeMH14Pg
NN4KPBqgjZEfN0i6m+SoCwbUPOUZuBG+51LsNPXwcOv+Stx6l/YHmV66XBAXWLt5HoBN8ol1duCD
+SEG/zLEbKYLw9UStMiXi9X7xplQQFJmDC/Nl/X0G+HT7NlfWBT5b/dMpHejW+bMj8t9C2Yls3Jq
NScbW38riFRI3dzYB/fGJGa0pwaCyDL+YJrWu+9+9T4gdekW8yQdWNRh5Oec34QW57IW+AhstwQY
aSKWBw2/HqtnezZaeJE4L4gWU7vMyjEQF94SKPOhqKNKwqCvllS2nMmrs5UARxDuCYolVJnVn67v
04VsqtxM49r1qNoWIqruqf+JEejnuhp8WM+vXa0vw+a1/ZtKGJDr+RPStaCyBeMWJ4EbXLbSflzI
Sw9FisHvrQcOi06eZ44E/t4c4igb+SlEcGLTadrrDIlx2EvEcKGy7BTv2r21rupaIb58L8qWCEZx
CKjDDF9Na5U2XhRy4eDJyGxYlhgiy3xBnG1x+rtykshOjGQ3/ZQIURW4aFmMfNgFOGmWze3AFCUt
CTgyxp6/bbNwp+OIEIJ3/zNeifkblQHjbqdF9T2PxjkADwCbPQZEZLLqqehOh49GOSjIDb1nRyl9
USiYpjYpjc7lLbZlvJDEf4dGTaI5FIcp3b/NPIbk4gXsxWk1xb6+gUj2eZAtbVK3kV3A+gx7eAN5
dcbKbwppRdmrBwnaZjPWE4BSvX9QibX6nKIjY/ZuCaoOt0toIgQvBPydV6TfHl9+yvkPH+misCc9
6UlmcpNn1/N9Z6yAVQ2IB0cGVstYGG9lDGUA7ti4kW5AHvVi8uUku1saMNCHVyDLid8dPmyfaL0h
0/HSuWE/buXv5tZVvlYjgkEJ10cYoiUX8uopEcP9+P/nPXUEZ0Zc6IJVc+g8zGogFlCKWqO2a+vy
zveXlJ5umB8is2pvSforlpzAx/htZgQNj2cCMfRt/Xmo+HdUSQU8JEjAwAuwvR+9vQh98FefbGzd
a59jG+ZerIdj5M6HUHonM1fSpzFJ9VNnh7V3OMurGp/geDD6NZ3qyYRySXIpeuUrhzHPqvFlRtK3
c4JJv1XG5fCOGnbxAINMq5EIkq694nZOYrdi8N/d4mQBIs68kJemXWtqc05FnTOOoe4qvdlwbvpo
AtGNXMarjWPUT3x4qebOolUSJh8B6F4PlOLx4kluj/MMzInt+xywARVzEQVv7Qhq8bGqCX8+WoS7
TgGeJGR/eC6j7m0sJ8C2/9A0u1SA5qErplv73jOeBKH9JXv/i2TCIBmXz9/j8n54aReja0JO/Rw0
qO9EXOf/Bjs1sTukejXa6ShF0TMQagXCa7C/n1zuxUl4mloWIpSivuRz1OD7DwaRxTUYYVkT460/
D0d//hBZrz/JU5+Jet8Jq+cXBAq6NQd9/bznzyIREodytX9jOAZluSANQ6ZpXkbMi9W3r5b+nnn8
hIdmO8oalCgJYon8CxHq+ccTgOpLxAw0gsrUljfM8Ez0Vb7/07nkXm4xSP1Rbmsn9ZySLGOnoj1B
CUnP8OAb3P6FWt4bh/gvrjK6ruYBVY6t5NaeR6BbKctrmBbCZk/K/ZhM99J3VDIr72eAZYZ4ICD4
7KwPifgIF4hsee17lh/FWu5W+7MkzefFdYQB4qAEJ2HCNPpqNYU+mFw1w4z6KPiSdpXZuBB91N7Y
QDqMFjEc4TdsqwQ7Ff6Jr/tDSjmqs/DV0NoPlNWwkZcBJ+qr7t7tRHYuF26Imz1P4u04pKacaTuF
5h0H6evhL2gKIk4BJ4k0BNhnpcZ5xjzwtdhpjM/gVKGmRSS0cGCeVKaf4npsQSZuJ/6vRwlm8zXU
BqH0zxt3sEO+spLHT+ngnTdBnqX29kmrivlvT5L7J+Gxp1syKIOWMgLCHgLiSEmWmNMtAh3QBWZ1
2Iy4M7NNo6yoU51rjZYGn413l46J/mzmBl8GUnAo1GEzmg9oAKzqa6zkPF01jYR/kYnrctPNz7/A
EK0kpVMVxm5QltvHRt/hSxCGVg98S4VRwQOKC3LcRJ8B22RSwwM79Ga/eXYJCvwhCgnMMzENfjpw
GcKAccNuRwvk0hydI1X+EFsc8tgOITFiHbPpBWrTD1s+MF4uwQbxpHiEvZ1nFalSidgC/FTugPZP
Wo1363GAd/FSTXpBzKLpvdvPLRlzHQqBRI/Srk9bd04FMInq8eWkruTA0mTeNCkRK4fLzGabC/NW
iWn1Yl7liirD/8+TtGNLiFTe6mSyvnEvojJz6JRlHnL/wwtw0uD73SQZlDMXDRoiznF0eSU2r4TK
3AjgDuNcIFpAt/z/4EcWYUwsCl8hmueXTJzCB4DtMa3N5W1dwcQpnNpsE/F1PDOJIP9bEbOVmEF3
wFXH7YuVTgQ1aV7xQnw7opyiHZYJVWYj4r/s3amZruK4ZphIgl/Iedj1eSOd1pK2feKok2aOEylt
iaD9v/p0/k0cRB/Zvq/12pRWftrfb5sR48NzLDaSARIKQ2w7l8CKjzaxwNPcsYv7yktCXPmNpUsZ
RIuLQTABWOE8g/9tprUGl8DehYmnmN+zDPyzzlBxIJUq08SungPUcgp3dbJONE5IHEKEvptXAi4M
QiCzF2ydUsL2KCyEXJjSv2kS0nyLGdbN2aS7GcJnOI129vB2kP4/Nv7Gk6TWZ/vA8lIQxchyLidU
SANeyjPQZUJliXGogAUC1WNxwnkiBW69SjbopZ1w0eWje3UAQB5seahVs4N9dXwaeAGA8LtiO2Vl
PF6LRopARjLWSVAlZaz3TzN5DZtvEEBIY+1lcqTPYNYQWXyoBre1b2xcEYq/XXT4XYVOAeevJRuc
9MoDuua+y+4LHJ85U9qPVEWQuqhwOR9d1fbu8AgKwy2eBGhWteRwYMuUIE1cZ6zMMa4JA17kB3b1
O0mRYoY0IeXp1yqgUS+Cq/whdhId9bpo4Vb5TZaE4cX4V/yYrWMyyf8IzPi8k16aD69FX2t7k8zJ
v+Yjo2jhpPRlV/XElrZnTPMpuTuQRK8kujZ1lh17loBFZOLLQt4p2ZWvBECkhgnJbBbi+MK4I/g3
9vOMMCNHJmub5JbbHQ+kodrkMER/c49HsXNUapoOjOsis+RjChG7iPPktUgf3ovS6/q4IH1cDiet
8p93ocB7vP+AsVdfg90bQM+Nd+jtuPsv/iYhaPAnef/eaDSEnX1kp56NZGhAA92PJzudfYHId7J4
bqBQidh6f9LOtxP1Q+vpKtelUflvWZjNTtEGZww8ux6g43Nl4Hb3hOZghY1cHs/mpqAmk9gdmzkb
aU65EL3HS+9l6kU/Xxi5rBAMiYYCicViD/4X5I2ZNhw2h370sK0P8RUA8H53T5Ky1vQgKW+90UKG
5OG2bM4/8xLEoP7Cn/GZPw+SLp6ESxJSfBgn+0a7ym62uihAReyxWNBGeS9HSNbn2H0af+fqfUOh
gQ4QI/o7/Gq7m89Kq/U62+vAn6StrSnSsI6YOJ9S1lBlUEbIXyO6Q1e49ivQYgNsDxYeGtu1hYDo
jwzQPdlnF6R+FdocODjsvltOr2T+VeWz9Fx36YWaunaIungyqyDMO5THWUweOYZ95IoXUixeSJBR
IkTDK6bN6vcnOCKsFi3yGzrsnL90GXBeliOQs0zFSMqL6RS9uqQLrLq5RO8FJomA14zExg7+HoCh
GnuX7K7itT4gSYfzsES+sjKf9U4rqUkY2Lv8dcrnJVmbmqmBTn0U6fDXj9mJIk5NtJy9XEc1K128
DQ5f/nVZ16iXdTNItvfjMUcHGNeEoHK9T2XaYuJELtSm2I/qBBeAiasIpFoiFPqkBysmrSStVAOn
WEeOpf9V1NmAV7EEuAsIU9LWPCgMKMjJ3Rjca/cNDgxqsKQ4bQP90aaPMZrN6xJanWqY6iab1vt3
qeULNX5TlliifhLHHATgT/ioxSOrj6tIKSjwJJMnPI7xg9vqYFIRguPw72WJqLMnwdPjNXXzQYPF
JOLUUgvgCohh2oYUX8joafmJ/1B5jyHP2OeJZNjosyEYzJcPSI4vuJdvESROnxD1EJOiVwcP/pYs
vGB0ghxOu/sn6d59835Ugg7asGFj+5Scz9T954kq57OMaKUCROFgDARZK9rUZJ3HJi4IhHJEYuXN
KLDPKVW/3+m4hPbmIOkJ4MBTgfomUg51CcLjZ8i4Iw6S7SHXZ4cCuUPmTNH30WxovnrxfkS/Hls4
GXFCA6VEnKZJ5U7/8dapByB0xpLCJBnL0nTBp9sRiIpWB436Or1m4/xL9H0tNQOldu2nn3tzys8H
QZT+z2o3USM57LCSx5uqbkydd91ny519LPIghIPXXKrleHioLYB9U242guTz6UguuxHYauN/6T8A
ndIgU2tnZUcQEgeO+bnH6qO/dbluG6pUfFYdkuX1hJMmMRXtT1mhSjEvkQhWJzx/VxTpL6qis3Or
vBkuG4Qk61v8KfU0x0ruRlmZ6u567ODBeaPcBnGhxnYQld9CQhdZQIEgk7aUh9rBeKgMHKh77LGq
gZn0qRiZcg7jMDv9x0bR11BtDZcl0E3cTcEcy33LBZIDpcwkvQM1JY0aubj3K/xkp/VDAnJ0DyLa
ZOGv6sT35ASAVx4GCRk2nZr6/LvHIMdpOsA05q7RSl2yYFtjuyyvMnY/hxJS+W6HrhG3lCcr+aWn
sKVvD7iQWacgKSIgAS7wD8/lwYvQpbPBsQGXoqvcuMR0dZVKMmmwDE/9fKwRUHLLzTfPNRR+G4su
/uNpGP/in/7jCEi6KprZAFTh/4IWl+QsKne/0lIGeRhCXkDqNFPmFx6/1JmdG7GWLFF66FfUHae/
YL3kg03QGtKJpOeVeLoUyMjcyz6asEZd3CBLPD06ctk/HIUrem6R4vLAMnoKh/aA5eIIXana47eI
LXIdFOkTR7hO/cZ2ncVOJFpZvg+TJKajSIyygEzZZkp2O1oBR81Jb0KfVM95rjWdQgdN8wBt2QGC
XMpYlweLGRg6xKE6jyWWDNCngVhUuwPIWHkYRupkjRDBikbaJWLuWIhvPkSaoxhFO7KJPyGkY1Hn
1DS0RfUYbe5yTbkWWawaW3V240WT6akVIW5CvXy3vy8fFr1yRjyWCIXJRjzrsILIk9LTVNknOUm1
Dvq3zGRbBYB8TM0hfL9W+dAIPxU75ZPbpUruJJfqNKoeAWzbiti4Sil2/MU0jnrr6p1ovprqTb08
iVJjM3ZSB5TEkI44eu35AlLouzKAiMKhqY6+JdN6MqxVjFB55SWVBCEtnMif9VlHTCijqPJuA7TD
vlGtt7e9DEzh2QEFJgMiwhRWn8Qic7NYzICJgmSYTlI+IQ31QmVH2y7vlFHwctUeFh2N0I9HH/NK
gjdgbfHm4QK4AjaYgNtRMuL9xWGsGYO0luF+dtY9Bo5QFgMwFkoFiV+6XJPE994wsZum2Jevc/bC
747z6ZFJALxnn43escHQiAd/qjRdId3e7N1yJ/nU8szlQnMbtakoxuf4LJwEYDqFeUgR9xCNCH4Q
dMb+J+BuJ0+Ekse1clDYb9NTZLGu1BViHoGYHg222X3JrCdkmW8HbYe2ueL3FM2+ly4Svxm7asnZ
0TkfV3fwJ8Sj34qGYBCbmI5643nJABLAs0NwFdvWdqM0GhfgQduInAIcCvaS2jVayEr+yGUApUlm
yhuSKZJNlSr4Y03deVkT2kq9iizYNl8EnJ9KcLQcnzMjhIfLOqxDLacwghw8EQo8yE5VXzMiZbmy
U00oY6S/dhGi7RPgqG2SLoGKbSjx5cTSOx8lgfxgWB5fMxl3D82dO6+v0xHGlHxEXxJIW3nvtY0g
NkAG0NGV6YYZxJjWZuTjkvP3fEFok6nPgkdG/MKkrh/+BLyLwRWlZ4oXxgI4wmXYTU57vR7nH9UK
ePMlux0PxHZqMosKFDY81NSXw/jWSEHWUo+t+ilFKLlqoy8syA/KFmWDI7Fs4C4SnCj/H8QuWvUK
b4stbvuCzmJkcVHqVqpTaWR5KhIH94SXG1ihG1Wr1XncTBlmYXOE0QNyY8WxMQ8piWZnNMyeqsNS
9oESAVJpLHRR6Fyeqi1IdQvZTnavRF+YrMWL5x6An3rSeyCW4BcxenSlocqeOmC0owoRZBxZw6G0
mUAdpWLM4/J8PCHhTds/UUyNk4IvYNyD8vbksnDncIJnO1r3w62gJw5WxQOrHEo9qbfNGRNd84vG
FqpLRLXsja5dvmY7i5RUBLm0HZeGpr7bg9FMb1iCWOJA5E8ruDpTlZhaD82pgzSo+3E9aVRsN3hJ
Qu7huZTcYLBh15ECJ66oBGv4Dh3XKCUHSPxFhJ3IN7nY2CAVuGpZPVLOzR/rEApIUe1pd7jdVLSL
BjetNcvW+lESoiUwnlcismMLJAUnunSNc9TCTk5GuHjz2OKgZJ+AzLPoMZUuvkkvkjsYQEbGrvbE
xnniV4UB30B+gDnwJUaPbdXJJhfzmMtOUvamf83nDghH1OaqodvugSFJ/HVZIHwd0XNNZWL8ykgk
eunkqwV/cnaeSs0YzXpiYjMEtlp84f1b6MblyyNeq+awryRPSuQQlEr6fMtITSzv6uaPJPQbElyV
+PBhuv/KoaSbL6SM76WYlcZklKZE+Er7CE1RNC2k71C1rBp7zVg7uYafljQ/lPzY7M55lSKG8KEg
OVcaxZkx2AmtFEv6D2QlFUFRJnSoprb3dKH4C75BqyTMiq2X8/GjM4xntB/0tgLXI0Yr0SoeMprJ
FYBNFGEylq0EWXZQkP4bUtv1OgVliNr6YqQ0WrJir7+TGyOTR8cZgwqMMVoMIvMUnbGpyTThil33
94wrI0Ts4lnIMUqrqRDa1um6bZ1aFS9P8mfSS0sAGpPmhZNrwwlGoKeKrgE/QP7C4Q4iAhdrtZbm
3BIB1MXFO8Qd2Sc7+uuJWZ/N3gc58Vx5BMID5hbg6XWCNnd3xzCorQFSv9SKOGg8svAGr1/pi+qS
HYG4u5CmpfMvrXUpquH45zPfXd0lmZflc2vkxAMiFHXcOIlX0gDK21L5nIfL+5wYjjVYwxNqgJb8
kq7U0InI0wAZm495YI9++YnmZq1mi5Sx39thdOwJLs5WVAdG2tY3J7f5n9ljf6U8fb+m7nkmWwMJ
3WG2Bp0Q7VA2SknJzwEtwlUcdrUF7LUAdWY2pZDTfiGIyoWy7CxHz5HUDkeEYCVhzO+KzlebhESO
an5kwwyaoPnRojAKcduwkM0CROuLBFbQeEkgMF7zaRJViS+v7AhbVOPiwl2e0/RWzNVJfUOftoJr
jO+7aCMfjHbPvHhmQq77j6hn+w27L2YUvE5cq98EofS2atPDB0My4P4xaV66OVwyT1Beud/jsJFo
Hxt2Zvc/ED+wbyIcS7rzHJ0x9tyU6zLtir3LjCb9wpSi7YuHlHIwfymoHSeNJvYBYaNlwrkOm1h/
8n3w3TwbNV8VmYyUDetjvkJLhovFOleBd6x3seLYGt13QweQrIcPkghzV8Y2YoU51JLZecdGn9py
/w4PK0IeAcNGlaROXgJlnPEMivYVWAvs5gzoQmRbMWfRssEpGIy4A6SoWwdJ3eYKShAgppAA2IMS
bNT322LWdtVPlIYrKuHqcKejb0GSeW5h/3ERWnojwdwJw5YVG3SMbfXSE2KNV/Xu2VZnK2x/wU/U
ni4+YPjNLy9MUcJe4ntR0tZMR0YZNWPoj4JUcTJeEzJfa1oMh5CC6TMXmRWTSUlOSC4BH0d0v1vW
H1uollsyZTRMGQ/lcmjzNDHqxoTNgkwy4iHwlWAo/6mnJWk1afNJx3jYbFXUK6txyh+Cu7KmL06U
Q3gC2rb/xOWtJtvFBjhp19Ia4zZQddrFwm4R8f00C0zWUXPVthiikIRynZ7waHCG5q7H9P0UCQ+6
0P9hyY15xm2mesXKIMVEMIEvXV5yM48ga2Xwoe/VgX3p45GlIM1fnGBqqv5JCuzw1dySltz88GOi
/rKEAQIUzRwvS6IGxVZjrcDFT1cVizVZH/umk++xOEjEy7P82VfznIFqJQ8F/0/oTvc+Bxeczcye
PVo1FZfzsulGGPPyAYbI5sTnMepxZf5g6M4fgKY8Kq4vfQASLysWsKsmAa1YDkYtmddNpf5y9kEo
UGwJGGQR0FjSDNrsuFSg4T9x2ML47O9UIIX3EFZI0pCO6xU0KdJHdD3ulz0EUablmjFkMLW2R+HD
Krh3xr7EdQVxLtKtunxwn38rVhasJ9ETxciwLvLd5mHjd4l58OrMjzIK6FrFVQyYWRjRKrGMcwoA
HgMJCmHpr83FitFE1/t2en4fmToq1QJyVE7OYh3VXqpLRwP7s+qVtAXLmMukLAnTSJ6LDA0A7HtL
trjJldeffjAE1Pt8ULcJKZJZszpbpnMcuJkTPvoWWhxNDhJIHXQTv6omGpYMUUgpjIamaLcoiNz/
K61CWY0/ad2Qx50qFgJ2wJpXGfF/p5S6tuANqAd3CjbR2mP+YRBZOHXnGDDQxXU6vLidVPw9lnet
pT0VeaBo2Yp4hGbs9E9Pw3Sz6SZnr9bD3w98CLoP2mejMpDBxyhphwUEn8qT+qqech5VcnOdM4sc
NNf+niwBDV8fMYrt9MJ+dipX3fc7Q60ld4RDFQaOlBVLCGv596lPKAqjLuOIm54UWsTL2qg78tzN
nFuNc9MuHF/G2TNqqTtUqWTIzjGgDNcllvog179l5HJ+nhZjZM7tpkghHxfMLG3gJu35Vpcn+dvB
PdFkyVQg2n2QXfE0jEK3oOopL/C3+PE0a0W2U2l58iYyWR4P103r1DS2tWcoAWvVKVa4Q7TVbS1W
8A1TjGLgyTArjrErbQekSneM4Xc59mbqQes/kFmIX6xeq4FDOfAN5W6Wfu9Ij5uy40URXnYPi9Zn
F2budo5y/K1l3XGvjJ96prhE6N1Ql/gvC2Kon9LCD8WypNXW8O44yLjbtS4ozzRyS5gJkQzbHcQ7
tY2GNCtXuhLQn+N3UYyr8a8DBNL1i9F35cYOusDkoug5h5a3+AYEBsFFJ80wSQU+m5tVcy3HbfBW
agnrAeevcBVMCQRRmw0Xy+YP93CVTE8wDx5pGUDp8tiKTejLdMQKGXqjh69pGFFwAPAbAHeTMGQj
BIfFwAOy7S7ciVjFw1nTbexLbP6JvFzm1viTNoyrGS6gFxLDNrom1KSGdPADmabcUrZf5FY88qBw
a/BsZLXNDh2+STxa09MCx+s5ULumlz19KJWnBwveMpPZHkHg3cHnatrPsMxMPXIszwtrQwrjyK5i
oz4PTz64ZEnEeMuUZGEaup0/Tte5JpqcNpFQmAucP4eOcMNN7gcPB8rLPcMv3UCj2Rhsln775KQn
KyCM+svJ+ZSV5yRtWI7M7zGue4F1lCgU4fcMM7lQ/I+8OCmWXxYGfWwsou6wEtBYgapFeiu/P9ZL
D9LWbQ+o1adoe7vs/SrJcNdXPR0KXMn2NLqX4cDudpGQ2voVkCc8oqEgNTGOKxtMpHmKvj9mIoKA
pjelXheVEYN2201PLrHv7rwy+yIkAvnn4IzYXlue5JpXlX45ZJg+afFUCihIA8/WTdcDN9WJgEPN
1Pc6ES/6J4XHgjmu2GqY4KoJiIuYe68YjjH77YxRttvjpo6cLQwNZyf5d6SlO9s1vP5mbFefeMmp
mdG2TZ0PBEiTtOEAnmXioub2xXPWdD6H/YqwAHr2axuxMTflyfyNFpDNV/LrWODRKpHTRDiwfKgJ
m4AuYS7n38QN/6Sz6CDkjJgVxG4R47PtmXkrnr6fJusNSxTWa94jzKC8xqhIM90oVVBhmRkm/Bt5
s1iFh46eXUnbP3XwKqvptOffUv/mF2xSjd3tXXejd2kMU4bf6jYQMDUeKs3dOJCggNxEmkvRuvl4
Ja5/cpxP/RdkrDHobVVTeNTJvVv2wx9LADMjI+af7UEk0UPmBxw34K5Zh11o/ZTHE2U7Rk/22goz
Iyi9PfFLmqyhovrVnUeHrBunsqk6U5pGW/GGoE5yj8GQEP5RElzidV8F16TqpCOLmx45r+l9gZiN
PY5zFYhNbJZ+MGb/g86WcGHQpSu7r7qSH9uILBKPVQ/jDEBaOB7yl1TGwj6uKZxAR4ZELfX2D55Y
Cw/68OP3cB5nTOKbZAlMkJGN2eEvwB7snpPfTihMl6uhTbRBjl9ixFgY3ocZNhbNhgj4D8TPLmZp
HESrUlBH7uOZM36fw5w26jvv9xjsoQbdsWlqXF5Nfi0Ke2e8TSagi+3+El3NqoaU+7S8inFtaOeb
J60/6iTj/PHVAPyca7TLvQYxQHQmagGYs6EUY843etB4jmTbeq0awXRSPZLIlHNmDdbrJorWLNNh
8VzWxBezdHpQSDx19jJM2epBwkHgWI82u9kzN5gdVY8bRr44d+f+zk8GbK+pBmsBoigPBhCbC2Ku
wNx2uDN7dVMB3ChmJj0qIVeTFQYSYF/aSasfxDo1DUzGtKhNocz46Kr18/aL/xAvhME1lnODP11o
LMLRf+AeUez2LAOP0sqxjp4QxjqBVLagY1GVzficV0zFCdTp9Z7KmZ+ncpYQxPR7EJ751vzCp4JW
mJgt1kP895T2c6o5VBmtpm1n0z+GBQisB7tkp29bfqVdNFsN6aL2liy2+SNpyScCZ8ArRWfk3AC4
sZkQLIzh4qTRPIdrlcwnF+PxrBxidFickexTp0/A0t/OhwY50CDDcuRRk9tjI4tqctaMzmXOXdfV
8RBhIpl8uy4KMMeparFEIRAqNYFcuhv3YU0S0gJqBhFEBr5/oYjNBOq2JcXTEaNTSiy/uKaggMn/
FxaZTm3Gtf7Hsq/aZNkOBfc1hJx9t5liBm5TT0AbK63nGi0X/+RO3k9qO0HE/5ZCqtwecUI5yXKn
0ITkgL33jXMQfGoeDsg6IfpoF2CvsnRLz29w9OiiKRlxkPLRGeTaGOrV4qNBobKSr6uBs90EOL6Q
OT6sDGVxhI0ELHEDRNyFLsz7M5zAqzynxg2IBs/60XnVfnd6GogYlHi+mk1udJynDI/fqjnsdFac
PLBx3DpPp3L8C4I4rmJ9i7WlpVgD12+4oUCiAHdKt5e8OP2M62f4JXXTYWpwUijgN6oj2hDjqIzg
suxmF/2D1Z76XfRgAB4kBVYajyI/Qn+bjs+oPlvix6ICkNX5jrcTnXi9W6VEadMPdNAI6JRkDv/2
h6+lW63D3/MUgMmpiUdYQcmkx2Bqo/BfaKEEpv+xTJ9zqs4rybO3FScGCAnWEh9Bq8/pKQFawrPL
8sJ+5TIvMDTN90lijFQ1snI6zGuknS/MarnTaPrcsqCm9p9EWvibpb0hrj5y9wgPP2eNBCLm0frX
VkdiJcdcJKag8XSpxzqmz1M13DNIjPi5NRWFJmnvkHM3HKT9WmY3s2Cyr5lkaIZIe2jMJafT7PGO
H3bH1ajWIu6oLdaWAnJHgS89xRaFT30ExOtHdpsaD2/FK5eAuL3VeNKmnnQpLKItvdNlj1cREKDC
snyH8A0FuaanShpiuLjHAfP/m4YgCUHxOZwVIBozOJqqIPWJ8wxHK1l+L1dRoMQKwILrk4oc5N3r
CFDND33r/1oWXUzDvZ8PmmJ5T71x3E5lxan4xkoFACFiopZSyG4Fy5prcIvb9nw0tb7qBjt2X9sA
WORF494x3zY8c1HelGU0GVZIOv4hKRkrejRH5pZw4ABLXTOCNIAMhK+YKaT1V1BA7brN4VxMMLmU
Xnnozcxrh7Db4XtPaDF3Xyv8rqAG72a2NG6cMRJG6lcWow/EvQzo8RDhWlvXtOKpALcFLOH+ztRl
GrlMd9eNanQrj85SKWrePHcaULClZzE95ujCNKY11sprtFgjz2OKLTf7kCznsaCoF2kOEIpVp7UH
9sVObaqLlMZpQ2uJHvVceZ4NEubkaWns134ZOMvOAbrbN4MOJwFMh8ODiOYurt6qcqtx0dIbhjyv
R+zsw/m9WDIfPosOZTIYkuUWvQO4S5QR30jM6EJ072Mxve/nbwyt5vfVucSzVPTuicSLjhds2MRZ
aN/Vblcg08zXZucRd8uEgQ7h8OLTIuzRLhuB5jMqpQoeAitfD3BxKzfg4G96KegmuuDlBRAJVnsr
q0yBf5xY0YWEOY8RAjyV66gGMyn+zogO2G/ZBVYiRIPWJeBqxq+VDLRmTuSZdyoHaPMiVqMJVQQB
yTKmABpUC54SolEGc6uBPUmdN29Pnu3AhtFO7bz98p26o2CSvTvCVubNH4qsSnHdBUiGve+7Xjzz
Cs06cslWbb4bEdAJADTVy1HzCfhWAX4m0g0bOj9fJ4dhwYmAfRjbNJ2OSLzXuWr8twbdgA83pNLM
ImL3tb7wFIBvx42pcdn56n+a4gNmqOK1fg6bc1pulYSRHBod45BSjejJlIqPuq3IZRskQcPC0IQJ
0oRTzqrmAIl5OGWoVy9VPpid1TNaKu5iUisYDpsvUXy3R4eKzwObrjULHG0R/P6WihonYHObCoxG
+N3FJHoAKxUG59WwmGA6gcVD7qZzIZlemrymqLZF7IWITnNq3oSqFFreBzPLvYVv6eRd9xkFuumv
3CyPYN24owHz2FsNT0oaT05am57rL2p7pQmu0t9Q4loUSlwN/eBRfXyj9qHMKtv1ZpRiHdSgPzVH
sS1J70+SFnR2oNV+HGa3ocxDvISufjJD5OyOAqgS8rzVIw7r3eRbOpMsUb2IbpmReiBVRfRUOigD
GfAXD2ogLPwiNp6Zkf1jjP+9YwsaA9mAy1QlZgHIuoAStlgebEsZLAJFJsoefcCfYbeNGHqCDICT
QQFNGvTEP7OnimwuQfMQXByS7aKl/ZJ+FUC+JN8ajJhz5W7xd6cXcjAdNOlJzp+X1ItmB2rP9Yxs
JJYC8w7jYz4Y7BYahmv71AyJ5w4tmJ0JApRV9bDjiHvNIlM3/ZrFfl+yI/SdXyJsb/5wafgLQG77
yXQhZ/IAHbFEXf8Ep+f5k2JYP9KH4q9Vg9aYKEAjJQlc7TaCtxkyZgdl2kGkuLiUbVOA233QHoqD
ArcJNosomCf4ri4Q72yEbtRmQif/yw/FAu8HBgDZqTlSndFbKwjprVfs7ve/K4XwBLL45z0qD+oE
dDVW1Dr+kRTPfZ+UNzITIlum7UZKXThSMU0tkHFF5Og/hkWvCTj5sAah6/16yBXK2vLxk/qPQjGZ
tZeOwuQ8rXulZ+MpZzYL2t3f6MuehKPX7AZHohEz+pKlRHv012vgi03SALh9kRLTAwU/MkS+GqZJ
QF32pvUUHZ1GEtRhiw2peKpJLluNcFT+tejeQlIENbBKe43E8bSO60qbmrfR6NStS8D282bIAl9l
c31yDLT6ik+I+gSji/sH+bAGoR8ye+mlIbJUqUHGD++6qwwuIwTIWiILHz+I5Ul6SjsrzfPlitLt
1Tu7vHrVN2zwJpemneHhDV8ThFLVeaZcmcgh1iCd88gFPenofXiCDsUwo4FKlUY9C9imGvKIO+JU
ZNEEcSjiMBXljRt+VksABP0qFIIY3TWykdk3L4HzZpiRzSAUOCjcbXTsoOMK1kNC98z9psVwReZg
JFYA0dWuzC5RzLHX5/sZs3YsJSHNZ3TNRgvyT4ti8oQ+S67T2enxSo9ubPObPPcEZulSvYKh4dJ3
jNYrEmPmb6A7noFJldg8aAgvW40d+kVRe2RSexqYIolkD191PYSMby2HP/0Jmij2L0+q84AZ3B46
1zf6CbfJ+H7eSzntRUCYIV8cLEQTbGmCmSXJx+YxBBhtFRRiagyBrE9KcX6cicql9LDlCO+bhgFE
QID7zYP+zk/4HoCQKcq6DUWY/Nf9/T7nunjQyFwds47hfJ1uuOnZWsF5xtVgZxlBml4+sRLcvgCJ
In9eT8vfSGO2j9fYS17F6/o/ElvLyp8zbmzHGV+lOMTLQo8/sEMRhz2/emxz9VDO4NKjSFWEgWoJ
XbJS3d6EurPAce2BGCyOtIUgscq6J/TTHYT0oy1VyDj4G/2GaHayiiHpm/eiNHZY7MF9xusTOhHf
3bA8G1f7E4DHygDlcbhv/myVr/QlZWwkSDQEnuekl1jUdlpXp8gbvjx33Hi4QM1+3452+S0oRSSj
vIaWd7PGEgv2fkX/0WFCRX2xqmT6ahIRsR9jMOBQw7PyVS+bj2XT3OEZ3jvFGQNkMgjre3lTU2zV
7xrCwkIDSJLbbshkZPoB42T0YLmM3fFvume2jwZ9+SKKWE5dG7kqTwofG3Al0itvX/iG9p54W2B5
67Wfk3x9rbxj3Er5LgmO50cM3iN3uFLnT6s2003O1hu6bU7SsAvl/AhhVD3dEFaIALhOk3oSzUFt
SRYj1QvLPUzLnPLJEGoo29CPrxl3g+kFKW088jkkdUu8TEB9C6XuR6Gth/nzhdVtl7iGWgDblHF/
gWROlf95l1X1fdPUGP1GSwwtCRfIrRQEuB9ok42Dd3fD1aUsbeBVW9cPznrz/ZKJyYpUIR9zL2GQ
x4auAWzNdVeGJ828aqNvhEmmtPwFbXkKYKV/PukXl9AGBVUwxnY6toQP0+Zcdz5Ms7NuHM+5467j
hhwVH8iLjf0JeDkFbqWyCZm/YZN7Aqef3GKinxzDCP22fsaPAdRLj2xshOiImM1yJwDsF88qT8vW
cpI92pysS7WzQQF9TU5r9DlEqSSgUDATrdyu62ougVjt3BE845C6u5LSFZN80qiW6zi4BjtL+WIt
uiHLvwBPWcEa0IKXEwel9LKoJ8QUB9HiA0zi/3MWlxO+uMCBG9Q4hFnaHaC7+syNt5nvDTQaeBSr
lSckwmAoo2j7+GzCH0eSMcsTa6WeDDvQysijt6FmKtgcW2FlcqVLh2JOe2rcm8o5BRtWuqE2fcfI
TumYsD7UcbhEy0qRhgj6ZpNeiiMNEisT6+BXS69l9UNFINQytbCvZLrYkxqvOz8a+WRCXt2mDfSN
JkYk1twLvOC2Oa+VLXj6zHVMapKIJpm0R3PkTFs54KIcDrUVHyokR5imXwLIy2fJB6f5ByhtH/8+
CfJ0DgplVyPUyaq19aak3L3NPdyZ3/MXnqdhS0LbCaWcx6u59ieoJxt9e3EVBaQsFGZLZMQIlYKD
Y+cjU9F6Z8t9P52MkYC7TpGrXu1bDB1LQp8p5qzT5VafODkMfctj+SwgP1u3YPscKDbwZ7PB2p+o
N0VRKqzZzEjNB1Ic1Dxz7Kxrfz6UurjIT+dZmx36c87tayZIxTdJVJLVWvjmAzh8VBwADaCD9nr5
13uoF+iqSVPLLMSg5ehgNdDNX7q1zOBSqTE2+e4PUYml8237qbCy07W9i1WCd5sm71kgVT4wCMQ3
sGnet2oLYvMO0GKeNHmhXM8s/0RGIB+lvEaJZVTTa981xRkXkhvyOcT/CimFsmUnMn6jYS4TfZst
bf7ionm9Y40owCAT76YymRO0/tOFEjLsbj8QXfFT61lcSSGJqidd2IAPrLPZv4B1vGg+VzSe31Vl
5U2EXHvNWcHz//MQ+rn57u/X+EOTg52Q2V/WO5fFv7rI5MEsOy9EOwAX64WF2Tc4YmBGOCC+YnXB
bwA/K61zt3gPfZQSAFC/OJR4icKSIO1a5yfLZyr/46Tn5M8eJkIJ7VQbK9Vb97f8Gk3aXhgNuDQR
JH6JIcI4PsdtlnzW8DqcZ9jC2c7A5jX2Y9AWrWsWIUgpQ/3LoxN3TTiGighyXY1uGPtky2jK7K8n
/QbhABZuvOygbXKuZl8p0p+njbHhJ8Q8CKuqzIZdiM8gETo52Dyn74BPwaPEPEDs/2lNadQaCI1M
xep635566b0bvIu8po5GOXHw02m0wn7WJK8ZI6Fwr+mv6x3nRIkGU08Iani+sxYoWXlc6HyyJ7ES
AlLBRZOEsKAtNl6KfqMemScaS4ovzg7R/XAuy/7sNWrrN4PkZUYOLl/ZuX802F0huaEYrhPAU0GY
nijZLHH1Z0zkAFoSTw9ReaiKYEFQABxMQZmThrkGvFT4ALgMLCvvwki0vnIj3QGKV82mNltyltWH
QGu7Ur9VUyueuKyKMwHuk04aV/AbBT3eNptvawDQp2sAw3U6oJ+Hrs/1qQ1v6GMoNmhSckzCLYfU
lcUJu0V8+PlSO+hP8rRmKG/qMJggW/ma72SRIDqD6W244XWppcwLUjKqNIT7NYv/u+seApxkjtRt
fAVcw8cK4JDbSMnv+3F4hyJ0DSVdgVYB/Ca97zeJhHmvLbvpYc4XixptgAkGo9sRQI34bxZcPz/b
3r0RrWMnD/2wx0ac8dylH/unROx1dP0Z96fn2IjQSxTmM+5ZEtyIJsdc6bckSkiwhn41GdDZenla
gazIui8Lqka/AR38Jvv1WOJTbBWZhuD0aywwvCMtpQA1MtvI4lAMD4mnnvyCpcVesKVxueMSE8AP
Bo/HOm5kOS4waiSb0LaN0TPe9Wv6kEU+lUbYR6cLP06eYo8C0ZRRDKd5J3dyqgS22mVmoCBqSjR2
d0KM32SldR6wV8r6mE+bGPIzGgJ0u9c8aF2x6evbkLgbu41teZa8KVp3nLJTYpJ3brY9hEFc9W/D
FnFamdA2fgD+uYwXOEBV7WIZ+gVK2QdQPidMuJIM0/mSMKrC6dPCzyI75xoRGf8dObDxU5HzsQrj
7d/h6RiZARtyAvPSbVqL1nCr400E9ID+iDOs1IW1lXdxiBBNtte9zKQ4XUTuKmiziuMiVai1x/Bn
xdwBtckY/RZ8dcWscDchCFpMcazEZH1KZojgWv2PrVEMFe+2RnYKGMiVlGhekhVoVK5jvn7wTvzH
OGmDbTG7WjmsO2EcHERoiScjotUE9wn0dIXdpsLIHWU0TMhydXYq0ijKfBanTajbip3nji0zY2NB
xpHSVGlnATv8Y3VzU6RCShUS0KaJEwKS3dPPR6KYzgBqchSyzSttWk4/m37HOEWsUTKtOqA9cUrY
rZPiQneojJJkLoQBlKUQSDHQYIxUQIHTfTcQBi/0X2AtRPvt3OWoVX4tGw8Cl0azHZXedNQ3TO/d
swHzYojGfPnJyxc7IZKmlIRnm3ktpoTo9e4QR2lOhGtU1Jr11SWeMqu+Xq8KzyHIPCXbPXlKfmkg
G2s+R8OG0diocpEiSc6u8NnUNLmj1hm+AZPHLCV5QdKG4Z+ZtjyChkKfUmwYLCO2obeVsd6n4PE9
jV18LJHpDqhGhrh1Kg2ECU96rHIGyt0ygkmMnKojZaovxDpprBwAha8SDrTIBYyL51bFLhxA9oVT
KFKSnkdAvWBBs6AFCQmI2p0QWX3jwjzAK2ekkVjcPRao2Is6h7L8SuSEe1CGp7u/EKfSYmfIKnHI
d6K6rmRaYdQW3wYDMlWYZbVjuXjQVH4fBupjEduE4UULlXzBf30Yne0F3FZkwM8q6JKcheTe6HhP
/0FMlaHfEM8WvVvKK3LXOxX3zDT5GSZEUXoJwx+JBnyzdvKbnqMCdTaay/W3zuRZwOXkg1uGwgdi
A/kbYo4mYtWQ79g463RSI2itJx224bSeA0/tA/EprZfkKkZ3reUfI8FoZc0OrMxEfq6PC6Oi21sO
POD+cLFx2PbDgiBXY7iUu9M3X851z7a+lAQHl5GvFf9ayXgx4Zl1FQcGlzVxqh5OPv93/U40Lz2O
Bg4K9/7Dz+Mr7yutebHGxRGcZ5AFUbX8YYTAt3lVWZMnza3nxLW+7mNSYyM03zBUd9W0w1QXAy4E
1OyFHzWhslE4mfwPgrIr6U2GJ2WdgtiuG6kGlzWzG37oBYKgwf5kuOb6nFtMDRMAV71ohWKJWwzU
6qHtu41WSD054Bhs1iKmLCHJBYk1WXjGPPttw+pIhwRrrDPBCAA0hbD2V2/86aaoBQIzkeTISZJm
uZTnDq8oRN8D9X8K5nBidOVjvuWFzEskVlUaal8XvVyhXTtb92Hzo+YFQPSWe0dJijMQlS1uzUC5
YYz8vsnwuLdAz+kHHifji2hCBOlFNTEwlJofZ71y1p2uWfGtB4VRV5TqF3VEsBrQMpIocBn3sezo
GoEws1ud5DoLdl+E154lOmt3X2xUtV7vuamZh4KWWQ5H5rY+pEe0xXH3uCWuAhAiT3heODA+zVa2
hGT7BlGC7Oc94udpSWjvtoLC45tpbRLBN0bkRBxr0OO5h/1EJFLYDxboshFxrJL97lkO2UDNMYuZ
68jXEAcjbEkeYyF89Z0v83PscP/68XKLmk8i0mzXks8UhMhQQGGHxP3fw3B3lx5q6pBhIY6lXvBT
x+lCrLWrYR985MjtHdUgzqsDqp6pK95VyWrmb3ap4Pm8jN5dtlgP0Z/9GvwnxenUnmiyGJsaA/sm
ZudBTECFDfjDBYWtQ5smoNNy8SHSH/tu9Yl+C/kPfBY1dORf0Ax3o06j3LCnfJY+rU2bhHlkgNz7
wo3Zr7TWOCGp+L+Uq1PljLsIHdXAaEXY9elcdl+RiWNOVGdN8kTHxuVCwIzJd+YQmt4IVNEnbNs0
vC8h0FDCy/dQx+tXA7Y0T58TVWqn4pW+06Ui8CVwzmYP36V3rPb3/c4s9Zs35bExbGZ6C0g0OIUI
TJCEpvV6+MhY3DHepAcI9oluPOrilgAcr7/deZty5SaFZKOPipFBSoEHrgh4jWmDPhe87DY2DKSW
wzTDzrB7Jo2U9jwDjwpYcXOltyD32a0rluleV1MtqXrp5BkJaBSakZZ77tfDNI/aIO6895oenSlG
HY1ZwyyRlXpd/jQmvUSZSTqOHYhJnR1qVZaZHVED9ohhH+TBqmE2oQLq/gXRarvPRmyZMDT3CEcJ
b+eCmZZSxXpF+AtrJguJpwCZweIrtxsTvWzEEZkhOyETRx904srhwsjW8RJ+3/EFcqr++x9VQdLl
Cp3kDw8yza6rbtwqcRyGdlAac2dz30ECFTgj55PsRfK8K/44Ix7UhKKajdihnKlMI02kwxZJ6cRO
C0CYBlaWO3AtHRWyyxGUvVAu9KA/iXMjQ1ESg2CQt2qxvbUvf14gIFeprCloUwihoVa/bEzoZhcW
Dlcm62B0Xe3Ca6u3fyd+MjJgFoGvf1SOLMtU1GmEuqBaQos14dvHWeXoqS0gdai/jfXz76vkociE
DaJB3qVoxwgmdABhR7lr802PsAti8H7w1uNZkYcDLwaOjKUirokPT/nhRaIg5nQ2DVYBMLQqVRoo
1yb9J5n0FXTmMh17fnb6qmGx08fg1vDJImZijLlJEM44SZK1CdPK5h4d3Y6/9ihgz7W9aADd+tqu
SqbmyaVSN0Irfh+qvr6GS5T/rdCB0dW4N1WUEh729Hg5/HxOY/cdRP9sZg4KOasAwk3ZNwaZSVMz
w8E8bEVwB0rFOCLAaTdVnPp2RgS1j9ZqVqVySSFxKLUDzTWGOB029KGx018YiSUOxu0VFg62BZ1K
4YscoGv1oxKxiivmtkOmOa6G4oZGqLfaoaeSLV4lKpT7kgaKd/jLCTdSQv5ZBOl33NC4AQmMSgiB
hAY0H5ok3FXJmns9mh60n10Kg/1gtk2342r8qDkNIQ7GFeEG/f2fePcO772sO4y75fSd4p4DwFqb
V/AVh3YQskjSisFPGYLix6U1EgC4byETXomRy+uhB38K9hi68iUu4VeJSnWn0oxfT+OfkEr1i1m4
vbUwna2nL4w/I5+pFgylfhM02AjqkjJgHhCi1C1WHaXdLMtjJkSDBurCrNVlMhFl/4DrgYayHjv0
4cgpVIFyhXaLvJyjiedUJogFs9yNMcEqNlG8bIUZ2+q053XOxmOTsZcga6GIrNxs3kzY+ez+hYUt
AAbI31Vh9f8QxT//ioZB3Du+ZVpGKLCMHpgdOowqbBeaQKzBrQd/GunoGfyOaxvJfh/WI9Z5fw4o
9i0xEzPtRz2mu256fUhH/1G1TbuQ+WirA7Jajq+1MF58L2uzDqVbhvcXBz64uXAZzV8YnJ+BpkbD
mmT60modhNdXMOWAZu3ARlFNdvAp6X26mZU/Uyp7B16BM14RjSSjbVTmar1lGW4iLbNvd1vYVsKK
Z6KN0xHAp+Va1jn+kJPykq3ll16pZ1p7eMpaT4H4ettHdEPbJgu7VquYVT6989UWeWeWA2QJSs5C
MS6FLtnfNXA73qmLd92G/SRwxKFnPtPjtloh8Gf6+l6UGjHIBZ/AcC+i4dTVXWhQy85/nof/F0t/
klNpX6ExR6/2pd3eDnOk7M77D0iQRiHFwCJJgtCWKGY7E20c98bxoc13G926Q1VLfbNfOoUaG+3C
o5f2SBup7MxapLa9a/wjmxD47Y1kOPKg5ubxYESShQKLzB7LRXjMlJXIE+PyKBtRBaCgwJUdSuhL
3Kgdd80tsuFm6mxqvSBa0PHFgamgjPSOCsvDAwxyIbxoosPISf5S/lOqnuJBdmL8bEtg5rYBoYdL
OWT+ENv9OGfy86O8L23Hf4fAnJ6MttqJBTg1VnHnbdAXoadQ8FOzpZjqZWTiAvH6AtDDjCMw/7Fv
cQJjeGOZDmz0CgJ7WHlo6NRnoM0JJSWgqS63U4BGQ80yrPvbi60sTp53CFvdDYPME7aNDkh88GI0
TTeusLwn0J/OblQc0elkJO+3H2AM/MpiT3xO5HZsheeVdO4tLFqQkC23MWkvNoRdVp2blmgcOSAs
CJRznrGnKC7VediGXY9LqX/6l8itR50OhYwZLFhmfgphYAufnN4IzfLvZrAj+Lj5BvzUHPqwK7H2
0b8Ugk1f+jQqNlgDy0RCuUQypPsx44zxxEIXq5lIMtO7Cv5tQSlOnQce/j77sx9WU1b60OeGAbvR
hfm9yIy3xhFEVgtrxnSfBq6DQFXJs0UJo1dGZM/LzKJH1mu69pJdIwrt682V983slA9ecCv35KCU
TkAOfvD9POmeiwvs0m4YdNQUXWFB1jQiq+qXupNwCdjNEMUVjJ6uCTxsDuEW/vmlpmGst4dfdWSG
e/B78rNQeS/hnbm6qZcgYuev1oRVzKIkC0vZ23Cm52v+rXNFJAn9aG0Y0NK14E09+/sUejbh1gIh
dRdevT4Wf8m2/42oGccR8cVFVnClMq0fU5n7coeol1QSGXqRr2pVy/k6NBlWzlP72oUgj7z48jQv
VF2NklLW7FTwX/bupxnazOYHZn6mgIEAUXhjC6C5TXuNPpZdwaCMzOUntzGDuz/rHYAuAQ6Is96/
1ewkrldYgwgzPapyAvDPTCV8aOFxz8rOrhymklVpE0BwTPDUfR/MtYBoJOV9FNXWput8pM7aa73K
lxEtZ6ntCrh1yJqMkAzTu/oejSVWKnUQW/mCOVb7P/f9vLWRGtRqctMu5VUnq3CqaFVU2wLXYI+g
e6YbjrrXoH0LbyN0n4NqqrnSsQ2Gf8Vto8WKn9eNEp9KZrzmmNBokmlBagx08wsMdRIH6L3YZhgZ
1bE3GbzTrdhwBiQDEM3cnNa2UDvafijm4TwagVhDoFtAWpBphAhddo/55oCeyqf/eijDLC6tAmfL
+F+M1cnJwHIbTDI1ZpEtptn90wottSM3/vqe8lqR1CA7ausmY1Hr/bS5q7rC8/kMn6tsZ6QQWj7w
LtaSY4pketuLkYU3mjQjlTrDo2Ya8aJ2GlTOM46ZgCFQHG3fX2YaNHvFWRThgLhVJ5HojDDjoWry
/iPP5G/dLEu33RiTKjgC4i6sQjzY+VDuVKjJolF5mLxuaqaKEMRYbmbbnA5cLrBL3T3cCkJSGY/9
DTANu0Y0FwSL4p3XHgJpuISXtsn/gt9OUTM3EJhtKnVf4MNM02957Sfo6OLwPkPBEU9nTQ2cXRvx
2wSi+35RRREKsPNahIus5PNbJWAmXatbJvnalQfRBSiIhlu1Uq+U0qN/jGZ13MxblbCvKnRMh4jv
E5ir/gIwyN7UxkbNztn2fjMfpFtDE3AEwY950U0SwiV8MnfGsvzhX1bEryp/OvCQ1dzlo50HMdhx
ysDUjX/filuy7Hsc73ZFpS1aHOOwkJH+TRyybNbjft4QT1PJ3Cv7WVNzTuSi7pc/O3YXOH3P6ZHg
FjW3q/QpOmnj6MNlXvbTU1okv3FBFocRodUVp1w6gQmGSr9H8U7yBtKuYcrRmpzUgruyh5L8XLdP
qFin+ogph39rSkBup0lYAPWu6wy38XeBsNdGy7Nli89hqzob6+WZDJlV8kUrM2En3XsS2njlgeim
JvXgIQChk2/if2vx8hCLFU8teLEt6FOjoZNwUC8hUFMQTX8k0y8ZoVFmndgiPOQ7mTgqksNSameq
k0ouz7U/ZMXpzgZTWz6itad/MX/7XggyD5alAXC2b/C8qAB19EbARK5ax0wWnSip+3TnHBak6uZl
qx4TtI8v1aKrdvBUGMCwye8mOO0cNTIYaFj7OJAzyUuSrEMJCjghLIpmyrMv8MJGGqWmYDzHUZL+
CBRrHI7RHbY1hA3i02MYf8hdPmqFcLO6XQGVsswKtBtle1Rv1Eb2n3XD8i9LEoQXS+8IYPSkeraE
dohZRFf07XTfqUDRKyQ3FdJeTLoholHEA/g/CPJoxAlh0fohOi2AbBPwXQ302csX2qRiaXUtSyXS
UmXsHGURF3ut8rpXvD2sbdreqpPn1DAgMQ0SPqqrQJRYjvCjml9gbwGnWxblPvGEZXDVr02+Ahzb
L85UEWnp694KgCPaal+RQri88SlI0zMZZFuIsQ1zXK79Xq/ezDQbFVX8NOiDBG4m6t/6HW4abT8b
skUpy9dRfH3uRUrcD+w6e1aGLvG17E8H0YCUI8UF89V4FCHpyr8n6RMbpsgsoc97M24qOeb4JiY/
hQgte0K/rxHOGRtowRW/S7+2+VbbXCRb2Wq5a67yMpFVzNIjcF5P4MXnz6XLtwUx3bhyX0+iqbkt
VU2XjtNU2hFNCCgVYJexsisaYl9g3XkgxzAj1bn1ugvJ6yt2utYyUZWEYuHATfUmAtqdI1hQoMFd
DButn5U+IMc6YiAZNGJa/z3UbGK5Z8GnCE5MVIyMy0joVlbQbpkfQL4A9/MScNMVaUKAbFECExuY
7DIOl+e/uD+RhGP40kNa1F62SGfshqNqr1ppVZn/iWzhWinOOLUj9jG6xcG4b0IoUKyyTK0aXhHs
XxaLEg8mChvZ3UuAlX5pW3rxQNJXbEbCwPOdRSUG7yjvYbgPQeewN6zK2GobBQPbt+l8jeRnMPTE
u9vOMWX4CGYhrwne4znprulp/BMDG24vsBUdp2+qvjzJtaBZBlhB7iPw2zmaX8SXU0Lo5xr/O4oA
wHThOlJQIv4ffcG2HD6p/ZofDxnwWM/9HCO+8vfzhynwP8pTR5spXyaxyLwJeebtn2b+7i4Cqkoy
nSHJwNIK6p0vKZBqfILDpI2uj9oFPfWQLE+RmxZQTOWux2kwa+gtG/8gDjU2wEgbZFfobzeYJIC7
Z5ON++8sweYc59gs/plFriI2qHgaatJplWyR4STmcK5K9UhKe3vSU3T8cmgUfGAzTUeHMS/7Ptjl
hbQBw3jlUcmIWkqMr7iZtVAW+sfUQJO1+1kWMwiIwGEtBoui1x8vS912P0Ud1doC7YQqNjcF9YKz
YqoMrMzLEG9ziRcRSSDrKn/Cz75EnkuhJjCBlvDRV73tjZfE03PTkmyObGVreX9XLOzEszWXoQDq
z3cwZ85wsAguaT54qSgAzw0vfL/owRR6lhRE5rMshKiY4kHgZFcAgIC8DmutIVHJaC/9XpcJmwc3
ztR9maHhzyQ3EaxBusax0/djSfcnblL5xo9HzK9HLDqdl8WCuWi4JRTiQSZwlM7dBHsJNgBYRq8D
Ngj78X6i6Xk8JWaUMVkn3pKukY0nyn9bRPKdrZXid3Vo+9a+gbusZDshehsXgt02hv3yigPwY+4q
18RbA4+G8NPdN43bxhxgh5FNmlmQJV63q/qnrvVxGd6aP2dd9702xNaExXy8PIduhVxNfakR3ydZ
6mOz0tj1U7HfXZkFWFcyYoH1ZGoyxtoSfQqJD0owAeYoLy5taUqVe8ttvrWDCNYhdieUDwn8rui/
UvKyMCqeRrMNdMIDNiIyqyiVEoTuBSITgmJqgPFO8Kl/NlNXoiTYPW3KvclsW+3PeBpffyGdVBvt
j/+kMWmcToBenhv6rZx3gkVrr2Y60nJ5t+A/kIjPGU80wWuwJxtHUpm9apdB5YCUhN8vEuIXovJZ
dFOFQlOk9FKBtRMHgZVimYr+6txIIej40n281LU+mCbtD7wV7lIkOE65Gzw1UPlc1EI/dmjm1PV9
QtczWPxCQtEVLE8NT+UlWaaVlbtc6KiR/2fyb0YGwNJotWQoXvzsVUtBXNlSzPjdJP+skaPQYMhq
ykGgC3t489YsMza8UDXYgMyQAuN1tN5Y6bdwMqTQbT1BP7AsF32/d4DLwK/wTrq+GGWt69crBiTD
S/FIe95cwN6afYGR+xuh2npZ+LnLMVxh0vMUZMoS8wq7eUCnoNg4DCh4t4pzeKpbmIohgbGTTK3C
hXv6DHailP3pSNbw5fZpRwgdZgyNX5LEOmOtWPHP4lKoqUcvGYDF5u01nR1kOHW2fO9VgRy3OEbA
sibXRN7kPDxJ200k9DWQYc7mEFrxEAnQ7HRdugkKSXa75q86g98acRuA6l+ET4lvp5sasDGQEtps
5eLJ5m/jSX0Fwxktp0KaVfttLdKI7YZwtFmH3xDyZArKCyQIKBh+XJzC8C0yItRjtHhCBRtnDOfO
qFCiWwNNzQEFr3tU3jbXDV8e6LMf07x4rdzMCTPK6tMpOB5Ngqz2eaMOUXAZucagvh7Cl8zdWMez
TXrE7i1ocUM1GnbQkWuMafm+Qh7E8HrIa9V85EiMMxXqY6hVj4QFNBV/RSzuLq7yDOaWrPRPSOzf
unJ+u+2IYajf1hYc2SueJOoa7FeElGBWqL92pOcVENTesTtV3mFBFsqTv8Th+iQTEY4Ua8lPai0R
rzQuofdpDiGVRUaoVobphvCVSG267qHGH6cHapOnm38SrSjtQX1S8GqRBMmse8FnJ2fSM8WUU0SX
gqMsLSAA3QvYiRxXEJn1j4B2ffO/Gij+d2Nu2yoMB8GNud6TlS28/ayHdQa0W/cRwvPHQnPBRv4d
Fm0oRxVKpP7NORBcy9w7K2QsxR95QvykoROYsCTricApZP/rWa7wJTf6Ch3MJYcX5+LwI0WTTbBJ
G8oMjSsVO0yxm09DpPiYemj6saWCuxzXL3sWuQyFu9dvQuHiK5n0DJxe/U5ZemHUkpsKD8Fy9XrY
WzHXkITD3M4BqWOfwDQdu9qifQf2ygf1TR3vSeEeTd9eDLCd55pDd+yiA+0pZ3h8aCmDdU+Ijyrk
vYIBwLzyH80MSZo5Pyf1JUiD+wtw81F+ODT5lv8K3EEZNpL2cuzvQzflXA6K3ERRuQG8P4YUq1xs
IricULna3hLZx96rgFU+6Zak8Ex5psW1n9MzWjeHmjpi7ZY/93zTueKwwbmPam560pWGEGMC3yx2
IlxBj8rzwc1bPcunPHJ5egN+V16BBwR1yv5VBCje6+0dye+xWubNji1UzAUs1G9kmpK5X84viaYA
iNafksYoEg++ZbfrFMyKrazVKekDaqYuf5e8TQuHHwo9GT8dzxbL8SUfwVqQ2vFZrp7bPy1A1Lo7
igBiIDbH5fiO7euIxhhB07kIWAaSsic4TmioSu5h3MWseDRK1FgGGOAWO6vde0YX2gKGblV9hn0O
Wcdgy7L7K/1EUY6Ihjwcx/YdwCsqkaoXS8t3Mi3ZBrGn5wgIkXvt4KttbeGcH8O0X/NWKoJ+k/Yr
Y0Re74a9UsqR6A7/lZqoNSPQPA79Fos7nj9QX8IP5414nFo88PWPFB2fUvQkCtTde03jd972Xefm
YBka6YRQxD4WOf+J5Mxb6tZQUIHjaOHaIfNhPV39ic+CtukpkoMRnbIAEVzbscC78CoaAQgD8myr
br+gO3/S+g3Vxjh3sAFqNUvRHF3nLb/k9lnY5sWaK1A2ckiCG8JUdWBvdAFTyANmmG2Xd76h348F
zRGrqVv34l8hEGA2O8UIZnfiNEv+ve7a8jX/SWDu/4ETQvD0IamOOdaN2JaNRsU5072ilAeW8Gsv
0vT4LmfVHtIWODS/eFN4/2k6mYmhKS1IJGag0QqmVZewyWEpvz3Vac9vzjqf4l0sooGfKvASNdv7
hFk/eUEsxQwcMqV11AJZDSo0iyk8MtjI+xHC25YtzE80NDZPMbJsaK9UToRZ8GgiUP0vEPP0We7t
qPoj/uUMZHJHI3bTvZviEcYpWy5qGF7CSnDTmDGwOOfzt0kzeaBgqUbh8LM4Ls4eUCnwgbeyqmA+
Qv12nyiBaFJ1Oox8q0tb5PDVONafKYeBii6ufwzIGz0JeeIr5SKkQIivyb/Ixz++Mrj2QcMeFX3h
mK8GgrU5jiCgx8tXl20hO7loZQ6L0RY28YFsybKfU7nszkWjmEi2xM/QFaURG01eomAWFN369Aoz
ACALS1YGAFYgyVvma7ztbNhrt8j/yDjEbOZY9PcPpXZGdAtgsEP2k4cjCBV8A5vnWhPmqdxaoNQi
k0/jPBrjEhKNWjI4x/8h2NiMM6Mer+ElKTfJG4kpSFiQ3V4zQ0TNaGhonUIWR364yTPbfwzMRxnq
s9OhCLi4CORcTh/3KFRIJMLAvRwcsD4gzsL/W1ETGcYfMdj5yXnjSCQLxtQdFcS7HiHEG+Z7A5n9
Cj3eyF9g+PKIlHRRKpwi+Z0RsgA83eYnXLiTWYut5bG41/q4pDFe6kK7L2qE0zyr/I2enS2BOlPJ
BL+m5sm1qWZkGQZBEUZQwYEEWy+QAPaxxmo397R6l6lzpOBBKPuLbTJRoFOptmi/iJUFGyGv9YhP
Q68dNtKH8r+GEdCJpz+FJwD4dg3Numh8hTq3+B4Liq909WMSX0UXpsmUkv5z+VL1ZVmIS/cfZ7nk
iv1SZ7w5vC5pgaK9y4ia3nNF7ynAeFzhrVAKUl/wfcWfdtcKI1Zbi3ptLJBQFDkKgqqY+c9XTHyi
x7iP37aLJQycdj3+7jKzxG7LM2C4SaiwzoqTP4UywGbYWzKT1X6kCFUTKGH3FXbUY5ee49rgDMvc
P3C/dfNJokmUMXZgkhhG1kd2zpki71835e/Oa0FHqN+lkrA5Okd78yUEXOaiL6km7xmTzmLDCLeW
KKtkA3sY0Pywh6Xs4iTxiPGnZQzBFXaZrPREX2wxLENDcyydjsgEwLrCnUxdP50UnYMq5/cYspfF
HC/CNUE8O5pYAzsUIs5pOETPlkEbCmgeEOUl07KsYI/xqrBn3wiI1FvMemHQqF0q1xATFb4YaqYx
M5PNBv3pmYPEH1PN2Ha4rrZJ8u4vSR/814SSIbusek4BFLMj8v0/4eAJLoviGqW3DjbzXozwTYbW
nzTF3q3RRufuNOxQ231A+SBzoHHrtfbx1wZR5iWyClemfPZP0PaVm3pZFOniyGpaCwL3Fb1mZkWD
rNlCR4anv8OP9jyG+BrIOkjte7p4RYyzcL73cnPpBC0k1c3zA9RSxk+IZmJsGpdVoppS1UN8OUYR
M6g6k9DMdIGF9Yxv7LKnSNp1E6Nubrvrqd5cNuhCtDkkIW8UaJ+4mcs14mz+r38xt37c29fb4/4d
L9lhJGPVcbTJTFtBLNlFmszCVAiBCuuc5L4gcF8xMrHci+7ml9Um+ToRVSzmB11PWOERFEyTt1VI
3pEdbznq9cw/k1xlq9koil5xHLPUs6KG1V0wtXEmRskI9cG6uGgvsqT97ymSG361TDOZ86YABlY5
++/RK9WHL/SaJc6ln8I1xuRuh4gbMIEmBvS2rVmutkJOShAXfeiaB8MNoj109d5fINVPYaANM5//
76Iy+3KxmMqw+qWoQlEvnJcAO6rqYAOn1WfJNkTM8HyPb6ElK+ghIiY9yO9aPtYlGRx6/uthQUW3
8obsBaS7/MRXDmS45mFAuH8x5rHAdJuwY7ksIV4pcnlmnSNO+PxgL6cdQh3XSfats6ueTpAjsXj8
XPnwERLKleM844U4lnMuLJC7ao+C0brOEvtx7eOniqI6r8nbEfPNWrjiB35MxJJKidT3aJUwrSuO
m8u5nA4eHFjUw/BZzInRNea8t/48jdWslkf+eB0Pya/vAoX5yBbmPT4oTTqoan/SEVbI8LzJYzD2
orEC5LMgAFeOW+W1pvCA4/ygJdQUQo6+2mRU//+B1WIWs6RjgCOA0vh+1Ata+1nAltzuhqRG9Lqi
A6XMruL+ExCFBCG67LXW71qjEJD8ZuZ9fE5bPXFmtEe6rExbflIiDqWnZ5H5G7vJlne9tgqJYHJx
vst4HPN/iH/4a4z+QfG4Fn0ZKx6TRBhOrnjGliFXYLtGZ5IoF3+3gI9kK58tsL2q9KoaRVYvkQV/
4eKT0Cg9FghW7VYUuTUAs1PKwjdnw6yy5p+4uKxUeVhnyEJ+g9y+bAyLOu3B1gQlpWyLmB0l9HQO
T5kRpHK+BOzRqlB19QUgB9o9TY8+nuHRtafx6t1iqUOMNon3Nj6ToIIvyLHby5HuI7vPiwyvDNvw
7n9aJMQMNgueebg1YNU0OhyJpMg6/Jaq7Rp4pNns4//nNDFHqNSvaLO8ihrfYNcObvEL8o8Pzyn9
Dj3hvDDdVPqL/Lz0B9PT9SFBaN19gbmsJUd/zsi7FPQzVrsKcVvUNYkjy9O4D6x8FsLW2cvtboIe
Tab6jVu1O26JOyPBFxWE9pgFuZBR6RanzZtOkemYM6HlngEq56uvPCCuR/ZmTdLgBf2qRc2RZBPO
91iLIzdCNViRkTl+q2JFU5BZkgzVmk8ZgwLViutfH4nH04u0QdhAsdOul1rhyb31iEssJn2hQSYl
LJRvYSPjNQ9uAFf8+YEBQjFM8AoRPt6cJv7pynn7vtKWQj4+raKSvek6zqXohFoOq/8TD24BdVgF
gtgQbfXv+1Vqv+x1X9kXqtjoEmPc02piV+trbwu04nJZ1WwVEGlzaU5JuK8ROXcivnzb8Pfw8ASy
Z2BAAJJCty9tIdwnXEOEXe+6UXv91HwSRdCVoyAH4S7zy/ibhBET22D2jqm8zrcdGiD8HFhDTF+D
oa8p+V/mjqt5W0or3brzVEd/UGdTBK4nd6vBHldpCIPXpPGwh10HfyGFTM2qO9hg5+2ztapEVh4B
K3OOhrQY/2xiSzV0ECiiDBTSTnA1ajcHGKxznt6krk905R9v+tJxkCx2xoxuAVkEpNsg91+hrPLz
hVZpoegKlQPM1htQxySZTuxi9hrTBzTMZHQLNHuTDW5T2XCDbY4IXR6dl1xMy4X2+wcozIYd9kt5
M2uR0UMpyM/aJZg2HFtyn7OcF50qhWH51xk/rn6IkycDEn7ihJ3/HvXPozGSWrebXuavIdYE/Obw
4ww4dYyY9wDIdTynsa1PYJiLnyaH9KpehD4oND9mnd6VqSPa24lZtnQbHQSvMsjJEqLZS2XPTato
YBNawGysp8k1S1h/kO5SjWAnDC3r5hSG8Hyjn04oUgveOBELpOXfRndDZUjFe8pzp0ylZ/PSU7Do
QCohN/g2JfwCH/a9+8wJiRuh2T6XIO+9Qi+CnqV9TmKnbENrsaoenRGMBMHYqWOG7qvyfQVphl6M
BwO8nBfALJBP6IcQdw/mifClZbgSQweVl/rmlDtlAxGCM9dC1SNK0g235MZ+hREPffZoznzxDNxJ
fHA9ptkGTlcivY3L4s2RDZ7wuhqxxOa4nlNca4fo9J7FIfsTR8orQa1x8Zm07dRoKRQD6mmUG9J3
m91ZV5toERHFd1UVdzcg9M3bdFhoIhHlrhn/9R7yPcF4vMDl1aMmpVdfVmnZ86F3YW0kESL33DsI
MfcPrxtX7kU4KDN0+Zf0XwrBNjf6Kdrxu8DkgGkQj99U+5RAfqGFbFm2ayZWEjpCTwSfoCEO6ay/
PvOwiAox8nJi7UqvWEWMB/WX3xMFB3StKpOj2eYTM+6OBrlvFer6MvYTpZtNDzpjFkM73PJlY/DM
2EsPWaxdQmDvVD44sIS1gEL1Ah67jwzjp53Q2+rNI3oy6x9TV99xwa/6EfzLqDZfYnloyxLyzue7
WzAwTJP9g3lvEgu1gY25h/L66R5PAI+JrMQoCzEWoOd+ENx371lsH/13PB7nLflMqskUnj8fNRRA
llsbPXlV4sX34sIhaoNR7KtZNAZEiajSaSjrM2FIre2VZOT8qoUUNHm7JiwD/gNX8LwOjVcL0EVH
ltotcqlR+I5956K2aV/xrVYTnREYByEDUDztbgce7Ctu+SNWIh/luwpnzx0vSqrgarn+dufSWg/m
2+lbsazdekvIWJFCU/7sateIupztJoLnFdWfa5b9TGBoHMbzwON+QWZVp6sxlkDFDACLLGqDZUCX
gXrZzhgDtaAym0v/qkkBS1k0EDWRdS/jxtXVmKCNNZUFoKitQsR/ks5+Z7Ljv/6imJ1u+L1qtAah
Wr9JOkvOF6BIBBONc0f95ZBxRIZMuOP2x2TJP/Gf1yTZHk0oHG7mgm+U0oEcPG7SMfrUi2utefFG
YxnC4wFka9enKt2AD+rNiUVkq2OmDro0DOc2yBoRhKAnWbvFPtKcGkpxOzWmaisA954snFBwxlUt
klXxMrVeT1fHhK8utPl+kK8MU/uC5ZVOtCWGV7zZYXxHDQbqtAUVSj1WHkBIuSTE+2BgY7xqwcer
Esa6FfnqUrbw/oCT9XqacwICw2wGs+0bU/WMJ/C9B2xcA9NfVqFWibAaQ5hkofrvGDtv1GcA/LrO
O/wu2/u03ix2EWia/PhoTGNfSO5oRhqKJ+8VM1vVf5qHFHJVAG5iHpGFR+QG1s4KCA5VYsts0ILI
pYaEvmugO5ogdGTvaNkTko7P4Wn6y9+ZpNiWJfA4+df9qba1/MZh1/Z0y6VgacnFp8U9o8of5aDm
BFT7PHvvNMVsDc9fp4MaKdXyWxRV+vfAgKY2bF7VbXlTX5d7K/esyB3mvaFHsjH4fjpyGEcskcNT
Mu2CvbJypSqYBgDwFO4GjWvhbsRc84Px1R6GevbxsbaPzHHRq86OiQSOrx+3oYt1kSUssyIEh//Y
hik5sWcg4kLKVnMDUMXgZrpqix8rDKGOb2IDTwtjpWBmuzUrrrF9Nmqloorm/wv7lwi6G/3bOJUQ
ie6b19bR437uFud8GSG1CXqJ0RwMTgWhrx7KWSud1vVh/gBAXUs5vssfk33YTvUkWFqXwBB2NiRu
A++EtekJ/o6nqd6ubyN36vmQTSICz2L+ST+mQXl0IcQwUqqIEXQGmEkzVBud70Z64yyPZg0GDeDS
tje/CWQ6q7triaWkuosduD/wQIChA+tr5eXj+3TGg1WCnneZ/5wDJ15fFxk/NQYQHiRjg54eqzRk
banM/oLBJ7ZX8qW+QVlLxyYwRtXCuDcih4/3R8yS5jF5PRRK68hYGcwnm4suaiFsT3buvGbAlree
jx8fyiVo0Od1Nd8kkZfSrZP1T+JgjlIeObjyDDG7WuH1h409EKJYQRWZ3QbibffwSdK41XI07OUr
UK6Z5MzkhA5oTyJzqwmKfVvI5bhwiDa8Sb8ew+gjYxksd75NH5zT4kK4BbE1PFI0puOYFxIN40cz
7R4Syc6LkJKII9Er3vk6flo9NCb/UZtVyk5/HyOeV147SttHEHpUDZ4q4RKHr+lEM9WkrN2i+usx
RlAAdlvqmwA3ehfs942UteASk/5/qxQ+C0atF5TmcpQMfyMHLauh42g3+3yVZmxQ8DE4B2MyTqNc
JEeiddJ+yXE+Wb4LEJVEomq8ERO1WXjHtZ01RUaOtHghiwH7olzL4xSeS2hkBdeUWZd9Uz7eojqp
TZ1RuhSNoZCVatXZQy81OxVWaYxI8L4m3DgHXGHmxN5S5v4RmgxLK8vLqymosH2LiQhQM8Sre5Ry
EN0L05CDl686pITxlBTPJc4jJEpkoTpgxvRCMD/xDB/y9hLw1cV3javrrIPQp8E7eccsmtUwBbd8
5V7HCeGyE4YL1S1OaKMUWfnZweggzn5WUXIiFZk8d7Myj/RFncschw09JKlqxsnIEt4Guzt/MY+0
IDU/tsF8kOkJcPaccTmq8us+eeyl4SagyE503xorVWZngU8a+IHstAHUMIuiXcJIDIzk9lTpmJwP
Lwp55Z34cquX3YBbPaQ5B9cBADGvaGW8U5PC51O+4C2urG/Ur9Is12dcXPkzarU6Elvr3ukQCUqJ
h7Tzb4qdN7/833YBlnQIqNILWpGjSvuBLd+lgxRzhglSoAxFkI1hfo7X0h1BdXa4y5ItNIFPmsee
NKhkxxFZm0zKCUp3AiztnUfEZcQHyAFK37INu9N72n8z+0Hj7nVIapf1Qw4oPCF+jJ2ysnkoR2jR
kuBCtpvny4iSqDSXRbTRqRrMUM9cxz3LMCzJ/TbEKBDDy5lLfYe14asNhYlw2mG7FYt/KJFnX6Gj
ZlQk2eWjoiYulAm1MEw07zw76A5x5D8zCNc1wS7sxw6fcHS5vOM+bMOo9zD/optNp3OsRtHf4PNU
xNn7lgzBczjsCrXiKQIqKfF0hISa5zJzOzWRXor/I++K+727rHbpq52yGIZ41b8pRbktEtW76LC3
eJTcmd9b+9zn5qnWOm8sY22eX0cKpCMeS1E1CmhemOjqcE42vDI4Z+Tb0ka6LgO9vsNzNnFuB8AW
qUQOMQLi1io8DlNSv2B4SCT6p3u1FunaQHexRqB/QCS454so4E9gM61xYZVUQLSad2BCxe1MWUOr
XSZ7tPAKeBNlt5sztz48nfS+jzPoiVztf/VDLTrUuQgSkK3zChhgzHsp020fnVrqQKjb6CCQZhMR
qz95y75Le1rSONVqZ2ezFx4JmGdbud7e1Dc7Jzn1Q31vMKPM5j32sXN5Hm1JAMFItT3U+iz8kwaA
WvVHp94VDtX1x36Ecf8BwO/DMx5ageWVA6ezdw0YX6ob/0XK9P4viyrTItJ5nbXUdStrAWsbrCv3
sZ2gq/Tc+K7oVDAwtv7Q1naJohTJ/opW39x46avFg0IJdbA6m0o6wHx+S3mtPCfFN2sS/B5NL01i
GQslP2bIY1iVINqMF7kMmwPRnCa4BzV++t69cLQ/gDC2NW3Hx3niFPsEKubD9dwQ1dE6V/+hCZ0x
Wkr3UL8rq9maZBgT8h3zGzfW48XXfxbO0ekv5Aeq6RVwhmgaL5n55vtgLzl0mHdV8ZWmHP5XuWFb
0sgTYWTeYDB+IdXLJSSmc66vwyUSCxQF7PEDd9i+WqA++hxPenq7at6h9uNuoKnrWCR5ejENEIo/
UaBT6daBe0+3R3aXLGEMcXG6bbFflzjPaDIDSRCowu6uwKd29e/tiY0fCReYQAirTB2KMvwXrKf7
C8cyk3c2TMJolVntErLO+Z68UAYnZNIDjMRr9ngoX92hFS/W0uoTlu2tfGApqxRvJ1vRE3sF0Xvc
dP5ZYqP5pgGNMx3PmBAbFNyGn3P9qB9x8FMvvufscvVgdaFW7OOArjEvtlwFbAb1Ntsly5bYPND5
dw/051NRR9qABmn5yEAwcIPa1XJ8Pnla1DoKgmqeZB9oRV72luqo3x/aOWlq9+IyH67NTG9USnAH
dt0EpNudwU+wVd0cXJujH3ECMY4CrIMkgF7XM/nlZM8IrohKYejBVWp7GfHrs8aT9iBTQf7F5eSV
WPyJwnGUbEtJoYXFiX4Qqzrg5nmSv4syoE7s7UbDczbpXkjs62SoRLxxK9xHdH1xvV6eUFBQ5Pmm
32KuXQGGMIOzaoNJuWI+PS9US6W4If9bavIdNRdyJSXsJlPubvlrl7YCc9u88mgszN12rnujvSGY
2GItwInz3Df0dBvo7lbcsqhvoiMI09A2mTuf1C4uJ7e3qcBr9Y9jqO+gjsO5ohq6q/fyKu0DN6nI
JHcYJZ/AlKESTtz8frPulC7XC1Wi0qvo+wEOnncSpmpZSdDgGVGF/uyqj/Vg5b18OiXJM6NaNeUH
m63DOHdOmgSD3Z9NAvZxOLKt1mu33FnB8Nvpa0vEy9QUAj28mAaWoxK22ZjCTEF+grwfJB7Z32Cn
luxq6Tw5VOTGNLW4blzLVx3JVadFTTz1qf+7nSPlw2PsdNk3qtPAdYE3kSI1VD1Z1ARJWxLe5pWq
qPF6Yx3PPdRC6cCkgkMUy/WSHlFSAohilvAUTCaeGYs26E5te8gBuKwKnf79/dy+Kh+csNNB6Ibh
SnBbRYoEhazZjxRA0jIWSo5uIIZ7ebIz0aiMx7LbKuGiu7gtCEYesixP8hUjLTUWO9JmPxBK6mlo
g/G0/I5aU7G50+UWjnz/vJkVP38IvlP0iIcE4Pen03Fa85Hi5sTfmDKAUMPLsbjVOFbWgvziF2Bm
lCIjdjwElhyMi2KCWGvafVMxZI9de5BogrC2fuUJBsfXq9AWdW2OfOvu/+xyxQmbVcx8toD92FmM
Pi+wNhI88rd8aHt/kfQObWnAYfdB+psdDXg2CfwFKOUX73WCeEMa/NPVsFW8OUz2msLPDXecAiWh
hrX72yk1Y2k4IwLnBelJJ37BaJq43sV/uqkLu0QqmmFsOwElN5zFBAc1WJ6i54sLOs5QiU0/DmVj
HZOEMSacIvMBP2k7PSwqsokpyWNxg1mBV0VIBxB3i/IjrxPRIpxski7YMBJvj1SVLVjmyzwKqHPc
SoJGhlmh4W1Nr4ELPDub7ewGxwIlSPx1+22vnnRJt4tpurgyuMUwg76BE1wu3UAtzp9amIXDVDVC
0QTZvjqVpVaLwDWmx59yeFZyEJK7J+Jf9stpQpL/mioJMuMM2h9m+7MSrDc1nrSvVTqQjkWgnIdN
snKHjpZqJ9Ib/ec+OQpURbmoCbZVe+yJXoxGRMk8Tmioo9Mp42vDqbrVttpiw82kBgd0wj5ZBHwb
aZB0e5xaepwtqmG7qFIzlT31XiJoPuVRAjnMYMJr5tIdHGUOoKJokLvJOZOZxftC2D547UxtG1Ys
hhvAX4KpfQiQCRnXmAZkMkWTyLgZ7xtAwQmkeTKx9Fegilugk6OnainbXNBesW2ZttAl6qD/yerS
uTe5+jEvNO2T8KWS0HvNTQ6BCTFDJ57Lt2dqY1Qo6OUgNiE1/HU76CEcZsfuwUQw8jKSCgWrGGSM
hKN+Zba8uX4jK7rmXRIge1pbbynNJ1MEhfuF7ElfQtmKYVzyjQth/vJ+mFtK7Xux8xYN/zA0fM1s
bS2J12yfPGIvluXEKPnhaQoGRGM4iMtD+SmXtfUBeYcWm7mGJeGho2pWXP/AdLDSkJXphlQqW/Qh
vvjLarCYP0Qa1QD2jsuMdbABC74KKdjU8nOe86sBo2id0d/6LLgdxGHrIrt8kpaCPn/TmO3EZO1c
MJ5+DJ7cw24KBevq8ncHV03S/kzCoVLyTQGvH40K0rDywMfw1lIbg1ndf8Kdjf4ZUWzKgUdjRNYO
QnvW6RiLIDWSAkyIAGBh9GuV9YEukgSL0A8OVv7jB1uiG+4xZ9JxeeMupEbs4Yhjb19I1MBTPDHQ
as4mnKkoYSPncF4K9Pi+oDZOho5e81b5YKVvFQL6GcI5DJo95G2dteNlHkp5SbkU4VS3KH0Xcw6b
Nls2XhQZ1Kk1QdKPoEwm62LEIh/OLwVZgonscHbHwLej9lm7Kv8xMWY9NM565Q+KafZYxcrItfLh
S7v3MKHHDxDv2HhzaloD+RBhcQoClQYv+ZUMyhaj7Z77AxCqvA4k15S4PBU4FaYPDXYUbrMJkNmE
HOZXuPslq/GN7rfmqSoSBBI9n10rsso9f5XrS8BhTLRAJjdyhiSnwOjNXVv12wK3jZ46lN0LcEER
0Tgjt9RjumJzexYZBkbx3jnZPa/67juij9sx16Nwq58st2UuCxtP/InhFRJnbPP9DRZSZxYX+H00
X2t0Ha22NtLhEekIQkgmsA502U2TKo7SdWA1hFZhochyRbLT893W5wDQBJwDUdvg+9D40koAGCDn
+aebJXADhvNkoEyawRj4IDC9f/TTXFz8T6TPPt8mwiuxivzqqmnU+wH7EuGG8Nj+XJ661qG77nq2
F36pdiNeKN8//uwZQo2tPe7PefzbY4YqTEYe8hY87nl7Q0NabfLJ7T8Ua3zwU3VojXPS53FpAiPX
6jjwujf0s9a9RIErW3sh8iEg1lrlK0n7akBNknbVdoRe6+FZ67Tx/3kC1VI9i4u6Q+tt6lXqQUoD
mugrSNPgNp0Y3ZhCUkX6PruSqsYuaS/1LI3SLe9f5RyvjJ36H1DjxRtnCC+kRAXuNLOKpvvbO7TQ
MHkQLm/xw4+9Jf7MWPoUyUBD7b6/1Z2mWi+e29zy3HWoUsvaxhD4dKtsQpomkbsXP+yCeNPL9DJc
DFcQpouvw/z7fa+KPDlI9wltcHRVB0CTCMN0H69BMxwzvE2bsfEWpUsmDlJeeD7oy9W1lV6ss6ar
p0Lkww/UfgCzrj/jw4rmn/sZXp6mWB+gSzps+XMTjjNhBJqBdGTQsyqwxuJ0Q0B5HKUu1if8w7Gf
woqxtkuJbGvkm3tszKGD6QBmdd4NmmxaKdNIO1a9YRYZO03mRgolYZoqS6ttMxUFtR4uYXVSZzo9
oW21LEBpFZahG+UZP7lpD8ziR3HtDe3ozD2rxFY+1yqD7o9hnRTZuDOjyJAYgC7XGjNld+ZiHMti
39ezf39/yvWuTVyLCA9e/IYFz8St0+OPTcWfpTgTk943R+KP/Ytj0ICsVMEWNMGpoTdArNM+q+Y2
yfLFS+zhWq4eS+ok9feJ8R0lY3AM+Xlr/diPb8hnHqn2Z3JQVLwx6R4r0jZV3fDjRHn5x6YUe6/q
eM+Cfzd0EqMB6HsNMCdUSHq22qp7xqYZ3Vh01GhQ38Rx/bR4bg+Cl3NlMJ4pdkwOo+pc0v0f35x1
gbJhVzcXsMjH55zfl3HawOxCHi2dfLSzfh1McfU2unn+Lfhne/wNFaWEX5myu0q5fC4xUbFL4Auj
wV1xMieIwH5VIOmakadwxutmL/ffc+bHEWaZymc6ucjd9mYgKubqUtBjb5bTDJaqDP4OYY52sH3A
DnraeVwjm2Ngr5iQ2RFIOHGO/+k/3KwWFIjpGJgNO8lV1aHYMiGFsDcMN4amK6+0aiiBahqoMfe1
kmU+gSkqp9LhNcXM3J+Z/DTIhUS5cxuM7Fl9d4BESQCT63dTyAgwieDf6erpsgcRKwWDXA+UhnP0
kjhtklvnWYZEVSXIbEDURGQeu1mokmsdJAUYuGCL07odvArk9y9+E1EhBk9hYZs7Hadw4qR662Ua
EVEt1ncA4LFvsXg4AFzC3FhuC8zmH3E4B2WYaHf5N45lYmRx7/gBoONg4PNB2LRDdu/BJX6f/WQU
EbmwCGAy8F/E6AMzR5l/RUToB0fnZenBhl2rh+WE4ocCaPozlj/XfZdomIDMz9CTlUFPijnpHuct
wvjqFt43/p0Cua0WXf+fg+pLW21AO0gws0Qgsatb1A7ZIoi89F+/jisRuFKy4AVcwpFLqGgp6JDm
1uEQeGzvSVAKOLxB5AoJQcfaJK6MWY1IIoaPyCE0wHiXTOPvs44uwzvY2V2Gdik4SQo76AE2v34v
fflaGj79qDW2Rvh97vMK+j0rMsX/pZZg6/y9dh68dmDKvTtONxYBkWjEf08T6kCDe5xJ31FU2v+R
CZJYRZTmjEqaNHAmc81Oa51ZDwyQuLjHsB/B6RlBoGbvww2U/XojTQWLxw81cjIvla8AhQRal6vQ
O0+e08hIlRpD5UMEXBmMlZ5BuzeVKjyFvIGucoogkyp9NXJB+b0TTxEktAInLkJr2PPBlrHpxQI9
4n+ULnlGbMsaMMlz/gKDh8+5Mxp6mTtAyKzrVGbi4A2BGmw+c1wL2GBHmZ12ZCqvf8p+epITaO/s
GO0L2mq1eeGpwU9F/hJ7/SOj2ln7sqo+THxmIW6gXWdyLugOCqSE9pxFuf8FNQx7H1E1HbNwwrwZ
GSavc5iZABdS0KkRXkcdSjapgUPfrkU1M3g1Pt/V7Zh9PK+rhb9SGh0/VJkSB0G8BgCQfmli/3Z0
95iNrl0axk7k5NNXqxdVYXbmCZu5P7lP4+eIKKn6Pa/ff40qXXfKsztnSembEQHLydWclbdKUtaC
ZhBoH3v6GVaNcRtQ7OuSsAmr2s29VGVXuHVqOBU9/xbHtsN9upAaozpmbXT8wZPEDSdDnQT8aTj+
G6Egd3WnjBmce0z2SbIxWRyCbrV2dzXDBXdj8DvvsgvlqxGvVHFKUvXR67fPD+uwxiyJlVoMUwhV
1kPXcyJKl6GkQ7eajFGdSP3cM6xwxCaLkFT2ZMAkM7ArQ67dV5ocCWrS4sHqu0GasbOrEUDPmYmP
Zxb7Irka7H9zJqx+3IuAUefCx56Zg7ko+oOYqM38Io72VTbXiUu9/fbGeb0SbsQcixXvanTSmWDn
qEzxn4AXOl/XAsQZn2RhOXBV+S85HnsBL/BzpAy5v+uphe1Uerzz+h0bB40bkisLjh9feGA/cc/R
UxwzkYmzpM+7qY0X95VqWInNQ0OPqkrAkOygNU1Nl2JoOI6iUW01QjlxuhoPEG0Pj0qyAXBpjY9y
0+20nW6L+86qMhVZe8H0abYMFprQqOaU+Nhgt1CFRPDSvwa9EZo57WGoiH0n+gSYdA4fAFt9beVh
L3NWJokP7+dE4NHn6PBPLryMFwnHLGoS1VFQ+SOwFTlUeX5d21fTYBPRR8hXfGAkwqpVD7TY19e/
a4ZQEayNlR+eN3Mgkm7C/6vCqnTPlCxP/RzdLl8OaiLZm/Jk4Gb+9KQ+zq9Q/5nzlw/sJkBMehgj
J79ZACPRp283jOVep/tMt0/It0i7ygO6G1ItGPrBqehfNO91DficvAHcu+pAKNDRTqaJWnsGpquH
pD4gMvWOFeWL+zsKOdYv9K0QkpBOBoz+5QnLMlN9v/soR0M9aRZyoPo7+eNDEhgPHc0PJ0gAKo77
VHCLtJ+xcpz2M5dd3bQ5at+Pu8tptYOZEi2ct03F+tXoW8gSfbmFNs+oY0KNbcaZS+TV2ifkq4f8
bo4AIRQEaO0COXwQSRarrQM0N0Dmnjn3CnPr7CmlpCzFPbHPLogt2iqTAVN7gzVUCdVu99f0seWC
OkWA5mFSgecTKYbqFpLc0LevJyPIf9PTrs6qE5Vvw2QbpP3T5rIjGBqJ63pr2OonK1gphG8lzoBR
fc3NX1x4a+CvYEH/5T7C/H2t8ax1Rrp7qCbHU6l+TODR6aDKbHScYyM6iXzND13K46QgIMQLWIt8
BfkkKYeDtuMMh3jW9TK32POmnS3GxO3ZKaI16elfQ3m2aImfFzisVnTFQWM7PyPEkTb87LblvQNB
Azoy+vvBBMIjiOmL/bAjuWnUzP5JkjW0NqZV36Hc+gUvwHdJj/dJHir6KQUjuXx/0/EI/ksbFpH5
7cY0DDjjOriO3Pk8IMwjk6JnDSQr2HmgWfsvCqp/SeCVEqYEVgrVb85r4uxravoYxBK+TdXoDJHZ
VipBMg2CszhiOjMdwqS374fQfmCjZWf+kzV9n7PmkvSV83fGOLTFIJrz9CAatRXmNsmRTMyRrfFp
g7PbkwFM51L/SYd9603BMm3xKMwPqntVvdn2t/nvMmvRqrqugySBn+34yCqbZjYo9VsUfH9RPmXF
Rst7TIpsWcLRNFgHY5Xch3NQgj64d3TWe0u2i0A+1K4e9+pNBH3sK/bJb9BBBSzg2znFfnUWBSW7
je4a+x4ytWFx/kehu4H2JGHRMN4H0+iq0Wk5Avsnz5y5btlkts/jjF0d9UA/F+gEz9oceAHIH9Ap
mIlZsVgcDpsnVibeQItaViOrXsW7YPmR7swWDRBP7NImK/aLDvc6rrGlw/B9kUYhwXFhqT32ia9e
g53XPuXlq7fpyhAzJTv33IMEH5Jjb2Q44GF3+o5ngQtsfFpDy8ji2SeYFmERz9Ad0MPF5xMWFIFT
oqlOWezLyjHK9xVjKyPCrcHaQh1FRbidFB3eNa0W1lCLsPneXhef57xPaNEhKWcInmtPOt6loF9g
VgnBDYJmBSeH8G0pGTzRG0Iq8CfdQRfFDDmddsOvG/JYbmb5NN53b0kU3rIxIjtQI8CgBmTYgpUZ
5+C/SYvGf5kEcjWLJy/HmfZnm0SrihlOn4Wl2yF2tQu3s0SkPRixFUxrfJ1VKmQLNNLz9uqyRD9s
swi8m6Gr4fWaOtA8Iz53naTFNh3jEj/E5mVR+C/UaV81AdbZlZRlJEzb0B54YtbXfCzdp0c4cWxi
5hFyTnJqovh3ea/2v+QVNrHMsC2Xzt2Xc6ef01yG84tY6GtNOG5LZ89nUtWnoe7cBbq4VnwmVxnk
6HLajKezviiHvLQU9UcjiVCgT+0HNKv3EVbylvzxQ/I63DEZBQytddLB+BHnjBpBLUvtNJo4GYPN
UPAx1IUV9rifiBz2D9zodsdo3NLwaw3VYcmRVzJGCJqUfW3ctksu/9EXLLqpbzf4Coq9DJpeRa52
wGrNGbf0LQK4nFlW+UEzqHfevNf0lqvifIK3w/A7d/w+EShSi6nR3OzFrVVKn2TkOeWmtAqdHhJt
jvCCQmZCf4ihPz6Gt0OADPFxaDqmElGGIIAwL1cHRL9FA80f2UdH9txz6epAvwJke5CNlSgIak00
ThFnppV+t/W9SaRDsjcwzwPCy/15Ss8T7AwumzD0feB5SjNkPGU6JFr8ncnQmOhXh7cXc1ha7NuP
1LtvsC0fnN3f6DwZZ4SNhMSFO3bsh0immE60jXgif4TSKjvYhPS29fBDi6u2CozvQJDj7vs1d61I
fioEHhiyTuGiZKtds3ish5scpuyfJcUxOcKJhrj7lhCNwQG22FQI0sa1prtNHptt3skav+XIJ1x3
jkQLeEXs+EQx4bYna1mTWiYHtZDswvKYFDsPI7cMCMFbj+AKogVcys9TmAg/kpgS9LbJqeMg9cHa
CRWbLood7xLL9rLVUZhHoEHpk53l0Z+HzEO64ZWFiO5Ye4SVRdcGd5B8NSnf/do+2+VXZ8nbmeF4
fky+7jeIUtKcRWVDSsD1/oxXIDzMUt5NJpesutuFwF5u+4o9koCfw3zJ2NqGi67NmwtHHnhp4ewz
5pBc0bspV7x1tzJPi45ZOIDdXayVoyW3SQMOwBwL6r9F4Sn8Gq2mNjm+QU0LZtWRp+fqfKOXZRdJ
vZ7hplVCvXAxHMKNH/kUcffLGqckyINC+PIqZWwo8+imG+81o7NIK9YnCLCPAI/9gRb7t9emW/hd
bxH6Gi/MS+U6yjYJqEojsIvFjkijgOkY4t8UbfrYVYM6UUAajGVHBEBlAneU1udILkpkc3zOzdPg
+SKJT24VvvWUpDgn+G2Wrz+/nYs19IKtP0VqF0XOMOVyF/pq8T7E/cyu/OjQ7zRu/qTjcmveEQgz
l9srnZIOQaSQEb7lIJe45/aMwt8qaHIqa0iTEJ5xpULMg/fJDzak3qiPEynCEaVsIXCHx4Uhqm5g
ON6NL/JXNDyhmQtWLOSEucf12Pn22xzRRFAKR0AFJ+35olKoWVeWU6d6sshYqv4jtAlE7S7OaQS7
xu2yU5uGDgvuEb/RV0MqOhYrKFORzGnr2v7xR6QgkTOMgn98fGDmkon5uwOTCn8E5nBw6papACSI
p0xU5cwCPPWGnBTFs5e68qs/zZiRYM+l06Won2nof0hRQcR4tAvNcel4rhbewiZghIE//lzK7GyF
2XAvsTqWmkstpnzvAK+86rAK1I22vFSKEyJzzcI+LG+URs9WSdjVszlgJ5gUSbgHF9g0typWi+GZ
7q6kltU9Zy008UjwQONcwMJ4iZ392CO/aeX9p540S1SK7VzIKmLkVj/t1FMkUwXkoVO6I9OcsX9Y
PQYKIEJAKMqonB4ZjjULVcRqmCybYVGVJAmsfMo1LqFwxCZQKdcj0x0I9hRkMg93lO6XWvO/SKgh
oAkO6rnenGQfCFRbjmWARlQwpH4NN+f59q6VLnvof/Qr+oerL1+5WGd09EdVPl/73nIkpMQIklVu
BKWLrgmGdYQ93+8Db90UrSTbNPl3+e4+bul6HP2QyXkUM4IhzD6l8ceTJBf+qvy13e1QyJWNopw4
16E0fuLB8oIkU32npYYE7ds+m6AL6UCv7+SZXZLzcxoeWVrvhcJsIUhHi6Rol5yQJLf52jiXNPa3
h87maS+3rrD8eijGr05Iu0F/AnTTiaRN9GbLHj+hrwr1z4mBAENQOR8rUTi8g9J83uTLaOM8yPLv
lOwkVyJpGt7nW4oO6mXbTsgvDn4ijzVDG07xl+m/B+5yotPBhksSvaIpEQwQNXFvRx42GcztOzct
d2KAYfs1jkTfJIYETzhW12WaFKmXamDUIUwv5Kz5buxIyL6Aq7jx+eNCE6drhJi4P/KSE4tjCUJL
RWL00ZQNdnCS42dA5tx+RqH2cET0Ud8fgdpPuv/C7nkpKcZxiX3FtWgLzxiZzJgEZ65AGL2DURvc
6+8YzJZWgai8aY3/1QM4tH9RLk5KELmLqdxGO7ULedoTLDdNVKy7f0u6hGon/FP2DF1lJd5A/2Id
QAEyCkjnTzYjJavnlP/UwmPnU8bXN2v8NvnlSTB98bIFxBoqn67MsQZYYOUlNMMfM1YfNXmeMWrH
36JJM/MKYK3UBvGwU/Lphr+dY6j1e6Ib7RLJDnsJW/Kl/F0dnxK5ST7AUROUAgC4LJ4ia55kxfDC
RmHqpqeOJJeISsOj5mUwhF9QS91EayTFfQHvGpy04OAh8h5FcOE48gAHXGf7lKYIrwHrlAtPW24c
2PdijR/KAPhy0hSpbjOYOvK3ZAOpPpNLZP77nRUTzimhq+l+iHlIm7DYzX+fMnhHahx7fGt5Pvs0
0B4Kc1PnE96aWs45bvglIohU+/HFZJZw7BMmD/fqn8M74T6DVXCgmu29oqzSR9IEgyWFZ5it61j7
9jhOqweVueFSRZKCWADm/wfMuK2mEimjAiq1+2pwIgIdfpE5SB7BCYK75StK48kaL/uzlED3mXjS
uQyyQWsx/4KZDg7mBW1Muaoa+mpyb0rucy/P3qz6U2vd7bQWm1p42hW4ifdxwAGUJxqHCbVk2Cpo
kZbyf6IGT7GfCgLJRCsG5r1YgvdsJi4c+o8DF6iyDsaikKg/baJ3oZnkrwDcJVqruh7SWBH5xyau
UPbQK26muYneOVEnGGOiHk46jg3FoNylYcnr0z6J1V8ODXkqhgMx3cKACLarC0fKic6UaLRwavzr
vgqrILr0jpGiuZMB1j4PftF/g9EQHbMeHrJtyrQcQqZ9SECsgDvIFzkhA7wqKZYb17K1vbCK/ovy
LDWoa4Tue5lNs0NFIZ5XEYhq540B+vIyTJQhbADvWQ0f6XGunHpD/Y5oNT67D8OSG6qG6nRQy5p4
lPf+eVvXH1EP2x+awxNbg/WbDW4cNu+/wJEqmXB+rwsCnbaI8jlpF5fFqgdb19ccI7ImB6+Odvdm
uSZlGL+XkTB25Eez2HKta1e4eitG/Dxy/X2OkFTHv0iA48gOLI9tskLjKTbAZwJ/3PzgaezT532l
zmkXQJGE9qCdgbAYD+5Hk7/DE79ZKiPSDxwNFOvu3BN5KYmiU1aMouuTJf2LGMhjc04Ho3S75jCl
g6Sh+g7haYf/OYHURBYaDNTErwbaiUYd/TCqUwS3wPii6/Vxs/mAJYqFf5cIeP+4+8AEI2gYAhlc
iiF5sodkd91PotcLQzABoJb0eNNW0ud+USMbPyRbLueOwxc1QBCcnVyOQxySm4w5lRXvC0S/tVHd
dIeLqQXHjC7uRI2wnaWjxu5QTjgK1UbM6zDbkwu5wIRaawZF3IX+XYqT29JJETkqT+kUzbGLYCte
bi1VnPjJryUfTd1/wdwqb9RlM/euh7S8dZPZ0K58CsmOkJCgAfgVWsyHKWCll0Z0g2ZWZi8x4WAG
nl0ZIa3BPX7kdDYWJj4AimhmFGy+MCJ1SgxswoaJf08JjcNX/yfVYn5X73CcLNWiDmEl5IKY7Zfn
/moHmsiKM/oHkjdDbrWgspzWx7bBCnWhqtQBkeEYobr/GnJsupL25Dj8jn/dmtNG1QAXOch+drgi
R0lvp9Ic5QBF9vgcPtEZuzk2u0TlYsqfzUFIkrWz0HGPNlXa8xlUmAUFbEuS39L+O8aCX5WoHSFs
2o+KoSxCVKyaHmb/+vbOnTM//8vxrBVdBxbbdUtCTph41UL+h2cyid3lygsXygo14Y+NfXSdUhXf
a0FL4M8DYPx8pEHK5KUk71zEAXZmVgvoJR46A7+NU0VjgiL4AQmCHN7ScKTTeycag3bpY06ZAZJI
sKlTbD+YQvjyotHQnBTcItk28+77Jeq/R9YAQ1j5Pdj7QShtx2NHgfqzNQL6phxM8dWcruXzrXD2
VPtCFua+IwTbGR37uoCHo4UM1LU7KqyLkXFvoWyJw6maABUeRc1hn2n+E2XLAot5EmWCL2J+6XAf
zQam1Lcozl8hf+wZOi1MjVVJOVMHnhoFOS5vay52yHalVHG+3ySzAhH0uDUHOJYJreTcWpOA/t5d
YkBRGyfgeSshNHdt8/mNlJcnxnS874o40j/eEE3RqJbkAunRaIGuC5jfEgMw+NVArAYyq8tCIJkU
ElscugYqFgTj9R6bO+DeYm1dCxZopci0K0WcvZO1lm4Usj4FHJ3ts7zmsP+ErDGBNjuD4RwOZGLs
egLTaiQb6x+7ugejbxS2SDKmn/Ft0LLgYEvqq3owWOAXDHmAop6oRnGXj1GWCZ6grTs4znhdEbpk
rp3ST2448NE+FPSwPc3kCh2f8tWxy4Z4fX04FY1WSyzJCiFAQGOpPFm7MKvEvQyuzgor3VUVVbAE
j/DBONKmKA/L3DK476Q1R+DjZbX/0QebEMLEER/M/78xxKdhN16cP/8AV8y+EZVf+PKgar9I2Hre
oKp3VBydVR1iS9+jyMhMb3rh/GFQNuoxmrOVbLIZth13KhPM8AFa+OSqOO18svMCk5XaS2kpOJaJ
SNyIUTBPLwjrKywoyLFIbqgAfyZWGMuUJZRdn6BmgRdecWQhY9LhAdJhHTGAEjiXdgLILb2LjSJM
Srtl6PjVv+HBbwHzEUgQZBizp6DGnct2s76Khv88OYUDEovQQfllOiBk0QwHo+w0TIievHcTFZM6
v5QQ3OxPLHB1Y47PxDDKirl4O4lsOQRVP5Dbfi7dzG16jwgFeHL6F+HZMgk80vm7aTFvPlqL8lMc
eUHmjDlC6WDz+1iiRnFnnPAsD8zSj+3vDq5exN+iqi+S2qsnLgkmeD+ShU3/v/1ZPnyt4489+ZV3
ndOA3X5QvBjSKQQ0Ct8WJi1OTZJ3badKkXPki/utFTosjOcK2zXx9rp76DIlecrrQqI2ezv1et0O
6hFAxFKeGsrwIALAPwEtEln62CNzGdmuhFfkJNjs7pNCrbmoqr/6HfuJCu8x+4YnFc4ChWp4YlIW
REtwfMTxTxKiMdT9v3wY6QChcy5z+lN7vI3JWkgmcOOGNrtr6r9pgNptpCdarMKplhk0u0T3FWl1
HTBw2BZXyv3IQgpyLDN/wWtVd+1oBsSVe/gJh8b0UMzHVJ3ho8/Qcrv5BDtiDm1J5nsoISYGcfGd
s8yp95Pp+7vZfpZ07pEFtHkrHCySaYOqCOBkd7hm0yxsFNbpuiH+LmZdcGNFjifCuWzdEGR5wZU4
Z5ZBUUdn4g+Deagy+uRHLM01F8TFHTYlih5i4AIr9Q21qGtrqtnynqoWDBkfdoNxWIiQ/M9H+Lsi
AQ7dbIjdAi5FM8r3Uk/hYrE8MgTgK9evAubqSxw1LCS48/cs9QWm9+yI+VlqB750n0Ywuza1WhOP
yuIDB9P7zGUviPKkpYM0/6cAq0w+Oldz+7NgBQS6O6lchk8+v0CFv6uzI3NIu2uIcKPnJdR5F83H
mmGTqOWOxz1iIE7ZAmnzgd9zvjJl2xjOBVmP+/lzg+3aZGsvDJ4GjhYxZO2HGmzN0+2Mr4kpGq2E
VnM3jJr28JszhfAwkTtDqYGBxT0JJbh7Oz018zQfN2NVw+6VsnNKR9hn4zXhphUad1js7ktGiCL3
KnKmSjO/4Iww2OZ5EIEvB1YjvYpe2LQaceXAEMlDh1va9eE5oMbX6mgxz1VnhZHPEZW8L7EriPqv
o7Bm0sRy2hUDw5WEvPK66w+DEWzY3qlv9jsBLy1fyPmaa530SYugcD4ztSnGwFBNv+lglDFXH14k
iAYcpCk4LLWnfEeyzbBw07vQH0mSNkBPotwvn8fMuy78clehU3lQCuNvBIpNW80Dw9RpEjS2QG5v
/8dJIYg6hmnIGjd1mbkCIFcC6TDF03MOvmem98VHDijzhu4EbSYCOAX5f5QfzI9USB5dZYCEvRBZ
u2Jk88lfLOEJgsRz/zXcope0uUIIyd66Pyv99+aBE36PsA9/2BpPCx6F9Awg1H8+u74mJ1bMovyG
Gt+yb7EYN8hmthWJy+njESiOFgRLDfaN6RZ+wmbDY5eu7NlhPMPt7RifY+fXs3iGjcAA9X8rYuhj
DXPX+lqb0QaMaQduyc/4ekr/CrhNhOPrQRygx1tw2djFPu1jYMbYCGF/B/OgkiVL+sP5KlqeTbvj
CdHe+gr3YhRnwOhJu9gsQr/XWbPgzuMI9nOILBR4hi3gnq5J4eTdTqX4nCJ1/ZNIyIYTBSUp+7UP
NnoqUR01JO0xkSDIB0lVdk5A8rUGv4BlWIeDSMEF7XaBXmf8YAcYtD/QKXlfa7uyefOQpioawuv4
DU7aLEGlNOWzeYoQ90RcIRBx7y5OQ31hzRm4hFWqMXsEAS/n7NLiId7d8r0ni1qBs3JUcWH5OUFB
hsKg9CD6v/0nAM7Clf6X0MdDWqkmoB9AyqZs4edbFmPt7gf7pgGquda/4rEKNRdgl73wF3XPLHw/
rke3DEc9Q3u5vOSaqcGh4xevGwASAoILVNhZCGwejp1hRizWbOhG2yvq4qGYThpm/uOIVukQHsPR
k8aFyu7+tBsPlb8+ye6EFgPNRSo3sX/7/OqvnFZ+ek+T83WKQAGjcBhhST2nEJEi2xjjb+PvigMi
JLQsWsOKN6PWT8x8oR4c4WHSW/9roYjnkgENbxUJHevowvdoA5i2ixaP/aVTckzejUfBCukdLvD2
FCVmCu9q+EJSIL2pIvkSJIGOLn6tsx/cbqLDcNt3lQdLBybWyMEldnPUwdEYGUojM5PKngX2FMJC
ofmphNRJp6PFz9QDG9Nl8GQ1oHyDlxQpbwnImP6EsMRVuEfxh67BR7YvVxPCTShph1OVOFRHOch3
+Ziqrrw95QoS4vaci1FS+X76n2aNqmnm92hAugCFKxnkTTXy1V0Q1uO+JbOnVN/YLgEjMdjDzoW3
Gd7ULrtcU6HHEZo62EWVbRk19ji+akr1JmUNl8FbVNUnsQ2L/pVC+ETy0umEnSHRqR7fTezQNNIC
SWF8UyLHs4Hux3dUuJcHCvrulHr3cG+C0nR/oLsowXpiT6fHeY/7hCgq8JR1IAfaXQkqBHBJ53Rv
6lo2XEOIVqMe1vMd0iYgUWon99X+oPP2lgClJcKtrAmsVHDHPKB+ch5PifECLxAF1jCri3U86eif
0TjP7ByYJ6G+iz2xfthYNfnAVEend4rc4J10jXW7A2iXbBTIYOmNlfdBio6WnoRqMlP0FDKPyBcD
M5AZy0E7Pd50X2j+xhi+dvMnJt116K8q3u+bne5vLUH0+EDA5oIT42wNYYLDcTHRBmDw7PtV8Vzx
6pij18+rG9GsvsD3thfHmEkLkg7S4zyX3hRRc0ahTGQx4S/K5b39z62+QWX3F9v+Xsi4i6P1s1Z7
OyeuFL6P0Y+vOBEhqsFPGrTdtnbUB4EVoHn80ztQZTs+JPcqxjRhaAFxRYTZPtwO703kvDrseQME
vfEx45siIiWXj9KIFO/f4BaV3CodqR5cwRG/TF39I21LsDj4wRhzs2Di0vmDaGIkOWZuy6VVjBRa
Lxifbe3SJtYdfvYBuJK0VQsLSlKbFSdCwfCMIsNneQVEnofy791AAigqGzBPnUtZJgV9e6J7tMKs
+r0Ui3BVs2kfl/S/e/qOt4Z1EqI8u7lLTfUa2rUA7FVsJV+H0Oz+yRRTgaJpVYBuvY3i5r91LYTy
9VW339A9wbqPsyTGKS8xPDuzb3i08HTJdUBdBaiLeFbU7lpmkdOPIe8uY+/Tl1MrQLchAWGsGvvv
hChsRHcY4M8omRyli8gloBv9DtWUqwiU4ZauH2CCOUMO/8qnr5AY7/eSzwNow9MGRsMzG3n+wMwv
242Udt0JKHrlU7llTd0NExnn2KeZ+jkZwzBJUR/2z/ghLntV54wpYHEKfXTsnsk9HVkFr93goL43
CHbuqJHaSUTWkCvzhjQPkfEvq9BsBxLM6AoPskAqPcepBP6/1mvGSbHw9zEwdr8KlviA4Wvcx54J
n5VCiAMDM18Gv4pR/CcfT5v6sgdUGqlmJZLs5/iqwsoufSsCnFWkPGkKcfwO8wTy2kAUG6xxHPPY
aS/X9hm/NECYQRmt89BlrKrYRwa06imE54Ib7hNKI7p8KUAbAxJbKrzSntMRZSBK9t4DVrb43ozo
NxmaRu8pFY+cyKeRaaY9lyJ9lJDDJh+ik0jBXs8U5qfLYLtaC/XHCB0lA08fotKj2GjI+SgXATOc
9VwEswESQhTKUl8LZVT6aBaRPNCovlFoMuuLLV5BQGwAnoVu7UXyih8vkrRNt0eo1HJyBX05lmC+
De2lUimjghfjEjLNQ6N32/znOhavED5hC7uDhr2jwc5MWSfLmAHXcrKGEEIon4w4QicQ6FQ8fI24
54lPpLssrSUwOoKUl0d4ZFIevP/qByvM/x7+Dcd/Vu3B0ZEolVOrcJye5WNyBACWKLMrLISQdCqT
4i8opa8A7scQUCQyIVqh6oOl06serz52b9qwuUjfKCIuDTEuJtwBozVqdYtTKSu/q8Mp9n6h0QcC
iPbFy0+KtbsaBz0r54aEjO6kPj++CzGtq2tm1dzYWdxoZtjBCaCfp8+VmuNlbjFTQdNrj6JgOj9A
+JmOHbscBh8pEs5EU4ti+Pam0ni00OLg8O2CgSIAqNbynMCJ0ttCyJ5GU5wPHEbKNDrDmAh3SOW3
HOaXKQiusJY8LA4LGSrRtNhcONvDUW3suIJ7JSwHzTT0LmOMLPFO/6IskdMkYKCB2SEm/RClxKOB
elWT2KFdcb6ANOapWMJqfxrs7YAQlpQlWO4ngu+WEu7LHW3REGjQGudkqbP25bCBAyzh9xMdBDwx
BsVyNjZN9oDC1uvx7K0CpsGvsq44geOKvfLmxuFooIZVCJTaSy/R6BgBc5PqjQGJGes2Lqwb/FxI
MQm4l/ZZcNRwTIjUwiQ9TSyHNEQq0X3M0ogNF299Ni4hDJFiCB4ahb84QOmwwmJQ8d4PRnuvgMwM
0Y2JugE8nOc64nIuA7JOlZCBuWljuCUVg7Yf89+EU7ZRF5D3GcYCYmFcPmII87yjsh6IHaH8ynDt
gDm+/yqEWRdMoIXHmZRbif/0YgqbhGUESvYCqIpW2Pgez9zNqrz473KvjvDGH3sDcHzunqwFmaSw
Olggsuy0+CaU12/n7F9bwQkkxE3JySN9BlA9N3iQfpA2uuSZheUmG858oSrPkIcoEajsMaSqVVVV
HCvMjmWGimnRkCggikTC2iSyIXBvtmaILIgVlxT8Fdp/W9S+pM0bcD7OM1D0R75Y3uNmMoPJyML+
3WjED1EP9lYCZZ8KjI7tOOXi8h6rQZEVTD7oid2xnJTLl4xKSew13nnjjddfJO7oePctfPjPdnE0
gVS4tprbemBaEB+6P4Y1LWIhkYM79KjFHYLBP652yKEMy6OtDt1HkoBB2aswC20LlAGW7CM4BSPo
njxkFeqGrzRE0MHBLnHrs0O1CCA5Ci3OET/pVXs4nCoubhqCuXTVPXWdSm8HkoQSHMCSz1AHS3rd
iOBwqJyLGb125EHygr5SlPSuj8nspreVmoslL/WPIPmF8z6rrmuakSiuv8ikdg3eQGZBN3le9nyq
ilrYD6wWeotevhfGetbEzfp+begME4XRLOSZ+tG62r2MuK5fY0t+NX8KuOh3Vpf8m1LuRZ4own0V
2pbJYqJVYwfwiyqC3pO2+B0JJoRche0O4Tm/n9KewUdNhPz43jAvAy7qCt0UhVbuOOPj++rIGR57
QemOsMR1hvUsGCcO+0t1WqJob9RR8HXdllNVAuX0b7K+VnVmD9C5KZuxw+RI/34gK1VPxFc4XwgW
uvtC70+K4ptqIIehUYJ/S2zq5mBH1acSbOxW7bHLy46tNVr37TjZU2cKqjoCNKh7Atx0z0AC1xEW
/LE5dfDXvC+igaWVOzW/Z6uDUfNMsW0/czlaTb9ieP25slRU8paerCQpgTgkNsk9QSPWaQme14y/
QgJdOMt84qdp7VhLbSAWyoiWhSXytqohk6FXiwRSqeh/Iyi1N5o2KxhhPDBBYzGr+RVo/2qJb+Tb
uRN4Py1RMDCujf3qhlCAWjZrCl83vOIIAmsvWBOf/pNVwwVW0Zn9q6dX96t19uwG6kY+F+lyH8hT
+QZUhEZxzFkmTVssQ6AdHWHP0eb4Q4rjZB3Sp7idHXi6sgl/aWqJSftUI35s7c4zGC+aEIJPBY+z
je6xurp+RLer7RyoYqz6NdTs7bDnvVu08klm1LgisMdJ0HxZTwKzxAd8NS7Aa3wgmGsIRZ9tGgSr
V1tsQFSrm9HEYZeP9BYZj1T+PHwwKIxePNMFCOEm4kNQQaIl/0yfTTvXiUAK6JWJ26XyYqA0uEJf
v42kbMvqfIBDVGSvK4ftGJBnqoYCYQLEmuqihuRZ2uNZH3NA83APhvBzlCo2pQitO+6VIVquA3IF
e3xkeyZcKWjhkTE+s8EHDwgPphdAgS6DLBpMOLZHD8h5esjBO1HxHPVJgvEvaEJOgsVfkxgKC52d
7zeH+XM6liMxXCKIKAqHJN6FNQyzJkNJJzkuTu/xV+w9a1Q01sEjsoi2kyl5HiCExCi072gsO0El
yvRHQKzE5pOCI19H8MLIc9DoZSAH9grpLEO+gqKymchLgOeBY/7kB17+156TUhEKpvln9uDNOusx
yxACxfFj5wNrI76A4yJwjsEyg/k8uzLtdVdW0RZoWXZ9L7PkCjxvSpw7UgA1UQiDDuLiz5tLpRGB
LxO07XYYkBfdGsKtIrhgW2kCdg4cFLPetGgedkp9xDLysZAZqYk2Djz6vwH90dvPLiEYP7DmIilQ
bJIFDkucCpBtU6XHHlPpNf0PXJXvqQNSWdeMzpEtJdun+qkqhw+g1kxeWRntz3CyKbuWCbMhYUmw
jzxl4tPZbdviLnHVH2Yqz1/nxc673Vy6fmSm4xfvVH7ycTuZx9/Qrx4aAkREcCpUn9m/yUqksjSf
NN+ZpbQnqFL8agAWjUVT88r3VHfI8790D0VYyWZgFapXpGycSldROqKEq68Kz9AUPXLIcmxAMhB3
vNbKAL7SbfMlGs50jcZ0OAdNXQGxyz6kA6GRiK78ReYmRX82y5iNkQCygnN1Zd8LODhl9zSOyJUj
6b6dS0V9d18NNLLk08aOraaA5Ccmmhm773dgWU9PrONb6bOTbFDU01tq2C99f66yoacQIYnC3/KM
PcCk6elD1qSgQ7pdwUoJ4P7qp4CQqm9uJEBhYvKTi8N8bFHc9UA1JJj+enEBJk31BcQZzO8krn8t
QHyDCzA6H06om8YXEKzURVJmd1Q8fg/IKXQU7zvYVgK0BFPePiVLD7QPIcHRl9oBeu48yDDl2N2+
+WvNdVyaPNlKqPWTzCWmh0MfxBEL4zQvdZybXG7EhwcyDIu+HvPUjGmgNK+TSfLWsgfZa1+4JVdI
BDEpNQnrZs3oiw0y86CnGPG1fI3JE+LC1dRjk7oV42LhQLwrmESFvIBv4BlxXM56iHaRVuFZVJ5Y
IOH1sisxtjcirJ4iEtyeDGYes06zow88EBWB2Ha00qUw67ILuo2rA7iQcxvUvJftp2QrkTReNFiy
9dKV9dFQBfz/LdiCqhwGWBQTVfwOUNlM9+TZEUC3SwI2jtZUj4gnKsxEZHSo8RzXym5QAe3RMP5H
5oAqu2yM4SvcCWgrL+Kbg0GJuz5jAWd1XJzcgYpu9QQMfIQjvxjZzLIaBKFOUZHOQTuaVWBC5PV3
7L1o4KfL2CJXrhiSZjJPSBkJg5PARyvzrDbq6CYShUKmD/GOvHn9UI7r55CcENkH/5i7vyyuCFFc
gl9kKghsqtyZdA2O20q9IKOAtFypbjGsNizDhkXVUKOZiDCD2g9WT9CHSrgUKSIHXlcrBcFuXC16
zohU+okE7IH/neYt4S/GXyAniVcfLaIywojXvaIWLGgIdJEVztdwJfNaR1DmgozSUfF+kixtG4yn
+cRzikz+/Z2mTIALzCu3TF4+DgLXyXLutF1aEYgWpraOZl325JSD5nlakTfg1iMvt0ziG/KGwHqn
7dqpMpUClJprEaLEfRX4c//Sj0f8+I+ui7gdQokhkWajbaRc6f+ocmM6vLvvCc/56MSqdpgG95Uw
LTR9iMNLv3UxUzytcGxWL3opKptWlU4uJSZaJqR7ee1JCj2cArEG92w6RDuxrPqYD2lh6KcnaZzc
LtxxdXTAbVzbmzS8y8/AQsq7Sh4dwttWH5D0Ot5op0iZOb2XNkeir5/uI5wjieov1oSoOKqqUDiy
Rk4x33hcoCGZk3tn1flao0Dj0dmQtEFGFwkRg4eaHwvsglPvqUQQ/259ZYlJ9WlyXZ3bNgWLEewR
84tn1WhfPSJTaRJ5/mglUGcnsRWHC0MM2rdcshPsAA9JpY5Mp6iZK5SWT0GwjNykag/LiyZ74Nuh
KKn2/ys7lXuPisxHbUdzF+5dJ+nPNYYdS9AZ9FkQfh/6gdW1NhD81qrMxC1nM2mSaQrtwvR7cE28
SMzNcBK76aC0w5y304mJdBE7lb8oJC0lcaViffhBl2US/vKshX712HDMJvTsTD84bfxxvNI+lm45
0ZtTGVaaIU4hVf3bMtBhMkgy2rxoR7gq31G749ewROLOi6iHyGIwHSsGoeabzk2UEiR1OkcPCQQI
EOiKdqRbJtco8HB5Xhdo6O5+kiF+f2GVcKRMw4OsMmrkGx1KpEduvRFxORxvMScIfq2nlok4n42/
Kwoeuh9ks4amdbSb0cKaGkshBx9AFZFowJkiptSRO3jeqSAWw5ucUHkcbEhA/sck3+apBX5RR9M8
vCvoFxRqLPVRMIm42rekgwAaQd8+6c8MBCNp1E8/GhxtaLacsWPlhfvINXP/sYAbGbN/qsNABysF
ReDzwRzhRLjx8OgzKau0zKIMMIGCmaF1CtxU5hTsWrZME3PJDhrgJG6bHzM0qpwfpUJI6Q8ibEZB
C656ZwK9zG8Ut/P89CAC420OPgTCmk95SK0Y2k6b6XnXXn41uh839crZQtFjABYNL1wRxezl3+0s
YMvRXnHsxbSwJR8OgKS7Hs2GA1D1xX+MvV/PBzvSQ3uV52A+v+W9PZp/v6CpwHDlfRHA4sUSu1rr
yC4BS8I1J3NzHAmCgncfdZCPNmBNRgXBIVyv3OLh+JGACxB9fl978tYw2voIpM9sCU4KcS7ukeZL
irov8s0gekl0oTZqH/RdYPAqF0OeEBY098y+FkYJMa24alghMvUNJ0u+o6QRKHyDE1Z/WV3rMfzy
zRAHeGJoWwnEASssWzYdGao6xbbHHVXheJAzcTOM667Nw0rYAd42qgTAP2zBoolmhbj5ARdUlXwV
bAvG1XUZgIbPWcwF5pAfYy4fCpfhE0bya9z7mkb7w2Z8xfzeM88vPIOg7Wfjj/rSgU16pOXVsNwH
3huGHeWQgpatqGHvd/BVI484ruPHm9zDbJpv6g9sIuumCx4zkNDxeNyS+0EwscTHXLhyiR+YWooQ
wgNOhlGn7uiQs20qcVc7YfNcB1Cv0AZ7fe52mK68kt03SVey11BFOQuG+HLqxXOC6Q9bO0v70mbZ
3VF5GehdNTaUr96eOZ7qkTEeJv9+uu78gGclHpsZ4MJwSAzh1ulpxqdN51I9G7WZo4ExuttDt80D
VyrqfMEC4n+dYTWyOjIptp5UWjmTF05ngMcApYREy7vfoZy413JMbqC4Ocs9BEnBhlgLpZ+gAln/
zD8eE69UNfayuoDpVx6qkpEeJXud2VbDYQBgwX6WyXSbNyxP1BpfkWKukRaDmH2qqeuLl64I4NpB
f5WNMfTDRVEMLg0NBuHfLvQQOM4VzZVjw6b3eYZEdvHvx0bMfsyirURGbCDge2HCea1Cu7q3TLMH
+Av3oE988jU8Vn6SsG9WV9nD7+S3bjVUOJhoPcZwOnplrMmJTAm3pNqU2MgbopwcoSp6A6A4XA2v
Nk9K6PraXrlm3UPeTgEm5t2EXPmFeaUhu2xeJxrovDJtsdC5fEGhQCI1ybsdBd3NRj9vKHKk1ngF
gDcuUbLxf5A9k9SacJ6WK5eeOiuaoCV7loiVYqdEyt0MA/mQCddC8Ka8eYGZvStASludd9J6u14S
0IyA/dFstC14Dgi/HKIVlF16Qpz4b4gYEw3INImh8PiMi4g7uuMQ3TpcTWd2YoIHEPX4B/E/1CNg
CwLfLAHowGEhv3n6RgYWD/ZVgKgBt2+WFZEHFVwGnA4A7KS8dk9kveUTbe5+eJjwM07YtxBmjKdX
m9eo1VTvN5KSyXV/VuQxroPwfrmQqBOSuq4mG+qe9tSzOQ0xSuEiAPxuDeCRq2qVmuepOlLsp/yK
XuuLFyy30RYZf+mauy+C/RoALthYPsDDVWmkrItHLKk2a7cxFmgtcH8fbKw5NoES+/1LdzJmIkui
MZgJ/sq28y8J6EiNClamB3dABZ/4O5NjljkQkDxD91h62aVr544QTFn65i/cIY0T2mo/XFtls9NT
ZCnS0noynw2k3A9mvttB4kpj8fzokpuFfwzn+Hpy/MrCCNfVfX1edu8c7WH44+1wze+hQxVuUK0k
UbMcsoJsZ6HEOdTP4IIlH1ub68V0K3hlSV6br+u2QqxOJezPI6bzyBdqLoL4hM1AYwl6oMMEvHBj
Lyd7anCXR5NSpnTd1/cYv+E42k+/hfPBj16JIo+JtL6KsxylRxJkRho6oxl+HweoqXMB0k25LEVn
Lc6NwVKllXuAt2oJ5ucbERGLAVjC9hqBvhJmRhruvDBesP8Lf2D9JF4l1ljVXfOMEfTRsI3FedaT
EyaBSEkh43GLRQRsci0DAvgyNWfwY0t3q1b/yGDvbIbw9DkQwy/yrmg1y5+qTZjaipiiRViG1CHw
UQPKEFjV3IbjkQIzbtxWn5D6u4gLjGD4vPqjqQFUefA9OeK/oDUEAnX1NRp9wsKlGbtR1p9B8FLa
mjoN4hOexYTObu8rZzdmGtlxr84S6e7sBETrSU7M1+J/ATX1TLXTCxGcgoteoM07l38LaAtPGimh
v3l4dS8hzRnI/67C+r4rhhBVmg5fDunHc61tGmobxiitYSpOmC4zB0nfoNo4X68WIRdllLWpTCJP
yrfKPMSJjeo3AOcS67xkYm/3HGKxgTGvNSQttHtSclJU4BtJ9GMu/MDOjepQeItymH/beOmPeC+R
/pNdh8npOZoXEvTa3Ff9OPl8Vm6xSSTOBEzhCRKsBI9aRwOkCFlAFS9siWCGvMGEEP0ugbp8OAoh
2mijz7twOZ5YBaAcoRckRZUHMLaLPQ8R8pezIqsE1dn+3Vl/GSFD12p2iy0bDDEbKJBicHJ3PDY8
PhEH7HTiVEZJfOeMTv5nQHH2JAS9TBGZfJl7l/Gfncmy0Vb/Fv9jGkoZn61qoopM3WlGdwO1LgGY
anjZkgda7Jv8LhkyQy/dq3gezLpIzac7M3L6+x4B4qX/aY0VBqC40AXqokGH5eJA2BTrcYU08cf2
V9xAIfrSWEMM0fLIemnYLuEWX6gB+XvTMpr+LbEJT+tKvaq+0WseCxvOkBCVHII6r81Qcl1dYmag
YfaUzOWQMUyodoQf2llzj8HJb0pWj6wKWRhbXf9TXu+oItx/dg9c7o7AeRw8RHVQI5aU8mn1WEa5
yz2SIZQ/9hrNa3R1a80X3MH2PvMrNFvwCQIGWX2YKoo7qUJyymhiMj9bE9WMcTNjETYqI3KXcFeJ
TC0DljYO1NERVof/qzUalo6ClXx2Iv1TRJiDqDl6U/9nBtiwS1gBrp2F2CqNLr95ng6KUX32SKfc
brDL1G3KNo4T2Pdbcor4X7fPiljJr2ZW5pneDltVNqisnZXGbyoQ/0SBwd253eWlesoEecDh5VWd
mcN7W8sruPWakWjwyXgmKHKEljYRfJAokAv5NiQBPf+1fzsHchlwuDamDunqVV+iObE8vamawmk6
rsXdVQP//2dirv/G1E3bt23api/IbqiJeaRmgzrud4n9n+MtoAwp7a1xsLytis+ZoJngj7A37f+6
2iHMgfRfUwIwQWLmtt3sxowC9q8FT3KZoahBPwqJ8/gTVlldt3xAqjvMsC3cNbdGjFgQyvkBA06f
bPW6UHOFEjHHLRST1mxa+bILiHYfVwpc6ZP0GFJo1pBbZwv16uvSlP6LhHNjvimIhEmbzzxxbmVR
Y5B24XJZ67XTzv6GLaiaBAwhYPX0hyB8iKbZxufzs5DDYW9uYP1RSwQygTdQS96fena6PYAJ/c/R
MHLKjhZF70NFa94734SyZUDJRrLABFAlbQ9LzPHVLfFRhjpNq4fZIjni/W5bHy2Du8jteN+fu4Ye
v0Wmvy1R5crBeQ55v0Z/rz2anoGKzQW8EIykNFBcjgfLjmKKur//j2MjDwKEYYCN/1h8yYIonPlH
Q+U5EH7do5X5aF5CDqUiEE9qztn0RslL9PSVzZgmkmWFXJesQ7kgo0yTHHmYdyRZ0Er71L0T7tsl
zfcKXsbj2MqiEbsv2YcqPXcZzekaY6UxhykSu3MFiGCcTLeojtFojjgThBUE2TKpAzCH9NaCsFfZ
Y2ZduBH5xsR6Uk33IbaqtvsE9GR/+2YEbeLIe74RNQJNIyv0FZ8ftyTlMWCpljeA6SV/OfARPDGU
40ByAY6mjN/MA/84EshDDszvOMYvRD+xokpw7W9298rINSVAtCQqYspJGHiHfxthwSQCQ25+/9yr
WQBf17l7no1v2jtjR1spTkz+7AnGdp0jb/FBfic2YS8z2aRBz6HM/AfNOnKmv2Q2LHGz1826YAoI
kBtsaqu5JpVttgtmaHK6jw0uV3QLh1PslMboFKAncCHbsuA5N0Gdz11KzBfyI6esHs15MMK3euZE
bakNv6ht+Y1fIKoFoxWHdo8WYl+nV7e2aInPNJgYEQ4K256aohVhewCs0l4BuHlXkWP2a3K87Zc/
0iOvChN4E7hZuE6MUi09cjxh0Qh435UZKdbvXzpXKYPIHP+/k9l5MdpSmiftCOUqPcTt9oGobKS6
AdEbJs6Jv7A0U27z9BAgitB3nbrG4PEcvG9to7LopVVZHPLzuRNLa4KmD+nP9nYYw8G2KSr1g4QH
gYrAPsyQU3AQm/IMZyF+B+vifKbYMeTUB6wuWiqtAC9gY2CAOI8pxHoPxlVfwBlFVx6ojrkBP6OM
Vg/jAEykgPTJTplZ/jWW/B5gwWeutTsXT86o+m+hOKJHm50M4fEQggecs4k8ktXHCkfUOwjYQYo8
9pL8P90cpsNACX9tlwh9q0BOFS2x0TkvmlrNHDXm3HehVpiwZ5xIvTAVxF6ebb0V2awzsUbI4U7F
PAef6Cx4VRE0iWiVQHoulu5bZU+f+Qvm6FWusz7IbMmBkZ0WVJd0yqIn0zCwCLylFONOE2NHwLCj
1/JH4IhiKVB0GsfODzktJDJcBxaHrjZemTrmR5aZrCJ5F5RiPR9XAZNt1Kq8eufUZHl6hY+vtUKG
M7yrbXGk6gMzBZtREqS2it2snpKgE4OOJhm16TK2XrJTkXeudfGgWU/a1IN0CmVeHWgv+bIvfuED
Zn6vHJFTWp5piZp/ebYlxapYELJvF8bdbgtjIhyyGfTGzZn0c6xsn4q488m+FYDrvK66gozoJpM0
9h+MF2BN+qF7rBM0EGsP6kXvykeudJxyKhFnz2EG+bJhSgjiVQIHKs3RUD/i8TuynmRjCM9WXH2w
TUx8UXZYm2j8ckJ9X1dJVmtTHdBSXdiJkWbfnFDN8TSULJm0Nq0jA9wir3yIx8hkLVck/LlhD162
HMqF0uUGtjJxnsdjyNxZPrDPvN6nW6xQT169jBwxxMtnRsUNNBmUl30902b8Gmf+TX8SH7ZEDDzU
jgNLm3qkqvrMTLwHBhExnf2Cxc03bkS1Jr278N0xuacg8JTkq5XucEzAbC+A/OHgJb6yj7fWOt4n
iGeCr2W131cQNxev0TyWshmKGpVF3S7ZdZPcUVVI9EjdZ2jBNOPKjov+zRoY9UxFSTHTIEOHWi8a
VPHZa9qsDL7iYIIKd+hLVb3h23oQlcziNOH6HvblgYP8p5MMhfxmYKIzGztavB0TND3d5h9BsId8
Ha9D5Ho4mKoXSZaDcW5LihD1L0QtcMxqio2KLdgzNcWDp0kJbQ47on4Ek1uyjsIGfyVG93J0Hd4i
tpyanLr0twCnt0P0eK8HN3/AS2oDbYMbV4T5sddJfvuv+eNuNSFoBcYpYNwtU9CouxY37RVUTrJI
HAEGsoY2pG8+ZOIc2dGAmX6g2hLJ4RZpCL8hDh81Rq+ZvhN7QMEI+TJrtHWu3Ccdc1RG7m0+vHgm
vDD0ABQOnLGksW6u7sAA1m36D9r2mqOyJGZWyUAvqc3N6ozMc00tIgpDrxBiJbhvLE7ERpkjqz6J
MTWjcgaKbSZS+yWePxXGaPk6pIiCGuZjIHZ4tNZLhwIC6IGsmPRzLIaalYW0z1CwMo14HF4VmI3I
CLPGT4E2AvnVcMQXoOY/QE+7Oh9tjsMru0hM3fmAPXMzFcRECFpHcksO0TeAFFAvbC9AUF3R9DR2
yyjFGMfZzm8CdvQS3mqNNB6feiVerjMWXhc8LapfCt6Glv43GObGZM2FEiLvPSNFm7IsBwZSlTv3
FwZtSKvJoB73/EO6c2GVeioEtJZb8QcL00SOJPosIhSyrvviWy7k6nMfx+o4xGMJ2w0aicppmYqU
67RV00i9j7eB0rEyvWnkh7Vf3kULkvEuohZY6+MWiW2ZkkJUmVUWVvDFkh5t2ylMJHJqNJN1MJcA
RWvwTIeyahSY4ZV6x2Z6dmMxxWqv81r/C69MrBfKos9OXselrMF2Y202WeSzflefdPwgbZkFNyLK
2qWZCIan6vjT1aEL6yFHMpRo8vGmNduV32tfaShZ9didfKhljnKamdok55tNEn4gAlxTnaoXp70M
hqehh5mo/S4vac/Ohs3QbIkZ/q6IQQcuhl7kqlymGw5cSPW1SfB5UhC8M4NUDkqrnjP+E4up00z0
NEYCp5OD7o1cwo/hYv4VR2e3vYMNdgu64uU6DlY8lwrXPjJ2/c1Gl3h2wsg4UA4W3S8rjmWRIhDm
M1QvsRKV2XNgQKx4WpVJZf/+9xECrzU2Ybxxab1kKjcOjgZxw+kTDccTnN0zPRqmxfENJdCEiJaf
Qlclv/PTRDzviw8heYGkCzqTHtMGJNG+6WI0bYYPPcMPJsBlrYE17BK6Ym/HXJNMfWqFMsd6WuZs
R3FhvzNfqSUM85M7XaTEHfuABorNzZtcGHUf44upw0B+ZMU9xFb5KKmrdnm7OxxNbmJLZ1yKDUt1
LLqVDxZXHjSdunBLPwH81P1kKWQ9uiKcebBII6MvfQfxUNFyrqNFapZFuwggORrYwNwrg5VhV5XC
8tOchjs03aEdMxM7c/YgMLx5sg2ywe5TjcorZiPXH/HBkV47rh+qfnca1kFNry/wTIKSraF2fd4I
K2r9ucPV6f8mGbXCIRLLi5uvf5N7h/0JKCigoBpH3RA/NPuMdvnvygcwyA2GbDcQQkmV8Yni3DNk
jpKPpN5UkqRohLAVLxOSLx7hEDHVjnN37MuL5jrD47WFPq2oIKD2Ftki42MsMUluJfgQIRim+ix/
SsYC3BvCDMMq4z9iUwA/YpGKxaHt8KD3YLyNoS8CY/4HEptBEKkDCptB0RgLVN4MelXsVrkjvGtl
qDgMMvfNb2AhuQLj3pY86sL8ht/dCe2A/51DXzVOw9G8BixEtBDFI+ArAa6+tpL9CHQRcbKitMyQ
7yl5ktvQz8NWLE4q8KtYDouB/8EZDS9JrHy3bv6/s66Ph3dr8sIxOqoiQ4jVEIu3iD2V1F2okymU
HtSduox4mKC0DpPD3/iClK5zCOplmuJjbp5PRxjoj1i2RkGepy+Ryxvkgsqt+XmxQqfvWUE7O5Nu
qgpU3ORxzB0n7cwNB4D2dfUWwZxpHF9QHzCwOMPeGULLaxh7iuRT6Upeb3hLvw0m2bA5Zecd7Mq4
UqFjuY4uYd8LMuo4PHLRiLHpRPjyZsrY+vF8kc6BuUtluQOPS/DiVuE/N30UTvW0qAIGZjWl3ujl
ZnbZl4LFxjv4O3MVKb0swrTqWKh7QK/pFz6V0PgXZwYPlKR5Yulc1A7fZbYUgTKKQ49tcUtQ1+xK
TqbrtbpOLpeo4kGOhpEeOv+xqdHN0etOlNEnLYyskgndqQRyRl3XVqooWPs3I/F1woQeGm5Igs0r
BpI9kgGxhsiu2Y//oyycMqK71YHnjzQrniZkBL61YkyezX7m6KE/QSKJzXTv1OiZa30Hq8PW1FTr
4+WP47wb3b3oAoQFUQLiBVGc59T+dh+MCo7+Yx96tyWb1cA+oloiDBCv12C5LzVJrVryJwhDrUi/
3H04QvBAO8EGztOKbcecnWqgdkAIfHVbNjehjiG7YbaiiXQ7OvnJoWCO+X4rWBMnME2YJyvKabxO
QMVXuspPhjjn3YBPB9osb5bBx3bACOref5qzaEftUrexoFs3VGIvPE0/UO1YYZ0kJMdbWHFNmFPk
T8MYDbW+i7kkGFgckadD4E9kmf6G8F6w26WSxYlfM3x9UurR0FXpWC+gY5KFGVkCAlVEF5y7XFcW
JHZWR4M1csa8z9/VR506IwH2mABsmTtRBKR6ZXUEe5i1XZXiISJb8R8+Wv5G6qsEPlVoU6pjibTj
D1wyaMwaLoZB+tpiZ2eLoXZc2wfRqLswK54dRSga2PFonkTJEOBY5hQpTeNlIr0y46K+U6oMXO7R
SoWKc+M4dCQBEWDdhZF/R42x1UcTF+jaBypydaSIrAgk9GcguVJsUCL3TD+GYGWr7ZQc0ibATSYT
9T4V4K7DcHSGPpMTHBeZVVr0iYCNHppF4iAYkDo134TLs4+zTxoLrbeXkd49JwhYuB+dipkg9TdV
yz9xgk1+fKeUehcjQWokbU59xRDCFI9u1FaVUL2RXFD0AnW7YwrbJ9rPi+AoLq0XcvlEU2ij59lR
iIJUFO19H71TfWj6A2yrZiiwjKGFhlCGupxWj82IK1ajH242Rx5gqHgkJbmxvaP3zxfpeJTRX/ii
i5eCOyqOpPSz6mvc1Fulkh7+SebZfmKD4u/9Q5HuZ6yAZjYXSTDj9LQsDgSpByBJ4mkeAMrP8whY
h8xUK0qkloX+rOoUYE1aozq7af11sIq9MjSMPbMJt3WYc72G5BmK9maBc5L+z5xEiYvVLZ6xvNcU
oInMgJjYQcvFnlu5uJlISFCpL6roQ1ePClfY72Mr7UkPaDdAG+CF0QoE39N9qBmf7g3wJYT78bOE
lqk+cmaGH0baWh1a6yIkbnhbsr7MLU4gVRbOTLELPrg+yUyA6XuIzUD6cnFN5qHBV7z+U9HaY/zg
wG6hJ3gVz0wq3xrXoqW5wcOOOA5y6cskB/u2Es5AYd0irhYFIrKVoN1l1RHNty4NNwHFf/ftC/KV
tVVWxbUrXuQOB3CJzmd6VfB/Y337i0dAgn+rwMnlVDmS4EussUG3CoGmrMA4MAxqPFXaIJmOHEEe
HZwknK0udYC4XNANVoomKiUtvnO+d818YdejCq4sDILAxlS2kiuOgPnfB19WKCB7fbl+iJksRpqF
rnWlFdgmxUW3rq2uBQadPNUbFGiC2/yfiUQsOzN4PRASZOqpcE44nGPk2PNXbzzmDPeE28FIjw+z
z+uxEcJBb35l59yWweciCW47D393x5z7mBg4aOv+C950mduJIZrgkDwgg3Nd6621W5qrlUhETTgR
//yUurhxoKaWvGGwlmS3gzV2y44aqOaqUsEz66m2S2RaXI2Y81KluAxPFMF6xvkkpjziABaN/eAO
ZqXfnf932JNGsf4o0QMErofySvRcYjo+4UAobRY5gvmQ84BITYj09GfkudpumGwm5NfODc6tLWIe
TGxlvnaKBc3PY6JfBT9OgGmouD8ZUa1qEFcEoz5NtuDB79LUqo82WNkDaUyMeTakDSVuvVgYwKO1
P6/e34aO98SSCV1eSIw95o8Owggl6Vsdnf9RA5YSnk6vRunA4AXO5LVMM5Pp9WhpsWcyLqqxYMv7
8WisVmoGJWhQASvLBkLK1v/ffjx8Wd3V69AWyVs8EWUvQ3PkLfS7hrOb6yU9uNrURH7YiZAP94uv
gYPnX9BnliXRLP6r70yd1J6G2zPrZHqis/D4k2Mg/gKlo98K1BRjLRBSgDVJRosu1SRhLEn7XaBG
fzZbCw5Nrre1sSrHljzGm1o/OPmrHid2cWCoOXCZgS/kV93i1obAqmcJVRqG4VMiP7Qj51Oh0qrj
qLYA51LMhmBOUZLpQZM7Vnjzah51IibCzhvurt93Nz7WFhkuIhm9RoX7DMTvxMvBoDAWl+jFhOVE
o5iPRmKdMrsVray7N8cazpAXi3oAwxxDVBrwyy4c4RYr21f2lpAeD1hFg+nwtAhOVFZS0BsF+rw7
+gOueqH/fs9nmIHHXqfycYLHCwCG9PseI3MHIOhjZTGJd76nTeJxNcOHCIu1iP95KHMTVaLUOBt+
8Cmj828ZXx+IjSCNBhVAX9FvDImgYj/5TG6VkHS09ZzIBMWYvwh1o5WFmkjq5f/FE9ZYf9/Yo0VZ
lp+5NhKSZqVjJKhKBY7rhRwYYK0OrEOELhIqbADLqY0d8Cbc57hQyMeTX1CYijOHEc0RrUd63wz4
KtFfpTWrVKzvxB0frif/TmQrW0mhMgsu69czJjFrRV+Sz5LiiAoVru+v9AEbVTyQYkOnh2rOyiWY
Ug+FJ0Z5SIOaIt9gZKxWSIZj4ZUQhukASi85CdNDqOJ9Adde3eB7zOwIJ2sm/dRe/rYNczPKgqwi
LCROrs8o/1evxYGDmu21Cw879q1F7gtxSMms/92e+YCutl3qkSlFGaVRTVZbr8J1XGjbBT9emvwf
F9qL6LM6/P3py+Yen4D/ZFgc9GGsSotnRlDs44WwW8DBRZfxkXzPVWLkQ9PFubnQLLF3mG88LdB0
rE7Ym9mgy9hbC70d0N7dzrsOtR6gSYS88KL5GFFpSC4da1+YZeA1NkEuLnXsCPE86Tclsp/4pN8Q
EqjHs3e/T479XrokhzoO8fVpvMFRbkLEm153WNwtw707r0N+IugwzOBve+nc9pKfiktfHUDQRqIJ
8hVvmSxMdk2j4mRq5VQOAR/m8kbBO2kQEldC012gn9VnhQl6jgo6Xgc62UnwKFsa5/NHJCaZaPyK
CzptBF6ggVAHExYkRZRP6I0k4VVNqdvYuuD42De6dfmVH8RxsdWOfPcP39TLxC54h/Hgs5TdE2Zt
0+OiYckm9y9yc5K085GRgjqPYZD+tb1Ghq0nmPIwU/2ZS/g8rX9CeSy/gXhlQk5lRH1/geS/gpJK
mAdB3OcSbb8YSVD7KyrRlK3zhhJvHWkd0NL+spwRdeibpgI/OhE5KxXacy46JfTf+RsZcG1zav23
xSEgGk+eIC0YMw//b8+UOPSqQ2AAYROtW5fI3RdgJBPTV7cR+7Wog+dyY2AR1lfVoekYk+Ys1qF3
Mv4e04BOksUsJikDh05V3p3ggJK0AX3V4+u1T2oTZQz30J9WEOZ6cJi9GmlVXhSbii7R4QR6PYDz
pt/YsTvLrMvBXhUXSv32ADy+9VJyZ+kkplUGGkhMMyZqBquzAkgkRX4eCDyrgoTI7BGizbwGcHqh
RHU6u1tL4jUOeH5jwWjDQtmyidELCNqN8DF1NlL0CioMS/C5F6E3wUKpOjkgRhEQfV+ooZmFaq/8
HDcuMAjSao5cF42ypBKRSFQC8Uot8JB7EtyAl89U9qrEArj84ynLenntpHcnRSILl+dyRoy7E9yO
6JB4B8Gkcyq+mQEbbyDu+misSq5BC7H/wnKP+xggSsCXJV442GB9tuF4tghft0aoYLPPbXBEtBab
rnWR3ceueVP/etLm/j1p5COUOrMancMdQj3/9IZv7IL1SJhTb/J4agpylU9SYMTGP4ELflVSGksP
Sdaw1swDVt2dq6QkxfyvuAoYIdbuikBIk1ZwH7oGUhAa2RYTXEpRbb+vEVrsAXlvDe7Pj1gw6Lnm
fAbeUOA3c9G9knfMIBNlWt7R/aApdKzG+msZcffcUqNCBwdvQCnSas7pfP7c9h7keSOs5Spa1/rN
0o7Pz2Tx8wRjpJEUCSktCG7LieVDKw0IADdDjMqMUI77P86T2zPHA8z7E3RCCWYcr5jygj8Zk3N+
325UcTf1AD+ElefIhr8epLX4eoq6+r2xX32XFrzVk6G7Dcj6XXWpfd0QT9w9ZEIp/tGQWsasuipC
sFVB7ImQ3HXJK8gqWiVnsTmw5g4K8EW85WtZyhjZV2C/ypYgFATuunJ8qDKNm3L8VsNdISD6tmGl
z7NXVG6nrO+4AMtGmCDK5236X8zTcqYyikP03QW4GCmcTK7TNsP7tW1FJahCGWzDsiiO1Dwd+up3
9vmLClJ4yYdeItxCkKySwuKU4NZuREpeKle4TPUP22BCo9bE1MtH9Y7poQTEApopTuvRWfrs3dOY
kWaJ8n8RG0hWtY4qdBdS5pX5GI+8IBuTSa0rsSIZ7iS2STZvlouh0ocrT9r8bixmXICU/8HFtvFM
aqP6ikBfPlNFipcy9QxyfVzhfk6SXurspbCIw1bSPjrohC2gHYGfLRQlP75GoIidbiDcr+yokRjJ
7s32Ui9V9UERIb6wrMDmgCQPSdjELyaM/6MRORaECqjghL8ZzyrQPiEnxK9ywSQdHn/rbcfsuQ0O
lmn8SS9elStbiiJ52lQI5YJ6Xk672poR0mUDvpqUOUmhDJSLJ2v0xU+TZfC/HbVOh3dWXEV6jLxX
PIvsU4E0wHhMFrKoqEMNmptGGt5mBN95tdMyNjdXqZ93t7evT/64bob8D3Mh5ltE04Ah92kGNkmp
yy00gfZr+JJgS0R8uVv7yuJdwrTErbi1FXqpEHJB9J4Z/J7Un7wequlFWklQeoDzySce3uLqKiQ4
54rXN9X2B2/jWpx/J83GXWSbz+xyX1m3n3cyq/IWt2ndjr8T8QCvB1XKqYjYLiQH6BIo/U2HkmVq
kRm9PalYfjZm9qedNMUXLTuIktvOSWvPdSopWx5BoIs3y2VsUNhhmFiIAiMk2r1NjAJeviU8UyFS
PIXVZOBIuJujMPSClEF4CQ8uHKNpuxhMr/Uw5tt5VH/8F03fTeU2hZBVsHEvdwH5YqugucmM1FFB
LTkY/VzbwEf33gKm8WCFVHKAWRSje6mmUtdQEYs3QtuDdMJh4UmSFDfAktev1xj+j/z27Vsai1oV
Wb7EK4x8BcZNdBx3qz9bbNXxh+wjCiM+CZipyYyJIAURZR8RSUW3bSkQZuylRHV7+q+m0dAoydLF
KSwejSlDZ7J++splcdKEMySDoXhzG6BR+L7VfMjrxfYlsPEX/hHaUiKobSzD0Z+5g8QpR54XxwEx
Aav1rRsiboFvj0kQtLCSMTACG7iuTei1zdUS/x2OSxTdj9hM23YwROVzCEWlHGsasjpujlVvGc1v
W76b98HnwLznV9EZZmWDq7L2AyHEFX1CNsmlMtyPsy0XhnSwIgyuBlA8lv4XdB0CMAjFZSAIZOlW
1PA6DrLI6j3T1kQgueTO5MvwwPpkvOTLtBNwjNnRKmSa/Mt/a61e2J1FG0Ad6lNbnwVoDKC08QuP
JxrLo4eWxnnE2EjD1ROps7x26d/c6TjtQOQVehVJ9/LdX3Bbp80S594F0Yqjwoq1hwCiBSiQ4N8U
u1ys43hF+kq5R57+TX1tHWIV2qTPl1QI6W1rvp4ic4oVDKV2US7A5ceakaiRwcnTfrEDwnvqgec2
b7EdVCKvXCKzKjq+OePUHd5QjCNjDVZ9mWSo8hkpexEhbxgqYaldl/HLV6Z6SLN6XVm+8ILfW6SA
N3gvP2/WOyzrhK3O2aCOeWkP+kGoVSuhYSHda4c/NSI5coRrcb2PBHnKzqtQWJMExo7Gxlh5yWxs
+vybhdblMZkgozrzTxz8d/jK18kP0DSU3vh2IjlRRqf4xRWdWJ9Oy6qDVcEx1a1wf3XaNZdb3N31
xXOgYz8zU/JPl5Ku/ePxNcdnd0HkJmgbRWBURpniTlQ2gB3nrAK5YOHblupH34JSYqp+PQRn+Qyy
464eW+Rifo8f8rHSy9mBSnP+F6/YoGEmHl+ep9bWDZ02ZBlZX7Aje6FMM3UXiWGVl+I5K0RMn5Q6
kjIaOmaCrIWQL9SexFD7zjur2sFfN199xzbVed5Zt9hfH7x0gpneN0BdPfqJMlzLV1KTGVDnzQIY
3T3H44W1MOaISe5z0wYKE+Olwhzu7CHvIaxHjK09/bbaoFb+ndQd+BDQr6ovBiTDky7AMUCA3PPP
86nQ3C92I8lGJ1LGFpRCxUaIDMGyxmUU8cEYbmx3OnYbEGlrx44mK+T/JSCj3AhNJzFRmHSOLSex
NUe7/DRH3TbJEYvsMqBew9p5TYlzK+SFbDepIiaqlH8+22oBi8amB//y6eNKTTaZF95EMdv+Dg18
RuDM85TigdUnI94vh2cx0D1Y/mEwJtNYi8cg2waWzgYxA44QNtL2ahP5vvKCgGDt+fhJCOQpYah3
maFVQYsxAjV1Ng7kyXtT/3hK9wdFJLEdE24TBECQS9n1j+ZY/hgIPawq7ja76tU15aN1lvwfiYQa
v6FYsglh87hJQDmn7qSsR+z7ctWQziMjQVb7GQpJFOLuNXp0De8+cOZf/MnF8AewJdw8xBpetE3e
EIw3P/iQsz5YYIYQZGMAF+bAqOEyehqnu62qtdCmGnj8CYMxUlouIiPp1X4XTVm/jQg6I2jlK2un
jpgH/L5O5lU/U7iZ5gwWrZ9LA6T3PiejjtH3RqHhWqAmT27NBaGftCCmg4BC/jBj4DxyfTfunUWk
TGT3FvO1yH6O4fyzmcD74XCrhAcZnWOfB8lWth3d4lgiMoj8XXhgkieADx0ka2C+kSvpo4YIIUJj
INDPiQnc6VUF+mNI81GtzwP7O1YBVdN2lln6LMQumla3TN7a2byOXn/ejIdKswIWgh2CSjCmjKpx
dlgxd1amLzRfajPjVsYPfA9+URZCw9aM/5yv9FyjGPkN4MZIPeu9A/d//fjUKnih8hlFlwC8WRxt
+tvhg9OuT2b3uZ9axKxjDUL/VdOUZ3ZanlKPJYnJkAUV17kid+YHlzi7gn8yUuBItwxExRp5xxZH
uo94fN5zCvB9hyaFWTD02dpiyApwyI1VzIQcSx1mEfO1VY7BEz8OVz3DZUdJbw2sfzHDN+YAL7yA
ls2X9Nf3jGsnD90h4G2Lqx2YrLxgrJqmW8FPX2M/QRLNeNRVMM03bwK7wvOHNayqdo2ibltkwge+
hzMTGl1vwEY0MhBd99V8cQtO/XZHE0du/oTEoyBDfp8qKzVLInyGEcenFYckajDm6KwJHgQnJc0b
8t7TQJyRW+Ec5iJrEJUPtCUJrYMxgASGvXTd8jh1nPkCj7ZidWQT+xRknD+IZtd6R3wR0l3WZlRD
rXoxhZ4yFBlF8C0cVTn+Us+Fklqx9Zj/jTESBJjtLkb5q2OTK2Enm5yk6l9+M9SG1IwtkrIMKfn0
4FfxC5tLfHBJXQbcEuE0EDmCR7GB9NbBFQhHDBJ3pT/Bl5+69EPEL6yK/G77z8LOlM32B1RaX/kO
uB0dCkJpLdsHKsfixT9cJ03wwli0YRbanJI4zDjmdOeI0qzird/AwNpyPee2C4jtcB1G7/jn/igl
604m4Q2/PJC63lzRBxXgm6lFeKScQkcrLUGMoDr0Vzf1PDKW7TCtKEAGBrMLrjypTVD7qaFBzPKk
dy6OxShYMuCau6Kb4q0FO5KvAGBckniWfrjHudhQelGrH/Ndewi2YcL3IrnsO3BCy/MsQ4vvBfBF
RCKYVKuRNAu8LBRjHF2p5AeDkmnAut5mqZbeOyNFMSisRTik8/Ll/pL91JosCN+UzTTWwzRb3MaQ
kO1RzEc6XlH2wDHG8muF5mmmmqkSw7LiLIlqr0KYKOgJOFHUD3gGkRfuyOcQST+ZB2RbyBgbMQUH
gLMHA4ymQVg6XHgpMvKM+h/xEct7eW881XDviSSaadLTpQlGIeCTXdiBaLmJGtzDkyJQnonkYmx/
S4qDC3PyGGfi9tI/IpOSw8yVAVCpUYkFxCP6YOCxuPM6XcmEq8mQrrzN21YFE/pJlftjpXEGO6n1
cfrLDqBxVwPgd5JnnJXlqkZPryQGdwUZCtpYWoFUf2beXieYo+Gits7iPposarw+faCLm+ZUn+dV
GA3S4SHC169A2wmmYqBWe3GHKTNgs1Cd2zW10EWl7z3P2tXkAv3UvfO2jFakuEAwMe+7C/SS/d/3
PXZjW8WJ81YYjLXnjH228SlX8VgLmyUt9bKkVHyZSIWrVKuGldTpAI9Hyc/HPbRU3UEhd2KHBrdE
H0ug4RgoGUuD8BUaP5xdZerlcFgcjrFsD556cHztWDmrgzlwNfE0vw2xDjyvlEBsZ876PmXOOMAh
bel33PMJaGyYoicyc7IJYX8cr/bHXDSThdx8lH6lgvWkJfOSRozyGh1eFsBwiOReiOcWy5BBL6Bn
oY4h+8WSvZhI1AtM9nD3JNfG7hccpMDxdChgAsrWggBVLfmulfI1ta7ob61hCEckmS9hq0GJkduZ
MF/mkvW2Zf6acvU/rAtS0SrXBCgRfM0jHwLChBts/j9CuK0rd9/slOz54qE+q9qWZBm4ZdrSyxKJ
TRt9NPcaWrv1JnAQ5VQRlLGE9voyuXHPUEUGURwRzE0Ls3FsEQvFZzdNmSk6VgZjeJlGFVJINvnL
svb22KVrwp8692brDJ0kbWAlr/IwmRN1CSuiyLpfOMaNG6FEt1IGT52MRf2X0S8ceKWZx3dfB/qd
N5wdde1SDojRY8NSzH63nU/cUPLASJwT0zfLce1hqKchWjbotwCWH2okyxf3fancNa1E3gvL1Rdt
AWy4mez6Ra9LenQHHpTKe17NjjBKMYD/d2qjxBQ4b41o0Z4fn5EVuq3nH77RvDyd0qdpYemj/+Lw
skQOo9vFS+CG8Ll4a/gdPCAR4So7AUbpB3YBlcTcb6rzXJvKx3emPAe5Aa3AiNk9KFog9JQkUMVe
agkYjpxcamPh/uvogOvAs3sAhtvspDBUpyWclMZUtl+/ZyfMe4TwiWLhmGvGZVzbUDVRvChWxQcH
2K1cV2Ea0kcawMTOKUkriMtIb2HfcPx5zrHSeW9IYaJgyxiNopDHZB3rJh64RdDnUdU7zL/VpMSc
l0AY3GgMVqo3YCmR/Blg92cJIeLZnazbqorxvCyYBoKWOwESVd39ONqQIn0yzUbGpwzmj8a4qWt6
6roTVOYkaEAB9yodHFd48MfNp9nAiNZBnfMtuZfGz4QQVuZd6oCRjzXcMOK7NIxTPSTz9meUdeHC
kRCU2BDc8Je1BodgT39aNlOy59lZztVOMXbAzPFBClbafJbVBvYTZsQ3Z/1SpnFNZXgwZBxxijmB
GegLVpJEDK0IiqFdXnZBsRIyEJotQKSXn/1nUO2mrh3zNoy05sQNBTk1/X68h+tYgGXAf9sYP2MP
1aEqD+6cep1lCAeFcVA+AAKpRKmHPjxCmm3H8f1kV3bhhlyEpqBE1HZt1S1bye6YRbOPP1JsbSrg
WCaSuDshSvGQdZqAF9JRHKsYFuSSEISEQwyYJ5Ypk7ZV8FhUGzpB2AxU8r/xQsNTIlnQAvpjJBrc
k+/wu0KcMj4EU9e0p6lqAb+km3QAJeJLCF3n0FuW2TNtJeChZUAKyjoyItkBKzcirgvOBZMf7LF9
vUfNszb0e5vbD2RyTCYSZXsxRa2FxJOxSOKdswWJPgUMyXuQsi2DWbc5zkMeSldAyVSF8o1YAHdT
LWjLBtpkvZgXnxSneHHV5qE6hYtW25tG+OdS++YTzOLxEnocqXhrNoZmF29XFHNyY2acdDCGRMEL
evFYKKWZZkKo+odr/rmZcMqKZiDqqSNp07KB1rTBF5s1lAcIMPTpW402dHomz6TfkkMVsQWq249S
lWMRckItkDK7N0SA01Sj5c8Urp4qpn9FS6+z+zIuuZK+8e5NnkPUypYg22KJ6ui9Tpo3eKvXU8jq
TRT5HYLd+g5qR623LQMIzdUAoFnkfPavL8ElVbJJgLEl6/GoZjwW0KaBl4nIbGHCS0YsY/MgMl7x
Jrjdgn7RjFq+4G4mjHPTdPNlF9qw/LNFN7pVzIT6z6Ea1C5/tSqTu5p71r05NI0xUp+aJOowWqvC
VGEZmeJ3mk64dbnHbGYk6Ho7u1BmiG1V+QcFuhgJPk7Ox2j8rTcOqbd4zHPV41Y9YG3s4nmne3Fk
LhR3lp00N+EjU1j3D/OD6r8CZkUCZLCPzecU/w+xHCoWui8OdMw2BFKIsW/L6PLJDH6gdlk8vUoG
pv+uvoEOZ8h5q+ROt5/ZLWckVd4O/wf5fODIfKo/2NfZ+O4Dakylc3RgjlEJ5ky5Vu+QB0XH+5Ao
CZ/925OcdgezZxjlQOseJKPUNH5mIgcmingKEH9y9bpukPjNDxYVOwW7E80sFHANUEjlzus/gz+e
ZsoAUTOnY/Y5Hj7TluIFokddILf3JUOOrqMGPaYA948FuUHPipu2eucwfDOZkScobHqPcqCkcnZN
YbTHWCpBP0GY4PUsyiJY1p/WejaJRnz69yxy1SEJ8G/ZlTz0BkU2b29fXv4Q+rmBTOGM0+Yj3EzJ
0NAg4iwyeWLUd0Lsa1XWt35BpqXVz8q6p85ck4Oter9IOBcncYiD+JnFgYxgxrSlwIiREKHBvsmH
GsoLZPMD5E1bhXxYG8wxY9L5uAmXSaC4lCD9ml6kl/ej+LgA7oZwMdSk5fGy9YdpJsBQT7VDmkfq
df15t4Y3VyeSJtXj0MGUxLaAlZVdsASY7F+wJz2e5e0M+r/vqDzI/1bCXB7K7WdfyyWX31Y/Q6sN
JG+uOXnX3FHKGELq2Q89VopxPctTpUiVYaj0CXQgrQsOWaBGMt2d49XMuBwHXyPtu1ogH6QevtpE
ivp6+hvLskNRfoUsuKb81n2Q05JBY4zx8oZ9W0bhBREiI6Xfjpfco8aieCijo4kY6iQpslq/HUDO
Cl+WNaBQW8PjxEQYnOmGYP/b6vAu2FHFySqTKxeSmtIVpwJuZtjpZA3g/hKIwW+wg2F3v0iDrDvJ
dKZMrJmWlrPDQsBUEUM0qDaKB/v7nowqAlvezVi+htIeQMed0X4mbQRJg/veodKgHsXxyVlYqoVv
IwxtxdejPU4hv5C6VfHuW9PR7v/M2Ofd/vrNanJJuYtn00YBK8aOZ+xs6lKzrwlGV+TEV0Iua6at
E0kAgG2HSwmd+1fpbSvfFMVyes1W1ztEx+v59RkgvgW8UZtdV5ulFH0gKSDshxsrBG8nsdIqVasU
BUP9EzkRM7McDNxD7TOWQMRLIh0EWr9Dw8PX4vTcynzB6OW8qjUZTbhmHwWIlbBB4MObnqPfoU2Y
qIFjUmM4jQ3M2hO1KBoz6MPTfjsUAQpfQF9RHasttNZmGpJXCsEQ3gZ4zIQWdiyZHdU+Pnvq0mxc
h8irxK+j5uWzS+GCoN3u2knrT6Ou52IIz8eknvxeLBVDU3kl46Yk1Ahcp0YMzGfgCsXwN2hcJI+K
PIyG7ix8LrEiN1E5wvX8fZUkMEB5IG73GuBe3Kqzk7tK504Gn08JfR2nPVIUJWPxPgdRtFBBkC3Z
KAkpNWu8cUDlm1J4qe7TeFizay2NNDvglhIID6Y9NFaMDciKLgLY4ch9tHCe96fjeHT8eAAJ+vpY
D1T4DkuP4DiSNWSgII4Ho60L0fiRdrBcaAlEOQ51+u2hYGQT8DHofJDqpcXzE4lVXKPlK00nthca
G8yKrGKArDCgdqHSgNSzLH3XYmDheimox5sZfr8EOv2OfenW2LlcPcbg3yfTSYeaTUmRX0P0VnzJ
Jm9ldBCa6Cx77EV/Q/DVwPV0ney4x1optPKug1PzMERf/VeREQaODvr0NWuTZ/8fjpzRZia3n9Hd
t1cuO6t4vAKooC/2+zqhlBuwjvUoEYvDT+VZM64s+BqEOeURhzvc+qKazoT5U+veCCYyK+66btyV
JzOPk55ouo4wbbqg3oYPX29CDhFMWBzIuc56kcr3yA/2MP+jvI+crl8VTg4DZiADy2h9VRM7iWzD
LDZls3V2PXNRtK4y8cFkZSEDW5LgJ/oXOO0sFqAMkH4KReP+1YalMpK3tRNzsHTJtdDh5ucp1yOu
8ec7s8sH9n0HqUgtJ3JactkLh+NeNncL7ml8C51Qg742aqptjEu7MzGeMvEoYVEM4jOYjHiIriLU
bM5gGAFc3ioBmnIb4nCMLo6tjbTVy42RlMq4rn9tVvxVE3G/SRp5xS70kAid450BrN6YQ8+WyudW
tuOejY5wfl9rLKNIt9MmsRhQgWUmyQ2pHbJYcSL8DWlnUTpIAZF12LrxVaGXkEQV6E34VdtVwUmg
Z6M2bKqdk0PAVSsJDkIzBR/sQc9hhkLRZLUW58+lRJZVefp5ygsKCRl0CI0v6vpcq7+Sbk7kEgrr
0iLk0LVgrwSOrMa2CuW5GCtB81pmCRzUy168x/2e9twLdj+pZT53ZMyioLVviYHBXcWDRT5YVzQR
v9Eh+MmgtCKKzx/OYrulWtwEQSZHBR3hcFJ+Kl90sPsUHzC+Jv5UN0XnNw81yMgmE1FGuZrMaSs8
qSbr6lIibwoCL21I9PtUZ+Q8ajQFtYpCK5GMfRxFCcNE0XZjSbtQHqeyJ2IFzW5TU6K4l9rZPsu2
Ke28B9lKF+S+dQoCd61wOw4twGqeLcTCojG7t1XHUsei8s+xCzRxB/hb+IRsieUnSJuvY8OaAZLL
VYx5Whr5xzPkKpJEUXudxOY6/t4wX6R7PnK43Yzg2mPkwYfy9x33aqtfSLUq8YOnEgRniYaLR6lZ
96Yz64Cjhouw+fgzA7bkenNRk+/L2b+2wAN3DZauVmvuv/sgnjw3LKayFieYgbyWcf/p6gmV3ekL
dTn4GBmWm1mGG/FxtWjUjbfB6zUUGCfs7VWYmvkz4GL2f+bOQeIEomiE8BnM8Nog6lHPIgS33keb
rfEyh0RvHvKHEPfSkfGBqpFyx6ZblURRWZqj/tX2MNuS1qszPNS7Tax8qyRlkStasGQ11/RshyKp
sqP6eXR8ZRk1vIMnHsc1KgrDeVecLFMYO3KV0uJ/CTWXDga7TDr3Jm60YRCROrCJtdNgbWw8atNy
IBKHNmbjLNGiDQwaBgBjjPAYDgqxYco19dk48bdTXi3eXmCw6A93KYQ8a9DZbmpNbZ6FBLJHcwQ6
clglC2Y7N+u3bMKPBQitPBr1sIOKBor4Ed2fAjyjO5BOv8Jwq4r+nEpv0Yy5AZvc+wFpv8U8Id1q
jSJln8+l2tcvpFReBAIxoClPpNEb3tuSYlXtIishCIR72LQH6gPsaJV0hAhWZwDAUUo83rwGfi1E
PKuvY6YJwGKypHBVzl7Xwrpw9MIQoVNqvvqlLSgkw9tQqmVxd//b/wAgGD8w41H9KFCsyeysUb+6
zQrGbabv/lGKCOycWVCBvN8NwRg9CkvgbbREaVHtu3l4dj0ZS8mNTJqKRhlSjadGY38EXQ0lQ25A
kU3IM+gfsZCDJNXTKyjp987EybCPhQcYgUDvzAmK8yf0rvxQnvgYAs1R/N9Hg7wYT9mtLK+c9pPl
8uzJp4g8qoOBq9GMqA+77DHyTP3oakYVy0TcZtyCC+BnOJHDAvVlwNZfTekhBUUnz+JXgQGri0ak
1pP4kosFRr/LUrSaHg5k8LeVfeSGH6tgPpsTmZpxJzjYkWFypkGnnuaJAt2WoG+scYJrYW5p1z8c
PRSB9+LOZJM7BB899R/SE3szF8M7DszxXKGOWA+XHydKkigBWr2S5lrskhuSlrvM1GEnwuLc+IXJ
+sABzOrc2WgF9S8zFYsyTmtP5GKgtu/eiGXD/zNjR8dzQcupimZOBX0fe/G5xLWYglw+ScNwLUx5
vpH2J61xhn5B7TY+15jz+XfryTbfp+tMxWujMBgkhGy5kQKBlh0xlC2A8Q+ahwcDIhOEp+X151Em
nArjtlDcaLtaNxQM+kaKDAAAf7QKtHG5/NKhd844KPOfFjfIqPGArGuiGzrrVkCzzRbu5trPnq/7
uKxlREVx0wkwrEXbiWXi/nvQY3zN6poCdBo3x4T3jh1A03nfU9eCpdh1biVdfXVmBFGxCJKZCWCL
a/puD87aB4mR9nCcPrrH+CbjiXLqhWWnkVpLcmc/3latjS7dpel2PK5f3jjpTEeGljg8Ril+9Ry3
AXA/cY+3OC2RT5HY6LWt781kfe1NRo64ZsJL2NT7qA4cZIQL/raPEPsJy0pv3SMaOTXm311RYDoQ
DvoEeopObonNrJFx8k9cw9MiP1JoAFkqyjBHC9gh9twgq94EZ7ip5Cm0Y4geO3jQlKReTBIs4gId
PXiVTw1apcZ/hRzIWS5O610ZqTbbpAwQMcqbe1sdiAvy7XnLhAyjJ4SKIaWo+rDpZmuk01zFyjMi
GxH4EM9p5mawSH5mBmfWpwdWjvCYYkJK1TqMKep2fYIUaOPHzdvJoFoW7zAWic5W1IrRj2GmpKSd
Z1tzTMy4xRySPGyfZzUYFTw+KKJnbwib33z6iqcyw7yX1zrwL066vcQkn1e/YjJzax75MzwUwf9C
GlsmfECnBvBpK99079iul/+XG7pSGIeU1gCBIx7SbJqvGtu4bRcZnnAcsV6PuevPigFx4zt9lqtP
AHRbiIcthJkAfZMbM4tmUB8bxeqe0p7SA0ASd6bqldRWjIwtP7SXGXMcUbeYiVFQZ0pO8m6vOoOf
RkjRwTS84iEkcUJP86WzRLmiiYgUCrsA8jTEtkM2GIKkDLJZY/b2xnIcryVhl4FCMPDkZ6Er84Tf
10FkJYn65cR0+y5xcJDShP7QdDRZ2AOfM7BJYQ1ADbVc3rFIk/iCwQSZUd8+Qa7bFuo24YiyvCWr
J0N+EB7rhCRpU+mVrRi9k99Lzqh0OFwfUPvbhJij9/LLLGnY0n0n8513AsWRURuAHqtX80S7Faxs
nwxbQVRXjzkPqvtBtXQIN7QC1eKb/dsvnIFynC7/25jIhKnfkJ7kYD7eVuf6Z2/ox5r4gQjLnrxf
x/y65yDWsojnsxzxmsiGs4hEehTJ9o6YePfzZnnEUzmL6C73IEzQq/7I4zo/q69zZrF3YE30gRyn
90Iqhjrn5ATFOLxYFNgbqNPkKM54hDkuJSR24q/XBHDjzk/lYOCXR2WRl0oi19xed5SqcAZUnLcm
Ea+rWgbY4GKidPFFy5/sD2UW3025tBt0aiJEmi1kWTrz7JfTmSfPXrdJK4DeKmi6iR5j3FpPFuJ5
7yXpcsArxYmcOX9rTMyyYJA5ES11yzWj6xgGj87+5uoDPY2guupYTKG1wC5E+ROgulDYmUblVLcp
TqZeyHEfifOetin6oT98xlCZ0gZRmXJe5RTp/M75d6qXCMGyhVQ1+g+cbpS1KFJWk9C6gGeopkXq
Ehs+aY/TiMd2gm+H3UdKVeNmv2qRxF1N4iwo4N8UrJM+7AZSQ1rpW/CfH2foBaqwRZpT7ibrCzyT
eFa8os5G+ExlRcj68pT8cPD38eXB2e9lTQCWI5fUPh+gIZN16uw5UL1x2H4PR0vlGXCuCkLdFcRw
P7X8RL/nHzAeY4a/NY7V+sydiZqJPx/ePgh47tmdcKVb/ixbPsj+IvPLNSxRFBkRUvPG8cN5Yexj
/PbNU8FVqAM55SdjyvUspbWOULjbsD4GhEwTvmf+z4PgY11LnhTI4JXlgte+0OB4JSznvbJrUCUH
QbLndPppyUPLLm7RUoFqmcTyjvMm8ND9nkJdDWWNmLSm8Nw1P1wB8MfGonR5BHgf+Fr4afCjmVuL
urRbSKSV1MLfccMzaSWsbKJMaSKgHAqcTr+xIeLsnTpeuoaapobKV9mV+MXcE2JPhAi1Cj0RoxEW
ZNdTWnY/TobbllaM4C1ei4oLBqab6SjfgNtk9lS237SWu0FtIARb+92tu6DPiB6XhdSbn0JrElfq
PS3dc7ZnLaZg5Hl7Y5zZgVcRQ2lmi9MkCbE/HxGMInZWmDra0NRnlYqkCpilsV4ql4Zusguu3URM
AwB10De0rcF19nyl1UC6FfH1DOsbaDk4pxeTmTUyeUQlRNj2irtt1QZKXww1g7XrkxOUrTly26IK
kpz2Vu1BvoRsZj94tykUM2kQv2rY6UfGG9uuX3PFXV4Ic7CPkhTblXnREE6pn8LPWelNxJKZYPXr
tYD4pWJ4VzTWdnCfPw5I9+xBezmHnJX4U1U+bdjwxmkK4DwXBTRB070OTKLWfg/poc2m8t2vR1s1
W4ub19/73IIrOymq2o7ztn02eOwfimhxUTqjgcooAFWWhjx9LLOG/OHf3c77jc79JonRAsw4rDCb
U0QhW/WMFRqKWdEuqaYdrqg3QjCkrUm7hQIOl630LY3dS0IbTX4P9TKXKNvCUKQaH6wdRtdhirbq
q+dbcRTdnByplmFDzym16I72QfWsWbb0J0+V1kkzb6+3VIEaylIg/OaCmIWYXo9RUtQtbkVSVqzs
urt3W5NsEWICKSSS9zOkguR/RYNAUGXPSAFufIpNLwqyCRju3tvSryrSZutqSQ2WqxK908PX2LSp
nthwtfkDT5ylzJMpitX/p4nhDvUSbucODbJFM8YgkfpbqEBdLl1gl5KwwA3QrW4FeRJFG7J2AUfB
A427x6pttTq4yStxKvUpylb8aXTcGgNqYk5ZyYLRZwQzk43blyjFLSfzOPPa8yA3VxNyw6JSY+QB
oDET7BkS/JQ63bnBQ5gjKsFIASoORoSresgt7fSj1QVE4HFU0HQPiFnhjXy2SvfQf9C4I8U6Jxu3
PZVMcBDrBvcILzHpA9FQ7vLVW+oA6hgbAwyzrs4x8Yadd9hGMK2DHiVjnI6mJCaEfWwkRpQtRdgJ
l8e1HisPyiWrrw4XbJG2LleTx6FAh2fjk5efAt2K5iSNR5IVAWb7XxihtmpSYuDb+ZI/oGGz40iA
9smZQvBbUhmY7lhE5rMazpSP8o00tYgIYriJjlroIsF12sR6NGUd3a6+DHp/ha/ScrchrEZZ+DHH
cFYPdDiJOU4BKnOiB+fNQF57y2Z7rw+a1JoffGB7nlVV9OK0rZZfQDulNOFgUAIg6MHhSqZbaT/Z
CeUUTQo50uHqrpBXtmkquj20T2vABvA3IZYYvCLCIXDTIQ9Doy/xefcyl/s2amx/NNtbdkYyHjMn
TFG+VWj5BY9Ex+5SxJRILRciOsl3seLkim9V9Bduq0jUnhf+IDkjyX8YeG/3o9lX86XGr38s/i57
mODy+lVv3gUgIWII1qNdtWEXr6qXG/mCHGjYPX3zRejT92orip662wF4JB199K0MRbBX+dwzf06P
zQJtVJfH4yhvrInp76tDBMYZSDMSTD10pP5Fxugyv77nhE7XULPPRflXdq+5pYM2jLZQNHNP+ouE
JUGuAm5au/pgcdNdfg2YW4CAIPoW07dnxkNIM1nGHDpQTmFy8WLiHuhFoNO3pSH4n6DDPT5uYa2b
uwjw480SI3+1uHlNGSdnqowH2Ga1Br8scv4F+GognDlrb/O/UDnFX07+SyBtPkhV4YkkADfdh6sY
EVhaV8iul5L4sjCzMhQ+ubbJom3G+YE6IxqVnWXYGZdltzaVPY9uzLS06rvZVNGVuyI9IuhY6+7/
sy6vij7I03MuSiBGLHxJCy0s+oHwqWNrYie5fCSShRJ4aCfaOrbLWijQWqLIJvzQv5CeAGrbiGlH
5HRlocZV+C80yxcRzoKUMBVrcEnvDL3wJoOwK9x47WVJY2OYAVWaaR5SfQgL3B/nCfWk7dFFTqlZ
piNhP7bj+MRYbrFXlmW+ox8rV1grLnqjOVN6A9gWm2WZ9ZYcpZOZ+8fm1lfTWLXbJrx6LJyeVzPX
nn4trUNFK/CzOCwac0o+3yGY35togZuVs1ZhlhWJSE9c3LrunGXpvSd+t6VJzG/YJLgl0AFed6Zb
tRWLbo30LIgwxgH80IeWJU/1mMnZAuW0Kna9fq0fSbGCZutcRxn8QSnZEjp037zWJl6C8+xMyzSk
n0aEDG1W5f5RdK90mEhJ2PMRNGR3e6ls0iigQDdrVx6qz1pzX9haTbyA1BRMc+VyIi09UMTmyuwU
85mr8Qedb0sk3Ce4V1p6As9UrkNr/D8w6KS7AFIhutRq8tXgdUcB+DP01heHX4Vc1M+rkIkqaSxH
O6tS8w6V5TaKEGWBgfMd9w8ncs5noL0py0yOJ92idk/fdAXc/kc6fTO3LhJnHD6rCZUiWUxHGe4V
Et/X6n0CcwWXef+cV6rWOHiHObLr47cIHcXKVD5V7hXAPQdziA7LEYPDj6aaA0mcDshwFhp0TAZC
Nf9OAOIcGgD1C3a65TPpf+woCjI7vpLX+fA9cANSEtaabv1skWXPdQIlNV234d+ZrI1BONz4Iyhr
jQOouxpklx0NfTNWu7ZcKanaIRTTQcngvQ9teAexBy4DrtwLQYUr2UR1azGavi9eRrsxK9aPVo5M
hJhKaiP7NppwZ8wkww0aXg0AKp06G5smnJva3eslCvzVUo9Fkwp205JHwbVQxulCJYSIzssBVQfD
Hpup3u1/7Lq5mX4KvCHxAFnIzT20Mo/Jy0YdSkg0BFr4Ov5PtyNEip3m34PnzR9f9wClZ61NVnjG
09bAyz5eV68+N+xLd3rQ6/TtgSc3TGu3LPWRKFb2m9dKUoufivLonDDzAPLCCSjj0HVwMcWhBkoZ
C6CAygxK4pu4aQ7Y6kjc6WWVHHEOn4iw08zrBNBQ5ufO9HB4btXwpO/0mQOIh5yZCdI0NHZHYcFE
yKtQzbsihN1FX9Gu8hRykzMl1aS1JNOesRa1BQQlfj5wU7H1dexjB44lgLzB0IIw+z7NXtpReSjW
yVlSeOKfk41XJ5L7sqSmDkkelQeVWd1DK141h8Bkq+gZgH2pEjcJncEGuqFr5PmeO/M7P2wiMTRH
egzRXSk2/AIywlk/mRQmhrHiZqWVJxSbqSdNj4B2B9fjalLdDj96dAXpvkGzN9EtOdduZ/LlIPmG
CDWrw+vpcJkyLbfqmc9zlZgWaOx2NbDgttZSRY9U82PxpSBY2+XAD+5+AwWMJYclIJwHnAtkZGzK
a44OzGO8VWr4YSuTUPHfQdTTAxxA5L17W6UAUXIdEqk6PIL95Z857dsZdKR+DHMA7k8Sp/4RdHbj
Dl9m7zCb5MFqIQ4PdD283Sb+aRcJjWqpy30jAhKxbDgTU23ZOdjVE1w4+nT6rja1ZX7Cq4B1BZJo
ML5TJuffbbJb2/chCfqhCQ9sKPNsYdJ2e/qJejBs1PLaBRRMLRQhzYSv9MECeHuAfdtzN9BwMnyw
E87ylGOAJjTp3F8E4SY49af/zRWWlXlJZBaatdF9VKXnnKTGM/+4foX2GWE3dgfgfKCeOKhtbKaQ
ll8OkExCVhwCUmtGKg5vH+O5uLvnU+/FZ6LoVxV4vwSqyUVM2WoTo2Haz+wPeBtpLM8JzhuQpWg8
vmqn7cQjoI0VSsikr+asLwj8/iGwFaCZEFw7QOu/Ec6coEf43tDP6dP6pG/GrnJiUkG7NJLlSXzG
R4Vc26/JUZgZS39h/sTnZfLW8gntOSQah79rRlu+rRIoZ8M5d3YjZSoixrIy4TutrLP6d72VmICn
c5PYB9yaIlGs3xGGzE2L+yFJ8+Pm5mTGnOzyIXzvQj9Ia8e/t3wrtgvnivHAxNuiHgDPpkHFv0ig
pYiMC1Xp9XQ6iCoFJnOB6gWhowhiR3+oAdVjL/CJNaF4xs1QLiVSwvYOq5rAnxCSBrUtClI2xi3Y
jW0oibHmrca9QErBM6sLfgxKgKJkmePvJ2yLX+K9Va88/+ZKwEdXRcMyWVb+GXyUn555we4wZW2a
wfvWX/q4HDMQMabeo6NwBefnqn5k71xEMO3+ROmbukP6jO1b9j9FHSs60zajnhRd7ewPglcB5o1P
HgjgYgn/8NqFE4xj5h6PSesn34YTZ92LWknn/xcsT8rSrzV6wK1MHPN9CAA7ox+m903+7ljwwnyJ
v6KiyaOKudwouDsru8LHuR+hBwkw7YW8QVp8qKhXAqIVYZCo57Qx919A9n8JYvg3XigvRUgS5nRm
IAGM6dn1yndd/Tll9fW0jMKJYdiuKkYwG8u/FOcSesy4HO3Hzf4enE7pXwdysdDhhT8Bh4bOGTi5
qxI7/HbrEVe3nlS/4kbzt+gQkYNmp7HIhCW0HzmwDmrp/slkWKjusPomI2UQZcKCu7+mKMjlWpJl
s7oC/zPvQt1quLyF1DuAFkER32D/BlXTstR+BuoX9vdsE90zbpNcijxzFJkIaKPhwF8xQEreF/Ei
NBucXhQNunlfguTN+bSfA6cmR9zrT/fAul75QLYBCtb1U7zGvFx3fRxe17aCFoYJPw34yftyCEFY
GnuE9m4ISRaYzwJAgjZFdfUitGb+EKxLkqWRajtHg1CjXGY/rCSz/F/66fociXkfeNCokqqP4NT6
iiFJySkqyUDRqlFMOYz/0UMDFHrI0I9yWdODX4MGzyL+P4PKbrM0K0ckvtKOxKlCXXD+lj6ZgEr+
8TmofNRlTALkIrSo83N3644GsEE7QI7w+wQw3VLzkeUtXWhq1A+gNKPm5TePDgYKszbmJSVzPCzi
aAemWYvtRw5Ct33txp66IfkyMmZTHSAZ+zvF+0Q6G5/oNY4M37wmwrE+WczaM2SbIo0gM7Gp9Mcm
BYrWT1TMq31mYUjymexWW7CPLpj2xEVJVQn6r+iKfz5PeJER/Bm+JIGQeqbf/5nQcty2vujU9+YN
MSVD6CixUcJLKxmB0fD1nWkLiCDMq42AZaIMX5s6tshq0Ejgm+2XEHL3RJz6KD8F+YGHJceQrgkW
15/6/G6QmlOtSXv/unuIdXrDRsnzzadag5kREfgeIR6IPaWK17EVgkzLeUSFNl8bTN/AA7fpfypu
JewQq3GW/LEurTiXlr5I3q0xlCRiwiN7JX12edvvplw64Zi9mNaxoXGvM4HW1YagDwdChUplR4LS
PwtxZ7bCM78ac7lOscO4ji8OUlMB28NNYsgIxodinR74GfQZ2ZcBb32Ukhzv1b68OgiJmN3I13TO
TU/WvcLvI8Z50BBfa8ZLkOVg1f9ThDLOWH0EXBpKvSEC53VHfV5uSSUNHheD5vRrivtzSBwXycuV
nQ0ns9yqxzu9a2blG2Wi+kW4tO+O1dFPnrQ/6CoCHOfLKN506casfZn1W+YErZbCXANXOuvtqlD8
suRELR8nvX+JlzR/YaVA3xj8AgrzL1yyw2X0Tq/ON/IUpvBw2u57EFtszjxlPbBkkodRe22bJDV6
InWonRk5OeCEzrniraB7cPj9sY/+WIKkXv3FtgdYWbOeecv31WQADyjr/onS6uCLgetFfSbwJb/g
jmVPI7NysZjY3HaAi9pNR8CGlL37cFo8lQwtzyeVXSmv+TXPATvlsqcdDgyx7rKG4u2l6US3WR8v
tJw125B9xMtec4wqJET3dvLnKvb+0LaMpMcbrfZMol2rInlCGtjCE+NWdbVC4p+PodpioeuMehFI
P+xh+r8oWYu/yu/8OiRmoK0B5e+rrsPrKHHXC2599fIbRy7zB6WBizP/sEfc4hKo1S7xWxesJhfq
st533TDvGfzJ+L0JIs13ECX9F09iKPGgeBEv0XQw+JNpg8uHRj/F3Wrp+c3S1b0/gwpaNUOtKexF
IHdhZw4q3OFykOXdOGsuz8e8O/M+nU2m3EZJ6pLkx3mUftXnD9IUGFTaOaTwtplNS4wCFVmHFjxT
KOgsVd43uTLdd8/E2WJG/ti+4q5JDfBh+JJ5Tuoh5/F/8CDtmWVq5M0EKHsREWUuQWRFFjdQ3Fek
1ruVg7lWHQ+kipDnn3TwnlbcVDtT+9qlWySBt4nOmKEGt4l+OGGqnOW6ooZYAOlkcg8SId10eB29
MJaMh+JxYAm49t0ldD4NAuAv141sjYS7dyxYBGU67ykTnr9Rke/c1s12bdta01/FphfoA2qB8wot
9PwBc9mVpeUiT81tTtwr9n2qboNYkTl6SlKTIr63K80ZT/752172mpsa2J8OvpEB8MO7iO8duAuW
TClDlcOIWPaaYtkE/CjDZqLY/mQvS4fcU6ZBlmbPocVK2X6kD8ut1OL3hQugwjFF6b4mJup8AEJm
93IAjMj4Lkec5tN5CXftQhZ7B2Z+4s/bx/ss3uHoIEaCv8QNgb5ksssuWM3g8KJpmSnW27m7xjxP
ZQfaAvMw6D2JZ8J7960D6bxYxwFjmmTmoI2u1o3TSZU1FBxu9eIGmE4fPOHHi0CKqYUA5cr1P27I
A0DlaVSOQ91e1gMr0b5Y66uuT+yAhnQVQKlSzZWqZfqw4skJr6Uy03PGHN1494zPBoZdPJ1c0BiZ
IcDCSaMi2vW96AYeDgZ7acyhL7RdFp1dORmgC4Y8iHQBBNvjjQfJ2fS3L54tgl9pC/cwmnQi7sgg
uNcG7/antAHw0QLSdf+jkWNjE8Dy2tMlMiFHnwHNWXyO4tQfdf/s1U3NtgkeHmyfYMMiH+QtAL22
XTBG302ytWHWstpxCkqsik0eJVx9b66LdGbOCGX6HZgSJWL1zFkKRgvjmmi8JF/+oVPW5u5sIvri
1fzJBI0dLorZ3Q6czTIl71r71YkdsZmthWSa+j9Si7DGLGzI42xDAXgiSly9CWZWlv9norkNbscW
eVynVuyJmUS1PaArJUElDj1NLBfwhC3OzCTc7np2Igf0Qj/cSzO9nlcdWjy8FaTb3DfMnROv0QeE
a8gw8DFP9l3hCXw3OHGblkEtENZZJg0uTi7ZjiEi1YLC6Vh27m2rkI+UymeEda8zJ8hCa/5AvBy7
G/gjmlQivG6uhsE0NDjluENXRw82LaJlu+4EibCLPJdilkjq0R8cE577QeEvl1/MuK39iKu2NWhG
KdkrR2feYGE1keLRwQ7i/DQu2/Ev3d9lJyOgeXtwfvQVJCDukLvdPGFuvRRfJSU71ysgvSmDlPnq
l6ev7/C47tYbinfoEpnrirPuB3T93tXAy9Jgm4BSTA66esVuoDPY47PFVkgx8Qn5aTsFHRIsEi4Q
8eysN6qoEZo2F1HgNT0/F366u9wxxaEmLm3QySW1jFy23vRHrs40HgKbiPilO91KN9vc7rbi2xgU
S1EpvcdfxWlldOF1JvygdS6hmXcASQBjkcIwBBcOE71Oxoh4sGLn9cIW6nkeHR4G48eyo1gcfb7l
FXToWmywrM49NT0s9gfu/SpPcaROZoK+jTyipSYJuAFnnBvBqCeoZZvkMswcJPPQbKMHDulc5f1f
LcE4saXaAVJUWfKJKjzIA8X2uT3nsCH+eB57AbBwBTCZpDWUvbjPL3SPbB+/hAA4Zu4v0xXRqTdJ
7eBme29eYGdpSaj1FAAm57kIB9yBgHJH5qCD9JvUhC1uXNnOn5rpulXhrgSg9jlsOikav/j/dg2M
Nfn3fPBlgixXdQtqtZjphVDU/9Edk2mASKgwEBvV1fhiOs3WF1KiiirHBKVk0qioc2ajK5c+026m
tbNutToWZ4Hdx+HY5y1gV/txSVCeDlG6AglRy/t0DKKg99p53rUaKBas0QIGSwFbOa9ki3XRRsL4
sGorZ49niFlHcOHXLt0Y1zwg+LeLCpGce0TvfApU8KqLodP2DFkx9ctRUtH5x+utUqliNZdX97xm
1E4qh9LNb9FlLxCJJS250wy8pA+oKm0eevNFnkDEZ2gICdx5AMvqEXECjPyR76AxlfS9R3C20e64
4TV1m+UtejeXug5FmoDIWFCwG2Lsd2souziechSYxzCJrB77vOHLfow5GIO3ZUoRzhDVXPzISNqH
CP5iJuun9To4ep6qb5nwtR8GXmDEzPyLMTTkFUo1Mc2I24C/RZwzkKmigqIcFJCGZH7ddM8jd6rC
DSII/zBYg6IP/2F5lClAQGS1qk9etou0pSTHX304/z5eCGbnIDySKz/vCxboSMPBbc6Ce+kTUntZ
Wxm0d9XMBS2cYZ7H3QLGvlYBsltPIwKbb7++Rv5vfGDCDC6MeajfKbHlUnM0Wz+jTip+8txddNbm
jE4rXkbAV1V/Kouq9JqfB8HUjB/bCFPrLs94Fgc9p/t0EQ8Bv57PHKT+yA/sgxnArR/ARl94wiAJ
LRE8i6w1BweM9G9OO6OCJ0DzsBBl+XatGQsHUm1A812LlLVCd/6iWmNLN82FtaiaH742CBn/Y57q
UroHvY+Wz1Wd69PXhBFf9p45p+bGWRAcHTUwrUkH60akQpDDyTOKyRlXn12jJRv418vqKr860wnh
AT3q9hmXY3dkzYN1fUtGSHrmaN7MBuGopbnDFKJerP963Hs8+p4np6wwnHpJEI9jzS3C0uaaF2sA
IpMayMZyKnX341fuL9SaYmkKajFIVfH4mrVe9ZvkjHmodfFQGtRyTFMZr+AUeUb9NBN/zIGh4PoB
iWkbCJkAtfd57J+cjur5AERwNR5js6qy6cF/GN1nuiYTKfDFMT2b3pK7Jc8cy9XgFoYsR+1AtZgM
OdbYUCQNnjuRZ9bJREQ9EBnM8TUqLwmBAR+CtNEQMiupitSvx/RJISTpR1Ih23wfUZB2d4C1wtND
bUOashMBlHm7wmpsi91fIYYPWz5P3aInJSBOl2opoi/Q1Id7xqVsaxOd+GJBpPE4kLtnSpmBIF7o
wG25x/6QtnTNCLSqXRuWEjGM0ateUzOj/6ImPOTS/n+TTROzJvHpBGB3oNZHouxKdI6Jx+bpKDIB
wRLkonGC1wqtjfbxc6Fr+jyL7vsOKIpIFJXH3kNvwdN1SPtrKhXpPgqUr+xKux4Vkq9yyVTq9JIc
sxWsCr8y2TSm4Z3mgFuIK6AyQlizCeYWUHta+FFHnE5er4Ixt0t0sh9eD5Gf4NAI7WwgJ7do9nut
zNX3GXbjHDzVYVXcX4YVqbRh/XjI4fNUspepju993W2Zzk5LCMB4btCCPoGGQAp8twVPA/OT7wcC
oamD5Y7Scnvj1UfMRD0X47BqUv590Z7rbF2+noROdnWqpn+/lsyArsmJBmhNylo8l4JEEMLUq0NE
oHzML4rUxEQqhzcYBZaY42efwONrd7cf0mgiugNpA8RwRbxgYVew85JVhN8xtqqSteEKqUTz6uN3
qjfWDQ6kRVEYbQkAzGXTdGxRGpP8tNcqxcBovLF2Ud4BR6mmtu02eAx0vo4LwLqeSOPsVQh8bweW
RvJawGg9GIzsYjrZcMbdJqtM+a8ykWQvZ3Dx8Cz//g2uBYDPqSsPf/peS8C4IzJOs7Mwfl7U0ZEk
wfJ7fqdXOcIW1UHZgHSilhh4gzSa3IQLodd1pmGksPqMOBT3fQbMODcRhBRelYmpsUX8FTGIee52
Bx7Qj5FC6u6JfjIhlK03Mvr4pRaG+b8vbbSV3SXSnoGauLTw+ceDPpdcZNwv95xRk/NzsaU5ZHsZ
BLhvBix/1Vy53lCYJulovrln7MpDHr7IHP3e45uxYhBjv7IPcp9PV3pQEH4DyqP1nh1AaXtT+McL
V5AfFbWh1tifSM4nwzQsgcCPY9Y8K1ZyxypvnOEvqQu9LQwGUrSDPLltbeyfGfBBdw4wpFS3qNO2
VDgpe38DM2znazc+g+HlMiT9XB/ohjicdMViqbM/abmvNFnhMmad2vJsWHiIIy1FpamVR5t3Iwnv
Tf00+otZg5Skx4n3jfafjhFiQ3SCciHBJdu49+rewzwgIvS846/35x1Eli+malNfAnEYhnaAnJ0+
b89shW4WA+ExByWroFCEvOTDbYmumtA2J3QvYvldzJYl51L5pycIEBGLPlXXnBKZgbXsagiKpa2E
a/bAtX/SLZ0jR+43v5R4DVbANuNZj/NL09gdzxjqeBhXU+nS91o5iIgh69QtPXUC1zFxnpyL781G
lxU6+rW/Eb51f6fgaEEmmy1CN/yfRoEOBbRVKnwHQdv3VUF33l9LvCmJOeJPPep5WGiQXX2gr4o1
+QwcIcZyjsPnONKJD9ce8Wo2yDKOolEfw2F905nEdnmJcuueii+ak550sSc4kn3EEwErcaC7yAoQ
u8SncCEJDTQTHODDyx04qtmfOMHEALx3HY//m0xmh0vVEunoV1rV64L83uR8er7M5jRU4ORtQ/Tv
XhbayEgSZecTNpmu0afzQQa6HdaPpLLLIE9n9t+yvsaGyWf3e2zqbLs7r+GvaYuK6ZhZg+CxtU6g
uFyN2brM2sotEQv/BvLFWlkrIy85gDSPkzjFZzq39vyb7xay2c8P/WU87J26Tyq8rcq6KmvcrV/a
oaU4BCRT0c5cJde2t8ZZmFNTjOXBRw99l9GheLENfSTntGdLPtqySU/APquVD3cYVYjSmaWEMcUt
3R6JcifLIjtuGJqBufl8EswjlXVFMyK3in8kBkaicnAA1Uwrytnam6zSL/7XJhlDXaqivMgqyVJQ
N2QAx1WzIsNWM6QHKI1blbGQKzZ2pLaarp0pGRCfGiguizO0N8iCABwj2rrq/8e2yZ7/iwDIK365
zCf4dg/jHmDw7rRosdk5B5Fep9X/FXN4G+UeiA3n1+zU2Oes1oZOuYs1ul/bH19s3Z2OelyYX3vc
pKrzdvfRpnC4FT/P09rfmpRcbr3XMziO96IR12pKgAwwia9BGzU9IkyscDmrzM03505R4XjwC/zD
XD5L5Kh5bO5mlaXmSV1pd+Acx80wFCpOg5LEJN3TGAq5Vt55nxTBhbYQKmTOmE+W5xuGCUft7A4B
dKbDB/nr7/WBlnHSjV3WSvrTuc19eke6zYNgmrz5MoHbIdS33Pz66/N8PHnLUxW7g5ZDGbtfY1Qf
Q/gnCQWm1ayKbBMJw7PlO7ZPen15LZQwNTskjJSUQUMMcCz3p6GPDZPyaDyrZiv2aajSaFCkenmv
jvAcdMKKypH2ykkJznHeeXyaBcbAeamMuXAULiHMaYEPvMZvpC1At/lfeQqU0UcAPwgp23/2To67
/h654j1MYumZA3vA7XctJ74He3RBzzoviY72xIWkS9EQx+zCNcdIK8VfLvjEBj5Osxp+0M/CLKjW
hDpllYRxyt+16InmkdgOlyjg4nlX9APiHLIlvGm6c6L6P62hPZssdfE/hwlOxMbVl3qp0EP/W8kx
tpjdffCj6ZGWwY3sI4O8euqZ42cpav3w24gsUKuAtkcQKXjBBmk3t4MkSZAthws7siduwwWwDbgf
lOpfpfbEQpjvXETgRuEm1HmtUVo9uI7j16ANROrANxXV+0FzUFE6VfYh0MlmjZkrcseYa9D02DrJ
U49ubyIkbyhq/Kz7ZcrHn2gRIC0+aS+qiLyMVpEHaFTqwOiiOGf+5pR2za1JOt2hbBadvin9K1ln
4EB/c3aDyZOardapkCF8DdqAc9J1c/L4y/VTvOMkRVH6mi7ZU09p+noTI40i5i4NCdJtmY0rA2Kd
7TPJq/k1CEgJZ51nFnocieCJmMvK3grB3nbigGldCY1vfZqLyDmfIVjXYzs6YGP61HJCDDSS4Er4
gJT8QkRD6axO/pIsZ8COfUBHhNPgJnzRdy3d0gJEj7hLaiqMJKGQ3JAkGpfdKXrTmxyU0BQ1Kx3x
vV9YktG0bJjHFH2SkwrThtu4mDydf3P+tsqVCJbSjqItHj1nmKSiHyVSWaAltd+6KRPC/vfMLp+6
J1+byfFAc4n3BoKEVmrbLnp4my6GdT8baeh0ipRnmWYGyFHUqnrxxH4GZNV8FXefu/JX/n10B490
dru0xIrQwcbLxIvLiQcWlgGnnK9dF/xR92t6wfw/gsEJEhcsdXZ8V9LKFik3L0KY8tmLZ+y677c9
2mw/UFEHB0BDBjg2DR9ABeLuewyw8XKZa4LN9ZRCRkO1otMg1yS6VXD9ZfVsIn+43j9kZ2AWjkaS
Bq5Ia59q9lV3aLQ7CXTKsqyiNv2Wotgo8B39wwML9yrt2xWIeBaiBkbF+zzSrCOEBQJtwp4ysSRP
MERQ3KB6wlrPCVBcmtG4O6D/ge40Z5dy8OvfOVs62iZk+LGRKz1NL8e7iR3x9Yb44Yt6TKGeXoTR
qx2lrCV1ML8O2NV3ANWRMDTjxsiQe40PveOdOa5m61tu6xvz4mHG8zLQwK2Spksee4SLot14Xomy
NqXA3Zo3WLOuii1UWSJiBvlpCmShOTPyIsSQRcZuI0STtITHw1TcOSkuWd/Jzf9nzshz6lQ2pDCF
XlY5TwmrW/rn3pvM3efUauQlxazs2kGdHt+AKv6zpkXTx81iKyoV+e66PB0VxVNgulilG06aW9rO
qbaLUuHdLHaj8ftnIo+lKqcb7R2XMWdAaWMQ0lpQsbfy3+igTs0nUwYDWoGOfqCWJr7tRCymvXW3
a+xiYoZyQawoN7guS9oGv2//A0KDKbqIuSwrXB8AlSfr08362FzS2FLnyaZzHQFWv+BQQG+GR4CY
Mb7hyUUBUmlSb625C1gsMfE8zYuzGtmdPgJAjSOhT3MUNgixphvP27QlaqrNbSd90LC2nZdafWt/
GYH1WvsnQf45rz+lnn/1G/pVdwkxup2ymD7VJwSdqvuI3EToVXfjuAeTq7YdkMS4HAfQUgSJmMt+
Dh/E9p2+px4tT7D6a3ukFQhRe5p8cDmkotB3moyebMcjxpFoCgEBPxt+WMpSdeU7lDC0UU6RPPMo
DhhxUxNMWKnROg/dG77G6O2wW+AAtEkIDeyUUGafAaxM2OpCW5TgNrVRqcMAVXHDFoP1ONINcHiO
xujRkBg5Qmxbe/unkWaxmE7DdHYoqFpLGFtwKIFXT08j7/oQQz98WzJIJ0XIMPJNWohQfqVINs/g
yFocWhajQNZCxBd8lYT03PXFV1d5GZN9ECbzdEUT/5xUP6PURwlxIsiNIId+AJFrt+tKmq663n8B
oP6gENaPhtxzkMg0Q0nJ8cweKJ2dmITO/VzWyu6oHTz8GvH9E2w718pncOIT2uVeeOAyFyA4BwbE
6aMj4+c/sIPNLbh/QMHElqxVawx8/fQe8PHiN8Yud29FjiAJye9xtQ+STAZdUqGIF87hMr7XP2B3
Z+y/FJFAqK4F3oNrlqHXqIhGmsE2kFMUXECIZZKmzykB5A1/2IThWDdQO+eyXbrzS1XSDfZEOpBb
Y2+D0TNINMlRoQ4ZOmmp7es6a+eX3How4zzaORasxDSYKJgJgZ1iCIlWkGR5EV5mhUTBXJ0DThD7
nPmjoo+23rXEEcaSC3Mxaz7lXqOhMJke2/fumdTuyjDuS1o7cfpWNKjV0JjkPlLkFxeljZAd7BLY
GdsyJ58q/3PkyE0OCFVucSvsjtLX69lnwugwclvVEWv3yxT3WGXhLC61z73rsr7AD1XiijjkrT0Y
Ag7HEdj7N75grPquWuawXk1y6GP8WKcuhBWb97Jvh7pgriK0ze09Dxc7nyM5F3DgptQLWTf0V1dA
EQ5HdL6N6cuieJ2pRIP1XaGK/+RO8i9Fx8rbfI7dsmZIABg46X5btMaEMnbm9MATrJdRo25QD8QH
a7E7hy+VhbfSr+OA+9dIXD7g7FVyi2qLH2zUcwu+KV22CT9v7A5/ROCJ+tX/tQE5Gx//9Pv0z2sl
96eJ8FDrsIWKCQwhYcGCue/E9x+IoCIZI/2C9oMWRITOS/qli+DXMtEZIIIByK/MRYK5R9PybH3A
8vxQyLjeJ1kpPFftIwtJ83tueI28llvl18cPH4V38KJzkGCdv/CY/nqMncbmxro/c32tx8BqSHWF
92hAwqw9nQ+jQ7oOPvkNMcQtZhuT8NnmS0I9dcCoYQG7uSN+1WY2BHd4SmRjvSjNq+e6gOkNYiIl
kmutew51+LheJHC7gCQZKSUDD93PdkiJ5p4Pa1Js6FRtBDG3m2ZVGY/0t/v8VMtWpnxhZGGkfo0z
/R6Fp4RHN6KLOVQP3hXcJYzTMotphYX2lEDfqX40OQvGytHMkXc4EoECh3Wbsf+gEzcCzlokGQzH
kAL/vUenBjPUZ+CeJbnDvXziNsiMVwMkaMYkq3L2pDvjNuhsHkr57A9FYRE3s0tWN7EhCNgDcXWb
a075k92VkQZ2O5xMlgWMEVkAkq2wFGfW58HkHrRCxSzS1aJ5GjiiW3nA8e2iGiOre4/tqMZcChI9
eouwNyTejT81BhslAXyfiUNh1psdR0N+fIEbN/NlvZIwP77+sSKoYypWJBlcUJUKVpbSkIq6EVAK
OqpjK11acUg39MSoN1Y8rm1JMrKVwcdVOYAOXNWJD9BHsRtq++zQdKm5+VC0APtT5p3wCSsuxKCU
KmJpAuLYshqbwBn207JVyLPQI6GxvW+8mO1kv7mozNNZgj3haJaKMDJ2Vs+93j4t51CXgC3sSZR2
gWDPUWZJ8NiXyi6AL02db0CC0mS2HJn3XkKmo2Kz3gQk3wwC9UB6b3l/vcNSVP4nNb3TnN1UwcXI
sPf085HZfLy66X407UVUoUqjjrAbkozdNn23NjOvpHMk1v/fErpnvXui+5Nogkbz70B0mj9YpXcz
W7WVbPb8MOf1f8v9zQBgIY2ImUGYmMz4HslnC3iaSl52FIdxmxTfdlcxmNozBNhuDyrd7MDPESH/
YJhiM2jVEAoIS7JJbKgPM5V76A1WiOJCYip5eBAC0Rw8Sc5VYJ6QPWeZL/HTqD/HXOUU7S5x6M96
M6HhG/p7IBFK5HcvU5B+wNJpTpCdMzZBNVFzucP7AtK6/TCKWrUursb8hm7YGRBV8/37EcCtVGdq
osWkJ+j+JBF3CQxU60WfpgWFcuWnCUgp2w8iWxbb78KieoIXGA9nMocMvYu4WD47EKFuEG8mS3Yr
EP+tF4TVG6ztLnUkNbKXk/BYo+nhlXQgeHKsS3wUeFUOlyLMXBGCPAZ1YPtqgF0D9OJqFYPgyqwe
FqxeGDGqTyovepxmsoY04K4qLGTWpWxDw5Zgas6AzLzyyPyZunmZDqkiRCGYnpobMojzlPJXYcJH
/MmsJXFB10WQNsy4PpoDSyi6fLcqpKA8mXAKozcCC1uopqljLbTA1R9O5mzdLlvykIILmpPnKeGJ
LC9os2CG1V/9KnQrBrNMSFAeshputcMO+fVVaGNAIkVrPLOmKEVbaXPRWakSv/EQ8NS5YBNXvTIJ
rdm6A5+vWGnTepUKDf4RhFaDpN/MmM/FH3XaQL55i+L6T6X1DZM6DcR1jp/Ll/0w2RmmYrt24vdR
RM+pXI+tOE8TvSGNBMDpVcq3uW+2eUs/hjTavm7AALdmhTsZbF1MqBwkM/pSJqmlVbq0lWbtaMT5
7vWh+HJmNFp86J2VHQEg4Qc7ntJ9Q9fwEb524uFfL/xHuG1iMpcBsFGyacEwpxCocE5fgojx2Z7m
iA/AkkNdr93gm6Q94qk3NqyXNwlYtDVfXwtL1HUfKO41o1+Yx39nQgyHFCbtdIBasw36gvxBRv0d
XnHBGj7t2UR/i1L6ICeFdVlX1oUlnbrh3IrZer5+y6dFV9iO2CDwHomWs2oDoJpUVEIr4fqZ0tul
6vK4mPsajujoXZIrq6fAdvKJizYmj8Ge5ytk7l/kUCeYKDu0O0zhUwHE5JiRIceFWIndtvlWgT/G
ofl2zVshxWhUD1TSfIWhPGMLrG4qW/WS2T8pX61e+gYuD90RHy+M0PLJxmhEf1+r6eGMVkSTca1S
6IL3jjjknZmO99fXTUFJV65G62ocSIhxav/aMHh++gcl5IlLEtcAsRjR8nLi0LUcTaV2Q/qcanDq
QW2iL6ljrgtAD5c3r30FHQNNBIdWgKXoz40kG+6c0pmm/YrQj6hA+bFIP3hf81LktfrWWpSkUz1Z
VGzAPHqu9Uoof1mE4NSUTomMSpdZMM+PxoFuZEkiSswCyQftD4CZkRWNoXhITp6Bw+NsM74sPm6P
aasoNaN2XTnEVQhtT2XMQKSmjyUmpGpZpgE6lKRzm73fbRL5YgkQX+xwxViuSujIcm48r+WtvAoH
MNblMy0VjtFx8NmnlJsPifb1hS7ejNFplN0tmZZQNfjs5RVa3EGpkP+1jvT11gwoO+hyvwhTNjYE
N5pN3vKcxuiTBfkNF2jPKm0e0b53H/Q9gi8+gSwGXFwuaWtYIfbV1HFSDQiKaAU1CsGuSAxXSqS1
CbEoQA+Ad+O0TJrUdf3mDpswkgx+kDW8/fLBduZuK0OUx8coNibJoaCwVzQa7nLktH5xhmlRV9gD
1MmrWkzlCjqC7DPbU6hCGXiHknDVtytBGaYf5MqS6Tpa3XQtDOw+cyBylCHth5Q5aH4X37pAyeW4
QqvH8rMWuP7xbibYkVPej4FogiP63HxEdC5rr8z7ekOgrFUVi09yVVbMKHbO0bKEmDrqu81fK7dS
xJJEohH9pIVT1MoCS5oEnxEJCFhce+4gYA5tAzwd4SIaGblf8I4B6P5KWXAD5g8q/5xmRmUJEMfZ
mvdv2kPZjyisYPkAx1ftCxptvIHMHmZvcmBrPry95QTu14+XjW8bFgy1OyONS6q9r0Jz24gZq6JZ
jMEgD+rn5WI/9P5bgqTBPWjMQ/43Y8pgNqlA9DlSBS0P9tf5EDIUsUU9vL5W9AZ98sLgIPs2PEDQ
yG9HkNg2PxKGKoWvEO0sNWcWyDKZTnCrcfWFYLLQnl5GjVg3BXPuH1pQjrUOj/AJurugq+BuFg40
IHA3jxrrf5ZSUbNefW4C4bTumCOX7OXWEDnPE22FY0LGoRplFP7jaPdlACOHWlCxNpr3pXHz61Mt
Tws71+fuXBHunPD5uSLPtmge/MynoPb7X58+cy/ObZNwAYIvAK8yBt2GtfOom7zOe8lSnCf1RFcd
7LluO2XVnYElxZYQxBq30He/lP0p/3A7cq2ZHhf8oTaz6w0hagRNPQw9Lj4oPeG+n2GHGyD0In2u
jENkhLB2g5e0IT5NmNtuuAxOlgqnNyLcr3jnXjr3hWiadZ4brXxGoNFf5qzms6o+wqQZJtOVV4Qg
RdkzbYtpeZn/MjOq3iesqMfAiy5a2ro20I5sNbQmwy8xmQ/eM1uwFwi8jq1wmmt+YPYNvFO1JBDN
8cftwB05v55qdIt/DnsbsR8HLUCKuziGvGHu8qyx9gTJVQO15hG1T3RYqPSKxIeXl1+EKVwdZd8j
Moh8GDgqNuHN49zXsn57KBBcLywT6vOCO3Yge75CH+xrfFbnDlzhCSpC6ZjvNTlyyr6H8+XxCTj9
sXL/SWR9MfGNaB7kGeoLpLwqR8ZcH1iPNksnNkx5C286Ep+XCwX/CglkfBVOcvt67vuYNwcKxhnM
Podvsq8Uh8Ljb3KrAJKKUOBSNRD6aJDMvEDmE8Q1r75H9LBctQHmqtwUG+GcI165pnWC1DYSgrdU
5eQnmsdC3ytBbNDha1ZCr8hMs61S57QQU5P6bDnKev/S47CZ3QCJO7Ue85tYbMkZtU5vkFjRyOVY
evtml2E0fZze2w5iCJwAXRh2Si7WHm1LzhRHwzIMupCb6ZuAxxUqUmAkg3YwrKPv3Fvfzq6GCkLK
LMGY6Cp1wdXY+G3xgZ+bEMwtjsu7zE1+0Tv9vDubUpVafrO0+dhwu5UmEe5IZkhUhtiehz+4jnLF
Z0vxaaf6zXO7bMuyfmsIpgadj7T1vrnSJa7PHrMvjriaQlZz3xqe3viT+O6qMupK9UDpXAAezau2
QaJqo6vqupn/OYwC7Pxo2lIdX6qV/hcVSTp2bo4ktDenpOyJnkXiHq0WA39LcQolKSkHmnFR/dVM
0NIxGzfTqY/BKUpSLzW+wz0GqH7FiOAA+LMfIsGfqaxdAwm8jDGuOGWqFAYZno+x10YMjTY6z+Iy
bLANueMV1Niv+o3OGrgrWvJF1ZGfqKpHoj8jkEU0X902w5h10WozB1fpFRzNWC+Uh/EELqAH7y7g
dyHwUC36fx2L3QShs464jGhCFVMva7e9/tOwPeZbeJUSOoprKtmn/Mh0bH/2YNsSzwL/asYXnlZz
jnQOtqiYQO922uD35+0zmG2b2+shaQ/Fu0vZtVF78+bPbw1zcD3+NYariTizQFCsgDTehgpb7fuA
R0LwLQTH+D44Xys4T84Zi7KWUMetJwURmZ5vLWx/noNtE5r1NDl0XY0Yrcvn3CwOjJbR1x1t2Ls7
okFK7YwTZx9xBimaZ8HnVvZMM9XL0r08RpZZOtUhiuvjtqtOSUcRn97WRqa+u906U/5r1nMb7au8
VfaGSJ2IgOR6/MwaUEYKlSw3JR/3/vEQ5X85Y0zEPzkhfquCbI5IC2gHn1e6JKpZjDaTXPE0v7sR
pHTsBFOflJhjdsAfo1nJmy3kmddblKF89/mIXl0SrR4FwQn3JmpFktpwSGIEF+JwLFujzQDpdfkZ
ozU06zYdrv3fRD13QkL8fUi2Log2NF46utOoJyymMBjbEXne8bKEhxhQLdw+OOL12ohNi1fk/eHB
cwX4xGzhTokJ3HCUSuo0OYITqs9j3LtT+ADORWJzEeadJ+4/yBYDM96PH/1yzCJAtSONw06zMHgy
scoiIOWxvAwV9bJbY74qz7h0V55Jvr+pwzN5coEVcpxbV8dWDQJMA/6BHNlM8WyTTCf/HDDrNyPn
BJvIYWFXAMe7x6IRFw3TBT+EvzURnIRH6sib5cjzKHSPAdFwQkxa50T5bmjiW/N/WXElGrAUQ7Md
KWgc0Ht71+oh+2G/tVS9njDR2sMFePCvEFWtA4kgjN/YlKAzaUu+1fJ/K+2E03ecXeckRjjnLR/Y
bDVZtIIT5bBQ0/jf/w9fpplLKOU6MrER5i57xss+yGuONa6/+z5wt63Ojwg1jS/3aenGu6fhgxkW
I91DoOPzfzsuwOhsnozAyJMfu9kV881kYcmVLnL1rG8W5Z08mVSNOJI5NG070O+4EOuuYdeXBFmv
uxBE60ALeccP3Io0ZboM8MdRuCG8aHLLNGoacebWH6wpwhcjJmvMy2+t5l+F1BlRiNYWDDXwgFFG
cXK2QvmSRSp3XigVYYFdewOBO78Q+r/z2hYiK3Oh1nYXG491LW+ysO0VlfW/DU9/olKlDkKBc/JJ
4SXm84DfkQvxzugP8tdX5+avcP90y0glOebOlg+Ma5yNrOGlpViX32Bi+R8IMbQNuTz397Gwy8ek
E4kV+tEEczoiieshJbQVwWWpDR5i6X0FVsPvissWfoZoW9f5u+hLoBntzkrTWFkzT1BEcVRu82Qd
XbzmHlhIF5tuURAZ1f6oEB1Og0ZkTY6fj18tFI8WoJs0/s9GYmbI4h8XfXrgSrBkyXsy159HftJm
w0JZ2QpgnCuKQEhGfj0TrbRneQWNThjdDe5NQQ5Oor3XDTmy7geszjf9kvBoRdAK/Tof2l3L9DSN
/dtHATFAC/EqY8pSPBUlKZsryKPwXxWaLEVA8o9+Snlq0QwQqwBnqY/H7ILxVHUjdf/pRJEKFIii
TtModGBJzyqUJf5P+5WT1rqm/jDaFx10NkpIBjEnzU9Ckccc662yt99J4KETk/yy1exzkKl056S/
vPh5+zvW4S0y2TW88+CGc3urF2SSzmwWveuGjsFenCAu0x4z+3qV99Zw1qkWHgFxX3P6/7fVU0lw
35sHEIliSKvZpaB4HBs2L7SyKCRaoZQKBQr9iMcnv7QrMi90sGrRA8a8p+AMbBHyAgbC5GOArxY7
spM8DYwrWxq1dKfcTHa3lwiARnklRN4jK11NkDRs6+joP1IBk0E1BZfCL6JVX6Ay+K8fZM4UdGRw
cGdCn1V+HBQt73u6s8uIpCcG7O7B2qkUSZjxR0PDhLUpOfs7Ad5n31wLrrJSlN6ugl4qL5AfW/Ht
pmyBRWLfw8fdO0KDiw+2wajlt4d1nXYiD20eb87gRtXfX7qmDpgSpBRUtvo1P+F9LnXkB1gJ2bRS
UpUZw4SqJAHynRD+kCgBzP5fVNqTB2w6Vp5ba983LHBE4X2MQQun87FSQis5pTVk7hRVOJoUge+l
DEjz3bB8gmzyq2fwMNrNb7NpGrudtgrTm5SfHGgbYR5OW2gDo0zRb1LV0UIXQASQx6niY9AAMEkw
vFjCkOa51DLztuhFVW6H01PoGLWO0a1gmgh89asv07VpFpS8fGsReU7IizCjGj5udetjHxHWX9OB
M0N0Bi0xDfyZtJRzurIz6Knz5r1wWD3Y+aXhT99MElUTdCDdEYNjR5sBM/IJlFt67MImxnpMCwGt
HcC1IoSmQOiO/3YYjVBpz4kr2PAY/UBaL80xjunfTlYVjW0GCbKTR9CbtD9P45gxGvgURnpYLroi
Kn+m1v7CZLJZBJE+X7GKJd/4x5Y6u1F4jyLFwvGgw1RmZRd5KTCX3EzAs/CkuOh8c069K+8I1Rsn
wcCykhDE2Jt/vRN00+4sda0lEy7DMwkjxxcyMQJhI9ZTboTh++bJmnf4hPJo5z+o6UPifVUra505
1pf6agpNDaK90xF1FK4R+P+YFacY5fIyYhI4r+gFQAO3RyeatpJCUvOXQCQ9SDYm63VEWeMtgjAW
oyfHRJ+yU8pN+qgMb7Y6CuzorIit3QndGeZ707gjqQoepQZ61aECU8gxgVThHywMoV1QIeTyHwA4
RHhxksjYgShRENLslBYjdHoXJHA/2WoFV92oUF8rK+KfyNehBt8iXQf5nd4tUEb3pEgUP3qhbzka
KuAlzkNIE8jGB2NOqWe1Wq8dVDGqUby0afAatXfbbcfC9Lu1WfXt6NZnBJzGNM2HsiZszElkGd80
sopzOL8vz2QDruAKPfM9gyZOg73rbA7fK72QHtawChJsoaKVue2uD2eVHfdbEXEvHntYtXNMyUCM
jSYS5HbJqRsXq9hlhHLnKWCWB0MlrCZjm9z2LauL1c21AGtpY9IT9XuIjjeA9RWTFKB1yimwSvrg
MFpwMHejAT9oCX9wF0HRrEdPgCt8Gq9p2L92lzPwSmlPUN41idc4X7OPaKE6Td4QyoBtWOWUt/hU
/jkIEOZQVnh9epr9MmTeIIab9rLwEE2+XpBtgnsbLyEyR7O6/QAh6bfp3woTZahECv+/3JQMX4I+
N1FOCm9wVfxvuFbIiZO/sYMdrWwoi8DdBkjEkSxyfBs+1WuGc6f0LfbikwBuoYObPkjQCV7ANpst
ea9sUEYZsNCbkvdWU1kQDpeSdPsDEJuZuWeskj9QUr1iKrO49c99iOB325rmYDWSWnYjXhjVc/ZA
VZkobTeLFwAiD6XlEdwjDG8IrtsNacOVdeUofNj+2x+t1kzPaoZQLN9bBVrmCMq0+xPb5J6uZdEs
J7SSknRcDqxSE7BTQBnj76PGs7kb1oCuNkaqDwBg8/JjaNlqa0V/0Uu6DIiDB0TmVPp3guPkuwcV
KyE/y5mXwAh3ZHg4GFzNsGTP1nresnzcjuJEnih6XWCyCnhU/6DA9X9s7pxPxGy9LLIi6KpdzCWc
50V1NXLOVKKYAYw+qg0HaGQLvZ7gEHdbINqhffxITk1MDXEtq+LGmGipvPAlA5+tnui63bvWzJI4
Vw1LS9zNDsf4mDTqH/Gzk3JZFhoeF/wGwGPcFsnAZ9tCJuohe4Y74dJwApURavO0y3NfZjIbA/Ir
jHmMVPkI6GBZtayB42CyQcNUhH51Je6bveFPKt4MVZjs2tQu3flglBy8YJDz6qp5hYBbcIcXugjT
YkZEDz8TAXZZDgzgfXjyQm+j/cUhbq3ChzsWZC3I2tvpLbTTKDTaFxaEd6mhwLFcOypFdSrjewum
BWeKUH+6+vJM7nJFf8Aw2C98CCI/RCoT87suohWlPXe52fTI85c/erfe1uka4HIV3H6fM+TbyA/n
jXFG9/bIeNTs1gFat3YygFq6xVCrFfXNqG8WFBYhBSoC7K8mxzqUZPSGWK4SA6RaNtLlti907zO0
ttnGj/RrMZXt4Ct906cmzzQD/ziH8v4U9/tSDsgQ1P5tcOPLJYPesCVKI+O/ngFhedYYBZHPhH73
ICO94afhCdxegHq/kSgx+bDTVcm9aulgi3WWU/KIQetn2TKwl2CF6GM+jllzGKxk4eAxjmNDQN1D
TT67T+cd2WVRt8Cy8PF8uPbIzd5M+9fIDE00WuPAq6P9wcD39D50/4ZKlyCNaARlSd6iuJ9UdLkf
rfdqf5Sto5ujNUtxS20sCuybO4uyrYoXYvm7RQYJJ885J/cMc7fsy6fiCAuoxlZg0YnD3Mt3zxaM
Osg12Tczeg8cmiW+AFRvoukfl4S+p5zmT6gzQfyWZDrYIMOBdT01o9zl3+JFA9htvu5IuFCc6Lqb
wKK0vy9+pXlrp1KLseCu6sMDloLrlWKGsBKerz2Oti+TR35z/dFgEPLuDhiHifrurhfBseWATGT4
ynzpPhFUrQgzM8O14I9QKNmw3tqr82j9ZuOzn7NalFVyjL7OY4zFRGruHqCDgBMF1+Hf37H9LtXH
LSvBtzQUUjF5Bu/BLZSLkwXN8hwDONI9wm3kWF0ps347b93xdotPv8RS7yAVcaTP5puYvNOznsT5
6AgfRtREidznmJHRC4oIbXKrMaOeo0tojhbEgBRhqElowPSZGs81k+FBUzvgU5p8hCMoeilOyub6
Ot4Alhv5M9BJHvOZJzSq6ap7vR9c5b5wzirt5LwzHb+nIK4O2d9mEzc0dQxwIuGGiGCZjvvIwfHY
ffhIxO8HYFr5ulCVRFZki1cRUCC3LdfXKBAgIizsqBmUmX6YnbCnPoK1ZkM0o44t/oVPg4y67CAQ
O8lpR1FDWuwwkTjE8y7k088aJ8ttgx8aiEiY4mqLSc+ue5kWMyJrfPXiS9Kg54q46uw62YJMkDIe
/ZN1Oz9DF6ZDNkeNne9y+WFBdA14F9C6fusRY6IpYGW/wmO568Wa24vn+W1ZiNTRLz5N3EYNIMFp
HmcItyxgd0P4JapAoiZV/gx+sD+3iDdZYQ/DdSapFqZf003usH3TIk+TcdDwhxeETa1BH4fvLaHE
DWzGAcOO0Ulu+KXAbYS6j5OQB7qqepsshVBwKBP9YKI7huGx2CW+hK0T3MHErs9WTRt0r7kmeHzf
3v5Y7n8Fw0vCPPkcW2bjRBfHty5B62xvxkCx4KJzgqGu9UMSH8pe/oryOR5prqMx0ZbA6PBTe3AK
cgzXk809s5YuxcjMYdckdl2y8y4qQRfdmHEcY+mI6hZ1F2myXf0mrK7W25TWaVNtAFvlro1LVQlC
48bpQRXAnp1jpq5t8ldxilJyUmAI+6DWOv14pH3Gxc/rmkRRcMX18D2GcifjIJyAA03RSojO2MkR
EX4N42ILPEicLFHauykt3St8/ylM/Y6URQsGGQivycuNuNsfm5KGj7ACIbbFHF88pohgNMphYyaC
kxdCptzBXrFcryfZGIl3+6XAd0KUfOrDAdkld6DUwrBZyKgcPMLLqt+jxx0jubN1uJ3TydsSBwOR
oS1M1LaxhAcoFBdfezULEVRiW6EqVwAxQUXMuKcs1VoK/tBSvQ87IC7XTAeR4LqvebsmquFsT3XY
jHgnAhcme421tZ20MvzRVTqTILPFQvLlpaXY28eg9vZ5Lsk5GdaGyVgrvSzxVK2sKgqyi3hJpQqa
jkPqd2RsOv/ai2OPqeyHu6Wh/nekJpoMQOEoqSl6xHofXlNwJEq+h2lzZFr34DadiAmp/JdLh8yO
20gbq7lHXEvaZGGHAK+IxHWyGhr1mDQDv2RXe00z2hmwee+V2MXqUwG/v4ezmU1hbgywOXAieoZT
ngXFdbfNCPMw9wLAAQHbCrzRAYZ5TyYDssCBd9lWUeRFmMnEJqJpvE3zbYKkiR+gKgspGQxo0Lco
WbtH26kVu7EtBEbnc85UJzk7Rr0ZsF+0a9fddPbAXFxcqYc45YsPJNbhQD2j2Bzz5NSGZ2+IayYW
nzv1265eLwf+9jQzG+fi7JMMXFzbIgcKparJt6RnBBC4lC32vnshxvqVYq+hW3k9Qmm21DtCDsXu
tUFfetneiYkWWBG15yMVLqBrES0S1dcaDKf5fahiNlENgtl7swpIbPOP4JK+BB220YgguMHFWm4C
0Nksgpwmg8AO+YH+gSisBlDIBNyzV7m9ObhrtANTpeLV379/8L2xCvxqzJ+e2+wqyoahAg9VmWOL
tNKWTatdltF4AXI9tzq4ESWPUia+ty0RnugsWy/jEj0h7REOnBwH2eTGJDqoVIJUfKB7KJhfIvBD
qdG8KL0E5VYJvsA2bxJtu0iXewcVGUjJULhUCNL3M5BKlcGiwm3OGvC6BqpFpkA+pQQGfgOVC1Oc
w1TCJgHRuzg01ctSA5VunlBGKmg9a3gj5VjwrLTlOhG1mren9gdyG3zcBf71S0VsKAsFczo7iv5f
dvl7l0H0ye33A1c9bLpCZyNBGso6fe+NwNyf/AosazOT9At0su47d1kD4SqJfuSJpXN+sYRakzXE
piCyFoNRTsGCAFUaJ3btZnYjbKBssYxi8Ii7n9qmE9M/5K5GjHgD+W+xdS4040LO5HkhFpvat9u8
jbnsDkpmR5Mv3HSYOxvQpPXUILY/KL75w6YFN/CklIHgiX567YWgcMlwb5JauEEvauFOl9/gvspU
jnJCRSo0zWnNy3CVeHsH1it+9HW1IRP7bCY6g0zqq/zsQAHc82+63kaSUvwaTOJ0n8b8Pl0Teega
d4BRjqVZ4KGHWPGwasf86CY3gL8yWerF/ZOgxir/xjmnVXMj98D66zJP/2GKwJF6uQiNtBhj/Oyh
LmoyK9zn/mUZtTm3Mz0ZnzU+pCZpIsbhLSwI9nNaGHi7GCHW7cLHenIGQZV2TMLXf+lEjLmwlTY6
hA1hPJ8S1YigtUV0Bx/nhSP6o8GmcjyNKH9BGSMX/pWuSDQ/c3TtY1pboCejk0D1T9f+7um3B22O
1RR6y+pBEEsGRPvcX8dnKCuAzwbOM3DGX8yx51eaXD9MR9M8fFvq5sdn1baqATOqGLeP/pjgFu8I
/j1y7XS1lUadFPyHD5Wn3lrNeBb+GS/WVRZLih75Xa2OEX4ftm6maO6yFIDl23Zio7UmxSZZ9bbx
IfCjhqHt9Ry9gIGltn00u6p+A0ZuF70HA8vORI86HLvxMn+Iay2N20LmMh6d4wCF5MdZHoPKvQir
SKN1vQZ5kfw8EkAHm3tugVIsLB+mBZyXOFh3MDmrfiZDqxUqmV0Bwe/FphHMaa9SHWMKdCiNRFpT
b/aKwwj7oXxcBn4MUR02J+mXjowGqNktITVhrcpgKZ144g9OYjwRvR2X97pJ6OukqtpCHyMfpKZ5
oUIxKR/w59toSecgPln5ZJEKYDit79Yje2lTlzBZ6Q3tX475hKlrWU/bwVDV+7Dp9ZCf7Ivp5qxN
UmQbbrlSRAYMpXXUFDNSPAomLUDBDcaPpZIKrbITUaHLISMxwVSi23QPL86DhjjWufpbh6vxRQP4
AJ/xDZx9G77Ys1HVdCFMqiI4Hs7QCI0TIjE9fo83DXk8EI3aTfNyRql3/EGt+m/MAYNqB+/gnEwi
1Wbn9J0eUEWFLmYyVvt0JuYdFaUZ3Euf2zKKLx6JxF5dkMAUa7vUDyXQBVUTSoFfX9XYzxm+oWU8
LSzw2CZWEK2dSufU0czZnk6TJe68jGnz/5vlpXJSZZvPg8or0XDQoyJWG0nOiOG/inVQH//Ds12f
hBIpJTABU0GY/SMRkjM7Y6zDHxlDyfwYZbJNGICUkQ1mXbsuumoT9BTNvA99+wWBg0uMPkaxBInK
hWDjtcxFVpvz6lrkF82gSLVWG9v8Ay0ZTmp6L7Y94iA1/2umkbm6wLqGtqwDXdtotGja50LpayEC
BtaXp/LhH3c9m6Yg8payPkeBEzf/YY7Bpr2c+NERaSYyleR5aVwMtrHP8Utu/dp9DgAGhgvznTF5
EjowH6cuCIsam8LrdA/UXIADLzndqcJpMc7/RIhNqQlgsMcomgxsOTaMhzh5ASlwmPvaJh3JHc3P
kIyGmCZp5QEeV7Tvf8PMOJDCgazcWTqlR2eOWukn1kKyJOfy9jTiyboY6BlVjWx1BoVGEhEuB4Qg
WHYyYNV5j6sOVI90jIdczKBpxfWi+l0znfH3SiFYb1ZvGtPXXwIr5Sl59lLdVOGBKx07ZZyZi2CM
AqOlKTXSZ9+JypYQdCpNToTbdMWlMsS9iWOMREsUvnRYXtwNO7wcq/Q0bV//uQOrlnU2S10yefzc
BCvoig5qBSgvxE7K2HA3WEPzhJbKmj5e4LO0/xBf5zeDlnMS3S7QOhat/mqOaZ0Qguj8I2u2DieF
F4iuGg4oAvmlg2HvIsesKFj6RzdoC3sElnkrL/CnMkbNVm9esTJe+DX+ymgr5gEaOe+TG+cMNspL
jnnmYMWEUGwt0YEum+WsJIIRP9bfPJWrlVjAo2ccMNvQxBdQUQMwmWNcOy+evDvBRFm84ubCE1V7
eBIu4f6ubussNnpohh4EgbhAWGoa1xKjSjHyXdnEAkK0mBDD9zVl6e4nOTvYVLQntQoWajNLtyWi
BK9SPQtevmDzs5Db0uRsZDuE/s6kF8X6OMtCzQTV0mjJRZ6hVCfdpsUu9linYus9Y/wvTqFSNMpA
zSth/OFiwk7LpFdjVsnwncnTpytBk2K5thPKRkLO1zccjWndh7EXTz9DrLPoyTjqbbOxE3K4VHac
g7kNqQURDrH1Kbm5nsKoyMxdCm07ddNl/Q5PxQzYCvYjGJE907xIMSqy8DkChKqrJPmO4MY7PHDt
c2xd61T38RCo6j7Qw7Ip5S/ouvFBnN4GpOXzTKbsLAod9IC4Z3IY4wU5troNSknK3JKuFZAps3vv
48c2D5/c+xPgquV6RsxIb3U84uzEheO+55dOF45g6OPL626EBA79qQdA4nHX6DT8sJcexVfHLdaU
xAyo6L+93Bm6AiVojm1E5+b4SePyI+VgELDGvEMUA9WCNCbcSsBAq5SG9dgeZZaaXwjHSxRpbJpX
afnDZd9NgKdf85laAX64uc5/QX4X5zYUGDuXh5Az9UF+hE5NeIi8RBy2oTMg3NWQBjgEmiKJNfW3
IG465JAeJvSdEr6YKdXKjoS6JbnKp2K7IiAySrf4T0Hh/nIl61X/bftBBQEKzw2DPp2wFHvBygYQ
qnRDfxQfWfKDAwIYtkwb5NprClDBedCt4AIvCyJNkWsNe8CfW0ypBiD0R7MeuTlLHmWNnXTpZpqE
e7Xjd8aAK/bKjOuvGgtVN0HB+9yXPIf1pKvW/bkrKApBBs8JziHsxh52ms4Z5ag4bxzjXpBCubpR
APldEja9vDqzMw9FgdFr62dYcYBoFebocyGvriNXg1uLE73ucWMKw4eUr5ISTJA4fEtysw+B3Kr/
gZ1lZb8cMd1DNjg88Js7jj29rg4oTGW/W36PirDtsxgcUjB0eq/tL4oNSIHVd/URfKOeD9H8G+rD
A3ozrC+XFzHNqhakRcfPKMaddYgfF6T9Btq2OnQ0WSh8NfxM6HfAqyslazROKZSoYJRUd0ZScgOk
aAvDBsoYo4QdSMZIYfYsWC5oBpW+mGlIhiX8y8ZRlcpNAfQF/45JRQqRYK4fToVcKzMrKoUMZMmy
1Ju3LIzokBm6F4Twzrv5asFxr32udMKYFN3sUAw4735ru7sHQazs+nrxouzYYQ/tOG+m6Q926bpf
ZuDgSOzK8EBh3z06dAi+LLxpWB3z6YnmdjzEj9jX4T9B/2IotPDhBazLLhWzHSXnggcyf4JIVrtX
bPnWWicA8PcDvA0+qhn50BTrcqyW9PaB5H2TS5YSLRasVNbtRBgV02qyD+djoLYC269RXS++QuGH
RyoEpMclBitIQdV500ANYi1YrnEHdwCpfT9XX/YjZVDPLzTnHBdXRwPnIeSvCK6J+lBSKDR3Seoi
pCqlYbgXAM2n9ZZoyySwlm7RqGSyc9WbLzJoHY3hLHgSHVMQ2cTuYixMX08ivLc8UxE3sH/SXZ8x
5esPvC2rnzltrvq/Cx97jxxxQSqkrM0Fogwjk3MyUGkVakQs/DjaROwMJlJF0zQiEMuRu1zlTxXe
2WhHOpybt9UBfGnwzwjqo9D/363TgaftWfTVeHvnKIb1E76Wkz8xP/HTH08JcMFfKJaN31DWIjEd
OIq8REfH0pbX1sAfmDbUra4Vt0oPHafGKCtuh+DfEgSHoERAqUU6OT9SILk6z6dq1hEEccgK4egK
bVgM9FujN3Lb1+zMcIPSNG5EUERlECUax+Fj9JlBHcuqf2Dnuxvk7VqO8c422MTVhCjH38rbmnws
zbK2I3oX5IIAECJjbfTKm7VSQs3lIGwErP5Mcldq7Ek5EwJDwTTxOp/Eh3h7TZG+Ay5RCvN1wOGb
ettgJWpiqFJ8nBj8r5DkcDNposxvolZatfn23RGPvmiw5iqiJuGZd14nlookw1hEOWyq7Gnp5eaA
NzPQZIs2eq8YcCczT2lxeNtTKsFlxC/gUmPclpw/fxIpzTEWtS6IQdcOOvNt38yyKwqOsO+UXlHu
A1fcKHYpsuXxBN6HduStRNPixQNiBNkBncSvRHjIbgnMlLB5alw5LkAhSn6Ukcuq7bODmlbl5gf1
bZ60PEaxOdLAOwtqbZ2nCSj7YY8HU8YTtTYhIMgXWscrUQ3qJAhmKVNebjd/Pi01a6LEnKdi9VWY
LXY0GfOH5KTw1MiRx0grMQqnPjdC2YgQXPtJvQLsCpbuoQQYli7HZogxu9L13nYGI8Z5e5kfVudD
NYSoHPOeA+un9nmvPijbU29LSM8oTo0v/hUB2cizDES37PYq6Zx1eH5l7pQBZHWG8OpOoq+xjYet
JtzhwXP3t9ejSZfMpH35UpkIFVxzxOReKn8mbBJGla+FfEEbTuY73WnqqkWwsc3ORE7hqpw2+5IN
NcTUSJoZoXd0eZPHKhxIW498GoIHHKcvjtIpxToUCThdyQGk6lCmahqJgrMFosYelb3bSemJ2e3m
xen3TJDJOKtiYP2W0jgBLcEqf/Aqs4z5XSfkP6rwlH4YWAWoCfnkSDqK4NjnpzBOUfAdb4crUtaU
ESoW14DDJVxaIB+JU2pR99zh2YuFjnkgGsP/77ihtyRnJBLl9QI4j77x1rl5P/Ah067ejxusiY74
ASuD4vkgw2Di+endr8bBjlnllninkk4z27EYHrfN0oM9CpUKakYy3kK0ieUq2kPkFdMMqrwekNsw
KqHnkGYqapj7gyustFJ3gw1rXQMscSZMaXSgv6H0wJSdkvyl7erR+5377bRXLQ4WmSN3zNjvqhYG
2NEF44ponTyE9zF8kJQNjAMRF5luhjRBKCNEFoCKXK045YAUsb/qxwYhGcruMRBGjkVqv48DTIQM
Ik58eRvAHo2JFIRzi1WkLDuGppgn0RCR+P8aLvdh1N6x9cWJAZOqj45DdMs8b3DWqncT6NQXH78h
kcYCSYzpA+hAiyHKJUbMgaEV4PNP7TGbHaV8RoZPkvsrLOnHYXONSxKiKFp4jB41zZozrrFoGdGo
YMh11X48HqToPKgGpCYZKysGMaQ72EvjH3qYJ87+ae3rZ88XWUWmTewrfXrW9rjl8tDGIPi1ryWe
8070XWITuu2FTA5oCCrEeEiXBYXo90mD1nhizfVXyXPdV7ooFzgLLzyvQJr5ulKMntvUeMRuqFTO
cOCjr9DnwGnd+DHmMOROXWPxhuF3rpBTyAEsS7StJuPH+5CoMj8ffnOQgF4eJObIKVWu2GuwFfXU
eK7YIm4d4EvoWC3Ouq0w4zrpe90fz1xhgbqgstbdjPM8fHramUgdTDZa24f8SeBBFqgwx/0TCA84
NoISvk93kjLD5VQctDZ3wTmTDWcO9sGETnt/4VQ88vZcWdUWo6Am1L6Y7wrOcWdwIbxZmLCkXnV8
b//9lEaUbYf510cmE0JX1mrW18FUbaRSqzsPRARZMvvo79PEH5FNQMPbbQMb+fcfwJYtYUPxaO4d
87yAU+IUYVMDsxwtYGm0iClO1fm59sTAmS+toPS8ij0LwcngCAHLKRenx5ZJoGu7U14niTC2kOdo
Q0Zabo+zgwWUB3Y6kbgp209qz7d14yzd3BUS95ncaMg9+5rk9o4nKdqBF+ssjlvH0zZ5ofbaAQWF
BnFvZV77YYWtC6lPSNt63k8teBbuE/5CIDYHH3dUVNvoaL0yx6+atcQcdGWWfX0xFSzWeU7e62bS
CUDzRDWAyVIRXU4heT1AVfD2n6FeHxvkahWUj4d+xGF+nBIp7G2GFHhV7EfL2sIZm9AJ5a1qAIVv
9z8nebAGWorfiQwPafnq8jBRgeLSw4jTF8KMVhfO4QGriiOZSF/iRmdqkd/Bqb4HZeVkv3/wZnuf
fuu4JzY016guBxT0TSGRI9cq+NJy9HpdeAs4ZMwYpOshJzEF1blLvL9zd4dyq0CoviCfZjnKhYkp
IWd6tykch11J4k/MTp79e6G77ilYvzzOTosMYYPuLoQrcK2j6rUGdIqtUVInI20Xa09Sg8uc5ajg
ubqEjrJZTb5PhvhEjLvA+3BgRg/YaPiJT0jjv11CT5vK7ZW5gpWl8AbeMteNrrSbivsILB2Cc025
/zYgydTetM5BqJlR5kehnNWcxwPN8sNF4aj6KDiSsUQSi80VxqjYpdiYu0SkdY+UaPgpFA+etnEE
us1+RnvrBGGjiMMkA78UPtMCYPFqobbMD0NkVlbvhp/Oa83vYa0qrhU5jWUXlCvmdl6mbHB/qZYs
1WT+OzxBffUVxlTC9YML5JA4XSOD9dwO4QRNJfYmSxQjQSBtzuH0UkMWE2TcNGdnAF51wkVT9NBD
GCKi5SiEsVYEpugAEOJMeRpjDNnMb0e1F7o5E/QQ6eW6XiQR7HkloQsZMUFK3838nWDpzIKD8IMF
5F+ZiBUFwOdkSsCOIc59+Tpuae1DezQ7KQG4xdZI6RajQ6yGJ0JjJ8hFh1UL+4qn6tht7YEjIQtQ
CL64iDrAy5C06kGp7GYzZYjZcgPnCzZQPq9GDe4OND35cqMfHDyEtrEE4fyociQwMYlVjgkEBVkC
JRngUgKDy6Gbjk1ZVEYVRHp1PgY9LhhciGwXl9G6BpmydmnbdGwaVGBYGnnYh6R9gsAlGAPMrv75
i03+5ahO9W6wy75JBkuNhoxZY1rvZMAwNY2XUALDyTlDW1DzRogXLcLkB+mFdatVcI8ed6lfbBuo
ljcKt6sAUVP/usIvWdN2Z83J6W9ThHUoPKApHCfkE3ijJm8++vICLymgLYVFyhp+6QVMgldDvpkp
2kJx60rr8vaInGMDrtkE3KeIs68JBDoqsYHxcGJRtjdevhItgEqaTnnTaQApMnwQRQwcSaAlSMVj
1lvKxSEZG+Hamtlj8yB0XkdqQCpeT93l+Lr6uoKgepmF0n4O6a7ywl8MxXQ+OIq3OVnxoShrH6Zh
A7agL7tHqE/4iojAz10I3Vy0AUztQfVKgncsR7Wff9dcoQWjIBCAALac9wLSkAxGykjk6lv4h/VC
mtvBJ6G8ihL4PRCJXKgsK8HrjT711xEQWIydmXBwSmCxyL/5TElKe0ivBHUyuPYUgkJ5ZGz9kKz/
j1+UX4pd30qilzgYCncnUIK/kjA+lHD/AsPypt651OEapKbHBGyMQP5wxRFL/IBs+ItTF2fUllFi
FEqfCoU+gdII4JJBhUaCTRylNN83qtx7lp655VhXlXwYqNCgAPVGm8L1v5RcY6n4thSB7a66Um95
uHb3aJf/1GHksbqKTArW/njCDbdA7jrsKL66O/M9LmsHY2y7+oSoQJ+42twbEdHglmyBDHAFDY6O
XLDs87S+Nt12ezypsYV4NG+sbfcdDrSYbOBH2Wm14phB4ZnOnlcW630k3JAYEJbof+vd3tScQdge
GlXr+pHk+s+Gveg0ftDRiAwV9sZIPUTFnSW5ATJf797mX7RC8WD621SesDUJeFdPeOcF0E+FoR9M
jGtOUNT5nysXbk2H7tuOxiCrGYFgXAbaiOYZBNfX9v7x3TVbER45wT8+ery2gk1B/M+fMjl0G/6W
QBBD2/kizxk6ZTKq6wSRqlWCkh2A8yvC5grWxyMfdo9Ujsd0yUGYRLdVmVzQ5Hk4REIdqYcGuGRz
unUottHbAW0RwJ4Lda84pR/thbenJd+UsVeN7EgzOGL8DXxVxeAVYB9KHf4Ba6bonTt7CGHbVHCs
6l091taUnHAB9ntfUYUaNZrfRkmFRocjWtAaFEsAptJx6HB4nZ7eILRqUH8o1IGB1r2WpzToNd6F
HwdH99wGFl0yI2NCcJ+ntt20XcSBHPPqExHFRHLxobTzdJvSjDxZGd0Hz7v8j6bOytk/jIAH7rMA
nVphLoB1JHH6WAmv41PayiVKyEpgN3peJ4fG88cVNtciFabMespHPl6V5EaHOdXi1I1ca1X9NUNp
PZdwm5jw7UIlnobYMoVwMV2UjC6xAEqS2vTgvb0KY2IUxkgLozU7TfoRijF0cRcTYNiM5pltmP7/
skVmq1mj2j7qNmMzMSETHdbdxOK00afCtBUnoTN3JYW5l2g1NblrLtMdfuwH8UUb29a6XDGSw9pd
daRGLdW8EkjNf3iPfDgasvlEI4CpZEZ/aQkoBv/vfMqXVkB30pVhf0LvkpdD5+RSEhCTgkr5YB0G
hRUMgBauxF4cvj604VKjAKMLkmFMc3kAzbOk/uDmOh2L+z7ZxUuYolMhJZca9PVk/SNyhYvhOhIt
6pxfoujEr412jGa/E7V6U4aVCQGm2RJDKixJ1LkJk1z4nFNjznmnxcT4Q/AiIotgEuhl+esgNAgu
wHIyRAeGTYhW8PKw1qjEOtwhgta2XDjSrQm49VE+yvpHCL9lXm8MwWl8Xt9DNI+l9FqMShaHqjDB
l3fHsmgoTTepiWVv4IH61/30Qp5pD4zd95m1NO9G/4oR4uHA+gyN92dGO2r6t2mMCe3b57XusmX5
ms5re4bg7NAi1oXnXawkXucadnwh6Wmu/GTr0TWUpFJVYw6FaqlOOu7g/kwRCq2VfN1gNf7SbLwm
mO29K2paRiP+lKrvEz8mJlbby8qmhZ124Uq6VcM/hhpTw167D43NIAKIGHLwLlWJJRwyK0TmUaZX
3Lw40qlxMlbrcGETmDvLDJWrlO5lKICZEWfuSKDAmhLVrIVle/bcXukKHFyz1SjjPoevJqa2p4Xj
IOQNlE0HYo/PykDsA6QFCI03tyS9PegwfBii8kQhDjA3xwaM7awmhm3a6CLJl/rmLfNBGnSLzWMM
qz+wYalFGHoMP1jwvBX0STjDNeoos4aD966XprLvhIO8kNsYiTgMYLwcj9mgoy+xOBEjcJpvHhra
uzbAUl9PXVBDmMaLUbCTh2T9TlwKM/sSt6fgJM7gHHflwb8j+caKOX6ZgAn1ARiCyLduk42P5YQg
M8Dvccp+l+TjWc53Gwja4PDf/jW9GvmHPHg6WXxBxMT2AX701mMXcNi3diXKm+LvAJxyptnOKZdj
5giGBzPVtQShLWoQg3HceF07Z9Wj5861oG78Kdna2JYpmv4aJrb5soykjbXSDP89MC8wN4oMcf7C
BIwVKvWIp5cWPzPDVJbZeIXaug9C40NiHQ3PO5NM+4qxgRJ/PreB9LaDIV9Zvir/FkkfhqOYCtB1
2IPiYUqYBqgrk06aYevIFQRndr+s1q+pvIBzDQGu3RWjbvfD7cBTKDHOgqU4OkVSaD4zp1+3gdJI
32SD5Bjiy6sn5egA2Ix29B/6mNReHsHhPjAZJidbi77KgJqAZcm6mWOodOIplep7zlRHJsDtgzxy
m71m2O29c2DRdWy84dYunRTtEZVw3jUziCB5Y6jUeTlJ/bdIKsgLy6GAT4SJ404dWraB6R7wji3S
kvyqw5XtolqKGxtvhZtWoLSToZz4N0cgXRUpFMdOoBeFLyqCUP0eX3WJT4+KCcv7I66HYaQnNnEW
SKnKFPvlSRj0eSVinUo3YgBljDVuXI9escSnbLAaSGfx92vzL3H1pXVqOou6VivvTK3epSNOi89D
iuQPmADdZT2oWZUlYyRmOHFYFxjU3KnofTCkzVRa/t+LrDim5yiNoeCYDG1/iuFBXXfjxut8GUVS
O0v10dh5EGo654LeTYawtVS048sd4q5bGO+AhYE4QVq8j9V9lZQ38zW0sLCwOHTcAxcM6SkYXo7z
URY6Lw0ldzFKN0vtkWZh/cY9sgBfKWTO07jGBidsPlgQ4QwZaftSNTjw3xtPYaQinzlu28EdcHO8
/PgsRe8m5B8KurrTQz5FvIuB/quZRpFxrwoF9RPph8aLaMcFXMrkwoi9SOm89IAub6eyLYoOXOCE
6JZAIk1bJcWNwwK4qSq21R+hT/0QQD4y12+o+pVaRakzGhCr4PmMqUz4eHb7qZn/f+Z3OlNmjC2B
yQABoIVa6FC0Q5x4kyWoDuIY1aEv04ot4DjLhcVqeCsq/jQXIVnBH35+BHKDJ26GpUYs3j1ckSuo
2VYUpwV09qAVdcsUEAu4Jxav0deAkcyTUG8h09DSriTaMGvwQrb2CTitjV4cNATvVjWRXiqeEGk6
kA3PyMd6c8ZQmR4bQfplZxH52FcFYpP0wLY4lR3KFK6ppj6jrEFW4Vo2s/u8QXJRLiIFBrDGI2N0
q/VQC+2f8nMnMzSfmLp31kbbk4V6iwMJJSAn/N3d8rgEi0c6GsuPejJBOzjqMv0wG/R72ZFRTy9S
k/473JSPgQs2j0UTeB45lpVfaAjDI3RuM+rrOFkzQgctvXRetODtAnSIGms6ulXVpU1TQRrsWoYW
vyy5YDTmO7/WQPJt1/EQNG97u91JSHXZgWisaaMlQOhuUtK5+DU1vF+B5WUqXBquFAYzs4r9v7tH
+s6rXb5MZwWwVK2M4wnWqdOnWhnxVZYWo8Kh5Cnb6r4EbZaHUd6nNeQcGqKc5/Q+AqTH3ExicEwW
gjk9/CoN0d/Ix8Ka/ZLSy8XWhWitAQBzYH2h97wGDJ17655Zj2pCOf+iHiGgyDF7b884ft4CJ+R6
znO5wEGzXs0YCO/2EJOeDRFqVPB2+Qii43T6rvQGC6FBGIN/3xn9Bm2v9tsUP76a15ThpX33V6tZ
/nHu+9fVTENpQYXnMuenh65ztA/2J8cQuKfkHoibgC2v/8D4dSG5wzjkZmFegVH5nf2EdNFXighb
H7qrbSEu6QX7uAjB7BpqaDl2mVfKLM85TSyGnLVOLqIZ9VndL7MUQv1Y4Vp0QSCWT2OD+5rGzjYX
OCOCYJ73rGFESYzHZNNs2OVNsIs+pVnOqBDRi4rqDswbAs1wA6O3QJbnZ00BnFGsC32xnRIMf011
I145l9Ne/9jf8XbrvdhJO1ZSZrm1gTUmYXz7d7o+kveRjWcCjqybc+W1U/u/9xoyzQGRs4OGQC+A
3jmczdfFndfVCxl4qkm3SuZjs9h5B9Z+ZJSBVAyyG9LgNzhPLvTEYNZSQHxARoCeI8AsS7jE0Zcc
Cs0L5VeaUfOC/pmzthjRkDrs7HM7gctDKp/XsygHhOAjx4FgwqPO8zOCNbpcBG5Q09X+DkHeQkvm
KSNRr+8QJsFEStpbg/iRvcv7hAf/KrVabPi9MJGlV7e84KOomCLe/KauzBW48k813hA+tlJDXGJX
kygXMehtD+JXWYqvljCNgFzJ4D5TccEXtrECXi59tw2pmVhfaEn4JKGkTA8qb12fBhskFXCH9LuL
r3FgsPiUrGKWqlnG8TDUNNyCGtk3oYlnx47XP5ya/nZhszx3WM5VjnSNuHxI4Hcn9+eevz0X3IHK
Xmwjuwu+s74i1Ec8ogYFBqWvM2Zn4Oa4+75Mz7PrsrThW8WNgA6jra0IQyVpM3ctG+It41orzz+z
ereLJaxlamcyVyu+Ym5fXXh7Oe4FMdFt/RCUTb7rKMAFsbm2xAJpqdYoD+lxz35ovin/j8let56x
Ko6vou3F6k+Lkc2QLo8nk8hg3XLYg5134FNIz0XdJX98wuUbhvJpaxBj3r0REbOLdceG277YhnkL
Y7VUAzBLJNSvU/mXGXRv0hAyFleWC4XX0BBPEl2D+TCpAQu+MiHX4nFeJi3NHJoz6wWROlDs3y50
w9JTYSTeslWIixjtt09BesWhtWQwA2DTFlaBGs6yX/pl3VIpj34rh7YLpBSCC3aovF7oEdyfMQM8
ZTJV55A9hByeZepqDMDiTKpBTT/O5ZRRjDUcg2Y15/j8HLwLHHAIwqzajHvdKN6xcUq7+jYW+QHW
pU7Pro4yGkDya6922HEkBrA5MpwItYxP87TRDLuH8FGqULj6CwDF4Z0jj0MPCyRG5xIPnoisgCYJ
b6xN+Z3J+lSD7XKXa2eeQu7YhAoyQ1dOSMnZe2JpM1bLXL5uI8Th8yovKtIAiJBw9L9BfsKFYW2t
ndnKmEQXp5ZmJRedQTUYNuypHdCDG6YC/tJ6KFXI+kkNjU338GW3c0vMlRsdzTLJ+WFPDAOoSX1b
KNYzCqzaI5FIlKQYYWeV+eZj49C6zQCp/M+LH4WSlOAswPVEdj4/otFdPPGjKxyzZzKXoXJRb6hT
VAG+qGbaEwwi0AdOooiKm1GR47adHfL0IVKZgIMPt5/EVZceKW6oonJqgElREmsb6lRTQxYYt58Q
CHUpUTjbs3Cs4jKXsBwoGu/rE5q4f8uYvbs+x6mRqz6eVZ/508c2C8Q/tw2davKlSdTgQycsGD+R
6/s1oa3826kW8/LdvbLpHJhbymENGTz5gE3PpsS7cca5WMmYOtUupz/yXplCKiYoiGDEnzjk95FF
KSEmUL6I0hsDj0PadMoaq7qgDkApLkx2rb9+1zrqPzlA2scKqo0QtaQvMv+cpCrcTKjweGEUfJxz
OdBeUBCj+FT0gJgSpwrE+p3z5SXLbNH4vpnYMZtLVY+oqU9DWI5aQvftc8qwsSZPspjPM8gFb3YR
LlXq1CDdJWRn8EZr9+s8vHpf+0fNemi/vphU+K21tP4x16tribakScNkvAfYJD1CQwAWwuCbUytM
4IT46dBeQzkoVqXWVe6rtKae2BkPkgABt9JNqLsmzB/zQ2SHRfi9Vy0skUuymH9N0G18SFzU9KDa
k6aL/CjuSdBSE/Xsi8lW4D7Tvazd4AMtontVn6du1QMpVpP7J7zJnxJbr29YbYdjWV1F6oJiihMt
BfF6WtC4Y7uZ/qN7ek8ZexzQ3icM6MZ3KBiCA+w1kTJoFpkqb2ZMfk2e/5ArdMd6hlyGIBSR6cNC
MGrUl8Cb1/7vLlNvLdJZM6gH/ZP/KYnN0MA88W9aiNtAhRS+fNOeasfSKC8f1H0LaaBb4MgS9nzC
3SRRQ03nu9Q+qucJtP9jEGkdE80JXoQR7wxTuYYD7Py9hcGClJTPSeIzDwEjLHJ8vRbmw5Vfhdhb
aiJd0p+CgjubOZj5kCDyqAuQMbukH5t3sisvPSQLMIqnxfs3cInWfKpZIo7drgCEcyVD9DwDRGPk
PHoHlG0ffoDqWnncawadaciCeRcsk3hCRnhfTNi/Y5WDrMWFHAWyCLfirm+BHZRde8vQNMczVIa2
BOA/v2PogR2NntTws/4W3Rw0y9aNrjD4YunXME3Q7ERjVkNJrq5Uk/+HL0bIoiw7MA6W9/fm5SmN
RmM9yW13M+//6llIvmcarVa3CYc6HOfNKtcRmd/WeoNL7XgHQikG2W9vYrmDDb28reJvutx6Ukbl
lEz696oIjMzPpxwDNPF9qsX7PB7K240lbZl5pHAgEMJ/rql6HxScOEccgrVkFW0lKO8xx7Dxi42l
AfA+84KSIacn2raN1GU7+0b4aDbEwGjTcHbvfUbnh3rB3sdE+GgNQcBP7kClOCIUaVVIP5p4h0e0
ZAHh5B7xj4BX9ux2d8ci3qB33WXxS4VcBPMtcuD0e/71BBafh9+5e8oIN4px8tgUqXo5MC1YEq0L
75+UsuOraPh5nYDj7NK6tSR6pw/N5RWOYDe9DnzJqdM9EJ6psI6sP0bMy+NzdH9iGAZiwQQ5v0s2
NqACrG9fMYwZp5mvtbTsg3U03og8S7kShHAbhcEy09vrvqfLQzcyQPoTEIMdYYFG5YecAOcvDyvg
JwvhlHTUWU6MwmJ8e+3VYRvG5ptNAuPEV1TB/SAsf+CrC1XEUcAD/H2RswS8KDyQoCOC9ilB7UAQ
42yFw4Ri9eAN8PtWUJM3WVjYIJ1HF+ZuPVlr0GL7pBUJL4HRQykkhvk4/1WZBqArNV+64cZAQHuy
gHx/X5T1NKqmaaPAYLhKRnqsOE16JAhs1u07HI/O90pSKVY9fMRG+xA6IqRoYGKCBRQGsEA2BsXj
szP5ntlbk0lkPAugaHfTGhepRhff+mgvdhnugO4NQI4x/+ISikmfS7Mdt9xgYNo9V75ZZ5ojd0Uu
PrUEeOHqE6aSuwpQA92GQEMzPYunnRnUJGBDgxb6z8x7MP4jaFiyyetvwsvBFgIumGyRlKgccUxR
WJtjEVIu1jyPzJx0c+fhsYu9ZjXHhXFrATTjeBH8AWaNcpCju5OvXvM1YeX1gIcN5jcdeJoCx/Q1
NkahQQUl5IMvr8J/n8Qu4FhBMJNvUiD+kNGKzAgCQYqlrK5aQWhPSmbuaY9KVF19XH4C+eYNvsrr
QX9gKZwUXibSDQYCpEJaBzx0UJqdszwDj3pkSzLZTRbGflatqpDhNAbbQiu15jyYRo8hep26vG5N
V91al7NYXyVnmWmGpk+FX/zA4Heig7qzNx3SSdtiW0nEZAfHa6tI9O06TcFA5F+CWYvUJzo9p3JV
vp0GO/JHRX6YbZpeIz2bpclUrY0eCya0dVayE7fl8U1phdqFs1QMg10X2ZLwemfU0lqLNWbV4Fjx
IUceFvqGnAf9D8475bRhgTvf50jCSphAV3XFhD6sNcCJ2GklTyj97e73pHEGGM8JVSPfD7dqB3ob
yzoa7M2v7pOi46F8NFCzF1jUDHXNqiDw9YgQfTdRy4qcD101TCFIicMBeknjRIHYKzeAcUdM9Hyz
XWkfSx7IPOKc2FOFeQDxluKJdk5rsWzq7IwKmUSzF1EC1Yw5drdih3XyIV+SeIscsElnmIwKZJsv
0YClZRWkvzYPQo/fpZZ8K2AvqFllAn8ffom7pVLawC2pm0aicORTyNgGw4Pa9MUxV9U9RXk/8fDM
oMCWtJwaGU67fdapxEdSzin4Vp2eKCA0TcPaSLuqb7+LWUn+BtxA82MySob+vie/+jjYzlryBWd7
gnsMuz7pTA1PacawA8KuHzY4cCiVLCGSUOYaqYGxwPiy1Vs9fOctlqmCKqikYrtXJp0I4AzskKGL
MNC4ec3AH+0goMifCq1J8kZfB7XGKUrkFJ5B0YHIsISf2OHNGfbXSQ4fjw2OKzCoVzxw+RmCxTFt
vHQILcx0N0Ui1y+hIpOleZ+OtXbUW/7UIOhtm4imYGT5dzBFJct6LLXNNF5CWOzpi/ZwFY46jO1A
b+aTvcdWh5uS4oquG/LJafC/ZrEW1gRMgFSK7cO2Eh/FTFPAs/2uBgU/Je0jYtt8CFa9C5unSeI3
McYKs3jjZ7NQzZmmQrzqPv2fr5Z5gZCf+eMADzvJOY3QVoCce1WRZBV/569i75sQYSHEuC1JjEh6
w679/IL5CMupdC3yyIEXV64b5p1N6juBjFWrVK8kb9zu6QngbnXtAFxpA3M0KWvIvfaoQhVywMcx
6JQ6fpro7MqJ74EenP0W3KnRPiv1p6/NzgDLpJ1odYICPh+2g6XCT5pPVkxWo3qKhvJtnf2EQRva
JJzvIoiIje7wHsXdRyWcEBocFT2E/83wROUB7HBldtBnDr6291gBvr44putu4Kmn0SGEi0BY9u9e
jC+rTtNRewYGoAYL4ahKBMEF7oV5z20N/sqnKLi55FodjsG1RN1mUqINiOL1zCy5Q71gzjjvwx5D
rkOUXMxcWp2VK8NQ+sspx6dCjws2dXOXWqjtVfTgX+P4VCEuqA3TbnkrXYbAUoCyjonvWf1dWN6L
r2AYlSpErGNQsp444n6eOSaePdZhO/hw8XVamNkRX/0k091virSjfb3wsdPN2InVOG/DRaarzCAZ
s+f+QvZxoK1h8zdln/rveK/gBLNsa4zdddw/04mUI2hrxd4Tu9dIg0f9QuoiJp1JMOgb/f58zyi7
T0BOUrymr9gTe+zEmGdYTodS/e/APDpflTB62gAg9i+NXjDGyXTo13CJxohjXv71NTw1Yyg7R3UI
wZFQcUED5joFxHlVnQ0wdxE+AlWzWXiDTSqU/aukqmsUksLRO73JLBrdgLMLWqvRiF+tPj2R9Uy/
xhySy2lvmZAF0ev0yBCokFYG6Kx7aPGb/HfmPM+bT76/VikJXau6tugrw6FQ4EDZPUzoBhQiqtFU
minfdwpB1ffrXwjoDoy5uUPLusJXi+250+umt9X6gaw9wm8jkxP7KcD0gWKC9rtzuVnK6xhnsRQs
TIPDvu5veqbZmhzHOMd/PUu1FtEnBc2xcX9s/5AuAF7eqbKDWbBhpwuxZ5oAPZ4f57SOawzvVkC8
5pHo/wWiS1ygWZ+GDK2iHnhEiUgSA0K/0MhtTbwKzrdSLUFQwCSA8oFVqYl9lA3lth2OY8jfk9WF
ECndYOO7mmWeh0VeZ0VthlnpUjRBV3XLJ405PZ16BoMQ7ntR+sP+Ml0bU6sgD+p58bAyAE76EWG1
6k/j6Auc/Ie0eOsdylnBSc+HibWv3ZStY5gbwiCfWcpdeK4zslfyk7JwD3gKsT/feuj+Ar2AcUDi
+4EVdJNMVGfXKvZiZVASiP8iLK9CD2IRNXR+PBt0AHa2ZAXRNVDYUBFGH/2v7V1s2i7Zju01XVYc
pec6NCJGCt8KeLq4Mm5XFHPTM0a4ug/f1g28dvPipLQ4EHYrz4mMXl0j5wBl5bTvB/7oQcJLvdrO
Ntbvwjomvdp/zFkdTbKSU66VTMy7+I4pzihAssFpZbcb1q72c5wkZ7pTXvivVD31Xju0uex8gZSx
RYhW/10cNHDm/QMi6R4sMW0+yXERX2X3yjO9JSCVRZfUNQPl4fVLXsIIgMKWwMZm+1cMdqhcSNNK
/B8gfz7aNlz7Rbz29kUdr2NWnIZtVV7pGKl2Fe46kTWgVQ3hD7RO3hwkQuns1a3mjZQsh3l9F+58
Sla86p6YinC9G8oYncb15J3SqRpKLmR7n04jNMc0sY4pw1md3v//ICaqvN7uPVBC61vkOaFR+PqR
HlaBdRJmcGHgIndA19knXxo03Afb2jcuZLe3080lR3XQh2wmGrcRolYItTtWlTevdwPbmjFbMscv
yk1y2hfMH0xr05p2cPJD1SsnL9Tm3PfRpruqeOofUDJVghPPwJudSf0DlfWsd2j2CORWgZgVNsvE
N+Op3VbEqPCKJpFyX0pyv0gzL08Qjf3maqIzdth0kxmvhPT6hcY3xtmTakeK8sJnQWLwjwzG3wXL
ygYOEeJoUmMj9aU4Ui/X9T7SCCPfuw1a6d8heYdYJtwDBPcETg+tqORWVdpQNIhcjMrnbxkgh5dQ
r29a8etXlDwziJ85ZtTkGa8aiRjlzXIvVocSok6U0RHNcofg396kYK+xiZe4/iL+gFQBkXlmYXeD
C2fRdgST8K/OJ429ljpe93OU9Vc0qm5DSdj3VTw6bVdva3wr8cZjtMdQfPwdHvgSGEOLzh++jGg6
Z+iG9jP1Ddj6f+rDX4c6XvFnuN50tJ8lXNguRbaoEuVlLH4hEcwJBB86WG6VCjcx5lZC9s5Zx0uD
Xjzs7sGowlJyQsuRvh+/j/RZQAvgIHQdo1ucOMTWW++mSVDPtrIA0LdRhHebcvtasVHs+OMahENR
jSqmvncCgtzvV+XBGVZwz2xcop59et1xVbpBKUVj03A6yz1s+70nDQXIFtXXZoqXhOz01Bcn1swP
tzEQ70sQz5/42B9vxroz1wpgeF+wiZRTJZ5TsZlYlHSlL6mbeTcNLdJp93eRFP8cQE7S0uJ7f66j
V3Sw20xukw62YGzry+V+v+uSYZyRF7Zn+OA9uJgU6pql2RJClXhmLBzHs4vRSDw0Gtq6fduJuk12
cuBp2+nYxSF6iL94lh88XK6TD9uLmVxB2MI6tN2jeU0fgNsd6OADSTnHUgTlCayB1V804bjczgpw
nD0p5+BIoQzwHt1S40q3w2xKfLljRwx7KLZAinl+J2Jhn1piL+hwx2mO4sLKOgYx9duUTTssPGYX
fQltqBkfedyqTzgJfe6PeQM6owesSyW90Y0Bm90cvIM024zk3uLSOm7WKZtS3ztNLsxO0npNg6Yx
WcjhFpXBKKEl/mEeEGe+VpXNd1TScq/fE4QsaN1aGkLb7vJf/kD4+j9+g69Nx0rkwpgg7XrMeXvc
kv+HJOd6c+PYIKrCA24IoWJHbCVk0Ah7oFAYv11yYDNK5C7oFRgzPSxqNKRthUzvKQJLHV9bJvgS
lFPBGL49XN/k4CZ/7HFHlKCejmZTWJigYQ9hbwQnNx5Yjie8aFeWrcXIxsXd+noWHZ961ZFIHSIc
ecWI49fNRb7ugOjLxSGG4LDhaULTFyr2djkbXr7KnOVEZK0/vqBEGljdI9p7wncGTEetw7Xlpt4L
rc/2kfa/3ADtJTi70dfbrNMsN8Kzq1XaQPklNqxc3TM6fXgnNm4l0/U/oXhgXa/idb+NtTDSipVU
XhhXRSF8twOmDUMouzEOo+jHwly2Y6XlIty+/Lmg6jp2uwVof2h7eoayTR9VxpGwsahj2h7TJm+Q
ebFStMJIz7X9AQGhc9Ih7xvQZMt6kFnyzlm46fZmNv86WQ7l0twTXtcZElNrvXoHqA/Q6177zlz0
gLAlxF3E328lJboM9YPgaGChbhSM1WTRats47Sz64soTYO3AHnau5AM9tjyyGp/p+0GCo5dwcr74
ddJ84U5GBesb5pZjwxlyZQIGCOlpetpy+Ej9ozZ0pENKMN73cV0eCJtZTrl4Rk6TMzC1beEq949/
Qt+0fKQJwKxDzBCuZl7WtJMipe4KQDVy8RE2WN/3rPmZ1FhzGuXPeEH4gni+/gAi3KhtKhB4Ptiq
ms7Z2l8bjUQMT29ZM43TLRnCRqeKLCMPK9f3mjQ1byOPWg59R1B0AYvQA5QMlNbyLcsfxLwL7ogO
FWasXm17JGMQfJ9eh8CQPeX9lbFCGa9sdFC/OJ3Ap3Jv3jdUXXtfNMzp08WYFo4JSlPX0mcgSRfF
WAWgFnLHAHmDqwhd0vr0fIgnLQEB/VS98/ceJ9iWcN7Sn9fIa0eGlqDWwtkdNxJzzQeGffz20vBP
GyPkM/KqW5R2XJZBv0338sz8VQV9L/mIuiS7qzFkoW75HzIR1WldgFlAJ1Kdt4wQg8Alb/iwQ/q2
ebin4CNC6WgNWl+OTmILtGnfItARmpiqk4PTqjKA70OOdQ6BLdPrZzISV2ckaDOHb9gF62C4XLAy
4T3Etna/ku42DgTcZLcymhF4az+it0BcXf9SjJ2UbqJfvobKwwy4kQW4mKUYnCOgPkKcsGwJPfQR
/UtoGzMpzVT3hyFuksFO1djzKZFzDZ7t5Jnt6XgLWeliUUfByiLFA3hsuZhgnZPG879su6vxzH0M
kBCRlViNA5qVt9v1B8KqsgSIsbhKNDG4r268lM35ozLdusi8Hymh3AhB49CXDRD9WpqhVjjtnPbR
sevZBCYhUQ2BZhUW2eiCy8ggUDEitai9Y5/91NKtTYV51sjHDYebqoaOm7dEiAe5b0QHmGfi9WX8
qaDkcDP0uHM7T5q2IwTer0RQcYKxUellzvTxhRAjhWTmtDdZT72LjsW/FyA9mrVHpx+ct3h+Oxsw
D3d/6kvN2SCGiQiZicEEXMsVe904hG9o37fQ6J6gzCC4i+2wJ+2ROFwvUJXVGAzQ3e9+YgmMfoFQ
XBrVfI9KPyMWgvtXfo2XZw+sv8VbCrk65O3TvXR0tujMqJk6QxIWlmrcdWKRmlinaP5TjJMZpnst
cBva671QdP0wD1VyweSA8iL+fvojWEhSFRXlv+t8TY2Y5827pddy4mmr6fZpw/dv2JxSN+wdkwq4
kp02PjOBg8Umhk6Ff/WGBKqVTbSaJ1LZUtZfLES+fhG9y/28hPFDF8IBM758y9mdQTYKaKfpdcGJ
dHSJ59dO7uSwqhefUVOrAE39hFdTV0jWrlHLZv+Ffu+lshURcpah0RQgzQlE5qfbLiOm+GWZrpQc
p8RO/eCTHBS32/xPmviJkVz9+0YzOcMwcT2QFx123UVhWRBJ3k40JBOqy1+caVZ7RYKd4vfKjag6
lG8Ko4rLcJT7cp5QHpldQLrQQVFHsXz9vjifInkICEqzHwImsW25kZ1btGdQm/ouzZipMuOx+ZyC
HeqZwhFjAKS1MU58XYw5vG/fvQrP+pL4cwUSYFLUoLBgolZ+S7dFs6DpVPZGOSHe+91sVR/GQgGD
p4wS3CsgZuIkg5F+S8IcNtW1tp8TvDSgUImdEw88H1MgYFonzneP3B7HR4vyIzRhBkKILcJobVSG
qSa52jXlbKO46NO+Y9Y0XvUvbdUJsNZwgVL6FU58zWaYYl3eQV5y/hylXH2T6WUqol0RtQ1pFU9i
S3UFdYEDGo2wiVaK6O7kKWdnJCG9jWqt7rmPlKpjRzDbQXZw5pYwVm7iCMgbpVPqDZes/fi3Zy7y
qjQdkuW3OHMV9N/Ht+CM8kCz4ni8s4vRj0Ta47Ia3fpcvBjyOHBubBatrcTrtM2adFZqmm16U7b0
OvRizmqEL9atkVEJH43jbjynHU7hNHOZNeIEFWOlWfCKDbqo0qEmp/t5kcEVe3E1cmfN1zRTWWXS
pDVCfkcRoM7FoCaJdf+cMXmCZXTq45QKy9q8X8iCZTjH3WG74sWYB1mSAsQxKpcrZR1/BBZvtHAr
8I2aH7xjZtwAjEq5DUyuOh9EVZD9d6wpZKsRx3V3cdhPfDmWakiNvkMb8qywVCBEKMmRS2/i/Kb2
laxExWvN7Fwt3opFXsx/JL7IYhw8gBp4APLnA4/uG/s/CT0BAZWVsGx2vvb7tgSNz173nH5OEftQ
6NQxrnbUmJYmBSTQ5XDI1U3G5vl3LaaGXTtw4FlvaO7tyQf4YcQ3/cdcERyiKvpnPAYoCQyuE9WX
HoaeVOVpLDX/TfifHroic3DUIMXiYnsh9wh1UzAmtlYEurKtCkl9glkTb9tDFliOY5/9K2jaMttp
QtzqGSTWpmO8BVoG8c/4ae7r+9m3HxrVcCzSnTclsXzCXWGnG3VYf8SqfcfmIDp01977a9mzpG+V
taWS/W4Yk8BLecpF3MpN8e+8M6tfL26Qb+botq8pb3UJIXJRu2sJyPYzgdhgbjL2pjRz1/0kn/r2
a+F/ieJqoQIy/zsBgnXvvyF7ptEm7RbWKWJQcm1+OyvLC1rKK5vCQcMw2T3q/giyU3o9EHPuNLma
ZWx0VhGnQu3y3+otUALcA3BRk8Env7OrPBOEbjVZbiAHVS6T496fxnRSrHqhFrRSc/2/oX69sCM6
xRxzQNF/rzBJ8qby8PgWrpGwO1mLFRMfz6IbYCK2IdmiwTKadzDtCz2gKUaPdtswBBQNYAF8fcyN
4xkt7Vj4X5/isQG2TklpjEw9GhmPMFif4ZWZHKkE3WjVlmCk4ofnBDOidnn3G+XtWRENrnqXxjZD
oVbpf9/sLAaso2M4b7ZtERi4qgvBmRuip6sPldEt7Gj/C3z0zrhuPvkrAVRAfuKzLeIuohIAgcFE
0tEV31h/UwGsOIRPedyqoJX9f0Xlj46WIzOCU0nV6JleuSG15WcCntIekZWxX4ux/0LpV4wGwJcr
R7Rvro7yHuY+KuhL/nVbLcjDf97safuJPmbBpSzO321rGl6NAiO8SIBg8Vb9tn7ishf3olSyrx/S
8cCxvzF4kCu7lMlVhLC5Es/cEDthzptMv34M0pbINPznj6dU9Ky8a/sM7RPsBkZC3Ss3L7YICexP
ukWTc7w16dOgTpocAc8DDa8XoWzt9D5GZ3Tq8aZ21Haz3oSl9D0GKkJq2ZppC/UChRF+KlZOh5zh
lkigac2AyV6GcQezFjzIEuB4QSBjM6KBcn/jggXal8Q2+e+EjJb4yoJX+o5uG5db/tmLfsfHAshl
bmtE1oVm3+d4bhKSXsp4xjJc+UAsvhisrYn1tgGd+GDZdNNDTgcf3lK2AlceQW+ewT8XWB06HeGK
k2c2Lxzc0n2o0UzMsk+dnPzNzy8UK/v7cxpC9NYpa/fNH6KFVH3bmZ3+3SoFmjfOCChTUOX2/cUT
gBnKxkdqt05MywggxEHXZOqNCekmJcU6sk6o9a0uqBw4dW41dA8RwxlrwLZ634LeIsxt4XCL5RwH
Dgn7oAUd2uu+nddRRBDHAEpmAecG5aTV6mcMyW8JMXzp/3rnFB0wEzemDgbHWzccpH3QWnX7nfTq
pS7qwHNeQYxZFsKEzMsNGtbVxjQO5SuLZTjFGJDS8ann0N4OkYyu3D+iT/EePa4XEij0OeH2BdLq
wQhDaMdYpHgqXMnqWXQR0ShRtEbLCV+NLk6iRO/l+8PdQ3dTlEIr+JbSJgFJS9fgGLc0zEzglqTF
fQq7IVT42xkO0r2IDvVlPFiAjgoNZzZEnVDFt/ELo3Dwmmwbo9Tx36XlMp+UvfBvBlJLvVN4hlDX
Y4tazW54oqKSss6dXWuNTMTgJ05PyyhPv3tdaVIlgYs03jtOp4cZjOC6z00gp874dAOEOp+0/aEX
CRQymAYAv+pd8ljEY1rs91Ks+D0FiN/NjKFiNkCJw0LUrbpeBSRGlw/zyeylKJrDodyBtXq5DAI9
DsFq4O3mCBMssfgBfWUaDmiy2jl/fwYC4wiQh/3K1z2KQvhnt+PIh/ybfx+VEs7gcclK2HXIW572
CvKVfJAz6SZVEV+7Z+AFBIeVIheUrsTaUZChqs/JtD3ttr4o8q078C9PW5+1FfPHXIDWhpQRD81C
Poy7GOWA2of3XNBwkIiyGPyOhCPdnbl4m4k2YKsA+E8z0eeEVLmM9/keSmLMf6d5I3Nn/knFE5qD
9bpub9P+xg/JDzhTCJWxPK3bhJG//JaowaStPuAkF5lag/bca4+rp1U10YZla5oBeBztgrvD44j5
7nn/2f6DP7uI/3eGb/Nmlzlhp9tS9k2I/injDSlJAo3y7oXQz8841bI1qJlyK91lKpq8M5JQJq0C
nzfrgGvvhcshvwR52j3qwomtRTgIcNKM6u8Yg1Zavb8tZLO77x4DnjHeomvLyeOTo6pIKqQD44df
O1PdNlNDZhOZtTAbW61Kkur/5HDmY9K9L4552czKQ8h41Sjxc0Eyg4SdzrCTJiCU2MDaoMlbAIb6
BX9QC+4LP96M7zW2pJoS9QFoRDh4t2Eys5uSaHMu8lcREjvqEFU6qdgf+PVAa0eXvXbccVMEJW5S
gxFW01IKeloFpj9s5ry/DrIFCdzV5Sg/oAiPAybOb1/GjxQFE/CjoBXfV/4HC05C1uT2CH5T58lJ
jXE6hCPPtIXr9iXoWV6cd7//WRrIY+dw+obLvnQUHiYi11OzWhdClbGBDK5VxkBPHAaW588sKaLU
Re5xBrkf5tFodb0dDmm0zHBt0nTVcG+GT45DMgpmYWwfI46evAk9nkml/p4n/ee2am9OK4waBNQH
cs7F8nKUNbnflSXbk5Vt6uJjrkXOPazZtoHqgyelmedpAg7ng6JoSHJrM7JGggNw/xEcnI115Q0e
AFvh2Wenqck+95/VDYK5sA+6pi7KkuWLj2rDBpggSmeym5UP2hCBF9Iwvk61vXAl1g0ok62ha8Tj
+91bWbFlH8er053ufgZz28nZLJo5DbKC9s64mKKpGlXekmPunFYT+hx7TPmqWp4YMoxs2fzZBlDM
ONwl9AUV4KYVj89LNsjocp+YcSMcwtKHPwen1QSy6SZTpfcgOmeTQqOyeaBM+WL4Zh7JHJ8fgE2X
AEFOUAuXm22WQ2JTpxaOp5ri7DliVgsbTQ+MpvNq6TfJGzoKvQpcx6XAeo9mPfJj5badVkUAbNmt
ceyfR0Zh6ZHqGM9ubT3vvzf50IXaH3HjVuVTYoU/zOC1+0cg8mxhqpOQ5AXCrLf3C/uc+a2BLWcW
Ssxt8LotC3w3I6G4n/WauKY8YdKQ8971i3UkOzdy1kChe+weQ4pbDZ73f0ro0WTJxd1EmriMcKgV
CGPSM1cwyENwCZNvXOIPXr+oxhyaSKl8YKABU8aU4UcYlGLn1dqdWemfWawwbIC1DrhlVxQ1IQhs
Fa9Giuz6lXtSVGyAHS+2IjzgGYuZ7jutukyuva0akKEhxIDmw867oCSsL4NVycBtCBhtG412cJae
g9RWrjAgv7fSuC4lOs9+zYy6ltAo+MtR1+GRqk7yFLAzpBLz0u2i3eRumHs2a1cV6nRVuANcjVR1
/3ilAnCpAZCUTEBj4yaWAGg34rSeTO0Z5Q0H0WE+yHtDIu2UGTC0WhyCFgayK6rsk6EHA38aHupn
BpVPZsBgBeaxz/IKxgQyz5buLZhuCCXm3V3amd0whSTJptz3QYLRPZk0wposVazJ40BF0DKdf4p4
QkxXNi7sLdLX5dgHcE3sP7W/BBTdS1tFAjyIRWaaeSoyaSo2+yxTmwDjXqZIdENimfDRNGXDYqRB
3F8Em+NOOq0GjBwd9xUolE0ARAIGa82Jf7vRF5h1MinNThrJpKxj1Otp8W9R8bcsP3Yqej9niyKo
aaX08/tJMVYBE48ondu+Vtn/h6XFaTMoqhHA89UwM94VVCwOZSXGFCRGhey22WEHkJH8oH5/oyOF
BESsqe8cnGlXIK/DVMozMtYtovOvPQpNY1i4FZyGrGbUWWeogFqqTL39z2y8t6iQi6GrwendwKPR
XuAYjckCJK2nmB6Ts8E2boBVrn8jJaq7x5w62qOFK6qkLiwJ5PO0/tk4Dxcutg2bBC8nTg5XhkiI
RuVM0zYmveZIwwohEjtTV9jn1aOkYTTy0wzznzY4RWqqx4o/52NYygW8wI4x3n21+woTyMycdRgf
Iz4fMQUZly1+6hMpxanb8nLKzVTzYfilESiL1PpoEWpUI1nPLpuTsk2KqFaBUysZleThCPhlyXuO
u8MZ1vj6N8rZD7/1WSMSmb9DtR455Su7Zjnar+Mtxz4DgdcGXVjt06K4ttZ9zUnVAzMRSn4g3WcB
RjRkg9kSn6TpaBAgCPUtbxMKfk/ejTDag/3e9yZo2Kp/PNjH+/fQ6VnyGuQKh7fPbVZuYcbY1lqk
K7VsGn4Vy38y+xqC6agUFe1e1b9Qi4BKDbQGbiVPaPKHKjyorKP3Mql9Gnz713UzVCY5ic5KZqG7
sqTrCiIZ/Z38vTRME2XzUfdl70CU7T5Ht64SX45WyoaqvWa/scGPSOaShMuHUdwaXm7pLFM6tSS7
/H9vK9Jmadk16Cc1dBXCrK3IUuDS/caWimPE8i9iJ2Zoz2FG6yOLHTnYUQP+9xx39GnuiM15C5GL
YJh4sR5P8JbCox/waTWst2d3DIfPpGBqCHP7a5FZ2BY6Mo9NO2IfPHSkapJBqUiHAvOaytKclF73
L/HtLW7y7tiDgtePekfUADeamDw4Abm0CxZhG0cYppSSOaB91SKyn9o1ITiohTGuG+WlcBErksYM
dIAs2ZSnX448Lb4Vqqn3CYybG+nxCrS1AmWU7F9/NmAvpmUf8jVEqahv0CfQXQAgLdvI6GH6vxjY
IiAJcItp+gU0YLB7BdlOXvYjoX40vEHAewU3vQo6QZLkgxgw4trcoPYayvp13+F3WBxx0gD8wkjT
AplbI73wBAz34g0uRVesW7zB0k3amHA569drQjlFzrQcmI01efv8BM4iCHDgJKqf+B4xRgM9iLXG
CGdnJaXU/ZOwvcVdFYAjRk8x4v3IvWPXc9k/m4koPJKxFT7gRdlmppuZfkYJOvVIRw9Sd7p4ZZW9
y07kYA9KvVVx4g1loLfxgOXR52OIChf5e4JIdsj9Aiogps0ZUMhyBazNmLge5whdERbV8Xlx83kH
H0iZqrAQbfmOgYr5bI1lUhznI+t8C6lOIUfk9y0FYmURZRL+CnbEf8+aMA0gwoXwW4Uzj4+RDwZI
gtcEe7hE+LHBvXc1OMdfOpKsNp2Ph2qrz9ckBJRJ6d88dT5/EvzqEpAWK/LA/kfnwXR4Flxe6C4w
f8cgjIaLeJu/retBTVIstahUqWYoTc/+bDQKjcd35gihOM/4Fy62aPWotB/3L4IP18zKYcQVua5C
SmH0mSY5wOIbY9bVlVPh/2hLKF2BInUfMGudhVbxbeQ36sNVJfffyK5a1EGm7VR6hyMRD3lbAqwb
KJvgGnXWJ4wKDxJlFUcYUEceY6FSRMv1FuuyMk3wlH8HBhlbhPLDEX1BCOfIBgisONXisI9JzX2g
oP0KwvhZPp8AM2F2gDNgRlYz1lOxhvzaLI0ZTZbeZN1UCuwQpPnwjTQTD8HcW0t+7cFYOHPKZxE9
LsrMILpdcKzIrR8O7JNdptRSvzNGFBeaHNkvtnsL/gIAySfdVDu8J8bbOzUDJNNZu3VTAVZHZMMo
RdrjsDvRwb5jGKF6o86Ep1kg7rYqf671GxN6U/zywMvOReMjk7yaZUiRBdkf4dCS1TfyQi4Xvr1R
UG7dsNjZgd02pb023EX5fJrNz4ghYgDHs/dOc8OlLDDHFvTt4uISx9TMjjXnjT8L8xwmHyEMgc/2
vYju+mgzR3QDepZHyRmwwUlZNoqeq9m00vvmkO5AxvKRO/pKi6fcRAi+n3/vCncleFyJNUwKFXYm
i8HwdwZfDWcmUVNTa1zo7ayn/Udpf6WZUtshb0S1PC1cbLRhcqNat+6iztb4V2RAac6R5mCxhhOt
qq/wRKZulhyKjPOsAgpptv4mlwX17h68YWP/VxAby/wzzNJ6iblr0CH8YSXAFi1xQ+R7zjlokAu6
WLmeFXubViER7ECGnv1j9Z8xXN9q6GbLscHxuydyOxB7y8jmMBvEDZO4zOG856eqrCmoTqs9asQo
tSQTw0A32JuqdxBFbz9AP21Y11M8K8C1m6KfHmTPgxCckqH+nK3Sk1ulBMT8eUSGDkLHaeQDAUbx
f8KwDz/udgYhaEu5bR2pryDRkwJ2vvCyMJbp3nvPBrufsIAQ+SqpvcDdiKqVmXL+qMeusHAYQAiJ
eyEJTRpAhlOTkblIFVExhSGkoNd8Np5YEixgzGAPkNjhb9TqUJPdbYrTCb+vv3BlIRf8nHJ7nAAh
R0kKx7/hQ9aiKw430XMiEh0SDCFa0dYyEb/WVS5NFfJbN++ljR2/OzeY7GahXaEsHvEAf4fTG41r
WTAXcrsU9pYiCsK9lUAi3QOGYymDfN2hdB8xFF8Ls6xzrLSRC3j3txJoFCbt2rrsANlCPpJf3Osd
lshZ55q1nuH2eDe048NKZtk3+2CgAJYVvXWXlOn7OiD6jfZp1S1wwC7mDb6qAmtOYjkqN/rUBB25
Dz+xToDe0UKXKAq1NMeATJjohbh7LSwA9XVClLo0NE9gHtWMMeHWNhB7JvTPRtLI80Hu8BxIbYHz
hVjb5KDWvxlYjFAm44b6brQiMrv1yJNV6lc7tVAlMKmy7RQNCSMvFcARtFgCicasfkUB9Q3ZY48H
n8m/uL908KrE6iB6BnsjktmZxRPYMaAGb3o4hXSvVGefe0MAD7opyZrpcGDp+r+ONt4T5ZgKQyRt
sLLKR/zmBcYMSAht7xBUEvWEe6EflzCkXicjlVxQSZ55ZGlK0Q0bq2eUzBqv+1PYBnd+kDMWlXcw
Z9d520AoED48d9LRR3LvbbkD2NCp6iwRsKOsRjrUbJLh1TcqixRUSU3IqTAWFR/EpqCYbjrjQkCB
FzmDYBn6WiQ2NbSSUslvJi9NhZEEczqFEN4ZI2BMMnvccj4Vfoq17XXcYQ0598cm8Ux3VM4nX4Uu
MYK/qlftvTKFWQhncbnzkQU8Dh8YoBXGeLvhqZHqGacCTzHSOwUEcw8N8tIURcMjzq7k1yCkK4/c
dNLCJrHw8BKANrebAoy/m/i3+4DVkHJV7u1R+mClDN7YzMRKmHMwCl39LE+lR13E7uUoikJ4iTEG
BME4h11ro0WXoy0/S+bbXGWpPyyWyPbmjsskx91F+9g9/K+Y0InHeHuHwm0cAL4GRyQTu5V72A5m
7JktqUZ4jlyBqlWZr/PLN4AdKNqyhmQhcI+6SpVeo+iArJmXnT/T+tqtxmTu6g3Bh/gqDe2CEa9a
Eoq3nIHYppQq7L9o0mp2tlIRW6aHzDXor3VMMlCmYK0h1+TcQ5JDh3N2dpXurbA/ueyceAJkJdxX
ygPPBbrFCKeplNhKnKgQzlH9TchlhV3vPFMeYQPVaj2GIWW5V9/85ZRt+i7dLYZlD18Jj7V9vVUR
kTje9F9s7RQ7DZbwwIupCfyZhiZ7N1i4Yh02yJ+BH5P2BZzM+deAQY6gON/TfFC8yYy+06YV7bXJ
jJwVGoJwwt/bVnce49OQk0IG2QKTybCg9h3ogMVyl9tJjzJ9yRjYmcgcbH/L3c2vFeUfTHMBMcNI
5eJdROTq4LjTgJtbzo6NCYymGH69kC28b8AX4LE35d8gaL8kSPLuPODRSgLuEwsANnXuojmQ6/MP
BGnfXSFN67G1ZOQqj9B6AT6nHr07sOanfnbscxRFKMCg7Ufy5pJvqzdQPWg98Trz4arxW+VDV/Sv
nNn8EiJYyRSqG5avn69QYktrgs1NL4TUsyZmYPY2hMtGo2rQu2K9+Ztp8xiqE6pfgSVfwaIJ79Km
ppy8uaJ++QMKiGfoag8QSZoBBMLjuInmkwhX/JHa6g8/rEspYQZTXuB+cp/nxPlImKySeH+aswHQ
aE+eoW7FDrKeCinYp/U+ABmhqul14gjk84AgVJKaReqikoqej4UZ0Psr8uN2fcGvQ10MKE6Ud7cZ
jvb3nJkchujVpnN5a/7DwLZUi+GWLS3xKIrLzM+4T1VlO1dns9zrMx79c/GcE2BGESp6GB/1e5a/
L3vFbO2KeJcye+My/tjfT+Y7yKVdMWG9G50UU+g+4fXpPb+CjynOj7qm+D5YNE/GWOmlP17COSLk
bdAI18pEb39CdgHaYX7B13V1CYyqFWVT7b1FM61xezm0oHV6CSnFi6VQbUh/nqK6X7Y2TZKMtLwF
7OLvXTk94wjIxaBhltIbjWk9zclNSg7g/fdLIVFjt2RalsOxxR4OIYpG/cSznSNOnX5hkwq9Po/F
dQH3+FDYcBVeZh1x9JO2oTlRwI1IUILkdX5jPe3DqKJWeivI60B8Ao36F5rdTDjjHv7vdv1lh1de
WJC+Oge/l0XvMvM1iBOCt+g4oToBqV3P+ywldEulHDq7tL1A/Sy8USMred/H3r+GvdXpOCwxJd5o
T/RK1XwIMG3vWHaHGvH36750GzRE3J2Cjbm6zphodvJCepJpxAK7ogRiHUuU91sKT5eNWKZAzOin
gvBcDdWCU5BzyOqvkqQO/A3xjcPxIvsbIKw01cY7ZsXgrgTz8bBVfmep+rhCG05Hyo3exVZR/KKl
dzCmhbqpsLr92eMmpcCv3rsQUHbAFH94hMVY1d9ZVy+UFtJTv/xlXWdxE5WUG/s3vYa4/yAnlZkU
PKZkPuopwBfAOS93Lkc3SvFNNwiCHkh0SAncUeZVMvFO9W0lcH4Bchmw6bHKMqMidjJZDpC4OE/a
yTJEnSUQsMvfpg1pesD51sAFaf2ZuLaIwZ/sgyacLcc4/wEmnHbRsY274QrRRoGRRWhPZca0sese
rdws0VvPxpvIcLFB7+r1NyLlwivpyWA59wOUVvXSsvtro2jk37LEXz2FRUpGrutVefvLRnrCecyg
8OVHJGetQNreFX2Ji2ayn5chOsJjU42sLCjWBFpggNityk5HVvejidKKnoA21FbXt3e8n3WUAx4M
i4PUkcOO9OicfAdR++P1G/3xjKtsZUFfhzbzOUuGEWNcjKKx8Qfwyoz+6YLLqMzVQVGvqFpoVEYE
n7J7VVKvoZi/i/LQy4ej1GO9KsGJevQnsjzPKXPD+JYeqPh2uaJOLhhMoclOiEoDdqn0JLweqMOd
6L2SQw4qz+hSZlv8UHJiiKrSJ7jmxKnyLeMJBKT8e3Th7FPLX51wF52TAFaA9XshwbAO6Eun9ta7
RGeZzOCdaYw0wpRY0ycdDzsdKKpbHOMKIP6zNWHyXFyq4sZH0A9Lkiv6WRaxGToD9pmA52PjkO+S
olm99VI67kV0a/O4G5F87NPPh5+pqCtwrsSJxB1T0CFjKZ+BHr/eXjCLW1nPYIl/TUMwCfzDG1WJ
2kdndtNl7lPSLNoGPOZvCaiSaGaY+f2DC4FprEtX8sm7OCaPWLGw1bGgb5JOjSuQhh593DHzYiCQ
nDf2LRQkr1q58CZNlqZaNIPVQgA7p3m111vrF+O0K/4v0yAa2Y5QfSXMLZJM7WVh2Ct/p0eOR762
mNkLJ+zO2Cgx6WmEivBASEMeruC4d7NdJhwhacZfMYWaMuQURWLyz3am2s5F7zKBUHcHq49XoYnB
l7zBmVXxrPuKorxVWEuRnJDh6rwP5Y6/5xNTpdFVp6HcfgZRldx7YNR4XYf2gNujbmqhigy1ZfrI
B38kJoLIh1CCZBBfWwzDLQrKyv8Hsj5VedKzyEc99KCJlcWtZH+2eS/A/YcD3LWulda1CH/2SCTY
8+749QRbRXkr0PviQ6Fp5upPIjzG2FN03XMHoRp10abPDrEXsw4ZMTetszo3SjmKYx0Qiskx3kf/
dTQyNhpw5VVlHxQXa6RWL2FdVsCrn5L5DEmgMQjSy8cAqqMEThtHOdqOBefvAf3GVvOAORGjNPsZ
2WPvfciy0dzsaHbQz/zbQ4EazR+s0JmDYbR75sZd5UJj0ofNjOvaV0PBjDbPyYMgIRCJJWzuhpIH
kmQfBrPQwfJzGxNyO7iAEwyJZjlV7j0tc5XlKNdSVOmMgPBrNWy+7YztzxPlpkEfmKYfP3eGgWYR
49CNhBFoR0VhDJKiffGMl48xp3rTU2Wl7mXe2KEkC2OrVp8eLNBPGEBgCN3jHAp9KdPUP42YUt3Q
KG9tsRzpMVUHnuIJm2B8db6gySo7TOejyJEwJPFHYtnK4pZWLO4PXozqDfQ9HUnD0nuLAu1q7raZ
jF0bA6WFRcCtXeUsVpoow0jom/aASjaZ1QTTQDmKbsEcmw2vDLz+l8ddC9lIDnGpaCziTqsKOKHK
yhnDJS/TTYMwnEsUy2McJjbsdlLVg5Ze1yOojdscJieUJhEGNDmraZWXS2ats83W+VenmjF98Pz9
kizkeqYlQF4o3iUHYpTy8oRznFfy6h7sxn8zdHZpoUik00jVJowzzpO62uj4zk/ToMqt5cRnRATI
oy+TBg5WyYRJ2TkxuD5O/A/OqfiatsNuXd+F2PRaWFFsBYXyaUrTpXLoRqLGkCRTTshLApYSRUXg
LCC3r17Gf9jIBYE9xmudVMk1NqKHKgwbdJ6+d3ME4zMs6c3nMPiBanGr8mNMee+8rtyjxqTtD6KW
d/JFEF1DAGl3kV162GH/f2j9myPX1vhWUccovhMOKgW3lUR5NYkXQ3AmcHTtnYHWdvktnIqtiXzQ
sZTr1TRyKBp3q7JC2hLmz0Ls8Mp7tcm6ESHhykTZhxKwjf0NJlsdR4F2I4zEs5VdvNY8kn+eqo9q
LD5NJmb6BQFatjlp0fzy0TWGS1YHPjvV7VY95QHPkwtq7b2iy6q+RwubwiLLTyshpdkLN7z07JvN
YaSjycASbRmQ33lWz/6nnjMX2XIR8Cod9n0x73cJF5JtuQ/DvOTJy3w/YRMlHUDKJwANSkampNDK
Zt73XcOaQh1y9d0VuqJvS5rfqjLh0BMyat1bY1cfEsVE/xnpVV3F2kZtFkQ2mY8Gfz3095QTmc5W
TsSoz0IT8hrN8ElLB5FNBeWTyPTB6EzdSdXSYlj3WSeWBnSvOP7aX9SE8DIYiu8n4NA8zJHV2Gpx
S0DknUM6mhI0/41RQ/8KiBfzbjGA6V0ZwxVrlUQX32PGZWHOku4/lqKrg3iie3mqC8VVOZ/8yY/W
xZ42ZWoRKYpT48fbgMN+8umx2gh+vKacwrAasTOmN4NMYAKn8FtRQHEn5g4gkQqhzY40DZbIoMye
S1iFTdfYk0oLApffzn6mX/rsgWDcQ+8HdS7zXPgxqSMjlGqT6U9hHqpTwnnElYx9cNOoD7SxlPHC
3g79mlOPykPg4l8BkwWajib2Qa5GLSlh5hn+l52+IWD60pFVtThojPBrgMxtnSBjOv563otzsBQ8
pUemrGbndD4+32HEjqEXYCKwS3ZWdsnSQsf8dFOGx1QN05+vYWZ9fv9wZkV+Yn4cY+C8Xp8hKpyA
mmmk8UinuvAKqY7yaEhgmhFBexm7D95ialORHDfFTNDM+vLizq3xOWbZIqJ95WPI7KxPAqDArE3X
7rn09iYQMJIopMudyMJYxItUOtVU6TJeaC9A7TlQWaF9Y0tdC1+HatfKfP1OfLDtgFQds/YkBkRl
zPrzpfyyTh+U17nQx4tvxhV17aFfMm+Cs3MT/gCd7R5oX9FbYT261HKgcLgAZDBXXLT1YI8hwL9R
y6Th4f5Wux2SkYC21P7xy9zect2Ul9T13ku2FKddwgL5d+fLJZGTydwo4TNKFriAomeFevsybzd0
OmZF1yHNr9gkDRPZOBew6gMMRrZvCUzAt2r6AL4C45a3FkIN1C7CayJ+AOeNZQ2+Z2e65mh4vBHi
MoscMnkWRMciW95MVs5gafVHPzFvIABVV/GC2U3Sqa/ZvNab5IWaMFlsXZsmbHHeXTnYAdHaxu3C
A57GfaJKSN5wMMDv7vW4v8Wo1Os346ZocjKHznDL/naPswfte66yDiEhbwPqVOmwzBmNUQkeN8dg
rT29wYeVxYXpxZYpjJYnC9kQH2rTJPq4cVnb0NyQTbsunZUjYr2tPGiborpR8DR0iOcjK35kang8
AbIOn6IM0pomdzYtzYK5B8Ju0V8BEyeRfGNwHLLvPfB9/w3wFx5GuVW5AMYJepyVNNNtaIS4AWy4
B2ww/oxOl7UeHItkzoy0dqmhjWONMrruyycm1PpvgmkyDLGAk2SPdnaGjvKuzEmFK6OThbuIDKja
amfsKvHcqCfvvhFpCYZF5Pyg4SpR9S+CTLUnx3zVsOSvCKpgO0ZHyjTkAav9DuZc8hJ+b0aUvsmM
29ieL6QFXoCsZjvZFEjDw7CY5zbVHroOQZ7qjDwIqRlynU2a31B2K0WxZc/0tvTx+IsiB61eCWnQ
AkRwNAWhO1yzC+zJZzkEVGIa6BlyVXi4n8POVHbxamZIawRiMVlwUI0osgJuCIgVUFgXaO3J5lhp
p8pTgGtKpopmceQhcvLPVqrSk+KXjY+qxUuulxvDtrn58MeDPuLlXgq3pF+8rvvq/8hXj1s0qV3O
8r2lqMgtrfgKN1Jfpu3aAwfJXYbzpDyzusofJhiizFJrp/c6hSGzWcQuTW7iZfnjT5YRQ9GkJveY
v0LK3f2cOBV+5KdMZFsfJYTkyd2v6igRB+F9QBihlDeht+hkNMJpPeUMhk9WFMD95DbiJmgpMGkh
RNNBVcIthPGh7ox7HmSREvb2cZNbz34BjZgBueDzoDPyCX+4o1FWzYlmMlJsOtHNvOZ1uzWlWNjw
/w70chJU+gqyUwLCBPCobrgwIv6jGsBDeRDzytNpTmAFli/SAQ5txzTaJMgzM9QzH5YMUAoX5mND
e7kbD0uKYPFgYBeSaBHcNIv2lpZvT8tva3WczypevI4nSqmSUkjaRMNKhctuMTb59LH3u2ziaRtV
HCA9kQfQesgUcorW6s5Fb1GvnCnbY5AnaMQhIGHvNtCJttSJHSxrYWlOMVzar9jJkrjREriWYJKb
cR/mn8/tG64KhW/BBygKPw5h/fZiiohqrFXeAQ4Z4uE09fghFeTqpTUbKzAD/wtqxvvLjzqeb9n7
PTe53pHazsLLmHsDhOBHcQkcGzl41Y/aJ9ZF3QbQ2d9vLK8e74xH1XnNh3KNlTOEaO4yFOaAwJ2k
UraqZGWMQa3PKuE6ADXDt1FaQx2ulUNHGsoXU2wE2sZ4/BzTGkdwQ3Tu+Vaja0qcwlp9DCJFmxnY
x3UxSSV3iKq0gtcSS9RQwntu4zqfsXS4F/bKIYta8vbJRHRL301LFfzeyeKGBxt/hUtvneU5S9ME
Zr7dsNMEY9e+5yCiI0lGqoaV9gVW6Xxe1tA5gvDtoGa7Uyb9Prhl6WPnPCdYbKyWhELXg6UEpMF/
7OQCgPG9a58EnHpEmtpzGeLa63SGiac8YPpV1dIbfX0G3dNX7UBdYgIXwNmT1TM7mqskEZ2Q38x8
iJQLwSg3H4NheG2Kkh2PLsfpWm73IiSi4GvI7HwmsezRg/nhOlyZxseW3ICTp7pRFIS1NGrGx8b2
lW1HDggvmkqAwqNUq84XbiJznAzNl5gm9d2/wEaqLw9GYSPhvu2BRPr5v4xZ6VNzx95/eAyGBv7m
y6u6j1mXasVVMlTPYBQqvk58bDqORNqz/u32XZQUlJIwkLoINKwx7m+5hvwGZrlaHCN4exodRypD
Q7hb2OlKIN02BAPWskDL+/TQN74aFOYk+ffKD/VxjQf/3YmgaKkQ9O6YUjde8ExGps3heXsQ4JWF
r2YERJ5hSmVywPt6UnUcUTpqBxoajumEjMqX7pV19swnJnsgbqgyMJFl6j/Ip/bag1cwjQlB9RMV
qqmsgt0EVNTYo1Tj+UkR0rrf1R7iyj4Fi73zqmtW2a6fn4r40+3FiW1C391stNI5mLnXL+QY/Y4E
kSl8Qlat4p84nYjyyuXnpaFH8xBpMk+UC5Ec/fsRI9MWunBmb91HYOp61m+m8/j4aEMMOseXNS79
lDUdWxf2VqT9NIGKsyamAXmcvXVRc31E4biQ4OBg3SRJhNfsMTE52BnEOLoCSwpaZzjWTyEEGjow
yXCL4ZlXkPJ1T58oGGPM07yv+qUq7z5jJ/nDaFaH/mwArtHLf+oYPZda2H3ED+ba1nB4KAQOLWTf
wLBCAPq/ZOU8AtsM/qLnYojPI0iRbNkGRca/oycRytah6Qy39O4anENerVSdTwwsWDXIPLRuHNB1
BlszfNGOn1fjQFZj2JRZhFvKqE8VWnNjxfFa8rP9HlRwJu327noOLbBeTjpSqnUIiGoiLShZ7yvp
waGG8bgsqnXKVuAjxi+ZWmkkyCg3gIoGsrYaN0IynU6SYtRJKEia3vBLeFgu+E5Zk0EyMG4qn450
w/TVxPn9QruZ9LYH1SRufuaxAFHERwVFhXAG3BpUwmmTrYb/r2qljOWm26/X2rXU4h0yFwQjTM//
gMXbM/IxcRUq9dFGC2GbAXlCYoLxhRrEoeyvWzbuWbsc+O8HmQJpiNwMC9ulAcNli0VKi1PiVOMe
K4dCbn3ypf4TLoO8L3JxpPe3HECgafywNGzskOzPeVO/Kvd/nEUM+9RdssgmuDlYD3OWtdvjX0fV
3OG2MlzDZVSLCM0klH0Lp0DgP3jjH24nu9pgCVQlKcfGzrMnuN8xU1PHz9ZCpWDKybd5SksYPvjf
EOHIQ/nC0OsPkegASAUP6F9TyfBsaYjfdSrRAELNX7LvfDPOsRsjbwuVC7j1HVCDvLns4xgTiGqM
5qhPkD7OGISBGVML7fr/hdguz0Fw601c7+dSztyzUIUCrWRNleCsF57sB17ZuAlLT/0NXRvjW8q5
qWzmr7BAaD/WIuG9iOLsveebzHumFXoZKJ3G/gqbLaoZeI13l29IOD/JP/gJ/iwWEFUJzJOhXsoB
slIjgXPCobABYfg1mHt3F/7fQowb9KPxQ6ZmeYDUhs2oiDdQdp61o226eWVPLKE+8O6uCUuCyH+E
6YjUTdAH4WD5Hr2nUXwFvDLfnh3RT2CsUEDeWa9aKS1v8wN3xlM0wD6IL+dAt4SbxQyv1WFbbj2F
De66hTf5JMeXOcXT5Hoi+P6pS3XBC22Yd/UxOrj5xiLM3P+tHp/IvALcwP0fGQl4gZl6yq5cKvji
iUW6bdSNlEqqWs36n6cbwPAQqRA2WXJjfXW+O0DTDQl92lYqeutYi0ri6cUqYx8Mg02QvXWCyOUh
f53dX5pcoexipfFZwQo1GquKTCKpldhorHHIWYjBRGB6J1BRtfLTXm+xZ+SHsCU0OpZhqqar7781
xx6/yZnRhw9w99Za8VMId6r158pQNlcxcKKC/DRqK/a0Leo+4I6yiBWQDAQXG/S16/C9SsDeoMGI
Pvzsv5L+uOJe4assXdCbaxP7XdDQFJ0RaQ3HTEzzvX+0yQ3VIqlGgSQpbu2By8IVqQrfeDxRgD1b
UKSqXgI92KbYKi0/4DRCnVfBo1Y3+QyM7fsTocBzSt8m7ayA/asy0NqIi8gEPy7mxhnCS8SrRIjL
E1VoshI3h2W6FS1Xcnx7+7mhilbWHRGMjsV+IEHcj4UBW/dW+27Oy23aWHv94+pQi7XFrPK5Vvpz
oi0UZaYf+cmy3jfMrtcIlpLNAo5rgglwF1NDKCmnc8npcfjr0KHdnmhQarpEsIRWMCzV1wua3+hS
e3l2MCaoqUrh8b88MvpmE0tW1NvyVXmXPoMGYFCNImjihn5nQbjVqwNMy31dT2/PG29PSIxPQY4e
l8TvqnDUC9A2PEfGuVYUb54aFlWRzFzjL/McMFkG2MyPky7Ppv2HsCuMobOZJ6TnFCq60NGlA1Kw
imdFivGmY8u8NvzLNBAi1qGEhCCCF8HdhhyObHxzyux6msKK8MRj6v2sm0ssP1j22a/lWsbWh5tD
OdJM7ECoPPY133UPssw3YmZfiKM82CMb6GxJ3F/vjilXoLyFyngCf0jqB+XNTIXZFjlitnmm41T0
sj8Fnlyim9MVDpl+OC6GkQVvtYKaFwyM6IE21w5utTDZ09Vb1ZnZKIswioUK8SoZfvC5dKx3b1fd
PWO8ROVtVYzNesF8cz6GsJTL4UcXnC3HNIM4IEaaUftQBtT5/NmsfPwaJGMELsdoXwP0ZQK3YiEP
t/4wtYG/w/apBrp723dDPBOOE3/4o6yMJXQc3w+T2ZAyxv7Qnxlj3N+6FrE8QTC5AxHpZF187Qux
O4r3K0MgErh1vuOkk9xiMpYYtydqYE7sr72/ncAplUN9MiTCJWl773lYe+3sNyOqOR7W3pULYYEc
Evl4nPpUsKUYfMA/rA2boxmBesx2U29WxtfHAVJErRHsuPsH1yYsKnRrBHtdstLdl8X47yZwTzL0
ZVjn+7bPoQ8+cgl5VnMej0aJrCiMjULK1Dw8SfAolLaOs4GeEFrCflPW0VYYjibuBjScpjcXTCxz
asFIyVmXj0YWjApMjcmwLyaKpscmrR0s56oqfRANo+NAWUqLQuElnL2w0CiAuJh1HjHZg6xice8n
jvGAQjnqWKGmYUFdaDh/rZgzIlNxXMzlFJP6HPhf2R2NQf9wUeudDsghAzpjXT17GcSJT57ldvHU
eiikNy5bsfHSyR+aCE63lzMHzm4CP5dxS56L+UN2PXV8JHRH0cSA6aCetpPFf0m3fZk+aEPcUOk/
Ny+fMKEAOEg7CgYfADRmbdU0MnaXTn26e5IkSfNP2n7pbVJv3KDouhcsvOy9OCn/9bzkrFnWP+ql
d8ISEck3M82sKnP7hxznugucKrGIZjxhPXsorx3xZ7cG6NdxJ4SBvgVVZ4ynbTbKvJVF//8CC9yk
Hynq8QGdUYRnyaLwTQpb0Ue0Mkba2u6d+jBYH35yJpxev9LZ3el75EIJSU0iBTkwOFs0qUdPn8Qf
44dVPy3cQvQ/mlwODOsy85c47AJX0HbxTHKTr790snmz7RSiUP2RF5p50s7sMRix62j4YUJrZFpY
5/Ag6lic7X/mwYyawNa2GHXuOvYvGXrsG+rg23VY88rlFhLEIrZRKzc9hC6zIXgtVJLpL9qlwQAL
UPjOcq5wSaXEi+gR5wyWCydPXknVApXJ5wM0pQdceSGEwNVfphpMy6An+QilmA3ETS7AHxEpVzu1
anGjKnGZ+YH60wOzUkUUOzEacm4txlQDUueUUun8NdnY9ILBHr+/uncbYn/uhaHR02q5AQngMeCO
Yx45v7AHZww/i+XYkTD5ee3GMmuniWrwlXx2RSMmatHHdWea9RNbfIkCsRi5tNVxfPHY9L1vntFF
9Zhuf/PzbA96gEd9Gc8DF0y9sSIJIJyaykrRReY+DcUr0DyHHzyyqEau7o6EXOU3UDuTxuPtDsGj
DqknB6oTholMzDw6DRV2Fl8BQ9j26a9T5KzCvlbcC0kRF8RVDRc9f2pQd5j2A+tohBszV14y2jPe
tKwV4djq9dd2s6sC7QmKWmDHMWzzkNbGfgx2L0WI2UKRpIqvxczNIQ7dPH0qSHwccAst+Gv9Jle1
QesJnjEHgb95JFuCs1r+qsJa6KwtKngndOhAzQ8EizmsdGuuiPTXOSIBga3LCy1ylVxB8IHdwY+l
J0Owk0VQaF34waTPmJPOaVa2nrljv88i7C+EypDvKj0yy9+BJboaZd1QrVmmA1zaaEkYq3ePtX8r
mri6WXuXXBbm+kWnnDVXwycfF5LlgvKyLCrkVEdII38cU2daIs4mXvqbXqOdeBCNgNuVLHbhpoOe
DnEyu22hFRBjoVo+e82PG1g+pedaxn/a96FHHKayutUGJVIz3/lwtqquIVjHhCwmF+yJtECifbB8
47aXOzsF6tT58Z30ZltNw9lNk8yookROMH8GfxAOvUmGApZXk674lsHoqezpKA4KNGurOcvAH5wf
XrDz5GxnL9boafusL7PnxW8nTFVxDFixm3Kr+Y41DguId8laEM6KO9h3/7tFYs/jVrtOVEWPCgbm
f4IpYPu5SR+zuaAeJOSFSDtYfqd+6uPoH0gIp8Nwt3olAKbboe0ibru24xn7477wJJ1wmifoh4eI
hLk7Zq9ZsC/ONx/s2PlZ3viW8B8j+4DhfoGeHbiV0ROLqeXMSax/Mcqqv/PB+rxXuXE+n1x21SnS
7HvPmqm8fEUDqgIyQsYINywddUBsppip5a2Q7TOl0oA5F2XHnxaH4o0ez+6W/h4Y6usTjXIouyQu
aI/kdhvIc47QgZow/AbOWtNiGKFXGXJsIsi30AEn6ZVy7ljqi9IcvdEMJCeSNBI+5WLGlkNV8UAP
pO6UR8FKZmlQipZjcu9G/xSe5hGaXmX8I7UrUGVyNcCXwwK+LoPIHFA6voc/dfgRXAGqwki28z4q
yJCpYUEkjmSz6Fk5D46AJVHWi518A/zcvpeoE9qGAhLU6qq6WW5uFXXp1MsBMJAmWhIvNI+CVaTU
MOuLnSsSNgqp1cgzSTevS+d1atT1BA0VmLCNTRxEh/kx+qG3t4/ZhmslgmCngHH/4QRNFKA0vAO6
VbLYtNycNaDlPNXIdb51/vVbp83fBQM7EmZ02yIdFiyKMk8Y8Ocv1UUlm5bc/T+wxy9504/+4eeU
qoL6uTUJeA+TaQMKZMzI/tJQeEDsdAz9gAX7MmRDl94FNTnj9HJPbBZJ095iAitSAHSW6AmE6F0g
Y1pCU6+X2CJlCWpNqy0DawyZ+vzpJOSM/zGHsrQsCmTOYFhObfp5k40hSmPER+dyzTB439j5lU4+
WCM8X4twZjaUt7BxmJcZ6YIEatBdVg+kWPQdrmUxRFx206bOZYXdluRZETHHvNy8ayovsBpDbNne
GZTTiUD9r17usrKzq1Iu37DxDytMTpapeA+wqM115+P51EpY7CUsIhJfPWVdsGHplfxVyvDEG8Iy
ZJ5go2P0iemId54zx2GCt1P3ZlDBTWHOV7GlhjMbjOKPlsR+CAiLODGWt6YuVMiR4QAtzX47HFxG
2tWo5ZkXn67vmQMDMiYOuEmug3KuE3oAl7m+mhyTlsLRMvDBxc0fcsBp5+ChMNOJ0EOImFb3RQgx
flvDGgak4T/jZ+/BiYVwl/ig6z0ME7UAvR3/LHhwfm16l+y8hYE6lMxYei5TtCo8M5DEm+WTBjaB
gG6e928FS6k7Oibt/HDAO4QvaFDT3mPfJYqUGoL66wcIeGbdTkjcSUUth7GnrIVozuKWtHCLvTlm
1nBd4J5pf83Q+77s6whKlWpUc93pLBZSZGkJ/YssFFxyvXiCrQTfs+WtOtGKkkSRd/hS65ljAzuo
+Di4k6iZHNNrCo0SOfwRbB3m3ZUOwUReRgNe4MMCVNM/Qs8iItliymUdxNHZfVMWarXSYs2QHUaU
dcqSoYarSBA2Mh0hzuzMyNNGJgLJqXPH7l0g28n+4RbH8zkH25SSc87NLc62gkMgTiCbOP1Gl1q9
bo/FVzCH4X2WijDYOKksdvdOUkfxxrjh9uEe8BXqHBeqLNSNf7HQFxjr/FhatDlJFTsofLpwk2Zt
a6nOA0b47n5uniPBckGYVPO3CheplAm4fuZW6Y01DAI9aYCwf5F4dYS0hmENO1IORvJ3xHNaz9kB
TA1Ey6VXKcLksBjpOCbrB5upTPoRXj54oEDzj9uGtmiylI8Xrhp0FwzrxlkOxFJGi1NZVGgIlgbf
kDkoXQAUxGfKslLD3TRwzKPsoYkxkDnnLkDRTO4ZO3J6j+K55WNV+1CjmN3KeaujcapyjuKnQyj9
Xo1Tbym6lx188u1Il4p9ltdup2yUmq08OMVuacN68b3sb+i04LQGS+TxSS2N3fzdUKGeXxGDjLY1
vCDr7CylnRw45fuMi5r/sP7e0mA+XT3FiIyNQ6AeCmQ+d+3J3RUYYVq6GSqiZ+j4wUWG/jJcFNLi
vJAnY5sVzazFoAGKo/Oy3S0YFPDUWgt8re28QlwngbiVEWPkKvgrSQ7PIrtnJRbK5gHQFb1ff1Mk
OyI78c6HQPHnUEvmNzUGvfMG+pwE4psZTaUOrW154yR8G4AElf1E1V9CZJ+aT3TMffLeSEB+srYB
BOn66k8LNHUJ1D+X2L9+DUubOliH64/pF3Xegal61Nvns4eztqpLGRkx/xMqQkDdELC6bGTj8lv7
H3uY3wfnFZ5qa5nhOE7Gu174/eMMk8eM3ZNxmkyjPN70Yy2mLGKcfhA68GTRj6tYw0+t8icvmC9y
mwJp4ycanqYF/sJvR5D4MpS4JWsBPtN3Lfi+aDsoBydn9kHnAMG5FZ0MTHZbtkuygM7ctEGTtUx5
QAPb2fJ8lUI7A14hyg1ZGvEzYQO+DiCX28JrX+ozMNHv8Y93t6N6ev1VJQQKUs5T3oc7HS5XgGBz
2EJk5p+91H32xWvetXsS+ku5oFM5ZWkAyMj1p7EaVM6tvSBpcUXeKSi+g5h3GdRtIaV6bi6Cey+q
FlFDxjeILf50Kzw+xj8s1LkDPkAghKQ/Vw9xcoS7gr0kX1noaVhSwc99CanEgE14qL83In7ut6zn
WGnRKW5AhsnilmJ/aoC3KCw3elDqfSHFVbJVi3WAxvwJjEUjlV6fJDh71Ok0j5tSUZHWx1UhvEX8
gOEi4d6MN+RnuPKUlueF66C5V4knqeHdx/FIijefr4mPgd3f/ov4ywacoqsR6HiEgLLwHXnomRSG
PC123Q1bhQxFAMopHkPsX406FT9wkBqfiD7PtYPqqENFWawVtf8HaIj8AfWHZOFiZCtEW3sfRVcP
5xLCp1RVtvXsU8Hej7SYKvxzivoLg/9OhvEnun6aO170/YISmyiouEYZRejHv9x/4GWfEMZhrE9b
goPUle9Pbu4OTuMZUf238r4bDyPc2u1tOoeu0bdgBQXWmJmF0JHMO6C+vawBfodwbNT49DB7q8Mk
bEsAYrjyaJK1oS7eJPw2xwRiW6V63LEYP4lXBbD4PGhMEKqgkm0NF73rhruDD0Vgq1+GXUbMJNEO
q3JsPhFfxTujzt94KK+0eRcevlizvMRWGwKk+rjFey5qFHf2tlWcDbrM7TBR5h/bRix0EaGw7ur5
CjY+yEAV7T1HDRtVsmRO0mCCtY91BnMZrlNSel8wRm64jaVQRCkbrVk1QHi0I6YXM5NMvHSv89l1
hKXBSt6t6NntctY7kZ+qOkjmHJLGwVzVCmgAxsNMZ9CzGm2FykyG4Y85NOVnxhbwZ42isRbDbjCV
OEJhWffyRaNiqyF/7FbQN5rk3fc3Pd2W29bxC+a1vnaHkVwcEC1o9bt0pRsrn4giJHmoDK6mpVI7
L/T7+NT3NVTpJ1wD4F832+rnuxj+wGNU1u59DU2m+I/XnOBmkjBnvpLlp2Us5CKMfH2PUgUUD6ot
MkNUxni96ZU79BowrMap86KAYaysBrRiN7yZmMqw8CAZMaIoYnP5yjiZnleS+35NdAJgRirR3/j+
KFzj4JuUox44cs/BkBk7IkI2MJxnTxK3g2OQEefziV3Wu0HmUIqPGvdrrsQyUw3e/NsOSSk+aa1E
B+IU7C+hTlPucZOQhUYRZtdwxW7K5Z8sUJefjxMc9eQIRqTEfFKj7snIRSGMgZpPdXBX0RVP0Afx
MMiTVnh09PUdzfdwPZxa+dd+V7jsx8SWgsWOCHqOpCsHXVtq+s1BM7Rc+QamnyCb7WsGZnWB41xd
F83cOxEBW6tR9iVBy9kOnM7G++gGJliosxKH5/2VzbqnJqjAM9SD0QMlNGH9r781IzTRdJ0rmEAv
u9Ipgk6HodXMmMk02Q/+EiFVhAvJPDv7Gs8O4IbyCeCG6J6jwRhelirpKk2q42P1feItlARmxBrK
uIh+l5U4KcFQiOP/OFAbz9SP9ypHElKxRG+mMTAR1j59t3ETHD4i5SUbl1zLE8ibDw4EpNzc+70k
dNBeVg21npvrFoCci5sjVhMwxFghX8fyd4fN34GC9Z89YmDPb728BS4PbCgEoN/Q+D2TgMvjuRm+
FvIMQf9SggS1hSbP+Rlft0cwxc6Nd26BUEiRm0qrl8gN0aeNmpYbNb/9seihb6NdsS0L92jjnU+M
1AAIZaRMy6KABqkOygXFLR9cCHBrhuDIqHUUKcZz1wfAV1nSEnH53b/W6utAehrbIaGDHND47eRm
Gd0gKwWNpRD6v6KXJsrKV0PUPuMvGKwwPZOrXEwVChb5WEgSmL+dpR2U7LEiH9j4eZd0ZTeTIMfg
0n4FNXIJRy7yQbYNA4nc3uINByWSIPQFY+ypzCsed1RW3rnT0TVpShlR7BACkqJpWRdZ296nDp25
7cW+O7uPZZdLLS71qFLCz0nQQswlZjP9GHSCjlhn0sSiRnw76JgawvV2Zr9kPVi0Q16MGWHUGrJI
MINpBir4gNM5AMO4JyawnaQTxzoZ05fg8ScknYAisVUEdLBqiy47wNVo6rVAEUomDr0Wne5KcoO5
qDer23AEqmqGnC57DuiIBgjl9R/GZi2bGLX2pG1kngm399MLB8MZ8cYu5MWWKzLMfloos1kcizZ+
DzpGASD5p6k9C+PcLlDbWxQClLgcEH4alNfQxt+UQ/dj9g7rsXG+QTywGgVXZajDJqe3DdKK8nwN
IrQRzaW5Gu3Cqyjc3DaxAd04Cgwc6VtdOFmNTIM+sZQKWEpFbW9vjmmEORpEUNKqMP/Jtr5eNXcD
L4ajjsfTftw4bh1sr9ZQAk1gr1eVxUqFdjUkrabo7z2ysLFRIPJ3Gduy9jJP/CV+XBcu46x4U/3u
bAhvFgCsJMeKzl8xuVWsbU/jEz74zjbYAtFZ+r2+wDFJUo3BdHTn5mVXz0KU+DNw+c8OgEWyj+KU
tQOnnhu7AmTMtl9JsDEwPPsgkF+7QHI5NsCc8KX8hXDSilZ3nX0IQ4mNSLFDc6QzRNrJtvpTgcDY
ybCoHIaxBXDyqW/rX4mq/gVK1ETDoSpImKwQf5V13Sxm9W5FGJu655MW8QjykiPAUY0bzSeAaCsP
Wj2En8igkBrabFTuk/YiT7yJF0ZWOQaK5vZBxEKcdDZIcgKNgqMIfQe22QiGJLwxs5pNOlnYypx5
f0l75ejwiNKZyJGp+1VKnWweWn8zBU5qgDEQu++pZwzGvMZ9vDdAYpSWPC3elha7fe45TWTlLHR6
tMLDhuWP15UOorn4OYhSKCEg0nlKazk/PIa0Gk5EDGUHkkTeT6zXwiSWW+LNR8bWajtOjQR53d0k
mYwKYKFICBiMWspM9HFnXy7daE2hTbAxdvhrwBOjI0VWf6XpKL/EBOLWcPj9jh19ZC87TG3Jhovj
BCI2hLm3GfIahLB2UU/Y06RMLPg9LNLHS/FVuddRscs1Irt7ckniXAzOwXS7iml0hKzHKT8kPM9B
JwJXZwMHyIDVoi5Yp2ck/6ECP+Wdg5CFUBHhavKwX0S8VT0IUYjJ2UwIn5yxCslHCFz6x1Ar67It
l0Aqfavo4kS8pIImmxjFJAMWJohC3mKAhYT0ckQuwAyLK/HtPjJWRGK6reyQfPOqCCDLz2MMzhi2
XVCqrDbjdl8N6mXJFyhrrdb7FIjUcGOz4uaVLoo4FxvxC4T+KG7pK2YB4jYUz84FC3/jh9y0ooHG
Bu4cJTuFtcgENFGqyPgIUVcDaNc7LTq45xbNywBYS1UU9MsY85UhWPO//yMGLRi8aKvDb/RDCtH6
NUvQt1S9EMikrkKzlzCL9S/LsfJWxITWY7ihqa2UOk07cCVJocXtTr5ru/H77Iiex6B1Y6Gd79RD
ALBhGZZZsAe+Cip3Rp6gAz0LgaRbOjVbxKdmejV8ipeOPCugMh+AT+CXhxw5hrQ2PSCmEPPACAvI
nZHLYt+x+Pw0gdemm2fZ8sbmi9T/bG7GPxD2CTKEncU7GgnFLHFyRjcdBgLwb6HltOCCIfpkPm1S
JHpAxNrwVEnnp7/RajZ1WRWlIdTaoe1UT6fZRWLA8qZ2jrICLEFRMsO4JYWgvPumkDxpMhH2bT95
EYdwfppFLfSyDBwl6Xhr2eVgDsaeA2MhIikJwRLmuEgLPFJ+WsfA8aUroP6+Oo1vNCuRxAUOGMxR
QjG7ovkaKLEWmbwNl8oDoiP9jMlpAAo3KHII+ZUjS2V7HFlNN8Iqsz24v7p16MhJbzEkbCM5zzxA
OvUaMNOH6HJH8W1m6/yoXKtB2qJO61tLr52fCWJrKdrazb9KcXJTuqobp2DW5IOJWaQ/HUQXq0L9
Lq6P/C51q8G9cLpWNLa1zlRRWyrymLdVUVDGu3x3j8zS2rzjhR2bR8ZhWGPDoNTOEXVSZiYEfqOj
tJrzBvouVss9GDMo0e965lP7uQoaPNuT1o4l/NSGkQnPAw7eFjMzoRy+OxJeJVY7uc1Z7SZK4x5i
iM4c0bhMyQCmICrsnZrQiJcF69w72iJKHL3OVOctVL4K6GQkIV5PODmHQpo0AQlCCjNgCOx1dHtx
x0U5d8ta1N/boUI8V+o4cDA7Sob3zhJPHKo4qi1l/N0arTYwXXd707HU+VCbwtjiGGvOR+cjM6/P
PViFOA/ukIhXIgu6XEq9ntorViGMZl7+M0ynTv9vZOTxjNMLqlxIthQaIBD1pxJYYVUmOpWJIleg
UXp2xHIElUmtGTf+/sLY/7Obz2/QIGf7HAS/kAlXND4C91DxVnqtdMOtozEL2Is2ViIrOQvmEhkF
cpTaAah3070TZtdlTb8WI0xAer/qE2ov4Sqf2ZMCFhNy3R8IgrRqcZh9ZjkG5ilUvvu15cxVZWRJ
leht8a30m7wLp/phbB8MAqz3Y02TZKbN+JpkXo9oA7fjPZ9UU0dCQEedF/srjGHnY3U8d4MxJGAR
aSgtfU30oAUfH3YSj0MycPOiDiKtnzPAQvALN7VrxqVI6yRf/8ipgQ0kjYrPS8pfSfuBA8wdiLLQ
haE44+QW3pt8Pus6dFmXNrQFxWQMIrsvTFs2NHzlM9kNWJONbvLOnbjcBzXKpEykhcknMI8Hq5xI
2Z8b/wA+OIfav7ISSWlO059qpsi31eB/95MsdUEJL8MfhXfRvWe85aFhpIGHF3J7zSPwjYTLbXcA
Jr5LftP2gHQ5ra7o5oBhnt0MH0C+yb5l1sjsNwmnjXH9PJU2B51YBWaBs2UT9YfbqxKhLkmRk0ZN
h3ftiauc+h3k0AXZC9Y0YRoN/aP5AD6ieeb9ctZ/r/38n4gz/B3YWnJKY58jYq9hJFf/oZZOtqkr
Zn6oNB2HhDDBy23oLoeKzpelkx2F8z27TJIaZsBykmfHzvIybTGYjqOmYZudk1kGJjGnFwFfImdM
URT8W6cPKqFea44MU4sb9/ki1JB6yFcy+YJxhPT9aHn63OoxKaaV2RV902iUgtbun3gWmL9otgTq
hGRkJzgVNifZCvfhJFfLFSjhOJGthtDHxoTL44miKY3GGUdTluanuNqcTCe+9aggX75JCJsZgWZf
i/ubMzQuB08KyIg1o3eYK23EcMtu7rytTtNC4/DmmMQvecHRLI6n3L9Ce/+U+r3elbAhaC4miRSu
ffw7EwLhnCGxS1y1csRrSX4dKqFO775jZBBEpsZ5BT6PQfcwh+ZzD1k6kEoyMEHv5bA6z3xejKTA
X1pfJA1ADWd8rnf0PXIaikA+c3bAHjN0gSuo403eitazugWkLQer/Lpz0djDhPtjHDVO8CkacG8u
jNErNXIQnQ5fej1YuTXCfpxUBSogs3XW9nzgZVi0NHTzS8fB2a2bNv0YYaFLqik/4bHTB1bjaxKq
ApjQZObwIHbM65AWl3ouaBDQcdPw7Y2qO3mQD6xrGT5MC7BGlVbz9FQJ4dPQIV8+OampXZ6cWdpA
rmu5YoOJyobkQ8azJ3YPa6ZtJBUD3BUys7DnEriLgPISFJAcVU5E3LMYR9MxunTjQnxuwJ+/QJyg
XX1J/y3soHzQJdhcapG/Q9HpD3kSvWoV6wp4a4deNBvnjygv2sB29WHmstEIsbiCWDZgGOxdMuLD
EIYJnq7CLHftiBYfxpYwTEuLwZ4DgM71v7rXBh8mj9yxKzxYaocXWLcnC3MN55weL++WBlX08mER
bqsuz+KaIZYf7JlVGHH6QDKqmPPazuI1kfqoBEywzqgKPoGISV7s3zZzS+mpeomJ0g7a2H2Z0nMB
WXJXXJk7G8tk/joedOzgtGEy64R/7AU0I/2qtpPlSHwH376hsYxssf3fZBluAuPy9AGoE9q+Gm+I
xBNoZtJnGvFeawfNUu1BxP3x6NYytTwmDt15o93uYgn5djVyBNMIPN/blvWOPa2EJeNrFTcpITm0
XHHSKp/qJwG3D8b6q8vkdbRDRXYI7JGY7/2008us1AOoh7mmoqii79IID3Ara4zqM8q1erhewthF
xovunlKE6szPtA3+j3cN2RAoFwtn39lpt0DyvocseWle1QcKnitUOeCFgNmSBW2UJzVunQJU0QQZ
ulSi54aYvCmejRwS1xKP5fa4Di0QGsUb5SiwjtcgUD81YbwePq0bqcb7ba55bQqooMLsOmDfVmXZ
XJWCNa1KjhO3VP/qT+NCJxeG1u756wExCpEklqhPLTkr6sucueqh7N58HoHoQ8I+Fg9uaKNNQUP+
kZvalZv9GbVr06JY8cLXR2zva1BDu1oj93INm38qRHq6Cl2VdkqM2+2+OibkWmZCWCfTlkl85XY+
kRCQcaQvHmfmt3xNMrozx6M5HlIsb6OZ9Dkt11qvk7tqxX2GYxGRuEqvt4G6sobkPMYsYF2FcYya
I3ASYO8vbEHuJ/AOZ+qTaO5WgtB9p6MTki2LLJ3fCThH0CePhFFyU6KRnr0EPjvUpMvjI1rxQn0j
j7y7sqbap55ujgzcukgja9FSepU+9kf9j7VhoDS8vmq5u3LW5pGbpp+7avn/aYhpzXOYJawrfirN
VGSkfNj2qOHxywTJsPjo7N/j6gX/He3CfXOv+1Nte0lmIndya9S2inFWzHc9qk+Xvqii2zzfO4os
k0JzyjFG6hPU5ykUHmg9RzOPw10ISv7Nn2iDXdAGOeDDpkGwqBUZ32fFXansAt62j5Lde//TKiF3
oWH2Z2QTjeT1CXsB8nRdjfgXgbYmHMra5jgzEmwTk9DnlB/A3AQ+nvDUXKO6KYYin8GSx8cMNuFK
Gyl4kwAEkLbzFFaE3OjpHd9mn+ASmjqcDe3hNi2+0vsAX5zPzRRMx1/dYSdI+vB46cMUUqRPg0xP
Hu7+TtvdjgWwBIAVouj8ieBTffYcmVACgDn7b8ABnhdD4Ubh9tUGdc2doFop8cwtbSpaz2isL+th
Qot1a4JRbzHopprmFIuCRbumytnvI/Tfdsmqz+Ho2MNoNk4D3jzrOyuSabrVSHlpJzfxQ6K3w0Sa
g0pv34M65pCXdVe5nHY2Sj1FaL+JkndsAW2nDSq6xd3HnWlZSCFCLqDLEK36SAg+e6CoYx47qqSY
2gWiXcEJKGV3AyFcmpnHaLiMsClIjdecRfr45l4Brv3Gx1lhtsC4W7XCTK1Dwk/vXTlQilARZZfH
tjIkYyJTJ9iS0nq/8fwYqrO9YXbIyqhBVqePYNHby/xBS7t7LkR7vbr7SypTz/85omkwyLPUlA6K
yhoHcCOpV8Rswzfo+KXDoYOory2Q3GUecTG0q81lTvr0r41aEeAD6rSkmK95RPR2/oNUJTbSqmuG
duQYGeKpXUryg20lIf83TjoRUOyguJhsgBLqcTpkC+o5sYsohjrZJw4UtZ/azTcqlIMA0KSZAWSF
zFvJnp5ETI9EagwpyNWNaG7A4PxX6QFTl3pEmSylrrngL8W9RiXW7Ch6ARVeWZHRQ9p+q0f+pTDz
Z/+HGCpaNs0/8Aci/jdYt95nnM6q3sKoM7s6cPFptGZHsnWgvwmOE2oqN0ygpWVbK/I9kbe7sPHP
FcNFAbS9vQcmX5+bM5my3fVbbxGEDRYAp+THja5xnxVhxvkBKoU9GoaIZ1eu4vmDFv73pAdqqCp0
F5Z/LZz7m6xMd1kqZfjYrV4CNl3ZwvathiD154Y2hx+jAwKtwa8DHswEpd0b0Yg9PfAOofs9ShKI
GWS1851xLePid20FuoKt6QjTP32zw1hqpGoMx6ktwcW+HjiDhrKn9OGC1GAH6tF4KAaBTiH3yvqr
8vOWRhqt090cLQfuSzfI2xxcF5NoJDugc27f6c4bCgFusZNCsFksisCMwTlr6z46v/HDabCgQtjg
cngNU2e/8M6SM+dhgMnWpqcncSUf7vm9S58pbaZBxGIHKru4/BFDw7OTodnijsanP9mwknsPXzQ3
Wr0/n1V1XvWZlQX3Zt6NSFKBObH+8wadHQNXQmp/HUzGJ48Bc3DfjW4BcP/Zntp96i2OpbE8OizW
7xncu+BfSoRpV8LcYEYvr1UEOnLJ19oE2cHeDYgmDf7EUA7Ks5tiYLLkmPkM4oreAlwYXDxGClRV
7lj3YrvIv3XnoeNVUBur8rmDdXhv4HkKLxpUkzurZiXBcjHsustT02fBszYZaSoVnJF3AxQK4MXd
zH+NH0HnZ/VU0UA11Z/g8Pix7tBAQ8NMi24MBmG/VlS1J4rgXGS0VR5uKJk/jM4n7ynPVJVuckF4
Wf5DGmQCxM+ZGi2LwuGPVcqr76RWXeMj7Bo9gBIFRmoMWwnrg/rkWzCE79SkvBGdkVd66GFc6S7a
HJgaipJfzVLJq4gDgSO4exW97CkHowZbH3Tc3kTRB5vuVqTAjVf2oIGWlCo2/R20mgSoW7xzPzk6
HDAXU/9Z27+Q1Quv1bqXN2vHDgrL1RvhOGEYVnDhB7fgyXxWMzYbQogJo9e6ubh4KmrUvZCvqgD3
76DGNVviRn2kYKRXAz1AjfNFzJhbmWT8SAauDfU2QnpC55DdiTPSkk/itQISrdtuKfkgMzapvlTY
UyQ/d3NBov8HL4c6nix7buaxrUb2HHxKRXf+pEK2eWMF0eDSRcZ1pb3NUql5Bn1CPW6NR55XuDP1
bBBfDpraQaS4GBYkbbC49gvo9lHsyVmz0GkEEJStr89/ocxWpL8+j4Xpi1GvOFfhb7oAnnairA/u
ooHs5dro+Dn98wDeoEPQlvPv9xRDAWFTJHSR3HVA65St7vNc35FliKF1k2jRJYpAU1cYESf1HgAv
F4kYn6TSGowHo3Ih9LQZLFgi9cLozd3P9MJZ5jRPyT0vTR+dmCbZHnVwT2r/14mfIidPKE+TQXyD
sAhMZLe7AJyAQ00yAph3BFEh+GgHrCoiF0FYJexf6BvkcGQ/dl5Bn/HixByAs2Vze7NDz/wNeB/f
uagGNmNR4UQ8iWLOOAdOaxloX/HC/bCqkXytiRcL4goeCmD9EqXgpkAEYlmoZW8knPsuR9HGrbAV
EPGXWI0TeAc0cgkTmq9rmpWT9WsHnI63TxKx3/v2/guu8teNymm7NuB9b2jtjo1sE69JO/w+J00q
sxm+6I3KmndoeEXVl+8apskmQZdK1huqqF2Jw8DavGk6Yx4cweJdQSixyc3koAH5YNcu8cw3hhRe
aQOu1m0mlayM7GkiHypsSTG5wJkaMa6yy2UHe/izia2+LDY/LB+R2Ayo7fg03v4zi+Ekd2TdOB5G
qkRoEDqeDga0JuvUQHf2O+yLbGTO8OvRaFdxiJEn+6Au2y7xdyuMptMqYCrnJpp6r2Sqv2eBYr9I
K+uLrBVHiDT7EtJnadKhrSPEGxgkjo70YHYBXgugSYX2vOEjxnqDgv5HyxQfoJQ24iQPb6TwQI7h
gJjlm8NAn290yd2EQi0aSiJsdcAsMM2mOev0ItULP8SXoQy9vDZ7BXMO3EyTPzQikOwJAgcF12Ue
kP8f2FuB4Mp0v5gm/3QyiwNR23C2Tt+Qa7U/6C55RMKoISPZtP54FkpU1dTZit7spcpfuZkwvOyE
Xi3PwqIIpCDESVGn2NQatVFj7/jcfsUiVFiET6vQocPfccdgfrC4SV1nmw/xZ+68uRgV2KI9MuPS
YdYV0N8RGPXGJlsIAbdSnds1laJKW1Vlmfuqw4sJwNsh8G5uJDfmpyqUvx/hb0gVwWMtNX/ma0eB
TxgFVTq4mNTGNDHePb+MJpgnMs2o1Fcl1ih1mSJ8B7JYx+rWPke3reaPZ6CIJ5zAMkwrcHdFZMxx
DfnCQDDFte82Gk7odjF73GcnAiwMMEiVXszw00+sYQ1b+FLW7ZZTq7A/es47oDfZieR05pf3nynO
EG+olUkuBvKWCGIKsl6EwQ5MacKULt9FqW2y+LdVEjkDGPJk1EYNgMZkCAVv2dG120YbnnX8zhFP
ECNlYxVibr/FfXXheHWVPu050P3HN1H3JpiWC1D4k8X4Y3u7x+GasiWV0dqkrmaY+k+01wcMofvC
j30uQYtfbrs2iwhEr1wY8u5vJXs3M0CNOTExWz2LarIUy1gsxw4Z6lalNmwwDX44o8TqaEeipxQS
3N4+FiOdHds0JbOQPmGDprjrbFTI32hNaOE2GR9uiJ4MeA32UYw4GbRnH4zFlJ5tl7whrLjgw2Tt
P5ACfzv2fS3ScdPKegy3G5MPLrc+/oilwzpEgF8J6Vo/6zd4PaEPBa62ebV/XAnfEUTqVwq6eUY8
86W7JTx09TrDjAoyuzgAf/HLb52iPHNfjOXF5osvIQ+2mySvH568rXkwLSkNH2nEbvG4QLu3L/vA
5L5OByd1N4Wpf8MSjwi5tg3VWxXDiYJT+xMehRn4fqiPEXPkI2DFjg+6qczWpyP57t30zWakDf2O
8Z1TBBrEeUl8FxZaxBweQtyuIM7IeHG/ki7SmQHq9HJftEh1IBDNy59EbZ+DSTLjV8h4DhcwHV3z
DV/seu60axV5jq9mQOtiFOgRhiK1jQbY4JUMwIEAGIFiMu5wAjJJvpCeWaKD9ugRBcZpea/XUK/3
JhGL3LgNx4Xq+plqnxthzKevPrz+7n5FXfS/BMkjT2HEGE2MRPp8MTAdLgR8t9cMwcS40gLAAw/B
N0bH+h3rRKVIWxsr4nd1XFsUNEsN1dg7WaK4lp5NtKNwc4fslizG+fpwonxBbCfI7a2Hc4Glxu0j
cxVQGnVD2z4cJ/SQfy6Pf2lV2KiDl0hPPujWV5TVwuCz7DKTXkrk8OshTMezfw4T2QzZPCdF9ZrG
XgmjVppWPEs5nRz4CjsL7wX0vE7a1xFSSayEZS5XvioBCUmE+3w0g58QJDXYphAg01+qoxfKnmy+
ViSz+aDpzOgqVlxIQYYtuaYQPIj7SEY6OovLRJN/NxzoxqRWfxtUdGjwNqpHMBBkgwIEMRovwR4s
RRbALK320BdhZZURvEXfSRmi0HL8e98jcCBDc2lxBNwtOJ4Lss38uNPoksk82PLACqDMgdbh5v56
fW3nWh9XX/PjpASb/rkYoCPL9/ollWIxqulE4xMmTt5F2CUzA2GLzw+LdAc+jKEPaCFF+PG7DcnY
XN5oF9rv1LtTDa1wKz4mPR8YY42LzxRD+TmANwXlW111WGNRMsCZTK3QqsaN+4XaEC1lG3GcNDwF
ja+sDBtbbxTmncvgWQC25xyhzvJj+S+DvCTDds/jDO2XZnZMmnIVeyCxyrQp96Vu0eFDF+W97Ul9
/VKFMliOSDWvWLTLSPVICxGdEFVyiEB9/WPy5JH5TFhyyOPpml7lBFE6OsYUcFFSrAn/2oFbMg1K
8H3/GvI7uYAhAfEGnuEQdBA00WspF6Tz0M0MR7MfBMrIX8ExSG/uqAC0e1gmZD5tJjK+QEe+X1bg
ncQeVITJtgjybbYCjx9h/2VjvWWWlOE1Umj5spk2D4SbQAoeQ6qMB2ZGm9dy5f/VlrOSJ5e3gJYy
kseCYYS0WrtPeQcNI4gAI5qmwT00UpM0Zz2amLU+Q/qKpngppnQGPXdQ38bR4nkiT65aqBEiKJgg
lBmyL5iCWdXT8VxWksFnLP7PSw80XPeci+q540bQt2m+wVtE8DRibvdf8xNjxIdS4T3S8NMkEToU
CnBDrGMgE+WeRqxCW0m8GS/jIZC+LYZiNm3wbCMXSqCn4abBpsi2Dy2U5iGj4nxZliliShPQui3q
2xC+HzbI+Ye3ERlFcGK7JAQvp1n91VmD9D78dvlH6mVi+0XFqEUdzbh5B5dWyLWxnXvCFojXYS+g
HLssIpi99og8gSaGO/BPeG/eV79EWctRvRgwiZ9KCfBE3iUVDv7ccj+xA/SUF24tHsznoORM1sFj
zHLFH7EympoyPTHCdUZgP5McfBB0PzqITWRhEbrdXKn7YrJ0/zcpSXaFM22l4Ru7ND7/D6Wa4zTb
N+dfFx0gWQYe1dK+dcH9Zq/XabCbeHJ8Vhdj0GXzJVDBuEu27KNxnjBzFQP13VJ2VN+muh6SNGhG
0aM4A8QtLe3Em+GcG5eCQKrUWoBaMrV3L8+sCYjJdAQC0DiX3cuo3hNZhX19/8fnVW9rayAi1sfC
x49oRnZFKDM5qb8GrEG8JVe+CFus5OaCvhwbKMrb+T43t5FGp4DjetuF2cTg4hhYEYKP5R7S3hNc
9lVdb+pL6sIxLYP86CYC6ZjnKiEFz5xTQrGGEjo2h6HGSKaM9IJcdozNjHDlb7e+9eOU3Y7JNxdT
apRy6iZ+JNbA4iQojDWU58+Im25I7lhy0RlCh+zVxdf0Qjo4qcLTHQeyxET9AexlbyeYBXeWN3Z+
QXVAUGUagL4zZ1yp2dBmvgJhhhpjxdJ+h1Pigko9yBDRpXnZMna1rmVMXohnqsjzNEgBlVleEuta
BUkK4jLmKEltnVWAm/9Tj2hSBV7uweB+6OccFOQMXMT4kSXA6BoYt4TU34Xhx0bPMaWSWBH1FNlR
lrlaLHwYxf3oZDreNHU0uu7JXIhgChRuHwrn/RSxM/RPOtfLFvg/P3CAVx//zCMRcaDxLOviqEEN
AiayOdYtRsbcuZxhxoDs/ocJa+Bv7xUrFibOLOtyrhvXxFxC0unCRsSS5lyQ43yOJYtsL5QWtK4f
EXViGsgrpWVnY1bihqcLldY01IJiCbhNLnW4U8MC/Li4Waeqz2FjDbOtUA9fREpvGzrKhYEuUIKU
08BahRH9f05q1JEhjiCyB028WXP97rbJa2gVv9eneokNtgOrOZ1RdTL5bawHwP28e/g7iqP/wcBx
JdVKrLN8K9Wl2bSUO6GNzj0Wi4vDGoOI8J4Kggo7axQaWhmdrVilDcqcBhonDzIkiJKA/Ep1bF9H
KlO5HIMS7fUT6hcdOfqknwyVgHWBPtsNFZEUN15E/a0g5Xon0T/YrpIeDtIPN1fU+wmf2OPcippB
4ZPGFSfltdZPVNvBVyj5PhQ+S3DPuLFaVt0LeV6663fFwZr7DVpgpA/s0lnK/bdGkq/VJdlj8F02
Rtwzk0+KoUUDMzw5qTkQwwkGz+GBxmW7voX22uUkkrr56zgKkidKsCH3on0sx5wE1mvKkwwL8DOw
vKl0Yhy04edsWKE/hxVstqf0WblV8dqeqLwMuktDNtk6y11usjSPhzsbNciXB9Qz+hBtxCu/waaQ
M8ew8v44tjKQCSHM30I6ClgJWido8DVn9u54JifEFUonLKr3CYkh79sx5vgsZNlWcKakl3b/Hm2/
UtujidwLJmXgH/TwYhoZmWRGhaO3bofDufjIIfY4n6mECcWlO5m1ZbNyQEahXYrwOdOt+ZgAUT3X
m6jSlFHi78onIFTdscUlooyD0RcNj5rBkFZhp8gp7hYuwv5c2ZztvYlqRx9UZPhQV0THWT2VkxtV
dHe9CzDBKehBi97OuTRH5gTpnHuK0LLrOnFF+JqCYPywoB6O9/zrzbk9Xw431dsdi7mpNZULMQco
MEXZpkZIrRPwFBaLQ2RNrbak9usFmUNmMtkiBwJYkaWwtkI3AVJViaVOY/n1p4DQZ19jWSS3Hp2R
45z6TR/FjS66VGA25GYZNveO9ujNLnN+BjDK2hTDxQt3dHgD6wrZxrqIGshDvIi+AgRPbcnxzmIm
C2EdtxOMYZ/iXMTbnOwFp00BO19/Zo11lAuAag+zASbYOXJFWwEANwTfSauQ8N0+UxZpATqJbxn4
rYRsanjjI2a1Adgbh7gd44nh2wv9gx4xytl5XrvUJNNOaY5DSp+96ul22vHSdY7mOjND5G62occU
k0N1P4pPOFtQBXx5++LG+jVxCuoHXsxYONYwDBrADSgLjdLjGLl89ShAd3etEHa1vk/m2JY80pdZ
8GA/xOPouX8Q/7b+CfkMLTlRBM3mf/Oh91zs7V9SY4bhZp6tuT9kAHqbBwWNw52DZ82tL3qGjm85
zE5wPs57dUNGliZykdG/3p1o74UsHpYtYngEErekg3ESZyRzz79ddrNqCZVdJU5ieX8QcSrF/kMs
UxECW5vR/euHsr40Fhn1OiGx0wah+CrLE22NQjWXj3SrpL3vqwhFGKJC473vcrycTgQL5h2z7b0C
I0pcrJgNh9rx8H9i21mW7l4ied5lexaPnVp1PwYiRaXehjZG5mhrKPBpIByl/FgYheMStLzCM1o7
doqf7WcJ5/i3606X3jLork5H4wnOn86ZGKLUYWq7nN0AMr/KdZ8RkAfOqkUthWpuxS8YrysaCiHa
+Hzqkz6QdR1JdahkjhfJrwT+S7EZOV+4M41uf2JvtUoyz4NyDqNFrcpGwFN4tu8ai1A1Mz2/6oLP
emBS7CFHJpRQhd0ReYw+9MNFSphK4H478gvu+oo1rxNqVcV2IZC0+xaamHmKElOW70sEI+Zkph89
P3I86M5KqBQyJqkgifgNBDMaDrc3VAN/ZoZK4gHh1CGCDBKi3k+8PlKIFJeuJ97Fp4cmF3izJLc/
duc4ychyEM/HXi2i8n2vJGeNsNqQvf3F+IOT4i8/O8ul5XAD6VTpa00mUCom7dtWbGofzgrCUIU4
lz5RbbRL5aYUcUKSewmKHVZBEEjBO68liLGZxMrr6nG8RABGHmfedeMOmS4rc4OIxtefW7sGlQZu
0ciIyePEGT5iTxR/pW6e/LntdaPpwv7Rm97M+L5G/o3f7PbK8eiZ1478beBYwbgK75Sx6cmw9vWo
XHLRdDkRPjnaBRu+40plGzbQoyNJpiQM2VGnTJmSibPnqMWyLRKYf0zBpftm5dPyUVBUAjJeHrIb
JpDh2RdcCVRvbVi2E8gfwd61E5fzrqok41HIoGsD7nQS7MYSr70N8jJMB6dFOdRbGZuqg38aBQa/
mpwjyLKFsmnTQEbNG86SwcnkajpUg1UKXQx0DXcAN7k4rJWAKC/CT1wax+hDokVQOUcPdxt7SHqj
3LeMNj/3n+7LZMS127Hy7T32uM4McMDo88BOJtdQ8KLMTTSSkuvf/AvO2zCttcdIJjIAJ9tYgUCk
Yxxr2NvPn2vmC9Oufl4zCwaHdk11dh4u9CkZX0MsiwCOhd49ko54uNS9BGwozQlZG0Eo3bXTRN8v
lU2pC1wEsl//AFZOqxHoI6t+Xt4yEUCcuFSOUv6EejogPRedHQYsdcEFQdonuZ14zbYwZXPIH2Y3
pX06f+6TAn+0A0zPrdPnt18yFsJwkRfNUVgcCnuelZK1VAdu/lNNf20oWImAlYzuJHDSeXbMZv1H
1K0Ypk7PtxYxKU6LYD0kylTYc+DJhBkVkjpBI1rFXmglDA3OLFKjR8ymyp5Zz91wawqjK/pofNQi
oh2R3ZP+MCDamHVu9TD5BgY6k/Z2xmmq4f2buuDzEShOD0bBYUiTm5aMJEmYMzkCAgH/G80gJGKG
JIAoin+oNx8NtB1muxAIhf7hIrMnWAI/cDmoSYnRCj3KUw3UYDgMCCqcmfPCI7rRy/RJqr727ION
+VcXKSq7KiQi0vEWhnsm/32carg660IvV3vlJ71BXlIQqR7eYpy+1Xhnt25XTdcLDgVi3Spqe/nn
pN8FiNnlxryQrBqGERPZ4kQTnqG7S8Gl1NlS4RahhnOfccZz6/bKTv8YjM5CnsjRbNRJebfJe05W
qYUFm5OSMGW/cfqWI7e/oc7W872sYEGAmpgPZRof+jgcNfFA/DUfEMicnk4ISlczolYn1C9PkNLx
Ukf56c+5fxoyt0pqHVeWTo7MhdDsTm+FZEktyKJbshMvVa33y7tvdaapc0k8lCKbqxmM8fApha0i
kV25Us1H9kjBu6Y/wSpA+EiuhXpGnqCkdLZAJw3WfWgHBLQcKmDNXSS6USaJBddVUxJPXMqYTmmh
VVaupPVvHhKDHKOT6wjxvto07qDjXuLQV+pgOwENPNs/lxTl2ca+KJX14Lj0H1+jNoMnYVMN4IiX
smPBjVExjca2mKOw5y/A5ysoPgxAz8Uz+y30iHxb4MByOZMoJtPFRD5u6uy1e7cLAofT9ZInebuz
fH4V3wUOOmyds1QdOHogyRPf28ZEAwGnJ8tRagVidMcJErIic4yHMUKeVEOr276VQ1mRVHTRQLxQ
dCPQXkzT2XgJvUcgG2R6fHOv5CBhOmSfRZAA2U9Z/ASjsXobKwwwXoM/t6dEv0lh15LKgCClSITS
YH8qxOZ5py3o3/7wYAdFiwloInCl3197caRsjcAriMI5UmiPuXF7fRvABblIPKA+rkD1vTOcyjq7
HQkbY1NTe4DSuX7ux2kUb1F1mN01lOG47o9PiQU8vVM6TwrYbpOexU/NCyw+0iq0CaueuxDgRrO+
thY+bscMtLSr5f7FBTX6eG8FTZPFEle2rxpl+3ym2WGd5Z2E6wKxD3RliZYJ3l2OU63E9vgChhZH
qE2iOUr7XPba6IIty5kraQQGzeBO5x0naf9LUjK39XIIJ2MF6TSeneHDGPrk98UzYZqKic+5ueC1
6CuM29GWlK6Kv1gp6rN0FxRi2RYvYvQPbkJOYxvAAaF1UoOJjnHco1dtzE2Zfz+Z8dKD34c37X5T
AjbKjyZkFapO3pzlFnJ5atRtaosI1EE3AQPcfF97fm3SdT6OtBD4nWJLgNYdxEzyu5deLcxi7DPx
1CalPzo79xe67Kn6Y2sRr24O1KvZEhYzd6yiLn/kCoZZqeqpb+dckNfUXu/blCRd41GipLm60zTV
WX5lCX3fhfSTMmENeZUls0bhB0YGLwROU3IG31mblUcGv1yHB+SWHxbDUZDgUwqoDwWQ8f0ku+ZA
Loii7OKCFqUHE7f7LTeEa+QN5Hc1J3yItgew8pVHbAFiks0OzmEgkAK3LKGHctN4ozn6Fvh3B/Rt
bgygXkkgX9yi+gcHfxe8lRuXgk1UYeX/AQ44tB0ohR+Zuc7OCMh2NDeyULrZb5CZKkr/5o+7grYp
WLIjt3Iui2VGOuFPAeXSwovck7M/K+ZlCfUBO5fJWRKxJ+8TAaMspfiDJwcLIBeJdya7mhYu8dsQ
b+/OgNtALZ9PJmJy0p/TF+J3uJkqXP0tcz1JU/vBYaPXrjWLw8BOlPvrxXkDapFTXIstjEf0Qwde
wZjOMvhg1mcfrXCuH9Hxu4btAgfUrsi2JhiCg7sqsJD3nB06+mz3C1foPdvhTtOmEn5d8fFixcPg
/u8zUO/l4qTILN+P/XvpGFJaoB2Eo2QD9up/mH/Doea4g9VLs4IWOcn3xM5wioejkos4LGlfkCG5
eG0nsLG8NAiPvZk/REoJ72sokHTn/qYqyf2XJd5it4X4pqFpuYsmlNu+Xi/5jhn7uxdw6ogjAc37
P+ewbVd1+yMh9W3VRFhwpUjMEylfveyQmwllTvLaC9zwy1ey6dXRPXDY6otmlRl/yZLmRW1qKFsm
9NXm6MWGaEdBwBHE+SIF6LiXcmvEJg2Qlr3uDMuvRVvaDHnvZ4KhChiw8q2ADUszMwYISmXx/3KP
XGOpUkosVpJ6u4isyD7GWfXEoaGfo70WQ/IqbPeugnW3a9PdFB6GfuVzORoEEwmnjGJlSxnHxuWC
PoRzXRB18LusJ3V+6hrOHhRWq2wZs9wCO6C/fxT5MltKC0llGiGrEWsXZ72QuPUJqIbQxBhxay1m
STlg8WUyVsYen98AePd0FPAMWOf9dmttct6JHhywDHTQJcrAFjI/GMxs/+1+FSMtTaCBq+QFtVXK
/0KKboXc1qrIMKfcLHxbIBoPf67CeiCbDNrKDjFA8TIp8OPL+hrsM2rlBpOVYkYtrtzr1QkI14Hy
4zowageYsDykGRfguWbWKXqDfAblQSJK34wM2fzKXdgHuzs3O0MlglNKZnru7C1J3cYa5200wVez
PAz0nk0jkhkd1ui/J6Obzu56ftHsdoItMOITOzCZMrweCl0WlfWJkG2fHBg/v+h77Dzu2NL3KZT5
SI3M4btjQKa3Ni7EWAMdzevAMna2rdERsQafPkmWzITWZeb9bBYZ4mOpvKqiY+3q5Z8GkFZfAHzm
EmDBXUsWN2LPHMCrWf029YJFuSjPLHJEfKpJuTN0gJka6y+P2k5miX4xNb+egOnC+RXIcIILIYlR
PQO+Oj53dVB0MMRB6TCOzfgrDQ8dTY2wcUKFOe9YCZ3p/8Sa8aNTYxD74Hu6bycBNcSL8Wulbz4W
VdE/EauIbjqi6gHhK8IA9rtqw535LcNT4hkP1QT3zZcJ7G/Q0P8tMXgy++jSaas6SU3X5b/g/rCv
lg2ZlxpRqQtrkGKLzoaUi43AGpfvGXykvIZCbXSyV+6GXgKtEKIAis/woq+0no0UoBn3lh7K3GAN
TlOoypT+QVNPlb2IaoLPcdgGjPZwPT0riZYfCpD0H7Xm19lwrhVmf3cTG+ULsK4i66Zbr0/zdhaW
UtmskHOOp5IXzsbWcE0exMM56ihPn2TgESM50a8TPt3joHiGvuSzdk31UiFgCWPcwv2Roxi3wTyV
o4bA+emCVnc5EeE5mrGJk+8MMZRpa8f+NN2rcKz8nSvQuIlfiK6YrTJznnls6oiIJmXFYd5YbXB+
7KElrXCRJ5cdDkSZa2IEBuHGSzHvC02G4qZIOXA8wZRl9Bikoo2QlV6TGXF8W2qWCvwPetI7FcVm
VoKaJqVk0XCWwymRNMgHxV7dU0hIDEQL2LCNzQVxFhFEslUBFU4wh4iDtgPTsg+BdtwzTCy5LH/O
1eYuBBtrB4rD5OMY5VrCTAI2ZlRGG6KWNChS4G3B2QCYbPnitpiuYb5rXrjcSVIO97bwy7YcLBhM
w56+y9ADly+EBWzrRgRW1zOfWp0NcHsDg9x4kR0uFEBMeowH6jBwsQlNji+/xuEbyiiStrts3Qrl
bK4qzT2QXxD6yorV08zi/lBGMXovSPxuLTq4Va3Ho1ToiLzb/n0x8Ywd+J4lXMBM6w01+kXIOf43
vQW/ILxUwG7GBvpX0HBE5QFHDH8oXMFkWNOTpoFc1cufzU4NpDlhjMt9+l9KRRAhUW23mOSPD51M
iIeuGzLqhrCNS/rcCGxMjioizFn/W0nJPvn9L+cqIqe84KE9D5EUMXGlh2LCqW3VMtXl8r4hGyDA
DtMQKAjng4KQcqtKm1UefShb9aomCaqe3DrEvIYH1NRiY/wiwE/WZ2Ik7qLJLk/EGHVSMcwEGOIk
x9jZlM3wXearQKb2cMWZCAVmrjIoHgkHTJYL3fGmwDSly1PGxDGBroWDLt81R1H5PDkfwFP1/X0V
J++AM9QTbpi5qaHYlPTuV+KsP79kJ70m26dXcy2eKEdYWXfrWtXqTN8hRmiL/qpXd8xYuk7hQZbn
ITwc44gJPN7O8HF3CFsY0s7RDqTjqDZ/k4wCzDOC1FkqhrCP3Pce1AHtclAtxaOJfmsvQsZPV46y
P/19wWLjoD7/AXIOpfpd1yCRdR+OAPypVc6nHLdkN9/vgwq5rjTwwYMybkhR9bKT5fLZc1+MaTmh
2grPL7UEHCSrgIBoANCGZuaJGJMsVVyzFWQ/aLvEf3amu/wbV0XHnc36isO5YIGCuHXgMYxGKlsY
p3Sy3jIF75dgWr6cNmZGnXV6ieoeg/7o6Aq/ujHLzMWeVL6aYmbTzq+IECGYXlyxi9A3GY3LtaMR
nuFypxdwieah+6n7HyOMa1Gc/bojq4JGQ42X/ja5D/eikyKH6XitB5uRa6sOGbsZ3nfHzaws8XzN
Ro1sGEOAiU07ztmsNANaSOGSzarvAupKbbx7iKAp+1uzYqEUiOiLWtzKUFGhoOkGbpBVyMs8xpbt
Owkw1/q/5q0HlC0VNXxKVmSebRJ85BM2l/H2wFTwFvSsEuFeN3siU+DUo2wrUizuoj/1JDCmjEdv
rfL01p4oWdcqyxJWVJfC9waqikDzcK9s8S3tlJKB9JLo9PLYY5JYiEID6rZObDP6vn419rJrU1Zp
XCVk5qYzFcXAl3woLcgWqSgJWq1sGpCG4lAUP/DuouhfaBYmo17V8ie0kveZmGQSlr5l/J5bW5QO
QuNt6ROBFE/kefz84iaMxHG569+mJZK46Hf0bWQw05ckpYJKpMNfl3QlLi3iBBSJgcFxLSKJRF+a
gYxweU1NOnhSo+InfYyIoxkvG4MC/qLLaRtlJ1Gauvq9Pwch8uN2TFqh5S1LATRIMDXqe2BXQjZ9
VINd27c8qcqwl/I+hkWPwx5zVKYOR/rQ5SynmZ0eXlny0mGBySgxaeZuz5eSVScx3hYtz7CyW1Qb
KOx188yiSJaDYKbIbgM10HiUB/kmUXl6ozVhy7ICyRuFQH3vbbNmuclo/ELeMTqaC756Vu9vIOLH
8U4o+npQFRuziQFRfSIi13C3Jfesnsl+6tDJwjFikyDj6VRMTrea6j4ok45xzurfgYCzd+BH3Qrn
9rgnYGg6gw80zUX0WSHdp7mTf0kwQA1bANuQ8VCRiTEDzVW5AX4Neamw/JMziO5pgJA0sZFJmvAu
xXjDuYuwGGIgSOPSC898UiLOix//xT+fZQfHa8Cj136NxfWoyQIAXcmEM2c6qfiDhCbfAWFp6tzz
pYTKapEJgbq86dhij2ggvmcdWwa+uO9xECSdsKh7R4BK3Gcws3ieyvNozTl+C4uroSdAOdkSLK9j
6AWjnnyOExlx5py5GJ2FynY29/R9ngkV0rdzOPFrIx6clWspRvoyuHD/35JXvR22LmHhqFMILQ/q
3NMu4VmHJUTijlHofwxPXFAS2mejoOnQDd4uK85B78xLdkDm7yAX3xX4PL731R0I+UqVhJOonX8l
sm3wj8HfX9IgINKKuxDUNjbHxz8PM5AECNKm698U5CAZAv/DNKBwEvVbmmc+pkJ948/NqlzTywnK
uyXtmVxD0Y9fROVfgvCsO0kX6r+hdZPr6VFHyxLr1URDJtMgzkEGRyflJhNr6GBdXDGCVNCixBQE
e88P3mszCWH1m/OaFWcCZ2/TYhFjdmc9d282nk+mJvgOgTi8NCBc0UN/IaJV4oYwPpLjgVk1jODh
bWhxoF9EZNNUACVuyu7AXeSN3SkLBnYqLRRw3xIGstAP176+3Dh88yjoBBEdIJ5PhP9Nshd2Suwf
6sZSuz0VRQjpjesDeTfQ6zGUeoZ6C6mNmt8LJux+EAQvrEaTqstSZ7gI1aU6tOQt7t1bN8iB0xu7
UqFn5ZGjI/IGyyL1VrwSd/pPRfv44rpAELxQfFcMgoGF4mEi0NbaLAIRUX9ewzoWCc/lIzl0soCD
wyc6ZvbZdEffzp/EqztuOeS8jutjCgENONAlBnc1mI1u9UiF+uuKHtBg+PBI1kuIgosfoPe0l6y+
bC3/+uAH0jBT7w4KqrJno547zWjF9OU0A/jVxWcxy00fB0oiMhZPlugSPgtY61B0I48OhiqrhLCF
WoEhRNzIR7THRpOlnUB7rlEBCIgQCji8KpBpldpOKPoKAf7V6AyVYYe7DxJ8G6Ph/cVGvosXknWq
MBM7mfAoQf4pHJfQjv7OHJsUiksR5RjsZ7qEx5mr66IW/++C25vslS5Wme+vanh52Fk6dW4FYx80
nkSYy7SAsc1RgFcDWApY/aBhvxHp46dxPZHT+vrJzin7PDqxUUGZMX+4pm0Qt8i9YY+5Ro2fU+/3
Kuj2GdTtlNhHH3/YJHA5AlXzivraq7DW8xpCqF0QZTJNaeJgelArA4mQAhk3wBGtLId+35BGrQH2
jB7EckuAcx13TrhpL0WGYb3yFfV0mD31475dieNDAdUaItZwmdeLAtSZLpVSGBpGoTfx4SHYYzPJ
s38cLS3ZMa5sl4IVi0lHSyJLiYYdRaaxbFnlpQ8gvzH6k5g53XPoMxsCVikgKC52yuE2CmgggbN8
rH0J7C3PMeYyqaHOdbMgLc5i6c1YHNJUxpK92hKRS3rb9/MKR9twEuv9SbKCJueOdeRyO46iZOyA
wx80Rhg3cQbM3jvlo5RPwGiqq4t9Q4iL8YQlQEyk7MuHSBvAcjMUPXc9duP5Ry6xI9XkgzZmOUrX
HsiEzZJeVkWCf9agEBGPKHjQmpSMeShdSChOH/7k/p02viSvONp3z95KA995V0kh7CurPVy3W3wZ
R9A0JBTBEGM3nXRRODwbcQvx5peTfntfePAoXle7aO6iWSFe8/Jjj0V9HyoyCnQ5e3g7bIchRYU2
tXdif3n1G+1vLKOV+QxZmKVBV/zvs34wVOx9g/Mxq0FWgEKcUgPGH1dCGUuCy21GunCAonTIE7vh
1fTkhb5/sdxlZk2Rvg0GLtG3COzrnWoky+8ErSAm70LE5kkybRln2saFGuYVewGvlae7F2S6djRb
dcnKTXG2og2jxM7PcN1ieugYYbkrsmrBoO+RirSpIKWG7oYOs71Um4A+KoUNlO0Krr6Gx2riaOJV
cgCMjawlwZWs3WpVIOR92sc7CTQFofgLEwQExRgl2mo8LE1tcgmp82J5J8f66qYHM7h7li8xRwG7
EEr8Z56qZcJ7j6SQV2VJts32AsRzRVTBUDj4kTR/ckOzwCFKuI4d83ZEM+uBIXbUpwYl33T0oJUJ
6y4HgYZ9eKU9AF3P0nRkH1PVpycwpLNmY/0xMOAK4kWjXc6qK/sogQCyhiQxXJhcFmpmsIB9KgA0
pZ6jLhdBUVR+l4MOPcojDOfBjVVdPRcxTabFM6U8IQj+ugxWDH2QdujMxTOvKIko4VzA6342URk/
I3TKeCI1vtAn/jNpL/vxYqjdyiXK1k8Kq+I7hhU0+xp8L3nv7BklzbQk088KKeicz0VUQbKhxiNp
LqjTTiy9G79Ehi9GY3GlGZ+0HFmml5MlU724u80LR5M2ppj3AuPucw6D5iNqwmBWsnHrDt74kUD8
uLmEWLIHAgMHPtsVMaPRcCjFgEISkfr3KHqUDVxleaN+z+ZOj+eSpL8EOCzmIb+OYZE+ZBZ4WDJV
ftMO3yrMIEwFqh38+fnun5Od2bzSK83NjSvY1DnrgvJ2Y4YFedku8powYCWjtRK5j9LWxGqepvdp
q99RTcYkK1vrqbmsyPbz0q36JnqWAvp0nx4vnnGpB5CZMlALXXAfe/S6J8mR0rVGZwLdbMyUGNSa
eDUyMDgQfoXTNUicB1YVSxCNwRHVdmdiQ9QgNWacLSHGLuYmjKxqn0PlCX4+GIq4yaswD2k8VsAz
j52h0nPGWvT/OX+Iic8MC6RBLnrwGaEqcApMk2B+elJAlED9uC7Xke7j69A3F9i7/TKDYb+DBbDP
+u8oE3IJRSzTHfM+r1DNaWt1aYeIw7CsoJ/e4EApWvagR7rNwoW7n/O6n8VI/udXqC/BVYzYKZzE
c4LfQrayHtlkPBMOvpwPLqFipOV0P+ERYIeOjmKEDSAyzBSUm3e+BO48A3BOmW6qRp2OBxeM76i4
tAeGOoYw3dUZZEa6YcTWPzMqryR/v0kOw4e7qImw4NAEgDiIvgdoQCWZfRUyRyfZe/afDsg+GXWB
aymtNng/K438TavuGQRhHmnROAmwKgpLUEYlEo/Kp7sU88QGRWg2+RutgI27l8QP5Cb3AKMUs9oq
D/ZazROcTY+ckM7hJARF5NXx+UzGXQNwwgB0zCDl6U9AMWzydfheaBkx/y9ZcTocC7pvgjQ5hxJ2
9Youg74MWI2e+58mTi8pqD5Qd4OrzDno3PswSv2LMuCP0ITQtSFu/iwQVfnzguxOvxSef1JSiO63
FpszIL6GLk4/fU9Y4gcT7dUYLa6OC11Q+tD59nJrjbT7g7L8lv3xUzAf/xy60XuW0vv//90fa+M4
Df5G1hy3maZqkXRobWhgXVPdWhoiEW09IID6P94Kpp9fxiGB8KI62oTPEJ8bky8mdDBytpq6xE81
6TSuxpZR2uES1QEkPxJSnYuSAeMSHXXG3kWuuM8r6ajTkjZbNAW0H5KuigtxfHAb+GKQ0Bz2voeP
kMAact8RQbNFkVxG2f65zSiyx7l6CMGDmJVuqx1Y/x31NChK1XRik+VuqWVr7ERZBD0DMnJsd9xv
sRpLkxcTxaAm1WTlLaWb7jKuYk908WzVfWc4TaXCnQNJkCno6AC+nDYfSQ1tQRIZ9HnngRe8WSjv
x0Hd4QXi1HyGD5QMoJIpYurUGYg34KOSgECv2okymzPB7GvpsKI52v0xs4b6jFHfUwHg6HS2d77E
mkE6vWgeQAnvMbkvtlTI8WveZKgzX6y8aNE9n3oKkx0fGlQ8hj85ioXQRtqx3n9p2AK40gyEUpRL
+FwnpcmPju2bByRq3PhxyujedkuuI0nnOJ3DNm8Q8LmjsFOeMYSw6HC3GbRvGQslXIN/aokTLXc6
k4IsCxOgbwYGZ8eboonS4QS7hQvdqQs3QMCE6DzdmHDkZ78Zl+o6qtZN210k4+e6Xx1+H5LBGRi1
ZxcQKWa0W8ues59PsOnnyRlGZE5wlu2RspvMUvEe2oo8eXQLvWc37PRYf+chu+afTp+3prxM4h6P
/K0/ZFMc3EX1RNFK+/sBpsogBh+wiqmR8FHgqUgRqVy1L7/8dJvDXrC9+BrRKuz1SbTiwnEDGOg8
Z+qBuiMmcNJ9PHwQy0YouykNx9g/ZdR08AwYhAUiK+OpYjNqjOXIG6BftT5M3nazg1PxnBNSOaP3
hwVD9ufKoTctYetRUQ1C8x1If3lp1AUPO1XH/1Kn7FAt6qBexRGNS75xPEAYfeVeJ12A4CMwaXWW
UQlPvZInDsrsrgfgF8WiyFIMorPRmWyZjpRsjT7O2y8oISu08pwuShI5rv1eJdSkVFqRVIUDqPF9
Ygb8PCwLumjErwh3FfMiVsU9TuNM3lcooPDmYaf1dhpp87aYkZEx7dZxtvb41KKvvcaqqFsbqYFo
W1VPzLxNUW9m7ZsMyibVy8Vz0t85BYapafYWV5SEaVWU3DdrqujVSnE94qEMmcy6OFE1vphnKXgy
gh4LjB1Z1PVPV7Kwb2n0W7Xmgbhy8FP/TkkEsGXn20Vll/eYHbK+JFAmbAWAGz8dLGFWpOZWy5qE
RprBGmqhcEPPePwWO6ABV8lYSVm/GIrIGrZ/Zd8AE0xBvoawaP0w4BmayOBfH3DifIUL2BeoVvEF
ihnmwgldkcEBaCwt0mtoi3G1pgJZ1fUBK+vSJpvnUA2W+Ammqi7hRxUEuH+civ+CdRQh+RFFs5jY
YLDhNJ9tHn9OUZr1ElQsY/v4V5fO0xrLtkRvTd9U4lhsBdqcxWOLRSG2/oL7inXkshq4JUX8FIq4
Th16CxdMvSMSnjKLPPtVeMrjOrB52bK0b0ZUKprZaFROAkTvVsbJLPWrAelSjGN3OQEeovgZc/Kv
Bxn1EVDUAS48mkrdlR8RBhGWRPpoBZPLfnDHi1ON6xYBTkCwlBAKYCc3R0xGdNXfJf6gCIC3Oa/i
KuF+/NEKNDS43gHr9l7bEfYCq2ZrMMyY/6LmupW5iylzAMyIRBkhvfCfXqqYo0xlj4xvNmr1HBet
XwKOoqGjLBakbIm7VHtpA4/7PMlUEszjyZpvfVp+3+Qle1YZGwououieoD0rKSK5uQ6zO1LoKDuh
Fh8kUI2Ts05qje47iej/s7iKAnDpQYpADZmcRgEnkaNuSW+aX8QKBuaSpHeGFzCvdGr9BCUISSg2
WGbJ+K9SCp43er0Qun5urN6xx0hRXD20N84pNxPqhmsmJ3/g3WJt2Fd4Uh7EUCYL3q5NKZwBzd1W
Usaby/3qEttYtwXSJbPmrdJc75pZIPQbbmv+uZGbEeA53PzwYrfeXYFKm1CKDToRRBv386uR7lnJ
PYMP5Q0DG4LnuyTDok6NYyM32UpCzb/RQTuHJsJA0OH1Ktblv9F5PAeFHFzhb8ETtBsPq/U6UtTx
TkNa2SrxWC5B3exJAwFbZXRhu0E2QGbATySJED2fsDAa4FmVVxI4h/We8wNK2YOlhrmC1lnUdC73
2fEqBFe8xYQIoZLePO9PA/sVjmV0RPqz4A1x6nLoB74ICeWYSbseF5UvvuwNdt5tCFOa+URWVpl5
trd5XjjruWQWQ11dlhDkj/Zg5RKB4d8h1QAbsbz/n+aR41MIhP3GLIck5teeyu70qc813a2oCm5q
btvfDchdMRu86Pjp6+6xqPLocQFx9kwJ9vNsuFl2dhuNGy+BxXO/hGvt6HAUk1lyTvH2SbCljKYQ
Dhw1IHZdiNtRzPUOhZ3CUmn5vRd62X6Xf00YjnlCoGWLHta3E0c957MygFs+wskPC1zoyNuNuV0K
wg2gaPhSSrkPyatIlgYoHVpz1D1nYrbCuK0XmD3L9zmVv4f+uTihvnH3ViDLXwFLU6itXpDeAjXv
TEXYFhO5oDNU4s+3JIxSnTQntnkuP47UWpPB1eeInLB52VViZvccFcYKTNSbsosZPw6MmyrMXrK6
guUftMezodumPTESpNu1wzfvhOAAyKqYFe4liJkpNB9rUWpJkAI7i+VSirskHckP/Il6T0wxBKOu
VhR8q/NXC7yeJVaIEDgqjvr43+G2gQPE1yDbO8VrjAahjhCyc6Krd6QF6OchvblGbCGDcRTAaJK2
LgdrX5TndbCRLrtL0k1c0qiwDGwrEBM8zZD5cT3i5by/VGVOGNa5jdG5fVjwR5KnrtJGTBf/LYVR
F0y5PeLdYQlzn7a7KL1hoLpZFMg1Df415Vi2HcCIum5cdf1fE/pLpa3s8MmfxUd0svEf9Os4nZtM
7K/6uKD1BuH3Rvg2801s++yt9HQOaSTngBFoxhyqTmb2JXxFXiO4VqOwrKmGnzTrPCi6ZwHaVh+a
2fEOUW8E+p8I3aMyNtfzZ4p8K8cdZ5OVHCfklXsa2PlAOjToxs9OSjmtaHEiaCVsvJW5hmyAS8zG
NKQt87scbkytlR3+Pwmh4vJ+a9GMYp9coPwwsuDlWgaOnUCWMa9fHMImvLLH295q0SlaPDf45Bdo
R1Jv+NxXIRWqR71lWEnAAPK0nMo3q7MwpS1REe/X0v8Qeh912KEJyuyK8tSLlGitvFvdDKsHV9hI
ysav2jTi4wdJEcc2xPnm2b/P2KLxbMGWqvYLPL5OCIXrwnJFDz/rkDFQNrHT/59dLDTSu2+JqPNs
NDAsLrLNzOxo45sclY/13AqRImSCN7Pn/BVrgCAkWNsAIE8YfPT5Ou1qeTOmNSNsykH5YQHD6+HN
p+GknVUvz1v42M7dpAMs4ZY5kV41hS4xkZCayzj+1WmLVy7FqLC6sAJQ6Mxt9LaA0TuuERoR1aJE
9catKZq2fGwfzaru+HGrS6RyqswWzsWyX5Ddn7o55QQCGLUQXA/b8eIGpuwew0jHFLN06OJxzNlV
TpJk88iEJ+E//LAiqkR8QH3nJfIAyo76ECPtHU0Op8SySqApAk38Blm7khAGFwFPPcfcoNX8wBaA
fW18AY2vznZ9LmhiuGdhTUYCwNXjrLr6PVR4wIXumJpaEe/toAjM/2XfUDfvtAuZKDmnJt2Glzjt
nvI59ffOgLuqx+BeusxhMZ85xQc6lNQXxEqFYNcWHxU6ZgCXpGe3sBkaM52JzoDjBESCAs2a6Sd1
pGksfO+JqS46NtAZ0EBsZRiJqgEIoz1eaPepDh3zNSr5/Z0t6Ureso7RWyVONPfNeHEFuHlgM36F
dqIVeKZoAZel1VcU1tV3Be3hUvkuBwTqZ4C2vhtrA2zXh69CJiP1y76jQw7nRroDqd9glWUViLEb
BrONVHN016vPOEkMaM6W4/egO8wVvsdioz9B6H4RWUXYXt7Y0cjZfHeaP1RrZSX/w3ZEnUo+F5J1
Gd0f6lheAA9ely/6j0H2B3fCCIMubXXpc7CE7o6ws7OqeQJ8WXtdK8Bl/nvvuwk75PJfChs8tqzc
+nz6uLqa+GjQ08Wnf58+nZi+NiHDKG6xbHxL1RVk1LT/nOps76KKb2ZBEblNXR6aFN0D/oEjWEEi
zWDTcZ9I5AvKCXHYinkkOqNUlFaPL/QPurdC0HkunfwG6kKoVNVYkifC23hmv5n+N9eJBWxJKG8D
gSujXbbh5Qz62TrmfXXGV186t7+2i1OWGO0PayRV8DnQrE+etYl7B2WKxxZ1ARdsv6tZhFc/KVJD
tt9dIBvEd3S1hfREKnI8FV2lmA+4qiEkWGQ/NnkP8Tcyy28CRSulNJxqJbWtc38i1lSRtiH67IaV
+gqSkY3sYgbXNsricFmHPucRsP42ZDth9re/cg/g+cC8lN7+iKJoNItVdas+HTezcxtS9j77vakk
RMJX1TMsPuzbVpS+Dcw22HeTq+gGj390WQSbZep/1hfguVq6m7aT/+L5/ZYux9B8PTQxui0kVJYD
ZDi77og3s+z5JIWJ5L/m0wiVsBlQomg0J/wpZEhu8U0UJWIFZ+kv9jAc7VQhSieGdPJz5LRSiq5w
JPRH4+YAVFzVZQAgiLZBNbuTFyz6bIi/E6qDLGsDGC7UCjwJT3OuzbMB8JlQg9HesNEt3igpstr5
995DPfIK23jApxtwho/88snq7Odbha/x2O+SxqCVWKMi9jK/1c2WsJueGpOXYTvVV6XJs8c0nQcK
Lfzhgd78lH1a9HA44PBzOKiQ6gswVF7tFrX6cCbzdj5eEKHqma20EsLDv1GMQiTzfne/3FOOma20
Gj44+fMryVk4+FJcCfKA2azO7cDEQH5+V2XzytK2LXPizL2nDfRQeOiDSXx7g3xPz0oteMGVAGeE
H8MiIpQM7Y0zGLcovgU7EftkyHPwBLQAGAvMw6AEC/GAzxB6gycPHmfKM3KczzyldQFp5rMQnFr0
dR80uPCJ1kyfHMA/bQS/s6/fOkdSp5PFYuUwHAB8CL7D9cGS1FQvg196RFt+jA0R+WYShrKH6OIR
nqK1QkIR4qc4JXP5Ybc2cVnpDqFC8QS4/BHvhNFtpyXimzT4LWmNSlI7LLG4Z1O6HpQssdyJlDuh
TZhj6PLxdcZNQs2CCrHoUhOuS11itejKBqOELAW83pLf2k/yn592ubR8sCOUCHGihc1tVR7A6TLH
5989ySek1xL5M3HXMH5OcgI+bavL+fliscy/rJBwUJqVIElfbcSCpvZcvKnuTHKTS7tEwf8QVz5j
CWVV2EngMz0JYn6+6gbuQI65jRM5gkWx84VNQnOCluxvJTJNLvKroOZj/sf5GDG7/EuyHWVos6SI
Z64H99/t4heuMEHaAdqBOgbGUL011Jx4hl9T3K6WjinLv8NWuopQ1r1XYKcZnVpn0Ge9cq89rZht
j8yOc6JIaZX1m4xMYxsB4iwOvDj+mtbcOwXJyg2m/HT++3n76Q5pZcC1uQ5n10hA5Cl9MtEr03gz
C2F7r4V+O/pAmFA+uwuWleVI5GxM/c2zD9rM6eLbUjhTxQA6FTxhBzim5B5iEXJkIKia//N5AxFv
8dfRwsrIO1QWPPa1MwM6DYG9xuRuI5+h+qoiRq8M7bmBhnuH1XU6N9SYJKOuziZ0okuTkaD+ACng
d5n6nKAyqruf8W294UXND+haaLes+4q/28jVp0rbD0Xki5wGv9OodOl0kTl51O7/O2R8VRc5EgfN
OoeR284Df9ktEmna3CGrWGy1nTH4k7vhxaI1n1R+xbEC57Y5DIQ1t1tVr4CJccD4AQdZgrz8W2RS
N14d3A3aBiZ1KLLUkMTW57AuwyZGEpCqcphr7MZ6ujzIez1xypfeGnwWe/+rAUycCsFKDoCe4l3G
Pak6OJhwZ+KQ2tOIGwBoY6lEhsyy7EEH4xyIrIdRItfh2Azj8+cCHGiU2ffKx3v3J7iaZce5OHFg
e/mkhuc0Ry9q9Zh2O5Z3hyjg73VFMNLJnitPw5AxWtZ/ZwHRGaUjOub+i1BE0jrkwNa1boEP/m7z
9t0TMOK3VTnuL+pV7LS0l79MB1TOMGrl6imbjtHQA8N7BU80YTgd4v3EdgvpH2Vx2WEnKc2/U9gy
SPdGwfLR+LYMA8E4C2O54i1zVn/0aV2j2TCQDC33hJanNp9/X9/4BYfUAItD5Ah+w9KkTYhDqVjs
5/zu9dNy/mjtY+D0CzW+FuOnXwnBe4Ie5GSiHAAlsAcm+KSqVRps1AndTdgIE3ZeU+vPixtSYBJh
RGUiQ2vHO3Qr3LP5Rbb8I7nIHWkg9vX+K9eMAOAQTOu+tVJDtlRc7THoeGXkmMqVtLELtW7xM/AQ
Abl9EW4Qq2D03IqUr8p9xZn71HmTuVXNtQVMrU3IQCG2cZsZ0MytHDBARiKNQiqmN3SHb25yIP5q
Lrm0FOAdMUS2b9DuUkukBAoiQ0wYNAeNx05lG9V3WvFNhAZHrxChPaiykuv2P7Ti7++gycA/awf6
XYOVM3pcvBNNHz6aUunXGRQwqGSv55OJl3HEYH4+NQMBPurkIPsVUNx29dooNwfdRxg8Mza375/U
STiC02mWgYMKCBvOD+Lgwz4ifP85l8VRGWHzoYt9wIMivbS+jVAD58Ou1P9BOmb3Vdw7CW4MFYJj
tbcP8DysFZMcuFUCHDeTblm2jirD+0KY+BTpWEC1lnDxmW39D/msuHXmF8fowtxM4aG/y0F9Cqj2
TXz3FW/q5mG3ULXu2VAxggHaXS4ICUa2KJhRe4Ca7IwBGDgvR3MF9QJLMxPAGbbMd7/7b4gAaZem
4OMHjQ3L4vhc0prWKNK23FIg299k2c8VpNh+anT3cshTvZgNObgdv0LEnHZ3hF/npCabWq+99KKE
rPtjxMSWo03eLolVVJ/ZH3dF4Re5R9BFw826R9aILxLXKw3KtU7tsfh6fRvFPPpDLo/bbswAv/Mn
Y8++hruY31ZPGHRna60j+yGoCqXVv18JnKAhNyX1j1cwq4ao6k6m5eDH46JqNYJrEz32XYOT9aw4
DyXU2S9rjx8LhE7Cwkb2RH1jtC48nTeNumSYewDA4QI/dj4RXeqdErQzEb5gXH1tAewx+C6HcOcz
xHS+6U/tk0JOEwIqD2trWGiLzS3yKdue6s/SexZ9V8Taw/J3EkADWsDBJzAMbrbX1OA/py3VdtNs
SSgZkamClzTv7W1j+Q25bQJmnoSSLAIhdc5wptBmmhJ0hO46zI1s/tJR5wSZCAQOTbND2IQ3hFBC
9BS4Qimtipp9e02o8IwaRE2Ha0mpoZ3aaEanVKdqT02d+MQt+DuOZ6SkM26iq9XptGhaXv/+uwpw
U6n8oYabMvHRPCuPZ+XxwmzMsy8AjqwM4NLQoMDH2oOotEuRrZEv0eP0hx6AjzghJ0umxXfvUmEn
CBPKtpyd9Ljxg7GSMxXoofkvkUF+pGIDojkY5dCkLsijrdh+BestWOwbpvEZ9Ct2k5b+Y/lHZf+y
mCZHr4dex+QVd9YBOfKxLWIbRykBnfROH2UthYD0/l2Yi8FZTqiJzMbqvIDk+vU422mIrI3eYxjx
NyhJNkYhRkW4h+muzBig7p8k2FDvXXdZFH6y7HBtjXo0eGVtoL9P/ZaYesV7sA/W4uztU7zCjfyV
Ta2wkI32ABB45r1bSIQoBVWfhA6d1/DZGdrOrnh4e27+TQ5ftUo8dyTUs/nY+3cgygy8CFBm2tt4
Ga8ekmrm6CuiuHnZ8tMtYiYQ/itwG506oUGTaWzKgVIiIptTyfuFZiNXMlABFP5RBDR0m/tw2FoF
bIyUP7ZgP3RkIYll4h72OfX8jrAGAEZ3/MVgpE4Qbnq9t6DOE5IPHD6QJ/myhRMa5k3JrgAv4VFu
QMr9V3Os8ypbRvnHVD+TXLl5hO/Xfw7Adk6kPzkiymn/rZDx15USUcyVug+TGu8NfN/yDFWodw8Q
wUOkhrtGy1bDo9nUclg84rcAvZ5DPVNo3zhFNzlm/ZBtaNKJaBCBMQQTYEqNtaM3wv2Qs7x4mioV
A6/p8eWt81eWkOTMsDumdLr2LlwWIHpyZ6hSacp/DlDC+n3dFVWv3g8iCzBJJOlZQ89Jt4Rr1GNt
M2fzDGIjYfKeiy7jpZTZbRpEcaq3RCn1qFNQO0r/4ZKVz7W/4EoH/xnOSNN3eqBK8KYgUlyaz/pB
Su9gRNddJ04VgLW5DlZc4yjEginnxW0ua8sAEDI0mW3nqtAgv5NmT/8mMJEkfQd7PyqlwcBj5tKk
pkxiHKdyREbcXvGCzvam157TE7VjUzhDSGzlqTKyQPIrXR77sMsrNhhnbNbIE8TQGtHWgzXhnTT6
SqQLpwBfn8pYB63tFD8UwGA6cFJLTulHj99P48TwUbQSCt4Oms6VDqMzvVQ4sVlFNTdFAMhh2AsW
Z+PXSFICWbYQ4jJH2xUWNEJZDsu5h0Y4miHBbPVYSLoI60lsglbhaL+ucLJ4W/IWT6rhQkznVPya
hkolL/2b/0ESaS21OGlNwF3pH2i/6+Qsx+3sEr+cMPLvnqSW37AyoCnTFTjlIy4Y2ClVaOyv6vO/
74neKW/u2oQ4VbQfZxGcIIyE63kNziuLUKsHUZQCr6P6Os/+Ze2Asobc3HJFaa3wwMvc9kGfd16B
GXgCHJXZr6KOff+r48mUGQeFv1nfIBP+a14Jqw6o0dGS0JcLsdWeo3rDGC1ZTipa7DCJHAlGWaj/
rgjM8BgjRxe8hSvTyxgZPXqKvt7ahc7Fga6gn3I2FXYOI7lcJyV5b3peCYuLPGgCDT6pYIablQmA
1WdySY6Qvfrsvd9MFZuSS8jpOL/Qzu07kd5mwOplgLeH6piceuRCkE1Y0ScN2HWGJLa4rM2mvaBp
u9u8rI8FH8tYSKZnCPru9mD6fjfZFhLOyjI52tB5f6cvnLbneJzpHAD1KBnkCzAUT77w1XSj2Ndf
5z/tEUFi+ScNSMtoDi45oY8aPHyarkflZcsN5iSNiTJgNrhQv/sqBPZbd0/t+f4fUhi9jUFG3rcG
565PoF7fHy8r35lngqgqo4VWfY2tuN6uc6TC3BJSOfn6wgq4af3aXnvYItzNdOGlQnsO/cj8kqHy
vaOIaq6kbpkMBr258XiO1ZkDsYCiTaV+iyMXueBt2XKQp6EIQH0v12zECLLzfp4ArOv24IkHN7Pl
1fRpDUA1r2h7wPxe++6GlLwgwMHMsJ58UtuyiHWu//Yg0kx9mpeqYaWuMZXnpRtrzKsCeHEbDPSo
U6PeXHBdgbVJs3Eafs/FOrpDkocpsE9jOmipWggc0a9tvp00uS77gbTR2w17b2fYWAeG/bo/rEWE
mq3CvHUlPCmtM215AvIUEOq5J2pb0JDFWkJJyo9LEApBFsZTN2jnTr4t57Mq2T2QyjeNOuO+aXkR
ot3T6FC9j3l8n9fRkhhwXwneNEY5LJzOvGI37RF12Hss6adsaNMAk+HTNVPoB+gfk+GN7ySBEVuX
Qqn92qT0p6NmosH5haxtZAv+vZAsRX1taWctUHIst+s+1Ipcfu4CLi55vGiZc00nMkQUMrEA/tV/
D14Hu2GdN5L19UqcDeiEHZLdKQkmnibxjN/kGLOzzIEEP9faxipX2+cO098ZNoeESrytglpaXD27
Cl6Xl9r+uTxtcrxAVIgXVTBsE27L422Hq3qTPUFMIyKQivSk9Y+0/Jja0H8OQXx0YHd62piF1rF+
Pt8K9nGpnnlsIsPCM1es59gNupB705U8mJB5JuUYE8Qnnmr4WLJ00UQGn00X3tkIFvMFOTsEtDlo
3RUzUh5T5JujWo9vQOU8EJYMPgPIuGU4l+a6o9JpAgP8ir2FleKtaKZaVBjUo1XdFI+DLk44NrH1
RowKT+JMMkUCAN4+H4OpZzjWzFgwVtcts/Yf3Zuac1e1xR8t6cpKB2A7IjJMc/5wmBGDSYu6xy8K
Fkq0Dm+T45NZ7aGZgYcDWN+L9o/WadSfV8reUZai6A5yFfOUp4CYTblx23+o8jzsz0k4lUC+9IVV
kvzJ0yd6w0S5y2GwE1FJ30yb1oXm+vqFy4QC1uQ10wkfz4yCG3xAI8SMFvakKBizjbdYxUhU1c+a
4WUrPJdHtaB6gxjwKSp/ej5ppwhgaj0IY+rOaIA7TguzJUOHIWhjgX4WwPPH0VDxIu0IgmOcwd8b
itg0rNiibv7Hh9yqvkg/tbqRnqJtE8uijSTTRfRi87wFwbH2SXDHWvU03vonn9iw52JG5QfVAPvD
W+5D6XBZ1xFwUlRA6o4m84j92nsvgqB8cFDt5/n0ZVnUtAp+eDg9sWCcQ4n6tuAzvdCDavlaTxgN
R32HkLcr2xNg4ole7XekuoyX1q/OPStPLYLSQOPxQnMhSg6F6VXhi5qyu7fpXMrqQC1bnmHZ71RK
Vl70Hg7m3KC+y05su+CZMDypetwjwMH88jA6487N/p2JGVScYRSh4MG9zxcZt5ulrJzSmSh6boef
OvOgSFuwADM/IqdrAXwD6DBj/h2aC3sRW2vtmJAzps0smdNDjHKeRFnfReYY23ZLluC2f5J28tH4
3XhUM3EPpljQxB6v9x1nkIKkdHwKKttXVJY4U87wRZOXZedli6Eb2Q+gye1nZzegRfP8+fvp4p2u
LhZ0mJMphWRdyPrIKXZXL1NQyvGEez3xplQxIl/56r6BPVIXJVcAVlMYb1ay0CMkmYFfWqnVXWFk
+2S3sDi51hGu+mITQiRlgmyzm/4CYPJjpNT71QC7LVv0h0EbwZCTniswyk2XjdVijDbNFDFEU7I6
vBUq72sQN1zEEB3/kNB5rkaJQGfxx940BXj3O248Gg96teMUwrCPFXLmTqNhprWO7dcybPX5vHRa
I9drvQGiBuQoNQ5awFWHW88epT95c42rq4mwmZmp/ClL6umJRVJF2MoVVy1fs/+0xEWUa49UYhoC
vLXE5PUzWlhYXCaIKCcriuFpg4JnByG30vTFGF+mVDTZm5CjBKvWr678/6Zr3lAYF4WShFHadxBR
+y4AtN1ma3HU0fW13pYtXVTyc/xQNYrH2QwpLUf1GEFI30Pb9IpajbYcgQBGBujgc4bBI73Ce9QX
PdQZH3lnctWycLRoYcRh/6kOq/enWUb3Jk+c4rjrbZqlEb+C2NJdAm3843v9++7lsYRaGe/54tqv
MicynLgYtU1pO7XQJmmOnXQ6LCEFmOOKnzsKLlxif++hFiSNVyQEscfZZ8j3lfRN2jY7l5zCrZ84
80wZp8ZEH5eF+yrFTdaurg1XspHUiCMfoWbpmH70fYvTJJ1gQebaaS1gXm+Zb0p6x9LUXAx7brdm
zIpg5L0v4FHBJgNXi3/zteXshEYj8yODbo1ZT3aZ0q2S489nd+xYhoxI5R3ERGvANYnCAdQCqROa
vL99e1zxRcMUkjHco9M1JPjK/IWfYld+BGk/geaajwNGb8pt3bI/fk3pbqLWWDVZRZQqIYcsxMkW
wnLZqPon34yy/ydDm8SdffKTyX6zT4Zm6l2TGy1cJYskAviO77wzlYF8GotZD18kBAlqFU4Dsfyq
BkeMlBDRdeIQ8PppTJoHuMgbl2XE28ofHp8wSjALg77oRNJjUuTnEFrUWvQihxYUWbYMOcm0kBHh
Tntn/thCjZSndOQf6CyztWl6RdRBiFJzr8acn051oyc/HnFfwtNnwl0NPH9Tt6hiOnlIm+qXlaet
76LvDZic2EtMAehKyhpU7hP5uiLaMFPVwc2j6h9Rj74ITyfS1UFylQp+3I6DmMXpT0QHw3ekZLby
07/eObfpY9DYRiZA4BYEmh9pmbjuAyF70EpCLWkF3sPco+N+HtRC8noNrCNG/fYGsK5GeReC8Q4R
SOWLdgaSRvT/QBysdMQqY0HtO6Ixz81pXx13qz/Iqy4PGkMumrpr4Y/NcK+VROW6ed04uZDHKm3Z
HjF3PyJekuRnrqLuzo0EgPfrUCWVOHjJVyOdA8myFWcpQBhaJcxI7BsW1hI/85lSvLF9DbwQ3xEm
znVARllcBCnxgK4nUIXl6Nzz1rmewo3ZsfBICT6mHEr0EEL0TF3yKb5dfpd1ulUIo7SWTwJy8wEk
F8kQlR4f5ZRzN4lI2gJ7FmA/qaYn6wk+Ur/hogHSwmLkqsvhAx8sRsOdP7ceFkjfRixF40/sIphS
tv8Kuk3LTb/Hi4BH9XDhkkrDM/VScR4cxjvS9bXHAanoqfvAmjizAkSRFgM98ISh86kh3pAWQnnI
HgRGPdOHnAPlHNamKa4jhVaZykNLOJmd7mA2LGR3o13oKlbWp1zKWlTADiz1ToIwHRmBjfXriwR/
jwU5jcmduEp4WI4IcqvGDBSUsyCL2496YaVl/xmzmuBqLQXcpnTFX8CLbKruCn902HTf/IiGWJI0
qm4S8gRNTZL0mYijj2OH40AbcY8IwoQYefHCf3yLZzDRPkqPZXa/rGyIy4TvzZTBj8bq4A8v70sM
3qZTS87K94fN8LheI3cs4n1p7wQrR5mxz6f0qXLcewkw6WITG2NWzS2lrYhgF37cpP8AWWn/sZBh
eejHdCRFK84IaUXdvrHQh1ajktVYzc27EMSDVW445t2YJc/YRSySWuWOGyq5hwUmYPwbiw2nEja6
Su3t7dJKBa9GbnloPMnJ6YIa4Z554x2nf3kJbnBkipM0y2mMfc483apYvXtTXIiOdT1EGp9jtcWQ
6NFWj9RYQIP52Rej5GhgDx5HLSHAN02Aa/cFVRli/LIxyP7j1iUqpm4apdBG/HT7PRZ6BH0ttlG0
7iv4kBGPbPUMIT0YHc2t7F6bmNuXwUlu8KTO+hI6/aEz9oFunDJDqKZ3oe4vC4A93mZAzpGI7yfF
f9KuIkcPL7xb2gNri7oTG3Xl3A2/1ob/Kncf19+8urWjuN/jtdriVkz9PRXsMSN8PTziAmzt4vse
/w4Y+0zzxJSvZXIL+c4/MSlIr6Ri+wg1bw7VXHO8hWVfPWI56a6pW1QsIq+HfYzsiwevaVfAI4AL
/MeGmRmr+8bkLOuLes7cJymtgDvX3mnto+WQRVrrUGhN3/JeLJ5/AZLtBc7h+Wl8MvVKtGEBUXjq
SLJisdmCfNyFciJauubr2TTVuXHpqAfSyJ2mpxWWMTQcGYYki7+lTEdb+SRGpMvV8kOD/C5sZOi/
kbmo4Y2TyclBLM9qEr834DKFt0vj4/yL05LiOdRYktA8p85Uoks2IcPmTxa4bfN0UUZUCl11xJ7r
SjQMdmHfu99mGjsCWvgoBNx3eo7j5OWnv5iizS1prmesUMvjRStvcBHhKF+DdOQdxmd5O2/UccDa
ICC8GQexN+d4ULz049ajGeKI1nHbggx4zgDRDSSvGmJR9/qduKojIL05w4oazOJ2yfRvpSM1Z9ew
hTM0qilv8wPkW1gVoow1lZ2iMeDdqAjhDRWW7dMgx7dAqj2U9t39CW47cO8wPGrZy/Alok9T9+92
Wt0N//QRyJhHhFnsGDqV9Exk9j3vZe1xOkI047GFOID6X7RcYDfUao/feOcEIgAUTqKxI/x3135U
x854FZjiyVo6pIS/X+0bp5xTOxvv7UIokIfw/+8egTBFzfK07JJpmrP1I6GHXH0sJc8PDy/wFe8f
UIdJEj+mr61yHCiU/GnbsMiOzYoupwwS6ovykPyBAecyXHjucupdW1Zxthvb1HJi851RAxyn2yib
wdIVjD39pgLte+f2CXFMYrYTzlvt6TtHmTstNKrFOz0TXsKX8qU7K3cMb+IdDY12wnhF94SOKI+a
B2tf/x9ufjvqr19HIo7Wp3wDo4UrqJ/tBeCEsqmO46GHOBYXRbdLoEkwEu5vx3rvFN0YTWn4Y/EB
8YtB2AxjOkbiBt7QgiCM2cw+0hNkHyvneHaSbmrvfStNL9rJ+ld0UWy2Lx7esazn9slnIAd9X7ag
5SPi0ZNk+gZcz4oUOavOdgmt1wsLiMpxxjI1VstSUIWP6oFTjTmMgLy2mf4mw0c4XSVa3DEEEquf
vFW7ioooZC/mRLoEJCuuBuo8FffoGI1+fpHgrfV/sBENDCHZklX/irKaJN3U2J0PNISAciHHT58A
CF/T82Y9JK1DaH7wbDGJen28LI2o1hGnsKZ4XppFcwBd1WUbgxJiv7tWyEfJHUlFBCcSvoFlH0R5
uEFzmK7elGE4l5o9I5YA+Oc729OGO4BE+OhxvAhFZWAozgNPHOHuWOCu1OR7EBSGTnjMKmptMlic
ZErzPcN9oiqkKLCHfmADQrnNMLN4k+2pmrHwxccloMuxjcCqfCuSEE5yrAtzMyZF9WDrGzdp+X0B
kFdFDn1TDwTzWgpMclagfi5TFIcbHdBJ06rLomWnx2RqllsK+IIeZlETeKDJE7rptCuYWgkFhO3A
PPENCQ0p3ysB7f7UTm19vkSSMLgmttIbGTNjb0DkA8TOAXyf9Fps+f9PnFs8K5ocyt8F7VVbCAj2
ZSH5zg3dscak4G7u7SVKRxgTIHnES6pIShZjs/Z02tdWLq8wUCUcyP91Rpt2qLSU6YKOtn2HJGDg
P3z8QIvQaw83ELYCUJmAVvUR6Kyinv8IQ0rQa0zPG7m76gtbu6sUGw5Ih5BIcT77jG7cB7BpcdXb
1NUt3+vgQFINAg0HOsnFIIuLEtOggdrdIIZTX6wWrWX6bOIwVPndroaAlKw/NIFqgH5Q2aFcLTr3
yR4IFopPLUcb8+Ltc/Uf4VfJM91Ltmm5hqWOMrZmoafC7yhe/iAuLArEZDBjoHfiYX9vF/ERc4+0
9nEswFoRXY1RyFgdMiRiulS5vBmZIDsPnqbqClixTULnpGYnoGj7JGkyY4EOXvvtPBRGxF308Ps6
FzV6uWKa2q7nzfbdJ3SJWxgVGhDOEgzRAmCeTqh0Yq12N+su5X3/SF9tK9K3uLs/PIvbhYk8zZMx
txfjUOoo9PRl14cTxsjw35A729ddF//Quz3ELkhKgCbXKwRVZUsoZmG34e37pLTFYm4t50oTDbcD
n3liVCrZVEnqNBqR7MHJyJ4O2SebkOajs/ilZYQIZEJyiId8G2V+QmLYuNTiVDrC/aQz3vNOd5js
m5UzfkXQjVdKpNwUDrBwvQsq5DcxlEJ5lKepCDHix7P5kFWI6pJRLHOgHArFaZKjk9CDhMhUWzHx
aLksydAuRO9GJPhKQtuuonXMLyV8Cfxb1U3I9hrBDG2zyhs0F8gAhO/nylMFok5kE0jcPVF+1y3p
5BVDjzlUdYnvGak+U197v03HnhF0Y9zWBj+yYoykbzWor4nUEsjW+ZPymsZ6yhO/M9gyhFQDcKew
2c9rbwQCOJnnK8KEgN8l+kVGvqeyde377HQ+LvL/8crvD1IuqQ5tYem3q17UkgF3Gl3JQHrd1aeT
YfshnflC9YcxH1+hcJKNHgp/yf/yDsp70XjIfOJ4pLdqBIOw1gOV5qMW4X12koUoY+F/RBBUItrk
o8m6NJY4TsYPz3K6dnnY5+osqAG+jxxtgrCsp1ybarNpxqa9c59ZiJQ7qfpWs9HjIpdmeRsQjkQu
KGewbgAZhEKz61lZOifeu7sUhCMLfuWAxmKQrTmLU2/JS4cL0kQrTK0buHTAoBCjoUzcMlOGxzW3
Vj5Uim/8x81FkTaGr8iudZ6wkGoPGHyB8SWqQ19j/Gg5oY6mfcLTV/yWdiIjko+7RgTtWmYh2iY+
wlOGzp8ebe2lJPKPATwKwmI0/3S9Ia7TIOuPo+KXvenxiG4ItmPfBIryWajlMLfLZW2689ojyzzm
9h3JqOlOnd9jxaSPpH9eKVFIIFFlI7jUfEtcsIi9q95A7o8SodAU74SfA3v0Pb+Hgt86poaIe7EE
5gbQMiUPLNtEwy2wf1ueTsg73RF8YXlJ544ITDc9cTTch6NipTmyfDtbB35khnl7UC+37i2C+3SI
C9eLW1/OBcvW/npaXrryx1cIdf0FjR61SsJWZEx43al71qqTQlRHTo3QzKGJNk479ONPBlt4EF44
ahus1HLoe2jX1Pt32UeqMJcfKo6ICZInQd7aiZIFpZ2kzVfARnMWH2VM8TGR3VUNQiXRg1/fEgLu
FZfs3Dl+sF2SbV0g9UUnv7Gs50rU02G49aPh6hg14mUZrRUbdK8g6B9TuHqfWNSaLvar3BsXgBya
NZpt5wQhhnOkGJOh5RQHQ21NN0OUGGQaEvjvkzdKEt7ekalMdyp+0F+eq7ma+zua2wLW/MUOoqz0
Y8V3elJtO5jniDvHGuMl/tMJB7c5a3mCGxmaLmeTCFgr8awfeVaUXy9W3rBPyGqqHErIVX8x0INC
ysmXrGvrCfHxBOKDvfrwXykpub+aacacZXeCsdosX3y3PlF7iAiQCk9ISngxmqqYPoWdvMP0LCml
oKz+kondqp/MA64tahqSgX17gjgtGCGj605AxAGftJGe4hs7gnXhKA/BO8jZf8v6+qH/sPJEaGL8
tG1MCfcZDhHsuxDtPH8KC5p02lFtImg/69y8+xcjU1xGZqMihnxh8zwn1UjTtWCoB5aX0DV+e5ZH
nNayPvl13IrTwWl3lctabJfDjMEIy6o7g3lUgJXn304Iaeb+TDZQcXTdCUz+EgecudDTuT89P3ko
SgzPL2Ag2rJc+nTf6rv7yM4CCvV4x2yVrED0ioid0XU4zYQBXJQ5jrXro7JxQFi4G0mbpuuaKHcF
IUGbH/hwSSQ+fObsiDNlc+x46+TQtRWZJWlWtlQDo2XnAUiOWw0QXz9hDqACeE/zeCuRe42sXWNu
ceWC51X820W9PRe0n+/2C56taoCFE4pG/Ic33I+9OI9Aysjar0WQDYawimX50h86Ce/HJuNXqBIT
7vvVMJZ6/JtufEGrXzG/FzoVH5lMtThd7DCXJ7fpywfvqoJDnN+vmHOeGfUgPveW7QzcNlssH2OS
LVkfgnrkd8N3vCNBlJwc5047B1EdO7zMEJTVgvB3tZmjjRaqJR0jJiBrQ+SxMOn9uaLQ+4LvPg2Y
7TpUZrMjKjcwKtXrAHsl+EJZbOivbIFY5rbVIbMdxbrsiQ4WstHBGc1rZt3yeOtE9/QhK+gLAb3K
nrUg8b6/oHSm5M2Px1JcWapHYIRQvowomdw18ynrZkhDSAjC8H+ER1X/1ErtKvVgTteFp+mkDQuN
N5PbpHQecXoICpZt0/sUdpnt7H4FWP0M7z78V9X7x5XEueZN7DlyW3IXosJdPxP64cRZ20mW1zLT
mN6xIa9XzpyKPAyzL2dpUaUZsUSH+7/TpHILFE7yetv0MqAKboGkatykrXy1nXFQgKXuu5s9op9e
6QZxAveNaC0qKDcPzRe2uEBuSforhmD/Smp2j8ZPDYD6ovy1ydQBniLWE5oaTJppsHBhfQ7yFX0R
1rljDp6XpFeGZcfGmcabJlmTzI+9Em948f9TmQn2wKo8ODbGEc/JWjsxU+XxoGdQ1j5L3a5clYKa
d1PbTTTZTZLUU0H0ZHj/PZ7nyfP/nj/GyP+ZFN77d+U6s1A9gZ8azxZyaZFT1d0N5wgw6KXQnf6U
ths+kWhidPwbKDF5xqhvVlAImiOo8oAH9Q28zkkmR0hx8J3P0wd9VYh7Y41z4Tg54sF+hCiEnGYz
4yvTsrcpuO4tYf2asyHMksDWSYVGuYH11HdLRKgMwFPP4oqSlAJ2QYb7pYM2bhNfvFkGFlmo5o+K
4I+AgtxWzo2zpmaP9BbAJKKpQLSPdr56zxYt98bJOX1PHp1MHBo9oZbu6UhKV36HKZTeoAVVVeSl
dUCGhNIxT4/MfToqFv8bVc7LTRX5+t/bYEkvQNrGN+a+toEktzDgUuF+ytxd8iBhUQS6ymLj3/zV
zLY3bAXNBk5coQJSvqX4huVwtsbXvI3eC+DsN7LkMguHLjZxlTTiELvLdWLOB/UbIbR8DZ4BEmGK
N4Kz5ewe/53w9yMyLFImZc8pWeDbK2yUlt90FOxi7TlPzYNyOQrpYX0JrR+FfFyKpNNFn6dqKiam
QUfdP6M2CyTKCg+ymFmV7Nc+c6YNO7y/yUZWpuCl1f1B1zm3SM85YylS94JLECG7I1ioIQgEeLBG
MjqX4pyd0T1JL/QJj08OjtJz18QZhsbZFGY6yzcr0AhHtaAJ8JCDmT+s3NVTfllx3f3DFLPfJXMN
SCAUXasnf4NR7mf4NaIHqVh+YpqctBZ892hmeatTCtkeWmXYvMfGeA+yKaWKtpdjiyrTpxCxgTEQ
0/YS90s5Y6LU0PHlmzL9Sz38K7FznYuqnU9izb/Tl0VAGM8C4y3bgrmImWD0rCNgOfTVj7Uigbdo
g+EWHUtHcfxZ61Pn3AB9lbwpnBn09BPSNZQiBaMkkqU4kVj6VduZhL7nyFmHK0Cjiz2XS++fz8MR
qglLs03vYPqSR4jxTUdLWhpijGBoVOQqBroSO0+ffvY28YD05PDTWeV3UmkY34E5zq7QDVczmckH
wVWTC1BPvoDyduXJzWkZvlV6zJD1+889YQ8HMTZg6ZSDUSQkA0b/LhgkXHPjjl9gPlM449daX9FO
RJEECvwW1WYd5KhLbHzW2irO9TtKZuj06ifvQ5inafjx2EKSycYTafjdiUE+eoukJ+QMSNGob+33
9FFm/DCWllwt4oHNVt+NYjKRKL4GnBybKh0QF7aJcundRpTHpt7tBQcyKwgYhxnUqpaO2nPUFJXk
keH0gAMJmoDn0717guPTn7b9FzH9ULfYl+DVtlQPMJl4oULk1nBMGH5QeYn/a04hYtMnmRlGgiGf
l5eOkXHnHizj5RJSNxmHnZM2Xv0zjIWQjdY9J49xlLKYb0WkLSy0TIbSztPgFZ3XDvnw6n3khvLn
Rmh6o74NcOa2qVerlZPyLv0jNqKsCtVejE35uzVch/4RHDCqT6UnFqH7EVfSsz9gX3TM71b5u1z8
YBQ2RA3M519Ex4i2U7prizhJk8QOsem8m/fRjyW6JH5q/f2Zo07SnRihu2QFkkcFfWRqTZHs26ZP
9Y1wxQbXPK99eq/6hh1iUSNGi9CRNSnQIFSq/LbNZBdNovtkrFmPFhE8SHIO5dPtauH8ux8A2TVO
I8iQsSOprNuwELKr+ftbBoZ6icSPENUFEEQKuA4OGfzCQOLulqT8P5QMsiZx43zCHK82Z2OkrWD7
F9lgcbYJzAQLh/l+KlLCVcGvmEWgw/QJfsbP1R9PPCZk7sAMbBP/d8+NPfw3VmPz0TLP7eHe3u5l
gbO48sV9Cc3X82HhjXoW0PvtoyxVv8geggj2RN4KrMUkhkToGuPs6CmB/o8osNeJNxgQTuX8tqht
Yp082DTIp4Mco/3HdwznhxFjsk/WhEnd+FPxOienEOkq5YVqsiJIJ7m6XQcWVC1yfvl0s9PJ00Ge
VCiG8O2NDxH2qB/Vw9CQoHxgs/Iep9XrtHSZogJlFUrms3NmlVo3+eXUl59Sk4sBzbgi0P/A6/gQ
iENWfOoyKqff/L5oh1PlCr0ZNasOHjqwOIW5z/x9JQhcjDN2M6NzJrSUJr7TAWC8j0bNd2OfDGjP
2apXNE/3o4dG074GP2Emmaq9Pjgp2IRrkBmVtW4HMlAbMaumCqFiqaGK5C8E2gH7gifp4e6t7w9N
uKTpglu4ES3rwTYsptu6H3Vxd5jVDZYSfemkJuSyI5j5SBooFpYgEK0lYFUbEnCMeudyJrB0M/Cg
xJtPCzB97Rlhz5alS4VhMM13rAY+OSYpg1emVJG+iJVGAqxWyfcJVagjVy0RhpaTSJgsSR4fTqKQ
zKsU7bChTxSU5WZjLwhWlbIFxwC6oG8fEefzVVPrWtJn8EnxGx4qHA27E89KFnxeaNkIPSKSWqm2
RRY/ePyseer7iv2q4BCcgC+9/JGzCxAekxqgUq61xgXKqHT3fNLxn5rnCVVLtR7U0TKTPaWwUYrv
WwVO2AaO4YjGs+NOCQe/uAFcK831hdyd3O0G2mxBvat/p0/mDWyWypweSUi//TiM10iShatzvm06
OhRCniuGMDBMG6mvRlJjbHgU8BFzhUnNOlVvZAwl1KyqleHJ3ZZpY5NSz90D/yt73wObB/dp4AeM
Xh0GXDwTenkQRvPwh5TOBIylkurQleP2FTSnYqgdhh6cK8SqtWuqr0qc5twHSKHjekw2z4JsHi+D
JLI6bSO9eFmrN7oG2abxD/8nyw/9fpzDK3G+dI/WWOzt1UPB2Hy0Ve8BYzh4eIzslY/uicd91jWB
/q+5YgO+lnhQqAvPQ9xSU0i/J7z7lCrIRM5XX23ZLI2chvl6gEHx3YPsZHWsrOmLk0dO4yTWHTIS
oCBFw1BRC02e32+DYe8XJZIhCCUEM81a/3nP2XedP2hcRY1WcolEOJrqk7AUcNwGNlOYZ8/wLrQh
ePbjPEm+029q7wpmdHKEUJkPFa3ejth9nBVoe9t5u8linONHev7+Kf3nwitNsuEyfD0rTibcffqS
G05dtu6DbAkpa1nHhca36VOH3n22G2jr+8ktXWmJP7HuupL11J5ulqdD9ZUsP4B8hCdI7IAGzLJ5
+3P6MdpxUldFuxK2ywsbhYhK/6iFjFS/8fJlHpxAkwD2F8Jdrjsf2C1nfzQqNoKWBGG3rK2eUEnZ
2KQzIGE3Tpk75AceHjLJd0g1Gw0HAVdAXb+TGTh+lmV91mTFbZI2o8zaMBkX2vHTZaau1svczhFZ
nAC536ka4strTwKSlGFCUsgo8R84t9i8Hm4eR1b5ech3lgc0eFdPBRNynp8DeNxPO5IJ2SjX/SRm
4EnPYxEDjpDzsstW79PPNbhDbvWkQtpL1ZMPmg70l/BLK3ytUjkzPnsyOj4apxTMgo0gSXszZuQD
THflOUfDkj063F+tQ2yvyTuNuW+35AOKU8b9gXRJPac/6nAgJyiAiBojm+lF3KPQmkSAVM2kuAV+
A730gS0nDr8jdE5RTl4BdE52JwCPfnMlJsQCSOks6dCHwuZde85XXRf2034pwWsU3cA1+BxX8nBF
Fp2U+5rW7nywSwvv6/Gv8/q1xDeMimbolkwJsr/uEnGix4aq6suCTY2oHTvwkEnFETpfaYHzx734
b1MfIyb2U+Yx0fQqB/vx5QLU9UidOYYuuKL6AyqigHdbLaBHiqxjR/1Jqt53CGofBHjMWBJSawf5
vh66Wm6oMvpXyEiUzD2FTjG6MVmehSaoE+iV1oHt3Z+FobSEyiJvo/e0VK2+tw96awEHME2N3Doy
w7NtEG57vUQDbmklP1qSm4xUbUnrXkWSZNi2B6U73PbOeKlFBAflXbEynl2XvWENCxlTEdxfjOBQ
2BlsK0DbvtTXv2X33OhRgZP7DYSsAXWh25KThHU8GqXJeprHxEz7jwZIq2pMHR7/OKKyTTPEgyRD
13s9HUQWcrqK6o0x3G3BVJL3FagpGdbHspLPABmgsEKCNDBK891nQ2SAMxzyt1ppUyZk8uBfI/Yc
ViOrJXsweHYPGg+EmC8ArwgeVnfO4rweEsgJ3Ajoyfg4V7k73AWdlfjjK8HexVHXGQg+7SDPQxL9
2+2D7RzVk3ZkeEMKJgr1of0ADUk7/Rqx9/icun2TcVH4kzQR7EgKjDxkwaQjgWtxmZ3tiP4bPrU0
CuF6Wrick2CLafbH1wC6tzDnxykyIGh5cKlwrXmLQlOu4MT77Xhxs0k8Rh7lsHJwGDLufQ6roNey
0wxd8VzEljIHnpZ3XiCYqnOxyI7ccSq91RTq7O6fvLz4aQ9iw2MZ7V52Bs1rSqvNRI7X/f/5rmOD
JBrEHdmSn/wzIWTs7WutpG+vU7S1zgOP/xTMgJl8kgOcGLq5dUSvlJPV5yxf8MTtorPi48xihYMH
foJVrXpk/DTNT+ZiINcRPhZwevKI4keo8bb3n34oj8iaulj9seovg95UyofqB7JPS7jbyijtLG2U
Tambs9GuKgB6rSa50mLeHuzsguvA/sGfVc/Zd+LjclQnDed4dQICkiEhAR8ck6bnZBbyX2/qdOfj
VXFItywOQWMhTdnQP2p96vFzRYLimWb3Ee2Ct7u1OhnXi75NckNho+gM9jg+LdXv2P6ycoFtmPhR
KnKEmWnTgwhdsF9I92HLyToUFxKvmqEF6m1JYEddhX8Ca+VFcOfECiXR1dl93hsUX8FdBON+zvih
X57q1kSIzsVV2cEEr5E7N5l9fuJQJbOWEwud9sppvnBnirMvQP3G2Z9dBs2Y7TnnUXPaLYnPYn6h
0w8ahyQoTOI3z1PghTwhXW1vDy84fNEptfc3pGQbu+rCxJrcY95gMSCUl1Jh5VizlsvsDyBo91hH
apbcQY3indbpAlMXXR+5a9xVmwbsDz/VGE9eIashvQCgwaR2GDEAucevXt1DNUoMxxzdsRnfwifb
BhsHaOmnYjaofFgdwV5I9V1r9fYfLLluwn3yj6g45q7rAAWfqhIV2DaO8Ic9tNtoRR1atHArRuFu
z1R52Ak+LmUGbn2vR5yvhJ4Gd/OoqrRs2+O0Lr/r62U8W6ERnwLy81zJTjPG+zPuKDBWgxLU92HI
UbWpu4mmCbX9JLcWvfiPTYOoxAnC4COWJ2hxV1WPijIuqTvDu+/p0X7+Q2Ak2c5amZZtcE6rHJQ6
HGLk1OHvBrNbbYF/xaQAtxY6PaOAGd9Bk3aU3IJoxVqleUJiqNIgzJK4HPf0mJHC8fLIOVMbuEjU
OvCZXbOSZw9z+WnMVkpTfjCdcUQqqog6wunSgzhJTTyDb3FaUhCBnwBOXGP4nlAYr5gjcB3sPSWL
3CQZKnAVNT4gcZvwdNGf23J+GX+hUCi6x8NVbVax1Gvd/zAvHvu1xcsr4Fn+XyGTEfj/LcVSWIHP
EQIe9xBPlraJCMZM4FAxQBQ7kKZ8+xkJx1Focgn58HF+qy9DTOU4i8ZrK4QWCGSQSClfBoMPwSvP
I6CvXnAgD2nWo1eV0s8f3AUvXYBy/8ZDL4CyBihQTBl8VQp1ArTv7pqSb0GwIh/bfYeITftQk5gF
sGn7D+yu9//awImIytlTc/i5mn7eZZD5fVeJHi3xMRmA5hNqwciDF/DDBxvupklQj5hBPhk83gtH
mCJYZSRkQ8UJ7iNv3WjsHaoX9hMkkFR/ofFQ8Dr4UrD1S10ulYNR4yPQna/nDATtFpggL/dzhEG/
snCnazuVcAg7VoroJiwGGfhiH0CEOTNowZf4Mtb4u6jacw3RzKG7362RX2zT6Kw/r2MXVSvHGUBi
cM0jM9pFcvY/xPNQG8nab16BwggLf9ef1C3va3I9jocyNdxHE3PhbakZqFQ83NdcUI51zpDBKPf+
Azcz4YT9+RViB/xFUiuYXUJo3+D7f5DdsNylbGe7KhZha8dMNf08Y0ATsxEvL3d3wPpuePRPCu5A
XUv1hZSptf0XSYb8PnYqFkhqxZCdoEfpE2GYdboxchpv9GTCTDAYnki9yHWWKfsYE7mhR0JgntkL
aVrS+vr0ZEDaI7qCH11k5NxIVCSNoUD63y+IBiKEk5SXj6plNvqA5NN1fm/zTwY+QpcFCToU5/cu
heaouiSwrv+owZ6WjuikeKRYEnFme3++MOvAw9j1rylejwGPtfaHNxHi0TMGePDT1Hn7fwDv76Cs
VVWf6QNung3pqznvn/r22M00KT7RimTBaKLbU/a5NaRP18DJXVgFJj6XE8vBOg++JHtXOv0rE0eh
4KsV+8iwbCEPZxJg/nZqQoguzPo7e0YYOlyfUGXNA320w7irORhi2Sq630b4ZpJXzd3BEPGlsv0V
GLC12icwChftTjY2NvB5c1DT2XQqMkMlZkKSFWY/sM2Kn+8fKBbLOptTL5wTJ45QqPHsT/uyXqIy
Ci7r5e0dNJO2wmD4kjM5SS7XMJkzcjSaf1KC02h939rakiMziFDaIRXYwl4I9Hr3zfcRrEt9OcIl
2NQJnZPsRFEgP12w5t75AbVrp6RMx9ZjiIWFpHIYNx7S0Wm59vDz6LoWADXwXHt4adw7YxzcC9hO
fStDs5H0nxgTKsT5A4GjlrAkXs2hu9fdP7mbqF+kXxZLvdyPNeLtoI0nCX2nOW2Qe+mCQUWpdcw1
RLsHSMOmMfqbhuz3xg+1jgmILFKEjjSikmKeJuwudMCngtLF+woAtkaxB0jO7MGwrs1dgP1w/c8V
GZA8KMx8Gx6rS4F6zdVpy+RrAaXh/fyJi9w2dlKYxduNCwaW8IFOhYgsGr5y8L898irIJEyoU7D+
ACWF4EkPr73d+4SHGzLRK3sqWZjbl4ltyjDzTAon3kZPvTd499b1nyHvNqfuyclVQBJn8tRhvS3i
jONr+8jMWamNPiEw+2EUB7lMEEQwqi2hKR3WcFK6gEDXbn3POmRCwXjfVgQBL1/XPgRRxAHmHgXr
78GImLw5KH9HFGf8YSTfHj23R0UTKFFHK8caK1er6uxTVJia7x2lCxPWGj6n7xF+kUWCj94y4lqS
KIevb0ikl85Z2cne8YIP5hLjX8c1O5WYZMZT3r1G6Fzixd7wUaVTMqhXC4AkXDkbmKoxvWzIUhDZ
4oAUJHqe0ofJ+V6w/PMeTm+WbDZZC8xFN26AiljDnShnaEhxF5Z5f+wpUP6fyPN6s6BbSsrkrByS
6fHnpynzPBPjh0kykzzBekbDlTasVat17DeUsI5tVoPItWyXKPWF9JeciJuRRvvtShLkQp9WYgiG
lqkz4ezneQJvl2AUtk6Da7x1Z660LsnEIwKzW12n840fKzmoljl8TesT0ZqvC9vX2uYn6es6OXoB
fykkW6zs/9+VuUR7ShKnxM05T3UqJp+yECrBQTi6g4RqxT4sH+ukltNQLcNKEGA/qlx1a1KtYshi
E1dn/vhOID1WF6lNL9iKw+AGjx2lfBRS6oTxEqc2yHIUpE7th6Ske1YOeZuBQ2p1pwEg+PoNvknA
3Hy8FKBN9/We0juDdF/nvlF/eB5Xs8BU2JlwDUJXolxKep6qZPvpFkeqqw9MiBOCfn5fMwTy95jo
uG0XS985gMluIyFLsBSMPbOCdjv9qkTiG1Yx8K09v141Fd9GFIt1c1rCHoFjsnaoX/q1nABonuSo
DiKyxkA1yvW6RbEc9JkB8O/whCvVzhO1Hm+alZOZ6N+WU/3v4RYqBs364XDVh/66lmYL5h4jjeyw
0+F4R1ZNCDQo3QjsKzgz6pFcAUz/eGr5MfAbtcGXPvgEnn7jWplU1M8jxz49ESIN5LGAtHr1SZkk
hQnsxGfeU+6Swv+15a02UfD5KBT67BmM9RbgTkS5utN5AzbM33aJ2AYbB5ZdhtXkBd2zpAepETXk
DPpto1U3MAHmE4a3174bjqP3qloHmVwyAIuSGZ7b97Oz8R6v0AcXNOodk2reqS5tCHu+kGF+QIVc
Ud58MQBfxcWUcR+P6U4wglJUWqaTQKDPQhOK5oUvn4tJH2gN1DbBAQR8s13HL3Zc70SI3epynJFj
4L5oMtxl6q41hPon8brZjnGuUKdZvxOmcSDJmGCsN8wvBn19ck0RtEHluU9cTDpsKiuDJADRQ7cn
3ph11KeBW8oByN/VqSw6pUtBhvi+SghtFi9Ajxdqi8KOgCHWS8DdFmGzj/BAWQRN8OL2eMWhmos2
9zq9Uszh+LorFXiQoxJfBZjt7PSLgMYdMfDbowO8nwnwzCZQ+GUg5Mk2ByVGTq1XIx8n/MIxTkQI
Ft1u/vHH1PS4iiT9O/ERAJh8+n24HA7TVbqYllr7cGGQhCTgu4grgNZK2hFaFnQHCJz7LHh46yA0
nCukYgyd9+kSdlyRptT3x78NmQOk24VNDDH1KnIWOKj9UGrHdsDr7RCzz4BUjvZUuxkOPV3sjQqg
R6bE6Ez2R+xOeHnMmJmhyVazl9jf55WsoTry1/+JK33kz7C0wICH6RaVqUviXGiJVkSrhqdk0MZj
lAHQVQ11u8M5lkc+2AvOydwRSuj3jf1Lipy4WmBgc136VF/F+caBFimAMkLBKbpp0i2P8zAjihx1
uMiBal9iqtl9udNVL4DPfpAqsZkNLIp+KP3Oh0yR+nGO0P5c/M7SQQSqHW6HN0lCShKOoYvOcNHK
h+7/ENGdf8LZ4nX47oPCtbKP3xmSLwc42CU2S4MfEvzWs/a6S2F30I5FIyW2lVKnyPOfHrJ4nx3X
M7N+w7bLzMUiWty1qbQrHasWJVhR+J/T5WMGPuFQMgctz3Ds4eUzeFVLySqtXhOizKrqu1ArscAH
jz//jRwm9aERP1OJ6gYWZ/lGS+v3G3AfBlwvDXeBnCUVhC+nRFpFWiLcuDoJNGOdUSebVrpj4UKw
PuclGhpbwH/360jVFHaUo1AsKlMhc0Ev71BiLtphei974Pe0dIWdPqF75XmvDjdRB9gC3q6CPbsU
Ns5dLZ61zU2h9gW7ogoW4AowCAGjQSDytpFFuo1J4XBP6gucvRt5DO2wGjpgedD6CzbZlWYXOAAm
MckTrhHEPIkUbULAHebP1UPSTsZ5+aAvTiIoBoBoCCoQKJDKhkjyZ993yf67X/8nA6SunPdGOy+N
4IA/a7xxymXFIMEesIHLGczkqn1cWlTNThQeMqkWh3R9goA3tbkZwqrzAY9aQBWC8IllbqSC26Xz
lhwHdghXX2OoXmR2SRM4u9evSACjzU/RtoWZa4+2Vl5P+YtnurDm2U9Id33hc75TbsE60vDk465L
u8oUP5CKfl5bNyX4YGMQKYx2g6Q75we+APJYPHWx7U2HrjaeuWP7PLhu/yN0/D8jCKdRNFyoQNaX
XjuQJRc86jec6OZ20ygyeL411VnBTpNd7jOm9dhuB+BY8seQZKdHInyE29ViKbWKVGgGCht98vv5
i4BXru6iIR/WE8leTn0aawAbIFfY51aiGcKXtAZDiuozDZTMyyW9F42aKstaMvKp1CIfYXpFg0TK
K8p3dr3CdALOc2HTgqHJz2CFCkrnF1lytTnheENRxNSQzqPd30DwgS6rrQmixn53iMlDGtVl4hnE
VzgFaoAKtzvk7EHclkJA5LgolgDkYYJa/49NGXPYxlttkgGDeqZUV+6I5DwZnLvPMoH/VvBQ19tq
9EPTe1Ni3Yx+ZY+7texbdALrAfhUHNZm2buhbxn1FkezsDOGi19ff+ZyC2xzvYEkyOtKK8a1r1Xh
HK3ask4Jk98u/2YFXE1Im2L4CaGGpDZx+SVwuBvSvfg3rB1S2ABPNCHYdarrAz8kKkKNX4998vWX
ncufjljJWgOwiSAeFo+9ApMlaJDDaixRjoQgH4aDIbEqeJntMygd6I+SRMiS2lHBmdQuNJ1qm2nm
CdRxLGctv2yBvCptVEpHXvzIbHF1AFuiKAK2GtG6J5QOpjbBS3F9x+Zfd/8YL+wjxvQLQPIjHcr2
Ho3XTrePOvkzlLf49oGu9KvnqVmUHCYd8qcAXvq2QgW1+ljd0Sb/zT6URnjgG6455aYEOGD6LD/i
MPytl+0K80pj2GmVZPK88dSrPQ6tjp1wbGTmEW+VgInHzkHOhuLiRZA5TdQCs6GXRZIclmWIRfqd
+gmJjNgnXxFqPa/kaxsZwkBoapeixI1lws8VS2oj90Ef0Gp87BvnuFWHDfx7vdiw0sjtowvb6S1x
v/rsskxaFUBFxgkF0Eo4IIavOsqgXB9qzG6tmj+JXZMjPOVwJQ8Gl4P3Lwny4iYOWhhWAwde4qhf
i4ju/+TfdS4FtKRznBoEW4lX6qZBFVzLmK9/acg6wKvnPjQSPNVJQJ3m/i/5Av7kJ9x2ToF2pRa6
Pv0vJSeGNNE7FZjzxl1bdW5VUXArk1G+yvEHKy1qMi/jYTlecNXMAj0B292XgZ/16SspZheNw0i8
Ba76FoPa3Ds7DU9URPXQsHf+XfklAbgZ/AtB3Z4h5B38bXAfnHylmj/YPegeXSLbncHl5w+knOUF
Qnt/pnB5ebB6TkXUNjwH3tWjT4YNlVHic1GF8VSdAnew3c/43xDRXKUp6MMUPJssAn8hpbHXo6/s
NvSpKBH73wT7dgrgMzRQ57AJzv+LzqP+QSwMJCI0jY2Zex+p43hGyDfXSklY9+MR243mJrNKKFjj
ZjttUsZf9dWhtheqc0p/pkTQEYPPC6WYs9YLTV5IXDhh8PMcH8uj0yKMludF2zqTwtI1f3s6U8R8
rUtMic9vjgQ06yC7qO66KqEk6yxvxFFO6h/YzH+rTiZUC7fka8Exgs7Kxnlly3wJqgngm13q4B2X
HnhGL2KDdV3/o/CAR5bH42p2mKp5gUNpxakkfF67EGxQsr08hJv1fHWbwtTtRibwcRlv/50QECT+
FeGH6HWDFOiOzcdQNe3Nxa/4huIkTH5456mv7zZB/3uQ6SCoAboQqtdZqCbcw2DacDuX3A9UePBd
V+THP23ztnk6gOebcVRARlOXPldQ7PtH7A4g8N0VSbP1Ed6Cd7jxn5tNvySSr45DJAGI9ifd/bGM
/skAYgS/UUwEtirbAvb3NqY2JLSUdcQQLDpyfrPbUjAhS4PyFf7ftavGyyQRrL0rYrTAUhgWZzBZ
0hy2sT0gHg2iZ2ekEJnSyB5iPvyJ+4QLzbLUk3glZDsznFJzpP53jj9NX6WS8xgpWatZAVD0F/E2
DcfqMSSAkj6uz+9HoYdrTdSNBzxADyzmLVw0J+7LZmkretlUgez1TfcYo3GTQWK3mZ2LYTOSvUev
iwFXGMn5CBUFSl6K0dmz31TLT0HMkoXoDTPxlb2PdJ1n0FCOVTuAV7koy77oycwFNCj3oLjc1xcH
PJHT+bMKxZ4TGJ4alUXpPSn0UA5mQcdRSKTwEVgMpJ95VRZKt7J9jzyCFC6fH8RUZKYtj9+0a6II
4q1QH1ta52MBwnVcsBezm8Hg6GJwBRwQ7Cftg+V/D5yCiIQ0chEQ03fgn7zAH761GZcS11+tWiqN
Pg1DlPJVf9XEfjKNO33Dn2SxL1GCsYo+vcfSgtmOmp+smg12zSONLHLl+k3pkYbDhC0uY1X6qYTO
xSsKl/tkn8rIRxcVfcn/tRmx56asUWO6rSDFQBHwWSWQZxkF9N1TTC5ZK3Crde4wMED0MYJY28W1
3Tyzt/pIvA/fsuYmdoI4cXilwKBKm0yIMnNGXL9TmafMeV8TpacISspmFBlytB0mM/BVwnLKiFOF
NWWfYhlS94ixM1ZQMCxTNlqtvJb0aTNecgS8yG4YrvTOHjKdpCZJn0SJjXmcAv32L5VOgnTBV6u/
RTXb96PyUj/2E7Pj+ppW7DQ/0pz7AHeUDtrVIbgL83pHx500XHJFTM+x/atWt0q3kTGLz3DGbwDr
/kNeeO+IqCge9zCoYKM7LJeycicZOsda22Prkdb7ECiczhhwHA4QmxhSP/QtkBkrcd+8vREmkMkR
TVbOLHefCysXu5qzJbTD7B6q8YVhAAZnc/JS6fYKkX6Ph8H4KBNspdpAbJA7P3bUeUoX0Rb5oO0H
Ci1L/rhF3beCwU6VzjSdM2t+sYWwznJant+FCI6d+dFgSiqjNbW1d/up3ewsXuePu0FG3Uo5xLZQ
ZkdtHoRoB68k51iCjZR6SMOGiJiykUQ6G5GMZMeRDMoieI//X0Gdc3XIg5llDAKqYQoj7lJJsvY+
aHPnCYT82jp83RJw1O5gRM5rGiqHFLR4v8UScOj4Zz1wEvU6w4I+iT9PgNmLkYjMOhMd/UiVVxNA
Dnbh9y+Fgic/2YR5/HZlW2qrkuFjV7aCvgEj5ZlSTlq6LCir/oSRZM+XOclmXaoWQxcqsn9Hk57g
ejy3BPYPVVHzVHlr+E4jHRxSzSHt00j/OjeDS7NYNipHvtTGvf6SaSa9ssFrpGiwTXqzBcIYzVNs
2PJn8rC2gs0f4AL8txL4ffZgwehFpAdohXCqlpBk3+2bb9YZcXeOCd2Yp5XeNFXMnjEdM73XMQBo
AXA4innOg5i0givIHRVGYhZiQ+kfj3u9p7UiioYewTFfaQQNS2NF3Dtph5c32uynLRT/1WGP1RQN
1cn23XmtqlPG71Kl5txgrNB/kQ54U6ltVenEXUQF0mo8vYAQDZMqLQR6Q7gX/i3PUhj/eMe6Yxg8
SZViIt+v7v+ypRf6zWEI5OrarQ+eo3srIiWIonh1mXsXF2xmibj15wYyFJCY0nJ15BbSAsELats7
H2JFaYx1s0XNsZ5xjXY+ddrfX6dPmpobaZvhKgINMBRLUDWSoSZlIVNzYFkWZw1UGzYn5A4r4zqM
HYq9w1ypFazvnwMClzgEulcfI8//C725Agby7rSlzEQpmQdl/blNageu9s+h8oL3GNitxnsqOcA5
CqN5OBnbzh63ZxbWK9sOzS0WhvE76eQkJJ7WgkupnnWy3X7fYhBU0vM2efHWosp5IlpdvPzLCgVi
eWImLwNG//5WEW6WKipLpTGhmFKlhBbAegBYnlCMUtOPOXE6BP/NEtF6Q0EBAWE2YwPwPOU3cTf+
rG9JMuwlzjKIfnfon4gWeJH2AOVEdaQg9FKeDw8YRYneFCdO7BlGBs1BNslD6cDGb+CSphzw4fH2
PYaXH2LslF9n7F9uq1fLXGMEI87lvYPfesUMvP4SCh2GLNNGK2fg2poqYw7iMaE5KogvS1m4FwM+
H1SE6XfEApUJrIe7MFgn/EOMJMCck6lkjCkxSZ710UBIbFcfKBxHJ6RxpkPpkYnkN0JLQdAOrceU
/tzc2+Om90QKF8EPly9L4m22oLz/Ym5r6W2H+G0WktGXST8VvSqROLwRxj6I2+eXAiwa54NdB3i2
ELmT2oCeCFLsPE+y3DkPVH+MkXC/pWAb7CYakUvbl0mLtvHDesWCyriuZuqzo8mbjtdUShZ8Q/2s
NXCiaTO7R8xvPYrxx8OSwTi/rbE/Im3DJiBqNYfA6TaPWjNnG1OTX9xmn9XOtNDcrd34ZtWnwGZZ
woNum4/GGFBU+dxPyA+8EDrVGzvslqTg9sHqBNgjGkPuQ8GPYkaDiDDIdq6p5++Bp6H/Y4Blf71v
VhomrdAR+puJOHeU2m58FODrfLr5tIfFKdMK+xJBRLm9/9/uB2HhtG+S9Tiqh15L/cdYNfedU7v8
T/8ol/a6JWM2STcX/P99ECbSx4EK+sEdhn2+H+4o9h4IB0JHv/iCziTlV3QzEbp30vgmNf/kJsSd
Pu+u5cCCeUAitXaodL6slCEUfCB2XY9YLk9h4EJmyLE02Gz0kG5pl72nf7R498L9j+5kHDPRMeXG
kLTBJW7jKhX/Cwdj/ZuKPmqxwePLaXx6NFrZHgQdL3VwlPB2aLAvfa6/jiUUvFf7Tl9zRN58IyFj
Icpat/qCp6SmTOjEuCwGtzjF5ypaFNPYgzt6iT+LX1ZB5HjeAIYRhs6kcduSpWHLE7udif9tQSZd
mMLcjShTU+CDmmVas1QXZUEN1yN+9v6fsS+Rgn1REe33DhaPbUhSjcUAOugOabm8EMUqAxcxFijk
KAaFyaSTVp7Vpi8dLeuFr7oDdgvx6mS/RQQ0wkO/6fqs8/bzVn5KYnd8g5uPXdthSN8mGXdtpNYE
1C1ag2H+FrJ8t3jTbxUwXIWXd8tXRtenAZugU/KZKmZfEdReii90n7tnCkd36L4A2PgVWi0+v6qj
aiAlwmQ3kRTJpRBR1Uryo5c+sze/4LrD2zyjXkFwxXjrMQBDnyzI5M//gug3dLHF+S7g53cgvVgN
J7jm0lGYpPLWczqmTOlTBBjUC1EMxsSRrQzzjCF6EWSbGAGx+QtFgm+/rFGKgGD/CoZPUVWvMtcf
t0MGH2DbK4VDjw5UnifdjMNXTS4i+NcnC+yfh7WTqMe3SLNcRXX2kIhRHy8SaGfHtB8YWIx3/sSp
1egRa3JYRSEReVEBvtDvKtnLwkDDGifWyMq0EnCNxJpMSMn9m9PkMnFrIrgDuHQicJIv15ZcJESv
Ivf2vynju+7hJYFFKkz3rl2CfPbPNIjOhgqytZ3QCn5SkbgjUp1QGNQ7Wc1OStLpmtmGh47AUw6T
BGpDWO5/E7scRSqa+BTkUzn1sxDrH6b8SRdOgzmHj52T7kH72Wqo2C6DEqDXe1cAAPXhDbC6EUGA
QQw/3vw8rdKw3QQ+g2N+0wi3vCIJ2mlKVjcce9kEbrq//DW66yjWX20qI9IIoaCqDELL4U5Rhu1H
c3H8IN4X7FpTlh+PQiF/xodox3Yg8Q9vUVRSPSY8SC3YZknf0gB1NJj/nn5eHSy3MWR1ZdJ7NzOS
ojwqUfjQei+VGVcC1HUfWUQQm53BBUEx9j8uPW1/h4F+emxXKCfHJ7L1sbxbmADbuYki3G+hXPtA
/HiMo2S84E/p1xFF0d04dphrsZUDzyZtsnlaqy22Go/gPEdSec3g9xg+W2Lm5w8MVmj4Ap3YnYlA
OybYE3qO5jKy6iAN7kVe5R6/koHGza9+QAMcWja5TfKhpNrAJw9S4pBO3iKyiR7GJJPvoEe8+cAJ
zIkhFr8SLZT4eGYyXAyDIFpk2PtSRfqMbU7c/m7ENZyRE6toyFaNcCHZUZUgMy9BNAkS4NkTet0U
Fq3JLLYZZAoy3VVUd7cTa43mJjFZ2LQL+xRdipLeX4gRxopmLO4QjkBcrjasJR5XDBrJzf9ibUGD
41E/9vfz6SSecE4iEEZOsgQZ+qkIhvXbph0UlN8HH815Glcfjm4EpjRwkKZzqA44iGwQ7xEHDwlD
0tkw1qS0wImk+RgM4I9ciW+pnMcBOYl7V2Wz7fYg1Lr34G2i50jTn52ui9foMnOhKFBjWdmubXq9
IOVVOWzwzCaetyCWB48Y30kXejGP0FtZtLipeKJUOctKcOIpe29tIzR9Lsa5aAJpfwpBHS+uMvbR
e+DHuSKQfQP0TxTj8HfUniimeP9uaIKQfxOLI8q8DcuzobWFJoHFTk5bpsHB/4rC2CsdNmRNsL44
2LgWH4FaPRBz+q2E19hbET/rdSkYl4uRGm3ePOssm91Dcm/aavsz/tnHttE6D9trKzKRIMjeLaXM
5FuhwEsfh5ZmpcFxe55HJ4LCWI4bHmRRwgkA2yQEX3I61WglJNp/VjStplniAdPM6h5c5MXjz9Ff
w+XjcniLUs4tru8LYgW762yMFoGL09hmlj3qz7L0j5M3PN4ytNoVmZdHmNLcMIqBxEJndd/HaUkK
q20KZXxkeiSaHG5fM4rQX/s9Z9Br2Ia74BnfV3UVe4vzNVaYhgvBEN1Fp36crOiLZsLBFdKknUgz
+CPSnaIJxjYbIWcM2smJ07w41XDdSdq7+SdhuipyYnWya85XcclrkZL1lq6DGOBNruuzD4LPd9WM
r3sK+b0y0wk6Jc8nkG+26MLEDCWO0jsATowcsEMBiMH0c5dEZLQs4h4EAYvdaG1mSYtI6xN1RqpZ
LsQ9LVadKAcePNm5RYdnxwuP2sO855QbniLgyTKV5Oh27IQbmg3O87e303MzcKTlI5OeNirAYVJn
U2ZYM7cm8TLLBlLRSjXcUwaUSlnOp8Rv7DSzOmbA0pJtA8UiskBNrkskPXtXnxvKuaOUqm9ewsFm
MiL4DFGGlQUfsEp6Z+khxN7+TiMcZ3owfgecCG4x1cNiFtNku58Rw+2DT1WkwsVDZQ/n4sryC52Y
7ABEBGCNAW2l9UzVx3k9UjY6OssvBkZKmcjtOgptFj+ZGQ3zlT5kyEgbd4x8G/f2iRGaTIolHgUb
dnNXikaKmnNGs9kYT8y0Is6kuDZp04XH/944FW38xqq+w5y9gQE+k22Zkflee/wcGCqbRz/pPOu9
jUb5LsjJu0uYLy1FIuyxGcmcnzOjFsoCuzTWvCEPVQfidhA/nnevQe7oUyaKKzn4jAFoj4zMV/E2
Lbyc00XAnr09w8cVEXYiPpyNj2WmPHYAcUudEeSzWQg436ZqWLroH29we8A0fXUZBy+1Oyjzs9BI
K7553ft3V1skE84B+R68j4HZX7zDZV6hQySdKFlcZ9ioTT21ZZ5FzAqF0qQw4s8l9xwQiDRGvEZy
FTTshpC/IG7ivFQzwtgtqVPp8AcuuXqimRwoTagidQ2T4yOqplhLRTWHBehJTXys/S1aBQISGdnJ
vDVFAZ9XcoJ/Vvsn1vG9usfr5fZauJUB8mDWAyHarn1K1Ahy2Gl6F8LgSfNb7STdrQ+eB8x89n9Z
Y/xmHXtHcgHemo/qbOWh4MPIL6T/Y1aVxmrk7Abe1C2imsooOUD56J+AjUnGXueHhq6qJE4gUjgN
zm4l3axeYPBGFgurUgIjtI8fkbNkIz0JVWQd6YcnRgxWAijFeA1DmZiIO6z14wJmiKby6L3hE9vR
CQdoWOl4lt8lnsDQJl8iTYQLmg0jyCj9m8XNviDWGGMpl++I0Rn6PDrpkIBmOlC7Yuqtzqpemx5b
vdXJWJUwc+BKYCLmsRFIY+N47rk1voR+xgOZF+taJUGBjEbg6JnXIvyTd5NzY8c+R5P7vRqVq4jR
9uYxxhs3jDwwV1sHZTKHTQe4vEGHgGZhQ4C1K/B8WyHnf4K6tyXs3qPIIFBcH3LVAv54lvexxpgI
37Xlr+lQH7JKOX/46uInOwIsRybMbpCaQ7oYS0nQURprKYM7zbt0baBXfzJ56GRTDUQ/GbFd04gw
Dmc4IxeiFnS+aHC/3EeiGU5bxJThnwcUUh+kU6C4Vbc4FW1jemyoEbXp0BjuaI4SNKIb5M4/Sxff
uMIY7Kx2sgxLoS+Yz/m4nPv0xFZE8HCOUfuTPUuFZqtj/BASsD8YQXdCO6Lro1s6wS1+VOxT0YDI
XOQD2FVK/rD6WJPgsL5HQeUyUQ17Nv882xvz257+HWYX4UD/p78rtlY4DFW6LSOqIyV3CxEx6MzF
HHGXXTcpOYhe2K5OZqspIqSSehjln33/oBMjRUgDz1LfFXp/EIVB0RiLZfT1icwbF1K19vC9ohO0
oNk2fBNH5Kh0b/hKbIfqundFnGI8MgDHSvVWiranVUNWIsVJKdtgMGW39l8MgpOMQs+CCCLey8rh
2eiXijqNxCRAf48FVFer1Rae8Oxz8Cvjc64kwBkexU/bptpsZA861/11t1Ev6+U0gjUoVK6DFH4z
3q52/okhxWZet6p6bPx6HRs0UtfJFG0gYCwcpfat2ACojA1ZhKRLdjcWM1LjlJj7FHb3BWAZwbzO
zRjxvCbFcMk5R4BFqdUsL8No00tbKPu1yLSXGfmertJQFK8kQ6TXJFQRPgBiwZzRiT9Im1obLH+d
/VGnp7cbDI02HNOlV4QHV/aVsv23WJz8in2oTNYjMUNzGCTHdslq9Sg22dF8mY+5MQZlrfCW3JFJ
MBpS7U8x7q5AiO3a71DPKOxp+eUKa58COz4ommhHgBHW3KaO12awK1DeT4uH25GnOHor9WFFAC+u
40S5q8vDXQdXADe5CmA6s8h6fHjxTTgvVUERJmNCcKnHUOvEzwngtgAr5RmfE3feVVu7ukxWsqJ6
NYOBOeZUYFc0Dwv3D+pc4ZxPAyf65JSLQ77QsYk6L0XzO//i8tWRWrvlOibD9mV53QfTQGIYj+9N
+hWyveV+MkusCqLLQfyFVOeyRihFrIoWtjZtvUbAI1mdl/6aNwC4qCJbsfSp5F9svQMwKfc6z6KS
afQp9vy/5H7Ye+/+DjD6PohZ8PuLjCsa2Z7IJMFT5ZlX1XSwAQwlHZuJuDWyjKBspMqmtTaDlzEn
mdED5Ubl2S0cpHXzbTC3HqXE/+OAmmSSKjhAdwJnrqdmD7aGy0sUkplX1SZu+EpApYvKrzdx0kZ3
qs3Ybb0wSbmUPy3Bok459/59Gv4JwMg9XUmNeBwxSBhc5DJPCD1NCFGwWg1u+ozhB7hee4tjSZl6
L+lO5SJSzvkQzN/ZSTBiU/keGT/K6asUGS4COVoCJhZ1mrnWN7A0wPocCGELs4w9zh7yWmxadEj4
5jC84H3MBMElcSGkrQiWCrlHcnUOQ7LosB575U8eelGN1Lr/UOjMAHSB9AXcfF3+diS5cZQrpKvD
YSAq1t5UlRxp13Imk5rfe6XMSWvKaB3mFpSBTENpqG3RBLdUmLVj21N3GdeAl2LJ3WBnpoys5V/W
pqo+0IA2tMoEWA5bjjs0OhuUoUWhRtKH7KIpoRv21bu7RN6EsxRw7N/kuTOeJy1GHif3is9JPPVz
LIwohk7e+STAwqYQf/Mkm9hVCWxY0q9KW/+tB2xwlGcL32CdM2o8UgYBAOeUWvejlPFwrD38QUZK
70fMpHnrTfZE7xfWKY/zFLSg3034G6o4YXvDgMMd5+wfYzKSemSpykJscfwt5sFVTF94d74FNmaX
kNdXjeVDdYgB+KCro2lhJYuVwGMcn5LhWr4y4vIayBJpfmeFXNpojpyqSU7vwQPBB1+ka5TZ7WEW
zD3CTDWyDGmGMQFxFMA3kiViQIsl664CndagmH3ei0xTpz0Uouj4fEPuUt1syqsIPdnFsW6S9jdT
qa0mSEv/aYbaIl+ySNMCcIYSCk5I0/oaoHxwXAJD+ncUQop/w0XDXoY3GpA4CDoiNuFWY3IBPF9m
S8cneVRTi9ZI9n2+o9fQAZ0N38HfYp/qPe/RCKt+SZXC34CZXTolEhyLQaBm9X/HjbVtC5SVE1/w
7ELriV2MA3Uwj2NtjxkTBGBOXCl5MilA/UMQoOKHmjUfzZWGgNnyh8orzXdVvpTy2Q+De7LB969P
hWXKl8N1QyZtXZQf/5AjIt/w1irbuJTnVnsjkZK5EaBtbqu61Frde+ML/5/Gx8XOmmkY2xqhJOF1
kAYHP+vjtY9JSSW1QKRQci1KK63lkn0taw46bLovgfSUmIpSZyFkMDCGXICRmOlj3zaLRWF8/m5F
XKV/2r4FbabySlnYP0XEG9dCF2BE4aY9Xd3k8s4fNZQ9/Qb7mOZb8BQAyRbiekTqCo64FeiXG5r6
fleiO+x5sj1mfrwPNuV3SmLMQTt/2so20gXMhimtqtm//0YffdU0JKeKHIU4u1gYDK43U9VCR/Qj
fOTh+rGlcVdnDYbkMODSaJy1GdIEyuckqfdjo9+v3sjoIBo75HDVZwz274DhMDhqHfpZMYr/hRXn
uPQL1t7Td1WOxAI/+FCdD6a1ixsMtgVuvaDuZIW8M6S1F8iLV8UlermYGbrxdhgX00F1iDcXQ13Y
wucagXZ3QLgZ/XJrFc0+5cIqvqqEXZGS0r51wMPP/QTswSmCSNg6urTCMsCHqFCwQYnd50iDQk7s
JBqROlgWp5/6cfB6faMqbkCjBUQxoOfKkThd1HrlKwZx0ThrfUv6/rzDiwcqCGHdqEUmrTTrKOBr
g4QV4U1RUyAYVFLiu1+b9+lhrbRk3VxAoujQBZrjy8/rU15iOeiZBFRk84WcTnPX6vUIiMvyyIs0
A5wboP2RvQu6XXI9sXLu5p+p5MUWOH9EUbbjWuzVzS9hGATdybyrquNQy3nmm0UvGMAbCTarGDpM
RPj7G2F5ZlCcsDICv1VY5dsoOVWPf7L7CdjLGNPoEdb9lHl5MzGd2kusIXNTHkxwzcV2mkiNrzYq
ri9uZXjVCdIhQL1gRKkaTyOSj3xstLfVMQUBYL4QdBpbO3F9I8ouVVl2KNIwB3H06yrg/raACqq3
Kzq1FaD+WPBQ/maNNZEN7ExH5q4PW9A4PEojBXb00VCx4PKW/6NQuks9qJ4PyE4oTLYiFqOigW19
AcEz+rtLSCq4PuCm4ecyEQM6etkohcR3QetKEkYhZUwVvyWjax6naopZZBfATwdyIpRMluJv8UhL
96yy5Bsl82pAtNz0KDi9bGeHXAgTAvsDFCEWQnlOVAGjBkiNGWpBLkdPwerxzc/249rAviN03uDF
Slk7dAS5C9L/3JVs7R9ouv++ael7al1B6cl4/rKd81bqaCp52iivfD9CEvNa19VqtLoJNZHsEKJC
6ljDfmzniKFPvKwzPUXE9Z+9yl/2pAmaaP4nFN88hBQ8rwfuRtMD+rtgtgFOV/riBd4Qqa+Adf4g
G41XqO/O4erm5St2KCkZPY3VGkJLZ7+N5BgPO14OaKU/NfWBCK57qv5pPVBh7sg+SGdqRSld0VBc
aB+ctn8yrKty/KT/iP0i+t5Rw4xtm1SLbl0PNLoz0uRDBdb8pK2SBMo2JtMbMKb+Xss85RFFRhKn
ivqlAKuD6KGMr9YCnX2jIITpil6grufYdaL2ZHi5gyXncAg0UiAweOypzn8egvsXHHGZuuJU5tnQ
X4q6FPOgMJEWWoKGXTk0UmbE7HW7lAQzHexfnGdKE9gyr1ctfjUezuztKBO3zWCJhvoL4VT1wV44
VLsiCEUKNfqeLayUHCH++6+Z+OLUV38l5jH72rIEni5gflZoifX3IYTzKGCeYOzv804lkBFtQXw6
aELo5o2x53TqnCPFBb5rijK6Lxn2mjx2vzdvBZcRXGn2FV9Jn7/c3TV+PD3jeidDBQdLTY1Vqvz9
fAY2XOz8T3fmR7MWXpc8PtqEKAZXjJUp8bvI4BdpxFPayoyQI7Z01DGZu93ApSqmYT2u831mR95Z
XUHzIrqYWQhIGoCDkmK+gSteEkffM2dKQZXJyPlApOAiJwkQQZC1eYqK8CL5yIxjTVBc0O3NG+46
f/bsaRLHhzp/Mu1TtH2xbQEyojqgRL2KAr8pTOV6SdZ9BoY/AXNddAkz5tA8Ufk+DhfMJUalfsFI
n6wSUck6djc6Ogi0EiRJbD1/4xC3Yaq3EJ8pyWd50FG5POKSvk9eOkXm9osBTSlUnQ1dZFhbrIFg
PYsi+39NxpXiqwaoEVITKvqfygFq01n2dZE9wbRCRJSdFZ++UIJ2mB7Vs/n77V4a1Kgcx4xG6LXY
CYKkBNVGxQ9V4JDqe+ygISGDgGJMlYqR+O7//BmpjhzvOG/TIWpDKJRHMbbs2KxbHWDnCryKfzKG
S8AdcncWlbnPTTWLkMIHsZAj5YIW3oCtRU79iITaXNzTcN16fVCMyAF37r9DmtW8p/gLjlEfRw56
4T8Z2pBMz1mBoFG8cZfv60/EPSfWe5TCndyMC6oFjsnKy7GXMBj0Q00jPIu/DU66u7JPjWguuWcm
EvLhMscVNObmREyVSnxE+Y5NE3utaOxPK2vKDn886cIE9QFoXsXlwYPyqNaqvZDAnixmvAbjJY+k
w1GXGP74u9QKyrr3ZaHMpJ/cmXR5VHMxNpAbwomfr/fMhk3nvOcIkepkAf8n5MtKe/FQ4bIwv3kZ
2p+W6DfkOWbi2zCiFxGyBykckcEgErKb/gFXlZwrYSaQrwlNZIM6QTdpoJcBvakJVlSS+WyZOUR4
u/PdYP1plj0iKTKc1XZ6qF9y+vzlYdyUxDgJj9I33eca71Z7F3RMWbKZLvAgoQaIMVDljEB5NGG2
nQ05gpQfMAS6KRPeLNbPnDOuJ9oBHMTwXDoiGeeAoydqb4z1Ab/2Nq5JT/zQAe9unH0jj2pWCa4n
doS/hA5we2CjKCpeLcRbQPV3mvfqVQOuweH3dAp8xvnlomMUuXhaLlpSHH0SFYKffZBEKBQb2SUE
nB0ChhWhXuNUooZYfBzfchXd5H7WLoQxs6v0zYp6b/QBMVfNW5eLprv/icUdweFb3d8KznMAJ3QU
EUcdneKXqufqeNr52cQ7XGPnDH5n4xRopUz5lrJQteSZLWzIF9wjHcHCKhBLTotLHES3mJHkTySx
7rYZk8TDJFB29y26Wthd/UjnumkOWtnUEpbNuM5LFVD/PPvb0C6nPOGU+IchCBxAnu+0H2/WIKHL
7lqL1CWERH7RHBDO0lAq4c77XdX0Jc/8y/uveImE1ggcz8fZTPy0QNM2vgL//Md3MQHgMtTaWNA/
TmDxG1O7Y3nW261BTJ+tDsnN9Y8wXc4jlnYx3OYGiSrnxifKauazJvDU1y8T8anagHG+ZL377YGD
gqlQxuRYgwphyzKc5vQhwUIMiCuYB4v/PJjH8UYEpGRTiRGt9yOg4GxdXEFLRt+zjXDkPj+n1Fj2
DuU9fyCAdhfPs56h8Y/GWSgNtOgGao2qODRUnerFZHf4vjSD6nOeU0n5hm0F19WgLBBCNnVr/1OF
WuyeSf1wU1u+0Ko5I3kDRX59wBwoyePSyhnHgunNRiebqSn4yN3GQIEwaLgSH7ujuZQBSKm4/OBV
PLvLULUqo8CftbRw1KocPiJOShZRJ52Dje9bKCgxyhuXzl2WraubGe7JqXZIEqkzzMzYujTybHUL
5RoxK1vFtgHORGqajDm+vED1205spLwR1HgWyqdxW47HI0YcI/DkFX0j6+sDhvhyBkQwi8qxQigC
iWsQWhe+ozll7kGDyeLMoBxjtbKp17mHgPKAJ81KQo1hHQu7igF5/9XJRpU+KjovXYstZXndvMBf
0HkK+AzVI4AV8NIKiEY1x8W8HBOnULKlVZt3ktUq2ckcWTQY00HuXXQ4qTbiqsDqMq8ZnsxceMp5
tVJziNXdhk0xOhe4HMVICtvBhvg+d69yN8hDaklJitIAT7Mj0wAu3Pu7sbfOiQEYUs43+u72Dk6W
Xgvfw1SWoV19tKi2kHwUWnk1uYPTuzTRBPnkcuP0LFJfBH4NIGHbKVGvWJHUwKNMHoBpg+uoJaDh
5Cp6a29xr0xX//Cc/0RBBCizfAOHYh7CHr/ar5ac+acyn5fhXXLaZg8P23UwjIb6womlhEOtxH2m
FauSO10AqRyc2pdXkZcuWO1Jo9hnsINgE1r6PtI3MjbsbU5QzqFCHEoVQJ0M1wEi7d934AfmRox7
DouKaFHhaNMZJ9h/KzTNzL+C8xSPjyy9LYqHiS8X4i4jDBg+jsmIu0ZcEZM3UoIGUresGMFV2BcE
Q+vEyBPd/2L2mnep9mDH2YeGj/BLapLSSJLsUj3jhHVjJyBm191lE47znle1mxeqFvrqajuoml+I
tNq5ISeXAgS6rsIJ56hcHZ8d+D8y7hPplpYdcAqPK3XaE+afJ9kjHCyYfhbwhCnnWkGbNsT2ytGo
rro16J1fvLt0D3xYt4wxiT5pn8MaWseYuoEs1OK+UOC4toggsqJrKzOpHgDV8W83BYDK+JCGNjXS
D4qzN3TPkwsybCaAHUDkv6dNFyuBvJSJWyUWUp5FzQdliOF6ut+q0U2ygbxF35cqFnpxuvoYszrE
JWeXn9Q8JjVPoABpEb1u0O3Cq45KXeuXAdrOPnG2Eoq/leejpE5V1DzeaqA6OprbyyqjsLGdbBSD
WD6HvWCiwGUn/Hspz38A5bDoBO0JVBuHf5M2LejSL1rLWNrQbjRFSP88S7Ua5AkIGv9vIobgZRK5
F/XCn09QkbDaEuvSoNTQDuHA5F3uyib6kx/EDNtS/XSxpFcdJJJMukDz2SZkD9INpLQwBfOCKJx3
JAfZuUufAZhNLmXf0VIBIOCQPQL1e0owHl2LtUGhXcyHWlfz4+M/KRww9bN//5tgQAeLT80FV+tI
quKNZQ+x49FYEwcUYdqQ6nB5qGPwytDhdH3bdYe9N6Vr/SSiqqUNP5QIzxszqEFSYyUyicc9cyBE
VgJSPd3Fygsp0MwABDFj78uTgBrClbf/Dxw6G7IPX/HAi+mWdpfaLfp2FMX48mGW2pVlVcvayZIL
KUN4RBrYVJiPk58Hha3cqfTLnpgiWOXdbLepjv7nq+fr8D1ItGnETCsl9tSbsE3Pkmnp0vNF4aFh
tbK2jHW0bOzWkjHS+fMg1s4Jgv35B/04os5+tn9YoPFYf1KuR4Vri1KdFZlqjaY8bNbwGL0UuicI
x0kqa4M0dB+4+EmVyiCxbkOJ+Gx0jRaRyNaRgYBqFrrRObxZSm3Tr4bN4mGJNZOQ++RvFYCOW6Y/
a6RguMLb3voDLmxDN5wZShF36apfiYLXIa+8TkUdmtclQooOArGWPxj/Zi5q8p8RPRRKt+rkyb/n
SPyhsWEb1MkQ524lwsm4tvOk/YMbAWQ4AWTiFeemI63WPEZ/2H0YN7vVl6NsHqSLlajVjw6eYi43
V3uC0ke4oh2UUDYIp0lO/e4Ad1wpmaz+ZX4qmRx4tQd77WlyBKUesCnfdaDsHYdh00V3te3mBf8B
MUNCib6bDk3P+KSGZ14YnF4uFHaJeuXK1fHxK6ccxWXgHqowGfsN8qa77LTTQ0tuPN2T87RKzGZ9
c4VmP9xLG/NF3Ay8r5SOdS6UwPgZZWpfNnj9tNkb2vU2EhR5nVtXCbZJeJtaTkVJ6W2VhX/G8Ljt
g1kCtwREQSyw9pgdGj08NcJGVSK6ukir6UV2gyVVh4VEqByFqrpsrFILSMLJQYA9reh5dH3x40l4
YJ0qZ8fkbkFLOJAE8EAMwlNSVDZNmCkLlDm1fk1J0hlwzdOHvP4dIN6c+8s6RSZoeL7wwn8i6G3r
nnHcC58vVWccq87TOsuI+FiANTqnrFiQcBhbpSQSBSeYPVIr8nZES8WjSba2JKEMsb78bsUevgnP
F2h+R1EJ46F+E2QRCHAO0JnggVt9Twgy4irdjhlOH7nTRFWuqzaTR6AOMgOp6OyJ3oZV7rZgnvvh
y5152Sc9+PLUTqrjkxfduy4ItoFmBnNZdTmI8cSzBKjtL9BkLJDZOOe6izWAhnsOBgN9wq3SSQhr
TWj3hcPGytk+TFHKZ70E0e3wlQpHWwbOK6d3flOPHbcSy+n4XpDBzghalasuiqMhAgCb9iNSEOZU
ekjWGumu4SYO3fFwH+9mBpLGytzmkzqeysJKDbKpTxjvtYy+plMFHY5sHVe7Isig1BqY2I5cvyIx
tidWVO9wmWFH1LKDJ61sQgO8BjNFbhH9MmLXJgxCJPog3Bndd2WVy0DePbS+r5Mh87iJ1+Sf3xSg
F3+NWDoSGG0xz0/OJiTIK/mRWkyuzDWD2ezMIV8whOMDXN+y5AdNclezeXycTvIISM9wzBQiocoi
86e0Xand4d5qwuN3sWVwYkt22gVyBijHXz8p5nMlRh0c1p6OfTkr3xe98G/8eGy01FY4XlaNIH8q
8XAJUScRIvz3onzxFzgUrJVt1b5KQVhEmyru5PE/wD4qIqR3tWyJ11oCaUjzziEj/80b0sQwfYCK
mHLYbKFHjdSyN4wx2qaZt9H2e3BG9CaQyZyq6sRjmyrgpLt5FdlZIDccNdYOQcMDXfseUzXaP7tx
QDOG0oQ77D3HeJFyrJBwrnQ+bGfQRXJ81c6kEv8zD5FaMjiKP7ZgYl6NVo4Qblbbk9pIXsdXlE2z
VNhokw7Iel4BBn6YLGvk6He9q3bx5sEySmxvJmVPKS74em2Egj7JfBt+n/FwjK0vEpagAyChflLj
jwEjCKfpbO7avMRwAuDEiZ6UnD7y+I2s0oskQO2opidq8kIEky9xDQZ/yW7l6QWp41WWUbeLUf6e
Bc5yV8QjDaWvARaX2FNCXC6BbtLT9vI1ZUzlkVqJCC8vZPyI+DYgQbS4QGFRzj6hgcIPZsSaGPmL
GUhmXeNFZFKfa+MRwd+0bq7RTNgTSXqVyc83Wk4AvaWyYfRQwPAsTRf9WQm0Dra+Vykkm3FHZj3s
Uze+9tyNK+j8Bt9liBVOi/nNU98djuHUmSSEkgPNnSGCYxeLnsvAGe3E9DwiL9XeFTCIk0jX0cjb
jN24If1sBHMVjz1LKuFxkpnJ1FG1SKrHo7NHlj8lH4AHWx8P5armTYhGNlwO/B7Vgx+40rBvKtO7
q7hgeUkKilnC4We0SP6fcMDtrpjpakXRYBMG7MIikyXL37eQRJv8u753tjbUfUPZg61VReqFaz0s
QIvguxlnFOevddLflRbrBX1qUmLdMhQsNZVyoW1oEqoBtoNRzdDsrtJLGJiFvas3pVU5J60NCrjs
68JnRsTzJXH1CZyfkveclWorLJyF1UTltd5vqT2jp7o12zr0Dyz2cqBV44IROO/66Q7cdsMFUucg
lMpF+jj5d62xsIPwjaSBIR2TSfp8Q+Z9SO04xIu8hPRrOHwAPuG0ey7rYjH9MN0hRWqJa/pkez6A
sso842ARpXbXjCZeFiPbLExvA3a7rmdc0kwhitDcgpD7LwfcbnLjmFP1//j5mCpDFENg5w/IeYDu
Hv78pRoOQXSRojAbftx/6dH9d6F58IcAIjUd6DUoHnYnoG9RBLYiX95xQwHslvoqH6/RdFy1yTDk
5EsOycDB5f4XxlJMguNVVbCGBAsOtMx6BWLQIdY9GktJRWem5GEUFOGBSOWsxkdXWGo8zD7ry7Ab
Tkac3/hKiuJ8AjWpSW3tMO+Mw8QBNVW3chPtzloAARSun0sCIY75VrW0BxYSh8O07LYQai1tuV/T
O7Kej0viRnxrZs7F/o7sFH08cMGYhQz9e92wfGiNnuvVUan9OXJvvErxxrI7tz6O3y2G809LYNnc
wkphloTNhjgWMxWmX/3v/x6Ign37BlZtnbV9ZzUIcWNgOKHrf5TtUpcF7GfeF5KL+Itejpk7EXmN
KPVYucxS0/EY/0J8tWmL68rYJJc1UhDL8XiszFWs3+vAzkjkacsNeMSauZP1SRteQUrJVZkbASu0
UoZBjOWLOJ9zl7DOuE0FGNzJO1Dhfnna/kLLPt8EaSZe2YHHIIee6O26j35kKoBUMt0uwF3myklZ
5dW360BG6rBVDs+U2kUjpI8DW4LhByC4pLfR0fuy5KVJTvsJiQcldemmjYVXrFgbNaOX8bgj0V9P
zAHtohTJsrJsKUxpwqPOzAvV9HGY8lRNTE5mMaAZsILRXq3EUqo31QrIEXN4gGsJge+OToXijW4A
iw27oq+xlS0zm3kRrAajDkZ+S2byPOhlaXPMc2mV1GxNOjVeaidLDcVt11+gBF2WasYWJw4qqu21
ReilKhiIp5NtAz7hdxmaY6aTZ4myaRi52i/ECw+NikVYGx/jTmvzz2TIgWOEo8A3SKrz6xDhIRb5
VS1V2TBDDQiHGAPhp+/vvcYQ+d062x8ieintEaZwSTA/B20ELTy3x3NJZO9Pv5ICcWFG6zIkR6tc
aHXNHYLms6juB/iSLL7lT8GL6EZyR9W3TPDDNxhKMJtqLB7+Twnor+NlUjIyP4hGQR4o89kHax8w
62K1Chq2tQ/xyU2UsFhJ2fvkv3GAcKa/VNsTyCY7lgn8iVx3ouOgotGMVlrEhgf+WCZ9fBOd8r7e
CSHMnxhjmfePYZV34BVn3NJux4J25U5U7AsvyH7Fnpgxz2AouiD/hQEn398jdoJitc7HjKoQ6ES0
8KJk2Rbrj2bQVoBlb+WoJ1EBM+6PrtDkuhGOFlCDBCIKCQWxLNuK0NuaLgA+HlUxKQy7ODbozToa
HcOzES3A33TgSiYTOegHBdn6TmmGOj+9Vm4l6l+CJsmQR00zvrzIHU/DNQG3CtBBronb1kj5ezhQ
xJ5tgi3DIm7Av3y7dxoCPYny65lGTV/+w+hiKZnjG7uLwXq6lGWVAdA2FufLu09jSRZwkjYEhX3J
iuqXB6prVImhJALhWoSfjAJh8262+DkYLkAthLJ13JQ+PApJdhl3V+Fc4oHNx0p4D/V2kcbonxMm
JVZK7njLkCBtC3l93vR7R7WsZBIdg/INcywogBm53pDBWmK03hnlN4TVOsRrMPmeZ6/iNS3dv17X
szmjdKQW7FD6gjEoz5FPEo0YfwdGBrjKMHPHo3vqA1wKnFNtJP6HxNF5vALp9k7A8yUJgJnrf/KC
677u2CMk0lKqLytyleSq4pqF7UJanF32ELbM2xiT/H+Z/7VCOhoG72xY6PIfnQyAQK0bx0ImBkXi
OuEoPlngyzMXFqvbEkbdOqywh+CkbTbsk7QVH+rbzqiSZMPB6yqFpNhVHEtOGJ5wVqnK51Dqmg1s
UXpyymzLm6ckNLHw3ZwdQkpLqdTGeBWsqGLfKpho5MxtzfUTXI4rAe55psfB3PR9d7fl4Hag9GKK
lFTfrvO/Q257uo2ypPyR6rr2P4mu1jQYHIeCIFjZmrpt8ZqycAEH+vO2vJmexUrlO7sMeLW9jt+J
4SY943tNjPHrCVepromLnYpPOPYA7Dglw3MOnQ3pDQudVSg66TvBQpJScCXQ+afv7vC684dpQh9Z
Cr+Umo1jv+okTZcD9gpsWFOsJk0ijeqdTWHH4I0oVFtDV/TwZuDftqugdbfxwDe+F24fTbphu0fk
ryO2wvtbioKFNGFNPXkSvv/kOmL91yNomXhHH0PklroVHgcP0b7Bv7cWgjd16R6VH9mRl7EODBFk
mHwVp8rgH37Sp8KmJKNsB2I1taxAWCyhDOhdWIv66egne9MCDap2HAyIK9+zJ26xvw8kECzqQFbC
MUA6TzRQRxBp+xVjSTs7et1761HQB0z5HfF1f4650/DHQfUda4pRioV8efynCPaPsapXMylb9kwh
JmD0Bb9xgEJAiDdItP19aRX4zEyXZKyKbJVKpoLfJmfq5hemyBo5bGCIlwtC08GiuGeLnprpDRUy
LoDFRmBa+8YApHV8DjlJpcFQuZd8Kyy7WdpZPGly3znLtp7OHAx8kHOUuLPuM0wsvq6siItIbTsO
2zVtjdeGSQngW9iOQ4RAlXhVAsPD4v6WsJkTABHtc6G0++TY9t9ztHiVM6G64b+GUTo4tI0NxXoh
KST/DPbftdJV90NMOcaFeTfG4V0hztAr9J8Gq5hiutTizRnhwpirdrs9fND4U23oAdaAWw5gdQ7c
1TrQAuqmWptzp4j6822UpJYCqGBP/ikSjBwNgkmMtgfpqbH4On4w7Kx8JEWsCjqpcCK7VxBnZji6
UJm7fO9Qrhjc0vHZzgSF+1DINTUiqUoEM6P5bnrfNEPa+Tx1JcDb7/tUlKedkGtyBQ60vY9KvEoj
R81n6qSjdtnnKBoMeehLKSABJOfXbwskKJwdrzax134p4tJ+hm+3edsfSWg5rKV/KDL57gqLIhxP
ConZLoYt07HFdjQgtww2cMC4o2LgwdOQcvWYZYuNzCCSXoE4pLcCSiDTGx6AaRMmBPSh5PQrAmjf
3z5t80xR4UVi8FdLkdvYppHutWnWAqcQ5fMzY54l9FrvAo4s3p0nbrno3aHyl7ryUlr5u2LkCDSZ
uRYdWHH86DufaQUdgtSR5U/p+Nwo6WvftFEQBqstoBHzAakBcX7q3uEmBKFWvdrvqP4XTbbI2/+m
dd9eOjWHzVtd2lRZoYzk0EG/Ulmn6AYIfZRVc7pmLYbp7HeQHiASeEFU4URs0XdeReyRQM20alRm
NFbHOF1BTOiPiHrt2OPu2PuzsbAz/6Ae54UMmxJifTbfxFN83dKh2FDMH+RJIJcDzYs9XsURoNeW
hYxf3ptonCZyWLA7lHntaq+b/59LABdY6lVBTzI9Jc1UnTSckej9ey7dQqVVEuWNGUja4QbUZaZq
hbe6bXm8b5g/ioC58s5QwaPpKc47MX0EQONGo0+Qz77wzmJGgQ7n64K3AAOjnQN2AWJiZkXxkHI4
H3zXY6k45Zklwz5tPz83LZ/oIY2maKmX0SnpWyjOuniVvOmfJYFd6i3WPOxYsAspi0LlnTQONyrn
Z/ngguh2hh4g+SRlJHUpnI9Tbq2frqqg5WuGmi/vYxb3zayathTxQXoKsPYAgO5WE2ST0KylNZ31
9lnICiRSogRWSPWI0Xf8yrxuubq/vSfTDUgtsihuVkzYayk7ZXAVVsH5oQLgmBSr1R30cjRHskIT
jTcIwr0saIRZQbf3Wwhb4ZbjZCHV+gryPjU1OMQOGxkHA3OgV9OkLIcWgPJsyIG7RXj9kKyyUMSH
tEhNJBdUTk/7nWCgxnFLCOyJ7ljFlNj8MJSDk6zIcZAiCTHsYNntK5RuSBeN8dk4w2eZ6MUPBftk
IKTqvKF9yAoc9DuktfGpnVeruAcOu2+1SfG7fD9RjCNrpSnjR+daPqAgeyXlm9/VYA6SAsl0XbaQ
RkiGtRY1qskgzOWKGE73kCKfcHJA0qndarPLU1u8zdd8UxoLYcXUTtr5fLWdliuBq0OO4NHPgqR7
ljUKBkFt4D39hWiZwAroRs+2E8hi2vN03woaKs2oYiUznXlsDS0zK7oi1K+i/+r39y7UhqYEwVbC
PMMpugHqvjgyGrilFIIfIPhARjZ74tEpd34pJNAciHk2tBAHnGjaBL/hVplTsJvJ1tUuOW0rd/qA
079TrXaDDNb42YOpfZc3GqBmrOyzoE8YKDKGXbi88iLfps8zzMsGrAVosnj6cVrYYA18+8DENirY
rZimcSi1s6ZbnmPFNbQ9HeTaQjoUM+nBag+6etKyuBJ5CqVD4TJn7aniEJxR/6El8GXZvmz6kxc5
GYBa6UJOSj+vcsEXJeWpCrv53YnYndgTArCRQ/isTQYzRvhdN2D07mGgfQ2RAMXsgp7HxuAJlwtT
sj94Z9rJHUIw3RahPsi76g0m3yz3f5Zb2W/e3QrqksPNuEKhgFvCSdWIJHyijzIpH2kgU9ZzQJFb
fm8ReF50M4vG4qXWGcXfMnUkvZUZCt2Z2xfcrQx+DnQK8b1SyAkGmlf21yRwMa9XYP3hiEs+xzqy
O6gI/2LcAVRcarbSLaTMah1VK9DIfeCoLk6Lo40vI1F6jnTWGTflgHJAeUOWQDJYw5+b9dGmpXnc
wNsOpUL4tuIf8ZSikFiJAQKtoZFou0Z+DQlPzPBm2DEetg61VYK1C6zBbO7js+t1/vKKK6157Nqn
xGVoh4imIb0Q4isLrROdux6Z/o/i+SuNvKc/hBOrcqHMCddfT+e+CKP2iavqTpzd4HWMNYia5pze
lj6bp8z6I8KbS/4XrCqYvEe9noH8XmCfZZqhxhuv86ZTCa6N3ZjJJNERDaU6EhfEgIZ/7Jwgv1WB
1hoEoz8nWQ008Qsc97BFxQOT6Fd0SKcCq6JP4bUz0dpaEji5oZL1chWx5FDzZYj0eoaZxq4p2BJ0
cmlQpIGdxostA+9Q3X5uAg88cGLAJ911LHILBQ0ULw4Aq8Qq9ule/uintrWo3nV4WbI99WxaJQGj
xwykhYQ/SjV3lZx21YqI64tyQBMtAXGooI2PSFgZaw5bUTyYR+t5hn0VfrQtL1itqqjPwEArELTb
CaQP8qp83uVT3QR3Oi1h1KNHn4ahnA19bQWi5s19+J3GJyEhpeGiQiVNmbunlyRAY/gtS6Bjl3/3
jHT2aj+r+zn4h1SOYjn4kPeftkM4wIQiGeS0v1mbE6h5Bl2bC9QtrJw2fwmGtPy4EAvoSZJ2gN9H
rzmMFwc/kvzdDxExAKD9RS6O+Bnou0xwkEzrXqNAdYBjIu9uzdQwV6tUt6dbtSvdTL0NKmjDowPb
IWrAXDdB9F/DpY7qcgHfY5aaog0nShDW9S2u71N6QMEGiBA7vIT1qqCRQZrbC+I+t6ax9mnjshA3
Gm32MwDG51OdkB3MbME77tVdjGvAR+nmz99nSdg7OoZZgBgZbeU3jRI7wKE5ZyIuwNKXMzSD1GBO
vRB7RJVO/zEyfaoJvahGNhQqRdDVYDp0qxjfmhEneqHRlumK1Yyqx/d/TlN3C1hqINQJjQ5I6mpR
gh6TIEf4SyzR+BGUF7/ct/RfOXekGrH/M60LuY1yZhLKa63KL8N7+HTeCTgRBXPuINDiDk1YgOKX
8X2rp5z/bWOUDHaf4oMkm6WZa7lYlOH1eeW7OnztWmhOFYpyhNVmD+CuccLxBZGFTfpKS37mJGS9
S8S9Voc9Vr1iAWVHtK4NZH3QDWVOAxIoHVmw0acif1aCIU+BgQ2H8RXUeorYM62NDThFWMUflzB+
WBr0zHmxkQD5wvHodkjbxC7wVNM5A0xNcMweyhgIZJtaAWypF61wHRshdpuLkmTjW9r97tEWBJyw
sxG6l6u1mGVXGw2roOlQXR8ZQVptA88/rksKnFwfD6/w+X1+cby7zv5vlRyh+5pKGkhffl5wzR4D
BIlE1cK90dVaBHxyuA4YWvVcsObwQnoPlAelPzXbNVGwmbwV1MjCGC2yhSHMCiuHcsYPJidTswTX
pxrnUd9+j+naF+uU5eVeBnRxZuz8FDQmhheZRn3K6I7mkdYVWwnSO1LBdOAkogr6mXjn2Ia3CHsk
TKC0fvI5uDQJ7Wb09GaX4QGr9fhQnPrSiYreWRv412ZD9j00QO5gkdLaeIv3fDT7rPZ+UDqyo/A3
2NCAt18uAebb82LD7JtU1rX4NiLTFSD4JcS6C+S5EOHGG8wWqt9CbTciIB36ZFO/DZZI5YCums5x
lizbokR8CzY25zYIni5+Wv+XOzZpFsYrz2TcOYS+3Hasm88bkJ9j0nr4vrD9eKzEGbojmhRYgqTC
ZOCJLiPG6xpU23rnQ7tu6MDu4GUzD1sWeMyOp2TBjgZkENHmKSlCUDQIzvi3BRujH/nNzKml6meT
dJX4WafdDjNT/XTjzmuNw5Dvf/WK2nakENXVpdxRtJVjDgoqiH+hNdeHIYcuKsFoU4tzMGNVXNCG
H+3rq5VLSHbWl6aVob3eBdGy0gymjSycWftS9ZUoFwUFsUjB1mUsbA7vpU76thxT+kiq0WhisWkx
05ThirE+efDUqFptw+4pcWn2gslgwd0YOUK/77SGQDVznJO8EFpN05fR5U1HRea6LMJGgysGDOj7
A8E2EcpFeyfO1mailqBHHARFMBlZePU0UxpD4whcRYNtH7dRk7+bAGNs2xXUtoQwbTlEZuM4VuBR
JP6Bjf2f9crwPMJ5Jxs+B9SvQmlQ7Ee8KSt0XqD1lOTZBFMEBeSV+ZotjeiNWagKm2UJybPRXQuq
QHbVLC1fMQWiQLwk5C6zjRB/d2goQ2LcuLmYlWPSkHpaOJLYyAzTVR2iSDrOT3t4FBComvZ8f/DJ
IuHVy4bz6ROVYWUEQ7+lS7bozkUnRBX6udMje1scbMppxcKekDHgd1Qhwqus68yLpnroFL1Z9xHU
ispaF7Z3OsD0V39AQZ/Slks/M3oKeJADxc513eQbmnW7qwsLHpM+qMzKGfqUdz2T1m7lLhWlXGfx
+L/D7bE62Obxyf4sIUVh/bfVnhGdyDFNqUDglkLJskQRfhHGkfneT4AjAJhOl5tBaB/5UH8ASnMA
wyntJDx3gMdNs9MlAVKhMh/I2TSn+LBE2uayueGed19aPxKMZkzDBRIzdxrebKaxC4I06Tf7GA2I
5Qq58oPJEyj/I6SBm8sq91N70iOJWBEZ8383ysfZ3P/iFmNpt2OzeZE+O8wc+6TMonZ18aQS3n5w
eivNTPRU+vramXzMgsbqF9MaKBdUzLYsFExZPuWQMW4R+MJJJiCeZZww304cjv1aqYJtmbID+vPT
IKAYon3xS6rk/x+GBsF14zv+Wi3NtAYUA6CGc5Ga6tJ7L2DIXt/Z4igsvIC5TqRMg9sk/NWN6OaR
C1RdkKA0QT14PCrvo55BX9diRcQyDziG8tA4IF5i+9xUnJJEUXNS7+lGXDWUoVIdsgQTrsH/vXcV
GiZbYJVTMKIRzkmniAMOnx894wZyqDFtZQjzdw08GOl/RKFHKJ/MtJT5slRc8f5MMyfQ5UcqzBcM
fncNmkFh5uzpxyppJuOiTKtsftmxSFjokvTW+UO5G+45mNTucJgyDWfGmsEE7dXtoyJ8J5wJJ4We
cxCthOAVTXOIClDlVCo75bs/3OsGmuBmXenio6Kb+IAooAfX9lQb8yNY9T0Zd6xaP5JMRnXwTeaP
1ih2thjFJQfoI7+0fJhHrBBTKQmHfEbH3+PseFpq4jyxzkKR6YMxkR2FXPwy0xQYcdrgJe5ETYfE
a0UylE2qSULHBQKtj7IijVntnyxO+8SjX39LVxf4gQpGJcLx8edxvjLy/7Euml5ibDmFzgDSE4Je
F2Jg5Ofc/WVYXbO7DI0ozlE288Y6+Wh+vml1/h2snS2EXfHpqvUSXRXfmajcXKqnOWCYGMUf/0Ok
r6xYLsnehZiYYIPB7KJ+dYuRJohUD8/6D1LhnU6ox1rOaw3h6RoLZ9Z4/bL3vz/Yf8DW5uqyju0w
H6IQm4Vbq5v1MviE4mOJIba1IPx5OYSPpgn0kf4cc/xLGL4+l0yrm9ldhWO7NC/1+XTs/RH4wlOq
Z2JVv5KYIg+SjqbrPuLES/iEDO85w1/nRo1qI3/5PAE/k9s/dKSl9s3SqqlzX1bcTxza+Bbf5qX4
ETvFN5Z2kzEOf5D+r5UBhpzm1GTYy5yESwgE5CeHmVLhOPJIPljY0ZnByOVQIjhdDt+5eKO7nGpW
8t/uTlojlEipCG+xpTlpkKGixfX+mvAhv4O8qU7x2h58ECzRPQKaBrLfTGYMiYf91T1VUR3VhMoN
+WSVqVObZuTnEEwTHNAqNpxul69NjLtzv8YVVqCYkACh9jKsphe3URqY+/biAWi0WfFGlcG7RRxY
ap6j5G24aPFXdGulJy8X+vBz6dIgmJjeHH2tiGlvAKSEyuPDDFDVz3UG6+Z6BYn6Q9SHohrI+0ps
aJmNfXsBec4Xsg5Ybl8LVAFGmhqqA/0hoQt1mgJqJf+Yu6+ARR/g7oBS10Gc5+XRACKfQnHIiLjN
0fvzBF/IUBA4/DWaE1X4HQRdlLP2zelpdpf9G8BOZNNy96pCAX1tFrH5YFLj2xIMWA3f7pOjn77l
NLmFIEqYVcWOptvDINlVDlpDlcgo6rM514AaaBLwwNP5F35izZS1ai5ouwjFzqx1bV6vDmCdA1pQ
2UrKE0wScXeq9i+RIUoEzZMfQlhE1xrtl8+oUskhcsWoqSxUpNyII4ncHkPkXl8Y9nknHBeTZqQA
TywIEdbW+YuaYt9nyKImeEX/AeqpGCmx23Gwksz0y1NhFbM6kRSWSVo+cb5gG6HFLVZxnbGKlkk/
JN78etfot52XE/zhdFfhzPKhSHfVZx/fmxB/D6igJXVsbp4xeeZbbKugS6oGab5WK5ni/cnh0YuM
Ajf2zzCUt6uXv92NioIm8v/kJh+KV43iGG0m7Oa6nbYzEzwz3cKiqXxmqrQC75oJngzRxM2Nsd4F
ip1GEUXlaPm4aXzG8Kd9mFZfSyTx1S3fUXK9vM3heaTFsUx7ZlWpK/07lJGLr6SPSl8rVap8M6Dh
OhB5DH6VNDZFBWmNnhl4Zrvop1G+HOdns71c4GsX2LIYCre/TO/6qYgaSNGDkec/KQFA3q/DrXFl
uo7UnBUGUAIoOtDCES4p4XM4PooruJ5esf828wDNaCo8dSFY1ZcmCLrw76DSyHu2rst15MB2Cppu
/c1wH/4bc86y6X3xEDXSZ2fHIRM3q9z/sxbLgjTqi0qmpFpXmOR1t9tyKiLr7NrQEmXkzkWf21wF
97/XofN7eloOAEJb19j1OZkW1hHseLvNBgsCkrzRCTZe75EhSJuh5TWaL7Faw1l3oXqJ1jDiw6cp
yWuUhFWkQRXLLHmeuVoacrpdZEFzk02f0coFPzWbuoRh3nfSQhJdfQCMOmON6luLqvfCjt7r6/S9
f9aja13p+33Ei9FT0rePtLQ31bOnp9D5b1hE5ysbMDcx3tTE+JRaSo8293YRIfqPfS5l1rP+bbn3
dYBG61B4G0Se3sFx0c8VNeK1tnL3O8qR6r6Mia1df9HdQhDgNbwjfarmBUbcKyW/2h2m/JaoXOJh
a907kiRH5r5ud1TEyja+mmmborYOPXliK1ssbN1W+Jo3l1l9nbGdYAxOSNPHsie487dV5mkOHrjA
YN0WABVH5R9UaKhxL99XCp/7LVhUMXHrISqiBEEHbjuR1mIdhSaZLjWRPTqtsXESwBdZ12Zk3PN9
bzyTbk5kqDCsQhmJwGzMY7fkWWP2sw/pgMTEnNQ0DpkyUY76RA5ouLyLZ99zrRLfOGNuJ5AJdd4s
rReugnrHrrL2McskY/XjAaTtud2p3A/vAudPTBAO56g2iefvX3e4qKQxYaHDqQNzhsF9+sv+zKbO
0EUvkc91LIhaQ8S2/NJu4S1ZwRfyaewIuoE0LXDqS01mmRLbWniV5HT+bmOmBwR3vBlpM/9VFgfR
FPFVLYs/NXnv0oppPP8GOUWnfCnAq3BTgktAVXnKKzHRUjJSYTdunRY0GtFIXKt9lhwVmIPnI6YV
fsD6fCooRWvlKGp3In5Ka43s7fTA5LTInuenxCPMv5lN2rMakeMh8dsLIjAMx/42OTezWegj0bX/
KIeQTNIEpq0rHxCJHc32c9p3GV2Cfgv5eqqdT6oBGdPkUQTPVebzkAwBXWqAKak3pwoEgNLa/QMh
/VexPnq7H6RpohiksbBapNg89xJbOYD6MwWbXrSstL96rMnTych5doOP/o9SemETI5cUXxS7nMrJ
HFVSBz5rvcas+sIdoX4DPyB/7HgT8Ow8/1ZDqoxUnQcNlnDYI+Kp0pSWBrlFVas4WNSoMXAAZMPr
cknMoZKRBdORPW9vdYzOOtXc2SriBZG3nILHwmbfLky9r3ytlkxg82P6WL6UUHy0mndxA+quTB6M
ug/hyLeEoaExasJN/e1VI+JgX3uH7GQyLkRCNFP+LNtEPlPlm3VBkwncRXQXx4JCyF3j3pnyDOFY
pWlAz3sSprw8m3YhSDc1f4ObYNQi5vq9g64VGO863/v7LOPggZP+TGi4473bFnSltg28NSoqyhPU
B3OxT3wsK0rU6dDv5cfhtjrcHGskcVbeEd8zun8D/AJ+CUlTBQ2hLBQ4ccI/8i1g/ULrUJZ4kk+q
bAa7Rm4o+UDIbVYtsITlBX2MT61wB27L3dWqEEhXal/xYx5IzcWSe3q8PfnlYy4D7HCPkWMiC3nt
8ijGs8Cg5zEuLFNGn9Msx4LBFeZ9nPlj0gdWKB0Q6iXfLP/Xu8CO0IoR2Uceg3sE9q3/idViSzu+
rYmXSWVEowHqZD/lYcoTkT6BlveeTAPqa7oiPs5xpejWAHoPyRMZ41D8qXtLkycN+3OsWxK5Q6ZT
iNJvWFuS4DYlcIMVJi76gZCpKKN5+trqPEdgXqaMSvDFl31bRKS17zm2Wu8y9oVmEoZK2nbtaov+
NTevyUUe8BLzJaU2FWjHy7QKSpTQRBTea6x62RsuMr6pFw8UZMhIl5bhPDJMacAqF+jQLnozDiFt
pBMzdrpyangcQQ9s+fG8HXmMpW2aH5Fpi6d3obZ5LHuKiIjBIQ3q8EQ+aUXkU+Ceh9z30GZYosHV
QMzDV5/4HKS+uDM03sv8uEg0CPBgv/rNg4HN4Nonb1pyQZPAGt5p2HfwVjIv+CVrPWRr/cPoTZZR
sUpc7bjFNRRSk1cqGMvFo/BM7p08Zx19sr1VoBQGTjZDgygnTqHxwtVNLhTZTDLGbdnsC69vm0fQ
FfXuEF+y+vC12EXAqH/bmwaZMX1dJzXwR5GkDF5m8Loc6xUAIrjfvoT4zglbOEw6NRR88v9iclKf
3BRGBQyyeCXHrDj43CCjhEccEgW2vWpNs3ZKpKeeNnEkGiOFqN2fKCtDmz7aj86eMdvK6m4Qvxvh
HLd8Tk9mbSZNq04XyRe7H5YjeTja38k8pLNoIGP5bUgGsNxEoQMKK+1Exg48nCSwS4XRIbhbbMLe
SXHCq8Dkoj1ZP3pDcxmUUyYgwwlQujGeAbzlyRA12+puas5wTjTR6DhJvdTffYCZ22UAzueZaUI1
3peNfpPW7CDUEbKno/08boKJHAkYxE+GTaHT7jTthRJPcBNzHWNMo9tk7stIc8OaJ5nm7ryDtgb3
4hS9V/pG84GYlRLpqOJP8CqG1ibXKMC7dNqe8G4nE7Wn/NyZcb7lY0eQZI3b/mqBqMCwlcTakBDL
Nws1sJ2T62cz9eYZRqFV7QB4daqFi65WCebf7QUsA3+yEOilBbzHsAWE959Fn5HIOugFDCV5xsI5
j5a5qTo6Os21n2GFBkp2Pr+eTrMsupwCHz/vY1/BYm8qi7JO+4nVj7K5/USalqK5jIs3n8JVK+Gd
a1DgkFSy72NCTQL6G0p6W5b4SQg5F1oeOOE0PmSwsXq1UqNNJxW1xmGrNbJwye7vzGD4Ue4khR//
nmJ548eQ8Y88+86xIFtcEABqWJntBnKBT/OoT9KB2ow+DyuQKymtncXBwoIMSO4TNHtiTo2tS3xv
daZ8Sb+DQqbrYsPoIsoox/LL4lELVLEe94mwCa6SuZ0lDSHRly3bfZmZ8aWIq9oS2kRppm8/4YNX
WihTyJQVqHoYdT+QWl47R2Y/zyg8CIbIBqYFKa8V7aJqtrmHJDbXSKSS0Ca3mE/S/bGcWR8ZJGnH
kbMfWw5zA0ZK4gryn2nx2Flva4QaYMRCskEmB3Ht9q4DZww/Z47eCkCixVVUFEyKckCFfRVXapqi
NezoZ3HND7ukw2fHiReHG3cR9WdLV/3m98ZreExEZjaCl7LIA2SemuLUiGoMQg1b52xc5GU/EG0J
13+9Kv5fv8/4OhKT5rydrNMjzSGF52egz2x10Ax2JEBX6IDotAXCw+IgRWrd7bTJdK9YLHIEWiHL
PorL799cTBiHXRTz/Mb7rc7FDqlkdsRtw9CwQsii80DfgmGRDDDYn5S5IJQgr77dU5cZob4Y9v8u
uqMJHSURS6ofV5tykXA4NNEr8vhYKGK9wjlyTVbEhmfSnfChjsF5RWNFBhfBBWfz1UkywD0yqvxu
/SyLdLYL732EianoWUHF8cR0tXSQ91XvrzXPhc0U2nplaKSvxq8y2yClzFwWduB9t70iLDU1MfEZ
wzyV0NNjBnWKINHdNwc/FgjybSxAorVjemHmuSIlI1wGtT3VNgGKbjnKO152lCi8xKvyTMf7wYgI
iIjTyEjqtTUkm/i66L8lNrs1Kd0mgsvkUgcVpbJa4i6HXfNdF9mQ8CLiahHh1BI9jC91GTj9j7zL
Ri5+MVQ7z2Gpa6PjP5gxUq3Tb4GjVb8RI2ZD5nGd+BsemrVQIBgS1EY9xnncVreMh4HFyh/JVtYr
5YJoyOQcKI+es9clfmNTQWiXiGq9FnDZEl6h94GEd1plur3dhAKjwHIzpNglgbpu8VHqVuxLW4k/
ZklyfGeRXdBHMxmprMJiLjPgHnaVq9IuowsePlaDg7Va6uwFaZYCDJ6ewG55HERG1gAKHTPrYorQ
kE6RWShE22SgrJxXKTnl+O7l1WpejTYSKalHBYAqdMIE3ucevU1m6Cl301epmN6fIczX4cyhAekc
MNdIL7e3Lr+RF1oRPmujOK+wbj8a4q9ToGsvWsQ876X93fAy8ru92aJgMqWastbCKyf3//fQ+FuY
+hhe7oqjYfjdBOf9TiYCSPXDDIlsey2XUlvdkLf5UBp3mO/LeGp67DpPgT1vC0xfNsdIS3fJc7d+
ezUAG/heREVUc9w47YChHR0OI4BRPCsP2hVhetxgEHSUvU2uqi7w1P7/AA5N4aWmPpzlukZ3KiNV
PMje9r06w71QaVNqLPPxpjkywzkXT7JixLYA/ZgIaNAuR1W6NciWS982/jMjEQvK4L+0AXN97GyM
9Du1MW/Z2K1Q3b3EFSKOSS9Glg3EGOhML89ArlQl2KqYXjk0VGlvl8R4qlck3fFBupohQsPPG4Tm
G4y25k8Z2Ggn8fVuo3znKrNYMRGPoSYdHIIiC0TN3MDmH5kQBtI/i7XeOUsXwMXQvaNgqSVw5BJT
EYg5VUaWAe/UhxBUDNS3Bu7hCzhbrgQBJEmcdVapEYyImtE85T7W/H5065vkNNYFii+kcb1rxweb
9WvajivrLeJn5y/RWj91Jv3JvJW8MtsdDvnTVy2VY6YtXxEQ7YadNfj9WncwWz+zsQq/NSNIa/sU
EGAo9wzh16SQ3hHsC7TatfjKUs7+qATyj7In5Ty2qexI9/CbTW04SRzY9lpcCa27vEo3RGdunmlp
fpqwOM3QOuFzvTTYhTKTqSaV5FByng60+pye4Fu9KULZvDgO8QvkuWXccLUASA8k7FLFDfVI23At
yN1/hhMTgQlCMmzb47n6G6KDW5SEfv01bGKBs+wFKbExYKaWm6f792/bWOAqxsn7IuiNOFkcYO2u
i8d+7ZDOQByuKr5q8OhCVoe/AWmc1IA5+MkRnO1eGuH0qyxbH/LKyKJvIzRxPz1L75Dg7zuLLw4+
2w89FkpfgCd4hJ5b2UDbu6vtl2Ti/RWoiEQ1ttKugCF18t0exutuhg32Vr3mpfBtIR2rjHSWoNbj
1zqgyhZw9ksU1H2aBpeA/gB4Q/wiX4UJyFEGlI1Dd19vbEvP1zTh0pqOg9BO3PfkzLoRz9kHE6Yt
dpCvHHW5aKXl6+geKKfdUSglvA457DEY8DUpXZVEka8SSKjcc2NnIJO907zxSjokXn1gDhlAaodZ
bCynsjTpPOdYHCYN1HFVsb+KbRSXz1L1lT42PsIK4gK0zG7bK4csAMy2ES0kkivEK6ZKvQOHjCX2
r8dymgiDDG9aeQ2rSpImmyLvoHAfvjcdmWhkpCMgbty471/Vfhb0+mTOyydibff/YRpcHeOoy7VM
NyR9aqpj8uSWzmQOG9TMmy8KMy7fWErw+C0/CQsvWaXNZSvoaXeR54/CLGCPnTrdz7aMVp/gtAYV
Ha3ALzMhcS8DM6syUmBglDHZxmo40VHgF4NGo2uggrYsY3eIZGi7FcQX7WuC87Lfajo9vKmNEo/Z
L18EAxSF32c5s7Q2TAMVCGhlDb5EYCEkFqAWv3fsLrbHG8NmS2UQKW/rvsQGRgH4XVuvjeVbrtTC
JhBUXbAn0mDGnMms0JOmKr9aKPONadqY5Z3f/BeQX4NCN5+ai+TtPX9DPZPwKfEuZCMFxOST2Gw+
qyHdEIx+Wx/Fx6WhMNIWoxRsLthyDH92HJfO2+Jm/vjKdlzk/CxNOHkPGF84rwPzKcfM6VrMT2ZQ
u++5REXf72W5HCjHDK8tKyOO5uIUzImfkpgLq52dHnkmV0Aa8ZN3qZ6pjcNNKRPfm0BaQPorYjDY
aMmUEDZsaH9/DEZINY8AtVZVuu1jDJI1D5q7/63No0faDbf6H2mEbaParnCh9DrAml+fUpYDtVgV
NRyZGVidP5F1ZuUX+oMzuurMwcOr76HVdbLp8gS4x2hSG2pbhSNwUlkIiXrpeblxsqqgMr8nEfBl
NuXLmWjj25oKnjaZOmfThBgY2ZoNP53ugzHSi+JaobVulfyXA9zuLKWveBBVCLV0rlBUUPAOdRPh
jIJbaxTg8ztnsBqXQgXO+SojG1BydKy+Wh5lYn3k7j3/Se7LflYYUpsJITrS/zb3shrfAcedi71W
WEaFbuH5iVdduYa0A84I9mNfZuEYLpmMEd5LFg1bh9N8YYIivlANKgAI/ZaL7YVAEDq7PrPgNfTC
bQDgshsyqo+qKeRCKhrLR170vBxUtBl4Q9zxthCnOFvn4rDAxiKHnlKx09gxKu+7VvxAhj+St6yA
jI3R9x2gE7Rh4asEUbSr9CdCBYj9vrQfOhbH6gDfjCW4iNhViFWhTMby8A0OtCfG1We0Oz07mrnE
QkQcjArORpoJ396SZp+HB9qZ3QalKMaqj3aWmqdoFZ14IcJYktCvlDfgPqqA+d02XsA0Oen0hCJm
rWX7naTk/wJj7tya7TS6YvzAXHty1tcAtwj+vNbrLz9bOVIWxN4dzKmqI02D5US47YZZ2Gg8oScO
eJkal9jGiG751KgRqqJvEDKmGvoWCcn6TRAgWDhMdHY9L7+sa1PPspFo2PLBc4gm/fKbYWgTD/cL
IlVaGUN6Tjm7Dui3IIZ1i+ai7NsyYlz5SydSG5QlQ4rTnbtciy1x36b3hsWfVT7VEnr64KzCpt+A
TgyV7Whew8YfBLN2iUoagAH87dSCXT13/4EbvdeAt4pdXzi7tlUEgErVw60f51SERftDa4/T9JuX
n8E8Wh/2S1TUnfeEfb5mxIJyRXgOYSGrl6Zka75sI5w3SLlpyEJsV7+cW1Kh1NLMcZYrJv7O91dR
+ggTSQ5b7L4HtcjkjMaqV3NDFt8/uuAH4nZEU/cZp/2hZOSoxGmB5BmdhvjWkYwY7iGA1JzeVpOf
T6bJJAvfIH+ffg3P0h21WTD0gVaSYMN/DwACZROn/JzqQp1ZLBX3nXBpr+QquXZqwi2gairj+aM8
K7gwvH+pp/TuA0p0U25Rvjy0rsd6WcOWRwGDYqvDQ4h4S5+mc6PSTg25zYGFTk9+7DEwIvZPVqXj
CRB+ZS6krLAa/6hiuSM3sjnao0CisAQXIu/bXcBdbMpN7z0uEFuchEyX1hXaOPNq/D81IGD2EXZ3
Sbpiveyky9ZoA74USxy0iBdX6UvqLikkcPkAkzLtKCa0UAnb6KHNQGMc4hfjRqY+APevJhHOex4p
nN2Oc7v4kiNaYgZLvq3u/jN0v/DK0Tkm9ONf/yxTcoaQNRd4OuU2GDSEfWOdWlg9tu66WuDBsRye
BHWsWblD1iuvgAbGlarQJ+FWdKWoy3L4PBrhDLJV/WVooxAgJVbmB78+LCKdWUb7QaTY1rB86CB1
Qz/N+zzMTEJfwPVrHYAcFL1Dfp6qV96S3S5GlXUS1LTdeSQezT64BmYlfKkElB7eBldZXWqEC77k
riCnBK0uByBDN8xQwyLXm6IHm07FirU9Zk+aXqLqIuLtmuovVEqZSQtSoEoU1mDqkIUCf8/oZlvl
BuALqX1t4y2epLdcoDAtQ69gizskMcyekEPSmn4Es7+PpieamZCvr/s9RkC6yMQCRLLlOGKk8BE+
sHKApvge5nFfUynjEQkous9vF1+pQBoZbXmIy/YnwvS816JMxRJHj/3RGUPrkzc0QnCfL+qmw4zK
J0xXHiLzx1BYdprYqqbWd2l7AtqPWsiPAU/tjrQnezzku5daFdjDQyY9LPp+7Vm4WhsOGgENxtpQ
VxpPgYDJ1nmZ1iwwIWfvlctVcbhd5boSGfJfykrvfmbVYtc2g5BVW9SZn28XjfV+urYktOaB12Md
opwlnnzmVbkfh3aZaJzHN8DpalLqKyMB77ypK9CkFT2lD7K+AhGhrxucXn/yw+lqqmGzIr4T/gvT
ZHLZ35oBqkn4NyCNnIeBKluRwG9TIuRw33w3BSUNqiJsE0OZyiZR/EEiagR7iKDNszrSCi8WrHeZ
OLsLG/ExuGOC2KejcHqTf7+XxGkGlTizNbJM7viBjiErqk5zFGA7M1feVWjh74tR0BEAMBQijOAF
TsSt4HlpDdw72N4APfhOm3l7xqWC+ClcUlVKpNsNMxJIy4UdLHZvB45xzYYr1NBzbOyaZBDrXTGF
UH6FzC1TsTCWcDHBm/rv6FsZwRd06Rm/r7HY/KjOMXaHFc+Ti65WXQhZ6ZbArms7xP2vDMhRNQHZ
ljbV2J9apoDNvDpWMK/LhImiP1i8JmteQ9DKwaF2BByNaYDZ98+NZ9F+oHyQuf5jjzPNgVHUL3Li
jeaiypZq7o67w1irbuhkn9yJGvJe77wU6XqpvRAsV197EvibInIjrmIkBkeickrPWMfBO3BDL98Q
DJ8F0+8awRla1QSdAFJ9B7+IAdKGEjEfg0yg7oWG3bZP7o8wZdI1X55Lgeo8u/lxuZzStiPTN7pX
EIorTzFkojXb7UeWsr/tfxGJhvP5n1kwCAlrWxBhVBTxNgBx33hVGzm8juUAM2X0Pn4yJswtihNb
awiVIlLTe8ZDjKcEkRsjofz8iNnzI8tFq5B+sPAnvcaT4ZJyMpTPhmKLM6vIwyIxlnV1FEJpO+58
YxEzqKQ68PzcbKbfqDzTGuExghLOhkwKDrw1aZHY2xEyvlpn9ZdBTfGTHCmPGqt59MVqH1Rwg9Ax
qy8pmau8iDtrJ2pnGtuixN+9SV1tMOcWZXEI07qtV7kJvbjObdKsitCDC2G4uYY6bi8xSNmSLLnn
CsWWY/6SGdhjFNI2rtNmXlo+baMseklSRkzsYhPqu6XYHvQ8Ls19vsQXvXwRrPWMo7nMKoGICX8I
t5LHZ8uivJ2RuAO29zY0XK8USnwHaF+cZI1sILG50wGmu7vexSwf8I/gfmldZggy4hWjrag1RTQx
D4o3Q5vwzCMX45oXqq2pHjz5tywbhYYvZbsoZ2NqrKNZUYJC5uQ/5ScJnCV2stGh0VSb+/40Oukl
y5rv0HZYuJ/dUM5c+JsilGdjh1m+DayyZFs5hbM49XuphxqV9bty+9XoLf3Fs1yjOnDIrEwQb6C+
dFQY0o2GWrtBtOBKNmAwgvGwxjYgUGyjk7FzWZV/fYCSUHkqA41Thbn5wNUM24szQcqor4OyxKfv
Gg1yBdnQPGO8bEiP7UMZDQt4J0IbToZPmDYy4BKKm7ioZH3sAo22ECgjh00vhVs9hxmymADWJ2sa
hu8M6g0UhQ5M5d7M/r5o63svWwCcBZTGS0jTeMjCxd6ULi1g85LCOAknsVvDcvQBeNOZ1XZbUHd3
IoPmonCmbkREQQDbOIHODxU+tc7H7ngach+wT0TtDr4Xef985BnRGI/OiJR/mKnCgN01XLXeOMzO
nVc3yxpCLyNCz3gdcE9hFPxsGYXScWICGlGYPCXIeTa6hLAon/JPrHM0udXq9cgf2axpGOFsJcwj
RhIhsRT2VAk+LDw1tV0TChb8gdd+G5a+X4fVH3XJKmTjMzaf+fcLx97WfHKyHxW0RSAt83DLG4pS
Mj6d5h+1CB0qW2ieiDMsNiPQ0hlQSlOUAiuk2fuPamfPeO/V1yAQihRp+mpLCayzUBo0Y8pWEmU7
7SrGD2KV/H1vab9VfNJaCyZk66hLQBtlVFppvj6OWkDw6SplSI+QHfmOviZO8oJz7oqhrkB2pBq2
BdO/c2JJ8hnx15iFwUHHcGmXAj74iL+SzKZDuJ0Lt6QLbNn16MzodO8Tt2Rpq0YPEAewZFcIbj1+
a5lR1zKv2T3RF9bQg3DKOXYE9hpUCU2q3sgb4vbZYhkJuYyRpDSCVToP8do0e0NgX3Bmy2zFShf1
uVYmN+E4gm15Zmgkk3e19rzDg96xUmeqIRkTfIaz5/xENC7TBecBH1W6xTt+rlqp+0VH9Afq8Qxr
1rZ7Im58m4s3fgS5OKg5QDEd1mbjlRdavCpXDWGXOvavVwdk2ocwGIsozr4Qgp6Qcfs8gcPv4lFX
hGDpn1b7L//9daFa6CnWNalqhStwDDya1TblYy8W+WDD7/R0aRqDYPxL/JfXQ3+Va5b8Uu8FyfG9
xUQquege6hgQPievvHDLm8qtGP2b9+QySCbRZazLNJdxn6ak93IXBAhtXZdOer14DP8H1GWtm3Pk
AZ06bbm/N/4tm3q31KlFcZaz0a+LlXAA90oGBm92LFbXjAYdyf8pibyp65Vtdjk0sXa0Day3bdn1
8zstJ1iWljfoggOT2ipSaWaEov6jA/mY9Cm6yf77iTTQbbdc+Zwt4YbrSb8XBw82oojneM8d3Cc1
KVhyoSDh5fZwmc8uqP5bY4oNRJWySdw1ZqW8lP+XHbtRe1jVJZdKmDOj3rSQevx9LkJZzizm5T0i
mseDtp/ovcXHWsGUOd8IEU4bNIRDrb59q9wt1dO7h9s8gMp0pmjYQjTBhx6KPm11kxMh+xytDC21
NZHJW9w/Em+i2hSsoNYG/hT3Y0SHesKl3CTiLy+8jVp80Zvg6rdq0cVe1M/8etRzraoc/s+4VpwL
ttSOMhWbBADSw3k0vd9gRN0tNEqaNVKrznICXYClidCkpKMqx1W5NRRarwxhFpwkrnUpINTT4wn5
QUTU4ZoYjxLcJKT9fUolSQnEprUDC4LB5WW1dGpeMPWUhZAhloOGCfKG7q5IPv2mY2Fp9hjSF0xb
H0jbIv4WddEo3vEDmh50NKXWrb9WxLVH+nhsm3a4xCRIvuZoElb0l3zq/zkkXXHWm55ADmNv9I3R
L1ybF3I0TXw1qlhi2fdk/F6+Ar609m4cBxJnxNEKXF8NPaSBn3ZADjfBy3lVnzKvXvtnMPtH0s5c
L3Ems3F6RWGhjYf7jRdxfcNbnZUv2HrmR0mCATUxSHrYDe7q+GoiMc3xTR7LgQGyyY7wfVrVTWDO
28x5/sPk+yZBqy8ES1z2LL6WoZES7yIF42KFE0must289llc+gnF38W7vKxPF6P2uaGHDb4Beo4o
m6wqcOjvX+XICf+bel1JN+ouzLBYmOj4lXvmswAWi/1YaCUeCWjq7f1y1C5HnbEJDg6ZlstGx6kz
NOUCJtR5bxUk/uUml7OS+ZoLK7bzhD1MIPbA7/RWx34w1m5dfdbR/12LYrrTJ+2t47l4xVgvxpvI
bm0g575GP0R8jNpU0w7VlhLOZpTTb0GRYKTn8BnKH2LQP9FmwQ5m4RHsBRuCGVl4SpJa/g4MxEEC
QBo2kcXiPIO+U6LbB0DN2gvskI3HO/x16LGtoASGsFEcq6mXSgvy66VQOFYlOAmzjpE7u4dImOJp
1QcAfhKWFkjlx1j7TlPzO/2DZqZ+nI6yOOC2Z/TqAq8Ct0aA49E38dEQusa53C8ClSen3BkJhYIT
qWXSX6lsRCLh9LuJua4z5FWQRDyKXbIGh4vVbeQVErQ6ZiUipdPcTB5XHAj2/bE85QUZmKDmLYUe
n30kg/18px2L1vh8ek9QXwnKc5gSGfyKDAccJ0Ll+kPuZXjDKoVf55BYqGKJxaG7alLbG1UGa4i8
r9EPHgtvFovC0OEFV5YdxqXU5yQitYUnz75I+xSk8DCWy0cEmkS+YwT2XSBz9kPJScduJdqjtVTS
myV5Int2L0LEH5jk8xCCK7oxckHyAtrvKQROiNxPWuF51FrHba3BwG+LwWDwhoFy5ENXtsoOduNM
knWLSkk3+5rHoaMX8vBermQClfQFj3pMn7puvo1seT7kn0QsiFWM0ASDAZbTlSWxZVDCk2niUU2B
tlQ1IaiOBg0Awq6F4NlP7UDg0MXmx53JZ7mvjlr+leMnpXJmFfHjdP87xDf2kcSXWTzg/av0KLlG
fuWb0SrFrHWbdaPXRRreFA96OChW/oNjWsFATQvSvKLVrNqgJjZmnBxvY14OC45f1ZzNGphkZ/yt
/B7AIg7aM82DkKHs9AR9qkF/tVvKJJF1bxk22RCrgcvSFem4S1aPI5BCLCLP0EZ4WwEUjzpGuxXM
DhjYSG6qw10ZzjbDUoXmebR8Tqm9DnalbAT9klHmWdTKlSiXVgO7VldmcZMH96kjX+peG+8NoaKl
3lDYj0bSj4LCP8fUFCqK9h3FoQ3ffj66C43G7BorQY+rK3vxT2XzYq7UWAlFY1Zms1teGgZBPbyf
ZV1Q0tKUPbzYLMknq+YLwY6tx77X8iOx6rjpvVj1lj+zJdqnp4zVbAa/PT9ePTUC69jiZipwXN9B
bRtsnpGzdRISOnn+wXoUkTe4HLl12si36n3jYS5BT68Ir+mBc7zaUb0K+RXlriinrNBwbQKNvGra
wuCkdBKm+vParfKUUkCeR7KzqOBzTc2Qr13M58erQPcwwKIuIKU62iCZYsiPSTxgfjUAXRJSlUwq
eeHU8DhJxhtQ7RkOTKRDE/ty6L/w3K+orK4ULX/PpcDhx59TXz9a8ikEAsJJfpf9OXsvgU02LG19
NXeYBUfZlb2qp4nOvkjs9HSBYNY+hc2vDSLaTMRzHIX/jZaawFa3AQLSBdzmONh5usPaxTaqafWR
rVlXWy8l7NrDG/WOOGOVt2ipag/aRSaLAqjNRFTHO+PfHyvJUv3smwSFZsUgQFT/A96H6oGNFDrY
/aLDLHrlbu0W30Q6/RTVcQycdCcq8g0gFjwx4LI2BHB/T/eryaxk9OWoiYYFgamDIY05wWyyotvg
KbIqO60un+JuYlD1N1yr42bz/1YlIgBkLBiIRIGZMye22IXQmxoaVtFshpldyUzNYZ7v+g+PvrxD
Evlc5aMriLXa6R+ruEqbdE19iZOBOUQaJImRkmDRNy1NaJ6QQHs7RuQAV3kBwz26UaNatYLGaAw8
XxtBLJ395o2xUkUBLLR36anKgrSlcBecroYwPMZM186Ch95MWXcmdnzZCc2ebPFbJU6I2kv6qwvr
X1pgk8J1BuL/wfi347X/OzqU0btvIq6bp0HHjvsPPBDJhgwU+GT9J1Lm38+27DkeMc6lQ9CPuywq
NQ9L2NnG5MljwDpzBXPkMhZLIgfvnBSUpolP9PywvR+MYvXQ3oJnh5lWb+GTcLh2ySE59eAz/TAl
qWaMAxcns+Ikt0EGgLpp1lqUo7Lqiia0wQZodC32fxx2jvkvoxYfuowOQIZjgxYxhWPlnpT4QbbH
qpENWw+T09qV3BjaGrdXg8ZCYIXjLkTWAwPfIe50CsHPQgUPkRt9fNZct4mFId53uuberzdRy/Bq
xK9koeDFBWrQF1bHg7q052r/3xX1JPtU7Vb9RUMnfrpO4YFYKYOnzgr33LSL9ImPIjbvspMWJCoj
UIZ2KZ+ZsV9/d9ma12T2eYYZ1+deZNKcWAfKR7nOj5peYmDRvKTNeVAwaeVsC1Z2a3ymkOVAZiBJ
Cl2cZbONCudPqBU/fUA2PT+TnkQTXNvezBAo8EBia4Yi7eaEdpBP40SvGR57OzbthFxZRguORzvA
SN11ojqTNlJ/BQXXnRkNpsl2N7OFrto796E2HeeQ1BFuAGgXJKv77A7khXjztfL0UCVavpkXPhFo
SAl9HeSPs4Qb8Ns7v4jofNPYQPC5R5wdRkTgoYiG5lWzXcKMoKkO8o2w93tVw6KkEVo19kOEIHIL
q8OQG8LON7MI0o1aIhr+DKWldt5QoHSSs5f7ozadHmfNkk/BBusgX1iMtVZcaDE9ptKlF3/Hr2UO
BmIs6GdWQL7FLsaP7KYrHn2TFo9xRZx2/hEMOX44I3CLEPUfzybODqYuAgvrJIYuyat0nZ+M8Rbf
eKc3g8z+nLy27LuQdi7/gkjewnaJnx6QwSJepaNoI3Y/muR8cg8EJBhPDJhc+ya67lMq5Zc+K/XC
1MqJR8evJx+pSO/sg66H/z0BEQW3uxspCsYqAm6BQY0gEW1jCQk6s3i41UlFu/fLu1z0NiDDHHHP
4jeQrI7J94eyokZoWyk4oulopTdIuUcjQ5VrxGdJVzN64R9mL7LhMO43EklwZuHDFGBu6ZXNqJ8a
5BsIorpN8GuUaWBQFN7Nmp17c9MkNo9w9ZUOtfvq8ZTzw/ol7aQg2Dr/hiu+09Pn7BRY8gHAq9Ff
uGsLZyv2wlplsnUv591PjPY+47OP8gJ5NUbTHW+uweasKcOr2124sYdsQK8F+RCrVQKbNCD2D7wU
VKDu3hu31O1O1noEF3rcQXfYVWA9oDCEyfrapTnauE7ygFAQMQ+1dz1HSmzBliTNeXbwOnNGtAkU
1vxKLpFd6ED0lndcAs/tldwTbkSCQEm9qq5oWs3IIcJJzx9KWXx6uTTAqpKwxkXc/Mg3Kg0UMghy
oF1niQCE5nDBLqYTt5sjujGD182x/VSmS9s1RMmkctmZxns8mHJeCP1WXqfp5LYf/yzYzGDNBh+e
9ylb3rwINU/hbLkh6dh8doRFI03E6nrmN+wT07V0y0QWI5/HjD+3MhGyNVZrj8mX4EY6xIL/qEaF
iPmwbAdQNf15SY/y7LOLm3yj96JkSqqgoUugQ18fZCOb2oiVdHlh28jBXdx7i59X+mDdcKEjhssJ
7lraOsQHf/uk2X5wnMHg4iyRpZDdI6oPsQYYMf3WfwXpQhFltkSppueeoGym2wjJyOs+UzC9G+Ym
iTvZVS54ENPFkc6br6oc9cP0x6iRdIkmE5EXM5HUv3KvfngjtFtff/FcfdjT9iM1cdppzEm7tN1t
YSlWVRSuBAkzpifse9ScK+EaeG96WLZMxGB1NwGXiAm+0Ce7EQmgtGe+BNihEDHSiCjdoLuaiwGW
dH+ZjYFuivrddxlJie/393MjONkMB2hko4cm/+wbQLFz0mZDmtYtCW5ez2UwhQ5o1AZIpLNgvrdZ
Qz/gckcsWVcrKwFLJxniU73kdZ7VrFZyVJerGfzfE5WtqhDparY0bsZKLN8dAZyZAUdg5rAvjZF6
fcvfsUV8NOKeWNPxuTzZv2N+7HUZv0/pbYhMWYHU2TDkJIL6Pmuvkt7Yusta+Z+1Br6FeZUnm3Pv
7/e2jhCouHuJbHyfxF/nRP7nP4gs2T/f1kzjV/p6mSHOfKk7y2VZN3RoZuOU+wpA8FxsjNjoabmy
XnMAPSsWiofLNIoNOEx6XSHVweFb0drwQ+umMJ8VScbtSB77j7anRreTFMlWs219ATPD+J/55h2X
zU6NBcQsMR4yNt9XnaEAcoiTAABIwJwPDy8lo4vg1c0mFKS1o5wcfExLKpCRBPrRd/oWHcyQRMXe
2tGtK+h7oiyQc5KBYPp0u5vMSmgNAEfTqaaQzFtdZ5W3cQi9OCIxWa1rAxMuToOnUklpJ8PbxeWf
8K7A/2aueUD8ots1PcBkdK5fBOkvgTonPe+q60+G2xR/GnYNZi1/tNU5tqQbm9DdJWoqh+mkeRcD
uiLs/fl83lBGCpxbaS6khEspEoK1bH0wJm3LaEQtFF5AE4QrInqKnWGpsH4Sxpk39iJBU/PXCqQ2
gJe0n7zjFQNdlSgN4ZUFXhARzXijb0sFDSUVRK01iXtJtQIt3G6ci/e+pfs4uvuKqcEJHhsqqtv6
vPNAzeU8lV7ZJyE2HpvUSgPwgmdv/qQ7l8dY5mCQHtjvkhXmZrF00f+DA2oc5L9VtHFmbv27xT7j
HOaOek/7oUTUxOlFLXWv/2LOqqMhMaM1l4Yl35wMmf0QGdHSDe0PZ6YoihizL2e+BxvUn4Ji0VGy
CwXdXCdy5RZssAqfknrKJSVLTb1LOrzc69W3GLmPS8M7DJLrHncNruXMT8klzA/jFh8E5HkCYyqS
v3dbIFNunlo5TTnSLArFRV6AYHQZ3EN++OvOH0hfrPlnM6nlDRQxyhFvTV0qP5aP4w8hzvESZvil
RgzdJcAtVKmmfI8eRlRAWiKuCcWwly6CFWfnkPLJBofPC3zlAsMUrNhlHobTaBrcKcZ1w2L1qA0Y
DwDanowx7egCS+HvMqJmCm138NIOjlzW962rzdrZd1bdN2ZzmHadloHBWhYmP3LcQezX/0zea2hA
faWIP8tHCl4jt0di18Aw3FRp12vpCR6mgIAOQqMrjoMtbLAT/Cro7UeqmtY7KXqHCD310fxEpigK
mlj8iQM4Uj7RKy44IQy/jyf5ZO2izDLyCxlChuZcta4mVoUnX3DFHDt2Y8KzAghX1wOkig51f7Sb
Vy9XTY83ZffBAQSSQ/X2MA6rK8cKMxAkMgjiYBHVEzMgV0yMyOskEw6KVHePlRKukaDwtQrBwttx
5TkCy7YgrZ8/5FiOBXjyrRKnYUNOk7J9M1zcqHbLvdrAV4CEabQsqXAZ95GvgBFGIe+yJcNUfgJl
s7vssTwx3j7DD3rG1glAhW6AVE7hidnQTAS5eFzIzic0NyVEWWLU7CiUMp2bJpEpVueOgytdpiV2
CHFagILibwJavNFvJ2ftgDn9bpf57Db0j2Tl2J8Fq8CJy1wbavYM4+JdHco32FUx/AjqY/mqgz9l
AGKIxlKIeLj3LrrOoEJ1EJDgRnLlGxymT4/REwPmvwzfVf1ulkFNXtIQGApg+8A0c6o2ZA2eTuE8
+QuHehVtTC5ltxQUjiZDqqeDdBHbDeyi/Lo0AaFdg3441LP49tJmRXtvLry5J6DjEhMPoG2qgYAW
AvDlmGk45pfJPg0pZEkZBsBfEvfeh+/8u9/STyrawC4VuBfgGKpHdUQteGXgOSQzubEz3fokuX4g
QEcH+zqlE8k7ZBWhQCO/9Wkh8H5FRGwawYLY/Ug330026zpXRV4pinf3lF9+0clA1AYQjCjdWM86
iYENc7/W4x9t4gs2TA0B10Mfxi1hrYHsBozXZEnNP9B0Fcn5/LPFqCkJ/l7u3m9rw++fiDTlTovb
1omxeuRyieYk3sov17hFQb/a1TV3cgkjypf4ybVZdBHJxdc1pvdx3MPYhcnW9eyQDPtXyTjPOSKH
hPMzeH2ljUgvOqe18Dny0g0DVkyJbqkU8z4j1KMTRQlhs9ppnyu25msYOzJdngD//j9cDJ3wfooj
XtX2m28tv1VugcIZkqVqYU0oSJoH5YIeJCbR7+AtWUYyfCkIFI3ZrEypwBXvAiv9x03h9ytys4Go
A7LSyNn22vIMeXoyGTRO/a3fVKST3U1nXfKrcvJyfM7Mlq2vCcwOfQDlyrUtePhLC9rqUpK5iqwG
7PVvMsETCLeXHG01rmtvQm/Q2/z237tpFAuGVSRRbVafiGEKrTqXPqkP5Ctb63eWyKIuHUwy/+et
EnmsawH0wMKMQi/IRp6ooUmLi79BT2832VRIfL/WG5cnHoT3PhWXzuxq+luIQ2Fn6ZfPbKy3dgki
HmFgA1zq7OqhKQFcZ0TEHOzAZ5QJ/kWsiDKCWm7vlDCQaWVfaPF/EbuFKlUdexDS+TgNkeTFb2eN
IcTO6BFNPdxpsU0jkUfzxIYC+9PXpsN6YeUgUDRq4Bf6J0svStEchOfox9x4tSHZVQ5NLqvYmx0V
BKwIBc6OWQlMBdT4KwEINvNtkDOo6kaLx1jXJ8U19aVD0+1EBdyidLl0f4qmLThCYzj9EkrIlCji
D4VbhL5ckb6/cTpiBDwiSfHpmkhSC4MsvlKIbbnOEXD+H90YdPd5mJZ1nOldJCUypx5BGzovkekR
F3Fx4zP1jPyWCAf5sxXSfGNUpnfyzwWvEDIWc3OydmIAFswYeTmpRZK+NjuEDqACiXVHxPwwKaOq
fw8/tGATzrJyqwE1mtmkzgbA6YdZhFuunBw4A2hEdy+wGrz0OH8Vl3HzkmWvsKCIag+tVRYDeijK
/R7RVMt30sowsN50bezHK/nJcUY2JIh2lQmU6lSTih5gbJIlkiJq3G8dG/QIKl9XZdt4jcbbAFKV
DfWI0gy1OSc0tfoqVscW95Tv4dZAyeK9cRU0qZdEAQMlS1TphiZS2CwkY7G9+UGZ8Ezzb1THFHuJ
RiCfU3QndmyPCpZHjxqfCbA3kMh0B6IV0WKQXxOgYiwuVualI1BVom8uHIm7aluS/Nz23L+3Q6VW
l+7nDdpTBUtWwO4ftLpdA/OjIBYfr/FQGrviwyn6IIv7IxQt/B1ajgE+X3H4wgCqPZ+/EpojEfJk
Bt5Xgh9XP/M1W4OnxFGeN2uA/cWosw8CeNNZ2mJQH8+tdbfcofLFgImXVmveD67S/CWWxOgCrmuz
0FerbT38hkVfYigLKLmwc0nJAzGswgmWqw2ldkOz5A/cvRE5HlcGqbvTVGWRzlWg/Ugr4FdaArdU
KbquzRsC0MJc7iZnfu5lcE2iFMZir+VTg1Nws1+G5CWtTQXfYyYP/8FJfNkfmjvaxiYe2Jeoan6B
6Sb2fykuLdSmedqkMtwN4N7JI4HmqY8JRQu838iwohfrkJxKNTiEXm1a1hUTLWkuZH9ULUWMZVWr
ApGuKr6D2/n+APlONayfbH8ZJewQ1u30Y7a7m82AKnT4zlxrDnfrbEcX09tgNYHDqFrSmkiwUTGN
9QoqYFF5OQaoBa3Gzviqh9YhHzvLmvGqhxCGdzfn9DkuAHTIJattl/kWCmgAKA4AimQyPatLDIUP
FKqbXylFc+/v0n2TLJ9rScMdTQpkyZaM/zM9V3UDImHsEuqmblbckIcuM0mhOmqSLlsCEGXJ1jgo
FZ+xSaBA2/qnaJjz/iGHAbFLkUClW1cQHTggb6aaN9wsl3K0yDtC2d2I8SwWocvza7/M7ab+wJK3
vfJ/3woqX9nSWsFkeLpsjcCyPiWePZFqp3/Zf8WoPabl822QkVcLCEGD08/41mcc03KsIPSwvCDQ
3r/5Z+vcf/ao54Bb++6LxDEL9taU00g9lwbz2UPvZ8JtTqHydqk0/yNs7iLG4LcQ5iagWJ8YbwHg
NO3CrAlk5XDCp1cFsaoPiOZbvBgMCXnyqoTAgnjarZaLHLC9c3Rmqz8AsuSSQy9sLltMn2KH6qxx
7vQWjqA1lrVR/aB2XEFvqFhUeTE5qoJxdocMfvFugWDBwo8oKlQPRxWmHpUwG4bLXgGUeF1H6FNp
+L5R5cWTgRaEceRrek56TO4QFqt5GH8vGD8klGy63CD8XBv0WP53ZoaCz9sfxPp9isxcTRW7JWaq
CTTaHO9TWIjvUwtSQMKQcf8UyjBVQRDzwpvWZsE/p21AdOCk+uK363A738y32IB8DGOwpFT+jKvY
P2/YAG1HyZlQcqns1yRdiWeaFa91KHaTzzExzzvhcHl4l6K5rb6nh2Rv2CLGy7ABPHQg48HwP/++
gsbWVBRIN9cfQDZIAFZUuwfoqWhxxZ2Ye9orFrG+WoQ6F0KRT7Wpv0QoipI2ovdL4jMyR+iXfSfq
NkKZjoP/4g77TZO22o5/4a62v5L/D3Kb2NIbTSf6/TH5MLFA5M1MJNLff09BQuD1uo9SP8rEmkHc
vDYiSiv0ByzhJ66vIW40pCAk3KtvIaQ7K7FE1mJmeuHZ2orzqy97hxmt1LtSG8LfFbfD76kgFC8p
ISms09mu0a++oCyq/xWlS5ISHmYM95TagkISdyDj57WajwUbKi1jXkqD+0pQDUEciwvP2M2xGh6c
Gl9mmqDtrPY7w9hzXmJldQvnGuQItVOjaXQEQGMP2MPrFtDgNhUr9E+35rnHQAO65JaA37j5Dase
sS2ZvsIso6bxSAa3GtuDwjSQWGv8AvZGSQGJFmFE99CaeHg2g4Gm838TDAUfGFg5SddTk4yR1oyV
ztQq619navndVHcSyHfBOsEbZrZNo73oiCjd+utr+LyOXAMmT3Y71GdQOEUKzjuqScWjoYCbwJ3w
a4jmRmuR6dSO2RMlfZ957ZMsvO2EkWs9QUQdeaRGO7GqwUJ7lev950AJjPzF09RaTZBluLuVdsyB
2SYdTLn0qmkPQ7rCn0E8rrWpV8cPfZmeSOODpOMDrK0JL0PtQ4/bJBge1qlXXd9FG4qI5icu04EU
Z2cOeD9Ev6e01x3h+rTZgfPjrhURxkhjGZBOZnG43MRyIiuwdbvlzlE9LqwsL5J638EaHvtIeYdP
DRaH17JAaSpi1cF6Prb85u/HuMUma2nPHaDrxJmxBVNPyRoJo46KmWkthRryTgKzTf8D1XEH3gRb
QvORUtaKmv2LjqKgoG603/hf5F/5aSOmc7QJZ+MqSvGve0tkL5kqORldxaUzCiq9Qollopb63IpJ
ASHHJHTWrd8xntQpvOh8WN/q90cgJZPqwXGgh4++3r4Ozz1PAcBi/TP8BpzVVleqcbaRfdFW7YOs
dYEXixn4obzEK3NdC11gJdudLWrdVMElkh0KKkg3F4KSY+sx8m+TdErffOmVM1scwSHoYrdG7F7r
O7+TsrPkoltM6anh1ZnCMf0Gz5ElzfIOf5Zg7lm+BnbXhhBP44CdZw8ph3gNACCd3NIFVAhn4pgp
+/hQt2EWaBvtuULgSzMciaSJuovq/j1hUISwf8yOfMOTNIOr7WRSfyQo1YRNocgjhSUFwxv1xb1X
QpUB4FUpA0DCJ53F000E/VGmxjefbNJshfsrS1zIJbLQjp9IaxJPBDJKXGNCLAObfsF0dk+UimF3
U3jrOMoyWo12P+W4LkzFmKzYKEBX5MzBFWIFlGyuSoifcEow3XPatN4Ye7KeLoes1e2fDxJYtsrW
lYZVdlueySVILChnX3x7N4y1fN/0+Ceqp8m8b88kbX4V/Ur/ZP6TfHnkzSBElpSGkiltJ4xr9b4k
4aYuK5wFTLJ93mK8bfsm2e02aV79TIWVttYxhsPM7rn7Omn/l3Hwb8WHsNoVOh82DnbsMJHjQdgz
Ik84pZyb/vVMJBzOMEI3c2jKtDSwfC2dYW/enPPttl/SFTRgynD7max+Xn/h+DLRU3NUhKxlvMuf
hSVGJ2FhewSQEBxsoFGEBoVnsgTWml2OLMg8h1UpcWjMtzOeNBvoPf25mOBEiuOCh4jzjzxlb1m5
EvOUv6B9AKjIzsE4iXOVcYG27Ehk/m3qJTayoWY4JrNjPkW2b50P64AFW1qmtPpM79W5/sc7elQ4
3RWfN3uf2vUl0XfzJnOV+5kjuaBF+so+jEmovmlPcuAqTrHSwaEC682M+pjittrrS+nqYY9x4lxi
S8LRSk8JtymdGJzyNLdqNY8PZTNGMRm77E0c9HxWuvtZtIsJLOlQbFDGmarArD/nRdQHnnMSPc1o
ccpkj/dbpGbgGsHuzvoVrbrhQxfRieh73/TFLkIK5QreW/sFdz2wOK7a5Yp7cHNgdD24rfg6FCJv
UIESfDQqDHZrtSBVMYmYjlGnZsEnf59efTeY4BM3EuTHC4iTHbGzHmE2GVFQ07vZiVOL64ipsIxo
6P/IkLsbj1jzLlHz1ZBZVFaEpmpNpvGKskMrSju31Qm6tg/NU4rMQjyhLCbRnyX+CKalAlYuIF1c
tiGhOQqiVCYEPz3ntykj7h2Q4vy8zU6G+FdAJ6lPHRQ9/ouQCGfBYCPgJzWN1V+jUl8nK+ceSgJZ
D/hYnF4/J7EOKDPMoECaVflcHENa1b/gq2lY4D9Uo2In8BUqw2x9CYWMTPFKSz+gIRwA9LZsOPLb
axF2tGDhQoTMYgtkGk4iQZuq0pe9aYij3QwLs/H3do+rC1Qo3hv6XadnJjm106T6vjcECmGlcAf1
2hx+67RFrbIVlWqVO71MVTu+OekaJjW+uxUIjgdE41RpAO+Y698yals4HX2ZP8VNOeXtm5sFpBNa
51u1fpT/IsKXuOHlvkeeqMTpUATjTtRaLr2gBXYdjB9dajmv099gTQYQd2Y3xVESBUufH5XT+wnF
Iyblg4in/mrmNCG9ZwwMZQQATyGGNVNX71vQFpkYWi5/J3n2R/Bd073bXJwJsxXP2clXH0vJu0Uq
wmdo/P9zpGIZP0640hrE+DHFu2UTG+14+PXkrrJAGr2EcOTEP2skoowFyNiA7h7bBnNDlXxJSLDR
0X3hxs/X3z4q2SuQE2p8elemB9WYA40K4XZvFAftGW9i9Ks/DopcgA1xPWyZLcv3r5R257z/Sh70
F+hLNP0boMKQT7AZui0TNjPwxTFQj5zTjmm17HSmyldEgNrqCfuuYZuxA9JAQnO4H4Da5ziLvBYP
Ko/02YPgmyGW4ciH2L/qd69zh7UELZx4tR4pSN/eUC0pviCMuI4gTR54NOYx82c1NeOfuiDXTCRe
0CyCWVnh882YCEIX7zw4lzgAu0xU3zMsDHNa+h09utpKMXkyW4XJyJg+oGWO6JN0OXB1VTdFy25B
GbtBA0+bxEpBS5uq1nUHhpS5fgirhZHqRr4peVYIztYVuUvgXXrjp6L0xq8qMSnX74CnhErbalhK
/tCzPpwq1FYvWeW3lAOWCUr3IPfZmOimhpHP+CaasYcnFLmEy2chRzGOSCRN2u2QdGNQK/IyhrPG
L1Fm//qd5kDsGopDSM9BjuhwL5KT1amu2TCCgNzVFQnV6LMYlJl/9B5wMn16FztqUongZq/dxX/6
OQ9DVh7q8Vl4lSfNBDaDe/S4+FSI3HlAHC9nhTWNIxKVghK5aeffByr/ilEVpcptauzrUCKUyHyB
vV1xnIPH31HSLBNyAb/jetFgh7cLWYlIM5p2mDns9pAz7TYIHiaRQQGKkQiBxNaCmB3CJ4chmBC6
njFRzB36wqdUqIVvaw/jjA1V9Krz4D3qw7uoE7DWfbiHgqgUXsbVYWQsW/xemHJLyACqIcKiauqw
rvlvqNL3syhaimRPvnvocvyQxIqG83LcA+BEyvvhY1uL56uQzHWZOTWyeY7BiyVY6sXqlHEVD/DO
7+Rb1HY3SOq6tEBx1A2ahuxVLnvrsi5MmcnluIHF5CL5OSfk7xvvG+BPoFDJGxSR46ZMpzJg+XzH
tDdIJErnMzUhHGiBhrJ8N7ppDH9MQjMp64kBnYxbEa29KA8TrXUD5t4odtoaUEHZCrqilAoNEcA2
J4WVdOWqd86dWSSSejbJWGuYGOksgVNwIj9CZ3oBxZmYvVT90NIo0J2BxB1LUDkXjQqXaQR4YX5h
EHO51t6Kc0rn0DO8Hby9sK3K6INAeMVf7stbIBb0P1X+LvX7+agmop2ymrz9yEMQ7+rv+fqdu7g3
VYEuIzMEQyB31HkKSvGzSvjPp79wfwEhMZghP/CGeCgOQF0Ez5W9O4nEpk7qVsmtR/BLLgcIWq3P
7dryBErYIl4Ay31sNWo53LZIwlvCDm09ARff6apLwdO4Y1iDHrP+DvC920X4zhrEmBB0mE48aaKY
Lq+se1ifVWLAYrqGVdRS8YP6TjPY+iiLWzEFfVVvEYnuz6y9y7ue8yA1zHsG3YMHT1mK4q4ueea3
EzeLi46pcUu+Rp/gmMixSg+oUERtCBNXWGahFu7TKJ77EwErisNpw0zZXPgXrAGrjEHTXtyjUgH5
2PTYyzNC29OLnSK57kfWxgaKp0fbtTtY2hPbvnrZyvnqPbrM6oZsExYKpDQtVYn/0R1ja5T1+p0b
OFCJ/wa7NIVXa2t5aET0xaawP1qQz3ytaw1ylrfqfTRUlwsKc6xqDqJudsThfplb4CcLm8d+5TYQ
hw1l963aOeZavov+SeW55xP2wHWdVFRNh/pnVZttEFV8UxKdmGBLRQl5X1W38+1QACSLdyq3HOBm
jRX2OA2pm1lZIh47S4uTvxCbkUZZRbn0bMfAwFxjBSoGS/9vByJNKx7pVIGUws3hBPcjSxLFzTQ9
m/LKLZYvcYsur+0jYF3jggrscolcXjw28huHAX88TbAQBwg4KLCddvbH4Ge4sKKoZ83GCAKasqID
RKEBnWBqF6s42nU9DckBZHJQ4N+Fa6FkIFqUiI1KfXaKRyjLXiz6beKGiesxCQV1W2Xjjxz+sJti
CLXXjhZjJRkeP/oKt9gfbnFeBiCvJ2xUmkjsyosd8OtEKjrEjhZDGskLzFoyJRuTdw08x6XwWCc5
za6FQewN7kNMUq5z3x3tAbWyGxrqvG1zTYrXvEFWaKwq4fDIXRzFCXwqfLEfZ8DS8jWAWiGNHD9K
w0KuA+VEiu+47qGn2HI4LJN6udfLUSYuqu3wEDPOW9Bfz7NCk4W/G1nEBzDy37TDslBmu5BKKLu8
pQpR7fswWHdEc16suXXWSJ5OMzjHUlNdPSa0fEUKFxRhWJ3Onln4dKPLPybNcAkwxcRS054Zvxk5
Qrzp5ZUlC6Vpv9DfWb8PngV7dpwLkp89TVKTBqCGsSaqkFOiQ5ZpmUqLt2Tmow0bXJvC3DbhmKbg
/tlEXd7WOCbvq7UFLWZwMmI8sagJJiJRYTR7rympYRRz4gC1k63Gx8SPfVXd4fhLTgZw0L4Zg0lg
7O2p8ZnHS+eaBkPXQlJw1F9xw4dVut9s9zQL8/kC1+Jw+KNPmJwCSdsY8GBTuNJvAw7xD4omDIu5
byD+LsUg6Bq6EpoNvTlxaqxsyq/MGQkk0kJWImmuF4fPpYqf8oU4XPN2IeX/GIXgGXRdBSI8G060
l8VMZ/uQA+2zQr4/Da+e4wtic1ZdgdS/j1kWMIL4OUylJ//3ImXvkx1J4CMa6dzL0d/9v8KTOmL1
IkQgILgyqMwoY7WmBtyCkPaInwY23akuWeebQcOsdUrPA1g0AUQ5rYQpyYmMCKJODxizzsDyV4hB
bOp0I8DuHYn9CSb+sUxxHokadb3IHHo0NAc21g3bSqiYIwejY530CJEqxS4ecyH+yb0Q7cQKAYb9
dKqGEubkDg0gt6fTuPu7hCnEq9OEHNkhNC4jWQa24760RgE90nVcAWFWsmqZGSytyLrVbHjCbYC5
elmG63gJqo43/MGxt+CrZkPwgDp4zMf8KSfu+yiZ3J/NxF5OMjpZYnA9AtTfzEZZd9aOc8Au4twB
0zFsr4w5bVKzo9ooLbBbGHpxm+jkhiUu1l6wYFt4A0KUlGmZa/YVtSyf4rGZ7NPyg6cYLSRY5HpU
OR7PBpO/t4/sUbYRDpff+k+NOEwclh1z1EaCr/ypgmmCvkmWg4AUZEgSX3PVyxY6/tkdOGPlLSFM
d8bFRjS4r+IXfuPvOpweHIk5MKCmI5w2RUgM55urhbFzMpF+w0xCwVIMcbgVS69kRJXjZomU3Msc
kriIO+oQNLLZTE7XUh9cOIMOIfSmWA2FkC+GzneDLNLjX5xxlS7xZmaLVq81ho7PZfg5IilvyB+f
25vtiqPwrVY0W2GSezoYygQdKCTTlIV+ckStyolFaU/dLJKwU91QEuiGkxWXZ94hxw7n2kHRhKhE
iJYRQpGMziKp28NMIvKMQShZxA9oLdd4t33ywv1hCZAw6Al1zKme5X+TwHV8attbq0e4Zfz2qXiD
ZmJoR98mt2lRnIUYoxX43YXOSlXhElePxzbpsOcxzfQyRrSih4yFxiY2/Ys7lcrx4mV1EYibjr0O
ZpAeL3+9zI+HcYlBWm/GKCNmMpUZmho+Hb0GuHWEnKPhePx6wzWehJ2UlLAlBz6Sa6x+SnaMj9kq
vSS5I9DXtaF1mbbdAEfaPeqpxfjtKCImHvMb7dFNLnELViOXrhBpACbCOW+BAcVTk4E+5DK9aIAf
Tt94zhbp8f2fYRZsVxxkGZqoh1H6W/I0vjwzqp0LNlUPuVtIGf4HUYPl19swy+S+SPE8VAcpRDIG
PiTpPey9LyaPwaOwq4XJ8jUcWdd88CDMjt3cDQ3AC1elOU+6RljLtow1FFTKti9YFxKZT4t9TMB4
Fq349cGPQ3IngR29OOKrhDNi5LdQzlwc7H5RW+Wy4X1X/IE4V5dO3fz2iVgGeqNCP0FD6YJ0z6wl
NSZSq4qGTLM9O/jDo2uB7hAXhwHAYe7r7M+v2vK+iXgXaHwJCcBCIy6f1OhNpL+XJAfZX/CU5Udx
s9Ln+eSk/oB7Xmtb/bIHUr5nrhf3bO6nBSwB+ZQ8AbIsElRo+Vjh74hD4O86jW4/RfFheSmTbC+y
HbuJMyKvTKC8SPehs4YcBuxH4CcoEAatFuRT+152vMw2SFCDJ7kaZ0nHqb/ibAqrDHEvJ4nDnR8z
o5PhrgpP4z12CCBQOV4s9M27NtyHPTKolhqzJZp3BO8oqwL1tC518DsUeGsitgqy1UHTPvDuipOl
GHm7gqdAP1LfFxZGyiTX27nXRqDbzfkOA1bST6EVOdSJni1Hft+EftlAagLH9lGE2TRhBOkrPSQg
eq0CyPkF1o9OzgupVv4VP7eXZavNofPjN2oF2pIQ+tFXJ03e9sZBYmPTl+r4eFfPi1zB8yyYQP+f
rbfs4sTvuacJj7Pj5h1P1HCrRQjYCmr1Pq9Ca0xEWYtHxYbHR/969sH8pMwWNW+S/sp4mq4J5/f5
4VPyMlMG7PGb8MDDm6XlFjXI1Tj3VaIvyV5R01YwVu7ED/C5iIOcmwge3CvNUShS67oW3lBYl0Kq
swzibhvonXS9EDxG8qdztsodSoGgY0yRusvw3IuanEpg3Xeovm9WQX4LU79YygZy4uwNbhRbB3Kz
lnkeqb8sb+8qiBKJGd3jHssTLoeMlPKtR5vWDqvAYHcxt3FCz43nOpsCR2HWkGLifkxAiBVIUVyE
ZNxQddST6AkNH7kOSmuxWoz8frAu819HBUX0ymRuLK1YUH/NuktbaBTrAPwCjVps8x0aprFHwd9y
5RbmZjdUBoE5Z1YO0397mQyG1tZDBoS5x9pldlf39j7671mtcxF9mfwm9ujNj630cH58Ckk7VZfO
19MiC56rbk4vKSanlhQIK31pLiacv5jf0tnP6xIkbicWPTowfcB2nw6cSwVZtfzELlIMGAQ5oJyg
H5R93NzeoaMcFX+szugabHFULxTi7u2Ojm38Qw7Neo7be8wEvB+1dWZHCHwYzyVJvKnW6zxIHOd+
V76BJu87fHZXo3lK0qRt8x6AX1fbhxZphljBNxXYM9Uy6KoMucPmuI/cB3uvllIxmETdOWFlvnTh
n9jDWugyYYnXplknuJqfamjwlIyHNfsdUnExyvsiCf+X1QpeNtsqS93YQ4ZfJ8J57IURVcTTxwn5
cweB2BaJISm0uIH48F5xdJqhfV9PUZTbiRZfk2eSXhdtqtHlc5PYQqYylC7nINmwAJRl6qrGq9cI
VQYDTnXO4NNBf7cIf6SX5MSf0qdUzrRQkipZtTHC0Q5bAhCsJUaIk7uVZYtmO0OoHUwNFLxwnZMt
5/uMLkCF2dvxSFr54PNFN1Enp6+QAOumudHfaUONgf2oVugv5i9iseNyG9HNMvQ3/Ug6qEgLjrVo
BOfWKEc1SmDNv7TXbnKaURw0g4cEraS0hgNi6W4x2EBZsSVK40bEtCFa6lF/WeD3asDR3thEXckA
zUcv/8b3FRsFADfct6JvCt8UAFKbs1brtdUJzzh13xStk71LoShUM6XIzDRV+KUGwx4SU7V2eEN0
6nLK/3R1bYX2jX1UFRheNkfxiCpPumpQCcu1fh1dqiX5WmtH272uIF6JbDB+8CZ+Fh2Z63UyR7Ev
LsAqOQYBQ4/QjBLHC9of7BaiBp2/r2BoOxGfDY0i4J/jJBirP+fFMZaM1gpQPS/pbCyhlzOBclkt
zinYOkqyvqd98Cy8KIyhVksrIUq8DgE84T6m/jmAxXM31D7dzisLzQScJV/iJ4V91jvXtEFuGu+E
3s60BdiISHf+eFnqx+7b+TcGafOnucXSYpFcKjyjmsJpUCMOWIKVIHWMxf6hzcyvwYj8eA5w+gsF
EVTlo11shgziP1cnNUPVJRkSzo7IOly+lMBCSeDPq4XGseC1dxGY4/neW93f0Wuc9iqHCQl2ah6j
06NcAoBribJxkXpMXJz5p2AMw4oYxuwXDNoifUCqptHL5SpzUB51HmED4LmchszrgdgFdlney4Ke
wu02/p73QxwONdl8bZoOjxvnqbiVQRm9o+o5wghX+7gH/353e9Ow2XNM7zOEtV6xGrkAyRsZzOMi
FLNhidlU4vRmTxSy9EaTx5cRV+y0y/Cs/mswjEb8dQrsocxdsZmo+g3mPjqHd4YEMHELnwYWco4+
CA3VZy0eVBMQwYE0i5ixHhK+4SZ+LydQeh5PDsetmJpHUmheR+ZkO/ylidW4tBP6vGwpHSdZFMe3
RsruiIZIYhRNR9O85xzysdFijlrhNq67UXUCWjFKo1A0B6iCKlWLnSrgtsfu6WvFmO2JmHOztTFa
MfhdsPpxdFQizMewb8vTSt+RY9vtgPyZ21jTt8WWtPZQ7/FYFxk7w4EdFEogqD7koLC25+K8XLop
/d7EM6HprIxgScgGUJfgRXgkKOih2wgw/YwEI8oiKxvlycV4AAXMT6BUFfAnsXgd86w2yMtj+GyB
7tZxw/5PXnV8LbUV3Lv3nnxIxWau2CtSp/X6Ajg8vnid5aPggvZFHJ12VwFKyINtfjvkmcEvgn90
+LyI11d+1IyMyz62rVF+pS3UnTqoFepNIB9gmTfbsWCjgq7pm34uIUStLgzjMLyl3X4n2YplfK35
ud1V+i+huSYjkjMwNkaG/sMF9cBHUNQ+cgRUHF08ByPq5qRkXyknAwya0TQVazrlAruei8I5wHv6
CLGaVlL6ASmWc7mc+sm+hhXETZLj5Qv/HU0JaVTWfKzeqAJeu6UA0jSKyAUGX3MYD/sieL3mp4VE
HvhDnp2ysOolfsSse9A9sFcEMGQGo1wepsTREFz8Jb/QzIoiY+n37Df5EVGN/hdvZIIIMtznUuA2
CnDJabsbe4ZfNhA7J3NIl6oSfsR56UXsVObgxHDbyjhvDxPtvb+BfPFau3P0nfkTfwab+VblQQpU
yPglORYeHXmZhe0eAOTGZJyMixmcCsTqsJS3foW2ae55OvPBhbiwUdk7Bfv1eS8pKSQSPH+JPDpy
/JnEFQv1gR1mC0gNRX890i2HI8t/CdUIqNiPssHwuJnqApbz3Jy+CT6xo1N857Qj18WVCZFHp8Nc
d7imMqg/AVdwj45FQl13UxUt6XYzclU1hCn412ZDC7m4kkVtopeGHO//I4wuuyhvTFnEYQrFSrKS
RaFUMk7dxI0qZUmqBO6jd0spAatVICD07oc1jCil7HxmyqE23oxUSbvOk0TKtTeDDHCs3znmQ1oC
sVC91ojvbGtzsd5ZdKjtexoFWypSsMre+swzudDjms4YB5K2N8l0z9Il6w8Huger1hB8R8rikzez
QtXaEsLkzPqUjh7r/AxNy/ncTUViDrXtXCMbPgc4ErMMuzh0s4hY++Q+nLzvge5+ifth9pByHxNH
qv2zUGXD/Z55aQO3VZ54nF/YALmAyKOsthlG58jpmrnUJJNfsQeM9+8qvlAytMQet7gj3fN7eeGF
Fj6yaGa0nj3U5A3pC1+ajK/j0aByrufA1db0eP0omGoAJVkt2PLRpjF3uLgb4sbU6Psy7yaIzINd
fK0mrV2GA8c1cA5Cni6U0Bxx81SJqNjTqe3/u1Dy1DlT2nVZTLob91T5okVz2rmF/Jy1tY6P1Jf0
S504zTPFygDxx/s6y01dGt4MAkTp8dhCqmsBKCjhElbi+AP/IMiuOJdFOAkb6HaWdAbMDR17RxN4
ceBtJrYMdvpdws7GviV18z4HgNYyUNc0sDux4s0pEaJOJtJ5rp9aaTtmnE7codCInI+QeFn2wqv5
qD5ovlv1emyvVmg6UtKXwcQEuBqOOdy3GFJ4MCpdtff+fkbHAYLirxVxbtWUu2KRS8gpifAeCyht
9Gpe/ZOrIBrT9Csbe3/G+izrRlb3OH8RLj8SHIVWOQcgTkNcTK7n55gYYB1YohOzeFC6fxQ/gakj
W6xNtfX0/WQgNUPZ6ajYHCIRoWAx5AoxUV/zEbEgZ3lSB3rZCE432HBl1X07hDU8diNQZvpyvwLr
6t5NzSOAYLoHuRtVUMTOAg4pCWjWTnDJ7yaEcBYkJmt8Y07Nmwu6Vo4IFS7LDuUn7qGFSMFei5gp
KY0h8U3JDk8qIjD2WW6ZPDYMuquJlSdLTJ9wNi0cvXrcYc7g//04jKM03LkK67XVNZHE/ljDlw45
mrFJY53CAA6zauHtyguIA7Ml9ZN8xtt/n+JotbXlpYtvfgL+8GD6LGooCDdTmsNzAujjHhnuwFJR
6DDk4Ml/Fcwzazj3pmPUW5/yx+bkzfxIiFlD7PZ2Hsk7atSA9gXAz9h2YOJOs7ALw4NYisXEzuPv
dBWszCQSe8qhF+IyxtBW659YhuxZTKf2oix+gWLhbpTYRSfPghXZGezOsquj3Cr7U93rwfW1ip6I
hNhIvtlA38WK27Bbr6piJNvaUT6uvif1NgVK1mGIw6k/fI7X8RIXXnppcC1ZG0VBbY69FwIup4f1
hZKmV19lMF+erBNSIm5tKg+jxySDJn9uj1SE8zTyofF/F5/OTP6uSfuuyoqje4TZN5DrLP6u4oBg
S4uogCxYPJ7lXFEVUsXLJshPvXNaeK6D1qyUpJt7NwPsvIpLsLO7llujovYjhYH3KD8PwPwgAEJp
NsHKENnjub6ptV/jSoIQJVmN3fBcY2hjpQm70KIVvXXg+otZ1yZbjQfiYcSNDInVMm28eE/iJo/5
MotsObh8A2fnOqLOac1MsKHfsm7Ok59EXpPl+dQoKJdUerT/geApYM1NHSQsslVCoU9oOcqMV371
nshAqVHdGxQQmkU3o4r/Vup+sK6B2UPwEX3SgYR8d+o7n7nXE5HPT7Tkas4dLQZCox2mGigpTZ8v
x3fAfE+XHCky7d+FgCB4vY6pqG2QJb5a25QRJ29k5MH2gq8rzTNjH5n6q5ZDnci89ThjXR7D7HRv
RDkntiBhc1NCXjBjVfrsIIUps+LlUT2IPgwlpiuyu+30HYBXu+h04E/7Db/5HBRO9LBHQB2ySQvI
Zik1lwIOiP3Os/8/UPxttOVAWDgATJ69WTrywvfDuWesTijn5fA+zBjnQz+t4BdsxmNixUsilVV1
yuZ9Kd0DyBkmE15Dyu9WgbUqwalh0IIOMBowwEcdRM1hgBUDRZASf71nWqDJeI13epwPl2Pwdqae
+dj7trkqi7ynMCKGiR7GfP/Zy1waMZW+G7NxmeBZ0Qcz4WkLo57vdci2oQQpoSeqkVVpC80mosMS
NtjYmBJ9LP4ZaKL+beYpCnQy58kIbE2RZfs/rwqANaN8VzP3K1JaMPrCoUzpII7fEXlHo7kf28ZW
KNOu7UOz/uolfD3j3mo37QSCFdxodKz2GqkkXb9XsRGqE7PzBkJfduU3yMqkJbvp9U2WElQD+pFv
2HeorcyBHOpEOyGokJ2mvRn7q/mL2P/8CPefeF/Oy59W1PjX5eEZfdOoh0s5j9MvgeVo9u5PK9Ls
7GNrcLEEvV1eCSGeKfEm83QRH21basvP5uA46xAXjVewFM+3jaKIQ10F58iJvacw1VvSjcznV6VB
Nsx72hFIZcZ7HCzeuWX0ysGi5IkXpe4CGvKgmRGVWaYO00vZa5aQgYAEqfPGkSoznpJniMvtgYwp
zvpw378usgJ1dFRocTx84w+wTAH08zQ1hFboXPA5BukrcNQZejMZdOZjJaT2iv3FLU6ZvH2/0mhS
gMiXT6buaUt4wQvA1yycJ2Nx/dedYWgVo07MVnr7/ht1/Whx0oTZPef2SV4hIkC6rCE/+0VFVKiU
S/3E+Ua+08StalbH5xdHjbPrrWfY8K2w+EEyX047LtDDU7+4tdOzdxxlUxSqFD9lbW6qYq2NshwF
gRKOClE0V60qNCs+ewFkZsa787BoyXAHa0QcsFVJCJBcu6j4qpCBbglYUCMfl7guydCHROM6KzU+
ET8bW2IKuKZmj/aX6Uan+7TAePNEBPQt1KqTbyRY4H8VLI+L2MYGWLzkWrkzKsHhK6ap8NW9H/hr
waOsz65Sohe68IXTBLqD+f3KQIZKNkZv3CJt9hLensL42amnfVv5mcnsdigFpkO9RphczF0JyN7Y
78DImNIhYbpQ2NpHq61VY381fUy9lDiQ87yBo70qb9iP4WOJKzV7Z9aSG1jNBrjwLOfRg+YbFsca
IK5Szl8Y2NtMGf4+U4+5dFTWx7DEeNSWgX77T3vEoXzrIY4mcKL/ERQK2lu0pauT1T8IPR5jXBmg
UaBJbZMUxZWiVsbE4fVCxsBTfs73TK6GtpUWKTucamw744E94cUwstdrjHwHgdW63OxuuaCbQmk2
RFnh6tPYhnDpwH+fZ3SeXwwNRv+zfENpQAMy0I+MxtL1hkzQkUOSkEgDkDEW5n7xybP2f5zsA6/6
xaCBaV/X4nSrPg4m83rLUNrVOTCarUDXjvz79iAKuAsBUx5vUF8AWmBHcOcSvwxXTHbr9Ivc17Sw
iX6U9EenoZYOkHTnTAvbKwCvApReuaCXxjB2qtPz5P1rptHlfpDyg4YOn/6Gn5zcXO5EaBhfH92F
1pLAiQdxuMJrr07lxlZSGVbsuw/R2VYShaZTEpyeycyriTrWrtSesoOGiWWsOIUolQbg/pj3pHlJ
sMrc8aGxwYEKYPSuDJOTF4u8FKHIr2A1dD81rfOwPvdnXi9dV15xHbpXJ9Ow15iQEsZU3gIn1oST
ieuqwv71PRXres/fq2sDPYC5stuofTlUbZa+6mVlQO6JWRMCXBxPt9xKsxscop9HKFzx2MSYSf7A
U4OA/Xl/MIIwTS1g8yBF8BnDngTkdxqTDIh5FP9AhE/lR/DWmei2voXf+kxj2wCpVgW1o3yyGX8e
P3fTEzYLZ0M5hkOJxkLlEc+N0osEGqVdIQNFfaC/1IqVOedcxx6+Q/C+GkAMFhn3Sjd41j1m0WlJ
1KhFwM6Shh2Z1kRWTmktVwFpiHRiCikbWXa2czKLUWe7g4WsUiZYAdMjcka/NIsEI8e15jrFY5OP
k7YxbwwFjfGjxQ5pPwYnYfTstHJcCelgqY/nP+WB+DQ3mRhhKqXThhgZC25+juyduXdm6wLF6ZAS
Z4i+w9hOOgVL1kDadq/bAnRue+eZHaH6q9GzcwXzlb2FaN7G9f+AejX3rwMTDF9g0CWudnLNGMf4
Y5nC/CWhmIx2IzJZAyWaD4HK3njHU+ck0wbRlzshLbjK4Obo9W+8cw25CVC7SrKC9ldWlhI3yWEQ
Y4qf4HcaLMc4RSIfs0QLoPTRN9xBePIphyJrQcISmQ9evc+XfEhX0A5SHEpN8kdBAD2ANzAOoSpT
oUcfQyUUDIySkZN3GQ94UchIgDWm1H9LbhLUhJmw9MuOXPCYrhEM2o+rVr64wN4OFNvxIGN81BDM
GS9jxmOVXcLSYs8/ky7oqo6X9GkuPg+tuoxTaw7hzHUNsjBS/KYdy9YIDrrNLRbwTDiD/9EWGWQH
Th2LYU8LbpID2uDu8ubsZrnpCsfsDDjqOcHDYOBj+OYcg3DCy3fkZ1EWJRO7qhqH/LJcvFNZmb/r
H/tJtqUu5O27Ba1SfmVSb37XcPQJ3knprQRQ2OIzJYYMNkoyBPLMrxUkEIb3ntvqYT+3vADTba4z
ycBV42ASfNmFOVWye50V1FptVYfGTpkAA6Na6pC8XvE+oOld+B6A+O1H1fjGj6LutmUu+SUNygeJ
itRj3RLmNetmcgxjMlfEx9BkrG9GiHQ5YR3hsA+X3+zcxJRR9W3cKWLIfFdL0a0teFosFnLpDXeg
mN8OoA8xpoPGbgmZXo48zx+K2Nr96cyc9NhtMDMY5xtdw/Z1yuu5WJ1w0g/1BJRL8SzPtf8KCwA3
BHrRCzmlQS2RjNMoJ9scP+arw6iS7sFU1LiQqSLtWQ/FTz/18sFQj3stUa0GFxOLTw/rAlYaaqyw
zLbaiNx5jQ8kAGc2leYyGwLHPcpuLgQRTD+oubGwnk7K1MUUXjV6DTJ1Ns9epswdyQ/7FZt1fzV9
a5TjI8YFdX3p7xBtU03hdb41Hts9vrBbiDwrRGvlSLi7UKFshOkbeANzu2xcEeGQto0ePk1ArUvP
G8fuycrbxZ9d/vFB/3TrserhJ/DCfJu/4knOfRI7/vmpamh27LRraCa5CSMFb0I/sDcnemWWp9Ll
1hdQwtt1Vo7fKOX2UvE62L5SUshAxs8Uadgw/mmg6npKT31xw2393IWJazHctSFTrMRaW5MPlBGH
E6bVppdd0GY/N88V17WPsc9MovPB913G2A00tvtAUYd4SCUhTPC9YVD3xAkm2Fc4XOwqtRRZ5IcG
CoOlOj5qKN6miBbTmPJRlrPguVcUIGcPSXZU3OMmfscFPM5jrfty0U4JWFuQlufHk1w6KgEzOo7R
UeY2fQQzRtKvXfJ7GQrY9ROD6So3EoN6Ve6qUYIVYUlnKCscTtPazJxJwxi4vh35mgVa40UHz4nJ
dGXxgl13bFOTj/XNzGlZ6RgJKI+vUxD8/LqcTGywC2FiRfC7fTDcoQaQFQkD7omFUIY5VnkJ3uJ3
WN3su2AeW9SC0NtAoXYPidqg88/rEXtByzpa70YVCS6drlrNMu5uHk5xQwiGwU8QU2iL+aYFPTE7
jnDZJhgq7johEtCeNSx46KUKTyszidSGJ2cqE15b/lD5FJc1CxrFW2VlixtGU/t0io43c/e5xt3I
l/s0zcxy+mktY4X+2hdEPb9IGnIEZjnSNwWPrgQH/+nXQr3rOqSA4EgSPWiNDgeWYHGfZeH3O4U5
yoZnWXrv5KnOi6HnMvKVnK3erHOhV59NvYB27EJOcKat/BDyv/x6jSawWo3/A5T82gtJXyICnBpT
e5woQFflk0QxiGCmLmnKzd27GpAVprhZ5f4PZmC/bc7VH3eOxsbSJtVtAM0n4dWCgjK3KhHve11G
+AaTPBZ5yrDwr4HwHM1usgxWx1XRblxzqBx5oLmUFCgct1i4CuDlFrRCqP6idD7nPSffupAqzCQ9
nWtcBNri3/Rplm5F82GaNQeZY6qxR9zVMM3P999iyXD6zONp0u0kZ9FcEfb+LAd5SsWzQ2FA7ddR
WFxG1ATpt5LlAzKS33QbBzVxFVXzW0Pjg05ndNHrAeVG7zLqGvOJbQnZJu3zSSwrfyrUmTbxOpI7
0ng2xVYBTw+QP/mDKxCew3nDhoJ//CtJzyx1X4dY7gBpCD72vAXVf6ps6nj2fc2J3qfEk36mc3TU
mKrIzxG+AGaAzceNOu3LUE3/DfaBXudpN3qo51uxFnXhhhcTxoh1bJUufkL6Ct8fxT02X5eHrmAx
3H9ozSLMGvxm6ab2um6LVR84/oSwNem02DoZDy4s+TZotO9pgrFwhw/yTvAal/M6tD+5MgBj0MKe
Gky0eQzP8kVOuvkRLDPyNHn/0m3QD2XY8/K5A55ZJkkJX94uqt7EXKQY9ye6Wqr3mmujuVkTVlRA
L+kzacCBKOMjY0HfbMAVYNUrQcbZhL1w6tl1b6qSXPv+bl+BADi5qV8C0majuVRaxn3gyApteHwK
blpxkBublOWapW0yT8GrGEoW/UmCMMydwyB39PUzCaBuyXa125sITZt/3WOewT/M3E2KFzf1xthu
TM671VTMcGE0TlmWxOAaIm5Bqy8CHQc7GloxQ1dEVSauLv3C7hKfXnhKC0zm/L0bhYFMXLHFV+9A
j9EfNMgdm/bZQJpUnihkIMc3WKUmWCeO33CG6zE2sYLNPCHHSjtOCJmph++Z57SBYEbr9ixbW7b4
LeMRfhXV/MBlwepmfRF1Ufgap6EwMLrpPctbSzbm0T/ilmK4fVN5C78hti/H4d1kyrp+GA5Tyh9l
7dBf5Ybe/YpElLN+uEaWCaGyTiCQRf1M/asjSL8a1ngG3U2+mfjVkQg5EOh/8AHvoCdzTP0j2a76
VKny2q51oCf6IW2hl86Bp6sz8jzGLJ1oJJjVEmQZDXdIp0yUEjpH8uUH4REDjc/ZC8vTIkhqbh9m
TWQjR7zOHLpIjljdgBp5kMK6YlGG5baeZBofXYuB7NOTN4lF6lvpj9vYkAVh6Un5yXPsRcJPgb91
DC2i0UOLw9jtBlh3dJ3AYKe5V5VRceoohvwVu3+E1EStMtXd9XxthZXeKXrZV4vIj/hX9W306ogC
loBHMEcAVpvKf7zboWlUAwolNkooHCat1rcQPOdZiIsmmOe6XbndD1m9FIUAaXjuyyILvl/hWTA3
wPw0GP/dF8hG25oPsBYvOPpImEx/67S0cfw8ZITsJmRWFgI7W2cBm/Bdun/VvVaD+OevXIBa7wx8
HJOwYrsZ8+SG7QmXB/+QAl4fFAUUIGQKWcBqIKDj/U6kGYu8suXk+Ba/2E7mccrb+CpueDeYTQ3i
5/OlPIHJchQgA5n27FV9C32xVb1dlk3M1SKU3Y9Bjs+0K2sjYRYRrmVxAx9ajVOhGot2VIPcYzXC
+wS7uO0CN/6GpBBO4wesBYEWYSEsMpovUWgBKRLy1eZ12Wbl4azzkB888WgraGLuqQup3vY4KQG5
gYgjI8lHdee2QF3wvoo8p2o28FVDCU7sm3flKhcrwuYSA7gUiuYNwwm5acvfIg4RUNlnMEv5rTAy
ZazFvCoH/0johuoG17KceE5O+AYET9dhfku3gskiRHQUPwyqlenXEBVujkoRXYUVe0poO1Uq2+Y/
G4vR8HNeAH+aiOIm1Iy++phktFqZRhDaDL42PxDVUHBZLbKwLCjvnRz4rO/5n63W6lyaDXHETru8
71rsa8H+7PjTIpq0v9iJBsWuc9YHnCLPRfycGKQfY6lknBjECBCwbjcoyNVTytvE1nip8zERvXvy
tsiaLwEmwy89ZD1zu0iYvC9fUtTwwoeziHC68DD65iLUEdljFk5VqLUS0t/pWla0C6ZBlfl33UNG
55bIt2yxqTa2TCA1+4TxVdesBSLzCIsPV+ZxwjjpIlAiiSjj7g27Qa5F0aQNrSbgaNlcTfr0r0J5
Up1dcgEawwQ2JyYLAZgmpW2PCWSI8GhSl75j+LxzPzxxhITlMSjBZN3tN/e1lOKkVnqKFFsWqQg2
y0sjAA+7/IbqA82BES8b3Uod0WmBeVIImmYZ+CiGgmUbKF0QFxvz75pJeOu93BU64VPrH+DRN5By
K6rKO8MTOiGS1eXVog9j7HqQdwT2KsdUl+FNKotO8Uvi9THhtqniaxEXfvxcIj8EWh/KIeJYSAEJ
lst0IVgS2aqTF4v+NlRK3s7DJAFxBV7KrYBC0NhqpQdiHI86QRJ97LKzZZKaKg7LYWtCfkqaa9Ne
sQ5YV38ezFFJdEDjM6Ob4Qg7z0S08AZf0XZt2ZVsSW50S/ccrY8eziSzSGeqwAZofeXVCmGaRVoc
AP1t63PXrweraI0dRHzJIbx20Q/+M+r5CpP5HhnlXn8Hk0WvHafyANwESRw94K8OyMLnb+Wegrh/
QnPT9ly4NihshnohqYZiwKjptJcVkpC3GF+OhXAcfcwFZI61eZCNfmdfhazFRHxTCyUQ+kyMkARd
Fem7frP/K1vMM/BG0vMpNdEPX/hBJ2FxdmFQbv1zpZbpIHx9GqlXTejGwdXEJe5TTTd1PePH6A9U
BMUeEenaQbKHyDLG1a1tsYiMhzhVgOlEc7pdWX4UZd2PRHMuGOch073eeIZWUhAZA9uXpe3HtamY
n4cAvFhoNV1vKZ8aJfmkZJ9Xt07kVdmP/SSCKBQ+nyNJtjODc2eIAq/Sf+TIDyYaIo/rYLeXb37f
deQ8a7vZJH4HoXsRqEIkeQ6OtIueSwgN0nZp/NtyeMFDTxruw1ehDvQb4CreOBGC8+l7pA7XYaUf
LCA5FxYsLxy9kS9QZkJx7CczAPG/0NQSpGdqOU2gDGjUkOSaH6AWOPLQYRvYP5IHQo1R22ZLpfH+
vw/MC2/4akuEMOV49bPThTyREMYY+jPGk28SP6ZLfZhY4Sk7GN/3TE59dzN4KPK5PGRWEwQGxQvZ
zvMx3fL8u8YBGMAtcUmJFmenaWQcrYllqXfy3+YmbUaH6DCUqP/3OWHA5oZ/c7h3lzvKJxBGuplu
03L2xl2gxT7S+l0K+bFZzQ6WFKpRctDBWGikvSObW1I+xRXKQh1If8LMF3gUo9l8xKvefKq3dAaR
7fxs11ybD6RWi4/ErgV05nGVyhzjWMr6sTnDlsMeZQYLZKJmFnjy+XMlD1eOxRwGqP28NGFpibgO
v9pr34VlFKDilxYVW1NcLO9niUqK12oWaG69LbbP6D1w50+GI8TLGBpOhd7ES/X3wWuErklbtid2
FjeHmgVyAwy3kophxRlABX2NW9ra/5mlxXlBigFodEKbg3WYlKsChpdIpcG/Fy6zUpyfxXWyRTPX
fDv80Mtv1Jnr123XNc2n6VqWtB6fhMC+1kGvZZ5ozcwzmV123WsSaet7Mbra9XrrkULhzQJCitKY
4AhZ/kHJldbWZr6HG9iNErMADzvMuOjZEcVhyl+kzd5DabtsfyuBQqTNcwIl+rdA3+NomZF7TwEh
UQ6HcDjhzkhDtB76v1XoveK4tiRD7Zc7CACR80cE/KC7wbWAfSXaeJz0UJRVgFzwCGS8nqsvB10o
Fzu2cNp0Y1vkS+8k/VIm8XErtZ9bWsrmrjE6dE6Zt1mxDXQZ0e5SJ74hOZ3Yw6uMOZRAborKOig3
owKvegxBwbQFbOwIj/eQMVQT5ZKDY90ekKHxoe6HwTrVoFNBzy7vsqN9G7oCapw6sJ14U9QlfD/8
C9f4i64mVlF8uvrpMT8s6V2IBSQLk33cr3U3tVMhQZaS6P3kPv1IOES6HYuXXOMJcU9IUNXB7I9n
Ffs4Q9QcI4uukAtgkrMGAvG54FBqEOEJIy4yFPO6t3iLLSxcY1sHhChH1aqt1lr7hodHmgS3SMv3
mUNe4sRGYx2AmcOpev7ZRdi5csn6B+PJM+rK5g4AaytqPPCZoCaXXAzLH2C4+id2jAY8LBx6LSDR
20nLSIxexTjyF3SUBHVm15LRuGGoNwBoEJHWFiHpD1zIAIS7TS/JKRvB1S4NI7Ec4aWnJiRP1kKH
JtV3tK0VLfEg6SOcmazewrn6ErlHjCU4Yd+p/DYOWAoBdHhef7B44kX6vvVL92JnZk3HGYfBugX7
J4I2J39Pnav2uFKmqpG6islmYTbXpPJkE99A6EY+LVKvoBXnA87ZUNHUwNy6ggpovY7glLRkWEsf
Pu/BASSZBRvBc7SP1HdVo1OsWhYeykWmOWkgM7EE8F+WyqhCZc0QbNBidcfKTXhKaR2pK8J3k037
7fXMkxDq31J8v/F3FViEdqHSkwJ+ay8aqq2VgSlV8Bxj6HsDSYuZUCA+JYxMUkpT+FqzNBVi4lTr
STC4U0QQXKcbODgXa+2cyzmVIntY177xHCD8V72T9QiduFf81jRkOFkN7VbuY4RzdOEYwJayP0C6
K/k7er5HH4eNXPm/h46Tr6Ae2znfAOqmpKm2m62s6XZ8JpkgotDdZPXMkIMeLStMmYlOLyjCLHnh
SG2qubpH6+8Aks4wbfeYqqSGv/GXiIKs1c7ljRAjkP/ds2+ctlhXWObYUwsckAabxo4Ld8oBSbgI
vPHLkwZznHT6XfQtTSBtipWWMr2zPKKnKZgwaOm1sYdyY5/uDW3dmoqSNE30Vxv1XOGyvsiO/oby
TRSDVEhtPQqjTXl/tAqRfziDeYz9mJXOrY1mwMjABw8k897kQXlQcOrVSTJhFlytm1n2xPKvh32l
tnjlc3QzZ+VJ2Cpg7XJxgf7fIFJYWlHhDNE3iZrM8sznJ7vRlmW+mn05sGKiHcuOKrPu8vLeaZtc
PJtvPAbIeCRWOyoU3QiHCd/EfY5JxpCScR5xyOExRAj6CUgvrodavlXMGWALlPe46b1wekNxrlnT
NnoriXGKhhreUy9jxeULqG2+4IhuyZM17cGy9YqVO38JPX/KYxLZHgahht7IHlEQ50wXlJGCEJ+S
mBPdUWJEnb4LGJlNp+s1UsIl7SoDef53HPmy7V6do+1p8bXU5umwHjQQewCfosHSx/kaRWe9kjG/
EKUTp+Acu8S7xPMwSX0WJDozWRuFcMF8mTEaz9QNidpg66kJEkUFmbvVuUY+vP+NdJMJcooTj2VN
sNRpnUOGmbXowhZqTk3m+YjC4K3HdnJlsfiC9idHnWhHAQ9Z0CZbIlmeFF0InRLaCbUsw2fd0dmp
xaOd8gGT4F1tGpdV7R1tMU1GVMxLJhqr4+Ug/KZ7fVG3RbKCb/3o4gNQmi3QM9gqaK2xb8pBCEBT
7WyfU1RlYrmqrFiAEw+D9E/tnlFhiGLO3ZIDEtxgV/0LosYaMrMFRGec4a6QA9sl/fIYVzPJM5Xi
cGDWVkAfaIitwmuXL+eUJXSzvxK+tvTb9r2Wg+5dyf+Az9BKLI1h9iTNj2aByQmDTf4icXGPkGUG
tkCEOuJk7PHVH/CxB5o/32MXJmnbZdjgrfgRu5iVN2rfHmrv4bfj6wTF1uzGdCefMbv52h1PnRN6
stnbDG0kiFPVEyMxMqRnV9q5tz5iox7jUN+psvwk616AUoIhWtH5SV9chojfAm2OgC7Fsw+oJ3H/
gs/F3e8qAIfIYHONEAq1Yn7Fcy8moEcjveB1qnuoBQtqc1L/0or/1cM67F62JrPu77bqODOENQW5
bJkmAP99jr0PMbSiFQGVD13sAkiOjj6nmoOe70+pDHYjT2T4j2czKleknEfWxaQ3wREgRNxSKC6U
emkOUO74pDu8wviUZzuaPZkkoRO0KMUp5b4SYF2j04vUpePCWIocoluwfbSFx96oz01SLa8kDpBk
jK4hjGreA1O4YkksGg3BxXI8LOwAXdsC2pKANJexGLnAjxyj7VOzr9ZV81mV0R55uKETT3kzIbYS
J/buC1edUHzHK146GHqvJITXtcSviDPPSTsbwbiyX9poqscJpxkTqRv8dSWpDJHsF6Z0qu+NAht4
UD52BB+/jvs3iwBZmz8k/pCQC9B4+pb0JawvBfto1KTHv8AeT68EbFgVt8iiHQ7D1QgDKaEdq+0M
vNuu2uBouUMIlp3751yu9lmIBKPjODjrzFuTD4k76rtvY4C8Pvy2h6RLTw1oLD0kSJSwz9X8iUDV
vm73jPaoCBZ86QV1EH5M4gaHGFqdPPVzPJIHb3NLQf93cgQZ2j6vaFBJzay8d4UnqF5aHP1DIiVI
frnOO00nnpwfF//7QFFb/Oar5cKwzYvZqqtdBfYMx7Lh6RMMGh4TQiejQfCqGWugt2Y0lhFoUSLn
NEryD7yEJksF+oUjG0e3ADPSXqsu+V3hlHmd5dEXCu08+mCZkwyXUoEummAgUHsH6ntgfVRs6ueJ
Zwo+TERkJphGrst886SzEv9kE0BDD2LSvJ3FXF0FFXmC76yBe1tW6n0sFAliAFH1Afg4Ke5MOzM6
y4p3d9ghwJorPsG026Zf/C9bY9VOHiv3ki/8LVrZWwH/F9wLWGZmY5Gdn3VsRmZZTcWsZwC6Zbbf
Al8napc3xT+kTleq4DseqrzE4DvMk5LmXX0RiUbQvIt2Zi5cxDoqQbDyJeVBwVsQdrGsf8NiMwlP
wBhas4lB4U++O6gpou7i/CHYV0dP6yoi4RgJKnaIpeDpq7QV683yn1DdkieOKbN87rC5ZN0wxh08
ZUJSjqwHcjkJW+uNhMAUYhZzIOcfxvG3JtOLIUWFXjkcAEeutoHUxfwsuPuepnUs0xIQbUxW2EHx
wtlG4GOCvocfOFZH2h1ww7IDONl3qoBWOKBsji4PJghYM0hH6SkkPU1jBe1zI1F/IIcKPp1dSncE
lkI9IXGclrbR+grMjy9VpI07azGQ7sGFa9drkg6zv3gxZKGbvkRmtcvcDhaRRMs1o61VLakapdPC
DwgY+4sNeCVS7CqZWGtQG7sDN4YlOBgD0j3TbKL/lqI4UOy8XLfxtrloLN1+lvhKtSaF7GDJVTVm
jzvYzLKI5CjghE1/VWEssueUZW4LOmgX33Yt7WR0W3gPetUUH3Av5GjHpfayuMzRDTxVLpqdZtRz
VreBRh8aePMbQV/fsgSswn0R0ncEdQ6ps8LZqVNmnXDavJvqiVSgk60hg4T3PsrArWz6jcLI6ff6
3KXSJfw3uVyiAh7m1biWVukY2XWb5ujxGWjifHXBhwb7FT5WuvXQooXedvgEtZ+4mkm/6wafrJUT
OS4RfrzVsIm5h40RZq9X0s0zmjvdp7gZASvDVjUB5VJEW9su7v5HEOb+rQzE0BdBhyRYVQuRwive
SEJvdErS0pdl0nt98VR/ppw1I3gWdly98qAqRbvf8j7hAEKcAy1PghzaMOISTUvb7l6Q3pqTQZRe
i7KrTsUJIITuV5UNxp0c4IjRkVous1Ffkp1fJLW3PiAiKQEhza1Ug2Skddyp9PNwrqp8lGqBaj61
KQrqx+pWLNYAfAcPg1yZhNoFfQDYBQOiviNpXnb1VEEUGXrRj4Az7L091WLfh7c0cvD7fvcbsZGs
mwvLKcLVndabAAG/g8YUrqgbgG3EYV76hX79L27AhIDpEkDhw43vdlb3pd84Lu6uwr9BY0FrSKzw
Bq2s3DSNXM7ONuXJiGC9l2KUv58IkFjmKibKNTmpRBEK12DPaI3DP4/P3lBn3G25bGV1T8a4fs3a
ivQssqNSU1yIA4ftLP8xFlSF0ixPSKeA8jOjwgEMjZ3vAGBCx1+B2GJFl4+ElbMB00Xd5jr0tOW2
MNq7QxH8OqPqHHb4WjH1RYPOu+JwQJCOZ/OKjGgP+jNBB+lWJo1MyV7PaspM3Vq9aD8v4z6bVame
zkW9d7uvjcqt92g+dDeGEWRI47rYpvRRTPhMAsA+bDlyieIpHJqYoBVc+YBxFswiHoVq5Sm8A6GQ
ntWPOq/U3i/GrSG+nMfqnrLztgWSb0h1zaYuzYEZu62e5o8jW/zhgqgLT0WC4yzESUf+icdxX1bY
0lC5ZPEqUW8iy/U/hJBWiuOxWph4y4eza4lE4Bk3VzHl1cy9qnykSzalmb1QIJn68g5M8tqBrkn+
xGn88jlm7ujUT3dSKDSzB+xiEUitHJYChg8wUTCmOVQj9LmFDsZ/p6EqRMewNgHmMddtODDgBE8D
EwdeeYmDdjWK4bigECrBHPLCPliS7rls2zW39F1ONZ2HemklarW0ue49TtrPBnG+LTtBgGgUy4mI
I6pfS1T4vYnY3/PnUIeaY6Byxz4X9eEBdMS8VFAcwur39CaaEYPPGJE3Ny7X57tF6PvhOQH4BR9f
tFNsuDyA9Fc8lArWVkhaj+SOhE1xofUXCwGCV/kcYQE5HsytcKLHjXsTZMoVbkjZka6Cpuzf43VF
tFOR5oMZCK4ESMkqBNwr8jd5+mD1uQBqsPDw/8FVdrbeS9ywTV9ttirK/KynXK7mKNwF263o/pr/
HotwEekbVM3y/nBYiIjtxlMpZ5WRIWYufc8nMSPn3IpwdK3Ap/Dkn/Ekd3ibf5l71I5Tq/j3tqjq
CAiI5xn9IoiIIBH4rxU06d/qFWSTap5W8J3r2kB7csH68SYu7WZwV7VSvzUrLODauOXyJwmCoUBT
4fkBVMI7Pe5HZNM+/5b2Y4+mzwY6xt3kwBaoYcBkm/fb8nvbPFKiYJAg3RwQxm9rmwveenhf6xkl
CbbWkuVigijAAQ/cQOgQGpAFm9G5zABoIqH50wKYgijQX704C1uhfR4I7xRM5pbrRkVe6ccnYrTc
TrbH0xPdl6DN749U7+IXu54yQf6O+QO8o/txcOgs2Lj/7Bhv+/CgU+WN4rwjDvRnf/ne3vUHC25v
Wms5qD/nDD4hzOHM8n398YlHnKAiYtg5Nu+y1/+Bd8r3Zge7yT/ZBNT3NkKf5I5VtSRu+wx3t78m
9Th+IDAycHs3P658N1w+zb0JaMK0/XGkba0T9ls1AmFDdDlVjXmereszuRdDF7622yOPxBNJCH3N
YJ7024vDV+LekWufn3VHXD0Ht+OpF1jOs6bUsyZPODzUUxmmJ3Im57af643uE5IMeq0g53NGs3Y3
gB6VFQIfXXAVRrm7U5PJhJ29a7MHtoti+tvgGxnLJaf7Qt6yLAtyXmomu1ffvK7m9EH7ivZgq5lJ
yjfMQfRi6DRddOQOs9bVo7HD3cJf9yCzfwzpPu2DCkqSnEVS3TT+FgPcYn2KQFyhjJJnir/7pK+Q
dYK0XWHuoc0pjGU6SRMyJbF6wWtMlTfobASFQYQVXtK6GCiFFIIqnGLv5HTk6+hj1af1r5/lueTj
7qVujRk1w6klXnRSnlL0PY7yb643K0JsUB01cO+lNm6XQXH3Fzz4WsI3rL7zJzaPvtly+bQxX3qy
Flm9Zzs88YbzCoyloudjL/BkfCi+5NuOF3DdePBkGFS9bfQYLarUtQrd2AlHLeGl4w6Try9Enl13
y8MTEqvGTyM7G8QY/DJe3T/irPOHxx2MmPvit2DekvVAI31syEo82C+RYNonO9PK9aAdzyz05tfI
01ekOuhT4hLOWgE+qBIbz/AEoAFlMz+swzqxDb+WN8SjHo7H9RMpKpC5oZS9AQxlWk+CW51XzBFo
E/z0AE1z+jymmHoc48FCJObx6GfL5Vmo6TocsjTJK51jDgbF5BDPVXaj/8VUBNqTsrTKFWNI1Gl5
1jIXU2xAQCOfBtVsokAKeoLUGDEMnVfOYM/Eysnd2ivuNSBfxZN9cD4UL1fbXrlmXHlj0/P4EpUK
owKNAxiX9RjiXRQUCMg7DyidxT0jG+J7SkcNVvU/druNOxzZLcYRNqY9s7Jr0MCFmvaRAwN4ys8C
YKNdc9P7l7GHrfPrmUmMNh4YgLTtaDr+eVlEGwzdriAdCGo2Ev5W7pcZd74tKj6c8ifM2GL71E26
KJzDV9K+f17/n9jXQW1NmEInYWODStlf/X1tl117VQKJ2ebgGtYUUSvwLBWaDXU04ybGHeyuPSYt
uIsqVnngzdoEeCGbsf08PIYY4MGpDvPFiTG/bvz0egBjRvda1kbegZSC0WlbyRdGBYMQLFoSMM+N
dpBY0p9m1vlmWpQ1NB8JhY9GOojw2iwv/w5bnx9/vUhwUbcu/EVWc6zk435E2gvt1G7I1tqovzdI
fReuHqgc6wUzXi5cMgS2G64igsgSV+RbxaFdmvErVG4GEaCu3XEZZhhO6WlJGQz6vbJ0rA0Mjnsq
b3ox3Ub+NDdSN7LPS3k01o+kdXqWwlxSxAWX7MQRrtUc1rIC7osMLbfQhMocV9XD/GmgwGXn8VQi
owCWAnnfm3zHiUoSla1gh3qLqviSgGIOdV21sasl7q6Lk2u0I35BQrpT9yGvpa6PXupTYrMOTXK7
m0g/zzSduXVYX1MSUvdEAxnfwk98hehyHeHFZvkJnCk6BfD8AjfDBmZcGfnzBNb5wbn7t4bRuzrJ
YIjEWnw7b5fhDKDOx/r8UUoRPeu87vGBP2K251DoykYGyXbGksUCYbzdQYpwuyzKLCluRe74nB/e
3cEW2pwkwH8LvVmRT/k7NJrWz7afIYZgv1Ygy0+T08vgOYqyE59yqPpLv3UPqdW9vwQbH3qZ3Msm
0kMD/UmWFRcrJixRyGkPql/udm+tkNThkphyYAn8nH+LitBP6zECnauipja6MnJQjopMV8ui2eTL
UsfHJ6gSscgnI4zWi95kukPlrcxSiRSZhWEWXc1+gu/edUny6DANj6jB+0Dg2PCH2bdgKbK53n/b
FHoBNmer98tBz6kA7FiSdMpvZxXniciFhbxT4kDAVIqff1+kUzPKfFRzsMlMXBvj6zHsBLphZYJP
JUwnbNsXQYpfYfiDoaEaXnldwsiReiPlweeQI06Rdhu0aIsZoKEl2Py8eqjKr7HVstgDVxuK9msd
tBY1EjRmi2s560dfvbcR2z0sYN7BAQGog9hhxHo7+YQSRwzgjCrktpFvkAlYWK9PfrTSqsCwxbyy
k7HQPKbvsDzzO/ty/rAb5KMiw6JtHVyfDymisiBwOd/aqSy0s4KveukkKBoD0n6g0DgOFPXrwzIP
dCi4DQD0ag4bHhD+sSDiPzAD0eIRp9OyHhR6H8au2O6ivycXUh6UCwzneu9zPfIkLvRREeyM0bfq
WeQLkXjpvfkakhkjwzubIuZHbcI2tr31ulXfrjH5mV8wwmalJ9SXbHt7pjYmNat3FVquqp5a92XS
X1dQ0Hma9lzDAXNHJ/SRUuOiNTlmSfiGY/jF2rELdCF8C+V+144QPXLoBZsRk84E5CXXYE4caASh
qpIVe1O5vzSk7eufLOZ79HShZIIa+UaTndPz5bRoQzCJpnN2yc3YMzBxzD7JBBiFM2UqwRV6hKlY
7YwBxvas1TJ6FGbkFerPPSJLjeif8kYKnU9kNkhrnZf/N4QOyJBNKPDeW6dJa8xQaing4OI4uG8h
dvbxm0SdgZSNSLt12wUVCKglcR8J0pMcQFlz64EzPHTZqNFLgTEwr4t+dQXWI/kgVcedsk3aTzjD
vdlblFz8efqfu7sNVeAW7aPWPlmpegv/ayBmD/koIaOns0Qly3WhSq8SLumsdHzzOR17Yufr+TLr
A5TFAGN+HXo8vwVzoGpNaDwh8vS3DRo9s1zEcFn3nrtoDLbzmhwusRiu0GDvf5+0eMsmrtcJnZ+N
P/3dfFZqioxvrpmKyKigmhMlW17d8S8TKVTO8sPs+kDDw6JPngWSVWdeRkHTgtoByPlZsHwvfumR
KYS18/fkEZCYJAeuA5G4foIHQu99s7Tz93lq95HT7aOZBu0hirwDe03T71T82xg2FNtEkNIFMpus
OJQPrWAst/fVTBiAtRk+vmkujWbplGNiGcVItEjTHtophx2xM+a7s+KA+g8MpokvFsTGCWeV8/oH
OOt+UF9gx+fvQNAARS889XtVceG/IzF0lIwCbD/StdQIt2nx9EcbM269+X/BJfx/gCZTeuHwiO3d
BqCRdYzdXWW0s9nmpzt9CnZObkU0pjcyE7/Mec4x05h0ouskzk9DFVOuttt++B7WnL02dnWFohHz
E+H4eTIMcY4L978RnNicWIHI0tmWO/StHMWn4bkrcYBvPvmF4fP4Uj1qqRG1GwUUDCOuaEKK5khs
MXK8iJxFZTvOJRpruwHyqiXllvDnoaMbtfkF1dQqX6fC0eBuIE5Pq482NeX6e2u2cG5UZ+k09JK+
mgFCvCClrFBlArptBq5fZLD2Fm17ZZPqJXEbSr4GPJTekLu7YJbPf/fUilgx+AY4yb1j6nev2Om8
g5P7vJYSyocUgJsMcSY3EZTxKFSMbZ2Xlfa/NeabCkkdAcWZCijAggJw55W1ltRv/7A2VlRXnuyR
n6IkaBEHUr13ALpLe/8Wq1oj/tmXVsmQHwD1lghze7H77+B0FKBxXMLdlUoanzK2LQUa9l4H0c3m
XDQOTNRrpkNoPQey8NJ5lGc93YXwpXH1yt+zGq4m+ugJvDNTHpRRUkB/BcqVXflwrnrXQZEjHDJ+
xreorxBVLIYymfVSCBuTRzAbs2PbJRBkpgTSYNVzfUr+ymi0RJQLk4LUaTfhT6/4XdP9g6fmEUrs
LjkJjxU6bN91PFDD2f0gwdXcj1OZkxKoumsDqlCSpj0YlglT/ThHAYCl/xWOg+ZZep01pUPO5Ezd
NF4h65+keN82x8947AdAOOrpSM2k2f7yIa7rZ9uoWiiBr3IXxCb+eq+QLSBpENs3MwQ/ofMJB5WW
4qHGSooXnkeAO0okop3euNv9DJf/lt5+hocE8gRRQ29KlGLT3uYbf1Ci344rQiB6IKThW7rRO+As
zehhTIBt+DJG4nd/0dEKb7zP3HwRmalT7vE8sZhOVKn44PzlImxnzFYoEXgrfqInYH/GUGC8ZE2x
x/OvBByfppKPmSazji9RjawEeEIDi+Isc7pk84/XStjdXpB0XWq1OxUHqpfopjJ9HaCIrh9/vWbd
g2beVNlkiWX1i3misdotfxYqIH60pAQwzdINtk2KZ2rmlaMv2J2BeeWb0VFol7TmI6BSDMXit4sX
anBw+70xsf9zlhq6WHI/BJSYHstq+3TxGqNO29y4jGsnIwSqEs0JjQ7eVickfi8lDqggREtvjuYv
TNoDbW3+eY8J+QcwVvoUsRUzo3PSlwpmhiagR/03odQ0b7DAF4Ff/W1m/z1SJVzdC2Md0Ecv1gnI
J/abwIa7nMNTIHmpFP9112k7nu8XxHPACTgRzXyCLE9Tch5hcVoUWM4mWvVkFpZ+mh0Yph64j/H0
CluqAf9rDIVTD1s4vr2S0xDMemb3VdYDUO77E6kUogJ5fuxJ8b657yyXG2NjV3JC+cyBlXfhNgi0
9oyv7uvKP5JXFeWbb1Olp5+J+w4ANQyhdcPwgTYuTZg3mukzV7T7g1Xc9zAZWWszehr1tavA8F0l
07rv4goQYxZOpntvfLmhtpge8zVmruqe2U6wDQZhIuyFxJdFXlNNy0uh5je8XoAU53Yl8croZLyv
xqfgQvwGNB0Qd4mI8Jy50P1IjHEFZW0cDXAuiRWyA5c49S+MUyfSqZSPe7z0itM/10YsiOeawPj6
5AEpKT+HXA1pHycBzZofBLZ2Gyo5S7rtx6lkS0gb7OggETnW8XAStH8dZp1Q81B8eOQViEnUE4TW
MfNEOpZ07EzIy8CdhzdMJtFIu9kEH/xramaLzapA4us2og1aVum+9nos4/+2H7btj5ZrI2aMubqh
YYDgYbQefIiIfdJZDTr3N5lJsVC0OKDVYh9v89NPlFuGxMh1ygESrIZuQdG/oMfbPzQW+ivGhCVt
y3p3tFGyGHqdvX2Fx+zvBwC9+Y+6xbInbKLo5ciImH8DKxOz+lawaXhzyO1vxA87E+uaBw5+CKqe
I/wuz7BN0MIsJrbcqGIBMQ5N3NA+vJkZQ+L1ts/BZjJgsCJyYiTId4XnYLQU7tRLlNHEBVEBDC4F
CiLolxl1P7ldBApfWEILP5pINOP2ojoCaaz3S6n5UkzPF5/ttFeCVZncZmGJhPtd86tHYLR1B7Iw
GmgOWhinpvJJ/f6M9QUhkRyM/5VP3hksy1EuaMWrBjK+osWgrGaW3EbJkvVfponYyUAOuEEeLOcB
u5bGvMfotAR61H2xgGyz3wDTv+xDrwqoib7228d3/EH9KNYMq/n4wvPIg0EyFNBX71xVMFBhw6i6
dp/GplJZGcKEiT41arQnEHRaHHBxYYweeHhjWXa2KQqSjOtKCHeg/pgp5NeM4s87ZvqaEAG3lAeW
EXJMfu6TffALOXgPLSak9ZHwqy3WzocjyUHEGYUVvRpfqVyTyR9iRwhL3MR74mviZPe0/b2yAzQC
MTCvPg9pE2hoy72ELsLVZMJQx+gef+gCLzHqrvliPUVX1xcBoRgf+oqSh5O4Vgnh3AveA+P73h5z
sZhPbpirQfBdqEVXRiq7ATIYE0GZ2D8/1ulXkxSRbC41f30HG5rgSoU1WBb4uCZG1i1r7w+0EZ2A
4nweOSMo4exEHezTBm3CUv41AqcCuSPVSlIp0db221VYDc+4cY5+iya36j/R6/zeS8sLefBsfWvD
k04Fiz6YJ5C6TSolBviXTUahcaexJDLnEpvvid/yWM+2sVcnF4UW3sXQ5RVfWvc48pD4Dw+PcmRq
cZkyoRL83YNGvy6tvAbXVGcRwy3JBzwyS4gC4OPT8K7gIGdnr7EucA0dV5fv4vpn2PvduwYU38pe
b5A3Ck/VRyNRUGt4I1NTrM21eUTXOgD6z9k3qROTmXpncMe3Z0HahOahn8rSmz/MV/9zCxdflji6
xmngFgKb2D4KHcyJmCQYBpwxuEC8b7tJZG7nw8Pq88EdPK0/myMpEfq/YNwgVq39plp/g0mRr9tL
EMHVfBhfKJBrXiMhxbsGzeLz0Yvc6EhIBXbviRTMOwx45nRC/41DcAACz4FHjJp+6w6uOPc69hrr
0/5XfXtwafM37huqaGXsN/ZnoXgodwwbUeQyhucEG//HsppATLSaGwnh+/fUF1KdXXpNe548FycG
IzK36zRhvZW4/zlF/MjXLmSIHISDQCGzO72eibCjiyFF3SLraM6jx3sDQE87z9WCbG+6KmoR8uH1
izIc3/XRy0No0wbh8U4q5JH1jI+JMxzs8qOpnv8HJxWdZnmSwakn+eVRmHNl6FCNOX1+HPHljq7f
Hf9nwDZbuIIzIDs7bskr4ufFSRxhh+mqWYJ8nH7VTBkFtMA58rO4QgtVBLGK24GWpcmjCo1eq5b6
kUetSQnn+C+/KLJGm+2Bx/wSa7oFSUdaH9emAjHHegeJCDUPsMmqEoRmVTxIXXNcr+GYQvWaUpXr
oehb8T2Emg9nOcYLzjg6I2LryDcecPFOjHPnRRlM1HY7riB3lOO8GQ7Xu31Nn8rYh9zUOTgTbAHG
As7R9OQgpe8Y4xXNet8UbYjyeMfjfMc0UDHVsRiYXoghhSwswf727lpwG0iPqgYv+sy+llkIHkRP
OE14QyN9I8LmxUWmPzNMSP+FeSujbZPhbpiuMC2gt8eH1BKxfCZZiQe2qK2U25U2S3dKAp/qkIs6
titR1Kl2dBiATGX8oYQYrUHAmPotTrFNq6y/qhdUcmH+I8KAWn3Rtd8phMtYjSKlS1cD+Th828Cn
HHkSCzgYqVtbDebfPOLm2waHt7CAhkayK/bdMhCcyRUCiQEui/nUCbJ73BjRMLeYBvAfAF0/bqs4
FT3FEV9kikjbdN6kjZeXg7IiHLioMXZXyNlK85TnXfyvLF4WHp1EkM3NcF8RRDbSMeorG06R3GO0
HlRwvGH96y2573db+IbakkRClO6v/osxUu25t1CNjwGQLQmnOtU55T9PNflmQVTa/B+rHUrhGOQA
2+iqDmwgjORv9e495NsBXxCRuhVBM8Ql5psNysJMmj04kffJtm5dSow9LRyKhEjU0l3YzsrnSAIS
Srg4pJTLZpncPxeWi+Y5iULKxq6fhvuIHHVYp+DzL/xwA+h60uFvtJvqxxljl7SA+02AWvtuyX4K
X/gq9aiV10Z/QnsVwHDTafVTquc6fDUwHZ2gfDZHuk1lfANVCFSlQZGttuH8dnt4Fpp4yaOxkbrG
1JwKwskp5bh/hP+E0cnkllGds+tPJhJcPZtOm1pMA4AC3DGhi5NgGoAc/pHKx0VBZLzaNtqvIo2x
pvSNge5sjH9PRBEq9BcumdMxNewOm6nH+jShuAzv4lucdMY3pfF9/rZ5HKfmzRRp5fUAw+ynRiYA
AFTyvQ0BEhF8jcqmvwltThRKwks6vp64qlMPqRyoksuCLW+BBzk5HcpAc0I2IozL6xsUeuC+5sdM
0IeIdyO9f5sxVqRkfnF28AdttYzMGeNH+9NQvFner7KAbxjF1Blkmnp3OdVQ+Z+xHlxUS0QNXeV3
e1p2OnthVcExwBpvIOzX+3T5colNvEXheO4kCDq3M8dOpGUUnIXddDxo20T+XnjJp/fKQ2/vVXh9
8dwEIwu9bUYGlcAvb4jY8KXxa4o0Fd6LmTY3/9lfPXVV6qNnQA5gJoPPGzGiCoT0/G3qT9x/ReQp
0G+v5BO4AtrmGM6wjXk66+5XtFZqL5pAKMmgqj1BN7xH2ey9aDJ01O/y6uYrwBSveQx8a9W6K9oY
jzcxXgt3q52F0rPfVA+KnLzrUpPlRajo94MqSm8Tpr7otFCJE8AbDwxW75KxdZFETLAWayI/pIeq
W1NziE7LFPKapyHu+L4MEUYnynb3imA58JInJ3HE6HXlJYcFo+Xq43Uwf6qtbmyTlEIvN38ZSCX2
6aWnuzwuR0Yjzsr8Ys9nsHWhakaMMk5TBLeF/NrANaltzKQOjJDOEZUbyqAeLD3B8Gb3FRsopN7K
Eb0GjV+quES2eQH86LIm1akDMJQ7ASKky63fzQyL0/SReXISR8Z9OhVC2KppRf7N+lJq2HK+XUnG
JPozkKAsaiJkpm4C3E8q3ekCYir0KTN/GFZ/FL1zL2gmg31oRZRaKUDHZsQlQawEUjSc78fTJYJ2
/bWBBvprTBdqA6dRvAkH8kXKLYmJg9lhQge4T5nVRdQR2p2g+aUvuyyyvh8Ax5Eagb32ot9MW3Z+
BuFFVRvLj3nTtOpYu1E4MiLjVjzKwc6p2X6YMJZuBL7ihsBZNmT0nqARSLK67qI5ArrHbMxCPEgc
5oU4nOOw0REtEZw4/GoTCJKr1/U09nDQ8WBj7ZDhWo4PiNd5fHbBhfUmTSYOOT3NeQN4LKmKc9av
F6sx0bO7mFfhUddxjKPquDMF+kGQn3NXaAV14DTVrOsyQekeBmroscVo+AgF4Yy8dnKMt+R30jju
ECSbx+OD+r40L/l1H86LwGrHfwdNjlHzRmsqD3UUoNiZ3YN4QvJ2XRlOP35dh6V6qbybUTkMohbe
8X0kwvoKP0FckVNAit2VZOrpOdNCns9LxWurWWouBSbo3AQzcqd/cBoTypwLeEMLJAlQFcDD4rHO
ulUGuIE5kYceBCs7TMfG6vRmL03yBYNN81knOWHytXDOdPhtEZEVUl99rx54jIFJb7bjRiXNQdmH
am13Ut6O/SzNdSNicL89Kvem0oS+LQzCZyjBVJPEZ9rlFq0g9ma0PoV9N6ZN1XkDIKRvxLNRPi3a
RQfp8ljtKgA9JCOtWh9vXRWqNMMmQKZkQsznKNYhHNm9S/hH3AMlY65u7P29lYE3GxvfEFzfQSvX
rOzSCOc0NAmBM93ykPdLZJ6nRJmCNZ6tTjRfPRsyaS3Xq0fh/T8KTSRHpYsz0dKWfqyIEAO6ZajL
9OLeVLv16GJxRPAVFstNxUuUb+leXQBwp/aE7ldYjdboXPmD3QOjMnOvx5WBikSCXLEGXiUsY3aV
vQSXzTxaLpPPC+GDuso7pzSLosXywhNYyfWyU9zJK0hDH0KZySUPTOIIOE0rYKXHGDtVg2yC2i1t
a264YxYg6EGzGMz9ZdU+14jnSN5UViRyKzH6VgFR0gkmmaGdsm1sQEOCYqgmc5FB9vn6tNJEpUQJ
cBiEB20ogNbx9giaXEiEFqn/Z2BgAdlxrm7r8b/g5ISPIBV9pHoROdFhC2dtTD0EgwF90aMjrhy0
ug/wvD09P1sbuwIjYvW8A6ylCWjW3VhUEkiv2dDmNQYT7ETnHMhST0H8E1CqaUUImu7WcHVB4eUt
nmlaLTp7CWSW+A2rtKLRJsQ9aFb7mpNLm5bCzlyWejvYIi5AGTJ7wNbmwKEdNcY0BWbTq9zv+MDg
qcXrNPvAqBUrwbxMLihi49SaK5YXydi7yIfZpDnBIw2yVtmyTSs8kSNwbmop9eBJRTwHIzyPKUCc
0HM9t8x9mmb5QbJPzro6efLj+1LhSZup++nazawsK+bwZPZ/YbP3JjfXq/5TM2Mmv+iodmEk3Vzs
UYmFdVcHGcsY3TtlCDk3ndsl5p1EsFkcCHMI7ADoInqO7A4tV/j1oiCopmkjbusYBZJeHJtnrsWG
fgoFxUnIpZCCZsN7xsxvr4pGXvJRXI+ezuzxO/kG1/Akv9kaQd44kzOujEaJrDqhIyTKUllWk+gF
imzEWOFj6oekDIvSSAfWurQbYfQ/6qAXgFxxSaQ0ggimysfc8He6n5nAijb3ksLuPlIwzjlB+CDL
xVAJwqLiyu05sPZT/cx1M3JFnjo/64t25lhtYZ6UDSh4QPzaHHVlyMIX7M7QwuLr+LEZ0OmvRc3e
vvw2+SjMLZIm3Nt31bZxKoZFfuYWyooyoP9T+YlnsrIyCqC7iZXgfJTMO/ao9O7A5r+eVeWQEUnW
9TVv42ugo+6NwlrvvzcOR/6FGSoTrRcjJcszE8Q964EMdxxsHlSbkNbj4DrJgZ9yRXCgtbq72CQI
XZ7T9lv9rTTSQWFvybs81JqBsP2aHXDCYZOfSL74S0Ke9MZnR+Wqx4dFIfILtSj4phw4nOlGtSYM
52zBLbr8NYsrBJSWxKuJzu+z7IQE+H1Z3UBw1euQRqOd/5b5AHUSWvrB2duj5O4RRNnUGA2WViHr
Eqs5CdnIkWbbke5onKSeAG+5CaPafdj1tRcfvF6n0mrUbrY+rD3riFXhJ2msXZFazF6AAX1jnuqt
cT0/YsDhVy7OyFSYqjoFCrT5cInyHSBcA6QZtzs9DOMe8DUtIHnjbDFWWYB4R+vpmGdXfzkt51+J
xILuuInM+AbFwzSHP4AgyN1vG1Gue+w6c5eOwAexxwwmcyxrSTwVl+ujVlomfxzs55G42qOiVLLT
/gmDsX+z3hw0jxcqt9Sf16Bay2Z/+dILgUyoURpa12cVDlCYAlxuQ5eR16qFgHP3S/Mf274+Gd0H
gHX9caEWKJb/15LEHDyBDg345auBTMQOaN4lP7BhS84gfcPZSnA/+tRp946mSbpjyjlZIyknLt3i
Ll7OMQspF5eSgbsw4+zw5iHdPuP0FtsrPmlbURx4PSkCv2hyYTx+IXRjqywcsI19kn3K7mVBLdlI
dg4VcYgVELdlGrNA9shjeiWOWDeyjezAr4svL9hzz2zsOceSPvRTGDCB1v43IG5s1sl2qhhqN+31
BQAN7Mx0br1kpE2k/gBpJmRQVlSIv73LNXwLdKuWihSyEiixaSs7siaofFBglSxVgV2+DmFI22+T
716APk2zMBhdds33ABGy8+mhVWnchUT/4sZX6bcHVOLeE0qhj600x3aQQrUpJHTAQb1Z6cew6lqc
P1VhchFrCeOg6tFvsy8NLUcBPkg6s2iLio7t+murPzftIvc1ivpvmTkqiXvyHHzNGxaufYyOSkpH
k1KbktL6U0xmytY7UtSS3Pm1A3704oYsZFcES8Z33C2xN5J1DTqyLmvSWwSSLFbMYFZdNkZcP0GK
0P6hiX5dycXHdQOnxH0JFZXGh1ji3mq8DjD5YiF3XMqpOFDwGWP90ERH+t3Y4IpCpw8Id4s+DMbJ
nh5KtaUiT4a94EhqbybTJaO4h2uFC60UV7SxdhTijiopuZ7R3blCrgr4Y95/IIH/9Lx2vwORS3gr
D+jMmk54uy0eHym99LoIVP+LitTRnhxtREkX/B9QIq8DyiiQvEXwVc9bfAxrG8HMCxpAPXyrt5V4
ZgfRQVZjR7TlSzb3Dqko6epQEBcOGJ8k5J6VcIRHPuyWcgVdlj+/7H0KavhMSkZ0ETFMKfduce7i
F29KzMReSeKw/K34Fzn29Xjd1biZERjjEEK8YZdr7SKP7sig7JokEAUd03j7c1ADWRwtc3owKI5n
52ChWwR+jHBUMQ8lg3hYcoRn7vSR9sYenkkad7VQnlt6G+/LTqUJNohSaHBjdakLdsJHyJxc3cfS
mmUmD6BBu/fCbAYbUUjore4yKryw4S0koB+5nWne2vYwlv0lk8OtpbCRB2pYjtGK6sLcUkvHhQkH
CIjJ8SYV3icX4naZkXfgsGG/VZdef3kg1K1kQ+yosL8kREOE7eDIXFofFOkqWRVr9UPdbcebfRpC
U4d6yYN7K/5r0AqYG7BJajS0j3kWZZyzYHeyjGVaz5PKaktPpsPFFb9R3b9opZEE4tSV4eEzVADd
mvxAl+8MfG0EnXUq80NtZp5jgS3HO5NdtDnlNYHoT/qSJO8DTS6FZYMcJXGI5NY5F8/z5XIVrMBH
TxASl5zAs61udUqrVQQIN9c0KdIHzPpp7vbjdQ2+eMR/OqDjanF+d/lb4EyJ2grM6BNjboUYBsPb
MG3cXde6ATQj/Hcf5Lp7n7vVW/5o+bgKwfrmmzYKYRryY5Q6J/CpLIWmfsda57XH9GTdCMWpRYzg
BPbphHwZhqCrxyliTSPXOP7NuXGZOHHLEsDt7r1041dw0oEYqXyAbaGeOpGjetW4R8S8UbLS0SC3
W8oWua0c7k2JUKKNWq2LjwfncdXgecPPcl+/3dzZfDuUqYEiCFnOB8ZxndbEGAfU1KWV+KOoLI5C
uiBtujpnQz53MXJ8oNo9aZ4beDxIMlLoOM2VOOERGD4nDluAenPhl483Ol8yrWWu27BKTh0iaiBc
eP81fkO5XKk5UA3iF+dALE05lCmJ4C3JbDlfrJllB4vc4xNaMEP9Zb6Naat5MExA8GNhSBQLQN4x
LpvoZ04hbtW4naVnvA4Hhp4AJ9o8QK0nDGtYatsa6lgFQLvmNMk95gVdBsvbAu0e2JvjqwYB3n93
V0rNwBFUJY8R1NgEl2W3PW/VW/OGKKQL9vNke3rLjnaRCQSUcVNoaBfgd9curZujwKgAn8m/5Y5Q
o2QjAut+PFHtzKxXobSfuaBVf5RKLSBkD0HOtuRat9wHS10rMk/QB+0nEoI0yx1AkI8/w3jH1XWB
/TPrKndbteeGzsPvTVTkhXaBQ/DUresLxbM09ts8vu+pL0O+a7a/lYsyjyUJoY+nwEQ3adaXrQRB
Hh+79ZhwDnU7JF2XxlyO1mUuocLR3Lc0f5CgVUvwczmufP1UIIm+n2AFMuqnbPGJPbYfOP8WkL8H
GCIbloNxEsKSA65BiJll5YDYpS1l/rbvK7a9079l1cPJ1Lrj+ERFKm3EcIS4CsFNgPV2bmP/zSlT
JALGc9idPknRxmro8M5wYxPqLJ4YXGyy/AmrO3Y+CQmL8KerETNXslRiL3xjaG/pW2FoPUTa2aIc
tQqaXEFVpz0PTCg/rmoqvVasuXZJszdrCvw0qRwCA4x9oxN6uY4aeOgpwoXEicXp3krDeUe53tzR
rZZy0Tx8hRChb+CUn2PqkDlsx8c6ed97S/OTqEC9ncx01juNnHF2qDUP0bnBeJBtbUXCXm8zK7dM
c3br7b8Fw3ULwqU62rWwogLYDw4G7a3iadQLxQPxzvVS4F60Q68Zky8wsPi8znwVYfWAH2Z4ZkTs
ajrIB6BMeGNuBRLriKMH+AMvhXH87JzdsozYNKaTZEb6VHZxPLHBnv9exuGdYsvG0ph5gb3Xp5RL
jodpRViSV1erEmUaXBlvrpADQAipkVYBgQYuIOr760i5TTAzEn2rKc6eoTmZlILqDhIezY11fj8B
CjuZm0nkFUZjQvyQCbYRkpDDPfJhErguYuOHYucJXtDhmcAiPrCyeNF1a9MCt/tF0A/Vl+6D/PcS
RNLRCEevHzNdcc2V96VT+x5HwRLwaGC9ySkmVBTSbBguHMMPPSDugXrfXVbFmzZ2TRUs0OqXEhZ+
Xkn1odWm6VOqPnLZrHCMnCvOcCJXSVRUyZhfkpKhFa4z0QlBX+V9Tyz/N67Y6hrWi+F1TMPc9cqO
z4zDm5OEI/Gpfn71Occp+3D4/jmmm2M87AMWILsVCPKDAAFo13oT34A5eFkZk9IsJacFjE2HeM6t
wWUu99Rzx/TOvgc9m87Cev+REPQTqfDwnips6Q2hT3PvroR296Bb63DXaPbcHTDLEQYM+VV6olfB
j1Kc54b65iL8DOJcQ/Sjb7WHV6dk4CrZdFGmT64H4nww4Y4ZuuhDNjhXD8Ak5RJ5NyJAx3WVfQmc
vwuBmzzMwG9w9lOaKdxddGZcH8rGiaOtXWG6+AbUmV0Ew+T7GLbhMQyr2CGfZb0v5pF1TrL5s/2j
kXt/0UWwwyNbvfygoTlvlNqRZTUoOkaGPaAftDumETmm5+VD0SrBaeWNLVyhAyQH5f6HNXc7eHt+
H0YvlkGlbwpK+wOMwDGOD40O8enb4pzQkdFuc7AMdkcCXs/+IQAZ+9tQxg+xOAb1EsIzUO/WYDBh
m72XfjzMNt5AaRtbOC58edkKDv6Y5GDCYHodRAUYNYw6aR4ZAcWktjiv78rEDPssyuLX9Ob1y+H6
spqS1t3QHgPH/60axm9qWAj53hfcIfbBrkrINBPMwXVbMa+R7a7cKvVFUg4ewSTtVG6exhf7J8XJ
XzmRL2ORoSv7zGllgdk6tOo4RZKYqyizNs3DgytMr9H46RzJu3ABNrgmerzn0REtclc0a6IjE/wS
YW9cAWFkz1StcuIWe/Ei7gW5bE7517HBo/fMTSNTERD/g23SM6cd4k9bvobCvWgKXgPRGihjOwha
1NHIkZe04NZj0BJQopRDendrPx/HYzRv9TCQHEifqhcSWbv8x2AVNTlkvbO+1tG8N6niA9vzNpLS
SgVFaCQbBKaH48ytErfxQV3Iau6XVXIVsVD2lR2eLmPGV69JMSBCZdXDMAEtr94fLre8OJYtV9Cp
jEdawDgBuXWenLzOu55ait7Bc084N/Htvpnh6QmQUb5vB+6Y/Gu05IYvXBv/6IOeD1VQHvoy0DpA
hYwiPNS9zuOs3NnJDnBFIHQH4HDyWRouvWvUHfGmpHw6dKv1w0JyDR3Ve9rLbMacyRqoF1sH/uDq
1QeDc8/UvrJoJWG+iKzYLQs1j7VBAd2PqSdyNrnzD8treypskRSJgKJnAkMoZZdql5n0HLZM7yyj
/tzkG8265JYfN3sjpczgS//t+COo6IwJHeclF+LBsIWL0/IlHB0VC0PhcE1Gwl5qiFChfjI6e+X4
oVB60YtP8lP9SnRJdSi1YcVJ1UWmOKq3z6ueBZmf+S8UzMC14OU/aPAmI2Nb9loSHLrM7frcZwpZ
m/K1vSCauUidJQKknw98K9pTCcBfXoQhf9n+82UJvhowbTgtGPI70ohGn891Rz2fGY4qRWaGHHf5
N2LfPBBHHIlJPC5yd+CRsuGvKxGcQMg1icYQyqwlpcumqXgkRFPc7pm0b6lap6kTdG8JBRiHET6+
pSYw5wRlWW/Ysy/scMmcT+yMOIAqSH03sdVxrbnMXzZnVpJvwo0hNfpuTXk+JUTz7stVAUo1O3PM
VgNZZJdmfyJurm+JEiWJTABXiZOnTbJ8QI6goUGOQcdHDDCYQDRMMDblJ3FspU6qWOPhxgiipBLJ
jcFdVISrbao+AmziawrDWW5GaDU4iC0KnjZ9PzCUAY5qFu9fgVTStnMjZmtCPGFn1AZlf4owjWUK
OSIDclX8G/XHgHCZ64FjBpj8i/WOa/a9WWOSu0IjNGG2NWWANsoIHwxetEfAM5+gK3AN1GB47tk2
frkK6CaDS47jsn/E/yFVCx6y9SgH4FmxvB4WKcN1SL1JYubBZfmxuQ5LbdlLGYxSXUNtqYsae2Kj
jp+bzfW8I7yclxsPusEwxSztjtwc0vWPHbmUbX+/f/hcHw8RiA1YDH57XsSTcUJCWdj1DA0R+SAj
FsVTpTn6/piPbSnyJx+pi+xJrOJkUp7Nlbe3lRs9M3JkMoyARvpfxSKEH2BpY/BG2MKP9jJzEw2d
NS19+wrMfm3sOOaqfVhYTS4fSWnQ9YeSmvPiM5Bz2TgzcOc4N5QIpZcDUtgGlWUwzuu3/dEXbzJp
grdTFWq3PbrgXWk9ef8YqS6vBGXNGk4aiQZ0VKWu6f/XBV+On6Ze26WIUDcpGvCOJRVIDBOHGHeD
LKyJm4T6j0lZZIoPROU3ADc9voonx2NJ2/UxxultijBLcFYF8SRrfUyCnIEJpx09MIZKbmANjMq+
kDuHAsJBAjW861r1842ipTYlG2/efG/dNTrKcyT1k7vGWilBW3HslOUSlfPFuxzR1BMQPthhUegb
2n4fM41BftMBKiN1QKXHeGOW7Au/KVkjtD1NtQZfGTsQ1975is+rtGS7mlbSaUyddVhTIROBAw4P
7LrVFB/guwzIRZEVJLrXEMmklcHAVoFSNgB1f4AFuDkW38nbizzdUdS+svPSssnLKS6jIsfIkG0E
rYzQ+/PXh1A44CMZI/sbjTu10fn/TGAbLcawMxwId6pyEzS5rqJJMkYiG4K8rFdujpbM4IkQgvh6
j7m8Xsoace+i3Heq1kBi+NYxhC+MbhajmvofkB2NEn23FcVXisRVXU4dpBdXsLoS9aPVC3sEOEPW
N9ZDwK23hDLu6gxok7dcQ4Wi4Xk9VKmiZ+cBuj6+Cc1mCqGW4eQ7Kyq17/rsgjZOwCtQBo2kXBAU
g8l5n7we+ZVjQfb2ON2TJnb/ExIO1WwTXMYihCUEJEh/wskot0kJ3beuRspBqnJbJj5Ij0CKUrDs
bnvqbsZPHNK5VChni+r8BMXgLExb8OOyeCoXp1gfb6OfQ8fwXuxrX3XS7+u6k4MZl0F+Cb8cJ3vq
J9Umh9X9HEgQugc1rpKfyMKxQDiZB2p3qydYg+nobRiUbOpeCizCgPNbCb+jTLFkNHbQZCtUNXOs
SfPtYTk0b3h/33brSF30kf0QNyxFz9PS9ziF3/yaCTIf2f1UjOYz4HJ9mkeUUGQU3tSqU5xpznXG
ptcIln+8zuDR9G/cJAxhbEtj1xiV1KUNP/zudcBSweOI7bp25StkCH9qsYOHIJbH0qmWuQersRp7
qJx1dcUVZjwyjKbNtIo9HIDoo0Y8hzSrS+QljFwQOJTd/IketI9f1itJ+Se8N8XFAdxGxKe0Qnw5
B2nqcFD+xzbhFjJKcpavMc693lLT93ovSU+R01iobRvCr7gj+B8SrjKlpdG+94ke4sNYqi6Ktj4Z
Qpt4eQdGDH8P1YsU+gK83rlQ9FZzRWpMpZmfXXNL9qyVTqXWP4WNlG/oPBWMFQKbCfozgzRp4Qy3
BTQ4+cjfNQCp0w6t3bwu+bzOGn3sqd1rRZ9qARvs+tfWPt7ZPszJyIjGptvHpA+GRhqygimX6wIF
dOpa3KJwZkSHhG9RZJQBdG/oahS53rHrXMyujUpMRZkd4LDt9LlNweCKBfrJUcYl+3WwrtewFLiz
8BDR43XvjkiX9MSOCmOBWVrB/rJmIf5eY+KZ2adP/PSVuqqwfWjEaL75d8z/owThl5uP5MTnVR1I
TEgLhu+BFeeBOe67c8rxH29gqAxOzRphdXyD3zQCnrp4Pk6xRBNFOfSD8Rbz0ugb5jMoN9cVwub1
BMSoj1TbwxeM21SAHDo84jZ7J8COE+C6VJ/3lEYA/3jdV2wNUyokTO9ER7mhse+GdFx0A4YTj/x8
j1cMQGG23c8TlWRoZEaAwizvo6s33bt89gCLGYzHrmjWWuxNtxDVyF4ef+lGzJ5Ibo9Hy0RA6ndR
0z84vi5APBHT/9DvbX8sXfpbUuWcjvOZRr9T2HWP2SAk/D5FRAop/P+9cc4u471yF7xNPdtNN84k
n3SOW13s+RQi6knFuBu7NZXw7Kcy+YRm7vh5CIPOqWeq3a/DBfvSkm3Aq3ntm2mUnlq3OtqmFlul
duCIH+y8W7MwsPZXCMntH2W2t1YQbl8zNeSPAwMqIYYO4MUNDgIEXhuHILLKMn6pDGx0PmiGagEe
LIhNyyJkI+lW52D1YeEdY1O4153MoBWY7KoTpYI99u2NZzr8m9khB8mH449mgHYpJKuEfOoFYg/T
1BnVLF1ab2mYZr422sgT7EKw9avSZxx8ZPod+hYkWqM9n+kriK57ZjRBHYmLs0zoq6mQ8aC/uDdW
BMMCIfd6gqdrUkL/xrFPaqwCOIFAzi15zwwVkjtJWMRTlCIOgfUbug/cMGYtw7efsz731BfzH4YI
rlSVwtEmqnsNiPDGH/jlYN2iExeg9MttpyZ08m30ZaUy1W7JhslZr2HDb+63x5+221A1+Orj8xu6
PVSEqBpZzXyy492JgniOlL0U3XbONkhlBOgntEd6QjlsQfI58VNF2W62FB+jIsNTT/l6FKOpbXnW
TzoGxVSRT7KX6xrEnTG27kWs9TLsiKliue/L/2CV95h/5R5DSlYarlnz7MUp8NfnGDGus7NjJ/pu
ybiPA/hd6NlDUoj+ZzXYGKInEII088tUef0KU1/G50JBmtbtPkfZ/Ax0CmpfCpEpFGhaEJcNMaTF
6GdNEeqVadQvTlYfvtzsNTa6gFwCiteQ5XPjFbuEYoZC/n5tGJ6NXLZ0uk4x0HPKSixfQSongOtb
nQHR1kdB6yoVXywaLYayDaKMHtBNMPgcHg9xo2Sqm3sZAg2BH0Ih1yvEWNFDM/ukfQbxEsw7TI+M
rklU1l27fX8t7W4soxHmfZQYZe64XnkVQ4KFVJpg6cjHgD9XEV4RZfli2GUSSB4U+xfp3HAb4lop
+w5XqXeVsTqkjZimSoItq343RtQi65h2xXopkB7cF6lVh8UTpLWoXf8iAgf98hRma8YNlxWyfyP1
VLZfU0WrdytUAOpo+awP+R6kJBc1ZH2Rom4hEM2o1OQorVmkaBfV4iD/afb6KTPHoA8wZNDg1uWC
32xq0KH+KkSpMjSSKXN3EemBWFVeSdVj9GuVpI5RgXyEEMuas1zDUrqcROuk1FrqFk+RfAwXtPb8
Z1xpMoHZ3XphknimbaAx5nG3/6y9LXjR37XITFcFGfOA5LA8ogMKTMH0p3280aElRuO6hqXEONsS
N/rQnB+WMH+xnj0qn7zd2LcpDtKwigqdfFShLux7TS1VElaSFRIJC+KTk1xocs4hwb3mBHo5iYf/
AKQTm3v0U5+S5d7s5Ysa2tou6if0p9sSSHx9SsEeA7V7hMwa8x4FD/5u0PtXh6yQdsMlhuP1Uy1K
k4IFnZQOmp1eQi3v0/1Vg/uwLWUS8Mr3ktUGAQR9MAllPYz8/PCSfbhPTF1T2LyEn5FqnDpF+Z5z
kFggqET90E1daJ67hWAqsp/GLG/jFf2sraSJ7AOD0jYTIT18wxXw9EoDisqrA9cnSN3xrzs5MTg2
TXa0H69zJ3Gaj6c/hjOLQHVlNx8CzMqV+3PIiVYuipzBuKcOHtCNH8AsPE65mKhwmgbArQhOGK9N
D87YD9yFTk21TffKKjlinQvaHzWMkxrk+ygMAXmz4vV2obmyR8zMkd7P2I9I5OTdq6eAqBahCCQ5
uehiVWztW0bJBbfF0yqwKDAggxS6E9GsX3cZuqEoXU3N7Rj/sRdqBxT1esUCHBEag+YGGIj7yJqw
118+hehQNseE/22GOcorOSi8ZqBx2xwRQJGcZlieLP+4fwvgIZaK6t3VMt2t5EMsOCogYZz/ZPZl
cL1W3ikXEIgKcLp8KX+kGD057+EzJPyUe4L+3BGZrxivZsT3xWI+WO9lzCUtcN/ZyI5aYM5SS7CI
SirITOrvyonw4iREX2NTRywGcWo/+K9CXB58sQIzl5MGfxQQaV++fuE8h/KgYRg7qW2TwXELYrro
BSiTUIdkEgW0pZVTc2kfFOABHRhb0osouZGWI7fXB7ANTpumpzQHnCzldPKngUnVl4rN4Tyo7B9x
tx1mUvWP4FvmxBIK3+s6jeuGvHiykwPE5YJZ1IVVSBwh+JoJh08YxyxTAFtAOpd9rTyfYwwfROHf
wUt7lEaBR/NPDeXIYnoY1d6gwnU6yf4sBMTUcqBWvVDHxaXLnnGUXLiHkCFzBbYQG6F6z7jo7DXJ
g7ozcdh1qGbUWp/mTIvWMeTKyWD/vY1U8NogW+yH6Osfqa6oLrUhaNhWIC/83kv3VTuyIouxHltm
3BTnBR1d7EUGYoapDvtamnjdOucC+n4xHUgZmQ+DljBp8Gj6dovWmllnGjUK0H3t7AnJO4MLjmZ3
dKO0dojY2UmNBmK4T6LB8v5ikqsdKp3sQoMQ9KbsGBYLpE1jh0FLUdQo8HwQwSxxsinBNdq5g9/R
24gIFgl4Xee6LehtsDepJMme0b7Qzxtpg0+ofoIVrll9gNUcNdCebaup6JF9FVNV/I2f6tnuVFJB
vpKCcPGFBxV3aGjU5pjmvTgZAC+Wj91SQIXg8Vfl7JGeBtc/VgaBiOKixSAWtkBvgi/Qd6cYCmZA
Fuuyq0Mp0Gqji0TpL6XYIjU3d1NzwKOOsXmIzS7Ayrug9w51Dg70Yov3mdkvqJzuDnhCVLJxcqkl
liMF2XxOtMPdkjMHwoSo3bMNKgjWq02XxN5Jd734BtMdBDp6hUxzfscNXWV+3NApFouHclhP/4Ei
skMguQw9qjP1BInO4TGTFVp209Rm8KD2Z44+ZY/ODy0YXgtsYMA6xEg6y4VMfPXDEKjjJhdRGIq/
vpgT24T+smtPTheTgqAx8mXMDm8FjX1wNYo5NEQtw4rmsiX2FkWgo5waXApDOGrUQ5RkcFicwVMP
qfD/0xN9neZwJgIuokO/DL9c7RTRjsBgR7qDg6hn5tLwkpr3lhDuDFhYV/b1p6kVBJYPIjArPQgZ
mP9Zojx2ly2JOQtgqoBO38k/Z+dcaxTHDCouMEhorvLXjXHp4nQpgjTb1SkYwg18L49gOl4NFIMa
uHZfv0V6BQrzRG9IIysGDOzyb4wHfcoFYRXx0S1OPO3jql/7zwBnDrmDrL3NYg2uvK0iymzH+zyT
r2L77rx/DxDiBNTYV1qc/fN3yIyC8ATWMdiajNqQfOXLxhLnGRyTxXfx2Fo0/VbIcL7wmvDb7Fw6
uhKgumzRbNmFY9tDVMzi7xtEyDVMUNGYjZCTl4r4TcV7rEoK534C4BWuc+BocFdhCfrH+JyOdMQa
CiG0DYrO6qnVVZbPXEYfI3dvLJtGwnNQpRms3Fapbx2Lk4yPPjZ8gmTopyz1OVsl2SO1W5sNbkkj
N/5Rvhk3hhUeRhjhVzT+YwvNfAfsnaXfxGMNTwRw2+rUrsQs3LlCqei31tEH7QQaEw9a1/eus/Ny
DgT9DW7lRCWrl3WdR+0AiSBScuGOu1VENUhUJ7WxXIXWGOpwj1CjN34QMY2aCeok4zfLF1nMs6Zv
Adkiki7y+rsZCw51FlUt8oYU+wJZPcIojOtPLmBiR7atfe3nJhP1vN80OHjlGGDZGmKf8C1xqpkc
HCjHDVsrVCY/7KitOM8jfoWRaOyEXEaDUcSkFXZirT6WRJrHwx7Xgd2j3Y7qOEcVhllVLWLvqOoF
XVUsKKPdBuOkpN/aiHFjhfqQY/c9sizSW/Us3eBjqGUab4YkcmaPJhlLUtIKRTNKmjLd2tAROD1o
0LI/Odo7eE2bK8F+EONZLi9BzYe7AsdMhlFTTGmoRhlUdaojPwSKuLhDa3+tcdlL0CZCI/KrAdf8
OqqaLjBdZ9/fFgHFZyeOsa2x85mQurkxH6q7H0avMfLnOeIze6m/jfo2vg2Qd+R7CTU62B2ZKWl+
gh2NfWSCZr+Aflp2e+dj1kg7gyI4j7EzMAZE+1EUeyuSkf9U5T9wwZdPhJ9Qcz5jhxYfWAPIYrVv
0PMWW+a3M7OZjo7BDrRRx0V4Si8v8JE8L7Vv8pTGzM+++6ufXfPSklHajxrRA4Pn4rg+t4amOUL3
oW8AKJP87+7uErjZVtqH+1zIZjHnA+nZu73PdcL6+nh1xw5/aD4w8p92ZkkhRRqrKmDIPfpcMfXQ
gZj5S7kLHK2AMLmpKlFEpSi7+vaFpIxWzNVJPe+3/jubm6ZWNBiuyoa0Goe4YxlS6acsNPvURchn
gwLoq99+9FxCOjCJ5PJsazUpmnrR909VLC3EJ+qXNHzuodwxzp61IuWTcC5UBm3lO2D1zStNW5yO
wpgey5trf/D86XS5bwPtXndmUL9o+7brOPSRRUqJzVHN0wBRGP6qMFFX3dwHFo6x+dpSnxaVPk7s
T3vAVDkuzem4ZWNQVH/i4iarDLUxI6UENXtAaqfoQRTaOGoSz29p7UdKN04rMCiWVdlA/SamLbJX
XVK/0Id9LgBrQEYV4FkfSO1btIw/NJFYDlrsDeKumbz9MPCOgSzpvHwm+aELGUIMq4bmoFy0LTCT
X4fyxkQLmBA33kuHIcWRd4r1RWGGXKZdv1wiZJJnpVxwV9bvmfpoqf96Yxdm+DZZavJ4qfxc6Igo
0cvliAAfRpPlsHXTfhP7tGXCtg/q27znOEbuPw8tcqoWwmWkLmr15j8R+LvyIVzO9DpeJ+I+Y4Vi
niFLB+/6MJ6VR2V6jA9cklM9aadk23wdcbF3KpKp5huDKUJE3PMqAFsuy3NcDJ0PyjaC5UIo0IsW
XarHw1rkW5piG3GMiykA8oNshZRcc6bqpadf2c667KtYVaHB1TJ2B41b8j0/K3Juy48mUzmNtWb8
L4RQQhP+nOIYeFMyR0RGleRmWKenZp9QoPNPxPtD3bPf583eKHj9Cna4HcqJOBF1oLDz6Bw5w6Ma
086liYPZiz1kUmPiESOl95bh7pIB5LHmZe7GNS/eeqgrJxajMTXTt4MJbaUjZ8RFA5Rvvmwfu4tT
0H/QdVp98O00bhyrpLB9W1KFvFV30TTW4MSoeL+my+BlY9HH7pQ1xPVozWn5eCWvjkOWUgvWQ+rm
/NY7Eygp1qCAbNOtQ8hLdtUYbjJdcjKyDGSVC7iTCDATGZNXU4r85k4qeO6MAThYOJ8dZiIoVFmi
uKaQUd2zo64K2GLKwWP5M5MtkEtIuRVwqwcB0SCRVU3vdjH9hVR7flZTzoiq+k744JnH1Sme52oR
Fu4YqHWU9ZxIrDmWmuY+8D3a+WxxtH8bieV1tPTgT79UC3+qpOUjgwxhlmNLDoHb6rjgjsYaVeHj
D2Lzpl+cp+NvoopmqqZNgnnPXdo+KnNv04vsrpeNRttzQp/m5rOKwvIbTqwF/a75X+UnfRrvnGGL
7NQFBFXZMD6XszTuOW3fEcY2SWAfNGNAU9dRVmgVoMe84X/JHlsg12DP/GdGyJaJpT/K+qaAxn5s
xaRd0cosBT/RZngPg4Gk6CeKtw+EZsAyl0YyTIlSZbjGUfVo0GN11WdZCGTlMZSqNwVOxlwY/zUm
caYpxFf9TP/Kc1wa2v3WXuIhBRiMjL1wcXv/9pfNjRPnndR2Y+GFn1sDC4McQk+oFV2VMmN/XQwa
MZfNkaTRaRdlZNrMFvnD6bHM1y7GT1lAvqnAm0cpcCh4ZxB+z6gVCz/H0JD2h5bCmVrftkDgMkxX
H5y2AWZP0LtMEFanIG+GU/O1vA/2v2mlpNHFw+VDDs7pSZlcNgAAHEUdMp1QRMHBuNbbIp5y/ERZ
tSvL7mI05xp5JhPvibp7sXw2sNGZNOjYylX0fJn7MKy709Sr/6NRhCcvywOch96ne5hCGugoLcZk
kenj8PBOBQ7cUekqiybH20n+MWk7AJ1pDXm7JkbQsq6wOg5EyqJjuPUSA7ypvYJWpIbgO5puZK/t
gXYkNMnUIbmUnvTA3rx/hA9vmNgelKtftpp1Qpj3xZyzm/7cOeYToZbOGw6PruqAnEvKdH25aRCx
5OIcSfZ1tsrz2uowpziYUUxmVuUd2nAF6TcJUuvQaqrdsfxJl2ly3p+l7bZVywZq3ptYddAjDQur
LICEb9OiVUj7taigePZ/gjMfN4nDXjVJA5UFMiPA1GWtuvgnpJxV/txHkUT4ghMhMaPGyz46GszX
kMFbLwq2H9kpohldgGlUkMhe8DxYNHSoFbXl9aDbjHoz3pKj9eWvT6394z/iBgOAzXM11vwZd4Ur
WOq605cKRCnu6jjCKhRNj9MZ2vP086tC/LXgO6aaQGcunRDlPhRpUypRk+aS7YCgFyrvmWSvWNAO
ScVkCPiwxsMM36Zp/i2eCv5LjhWwgnp0+YRtiKry/JfM5JS8Ai0j3Bve6ExnOixPbVF9MHIE8SC9
ldVLj0ZdrRqI+q0DFZd4hcCZFS6BuiWMfg08to9drXYpcjiSEriSw8JGMVBAqjOZSjPTy0XvldEJ
suFJBj9zCB6/ottrOZ8qujJ9xNGytpFk17QlOSJIH+JJZG0WF5WX+q1h18ys+OUro59kmLyUikUh
lQ5IZlspjB9dKTkk2IalSgMLBc0JuMq7wQ6W+ziGvp3zFC6/r2fgv+pEupBEjFHfEYsExaNytN3+
eGLwgawMszV+4bHUc2K9tFp9CWlyioFcbYnbHQZR23fgxFdSPCRffaGv3DECjQQBghFuLbWjW+ic
tLwoJIa7KyQqHAxcy3UPH8nyasZgM2urwMutkIBNjN2Uu1l5RwvFnAE30jT0OzJMRot6tnKZqp7p
ONyhjQx3BQ8K81W4pJ21pNgzSL6pHpSsmcjVPMjlqmVCTg2Kk2eVSeR28uZ3/VCzruJ0pBWwTPiy
pZZJDCxFCuiDYw/CxV+t3bIxa3mbwzz5rA51rTr8FC5xyFjkw58sfjBUYQH+G4b0yiL07+/U2ZXu
dCplwXOuHWNxB5BAMXlus/0myRQ8aW7d4ASkNZil7UL1R0BaAxzNDSdxrgRym022ODdAp8gNZoXe
Kk0vdLygkClOqinaYllsEhPuiSrvisVhRiq8Fi8/EQyYUEgGwN7TNX+8098WjnoHcrQEuJCnrX1R
I1Cn1RIEqK8WBx8pPY58zPBZPfPvEwElHR5lhc8Vm+annX49TLxG4JRJ2Ynno1pIGqxOyuNNVL+y
DVJNUjwxfOwQGXDiUXwdQi3fqx3wESYe8v6eX3iRZaHvFcIS85FrPlC5K93pA3Ia99j0HzS+WBdb
0Tg11lp5K5CuZX07K8k24F4u+83cEtndmIyF7AjP7zH9Y+EH7sKOpFQSQFuQNCYjd6kv1U7lwhVN
/bf20OchGyiDb59ZCUMWq+0vcVTx+M0s+b3WUldAxI2lrIRTPu+RFvGvBN226QgrsXc8v2ckf9p2
Q6kMjW3wX8NVqLVA7aWCGJEf3UqO7e7vajvm4RLgLsT+2iN8mRvEDBmAzTqScYxTqSODAubr6x4Y
K8JXxHlqp4R9q1eAGTbtsPYXyKAchgjodth4PJYtP65epY5w9X7nqn1Z7TCtweeT8dmUx60NO6VF
siCKErpJzI6S7mKn0BrjkdSwerToOqkiUWALikMR1Sg4gUX+a5tyOnaGfk6HHCEltoHlmFq8u0aG
ccpUNH1cz3id+qJp3LHVDv9m+kNH/nVlrghwJdfKB1UMwq6FVOs2d4t6ScKURDfHEazxbqupmhA6
Q+2yzJmygFCpk6sfi4hOqjwFDFoUINNZJ1Rf9rwmzsFCWk/RyltsvKEzbo4i8Oo3Dqiws7Kgwvuz
gIUJsEsOqwPBjsmpbrXG6AS15G+MsCmQCJvkxYFJnPtcYrYlJZq2qSEaAnrvpZEhOIRs9Ej6W3Sw
UueyFx9EFI4Ry2rtb2VcAS/10OGueLs79WrwZsBceBj/zmzpvnCGwyw4/aK9CEoN9UlgH5ULoKSA
Riv5yYqHX8RFtHUzR63vcBCHLQH6VGmIRZncfejltpvzi3rEzTDhATnjJc+7ToAQgtk6m04O6xVX
4JeXuYc+A4jJ58d2t0NxJaQmSsT8EsfZSgFVKCB9t+g/9hKmHsTSuzrSblzTkiOcRqfsL+2EOLuQ
RcxtGp95R3soP+vEeQkvPqcg0QSDbjqkWA42Xd3vTIxADJtRaP9kCKnmHX7bR/SwB9O5pTQ1hqdj
/FRoidoDn3nN3jmjJuqIZQyrBPdWs4p/++e8VL2EsLxfjQDJaoEr5WBpZ1/9SvHORdn3+7UFEtCm
2kzwDed6hkSEQ87+jgtWyiSp7mzscu4iWuWfiLqDnm8N+n3VVLoPYwiuKBxDdWQi75IiiSygTpRb
nNMcvKaqGmtcRSaOYCX/MptxpHktN/2RIMI5k9Gg5TzXFZQIngMQsa3S8sR2YYduimhh2SSYvB5w
l/kXQIYI3sgr7ujwEfr29Cr1m8CuBz0RY40Mbfq1s5w/tRBtUC98924dXAjA2t5UMPJSYdzxKODU
gRTB4lAK9XS3STbrgfleWL2WBYLlAiZtKjmX7ivm3xbZSGzscEGo5AqvZQjVTpA/Xdk1b2DoWlN6
De/f+ik6UlRB2mbLQuehOwsB7HcodlxAwoBLbrw1w7sIH2EafQ1Wl6lSddGfbixz1doDPv7M8pwn
hApNkfSo/yxR+45d9aeF/9xVhKzXL11OxMx8m0lsBRwgfNg8ERPnLNrvZuXdVTbIJ+uUEsH22lSa
0Uc2KcSJo9bbhtn5AVOvOI9GJZ4iaUWgzh2QGgIWYA11EJvcZxTVYu7MBtSPZ3ukfCx2OtMZGL6p
GM5ZdVt8KE7g1hCHoEbDtL1nUiSleclc0Md7IA4QJ7iN3SJGpiblNYgSqG/kh6ocQtQDZkNUNce0
FxwgLwzIY/b8HzPGw62/4YOBXmwMchwyftGU0noI8hNK3wgrnMYHtvNYPCeJPpoXKRnY4fu9vufH
+3DOTasxiQqK18DL3l+93YZ2CxddEZWl6rRC8+gX4jL4qNeV6mCqfwHCj3XI0ftGYGws4BcpOD+o
FHIa+lAouGjZvNRPQOYh5YFRRVkUF3/FFklxuZP/foN7KtfIn/AbMbFm6oH99zgtkK1SlmSII5HS
rSo7BbbJVjpCyzdvpvUFzQ52ZhLgxaVFqWEvMkjd02ssroyQih43L7cpgtRp99Iy6FLuOCvvULer
9bUxAjyfVIXNEJUXrPchSiN8tCIhCIjrptQbgXDHhYaYAIXpozU/TIY/9JQkXqd6VBIV1YTEAqF6
dN0ZGo5JQbQkjATE55ib0tUQU3B9K4Ua0quANvCDwcBhJdYFDeZnE2X2VCVl+GMtmlqTpD8FJJeM
P0pHdXGwXVVmppfB3prgQ7ZyrrOrztWZ3/hKIrbAAvQ9ElUx+do1mhjq0I8raV0FuLWMGa/bKES6
mypQapTkpEf7zzqKv/PNMxL6Q1TZPzDjJd0kSkVSqNnGuvdXfCZcSu4atLqhdH587lwK04jw1OvX
uHm+vRgTwSTeSpHjpNPyfHK9ZPeD6uFLE+YJ2R+ni9cTXXFH06DZf+P1WJupP1XSUxrGZXoYcsIc
lOz7va9JTGMf8PsOsmE7ljuk01tsRBo8zY3D7Wh8FT6+o/88+FlSPyMEWFZc18cCHBjp3ThqCX0D
YM7Zuy6KvSP+FQPQ1Ss/cBtWsCdJ7x2jx9zZZFgWwV2waDHlq8N1NECdo3kJNl8+cLnQdyOp47MB
enau1458j7HgXAtJJdHxaS3eIidhKaTAD4zkG6xLEJkR6S+NzuZb/38Fnpccl+w+JhL0VijO9g0o
965GDkoiEMpikuDlRWffAgY38GzTA97oLPe4TMfp4pI2X93MoJxhSMVuGq2pU02mxAG3iQwWmzC1
9vRwMHTLmcyg6WuMSURHO5rva4bcDmyKZ7MqIU8voE8lNkIZcSDlQ4moUQHxgr+OamboVHPEBQCN
lqfJ4+hCO/bHfYimf2ik9sVXdu+yiQUfH4l0YVOJx6pko3QDfTBh1tZz2leF/cOHeGervuKhcQFI
80SB+WkdU7TufwsQ5VfyGeSqU5zoq/WnoLb9FxloSlW8jD1491TfkvgFKp743oDkGzglunGfBUvC
DUJYwjtkyZYogVRCSGhAspy5XXrofSODSfNGyGdWlaqB/Vs0iTbYQNPWuMRWds9gQMXzZ/MZEmuv
i68v1oyKCbWxLuUtkB1KJiMlsziPH2njd7Lc6d+OXtAPggzL306qxwvlNXp5xZ/g8D+zY7xIQjrq
zm5e1rVXSOoF5giQEDne6Fi52URwkczIba2AsbzZSFfy63brYaWe1rGVhqd3rrUPkaMhDi+U038f
5oaZ4m1XBA9HL3uh391PJ4wVYx6zgBqE38Y9s8/dWtC0/eIPn0r6FZPKvmTboGlRE8Md+IrdyHXf
q5cQF312Mv4KMzzvDYL23Bi88LwxCbiofIZeN0FUsCtMcu9hxcX5uwQsXzjInP/bAKv5rWZhoBt6
HL67sz+jCwYZ8VYavb9mlGXpdqVibb/avISlQNfhFG+ST25+qUAGTfvFaqxO+evaLUUcrcecyY/6
ZBBTpU59ufEk2CRabMdEv05VlLb4dQDpsnHDaosMSn7VTpsxmRs6UQlE79IWRCWyB/w+SMEJ10LV
DuObtfUpRa4QtSzyFhP0+UhNlXpUsz1dZp9GJzPapFFv0E0uCm3MgCIMX+MLs/67A+2y92NELN96
jCoptid1A0U/4oNxmSt1ZKVwegx3Lx4Vyth48GQBeyebZ7753XpP1FEuhBtk9ULVpCYimNuKwCtn
MKJHOdMEVHi0sc4ZuCwNpudyfHpda3spFkgC8l8fet0t3/UNM+UoFNfDkDDX6RR+If9XLXqbBqVM
UefWK1pF1ZBGqPBYyA4eyiZagXnXFlcJ+XRGvk/P9XPILX/NOkF6l0XVRHCHjwtoSlRyPxaWzDl0
qufKDzLYevH9GU6e1coNesFNOyDSep6v3wS5XFNMolUTW6EyYcjIPzIgPjfb9wyEtTRp3XTFw0IQ
TbBsQ7eBQeNY+Hi+VoId4r45GJ+hlbKThTfpbfrD02xayyvfXX1i8zGreuLDAHIGNuyCZzcPdJKj
P+g9zI6H+CpLQOoVkXHgzKJo5zZgylK0LXyRf92YXkQQyzXsxzL/lDrkYop7lyqFdtsQaWvYFmZm
j0KtncG0ijjoKGk69srkjzXy9HKZp4ejV7psUftCXw6ODsZAEno/BsbqtVrck7VqiZsdKSYEQgJx
wLYGWc2Q4wVs1LmD23DpECMgqBtWNa/diCesF3i859Ou0xoUGCvQpDnfRwa85nin75prJ8+mF5u4
FATsvOSS6cSlANym7q8e39kHSuCdy9tkpvFz764TusGvg9r1x3ldBw9/Lx2yI7thAkUBytVULgzm
Rk25ALPIG1+GaE4WuJdqp5866KhAqRmhKe1rYqbFwaYuqQRd6pjROYKRHAI1ETyzVYl2LIBQyMWe
8fgQCJxy0XDpq31y8WZ5ijWJnfinzDB2ndm0xL/atnDwwxymwru82ht1Rd36zZz35bT1RrXtXmDo
AQ306hlVPDG0AJRlHTm5K52BkqZFXSDzNtUq7lhKA6ajw0ciN5l2g4E/H0/6lSQtaViSkxNTed2R
KcJueCf2B/NKxUY/LCzpI38wKPK69jtNcFcqG2/y+rIpTpKXSOgSHVDNtXfhqZVIH9YfxYdIpgJ3
03EBimPucnowITx1dxKOCD3y3RLBZnhnEHkrnp9Roxpk/RU6M51c8iEHFF5tdgERYLHTx8y+uooj
9NMP/7G0ClYmgeIw7OS3MXhwZ1DB+giMegPUaDL40l+JNMaiy72a2iINuC9HV5jZzHQ1Q2m3NeAu
8ed3wA8AeZwGyoc0g3fKJ8PjpP/+CVtsB+jIkLbrb39svRFaB7QH5RehCnluFrnp+RgREcMU7ZeG
aYvPRDmJAG6nY1qggPIRBOUxUh/OF0g5kD4SLBlVVTV4fWr2wOUMkwtry7z6/aBmS9nm5j0SkxaM
gzVv2UsQ6EiR5O+sOFe8wMHqp3K1pg64TUeHrHaj1NuLAAg/hJ6HVm7FVjsl7jutKu5qexIY8Ro0
waWM6tg7SbcdBj12F/YX6LdhPQBFPrjmo2yIO68WARi/gEau493FYcPMSn38CtdDDz8VFNlfv+5G
0drCJFhuZyG7yCKTG7ATaOYhZD+Toycsb3FNxc0y3NGmcpHuBk+4aoOjuDR6LQvZcby5Pp+yFF6z
+maSoWC9rMxUFC6AOCjqbiM9VVr3kiG+8n/JlwzOQPrNRJT7TR0/9xFtlYc6uwwZ0Hz2aR46h8yF
rwzIqQw+m+VDst3WPJGAnL/77rIU/qNfgRE8NK28Z4fvujWtzYKgVGsjGo/g+/ps7FdNZ8Mof5Gq
TpfcTX8HG1yDRdOXea+lpWaiBtcbZeJWC00GtOE5zcTnlChO5C10wZQ8JL5E5c9ik+7GCoQlusy2
kzbVG9NDW49prxwNRQGP+DfPYLqfLRmJliYh60R30sl/zoe+e6vI3y4SKTI9cM71j4SLrlGnkkTm
i/B9Eea6wK6ltswkBHXFOUJxZ0OdGPluW8MVNheZFa7JIaW1drwbAqSBRq8cYMCac+L4pT7qRaiH
CSifb+sOjlDMEA6yinUT14WOnNvc3sUdy5Z5WJDJmPMxNuCPpvPJw2VSGAJoR5jivT3nhU8s+5su
SQEVE8FbskWYnF3m0S+MhNOWdSMnJU3Lx9rtByt1hGOakRhzOaLdlcKMH+Io8jYXSoCgwbPPooWg
RJyV3e6iaeLXy+jks2wQ7N9wyamNRvyvr16dozpBOrnxO4zjU0dmd9OinuqUgXy5/IVcr2ddkSVK
pkXy9rkIF4AwzWW5+uuh/0A21c1cQCkAUy8WetupzqZIyDKOPsciGiujE+ktvpCc5f5HYUPjiMJd
iSCcLtcLadNFb3H8EhI9T8ODojeu8O+sEPcEf24bPCfnjRGexFMol6nmC68xXkh+raYNW0tajnB2
VPT4uM/f02r+1W/yxtAgBvOUn1kU600bcMKK+yC98bQys5pmJFya3Ln7neaIFxSNf+N+9AIvcqTe
aMMPiOZK4Id+dQpkY8e7aYEyzJDA42Bd1+AFgYlAW51fZMlriWSeSgNs9bicgFytbzvsWFmXQ2kU
+3m4COGY3CFvuDwIkZq0Trp739cB63KD7JKVTrXoLalRvcVTfToaFuc9ThooZW/aKAWDXwPIoGYp
VNMSfJrr86AwhXHkU1UjQxPqGJNq1WN72H1GipPZKydx6Eri02ooavcmcT0UzsVzt0BiQXnGFfZu
6hEzk98d0SJBIgi+/l7n87EcOPjlGVfQFKeLV8ZR9MMnv3FXtvQGJUBozoTFmrwcJSHgPPa13aEj
XR1FwZBjCEJpu/nRO2CFw+utWwblWYiXCStXoUhpX4v2c6dHa8+BjC6Eh03os2Dd5biS7zZo01PW
04txdXEkrBJROv6dGSO/fcU7ySMwL2pTS+CuRj93pZcbxvc15+WHB4OwbikFx2qQDuP+84eJhN3v
bByCR3AntAI8WHU81cdKkMY2ypyEbD2A1bW5m3fFpwIinwGZWrIOBRpwqtGdz4LTTWdrags9B8VJ
Ip63KJX4tthS4uE2D1/aWsb/zG1NiBtu2ujzp6ogBwEiFQhZqZnLkEkr/CATT2KJS5Jcj2B+0KnZ
Tel9moClDdZ6NZ/uRQI5CImN+f7g0JIAzLisPuN0HV00KJJ2mgOMamGAbBIbsPtpPk1+BA7hSHwf
RkH7+AqMhz2fTXt09r3VjqTKS/bdyc2vnVCHpCU1vwAvW0mAjOTqtwW8EHK+Ya8gC94Y065fK7oD
mGkyUFn4AWrnRM2r1UHFvG7Ise8BDSEk5D2ZCw6bGWQDQf3SZZvDgJkAaav4nbAFHLGcbmvDpCah
7vqsenMFwbiwiZiZQCaWygYlW7rsvRRDMZmFjErW74aVmzxcrzSjNUudSNz2sfsuGOoUZlzFknZZ
o/BWGKTovg9i5wN92WWOvCG12ZEptUrePsAJTL/QN5ksJPOOk3uV9nWfurm9OilNSGVH9Q/AcWtU
8Ck4of0y9bi++fFxrZUQbTA1/QAWUdmjhyWrCBwA8aO4HfC7c6rYCxxFg3i0pY0604nheSqIWolb
cwQ14vRBs33w81RT0JTS1fc3jOobEgI2Cxy7eOwgv2XGHISc4vu/nuSb/zTRlgX4MvQkgHJducxQ
zIjvvfNnNaAD/ehx7rNVN7+5ah3FucM004OhBqS9xAIBTBdaCneg+WXAf/o/6fGm8oXHtCeUJR1+
ySjASnEejbMo8vKODPylDbu5I+vRIgpcI+8h/tQ2eKtjNhkaMkJHdHxKVePVFFUQ7Inpt9f5pydx
4wlLfKjuJgokPCjXl1o/H9X/aAIratXSwbvNfHiiU9tdHB4oc60GmWuY3EDywjQhutlXAKuy2vIx
lHcvUumXvgCpTnxdg0sc9eJmVN6gSvA5fw8EPtMwDyL1OPHPT9jH97IGRUxe6V6vossLY6b9AhYD
MTOKUcbUHI7vGWW5CNcxB7+RfMX/aeGJxVcm197BOtaYuLS7ovxXK9NHSfy9cyGcTROZrnfvfhOh
/9j/YVv9f49+WGAoaElXs6DmjByU2nsIMN9ns24XnN/EV8F2B4ZGzD7cUVmceRKxoKX8Ul4M1zRC
EXK8/PjwFuZ1E1c9Zs64mX5czSWS25Njjde2ZvPrcA+icOq3K7GoUat3f1D7WeLcitQHHn+HrJaO
FySObgOPdkd57Z9c2IaKw8UZUUX3HepvGNxKI3WB8kr99EFOyuKoyJIqGil1fNEHi6UOoK6SrkrG
/ih/cDmszuZKbljriMJYJSSpzn+pXgN7YlZ7HQxYION8T5TG/dYsiIHBCZ8h8QuiofFNXgv7CQ1R
x8nQBPPH6dh3vVdl4OyBeLO79p3Yh/HX6SVtHzmSRBpv/JJXu6eHMXGeoQPg3Yqp1iG85OxpHipZ
HstEU0sb/GthL54sUO/vTvalofdEI8DxZcgnGppAVHJcrhEuV/dTRenYQ0rQV2rZvqd0k64wgtei
/i53+YJCTROgzJA8IGg6U4tkO60DtPcZlfbJbPgq+KvhTCKGT/Bb5Cz096Dr2zK3dFQFiYkloXxt
Y1geOKNApC4ouv4u3G+VBqQKduANtykYl1Wtdr9eNQb1HC+pDeEn6rDBetrfC3QC2YB9wjlNZddb
0FxGu1tanfbvrkLlxgsqncC1DAUOSzHHlBRGjSrAFpaxHP4FYmzuVCYO+tQrnYDxrm+XoaKtOleT
Mk/8/c+r3d6yMg5wgRcTBHhuE2O7p0FjOzilh8PmCoS0lyzSm2gCyKVMvzYmMfxaREbn2PbEwmu1
8tewNHqxPIUYW23Yyy7MGLMXTfigPYE+tHl06GV3bJ0CQ7FUmvUUEB8Al7DWIKbevAGzzQ1xGD6y
OMcJWMZslbY1kmnZp0ru01mHKTBTqrcXwtvmhFS8HzOCPnDulNUgTfTO7CDUvOvMsSKju8kZzal4
9XM5AYxgnCY8YFPZHcF9rSYchlD1NRSZ3GKwG3xhg1gzbiA2u4cbQEMjPkuutknhdMy7gVUHeXVS
n8I8Z38MCRCUK8X99WXaoY2zwdRs9YBmi8Rem3Ukdp4X1I35VuSoZ/hrr4l4fCmCQy4amAHhvPX8
HlHSS3C1Eg+qtsJEQpkQ29dzMHEiuWbZNZH3VVVZ4ckUC6hFLUKiSED4wI4MfSsAjreU9rSX24bq
52RVooQ2Yt36RE5tKhbjLP0oyc0UDI8e9O09ZLzYhM1m1hJU7HV4RU8uPYoNMY/q69U3lRo3lBx3
gwmHLYcOOMOojORDKE5xzI2tXWlfkfNgswSKkOpoYFf1v6t6h/6XNlAEQ1oI6e/uL5UQkFBxd7wh
XlNKO7B69zghj+NDaMUKODMXZZA5iEI2FfisUOHT+e7Gx1h3vJvB2VvQKOIfVrhvCXXrQKItbOpg
XTraWIFcdeqxqpAWaDFIOzvhRzbVeFZQh/oVAzw6IBpNkinjALa3fl10UsMHGZsU6YaSbCkMFKw3
r7INLm3LQzQ1tPGrTkYKKA/v4RSL4Nq/AfstcIS16PmUhF7B9gPI05tsukFsLRg4so7icPv6LjHi
Rm4pTLowcw1xACuJUTX+NjpBuwpbYYE1u8BTvDG3t4dLyjpLksApozjEteAGNoc9LY9582g9f0+c
bCP2ZUR1mfJ7Ldr+eC/7c44ysc9JtcBsHCXjHLJnnaWvN+V8aW8gQ9QtKbmEbfYdf7QSKdB8zvXf
DSJdtgSJOQGPwl5uFrohABlBz9tCyDUU6iPzkB4d7c9ieqvSU36e7xJAUXq6HuCiUshzJcfC+Dpf
SeRoIeGlQhjEQRcEyzBIOlCHnK6Stm7cXaqSWjhOjIYZU5EtxowXIBpk97AVYpmSVtAAPNg1p7z0
++rc292Bk1BshctXPc2v0w8uuLJAMLEDt9mPxSM8Kk/NgjEh/eNaIX6pXNJkqYcMiqloE4oMJDX9
DKKVmmUHEjBS8WslmTVatWsw0IXSnyOv3E9C11Qq1fKNVLu+jpXE4ZhAm2A1PMVeGhV4iQCzFqjU
abiV0phJm7sK6El2QD97zCTY96l1//LQeD5DxWdBryUrQnOA1Gv9w0BRBgEHhhD+Aq34i4Fi/Tpm
8rifXkwtWwqqYc+wr8Jp0s6a9a+DCAuV0BSij3guEh80ZfNzUdpze3Mx4C+gGVWVivdW7RqW63bF
RN7HrH9af78Zy+8Atu3rlQAX8AxsZkma/D7nWUhOPWO/ahNqM8lILV4tac3egH7A1hZjA9HyYiXw
MWN5mhFHxsTjmIcHgZ1L0t227GQvzceogbvSNqf7jKD67f+al6YZ0w6XY/RbQPpOTQGcGkwDfX2C
pETzN53lmWvb1KorctCCKmFv8t2u9+xXJRFlLvxZAg3Ht4tCZgBU+3B8cNqGZAI9holeM/ioJ9D9
WkagmJAFSEc1h674X176oYzbpSUm6HYGBu+20FZtbj65t+6jk/fhKQ7t3hZHRI2qbtDKPdFZTazV
gO3OOvhJK2ZB8MTg+MqcGLBg8Ml+5rV6Kd8bY8cFL8dxfrm29PcPcgizmoyzDm6Spi6EnV5gL88Y
b61CoGTlzoPcz6Eov3avjBxXfCWItT7CVnV6t+tdN++LzaMN1LdfLNGcr8bRnAXxS9icck9GzydD
H+Mam+zEcMDT+7eO7YyEAWV59Y31MA0mm6VhjlEzFjUltq6GPr9zRSHrACyxJODXhtK/z3Yb5pvC
SWJO6fUR3SySIdMcT+Olgxyry2TgRtCaQQsbEU8SCkJFkko6IrA9YlFJJvOOJYK0lLo/T4M5pWkN
q0vKvb/CVxWxJphkvVI9/5Bu1dKdTdtcu8QHLCfpKC7mK4aN1N8GWkbk3pnhAcGbpIYNEZT3+U4i
jrSvLo4X3X9bNSgv9TBDUYtVjjztudJcRj7zIGKgAatJ8lVNdQmGx0keCimjIeg4aC4+tsISqs3V
OJVvL9uUuawo+i6POR/rj9qN0bIDuTUsxHC6zOTeiiNnwSxcjVIuO81TVMHnMZG+HJlS8Kt/pvzS
v6ebYLzj7jtmWfJxC/x0Zl0fvNeKj/iZ3Wbl5hokJz0Gpfoykq2udPCG2059ougeJe94ahz56jvk
5nMQVlBftMB9ZTTZmbqQqcroIqBqBjIBVHlB/qw+Ai1nRidLUTUlTWp2e486/QATZxC8WrIuSTi/
IeaLLblM4lR1FKpS7owfYBdAmhuSlVwoRGXr4xnE5ThE+zHGgi7wkzB6j1pEGeP3vcJtlwS4mO+F
7ZFxWo+QB1SC/P6A1PNBNnHcms5a5cbr5hNfGqEx8EqRpxK66DlvmSwq2WNT3bnQEA7SRRSMWU6O
XYxFG1EabEXkrBOIlcUOfwffCsLpZU46MRhYXBu1Pn+RJuoMOUmkTyrf9aDNgWs2UtXWk77iz1YY
dwybXohrIXQY/y/+1+AeAUvAy79URHEVfpyZ+NBLSeVsUSRVfHgYm2HqtyMNl09rS3UazNVhWXXH
cqirfyOiPicB+JxUvR+rAhev7t61mNuEBFWIS7xwIgqOIa2s27Nia3gJEyLnivZ/B8pL/OIK5Imr
OTBfJ6+ER+o+uY9wUirUtGw2p7c44iVNwaQND4QdMFIrD6/7ohVCNZFjXKc724mJpR0f9+SpQ5+L
rjOHZofJQUY3dEt1oLN4yvF8M8QNC+ctaGV0X4rKtJHZL9UtftFssTC8+kqXsm2koyFFGPAA6FgU
zfCvW8l5YSmut5FsOm8TUqXuzipVZpS6zcCCMLx2DjDUkPbZQJsE6bJnmWb8bd9G7FY4tWASnHDU
cJqHr00HL/SQq0sUQtbzK6KPOIuPGXDbsbDKJ6jbPOC6OtFTRB5twF38fI7zrcv8xPJeEj+/ldr7
MjEehAqrOqqfJTlP6FSixQJ53Z4261Z8aKAB2WXdtuiW9FAhFWJAFcpwo6SDgZ4r/zsaj50h42WG
vYz8Q6Me26CAQhkMFGiuSGuzW2f50waD5AACO9foYWtByoFheaL9o62QjuLSyrJ0j2Ryy/j2Vsv+
MdLmbYkpANX0d5AViK7gTeTE3AeOxez4h7hH8AWvMNyAM2ImRqlSZeW0XgkwRxw69Zs7UhS3+7xi
6I3vIsXuEYmfvlmz9ZAYZWZ5yYJYape+FZu3gXpn97hMzwzVCbP7NpjuveLeIJTvpPm6KGYIyzgu
XXYesKZCwDsQV7UKV0fV/vgmzov5w+FVTQD1rDv5Hj6supQfQ9wxS1z+IAdUiPo8tPvL0aOD3FY4
Ncn3fQ4y7fWQMKVjuME2LdGtr1OaeoZAWJ1RKPCy37g8/0jFbahpK9B1PgDnKRqdTKFndnTpcLt/
Ff2nhcbNH7tj59/n+8CLAbKq2UMgyPU41Yuy28qIozZpx78WbZrO3NwWqvMW8Pf7H4M+fBOEUP/e
hH7fDN2aqCauqd+vE61lsTqFk6Is/QDPH0TXrOe42jYMw/bUYIGwSFWLImiootkbwiPM5JurTTYp
6TntRzU1BclDAPZU7qmQMu5PktBsAJQKICIMWAaw8XlpNM8/J2n573XtZSKk9btPYXXF0uesv9JN
cV1tefW47jYTpBmOGeLyKBvPJZgZS4iWNljs2xMwW0uQrXTC377WEswB/RXkoNXFYSU8fDQfFOEK
8hWykDhdi5z5RYwuJ3vQmykXvS0F3PjjlMciXoRE6CLAP+q0ajAJPZF8F3dwidGOVlhVa7l/CmCD
yrz/O6pzCMnSftQdQjQdrfn0n5AYzpgHsgPaz0bTopv6rXzd3nz8ieR5UzZ1OyAzZASEKbbjE3ov
bTFnCw/GmzsAhryf/+7tpFONU7IreNzcBrNlDeIDb8oAYM2+EHWx3b/t8ZgkJgrmR5JZYA3uyBeB
2uKzNGc1jlYmsgscZZvz5E6MDR8LqeRD9NGLtAn7G1UqjF2bbejQC4ob637aMJ0VdQ7Mx99afpYp
VKIcHrb2PArjJfLVfB+2rX3E7+BoufDFc6avrkLJQdQA29AT5pWlSscpi8fW9lvqLHDeKnQ5B6lk
3ErMeQO5gOcqMzqyMvVNMOUXtavRLi9sYRZT6/LjaZwAgyiypnsnHAdPVuXv0ldaE2zHAmk0mQW1
dmUIuQaUWWbiO19kKzR7XcAetXLrUQXhPIPqZSOFdRy79AmwjnQ2rbqaFgqb4/vdoMWOvVZ7YT/L
W7dXwv9CjpM4cAW4+XsWU28SKNhwXSlxX207efGAe4MFGSPI4+h+DdEk8+p1a20KRMc4lTurJxqt
ZE1beojigYAGPxJbj+xk+iulb4t1He+fdMbXuxi66qBvY3172xIeryqprpBqFHctUhtUBpU6UmXT
4QW9Ggts9hL8for1P6soRbJYh/m6dYz6LyEl+X+P56T9Z7hJId1/UlJSlaIm5F6lsrMsrAu8EaAF
I1eEexJsijtr19o2OvO929HRHiGMy/nIm2bcxvwNHZ4BIevi5jGYZn+J2Gwl3hOiZxVmmUweaJpZ
4G3YqcOXVS3dqOLIGUpmlRE69EtAeCji4X/jtSkL7KSVZIL/y0alMh8D0ttbmhNiDZJO8IkBsMwo
Sr3J2bZ/jhwnUeqoTsHDHKJKcgM2LNdtEgQwYk1wF8Ya/S9p+jJosBcYtiYn/iguWz01x5E7zhgs
ITFG115C9eE83F+rk/0kXINMAo0AYa7czIAAJ0g5C/BCokDoa1qo7N3/WozuXEOc9p320dVYkSF7
2xsHPKwNsHYtUImSsQzGC+0ZMvBHGJDF35Sr7aVcbQKZJsWthUVX6bN+I4iknLvOvknwSSKTRvtC
7d1+mHiaDrslLx77VYEFs1ANPGhlsULQH/tHTYGTwOAEQaW4rg8BiSvnoa/+JH2GFzbsTnrsy86x
Tedvl5ZU9g3KacvuMMXlDouYJ1zqMbtapxCPV3twDitiVaZ44oWyh2A8ic9vwCuTPLRGy76uQCjJ
uAnvIo/zP4EGDbDeYpsfK6xfdb88XSj5A/yHmkD8BYkkprQyXTL9P2toB68Jk/q6tBv5vgK0czZy
Ab+SBpuOQkXdxWrjQnunomzuQh2Fvthjyg8IW0tjnqYQJ87Puze8To7Zg6Z+l5iVZHni0XNPbB1O
FthLkGYsATw3MMJ62b61ObZqceSmtgxkkc+OZBWmo8CgsAWg64G6W0YqwajyIpoV2dcKYlLrClGM
QkQDpNVxAcIoDvF+WHCpkpn4L8qM3SUQ4iO06JxZZ9OaOpSU/+pqZoUFfyC6yWoeODimoghUlZpq
E4ZLY9+Brl9Y7gqPwNRRUIfiS+VYSI3ZOyBDk8KFkiafLi61el5o8TifhdZ6gLPDp/nog4gpY9ze
zA4OEUCKVaexcP8mOF6cO0HxNU/tHjug3QRY7ULNURKjKOQhUK6WDC3No0k7HwBH2pMW5f3udwf2
Afr9csr0XLa0D24eZfjc1Orc0krSBizeQghoIXhrIT6D3Fzqyvm82s+o5qimHpuCJWtNX4NKYCgf
IysCo9BkSF3TLvZWNY2bHS/UvsToUrdc8V2ufC529990kCYk41HjwKTYm7CriXQ357UKeifYwFCE
JAzw+KFsXNWEgL6KiKM/HpNHOm++ZVjUbhz6FwuYkFartX3iDEqi0dLY2sP9AFmaJE+UfahgQ6kc
HHuce2g1L9VIvjlazq/QWVcWEVTVPe8UB2e0ZBKobKgMxeUXK/xJVqObsbWt1+ee9KOCXo1I8xZW
ej0bzkScDQtK0qtcWYluyZU1SCKYufjlsUlGYL4P8DNGpHbTULmkg7QylRHnigXZrOsotOGag/dt
Wuo5abXsZZghxd5he98TmTbO9e+nZnEG7vBxxUaNrYj1vaqvIYjqI/WpeJ5MNne6IadtrvU4jLtb
I6pWVrTZgJG+sHH12YT4I7orOWUdNTHRoIDaSQ3ImiGHlCl7g+I9Ji5ODlSKChYMCHDBWTyE8Q/A
kkX77uUaRj7UhjtWkiqlolFtiZTkUHHBPQaBf1yHtTAvobqUmGFpKj+5x8mdTJ6BoDAA12kvYvg8
3kScGU6Z6KiibUjlcVVuN+K7t/qjgNwD3Ud6RTZEH9guXuf/m0rwTLHNC0UaUZwxwjOZItRcxrOo
PZWoyl/kGl2KWWezVNqxrewOITUhCP8baRyg1l7/kGE9bJj977pRxdMldhXo+/LW0cwyNp62d7BX
tjI0B8uzW+ORVkT8ixtR0I3qG3wrxycMxd9+XweN3GPmK3T17ah4Icvhs/giSqGrOnldFcxJc2Ia
/3MVB9UXgszkazvuYi9h3OUFbyK2QkIYOtJY97Tk3imjh6JSECeGIq9qv747oD4utKr2Fgh460qg
KzMdpj8RccQCZM/l/Df2rfq/5Z0be7zaopRPoSVX27OPs3CgdzTM7TnzvmLbh7BIbd3oufbmvNK7
VmWWlCXYyji/MTyg+ZsPTv9XQpE8o+IIfF61v5JcGrAWBoMcbatmzLjcSMCXdalt+ePEdGRyAplU
J06Xs9ff6JpW+l+bn/xzM1WkQD0EQ4LYP623aas1ECP3I9YmsaxgReq3l8KB8CsnfeXf7kclb/8x
UTBWMe4W7cSnQ+aOW3GzPDrcKZrHJAr4qmHbmSWqwqeVMUdbWrnmGOxlOKCV3QPCU1aSnjMqm94b
HCnHhocH7LfTcER7KtKwBnBKvXMCZfz3J3k1Np1B2pgbU4Md1jaSNdFeRHZjcfZT5jYLIwmwS+cE
cvfuOzfQqE+tAC517ZyK82EYjkBOB9JvZkQBTyRZmVlgu4JV2ehpCDOICVrrtXKFxx8XkYyh7a0h
LIslZcI3sfUcjKZAdRk89YYB5rjnqxLQ+qaiiIJzv5KocJmQB+jN+a5LqbqBAg7O8pUjkB3iI8qf
wht766SEWidbLSWkOjuLYaB00mlUmEI1NzI2X5gblD0RXeeRi+AlvB1De2CBvy5iQU+MKUInMqk6
N38vUWQHMONRNC77d/67kLg9KnL1vSZOqZJXBNEOv80NmT0decevfgkubecNg63w8AeYOmI6DsVo
xp1gCOeShYZ2/WmcfK5Uv2QDHkAg/8FCwuB77vJ7iDu36YfPiwH7AI3W/Rfof0qv7HLYenivH8n7
fWNYToFkwaavO6Lm/NgopThNhjULmwYYkpyfN+NuZ7LNDU7uB0z4TJn+tO3Fnh2nsJZQ3xTIi8y+
oJwsvQurXiijOSm7UcBjCBb7XAibZV+gUoY0XGjaQip55P/rNrHwVzI3DY3jaQFJ6t45GvXh1C0f
mkbWdsnp4Or0S6jrRCMETtP+MkwY4+tKXf4X3bb5SjysRhiGwbKAYriYLNxPKVmtaXaK8HesORi9
++GHHkNDuvjtpQ3PgccfTjJVempk6fdetV4t9lygCP56hK4tMk+1L3f/C2cNE3SUGh0LgZc7ila7
hCX0wod6/bvVTJGTLoHwJGCdVXiN+CJwLJu8QfpqQsfXawRrr++56FF3AqnFQMxyODefWNwn8adT
b8byClnBxmOjlHQDSF2Ia+31OASHFmlEcJRZ8GFSI7NMAz4xQR9CKhRztGqpUFve4WzYOtmcGIxL
z8dhQL+6PgbLlDvkgb/wSyXBlZGIRyDz7Y8eM03ddnQo93nBQsE7lLTWF8TboEU3k7girReS3o9J
sM7WqbABYaddqq1HHgwbS5Sv74GWJRnchehzZ9tIxfTzBM0erjIGAYj+XEAIu9v9W/pGfN22vp1v
dq3X7Ol4IixVor5ODpyqRgAuQTU1Uwuv3raV8c2n+f+5xrOWVrLr71ni3oRDrH4E6ieSDzETj3To
qUkcMqJ16uPRDaT0K+m2oeeue+FNSydlqRVgVdlh55h+2RxoN37PAWB+ZxLVIGVCEg3sZvBZbYEg
HpTtac4r/897x4SYvws257oT9pfH0O6rcwqLRSl2vncmI/Op/Djc8LxIcr5EUN9TfULO8ih2u3KO
vgaILxLIhHIp4K66vIAhzx/mXn1m2vJcJVTwsHZXHYOQ411AJuo7erdI4lRCdlvP9/96dDJ0xBbc
tX5qpQrTej2q4rMWh0i+n9OFWoDHFm+AIU8A+SzXyUd+2Q77rnB4T5BPN1Ds7k60I3Agwbud6c8p
mgZtUzrKpui+FGW1BE+tPH3Eu43Izo5P/DgmuhTt+4MdOx2xnBmCQwj8DqzzjAauQgFvSMpVI4if
/HFoxgHVNGdNKfXiMkSNhLqSwOyBF0wOb4JQmRgWp5HPFzFky5DabYiJ5PC79rdrEIiqMFUri+DZ
NZ88O3awgOsHj7Wm/3PF4+DiGenMCRiEcY9fm/mxuz+FS6hf3xVosOABfJuQgS9/NOJUsyY5FgCV
c36y/0oB6BGAOYyb5tjFlHbIISOHyLVdNHjWEfY9g3ETfZCGvAhH0BfCS/gwtEepd4Cq8f4YEcFW
XZcUipULsefH5LJuvmxwhSh7r1ezpS1xpnWo2fUWF90vyiLWXKSRom2CkQJr+CVcg4aCyr70YZRF
hhLIzUzUUY8EBeOSNCod3gCP6ORboACSNuX0+aC/8uT1/oD8kXpPwWOBNNdy17iM8kyB/Ooz4FR8
kY8AJxUP9+ipev56epe+Q46RZYi9fZPUonOcZUijIs7MNSBoHNku8ir952W+BFx77h9QQzolyTnG
Cp/tDEvS1InCAeSROBzD3wyRHUq38/y3byodbpvwBkE0W5CMSCXRFrYKJLEraBMbaHHqE3bxKxKA
6YE2gqW9nvGQyLj+SIo0qBLkXVQ2rX1yo0P1Q7uYCakGZM7bch5lm4+R5wBqNBvWXGuEeP2Eitac
kgF90Nv3Cfm0+kdTFBjN2UDdxvC3pACjJjRziO/hE9ImkwVzOC585Ljo8+8hQILzyokmHVDnBtWZ
QHPpImPX7qbUUK0opyl6fauCQodAW7by6wtuLW7tKItWqRdbz00LSzZjBUYmdFR/LS762VNoGqut
eDCQoAmFBkRU/aUIO6rmcQRiFdmtDx5gZCcar6ywIw6CMbnjvbLYpuWFLZW2kdMbXPdluzs77xU0
2Hi+6aeW/FlRxSGgwH3AGXQFW6+yaVriGyTaxOyxooyT6nropMgWB1wq7nZAx0IwpmGVG4D9ZtyH
AobK97j7w3cN9KE1RFklKITeiyW2G2B2G03j4HFHFgLDFLefVA34ru/brWTcDcOk9FwS367LdppA
7bas5S7L1kQSCsTFs4lvdVrL2Ojr9wAFHxOoq7bwqxREoBAGoibDAmuyTL/qEa20zYIh0zkcIpFz
sN/m5U888mS9aMqLlFhE+e/NYxyFbw+K5TqdcZVcYACf85EPIVfBSeVdsjuKDgx1mg7tPTdeCyi+
3kq60xRmrU69LEl5uSlwgHxtaw427eJ/g6a5sqc4F6Y9xxG1XDGhWqfQ+lTAuAOq6H8PWmXnWeXD
v4epHjX6vvKiRIPf+VVp4FQ4OStR2lgadSmDJMQJ0RNId0adzjUn9Q4muMfS6uP21r7ft+JlE6ek
fimdrlVMGzVDoSwOsfO1bNtK62LqI0A5+msBRb57kQCd2aSg+Z3JUaPRj6fyvXcYmzIR6ba9lv1M
slaOnyCoe7NYSf4rjW6kKdDhi+3LnhONqECYVYYKVnZ7waLl5uYwMVMz1QwMhFBROCB62QXiAGTh
ViuRxK+flUlsDRl+hMbSTWIj6IrBy5dGxk22sZoHZ+Y/4ffGR6d1SxuFl2h4A+W67pQc1/by/Oag
O22mIFRBozQ1e/0fuMX9gHx2kbdnNN1/zkRUbBfJ/t6g7TCnwzsRVihldxmW5MRsQpNex0QcTDD+
AY8bbiHbif2HLcjQONnOvqFA7EnVh6u6kkq9VY+97vu7/fzqzOPrzAllOPpksDvXWmOAbigSPFX3
aJwMncEgbOuB2rJjuduWLKbZGrwTfUdoy980FAVkxsZ5vd3rOi+pXnPxN0wsAFNYVph/s4QNfJSD
7FMMuade5+TBMtVRcLAtkQAQOp+P8MHrMedua45rcbrdq9WrJ3lLoJBX4oCFQNG92yDmO/iRqA1L
XFu4xS8W0zhLavo8hs+9h4CGG8YFbU0BQ7PKOFSiu3A4FO+puUuVkHsPIwHekhtDFKq/cSBYiHv2
9udN+TBOWGJiR4XVjYyC0AOkZUEDpZWL2dqH2FQwC4zKFHzj+3xAsWZXBP9dzJOafc/X0/wwH6Gx
fMzOX5s+IdLghWebs4AGnaDE58Txg/PY5Jpbq3/MmFIfaF6Mh9DNAEnYwYag2JNXGXcrhkKH+vEP
uVU3uCixqekA064suP0ZzzpWOl/DjyIiYFlOIJM9Ncn4NDkImErhPPLPL4KBIVF8Gdz19nIQ0HfF
xAjz+gUIj+zXGfIrquVVCxrrLbe8jnwFNemqmPfQBxtMvHjDdxHWP86E3PlIN+FgF4JCcBFrwsaX
RA0tmRRKFnoBIDePWJLOathJ/RwAxa9/74XK0qGPGJOM88XpfWypnTMojFohErICQDGj5EMxx6Gv
09d7G6jPz1HdSVcIlPnY53JoJwtOBl4LV0IeRF8FmUFCLAoly/A9g6OBh3Mud6SVMB00gca6BA/u
ldM7heC9hkQYthkrZgDPtZBSpC0Y8ZCjwQ1QjwJ+FSCDTXDK0EpN2uX9YwWLVunGMTgu3SBnE0cP
SdzW//Fo0UkCJlNj72ncfITgN1jl7BLUKXP2ydHdXwr1kAyPjE64X0usdhoj4uv1obE3tND+fxeQ
tcyZpeMRY5JyfXFWxpsi6SCaB6ph0Mh5fJGi1qhYX5iepdbRbzNZ1I8Jj+IWczBYtwUo/WB4xecT
v8LgB//aYZmIsG33/n4dNUV2t256rgSAgWIRuw9JfR82p8XPNkwP/6lTgniLqPQ6U+fnhAML53mk
SLOR3+gVsQtcHhIHroRnABq/tRPEI2pclXhGddfRy9OVDDMkaW84PmE5lGxANhprXuXBNXhw+OXA
XG8+A/BEVb14FUe271qBoAWoDIErfeT1FtYTevQzxSXpxaapnj6ZzX8NKakLUecqufAa7hkt91eA
6sjR+dN+ZGroKxOxXypoxijFMpHuA5AGFKSh0QkjdVZy5duCcGKUT3myOMDLbGwxwHFEANN8Pbbz
xJcvO75lY1oUO50qidIlbXkpMRINVrQ4FxWiNjtgd/MwyMYMQHd9ZZy/4swrpuI2ZHa+7Vxpm2j+
bnVSo7fnfE/c2WVahvWbixEf7ZmE13qSu6cMQhi5AZ2osVCBZtV45h74T5i0YaIZCuu8wo+AK5E0
9sv0IOlgU/F56JyrRxTrIykbCUpq4csqg4iy9i8hm33dgeA/TN9ZZ8Jr0+T234XaQsin3rAAJjxE
4h3ZVNcmRVqQAYcc10AEa9JqAMDbRZEQUmuhFVuwyQBl9VtfOIBQ9o62ZpW1+MMLxff6O1vHfE6Z
0NZQSuVECmch5eePwpVuOYCsmGd+wMpUKXI2CuRm8sWPjj98u1UDAn73fnqJd+M7pCeYwMhKoM/Y
//UxJmu3jSmoqk4HvXrJH4sr/VBmQSbS83HCzF2qvUrVWf6J30hYJETvlXmMtioyC7iSRSitv5hb
zJ7algQP/UphEqEyB2ApJic/BM+e8SxOHZX7bY6XEuJdNFeAQ+3qXlMCyPxGIhuOXeBsLxl998FA
f039F4uIkcLM4Lu1GMHp5iZhwYt1MrqussckUm5D36lKGeHgf05rQBknYToEh4G+bk5h++tOUEvd
JTcsYLQKdWQaTVFQ7QrZYZrXjFKOy7awAr0RcnFH6fB2rrOZFCGGZWwCPPO9OlC0vPgRigsd5ZX5
nNuV69QiurJ2Bze55FbMO+of83zROpe7eX07gLm2YnWUGPdhHPeXGT/VR+usOaXZ57G+hdvms1/r
+gbtndfBFJUxUGmH0TqSUzft31NVs6h+9fUu8QS3hca3QIhHfaZsXuSqF2QhdvQnI3NkuAwsB65T
JkaTnHcllZstEJ+1p8WxpHHB7gDpEPRv0IBhHM5SdTTji3nOAPFeTbk2vzkIbu6/bffI5Gvlx+nm
4hehMFf5HaNpjLkEoGpHWwPPoPg7PJ29tr0n9eKFbN0zQv7MV+HjgJr16E/OrfAbYTs0ixVMZ2UK
hRO5817TmP6OU1o99kBdBh3gZouyOqOtgehGTZi8NLbeTm0iShxRoPK2BO6mzj0iy3nDMZhutuf/
iWKnpk9AfY65aONawUKuancwwDjMeyxG9n92STbNAK47HlAI0mEvwNeexVoUVru+vyLlJLXLV0dl
5W4m8EM/EXbo8WdORK63CT2pyf9ydEn7+kFkwhRXn469f67uI1HZ7kMP4/wDYp3lgcLDwap7fm1J
0ZbDnvBEUP06jMfYpsqpXuB+mQowupZBC/LJu4DvN0RGordOreyNXF6Hd0f1fCBf4rcmSrVBQg3r
GFFv31PPQeojf9Ke615zfqDgmbEIspGBemSCx5OBJjPM1I2Qpf2Me4wOXzbxVoEBpcDMMq2xCGw0
62iVSpuxzDcI2zbAmIChTNKYn3PlD0Ud361V7BA+0W/d+TUcEwju940cmJQsdbV6lmQ++iad2AFJ
nFa9hQ0NZJtTnd5nK4vyNDZSGPhqIcmmebxgAg5DdFLY/INRCVyje1szdYwmDEgnol9jJ351CCp9
9gNtUTLdmBqS/S7QWkovIWt51E9anpGH6XzACsCEia9x9tikHfOAGZBFit0lkpKvg1/sa4MDLBg5
TXr+kE2dTF4pauKOlLU5h8gdCxtUdhFRhQKiLJgMYclqsjweIuYh2VnGcqlfyj2ipRXSrO6rp5X3
gQIbHKhqNqn6GBkqiey4pcGYyOfjxMXhn12lWSAMiglj5aR0CZVxEsswrU/9xWzde/aYjoaXGkh3
edqjFZ5k4zml34ceLzvclQwgPlbJMzeQ3vWFGSyuOxsUDYY3M00/TNQvay2fBja5k+P6XMgGwjtu
6zVQWtT8ZudUbqguC1tA5TrHFuhUH+wt2wRhgLtSmH7VMqbKcCDP0ubdx1bafpeHzmjfzPgxT6tA
tMsH2pPMhIIV9m/SDQIwqSSzb8INflo0RIV8e3CtjZhp6EGnw/5GqVdKvqURCxZefiH3CbrJcsJF
xM0E5wDXIddd6gX5qmvSYUpyROG025hy4704NVE9KZjad2gWV/dG8mkLEcvTLF1wxHtqICmXR4MA
MbBkyqIkoWAkL67I4v3ZSuFEpKHzS/LmsuoJpvq5iKIFLs/2vQdCrOg5YcPym85N1/RJKCnrTTXe
+UAhWHWmXGtxBDaxZASVi1YM9uRXuOPD3hk7bf9O/IxImUWrBZkkhL2hcYXhu6p2SRC7j+uSZI/P
T8HSFmjzfFJwcN4M945BJYSs3uYa8wB+ToYF5k0IJBEz56tmJNV/vnOVgRtQzZ9UpTaLjh0vFtDw
I2j5rm6C9iIv8br4uPoMzSTNuCfGzVeciMn4rlIPNSiPCKinXCFOJQWeyPCUEsWaf4k8JEl16etF
dh6Moq1+dn05izaZn8ilCSrqksitTgspzwfGpbkDgHdB7wUmzm7iTgqB4SVInt65P/AFE3xCKocB
0trcEPGo7hBtknRp3NIapqlNrY8Xsroy+UgH4NAVr7gfKIwynukACDeKXxyIZOlAMeNKMgVMoQcN
2wuJh9NGC40NoPXfWrzyng8hDycgrk5qxoa+ZWJRzPfXp/rbEWjvlKMOTWsnwfuV/kWW3E4dAmaT
Gxv3606aRYX9MI/9uQHLvuqcgcjrdmxeojQcYBGHbXhvDQfdafICkY4ljB+HFKGP7AWufTy3psLP
55OxVW+oHsFKA0hhAcSx49CHDK5+xZL7xFpu1FfbX/4QYueqEYhjHKsLzHM3qNjQTPParXHiMJhv
RiJp3MBLNSRyaZiUUQglh1lX39Ab2nTzYuuJRKiyqxQLrLbQzLTid4my3VIKNxLhDD10x8ybE48e
D9htN4DWO2d12gYbygmXGOpXEN/s9bnOKnEpbO3HTeg/5d0eChuievryHdcTrF65+P0VQMi8FUEB
5zVKtUJVy1TXdb+NjAmxleYwa7+lbOCZ4oe6EZcpwTmhhihXf9YZAgt0T/VjcLg+yAKUYZ9VmWT6
5uyH4AzS9nKJGzBLqsQvv5uIURIG+AN1iMZ7My9iV+NKjCs6KSE1CTKY9z8LALvaTp1/tYdykcK5
FVXMEpgTifNOMCLOWMenYtoHIgh/mHJdBNHga9J4oLyqcCDY9P7RJ9Zeebm7yUQ3fd/W18UUDvI3
oQqyS73eMA3Ehi2pR4hsC7b6v60H0PGKoYMVK57ksgUzDEroRmWxKdWbE4/vKR+qrxQLCQbH6oev
P4CPSWo1RE/nyRL7k9y5ed4oZySqodk5igLB+kmeRDsfCF1GPDgBhinfKKOx+rxC6hR0p6zSD7Jx
J8BMrDbKbX6LYhHrTU9ya5UfdE55ioc4tD+8mAi/NBDwEA7ZJPlnVCwoH3c9JEwlP1iaimR5JUsB
zVMAz2b3pufyotN3ffpFEH8mWwoSFau8JgYl22PMMMP//+V9tCg6u3zQPYyA9h7UVZrONXUiuRnS
AGYw/WqpdKVcKSVa+fx/lLoZJNAyUMN5SivBEJ3q3sDQWdjYd7Sy0hT6GZZsbU5Ow+93+ZhrCZdf
Q2TIg8Rptr5Du/8gtAGJf1f/0Q4GZ03s/DScY753WfdpPv1ZWQHDZiiuxL9kzy8G/uzg4fuvpOW0
e5WDPj3qGEe7msaacMCMtcbmzbduUQ/JzEHE3N672Z0HAILK7jpFUw+tpI9S6DD7EzHEz0UF5FiW
dVbPEJz7dfqN1UpfK4PvlQiiGTYsfnu/3RhPiWl+FSR5nJgTvZ77yJURmF3t0VYkFRbRsG272ssw
Pu5VqQDVKQWiqyaZx13zfs+p3202eqnYQhsZJrFepfPPKJN3pUG6i4c462KmhDyXPfoqiOnAIRBO
Sg2NMKlp/D7oYe1bQAj8BoPAbB4qXBdFjnTHgepB0HnHwVgAd+54FMpoWnpe54rTgl16h0LrKTvB
Lu1VJO5LwUBvp4sZsRxTav81OirMU9dfLuP01Z8abZ2xfBb2SMwWGYbRZmpgGPFlCIT4V3Ji2xoV
9TYdCdvnSpwcTyJKXYj80yb2Sj5OJKtB1ArKh5qt+OROQNLjbjO6aRSfYOtfXs1XzXNmOStXICVn
z5VoR5S9fSuUeZ8Vr2OD4qBIfDSWS1u9rUPM/7M/X0CvC6tEBxutybSZR1twLjzPWDzzsl+oUYJP
EOmiXneIqqpA1k0lziMVOMj4jil2yw3Vb7ZSJULmt4Mgnbq9UmfMQDkfLzNDjwb4yd0JNfdS7V+T
DB3h6kXatQ6X2qJ8pckqFs5x6WYI7L6BUsEsw2Fx7FhDyGmXYtrL3ek/rD7AKE/DwwkgY3myXF2T
/dcntNyHf4e+3UJ0xbpJCKXxW02uv3ndfGAnu10mtxjbSzIJKmGcXNDWsc9TKarrD+T52GJBP0HH
UoDOKM8T34UsJ9BGInCFeC1dS2EzvYu8jOVo695NxgslLLJrw/GyxSS1xyBzGyHv74NK3kWSJL7N
5QRoAsJ/vJSRK56+l8ew24PculwAll5gxccEeRe1Hib0nUR9w2lIypFt797eid3Ru+X78hZxz3Uu
WJiQNOdSVW5C3lnfz5CBe00wi4MCbKiZUTL7uAbWeWBXIb7BQnVaUNY9in6migjrSI1fhw0DyHU9
fEZQd+StwaDbVz4KQdaVbqv6quFVWYq8sp84TpYmPAAvfp4pZOq+M39UbZAkDLirPW0hqx0bw38K
b0mPmVIN2Wy/Zf+YWzW46XcOthfLl8okSCxSmfR50qpm4RapsZCC7i0Dib5HBwGwXcGQk8qkJumV
rQUFKJrlBYgxHH434GTUep2O8n4eZgKGTiaMKfLAWo4FdNHCaHLalb7B3FBz+bxyOKb/C5ePtHB2
vW8r2zOmbxu1Z6Bhrl6wf1wOI7GbQzr21m8TBg0aR8wIa0ynSQ6uiHPTQTloPuOdzXCVeEbNV8uM
sUsBTfpneJ6Bn21VK5H/zmdkVnamkHly4v8EZHBaVIKQYo1aNVxGNB+Rd24SsfE11e7lN25mpR1d
rJ6o9oMMbNDVumN5WtpK5Z4ZPPyOGVGGCkUONk9BVEqpuzZqPJ0yNcI1wW+JKeQotcchznnlXQpX
oOC6zkZtuJR/j8ZyqifYIbM7Y8WZRFBg59y+nsr56VGthMqL7KRtOgAOMwxjS2pz+2L0X9ndfs+I
a1gevc7+rRh4cNkfDu2qMDFr4Z2WAh4QCA1f6yldy5EYMBHXIO/1//oDsls492ZgHkf8rWunqDgY
uItE3J67Wb13B/dgtjeDRgfFgwOPz60y61+C2ALJTuR+tkTPpGmkOeyB2bRCUltFpeyV0/7wQz1x
h4nC7Q1zhrQVWIeLJOJ3eWfP12lq4x5WzHs9JpdukLCYeLMVV/LtI6SRD37U3MKLgijrL3G1HG1R
/aX3m1osHfePYLJ7gAzXGcLp84PALQ4rswSYOluNaq8fY5ZguYnBUAFjWm4ITLaefoivcFgFZjtz
1hK9yb+3ziMTY64exwI4dhaQYCKHaqMOJ/i3V78kmIlSzgCzaJ2t1DTYMmUVZ+LcyIkxO0F/sHxO
8ADwAUepgv/7qhv0jvxgkyYnkME6LkbuZw4c/mAX++lcWzZOII96JQBNqdjTeK8PUiLxn2HBTDlg
IbZa4P/P4f2vTRBaljiR48+PDWkTjIV/LHsJ77OMooKG240pQAEY4dy99Zivbsd4nBYcmvrG8Ddq
bPuDgYl4JC6H+RiARHeq0pAM2U4t4WYb+9EXZEW8M8kN/NJ3Av7P2oyCR8IJ/VPBVuNbwXBl1fyp
xeKqj9zUVL0SiH0KmRnoM05O6RFJro3YTrLJizFe/hcccVWAmyTnVynXGb/ikQ6ryloN31KfNhDl
ZXYVG5GvlcHdxKoPGTIBQfCcPg3rffYa/foUCoBhbmHxP5xsmTTc+jvDIpVno7mskjNmHEkAwcUH
BxprZTF3hus/rUOT3z0bHxT93cs6+0tMjFQM36lj84QH+V5qbV2k3w7K5OG8RYdSBmrkpGflpuWr
yYoFVcR7UHRBa1sdfRH3xZGCYXmWvGm6Cx6wN4mUDwgzkBjY2oIf17BE4j5ZrXNVdZj7GRvcT1zx
b1XVU258FeV+fJ880b13Ndp8tarkfmrZTfYZjGsnnArKwcTN3WblUXzhqKRqNt2fZUFc0ulRP9JO
Xe4BgWB4/7SHe4Za4l7qwCi78NYTKmnRrL1UR+mw2HvJdkqQOJ8sq10tAr7D4SGgX0YJtA2pIosH
UD0XYDZCRLe+aqdgNgq+zthKJ3216AwfwahMrJNCLs3NagLVkTo5a1ihc0DSuoN/xs06Ervc9PjM
Ydc2yMUBN26QqBJdCxYcWwCpifQT+fwgqFz8v3Xa4piC9ahhvrvi8HBghtH2ctE2Xc7bHrJsBEy8
EfFRKfZ6JZWNgasZmZ6U6bHNaJF06nV6sUwgzqmrC+eYWpQzwie5oAvJ+ifdcpsQVlK/q5eE2Ut3
67vuv4BYiv9bw0yk/9SfZOqc3rn5a/YpbhpJAQeXawxT40ty5lbruezIL6o05sDGPX4QrX8CjHR2
1cxJVHy2cAmwtvnKTMiGaQfPS4Ho9wDLajL0e3pJBcd7thRl8GYTGSukYKnNnlnmlYDWgOLdF7D+
uDJhCQ2OGGBkKE6K3zfAGmXKFwfc89JJS7XYhTurZmEoWw96zj95ddB/RSjvcPXPjLHiD1SH2Cp7
UturmfulyyyUc8oR+lV2x9VzplXs9Ex4zL/Vyt2ZKIYOLzw0Gne5AFZFkn2NCjPjhNwjgyqIuzqv
4jpAUim0vQ3Sasp22RtRpmwIMcMd9T4So+f7v8yaJ69t0yzjL8Y0vXAC7mZfkyDRJggSQ5E6bxTa
O+Rie1dYHGwpIabioYocoUTnblNoV/17HyF+LmVc6aMkoIBvci49w45PRNJ97nSTminQJT+eYeOe
8cB2xzG5f9TySsc9e6/8NRxbiKNpiATLE2NE6hmXPBYLfH7dJac2pYWvxmjBKMtdArzuOl4SxITT
COzSP0/yEMOJTlfE4lYjkU0G88rS3HeUx9pa+0Tm3YdpH4WPkNV5KKz1o0SAZScmjquXzyR7zY3e
G+nViQG9RKCa2KsEsrR+zjUrkr3UMvOwqmkvDpy98zxFfCGhwTjoMGL0JdK2t17hEXY81rzXB3sB
hPh2+i66ZA1gnUlfWC9njJBcmnkRAdLtOm1OVPYAvzG9nZ8Vb1Sx+IvMC1bY2M1LazQNZhfhacg+
FcnvGvFgnzq30aAil5yKkWYHVWJuPAegBDx2xB4TxaotAbnA/BJTy4yuhf5EG43kbIHTr1saLvR6
SMe0D8WdGyBzbPHNgf5YaFnWG29tZO++h/pZhjoKkNDJxSVocofrTcapYSht2CnD+mDN8ZaSQUOh
NdU1QgeRe0H2TtfYBo5gxcHWld0vpiL/VUQHDo2VoF0txBt57X2QHaWDD/kiR6tzxLGJIbdOH8IN
M5haAlryM3qVQaf0Q4gQNbVh1K3UlKEwV5UccYDprx3bH27ezgBahE+46GaxeapWresHd7uYAdlw
5OgAPeLh+PR4OK5XlfC195sGiUsCLgGjPV2/LdvQnQUBGjCN/Si9I6wfXC0L0+85YczHQf7J6q8j
g3EfVmaU7uceOGdENSuoRWleSuxJnxITT4MegskcV99l0dq+/e6piBoBFLKNdGyfuxPnmRqn+3/R
kclhREbf8LTJDp77UBAxxxojfui/Lq2pu95iViI1xg2RaPphmkbp2W9jkMB2i9xYtsLzDHVg5HIk
l2ixev66N+3Wr96V7mdLC1VMV/LRu/yTM9PQZ6sx1C1gRK0czeYeHXgMENo8DGOE9i8IrbCasEEm
D+J8dVuqr1W+OoTEalR2u4KCySj4llG1Mu9AArJw69o9j6HP28hTNi+1xOjo2bQuuqvQEduLkVUv
Ik6j2HqxbPuriBq49oSExuc7q1lVXbQ8NKpfDQxt6OQEQuzuQp1dqcFM5ciyc4+fzk25D/VNt8Re
wpn21eoMTvg1Jusxyko7DSlqpDFEBMqSycSwk2N3aW1xw4u8nnmaRRZit+CHa0M7XfuHfhhjLgHa
I9dn2HVaDntw3k31N+CMSWmqk7+D8oBN1DpzV8me8YK7RynH3PNX1+M2HWzRi/22bLdE+eOv71RC
X0VF6A+jEX9TWyemGH58PDz/S6kji6GtoVvVugEDC7C8gZpbldjYkmdxAwcOwN/WyQ8OugkIHxOT
CbwOhPHsJTGBKUcryg254NDMFjIsCI8AO+tV0h/wNhrmwt0DkJBIryEpP9CgEX9EdTc0Mv325M75
yFRzRsoqJ+nDKfA2MTFdYwwO9tebSnbXMTMWlhd0JA8SS079dcAPJQhfZrRI1tAgJlPux4NAEQOP
c8PpUEQZWS/gbVYn0HrSu9YLhySBLSAhgQ6B9V3QYilvHuayL9fOa6u5jDuNWTNW8mSRiv0fL72P
Lp59GuI2s1I6H89PSJs+LTDoXFi36GUsBrHCMca9P7E+VNoYcF5S3PF7c2Bvr3hArrN6Xp0nwJ6X
Q8LXoUJMrT4hAEdWVBFDLE+S8f2AjcG1bAPDqzDWjBfthqYO3T+Edyg/V+f3HE4ldTunPL54CrFs
466t6J5QiNt7OvVPerwe96ZKyzQcaA8JG81AF3N4EesttlcgG4Z65DvdjWsTnyZyB9BgoWyHytr6
09Ujq3kaGIV7Clzvz5qAILD0FPltwPCXpnaS3X47tJtFN7JtaqU7jZXRSCTHBPrgc+7iOWuZf5Ly
Fu+pJQkH63Nwh/VxfZu9yOEucg6DnjxcdV3vwhrdJLrzEHx3s5ZmpydFF3YfSeOur7METUkGQEAi
eWRCvcSwdkpmyW2zHpA+VqugiLd50Hv8FMoJqeVBMpZcCkLzZIs9hgb6EihD/HOIUvDC8bJrO4kq
xZ+hW/5CXo5SsGa/b3gnkLzNoo8OzOyluq3ECbvCXBlgD7MoiIn4MFy3gv1TjA65vbGxWo2BnDv4
A5kxe+Z7M1vEOmKhYdVMzwkHnHkx/L8hcoi7rwqkXYrG7uvCjn4A0Cv4m0G1kNgnHm1FrOBa++So
4lO512vjeuVc0S2HrVxptUb1p9Lqt/tVBkh9rSfMPwo9c1eDuey+HCy7mqSEQYRLY6Tzqca066Zy
Y4fuQKExgnJOsu5o8biCkI9/Qtk07YNcMBVGP+qVtgmR3h4iuwOeWhjAcPCP27pzT0E+CbXP9UtG
1KnrsdthhvGLx4vcFGWhVzS4ks1hjqkG/l3Q3+Xw+oO+rvgsE9/O7NTDJ2kA3G2R3zqKdcEIXCTk
GMEESupPZNLY+7mCFPi6ORkkAhcTHAwMuiVZ1BssE3GxrGLGg4b1c8eYeiLHPAeYzl7EOGrHxvb7
cB6qLooSyVzN9e7fb/Y+G4+6KAE8sHaD2zv+qZjnllMg4t6HL4gQo0KXOm9/RaKokBkAEPWzxKVT
K7w36LMiC9Zkj9xoTVCGyTlMG7vaM6eMKs52DntkwyiUIhIX4JM2bwxDGfuIN1bC2RgeTllk9/j7
NHmiKr/kVRfQ0Vs4oR3MRUx6/rqI3bWq270N6mwgPhoX611sP+CSt70z85vfoyMrAjFTBJLweFa2
J3mFo46/pE69/KhMU1rhXVKIIXXhBrdoSbiBd4ACn+IAbg4UIOyNuNcKcv3Np1HA9fGlnHEq0rZi
xqvzMtR5BXrebNomujpFnRQmo1BM2VEchFhUYA1LWi8fNTarzIr/WtFCI/IQ3f3T7s2JOE9IDWPM
1jCL8wgBVjDahbLgYk1YAMK6quXiIrctVoFIpR+eGiR76dETukmV9nOvyN+X1XGwR2pgUi6T59GM
9kGiB11OGPXLU+YooOyF2jNwaMCW7lvYUHYl1Bw87OcdMnT/Bv+Ot/Ym6wQAyOKve6YQA0MVbbeh
gqBWQVtofP8MCSkgsWXKFTEPV7nTnG4myUnZlRVY/m14OLpZGQmFrfaB0UNUews3hhH2+PnEfaTG
0/Y3I17YqQxk7WeUhl603cYhoMiMrOb0gabyIt1txp68U2moBlA8vRXnlN302Rf8+wfn4AX/RTZg
qP1wFh8ERDvS6c127n492lMmtq4x/7wBhvNHXyxVQW7jmkPS1RHilQpBiOkoU74VmGRVGNLD+W6m
jugvEyTIvPmfDAVB30NU2Jqz0MgPSZwuOirT7gGOkBk5CzByFKS6J8kTrJFQz4XNLdWggDm1fbR3
Bz59n4iQA0wmu0qPZ/GFIZ6CKd3GDET36YngXCMEfV9WurpkQ1p+apPgpAmWgW3qD9nEvSowJrOi
xgTHhFJWDeKreFquXQC/9GBKjh0fSKN83+3gb1A8g7u6hppKUH+Ec03bQMTBlhytA/fWj9T3pyUy
X2Sb2c+SvNRT5+XmGBbSS//NN5sbc/VTf43ssW71BkfBN7vlPynQyJeakHmtGEavwgLyhIA9kVH5
H6F7qdHennI/919/xe/8ByMfnLlWfV4hgo17FRb17qwwofnfpK6JmZbiDgLYL4OWiMQS304CUNr8
OEDJ9UktRsvBB5MOVxJEusI/vloQ+qMjmrSB+phrpOBYSyOgfUbnqrjSI1OOcGU5fgJw7FXalrRn
ESmM01eUcYlVY25WNpo0J9ZlUICwFPftoHnoHNPnR55jlV0LduUjX672hxSFb1+jia0DTibfzflT
MabhQ58Ksc/4YRhSyj7T8g70v41sJuKlE/nei70GwT/UELKKwACP/BOuITveuFF38T63nACduQEc
JxRMLpQLAoSK7iaAjji8U3MFvVp2wCmrAzPdi4gwCtE6zvbigjACcYy+VpmZ3XBiLPcniqng1reU
ZxOQQSlKdQO4ciC91Gf9ouLTVq9vPaOKauDsUYv5Bg+Em7ERG+a+Ws1IlDZUOQJE6QUqSFgkY8oK
ntNOGPcsRiQaAmJ2pNqA+r+kdOSVt+ZwwfM4U1Z6qMSi6VaLVnRl9F9Y6Q0z/aJzT9YsIInO9Vml
0eUqkR7fXZ7hdnVNBkPK/kuhaOANcnRZNB+UfcpPhLp944rzoUPXpUDw4NiwkieqoC8cDoqZ26Vq
zzkSx1NWvO00JzH9HqFbbw2bD9UF1WMZt75IR7Yye2cBJMYojDO8uUPzoZJYjiNnSMHCJfbsm8TY
ae0e4U6psT3EqIaiB62gSGH2792+MU5x2r1r/UfExdPxalLz8TwRRrlPDZUyDjPVfhFAnsvGdlJe
DfEyl+1KBKauDqFsDq/PcSgQUxbnNTa3U3J14g8HbHYiR0Dzp95niQ7a6pt7xrBKwyn/F7F92b+q
R4HtsqWeGIN/2DH4Z2r5Ns6l7rnMVH2ZdpKosZiQtdHe9vnjaQdUDlyZzGTiMKtmwyv19sk2UeF4
+aj82FL81GMMAC/d3KneAbrBBT9xnEQMgus/0hv1MfNVBmB2Dr5TR2XsigUA52N0qrvmhb12IMf+
YMOeDQaW9uEr+CUpME8cO+XXUnsl5JE0U1R+VNxF8FpkP+3N7/y56t4M1roHiP11UJXJLsEPeQAM
DnmbBdeGlEkQU1YyzI2ivv/tujtV/0YWfF+TWVzMV1hiI+gY4mH4X3KdVteSEbLKi/dZjzVQ4VZv
C8R+OkGIl8Gg7WC1CKeusj5h64kNpKY9lnHOOh1gx6fj0M8neGDkpeFX283SBNsgBeJvjzwvRDQy
wY2gk2i/372rH0MnSvlKnJ3z4r8knqbZxahovRjQwwN1kZGWgFPaE7otG6Qu+9tHGz5VCsZ2/B7a
XD21BuOSW7d9qFf7is7qz4DY6ew6OdI68UDA/T2gSzyb8bj1eMD/6jlwVqMsNxoF3dO1KIGoMbCu
2vN74xTAtjpC8IwGS8U6EoUeaoarC0/UtfCRazle2JzSEDJCP6oZDLGd16zpOE4eT8UnSS8341XU
6SSKanHQua7jSQTvTUMQ9QVAaBPRdLn33h9Wxy3d1pxLzI33SIMV/5Y/A12Uyn2FhgvN88rmvKSB
lFUus2Re31DcjpqHx5DbEKc5Dfv23nd/w9sSeEV5XrL+TZI18Na6+LqKsxMLxJK+YhdTe+yJa76z
vGPtBs2nRSiAJbbNZf+tWfIFUBUfrDuKERwGukkzHr6+TezQ/k8Y806FPHMqDR/e6/vJheEYoso+
rKfxgGRMND4m/CJ1KftHgaq/WYQZSVE6Ma3sVU+dorm+QKK5rDWDksfjL7xgezsMJ/pGg1/xXiRT
oZ0Phs4Yj06xlaEFPAl6/jGUyhOyO8HPNws/F3pUOVoPYN1LVKhbhWGa4XAuiw6yzIX1blUBJ3wB
h9OzrnV0sw0aM0xb11aahmyJ58ZI7N70WY6lQrFCIo7gtsDQd3n0c1sWHpzfhvV6H8Mz1036z6gS
JGDvEdXOT94vde9OxHq907Iy1u3P3O4Oel+QDSmx6Hb3bK/DU1XQUcl+EPbbI5aL8iHrmUl3clBm
EfJv8c4Y/oD/ZwBfKLV/M0QAn9mOM+0vRYJZuTPtUFopuSPGJTpkIRfCSzNDHlJi7FBB+J2Ygt5S
tFcNLOZ9VDEd9KU77leD0pZAhr6eMNRZwX1pR8N+FG0HLB8dac4A64k9eA8of23S2Y8Uivg1VmBi
WXqdWasQXf3uqWfvPCa9g3eSN6b1EeJk12K2tr5H7LJJ5bpusaOj6EsbO5TqQcVNtzzTz5ZW6rvA
qBTYW2wetlEtM//RO10t8WuXxja7J/h1AFFV2AuuPhiyrXbrxVSUUI0ee/47deIi4jVPFVKjXY+m
ol4ZgypyANB343d5L3a1fR5Mq/QyG2RG22F4k/10q7K6MSlGcYE512Kr9xsqJ7pq6y3awzgNuxvv
mbx3U1kflL9BHCYSXfvD1vVuX7FNiVAgEP+AZUFPtG8au0op9J0+NHqjqopyAi4JT468DqKX28B1
5sg/inc3IeToMjVC6J0U7e+/t8dPbuczrOW9LQytGIFIuxDCysj0DQAIlrWoSVeyODobMU55jp/r
4w90/WreaThKwOX4LSH7ikU9trjz7rvky49YGD/zBeB6Vcq6vW5YT0pfnHnyTjXNZ0HSabOUAjwS
li7F/0xtIRCTlFrFR5jdrmy8KfAAAbaAQZyif9cvU3TwrT1l9Q/dyJiFJjnUwHjgF+lHpDthq6t7
/BwZyLCCXC5GfYjIMsD/gyy0rCR9CUrHkA7RckVGaeDEnTPiUCV7lPafuJGeQxbPfXReztA1y+K5
RDMdGqxGazb29tkqkKRsaqccbXZXZVkf1MrUKyZO7kDLobVyzw1zDJNHpH9o3Qs+XHjlJSwKqm6a
/K/IPtIdbSOK/hoaGn2jU35TYdFYbqYsfvXI/ncHHtjRUahDfdux46AMdwm8jQJleUIGLNAKO2H4
jClNndcVbXOkAlnrOs+T6tVphofmsCGA/82lStNNkZDHCoYtp/vXh8256coJlKAmKO6Yomq7I5ts
7IeA0vQCmNZyhl/0YTToH9kAYWE3luvPWmh8qNLsuB+E1lguHrskc3/jdy3cwwEE9fMfVHQjkSBc
xUcrE9tFPuPuZPGnNdWm+xJAoIYfcRHZ/tACCgtT40f8FvTwkMgYVY4uaeAJZvPxUH2WibilxJlJ
oVdxvbBM/CirZ2bi3VxSdBpefy95jfDu2JZvp3lNFGLCctslXwFDeyJXPLiJz5EadIT/fmhz7qt8
Jn8B9uTp1j9ZRb9jqBNPC9MiKBZ8VFB1wcy25YNwCRWKcn6eoCWnQ2ygwIBiUTyjjd3Frlomh5Ge
zyB8dnaC5BsCUo0qswgP1BLN0sCRCibGV+S3cxnBXjs0liWQ2L+PbTa+oPsWb4SWhscB7a3XB/bI
KE2iQL8wHhnUFpQC+R6EY4FhzKGZ8L+OGxF24oLAaiKXpYWazPsSa4DQS5/vGB4Ud4bia9VSP3hM
DPb2UPbop3U3CnBEzUgZuPWXKixwpMIhbfgNHfSAoaaVjdjtcVcrdnYxGi746M5F7RdpDkCUqkZn
aOvs4PH+DC5zNRI4h3piWz/q2XWO8v6AMgOIeKiqod8u0I0nqyddOu8yk1A3OayQjhO8elYSLiNS
tRsXr7NpsNA6ROMHL6l+qhLocXff/DI/a0Yy84tXv6R60+f7GDt31kUCDIM6v3b2xZdGUcgZf8a2
MZMkfMHlj0Xv5QmxLvG4/1038EcLP0UL25QVdeo7/1q6dW8SvBKtf32e5rNgzNu/LZZSIR5DQ8yH
iFxSHvNvNI6Lq6+NO6rtgvMRMqRJruelyE6bAMcWqgDVohBW1JMnxqTeV/u8nS+m2+TJsbFc2ZiD
asZnbPEcoS1v8qcYlknFbM6klkOWFGeqUhyJ6g7wbd+JCTVloYM04u2qLfB2SzPIsInnQjVlwOt5
5W7gqNGspYJpNTi7BkywRq8WZGJhejuM29dmZ1FugFhADo0CHX53t7OVhVNFMKjigy/xym9VUNAJ
7Fr/kYB6xht/Q6Kl/EHDnXq+pkZy/zJb9t8sylWLZnQO5RrGv/PipuG/PQ8SKf5tXG1nTu3XMrW7
EIttv7IHAFdHlg66+ANKmUJq1L5uunjQ9jRdojjZWPLDJLlAX2+9wrFFJvep5Awce19kKHK1Ox7i
vn4BXkphANnW1bbxOni+YCUu6PfUS1iWJeZSL/j+zzpCkHJb0gNuH8fpmr4R6sOOsnlpEoPxCiyj
jPfik02wBd7iecZTK6LqaFqGyHlEj+xTayPnyKin0Fu0PlQLwL/Rr7iX0Qdeb5qsj5ekqS8zizkq
gPndqt9H77yKmWZE4Uk760i+cKPGK9Pj/XaiayB5wEJMR1fuMiT28Q1lMAsqHQrj2cELJZcy604i
JiTxgUhjjjK0DnB1Pikaa09dZBwB/EYCHjJBXHoGOMK/s/HzOGCKU8znMt8FXs+fadDhtMzhZ/rW
WkNBrZEDTW2V1pk5OSpUWIQAFDmF1lPizPv4yCIHqd7mrfc8/P4EukuPIgucX6//E0iqW6XuPSBJ
/agB6eW/3IVA29ps4UFD52GVfAmliM49TlbQwCG207jescRER6rISH+xw/JTYaZ/QZb2S+ciwCvt
6SSWZKATvTVgO0kgZ9w5zeLheodWHWHfilxhIRU1Sg6JpqY5dGsSS1m0jWV84vfhxNTyMykqNTYl
E01uf+FIaDw9V8wZmWC41lAQs3RbhI4RcfS7KAg/Gru8cWYI/7Bn1LrAGxrcn+fw9VhllvaFoiDQ
e1gBKs7ilYNNgdhq7zP3jHTD8eAE3DLFUa4PIAdjrshZsa/hMg/q84brUz/b+6WVl8cKIiUG7WO7
hp7D/QvAUWaiEopag10+/PnRBpVCXYB7yFDOJJaVR8ww+DbOkU8h2Zi3oJ+HcuxMiMg8n8HNHXPl
a81YiH+rjFeu3phliaZok+2gyAkF2KqeFwNzJpCEdUPdgM50iqt4mnKK7SmYY7eFqhUfIWghz1iJ
TR+ap5GI8lWmIcctjFL9iYt+5bPXp1OfCXZmn/KCvwQWOZ1iTtqcg+QT5RamEvjZyfQpKAsnLGkc
g3Kpw8g8+i6Kx6VgPXwYjaIGnmnCmh6mt5cd8733cdIfpLRtZm8patqF1kuK8/i9GiclDyg43eiL
BetOkenguD1zmYxaYyB/R6WgSB37VWknLUxnfMT6aavJ8RS3xPScZZAXKUG9dPqRUZqS3/amvcp1
0HvZFcsd+MLTrGvpTkXu+db/tTF1tAul3HqnAznjTDrC9zVLUzEkVrEsyFMLw1U0L2YrNOMXSJjc
L1Gj6XfDmFpYVyHITFV6QXGB31Axu7GdZM1n6hSdacJjsGgyaCcg5DRVrPBo72HdeOJjFRo0TTBt
92SH5HsW+7m4uus5uZ9BOtU/HF9pN7/5irD3V7aMXALLpMt7CiZccnBpk5NIhhiwkxyn9r/TLTI0
ILLvywLZnCsjIMFjKfGpFfN8tnJmrxkN0lHRpU5Hr8+tERnQPhqhPxL+txsr0FNA5hyVCKrwmZbV
XAXv9Duz1V960NuSfay2kniTCIMCfcfs0rSMFXroBauFkHG5MXiNCr9Ux6a5YxGsHVu5EfdT14VB
A9zChb6cc2ylXHj5QmvbJiUuelCfvaVzYfrOQNJusxRYXU2Mykv2mDIpvmzD1sCLJADV+uzZi6MH
5b4c60lNwA21k/3lPfZaKV5nHxP7+YjWfZ5kKQ+UjZGuWb0V9iXKEl69KVP0S1cN3bjIztknn/K3
S1AoatZ/qJP3dQJJQ5fpZugJO+c/OHpd0mHywf8DiWtq9E4/ihMunQpysjewyO0HIpIBzdy1me1a
gLYYU913VGa5CcWW5FdBq6JZZ2ah3NvLC0ApHzjdlFHSEMxHNMk93H9hff4BDwSTqE/x7iwyGvid
3djEPbHg1GYxzym+enRA7jCIwlaehDmq1k2bNcibdAsFmcc97W+tdCukjRT9JT/8hPZ1FrXEBRa0
2EOPIa7LzgFCQAvL+f0MPn0zudN3DVrcSf5wF42pCp8rVmeTEhxmizkvK+aNvAK1jNiOH432p+jd
igIoZHS7m9oRKxdqE5kFsb3MVDtdJmR2f2FWYPvof728JYzvFYM/5FlGsyIm80n3uZLIXssIlEEk
Hog23PBle6plrTWbPgTxqU/jl9/3auPfz7t7ojp03p3o6dB9j7XPYw3hbAtOkKNMmm2O2GOiEsr+
hMlE/4Twi25KRT3bjnbIQJMsqiLVtZ6z1gOBRNkB7Dt6dwkIkhPPLE+NR6NLEMZc1Dp0lEj6dW/j
PFfptBCfN/Q6LcxpY4ZeGRGNrwVPBG/mVqanIZwHIBoxdCNGnQeNNkMF1qMVWZH2KbOAS8zaflp1
678bD4eYdOd4SfJw3WX9YKER+na7K2DYR3CD75thkwoLPZf9jCetQoqFxSeP+Z1hDC9tkWQpRtjX
LZjd9zkTWDxJrhLxJ3+5WF2HcZ1/vf5bEQmPKBLoRj3JtTd9pKW09Ahke6Hp1DTHQ077NvVclhtg
zXaRJUZ7UI5QYp8h1u4o31HU9VuaZZxEKxbCfjDJdtHfrXankWzT4RsnuLEvhcPkX2gwQSk4wm4q
O2pSwvD5MTntaxCauAJCoUfkWlkk3Rvgeav06x9MgNy6qEnmjUVE/3g/WNWJfM6fJ9J0l96fYdiI
VcCFXheC076iS9O/gw/SOIQP+CDGVHVt+iyRO1dfv4RM6io6dvTEUvZWyiyc2/CjOrlFX7k2x+9h
MtIP9qRMrjczEYYNDlqCGrehrhLFw2tepSovsD6F/LUuygd0pe0TCPnTtePe05MAOh51WbtIaceW
3k9PLfFKzC4kLstIbXEhEyoIpyJa2EAmErZwgQbRHC4K78r9NRoNu3Hj1yjSXA4mIjO3cxJhYDtr
ujHmfMf4/DFnMGcm+Fx65PJtVgNmqifx5dYfFcbC0h9WpRksbAxUcBq5HlHIBd836ZEi0eSPv14l
SDJwqYmjsefzKUOgS4yruuxo0E7AzF9kZwNqvEmpcuK5ig0SUl4b5bEBvu4toEOnLu5Vc1V0pEnu
m9EaFef9idl19e5d8SwhcPyQl7mECzM1aEMDqQZDvF+pQFuVyf4k/jvoG0FHK6bi80bmvMct11Gd
IphCEnv5cgyJdiQ9pkfgzyPONw38g7zHTk/nXGcVEAZUwJHmaVwp2d7+t3zbCTSUpYNszo4x4888
r59CRTz+knJ9juurd425XgGIQnEO1oToTRSBYLVqfZKihLbN7Z83sFP6F9XYG36wkhPhuq6KxYiN
ZcIa/qW3BmKDxg3Z56j0GIJl953oUq67yotba+dSbUWE0hIEySYFZNNlPEWG1iMD4DB61nOoeveS
oIFQBQ5d6U3+67jEr8YABtQGTydomczA1VRVA5o04mN0EI2pHMcb+jYieHuNTVwWt4MElruBWNu4
GhYmhOxoXrGqjU8zQ8gp4K0br43wGnIrHqNA8vNFASqYYm7V2hFdDvP+gWb9Za7uONOCBS6a7LAK
BphIcGD5RmapneuAhM4TVqB1RUkm6fHO+gIBvmeE634l5ZHKChxU9/bVcUbBXUt3BAQLS1GC60Ph
n4DsUP5h0d80r36ZAdDP0/9tUZgCbfZIh2jS+YHEfakya2nPQKhJZ+JMTzuwNs8+zcTbhmINkrIY
31LvBZqpSC2zUmsWVP5DM5tdx4L2UWWAFaJ6skRICYdIKQuDlqawVlCwR0Uo+xxHNohp9CmlJFau
aVJo+5FZui0NFlUBXls9FI8ouVU36fwCWtOstBSIEB1KFFz/heyXqGj9gEV/LUTRSyzYtSN495/j
dCL+pM5oPvK3bG4eN0Vdk0zb0oyI2V/NslfSVvdcUw+S6zcyOo9SsZX17AxGVAncoVMs8rqvvf+g
/3dihJibx7Wp+id/jp0VBKEzwsF6xomn9exDYSfGBAgliq/qFxMwswj8vGt6MJUBTzCFfo7nMB/f
4l4X1hCG3Qi6cKAtlbne3C2aCaQWdV5gKko9MDrNug/8NeNp+WHooyN9ibjPbUNKTWUB72QZVixX
rjXIG3jrRU5MnAwk+E/P5kDH2icNZso3j0Qmfga8pX74/pzVvj6K9KU2yjMw2lJQ9sAYZ9CX5aE5
4ctCkQx6jSNw+DAcLszydDxQXmXrriAR9SsT968NsUPGflfe95hnbPAs+e3SELLnvi2MxdFwI79I
MqfcmJq2/WWJywNwOS/rjqbX82txTJaIUIcqHHTm1yyJwhli4xlqBez9MMZI+KR/dzFKWQwYIHEq
4kKMpwSh6rO09jIDfN86PwrLvjCUr4VYFYE9cRIGzjqEqzV6ZkD3tRHIllewKaKxZtxGdVkOC/qd
uMfGESvnMLZmrgOxp8c5C5Yrp4g+I73OlvvP2ePL9m/0UWbkWsmSFcFwH7W29Ye6+SLI4eD3mr4W
Mido+Cf6LpvT0cMH/Ql23r4KAkDzjH1R9p+HXQUtXkpN7UdO2F7OABJG43mdcClXpsNevheIDHM4
TPirfUW3ZXgFo+Uk6D2HzACtZXU1HQ+Us2CQrchTb9fcYQ3F6ZZzjya+x+EsjT3vnuTwcHnuwXFD
IQDd8U5lu2svT64OjwhzjUtyWxyslJThSvvks5xV0zMV9CSr7phO9SqKLioVOBIp1j3PB32u2D8R
qWRqC4vH48PVbSti0XnMXVAr1rAEekVelmFW/dphKOa79B09+G9ELIXcgZPVmRkaPiuCbCgy5yKh
j1adIzb/GANRd7PAqCrm5Bf7QDoonaQ3TX9wC2D5jNCu8bOrcizsIKVUtYIZQVWdF7JpxrH3qPgX
TfPEfRw5qjrUT+kZIStDb4gChSF4AWFD4OidMbGfe1gJpwJlg7FcqpQK0Q5pPPGHB7bGL/lfN0na
EL5TdLb4miheiMXHMMQ+t302ke6SYQ4WMuzzVadCbBT299vhmcTaL1CsHLZiX5Zk7mHPfqxGV1er
rix8D+s3w5jO1e08YC/544tbJP7xaFjSg//87go8fLlFabi5LPYXVMN5qZsDSkfMsuwr9exVPePa
9nog/lKa4hxux9As1ol0dmNgWuhKAHFWmH8hCurLaTx8yn7jL3bnGdbq+EYuetZ+o6ywqBmAwxNJ
WZUc271oxSLMQc7K5SxKcNM52fSRky3UFcsgHvyeC97OeXriRgMowwLWKsWYDeIbVsRu8LEYxQ8y
PA+p3Y0xc/FYgGvoxjPLwCwfhFTW/X5Wr3aLnMvHZklRdY6cYKSbHMD/3Tl2yOGe2AemsGrXjOKS
2jn0WGN1mO+VkpAqyvkm0Z1svT9Gr0TV3PB/zAovNgjkKDE+s4FVnt2yHmyzT5VVIOIju6Cl10ot
UfqzdluqI9Gape0TjRK1QfOtLCFv7b2Hd8g8JcsRZBVOolTyyecO6kdOf3bw63R2aRUa0iLAEnVI
LaZ+FHQX9XQuRldzk5BsJvIjpYPrSXYHoeDVUkD5VgThpz+Q41JT5Vf6Y4784sNF2V21yRWC+JtP
Oq1Wni2Q0KsOOGvtOK0cPtdFqNXBLyFyV4/6uDDYr43KOeWj2f1OQCR94tdzCfWriw3BTIm5quF6
yPRYt93MbXGG8v1noxdQ+judBOuyaPpxjhbEY2wdqtYWjxYHcvrrXY8jVZgAW532QNVAfVFvhjr4
rNSVSfDUuexHzBkDRaEMsGr+ll+/NI/LGV5sSEpDiCzQHw7dT+zdUQLGhbAsfF8okVT4UPQqV0j0
OXkFr36ZdFlxmu4TWVIHAl8lasrGlROvAhPjPH6x3bNfjIhBeMvpwhR8pOszLluXmZE1YhdzL+ca
zUd3wpq+CNyO1jyURIOmzYH73Cl1qR4gtIMp9GLAjBqWWCj+qPcHcD/k4umHBWcmIa9AXRZLhmXQ
Sy13OwHEuKSXUY8Q3cTazlDownkrAKSkJbkv6iZwiYqe5vAfDvMwWj4bxeclziB38AVHtPcxc+NA
Z2AjTLv5tU+gLvMehfLrZQ0aRnOlDx4ANLQn5KospPbqNRKhkqbwWRKy2GhD1NJsktnh1otVVg4v
arQMe4M/pG1CbOwDcIW2Bulo1Mhx92Kb46Y0HPlLOLFxBc0IwIo6JNjlGlp3ZwvoIvy7JVRWxqY+
R7FHS71v8wEHOyDf30M3aKTCjhcEe84cMe6QZz48K8SJFbe4aT6aH3kYwJLYOEfhBXcE/3xWjwjA
gFANNhGhxTrPtulaga1caCl2PE7aSN48LanVa7C2DSbgj2VmnNS4oiFlmVVD/rx8oDE5kRamaVK/
zHcEKzuHQWu1mmTGlQ9QjqgR2xEd18juTgtLwoZr6OKCYVvxqj5ArKhz6UkcuSo1JXyfLgb8EWRe
gcymlProoWFIiDOOXyLrgTMWKS7ClT1c3r1kWNS2CBpu46e6tQ/Duq40vrVHX9ZAkg9b6aiANxMQ
P2j5adv1sF+HqTdCoQ6iX01lCKzwTPyOgx+bQe2VSo7neSwf+GRoIeRQ3P8X3kvfvTRtHU3frJdJ
lSvS6EJKgpbtz6YU7mY6D9iBPwZsphsq2iZadIYGk+qjB4QGqLqvDxdPpAPVfschdyD4ZmsWBhWv
zcrZMjRpHUmhBZtD1i46ASL85oNKcqSB3zrZqar6vZzbBrAZSghNv8n1ynG92fMTkuZNWtqY0UfX
DV8AWUQpwEHCvY+sYFpugmIfcDpHCNqLyJE4iRZl8IXKNwqw5YNfnSc5mgbepY0vB3l3wdfOTHWt
BYmts1IEXAuLSTVAQh0TtqSzw68USfVnQsjDnjiYzHxemFKIeZ94RNqOjhbdH5eB9vCWbvprJMAh
nJoarkwlitZ50LyGHJw3fDjqdpf4GUnqpmy6aU7ll3s5qRsMcWTcIeTnBUDZfFCW7jC94NpzZz3L
ALTntNLWQNAMpGbRwEB/fXe1+M6jDe1gs+INievYJkWnbIAwIVS587lsJBXCi+DkI6+Dg9FH1kOU
QUducvU8kubVPIx6gL0iPdAAep5BekWSlLWToZVjl6ihq7SdwxCj2NwxfZGwzo4mTcAzj7r0w/cA
NBePRC59r5OINxlaiWUuR5I290boLqfOlm+FJ+BUMCKxWv2d9/rEHR4NYhRdmi9LfawmcWpdaura
QsvjMqJjJXGKqD74B6rX02Ow8maiQ+nTgWK+jAMiGdOZv53AEwmFRO5POzyRHVdWW0K+Avh6tLxJ
vhkAK92olL6NZRMh97KxTJGfFVt65eq0aRNAQzAfzMZhEo5eveBB+8yQNAWr6V8hoVywKKIrKPct
1xEkb7JFiLNoOseuxdRpNly5Gu5ugSCavD/fWl8XqW/W8vXKLzvB3dgsKhqY5t1B82rjNuwZHDSI
Licv70I8jtJu12uDYobo7fzFoyXay1XW3tqv6AKGRfvqfxd3zPlLm1aFUPPSYxHnjdKV/zseiYWN
43JcD/P00pBkYeS+I5GEtW495jmPDkB3vc4i3gnZetVCbJnUOC3g5mv0mjw8/uolKbOL7jdA9/Gs
W2uHOfe4k3oZQauprqVGuppPMpZUH8phQKgx1QE8KQ4HhqJVoY28nsOjniaBZgJPUhuJZ0U3HnWl
WEJ1blH8Dh5hxZAULxAWWSaB/SePiYu8T4uEmKDi/FZACQC9lCH6Znke0wu2ygM3FHs/Z5M7sgOu
14c9kuLv768Rdz8ueWC+gVl8STr9jD2ZNt5JOjOUOx6ceJw7tpD/iEc+ksKRRLe2PIWyC8duiCJP
SnNlMsa5mZTRoGCPcYDR9OY7zamO0aMwGb579gravtMYAi8En61hYEMA2I4lJRHi84Fgs+3mtKPy
dHR16ZxowKeyAxY78638qwoIRTZMHqXqiw3+PbemnqwW3Bz6TtoM8Y0ncikzouBoPgUslDx8jkgw
F2gmWGTlc6oi4z1emHK80QgBWp2Fj8Htng5wvjb21ZUbw1teltTWp/kWUFFhkUkhDPwGyU89ARaF
cZmps+qrtcOGZ4n9SyFWh6RnBTeQHlTbt7+1Wc9DFBOb+l7Kbx3dAQe34KbIgAr7nzJUrx9QvdNR
C+5Sfi5T5aCVcPrQwA8ryPZMo80b6NdM9tnLyitnTcXIjq2WZwL7m+XA/+j3WLT1eZVU38ykZxMe
xXtOLS7kkrp6bGph5N9BzhvIQLZ+RQDqn1p0iy6FbrHdonyQHu9PT+Wynylq9/vV0HQBw3jKIgMt
wap/gsZz8lte/XFx5eQPAw1ksz9zQxwmPJMEhH9SR3Ys6taCNfGV9JQdefwfY72e6Mp2t4vwioNM
DzZ5HHL+owGdt8SD4+IwgcKbjlXkwWC7i22xe2Dh0LV55gz3FPWU7w6y9bPPnWFE6Yo3Bj4/1zwx
3BuK77wdqpx+DfvXxUF7hbK9lABi3q2ZwsmCNmkWCUzFDe0NBu2iaTsJOW8UGrfJHxcJJcXoAV2g
rIRPN1B4rONM11X4YpH6Sj4H+9vUmkuO3M3Ntug/IJ3xM2fhZJq4LJ4t9r5+/vAa1TgdOjwvUqYq
aKQBIB1HMdB9Vm2Mc+lNLUbbERhTurp6Zuu5ZHpUBVWZYAwVS0cmbcbTr3Ucq2ZlKcyzZI3NN8tq
DHkF1XfHtUmKE5+i27OCR1v6odraXyHEHciZaQ1ZWwtqu9D1TLB2TQCC4eTtz8dcbE02aoaiulPP
PGmiLOJA864H3INFT+74hXSV+/t1Cf1v4Oi1nD2EZsrGw11lDr+nb7YvMfwEhBNqU5LNpoqalo+a
l4mZexGBNMoACCay2sun7H6xtE+3QE+qMNz0ICQHlQjO+BYLOby1jUiTeKvzJeONpaqf9YNfgsrB
vwy8tPAf2FQibbRFpFL4VLAJgJWtXceLYDxBi/xfL28YInZqx7iYW6Fvq0CbFPXPbD5oX0V4rfPd
DFsTUgfvi/wImZUMZDH1OnRq1MLrsl91a/p9HloJ8lPxLaR2jsB4cDAVj//Ib/2b7+eaycKe9yNh
TSWy2Y+sUY4zXRLB28sezUp8JO1YZnbcl5O9ZgeWlRw8q+YCPEgarbXiwOP6wKwEvmckhez0XBn9
FbuJ26YcCs44LARwJu/q21wV1Dy6H9urw0QpUMAskpMFV1A5LTOsLJyJi7sQpUyFkd2IO+qOCWKl
i++90MJL7vDP9wJTgKCQqmdWEg8TdkhMqyQQ3PT80MDkyLolLAFMgKISySg9UhMaZFeeMWoyKP7/
GWXf02dtjbwH9sOrIjdiLKuEt9GPngotWDyTBhiez7vG91khDgU1W+g+mH6CKIr9EPkA3mPGNeAW
ou06pcxF7mUEN1WZo2sq/dh2QXwfxLESqhI2g9yQmqPfsCUtXZTwbkqYx3IDrePveVeFYYp1FMod
RYzrpAECE2zK7r7EkjrHDDJxItie+2HZXW+Mcz4iJdO+E7NlTzY3uRMaoY6YRf7pgfnZfysaXTtK
jT6iiig53qU9VnvVfE3sa/axa+Q8J+ckKoK7Ga/FjJ51xqUCD+OwCnXnn2YAWGLkslbq0j5T4TZX
5bTVbUU0wwh7iFFYmNEaaPXOMvcqA9rGd1naRm3WuQYyhbBZ4P/MlZ+GMLKDTRWoZqSPDAzvQVE5
EnrLwqXuQSKlGj9DZsza3ugBjLzl85t48ONwlI+HU8+ir2JmaFxjzmaCOxgPCK7pqwP/2ZLbpPFa
oedFTLnu0JnnkHNuhvUnFukffRCb3E3tqmEs5SAdWTKD5M3cVLfEn1xIxqQfZrdWtQ6Squf0BwLM
fEb5e2bQpD2pSpU+v/BqEJLbq85b5/A7nKodCywIdcW9X9PKyltxfhH+Va+AHUBqWryvf3trqkhU
Z9GZK6NvxKfNyi1ybTZ0G/ZelNYzigT8ytDLO9XEhI2dT/gow65CGKjKfKuXdacFEY3zA8UI2quf
RAxnSczon0gUf7J89+Nbab3fu78M+gCOIBnollGgqOwqOchkkQ6zarWpc94QwHJ6i67BTfmAGWJ1
vfHVlyJ8g/KJHspFKaXQ+tn5OFuC9HnF6WX21jjcjsM+sv/fvaZIzAq5g0077hpKcj3PVZMURNr5
HNWvsB/YBGTP28ZVLJRq/8Kpzg0n9P6VBv6ucoZ9mylVlfT/XL/pZuSxFT0fz54H6JTLgeFVDlQu
At2KucfhWsoc/q2gER0G4ZtlBeZvC8hS7V6fq+ThlDz4Ms/6hiExN5Z2yBhDttnxhLIVY2CW09v2
EFQShUQMU1AAwWLHwgGFG796/CXHl27n9H4PQEcjRdlSKL4BycHvAQfViiuEJMzkPGiXrIwc2me7
dnrXSt870GtJC0Ar5TApPQU/zG0fGZtw5HBpp1b0+dSEm1Kp3imtiHdB6rZ+s3wHmEK93FjquJ3F
CjWgNgcudmy7gAqY9zw2Z5Wh+bKwNPKBTGfllssWK1gcReNjRS58HmgX5R529ZQanRlQHCNApmNb
cdWG/P3qYLsNpTFdYy8W9Udq60LMzNYFklK2z0ICwFbyAmV4XDCwQc1WznB3mlgh89mm3FVYiSIH
KI4IHyPOpNiGKHqG9/emin1n7BHXFFjB7RYFoKIxjocMPrXlqSwig7LJuGw1cilc4m3KTL6KgC4z
0gubUlmm71JDUjS3/sOoxds4oKiBD2GCtOtr6dPH2nqapbcZSlZCEtiqMOnQsaGUDUccaUNDqlw9
gUP4F4AFkF+SIQwTYeZxRfcFa2G8fcwFRbpzT1lQ5ZA5OrARHGVorzLhznSTAKcSQevSrs77Bb5n
V4ZWzio6IU3gdi606mC5NboSOA3MtTQ87+Yj2qcmgtDvcua+0VRGW3S9Ukf7sdiVq8HithIsixvZ
/1ZNRUqM51NkmYILCouDgWo2BsjHIvNhhylb8rlYr201zYFydd1G3uBWzFfmX9boj3/XDWIF0Klo
vmWOCCQv+d3+0JjEWhgBsyykwPgSoPJeiqNhXX+IWMhhKYWNNllyAcBouEEeU3qUjRd5AV6fkXfn
lYV/x4v8WBnHiaODU0umnoI0MbN1tdtsF0Y5wx68oqpQpp/2rCDJhTRYtzt2yJhEI6hAzvNdc0mY
bvNseeS8CSL8tRML61NMY4izv0Syvhns8H7j6ZPvFwCwXNEHKknpaX94U3SLPaeOWTgaLhThseml
oJa1/4UDQKDdKZdH44d0deFSzqluwwCb8mDTz7tH/7L8Jb75oCDt6DwetRJDF9mxrEHb+A+4TCUv
WZBHIbH7bQ8GOnVCQt+5Vq9vXF+0fsYtcPkkBppcGjCFTGc24dSiOXzKRKQGxSQywyPCaPNA7jhO
azigXhdxP2hP1WWg/x7GirvKs4and+H0x7NJ59reAK2Jppu7Mw0gFx4ww4tdChffIxt5rrbG8b9B
i9nxy2crMwit9yFqbzZ97pyH6cqkjyUCu5597PBKr8Y0Sk8xAHRtwKtWlKf5v37er0gSSQ3utL9U
+FyI4ySd6YBOwwrmtybnLbjUAD/nsSvApx2Fw/vccicrqbtLOOfxdvswZZiSJ5BG1JCzMqm6PoU8
Xfik61Em1dWmQJeRBO0Qez/6ENCPMUmMTuQFUeHdb4AaUpUvW8nmq3f2Wy91rkZ1gb4Bq0njbGub
SMqexv42o6sukuN6TexO6L4rczwdbSGzmatFpzKlGVvFDPH1AyfzDYnsmGnEMUByVjkd810Uxi33
YIqcxRVxM8wjkdST6GFMh4oNyeYVMkB9d8zUV8LqEVA2H2wQFiU5/gmQk5V+gFtqMG/uEUn16rJd
5+aWPKKpJSOHVALuJMyrce+qyIVmwYzsu+xYOdQLSP9zmsY34zXnQ3UYhO+IZN96lE4R/z4B9mfj
YsM6bxLOKBFRRJGv3vGqtyt+Sz/l467ay0Qag7vloltUXA7Kn1WLOTZJQAvBPOid7qUlMbANLYXP
RepEErx9UZO6OOds3EwgeL4M+5ynWaLZYyVh19dUDN14GpAGCYMQFtov2jIB9jFQlGz1wULqHt/9
kXvo3L7/aSwIfv/n2QZSzhPx6K/raP/eucJUd5mfSR6jyH0Xe+6vgiQoMkZKAn3o6C3DlyMEh0a9
0bDgahAJUnNnGaIrM6aXN5SLusHp7xFo2KqAFXUi4TByA6RCFpdOIKMgoRyJVzDTxPgzQGncpQI5
sOm12PBkCq3BpOTPcryLm3MJLc+/UfT3RCIXpyd9vpYpX8OG21w8wmwWbVYg9CAatnz3jMvbJ8bK
6dQ69FGdksuSTBTGjskjAYDn/U/Rsv/36FvW8n5a6cnh7OxH5ZuRi6fSdz+5Z2dQLn5hxx2o/ort
E50/ib4GDFyyRstDtGotYwtNcM3JR+Pa6eZNfGWjHvX1EB9E7APcNh4s9gf89cKYW+xhO6FYQQyh
iVXh2bZm4XnwmDm/vdUfeOrclRPVCBPIO5dcR/tnklM8HFCuuLLb0rEIpPDaIxHAA9xskk+t/6vZ
EOC8fVP8gw9h147dLh4LYgmPbiM0GGhzeM/i4cOpCQ5CE4luv1hdpMhUYJkOYYs+fZ1LVinEFGoP
b+0KLSrKDq+9SBy0aFDCLE5zIfm8hoC8Z2I1/0yJ5JYo5d5lHJETKbLBh6Qds2+DgEn0KjXHORFu
JN8W3O0Y2xPXsjsetsE0Mg2VSmWfDlCsLgQV4LZ7I7bnwUdatK7RwaMGDPgXsrZyb/hXkEVsA/8r
YLjWRdpZ9U85EQhE/O8bIxlQ+q0iyn/oVEx2qSpwbjLXOpXLR2d1viE1vU2xR33M+p95N6ViuWM+
SsWifqPOrZEBQ07UUPCkUmoG3VRtAx/esrsVcLDJeEi3xPD/3mY66h1FEJa4xUeffvZhBx+GL3tb
fEkvHo1/7OsrlPCnXGtQbn9l+u/tm+2NlSVrjo1PH+Hlr0b7mm5tX6tgkELF8U2A+xq+wwN83gYt
jNomUw/bwbewbdPtK9F/lRxyHtrRzHQMCw9AOjc2zqUm9pRh37PTJ7EEl26Y6nkIB5IAaEzpXujy
opl9B5pWeL71ZF4hB/jv8VZwuBVIDsaizt16pkB02iQyO6I1VDbhTTNC1i33hRd7myNXC58w1mC+
NV2CLgfGw2Ka/vKcEWpStoEvmd5HOs6X2D1jIRuZi0PAi2E7uC7EDJwMzgTvbcarVi0+T9T+sGnP
RRGOoquKrru2yVrkUNC/6FtR/Svcru7LRzn29gFfjp+4Kl7ODcvjQd5kS3rhe7hAlHMAuYJCDlxm
C55mDCxkvG1Q2KrR4uh/j3ohYxh04E2GjWhIx8XM0S83Hne8i9LvWf3NBurGFbb1LZBUZ+wJrees
zcJ9hq+s7qcsvbAbyOmVhDxtdMSHQu3ENKe+WjYueWfqu+6MUCcEwAsm8RSEbX5jEGo12XaJog+W
KAH7HVbg0kINlKpcgwnW0/eeNA1qFMyHfrN8KLovImuEUGJERcnIaWGld77WS8QVPAZ8TeBw+SK9
JbhfhuiJ0RB5fRj2ghgS6qf3VbpGNy2m1HxWlp+DPzYJoJ6Mn6MTg8nFyMk4IJ8OgDS5NgMoJXlJ
jEALQ/aLJRcOHC/i9zdVxSFsG0pfxsbVhr65F0PIW61kkAKJYBqfoFsS263o9f/xvxRpTUihBLRU
6IeXTZN05SBsxcJF4O/VNJFVpcF+qsEdUgRWPNZlFtZAnjKh9yIeCyfNIPDgmrbt/S8MXSMH/bRz
Rs8cEumKja9JWeDKl0nWzprg0PiQ8EEkgYljUNlXTQRiBivxFIKHF2gENoWLca+9rsiOu/lysprM
YQcqAMM0xzn4EmHrKQnPnKNrKD+1tbSL0cgDt+47n6yjtnjbh23TMAPb2qiYlwIG3Lb5Q9cQZd+Y
TvEL9G9yoRag/6cHxKa1pEbnqURPBsoEG5yna/N8aDTvJP81d/wU54IP7lfEqDVfYqUIlbkd0T01
h7MSwXgaz8BonYIvQWuS2H6l84GdMaTsAo9ZWxhKic0mBHYajCnESNGq8II4V07n+zp9NRymhCck
yMzbRNeGMrlXnpq4x6OzPgPnMQgUNu9wFqjsFlv84QG5RxMlqt895CvLTthRN89eC/ZnrsunjUTh
2q7CWfu2sDL3zaupo7u7AkAmH0gLWt6xcGSSMtneZ2AKW98mzWUeTRsBFaSUCWfJhoDheULU8lgj
Jaqf9sv8c8YBpRsnk29mN8DYabh0hL+JEAtzjovxCrcKkbB6cmnIsFDuUDOBB/NQL60K0R9l+To7
xsOeUBWFmyhdFXDGxNIWR51YaGafYeRKYDcma73Hv9yq0GBWQmQPZLWoD0Q26dlnHKQrz/z72ugc
qgaKuvkfiAkY89TDc663NH/eagvQZHHjbh+7xRh3FmEk145b4GXGMzWHjn0mEvb0guOZW0+C7KPe
H/JQdtsfgP/8Qw7vn5SeLHl+mp7kmd4CAPw2iOnJvcsGvD6zQEty/bgOZWe+dX2bpWZmQiTZPXsw
ZLKgOnQWVrF4GzORFEw4AxEnj9rAeBo7ZUGbSE5nmW0lGSBJJlkYD4iMVXaK/idKcHOUIrR0gV8b
Q4fkzkp9qn5KMSpDgoDDHFuM4CZ34dqgwxmSxx6NqWC79Ii74Giyx03DRZssnsZz/QfFH4NO04y5
4S0yDKkogmWKkdGvYHDLQGlGtrnXjnAKdsp9u/NQyhrrQV4DJoxEN4hXI+3vZphKbZ9BgpoJxQpK
2UJnIZH8QOzjBG1hWL/GX9hDcVvQ+HHtcGvBxRT/YdB+5lC5bhXr/sZPLCQIFnQjFvtiH6fHt4CY
PiNZTi5Wnbn399frvzy0tpd0hbtuaL/IPvX3UhZjO0VDekvm/6KY6euV9xXRTQqCf4rcBuqjiZeO
0F0xVTfJRZjNmWKc2jR0HRyba85qc+yhze0B4UMcJoSbYgVIufZlzNHzPFo5v4MAOyd3U5uSHUP5
HAYT9EUzVERTaDa6LTycBmQLePZo4YmGJO+Hj2OHXabzorqYMEu8OOnRsH5JiBO1igq6e3LM68wm
rGMhjlD/8eTFit8trfLdUmpLPOe+rmGNcOVWm/bRylZXfMCV9nJc2CvZVAlbsum50+lSmNIPJzSG
S5MaxxsuR+XpbyzRRWSEAA4sy4puLKCR9g3NC12srrT1U1EoJ4CJUxSGmL9QJkNHYODMyO0J7YwU
ueKfhXGgVDNCtTGWYb7c7Vd5OXd5GinKfi0/475O0yoBp9Kuoh+ChIF2Ba1hlxU8HtUQ55O1reUR
Hu6VtIr5o2mompDxGA8yjv5a18Crbgb8Dt0RcaU1qMnRBZMOJE11SbjYV1PVKXxT2qzA/r/FB7lU
ZZlbrq5VqIpXxUaYXplwppzUWF8XxJiwYa/0lfS4JBeBAcczJBsMXjo1C/WuMtuZ7QsGh080xNG9
cFDCOd7bNBNuGWA9pE6FhQhWrot7ZJM7y++vaMPbZyv8ahdj56wcK3BzrJO6mrR1y+xbrh7WPkUN
n0MfJJ0JRLXDqWAgEA+0wlbGYwdj2YdBEe+G3mY/Z31pQ8qe0vzBs3uOMLe/Dmg/IVBkP9pOYTca
Rzi2v7x4kiUnrfnlfAf+UC+UdO/p6pN5g0hob8H36XgDqE2ZKRjWiWwU0Rbx9FT4xUvHVJY50cQb
zbQIwrWunkIVPMchOzEd5Rf7M9cGq47ENCh2/pzKRtIBSlpUpNZtIp98n7CJ3FqkFp7s+pJBT5Rv
ZfYdtQ9kKFRlxKWOzGEfzePJnNeaKIMBz4HhyVesg+OilmvnsPjmG41NCMFCLGZ6pmCnToYthbgm
bk88pVYJCHDrz01XH/1cTE8EaIupYu4NVcsb1VDtm++hVBCAvGZ1hwRxK5SpmC6J+mtJCyxzu0MF
7/wkyVj8Fp9KsfCrWPrhz2cPErRqdGJKKgWD3Kcp4EVfzlkJbF/KLx2Y6AUKl5i6iBVp8U8KGRpZ
8W9aggHN0/mUEjHn7/blj1kTd0a5pVJgTveHiNkQMCudcv+zrEtdKAR/0KS1BN3OCROGv0aoIiwj
bQFNEHCodpF3x8XrOFYxexHoHHvJkwpHWoyAGLC4NxtODfW5aHAd4/TO/T8xAnhXjrfEtJaoxhbi
YluFoI6rn39b5yHuuvIUc/o8je0VJH4PhH4deOp7dFjh2hKfTKHWnW4I6M++7H14omdB0lXD0U4Z
PoRS7x4KAGLGHdb2+7t00xwWKhBeIPwrzQRqxRufuELhV1eThdZZj2qRcwoLtmAOCSduB2rTUfuM
DXXiZgfJX9aQIX7tZabiakPKp8xU+F4OY1F1U9r8SwwxF3yyrCTzEbsaP9TKdLvznsuIAG5uKIDZ
FlvtY48kND2MEVdke0PmIC+L98qi1RmNAw7uIiRq7pRHsmTsCFOxz3DWVhRZCKRGu8pYsXspJrv0
9Psnt9rvrKvzr8zD4VGz6buKuS+ts1lm/+KXgnQCpQD5pU/UjC4CyU5LNJ/qA8TzuRumrKZDCwXt
tHbW6Xsyuonhy/ECVYaK1QZ3J9eC5RI0aE7v5r72pme5kTFl7qxu4qvzP82A/qQDnINIv+HKeYFw
yu0wAyLGsYiJbcaGu/AIS1LTWO5pPDKp+rlvATQ4aFclpjs2fA/CgVEsPhu+7kFLgkpJuM0bWn0J
Yesu5jL3lhpAjCM7L/cTMii+0n1XGX/YKs6ustH/Bn5DbafiKnN52f1irf9DE4nG6cc1fUk7fTEH
Oi+UsNeQSUN5xGSO88BTCfYaWFc202drl/OnGmVfKmXF8ngtJ3owaC7SEqwQZvTzlCY/fgNY/YbG
MwwZe2LESFcbwuVIvaLiAeJDbGXkUSzH1GxXxKlONQYm4ZR9lrlf35xg5tp7+jb7S7TT9RZ6PCNE
xBj1xlZas1sUQZA0BDD2fk46/KrrsPbcHRI1VL0bRv2/UQTXWJdukla3WmB5c+j9h3LAczJEJTIZ
Am1ZESpdK1LBIebAmn6yCosH6IdobssXahsLSOZEorIgqBSjEaXkHvcDbvnIJJtEi8hxEkq+rtmy
qAtXB8A1/aVkZ1QcRcRe6DyQxEMEnrYKMi3ocwbsdEBYDPocUlGEhT/o1iuJJxIcfEqg1KiMF3L9
adxQRcti5gGGeqI6oZ/ayYvfhw4B6XljTuyVdNcY6fEei3Zz0bLm9s5oiLt8UmdBjhAuI5SO8s5j
UjfVTPkKm/XYwQON44VcWMywkzK+SXJPA3FOzd3bxsyvgev14+7yB8SoMUZ7mykSyZoPkFQvJ3JQ
SzWiqjcFA5WOnjmH3yWBz0LisashiRmQw6Ek76ZR5dH5ZyugtJ11WB3PR+RxetePUPGcDQjldZS0
gT652qlfb5hHNaqIJM3f/IlHwVoyDBj4cfDrLANpMa2N+PYXQF5lfqF7cE4lwq9o39Y2CHwSYBLH
ng213PMWbi0yhnDHuZElhtIdgXHUP9TxNBG4xUdc7kdkBT/LzvIbXUtWs03PH6nDK3XLHaPWWtuJ
/EActmFdS3ylDYbzL3UgsEKY4bp3J2Gcs2RH9ksQ/VbIub7Xnh58r1LkNp4aw33yvCEAQyqTHNkm
QPdwiY2So1OGUU0l2R5DVvbxa5c6Ep7zC+lRPYadIuP0x1ntiLCSU0sqfAQNJ7a5Qtw/0n40Uke4
2cmMU09VeZqwfyJCoFoKqTdK9+BUDejUISyT4KGjwDH/T0JtEuQdel+C+nPTpaW+1NDEpIFymZSw
niadWoDAP641m1f2p8wXCmt8Qaxb+Ledec4bKN9WYwJ4Qy6tdMwqearj8IM9nPOmBaEx9LA7oSdb
aclbuMaZDMvm4tKhBCRq3Yy7pibYdCOesQ5vi9XrNz9XxHy8CEWarDA9WeEX9aDcvpoqaDs4ndcb
TYh34WHs4ECkGdSKkgNBGhHUatDRPHFhKWik4i+tonE3rAnavTbcEdy579iZKjUgnFb9SbS+7tXM
ke/qcl0YMA74jbOQ4Fazz7Z9yY1jPPbS3dRxhS4C2/Wk3VtXXBifLm5Art5jYSXpcvOz8VP3Il9L
WhUYisIIqlQizIjCv70hXlZ8CpuHGMdUkOVHVf3sUlEYGst/ccyb2Pm2wYYTekOznLL90ABA0oMf
IiOqBcJPr0ZdGU/lhUVj/BNCym/6Bn8qNMgtAwhh2HWA9xJlAnEBdrANwhbiVOmsBmvwcK4GR0Pa
93RusxWn+3ifaH30D1SvtDZh6n7OneXymU2E73Z/fLMJTUueiv9aeApcv1LYPXX/eC5DHFoc+vw3
s47JDtfYLjwTsThSJNmR5PZftqQf40lon9Om9KdFAkGQdjCNHSXay3nGZTe8NJfR1+v0FE5fBhr/
a/hHAnJXU/Bthg09DVRXID4wv3Cqk4bfhz3hwV9AaMTHXOastav/527oVPWN2A1i/peeS7JuFO/c
kCcaONMAQfyGCKaH60QrgH+j5EkRRseT/LvmSl3bYZrLh+ctqM+1FVAhgi87JJcvNpi/h/+zaPwb
n7Ry6jl7yKBl5ow8wsPpYIQaJHU+1dV6t1LP7eysZOTmx4/89Dp6CiNmv9/eEdhoVWi2zfzNhSQQ
+ia3EOnRIv5scRrR3/QW/AKVArgybOdJaDH1AhgYIbJk3F/bBO18OcBxcrhG9cWo1KRQsYawgr6t
08fLtlEf320nCPCxvHYMJhhhHG95gRMPZziX4uPOuyjKo3ANqFtlcaX3HXi8x5h+KLvPP+cZ35aU
Ypv+oODSCjqv9Dk+cxNKVXhUBT8vTqwwjJSv7JFw2IAGMnh+vnOW3nlswLXetV5BdrGfHuV/D2Tp
ZnoZpqWBqBEc2yhk3dWWrowzfx4H6aOXRoL+yzuk8GkUyS1HXNTtCQlP4vyGUgFJznJzxH4A4Cxl
3in0rhwgYVQSKGsUehl+2GY4YeGTu02XfHAr56Ybn9QeY9kkcq8EqhyTfggWXNpiDxB1AmcXyZ/q
cywt+P3Bjx1QLKGvXzd4x01U3lcVIOQL3lEwCsTJ/P41rBlTRfLnSQzCkD7cw60xlJAW62D5h60X
eKE0FnGSEItkl/osjpEtHtwQYr6d/e4fe4OYTr3IjoJnRM5HR5xUd5evv5pZhnIAUy3SONOxx4sm
jCg29MQZaj196AlIT8kbDPvVSwZZ5Nh05qiwDEr1o/dxAW1UL/bjrsqgfPJz5ENm0hQ2GuGrrsbZ
j5KXww9e16aXgYRQMlZ/fIQpjI8owcs8a29El8fKvK2BeasCyNbZuaLpaq+9/fzu8dmpdTkdsg6Z
Jfb+y8Od0bYKVIuGMdgl0jy4aBxjvXTH1httlUoZsnJRJOV9XNEAL0f3imP7Ugif1O5OKIqkC/io
MH7r0sVNAb405ulP1unjc99U5xZKBlbQfsRQ7MwJ8Jpl8bLR59XP/zIyy+JxYpnbXeaGpH84w7sW
lAJZHh+VQO06+VF2Y8zpR0pptgUJQ8BvAjsUNDwIGpflop+dbFffVOcggeBSOlQwUxMC1pVP2sVi
+Qb9HSMA6duJgWgJnD8eBOCAsDjmZg3k/Ld9CJ45p7qPlcmRJ//d75t863ed7OnnzQVa7km4AWXa
GiKVl6EE4g90Eov5uRvOz2BSdCUwZA6WZMIcGBLsIH1ujjMD4r2jxh8cjB1oaJK6BVpGfuGT8W2S
5gX5CEFFNX7tXWkoPhJt7zZqUsJq29KeSJK+ANCH9KM8Oz21yC+0hiUwbgr99OmyU/cYZWek1qXX
Ctsotg955R+Rnb3TN2QKsaGoi5geqPUYiaTwqEaVk4BASBJRxHnhaPWAghakexZRyuuHFYA75k9R
CDTTCHzRnehpBrV5fitsAy6mVH2PPhic8a5ajqJJ+PtnugIl9VlM2L6y2p5XLnFSlsGUrxOY2gZJ
dWm3F+IvBx4qpVjS3M7pmSgitoLbR4jOAVl+FxGvbZd0LDwAAzi3zqGJFaU4n6Oy75y/XS8GZJxe
wBrmcOib6vUTghN6y1pBBb0BMuONND0CNOPQa5iFpik5BfRBgvGlr0oFjd/pyS0cA3vVRz6xEGzA
GuFuKNE8kEZTedIBZpga6CJKXNz1IBP9d8kv2yffoN79KaZ0XEo/YAZJIygI7bfhBwpsX2lJ72Ad
skUlYaAT3C/qH9GCF1H7xsNrRi0Jm2QvzgsnElLcomV5ux4e8tZfZ5PzAsmBZz++bOsUfcXDheoz
wP+0zyVvheCOmxQr3d7gF9RCa4p4VE7Z308Ajga7+Wb96qN446b/OkbBwUu9dm0gB5d5hQBDyJRM
wY7u2VgZG3oqlgFlQklUODP2XFVDuuGuWAG/xTis+Sk71/rcQ/yRAYc2rq2uQcSI6FNwlIo21n/m
pFHkw0GVKIYusGq2PaQ/lAvX0aXMFiGdJNlSLnnxzyELk/XEJl/poA7HLbTsS/jq1uVHb0n33ca+
7b1VWIp4sN6yghIQY7SxdbkOzjAi/E2GqI+H3Tov3DR1MxbSLz9DGwkbWPkb79rv4HYm5Hz7Y458
6wMmJl8viMw0BkpR6c6VbulfSxHu7t/XTqQVz/o/sLtG7f/8uPdkEJzywMgZhcmvGNl8P8qtoJDs
rIbHg+eUrxImxOe6btwND8hFl0wKpTgWFBdNJC4bjRDaZYxIAxDGETr6WU5Fh3RAqM5gxdLOGw5s
5wY0/qZf95MaDhPEHV60HsLLbiI6XKiGI80MA/QmSJbDzxjD54MdAbSpgG5QhtNOeI4aIJSe25WF
9cTcgLk+ecNhOi00LINZK9xMLJqMhPYREIJz0woNHx666SxNxxuuW6rI5GUNriCqBPTNKT+FVTZN
zHg9b4sSZmuJ+IaJHdy9FHJFwWuBxP9u9cvwwpjyI7Yjwo4sMZ0LzgXBq+pfbHVlkTisEJY5nhA7
Bho0x5p3PfBHI2U7KFv/OtZ93/d64iuHh8OCIk90ibnH8AmIxo4A1njZ13o3IGg4KO82AD0tUoD2
4nTkH/7zIJfwj0AFrTPy+XhzmR5hXCD3SVCkOCcfSdpptpSfVl4rF7F5efB9LuzRt7pFEIT1wxzo
4eDtmbUjK7xK+8/VLVzcl7l4Uk8LqSq/JUWKjxCxpiepWsasSPnr1XtbsrSMoTbpafrmuW56Bkm9
W1NAkOn4y9qYCOyXd7XdL4GtWZk+JzkUL1XyqGysiGEhwnt10+CMsAvgr6OIXITO5Yatko6IsVZ1
XWVhS7WdzygGFsQgjfalGxqKlUFrqlOLpSGSYpcZ8KPmmh97/IxnxuNiS2Jcrhbuzj/bFMn74ITM
a5KYZMI5yUeb1Z34vnH84wEYEqXvm8C4RS3Ciny1et7FdM0b7/bTu+N0163BI9Gxq/AeGO+lEKJv
TcEbEgEVLqFImhsbHf+KOEqg+/eok/kyqxHJ0nL5AElM4bLurLALjfySJ3fUowFnq3edgEJwdg5Z
VLg/ph4sN0rv06CEOnCU+b1wSHUuvkeOyfp8BoD5eudbqJBBV2T8eFPxZhr7bwRmlI1utZBMCQuw
bi0jE96oBxagO3v/GYpa/oXU28hEZ2DK16Dz5wN2NP4T9e850z4p5HChVk2c1n3JNBfhny//t34/
JQxMfehJ5Y2laj7QgFB9nRywIxfmhBLaHnsMajybVV7EuGDfXKASmkSPO01tDfjz5g62jN9rG0u8
fNySdht7YfotiSX2vq/jop2HjogBoIqK8+Oa+sOiwfFnQLI7Lt28gCat/O3oAhwvUwQOieUp0OWy
RRB1gWn7502FcneTZP6882l3S/ns6vlSIuAidCk+gD1vKyEhwk9HcfrV65IR79G1MPmga7X78Dho
+xBLZpysuG0V2rWrQEqWJM5ul7wqpEmGeqTJX9e3MkLZB8P/5Pgz/p/Aw9yqoJfHQ5IM7HZ6zegH
F9OIkdtAmIV+OJlYBCDy+W4qP+cvRQWGTU9/mYNA+Rio04IqX0nP+6f/LRVaGagGCPIGCHzBvDE3
fmbTaSKkqlKcVv1X8Q5JXxMY/q9Y+FDOWIPvcP8sMczlT3g0V24/J3LfJXGU68VrFhIAsBQYH9f9
3RRlcC5pJUQ9PQ9wDretYowlLZ3CZFILMavx+gE9RFCw7cp4uYm2YMmkB375+/o4QaUFlDsGfJVh
Tb/4I6AONmhvCrxc68piou9UHTKdYmPGoDwGXM2xDXVoI81KCQ8JKHcsTsqdlRVFsqaE1q8MncV7
e3S6JE6tnyOmMn0Btd7VSDYbTsghA0FWYGqai6eDMDkbgOE/Uc/8nl1fxF3aduURQRL37cqK6OrQ
JICnuluVOXwyiGKazUK/PMRSaKoLStCoAsafied7aWUT/XPdPwim9PZiY3eC2OM6yYjogpHz2mFK
o6byYKvUbJBlw8TGsQDXUeUxLlREJhyUTshWGLZlN817AUitwzetL9o3hci2p5zcczPHr21Bo472
12EK5iGr6ouSFkVxCv9ayyre8r/c3/kvnegKXdTLD3+eBAYFmM8Pg1wNm9P3IdsISOm6d1Y8k5Er
tlhTkSxDJNkw6/EqoG3FPU2MDJ6mldgWLGvLKlY61kPFe1KHlCSWgcxvNyRg6QZO7SLUMZKiZM43
kuS+5As2V0X2R5O6NzAEbsucUxEia/gce59KaQ4CG8pPleYNm8Njket/OAtR4NvjKyc/t04B2lA8
EDkCWj/Y1zdLnhDmLI4QD6DNSCnL0J4h0+gxaqpgzIxhJknOVoiS8yKhw81dUjdpKKYP2W8+ms1O
rTJ3LIf6ViBYlPG8pM7+8ZvNB2F/Na7vGHbK2/EAcEKf2xHIOqvtMSmoYzadF8b5GTgN5nXJyMvT
hsh9rPxR8Z4zy4gk5HCCD1yVncwLDaOcNbWfWfvZR1F+yhodFHDNR7Pnh2ygZCgznG+JtzQTyHck
ON0wvvu3tzKsT0bDsgE/DuRIe58hAr1IYHjFMHL07N3Nfbo9Ug6mIb0p/eWzVGC/yGGMat8HT2N1
5PKyRDQ3rB+XMOwgGQBmqq/oJ/FzxH5J9do5FwSix6oq18axnX0K6PEg9OcVtI4Ig796oDDHq6OY
g8yBdK6sNQ0Ed1PHQLnckZPJUvZqZdBdCSEzXm4A2la9NIAwh17s9q/82j4KxDiuYiOfvHWaP5F7
oFTkLL+Jtrhy3oH8nHXAe3eu2AzvFZ0JqCx49D0Hv7kOpynCLvsN1tBYFQr3KLyaSycpGiVBKXHq
MrtcO3DI0EgDBmAxTpa7/Vjsf+DwRHFumAHg6BLldrZSnPa9Et035uAlNHhujx+Vn4ScMHmwPUGC
tAwJiJWF9TUbSoVhkWGtzPJZKUqO8r2STcZoVt/m9Z+8tYG7FW2yCh0+o63Iwp6BkJrZHTBf28/n
+KWObGqEw+3fmVoxFrxnUQa+4iyLaHetyetmaZun/GlA1abtT1lFE+vgiKw2Yh6kI8eHsQvoFwDD
/GTyqnGE3FEP33cKHaxITQjQ8VVk0MDuYob/nnXoWLt1Sw0GhS/wREwgAeViejVfomzQzbHs9BPp
epJTpiqreBqj2egRHBn0mqeIeokkKxVTgUhHBrn7RabPzVqTiqjr9AtGCUyrDK86zMVLgGGmfhRJ
sD/cB/3iuI3uz4dQGgqJjwga9lJMofRYLBP5pgrqEK9lXhy+6BfdR0Quuvs/XacnTrjFK2fR6aji
ckY5aiYbl1O4IWp48X7i4l10SmXcIAr/Z3LQtaSWIxJuUKZFRF4b+kH4cPPvNlr8R0rLUs+8A28m
WLuxGGS1FJBPtv3f+bcgsOeieGK+4sNjlTD6EqWhgGTkEtQBG8qRjUzZkO9QWIrxfKxPYCrzev8K
g4SUJK3TA2Z+4v4bv8jngiB2Zp8nJ4cBcs1PQvvCtfNgaUfcT+mNs5PsmljF1mdn92LwKBbg2qFO
FEfAJeCHyc2lBUxfPTOFUGp62cUIvGN3j7iarLDuRdf8z2FQ3NeUaNujLeA2i5mbsKnH1dSoH6qT
7QAAqT9x3GifCAuApTNuIB6W3qW7CbRnlEtfPxsa2IjS8Ngl6HxJgzX1mXkZrmgECVHApBhYevyR
WTb8359X3jVuDQxECgDKP1gg8p6yn38S7afrhWRGQliXMkDziVZFCSNzB4dXZC/wMtxRklFViK+I
KiYkyJrMuWMmFWyhdX0TGPu3VyskXMsZqQt5CmdKmTFdwHEHkcro91KW1J4THxNr1+Ztky0046uK
GD6O1v5r/bIfMy6pnmhnMYBC/pYYmE9LFq6cBOY/YRl4pPOe9yin94gIEDmHGfchKTm480zA18Cz
l1DRmqvAnaU/Q6ElbRrpn8y7muHps7P6uDnECYLQ7kzWI84F+KpvF86v21D4wDfJA896mv2Hle7s
AF4G/8DeS++G3L5J7QzCSOG/oFijrbrDdwtyoUpgIghsVjzlWNsE6u9klrqPQ4S/menvDj/+9uy5
OVfTyMaZZiBOSBgKN5eVM0SdxF/0HGs/KrV3aL/VbYIT/r1J+fGNPbRuC5uGKX/htpCQK7W3Tsf1
FGFtXqv3hZ0+T3ze7BZN0rWgTfgMF+Vx24gaTntJsHWmlCxOLi2n7j+QOUps+rram0Z/1FLiYy++
+01hIdrjd9XwacaAVfk0L1u1k70lyNOxOFXf+l9CgKA02fAL2L2s4zOWUo6ggV0VBETDpSLxpIeF
CxLQINqZKsijkJL6wYbjeu9Q7GCf+HKa8PKBoERl3YiT7tYzMMSWaLNSRqleWcWhDpxk6RrfdYjq
kvwMwqwHa0jjFlTrUiuA/s3CLvdUMUCiIeQqrQpPOQ9J+dGGzQ43zM8R2d5a/OeOPZV44ICZMsRf
X1dZIZRLEnFuAnp3ud5Lvk3rg5MWb9SDuEgG0ybLXekbXQdogajkCVjNBaULu59qKKpX7v2OvE9Q
56uyiBDjV9VTFK064DzmGtoxyphjxWS96XhfAQNb9nhf0iQ1zhyyYxsDa4DbfrFqSAmYcyfkavkG
1BeUqchA0Gg80iZGPh3Vn+YES+0idULcQeTS5eugL8k4Zghmibn9ifLWqLAmAVY+TtNT0VaCdXqC
c7o4x+n4I4xMdTWu3hnCdhHp4Hx6I/SEcdKX5/jQ++BeX4zXWPtveSgL29y14M0rmSDC38gQH6yp
xqVP/xLi8ljTjaHvEIoH9zeY20hWGqSiNk/UgcGD+lFNxEwwzggvec0Oh5YSR4/MbOdOjWcUmkaH
xUOB/KxIq9orUSYrDyrtsxrfga6YH2S/a/uQsTtoPKqtN7XbszEHKyN2TKn09KOz4jjzDjEs2tEF
ILpb/JfmbVAgxobUdQy3b9M1ulbl67nyCnvnfZX/rRkCao4vFXbnQO4C5tI8IhgryHJs0YHICDRo
YT8fPttpCxxaURSIwuRPEHOf7emELgXTkV/FQqLRDJg3a/9RR02CkvNmKHCvhXdbO7bYHMwPwyli
+1xEQzLXy4iV4cWUf0etEccBD3xajJtzYotl16yRHd39EaTYKT5Du93XVbcSTc9tAWKxmr+p2zbu
SgyeH+QDZ7pJ2bIl9YKiqAhNXJsZGdVn2FGCknlM6cIJrBM9pbrlLL0jjpaTQkhdsfYsit/DD3Hy
HFm9LSGJ2aAzquFwiASCPS0aZ5UfiUyo39ZFYFqH6mblHpAlzoiG0rXLv07FgdxM8GMMBeAJ6EAx
7aGJDJwy4ww2sinwbHB84S7yyAEsIilds3cMQXCepSiixFevCj8EYkuHv81H/nTrb2u2xOh8Ol9x
u76Lo8bXcz72OvYElhzzzej/dEsJ7Ftj1dPZ85kyT2EesKcjLA3qat9C1jvBnsO28y4j1k8Yw7Di
HAD/cHPszXoTHU8wmbpP9KsckS9345ZBQBzVdPYmh7kEwvCPeqlrJZNnjKph5iLj4KeBOwAOyrJh
c8gt7BgMNoHqQtZR9Ml1h0FFEIqzD/FxKwxXEaP0qfhMeuH1PFv8o1RYPRAqncAR/hcyU87vNPM/
fj2go47w4f5S3/NkE3PeqyPULMfMS6NKwvoXGmcxV2mnFrhnCMdwvRgbKcpasUBUf8z89y+0ZgxB
1lXVW/hDEPhzNZY5IoYALU+bGej2qzjtMKYIfpjpmaHyk97m2mDm1G9t8Ci4i3Q7kUCOS6aKf70y
F4w4lVq+HIza5H8HxeyDDS8PmbAzypXU0EadO1O92a6PY5U5FzAIjJNdi05wztQKXN+N5KtV+oZa
vA7xCnPPQIUY44x+CMNbiLtjgcAfOrJ8EEHf5brBVfiGZ6bZpjAbKtTzERsOOAUEMNi5JgR4rjnm
j4N8g/9vG8tbO09UOxW1Hco4qRk36m8lXOdqyWK9m8DOmCPhFgTwFKz2/VjQWceESgz2fY0IKxyd
dz0xPxp9UCXvAh+VmK4jRihFwn8m9WuKsAYk2WMV8xs9Yty9lLlYbFtOiSkRwbRRJACX33oO3D0Y
9gwdyN1V+cJovJoqTNfBKMzlldEI6xX4KG8QUCaYLtZM2O+1PUgblx+pgUBU2XxA0Zm6A1/dxX8H
bsGU/o3OFfDuY/egp0hOxbvZnWhNDa6bNCpNP5nfncWXRnYdNQtNBkDGGPQ2W/xJ2yb2kRQuFtd2
rEe5j0MDfXi+Gg13fBvI2q0TBQOeUBG489V2D3x2kvYErM/9X9H3zwUB0K2ojz1tbG5wmGl3qMJ5
tFE8njXoQk15Tj0iZNQ473uTuJitFostg6n2ve0CFNyB/0ZvzimQbwMLHP83eYF8MIGQdPlKVx8h
/HScVTPDX7g4g22iuRVDccBO5g9OtXRBAdXbEF5AKRRTouFyDvDaEloB9wHpJ9pmT3/UUvHiFP+g
bK3djONC3NoHKAAfHFYROnlMBYNMHFM28xhJ0+jVpUWOSKxgQaUikUtcFyFSw74lL8gHSb+Y5Nuz
wJeyZsRBQjbuT+yabO5VsBIPeKOTkFnLirWgzttySMMTrstcBxOKTY4oLtOjNX7F4Lj7VI+8ZEvt
gTrsFtMhWcL9CSAq8SEgGQvJU+VTgE0kGQKluhHtQFYTekj5FEZ1HFZFAyWnS5QzL1tHGEP8yh5V
DiYyggd8U8dZhXj3NEJU72BD6ZunjjxiTT53sN03Nou7DXItzBfRdkV2krCTVtehO4hWGdr/feGl
7Xea/5Lyns9qTNTjF13mJP7s6XMWmEUsUa5pe4joW67kPZZ/W4P7sQFD5QlexjNuULc8GODdp9Hz
YAXVpaX9FgukKm/E8UFFXb8kJnMBYU6w1l6MFikgKOi+Trr6GxiaMFq+7XzA0P+x89DPcFaXB/Hf
yLoZVoYhnxEZtsq2PO/2nmIqNkTyhog48uF7BKQIflyua4IoyWaqbeY2O08wQoAE5D/OYAnNEpeD
HA0be10efF2Eu5S0c16m97dpQWYaHG/g0TGh3qFL0XMF8pz4DaW0/A73M5rRh0jqXkC0gCvzwRT+
5VGmI9JmZqn2mDecczSR8FcDN/S+Dp1p3D+/s0VzwThCkVFYXdMfelXi0QtoWL+XKdm7zSGSCx+t
Z/GKAYL87uhlNStMbXkyd/vJ3B5jiqqdunRrKQsoxlj7niFnXKAHivKCSuuWew/8Jl/MOFmCu5CN
yviopSYHufYXwgWJU3uofUgGYEGIcosAwNvIMsaisyr5w8lOepmzMM7O3gBV2dyd0GN9ns+v+mrA
Tw88nqIXx4L4JVpDo0XYZ4fbnDe70sOVzBtVst1449UXbO0OtzwdralHh989JeCzeOEqbXiareqh
Qz+84QrRfJD85lkp3VmZz8K3m7CQ6i12IStqiNJ9HzlHz5utk+2W4lpKT3WwYTfMcQdmK67iJv+W
DTZHkuSmpxc570ABiwRroU3KqzzN1rT5wWU6kD6Wc5GQA7Zhu+Oo65C9lMjiR0+rESpilleIpGHU
F2ix40NwOZ8/FNNpdM0KVfGLRw4/cDybS0jmW7EhKaI+HNj03/qApJqo5uHXKLxfv8yoYSMqMy9r
yC6xcNPaQ6krhFqDuO0bM/NizC7WO4B+Wu08PTcwrDACVz4LA4ahWNT+M1WqY/xWHX8EJPEk5Cq8
aI4VkNf0ZJg8mfPT9vtDsg5jxaaP/rheLp6MWJdDk+lxr0LVlq2J5YqsLskPc5HneDgzqsbchPlX
UQupeIGCrKI5cOnAqtn3tFRmdGQX1j5MQads4W94cUMpYElrfVzD6GT1bBA7PCMGNlOAL02MWrWh
/Tn7ViB6jbPgGGYpaKJi2PSFRYyBzt02g2wi1WLuSjT5DEeQqJepcBlOzoAhDpt53Rzga3+/eCVd
74xyY6C48x11H0N+pPn4OEFOx7Fsakk0TWFcU7I8jB+eBvWcHKSjdykEV/KG2WAB3YF4jeCiC6jG
VvQGW82kzzCC2Fk54uljhklAgfUmsyp2QjxyS83GdXJDR7I79qFTsMa4sJX+bWCwoDz2JlmYIyJF
TVXyO9jrNm95J/bS2Z/pgmidkx1QyZ3qQsHxQy6/edFZOc2YGjsH945iIBtKTgxIeSj+dW/rI2Vi
ap9gjtFmM3+vC0LrD5HCHLh6kUJzTBPnT+ofyUXlRRg8dAX4N597Cn2xsixizOjbnCyNFvagpw+G
YoxY3AiRv6aPeJkKfolNpyWaktQXqHYEehGDaPoDfJL/Gl9QQiLfkCLJ3FJGsuANaeKd81qt7jqs
+JxWps2tQdU9SbwQfMgI51GCdxADnYXn4ju+azCAacxRPI5YvM/qqkQfeBz/ce1D6svIdr7bjAa7
1MHnOaWBYhNFCSsFSX/ZhKOr2YsUa5x4m01f/tykD9vDXp3Nd1wWm5sxuMa9mTToO6pNO/4OE/sF
XPAFtHJ8S6MrwY4Jadu0QOjmPei2tOlclYO3QGTF5MPIiMuufxDuOLIAsh68nGSBETO0nRNIZB62
1zEVy5TSABfGIhFHYAwfD7kxDTkxXpqq8tpFolsDJZjcAq3FlcrhHF04+93rvY39Ws6oLF0wNN0q
MC1kFP9WENYfmb5kbVLPtl81nnogUH8d9C3aqgmneL8AXxtESISXX0KgQ4VJJKQn2IMcNED/t0jB
0KHuHlakuhZ6S0PECGQZjBcdSsnIL4nNXVKmvvOUlGMf1H2sCKuxI2hr/dOcqTrp9kTDN11CVsDM
i/w+TMIj5aZaC+WUz5XIrFyoIjojJgUtfwr3Jg7u1klFaRofO5Yd/2Fcf+00WpGRD/j/p0cfno39
5h0Sn+kd91/anNOf36rQNtQ+K4MUdomQBN33qaqdyEHL4H0tPex+meeQQ25YRF9/F6n1+Tsi26F5
Qi82h/Jf50abbEjOwOpf1OAe669bpY1tTdwFRJZHbgjnTNLP4FKOqc62H4xQrTPlLRKYkPtDk+LB
7Ew7Fxk1lAgZ7fadMxnWAEnJ+XRlKs11DyJrEsEYb8vDtWcbLBS6t2FCIFT+X0iWqqCcNViQJGjQ
oVC8QKHCkgH7NaGXxAgiiOhLKoW2FfPJsMA24owWOG6BuSEGP/E+PPbj1sswVRzuYzlxShUMivqM
Ab6aTHcNj28cXXCLsTLjurAxqOb4lWnLI7GEZ6jOxLvQeV4g/7AM4KuTEtNJML3Jm4vmZegfSmPH
JAFlX0qgsv68pTKl+8fDne4EA56dLeoPcejnl18+tiZm7KhFYXvd9Lfhqol8jHJmjaKvJIN8XKSo
BC4+Dik+OgehBhxpQ9V7s8vvJuHFcjE0xlmLKGkD52l9qhMYk4X0G/wb9TzLPvK+khBhIC8dnxi/
aWtU6t/I1u8dm5G6WAT2S27m5yvnkjVq5F2URUptiNvyqZGZOkZZcIaAUh0rK2TAFp6UrLdi9ZXn
FDh5pxbPIolHHtLzPA+DO+Bq3Wv/YWGQCg9GidMkU+I67FIKwXAoZPTiR60mqlScL/X+70TOqLlC
7HmN/xe5MkD3vKFEePWBIIZDc4gyyvkFryyzPsLEHOQMjDHSgc36/N2dAyIK4cBDDO2/HBVkbDkj
OR6ccU80YKjUPw2LxaQ0iQP95uEpp4KvaSuk9GK0/C6H7c2m5IblFWAewtL2AeY5sNZBxIoL5b8J
O5+aECn6dU0y1K5NdkJQf65FO/rOqNjcJfH3DvZGroeBiakqNQD7lqEp/q9P0kXDufinADPnC+dP
ogMIrNC2LtnCfERDGjPaBREjW7o4SYDgD0wutH+NzMPhdmjVscO1R3gQH916kgbl8yeG+lrxczqK
UtvHeYbEIpm8TTTiajNf+Hyouv4kkBbZYiW9e9YO5oK/bLs9UlHo6kQP9oBeH7J6VZ8MhPl0qVGQ
1DaJUs+EkiirHjLv/bBEZTpjKokKfaxoeMG1WBAjPpWIyrD9gmAT0E96LlcRByoNzIZKtt7yU2Q4
9tD//MCLqBaXbR4gjE+VaOiQQRryGe/V3cGiI2KQ1xiBQgMWw5ZRi2NUilKBYqglSZrc3mTE6Ucz
ybNa1t6j2iBLujno2GlW4W/ndLMj8nGU1al8JyOmWcUdSNfobsaGOLWvG6hScNVCxbAocJuMwb86
zHTqm58QXD0O+jdUFtLzQloB9yYJWXJ10DF42d2BHfxYYHzmGYRbxJTKXWW+128BY6pNdHJpiGd3
AKeHDIJ2BCXTCJD2S8XUSsW+8Gq3a2IHUelhNFcsZ/OTBGMQn2rLjlq2KM+Rhq0NpJFg9bbopsr4
1GYNlgiIo0njl2txjhoBnGBDKc9Y5mvK5OwkURDKdP2mxL2ot5tpyMqq26TD78f5t9Gw4y5H/zdx
7ARXf2hCQ7SaM4Jw0kIcOJxLUr2PwsdiL8ivB2QGy2aIsv5ZQVmDd4ogWqFK1U/WgrOdVlmgGysX
0iz78F7HnXGYffqvV26/vyBbnWXTnJGJXDS9+MQncnGjcu5lZNq0F/sRa4FRIdR/SSHnq9K3o8Ab
SqkWrbmJY0wfJXAPhW6K53tIZ6J34tUU69xg+6gX2RfP78ISN9qFFSnQ2vqPsEMU4zXlvUxvDAN7
BoN1XuC45nP8TMyI1P86iZbJL84a40bOVzzqcOL1V+RNvUeUwiBUricL2HpoiTRz4VnTmq0Y6YHL
adL2lmOX7ILy0Tp/O6oaEdA1AmkC3T0UyKH+qU6HS7/Dljz8dS86tvlEeiyPi1D6kVD46PSZ1sUk
A/VsfRSOfJdYL/6z8ZmxeEpP0cQtb8yJ6rSGjthtS3AoXyroTZ7dzgYdMjMLmavmhiU9z7jD5Qur
DjXH9g+FvGWYDk4Qj5w9JZs+ATlrSakx2rMudnu96kD18MPSs0y8wVAik4WWjeutC0obX8FilUU9
27jWUhWmrKdHb7meVu1L3RA4PSb1qnK7TVTbnj2aZ0yMLOeAB8ggZKvWn4ixzJyGbhHRpKpiXH1H
9PeJ9hluTZoQ+VBvRPZoTmHa9sw/1SwPW5YKknmPEqvMHwOfu421WLTvjtddwSN9p+Tv99RmO5IX
t5+yP4td9LhLl5JBsN9cpULOMMb0d+/EIu7AF0S7LWJc0nx40ttP0By4DH0iT/QS11e2UzycMdcY
Fvd8n7qeuOSdZral+N9z8Q4B0ru33sXhgAbL4onvlFJo/ukT5kHGyi/P5mugKBNQecs2J90a7wh4
Xlgy9/Dj1SY8l5dBh4JCsCXKINXycwcINlkRNeyL6yMYOgSfri3825DwdlR+3qWsdWCdlBlo3L2j
RPE3xD5/TiW4jwFURcgQMynOrhEQXFCrguxwlcAjP2ZU7Uoo4sIBK9pGpOkxy7eoKkusC0agr0Yy
JFzLwlrPo8N1c9bkuSE4k2HzMJJ191YnONFV5GqSDi7l3bTZ3vcclh+6HOPpT9h3XqZnYJHjzuyd
XhOqnBXulQHdXZ25A2rYtPx9QEN8SGq48XrBqkQxXamAVk5Qqh4A+z+0xUEZoida0ybKerrXE3yL
lucun8OoFVCGuwdNy9I/uOpubc2tAJonQ45Sualr4UEQnumLACxSxB8IwxHy9W7+1n9cENACIJDF
jfhCPicnqd5hQREJNLFx+gT22m9xQpgbTOEAHBa10BRGwvgZCVHQHD7T09hHW5DjlvXEzhgZr87l
+sKhi+YybpP43Z+nghC9TkR6CMNPt9SyegqAk8iMelt0AjmICxqqhIKQ9l7teIT6UphlszC8CxHn
ToslTCHuM6cNrttBUWEspKiXUq7sChx9jCvLcY9e2463i7nyKC/2p9sMMT1neqW2Vzdc6v8s2NSj
5PNiPsd4UIVdTz7F9oUUqy2vo5VeiAalOeUv+25MTEfQQWh/kflyMizKlLjbQIEiqGMEuuEIVQEk
2uVkRSLmI8yZIVtYoVDI4TGsb4cZW80tZ/69gvCvDkcs8WX3eWuPZk/+h8DIB8FKharxxDCaxZHq
GEFE8o61iL5tPsJ6WVq32AC0OcaWNh6SwgFH1hkI2QTsp9VT0VyK1MEa9v13gKhG61LVF7U3v/n1
uy0P+tYzxPgBF80UULUeNM4yllYUm9+mIvmknb8TTB7fTbFI+UrebLF0UvbzZ79zFfBA6+Rr7dwv
NcYp0fDoDzfVIdRnd7Gdki7Nx9pR6qCtY5fx19PVZ83mnS+Btb/P5uiHWI4Hyl99yEuUGoRvJ603
MqGGoI4EL8CtEcfwGP9NXIQTQhzar+7uziFqXov/UkfHCdCDHrE2hwJayWKAz0tkRweDVA7bxjj1
Sg/S2mz67v3xNjdsUi6EOsXT91dRMfIul2vJBTDSXjAyP7Cnx/Px5K+qnbrq5rGXrV/99WEAEL5S
i1BGQp4OGiW75CCfGc23RBJsMqiIOtNqdiLonG4zOMf2OqF/uY6LEHVuRgqtv2sMj7rBM4J3zRuW
bZXzjvfuRsnViqh0ztXRNbmaZ/p0kC1EItqzNJ9lRNpxr0VU4q1+1/JTEunVZYzaPEEBr7Q1GdTn
2XbRwtWgUQAwtZEA2eQE+ZV6SvsDNHyQqCPlhNEMekB+7+F/AL4uV1kTSdv0XUwD+ZXJx0M9TkWl
XdMzaHqMdWTgE9+M8G74UEfS5rBHsKIQQjbBOgcEV6BFiVSCW4ElD0DzOnLDrmZyl8A+QsS1j6hV
NAN71a1qZmSx4SpjFfV8dHNBob/+CjSW0uaxE0O2WbU/xpUpox5YEiUfX219C+5NNxOhZad7Y4Xx
DHId4u1zQxrTWMkGC89Ngty3z0gb7lMSSYNtglyBv94Rs28TIo3OxZ84qDDEqMw6xZ5DQ6GIgD+V
QxbolesGCzQggeRz/eAGm89i0q1i0wdP3srwNDWYappRznqurMUaXNeqDsiVlGRqm9lyVIT+V5BQ
4gvHM5Ie1W3VFsqrQUDaLgzRdiqr6LoxphdmLuKW5TWRXLjTWaOLdAqvmjMhkWhzIId5Z0dUU1ec
6TlnzYXeu+8oV5tMQZSpSH8o9YA0t5ZEyixJpyqFqbujvAYSv45Rtlit5dbivgEjQwM3SLCXuXyN
vxjwtubuw+pyl1jQ0/i3O56L0LO8/KmWJRZ98aPc5jXaOrYNCMECaOxS6mMpai/igIc3VfaeHiF9
CRCy2wQ4UaFEHlM/xVrNAq6DnwFQy0XB5wuQnpF4vI42WBo6b8MRuV5EraF16C8e1EQ+JL7oDJBG
P6AhgF99+U5dxAMDexBkyef9ZYy5YJ2WseVBEVH+Roj1IxoFz8lDpAs+je0GCCL+9LFaILcMDjXm
kfertIPiYvfozSznBzWbptrGWfNxHb8SKvf8OQ5yjDGSijUOxBTxdjwQ216A/iaG1GSr0pmVUziK
q2qP5c60AvrvnQ520wksDuFJmsSxzwL2bDQBwvoorJNBesZ+yKF5c57SdUdikOy0pwZ/usTXLp2U
AoUiWTfwBiIdi1FG3TzQ6NWL7fnBxy6zPtCl2RVSWdghnmPOhjvOwQX11fg5720RPEgRxNLoz0y7
10zvnpkK+FZSDxkQrS2j61k3CGhrhJysiYKq8hzpc9nOWibhaYwtiGaSXpMMz482inUSkvXoQR8B
nLelvVTK8qpmJjnwkXS6suPx2FrhPtkcPpcRWRyioE8UotAcy+mwRL0JoGebuMNOup8Dbm6s56iI
FxmeErhf3YftWyeP7di8PXn0h3lEpO/uglmgW9zWUV2S+sB31ZlpfyciiGJDBDbXaIrrhBMRDoF8
HCa/nUlnpYX3HKLeLg3b0UvhRPbcL8FwvH22WWfVFdih50Z19X1M8fNprAzUaQKxnWKkgZ1ItmuR
OlIrDgK24NAvxp79T3sz3sQbUKMU72fslR0QEdPYK1KogXKIEFTwErINt558vp+0gIAgV1bk9rR6
W6SyvkgVHvhJ3ra5rGQHv3rvx1SfjpijX9VcoHIsNYZ+kIxekDKmm5cf84bUPbdV7kYjv3RSJxuV
0QSBrVpUM2oTcMGz52pmw1mttLzSjzuGvlIfKJcHrkY1mJ3LG1ig68m7pSPk03UHMh8ANIzhdX7J
/qW5mC08FmfUc1CQqGHMxSO02CgH+Nmb7fXcyGxSJCRvWb9w1kf2Ll4wcQI4BAJRNRZObURjb2r9
t/aRPRx4UtFjNwhhl5uUt1I6UBY0/rVqmCEXI04Pm4KtiQZ3HDGMXqOAls9uLhMLbQq6GdmrcwDn
8IsELPgpCBrnsP2r5fGPGF1kAvkxKmbEi4vHrklkboSuOqfhSAujRzRIO0wvh8iKTGCpyIgKTdAA
Ul46qob6NzLBo6M0abNn8JOLlE93AUkVmEJYGvlvX8FGxx8qvs/QGbk1t5PWUbEKQEXX1RLtZkm6
Az7CLoYwUAJrc5hXQ2/SkAPcXeflBkDkVvvyb0zHXGZRw7LILkJiW6N8e8OccfRLx4svKWxRDa+G
1GRtOPEtJqgLSBPkBL1sOZly23+/puAE8Q7Sn5Nj9X2u7Nb8si0DjOzAZrs7heT2V0WmGFa2gCyN
4UqqURomRS5QuowvNzIQ4hPx//qzSsbQ4lAHCEJ1t80wxmJKrKppnO13tLXQyuVU6TokHkVQsL9F
/V+vjG7F0stIO9JytEY1V4/uzcMxSZ1b7rs34cJj9Pla3clQcSjzPLWQFLoRXHReYFAK6J/b7Sg4
vSl6ncYjsU4qtbgH2k0oe1SaLyx0pS48mizbO4rynp72N4ndQM9TwWYJPHF8hmeGLYBHYsVXgHGj
j2ufkqIrRdyFrBjAVCsqg9SIcKXUvXk+Af4V1MblrWpctJhVDNUBZpFKHd2YSuB9dCbFR2W4Ob6m
Q7e/b3a6/9oi3QUsef2z3B3yzxcy2kW/P+si8rEfuQC/A0qNOw+AkwnbInIaa3M+C5qJ5seSGTIP
fvSllIGe8dXwXRuN8392dJekEs3wDu4hxcbQnneAoM4cN5QNNKpl6ZGpLI5lGz+Ppow4+Gf4wLbZ
xpaPnmCYcQ8iAus7CB56kV9If5WX0NdMYZo5bRVCO88F20zXx4uLR2WBkpFuks1sP5EI2NJIeQwW
redpITykmNZjcuf2t5BueIDAEezVuzsDiTygpIrWwW8U/mL28xISlRPuY4iwaa5aGTTdsc5opiF+
8w6p2XH8xdZicSA48gxAYZ0EKtsbo/NKrC/RD8RNeVPNTZ2wyQZGF558rRI/iFBCZK82cF/8QMyC
q2Lux2BuaHLy/ducsNPVvFIHaIX7fqmREQ5QnWgMmoo4YdQzr9PCJHkVDGtCPdWlGjNRntGL7oXB
YXF4lxqWAeIj6QzrVFbmwi8wDKNJTGkrSyenu+SWvYl7exkMrHBj57VQod19isHi0v+UP2y2iplh
xE+FEnhjtKOPrB4E1Re/k6eKONR9yOGMWuH99EjrKFHw4961gN4BK5eJSwWKRthSqG5JcfqOYsCO
x6EtHwrQurmZVIg8rPxnRRz4yIEX9pgB5iIKpq0ovmr2eBVeU14njFdrNAx9WY+8QZpvwfFSdV8L
++6BWTnflsk1IYdd2DfsedPQId/lSuR4Gj+0yaUYgxiaBIjnUJ4Rby41oNInLiEDm2EDDq6R0/we
bLW/3bVs5Vtaq7bg5C1HuiGDCFmSEujoInXZOnvVLzPUeN8bPizwLXX4SWvfH1yHFD1ClVp5szCk
Y+1ZbqZUXQXfOXV5AwQ51g7N1bP1In95kPLb6B+xCkIigcFHda1G7WjBFxZimgHPq+fdGRvES3uG
pbXgUv60WhDv1g/lO2YoNFv39DzvZGFrluSjtWJFnwNRp+zt6ptBEQucysntfgIm1vS9eo/OKFEN
4vQel1U8p8lkiJc2845xQW1LQ1wZb8nQixJfiWJUu3NkHhVklNZ4LUNzEe8u5QrRexnU8fhA4m3M
NzXDj4K/R93Vap6oXFiLTcJvsGf0zjzmOznmybBxBtqVRcp/fs5CmqFJkx/BNmp4pIzzNFDU272C
8NHwzDIoH8ohPSgCn7PEH3l05kUGu4LgDW5hQxhyxEKyOnt2JzZ6uh4HHZ3BwRFDnTJjedlA6N3t
fb8z7viTjtZSNVM8gH+vS9rcC9cvkCEYyQH8vL5U6a4ZTB/ZD4ONyGrbcHsVnPAp3PdQGIcXPH2P
ReBdsdH1vJ9L/ADY5Cm36Wk6We5koAAJAW0RX9vFAuacjgw6jU4jdQql4DHL3ZmfolxcGHsoVfX/
GbdbfTqv/it1p0GPECYbW5NOGQlywHusE193YgHOe8LsJQPKMwgCe/w0aIdo0pPLJjcFaVQN7s08
89WkAQWm3DGA7YLLzK8Fw6Erfht3bpnstubUcPJk8bobHw69570KghI6mcIKZkEOhq7fDOSKjXvX
wEq1YrvS2VweO+l4IYmlwkl8nQJ6PpkSxwcJpXGG1LpZsJlcRB6pG+aZc6WSjm7U6b1sNJzEimo5
WAqRkIBMzHRajN0dnv0s0ITj5AsBazlvTjNJIAfRE7LHAL6zLVb8YvuE9wMltfSU1YvGLmT2hn/S
QAS0PVhqzQWlyrCn1T9U9PU4QuPR1N5BURDkP8ddh2rUIgX/MdxtfkCepsvIRD8bTrKN3kbJ5kj2
hFzmy6rEUJBdEui+JAY76dA5i4gWbhG1cs7GGDJNAp4bRHjUFxhIBobhUK01wqdPtwyV1+MEZSnj
odY/Fl9xyheGsFM4/EbZsIzruBlYFbqxNAzcfoxpzKDpNCWR0NlETM3v+3bt14kr8gGbUvwqriEa
cr8bNSdnJk0tW0ljmNMU9fjSqDieYFN9DhwReJorDCFf45lMacAJHp39s/WeBbDbw1bvsC4QIBE7
2lYLiqQ89DghiEi8V7umoHV9z+aM0pxKNkQhVX4YDqUrkFXBN5WBXqsx34jBLfWB9EdirAjUx80y
DAVo1052wQnQQ8SgI71WwgkgREIr0Cvc+jxmf/cv3Yyh0qJup+9TTkRXnH73vlWSRhJCYKJt4ZIw
q33cjTzm3vT3CTWrWzvKIspWoFGKFJM2fscGARwGpUOO1bCxW0ZAb/rE4DPIIQE3U67WZ+ZB+tHR
BkjOTXmtqioDAFah/9XdDb9bqMy9DTTR5Cva3cxFhREfhn7Kl7+tBgCy/qbJ0EQWfDjQgJu8UG11
2UaJwCLawEOpKhwcQxT037vpl5O7wC5621e7raXIidcga9I7dHU9VO1Wlpsr6P1nshS0hG4TF/Fs
OXNSQKXg0KpfesldCI+QTm+eKWL0cRWmPrLhFggGrYzoY4csBnTWSUn5mZrWkRQoBBxJvqgUgohD
NoJLQEdHhdENlSSgtr1E3bc3c4QdLdxwBMQ7ISENM+td6Q+75W4lBDYwszBpZOIm1UaImq0Emiza
D7BwitOlYC/FgMv0Ln8ggEV2aqpB56RIqa3GErNtWDFg1ZNWBYr1jP6SfqS01fKi2OdWzh7LDPWj
zD5SEE+81b1LLrgoBoLkY03ABHTFjtZRNHV2Tu8YxjhCavlPNdJeVjkbLpaL3h8Tdoudwwdq4RDb
rZiGrJTN44y5bj+rs3eoQT2Jwix7gzdXZKXy28pK/xK2AwgdPuDF7H0CYmtZted00BENFrchimcH
J0aNiTIOFLyDiS1VY2fMvFx/euqRpqwIxfo4vUizX891h4Znu4i+PKYaqcU+DTvJkS9JynuIYSND
kkCLDjr2lf/OAVxemO/Pgy4y+eTkMczVeSZ9nJ3n98Vrq30qKZbbt1k58aIHMlmpgjuJ8kC7FFny
tH21mC8xgohDgx9pEtztAlQdDQsFlrCrKAH+NTZyhGxmBrO7Eveqicpf674UPCadBH50sEq3Xx9F
AIMx+63hbKc72pqrQLPRmfuAcM1W6GKywmtLJcIMkGUQYwjBdlLwUO6qdx65izn7JUWF/iR3Z4KA
RXCKxkUaOQ6OFLAK1aWOI2pbjHzoD90quxHsgZxPs9nxk3/rHwwJfmwz03Ci7fXqTzRlHd/4Z+8j
1/Jn9g7yBPnmS8QFSCJ6z5Qe2ZXcUcpivL/uq2i8Dgy/1UsR97TIZ0+nrdxDi7/IhcmDPWJk/l3+
hR7Ai0XYRUFev/dCuEU3HJjdyRwO6z6v1NevvlZJc9bw5fYdz+hl4pAKDSPcH4juxP/jrnFxHLYl
O9smqysoI/ZI0MqhRoAwe+lWctHoe5ZnAmkfqZ1it76w4bNa+w0hITpXYTDbPMHVFyZlBszJI1GZ
qmw7cVyiDGME53aPOKxj4PXB6iuT8+OcvQpSDwRvZRWbSygHgL7y440BAD2GcW9Uh5h4weB3pAK3
O9k4YhndTKxBNMhG271t1Ew3G5ynP2YChGDTjrXoECYsEZhLevPPlq8K9GVT2+aKXvbieuYKEiZi
N/VSVbeaP2uRVjoGJvNPwljCzlyoBtTSZ7BDBoJvDYyw56qR2uPayJtCeCUoCNwgQtuLNYUh2dmP
DBgq6i1Wk4I5Qev14tXLOIEr+1qqRpBO3SkaVcjsC0q9UGWEs+is9po+CpPPQpkfrc01kG3+kAdG
2vCBFMhK0hGDj74ir5m05eDDebZPPOG95OvGRNEleUbJJMJztciM6mThMvGfBcf7FTdY2SPaYi8g
9/9BO6spH2JgzjMgZSkx1FK/OowFG0ThU/oGDQL/pZfdzBL5IJJoCueAwJqzz34zhDUYFbBlzPRr
SOlle0Vwj8WspswfB+KMlpQSyorv3K8R49Vz6DnZllN92mqbNWhRD9EhPZYx+GfukQ7fzTZy0C1n
mBpyCJus3fFk0yOppzCfgDUq7rMW5PMomCE+LxiO5kDmoVC1gkuUTow0gLgb5bYRunqhqFC8qbn9
yD0j+VZJJXXgwe3pSxGEsg7LMadxwazPVp/h0AhoyM4d+BVuXVTHdrW8B/XsZZpIz9R8dTiCANys
ZnozGyZjqv6vGYHGWduYzilj4SYvMsUEnLecmHYwTYTA/bwUhc/OFD/RTeX/x+N1FeTTgmOmvuGQ
KYvl/2d57CbQ/r+PX3J9dcogOqP2BsuXM0X/yIYdAm0ue4grH4Dfhr0ayKLAabEg9PyldlY7RDYO
1tM/9qxTeE4AwRODnSpFUG2U/x2l42/BZN4Cg6675GIno109NzvVurPfWhabppkSG4A+aAUnREEd
mW++CXYaiLu9NUIZfdUYMcO9gISG0HNoLcUdB863qymlfwdc8qJUjKjXFoLvFjhYxqITXqtXSryp
ZmersH1iLxi5b/5CPLJFaRGqZPw/86tGxsvGS57qNGh9s8t8LYXhW8Et7Km57ZJxJsdPLV1TJn8C
liDpIgmn8YM+81DqoTxEDekcUnlhhW0AkqOhAHBW/imt8MiubF9ebogOqY87Vzje4i/J6g5w7Wkn
4m6M6doBbpHGYo4nTqaEVwP98daB7qMPVUvZvdnF9j7lN/LpLEPvOWjt4YmGkrcdszbeGQ6Ky0vw
Teqd+UKC66xqILxhqzgo9ZZO9P78MIKP00/X5nN6P8kyS8h6M1ZSFJi85VYtpxFy1A+yG4i1dMCS
CcfXE6OcKBnJxnCuT8PrlfbLu8qNO/Lzsw1IbVsHRl/zesmAnpkGJPusGJ/LB3Tk3rFfb/sh2SaA
S9OB1v/46QaQU4K2BiL/rT+D7V1BXOqmExWXOn5drDumwSATihHJLV9rl11X/fjXFqOa+qINJ/HP
PQ4Xfzs7K0ms6e9BEAYzbutMbTflrLQUxGH5uadgIgH4yJml4n+SQEC1k4uMMBXq5S7i5/kpcO+/
2Pt7yHlxlgPdRnGh/aKWDiDyb3DxiBilPfgEPtCvtcTxqgkQ+j+QkMQuuqLLlIB0+aCZIUcwrsji
PBiu43t/mkWN/Ykb6KuPdXKBsofRDR9MhrtkRxo8kJ1IF9NETFXBt9ywKR4yWw7/nBL6BXlqmLrU
Z6MN4CfpGtirlogPr1OsXWgGY9Ob7gFXKT4X3Fnjhx+EiEhUhtTk+Qfe+Snpgv3ovlSOmzZfeJz1
hsAyYXdBgjLeLXTo7Beb3ZezE7yADOEalP4gdTj6UzClWBWDA62uxW9dyxa0Ep8h8KhgaD/yFE1c
c376ynAH3aSeRIM/y6+DQYnC62nwuii/tSxe/rnX+Pqv3wo3TIpdO1kDA5VZTjldCHjMH4rkZsGh
a8/AS9l0MjXLVCcAFtWNi4tHMRBjhc6SJwl/QCEB2kh9fLr/jK5OKGndOrqXKsQvC+bhfprz8JJX
savTIwFfq86s35rnkpVh8VvPD9CY42JmUZXt98OCuKXks0opaK1z13t/cZIE3DP2HXXxyIvFjuj3
tiV09mIHTjNG8jGwWVd9aE37l0GvTDLsr4gDja4UASPsXzK8rCBkuHeRou7XMCKYD+5F9dP9oyAh
fB/2MtT39YF7Bnq8XSdsXuE/rxr4BcLUDkEtgq7bHDFeY2B88gs5HEmkgDBfqQZdk2TDDI2DZQUH
j5KKGXRdpNemhyFYO9kgy+iivYxR97rb/TqPllVF6hBlpbDGc02b5s6WxPkxBPBK8zGsr6stn2Qp
A2K4GD/epJVKuHcPHvjLxK7xzsZH1BKNCUXPsc5UmxJyXmCVoHqRmPU3KzTiqovel3IjVW6b1azY
TJBSjeJxW5hRFQze5iLJwZyOGe/okY9vw14dHxo5asWt8kKnWphAdliGVHeqef/6T7Xwo+h4iTyw
XgA05WxvfhcwRCWkjDhUmxYdmR1zNDSEopOzPueabrZxOfrGczWg5Ci4v3HjnBBUhUg3V2obCVef
firqKW3mHbKNnr0DnuqxuVmXXtD1TJ45qAVeDhTN1HndPWBAtzCxmC+5qd1e/SYIyrWkC3z7NwPt
gu6xmLEY1JCBJm/s8de3GLVRDXfijIsh/+OMWEqxLwsq6CJ220UGhmBC0VQuNQS0tDlLkUREECyM
yjcH3zgI/4HWfIYY9tsOY/rfKcxmArAqnMmecQv9D89TMn4Ap2rmxaOd8CPmG9Wj6W0bVrXk8ptj
wnrJe+BsSEv/+bNYPzky3grPKpWa1bJa89c9dxRp1cz3ORN1G25/L3rE9QhrB+ugdQvCl9shmKJy
XG9S4IRKy3dRFsisZ9lL8ndY5pYVh4G47HgO+zROBsPc9zctQkXI4b+rNDIZ/mlBLEiMR6CSU2+C
qvnijozMx4FMNJbfn4xOWFwZXQQ+oCWYlziXpC196GX98V9GWi5xYfV5C/f3SyC9IvfTyaKC63xa
3bcSIblp+KxZJwH01VZ1A0ywIuPaSeyUyiY7axRrEm0h7eIF/tB7Ps8TbG0V6NDXdOPT+mgtU3m7
EifhZZnOADzffo16ERtAQhLAWyDLFIsFduEW4yQ3v+H/ZMb0+j0vxQzA0TC8qL/6UpQLCU6tL4sL
RAyOxjzWom8o+vlo1Giw5CS2JlVzXdshklhEzufAkwz6kGU6AWP4RoEDvm0u+vwh3V+WJ3oIo9mb
i3u6+vde8VNU7lDl3L9gYfS6P6WCFDOHn4OUt6olOZWBUKJJU0hTOaxNUB2RbS9KmJnrs8h5qoOr
fRMxi0zgYc8hJ2AeSpdU/pTQmwEpS3Ylt7g7u1m0FkZ47TwPAAkRb2ZSnZuOgMpdyf0qlc8IiJ5U
0PfIHN9LZWfA/0pFxvhsWuVtd872CMlFc35AQ34rGG1l/n2fg39goT4xkcB0cUeXzirGD7ZYVLRG
ZVQiJstkaLu7E8+Hr5e8Esw61rKP9nccGo8Ud3VZULrlS9tvNEsFZvVTW8p9X+5nO17kr8cIiZF+
/8/OvrOHcgq3OXk33ulJLS2iXVBk5+7fK680ZXmuaGf3P42B6XcNAjpt/+BKpjal6G6BwBdx8uIA
k6H+Tj503pKW/EbQLuQREU2V3+z05EzxS9bHzUc/LJLJMIMnR3N/kXTfmGU77B2OOYWLG0FFE2jO
roE/JPVhKfP0iJ0W9rC3L5dToT+Do6cDgd/isKnmuIC7dfLK63liECJNDt9/158oNJeEhqrmmFxQ
YEstO+odLMe/fN2bx3INx+ojmDUd7HuLtcNDRANzAWg4P7ZjDfVbuo4lm06ExWsv2NomyzOs2dqx
KnkkyAuEwG2/LR8WQN9YZejopze9l7uWI0oc7Ld50kssnAhzw5jk+FIc62C6SHT70S+DWtkucPkO
n+BjSjHj2RbJUsCG9xIxk3UoCg3XnpbNsuDGhCBTQkZ6VsiZFiX+qdWCLoIQTW2AwlTC9+nkmDpW
fqIAjdOxRjGkUqyGH3/59RZaJAeKpsjOh/9SnL213Jg0mNesUczShSbDDBHhhHVhSZ4cYOH5jSEl
XxPmDsxjWNUCpka23bvVjPLtClblow0DVYL6vkCRyPGo+Vflzu7AbuvD9uYq9apmXypwDK6ik/zH
VuIscC1OAysYBOT87MSXEivP9RsCM4UjxjIMbOa1a4OP1DDSupOBGtRjj1URYwAkss+SidjS38Q7
uqoOaGxMMA0/b8JS7uMp18R5d5kIvcSXuB7tDhi2u7imcjKNjSWrGAPErqtprSKKhd25wINRJumc
Y2QKATJXx2x6HOwXFjluut/Kaizfut848kHl6spSVVzBEpn04LEg06Ez+XH1Za96iEEqZC1HI8L+
/KXGLPYsuw70iMkVkfZZvWkr9h4CKk6UgLfZmwTwX7vRE7nEkti/7F8ZJq1YvgCS/nwfT3cfCKOm
ofMEoxGw1BbkRl/s18WsZWmqFk8oUrq3THvDvEwhFy2AiqEClxju4HaK52j4PyqZs1tSxeegfVS6
dHS6WiYdL2QnOCVyOR8N7IQxnRoEdxlqyZSPzsnFvi5jxtUREoo+4Bv18xG0iSbHpRxlIoz4x7Fw
0GrBY7qe7xv8sF/esRX0R6CbxAtn3lOowUUmXbnpRvw6iaCeoRZVJMsVYFBdVO7wVTLIU7bUmAL9
alsRNQ+Tcgh3mKsWHudRg35oUXKSwmeGqsDBy94WjBgFn1qL43tB2ksFPZQt1+TmMj2oDtTGVgsI
ATpqbIYnymlnO8l/u+qNbbZBnvC+4rTFC1hPVeueGuVZepXbZcr17kcyFTCYKrAwm6JObfMDRTt8
QdPtTKjs+y8Lu98dmX1JOcl7P/wVUV4HgtBDxPyD1aRpEysimGnErdKJEym83S1AnRLTtAzC0wsc
tFcIKNGMDASe/XW8UXOCJLdQNFWBgWCmQk0pcWg4kaz79TM1vRP8K8qXhIgwFzSkfi81F8c8faYS
/bWsbPYU+6PKtoQvvXJTtK0aBDpkPclXdKLLhlcuXwvwR8t1pbfgE+LG5Hx0G/AMlz3ZkPMQUIUk
iGHTQ9dXYoZh3v4UoZgeyQNdK6lcGmhSOybuRR1wNnZNGULEWnyQy81rQzXVJnfzsxPxH9nap8vk
E5yayiGxKG7kedtyIY4cGhmXcNSPIJFJ1+LGxtk57dbeaR5lCBUVIvHdth0uEReYJYIYQAyq1xL3
r9qdZ1sRBWe01TltVKP78bSFPOZ1huPDvFLyp/FRkZonGKBwl2vCcsjMCavbJJubGm8j/VHCReYE
j7FU6ExkFwDzQdIY82UbY3OW5C4YD5cPrmI15Df5MtUh4iTAfT7BHQfFPJHYHpk8dySAFhaVCaG8
yHnvHm7kDEvdsLpYrm03+C4JwFwPrtX4eYMg3nL70g2VaB0iaT46ByGg2jYmVXD2J4J2AJ+PYyvE
6wzPCjhPvpgYh403RxkZLHf8fAwDFI8FzeFlJDqLMCLswaxXGNiLP+6ldyEkBKnSYLyzCf/zKbfF
SPYiHxmlAOI2rFNcBy/d21lPyyc8rGsZmnXN+S51bsxXQ2dLX929omBkiGAqV0AW641VGUTNKaXK
nnPDMzKM+7oBqc1J9XuO+6MB3up+FAdoDk2DeP0s9zvHJ4gKfn8LBtpXxLlpcj8ahLYAtwqzNWoo
EnXAl/an0QyC20yBm8gNSf/Xs4Q8iCfWIOWhcYDWrUFTa3NVu0yAV+mXRA6JDUd/OE2lqwxnP22f
G6DC0t6Be3G9DbldXSfynehssvG5mCvTWoGjC4UAIsKuDi0KW5P87/WmZ1FzDylqC9yEJrJZs7BE
lxuqIbY25lrs7Wsicv1ldznhF6n3PV8BbMUvuoksI+ZIgdvMHjXaF+cz6juKSypY8uJfHGgJmmr1
yAoM0fyCilF5SLZZAg4r5U4WnSZ/OaDZo4HC15GgxdkBi5vvBVpdXqtc9bir9BPptP66RQvIlPOZ
qxpb28vxfWeWH4ukHsqRIFleHwfloaToXtVoXFpsfdum0l6MxaR/MkPcqFRLCvkDslIha+vpbY3+
KqHmwkPPE7y/vN990CC2w6BAinYwVHgkOkuFN8jE5uVVjn9kK2+dgoatL4ACPc1b2/hNrzlSnN6K
7VR3eDmEJuYgiuqDexH7RkFwVGCBGefXO8zKxEJe1c2Gb+rjSxrJLmY1A+fSvAtkJxShHRRPyP+X
TpmCjmcTNkF5qgQRLZpmBXap0RD7Hvnf4aAzGRP6mMWCWFkXpuFhT/5ogBUf4r2A4Qr32+x9QlAD
jYNHl919q2D5SmG0JCWnpRhLayBuKQdftj+s98ebN8qnkAB6MV3ts2I94TJ/OeZ5MvWxV9ipMS0G
QZW5IPJYlSsT3wwPoGpxyaTSXeq9Mq0EV+hbPPoDlKfJzSzmDubR1Mb3v0xLLG2vvXnpC4xfgP1T
QHmjRXLAf+fGk9A1WVoe0B5KrCXzaM8klQgs6+qME4ALIa+z/L/SwVGFcorr942E8JEffkD7AuxM
F86Ygip8A2Vm1shlGI0L4euFZVxSktPDZfbzH9wNUD5CouKT89w3gLRMaYlthAzQ/JGgbAVBkPFs
pzpi4q1wfkOkG3Fom/TMRMrBLlQ6+FbB7QcQxLBPTtNi5oOF/D1fswm8nX6uyzANyqE3arWMZ185
0sdqE71eJop78InH7g9dbMuEb7wmdG/Jrbq965WFjVFrKaTJFxmBpr5uiqMVkIdot/50cysyiYuH
/ltlqBAnwUdpmTsfFf0LMiI5rmQA8Yg+E+Nu0ruFXj08y/xWrh9UbTcNU/KhHwY6OI68GxOmmNoW
CDhlK1UCIi7qrLAt+MutfkuRd4uLq3M41+ZkpVwtNH3VKIXhx0Zc4KpwtZW4u19+N/8Acm6Ihv96
v8aVL+PndF3LZwsOfBwxfmZ9uM+m7oz+cmiYRM7w4XK3wwhaMTiZiJroMNCOfY6B2BSsWtXZ2G0b
Bd7PrZ3r9ptbomwLaYZCUBxqxb0zAuUN0eLjtgITL2V3FFVzVy4csBllqHJEM3BRwJMfnS033Lam
3wNglHn0yn4mGKfAdlbeynHP35c3L6e/WVdablXsl07mT36GjKHY1gORUuLAYQ1yIy4fMI6x0fl+
tOrYfH9+rz0YXrlgKhAPVCUnQPGCETus+QTFYqirg4tZmbh0MGZptObhtECGoRzc0/fTWE3qNRF7
Lz8YPeXOmo+8GUwyicFlkRF25fZIfMpal9UWKReG6/W9ADOxMHkYRcPHxsza1hFMhu4qXsWc2O/5
r+0+rYoYmQ/Ub1th4MHzQp/cXVgqr1Zc2T+qVKu1nD1OEUUjfVsHSW9v+ApWliMh0YJ8QqS5qjGc
Gyp4b5+ErWP/lT4ilUQ0Dej5KqWcWWn32omFsQnmE7JYZcqlUZlcBhew1on5I75hsUphPalzNXbK
P7bfb3vuXJZhl3FkQ8GwzgbSEz4KkAOp66vjMyas1KDra9k9uIKCmSilHuxBVHn2l9NCgFnopF42
xQCjPlHvad7DQHHV2xSABC0HXRJrxaY9uvpai1mzz7LyZcRHwrgbaaCYwO3/pE14AtyeTMHSDSCM
9v33QMXij2mo3REQm1CmHXRd6Lgu4Q4qagbIOjnOwd7iaemLvl5Q+fCA+e3nh+Ngq2cm/Ips3hAA
Zr0J6p+gbjMaY9cEfevZeZ37rnja1qsD6dM7p4a3IKfn6mXZrv59NyXjx1NcnCMXaa2MyHipeyoB
ef3oqRTqmMHsSRlhjuE2XY95Aaj17SpUhj3UkDLcZ90iGj7PEdfDsRS85O2QRCiCsNXL94mUg5q+
GFl1SGWkO3KsUcxBh8uYj0FCLZDBYN/OGxFpLiOl2v3tXqpx4HVZuzrqik1tzuavVhzzzdwdwlGp
AhJL80JRwJ8c8jjpnI8eCbGRQo+q2AZjGeuDHsoJdKIhNxjLsDH+tpObwxKRw3p3CYYLs89j5WgI
Vf7Qk8Be9IWoj/xs3VzHCh0MSyjIKSMlEGcjSOOtcFFm846wH+dB1zt+P0Qq/lTExXgQp9bfhH2G
t8lOhr9YoET3XJyUzTzJvwB7l/Uxac/VNdfX+TkMXnpDffj1/0OsN92ta6xXrfGK9IkU/8XO4Kw9
s0TniM9ew3GFaKr0Ix4xtG131UALMXRUBLoDVB9OJLkQwwAA857hzGYZKmXSMo/LuiuMHUAtgz8c
Hooq4lQ69dly3ucHPPNUskN9yjXjZA8AoJeTMVdI61qG1wJd5Fd0LpJtBLQu8h86tkAmynyx64j5
CEvvgk2eotfyNNQ8KRpYgS8E4ukkIXaGUiAe3mfkTGxwNpraLQcV83BtLvjMag1SrrZq5MHCgbQa
LbqN6I7nb5KQxs6m9/SJWulLo6KqoLzomgNmV4IS8XTP/rFIBajpf9TWP4lBoxUdNFds4mQkdBn7
cLLF/QEU0r/D/N3zBKeDNkAnEnj7PmdrlbB51nuJsu8r+YEdpWwUGPppkFL54feWCVfcf2ZxmLfC
JzTCJsXtHm08xX/a4mUg+prBXpxyXhy/O7WqEbTmantdY6NokNpcSnqu4xgrAJ1b4FRJ42KiEx7o
feGawCmSqL4S9x0R3lRbLlrGPXW57tKorIXAjVN2a+PxTqK7KaV3AjqbtcPhDOJMAuaBlaf59UFU
LEAJ+bJirkKQ1iCbHPJ63kLlG8uiN2IkyWgrg8G4yZmKkqsKIhxonAjp5UJK5SL+hOVEzp5Rb+MZ
Vixtq+ZPvRLP0aOAvPVLpq/NXfsAfpJwNggCyS8JUF2SfIsGGq3A3rqB6cEmvyWYBeSa5c+VcAj5
GQjXW8J5zEZQX+HFRQKZ3Jxzbrw6XfNoZa7rajx2V25BlmP7toFD/wLJ14LQtI87HszMEVou8k74
mwjpyCl9CTOALS+NTPnH/1Oip7xFIHXM57ZKkw2qBosOZ4t+bgyY3z7eW5eDqINNR8tsmDyUBSAM
9dwr1lFoGBXdf9RPfUe8pYJRZStHCMfJdnK6ApfIdFyGRa6yMqIl/NVTpzw/ijIv6PV78bC21aBr
sjOAi9YwDdX8hi29kipHAuud36iodAdqrAAZQTdB3ABZr0zpJCL94iR7jV7ptlCfN1BGTW+P99hS
VRsdU6b03oE6W6kmdvZRvXuS6fcmwwZ4Ow9ADVpi8ghwsKveZ3MfdTkhRlhZC1fc3IzCIqtldVCl
F4e9hHYFC3NtNPVV5s7+fm2gc3PsxrpYI83wRy6YowXxRcHEmOE9s3MFGM5aq3ot0rEH6WiOr3sf
iHclWnuAMx74Z2ZN/5sz9rLAHJdCYj520A3uralEyeZdJ1ag5pPoyJyBq+rx/aXVK0mnzVXnJ49z
xjhouQuCft8xrACmcntKVh+YDeSpQEa5rss4vF4MkcuTJK98GUUfInk571kFssoDSJmRPTzyeUXU
l4w6taq/NmpRih3WELlmKHsgD1PVlNVqriVG2so6Y2BjBdKXIQUpeaRwD5S63/THbQWnmLZp71Jq
xfChUV2bTxifRzqLqSuTTjrAx+Z1vOKDZ6S/gwE/3X/coh81Zaa2N6lV+HQR0JfagLfnx5w3cbIe
ej1AMVKeFbT4B94wBMHElhozDp/B32TcGCkb+dKnlc9ASDZcBWPLpo1cxofnffw0uDWa0h6/4lQ1
Cy3bwaUjGQQlLeP9n3CAPSqgjdp4Hh5CA2YI1yOzeGNI9VVV3FBWRI5u2ANktedah+t27OtYlV0E
9FA0s38X660oBNCgjokd3J60LmbEiWaySsXO0pjFDMhoy8Lkm6DzDwJ+EkM8qM6Sg1gb6Tc5PMGW
dWWXdQjPNo/Y//XZ2D3H7yvS/pMWjuzVYC+dct86S+uEgL8JN7e59QaWAF1pHS8zd2MDqOaxhfbs
z1g+by7j6dbJNRKKfrPwATzt4tTjEaPE3oXJ1vIS1wJAKZ24db0ET+Txj6zV9Dj6C4hbmbidjENt
36B9/iHVqpkUKgIyjmrcIDc1tesuGY0Bz2lwLYRlaKRJoRu5mb2OIqa0unyEEAHUeVUWyn/naR7I
RjIyb8vs0Mp2oeISL4e67CeE+DlILaCjKxUfhL5keFap5V+i3Attr5apOijFWi+4VkHeP9HOcns1
eg9x9kXHkAbDJc/0kOy6tRlJzodDFNTivlhgvOh5XKT6yGdHEu6wQCbySDnwJYYIClY08gxe+ztB
szsX7qWGxF60D8M3K2qIrWoyJNSbXEAVAfssLJTZO+H689Xs7T87r1aGTFsqHKLAUy8jQHOAXekY
ue/i4ICWz3Q9bgaAMtkdXh/GwB5C9GZYbP7kAsqyHSZOfXsswKujbv+COZLSoj8AZ/jdK6xH6FVx
PRW4fVkZSglclwS5XLCQPX4Pxi/naJ+gcBPlRr6HPw8OyrAfncrXv6XO6lQ4T44jjknVMcneMJGX
nciqDll92xd7jkq/UFGVwADkg6aUjahpmIOcphe4s9M2satc+SWOk5Cd6f2eA96Bfdrya0Zznz5E
1C0+VnQCMQp5GzgAZaSMm1qtEqS7NlxikwZmbLP/g8H3utIL66STWHVdH6jory9erxZA/KiB/FNY
3MVK02y4A3Fb1ipp/VmUr7LJNuOQP9Ba0E8vBrL/PIiUrdn8UmKdCg2NA5dYkHIBR0Sp7zd8x9eS
SIktRn3oeb7gclEra5EA8mx2ces17JgjnsMBFXqelIvn2RF9EBn2oYUEwFvkJuoXIF4RnIsxjTud
TSacuXOqiSXZNvb3Azes4XLIeK2Fhjb3d05CaSBjWbsCG2RCj6K4jT7yQu7dOEXwD5NSC2lHukwg
R5q9cMabDDKezew1rI43ZgQPmJivHyF69YOhWFT7ETZ0x5j4LZVQ7Vr4870MtfGRGG4pgJ9Sx5IL
NAuMmsNcMF8mw7QBq/jZUlJCNUQtFF7dsX30WhdNX3aGQJ4jrTrDzXkBTh7WpJTvKah6CamSbMCA
J06plS6ddfJZMiOaPwH2Th4pz7epRsu2sgr3pAcQDQQpKxEITUYNLMzNZKmVW8whBh7rH2k0lM/H
L/AVlzHhbDxXCVhzuLliO6Nvw49ZrL5MrlfGeNwSCg63JS+llW+mORrlFNVo1cCZgRcJTf3CISou
9ad+JgS04EQzf+i8XqklrlKc83vPlwmNWpjvr/JpUFiDsIIQbfoisn5ZLC0Hm/zsVMcbm92h3HcL
66PydQ3w/cykxL1dqO8fDkFFJC65008lS5DGwpBaokBmoULybieye8Cm2k0RytoVDUNBgT5V+p9F
DbZsprUUk6gOgkm3fIp6tQ7RS9qQjDqp/kU1l95NLwGNUiOhRpor6rZ0UJp+Oi4G9JNhW5EO8dG4
paNGNcEvcHihor8ZUqnNyWP4+aChiks4ctCX07+zVWcSyZg0tHoGIoD493YuWRMmLMjfbAVwZqR+
u/+E7GK5BEKcST2+VCm4jMaxT6jD5tKvk/VziUYc7Jfe+gBg3pdIA/V7uodawzwts+jaLhtGYPjE
9WyEPjyA/7HMKDazIP6YuT4KqdsjUSu4spDrFLU1NlQg3yR0CEQb0fYzaJ7aekXwXWl8xyMSMlZB
Jw4zHRye2jhEXgNjGBClZTgP9XwQ7OtjSdss3hsSliHNgcyoQewsevh3XyL4AlMnyqfKpJuQtCCN
iBv4tEyEe1iXkO/6VOflvvh4Cc/1BF1f4aTQPlkqkKZ8/C3WnfqKSaUPEqs1EaKUvdu00CoZaj3o
4mviJLRKLaAaQ0dQzQvXJNf6xDgh7K0P+XSG7QgvJaKHYe+oGd4VQxFy8yH7396HsR3M0pTcRUH2
prLWH+VZku6PpY/7PjYEqFCHMekPlh8/c0B4OwKJRMeE6TonX36NAQuHPROa2GhRUmVzGuOpyj1y
YDg3qts0z69F2QL7/Ixuvcajg30tCY6Iba5C3LhnASOkfHhtlqBaSf9NcfnS4Gr62563tSpMWYFO
goh+GUZw7+SWwsiFUymz9wKxK4SQM7IeiSeWtFnTgutdh7NF7ms82D8s6ga+H5iIVk04RTtODOsG
Zr4G0QfvQZ+A9aw3cElDttziAVAyGGolPQCX9ZmfxPHBtlA5ab8E37GnLPq44f1Ggw91itb5pNky
Lfuzt/OaXg/ngC2UeAlbHivCBHtfSOcsfe0zTkxdjj2Miw7m/nHsDh4LjQTMs6+/MBfjQhsBWC7G
GsFaFuoeddGKLSCZsGXOdAD3+oWpE0ujqlql9tUEmr969/pHZtc7dFtEKhTOe3s+XxFaBwiFciJ5
oDhI3TRPgOGaJs0gjYdsNxowB/pIYNbBgUMplYLU5P0Y0YPN/m3El+nrqs0vumAsuIdeXFB01VTJ
mh7huA0H+POg+c0d1app2jzSLPmzs5/dpgJYeDkkrkYaldb1Wtx5io4FYby73aGm+J0BhHZWCoQY
1ryZVOlMJJnc39s7k7jJoy93KTt8QZ/qtAiv82pzX7l6yBFB2gKnB4pSSjOOv/KBxZX187JQAvey
+8HJAJs8AApKv5uUB45m4fRefzdhKc2N+LOgSE5PblsR33eLbOZ5tovEPX1pb3hlXSFvFdPcTIQZ
rOoVpyoIXdabaK3sCzve6iSt/HKkrK6qoqhV8Y69IbCV9VYjMNT9bMSrq+1n8PYUsEZLwbUcFXq+
+Q2oEeKMLzT13PFDeGkOgnVaATyCAGjBwURPtyRBZ4S6dU92QOG+waqBitbsaHS3CI4hXiJSPswC
nQjX5UU0IwkoehkiTIEoyi2s+pPJ7GRJwKv++beNeCRJIT0Y+SSeDOY4U03JOEqXDxAS9yO5bQmU
O2Fg6tLN4rM4PNfbIP0UgA+nDW1vgL4fv1h+i0BHlGXzjyf6563qHb+0rpHCVHZe/LWNsb1LglZK
4Ji8mg42e6IiUYX+hGPcDQb9AErlwq2dHZGZaKxPwx9j0zZJ1pBOQ0rqPIMhEHi1nNut68A8zUj2
A6nnl7re/l1CvyaQUK5QRb1kAyH1gSrbI1Us4gyenPJ6BgVxFzwHumxJULF67cxX/ymoIiQKOWo6
Svsqrq7Q9jSvpaIynAB3e7xIyovXrpQVGSDCDdd0f5Up/WFzjAe2DhTv5IxHJRsYpCsL1G1nC5Dj
CivgexhPrwx/dQWfZSHgXTg84qR0nDVUA6LygNAHK2HLCMYsCVQFUcjYyso8LprB0BR0DMeZWCfQ
rWQurkuPb7+KuurLXTZV68gQxQ8XdyYqZ++1UEjHD/GxoTH0/T/a2bPrnWqtkazd+B9/2DyFoPP6
oD3TuDrvVac24fRX8jFWnyx9WuHdaDjom5h4MeK8phc89sqBatwoKClI85f6LzoTZt+TY9QV3b4z
8gktvfx4jn2lgV1QGc4DeEHyzVHC29CcFbArVzq8ZsMUqS5LxYYI+8NSympTR73aXnnnl29khrEh
khNpOzsk/Zy0MXJH8kC8czaK03DKBsIHPsUp2jnxRSqRSKiuwn4WsmWJLHP0YggT3Lcmm6wcGoG2
hY2tfZpEheWi6WH2vcQuUuOC4TJkThP3/+tflKu+Mz06aYdn7u3l10Y93RzdB9VAe1+7RDynJ7GC
oBVRo8rVjypKfb8clplLMyVjNBPTN/792kRcA0oIfyzKwK2QMNw3XYaLaZ4jBnX8Iz1X326KFWee
dcK3IogRNt7HnSHAbYZFWwO30O06Ct9DKNNjVZPR1o/WrogN/wGbDdm1Nog+T7FjbFvLcmJ7ptl5
hDyBx9WNA0JkEbqyBpXS+7LHrK2aiC4V3snjROjX82yApTVkqg+C3DJBkdaSGZd6MdEz59YapQax
0pBN7pmsFHRXxzLiIbqRhfuFSlxXE7I9ygCicqddlczIEik/o2CVz8pWYT1fGLxxeOafTMhzIca0
FTwro0Euam4tKplxD8b2c5DTso2hYaJH6yhALLPuvSZdp7re3PRF0+EXLcAPuGK00U578ReHkObJ
lxF89cROZWzDJN+NjA9Qr9++68tZAOZm5gV48DMUh7V85pn1wmrYDpxZAPKJaw97TasIyiltJ9w1
fMOEivGwFDxA5X1pLht4iRzEZCS4nKFTa2RqE+rwwqNq2CP0PT6U4fgkuZHZ7MiiVDy12Fjj/Hpo
tEftopxMjwUfH62pOjM2vnhhHbZXD3Dd9EsXg9dTXAyZyUMnwZjsRbChwwtltjql5oaQW21fa07p
NS9ysNq9951RZsk7+ZX8gNQ/qrEPUgxPtxuvDiiJ8+JxOg++oLaIYWRYaqXr4vmUl+XI3zLtOB1j
1y8KO/i4Vjqi88p3BPe9Fw+74mTesj5CDuM7RZ/D1WPuRt/dM5rWC22l13pDF8wI7m7pz9ibkJok
x+4whlvgAYRFq0F/FEy2f3fRW5DU4keehr+JudS5i7ST0IBUTz9KsmnGWhYRjWtdLNT15Ti9V2/a
Z/n3QIg90dkaqx0DeLxe/hmo2jNUANX9tassqOP7HBF+pXW064ENZdON/vre1BLQuoWolvD0GER2
KCBpqsWK1JWly+Q58R+R9hQw/HXoNPBdOBB6DUdL/5l7tMUuAFa0dB38IWiZx9ySJYhhO/2KQMU2
jv13+cQgyHf+rMgT5id3Pu8f0Khk5Zz0GkDUoWIpKvJcLH4dr5iRKYmioh8J1iJ/cuXEdXvGmJee
4Jm+RxuJH5cNL2gPlwCzAZ3mpnk8umzjuIn7EiReljzribgLpdCdbh7Ty+OL7gTLqWREJjphQ8RJ
hRua8/OOR2fVWgQ3hxx7WsQKiupK8XlefGJAfCyIq20VpA575wTMaHFMM6yLovRv1wi3JZppsM9b
HF7vqO+IoJV18aIru0WszLc55qw/cHLt+a4czk7n13Ne+EMm+2y3GtPZLpLS2CX/eALIpKlWu4aN
CcNLE/iGWeYufGnXu/vSbX+K3OY9ETaEt7LHA8mN04kNf5zegenh30OxtEDZohI+U/rtbJA5v/MZ
Iq1fjvrM4DHZyVr6YJswFRvYsWNLL9u9SK7P9Bg5502frwIlNYGAL7dDBjHJvAdSEdCWui2KmHEo
A0uzkbNxXYpzv0iX1EDMuSsP24dLebUoNo2fY9HLaQStpyeoDYmXoaG2pPU43FktCqnr5clDnsuf
wGtZ/E6yiYY+KRV45Cvv3wzLbQvNCrSSSCwqYUTiB9hXio9RIjt2dDRkhqMdSg8osaCV5VEJmtEj
tVdsy5tK3vte5sEkgCYHMXnUjp5UBI4Bi6Iqx3KLmEkEixBcvRdPlGW8hw4QfNQ5vlGWBSRUehiq
hlVvE+joJ/63VFyjNeh4NdW05+RxB4n+hHTTTXCNDM1FiWI3wAJgloi4pxT974xv+Ja83zQOy6ag
J1ulCwA5NKmB45iygnASJksaEsUPnBB5w+sa7kCH1EU1dTuJik2DNJoxIekNwqi3ILQhAqcLWkFr
ugPb1iizokiqa+O/A4DrBhQGp92bUiJh1wZiKRqS9JgrYBkk6I6iL+/SlV+SaldMA9O7LURz4EjP
M+C5z+65glipbp+Hnam7uyAKxzYvbuFiqtlQxyl8rgW+6+ZCW17yuSRX2ca5GwdIQU94pI9pF/f/
D8+ULbyUC9r68l+S9vll75Adiw2htXHvlEOiCuzeAOFyNFKMe49I6jnlO+YfGl/5NI43qjn5Ipj2
5CNRJETdmDIj+s6Mzi7oQmB5wMsbifCMufbT/clSk3/+B6xBbLbpSuYwt0g/0jr22A0fYFSKlYVO
tF1ZzQNbHao17a8Q/fJfHcSsG7XbE6fdaA2MZjfP/W3DDHgUxZHo+WRoIJN6Soi10x5UXN1c3bpT
8CBd+kYypklUuV1iz2y3k8lrqIN3Hf28ZIo9GCWkZJaUPyT84+hhO6pwrYIF2wFovJ6BIOYyDZU3
ynSbXKKRlGx1s0wYM2K8P/Nj9ZmTBlYfC5j2ZjXzC+cZdXdEUaqPthSI9dsNakEjyJFgemtXlsEH
Vf5rMOJ5ZcR3BPUQZ9E9SLrXhjHO0fy6L5+DDlMc5AYz1W8lXibYq9EXu00LeXWGfdlmWePn8enG
tN9Czu1ro5Lglq961zn6U8sBzppeSwG179EifBbBhwrXoCIJX8OlN0YMLjfdnxbCCsaxB7l2M4BW
7vpyTs6ZKEUlCVN7pqFZ3ICF1XbOuBuhZdaQ8jF2Ort3erebwOC/5Sp4vDGHT2iMgyeeOP0t2ME+
2XfT2FjLLna7sn8X4hJkhUsUK8qnjFoGtU1ciV+V8t5A0VfHxGg28KDUGlbOR4U1oqxmaUEGyOj5
Dd7lrgUnNLIaLqG9zjAhceQ5FX3+wgH1qzTD+nyOoiwBR2DLYZ86liLzI9BsgLvLRY2ROqOOJ2sb
u+pEx4GTYL8xLur/tEfmbXYlxOHgvCV7D1fDQbGvR4VmyQUHmRKZuvKOwImMI5xZftnxkHb6R8bf
SMwSM3llngHqAgAgc4VcmsjX1AnHjdTBxaFLqddRWCQe91gE5ECjaEIIxlDoigyUdK7Dm+8s5Q8K
guFHOYuHLAQ3quzgy49lDKovfhIiPqZQGXTa8UpbwIf2gU4WqR5x3cbDBCAyW161cIrhIjsH5Hqa
3BNEscG3GKMtx8CVQMy/zy6cV5jQHhKWndtPxmIKN7rP8m3HC5vnHoeyOjh7va6Bklw4r6FCvXAE
cFlk9MIoKgPEZMDa9JJou/rbZxp0U1rjHeXhYkybOq5mVw0L2OELRCJaxKF3t+cUVagYOLVsBkAY
9g/mWrUcBhxzzNPYlCpfTBzjycpwQLbV7lcQe6F2atHRsPWQdOJnO7dN0g/lIzTkxvhxQRMXSxJc
tY9DPzQvyJxNkVPU6wBwfLby97AzYvbAv4BhPTS1kwjVtMO5XgalsxeByWw50ORAl/A4HMh3rS2m
9fVYAz6Nt3eHLH8M7eYGi03xfA05o6Z/681m6hKkNWbYuQLZjWnDSxyxKegDaQZM+IW3UMsLDrgM
IqDtb2BIrD+KV3hZAphpU9FhRlXy4+H3fQR0qy/+JkM44HIlSaOIg57zywUd1uoK8XFi+B0Fm1aj
NuTAGoQfOqsCSt60TbpDBtzaNMDk+HJ3aFvshDEr6tRzc5N2urPNCcyIKj9xF/NHtTSo8aBMu/A+
/QUH9dY1IWuhHOu1i0JqhIYU2+JtazZmP0Q1nNYFLWkvs2of7U8TIpbDeJzFHTHxP/QORboOrvyy
GPjgqHj8+z0rH3XVYQbBzNDJ60UmHO7AgkVTOn388iIExvwpvbHoz+QBDusPgoQWkJ7jOgzhDy4u
p5Uxa2GFkUZnRffSlxyu2bmaEEZQUjb0zHKTzF+QQXQJUXEnya+ir25Bs05qKzQr3q9wFxABsi0E
L4unOQia/MMLAz2inZqDoB8tpjmh4TGul9f3wZxgXPTANPH3CPqOAnMsYmtSN46MwfQKHpnBuOlJ
KvHUD3ejXKiZDUg5V78XDYG/6L3+LUso6MqxMFBjyxtm6QMXZNeF3wffk6OQ7LGnNQ50Msf4H61a
MJ14QMA2PdZiFv7mzNaT501K0JcM5M32ipHgm/J32++gw8K3ImXncsmG9Eb1KhFttgVfFxEpIAGM
31lgmPl6+m++O5mPnxsNCqplEt368R3G6Myz2/qjPOI4E9yaNGaQS1Rtq8w6UM33bjtYDO0gWqZt
zMUw+HPl11abYbcMKtMMHAdLxqe9mfxZwfToWZxS3Nexp1MkK07dbzxCixLyVkflS2xk+nuiL0Ir
mDasvEfDiz/dAVBKIk8wHXVD/I+3QAHgtv41gVXLfM+4QmjKYsS4axZyXETNAVqdTc6hyS9Qf6GO
rIkt2Kt04S9gp3vJCJBukOvSu7cMR29tqig3lswMFbRZAgpmNtg7srAudDjgpr6BiT600dasJS74
914z3JQHfxEAp9SLuyLw2pShFWCeVw/0M8JiMdq/4B33PlHGJKUWNbObKk6u01Lk1wfUC88wM5lG
LELcJtbOAslYx7ycOaUQ42SL1FKpiaODtEjHrjhvtNDh/gtU6QWTL6bVNubVfjIeXl0kyc3hk/Ow
RTt8R2+fvqnuicA6q+GKVxsKpU5bPlUmE2FhIG9dujHgDbUCgCukaLjttlzw6nsQb0dj0hPOu0FU
2Qtv7AZONsOS/QQ4DBoUFvaCDBQEvkDe7xJ19TX53HMsCqJmH6tS7txpjKaclY2bBX6Qw6aSu/AR
8atGK9t0rKOC0FmRnavGHm8Eqwgl9ZQW/xcqpICnCaFA3OaSQ0MAe6vCfX5i2kwv41meiFu49RWL
qC7xzCxwJSMeSF80o8PAe4oufoYVSzzaPcSbEiJGxzCa0Sb+4+nf0hukM5EA+q0WiZDmNjPa9OY6
+3F3vqeVk1p5dcJUo70rTrx9UeIKC8wNG7FJxH8TVqOLbFjMOLK82afsNcuh+tpNkjsWa5v47tb7
Pr2fnynrZ1qqOpLk0AHFBwM2//herCl2i5a99NbzkncfDiZcJEM/NVK5B74mUk6Pkp7fTwBjBzNF
DA5pgkSqi80Tpqi/ucD87GgBwGawT+O20zdmvZ9PWCBdDvMBQvHxV9+pjvxTh9naehAgwlncIojH
kTiHNh9lvLIXipS7Yswl7vUtM70t1rcQCf/Xts2SJ+Z1Nkb8JHm5wQXc+jCzJLU8g8AA3Vq6JkKK
Ew/Uxks95qpV+vZa4EEo8QweEJwY/gGFQhiDt3FVejYvh8Cnoa+KUkjlXhXWTpZg8HRkjrpupgIy
qcoVR2061ApO5yU6iC/Fg0SlQ8MM5Dx+PKRzPEzFvmpgi70RGG9fpQFNULSoc9E9Fm5wxY7M3TEp
DQ+9x4AEnI4XQLWaXYEU4RsJ0Dn8Udf1t9FfQz8MeaNDnHNK9P48opk8TtoVEC4t0XcMW2g2KeD6
JPW7JWgbE1varrZ+gIFTKlV5WaffScyUK3zee1D8uNpnjFZuiM4F+rjWSBhG1ObwaMQEep1aXGIK
pkvBUylgm4x6SxhcRxdDkza2rmDlaSFIHpNnM1jPJDoIRy+xvWCnS9IFDyeQJmlNDmXVHlVyMqbz
3/Kz6U2UoeXXOQA3Oytbj8n4owzMd3tHOxPlZnGVGxQVZa8+4W3nv8Vg5y0cRn4Z3/9ac93OgdsH
Z54ejPsDOtmdj1NZ3PSzH2mbN3v4OVq0sVm9N1WrQ4vD7d63r6R/TzH3DWECXBccefFf43MJzmth
MM2Eskv5H+vSm3/OSeImaAYrurYgw3+ypGMekqWs4Nhm0c88WMRjavRXwwhr1rxVHn8VIozzyPde
u5AsH5UHmeLXZxCHxKcpIrWx+UbbU+cwqI90Rp06AYOub7a4nSmMD563DJQb1h6Apm7BRPl/VtQr
+v22g8/G6z+RMb25ZkUR/q/nTPUneXYUtjVRdgJvXDgWYKGUXRL5z6FS7v/+eD/xesHV4zm2RQCx
dC1/dV2r1sMCjo5QuAeH0MLP4Jega9vVrzaGKVvRCGVYIzYmKUq4MRsMEDL7xqjBgmXTGZ1UcaZ3
3jZS4aYFJ2wJiW4PBzzg1SBntN1IFWaaI2Gz4UAid7vIHMgrYypgsXocQbs4k7FlArDwZNCHQB8r
CDDQhUNOimtAT9f+KrKNFh/vnecZ16eDAbTaA3hYYLdW3IIwsvA7JDvQQeX8Y0+qRmU+Wmlf/TAv
gViyQHNJ1j5fYQjIrJEZqyRsZfjLXBkOafwZ0BlgBLrdH2Refl9uETNjHSCcdwp3CjSByCqYEQce
1Ah7ywXgc2sBXRi5/0XGx8+sj0qlQooTP2uC8sab89PrqJkHir8FapvOcphwhwwWlIi3Efyyk2OQ
Wmc6P7gSoCdsOdJBMyd29LrJToj/12yvfV2ouOi5Ped+uQ6UAqnhsHvL8HLTrqe3RSI1nSZITHgU
9B7h/b6Lm6PaYtuTk8kNcmFdWTUiR51A6g+6yKEHOINoPU0a9OIaE8EYEc0uk0xDpyTrlPUhFhQ6
lQGOASPbN1k0bcWRHFt6hBPmVOcDqqlzG3OA9AFwhcLrhjLPeLytNW0/cgvfagWF5wgGnyy5WEBy
V+hdb0/VY+Er3QHFDkYOdT3hpK1xQjXDNa4tO5h1H2lGGICaabYm0Ghd6Fdnhk+BK9IXsmMJTabG
WPMADRZx8q+FhtACxzm9ymc8lLLtwCoG2PYCH3gj3aGJ449nD2sf4GCo04dCFmMv5CKLwsJetpUe
4VOWk/KPQOqZ+N0xlzvF8HORHnFTHboSbmewyeQrbKIJJDaVkeyEvk66Z3AmsmlRP0j96KriF3N4
r0ZctV4jp5IjYjdNmwXX/fOcr+iKjKfYsOeb4sbT0ApCjpnIg1DYo02QNjqIgnxG82hPYwRvCXDl
EoZ4VETdOMtpDonn2kmRuv7KYrJdbfMZVlFhtWf1NjrcqplUbCRJh2UUBYl5qq6JtmDrqeKodxqU
dmlwhx7b7fALwAP7hp4qWePSjKKtv7kSpKwpMjAU6E3MfcbcLydoXNM/O3sVwJn2bXl0vzx36nVz
ciMdmxkEOi9zevd4V6huukpi8HVDh328YB6iaj3WoMRyme2cDNtQxTbgnv+jpSVGbl38sCT7F+CD
f0KqoHWJQoon1XBUfHk4hxXef6P7eVV5zK/E3dVHnoLMCn3/TsrvHCD5MHoaInVruFN9gAwstXJZ
hUkKR3MwrwwP7zhAANSGrwv4vABIDaYOGUbME3+z6Vam3mL0M9YSl4bmF6Xi9jdy/dbBNfuOGdho
X2viH679upA5q4hubOWbv1JF2icJsaiE3T8mwzRpfInfii2fOBy42AF9eZNTkcssh6pcbt8FDBsB
ocok/nkCgC+fPQl2GFncRaPAXx+kGO5bZNcdXuBgEeRckorRT1WjA+oAh2YYm3VUkrNUDLUua6QF
i11TomOjnkgSpa4tAMcoElGS9gO/t+vbmbrMS+DKbmRuYh5QLqsqA5eZ2z8Y8k9Cjcf2JcsyA/xh
mpmEKX7hzd0QR31ct8/qxKp+9PXceZu3kVn+/hV4bOFZ/4GQHFZU+SHhtCxb9U1gSoqDQO3zjBdB
ksB6DHOxfS948Kft37sCYddyai0WikI95TTkRGIXspVE0ZmIr86aWc3yNYJmdMN+N+pp3HJ7pBxF
zueD1YAaDG+74yDGVOVz7zEoGO9O598DdUi+0aAeVm3yPhQUBAj9da1PY+38WH0fzsW6aBuyhw1J
jfsS5GIkI/pQx+hOTeY7uUbwJfrTs4HByd5L2qPSEgq5jnZaVlD1LN6XuPC1JTkU4Sa7vU1+cKXl
YIBglR66Q1fNB+AL0XwN2UuPBhz4+xU8O3mALIaoNnmaHYi0nkhRn8wdX8p7pbY05nSKgkNFuBw6
57UkZN6QSNmoygUh9Q91tpIhxedgHKh53OyULRTV+qfIJq/6Zn396EX457LmaaqCkwQbmONQ2Z2F
Ix++gkOEUYAmp0h6vlhZsHGT4GMTHNgb64gwh9k+CCniyPwM/ClR7Pp/qzSG1CEuWyecl4Q/b+mP
RcNNBdc/3vwNpE+Ne/8VopJmyc/C28oCO7R13b7tKXEm3SS6SWJ7NXZ1ijeIW72nfnjRBzB4/6Ps
VpKdZW8LZsAoGGD/w43vKlF/yU81bDpC53vFoY4F03GZBOoIBbvhXoEs3ZNQeUruIXl75x9EV99N
W9SBX7ypZwTean/mSpgq7fzcadDktgOAbVxzZEo6iAF9riWfVXCKK9cyWjbPUWZ3lM8cmfspNEs0
4gtL21IJRBjxeFpsGjAPZTZx15fBOznCZtGOjtPGdqqXmhPoFjwH+TqMPMJRlv1pkSs2V7f14Q3B
kOQRsy8nkxycaCM5RgQ0vX8TCbFniuRt4NjVH+zSkRwkij+4Yo/GlkEIWGLu29otM3IN+iBnNn4M
P7KOrTN5EAldlgwItRZnzHGSkzp3qDG6FKgsluWReA2t7/PPBpJ1FrzABZo634hVpSP7gmgS5Ntp
oDXUKI9uLPdWtWQmzclL93XLKwIuBTk8X5WiSywG3r6llkxoknm96Mac7+pLLu+5fEVO+kAOtFWH
qcKijCc2R9b7aDRfSnLNSDC7bSbJIdyDFZtjz9KwGGe4NLZ0EW0yfqiPKQrnGexdf4JRYz/B/tLJ
LLWDKStyUuTM5DBF5iGDJi8fpxtGQtUoNqqkR4MhlpxqH0/VuU76Dxv+9ZXK9kQZ9kL+Jq6zzrx8
DEi4vYFq2nR3mRhb2awlDtSTxmNYcukrtDyCdkHg0aI9hOmeViffRnK8aHtjchTQImj4jVXd2jYl
Ak5A+Sc2f11jt1DkbtgTrK9vduQl9Tuly3FlFaSXgZROrt8Yt25xDoIU+BpewJLmym5ziELEtlF5
VFIbgaYU3JO0YW0dbmQxosccCwDfjHnroaRiMKzChAXJ4eEZmfb9axefVqZX5GoWEKqB/7r6/Gcd
aM+4zCNB8ichcsh/QQD8ZTmBBbRVFqBuz+QLRK89+RKHDhY5dV4bhlxHu3YT+gtT9Wet4Pc6jhkC
Bx9qAMKu0JDHwhg/wJiOQ5h+mAVd4Pb4DWfh88Bvjy2/cw8nSYRTCwc7f1LBX0XSMV+XzrzHcWYy
kRl/hBy6qcB46qMZ4wuGHZzYgOSc7MhMKJeBMMqXIZNWiD+meW7yN3fphSBJe69rIhOOWJL+1Ybb
dw/PYJ0x+P2XVE05ioQYzXj0CCrdnQlaQkQUTY/RRUX2EM7ILmX/Ai68x88BBBUA1nWFjQ+tHe/R
Go5tPT9M6OGq5eGm/CD0IdYdN+ScQWcfti90MUfIfAGTo5Dl8ktGlTrmmagfsvpuOejWEPT1D6VF
oL0DMswJIS/JN2em66ZGT5ylTHzjiFe5t8ZkOn/c2itlU6yH4zL/tYaF38C70gTllXZWSVXO3OXj
1xF/S3x+GNWXseARgd3xUgYHIjDBhyLHR/GuaJtnZMf1VDZ2TrmZQXbHTc4MDELfVcOeYNArIral
wEjQnRBjSLW5HyIARrWy/o9H6EVDG0Qk7Vl2bGjWUOvw+s5M+ZA6GvEZLD09fjhsnCZKti5FR7JV
/xA0hFKnIKlGjN5C4K6ngn8isfhtr2YA/07DAQ9R0A0KWS3ymaQWOKhHqakOwseXAouWjbUQcghv
5naVjr1mIk7fDkWU+QUJxx3w7OCq8iik2zXTidjcgZogfSL7WXPszEIr99k3yStB7HooAk+r+zcE
3rUsal6P8X7hSMWpgysMgxYGODXUEpOg2EYv1zIxA1SVO9R+Okq2syJTiTUIYvLm41i1D2qlrMqX
Oz3/JKjupN8k08KwL0OrLF9MZW54a6RbytRObCeUD0tqMvfqckBNfEENyUjPUTKUHgFa6JyFnG9B
EeGYjYXKc+TFE/9LvBM9LxhNoxovfkBYt+u2IZBkJ2oWS/lXN+KKWQewEMeng7yN3/l/wNGgxffL
p3QFTfajUTTpNSpCN96KKZHNefStNq5DQQ8P5WFR4YBpHzkopS6VjzDzQGn85LpVl8eKeE6TAduW
e4lieqpX+skWyXgALoz09QVTog34dGc2uVRxXNPVKj5xb/nkyZX9ZkLnaLxBpDz1kl39is6MjLLF
hN2CCMssTe9F0p4UjjGhcvNimhCp0CopzifmyI9qYwFezX+A/gm3Rywc2hbjKFa8jK7O7GTo+1IU
eUqP2c5ChZIYyyrdwBmLhQH8DAaguoLiVZdNTk9BJR0poM/CuMx5tG0xDeDemgcB9vXXaFTWuoWs
BO4TT+xlpRim/ZeBZLxj+36yNhIY0deFutOKf/IASY2pj0AV1YLwjCzW3TG6G6xW5dg4p8baP9db
B3su112VdR36MUV3SAZW1UR/RkrHiVRYtTfzY3pCmzIPO42sM5LUmfUu/DFrz/tNM4oaOccDiKp2
J+GeOeAbBt4pN/6fxojUvjEMRTDvJgKGh8mYz2GbNuDLTJLJmWigv92TyIGnhwCdkbHEmiFQAfT7
QOSm68Y9R7VGD6jQKTT/BgRwcweW0FqBOvvXyuYIgkXbb7n7iB0VSmd/3idXgjVboaB1UC3kBnnC
9lMj3Hcs/1oJuOHepxkWHoFtFOGrOg0tZ50LB+YWi2qh7bhHWo47KbM1yVINORustzbQUjIxkQ3g
4FdCPUzD5kR0icpDRle4ifx0Cc9F8/Qj1t/kU16AY0g5xvsME9WAArcnQV5+6N+nCVSMaQXlusgr
ei/eZTLMgSdZxG1w6uzdJmKKWQExpw6h1UNKEKToabW06NcxU5daB8lT5JJO8ZzcV61ywEypeM13
XLB2fA8Ew6mDvn+wDlSZSswxBzKkpDx+PmCNV3dNR7PVnnUaB0kC4HC6MKgUN91+dkqASl67Gbxx
G/zPAjFfWBZY2L22vbYvMnqrgGQpuVz+/XB/fNp0OBsGYvB7eLZh6RaVYTIgjWmOgRo0Bx+1Zpza
4aQhAt9qSK3+2SSo+Ieq+uKjwq3chSV9lu1m9KlaxkeTDNQ3auxN3oAEomEBVvQ3oL1Ekmy+qNa/
E9dyxIdcZXLW0njyH6MLfBJ6cWi93KRExYAc3AHbwK3cOMPjasgxPGTvq4+qZ5xPIuhg2nNjDbAs
Ja2wIc3IOcysOBr3FQ3VNqUyKlXDiGC3cUKsnlSoSD4M8mRkkyIGnv0iqJgYSBBFYqUZ5fyT+DrZ
Z1Lhwim1v+fnfYBqVIFsRfKVtZ2apUyWLWQOD7KCSJeLbP7EVamnJ1LzFlfLNxjUy45Ejy+qRqhy
QC8ONfHMMn32rfFu0p9iY0k6Qglul+1K7S655hVSs0VNMFP9C1z2zgP9hsNEOKyAT0mgn7DQzrpq
ONAcqqY/gB5kfA8Kzs4wc23uIKgCpVUrsn/CXLFTAYfrORJWYmj8kc9CeL6aE6hvo2bqiMxHTodc
gIO0H9YSZTihc0VLGJTU4riqp9BozxKCTPbdKag2kZqr3+moNIohmE7v8UDzrme2wo7VAGp0OvhI
n3j/wOQQUW62HPvrbwDg8K98GvoDXGg5liFj9VMT+9raTxaWnV+8GAJIqSkZQevtltIbTC0K8aPh
BE4opVWvQ6itSRHIdKnYx1T4RWPxKFLEu497bV8sIgIgyRSK4dk6dZ4VjgWIkfpHKxGMeOAymFl1
GxICtnEW7HlOsc7xvov3W+IpImjh+2t95bfQ6xqxtM2X0424qOJ8LOMfP0h3UmdQpsZc7uqzTxFU
hF7IkA8Kcq680RFl+SnA7/bAXI0php8nQSwkU80c366bB/oMvjaKqlPNKJM6Z9GwNJAm8XzNAh/x
O0F/jOCxNXQkAhaLMEd6JxY54m2U4ejOUtwSgEtumxduLYtEfQQH8LySeue8mNugmDSj0GMLUZDP
Ixy2PsFbVYvfOkiRobOrBmpHYkBnUTCiEVO5WkdMpj4tyJWvtjZS67GFDJ9QCmRuOBS4e0jV1PQ1
fUVbp73NAyGmCvDB4YMp/k8KlSKnHpGfOVBoyz2nZXPszc4pfoqrzm2rYqjBXSWhyNbmVvoVAIy3
YawRjqdT2BPWKpDiTetaTcMVWZtu2yLYuIQwdakY4Fa4sF25XbG/qtwffdb7uBdxMm79UG7rwbMW
nGpxpabDzOOzOn8iUNArICZl9hlvLDtS/FkcEBfR+wwm4eVCvAWxCtoNxo7J+VmZYGF4KXKjKIoo
ao86ksXkHYfxcM/eDbYotC5HeMjk5tDntpXGC7CvyLzHBwk2Io5S1jx0EMcedfb8ZprULtZ/kdGq
vqxh3962BtUAzKHlwzGNPNJU9JpNFcfWYoKqBtPIZqTr22NKo3rnL+fY3f7/ubUApx4+SgPvX3DP
mtGN+T+ub9T7kJw4JxHjDuSYDXXdayD7VncpZpb2Wt23QDdJ7l07spGXKLQASnl543GtuykGKKhh
GQJSjYPUfURNgHBvA6N0KKR0VC5kp6aMxQ+kGZrdONArLlq+7v02esyms/FF8TUiwYelQAfoZw9K
Bq4aRWTk6lFuQ8/MQeC3jQpXaw/aXBooUGAObMlLQWyizVjfT9VLIinvvyP7pDhpvYXbj7fe32he
osQSeJptwWAJ741UTnMF96DGGS2y1ukPu5/0nMtARnAN1sht2SxJXHpnyk5D6A0RlUrQ6IQUcfeR
pDqcs2cy4L28a04WnvgPMC7GnGqYXRry4TNtu9ScQ/tAvetgQFtBmlAF7skoEfWhLSaY2WsoDHHZ
v9HU6T1KXbBOfNJEIjw6tXenUGjZy7bWV0Z3oJludTUFXGCqyHUKcJEI/G/zvfp2vVOil2aAcOwL
WaInbaVYkLP2+ivhYRqegHxArmR4Sze0390z6f+6BZwm4ukN7Q6t4+bsAsWpRFVSVqthXPo91wxl
n6liarFeL6U894gCLVKeodPN0b8YZjjkXJdr6/uY88TkMUmvrTKJiu9Vle8eL8N+yaXaw8PTVlUL
2YesRJMwfb5ap/s9uVtSQyc0EmkLKZqFVZGOiGjnRk8X/71qRTLrfm3QTd2GCdkl0dolzasZ3r1u
106/PoM5F1f9xIZ8CUsUuyem+oV+haY9LGuzlkYYzYiiyVW4lqngS19bEEqwJ2DxMOwQAgiEwcCf
zPJlU72gsuRsWR4arNPhb2KPnYiWi7s8gPuc5p8LnIWXa/olEUa/1ommw8WsSsUCe96LdCMaoxQW
a3LzunYbenqvhL/GLmtbUQWHo7sMjL+M8x8aJCuaXdI1jag5r6Siafd4nQY9bCia/G3KZ89z1n8W
80soK9Lgu6QybQgDqelnElE7nGc+pjAFyfbAf6LUVXYbCB7D0XYh+8M0Vbsq1tdJ9emMRNrDkGhz
OPl6EYfCD4D+KQmqs+jI66eoEg8TFSIV+kBbROiWwPoEOZ6PoiGdaw5naAFEqPRofTiXRnKMiAyc
Yu1fI2ggNJ6AH0XrsA6wwHjjvB/achYlwQALBo13cwsXWnalq91mIbdx1jpxxNPfJb5v3t9+z/uj
49rgJf6J2ydhDmF8l/07eE5ILgugUFH0orEQHTALjt3ADOVi6EZqcjUP9lp6BZ0AdAs63bMz1rga
D1vb0EKgvcXVn5fXrpAIm/Pr0n/jhcdNKGZH3MWbe9JjPCyUdUTAriOuchW+s+KUWqBZim77qWJO
NaL+XU0VSCoQYV7LUNmLoOMQzECnOwN3K+lwtZMLH7JZrOx4BTF6sGUNgq3tNl4RTibO3QlJ+msF
ysuxJ1yNgJrTosjvpsde6TvUTPK4V+kgYDtQCiyBOWhTFvFZNy1asynIToRJzPnZYTLe44EoFIib
9dvhs+93/r1sQi24zCpFP+Z6McCQm59F4SMzqyo9dsB0SCKr/NIEDZ9eq9mcw9jU5W4eSITU6L3c
e54N40AMV4lksV+xwtjDkwh2v1pwtO1O60KC2ktWCuIE714NkGkZgLZI1h4wmaMSkj2aIFos54co
zxH4r5ZPm24bxeslXjlLt89sLhRr+CDanMr6SpI8pjm0ITKpKKamukue7drfuucN4C0WsgEoc81X
hS0gG/jqOERhKF7XuRcwWhRDU1UcqpxTUhHc2NXo+3nm7A6UZjbOGmJCMqCxIS98mlkERJ5z3lxA
+Lt6Dem3E90LZ1aK0KJ0vndAeuZ50sdTRvqVr+5Ad/lKkBf79jpXFpskfRaCxXzKrkMwfPOav9pr
saXcmxA9F6Sq1i1d7S05d9LdXcbXg0fDOs4sgwZTiXlCnqLjj8q+Bpbmk+rvGIP8IHQXTm9BSgvN
p6w/VlD26LGc7KSpP05L8vD4pAkdX63THHO18yKZGVcbZZ72oVzDWRejjETNcVo8/j4hKHb95ZfP
dDfFTuKPtUfIPfz07vPjvIrzMMrnexsozXgaqXpErHg1NdSpee3u9Qp7y3al7eC1kbCSM487YycV
9ny6+egQg1L2F9Y2qURFVDgHPHyYplhQ4Lfu5I9W6dUV8QCajhJeNCZnB8kuh3R1aPCSyX8dqAXc
WNEO8B2Za6z8bTg6uTW9xywmW69g66b1O32uQtN+BHVrI1Xqm76rEMPebD2VJ12CaHLYd8U8zMLm
DutV9zw57Zs1gBu1OKknTRHfJ0Xo5SEZFC0P/X/i4oJTmI8ByTUQQyhaOJFFWnA+pS3NdShSnqNP
YTEdhrkybgUFDP2yMtkziclZnJOsm5aIBY2xxqnmDtIU7WuuxQUfWkv1FCLsm1epRIjDtbZvjTUv
althU2BZzFPa5H0UU+hyuHSY9RkAU40k3TsWLn4N9YACBl8VNe842kTvbAguKvFTLeyVNJLFDhqh
Qf+UxkGvE+KToTXzUWDsVBCSEzUSZw9AA4E21SDXAdaVB5t4qM1i3t6S8QV0NPy8y9yG/ie0l2tG
zSB5V+EReICTsr047gj0EVbzTrghXFuxZ81v6jEwqCqusE7qAYPvixrJylCPMHgWFcr9eGXdKISC
QNGnTE8OqTlqgMNISRwBb190vSjdi/0iB7qdraU7qMBeA+r4wvl3iorwD+IgNMhRjyKflLTSCrGm
xSCFfx6i82EXPQ8Ywl0QYT2NlMmHs5QkwPxWJdwxFY7eriICTiXLzTKrf+xOI58xK2rVNu1ESgNe
BEONAbg8pAS1WT1v2T6yeapJsCioOWs6tI4gHXzHxqgRimmMnbyp6nmV+3nQLPrpJANanZGtSUqH
ISIdnKRTi23jV8WD5mJehjYhKeCfQV/P13gaAuMz+EW7f9DJwv/9mXZ1MOozkIL5H28CqY69alY2
6nq0uOqUie1rBh7jVJE/ckAY6Io+JQZqa6gh1hIKsU4mogf6yXwVquRdbBsAZ4xtYPxDKJvwrv2o
boAv6DAO+Oax0HYd/nw+0jUpZ5KKD5+8GkDAZymvJkYcfd0koJV8WC9deoyafHKa/iWL/UIaE3KW
7ECgt9SAgW885RUlu0H1O2gW5LsGFzL6PKaYYN8N4dsGClC8c7/A4Vb4/c3hJQlkAumIhU6zY2IW
6F8EFMQ9CE2t4w0gsC0EtJAYJnaF1BAaFwKMdEV3eBMN1XB9GYO9E1x7rrDzD7HZbW6CSQlyptCq
BI6U6RkYOv0la9uOMSPfyOuAJa7/iCoQ7F8AVMnJHCg67V4ru4+MeYg9pT7rJlWdTqop9qavAW/8
/WigIE0cUcaNLJ34dfHVAMM6XYdvPVP7CxMKGIKYIcBoJGGBTd2i6z3bNQjssb6Vmt0PmulTyJPj
2XCSrEJ5tcOMUWBWw4NejP06DfTyawzKzoVw5sA1ZEwQ2JF09FBJYKgI6snv6ucfSwJom2Jsgm3t
kkrZioDzE+vHyZtFv0Hy6eCfmrNmg6nBIuwtaNLiE/LzHmoPCPsQwXPp53xoSFPIJGUVl/7L+aGp
G/SuwpolC+CLsCUFof7HqI72sjtucVU0IRxYz3bUoBkjhxBgEQGLu5WrLD0UDOp0/VU90rEZ7CSD
1558O++jz0NOX4dcYei5121vpkBMxcDPKcZnuS2NYZDU0Rt9uLVGkDaE6rhvIsaaUevHVv8QIlmN
2/IrG5dUkIJ2V3eiwS3/KjAFcCslMjuHVnKll6C365v0x3S9G8CX0k4LmGjNu2IqyTZ7I2S5iAr2
rvECWr8LmGRlxdtbIcBvNyKt8tMRxQfGFKZIaqI9naRm/8MggoLExD3iLnNdyRpWgzzoIkzwjAfR
umOzFAzM8i9hrNP23tYgFRXKgaYj1pQ93qxk2QmDsr2nFSwX/4ZcMLBVAoStv3WeUMAJtfrPQrGf
aVXaeX8fB/DGzW0T04eW35aAaNQGIFEgEYtg91dGlVur4zoY6RZwrXAhmkTdZEJ9yoRnYJACwwBd
O8BaqljHRvJqSu/Rj+QmECdTBoYoF5xLs9k3AI+nO91AOs5aLT83ZNmjyLc/4pF2DCtvln2QxsDn
fQ5L2KPAYxuu8dqvEgIRHe1LxkutPDn65VY6vEKWKtcuexBhVRyrAQ14l01RBC2mXSn9ujG6nLSu
pRUqtYKmu2VCPvQlCGAxEoddM1zw35f/CWkqu9HFhF9DLRglkBtPQY1cE3B9hHFKNXbVZrahUBfR
5j+B3H/IGq/6ORD44/xNpspiRC3x91ZNAAOlfXQ6r8uFgdOwvegLv5UdSVA/D2JmwTFTu+jZFas0
qOSLDfBoRNMFzrsJ6obHGzgewugvLZ8O9FMGlo3l+zUcERkGrJC18C51r82aO1/9aK18Yl538mD7
J1liUoOeRRxrcod00vwYUu2OIUn9OMGRQyrEgxb48Bp4hwdOe7lufz+n0IhSdLNe9aHZjaqxKbxs
r7CN0hnQu0VWPF94WRodD57X9+MO4cAtPcRPN/xMCOS7gLyqudIt71yz2zbllHp1K0HLYDDl7ydz
XkCk0pnCowjVmPlIUJwX1D4lh0TbQRfWZB8h+c075FNy1v8O7LbTv7zW3/MyeX4sBSsbbMWLjURM
zs8MCmSZrRui4pbuUX+NLux+8R+wbKvFmet0VzxcexxF7Y+BldajZ1u3Jq//ZzfeAwumSGoeIvVR
wMTgfAgB5MrbgOBf+vLYaeUAd/iDHxRKWz19FKEVVvf9jDeH6fXSw3KFFrvCXBPxRBoQp8FEkWlP
4I31yexAkF7U8ihbnHfFuLBOPVn0ia7nfy1IX2jsR/sgHuwq/vWZIEmih3VZ4tABEAnYx218VwCx
OrLXRs/Ir57nmvPDcqoGt/8r8LdWDU8WMS260V6iTlAqcm+7MrzHAboOdDyLSczM8kgQmppxsoh7
p0UgYVZD0HB8NLG1PCoUqoriWuAvImRoSwGmWbVf4kD0Fk1JtqdJb6mrEWUGKDZ+wh1rlkuaG5Xc
jS1oStvj6Zw4ayNPtj8Q+fUTTVDoz3nYE54cxiANDbVw/TZSFp6VlsVuN9xaRmIbJrMOuMTmb/UV
vjb7+/iTwKnypm7I+HmVKqmF4hkIpIczpBLa67cJeHmmBMU0mBd2e7bfHm6RI5Q8uXcQgkBOFe+i
IlRlThJEkIhRqgqrf/aw9LEHJ0PheuY3MbR3nOO6ShJ4S5JuLP+bgMccdDK6RbMe+5b9cJbxLmZP
v7M0PpMqzX4imgP1XFA6WQR3rkNDONiQZ5n1AXuytziy+NSBi7WZX/2g8zGMKrzfMp7W87iCTG3X
H8FchA1zlvuCvvtQxXa/bVvwZJc3+XeaartWAYidULryELdjsnBXPHrgroQHxM4Iwdc3d5OA5Ee+
EQ/QknFzkk4El+SYYHRM6djQO3bntXvu3UBK7YfG3yiwsf8DpCQ04Org156XMrC7BJC7MpPWtlUR
aK7prm6B+UN4StbZ/aqCPAMAukoxRKvYJzQK9ezcl6mQvvhJyCIvf+tme1heFbTx5hbIAUa6ErHQ
F9wezeNmsf7KOyLEcxa3WCAZSKibm1z+if41n8hMOr2APGZYTYbQLDu+Z+hRUFAybB2hSlQ9wBts
IRHuKf61GlIMkfS4bpHTZblsK/Lb/GjdmzZ5HgFWXiRIju7a/HgS3w8M+7inuf4/8Q+W7Fi6D3iH
2cOVHxv9CO+K9PmUC1naiTPJ8CqGL5mApv80QMZ0mQG9ioSGFJf2k11MKLEJejecYHwvYFuaeuwE
S7mKhNugnZIEHLqrDqFsrXeA8u5sfAExXe3yIJSzRcJB8Qr9pNq1IjdQK7cpeYMrxpMKtJYeGH03
qb3+nZDIYbK0Xef1nU3B3JWNnM8N9QELFkOGBmDFa9yBsmd7/NSxJr7Mdjv5oWRZmOVybk1sJvVs
8C4mwjISsk7jfYKvCZWDgLHcKc9yhB0jKN0vHGgVB+ep6M/z/BPxyT6rzdKMHJTeMBg0E3/grc2V
yD76OKWSyeQsWRBU5G8xGLO7go7tYFChGvioopHn/tb4AlbmRc6flUfLpRPsSL0X1cRSaBRRVLsH
Ri3fIve+Ju5l4sKjdibA6GDG78u5kBx1QpD07Z4U6/UlhO+/SrTmMZqgCGmIX27n/iEg6jIMD6hP
y+hEY6epSCxvBziYCRY6ksk909kAK9e6G3fcFt6ErKewB7Omk+HySgtIJTbKvDMsZeaPpg1xQVrr
z3iNr35mvaV4Rtu4x9yBNQd4eJ28LnNyIJDznY/XrT4IhICvjVJavo5mp5J7yklrWU3RAyVCAdTD
NkNMfdJMLb879r7qI0pJwyU0vlPN9U64HPnCEyQ0vzLHpIHaPyI8f/+XYqG9GVbqNQjo3uO6aNK7
JIIZ6yK2Mo5y1Mm9nrKWkKouL6D6G74XuMMvUyHJqwwbxntlceUlkkMfHVGAu5Ov5nBO4hxQBUfG
VYpXvHZYoAMnZxluS8Vg4CfrsPGmR1izPXBRAc4R45LAQsyiB2CxVSjCz0zHvngoN8mO9oKHXpEY
4yBR066PtCBPRJ8NyeosvLmTL2w76ilxIZoGuZp6RDnIOAXuwqjrC8IOFt4rPgpMSmgY0tXyKTKp
FSbt9sPOJftnruy8GaPg8G9y0LgIpS7ISJD/qgbgtRZLS+VSB6hWZsL1CucXpa6NdkpGhaPT8NTX
cRjWOcVx5cowYOZ9tn21zcWBeeWCvJ9Tl+P0XCvEvrVI0TH2yFtGSZKJJeSrNKLM2OjDpFmdxKlY
yh3EdpD74j83WIzIwT7Xr8hZeqY3Dx7I4RPLu+U3DYWPn9mb8sfwFiwd1J6JzRmwdxNettvniOF6
Wv53PyrD1XY/WLJhtGEKuOkpVkmyyo3wTCZFRRjJBmRyr+9g34pImm5wXEapARKkoEurzFLWXP+g
jOE7mghbNhu1r0MuUvdT9taD2Lq6VT0hDlUW7w00fyXiO5mQuS4FWcUrpIbuU5Ti9+aaE1kF1QYx
CilEqRrIb5nSTrNoSw6ID2u+3KHRdnmRgMWJ6A3adb6h92x5F2dMtXHQb/UOIIbYtmxYSXVtpn4m
d2NyEvBZvv0ujSTmD9P0PVIRrTYBgXg5aip6rbU+Z0aDPoxAinHmntjZHKAztzwuLHkBVz1OTeVW
bEaHpX6w3ASK7u2Aoq+GXahZBLTlQAycP9f0KARcs9PPOSEFUAWAtC7Sl3CjyTZKU9roFnUSdzS2
V0UPkDUUM3WiIYyOZcDkTuUFomPc450uRSvSgqJIGyOPkbA8ppkJsyNT29W2t631c/0IIa5k5hm7
F66vgb4yl6t2xLjgHTrQeFO+G+KyNmI2flMrJKb0y8W07Jl1ui8OD5Qx9RPBtF+ZYsq8K2K4cERl
psW8SstSTF4ZXECWQa4CnxcKHWr/FKACeq6YezwSqD/DHHAVU7/SUlUfi+6c8kaiZlK4TVdImtz3
9wxOhP9QiBjhmyTSDwDqqY5vUjucf0ltTxPwC+3CkCt9wonr7WgxvBqd5WgZiQ9GhyDsS9/BfG4/
uojL6a+h83ZjGqW7hDCeHa0sFpNJg9R2IPfSp9lhy3LN/2pKp79i681agV+GK+/P4UpQQ/2OoOvD
R/LzbIRW9ybKbVW1dzbari1QdtWhLiCL5EfCLNlcNHUmkkYkXsBi/Gx/hfLVSLlx7kMN9r8mPug5
jFtN0PuriIpua1r/c9zJY6QejLU0PlPH8s6auJGZNyxtkutcaf+ynuheflS6fDL4Zq6R0ZTd2MyB
blROSUbIK7ts5IhSzT8p1oUy+ZMPxhfx5SF00sdiDTXbf0QHdXkxprCuBc+WieV7tcZvo67/bRVD
WDnayfYYawF+oBRjwvxbagE3ZCmNndUDMnhjZg3Onwh38/qNC5THmHvIXE3BTKXTtzN1uaptgIZB
QpF7iI1OJAPFgd19aQeY3qW0GWA/9eCwgi7Os+DiFK0QfhQUWpNtSJuu7kJ+bSdPAWwNjrZ22JyX
Ce6HtQxIqs/dyRaHSPOSuJdiYiK+MjX4Y52wCKWHAjPRW6XoJBACQZuTKZLGJfkXPuItzFM+9Gz7
E9rAC7j1UtekPLWhLz7diDhBCLh+ZF6xlhBoEFwod7Ga+8rPmT3H3oykBkw38lt4H565VAziJrpI
cuYOcx9URbzb0ByIjl/L7DkeOSVet9uTvTs5YMBHdLLOtlCZZf2vXsxAxbZVeD+7bzUvOJpMvQkN
dd4eh1rbjWgi6tcth99MlzAtHYFG6jS6Cq5dbjiAs6izaRasmALRxvcmlVyCmCbSy3Zklydytsw3
WKiqgx0SxttGGUebejfiEqLW0bWw/n/QD0vJftYLEljMwh70vwGOPV8ZQgrB4dyq9KWiHVb0w03O
trtwZKSCsALDWd3mARbajO0wXGfznUVAWxEz+FI6Pwtw8k4IWrbgQtAfIxZgDYxUoxVyF/jfm/xP
iwZ6rmYUIdLs0BIXmtEJTzU7O56D3jbKzuMLwrHuxedwRpC7pmA13W+k7P2pICVEUNDiW5QG6kJi
DYOegpmrsvzCz1DwB4lKHMZFOLSfITI6MSSN4ps5mwSsjhivOJ98bI57zN74chyHyfez39ul0vTy
x58Iwj6Y4O1EzyH7mZvJoBejcAnd/HMGFeCl4fl4yt52ZyjEg1VpeVIKYibDXgZneJ+NeudNKO/w
qnT21o5o1dCHymOC633FayLIjbyEsbtkMAMJqYKNRq0kO7zEu0Xd6MQC412M1GN/fdoiRCQxX/I0
mHLnJLFEnBKD4MvzsZG/IZm6wkuhOHDWxbmGf+BfkpsgA4Bs2/ma+0b0IowJhkaN7/YspCts+EHT
ViYM18hdSq4dQENeE2dnkH5xi0LB5lkAHfvuz2YtH5lX7ddqPKK1URVak7hr0cl0UhZzjXe/CzUE
RphwX183adWpzaVphdQ0OSxr3Bl8coUG02QOtyxx9IKNCiyNPjoXOhT+aJKH+t9sZ6hw2T3BjV6l
ygs/R0BhaULP5cC6fKY5OV6HQTVS9YlOGi46CUrutbAZJhL3f36E2OLEitXBrEy50tUFyWnNdI2j
OE/UQuhWpRJvHxlhMzH6uaDjNO1lGvg2BOuSYylnX+Lg+8WZ0Gi8QBF6gy3YOB1c4acmOhnOjC7t
swNuJnArUaNg9VHjMf/Lm7/Xo9I13N18EhXrtdO4Ll0QUDeWFM/XN/BwgVcaYdD6rOnoZpo5m6NL
4Egv6mJOiXAP4aRKlEG3K8nPiL+sYmpx3PxR8bssx8+fPQvDcTpHFHIz2UTkXLAiIMB7IFA1b6AP
A4BlLAdDq95YI2oo7FiC740TmrtyaDGIS9An7r39By/WsXc8JLT0mAIE0KXcJN//fbnUNst/Qhrw
vbBwMKvA5iCbNslmfSmGcro98T0f3z9V5TTaKdFWnCn40wwC55ujU19UUU3nzrAbAXWRwoG3RYyh
pMd2Xtqcm6DwMYAisy2rpZO4TOf/0qVtB3qQuegdjf6gSE78cNlQaSUOLUni9P9UgPhT3WfQqqKH
ueCcq6AEeYeFtXAyRNfY1SvUL6k5iKY5YeDrzowSr7w+A74lG8PupbPuClwccHjAVBm7vCYC6Qri
iCtTz4XP2Xg7+zfGldlQu5fW8bwBtfpC+c7F+QEC1GZ2mNSVQrw6PQslKeax0mdUN4k0uSDKOuKx
12ZsITJAISpUHwZDxaaFzfpnwJDuluf60axQrPecel0SG3llSAunVMhCKCj3ndXstTKRGDZsvy6P
0Gi21xFAz/fJzfuZfWQcLVYPg3tMbmJgoJlVOiwjBKQ6upymHNCyZZE2nYCUrSfXtYQx4uCMPU4Y
sawFuoYQPUBPn9NvedJWBIq/oXdEk/OJc8A7e/Iz0Kwm291TGLPk/wOeA9cZOF3+BNyPcIfe3L21
Xl4yqDo/AJ08FuHGbZ2aTBNqRLEoCSW3MmR3IYKVOm1j/5Z7R213pSkjEqbUiuZ5hKncJpTqQ/11
BZFQS4XXWZ4FZflUtwaXD3eDV0i4jPShVutz6ysGy8h9ODjSd9u958K5wwa8PtujoivLh0C6oS7S
C3mBwxdm/fmVeXLgOYTeG42ZdbHIJtM2kIRWlyAZHqngIfWzW55ph1NxMUMPSQxXCQIAwOHPe2ZQ
53zO1ncmhYaGb8IwAa9u4b4YsowrvwqkiA0BKOiS5/EPNHYicRYC8MtYhA1uN7BIC0FfjXZDPnZE
08ITMWMXWDmBe849474KhbMyE3irbO4dpqkKmKpxnFk+6oSi4RKQgyY4Cki6BeiAUxNLczXw2XyU
GwWQadouMk1p2KNR/DMVn8a/hRbkRDsVKHH1MWn450jPd0FVX72IemSEkDsHmqdasge/9jNCfMN2
gMYJNBnmXeSYjWXPMXe5EpkuM614DwkJUm4oeMdaEUbdmrgMd+Dyai+AYPsXP3hgbQYZDEHbztgk
R/5G7qhVmGdgzsbHUvxrsIGaXxr8uN3y5WcK3GhjJc/GiMTmVwUM205lqIYcUVm8ynoLb4b0JTAb
j+p00e/jll2dli46XbqmBRP0XnH4Ep2WhbBbFF7s8ib6smJkaSOO5Uh8rEMSZM/2OTESB5EKWCUS
SPM5bppU90EI09lyMljIqlu0J1SetU2SjW2KTUNaajoCX2W7CGfOgTgEqtrxjdb2mxHHky7LJXZA
nfEDQYAJdQ988wooulI50xYd8vtlb/yVvaH5i4490yZSkG3+sbrP3Fv3GomFqOqTyxipNiCScQ0g
lHDBPdt/DGPdcA55wwDFVXjTMqiACpBi+gTcf4GbmmXj+aNyP54OuD7aybtZ/7FTEXcrc0mbSeXh
sWbRLjEFd5CtVrX0a1p5NBRqXov7KAAN8PCVwCfV/LqCIdvLd3QvoAFClyFXERCt7+vCm8jcllUh
TTPhV7TRxZWqFMvA3oju7fOGrWnZt45Y8aFXmvsExjdcmXRYc1vi0HDmqpO4GXt63iL6RjrG+Nxi
rQUQMJWP3e964oJlFnQXKLnJ4NhlddarsJFmVj2NJYo/2APksO2KLYSV2rV3gybgiRB+w9s3XVrq
kvaPrCp0r41m9PD1dO48eKvPaoOMl4NRX4lvdPWFRtLCrEOu0Fa4X9Qb5baxJH032rpi7NyC55fK
1tTr1O3xogjdkheidJR2xIv/XCIcxVA0RPGV1IKrdVVxrXfVVWBoS7LYecn1Sb/qsm36TWsjQBfB
99Tqj0N7br2kapndUrlnVhs79Svc88tmfNcMOoKj4MBd7c0ekvMrrjYHGPPYnLp+Iu15bQMgGoDR
gKKtaOmWs81UmyZRW3VFvC/UQaMaPeYkgXHfkhtkImCUfwxvq0thfT9MA8Jm1/OGB8YJmxLJvZJg
UVClPnfKSv8qY7zu0SL8Q+fpe2+Bkfcug323rDNXZjA2IJf64GKNYYJmW257mUz41x+JHXJiqVAQ
L/0w3zqgVAKQnz6JLSRDb+5Ia+tMesJjQuBlAmUlHzQe0JT0N1B6ZcgVSJjRAWm25cUPpdD3shdf
yaUmegsbdQasnJrh/O42qSRSZNffeFPHZcKwaKvwqBKf3NUlJOu7Qrc1vXAKbdLauBOfG6GRAZbe
U2KbM6tiP0aenRcaRrKTmnNpK4ikc2S3kKiGvg1Jtn9G9hrhD9Aq7M/bi07HiFsu5jef29UEYCHl
oBdVzfJGGUnBtcipTKmFNwqTvUqtltLTJeIpXfyPBno+d0hiloW2ftcQ/DTsBExnN0fBuoveZ/F4
DybPhCeIDr1Nuqa/DyvXwV8yjbl0JYjqlq3JBFKoQmggNGYZ+DjpAzp2UTKclwCXfTsVGpNEj/Bv
dbqh/6qpUXgIKN3Bgn7peXZjP94pp7WeudIPZ2dM7adf9597JyrogfzWUKwspRDPg3/96Fr7flrH
36/iV3QPhxZePPYxjG62a0umIfaEbsZDva8mqFbJCLd8bs2QH9qOlC8sZFWoF7wzRnUbNqBqKdEG
MsGBhhiRJEgxiq0dMNgMQiBG7VPLJ/MYmZHT717jSAmy1DPBy4wYv50DJ+JLomTx0MOoXi5RqUK/
8IgYXW85lwttCB116KiZQ7gCzwWGuR4g167x+A7cThyfHaaopX1Nb8iMYRfFqLJrmvmdllCHSI/f
6cArShSLPqrBsa+x21Kc1ATm5whwCBXlrDu7ZYLsQ3/364asM5UVr7aC7oPsw18hdKM1zZTiT9O5
0SIONhcYiudUpBmq0AGFpKbxfrFNwxOWtkWu1O79wvE3QqcJH6cL7WkVuIGkNfRM7e3JuQ8g199h
5NtjgmQOd75s8AzpRxT1P2JyXTTc4+zy9e+Q5w65/sIsY92Wp/BQTE0X04M+iTpgXKGtKJwDV3PZ
IfPNlLApnYsvsGh5mqx6FIrRIYQgqgCrdoZM/S1H5rixRACfMQVndCfO6sNGCX9SeQGQ8FwxOuqm
dEc8gjlK1p9fJ8LA/2jasPFh2yGz0naOzgaTZDAOIxb5oWIYg7ukIBD4yFaZIQ0x9R1AnvH4h8ku
9+jBSsA7ju3LtEwV2Am/XKIrXvI0h7H3iZaso8aPDIzTk3mXud7GZyeBgt9lQfnKVmQKVxzOxu0m
mnoioSb91FsxkqDbKRTj4UAOhddkNSI9iv16VCMeYsRwagqGmuEBHWLLFS1/ViiUTLYAnPwuvmqk
yfomj3dQMTBbFmlJu5BRLrO+C8/jbhZPFXeDy81u1pWJ8FAARor2KLo22RdsjthnuIfnUTbdi+KK
pBL8yrW8kOL+9toTqVNI9+LqxaEGQBPadcYV5KK7Q5455cTbijPO1CL3mFWIK32DDQ4msvEngDv3
9tpo4RbJnlt/G8iOBlULrHgYHR+CaZMQv6qyDrlMQChF3Zr+Hjloyv9T2BaYDCgugxl9tmm2K7/r
S8sfjzsXhjbOJ7ajnEi+MU05nqPvloj/c/6yb0YbvT7crpWouhu0HjwjkOw7vTKexNqxFuCAroJ5
QCf8TcrRHpRUJBUelDCwfk85Ja4zU6QIKirehS3NXAE+Ng66GKdrRfcOHn5ElsnpeYGxleZc8Llz
IWJyDaUW5j3u2ZbKw6sDs6ryb+ypc63nk+k3RLLjdb6A34ruFUJBQoSxVLSyCrSKNnYlmvX7jlNy
udmwIFUeH/K9o7u/4xKK6aXrYMm4DEJwxLHu07u6ju1y34ovf5SiQLSC/upRn1BXy+fUjJ+Ebu/h
jodFlZvPJOCTG054a1d5ssl5VAp/EeqzQTnOhuP6oXEdSf09/z29v4hiB8mrvXJkNMHousk4EIYy
pO32sTZLkhur7jfLUbmPER5e4R2DxaMFNBVO3KRh8TH/MP5tAw7t8Wi13+9jZKbqMD0GivJ7oqTs
gyfO39Ra0x0+/IxjsG1+S6PBIFYdCeYNgGBwWaKffWxAH4libXLqWFZ0uVbPOFJnAsGqEqqsravR
IEwvmTD57l1Xrf+4WtS9kqxWnVyclwOysRg53OfC3Joa83LGYjCTyxvKE2qbWjaRgFxd7wcCId/M
yrvAr8UEqaSsvDqyjgtav1NmeiwOfmfq1L45CH+ZGzVgJuApmua7mTqlSZ9sXBfpEtqR2YmB6h68
kSMvXyBPxV6h9Tk4GBP2pM79JC/FnSuNeFfKdZGOa6VksBhOmpJ9cwELzXX0P6Md8SogHgEii7dB
WWTSZAHWqc+GwnbztbeoOVC/DncTOH+dhvw0xm6/itTgDEd1B/ybUhGqFoExDTvGfT9S/urbhoq9
G8x5mbDFQs4sMEpi/RTCSuO8gNkA0voWKFp2SWOfrWdUBGjkypjHUglaspL04C+Y4FqfjZInoL9N
lZmnsfUuX98BSy2KlpOFY8I/v2UtlaHwfABrIxE3ltrvMugLTgCoeIz+mkLE4Grf4NZQiK/FGglr
XtK1oISa3yuxZaucLvABWiaE0hpMdxLK7dsTnNZ/TPRQT6FBUrdj2wW9Inkmh/nkKQCCkh4tmk4h
fk9sigRRx8bMSbp2b8KnZKiwj15/OHcHilIKK3bGP2MQMrhfWVliaX5JgbZ5DQYeKOk8b0MU3ho5
/aa4zKo1h7O1wBQVi0uFC6hstZv3a0A0dCg99uAcXEDjQkT2vL+z0WkrOEUnSE+bGfk636kHe/hx
b2/Khlfq8h6xnvYY+y0wgtoDfCM1LIjOhIMHy+OyhOh+sqb+PF56pGJiq6k3AolHHQ7eLJTeMhD5
ulDkdc393lQqwP1iNXHzC5mpmtRmq1uD101p1AKPXWNrEBKelx9C2SfIO84Mqflg8UvxVBxI+s1c
GYqIiWQZRXA6hLw02TydLOM5iavk8YLh8mrEyuqm2P9xWZNApVHikU/2AS9PfVqAJ7irkvd8rCzm
JTJY5WplpAoqkFDyI1FcQjmnZ9Um0K2s8sUZMwuKxklp13YnFJnLQ85WAUNtW81s9Ww+FhpRkCOq
cT6GziWGV1IhY5w3cF+1YOcd3ndnkvMFC2YZW4UV0lawq8ZlSRfkUF7/fSlYjbOepGcu2tKW2ClN
TnlDbONE8wU5M6B0BNn42r6OqDAW4N/3CGmjT/+RzqIccMTG7tyJPObPKUd6pwenHfYuY8xPqOd9
g16DFbEsXaViYpMilpjKb7RfRkn1kb1o5XCSa1O8YC9Hp6Jm+gx5UzfS1zZDF+XN2qhFGV6aL/Uz
58IX2y5yceMELByqgVGWvHdcMh8KmDPVOi8PbYGOcyvD+NsPO5B78eHd1cOKBH6BsJjtHDobRCjA
Aue0oZ8SRAIheQU2Ih7hfrObv3+IyqTPW4aIC1DfYLvd/9aiMnZ5K4UamcIbRevHldzZdLhdPpt/
RDnygnq6paPQmBBbiBB2fNkE0SELy/uTbIUV3Ew+CX4b0Fgiwl4I8NgywIOhZkd4WJ079cQJakdX
yVG0+L/ozzyjUeBUSItRfZTOZG6mD+wIAboPSX9DiO38QhJ8AQu8VAN9jfGFAYCycl8RjD22hfrB
++SO6KqKsBN5op8RpkRbW0JSyjpLeks0Yumqwql08eAMQzm1vPmrs3uLJc74yWFaR0IPafmBp4ZO
NtiC5PCyvAgLy+ictP4m+cA2gRnqSyRgfYP/Vg87UzWiXfArqKTrer1c6mSU0NKTEWHUCWQNHjFu
azWKYqN6shiCzi+1wrbzYKATcYXKfGgJ9VIGKQ46YXWQySjPeVdk8dZPL9pAfqxifo0QPP1EbGeB
uewXtuNd6cBMQF9VxyUTLwBiaFC0MgcILNsZCq0HLfCLj12lJg+9URNXPmeKwuOS6Wu9po5uPJg/
80WSQRMa1RN9Jg6qrlIbhS62JHIOaqZU3PtRg8ZmF9y6abT7GcHtB7F3GZ0dlrtOqej6uBx1H/SE
TkZ4aa8SeVl1gUiRTHEVWa/16g8mAHI9ecTmVO2j1Lm+WZqrKHw0dMSCvMEBjGkTGEYrUtE40zwu
TxSRgBYyX0mARt+nSoGPWGiXribF/wrlQDhOXRKGl8krhNZ3GU9YjRdWHR+d6WHJQS2V/lNRlVR5
EoOXLPrMHMHBnIqUEPy2i9rdG/LknjrZEnodhhtcRosZVzdSodWGcxTzVWN/2uxL/Y4BT4RgH9M9
T2nsvrvMLA39/P/bIDPK/0NmghXs4FntlNdYQo8jURmAn/6KOtFW+O96zLfFiGFOjuMKfYpDyIKH
SdEXl3PQ6oNRgJJ7GvmhUjDZB2+lsq+PNcvNxUu7BmHk5ORXsCKfroV1rycr8ovE3iyqniZNmNDa
RkiEpw9taQo18nSKPvRngskqejrbAClVSlAUk4QwboqmyNyfYaq5sqjNpah7NlXokBOUiCYRTLBe
MVWnHi2efe5SPssSd6sSqYkUnbbkyj2xsJURvQ4hQFFhTj91LaikVJ5kHIxGpxLstMuUFdLmUCka
sLo79EK0wTGVGQdA/lDUTxZck8yjjxecevb0qTngtA7qXzfDF8PyYTgBkIJ7dZimVHYXSVEb4mem
5T7b98A5nMg67UzZJOdZtWV0dHWW2w4Y7VKBI0Q+QU9v7H2ojjp/VJtPEO/DKFNmN65QljTioCa6
WUjUYe31Z4BRggrSN7C6HosXWQGwpWVf3Xr6Oi6eSHpAwg0XwvY9At3qSxH7dDTOaQpO8q1VMxPc
SSOUDrNxCTQZqdrUIA5JXx+xCy4nrGhzFuuQgt1nJndIbB5HV0d0+AsXSIRPW3u9Fv8558Jjwwue
ypcW57N54eD5Rd0CWizKhRJOKp9VkkOX8ngGn9FtdzRp97g6rObH0Gh0HHElLELn6adjyONPEB5v
FkBWFWjmYjt08sOUiBZKVEJqlwL6sO+Gv/SEdIGrMqnrLXVL25J6AYqKJuqwnSXkbnpgLdRA66Fh
dlDi5G7fiKhrEgxGCQrOQFUxy4HOkY6CxAyonDzu5SoiqhUSbqUH7U5c6FBezennZAo2T/4lvl6z
mbQNfFTkEpFwqV2EggiHz46RnYjtDFhFdsmaydwaPhSSLZJxsAYMg0Cn2m603RhKNgqrIRt9bjfi
CYK8KCGEHxp6koqwrkyjXfqUXQFrxTqZ+v84LDS++GJPps1BKyVLLXP4vcgxIjaeXppZJ/7l9q02
ChW+60AoL6nmcZzSvDL25H7bnx+82SfHAvZ5zsABjj2IjfTZxs8ysseOvy7ko4Nm2JatzB/COqLZ
6Zb/A6HgehLPDbTxbSDUeYbXxxNqP2ahLGNzO/4C4l1Q9mkH2Vok3ve6GSB3Yn7eKO2lKDdeSasr
ZWjwO4RY4ik099rSqUiwewr2HfELAGprI1gErXoWreTkO7IFLtzUE321u/epR15aGwJpjIDnbt3T
or+j20h8mGE+Ydo23/6XVYFejNVgEMdgdimStwHlltyUIiZUOBjyY6wkgXdizvFwISj54I65M4t7
5Z+a+eL+Ro4oIaV2f9pquqysYz2XD1CPAGDLIU8pJhFEghVTh4TX0HP7EyDXXWZg4KNbmP2D4rEU
sXcRg6pGuRNBKvcwyJurRuvo1S7f5M6s9fYe9MzXkm3XqTT8P2uryyMDLCL/Qayu33MIrz4ophXC
i+k4anD2vSgHqJ9zglBuJcKs0/6d944jFE4FPyeq9vDImzxqXYecsQXBhYBVotZ6DTn5L8nTacBB
CppZPpex2b6HQZfB3JuhZtTTQturmVmpyxSpwXu+Rs0hJEL7S8J4d6ohXPmlDJfTqoP0FKrHkVA4
Gz0sRuKb34etHJlHvMJeJbXgCeyeDpON4obotXf1Ec4pJD3/CaiQv8ghdD/OD6rdF92OSKFeiPYl
3ppOuCL7dLXWxZjP6OpCgkPEA5OdNgotUAk+m8ixeIhpeSk9SnWLv40lzjdrSFDss0k57F7Yhz4J
oXSQFta8sndJp6WQbueh4j6aiBXDQkfeR+9+ahy8diWx07cRtOAwKn34Ya9G95HjNWKJo8DTZo79
bzPoEWQ6NVRx6o3p/bkA/oTcLIWXUKWlOAdDEeC8Obw8+5fWZlgr08sKGI1CkBrAAAgQWvJprPZu
3YcAvA848riNSMs6MmxqX1O2UzoMspPt2eQOmj3vrLoWE0fiT+HvKdkt4bUpmFOJQAq/3+ydsm5H
FAJaetyBLIoS/2QBoejS4VyD6Lqd/64AQMzkHtXpHEGAoS2fTbdChwXm0u5jXgL+Xm63uw2HBk4w
SrDwzC9I8c41nIPWbs4MTkQSygY9felgH5TdOGlRmn8Pny32YObAbtrzaTjlZV8Qo98eRrdDSeB9
3t/oqzYCQkVXnBuDiETWebmdC6L/KlHvXinO44xoh9vZm/n8ddhnfp9zKS8Y9p1/GssEk4aaj1wi
JNRt5iMRRQaoM5CvrL3nbYvdHNirO+iOfmdSlfe9pRsPs1zfBlPj9PfSHjPdGrHaRfSA01XWJZFi
tS7FA52Bwqp+YJK58lO1ekAc5Uzk/8TwHYy+ijR9/o35MoEGe75PIKjtOqGOuqJWlXcTN8yG86IU
udeVKW8cG624xfaLVxe3rU1t9oFAM968fY+IQjmYDDrQWbnrWiQF0KtJVFLYSfNQn2V7uRrqgj6/
UB3rVkiT3YMkCGO8o2ZMTp+vi2IrIn7y73OIA423rXMb3sMdmvE/3KjXQ6SMaFTpwkgI15/iYTNr
cWvFmaoCjht/UUiugXB+7JaU20dAOvPOIGEwu1FHWU54+37EYEt4EBq2Bbx3P3gTcClYTmOjoz83
8ULl07ikchne64h8xfPI9uNYPm6/93sRxfafrDEMEJVYe7auHKg4gimsSobu23tbsuYRa4UvCWko
OIvOaO3OqZmWWQeFSDRWJclE2bvdzR9fhOxnwiSLYx5mckh34W1dstRNiPRnl0IetrWBR+z8Q2q6
xSbNfICXnNZXu/4iW5fkqxU4WULVkZ9vTMqypxvMtDqdLEnjn+vQRlwOGBrsdegnM05JtjHEHYkM
iDGtIS1RvhR6cXVrmsyTqh8Asy7GLvcA5nZy7lUTAerILvhZa1tqFEfHM8G7+GHXpSA8sJiXYPcn
waJpg+nhmhMYQkhPjQkkFomYSe0cBc9HOdqP7cm7yFLxAEvtii0bStKoQ8yq6BgOgvf6+TxUE443
Kdz2999xBci/iQkJsi+fVtMpYP/JUIoC67P14wRQlEQNGeJb1UJ7jH6oC7wm8uR8r9cygWysasvT
SxF4b4Kk4F5D3wl1BfmWaKZQ0ZGFZmzeUX6RjtiJ1L7S81nKw+172CenZn+d3Pia3lFWgI16Qbqn
MBvYf6pL3EmKygVhpBgl++ozZqe03TL/tVbu41D4u5XS8LOjp79YwxcDpYy3FMKQ14TB2HC/fj1w
2tu2uYxCpfmhKYwws5sFAKn3XLPnPCiR2nZR2g2uDP+gHP1V5iLg6B3DINjGqkLj64lbLfSrt3Y0
iXzgN4xEWXjbvkL8o2RY7+WUZ+SInFCA3JBfrzUwE68HW7siolaHaZlHsXCGLHX7DU4rdUpQ8IyB
7Ga1PDfPmS7To5vvlRy0PoWUXMnqYkMf4gg/pn5OFO+QsOOvEuwnTcduTUopIWn/A4wh9Po4At5x
rku7Tox0iS5OaGgRkHkwJvRZcaQNJ9k0bUzMWQYGNN1/5i1nnzNOoGVHTpbZisnvTNEC8EDHI76s
tmweiFzOagwB2y/+srMWYhtdSNPd3Hu5r7p2plRJSBsTI4tpGUfdsbtjHJWD6amH+TgtiQW+7Ghv
RGI05QEnlZZs39Ftr8H5fQmn5dxeK9TFAucM/Asu76r7vXiwoZqy5Xhur20xLmyTuVr+MC4IsS9I
xsjCQJeiNsNvxS9zEQQ71nTUCPJKGf7SCNseSHRAiwofgvsBnd1ms9MPqQK9n2l/s/LMyNHd5pnr
wj5YRse/UmSySQo9b98SRpwqFUx1KrU/m3IMLlxUL2hptsqsxVBTESLMPrnUM0HfqscAhJbbM3vT
15w9PamlRZ0sXgT0lHS9hVDfujkupexLwnirB6qq1gdlLfPSGvbCXkOLnvF7VhdLIGg4R+UvQDag
yGQ86vh0ROkgdEKEiRFCeRyMMVOlBoYGumBA6Td3RP6YVS39JaF6KN8aoOk9hkxGH66qr0vIciMK
Zq4ZmgU54Y1T2+go2rNqgrqNWlhMDiUR+8BJg8MWEygA8gjM9hhTnMAGMiKVC7H2K/N4y3wFqJvi
+aX66Ehf+GY753YNIqkKLUp2Z3s//V0uikwycJqfvFAw5JR40H5daW1FxFb/hRQ+W7hmGWHWSjO5
P08z2RLGSl4HYVH6T65iOskJSrsu9Zh1Zng3hQ2H/dAgknISiaGVg7IycQidwuONevuIA/tU+Xfw
3mqtHWH0oBSfX73mT2KBMTzXrvQ5eyWMJ0jkUCGlVJOyOukPUTYn6qs5QePuMtVp9ZhAqmIgPjww
aZEQK3lWirPPT9aUNPsACV0YA62v1w9mLdeg3fbn14zg4+sYG/ha66wYKjWVITcsvyskn7jKNcKA
RAs18Lddg3Kke9NsfG9d0GXCCkq2nhdeIw7GUk9RInkbmdTsZ8K5xfkXLvztVeR+o7+DPuc+j5o9
JqYAa3JM1XZm4ttWy+DsWqnlBgazxgSuNjshw590eQ8B8VzNT1v7oszB2jN2p9rF+T3XNsfStHln
OtmKcUFTiq8PjyOgtkRrmOBsWTjJcUW4ul82ZiC0rMr0UNyTMpVZL0neGrMIBLrHR0yBFq8QgEYR
pipV9qZlVDCT9PbmUY/0zqN9jtuNlMR5LOalJjBFBSXwYJq+4An+ZFEqpC16s2TmAWHbyprBKXE4
5/zX1R24Pex70RjIb+EeYYBdAyTZHh6oxWQABh8BBbg1pNnQbxbD1VN6sqAqZFzse4D5f5bX5P3s
r4BILEUhTO+MFAO65TDkI+CKC7rB37BSkRVQAK/ikGwAS+K7kjkfW3rpZLEqTiu/qK+QX9IzLqIi
iTaUblqntjghPMPb9bKwGxx/lPBEM6Tmc+06KdKda+Ru9NQAZ/8ohDoQX8TRmERfxzII6gv2bcu9
lYBy8jBX0Lp9TgqHHDDyc/AU9j5Y+4q1msLiJfxgSd13UPIQvptlM245VVhM3XwdF5cnR4KlUHrv
AXGvx6ElxBj+o98APWrdFa0iyr3QlCWLa+UdzMt0zdCzconGaihiR8SzK+Jhx5a0WUTft0fZwaGn
zdy9UmzyMKR3JeRGLTIAGh+ZoyImtwFSIwEuog9IY9VDF8cZj5xOe2TnPiRvdJbHcB7fadXgRt76
F30Zg6O64W9qv2SLQqCYOWeb9iadYNshe1jBp8lky3HECr3mqyZ0gzga7+E11AwqhESAfXNDexWm
6zZHhrmHmBte7z63+82lmL7vl784ZukGtORkpdTsTwX/GQoqqusmThlkDrK7w76Q+RnSZpfVAiqT
+ntTEY728BmfcskbnoO//XNOcPgXi6aDJpPTa9jIzAcGbCDugi2xx9vslf8EKkyqz7w2wcsg3Tcb
YplrjCnDIIjy4i8d6O+PYbynXZ+MWft8mWtvYRzYmjTMy8vDDSdRXk+zEskbYr0CNHMoIvhCMxpe
vTZa3yojT/lpVlsY/lCY/kYVi5f54OkM2dkrwDw6zCdLpj9ifZ9vePSIx0yEpzu2akuQIaIWHnn5
QpIxWQcCWLwtDzRoESFYk0uiIbM1OH+Fg2QMBj5BUlvcIStehIiBY9IJT2fJobcwVt5jgg/zDmDn
mjlItNlfGjbKW9rqSOamkjwLG78nLkuZuAFMrgbmB2l+g60uCxZAxN4jiskmYx+9u40ZStK914hF
cUedletyTuNsXsTbm7T66gnbdzm69UZZaWucOeBN+1APBDSdJrBbC/vYO0ovNqwGjOF/+AFLf3j3
/nYws/H9rEe989K81VTWJnDHo7NFCHroezvrGV7MMmUKaKagv1hJCNSHpNHJC6XIfAyIf+/TYljG
wkW51XZyj5cNbBidbYKK8DCewIol3VWu9l/tQTKSjpkNKKOA7bMnoFSWO7UZSmN+2nRTsged81XQ
gDYRmBNNY99liWZimUD8Dk5aDlNrQZQmRFVGjDDcc7i59UQ9ZEK/XdgtHYYG+jYvuIafFa8lbbLR
PHsWPj3y2r4XeQQWZQn7EJRuhC1WOnx7tJhIDZyiV3XZ/z7D4u6Gm2bC4x9iX0T6sahOyy44BrU7
doESu+xElY84KHNV1fFgbQoXIJymxQ5Xu/2YWioiLkcfJ/7Ii5l5tkfI1o56X2QURfFQSmIVp545
CqgrM/npcvWpZvTGHAhQdd1lKUKZPX2Kl6QQdhcJiw9gXFpaX5Arb8BKIuZAgVMAeH5nNJSEa61r
/imbroS37nc+4wxrLgy8vJSQHc1oN1RuojvTT8iXsjFM/i+YctjWrZOs6PRfXyW9QZy4ppzPaLeP
CYzo0xZt4ilUzssuibHPOziAGR2HDv9+02HiyQ881ii+chgW06M71otUq6lvuHxtrioZ2ZJLy4ed
HcHeTaZHZX857pVEv6jHrP5AMD7C7ex5KP2DdWZ5a2huZxa0uNCveXRNiLn2KsKtBWfCkslHxEt/
L1IGnmJfsQQajjLarVM9+F0EAVQ+t21gum647SfBtXUIgoEjqvndGHa29AzZtPJnKsG411oyS8yr
q73HLBkc1ZKwuChcIzfegSdPa9CjnHbVrpF9mxymoeAy/if8bNCM9q7/6Mc+vQiSzEkzI5s+SWZo
y4vy4NKmu+cwldcWAl5w5J/apBll7eXosWbWcMwrrmlza0tWN6gk0vdBxMWX6Ec37eQMKYiJWOAb
ZogBZqi1KRfbobctJslIlZcxNi0YqU9/mQKkspUZaSAMRjG6DPBNHItMmt3PjBJC4qq9/YqgOEFK
mJxekkRMtMbyJM1yodVluqSw+t8h3BuLPMhLOphHneKzRw7JlNpZwO2v+3O/RVvcL1n3uGIs1Ndv
rjxSus26MT9Pv5QsENx+GhY1gqesL1hr6w54L0pEloB71WP6ZcoDcnQMpNKqGPDP6ZbkniNtNazg
PMErIIdJC3SlNbPT2pd5cq5OgJUT1K2h9W4GRQVpgybrb0/bf8RBJxf7BT2QFEVOF/Uv1jVCZivX
eFEk8rrwvqMYdDcp5dUSLSld/doKfpWVLgcgcDZjHUqtwnMvvsV+SrpYSzpuiSRRg23X+xMRkfx7
3IJXZXgIwvC4XFPluZAq+G9Vt1KbtUUpfO2E2vY7PMFqmjjij2ky8Cnhr6NTBjntAGZJwF7wjfDm
x/KD3yYERSRhst8sf0ua7NIM2GKw3/F6WLo8HCG01V25TA17LUzJsbY6oDMehYxKAbp7vt/+aGK3
ccu7rjKCzFZ4n0VmBfeO13H5vDF4Tau4OEp6IrgVPrqAIIG5gm2O+eMwDhdvXWsQ0ELeHI1//zBS
ZeyUEfBYzHfsBjrUTPCIv1Ki0KCYSrCPaIYTfQwSp3vhMqVD4Dpyu86w/HSG1I/tP1sa+o3LEE4+
e+kDJpcSZ+NUt9/iqZUsKJNn7O5RZNfOpwxyjvJHN+av6CIGpzH/yyNFpUC1nEcPOZByYl7aQYTV
aiTwcU2O/0+hZs9vV4VJAJoAACRDjwDR6VKEvVAHg2mR/+ibEbVaES56hXxF3f1ywwf6MA/R34td
OWMaJCBTd+28g7t6kKux/w7kv8l4MEHj8tmFIoSe3bw3O+OiAJ3rWkW30MY/0uupuO1fBg/3SasD
Xp/qOOBLIv3qojxBSF/OPUcLYfb4VfKh5Yt6rGNe7nNiTjR6YsSGpA76PegQ/4+JBWI+e2Zydi/F
d80FPw0w6rxM1NGZpi4Tr8xxs1uLE8j0cuGT7zmaT/3KR/7OSP2Ccfh/WjzxrRiIU/cAHpJw+SGa
dPHKmz7J0yCKREYVIhZaIVo1kYk5LI/xaUbVcuXNb8kOL1f69ci4DV2fOpbiWB4wFOOWILq4g+5o
cpK6wUgEjGBT47Yi5RpTzwFT+p8nJsPd15fAoa5yVQE6KJnFeU8nViX3Brpy0ljja5lSLdp8frSi
IGlZSD58Ah/UR/TwdhlnNub+vGfeRO26QuO1elVvI6vyfHmnKCmLXVlRbnboMziP0+OQoboVpwGa
ENnLqK09Vwzy4SPn1GnTmmb9j8MUCKuPswgT13E3pIVIpjKPh/Ldpx2WN8QUWyC+bjV7AfHBCSy2
sHD+vqcLODB/GfDWjCibuO/jzP26ynqmiZ8vLcQ03u9v0Qrzz62wEtGhCuubxX2+kdebDsQXx7qd
BIsPLyZfPr2dG9+pp3m6XsXJjeK8ajel7ttIqSRbunfV0z7zEwFlrXLnjNnubDqlebOXPngdQA0+
UNbXbukQVHosYoEI0F2zlzHIrFKLTTbSIB+rGt/4V8B7oFptECNCNN4DOb0PskXVrg6/O02Wk6yG
PORuiQ7Ibf0DliyOIx4SxDV7yKlM2Q/z32uD2O/ZZrGv/nhQYLuKjDl4ClFP1BbQi/c9kIVymvDm
wdu2DBs1wUPrnvDrdiWcG4TRTTYHeqLfEoZvGBJ+3bQcRZLbEY2g2CUfg14OYKMPB8BSclzFpcja
mRW4vUeiCLQNyrg3ZGkuqEjm9KI7aO13XPfTQUoEs53DrF6YYdqPLP/XiavPxIfRDDziS/STqT9z
8cZ5W/bUq37Ec1R/LzzLKPH3TV0hsDAa1rwMYV8MyxmCOTiyfZ5atdCjs3KS1tmCgXQM5gTjVzUC
ktHUlt2R4bBcxKo2ROPiRagjk4EKCdcmshRadyrFo0+5fFT/CvwIP7O0cMuSW5rKEU2EUvafhuH4
4y8d7KxDv+GFjZIPOW/PAmTGYsri21lmweBdXBwH6FGWwuiOGxYwbM+g+xg8Dm8doLDBEFhskWb9
3DDkcmXqDE686Jub/jc6begdh95jY/K6lw1q+Vx6/mtKhZidj+jCZwDXB70XVpB6XPegP2R5mmO5
7k+//teWaNGn4oSzjU12axawsmyaORFfdQnyUlGKV3GT/9RZfS36a999fDHZbUd8h+rJjM6n8qqI
RF96EChDx1+Z/tAcC8yjHWzsowMaUJB7oDU14pHsy4FlAyzF7qxnUumRCxiCN+h94Gg6m6nOApe2
aBMmazHwvMOGWDvX7RvlMPaRvFFxG7T6uY2WEMA//6BB8xNOVuVIxeyozN5JWfvuYmX3wTn62A7x
e/c0v6HpVK9Jzt885qRCVSCrCmireX+BXvfXqBlaoayyhyrEEYrjHT8kCSGqV4O49zp8tgOWF7Gi
iKx1S3pnVw91hOjduixT1oMAm//nocEvMeTACpea8alDGXgWWY5ayo/MXFpxq2+JVHA90EM9ABvd
dns1LijrpTVq/+W+xtAgUvJJSfqFQtvfwNTJ4dwyLclj915NIuckLckLQZb3BtGFFWEtwRehkv0r
ZDLA+0LBiWxQZAIXFvbykIv2YUCuVBb6/qv9RufORfuRAbutw+d+A3EUfsneaLNy+822V+C2ubQm
56HsRFfiy9ZhWKHm1S40923mZyF+xgIyrI/i82tCsjf6gMgmCtPa8PJ8ZCtw1HRcD59hh/XjCb/k
Hi56xAuYJaMsLdiqxmstIeascP0hxwM0q6J9xzM7p+3tWehIOI+sZFbWUCRiDbSLxdAlenoAcd0V
H67oaO/VjGG6IwBd+iW4eSQssUAYT0Yj/kDT+V09650ZTfulSsMkRBdhAHgtJ6DUA+qxkWnTTtbi
J4XFzWE9naigJA7hpK4tr5A0REUXcljL55GOmf+i05fZSXmbB88uBKqWcMiWBM+HvjRsOFA9oIQl
Q4wCZZDIcdgnLkp9iUk0i2nhMPT1SvqTLev6qMxvKpBcbi47CCPArhBRlyJEU2p4SNVaQFd2Iq1m
Z3pHQbI0hNaf1JYOY9vQuGYix5m4GejrUwFbD+HgdUm9Wc3qFZWzGW4irmSLPlEqWPGKYdaWuNAX
Pc3uDGPqup4GQsRASNd2i0OfI1bSCFyFPqZZvWG902fRSrU3I1DAd/a8Bvf4Jxwl/lrl10Iw9wKl
cdguQa45Xd4krV6iGWhXuMJucRrk8IuIWvFPEzKPojlaidkTjYVDKb2L3+Oz9jg/FtqygGz0ho/p
AXvvVumEFlzIFfsK2lJjpemuQvQ88nB1guftoZ09dN/f/y4QgDvAt6sFDaM6Apoz3DEIN4LbZNS6
Ri0BD5m8TVXEinkiYNl0cy+HLXPxoulx0L810xhJhVe1MAkbtBwye80E35upWnYtQz5dSsSXzaui
ViU+XnT4K+cSP+bayxvLzcJYe0z0kI8OuVtvWTUOSUPuvXVSLSlQNW/93apVAHObTvFwJbaX9MX/
IcgvxFKEuVFRMDfifUHq0jBQJweB8rPgb5Jixi3M/GpJtGsIpm9/70p7fbmRZJ0Lc6VyWIjggAU7
dCA/Jzjnj/HPKqM3e621ctoBDqJbMhG6rKg9DfEBai5JeotltDFGtMkI6CdqxpAf+YBteQUlxJAa
ABDk311Oqjz1PcQnIgosH7tdpW2DH3D5iqmA6RxUaGefR8vpW/D+5TghnVM237kDFC1G7G1DhW0F
8lLD+UhtZzISZdBkni4ZnGOCQ4J4o7jPQhh+jroSosVZ3Ah3stDHa//wpmBHtMO/JXCukEtcJPOE
a5TCtXx9qdctRyLQMoLpkIQUUdxXzBAKFxMm7BF0ig4x2VJMX+7G532j6khrRNmdnQv2YUXHCIs5
JG3+Lxgv2/AVjr1Sz81nY3t13qhKPKruwzoZvngYco1lLYkpj87WrRq4k6jVlpE8EwferMnDstQ1
zO/xKqoF1qZncGXpA+27drLM1X61zfIbGjLgqlFHK+TIhDNgLI7uLSFRUPtP4W76Q5ZplwvFodki
2h9BX2/2IM3ee8zrNw+BjuPBEO5JvdH1ixmEETLq+Vy3Y/yGgQY0x8PQKWhe84XsX6Nbf7HAbUDQ
/GGA5Gou5figIESI2UEVH0xAFDeHhzA92177ineYcoR8dYen33J87GXrypcXzRvef4Q3JrBPs20/
VYQFSv9Es9QIx/GgTtWPjl0bBOdq9npNW6mM0ku4H74hx7mSfKK4/2ceC5myKOFFFfGdQiYrzEtB
m2cKWbKLUdpf7VwNyR3MwQKyr38PmvVN2I7bZovA6Lzpb0N7iAy6EcUizs8+JU+L8W420ulwEW/g
ZcyBajHX58MKUYGbsydt2VTSyqap/sGw093OgMKL9JsebbGDLr+ZLWmxglvdlcjK+5Xmzpdr08mG
8KXpaAm2r0JnjwoY6ohes8vvDB9AxTebOHWpCTzdv+lKWQvN1M/wh10GkaPkF1+q4PleXNH3LGT4
6CHTtOsjvS7cVL2B5hTE5ralCjjnIkURaxAFFFZDYzQss5dMmuLmUl5Q1ZHmAajHZ6rTHc5gFWkT
30VEY8DjNDrl/7O7uPU7DyviE8KNYgsYXyaBQrbJSyjA7dGIHwtt1rV3gDvCndXnmkkUD48a/MBV
7j3KeAjIXPZM4qM59fzlP69s7wmr+Dba4c9289PTXeXt5Ly27aObC1dWp4l2DDNmieB+bH8ZU/sI
Ki/DQuuyTyuhwazAnuvB++CAPaieJjP4nMNk3Wz+fE1nKDPnwE2KcRsAZJezE+mSl8qOamFhAFnY
uhtiGY7uLwIRwBxpUHFzK7Sj5Ev7ztd3FHgk0BZOW4GGOnSLcMFEhfx+BoQ4InolvgXqeskMKl3N
UvOwtAVm3N4u5UTvZ+LJBxjkHRkTe/AfJ3axRCwlIWTADYx0BBvy7vKUJaehmTG3V9nBq3Ye9Io7
5t/Q8u0ELSg4O+c2aWlIvTdaM2FhYW/zyUOGcTJHy098fJKsdR/Evm/qlYHNkTcN43Y2GhOcnN7r
320Rno4uaHIpGwQ9yk4wc1QDDHOkLD7mTyvr+aI9msTrAN1fmqbZL+211BsYlHZ3nFdV2SQhlR/v
H/VLr8nORxykxyhIgmc0fYJC3FCmO4dkiNBGWVQv8pnQCT7FtYxC4oNkZkjlhrD7dOXZEsZCWDg5
Xi62vG5wZLIK57lCnqChrnP9U8q0bCNMQHU/t4CKtSLdQBvxeX4zbSyoo3uDJbkfSodxSW66aIIW
lV/PhkrrZ8jJEx65T85aj2kiFEn6J7tvf+0QNqc10zdJnvn03fRAP9KVLFsRZiurMZ3iuYt3q4EB
PZ9IXQG/qx6cVRvZhkzZbg9V6sYgnOlbmXgjnEy1VOsMsauEmG15AvtAImu3H5CdV62QUZvg3aj7
tsGk8sqI9f+N9Kd9yUBC2eFQ2+Qnt/fDcrd2mQqYWWDVMZjv7G9qsfLLYRWy5sCJkxW7X9ZaNnCU
MfQm+kcnKp7j377EE9qjhKl18+WKdNDiac2usIJqa9MO7+pWp20qySPTUktAQKaV9qCo+U94je3E
F09amDibYcDHIcseH1R4GouhX0xyIjZ100IRblIKoZDpEMdcRduSFp/pGJsGYbJOtFpBohLg7YAg
xdCr2ez96v4HshaS8cVPwCnVP+E3l4P6Q8FkA3nge5pkMAM8LGc2gQnGmorJ2yPhZUB2/mTCBWpn
A+Yk/2HNtgC3Jea1HpObgJcxjhO8P4zeFOy4lDJi7ZyBeD4esESk5WNfuzEnD0LD4omUl38a9z0g
SWj1QFkeD2G+GKrs1ab5vGbW6KSKQUSqtmY8QgNfcH06nPaU15xBLzbc/CFBFKuBhuME4QfCeFhQ
nlE1RT95LoIn/j7s/QQgVOr3DMR6d5RDcfC60HGQi5Ssuh6Jsf9EWVGRuAEg9/9Qr2fuNYbCE2k0
4zdSxAa71Ml5arN4uas3vYShP6WloC0Np6ALBk7gwXIAv0Jhyw9EOwdp6Oc8J2fELp8DXE2ZKS9x
OLRgCwx9ExLlcRKXKmAcdlhr8MxLiUI0ZYi/yGTMIuAHgxSHyu3DCaB3Dbx4exNn9GEiwiau3cmh
tmiGeT1vqrEzDRMkhJD8LFqAPIrnByse8D1SUBDaE0g7+Q1k33yO1WucrXbCOZCMWOTEIZzsT+nJ
y2m7ruWGehndtw4M8v8UiggVqn9XTuOG35XGFAJBx8kTFHSdYoN4n6+oWq5/Rj373uJyktDztkp4
pFyBenI+R4jgklB60rT9Pl126avrubszbvcPg9Vw0GmLdCz/slXKrf1hRCMjcVQ/gKnFAdXf7nfl
C4mxXDBjuuvydgmBdWMAesl/4UgnD8QLeRIwT/LFLO5iU7J/yuG+olfwErHMdpJfx9nVry88Ntrx
BgYbBrDEhiiDli3P89peLppw+UvQzDUlWSONJhVMMBATnLkQe539jQ68UrBG/SdIS2xU/mlGSVXU
zk0S2FVZ/IL+/xpo+ZSsMmYQZNA1Fp/ohkCwSw30Jvv+k4jd2YnrRQAhrlcFCy2jU29jklZiMO1+
YWlFoOaQeZkhJwgpwndz6vyHKR7pUjRSqXxXqXpzylpQxZ7T/kOQkotgR3P/fHRzd1Am6RwJV7v9
aKMg161d90Vl4lAbggzhH4do4DKGlTFQGIqK38+t/BjumJLLU6vJxghUz9TPcgHsYCOOJ/kgWhb7
n3el/RLExW2T/1RWXhIC5vqKpkdHXgXRV1q4V13gvNtm/s2F6H9Q1hjsTw+W+ylcj9sG7UQA2Z6f
l9uKbIlbcOLeKDIUYKlWaNUJPAEQXT8e7dqnpJ315k9x88UUTO7V+Fys64j6QyECumaIdJY8tiXU
jARuwPlu1e1XBZA+X0STZuEZz31reSSFETd0dR/WZpQR6uctq7494PkI9HjCYZkBBATD2+LHCuGC
bZvyuEY36quK0dhtFP3DAFAK24+HIB1TsJiqf0rpDvqg9UkcRON3f5JpCt1Rgxxldnaft6pk93Oa
VKV77fk3AmnALtfjOFvknsZiTS5tESlwKBVHcmNO2XPODrnoNH4za3m19lcY1nT4MGZx5quHVq4q
eHeta6CywAgSxuMOSTStBz3lhemXxDFkMTpkHX3Ui8v7Nr5sQ+GO4ccBKivFo4pSrYfNHQq2uyhS
gHzgM0cV2NNatzGBp2qIJs6MxpETsnMRuqXTUj/zAX2FDznOJJWRl2be8C35WKiUFDJbqHTkqPQV
GF5bh0smDhyJh/dD/iZ/Ugyxinp90YlnAWrddrsiH3312IgwgPuq47l/BDpU6wvlqya/K4hqiCtz
J8MfLEjkVaqHNHVG/SP8liJays5irr9yAGKpfZEiRaFxgejfKFy+L7eYRHiCbri+7Zj5ywcOgJkP
WrY0PTkaR6e9Thn2b476TLa0p+BVn2tS2J4LwqOVhuLnL5qw08Jh7hGVlrvdpLTXvtj/vfV5Ay+m
Hw0YVb1OmOJsgDNoLqX0RGubuz69A4ZpUJQyOswiwVV2YVbHWkGGYnEdvDAmBCgc/InQYRwHHQwZ
GZI5EJLLTSQXjMFe03B8bdf4852LTtcQ00j3OhxVJnopc6Uzj3Q47pprisKy/TkyhsW3ggHnQDGl
ZNgv0XYMcRfJ1+J3vhKfGodk09lU5Nqd680YJbWC30PtLXZyMtLfNk9/CJIRt15nKcItqb5n+KtR
3eLZqqPaKPQiklZWDr/RYA2Xpm9s+Ost/nk9gEqyPYjRo75i9rbN5ebGIQIXvRYcqwPLPpY8RRWw
7uaL29oIpkV65pe828bSs7vFE7KA1m+KwTtm3sVM8dFjSTUApyxHUsXy1wRtXbrtTh2k2f/5rXaj
eHI9t2+wwKqIfy/YeMvkctwWU9bXXU/U+XTdxBwjOdMSJa0mKwmjA7aizWbOUPpJnwCl/24ZKGli
jKWJkw6ehkDdNqfDRvJKt41sqS1vZvbCdI78HTdBHdywxasMbqBv7N5/KFEBdAHLLjfVyHFtg8to
7XgyGXC2BvHymwEq+eKtXF2OzQ5BBlass6d5y1m8xYdlxgvp6WB/4fY/OhCg2eGyiZe9vYkG9JMn
pOsnR+Gstg8mcrQN+RYfpgow4+ARRoPmBIu0W9Zja3IRCUT55e+yUxFkrK/DohmK0+qLncHTieFe
zgduTNg2PyNp/PUIaTMFWyq4o9JeeOT0+DSw6mEF7EjPsggXkKeuYXnJsmYVYVAw/iwH9wH1orHD
RD9Ovwqd0tN5e/Oue5f+Sk0cKAIiSkclCHVO2ThS9IoDOGvClBpipmd+fMJVmEqduF36eLl73z6R
g6xyC9niNr9zwotxHqBfTXukfPnfhDnJSO/yyu/gS/yRH+0C9lnq9wmP//3PcR8FB5AivYFmW1PK
Fm4zx4uDkDdibwYYkcQ3GZjMWOMUL7dmQybILM5E49T5YDdAXyQHjhjD1du+9iZU6MkHmM+UTrFx
gYM6HHmOS8DO8E0ncrsJKdqBPpXyyBHahZNJ6tiygygnX4vZgBLDDJp1RIagtjEnJV1Fa98IIIW7
Kwoyfnj1WWcfjusX1cyimZAyGDOGRYHYagFPU+1+ow9GTqtYJNQsi6KuIGw1CMWv26NoZ/qNv33P
SBqDygjGBytn3tpHoCp3w2LkWixBe9Jl8wP5kKoxJxFK27ViC445sYba7QIArDa7vH8DUQfRC4kd
lBgKddK901w9BQushsud52kLFiKPivlH13CUa55YOGDrZQXJLIz00es6hYxzYVRxjiMOOtY8ke+P
g+TpCqNLiK/YmgA5prrqUSnT+wEQE/ulhlz8Md1N10zpw+JFmXtC4TpiP+mxg09CamY3D6QJOZtK
ILSrILlMRcGCLzMgN9YsKUm+aQcoKTYcJryk4AlXvQ/41PMFHfATMEkQGbY40Mmpf4RTxfWQ4jj6
ds5bVlc8QljPpO+bZaN8GCGqErenS+1/k934ZyHjBS6FDmAOjLkxlptQEVJ/RlrE/3pScLv6O4Ud
RJMNAYkAABUiqAL4p2JeX2E7U3C6ptUghpWUSIuGnwhiXWtByxN+CrZMyPSYpfQCEsfijQMPTDUN
qgcEaWteUclEvsM9WXKnb5JGSIUqg2QKDZ/2j5nfdklujJXtjTeuzDMAfEfTpNIaVuNXp1PispJo
NryMmGfey9pN1Pytn/nwTZvwRcDswAmndX8OglI3/gYcGDZGTzG/QxYHM06pUIkoebOxf+Sd6bap
7tgskzvKO+i+FcJoTXb0uNbL/HvCuIRGYzTQhkFgsX+37EoGvSqwZz9XXJpKnGSZgU0jPxOtqjDm
VvLrcBEo6Ot2bgGmTWGI9BJ2zRLXYIDx2uXqP0ST0+AQZYAfPbz871ieeLQvPNGW6Vyycw8i2r9d
3RAe54k8S8+fLHUkSdd5iD8/1lATx3VqJJLRYdLTweEoICRIDp/ChK+3Hfi+xxbccE1H214bBMtI
PzwsPwKreI5EajCR3ck8TSnZQWD5mEroyYC8zv841e0Kq0HyHksTcKETHa308jCpO8E3cbcwfe0/
D3SqhwzuVLHf/ReIibROMTjnD49uxDIA3GfyHWm03zGkVmka3ICuaTGjdzYS0fM5yE0kz2X+I44t
alBk1kvU96EzTTT6pVp4++qRrAzu6VHMplQoEA0MmByqePn/oxM7qLTnPfIC5G3rDx8/NtfBaHJi
AEl8yahVwFWCK7IGY88oE/5Lkr9WqAsT+JQMXL817tGXHg0HwuidWFuCCmMRBqhVSF05IajMhSKU
/OUdZXuVEnCFb6I63kyHVXfTSL5BxR/5xN3dNbjXHRHDsPIX4hNp92YZwCQ4HLY4rA60HMa9x7Rm
ujFBgWLw+Io4G+igzxS/jixc+gX8E2bkxZOcWfCUNraWNBk+0bQYycsF96Y8jpfgMYCmL4GQo7Hn
vpXBZBSW/2nlvopWdHyC7pvssXI62m/QDK072+JaZuH/jVEupSR+LHYEzqbvdEFxnWTJgQyi0YxP
kP5SeZSyLeTcb7FB3KpAbdgcu1jry2fRBZFQHgL3a9gLaWE16yTKkBMOg3vptdzQK02KWi3NtCu0
mZi+K6FuUEKmIPgqRIFlDiLfo2a1yvehkTzwoFIVSS9hs7S6jdBXprXSPb1x3iCdCd37mkTK0n+7
bmyvomnZttbl0mWGyfdCojpmhlQBInLwjhHAe3uIE9qykmwCdP3GRTwG9R6UWk/T3HWL4vybgYzN
ozAgDKTHkU1ZT55EJZ8c19XSoUir4+jugdDwpPgLGGvT3vFX+FGiSJucJqUWqC4q6BVBvOxEeLHv
mG0kehKg/rwBmk1P66LFGqeEWLdZ0fXIMIiWXHdPiOSLbyZwSsZM/+qn5KBHRsxZkRlY0Cbl3LVS
tSMfk5aqUYmxWj90YDV1XR5oAN1K4aXd8fVogOM4AsxuhHTiUIG8yZ1nr0x2Pz/linru4R3vQt8M
aNQyjnqelfthMiCoBZ6o9ng66tE5nAQWC8C8k/Eb0aDS8PyGbxRL4znqnwUy5IXV4djc5KYSItui
QcB0+FiSlQt+V/ooDfdNKqqq6AJqIHujMlP3S4Pbua0+vCMQMnjnhA5yFg+zIb+r/fw/js7o7GXi
iW6xkGDOquhzp6b9EAV6om5+xqEUMhloP4+Ukr07MHctraN3nHk2VXdWGyd9h+pE+PULnp85ylAQ
fz/DeUvB5CpeI6ft5qjRYwyRbkw/xt5uVB+kQBuJvw88eblxcNYLV561f228ANJKsuhEdWSe7TTd
wBnWLUMSRw4/dc19TsGzV4UFfm4A7OM+qZ0lv0Qmt2hpC3ZPcM45uvX6bBA8avaAR8ei/ANOT2V7
l4XcA/uT05HFTxf6gH2A5liK696sa/5Z8NPSQ5j+KaH/QACBa2sR9pvBsPhTWGxfkH+oWvThkryn
V+y88+ZrlzCSrLVz0qgb8294eHCkVhEmCV3YGI9uNYfa4RW22X/dmlJNkfnVCIVMzWv23pqsPvSe
ioP8Jmh/pw9Aj2AjG4kvR0mHZw1Bw1c5MX20CUUkMtSPJF68+MN9hWULykqlTQN1ha95BB9N4EHh
0YgmEgeAjA18zhMm9hlVoXOxeju+7LhjZ5o0fNVmB9t8y9LARwI53SR7AXw6rAw4BfjOumexjnwd
UKjDmqyFhpzIZ1CeTum/r4S1/JacMQvDy5IqXlQsA2CWdAZOCAVyyHGa0WN9eJaU+JZ/ulw87WTX
7jHOg0PylnQRjRKDa1E58OGqGJutYG4N2/W7BgcLSx2QmMBaTRDQXA/58H2L5fA26oaJySwDokJl
zg4DcWI0BliCRO0o0BFXP8eoZYM7jP6sbEwk0TBptGZ7evknXL+WCQQm9GTsl64tVzi8fRhDegXo
5w9Yj9hiGGHGPHHgSfEkSUTG0M2xYo95VIXP9/XHP+M/lW6/gwaHvA4q07JANaxOxo9VbiZ38bwT
3qPbR+mY7IybDq5g4PQZOZhVdJ64mFdZ6+3IiN71d7y7T/AT3uBYJu7v+RJgBI5zyjjjxBRJiEzZ
GqOPrfCPr0RfOGjt2tGkcAllXv0rDe6QVJZ+gMtDIB4jTedVvUnj2SaeGPbMENLc/JohZTw0hEDN
jKdSLqO6rFCpmis4pf77bp3Bx/ns4gbCpZdV4F6ReHhXDVfH1XQuxWdnb6kMHHMLI2zxvdKKDLW3
DwMkQ9hzcQTC6gc4qdefq7VZWTCCLczO91inkSr4zrFB9sNBBrAFr2VpoFzJ/tCQHOHlZRZ7wSau
5o0PiSevX9huU0PK4luGSx9SCtr2MyjQ1K7v3KX+VAElYX9ldi1rdHTVdUXH1yzND76fbsdbnxM/
ckQl8EiXbdehMBs/WNABiLF5h0685iphde4FQPHug9XrRb8vQPRTA9zFeN1CpsGBtNNECU343CD4
GXptNez0MtYeFgz8RovV7Q9K6TInogxcRCKLv6xLACQGRE2gCG1JPJIEVlaJYF1CkaHenv0IsZDM
Eoo3QFxsiM65UMS/dtIXysZaYxx1ziRLu1dXADZhL3RePXIjdVmafRhfuKwj+THUucK2XKeIvWKl
JisyYJTIN61hG1VKiszd2+wjSiA4GCz5y+068SYpc8jNmXyJN+/trguunrul+8vsy542vnZsv8H1
TkHXVOMoPkDa6oXjklh/7pEwvGTtzVdTlUds+uvD95bW58DORwnvyz+nmKqUWLcEq65CXn3TEb52
LzPCZ/4+S124Hc4CcATuHADfl4sHcJSe8sJZY96Nr9jqjTeif45Nvt2LqPRoxfItsB1TV5TMQWSX
0Ozs+I98tmWHkp3oMqAr6v7ohIqFfZth/rJAGqRZJbA9Rt+KjgWS8/RnUsxkpabOvzni97FCyyNE
jdD7FDSJUfbd2ng0ACtEWppLe3rkRq1nKsty//fDtJSEICUYasBdkRMxjJ8wxfDDKaKNfxQV23XF
4DNTAjzSO9HmtWhxQPMjUmLrYwLQ/lLaRk060VUe7lXYo/atOf6o6lOplP93mmG33e/UhTmOrCQH
LjkwBr0+x30fDCghSzAmd5zSsJmYjuSBY7oujqlOiQGkX39kXYYrhkvXhBH5nL+g23Cwja3q05T4
cAXaxjTZLuHwIJFup4shhQ53v/tT86zOIAhfJn/mIKq05TenbM7CHeuZA918dbCHNO5VUrHsY1Nx
UZ9/y0+a1s4pl/duex2gZsP2zHo+kv1+hpcPnyDESu/nliDG32Yjde29o9hRVCpRChqu8WJWkN5m
ngkwl7s2hNLV97FJ4NFteeCijMHqyvVCB2AEJx9W1UzysTMnbamu+TgdQ/TO0m860uPJjJ9VpIeY
pvz3P3Q0K0oM8W16LT0y36jybwkDvecn5Ae+6p2EhF/dcXAM+WptyKX5QL8rKrk0VSpm9LHa4P5e
/L5xNVrmpvzfmjId4hgRdBI7SaYswnxOzdvi9caTS0QyHYEVFw1CyP4c15rvrBRAYJ14FbS9xt3L
fREQ3pwnAwOqXcvbxJ7DkN7vO0uutjE98R7biGvTQwYFH7ow44g9mtDwNxLK7cj8daglM/j+vm37
dKadlwlLPrRhlI+qaJhbDqqfkd+NSkxp+8OXCRf+yp1J9R1O1hZYLmRipfnptZZm0dWJIvHPV7Hs
orqS5bhbc2iDLSz9Q/W7bvDM/a22it1+MpznkG9p8Is16oX7ZPkLJWTRInEyEybGcvrzyP1rceRz
N6+dEMLS5DOviSW8LkMSUH6lFM0XJ8m5zt001fEm7puyEnAz1gKm2cnsZma0pFsrL9Esq1WaPEBH
kHKC8bSDC3EMT0tk0AcqHSmC8CTLKfNQHrUgeytLftFiSV6aZ4iGG7xlQSQlR5G7U8OQy2yFAX7H
VD9lbh0X9ZGt6HCU4abcaGw+omG0Cxec2K3OqYlUfDvYIswqaHbVeZWHAye3XzWRJ2EYhwP7kKHx
IBcllcHQxuJZuljKlKtQEbut5RTvASOEUp9e7xMq3nDwSmypF0hRTLl7XeNKSS6QB9XxQ5dbRPBF
yW1NdPpBXlubYeYWkSFGzTq00YaaCGAxLUBbh78qnLFWO/8ooPNFbC4vdC1Z+4reRoBE4zDz9wvj
Hpvr5/jwu3Vgj8bhUPg0AdfbVyKJaUROwa7v9dKG1Fl82IJdKhAMrB7nIdh+PfxrAJNxgQIB7MbW
h/UQwMTrudlMYEFG6h2VGvoCkKeOo40ClIR3kBi59Edjf57hVOJtPrBhxQVfVO6su47buBjr5JcO
/hjLWZcx0vfh8XawVyvbpnv/xzTrTv6ggJ/7Q5D7FLZJp08OMHE8BrCf9xhd3GMz9Z1zP7vRfSYV
YEkXa6sZ/P8MiP26/LtGMrunlE9rPGZbZLAehLoRt/4dMjYP3UWiM5Z74v6KVh4+fFhfFHH9MZzP
3ed1kUxRBTokc577rEwavF6wKES8cEIrnOvMJtIVwkgy2tJ7TzX+V3CTf9tPLckC+XA7/47lVXPo
236ttxB8+HaeIbFlxn7N41s3CIaSu4IKSFA5/EyXZpe2q8itTycx2uJMVjzFPjfjk8U4o8i68I2x
bJWj7tp1Eeo02p/BjNoHY5H3mLDI07FSvS+rzOIzuv5Y589alzVTGN408Z4WJVzpi32q155493f2
EAYG/mLSsAn8HJ7k/Gedh/I50qmoB+JEF2iTyI+phI9Kfw2kJUg093JKCY2w5aN5jWFo5yKq9Knw
dvQxAlGotdSDZDpBthzUvVP4RFokifCdljiT+Fcl9Qned1rpc6VuJFfYEQWKs6MP0g4yPs/Dj0fA
5dEi4D+gD186yo1AgrgoIpFbCmBIaI9A1wcBLBzy0hK3g70ZcUbniLWl/gwDPWagjckK+aCqB7Ks
wbOHN7Is3UJBkBAs635p1UNHwNXXJPhqrcSPgl7vqAWcbah8z49GDBukvv83Czgj3djAVhePGBE7
8J8hwp2E88Hd/BLdncjE50/+zurDECRgG0+YZTgwp9hhJierGB+yHozYdbWvpr0KAdMFOHOMXbn8
qP1ShvDnO0+5/sDU4UMpz0U83kAYr7sUIjglO3D9mqkz03pRjj0C5nTfAKTFs9qWjeLiP16cxK6K
jX1VwPDdPNfiFgqdNXWrKPEcIQG/o/f9+w4rIvjb77oxgyooNJ48qyVL6QpYVfpb8DAi9C2x5ckA
jqmz7L04ibsP6swZy+9lj607PEFZljYn0gZkimdgqLuB3m3rky20bHl7hivmtjMZj8u/UndnDTf8
6kx8vjaqYU8VRbj6319O7YK2Amk7mXyNZMXu2/+yDKt/h5EW24PUvPTyMriShSgdRZMR5UD4JcAl
xgtX7cD5+T4dArk4uKeP75F2/3ttmrzHwP70BsV82U9y4zfyxVnwn+rbE+EhayJ2fUhxzdrMv0co
o09xcq3d1GllYvl//bhOAv5hLewCWqPmOPrBh9nzJUpkS31muppMR4OLQZ5CVvSJt8GUh+10jvuY
fhMGQSIWX0zws3spJ02vbLvHBmrRAiC2InjgfMorEnCIUlYbIsxIkHMALtwylNYIeSUykKjLWmo/
DAuAFRD6Qt1h3QplehBMfcI8TF927kEGw0q2Ckm9smzHDzdIoR1lwVLQrYvFP/JpGuGmsQLBofWd
iy3oPyTszqh4zNTTCvtv/h+5RKpCgEKuZzSDmjfslUZa2F+o/hRG8zIcf8yqjOOxv1b/ef4Kjve2
O/1sHF213odBSKU+ycECJDBK2E8pB487FqxyAMi8hF9Q1hIZlLnki6qhE6dQ1QYzhHk+2fqOZsml
Llw0W3YhOppiO3L75HhMZpT203mY2+AP11urSNyLanUjhJl0KhvWjweh/sMPylQss7eMMfeThVmP
RAgMhinH24xE1fR4vbTFMgAR+EPO3s39VT96Fnl6p6GstsRA8SjJpyNZ66a0NdvuqNhBU0aIwuLB
at/eoUcF5+MIxmGjWxTNuy+u4f9UVU3iqbm2fQwNtUueBJo3lmetzFlaFSdRq9zonh+KxcXRCiFm
YP8rJpjDJI439MjtX5VLuog0S8O2KC4Qu8cqFijO+G4j76F94oMz+rw5rW0G9xwB3UFlfEecybaY
1swD3OkU+DOfhD9TvOMhjAvMiiRA/2uVErzTsWoxn49rtCAyQ4VhXIQqE0xVSsOaF2HlXA4sdtZ5
KFhjSv5Ye4pNq9iJxnY/MD6zknXqNJG6+GRdAYZkwinRb7TS8qAY6QirRVIKFOamt0HDJhR7MueK
Gmd7MmCd+cdWvjNqKQ49+WFFq/kfuBY1v66/7Hmv/B4Wv2joKEFoNi7md9FbpjcQfb+tAfMxHNbm
YlSramCTQH6aT2OQAGuGSiBwFHfVQyFsDFjmyAWSmulN6QI5FxDMfG5f6RrfjmjFfD5eAWkZ7ZAk
bNne8Jzvu5IK+d4NlQfWRO4+UQ3f7TrJiOiiKDJ6YgA56mPDqobDbs0aEpQckTuaOIjLJeiKVhQP
TCgH8fldz2GHFqD7d+6wygepldxHR8Flmi6ChsnnZ9PEMfKuSx4cSKV9gIW6TgOnsQLQCxgAcgIB
c3WDKX47+gBGkj1eWL+jLdmGCUYA9JfnjJ4Sm1Is5LPzosJm5EKrIgjGD1W6tLxnCAsyhb/BhZba
QNUvTzWTOVcRAtbLDaNVV+MhNvogBob0uggF8jyXADYsKjXn8r2LJDFRddEh4jETmcALWREoUXpx
aEDB/XBYIvWNEmRSk8BNIYzIE46MXEw2Dos4DzlAbu4Sr+z+01WXtTOrtFDfOgnkyfeL/1uUgaIR
tgPy5XZg3OzJGiugO36jpdysBd8Tojy/tCzVk3qpr9xzgDM4W/cfRaeSLWpbiQzePEg45EfH7T6l
OmrY0bZ3GD7fP1fmDydeo0/MIqVLjkWX/tDMNuS6s6LiW1ylxjs1Z6iWFcbqQMwCvQa1D+IzeagN
+tIj5J1ShzNne1h++Dlw5EXk9moNDs/BMPBeBcNQzRToyOEcuoBijaC9a3LAS9O1DhV51ip/y9uV
o4N4w0RI5eReG5pikmUA6uP1CjxbPm61sxbphYNUhSNfspm9CiGa9GTpYtKyR4i2Un9Xo3Sg6TYI
NhOmFhcY12fI0LuMzTqHD3/tmVGRwQrqLztDSqGeWt8yu5txDVQFzsggs00iAZZGN1/h2w1Q7GXR
CbXp0trxDt8SIbo5rZwLdZ2vu+97jqTuVqjEo3G3TDvyBimNF0NhLBGTNwMf3RCQMbk9aeceQaiB
paQH5UQbuRyD6HnBdlQWuu7lmEzx9FisWG0foGGCJxYcGA8b8DpK7sPVXxIIdEb8iPOZtaFhsUQP
V2uwfb1DhE8gFK2Tc7aI5upPTDtjtU//rmZCEUvBgm7yB/8mCkvqgjQ0lhy5ddehErjHdRZcP5uf
qtZd0l78iVi6MWYDPTeeMRAKetbSp6TBeOQQt6cGlIG1c3dfmFzzjHf2kJJKm/BOOToX0au5y+S6
69tGux0x28wo5VuZ+GzVZE6LtTIlLxlPqhYkTkKOMQ1VbgdlpV+AmrNEyBMq4XlFvM+Br/VkBa5V
7ALTls85qvAy4JhaAungm7+WLX2Qn8O/H4Kos6JoifsHINiTBEcJ9tKps72FcRFQX0ZBwVAPe11b
JB3KiNiSOIPE7ecpIQ84YI4uD+UqaGKn5gBCXA879eP/r5oa7EgIsov1JVCY4YkfZNbGtb9//Pc2
uxnyH7mIUQM8WUvPVxiV6xfRZQ6YCffrEBtDAPT/WO81MO5zq3kn3bEY+QfIHsWBHj/cUj3w1NPo
t1AzB8jLidkPRN/sn6diKQSpMxMSwQQV/i1rFy6tI8pNBIWMUufqRdaB3vJO27jFJv0iqPfoqHHy
UNtj1/qe5c7c59N8gPNkeaDP3lIW2n0xvy19avYGXENyiYUfwCDQXTPpXQdWQfH33kQfEAgaPOt1
Zud27345SJY4My+COuOX2nmeGbyGwC12nEAn/Y/sp8hKg2cFi//7/2iNGm51lPiQfCYnuznU/M4B
zb3miFzl6fg4wd21xJgI7O27X5YLyto/Tmwy7YrdIN+Z3U2CKN1M1j7dJi1crMVush63iGs5el87
07zHK6MRDssqHjdGgNzamvrj67YBs8WyU+ZmvX3p7degacFbYULEXVcfatNn7MmLJNbDMOwk/+i7
Y6mYsUd8l12wdaCZ1XEktWpsmdZye8+h34EPPQ5Dw1xhqn5gQ2PNJzLBNPQePdCpmI4Cr3KHgXg2
id5/jTT1vZwUGbh4OWXjl0SUMLgXDesTdv/hjX/E4F2P+mmczU2vTWUwe0kqkmoiXsp3JLJkUN3+
hx/j7H3ZsXN9xQG0t2mKB+j47316kZ0b0Jcwv7cxRM7c+ouX8YY7+OfBQVeZRrhGlDcSAUym2DF6
SCbo7wKrZxeu2OeJh3vWMHleM2BJETiKoOe/2eKVf1HNBqugyckfRT7Fg9EOu+QA55XCbP/7i7zn
sxfpOgxo5j3QtE5uwXK12iEJxSCHCHvYy4zxltEWD4SbaqxyRNF1SFQsRli/9XKG4FMGWZA9KsWP
Q49+UVj/TyS/zLrIWqs5A0ADgKsTCTiAitEkt4I5DU2eGWEea36vvi1b+ROQRZQv7KThE5aXZmqM
cipJNg6TCkOkvIzdXDeJICxOsbshcIPhkRFbQnKXxtHduZPTRCTGyHMDPbf5sl5e3wKUmQsE3ShL
rEj9xAoeLhqgD5MGMLbfjP1i0xcD0TebhJ7BmNVKt/yBQsNXr6Csni15JjdEmA6Uw+hOB21HnSPQ
LnJA8Q7rRj3RKqJ2CpSIdgULBgjnT8nBAJSpj5/xUnQkh1vPCuHJ4EOoAHTOnHtlolPjpcHFnT+5
1UIH0I/akKB/NhMfEHyDeZ0D7bHC5q7jIlqqxNfbYkMMV+8y0OJH5Em2PhH6fDiSXcYPXDOhMYkA
7uvwDZGX4IdlFzbETPFC3vR1cKeYhur7BroWY9j+rGhnHmDuTHBVM4+i6XW5z+xl6ThTohNDp947
NFkA8F+3CbBdPtJT10Sug4by5Zv/HmzsPY0viKX6xk1Q8yI44BaavOq3eumuZi2zixMTSLo6J/bK
ntdR+iFZxC2Gawt7CQpCgYKXKcoRnDql+zV0kXyjJj2/VfVgJRy2xHAskjs9hzvO51PeNk86faxh
YqA2AxnmCYGYs6HW1XJVb19aQ4B75QuU7rqm5L+42tInyPKyZpu8DfHbnBNp+nLLWxGeMb5Jep5g
3HtMixRKedXwO3ECkws9RAsc5/1q8GbtUyLZgPvM20oumcYV0vFtZZ8PwCtctOW7AuCvnsLlmP/5
L3ggLMZfwXoLrONOakH3KCj7vRDTwBTVPNoiS9F9+sMruX7py9IL0CZ2PFID2OBxg9VLdAwXYuCM
fyRn2ka2FFGJ96DIrazqJdLvw2JG3x3bhL+lHzjqZY60bmP1UZnPMyptvud4Xm61S+sZPYjYKbUF
fTegkW1FwLOTpoZBg6Dh2kq24GQw55EYL5UMx/0U9jEDwm4JqpwrH4fYEaqALlyR4GfqnAFVn9fx
QFUVeKkxgesUK2cwcEaChKOhv4Ycz7h1erlG8WO0jCWlhEAh5ZvfdYICPjl+p/I5S2ySXuG1ClVV
zooZi+a9SuNHG711IL0JeONKxExPES3S3MIVpnr+POfvCXBIPcDCTt0Vd+OunfDE6i8vB+IVXpAe
zNFQ8s3zVqSgUp6Dux1lolJ2HuIQ62CkmVPCfLOe7Cr3yDZwEnNMYRhJ4QbkR1mvxJrRQ63FMFnp
HNHBhN0Cy1TYMF95jUaTQNhnKCSDjzaacwMmupyJQusfMt29DVQh9pACjX6sD9CaybNWrTz2JIXR
oNCSwN+27yuFToE/glVHBxGalIo9J3P66GRJprIZlgojXkbqxgs+T7IHgPWNm/YwMsvXWU+PydXR
GRCDMdyJwIPeHET8bs21mBXBkgxAaY6aDn0rwpJi2xBV4sHIXxGxhlb6QtqHUaiMxfw2zEMUrbhI
ldIscRQXKJEpV8vDN2D/XBYqP/SQBOJoTmS25rpHyTI7NckbUdGAr1UFTfhy5GdUitS2Z6JIdQu3
pmTj2W557153bqaT+9yWTi1Z3lWVrbGMM26ivEnTk35+1V4Ldid9saweojQ0IpCg3jMkeKEegWq7
DH74Wt3O8/xP2NsggNy+vdJoSqb8dNNhWLjn1Pjz20kT8Ar3o9nLRaTgipncFowEp51sjFYmHuOi
hLxbMlCYaSadcQaW69/HKGiLReWn37qTMaNsjJupbdLjvxntfxDmDQx7OQlXuYvelqmDxvY6JrKO
HNL8tLR04J6HjBBSjpw1pVEnN9djvRiA0AtZMGOE/8XLKeeTWRurTfjQBE0opUPr5o9wl5NlioHd
qvf80JoiosPkyge9OtLA9D0YYos77eBZG8VQ60uW4s3ah7KkgCNY8TatTYwhSZMhviHkZaa7jVMV
4poQRQxIeniGmppHJMJ/EZ/ZAVJies+zOj/kHBL+4eGLABN3QEMWtZ5ENOScSXU6PisJt9XSdsey
Zxq62hU3XZfwmMcxk5y+6XbKVXIu3gdfI/45kEOdRvykUoPqvxz7PHhhIceL4kP9+kyAH3WWzsg/
ISiwJE09qPv+Vn3sIecMQ5OCNMKF5sVuEJz209usm9Qn2FcvFNUjtuFQRNc5zj6tfsfZ4yUmG3ZI
Oxi7MByY73iby71dYpeYb6uhoDHv0yomM9dG+Af3VKlAFLIokDfzFuVl2JyIdzBjHDvWUhwTuSoq
f0/iMDC46nFXj9CJ/KirzKIPHur1nRrYsUV3zfScr5yN3b309/bynWZeR+vhtc5VnID+Z6bkv2FV
yGrG69jmuBE6fDTYiYau1WHmZfEM6i8Qw5baqOQ7qag6obrE2hVPQiwiv6hQD5DDgJC0u9uGDNJP
lo587vHNdgk8V0WdhqdlJoTk3HgIEt+JpZfflsanwszCBp+VuM4LQod1f0JclqQ6wWRNKdO9MYDq
h/aD7ZQX/mfmOSpU2kxOPUbiu8YOdHgMahwT5F/LiMbsCT5FafDF1fdF933ID3OcvZMhE8+/CVpt
C0SuwYDvSji9aoQZRPVt8Z8MhTHyqRVflt9NLh6HoX8XIzq+xgin4n68YHcFf70J5bLn8C/1XenM
5rvEDth1n/yMYv+D24mX0eGDEpuCNDYBfFb1jdOhroHzKIGXF8Qc5cpQ9Q3TUnQgxwQens2Sia+3
TFLzCl6GrUUcNomsKaPS9Do3DPW1NgQafOyc1foQBnORkzZJv59BAyI/a4X9nSa2x8c9fz+iFUe+
XSIronyNulMM4s+UeyX+uNeX9Y3j6XshZbaT5lEc53hIWPtrmhk2nUOeuiv3MgVUYxvVlOT5wrSG
ZLiVr1IzZL8wmlooqPiQoMFbBg2AWI01E5nh3MkgsZ6LUc40IsaSHdCh1BLZT1CuFZChSwUwar7K
8MonaXS+HCBp+9Qr7ag9LQ4v1IEzdA/DHsEiH3QejzVu0U1Ipk28HMUSC/0FJQ2Fn0ac2RIV5cfN
hnguyc8NJ4KHQbNSzUEt5Gns4vhvRmMc6mG4/eMBlW2zJn3JbGUnt5QrcOSgPp/TEZiQ8hd1Lu81
oZP62343JOoSqJurLy6AurC9R9mviIiLz3DXWY5rImuiMZgK2tEYDYAEx7Mzemb1gscrFh8Zdrgm
KcCVaTOtZhFCWrecFyAyhADq/FssTGUBVxGtm0nF4WdE5i/LCYERV3lHBQNINOa2SwOH245S6dC+
OA7+LmibtZ0CGMVWsAkdEpSDiJ+vi9SPxTbYplC0nR1E7YXL3DukOe9bB3j/a88L1/3eTYV7bZdb
ROK8/vCBeiDwpTwp4cPG9ophO8DjvB7Y41hTDXetzqJEhjmkPC11B2/S1yC1TcfhLccILJCVKQ13
CsMfp+UV1eP4DXvxGkbucSu6//tfqxAzIHuI/1LwCJ2P7pUh8v9oFaCZ8Wlpxto/eIDGXYcVyQ/w
Q+xAKdk5wBN0k3zRz22cpq7qay65R5LGMT+PZum7cBS4mAtapy+WWqaA+qVf4liKIE7xo2xKScl6
vArUamdJAJMXZ9KaO4wXb4HCmUHdr5wrgr1/FjT/07coXXHENO8E5pmbRe5B0ATd9B04zMTmoWcq
ffcCgtjjpPJY1TVg41Xdf8x5NkEKxZkynPzof3thDcHmvENoN0DfCTg4b7eX8RSY675NlB0V3ZeW
BJlmSr+dIop38B9fQcR3WftqewAfretw8pD5yS5UPGowbLtuqrz6tH5RzcTyk0uy1Qe5Dv4WDdrv
Lk8SHJxDELMHitigil6+A2Hd3RvfBgjXWuePCe/BtuwM9vxQYvyqe2iXYJRarChgiCQEYrdThwPV
iwJxeHOlkyGl8p4gPAF//gJCu8EwNZzma1geegEJ76XOUE9/VGm4w7EkhB8PYmmcnPWhlfsSaMq8
2pRGuY5DO3vEkOfwEimaF8nxyqEY8t5WRve/dxhvt1XkDUdSyln72ktXF9+rh/cvkS6Gv8LKH6sJ
0UmFo2PKE3ovxteuBDWMAhbHffyrM2vwe28FPc+AaUrI3o/Bl4khYAVNphuedkrl812QF7NHDyFY
AV8KKrx/BimAaO8Td7/v5MRcXcjXqn5sIJLApZnSaWSVeaxTypsP0g6kYXygk+CO2PPhY56ZSlOb
26zjNC2FKF+4ThC578vj3HgCnisfJxXlNO1sWDXyAgTbm51CYS4jM9JUr6zJZJ3nx7W8F2VWpmMU
9UL6pPPsTUP9RVXITcW9kuuk+pLuDWDTqk2B5nSokB5JcZj0p2tsuDSfkaLQQ55RETwq1qmQ+pDV
EBbLhVfB3EW/NJKJm5KXYEIMYeRRCh4O3iPBTjaxCEA07DJ4eMqMYJ1EfpeEa6r1sDljh6bmlv9V
zJFKh8ZxR809xWtpUGYnCjS87GHHyb5h6ywXQBFbXdfF7jCFZwOQ5QruGrl+UW6Q/LgQHvGPyKM8
29t2qlhtxhEbayCzm8lyr7rCqhlNlYyTUBLPydiYJDDVgBRnB9w0VDrWOgLjcYCFCfXtyUHG0HQl
hsRAiHSf5LnlAVtQCdZl0L5UZ5vcFwgAjPBeZM3hfCmOCiyq0hMgYOUHoRu9fN58QNgfUFHxwbJZ
kvf7rUWBQbWwMwUfENv4qx14U3lcOXz0LSmtO5Y4Uq5fS4hnj9G6hlBHokl9GUtVy5XGS/HtVJq5
zKQEnItWTIsZLy/2ilEDrQKz+AeTA5wE8Th5OehYjrurgCbLeyER58f++ZYTdxKq8oblJlZuDT66
8kNrX6LC6wWX4JkBfZEk5YACXsB/PF/nr9DsiurZx9eKqKe+0ioqH+C5ILPvYz1OJyylSQQOkQdG
MX47pboRz7xY8I+5PCxAKARPAQrjQNl5JMLGojuwfT2v7n06H7XBt3nfxcEaI3fBbi0XFKH9zyft
trqtLdu2N1+xWAxasKb0Hj/H3pcT+i2M050/HcCgWJVTiFsoi4x7T96xn8K9qnyXgBeBf+LVFCZr
CjV5LSy4k7qpOU0XwzvmOZdA1eTfEEjWl+zw1e/6hiUMWB4QdNXCaGSG38wUWOL94z5xtkokDjQC
MJipZuSRdOhMml+R0nwevn23bvECjJMteRjQmPVXrVPYvBuIyWgaLBdmlWanOoDFJ4MTavFrBRmG
NwA3BURLoi2rvTZyK2lz2X6rNkuNByNOes4nnx34B4/uYn/LyDKT2eJ4GKnhctpehnQQhUT1hryt
HGAxuF0fI5ggZkq891bOIQewsfkaHgIRd1u52DNrKDrerkCnUqIuWjoYQoIJ4umFhXNtTWelKCEt
4D21u8ZNgj9cVO1AIAXyDvziA8+AkVPEBFbBabHjttqpkGXW2sQREC8WAfyYaG5L5b4+3iwqzpZH
xEhctaio8ykAEWLllV4Abmnvtnv2OIRPgRozFUTF/YmNeS+rGl3Q0GWVqyiIMxcnoFp1sKGuHTxG
t3LWKAV7D+jropd3HPb5gJZMZfbBcJe7ASykRn1MkhyVbAOj4VvY7M6x0oVq6GIqA2voCeAvwDvv
B2xMPtXsifeuSfMFh7ZrrwOZlmsyjq3/DeMms1O8PbcaV34C2pUZzQoWxOYByDx0fz1tNydmeT35
seBu3UBIaTCbIcKOksTTbHVa9fE1j347t5majrQAxVS/D4jdRQGbqkmYYBiOF6qh3npZE81i6EDY
OUUglPGSAqT1E12xyOE51DlApFHZ29ZXKt1osBDx97dYUkxaCAibs8PKnS+Y3BmENZvpBZqHWOH+
iHd/7Xd/YePuNmOZ3OyCX+/y0O2Dl/6CnueJeFsajBZpUDNdgwCJIjF9+UIe1xiwVoMuX6+5zogO
G6zHM6Lu3SsAhT1LfiSaBajGOl5oi40Nr0glsV8Mnz8u8ZP3dEhzOumujrE71K/ETbaxqKPISJbF
KEmMdlep4RHNdKto6vZkiV8Z350eCQpbDusWy8XpGSm6JNuN75wtWboJMHOUnll4INAnfEeklrd+
LDeOQhMrU+YOx3ki0djKfalROc0SlH/vBzt/lk1FI+g8P2UXpsSowRLfCxl266q768opXTXjuvac
GnAkMn5D9U8qIM5yKBGvSIHLCDAwcFYh1CoL/BBOTfSI4DCpsvW0SyiscB1q4jAgQ2ls1fr1Ryad
TmSTtJaou0RTsj+U7xM4bhcspJsmIchyfmD2VwFmeyTXhNee6AwlKjrg/2EdW3inGt9VU+1B8qnv
t8LWs/ebCAgDkgCti0v7L6Ev/LA2Ebekfwc8EMGePhhtTbkduLTAi+TYQClUFPuqRQoiLUOp5xhf
lfzyRt0OTj4YJEgzUPNLWbo9I1N7sRTTp0ulibMinkhvq6+Uvcb0idkxECfKsXAYKFssd7+jfRNr
TRaMv//m1TrP7zRAMB86XW/vP6ughwk3jUP8P9jUcig5iGQbbSQnh/zHBAl+ioAuV5KUq77gyLly
Yo1ueDkdRllc01JPiCEeWuoB06r6opByS9hzx9RjNyrH6+JXh64aznjwcWUDipIfbR7lqXQ3UahC
q+UH/SOy698tm4DTAk1v8aZ1zzo5mEPQzj1hU14xvJ9FT4omyb5JdQlcLjzND2pHFNknYyEH1uLL
ar++VUtqOi1Uvy6AvM7H29wy/QEhosMSJ0wMfPJZBEOw4p8hLbJxQIgwCJZWI/cTW/vogSi00qd8
TtITJDh/PxWOyq2SxO+XP9uce8+wajf/jkNUN7LyD99LNDK+cJ6JakQewmvdLrXlZNfI9aB1vMfW
YhQudNEMDoBlsq2xnlhf/AqibTVFnooe51hWKpzQ0PWMUi9Qo7V9so4XMQUEK2+c+4G3xxZg9kU8
TTsk8VMeBkRxJiMiqiVmKNbVPmHqhUa4ZKd2ZX4zwdSRDXOKeAtGB5fh3nUj8M2001QCdc912bWL
xn2l/DZQ8CAid7YLawbgd1RVoN064c0xDmopOwGTdwdDBV2erStwZExzYvNRycwbU+osGtfGgX2b
dTCs8PRPYQ8zw1buTs8kJouExl7TXylezS0TBlkQxex6nwKzcAckAcQKu09KpgAVWDJVDNlMbCIc
J23XnCAeGJzZ+XA8Ici+6Z1rZeA1Po+WqaBEBN5H7rEost2SD7PSpb0WlW393+tR55e2Ggdzqj3z
gAO2FiJuAoqEWIGjEnP51sgcczMdGXrIYWtbxX7AqViI9t5hmcDPPGT+FzJUFLu17tqHnMbWmd9A
kPGVdAYnA6iouGaAEwjd+5tnD62dfiAsmzkBa6JPE4IKetTqNPXL/vEFtY1BIbq0wWPI1PC46EWX
yQYhShazV+28rP155PGV4SXNahuwDzWtRm63mFRV1LKKWu+yY0zyTmjih+fl50aazl6IVhfiUMuh
HhK8AgdTh6yfN+cMsnBxN/XL5FiguUqxXBpPNKrXeKzE4zpM4IhpleLeOuzfNv2V/WcsBiNEjh5Z
yORpmFC0yfgo3wGhwWuja/e4GEN9jtgn8OPtge7rxX0scPbCcqdaPwy/1y/vxYY5h9LJvyFrhqu5
vtenLNhJc4EPGho/gIl4H1kNN/e+EuarN2XfwcDb634Fvsgo1xLJzvHOrUe7GST598LJ0nGbIvoP
MsDl+kUkly3OvW0QgBKKgjGQGFl89lG+JWgtGDYAASnwUYh6yqciCHMbpwQrlFBIoNjGC22RvjUm
pv/u8i+5pbNOhawJB5AxvH93d/13w9q8aKLnUAT1KegHfVW4R5awiGo3uIE6GeolatjbLDO9MnNy
ERoVMBR+Cr8UshMm2VY+CJuJk2rxvETBvD2NUv6dc4KBsBZAAn7TZeJq7Teiw1qixMq1LsHUsOhV
ayaD/JGDasTJDk8uIujnw3d64Oz3fElEFchU3veKhHXvDdYiMcK6+9rAdmKmm7lRVdtXyo4eaZyR
rRf++AlfY2CXUsXrTO8XEIU25R/LNbCCtMN2EGFCZgITg0/q46f+bhyOMqOHX2gsMbiiOln1rurU
miGX7n4AQRbYe3R+ZcFS3AYamxE3eO4oNh8Q0YQIKadoz/Oi3++LtOUvFk67FR5evSnUAUl+9vYw
x+WZltYFLbcm/ZeU2MREw9em34WimzRFtY/GKIl1k+mStxY0Pw+v7BTcFxkT2q4fOgo3Hd5UAUYo
PqJ2R56Qj662/o6z/8mwQB/3aR39LsjxstB1f8sMKYfqmoAP42FosQnb+mxmR9C5/db/irnbclqE
oJbigX8cpvFq1DDD6oMG5Qyj/vFGmuc5IxtoCno2folI4a0nhagr/BT45XEDkW8qqokUhcloRefY
uBzSF7RQNYR3gbuu2WzlCoaCi+D3lN2+M4BTpUdxiJkh0nGLM9T76XD3zPAvQXL+6D+vtPvZ+uSo
8jH9eAbWTIv6BQZlzs1GMSawlJpReyYZfWN0V8O1y7VcCMTRQB8EPdCzLQrtSy4RqsjNEdKeQx2r
HAVBS+ylqkdLVrjARuOo7OSQ1x9cGXZSlR9NrHHIipUVmkwersgkw18jJClJ+9orlVNhLpJYCJ9m
iVoS5BNCjIGYiznvrgtMcV22iPbDdqFegqN8h0K/YCy9k0LV1CxFcONWazyha8YXlAkHj7MOfqzF
zVkEl2QrlpxewjxWfON5m7jvpWqROPZnEA6B+7JbZZLUpp62vbht7d8KZYg88bSNcK/OGLcCh2hR
+fjk34tI49BGF2tVP2Xop1IRA1sPcft8b5reIFfapG6bM1TD1vY9vgI7VBfj4cFMSVkjxx0RnG+g
Wa05AenMv55GSgT8xilTC8KOgXOZF7ZzvNI9IRtD/vmdiEj+dDaRDz2lr+xgYwtQBXIs+bEEIEFO
2yrucO9o7EQi1Qn+r4eiawQRkPplGsfh534w6p/r8hqs2snPD7/Kbwsvdzl8Ll+3r9jRirZHX7A6
l9pUXahamalrGWs1NK7Fej0uuCzMt6I6k4zmEfjzPDpmxz3gK1g5rHrAar+XEPvF+azat8X+/ZSe
tITYtOxtOLr/Qr3hNY0NerQshNhD1hpTKNzW1hKvvHt9iLnHz/WuSuHKgqDgcAXEDjNeKgUmWgCp
VMX+85/fw5+5mgR+obAWZmtu8i+ttNtfu2QAJgAFMm2s46A3Lx99H+BE3xrq0Rz2lQTGQ6kVBxPj
XU+E+qzx+LIdrwnzUeAdPvcsi8v8cT55gUliyDPH4tFkBgf2/mfS2YwcTHZMIFESrlRqIiTcPT20
bLC9rWb+MfmWyjQVDqSaX456OhzXdO+uNV6LkLJqjP+SV7sJog0ALWm0hQeQCW0Q4lvna/aOqfTk
fLzvkxlOEhUfa8fAWMlUJGRRBu7G9Gzlkdwcs6XHMU6btPkG+gkoJyCiIIYq8pEt4lHPJucicJV+
Bbk/w2TepcGPwzy+CkWODcntHJGO4v3vqBygYYG/5SohuQ/qYhnoP5Fv1UtkOrSql2fCLYcSxYU9
B7rTd2/8ZaI299CntKEMpDT+TKxcaZRuwl48ooKCW25uReLV6LIMHRF2v9+kn+9PCPy0Efsfxa3w
P+ujJaSnrzRc8vvH5Djzn0P+3lVLuAa3q3rwajPkoO5jg1RhoCsppaEYaS+mrVUK1g/vVAfM3dDp
mVwZb7FGX89dS5Y/zKOLPauHfKFU8LITxmM6c9/YvpW/Nf6hfzATrqaTBVJeyW2mPeP5k6JVUUEE
2p1f0x1JidD/0Fw+CdLF1YDTPmeZwFLNPsYQqNz+cFOo++ddV5ZBM2NKGl9wSosJ2uOEnFhvfChn
rreR3Q+u9IpWHkrWTJCVphBoHs18Gx+HRigtPE4P1is4tTU0C1vkaHcBwEsczJCF4gkJV+hXtNak
sjXrG8R6AnYeZIM/2/mE9xokTxLZdeiws9dgtcZxIyf9kRcq5BhVMVWURdxRgCx78JBpZ/SbNMhB
tfVJJ9O85G6JluXFb7bx8y82z60bkjkyxXJRYRhslss/ORkd6P6awgi1CoulFv5jqK/DEItLGzXq
ZgnOrkk9dXLq3iT7PIpLFZJegrNYqnIV+CA32hOgM1bM5NMLqabsqoisR+x02UjzcRjT6y/v1uWd
wQLhbDkSoZzMGPpkDfmfYwl/YMJ7t42aU7At7D4Nlstaw/RLUhmB6uQxgJkctg2amEDiJO14SZX/
aPD0s0LOdK0jIAzoJlLqGrzZdthmypGbktCMu78qH1xO/6RaKs4l7zJWAF8qdJGybX0241hbhgXE
MUDYTsPXDSFgfNRCrsB3O0Ag0pFcx6hRwsaFUAvocU1S2v+xdt8mmjsEzyWHl/kODXQHnTUuO0xy
SI6/ED2LF+qM9nPJML/YTWByS0e5pr88xaur+OwpEvThEMP5x/pLGQeNd/FpO8NcANvhhMor7h60
BoJ7C6SqDY6aQKKsMO4wfnijj9YqI3jDkLD4FlkXwQwWuzIwi9DzZeIHwrH6VcVPXseWxSFw3u+H
ojOPvBP6JE+mbVUsVuPpX1mjO0W92wFrYnVpxHAmBiJXw06ZToygs13oiF9ZO0QjSZivehbGDFhL
v4fZAVsYnG88J4S1SkhNeuQ2WOm4eGFxrHWvCVhCqigu9EmHONu81L7OXEEFBolszfyhx0YipGu9
hQ7EMYeHdqucBiq+hY8mNRnK93YqhUTfbshjo6M7QynI7hB7q4W1efCrVixfwpM7ai1HLxiW+qpd
wuuOiI+flR3jta35NBgLMufRYvSY/sHZaLEZM0rVuoWup0sn+w7oiY4LJdrQWeRABuWLdQZgA0PO
tF+dZ2oAxcItmIEqPi99uKKg4GDgQlUoNXoDxLBOrHRluJdsvpmX7UZ+FuWt7svp/aucivF1kP1C
ha75yh3VGvxEG+lV4dbA5UtOz33u41DXR4REEx6WmVu1ynd6+twGyMS10z2bKt96TPLnIbdO3dBl
DhXAD62Mbk3zGZNPgjWCePDPa1l/ePmf+XIr+6ml0NvEAIFqL9Q+SCq9fTdtjdJ5LdMOkHK95gC7
151xM5gInAJM2HSFNwpGQTK7ZiI9K01GSjtNP6Rfe08eGjyMyACVqCxqDRDfe45w4FMm1qvNeslc
RQwqacqD9TGJ1kXi06blPqgc4m9js+43S4/XVoEHA2gAM+hEzK2/vPcWlppuYuV2Y9uavhDGRhW7
H6KJkd5xiX/p0L/GslYaw8geyvfKDf8U4eFVgfe4vqRB2WoizdzWNl8QfyMfK7Y43Vjnz4ZFLOqz
rlxZ+lWjeFk8AKMHLhCS91boyAI74iXoHtBe4BvD7fZgtaPgSHDPvT6sVdNWSWz+3zhuBnygSC+e
hcotPmgrXn//59Hw0N1fliclnTT2jE5Ysbm5BL9G/DyJljgw0d1Rvu8X4TGmvyCJ+FpMYkbOo5eW
k4vtdhqyY646r+whVSNujzNiK9p+qu6XmuW9VSnXobcmI/j8zze+k7rR+u4KsLAYLAzLoZNyrP4T
0anWf7TizuVOiILhHZgYkKEEoYOYHEmz/J1T22PX0cf7YfbAVad7ZfMZotmOP4C+S8A+zbNlRpEF
3jiqoXWu3koZUMc9FvlI5lz8/mCzhXnTaWe6R82gGLL9o7D/NTUT0KMT+gPPnt4lMtxeZd3Qc+Ad
VlkKSXJakXsQrwGuyn+6QsikN35/HUcPxefsEDQLPgedIX0Cma9tZihhD+bkWCdkTNNNai2SXRp1
8+e4f4V+uRv+Iho5WvaGwZcfDCyyJW+enDKjArwa2lfpdrXVEhjXrTHTnOGjki09lDoVYA+rKPXm
WU/8hQ1L8Rm0X+MEjSa4z5mjxdDmch6fgwkMisuyy5pJkxKOQk5daToXNHB8ODEnUevgqgwwjS0x
Uw/R6V/v4g+b63WROTu+fRDpfRitrZf7fsV95B88+JIU7F3H+w4/sG5p6sXOn61Dk46kC6xgszOU
8fU6EbCLJGwGnyGt0wsapdcBRBhYv+UG2x2g4xdAj4rvB9YbJrgyxg9mZbbdsf9DvNkenGB2Ku7U
KKKNx2bJhjlme/LNZuzI0xFPiYe/x8ZxEHF2a2KvU4V7+tA3eiNkO7ryVWqXP8AIhZ9v0VsIV6iO
VLFuKv4w2JHXl2LCvlKAmBiFRGMU6T/4ZjpStcCKtKgKuEUFh6rUjH8Flw8UQLQhSiKF/E2O0u+p
UWj5btJIvYK7jwqgzT40Z4BQZ5LZHN42fD1/zMMa51PY0g+uMtrLTXqn/hZxmZDnWHbJ3czuVWZr
El7hP8xmqSCs+DwC2EgEZJ85xWBJQN+4uOlP+eG4XRREimYA7Hh7Fj6byysbAeAuZkUpi2P52961
hhWfiTwGJ9bvdgzdmwZgvIpq7Qj9RPW/ipQIlF5aHkn/BBebmv7laaOT1qB+7hIrzZ02gCww03A7
6SmYzbIHOPOt1pYkOP5gG/Cfke8ClovOd1i/+TnWocQrxdfvWZv77YS5sCCyXHW0WXfS1s0PfXBx
MZtt/XGGYBBigz2woG5pL7FwXC1+7xXt7MszEHVAQbthyUm2HRCsL27ph95Q02wCTTbIG89KsWCL
HXGhbNebiP3cAN+OTcDSHg9+NNrffIEibyJMURSizmJt+diZky5Cp4OlXAI9VHq+2uBhm3t5jVet
y950iO3HF47+rNa+YJKjSHQME7mqw7U3TC6etwT+jtW285/vUS1G583gXoS1Dn9C47+Qdp/A5K/m
HteVFWKN5JsXgQ9AyHU5X0dE1/l8ECz+/iKaFEzRz93nGKV5NnwlIUSKsYuOOHb51d4ZREEVgFiZ
ZWOEPZfe/j7+1nmwXn2+A2MPM4/wOFifLBT/q2f0XgCNpme2VF2crGQaxtPTyorukDsSs7FOgmaS
2NL/lxiS3ay1GNi4lFEmyg80hd/0jBYJGZoPxVDME5dK7ksC6NHDOgcmLQis+BmFc8DfYisW/mbc
sxYgyN8GiTI0M9YoMIO7QE7rDPcBA1Edjobg9NVtbZEjPNadbkXbMMXlzi2F7Nm3uO26QccTdSY5
UeQZQlb4Qd9lSr99d9nwC1CKAweYc1kYZYq4HbRiXQJSbctnchyNysPheYu72vCJxeJ2oer3uAiO
gpG9temr2HGec2LYROkppeTrgAltu6fztkQFRZt3dZnewyLHUTU9k5WwzffmIy7Kiyor+DmatuhJ
1KmaxaIiznJKJAoDHJ+NLsmT3EIgMkTz6j4vH1WDLN1Puwho7Wnhkiy/+gOW9Hy4eQ6YiHtDtkJA
CIQHUpVEqsKhVa2cKV9NhOVug/gyMNQAzpBDk7lYDu4+ytGCaaG2SjJIDsT1npSagE8uFR4Lyxs0
AyAJSUu4/TxOuoentol8bEaFcZoKRupDBsWf9yXZ/j3VxLIocuPT4WVnB/u3mcxl/nnWGclZrYuB
XsLjvMrow1CRTWWj8UhafsHo//u7Tj0sIh93Q8bxk4/q9xJfNmx4DiXq/H1sB/AamfaQaoi+6Oax
c76z8o5VqvN15WKuX/JOFMjQovTRX5KfATKMg8z07YYc8WqWCwNMEpwA1u0pCDUmjNf9pkT7yc7/
sM2dnp6LQN+XJpmC1eXujh/L1N8g9g/iPpTyK7uJPiAjBjqC8+wu8gsVEbUs9w7JAkdlAPaRMDtJ
I4PtmUK7XqSM+tvrZ6kbkEQR9PE/wzOcEB1LcQM4s1Kj+lm/OVAS9aS1kCASXEnLtVrj4MQT3JKy
zuideWAIgyxwlfQeeXqQkzZXvv2HQxWZgf9ZFik8uN+1RBio32/id58K8Plsz9qtgJMxagcVbB6r
hvmTVjLt/DngyYx/63jkMDEU1WNyW38o7B8C2svuTCUZjqnvb+M6j8T315RzmOUq6ekba+lIYacB
LX4L8/CC+atflLM2hg7r+gbz8UVxc1eVnul72ntvuyphSnbwAE/q/4iSh7L8oZqTTU8B7Yd/HKa4
OCPU2dQmsEY/JWbUV7Uf+z3Oa1odoLOZAVvO/sw/5vxE+fg7aRitKbOQgNzUxhSaXymkLDDEDPEc
vyBlD7eyEfhDgxneCwzcyhDB0XsUZ/Vf5N4d9bdX9aNbzGWR486SGucdJfLeeUoq5b2f/cQ1d+DL
RK9bfbYTmyu2Gbm8vSRkP1cN3CPtU2cIsNGQMZV9KW7NP7KYDplhYM3BEaA3P4IEmk3Ro8Yujtuy
U/LiOTCsfczgZFR2HHICJufxxy/aXGZ645cQ0AqA3CMk0P/r9G6MxHBOzs/0zCjtIGRC5+GJIFPX
nA0f81Lw6RvpIS2Mvt3U270UrkE0H1fa5dt+h3AdoZy73QTzY9+nDigYuDSeg5CDiQvH3buIv3fU
yC4M/ItcVKNQHvEttm5Y9Oj/UlT1BbZZs/pXifnUuQH2Qqxmiz/m3VGHS5OJsYawtgGPSBD8rmtV
fOMalzbr93cZqZfphi2XFU/S8D38wvBULNCMDr3abGCtivXWJ36STOP4xJajmuMiZL7h1Yr55aK1
xurgOOJzsK9MBI8iVCjKDhLpUfUN8guOUGWoTF0STFkn/fgrmO26JfseC7eo10Siq2Qx6myEXLNR
baE7i7S180KIzLTyyR043wjn+HsxlL9Zly12JqLCZckWQ3uDKq3k0QO8zQYwAHAnr9MHxkbuERvy
Vc5Brwp6vGguS/0aeLVMduhUp+BivWrLTnLvINjYQ6HYV1A6n8EXw7dm+f2bfoNYzu25AZf5nYuJ
RLnRQcY2D1GanPp8Jmq7OVjmZPyXzNgeM7VjO0NRahU2Gi1hhkQWh6hObeIj/xLAweJBN9hPJtyu
51gTw8qaKsH8lb/XYYeJThWT38pb+IEjvPkrcHTzvd3rrULxwoq1c0ciUFt6P5mvUlr8tq7a0p+l
EhdMlCLPq0wO5E1JNwFKaZ5zXh+N1sliCu9XELbCZj7OXYTyDY1ZE7CC/xMp3nSa2xxwknsFPgel
D1mlueUqmN6ZkHdQTHcbgGBfEpBn0dGzIoy5e86RbWlVgvWdvmU+LU0RE13d5icDB/tW13zumBju
PCQZW8e5RtKIifbgwNgsX3drPb6qRAY/Tyeb4nWTy+bkSFISEFzZ0Gt/jzeD8gv3wPEWZInBSWR9
ixFp/wzx05Ul/IRb+8fOGJ2VR4yq4kH6/VQwwefxLM6VQJstIPY4jpxP0LZwFWQC6/KtmT87YuMf
BNL35v1gGGX/9V4blxPjw8t1QYa7gCy5AB5uVFZ41du8lrnImSLA/EIEkqGKl6asnHs7Zx9Jm7SE
ooEdhVBdGvS2Rlb5vHfScAHneevc0ekDTG+vUSNOy7vJ9dgEqdYlFGY1aCu0kw+wt5Grg+SsgkQN
PU1rTYw0w/ILUTQZ0bJtKYn7SlFiY6PPRZe0SAYcD6Y9pOmaUPnjOExFjlY+HI+R38S1pRdlNOde
G6c8eaiItPYj8+3t2ufBV/Z7xpBbFqshKOiPmjSIA3OrtDvrbTtcB9PFc9cNZKqWD8Ig+PPMvapD
3TTSHheNr/s8l1B+kMzxNF9Li32H0UVMAADHVH7Ij9/q/AFDnJ23FAOp6E733ekP9BE9BFOrV+BE
0KRTnfjfb8W9f3UkXpMfz6rAKihBsz6MJ+5TdZMEE86i1d7SUwJYi2iK/32aWIhrHe0Ezrf5GCbp
0NLAyoXatQgtXEW3DEFrnqXGhaL4EOiDBntuTedO8ZqfFB33pR0e6LDyVyU+2mSZq/kBeBWhLjvK
sfj1aMgZkSU8NMA16xVi+bEo4gRTEQjCqOGSmTQbDnbYwzodbb1u0xltEVMPvLVZo3fJsLMB2Pd6
IBHCQps51IzD8l9baRYuCoT4GSxkPWZkOCAKpULMrUGJHmPdqHZMcfqTFfyofahHVY3X5fK310mQ
oCV+EULwnCo8DOaB0Gk3i7s7L2LnFNDKQd9z7CEhUG4Iy6XLxYOS+aHkP86+LpWi/o6uXZJmOORj
caq/hYV8xr9f0x2ya4oy4StwesYwVksXYdhxJrjBYDfFTBiVaG0ad00hDM7ygWOYY39i5+qdDDAU
sS8nvjdoXQTKdxjI626ECEaxd6IkH8lZdSOAyrR86DAUteEuyw2S1zHDoN5ANMFSBjA0kMW83qRs
sDvfsdUY11L447uXYklVD2bH1HlJzuoC92NUoPRkm3fKyTFdLdOCkV/4iFStAi+Fvm5+IcZeeAOp
fWlwez9hSc3UkDlsITPywFzjyesgOew+gr8rQiw1DjqtVttquFo4bLy4vO63RvhA+fXQ6tjQhj57
oSWw9Jbukg2aqdthtJFJhDG+5FT4BRMhtwK8cLmRk1m2QxphDGvPdBnoIniwR+Agp+oeYpRnOqEF
TMfcvrfOUErSRDUUBDgCMhFxVp7rQgclV+GUQdiYssFLe3VdJqEDcr1axDKtgDWXh1XHwPqyREt4
CLVC82xUr15FsqwEJIqdFQiSvXQHFHrtpHrway3Nzjgvd0m0w3p0CXb3xDIb3QH3Qyagq6NZZokS
Euw8BlFu/+jN9KhyzOJGUiZpHvcnm4ob6E2kmelG0jXzustIJ3IA9TreGqT07jpcYKFufLRIVc4s
g1N06V74B1XVPyKJQJ12QF/FxBrmM995RhyLH52gGqq8uXE/2xPoxX3hsA/sJg4PmXcjnjsx49MO
mityQQ2pAX7Qi0BuTQNzizkMoMaVjXZwFKqyWVe0hOj/VQoXTWg5OGZ3Pv28WNbNdVmNyqRtpRep
4+HwecnpGGoQfaLwL1KnZ+uxea4zP0nm2DDcQaC05dDp6UCtHfKByQOLByrwvGiK71mjYfZ0LYDE
Kss5au65PN/CAdEt1trRAwL57/MENxwsIjX+u7ucfDi5lIrKviu6TjYRabdaiZfNtDpSlQ89RVz8
YFO4Ayy+ifPBfziSIDJrYJtNwwLN1gV653x+t+OlzojcAx4xCJK4GyVwH/dWjCIQpImscgVf7zfS
pC/C8lOi6lyPSF0v+rzE5ywc/lUHyGNyS/GCMr2Z5QtblPN4u9Q2TzIlxvpES6thERFqEJ2ppoec
fAzIyh8zBe+GhJxVIwhfKBZwR+H8tZ5gv4nxGJl1qhu+txXdyXv16Czm9tFa7t7NM8/hoSt0Or5J
ekFZnCOjSwx7Kv6mnGOB0SdIr/mtoEevLV7l1kArHjKCQAseA2kZsM1rZb/POhU4OrsxZ76Wf50q
NMAKS0F6bnU5ztE5QqCXWTzhd7m8TtGzggMJCL1SkfefGXQMqJ4QUKg2noUfEOHq1qkXdWATJblz
sBjwO7lOhDeT7lHT6c3BOlIS17jbwuKdWIfG39BRoKqvYwlpBR5OvmW8P0oylX6Z0LrG+7qRD119
5rvf5XSMIWUNWxUBKYl+1Bj7HKJD5jQB7vE4EgK8Hm24iVRxFn2EulV4lgpua51F1X/AzjID1NG+
6+v2YFYNbdMYKUfi8dCe8URfmE9Ois+wyrgFQ7JGMHsuynwNmwmAg1a99L07yfS346Zj6KuKVE9u
WlE0lTcsZWhffNWnDxGzRbPny5FifPj9peqHUheFfP0kPSmx8gE2OVVlceBDV3/Gxifv23R1XRep
UKbNHXiLDqOr0koOG3SyVSH5t+8/Twc3vTEWc5lDVSpv9CcGh9KuMYFW1+OydtOKnmncOK5iZisv
WqOFMsFtMIfh0KqsZmUu8k/kcNv4bVf0dLRaOHptWSvFbevBTo45l4cI8WQT07QZ4NflwZDSHzaQ
Qz7XzAgMLpbvavDy5Z8RBhISpTKlZStNplT7f80uG4asxoGdQ+C1DKQDvUbX3xHvzzGfkHe9dmKv
YJjj64vB7IEeFeLGbFVIbq+TzyuWNDwjkPlAJmHQtKhThbbUZA4dSlguQbqOyh6hU3p0iR32a/O0
KMqPP2vQd4mTgbY1YVR7WS8QiqBxLVaSn4eO+RAE3QVfFcUPi4bYDF5pTIz6bMEF0Ie4MXR3WoJr
+ou7EtvUvwe9BouKR6L7FXkUkyC1DEeIrLedVJb207jn8iQeaOvCgIoHO/IDlEwAuTt668F6BmyB
3B+HqjxGKCEZms6MN/3Ej9qV8dPwLiQVGBRN9ndK93B+41+Q7wDRvsdWK8mbYR9pkptQR/mrLaYK
GXixEuZw9nKa8zjVIsoxkH4ezLmNLCOZYGu2fqYl4W1Ge5mwb4MaEAFHZBhO34zeQv7m5f73nH9U
pRMI/pvpHwZImKqpAQgYvfOu6yTNJmdPlWa4NnRWJAxrSqnCes4kcHkcKDvMPK9S8Qq+72p6vhSG
xQ1bAi47nlv8fqkua5UpQMqLEAXoqxjZ7BYDqFdXWUM3MoC1UxpyodrHKA2W455BAoWbr62ZIEIe
afjWF/jVfsmnG3xLwvsmR9OgriyBpaaDS9tEQThXel/RWaqB/GZnaRj5L3/g3wpoMETAh7oWZboL
KlcvmUZ44aSDW+XEF+W3v93eV0TVNCrhB/qG+4xC3x/V2w+R52oj0oyh2PMLJy/oKrkAfd5/+Mwi
HjTCnayYJqPC5zRORQieq+WLav6f7MFpj3I3r639Dd7mAjlxjjA6lO3/zsPM4aMo8GN0Nd0NXWaT
whxtV4t7z4lPT5wKQcLKDp3czl4674noDJA0qB/jFiKnxlC5FG+gsILni0H/EYVarRrAv+mhXs3Z
wbLTN+hi4aOQnAL4Okb4g/ukiy92xJRKfhL+zQhq5089lA5DVGF5SRMpqOVuJ4gRQ020E/ddgTvN
0Wo8Un00AgQPWn5uI7vo459NZ4qbsF15iz+449rfrcAZZ+C95NnNTjerwpkFan4jljaWnmJyDyHC
bnnLnu3Ir6KHK/9DuVXSIqkDHoc+zrM4mo9cXIX5hgBEtIh8xUyvQ4QA7AfZi8FDY39Rm5GYfvtp
zn25LSoqd1uzKP0dsIK7KJRDd+2lalI8OXvc/rNzRsIK5mUfomNJiDjaGWqGjiWqBp2nfaSuHy+0
SzGOIj4Ok15WwQY55w1iDPzQ+FUEgiRnY2nm01Hkbo2Z4Es3sZoqD0RcPchKgkqIlrlwt4//+Z27
nwi8ryFjv6fv0CzDjGCfB0xRtC9egtJ6owa/8dBkJtliQ7DV1K5W4NDlOO50Gj7TYZKca/twP1Qm
KUiqGxF7x5noKZuW13qvLH+hSwbMNERRRcCzr/wvMFkxl1azCYoUg97OxjOMNh0QkjbwZ6lWiHlU
KGnM8TpoKlPoi2dQ25D4VqrC6RJ0eb3rz7pOnvN+xwrYqrLD/rOIlkJsmicCqV03g5oc/z4aR8FG
erYjOjIWBomIMkHGf04H9a0puHNCX2Zfg2l8cnWkKtuDWusHT5jZJCGjt6siet7GmFhwJPusVmoc
xkhY3M69IwcrReHW5B2DL5CfEb0xBCj9C6WctEPalthCHEZa+FjJ8LLXYP3GLnnCEXFim/N4sxBK
IXxXupvRMss6fIRi5zP8DZYl9Vg+osSwflatjCqrdXNoRdEhm73LgxuBnH9J8AAJH2PhSLu/xZQz
N8EVkhR/++M8P1S+PPnABm/BeqeYC9OMvu9CaPOSnKvwQytC7vJ6m4Wa28hUmmoA6dYNrEnVHwO9
dpx4oL6mVgSV30LLYJydleLE4pxHfo9W7dlhGslYWseaSWumpqkvD3K6LIM1zR6lKUT29pMT1Y1a
otKyiH9PSoCHkyvKQjAN8VMBQcb0IEC+lFzib4tIIOqcjIwA5t4THibs2e9GWCVahSkZCwCCyqnD
30LkV1gH27khhuILESl9Muv6U/BZUOKCp0S4/5Mxw08uNrkzYhshPSizVZE6k1LLLfX5UyTwAiei
YwLohevnxZ7D8Su1qgqILQvO4jSc4mChpFQYjimyOTuDo//8RlpcIRAm9Aa853qMLR8QP5tMH1im
tVEcwQVX0KySCPDjsUpJSxFk5y2KH3Dw0L8bfh9qo0rtcb/0Z3hIy7l07rPR96Ui4RZKQIhBb3b2
x6BgXhOSK4Wqxz5zB2mBr6fZJibMrVGi/tLz4SPKJ8Kdk3AlA5jmx87xxntPNgeN3Now6+1f15WR
j355EmPqbKu2xary6+9oJrajUonVhcmqRGag7FyQGyiJAKTAktpcUhUZQ3dBASd3FSmjCrHVw7A1
z7t3lb9aAMsHhBfl2NNEIFhoRNSLLbhvyBeaMOMxKQhsTBtNaLomr+if5P0fBs9wcnwvf4DG3Qyz
9pVPtCu3zIrrJqebceHLuO5suOQz0HH5pHyXKy2TyouIA+8VjnF6BURPdYCSiArTzsMwEVs9XYaY
yt0Jw+BNKDOY4SJZEqt9CScwfcFAIrOGYCAS0jmwrLEb27biEVI1mvSNj/coj8BK7xjhgSvLowC3
pr9V6uaivvz0vmbyvaWYNv+RD2MiNeyN1RC2Ha4VyoL9aMm/+fzugstK0xSGp6ePtu9n7Xl45YcL
/cEIzpwpzfiModXtKVJ8s6kq2IWybGJD8eOFmBnSxUULUBj0YBxv9pcWu2lQMFpFS8j3FhzuBUuw
SfGmKqlNIiVu4f3wyB7S/YuQGv8OuScqAn91d90YADgvEX3OEF6bYWBeJzWJl0DVoJmWKSeVgQEv
0Orwo050CmBfdfY0CMe1yy+GgJUv+Or5VAagT+Lvy5Yj8kwdI20srYVg4YlN9muBOca8G6kIxcx2
U0vnHThn/M1jqswWm+MIsDzX+1v1TywroIfAEre0W/Ean9W3yUCmJpnQQ3zKOCtkfjhZM+f75xRb
SNNmL5DRC5i67rGkQX3czs1zzkGl+GnWWsvzGC7iC2N4ZHl8KkSkdQveveIxf2KNxfEGRltsIg5V
nMlClQ76Th5paoQTZIf4ouMC/+YwVQkGvhFUn8fRNZlY3me7aAnS4hnHDQr5QzTgfUbSVKpPzOcc
NRvH6pDBpeBhTWMdFT6d0QyKmjCEZuaE67FLX+UnaNcuBkW3chzooYhDZmCdHN/lNQo6o+iI1fuQ
Iw2dOp7HNu2pW+0+GWYxQjWi8BpS25W0O5ti9TdqOUm0Mku5wuVj5TVGBlKk6TZ+ycA1kjOI1YLJ
EPVcwZIt/qTxKpyq7Qm6Ohk4LE3fv5yYdcMz4mhXMr7WKE5MYtK/9SxNZFsRTFbZqOZYpbn01O2E
tXZe33uFTco9no7A2rqrrk5en/XLQzZLwXwYEuqXsMOGdLGQQhPs82aXAVd5ug4tcuyPfHTvUx1u
zF4lb8wJ5GScWj/rlqff/TzY4pwSekrGoSzBb94H67qHc2XGY618nOopz1uXT9gk3pt0bMc/3ygJ
scgyy35V7iH0h1ZeOuYAPF8RT1NrZE3fjisKHg1pmJesAC+9xISlBxyLE6GSlIJi3PgqTeaKQSuU
1hSf+TjouSX5nS3ypBmp967jb+PYUlvf6Ytb1H8URC0P/nNrrA5/n1GenCrwDGkLsa3uLwazegaB
bhQi1/D8E/vzQiRDbHtFgh3u+/pYAVKqvxzzNNC0FCj4pSAEy5QwVXvVe4u1RySTzRTC3QiXilK0
dd660YHd2ykDBuekb1a3t4Hkw1l/X3VdPnj/U40lLiZ+wR+hhT+wSn8NxXoWb3Jlf2baT5xFOukt
zBrVm1jtt3+TSJKlhe+lkNVTSTDEGe5FmIwOKjoxrOHwmMMaUweD1/1lVKy5UI3yVFDBQq1TBRTv
K7z/Yh5ZAqCLQsQ+GxGomiD5grJvZGV2PT4Kdjlmp4OtnheAgvV4v1Q1fcWjLrCzbyjkHD58vHkk
lEe+Z1GjMRxn5OJ1E8acfvw6xHorQdQ44kj8PBa96jUzYBCOYqZMoYuMchFuYE3h1F/EzWmf3xZE
+/1X90yyZ70H/GgioD6KfoISRPgUW9EvdKZmoolSEM8n3TsUJGgfqDtUkkEpULldSzyuCywACg4M
Y5vlk/QWAz7ciquoKw2W7NC36nwmPa2dINIMfFML9Pq/+1NaaVktAuvZ6ovW9QWfaAkrXGVURe+2
EKsAQO/cGteCh44jzJB+GQkhV7wGsH3cM/rAa/VkYlzoFuW8IumioN3kUsHYsUv+oOj3QlAYXd3R
NVbXRterGLGLHS+C71+XQW5pYB7b2pWqFobNXhjV8mpWYi8l6p28Y38C3MPCejHS65qM/kusWKxh
n9N3fM66AK4yCpwgSqNi5BOVYSWHl1Dfvbg5lb8M3t5BPfJW7PHqnkCh1manaNMdqXs3xMfuIiU3
h59BbhapohcYml7LIcrZWOavs9w4TTn4cHLCUtGJtKC1cQX87JFNorGY8anEWheoSkEkcj1Px9Bs
D+ExbhbROyKQieNe5yZRG5yp1nKONZkxqIz457kF8wpqD7AG9KM0no3QcoSYVB37BlJdd/On4NQF
jNY8sFwFdy+kaPHfm+V1pNxIKyUDL7AejH6JOmnMfSw9cxRvDH/U5jOPx8XH2BHCMDe3c4kZ+Gro
+i7TK7WaiqPGM+zfB50G1vFyiw86JAIi95IXukPN3cYdDSTFhCYx+2l4vLj8gOYGf+yU712K8Ic4
1s7BFipVCtkYUsKRxGIL9WlP7Un/xmSI88LS0uvcHsvx1EH79lGlcz84urodyrud/8JUKcVqwdyP
L//ipvXE5LtAMn1r1nR8XDQRhqIf9X55MHVbfE86UbzvY6xhS2O4DULHkIrSZH6Wcef4irqBuOWa
imYg3fF7C9/kxYBqE1lVZv8/TNNaZYtAjd47wrzp/QcNr8CG2bOnnD660aY8VhBq9wBBPF2dGnI7
HcwrPWuqTGL3NewXDN96cCZF0Gm9vBNjhsVvY/sr6LCv5cXpTk4c+Ppy5WUdZ8ZqyEkexX/fUdyf
MydbnjESfxjpK77F0W2fRY4HuA9QolBk8BU+tdx0iF0yylBmsNLCYr3YQnEUTM0nJ+O15Nhx+QBN
8TJHU6ETbU7KGiM3/cBEtPhk2yJA6r5of4lv42KBkKasfXfEEGRboZGpJTPWDivhuZfg1DuoLXmB
DdaNgNVKxFP2UYO3o4kuBCrhXHXhxxtBqNxa84FnXTZDg38oZk578MF0OtYRiLEBmvq6jz4NHPUe
mQ9M7GWcbC4DuWcaUt9cJgQtD0vlatRtG1rnu/5PhYwfZi7rIkrpGBcn46oFZVsGLgqZx03VkaSf
4LEEpd8iMEegvX0IoB0Vx9M1QVx+/FaVY0nz08XZ/jqKxCSrF7doRO02T3pMN6N0A1Uj7x28mgL5
CjPE9bNr/K2j5djbugnuL/tf2HpWj9b/SO1DlAUmHjVT+SgAR6W0DTuEHQV2JViJhvE7sKlpDhXB
q7flxSxdDHEQ64gejDT4BJti23Ej3bZVTLEVaT6bZTjHG612TUK9CxLe5Y3M3p8Ue2lQ37ydR2SS
Vly5dIvcEYAxMhnjMcOwgDduKI1yaXO+/TWc1VdLeSeXnEwZuP1pFbM2y2WFIqB3Sk/Mhqcd9YQ3
E2qPlx+RtTRxhX644JJxMiDisJokzuFlcF4S8t1r2IlbZ7UpTqrMGgMEkBY5xt4Acec7eVQvSjPX
aV/FQb1hQ+/nLOVeKB8yWszCarpd+VV2WnRnsZ17Dw/hOnOZzG6yxvJk9d6ucZ+oyTOBAc8mLqxh
ac6cTulacivMq93gz1JUcGDaxgIRmXUHVZ63u4125T+jftoiVO/Abl4NQKEa3JO0j84BiVbw7+hC
+9FTLpbrTuHZZoxjpkQILFjeWLUHtzzjYhckRKJqkDShZ7U97NmJF9qCiquHCDIXbpPg4lXj/pr3
WmKOmbBYxuUjcHuFT9/m7xaGIpsv+PwrMoyG019txntwRUvdY29EKD8b+h3/EApUogkkB+Tw8h2K
TpCWD24XwoXvRxxkQ9Tfdm5ri3mMCBKrgUb1VLdKgVxFlJ2CnhPGMVJtG3Vs5+TP6H3dijHQ/8ys
gOuvugBfnt2LgO3AbrprZ6QCXf3N5LE8dMYhLxpDyoR3c3XciLGGL93sE4h0358z1ao2V89UTllr
7+vloo1w0YHqtWM09SF6LoeEtSRkS4vWVUVppFKvJpWr2oqQernzCcH5F3T4qkTdM6Im884SrypG
wTO++XFP/rHwMMoN7fA03M3ifJRxGq0IM8dX8brAyVVfdPVB+LBlgY+y0U/hlPDRIOTr2ZcEl4f+
rUi0SvYFNVnbDpTRbH0WHEw8VwNhu9cukau7SNf9ysg7apcbaLm+w5/QDM3byX4x4n5MgrvPh4H8
y2wBI4wPiP6bxKe8PWguYVxRpYMjDRnOV0hU+UnQi/2w4FAbpxj+Nkf2ZJbyfwD390nGYuhrQ/8f
54ZrJOuduRTS+1CAYvHpeH8R0pKakO2TB+qsR8CgwIwaVfg5WepG2iUEdGJBjYlJYtF2MVk+wt8U
Mm7nIBJdLX3rE2xL/W3WpBmz7EMMQVstHY9JU/ehH9Hj/KcIwPZ15Tls6OMrvrEwJzIA2J5Aq7gf
xK96svOs66d0KD7iKPTPmlDkcMmfNXYWbEXs+dKLEjt6yrBpuHwplr5Ajdsotv0xrGhN+zZNGyQA
+sDHj5xQW7F8xWULfy8qM+B1m/ezkp+IO2EkuFNaEmoF/k+MTGgKeUgFiVlYQyrETfYZhJvJ7jzK
N+vTsi+HqDdCkkbZBd76ICFYqbFwUjeHGY8PhJTF2H/7B/3gMno7/SlCb7QIdv/h8T2oz8j6rHoZ
kMGLxAosHsktGXBoOqvHJp3u8pmkj7ZIypYvbdOLjd0nag/QODKHu2Jsz+QpTn5q8ttSopdMVsQ9
m+TogyDT0qYnvNUi32/TzLYkNnV5g68k+qwHghfext1T1bFyC2E7H4778xvaJcldzhBTa0XlyYfw
k77bn71DsuxXazPVopEMPZJgHko4tB1OTy4J69GG584T0fZx58JlOscHFxxRWcZb1gVhyd1r1862
+dR4pWXVF4VBUIFqw2Y/JebAiiqFD/iJx8Il/jiaP7Yes8JYY/s+r+U6CoJZ9qGOebIbQAOzsCvT
LeWpbAjiTzqnpWbpMu+cuSMl4FwzsceE6ugJ7OUq7j1jqd/2FYe70PQhvB1UCiTIvf5wuredkJcc
0P3x52JRHaeDLc6o81+nZ0/KXCV+GOBv6LiYriR8yRGO+SYrexT6uOWHZXPvoNoSMOYQ5BjkyM1z
PEUQcKeNSoNJY07gY4f0gZOWXQUoSU2LxBY9ZzKxCF9a+Afp1hJv419P2H7wY1kalsg6Vwg4X2kI
1wUKNpPT+xYtaZvWPh4zp0V14lPhyIVV1nWKOdyijIH1Zkaa/dlJzjJYRjepGkSdR0Wut7F3YeNF
vCF8IOryGUuAahEYofOsSXCn4BamsaA+UvBfIxg+EkS+y0FuMVVBz3JWaE0D5FU04g/lvEDMLcj1
R2qkGBVSbZtxm/anh8sOEoUnUCpPKvL9z75k/LT9zVw6jyFh4WNkz4Cg8Qb1elea0dOxgEj+Xhj+
nu8/FxxJCamaZQw4PHBNtJzJGlQZHOfbz1T73IKkRVrs4hEsOVsO2LOedjT/LEQwQBHnCUmREBLj
050m9kMnGNwSog0AL8VyVM1BVzpoyCyhoP4pXibmCocglMdQaaOVQG2WzA7HIwp2T2P42ptFc/sc
UYLp5wlbw/cl5JLv5PSKjA8DpGEA+Hx7DE3BqzwNCTM716ZFlwex/taZNNxD/3j0WEWt6/8ETZFS
hBjtgXy1kF8WkHUG2lsOHqUAOw5fbViZyKFlaEhC8dwi/E+a6/oRafcU/VaWjFBNPMQjMLV/mvpq
0pDycR7u0GfVKUHY2rXfAfpbDl9BQZGvL0kq0P+iRNtIHhVD7TxT6ZAllsVllo/Ka2ZRRTLlB56e
Hw3xLAw+7O6pjNIkZ6jjalSBy7o3IbCBb/tMjEHZ4gy5vnxrGq5YDNN3T2FiPKbUae7pCu2d1/oH
1+nTKLbaU3rKUyVG8c949ONPGPPq8yIuWE2d3jJc3E9yeVaXp10WrDHra/IUxZT3OYlsTNFfarkx
LFHCottjxrEgpPSj1U0xdvP8l9c7kRMSuczvoRXNtL87o89N73YVOeqMViORWApkqspee5akTFjF
hsvdOxmAOV74yEMx9il/SKy00hi2AD95HVXynlnl8hW05FSMIRfBFNSlTlunxUrm6Cd7PjPkV/dS
6gwpDzOI2eBay5s7GE58ciZOqZeNMiQi41zNQXcifKnpItkiuN+YC2v1RXx8b4KurZ2yJcMsXLjW
Zdx0YeNFlY2bqKVLLSEKu3zyL6c1foObgN0hYwgmfiBrKNfLVtO2J0tCPfCf5LDGRwC7isq1OO7f
U/20FhrCvnAUBRV8Z9U+WKVt1A4k8Lv27/O3eNnHgXlx2FhysEPTIAEnLIhzedkGwFASNTI1VGq1
anxxi6fJVv3ZGviKOvL3pco1cmEd7l2UZgehmlE87ojRk7Vqz4Gf0ANdM/6xJYxJHSXchfVyaPcC
MT/BmZ04oMPATRnsbA0rUeBsRWt85WcBoUY5nuRuXPTwm1UIukpDwqGW/L7+NvtusBnR2iFXwL3E
R27paOcEqw7QvupEi8TEcfCSzBOkCoIPrFwpOwL0t/r/xtOGTohjTNhjCN4DGLHdETIP4zscU4bA
w+AJ/YGBf7ONbHLoOWXTDs6HdoEvVgxOA95YRAyt3WYDvpBkvmAR9Ro/XZRhxqHDEWhJHosOI+QC
DB5AQYPMJxZjALw52Kfeys49v/v3ccI7aCLrn7RWYe+aLIIDA6i+pCgFi5+Nyqucum8vDG2pWMmr
Hq4agu5UJrSzNNVWsqUqWoGFlcMW6+4Uq8CwzQRNxr1Bu56xujpycZ1nJgyi+DQNCOlKU43wOE+u
jBo5pSzVj4ROa35R9sBRG8tgP3HAi6UIWHm9w7kRyRbjJFWqVPYdW4jHj56F0777AHkF7WHpRQVL
6B4a+jqkOTmwlQpEiYL531n4D+4oJ//6+TdY2ACmaqTJsevp0FsaHLPnAG8aHpG5SSlU0DXj1acE
3b1wzUWCuKOCLWGl1A07PiopNANySwvfcw6x79ekNVJHsFgqG1kEUl7NfbUsc4RnrPX9rywt8VjL
k4YXqCIky3oogg5K0VlSXyG9zDLRqSBGHS2ZwP8LR6qckU1vwnwEANdXyml1PWWGFKXGHIf5Y/L6
eCLQeF+ZOGV83NOF/fVoq+u4jri4g15thP97PIJXsKXswoN0ljvEWtMdx4YXTHX2oo4xGQ4SQjl0
cOOz/VOcrYs1Rc73NVz468GVxkT2WgQxVCf0mz/MAC2EbYZWhqdqD7WNsgKpvs/Dys9Mzahsr3aF
lpVT3S8jTwc++YMHtWeR6O95tmZSK0ifS8pCw1qMi+lUTjTEXV64waDG7zt8ylgWUJV/O7VwE8A+
0RCaDQrvz/AFPxmSMFwXmCSzMrMGeQn6RceNX9dnVUhSpDMXe8nP1cD0Ypg9DGJcbhtZyEWYrE3r
adHVj0UOCr3VvLkgJ/jFRyTv2Eesi09+JBfghbs6EPkIEbBHjMwL2mWBj8Ga/0fxjtTdiHAGprHM
yaFXDAiKe4Oh2MJmWzt+YkelRsIuDjQ3HuVnuHDm3ILDh4Pqe2wu3VX17lFj1trf5La7EpXwavwS
WPcxA2ATECt0RnOK+t3lJxUWj94siJwEQ7aB9yVtLMoV8SCrwcES1QIiogQbbD1L/NRiWQm5R0v6
roKLxk2kAUz+KUTBQUee7XcNfHNEb1led4eU23T+Dgev+gHHPB+OsZWphLsghXaLLzwPV6Qu/MUC
2E9+6WKguqZJ8bbuu2GN77NBx1xQ97hZ25pp29D1QY3lb+31BRmF9YW3ldrP1YFodMrWuR37huel
snMnvQmnOmMYEdwVJSSpUuCxded5T6/Y6vri0rYUQRmK1YQ+J6M3zY8GobW5vPyqtG38nRris9XH
JEuoR2Gf8ABSe52Pm5mmHKjUHIeld8+KpxGBo07/keQf7lEDqmN3Ceg+mgiPBxAGam6y/xWCryDh
COwiWvqFFy8/xuC8+kTR4yB3g/ljzG8fcyGRihdaIhxdZRivmLOj9X4NC1RIQTtHgEoDJJZr51pK
/AgkVZI99WmYqby6K4HOOsH5mArpIxlBNqSjv2dt+IPcvE3vA0LdYdtdVQ8PxRJJX+lrBKW1WP45
Hj10dXrRZP8YWQcQKriebJVe1xnvItpA3FWXI15a8LlecqXgPD3SaokNIKjxw3KzErkTJZ1PY0xL
ZTP57AoIfx4h4zFuAs0w5C3b1y/eJnDr+kcZgOmOGHOXIeM99izDxkOcWrVqeSuxN9uf9PsKMLcP
zVNQE8wr53WjHcKpOw634o5f7LdRIkJw11c86Yau2GO9BEo5zqe+m4ancij1RUt/1dF8w8eEmR1g
tpCw6gPUbpW01AeMJWqJR7jAGaaFKLpk9VQqyZ6r9d7nThTYBACMYTqR06XYjlFmQYVWgHVTNLar
GfRSZSVg2OwrbHIS0pGJsCEHgJ+aFgohHfpmP3+rptxjocN6JUpiibkf+I6KrXlsYQUc72i0MC4v
ZtWX9K+s7aI7SkwPAEvshrpDmpoxruWo6tY00U4jSv9dX5QKvj4X7fNCLU/yD1oF88qBg0YT/SI1
W32IJWBI8NesuscIHZVRyG2xLeIgM3OZqbodgqDDcCLkg8elH+FMk1bibVTANM9QecuBE8Q3HU5W
SDc7RZDZAkay+TKgDP/MI3rqQzIQipAhyhrFmi/y1CZnzYSuJMeTz9URR5hrypPpkb1S9TN/ulIW
uGlX3Bc40qbLYwrB2QsLIkhQrvTeplAQg/UdnlZ0uDKb33zeW0oSlpdOh8WgJVPl+e1BQ1ZvYq+U
Wu1NAHQNE8RBy/wgEDI8RjZDVHqCymrq4++/eQ0nq4SHslKTTX3863Wd0cnCyZLFuzjfz3hLjjCv
c4GX07t9bMFwsLM/Z30XQuNDpfYqi8at5tYjEJ9CNpEe/llg6BROK8OQyybq3pM8t4pADG5LtzTw
nvz5S9zDgcXyYbu6q2kcGlxnuO5CXDfm5HbQEgClGB7yrFSrODdbdz+EBZhGql/Q8SEbrLvVd0Bh
keJ0ITQSS8bfh8HxopWvstXqKsdK0ZoR0DwYPnCfayhvBEvI2XSf/F3Tevw4YFau9OvDpUEA0tLF
1OIWxdVNS1M3qjqgCQChaeqjP/LZL/yi6OZnu5q3smBSP15zl/nqoSxVX/LPRuvtGmafNBCHCsGS
zzHUTd4hqnaJGNT6+05d63RHWddqXMH+xI5AY1AGuMrn8LyKH3eOLTn5T0+4UuvpZw5cayfREa9r
0ay1fkqMMnlg/3SfYXqTXfsejNYVPEi5O4jmglVyIJ16dEN6hRPO/Id08WHkzCgxPkuzPndBIeA6
bsgI/vF7cYVk4/NoMIivU/GwaSoZVadFgjF1WwXTe5Y39JVbVrnGpU04hY0ipPT25+iIVVwdnO/z
aD7QdUnycfc7lv8Xbfhn/iQy+S/Kohp7GygzKgi7WgtzB+T+9bO5vKWW5O68LrLW7WAsl9eapNZS
ccWPyhtwID/b0/Z0lRlvmgv5dNM616YBodhyk0MNRdPqBoM996jgQ6nMSH3JSAhjs9erOpbiK/5n
JMEwCsuBSPu8+lO4gHpoEPEkK7pgv2PGCMSHDF7TVo6QTuDgcjrqlEyUc89gGEBY474iSifurzd8
/WPjre3qeubTuMbi+/BTDZ5Lrg4y7wIu9y9XnTsf3dUYLWdCOOU0jjpF6mVYsFjQc4YwzNBgpqJR
d0uh7BLt5g3yIeyIkviODQ7mAw3TY1G8yoDc8TNc53WJuibEt5mJ3ODJRLqundiZd04C0o1S3J55
WoY9AEkghLfV0RTvuUQH1R6W2SLCOCl6w01zoB3V0XlNXAEeWUAKFcj2EbpAx7/Ttrkdo8LFUzfH
u//WILMOg2HaJhb1wy+JRPgraDXhBJuh0LBAJLckzCd/Gb+m1640nu/9eqBsIZzuQfh0nMfYHyno
+MfIy8OCNGl9EN6zIkgT/F8C755/JgTIm39gI/ueWqjJsQv7E1RlhJp/IldRI6f9DcdamioTaCmK
jV5sxNJUGHQ14Y5chthQMdS5AR2/s8a65mths6iDHS4jS6d73NsNn7WsxWnVS8V6iiSrpJWJLgvj
Z11MWX/I+fAPIyIwwQELxbfBjuHW+bWq41GJo2/FT3Z14YK3GD+SU/F7/9eDZzReuUwdhiUSMUj5
hcLAo9Rn0m2Cgr1fSS1JciMgPi6GP4VnSYo7aRJdENS7itvd9OkCp/n6oI+/QST4UzQ6Y9SnUS+K
XZoUknrmnTV02QVm5awFtwLpSktBakeVmv9NZrhcN0HoONdup4jv9S+sIn+8n1MepqhY4pCZu6A/
rn7KIB0St+jkHlcSrO2SfTbm77xnejsFJnGZVmTDxm3P13RCoCkNAyX9vX733z3rQng5EnXLhPwo
gzUt0mpKMJhYlNK591YNr/k6PJE8rbwsZ/XN0xZbDTHbgjyuOjpMa+psXXOtIb9HPNct/rBBKcR4
/g3Q7B2lCy4TVIoRnfhLSDZj55UtlnN0UBxmJZs8wyUGIazTDA9d1CrQKBaiVEIzp7yzN37oIkYE
XJCrw+Q1n/fljopS6rmgW8Kz8VwI+pVqNpTG8q7QsWzPSxEsCbl44cCF5A/gQOH1dr+HuwidVcLj
DLscGax9TgbbNYF05SGyo0aQ4imEpIrrighM1IX37eXCxTq65u5JrLIk8UTVd84RAUS203h3Iofr
nIqhvUtMcfFsoM1nmxo1Yp6GwOn3nTLZPsRz3XMrbkSfHP2q/fsiJDM4WGXgS4lVUX9inoUYphQi
SuDTRMe7h6PXcn5pyaQzQbNWVili0ne5RmCPDt1lfWSryGXhsSdhVCZdHQmn5sFJVEZhSNCgJguX
KS7DN1AtZj0iVBWw/H/gxta6xhk21Rh5Jhrqhu+btnpholXtcDuQgiBT4oCHpxlgsVDv8veNAX1Z
w3fdJOvNfTTouFfLQEObhuncsoZ+dUm5y56V6wKhrmGbjLYG3S4Qk0CHLFG4YZyExwMa5rhdrPNB
4B3YwyLJ6DTNbdGzVZcxt457xpC1d9+bKu/VC9Vo1MbJGPCYxOTd5zq8CSCVc1aO843j0sazXqia
wnyUuLRfHAGRe2Tvl6lAIZp4Z7751kYzaS0VmkYGMosEg7SkE6mkysPe9FmSpWr/b6cNxO8dLgrT
sYe9U43Alj6m610dD32vFMCPR9EvbYndlUNIa9HD2g3KlWcV/uqp5xu0cIlgptQZ4fnCzqVTZTyQ
0d+O57iWKSKokCrnq+sqIERT2KpSFStaqvOdl6VYprbhhwAiH8jv4SkefCq7IIe0YfDlBbHzKrq0
pNRQT+QAdAuaKUnyCUm4jITolv7A8pv/k8Q/doOT26jRNbYiEYomfIySXjj6npIhN0pHeqpfnfX6
IE5ppS3YDcxfWy17Wh+wFjmIWpnCFca4mu2mp7aYSYigLArrHe/Dw8LmNrxQbfVsptZ77rtBVZYy
r5gmuXp2HUxrRSpxW+bLjLci7M3R0ik5RS7pDZAx7OfeoTOBb5ER0wO9nzK3KrAWIgf8KrzJIpTU
shqr8SMXmxE/E4kgcPakqNgmlj1KJl2rtB+8udRafvzF79tIlkIBrpURedWMy2ophMhXZAo5gDYw
FI0uKsH2eHgXnHlqbNXJ2j8ycqfo7ucJXjQDoJ3Xc+RezbnSJvHDf68KeKjcVspuon50+OFyPTD+
HGs7Ob/LCgmAMnKHG7/OU295Bci825kJSWpcMDownphtQf6zHzBcZ/P7bngIdF6x1h9bflcMjICx
tnVA1gF9Fmip5sV5otekt14nEun5MyxYvy33Ip4y1keAiKMTvxnzCS1P+6w/WalVbCWUhwn7YwK/
hNdRpyMNeYoaCShDQesPPKF+NC3AfbeAT4vvd+YAiLlhNl23cj6pcFB/uq3YU2aO44ZIXJwuD6XL
FZ5sD7HLTp17htD6bizABvs6wkBl+v2KeV/7k3VvREJKBkz+7bFU+WUtRN7WcpBZ/1ajkv2i0hh3
J5Vef66ir2dUIP7Pev3T156XXz3/svE+mFmDdrUamEao694ecogq/szoyJA92rZDq4wkSOLoHnff
AQwGlGLqvNDyJLR1Ab+19TmrL7a5czPYOkIDuRFC6t6QquxOdyP6OZomCY+ol+WCS70cBJP4vwkl
HNI04yneoi+Gl5n8i5GiU6GXym+9VEeBByNYVrcw2uGPiw9e1wlk8j4vQhrrem62+0D/bL5xZTrr
b+TvngeRPnwEJMRqoZRg0bzRcTbengat42qAwaUnR++9w12HfHKm8VZnoqaIZ+0f2A5BZYPSyaX9
7kCANuBLjEzVvzy04UM36ByC6+ErBlBMnl2Rus6Z+C5r9NGf56a/d0fOZJC1FnqgN/QqxJawGKOr
DsDJtJkPfQ7R6uF0V14rRpGW2IHj9vlRIIGtViv4zwGEJqAqzhhB+YByNwQOoFfG1Ez1h+Dgl7aO
Ct/6Z/w+k//r7QH33cQSYHjUSGfQB33FOUOM2+eH8g6jz/XQ9+56ssbenRVTrY3Hg0tLj14ClVAB
2TUA4jLIoJyPFva7SHEO6qkjRtgT2XftMsIdAQyYxMxKWaSr47015xcwuxAhWEnP8zmxPhN6lJdR
hg3LHi5XqIlbN6RABMD7mHqT+PH/WoT+1EDaGzqSfuB11Hic4zh3LURGF/NL59+YoAzy03WAraU9
/GRzm7BlAoL+0vBK1EK4ehOxsWiNo5FmNC2qAqyEXfujL3fimReqivRVH3sCLfwlRwnLFg6E2DTB
SlGYCmLu1vlJ1bQxZAIrwQfLH6PTfvhWbVgi9vHR3HmjVbZQEvu3HRVlFzECyGP4PtZcjmjHEew4
JnWQMSspTvB573V7XOgWvTLMYNf6RveX9XCTTVh2Msg9/CGk5lQxO4Y7Fp5i1et+tVeAQe4DSaj0
LBLUEQ01CXqcldhfmhy8bg2WFGfER1Vqlb0OmAfJMcxZGRlvBeV5oDTV0RG1lFlFOXEbiPLCemnp
2pirZqT+2LE0jiinzgn85IKZme854KC+YccrfAq38NF62iTFgLEdhdbY2b2N2A9LVzlY223kWE3y
j7+D5NrqMu8yLWXcZ7VazE5cAOLbCoOoWXXJ9Gsfoi1MxYHUVl0CLgfAPcB/oUD3a4H0WubbR91d
ateTIh/ibA7Vc4XrJ07KwNSFz4GuFNA5PANBK5NSWJSYyP9cYL1uL1GmIgWRjPKPZubhtukZ3yTz
JQmVPITKcPUiZy2B5FiChN45GLUmIUOKCBv1WbfoMdILRZbiuQrfQXprlt3IeQLVJS3vJivWNdbJ
zehF3EJbQVvD/PneSZVpmdxaIDmisQ9HgbCvRoqLsiY2JlgA6cZQZoezQZL8hUIn5GBkxj/bY2Oj
9j4ofj9d0tcHu98Xc3/RfdXeuNyyM6v2vpPiqCrWpKsgOxvxu4onTJGRKs0aOoVMo83MeqI/8rok
JFn2d2pT4j7Et+scRD2WtfK5y6o7JhvvC5j3bqS7OxxlK/hi0doZEbzEsaTq/hkz0j1xPWEyyglN
gaacqcYUMHfEwYmWoU8ZqOjim32NOK4iekRBv5Ub6pZHdB6b/LCwP9hRjqms63u1SmmFks7km0jj
S/WjFCuaru2CDZlVmTdOiATIeb2HPAft+rJ3sak/wPpm4pRxDbUWgkEbYuV8AeJxoluzatUc/pLv
JmRptQi8fzBoq2FD/5wUPRJC9AAQujYNQraGLU1zdJWAMD6zQtli08UYYnrZJJY78+TdFWCVwDkf
xR9HL3ITMw4Q6dPktSOmX90Np0BiBQi0qCkXFie7SKOitkdreGXE780mBy8Kh87YJYVeWMDd8TxC
sJEBQFxkyNZAR7i2O84oj5nksnDxTdrz6ILvzZTKej37VIclbkhnR4XFdfsFSeT3x8kstRhEEuZ6
l5PuNOAcZfVcWuMIDGQ0ytSLvJcnwvkJIG8du2xv/NMRT/bXAZmspRHhjLqJFqW3fNWp2kw9RBsQ
RH83QWhuWiDxHYPCaKNfCb4DJoCDIzx3bqA6CH4vUKUQGU5vgKI/UQ8ga/qHdSAUiUbBxP+FZYvB
NMwlRD25/hLA9ZixM617l1MJBeQo/WYvoyGuqYQTo+KU25+x/9bJxRC9tTJMevSfon/ce8nlMpcI
qVm2JkEfEzwcek3tx5YB9NIuJkGTYihNyAvEnMgtz7j4s3P4jtpEqwrsdenKLeDlJf07NLMnaxqM
48lHcnNcDJjrDdkvYzlGOEkxY6xhgOB48UxB4m8WK/2DcR3fjzNV4wE6DfBqVPhuMg1IQGwE1TeP
3oD4p3mVe/10q4PQS9X+qaUtJYFTM7x/s6nL8oOPmFX7CQnfKZaUbzk4USMH4qCbggKh2UpxF+m7
a3pgjHEccE86+3IjDDbmW4azQaVtwPxzmYauBH3SA+60/36ukBCuDcNJgOGuY6c0cnwsel2Bek+y
mEwFNzVzSTeaEmsB4MBkSp9qHTpOV/9XROptN89ed11FsGqA9GM7bmxnkOPP0XXl/35jYyvKeQda
7BzyBEukCrh2GV+i0bb3xR0MWBGXtW6nzUz7L1PzT3ChH3K0nkx9qM2wzdsVN0zHhZAtGJTUNb38
YgQ8JzwY4mf/T2sBGeHUSMyO/xyikTvj/atek493E+uxVn+O8TwIIyObsR0x6FzPUd2XHg34M2Ds
4Y2YQjVv2tn9RB2Ruh+oYCxqJhrS/Cick4geyF8MyxOtKA7w1USCGykluWeVuZV0RfdJt/2xb9zu
v1zb+EPR7QcC8gw1DUxLeecL95FrfRSb3GGMASZEgyxYWuhgsaZoINIUHtl4oizHdtM+X08i3FwU
cwTbY1xhulDCpOtdjlFawm8+2OKYGpeddfeGS7j85MJtniMNkk2GZXh3F14srkG41KOnb3jV5TnT
6UxcRTkVWjRcsYkwHmq6P2lj9u9AyXOkUUlmkPi+gj7nrcKbwvPOxBkF/qBcLMMQ6itEn4Ti4p7X
T5O4gGEIt05wLVvuPoSPKFtcff4TFCyCsJ+iavJ+lyvF/MQg0eeimZvxfKmL+HPLT4ozytploYKs
1hATFz25tXnYKtw9+RzFuKynMdRxFmgIv4aMPsovdvjHXVoUuXnKOPfQHnzIRwxpzjApmFnyLRPO
la+pQFaYueEE912vxCvVLk4Buoka6ynTHOoofajNt/bamgHKpd4fG2NxIiA1k9JE+g4fgZRFv72T
ueMS+sSoYWs9XvGimXCx6hqofIzN+pRO2zDv6AUy/+MI7kl6NO7ie3+aVlTas+BWby/C5+X0l8Bb
15itMb70PPm8o/IN4IbdI7tNAkEG/kFmdmvWQT4Dwn5ZWkipiwGdqugRyvI+AopRFMh+LxnbT9h1
wrkQVOdRlQdzL1wU3rK5+t/p6r7slAB9Gb0scfXdAzIC5U3Tim1+NxC58D+DJOYVKE59jnnBTWhF
mDDTA6bCUODq+rAnjBEGX5P/eQxDzmTsIKv6wxv4Wql3j4f8ejliN0iJ1OBXz60pMTP5/+Zer8gg
UUutfwtTABekKi1hLHyGxdzqRJx2S76TwsqvGXZG2fytAS1/1WXDug+KrX20Yly8ldxKW4BeN7b3
Ofkx/ItUrh+/8/lyai61SwfZm8hAZQU67jCgFroL2mtBR2eHRgOU342nPKIuVbnor98zTtDVFyqc
oDqAMUVnHAceJviiXgHFjh7SR4RhAk9AItztAtStBYmwl1TtQ/4zY/iDXE7J46LWV6YzixpvPOB8
f1H3/8fNxNEhHbSlqPTnxT1e1YvFb76j7fx+M5aG6JClNIC6RWgp/kS0cN1MDnnudG/Mq3aRRi8T
N6QeNDmL2t26Muk7PxolU9SbtroFQj07anoR1Kb122dBwow6iOgMDZNegL4LrAJBznuW73NGCQ1M
B8SqPWp4ce6lg5s0Z82x1mRa9w0CJx75tv4Hqb0Gx2SfEDY/vrowyA3buEOl2hiAL5EKHvPzHy6C
MQzmHU8v1Fu2DT6tARISnMgWDZG02JDvsBjQqbxlQq0OjQ9ZmpEG21KCdxxdY8/ZuvTLgYhBVcny
hdKhiKMK3E/JtIr1L2qpJaLqVQmvhyYSwFtd9qSTWT9g79wr4lnc6LB2W+blSzWlducGr8zGCGCN
g3xaZTQl1HYYhCkWwAkWAPh9OM6jb/yahfiPvmlHzHA+RKVRuCIG/dLa7juRhLQNkeMuk7q3MSkK
7DxUyeZ2A4IJJTVl3S4xZTiLV8Pa2kCrYFT226BNW+ppF2eUGQGOl24mwNAUMZkGAx/ARhav3h+x
V4b0bY+cmHmRxsBpTfDYBl6ZN0s+NiqVcJG9L4oQHodh23gnHnyKNueHH1fTba5DwkZM+r6+gG8v
cazJf7cC2PNewE+TeeSm/xE6DfSNLgs4m4RbgsCmlwuN6u4YYTUgK1XQC03aaqfIYaLi7Y+IhU9D
PlKgfydFKFqtRi5iYZ8Hhttn3GBGbjoa2rgHsJuW5SCjDIV/jFNQKcRRhZhuyetLK6rsSdwlQ7N0
B4KzHie1FKhHXuEhWMKpWKJ5fHCDGUxIJjjKWixWiISMXEuctzkJM3jedyRayT9+DQZA2YKYye7L
AzWZjAZKFSajMNJTo3X9UPgy6tYCDD9IvbBlP6KMfw7Jv+RHqNVmFz4ZutXS52oKG93bUoYcdcb3
RlsLdnKGNHhRHdCZS3+M0yGqDJ168e90/vYJc2uVvSjpYrWYnvry0CR8PH0NiOSabMV97HKUFTJu
tC4scnhDMRLFD2WEJwa5SfEXocRe4vyaulDHs6MJHCS1L288MB5HswlPs2eOYa4oe9eC9XX5yEZG
74tmQym+SfRoXOMgZXNJQKHyhJ1xekYrWjee/VXOArk0fhyXjpLx5KLuDmOSF+RX1occt6D5LLVg
7iud5aemwQeCnbDE8x/k/Tp5mUJj+qK8vF3tsuoAKsrdrqfmsgmjlCcuSzrKnrcu0tIQaR+dbCST
emiEGextG1LDHoExoC+jMuHrFDVwqSg96naJCOjtKvutz6OA2bg35UTAdHGNG/F83Qj4WzzWOA7u
INhSQ9Dj7xoRerw/PoAdTn6YfMln+DtIdugp62ow3aoa0TuULABJjBj7YoTQAnaviQqcVTeyOQGK
tw4sePTfy6tdGp657hMZEmEM3LgJ4UsFp3DH96HtLkhLmYJ3U9SEPdeAYHVXghAmlQ+4ufrno3XD
t/T32Tk6AZRmdGC8uxiNDPqd1oMQ3SQ+2OUxid1eacE8zsLITzn4lPJbQpETl7Y3nUelasWA5pYs
Hd0dLsNJ6SgXW8YsvOlyAAV/a+wueoiQhTkiZ13MtqiJJLnBJKOgJhovR9yRtp8uEgxbn+BgqIRd
3frSUxZyW6BbncRtGRLPC0gRgbvJnC2s4aszcaRQ4rIRYCyD/qUXGBMNlMH7+anRN8lfefFEONK5
jK25D65d4OpOLbvO2R1WWreo6F1Rq91llp8sCmvcZClfhfd4fO3gLCYmcE9aItC2p9hzWMekzzBQ
fioinBoJeZkJD6NImypXBfayM4QYZHerVNMc4kzcxqy2llDbR1J0hAz3rRFGoHakncLmvXiZ/dYS
5eRJqQ1dhDXUvUdaSDBx3RciVJ/gqb0jaxX19Ah+a5AB6R+1giSWuhKs4ygDFEu8sarNC9k7jNR+
uNcrzwxHbsfraikrX2lsTIXd/mX0xYxppFjA4+kWLvZD4vxIpxciD932bZYLMHfnRFBT+ZLOwmpp
GqJCdtURFVgrq1rUpmB/fNFdx//CS71W8ZXF4g8hUvKip/rwTgWMrdP2cIFkbheDFPI+YQus0rI0
D67NEdtvFDt3ZL33mh9LNQ9N2rhEwm+tbSTJZoVXChNjvNezyEGsxyIrhUMulahXllMcNKyLPLwo
U5vfio4l9SM73tRy52ExnkqsjJfb3iVZMwIbOSbsz37GnzrjlkJ9rJcPe2y84PHDdhE7MLip6TRE
ENGXq2C8Uhhw7BbwYccJzw+61bDDfRKlBFUwVv/gPHonfIShp3U7pXzJl45kOuPKUWlAVqIrrYva
21IgjxpidrjTrK4e4OnSOvx5tKzh4A2yG8tjHDzwBoShrRMNBYxNh3jPZS2bM7LtqY6CRs0BZVpR
UOnpHERslMp9iz+5C1yXIrICYQCMMQwOXEdDIO88QKPYShmbGOWRiQAzl5cYWDuEoRsgtlY89WiR
I/qJIsWofwOqlS0jVCgyduwgidfMYW6ALEZ6EPNgI6btI1aKEAR81CdfvNVB3Za17TZtY8lmIuxB
moNdkuC+bO5HI/VLKZerHz9KofN3/t5CsQd6f0W/tLfd+xHP84Wp6GHRa85JS9hHRn9L6EBOO/jf
TI+pHKEMT9dsfjezbYkh+ZII13nvoyYMbqBlAYSB/YVUp4muSKlP2fl0hiNdblyUZVxncb+KUK3a
Yv/ARd6vNwfeYBaz3cHkQ/hxQGW0UCF7ryaAVOg3TJW0HueIGJB6UiXrZdH2EbC6LUI7fIeK2tpq
fHspinehvzetvwbwM0wUuvAF7jFrk7SrsQn5z8fL0dR3Ro7iiPhJsq6QEIYVgl+Zedneype0qe0t
7pmOsFgOSSYZYnPrIYRbD1+LWnfcHOvds4mxdfBktXKRqX9yVuav+nrTf1KVRA+iNQ7C6q9krgH9
Ze7oIV9n7ZhUdVkMpc5TUDSPvA9GtaGHyWcldB7wI7D6ETADu96qL+Qg++D7Ek7KL7EBoBestAKp
xFGeLEO7HKhCgGvkcYDukYMHucEv3aqZSsH7utv+BfTJrrQ4yy3cY6ojqUcGKXb8snTidObb6RYv
RIfeNgqT5ZnFR/LGMOoWP5zIV/o0WpmC/qUKV7BpNfgHn/wGaXKAS7yU5br0eqb6VatVh8gS//hC
/u6p8AfJcFs4fLP/5yO+TGP2fUUz7fUb2WBcuv3ME7AnRvZZRjeY8TL9+KeWHYP5ZDEOOF+FkO3k
HohlRReVK/IwoQPvuiqf36Rz7d4FlXn1S+SPQl3UherBypwJTMFxMWRP75sao5PvGGsPs+IAUiJn
vT2wg3OcOKXf3PvzlA943QmREW2Ndcv7EnA5UcjlM2QVMlgoTP1sACjJpAfD+TpCGbvduz+qiUcs
rdkbzHOzSGFtmjUEsESiCOyniZsN7+H0r82lZKNxRRiv4ysPIhruUpVgLVL6zDw15N2slLENNv1M
cdLFIe3Ew+v5Tta8M1jWpRHpHop7B+g263b9w7oSKeK2+Mhn549uAjcpjzBqBRGQeXp7bYF84cPg
rKH7W7Q+vPWAmdicH5z5cO9ru6ak2/Gfpd9bZwSp3y3T5oHN2hL/CQAil9sgn010US5D9WeAASAI
iUsB9u8h+xXuo2FMGg7c8CXBl7y4FGwFXb4l6e3OKPu1DAcsWwXvkyUQqtpqkjW7AeM2UFV38v/K
gIfxxL8jcdin7BWpAb0Il5kKCnUbhygh+o+2ioUirRArkp7gK4HKTJRFrnCZA0QWAfr6PlA/8Zzi
a5j2cydSOhMR3mVl5zgDx64FKTvLRTakrCdGez3aTxXH9hIqWay0V1o26A8nUr+KLkqwUsTq2Bz4
9HNFLOdCPkJwGuztaafXUVyJT7qwxycWwJtFyiVDGY/1xmkvxwj+A5aAOsZCx9bV8TeTvPdWNZy7
YNeZt0lGY46AH55o2suFtKz9SLH6A+YD4DgMwSboeM+ZUYKBci7JEakuatplSd5KfB5l0528pYsx
hoNk0UkECsoT2b4SbuDdosmdE3jr9pkrnbwMCeidWYwP5fIkmSlE/CamqXs1ZP/SfH7IvW7H3gsg
EjucAtz7hjB+1A02h88RMYvLTU3u4pRlmE+z5KBgd3+zIXtIPJ5qBdKV2HS574N6Er5tSDTXgNgI
oZkNcJAaquqeMRa74ZyHfELdx8x4GmBJzyie6wTr0gKUxfuPaQVwKcqaf3yNif93pKNVJrD+274o
MfvfTtHc+zlBP564MPHsR7NMN0/F+EFD+I6g3IcDBIHbv7qWQOgjxr1afPS/bQ8C4spNhDDhgEpq
99wXL1F92JC3Rn/TsZRti2uhSWzqHdQAAPaDNTKEH1JglUw44M3aDoUYXQG5jhBpQAj63bdKW5WB
4UHYLKhXv+fNFBOZkp2OxJ1wymBPGeBjqV6MZSaNrNyUYkoRXHLVMUlxkHEN4gx8Um8KkFOroWLI
1JxLcRvP3AU+gqtotYcFnmJ03R3I3OTNfWbAHGBNc+KnQL+4PWAMQA4TUVRN9+vabgWBxGzyA6tc
3jCSE0hKx8LlykKemcQ6jI1SQjK+U3CYFAFwk97wefrNOsfQV7z9I0Kc87LqipfnsQMa+wTGaGqP
PQXy5URRkaDuq3u8PuymfkLbrsZw3UPFKWzWBahlXzXGqqsVwuMr78ToRs4WgF51whqgHe5bE5u9
9xVQCk4Yl2zX+JI8oW5ebvGp4za4YfmGi9vHRnMv6HDQIwbB5CMHqbEMDDIKop3zu2a+LwwgW68G
n0jRmqiH7P3v8CkUgUmBYFkdY1KT9oCH+IgKF1K0SYgWzj1LVbu1XK40u6FJd/aF/szuBB8Fb4sC
KC8U/2quYPl9rpS1mTK6anvANogc21Svqdd/BMvTQ2A0OuKhCU6mjXe8Aj+K3IO2JozoMhGQhxI/
5M5p3YWxkB5DSqGN963vJaSxd/nvCUVbE3VhtcmX5DRtCpplvWODdwVGCC1Vq5eamCxJE+r6HS8I
6FT03hAWaMKWkWHrhn8T2wkOTOrnjoSQ3wZTiz3OOKsIEYAOQq0U6b62o5+u0IhI5Q5R/CTP12yJ
VUCCKCjnGUImWAC8JICyzOJCYqmPI5cR75V/HdSWXF7fHYe6Sn1PcT1pWxiZv0e2tYuOc5VjEUdr
OXmPg/ODwBt+NROgaGjQVc2ZZLoT0//SRkJathhS7VUflyVzJ1zOwPKWF63B4Tk4Xe3MEXThxURV
uyfJdObJOXQfEFBBcFx2sQP/tLW/DVc5WOB4nSV5yKGSDNOHLwkBh95RntoOFvc2Nucbql3L1Lt5
LWpy1U4fTLHS+bYFpm+N/++8jrhON9mJMFm+vIrOZomFYrlOPJUOwGNpmMNeAC7bj6mK3wGwYdzj
3+nTvwjkSZBo1tl8D22v9ArunTHVCI6aj3uOV2NQCEupTvNPXfhTFmXsbiejXVy/6lC+hk1PUk7a
/xbsP/7sAVzb/hpUTBNm7tOEODY5oDiQ041mOipF3zZCwyUDGCehBiD1R7RbVm+Gshm2jqp4UGS4
0lqK8qF2KYdeumS7fjkMnn9VY34jrSvukxDN7Avn3uK6XgOS0hRoVAvG1LoUHDkT9WrvRnho5fxX
yuLchWiHbAbFdCYy9YaCCCtnTzwLuQUyBOwZ8uuI+jpOMfXVk63w/GB+aiJplPeeoGm3zGNhLx2f
p9LOLcYodocistCEnwsY+gOpus0Xq77X+I49kKAqFnOQrW6URS6Nz6NJb6y7X0lHqt5/+rCk3m4v
p94FYnxFgFsaWxpsZgUTXjW2Dt6FcorQDi9qTnXmpUaKxTuxuU9mWwXH0YQLWL3oX66vmSXiqhhO
pqOfAVXjyAg5ahWbgMSah2jtu0vsWJd50fVEed5/zuUunNl+OlmoUrBCPdeCUuFsCqwcKEZf5yK8
W2mMWYkCsA8DnJOnzhIFhm9TX+6uiH0/oW6VJ5YFT9LccMnYkVtdTljdw+R1p7+XUKYMzicP0VNG
xQgpGvKpN5x43lvkefysK5ug5ugxL1q5KjDDpJL2NXo+pLKjE+3FM8MEv+Tz3ySts/Q/uY/ktLNw
Qw1vHGXgmEq5yy8vG9tOUHtJHTGXCbjMeV8I3iHJe3VxajH6KfXTPKZxeQ3p4YMitAtMSQXBLIPG
8gIOMqWA3ik8vHpS5srGRbmHMbBiHUIAGyk8w08p5XcQqpjTodWkk9JT3r/FNU++SwaFCpT0FCjB
EVc6trAAmMjtFm4GiyahY7vTJGmRoiEpDVQRvmqGjRqFykPDbvayXwgzVh7wGXv0evVHxwyR2HcS
ytnz88Oz5YkoJFJMF/jdo58W70AHbh4fddYS/KAvGujx+f8/0k1cSr38YBgWK6LSV4OzEWB83q3s
4Ykv3lJzwoSHxuGSfE3FujNfScvav4jrnAPD+Ewg14XDC3Ca0a+cacV7fXSegCHqoVueJX+nbT+n
tejds0Z2L4cpWguuLYBIoJJYWtqWds29m287uor0K9RsazKeIDpLCSLrd4x15HwehBH5XH2hzLdU
WbHR2a8f9cmBSNZVZPI+dYCNvco/K1QbpLF5rcx3mbmu/6gY+yPy6+1HBttru78Y+JTRhOm+nn0N
C+pS/yTWLRLo/RILQzrAWqIVjJDmfBryr/0XXE/+tbqxSNG+sbl0FzW422+qH9OJCMEd8ArfOM82
eraEsOTzWhvKqTrS2SW1CFadcGzx/EsvCzh5OU6PwEMDznqYAF5irviUzwHLYAJdREwqJzTUnnmv
KoA+cyA8KgZrXH92kDa7hhATzdpFr4PCSAnb+sz+GK5uATiyPCIpXDU97XH6g29/A5EkqlpUdxjh
FVI5MaMJ+XdudLEGXnwwYXUqayYCilCe7MGG8XuwV+Vc/W2DElgBEFBhxln/ljLJTG4Y8qYrnj62
ele+/xmQiL0qp1a5P01fLy9CmE5D+dgsmPL7lFW2T8lRc8KX9lRokyPplTTV1SCcUl+pQWRE60NR
S4FaiPEmd+eQ5tgd1c5jedILtszxnD8aaJihRHUmXlvvFdLkp88DpW4xCo2DEcbEcUx42PwN29Jz
6MQZT8JoMtl7bG909vSoLPkq8/cFufSHYjvBQn2heCapMknbrt68+Gh5MwhTyJdK+dKXeIn3DrOL
lurGbdIsIsARIJJ4GERi8+szfbetIqzVdsCvgRDG3tmACIGAmxXrkXIJVtzECSZ5Wl1JuXrYjUYW
T0ouGP+f/MUBspHF/5DhAuNl7ix+O16Z+mXIYTSVxrPyTZimcZKBqakK3X+UkYMW+OtP1IejQs9w
MGy5tvXUSEaHu1Yhe9dwxqYVXtlH+IdSV7N/zMXRLvb4lNRuPXZe8CjxXzcfvY6ZvvABjxwisiJx
HuFdp4JIjZ+gVxJfYnxLdQ7A7e4mvwOMaXRR97iVe70mVNLzD7XlvKI8JiDKNavRRHOW/FFiUPsZ
SkOYA1JGE2OzkGNexjG7hGnkK4teyewTfkeUyjyESff/5UQ7wvCLttTM5Vf73DMyZPOGJS8jgXWg
TgWo3MOPbgHlTvbaj/HhOnIDhNwr9DhyLAzhcZ7nz9Vh7usCcNgpIAVHltPGcRpm32fxmepR6Bs7
AEHz8+EKvM+aZBp69XSP+BkPOVHfovZ+9Vj53e6gHa92goTU9hivLnnH9Z4S4eP9xl7WhwiJ58Cn
NUhCSj8heetOwS9CCGPx/dhjZLcM3oeAMOj93Tvf2oRcFhQBooS5IVi9yDCbR7wGkK6AgU9tJUic
4rE+OkyHmL3kHH8Z8/SUoltkcdrrBhJ/avxzUQjOzWzAwXIclnQ7eCnPK0+iAoQl1o2hTfLYreE1
6oenFw2LSauiqxzfKp+MOnyAjcRolsGw5zmM1MIf2EW2xEIFAawEg6T00MuVwG2DmJkW+ZkWOAiW
34A5rpdhGSJVZYSJJGvyEdps192n7ZDDaqE2i2hQNvVVKkLwjpoMBXP06R54GUDvum8t/U5xoY2I
lIXMgLnADkimNzA/KF3U5delhEKobDe/6OYVUdBKi4uegIZ7c/SrprfsRyhdCn6pTNAWsSFD6k9o
C6znpsHhuyJ3zeFxbFAI5wU3+Az5ppQW5zTIyAeSYENOdheMIbdcR6WdDVHK833vM8cTdxaxd9Sz
PCnY4GZMzHT2FNhWFUzJ8ZzfiD7JGfSeNGFBs7eMZ4ko2KPlvlMCjhAHPfi9ahm1xEvywD2nV/ks
CSnoucBgwteAkvBxTNAZ2q5pgKLK8ks/NgD73NlCb6zDWIofu905bxnYYKwTV6GfJLKY1+iZv3to
SpHs5ex06il6VuFJD3JBWALfEZDFDDqaQPus/NdWYEa5kal3FVRWY3ZGI1ICAM+/lCSGVTpX0Ma7
Litz8DCcoZmnzvNvHVxRpAJeab1QALyM39/dwvzVvrKpFQibyghe1XDSWJBZTnPxTLfg6b4haLRv
4pWAPP98OgLDVSYpabq+ikrgqzWkSwTz7c6DltxKibpo08I4VTbEy9SZEhnnhBx4qv9sOMp7TpKF
R1ikxGLLY0ahltXzaMEH+7rhfnpSnsT2DSnsNEF8JfaYtA7ME2gMZpcYOSo9x7hDb8DlJtIvWBNq
S9RoeZMCvm9ENOWAzjn+2XWSKJdgy7cVBCkW3txFZ3ZzhFL06dx1GN5sKYzHYLck1A+xEkiUSUe9
q00lfhZybr+TYBC7G9R2XToaq8jqAbq5hFZ8kSWyQMsSae7V0IAgLYUcYKhYKpDLjQLFcGDKYYuC
yl2J/2v5/ztYOiQ56Xsts8h9ykO5qCwLhjp/3rm636zgOfwZA0XLrWBhPTnn2Nho0a67dCiNIQoN
djN7XBdo6HV8n9WgxOdf6lvrr9yJs4CgAGmnrabsBnfDrXMWhjS3QT+o7faJ6BRZXFdmAkfzPTDv
aSSkcnwfeG9dKmIBnVUwgDm0LsafWag714HFtAn5ijVt8+PdeYa8NjyhFLff5vBr2IHLE+/xiQSN
daE7j/jtQuAayqK8i74V78rxQ7VOIhHE1Y9fgQIxg/vgeWNhvx0gXUGXSGl+9IAL8EDhRIXQ+msP
5XWlkwQCR3/OhXzOGTvYyOV59utepQ29NIIHmXyM5xCjuueaoQTHC8VRZrcFyrcNgac8cqdyIncn
VBoy9/U1RnpxdewJi1epTEMphUaAaCGi/NBLBHBOyO/v3+YjTgjjHDU1xzLidbrvciFv7jn2U4Dv
kXPkcTLRv3xLqQME5kC7FRwc/O0XvMcp05/8yRuMlRu9AHLKu9r0cPxfXvDkaXv/qkZCuoBDvCAY
o8eLSmOJan5JHpSYSP2/j8ABr/QcdoHspuzQlwuI4OaYxDlt4hVVDntT8hCCiZnJZjdSzGW4zeYs
WmK/xksaiarXvxqrL6WDmyxvX/GNWHnCB1XpkCHqgV6oRD7F6Ya+dV0t/W3ZQUdIQXLnuJrkEiPL
N/tHd3ZLFlSEG8hd/g50Uh1y9NaF73hAK0pVXzvY6TOPTAu7v/0WGBZ/9TcJvswowfUlGfIJsjYE
3kQK3XOmlNaPvJl8iIEtsfmsxe5WHm0e7zltw7CL1UOpQIZVHohdgMvHXYizf88TILQ6H/7NXbrj
YJynMoER5M4xxH7hur1C7sPPDpFy9Apmj+36/sV0iptkURAfalbssp/ZYdnc/I587chVfJXSWPpS
aYsG2rTzZw7ilnzojt/9vFgfiYzEY92UrgdKGn7jwpwUdI37+y/fZaNuHTziYcZKEg85/13ecS4u
3KbyVsOdPJTjsp1YxWjdVifetKXngdpS1b6awAbZyvG9V42Ix6cUjygLJmEA2F+mLvaR11zv5B3w
ORyqq9uvGad+Kk8ay9oUEWhBv9Pc2xeyghAjcPAX5tUQnpc3IYi65SY0q98HUsv1O01RQsPmKK0M
qTgRjO229Pyo/Coz30pADguAf85h6Ede8A+TJscsiI3ak//5x2EFiO2t+ADMZaTouVmW0NdymERc
fRemhWXvklqXp/r+M2iVwLgBnWCItlcmtXb/JzMZw5IdeB2n1g/L1ahnTrZB5u1PfKU374YkwwFf
WoXabeEboaAFQ+U+wPhAC2TDY3AlTgwjSwfcEs0OM4VoNzzuSWv25uHC/ehwDlECGdLvsfd66XU0
UAonQL6r2VNdbyLAUhaY5uUKOrzoM/KBJEKNp8WklCZ3QAggLX9O69kql0Ye4exzQjvqu7EowEZp
TIbaXC2/2QxLyID44p81gLsuKOloJfG5Q5nxwxWDWrrjgRkteNBnvWLNmundUJ+zNGK77+3HCFe9
vYspG81sk8Kt+IGaDvpQla6z02TpvhIOtgkK5xTYnqb66HcIm49dN8IO2t8RD9gv4S7naMGJgccP
9yDxaO99DzTP2pHnG81zqjKW87Z/EQE/F+P7t46+CMAMSf72D6Uex6egOWnGUnRlL+R9StMJ0Q4G
+ZKlUaRColkvOWEWaSbyZ68oWc1IcT/7BeTCGC/ia8DMg+J4WCs8Ackb1L2RX3fWXK2JEehWo315
/4Dwfsa71c+Tw0/leyhfVSWgpHKcAnNEbJrC998iTgDvPMCfLf/6OcfC5dTkShkuT0oDQvuaMxBU
nYzx3xmOl001tXMFrm3jUT45gg9PFnJGJPxZZQeLZjYs+wIIp5j6cWfO0zgGGy3hvM8aKUCAOWaW
I+mGRERmEKSF0TtokwywwmWVm0W9HysKm+BAb4lqy09zvEcbAS8MZpn7J2Z5XP0saIsJm5Xfdcqz
gZiAKcXTJ14evK+D/2QrkiG1C1p4B++6de93ApLclh8q4KiCHD+HQW7oLggNFOv5jMbGMrgw8K53
N8TxSJo4RN64Oda1wm9TigRxLo65iZkPMFsV6esLV/xoIbdt3WMDmwIyBO6mAUZPKUGnIijdDipu
OBkUMjbCJtW7cz5yaTNEQWN5lE2YuBJFdUOKU39m1pK9FRuAvEmUCZkqqTmOJHLBek/kOm8L7yGr
+9GX1IVbi12CIQ1zQnDp21jtkgEQCf3r61NaX89W8AYjpu7uk+2jXBGyFVFuKHAweva/8/yW0hb9
MLG1InwWTFcoZAtH7jgnimrbnuorYkKH9w6fLFeLn0rAVRX1Xeb3/F++ATxROn8uYnkcHzydMV35
eeUatBF56KdfCgtVWV2Soh/8NErfYO4kCZxZermOPcF+/iwXmuF7tZDSHNXVQnfYSGiJmiWZhbxO
jjBgNJrjBa4azyp3k6WpzLqplP+hGrxLHEIcsZ/6hYiyTbolobG7H/tdAYEdOsEuUdD1YBj9R1N8
OJjh9P1xMwZD9Qkn10Sck6nrplwOdA6zJHoYB+CLqnZQ5UiMQarq1pljMMlsQuQTzImNOK/7N3CR
UgEzB6jrbqtL3B6EopC/UxA7uhjk12gVBR0V+6MX6RSpH+2chZVy5dCs1y5gIhckbqwWvLRoOBSB
ipXnDwn0rZVrhaZVO3/Y16R7ZaJxcnR2oulgKp9XtC/d5C7fbYYb8KzZiBEKG414van/A8nRbdi4
0npBymHdhrS1jxDbwEmgpMHN4sAU9r5KKS5W3AqeU8gcYNRuZ+rdgcnYy6H7bkfoFmvSPARC/nvt
+fnNA9CRLtG3sjTzCt0RroS0p8cknhjMZMCTKILiR8HZ6V/+4uBK+KtwGEvdYDeuyMWAjDb1wXCA
pDHl2awcY4dyKYBFeb+ccIcwPN4R/w3/RFxmseuhh0f1q8MaWsraE4m3gHCdUr+CBLUc/NPKav/W
gK+nIJ7IGhkocvMOXN20G6kX95qxnCsvQFNHIrGc8tlUL2tA7FhzeYN3hXSKtbtkjyTVS4rtkC33
QSluFvhbMs31OXcv3PDGe5cRGe9h1s+NmjV5qXMv3fKC+qXlvlF5z/XHUq6eUZdAY9dH/tXrybnC
MsLLazCLC+I7MloZp6tRmLZiFygN7TglVy8rEl7513h1lwhhCOJLMXrdUKbJApoChEbozqlNl8du
Xqe3ARAk7MHuTC90to8f6/7d1hZTDU4EYmymOyD4tnrHseAo2tuvAz7TBxjy5uDAxQnHSonnTDba
YoNWhjLdf1H2mOiP2aGxRWmXFLsnVWNHRnwmpvhzQQOiD8aF3rHffNCPaDXpX8ct7jgu6QSPKfGa
cjLBKNqbxQT3vnq5qS6xE3AUAA1vgLgB1cOLEpi9c7fBzIxy+juUCxtMnaYZBJje4c7EV66CMoNB
jut3P07pGxIb1DmGirK4AoGutvuWXcTcv0MhDuBnBApGszZMd/joM6m2SnBlOsZghbZscTG0sIRT
bj9sLf+UJd9dbb7X8rqBqTN1Bw4+mjNbO6vl/20yRfD1QWz/4uUlV45GA3ZYFpMOQ/7WZ8OnC8Sr
j8Bao3RUWALVAuzyVCa7kVDw/T/+uBMFt1tq72z3bAW6AJMEdu0PebNInpVrpXDP0mkIY8xIFdH7
mvsb8sCsT7P+i181NEx7c/AS75G3J2HiN6zxY73LXtscqbTcyG9I4tP0y4YiWPa0nM2rXb4LbDji
c15Kbq6J7D73jbtra43RKgGCd5fVXf9HF4ca0lhKRb4Jed+6CVhkqHqcd2y4Cm7GiejoiVFlcnnP
TVdAoCqiDZaJP3/jP+xGGG2QhZWTDPJpas/VBXCnMp/8SSD+o9gtxXziy5P2lp36Yq2xszdzAJpB
VERs3bIJpwzPC3ZBuYcNbwWPv9yveg+frhnlSu98LU9pmAc4/sHgwKLRjq+fqUUGhRjWWT0cUOPx
2FiYNi/GHdEngev4S7MZN2QjrPjCs0nrzjxZ7REvCiAbuySYePD5JEiKCBRoHcllwVQ/9j+cs30/
QwOHD+Z0XzxcACYU9bRV4HMEfdYE4q2yOqNz+6PUut5x7hgmRzcvEq7E3yfo94/nqB/FSrax1JkW
8S4BqwXuheMX7xSdwk3XJIUTpo15KgE81r8aOuTf0CVfvoQMzhq3qV++rCWP+ZczFx9f7xP7z9uw
7WVBLq7Fu7ZPhZwKx+zEFf/NxEJbIZzjZLXuKB6spyhw70I44b7a+FHgtqEfX45DL/pI6t9kH+uU
NEdUG5Sv0yltM89QZ2lXOm5JDrJOEptfn81ep3+60eSRFu2enGRX20j74fxdLJ7VRsbU3wswagK3
Pdna1/TM4mUm2JprBc5yHTVHLdfKjmXPVOxRwpvZcuzkZYGUYH/6lXb3DOS2YlHGdx38f4OKO8As
T71xcloqVxA3GuNID3kfyfqBAnqtQLz5FBIleTp0s9xQQgP76bP6ujmA9z/tCME2jnOes5tol4xr
LuIOmagCdo2yDlxpaGkum+7Z+GIBVZ8MrQ5S8UF5WUaVNgX7cTKQy/StUxaW6AjCIswfJGHDNHGR
8kW8pUT9lCNSgOjmBPApHLuKvTsx6foX32uwmW/P9Qscaf6ZaVTPLFQU2GG1SepPB3dcyG83j6jO
mJFNJAikGdNp7HDey3wFxT4IDbg4WMhy4jhYj9dlt2SwMqhcOGL1J6r/PyG0P5xPKYMz+xq5e/hu
V0OHApPpxXv1PDT0ylezdQjsyKEn4vEQ57MLl+cHCKtnnFjaGypjooNQ024ps3rx4Aq2mOrl0D+g
FyMKpJ20mwg0hQD9Rd1+BGs+DtHia48vX44ddsNxOFSN5409XQz8vcPvUhAmGvVUBESDt64TQTJC
SZHsQEhOA4Js6GXkY36beD4DwRIBwVLV2z0xEubzcO+iJg9Iq+BeUuizB85/qcx2PSSa73XRJIzK
fc+fSdL4n7co0R1Aln9oIOoGfk8TWQrw8AWYJ1QFJAM7/U3eGXje6ojpE8UcUV6t3gJNlvN1MIMi
AFs5KaoExn/do6ijWn85vlarsZPiwWvOgTf/GMuaatC9mJcYPdaUl4lVVAFpTIjOgPN1Ul9wFdic
gPnojGg/qWDCHD61yY283jZnY/JXTwuBSiaz7o5BghekWhJ+LWloQMB7aDlcKC7RPP3UGSpvm5iY
ne9X6o0Ft3K+D4DjOJxhLaLbrUFpWVJUPpBucLbvSjupOPrJYqLylVMweyIOJ3T5qTnWCEcuutV8
s288LXKDc43UWfmh430MRNDHBep4F/LdUFTWRL1HX9XeTHgTRr5ThGoxtEBINwbHmSth/i6QW4xD
763j23g5QyA441MS1J85NpNLYYsBiTMm/YeWyS7kpK/QyQxnYsn6EW58ryVghwOuvy1vhSBeM29N
+7lPBh+OB513LWpf+MKGoc74glq1clEqOedOZK++6SaT0rK4lb7wStbSyEboSudpwUGNSXyiB1j+
3oX4yhLqWy2s22aUos9xHfLyTesOxIid5DTSpDrwxy7fqiJeHqCX/rch1HQFFPxrVMiKcrd/NYGE
drqzzB8okekRsNWNunRxM/6GObeqLyJTKYMCEjtJ0iQn+Acu+xsFC2fS6kJI09aMQDFcExNrW+yI
QowVzvfluJTNtAxHQWJxz8Z+xtBkPxg2Qcdt1BvbX7DLt9mzaMuWoLR50H+dTmeJGXngz4y7iJ2D
ngNBMpimRMZAk59+jqbHvlcfnGSaOjnQNOnC/UUUD9f4n4DQvJfNYvb3QNMsS2tMcJwSb2yKmN1t
4BwD3fJIZqvyZ/SUSl/kfaDX4YM7DyGX20DZX+swOTKwgaKJdBgEUVcOJreloCw/eW9VZs/VClRE
c1peGI9QLj7bpIFF9eZzED01nlQASnS/E/9nlAj/4AxHmdVCSJ8SotQ6sbeOyJBqt0QZEHtkT2v6
06vpao9ijsQLeCqvfvke/ORFiZ91AJJUfBZHkbDeKg0WvAodZDBRebx/rw8EYHa22rCa1Aqu5CHP
XMY/zB42HEunGnQ1SW94I0TO3tKNvD/xVeLub1e6IsMe2/n0ZFKH2w2ymaxHNDvinVVwlVeHU82H
pFxuZzB74Mx4xD/aknayBjh2jqv7Rh2f/XEU0AciBCtYxAXCgKvfUVFo0zCvWmwm9LY6mka1h7O9
MnHypQONYXjVCcNFa5YZZAu2nl9hnLNukakdq4cfUrz4I9ZT2wTSv2yoRpgMXbCKBmUt7ilhXuLT
k231FlQIyHK2/oCR6sDgppENOmRlsujpcLiTt2IBDsDe3wa/hq0lChEaD08SoUZx0CIlsVWtIQCt
CWsJv/i729EMxojshXes4U9eJGjdgfREnBuF2/+IFdv2VntHgcAO93iTPnarsGoNh0hS8/euHf+j
Md4AcioQzDZqWHhyGklKT7CsVCjPnrKajEIv1vDq2ZTgRRnERCkB9f9EhR+Ih5A3uFSA7lP8WhHs
EftWAHsqHZHaD2k3BIZUluHvC+/LKQGyrUDRajFaNtpLhxCFtq1wzrLbGvzBOs+JRnA3BUv/a/LZ
OGwQ0/jk0sBK/dDieWZpF0kw0PCax+gnYMcXALjvzSDhtkYCqnGS2qmlSPUyikju/FxK1hraaCBY
QHRYm/+ZwOUiQRD8ZBazkFxqFxDIYDBgaU6f37Pozz35OPXhh+CLx6cn/CKBJEVgt2BSZug2ERFI
rrVZcWlCOMwONSMMJXCKhCJHcJ6Zm2ued7GMI0qIMxnE8sE3GBFUkM56Um2rnm/UN+Cct+w7Vwh2
k4s5YxaXyiw58a96NK8RUHhoPQVidQBEKXLHWP0u35YtxMEJvwErobuonxX0zLsxfXsY0q+C4RA6
AUsUTjDlAptqMR7AV4U6Kspv76CFyAIkXZaDaZmvrV3SwgUsujV/GzQfM5S37hjzYYDv5HSB6arh
tsc/Dl015z4lsSLrauoo6tZ6VlCOsti1H61D9qKEF6CuhsoiOCYMm7ZkHgiLLFbQb3oM/tOib6hg
tWhU6l/BMLMqkgdvyPnqHCtYtgq3VM/rcB7i1F+enhG4ovgDYQ7FiMDE3WYa//gJaxrKij2Cw6pv
dwklqKz5GoAhFROmZI5LCn88wgPMOP5ic14oQNe6AV+4AOE4u2MezsIXdqiRkq1U16VwZa39Yyhx
HHyLH5F/3T0X7VrNiHJ1BioIX0Wu2asS/ngN58EUQLameiWnaPjHl5USiK2e5w9MCuZYPkD/m9/I
Pb1Om3mD/Y3pzbfVG/BcV51xCVkzJxuYCN3KU2WDBTsidlJLtDToWKTdDiBt/lGZltsEqNSGBn5Y
3s3rKK+BqzGaaa5gkhd62FJ99x90HF4KDgiS50Jg5tHy5y5GlWzdJftRRma5RzX3ICHEg+lkFFVM
UhFT7GB4rZ3rHFNnRS1QZQHxrMFu4lWK5V0DaWZ0qNhmZ/1rXrdleG0QCNc6rdDe14VdQZmpqOHS
waYpiKlx2Rbsl6KAjYlMYbnFkEIUUUB6bHGpbG330AXTJklYIkJsrjpfYv+dKIOMiPqekYiNtarB
gOO3UAaRnynjBJ/+Qo64kUP9GM8MR4jch5ZR/deFsv3XiPdROzXvbWDXJkyMaq3sH7eUCR+xyrAH
UcOvNWZKaixDvWcSsyya2Y4OaHV4mpZoJssugCi2iJ9gcJm4GZdN6CFqkRrLJAndIMrPgnn+/bQN
wj33Dwh8/t6s/hwVI9kPgbYoQC5s3Hya4CDBmHRq+fR2GL5RrG4P5cues5BOCNiLNdoaAImygT4X
lo5b9bN5CWpLjvPwSwSfJ/FE/lbzQIBkUg2WtcjTnoZtGb/FKySAk5ZGubmoHxiAuPl+ZeCboOgy
0HhpquM/v4xiRm63mw+THSQfEgEybMTWr2pcly6tVa3pcLFPVpNW6AnwptPqQ1AKQg6QAPpBJBKU
KE+oEaVG53JWaOgplRgNmtjrbYs4dAym2VtGrSCMzfmJB9E8sEJICNlF9Vu4spnN/UK0aL3yrTRH
T1FoVKcj2Wnom3qZsvpLzUHb6T6pyF7zZ2Is1psHhay0acKsVgS9V4T09mABdPrLrPjroQlDhp5Z
Htdgygbpt35nl1oEMKcOQlBqNjzxe+ul8rMqXORoHYX15SDI/1guDtIMcKILEOuAVeul98H77D3C
u9ukw5slgdAbukaC7aF4DuzEO3noALQ7AeTeG0gCHK9XojuegylFHJFO51u9JJFIAtuSUUNbQy9D
OLFa1fKpqv66Sk5ZPrOOlRcWOMys0iridMrkBjiIOKOrciX1kAkdwzeksK7S4oZ/PeG8ay548twD
p7Y0cUGvOwp6Dc/MzPwUWLHaSHCT2b7ycrrXAx47zooVDaQnm4JpsbN/9789EwGaMJBX7SDleMFh
GLD7nJ+D+dv2bYkT6LrleTyUsrlzME+eWhvf/swQeoMjNra1WLWLi9vj8pDo812NY3Dkc7rb8Yvv
Bs7LDnxHVnXE5wr93qBl6D8QlTunRNk5msKwGzH7cg4Q++slCqqsEGoZ381p1z21GmaHft8i/jdg
z5jP10wgNE3Lf7BARwiwqQLwdyfFQwlvwW+FLZ8Sphr1dS2HAWba/AZ3DxD6zQMJwNmYkqNGB/3x
QaG7nOxaEJR1L9v5l6AE/2rZGlTTolsVmoRXfeF5tb7d8JZC611oo5n2PbaPdyz6h1G8+uVCg1dP
e7/2alhBA3obTeUkoNJyAh2xoMcxWHy5vlKTtSRfuCb8o5S7bBti3q3JWTc5+3t2a+J5O/vfYqWT
TKfxmUzk8OCuZxd82yWmRUgkX9KIyHBZzCP2mjmrZ11+aUXGAl6yijqukWku/lcN/SqaSeqc2iuQ
ES0vIb6P68HrLOPIQEeataI7aPtFLTqp4mTj+YR1WtcXCeTCjL6lkj02tMrca8VwhCCffNCQi36h
zgKXJBlP7mBbiqJGJMY8nbOagGqv3Brgj30xvCBXN+hzIlpXNroB506G9dTj5MYkuCB6ekXCjUlB
wwwFwwh4asFTMmVNlqGR43nJg1DqOkITxYiaJb5lwOS7XvsfVFAk8SQSxc2ZaW66o8JxNnrwGOUt
s6ZIWf48OkSxZHPjePUser8Vx5blKWnYNpKy+XH2Qt0b0TVUaGXfYFED3+ad4PuAadzs7sBjq4JY
TOTiZq2b/9yjWI6y6A18hP7off35qg4q6XcGP2z7HKuY1ENBFaJtIr3FWoga1aYi1vFGAqnIu7Hh
YR+XG/UlIJ/rUG6cD5R5/iLzpg9dreaVmYHiQGpokBHG1v+yKx7kZpxorppjqcOrvqHGlU5RTIlK
5h1Ox9IqVH+NSuDURm5+KkYh6Xrg7APemhQjCJb5lSM5BRLBkU1QWMegt0WZRg6EzxzF1EkScu5A
Wvdhz4fW5ECY/18yvYjCW+HuXC4nTEeZACR3LGX8e3CcNRghQ11cesmmbNslDX9J+RYJO/rCjh6h
q6vwJ6yfLlLNX5MYty8m/VfcQFQR8WvZFi9SLp0y0UYFg0+/wk+uxyAlqZi9ssQd1jiYdCCIyxkY
6KlOZBMDqo2fU2gBUNrmu1YRmVAetAPAi9G7jOGGIIwdgjRFuJhebsBJwFVsdZ1VX7gfeR4Fg86O
mTUQB9wi1sYh2D1X+n+pVQWWb15ocOaHo/4V+bVG6MeTWNtgKK+/nlsAFkKzpkgxevh0HcMQNv2W
3GR+ySdvV4MEAdCMhRVou53ApWwv2GDYHUHh7X9If9HogcecsHwfxHY5nvtGRFJNhIMuDvSnKOiK
l+YXA9hTavOsNMeHmvcuQ4tThv0oRb/CNSaNd2im1/mnTNjiztac3UxFGjeQkA/j6a1iXAUPNaOu
w16U4YaHnZ73jtWMpilk35JsWxchQm6JlzEZbje9WPiitg8lrslVmrPMYJ51jFjSP4/pqvTwQBtp
mJVHtBWweTVyDHK48dd4E8SuEDMUqtMv5sGfStG2JH59jMLHYXt4evXMzd5IAqswkyMA9X7PP77q
BXcqcZui6Nn1Ns3U7jXkV8W8HLgOWaVnIX/0E3SV+NJViXuNhiv7A3zbk4sQFXK2Iole7TjMSe13
YV9XjuvgdyYypXNaxE2fM2Ksw7ULkcRzcSwtN5JHcu/S7sGWiHM6CP7rObxln1KmzKM9Es4RrcNE
ja32p6KCPl0j3cvyhEjenxk8U/60ifi95k+nwbvsYODSFDETy47yNTJCYKxvHfaB5lFE54SdRfL6
mn1hEE6AG15XhZk0GOTGN5e1tgquIITay1ZCDIj4XamvwbQvbO3vyJygzczlL11JbfHFBYuo94/d
ra19Tq6+8CONTu2m7eFS765oqfBbW8DxBF8q19lkMmDByWZCtZvldB1rQ8TksXyKbsgcJ0G/sIcH
21bgixNUnhBePuaBDbYWU8umDVrky7MIm+krCd101XQyXLmLeH/k+hMZsqY4MFXjsMUE2oxBFUac
Z2DnHdCa3I9NR4gbOC2dBjCkN9jzKJDxVSsxjf7mbwDwnvSeTeAPUuWBj7Onc28+VlPSYYcfa7ef
xxjD6D4yd0mjah8zKQXmBpfF2seDbjsdEFnfV0u1NbI+bd3i+VeVC4v1bkW30WHnJuHHj7v3UmxP
Ptbng3VS727M4M/gA6bIPt+3oLVs3rpgAxd5MjqRRyx7OaunauI5wJQfREs2EOAHMW6Rp1s7uxtb
B0U1IVtCpQTCH5gD0Rx0NabJgGr0K9BY+SV8f0yhb6YNkeBgA3ymAH6//Cd5yymIyG7o16njAhC3
wnnH10XVyKzs52GuG3CEylsvyIkierfj327CnP/nctMbzKgFNxW+evkb/AbUaF8kTufDD8SEMJsD
kbnIRDdKZMWO67NejnwYcSyaa9dAtHUZljK1i0km5svyFQIWe0AX5J6u171dZeUiSisKShroyB7b
+4GC2KBrF7exwxn70e9UfnfYwvA8hBbn5V9K77UaovhdL/s5eeiipKXJ/ROocjfdSH9xhW652Y95
4DfSPZmQmZsl2Q61S+q0jA3mHEzBrJJY2NA3QHZd9t+QrpFQ0+EquD9J0dBqELdPM+uThXhTZwzO
G50/tLhbMlxkqqo5d4/AEiYbHkosyYMccukvm+EyuZoyR4f/94Ek6J9XdPP4+HIzF3IL8dMG214+
IOddDejFDBcH5okcBZoAt6rzFYmFNad7ZhPOHCAfO0Lq78F7gNrl5YJDtyN4U9biAQWGs/OtvcZ5
nk22VYEsWIg7ZDwfpqwzVBReX5Uy7zlRseWMHawuEzSeb52LlHpldwE7iUAhMxyYmL1Zh8N1eXyH
ipQ+PHAINKwktVDD3EDMqaz0AtRZS5FZHuIOcMHxDkHJsH9ZR6PyXhoVPcGkYs9MW4MbSqOWrrxm
VtOen2Miu07EUntY4IZZhSdW3BZXzE0qxavJ4CoaCMFC+UEaJCK/NrPOdt4bMFW09HsEeUdfk8Z8
xb3ftIsFAEmuVzZtxuBz/MPBpX6CvVYlIBoMPPdyyTFMctVjkqqbwqlrjDjYUP5s9aufGGTCxlsm
o41DTQoupZDGnKh06STlMoI+aejdZ5BaePJYexgiAtXfGiwmMxIrtv9gjlo0twswEkKIAsyHH79A
Kf4SJxmvMj1Zd59mPp/rsgeVX4xe5vbI13deRJjkKkWcS0VxD6uQI3GdDXc2lLM3jNL/lYc47Us8
iQnykcQH27rHv5SojhEUlb4Esb+78thTC4/4rrH3yxp+eE5HIZRAsMMsn0fG0kjhE+uRf2DLBkkX
c/G8ukZoSeBgLRptsMqIHr04hGPCLOTQCardVRb47IWPl1D6LOLA5fuad/7GQcpg213XmJzRcNMi
CZg+9t1a1I0l9H7XWxkP7SgybUpXsHfRUVH1jI2e0FSq4FI9Yi18jVFmwRseJaldnh7BxRxwO+h2
EvW1ACl5yblpVP2hXLZdRuv7lWNAQQviboF21Ov3tSVPgwsmWFsBjFksDPkOzpPcGGHMNAHkegf6
krBnFJkfRa16AZe8j5/sL3iKa54C5DPLB8yxUsHFIzdkuL/r1fQwOhOApxQF6Ww6jKfrPoj4c8ia
T25EHH1TXuKmVtXL+rmOEdLF9e6bjzgdJasc+zEeDS1ZavpbhdTz00CdSsmiH+QooIgg14Kg9j2F
ndH4bcKTL1lcrmnZjYh+ptob4MTNscZ3XWqDVnB/qgWlSlLa8iYn4gN42mJYj27ZC4ijEOY7epz/
GLLt+1gawPQUDCQhz9Z3/k2eoAlrkfVVn724cv+snrKoJ8RCMWnTB7csJaxlGFOcwlzbMyd9HgQJ
ez0ny3AogCahQsRjOINQc4Clt0ZE0eLtsmR2/dKlyVaAlKqSDfaoyPO2T3kEzYdrYoTndxyk96Pf
PVM+E6n/QouOleAZUaVpRZrbp0L39QCxi3B0Z73Dn9yB6wZwn25V42QtQJzlELEiwP6ZCU3xZnvE
d+/WKv8F+AI7lZ3YBBVHB8jMcC0UlM+fLom8vMZkUatIe1YXXtPabxtQ3jJRfTxt5Sik4Et4zGFb
IATTkaaA6tV+lVze9QRd6/5H9s8hfiM/JNmwMk7d8OKuAjnb0awIGLkQhgkDRepGcxVBuGvKBitp
vbJHvv3zoFPnOSJhQ96eOTGD8bnocjHT+c0yPMf63ugvTUJkWi/WW0zy4q5qrYrtTiEhhMvsgBd1
sTDx320ZueuPbo1yoevmLjFoi7Eg1iFIuvboK+Pkci1Lu9ThNOj4jWKLTeMXrPeZq2QtrO/5jh+g
AE1n0lxpK7nx6bQUCod2x3updnAXc1exRyCBlSI9nsBYVqzfsiBzFK4bRCdE8tnhHenhzlpWp6fV
cXBh//iJg2A2p146yZ+mSz5aYPS+w9zlV+NDrAveafc7HXgBDOfWohetINlghofAh7oBK5DbaCHa
3rePXpMmKjiuhAYRKL+0Qb6B0JZsb8J7RhLO0cHxBg/fyz1lUFwb6NvdlzMPviAmtvmZ+eAMECOD
PVkX4CkhLM+NnKRF7bbN/yZrU1ze6/bH8XRpXc+3IEqES6hMxv1TlAKtItj7mWEfeTAyb6HOW1Ia
lkJJ9bMh19BcekqlZXzLfWHbRCvxomNIHTYqU8iIQ6rxqjx48LZbbJMvM5QrNfvi4eEnbivjpA0P
fpLZNoIU7S4fNdCMOdJFBIhQuCMG3cq2W6rBoKrKaIAwupq677RnfZ+KC0lk8/CEr/LcHD46In4l
fw5a64izopq3bYWptSy+CxAzwOPxIjlw7fEjCe1ONwCNYXbRN1kmvZIn/zutopkDhBW/gLfnbGqe
m7I+633VyZ+INtyxl+nuZfwQnbSYXf00bdHmJw7azHKTuk6nOAhQTUW3KYZADrH2HmEbV+e38OsW
GupoXmgcBMi67760n1ZPOOrU2B6ZaPQZA9gEwOvB+BUG1OU+Fhwe3HFKhD/7BHtvD13df9ozazh7
922PK3eCmypZtv+EBwg0e6mUn5xJqchU0kL76HztzFiQ1ucbPPUwr5pDzpPE2N85mOJJRHij5XZZ
MwrBjnKhJ8/OOT8QemNE/pYIut6I1taH5TpS3/C1n9m/VcyYW+tNfkJZWHa5IST+9ZERm1+OoGhs
GeVHOwDWchcpuOAMlccw3U6XVagOp3wkb0raZmenZIpC17hNWrDg0wzL7q4h129Itq+YyZkbTLuN
J8NpIb+vA8tN9nk5MUud6DAY9VNpfayIYLfMcyLqzkOT95Wg+soNQWmZZlA24FlxiLfXHUAN9BkU
3zbGsekyqxhZyufNfoLndNU7SM/P8/iAFoAfTsvXIHf+DuZiYqv2SyOOi7Y7XKCqUv1LrQaNKw6o
H34HBcllgnWKsy+wKnt+ItIOosB/etD6ZVAw4rhNXZsP8aCOCcGCasLTwTcFm2jXcY0QptmKyKcA
XX43ZehTlWDGCR0Q7QNVpaZfJg/EBTliCxG/2hPMXWjO9SIC4LAyaBGAzOqiNRCo6TyIziYSRbNA
WjPf4xg81UmUWz4PwjKCw65TAq234NFNjehnDCBHn7i5JGP+brkDn1M0ZpauSVwbzEy1jOOu0GRt
7M9T6F7vtGVSJ9PH1AOmzJXJ5chJs+v3sN/TAwadMGiNL2hjlPLF5//QYKOhrmPm00oLrgeuIYJ/
bJroqDi39LF0Gqiqhtn3g0iNQi9IkT2eNTSvxDniJPXvvQB7Ecw3Fmu5V+Gw0d2g/XTAaAbaS53P
kvM/lzAb2qS47N9SZ5FXNSgxwDTV1Sd0hwvTov2cwglAcs5j7Rpcoe5b+wxz1lQgtIr/z8OV1RT6
Yz6crS/gn79PnmxPrGOlkR3K20AngZiVxqWflhgsObMpX35B4Wsl7mE4tJ/uiDOG2/PYxAji/DSb
hHyG5piiv+bEw3JcWlM1K9+ftrmEFNE0kCUBqAmtQUNcsUxvlzjUfvNL4NsBEqmt8m56ZpSx+U4y
//DIY4lEtUAxu1OqN7UnElx7wqqqWWfYDjKGgTIdyElUZjU0sOSH9mmZdmAfrmAkWi3LsOS32Hec
qhk8Pn/iusWOqv4AkYnrkxPY4sUx76N7p8itIv+Kzuwc7mfZRkIBWvMeNmUktm6jam4log/pDbAV
pXBEkFvlXmmUwFHcM97VmRRx05wV9p5KG1IjZC1zt6m7V5rmkUpPHqFl8BocbSo2ZF6GaKm9wvPf
uaZpB+djp7+buUBuJ8vjVCMMM8xHT1NUcdOkwObs3c+yuWofFTfN9wj2lNpfd5BkkT8Xg0abFt75
ix/OVUiZXw3vGD7Fs5jelCmqT+vGk+mThvhwM3VW12fhRCUc03nfi7vz0ocb8pZhzgBt/f+dhGIk
t92WMXc7vRnCpfAH0iDbicHr7DcJUQ/BPnvhOFk70I/MTVtISevq5qIharL33/1mPvzVgGqpvSQb
G6UPX+zc0uZtHC6HGELskqVIuEf5fU1517wcnz1kdHXyWRNk6v1ecE7HH4diaPg9nBd8npVzPvFb
vo+c+M58CPbL0HK/+okBPA96o2EfhXE0wMyVULuqLdKegkOsk02EjaBqkGQcSOR3CYgBMzarJ9oK
1Kzd2h+Q6aqoK4oyp7yReaYMGkv3E+EVMBYu5jQ2WSu6wnIM9j42e88SJ1F3hj9ke6dxJFdR1qss
qbFb3GkicHxw9cdlQH9KTyvxIGMIH/Jfzc1C9mgWQnQew5QDcQ3m7htekBV1dN9CRtiMjTUxfEgE
FbQmcDAeVno84y5Opj+udhDpaQK5J0gVoT7xeV7O+DLxEhqkIWE1a/DS8Gga73gPxWz2oWAeVlW4
yfwuujP7aA5ry56zvNfBiLx6/7/NzO1nlsR2xDBobKWHtpYj59hp27HXCn8hwrc9G7rBlP/R8rjo
lFlUqO6v1uF2kd5xjSK05c4DdDeZk3iWbqgjNEd+9tLnzwlqtpIVl92yzk/GVl9D32GJq4kyOyBb
9Pk/yAfQsmoDqUvDGs28MmV9RDayLdjFBnfqq82XIWNDydDh0vTGBrzbrbIYLZGSJkQ473an0cnB
Ykb1D5xCDCzIheNJ2CkswRf/UTF4puIPklH4vgh0ZQ0ybahfv2Df0KmqI4HaXwJBTC2sE1nICydj
agVec0pZv42uK2ax92uqpqWBfDmPjXj7jR6DSEWY806HmoEl4eXyGtlSvSM8ObfnDCGYgy+ABbod
WYnDAdCBxzo9TWgLpLVqA7YgKZ2YmdkIMi4hP5zdqPYThCNUIHahXDhqED7b18f64yIfaDFEAlQw
eh98GHj71ClC/mIPeNvSBYKJRPlikbWaXVU4uDtptJ3gKZ1nOVdQV+qzk1QFKwXDkhMQ1N6eCQDd
YS9FQrEzmp9pfWhG9KV+FLd/c9Hv8isSPgeezhR+JSLWn+Op4mulWfBvqAwZx7jGEGQpZykc+5Cy
zZ2YmlcnK1Jvvixx21MKHj/exClhFHH3KvYKWD7mt7XZeD4veH/w/LxW7AvZpKJ130xMXnj4ETLC
231RC8YvtXaRRXG+vGRrMPrcaTxf+KYpgf4K43luBWlLNCFBvTQSLXG7fCa37LKklmuy4XXSdzpD
ZR94uAJyRPFGAKAGNGlNX6A0559DS1vc/gOLB2hh55CxoIFl7zfKc0O59ksC9OJVDkAeDIKmDboF
nC7rA0DYlYKCqkJHzTbkMorKUv2v3uPSFdbnlZSVJ+ZjUcvEcQTg6sIrSJH9xRCfMyo6tjB+LBs/
o8ie22TZg7s8I3tfZIUYLdHQLL170+/0a0jFTM+s+OY4wL3A4jNF4D7B2dmuuCBbOlWmZFPt+ggT
M9BQmNzZfd9PmzVaGxu25yrDuA8RfXtW6wy2AEzWZ3ZBkB2HjnTH1KCWAu8wCfj/x1UN4aWcwZe/
jkOJbWzt9jclN8mbD6JednTHllOfjiVNH6ippnW7p17ZgNmx8WDvs0vfuQ2Hn1b6LJ/q+WkZeERn
BQW6mAVpcKj0cnwG/bFadkXAMbnBr8/HFNzol6hkVFTwhLBu+sqWPvaF8YSLB7rYxMuWJQadQOr0
2GCeWjXLcv9zFGfBDwWSGCy2KMcWA5o17gW2lOvbRRvd19V10JIa20bmys0mHQnhDQIANYCx4Zjj
ElGemzZccKl7bpfY1zXI1IPM8WIzBXxSl5O8XfWGcAnDEgN+HMkWEo6DUriwvhT7Qwt8DySdc4vP
OAzRpcQPoepacn6trP/Q7HPjUTDCiGfa0zcJDHgqmbJkSTtpBs15Zy1DhSg2IclCN5T1DQbXD8jx
L1v2u3BlnECrZTYdfUYXmUyLzsryFk/+Dh2fPPPyZxFEAV6Y3ca1BX5hYV8IJ0t3/DkDrOqvWPst
vhiAFjH8r06BUytXWSYdmWFC5gd8fZ9joyjq5222RLpkfHVznATwQ1XfhBnusSMIhwkgIsENNRlA
cPpsGCStSvSIamfPDpGmrVcQ0e6y4bawAEo6J04gu9iu7+IQ9DkoO6XHsVFZP44g+ttFSFDuBnm0
lxvmdOzAeoJWsl/3MUg6d8bkwfq6L9bVJxNKP/9YqAYK0LQsjO0xJCTqJX4dNYN55q4lxdSLhn/T
jtkjL84mzc9ve1TIf0x4rIiNypBVOJ1UuJ33loql649eueTYwekgFKEyQZdOjVxhnYKLGuiqM1x4
jPHjHmEHxm5qt/Rb1oNH16kZtPtXbNtqiRxN1cLSamM2LicKA1HrknttMOkUgKrbnrqW9YkZ+RW9
7K8aoxhY9B1vJ4l4vUEA/Rwj7kQ5Vug/22N94lmSMY0xqkeJs1JS38Ge//qDzX259xCmmGiF8arR
XRCuRHq9xKkTtENA0G1Md+EcMLJqMT3ajQd8/Lrg8P4urHtg5BTBK5IFaxulQhYD9vP01s6rD12d
/XqCndzmakvUPihUV5/jfoQNne755fjtvnVJr2ugLEwid2WeoWC1ymceuHwBnGd6U+Vr5rdpyoKz
e+gE52IKeYygImIMB9AddEas+PQY28cEiB7omwDZ9JrOlrqMrwPLmMVQevbelJTF5kQeKtexU1i/
8eTT2ViFyFNPHIcWmrQtANUM/2jgP5+2Qr3McEriuw527g7eVcrBlD/QyXFr/+GSP+o4m/7wXC5l
8a3NuOAgjre1fyE/IMJ/MaoTk1efLkV/DlmzGQzT2obddPv+ppDa5/FskygACCAAWUJac2b4Hf/e
UfLG/VN78iG7KRC+MMrcoUN+wFpPNY/8SrxGq1RbMaC23v0V5NkX9DAXfSouTYDlde8SB8ct29Zf
EVlHG23GZHH2EsZI4s1yNkTFAPujmaQFQUDg6gK3AS3t1Zp0mKUecLDJ22vie+tZIR4olkFI0Ytt
4VNYYzikaM2h5vbz145djlJMYrdVvmaEpY50t0KJySskeLULCdDBWHsu6Eb8fAqQyAjuyCZX+DjB
9uSD1aMuTST9Vxurj4TzckbNv4KbCPIZpY+UiKj4z1TZ4vMelTQR5cl9vKMMs2Z5wNtfdQC0/hcr
c5RO8O/JwHDJsJS1DIRBA5hiv3Ul27gotdYpJUIhV++oAFggkYCpQ4uYxSODFSkFZJ0YpDRMYMNf
NN2tpSmyT5dX3HyLKqO7hzp9h9udLvMKhl/k7+312mEWFttV0jMof8aQ+UzEzoAyB4SA2/J/Xycf
NjL1LnZtZpUfuGwwQ7LBXTdLf8ZWX27JoRputeqgNTQUWpyLiNxw0NBiqKGDQ6LSaL/EFu1F4Kol
vHkmonc8kdrXzQsFPpABMVqpYka/an7f0a7C9exNdkHV8cPaXlN/1vKW1NpqX4JFnM25IN4eirBw
5zrXhcG9TH92Jzq+uFkakfpXh/9gxHDT50p4QIyll5P9hJOUgEw30l1N+Hb3DJdGkexw56aNR6wd
/IUWglQsZnNXIp0LRbmTMTa3QoU3Fe3FbnAowTDSeRaofy9dgg0TuM2twXVHsmmbjgjL/cmcg+ok
JsYPqNYnMUVb9yhyS8MIkWvpA9LrjWDrh27W3gXY8MPPA+zbi/xgWoondjMnDpbMUkqLIArA8byY
oFH6/+WNjrYFrFDLqIhaFAJHB+Q7aMN3P3gDgwUgvgZlTsgY3TJniABpua3RVSG7hHXvDigzdTBD
BpYT+3fZzsg+jhzSdwvgxyX1JcujxXhtZVN2+Vl7sbqPlzyvnIcxw60BedP1SStSE5CaWCFeeg96
UwAdpOjXTSyQGic6ySf+GhEEwMr9sCB1txtpqDqkQlXM3Rkq1+ClsGVOeMsZqcKGnJaU8yQwGU8i
hkyXz/BSVosUuBzuHy1+vdS8El842+DkUJ2vB0TgEOfn2BhSmOg6rR7XJdF5Lw8MOiS4rTKTXxmN
3mawdhlWGD8Xg1VedTFxMOli4J0ZGnb5hIx+eFte7LSTH9i7LN89iSj5nMLL2ng9Xs8viOILhnS9
5lHgrTj7EwhMy9c4tjugwRtU2jaNReUJPdbFDnrghdwxlM9UQc2bovoKZpYqor/S/JZcVtzFlZp+
hAw8/Nyft0WbV4mKUZzcoFR6SSrK3+koEKtiNFfPJ10NIR3cTJUjZO5pfx2cYa45T6u6my71tpXZ
Sc8oj4KgNjehajRm8QDCRDSpXAQD/8nDBEixTalqyy22srWzWdAL5NAAsqFjgXU3XqETWYWZ1vdl
MVLd6aHIlxL/T+N6+/0T59RkA96cXWEIT4duFUJW2Yt+iRECp2P/qYjL1XCudlmECbhzL91O1SB2
DJA/uVs13uZYR9lnx6RTZLiDnWSbMn16xAdh5ARuVyq3n9ArwhhyCDukrROBfiiWuJ4y2++cClcv
ib0NCRKpB4UMfKihkCUcYL4Ua1Np9yMdQSmSB0o4LIcfHTSdH2yvmEmebFrb2nyJKPz+mZL2DhIw
RXxNDutu2Qcl5cdLdSm7EO+IfbJqUSwV9eOsaqaH4VY3jf+0yIV4aJ/vAE0ch6OE0LHYX10Ew6y5
4dJdc9m/KjNa0XHlnLuCaofjF7l+DJDqCeVHmX4XTYiXeNcpQzVHwmvsfw1Y8jDZ74wP602tvJAM
THnAUmiP9KUth/B4SIVCAacGC4UXNjYjlTTx22RF9/IJW9Y9qkJJ55kSpvB88iKfIRQ9+/bCTXSl
QnydN/4s9eJnm9Mc1H1wmg2JyNCUG4nYpG8QDfAxryVnsEDoOnRoxG47bFrlVHPdc9alRz/D+ATU
xjSTf7yUIaSH66XZZ56QwQlUnWrAF/X8trOZEZJPDtK+B19qJG+B5enrc0Y7URo7f+f2LhYFd7tn
TowcSBWDUAraSW5Bz18dBDqjU3pg6kGtIoSsQxOywrbP1RhAj5e83v3Df67T0UDxNPvJWD+Co28n
86in09ADnFgJin/6WhPhafGSATpEAd1dZMKpYqC+GlH/fB4Z3T3CcCC+lnne/AkasPPLRFNqEKZ/
VMakfyI5MDBxQojG1+0kIUvioeb+ORZd5U1eRrrSqQMckh8nBxoLfqxdCajoWdrjdACwmn+qBfH8
fodo4WrMebdHrDr8w72jNN8ZSLdS1gHHakxLxMLxJ7JbJsg5GlC9JlFJEXrnWwJAujiywivdi8Cx
tv1aeLUUtFA02wBcyzA4ZhFOPeZXLRxWwMu6bHLtsv6pD9UMA9/oapky1HIKREMyc8blkUcR++2+
b5bXnf9QE8fXZE6NtwBcMBNiI39xyFKEvgWt2uGOYbrOdtxACLhvF21gMjNJ8yCFXFKWIZvGQNW5
LchT1yUygfeUJKIf1Nox2F/SS/srKpqL67MOkcw17GElDbdMAk5WIuDFaSiK6IKZiiY0zSbFwEq+
yOSQBuYUN/yjOuRIm+4bSJxe/GNXQAYv5BsFVSMq9lbP5JEw8IQ2EAzkIm3YPN2KoU/tP4ugAS5W
jnh76jHGsl3ffHxJrDdjZtmhSsfs2RLVE0uanlJEpRKMK6kpD5ft7a3E57rdyeVjr8R2YHrgFX6R
uw0gl777JP8cWn7zDlqSXwY2HzgPxHzLIaIIo9ShEVa5qBGjyeBDvXucbIr9irVg3qHEkkyPYJb8
BrznvME3LvpSVMa3iLf0P/p8ia3COPUdt6XUaBie0w84lJ1kZSG2Hgg6D9mfIGeTBueoRzUlkZZD
HK9WmBVKu/ttdrR1m3mJgpqIGVE3wwz2vWbjRsSYd6F35L6aDQKMZcAXLY95AweuLmcOrcyR9Frw
ylPOoOg60OOLFpKXkQ9VUKZdhL4Ep0TphT2y/Y7NSI1u+B1EFqTVjOrJR9FhmoQFuLeRqvyPkSB5
999r0Wzl9RhMq3maBFNeJdfMG7Oax25PmyRqAMtPUwd/TZoZRoeCHGoWbrvw2DLJF83hh2ju8SEX
aMQdTz76dAP5mHz8YoOTQAdaC7843fvraj5ZdIF6MdpNqJIvxW0YVIO9hkRbnZcOGYreyyCMU6Uq
vGCMvK6/8c8GJRUChiOrBLRIqpwaq8ojKZU2GeqlUNxCQtHFvxhr6l52iHp/mAiclOsEJB/TbLK4
sn2F+tvtfKnPUgC8BL1oByl16g0pfCroCKDtRJzx7eNK4SWWqlSJJsq1eUsPJlW19x3HkcI0G4Sd
TNzpRdAXncJItfDH6r83r0MOvw1HSDoI2gcpoZ8/2CzQRS0RwA8KnbBTokzMQaq+soo46VBfAbZF
mLO6oVWAdkLAhOFn/eKcluDhRLZeTS1xLx//phWt2he0UyJlP9d72XXzvMBzO38h5i/j3yQpxpIj
sOk4EwqKNXXTlWQuLVf2Bla9RHJW8FcBseSPjgpseA7+7b2e0ensyHczkyrcT4OCaLrlSSBjVTvN
VbPOVSOGXwcQ/WB8M86Xtai/3EGFJsJAn+ae1Wbd1d6R5HIv8T0g7d6CVWP6L0Lda90/RMniIKqV
o5MgCHKQUvPObSVDO+5+j5waMwVFxqmKxwKy6smQ1TkDK2oStR6Zp+lsG3L49Bca0IA+9+9+Gqme
SIqlepeKku0qyzk5lqEMPOVlt5WFL1F5EEdXbvsH2sFbG/EgiE8wyD4ku4kF94YKOQlCPo5X8dyJ
jWiTU/4vKDYFoPwdbfjkoaajqKc2tVaEjimurEJ8vNR/2yzbW3NUUk4y5fknTqtbIHx9zqsuwViR
+71ePuvO6c3so/D62/RVD6tgefhRvwifq4SnZ74hs+v+PiaQqMHSM6momRbLDKouVM+ajRexpyZy
519d2ied1UDll6kgXcw19rG/sRWGxAA9ivuYjg9wmIFEKrC/71ZdJ2wi2bnU9gukKvOjeEozDt8G
9QA7+zTDcFQSX0qQbcLdcedWTGgjwSS2XwAREDWyEi+EoxptPKQsNGLcY/u4T5udzafgUP2dt2X/
uX9qOXdNom69G5B0GxPeUh62nP+qImac+ujTuleH4M2pGjUVYQIXniKUQ1ju2f3blR7dsliqGWoc
eN7LPHerybfbfKbJCRW02l/WL5mIIbJlW9HqP/owr8tFi1nap6bS/qfVd3hvaMANcFciwDbyXhfs
iiZThOcMJ8gdcCdf8T/UIQhTtIjH+ODKiq18TV3f4Vi0l9xACFbOGzZ5CDKOjlqnvJ5LaMCXlVYW
XTq93E2r+L4OJsKjA9+hJAYLdL/Jam6RCjw2X+N1KzcjKKNm9ixqjUCNYvPXjkPD7OSJGPu5vozU
BIA1+TbQxj6oB8MnNUIeBzvJJTl14nqiHt8yTR2V31UVpuMDYFQiaFpqhlD0oVCl1lJfDNHEBuW6
+VB1bwUXd95ObSBV8j6PFUfr57RiBZXQrnTdDJDiL73R4jkUItbz5qiyGVIFK/QsLzgT5AcXNRXG
UfLdCU282OIlAovI7wqiEktHHTVqdMk4oZ7BRRzFAo0s3O4Zw60uESrtgqKtyFmNOUtSh8JOl/5e
xx0kIBK5OXhjmRA6YgOyhwO2U8SGh3S3L3oaeM8tmxBTJqxx/ibwFc/V+AvoO0jIqJ9QH0zwzIuc
Nd2M3C29cyYjx8DZacU6ouZ4t0RN31OPzus0crHzvrMAXojZi1mosatIV3L8pXQMSiDvV1+907dd
HV6hiBlBvNA1l39qBe67MsW0iPT2jTLcxJgjj5PGf31Z+qpHcHBJCz4vR+DPmNxcs9d18BDeU/6T
YpIUzFTHU+JbMyzxy3lOfVJ0EuFwj6oQht+QpjKOfxqihQDBqrU7OSEh2U0zIDO2LwzYWG0Vy1K+
mFiQDpO09Q4Hq2SCQf+27f69Fq7tczHNK4v4o6CdvXHChmkri7DMhw3gPPUv0wAcoezsZgEYdoF1
xQgojB7ts6meT0Kqj/0+8gg7iLmVwmfvmziw2iS2NHV1FfJA8mn0Xq3lzwpL5A/TofvC0zJJk447
SYTp2tGjUA+7wxggb1iUe+hwPbLCBOyoGgEjYbY2rrj9kog3LoDlGdBaAhzx23j8RkKoOltLsscX
jZvCOgBwU5Jp1aH+B012N4VQpzTRX8NcrMwCYQ7DCL+k1L4u46HgehF0K39hmqUWcXiRYiNEzexi
cJtgBsyyNjtN5KGO+Ou1ozq0kCg7H3UCXNnuGbcvto35T75Ij1UigCIl6NkWLVe1s3w/3vyycK6w
0CxTGx2Cj/Ge7JUxcavsAoiSTHacc3AoQSZDzNgcVX8I2IsjGLVdjvrkUfIphqeSufqFI+MEKiyW
YWi480+FJkJzOSjvOm0wIzsdli60aKFWu2KB7FiLhfbFeodgfQRGg8AB8zrCEjkCjnuHLjv7+6Z1
KVzzt1Vgh0diD1euyBfw6opteRchcHOJvKX+nB0+g+ekpor+mg1ys0Mjg9mPrXu3l2o5dE+vxQvc
mozKdXhhNFNG8ekX1hbBe0hVCMuN4/+XQjoxu3PU+6JKs+AQ0P+gA6a454saPkvOpubdOHgPWCfB
8L7FJ13ifCUoOuVyXE+bIMv5345sL1njJzGTnmlJ/5q89nmZk0vn3PCMPzZOykPcz12HQ3Q5X0V5
4leakExEZgFeBXFHVXyySlrsrCX62/B/4f+N+Ejrtae8xxFUWnnuj+3ZaLXUTB9oa2+kUNj0mYhU
5ralZoYQBa2lL1i/hDkxthwwqrZWDFJXHpJVe3KQ/kH52XVzGw+1RHQkBB47lWfADrUAXJFHHi3I
W4tipsZw2DsDiPfdXboxpqIWxwg3flsA29bshD6y6kFUYdjRs8PpKWKZ6jJhxhHZY0nLaw3/g0G1
ryI7BYzyh6s9Ek6HvrjIzIeZ/1Y3JC1uGQhPnTBJaKsAGx4JNm3JrjxWgLumVS/jnafMYuDlsyqm
Q5XF97Ue72phI989wO88KdwfGPoLnfvxaQ3oTxdvS+VP4vB6lPhFdm7h2IvaD4dKxRFojXzEG1Kz
YcYHzVdEHYHWWpkS6PEPvgiten2Jx1Fi8c+1QHgRqEazW89OSr4L6KESe/bFxu1G0PIBYYtp3a0a
OR42mIuph34GV8BfAEeoFSrOSWlCddYBbecepXa9X+TRQdIN0nTpayfmWdFJx4epYaezXPS2nIvu
l7UJab6jC3tYpr8VREG4yh72BkRVXWjV5WU3ZWEBTfwzsCAcUjf0wn1k12tsbGVZ/Xk63qhJ6cyV
5BmiFr4jbcpBzuPIpmsfdT7qz9/DhHqPTwdDiM0SIRz9iwIE7DGnD3xTHAg3hLkxIgad9at4dFGJ
aRQ9QJ31bhaRXmrSqvFyQKXfHt4JLFVqqICBTkSRZ8CeupelFJB20oFON/erfov38jvk61VShaUW
wqM7k61w7MMBchKpDI1EX0cE916M0Fb97Uf/hrtAYxZq8zT7jLJOuUOrZs57B0Y40g0ElgBWwqVJ
Vk4LTypvv6sYfprkQHXZ4flzucfHTTwKYWX3m11w52w886jIHlrs3B+X5pIFRxEbrxxyRuTPuy7l
cVLraBQ2oRhvu/Esv7vvYG4cD121S1TKPs5+sa1qCasWokVnIV+Oh4q3hG2eGRbUGjqWyDE/fLwV
c1uWI/vkfv4cQZIIIktG0dtc7Wv9ZjRNVQtMw0R7d58T32qK4HLoa9oQKjRk8rNvYYyyQY5plCoA
ZGI5PUabmYUU8g0CalAY/a924b9sOL/eTbRzLl5Y1ZiGSj1BdycpwnJLz5M1iGZJB35pQqskprh+
k5N7MjkzPObE2U9re5GRK0GzJHNvCTnwif5JDpTa+OsGlWfjj1VzeSu7yI+Z+JmZJhWHp0j3i+/J
n0s3AMHnNVYhmcabPmCaXBUV5KyJDnyZTxCA2LW2MSNFRDQXeLE1nEPmzjT4/SW2yObQFrReh8tC
ydhGyXRROvQKx8Sc0/VeD4KTIV4rdyVMWSG+QxSGGEPz9fB3ktkYJ8m/koJULLJ07rJoR+9B/dxE
YaNCgNPdRyNaldesI7qvHuWJUmiOqbX1tOP6RYiKIRWhUTkWg4I2bdjJdPsSVrHpyvOwkhz76odb
N9qqXmzXbGZ8Lx3K/mLvomdjjjpNr92JQWyL5In+ycQ7Zu/A/VaviDV0VVoxQP9aifPP8X485P4S
ZK5QoRDMIKPLDpgefnh6mao/+ep5gm/VFtO5ItzyD+XtmlyP7L/dmzhyehlQ9ohBcATL4EF1Sd/i
KHHzqXU6dWqJAdQL8cCej5J1v493oXbcKMIG4tQiTLYatORZObHtE8huFfqpn+wde0V2f+KmyFa7
8+Xu/C5CrL67DRlq9kLaJwtMbc55hAbY3TMY6vZDi4vD/Te2WKKQZMQQIOcoyDJ6hq2JtaqT+ejb
NhPkanFs0KdhbuYOQHLG/ihYj4KyFyGmh77UFJ+Bfp92/HYiOKom/buWkxCzEKk+0d2IghLdP9hD
ZYjZMaPmYAHEkWlq40RMC27lYLzPVY7NQ5gypoiPUZW6NQcCZvFozJxx2pT6rs3Tggq7XhXZzr/U
3I9nrXLzJJcJ+JHzB9bwJETARwY8Khweono///vsKr8zBGNorV2uTrDzPpqGBP6te3yO+QfRAMoO
z1uIphogebCx+p1fxDGYVlKw5Ex2jZas0hG35UPLJ5igEvJlGaXiq+BHSAgLEMB2gQfXKETctr2F
7i1Lo7ASOFIRO6Gvi4oIp6MyrFy6MB9ayQAam1mrWuOuWNOK+ELWR6jplHDRF99G6hIhu/Yb8kDo
8Le0lc/RtYcGaaWkO/7D6K+g45fMXFu/0LAxsou2LthmTQqrD7apmsKimalMd08glUWJ+++UP80J
Ngc+36iwDcJ7+pseAgtxT3p0/nfup7HZLz29dNeARgVC808FohPJDgIQiTXz0Uadyan5eFXzLHce
PBzK17nLtLFCCYDZ0ZYzXomKkCSZGhp9z5H2++fLhqkXKqVxEpqPQB7+ZQcbeb+cHmbT3Y/LhqB7
+9nBCJg5J98OXfb9HEfo/vqs0fuTOGw2+HXaFZPPCnz7DgvsFXJmGU+/hEidiil4kUkGLP9PSFDi
xEcm44vkHIFzP/cD+RAbMSH4XWtvyl7d8Xh6rSfUBjIN1b1V3O/qImr0DXxkZ62TsdxHd9Hs+BxM
UsQcgDGilRD+D36Rt5CVYO89RPdVV34QF10w1h9xH0n7ASLYNqTR4Ox8YngonUCJua1LWwBgCoug
u941AV4qSk0aPDXA9MHTgDlR4LMO/wJDqlhW/68F3X0llQ/W/4OYjSWTSNITzFSZiWYt1PR95d6L
hP40H0hEhj2OSv3SMnZ8Lk+ZlA5QTR6/2MTq38CcHtK0CZ0nPyi5mrMMFKCi8dznFvBy5OBPY3IY
nQOEDQO+cJ3ul7HgWlgypxfFAA+dtIPBDMupGSfHhwP4bYLC2VXL32ARo0+CRKi7vlNZ1lgP2Vos
BQAm4FSVIwps5QKtoAJBXj5RYrdkyfT1zqSTh9NeHOKIBHbyj+4e41Df6NC/Rkuc6vDadhXGBRN0
NIVvQdi6uJpokL9+S0YeBSQFLmjJk2n99GCmO4kxiMrZskdgPblBBgKtmzlNWR9LhO3BaKfqFo5v
uqEKBc8KdlHDPytp7xbmMedN9rpn20D8xOJHBb56lOhdsuUKyd7Y97qE+EFkm+wott3QcIEXK+XV
yp8eV8MW0XhgXfUxhL9I0XmmeTNcPA07M/fer2nHMHf8xEPyn80RlUfOXFhVInKVrtiJ9yrRVwNh
HPlQOBZH/O8SxIvgJ1srwBokyN2Fs8gcrimkCH+hlNq5BVlOEOFAZ/ooEQowfHwoTW7FlJOw0Lez
6/XFNAwqLFwtY0DXwpfvlB7aEgKGOEhVKvSBJ8y45J/5CLwGecBg88FKB4bc9PMy/2EMqiN2Iqu1
N4VtSKG0CjxWtmyLo4mcz3fRJfla++fTodHHlcXh5nsTZ47n0PhdLEtbhqEtJq1lo/Xb7fCTJ5yS
v8+N7dxK5lMbgmuaGErG43IYCi9SZba0NkEY6oo6NtXY9G3eS66RLcsEEPg1/B/GotJ4jiz4s+Xo
I9HYk0ISNHtznN9l5mBEdJvjpLjMTx10b5e902VTjRakTnqB9es7dH0aKPNGN+oMkOivP5DcG8ZL
/qt3Nd9wB4KTHRMJC6oJUtUsLoZkrDnmSA8PZ3rv6qSukQ9iejHaARrb+wMezf2a4N8H5MR2s4lN
lwDoUwTZ3IM1IAEfnFvbWFmCMmae1GLZcGlCqnM3Pgzr69rNp9sbc0urCUxfh3wcPJGKCFm2bSXL
wbjujQlzGeUQIP54csA3pEvkfkHFqTqSwe4ioygyhbZrGbpbR02wwvfNgFOwRQQLI1GaY2I/AJFh
4XeczYGMwkKzEHqb4hY8FxlX9bV7H/9ryr8x/gwds9OMxFRPJeCdgwhEfiwNaFLUa9+SSNWneC8s
bCQT6jzcMQi5wH6hrr8isBc5m57KdKy5bz2+JOuuZIaTUP80VIk3RrE7eoOqFFVgisbwA0gIrUbM
3PPV+s214zWmT1pg5rZihfPCeeIj7lewYhUcm1noKeEhanhOGhb4PYdQocZQOgKkHW3c2AymvfTN
6Ww3CtEyRkNpH8unLkPkr7kJLjvRy23DBAvNKhBjtH3erMQZU2TaKIpzLx0uOwlXDuWQfzFJXhSG
KV8sM8yJPrCjd+sVu1YmZmdH0++i24e7LXI4k2O/jsD2gpPukXcmUDn9ruoY20igNNVxzWZid+di
VJ7wCk60hEYnRM6DH8EWaM6Kt5umlPrzyeXh/OcF2j4dgC8cOuOZpKDjbIMcIAbtM/QJp7ED65oo
1Epb+HJZpfmP8C/Sy79C/4/73QxnbQqjbVmv+3047td5Vgyu20Ni40LoPY4s4d2YAGudT9t7ZN8t
VdDoc56fFOCxZADLQr6//1pby/YIxyxKVHsQW9E4eVTTxu3aveSj1hN4pt4i91WB+G/xIanSkt/r
FwllO7PmGBluu8uEwcFbWTINb19cmuTMRynA2tt3wOWvlSgy8W0dQ2nHX7CWCsXg1Mu3c/y0aTNA
RJ4diHzRSlK3scfeaML0+qpmr8uzpeUtpALHs8u41S+8qJZVCWhdbIqOMUIz15QrUSSvOGQ2ELXK
RsGSGaER/N0lqjv//UG+4E2wVnQl3zupmF0b3bF3BfXj5EKGoZN4j+EC21sqHnfYsQexwohAm73d
P1IUYorFcsuWneLQnJXFR10+IQ8IGIrzYYQDmkrYFV90lOu55oi1QjYqBENNKTd0xns72wCQwOh0
d5bzb0MDmjkP7/qW4FeTK9DiyN2LK43o74+ALIM6S/B4/XJ7lbMAJWL+Yoe8qe6kM6XJWr9UILYE
XzQRktLpRpC2uoPtpt22u59/DggGBFBELFUd7Fu3cGNFaOphkyjr1JLcw6KdiU3LyKGHDVujRKb0
O9LePlgt6WrZpHogp5eL4Bg+7rxb/mNh37U93AU3MOmlUlIgaYAQxPHowMh/YlkmNJJgMNpvRXHA
TVQ/Rvs61S8sq7iiPa71OR9rhISEPdIMVv0CGpYg5nMsxlXSvNZuaMf/WtQHpX5TKO5Wve6s+QLw
tx24yGeAHkmm/jduhdhZIHRctY5d/eugxD10ivU3EmfeSIi341/nCN43D/aortfog8/PqG+rj4Yb
L3LsRZr7InkdhfxVyXNng5KFH+n4+F9fAYl5MIliCK8yv5boYVJagv4AsWqLTY8p9OmFN2RXC9d0
Eh8siqKhZgv3EitmtmNuA7h1Yn0p2Ksll0afmpMHQ+6HTEeXuP8DeXjOTXVrJJduc0O6xkiVkqEb
mfYL9HuzSErWvixvp2aqMoCOm2BHaibWAaa/yGWdS0ZSK84+5C+zmhVs1m2+J2A+wvkHVChWsgPr
/vFSJMJKbWeKUzWFijlHr45E1/x22rhGR+D2y7bJEE9JCfiZVOT5SaJtw1g64jCkSjykRdAT8+uQ
fWF7F4KwlPUZRZzjdi5jGII4zt7tjZVSEvFmoZgDrYrA2zHF+lT6/emLEuFrXYN9lkbLf46pBXyV
8ndzTrO3TbKRyapdIm1krk/zL6/d22q7rmzUeT0b11QyTdkKsX+BNmZ0fePihu+Uv5uHFw4BMVyF
fo2uMoFBXJNS1FqQkV25JbgAuCmm/WI2J5ZsMc+PmzT0YLWxP1qmt0yN1XVuDjd/jLfb33Fs8tk7
bWm7vJkiucGtDPGIIrOG5kn1owmK1E8i+yPli5gjVPndnvGkgHAQESRRNIa2G+mr0+ZfY8hlusti
IQOAseSON0BKjHB2CD+3GIJSvmI9RmlU9FzVzKWn4MTNOVlnNSSG6N87Xz5y1st8J+DzLYEuXOaV
yvMUpp4NH/OYYEmBSF6U502+mDO94SV2OxAU+MLm9eeqvdmxoozww8AcRJO+lw9CFwv9U/armGFe
2THYrQeX8Rsc0m6oZWqTiqAU4LhgIQSYkj3UuDAYc3KDX9nWmAsxiHubcDtQTDej7HAcMiI1PVGH
1HUWKfPtvU7pd3M2O8RXHNCcBPDbRUqPnRQOKEDeAIeBWgGyM5OrV4d/m0kUWjFIgsWRnTfZd2jl
5NHlDKRhtygP4Zunn+q2PFILiI/k40/8KurahiMDoWD9myfMlwfyIGVGTHXT1uHyBR7b6/aOI8Sl
qxJYTBOdl2dH9YKkdn9g4SJZ0RHowG72/GzY1vaSu++zss9LY9QlvB5ecYWtiVXagfkPwmJEx3oC
1BX2UXOSOaWIXck9Od6qIZFYhln9ceewtaL9yH8tn94IS+mJsvL/2ntd1YyBzcvxMEmwnGVVWBhl
oVX6yJJ9yl1JUrLc8Xjfd9KFwUFREWtIk3Yrq3oD7Yqk3yloSjWvoLkYm8Bnv++IO2As7a/068i0
hzjfFejTR4SvMEGFmCDM9f9MkBnhFGQKHd4MnPAbEPRYQI7AGl3+T+VnATskUYnYRR3C12FcYc+U
ro8f/tj/0g6IZZ6vnSbGLEgwHHDbNAOm0/CSLMBUc3s6cGfI6bAtTL3DbEzknilW0Hk+l1D//6xv
Fq4ZXgGhVyclMowuHiD2QtokuaTkc90Idf8lKPoc0OB3o7ba+bvp8FdYQJfpTKLV/M2R+RxIyIYK
murMOif5120d7SjwR5aU4YKrN7dxQjkRMhNp3Q1VX0vfoIrXMZbBwdAkObjOd9qeattQovQhZTB5
lWwfGnl+f19CLkS3+/YQbKPCSpffu1oPNRFqqCqT8P0jjsgJutGEAVyrh4V7UCgJfK/y8CKxXO/W
3LpMUGTQrfATo8rcUJ9rxvIE1xnxA8CM07DEpu3wImDYfxx36obyNRs3wks3YQ1PTtyo7y48YU25
RbvzM8GiU4VTy+we3hcAMICACia+AAG/r3fOA0GjybB30Pn+5fkmWaUmdP/XO6qIzriuHeaXgzoX
2eOybQVnCTdJser7UkK/3sfrEk4Hc3dJsvpM9irXwIhUwFCEcbsmPqesZHd+vW47Fry1C8bD2XOm
9P+eCmuVcJHrxMb9V0i5geyvi59qQlYxn8qaEfgRfhtX8y4h+VeU0Ag/O2NMegPOq2cgiorso5UH
5SWYbCyO1ZypOmrgH9aEBfg36fqTdQs2+FR2AT+JF1edJ5l+sdaoudCoGaHmVby91Kro8zqB2iDX
KHqhmo+M5PHjU4maowu7epn7U6sEk0sfmpWIyPm2f/YtsgaxvaNsMQbDfQk2TlLDalc012AXUQ1P
3zF0y7sKnFwbR5mthRXUdfvemf2WRCdWRQGXzVszVyzPHtaylvmmHL6W9d5ZT7IKdZn1h+WLxsjc
xktfp7O/yI970n4wQAWwkx8bGXXGUMNWP1KPL3ib5S4XEBogpKuE/HR+agUuRLYLGwtt0nZJQmm8
LqBxQ4IB1A8UKpzMUzJTCn4GL0pky055ZMjlsp2kAvyZrxM5NzYsTS/79Y228fhXiNtASStJ07hQ
kKNpAR2321XQqttH/8JdMdddjLRDTK8Fu1h+DJSqJLOIGYD0UeZ/kt1bTQN2CpDAODR8l9No8Lk8
IMpl0kCC81zQ6a/Mq0ZSwvEdvd+QAg1kmaen26/PpG4GEzrMkH95oqeDx+dIwYLzfnxmjTcEibJ9
n5ltdLEfULN1qbeEI/wEt/Cqo0gJ5KwdM8Tg7y+QChphq4I/heaTQltEeasSqNlbLDE5+TCJ7wCj
gMxZuuobVznjK29lUj9iK6EmGSYb9GIl2uhoojRUi4YwrxtwUNvV8pzblviPdHWqYh/ZmzCsH+sM
t2B9xcBqAJ4CYqmUcwRhrAuIOfKjyWw33fH4B3g11D3avj5Gf7G9ZX2WvNGtyDlIzFV2IfHNxPTK
tajtLLSXzDbxtiKn5TMm9L0X479A8fueSRgatFlW7U4NdDYX9kuj1JKZK+t9dvkdhWz5gF9pwQjh
jNB2IJtEvw3UG8gT014oOTM1G6Uh2uNQukKDjjhhExW20vB8x69xuPzzFuGcud8IXzqq82GARncw
GQDBbzRjLUFpozzQ492ZpKkEqLgX//vDkP6VIMqAxl2z0SjoT4Su0cpLBn8mGvDoeSCpqM7KdWzs
lVbwkE1MeXr3VlJZ2gx8SUJ+ND5Ywp4gJAbrQQUhzbZ8B8Bf5n2CF+W1BfCncbQZhW+KA+3DnSi/
FLM+g2LWFXRjGnRr16a5vGuYtEolqD5QpZFhHZdw9BYjSaxmdD4Z5J9VBBsTjAIy/ktM+3sbzFyj
xyf1GUeO0dmnvw2Coo0M8/K5qNQBKAYOURui5hQZbeBaX5rXaPmFPIiXY4MK8DyyWur9pd4FjvoI
eu9Zr5ijf+S43e4BgMmYP/m2oVoWIEWZ5cjmUfd7kXrbii/YxhItKsKRwhlaU6UILsB0YAjOBcPz
YtsoRYEo9+xtaFgQE/xg7KDOU3hYHBErAT3k85hM8DIzjf1a/eSZYotp29Jer4dqtWiO0FLbDP2D
UB26qTsc8HMFlOxLOfyafGyQ7ITIiMiSF+VkRPPw6o9HMrw1wdQKuNi/EXndhTxUyukNIKaQKT+r
4jzgUi8jM3ZlK7FmitEtXZc8GeMRDAzb2E12qfx6/M5rRkUaXrS0bOEckQcGp4VkVOAosC0UhU1s
c9J44VZSA7sqFKOurP5AbqyxvBcX60IaTnNnfp2yp28t9NKzk2RqnD0jUQatoDUtsmabRpbwDZVV
+6RhSAinhk948KtlOKh4xd+8dHaW3aO4w/z1rq7bEJxIHfUm97FodsDukSlc66UXcAHsagrvlXrd
OlgSHb7GIsSL+8n21DY7ZcaGL+FoQHGE73zd844SOJeKBAETYdou+nDuvhjKD3q6DppjIAP+s6Wi
alb+2FnUCSzucCnEXfBA4LZRgcFDRpi9XGd8TSjm/P7vMAk6h2AQbkdraVGaN9ffnCGCxAvV5EOs
LU9fiKnKhn/5rf4hqzBABoKERFaUbzVosw3epB4/eKkGRKg04SpQRmCMF2fefjZM6XJxMGzMYXQk
e9ufmS9c3n5rY4zOaBl5EmanxF0bTxthFUHxLHi75m7xwLo+rq0D1BM9JRCjlb+3I87m5cJpGnKo
4/zsMmAEypDdedKUivO1cjWxmGVoub8SBdW4meOG3MbN3abatBYSFIli+6KQa0cR74MA8PZm4bp/
WMkQsdsDX5rnaqF8xjDei6xXBGBpS6f0aEeas5RGse+nIcz0db9n5lkMx0n+BdeIDGgVNGy+OA1E
q3NQfFbktw6SbD63Ab7sLDnWs2VB03RnjNcrinzwGl9E0tkqtGbFyKtRDFsGD0eXACfDPXpzoEwe
RuKcn2GQzkiSflilfwOT80MtPDLrlXOtxFde+HfB94aAiOOryfgxttVBkYDgW0rb65XNrPWvLMDs
HINsRo47w2nKcRFeAshIt4XrmY+0fYJB6vvvLihVUISeHtg+9edpT5QNaXcjIO/dJGqdMAuULzPM
cpSSm2h4i8PsxOa4yArw7T+qMWtAN8XcATPeXP7wELsstV2JCUs1uKz18Fduo9c3oxzQB4og+GMM
2bWMypYGfITuUkAQmuclG6oopdBcO/wIbW1HnhEC9RHS3sVyYzYjsWSn4P7ro91r50RCgcJ0mUX7
Pxb461EJ15vNgRfjf5XBucHXbUQOBSTu7pFvjmV/vtGMr5vRFwZK7kuKCCYbeHWLr1K+VJbj8APS
NWzjlmWR8p7ZnGiSYxtEJ1DIyBoUnGrDBxhPSFf3z+VxkBoD1/NTeqtgXXfOTtTnb2vSNjqVOaHM
yutxCGrLlInIB3NKpeZLX9Az32k3MeRaEv+G2ZI7G8Cd3KsHmFqX6aHfL54bGMhALWNL2c6uPRsi
Xa0MI3EKuPodfNT8TH8z0vHfYVW3qn5Z1AW0Ovxjggqmg6McoAevBFdXcgNYy/F2wJn0yZWhDE7q
Y+rrTALLSK61wU0TbnUI4faRQ0ur6NG/IEW4TB0fQ5STSsl1SMDUzKUvd4DqMNrYkB+LWQA8A5PU
RoTCLUNNo8ElP6glM2f/535kiV6SQldgYvO5suoXeR95IhhxT7UvdpcYotNhTRIniDnyP8Nq7V6A
I7/SMRPVe1ro6WtpQ9jhJuKgZh2HgcIBfOc0LMVlLK77v/TiCp8AnXQgPg50zZ63ADG1AwReSILP
GI8JZzbLusKFcZGCQVN8A0flWUP/V0OyPwDr+GDRpS19DT2X8bWQ+FPR7enP4kQfkvirdnEuhzpj
XNgrYjXZLgLWv3tA2wv1mFHXIp7l2jP6HtoEXq7uAtNrGQd+LvyBnmxDXK/ZCmRMl9kP6VmfNV6Z
bMzRei1HTjJXaPRq7MPXodkeqI9uXCYyK/MFRKdlGJdnN/vSZ4pTM/VSnpezny06fWvPylWGLEfJ
XBREaArVSc3g2JeCXBrHA1sIR7g4g7XML+keuCihtuDtKjVLGRKDDlPIHvtX897VbrSBck0lcm8m
1whxnWz7vNU3WSyJ4rk0c6b/2Rnbptvtr3ZBTEqx4PtLB75wnI4oIPdF0Xz/thfdSqmWbCVEcJDA
3yRp+sFn5084jI2qD1BYf5fmRfD6b1oAQa9mq5Fl1fBK/u+6TV0fC7fAnBUOP96we8yfCMZ0bWgF
Y9MM/7FAT+NJY31gRv0lkZsdh9RK5CB7AScBItDvemB2DJrqn7Uvoipxntu9DVuZur9+6+lbjrUn
O1HfvdMDQC2cCszQc+QjYMaV4eSbaoauh+uvhxCeQQFIV+l5BLL0pE8p5ogyzLKavjup2RRtk3t5
z+rtXO0wpdQH/QCE3Dhj5nsmgacyqGvOgO/il3eKu4JOeZQcX6LumJLcR/MDplvjTzvhNm/b8oLb
4lCD6zCYg4qC6XV0B/IoKmseD5yGVHj8OfdyGkQq35mH68zF1/nYCIZd/SbyMkZFxaGeJmAukWvs
KcL++nbSxhJ9V8tVFXrqe8O8vRiLMW9IavOahNBVlUaqpi8boZNgg7pitU+KWFHOPZY3gZ/d3QFG
wPuDTLpkFIeWl8upNkRriNkvfrOycC5gcwoHCGYNFhdp6/pIkaHDX7CCkk8MKP40PGQITndwxM79
Qis4IHhjAvS9NxT3XEJ9R2wTPgZuUU2+UBHN5ybCKQbB9x3hiQ6Bo1m7TarE/4bHxF2xEnUSi/Al
q7gV4AfTdTgthh1MgZmHyjn40NkBwcYoaTwptT1wGrHuF7YahiYcKmuczYXrh/prdfSvb+nOQBgW
d9HejslvYuEexkvtxNr5djOKbXVHcpHa3XCzTVx7SJT0WO75Ue1cVZfQ5H45bJ+mmo4uR9ClWR7a
82MbgERFoubikEodqV1s45hxUbt2ZGrQwgOETw/b5f68uLs7QpcCAmge6Tvj2Veiw0OaezlDv2N3
+TQCCIZZ2LDIsOtfLdYaTczipCU8V7vvPOz1aYbVs+LoeE0FPWpSu+R0O5jLhQLxZozoJUtQs7cc
8cZKb8A/jLnDxiqHGi0OCvclvGD1OUDB+pp98X+6ozoo8F4GGhDVK/3hGOIXXwufGBRdvARYw6A7
SguJjM4NQiY0E26R32WkXqal9H5jcjtF7z/0Mm9s3pfbpieIM8a4daprNmV5faPiB1Dec6d1DWaL
ImZNi951AIaWDoCRWpwXdsnqLRCZ13PVe7teRusKfPXNamSCWSnJBsuB+5cjWHuIuPFGwMw7P/Il
jSnkJ+Sgl55hCuoKh2UP2O8+YpG5Bsn/uhZmrpLqcOmEERa8s0NDlnFnGEER7BEhCWNtvyd1m52V
Q2Z0ZyDjPz21GC884kz6fhf2TGQYghzTG0mkm2qM9Uzp+MrT2YAxxVHBoVxhbO0JRPcw0YcoZJVq
cxMnCun+soL7OYPrXIIQR+YHOVQOcVUV5Vjs7QZWSCJ2nVwrvzyYxBCW9sl6piRqvmxtPvOLrsB4
SA4jcKKIOJ5UFxpsoWAUbywArn8MEJtiPjCLs0W5CFlByIoFPHf7yocQjtBR2cIw+gVmvS3I6Pod
B+To1vGTDWnC+2JGYb9XQB7CAJSW39qNYW3awlnsqM3ihG/+FW/fo4qktD86vvGI4eOgKSHqEGa5
sQLDzwjjhSvoY4QQhYJrYf9FMuNe2Hc4BDkitvbWrds+YTfa9eq5wW7nVF+MqjLTX7zi4He5Da4b
81V9WMDOnTSCO3pD5buCc79giR8XedAYjPTGqgcEDJHTwoimQnLZ4QCBVjlldsuuK/eYQWw4Ffcu
aAlZDdGg5k07YhBzTHnrPIo4nr4/GqOUQEULtPS1OPe3upOGG+aFVZMoy9tsHwZi4ETgNB2ZUrkQ
KAUe+PaEhIZKkgfYd3c7MscW5ODELu4BBxNAtA02aciBx9Sf0ThTtf9bayRTSEtbqLNrJuuVb565
HQe4LHFvolumbu5JcDhaACrnww9xlQKQjVCdTtXwsa1CtZP8Au+fVlleOV8fOJlCCCO801a9EjDa
RWtAY8eo3n2xIV25DGQM1lIagP/eb4t41NQixStqDUv4KSx65EwhDgDg6zp0p22adf3Qh/U8M7eC
NHrPj/QQDlLF9lmTwoZ3bZQbWALMIMASGPUzX6HM06aUbfERv42eMXHGFENNuC9fihe/LaBoxebh
Q8d6TuKg3oPFPYTv0bmVUVZGGk/BPnL0bVP5Y8v9G2LAhuzRsQBRQkSSbc+xGdKeXesNu+g9W8+r
+clpUXZn20mlWkx3Xtwfi8LxaRu+Ju2hHbUYKcS3ez8TLUlxLEUGd4GcmBNfW9FE2OjYxVGZGmzO
V97fNQ7HY8+88HxQR3mcoPR6e1R26KSmia6bnNFqIukyCvplw6l4BjNe6Dkvz3f+hxXrCPCeujTb
PqWBFx4WYMrY7F1SNsdq+6HHOe4WvaOfT1GVfzL6CdOIm5cFgoK09DkXM+BYXg9spBZ9CNPRSyjF
q/MjRV5fNblDP0O5GEvpdfaRJeHTIhX+sPzd6ATnJpUO/BUCrjXQWF2q6ch36+AYAXZHp4tbWLxm
bVNmiXPWnYC8XztzCBh2IC5lNliGbM9hOo5KiPM19xnKit4hVo4EXtWsB4VTinT+Rs8N8uHqIrZg
OQqg/cyAZalXPhWiIDcDnijYNr7zjKMwSdvHvRiuYGWu9iAMfu6ndZHWi9tkbUJ2Au5w2tcQQoCa
mkJPlI+F4KoDt1y4/KYqFPmG0BCwKEUubjt1sXD1VFN6J0/XfRHzK3+nSqCRKWzaECvC2gCIMri6
P7lGA5CczZ9ggySXt4g6VJtpM2upjVZ8uWuHllAw6ogWYl9H/ZGLR9IQXlK0xiv6x39XxqHyWd5R
LYbY6YnLliEt0+Nk/QdIgfQkBn68o+KhAuTGXhcSUYtZExjclpanCSG2WfDogSjuKxly28YyLD83
lsoQ1gjCKY1dml1Yx7Y52NPex8Pyndaw8xykPjVK6ZnnIOAORXNIH5hXqk64WLMP/5jTdS5Iwr/S
WQcmNSo8+w5Ag3jZb/51xdf76JRkj6rZNOV8njTu1OMYVzFW0vhnNfmS9eWGF66NQI2X48UgucxL
qq+rjDuVsD2D2xT3HkzkNmQo0Vwq7U5NUuJV7rT/EEj2nHcYS6sCog10+PVH0DeJpx9HZpxnayrn
1MmUJS7rYMMzXgRcgoWtFDGrBo4vhWH4GkpXT+xr/eAXpNK8BPJ4Oina7lHBG06BOiWpHdABICU/
nVqCzgzmH0C7TotYFj6qOH7tQqjvLNOOFKi8pJ3YQPZlC2zH53fUgtVGAQFf7G0QJRMi689N40ex
wk/gwVINfabUkgrsOpM6V0MBSXSUuwG84NT0sNsmuiJb/htPDlYMbYhFBjzmUL1d2YJpTuax6lV8
R8CCbsrDOAZCRM2gZpRCCHehT2GCT+lyE5vfTLHfzsFj3lNUS+PSccPvNNPei701gXwNmODPBDRx
0ZxDLXtHPYy/+UQFNlB8FF+fo+dTn0RxLQQSScP5F0PIaWo4kUXe8S7UcvoqI9vSxLcA3O97zJs4
LbYl9a7zR23QaLOO/wsWZhJhrYxQ7hbtav6ko2nrlLlcqpTdqKdkQXL4kZXhO14m3o4n9OepeuC3
kKfsg/S6qObZEWX5U6EN0bNL6HOjk7zbmE1h9Ev1ASW1HZXmZn1GSuPy5QYdz2wvIP53fdWZPRcp
3z8xJaS++dWi1RNnPJoMNN9iauuy8ygnAfcW0KMklcCEZaApE8ba2TLNsMadNwwWiC5gHrQxLag4
ic3e1+gfek5Myhx7eWEBSg1pwzfq8Csaqsq8w/DiPsAfcdRLOJgmVn4NIy5GoQi2Vq9lSqTa5QN1
nrKsF9dXVkKWz+wpzV1gy2VlpUdB12vX666Z2d3xlxSo/lcCXhnFgt3CYmZ0M/UtruNj0BRuw1Qx
09m0CFhuYGD96jXdOlHog6xakBHFBrnCwv2KJB6RRm4SZ3mz/qU+YVhCbdOE/ER219NxsigclIUS
yWrQLYD3mTGt4PVd3frFQDgnxI/XohtC9YuqxHf7AhBCDpNSXbprCkZLwFrQOO1uX6YfUq6RCXHJ
tSX+kBln+Qd2gvmmRcE9gMxAb7IUCvye9ydBDtYwVdi3oBG3u4aFw7ikpa+g7AhBUp7jrkDhNpT4
rlbq4K6af6P7qnrPFHLxCZkQEUWVnFatuwWALbt0mapGCImQVF2LTq0bl9C1oFp8/Ce6WCJhJJ/6
tSThuyX6qHwOre3w9ySDJMF1PwZXn4X0ApKyS+QbKPtp/mfBfJz4OAYCaTTKeyV8ra4LkBbq/Abw
F+xV9HgMMtNFcK/b0/DeqsFs5ORB7XDKd1U6XR549SBLbcNBnbt+GvszYA6qODCC29zNjANI1MAX
JxalktxMf+QzQ2o+7V+cYpeARzzHqVkAjcJXLV0m8U4mtnIPy37C1fY5VZe2CzxeAHxW/WYm+hiG
5BxgerZ673HW15jRgL5qnF28F3GzgtcsRJdtbs45NKyvSTaoC8Yj/FwzSJ97GDS1gGXJhOjMikc0
kzeWTEuJDfOxlu2SnLVMKtkZ6Qj4PTbvOTcwFqbT58Tupp2U/Fx/FAH48YwT8YbgQHlspZGNF6yq
joY7WkZMX+1h/2MsyYRgDhtjAT3AcmM++V/DapMpRFnZpTnDQa+PpWbhtva6ZCuV/1rQzdxKSvXx
7hm02cl31ZyN1s/kODHwfSdXd2pccGv5yLYp53DbTrJBeVWYGR0N7x5AGs0eT3UZ7BUkQNv6iBm6
kRmuHlUzmI7xD1932/od1aaihnlErH1FTRD8BbhKJabl2IMwDWv/rIF3A3AiVDADaYn1UNkk/NPe
ULc5rVb7BBe3Sp5PzAdmLUBP7poENtTfw2v5uivnUpIAchT1jeZs56uRaUo1CahgNjM8JKvwT2bn
fRgvkD4ELASOx9Q8bfpACZd4NUAKTDBZ3OLkTocHRwnl0JlX/Q9rfOK8IALh4KGB/vKw6hnO2CZU
4+yYsC23Um4Ypfc/5AAU4TnVapAF4XK8U8tc5w6XqYLuxhWV9uR3zJ4KiNKNmLt7ZvY675xdyTX2
TQgL8LnE941WlwkSNBy5ZQggFbfNukOIBMWg4ckUklZ/mnqDQ/Gjht4WrMlFqDrap/BOYZq1qAam
RO0Kjm/k4g3hxIcma8NkobL4MBSPBViuREEfpjhLYQyLeWChSeOJAz/1BYfXid0OYpwMOdDGaxZy
iVAHmqGwmrJKxSqEKK48G63b4ZYv4VmloE1rqKTdyBEVnS0xxYEkRRYdbrJsGUOpA65s5ed+HC/S
uOQssFdZAIZXkVhhArA9cyrOhaVVznQCupiLnL/Gn3uOpTbgGgJOAaGZ6OmyDMbdKvi7oyua+0Fa
GjC+0JuyxW629+uHZdVjlkg2AL4jTW4KecGb8Fce57H0oqaK5XyRHNHGzdGDfTszrgNMiwjVBQJY
1kzrVx9L9fyAMRzRBSaNhMKL67/imND8p86db2CAvLdA99oj6d4QL7P463CX6KNv5Vyi1yBtYRn4
8zEBtN7zNID5B4hg8LDU4jzqPodVD0zUkdP4xogd4tQeJUXP7DSFdBT4rNAzScnSYEFSmt6WiVy3
MRGitDg+Ds5uXskpuVDgF5nrfkd3BC/Pam/HyjPeJNEAuRCZSky1l09QRs/oQGxT9GY0yD+jNL9G
E2zSZhdsj8nshG5pzDVPwyD5i0Fw47lzlk1Y0T2Zj2NGrVriVfsMJasu+Ts948H3hsgNwZ6L9FVT
dw4jQ1QtQ/ryMMJCZ2uY49/bY9Kl6SV3fa2tgyJK8WDLasy7IeDa8wGuxcDsCYyR2qGFW59mnPez
4TN8Z6dTA6IZjJ9thVFJY6eiGfdVRJGrcupT64zj3TrHxAiWZ8yUUpI5yiQk4f93DYCrkNrchCYD
Yq6ni9OXubciLw8QudWTci0W+f9yMt74SauqoaeXbXhrs2kdFBQS2GSJ6TVEOnr0pDDB9xz0x4hZ
UPgmyjpNmFEotQ8crCSZ7V04ykZnKTEhayKnDzxIkzronKmxEuJeYwvcQV7oWQijTShzSmhOJqER
xI2orYJT448EG1PZv9o7kzz/kJiqCjsM3qBlo7pUbP7fFnbG6aVLwmknxgeKVBTzvZZyk4k75/7b
E6v9716qzrSA+fBx9HYZLiXWx++YaRWjHjYt+0Gu160tFYfqLDh0YKosbwl81bS1vPsJiGNVtzGF
w9UgHt/fM4RKgT0yLhBZtAUU2lv5HpIcNQ1kdU27LeMsm3bQieryfs9PyJZ+6AFPBKEo7kUPrzfE
GcdhUvw1ITci8u2tuTqkV4d3/D8B7P5wLfCoTurL6h+Q6UTjEgQOxLtw7XaDVl/2f8T8etDBUsK0
4EwNWTN+ToCuLzYx9SxB52lPcXdIjJffzAUHq4sVDXjZTUtVxvN20ddC7frbZKeYCvhP2v3XXWnl
40CJICVV8thI5m4sSuAFz4zLGYSS2sklSkJH+X7VP8tPBJBmL6NTSB+vSQhgCXxUDQIjVwufgjOR
X2xM/wBTG6sH9n0/+Mssp7VD/x86rKg06HHMUyjJRTwogwPYWDZXxLibAzGz724gO0HPjiZq2tPX
FX5RzRC8y/Y87wLuNSrrcQsfv02OM4UUCvHU6OFcrI8yFpNiFh6cwzZMVrINdpo+j1978BD5/ZIU
kQGHtr/PGq0cvuS3V3WYoh4ZLNyfGWPyBD+zN+d75wyB5t8/Y+b1XxsXViSrslDBzI8X0Ti9PM5a
6uehrWQO5jwZz14aWIhNZCwsD89P7TmqoC5h+IqhYIPSxO3WWsVhJW1hRkPtHJ6+dULhdYmZXrb7
+w6QrxOgL90TQaEAbQwpdP4frGTnWB+AKylrh0q81Ly3wth3qK9Uxap7uHVJLDHxEdSX1E9Ef60/
V+pdlVIHXCcNt8u5TCmrqi7EQFSvd22sBzoE8w1zk91g1h0dk6A3jxkghmsUObDAaBLcKVMJluTg
AxU4/zE8YE9GA2Eh7GTnOZz+PIEG8d5EnUn0i5Zv0vEVdrcxJVLV5Aravpfu2Q7Lw5AZrt7EL/l5
9s79em0Z029INNRqm9PdRp58ltl4VasjC3e8/SGCVad+paG6FAghVdGQ9cTr5AFYyuOULH1vNvfl
n+UvZaKrQ8UR/QY7P58f81D0DtyUnW/LOHhIAgPCpAEn07u4xJ8fchlLLZlMqbHatC/xdlZS2k+P
dLmcII43+NLBYoQnnHi4cuot+R2FxTuA+PEZUQLDGcvvZLsNGB1V4DBZonNsDGr3QtuK3V7WEUfM
KKEz/iXqV5Q4CYXbZX4NIdmc3b0c57ESl+wHkF3YvE4a2VLXKt+BPx8HY3hMfuHD1ho1DJqY13ZO
kDrtAVTLAjaG+hV0GEBbpxjkHmTcRnw/jbh2sZfbL8n8F6AHKxVdhACi79Kq/a93W8GfY1UwiL9V
SuMGma4yV9anQNublUF78m+L3G3UNybpnomGcSfXxbm5KUaqX2OoTWeZUB9l+ohxUf6KU4L7jZhz
VBSaNTphvi22f1/jiDj7msPpQgBExBtsiGH4/3L0cBmwOpIMlSiOBARKdXuTdBowU9YGeVfa34rb
vYng91ykaY2Dbo6FbniFDdWyp56XyXOYXPorKWyDd3slzvGfyUrxHhoqzqG/HcH3x6UldCUt+Oum
i5/QmXC+WQKZYWkkLbY65mcpy/MaXO6Zqoa95TcisZRjXHlEq036O+4LxmbtxGScFEB0Kut5ejZB
SymDtCQnDjlKkXE7OcjKRv1JfjyD/vcGn/Gsx2ihRdMreoPEUHXWE5xZPTNYxkFX9HxwlX7tk+Ay
XKbx9yo6IHII/e5Mpp8SpwumDF1GOm7Nnjh1uM5U3y0iph6E/tQy1xw1zulGMIp0EcCWT39pQgPe
GG4QSRhv3sEpC+9+YAZp7ZupPA3kjNaLxa+rLDU4/82liHdzkzn6F9f33qF67CRWxvHEKQOtqHYg
Ofh+bOfahsxifKgyN6w+qU2peiB8OjZjZc7mbY0UA+L8PTJ3nXoinRtUOv/QlOXnuwqFCOrQ2tLO
S43NG/M2T9DeGgIsbL/6SwQuq+PxGKmey2pCrMQ4zZx3hzvqhoSUh8ILNSAZXPFH0u9wjFu8KglY
J+bJJ07cjdtnwsskEu0KrI38miHBpEN6qwNcdmNs6NEcjcA3Ubqvpzw0T6s8AukqE5WN7ac1bGri
fFoFYi0rOFKOqNGkepQx3pFl38mR2NRTfao0of7RjSeaJzs67+v5xwLldXviSZpH9EKylKiqh5Ow
ESnuUGO/lpRnj74oIGhKmSLj9rGiHyokfYOghtNwUbVAf608FsF/fOn0+ovBKBQY+Qa5s/15kps0
DzRSodVeyZfsaCRLDYzakHQqyhODAQ7scxjReoT4mMWz5zYNRkgThRpJqPv1WbIXmfhSxJV+ctNb
05ayb+IGHyaxp5FkKVqGwgfpZ4OkGLSZ1rRWHJWOzLJaC6E0iV/Y7j0NFhP1AGEzldAYBhxX1vZS
RaZHpDRdC5fmjcDLT3Jfkp/7/x8BMzxYjKQPRYxuIW2ZBQZ4lQcENeS5REb1dZUGB4oMnQIJJ+Hy
UXFw7oR0klNTodVBQ5XoZ+18A7ESBKBzZwYwJMhs641yFYnebhuSBQ00oT0VQ6RWS67s/IN+95Gk
z5vmzXkBqhLdn9LzmndUW09lLNjg1LN5mdnPYcu8tWJM6UoHczWEdEaBh3nSplONiRYQraMay4AK
634KpFQj7dmfkAo5qEVIhcdUWd5muKZUeojb38sgAWoBZYl+ZAmiF322Rs2kjpIaI9tyyqk95f0H
G0fRK3DQs47MxOhvQe1K/3Ziyo2OsT65DXrPlOmoICejeism2A4NJgHjdFfwfMbPYlnoQZngNw+p
5odE0b0/wgCHMjJ9UU6UNCPBMG3yGIsXZ/koR5xFgWl7YGjAgfmkZjEjdzAN5upjulFXzuYPsADs
QRlxyUHbe+YV1uVJRlEVIkUsaYcSj73YacxyEl6N0Rk6ap8JtWlY7oWZ2I47J+ZCV3LmCvz+qE2f
cwg62r9qmvWcclD9cFDP9O375o23Dr8bTrRx+u23BLQsO/cm1rUsb7iYRDrkXr1cC9rOH6qHpBVT
uMa/fMGnUAeUd+PHVRA5j+XTDBGNbtnaFBdG9y4b6/b5L/nedcChnF1JZsrBT7OSH8MK/rZ5JJGv
fyXpAWy+ubNse3yiKBFDnVliretEzXuskp8Q6HHExODeevz3ZKxMy6GQFO9QGvkXYJ0AzP6jzTpQ
VrP8Ph+Oko2YV2uDqZ0HTogiv6zF1m5E75X0Nh7w1pas6Si+26HoheguS3IqfwcWKq3HtAfq2dTA
yhrFXNcWsQ8WRFFbySLH3Ujtb3jfYqpEo0NU2Q8e840jvl4PPuGhXtHe8GYSAibZUHlqEcr4C0Ul
CxYp+kMNzkyCoaPug3NVvi1SViuk+T0SaoZFbXbysZ8eXXIDOMRi59+4L6f+1Damg9rbpJpNJlXZ
t+hpRpACHs0AkumMzVuB0i5wD9Nrsu+iHoKDLEpFbCkL5l5SaDNRuieu7hQ34omevYgEg83yvwS+
l0hCPnwRNTAWa/oUVyd+h5kQ0wmQqgeHNYcyGySpjhOyDMMevJIukvspxBY8HtOmHb7h9aQvIB+J
VPctQAeU6gt1Zmm+ht11kOP2DP6X4sLFqa9vp1SdBpuZUoSnBCmVMNT+Rp1zvvG1/9jEMT4ZlrlH
iYcgS6mK4hKIMwH5JdW9FUO7nGn00rUkVVC6bls//+JL7FpvUPTTboN0S88TOtcjrsDXrbKlLD0D
cwN2Tn5hyZriSNveT7pyn0iA7U0qzE1x+6r6Nvkcw1s3eEaIWSQ7bS5b6wqNvhPhtnbhBwTeDICw
/F+B0s8EbVU/D4vgIyJwJBn6VAvU5GhVFMxOQZqxxlTnDKjFuaQZXY1gL2se9IbAXUWnz6ZwOO3e
A/ddi8NXzsXANlbf1cg9XDm/3DPXaUoai0YMsL34Gy045vHJtPij4Wz0L1YwdGP4kKBy2WsieNOI
ZNgCPFg9KnyGsxA9knWnfaAROTd5Lzkv1L3YQ2VGTIxKfb+1M4S9I2wcYyR2A6zJxQh09ZEgLHkh
Ne6sB2iqBxi+gGQNnJ+0z+9KvkiFvof0EeL/Vp5xm6HczJ2OA3Wb/WW8xCgJwHLcS3OCAR4QYx6K
mKg7nY4t3wTl5F7Gaq4GfiQweMhfjGdnnwZ3hr6PLhp75YPaRaySYr3g66igCh7Mn8nbTID2hufu
TLBTspIraZp5OuIzVYQVV58RjdVKMCa/piqNRsGsO7IsyYGaOKBoR0cvdr9pQuOHOyFGQqzK97vb
vjr2IHuzwDYXR3k149eRUE4WwqKZMlo9Bpf/dTzwcexI4XEEnVNvU3XtGw45iFq82INRAV6D/To2
ElT04+VV0PkdHebOBbUbPBYftcyKCOi/ZF7GJGhf/4I/dkPhoHmwwNKleW0ZZQ/7tO90ThlZqoOq
DMjGaXPS5D7Nlg5YYYUaBCAKX0ZTTGKOHKhG7klrJgkNTmlsD2D5+7BCZiEfWcd1oKgm105GDMqW
DpFmanG7Ku8PW41aGclPu0NQ0vGPidrAxL5xrD8nwpuATjL4OdmK6lqRYGEx+n1EAxI0mF3kqSCu
BoqkYNsLTZnX9MTEviWWSa/m7HKl7WJOLBlDcVtBABf6BMNr+3yGICty60ES1qWn8+0ZMHmZQRn4
poNbOr3uvehCHQk0lFbsxsliQ6NxBYOQdNs08mpd8BPnXkZQa88YxENlTiya4EHwc2WOz9vpQO4S
pd5OGLMQODcWQyKfAq2E8XOHtvad3xHJaowyZpLrHkJ0UsfvPjSQKgyVeZc0g1+I03LRJ0RDSZ0O
4avunKRb9T20tE+xbz3xjX4Zee5Fe+6KQYNbm6i5QVhN8Z9ggbGIlx5GQvR+KIL5aGgZ+Dmn5RNL
ZMw3jD/GdIMnpyZqSMkVx8QBzWMYPeDJnvuihAKuSIv3abbKRPAWaOyhtc0hm4j+LtPyjVTIkhEl
wHEFigtLrUB70mriUW/HjU60Ozzu9wx+YJHDHLLzyP9R5M2uoiYi9kkTCCnbRA/F2R6Eo2hFk7uM
E76ir9cO6l4EsBNhA+2njY1pi0tYsIw/7Yy0xwaxrUqoAK9QXxOWwRSxTQVKksKZdANtbSFhAmcO
yKvfsbJM4paBp5jl85wSD4hn3IK4srC0J1LaVssKQPa97YOWtkf6n2+mRlHinyarhdF/gWtzinC1
f9CyseZeAC3U+uBPqKfJUejdCSM55CxZz5UM50md1sshpT4YQf005zBgkoC0Px6j9ev5EXOh3Jtd
cEpA6mHhlghsmxtdjbDjXd0EkhfPZh4cu2Seiyhg+Ah7w+pCa+p6Zr02d6XinD0sFduJOXHXS8Hb
UfBltiwnXqIW3YgU+TsWPF/sIczTdFWka1wijCYci1KLPmRxtx3ujMX296X9xr78bTtNmATSiMGr
LmyfeFyoOfnFvVClaAWLy8xlAIG2cm0RonR/+xY+PmQAa0oV4cbXN1Xa+ceKvhtk13T9Ny5gDzQx
2xbPhYJ3xXV6BYQmpo/7E3mUDigtdhslNfUQ9Y4vNf2xFHCXCfniU6xqKakiW57VCwGHO/t9eWg1
+x6eOstswTN8qhhQjLZnjIVSK0bdoNrjun4zvVPPX3jaeSFK9owKu13kAzwgFUPI2eR//DU09h/F
DFq51geR+258M40OiWn5zCwkPhztzFrPYO5pygd+KX+OYDtunrbPgykpAdeFa6DFb7ZYWIYa8nTe
NyP3p+oC1wyyHMcLOGkdp5LA0m8VYJLMl7nIJ85bh9d0dVGyVcDbvWBKKXbQdaRBVojt0h+/xtia
iQCLlu8I/mTuN30EsIjXKqMi4KNzThMe9fIuZcX5PiPC9c5B5ikA6UbvbA41AaE8bbOQzLEqNrnQ
7jTPzERx3QTqAQkogI394XpNrynOok4XTQpeBC8Q3xAKZ8XzO5vhU4ulHVcXI3jZO9RG1FFLVQ3w
HJhF6WhH1zrrZjTt99tgs9L45u1lr6IGYyz3ivarDrJ7q6/xAAkOhPG0szzolcrUDQj4j+7TPaUx
PzDhD+oeusNsppiXxGxn9ZAgcVREJfWfALmIUcMnNO7bDlO3oRSQWzYJpuDOG2o2ZmzWBD0LFiWd
kjdGLawdi7HxCM5x161+1A50k3yhrQD/4l2jrq/9sAWoZfbxnEXFB8TRfEu7OpZfcnAcLfLYoyuQ
mN0gtFYFOPWPXeYX9T48deR4Y9/cQFS7/nzzQIDi07uBqW5dU4p3KExvCbXoALtxUp7OWWS43Xa/
0nqIhz0ItcgVCTDnJ6zHj/xhNoRcgtm8kpeCuJl/CRqEUErlA4PY/+71vlhkoi0JwP5Ao8lG4pUc
Ybu4DvSyZJRsyoCpv+q2TR41qZ0HmY+XO5hOTXTXS70tkoF7ZNiMgKq+HBVqciiWcLJeGNFDo7SZ
tlHnLTYraolBxyUoa5uQ8Ttc0mN/zMt+nObiD2Kt++7sb/pDi+BJ2MfOj6jPWE2CbDi7675grjqy
8Qr6zHeW0J+1efTvvsXpM/TnIvmb2DrId9t0MLGg9l8X5YnCbdhDe5kvXPsv+QUzkLBk1YdYl8iV
cz++5M68L3b9Yuabzgl302t5wgbHYsdyIemRhC8LUpO8yxxjBENAHlbWJwa5wp/xntKLvoUoAtbg
GBegjI/pX8pcko5HxU4/xvz2mpqlUIO05r//FqDfaGnzvfyTGnwLJpnQsIz4nMJ7NOF8OIHgge7v
jSTvL41jeOGKPPk8OKJW7U8vZ9cZgr0HNxtiIDPz0aKCNVMrKfjuWl4KODNIduIbR9d8HF5XcYmO
wNxgJ3qwzHJNvIK1PtaY2K6u7RvGWlc6WofI0zDWRG0xEO8Do3RV7fs4VLTfH5J4gPTacBXTrwoz
oqtrMpTnZHSTeMOvV2DFB59kNeWb6w1cGltV//WnY9OcbOzGqI+mf3ijvhmkyJzOOJ+CLwQwp+8Y
8uiPjTYObKU1YNVR0La1HeQkDWt0XUdyV2jlhqIh7tAYThp1gxys6uKWUGPPHIk/zDQmQ1z67om4
k5xie4rETRt3EEb2hzPiU74m4M4HTXTSEyVIRQcG3Eo8VZEmgR3tqEJK+Zynw4VI+zo2GhRIUWUH
W4p7xlo+S48uIs8WdQ1byryjE57yj8iwb8qRusCpcJ6jn/JlD1UuBdjP0anU60QlcVe4Azb0bu6p
4Tv75wisHSeetmGAEx2vfXiuGCUj8tW7R1SgNlt02kRSI4dKaR8rlOTTtML0RHwLLrsTIKS37OT7
i46urkB16DQu1wzc1gDz0yL0oM6Xb8iZiIOVEGP7dI/f4jrc9C58nLNss4mKHHHWa7UZ25Q+YM86
3V8zDBFQeftXcL+WODhtBlKviaqSfULHptcSxxY18bej55EhWQ6M/3KLRtWFG1oVyLzRDboO705x
ScyB4qGw9scGNB6N36/zKQ0/YHBea50OCOleEV5ITUN1A5G/li/Glp6fvNvRx0ovrOWqvjXfRZ+Q
BuxYmVwr5LW5FreiY8IW0RXRmS9Q0fvyjS4lGnVYV3u39IqYp+PAXUoZHXbiAsz7jwnvgolfC/dn
E7lBYaY6LqivC8xdAYELFBSg7gZwjGF3S7BSRdOVXHOuSz/sUrXeImhQrOe3jr23725aPo6enLsz
YGHvAs6WHrf+QwXFW5fWiWdjlsQGqyFLzX7ZrmgwZhcEo+GPWHVOtcPTUhQpmtmQ6Xq5ZFK/JrZT
ChLNg9HeA216KRuPC6jMXmBqK332b3QT/HQooc9+pH5ABG3k7yx9e8XtTro+ud9WdPIgydZOfhgK
OtxBQvcTYFoZrBmEYVBHempqdm4MSMMBWNc97xzAiTEKKrGUfRH9bFY2LmVc06Onj+diNM22qk2y
CUqSkPjeZO8Pce2MnhzjsWNTnl8dgJMoS52S1tDWyVqq1vjFXymtf40OZS1HAQkwJPDV+WsgSEoq
G3uIrqJAmQI7VsbN4K9ugAVAVMPKmgloOP/3b2B6UOU0CcwuFeUF+aVVXU6gkbTeOfPa/nmk0//d
rfr3CtXTNSsfBCjTuUEJbBw0BlO3mMZvVgSrh71W1p4Yo2SCWdNhYusjP+XZjzEKqTcacGdeacqQ
dtiqQMiC7dyEc6rssZht2QBQUqoz+1DQvAM/jv+4p27Uig/1csCGwCzYMikUhBIszR0Ju3yEWelk
0Tzb6yR1VDXMXdQ70T4n/KND4XnY7G1m4tLwJoCLaBc8cr0DY4hS3ZU3QUpH7+IaT37JrvaHoM/B
ARD3h6X8QaEB7tsa+BQDul+1M3Jwyrr955bmW3ioGGqtWA6BiDc0AN7YN2xhfnov+2lib4KEAjiM
h4ysTna68KXGjOvCawLM22S+wsOSHDS/uEzEijwf2EEx1Rp+826NNfuwndmaGLI8k32My3V/K1+0
yukW2kYHoF1gN6ju7IXSl2u8QNDoLpeTwiBkb5hZ8f5kRjvNQTc06Y7FNyXtP+sWQgYnCF1XezBT
OsmsLzlQ5lGbrx+/prUZwHs16mCPjLhhFf1rte66SRQrj0mNei2cPZofnMrtxDQmgPCGV3TggD87
UYCrP5hSU5M2qqnXARJshpycQ3DK/gpiBUXVtb9HU3ut5izWaaikx5lHQJq9YYMz4kcwtPoAZRrO
toDOE/Bpibls4uWIXeibE0+O8yJbhARoPf2RsxcARcO7LTWD0qIFqkMzfTo/t7WCxPvCZ6Ny1FcO
mwj3J0sJwJYcspQSiIqUIlndVTM3alKp3jRhedUXn1YzEW5NG5K5DIyEhe/06dHf7BrdAqevOsL6
6stZ9oNWrptTzikyOBLhFbvV5FXk7g88/AcDspQek4GsZ7X8wogVJXM+LCc5NMK9xryufsUjSKa5
ScTVGinYiDzH7eKCTD76pdJqIIOoHJxPtydgyDvr5Qkbs0Ye5Iu4y4ka1WQaQ5ScxuxV+9BxDXoy
KdHLdSRBOiy+PHuHIdSK8g19qrBKG4duKHVlplsVgrQYm04CZ+boBDV1np7whiiNeRIMe1UOyyy4
2svIpiOdcUc7g5SJ+JE06Fx5ruYUf8Xyw5EH/tujwLOQKCwIVKdZAM6TFsYkbi33n5WAGuSpMllU
29LFjskwa5pYCtb6JOQCiILL/CH2aPHOfjaywYtsVlTOkNebMw79G4zPS1mJn1g9ZcQ73aqwUqKu
vk6EFipPqO/qG/7JZlLW/O+XObayPF1Aravm+nZN5i7m/FlLUuwLsg+NWEpd6mK30QZGcfRVVsV0
yFKDxU8xM7Oo19ycOzHDFigX//ztxCnSr05/3eZj5GRKW4nG9BCJEcBc3z/7UvKjNZXCzXWwwcgC
d6P6HSAR3TIL/QstBMgQrQGTHIMRwlYXbUonqkIlHSwcRstVV3JY1uPRFyeeedrkkAisyM7tz5Nc
bd9mxUwOVrlG2ZG0LVeo7+VtrN5g9xP+V+++Oe0i4wDArpDv7Qcc3J2KTpwVCQ9uA+y3Bv8boNfS
P6HoQ93+qyRqTDSxNAUth2YsQchvZEa7c8veQ9G6093QRz/ekLqG0e8RUndPuC3kCCFv9uUL5QxE
M2+jOYAziHLZqJjKmLSh00Ao+lTjsOUPlJqfE/OxhZUmPt/jdfN/AUJTKVU2v0jDae4SEAmhAWrK
ROvIo2AI42Vyz9ugnsJv1MFR46p8Q7q1YMBL8H+cg8KDxgyTvRTbzZyo4GWV6AHeNDBPf4GYPiel
2AN3a1JdeIwdUpshQd/A0N/an9b8ryUOxQv6M7hHXMxP7v9UIYy5XTQZOrr3bjl51IOSGhwmS8tE
Is+yTp7PnG/TrajJldW0aRBPmt/b/GYZA/+e7rTGyW3loHrs6B4xdi7iC6LJudmDFo9l1pKi7Ezo
pfCTDSvrQABfSVqD/ZhMMORigZ49PQZ4nLF8v+4f2Q7yfSClX3kF7U4PVtVnr7Qf3/xH5EHYHK+S
+mdWYV3VrfsHixONFd/X7YOKmJFJjuMqglTN/iTkYK2KjxTGrD881bYGXZEkfH7gZZBgZ3AcNJlm
GfPJYSEyCIiwOiOerFAB4yG1A7D8p+rV/Zd+w3cFSyaKRF/2xFo8qU3BxHzQvUYDcfYlQtqJmFhQ
kFbXuECGWeWnN+X+efyKG4UAPPihU1B6Lm9wCS8IkbTdjCeBUHk4TLQZ5vbWbU3WHA/x/TVQe2VK
VWa87ABvHPgBpUIW/sxRqBG9OcdOvQE1SA0KEcz8U1ycByuIh/OHUo5cEb7QpX1TsiKjrbj+JU5H
r471X4PT5+GXkDxWbutTNGSwdZGDAg2GFBnOnyj4wi9E6UO/no+3TCmTps8JsI2yk4KVTgXOG2ZK
XsNkkVd2Jz90sds5uepPWVaUp8R8lvwjqZCkt/G/Mw51wTTXeapfqfsel/gC465g69HJUeOI9dZR
MwIqBUkEO4Hp2nduKM1TDaOksIZxjMo3U1fPvDdU2OOFXSAs65VwNmiQcm2Q150gwy9fnPXFXAf3
tyMfrabIqWqvBTwFSvuGm+s122ATiJx0Hg/+J3bVjztM+8wDfhMKDwBRendSFlFtfF2SCxPJViOp
QrTDswegdtiLfshlDRJXLwhRi2AWUvlEheO5xCh+YUlJHfWGBLrUdBhvOrrvDGuTHI+2vEMpJYE2
vlueWs4gzFahKkCiwcTVmWlV6e5pqhXAsMMD+6Q47w+CjqaFa8O6FX7PryTPIwf7YxaWUzMBCK67
eavwTDz1msTQxrC5dcsvCKnAkvCMgpjSM+na+KsQ1MB+KW8hmSivXheUeaVM3sdknywq/NQGhSIM
ILDoIYkzQ9wc2Pa6Vl3w8xE9+KavAdLXfkPterRxEbGtpDVIxr69eMKScMrtny0eEIRFCGg9LWKe
A0fU4+W9+l/Cabgi50gR285xd3IDerrZsS1H9iqtUrJwhmFl1mk3h/V/eRbGczESk0M+PuXoizC7
hUi/sfrwb3PU5aWgShOdTd2oF4DZdz8MEReIbPo5QFCi1u/gitl6vrD/yZpSS4TmS6qJQOQ4O/d7
lX89P87+kCbDCosnVNPXVsMdQKv7tM3esKdAPgxDF2LncVtaDF7HK8Q30ko0fN/nUGg6TYvyx+P4
TNgSEDmvnZ3zUGEei9+4N5sOcDjq/iuSBzOFEHyQ+RMKZzz9FtQGLFBldk/MWo9aEAN4EnFi2q+I
LqeLKa12e9VoYiMualRkGV31QkdUdzQtpBKBQ/AOX1ipBhalnPyuvLlQKfeHoVLhxcUlqAE8ufym
DrCTZtycjNsFDoYrAeUtCqgSLbWLZKwz8Oz/q/85nbrzNmoO6LgULwhFx3yNWL+UJMRThFvTYyxo
Nje2w6/klWnEm/yHu0aQ13S7iwcfAD+xJMKvPSnfzhonLq17+N7U5EKrEdKvnCsJe36+NKWa0HWl
6k4daB+HnCzl4N61TcQCY8y+6SCcpfkVqyEreYs1ziFDuQznobrJ6iEqZOmUUvJQeBdLHCyj29Hj
SfVjYhtSAzHZkJHBs4WadTSkaJaswWov7LySKK0Q+l5399JLeAq0z9TxdS6Oj+Rc7x1ZkhUbWkW/
emMyBvdAy8jUX+4l9w16rbo9gYPFCV3C3VaFD0dnF56E9AabyITGUgQyla+Zzg/tAO3Eb1L2ztdz
F1jyLbOkVEd6grj3rWuDoKnNxfnMRDN8VtDSLTn4RhFDAzvVbHPlqd/EkmhyQ086AC0K3afNVFgC
Gnm7b7MLAnCJyZ1h02HnUuoQWj2+tl/mt17rA0jbiV9Wp2npWXWyzTmIu9iA7RilUpL0Dc/TSz4G
IAGozEJ5HykqK4KaCtp3Sl+uihSKeFi8Mh1eybSAw7QU+BErgDRzs67UebJZ8ciQxJ3lRI1oj+ef
Xrm26fjH/7O7Ptl+cQZ0MujRZRcrL83SC4gvVjSOBSgzmbMuvw27V5nyWBicElD7BCD3Oo0SNteN
W432UOSQVHrPxbVRu+lgmhV086c43HzsNH+UXy1NJwqr2oY5+WnfE8MwTxBhtyg5A3kY+99W0+gU
xO3zOp6P+IpCo1VjMqiN6BSi+SfSbS6xzlb9m3QQYietXArvG+DhBoDeSrNHSZticOgH99RP4Qo3
W7acNNBS18Wi+VXg+k8oaBI0PQ+xPOx8V38WqKl06/dEHecUUbrccS3do3aBqzmcRttA9rj6cvd8
hgjUtfo+CTAkNsJo9rzgbS5ja/l4Sh8T4dlsEgDkKYL+YqVITvYjxMAnlqZ0t8hOjV27wH6jTQZt
mlWRj0jl1Ju3OMNbxC1V5iwInJNDZ9DonlFTF3ca68qXa8A194v+jn2E0cmLiRXmWN64f/SfXVLY
lhjlAUHZ1o4AdXsmyxkg+YMgYd7r/hzqeMuzHmVCoBXrJ1KrcwKdqEcmLYxbLCAz9KZb2kVjouPy
Y+wKyaouErieHO8aJHCEUmMevLWNtbrFwF7avQSBLLSHc9wfQtedsZdK841LF38SPi31E5GExCXA
iEm1SVsbBYIq52IOopMomUmFyRdY0sQ/1BFdGbN/6icP05Nqw5aCttdjurLas6ONmL8EeojHdsbG
CtMiXwjkkTF9QjVG5Vx/5FmYkQ2DZoywi7LfpLHc2bb/V5UQOnFxUL7E03s4e9bO79mn9AbTrozR
YlNSqKDalDkRulgY0fwIrsQGBv6ZAUVineGpmTBlGUME66MvRCokK97e5qDvKBSPjQq7v0Bqw1yp
iuaxJU0CvbSel4EVVtcQ1B837kQlS6GuSQbMYNmxVn6grQk2lacgnskVgK6I3nlZNz39sBvGaQj5
s0/sDD7OIcI2CUd1aF4NugTjyS9lZMQUUF9qW1XlysXZx5Y5uSqnI63rKwinNTIhoojGbwG3BFl+
wBPzKwhbzE7/1fyjrNofNraYis73gGhyd/707Ck0j/wZH8fMyzHG6vebTcjRAwWjSOny9WcNxiru
Rk5RH9IQkMyVCOB/Jw+zeEsr39+Fp47b+LeHb77MM3dMO/qbatTTSroPi+4lw4Ey6xMjnQts274m
oJl/enNEuAONPMTrZqmrNT/Rb0FiaUUx9L0crnAlLw7aMT7KguiMCZUJb7AgvmDy+IGZXugbHO2o
QzkZ5BENhMshyipDRHCKhKE09BvE5hrHaAcI74+OSPgdLA/5jI/3AELZAFitYTnl7nxVTfIBR3YL
GdpdhBeEvQZXn0J87WXozO98si9O9t5c1RioJKfv1xwMzyb/xp1TRMsvh3N6bl6NfOgG46GiekCp
45w1kv1N/Gl4Wrba+6tfV7qbDQzWao5sIvbdAMEgIXO6KeH9R+l8LFgZMkUj/yi1RuphlLz2GBrb
g70cYIwzEzAgGcTXj0xCdCvMX8c141DyAgZ8Tjf8qRzHZgYv1AlwnxS7UTKCG/5v7aL8NtIUAF0y
4UMLGv2CRtpYB/yDPIhVErjJGNf18EvbRuHnGQdmgj+U+euVjMYOC0qT9zcTRySwW/UeBEbereUp
/wYHammm6jmbQwyJu843ITx4mEw2jUujYVrxd/wsLOUYyT0R+p7r9hJWFwyVf4IR4T8TPOfu37J6
i9i+jMJvtgC3tIGWyd02mv77kILSyTAqSQECWXBW927EO6Dme76Hifkwckx9JZHq22qs/6IGMVEV
f5nQ+/Q1zw7JuM3z/SJmjRDnB2DjisujtXQSki1RxZJBMMZh+z5XhXKcwmT2CwxxxkTbofX84yH6
ph1dZITNBrK+RUbhSYHmkLs8wQcVNR/HkITRGUUCOra3DxSHJAblHKemyOnbU97tsnsIXZJwnh2d
SttOSCzVTxboBTlx2+e/OiiPowaIONGJF7Jwfra9hNC82BWPiND+JTOVmpwLA4MQrVAB3MH8M6Xr
V5cH2YNemSzFDiBYEnoDrrm8UOM8CwwT5jpWApSGSVIY8+WDGmJBrcoC0BX7c7ntDYsBr9Q+41QH
odW4KUiBsAKpmCRnjc5EyJVI8WoL3ktpIsDdcnHNSjhEntZ4j2xoZYF51Gkd21DJPQiJr9NbleAf
nqx6MVuU2fXiJIbbKglHRD5UTfIkMcCdKUs35jadopkb6/sW+cT7P4HS3DVA0J2C4NYgpW/YWC0s
IxjVRWAWGGrQ7JJrfd3kmqAmr/IdypEkGj4oIPC+7f183VTMEh2MZdjqwTfOOsW4laFT0MIjV1GR
vhEn06WV/ChR4krH9E9OKYt0J9pL3w/rHStOcjms0ihM8x3xv6NPdAGN4F7+kT1iUNm2XWnCymyj
tZSfoQpvor9bW3qmJpaVa/mt9ArnmoSkqB5WDtIVce0oArwAKMQA8pmrT/pOni64BInxIM+tjpgE
hrMYFIOLMQqVlZbfI4u3gEVUd1h0lOeX0lFZmnAYULThSrTHxikATeXMO4Cj8IVWNknwFY69SQ4N
x7YKW2Wr2bv2t7XgcIL3YephAGizcf4TwvjcUfzTkytQfERxGgBHqinPHFBwvwx9QW+ZKssdKczc
0JeBm3YtPGkTvN1fKRDaf7MZlVJN6Q/OvxsIL6nH2aYVtVZwHIz++F//Gu6a+hXwWnxRKFE7JVdI
TeawjbmCxwg2AkZZEAjMO+eELuoLdsGkXqNwACQUJwL8rEhqiGpu+j3hI+k5hPmB8dhdR8S24do/
B1yPlYj4ZVukpV0owv3GMcQLeTR9Ce8neTR8CjKgtXltTjBQqPgFvbkVPlJ1F6ebi+1YXgrp/HYC
6V5MEcsAKmbSlZTzS1cIVnqUzJZ/vMkUPMV9Qk7SoXo6K97H2SGsNwEvZpsHRT0QfSPYZwPVJlV9
zmGlRILUDXWVtATqTiGpRH5vQyKOUQRdt86FgP6w4OpGxRfhgmyu63rXB8gTZorPXy1J+3yay3A0
3r6aRSrOsRiXGBrUTkyJXBjzEPcMjqa5y22gaXMvIW9NMK1QAmKyFBdZEp2Am44k4kV3iJEuOqH8
kAWgO1pXgRYFk4fxETqdd1uK6Wp9m5mnbLsJMz89JT3nCPFlzIEvPa6mAiXU3pFeIySy3BCIWvt9
giKJz+qLLOobPcLKSU69or8+AJywXHW7/B9yN5t/NRoAwjgvOcIWFvbs0lt1n/TkXgo3n4ylU157
EtHUi7cGztNQ/wQOZKR6wPlh4YFVGBUEuZO8zFNBAqVcqn0FlUt4dLxvAEOSoKjXI3qmsKeMBQ5m
Hi7pLSfWboWI/Qks7VNCjuCUII6SAsCubNH8MJ250F0mojqtm4v9Rwa4xjePu3WK3xC6hduHtpoy
Gjy/i5Cdq9GcA9mrYNa1cj30lq9mLHXyqWXLZu6WgrmmaM6rLnWi1b6wAowbaR/5jESxxozhdGZo
3eOc15WkGhviLVwa7howJRQFp1/rgzDH/RrRVr1wsSA7Czaq3P/sonWlbDk1RGAHU9Z6LqP8a8EQ
iW5B6PyNGF6yhbsJE4buca4g8qW7beIeX2qMcmL8Zn+pLdL7G56EUtPFMEggbHhaYvORBUCd1wN0
dw7qD+N94IeJ8C1iR1Q09Trk1lXa9nZShCKIyZNTqsZ/IKxa3Ezs6AFhlr3lklNezQJMNNdMvLxG
R8g8V+uJWUD+vSPlR128i2mH3ICeKKZntHDtJDtjazz1Yn0FkW38/9ErtOh2P3YfeNqPktgAQlV8
4UkyFbFN1hoTOH2UB8N6so2MilemoHqtoqmVB1s5GpCONvYL3cgeqlAxxRwg2WV8ZDJ8AY4Dyn66
QCD3EEMgHa5jyMaGJ5fgcwTW2APcsCvQ97KNqIaw4gQ8oOiSB+3nuvmTg83hjD2Qd0tOjSjnOqX/
pfxW2qloSqyMNag0n2BfQzgMluZd7UJDWubqpuRMraso7o4cb5gAeKyy+16RWKOjTgONDUWEEQdd
a7ka2fv3fg3o0Gd1virKpDlqj8IHXfofkbdymD0nYUe8N9FuLlPnaAZqaGQcOm2McxT2UR30+saB
Nb4oOcgkm/r4QTBfoiZuXBkaUXlLAZ2ijFz8eBI6Bc2LGZulvWFECECyTYh1z08+AgLhJ13d2A/q
AZIhNJdwkvjwjEoOowQxaFGu4NXjm2+8g//PTPze+jajSnSE8ZvsjA0J2UKJi8I9eYVv4p9DpXlT
x4XNPqjOmoZl8C+4DHoWNlDTK2Pv/nnpARgbdshCkGyKnBIMde0DNu9RQwbzkNVFVqeo/enZMkoE
hmj6yGARQltzYlvzTq/puLHYhXImYC90mtQmr6ol3miadRvPPq4Dsjk42x1TFB4PCwTQpfz1eB+0
lz14ZpsHEbV4fIGHMF7fXVa3wrMOOwefzNjH4Yy2HI6oUKzaD3lH8xwqiajFcaLEc4/h/T2GJLAW
ly1yJQIZ8pn1HbbMRAM5eEjwdUbX6Vm6VojEWOxbVycuVwZiWxGR7nJpa2izHVHffUpNuD7BBZkO
7o9/eLF7mhFiT+lnk4iybuHhqKgwtfDn1Y8KbhhC4rSJlzIuZk61BULx+xugAQHnRDMg3y46KDK9
+bg7XcBnSRi1hnUrXdE/DwehPSq0X+f+WyavMde96x2COWhOsb1C7iMFqsZdEyJSJr1OuF6SvP7u
H///BAponTbOparlxXCW1ehkfP0pNZWssOoSBS8dRPfpfCq6tjJ9AO0xvPzYcUVPlthQnpfzjC+s
88cqGraVZFnf2AMfmu8XvePXWm9bTq8s8pSGvxDZ4jbhrKDvoKfTKFt045jnuwLHboG2RuJiCLaH
BTIM3fW7SigQSuG58FCYTf2xgaioUYHRuJaUfjx9cWwTMABBS4jccrdrZMLas5NKLPR+H3lBcQD2
06HNcXSK+N/OFE+Eg7QYYm4QFd/hAfo+Vhe6RjOIZlXz4q/MKFqqA1ZthYNv2wTUnUF22o/bziYs
89oNPBAZGrwt50aQfn3aTUmD1nXmaigC/krWc3N9jwsoz6p8vA/wSyBF/jV9c52A6kkMYscypuL/
TWL47k20XOCoiMf1ZuOKLcDID1PJgibyASlxaexpBWVaHooNcat8LNQUTGjU4Uox39EKN5Clved0
3jcELBtkSPaOdE9m740MB9pwEChnmcFwCTTlA72RNc6EvFTRYLoChi76Dd8hyf7/2ru79z6zET6b
hvVAM4SPEVyiyjBmzkNGe6cpW6Nsrf61S4CFF/EVpb5W1Xm4pHXJSlvB2gJBNnVXf91GpbQRljh2
yQ/P6JXZwIvhHHFt6LeUaog5LPltHldvvnvMBowxUOeG/r+AP5MhWw2OugUSzJHU1pbe9z8ReKvE
Mo945qkg2zd7hDzumhsJlCp0trCDXCOeIDzrHgIcUrRsVUpVnCFR2rdcSkbE1x4f4xevGXu/sxxt
5RO21uou9QlyBpj4/wToBJdVdHhbwCLBZjvh8lD6fl3+UUXY7ncr/anjQasDPuhkzd6yEF9s6UEQ
bW/2sYb4N4DX+K829ct6MUf1rYpDRR2XIp+rkscAVlK6ArsdICZcv2gp/hjeZv4gWiYNtWJf9KMG
9F0/9BQY4LHWvRboctynj4c/IR/hXN95/S+Fk4AK85V5XCBh6EqPTdkqNccpAcO0A7pmVNGIKQIx
uM5Kix6LXIcDazJ+vex4brCucb9RX1sekfQdhRVJJx3bvb/QV9sXMHY9D0LqZJUKx+f1BBeK8k2K
8JENRD1ll7+h/nIjBYG54Y7n7VQYKJ9EJyMtmynq9Fsa2TA/xDQWps7gUL6b0ZsvLlAF6Xl+Ou1t
JoNEpcGE9QoZLiLTx0VvxH/ZqvGl0oabAoGlg2wqdWwiYNLOGOlH0ikmP4MTvGyzk105FlelCXYy
Be7yfY+6+E5fwErwW5nZ3ZanvEPIAafUwzUrSP8kP+Qv2bQbpxt23efXXPdo4IVgyUQMZiVUTuDZ
ap3HoXsRQij1qHgGd+WXcos+CT6nzm0G+x0P+v9abe7P1oh0gKjRkTl/41vqZpNUzQ0WMaVlhg3y
a8jdXvdiT0QIi7lrtNBpqXs3ki48mFXJjq9Ob/CS3neKUzS5x4+PnVO/fZyrTSvcTDpAKtDKS894
eKYFyztlRSsvZjNxDNOAEjRVz3yJbI49v56XZIiAL+zMZbX8Bl0BTO9ML0IoJOChJyWnLcBgxNV4
534JdiNt0yZAQkjXuWpPm6kGXlq8SsWao40EbjmOWMn4p5i/qgBYWY2l5VfxMc9r29vJaRppMYRW
stplzQ7VRNVNrfLAve4XTFmEzHNnOZcBstigT7YSzTAnyabFgRhY/uKGN7rS4tPpAGVKqFA5+6ku
cc9ZFJfAwnzz2psLtoxmYklsrZ5gnwA6EW5g1/8cOzXaSCcx2k+wa7At6CNBhsLtFnELsXY/Tx+w
EvqbZed2YnlDuD/GFQGmoStcnNW2qnzUNd6OCnfCnSerBLwiVYR7S8iYbI6cCuu/cH+b+dRSY5eK
kFesYUHx2foMto1I+fjQ4tVHCmETrFn26m0n1Zca8gzn6sDiIBLMDUNSYS+pq2llFyk7RSB8pUbJ
J6dJ59MQI8IJeCBncdVS9qATTqz2ZT+swgj6h7wTuGdcPka8KQVnaRoUBB7Ey/Y2rG1BmjGsfzAu
QS4MfxHWS0kkqBuC5NcY6xc6HKWeV3/sOTVXGV/fTCdPfH7S/7J4/W74ioRALQWvA4vc/HpV8Goz
ELiEMjQ2+NVO7r0hHExbueAVekc0WY2fi1OYPYtTdvjW3/+7BQZ5SOqRSSmjFIbG5S8UCfo60EtN
X7CvpIzWs3Di1/k984DansJqTDiG3VSoFgZU15hbtAgZKkZQcnkr/5Yfn24jiM1BycYCgwexrApj
WIPwoFr7RJhj2Xd23hrHrMSz3Paflwy3F4MNZALm0SZzeqmaOrjPGECudArk4zU6iyr2X/X/ejnE
nhhCWTqMu66L9uJU65j9MgZHkSYOtfG66/YkRJa+08jF5eR3yQEhiXQQWrBq2P2rwyY3wLxCDbrS
ziclhE9DRXQk3f5IBUrXn8/Hd78BErbDkpUv4+eB+ldZUKnwpW3GEC+35ox6DkbEig6dLhat6CR5
9d8c2n0ICGa8XX+J3+qHM7WVNnFQR7Hp/I5dbe31yT4EDXn8J+c0w4y7Eewr7sQh9rAvXAkif5VR
+4UIPxn8fu0ziHkjEurVWJnJ9KWhbQ5uTRipEqswdhhmqNo4vr/PDNWuhHsRiO/+fpRpxx7tHzfe
Hrx3A8U34DrniUxFFqGj8R3TtRni9f7FyZKx7lPcuVtrRBrKi4HS9bJdoDQSNATIhH3apRxRLxtQ
DPC/+6TozbOwlelLvXevwrYiTF6MMUN/6wYjxIKYdKF6SScY4NvSjmwpZFwyZ3fEiBoSaE6VJXBt
3YfkJILOXkPzYd3nYz/G2GEx7CEc+u7p/K/w4U0w41zonTa8B2sIV6ENnkCnINQUEiNcPLj0j7aj
noWgHfw5lqo776wJawCcGCuUinsV9e5EAG9UEj8pNHfEDAwKCnv0A73IO8IyBjpXZNaqzCe7t84Y
w7uXT4qKPk93hzoKyYXp59PwADuYI+l95DxD//OxuHzRulbkEsliV0JgGAM6mTtn9oK+G+VHAAji
9FF0veHcGE+iSO4pWYmb8nk7Av26Lts8u6YJftosWBrsOxoVy3bRWFIrfQrAhCpxEEL6ol4nNbw9
nROGcgvZvr/jD6sFBAWNP8ifiTC2oHsIRl/xTU2UbwEm5AiBMq903HTiPR+/+zhmHtnTMb0OA4oA
RzuFbXMxUHpoKXR3hw6osGN7VljkjDYSO48bHpq8cj8eSBXg4BjlSEawvozXTbjLMA1PcK1xRfk4
y0CroKLUeIJIS5J+lZFycpR/fmVvy7LtoL8aM9WojeJGiTuOhraO3V1Ow431ieFWvt6H179TIW2p
0gUeTTyUkwZDC9BlNPn5OVl81o9WAGtS/K22MOmvFHy333Rop9BeSvjGddgfmMpnnwQmNiL0HN6Q
ZAS6Bfu9Lvd8YWa3fW+NKDwDUTnwtYFAcNqWjIhEQNFWZmPMeevf0A7eHHxV0LMsWVWYYzqCNi47
QeCLW2vnvalb822zpRT9go5GfCaHjJctew4T1Fd2yyxJXVicoeEwHezjYD+O5FpcoSrhOiwj8jj5
Tf8o0n4msmTKwmYY4GNAWYX/Lom5BHx6Kb8aCIq+lwLNuuXgO9l/YJMjNI9thrFBW6BxXtqwYQA9
ov7c+VuxNTlAyT0TN8WoTn/VXFAj6yBrRkcxOgKLZMs0uAuGeziiUzTgGeGVoZsEiYfHd8cCjjNb
X7tYs6oo9KRkz3HHiEWucbNRQNJdTYSFaG6hwYl4diDNvJvezwDGclRyMk60iK/PCm83f/dkxQbT
W4jQNFwOA6VZ624QGQFe1nEETl4e6cjd+m8tyBB2Au3JyQrCG1yCgF1ZDVB8Qxou5xVBqi8a629k
3Nv7Ue6TOV/tu9AOIOh3HndTUE51b9lPX9NOg8GhgLafXN+366bKwCFP/x3tvNsmsKO5N91/fE97
V365B2cSXKtBh/BlgiR8sahRkFtgDDyGeaooQECu8K+aVAe2ESZiqvS+0GcFqZ0hPfSQKmv09GL6
yaYdiJnV/0/TpDLGYnzsC8bY4TGO3KfJS2Dq1f+yYjMU3Il4lNL5Y2itMxUgBOT/5bpELJu+yHP3
F4o8bRvAL9XCZhtnw6D4SR64Ck9MJAg7aMnK0D9DPPKMDSy5lZaofaXjl0oMIPM1flmssRoH9rJS
Dg+hFYyWI9K9jPtCv98DRF8V59DmcyDidjAWf0LseA3I44CS+mIBgp4KAh/Zo8aoyfzvMal40WWi
WeQyOE3zVMCw/G/HB8XAhVsqsLZvu7t6n2PJROa9E+IV8nfalSvuiYkt9wvuVQ7j6Y2VlRmrbU9w
jATbHJG0AE9LYQIhUgMkyN3e71xSqp193yERNkOSgOS/rVYA4OPJ+E1sB3hMchE8hFlrWZxxv3R1
OqmtVtr4D1dZnEN3g9VDwSf/UCQORFVq7nWsMZZe3nd1lEu0zlhnhi777G+GUmuOtoQ+FNxgfsM1
5/H+4ptslpoXn+eep/Hjps/2r3vywkYkBGA4yMGkI6yKSthRFlOcNPsIT6K54wFaC7Ofm3Mu5TEk
m5bMhWsD6tflu/T1GI5wALGiA7oFP/b1R2+YCEi3RwAdWDf4AVd6OWKLlVP/bOD8k974azsAlHi2
UAshFNY1rAWSh3yDeTWw0MZN0AZEezwwiORqQ7YkyUPIF0WGeIYbC85tQJncfWRh41Zv1rcZfbia
yRsRzmRha3x+YULaRicaUNPcIPXfqAYkbxnQscerTvYOMpupsz17wfoqVcDCgXRKDRqzqKPWCptq
0A43J4K207Q+c3Op7KbOmVbB8GBAHM51GRz0Mi4GQfMlm127XnQlPMja5GNzqMnYx9n8gOl7X6Gl
nJDp1SnTutxhretvVt2YwxdjClA67jDanoqHd89zaGZLwzs9qFGc2C07JeT4HBSzwaOzqF+b8+8K
efTWTHYEHL50mwr5hFMlr1fBPnkPzQo1rGJvpVNPKLwK/vE5ctyKAA9ELt9z4RoYy2dUUc/3wxaf
dRKcQ1vciTEw73Augi7wpRX231QiuHamXWqmUxukb4vaAdAE9WgfO653k+wH9WG12meyfWdHoO4m
8ymRwe7TYm16GE6PKitsHK/wcAV2xvpdTKG0Hr8Saz+ST999i0PCh1z8FJYeh95yUZ9ukDk9MsI/
ufrwNsh3yPTPpbQw0nzrKrE2C4hayJ19A84ZXwPHbYyUEDgqboYk3w5oraLWAsh38Iu9TXUGWEL2
I1wblqYmtH0w+Yy6nx9CgKq+Ldw2ZLEF8LgZjOftc8zgcfnwZufC4QevtYQsOtarHjhfkdCVN66L
V9sG9GG4orMzEkt7kB8Aq65QKERaXp8fIJ7Ui+xExJOdZOsjEGq6+oDfy9TdmRKEB/fBFenFUxMa
6K1XaYXlDPLlK8Pyraa5OnRHj/VW1ktRIZK3RFG/gsbDNq6r1029gWtIEJeIclv7efD6Fhe6XChr
Q1gfuRh8TcoknCd2Dd8Zx/DPUyUalsDvNyPrynYCDY/8Mv9DXkUNo/PftQMPviokjzB3qUlSRxWl
t8qM5UyZ83poLJHzIzGIDuHxDmwykw+UuFwvwEwkwoG0AzBPWHUnXg2cqqw8EvuJW5YFLLsVQ747
uMUKlDn4+1UgrizlsX8EmK6c/IeLLqtjZm+EVQn7pDPBCrRVTcJrXKmrnWqlukWkNW38FxmIwQ1w
iZOX5e26GL1YGxtHvzF4MwRJSWszxRUSTenXH16UdJI3Sk+jcgKCT7hEyFP5CKOp3ZHz6526hzh5
tNvpQ2MkTaFsFkIyDSUUAQ8fY1AYJUCYR6nWiqXkHfP+tmsg0BpIPSWSj5uZFav3iRxkyM3iD9Ow
R9pPlWNTe9CsZkZgs9xoOFAo6TWZj4fa7Y0dpHSaLqJWR3KJP+YJa2TAeo+/lINrurUQZ35DGGYL
koIM2//65564OXxxl9egRa4wzwD5PPDJp4N0u3cy8E8hzcGDHzoSyayUu7yHRBRKianJSeqGDak+
JO10Y8W/F8yXnUFM5U0PIfADksIGm7UHQj51VBoH2M6hD28qGi6luV1K2qynfTmj8g0nwixg4zuW
Xm2JyEySlNYMNbT/Km+ld+3sbBh5ytTmwjknqyBxCpIsNch6r++tQ84DxNFBNJys5/PeWdUKroik
5N50aGoEsqoQGnjnZrRC3SkYeA+votAB336IFVJt7zkbyXxXm+OQYzIzXhWops8i9bnOjbjAYfu4
NzMl/CI1JrCGkp07+yWSShDZOy12sFasq7RT+uS2zykFXvIcrPnMUyGxcYrCqTG2zwIALjjt/4TF
PYiaxdvlny3+G2LVLmN9LKe5zP1720HCKvwvnZNFDqRd9saR/LqRv1eHuspb+aElw0thZ3O1ScgX
QzlcmtVwGm0+PqIdNlBAYqSPhrFjU/oqvnK5YU7F9bEFCavqpybQoRJDeVZ4HiUlbMCTg5ABxktI
R6DXukxOhm4YFJuQRx694RiZ3W0tbyx76T/WU5hBzdEHBGlCJ++gNp/r/roR+fNkWJyHMkyL3SdX
lRtL1E0uu8Bi6UjHCdOh+To3LODnIQBVFpkqEciR/2XDwwXY7848CaaTuPzkdHoZp/p2mImVip46
xrNkjTkkpVdnXQJz2ckXzb+1FPSCNVHAlPZGinH2gq0qyMIBfNorK/8YZdgaE1leQ8cj/gf/oaaH
zieRJXBHFe9HpE6TuaPlOWICqMP/5dZtD/ZwK5WNFx8WC64s9RVlhjSmSz0aPYDBElXzVqe+/8YO
ZPKceT7kpFIuGv62oYRyi2CWxt8l2pP43bYWkbdiRrGUU02pg8siq/SJhvDbeQGLG35sJwTSzsjX
zUFB7OHw5xIa7eG6kNywLZcseTf2KcpAzvZUSORDq8csuKvinbb+p0Qmp07GF98e2J8WjvVhYIyu
4djpJ0UEuxeeh/EmpqYfcU0q7wXx4HQh7ADGldGzBAjfjSL9aoM2l84LXALye6VCHBsZaxYH8BPn
e3m3qGrJYxlLfbifQARa7gVly7fM6ERXd3kgzEkroXPJPInWHNzcMjNfAc2EJ+OMRh0NLybMxCrP
GoH4e0uXPxx2rib5DQpCneh3NHk/yqem/t3O9QUbVxkPmZuOh93gBAtRx//DppFSnOEYLXwJoESA
m4ri7TH0OyAzmlNjcoNq52Ri4Ut1kv6EjmuqVtKhvtGLQdK16hkMVNIymVJoJYdWHawoJgAL/xOv
Vrvaz0rSY7H1zenBQZ7E/kCASjtWt52JYMm2ypMVViHJY9k7pzcYBN5uRgfbT1DffndbMkiIrMUl
EH8zY28K24gzNTb/FevNjuFRRf5iMdqX0w8TFk59UQeeUpV1APUqN2hdVPijDc+7GqtQiPSp6QPl
lsDOc37ZW95MfDyrxH1JZh3HeLmo5nRgtlPCbVX6Mdd6mqyzcccLLKICybEi8dqJaFwMiiuciajW
DdnQsxMYRr1r87etda5g3Zr42eAe+X9G3oTvkU40Eta0KKHCbxIYGugHJb8OrdBpoB3a8Iz5wlwt
J9VWsi9G8D0aPDeTqc3lT47tZ8cNVv7x9CumfXefamm+kNuAoL3c2Rlm+1mDy97xktQ4WOg00/nT
Uw6ugDCCezvIVchugYENbMBN6xbHGavSihZR/OY67gT8si9ZzizQUaAKjrxg0ufq9fXFt3r6YZ0h
GcGRgi15T7KfHCEcfHGKmj0ZWQrhRmzqeGmL+hESJiErj8X9JylwN1md/u1BXBWlIxlCBYxZIWyK
g8kz2s9foMcftmGSgrHiNI+9IRL7RFwmNf8qZJRBDJYdPV87ew0XVBfvyio4xojTtgjmn0b19wc2
8i1Ubl2GLcRBEesAzwJRpUGQIZbRop1t1Emx7WO/gRhogpDgWzYKLJXAvOqcSacHUkCGxQTTjpnO
AbbsKiIkK9rRakoIX7xVpDulLpNALd5uP6sXTtaaEHc552TNGNFlYkaeWlnIIc//oLiizlUOdY6K
II668MEs4XR5UuI0qKBeCPY8gCbk7tbQqWxEB5Kcv2ZvKYV2waFQ3rwlzjTJCPlKB9jmf1tqLxOj
TDEKLTzT8jsTBaquWyLPLamzk07RrvH0/Ck7Jg7aQKShnbqAGshs6sjEQruhRMHGIZmHmcnLddKq
LtKdbejtLVBxMkRkU+UUsDzffsYhAxSJ0M9nUe8kgM945OOOzCG1oDwdz/eq9OfTrCBFwITaPFWT
Y3aTs8PsrYJHC3Y/vN4NyDDDbwr4XbfUZ2XH7x01p0z5Mo9U7w+cCWnieNVZJq4Q/MTm5GXfWblm
4cn6EdHTwHQdrEwckxsMAG/dW9LlhUtWOyyTHCO0R3AN89FDmHuQsThuFRYo/5P70vTqrTMKVh+t
YhH4P53ZkERGDA9ccIz1/JpsJETnCXCxUJog9FzJZnuw2gC5theoMkj2q8TRipMmgtTDYj+LcHtn
rddab9PGPl8BwLj0TYmJ9TTc5mWP1bod0KCIOhI6YfQx/UU+AlAPdnLMU4nowNFdgSsacs3+AFSc
CxtBEBxqjt4sWbzeAT84Z9tH7xklI2E+P6mFmQvxO2AshmdixTgXa8sXi8S01hZjnRGVgOaLoi00
JKgOTV7GWwKmm2YcAQq/5ZmycRK2OTDzdiIB5yMl301sOdzykyw8D8Tw45zOCfugBN4kR0sTVPZn
La+TwJJp9AhzsM2dm15bjHeaOrPEytkMdv1SEVa5W2hf90Pzagh+BH06YhXxs1a9nYOWlcr1dIBa
gcWwFMfenk9g8W8hGR4SgqiNiKEcnkKu3hjA79VBMCLcCWS1B55/n1zRfxg+sOntj/C7ciqjKM0X
RcKio8tqK+WfMtdy8d/uoT+g4JcGDRPuvF9jIho9+7bJW9pDJR9PwC4BUKvx/tIlRBgGhGXX0j81
Z3BlHK/+Rc52x6P4dt1S6unml8ajiT7YlpZ8Z/ArJKLBb8m9Q4qTOu7mSmno0fVVEkD9hf4LbgQ0
HQVvZEBN6kgIPfA4XUbnGKsaVb8H3cYueRhcssShZdJZ9hE+kalS9czfl1aq47I3fjeSuf/xNhGi
UKndRY3YporWIDbvTp0+IobgBH3RKhu3Ncfd+0KPTR4oopY5os6fZu9Uvb/cnG/wfEr+yEuX0FyI
0ZhCweqEP3zSKojuZ9pe7I/qwLWnKSpR40F21aqQCifaGbDvt00DToanq0GTzLzrjjLESix5UMbx
JsIx+9IDMeHPp51awDu9oAm7sFRTIOZmCoHPoVqBEXdMcGNABmngr0+rWxGH1foj9k1bJ+/QX2Mh
sj42vFjM6QMy7Vbgh7qy4ZknvSre8tE7VN763f5ak2uKnSGocI8JtbFTTPnutXO4ZPmYi/JmHAgz
HcxACEE3GOgjPgW4gKSihac1H5fxcMLj6JjrgkWGGrYmLmp8UP3rF4KepcPH6EKK2h/vXz/uMovz
DhAfX+lJOwPlUQGs3VxTchWqPJYf5oj0udi0hAUKVYE7JEng1asfGD7oOpYNVVx+DlzVStfLEjzY
c+xyxIKRLSzshGXeY4D4X3i4QddY9w8n9LTGl+hPtzr+Tl9UJ8YucdsmIqodwc0KGs14RYJ84muV
nCvnpbdrd6lEt288DS1hT9nneJU2/bLOue8/Q7Dxkl+CLMC4JZrmWEoffhffZ3Hqp7XHoGjthe9H
XhGopvm8I9Cjv2Mi9Tu0m/FaxRNH72vzYKZth2PcUSV67j5Ads9aV2u4Q0A3ewJPrsOCMLZr8nrn
bFXU/iHYNIv0/OXf9aGz7uMX/9XRiOAJas34d7QxxZ2fdFA7Z7hGq/IMP0RiR+PGTcuR1mhD2mPx
jC5KrKXqlXgS+78W20cUDK+ZIw/XydQrN4cljQWJIFJIwcn0oadwda+XFEWJ6xp0jbsNf+kUKDgn
bhdcCO8B87fvVXahq287MaEhqmczSGMGNrd0QXVgo1UFjX/6SbPA+4+n80QtKGOzcEI6gTe8PoUy
iYXrksfVaVGCclcYkesPn8wn8mnssrXtKG5rBiR7bcBbH8GRzDCL0aN2eAR61Wkk+L9gJSN1EKyW
PdTlNXxto/Ud0irhVN+gOspGDEi9eIbevHlACljY/dy6k9nZ+Uxf+e5Gl2n1zJMTzAwooSBI6GWi
65abHqdOKtj1qN/bFXORbZ/3ldk5rnJ24kdXEBaMw5N7G4dMLCptps5sNpI9+Y3zIHw5dRNEXfPf
MNQVBwrmuiYSS1bcqDy02+ERtGUc4ic21UJk/J7I2AAs/M3OhGpKubZ1Hw/dNgKv/3Ki+fxUzxN7
x3u3qXDVDZX8DxbAfFGty5o3jTyPczMSxdnbNQlJ8UyLZHxjaDlW1K3Kry1VCA6eMP4g5cPOZUHv
XWnHaKfIr/1fQ3LApoVoWoj28K+Fm8/j6TELRgfdOkQ/n7playyS9rx8Is1MXxHOkPoTTeRfRu+Q
/DT1S2Y0Z0byPFsbDvujR3R3VLBKf/pD0XoKCHR1zFxOeY6Z+JQn0BFlHjB6MYs1tTGU7WP4dX2q
0hDT/ch50y/FHCyVqHqVZig5JaLeKwEdopIP5aXGxI3LfpdEB0vfZKvestv1cJazSw7B8aLOzOhE
eJHFCm+1yW5RgrzuwzvJJeFrgfVzL2rZr9Ruq672qv2T3YHRSORWWUelylX5gREoH9OgxhG0iV5e
ZMQbsVzbl5k1Uvmh9ToLQEjR2iEhe5wozV2syCBwGFcyWqbxXizF6d0WwYGGSSAzxPYYocaOcEai
CEn+oFIpicdI6AiDpurWGdFRSchMtq/9Z1OzB9MUMBO77d8JBMRRNFrbIdo6cXqVhB+PfvwtiQpx
mxaWovBxEVAdLW12x6SRwr2MwcZwVIKOKCU9eKH6EYwpU2RPkM8/FK0y7fH6ArpAV7pmefGw6nCY
t45LuHXVav9d3bIWdOhwFg9jCVq3XlKhhpo7uAtDXdpyDKFXypzanZmUSN5FIZPTpZmdPsTeTAEC
lOGUiwm9diZevRQshRymdvEsGew7Jvk091V69OABhzX3C6EDBcJVM5PxoeOs5hHX9v6WnYJ1Tg61
If1ei++rK1+HYl52kwidpi981O5k7wDPQIBJXY3T0npRrih6gBlsn7DlDv537tQTr2Lq/OZ9+lcb
CCNVwtTKuIGqP2WToq5GnrjEdwx0i19mFsbwhJHnFdFvPTiXnOJCDiIdPlToMHqPrLbXyPHL603p
qw0eGoMQmS5fvQlodiG2rmTxcGGhHp/mtT6ReNuEP5Vn0Q0bKj0RayKUdkUs4cnIaNfXoyT+j4rx
ryEvS0oX0/p2dQYOrwdokiAFZSHBT7n3mMDIJPQ3ewDMwV4YLkr7eAWZyT9mqJSCxl0l72LqxmOt
K6q8nfXUHyG+K/q986IpHVJEGXh0fYE0/OxXC5G3yQ3iuiYp+XlxtB5nujuLZQmrw5AElIaTIRrV
SiGLmHQoSFdnOYHkqYF/ODh1mfeOkUsDqY6IaxOGI00RKIRe4HZSNHqXtvsJ5e58+vszpbMiY+oG
mizLxJW9HzKiWxTkd41zJRyJBJNU/l4zF4wFaFt52V4NQijOlo1Kmf6Vok/ZQO4h2tE96LqZrmhb
Zf5CkTUoOSpXjkWOXeOFUkXnt6oVz6XzEcHPWqBL1+Rd8/DJSgvO+zpAiUMENhUfHCA47NaVpokR
y38V39M8GgY8ZyBU/RNP7cOAO29N29PvG27NP9JwnQUJG120MNDynWQkuzbCcoXhUqFd4RR+xy1H
7wg8eG2GCPfci52M/clVtM7nZrMXX2q1VOaPgR3ltSaVM8WLDiiqWIZZNgocQbaE4SnKKjzz3nL+
8UUQ8ja5+FDXMyCmz2d8P9eDj4woPUiZRJobLUcC+0UuCkPHEUokgWQaTs5ZXHAss9oqOhIRchF1
c+Z7LUqu9Hvlkc2hJMC6DSK7ZhZ6mDAu8JNq9GOzS0ftsoK3FIynua9xYjgh6SC/5PhQNoMgHwDV
w0Y2kcARZYfZ4bnO+xbn5gOGhTeIXRv5AabDScpEVkJ3VveHX3TZSGvNrDNqKOtTq21YayZI1OPX
8PE2O2lUpUCAXFNkj0XX4+JCKmZ99/z5arLqLKwFQDsRXzJVfU2FpzOS5Ksv/98NlGIkPZoiPh7v
AwdJN7wpbG00/qz73YDPbsriSPTlpivgqkhkIqxPLQM0E/Wngzy0qEBNMyk1Ok8Hj+aw2OkVxwqm
jBkpAezBVsby64sPo3E/Dc1E1yikT3vlF1n6tZMewJpqcfQZFQOWdgl+mOV5fDKoYxpkBbHAHk7u
mUoRPhzJ7LXFfz106f5eypFhp5Cqi4g5BpLzZvMJ/3KqFU3seznD4wFlHqOB61f6eDoc9K1TJrL5
sDaMd0Bx4UKdqz4HyjMCpw/PrgyUq5SvHyWXNDtDTFSUHFazjs2p0g/FROiihCJ+Ip9GvHuD4H23
dgjH2vLz5HEBSHB0C+R6jsBUkT1XWO1oOYUbXJpl5IPh6R5qNvXCXMFxo4RVClE/RnvVk5U+iKv5
sLDmSfHcXRfNYrmUs22dA2IfPR288s0gTi71ldmnKX8xMXxhxT96cfPsjqQ7UMKtjtVVFCIq9P6R
u9plWSAPoGRhQuyIn5P9LBN6Oak+Srh26Q3MzryX/HCKp61VdGOgI9HCwTGnseQPIBibzFHfcmEo
xaJXwOdL/JTEM1NgcWDc3IijI3v3OpgaIulIMzpmbjMRLqSeGBkCLSfO4iDE9vMe6Lqnn8rSRG+f
UO1LkDEomE5clHjINLnWGtCSUYBZSY+iWn0F73VKedGO8IhSX5ZNXmwmal2HVTuF66UqwgjRH29K
/j5rny7Wfli4iSop++kJ22SGv6/kfq+6vra8XPRqYQ4lhcbWnhwSXSaSpVlmgoWYRbb9Byn6Z7qf
7DypdtKHb6Yf3Elg3wE+ChZDqQBUQRtucFdaDq3OYqcX+99GLrAEvvkzeEApAt12ogQEgc/Vr3sE
Ykkq3EqaAOQtOm1F/rY7ONaQcG4yNPPk/KoB6wkjo3lvOzLuhxdyoVmjmWBntObE+TJLvMGPuhOo
ix2ZRjaILvo4SXj8NPRNVOLQAiOzymOfJrbCvfaAqfGa7+RBGF7bTOXuXB5xc4lequU4AbVhyhPo
oHHIMHHpq9NGyYZkplXljUaPwqTJdzWtuIrAhVkIghjJNjby0jOORPchbraW68KSPw8w25UVrWnn
fyrB9JJFVTXiwzCkUtfudqq7JBb+SWTvuRgzE0Pw6xQE/fSnIUp8WBO5N74vGhZinXD29OTz+ZN3
fCAtGDK9VD2PrHXJxcISGaVPql2dB0aO1nE8aIZ+VVr7neV5amac81uBAl4FSgzEFpkiNLPzolDc
X3PzeeWGN0pvD6RMAA+t6evvwVOET0mFMCAfE6hA+NCK3hR//RarhzaHohhgsT9nXbE1F+NJLW8K
6Gn9c7hRDcBxBAF9wns92TzgNvljlEg8wmddKoHx9FbeMw8bUqLX+THnz/I6gsd2jI8PvZaZsuE1
MK2k18oeVr4ChcDNugzCKzOSSBRSDxmOZbkgl+lCxvMNf2TsOOmnmcJvr3SmFlS/24tOzkr9fCyb
zhOgAiji61/XdwqmZ+6N05JyyIQ85OdbCQNMmWrorKalJrqWbEogHg7ckfzmpBdVczdkRzvyXy5w
1wIwh+00JH88K348IfCM3BeCi/heOssbCyNKdj4Qc/W6KZMTmb2H9Cs9AwKYpL7sPZC9NKwjAE2b
6CzGtZUeJCnyKHLobvaF5ydAdjueIbMWms44R8UUQUcVbUo3KLhVSUMNkokUkdxpBqCcBZAIAY1W
cOUUp/vQuxE/zNPgT78+d/1zLubPPgudIm2SoJAGNsZuz8RvBiG2ZjPC7sMpvUiEFmeswfj0d//4
L9DEU91ZwTmnvQKSs5GpoLuwRFxgDnAI/fmLKuQ9xAQp1nTmrNzvxzNIGoxTxlfIuWVLAMAor1Se
+F3Fx4e7wi17YwpJzDo0zRXvSRI4qj4aw/IPpj3Nr7+v/aeBDomPaxZKgi0iMh2UuGxs6Lue6wad
MZxROlgWHnGjP00SVfT80/s/rwWOssTOJ5HdIRvssxxMQup24hMeockrXb/AZRb/al/6Ny5QOFw/
ltuc3IfcUNj9EKbf1HsYoolDsR4ttmzsPsXi4vmtNGu9QNdvJK1UhA74xCejp8htwm2G+5Ej4NQj
6/OJPrFqe1bVUWjr3jWzJvLcS1lpqp93cp2IOde0Htq5XZjfPfRX/6qydVIo17fRI7gBkw69ElHA
Lzd2UINNZBkToxXy2ZCzsHPS4xE1f8GwC9WxNLXMs5yj38N+8LOQmHrHd5iBrUC6doTQALRXMshQ
yFckT4+4RkPaHdNEDiN20e+27G3IlzvmYluboOsyXsNrn5hscDTi470RR18aPLt+H1wmjbh753g0
qFo5q5KKi+IV0+nOutxsASu//yCMa1rPj6bZmsQKQYu7G3mwdQrzGN9+Pk6pNvCmqKQVhCQzAPsl
UdANtQlRUIv3n/St5buTL123NiqZm62nRRyNjU1tIy/jay0mm4vQOhVi5kEEKiSSvlQpLw2JTfCl
50hUyNKswZwo/pUzAB/YgWT8cwwlSo4p5fn7qrV6wPS/9cEyeitpJ70STxKQYEyMe3Y2FWYqtJ1B
s+osOEoGzdCDSr9Td8p0tixZvwc7hyABWbTJ+B67Hj5kiYcdYvezYB8LDHqK+yc4P1d1PSh5eIHe
8g2Jsom7dX+BDZIXFEG/hw1Eg8qJGPbkH1fvizv07acFFm4hbfwWYaTvNfz5dA4B6JfqPno3fGLo
BCNz5w8u5t3BWy7K8T//Pf0PCFkggVNfeRBAYOLp9sGygLkUcig1z8cRL7K3C8nEL9qih3SeYSXm
uXhIobhWjZ7MTIbaPhaVcebwg6xeRNXkMG8Y8jZ2SEhCgvxpWM7gobOXukSX74VSbuJLcUo6rwEm
p+Mz7I/3RzM6SL7ngDpffsU7o522Ionq1TPVBxMXPzCK359TfAPwh+LHNMeHQ7WLnj9obOjZMvSi
Xr3I0CWXbv7jxrg17Zd402qWphpMchnU3PzTvJU7HlXYwYCacUtdi87ors9E6gEeEfqoVsh4ltRU
lCp+fOkrCzCKYUnxE9Sgh/IVKy+rZBvPDylqvPs2IhierLMXDE6NbjkwMcLkmUxZs1DSMyKFKBtN
jjO/Dm2ALr5VD1Dl6SCbOQsBT2FWaoEoh6IqOoceC+jUtuoEfhOGi1sZaetZwi14hRcaYA1xQHn9
sdFPfEXF17kne4edaoaANfVfDaFUZEWPTBYwz3x2SeSnem+CwljvvGVbAFP9uWiESA/20/6tsn1P
itL48JwTa7rM9RamIBPdvmVfGoguL+5psXv33XVkRQMvl14Wyt9HOkpQkzmindLfPvdZBp0xA2je
ja4XN316Y+NzQlSPki+1FmSwQsBgQIYGMU3PAjCYfccGOccLv0Ue0wvu5QOpJtyQ0S1p6XhnOD3B
1Qi9fQ2uFtVLJUgvlNeU6sCXkry1iWoLkfzdiIR1ixIctkms3gRRqIi09CpxK3SE+yMVWhJEvRg+
R2lreoMvIZFmRNY1iq6hqeCd41fOV1bxUJfCwjKU01drvARuRxHLaytYT3hNdE7dTWoGEF5r5xBF
mW0Ex6PPApaBpV0iqeyKllb7b7wARVVVZY1RZ+BQyNtO+SjY3DSXtOrGeYerx9a1GsCDf285Rnkf
9ynBQIC9O/yx8E53S06STa3/wuqddp/c06Toxl0DknKbUROqaZWu2VAeQSUnVKREKoQeecvBXxC/
mPhZgAID9bHEAvZbSPqBp61dGyk4oyKzzxzyw7sXJK6TyjHJ+Sbvq4NthyuKBk/kDIdPgCEYcvIl
tWqivbnrkx/RRdM2tHeZRSkCp7mwUJukUaE1Qixh8Bwjl5KASv+pbImVtPVeyywPTIHe7TR/zMmS
TT7L9zqpsbL8R/9iU8mPGsb3ltMKnT3fuTX+moTmr3gptvmvBrdN489BXNE3hk9ykZ5kbxmlTlBM
9Chqpren/m3y0O3E3MO1phCaMONMaJBkVguAziiOcbqHhtbFUWJoWeOZxEIgMbpNTv2j6kZcq98d
geB4D8nDPyz4GuxYrIJSPWNNz09dPIFvLLwBZJaiezBGC6m1i0TAUeT1duRnOoCstUBRFQw19aWX
r8KHUXlTC/vYDyoyDpyjhqAmtO8ZYtlqV32PaiyAFI8W7p92Xr3X1SKYyulsROq0ASaZXJnmRkka
D3qOkWZIXQI1Uui3kgzKmAFrBOQStxSZQjkMB91RSeQfAaVWK1FAsJ7cMSgmqK8HE4biLtsQbqDM
Knnrx6k9fN5Mmv8F0MZWGk5aSELNlJ+zs+uIVL7iq4YfNgJBy3ive41GtMB/Oxlpmb3TiDhcRwgJ
ohk1MQbaUCe/IpDkxwiA/NMEdAeXv8OpZIOFlNL8SAw5MapQ14fZ0ac7T7OA8YsGICweSXtuhxj5
OHCJGmmqLqOilMr+QIkXj3fTKZXfNNUCi5MYCz8ICgDEJ2beJgeOpyVcicZtdte3Bv92VW4b2ywU
nOR8+TSObrW3VAEyGEAj7Dq8QLqzs64AYlNGJw2pw+qOzYDHEsLTX0BJotLLBWM0nkfx0MPLOUyy
TCbWHRi/jCSP8oArXBXishR10abYdB8eou3tTR/4wu3pVaRMC0QzoKPms+1kCAmF14lu5PKP4djJ
7pReWktFjAmusPSz5IyIBmkri++DSwLTner9JwUBZ9twp+0vvtqHpuO6i6+2+eXVO42Zvqusyn3K
3git1asmYPAknRUXK+OGAi/VN5MTsgVxhtLBJjlWNFWB9mJgNYNY0Tu5P+wLbIbeTBpetufLqiUd
LQDnHP7eKEaI/akYB+A2oA7FMy0b/gY91I/MUTCYJo62zPbQbD1S3Dbaq/VLFLjgzMrNkmH6H6XI
v8fo5n9lRCFtQPuc0KM7+zQAKxJ2jsbifIIuK/cTTwpsZpXy42B03Sa9R6MDpFt1STiFRoz8LNYe
t16oIqKkz4xPtpEfAnNIdo9W6a1QDx7nMWOzay1qXk4lifWKmYkTje0u+v3HNhp67DDstovXl0MR
QY8rEdJuoxZw65W1e1D+VMNTATEIPoPelLLgE8swgJoaaIcws5kWKe3Xt9IggQXZsP+rdSk8GXjJ
cBvd5gFjlZeCBdqL7jlvuIBSx1sQV8jDtnGL1z5Pn3W70UUx+LG59RPIBl0lGFw7G9r46qVeVxUX
xMlHwtOx8e3oN813v7SfOzAxiZk8W/1gnuM5TZdkji3aP900kC99/Gm5HdVxxZXdTtBkMFv89gl6
dDC45SJkNj6Mcnx+N7a2ZNBdkpusSLp/5vyrNILMzS8ijc0mupfduxe4z3fKcULIoBLL/7GLc82Y
dynB6fk1TMYLNlDvZtFKwiutdpu/Egh14RwW559L1pMojvw2A7o8qrr6d0Hldn6gpXB6ctucYAlv
YorzAbKHKCdxip6JutJ00eMgRzG1p7LqOWSGvU4Qmoxch1kpTIQHvbByGmWpfF8nE+cT7ovKrlfT
5nRVW0DtL4/r4FD6JexkYCqo8cl4ZFeLfdlizUI9Qu6Pwd6tGKGDV822MWDVTqOJOjDTHWug4Jpr
YKS6TyQYnCJSxGqlyJFTbxZOZXci/v4vwcMYjlwgwhbZGeJbnkD4uCQ/elpbgLAL1AD2DlSlQaLt
Uns3/m3tcFOC7x3BpBVD3pKeZNCC8bqIRttDOwZVKW4kCFLSxIYjwMENqRIDiBmXfCcfougSXHvF
CF2K8vaoelNRbLO/5yllEPIaG07Iiv0K4JKteEZneHRfa44PNfk5Y3J0E4SVtEG3Tvx4OB1dLdJS
L+zRhOxNH0KLeUY4sCTKQdYWA5cCcNsq6aZ8RqfHU8umERcPEBtrXlFjUhk0jAiW+eWX04NM6qwV
Jb8DuUXmNydr5kGIL85Y2xtxNOW9F81w182MvKtbhtRi1kE+HcR+bK7osVINWPZMOk4H/hAS7A+W
Y3ZMZoIKBsnVt4y6B7O1aTst7yoN+uGnoJ8pv3X98L+83nZUcy9BE6AV/4/6P6tLIl7ipAicJvuB
rTP+5yJdGPt/kxqQXa3laqpEXHZkdYas0yKKXEYz0/yWQ3IiL/L0LVkJtbfSQMk4SZ5cuaFWqHww
bl6tvH53NYuGQerQ3oY2fOAxW6AbW5Ioe3atCAB4BNe5yGl6oAEWGO8SsEETENwz6a/VtnTDMJ6Z
jTP0pYtMFM87UGHRqZPBp77sXLf9pE+79uqcmaEr7NXYYb3ujF3H/rLJ4qwvsciKUn8FHET1IxID
insBK+RhJzaTBKeN6EFEjgBdUByi5foGh8qDXNHwVXK/BJjlF3EZyOsK4FKKYew3ICZQLjCqYr5K
YjSDa3TQCGV0H0suQ83ur7v7FtxrHOmjNkuqMTZNqmzKJ5yot3S5HwTFMy5AgyYoFwAr0unkcmMs
89GKnOed3ml1duzAK4/oyik0pi9QvTGot1xNH7BmKdR4nRYU/Vtn3xF5ZrTpfiOqSh4D0SNbLlsM
NB8pIksPs88Ihmdy8IkvAXE9P7TZm3vfF3WFXvyINlkqi3xNiY4HGJrkXDU2VF7vYlgjRp2x1MCl
+VB5FADhCKsLiiWKGmX8pdd2/vrK/yokCL+xcekcnvs6Jr62VHwv1TvFUMv1kfjZ6XHW0ppCgmzy
7GH5wY0Hp+XxCymeJGxg7D7zF9Yy3Xqpq5wLkPXfrsu1zIxezjsTfAEBRGUfV3xlMO5koHprSqTE
IEofpBUooyuvlUmNK5N17R7PjVf+zsPBUf9ONFBPyUpD6NXdQBvnbAvr4oOe6xPOIiNwBI6QeZpk
XVMd6ZkGLMOVAdQDYuA7i8sBoO5nMXjeoGQlCbbMu0XptXlN6m7o+FcnIkp7dWx26PxjZOrb7nPU
azIKsl3+MX5HNNX4GwWVSJS1wqZWy4GD6aBAeFBpRGYm/MpJG41DUtWpr8ErjFZ8K2X6bWxv0syD
/FjGr076w8Y839TAuX+9nzTy1n2OZVqJyme+NtaKUccdzF5CEDp82jik6dqYpeYXxvaiBS/yLPsQ
CbARz/mF9l+X21Fm61zHltwZTRNVC/QWCzM0DcQI6PD3kKeNGPrE4QebTUbnm3+iv9Nqq8n3ttJS
Anpv1Z7+j6ABtmCnz6A7cimeAgnJ33XCjFSEa3OoQrxqqf+duVPGG2j58qAbUfmd7Sv7TrNBEYFd
HxXdbnu+154UVjUhIxVJRadg0S/XDQpDatWrmtueJ4uFUVuHMtplCDQM/DFC+QVfB7eY5PphbWNO
wb35s3ScFBgkNrDHejhIZrDeUj6i0zOlEuEiDnKg61Ru5TXOG9T7bJN7oCzuGDtv8hQGtbFmnVYS
jPeH4RRt0S0Yzw10wQb9W+4X+Y+ely1TtoX75KQF+nTtFEvxLtiP8eugXbnOe1L+/o+eMpSZY5Ov
nPj91VDdMofDFU4azTuvIJ/GMu405H9w68VZB09K4klyjYAHZeuGLrpyLEYL8r7CIYIUJJtoxPR+
UiKBm8uR5u2v0AeDPQ8fAFB/6SdfmebMeyRL9FlrNDX/9zWWTYdoef/fde65N2jea6K6Q3LtOIUX
O3nBUbBhcUz0dIAmS/493frDZBmCMeK3pi4NmysUVR+T1g2Z9cGs/VYwrCSxalbU6t/9iDxoSYS+
JRooNB7jN4QummkQX5qiydQF9x3jCIwX9qyaFQDwCUuSS8gt/O/1JdyTW1bI2lOXC2bCkf7HS0d6
yB24uyhkwjB+imtfPEXauE2xbHe7Jbj9e5MYYy8bP7l6/q2Fdk6bfqta8xMJiPcNoqMpK0g/D35+
e1hdB+BRE6I7DDVU+jNs9EMkgD/s0DoLZyeRH0axNx7/bCJde/OqRc/3jaQfP0UrECachdnJpENS
QKXuovBhh4HkD4WwlzwdaYLVXzko59bvElZqsPGDUJmbKNAhi+k10nOm2jNrWVAPtRLI+4PTdTZo
sEudn73UsNSomVxCJaUB+KtdK/yfv+huXbsjaV49jRy1uPyIofHtXagnpnzV0vwAryybHPI3Llae
tu0G+6d4DHu6bVap+XBcVb+DOp3GufFMjiBRo1oH1grby8OtNuBLTIdFjrUb5Q19TbNcZ9CqqKXP
MZj/D1UkrttKpwj6hwkMVgGPq6b/RvN3n+YDGQEaZyklXWlP1tduZxF7/rw/t/CZpCOA6IB+MP9m
lVCcUD3Odvwla3F0crCVPlA5y4L6rbkbtkcL5NE64VMVAT8ZECAudikL9JBoJnOGhZVAbK28kT9l
2D60Ws9oDI16KNWQMji7LKJeKAYhQ++aL0g697ayHnhSJXYZGS9XpeHuvi0EvsdgH31fNXc8Vws9
t212GFLKsVsPQ7cwiqxNKsPderPPxeebMuWkBfHD4AJM3aTqE88LQk9+64a19JpsaWiZrRgSk6N+
Z82antiPpSCTv+8/w+ifvzmaIUGEdeKqgkJat33BBxi7ueVafAOZHAqLN7OnkS8dt7kY0jXvp67S
WqitDekp0RiKVImXtL+BVe4ziC9vs97yO7cpWCiXt375MHLBEEwBX058Iam97ht+4Cb6rClYttTg
8RlidaCnHq+wqtzYgMVKJiG7er3jNZJhRF4rZH1wWJljN2D8vUMocqIto4buB3E9fwae9Fw68WOp
jFT5XIoz9/0Bbfm+B7Y2OCTm9UgzDun4nAE2kqRCASpqUQObBwStSiumAuRiJA/6jFQU8jv2TIj3
ZPqKDH5nX5RFY7PrQleiAZ/J4cGPaCrJL7L5Yz7/fVY13gyRkNphrkupgEWRq6IbAdZWIGm7vngR
A84Wr1+uE3Wfe7+h2e4y8BWJ1H0ppGl2fbFMa13dmMrVO0LxeYjDO9heryrbgTq5diAagroLFRPT
id4IvoIDYDAMeeio/NSZ5xetTatAfBa4dhYm5zgLVSMwF6Vk5Zity9jehMW4wOXLTQOygHq9mHCz
ClbLUNGEjhNSniqglFaJ3Lc6crVt+GcVE/pxFx3XBAIgSC0qEAb5d/yIR+GmqCbrT5/Bw8RYQkXw
lcd4+vR7d1Iw5OrKS0mkWsmh5gBfvHO9kj7kRzu5vCMEFEkvUZ8XlBjzN69HlyQxBDdQw59eCgBr
cSCm5HscyNFQdicDxL6U7WnjC8QqynWv0wVb5bsrYJegcSoArqpQM7moR7UWVGoLtW0MlXR3Yrcn
H1J0ZrG9ZOOrjvjcNB1OOjFinULCTtwgYvmPcOkawRzkDD0NHKa656zwkksGgqwBI84USxwuB2VZ
Dng5Qrb8crnZlG7oDGN2f58YOqZbvIpa3FA7oP/vs1ogprrOtZdb2J8LCnlsIrpqfIH6pUDMGv+Z
j6UXLlcgbAN8YlTvDEMRWYOHLWKeaCpBSMLwH5AU+Qn21wvBZWBaAkhtBEvGw1jUAPki2A7D+QmC
u6FJ59YyvwBGRIcNud8IHXA2TpBWPP8HTUcKIEyjKmDfx52/bI4LOpCC9cAmEM0J67jGl34SA3rN
Ud9iOEzQJCOS5NNbeOu53PzKmcmMbG1zYZfhSumoMoRNfO/PvwKdrFr/B+PJHQhr+VrYlD7LxWRl
yM9KQuUol8xUCbhPxp5DzecTZCyDdJEaVuA74G6wBlg86kkKxYYgmnFXjGF/Q8ofqJCCXbuV3f0b
98z4tkYuPUeUdGy0hhlWk9i8qAcmmXCdRe3N+1Kt9IdBRDxn5U9/PFXaTJA12fzroQkGgwMuwOwn
8cbfKXb4IZc6NYR7vXQO/VWEhnf5JkfAK9FNNS0ggYBH6Eg+DvyU7UxqYmGutf2gfx62g8dZXpQ0
VyDjFuo3D0CnW08MkjXrVyUXNKUAGUWnmufRhnoxv9SXI/ZVNZUvkMZZVUxgEyjwH8WDWGqdwBUQ
UUuR/7XPoOlY2kLKqd70K9mHEi0UCQehBztYpUnHPOjUgfWXu+ypGaAtfLdE+E4aGiWv10gIqoDH
e4iJ/FreLTVF0Np8iLuMcVfBlk7nthxVS5zGMhdXd/j3uUOIlU7/OV3BZ6aJDyPhgvyKZ9H6WHJV
v6Q5tewZ65JRaHIumgMitxxEx0OAchnokbctAxsbPkkuiR2/gf6WVG0sLzgK8x4e/02oqqarZGSw
z58mAz6vQB62Qm8G9LVjLSB+IyEiYJfUnGcx2UWqBfVEGU8fMjUS862Wbel1uPueD5a2ZxCioewg
gX2ZslyCqEdmqsit6u+Fuw6vMIsdGgIdmiDMA5kCnfFiRbYw+QhzYj/kNokozcKwSt7FQRemGFZh
ByDjygbI6dV63g9MA8NBo8/edwuWDgGey8Fr4R1FzII2PnExlpIytTKjyOYXGeexLdNr78bQqCpy
qJbySC/8KhRFcCFzoT+4WSQ12wa2B1QD/5Tm9Tl4nXrASweATc+SxMz5mfIUZ6rfFDe26sMIFxvh
zXz5mZUVt1O3VvGHIECvLUoTfBN9Al5WUFPiiVmvnkMYYzJpCvEwp/I2e0B6Odhgku/6CYMZw6Jm
2qATUNjZGqEJ6Jh6ruzAEwbWeffwbvncmeRoT4vf7ihw0ppX6J1PGkxxIZTYgE6mV1JyOOh8DScL
LyJKN0BhExNutjaWerEAqQp/TmmRD8Tnnvq92rLV1ndY+LRKMlq22++zDTn+BAqFnYzA9A4zS/QN
BU8BJvG6NLbBMRIDhfQGhQ8ekL3Fi9mpoYb/raDRoi5/1OD4Pc3Ar+tXtIQNXO+2mfZIYhJ2vIWV
7i9La6MIgR2jl2m28FDqqjhqxs5pbhT9+e8In5/El6EUSdyrIP7oM5xYqHPu1v/z4fvkNytLPE+V
nCma3JdBkiso2drjNl0H7P1z1Q8cmlAiUSWX4x3SwxUGzbibHItihKJ5UT7hDIf/8wF9Ef/QvfD/
ZrONcHVVPsRoSbmJAu2532t9QjKxQxHIwC8V3n4zsNogXxhBoEoRKRDavI30EuEwTW2cK73/Zngf
prtKiP/QV0AdMcTR3ALbIlCvPkWTPMprARCfw/zCqURxne5N/gX9HrtLkKc660Iiv0MOjoutTmun
RFX4eYsFkcLm1lyM/1rfta60Ug9cdOtGaPkS7329ROJcwMgmK+X4srRhqHXGEUQhRE60iSE7cMCB
s4vX6ysgjH7HcHVNsy/ST8NLzXogd5zNPEzkfHxKYI33T5oXr/u03CFe1XFISTqdHQBsERSdjmx/
XgSaF2AMMDl5y8X5X5bfCdX5SUWVPLU3QzY/IYlJumYID88Thbk2JDPMyfBMFaHIF7jbv9Ljddrs
qJuoSQ1qlqaYMkLLV/jijgPw2vbQGHfQfuLaNEAN0uZ3yAPB8nsxuL5ld6ihgXGBAmoMUQ21NBjR
x7a+ycV1bj0M2xj/Euc+nRNxatumfBnrmg6DaSpFD9pqbagqKn4kbn18R5GDrxiEcBCsg2SIaZGJ
PN6pvXjoJXNuDU6Q1aRrS84IB8YP4Ig96XaewZiMiPoNK1khl3dXOYNDCdlillu/zc27DOVBUvYn
SCwIot3aDdYzIWM23Qh9CR38DHrEhORelE5YqVcP0w0/2xqV0MB5FMma+kVz/it0BuKXU+smfhru
+H0PjnX9kVmh++UGslRQs3NuD9KcPAVBNoKggJHgGkQ/mDt6OgBnURjsi6/IEu3JQdzuMv49rkzs
2CL6ZR4C5eQnaAU9zWB49p53Rrv2EDLViVdHgarVrvuc9uBNyyvjlwWImET5XUjv4563fzyvED3c
xMm2u8AKX3ryVVkUKiM5WaV/b5KNxRLYjcjVaIC0Y/B8pU8ncFASehC1i76az9q9m4dCykgB2Hdu
t2zeVqZOeeyFNS/Kb8pt0z/vRM2Gsp58/ZKv5CLoTnvelc9wP+aD7RI3j+ssVx9qfObavDV9H3Er
YplJXQStcY0HjUOvuZUQqqbWiVpfb4/205TGGFFVddV/q7G9KL9f3vWR8fdurLo/xWPpvRi5gr58
lDLRfk/MJJSVviN+uk+Xp2afmVfdVGK8vyQvudpF31/8r4wZ+OIzqXYhC6HpwX3p/nYEtVrZJEIS
DjHhLC9fWRSZMOJYs8TL4OLokRFPhuH6MTiAtufr1HsxEmCIWriL/OktLtJL5pFKG1qpfUjndsQy
yY4j3KYh8srDUE5LdQyOxcwHG0w7qMufo/RliU+/EA6jyVIJhq2BfEFyVDipSZN2tv4a5zTxp5N8
zkgn0jF8UwAkLsWDMPgBzmDG9sGF3o9FTIMTLqT+xm792IJ5rLwJ6GzwAK2j42FwED3LM/n4QFxA
lmWq7fuilwMyovnOBB4K1TjQ5gzUvhUWqUZl97Ix/zLF6UrJhB/XVKgzG+Sj8ZA9fAIB7cseRpfi
Ec2vuj8rwWs81CnrzPPXzrTazu+i7Dxp2Zq4SGNhxrBxioWqmBaYn6Ghi65oqo4i38wU1Tj5N9j0
QvX/6jpm8heDofoJ+SthSwascQGwMLGnA9sOpp+VFsF27Jek0Z7KJzfhLixWk2ZRdETCDgKVKa+U
lLTHyQkq55CcoYhtJQnKuMuzW7SamOcGbHQCI1rNidng1i8w+hmi6VbQbycfIdbWFKisFW706un8
Eo3kzg5FCqFeAxzP1JdIysz/Lh2lmAya5pDT1hBIxPsD5NzK2shLoOid7OmXWfQ84jtYPt2lyrN7
sBt5nnl7ds67rH+QbYp4iLxa64pioU+vl9TgQl5x/XXZTVT8bo1E0sH0E3UiVN8Zc3RAhQPlg60j
B2T0ANDOFH/1lQi5Q9RMc/5M+QzmRMmGDCKrxiysjdnYyn71hQdTezA/8No4peMevIBgiBbqpgBE
cy2TRp7yGbivDzbwrU2S2OLKvOULEAVxfYiW5E0jJO1H/X12pOqJ7Hp42ypqzTjh8N2Y8OM5B152
Br15ELViFTWPW5exQ7eWbx4+FBn67oFaftq0PL9BZ3DagnTZIgPXvElaedt/WkQR9bLVW2z6Ggt0
CMyJi5dw4ZFG8kAL9HGMsqweZIHGgujm+XmijCqtNpSr004MGCXnlnV5RR9DkhzKTuqIu2/GwqYH
cViRQoIPWLOO3Ny72De4Ve5a7yaTfRQYANIo8qcWutWUsvGlEIb1guOEQcDcI2N58N9qk9GNYnm2
OFwI6pvwwWIavHIgxYrfYB/lmpRyKfPkB33/vlsSZRiaeC1ote0PPqwNtcNOP4wdxlUSecz50VlS
+9tCmLKmoAr3lFJN4lOPyr1apy14obtg+ekT+flGSMgY3VVOQQAVCYO8ugfc+Pbku56T0fd1vepR
Azk1Cq4Ga3zXr7GvOZKigcSpOCtqWzBVuazmxabZ8FYs0BAorbvLKLi0Uv6H04s4EJiF32e7wnT3
3DSyC1rECCuXYo5Wc3W4V8ZF4dSbvf4T11NqyfXeeINBsc6wO2UeQ2cqI+OvIxJzwyodJqYTikxf
qp1h8Hgmr5pwjNk1bmVY2uEYePpQniLBPgZXJ8x8/jAqYzLMhARhVymJ5Zo9JNLtjB0WZUOALNTR
bR2atijumGdjsw6U6pcQb8zBt2Ym5QTP4Mv0uR9DeajaO4XjEQ3TA1IynHSFm2oPzQsYUnK51jA3
kFzVKXPxRWhc6SC6KdQPv0UsHfrGBLLBymCQnFMQCsbKGQRGGWxJ3vercPdUZh5tf8diOzhVUFnB
TM8BA7HnY68WDUQDzjUj5Hfefi10FujmaxXAek334VB0GEzUvhB1CAWYKgVbPgymZlYQBT7AOchm
au0ndfSRHzLE5x50F2lxBzoc2899JyccR+K6RO4iRFNzRnP5N3B0Z12oAbYHXkt9HWqA2jnVj1kp
6y5r7gYwIVzdDUiie9tpJXoUtSuGAzn2g2qWgB5AkinxWLMHiyTyrZSfePk2tpydW8nT5/opHsAD
fcIIBcWcota0s5f5alGQtOtUUrC2EsSFdnoXbZueEaI3SHIYybvTxuDqMOfKA5sRhmCq/vUJ/xN7
gGnb3nT34cUyxJZx7nU+MLShdMVwGB3Y41Z7FE5Ktk/XasBlWKRei14UiiHhp6GCIF9zItousmba
cTZiFu5zJJUEU0uvdKUNfyxA9mEIvZXH5cXfrOtZppAeUGJJL20rr2LWAQnOSAnJ7BrA5jDoZMzT
kpYhkZEGnLNjor5aKZZtbxvFMc8tAG4vWz5xQpCNC/wY5HJZxDCCP+gyAD3bBQ7jKXFA5VrYoTKf
zyBsUVz46YTBgcsuLOBzgDDt/LFZBjIiQDsTA5hiFlpx/ZbZ0Lt8w4u0dH+rIV2wYpmhb4pjlZ2M
UguYwzSG2JVd8YUPPK+/AkVIyE2WraoJ/ofQ+taWs6SkgAWwg5hNDcogzUya3DyVke66abRhBHh0
gTv5jVgWjk+wS298dobDNLfQ5Ic4PHqK80ISBTZh5uOG8BV6hELMawgbxpI13qo+IzDDMvdzUg+s
1LODN8whq+fi9n6QbxYQntDbcSrB8C/1aER8H4Np0LsZ4M/RgaaoKN+lTE5LRf2DQw5pKVBWn7Kl
us5isL6FbBoWfEqWtJ1//JIGKLIY/UdjCaCIatBXIaOpyN+B5TXeiP6NPDFM3sRGwhE+5qwf1L8I
jZyccKPQFoIUNB3AmZbz7DxCRxxlCsI0mVrQsABdpe7d3fT+gk/8hXmN9Jb1sdBXbOBm+f1GUThi
GAFCq+Pz8Sl/esik3HuSdq9IQEnyUKCKJtPA6M9S2JaBcSezITpvyytrTzbX9+3oU/6ORkERaBPq
GtvrVrcSdzEQtb6J6ZWh+ygBAE7jM/uSqfh5TjRr9QDsJ4JhAjman7A2ENdoUHWWiUM81WNGKQiu
VYnTd6rASTTNpBMKDq709fo+9y65nr/5dg135bH0aWyf87Mz3Yxl6TnQQS8Tl/Q0HhmNVu+OunDd
RjjFi4jUAs67bD/61xK1DYr0ZlrIzZ1KMkREGaMOZkuopCQvTuz4lUSGqhe/lPmU0s4BUsP2dAC/
KQB2+n+/9KdFOPL815p/GmLTntX5ZCBsZTvNT1HA5m9YgFj0kvqWVMMksI3FTD83I0qOc1oBDQur
fG37T4j2uxGXoRUWSXNeWFh//47NavhKO+/K9kpdJexAgUxPL5xxSud72RCDjV3Iz1cMXZVvE56f
3DtbxRQuvULaUr9qb7i9GL4iOegs4bZtC5efnjUp6iGu1WfoYXymWbRtwK6bU05MYDEwyBg+To2y
6AWn3MJtCiGVEw1Wwo3Q3yWL2iWR/qgJ2vrjQTkOwIdC9spCrb/0uYS6sLmbs/wAEKPEWb5t/xtK
EgLGPCvLlguRO1sMPINgPzgQr3ZzMSr1sN9PyTmCyPk4+7+5PfTQ709k3j2LZGu+tQERT03BC5uT
z2MV5Kml4iA3rb6jNdYsSGyQ/2B3k4ir+LGUdAzT/7Nk/iQW2P0Qv3mzZJmIYRcOzzJypEqCmxOC
fGVfnII+rdc3qhWlLY94lKR1fQC0dKJuRF5sHOWNC3XMQcrEYXk81eUus4cffVZmoloI0QwhEdnF
7OoDU9fUAmMP2LKaNoxwKPvMAyZFaiWzOlEszOOGXO2mNjrwuCEwz0wNCwWIrMTVRmy0OYqx1DQA
qbNaGwJ5TZQ5jNaVrpDWPBjiePItdLQGb+aTv7vn35BzoVmCteBJCeelxbX6KeBQHI7Gvs4ETuN0
YK6dF8B/qsgGQaZ4CSo/AHfRUAXWmlG/I7oGOwxHhKgrfDOx/eapC98bd3nTDScfx5bx6DYxr5Ym
iTAGpeLSuhTWsXCpdvhiuxUijn8r3qm0YongIPfW4RjbIJnQDrus/VG1RcGT3wS1qAAThKtA/c6X
FvYCyvT2y6/1JgpEJCmqmr95UqjJhSvJYJNH+Mo87WaB8xaWRAS9XgUIGVBEQMTff7wtKEHZhyUB
p/N1YIqdcvS4NR6K32wiMhjgCulFNo9r///wUYYvgBzQJpflTM+eZ/5aw18iC/6ip60rRXWMe2xX
ErlViOR/E7RsY19TLeu7E765wIjlB6uVnt22rY506WIohxda+ahxc4TqESQ/X0IniJYdQ3RrhAp+
XB2NhvWQlZ7B0dYuxzagwowpTU1I1v+Qbr2hpPiJ7DERbHOJ3nGmHzXJ7Rck7VCmXBw2NbjxnBIu
Br+csIbCZp1ylGE5ywqtpC/ygyVrpJp0588yQj1jCpVSHDmPW/tpF1mqZHggv/xRAUjumbfPys3y
fNInlMBT4104KFdlawk0BAiYP/7rO/HbOvXAk+Fg+v90D98x+H4vvOB+jNO/oT4cBnngP6NcHWP6
83ia5Roq8kyO9pgUshRHVa9XJF/H8soWpLIIwHTyxVikeM8ItNO2SJVx7SHyyOOLKgkzUgsNprUL
thQXAaBn/Pf8XMoyNZJc4gKEkkH6AIVOVbRZIRk4ZRQqaUq4qajguHo+khqphpIdIMb8aJEYFRri
tWEbTePg6u8nGi2YQlvvQs7d7MyAa8PWnolYGBwOw3FiBpOZOWlQ2avlDHo6qJ6yYJH6cb3z28A5
rJNbP41nq87YtUUJS8WghlXfVwp+YEUhd8JXe6EcW89K+wGGXnb1DmL2S+x5/w0sg4Ks3KVIEVwm
JUx24FNzpygDnZe+1DYFqIQxHCu2tvngW0Uk2YEF+dvizCTue3VJw3cX1MGsP584iPCA8vY1qiQN
t8xgZIu2yf43nL8R0uE9D7rFR2SUyUZa2k24jLznMGdDxEFvTpSyL6NjroUxaOknr+s8+Ptl7rpy
8p841a8H2f/tZ7dHiGqp882houwRViAY3Xr6dfcfseBaSbsN6TKvoS0AaN3d6VHO7zbeA+kpXYcj
eRzyrSEqlQFSSGWEgBOC28fUrhQaaecVF6ogv9G3Y79BUj3aI1FqiyHX3crDwN0OOQFordY8GuqY
FqDT9bts8xJwrBE3rEnqw5o6fQJPF0xT3XoYnvIvT/VfZQcm2cO5R1HilHXtrjk+D/ANw5jp4lzD
WaiRNm4ScPVto+itWelxcrZeS1V9KnGKTZJN3Y9mQvb7WcGkV8Y6lPxvssC594WVMsqswxOCcy/t
VCI+SJx9eVIP3LtqrsVUgRkT3UFZXB0TTWBrzTEvXNNsepg5JgyYo2b1Q1E8a6LQh56POzDRyF3z
Y4VV1L3gGtkmyvWGMZ7EAoeUqG1GutLkgjP6FGmRkwvLBEPUgtbrfOJM4Ks0j+RldX5aItLCKflL
xu1xpL3+YBT8ux8EQYVm4iSeysacBpQfGoSjmLgt0sPyjEw5rNUff1SmDChvV7wnBT3cBFkkrEkJ
GDQlWtm9tBjJhxuzPnEJMbBP4seIFCozad1Ah49pbhhipJOYKGQrnBFrjt515l/FbEV0dbWlyCvU
9oVW/BB6WeghWFN13DMUt2FPoRukwCVrtCULS4oBoyRjJuuAKWFmgcWVZTrI8S0yFivL2bkzPbT3
Qz6cTQiljUzvl3hEZkrEXC+KuCYxOYNCfqwd0kilm0xV386sRmTY0H/ZwERN5twqtoTGhBabuV89
G4xuLe8zBvgqkE4p00ZYmAjdi8/FiIBo1A72ESHo2oqT8FBzWPv689xS0S42DDjBus1VLjzJRXJL
dj/JrmlgK7Y9iZaWUM/s2d8dk7UmP7VxAnjU1JfHJEXakIy8u3hnVlRwFvfDDgqNDIPxRVLjxPvt
XVkXAktNuVQ9WVIN2+kADdy5MVUg2gaWpZrNOhlIrFzD+Fn9z5rTMGtCbm8efQ6NkmRqn7Zb1mwY
e8RLc63DAsRVM3FltvEmaM17diOZClJjhH/1kQxQhpSOXXwP73F8BVcrKjkgIo1vKkrHIaHs2t2r
StJXUR6q1mD+RMBT0CUCaMhA/iEDHHn5I5aB4nQyaULMPS1H3nmL5dNLNoQhCXO9rf/G/ZGZ8eXn
UkBPFRih8ezVQQ7azjJ5BoOTvxmiNaHl36Gxfge8g4gnW6FRJrnhEwxEkAqljnruxxSfmsdUFme2
ycQueol5fIcdLRN8AjDKKpA+ddMWNxyxSERmFBF6HcAVIz5dIowe4a3yx/U15c/JT1EUV+QajnNJ
GFoq+CmihaTooUp7YQj99jpyauDeDqZDp0wCQ8nzEEJsgXZ8IQW24KIedfe6gF2Q0YRqouXPdMGb
AYAFHiieQ5bwDtDvCyDjdRZSOBzzLgan9vD3I4S+gnzr0ovlgYeYLTrcwuXmq12lYFW6GmvU7MIH
ig2ikhLfsSkemiC0w3PPmyy3pPnW4rqT6WKmudBMxp5VorU8n0DugTWCC6twxDqmicB0Oq0fj0K+
UywDRbLDRWZuWoyBivQM2I0VvfF6zanKS2ASdoVaYqBuX4VBVGZn1+h6pve49PPTVK0KFOH0cClW
QSSblNu8NzVXPHMAmCCLontluCVdDKyU/vO2ZdgwIvj2E9azCVQpC72CrCwlWJ2F+5yl2EqeQgAk
5yc3Q7ovMkKe6jPJfyiQp/ZlVad/2xspmNgvY9Vr9BwkV07/oumRZ2GDm9CWCJHUwd3+Inc/tff2
vabsJifJMiFxL9U9l1YXKIcw3hEibZi+7LAkARJaa7baMXz40fppR1zX6NzVfozJMBQNgt0VX7Rj
6BQVdoPZ6Mahvmgt4R0WQDVYF4LZM+CTTLLr5UPAZgS/3kFrTjWpmTFXtLbw6MUmKBcP9Ox5HtOs
CKqdguGq9iZF55m97b9idYRD6zm7SBKrCEFL7+T+gNDrA/cBrvMDg+BxorjDRhpWHf2SkrKUn7rB
aRZCR79KbnX/BnZFyr8ThbsdMdbEtkZI3JywroqMTG2XUIx00Q3UMqwgyf0b66h7fM+ze3fx18+a
yDaUIA7D8jyq7Pa9mF7vrwc3bVFKN08zfkHayAKUoFEmxxeTJnuwJRLJL5VsB4v3TZ9UOEFs7d5r
y00QgEmMj5rkp/BYxicLgPd/vRyEph00OQnxi7UWYSdpZ/ai7RoZo3fRC2V4zleVIGoAYof9ck9m
TO85nKZDKX+SRhMnFUzlB+3DMp5NdazUW4AAzoarCVvQTIHbiJyfrei9Dwdm+605Jebtys/mSddw
kLyAd7XyVsame4Yu5SN2wo/AaK3y38j37k629n1zG41NPYiaYyxDKX5kJwSRS2UlOewuqs0KXkAW
6Jz2cuTs5Nf/gG7zXjdC6ch1IoaRsyMdPJJo5sd6z5mhweHVXhuWBIsjr9GUx5pIY/ocS3pmCpg0
RVExc3iU3tmI2zndy9vKQUs0sH8yPZmXalK+N4qbZTMs6Z74N91WAm0TklXOx00ZtTSnDxPQu1s2
UPIgH69s4+Y8+GAvkUlyKW8D2fHnGCWAoh3GsxcvzqSZdbPoiDMbJyrYlWLPC+7tIQlJ8Uhcg81m
70lj9qNJajt9EIHpRMxRxgXLp36X2Me5WlJgOWKEwoaixIUbcUvdtWkqHw6XrX4OSS2t4oFzZjG0
d/cdgIbITp6mWr6qZc+MrS70gJIMgUMidmW6ysV1ZEvi+BgA85fqM+Si1bl6+5VueMRk9cEhXGhN
14wEkEDgOYk5FsHyC8MXEt3SHBQ8TdH8p0oly/U4VcfhWnrPJfjB6hvxqeLzfhNAOZWv+/hlRlnQ
qD/Fjx9UFfG2rPdQV3TKb3oa/wQ6P42rX5tE4/prh1sB1595tiHAvPjD2dQLBrdMNGxv2JDzDKOA
dn/QvtfJCenmGldCUUOVTbESt7sLTFMoPCUPfxNz3Q4OCF3gWW9Ilqc5NDqYttQkQGQbSNEAGDPp
W2ARu+PLz3qkp6MT67mXOGm48CX5kxUrOJpQbDoIPvrWkXz86xWsua9TtGXUYJH2VvKRipYFsreX
1r2ddjvXT8Zn9tB6hgzDociFI2IApeyqNgipYGcfioYtYSfjCGKC8Ln0e0FD4KIfrfBhizmsWgom
5YhxuWD4eInt/Kvj0Ip1JC9Fj1Y0Kft13sX8iNpPhGkFxhJp8H38CH+PYUBx5kpb24pISjgPEZK7
6UIjJQxQoX1BJ1cuPuK1uzzdW5wdB9BBCWgylxNzw7paCUT4lifRZedblufVxRmt5AuWvEEjTyAP
aPjHxNl/UM50yMI7Pq3/Lqwd5jxpkJzFlIHh/SxLnLE/t1uDz9xn5tVBO3rjqq0bt0s0YRfU+VfR
7tjWhxlOrAyuhz5nWe62yU9AQbaFUPa3urkrDKAlfe1Rc4znhucfeeokEKhL1SjpC5GphfmK9oUQ
634XwEG/XgibB08Xrqn1IMM0DtBgLOgXeAnrXl1vYB41/fE3X3FV6FENyn3LY5VCVDx4gwKrhCU0
qa0K+iSp7g+9LLj5bZ5a3nsQm9vZvQhqX3W/opA+Em2fFA+CbuRw+RH6r+lMwr6OsxX2iiBqjfr+
4EJ1oMTIJ6xyvBmcDAAoXipIKlDb/zBElxdr7FPBeMOvctCG/YJ/5l7J5qxICFMv91rJdG944MxF
fR0zPAT0vSJ9evBHeRn6fF7QtTsFkzcHwGrzRLaYBgIQPS/kkiDYDKJeamDW3BonslH2ZDZYHQpa
F10cN/UCUzwvtLAyPCffxzT6xNUlgYIS8iBuD/Lhria8UniJYm2JfUxxHi4LZZTFri3YvnzeRRIC
H3EbdQRChMNOBPdSqedN2v0Rjd2apcW1JOZlIsFdhVvidwZT2D5AgjkuyawVNJJIifG4iTuYdNC3
1rEmprJF3ALIH2Wx7Mhc+WwlPtDXyfKNZabFwYa4Xuc8KxmU1hCKJwSYqdmvrPDrLEukZb4WvOcD
QFh5MYBvFhgYghi2sklcIoQyDqUAA7BVacp2HwGwuI27TowGk7tdQLj6drgNzw7Cfov5koelXhvw
uIc4dzeOZvx9THLoU+dl9fstQ7gj3QpsgSnupI6TQvmCx3QR/O9CK6PIbtTgEmnhMw4L2E/KKDa+
Gu/5NtZMt62dTJ3utGQ46KiHKLnIh0TAzTbHX92yDPxQiBINQaufPrD7L1iBfeHbQw1eFHDgVsGB
1SqbEIZU/Vi0GjjW+iRTS17hjJszNIlUvgp32urtwAw4nZc8GUxBiIprRdKEy5X2zxumUhjNMh/Y
UTwL4NkDFJ7I9YuEd9NsVaMtmr4WbAC1WDItDYSQYwhKivaPduuW9iTXr30mYeWm39Qm6YZnrfWG
hU+rV9W/2sRjFgmqsCxbtw9gwx1lLQD1WPlG9y8TjCoUsdyihtiCBFyJpuARXe/mmnfzdHF6A96Q
pIAYD9KJvDF8YQC49qHhopWCQA/YaSXk63Ki/IV75d20GC4q2QE5Wv8minlviz5PUrIOmePijuYZ
U9qEqIq95SRM04zsIeOaI9yclkzXMPg3sMtI+wx8nDCOwic9azQElPzEzdW8C7vTNlCRqlcaZQX0
bRoCa20+oZBcya5o2uZKx3FnfYsOqnIajps/a8ssOuxPJ950NPbrk27n5f1DpptaIqOHoIH7qH1w
fvxyRIrtZOKZA1YwtZUkDuHhma3yCQ7dGco42QIo6bj4E409/2xlz7Zay+/Uyl/B7I4Yl07+5wKC
IDyoG1n4e1iPj5blp68YjknXqW0jzyNGIeg8E3b3RbVUQ9bZRGoEbKBHk5q0ySOIgOkfxp3VDBa0
OneCsg9E0RFZfv6RLAVFVjBycC+Bd3ffap55SaQbdu09rb7WlN5y2dFkPUUsNU3JBhI5C4XH0Xfh
n7DjivBczDXiGj5txyl3mCMq0OgQmmvR03zO3BMU8iQjNbCxdjksJMci/hh62HaHZNMZJfXYTfvx
QYYRmji1d6XFkR1+ddeq9MPCwQmyTd/r9lRGNybpuEitpntBY5fZSP5l6rywsA36xm/vk6IX+dnm
5yy3bomQKsVFV5RUzakn+pnV4Pc1wLf5uxtVDd5N20PuCEZT1YwenZLeH/2XRgoPhbXu7hM3KYpu
wA1sC9p/A88536O2QQhvmndXT6RFUVV2BfKU4MzpOlIDgIVGq2pZjC21DLQ/4EGLoe6JptBIdlq2
MNw9nTwraZZ+Y2aH9rHbpdSdw1OamFG4OZRnjFMkmtzKx6jCzOtzT6doCQn/GAH+k39A7E68G7KX
pvTAZCypjI7B7fE10V5nmPJ6JwP+2FhFdy4y0d/zD5ysLApBAzgN/hDmqXMRcf8flj2AhrY5B5hm
If5B+AnEMsWvUYupHZKWy1n/RJje1+yvH97DDNOtRikgKXpuf4yhI974eHBwRXZOEgrG7yZq2cXT
CdlMDA9tOEXZIZlxUsVeHLgX3M1wXo1h9Dqrdw8vRXD4nnp6NNvuVLWJAuk+509SFmCCKqiut5EO
+k+ENHFOcsvPCEKqcWW0fvzwQ7qup0J0mNmw+cpznt+a1xBV7NJZBzdP58bLdb8+E4/Kx6kuwDQz
1BPWFM1EmlF1Y3H3EnbCYuKIDxDw4hyg4sKN2fbBCAChXv/coV9PDyzwI9tJ81S8JD4ETTd4PLuW
aoKFMtfkKTDVf9FlPjj4MaI4RZxYoLbOg1iJIfPlHKnk8tRE6mGRWycvz7sZvNYHWZOLTGuzrZ9x
/i9GAzPpoNJyeZBGQu96wz1xefwMUfowWDRlS0XVFGz93LQNrVoVaG51cArfJbywIDhVnDfbS5BA
lqfcMVBvAWMsGza+PXfHCvQC452iWdRId4yWvFOtqBn8N432BOefECQGPX9YkxAQbFbwD6JQkn4I
byN8g3nmY08QATaXyoFtCGAWqyXaJW2wU0He9a/R6lsRJf7odmhSSDsLDokb76XCE2/U0uvZ3Hum
fhV5WCnSDBPrPXBSd3eg+7J0IMflaPW7Xbvb5d6HyLNrnG/mMb+S5Wti+eM9U1o9x9brNibezGg6
KGU/E2Tls2Gl9GV+yFKC71Pd8c+X2HULMbW2genFXb/VaxpNoW8a8LLrR4VPPaCwCxSiHOJLCpXN
3qhCHicCM961kFfKDsf6gcGePVDfF7HA9bEDZRSbePo3DEtYg5iBk9Djid+TdFARUNqePUJuR3l9
J2Hf1elhCb6EC39605BghG7KCj95irTcn0S5887sImIcDRttaTYuuuTAm3inwey+Aisd5kpQpcD+
4Tt9Wknjfosfm2TCEb3rm54lLySiCRu6y5FH6EAc2yvnDH7h2RJrdFkwM5EdD4xu7VCppdyQHrED
AqqZAWG6X5USMhEqY8ctx/KvCS8cku4gyZV9RbCVwOuglqF0OwtPIpG91BvQYo52P4qc2SuPI3fL
YsH+EwcOJG3/5/CpxsSSvEeYXnDaHiL6dpZ4WeEWmuTV+ajXkWkJG5cntVS+/I+/935wCCSin1x6
h695xI3nc/CEXQv8+kit4MB6CDYrdFUnWdEUajQt3/yrbYgp7wOabafN/m0dzt/biPH4jgBg6N+k
ochRPAxw7l7mNDRpTAfFZsAbaAdJDcoMDilV3dcqUJkYkGRxVf6HiF1OFEEZ+3GftqtRp3mtVp/z
iNYvsec9IcqYOUml6Y9pD+tGnaYq3vAVGsINd7DL/fWhgJ2xhcgG7tBUHN6t4KgOp52UZb5o6pka
IYMDItEHAf63fiKzoJkr4pzNKjY+SVmK16fyPUICyf63bU2yukYUwhlzCTlvkTcF5KLIa2u3lLKI
NmYwc4DBn/Xx+UkaY36WXHMEj+7E+pzDqTxjZhsVf2ogYHqlLPzWDswd+rkP+9Wdp0MNMPhZXYxl
9Lv5LAtoHjsXuISb2cjazm29+Xc4ciAIprs7AcnO2iXC6VCAwiKpOyVuOMDY+ltQ81Us3Mt+bbqH
Cz1XzGgyd0u6ife3l3GOJwmIBtRjtLKmJ5rhBlONdCTouu0auDQpYv92LJkr32TUKestefeukGNe
f3wt1IblDzBKWHoSpRMHdBHjPDqPUtLuWasnGCSypr2VhI8ubCPOMm28Riq2XpgOieNLRQVLMetX
feKkXbWd6vLxKe3zvJWeg9YJC9coWUZK8I4RHIl6jFP5/YArl6AvxCyHZNLhznUCSH3aExavry7C
jJhsvjgGTqEz39qJ9DGJLXfgo5nyJ3wjWuAcMRYf0sARSYtUG0FkeHm0txK910Rc5ez+T2TAA4B3
N/oHuKXxyE5/yK7hW08yqycVkznXqf6KEeSmbz7scS/UHawIdPA9ibJkuwfWgXu9H+Uzjs6PVM54
b7mgPr6aRMv4yp+9pBaYYmUFzMn7fxG3NOX3eYaTR/OQihqa+4urMklewXSqtqmzKgkRh2qysRbT
jMsA1oztuOE3AJJmEAndPePgLgdh5BSwpTL1lvLkldfylHdm2YJqs6tSOCMCqn2Ii468ycFg/WZh
d2Ltr+4xSyseKKLI27CcicclD+mlAiulaoJcwrd0aHMSi35ePpJ/6eiyDZ1PJOYjECtzFw2Iv9Hd
geUMS7R+Fo/glEZXFWWEij0rmiLYSS1dHxTZURz+qQAlcHMSf5ZtWvQ3oDQaxHgPgocaQw8lDatP
bdlFndppMKa/IjDL2gP9XP01uQ5VgMB3/k/ewVO/m1A3h/PwaRgoe2rL8NaUiqxtpZxH9AJUhQ7J
ZQc6YEhQFi8/XISJsCS0MWJTFlxemWb0xs7kjxLCn152AE5qsUIyETjyQFZvIb9v1MDNlrn0GIay
kbV7ahqMU9gjGF4O/I3Gz5uAsUPuhmGCLFNf0A6nIi9gEnjdB47uWWLmHRVdeOcWR0ErHc/OrPfK
fF4DLmk3rvelhqUPpg9QZw/fsagKgjgIxOTDNqWg7iGm3WwEE6Y85qsfTMtb191CXXWHB1EXOkJS
MEsAGGmo4j9uq3bm4tDFp+CqUvNsjJR3x1V/TU3kdS5I+F/piV+tStpSi18iqIaVAsomldp3w+WT
f871oW6JKfIESotjX61VShuEF3VoTtf6ByXUReJVf0l+lqSsVbdhYgceytJ6NQapmkCk4bATesnL
5HBhnkZo3a+HYGjogmQeSjLMEH6V84qrpDqpFeIpdQQ5YYSslES/l7ClzY5Z/rOBcAXlbOejfGad
GkMXD49aVnH75xzEX2+pt2oo+COrO/zkUWG3isgiTgxqMQyXq/tLLSMgg2VmiAj87yVg5Te/6Dil
YoLgvGJfeCxTtd65uMbu0CivqwRrkvzNVjm8857ItF4u9RJHymhEsfnFVMoYNKK9qhu8bDa+avJb
TzGfexSM+jUZ8pFHfhSoPYV6DcxMkdOEU1898/fag+ijp5c6uZn9yQjEA0xiMdRm/TWGhWT8Hy+U
uiVyhcJ+pSLtbFtfv0Hp9mPQ2U+AvNjivAfxzlEzE41TUhYcHuhZXci/81tbfUmUuz1eyXgBr29o
U7rN2EpJjNIAbTIbE3HEIVpR2m/5viDOpB+gva3PArSpM9HGCypxDkMkGjp7UFcxxN6AomwfOTvR
17Ss+VyP+hrJYC99GmeBuQcWHgbe48TfNDZsRdQAPHn7B/PyFeWL3BnP/p2k+alHU5f/3l3gBgD8
N5qWB9Uea2H5mTyltprXghKqb16v4c7zzcZ5i8to8iWbLgj5YrU7voT42BZ7nfD5/rUahXIRQf9c
4OCJLY9dseVyLxovT6wH5UFJQsU8zKjH6nCNB6ks3Ut2u2O74YrQMKa0j9hXL0Aek+f2Ui4S1YBi
1SPvYcbvl+gin5tkY2ByaRqncPRuekbQYI+KHutDF4sLnM6QaScJYty5CuGW6xHsTIAZrWrieJoR
7RUJmzhJY6V5dsmf428a6INjgQmU1xRWFvVDzHE16IVYuY5dDvpNyCN+XaQLzU8qL5n2qA1P7xXT
OMLs5gQniQE/JNbXL1pwe3dV3XGdOrTJudeTwEYBLYzxfnCiun1daicHsjT0ueG4Y3igDweDcCZJ
FT/ytz6fCByUC4u4OglAznOziawbPL87unwOPPUSQllD3ZUJG1Mz4XnVOXq/s67xZNi06HfMu3g5
r7UPY4cggZ2u6s12mPK2aCIRET+H0mT/dxEfXyIqILD6tfjXfwQvniQlFGN69kiZnkfkRZ45y0+v
hA645ucskxTFWreCYyfJpyjfHRCTmGP2qNC0FFq56xjc+2nigSSUCQSi3ReEDlYfANGkFqWFxqDD
7TxcvXK6cRcG2581DtGJDXZ2P6pdqZqabktDX6bhZAI00ObsoMqzESq4cQYZsuVv/lPqMO5gQtsO
EWWZAJKd+DbriEPWIyqeRZTm7RibOy01IF7ca1ViyCiEEH5oDTASFw+DE6fM2Tzran/XF866IW7J
vCUvaP+orELhUxyXZrz+sBL64W5UCjATi4Kj8NOhbAwPRW1HlVw5N+Po5BZGsR8MAUQrgXe5Ys8O
cvqk5ziytRGPASMSVRe1v2mDDQYE/xrIz1ghSYLPWRHbB52VRbdEqDkXOgZ6DbEvU/ZXjO51W4qX
GmL9xLuLNK8zouRCPswqFJc9ZnMGLfmzhC3wgXE90jSpmU36V4jhf+ZVVI2TAv7ZNRreuUQ4ruZk
tBAhq3Hnoa6BVY7HgUjV4qiGamPR1lCYtL9n7WIqVdbwH3n9axRE8epPdR9zGcKarf13XuCX792y
C6MOSYyvLsVxZ/Axi6BEmMx7BakdMVry/b9/NavM/PB0C21i1/LmNei6A2KCuORtH23/mOFQFD/O
ZiVf2Hse5HmfDjEJdyT9rfBAt0FbYAiGh5kfBQbD3Whb9jEGRgDBhUaNvY/1/qO9Fs7RmGzXdpPY
s84mcBV3xkxDA1lu+jsXqlVTxixNnLtzurS4NxqBk6KkwQeHVVkMJpL51TTf0xUBFuUay82SwAPe
+kIr4ocPHqxovAGqU7z0tprsk9ZYE/H2tZfrFokM/ZZ67uzqHuZleDGD0xa9WkDu43BNRsHyUC0X
l3ZXFmjHvzuGje+ElnWjGvsiPKBHWXCFuvdF7J+hZ3ysTexRMk7sSYiT0LbAn9Z/pMyxqswZCGe3
DWq2aU9sV6oBajM4YmUofhpvmRTdj58g/vYLY53TbjkkqsD7a+EupT3GVSfhXA8x78uiQCS3YBq5
l+eF9BlkMXauRLo6UToSwAFXrLJx9311YjhO05sn/dQNMQRrJvl4DH/8Os86cTU9p/ssEltoSXXs
oy72kru4j+050kpQt6zhJHDIKJ8B0vM+fFi7if+DfYHoDAMTbeI+/wyogrXmeQQPHEWG+GCg2Zut
JKogFTw+rYbfLzksrsh8Eh1xDuw+73QjmUxlwvmptuYMmntC83AMuSwB9h2yGP8DunenL4Mjlk/x
6khOklK0ZC0MAY7g6nbbLXyZJHvclAgAWSfF8qzA8MBGbexaR5ebcAQ26vXGenYoFcvlNnnQ/nX4
DUg+YQUU+wuNKiXQ0St70AQ/WZe90+SP9+zy71AVK/XuCp7R6cGloXRKm8H96PCh8y0Pqnxsn/MA
dSQjbe8qDOxh6049mlLlMOd6kWoOladXil2BeO8aUth88nVTne4R6Z0WdBzXZZDgpbC7T1fRYaQH
ZAgYE3KK+WyyzbhUT7PGXMNnpl37zdHB9ajDQu8uAwqtI0VJ93x2W+tXtnh9Y7PWbQk4jtjiOfNJ
gaIbOvpXLo6yyEusvvT9FOEucLyiJqAGzXiWSl7WIbM+Lp/Edzcl6CB8pNNfpHeBClBTMXqXH+wC
gYOX4DXb/Kz4pP+IBk3bD9LTlSFG+nawV3iCp6pCtmgpxSXjpsBV1zSRwW9Jr09n9QUgd0ekZlEJ
ofmZsjPi+N7/eZ1sUkWDUo4e7i38EAoOtH4/iWLvegCnrx+ykcObh12f1DLoT9EytqNsogdz681s
a/1q4CaEEtBs5KBv3YCl2SwOm4bn83itJyOcxM5t5g4XHyhmlKdAkdH4KOx9/5hUuUVUAqvsiJo9
nmwbmvcSXy9g72HEaW1vIJ0qyIhj2prs7mCc98ARKqFUfJAglgqqrxlv5SzHLcPGSpdmJsik5gx2
RdOE1VPGOPPxkyOeNGslh+Z/a5TLYK+PBlysZ4Ad5mlRwotHn3jPH+pckS2yTUNzqHOiuOcZ4Apx
WdKzgVy6gNSbN9XlxhvgL5GxyoRTFwCIBglUQ4KkQ8OJms/y1oG7oJvmn8knLbRFDuSmDAnasfNo
ns+dsjqhhfU4tN1IsWldIKOjP518vvHdWaaRXXVi/lJJhr/wKMFB0JZONAkRscUERjV0lvGubVOW
iplFEnOfc0Fwk7vkh98LkWPXtpBB2teVl0kK64wYNsrYaraQ9QrfaSbii7wNAsp2AqiQCgDllGCC
7voYfKe5CVpslRV/gcGy+E/lSbnV3p+trQMD9NbnMd0Pr2kwv5mwgUJQ58sJWf7kAFFWUVMeRw2n
+9BapzZA4o0rVD7xDamnbw9knE5WJquarVR/heJ6Oo2NzdSnG0teFABvphLo3vDJ0gWF43Y44En7
/p7lddEEYdsOoktIwqmq/Nalb4YHQXREwDv/uHyXiBBPs5hkguCB1fSgGzFpFtTc9SYzCo4yjBMO
e1TNl03Y79wMRnYO89Q/DjKMy/yiF8QetquvTL6mgxtuIHJRRrOTVOvxpS7Bhz6hKpNURfEL4PAX
fLYA7gp7+lsyFOf/YXxbrAUtSPNA9jrRvjcYzp53L7XGZ1c9BMAxkJ9W0AV9YTW9osXLs1HVYV0M
47+G+9FhtedcRreUKJlL1fnFnhbKb5EIdwOJirWVvvHslk4z7wzM3nPqjSdDtQgvYxwDKl75NLLo
JVpSVHH2LCEIUqZ2O+sfz5W2/kUyZG1D9SBTpAYcHbecP3MVOzpN74yOcmT3tLXcfQCPLjoqHD08
+yS6jwDp6mXsbJNHgiOrHnxw6ZZJGQREWfZgATWzn39d+FvjNFnTzPoPo6pEdue/sYJHKOLkSW7g
90bxqxiwd1js2rtGiL1SKKMR/JLOOceRG/Y44cEWPxxvY8gfxHOBpbzd9CEwCcrjjcMw+Kzm/1Uk
NhaODx7NMNWddOJex+f7SpjOfr47E6XtpImBG3z2l+Cfb+tr04scCTZrIKkoR1Un2Ne9izJI3x/q
+KPo37mRn48VklXzlFFJKTvKMrP8h/8w2G41zS8elvbqGx3QOZjw2MKbNaBwUfRs//ibhKdclp9B
YA9LI+ReF9D27Ym8p+/wj65jtUJ9zNidNGMw+1kvkc8sC1NQJPChZ+araCVqJtvoRpcFIPsaeh2Y
I2bo8YbUQvCeqAu4bJ1/EICTdH4wOoq6hZI85fcsBeybjtGm1LXDRGUG7YwS5hVxrM44qpu25btH
knNAi2Gg3ps52myIJuk+dC9ibx73fhH6ZAKw/wEKO1kTyIRxIswzqxTRuRxQakvE0BV+ciZCAUJe
4Yoemy533T/a23KsnZXJ6HTbJC5o2FbfZH5qq+IWt0jm/s9SgNzZXNUVrJ2bagyz3Kg/wy2PZKTa
tw/qqBnRhZKO10i0Ji2v3XhVgNu/OtJjDy2KCaUa/acwzcYYhajIJkjYQPqV1KUufdCzUyrzfJg/
3nLKUF8G5UoFsTzy9arPbWxt01aNZMczlkF2PEDlNQ0AqCx8GfQm/Vwdnu8/YJWUyIf5HLSFy/SN
1aKOx7zD7uGAOvrAUtkyjeHoV7xxkyzbPyhXbI3fRvXWKz5E0sLaFDXgc+XgyLqTPf90K3xjA8gt
zbXr5tQg0Q+0RMoGoVu66s66J5bUGJ3+/BeeCi2agOLHV3rqZhUONaOIegtxw4wjEShf3n5EnJ3y
aWXXW/w3g8SBwZ71u+NdE6AklNCddBQ1uZtyPX5CyQmhLNDjgXswRV/1M1Edd4dbetmR+YP9u7ix
zs3GWALVgnwiYKB4bWJn8ZjZHZbE1kk+J0Af98V2To1WuFtcYOxr1yYkarOXuEXBf1zgM+YaC44U
LYWZad6LDH9eOW22oFErvo3tTuugROMsjbGVTyLmpVIOEyVkjLkgrJDfEiwtCNHQ8fbprCVeJX4S
ql3fMYpk0rssrehuvFpDXaG0L+MaNiFEwam2mD5+xXSvHWxCTQcw4hxc4Av1O8+sEqNVlK9R3vZ0
RwbHy03zlRpQ2ne7PuWBFTvyXQ61l+2/ev2g9wnW2HqVzkB4mpTbhfiX5wBSyxnjIlkmahmW41a8
CINVpO24UvvADrnhHIB5iShu9W7fMKQcdy+/Dr5/jrG0vOR6MM4aAqUbZmtbqbCTgjA6FbhzJ61p
PKDLkiuSpm1APsL7OooMrq6BtoCQbOIHMaidR5eaGpMbFS0SV5+picLr6966Ne6gZqOnrtMPMTmg
DTB5h2E+T+NgMGUirzjyH3E/6LSVrZ3kvSE7Z05USnUQ8Dlqtc7jhPpdnxP08cvkX1YfSQOj1ElK
jAZKWg6+3hzhAuomNrj6x02OtMnpZTIlkGGPtwpuzDAlrbn3A/vZzisVHQ1mn4CzvAan4ivpxKPE
1a4PhVF9/zqSFo15ouAsEo4DBX5rl3yGKqJQt/i3vzNQ7DCAW0nqQweqAhk/aenXYDqxPZDZzKsR
52dO4V0eaDVTjiGLiMHPIdUyJYTB/rNSywTX1Io/Suz4sUUnfEKQymYGpmbYEIib2px96t5242ID
ZCcn/ml2P4eK9kvCTPuGKsrdudR4pPrXKszkQh3y65L88FfpqpShxDfGnuSSqRhwUGSOPrUR3KAN
1jISOX0LyFAWHcu3ZJ24v/wVkbHHcEN5DjjQeklucNk0aT0XlVOuVizNDNzEfwCQmhDKv4jPgXgB
yK5i7DdbaHQEdW3kvegrVSmZ5LlC3soldZhea+oU8SlHYxOSLYYQrlCnuQXIj1Y4bmE+pGWgBQKh
WJGpioPgA+1+lGWIq54nVRPbYnrbSOJmMcl5wDhCHnVNyZSrca1Dbn5rF7ndkc9UYOwMNx1cYGum
zdvT/EKgIqYr9gm3i4G7+xs4ijDmz1vrErzfPlBj6Fr4H92PxoUcuWdnIlS5KFnN1h7uquJZky9Z
C8gdEoSHBzbQEn1ITHYCWrwCPQgIzN8IFmhE5g5rQktR5h9Sqhe0cze3HwWFVBY0/q6GwdbTs3gP
8Euu5As1wGO1X2cGAnmY8CxOHa4iHjHbDPT0ZrOBj92vN7Xm1VK3PQTrL+txBG6LJ04faBmTB/Mm
sTzRJ1P6GoRZw6Jwz/dJH9dsJlWjv0tgrzW6NJ+8fSKpd/y3RgZdZ4M6oSBvLgBcO7J6WP1L0MGK
hUmoUB25jcWWUrtE6Bd5FJNJxMKWHOdF4AsDLrSckcWYs39L04SklFn21henF9O6YMRb+haJc153
/slb6gMLAalzLxYVbhc2OwpZXajZSszUUqS2xhFcDHo2jxWGZDLqOsN0vCKdxFHPL+2HJ4b41nVZ
nxklpkqiVlQbSR5syJn/swZp+VinXjiziwRk4KXKYY0Si4/RHuNjKqypMg6OMgKTsUNCJ/8eJ8Lr
HRZxNDe3J8DsArHz0HBH065v3la9LQaXZv8UjhIQ7IEIVlIzKv1j+ecVeiSsj9brpmppcj2bT6DX
8EpW9byWxELLVAHqjr+yVG7yAlq/d9fzLrVhchQJhN0Rcba72KOL1XPgYaVcKXWmMnUY5VOYZNv0
c64e1+xDH+Ud8WtlTLsWYSeZWEeDcyCmmBBEwKCUYzVDMNXaAX2LAFvdYV7MmGEV/uNl6iCOJHQA
+U3P0ZBel42Or+0+igZotKptKisazZ1TT0N9xa+2is3bIya1UqJFuCbhYs3QMk0LPrWJ3whWj/AW
o95J0aldOPGnwA8ZubWIUr800UjUequVcIJ/5V7Oy8AdtNAJFS0hIhBKB3Fsh1ETjFg319qDbLNr
i5luXe9wnmwVzH6TJZNHPu3xDJqBNaj1dem6Nqp0BkcOXLh7cxrNrCmCKpC/DTwjAsye2eMohKM0
nzFh/c1gqVhUViBLO7wM7Q7+Bix1d7zo4I8V+jUDFVjYifrLstg5FFtXum26enR6h0OnQJcDm70D
xrRZk6pdpkQh0HbzQVMK+sDCtrr2YT3bSeIbm7wrb0770d5o4GRhBG9J2fDZoOi7hA+R75Xhpaiq
r5hKVyrBCa4bH8LibmjWhUPWQQYucYZTeOFYEqbxiI4m1zBbAqUWuI0aq4oJnyDF8YD6iFVl0fOV
4dep1XyS4hCFzk9Ct7qTpfseGWI5PaddGPimC8WW8zFCOeEXa+4dPb1LHYfZF2Ss8/kQuN3k2jFy
9zcm/sAzvItgPN8e4ePNr2UI7MzoXcYMbS3CabSfS96mgsU2F/p+UY767WensAQEx0XqwbMURuwv
4dgNdHrFQIMynTlbTy79dEYhMzThljcoQCYWWa1RWpxI5t4QWoSgbi4lRn0UZV7Ql46dTu/6uHft
lcfQ1gMBH/YlOrwTbGnzbJoqX0Stci52pwMUgKlTYZRzWBDcF6mMM0PtBz2Qg8GPhyP1hjbKhjgK
ROBn8wY57LhgZ3qzdnITaf0s4rgAurHXG606UPLG/Ct1uR9+YdygBfzdN54RvdsW3fHWTbnDRFaa
94Ag3HvN1w/ZkPrXKYLQ2+4k+Mh+e11GAtTh4ENYMVjHE4rCJ2lpKvHRz/6xu4G87JSSxJaOtt2R
r/b6BQ0Re/eRvF1MZlZ2A8ybEZDWzqzrNjpqJ61tHCQbNp8WmudaFIrNwYIa2TWuktYSBUfRAiqq
vvyGRRR6gbK8aixBF6H+OPyrl48P8uJfSkjPBNQSbzxsq2VGt8djfqPNWmSdiEXgEiezMh8g7OJu
dPRtOAd9GQ5/mRA5ZQEcrolQjCeQpRsaPxay5u3pLo4zYEoPrwOyfxfKfV5Gl52iHQv3W9R2uSXK
XWfC1jR3dHh5piNKzImAjY+cVbcobisUOfy9c1dESbQLksowvHyJws976Z7n+Y0JIQB0SZBWn5/q
M+1r6RQ3CxclbrVgMhTWR9I+RWQNjHOPwiK/2jnuJQJTEiggN48GX+jCz6RtoAxv9nzU+n+9iLoi
JubB/NFe/lrxy8GRul1fDVFJ3bbWq2Yy3q7t2dMkbOnrd3xRpyTzMYg1VJQ8yqzrRbhA4Kq90Fs1
zfDwHIkCWNtdETDWVrs8VknavtK1D6FHmfIQh2ngVsBGbaRK8WuZH3k6uGMZrrXZwcDuVpcAvyOG
JSQo8RN+1ZJeJKqUa/zUEYsbS997Dz3m8jZTQ9BDBrgnyDCKX5wAcRDL9dD8MdnuMvTZWyp9RgEM
nHBI0wXenwETMEJzDF0KoHE2Ggf6B4/lTwkgWpxarroO+uLyIbpRsWHD5E0+tsr324+oF6zt/6Xj
RhnlbwcovE/U/KRroXENx8jAINmvx7mqq0hOnrxitL20EcmVHjSKCNsjGS9R5hLQPkuvhrS3fJxn
PKJ9OD3TC7eP0r+jpycOs+xeveLv7tQnSMI5CnVF5X5VsaIPo+cq6fHFlnmwpXDgG4G0D2pjFSQB
NGFBuVkkfrod9tWFUWL8SvCsfK49AKSWcR7Kk8IcjB4hE26CwH/5P341ORwBtoJQ6YwroKNPDbkC
aYdc5AEcrjt0YN8nGf69g4iHExmYnvbT2ZtMGiFBShMhND2Z4AlTFZBI1RqlAjoKkEJVZ/hmrq89
C8mcYvzd/U3Tzha1T2/OdV3v/omzz04NG7oszBPYDtY3swd1hj5pxQiGAD9e4bXHg54B5X4PW1+W
SL4z2jldWY22HlvlLh9uLWf9Y4ByZ8nMC/BpO5xfLZi3hMLQIRGKnlm99surGMuaWOucXcILVnz1
+RCwIWGIrZLzzvz+5swGJ/9Ogyke1x1CuS990JzdSSflF2gifEgQyN/FEGAMhIn7YVBWUv7qVRcX
wU2FOpWDNFJ2OfihhZkMdI825A6yX7cg+Oq001TJTh6dFRb66LjHOuEQGHGAj/pEwUVOkQMUCsUH
49PERekvtO9+DTr0qOZ0G/osaRaltR5pTEeRqGRZQoIlXmpEF1SXUg2HlvkmHvuKbiwaB3MRFewj
0Q/MFUdXQ1JKtxa7owdYcd/qFFLKWzRCELhxtPr7lak+VSNSN8sGMH0bgjuhF5Cb2Yh/GruGgC3P
doWDi9xD9Jsh8CNGAiKEbTPu7VPBegdrcgJeWX49hzr3xU4J3sdG/NSq+XG+hOHkBdK+Iq4KRC3y
0m++NK4yWHVfHSYJM6uoGXR3HCgway8DH3YO0/FIVov6hJi/urg9k9+j5toCBn9qNzgewmgqjmJO
lEFtLOPLC93bm6iPHu7bVGcsMR0Dcz/+hjr5YtWe3GJG77fpl9CuQ3HhqAAxiaWGWyCzXIV0q7Ke
co9vT97liZuHvSR7mqB0LHN65mDJDZJY9cxpHMhkUrOjhHW/MuOXFcTbZKBAxhT6seKq+DSz3byu
+qMZQSNyYHDtQNCYw6OY272U9Tl4JZ4RlqvlFTTBk9lAmBZwRSkAad/sqNI/UQ/gWrOptfvE5Yeh
MVlV51H4/LsYQP3mj2vZ6iq76U9Z4hqrqVVLd3n7/1kOtBTrAVXod+vwk46uM0xtfKakQW1azIuu
LDj3O43EDmr9RZ0Z0zJXJIozADzeekFjfuAjFKvYdRHSYx7ejMxJPg64xRYrxBMWu5tEOfiCM2UR
vAQha9dnBHhfxZODXbELo4sDzQycUAfc0OFD9U/i0cC5iY4dC8ZNzf/m+jSCzUw+2EmivRsHaUZZ
4Zn8p7Hnaxjx03NTYU7XIDCz/UNj6qhzAZq8GQfc3kNmRCrAhdb212AebOBO582/1mcsUDYOMO+2
OfstEUb2P1bcHd3QsDfSEsbK2rlvkOtkLdsTefBKawHHEZyEKExPvl+fTc4rjtJ0ElHX3wbcoUzT
+aIjJH6a181IhcLpFnDfxYd9Tvhe7XNq0Tehw/6uxYiX5xBVkTiekn99Fy+wF4dh/nTSz+XSbjo0
JvoLtH0EZfcDYXEl17g26Fqty7NcqoI7FnRCuz3fZAtdwAJqn1hVvZAlZ+AthTE0EBsZA8VItEKS
940m+LBe7jKSWyWnBH20T7GBMtT77G0Ml/K5KInpoesudtP+SZcqGpho+OQa5oCaVyVByzB2WNSL
Jy3lSstUIm7AppdjlX8m5bmymXGdyC5cjdQ+P4exqLVBdnBLOJ9kLq/zNzgHh7qyNLmuIkIEDekH
7domxXmYJZLi4QENm3TpkegmhRCEqckqddLHe0U+GmIApHy+9auGDGF3UtXFwQhSPQ+d8U8BSlQA
fgWSH5rZ+KgPT1MGvIeHHcgNqlG8gul453VekDVU0uJZtG7nfXYkE1m2ZLGBbzqX86tT8dqhcVVT
kis2egUh9f3ogSFW93lK9ns9fOHpvgF1ylISmvDhOnpdjtYLfTuVJ2EBo/f3wmN/v7M5wZZixb8E
mpFkQA3dRmiTxZzZrRRE7nxNqc/LFLeZRCC/MpeqxVJTo1hJqRj08vQLgzfuuGJUhAyaF1R68ybK
kKCiu0pL+OfKaxakdkMSPguk8pfSDnQtK1tjNACGvHW799dOKbbS+FFjAdWK4Cey29aFl8E9fixz
i6CGCzF3ocHLo74dUDfoJuk9HaV6ow+uJtEB25Jm2pX9VJ0zLNPSqLulTja9k0EGW6HLgrKzPJAa
IuWhrn9FolWE44HIRmFBoRdPAjI2tCED1yBy1JebwlMfEWIdy+5dwIMERXQKyo7L30emVi/1FHEe
my8l1ABUlnZI0CXCTc80WQhedMrPU83hK1x0FdbJdrlPPoQbswgqConGWSQ4fQDl2AIjj4QB/meC
ybQruKx0uTSh3v7qJAKP4UfgEf9d404kCW4lZP5zrLg1VLApwBM69g4t/W4flohdIsVxQW8cYo7T
O1lV2i8NnL0w4Ovu5gxczDE2vmN534SfyKue5YG7LPq8Qavimbvtf1ySWgRMf0vPeygzKrTtb1TM
JYrPb/E2XoGM3uwXOFMO8l/saMPrRWMENUsD9sRbEpLLNSTQGPw70l/ljR8OPLc103GNXFTHVe9h
5ucGcl4v/Xpj6Ojp37sWJW28kJJ6jlNMghOuB3K/rch9dZ1l+aPpXvkk+5D0qIa4iTSKo13FOO1j
Gsgkm5Yc3uWLRX4kP9oKg41xvQgSTxi984Nurp4aS3azlPfeI7Wg4opHSlpO3lIGJUaKz33b6wII
o0VyUmi7b6ZzrC86gE88eDaf9nCJrvC5gqHzW7P1Gug0FVtdFzazI63vgAULzNx+TK/1E1WqRD3x
3N0VOLaQFwRT207f5ZFY20AsqGl7GlfrHH+c3fo1oDWkJgxivF2IvlPfefZEgmHun/BvlrFfpoeo
24QbDTby4Sof8jeA92okzLdLF63vI3rEicCTESAPZsyNk3++G2JFvsNIntSVClrNN8PcQhvq/poU
ZB+vg1QEC7FCodPdMYh+/iMOLXxpUp4+9YabOvz4UiIAoadnreT6iPC35vwU4dvStmPYsGDKhtN+
tBbMa/47I8GsXYabr1V+ecdSnVcQIdWQ//e6c5ouqxISBTO9WLC7I6qX3HvvESu3Awb9E++nLisb
Ty0zzpDNb2fJzo2oOiv+Xv5rQ3rHY2ZWD9rfjMphNuzSj6WydvW1w5MK/lr16tFiau9cDF94/uIc
Rf9PNoNga8CHHqJ9lGomS32MqZKBXRjn4wlYWPRTJBAMSKFRnzI7TvRkSzr4hZXdeeYxKWiHYI/b
nj9rl8noDenTDIRV6bkxou9JsuyvoLyOx8QEvSLZxVnBgN12Wvcc0HL1P2iOj/sKWfx2hRYrwsn3
9yts6xtAzHhEoa8T1LrqzZleosYyAJEC/Yy0dNT/oekeyVD11jDrMNsw7aUh0fLx1HfrWnF7eNv7
Z2PJP/GlpmHEtetXfdWu3rbSo2FnDzlgnZM1/D5RUMcx9+kDPh583t7jL1w+WPRWB8cSqTpryPiW
ZbsDZG6C+YOhqcuIPGs02Xk0A8J6ibw6necCM8rsN1wx7Uco0R69OLmjXCpd76y2zG+W0ND5KaHi
8+OI+L/D0mHAmrxi/Nv6wBkgslvPmK5p1Yf+54e+ZD8jG9ffIIdwiaEthLC2vtkekc19SkLJUoWP
hlhCpPLL1c/mJ94fTyZQiz0LKmbiZ5HvbcocZ7nHyq28nbc9gWpNrXaTndaYQmcBI4T6R7i9Oau5
lM6unFrUzFzX0IiY0cQYD2U0g3ibYrAS77R2AS0OIy3gCnDcg2rXGrhD3vbXJCkjOV5CA6lyrB9f
ZbQQTz9udhoC4sfCrCs9owH9etskStbG/TL3rNepWIQD1VjkQgkVvrctpVU5PRjvQjX5dnD4oL/i
4eWWHRyhzITcBGXlbz/CkhGhd6K7iEbydUZ00Cu6KJPcVHGPe71vbZGwcM+/sD4tdeIpA3+PHtPp
7lAteRGyLt5CHLTINJIxgjSn8hP1UkJIG/kXXrq+KQe8RoAafguK5EGhEpn2Vr8yAS8QofgQwh47
NXaHCyHDnfKGSKod7xJE/r2LRmNJAovV97exm/SR8Azq6krETwh/son4zZxGoPAASkq4DGyHxZsJ
c29VdmJYxLnk1KMtj3vbOJVNrbmVI0ZEN7Ekf9fCT7S+D3G4C7octGNgesMKK4dTUZ7OGP0Gnqev
AwwmeRRifWdM7EgpAnvfRPeq56dOk9ZUb3rHFzReKRdQCOugzjdHdFaqjbYLXbzIM23X6gL/sFah
40X0emG3UVnhsPM01pgFwQcH/N30oF08Bexlhtcw0/ocA8uv5N1XlTbKYKFnEdbg85SzL9miVCRB
d3jT6lt6LrEqDHWzdVSNP/+e2DT1Q2RUG7c2TyPA2Y5GrAOfKu2azJSe642JYfep14UZhGsao7ba
m2Ge4IBmlaXAd6b/ZZ1/P6y4KzTwPPi9NefCrtrAQnIgBjS2fT7rVUiyfF5Ut7UdxehW4VTgtVQr
VZX/scDodBtHVslCUHThRLH836ca6pBgQhNvXV8/G7gzmSXi5rq1eSgqb47jWE8CABGfdWtqWAY+
Z29pBinClfB3iBGLVnbhmfRlh0f1lDtdkzRS+y13nLTGSy35WbikeiOf6nHt6sBGY1SJWOyfa5MR
sdSwEtPFxyqZhdq1G7qgljCZK1y2BSp9G0gEoG15cZYmXoQSSQWgeyOT07CV22qGfKZXMO05f0nS
FJ5++p2W5E3PI7ephz/rtKqCZBx4oZEHKM6Kj59DjBgHOXtHW46EkCWkaqinloq+sRRtT8zVNnjq
zlP81iQduxvg+qdMfZUqiFW6fYAXMIZfefxwcZhi3Fk38t4UoIQ/d+gTPDWR7q3SJEvhbEcC8kxK
80xZc9MR7/xvVE0+YJnzzHdsy9zVdnbPU+Le6YhmH6FqZhsgRzxMEWXQb0mtcEetIXCAOZfJab6k
3c1GCNFfhXEBTEHr3TI6CDe3syB9VvybhGaKgGFzbSxsdS1Iyl9uGnITXnpAE8yvNNzjl/R0cQfk
6FpBVLKVuFJW2pmZ8cnpUy7BlGOwjdNiYHM6HElyk0TK0wgZgGvOE7v8gbnFhwQsKTm/S9Lo0S2A
hDLxlTtRkVF73+Ro7QeJ05o1e+dPE7ig3nnQE3Sm/OzNbGICkDYgcnUrhuyQTCfJWpDUDSOguZWn
9b8tzyqSlRokoVqSXxZce4WTONlbY3fRSEUeQQopqm3gXP07DKBFiiSOIyJASaJFj537o/oOjnMJ
HZpdiGATn2ntPYAWjQbaq+QENfslPMmPjt3zc1ciJhjir5GMMzBA8Gzz9npMNA/rjGM7RtNWYwve
P3zuOS+Vp80cCmb/dJceXE+nUYfspOQ0qrcdNZt0OGugBGa+7VKVI37OJw+TgKVUQ6zQTCtzg1Yi
Ct/CgG+OcqPZYKbksivfM5toh87naWm+pbP+2AxgUDs0rP3smA0lgbKTjUB78ppJLK98uyb1wByF
xFnTChRXnbXsEtreawcIzGHlL2hwvQ63HgTC/wyFmVnHBFYsHec7eLt3H0E2YqnZqr2JXPVgHz38
C29jYzmAjggg5+/yxYBdJgTtL5lTXZfflIDpk1dNHrJIi0v8bai8z8JuD7zEbOBGbfAiKUA0zoNn
aSZiN/b+5SdRN7RJnTIADKQpC48doHqtRmJYE7VurBpCdborFuVWTvn/o6x6ARX8V4YJcw0tFemn
touWNQGCNHixdYVWyNjI2cipuwBTDdUU88WWceFd840BlT+zYiWBFCO2i5cwcu9ptP5Zy+luC4BC
Z22EQHwAFizLHs6fwtFYNw8EZjmC+toFuloOVPN+ZFCwSQLt4U173iCiJxQVXgY5DJC4oDg16kRz
oABn9ISgOSITEakWSpS8uAxyvGpJhDlYumJikOIm5I+EbSIX354+sOPfvnuq7mNkmJthpJje8+6Z
kF4C6Z2akwU3AvQVbOMpZLxDkaZsXPVOTsYl87pcGOsugxJSO73je2UPD1BOIGIej9HjDYujpm+C
6VCy2XUPKr/AuT/vuN4QIkZcNBGS/Dx3kBpqfeAIHEBlRpY0iWhwI1d3F4OqlAMJ47PTHokiWVKh
40lTw5mSBnAXOsH2hGKcbc0qlbjpqG+42V50PZuSu5u1myxv6XwNuQZka5H47w6p3EualkuhJEPp
8Thn1z2HKWa81IAkq51CzLygfACApRy9HRb+j5QKqDUiBnzySOhx4vDINtuxKVmWs73hd4z4OZo3
by+7d7r8Xur7F9rUUOFM3pp0L8IJgBZrig0zdKOJBayK97IS0+nYUOSSmJPCAsek2nKP/+8QnY3q
eXJBfCd9mu99RV5ug3tizgk0sgPeNGEcxIjLvbSzUl33yTsxFd4trFtp4BH8gA0sXsj7sRFYLREW
VPaIHzwKD9sdpfsexzXs8SQdnWsZikAzXNoN0mPsgne9nflsgAQW7dKoZOKQ7thsZSEK35YKD/j4
Hp7RUAsz4dtSP23vAcFIrW3LNT/XewTcp25gZXr++2GnTsJWBbgQsoMgfdvQNzAiYt8mUt8PdeV9
V8W3Q2H0vSm8Oj+sBHdJpCJ8VRbhEjOmxzn+8AkpKIVaoHr9Y7xVM/1iK2nScHVvLsPVCa9sUw8o
knhuQGqJwIOUlbrIUX9nPwfv3LqdYS+dmZh4n22T0TtzWoIzJUeZyBmvY+iRhGJiPD2CjCOezLcW
IxF8R6fmtWa3gV4rL757GvTUcpmRI1P/TAltqpCLG5/9ggwfcyLANR7gOdYKbES7x3N+sdCrhiji
wfwTAWh/ydKgm29Eyw3FM42373/tFHoyGtDb1Ns0fSzOFuaU/dMdTjXYBhKFpoT+bqHSNAvIwN/V
pU5XvAkrmw7vmC0GXMNXMjAqB4G3n1HsTRtbvzQYcWSUynHQ05/U9JKkRoAXj3AqtFXS1KOBhjzJ
/EuTHQsz/hx2kImbK5YVOeWjkrlHciUFLYi5yNyCHedHz9d7k2f/VA7a+9xWlPtVZROST+rzZ4X4
xPIrD93KpOQ4VYJQok6SDw0rw6Fplza6szJYaJbw5b/h+vJJ0a9qNGtc0Z3ov+FwMf2OUoTjkeZV
zuXXrdyhPph5J+LsbQoRfRqGi2IIkyJOAEy8Ku78YsqycBAQr6/jS4Sa8bG5n+oFDDqw+49P4F8p
xznYVNN68wUSXJ3QYonvuQ4hB4Lip4BYtENwta18ouNmATNgvgKioa5ZowKhU53fhoR/z86nFbPy
UB0Ouj9+HyNCdfNCDPMK4duxgFVtI8zMQEzZqMg6B7QwdBDhhmZg+FYCrKTHOwruciInxOGMbYmE
atBcl+rBjj5AR9XjCQuyaDolKSzdSk6ba/mWSqA+ItCaUBLuZ6Vk6XFiKVenAgK6d0GDbIy0yaZe
0Wx30wsJy9mfO37uHqW4BuE1boRfI+rqs3kgVRotqwfRobliYH8qEGw/R0oYCW45upixpvIaxWOH
AtUnVf5p6onuEK6/zWRtcq84znzAEkGbBTSHs5WaIsg7pYTIyQ1dP2J8SyS7U+tt1BUTKizUSSU+
+VhXr9N5t58w558hQGp7RkCv/NjGAutpk7BJiEl86nwhCT+UdnlrMgN2e4DPnVD8295OgmRk5Ltb
JMZtMgK0iplM2/4GPrZS7G8sAbxVYkyP8G/1ndZYQb+Hx9sePBZqUc12/ARXRRAfZpoNOUycyeLn
42pnRxJFmKAPq/ZEpulK1T7UekGYGQUlA2WrYVKVy0yhmzhmHu243z1tXzvP9tK5n7271ABvE3zv
W36zws8fvIX4vMfA+0duwaV/hnflI5fuC1HfGjvC43h8xJ+aBHKQea8pzDZpuIOA4SBVz4PF1rZQ
kOzJI2CSTHl2xL8vbQz9ic/LyqzoGYqXQKhiXl/kBsi/yX4fGoWSSzv/7eRMhk2xLiXDNv8AgV5I
InkmomNliRwPw6UDFng7EeqR7n81gA+O7Kx84UDNej8lCthmTbrcW6oK1PqcChLngHHGQPfT91l6
Kaz9xjkhT4S6hwsHb+A2vEkez4ZrkfT3yV+7240VR29rHHcsPTw4YIxuj23bhMRU0faf9OyVc4n8
N++O8pEhnUUxzSMX+F/qcw8+Zpx6rk5x3Z2TgNRi+bCLWLVrdpTtZeIrPNTR3t7qC9ulpv2jWn9i
yytg0oxAvWuIcra3fAATIx0s1m80YOH0RWwiLLaXDrK5H5z+23iX+I9G9J13NrlGR2RmgMM8Kodg
O7tNoGoVWkmkZF1x/anQIus2nHIJN1Q/gXoLh+I3UHIFJ/psyCyqUKCs4NY3smNW7v5XfISdglY1
AnYehZCjb2V+C3VjGdyT29MvXxyfty8dHm3fz8tZtnFJ08NOOsSVH5pRmDdRZH4RHVrY9Ja/+Jmo
JNzi7bkNRX3gCUxx66NMSalc9AjGqJY0td8N2Y54GMTXM6vthz4QBcmAxWu7kGIVMTesIiAd/H1y
c7zpIqu8y67SJ9h6J2fdnGS3S5GckQrTl80hdK42rcCwVX2LT6RDGQrfyve46uKYMB3QtVPB/LAV
yfhSfJJePUQVI8V2XkRVrOqehaEcZE90BkOhRVo142T+1GkveEsXHeK/rcgsM/sMd/EYMXLlNGWR
BLkXkSkoYrOw7EIDhT1ltRfdus+qVpCisJukYfNaq+rmjR5YTRM9iPjHHbU/12Ym6hRGLMvQsKWL
d5MnO/0twTv08WZjRLhe8VRmwxF2uPTYnWIHg7NHoWE46T2/f5bm/rJDkjPkL7NunzlkzbZpJT2B
m4t8Sfzy7uPxtAwiiEVs38qHlpDVWL8slJMZ2NN9Ze6S8jIDqF04ErCTy/ThjYa9USqUp3ZK4hdb
M9wB9u1usOFnMiqfkeTxKjvccpCReVjm/MF0jd1GGTB4fYW5pybMOzDzyuwy3F9xssE89P+9AnOH
5icwXcavPaVHP3a7LEv7L2aS8UVv0ctIl1SFdpP5/F6gzzVdVjO9VKMSpBnplzSJyzMjiHrpCo1l
Ow094vfSl/l2cI5OWRDrpRHSnTtPk9I6cnIqqvX2beIXiq6G/Dcb4nydmBI+T7li4xqkG/qLlB+e
vrY6EUjvqEfxZOvz3kp3jBj2oX48HUgZCm/nmhVHkLgMK59SkgPQ8sTeujM811phB8JIRKcL9C9N
vk5qy14fEmbOKvKjNayzoXjkjArR+faEBfIR2eShqeSQ3li9ZnJNTaFE2X38U+BQ9kTya5mdxRpo
KUYsazv75ng+WXw/HFoZ46F+Uq3MAGowkG1Fycjx//w7ABpEKszvRGfBMEmIB6Z64lj8QaIlrfhC
8ckKoV0Lkzyoo/BocKObda8Vobd7srfunDH+fpIHEKAy0dWBo6evZcOMh3QWt5D5F0rfYdR49o+s
x/t4h9UKCbHRQO3EKnsahlNkcTtGJiz8ASYDC9TaDsGHJu9UWntwXl5kPyMzlWcEKEhOiWzx7Bzb
OjTnPa216eUMyyyhpE8jR0EfaeskT1Nmb+vITgZZhnbQN/GS6PEOv1UWvlv5RIF9+9lVdBHTJmIJ
Cs//H5V6rZ8dm2QZK8BJrrpu3WPCfyttRfe8fvXXH5JA2AV9dpk7AfgKoPfNxJK1ptdJuvwOtd5B
qoCSFcuMuUaEmKQCUgzzUaKhlHZCp5iYfkE3ZcY6PFO8vrbIkp22w7u0UDKwynStXACIfp9r6yDU
UByNytvEUKvrtDV3GcQsH9Er13u07NXAtB/nWqJ5mIbTEkJvcYMm8qxIM6mpFZdLTNoedgH6RbhM
E5DcaGGwEAv0A/vqbAha952DhtjsHIH7kznrXgSZyafEcMSU3zIcClwM4BMFQEcwTDvm/Ywxw/cC
Wzkd3/XXgKgMry2QfdzCbSMx+8IQL3KlLCLvXTjxZn8fVeFfKbIOm6Mvr9dXN3dQAqaGKe906vrK
bs9ROLsMrK2w6kR3XLv9JGSqWik1IPsrXq3omWzkbs2BceoAgUmjQueqVp0/f7RnpgjZ2St6bg2B
rSwgomfM53bq3YdPYQccJeRK+tPlKJih4ZoAUD3Fv1TjdVfu83+w/S58uSpGyjysg5BOanlNnw2F
jENHvdzqz6NsAPylKE6KGmGRudO//hILTcEdGoj9dbq1tpIsKinz2jxT4et6YdvF5yFP4SLHOpUh
+TbjmjPdR3I6AtS9OYEnonNclsyVmz5OSNWL+CRkB7ZNhi3tyJUMb0ysGWrO/SIt9wvljWGfGReR
Lp3Yszzbe8DPasHhYPOU8P5K11qLg7mm3YsyUWdlGRXfexdBYpIMLgrCktVABohNBev33VFPV1zH
saI31S2LGaJ0ROz3SpIF0tv79m+vDqxI4qkOduXGvYEZGIbUKndnASF0xjPsVIra9ZyrmylVPYva
Y6aF9eobHXvJ3WV0nrrPPjm0J8sCL6OafbEuFP8FcYezzGOeyJC/WOBNVtBcZAP9b6cORMHIEYrA
F0wOuoQZUPW6lZQmPmcmEAmKzmZJ1+Nj4FiZyMPPxb3c+pI8of7fVJFE1B2xOGSJBq2l0jz5fvkf
h/GHphoeAzAVLm2sNnQzHP/XiUdye7cQ2C7pjeGa/XXpSeKKFWGdR3Q3ti6bN9OFQ1J42Ock4s+3
mwfWo2XoGbewad3B6tLcUjVdDfKUWxJ9Ov7jw32+t3wwD0rMG7ZdrwXQO5pkLqxPGlMM4FErlT7d
YHYFpO8FCQJBKxB5PXCwmmW37LKsHnIjhdmSN8dUyqlVzOTuAPsFvpi6nqDqc3ilYjteZo6xvXOm
9R3+UTqpQ1RtM/9B/zFvsFy/SzDy7wqTolOnSRYkZdDMc99VNNbZuNqNblFqkXkhivW+wxAIZikN
IRJSzncNsTdUpbtOkY0RMZ66GsIiBj9DL+nOV4v9jqP62CGsMdf29VCjhL5LLDbPOkdKmdctTTZp
KCiIJHsCaJPPElPwzmGkNN3oe/c2huC1ucA5Gu6FrZjgSqKZDr9NIznBupPE4IvARJVF9Bzx79hQ
EoAR8aFaPpQumeu4/HWHA3aSTTaldwKctoEiO4mxAJFZq4/BQvLVAiuqLUnYEH/RwsQ+QGeeU88v
IlKIWQqa3cW4wS/DaWz5T1GoNyTWwWCEzSKIIZbnrH05EO7cBjyMMWkAjJJeHzdWI4/tiJ5tNoF6
CV8wylPCZ5I4KGZ82vCYPAxaAs9rlKT7/F+LSs0+l/Md/n4llp7E4jHnTythhtM+vJ02Cw26XNHh
Z+YlKkoslHEEuXoLploqkXZYVA5uPqSsn7CwfbssMkKLknc/9OB3GKCBmh7YB+gBRFBrngeLFmQE
rJVPEatTrLPNLE4yQU5euSE3bxig2EFkOO0y/ZXdE3zs3oWkBH+cUdcgpkk35sj6EYG2whb5j1PT
mxwMJiJP6cT67ZLGEPzO6Rk38qZCMmRstN+KjqaTlchNSWeMIjp1r34gxWKUKRBwjqiB/ZxtaSPt
VJcr2TgsMJz4ARjTxN21fo4vba8Q3az/fYEijsoOKWshw+hU0HybTGr17/iG+cuw3bnxhj4CPnJh
vZbcPqd4ubUVq5cJo6+/z7wiAADva7qUkfZKUXgHY+SBNYqFWbfNPNZ+E4pIkyTXTW7MSXZ9zzz/
6yJ93lLp4c1/+weKybNho+PXyuRXMrGro9ePzyPOwNZJ4V0R3Nh2oaMRSx16ukcVyLo0f7Uox5/E
0mJyMwXtfAk2VqZfxXEHXKBBvgqCMpAkR2BmkQ/1GGVLjTovTpgfvuzHt8dZmpLV+fdRWBkirh2i
Px/IgiehDuzaDV/zVhUQpFxNWWkZjZJGYOu/5TTpComTEPXyKZm02K3IeNXURtdQEpMqPe1le/xs
MgMjL+CG47iAY6/EMYJ5Z4QoAEiRR663tFgH9dvyV2bZWZVrQtT1jYfUsdIKzCaqsTFRq7h8yGlJ
ARawhl5hB39PFXS4fEkA6tiWx+0oAx4zlVssGCfsM55luOoGGO5feav7NO9f3N1ynX75Q8TdaEP5
5En0Dkq0fFMF+Icm0yQNcswZxuabbAUMmT7SU0XcP+T7ZtkIKY0qIeym1hhkfEPWIy2oF3B2do58
WBEzMaCu64PCWbzmL3JDuzfQjs0/FV3BBUWxftxJyCt1LWFMonFTs1sDX0ZPeDzR9dBTBdDFuGMa
s5kwtKU7e4IZnM19JrBU6QYEFIco+yYSMjpuH6gvUI2mkWEs54HBPL2FJq0nZGa4Gu7HEeIv6YNh
IvvRXOPnFNtkbw2RmgSsAHB8Vr6wxlNAkqvGvmuMDmegxr974WqmU7jD9TFfNuj4Q1XTFMP5RPeD
YwsFqd4qtmiqOq48jZ1SWJbuP0p49fgVW/iljoiDWzm0W0ALJkFGQ3D/S/QGr0haz9KDe0t3m5S2
tqx+3R1C5WEAMuGFiZpMuVUJIVqiGz+pXGFcsuewUqhJAvMMmCnAM9rkNa0cFwuagRTo9qxqyaVh
emKbHzmacbj4f/nfsB60PrzzjdJoFAQSlgoW4ZfCaCoBrLwpPEdkv0h5aGoP3cY9W6H/mgj1roPc
tPbej2L6VOF7inJXnlKTwYBZKQNe4s3DcmcYImhZyOz3vVVJ1nonJivvTYRtbQNVTeQv1/d0peer
PV0Iy6nO6ei4zL4D33aNQbGNOC8oUhJeZ5Y7bUggA/Z79X9/8crhiiehIxG6SdOWEDKJsEOYbxSJ
nMSGX9r9LI9b045PePuybKEidAma2hFKty2/eMjOR0IDQKlJ5Scc9vl7g5adVjt7SfFqPBYThadW
3zgurjAmVWe+vW0wY5/373BThobSdVB7jJXQSOBjFkHbeOzaCQXPqpJQ0dpKkc4RqZxF0I1JiWS4
Bd1RLreRGY960jpLVI4PqJW9axSaTSsyagQIbYy+lrYDPB2lVZ96uNo5CHnAnD4T9IPWxaUkrLzL
/Oi2PV94IvdV/L2VvB1hIAvxaCrPmUOwXO/GOUaktz3aSA28sajbSRj4L24bFEZXnHn0J/4g6Yjx
iLDCz8fy9LIbLkY67NdN+6PylAac+cNWipPHKfA9UIXEQ0KPjzhKQmjOfb23qbUkFpJOCxVIcuND
k2SypjzNz6Aymohay7YP5zITgGb4pMjDrntOYSo2LM0rWEnDD2z9QNzrXkL0+eVUe2kuPy5IyZFY
9VaEZ76e08nXGCHpiJES8EYMGfE7ITc6q2rV/6R7pBgcC2FDyhgoyUTDkFMghBhbtuSfbJxqSrNn
wIF9qyy/qY4XhGhTv7EC5C4JAPoVRjrdSgvVKdp53bqkoZtcyJ6pHytDDuCSLdxGHib3Y53ToVCp
cf0iGT61pNj0sU9y0xiffKvB+uQ3Xia8VLeM3VcTOeCcEQEpdiiC0gYX5BJYtY/Z+dzSBJIicf5D
dr9smuFTVGjUwjI7extUEG+lrxQRBU1TexaPr2G8QS+4yRHAOnsxNjwFxPHOzf48KwBgV3RLc/5u
wRHm/Jynzzbyh2X+OoXZjbaHRcMfp0bsb0bpK0BdINjiUdb8tFJnJ4hDNIgNTS19axgZSiXiuLJY
OSYtZPC+zISrsfZyVTiBf2S4+Hh0Dn7bPMzxaU/tzUI+aHDKu6InUiTsjXzowRQfAJclErmACB+B
cYy2t+wQ1sRzvQnBo8Y0ynFCGPhW+WgilgUDEYZPALxwfRIBmwtdg8S+4dAX4IJIngbbmbFVIq0B
DHlU58TVquJhbQGXN7+/l3Ix4/V93EPa46RqY72uJ1quqDpudHkYESeVSVklkGuX+owfNJKR37lo
es/hfDIXe1kreGJFwttWfjK/6P0ig7nZL2TJO3WSCWDjKVD89vmYtVGW3MkQll1lEV60z+vQtgtS
UFeSJwhkZ0seDKFkmEzc5pFPoUlVUAPdysKYQKMwMujLoV0OWg2/4LqpDlqDgajp9T2bt/5TzYXm
YuI+6Eoo2TV6lRNNDClo40Gfvu8+ZOZX/DOiU3nycCXXKGnSYXLKnlVQg55SJQLrJ+eflBdJwOp5
S0M4gyZiQUgIot7KX1Gi81XMPFon0H6bsNLwLUk9KNu6HHEYqIVLDJ24EfsVlphy3abMI8u4zuZ4
Nf/l2WKojtAJBHQxx6hO8MnR24ZCLjFyZ1IgR68v23RjiQpNi0ythbGECa72SIqcXw+z7FwTGWvt
XHXrJbU5JCheTIoGappQC0uYqqUfRfuE1wV+b/c8zCyD6YYkbxstUn4PJgYk1+6azJQ5A101ySqw
nwol9X1nnJwa5bdEwS2s5xjm4OzQgr+OxZZDVvXMs3Gq791Szy3J7ALM1C8/Y75V6tW18iYSAer2
PqIeAJXQJi4YuOqPQMQgR2ysl92b24PNZU/f50Qt5//K5FT5bCjRtsKTN8BGPju9/xmhXOyO0Vg4
F7KJ6kTLZs5UcBOt4APHvwUl8W3NJ8DS0rCxegBMpYbY4NzKbvGsz90apBaxOh0M0hgM1XN2I+Ui
yFXIBvGea8BTlo1kWk7kpQABSVAErgMZ9RJruIZm76A7wepGXH2KRXNTxMOqQmgcWEV2EMaQO7+Z
j45gxz3J87XLNPg8XvF3TqJM/iSGhGBJ1xTxGQDnqoogI0vElIyMaFFlJ+N73hydYBX635Novjh3
YSarDRZsOPhuavyIxRblUFm8H1YmfMIkpoUgVH/ztv/2wNM0a1Z+UCrZvqgbXVWZhEVCqxvpiwrX
5lkFOHwLNLOzrLZxEnxhCd7XkzxiOXQm6bjmj6rZOMtT+LTC9W05QeFJl7P8cjLX1tfAF0KbxRqJ
BJJU8OSR9cNr0pv+CBZvFXFndGaih8jGTYsvFv2apzk9hlGuWA+T9fRTbnBrktnNkaswIPYcq2Im
ttmyEb7ySE3Jb4Mz0IiaskFwhpvk8eqjexbJXxUlQoB+8axkSReSz0R8A16Y5g+8AaggDC4OU+7Y
vHigKGqXomg/OkC4Mv5QG/lItMz6NfFalQ2tIWgo33hBVBhKydypRIC0Q1Q+moLAKDc45jQP13FN
rHUk6CX5+jpjsf9gJvV/nXZOoJWEB5mfL/eGNKCxxhMXzoDfvbqtxalU/FfsMZjeOmAo1e5d6RSv
12EBWEvAFGmz3uYkP7LEUgB93QxRA7DW+oMtx5Esro0zhZgYWHJer3JAV8LR1qxLBD6Onw4yJ/+J
S8zK06nMENKIjnH/+4gy1If4Z5+gl57gM1x1X7vHsNBh3CMNsII55qJ1FA8S5OkZSUjWMKOyrszl
Zm3rIsPrBTQfTNn3qYaw7t0cDojLFYwoNI6aD3YzVXlhGmrO8s+os5cdT+HvGYzORumFQMhnGNRh
QAreLZs2ZeeG/p7Q4pTY+rFuQL00oK4wYlqvG6BlUycWkUy8NC5UF6K9bQaZ0UCsp58jYRU7Ldbf
2QojMS/frBz+nW192o5ZRcKfozKzVgmz6wG1hn1IRCpR4HLLXwrE5HBpc27jP7QFL9BIBf0rQSon
r6YwHKXZLfqqO+Db5HVUSv2Zc73TZARNgMoob0lN/gX078GaCPViHWEG9jAe1Wf+liM54qIt7d4d
bNwP5UhW/wr4429BlMDXu4NTY+QulIN8gHOyiKpJv+wSLWMNH3C7rpedyM+poMku6PYZkACEB/K9
LcIp7zupUQunYTbYk68mIU/3ICmQ/1J01WmLmwcdpKSyr0h4aQrSjz68JteeK77TKMQ0Y6jImtU+
/iYtjPkvDBUiRAEYDkfAACRPhIYbUMRFWmbzFLccAsAMdheIH+P+zWtss3c1aH7uHObpgEZ6Tomy
8pv0HV9zeyy4FK26HD0e6845Wnr2hkj65oUpToLYf4Tu5r1cVcUR0As7vKf2rX6YA7KjTJQvvETC
zzEs9n8qndzAIMqBe/DhvUh/I7CZhBIONbWHNrbuZb+PvPleSQrUJaMAAnQxXeNn1jpEDu+gdVuX
IqMblkf8X4nbVPwsuKbelLSCOkuIoGgH33UHa89jRFgZ57CJ41zqibFr6Kcxn8+fhY4dIvvNnwYR
3Oo4vCjXo50eVfPX5n41gKUTMtxIsPjju43QMb8x82DTu1xjzJE30JsXCaDEjCzhf5QbPTunFmNN
LJE6KBnfrTuLYKT484GEBUmnI0hQYpYe3mKMPP3H71CeGIO/am+bqBszsoeZEELE0rt9sg3ZCWSZ
sYm1kRxw+Gdzt5TGb95pjIUP6kPpyTuMtkfHvXvrni5FNngvIQPbEFAvKZId9ioQOWREbcTy7Jz7
gS5F2+0bSm8RhRyUcLSDhTdZfWbGKBrY3oKPowXAxVz4ck3HcT3bHs0pSHwdJm2njatGJ3yopfF1
49b1kUgoZAMFnY812p5ZcXEG0tZmkUNSmV4uq69bP4KxaLttl4Ge5PLKdy9/MKeNlgnkGrcMJsX1
Rzf8a3oIK9N9YKrnqNbmSSdas1/vh9BWkhRwfJfFgB9bPSxETTCRlLP4QCa1mM1O7a6zB39dLgW8
qf1IF/xBVkLs5dKeyq5RqZbvu+PlK1t4TLJYW5xOQ0IHlfii1KLmilazZ4GAACnVerKbspCTWGyO
fx+yoGjhVrmfJENOfhsGt+wb5JW+4f0bw7ZHshjZJDjWUUNFinHbUd1SqyuJBxWFmtAgtHEKdcTb
069rkpjn8u5pgyuEpTQ7POcZWba4BGrg91qCSE/hBeRJYJQOtCkSo3hDfVwPdFfpxyijBJcaZoP3
adZknrqk4R3OXrRlaeFshkTdi0CEFwt7VDBO0ZZVmxFo2++jXBMaPy9OrINmTUnV8S+sYwC9EceF
pBUw3pNaMC/ZnrMflBkgH56IMqe7jaUZtVeXnqcEpBdBPAFQB1BJsZyikUmj08wRROg+OnlWn1Xg
xHVCcplXYbojhkXRch1RjUQyL75HcLVeJJdIJucuL7ukd1gWcac2BKqgaWYbyuoJUFY/VDeE/qZx
xLa2l/PlH5m7ezzJLmSFTvTyLf/7Ctl+E9xz3EtI6HBI+5iEZ3VcSzv9AUOIdN1Xu5dp21upBXJC
GOVAyKoe41QBH4vkn3g4eVhKoKS8R5KdNOOxX+N8a1/vYn2zEtjY7BdgSHDTMVZFz2FB8nBSYpZN
7rbLN6pRFPfHSOo7P9tTfelsCH2FnAilGnkDRdxEXM4IRMOP73mIDpr9FZnhWKMHvcnbrtPOimNq
2hoCiw/tM7TSujSLNHi+XyNLspOoMIywxyw741tCANouY55ZMsdWOmX+BgMzVIoemRqv+w+7zbYA
2ZQFHDMJ5o2rzCkv0cS0CEU9bBDGac2qfrkwE0oHcXzp0DXfHSvfx2XWsVXRbhh/RLZR3P8n87Tj
eJJLOVN6SZsk4VMDMkz4jumLxAUOdoxi1NoMMqebg1ttCsuTsqVxye9kepwE6yRUMH5ji6O9E02Y
XVnp1dprlXq/Repw3d3zcqQGJV/aQRjOj4JEo0KUq4TC2SxucPE0Pl0YWeqOjDs+lpDDxZ1T8K4e
3eV+ex4/EMX0zA2jKamAoc6AHTw/f7XgTNQ/neqnLmjvNWGLWyndnYGeYGS7Gyq9/b24PUE7NVZ7
u097qO7M4KHM3xZPgqkUXEtiRluVMcmLVYArr06URFLCVUvLBCR689qpBRAl8/6N6Kvhou/a/h/M
F3rBFflSa3OqnFAKTrfsjsFE06d/pg6MCIro+doWGnJNrgWUDxbBUlFbkwQozC+1Jv9mLTgc/IQ5
/6Ug1tVj5K7gF77d2t84r9aSbx/6QfqlsjQbJZCeHIFKcnflOLBi/NViXfWHLvWFcZEZIaxxFA4R
fIdpNwyQ3ePnd/86VQi5mPop7FH5JLhU0JnFqlFv5mqptWhwMJeIJicr0fl5yH7ASZ414p0/jXno
9GnlNDDm2LekbGuVsLA3c5ge7+5XDaKhORAFZh27uMVIQPe5jSAYyznXFxmr9QNUhWT73/1sHO+z
q9I2b2SmkfxKx678GHQs5v2bW7IurYjt/+UG7rr9Jv/oGhLyh7JA2hIaz2tFBwfzqagrkrMBDdfO
dxnnLuVmxYdE5NUDjMmMdlCvRLfozVy9yFN02zkjXasPQBskyZob0YOheeDYMFTrAsZvKDZ6PcJJ
Gfj7bKjxhkyLTo9VXdevxLUFQ/yu2YpJqNwaH4+dM4o1/5vVm0hKdOR15Z7p3VEdnW4K4nfTHlwM
khdy1zL3C2EulxSsEbiZ1OBpnZe9TzjANsmo54sAwQVk/6pAGff1WBxEKGrA6pvEXPZ2tebi9HLN
DdbyinDacrlT//4xqE6KTr8FFtVw5TmsktHDRlVVlwr22NW9PkH30aFj6UOndqrCE9/fC3bsAwv5
zqowC2UcUUVnugdduRijX2bTrjzKRdii3Fzj5ZBkuOth8gL3QncjoW58w4g863hYSnsL8n9wx0ET
+qB3GJ5SfbyZSsRKtrMthUEmLPfquXIucF9tSJW+ltqrVQBhnubZyNgYrFKfYYXa9AzI6qET9UYl
4FaDAGYVQKLPt1szuRefTsEOpGhN7O3l1HtVbWWOHGy7j4HzY+G2fW1ngHRL1IKn+zR87HsZKeaQ
FCgK8BqoDLstzSUxFr3DUEyeb854SZp73SOyXxabUBYkoALc6/x8WUoYgVHvZdvByOmP6Z91uBLK
7hSF+etzGmHFJikFmf9XL9miom6lTET6VhhtRFchzZBfFTe7XmvRQa8rRTTmirfTXxFIEs8iuzlj
UfI8eTLZxTesUo+v/CAjGUWEb+zN+kD/e27znnPVbCNLa2f9qg0WMk36wkrZKnnmEQycxRirEJKb
Wx3SdifUud+Q90OFX8v70gZknQ394uMafUqwh7tPrcx10vMBfo0pVN3bZ7WO3dNRqDVmUCKNX0n6
BnDqrYmWtHufcHCfsWSqXWUAfavcdhp7/CrcoLfC55IUZZTXpLa6lrY31CD6GP/hnrl2P6eA+5vJ
hd1X5SHL8XH354gEbXToO5xCHsatYlksjNw+vcMXuLs0wClvBaYOwZQ2mjdGEmjplXYdYwE/6kar
7272Vg/ArJTEe3iLeP1loG9mddzxlREVWTi/R6bQBE2S5BbVBqmNUyt9ps/VvJWgS4RmG+gO/hNs
nemlS2o1yOj0xDu0gas3SFyrOTgKcj7lGDDMDxrFwra8fn97K/R6WiWV8fSYGuNryteKWVb9091S
oXDGSdG/pAS4hEqCBP3Rrkh7ldVgoC5QIAYUC1bhXF4dqG4jAiUyD4twcFohXCkvO6ECryaIF6mX
53u0RqbpPyJRITt7N7u2LrtBZNwcsRX4fHNo6l6dEQb4A7GX60EjvWRRqWqmgAE9udir7WmnVBHW
it+Q86ZfB14aRsTKnGtfCGqO84HKhISKUKCt3mPJx0Jz4ugJOb6gaG33gJEwjdzBqSK+gxKPobwl
q4a4Wwi6FyouZ1yISJH/a0pxdcQkC3Z8ATIEyiuyLrdxqXJ69BdgDPdNIujWTmMnW9QTr7xBN6n3
CSpBxhAI6ih08kprwItw+sDCijuxePP1GOr+7AZo9dDqgp4d7Q2anD3TcN3TQF9Lk6ideglNgz6v
IqX9S/A8Nwbq+dFx46R5jrOC8naGh4J/3a086bKZ6nMZVQKU0Lc4DQgWxqtpzAVJYRmvRKvFASJh
/FCuFGM3L5bCcdyg4XfqzA9dN5F4WabcX8iKDMgmn1r/1i8JgIIxI8iDWGXMwxBpastG/DIIrzBB
Hp4YHZ9dircklGuqGrLj9d51GBNbmOAIh0By/eJIXU6qghgdISTTjCVxQsbQJ91jBR8kMaZO/kec
RGvl74hwZsKS23iIN5KrvhXYvQxXy6bh7xx9g6Rg4tL4OQ98f8xGoKSQdpXqRakVp58X2I7QdAJc
+E90m65Nh76HbbWzpV6eml4GBrlckiNNO2Q/bLsWXk8L9s2xZ5Xg498jQ0vEb5is12MZhQht4wxs
o31BYqt42I3ePy8aLWSKGl9K2BIY/arNb5bszWW9m2vqp+/4XoR0NxCc8+ldA44VpWRURTp3HeWX
oA25h4kHQXHXX1AnlmDp3wKBRwUJ2d8nk39rSZjk9h/upUZldw0EkLG89MQpPoYLzLGMmEkpVFk3
qKMs1SRI52pgsVE7262V6oPZaaoeK1MGtkxg73oJ7mHM2xGLWktBfNu94iDGXOcjzXb7hrsioU0g
MEjF7OZIJUL3VN+zSiiByBjfWEiOw7lAsIX/EeoSA9FO3BgkRi6mlzr+8tgATiLCR84Zu1H5clMA
SRm8/Nju2aP7Vs5ud7JIqN22hORtlzVSLxgFQDh62SFh7A2rXzpEhYpelD0/3W8YeBtjiSKEI1X/
iaeykRGN/MqSlSrtilRJIv63XeTTzhQUyEtWGM6wIIedpuUDCYAVTKPaCdZrk6Tk6+Faye8DOFt6
y/RfL4EECyoZcpsbHjuWrHgPcu5N/O4H2opmxgaLBoPAWazbsbyj5SQtCGmw8Wu9Z8dLecJWcIcg
AZFqUI7VrO/GRGHQkRjHVsiDscZ/i/NWzeHIKXHrk91oUJW/NcEJBpCA+FaMkCOqfIlsl5U9mpxy
ITUzF2IkLZFRvTUGUjZliXAJrGflJJJbGupazqOkEcXfrhP2TvNXfVj5/8fKRc0SqQL6kqh27ShM
ASeymQ52ZMsaTomx9SgekphCT8RNWpdJicZ4bHm64ii80sIaELhu7tZFz2zFMwaVhIsBPdA9U3jB
ToTk3GiSZLGpiZxshCKzZfvjzJ2U6Qdr0vdaY1hXeeV6Zadd3/8XaaXmJk1MpFa4kF4wH/FN2df1
mIFaDQyLK2nUwThHsZjBXj6sUtnd+pd3bIR8dR2fus5wqQWF3+tNjqCyElKW6ZEH4Z+YdH348viI
r1rV7YE0PUBF2PaOELj3EeeXFbaMYIY4q37X14ZjJSv8oH6L0ImUlW+V5Yd6YfgTjXb30JV6bXQx
5xtZHGrydC03pL512/xXN7ryJlcgrNTRtAKZPDMDO4lrW/jvFJzQEBqOaUtLCUMz/252KnVnkwiR
4GV+Sw1s3Kg+Tod6tvqLcbKs6qppt8pNGVv5U5m1f3ffEuQeVNrZUMEDDGvqr2sI/7s26piY7Er8
UtISSdexoXEDEJFDwgE/FMDwNw7WRKsLH6r6mCwysKvLz2LksX26o1Ryv50bAd89T/GjwgaTL1L9
b7fHcZ1Mvnvr8KMCFPX/doe2lDNKs7pMp/Ixda5L3/RLgDgAd7ryt1XAeBw2Dd/iRWkFmBpZe29o
8p4gkHKHyMW3LfVxsxKuaQQASfN9De1YohJeLorL3IVkdAxBWCacZC1XFI2KbTye7Ny7tXbIDLaL
np5zyN8zYfFjapCatH8+IaTJbdRfI6DIZAds++114EctogzpnSHFARXu8NjW00QQmEpfuRd+lCU0
8R7LV5xxTq9OJpZSKskgL4MksEz1m9dn4DZ3T9GlELGV3CCfvNp17HzEgmLlKXJ4XW8iJGEXWIW+
p9aHjz6nMmCN303NZpk+cb8TXgXi/YVBAFnM4qAYZ9vngBYLE3T2eIkI7Yq5jzotY1pZdNiTMu6D
qEy9z/d5NZ5Vf8D4i3FiQYwDuu1ikO/Ktm0p/mrtzkzEfxfisaajTmhpur0A7ERBQDexbdYBlzY3
Ljxi4V5IE92KkEDDnwU4DGnqFGccMXFjm0Ur6nHZBu0DZ3xu2bv1AMYBuy0ne+mo1IuYiWRSkxaJ
GUcO6jN6UcqSsCLjiXE0g8RZU3CnyWy8fr8ezR803zAQNBOAeMhjIuE5ElMtWC2GvrkrE4QU0nhw
gzJcgoZqYe5JpWku5TgzfelmxgZwZmS0+SaP05Pp7tW/Lvz+OUWpdyYLqDBKs1th9NHwYT0CgZ3u
Bs7q0lWywY76WT3+9wAMO7WKUMLqZBjSf2LiJOQRFLEUo+DAPLKpWo8Kn9dfxr55NKd1yl/PhAYB
15Er6mz4v80QCCiRerV/XIptMC2HlFuo/ohejVSx427GDvws7T/TBBTZnHiMIMUB6B36gwJs5H/n
Cf9XNqarX4M2+tmXsxShnZQnpnN0jyYcReXFZC4Rn+AJXvZl176webTzLZUe+kY4Qr8P+A0jB4GV
jx4xq70+Va8CNTUyemBEXp3hS40rM7xb+dV78AoXjPFV4m7LPycb811vPRCDTN/prdDtie8bUecO
AmCtlsE2N40qKNDVMpcOhuljgLQjrQr5GjMV2LLaxRbgadEgEg+3Dft1ILM9iH9/70+K9OOSD4HL
OMpc7Vllitb3WDgvMAxzEfOxDp8wctncCbp+ELRU0Q2RMNmEWYNLaeenZiU7b9r5hfWSYrnJP8Nv
nfBrzL+Pl1y/UgaU6Wcc7lGgfWutQzsr+K/slV7CnEm3sqFJv4PCjf+FQXQ4CvgBDzYVmuEwCazv
ZPGXauNv/G7MNjBzFRWwJfdvH9M08kz7tQ/n88t/eCHKSKO7aO/1qFhdUdAjm6Aoe5/cbNG6aD3V
KOAxsU4KLRXCjRXpo6iT5wJh3Bb4mv2Nse4lpJxHY+h3vzL8ePWOkWmLRpHkyvQhfI7ONRyctiDg
5dg+dasPhhZfRiNd+s34VkzqZsl4QPwhXWOq9XJrlkRDrsFaM3ADXQy3w+sfJaWSsv1FFLQBZEZ8
b9Py+HydjO0AqKygCzXUzSsN+tvntmRQc4V3H+InbCiR+/6JdVUSZOCYBPMml0LpeeA5AUhw1L22
EQpLcRTl1tOQ9VpZunrHsbauytZyoVfxoKQjC5wMY1IGcu04QwO9Eydd5XRYraQbhpZ37Q6JvYX4
EpHfEl4rPY7kTsH1qoFDvTG53cNFLFW0JRu9khGC+s5IDjFIFRXFl9/5odP57TMFuepbP887y3WE
PTJRWlSj0XyrVjaJICgvwHWhDPtcfP3g9QJijSaoxAyJDleaaolQbAfcGxl5eXu+GiK9v1PCKemQ
o5mCVmI/EN2RT4eQoBy5aRDKy4xJNg2ZtUzUA13PDvb3hE7LztiAIqwGC/10iHf+55rN0NchvHIJ
JQTm4ocOeBBjQF9z4klRs4oGn2mGo9W6+amxbsvVSBSga/kUp9PE2K9n5pjJQDD93b8WbGMyRh78
GOLz8+4kZzcAse8dZCHaOsejjQyWX6sxkZ1ykQStOncIXpRIGbtE6Syz+PjtOhVvab3mHKvoLpCY
u7rN141vstU5dF/KvhwH3KHNS0UJZse/sf09VKy6Pw7OpNGvsRpxzTT7aTRYuYvYvA2fTNC01DQk
Vct9CFxJxngnKWZ1spHe4Dp3a7GmE2PB6/UQUXApoHu+8J4UAmb6xpK0TFgESxJr7MXtcjGYLWfq
aqbd4Swx6jfb8HDbYhkpeqBzO5gK2i0jIepG47bFFRl0pzEXoGnfz9KO7+PYD6gs6TEdVTmpqIRP
BdMMNegqhDu6Bi3MxZHPyUO/0q503AZlSUoawEmh/rubHfpb9QwWdfrlItXc8vC9o0FDLvxqCktj
Dp4ceYThdCroNXWHiRwmvbX3THdp2rIOcGxkPIFcNIRrE5faCqXsV3lVF2tZjzrVFQ67lo1GSJd3
96q7X0RsaP++F1+q3QIwDuv2UeLRA0f6C4vp2rGaYQvN6UVCElNn/nDyuRZIIWYFS2KN3/KGRy56
j1ZQcu33JK0BcxZ+1bUrBgPrBUvwAlr1Af6tFdGSXpV7PWX16XP3PSQUJQD50Ydw/brhSeNginL4
DxvWsAYclN/CbdDq9OPyaWFz0oF4n7wPhSr74OPk1xwn//5fmn77iEKqy68BEqRg53YrNC/Uhwtr
q+Cq63/hNzzcfwrCGAryrAnSyV2upVa8h1vUG2uJzDGRMn26/Xrjv+EGEOQ1hWmttAsk28XrtdE9
k4QldCjiOaFtAoUh+ihU4nwAEw+LPkRb3Mw1UW06tMlsXbXXBN1nJsyao/jg/vfM/TtfMDLYLFf+
HQQIjNpJJVQ6taYrc4UVtJXEvqj5SaeDf/cTlyi/K66b4PMEODNzG1Ji5hhT2DZHQ3wuG1rw9Vfq
xV9PRZ/j2ti6DlIBYlXSLjgGP2C2UszAk2WQtbNsYZdhh2dYhjTm5pa3Y3/T5Rb9yWI5BlwTzRuW
tZvDjdLkIOSaLriYRWGkuOeWDM77zzHaxBoJcBjXrnEKakstey8wAHkA6oVIYZEVpTpMO9yCEFYR
34gHQvxBDwV1pQYOo3YuPhTdbRJshDQA8fCahM24RHPMaVxJVgSGsOnumf7kDNX90zU8Sx/y9Apm
GDSFV2ogkFa3fgW5BiqKn/6jWilAyeS+Qsu2EwzNyZ6NVn8dwkcoMSJL06ZmP59jGw4Nued0p+FV
VdDogNsd5YNiWegpbLLUhEqd0gm9z8/mUgRt6rSePWmmHerX0oqOGUhwutKHCNAoFpep9l+Ka/XH
zVfM70xVWSd4INn8xJ6zzDf6bxSkwy26WrHNk9lFKTwtFxkyL476iXDvVaf7+82RpK+zLMTwulnK
AstxePnoGDhtCOKhJ7e740X6Jxzu/zkeGfMBKYG3ahCjH4cRzTuLDEuEr8bHU/TwPM5fQeKj+uYl
Re4na/gCWAk2Dj7PaM58vA3HuAj+pfZXkcguc7cxLkffNVK/9box6nC1zNAPB2ydNIB6DJsMTil1
nD7QpmRiudgLTp+4CDppuX6InN5JTovInPz6/ZLejRc0vIbMl43Ehi/iCENwQjkBQYChqhM2/J7d
VO0LMrYNRcJyqbrl9YNh6qiFr0YrzjYTs7T3pNb3hEH0RjpPie88S27QAzdkY76QGeke4wKzxQWa
HPS5XHBYQYVW3Bje68IIT/fAmBfR7IDQJRMGYf7h0dKzERJYXpMi0xHpdW1dD2PaGjSlasSr5sCF
2Jne3wk7KhoelCzslskCiIIF3iTL3yob2iRyS03xfoLN/NRV6lwikP7g2z8RQQGurxmgrCD6fRX2
B+bIrukA1ObNd0HJf6HGRxkaxoyu8Dpwgctn6jKXhljwi4BqicWgwPFE7D88dBqjys3QBWjhReBF
M/fTVoFoSBTVD1Ui2koUg5yT7oPP74/6KbenaTjjqN1fOScflYrQ0+JKofZg81jKoxZzG+QxZXKG
ScIgGgzbkjzeQqs8amDc8jxhd2eCqpeRIr3hrwMvzIn58qAr7YTqPss84cimkl6ReuLjmsQj4jjm
EPnSF0tQ7djESQxbspqwi7qTiAXDvAgXW3McUoFJqhelelcUATahxG5UK3oy5jX5zyDa1gif6nWE
hKoyLMkvBURHHCUpZOQ/8dBAWXPY4mhU6h7lt/O0y8q+o6YJPl0/jYOZJsW1PYDav5Mp/MBZ0pk+
ZmeC/mwZ+uSEukrqhe5WzxjTYAy1imkDku2m3VvwRbLzcWjTkn+wdimALx5qR3p33pTPYGLcnKg7
bkZsvQcQbVJRUlxi1zFQStnS2uzfTuGQckTeLNi4sAsOHwTft25d85PdgAXcKzborGb8iVquFcZs
JQdpXGuBTOlLWdBME595uV+PKuh+KoZOjU415eRdj2p46GjA7Mumwlu8IaTWN8AHo+JhSsTcG0Mb
gSSqasZWeMxfH8eA2pf2dOb5dhroJCM+jhW/6qph98yt/Khi1K1/8kXODmYu15o3hMEFkYC6QYFI
XNxwQgCeYsZJSU3QrqzM5NPChe79Kuma3tJvf9wBAmFUbq+VHO0O+0t/qOoYO71p/+LgFFmpLlhD
LSXe3ayidV5Dud4H9LJXmcvDmBOfnPNJpkGUSTy+nY3ekFgwYX1NKrVieEpCbpNKhEu4lsrcExkh
8aHrcCSmbDVME7RH1LAQlYgkfpuhQXQ3qsdrrDZ/bbaSByjaW/hV73I4SkX2F0lsym69SSLRetUx
qTDjEO646t3KjetAnCkZgxRgTnvpGe3nDKcCleDUUxbT1WV5wLoa+HuZ4mpGF9EHja9veVNhJYB+
0+qy0AsshO/dmzsZ+B7PiWK17Hbm0AQg64vPRo8lKD4Z+Ebav/3gppURUiEkTxtjxtO43BDRr9mZ
gSrXRtroQWZ+WYZsuqw9yGmHJ/RzjbXTn1S2KJXeiShkRpxOljFHlHMBasFLSu9JMmT0znbNIM/a
5IqDYmZnRScZBO+rh9eSX9g6YccuIo4Vh2nIznH+tJbyWYldJ8GhSVo2Mty7dq4/Y/GLILdrsMyi
JnKM3pU/suUUfOu3KupDM9R2lPus0d63R0F5mreE59ius1Q76Hrd+MzpxkwtkBcqSy3O7bAFiGjW
w1AtZtdl3kvbseLPtKr+L3caRYdReqGNO/BGBIw4D9re+uC8SmwyOB0yFb2+jf2ziASX3AT9OEmj
7cvXf6VrpOL2qG44rottjDAPIVya4/vV9tdvpzMs4N13SMOmDXvjCIb1+NR0QCE8kh+TcrwzYYer
bWj+dYCwWrKr4V2X7T1efVZqbCxFBYFB+XnMHCzCHobD5S65eiSa1P9zluuG6N4JtCW2fixUfnzp
QGUXSWrH3aa25TDFB5EOjgASWyJaU/GsjKjF95+VlpLm8YvrOBEZAnTtfjh7bUDIby4WCGTAROoG
HLZyZo0AU9aVK6UsZ2l51mGxiJHWapSGwy8woTWq5hLsqNahZ27sfhyoihy6oD+OF8Wxu+WI0fgb
toQs59cZ0VBDPiL0FJx6IGEUi/u5ftFz7cKxfrm+Ko2LJQ9FWyLT+9tPCtB63U+7DDUzATEigOcj
6erFP/7Op0fybKVkkioi6XJS7thi7t+ENlOe3pCx2YfnqD98G+KfY1RoYxpG8bZfsG0+KFGXBCLl
JvIkHfHqbUgYeBGx65qZIDn4hSaWJWiNEdh6EG3sOS/7M8N3c2QQ4Ml1/35WM9CCTi8J8vYSI4Es
k0tY7n08HmFtpUyyHiUEwmd9/Poq/1PgdGZLanwrtrnRhnd4TvkFqtECTaF5BY3hjnZi2xhpHCNl
eCWwldupsVcmnbkf82JsNg8ZRdZUFGRF3HdrUYnm6oG4P3bVBcv7HByP7WBr8QhfzWLsmTC3uakA
2fgnnPBG/AtoyxJbG16PfeuKf7m9uLBL/lMVEZpRBPJG2jsDuEzI6gFj8UpAqOHfI+zy703D8WkH
vGbuqnYFpizR3uIUed6HZ1j2JTgcwKwhzYfBA0lpuFwmEb4Y+v2JgcSagmC9mxCkyHLZz0AiaqRD
jU4McevMkNhxTTsVuXp9gzTZwlRga86l17MQsrfuQQ8cPVwTI63OoMcClnXc6wQQxv+13PNbxlJD
WBv8YiYAmCV+A76fBPaPUTCaNFEcVOsbj7wmT8tKRcJa3mQ/gjzTFRDhOkBsHAmz/Oa1/7su9jED
L9+W3lN4TLlPcVbX6tXmF/9DmG5XQwlrYRfz9q87tzzhF8WzlT3SpY796L1pR7AqjcGCGdCAFGII
bstGdggkmWJ/pKp4V+LGHILGZqI0dsZFMAMFTYGaMXNT3gGr4QgOye94fnIEMUiSSO2Q37SCixBc
XtzVMwIhYFayrr6vuTjNpy4CJATGmNGNwpdChy2/Qas4+LXBw6mdSHc//vR5NVsPjBH46n0v5bwP
0JlYj2SlQ1t3EKXpWlHIEM4pYFnwYqqLk5ZMNsqnakSV7UejfIVMNiJ1KijnKHZx9+q56uJmYvYL
3wBmknKzd035xQXxwa4B45vehws2uFpvuD5NmBcFu8Yov2A/RKm7lUNxvPmKGanB9Btx/ejYdloF
y8A/BHXKCuEjdzrqui5sQD6B9QhynbRfkTykrdEBF66RTv+tKtSyCwqn8lzo+mdmP+X89XoKaan7
+SNWMpH7Uvqpf+yXj9znwliXDMdQ0Mt7S1/yHTC/B4twQATK4mJS6BPNpgt6RptS7Itzjsg2XJHA
KYmruEc+JukqbhDw9PPoau+MCTIqwp2dypg8pZEZ+1iuXepRTZDVpBHA+88fsfliV+6G+OhB6Fbq
IDXbfj19hWFnswJX2F8aGl7GD/5eWUcYbu1eCKjew7ofNilCq0bSRKexWHvvpt5rMHEpGuLCU+pH
OmmaOoq4mpeW2iz8Ca+dtDw82Fne7bpbUja3I+VUxC4CxDF0SULbdtjwyzBKJgx7hTDKOnPsgQiG
46i5XWEiUHsbJJKjlGiasGW+3GdLvKgARQ/xTeuGFykcpMiC9e/ng+fiWFoGRfNYKbMa4F3Ps/UK
SVcjQknxb5iwMXcqZGapjS2XyrKTc60n24BjdlGFnU51ZmorwytFZejEsYw6+ZpSCTHhqS0CxX2E
uLC7ybiQN6v9qwQrI92kdb8k/dRsCbp2ZLx5axfI8bBcd8I6d21/b7ydTMAk5To1Ii2iY2MJQRh2
fPHDr7IAsAqx9ZzxytW9sqXXe/qbSiITr1lGIz0mrf5G35uMhl1d1Zq36DnvIMrF3NVQGjvrides
j4yJIn6QjXpfJEpR2ZjTi9GarBVe4audMLxk3fAYcrEc18mupS+txD8xSSMW6sZ4WlNIlCho0v48
Sv3FhR2wDf0w8y/fBKulH6cUqu/A5wjO3qRT6LRrh4ACEedGnWkS9E5SYQZ3ipcewmOjh8Ur1fla
qNulP4xXAgkyMDBZoy/iXYf5pvTrT4174u0hSPu7XLYRKoDxDaYfv1QX3b8YXkmTE/x14dPAtmA+
bKQH3QyPf6TuRKVwcBAyATeLIVgtw0guAwbKwQIkuqgHsbtpqR1ZJVmNDwLhmz6G0pEQCj188icR
5En0+SKhruwxejN4HR0TSNYy34xumm4lXOLbzfvdqaPZ0F+kJuYvxPyCET7I0cch/K7YhrKf+rUr
M2RQDan1kYhiGBvgiVH8cHaC7n7G61iQ0Q2/04yc7c+U4te1ByxgTpfVIDIy3Rxm90qdxcF0OVi9
F0zQHZnD5zkbGwPK2QVtFwdSUtvEwwsFz57xnOWT3m4Ti1/CtltKfHBp0A6SD9dp+NcwB6opXggh
zGfIQaZu8W095qO7cpgr1ZNrgAKeKf/3BA9DDXYVcc/FSYkaSf3IUYqR3EdpubbpvgtW18ydUg6c
AjPLhBn3ic0NBgXTKHa5jEh2C2d7w4uuWvhhXKOcRVz3a58ESXHqY+SEDLBigsLIkgQfuamhfPH2
iHgfozUJdaXkbnX1V1R/CsW3lDA2HCe4S+Aw9cXPIzjJmamvg2qc9rVuwT8EVMegKP4YHNZsj7Qk
Cs9rNBrVbTAKgM5rcjgHbBau/s2znG/SJ8YzER9iwIBkyEqdypuIVty/Mm/UX5v41p6R0gCzHO5e
T/ZMeVAAfILZMqxOPfb3heVFuvlJBrzknmoEr/dzCBlTF9I+hq1S+53DHwSru/E00lVGjy54RvQA
ScwFZX/6C9jm3fd1YG0gTzNeh/sLWyhNTVSktQFE43EHbaDRrNU398CcNJWpP0onIK6HCW4JZZdt
lUcyhgoDCV+o9EfMtbASg8Mr7+XtuyZnDv4svrvW6uJdzmoXAvCfHwpMhyiCt2n72ofQbRZQqZ/8
8pgJfEukw65/95MwHVv2NEtmpIMBw6OJVTctoizB+/KlTp8uGas6IlUqzZw6W2Nv/2JmI6nPl4CG
Kl0sxaFeCVCjMk11kQm1IFBP+SL/IW3yb9VBrF9gX1TUr/LtZjTySRp4kRL9PzkMMZnjgoMbaIK6
hWwOh5bgV00bJ0DxIVWWsOY5auDJdYgVusuCjHgXW/gljFZDBH3K9KJejB26KI3kTHG5taTRUKA2
qo5Gu+1HE/zVu6L9zkrRgf+/WsoDNFh73topLwhWL1x0ItqOVUxLmuivIDMDJsIw3g7E9bvDsX+l
+CC+JcOqIXYZdriTEDXUOp618dj3aJiVNq4EBHFbwXZsZOUAENXImlBUiHDmZQP9Mos95aH4/Mj/
Mxff9Nn9GLejDPcRziHnBPA09L4ZDdc5JWJe47chvxuNMcs14rwwBGsIByR8ALtm1pj4Yl2u+x5Q
voYOM2eee0DPI5g4xcqnW0q3Z0aJyUWrdzSBh09fHpzCLSu49tYoG7YcySnOHcYwctRWa9U+uNXV
LgGuoznYVXkFrS9ssLzwfJob9FTAlaAupZQjT3ilTnxpAh1QjUaoxSjUMG90ghRiT5x2jlg0prZT
/aAzeI1xLKHEB3jTDXAwaIh9O2G5ndW/H0AR5lKYX9wsmCrmKR/e8dxwCXck60mX/78JAsUSsfEh
MV8J3insEFEnhEY3K1yH9p7Blyen835eYJDlK7YKlHx4W36c59i9C2l1pZ/8VgyoYJ2xPr9fnEv6
oQ1hWWz3quyhSKNLC1EKUppPHLYfYw31e2NAYS8xqy87vfNsCUoOO3iZJ0ATmIOv2q1qOMy4CBDC
kSKjzzf8xzoCYsvZbQ6fbfyuRSyy+WsFbIM9FA5TNkXlvHFMh8XcXlOgq3wxInxHuRF0rDmmpH58
phVD1kdS471tAmlgqAyTnsMyrA4p2DQBE34UnDxdYq/d4UdDn+CoD8443FKksc9X0xt1PiwjUvj4
2nIip9TKK7Zo/mGNrFrbizUYfmeOKDelRXANkBMfoFUm8yWSRTro/iIbpFzDR3e6GiBM0pGzO8zN
algYq0urQ5gvynD0w8ku74jRKxdV5H+UE4Gr1MLX9hv2mABoIc7tB7X1krd7BRoLgkaCowdWcwHC
NPBlwsDbc6KLExaSCwLFsBGEPnFPkegrfN0v5gckb+f794osF2umQPbHh/TzkZUWzFkZHry2ykHg
er59kB8SDSLeAbLJwNxH4UnoM+72I1oIvTY/gOz3nk+R/uVO0N5wv20orE1Jua6lPcx1W0y3blXa
4PSbb7sOIa6tLcYjZev5i/nqdvT46o0+5j8MCwbJjDeslEuuBWMibKLJfVbxJ9z1Or0YqwTopUd0
tZ1G0VrrtoCBjyI6NcIe/16Yu8Copg8xmfiNFaofbkIwcVYFJm2LdeDg8T9im/BSuUY22pLyNiqj
W0pXU4Vt6+RnyuXIXiKR5IhHdPSqkxl61W/eNwkLPMTwP8Wdvydn0CrTYn1tR6W6XITACCBZBik+
Y2OG9QjU/6ri6lxnTCe0CJHwKI+3a5FqDmKz0spobx7Jts3n6GOe+hC0u5NkjMNkqfA1LtJ6+ez3
Zm6XOArudoNOfpKsbYe9l50ujDRlE/hl7MXzmjx3ArbTOXNgBGiem7XNSP3M9WMI8/nyVGKA1mTo
3wi/wt/KTgCMyHFxHj9SBLEGhg8GHgLkGseQSzgJ1p32A2e7nGIXfzE9UCdXYjnvaZgEhi94xjBX
WWzh/RJAzWuKPRpmiHG59oknDAT0/Iq3w9H9nqsdCL3J9htvz13jdPgwHFhZHtaIwTdM3AKNzTgm
vSCuTJVxdL//sJ5+7Rc+JALzuYZV2nIOw+sc6MtdvY0I9cIbbhELHGh5iWEW3nxdqGEOpupOpOtc
GYRgs1nUlFhk0Rxkkjmgxwy5HOWXScgqbIJhTOTcOz/PL8xKeXn0UWWme39pCYqgq/ZsIYVyahhl
HMwVcJzbvzTubx+vdCbG1+UsgWZ+e1P554HZrId4mfEf7E8tYeWyD7VjXvJE2ISOHgJil6BoTc84
dyKNp/mSwq9fQuO3aWIqrQDDXkVpvoxh5xLAuremVb5x93JQAE54KANUgVPZx0uqJ1AXEFGNDTPE
kM3AeI4jLN6uCaJR6j4o0iFVmFpSo97osTknbSorC4wLEW/wYNs4mEHS2/kYEpq43Zj+1zuS+UVU
8Qrk2CVP4ZEkZVtSoJxCIWSLfOHjSJnRybOfN4cUk298Rua68xi5Ur0IBDM9vdEr4TylPbVdvoeY
0ZKJi5ceWbyDg9BnPNSbvhrENPAJzmk3+wkQGOvsqvMe0QahRN1Jlu0p7O6YiFAq4bYop21PNA4/
fpOvbqcG7D4hFmdyMYzl/j5fyrO5OzHhrfpaJr5KiWgAnWJqOXXGcrttWVWCDfrlJty59iQfje9A
bLX1h4x+g2vY9GnhrAxO9d1dvjy1U90N1Ymwv4LCk34znUHAEBXD6IcAeQxQDXQg0lAE9aRTijXQ
bJwsXvw4UmC3Ek8i5bVNZq0u0Arlns+onwbKKWduEKZ6Bv1QupQng45SW3I40DbVVLez/5vsrsSh
oGe4K1fwgzLTU03KG5Yyu1gRK5+rVTl33o0d2aCpVQqXm0KkRFLG6x804UBNm4oktW9jWalq/p3H
SUDQLc02AtNO8UpeCpYdswoVT86SRRYOqoBiJbWvoHI1Km3Pwa2qnZfRbWr45/Oj0WEJ5zebuUaJ
CgNXJtjfVLmmWF6emmcFb5h6QxzQZ2pGUJIWRHMZWu0OrUKzOx/Acxq9Z+JjW+aUaGJFtfTtT91P
v7AsZ3UlRJrnlVT0MZvMO1v4Gs9W9untdcZBgLZ+ft0iOtstHGhXsmsQrqnCBlnjDDQSN/RauSTS
CPYoZ5u/PHAZBEmU7hEmon58euf/X21jxk/2GDT6q8gUXBFCpWL+U/rIYBs35GjgJTm4MvYQjOHU
wFS2HwQfc7ekJLhLWstiBRzNISm0E6lPmOVT0Iuq9IFY9plgBtrdUpLZTbj8VdtFReGBYn3KdsAq
5hToHkD3atpb+9jCgANvrtxIAdyLdnvFteCLZ8cyKdUMwgifQDvX6VPxH1uI7ZeNbR+JBWexMJyS
YMnPq70lUczf+3jeeF79J6kSy5Ec+O+X3hdwGXNogv+rkVpqdToM8eHZPqqG+eD5FX9/bQ5O2EbS
jkkk39oCVCJOj+COcAIL626Rm+wOn0eShQ58nGcEKR0ytNPz62RDy3QeXgqHe/pfYJZS/OE4a1L7
s5zl+xSb2gwgehKGu09jLynNWI2UqunQsNlEEXKGNesAwU/H5uzHIbNHKIyVkSU7s0ZdNPrtAi45
9d8JcxuHX95cMVNf+HJrSJOa4v+tOLF4+o2tAa/vBFfJJKH6s+xpFeG9ThS5nEjfKly2HJfg1lsB
1jm2JyduqK9E2KqaIUZvVTzeXS5wmr8kdruGMNAmxCtUW8xR75i9cg97apmu77D1yto9c2fCT5CE
YmlefChMXJzsEazY8FXA4T5+naLl/y+Ywf5Imra/07wdnkbNUrfZRvNhZZvO9iM5TpBNu9ahHjGJ
uS5OchvYxfuqG9W9rzpOk8W5jT7lwKhz8bacQEMI63b6JQP3GSOFx5Beor9filitoDppoiJ/jIOW
OhMTwVXeZUN04NDIZN9kH140i+ga2P2/7bFvADDwRuzh0Z04RyA01hxOavup8+5ZAn/8MIGpRbwX
PVMza/s0rTbs4uy/hQIdGyNuYn8qUoCwW15gy1ck9qhjV8IuwtlBV5T1ofX1/uTZDUPYMTZT3jq+
pQpru3dcCFsdwSLzUyMWUWOMS8lU+lzMu301PhWYuG/4150rREvJCrPVmv4myvhTAY/NK2zlf39w
RnABNLPfymMw2xPuBTHK7G2IeLJiSfoEI9zkJ43GwNDW+CSByktHtPZUx093lCV458+NJyZPVrR9
Jh1BY+HDoBnf5MzTBt8uSuiOaQJfTPPKNgpql/ND/4AqVXIqVJ8RUGyoZFnkZY0L2Zqs8W7Eq0sg
pkHeu6bVduq9K4xQwo6eD2CaH06pEmlHbtrW3N+NmWzvCwDBWmRJxQsNmIs6s3R7hgq/ESqcDq1c
GmdbJ5Z+gCkSonoq5LxeK1uws05vjfRPltgK/l2m/xudQrOQrYQcI0xZiKM2cvoa0yNX6VaAHIIx
LVPbUcv/32DNaDRBG+dnHrj/tpgduEoqlqN5lNeI3W8hklI52xqjxdHNB7sHP585ObOhEDVaq9q4
wHrZJ1llx6yEWM2ttZ4WnDazm2Z22BesuTkAWeoa12aE045c/FBmjdWnPzgBad4u2SAec1WrpLPt
B5qUhl8H4um2sVn+ND9zRbaZiO2zMrIGV0lTvRsmpQFHogZGlyhqc80UkPoBiAwBoXkndeS2zNnG
CNY+BCJbchV1EMATu3NDebC/lRMNPfhALPa7+V2Kpk7yO+7sM8b2Mn5IPO0ZewbqVgUHetmO8oQh
gePcC3cd4mxP1MeP+R6ypZPnRbrP/IICwzVjM7Gt5Grdfm2Ew8EUXWI54NI/WQ513VK162hm20ij
lXZN/fKTuKcyQDwawVBZDaMEe11riTM2QpnFasISjiLQrkdxj2GpPhFTfhd0GWwzuA3hBB8xMLie
6QOpEYFbeZPuiKvXK8388mwYim4DuSd0/pYBDvAGPl/BWcDLTG2SkvCJpIzuDQN3YyILlApBFo2K
587AgB97dhjEcPMfYeQTzvTbc9800yBQ1oiiO57mQP3bX1yFojukkC2J7wT1ZCa+SSh4jXXo6xj4
M/bGaTn22zFjH0ETBFFQ3yn4Oa9JofhDB+7+Kfld1VyVChjUktlmB361cDWAjhrGdzGo8hB5+ugr
WfuoKHIFfxPmBMTwkG2Wk60TJAhCuzxBNOMWyT51Zgqec9BLaxGvTM2+GPW8t0ZnLTFTKmbvgWQt
JIASqrfwmluiRcJlQve+A8izfU1pG5/X3nBXSnif0Rvcb+uOg1725JvCkawesFJ3JyQte2UUkEVb
eka2gYPCx2l91UT2NbrExEq+IJirc1Fli5j2Ow3A7kHDCN6fk3aS03t5Bux/3sBJY5ANSwrX/0JY
oVAXuzOSUw0xUMxwgNivF+/bocKA4tXnwAu/eqiPHbuEMxDzIE9PPbNER9eIAJe/tCicpo7A9Av9
/pfVJ/IkQJy7RDKtbM7QiODMK7424dF+dwYhO4wvcx5YtLPL7QLyKnuOM/cWbLw/Um/d8k9rHKrO
FTJmn6fpR0mzjDO1cwglu57mO+x9px0ZHt93TnHTRzP9t4588ouQ61NYDp0V9s06HzR370aJJHFS
/EX4azElN2pLknb7s1ZAMaW7BL8n8/Pi+wq16W85DllTBYb6FAGkplgTm1inj8aqly+qLrTPZxZz
cOu2CC4Nw4ivNyvh27Vhc9zIwm2AEb3od/9Uw+21gmux5kkClHV9iuWOQHhOl6Kt+NDcPd7BoD4q
v39HGpwbw4V6mW8qw6bTwPTYWojTvPHO1W8o5n3H3bvOCVLsWksQiGoJArB4nLeztYf/jMpLLulS
yqXa80Bx1QJL0HbLecasH0aqAZfnqRZYeVBpktWg20+06npI3xtCbHMmtkhLOTmcB9Ki6Rp1ztCi
oPwMjPvTKsqwWAi7hvTDHEk7i16UnhWxXuX0vi0fXv5Zcbg4YzGFUgxjG5PCStmaJZTEosL8tf9n
TE2t37E7Oh16it+BH711GbENLW/xaRZ/YV4lcs5oVbSVawBUM5PKolCokouevcdAQBCrTaI+yXQU
KUrqjtQ089S6ufdcKSfZgls3UGAwwhop5o3XoB75IGvpaBq+u3eHRrT3qX9Df/Smaft4WIU/ssm6
Bra80KmYjt4VGG1zNcCEnD2TBO5pwCgANJe8WPJMHp290lTA1o1/j1H40Uj/9UJ9G1tql1ia5VHi
fwlybtYE2TvdZBhwKZsys7UqzEpJ/z8Xe+NKFwqydskyv+l+UKM4m9RS2dqsLniF7d/+rGOmwpDJ
EhIycgX7yMO6CmetP9eE73mYqx5o4W/mBTJqGttPwBGCVCC2zlmgdGgbGGmQpIKgYbchhh6Qc7oC
5uJJvBEMjs+2hvN52NHWncyPGh1Q98QDNPWQmuI7gcLEmws0FZzcP354KMs5PyTrG8MiHXgWME30
HeKnqqM+xq0No4mMkf1ohGH/ROMo+U14rflj6lZ0zf9KzcovT1YjG1M70UaNU9F+Da6+4wiVfvAi
5+fQBUBBWIOZurQRFcJghygOk/izba+GFCzi53Rt8BVNHOEqwTsbELOy8rS5M2KRiDS5D8ZNwDMu
FEB2apLb9RsYLtVvkU8SRNxyQ1MfH4fLNLwTcXdhoRjKxbMovCq0+gGtY6qGzIGnXekd+kEcgl7T
pGjXp/YfY2r1wlTHJ82/gv435AiWiOVgLLksiYOOrB7rZ8UvqDnIOdZwcgw3suhwB/UdxuFFEqc9
3/bS/cwsjh9OXU+OZw4qJluWRXeCv2pqHQXflvLkxFcfdVAtiKgwtgEHUETYnx5DtlxTUsUnuNlI
F+Yt+3mTQn1dnFnJ0EWsoZ0u49eblU02Z0zk/9TYmuGWhIE+nsAPfuKTYmmzOzFExF+vB2LpV8Dc
zuvOU2QCEqZYMOH8s6bhoiia4qJJ2/ydZX4afD+rv5xOOTUA63L43zPnu7kCo1M07fPfd0BWl+YD
b+aCeSFODSxYdUO2A89HTySOzl4YssVrH3eVMe7JqB2fEexypAGAnD+aLxOfnl/vBNuBiFLKpl2f
isK+wc9Y843TpkF9hs+6uWXzyXjMEwidRCkQspZKI0kcLki/jdOfom8yg8a137Zv1m+xpohdXUoO
jNRAdnPdVJvtm3e7q9TJdfBNqaD02W5wA6LlL96E195GRMI1v1CosAxCdGMmvEqd9fSk49/6noAH
4bcE4sGOwW25IUGJBrZL3pzLy4in4q7jm2+DsAxoZShBKl+ngrpQXEsO8hVfHySPdeHvcrRC9viL
i3pXZCBku4DggbasAAk+A97/de29Zw3aGLnUr24snDYezBJwZvMczVsdlBn2t7UEDRkT3KezH3gL
CcHJdLUgQ7SexzoIya01KSyjuqtzP/RLfxcqv/DoTRxrWIMK/AV0o8voI/LvD6BCHJH7FTd7VnMf
5PrlRhQxQhKGURuSBzjyYAgGZta616lBJ+fCO4EnAbY2DDcXrjfy3ACMIK7on2w1fFs69aIOHGMu
cf5giDeIHnvD6ipyCaTYbnOQJ2uTsih1fHU2+JwKddn6tm5b1GENfVO+c0utwmWUFilz3d1ixWq+
6Rmu4uxHclzZ8PmPBlyNBElDfSRSOpkp4MwCRLwMi1hw3qr6wvk4n5/coW7JKnRf1jLlO2CLfPY+
9z2XwE+0Sizj39txh2uU1P8tybxDSjQt5lg6XzLa/LJK62eZJ19pqx5uhIv5CLS9Itp+IWufIYCy
2J1zeXPdW6kGBAmxF1R9CLmMIkpghn4u2vwgSwnJgef/qTXLdx5mdy4Sw/RffO7HdwVQUtaVyXYT
nMkDA4D8exAWvg+ArqruoBolELuqq8PW1onxfkFPVI0vRAwiLez4H5Iq0bhSvy1u6E6bmahdVU5j
a749vN3ynhdOogFuYNdC5mDErBZLBuEpwJSObrDws1ewqcq1k8Whi3Grh1POlHk5NO/6vm0ZY3xh
09fmtSlD6lLKiqLAURZT1qADFyJIjzREOmDA3wYWIz58nK9LFlTuBUy4eUNQsSeyArcJjCK3Uc0m
L03a0TN4Cj0AxV1HeqnY9tD5zWNB/OjQ4wEWeJlN6gzIjDiF9oxyK7YL2t3XfH1QMAMNAMreKpne
Pex4rT192kg+1WNMyGdUL/SJ0row0okEIPAxw6vOpNGR8y2EL6fxN4c2MpVhCORL2/DUxl8p98hu
hcZrCFzPWQkJqMtvwmQcSVHSaIJsmDdT/L6+klF+AuE3sXlYtRW7a17v81tSZwkq6stfwcHu9jr5
yAZnA0maqXR/10u/QlLSlSNqFYaDQqIBct+FDUs7BHf00j2VePZKojaj4vIuudQ9eMNfAyGeElr/
K3GtAVtRcOdujRIhQlvWElP6Ly4tMfMFooJP1XtIdmQaPAaN+FpOfTWc04+1ibSBs9e9sDbcDXfA
svmAWWU/P4Ry1Us6lG7V6w7/JpYqsHDHfPP3E/7aAkDQ3cf+qjpsUj+mMDrgytjYQRIcI2sHZ6W+
Nv2zrWMV31SefZrQrSVr93BNMEHWU9W1y2vjiGKulJmncm8ExWY6GuZ2AAAh27XczV+9QkLQU2vT
eekDBanVxPliwk0A3dptXyYLggrpwh2F39yfwFqreX5l0QfEGAZ9APJhOQH0gWBRq3kJtZLvuPas
Iw+ZnXU6gFcd1lgBKZYqwKmkUI6SeDDwHBZ12gdxhs7iUFz0pI2/7XMVmBd76VBL8IE3R0OUovfd
jXqXurYmZ7bhRMc1lXpgXxNy88ASP1iB2aHLpGQ1ecY4dbN67rD0vge1Vd4Y2ddRj5kgYiqyYeuE
TPFCOf4hXFPFDfeo234Lnzic30a+I9DpKZGCUyM5ntAFARjl8jDt/R9wTIjGaN+MrtA/wydQ2f9+
m60bBMvEFHIHeS7L0XX0IfJu6DGfLJteJ71IVoXUWNV1G5WHEc1IidllED4K0yEHBQx9ok25dd/b
E57cLtgbe6yco2Xcq69Hn85+fqNGP9EZC+iQNGHUDxOhWVdSccxP2vtIFukDhqa5J0AjtINIkBJN
2cDwTwFpmr8W17/k7tdldoZbyG4VYyiY9lvLoTKzzDSKkdHafcUvF/ZazO4/1F71uTgrBbFOEb95
7zWtsuqNQ51WQMqrbJe02SOFA2w0BUu4naNc/3Tgnwb9IYsDPQ8ANCsPi22BhkDFxD0owEsGaWC6
h0IaAUj4JaqBXzXXsMNH0qF83QnHz4/669ymgbPoGoC2rAzvv3xmv/yoTYpvjpMq50DZarlyokID
roOE900gdk9q8GyZy8VfjK0eO04BRF4XqCY7Yi9Z7Q+1d6yBMFvttG9TCpb4ktVqhezpaiKsRj8n
NpwaIalHTijSAYXi4oC5MVXzo5JIShQFqs6xjksDmXAOl/fZXIlSSjiVXPoUdKU3Bdzm+0SvniSe
476s4aq5ZbTYwU9EJnmBXLVgJmXJBZNt/1wfCKuwJlov41aqboU3qTCBhc+rCe9sKMbQz3aPfHD1
DWj05gpehyH0TGTaVZ33nEgxODQxLXttpHHoScAEWwPN0E6ZPY7bbImr6r7o62KTr+s+iegMuLaH
fLvYTMFlJOSK2HQIsgCwcUa2P9L8f/LdYXsSqgv8gElZfcvwc9bbn5tNofyTV68LVkigZFn1DJm0
Ale2oT1KYCKrgAvtv0LPoPTRI16jv0WWhav+CzIlqLJ6CTp7sFeyEs4v3Id7ufyqWNgU7RbniIcM
5f8E4Yr8XBFJ8x/MPE1GLR1+0hgUHSfoOA4C8ewcE6UexaUHcgrXMaU9IFKz0+Bd8vQYYsUqVVFX
rHL9/an0wGdW22BEnYRxUbJ8wgni153qlBPmTZdmTcUmKEdaDzMIDmxwuv/I8P7Rs+hh+/svw56t
qVxVZIKw7/gjw7Z7P2r9AMKVEHuWS3XjJzUB221WQZcDAeBtwG/56+nqh3cFTzjbHV/jVQpR+fDJ
8jBe22ctrEHd5j+Hiv34uxVq3AkgbCWkVJ+7cE06Mu7lObVy5k5lYrVUl8oeYP4h861fALxpDcZQ
Ya9LdewofuwfdeNPQ9uR98twljVgqAyC3FRRCuzlIyuOEyJD+3n+N3CzRnz/PrCyXRXSJreEUlvN
s4gKrz9jO91rYgaVqvWv1oonP8CStqF/q3Ke8uTRvtqEMH37nyLtyTJmzezWp5vbgrC1bn9LerUX
S9s6sWPYvXRQJjWYOLH8fOxuPk3MMFFMwBmG/FsZ5h8PI8tNIzA0RIuZ5rug9DOs0a9fxwpIa1GP
qmznT2Ngv2sCOTvFmzrNWcNALcgX0YSWEt4RpHnlPTox6HCNhZ+kz0iiFoLfSH1vp1C3nqfucoRJ
jKvKHHuQ21MEv6pq5BR2OM/rCwPV6TcoKvnLcS1UNIFVtZpvr56d36bszN4mgJ9Lows9rXriEj1B
zevR3nx2VrGEnyLsNTdmDpLf+LRPgllEZV4lqEtq+sYHeNy7OY9MvF8VK9QHLd4gZdq0QCzqwQgq
TDj5K8LmXaF2N/IVPCN5fWqmQFFMozDJRyj/KCikE50laQ8MvAJ2DqAM3JWj5gIDpbSpZQ+e7vSU
Kg56dW6AlSsR6LtBZJi6eY3hQXYlpISmIjKid7isMyew9Ol3roEsZoXuKBWXtHH3uU8J/nlxzadd
Yz9wfx52CLk8ym6cjKfmkQizoBTZsOtNH1NmK/18s59xvFAWPVWdxJhitDIE38qiht/dhHgki8O5
cnq4dYh5n3UVMpPMR7Tux+L5uhA4wNdemwK+Ulx6ZidxOQPmTFGxoxq2ZFGVmwaI3OzJzQ4On1jk
aPAjgBIQK78sTPLraJg1WfkVEJvQULzyioRe0oOi6XAywAtH4FlN8NrpUcDPBfBGCS0oBysBidJ4
CZwPGcuVHyTVrgvjF6JUhVMD0f6qB4bT93gOITZhEFq0GOmUmJqmL2D9taNNHV7cSE8gWd92FRRp
Il3Z5L7t92DtaKfXnQehfPTFcB9uhCNlY9p/MSGPXQ7o//Blg/iwmB5hr8SyAtanD1zf7axPQtrN
bc8tuS9ObUU+AAORIewJGEcc6ImxZMEKQuF40nOSRZ/X2NTLtcQpwrfh2UUIIKdd1sGpcfwHIuON
3NAFSwbFkPJ+iVOw19WeRPS4zsco8PfBJJlxXBsGrZJqVZj12RpMKsSY9Gwvf+MFXeCVpSTzQ7LT
qbegnYLVhziqkE2S/vmPW9El6vbSiTJn23kHF/asf1BkpczVXVLPKBHOEAetZsAWtHgAzBLKGw16
V634+meQXloUIzk+xul24JkAAF89rgIFdJkZWMgxiVtqm/3/xUNFkpfmajFFMQlIhPTSY9eOibev
20qwk7uKkl0hx7gQrY7d/8xZ+C5bteLHZUB1OetIUPDgp+HTNOY+ESIWJ+XGF4ddML0MSVYpW68h
Oh27gkwJZMFBKHQC/CywKRQnn5VfAVAm/075OvUom9LoX/eGDLDhrUaolbbCvaZaa/epDss2QhCO
l5+WcZdQTpKH6NDM5HoLoTIItns75nydS81W6lpwi1GBjtKzhay/+zmfZ7KntxE0GQQfljkOrzSE
RP/0wnQGDaXZwleZ4auiCCwY9XKeygfEw2dbp0E0WAw6yANZ+BhCChG7exIYGg9ZpINOvH8eH4LS
I2Ph3qT3kLc5d1Ru+yhnGl37tH6Cy/A7Ois2pS8zQ+2oTc2zyczNilHPfKhnvxALrvLGEDuUV9eL
D5SiHEim/J6UJ1u8ngITM4CKVUl9BmgEsZ59y4F8JyN2+O9+gUcCATo5+PTuPlpT4qHX8SWEWsqp
MFqY3jFtl49T5cq52pp/jPq7kVl4t5YkqQeheSE+zmEqdT/qabb1M9FjD5x0hB2yValGx0ZZ91QT
VewOZwUTQbGbNKpzOYMBxcUf7ZLE1BE75tk4NQkO8iZKZ8NwMeNghaLjFImMakrVmnixONtoEGyL
K/PSVdowA7NOqOIZhexHLw+bunSQjPa2TQY/5l6OD3iHbGB8HrQ+VnK29bTs+GQyr5Kf0IRjMzO8
mDilzC/FSLQsI7M0mB83t1EcOQO2i+O1HSBBS6Vl1UBviKx8n3EcM1Vesgzm/gr9NejdXNVs3xm8
pKI5ZqsgRglFgjPqw4saWcvi/nKNEVAZsyOuppzlmE9lIRmbJefiQpdlnE16dojwOKjljQfRK0rn
Nglp3fQ9cgN37viKTItEHrLorsr7IGUviBq9EC1DI0huBBX9CeSx6lN5Iz87ZKNa0c1NrK8jvMSS
UMzprnc9TZUw97XxOwu0XgP1SwcyRqJ5eThNfAfCpkshyOYmXaFdJzlDTNrs8s2QMWFH+GdWTBle
CmjzaXtssdI+CCbJcg2k87vbaz384FyUrXePz01OiT9IbLnQRltHtuhLHY3TfarcAaJMJg0mloX3
hArSg6ARBGCc8nZ6cc5VQ/H/nKLykbooFUlKuzmNWjbrCfdf2IutB3A5F6iV31NbNSLMDcUX9bLe
qJdNOCivZIAtn4/MT6S60fqrCnd1Dlkd+RC2JKN3RfvH8nA0pBSojDndpxejrFzn7LeH2dqcBUkZ
v6oQrV3Bjfoe4QJCKkdjZ0z2Y8jPG62p3ylPhB9QzBvSY4aG/oC/gd0pl6skeItCt5tPzNHrudU4
6qvsmcGE/rY/qpO9BbO5XZtkQP8ozKY8bwklAJkAYOwY9HBRv0FGj/3q8tCA1leziVuvzS4RzAJv
andadn/snMoKsKsd/13IbKNjK/ckr0+60olu5+ceMxe1xFG1zB31iZeBHY3dw4Urtg76hHsj9/Co
PE9djKa6GvY0nvGq4yqy/pNLBb65wFAtRkyvmILi2bGoN10hAUjqMyEYlbhk2iwqp+/+wlDAOrr+
LQSH0j9pxR8a7woMQEyFnqEZd8kkfugXt6wfEt7qq8GUoSho4tggh4Dgv2+Htd7C0yBF+s+j1z22
epilizYubf0I1BAZGJ5tLG411RDU3Yu+O5Mj2dlWvq/MzHHJ2+VNlr2ls3NCKdB2Py14s6wNcYrt
uZZI7bksYQZQDsl7c9p2TDOE9eH4eK0q8m2t6xS01qM388q1C7MXdEhgy6du3sXPdKAg54rdWBHl
OJSgVSNmTHtuBalgyAfZRHWYJmrCrUIUF1rC0ZPH6KYBTTbkBKEERvXHSbA+6g6HeobNjo05YTZA
SaEXeEd/Tmh1Zy9UN7Ftm54w0HTp0V25hIaXBDgSz5Twx3GJbgCg1c/VgsUXDu5vKIQtltLPVtlc
vhK9i8BeUrCK5AfQG5F0UaGG3kUz90+tVEiNrCJslu1jRCyZ6kkR1krgp4mfugb6ODhV/cPAKOHl
uUsrugByGykUjwjSP3eDdqFOmCnRFkMf5CoBAFoQcxSkTwzyaLZk4i3DJ3TH1QQOe6oTUQTE30DH
vXFO51gpGj39LOJXC9X5MPPkBkxxoUmuuAcskOwq6lRJLd13bBdCpXpbqhzBaKifbcIFuFk0+hbA
jag0Ut849zeo12UnM2+608yw2jgrOa9tzIUjyI80q/RP1LtW8tPUTaVve0vr9bWtBmOVS6sFv+sb
vGbZBxJ83L+oPi88U9hbopyGh8VuaX0BASJcV/SjdTLC0XXax7jtFs06iNSCZku3p9BHhzA5PZXl
h8Skrl8+Qt9Qws9PyKxpSjStAaWcdjN97lU8qVhszOei4a9iopFYaMCr2ERXGh1y3l/PlAJ1v/MX
oVeDo6ZMLcabK25YwrRW1UQCv/39/96KejfIPf2ITeMnD2doB8AVIZMRGmn6W84Jh/U5uLBYAV5U
mlfKKGI2bsLbxr3cxlW6TZRQBRLdGBgiCqBvVUi0mrF6e4Lw6kYDLDAROHRkCfL7X+YoynWayok4
n/XVMjRy0SszIVVgyyFXIFa13oq0jczPVzB2y6aN2jdTDVLYzl6vU9qB5MxvS2EMlj7sh0u9wECM
4aNH7qFErbFVgdYfMBkqJLB2rg+2x1C7L9fB8tCvjw9O3B+BRjzNdlHX1tj4thSO1BonhdjGZEhY
hodd2rRqHtYzVIsKYJdYMwRDwoyjztRL+8Yv7oKDkzrNnV5LvL6ZyH1by1/HLGBmgA8yE3y4OJ2A
EmCo7vmRj7Byh8xgeFQAJuudQhgE7n6tfLrkMu0A8btjtYfplt3m6T6Mn1F7brkliWgUxD/kg8Ah
w0VX/KlEhs3oA/d/RcFDQlVkSySVs2+6TEutL/HLVFpc8jHiInX1u8Mj91zBCCFsBv3muIqDPpqB
JF5WTMOj6mXOWseiwoQ6/p7LgeWbQR/hv4xGlvHH3xpkuPGVguwWtwufTh5Zq777ZRJb0ZyEGu5x
cywQCNvaD5AfFR5RX+oeQJcdn7zupedbPYVSaTesyBK30FNyCRnqGpjbFmjyLdkJmAB6wEcXDw9s
j3w2cVrPpp3Y2WRUHbWztHCBJ/hZYrCfWoExjOTMbcbj6GwV8KgO1ZnNdmloLbJZ8TcWKdP+MvgM
dLBWP10Nx2AodUb7soMgfQ6AeBw5jzz0n0ahm7qi+D/a6JaOgSYjj9CjRl65+xGASyuo8cxIT2g/
lWTdM5Ox5EI3dakL/2Yieoxpdq/wLLoTUL7o7vf9W1iJ3Kcz5I5GDmvz2wqzKb0mL7vJNyFgHANs
X+XQtVk958QeUdtSZCOChplF+4FaNEmyES6IwSPrtUTiX559k5Vdeuy4IkAyMhWFOwYscWgi5Z4y
oqR0/K1U3B37eKg63PpKXg2/x9BhxUdAPT85VmboJ04W89ilwepubE3oh8T4WNymg/ufq9ljlo2X
GCqSOevmGp9POdijqOnWkFa07yEEQX0SLoZqeiSCLgnZw4ii5Zc+9II32Ghm/DtsUJirKpek70FN
lXMePl6B1mlfDScWYXYG2yQqLnt5u+bsEW8nEa7PDdBmMc6pBvlLmwSgIlgJ9M/c2jyFO2zRwKRD
BXNI9NZJH9ovy9xVSc1haEXYUvUYXm070vwB8mzM2bjPlaMn+RY0kFbKIUne78Mhc+h6mCtBXODO
0mAU3ev2EWZg0g9y+3L4zEMY6pdC6ozklOJtJ2UK2qI84klBgOtBwigGOApKiknc4EJiSd71LfnH
BVlA4ScGq/OZWp9OACnGp9Bo7fd58kPW3rQD4stNa9oudrOand2z2owK3zaP3rVLFAv/mkXauCj2
nW3kSlos/TJtE7jb7Lk6RoyRcoBSuIF7qgHjcUk217em2759lWRqjX65LXFn8xq9NAX/xkW5QeRI
Z4sAmddeGNFKRm2yuT5LNHssBTrAG/vEAW/HfoAEjZ9xhqRI4oECr4S8/S4LfHR/wKOfWDJzEako
1hf7XpONkYCnpQQLf3T6s5Bmg3VctIGMY/7kQ5tsWPtYbuhZpOIDsU93l9P6J2RGA7B90g9hGE2d
kWY9U3LpTMqKu43gGngryGt0ZaLPfli26jPXaSEtWedOjSt8w509Q+Ca5N+pDvHbAdYot4smbyvN
YoiVe9KhBAFTGtRHIkTKhrfp201cFEMtIwKVufFSGLgy7DKaNJI8dCrgCFpX6FCyisQfBlMBv3Y2
8TKxHFgWKIHSnTPSQW/bqAqF0Y8JOzneI8PHixrjYdN2E/Yerav4NqtE9ARXMSPM7EKrtzFfFNtD
YNUJRKjK000l6N61wmt1za4KMnGuXa2A0ACPGcThLcw4UDK4D+fdrMuFcvjSKH4+gG2qqADE+2NE
CzAbP3+FKXHm2P+eqrELj+6QOvT/6VbWT6ZaxpD86UerIae66ujzP5t1wmhasjqcJpcjRTZbO5jP
W4ZqU4w8gBaQnEla1J3+yW8xksGh/t3JvPd7B1WM0MtWbabWZD+RlN4lqaBc4Qd3PR9PhiqKIvyW
3kNlqZTVtc4QawOwaBhDYufTH/irDy/85tvHTb2JieGX22lcKAVV2Wxr02baP7iqGLHxIZtgbL9I
lgHkOzT6i5jllov3lTzh+kRNOKi6yvCsdud/cRSniVjqmnmdjbdal7pxkM7UaGXRbGG/qGO4lacr
mP/Gh8Y/umd9IxQk+dDLmQOtPNPbGF09wKZTvSYfy3x9QykaEvzKf3z3lWJlyjk9mtAXJfUt+f69
weVwzcCHUl8f4Ft1MYV+rbu2yrIKGhPe4a6JYovAG1YrZfQuHBtpfaONsx90osZJeYpuvmF2srb0
c53wRLWxzaymCpjMdA07v1bdR9f3EYbGP1aCnWY7Abfxkckc8Xfstv/PYNHlkkrpkbt9VVoAwt3M
7avtTN7kjl5qO1TiwxWHfaILaugBYY+97PvAtJYklC8iGj2b50zwbdLctqo5kBkcgcH4lEaBpC2Q
yLJ6xMl6Lz46Qt8IRlIS2Q6hvMK5kJwZ/1PlomPdFu1DJkM1H+gxltZPPo4BKtfcDuOLcNbPH3nU
qqfGjnv3MKuqVoI5AhEJU9ghV1z3DH/jC05CL8Y+2lx2u4FP+A7jnQ/v/NF1N253wimrjBkvJZlQ
GV2Me/vmDi4MvmBjZJf4eZnognK2m8EK87CVH9Nr7zUMoWlK1o3z7EJVc8TH8pD6Kamkl05c8DeW
Zgs+ZV3v0f4Na8FvqRu4dDDTvAX7DNelkr6RST8mZNscduxb+mlPFYYV/nBNLVeNIuq4vxLrDQm0
BKjjRzc986kd1EqsSgk/W78IP0VeIeTC1wil/zYyddd7uNSKSIQKP0LOoPv3ErZdKeCUBJ1UcYqD
zVBy+KByzL2Fl0joTCVh7jl86xfOeviXebL8MuWnXFY5iURROmh6IUx8x12edVQ0vpkAp29SojJ5
SBgG45rvHFPyuf4sS9ZfUXadLmAr2YCDqpnn8Y9W3OdBxVFqEXesdSzLk0VcdFFOJZ7NMd6IReXz
oaGNkZ98xS3JTaX9dfSN+YTt36CQJyur8+rQOLDLLhv7EKAUp3KOXdDChcFehLIaP/BXXf15rQBO
ATfKYQhMz6rDYInvyL5M1l6HYZ2cZboLhP7XNEBJeh8YUKs9cPPDISnCKOioeJZig4LUJtobqOWt
x/sOV/bCssLfoygFHVjFHY5QbbeXfZBfxE/Z4FFZ8lq21Rk0w81JhtV4G+7H2uCUfqNwxZVHY/7X
vkbiCCbf85uQZTwDJULFRKCirCAV4aYqsBvtviJeZSc3h1oWAgmnva6maM1Cdi7ay9dH70arJ2Ts
6TX/xqTdcF7DpMCBbXS/uy5+QD/xZkCAbjUawAo35k+JV6+f+jnrhdifX8vDDLSb5V6NAegiJbXT
9iIRJKPRdekY053plhINNBIxLviHyOktA8FFpn8ksg31dDX/whXgOD05nRXEBzBGUUEJQbdUnTpI
H4PJ4p9yNrl1ifiTdcmW+R6He1+/FY0cI/43bdmsctDkKBW8wZgXfC9MIpcMfqRLhxp1J9U24q04
sCvg7XrMT6PMoXDa5jTC+yEL3YascsopfqkSBSQR0pZ51wArqoP6yXyvCLbiaPhb1K3RaC7M/Zt6
B/V3zlpeoWUN5H53qvFZqGsoMxxrZ5KtwAj5TzapL+JIHBCacPVZhp8tR2ePZbNEjdRf06wKDrmn
dJtRX5WF9Bzp0V8sf0yi548L8qsoRXvtnoth8MWR6hBPV/SFBbQJ8F90IQ+lNQEtTi6+wKFKOdAV
vcS6owaJoQaMl6C3HtiUD5nROMj6hDRL6Nsn/f8zG4rQVUQzmBSX/cA+XBmigb3bwEFGWAcKAd9e
dO7YsQSlbSHU9iI0h2ccl9Z6y+Taq9RZ9WC4T3AIctZ8NoC+Oaq8UJR/3DrEHpWwrTTSqoQoj2+X
BgjlTRZsdewmPBWy2Q1WDEvjlfKX1tLc1Yy6aAO9sFN7B7Lxq+Xsb9m5RwMWOSJsaiWVHQQsOgOi
oF1k2NJZRCdJPDGT+etfJA1k5Qgxyg5gxuJp4BntDIpNvQ9E700pMzquyosZcdB+VtuppODpQSeq
6xrwoCkWMw+hWBEOvGT/Va6YWmyMvw1r7ZrdbaAMLYNiAz6EO3WHvxVUpbzgkUljhtdfdsxEm0aA
hXSTjeEzVPnxVVPpO+cLeWLtzFZQ+q5iK6NiwMeL4o4pdkrwHo0ysBq4a5ZTMvTAJeaWlRrp/be+
DgtFn78ZnPvjDtTOibt+SR3l4Qmk4ODN5OyCDXXwR2hauzAROX/5oPJxdutP4Wet4BMfmtkQxkZq
vj+WQhaUO+JoDQjQ4Zgnl4uxqy2rP1aDm+pX/tX3HhKfWhdU6ELHFz/3choXpUz9kBPRq5E62tzZ
7mR1oDSXwT5F6gGaJUMXIJtCdI5QA4LmN5QQs1arrxfjiw3rYVY/27HY7X4uwumgcOyw8SFMrrUd
9ZLOmvHSE/nBnHgld3nzmoLddts7zE24LUErmO7gef03DonQcVeAmyka6Gp4aP4xtJU92XTSFnfu
+maHt1jFywTqjyHuAfP5QIuocPx7LBuhr+bZWi6uLxXYck1804pUrl1su4HMp5eAp5rU8lziNu32
2NHRwoSGJ0itriw9IdCC6dhQAK7MnX/+OQ+auNn4rh8kBRfnprOrJnUKcDqncJEzw2fPIMI+Z0yE
uA9GaAkAWL0XlR8J22NTJK50Bo5dn9NnvRMqyQWL15wD8c8gdH/hroXIEeRVr/ZwJwseATJqKTnh
PKyLtdHdo5d+Gmudk74hjL3mQGl0/vWaKzFGhsikUz/LjQx2WDVgxF7aXZ4RP82XMmHxycpHnsd5
tNWo70XHd5CUuHfalXwqlz6fCtRYEYz4kOV2K0OVKNZooYEtHpI1hp/HebHoSczsEj6neSoIGtSh
LqFmh4RixJy2sRgvkHxGWH/N7KDYtPOwT/P+rNXGODhjM/39klfNR/xoD4dlrLdhKc/7kbWPCxja
JnlUSCEtMTOuEs8QiyrEleQGbmjh859ACtUMcpZYmeIRumfpdUm2Zdvj9D2jYmgJVVy2zsJBiG0W
gd7eeN0TZu6Kfh3wV0NkFskdqryjKuzYk1Oz9r3yV7qHBxFhdM1QRRIYZCea++Cp3aHDuKfojGqx
xIIw8vGfj9qVVeUfkXTV23OOudFhQKBRcbglstoMY9KfYy/RFxt9sy0aVdCkuS48lJWdjQHXRnCl
E/ygS2YWxZV2TJ6bXMIGWMlQ8OCT5Cc56yWjCOvPl+bLFmG7wB2N3kpScWp9qHfKGtZh9LEdKxod
Mha6Z+Fwz8myBs0EPmGmN66yIKMX6KCMhYZRwHxD98R6mJgGL7uSiyuO1n4VTbL262E9KF74hTAD
mkinbvXPRMrWEt6taRiDmDyu4122uMYOLxIX9jsDuZQd8HaTHMzbTC6Rb0hp8Nw1gdQ+JuibpxmR
CtXDk0PLW4IvOMV2dat3x9oPTnkEHQjo5rHzphWEQC+vwe8y5S7i0Ezopc0NmBZHHsR6FvzLFojw
8m83YMNNGd9BNRRmAnJUfOJ47D868kyXHcDt6RK5bgD+oDCK3DIXIWZytE0mfjf+3gXYjwd58Wof
rm3pV8o2QuZLlRRroLvVqb2irPKHylnEyPnIFtjwbBkHGRxXfD35v2gdvNZwt8n/G/FB17Lsfzx/
CQWxP9oVdWLL8kfJgcGJ6Pi4IXTBsDilhRARwC/+aGnLG+SXhEg0Ahc+rKH2DnxhfjKMCq8SdGYi
/eSr0XElZvPIS5NJNfkX4knWarcXK7OTk1QCVK8uI9wjqvoVHBSxANuyN7ONxV2vx0pURP2quP2z
F1BIDMCnkJv373oE3Rkw7sq1kWVfFNE4lz2ylDk8h9j5ED7IXNltWXiIHweVKOtVUmCe9pd2kyDO
XQM+FXGTUQw2rPod0ttqE3C3N49v4fII00KOLuARHGvEgeB61rhlliZfe7FeGLNDM2jUN3l+ZPzC
30iCaAtwRFL+7SoGMTB1+ezxRB8akjlqmly3nMtwvN5GRqbNF263ka75tYIHuXIUeE06cFYWKjRn
eD2fMmQNvdBN3j42kRJOKVHuAcSrOba+E56flDMKH3m1DNtPd6lkKuxkI7zS8zvE+lCtyglFvr3t
72gqT2HFRo2SEc9KQgDQo5vO+xThCmujLHSCHUV4dYvWmqsGO4A4W4ZiKIsWtceYiT5t+HOdt6io
FbvY28Rj7g1a8U3jFh0f5EGb+2TfOIP9Y0XuIVVzxMTXlAUcRnezDEw6326IGlOwAet5o/d4IPHk
jkml6khCdEukxONBJ3MTzEdJcy1ajAAyKI19QhqoXIe1SgF3MdXNfPAMu49D2x3SJfbDFLfO+WKD
7SswmBFqtQx9mzsRzrRIVxm/HBAH2TrCbxcqdCcavPKZo4pJ9Bw6SCv/OB+hNtyJb4IYAkJpvt4F
Mg3g7X7gLQFZpTAscXog5BBLu5nOHSrxN2Tt3npit6ZS8VwPQLUSXIOgZpBus4eTN5xzhaj+vYCO
qbyEhlpRjYuDh79JHF5L5/V9NH0h80KXuVB7wIBoIPLKDUBAzAsljGcq2KlK9zFKpvVvGVLrkL5H
xjwIGvbWSp76vUDuIAxsUZW96QofCesDWdhPIs6jR1SeFxH2UsfRXgNjZEjixe0OFJbDlbfal5Vq
KeIEzx75swYOnm6oAd3PjOEX1ryyU7yDWmEdK8wChulP5TsakhZZa0jkjTXbLyv1mCpDrp0+GJcz
KNaQBNggoDl6cHidfsUJ9hvNpqpV15tg33Xrb7s7mQSGtvm84+ieKgiJqUfLmb/IifEogq4Nj1im
46dRS9lurapwdfGKwAIpP8TexJvDWmRlaeqSgYqeoTg0xi4neVcKiSt0oSoFqwVUenNOZwlqR+ip
4v1jhc/hUSvTE4OgNBc0CeKONppPvuYi0V84J4hFAUmfwC9k0Ar7oQgF2koWKPo6aJ2qP4ROB57Q
zqzYcw8BWCTCBtdgUJ3xco9VZy4fQL++nsJjHeF3VBLlZVQ2sAIeC+SlVzqmPaU2G0vDj+n70IS1
gTz2nzvvya7qlgK3Bvk2z8GDqdFP+/lBNpDX2iyMOiNDwMHh9+4jQFv5urmOojXKkbSxwWQE1tEY
emEVPyMx1rI7Bw4Fnuri4j56DDobTq9MJnMHxNv2EagZeQEbqa938cUNXiH5oKsfuViWeo9Q/pnn
X7gylBCFxWNu+2BKiuMykpRf+hsUgVL/OfHeW+sJc7krBR1Ufd8PmJ6qpkl26nOkeVPK8CQnoYSY
HTeDmM2B2uiFYbYTRGPhPsVo5ve4zNtx2nYQBiIH8MW3zUiOXy00mmnX6ZpCUKr/aN9pj3o81qtz
rNaL8MQ2XSu5ufKYN/aO5H0iKO/F6JiTdyk3XlkTS4Wo0d12mOmFIK3FWQYckFh3JHgpnkWuOphD
dIIJ4nIzJ6vkmvYNP2e1O0ifDASKowZ4M1TaK5c6sC8BcXhKfg7R+rdfghn+lvrnPu9uYIzSG6eN
GljjmgHw/5BHxeObL/33k/E7CdGnjPCE6ng3S78O/wnZgvd9P1N/DxYDWatl0i1sgPEIZ2ytJAFK
KVj5WVrJsmRDqLnMuBYVcDSgviTaKtzemCO039JKJzOL/A6QdzbVzki3N2cPJiE067Xvzj/79U8l
AUkx5NsNSHU+yG0C7REvSZymeZ0HB/OesXoD5mdUFrcKFzbbb7ml6+jpiXPFIQOwPok/bViRmC1E
pSb1QNP1CBAkHPDsIYkpe4p4T895IFhFBPGRyaHyg0j9l3blzVwwC85SticBCwNjG/YpddIZa2Ux
yKMbSCQhlRpREKZysHRAsx/5CW8AiGt2fTNhXiaNsEx3GfeZMaWVjNePIVrjq7KE+etCHP51p9YG
zokHWXdBFcWhBDGfnD34SCE+nlyO8HjV/eM185IihcFrLyE/UqGEi0IhRh79lVxhxmQ69UsNNTJO
CVMzxlW89v1oO/bkQQLwCnU8HTQ8l6qdSJ+FkXB7J5rYYwdercY807pC1beKkgumApLVOyR5FjUm
oM2uEaTbZ2VVDR/suB4Prk183lphTJAjHckHxwoO3acBMarRN0i4/rXZ2lsA4mjnsh/PW6Bf/5ro
f+gKlwEmq6iaqefPWV//znnjnVosuPDgDejq2DGYnHpQH64fif2UZEK1ILIdYozJOuW1CbRQLK2L
+l58eDiTQUYknkxF9LzXO9GFLYHkxAZUZKJpZYEkMEQ9IO2pRszlpqHPKGHxpxPdEcTE5oYzP8oE
WdG7ReyRV6XYauVYAV02s4Z8v2wa9AjNL6AjuOUFY5ExwBSUm88GyqAmMoiZ1fFrQ6kLv+aaJLZ5
FQThPZKmd8FYdhuRwKwGPUHSdC6pNNPp45yXZsy7m5+S2TCOMUpKwzOdaaBIdgC5tPvLdkVuIpao
VD6FDWVdS8WgtDjxEjZfVa9ANjXceST3jXktDS/s7SHefz44W/9skCSS2IIiOyTDsjBUPr6j0zkt
BptY3yET3dCg2Byl3zuz+225delRBjLEJemUS3RhmG7dM6QX7pd4QXwZ+0DpYp8nvb9DOR9mMEDX
mexjD9FOXdMk7Tudgh6F6T9agiVWjAHC5SMlCaxgOvSOsbuwpPppy8t1LqgRofGTx62hudYMffBB
iwFgHbXtOYs4VyVFAKXPA8h8Fjjz2BSt5Gz7TAH5T+GfPQGkOxQpDpy5wYtu2nJ/MyRPODcCQr4s
F5WlBfzA+Fd8vsialxrUojt9UoxPQIkvshDwfcY1Q5bmnvLYBX16/BA4OWckJBu1UKXJXwUZ117d
aprseJgw4GU7B5Z593jszT7Yfs/ElW/aYCEc/+c828mkaQ+zL/LUv7IEFQFYRZE91p1H6wHn6KRY
X/fUYmOKJCqtSJv/noIaDCNrYQ6vNjmGLZa5rlb/xP2e91mPCmE7cD8fwvuVNAheYKP1kvr5VmYp
JSz0NeJzAlqLnVHfS+GypvhAeFBGo934+oMbmm6vkFPbTlh9F6RC1lH4ETPygOfgH1GUiXLOyuno
Qpr8GXXN7ACu4DFuWnclsNOh41xlQ/ylIXoFdY5bLaW9KA4cBQ1jJlC/PStV1riNJlUHm4SnZpV0
GmzNmAGqYQNuki4hfhh1TbHJhnKjGtYDUVI/X38cUkMhnGlz8o2OA7bpbZVmaoQi3gyc5JGZbxas
h9WEQTbCN00+QzM6ag+t+CMzVZzn5I5oqhGEJjj65uK/FUSJK1TTb16lqwZcR5tXdaPg0nMYa5EC
/3YFzGWj2kZvXVMSX2gifxLVm9I51uaJOikWeFPapLNfOt8hs/akib62r3kq6bCsnqgBVpnahqH+
7Dfrs/G+ZAqln9v/3BzsFd7gKHjLJK/Lwr0t/TbxS/pGPeJ3sicVkSDoy2vxHP2+Vx4JgUXyGb0L
09lo+Ey+F8L1PJqFxvhSTgBdXIpWIBQlOgYjDB3vaD9rZJMig27/3C0ZR/QCW6RjOTgSn2mj3hJy
kW0j0bnl8YGwtRDi6RZYRKpv9u3wrPq7EF7KTZSB+OPt9l+yC4d7srN2NXPwBj1eVAiW5KdPKgwg
VC4CPwbJ8CBgkcbLMjKrvlLJPk4HD8r+bs9t5NsCeX96nJQ4+S2DD0B6CA8OKz+g3oUK15yfifDU
reahjYBeZkKqr5HDO7Cp586NnGw10qRj8ckGZTrdbDXlronQmfr+gMGssw/ZFdh6g0IZC7ZiR9uj
9EiJ8Ds6fIU/L1bVhDkbZl3S2BLyiCEO67dIT4M0Y4k3qHVCt4ZyEahPx4OUPUf3Nf462b8c3WPZ
yKBV7h0o2OUqkGksNjpOvs0w3QpdVIju7Mw28oVL4pUJ//FpQy+YMxFe/mMf0uoJlntdCx1Kqspm
3Cr6TuSv6nmoEwfRWBd5PMbIAgoWuydQE4FmhhUb6OSBZpZ7HbM9dp6bCT/DT1N0RkNlouhUsW5E
307J/q2mV6tdcXdaweC42uH92wiJ3+CKlXom+/dd2LBKv6z6yIOetXuBw7Bp5o8W3Mu0K4uksVT5
yddk1gBlxV2peiKqvrv+S5x9IU5Jj2oo7HcEzkh886561BPf9KLj+sCEwPfaGMFR/qeSv43ChiXX
b5x3Tf9+6CbZMJ/EmIkyaJURMgJkdRb9ckVewCuJkaytyR24vtucksOWtypi4k8jdKKUN1Sn8EwT
NRa+Tv61OMYnBata4HvOfka5YmRWEyXrD1DXWcfNXjnLsCcC4lzh2joOmB+Q5vNlsin89ShkI+p9
3d66QthlYLWlFEHocdP49OT9VEmJwcdfrQzfUMB/gxoD4fFjaWrWLj0JOCBgZIYvnq9xGKa9bUX8
cFjkCDUvj0MNFvWF8RsXIoCj+061pZXnAlDBSvHpTGF2W6FxJU+W6f1qc4nFkU2AfBCOesyFF9AB
hjH0Kcu6rGwl153NZj1nAZLR3DkU1JN1hoSEuhkfMKr1ACvr8I40/QPekoGT3dONakzdROQ2UE6w
zc7U5pjo9YuW1LQJZKorNiRv5YX1apKg9e032Y9/6fW7iur1K6uwoZqx80Pg7JxwWZnIc2s8nDuB
QaadsLwXcfZ5MR654xBJ/IYxzVI398W9cIdbianADEsZvpu3llR1Z6UaBjjDM0dF48SvL1eqx8h/
ybiT8TXLuS1fPXDQzRuQ0J7RqZj0Fa8IJCUQw985ex2khaoh2ZogVMudksGhw5bLAIdrpklR3348
NiuUU0/BZF/xJ4KYadO2H2KZ+AiLpfP/pHPyywaUMEuDJoTqssNnIvjTQIWZNRm//1O7q5/4C/Um
GVx6z5mZt3KrBx3cXxtF9HpntoSoNAMUT1nG2QT1qvdZixI80U3IQc7pcdNdKZ9LelEAb62W4KCO
b5ToTOllE+Vsu6z+JwYhsSYbSS260Nzr22QyOSsvBLuSvFZ2X7m50JVXa5sdbmgTi5Lq0egh0CYO
XaUb6kZ+wZzYabWEuG17dXSVU97rQE6FtqfnIbfbuH5cC13BmKnxPjiKpBNJCsesPFGKuRLeNIxK
segNm8u7eir9cYnS+yWVMDeqVLPQDTqkBu2LMPopiCNW+WY13HQg19UArJDLxJDNhjIwX8aT3+zc
6eaSZvD8ylRM/khaOf62jovz34InA8t2t+ZGoMkx+e+3MYOAyMuqz0uI/xuMtZGe/ghIOurgGcFg
p2ljQ68uLI3DFiqxQbckA+7Lan71dUsffskcgNhVX3UG2Xdo73JQVhwyGpAq+LbEAddepQog/9fh
I6/58cVBuvl7WdeMQRuCq5G0uAa/aeDMIrteM+9NW7AY9J+tohGQD9Y/KnLfqAv4AE1lX0ezv3I5
Xa+TxYpB1QKbLV9skHPpDytg+r8+pZpJcH8kUPfuDuvXFdPZZGBMSZfW4+F0OQxsOCbAYdGA4318
4D5lAh/e6Id+SUjGnK7jK8OQbDLOCRtFuAjyxb2Apk7uxfMLkzTVtpXuOYhDkqpaSgG8qgSqI9VV
oKuaQJL424Yt7+/ncTjSBQf9ziXIEMt+U2FQcSnpjuaKVcsBqhDaV5Mets8++4/cTdAcdCzO3f5v
rrjQ8lREjinBIHd9X1C/9OanCIWUWjO2pf74NPBtfs0zOX3Kdv3n/FiqlSB5O7U4DY6JP3xxU4Rj
nKJr0yMal9LpCgUck+BBQYUFec9yeCQOUdQu2BXdWfEWpTiS/6LDvMLWNC/0FqlBxXBBFNIymo9R
tEsNFpM/ny7oETu1SwTIIJYRNjTzCk9kr3gyADpHA4RLNvonUoghKM6ROgKATIWo60omG2LYaLig
Cg+G6DpIpx7VQwwLGTg3XobEA0XQga22sEA3HbZeszvCI6okTCEl8WM9HNaPrx6eVbZ4YjBdB3tg
oNj6titUddX+z78MqAEdWSziGSuV4KCBZMgQMkbAaFJnGgKjheYXjlRyzSbDoyfqGpgsTFKxK7vE
hLZxG14D1TON2XG5cE4Mihxf2cO8G/kAE3CGz98IJA+97euam6XsJKQniC/YZzaQViLUDqt1tikw
PmFHlUN/W4QqcMSxaY8SASJ+iJ6+Sk+9IV91f0iQih93sX9J+D3ht8q76N1TwCheC5NLHtWCeQgc
fgybGrhGTFZK5Cw8xs6k1YfDO/4+gb5Byk05QTKt5fPy06/YR8Qj+ROVovUVH3Nrrgvsx5L/s5Xc
ptG3FqcVa0MV9vGr6z9C6sM4TiMEDl5B1wdZnsVJsAKTP5oJk/0XeVbAbsbI9taM0U+eS0HrpyKa
GuVuApCkISL2zHUKlZZ/usYFEKa4BmTlUHwlEKeFQwtTvwvRulhQG93XfFsPV0WVD2lKZejQPg+U
vohTxVt4EWA4orU6EmBBCOQX5cdGvPIMp+ZeK2nANY1fQLFidEFNzpOuhadAXBQISHXl470TNruV
SRqnNAIWSm6Ltcs4JgnVxPfo5GYYIk2QGkiqjiia1X2wdjAPb2Idp9bcr3RzF8MbE8GxOz13zprx
4fIffsWQ/5+hZ3nTir1A4UW3f49YFibA3wYUCcR56a+CK6Jm55+ZkrYrE7/E0e3it0IjsQ3flB/U
lolVWH4N7W+jh62AqtGjGqw5lHOzD1MOpJmBG+gHzwFQn9Wn38HPiHCeg5/kHgTn7Re51JqqWq3y
rJiPdiOoj5+F7jMYQMU9a833mc2QE0wExwQ32hfDHjcXrNRKU/FBGTPFtrK/zG6v37L3XTH1mqic
NixIhU4IqhAnqs6RX8KP/KgfUP6bdssMT5lE/wj39uzj2Jes1kBgr9EmjvIFLaVz5I1e3jQlsOGP
e1K99oDKmNQ12KuJy+szL40v5k+GVY9SaIZC6a3xxCL8CWgvehzfqh9HEWpeE79gDcvBcMrTHrZr
AJ4h1o0a/hW00czMD0plmv3khaeJryyUSO+ZCR3wV7OPIy45JLlGvvP+eJJFbjixMHvvU9Mes7Gt
HXLg1pMLaMu1AvK1DnfDyVMfgcMAdWkaTUeXUa5B2Asj7ZUf8ytLQyCOK/MYtWXl66ZBgkoBKx3/
Q9adK3mSqQC6vqutSESib3fm7tOGdr7YAOx8AQCmhZij0VF2Ni9LJeuHeFa6KAs1VfnDfkge/lYk
laMKBxbXFXpXTL0T2a1C7KqCt/T0pujGkhQ/UGPfyvjQKZPvyyH2bMZr0qPSl04tK1ZkdAT6MZ1V
/Lr38w7OTvwWRSZOVO87c3rl0x7/YVcrSm6NZNULLVhjhr3vNFvu+qIK47UAVq2UhoWlqd2Ns5+K
GbtyylgqxfmmhJ2mB63wVYqstIPW0DbKsRfLX0b5yBtlQUXd4J1Ah+2/N7xs3P3tFBt4WhikryZt
sbluLTBBf1O0Y6PtQCps6T9oCQLKJZDy371l/GG+lH+09TtuFjd79Di5njI7XoYjVPqmkxu5ajD3
Mis93YQieaVC/ScBBzJxpNqOHcZG6ytnk6SKA4szrxItr0572GEWNvo3KS+CnPEG0iDnEFWnWsNe
rXMjydRcaTRS5aoVfL0zWCQHSm35rXFcjrh37+UFpdeSyFsd1xMujt9Ya2JWbwVb9/RfFWvUtEDZ
gT44XaiIVrQV3O+rW6ccSDE8+xs/X59l8oN8GkRA7EzOxIIF8h1xmOFxJ7pd0OPeduiC8CPzDr33
3qMPX9JDSXyWztczFG2V50v2frici/h2qUZPGX7NAyvFvjp/KaQMrpbeuX258b1xQQVxY4Icj3h5
NieeDtB7Dm7ut3j2Jk01fVZFsakhFrnDjehZF2Pk9WQpHmHN1vJkYNADxIcYEDv3U8JGfowHQrwH
qApyqNXDvnVL0GP0pOG+xddqeMg2sS4OIwkSqyqmot/uYBY2WLNK5TkmXrqJYnmDGgFMPuiJINlv
orV3x5DlFlGJ/IPj2xl38LnPYhurXQCbfKPzcFAlWVLHXQAbS588ylNSjDGuOGdILJkYMBx/hEEv
gUiX5u41su/LrRclwvTB3v3NlnRyfoVOo7DpukfOBIzPTzc6PaNAARvstkFPkxGGn/PNa9kSYb0w
EVUDJHlRGbciYgJBS2faVL569LpuElu9U/GNudk+31deXG9CvexKrYb1pzduXAEw3utjGnVAjjiS
knsRWarWvp5sAT5Y7WDbXujmMI95UVmphqcUeUDyCMhcdkVq8P+6q0PBc6CBY2CdxxybHv8x5fyD
xfuOcS/1gdNaXN4yU5Ty9RFtMbrZFHwNldYY/PSsc/joidvNsFfHOSydIe2HGSwJemKtLrWkCD32
H0h1LBaJIorO7Cyiiq03Jjto5YJ+BDl6sQA5MIPmUiAf//ISMfaFSgRP1wn52fGvtSEYdzxzwjWz
i0iMHF9DwXNu4aY+ha7/yynvrd2D6wQ2gxEs8w7PPa80+LmTnnKOTukpwA/sIc7KhMj+PdTOKCmR
r+T5hEKhncGHMvofJ2ITpPxGuaqjAKf9pCqbBsZ7niQL0T1HuxJwAYrxdzRhFq6OD03wSMwRZe2j
FtkG63a3Rk0Gt94c1iH/lgnsfzHERHuYKZ0z+bmszgRCJnMXO6a7r8Z21Qx12dRclZsut1mpuwLP
C/rTiz3g3/Kyg5fSQ/TBuOlO9ddNfhDFHYhsHNgccZP7IzbWNtcLAVdKnF9y4y6h4ouoCWNne6AY
QTNVSvaK5mT/1u7GJ0jph37UUlG6WsYC6+TQ0w0RJUyGaYfjph28AmGISQnuDpdzIUohKaneXArg
wCOL9tshadGnYhIwLiRTErlgweC8FQUPlwryjXlobZ8r5azA+n4eq4MHp9LX0kdG8sHpmOixm8Sk
h4Lj2CUvO90AhmS1SGfGO3lNeASJcNzN4ei++TnlC6TicTI/yXhVjhXaDLNYsmOhBXafWxtw584x
PqXabKJ34vWFtfglXfr3LeWXWQi1idZxHGEze1CPsZCIayUjN8YwKH8o//+mxzHToCGuPAbC7GPg
YMQMuVcmJqnbOXTrUaXOt5KUF9qlk/LVRlgCeqWZHJcomYwOYnrLVX10LIAom8vgkFW0DC2bI+0u
76YYfUHEjqAQfMJ6PgD9JJdjMSFvwOsg1Er8/eGBDdhZjTSw9NZA2FlMA5Ug5dLl3Le25Y7OaSpI
TaBR1H+82WjYQm4MUWjRV/pDsB9S93ryERUnQf5Bh/KiBkchjx6PSguf+6+k8IdtOL6H5JYhBaLj
7x9ZvtPmLqw6Vo8dp5XIj/qrVglqavOzs61vj+q9fUq8wrlwaPyLW7ghNF2gGnIiJJO5vC7gewgg
Y4//233tbLXYw2M07OFrzfjCHNpcbyz8DkxHCMvKQ1uvu83tzrKP2SdEes8XnvIQtu0PxfLCMOTx
oGUEaBhqWnkBhFXcRha/jmH70ke/ZnwnCg897DOTUEL0FC3ohzqd141Zfc5xDxnPGb4BAKuY3F7q
GiUxaALvcTa90N5IVIrz5z25qeldrUXpTNEFKnnfMGOpefuvgUoMAG+0TE0gjMzPCudsF2lPSrZg
kI7GO/WtrX4cSikLRscATQwcTPU7EeniXRIJOCC/iZCH2ANdizEvOXVCFwciI6bZqZdLw62JeQj3
kDf3HB/Gxes+rScOQS9EWxwXucH6uYyoZXKX2J9b48oBXy70KjtWeuVTj3LKnvuTH72BNOZEofED
oAJRevKbENuFAj20kDVveuWCNmzXFMVevdPezkdwrOljpXs1aoC7l1QuEUSKymxR8KGky1fy5zPI
laqgR7e1YkXU/uBh+rj7nj9ezX5tIu5kinzbVdG88pZFVCiteWwL9Knez9gEuNPvZ0be6PaW4LVg
KP1G8gf9dkZYEjesqcIL3EF5OH7FTnOntl5o9+97NY1/OBsURuUNVLADCe69yjVxSBkE0gl9AM+N
IAj9nDEaCeOZkDaCCxStntDNeU92kpeGac2C8uG5p3Ihd6BwF24w0p2WsolBkEZE5cnHmZdvsijd
u19qUv45sU3i2v2Y7dtzTT8C1EKXBJm+WUX0taYMUq56sSLiTzXy3h2pNvLuodDLOXPrqYEqH64E
FQX4PfPiZxA2z89zS40Ip00k02l+W8aqV1BYxOaRXzX55zjCWzq2H9N3P852/3wsIwgenVqWOb+k
EENT9YnLzE/GqGBxRB/sis639WYFqdqrrrWFy8M6RWKKjAUnou4jEi1OTaLhvrsv6hAF0rEY3Me9
Hh/ZObQUCSZBnT70vsewHex4ydPgAO9Iz0aDBd9tDPAMPIbxK5Lusmrb910+1dOiPx1vDW+6fEWj
aYJQTfLongwlOjqBe0A5gssFI1tKPSnY75v2RbSihgG+HATjBIdpBZG2TCk5LO8A0clJ8Xt9oHAn
8+ZSQZdYtrwu+l7FoWcR7K+36xQ+LVusgoDqhXo8mJ7wLJ8xu9oLu/HpvMOMmOBfFvEtLC5PDWyQ
EPGPCAXdJdGTW7nGWSGpvSlUrn6fxMkHMTkBMjveLL8VXynMFAQ0rqTDzJYXLWDQbxCS01xv0UzN
jbdhGo0kOCex1mjXgtTu+l0Tjgta2zGE+d0UZaTvmwXssAjBc+0tnxRNRgvOQOupHJDiFgjMRerF
WT3WrVHYzt1iA6+dQ/qj/UrCKziqErjsvXqgw8Hvc6iGhC42m7Yf8PFuydjva+YZ1mA5wuKxL45u
/Bn7m80rqFKq3MlbJ61uxMKC3s98pREf0KaTbmkh7VoaJ70G5Hf+Y2j6yQcNulEQ5il7L7WlLkId
EU7TOcUOBYgbxnl2s367zux7/Exp+8bcWmSuE884zjL7P23aXzCseduHCXNpLjvl/mbLHIz4b+Ig
b/HyjkMuE1zT9svhBzSkWJ/s36nLsSKaxeX9YCrIOeCiVYagvJsDQlJDFtiwcU/w6kvkRPjSiA1e
CQZKWi8O23DnzXl/3gUcfHjNntVO+61qwiMQH7QPxwrTxaYM/nXYrgScmtXBPH8YT8MiaEgwQA0G
58YVX2P5WzNoUUIIEaVHRR7ETltEoxkuE0DHUt7zKKQXb73Ws4nftOyeXADMK7S8UsHHFqRhKiY3
IlWEokDtH1/1+NhjwM9h9LZWRiOdoGkSV9KCRubWup41yDDKNWvK85cjRVMxwzn3QGsLSbMqE1LR
C94AUsflKp3szOHoQ6SghMGiLOYRW/uhPY3wWanBZtaF/kuxKY1KPRDE27JYn6drjFWtgKW6KRn7
pkLjR54D9/ofW2UWui1jKtU87UpdQuZUV0XDKC4bCYvGwyaM+ALcLBZaVxShUfINfLnh9YpbyZFD
/3vj83d2tGWAIG0GWXka2fLBeYCLNzHpFlKeF9/Jdl62r7ZhcVyMtzY3e8zi6J6f4gNnqXq0u37v
3MGd7ymuxlxpAVsJPDUBWJeScoGQT+yio327zfoyc2Mc/AJYG/R7yjBkIi2RHJbqxSF6cnUsmr/o
yY0GJyMEE3gPRLQElMDnK+duiiNnO8e1NVkaewkecOr6NoXE0IMHm6UvOzUs1rZ1k0QyRsfkmgHT
Q9TgaqgwEy8t0U6Cx5uelgDrmpM/4P9y5hvyvnwqO2GT1eXxxlH5nRaBtxxtvSK9RdMR88E3yBOM
tblzdXWFVAX6s8yJdedPe08YgNf4wKylwfZy6yTu6myq+l7ZO6gcxiBVJ1naW/kljcZetOSE6BQm
xevZRGIcMPtFUF2Dt/SwGTwduH43AmFAoZpk2Ohlp+k96xNHRXMoS0xvU4DkojbjWQvYRp9a9CJp
mB4jT9H+gRBjJWV8HkhG2Pmy0zfCfeYq3UX4i34Jl33OwPqdLiHz66xoJRfnrlGIpuSJjv+pwwRQ
t48y2HanfztgbPEY7jv4rWgPuoDgKs+1QDxLCYyB0UjdQ6c6yfNtibcirhJdXa7QY4cMHMPUVv4r
H3CNn8V00UKTIQq1rQ6prERR60VlDAZrAb2MOeUWpw6srJbOPzx3C5zBAHSyqy3x7QiMuAZX26Jd
UEAVksCihU+ZJbDZ69Xf6fl60MW5gMyj5DDZzGEm1ecDPca69CB0LpUFNGPFChouKwkE+6oNxiJb
PPuDSxXgY4w30OH+grd6wosypGWxHP3O91yvR1IRhs2BioknT2jiwnsTRmssSIhpx8ig2qNebZvO
W0HBrJhT4o8D3whjfZoMvBxWsVHU5cbPX9ZnmHqTk+YAGbl7D9CipPSAboGQdVzb+52+ui4d8kuB
Dw+bKVuMtvwX0NP+bmbZZ5JgK4y+FyP9/IMKUuSCKdWOi7Xvik0zuUmWjLNhqGJHqKkyzk+5AQPE
utxLXVEdgurfwlmHFU0V7cXFbdVkAq7Qt+A5n9VsCy6viNdtaAjY6zbQIxasu2IjllNjr8E4mLbM
1ExEv1dinXCzH7f7a3MJ0VPkwo4FjLNFfocHmOCsV5tgSPf4a3VjUmXw5LZ8eOcnTxd1AoayB4Yj
j5KHgd77U5WHte/uosG5M2y32Iwv2j8JjGCn+KiufdXYaoCLHIDWQGbwmL8uTjOXs3szAbUozfAO
f9GlZXAvHWmByJyznBecqHh7Wc/L5TjEXA+tCAQGm48fHBh6JXxZp2nT25qkt1UQ+R52cus96By/
eD818UO0QtRPgQYq4NS3XB//gwlTONgYn5U3N/9gwhZHcDskO5ksqTEcGz8ysMdfZMdxWbdlprnz
Ovdy4oC1ph3TlXvKFr9C1w/q8LUUME7jzFfy09cSh2xkECKi39VOjq2tjUv1iDIwn/ryN+JkTk0O
zc6/LWZyBpTmEIPTf8L37ymD7MBBc4CgigQYRl4jKksMI8dUj1cZVqNMizsL/7nxRkYdB21/SHAB
XbYNjIJ8dVzu/7Xaco1EymXvh6Hsm9SfgA5kKTUP1PR2XisJKzhQnWNIcBvzlUTRHHXjdxjwidNW
yidZaSTDYEH+Heyhud3e8XH4DRFqOs3V5iJHBDmP6fbzYY0NsB8RbRq+ZNsBcNSvemfMSW9EHT9S
S6RIbV+uc3pxhFAdoqDjr77bFmnft9HW0wvxxFAhbEii4frQ0LtE5hZQGjkmyITE7MuP3U/Sx09Z
3GzWwfn1d8JR+JGw8XrIFYdZVHRi+YR+q/UwCrOLCaImRYIenlBknDpbMOE3yY3hSbZ+gFuygBhc
08H+CUQ6/szXWGkSmpbP3IBAVpz8PaUApuxEKlX7fhrCFPO2eWgfbFaA93NOFdRvXBPnsg/jlyeM
gkAnGXSA3BnkeckUWpIaS6BFmzhDbpVO3RvCTJksLFslaCnSJG40o8ThASStCHAcG9AwJu7hp2om
8NIgfCgCz4LTnRcyps9mUylopa68ZvFbLk3HNXoIakce/p+TdEUHkllcCo8BfdHRLISkCa4n0FWJ
0hSNLZlI7XMAYUMfJaOGZG62cXhFIUv5pyoUtWqOpbHIw9DhnP6HFw72e0HKgcaNboqA9xdg36cY
JBqEgooaXkas5HTFRWU4B0a06BcLAJ0wuI21lsA9zutRMxY0ISLt9M/23++UkzsiFBUldPvcnceI
Nhuyo86TCLfnY0lBv1HM2YLhfu1zmbQa4eEY1DLOdPzMiX/s0CPErgtyg7hwh4lR6cZ2labsyvbc
v72tzfBYx/s5vMKKM8g0iWkoO68TL7XrPLqcZ8xFyjGb/QmQP95xXNM5KNjE7RDYsiesz+rnAQ7b
7iBcfigGOhF3Hptguvv31OuA2ym+sXLvelVdiOXR9dT3SL42xEFHQaBSa5MoWIVwx2dloOtrXIfH
lOg4yHGb5+EIpLado9cW/cU967V3WR8trLq5FJblJ7eJQwn6EdxT+bk69jA9tLjLLMiquwFmBq6V
vgGEuv60SvdBar+ECcpR7RmS+/q43KKOfqdWMxepKlfLullnFSexSK+YBSZNcsnK+3CD6FyQ7c4S
3vHwX+0x85Z/SxJ6mQbgJQH9JOnYPoYEFrfxciZsIn1EyqvB/VVgIZMHjANh/FR9J/YqswfQwoGa
uOwF8eM5uO2AoYJfaudaPdRAR20mtE8OApPmu6JAHzGMh3N7MhbJPgug7rvOqyLj4vHY0mt+ZE1Y
yKYMOZ9Q3NeVvrvcxbJGRSvNSkg/uVQVzW63m4/6rxwr+aKAngfFtaWGIyxzG6yWs3qjpED5EQVd
Un8p61Anfiy1dyFX7ZzO3XU1vCbYIjXf9yRysmZbZycnp8puC1y0R7nJg5zNgrY9eEsQTb8CzlIv
eTVtCq31s6rWcyvWM6yUf9Wvmt6/PG9RUtKchxuEdFhaue+SeZTrbFtfZXCLHaKIDNfhbxSIqW4q
8vHOWtn/mAPZPzJ/ywtYjbMg5P7/gHJ2K7YjIfLHOoHBUPDuczHAfASMefgBdIPZy37/2Q0adGK2
2M6kt8KVyir8yR6baYTur2nF2Y2Zf7SDrDfjeAp4UGfa01YueQORy2Hzs71hkqh73ec2f7mAKxbG
H1z2rqddl0H9nHn7najwLh0j064h4rVe/htoeSrptrsJhbB7oC45l9bw5Q84ErIb3mKOw/a/KuX2
L9qr9TU2l9gQVyHa+7fLDonwEC+2yC2TBQEgoIlcCrom4TDoBbR9gCEaDjyaRoalV9DrGrhuaTWj
SciEmazRfFoEyJMszx03L8JgXVmQI7UmyYsrY4i0nwhKKZJ92zoPAFBO0Otzl4qJ/YGueN9/AXCo
VNPGlZWJ8QRoJQpMYziwS/qCNn6Ap+RD7oGJhF3Pz1F3Ieel0WWN80Yc+RB5Q0lrolQNXdpexSRG
eePHkT4txz5RYajzM9HHheCGUCHTXmGC/lQnlKHuf+nH2CMWfyPxF1CDXx9MEPZjvNRrkHxhbm5E
PEYdNx2l/ksda4AFk1N33NxLKrXBvCv+Ipxda8Jz/syVu4+/lRjKOlYUJflB/XwHG72dZm5r75KE
EQ1F2jmS0iGv3nxi3Aupt1krPrmrHH9RpNAJflWfO4C0xnf1zN6j7rqTr22J5SPaLiQ+rtV0bXI9
cdLOZJTdnAB15w0Y03V16CZYMgkHs1++Hcqd7wwgHNspRbVa6yOjqDIiQcJLqPGshMbb3GgJgoGQ
X7UKH6WdjyX8U/VJEuFJgqaZI9WnJHCJwRTSacoPVZ5vSwctQk1pKNe2eMvVsb6UkU3vVXndBzzV
zUuawhwNX2B1v4gIFwO8Mbx+7+XJFs/LFxRVMtQR9xmUaIGNOtW+yg/So/WsdGa+87gbfEUQNISy
cBX54Mns0rsD1vNLfsiAlGauKdszpEHfhyM69cgJYzVwjNLQ75g9+0qVmQ0tiFq47BM4N4bHH8Qt
8ihH8STIV8JJvSDHs/YGpJaBORqiUk3v6kQq+ra5eG2hAk9ppfOYK9DHvG5Z7E4Ta5gI7ex+gLCv
sN7YL5nT2uJrkWqsJR5Hhl+uBf3xgXwIcVGJXRkS8YCEuuqu/fKv729gorwAmnfhM1XIzniMPiu4
daifBHXk8O7F59pobpqZ7rmMLj6jpKmXoVOo4zjXzB9DTRfQ4xHsO4z5QGVJoAu/1YQGnjYwDpNZ
Q1fJofs4wsxPK+z4k/47/emxFU+cnp62jsQMmrDku2Pd30angSWbC+JoNkysD4ddCBdqVLEUWHb+
oTUPpS/OqBbtcnH6iv9Ig1PEhBkjJDNdbn6j+ke42HlPajjZ7jFpOyddqSqvaQt4YSMtBtU7Wv0l
2uTNKp25NfHu2UiLzNOjnxQGOtdQaYnen7RvozQBobctOiYf7moWBQcF4yEgdZNzeggWZY5dlyzy
UbaSTTAj7i4lpp2LbR+Rb58HMN8/69nn/wbpW3Nw5K+fM6nYSJzF8q6MvgRmeGgl+c0kPaIfEZ3r
wtRB1TWiI2KNPi3CBQMcN4yUB3Nf1RjwO2SRXBkAwKD6GsjQt24ENWYTUR5JWFDeoSmUpc9SpcnK
y54kT9bMUoFtCVDtU7r/ehCKKw9JnskNZFbXUGr3WxR5sxH49OzdhHkXE1PgqGVeZzW942zGG7/F
8MF3pnu5VUFqLlEpVX33oam/04ZLMBycURH5nulOrjCwbbV81i3UvntNpYzVJejYdlW+7qYEFW0b
3tiitojBp48/8klGJh2WwOgn0wdQuhRvuNiBDdVFlsqyk7fIWVlOjrWDH4Ak1bHnzrXD099lS5Vq
AIgB5YVs7dP16TifBrrZTOT3KJJwN1ZeA7DHNnqKcKZ0tV+OJowaStF9qcERYjkuzI5Lmj6je+m3
9V6axpkOOIoWqQEBijGXiF9FS5dkZZ1Tku5smhwtLVoxRcfqmdYRf3zN+A88nymj081AKAjL/Wj3
X24VZF8sRcOrStDbL4E1snOEBlib5gne8FC021H1ewVZGvA+HYS1/t3XIW/xTKqZHLGprLGtIZuV
1oys9GNiUkMXxAWxqY4UqupH7GvENh8ygBv9fJTeiDczrMAw6DEzKC1BdHD7b7/RVuKIOlKh81/3
PL/36/AICRYkDVcL0SPB/PblgvnJSG4xoKhyOBKnqC0maeqsvZgGyhD9UiUIXapQJumMygA0Ychp
QqWE15qUYo6njANKEt+2XCF3B4LwvaV7iBPNSmJuDOHnpfZUKz6nFtKJffy6TGT/bfE7WDY1aqyg
39yM4HD3uuKWFuq7fq1zdMN3uPbYOWqqlxCL0w4jqIlTfDmXKOfcETIotH7jNNzCXb4ERDlyq6B6
JMSllP4/Wv4/9U5ZSYdf8/m8dMH+RPDqCKnJ9cRMxq0/4JVEGqdnDoAXVqTIJ02PtnhnZXYfPtu6
CRFDAvi3uz97zdyefEkaih3mfXclcTI51MZ57VhgvO16o7QFy/R9/0qealffhnanp8aT0cQel6cq
1jgveRB5pOZQd26VFy85pDMBVuNm/ET26211Zu+TKi6lWtRM3e/sVM5l/gSFUQYh1Y6UGaa0Z4EP
auSrWOPyGuGuRuYHOTPyU6jFFURfXytXwerCHZAg11IMMXwQo87BGhpiOez8mb9MiuUYwrlMRYeO
MJhL4biTMeDtMu2C7zBuMNcD3LSBPNCpC2WJ8ipgUFTh2DyxIuToKdtV6BPwl4W1n2dxvo2G1M1y
RA0OhUen+9gsR9OtEzjSzWJcneKQGMuNnKWLuz6u+uIZOkzl3LUcaGKdT78Bh/ED/pQw5MLMJu4+
puE9Y+Prt6uyaoYu0T6wzfjf4WZZ8QCCDx8Uy9m7366sDbwb0Tlz3bfFczp3KoIRReQ8tPwzui+5
1AbiW4/55DpcuUa7jm2FhxYyEyilwoL6n0/PAZ46c6MlTbBzkqH4XvcKtM67A63ODdnq4dCl2b/c
OPWVZWsjm81RL/mMubVhiM1TmG0mMwK036msJ1pyI9clmIhM7pemP5Y6hS0DDjkjXGMTeiKHrTOg
D42HIWL4GLtI2arj6Ajq+jdqsakKkPySp/cbu81nCTFvpGuUQm5AvVxqa5Myop7XOnWzU286gaK/
ZXhIUp37lxZaz775xGqeQuG05NYh6r9avdZVD5yf+nuzJYivBREhE95sczjdwr+t2cqpjoGxH2Ec
iYLBm9fgiH+2eWA6r7DiH+Jbpvm2YUv7kRMRAgDL+1ZGzp52TPAKaCJ9NbegkaWZKgbxKfGUdl4/
lekw1qP7pY96FMZFlqr8308AvINspvxbplyIAj5SmYIh+RCxYdn6AdrrCKdP1vcl4udXzxW/hs2k
MwG9QC2F0I+WU4HHUpjzfJBZteoDTSwrlzLzCvvv4SAGGid1zItz3GWutFKGo27TQTFuRyk5PY2H
eMswN+yeSb8FrUf1oS8QXRh1EJkaiUErxikeefMUaOYLawSGeWZIAw9tyv4tPbrATy4OOyzcnXs8
p2nyRtac509RgIQ8Tr+/JlAu7kwIK8j5P6fsOVTcg93kN4IHFYzXr1sPOx6k7uYu1Anc9LsPBzxv
Ija2wapPYATg9eBKhZ5tp/duIvO6LQGmqPFmZ8OTH9rDlSVJnv7Ujb9SQf3dZt/2twEzvQYyXWTL
n27GoZdBCNMwSWtLW1QNVjK79TewXSy3qrtg6xATkvOE+/gATGSsBYbXfEcQ1CBJ8NE4sGZQmHBx
OeHWT5t/SZHZZLn49BucX/WKciPlN4vH0zovWmsiVyiIOis1P/seArRW01vnufAqYlzBhzQjiJz5
NUmQrJ7moasbDJBjFd7IZFAvCBO5ezEUHA0ehO7K2YBcwBLGoLKrHGs1fvzJz1J0BBGkPP/nAU04
35F8andl6f4rSsFh1qPxljvYLmnuHVc4i32XVIco3CvkzPh8hjNozgXUgsBwKxQ6fae/B8vVqiCB
8jDPwguB/82ocGXuChLWZC+2XAW/Exlr+AJmv9IfbCptzlYBChfc/LLQ8SRoTK4i+TrgiuYebGvC
SRNlhZjSoZoYSI4AQWY/2YVR1QEAY33iydo6FA3psintLUgOPmVb8ow6TFdhhO22XidfsyquOtLi
kgq77NZl5HJAjRVyKCbv44ulN9OeKyoEaNhExFQQ76KavqHlSsn55Dvnyq0KrEWzD+Z+EueQlPtQ
OA6s9KcJVaizgbk/Bx/mUgmF9XntIsXVRyacgM9LaPx0UBZSOh08fc13vfnv2ysY2OsWVA+S3HfV
32vVrH1QHB2R1h/wHOif1qj6BYYinSJghHiO1NnQkyDxrUF1+4rzJFfL8Ey2Xfzcy095/g8ep92G
6XPhXd+zJbHcaCDPWKqh6/nItjN9X6bCXTA8HQntYnRB3kk/FRwczyV+0bSiPe0MagRdOaQtLNBJ
vDphSDAVMFSTsCdvPUHROKM1aPRHQnmIgglEh9HYxVF0u1pOTmCNr7rpYvzWmW+Z26mmg97jod7e
goC+SFj35diSft8dkopBUFqFiz/ufMGe1RBmFI9uryXe3Y7GuKLIrsH9kkamLcJ1kkOe9q2/JlnF
iHBPK6Xw+gW9yIuyJb3hnMpOsOJ/poXNoZS4Os2AEx9XxmSY571DU1PTv5+a9DM0RkLswiYvOrSu
c0bWx/OcmoD1ZOmSHCoHoWvQczAhwmQ4QzA0gdYxgllCJqQi4BDTbVkMd4cVpztQjk4Dnyd27NRs
RPAqCdpnOdXnsaQH5x0IXY66fbKyWTYRuBedVy86BriCnWKwr9w8HSFeyBy/dmCWl/NT4F1v71E3
zql8/ihOlQwaxkKEhSrHTlIZtgQzYVx5691TkTxc4JbIXcxw7cbU0YLQ78HNyJgTpJTTVXltmAYK
oIDdk3wMhyKLre49OxQ6eY6hUiQxR1MwaXVjTjA4iJ7gjrg+vIC55t0xfVCHDBYAQNuCeDYl0O6G
VdrH//l0kdTnGhKooplVZAnvk4AdgIqFrdQ+3fu9mupsliEXp5VpUTdybA7GEP395pGDZVcNHIKz
KnQSyTxxmXbLIqT12oxwkeCpUh8PTrn20WhLXsO8dW773jYDBJGL9iF+3vMvwgCa136XTKTbJ7Ww
F/ICpWk1T8lexwNTcE668B6zOZtJI8XViQqVAjOxOH8nNGCtjs4y/OFfZmfOKqSNFLF6QFSBsQhk
NN4Fhk6K1QiUDq/lqoDmPF5c7kBvU6K7I7+/uSrFELTfVVC2iDFfs8ftcODEBitygbrFBiESZW3m
Uaa7N8AaHw/+f2mCWgq9mP62HadV1KPrTeIQx8rLYg1RPgsnqmNL7dRJXWTLyuXagkXoh17SPM8n
VAI173jggK2SEtth/y0CW4cT9RoE3qWrZ2pIJo1rvANZmOwYeR1f6l/ODlfl9lQhwAjaUceRSNbl
BHY205XYNWBNcOAV6aMF3I7J8nobCm+RlpgtLiSFjIJ5Fyz0/PIt22f7fRSFrlJg9XFAtLLdghol
AkSOrY3hUXdu74YZ8OFxE8wn1UwGsTB4Tmli9wVgJfcY0XHMBS9rAKsHhwR4/xbaEnZjSw1foafs
5lplWS9PHVkmUPFbPc0uQyi+LX1i7ThmUQXD1jASYeq1duEJgbX4oh9LBRjbsBxT11UmO++VtGYR
bwzbqOzH5LxM9jWTqLrOUaeur1cJix3PC7XGpS97OwMAMXgygXwYCEqSCOP9NhyzJ2bZlsZgJ/+K
OmRsqnoJvcw+W4IWWvkuyjq+5IV/oqoqSS+FOPH+Fwylo/xuwGtYPFk+UWXChKrMF7AVxL/u0vOR
1iv3SqPYfxggpTcU9at0r7Tz4jZ1+5buZpJgTxTtFDmpCRqz0lCdY0+UtC/38OPSpeOr1DXatQfh
wKJdlFaD6J0MeDqF5A8tiMe0T/L4D3tSgdlHd/pa7BrEFWNpwXSvUkmKJHi66uvWWmzwG3J4orh9
NnuEu5HLvFbjRdhV5Alcb4Qaek+WCnRiqWsg4iG/9bjcfF1kh0tH5ZKycZG/HaJWBXHTt8LciSZ3
boTeIHCzoK6wPhjAcm74TA796tBS/bFk9p4YFB1U9WHvftnfbRtMwvLvU1yFVNVsU+Plv0PJvwcj
IQHjOFyqALA4FPPVqQuxbd27wH5p+z+BFUA9FoTWOnQvwkWUkGQ2l56wpEpmSJ7a8xoBSWJk8NI9
RjaPo2WqJqB5MGy90O/BqU78iDvHJoXMmqNgdjbpkUYFOdWyk+xnP4pbVfWxBC23DxzYG9GoNViP
WXL7c67PEwfEc75hKudmKHPDisTBBxI/BnzDS8fohX9UymdESda0WwyDM0XLETUgjKKdRRUoceVY
Z1MCCAOsk2f7K2lFjWcXMF7A31NSg0P84IKRZ3mKt1SL9tKHJd6m7F0CRGLLiQK/0bEnJPJwKuX7
JgDiXlhbDTMvEeGwHg1lGOz2wgYso4R2kiNDP0KOkBz9wecuzrY0LODEiF7YaKS2mlNWvB3kDgwT
SCyieZiMbFItQAwD9ur1sKIDTZDgAKPsQXjhkR1fT5jZz0b7u5mNAFcXLV3utraFAJblLE7fsOMD
QcWoZhCXV7td+hnSwuEIiRrJNNanRnYJb3g3EkQL6SkWreG0fkbnEUEGIAMFuhU+dzIHsETZzZ7J
r0Idh/AcfW6qSzG9oO3xkk0JEBfP9uWslgEnQVuqZOn3lTdYx8yuIJatQGTcxY9TByUFCytcEb5/
CiHcaW7+mXEDlPJUig1pCbF2k+zOlLJJaa1nPuSYVTeDuy1pj91KoR9YpOp4TVsriWmgaUuy6ygv
xvEDM5/9tQuOzXxY9bVT6QByjp5NzTlNDakDx1I3FSCRIVVI5MllGTy/r4fDZiklo3n1Wp4DYSBA
lzdw0mCo9LPB9c38aZbW/t7SZvSQ5Sf+HMs7yFdtOlnfuCrzfW+W55tU3kLttN5w08eqjDFpyq8k
fLUoOYnhpSnJcDPPuA4mfKRwdwKcw+hpZRD3C+1t66rSAst1xHmA7r+/f5fzrLqmHwIJ4Wk2/Ap4
6YP7zIb036Kk/LpAEeRi8da2m++QCFNDAPHcLyyZQZGU7Ot9nY8jCcIIiNNaO4IQGRvzjFPW9/z3
+XWnwwKimDI68/D9ZZIpkvtNGaxooeYqoGJEPveJiH/VLfij7dlTkRcLNuiQ2AUmdt3Eq/I232Ih
8OioHrVqechIi34+FGr7JVrzcta9WRDBPcyTrLwuLWa6AJDyFqe37jgNT/gQJIeVXusbTqLMzakf
hIR7tzMjzSudf2SFSv8BN3kRYNecHu3Qe/BGz83AstBuJO1jKn0VUgda2+GhdW9W7I0XioXnSMCH
n/XsUVvWcl6+Y2v4oy9TrulyoQgS2TgIG4fzlqQymKalNJEqu4q8sD/WoCWMqYE7YE9JOnNdiXVm
aHwBVUEKA0QnheYg07+rNd2qN7woZIEbPl5TiMN/4V8+Wy28+ezGR4pVuHt5/3uMo6AQnnVLBh2Z
cxS68oh53BMiGF6mos2qXF9OHFdLkbTJLj+LUCqoNHi4qb6Ictzgws+N12Mu++o5RrZ5jMm1hYEQ
akBY945vTtQjq2Nv9drIrqr3ntDwiisfG4Akn7E9iiscyXbUyThkoaBgCc6AlyMjcpXUhdjdHFAM
3+6itMo7ywxdD426r1mIvzXBxVKcfwGSXvdF/TlBfcn3OuPsCmdatHmDnzhWjmTl+hvqkes3gkX4
Do27Yk6tWOCdIrYTgtFn23lthE/d/OksFbCH3y5xV2zeezVdwB32n/pE8SKD0i9ma0yXgs9B42sa
EmX8HSxHLDjt6fQpX4JOrJI4EpAZINkpnkIkFUVBuhp/My3RYndAUil8Y5cCS0ngBU2Pn4YiIqUl
5fQ8v47ZKMWM2pIshe5InHNmj241Rl8C6ir+dZtfcpnXRs9V2GM8be4vv1tO2qP7FOIPu7Qwx/3x
pqnLgGgh2M11nJuZqKvwwOYy2AxkEHKbGyJGR5LO2tJZvIIx5XX8bJ0KKhqGFIAVE9rMOMp1Spjw
2xmxUmTqBP032P+SQKXWvhjRAQm5LXeoWgcVQ6cTDdak3uTITQre2HmFcbUPeE9XefklMUKAi7jJ
1sd5JoNOdggFDjx77YC1RaZaoy80p7cSFyX3mKJ9m1ApmTH9KpvkgOOwvAPNIKdbPhSOy3IlAMfX
dV7fNUA1ANzV1FWhP0cGgjMUh3zA74GxC9a35uZpKiicmujWcwkDi1Weqevuu0TfAEUIjFiSl62G
QrtoWKPDJgXoxQvLwQWELwHrTraJoPPt0VK74hKBaj7l3E7eI6gD4aJLFuQ42lFGTN8WsOB9sZIY
9cb8rtcuROZuSLsZmnvhgLaytv8PPW9i5tlXq8H+ccwUr01PXLnT32ua7/54Fi9AahYGipBkRtnT
5zy10FHYuLPsEsi6JOnHTKrNWnj/X+uaOclGqjvtDCJ02kMezNFGv+zTp+HvcCmGZvnceCIPhXwO
mpFLF0XSqN9Pk9Z8WkW93N2MOqJSqXQWve1sLvEUQpvqunAgpjSRLIEYExCxnHyV1yF7rk5gvCKM
mOPIG0W5itDcBHib1kyj7Az18NaddJJw83RKz3xZSQ27ooVFH92xpf/CNUlKQ9J7U70IccWD9k00
xxwqNuK/Ltvbutv6S54mrAj2Er9JWF/fAC/mLG0OHqfaOHGZlGpJ5lXRmYGSCfmOy5cgb1K6VfzY
Fgqz3eE3rlaXe6wtTlTUMlH+6DhrfAnLHbMQ0RFzFp1DYlBJEUfxdKUC4AFMsH6Z6lBOsiXNLtKH
8xvoCsUffuV6n3/0uHOMCMvsfMYabF5S+2WO94zmgrvUsYPu7cICV0/j9NANU3XbkCXWZiDD41SI
jYMcUJw+4+Fj8HQs2+tVVbQVXjfK1Bin7NeWDGru2DsL3r/bUycgvLmVnOGp3Ewi2l38ZUF/eHar
3GAUtXhRczMRF6pL6X74kV0Om3jh7jBBVZbFgMTXuj7vOPLLccSF2wQFYwfEsdtopuTp1sz9Y66N
s+Rs51eccG6iYY/+l2v6UYrShA/Z8cpEwhF1HwgKRP5kEb9jJ1EkRjb9Y31m0ZCM5hnGdyTd7orq
Ai5qGUPWqCqZTjx/HVDWlhdPggjtg6WTZTN8YOBBEOmn2kR6D6sRB7YvHBGu2XYOi2FHhAqgffgz
FlI+T1+mtnSvWS4tNNeZkGLgtC4PIBEd4GArHPkfzL9SV2vTrJ+5lsoHPalfXzvXURnmyzPbniyf
f286m5ZmrRXDUtCZbGOr36S58+r9SyOMUqEmJRpVyGpg4yAt8a7oSG9aKxZa3PciM+zAwYnR/Qre
W0cfUbCAUITkVvSSmQ2iVeYFqGgpouk42T5Zsi2i7gPhIyMegOzeMxLzgGMwOZrvuQ8KDmwx6216
KvaXz/cwYNpHhyr2vVQ9P4Ow2Q6gE5aKFCYsFDEiE5vh46M5gZ7lIZOVBQsahKmTRquxxCpekmWI
r03UWB/eB+QCazXhhUmKXSAFHAC2oYm/ovH+Ava4KSQcHP9Oxv9EkC6PDwGim2Zyf2FQjbzKVKuW
6bmR0vI9Qs3Pjfidko1r+ywsbHziZpNJe8MXQSU06ifJy1Ut1kA/CcRjPo8bvGV/EnrS0KQMfdrx
b5z3V0GaUTLCFEX57fGw8MOH3KaM1322hceUNdBnTitjE0TDQS4qQ3YHwl5dvFVPlrSYCKOxzZCk
8YTl94oqeZeOMwfESxTiq7z65NtlqJv6wU6j7+7IL25X2IlNf/tY+QxgqP6GNR0L0sXu6fB5MGog
Uu0i3/0oEzfyrZSXE1LlJUbfq+kaXu1R5KSjio2ZLRODf4rIm1oGX3ShAa2HxIgVTNDgESLvwwb9
makp4Ac8jo4NZzgk1Mq+BVbV2T0h+HuHzZAU5/OCZjR8DMj7RK8aYq3YBQkrGnhVqhuKIgqY0kwv
v0fea4pizdmq0reDoNd440JR/h5ptuqhPRPAv0f7kXnNrUmyaHt8uf1bzkz5K/ccwSzT9zf6iPVI
fHE5R/Up5mnESqhPgPr5bGYAIGLXxZfjyzFgoJ+hQ8jvltiOsxG9yxjYVU7kurGNNJuRImMSkhbM
mVHXZK/wGNwriPc95mqmT5X4WoJrzZSm+zRV05iZqKG1KemUV1yWwpIGKdQsjWiA0YuqEfTiXZrA
jfKPwJWU0udoIH0RvlWB22ev7AHg6s7zLo5ajlGizfZCrbu3T20ThtrHonYrlvEjdKEuZv1lR4Ia
m8tXU7Yb9/qAb+/e4gcfaou8VV6CgzaYSqTr/FFXG/v1aDIGeKROr1V9q3TmnTnRIJtxRIrbB8DR
j3KGkPDc7T/67BkewNxzKYhTZhRImpKwbm5E3EXouqx5/ZIbjDCU/0fqqKGA1axf6JWuNxLLBAos
GGf93mnnLc/+fHXRSAlqA8xHDiSBdqzOzhYLCTQshZadMBW09znpBgvRS1psEoKtrUVkWlpEURqf
B1ELX/eC6TdBuqut+7jm7lzylbKydSJCQq/DliVrejDb3+SNnonTN3buchq2RyOL86L6YvQaxB6c
hf3TTXn0qBXpTaOKcIHPov3NaHtG43Sy8dvMTZnFkRBW5kUFLBUYXT7PmG9zEUZtdu5z9Ykj92pk
L6HHBut/2rNyChTVWW2n9mNYFWPGudmjsdDVwZZaH4nDX0Gcb3UPY6agy3hHwmWANb4wd6+k607c
/vOiclv3SQjhiWSRaP8AgnCDWUzhdExYoLUJ6ZdhiPwbZFZDQyc7TkT0/f9yB5rOyrxw8xQr6sIu
l6uRqbXx5xR4+2QqiL0zNKZPoJEDlYEMFo7h3oVa9AvZ63Via19rZMVgttn/ibfkK6k5OvX+7qOu
HnjhC/4o+TEEQss1YBUuOUdvu30g+i7XRJwSRdV3wy68iRHmLxeFczQAeULxeLZ54jmBHuCeydRf
GtyLqMkoHIChvWp8IR6rt9ZfqWlNIxTxKikyQb7AGX67jTWANx2Pk7X42ucYBEA2l69Cx54SPjSP
8uweGWQQccwokDCFt/eUWJlDWLadrF0S4+1v3EwfRv+2xEFfaokUih4uFPpbx72yIuKHRYUkaL69
bIwFIHV8KjJb+U6AQbhtwv39keofIN10l7pSNvAmFM2Utqb4a90VOQU/DGReo4ZvX0nQxKHkyloD
LsMcthc0rffUSKHQwPTe4fDDvv93ACeZtc5ZX9TS6fC6NuqO3WV3lTT/h010DtxcgG4S1/Wb8xlN
wtxdBjWyOFhj5PxAOgCyZsAEJovlk2ma5XFlPKVCyJ7O+dU5WxFtPO0V0+hyAUt1tYIsiS/+Y1Hx
Xj4HWcaee0vn/ub03qUxf4FJmey/uPIP3zz3VBTZuCeTrkxWJFO+qq1XVNGAnpxXXJx8m3V6WUYk
DX4l2ciBrPTMXQFXA8qSsbomllYfdmGf7J1SDI6jMtUyHbq2HFzflKUEM2YFfvscf6/yMgfHxuhg
hOzwFjbJdrZELmta/j9ix+Z4TiKIkPERiWlEcOmsBMOixw/jNQS77hTyKV8TBX7bb5T1pFkzkjhM
DnBpvHmgIXBvPHIAP3+9nFeLjh/XvGlovHxVZv8ha4BdSMBs9lz93rbK+8qAY5LUl+1R8LFrEoic
1NR2Bd5RKvSxB8aUFLGmz2FdQS28PMmSyMkLyvS9Ev+zfVTDwbNw3jNNBlTzMrLmDFF458QeSif+
87zVW80R5o9jH9QsUXP3zrHtlQE7AaDU1j+rrAX/1uBmbF1BOmnB8wzzF/1O+OonjZWM7mJOgzZX
Cs/4xNRY38NkcGS8PV60u5WNl0kN7zvHNLN26DY1S7UDVQ2wgTBBuyBqrRNF6hHpINoTv7Wt4lCz
X6XqGt87orrBONMNmXOjdIWy8NvQ7+5+hXu6uGOfeXedxcn1LrRXhwaxdKNv/5OfLvrmMOXprLJa
Z7fmIMu7TnedWEVOBLtEJtiO+q5ihwStg8nMBtr0jTt6fovpR0D0pNoM4aeovOoxYvsqOOOlk4Qm
Nk28eJ9mKtJxkxpagwQMEm+ZFQ8lHs/g09piQxusEdgsUG36dJlRuOf8BM99pQRK2iYsPVq+c7OL
JSDW09QyEeqT7REkIBJRma3AE9Sjpqni1bJUuTu/2ityEdFZuI54oi4s6XlPUMowC+FhvdyHtsCU
TcUpCLNEzVST1JQQvecpxTVwF2MOp0aL5L8hxomKNV+DPBsKMq9WK9OgLDOVZN6PpAa7PC4sfbvH
AWKs5MzDvRiVRIOgcJ/UBy1Q56TZNHmiq0gOKpkObV1ZiGUNWB3Od7b827kgug9jCIhAsmDpxapx
gQn5x8f1r9vWPmGAyetFu24Dr61xvQJCj3fMzHFgjaDJnG8bYm1q97F/DGyjEPN3Snn37TIx9v8W
TJydsOdRQppFrkU4zVVvMFeHjO7qRcWEt/v0pSR+6ld6m3vBb/G2RboD5Geo03zarAolojum2Pqx
Tk7ykgleepsC0WpjkXujc3modUSxkEyNcpbDnvrRNuyjEM8WGPXa8Dt4zutGLVVIrIDmhj+mmILY
zljRRH0bxLDUMsqq+Z4jRH/u6ahOMeAfNv/r0iO2hixYChKQ7RhfiYVkqwHlsTLRXjd+doPmyZTx
iZURDggVPrpAAEjlQMKSQL0nj46R/KUebtvBRlhzH14VmdX5xaao8NCDDUDlt7BD3i0JohxH3Bfv
Gaup3/RW8moILKm61NLzLBTM9pNKxFBceHD4HoMEFKViKzYWHZ/WG/1V4/vCGtziNebmgLKVSn/e
ZBkK1JG8Z9Rt5HVqzbvdRktXIGU0SujjT8DqRXf08k+g6+40pYSDfBbs9gT4WfbuNg/ZvgkB9hrL
dUbpNtDdemMV1mYhic1L+od1TUb4BN7pnVSMLrCkicAMyzWbR5PpZoRY+GBK9usfeSLNv1q2ge2p
SL5T34euQ7opPz3mz2Nlt7oQDTMC8bDrjfOcWpTDw/6V0KDzYXuPnhWqQf+xuBF0PlAhoCQ/0O3U
HCTS9RQgBFMhk6+B0t1iZnlnAFxaQCANlWUQCA5XVCLaQLOAbhpHNw5G1a5VYxCcqzv22K/TcYGK
UK8uNdHpmHr1UyUOrTKIzbW9LaKdn7a3CvzGREg9ycSi5UEjsidqZy472BiWfrC/dPzd3Tx0xBi5
NXnbiA+XHvMUkNdb3te5UXR1Qd/BMF+Nj7SftVToEEvFZp8QBHJei9TR3atjFJmsUEdoXlcmnH0s
cinIO3SIxxpjDBL2z8viLPwwru9vBvmOpn6tOQ8daq6aJ9AsrcXQ7LEM2glQRToqHZ8OEHJNLT7E
oJjSj6mdA90S9r4hBsKp7OOc8Vrh4VRslJBZ8osx7OB3e0g4dbCYabrbM2VqSSWKYh6dmAKQbdDV
ty4bAPbw1KvcZstfKE0ZOhseSUGlqE7DNaAaRakIbt1JXcwYp1IUNq+IwjaCMKhg9DUYSklpV78X
XIV9N42qGcCmW0C/3HQqeTLkocx+60n3zsS7Ac/eFTFk8fucFS1Um3k9gey6euumy99BwZ9t58Pz
WcXVZm5DWI1PgwlPuAG5tNgkDEkziEjRbebIgc1zxJ9Mbaj464+jsW1c0fSrCbd4qGUX7uSmeVf5
Thi7pCJoKc00WeX5AVguedkUVvz+KYen7zqElGSmGOOpk0LIKLd0NxPr+nSRAyBt3pIm1I/L+9R4
FgEzmkfL+v3+CiN2x55gSipCxp8uQz4W1nGGM91WC5yMCjNnA2f14+KWA/WM2NgSMbbMZg/B6oVw
Mk9h5kNNUHRfmPa8Rhv2U/iSMucxx54DVeIoIswhwjNG/eZp675yxml1kTyHkJ6NzWcW82+6ubIt
TUW6diVQc57Mx1Zyz0KV2WIg29gOFA8yrTqCYjGD5ro8x+gutRcMUgpWds1s7FGYuUnDJNHHpWbS
cY/oO7i/TNOLg/HZpb7UNQK/fCyC9LBcGkrPZ9sUDIJusrgkBIuLgaQhy8AouevyndxEOm7gKD01
I0F901TvpHQm4m9LHjaTK2NwG9qvRpfF998+AvTjkuhVbbCeo7snphogz92zx84P7pIqXs8a9Hg9
FHpZG1Kvf9p0Me3Ir6Z1JYv9BG9G6rQN+pwLEiydqYfs5aIPqFO0IAEXJf2XwhcdZ9AyaPMlGiZS
J01T71H1Ss8AS/GVE6TNCcP2DTLVBYHDNOxv8Lz0CISEA1Sl/M7tcLuS2enASvqETTLrZKYoO6L0
UAYrL80wz3pKdGrFK3wCs2+dYWBYBbDLUcy69Trdhv9TKdYYaeOZvxRWR6kdmWD7ctk6SeD1fIQ/
829T9HpXvhAtlmkauRoIx84DZSlLgnqniQpwhc/nCvpyDqkZjwLoOmfVA1Z251XMbwqf1BkRKj7P
6TqkqtOsckNRnPdHwtdyr5pmgL+V/20INA+kFbzDMWmuCif4XuDG3zoAclwGpsITVAaDbryBa7KC
W3U5zm1ifnfCxqC9bnMCeHDZQU3VGCCOpGC73ybURG32Lb2Ib7L7SUc+o/FZex8AiVOL4xvkJDQp
1AA6i2DJDD2+rO1NuDyWoPyAcUy2rW6HddxEVHrsBSmkneGzDbXzIqAr9EKuXKvpOmag2VicRkuO
QDJ9DCUDcvvRRlAxKnfcjbRNkTISo0hki0kFpYNf2F+OKmLpzBbz8FL+6YIZB+zmSDvdPi46GuTv
FqyCOdkarkKFPoD9Uz1+YK5PuUuIZqCl/kjF07t+EUlMEVFPTq4r8xzMwdkpFFLo/WPpHb+SUYUL
MUkYBI/bx2oYhiWDxvMpIBNU8KvN51eViefdRzxXlEN1MKUQ/16nNJ9z+JjnbW6JEq/NvKJmMAtf
G2hp7Wh3dUS25VJ7DtFS0qVxO0o4BgrPUMXPzklDXmKxnMDeZgNHq4EXdnC30Ql2dp5rahb7Scde
Jr5iKYJXE6/mP5T8qhMdlT77Jm2WEa7nIQtehA2dm0S7eVFpkhehmVrF3zUPt++irGkNha+hypdG
vhUdE46GqbIIG/zg/VVFVBbjQVkU6fMexMrX+iQ2mXpnwyhBdwI+bTfYeMwPqfj1nVZgTNbklFzK
s3+h7JGxwkL4ioKEnqFdvMrEautuevrzTCNs9rkSeL5jZtzU8O6lp2ZUPQd9hE+ZFkEBU3US4PBA
uaB7PAKFo4tWToIWRRYZVDpsRvVjXIZjUWLkZqDIOQ2zjuHowL7IIyilD2hVaeaQx6L2fA7Ub4TS
XWTdLDejZBW8iSFdqnWjeollwnAy1a9cyxgHL0jSc1s74aH4QJ/vwmO38wEoTjDiYdzGWSFXc5sK
JC9aw3FJc0B8jUuA3gx2SWoSKylN/9tdtvxeQ2niXHyUkUUel2B5/Tv/xLXR5Hnk3YKZOiPg8J82
nqAIJciwsbxuv2169mD4o9/K5PxrkRnFmyQAppvliQGHabB3wUCjEFFgM2U28JDzdX1a/pWoz0He
lbw3ETn7isWUlXmbsKFjeDVKYpKoTugQtnRqmZnqccDYCWltOMsV1GvExnUEeCSHwSLZ4p5HZ4Yh
LJXetM8nqsoVc+7BH1ZwA+zMs1t4uieXQg86ABLi9ssh02UXlAJyFE93UsSXpi3iWiHY8+cjweQ4
messQUN+xKIiY2QgiGms3fOvkQ2Wl2YRn8+it0T/VJ7tlhAnp9qWuItN24KOUSQc59KlNmt50pRK
X88DR0H8lVeCgPsf6qMS03U02O4GpHe+27px3Ou1I3h5Ny95ydc1Jc2QboZsSonl3yDmT5Nfncjo
nhYtJEHD99NfVAk/wQL+H7QGMTWhIHbkp3/pjBX90YIIoewj0WuPr0XlWbaulX9lNyXfr3qyWDJ0
rwffclUVaB/1zaXwbVBw1nll3pq1JHMxsnXYCfq2MsmspDnS6u/74e8vtUHa0JBzA4ZoC4fyRzjH
SQXjGrpv2umHKrsMBhRZ+utoPWyImxJ72sgg3qTullj8npwl0bPRcDm7j9YIfIpdkFD9APYu+8vN
f/4lH33GNCDoS4LxdEAi8oWL3eevCqRYut9/cazomQmX7HzDrLcillNBHxZMFVRglIX8sx2ohRLt
/HknnDgVvE8m1sa//Bkl9NLtOQ2iAG5xBY3XfYuEjC3uNuOw+UKz6F5FbFKw/K+5bCoao4+G0pUn
OEFzf1Yx5Otm43Vd9wqkckO1dAkVaVwfV9qELyj9a2ymJZAKmbfFPjdFjRgNzmN9kAR0nI1ig/7m
fafw/RUuC6DCFzbV9OuBcVRg5b2KUo6fXqkzX2/Ik4UzU41QvCHN+7+yHRIXYGbW7tZdKth1les2
pdZdfjpNJjCPrVBokEI/6+58xXjrv6sUf/OtHTyUT+aYv3hyyb+LHUsFnuaPWz5BnukjL54lhfdU
M07wiiGmDhABlHldaelO3x4gN3hlkn1nKMOZ7GsWlPQurVrO4xnclJBcrL6oOLcv13QmuuoSolZt
Hqw3Pb9+lDXjqZ2u5lTfd33Rl7DkAdn/Nigl06Nr0oCa3FpOvjHvHbrWot+6PqsvpALFojcPtyE8
CopojoU3P1FZlG0jnpSxtHGOFjReUvO1NCBG3e1StuideaEdrUUDoCyjj31Cw3FdZeJVbgGt4enP
66KJ2BmY7DxYpeHrR+hxKctcrMwRCplYLTqLDm/a4iIqSnwhDRLl9iEcGbN/9wj0/BLi4j4mmkLP
otTl4UcZQVw84rKNpihkJItRlhqyowiaQyagyQ6YfP1BGq31ogbeZZUxBVwFJPc9xIl6a2wV/qDU
p+CfB8QhR1Zj9nucOwEkwlENbs3JYEjHBHoARdHlGWwWJK1qU2r/UJGDWJCcSJwh19/QR0EvnCWg
tu5ZXbJSbqvy/h0fe6qXk5LBJ4FT+C0SvdQafDmWpkOyvRBKMgWLPiaOeNgT8cxzVLzRS9DjsdPA
9Ldu7DZ24tKZIl7MERpKO0jqg7/60nrQe3P8/fPlm6RbPCYj2K5ZA50+4r6l5kY2w3ta9noZ9SKr
XsoyRRFjdOKJIeStpSxX2BZHdcr9N12PEC+wo4pZlWLcgMBHg2bY/TMrtnVL4jXWkoxOJnVqR83F
2fC4DeHISCm6LpXFQHBtpBb3PAODBEa9cmsN8z0+esreUPRIHzA9UqLFy5bsPO/BgFDnm6Fk1w5J
AeEM5x7Mq3nVOcUDosjizRkL/bkFcc/U3nFQ3pE9xZb1V7GG4+62lT9+kKW0qx1T5BVETQkjTmPs
jqvS/71IL+CBQFpR7LlTpO4vqDUP94kuxb+Owq9kXitXObpbnU9wi2zYPAZ5reS8qtbPvmGjQPCH
3u9emO5337p56Zh97AwD/ux3XqdRZSzZ4+/and61xI5C5PcT0O7c/haNsNLOfyn239DuJtDBdQdx
As18iljy9lGRnSZ/+5PYO/SKcPlo/l08WootqECx9W2csylQW+zh/5RnpwToH+T93OQTeVDhVHcW
DNipD955SbNzf1OyWVgmnaPlppRlrjnrOrrKZecT8q7pDqleTO67/31fpdE3j6nUKtTtXi2yNsv0
F/+gV3CSkFS4A7nFebSz4DPoOmhlDNRNTD+c5scb7REldBTS78CMP1OaiW0UyqgYQ9ho6hM3tSMv
N/5RFUeTk18zJRb2bk8++6cxbDAXrebRSQUHwL0M8W381C8nj/RiuFVTd2RwDZs+ilCVf1f5gcb2
+Yt5zeoboQKfgWe7m2aek0aiDTxBPj740ny8tS/A7lYMFOLOQNpVHzSDp85HBF/LOHks9xko9kDX
Zv39yIg4LN+BOQvapPoaCDIISnSGXCv1FMvtMz2S0WqcFLC7kpV38CkbHjxTA/NwN6iDgOhk9jMq
1qrlvvxNz+JpZhx/qQ+jdPSs58SAnUbWJYJzZQeW7e4xNzsnlmdMETVDYdc9SZaHfye9KU6EGosm
LAiRlen+ubp3T76V+i/2uP3CXO/U18rLuTbIPF+MsV5rggoCWqDz9Z1zogB57FBKzWX+6Pg7dz+U
xdxC+KBeuXctZOfnwmyJprFqMhfZ3eFpw1SjZrvVTBnabYYOPn+hHKwAnOhczPOJ9CzhT1UlDLG2
qiCtwLO+FtjEgICOHs+kYhuhNQsn0k0+zPeQKUEZRd1PSE1LJio7BzuUFtdkss28EUt8kRBXMmnG
c4BGYjlT0Hq8anAfVCts69cC75ATujUBBo4WecSGZMiXg454zww09h75pKBsyNS9O4rWfFvtHlHP
l2CSHgsrhOxQYvs2uacOTqk8fxy/LfYpQiIjRSzL7UJmn8lBY2pnYTaO6RmeZpR6L22Q1U1MZVz+
G5cs2uw78Yz+M2gYainf70EcMTHRFatZ6WgR+oN8eEZr192igzPPnNWQX1X1h2KX5r0D2hRp0Cmy
MbehfWLbJBrcS2rY2wfT4BfEgfq2hEpOOe+pjRTjOqdBHII4ZQrf9GrFTu6a3+JjGXmlj0RfiDgK
JP5Rv2MivXrZh3wEu0ICrWhjKsGAF1DqMPt/XsmEm6w1FZcg6na2RQH1tx4u9qlfKl9VajBdZoM3
YzvM91r6LeKPC4wsJbVXYy+0I+UajBXIu8inycdIto4AMRhav/dlMJeDCrm85eaoTTObc33HvqfD
llz/CQMN5OmCvE5zOsxkx686Ry9+PM0/92cYGE7Xvs5w27+3AYlvWDMLXOecGGzRwI2insy0vQOR
7OdT2lZ/Ad9KzMT2W5ZGGLJ7dJckkVD53HQFUa4wSLSMOtesS6C+EvuW/m6Mu6cC5wWt3Wx6Y3TF
nU5hI8JAgBP7/DDVpngJg8HKQEsMhbX3d+dwJYFf9wdeps95ikf7+FMt+tHOuyO9kCXmFesCchop
y4UkpNyeQ06Wz4Ed2JWZPxCsMQMHhpykHSIxhzve5iJXbfvIfIOq7GI5WPsfEDED09lMT4bQQZkI
J14E+nnHlEDzya/vLQxiKicwFdNFxibpLI0FE5EsF2RitFu7YkK3H8mdFh8ndvig6TmZ8hqY4JWK
d6EeUaQVO1yVFgrELmHyNFoXrJP47ha/Q+FMs6PNKoeOQjj3wk6xOYC1LqZIy1fU+GVGLNLUvCx6
26ZM29py3LAkFurMT6CMm6zDGAx6xqPwF7MDl/m5QIn1ja8eULfl45Ogo8cgWZdgiBxVK7uBqX7+
wA9aGzbpgVsl0OPVF4k87BOaNESOa3JwlQh5NotRnSPRFJJfx42sxN1gDXVr3BK3AlO6i0aNyUDK
ai6O4j5V3nSeu5DNtprPPXa0ViOU1vF/69RY3BcoO35L9A5iVVuaI8zP2duFoMJaCjhsO9jzcYp+
+95o4YgoN+FERzw9rxWoQ9kyrHXOdbqpCzTD00+9boSwkk6REIctjISFFGloPf6SgFovrYS+Dg7N
utSi2gV3gQvdqQ6cj7/Kc00V47mjnxBoC7pJLghCV9HhYlMSkWmPUlX8fkXssG8ia72+GPKyAd3O
Gix6hZF2s48OBz1YsGA9qZpts48vV9b0LATJaeZkotFnt1w8zyeVZmOen3yt4gny1wspuJ/I2Z7Y
Sg/XH44D0RkW7TSvfTPg3zZWuPi5m/WMbHCAspHGWfru/ZawbTQCDVYF9cy6xSydjNs67srRHUbM
fdG6zNdvBAmlgRridMbJ2xbkPLlQh1hhyBcRZ2+Ll/uADWtNKFLwiI7Gx3H4JmHu2SklyHGYj3n2
vk4ZEVxmqIWVt/Ns8ytIw+yz3zxWc8e2eswLjgK8JZtC0UEdI1l0kjvUfY2ntfvOrYAfo+ChIxU2
0/7qoOYkQ22vtpJnwjdgNv4zN7RZ+vyFqfp2XzSKpmFnNsAaPTJ5QPwc8rukUk8dvWYwb03lUcW0
+5OomsdCXirhtwXsBwPADFnk9SU7jYC8EarSoYkAxwpr6FYDY7ko0QeFhzrpEd6CAJ+2psXiLhRX
5tQYq0qoOfeqTrKm0xuUn8voGCcLA3oWJBIdWG9Zkx5V4oVEbAixfKPSrYnWR5Cd+x2MS/vEHoev
k3B8YN3QQ2r+T/8d1FwbfrYMdAhq4oErpBjNPZKWDMAyWWigPKIlbN/IAhoqF5NJt4S1iJjwU61R
2WJKevkNBKRGoqEpcDZFV8fhGk0/vdgyQJg1xFcHABCG35suIVJJKYxh3+UYLTJBTeVaGRObqJ44
7ARtqjCZjtT3ffa/EYg6bov+A+oQrDauDp9mwC49tEnx9TB8mp8MfmCHyTNwefY3MrHHtvgtvq7P
zCGFk/BF7BUkfZWadpm7/sEQiofLcfzn2AFvWGCYtBoNtjeYNC+ZdRyWJKP5B9QY65tYc+rWKOuz
mV8jRvqLV9uSfIXWgroGZzn5uLhs+rSF6lqFmpLeUSb5pg1DvNAVw5cDn+f3kCVRjB3BEEaPde4T
kalywri5hYlXgrB9xWR62twv2wJecbOZQYOVoH14CzC2GnCWCnzJBMBjz1dOWrJFnEMK8ANKo4LS
jPZTUuZmaNi/bPvbi3NCgLG2SsZnoixWR4ApOeZAhpu4Sv0eiaWjTwRmjiKBiuw6M5Pw1eLrBHwn
3moJ0ONhLPgFPdpa6CBrsvMobaNJZ913GsHCPw9GN/GOEtUTphwplxIMM/RFRJbBy5DHY/IAJti3
HrNd/UNNOpi48pwWmOV5OBxJiq7T7ioHYjOZrFfkZxCHFpD97z4rZmne+Eb7b49Aco+t2dLD9YSz
hKhvagowNQF6GmwaHV46q8KCnU/81mINL6Et4fsvx5fO+HVScY7obwiuif8roRqjJRvZQ+0pIN9b
Fg9YRGqxNf4IUWGStwkQJkNYDpNo7nKUJplbOo2HOiAoxXB4n4zfhKo115Z8KvIkrxsAotVHY5oW
dmaX5+iiM464A0/rGyyDzA3h6y0yvEIW4FXIp/hCVgjdpV2xKqKGWtB48pmGNlrI4YIpkqdrpGHh
xUaf3bOywYzNo0ji9dQftADM7y/byyf3yGI4Puh5aaceeD77A6JeIHNanvW3Zs/ZgNlfm3yW+3U0
UF2sETHM0UVkEu111XD/0O21rz/BMnotqC+4POjUiNuaV3E0CuNc2zcejR4xLOSbdGrsWwrkTNx3
sPmfUBd9S4l21RmfjPKJedrqC+zlcLDm6KzYkUSQ+KazfmHfJfUFM1273GNjSHKzqKqNOvYjH76p
mIW1bOBokcKXeEytQJhgi7/aNzdStLVV4V76a+ITRxKdQds3GmZmrh/LZnLJnZdJtAd6+yibFUv3
mAYs2r/rou+7VCyXFU+rGogkAXm2dwrFgFK3hD8NtsblUhKR06CfB+FFiCxsnwx4tpWIsLUPugcN
s1nv6Ay/iALWdPF/ZtklT7oUjOAsAB4UFH7I/dqO2kSnOlvseyIkKYdiRfsjvQ8dkoVjuT3ZzBjT
LXWEs5ojY1wIwCKJKe+GTa4zPmbwfbms0rJ87Bo3D2ZMgqeIVFiUtU++p7QfTZ6vQS7JjNuHqJRZ
QmAr1fdoHVl4U562DnX4VHOx35PdNN1ghPiNYnzc+T00Hvu9E7kNU45V5Y6eXRFgZwKY+eMf7FPL
/O9WrjuuWPqZLmXIOJAixNd21OjrehFWGqwGLKBUdN++iouSp68O2sH/EvscPQsluTQcDLj74hf/
JJTzMgTT2Ciw7miRCEXTp4SLLfk1mLMSwCCt/lxEyzGI+mAVD3c+ooujYYtYos8e822fnlK0Zn8H
T2GX9TNQxVBcFvZT7Hjj05KEY/bRrLGuWvWjsNDFUsl8mmqjzCSi6GiMgkpr1yPbOzFORlIno8Cb
Jc1iTAS+Xd8YpIb1hV84T7BApbTHCXNqodw2h/aBCY0YkPsy2RPfFmJ/Xt6gH0LmCbV3H6SmOlYz
Dg8k9WcmbqS3jltZ9LsUVPR4yLyvaKL9l9utusbjQGch/6h7BhNEdSVBepk4dAi1aouJZnMoWuoM
jcwGaXuyEeJFlgdEa/fWARX52g8oaYkOAaHq1ofGvIGebMePPkBKQOWLH2PULFHIzpoQtciolPdx
hIZclRHerOfyAvSnNpIvQyI5KEbYGxTBbyeYlLp9PTQKHTEhXoYyC2K9Ezqe6lkLyKO7Coai8rih
Uym8D2t0Tz6/Yi6H1cOCGGfix2xEwCyIozydxnTUn8AQdqTd8nw6P4By0934FtC2Ap3BguGvPeqv
PzzCdlfL5uncs8w7ZS9RaLX7/l2A7eer13FabSylZKYqWB5Yn8z8/ENHICrjGNjs4QDtQ1RFoQQS
651sTfTpGeoqTSqmviWayMZLoXy2Wk9ACxD573O5Tq8sw1KL7YOjJBTaH6sTCvqVaSEUPreFpjkj
/cHGUh4odTHfO2vmvNektdj48DOXEVFKCzd/H4bRMxNoKymLHwozgaX4VI805HrfP3WBa2IUpQ0e
7jZ6oA80pS4yFzJbb4W8HCwLDRZaJAX/AW91oxEVVfKrgdvOgMsEWOWN7cJlV9xZx9qOV0u3y2J5
qVJecBZB+dAdpiB42AFXb7br8rDpmqoiFp0wp9RvuCtJHy7rzINwNEQt2vAkosgomGk5EzrUwNHM
eYoZgyNWyVJv5WwDUYsJmOS8LlV4auVdFgm4QrIngwc+K+80Uo2mrsApnfRI/CqUMFfBjiwLouPD
Pq6h89tKJCnYmMfQ6QpGmIfaysVG/BtaV61ZhOwEzrS8ugHtQ9y+/hylWuvmI9Ca3e6/5+BNmGwR
fzkysOG8+n3Stv0ozp9/mQCB1SdF3EyENovyykiaSzWn8KkBBYlSCcgJNBthOEvBBWNbFKj+7zvv
ShkU3j+pcHBR3vQQO9j4eKWzKSYbvmwzz/avcU1dcFcEaUN8gQOQBeqOw62h9qC80asmD6KEY9/w
ubw6cIglKlKBYo/x8F0yjmWdiQJDHdH6wFZFkGXZ4j9jqZdQ72+KslTsllRaEbZL0s4zK2o2kXkI
Oy8+jw2gXU8Lm/MqxX028rNE5XJ4iYAordjP1nXlPJYALlnhmgN9Bqeqz0KDaYnBwa0rwXFlqbz0
tvtYDuMI78jXldrGWfd9ScQVjnbDXL2eqE1suRPyz6iMH7ER/wIuW2jxZiLXTmCnYwsY5P/vEc1s
aFHnik96M3Oag1Vh44eP7jQewQW4mGcVfeJ1aiDrN4ujy//ePnNVzfSF3nbleXRPvFef6oKX8f0h
t1JzA2IotOlWVGUdGnygcQz4bjXi8lpXDLJHiWV/asR/QIloWCuz6oC8K2VVwPqBvrcxqLiY3Tro
E6dCgrwAHcqtbWLVACEyb+2lUO7It26JS5i3R2wviSBbg+pho5dVEemTC5ynyrITAjrCU51cd6yz
aGJinMta8vxGB4tBVg6ZYUI1Gp2Zgw4aoFJZNduSUyuwC7v82fP5N4DYYwD8IprI8bmOCJXOgdSU
kunJUsP1X6Wo50nK2ky1cAyo55htsUZ1C0u3FvWT8smiMqU2dM7qN9Fkp+YAlC0Vmhwsp03dkHUB
rrvknPW11ErmcjdfGUSlvIEpODxM9MbMh86+zP5HhBf/CI8KBcIVPF2AX/L16/YA1G8QoiQc9CEa
xW9TNkpIOCJxZ6KvMGHb3prRFfEQW0PJzf+JACHXsMxxS282DZusLhRYFTDW3mquhIQfKEJ4NDjt
IOAtubHkma+xOXRs/DqekouxbqzwpCgwleOj7CM2uVpUkTD2d3YdYHgvkx60E7jig++FwgHgRoGD
F/cvOWD3xkQrcR97Bj4vvhnKkHhxjYkmMdPCMnabCsLzdrQ6fU4vt6Qh/rxr+Xtu7nCf86Acrsr/
WfvBqTEAVlk29vPMnvDrnKhy11madhDlIcgwCiL66ar53BWaT2rysg8wW24TpP9dR77dMW6hEl7+
fkyoVqI3/P/QA65XWAviVw2RJ6B7X/48cvPQ8J5J+aJXUJuEy7Do3ydIhbPzJlK5hvLB+73CYODx
GpIq1kWXo0idgC1yNDYsL5hUCH4ZuwjdlnsgjpQis31BzbWC2yAG/5F+/OybZQl7y1CgK5oLyS32
916+5M4ziUO1lZBECrA4eJbdElD01zTLo4qoqJ3vBqNI5b2bB9VcPJqf64P3KlWr/5i1pf5NkrSw
OUcs3MQcdCW78D/t7k4oAygZneU3qMMAtCpR/bHKPaMHDxpgLsXObwQ/Fmi451M=
`protect end_protected

