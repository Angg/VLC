

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
aEqvcre4Lyvq+Tt5PXDTwx71ktTXYMy4x/0E4dKe9BgxVOReq4m528LoaLIP6GW+fVGwy018LBOH
jm1+bivxEA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
QYrPCp2aMIlbBfuPNfY2dUNw4w+QKreq1bwTmXohDVK/xUEdLBItloqXSCGC7+jUg/Qb5I85f/Ah
KtJEJyCziwj6IUpMayW9odpLYrmaGSusKTx06OZfHHMO82exXNzudcAn72ELL03w+v3J7Rw16Yaz
qLJy0R/MjFA4OGOwuMs=


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
WY4Zr5cvsgwcIO/1W7ZGRcuOPxuu6EPbRD5e9/HsVO16X368aWkQR33DvIRaKE6mu6z2j0ahwjZs
reKraTCWpXPIX3kHEOQ4G+U8/pfBNAeLu+gHRaqilAs+vw9yv9whz81+ixVCKNNcRWQOTvo30pDu
skLTcm2m/QQjNLEpHtQ=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
m6613vAd4+Ikpmzvgk61cQ3LztOi3BEUS+a/u62stTAr62ac1zeSm3L/nrHzan4UzFg0iiv0fkQI
HlLvWFQnraEvQEyI3HNvXjW3i1zg2bQV+yu1q5XCIXhmGlzOkz2w70qM5ze4T5v98BsjMp4dYmMx
A5f4dpYgpZiFnTGLeMS7ck0fB2IZjiquePTdi7jgm/IG+qLBUBUT8dNiDp8GCdQcgG4HweV/m/jI
vG3z9EfAXam/6EPH8epbQzdWAIlMPFNElVQWIXYwEK7n7IkwPHcKKy8h8TIQQBgfI3+K1o6wVERE
QWtvGEQ9KskjsTu85uDfcWnHbHjSbT9CjOWhQQ==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
akC0NqgvB/U73AVdpjoyhrtNQqSO1F1f7/iM28U3ok7yrD2+mcT2y/A9xisbQ06qgSdVkeeZQ/fM
UEmZFdpeZP65dH8ladxkyOXEBZxMn5HBR6Cc/cxzHpMOCwyqreDrscOV//dRgt/fMDUdAzVx9xAF
S3wPRW/FXBzvZQSBlmnr30bFT/LL4Cj8vJGIP0+tX4O1SFvZ4wHGKlU5KqTKs8dVxLyBzSJGBQVb
pymfPPn1F6nJ0s221XFfFykuFYfHfCrSyu+wvMs87eFK5xuSJUkyXUmL+AeodntlACtqvxNeG53J
I6QuD4FQzVWl4npAqVztFXpihv43QWWvfcc+3g==


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
SbRxC27qGffCE5dqvP2lAKXlQLXs2E8yapa9AwWyA+r636Hw6fp2hwwnmJLYUQJzK+qMT7z/eV8Y
OxzIIxbpnjsdHYaEBRYqwROlVe6YwnZ7L6xK5KKxX53MhhFuBHhAxWp9i8Abwj6PqlCffSngelnZ
dnsX8SbNI4PN4MqYSBwgphTtKUTWu1vfLq7rTdNhmsL/7y528gK8mIQQ5SkILrzE8DHO+vA0WuoB
gDK05L8J22kNnh053JxW/y8ZxHFerifahlKocYNdeEgc4mj1EWLlwOKC3M4lBgZJ7fZnJl1veWSN
xU8ddBWIU09TNJJQCC3Tzn/0bh/v6jX6rkbLQw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13264)
`protect data_block
nOcTRlqPcoNBkT5B1lUJpZZFV4narJ6etMCEGmQpWuI3bN4l7C/KVyS0FxaT1Xa79WUUTgKqVw0c
PfkF7sZw2h+RbhmHR7cR17Mq2hLUtmgszvjpo/t7kZ6hlA+SwNvdLMQ4Bzam0fhpjWNdJPuGyhca
IfYpxvtaobo0dByOXnsSlEsNqU6J1pudLc2VUgCg9G/umr8AihAUOtY/O5bxS84RizjpKmdS9BCS
6DJ9tQF8wK4VMKgPEi9aBc4v6C6MJvpnN19DHwz6wKLMDpbjB0YHUkL0Jx5Tps5QPPoD/2sKrQZO
HGLEEIRSa38Km+9H9MMXzOq1VQG7Jdb+rLruUkLcCVwq8do+AI2JRZgQd80gGvhvAvaD93MTENXZ
FzMc+4pbtPEAStv+gXmo0Gw+EQ2LKvgmAkoHUD20ZToFoIedd0Z89BLqXMeaUCZeXSsIvukqxnyj
fr4X62O/cNWK+EagjWEHlsqEJhBWN3r6HCikhEwc0A5xa2EWYxV59xZr+jjJX3PWESbP+PxUY1Pt
u9tzAFzDbopRNuQqIEiCoEEnW9gP4gzBge9YBqISh+gUj2y308aq4pchO7L+oMeViuJDhg6OBqpp
hltDz3P0124jn7jSom6tBKZZpHlgqvCGBpLRpGXH9qGAk1EqBYQYklZbPrvcNEQOCAM/sH3NODfP
RaqzCQWdy9LXvostlEHFr89TB32HF1yetGpafLP3+1HIJEY83fFxLmqheTQJ7Y1FZDdVRt1HD7uL
CYhuyc6WsgqCJSv6Bi15Ia2tI/fU6O3Lfag+1HdBwOo3KVdsYPT3h6UC9qmk+F25SqPFNyDLA4Z7
/U7UKHib4Msc1fmPtux+qdPzhtW7/YuAmOg3gTmoTjwSKRRknwYvbkOIzgVwBYy26rEIn3VHrOes
uBaCUDPwlWXW8H1l20bj3AyhrU8Ztb0BDVNfH3orLtzg+jOcjN08H/OOs1ZQm9Z8arFQdPnU/2/N
fWiPwYqe8ZiTaxYyNQgP/uU7yIbmsMlpHmZF7P0Svlg2LufOKCZi6P6fJSJa5k6JTQklIwywU7qy
YikDcQIcgmJ7byHsfurRd+fNG0IAkJ/gLdTs+RvLHCSeS1m8AjR6FVl8hrh+qwRANTul15C1bzVZ
rWF4863fYCSp9HY8c7mJAfbPIPzsj+sXoWMeDewAUrUOQolqOOV3xgaqAXOLy5SDRu+pw4UTD8kf
fz0PUsLrznR+2ISNjVpwmADPKI+fGmaXBdIdZTUccKSntip9ztegGiTWyxSEChc7EniViEOVuBre
o1TxatzsViMihMkEc0uxXniJ2ch6AWA4Nta8Mvl9xgMWW+KtFYhpsAeY+UZ1nvLkEe6mYrEHRbGI
RhD7aRRFY8uC1BDYB+ZfYHhp77alACR8ZVh1d3b3BpLMgwHXh4sW84x8elFIW4gwGK1BbtQ2wpMa
M/g+cwSyJv17qHPYIJF+HkXGlvt5OIx0DH2DiPmtTgLRWY4fTJp9qJBiXo6P30z/niHh5As9qkBo
kbAFG9SoqRndoRdg+atFPMTfd9vBWcO+6vOEcd5WWlT/EEyL0a5wHPgkrlXoOovBcSg6BGKlVOb/
BTW0NFXj1UUUb1ZoB1a9NezQN+Ln37YoHHDnfPvS+3a7G7iV2ZLWmOk38qgavUJ7JEbBUXUHwNGe
W87Z95jK2Ggs0t2yV8L6UemsVyHUV/sKnR3sNAOGMi9stN4Lb3qYPoyMKFszYwHfqvqRGi8WFRHt
i9QTM0HMefHpsZvhXanhp8I7exBWrYslZe6FoN3VDwhWCPM4KIjY0WBpZSAXjigxXPI/Lbflndqr
/ljfjUY11W2dKQRKdO0Q/xdv9axg7VpB+mj4caDuVVZu/yflDvvgKGt8fe2IXIrcFpKerq6+ciUl
q115ER+PVnrOpwR6Xf4QmcmtYlz7RrYmrBsfdwvkfBXi+xITEO2P6Qe/XmKBhyLhid480PrQTMBj
u0uFhE7n/NcTp1xPeDqqScKdUqvUuTz1q9WnHLdex0/vw1B8JCmMIqVZ0yADLCs6gtkgLwKNPOQo
L0y4VYAtZrwckUWLm0BJX1VOIHjhbbwQtND/fR3mVTy4PQhjM/phFk1Z6JUVBnXcnVzZ96PiYYFy
2plFsmqc2pFeo7MF9OriSV7C/2CTE/NGXV3jmOoUlI10BLrBa8VsUWtaL51fk9DKYYpJor4aGnNo
Ts3gh6MjXlau+37kElz3bmh5R8ec4EO6gaxMHPTfVBgpyFf4asS1SG3vXHdNxwF/hZkXxXl+xCJW
rBxwj7bA2qrYqd/2aZ8wI9MVODgqbWCUbViryYKPuBJArg8ehrdHGGwtZNVXdZ+Amz0e2PlrxIxJ
nlB2ONcro/3NKXMpmYYu51Z4J2f/UrUnnZcK1ntLNQ6Fxvh7NkUIxd0R1Wq1YJxC/8DKjmesjhPH
DlJynOlSCvYHTvkssHc8YBTjmLmdhP0qJAnFSEGdUpKSOpcHfoVf7+Q1D3AfP2xJeqg2W5VAsnKm
sEkjZ/743Gv18jxjMKPhGl4/tiHQN4pADo250xfcMHWqglaU5I4JRD8e1DkCUHZvPF8Gq456D2mF
7rF09BU9vaO852SgSnlfTXl4BcknibwtvNA0AWhI0+vEuoRp2Hr9GGlGUNyyAilTsS5MA3oTw/XW
kBJ88LGo4Q4owml0kBiNelePSLaoLg+rNgbwO072vz61AjLc3QanMGdP1/vVSfI2fGCUJvzg+TS/
hDBCnfDYBYW6R+KQ7sgWDWxe+MoZsAbJPCfXjzwp1d1axNU8/36baw3JcIDim1QN5FjjUqCDOCVA
7hXYR87yrLsR4VVCQeMDAOkH5234pxNHuS/4bVqbovox7+TfK+xl1EvO84oQxDqsHH/vqEgT5HGu
O0uw0A0P3n2I6LOFQxNCFqCDgC0Frqf4Wk5nu2i11nyrdYo7jwzt/rHRNVdT92iz7877nRWpqMJV
QfYrl/xKspG8z8Xx0ZKEIFXGE3VVLd9j4kDT3+l9vn4FEW/qgrufp0qFoYJTxuAtP/zUFqAQPH9q
nr+qMY/NO6Jzfe4BgNT1k/kDG9hnFKFJeZQqEAckIQSS6qoyyJ9c+kPixhtD3gPDce5MescQ9TnF
UhG7YX52zcM/IuagtqEypO7ys7EYn6/AWwmWTBZ8YTLCkq8VqSSTCc4Uya/KUMWJYD4xmfVfVkYI
mVI/8/4tw7otUlCUPlgLMphQDuQLprdHqV5WwOhoYkl8LBB9GKBy/E2lcfRI/WQktZdutzqEZrKO
MunNRXVNI1CUB7lOUrRSXpOWXGJHAJQpi0+u7+8BbF8hHlxuZzIJFYF8b9SpTIcZ3zkAd442yiel
yi3AVv31afNDToN0cRyh3hF1nIVuwvrruXXcxmbRGOG4rmVLQm/Eg6+rp6RtISrqbz4uSAOyq4yz
ihWR2EsN3Ny93Ao7Svpn+/TgiGHnj536vUyMg+5qfadjT1RyTxDiYziodbowPnsj1G5qPNeSwaEQ
avzTIcAPVJIn9scuLlOsnRSN2UUf1+Qpi9uwcYEWdIEKDRNomoPJpXzGwMpJMUWma1GDY7gElr3L
7bIDK9sW+gel1G1vpBEFLdpQWHUa7PFrRSFNe8xkc4EUfwbfKkEQgfrhkHjTdQEqasLR+HciLYDp
1w3DNHptXXHqyxYjUCAaQUXbD7zzex1QHLJwKLDN36XG/3a0S30/qB3cw1lW/FfUgMmb8P73+N8x
zEj4ZH5BnPiwbKoqdSgmHAwu1X6bgoAdHWIf2ZElHPrUGLOuSAYvn+zMqYbycuUdAqzPTiUJf1Nn
ff8BCuleTdPzCSeHZ+zFM+Q6jvLcHbLXCAKe7oGvcrTIE+H9soGJtlKQunH+JAZXaWHDpksAvk8/
QP+XrA5HweiF6lraWpeb78Dgj4aSbKIOVduXpM5E2dpYI8gZUMl70sRbqJQVrSrWqtFNZVgiQv92
ySVunMkm+1vMluZ5N2KP9RVBW/NFHhfXD2/fe2wPMPcWzk94NIvaCU351j4zMN0ctIS9aDTYXdSL
xyfmAL7YDV08fPCuUPfnAQDgki0jQdI7yijZDaPwnIWyGNHXGbIEZ1ASi9+dLqConiLdzlmmXUA0
KdyeGFpNSOKGhxIueVCP4jH54Js8yjl6KmD99vulCIGDCFePp5Fi86BZBZSpqbbsGO94fLMpYmwg
6PqJjRuoi9s00xJiMmvhfqGE8uFOoP/dJht1ZbdoSeQcLLFbrfLuEhlnRkKVjhR2/3hrspE4DLld
BDe+hXrkqycNERIUPZUY4P4U6HXfYXnB+uEoa0dbR1MutZZrw3XXI6tOMW2gtd9PINfHAYfvGX3/
m75awa5pTV/qv3TR0jezkU4WHnA6ghAUnKbUx6ac9JUAcTfvVRzVjMPCeVj9UwcZBVX+Olfr52pL
5IxuGPAizEO9T76fdW5F2iP9yyf2uFgZvOYxGvY9dwYzNDbPUDJIGDgrEYes6fdpuWBNBD1ohDVI
dzS8vsAqCmsNJpRxySJhhFm0sHA3f+o/PN2mdwTXbGgcxvw58sX4O6y50TA57m+6mOJSXzDWTK0t
bIv6ZaTYpbi7r0vO74L1yaVc6WrdbbyNxwm9daPezAa1b6z41SI3f2GsvS4SdhmOZ/1WJlOKoFDD
t6QGR9666ChnHysvFEIIK6rGCAXgU8U+cTmtqAqDt24v5lL06VJNW/9s7yQ21DUMnoRasMffCuUh
LanPXt9xtRdS2C95TqCKaFX6Qohc0BXPFe+Gw7gx3iCurpVWh1P39gsjj2XCiWvfhRCRE4mP0cWU
adKF97d6+Bt+vE03FGPBGuOwyN8ROo8QEVzRoNRNtblptyiPCUj+i3yYMUYis+5bVUa1JeIXntk4
0qI8YFxfBuvoSpU9dYf/Bf1d3GALbEwu/z/jomdRlxBArGK4gHAWmOGDOABDtcNMtRsHiArPiP0g
5tbP3Z+lgg/VoId4MuSdm2SvL2LIpN99yRGpFKcHNkmZ/JkBqJp5tSfTtz0Nr+jsUC3I4oATfzAM
/WwIX0e1ya/s3AaJgGDQ3ld1Vj3rXXHCDKG6NROO4eMDWKeB/N5QHm6GULgHojjpkuHFPilE/iWb
p06mhNcABLxCSnF625eX8u+VyGVxKhSanjmoEplSieFFiMHyJ/2ssTOn5nDnQuBO5eYNJBz10A8Q
7V4r3vy4B8eyJtXJ0dP0ws4T/KpOLaA2h/8yqT8vAcCIyZgTAEr41oUDzejiSW5uuRPA6r7iDvKm
nlY88sKI20gYtC5SGn3iAdlwK9JQ1PRIN6pzOKjYm7XFaWVb1cHA9OV+697wtjJ3PlCP77qZ+FJL
PFnxaFE2n2MyYe5s4cm9Wz0SghjnDq0/pkdJw2wC/unPG6QrXoa7qbB//5cITerahAesFwSyNr+A
tiSyMkiRMf+seAUh4PZdIEi12NgFwWv6dz6ymaGql0SPjojZd1afqzBZby5exMcMF1Ej6YFGzFzX
Q1R9K6xuOu+bel/yDXi58PrsbhV52oax2qhYzxa5uiRK+u9uxN5hWYLIaVhX3oMsLa+92NgE02Pl
OLYiZ79tL0dvbxMxYro2wvWhWYGRJTXLkplJzLIicBi8CTLUzQkKUjkmc/ODvtw9xLCn4cv2wjYx
hXvofUDJ61vo8TCOGiLAKyGQek1KJASApB1oNSIYmmFbGCbrzNMo1DKTvagWLaA8YxFOd40kVLOt
ALQlI0RP8w/weWK6JUQapY8eD6bBuaFpYUqs7I23S7CwMUupKM4R3oVptVqg9ALAc4Yh5AkgffSR
ncnLMvJbNy6zTa0kOFN13KLVkueV4pDMxNXpmONnV21XoRSkK92JgNVx/AUNe8CjdDmTyhdvYTVO
GA4Y/G+VOG95X2LcCgKDzonaWVdy39FflXQIcmiuvdK9Qoypyj3vpbuatIA8f39sJelacUQuP1Ly
cwvb7pxjF43KTd7xZzWmitSbTTeKmS4WlIwIeHJo+Kkf6ZTba6mz9RZPK8bRojGWxl2EeFxSYQfP
wHVizhfJiPDXBpFIao5Ad8cr8cK2j0ZLHqZp7w4kwXJ/0NpjJn+KeYebKLLUdPiyvK0nxMrHbuEQ
VwBQqadHHFMy+ujNBwc4vl7rnWiHi2IP4PuJGULlvtjKjQhUOO2A1jaKmL608In9+E816fdFlEZn
Pq9X8e7sXjDt3AQFXRqNuDoD5rGE4DsOhDn/RXc5TSAPaG14O98F01YUsqiIc9Lce4gAwgmgLV7o
ZUI6i8doZdAj84KQCn1va2KrtpDN2AZQGxAgvb4tbXTpdNJ6T+NPMcL6S428HI2iGyJqvjXKMBFW
JCQGcaeLbhGX1wbb9jtKag8VWLqkMTbTQf79SHJkVQvzaQgAmjRly2S7p5yiINBZbao2IlCz5XE1
kUpnjm9mEfVyDWPfEErvG6q45vIJ9S437ZROdbYTWNSASO46fN+JIVf0TkHomvXUxBiu8OFETrpd
seLG99puBswi/7SHk8JwG9lKjO+XEdyZl/ouaZZaiwvsLnid/lBMY75bzNKwOo3/4Zye4WzPiTNN
/w5XbsyFo7EOZKc+fI0YAEdwz3wnYcr9vpNKUjYGopTKhXGP1xI+fEHRkOHJTQoLCkUMVCOD30+F
DH/nHjgDSZIHbZtTRQRJD+vWVxb8cBEL1UcD1ltCv7Qtjr1mgggzSGhgBKNbDA9DWOCWvmhOUaaW
p9i9Mu//q/2oeOdY9fTYxabUlTqhIuoJg/e4xVQjBavyIKBtpdnjAYRZwqFQW8j8OL+BMv150rjT
LuLQdmQEtUxshwYPOiKYOHpSsxuUt3wpCcYTVQMw9h2DJHlwCHkUfgi6XH9cjSgWiK8A/vXlc2Jf
Jss83/My+YSLxv44cjoMqip8HuV0gI7DRE2/WbivNVBqi/Qcg5dfSrWGKDLo1F96FHJfZgdadgMA
uwkqSPDSxTeJeTLIi8BAmTifxDwrxoSoltU3ozJiodYPmbNMf0ZCBQPcM4wHoabt/Pl5JZ2D5kip
et+a21y3IrXB2A6R1FjU/ML9l1yicA54Lpk3FV2E8cbcXuIcdG2rBLuQ8FPRkzZ3KFkcCPvrWP1T
4JjkNcMUbYVLp6PsWYOdMz3uysR3B5xbz6UykzTgs4wXHYcLl9yiNwALJVzQBBNJKd6v7g03PQLg
zIeKY19fbrsD5/P3NyeY6irSaRkL940ZuwWm/00GWfYiWXmTAssh05QRIY+q9kPNEThBjSafhGsj
o8fYaEIWJKjGSkXEDfdqEPpJz0sI60+sf4pJxHLiafI5ZAQ+AajGSsskQiEcWQ5VXIMYISU9lsnx
2vs2oJpgtnrBJ9cjzbMi+lr2PaLfLaVFXDeQil+9sMsugtLEi4fPnvBYCbSusT5eKDvRteeNe2zD
fCAuMXcJXmJO4Pv6xi7JLY1VJgXUrled5whx1aHg2PmoqclnP/VWlbEORKQzc41uL28dUm4fpC5L
P1GhwfD0kh4+Ae2DE7RQNAuDipLMkQPfIRcxaXqMhTebtfTg4zBQXIORhdyHOz8jfJ54loJI3GXK
zvMD4KJ3yVAVCpugnhdKTDolGP06akIiqXg78zRgACV+xLcN0ULsGzJ2BEusmKKVU8qmGBRdfIem
kPZhNWxEotSkAHr9636z3j/wMIMQTYrDrKIJb2OS9Hcn3uyoDz5fjNgQVDTZeSz3LdS2Sc8p+DO1
5CV/NdcvSQCeEM3jgMEZQc1jkf8RBVI1bxRE3cY8QjRvyg4R3woJWnwsgXvvjOgC+xM/K4QlKllO
siZN70XEeUhUx0+hTl9YeVOR5krjL2cuMPUrqgDI0BdSwkPnvEaEd5EIFVH1tbNJX1+NdFYjEy9v
+Cub0DjFdGXIqXqyfuxDszlxIWE7dxWMlK+WiyUA3ciFJMABoX0gmBUR+I/KTmxY77nddzkaYZcW
JgmxY4obY+WZqZrgchCInpAmrQ3z5YSB1n+I2KAOPZh8zVvakqAhptpFekgB/zt6ri/PGs7esdTG
pQsBnie3uGYQH4Ki4ztFV+toPY70Rkl/VkzBjGZmaGioC+iZ5VMmX+fMcVhNiW4+YG6VyGMqWRXq
H1E6sPoUPs4kmQvZQbwB8vD5v8yj3Jqr3J8djIl6EvVPqVQltUFyx9WDlp4ySLazmKn1P1WAatmi
LaJAvoxpxSbfBwQAyl3J2ULNAJ5tkImEEp65OSdnTgWY9tEzd5D95bHrkjR+LdC9NyKLN3XaOeFf
oR1ZVNOX++mqVcXkoa6gCqz8we6BVy5ZtrcKZd6eCQrjPF5fqqIKagwn0cm5IPo4n4FLJvCnhmdG
mfkdhmKraaSkzzrt7NyEbSj+BOCE+VFJhxIxnueaS3vzyQhSRZdB79BnzD050KB7v4RPpgaV+JSU
CqTZEFouBDzIHXi3/OhHMEv1LQYVpCCC52aejq+yTBQR9thLxMNHcitBQ3O0wcp1WGurVXNVhUpy
N/PBaMy0rBAYrzU0Z/ahQQH0KQ+L5FsW5J8/UCw0JSMBt2Ooec8lLh86DiqW1O1JMe6mHT6znEwH
038NqRaY3PMPcC8VQr846H0N7IoIV6MoKGcXL1tojP4Ggyr7e0HZm6FARfN93dp784uP8FTLTnE3
tJD/+zh1PoKPZDDqiaSj/7qD0X3oqNoOQQb1w/GGYLt8viV9QhVNOYrs1mrfgeCDe7WCkyrEreO0
S629ggc+/H0vupzo5VS2ah3hVKcVpjQJntcrlKxhV+0PoVBli3L7oHmW2LX/I5V5BQbKCAyT2yCA
gP8pUkiDmAakKVTBVS57hYILY8gMFpn5K/x1y8H3CJXxpeKXXrY0q1kEoY9eqLBnL8cmFIhDzFiu
+16dgGzM2GMpmL6f5Z2EAu+i3Vmk4TpW5vqmz42azC+Kvly1sPIz/jZuDEFXcDHFll8x6+VG5/z/
m2hlCqL1aNtnLZJogdRIzXz44VOk4R4bQ7TFjUscFab5yU3ImnwiYPhfMDyx3Lhv/tgTEpAu03V8
Xa2/mMz+6X1102YjAWRXC0TphgtY2mkc1wrO5B7xiihlXKJrFkFU0f3IPy83tN/9oyGpgvUxrFHd
lTN3RIXaaG11Z/mTh0zFPDMCms7y+R19sbIDncy5c/epuYu1lBaFwW3czcJ2X5xXcI2cxXI+4yae
Nf6kr+mewFoy/9z9OjZpHmvWhNv08g5Rp3yIEeZN8/NjF/9JaMRgSvEsyVw/u8U3VD1I8+1GR1vW
Z+K5a1RfynkzZ7dl8Lt0oorK+oqxvVyAEtbX4tJkiLmmuNAvP0tQryVxAnNq0mNrJBXIJZAMLtKf
UUncjNFHBj0oJp0nXt3xvMmWzNA3aWr6ub+vhMJKpy2t/buO9JHS9oRgMO4if8IKO6H7goa651C3
SwJdTo4ZMcX1liiVLprfO06SMZ3+yp2DvImlfc7EkBrU10ebdwt0fS6j+Z3eSsD1ipq6PlNV606k
7xImH9ao4ZRDu0+vyhUNVk8vUZCyBMvEpdCZcN3yEfmxRSWhop6RguSNhFZXeAyV96ZWeuVXVAYv
8gJilzK2O40XFRUFYH0wu75DY+yEtmL0QmRrFc65wdVgXVPz5Q+ByjAiwYitG30rjcFuJXhxO2Xp
h9wd7L5A6spKc4c5aTJIhklVgMzJNMvmBMpq4g+Wcna6jOxLrux5l5rxddQBfbFLb+mGyMS+80wV
u/KC+G8MbcNHwKp2xEiraxZ7vagGozoEN1rzl1NaTKp2YsANQ6cCTdiGhXVdXtuIXjZxVvU9ePkU
2JmtxVPR+YIm8HvEW/tG6ICAk9QltbZ4rrc73v5t6k4Z7zXtLU2g7U5kmHdV5aeDTbEwpU1uNwgc
M/uSeu2a0r+L8pMPV88PqjAO234UJ1YSvCxlm6/qriMLpEky/QksyDQbiNTPcM2dhPiHkHb9A7C8
l3U15HCXNMeAdumOYP3doYb6OO5jd7O0baLKrAkgwYwMRWBxPxfR7+pYrQWM1oaL4fXFwHgToV6u
stRG6lOg/xFmaQacEmVgzz8hz2rqvdNorIKHVjTJF5Nb/YfOwYNyBAkZ2uJ17GqQnWHIcLmlYWDs
E8QZ1naE7pP6j7WhRWuX47y9EoFwkUB0Zm8hwU+pawdrGUNqhQ72KCUuO5gSR/7n5xnlOHTv28ge
Xh6vzg9SPau1tOnd4MZlm95wkQmDwfLt5DkNNwwU2F8+xVQVV+up99APOFD4yjjvtW1nIa8P7kAu
KJLT6Q8ZUsmBu5NiNzijpMm4fZhKal9Myxt6Qr9AJ2+Db9phX0lzGTVdc3uq7x14/CoyavZ85hjC
3BRA3raXezWsmRIEAOr2YPKXmrYHpC1IGxeRgYh1vjp1f2znE4LI+FQzi6ApPAW8cumspteYCsA9
+o1JLR+0BOHMFqS3jE0qaYtL0HxpRJno84b1XG6TnhrsxEaLfLJRh1ZsW8f7IY32wNCSSTRC5fpZ
ed2vCUyUEJ9vYvmJxDynJ8iqBX35cRTlHyS1BCv+KM+rnR8euj097WQi+cVEi/wAfTx6HGDkL25M
cVlO69dgBBvCUQ+d7lacL1XV1nSt5T1zsgWCzHZEOk/jCQR2uq1io0ss0NZ1tMTt4htpc8iTzxDm
uRyotJNzOa6sKenzgUUK7CjAcaQON2Rg89UsVPZ6Z/q+8bSjQfwchYiD1w0CI1WI3yjmaTUM9wIu
4zQPSJCx8H4b+Diy7DQMO0UhZYPBsbfqvCfUWJhz758noKS54HgwEPwCnmtO8Mjl7xaWo153SyGi
mm+C+u+t1DM1JXvfJZ2p1fg3asTI2qfSqeiDa7jOyim2Z1tET9R9A4VTrsPKq3ivj/WLUNhQ2R8c
fVxhmHeMsUh1mKy+irYlIXkRSI/8nzoD0bbtl9BA8bIM2VwgDthG0jzoCPjD/ZKBpvMltVr6k/fO
ta5qZJqNry6RKkXal5248UzrRJDhOKFNQDgilzrO4wreJgk3Zyw5PsOTAIGOub0borSA3TfU95xm
PzYL6tS3yRXlCRAgtu5yhReAZOTEUqo/m0YktYyON49OqlOHLQM1YhrzIcG2J1VcXhduAhJmWsZ0
vPF8eMEpzzk9RkfG6HTBy6M53hhnjO2PSN6co4ru7ya7KxXeI70JQpc//mwpt3ckFH7ZKG8ocbE6
6gs7gLenj0WuHkftmmigeIJBO+kKVYxfCr9TtfyGym7W/+sXIIoq/AqJlJ1AKYNaWLiE81cXhR96
qruWFaZErq1wx5iZldjnD0w9BM3j2Sr8qqvIf3TDCbNVybCAFPeCmS5KG0LkXyMc+8KcHGtivWGm
5gzta7KdNg0IPgoT5BDK18x62a8X2V3Z/1YU3pHx8x3cqnWrtoVPYTDay2+ygqoQ9IFPSWAZI/zN
mNY1B5iiv3u+d+I2MVtcetmCIYLvN6vMfqnQZ2AWcoHkK9lW+YvbmcKV/FPj+F4k6tZfSga3wq1c
LReMkIBTyDjMKXM3OL+wfcFbCP0hpUoXDTQHwDoyT+27Q/zG+9AQYwGr8ykX6uCAlXZtI2+Vyd26
O3v4WraMFTCanYix9I3K6S2/TWVMrZRmZLwpPRkWWn4ZvYFiySg5Cn9TC8GTAzMOJLaGv632JSRw
LYpEBhJwXDu69FJQ7uQPQZMN4soVVaK0TunFVdD2gPBpU8G7s7+aW3rLidVyEOthExHVjOXGGm8S
9XOaJ613RGIybCM/HHzHg4keo7c+LxY6E2EbwSY4WZBHRAFk/Y7okZkvfOTDyUtd1RV3bYxhC0DO
t/N1SG01Q/rXthTjeIjWhZoiRM3F00lFkUhV6TdK2Ik+XfKN+9ytUub1oA9/W7wazxDeyl9D+t2O
L4tPeoRYTrgtB6rPdG2/e7e4cwZxWrYgkbYT1BsTELpwfKYEIW5IDXD1FxEJzOyHN8labmrpYIPy
sMh9oOKKmHsCNFA05nYf8hJmWNh4E/a7j+IrExqf0GgWgzcfCEdUfBFGmVQC7Cfo9LYr6IosGrtB
uVbbbI0zuj6BwmpZbdd5MRd5aD6WfoUMJVH2HyDzTNjuBCh2udorGizAKR5V+4zsMRY6rUFthUqr
Peqy6ov/qxkRms3wxP3cK7ts1K/bhwP5L7HsniIQUUt71D9z43cfZiLKVTPzJt1VzGwKe8v1qpXy
W3LdhvQDMbJ55SyHN1qkL4MnCsT7JImcCI94UrLcbwWyXstyuXY4Qz5m0shvj6Xa2801LkQGTiGE
OvkDCM8gYoMFhfU/wOeDfiZNJYqKcFpZBzDie3zHb3mgRCMPYDBTYyAbiiShKoq4qQd51kP/oidY
AdiLUErZjRjMfTUmyKiMP9C3kzpcBLBQS7cm9g00SXPKQEfSTcJIFHZeclfrdZ6qo7NIR2n5XPfA
AYdeMgZybI0Twicqu2iWySfWz8cIAasPumtV40gz255GP3zbM2px1zPw56FanzYtrpulLblW1Doh
YEFD9W6dG3ZK8AspbSa93XtRCJm2UkGR82p+oeew/ler2aOuCyjGfFdxGmc2PATrEm/PZNkPjbHW
7jQnwfOaz2zaRsKiLsFa10HASJSe08SUHCEU8FHrN12yiLqz6KrYIhiKcmaACbI8Rrg+ifwefcPn
U6dguW70o8EVUVNnWrogkq/raj9+LMfdzXasZHw57dDATLX3zvYZ47YYWlFxTZmk2zm1GqcUwMgy
N7cESbX6iBUaA9LfqkjlOkFVSQbPXfCt0rmBs0chapg5tgOpWnszNY2xIJAUUpSoce48gpjozpLb
H3uJrHDXtlViDaOE2BcZx2yHsKDtRvAd+qeRegLTuB2DWwBpFF3l98C2t6wkQGi75ZtBuCsi8Htq
mOfsoBC8P5yEx0fazUVZojKxWU7GpTPEbQn39XfcAMfRNog59a3ZsstuMZGFxThj/omkhNQ+2ySO
mE3W9lLSgaeqCsJLNYktQiBokRDBeo34NkoPXYOfANnemZZShFX252gqGSuKDTC5AMjZfI7WSPSD
3oKh6aMR+7Hg3KVUQic3JgvXR0Su+h2U6LDAGk9GSzXnoZW92GINA1vJXCiOCFREHAGkVj9RzJLD
Zvh85qGiXjpOmSzBIT4++vuwdA/nIz6I13v9tgmWFTkgeL/Q+pGWg3HTDZMu17j8gYIR2yTr30jO
koC56O3DNk04IemoCUWZBAeyPSwD2RCNSQTgcqDNSZNTCc36tbPC8tnvGwWo3YDcx6NVE6c83U9b
8eqpjq4IJqYrAeZvxJEG4Z0rREV66Ymx+pCUHXgbImTJpjCgBkAQLrMu4/Dgfqg25MvA2GBzFMaM
nqRqoC0Oobg1xyuV/dt1W2UgZPtq2JvShDgDaKewIq/U8Z6KMUIgSLpXWcK1lUTV6DkeopLqBrNe
MPBb7YsMtNM1LsSTSmQzuJMwW3vXAYyO8bvCQd0sbL8F2tv3JYdGX7pDiqtibNXh1BiZNIKKZg1r
Np41TcCText0U1InsvLlz9E2QhhSnW0hTNBgoaUGTNsFu8W2OnHODQQ43CvmEUp4bVvtsoJyCsSy
TyGyvVQeID5xVUc3/oTjXVV2whqtxzwlKomVxDD4UhbalbHWgXCNqd7SbuEhecEiY7/iSBKwaEac
TU9abLAsipJGix9GyEmlUyW3/gnkILkf1ohmbPi0xl4u/htduBEdlkPbaS8qL6zu/iYRzsriKGCA
LzlM2xTwyrUKU33PtsDyLgnq9S0csDGKzWz137O0LZ3IyjhC2p97XgXbWO5R+hvD0Cw5Szk3ONU4
hDigU0b1sPyR1BbfKmOKcNv6H8YueXAPa4ewUJIX46iKWLjaGtnRq848UvEIFZOTLoeOvx/dq+3t
oDshIpdbA8MKXHT1uh78Cra8LExSPLVbHBhUPDIx+7kCxzTp1xC4rUCb6WNJWShLVh21x9i/2U+P
cj19HjYCpnDyC700jAPgDHEsYDQilOwZSc6tSbD/NuqRfH2rUmU9/XX7rcwjib9Cz3CRpJdJ/PM2
6YUw9q3SyIoYcmh33bKCvhLQUD5/li6XM3nCjpiZ/6BJhuW9xDAQ0xResg/QRRCyLnVNzFmzccm6
YeQ/QDy0UExRUZ2PhgH9XrDopKHHfmBA6nJhzjmKRqCJi16znfjtWnIsP1bi7LHKDVYC+IVePLkK
SMQWPSnVPkiwDHRc+1UiPzjLrXsf7i3KQdFGKp5di5wsLnSUfUnb6LeZpcP9WFYLRQZv/1XBAt5j
OOzqa5hgZuQHLwNiG1MEybovVtIsMJ0UGRUePzEg+oqLryzsg8IAdDzmBzep8DKMmPwVm8nRchCB
gxqaf71Vvp3Kv+Al83URmFndrPrE2VcidMDfEXwJPXjJ4k82vKDweGQTTaC8mF7s7i3TI0DyOp0Q
cIpc+8Zt4cSxdHVeFe6AQCoLJCfTj0k3U+UBf44cPX1TzTTuYVDWPj5N0UK1Op7tOPmUp7cZPg0s
g74fCpENOvq7hiPP+8ykrhPAnO3MbmjDsivaABA11tP6kBz8xzUWfUyU0G/h1dg1Blb7Jd4BGWJF
pBd+acECnXmPgxRWIVfRTXwiEkHANC+REjE5LDtVbDOS8SHHiF4qdr6hWjaUil5m/EZea//pW8Hb
ilFJxnuNRwFwqwuNbcmWAfVWuM4rS7mL9WYnwNM4jdo8ggwDauITP/zWyCg4IbNAK4X/qJAFdo18
zPNZCGmPgXh0c4oE8vO7JoInV16NErux8d8Z5uKITjxDlLrhfYB842iP5fmXenwn0Kpb/Y6dDZyI
US64wCEy5YqL2m1FXpmQj51Hhmonlvhvu2p7Jndc5s4yua5gajwdpbhYOLe7GitY9V93P0K0+Typ
8S6/N72idLe8zPKqWzTUrNA1oEJeZee9lVga+lLTGWJGhVw7IM4snQFxl1DEPrQUOdyo+PJqyUEQ
s7f8u0pZxpTkiPlqK+nogkQTcatVMgSSzt1S+KjNTc26VjkZXT3DORC5MOOqIGwS03dTh4xBjegO
nToKOt/DjqYKccKFnzXiCdHgiSYefvyDhQIGIPRqVKGybK9xi74vKRp+jrtMggkn/TIuwQpq7bxK
1zSmSc48SpJrvvn/PAaWce5iqj0+HERkQIopVQ2d84wQvjSyGabRYG1JdY5c2AY9ze1D8qoxv1eg
DtNjSp7isJpdMZV4ROSYhACF7iLtCUJCxUlMnv3DT3oF4nXoCPseAQIblkHwBZk+ZL7x2418OgBC
bPfuE7ssy/VcXItOCbcPwTwPfnwX746g06Hb+o2/yzEekafflbPhUp8I1Svc9CWUw8Lm116cudcp
+JaEUZDBCDv+eWNmw+EtGPiVP9syiq/n3ui/Rgx3IoEefWn9mWSPZNM+S5dP634PhkeoHhEjnde3
db0D7hDhiHWsyMfY+2aDEJm8s3j9GvoViHH0vMCucQtXm1mPmwFQgtOSRg4xjOihEEe7vPJVBbH7
X8qebnEtc5SLfHVktA/kuCgnafA+weVId9rmOLKml9MpFuJwEC8RAbDvaQo3LMo0+QwbjRKakCsD
ovgRhpmz9+8yWhTMsHf3Su05kuh1Ag/4zQ5GOFS2Sn5bEVRL60sU7MnU4rn+4guUjzmHK1gBc3R+
jDTQ6RW31c081u4a7aUELtmEJx+zIUULif9o886lN8levw0QL1Ki5aoWYKvP/wIdxUdzshw6QVu6
Fvv4tvwQetgTqRs0CsLVddSBwA8SY2o3DI3uihRKi1/JMmXlmZp2WIXO6i5aQmSIkfE24G2rhvv+
W6k9g2nJF+q/VjdBxg66zHyo/2zrTlNJ8It0G/qM/AZxMtT/ai3JbYvo/zpHUCF1kIZaHgasYbYO
O3kmjNV03SH0ywIuaKnUdscAqLVe7rFoDE/4K7Ah1jK4bOjp9J1qLdoeVvspE9c/PXlyZa3ml2kD
14dh70DrVBcSbiPZ5M6kIzU5LPflxIotDsMEKUpVQrqPewE9WYiFqJJyE3z+hKqoSxsZVeFiaKxu
qCtrlc6IsVbwmuYXz6xrl/Kr+4QpAah9xaYqt2AtwSSTu7XY3SaE87EDwZct2Y3946TNOyVpBU1+
+TbPyAGxjatbJrNRIIKycsvIZsk6JlPf7xa7NO3IRwzCiDX1lf1TIeLnpUHG0zzl9BhFQ2fbXCdp
Owh7EKkfy14nU/yv7Zn313qQ13vklJwrE9C6Hu7MkVBIwbeXgb9bSyWSP/zl85HVOgg0gnvSP8wu
dXe/b6MQNX34RxHP/cVY7LbpXtpm6q+tqPo1VlzkxzBUTm1M1OZCLbAEhkdPHUSwC7pYywLH5Qqq
7pIP161zWqacr3fjLaAclCeTf/fUdbhzRRgNZn3l7Jj3fW+7czH5+R8CiMMRVlntVAsEZXYxvMSS
IVKf64OwwBkaCb0wgFLZaDsjIWx08VvtxuG+Ia/oVkn0SdFLHVuW95WNkb2/pEc9MxliWtTigh8+
lopzLj196/yOwUGWk7zhZQ2EngsUf21SkDW5++HtqJS41UUIfCE8QksriFa92kkc+nEf8zmfY7ce
2pz5X4XSzA/WrmCVf9+2+5DLXg2EoVAIchilm7ez5qnJfpcaSrw6/IG8hKdQaZewCM0vqVglHr/3
0Vp6sBVjnaietrQ7cTDVyEGK9y3bjRzxn/EjhnSOq8jmnWvfdVH8P6jr2Nh8H9UJRVj768umsWT5
6aqzHRCfrr8dtV92XETtXvwrG11GkiP2r+6WNXAmSHuK2lo9vT81aowAbMFsnYqCGKg/7fkXl/Dh
kEuLgZ9fyF4RbstpdvmJaDz6GeRE+KLCsD63ocUdLKblKAD+GlC9GX/wIFetb7Szl45xY+tq4D/o
wxUHqhvu1Ruot9sX8bT7IBd8X73ZakqkzZfqAIhxpVvvgVvWqeka/XGkURVNhEE/IR6bWyXS7h8n
QfgCZvavkzpg1/qJLqvdhF2HPhsvYCNyItMjrRTDiozCYbt7VD+QQG4Kp0H9w4N7btE/4smijDeC
sYfyPpMjB2pbVnWNHPWxE38cSk/uwda7l7b/NZlmaF4W2gxK539P8iTYKxkmaCDChBeXzybNre47
auos8ADU81sRlEQiCIDINnjhcon62cVm7hU1pT4oyAeshUoQej7W8MmP5m/69Jn1U/xgzwPz6mmw
l3ie1ze+gsU8xeUw6QWmXAkyk88EEOcvYKE6OrzOaQ7l5Ci8p5SIGUvQWVTVvtyE/D+/5nTLf5yt
qpcrohM8RSw3vRL70nNZvHTr+n7Gcx7wutRYCLynzgHlGc3mf3IqORI7ilihEpmQMvN8hYEnRah8
oq5cbWpfYQMhtsHTvzFjTRIzo8Miaqxd0DUleZKq0GsgxbcWuYsDVw+Y2zv+PP1dXOVn0q6jVa1M
iBIgH6Mnce+0HbNY3Z73CH+ZwoCykOTz+Slf9CgAXsxY/Xuk4kewklx0/GLrjzZ3QysGVFST+Da3
fWgV85bJ52SsZk0y2/KZmePx7PTwU07Z9S7Gj4139QLM7rIgaxG9KVnRgwIWwRp2texhm1LKR6jK
2v+2AGxgJ/vPS8LU01HM07qBrDIFh0Njv5+9rt7/tYr1Q8AfulAkW17GPtFM7YElg5rNF7WSWIHo
RSRB4HGtmPYu9MbBj9MwMsozYA9uRO1qMMU7wLTyM7W8QcsjYTE5L7Z2ndY93pLvnh5otBWBvuqj
KATEvWrZ8Vjz8HPV6cVOznVS77ezDk60fbv3xIBraofUEa+fxcGZio9sqVkkzm4qE+ebnUnBGT6p
5LFC3iW0eEUs8prVZEBUtMQM20bANsY82qdoZj5oxeDfHMRVgWT94w==
`protect end_protected

