

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
cQDd3XIPPlgRDhqULvYHvwCty2ZrVwzfefmANvx1dZIylIMC/SlAcj88wfYJOEUSOPC1U3p3rRJH
cF/G+RPdfg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
hcwXqOGXIKp1yMXglvtwKNDD2csTguI/218BbAfP1Qe5YaY7t7J14bh3PN4/sY8v5SUfs5PPhYYF
AVoQ7+Y8KyIAkFOjVjl8Q3cizlaMAyaX6UCc4wmflvCCOjy7mkT0VJKPELyiFH5OE1gTiKu4NfqY
cLpas2QiSAVn/xZw83g=


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JJiSVarYWytdLFzHp3wkrD5+jxEb6zxCxwIxMuHES7X4vO/81ppoMZmSB67P59pBX5Chyu0EswKT
bCRha6XDZljqkcBWrrqj3cLRE57UCaEr1RVpDNBMw7hjNrwCb9eTELEwb3X0mZPKBqVrRNroBMN5
Mb9o7SPJ2GKhIDEDF5Q=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
x9rjekK3vn0E248BFQkRU8rm2REs1XV6NiMfscimCVnt3moe1QOgVJzTLPCcPYvThLcZJXwVyFUX
J1k2lVxuHKaC3FNNToKLX7girUcVANbS6jS2AjaAfdpYmQXF6epSjXy+KOWM7AfrGv2r7XNIcV6T
P4He3ZDDIABlWanBaDiVD6NYtB9SspFXaifjJ2faT9Et8gWmYJogYQ4BjXl960BUcxWS5faBudWm
MidcfsfVFpzH5bJ9L+thBkdIh/P3Rjr9ssCSzEagp+1l0DsZGX583KqMaKiaZiIsR+KyQ8Hrld0H
vh5k+kh3k9z7ewkJNwM0LCpa2Y0qGSJOxIauzg==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bMGW+/GNxe7XIGxZQsPwYg9NhBUySelE4d3DawPwcsMkcAefxMJ1JdlslSvSp+VjxIobQhkauqfs
plGQEEjRkhr+3m8iz7uiwT6s+TtBZQ509t+m12KAHsziCshi0m7JEPgqnpkYUxS5ZbKQCRgudms0
J1TIIpIIdBJiHjiJWPFKhl2FSk46olekE0MQ/LvS36IE6UC8sP+H2MLZpAxpzqHuZ9TNFvVcyr9C
pc7viw1i7pElJF0USsLWRjDFrkLdXdznJwKPhjmDvq2WWhH0UZss4B7FZEDrUrjB/HO8EjVy2Hj1
fpw3eQ84VC/StEBHWhh2/ovbE1xsoAsXeBE8Tw==


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pp8HZNaXt/evJqKzoiOa8A1cmkUh/1mQf/2Vkpam3N+hCoX7wAAqGU/zZVMPYP16RpMjeC5zeSin
YvUeVcdgv5x+e+joKUcjexTi2LwQorDqPIl0bCwYx4LccUexnWG6I9/pSM85Q6QNP03F3dTfZ+nY
q8I48HLVTNxhG5xD9+JTBp8D7rjXe9TJGi+hVikOsYhuY2PrwtvuAWhuicAfJnsIE23LJrp0i1cL
6oyVsfKsx+68L6qOWniySUGZ5yDe5zDF3WoQ1oHIZl8/tfnTJcGPsIRyeo3fpk/6/w5zWnz1pHuZ
HvGPaU9zIF3KNoE/3qKTDNhAcVbvP4+ohJfKxw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 69472)
`protect data_block
ufGjJ2eQAYu3yVAh9icN1qDiHHgwrnBgbUDddBKkBCyjFMjB+HWnzmAsnYyIpuveE+k9wCbsKycn
YMYMJaXx4smi9tU1eYUo5h6zak5ZC8bxESTIcqEX4IDxE5jrCOlbLSftmxzWmCmwQbVc2rGFyC8M
TYuznp/fbvYN+IEe9bq/jEiEPnGIRcad3jXBEwBfY1gMdW3zUi3PSbRq1Mbu6uIt3k9uDlzSQFHg
37nggNZYolztf4QCIC/2hXyzd/fJxxhefA8F3i8Dzu8qS2x4uX5qdCITYmCd9ehBcx/CcspoyyL5
5NyPqriLsgBidlp4w3/d5mXyKiZNnhyxf/P9PwV3vh4jIndkqTC9cbBPTPccuffrJM1DJ9RJi8Cb
EKKNBit3Mb0cSOQqCagYd+I8Mpd2q/s5WUUztkKNcsfIFdiiZEKfsEBrTQ88iZephyQq0kbnYep3
N5bfUdo8TvRIXEVw1we6PNlahUB0n4ZgzY8VgbS7MgWOmOtT2Hx/6YTCGk252ktpEJpilvIl8VBH
LZnfo3UUhEyGtfHWxxWW8EH0rplYsw9HbcejjT7UjXNJETJqG9WG6/zz349/o0r5jeCOExjPpVMO
NwcIbjqHK0yYyVJc6WZfqKkFwCf83dmMje+ptomi5JqMkZ778n0FM6jP+OUh+dBuSvH+UVSLYEVp
Xrcf72fugNpqO6a99AdyVXDLrxJd0dVb4XV7PPc6LOpf1B0doi35QdrVvRNoG1QvkDD4JBeo7MBT
6WzEBr02rCKzUiM8U9+XwbxmQB7HZV+ULqSyEuV9Dhl2b7clg7WAH+o8kjORq/1mCxZpvf46W2UM
3S40DVBBQvnDTEn+Kwmk5ksv7KMR4mnHEmap0C+fXnzcQrgi9ZI6nY22dYOQ960c5Z2Na3FnOg+9
xP/DUZteWtGVQw9iIoEHts+RvUyh6j4lagg5g4T91isPlB6OkFi0jDden4FKc4di3y4FTLqLcHG5
LC5hGPdCNyZGENV7zIIGIv8PlqK5sMJfkxuWzVjp+mai7vzLF6n648m0KOJOKlJFCjJZi0IpGBYp
Kgy0WvD7SAsvevQEup14KqRxg5NQZx13Wmm5MWd8JI5o9KOEl6C8eHKLtglwrfsVcI8/jaB1C6NG
CIQd9O6ZHfAOzUkkLSiZTcU1KNJZgY2/wjOq8pCwHGJzwp95Q42UoEqXbOiuZt/b6tFhtAMBGnU5
f+pghvTa8sEIIZNPgDdkogyoOtu7cg0yznZ8X45Uep5JcdyRsj1B2mfqv0BUPHTSUTn8xF0YJWVX
xNFnEh6lwDTndJ6cT8bSmgsTY7fhr3G2UJnS+1FcQTclfdxCphMoElMXhfu9MdjWipbtHshvwf5L
Jx6OqOeckyM+L6Eb1AKrAzrQMFXZmiLFCdMIv56z5uW/AEq82eCLXe3smnFqNtgYbdpyD3KQeGBz
7P70F4hNU8RP7oiWDX1XyM2yv3pJbvU+pXFf+Be9S+vn12BdpZLZdgUi45hoyIW+Syn6ynfsppex
uCgKEUzQruADiXafYIGPLCg0OD5M5YHvplG0+21RmVDpczlMxrvppMe0eY3sZ3hFyuNWiZqMxOI9
mTFjEfCE7RGTUVRq+Z7oQDLgfdpHxjJFME1MuL1ASoyUZUZOIqtUwxmrnVv9+vDxRFu9XVlz++8u
btNVXswDPIWEwFwq9F0c+0Kvv6JcILVPZpxy/fcFgK5/8LUTVeKZ5kGGBHeZuW04Za9jxsPOJs6V
sfg9L0n/8NxvkbSCmnWjg1GBsbzJu56CxSiC9rfBf4AXdYJQ6ywXOmVRrbE3kQgEjmlEeI4oIGJO
2onXOAWEM1Tih/m/VD42w5AjKk4zJ/GWn4Gj3Q/ApNRVBUb7lYF0mDleI7HFLAIupsLZbh1oHG26
ppjYclpfujdF1x+KsJhkBRnbF7Ma6SKrIniI/EiR85monrZRHPUBRAY+Xbf+iocmtEwE0Db2CvOe
Z9x4/Y3J/hI0U0Z8ZwR/bqixPSJhZ3WqYovjFMkroRrtpXY5EGiFEY6wNDwO0pbEdbz6oKImtIWk
mk7UqYu/Ka6dTv81fmAa/nKGSOZ5vLszVyfk3fOvr/iquThmM7nxYUEcaSDB9E61iePro5sppzRr
FTfe8aUcZt6GL7U8Vlfu1jALEdw8hVtkRIVB3K0verWNaAKMC5WRt0ZXHxQVpvee+Pf4C+90F84P
LUxajtVuTvHCpuUJX8fk1zkAzzBU8Cz/s3xEe6nIZSen9/c/xIJwWGzuoBp9vg2sZOUVy/bIdmPG
2BR86XFmJsmjYu4hrjYwOVGwIquzN0/nCn8G5J+6qTdX7V2YInlvY9q/0BGGOMQASZ/Uo9p2FVWq
iDEMc+Dq/mdK2k8UXPqOWtzPiM8nf0WwKxsBOSo5G8FZOCQ/Rex+DiWSMsGFM48R902pawhVd1So
0WfJepAlHJLrdGPpqVOFQIZaH95C5pMpUrGEjg9Zs5fgafp2OGMTiWZkg47MOzzb7wiNckAAKkmO
x5sAo//0XU1tL7ZMZHSKdsNvi4xx2YiqW6mpVOtOS7QxMIs47TXrY2kne1u9UGvcvEVVbeu0Ultw
D6mPRBIsOGTwkl2s8Vnlfi9y7dOm88HAIyTJoXbJIsYdWXu2s+eBMPQ1thzZlZN6LwXdLxiW4uk2
OOgsU9pnQD4Fid63us+fi1H8HMwaCm7QEcz0viyasorn+JcCM+WZOL43Eeg05Msz/uDZ3raZ/Om3
SQdBhwqdli5XC3QTSqfJIdd9mCg1exRIDa/cujEmIB/oABTYGYS3CHXscj+SA7jishtfxY/nTiQQ
vORRTz60jqajtjuRBXloL/JPeeP+C77b6Rb3JtsxhIyt4svHXIz61upDLjQ5zWc5G1Z7hQ2dARhD
F8teGP65LdXKU+iTvLT3W0vgU42HLxDQlkUCGgjTQJIEGjI0pFV3OIfWbwoNYiWhd2xyIKCJor+v
8SnCBXMVn8mwpp7ICvP57Ib64V6sQYNWAkI077t5kzORO+1SfEjoh+8PhhbXIWCNZaxPuphEmzIA
yYfuAFpT41+VmYQW5bexDg/BzoDRdHlu5mnWsrHr4M3fNX5zyR6rPWG2SO8SwTjJcvpwvZoR0r3C
BAwNQ98byeawV+zgGh16X2JQNfRBuaKI/qg1/Uwa+okNUGo2iekI5s6Eo5fxBMeArSDvImTmziJ5
8PUuoNXkC7SA32N0IeKbhCq2EIA2mQIlWmLCLfhyuCPa0KUPFcGEc9fhQDvRqfAmjTgQZKWTObmd
9GSwz/K8nuZdxMG/BcDhcVLgOcuMgXXnVw3NRtDQU4mKNHK79XmLIqn4gYs2Vcdjzt9+5Yxgmuwr
Y2g8CkoBwc01/EBWv6jHIwvMjAbHY68b+E+pNxPq+oWH1OcOvBA307WHJ+42FhA9YsD917koV/fs
ovTcnNp5wTotM1IFE88/Ytock7tfW/AYi3Po/jEThBkGSYBglGwrM7UVYmAqlkr+KX5N+J1GI7h4
/RWY2StWlhTUAdgsWmX0WxVXofCbF+KTBWB/YPK/8GMgsgWC3UVqq0VYXReF0vNIKBX8xjlGXW2a
1t8KgCiLPsNQMFA+IQliRASYtQnQJpSwKtcBqXpHBkSwXDo8a+YvjavBEFpR8S2e2kzReqw+0ASL
JqBFVZMfz04shPtPfL9GOOJUNd1o0srlqU4xsbD59Of0lpITJmTHjA0QujpR9ug8dZyhHjyzgC9R
FprQxEJBF5x57QFb6RmMRx75k67nZNeOh497ZeJplL0rU3rkR0C/D9uFUOdUMAfmaX/ycaVfWk7+
0IiQgokMDxsNj300G7wiwGKkMK5bIm9w1PuDMxnfYs+PK9jpCKmLp/TfljBlgVjguO3QcNz8EOqB
H0ryFPiXkJ8fHCIJw0PXUkYLKrDhLQG33CGtTiwLXGWenqEJ8dRVbTEhmguqMHEjRM0Zi1kt+dLP
ZEhWQgJ6aOoAZcVf2sd7anY4vS8HuCUiXuSZ9GhGYFf+wlQtiKjMq4P8DkglScSvhz0MAUKEbwzn
dhOAW2DHhTt8BUie7TStr6JQqSt4aAgQ49kYo3xbXG/pLuk8nn3LpTvFHci2WplgyHdtJFHYZ8u+
9GlpUO+RrqNv/gORZvGqNY/TSK76ikxT3/Z+XfHObDdKe7iLMn1rBX3lpjH8PGUjDnJBMxW+sH6x
odllG3UAsDs2+ELjAp6vstTJhqg2M89cE/GWNlk1o+89JMQhka0kSW63jRJoZZk+W2twcae1TAzT
FHuHQW/pfyobm9Mccs9Q+O4q4rsSCRXH10WNe1337XKWttzfIiw6Eh9vMUxC+B0g5sbbsKPQy6bY
bwBKiKpq/8AsSpnwQJncRtOgL5ovs9nVAjapxefshqB1C0keC91eEhfJUjjbZMCgYIy61scYulIo
e48XsBeYiGh28047h/VA2GRxTXrOT+alhrMwpkc8JBc+gKmdJ3TVQKuvgUFexW14aiW0IcD5TJbW
9QJqnmG44NDSYyV7a3fScff/VKKVVIWT7MNOFr5h5gRNcF7ySMK/Tl+AQO67ddt/W5mypFWM67Na
oQS4W+SOQC7E0ybe+FepFjSeu5cEm+6TPm+4+DUvHrA9ZqupLmt2KXMXJ7oRzMdbklcQgLLDj37r
NidKTEdGLSB2IrR7kqr8HK+JmFlqOKse84HJ56kTIAIbEj8+aXsQ9MmLRgt2Nb/DnSKwxWdbhC6M
BqQ+GCRAOC/6JcJypGwBBiksXvLGXttCaNnC4JpzR3pdn8M8vuqQP6aoiT0XWcKWQyZ1T0pLRtvk
qd02qZEdwjVb71sbdZcvmvTeWydWMmojU5Yp8L/aUc2CWfF/IoGQWbUp2gfAHwP+z6mpCK8Z5roE
ZiY9Z9wRqZEMkT1GHDBgGDxjauIP0GjoVQBmxG3USlic9oIueSZt6+SadMF8MZdH+wt79+tVOE7F
TJ0xwVTE3i798xzpWXKA3BEfLDUeN7BUnlvFvpuE7Ig3JwHYxfIh1gjyv96KpvVWUGMt/Ogd91Uu
EDSmK1Gaq7YKUI4dyDFAs9SFb8KiWDPxwK9BJX0aBiXnlqeEpM3Ns4138q7mBrJYZqX8nvQbE5q+
XVGNetZT0rcNN2BPixU3qsKl6IgFYGsV2BawhmRyir6DTfYHtyj2wAxHD0kPLIL8ot29pmUZWrlO
xt3bnmSqLFsmJX9QDo9fOnSQavUdAJbq4GKOJGwl0Z7gPaIFFTT9ESu3KYUkB6d9YsRRUebPucr/
OFh10eab3ba1mLfSmiTYBQ5yggCRA3Sg4R0yZ0tRQO6IbTiZJQkT7LGo2nAVYcDB7DW85h1FUmEm
lMSdUxWG6RTtAMYmck2Zw2gdpax57iaHaaexdfzHzd9jK75aKK4HpeyBYTLt6MCdobp3TXEoRYQA
QTVLVR2ANHzKExJRNjrXBJrp0wySsDcoPnhWM7DjQ9L+YT04XGfM8z/8B3lD2cmF6BWQNRZZyeYz
mUBmL4LLr9LiwhfanOW07bkLWu+tSE9OcqSgTONFUqhjsNWs+tGYjJVlVgOWfxn1OG7GPkA+GRj5
wukFeUly+9mxvo0CZozaluMtCWQPXfqhqO0g1CwGmhqGidL+TOxU3A4+e6UD+q6C6j+kt+vM9AnL
rs21plOlu2q1APUtExhQG6P9OUzf/wdU0aVeLhfduSGonacwxYgoEgsKus/v/N+wVvWJJpRsHP7g
7PXVT2h/aU6Wwb0ywagLgsCRRBQZwgaAxMxpxJyOt1ZcEgxJlPR0wbDWSrtgECrs/x9FKpE14KSp
1RM80avRf3TLH2o15Bnnmv4zJkYl3Cm0iTDT8WZ9X+J4u1AOD8KjvVxTZrJOZtlPUjfNJztW+MTj
5My621fu1XClhj3DpVKslk9oA0Y+KcjhldkqzSus/DHZFtAfh7PZjrmnDgUT94hr5A6UqpYIJTIF
tJaPQE40zYxgVoPLfhJSlaKcRJDOQ1rySYFFgup/Q66GdKgRKv7aO9cOx3/7aPyHnDnPnptBWxi4
feqHmoWwKjBPWscoAB01XdwNYcSxJyny1p9DDXSpUY914oD5HfNzzsHcRqNu+4KM6EaOewVll+9o
V4Yv+jpFKqC35FDNdw76cyoj8iRxQy7A7WwhzVWfpcRGfI2JlUENzA9/gCqHImLfh2m9x0Gni5ph
M3m/rCWFPz3XYYJ2pcN+50OouqMBIV5HqO3U52lUiQ/gNBoVzWjyQwqtx0K4kbjhra0pOpD/U9Po
qzTU7L1zo63S7Khc7j20At2QEvc2sIQ760/vnGh2EQPN128DTk2kOngaTrqjFbBYLgc9rIWsYfU4
cvfNSXG15ml+noMQAvNhNKYO0/58SszzKo5tBQt0WD8tQ5dl5fOZpl9iNQlenXHSG294q3OAmKWb
iB2Mfex6wcGYscCqE8fq3Lm1hwGnfFhPlMQsrUuLmNgTPIiTZUw9OJcUI/0E5xw+gQJ37CFHZtEp
OhHDQdySF7kDkxJMaIBJM+yjMdfecfZGtqqLOaWo2QXA7P89JXU65kNJgFEi21pe3TsnPVwhLUAR
hlLG8ICxTo89KJfyB8dUJDKUvLBSQ99ro81xvhNQlTAntNc98st+EklR4d6LK4N2ndOEQCYoichq
FgUB60UpBXzlUXkBxsdvlvVzlq0T6gokhvPW7o6Yb8FpKij1J4srokJmLn4TYxR99py/1yRW6OHo
+EumkVNbOKP4d8rTp115LHfD865cBib2cXBPRpGd24KljbvNDuPbpoV0zEuF35mfY/KiapA8NSIA
7408kD273KuHJa4rQBl+9iz9kGYb3iVjYOi5Sq0tAaOqjTfoG//IhabV7rXp384wEW1f+MRQ2c7s
a7sduroZlm4Gve90rl05nnujEzcAlULCw4K6j3KxgkEVHNBF6cHh14CQLt8knd1L2fDllytnc9Eo
WJIVrOnJcRjqKKxx4Xc0L9K1DKjzAvcnzGmXrTTX9miI4iNpXY3TQeQQ/v5VXdQmRHHqTeUORlgB
EaKoGO0UCFL0hOz7cTX1E5SgyOyoxHQO/zMoYiyxrL3jCJONYflf2UQdyTsW/M1XpjOSwDAHgiyD
o4jbgsZrZx9+U3gvUxA6PZGTA0JNnSQ4ldFlNv+ARuxIYPBYcRFQNqriLokJGTsObTXv49EaiHuF
1WNn9SN837l7KIs/uTFDjZcXOCabuXRnyBDkFWCefAjXAxCcuiG0PbTCqPl0WKJMYgjPpAEec7tK
TUzZ3EZaK4mQ7diSfuU/hxBMslScdE7bVt9c0iLAMihsf+O3U8sO6duTdPt8KZyA8enoKxjkT5iv
cRVMZvMTHaR4OJkUGBvEBKZceXZECKyqQERbqnGmOD4/aBZRAFY1pwjoUeouP+o+S2TOjjuPD/Q0
x2pGUHSfTVRLE2RiCw/h79ornHzgQpSjvGpBEHtylGVBxJqnuMo/VeFUbD4W+AcHf6Zy9irDcxQS
eCIeEpGxljf+DLwJ5ZBGoqc8GL+Afge/dHGJT5AVMRJtLcWNrayL0sIpFf6DUvZkasoEGcYNSFYu
HivuTsELQduxAbzSpgchfLpYqxNtPMboTeh9UTx5Q9vnPUKGyhaTpC3fT4b0QJNjXiceoHFhRqgp
u1l6ndIvnuk7A0ITMywhBIwnsBRxW6lW5v/k3w/RvkKnzxETmQguHF9RXOdHztAznJBBeBn4zTFW
pgYcftLNDE+IRhmmExYAxrb/H07tWAsIsNCiOiK3jwYCyWubt+2qFw0RPoVSNJIhEaS8nDDDysH6
iGigwYMpVE+hdTuvKCMC3wXkCL4wRKbgpYs0FME5MLZGGflE7MX/EhNo0Ra3dhSYRMCm1HyVFU66
5YTfrmSoFBV65c6JsVnhZW4xAY22ti2wPNAw2mr0Gfh08RK21SfzMRhAbERB5Qgotaax/DmDa5TC
eGS5z2FLnr9+FWwrn13JYf0nVShy3FMOA833CmzPlckngswR/itxVTJJLsMo+6KuA8RdGx+lAFrK
AQjZP/zccL7YMrC6ZMtU6Ph5rXCTstN6t+5JsbotoWM859wSUP2cJHxjHjSffV+8pzDhGF8xs8Ro
iYtMyAFwR/xRzXfXrd7Gs4KMgsB0VP7pkSmiz9ta3zJPbLzyVFjsl0iicSqpkGzJNR2mYWJdAoNq
VnyN82zBeAW4hM+GstAT4Jpu8rL8r8QAOLR/UUveffldOMWBeVojP7+Lh2No/+9gIi9y49+TQWZM
Rvq8KcNhRsidGyIKiFcUSOFxrkfOhLgEvkEBpkPf4I2CVeuqNSz0oVLyxCI6bmhB1KOUA8eG/zPG
wl8hLHvB1jSTf85mpf9QSBkH6RPKyi7y5lVtUgsc01RETnZysoYePBJICMrOB3gDPc/Hn99OA/uf
mJRBLRSI0cbSXsQtzuEPQL8UCdx0ky+glFkDBzu9xDM+Ue/agQqzpmtGhT5v2eIZTArMGE2QGQcH
wRbsvm0ShWh0SrAiPIBzMabWTOfSq7o4gfonylVZ3QzKaSQwMuKt/xNExaXXyuemDbYxGqoCKk2T
dSgxH5N7Pp8QAGk4Ijb5PS7yo6l9AKhGtqX1QJHT4JoqhewOf2ZL8lwoaQqM9S9c/D4k/50Uz96h
n2148gjSsl66+NTFzIhxiSEm5MCdhYVI8hpw+7Zbf42I2iiO8HxSZn5RHX722obRlYyzMeEmvJa6
TSLBgrSLSfKi4KDkEfaHfvPOYhVTunOxF3RwEJPCUrGSbauzCCfeyTaNLNdsB1VELlJMKbNJEbw0
i9rK/M60281NlKuW/tsBFD/8Xq8xs7J3kmdlOIjUe5pcApZwi6BfJeOCDtdQ31PnRbFXCbR18X1L
YFzq5uMgXh7jWGu1eExbtghGnvcLOV9glEBtGWAaFA/M+GfgAQrzVRzoHGMiNPIQzJpc2YDbH/UD
nKp8piA0y+LPW8W16R1YgLKMUCOS6gKbk9qR4HWjKGbzpYqRqUyGzmPJ998N301PjSZv9JMmCqK4
sSnAqGTEo1n61+bAiDU2WgCCoiRKVE0lwIbJ/LSWjAv/5oOB7bi69479Wh7sE7HeCtz5bKI56bNd
NnD6tdyMvymo8oVymLBCO26hfvdzqhX/GZzNWb8zy7hzRJmBAIqcmkeKa08C7Ky4Nc8ontBLcsu6
T2Lb6vskPR5kerYZRhogoztQG9kuUuXJopKZGYiODWmqizU1RiwYWiThtnEWUBh0nTI5Cz80MaHW
S7N3k6zFInIHdfoWTqnp0W1qv72rGTRjmS9I5dRLj2D1YeOL9icz3ASheByT5iQArv72iFHsQoIa
MNd3CXtKCIvjZHIL7aDzWjp5cdfUDZ9UAfj8yA+N5ZwZx8HB7oYMG3ZNPaFGzz3lqeeEjOfzB2/1
+IkpP3g4X8yCi9i42FgNUMrYHMvgwyj6ue4p7jL5yk1bNB1lBD4atRJq1hCg6t+8OL9uQDY3MVAO
2/THPHMGS04CHXQYsneo8V5WDK+O6fisODgfGXr7C1qYZ9BuO8vPTVnFEjmIMfRlXddGwktpbnxN
9D0BXtFMLRZM4/KdzhDAp0Pnh9RSoJZZfchVV8EO260eCYL8+XomLNE2nsfGQ6iTLwP2BIZkikhz
Z5dDu6akrEb2OCtBGINbjclzJ99opbg9GrjK76pLlEjx3P7tL7S3JIAPm+0UHOSKODhemgQPpQIz
RGVDNDkPDc1HG2vZGdg1FOqjAJb3w0SNYPm7p2iOr/R4WCLlIryVjGwoc6Ei+kdw55sUKJ9vhpAJ
Ld1+XfDGnQpAzLgaM1i0VAwI2zY4vQUIghhfOzw18attGRGbv8bAwWGzNsYYGEWdr/45jTGq8IsL
nGmBsjVyUbzt0cuoAzjw8Ro6bUG0ndQ4SYdemzUvccFu467uLo10vZwv+QoaEATVUHxZPAdJJkaA
CezlZob/SmxTRkI+Wrsk5s1U4glRdX1XP+jnKIIU3eKU/0VRavvsBXAFlNNc+MWAClNLeNHVoz1C
Y4KD2+WHk2ibGsM1YGC8sKBCUlHVVWMTxvWrKtQzZJuJdzmE4jEsX3Ymvmjcd7kO6bN+HCKFbnrz
KhZSrfBYBPjRALEP9hUxoMHeTDu+UNMZz5V7LgeCnBE5O7zflPpfrxHTfGZyJwz06O0ZgbTgl2ya
y+rr2MCip/fj8x9doH7XtkCnAAu7KUltcgIX6j5Trowgu6coOGVYW8Ul0bvO269gM7L0kQXVxd+G
BrF6chuQDKzMtRQ3rMamsZt7lvCVmwmAMlvc7gNEc1K5tNPU+qQkL3nhpkTVi5o0WJO4JT+rzq0L
kh2Q9DS4ublVpKlH+fwrx7iN46abgLUNWHhRn41p+OtlYzTUtbRSfyV1QNhJYbuPWoTPWI884FVA
cRzSKR6zmsbUc0isHTeQs7x5y13i2hkJl0R2CQQbAXrzNUyQo9yi+7ONS9nSAq8ASQn5asZ/k7WW
WaMMwvsNuWuTqc/IpvZbbQoXIR/waUI1NPlTiWkAxqmci+cKTdNj1sOUyZm0VJnr4T9B4802aKZY
H8KQMycdp4t2IfCy0TYlJHmASzyDrY03MK45zw5k39TJHs6kcf6ou51qsetvEKTQ1ly9pIffM5cp
rI1mYuXVn5bCE00f8EqAl7NqdLUbiRbY08j4KNMSSI7s736wQS2ATSjZcKyzoYgtd+ekF27utywG
EQlQ/KUHLlrEu0SC8rJuOUsw+HTP8cbqLqmYBj9wd4nOxu5BrjuZ/QklltHzwvElyTHWhjiGRNhK
OHIe6EELsex4iKXirXT0Hv7nZownPJBhLJ7/G41E2rup5/nZSGjsdilpEGUlIKVMZAjwFnMA2RVU
v1FcmgpmMMoRiVI+zEpgs3Seg8c3mWF9K/pflDiIuValh9mLmls2U0BXplyPav6TeFsNmdYPOmIN
ndCU9MxXD6lS0Zpw02/NL5aaYROKf+0UaRrg7LxTTSfcbcuz0aKyzzEUIa/Wt2T2r5ui0ckl2fS7
tZOFzdjehBRetBjXGfGAR4LWJTJpymkLSG3cXgSS4QMhJ7evxO+sDJs0IGNnHzcbGMJAmmnp06Y+
n21+/1ev7KgMTG3NOiq1el5Xfj348cyTcheBd1+07nuBBXLl1Luenmo30LV/be5SqeKb6hIoFXYC
iyOy7oKzCVHvHy4+dPL9vrui7Q7RH7flxj3Fu7oUy3PpXijLx1xMoOQhCl/xV7a23akmNSKVx8Fy
BI1dDzcks/VlkuAzAJiPqzzvJbXLcVVwGw8I59tHrJpBsMNunv1MtNFrkYMX86QlzOMdKOP5S9hS
/qfOyMlhNb+X17gZmw3umetg4U/0IsGlgqcMFyhm5ZNCZ7rL/gMrqixmYiTNfDWKYxhqoBAMETct
tGth+UZhYmPQ2VE/m/OiTyOb+0K3j7s/sf40eVsHwIpkkDa4Y/cuYpjx5Vnp5Kr4bXHJU+AApVH+
aU5msnC3DkCLGZtL1MjBV/v2LfV1RPOpCjUa6CA0DyHaFbE+LW/i6uv/BGifG+O3xMRqgxX0zfQL
XDmVdhAH8u6cwrnIlhQYsEefV2F1RvZQCN3GryDJ5LyYvrBsw6XoSW8MR3f3y39Ku/xp8KjKaGIt
OBH0lv9QqoOhva2rgjimhhiCxY/Kpc4Kf5MA5fIluRu8VfCwBEa/rQmsJdn2tgaQdZN8oOAbPV68
+eIqNmdzY8VS2Zxf6B9obYxm2xwtjumIZqyIoxXhCBEJtLUm2y4WmcTE2SErBd9elkuP9lCAMcQi
zEaR+fNchvPem60/Q67o491mPJSIkLx7oocR7sxR1jHUZhIXiKmcbOGtP1A4L9f2YvO5bApMIyY1
qefYQJHegiey2Xx/xTYkiw7Ba45xwozWyt+Dazse8EFY0ekBEK/EQuLL8xGonIBEcQlBnKUQV5aH
Nt61bc0ZwL897DNw16KFD6YpIAROCQFjPcl0idFvJzS5nePKd0H4YD101KksFG9QjlsYUgx60faq
DRZrnRXLmXEL4gX2PB121YDalhY3cHuVnEqCBzZrgJDC9UJE/628BUH4dZClFRDhBymLxsyWbb2k
ze+5oXMBaxIrHjZs7AfCcAbkUcm+IlK1kDUlrwKyCmDCGexiPy3X8RhZvMMkjDx5qxDuTPnsO8lG
zfqZMHltR4wEE8aOiPpxN1PDRC3+Iu+iUFyiy/L2NMyn4dph9YJEN7GuYRuqNLQk7qpfrVjRWkb5
jCAkBvMSmds0LWZdQN4t+QkTZctQz5e0soBEmu1sMTZ6MPhiGDLRIo+RtLYF+4tNR6F7s85AsrIw
QU1Fs2Ard1JEN73h1+hklxol81n9ok/ANAuKh+ZX56i8UYBXEGg4Kyy+XqluyJWc8qSCo1z3vZvF
vYHy6L86QdRd466aY/P3ogmV98N8ah3KCXByZhT8eQKIzr7rLghGhwGbVJZfAQ6DcdXbHDlBTI5D
q4J0dsx16hegLnBLdBqTZYoEpH28yC1yz7OxmEsDFV4UDhctCQ5RYKzR5y7gxQYt/vV8OiVFkkI+
cva00Zba7jTURbjX7O3msIYOISD6dY+5OotUMUU2UVn5pUPLEuLHrTMUZUQP1GjnhSrS+PS9sRcT
PqSWwP6Q1MNpyC9g5DBBonCrZ0z+V+mchC/f10VzOSzeRUhGJuX5tLsTjFGm2irtIM4navdvtrmg
s5CM/oDTKy0T/8aoIeBDyHzpz6QeVZp32AwuoHO6LERE1NPZ7YsMSZi22GV8eak82ST7A+hwsxXl
ifKRe382+qE5I8Szjcx+g7oKq9twU7QlJFgJBjS2VMM2nIrHgOil4B7m27X2/cuspS5Pn2cirref
3wYHbjgDE/XY78S9SU06suM7qJnkId0VrbxH3GB0tFaHJx2qRbYx9/dd2DRe4V0GROLUucMpLO1o
kchPxv5jA1PCyFutv5wyqcLBe/BjqF33ye67wBmzQtaA+e5SH1M9vHgp0REbpUS2ZK7lwea/rWLA
j9PJpyMK0IkO7C4yTHggOAx4iq+T+A4MzIPhLmXAvmFTvlqWySwlwVIm2BMc12dqoacFfpplZM+I
686KP0Q9mYgAenKAIfezlhfgMBc4TBrsLjA7weGFduFkvNe2UeiAbxdc29jQOnuQ9mVGNie6yr14
xLNZ6EGR+1jfQFsOfBEc8HSo3uD35BUgmcmhFsBqDinF4N8/t4sKl4MGVCX8glRR6h/8Tf06ov4Y
psgqziDV74Y2W6voqjPv8PBqWWK2OGPNGeA400/CUzH7Ft7/HVrRDB54+d+UfhbTVtOEcfD1mRh6
c5gSZ3lCWYoWhRhF52Q3H48TuvPQWOhyzYGCSwFHe5GajBMo2jbPu3FDy1d9sJaQCtuh4HMigWa3
wNd6ogwTpTGRyjeVB5yKOYTFirG6kt1eda1H2cQr0o4xK0COLPL5eC3lKI/l8+fmIBGQrNtO3GuT
tnfVGDKGtCe57mYK4bm5uSt3o2zO0J6BGxjj53B2ryMY9JMeI0a70W5LKvZwQpAaCD54IL9R+ThJ
Gb1Xmk1U7Ny5fmQ5WUSQBTBXVAWJ3hABGr9oJU9lUXA+fdz//JHZnNvAC7jCiY3/qfg6p9OvVX8G
3a99u8ROR2tEuZ3N5XDj5wHKV7QiAqcIxdTSXEkFvJlXEoh8VgYhIN2/yP042Ofwzy+jSnmzoEFN
EAvV/3RN3iRiGiiHkwgcH4Ac/n3z+UpcX2SWOukqCsfK35cyAlnzu9D/kRrx37dxvbkUTH4H0hkT
LwDG6IuX0rkn/Uzr4piUo14ilAu0/n/r++RdY/3nSCDEfr5nna4lWu881k+cmRUliGx4+YqFeapQ
nHp/o6fcnCrUuJz4umVZ4DlodSCSHe9pSDP8eGwNwwNT2amQ2rx2KTx5ZFGTQ6EYCc8uRLGo0TLz
ei90GnpSzHTgUk/D000NNZdUfsu8osWJfhgjWlpNjRf9pqCkwvTyg1pFC9o/j5C2J0PB3GFt+bKt
i751bYUeBYFOh31yevPwkyvYxi6VqvtKszvksEE4SV9PZOacVjKM+rAB+nrGI0Lw4nB4BKwUMspg
EAnDWbV+MnmdmEvlf6GE6y76HGmYb1+0xkp5q0gFNBCb1/txrLl0Z3TSh7DBi3LX2a8iGxXb7Iol
gtdnCzShpQdgXTEkWXPDmgG/1XrzdrEiPQE94Mw8WA2tHz7+ws7TuL+oAtPtIDFhEJCpyEOsQc8U
Qapjuz/M2oZq+VgvvUIzkP+4urftZPhFMeJrogdeYejb+suhdqpqUCF7FlEeIdMh3ijUDphHIq49
dV/p7vkgOu0Gh1SKiRQzBIjkpsb84wceq48qsQicw0fgFlDaD1p1Bad/RwVgf+ca7rIRsROH9RDz
3Fc4f7GAtM6LCU4GNSXDYb9IdTSugQhzmEOCQLryP302IAv4Ntfn1FTUUrJOP+gng6kH8AbW7kd/
RxWJoIvADSKetZtQkrupTUKT444vJ7DCJVFSB/nKGrtY9xyunpVf6f1sSPQD4G/h9RAzLKNMYOw2
+8RDBNTQ2rimWuU9AKi5PXEQxMErNXNyEyvy/9qLKuqNmqkBf7V0YQkcDPfP13/I4hko3HWycf70
c/MCNQmBJiT6Bmjs7ApOwh3FBME1UsrhHUTkKmyp9UYDeoCDzK1RWGmH6nFDlxl/QVVMSPSVghpl
JQpnBcH14rwtteh6iLexvsYrx40F7LPHK7a0qD6bBqcgHc2OYGfF38m+lT6YsIRvIUhJBQ7cbvLh
Uqjyeoc+rtQp/45zxezY2sL7gBfyHsSrtqEo84eSyyBPGP5R7nj8ZRZh48jLlOIWDTVJEq3ykF58
Gvoo1BytGIAw6GvFRfeJ8Q1IXOHyBD/U5S71w6WA5D5T81U6iCtQgqfmUfQ34J7aO6WnZtn6QWY5
s5b3aQudNTKORPV7gI9JGI7CBkJZloMdShuzZ2H2VLNvNK0v3KEY5LtmrzCosR4FyKWxeT0f2ZMc
ecXQLKP9t9hSW9uEhjkUFTpvrhlD7XmYSccYxfoFdUjoFS/bCQpE07Cj54xLGUoBeEHLh0M2Wfz4
5jqmOtINM/Udsa4jtxTADc7wlwrz/ZVoL2AfGRlPXlwE+rrxLqnaiW5Fvr5K4XQ05yt48UsV6dQm
otW+GThfeeu54trXwK1f6Y4LVu2reAp++ZEz3eLn0KoTMC/dUVvROEcAUM4F7VDWyG8qnf7VRcrI
WCf6xzCfBZvFAvl9VfIiXWg+o5+6Ei1j8qTbOXGi2nvJOoGsAAGaNUZfrnqVWgfEPq2drLF5vste
qDxDYPMUoDdkC1iMFhpo3v+TkEMOGKObez8a8Y3D7O7ICufAK/gUSizALaJMmI+D0BarlTmAnhPj
vZCRJkTrUZVt8HTLR0h5xFwp9/KU93XsmxrGvyu3FijLsTS9NxAnSrqpEh+QoccCS/i6xhGwyVvg
IvODQf/WY+FXSbgiSlGnWjBn0hBYPtqqNGDDlFvkBOB/JehFhnf5NFJZIHvl4Hxsz0QiUsPl0tMS
+z+hcviYwbwZYwISSdjrb2LwFHUwYlm4H3fUZ+xSXcT6qEbPZxtS2HY0doBQ7BP1cpl3bTw83YH6
RsDgcxzBV/EKTmXfNQtqmobbUpuBUlrLLrD6GkaFG9PqPVxZwjjMBr3P++xvdydVRlXhclawwy/B
J9c+njSwuoigPBiYLxCtnE29igfev/f/dmwC/OIDkcd47wUQJHIKbB7Qpcj2p/Ltlw59OFGsuv3s
y4xXABbWwWZ8BwwJCxDvVG16jzsru/dIYUnzeGWmr3zDFHE7HbhFjaoISjKlMiA5gmkArWJUf+Gp
DS3BHjcfe9vH8UGZukm4FVfTeYtlbHqGAjoGmzRvFcvtnXqF9XOKzY4mi0pkEMiLZzt28wJs9lx1
yRkjmV1a7a4YgDsk0EMb9IUL0VwgmYE3UFb6Hk44XREjOFS+whrpmBpJX34MNVug8HIgKBi/Kew1
LZnAzMHllCwyMbrmTbHaw+JkwoVNHpesSCUCHxs9qBnkMU1Gwq+FsTXcKfajzFWmNbGrLKqi7dyO
sOIhWoFdjh5KBLMRdIgf+FKyzEMUclrULmRRFGjGtVpCXAu3c6gh+/rreE5BojHyg3egxdV/NA8y
xXnTTEjapZEOJ23sdn7qpbgqC4J+zhULYGNze6w767fIP3h53wFOVjrravzYIXOEV3j3B5Sgo4aF
aR5vXtWlxlpyQh02ygCbYOGawbISSQweL9bVtVhQoZnpjSJjM9C7NObtQKqNj+ia1NgRDjQxn7eM
1JkV52jwuRAWkbihTynMORhnedzUNiBbJjDBloCPifoI7GPY6lQ3zqEnxSfotRL9Ae+zXFcm/Lts
pb3JN/9y8TP+kMjZQQwc2BNnbqIf8ivfTq+rshm8nYoLRXjWuE8ZqByl5Bcg7spZi1GQMu6vHi7A
HxngY9iH9mYG49/X109u5bJtIM9tGvGukJzzvFQxC1/gyriVW38iRpYSz9vlIOc6aq1xGaaNyYe7
9UPSGRke4ZuM0VoIKINTPOKYuyiU+oIIv1YuDC1XF5jVa4DvY/kMQAiOMBcHUegrv6aMsAcygpaw
n4VyDh5J9e/Goz0YC6E7aAtphUTFbQAw5AQlXcBJ4lHukiswXWmIvWIdK3YgBnc1Z0+8ES5ElETs
ZUrxKJBUK5M/KiesIDjv/YITMs79fyw42oVd7GAqhTkpmp6GmNf2NRwgN1DxdZrf/7UozlUKmDtx
c3t/Nt37zFp0jF3/EZqUE/tUAtQduXe/2uTADqQhzmbfsBj9jKJLd8FMRVgtbmNXum4iCaVhecoZ
muPk24JaS9Cq98/MV15y4yBP7xittsSQTjinbitp3oniTT6AcccVeoQ5UtPHSGfux5irLqURSi4b
lDXuoMObjfuwZcNM3q2qv6XfFU6G0sLGj/ILVBTfNGmyUu7d19eEX3Vr3F2PmI5x3hbYnfaZF2rV
W79aeab6RzgENpzIeOg+63W/zqTPh48IAQ+KWcPfyawCPxUMlSbzhJqZIDtZxagz6Du8EsWkE5EL
rxlHZTnr/CxjLWR875DLiMDu53fgR2PyHuQAFOaORXCd+d+giA7N2Z6igI9lDU9kF2hwjh3FDWPb
0CSlgjPJben5j5/eHXrHqzqTLQGR/W1Kqy+tQfQhTV6c8ICAIPGVWSdeYRICdDt6nvoGE+f7/4Kx
WLNi4fhGqBbMejTqk7TVwlBhXos50Rwv8ELnmJnrijeYeoI2KQTPEEPLLrXKvMGj7xwk4qgHQNT6
peTI6ov2n9DFBy/9aZjN09RmXd/R0ZvpsYFlPvNynDmEu74L3MZ04ggxpup4sdBS1eqieKxXljHe
ZQipOSFus6yzQReZwSaf1AsjLkAJf0V2FHyj4/NBKaW4GxMHR4ZcWDkeiD2VTUIBm+8+Gs4Zgfw+
smWhySouZu+YVqJYYJ1jVY9lBtjYKEEs9cMPlB86Q+qWXwGlmQYDW/zZR6cOr//JoeoAMoCjFssJ
9soJJtNL2ehoDPRIhcL2fyzvV+RpkASvGFhZ5RyOTRjpzgW3XnCYuMnRfY9xetY/vu6Inkv+J3Ll
B3n3qS1XSfyPxdN5N/DHp3k6B5S2maq7TcLzQyrdxepon+rF+QWe2azck/hAXr3rj3Y7OZJHt1jX
YUGmoJwlubuPDIJVCxmwrROha8C75dUwYbdUh7yWNzaBFQrL4/rBCxGAirjDyYDHxJBBetQfQGTe
+Jn3O7sXgaf/WQGT3370Biw8ucL/hivB5q1nTBpSEyxJ73UVMXCoIoMmzaytRCtP35a2Gwr+lLrk
uytZ03z3SozfQSOcLW/FjExGZH8rRk8Pds8rAQ6YaxA4sjMnEp7sVgBgyP5/uDroCw3he7NnaFVU
0NOZnA2/G4KsNRo6/VEEZ7ek37Z78sNo0mYSeV8TWxhVI4mxULX+rSbEuESTZ4GYqD6NU+zHqMFv
nhh9DcLaaE3Bw+3klkzGs0MMpLQtU+x4UWTZbqyFpW2edf7zQ6Rn0pU8+wLE+qPkRkdLArFAH3Ka
yJxNdxwwom2pUR+Blc7MAq5Y3tkbA5tq9lMx2Xid5NqNZYYjk1/73mdbcy7p/O/lb+IGwRk0Pc36
VvN4USJMlW3R1kUHV6ONFI9i/W3Ac6b96rImMECxSdmABTo+l66l2qdbzueFTMfRDcsOgKMskjx7
4KVb8a5aMCXfpW4SD9VcnTb+9yk9XMZ0eA0EsISk1HYXAP7kV1Vw4ZPJC6EjWf5R42fl9XWEAD2m
PsQ+RgL0SPT6SjZEeDl64JHmieUg8hgc07dOVyC0PuoJ4jGn738LnWksW4hJQq+elEsa2Qv6Pi00
P7pMBjDpB34tDm9SQkSKd0hs0gNcdvWNL5UxJ12R3ADU01Ju1fUVsF5BjMHZVOcIFxIjVy4U1KRD
MsyKjIEuzAnXls9pQ7MKFnBXYMbZi4y/TuAnCXDsFUpksHWr+9CI5HocfQ3JXZq4hIKRMosxxkRd
e2/q2mzZf/7slBCn+rT0G6wvnKHbTeXvGUGPXOAv6SNTBSdvEvemXnyibYH+mfZUAJPOsSEdZjqC
cpKQbXzEGUUJGHM8G4QV/bSyCkK4Fyc7NqFYoP1/t19euTu3v5tb5ubs1MpxEJb3BNvn85Ku1DnQ
uQNRsQh6g8Eo8kOtCMdRrat18yHYtd1M+/zg3c0l/DwxEhI5dsIwMftccUkNInRSi8JvwQCZFsd8
+s5ZJzpaeIIdYVNZIcf6aRx4VRSyIqSaxsA5sbSrumVPxFaEniWLZPX37YT9VHmaqJ+lnO/5bGJI
E6W6RPOsbcPJGyDpa4Pc/9VKakGn/Q9O30A/5JwwvT3YacESWjajt4e38Y9JnzGdPvMA+EsqH23v
2Yvyvi0qkWQRNhl5XY/D9ZVB0enIvV8jnhLgiwfBshXBJuA2EgVzfRINw88ZYY2GJIx7ae3A2GIB
waYuNmi/9HHYpP5Mnsqs/rbkLJw5rG5MGTaD0glEtUKbP/VwX+mZhF+SbuoaeMYxH7wQvZfm9kGn
Sa+OfPgfk/IXZU9zczvwRDkBmdnS+1ioPgEeh6HJsKurZN5A/kB7TYUqlxbkuugJVDJ8n94+BCXJ
H3mzGzUy3Rw8/jO7y+hRLCxcQgBKBFGVMg71n/EPVr33z9w13EJCj8nM8mV3cvyc6vTbTQECgdUg
rx5lwb2HLEZ3jG2vE4ESwr4/k2hgumQRfYEJz6GF/lS6V+EMbVQ76iizlXFhruixR+vng8p7w/rh
DUd0xLjp49wVIpdUQAWumiT3gU/t9B9S6qRjDYV+yk3SATKoQU34T4HJnk2izNitn32gq16/k3/a
kV2egY96qvEKNQ3/DIZtPA2wP1OyAlszvzIdueZFc3y/wh2cTsHM5bxMXJcT9MiMy29R8lsdNCn0
5woMpM0v/4WoWG1smhuIiWRaz9WBK0epR4EmtpUReFUzadZILaAGGTQoeP+x8To1xfVCFp33yx3e
Y2cVXyyC+LdPfv1d1nXk2/9QqGU9Huxe4xzg601W+GxD4NKetyrSU+7PzVaxu1jTf3dUYCo3LnKa
y8d16q9rIQknEwHR8WRU+EEEE13Ufmit0GxQQ2wrk4oOkhJpa5LCtlCK6JzkaMugxnYoKzUlkXKC
1BKvT3BU4vebaxOtRD4NOpL6GiddGHQFOb0dgwG2AXhuJuK/6J3DRhwRZt5GIG7yvn0Sdk4KEdgm
UwC0VwUyNWghqt65rLuIcw0NATr7OhtgDyOLG5AZRJUtB2LOY+3TmrU0zZpogPZ13f3HYlro4+ai
K48Sv+Da42LPvvhwxbsj15y8m7OND8lrAj5HLIS1RaRMsIi5s40hPcp8S/pOJH6gOQeMFOON0zXX
syDJp/JnfuXt/AzW1YBfZrbHU6r8U/yAJ7FAXak2ttI4CFltXdvDcu52dcGrgNL9ozwRpWruD0FA
G1z8kPkKOj8PxYq3x9K3y9qIKE5keht47GP87iES99ngno9IetBN3SbVp9vgjCTqkAHdX7TGgNdz
EJ3+EMY1oPe1h549QOmw3MuEaWWuhaNvxCPTSNp+oGG3o3IuCDWo2uGTvMUz++OXAUGtz6eMipDY
kbqomiEXYkfZonqh1j7VmG41nrwFFA2GVbne7s0LvT+2Q2Wp1EJ3/AULvDnuCJElu90Bbe3fJEsv
zb1bhk8r7PRDy1OO0lN2nhMGdkyDlUwIZky/PB2iMyRpDizEFToJkW+Qfv7UBQSoPp8itwiCH0BF
0Rlkyz8i3aid8Usgn0fiJ6ORPdmmaP6e7Cz68IpjruLEhmvcnrnHE7frx6ywT37MyEWCZEepmUM/
H7NX3jGoiNgocqxaWhB3Ab38oC/5o0f7EMfF3n1BoYgq6K3yuNtbCkb04a6cxmCCzuCVtNuudgay
e9uyggtXeCQTj9XZ/66jFEP0EAW8IDifEGRKSDINT39f4iTt04k5/KamTtfwzElPXt8/rfA7SYaK
PfnBnh1+341VQ9juzpZhyCO60Ra3JPFFIfO/iTCFdPn/GCk74tMIWipM+sQe43fMFGLSTqnLgA9U
WX4i+bDdrerzq/0PtXZY3M5o761dR/+5GjLWxiLLkI/KhyBgqaIzuu2/w3fYvCxkEg3r/FAKUTAt
6pgG6KbD/dBa4LMFik8Fmpe6sxA0qZdlxsPKklbEnj/RafdiVtrg80VAY6SURvucn9lQeIuxpB5d
AWBAICUCl5jn5KZ4JDMERY1gXvjv341ArM4XuNjijhwGAG2iW02pHlZgB0WqFogEG0csqR126lHE
vnqB66pJwnJhkUU+9muSUzSCkeNWf5GzXhAsIC8YhUAU/wIYK9a+1SaCO2ZMezJkuHztP/evQcxJ
k7aI8qeEipilkDmYgtLn/LQ35YJ2GlFKbGK/d7CNnrhjnCvbCh7ataXzZYqwN0LMfjDuk1FqExCX
m6DTJZvTxGd9npV37zDPddgNf5Cblom6psSL1AymMuvK1tVOANdPEooXs3GjK5y9BS9feq7E9v+c
S3svIcF0cMCLMPFXa9c5uzrfQU4m0mfbKubTu5vyWzXNiRW88E1KRNA+5mxf1h4X/qz4VJ78Chda
AzWv1Ay/RNh37cxq8/Kw++2SMqh10rEeaMxfDTNdE4CeWDXJBrhtTLhNkMR7WX4E8ObD0xZHO8Y/
6OUFj6oAglx3aKPM6Du46AUG2EnmA875CHYd4KOMGQNuqQCiIDbwZVrmk19GT9b+/XveQP94TXi1
rfn6pwpwuhRq+ALxvpQsbTGpk+YRhhrq+TyGZU1QPlm2x6MLjAq/B3GO7um9zWOeD40/mLTi3Kua
6+odkPTzWZ9xRfZnPQG7KrDU71ov/mFfiZfJuqNQrixzcvC5qs4TGzvbqYP/qCDPcsIn1G7UbAgh
J05ORtgEbY5U26ETdHhR2wEfKNgbQv87mPTnYM2zQwfSjbQu1Iuh7h3x6g2VenIo0GQtqSnGYwDn
P5mBgVjeIhZDnCRbabkx5bImZyEyh1QdbV5pzZv9TulWJjKsEZTj/LEHe8I20dmXDefvgg8CnOZ6
XAc2BkujObbpn/+ws+ku9NoEJVX2x1HuV6R70S9d78YiHZTxYs4GeIU93osD3aKt3C7HsHTj7Ehr
v7lCjFIz3rDMox/DH35rKd7FSuxKzt7nVmiJxDHq9a0RXinQOt+LCkwiqOxo1dr0C3w1o88xB6Ep
dvS6HppA0NxkPMszl/EJxjHpSI/oJ8J7/1H7yOvyMlNc4hFLRDN88oVovDc5npwzds9/nYQh6/G9
yOIYA1l2AFyRd/uev0m/dK5dVITvj2MX8QxrlWvwKLqdV/oDfuWNeLiQxzFoYiiIwyeofhhwr4Yv
nEVNMTOleI/dce8Hrmwi1o/enemojfCP7bMmx+P0jCRDYmlXgAmTDX5Gbi4So462sP8NPUf/e8yh
ryPRO3d5rNuJRo3g79zXykY8ehtgGVjDqeBemPScLxJpNoPliWdaNHU9go7CUcXpjwelyN3PtgOY
E8wioZ1YxhBcbvNpLtRtSULmX66+WZV1YoiszU0lIJ4hIfIIVhmMzGO24mFTIb8A+ArFguK9Cf0U
sLw6VVhyBeHcpiw+/2/pcrbZ1fDeicdPvgaIv4HTMTPxHTMvelNYnvztvwUP6ljad/ArEfr0aaOc
UZWHjmnZsnPM5a2PTzE5L/7jlf+uMiUzB6T63Ke+0ziEPbwH+aboDna7VTDPFIQVRkpwfyBWAS/m
ZsVDOJ7e3HJkZIVoxA2y0Au/jSVHMj6RPYA/cv3pFf114rmApljkucgCnnm8Svl08pBxtwuxdfqf
s2g/adbxIos/M6eSRtt5wQN0qjw7uoxzFXuyH8kt/l19pR1jxnAcg8gM4+2XvhXki0N83qMCTHgR
xniTXq/oxWAaly9cBzzIDw0gYDPFS6VgI9h8rTiMtTw6hePTiKb5KIdgMvKSEvqZhse2ln23Sxc3
8uRuWBi7HtYGP/IR2zyTd02l9RxGbrfooRCi7Zz/458ONLZYOQLGd5Y5GO5ZCwIX0ykTM95vxSty
GrrRrdumu+RdE+QCBtLUkMD8DpFiAGuCyDjvtQAMQ7J5juBxL2NgzI7WLYj6N33TM/QATsc/BiSG
1gkJLUOdyUrQk+C7c5tywViK4CqdPpDLo5CBnjlMpMB8DDENbNXodLrUW4n+58C6Wx6HMvuqG1hg
pHGGBXyBwpCSM7c/pmYSidGX1oeWAZzMJ7TyVIdC0otEmCGmSRQOYOPdq8/oL7w2wdhnEIKRP/89
29MUtT+Du/dprnUlObbcxRDvWY8flprNhlWS7pzhoYhrJJIWMAxof8wBQT3hcJpCnnVWU11hRr+O
aETb4tsDDBy/RCKmzpS3vGQl7jx+jQzUQCXDq7NsUEZyZjP8GsfDxAQe+YZzE6BVy94m1yCoMgO5
s5yte46oFUFORnQzyROh1DPtecYjXgC3/jhqke59UHFUpfzHB5JB2DK0s3cB9P1kgazorLIS9JUz
U4s1dCFlY4fmBHctFCzTCPVvcm1MrAmPtGnvIAujF6oFhwU0dvYr7/gRybPFm6bnMqhC/KlVQUBX
Pf8Quqah5Tg60ZLCopUPO3qKydcT5bO5Assm5pcwS1n9rC3VTZPu1IEgoCyvOmoHEksRCpjb+gZ+
lpk2mLbN4eUC245hsXpCjz2trK65NNJ8nrAJ6ljyuBugzY1iHqsP5O9mtw8ih3tGtGblN7Lcsf5W
hh6YeoBiCnS5bOvY17UPT8YQJm0raHUA21npC489AUEheKoRj8tYHlJxKv7paY6ODV0kKkFPGkIA
xTWfhBI6RiwH2RizCoMER7IHzsQ73ITQ+g4JHPjrKHKslYdEkwGQ6/AtaAV6dK2wGpxfFIfXwvN6
08UrE3Dz26foEut4CxhdzZ7OLu9K3b03ZPnSfEVw84YvdfZL5HGImBoa+lZ/d3LWUXt2O6UvCICi
LWge2FTYPmgKt1Oyony5pIw75JAXWng/CbqysQdUetX9kv2Spcof4fukTgOtWj6vtQ/oBfpmnLPM
uYd143nE71v/Fd21nhlb3oi8eXWKdD2Kl6wVqJv/i6GfG3bWJx8+Cn5slWdYqJXbEyl6znlY8qNQ
oPFAyB+IwTh7+ygGfWIOp5Ei1dOe6B5pzihFgivhwTVYGfUx7ehhoX+SEuqi5a4yt/L/CL48eZjU
bngWzNUECGhhFv2gJO2NstzkbzI+Z9n4T8OX3RxBDoHMDGPA4k3UYP0yS/w1tgOsjTo90gzHhTAa
ab7mAc0dq7SY6C5Nr09VnsWLJxKqA4cvFCz+KdlGa/BOD4rGjSoIbvc8XmXO2XZoXR+8qSl17VjI
41nrLpmJ4eovepZ2V5l8MRTbW0qEeVLWttTRpxh1a26kFTMatoVdb/TrmY3YjqoEtzGXNe21KIic
DQkEANROarcIaScoAYjIhI5P0iMQ3oRGfYB29xmv7jOaUbkHJw8uJidhXVKuaYRrEm96T4kkFdia
gsuZ5CWAAfjr6biFZrMrsKg94G2RBUmhYoBtMr/Rm9cFp1axJQ/1iNoeFGkml1Mwt+eThbriYOSC
knTXtCqdsZXJiakfF8/zHG4S7wjnAf/xLnIPLdhYOP8EWtRfvL6NTTF/ASHYhyHBGblrf/Z25uBb
0R+bOj74KUa6poiryTe7Vz8ri/E1Fn1xP+YzQ6Hkh5foudvurXfCsYTUvByPiO94cdNnpECwzDu6
jUJ+mGyyLRWZ8/JKpDEAUzrH4gToKOf5+YStDpMMbVPp4NEotefameaTH+hWjd9aTB+i8CFECTvf
/1EeZAoWtHxjGZFA++RN3UWRz/A2VGvPZPJW+zzmUgg3xLn3XlnMQ3JexMzteXyKT+P3nH7oyJnq
ClpMfqxsPuIYaQ1tveDXXahzdvDmDXTIWopE+AB7lXwKUhKafXv9pltPeKnTxFeGR5Zj1qbAdO1c
tNUNSMXjFqBG7Az7G+BR4RlJSzv1yBZ2BLa08FzVi675RvdXiLrxtcED/81jBsrvlLnyem2Irdkx
Ga5g0JMNQEUrTPEgiGwRse0wv8ZR1J2c3k4A8IAZLNANLWZlh4bOwjbLowMVlrthuTl/VFqAceJf
/gL5P6R/Utr0Wl531GLP5lcSojpOlUY7AWPGWuCfkQoohmzp2puOzzGr4ZlzXWzCV21FDQCWM2tC
fiErvkv82hdIs+AqpsPZN8cznh/sOW2H5IWaKkz6cI+SXBC6Y1KkkOasp6hSV8Q8e186VGBio8rF
qLl2AcjUZRYw8678yicXK9ciPIMxDZriInT59Yeo6Ov4unipGqufX6EQYA3tr3N5SuZFDIbnnqqS
zetwoNjMAbxdG70eyG8K9iGaHD0ogwXoAmRPYoZ/VAb+q3ADaMLzXpXufUt7KT1UQ/SfnZistPLm
yNRhSs+FwFbaKEb6L2DDS8pN5XYTyt7aEchuxRZ7Svhk9zEa1aYuvRhikrP9FY/4mXEAfBQ+Vc3e
snXAjswNeYyenNtybCTyKrBE0vNvGkGeGylANRVyPfZ/3xTGK3NejSfb0ZK3lxIVhnzWiFqlt/ya
Pry/+B7MLO+ITnbvt+yRXQSfWxedXLn5JiO4CInFz0o7/gDZqqg6VFwpsTMFyGajnj5p+3XW3sbz
dVITrGRNdVHYp4NidjhiJNFvNvC0chxUIqZ0xwykanzy3WmnYw18HZGtJ/Vo736Y3ChrR5kkSEwn
dVupqDRWJb53LR0TkP1BUTPSZ9jDs6+jcRQ18kZADkQOwALULJNa9G183oY0E3GtPQp2Rt4j1CbW
LXRKqlvvXv2Jw3JKeMrB5Eil7agJnbFVOoIN4cEq/lyCHHxYeUOj3HVAaiK/SSb0u3N8EV1swGGV
LwjsU2PDXqE062JEJetLq6U6yLzyFL7ti8Csgzqe1Gp896fyrJbwNo9aoSwHzHUVKHAjtYdigWdb
iIUyJgZZXHpJTM0YUiIyZMDh5wA6kfWUPWE1WtUhz95sAmBci3Oj1LuwfSCtthfMhX5ieTPFNF2a
YRdpsoVyQekZL741TrGFAx1uwUFbgYjIjHGWlnhItTEfffvI18LrpGt8wuniMJ/bkxNOG29ygTfs
F7b98gxHD1DlwEzbVsEAKCtUKw6408nS770hE7x4NLt0sl4wgj+6QWRqXhGOGpB3e/pUdhFIBqmF
9ujr9Su0S3cizvyNuRwmdJFCJhoNKBDRftsukqoGcUBXg0BGk/C3LxV/Ws8lG0u87e+Wqi6vyPHp
wOEisTI4RTSy0JZKP15KV6KS2R4C2T4Ctg8d6yrHQ/f+Qwl1b4GrU2lAlipV1N7GtlEKUhaRfMjS
NUsfnyYWgEkrwIk78CQ/4P4V7NFRCC1cFjH/nd5/AwUuweFgTDKSj9VWKKMoWPMP78F+KVKIZ+NF
PBrDzrpi9kPXqUsloKKX435EPJj3EgJm7fsIABwa+3kFDpnRKLjZmu4zU7/QZICihH1HhZNTaffF
TUONhdXzB1oOnEVe5XFIHsdhd4tX36vDjFOsC0K51OdFK9DugcB1vKpum3Eh8RrVAaPCNYEdJUhG
hSQ7UVVHIEkmZtFdfIK2uiGZeZgsf1Fvt/4v1UG2HI5fmrMaySRq0Zq/WajuQUWA0wneyg8Tvvfy
7MpWe+0UfUWsp03sKxrB5Fr4+5F+jrDfQgg66lUBCWBYUOhXhJTLE97cOZDQHK3bkBMOKzghwjr3
l0iLn3vZAV23u1KQxkA5uW39CEj68nDg7Q90I78t6WAZyq8tGeQv2SJA/rXE19wsPQ9ZqySubLEb
cA+fu7h/GliLIKsllz6aBkRZKQCUgs8xG4JivFE/S0ZbmcO4zdIbZhRAN73bwXWJuzPMcX8biH5z
ezqaMHT4+OSZszr7f1DnWaZwqWEQH344XzVcB4FjYoEY9DG97qr3rDpeXo2tK2W4+AQrum/yPXja
oHDph77GjkdoOZ4646+e841YsQDmCLe9vA9V8ovrOU4zjmyGg8R32vhVazxY8MASFjkKL/iLItCN
FK5RQA4cOJWPSjgb9q2lDI6NdYKjIuaWu4dg2Q3aja7WmC6ytNCnFhZ3VgsOwqcA9HvAu4mQHJxk
cV9uPVogIzqzPTqkylrQ65QZa++bVH9K5JQqYfoAQwrSvfowar33ZQxjwPNgJmITT9nXF/SMhPGo
5tc5+dYJKKIGjWxFcZOTcDq92Up4amPcH+7LSLfo/aW3aSCQNo1LG4VCTvG3ap7o7GK8CB2XmMch
PcLciRnfCMEZXLqhROaUhJ5OJhKSCcajnd3HHsBcQVQ0+83XmWb8uo3zovd0bbgz/t8Ru07G2pQb
6XGAC1axo5XwrZs/q55CwT8FKnku/vTRhFbYU/vEH0Dw8AidglZzQWPTVM7NGC8yCgLG17Vm7zMf
dy/4gq0ge+Z12IAsV0veWIXXxN/7PZKZIPG0Sk1YiGhyLCR0octUxwMTNq2gZonHFMkRul9n+UbW
JcAhKBAPs9eqTScj5N4k+ZJWGlUpEXa3zV3oQ/IwKm7+CTAsjQ+KeAVTUkAsYW/IbFPf3s0cpkSI
DD2obLJwyHrsm8sclvU9q6Nxv+GfpmwJnb3qJefZd4liBG/S9AUCjSbBcuke0UMrXV49Zng47XeH
K3PXFPHtc/4aeZXTPjfFeo+jfPYhUOJ6THWXw2/y81tGPuju9huv6GpTGifgoAHpImMnVZjBMcrn
RO5RiHs0g1MnIUvGNg2MVMI2edargmLU4/RvQEf26zeI57AFFJPRm3j0qQkwVU3msQXmvIJ0N56U
1olBfBbVLTTX8t6euYJnq+SFTGJNXj7jgSqMF0WlL/pgyf7MsSz7F+TFL+9AgBIh/ErXY7v4f+4M
8R9p/WLdGWF8Nrz6ah7r+mKOFQm5HK8eUNdoCkFCKCbtTtNuNaya4lOxXIyny85c7C8n7kEIYpKc
VaPcbCdGizgsDfEuTYQAII3266te+OAJHB5W5nj4/Bj70eVeJPtNpTJ2ffpBk6Wb/J3fEpX00hrT
Y/12hSS51HOYqmPztIFL0nbZNPA6D1EEeFUCfn+31Rm2q2udF0ic9IT3cq8551mr0cTtPHGjVrVd
V54Mt52Rj8f5zcpgySMarxGt7z3oDW42IBd7BA2b8j7ZbXqcOUbOK76QFY+wvDnfuMtHhFVYfdzy
NPbI3jymTsSOMg6C/ZMFdxRkquQPOvSq32MM18y0+MCoKfIyypcXZ8ZDUoq/Mb6UtA0/4LvljlCl
w5fsTittiP9HJIlN14YDVi+jDmSUBmtg4iY6yceMRk22DgGMRPxZ6DUv0dnw5etHlhgDiwWkWofo
Lcz7lnTgr5v41OpkH5r0m+yRjIvexdY0ecQlG2BBwcG4s8rdR4AC8H2bR4BOqj922iHHw6Jahpy7
YcVNHCV5N7sGiZ//8ve7+Bo0nZShX/YmbEGql3lPgQynnDaXY3iqIzNITObJ7g8nnK0iWSL7sb8L
Zc0AzjR9nIksL7s9RM+PM6xiQ2uDv2TztXIm4AIpAbjtf83lWcntiQoijxy89ZIvnuwTKJgyCsdF
a8rGkv5GiT707QJF078NGfcYZucLFqCqCUlMO5g2g1p+Ve6LK6oT4HPrR5sUAg+pPQhMUAU2KdCs
b9kpb9JpxzH9mbFOKN7BkvVSTqJM2hfPXinO1kEeb8k3m9x1c5Z7N/OWKEPTBS3UsnRnqiaAOsDa
lejmMQmV4P1iZSNMfXGmLRYe2tICOiyur9qb4Ay8USPXUM+qmU8d+jP4AqlSzbdX+3gw0F2fqE7H
xaWs1J+v13iueqP2mx4+4cAnVwnOaIJ7rqgLjW+QNdgnieYhof8CRB/IpZif+GVLUV0JPFzuvF22
f0Kj68XBxjLkPu1RbIU5Va5NnXKJJVwTIkJcKaUSDWQvIuEUDEMgacYyb/Hef5Dhnbt2B7cFsgDS
KZLd6HsFdsy3ZM/dbxs1DJEytB+vNFx6rZPW53GWYwStItbXWxn6ueXvcWKNcJhfgbmraY26FkXh
JKcjF65KTnZJLt84MJwaCJR96ruAS3ZaJxx1pO/MAt1Lz+U48QSYuVB8VD9lGPagUNzxcIzhpZm3
73nBWuJEjbnV/80hug0NPDsI1kRNc3LQlVd8rRr7Y838vvvtPj1+I+4To8wYaGaIhtwj00trO+nt
bmFmQG2CO8tkwwPDT7/btm6oWqUCUDHXlSvMQv44FTeYcVcVTlMnsECCEcZoDp/8ZirTF/N77xHA
k1s57mV6r8R/Ps10eaEmBLuELXT20+kTS0SrwhMcyl590zk4hQZeCS+Mb95otcfYT11/f3f6kbtf
bhjK39eA5y2wuj3ThEzErdzb8sByyP0Ltdc+sbc6HzLUNaLI4gBl61G9U2p/s5fXmOVOl3xStNxH
AzemWa7dKRBNYVwyRE1NzvF7mNEDQLiERdAAmYO1iRIeejMEBLQSoYyUf0lLnEPf7xZ3wOchJUTC
LxtkDUcY3+eBJ7EkRZ7C4MjO9KSXLE7BaMNRYVCY/uWNpYCjK2UQS0ukRhln3vRGUOC5cn7vnyb9
m/X5BKxo6LZdOWQxJL1JI6TXzlhH33/cY/XlzRgd4TCo3JudfSVDRs++3SLwxPxLA5UOlxSwq7BO
hAmgIiX795Qwg/QyW0fUnTyomLD+GOIxO9XYsAgjV7GoBxGg6cgjhZDraImE53LqVDXKJC4+pi4W
5j2HN//Pz/Dq6H3i+dqwrTfrV7xcNbjWommyN/Dide9Nn+IpbGZhWU/t1h/oupmqJewTU5nXxODr
xvOQEfLeCt+KaqgZhfZSUjkfe6jtCHS2ngPvbv8mJogSTohJdhut8A6WgUKS2Q89eqDoAhaOYSsp
G4CeRdsWHwCROTffCettLwfHYJU1g2IIjDc6wQyGwvF5iKFg64Bo94VAC1uh6fLW4Q3Ri/mXrSSa
CsSUzYsRkueps66NKJPJfsmk/4CEvFr2mBgap95ZMPwTvpjp4JHnM1ciLD/VHNhmul2DuN6WYaJY
9+7N6FMR5WP21HUMfb2md9wfL/9MwE+2r94v6GXqgAsGYfWfBHMotlPK/tvM2Zh/SIq53SWN+OUH
pFDzWiGGdrYR9qN6k2u6SlBbhdUSK6fm3LvnZsaDKupVSM+yMX7MYPLjxw/tpw4L5511Dk/KtLYe
AiS5DgNlWFNQsBYuSucdLAxi1pFha8lJB1umF40xLdiPtl2iEpdmAOrV6PxrDicONqdsbuihrihq
EAeMTaiOINApJ4SSDKcSrHIlUpJExv+kZEgvrRb0m/jofGw0wdHxj98xh7BdA+PRrXt2FlTNpBUk
iGiZvfJJp5kjBnfNUEufficrou5DkCCkgj2hOhVkykg4pxY0VhDWrzanxtvfeKZV1Dygvh5D8MfD
VPWBEcEIDbsCGXJO6Z5FhlwQsSKwqNDCVdcvlsVJSObXh8kTC04lYKriQPEbFYH/Hh8Q1N4i7sAT
QKDbjT1MY7M6LB5n96oB4vA19MUFwqClJbgnyfZ3bTkGGsn6lI2FlViFSv3Sitnv7/CSTnuJ2a/P
TeN7uZeQZP7E+w6oxoGbaECe3cOL5OvSxpF/7WoTRnmCxeWWaSUhiUvSZWB6aI0KXYQs9Hn0ab5/
K+L92dxBbITAyJENExeyPp+4l51N2ty0K0/Re4bWZSIHPK/EPRDkN4bGunnSjMsZ6/nMJbdVZ5o8
f3VKhP6iebDAoddE2yglwXZWJayTJrnMsKrIyR8tx9N6y74+8BWScwZNEv/ZXKyIig1H1NtCJHvg
0ag6cYWvRhUesRFNhBKDu89DocxwGbhakoa/pZloaJAvnTopGq+vR0Ryv+wslgp0LDGINNyOWNlp
lU8cL5aCZWZw7mcZO39sqzUMuJJtxcCYES1bmoigBdoVapqz0X+SCp20/YMrMabfv7bwVfrfTTMx
c2f/AEjdUBqV+LKNmMTZMjh53cvF829qfj+FYT7j2QMjcp5KEb19SRTYi1x5FBiGkUr6sAB8yZCO
dxOR/siwtXD9ec9FlzWwh9L6K9eXFz897CQZ5raZaCMqObGkCj8SRmO/WQmrehu26sBuhOOnobOE
PI0UW1vVrwCq0NJ+qI9EWxj61L7milBEySiXjC1n0LgiVoLJ1AZ+qXX8lnp3f4ggnDsZ6LVILrJP
RwM16roU6uGRJ2ZadWSSxAyPK6ge1lVLItsBq4SAm8QA4giWgew0NTKZwnrDvagmPKsgK/rwGVer
1HfcRYU3figW5bjo2m/isw4+XoeswtDOuVfT4UCH/tiraTu7/bX+Kv8Uoe0Er2WOYQ/w/rJor3yR
auDXhvTjVJqnRqZGWHe3Fv80rFDwC/1+Vg4HEh2hZGbGS4eDRW10gkERBf1P6Kt3UjCv7qfEzUlB
48EQ6Ue4bFo4N95pKqN9ZdfQ8Ru1JpJAewsWoa79+WjyoGWcaefsnlbnRQRZjnOJ1cUt8cpP0NAW
Ip75hxatJWfaqTyk1d1AVRXd8GiV7PqHKOopIdMCyvyrENF3pzf6wzWksidzgXniDScJyaATs0TT
I97H6WiHcRTmnlaXYY3gr/9VdUacCU/UzjXrmF0irBC3ds/Fby3M7/L6cTwJxO/0DKgHzDI1TBwF
u0iUDV9iHhBFOxAlaiGcSW2IAYfukdJxmT2hUmZb713cFyg2K99hVBl/KrfjbmPqa/0yCJAe7Udw
HuBzJHTAMRFIjk69YHF0OkbWSrZVxZMaGP/AklMuo2D2qx7S6gtuQXZAyCYqSlpbokIe62PjsVmb
YgPq6XoRjrKAKtDgheNPH9y+mDUd5v7y7x4kcd/tS4w41+PtGOB7Y4aPn29Pk+EKkVV7ovyXzzCd
oeYgMIgTzQYzE/Dz/Zs8gTCjNIm8fDCVgIryAJaU43yWSdc42UPfpezcotMzkTzYr98+PYp+xfXv
GWWJPiHrfdN0MKE1MJwmkSGrwnl+JAgHhCIBOYwLsqOz8tBAkgvbOE+3aPlmTwo++ZKetE5ghr10
1/Rp6zhs5NK/DF/dj8yJ0r7JXLbRLO7YtJr0cbVUI+BXr/Ll0E17z7kkLL3KBvOWCn5/5aiclfIR
rGmiNPcn2Vi3VMI8Cvvsu9X+VJHQXb+pUIFrE2f3hUFJbIrkjix6QptTZF2MWi+lXB31aTFe6Qaw
oPHBWyKec+CMQUNU+b5YatnfwqcBR46mMF6ST33JjU3RB4GPT7FBf5tEV2KPRToJ7WJTNu7evXup
Yx6Bv2c8LDidL+f8cvJiceJzexbYm7RJw8nTe1FLxHtDHPwhW79fJY285IN/MBPkbtHWQsnxE1Zj
2FBjMguDPGM5NbJpYnrrJ50DnHTG+2lSgoybc9pX5QaWDsbhjf3j+xXPX2d0e4HdzEvGXF5RwJja
X2iQ9LJLxU5ZaFPtTBv9EY1xU9x/ilnh3nCYn/rcD7KTeS9e3Kn669L9OQHXjB4ENoLunOaIjQ2q
yDDrHp52IWf+zvM9CaVubJnLQwyKsi/41BuGe+vBoGDMpfZb9Ls+FjUOxAlN80dkPXRwXIt2YPFY
9ruTuxOg1wPMg0bl2OYpn/HMyX3ilQEylVcoBMs1VQRPZcdFiAZCd+XD2qnpgvqgs6bxRH93hkqK
Lnp6LVxJ/mLthm2gQ1ynQPeF9LsUIGFzHReqfXIM6V5j0XwmDM+D0wYKp+SICeAt3+l6dQZ4Gq7b
D7JGv7aZsuzTfb0u4LVF4+hVl3mLqpxaWlYaZ35tR91cGavRrOdu3D7KpUq/YY+NoKmJOCbOr9s+
bucd3Hf2OAEw/R77uSwSqFng9mHFiBHyZ1lWHNiXG40JgjLyhZE9lcoeWsGy67a6QOp3r8FXXaly
MIz4LsuIweXnjti7hp9Ig3vboBHN5XHfUk6ESb7kImD8EH11t9YUdFzmaS4NXv5p+F4k/o3nD/Dx
GOz+12RbZhtQgdZM/p5bf3wDv0Y7ej22bc6a2K+6EwOE6IwhFOJelkHivo3bMwFeQiqRAnSShMEA
+g8EU6f4L/mkLAyW6hlqWVhAwGv8RLqnZb2/M1COlTZMuFB8+s/F8aFt1x8j9Ov0Q3mrWXMJIcwo
IHWHiczq1MkiuYM1UfYV8C4styPOMeGfObclJpBe0QR1510ulKGg1fv/dES0hdCQBilVRI7IlXYY
hPE3xUIDSVA4DhUHpozKQrRxGKnq4bzGabtJ6maapTpod4+8yxpZJ0pth9plUkylPfxHlYCn9GQ+
0MtgEkXNJ8zCqJZ9OEGj9qNgqWXHat8H672yfo8S6f9yw/5z3lK4N2Gw452eWPxQ0Ebr1vOUnl3B
oEQQWSXzoTQFYchDtzUKPxAdiwTpr5lEAhYEfqCGXEpNdqNZsLIJlD+Jy8gU2HlsRrgoepUGYZX2
XdDMAeTBx1XbUkWGdjSIMc4PJv2bFj/rQEmAM0cYXRT1zNbeBkwWSUDfRFVgK51mjAPkzDIrH7qd
jnqkyKm6yJRLe7088jDVZpZCoB10b/rc0wiyJJxarUrBFUArdsJDXz/P2KBZrNLLmxYr8ePDrifs
5Si8qankZgO2IS5nfrB90euMTVjmsb7afDsRdbF7fotKdeqcmmH8JtE2PSrOE9l6Km3/95EYXi9q
XVeDPyOofuia/qt6E214UlEJy4BRJhEs73Gj3Iw/4+WV8XKCJgltOU/Qow7ZK1Mg3DQT368Aansl
UXx/Zyl1W/UhoGM+HpUaFTh6faxqtKJ1VCLJtk7vKRxyOVTxGkdCsO+isZLt3Rl2tWBhKMFNWvJC
IVxBLPgp3ekVP+scWTIZAND/1sgzC2qjqjtFc52tFDLLx2B8FYNfhNXMEB+vKDsd2njDc3ovGgBh
SkDDVr+Js9AEVG9aDZWtZYdQi1Tjgc5Qn4kEuJSiokyVjJpl5lBTNYYVWJixTDe4Q5C7TRiEzEmp
xwG3ikWK19UeT6/nd5ONAqs8hg8ydCkHRkVUhzk6fbf3/Vg+znbq0eShnBs8NSA3BDo5srDi+Gro
iW5FobJiR8aGKysQvebln6yeT3iZ/+TJSpemoMDIpLkpMY3/vylJngUTbOs+XxvQtCzXFY7Dk8eS
qw6zgoEC1st3TpKFJOnXcoRVxFP40m6hHFcywmUo/32HVILBXxc38fUgbMjRa52MlNn/dA8H9Olp
6ZeWU9meSMoThaxc78Rg4RQES2CB6xig8gi0spL+mj+5H831PLeqQqfMCiCdQy0LORN1wXTKimtR
KFr1eQkj7VoETZqiaAcHODpioO4L+Ww7rpJmdeJ4j6QSk3wTWeBCRqxqq4DM95ynqzTjKIUwGFS5
X5jtmL+VyTHddqLsdqPgpg4GwnFwlYu5zAzpiTA6p6j6brUIaR0xywXaQS30DR/lohbSLvfEqpBS
GiZEhDA4MdRkPc6bmZUdPQW6/Ooowa8pxV/JTRSNDvj/PUs+fnnzkyXk+BzT8wbdUPAuXCMLglhH
201n8sOi1wgVOr4N/bugpx4zkD955A/iHKjMPnNS9PUADZNGb+GkK8jle6qBA1NM8DktWrNqmvVv
4nd6o9cxawQmqO6OIyxW4xNLeIhhWtF3Il8r+aXkgSCNdqFl9ekTrSnY7zYJ2KeMsq9/MCyrBj3S
qKDaqErgHf9KeKtUT3Vb3gYUxFmNFiHFgtC8jGLxtdQi0nMHg/UOvvDUSRA4XEm7lSGlojb+bRmt
5nEW5kxD/q2YhLZUSQjOhyAM2qyyEFOV1f7cTs0rApuSKsUX8ym1+Fp4sp+TANsQ9HqZEmmmqIrm
gkW3lHEeZIPn4RedkM9bEHJCgMw5n8/grM+9oJWAdBFuBgN1FAOTDSp3Jfm2+g4BSYgr+5Y/22In
yMM2sOQTof0dKKFXylV0lxeBskdPfi6a7l8HFG0J4Xl501zmFMMX0v0P7lZpDN4iP9o9/n6AWUzG
M4zfWw18Vv9M3EchbS1mgtbQF4uu5OnBv11AZg3DlASI/Dk685tZjmWAzVgz8BIYB0d4urI4dMd/
D3cQUxPXodPTvChpPQecQ0gNizUaH0HdfmZPkwtJuHFyM82wXsSEUFbrnu0H4ZST7COIjYJIk4c6
2rl7hyFSV+6YkOBMaUA5SIC6YjXNZC2fGdiCqCdcVyv8eraSowvoA/kQDRwgX7gFSltAp0Il+Iu6
mwEjVZ/KQLUnvnrNMkridQJ78DKq4v+0KK2xGf/DK6epgF6vfoxv6Ba+xRPxF8Gsp7IdUHOKg6CG
QZ6etzgKuLCFHO7/b/E8JBPn9xT80Qpl3Jyz8mQGcFZSkXJE6zJf0YzTjC/dt50b/xyyzxZ+/7oA
eijTzmM7g7ExQjFL1pU2R6uUiB8dhZcdFqh89173IBF0ik/Crvpu6qRxc3OIkqzLs8oHrusRXrkJ
oYw9ajmEDHsBM17MDL+cemfxzaqut9Btlh5faxiif8qmVbKCUFOIULZKzWgCX+zNoKq5vgdOpBtn
iymeUfGV5eVDvETljV1onl7Esg8rZ4s9w0wOrRQne7dq/0W6mw24c4ubnqUVU+gXSGzfOGabcIWU
MdINHN8LffCecnaqA88HZnoJoAcoAPgncOli/3+kTqsDKkRIjUfnCmWVAmxrrMZDFOCQPu9X9HyA
ldpcqL3vyLf5gWkO+be0tTyLr1DCrDq/78EBVcUe8C74+gnnVzudmmmOK99USZ3HbatQA2kFqOAV
friLJcPc/u/UQ+qNQVGI1O/BhzTgORyQr/MOwsmzM2bNncOdwHvZX2pXztfdqEV42AYSbUsOruqK
jVWf2Cw91TApS6xFgQOHxOhT8C8Wgf6iE1thP1S7M97eMZxPt/0Q8alfD7ycKQlsxFbzLnZcE2FD
bIK2K32P9Qqdm0ypsHCNDujkO0b0CIRfora3r6b9/jlEBwacONuWbB9vwZE+lFUdNXg1Ee8l8sk8
YldH53m48rpDUFSowQDppU3yQbdsKFeWdyK5oHuGovOHH/DfY8RxDQsZ7xKugusLCCSBLin0Qa33
2L9FPhD/x6jFqPwj3yuSOhXaEi5ejAjzywHPedQvML/+JFotan1uUZGpxnIZdsBxodqmtDdgaTLP
L5PIredusigQ6mUNyPwr0GjMRXEHf03JKpNQSNq0bP0YqcDaUYOl6xm1xOyGGBjHwMWDWkl27atz
2lFaOgkGXbDFIDvXofuouBjt9o/aT6SB34oHw4/GNIUE5KeczV23G2k+VXPGcfxbcKiuv1za2IXX
EtucXf6+n4JnRFXbIIfYhKa4iEcp2wUs5rMl298JN7Z8OnEFRoA+34ZWdeZAQ7AV9Qdi3SsF7cjp
qD8F9x/tc+pq2DkbK2Cn/Fs0TYXl0eNcEwNF7iYbQSafe4ktLqAh0gMTsMp+msTOwDoMz41sreex
7bhtEo6EEo+1nwTS1q8nNF0OWErqwMnL0Xaagdxuo5M77f65m17pUHf7FrltKKPcxV9CVy2g68KQ
oNvPJpgcqMw+gjgOf0oHuKsMfpxUHGLopab6Yx1OWOO7pBEhoS34oqp3zp/rPaRejP5ioDomfxgQ
Q6WInxO0oJiJ/V499AerZP6bqMrLe5jlyWeT8/TYGifP/766xr9Y0zly9WUAz5htBqR3bLYzZh79
4H+lGQiWA79kWdyfuhphvrxTMiD/vdylMje38z2gKgvWeu6ERmdYW1kVO/Mp3uXc6XGrwihgh0VO
7FQKH3HpoxLrYDU/xfF2caJcnWCk3WtvXz2oURHvg0Pe5dwTLl8JjxugfJ5C9ARnmGCKmisLwjLH
G9gw7EOzyJmkP176ETuXSj6yepObVHxBpDmMjHbSLEg823SpQTuISos75QYb5F2vypEEcnf2kGN6
L0HJZbp+czLNVMnTlBpC8HXCh1AuoWVsEZNuNoBEw46Zm1b6Fn03NDhF3EuEmpQ0y88OvrlmmuC5
3sCLmwQrZnoPhUOvw3gQGZrZnZz63oCBNX7+pM6LDiiW6jiyDIkx3LIMLK8PylG21sz+MgOa2QdY
5ARekPbbsLHCCITPE8NbVbVmQYKpMeDJw1LF0UzTkNnt0UN2ggEA4iEstjdNd1Pz63jWYNr/tlwx
2EqdGRdcukiBnIyMFJY3IphFsXQKHyhFMYjazBNscG/tdwztXCJYJDDl3KRRMMzcUxAU/c+9TTI8
IA7n0x+3X7lL0nALel9vJXMdy7/ggFMxK5TpGGkSkDhIJRNENsUqlFVaYfjLKhH/sHv0zTyUEV5p
AvvKNxO0B9QgKrwcfoSYTHO953BCFa02IQZG/eoVOHSqUQ6SSZW6S9pzGMFd6PmtkSeGOObTJwPQ
n6qxmVl++ut2rTmp0KQZcT4wWGDzOcpHkeGc+c5zsPyhA/FI+fkVBFH7k58q1lTQvhQlIeAgIxfi
449aHocUCIEkO2qEjt3TZLhv9VCEZZG1/C3bt/zPcXdb/4hSgVt0Rk/x0JqJA+WYrTkJjgNgbWVF
L1IPKTLwD+E9gA9HnMmXfnO/bh2xqPCbpp3RDE+DfSi40JOn7p9y5n+wjqfHJsfxFdWvhwvzEUJ+
AfJyg8NmUohQlE6hUXLpGqCFXuoUu/7P654Sr4/bOcL7l5lXTS83T2tgW5N2xgxdfjapMLSIm/WB
upJgCqfn4txrZFsFEdxictez5i9ifPUTuKVxudR8h3Q3ch2TZ9dvYfj+3W5vIirvpg+QITQ1OXPF
PoSpInIMDjceCNR1CvskltdjVIY1Sft4wDpqyxn/6q7xKk1OqE7xwu5QSbPb4kvz3F1lcGn+vd/2
F7eSzA/H1gDeVqSp8Pn1K8qarL46MJsnupn3roTX5+EIfUFxuDLZacdCUxHlXK490JfescTDL/kc
Z8JGoIAPVDRMGB+bxGD2bg8w5TxxehTRn8+CnnZxbpqi698l8lhgNK4JJcytuGQmvKOmrK0zzjS9
YqRYCF7T/LWe8d2R83AH0FCKjbgrPtKHx1SIDmcCi5D9mvpBgY5zsb1KtRV9qCVASwGqH3P30//Y
vdKuQfKxpWCtHmZ8n20icoJSA+VUJcCh5DEFeFyj29jC+AlliAJxw0QNswh4kBhjpj7AFsVJo0xu
ppsSFPitvbZA5qj6e311O5hJQkaU8xLvBrdaH7Iu7jtqAMNfsTDOkqImnJNV949vNujQ9Ml56Ftz
GVZoMfr+ZVTDqqiWr77Tvrf9ya6AS5+PRegm0CZ3cm6tkq8e4w7NsRIk8OJES+10DLtqJj/rZu7e
kvXqj4IxBQ62SObsPlj5pyWi+ahMtIrkX1n+kFsu5YwZskvecbjnyX5JLGAU2II0O9pPyjsu99l+
0ThqEYSfX1DrGNl2rONvXGs0betQekFvWA494B/8ixuQv28ssV35Ef4J0WU595shNCovmn7v16wK
fmNxUpJ/sTkgEqk6cmMvjzBH+P8U8DhpHO5Bxc/4LfFbdPE56/8DS8USKwU8/XwEIbgxTTBR9jN8
GAfBHrF6a8DEaMvOhvVdmn/qN4wHH/bjaW1coKuzJRkQl4Fzuqsyp0uR5e9ypBttQqfDzIF72gY/
8QyQ/IjpWfF6g1eA0CxbTgVpdk7lZxGxrrZFI3KG2MrH6uE3rfNBP+/YJdXkg//M5/HHeCl/pWaK
Sdr4asCZwQlN9GMLNW8RbMTZi/sxXVGYiQfEwRGgV1quAhwy/kEhKenn3+Ji71274F+IBj/84lpN
iUi3atxKRL3n6QKUPWrMh99gK2zbwKuBF58hmMLtm20NSigDgSP075WjzbryJCtQpPwCgpdYJ8RY
W6n++L0wVucc03ZNHckukk2FW1rKRg/xF5aQCh+4ySZcDUjW4UAOFvYz10L+N/M7jFzPvn8LHOgW
AqQfqV93OyOiA/tF8X3YIW28LxC15vKnxs/Le712Ylc18rrfgpVcYGjjR2MNq+re+fLoNWRdzsdc
2giqS7WskQ92mZwttDyaHbnXZuDR0PX6+4lubqpyAOlHDFyL4ZCBxeHKD3rA9CgedwYcjOjtTblJ
MeQadcpJ8cV7oxciTVuOQvjTBn4rhpHGfdcyFUIWg78QlSw8+E5Vz9LdIQjmrepiNCEgNGS7HgWo
QeZW3ZEzLltdXMm6w/jWEa4QZ+O+yJ8tp0qian4FXOqPrUKQ5n7OzpDNAdbpLMyoEcIPR1V/YTQA
11PatKSK2c8mZBr88KadegXcoynVNTPy4DYvhc85Cnt40Tnw+7h0oUL7FULrC9xKcpbcnc6DEeaj
Iq5EV+Va/xuR4TcgLG4ihRX4QsT8iBD8PqnKJt93GIFbcv7ahWaK103++lEOp/jibOC/qrXXRYog
BWGBysVeDr5DA3n4gVwwxoNDdqhI8JkiG/sHb65MK/qOCOBHNNZ9xcu2ZuKGC1gcMjfDV8yPHA38
EqKlDCelx4UTaKrCxMyvi36ym5mnfnW3H4xEPe4Z60pba540v2na8pq+jCBoCe3cQJFvrnRys6wC
JhPgrkbGl3/M1KTzfZ+5ozpCLGqMi4Dpa7uyMHbNDYWj4DjYAWEB2rQ3QY+xaO+WybpuI3VNqsWS
DzuVioi/vtyez86C6dNicS+XTlgaOByNGSnX5qrRr92STbYayH+u488XP/pncud//dQafYxhcG7B
i4vzpzB9Rqrvyz4rIL/ExIZ/q+G8zDujmHg2PwIcOcZEA+i/gGqooChd9UUe20CUHJZMrjZLkhWs
3EC9maKh/vzyNGvi1QNDTT85f1DiGYpNjl4OaXXJZeThkfjyfvE7XmKHWjnoDlg2d3NOW6+g28BL
6qGug0CWWpH83S+SCdWNep2JF2kiVWGas5QgMeu83LLngwel840fgpV7GUCfybFoVAa5EIjpIW5l
gb1xG4QGfqWI2zK/Tin9IVgs0WkgYuq7mo7d/+b2TR/cyi4hYqJOghNPx6Dn+xw27hz5f8NLKSU2
KC9AkmWyjcgxOno584E7rKWJ2D0AM7l2+2IUEwAa2QSjSN5IU+oMWoIg4wW8RC6NbRC4zfO+WrZE
ayVY+LlvVEaLOcwHV9070fKjGgulRlKtZJ1vlrmcV8nFxb1do2RrCCAPGE03EUniMSH2ZyGfmebp
oazBxOlJcK/1jHhsC7f4ozKE1N3jaov7I8nSbLsONpwD8kJVlD+ZXjy90hnby5Ddc5+OaXm0m2tc
t31o0l4pgsSob1dVL8hQ2CrzQfPp9Sxg3E64woo+Zl58wGQURV3lL/BAJIrERzzBKwLqBUhOc0De
bNpt/xR7EP+obB4sVxg6137e8+K6cMkN1kPEja/98ikZla2zSfMNNaSV3OgCkxXqRbJ64woCCf9A
g/jt1w4GIScSa9hQn7KHzFUNAzwlUfHwXUyWPtzEcYKsZ8Ih+1hv89xyOsL/IRfySNeNDgYZMWyL
BO9bsvOijmW6fT2k2c1o6B7xbbKRT0vU+u12vKFQRHObYv3RBuEgJBrxAt4DUloyCqyheeNZFtX7
6/kJpLXHlZYLk88XmbX9Q+IRFHYKrVeggxETM3g9b4+E4id7uFLKqyuzGlXwxthpQ165ddedJRom
iWcWp+Iy+6YCmuy4qberj46R+WtRiFt9GA6ZrRt/dkhDIY8DxPwZUlndTgG7U4uLsbjlHXhHTqKS
N/PQJdsbrmjPwayDrkhN1vBBi3MgZmpLfJNGPyB1EkJsfhLVsWHqNj+HEQSK6ErGEkG6xNgeJewR
apHBT0k0SLNDaxxNSn9nTE5ApPh2wMqErYqKLY4rj8iV1RitRtz58V2ROEDG56bPHVABlNTBVaRC
OoeRcfiopAkHKgno2N+pKfiGSJm52b2BY/q2uxDWkYMbnUDjjOUki7+cxsMiC6pGSmJoZA5OwNLe
COdrawR6ZijhoxBFulJJfuK5aCuhI0Qn0zS+01Y6U1SQ+cqACbjZhqGn7gyVr6zk1cEBQIAMZF8J
QFGekTukean4tdu0i7nACs5t0Ug/7JlfCp5vfCR0ve0DOexv1DTVQDiFcgsIpFuyieMOE4IL76uB
AEYmFpF69oDUbL2mMDM6xaFreVH+ehyUOyFnYl9ux+555knp3S34OXMS8MhDwksnSbFeyxJ6CuW1
ovCUFHcD0POgtuakBWvZnW+byPl2I3K7lsxztHlCKkw4o7KvKKGyWVI6cv0iNXjc1v42omo3HLIx
wjNiVkhrhcsBeG8Z5ApLlbItqvgbGDhK0MfyPBWknpC4ZaEcYqxcOAJVhMy8L2pODwIi2V1OmNLJ
G+9muEPgU9+zg9+zpp6SYq2qGoQI/LsyNqEMiJzksgBW8y4nvwARvn4RlaiPKGcKfT+DA4o0nMDT
n8oHSRfr31WLuLFBgNqoH9t8zfg/kqKA67OmZ5VJKnOnrPJLq+pXAX3Sah2wzGlDXPGgsSgrrMxi
oHwkUJz5yfR0h61TkTCCKeYjMn0/X9Jp7gjEE/PPDrcMVQ1txBFy6Qas3D0u1BYjG0UI3sHUIFGe
AsE4cbEK7aARNk39iR5ID5+ydNthaPMLgfMM0RnuUbxbwwDyjBGe5A/045iC2EG1n9PR6qPd0bqu
5FC1/3cwHIE7lnml8af/QtLAESq+BQ6Bif5sMWvbuarRXZbVvddPGF+sVIvzlP7R87anT/2wUHI5
ZUpNHAVVCUr4VhhGrKtuJwrZwm3NKxz60lcxe2urrnqRy39ZnftYmGK8PXLRPmXWI+K5yfoK7VXe
drQJFpFY8ghNBlP/dbj+mQwr+WPpYkqXYmrXDOcMzDrGzht7Md/PJFVMwJm7LyjoUsjZZSrBlWVa
Ply9oe6xc+xpaMHTRzK4rKI9ujFE77lmaC2lsugL9ZIYB+hqDYgKpC9b5vEzo/pvJ4fandWU7C2x
6GTmIGjr33+o1CJ3qjHTwNRF0DGI74FU1NzZPr1RZUkIxtEt/1viQAuzggccAGM4jAFJDPZDQbia
PtDuXsGQPq+w/Gc6QrYKMORRR4qIZbmn+b05RpLGX/9q7EPXYSAcvhvDVv7r/vwYAUsy59CyDDV2
n0MnuBJZG7QXmxTMHwTyBzE79/kZdvOq3OitneUYiqdA68nLsiXL9eK+tYz3RmGD4h3iLmMg87Ra
v+0IT84Azt12F07lMuL+6oAqkMuZcXVQz9HocjMYzKCv1UyooI6mWYkxA+inuQux3SWz2aR32NiF
dU41Wd+M1M5s/Ljz4mzm3KkeB6LwYf/meiFJuugMp8o3buTxyMvzcxCbqY00jOsaV6b8Y0yNAert
ZTZN70P/BmLRmc1uMHix+wSQsopJvwSdrvLfJE5t+OTSHTW8AR50l8OgrnOaz6r7oa1zsDk4OZw1
OYdqgfPJSxUIV0LU6vP708xNzRaB97wsVz2Sc+WpxOLlRuDtAJpOfK2ohNLktO3mb5iyQYeYkjgh
eEnhm/SWgUJMz//O1Ee2KuF3dV2CjFo5uonyGjonzC/34M1nkILvATTC6QOVkUYYYhyqE55GcqSR
fzRKnNTYIvLGFBjq2oWbJgIJ154slJNZkadXa2wYaQ9ggIx5Jo8aR4yH9rRHtSggewXNl1aeuzMH
W6jJzSmLkgvNVv4VHYJPg3oHHv1xijoDQSLLy6d4DBXEAqtfdKdHajAH6qONRaPh1t/sBUz8WfEQ
VM0R8Mul2YvPbJJZFQHrU44KHAVzjd33ghYlCne6fURIcQ1a2O51mIT4GJGnLY9ICVls5lbka2O2
8UoExvN6pbOxhZ3qcRAcgWQFNhI2giVSWkaxCrN6pQSRoV0r0ogmhP8/mRI2P87AsyHwvSonio8z
ki7bD3hD7IDk25pVmeID8iJ8TjszVpt8u5NTgRGSemvHnQl80PjsJPsoUnuXcDwzSsZQ5IAE04LZ
nCYoyBKFBj/xCl7pLdvDT7S1bNqyCysIUox7NShlk/MddHr4ClQhYt/hRJ9oJT9kiCXSDjK0jPo+
zdN4RyvomPgLAjoAzWKyLjqbvZbFTjkT1PRaybDe1FoE15zX/wV8j8DovxAjOIJ3hL+9hYjPrMUf
DNSHu/GEaSKt7TnB5OdNL8bo+Ta1roU7vVBkQTLh+gG1PS191DRqEcXDD5OF3CvNvm9nVNJyKc5T
3sW4s07UH7C2wi6+7jtn+PsIRPjC5uNQoZj86elNHHUFoNuV2CAcwA5gM5cP9JtgpXaNahTE6EZD
65VQcVEbygEp1imoqWACyZtrttawYxSVhXzYtCcNh8DoCGPvbaJy3dj4Q+EEIinooetEHB+MGOsz
sI73eDeYW5K+z+AIrMSzPVk8WxGpiR6RQiJ8kJzGXARl187EORceP25/SBI2k2Pu0dNtFn7EB4iW
HGzICIyTU1eHleVEdLfrM0XXp6XPvXw73LNGXwFQVvSJH3ReKnoj8cXcFnDqYBAUWiraK44Vwaxl
UdR3WA1Tm3zM8LKJEvRvJB3g3oveYX5iLDoiY8kBj8u8cTiFUmyFUMIuKfb9UWYa4NMADk8arc0V
DyfwOr2i5hz+p5DZRvc54WF5yotILzdkDBHlTjVvUeC4Dtzk7Bp+YFdEmOcOPgAlVN08o+Q9OGHP
c8O3OmchmYC/NUJ/VT4BtrNvKvsO/MdpndaIzcGh1rrQQIkGuyBQa93PHYwDnzGRz7EDbB2BbrmO
36YpAu+C9LhQtQ4Y4dOqXojwTFvqxCdrQEVS55J+eEWYZMThh8eIL5x/fnFpJ413bM8PiHRCiUkw
wpViuuP1j50rpSnOzCQug1OKVH04ErIPQUl1U/gO7K5v4luxwMm8+zcGA/HH3dY+6x7dyUZRDMwG
1QACQG39jo1sxmu/D4J6iCOnnDR3qXPSe0+VFvdxqpoL75R/1OXP+jeQy3G35i3uPZW5gAGM8Kb+
D3DcMu0KUtp2b3Ds3LLsddMV6eN8pAQgXdoxAdY133KvAUhH1m1d+O9g21OQlUysT8v8KDSc3MYG
iW2ClKgFeFDlZWn8Zn9QFK9YRB5XCHagGUaIMeJzzXEeWhUNIJGkV1/4/tsTryAoW051/7OCBA+Y
6/YI46MUizUgG5IdwYuyIDheD8kX9NDRXmTMnTg6TbT7SyexE8BnIzd3PU9EgBM3WcNt+0SDjHaP
ctC95WvD2PlqD3o/wxm5F5mePOBkYo5iDOAyB0W+/73twBE4FcsZadw7kGfoRjchCZtr+H7MG/5C
YHGZTW97PkCVp7zt5X9Vz9mpCCzAfzniWbhL/tSFT/NapwUcWpfXeA0BgkA+YwEv+HhhBnbr3oky
khSCPCXdfG5FOLdAo4arvm0sChE3VZXzah6ctpljjd16UL5ceAYRJ1vvdo0XImxKyJR1zAMv2c+f
Ys7bCQmeN7agN4QGdDTBFp2ynoFxshZpndNVowEGJJI+oUgRNbwtSpqMSwn+1J/lfXl1I3NlUXh9
VzloPxhyMidA4EeeNy0ei47CQKPVcoJxRiX7YaE11X460rMWbASzPYDA/TxGWvN/cPiCRJls2HI9
rayvs9lOdpi2F3YpHtOuQ61Y1KMamrjKqUcz7dXdvYG9k3NuovySONwN8L2dVCbFainaWdy6xnzr
Lzomts/HTYrjaNAsnKffAucyOg68snFVF7rN7XbvDsdTMljX8X7XHPTKfmoQYxX/kZ0xqamunOfR
pkeNm6/0g+rXRgEmPbLYXOJAa3EGJDApk+guk0NfSPLJ9RxYiKoujhCwzFOVF9O8/GfATv/xHKsy
SarSKx/XudSUOsKibfZdceBMFws72gGWyGDEfLEo1M3QvscbUXjGylnAqCSN4cybIZgK3ahsod/m
XQtlJZs4aHSy2xOWKvLAvYDGmSHK7OUhCSFL5wivr1X5tNeqZwUDP6/pH4uCoDy36ngGrjs77W5s
nOGuBW0LXHl8KBsQbe3oyyviuPJrHkJrkzcpn0jfqWAH5p18JGv8zsrp3Yc5Wsr1nArDpAtr66XR
0Hc4FW61DaWCmfscaA2un2sYOK/LN8XwPMg0lnWh7zXzS5nmV3IjNv1VYpuqp+0Z0qr/VBjl2E2P
gvStlf6XHTRiNlbWqp0CTwm1KX4qYN9zpQAxDb78noqi7wsWUSQv717zZaCX/12cQmP/vJ02tK7R
OCEsdnkVZTC3jJ/2lstatzHJ50nTPlTlyz46v/XQBMGywlLSpiW8Z7XP5ZGdovd9aG2wmBo5ejvy
mkx+6wectQg3BYQcetyLH8DpOdKuXWgUr3VJxrS86jvK8aIED+4sf9eMUHp8SJh7EXRY4tWR0OMH
Cr11qsgezDu8IBJo/YBcjl6/yUunOubDe6nxjl9lwxc1aWqL4HEV0CgwIa0yKzrf2JpNPalZadNS
TQA/MFP0wA9OnZn31S9lQ9TKtrU7DDjYbgVxCkV28pMmfZQsklaVFU5JVxmHSssxmiEhI8u2dhOi
+1ECR1hM/QVWsK/XXLag8t3TQz/xHkUjJ0bOk3PdDXxWD+Q90O0huyGm8CcsPUmqfoO2S8cbhqkL
y8zevn1Wqyh0WhJLbnanG3AFbBn6Tk1iddHzlAqquRRogY9gX4WVLkmwlm4r2UXFSB7SI4YoIbLD
royYdKzqMU4OVolkjrl8TSUIpU9/LLNiaEy/p6ZxIIXRpBjWv+HkdcJqYE5W9+6gMx9ErT/WpxEI
xwx5lC/jVne90/MuD5FkwtKZKvFgXQbyw88+aHqkGVyL0wSu5U1Sy799VX+j7+Enmc/zCJpTulTn
yOrSO+e0sqXUnTJRlYpIDLkOBIO4KiW9hhOZ8bu6SgjqlgWzBpEehWVgBW9YrIWP8Ekj/5vhp3Eq
MqXhz2daZgi+E2mfi5mJFASpEyh9yOZPyDzUcU8Wb+YNs+kgyApT45vPXCWmj9q1/evCA3RMp85R
E3KDl3+sk9zYTwYT9XOxhM9jnCY8dJ86rR8NiRgp9doIKsNmtfxpcbTu9ca1knmHDDR1O4jEu+rF
Xbw4id7qKgoa8i3r4UVFDHNhBk8U0gXxWdGnLXqyP8FPxi3KJ+NPZILqIHoG1ZmMi1mAhNJLZdGo
vL2W+KzOJP29JeEyXzxB3fBa840i35TbwXXmuaKK16HkD4idmshURrs7qNBHm35uk0UU6a8X8lMw
Z0Do/jItc51bOqP5CTM8HLKAgH73CmWWpaRrPxTgIOI0kSDN1yQKDDAWlos1KbhaecBU2KLoPiHN
WLDye0XboSkomFBR7R0kyNafNBQk3vDbSU99R358SOeK16DYzjcSdnB1HJA3jxOGVzqOU3iDoxIP
0FdqAT759jn2o0JWTXydwQUcYcukTdZAIJa5lD3FsdEHnuCO9CgZAZYCx+bELUOJDlNyNlsgvb5h
iD0Lh3hnL8ZZm9/H8nxnOYU5rbFBaELTDg3bPzLojoRO0ot5+0L3bW96QuotrnTiLt0sW8TZxHYO
QvEcZCLGzeb7uNA2nM6ovsBM9Np33tG3+4HT/X2vPVimC9q+X9B0fqGenV4mowTYP30u25lDlcgi
QtzO3cLU89+/iT1DQ0VcEm+S+qX4jbUYxWJcWtoWd9S2ib0Vdb6BQFuFDAbC/adwtngajnbQbs7E
DVMvhVMaXY4r/5oqR4eXG58TkJHrMDT/O7LuD0TYrN/anTl6Y21MqxBq9P0tcAAahqI3YyxJO6Pt
HmUfmiPTGBCcuZFOBGhRFsMXKZKUJI69m1s+gX5AILU+eSdLTm7CbJgrVNR5nTMoVO8eYiDQKjKY
uIaI7tQ16XQBzYTKTuQ9Qr15lGgVTOuGgKFLJTbUS9sDVhr57XSgezjGyn8HKJirFrrUDJLRgktb
kImk5o85tWaN/BQOS77IblPPwf8mH69izX/MD1ueli+1J6nRZg8CoXdoCjYV1K77k8To/TeRl6F5
EMu8Tz9k/qM758W+b5slCuKCRt6+5ZqMjE756jmUqAxdhB4stlSQcJlORzNgeHLPpOtVOSSy6myi
Cvl1WuKazwVaBPqAOGYlIbHf3giq3IMjzuFOLMOBOKDtXyUl63cA0tUKT6YduoaxqtsiYmMeH6cK
QOc5meSqnGZavTIoXuhF4tnyHRizFZmJpRaoxyleDdFlpTN4CFO6EKVJGBjaJ5B8eEk0UkDbB3qH
l0aIWgxS8Ub0SGbE2FPbDSxK5kh6W6Dz+FbUMEqb2WBzNdH61OL9yV2mP6lHt4+HysSGOFpmSZ5m
s4CBARuoZcdceDMH8Sf7oR+G4B/wUTJPzKyC+MhkTMDWjVyaJeynGdIFg9kqMnvqvERvWsnJSAPt
taoSNzYamlJomgH3WNsT08kGvPgbk8Aw2qyKKz9lXcZ7OLe0iHhTNIlIJ1j84TI+hZZjoXDuXvnX
k4lnh2+2ZaBUuOdxn+ja3r2w7ne38Q4fUA1BpBFV+hZxBK8Bp4t4b20fqe4UvUE52cWTXS14uuUx
sTWNkCMxVUjevbXGvN9rpq5QI9/hbEroT4sy/apKyeLw7fmcFAQIgdUeQv4t8+8YkpdvUoIidE6D
TDpcJG++ZUtJO2/llRwK32GdEmfrW0yTOHJ+Wkh6YKwrD1dhXGocCNjceHCnASn9fUXQbys9mq6N
9mIFaeNdX77xdfcrB9DyTK9cPaQ+egxgIfhj9FHb9GY4WflqxjQmyy5ePBUZs0dM+FbLXCk3OaAg
SmxzerMSBLIFLkicezgtNY9I1PIOGWErWODEJxCD9D3/Oerc0KIuc8ohmlbg3xE8sJoBjOTfF44j
inxNO1HhsSJET/PNTeck5adzgbeBF6L0jWcB8xFqjXv7a7hDtM8UzGjlUJC4hOz5Uh0lEZv4sH+Y
f5uaK+lZOqSqV6ALaob3jK9+jgcMBr+/otwAUwvgx43R6OFtAMytNVTeIAPFoB56ydQyGuJr+500
4oxYoefsuBgq6pHZj56Zq07rzKuSBtNzBFL2B7WOCCr6otja6j1gCW6QwsfxonDHUOT4DtyuvdCh
oPH6svC1G6B7KcV6yQjUZAB3fr06eTx/Ed6TmSlCw4qy6S5QMZEXs46UoJXyY171cl2Ofzty7M/6
1rf0QpKMu0OXsqtGAyB6B5sQ4k/fFN5RKgn1gpaLOUbdmvv4D8gXl/newgoecJL1FXv3z0kbnmPU
CLooEYukH7B+b/zJy7XQrZQDc3XzqK4J4inhM0XzGBY43Cvo0YTpi8wrMfK2GZ/yzxde9oUwswQ/
u5BbE7cZb2+e2iFn+s87F7HxBJHIbO8qQkVlAL/OcFVsB7zKWFEsORX0y+iBiu1Gk4CfqdOwpt1Z
2CKFRNpdKyLEpe9+QtEPfljTixYS+c0RcvfbaVSxLp7vRbQcQQEW49SOjKjiLUoXvXQqkz09yqIk
znysHRqze2s/3LBUVGyjO3t+gXSFZ+JEq5eZsOiw2aXOFmwMF6Q/bj/E2AnLe0tRcpjnBJEUuW51
UWKJsWmA75bfh7EVGsCfFa5bfyPdsbInli8lxq6N5fkhn1jkFq6B1XFW3BphoQrG/PRMpOGv3csd
ULAtFTei+ZPEIolMDDSiB3lRiiCxaQkgGzdlANW9+4fL9lyXTy2jZjc6VAdxZ3hw948Xsjsl23hI
IAsC1PJtVRrANeT0H8f+SUIFN+srgHQtr5/vXBWFr9TVor1MqX40MUaSR6Y9E5R/EHsWqLrwxdtJ
+w9URY3pyR8Z+6taAtajI5jD7dJJpt9u9f8kIJRzZ8i+qVaX6b1OV+ib1xK5aYWtod+h+gVKDquL
VAvpcqXHXzBQYzzBET/qO4d/R1xIEvTI7LHNLJZSYNlAVQN/mDVHpgLEsQrdg60AE4PFZaJtVhGN
b6g9NieoLuutG/gzgs274oZx9U5ZK4n9nvgNCjfhQW5IYm6eV/ha/J8FpRL4+CdsGvApLfho9ddj
C0Tp4TJJklcwPtRbRgbc1lNj5CY8xclmrG9o9wRr2jRZRcpu89HaoJIvaA8EfXijPgtnn9Oh+pFw
TjZ3VpY2huONEGY9fV1+cra+Mnz+4sE1ybLhhsSWRJKvQrpIFdCbUZFx11MiFlBNPTq6DG7gSX1i
BSUKaLGyrySOJIigZyMg2BN+IUFQTR2BgmYP6Uxc7+xgWfaJtj42aYee7uh6H+ZZS5YVX60sjKFV
LYMjiCvecHVU8Lf6XIZdsn7DcPalZJWRiuAB+o5nLbaQ+ZO2I0H1QH4s1OLY7HoxzVPKldG3EmcN
d78/3HGVOf5L6mSzZVOXna5Lpy4K5KqjlC6L1Ns4MGCOlunBZv7K5msgHc5JwpkmZ2/oakTboalh
aJarVNRemdQiwrDGh0tubun0cvMVB1/9bGTE7ver5JxR8MQHs9J97tEVdlZOeeNd4B3pt4H5mRG/
fUSDakatNSUebgp1g7dscUGertr7XJyfrGjtobxnvOuqIYeE17ZLpoSRJS30zmIy4D2DmcTQov0w
mpIHrahFOPYIzvguo8iSSSxxczlDNgbE/frN6OzlV//+2GHeNkWhlxN4TZzZsygmeeka0FrIRG/n
CWrV1dNhahce4pZUZsZ4gcmiuJWqDS28icLvMYrW9rdlM55KmW7JLhQdA8YGuj6VTIrFIEzJILQx
+xcpRnP37VGLSGUGGYEGchZisWJdzLxBxT8mj1rtRnZD79Yaz9IPspPZQsy9MbAS34Ro+L6J6uD4
9TUnccJScmLQG+sC+Ja8/2kDqgvtHpRy5zzLt3LBPkA7TMnrMf5CHq5WSGI53afXPRTgnSbnfHxF
tQR3vjv53Em765Xv5cnPZsnp7Me/UJWMA1AdmfkiI74PnGlRzYz2yTeqqc7t8mxEranFiXggppe9
yStW+P36vysBv+TceU8xRlrpORRx08rlnpzcWDQR3UTQNqPG65fHet4TYw43zkaMYZpPovVGBUoX
/9rnoROeim0Szvv0NA9XU9RNex64cKFF50kv2v7cvlfBouglaGsnm5XCKVEiT+VlImYrg/9HyOYN
YikfablXkjgjZV1/uDZpnNTCZyNQBByDAm5/X0nAeJ9DVxLndygvUImAjuriKvi86fk18O1kekz+
zVz8Y8m5FbbXEPOHgH24/cLxOIChW3C0fst4Ew2p3D9hN5fE8fHumVOdZIx6Mp+fk8L9XIA+RCh2
Qgkr5mAlKebECtxYGHdw2D2EOv+R2cm09CB+KIFtAcE/+ozOOtkbJrqQZNxJTOWzZ1QAkq0gL44a
6qYkp5nxxUZrfi87A4JewLUkALCchQ40WERA5mwqVmyBYWG396s8sdnIQiZiYRtgdCVzyi3CZwwN
n2UCD+L6zW9JSjtr1fVNIZbxggILIRpccifgOFOHuR59n1y3sR288Fmme/ZUtLfstJ7PN/4odHZc
wreQaArFVpQMK2lc/NT2HBkvl1qOg8ULAUGLcDXZtf0+LRmEjPlWJB20JOcs6hgohH89jYrb9E/4
ayYiKDOzzkuVAt4o4bqTFFUvOSYsCthMEVfLSCjRwDkX0KenufLcv6hoS/BW/wLOsKx3NRbgzdsC
r0XGnRMkmtRGQgLaTotcctimGulA9rvNVjQMar7z1NQrp1m8WC4gpjl3qetisO1u79lHE/2P8F49
ClmyvBYuDh7wqbHZ9PioMxxtKYEGeYF/jeNheeK4j0Mc3z0NsJx0p6AMKntdpntDJuWjoVWw1KEP
pF527fzaiX3EsyH/IyRi6k0BVx+OHQb4HDOznyJl0+PuEe6I+zxzJMVa1MGDBJk3HSL1P+YShU6i
gHf3yL8v0yizipytXvovAKyeIcjprtvSVmdfHrm64BwDfwMmgI2tlH0J3LI1ukC6sR397yZQZ7t1
Cpvh6k+V3//fdwNCrcKgBYeitO9vAWIxxk2JqhJnzycTYUS+qaQ44aTK46WmI72j2RcqLACXNXuF
aCa2mMoEfsOnuJ8UXhosvj/neeJNQ3F5To9i+7voL54WSvuLfhCO8XA/HXw3hyoTs4XuYD8qSrwM
NwdOCkT6/OPFOp1RgTMWg7UEkengTzAka0sS6HwkEr2nBTPrUEC9xRez50vmXtvTZI3Xg7VArioe
VcEqTBKOocLqdiAGs6JoWIS1gPhKwtFP3UYF0JLr3fNcOdRjfxCCO5VRd2EX/THXOZi1Npz9pINL
iXRPvRZiKF8b+rWmkxh3NsGLqNlytcU4zgN5XGJubyW/qS5BqL6/1ee68y47P22DWdRLZifnVyzC
0VNtAk5rjViB2SA85/xirJpiNvQ+0xOzcPEhqMtSDMjEHuwOvobgF/mACtaMgeVy/c8ao1b4nznN
LtuSh/IiolbHpXtOWH1L7w6N0GNx8YWODHkWj4k0GCvzc3a/zw2tqvJeqIRRYoBHc9KkCragr57w
nTSlp4XLYvf5c14A5XMM/bpy4ks6r4flpyVkNkh8YGcWkJgrMxp45FwduwwziJ/51iz6dbwRgrgo
D5/cL7sDFWEBa91ON77HiA1axwrhlge0lhI6vCD+eQMaUs5uDvIpqPBZcjyejpfnzKKVKiIznXk9
FeMvnFb4NrRsB9elBKG729M382PtgVK1sQEQzS1dnsZ41IrAvcYMSAsAfOtANurkeVgT5i4NHyNy
4vjH4mDyIU17tmGhSoH2QmD7iHyQtMMGWiHtHTH++mPzrNs+rtFT+EbkQatf5ilFTBXNr1+eHVBp
T2gr1hhK86jKjNorIynPHf1FWvKzJxuUI3vPqqfEJ+WJCLgPdRXbGHwIcjEupo2XUEWucwH9ZY7a
8GRUkZ2BIX51uikftTHEhFwm5eq9ReHYEEb3u5udhiso57lv2i51f4PFeWpkXvrrrtcSkTakqXzf
gjFbRxDah/eJah+bGHio2KYNS5KshWkIo/uk9daqsQpaw3zpQyYXjgJU+LZowrWC2B7Jiu8CIL/o
0Py7b1NUtZ45Ys9RYvQX6zn7kL5lVFq1pjrCjAVpnxElR607zMn3+eVchczH3oE29DnuLXkARciC
36TUsAtJ8qMME+3Tie9PtjOP5mXMnxaABhv7dXAIt3SWRngUQ3InpBy8ldzZK9cmWxZ/FKIIoai+
csRk/XOQfgNTBqtX4YxZcmwEKlihXYpALBv56uDxpGOQecuP2R+JtvGFuzLqf1iLh+H7A6aUAXro
ao8u0sm3WSq0cGEhdhQi52DNDo8HzRnvfmeP92yaXjxlHkF99CMGGkDqzhVlEm5oOO49kv05E67w
wJNDf9LdoukACciU17VTSUGJ3YmuPeH43upQtevLzdyInGajpcVye5SwH1KXD7hIA5/KBUA2uQBJ
SJT6vYZPMyZulM0E+SL5qhVVBIBboAg+M+ahJy+BwezVs+KN+92ZfGQbqGhiTt06WtXlwaIGQ8Jp
hwLuzYNTnsbl51zNZ4NhHEPhDOJsehRYCQYwTCd2tLUEa+E7+9DoQMDxvRYv6z8wrGLmqFtuKEgf
WmCQ1BMVWX9jSolHPPeTr75L8bYIEmcWE/U1S72JP/RoAeuyDnb1zPshFgzAzjBvejCkRyXeMxeb
mgAMFGwEYFF4Lu98PVle3dgdoIo58VrE0LdsI16J7/rhXu5DV8QgZCQJnpIhBPWnvEZAgQt8I4rz
qGQmI8CpMrDSXnOCWONp1o3JB08x17aqN5w8K2C4fOjKaffR/cFcGyem91UCXUlEu5q+UoK8dRUN
+LIotEyJjL4UxOSUYhc9Zf9AZGBHsglkFWIncRFRLKnI3W3E6TkKBoGkhzwWY2Hts+wWM1xofrNI
zJgvUx0CpEjZwU53fkMM2ERhMa7ofg2BRX8WqPKs25gQNz7z1J/T5JVJKOGiMrmIzDfzDzgz0SOX
MmUs56gi5TAQ2yS4T72RktgWsAgiu0pWdh4dpZPdzAJtcwj9yWZSrRs24cbx6JDHDl2zqY0VgbG3
S1KnhLpwKNBHRcw3ZRkTxhJ2CtzL58mDPh0vkuZlFXvpt4t4BZEyk/8QCmv2C0In7Jl/aIQ9Tpvu
luiuSCTlYAPdzYVLK9tg5MnXAVuVcqDivPAc03DBYC7YXtn7elchMFtci+wN1iUJadGr2C0VFH0S
EXXYYqIW7xnhH/gPRkNvGmbT3bFcQja2j0qGVP8yiXnnmzL6eTugQucd2UMn/E2C8m6vzukXnXKR
S4Mt5juMCV1zimkIxeKO8kfLmM9jm2qOw1UiHf4I8TgkGh/OHM0AIcWGKGZUOfe1EL347HP0ZXff
NV1ANDYNQ2+/ocADKjfMPFJoYDD4Jh2sASNIxf194C6AHEPKkPwklG2uPSp+vLhFrvbN9EcGvayM
VmY7lZio/10qHwiWCyM48hwqTIqS4cFZx/PfQZAOl2Zaok4uwMSMhS5zoIU5Ao+Fk3thkvRzIuZt
4GfjE5gpdupcqRNUdJxFF00w0zvETgEZ2v/StkdGfaT+WWHmVOmJaw6NrOgWS1tDuMvX2KnJtBCH
t/y6eN0dzZ8mtut7F/2uoUiK/qIwldiGsiOqrfvgBnvdIR1+UXxaE9kzwytTc1rHdJsfAWHND6cY
ZlO1/B/5yshDFhOOgVyoUrNhLWKvwGQcZCfmVD5KnXGtJ+iVWB6lvoHCkiw2Txpm7ZAEtomG2aTl
LbJffMzJrzyJJiiXAO1TmmdSEDDH0Yza9A8BaRyZHE2ubTKOEIY02UEOpxdyQ1gIyfgKQuISJXJu
ruqyk5p5Hs3rRcCFB4hoOMOOmvV4vJGituhOsL/RpOrx/Wlxb6K2+TzIvIwTm+HVjp+T9bAsdbLh
yb/6cqiwDY+Dg0RmJdLYkx9TbHq4cvsBaao72/pGd6340wcByi8LPRKxI5yiqdw2//p9Wh98Bc+n
UgUScwpfweQV2oKoRH0sBWo3qcJFs1CP9HWy1ozC1k9X7Xvxsi7NsevoB+KHNaLvMniO+RKXzwl4
iiuFGFxgQThjkLfxnG1n4SNAmKQtPt/h7V95skc9vMZEPVESxsBsIORff1htl62ltjsMakJz9Hx7
rCxAugQYjRv51KNWQBUvZ1OQsT3/h6B7sWFY+0DYYnHLyHL236fwHhr75E3M74gNedtTQu2oN6ME
eaQIebvYwC2Eyi/nPbCN/k4jrUbxp8DNeghM9yQkWtiYaGat58indLehuSC2wlWL5Nt+Jd2R7K3H
z7tnC0ajyK9W/IrSajdtllH/daFf0est12e8sf3vyhOF0ODI37ZaNd1DvfxTmGdt4KWnKMyQVJRw
IwlPwfn2U47db3Hh+3oXTLiUnuA36vPPMtRA4IjAlA71Fi55e4/dG9VCWU1b8SkhVcWPzOK72VVu
LI50EQjF608trFlfynAta6KiKV6bjwyMtc/l4vWKem9YVwuXUjVd9wyTyzp4FHsYQOTKooi4WxjN
AcRqYfXNuFjjFE+yXT6qqIifygIBLTm6L4YnLtCg9aw+GXahq90RrNPCcUdQxBb+NX1IMpZ48eDL
paHdilU6J9YuXwJo0PY1TliFmLe5ZUbhj0M25O2EYvBdHxG2K15EgMtIg7EtBA5bPM9y0ZzDburF
boGewjcWntiWIJNscY23VjCSFieacZZMx4HfqcMuLJMnMShjaVnBArPlpnpepZCrORXc9Ue8ZsI9
n02OQe32bMG6San2IZdvBIfcDu2LsSAcUk2SWR+cQes6sNSH6zIfhC6LD5cdL5BLuIoB/BWS+UyD
g3sYI6T/KmTvR0C3RE6l6+kQvNqXQE/JPuOxJhS9U74mu7RpzY12ffEkMpHcJu9k39hMMqs1fMfR
9LEs05BsVIJ+I3ytZiOpNVoyE4xM+i5LePvOOlO7sIPcrkQyQ0l47NxDDAzHtasELa1OQ/dX9tuP
q9B8HArqPwOBK749EzzN7pmUELJMqpHYFhjaRaUSabAxhCXOwiT2Qt4SSvvqWuX4+t+c5HHOGv7X
nyySltbAAT8Sz1UX6AVlOFHKEt38XTiGPV1T04jALOFfMCdtFPj/IhJGfHnp+el5EQGqzkd58QId
MFgBjnxhQbGwlM1egjQtes3vwCf63MbdqywUIZhZIQfwQbTSPjY5kvw76idlxFVaJsVL1ttEU2LA
0hsc8nNSpYjXbKyozUrxTx3lAyj7DUX/AwHrsZhwmM0PXwSqNnptAKX0ve+gQM80Jm/zFFgurrQh
YSq1jTHWcmGTiJodE1blQbWmqyFJsF+QJ56SMWl0DPOiKjGKJW7QAB2s2FXpKpJFsvQHyg6UF+R+
WW96KVyy5mWteuD74kAtYNP0rG9ZvRrtGTvNoIZhoPRjTL7JJnOlhQvuurTSECp6FIR9Y4l5JJE8
G3zMu4bNtvYx2l6d44ZTiVzQ4wm9VCLuXMoRO5PQ1qgNMii+wMbR08TtrgW5BPf07ur2BKCKyCxa
PkwzBfiVKzfySfraEo5EV7OCra1GbLI0eQbhSCzEj2PAGUEL5L0BbRLPbFUx3q7uFG6EPLgRPAdz
FeyWwSnpG+YvXMEjKQqSkwU5d71uAjpYAmF1GawMCQCYqEA5iqwQVv8I5exQcNEHjE/aFcByXimx
7NyezrbXy7emCikRcbPgPPeAWxslCiHsk7AfxNkV8RFVYtHmvB6JJDcoO2ObVq5me961NKCcXw48
eh9pV3fi0W4ZBFOclj4T5fVuocWXekZCxPCB/pMxSdnC2IoZYxre963SIZq/H3TQOd/YFp/oEs6Z
antML/n88cAjbJLUaUYfeFvmMgISIM61E9f2t/DkhnnA8jSrKCcmHuCCOel8HXlf0RM3Ccy7sxks
hF59Pg6qbyrtD1hU3nPm+9/NFafQPNXlNd8Gnc2+skgB8wOqAHB9wqz5X7JnWobgj5sYWkB5FFPq
w0Nt+DLd1BMPy4Zmkury6EVUOpFoeiTdxxA0WHkgfVvQnOIg54iHmQkEokDZnJBNaFKkxLZwd794
h1zipOsqS6TniA+VMKBZF0UlYar4PBp47Me4Ur6VSbj4NBuLQ66muFEoVI/bFIcxmCMRCBjjkt9Z
9V+2onVDZorJE3+pz4dgE7Du+xkVuYCbsah7CFn2sCrWzCUTwvDiMBgBjHhaExQ2iLVjhdnwm+N0
503wqe3YL8rc1d6seWecFQKNfpcCPBp4WxCsCk15hNJp4RNOXAF72i5v6hKyxeDebVgoKvn+uu3Q
OwvEe6vv9JmFLzhS9Xt6h3hgfUWOgOymIAI4yscihVfYq0C1HXBSxSQWqTCkKx6ctcoJDeX/fpU8
fDwoMFj20PkjZSizjGUkLe8e7I4lh8FFYwQbXSzGVrzGuKWE4LLPKeZ7keInaE4GBumheZvCrNlJ
GkheySbTA51e988T+asJNAyQexQLNln7RLXYMscFpBE99D+c+kIjyrFb9emOzMJ0yy09ZbuqJDV3
yGGCUOtidO/VUAEicJ09Ml1e87kG3x/kr6dS6GyZ1kWfbvW4n5It4S7sAf25Lqw5R5nGr9rtZ2O5
V3DFiC0wNFMhyby1wUAgwxy1X1/9ZzgN+fYSAc/PtIig6se7Skq0Ki6hUnfuOv+NzURKWVIlkEIJ
MpMycKwahKvoYMfqmyXCFvVKiCMPiUfRVT0f4FEe0WedhGYZKA63uwuvKhx9SrS+/86ckbr1iNEt
eC6aba1s4AJZL0fmp5fCba0n7CFZiKe1JyfuJBdSo/+rB3nAi6+o9XfETj+0iRuA97jSRlQmpyD4
MkGNwxJK0imSiKQFZT4GBIRYvzGyrTuQrzGUAR1hFnctXYe5dFv0N+llG3YH35myKmrBnPHtzh0s
0EvTLDfqDMIcvQegIcUDkrCdjyt71sMYnJD/ieklRo92TukL049o2DC4+aYZkfCJwyl7VTMgdcCj
9n2jSPSAGMgrQgKXu9rEHrM+BV5u8s+VXF5IkXbwcaDfaMAQ01RnV158JkveLdxa3+i+yd5P3c39
zdVbqYfP8U8xrAKIgP4hCTaHqsVxTtuC6gCB6YB4bcVD6FqVzq7nzhwB50rt0AMLUNF7BxfM33LE
Qt5oTKExPLOxrZLqJK1wNecyrAtRmoy0oQ18Ftl5BEFgwxKpmQGq85qJ/mfrFOphwNZUHf39u9Wo
Fb8KNV/0Xjq2kEUxE3YioWTnjb3wum+HXuGtWvwcuOZd7/AAVUALzsOExXDR04+hrMWMTczca8tq
QzEVLplwHflEoO8AOif3goli+umn8T8SC7MHZncR85vgWSDsQh+T+gzwbcC4czRSleZ48cSgA4if
rvRI+T0ImRQRgJ5K8glVvL3bI8quelBUzOaEuKFQIJXPRn+Ydb2ce/71dLFJgaujZy3l2/Oe1y6Q
Q88Vokc3IEzieOczXWd3qYskRZnzTHaiaA8IkASn/uLMA3JSDo3f2hcckbLXmHmUS6CTrcmeVU9l
8yHAOSIHJLgj9JpmOYmKVY1dNiP9we8hM1y0Nfom/1xzyk9YFcTvpMndgvwidDAeBOXtcvd71htN
Mo4gnRDDUAhZ0vhAfzIxQkOn8NBuvWj9uub87oIjd9Y9nNGZcjdG8W8UuFAFyA9MCKVihPLb9E1r
2NNjbyqpacqn1P0/F6NFAd0xo6viYYKCTaZfcWZ8fp3AVoRILfifsG6lBL1nfmyydlrhbkIwBwg1
te4ZQZFTlJzew8X9MPaL0/v8EDwT48hGIeM8cWXvLRFrelswNLg48ClplB3YxNcWguC86Z/JPMtU
EWJC1P7jokvq9iNr9y8B0YxxuKkPDGFhVweVE1Z0hhMDOm/lEpGJHy6TVrjEZ03q+0nT9eRhL6ng
VrpL+K7fK5CSpx9dZ8irm1pt2sPLror+oEDBa3ppbUdM3uwpbXVZYCOHoy/2ROBVYTnWbF4z1JjD
pHxmPAy4mLXJfsKC/A4GJkQrIJRHldILnfI0YQQXHD7RkiyrOYmrT3siSgePPKZQ4vQBlcZ23ORk
HXofogI3aUX2fET8DaWgZfHknAmeQ4Pp8gXSiGnACqfqILaJ5C+HqJyQYWYgRhY4aiLJ30cs6l8A
KA5D2UsKndLu7hcRXZSU3AQHeA9ghasXrFe+IngE2TStnFU7NUZihEQtyuTiv5ZUK6r8gJR/A/oD
abty0eIiYqlbXEctWi0I+gQZBgIsVOdzczNz40PPLQAWAVQkbKXn0EQHi5sy0xbgxiYggRF3/WZP
AjbzL+Qr4FMdu4zevugoxwVR4OYnZACjZRG82MkPkJE5Moi9XZ1XC8gKedcv0eVvX13UY0LJIHW+
apaD1T6tWBC9cZF8UpFQQzHhO+zsH+x5PAMy2tj/BAKUpkLVc8wPv5hvpVImbcMh8vux0UxR89mH
8r/PEaGUnM94+pvcCdLQkED+1WOBkPjJ7FCNh+F5YUKf43TlCzf1bmxiSrC1v6KSvCAi7H1IZHcO
j/3Dn8v30UEhVRe1v/XBElF8BPPUtYm9nBOZ7+48Mq6ej5Mkcsi9WFbqbW75ULdXHol+PdddJL4J
jj+cz3//y2gZ/yXWUhVj1mKK4rW2ib1E9D9UVefQAhe+8eJRKULwyrmegZBtre21hlp5YJzVTjN7
IZUUNeYItLYemIYg+gy3wFrJzi4lMmm9Tg3q/92SvuAgfhb3BrE8jzbtqLR1iyfviXpU1cUDH9LL
tXxPRhYkvSg5ZViSWcabaoXJzpDZNF/QQwLTHegYutk1uvHLLOunw1A2I0nyafATVlFb9OI/6j8E
A7Dn5dNWiXrGjRuHnswJOlvjXJlCJuh7znd9SXEkWGtEgZRrbOFkpODe6wqrbxLOyUw4WpzsSi+b
mU3mzZz3rtZeTff+yOao9/zXuHhqjH+Zo9L1Ms98u3tTKzY9dlEESfzy+1NHEMVNwhRojK1PsxEY
LCesLm8FQcO+R1O8nZ4ZY2li1zea7xR/teyI/de/4fjZWPrWwWQ+Os9u+9mLj+8b3tRiBEfyesfZ
7I+/mUwWePQ5sBICYlB7UAQAr7xJJycJbgKPEb5T9LqxWLRrrjYcFusYaz2+X2UFjVLZtUNvwmDd
RTlmVwKLf174xU5ZjvMMxUg1nPet++ikf/h73E6wLJS8+n+lLmXvDCl0GXSvVfyx7GFofYklX+5L
O/pL2/fzpqWrSUmNuZcMVyGBDaAqOEGnFBfyuQU+8GTR4VrX//JmZBNldBgY6qlmovqYjcy3Qdax
X/3SxeLsh3jKp4E6kmTL1QIlXwI0wjwLkX4nlFy6sjjNUIaau3o7BzXKf8nRgINVPWz0HbjGyryT
3chLWFfTomPIpm2SziyiRyhOMejkWa2mKDhyBuLTLgxYTBSarLEvAIZpBkCSRWTKtGvmyeZMMeKh
cSySUFdy+CWW7HnjTG7bXOSmRIgoSapipg/9ARsS6cOJany4dDsrWSvsMeuI6gV8zjuMBhYCm510
wpbZqQQKioZODe5oGn8NRnXjyvMl0V73tQ2ssDmkbWItbhLYxnToc9azlvhERZ5pJOP+yMINwxrN
nWbFJmwgshmOw067zdw8pZnd8uRILM8PxdHQGe2Kc0Jeh7NAWLzv23EujSRgWcrozfmhVp8FCAaM
uOSSUXzOGi5AuI9YAFDB2y7a8tp2eUEXV5KNRfstB/GZM90JnwyuiK9hXqyOm2iSaxsXFw5Pe6C9
pA/q1+iGvTXXiDrGA05dBqr5tueO4zwSMHTtNghPgwAwQ7m9n8PyEz50dnZOjTJTq9cCCNtqT1GZ
r1pp0qQDgS9tLH5KpVloEaD5slk9WcYhwk+uQ+v14422WOCgAcBlc+0ooImNXgQZM0w3XrEIZrqq
knOmQtBNmBhENx/KjlKwTwxag31vUe6Ddjdt9Zf8yrScgrSV6t2kl0EFoMvbCnRPCPa2mMQ23d4K
n1S4X4UZ/NoCipLWHeVNH5SXsDgBcIp0VaMxdVDBDInRQEZW/i9i9B1LhYwrKWu2aNWRe1JIp3cs
xMnWg8Xmn6s8nIkbugp0Frb8e9T3DENROQvZhe4g6DHnzai/pZ2+VbnmL8n44uMW6lhOR9VmkBQE
fWg/PY3dlTob0PDo8ICtNiQ7El860uxhQbK3sN5dJuTf8E3xErWrlgiww3QfzHxDKcvyqVl5dgkA
pQGaERibHyTeys5TbdTbHfilMzJyYPoYF4/XS7uWqqDk6zdjLfgQAMP56J6UZCVvkmP0e4uKLnh/
6wyG99S9SfuD0prL89a8hfLox+BmepnRcqiNKCotCFA5guo/4yvGiqFccHYOfYBXQmu+8tGV4mxg
FHaYzaGSvmbNTduafzYf9sK5aujhwSgtJeTyaqdwmPwUUiJPQn262wm2dSHvr/rXSg1XPPuO/pJf
smioHxqgCK5K1/CNBZ1lQE1dAVjye5sdgxKoSQuf76FtMJyPLMTeWs+IXCdxdgV4MCmesxFGO531
6TGsUfoAeqbJsVSdUlTlPaCBqjMA66XLk4N5YcPen+Dp/f0iKgvnI1fZKJM0XxW5z7N8lOX0HBjX
c3s6QAf4NP3sZifxEBUgF2ay62N1+JNEeLZVfiwko9fpUwAb4Bsbbc+UnXqs3bx7h42rKzmj0aKX
QfwNdGZC/8w6hUBdlF4VT3clxdKmp+E1C2RN5PCPHr6HOvXEv/4Umn6t0qWFWu1/vc8YhAv3s4aB
2NxNRN6M2X7MjZOqqUXZqktjEgruORZ5lThBYVWpzb2p5dQB4Bec791Cm+FV45VDA/AQeHCaNoAG
H5IwySJG3ER9hx1StRks/B3+335Yaht9pyFH1C4kITh6CyrRCiduxb4Z0fVeEKEXWTo+zSs0WmyB
hv/zYq1mCLqn8A98Y0PEoZ9v9o4j4GU6i88Pyczn605pNpYDVj+aHPwwU7vYUE4PIBdi3uGPJCvK
Cclh8NAEH9JS4x8BfEUsiCeiF+Zv/GUcS4RgnTaAR86/tXE19j13x2BFPjONamqY2N+emR/VE2XM
m33ajmzPbm7srcepCYRCC4BcxLhBmrwkmVww+9vw5UUME5S1lvH6/tni49LPDG2rVbSvDuVgoYyQ
mmf765ANt9z9z+aer1Tbpv+33Bm3HvpRwnnpqRbypfyrXM9+hUFlGEjaqsa3a3c7FRMRbWIk6Ztk
k/vQ1Au/3zrohPTyrHVr/Uy3M1OT5HtEKPm71cON4sJpGIKaLEi9u1KkPtrKvysjsrJey/gy4zN2
b/dZDgC9gsr5Cq7lCnNmS9z13p7JGEM5+Pb82//scEgFYCyUAScru7+2XuJtv4mJflyR3tbaFlCA
8SgtqVd7vBIL7CbxKVLUrHNEKVGRHM9CkgMkL6KX8c8W9q39Ma2o6f1Rn77vH6lpZ/sS6fL84YtQ
qqRu9DhQcZ1mKz1faWPV+d5W/+nNCEZpj/emZF/isAwl5ZKKQ7X7JddNr+9kDx/hCTAbs16HtY2F
Kym8j9FpBCa3XKdcKTT4I/Hj844HMC6eAd3o/J46XU5uWIbz0ckdApIdFIBC86T+o1UnXP1F1loS
S7u1a6393deBt8ibRVTZVaCaleQH5Km6nx29JFHpEcSYXqmth03g7j7NcEKe3ba+l7Y2jH9jWMxW
bh23h3iD4+zPyPPUBaUjAS3yV0CIcCCTrRyEQJCe2KdKR6NLRZeBrB23lUjfIKE29475JOFIA/Bk
ghYeevSQjuTO10jjn+XECpjA0P3rr/Xd+q3yFpGAYBUcg19WFEH3lFN0pqCVUVJtHt/qlG9ZMOsM
dKXN5WxJVlgI74rbPUgA1HJ9ypqU3Y8CyLbIe04/zSWqEcXeyK5dKNSS2G+zt0wRNY/HLrCpDqFO
2ofPuxTAmj/FDRa0tfhQMsRgy5CUzwyqpepl+Yy7EUn710M43l0pmlYc0n1cLrDeMslk2YdMk7IO
1Byq0ywDDWcm3/HUYOaJBX4qNS5d0c57uUw34J+qNbSASjK1NKmtulpHifGo+Z2msWeagg+vqHED
YI37Fg4k9aYyzdRlEJVzr1j20uMKzxCImQn19r1jJ9nZt4T1y/onGZT+U6PW33UiWkeKwX9nTCX4
t+XeBLmMLpROb9xaKo28iCG35+3OdXoCep+a8+eIfigvSZrRMSOVMqr7HfJrok7YDUdnmf74qt8f
lOfWokJfvQM9WiX2ToQv/3gE77EBd4QXDkOG3SZuniBS3LA9CeuUVHmbWuSQchM/rBUw/gqFfXT6
t6mlCiIKtt0jOiaY7pMyJNMuwcYt30gafkCO8h9l3iYSHooxRyiKSMzmi34NJlfGeMEaCkC2F73B
IEO5vX0oYQJEH4HzBUBclQAmVivs7g5dJs5U0b9EpQEmjbqATBXsR/3JffGDmOBj9ELlSPCpVhQQ
UqLEC7ZVqAqo4GaEKvY7ewBTvlerJd4igYEq+DakxVo20s5pce4OUbrBt8jny6dAK5jloCbMoZcP
t6hjDNZr437KCuLpDbNlp8jIGcLbjXq1WuAHqEbN6DLDW+GcVRqR1HWrZvekmehYGHtIDRbp6ozD
Hnx47oUTzIKo0h+xNty9pnKL43Gm/Ao8e9V2riz+ManAvRuljaAWjJsAZKISzbD/jkvcsuAYdQUa
bi/S9lbDnSqut3rreMnvLoOfoZpxZf4nMnEK+9OUKrp3yBM0Q+PeKMS9EsTwaKqw6jf6ef6CHn9a
V0wx5wdJev+DD+i/wVjeNdNMiC45m+7SOENeOO/N2qGCEzGcqiysUegkRqxefTP0AjnhKUNaf+vu
upnU3+C3+F4mR/Pl/cjJZJ7/IkbRM5w3fEV5z+KtoBNujnBVm8h4AeuNlj2yc0CIrP5w97XQkDD8
alLLKRytwo0YIh/LWKCwxlPvdHqpnl6agyAjWskEDws7a4G7jCI0xttNa6WYCYxbRau4vvZUxefR
AU7Iva5q5wgEbKVRNpxqT+fnoGAtt2fAxSEVix8gxc7Xe9RD3Kvkyy0aZFZoEwoagncq8gsDK1Dg
p3kguGthjZNPgBoQyrRITekD5a4TPRpoyxEFcGgoiWLpkQAV63S6H8IRs3Rx0nY+hSYNHdRjbwPu
MGH5gpGHxtFStkZhztQq50rEyq3UVI3iTJuXY7iShIk2s6YdV9pBT4Ir6DVY4hMuS4zrzMpz9gAG
LQna/q8h3N4x7wrCdkOBxg4j+brHz/cINdGzSuPteN4mek6JOGrC1RnHzRAN+AHpvHw4XGR+dVvh
1Dow1Zp5BcMhGMI47ShXVp1gpBskcbiSA+G0R+o5XHP2H+gRkO6DXASCUnvofyWUaz4Gtuo7Gr9w
fz8aMefytMkWLiss9XDcu42zu7hNPGAUTxgwdY6/ixlFtli/qzKD+F5IV6Ylz6DA1ZOzIiild88a
qJE0NnfeaL1x5p4Ncs1/DHGwth/n9sE7pLUabSEUESd6oO5f3sJser62s+nRzw3vWry20zZVWLqq
7CSJVWzeOZPJuEe1/5QH0ZbBVYJK+4My+nHgMHQHi78Cc4Mqz4KEA9GHV1pHR7Yz//pmaDOR0QAN
2qrRZ6axjEivQain97hnFoiuix9Wnuz8NgFudUHthWSgozBEFBc2fm6BsNO0/OcKsQ/tFc7YA6IW
J0s2mAt1gajXAcxSv6+Rl9SKhn1EGOXcxlKEKGSoH/JcbKGo+LcHncyDskCBqtknScievoWGgR+5
GGhPNJkV9UPUk+PEA/Py5R5BaGkF/T70iUCvrfXAsxVtkh4W7JT9mYhlB+OG/AM4QaDruEXF/lW1
K98VUQiuyuEP7bvmmUXemuPMmDxnXrvSd/DAIAG5g/U+j3dN/42by5/QC44wozIdfIW4xVZD8Zch
oKCcZa7Krihk6zZW+imqOuntn4VTv9jlLOUMxZS/f97ekPmCFHDbcl2mNaD4/IeSPLYVoXPX46Px
rpk4M9Kg5HsNLXOlkknlNkLKKand2azQMRO2NerA8WM5eQwBe3tFqYn2KR4t9sORmhtnEiGbO/mp
pPa98smNCFJN6QsR/I2PzEWPRHCrp0PhJ3bAlZoZYH40p452SWF2pOadUH4FTSic3fxS3+bo7JmS
svr99dPg/COcv/xnw7GHZnLgeDM0IdGyiZh4J3Y82L6fxwsmPdKSOFWG4+xouGsqOHz8RdLAnzHU
kEFGCwh12iPRMYztcJlyln5XwOM5E3sL7L9LLaqhurNrML3wyBXHl1N4hjGhIxZ98iD8bNHFiL5E
sQp6Xd/rKmX9CYLmBKPoQ+/h+eyV0n+MHKk0S2t3ar1IlYHFf1Ewm8YJEH/wl+vEGY+OxAvsV//e
qSbYysANEVMwnFOtGjka4LBoNqL+jlDrEyanyjgmxJYIt3sb07kxEqwqBlBSQVjLhYUuqfeC9YnR
n67TXdP2GHskgK82NOMpVg6sfxd+0p1KfAf+ukrrm3cf1yaZNwEO+jMZ1ee3CY1o6h9CPz+5ttWx
T4Jc2LqxX5AEPovNbYphhMbQLMdrgu4kHOMIvbvwq0rzsNWOnsEo1DQwAp/Fvt19LHJ2I6U97kUi
LDYPbAxqD2CxEPHUasGsnOn9Ypqix1Yw/p00exT8eq8WgmHDZVNwKumb9k5A8fSnbD04l/FwJzmA
+ExkgxN/4J1P2Aa0YP/6gS15YyZqQQ95tle1bAAKK1vfTvRckCo2YC5bwKJ82Wj26lfE6z3bHdJK
Zvb9DGi9SE+b24dCQejKsQZKgvjbgl9aD0zPBmo6lNoUTzVkGBCzT3CU2Cw34+xn8Vyq2qy6ztYp
ZkFBi5/Gg2AHMRBwDjb+hyVbj/BfIjIwkMocS5/DQit5o4SFDZ3WfF3wR7mXFDSVny6CrAPzsC3p
VtfyisFZd9jVNDg/+WOYQy5n7sZ7HERRjtaembWGkA5uXN7GJ/S4eoLiBs29TVpkjkAOofvAsxgq
Hc5lhCUXLe+Reo1s2RRA3SWBCbskZV2VaH1tSMd5bvMwHBokn3S6OGzIzSDcd6si8ErLx3/Cp+C9
nA2Sp0KxoJwy5zG1cRwdhOqj4u8e+QJBg9Dq7ER8UV33hJAwdJDIRwKx4Q7Db0J6GyDrGEPJgPLJ
pdaHAlEqxVuNUPrzlXfsoNXIVweNZp3/jSEnqtK0yanuc74g4ZRKjv04COfpfw8/YhM521LoJ3gq
rqJDJWAjH+kzz+AS3r/FNOvcZPyWFQM9gfZda/kJQfKOGfRiQru4rBVjK/dBHjOuF5bGvSWxrofQ
TQZdEMZYVJOcbwab1seRgbHpw6bqZXdDhu/V3HRKeWumGIjNo72IKt4VVbbQKNzYxPeWZdrfA/Kr
YcEbK5c/D1JJLkutGqNw+oMcUEKVQyqGHv5xi1kobiFunCTSwUecxzIbxOgrJG32H5jgY9Dr4F45
UX++P3YSsY6dwjFm5I3F0n/Dly2OB2DY5e3e3IOPwW5tb0TWL16/i7APfw5JEVw3qRXzSgti46vW
2NT10cRURHH3HpC/QzPM5kAw5XjD2PDWR8AOTw/vDX9mUXigpP6yuoT45/sxBgbvuiKbTdkfpgpa
n5TM3XG5ltP+Ql4/QT/7+DdDpclzD2smrZIL7YcM4fbJ2moNxz1d2PB6rajDHtNTYRoflAHWGIwA
VQ4yiDGmm93jYI4cjl7b+wAZar438GbZ/PXGMI0N/SDvI5+3I7kOJ94xVsrRLJtRFn81ZH+uj57T
VQXW1U+Qr74WSaspw6rhJ6QbRT0CbhNEc6WqN0thlnAXVvm6uiMDZLTT0vaZACLag8yFyJVZobVB
fMc0F//q5GFYAuwHCQ0nH66V+Q5euwrEfi1ScZaqcjtpQtdaNNCAy2yfDU1tqmYBv9tBlGsDU7Vq
o8Rk7eVhamqpCh8jvuk5Dr0smdew6RBNb5lvknRLtpmrs1HZdXJBNXY1+nvAv/DOLkfXOisEX+t1
A17C5WUhrPj7De4AqdHGRXfRNcbhaOvJUcNT/cQqYl2qfET25o7VxyxY78RYtUgUnXLVmkvmvaND
hb45NOkpdLX2BQdBJZqBZMA1alA1dJ3ibm1ZrhPaXXrXZ7M/9Do1LK0yGBi/1m0LwLQtEcxETKrI
tRq1LSjeC927VLxjuonlMb2Kjy90oUNX5Jo70WyphOq3dCps7hW9nXd3djy6itvDAElOJEy+ZcOA
MpJ6m4ioRVUfGZ7nknCGPrxV9+TPOFDSWM8i4ZwshPpht+ofQ4049cisLOWRNAGTKRe8S0jvDE4u
91Y1cKUUEYlfxisykJaTYrJcSFTTb4bX4CXgCQzebu3Gle2E4jZYGnzfd1/xRTtTGZgHIWAt9cvh
tspon5JW+t2E48PIkKBxacBkPURKPYpAyxJNMYP9K6Kpu110AZtlh+w6T+EOfqFdKqSxRjfXTt3O
pLI19LIqW32YKIzbP2i5uOBRiqZKVFAvXHa9Di7i+rSG7vgoLgUUAr1Dea5YJOhDnjvBIRoL8itk
RlU8iCuz0OLMG/HX4NLRAymWOxDsr95GEQy9zGCeoOG9b+WLOfRbciP5u1Rvn8/Pw6Sjn24RcWEW
gDBlZ+2ZoAG5Fct9EO+vFCMwfOPTB4EiK0e+8eF4FG5DaDABvABwGEKXLjYsAKOA03Vw0oho2Hsv
/hixYqWOJJmkKVpbu9ajzkY4NWPadZu9WwiTDgJnnnqiSIdDQrGVJ2tExLULNk/a0Y710XqU7w5l
DhrrXyU4q3QleudhIIZ4MO8n9Ft1NZV6ntVZtEpmugUFkOZh2Q89u7bk5kuaHHoZGYUA0n1flu4s
5W38FweyD0k0UeCTW7prEzKEcXUtplwGEXVtYEFnLVIHDU7foAtqvW/NanQa6Z3+Fq8KEO0LhEap
s62fapWnJNbvdzgU1pYDE7vREugcVTJj4XwZk6Bu8Ik1t6MLQU0yK2vqWDRMvzgnTJDvybM2hDbb
pVlvyLbtdPcazMe+jH1WlgwCYplAnfpYR4OUKuDSbZnLpjUjmGL6fTqUidX08rF1qZibStabB+qX
9bjyw7MvzDYr6GNHbUFMnguewmQfenKtuqnhyM92sGeo7IOwn8frp9dE1HaIfH9Drv6AkO8W+SIN
ibaTQUe/xzcFe5zA9CSJnkBjTj1DGOswK9BgaHoMgUz1rvl7noSefTxwUqy9TU8r2f5c+XFWDPbE
a1HKrzzi6yLjULFQ9NQyPNcStqRCe1RJinNIZb7fGCUtLtPIb3Sh9lFWko6xJU4STZZleP7YLJVW
Rsb1gWBaGbb8zAI9tUw5t3v4xU+RxnJ0DtJCk6tAr1iNuozqfUoFMFz5SPa0Rn0iHuRHsBqR/I8J
NagbmI50D98kh/J06nGOsbfFURQjQ1NJQdx6ias8uhGP7dSurMcUQRenyZbj7giAWc5U/GINMKO1
mhVbnRq9j5o6Zejj/dLxncubppJcSNY0y5cvNjFdzlSWSSFXATZcEk+4zE3HLvKMWSKvwOdd5Wx4
zkpX+nFoDXQ66HPGdDefnIwBp/T0nXgbaICj/TbQxJQTb+eEwdP2rmNBdhmuRKA3d7cYpMTNZDJr
SEG7/pZAfb7fvX+FHm9OD/EeDZEfA1I1Q42tGCeHKdsR9oaOAOqe0U7iro8ScDWNJJvpjSSnKf/G
StwFox79MLQ9yOGMZHq3tmhMt42BkU/xHia/krbtrUce5T2vinK2dSCZDPy3pchFeFKrwba4WqvG
x+Vii48I6TgPEJEkplsDhEZr/+gWUDtPRIiLKT6VV0CHzkT6bSTmhhnrEKCdn5R3G+8k8GOwLdOQ
TJW1wkMabqTmseHbhCFvcNFHJdHfdSlCXSX3sSUxskCN5ktiGsienqUjiYXaMtSRDFPEfuPAFxO/
IojUVJJq57eTsn86DQ2CozyE7NWbSKsejPMbIcpGeSZoYrJNOjdeo9rLkyDE7/Dyt4V3SZEl1UAH
JoSI15ZF/ZRAy0ddmPVFF2cpbH7LdHd8gFyTuaLsSmc1bEO4skTXs/a4MOk41aa4MCVEm0ILTjFJ
RDJsaSbpCRPEPMv/UrV/CunRVPIGjLXmgC7AOI2Kl0oENxyq0JY+pzTRcmbyIKK4X5fs6azTIz0W
ccgg2M1xk67LvC6kbVTkLTgbZIeBywROHxYZUhNCWxA0kE4gZE/H3882d8dQctMTQC+pL8dpFVLW
DXQDyNy7fzyW+wwbm68EDdO0FvYVrIUtTH7wwFs9lr2Ob43WxnAatbbS27zaD78DWMaHppdL4Wjq
F92uP4+oY6FT6HK40D6yt51H9HPT/fA4wsSOYFOM795221Zww85liP1e3uGf5iCEnSQRS6senSd3
f8u9p5Xcwx+CDqfDli5lsjB6d2AjH9vfR/EZGMrslpPFRC9z30XzPNcruSLFIMvmXFRacA9BF4j9
6uLclOBbI9YqWKeaXy2Zro46MGMa9Zb37r0ySjAGsiH42c4/utBYRcwbdLsope2RZbz7hTeSblxi
s/RQzAZnZABK5hmH9mPlswfsjq+mOLBrZlJXvYSrGelPnxkQcE47E6lC1PcWTy72Fh1j1QaBbVnb
Y+bjagpMsI+oVtq1DzeB9s5crB8DTor2Abw8ZRSRR8wC3oYyM6P6nhTmmtTeCgodgb37T2tV0inL
K9O/Q8N5H7rRi8+Jb/ByKcnaF96bBbsLjvfq+1++yr3wHhSxKNoWPaZ3PCA699TM7WWCQMCTAtMu
MEc8O3j3+YDpuzciM0MuUnPEFiToFWS0fpZt7p7H7uowDPSnaOG6WtF8kePCWJAAVUq76q8EvcW8
gF885a/kdNEVvomB6aiqcLRQ/zcwaNmBoyEIK7GQ2MIoYFEy+Fv9QkIb7mQ0C+hccma6LROCzPRz
wCOGdEXRDjZVxwhiZXFrgV0iTt4KKxA+Ia0XwuZin0idcW/DYH9pvGIQBA2AXA3ic4J0IxszUHdd
ya+BSTIIlb+PGa+7knP836JV5DfpJVQmwqvl86MTwOUDdiCFswIAGqNZDDlHZN49qCOH5TDOzC4d
+v1VW6XSK++EpyhLwwBnSU5nkm+GY2D7VMriVAXTi+7RJzjoF5IoLMdeo5M/9QQNfw2BX2NR0tRR
+fuzO+nDUYxwvCNzBqYOy0q8fL2iqoY5zRbPxKHBbvVIoma0ofTFbOZTtKMW1VTMnUo0b8T+nfEt
Y2qdV5Z+RnmD6u/U5WxSbc7NTusAON/ZmLnXZXDMRYj13LBwbV29rkOmrV9NVNb9pcRUejQHg0HV
LE1RNGAEySaxGzHCTBcZO/swr/6hscpm7JVsXGuH60nr3p59xFggdBMTOurB8g4VALMLjWE8Za+r
1+lOzI6QAo5ZWxhJCThDhWySFvvm3yjG29zMIgVhHidoyZD9YLsCxUkFe2r33/nkyiezX9aoKvlv
I/C4syHCnJMAu3czD7XHY1FyWF0n3Dz18ypVmckcIjENNPm04GWV2VsqMtt7+v98FeIOu4bcxC22
cCkBzlQLNBlBzK6NTFfmCizCqg1cX4xmPXgQBG695B6MD3S9BUWVlT7phDGT68zavPE2OJj4j/AD
82qFP+iMU+zUb1xI7ugeRoxJRClA3vdo1Jd3XmqJjBKPwhCI2wWahswhbzYzAduFXCQjDxf3EEdI
TdLi+dpTkbr7/GMFL+PyZA+2Z+uOq5PCBAXgkIeTX0sbsAF5OPJy6eM1V24fH0ig5ydoP1iHv+fA
gEs8DYQqkvWNkYtM+693JrM9pJ1rYKy4yYAmioif4840shYLhxNdoa4k6qp97WOc0+DXIWnfG/Nu
GmofvoCyWzaVELBnOrnogkefKRa1NmAP53VpS7FY1cERtSM7wAJUjSjQi5Qf22jUaOeeFdU3WVH9
sge+Xmy3AAWFc7ORQk4cZYPuAlLjoXqlQbLeqAheJtVpJ6dHXVvJLhiKermR7i8S2IViOOh61x6N
bWOhMtFGUhARpIRrq0RCpiEaN8dOZ3WpvuyVqiwQFyHGijyKi91/78BjyyfMNVJjTkA3Hif0VH8E
RMrabdRxa4WsdcsFNbF7AYaa07avM9yekkYFkfQePw6IJNSX4hrVQbkdF8mGcXaJFL3+yqSwM0fb
6CyCpfAdnJ72L+0pEZ+aZOedHo5Py/7ZaZgCTWQBfv9jjENl02Ekl9HACHBmaSggMMeTCB3xnJjT
dNQSfusgiOpH8Hps4KQd8Ye2Rq8GddQuCM7MlL6bBOvJZwcNp+TUabMfvmEk0E+W3dkq1T+csJpO
Epb/lIA21UDFi0JaqZy2piB+zdxUQK8jcHomm98P3IUlStksvNVdfhroDeDAg7b3WyWdIrZQyxxE
g0zhIoOPESZo8rWKtUi/0D4wan/4RwRBbzlFTORFnB1TZf+jhx/DwlpH7BSuKfiq1wo2C33Ispvy
aJKCw+XWr6zLF3yxnXVpimffsa5s5wUa32+k5uF4mRyaAXeV2pEsJL7VBi1zjGEP+SjS7j/U5IJN
/CXp01YEy1un1lF/RSmOXbItD/B8RL9JSygfoXHoZeOszokmQBkWTHykdz2vg7rBtMw/tzM1g4I7
v8E21f5cO5+qFFMppUStMDQq/cl1grQ7zO1RzXWRPleMtTvVjWgeLcSLdMWdfm54XvdG8zjBPoUC
i7md1y0Nj3FxXwjVs+RP8QKgj4z0JU1zn9FSYKkDV3dzIBrXkcQWWSvSHVW7yprYi0IP06Xv1CkK
W7Rr+SBkB9nUjMiBTzXL5dgIn4widiH65d3Ukgll8dGClvap/IRPw3V72BjaHs049lUA8Bt6dqWg
UivPw4dCE3IzQS1bST0l07wT3e0FDR8Y8FAeipmTF02QGH0JAo9u1AcAbw43+/ysFrndVg5cn759
Ca/x3eqTifA9mMm2CPyeFBrCbp+j1s5o4awCpurMUVmsPubcgc7tRmgAlFJFUTXAxzbPRie4HRd9
/ZTZrPMCVhvFnnGktJduw9dWjvoo5AXdr2HYie5qulzxAnnJ/cmA4I+AnPLowZtoobEu507tOFqd
OxmUNI9NB+IGEHN03XUQapI91hKZFYF5MbUQbOsLaZ1ycc7AZ2hcOmHlIFheozLRiKaZfylhNsrA
bDVvkvsumE8vyJjH63oJLoz5flaT2zXo2LdbOktQI+uycFvTz3Hm4BTe8XhX76W9hdo0uYYIiJ6P
sz7WGhp/MrkULAQp3CSdC9uo4c56HRmlpu1/OyQrGaU8ej03TqHdh7OoHraeBMrS8fx3M+/BsyT/
wM23qvPN2ZCNQXYcOhLjfYzefzXo/Dr+7L8CKfvhl4ZE6l3zmMCwzaE2QS+cNvGdBFK7BlYeLnSR
ZofQvM4NUAtm2xq9DbG/Qsw5xBvspt8W9ZR05BVjHT0tbYC5bRXYuVQPUNibu3OqJwK5fEwMSv9i
7FYZdf2XaXlM+W4NRih3JhWaZqo+UsBhD5lzrCRaW7YvGkDQcZ9xJjuZaHw5avNl3TWsH77Hb8B/
sAHFW/05bol0wp2QdQCf2zUbARpiXHNvHT37Ezen0Ln2vE3nvDAYZv+aebj/Js4pv3cVd4cI5DJr
ugwctVQCpAVMADcdZl0SqSR58Y+ye+5voghoL/WCIM8DDnP4bumoBqa4WgVHH6TM9R64F9VyGxdb
aK9XZo34mJ7TSg7D1J1Wsht+t1+gJESrqVuOr00BIPB2C6Uy8+HD5KMzNjAImOhiTJbE/8ceRHF7
/Q6f2TVSp/7gdaS9QBQ97jUE9mBPIUI887rKipXGDWGN+9xaPskuGyABknpsqtK3b5GB7qCYRDHD
fn0dAVFMhNeCoh4/zfFeNTRusybXWicOdeMcYfrpRcxtAQMDP75KZ8xKLen6NvDP3lcZB5Sa1AIq
3gALSpg0Qe40f3pmTO7q9vsEwEbYTegi1T9ykVO+VjmQ/HReGmgl0F9mtVL1CjzrSOPenBy0uCJE
mq5pxOwRzYBY8yVpWP1YECS5Jgo3Da1CsJdS/upcpj6N69CaCzwXiNng6zzY4LotnuCtLWsWNSep
UAxAomRZwk48XqNfQey1/m0zWTKKYSNVe3KvqbzqfRURuluXkpM4oviigDpKkB98JwsFsn1D0D+z
7tS/kXusGoDUPeJZ2409qMeXU84Elolc6wPCXmHaO0GX37uXP4MzM/A8cs20/FIxwzz7hzsJPYtZ
GgkwRf4b/KAJp4ml43oL5mXIKB8+oCx4u5OSflQofL3tVxfUihRlupyyto80/hdsKdG7pBVh8fir
2jlDYOjL/6HHfSqdCVZ+I3otMcyaYeB/fSm5b301cQnXeAFV3E612rK1Mw9EXjCz3CMmdA7k+ara
jwW9MbplUGecST24wXdSL2Il+6lU4XN7JfaM8jn2A0zNbKUPjxliz1X5K9m4rul5mDrC6Gl0uxDN
7jq+1jdb+PSU2+dJFiq96VSOts7N2sE3IaprcL3irm7lcGWLc/RX0nmTpYlzD1/ha6Ietx5o7Axu
4Zn+MB4HCnjNYb31oueh7zCZAgx+zUDHhCrf6l6AoHBS3OvbtfNfxPF2u7jgizHldYgnIXfWd1AN
wzfwJVtgVTP45gcIXsdJE8yNQhNqBq1t9lokjV+95W0CObDWcs2BkktHfkWd5WlWH07CYyQtgYVg
gAKUefcPg2PiQ0fMor7JTBBJmUjlPI+fA/uU6k4IxCSUL7k57MQN8sYuHzZ/ZaX/0DiRrcJKDAe1
0jV3UGPoXiPhEC5A2ScoR0pc22XuDMvvhZjamVKclqLbzHS2ChFSy5GkvIeFI1bV8jCUxPCE2WNB
gJhiSFHdWRpPCUu5o+j0iwxaZ+D5RSJE7Zqj+qjpk1HnscSa8b3QEq2kzBXlgtxcdEg9ei30WDOu
90a1m9Mx2ZLF+5C/Zx0aOuW9eixuLvQLpniONEqPFzVwx96dCdYopFgZCVFHYF7kdSPw0oySli6B
lRocflgxc9tdhxyQPSEXqkLh+69s8f73ulQreMWJyKiqAOrlUZZ/wTquG9v7ZC/e/HSRYV+y2anJ
vptLry9Xy8lGZMp8fM6pfvMYHCbBntXaubdvVdY5j0W7K/ZcGi3hGRYJODhh5IrEKo7Ystkzoclh
g7m6ZxU0IsvMzs8rFA+63U7fOiu3LWODtiCeNifz0yVG+vkytWqp4d0TMebQzY+SVsQ+p/0cqkth
XNActlmWwkyOAao/qCvwOkIg7x2439TUYh1Gx/5QyZFoh37Z4g80Ja5xDjeIvE8FJtAQqFQIhuCw
67tWMcuQNLpuR6fB7keIaT76Y5jdK6ia+IZL0qwlRtEFtj/IFsLBopDUnNUgpOyW412Ed4+FrWJZ
DVchNQUnjOeuDphcnLJrIDaOAG9kUlMJbJQ+6YiDmDA/mE4uFFBzD3jAbr6pfOIH9hbyjv4o1Qto
9Ti/p/SY1MjLNgcIaV4kDvd6BvBPEOXxTYDp2UQW4Y2Exh5Vr9mVijTnEzFtNj+EkuUOcAFggnyD
sPqtAAOp46mNxrL2Suu8GAeqWReUl2R8SXW7vK68MZSWPBkdI6p3AGOWerCQGP3KwfH+Mj35U0oh
QmRpB/vzCXE+YsbnkpA3TMTDSUSRH/SveFHjiYyZbLpYEWfW0RCt0dmQpyG+2whFQwTpI8wNGmwI
X0oguPpx+b8CvVB0jKEWVqjahAZWAgNmGRAQ4tjsoOZrRAlPdAPCmGZe1KedYtQUZea3YijkE6h7
X8SYMJe5/egQkUbsExYVLgNJ8laRBdvwg7d3O/CSIImyf3W8MA1mv1tOqjL2Rju6uhDmDGyFe/3R
9klBXy/Taus0NMBpwNEtrhfVpmM+IHN3BHmFdGZqltdEb0UQ0tDKDB2lMI0wB7elqPw1xdzK+MXL
Xic1g70MH1rzUd3dX/zUeNXm0XtIZr48/HmojrZ+K4bLOCt6hxPLjyD/ho/YRr0zCu9TrENYJnn3
GOf9O9m+vyFvSL+U5JaYuhc3i10W+tU9uiTtg5vFZSJoM6d6sbtdrKQBhDZ532QbnZhQqhAxuZla
fDEVHweQ0njWz4eUt52ViU/1kA2F+tFaiIM/smDvJmDApkCfgQWk+sFFFbtM4yS6a7puBjKtpj+l
fbB3d6bocJzgO5lKDkkmb1WXkPQcHlA3LgtuQRJTabn/t7phKKc6nzy0MyMGKhZHl1PLA2fe2ndv
Ow/bxPSNaWGcTW6GRaoSPUSliMriV5Sq1Gfn5UWby1tY2ZRxidRJOPM/XpGQ6KCZ1mqr2M/a5g3l
zRbQIhiY2FYPIt2t1f9RFkgxUUWJIierFj4xx1TNZnTVj6OBVkfeUQN4o5sKBXWHIAatOtXySfZO
DCwXRioKpZOpKCY+oMZYYr7cXGVThuZU3jfF2iBJHeDz5G14M8BADwY1ZWsSCIlKwZOKscNTlPLI
CyONxzbVC3PwzVw4FS4DgSn6MDxqBNNz5UtqTnBf7KG+iSnTo5yCghEkOP/UWQkNFmCvt513i6oh
bdZTteyl+c4M02u1CKcqYtH74dKTwnsXry3znDuLZDQw0RlN5XoX0mpcFH8Uliq/u8PeZ7DnBujI
kh2c87GD2ouxoBMfPGBGB5dfptt5/cZacjAniMA7h9SwXYMYtoinHhnurPyYabJ9S33iZ941jzB+
gungBevhsqvVik9We9lT2xVfNMGB5fcqO8eKCdLAl9UozxNWRKIvOZzjEDLCzDjRxUsCx8F55KW9
I3O4IhACTV27hMorOyvS11/9z9BLvvHFrJUVsIR8dWY2cc+seClEBp/FRib+avGqyy1R5jsFmZXL
EQl+dlIpnANFecQCUzYNXdcHv2kr/hivkgxR038NcLtu7n8tQRRX0MpXLYp0YpJfZLl67zM6+jqq
NB6QvNSpVJtmOKkPeMCSkoo5AN6duNR0dWCAeLdb2v9ZkdA92NNQp4iptvaJbJIhLlLd3wWcUlWq
++DczczoxK0sTm0v8welJZtRvnWe+4Pai0lOGS4dlFTe9auFKCklTSqbBuBSFOQUrn589Pc9bogs
/gHT+MIDPrMMjkihZ03NdG+meSWH+3L+rm02dM7CsOkGPYlj5FD4/ZeQTtmlVvnlczcD0JllQQFY
xTG71Wcr7osKvm/7I4daTVcrurSYLUs8WDaz4T8x9xumJ+bkxKAAY0ZLSNTloRgCkEuVs/Tybjx+
KyeuKEofHAFz8IFbK4spf0vWdm51FcGyb4hfVDAfu6JR1JHqrHTAfKzduNhDEUrBYLa953AZyfuR
yUE8rWUqTwjBq+hLHyRENNCh5n4Q+VP/GrjLHMtoR7Mm+DHfVMlJbe4T7c9IaL3A9n+/U4Wwsqre
givxMYXgNYeetAWVq6ZizILIT4aqA2hbvfQTcmRIS/v6osVlvi08gdAGGIe4kO8colZawzlBM1+V
pRZCuA7QvozieRqrRkyFWEp+6TVPbz5Ku418kMpX5Qlhn19/qi9z43rLOU3L3QYi5uqm6sK4FVVy
dOA8jPSQH+fTZ0tLRAplmuKz7c4qGKTX6tCYbqycaWVU7MKSkWIe21LPiBbHxBfEQpg3UjFKmhHt
81M2Sov04NmSA/s+Dul/83xKhcy/yr2wYP5Coj8pbkSinTUp04oxEMet+7nMYoy/Ab8NZ8vX0ouM
5JpShJcBfXz7b06HnyJHmYoNfFFfkO5/OsQ4EWCzcf/dXZY8oIEl5TCkHBZT0uS4WQAYEIWoQEtS
PrtHQqnMG3eK5Cm9sW5JMANaIiN3OqAkCpWcEkxIKbl51mHYbuD2iKricDFddXelTzqRF9eY2apd
VFxN7PANyd0xv7xYY9FnGpxAx/7W/X4/E+iA+JgeHoaz/zJ2UKlvOyv9jW+GOb/BdbNyy75+Iw7J
YqyjatBvRh0cWa4SclZISxwKtoNITlqVHGXhLaKRaBF/oFT/KOP01V2Z1JlU2Bgvtot6LWyY0L2c
bJsl0tfPLisnhVQ2/HbFSwHGw/psAQ0ID6qbzowOzz4P0UnFVqvlKJSdZef+yKaChPjX72BupBd9
pYKX0fayXjLgATXOxdNnO0wHH7MV75KPwlyGPv+FABnT8V5zYGFD2766TZUOLjcjAI2VxVqrkdwr
gJYg2tW5VyVYYIGD8bhmiWtut0Z/g/cRkCiaOTtBC1eB5/32NJLRHe/PUWHX9Id3bsbNiSKYxRln
y3QQeBjiJuF15ShDAxn/+HpwmaFVjjF5hEEd8zx+6EBRz3OiJpw7cB6qFhdrhpX1LEzh+zrPQZs3
jr3sCfCciyZchqolpZyC7FJmSpne6BRbBqDC9lPZuZzc6pVqfOrP6oeD7dc967uF+/Zy7xHGH79M
KX8z0EVqE/SHpnvIwsUNjr4C187BBPeqo2fnKGpVs+XeJLX/K6U5q/CO5oQwvhzM9yPSLg6ibqtO
ll2RwJbwn7Jk2J8nhQNdyI7saU83xMH/VM3hMyJfhb1GFy/a0ODFJwYF/zO2Z5LcYuf76n7jLAXa
GNW1k3FsXP8pb2M7+UHiVedC+BJQjCpC+1kjfGO2Q5DV9XsxBuWvcuS7srtlx/ixE1oZOXB91IZU
3ZFRrggnA6MwqcZ8ko1WHj/Y6+8fuJzYXPLIDQjyyyI0sW/7mEW8PVTDt+4tswe5aBerU9PRWGpA
4HYRdmlFdKxtXSSRp13liFxUdoo+HKzeDm3rgEV+TZBeKHLKFV1YhHSlHa/Wdoqheb+aZWKfd+fe
A+K3jZGcgmgbpVHZKnayA9FxsmhrOhPrbTEXP5ZCPjQ5kOjzbpZcj6BdIJpihYEdPSAA80SgU/1J
4XMv5fEGBOl2hNo28KzrE5zJ09oNl2E22482Y0+36j2JcOMrTAdQraSpbbxbcdSfY3Urwi+vXj0p
KCsml4HAEU/bN4d+exUq6GDexZ8b16MqfyP6itmYMD6oppCA8mBlHuScNvKw/qy+kM+bZZs0x7u1
j4F9Cy98KCl4/u0KmDl4qqwsOgVlE042SHefIaSdAVJYWDuc5KUfr/keH0p+x/L+67zUVSgx3sWV
74rYBVWhZMdjorGFfk99JoHZBe9rZ9Xz5RBnc8/MQT30fSFUjbLgyT20fvZQAeeYV4FzvWCWHQup
AqJwQYL5ZGIllMx5krGbxkAY5F58/BD4jQseWMTwzEmfhkIgrtHQdxVF4LJzUDCwcV17Z9Cv0fc6
noaqrsOSEXyq29/6J3siRw33ocswK8P5Fx4pxKw5nyWnQFsl4WxKtdiEkp3qy8tp6qexULRXRoNo
NumrtygEgWVSPOdWc9/tmhXbiGT8COjH1xejFmhMMsVMOi1CGcTr7z2fMMn16wgMY7VB0UUGggRw
BcxFke0mP6FV5Nnn88a8YWJi+yk4lc1irtBMfys2KaJzNiVEr5ZioBB5j5zuPbDIq1+ITnWtnKX6
LezG/Q32z5bhkhyJH3l6BFhSqaN+J0H7bA4Ou4Uz0p61PDrzNFvLBg6N2Vd0OD/npWgfw7d4S3Je
STlMNoqBSuAcV5nsehjKbep8GMBTSGZmxy37Hf1hfaSXRX8S3dU7sQ4nfqzfqyrtdDA5+dSL4F4w
hNusK7wBEmR2SAac6fVlZfnGMCBm37968lGX7QvhSFP0e9U8C/s7NuCYYLVn9TPnvDscxQngfCpj
NjXv9umOgjsRjciBVEC/pS5Gd+sNRAbmy9nc8ga/PbLnJzcd2GSAJECCa1Nh6ccKRFWvG2QLoDWJ
gfcGv+7fluxrpOqUMgKRP7IAZ6I/AXgBJ3kC2nVjuq3wjiWQZI06ps6CAK7tBcWOxHhhiENdp7dR
aVUbv8v+AsLZ0Pd/Pv848/fSEnJE3fzg7YgZb4YHvGBZtxY8KoT/Z/+grP7xcdatKOzPciuhhoIB
fFAoumc5ZhZIPy69MjcGWfX9Q/RQ+WIfIMjMPhQc5aPfWYgioamO/+H0lEZTxZzs9p0ouln+qunT
og9KmASU3ZVPPhbb6L09vCzbCUn3ZuKtXyaXV8csYirvLKFtbV2sC7SM6dp84//O93EDht6E+7vr
UX4Wl/fRw8sMId21Vi02Oov4d4quVDaeifBwgZbW/yiducXr1gkIQiRMsE1202AOa0mTtyPQ6dYB
2pPCgJwyV5ggUeHiptkjTRchgUxppvsfcfrv6VLNIq5QkfJgK7PlURFLmkPb79Em+/Gs7zYcMAVz
eyzy98giRRYf4BalvUyUhMbWcsm98NwDKbTAzq40E14XkhJoDh3TSruyBYIVScnTS2PqO5W3XAQQ
CNvO+HhQTYTynpU7lS9/tIMowbNf1NtR5xAHmz8iNTgS8V5bLhn8le+U2bQe2N98MiS7e6BIPl/Y
dT+oOCJmj9+d2ypCG1R/a7Zt39LeQHbV1tofScTOdJVu817ucqI7Pa3Xo4l8wPWneDmlJphwxW6Y
KMK51wsWleaTp73WL1DLQPVgFB51W4+5xQutJjTMOq6b8Fz0A7Tt9NuiUjibNR2/CkbkIQar/wUB
FRNURfhKhx+8lpYitfKXMM6vhxXKEdXmi6QAUAEyDo1yEWKX2FgK77+iv3STQT0a+Rb0nsAYlm4x
qR6MwKriNg3/uoW50t5vytv1LHWaagZtT56bJeJUyuf2XdKYvWIHzuMLSUMuk0wEK48dKDsFIQzc
GQapOBeQSW/eoUnvzac7iExjhDMSalaMCNusQKQmzENssWIaH7loxdxkvMZAOyxG5Bt7I+jP2kcO
342m6PIOLfub3YK60PQGzdhmpQJOn07LKz2o/krCpd4LluKl9VAgfD9rudcfzlm3coCkhqUC5oVU
P5L5OCsJ7PdfDnhZDT+0Ik8RsAW/tiJ4txZNNB9LDqoPjrtxKZs8ZrEzfewV16TeGWzMi+0fIp5m
mkbcEqjb9DCPjhBhl+tfVhYIPUwXL5W5jtE/gKMG5tpak0YwJoxSI2W8q2ELr7n44pNHSW/n+YVS
wKIFXk3aMLiqxqR2qDLkJW7NwHQCBiQtRexutCKsAtWBgD0qS4rCDVZtaD8FoKduiq4yLZ4wR9fH
yjxNU0m5A7L5ZrIeT/Oklag2udEso/xBeWAI/hzNvTx7pdrcH1WNf7p80dj/zPtpig4uNQ0RBtwY
eGl8KRvXoBRv5wGbInc3pJ68YGLSiEfrRhwnvL9qJoTC1OE+rJHK7qMKDqoxptmC6ujMzx7aYEqN
mLs50PegI7RmFNKbciCLmooyVBLHIt4QitfimRdcP9P4Wm6HA+Jtn+VeSY5Xd4EGR1H4If5XJca0
t1DfEW9WVEyy02eqW8/fj/pHsb1mbD3UJ0FJbdoDCKuyhBCnr1Ntn2Yqq8GmjfAzkN8xbpcsD5jP
5ZnxvDwrnXT+Lk+B13PLT5+qs/Gsq/Iqcc3r8R82tHzwbWE+PQpstBC+NMYl1jLxLzeIl3yD63As
B1uoRB1IibGox1wig3Fa2YeiF7r5wgtccMTuF0a9DzIZcdIGzGLBMO3f/n5cIRTDywHVglcpQKlu
aiyjOVAKmgEcy6e4t3HQzX0gGPkdeeXSbLSFuLUapP5z5y5Wg6QOHa9bjRggedNT4osFR1JYXHxT
dm6vLQ7YWnhGMgizb6mTKOs0cHOUZpvBNCnWMx4SK3yp5UJ065e0mnoki0pncpca8qg+bf73bdXT
Z/DOuZCu5hlY7FkfpZqOBnrb8ynol9rtYP58jYgTwMUOajArZLVmhhvF2FDizvPQO9W8Du9z7x2/
mGN30GPXhmWhUWVxHpQCg8QWpPSqARbKH/T2hhl7rWzLX/N0P5qxZbw84DH0uQ0yPV1BsDJMn6Mq
9fRrHJA+gwoyynNPRYu6Ss7/cfznmw46wFHoVyEmcjoTQJx8oTHzWmocJt0KbU9hH4kVIovJ/4bE
x6gh2pXrgmvOhAMC+hV5UdDYxVV0mUpL1Zo6M+drVZQYbnMWrUZ3E0CrimOjbJtOX3tCQAcWsiaj
DM3SfWG2pvzz3AeN7iheNlP7ILiCqwjW9JxFBdY7J7Fj6rNR4AKLWfh8DljDF6ISLNeAvc2DI2qG
8CdNpPuVeO3lXQ+Vvouo3e7h29xO9kbyi1BwMTga3yxWXOiPuuK0dNqlAfSL80tRPJDDW6zlX2k/
kg+7lEoJ8PvSq+9MlvDv4cvS4D2Te3neaHc+4zxjW05/y/EzmpIr9hM6F4+J3fQ+eaZMR7sAMDpU
2bN35v+EEFtElpZ8ZeZBq7dZ/XqqHtKfGiV7+F2mOW8AbqBPbebaxyA/AfDF2jC5IIeaUS+0Lflw
Z/GXYuW6xmzu3BdFLbWW9mjCRmnsB8vx/SXox2t2q2dIKousBPn7LqUMRN8EudYPUWaAXnmA0DGu
XjQjtepbr3TLbt/dVNXVOlUmRJN+I54Bi2kAvtMEiUKr9Kb69Iz0slw7DXDCZ1BsD5q2izzEP5qs
4G9LE1VmrwGHjH+MZ0Gg8WC+VmkMVTuaT9RiJHShK0TMfv3FrDu7h5Wzyb2hTXXliRg+UaTHIfAh
POmdAsyx7H1vLwJwErSxlMbMKk81ljYBeM43oSLdOyo3KFFCiAQ/eQh0MBWlhzJThCTxbTQu9irC
Es4AMnA+8sf0rGQd5tXfl9wjWu3k9M+rTKrk1UTb/AwzM8+VCPqW8JVA9Qa/FrGarka5LG2AkTU2
4IXAdOBTrsTU4m+6qptDjnKQDecnjCcDqPCLMuWru7BJ4rbq3wUypzwIPp5e8SWcFzsFmi5Q7whI
SssPmZ2OTJw7A1ylWw8XJObVuUQI7H7zc5wUxKj29lSf6ypHcjXHkqk+bf0Oel+VB+XBg50xuboU
U7l8jM5EKmo6P6BRuJHZfNpnKx3iEXSjV88HyVWkA+IWbWjPNO4LzUTmugT9TGd3idU9MSDyE7y8
RYUUjYmAcitVm3Gqcvq5w2+2xvspN6IgxjUlIjikW3e8onJRXq6o3xHXIpLpC9hjc2Uz5C4GZgEp
P8fWp5hcXYStRpuMCByn30RkgShF7T0fepmNJVs8oEDwIc0IaU/p3Cw8wB5yRx+c/ZVf/Er/t7J9
Bgr9XWlI3S2/pvIgB6n5RqBA5INn8LZuy5a2r15cIO2QnM/1WHS45FZRbe3+eGlmoRoFp/ec/TVU
SWK1G9FY2u1zC1P7pWWix4oW3LMBAjYVj+GCwWaNgWhQNSS0+9bfrSPDp3zTHq5UVWF9IbZ+tZxf
iCvkKHaYKGJH2a/X0LFq0bxRirSCWrZRiAPu5WUfs5zN9yGZLg25zSdggfQquOXjy+6UbWSnXHJM
vaUNIR5JD5ygQV6OU2wtlGXWG3SPMM8zN0toe1tmLice/2scfjP5LW+juiYpj9b/yoXg0lQ9jNq8
V1EtxDj4R0Q8ha3ANP9ZW5y9oQsKySArUjQfji62yE3sfLOhWMmGjeSwhhCopzWCZEvISGsZVQdb
cCUzGjK2Gajj2SpU4vUEpWk3UilvgFUYXDloOxNu8C6nuW5cmEhlF93i6xwC4/tVwznjAu3/Ife/
WPeuQXskz3ruOZN5XiHzWaQq1q72lm+9m5DS0qNI+MFfjEaH0GDy5yJrU5oPWLzigPSqGhDW1yW5
a7Mb6DUedfLDxcpcyv/04tDicyH3HYaPiei1bF2p7SKLFu67kmKreySWJty+y6Bxv3f9Ng5ItQwu
XVUqWri1QofpmFOgS9cX2pV488Q+UnafrIkM4aKBSAWaF5ECAdvwtgkDVoC43iPzbXN3UmGTm14I
aCouOep1GLuyg+39+nqDD6L+ntggEpABtmTlJ5W5vx26UrxBab6Rnlbi4z17+CfEaWVZT/jMjtxQ
OxECs5iN998hF1JL+sxYJoe4iYrN4Zq9NZLC1FhKvOvQsv/oz3dMiX2zXgyhyEdtyr4uFrSsi8b4
xtCxN41iAYfbq97jOcnoz281qJaP7wD6aBStyhIBOk0jJUGAF6Vx1dYBe4G+z2h4BgRe4qGDq5sj
I2jUHxZ/dDd3x6/BxqoUv+4dbsKpinWj0tX7n+apDJFYKlT059X+5K3t8fTg8OA0yVyKyC+GSbE7
9MhSYCFJdIVP2U5ZlQBt2Rbibu8HQZP4gLNs4crF2VjsO4KJacWwHdwewBsx8nW1SUlPYxkx0qdf
atr0P2854/WKyPtthHGctLowwYZZAjAoG7F6Qv0MBXgbgt1tW75aXhfaXVNxMzcPAQxqvPJfNhsv
A5739O0iZqQ7sBX+i83QdYt+d1CvDhJHudnu94yOxduuP3FPPg7CH2FC1PXKEKtuGs0uZyeUUVmx
buKj+5b051irGpmMJVeL+B8JVBAfxacZWEWWzETbm7FzE7EWxoCdiddKXCHG7x+JHo9cjGZibn/r
jUqmSFWr+wfqOa+rVzSQAgoi+IYmr017t5KHm4bu/6DzFH4RVg8l5eeGLsvicKB3U+PI0jF0gBBT
Q7DOByDeSZHdxgDjN6KCJu9zkO7mwHHeuTSVdRk9DY+GvYaAi7HGrIhGDj1rsJZUuolZ7pqTJNy9
PtR9eDYufA49rQDUdgMl998VYiyFN4VF4I+V5o04q/ENLolzRjakV+2jS7FclTVgkPmUMhJofgce
DMzR96/UTI4YV80NNmGvaL10C0+t5SJvV4AAFqPN2gRvsPdy0ixEDBUqIfjs9QBWSKNGWNiqMdeo
jhR0+hP75tNAOwvNgPbhahgBBE5j0uDKVFvitoAyKlDYXpHPsZNFm668iQttsPjb9EF64ktD8fZT
73vtjg6G5P2P1+3QISAC3Gi5XyBMjPyVUxA8hmBjgmgaooHw9GVDJM8fXUrpd6BNoc+VQZps2WLT
WEE6NNLoUoLK46fVddQIMyM9QzZr+YM0Qpi1aEk+K2thMR4nh6HHQleaifIFE4DLnaMfS0RX3lJx
hBzsfwiee0T+Xbi+tvlaEC70qpB0ZExjyMNjmYnX5fCMnr8uzJ/RaDQHOtlT0kGaPOoWfmK8JdAF
7GpFolQwuXuyWSyKOXkd/RwxtGreUpwugOYaI6P1BrFtLMJhwKY3zyEZDvLnnrNMtuA14re4DpsN
4ANIYxuuBdTZ3kjagX6kMmP96xOXvFZSA3pfD0W+MF4ZhmY7dRzzvP+r0yZ9rs3lWBXFvc81ug/c
2nmYwPWscy6J4tJ6Istp9qK/HjWZGTfHA6RhB2gyzSLJz2lsKILrs9UxOX0yx/INoZ7QAe8KX1m/
A4e9Fk9ojg/MBOZP65RuxZapyZx71gMLPwZiKx6rucuNudlM/6QLWGHikOrTGwWAd09NwWykojua
c4LWnvEvNPsFkyYFKkORZIEbR3HheQNaVZ2jQKaJfH6m/yYPSr6oN4S2tLffS6GFNlsLIy/R159P
Hln5ToALh1mJlLok/2FtLLFjjMTzvAIOhSVA41xSVZ1OQEJ02q3gZE/85Hisv3hcBDGimALuYvzN
EiaVpDzs5KLPqE7Kh9R7YJLQX72/nGuw6b8bQVsg1TBusKcnZIyfkKTQahq8D44Zk+etyfbfP0HI
iYjhtfSSDaxq3CRonlcc6CwYKeZxNvnqBNWbrpSDxwd7u3v0LUR48K5GQ5Zeim6f7WsXmi2clcYh
pVhWrhRUkShIxwCC2J7Gt554JQ2U4VLQexXctUgwgWFneg1pNRbSu2d5CdL81nNbDTlYY9H6276l
mg2NKd02qd50NIka2VVrYTXfOl3VhOdysvM3IetN5sJo/xEA1ZYEhMWOZahcGjboUZB7pvy9HsIF
dvCh7yFhg2NXJyxykx8GLXWLEl9hVQifxlaivGAOESvdtI4PIVgZWsr7wItxBgERqrpXveHqhmJG
Iu9tdAg72HdSx4l3tupVCQNeLK5nLDco2dbmT6fMoIuDXJUs6VYAa4EoCl/84mpBjbwh83nVB8MQ
D5ttyZLYAZGG5fsdNBEE9YhLrgpKFuPmkVr86X03boTsGbi0Q8IU/v7mMIFbGp4OgjrvwMxo6GIs
B0uMYKdOsizrkyq85rlG4PmAGcYDun+lTT0OY/YI3Rs9Ow8pXpjqosvS54anjmJr+k/QaaF/2QKV
w9IHlZzHeKodnW4ggmgCfQyHvLxK3RQMzu51U9gtukFvoFjNT5XTJhcfXWaP+qTs6YS7J8iRETHa
+A4bb7OC/CE41ITnOcKM+SFDwEzS4hlt8KTgzdLe+a2uEsRFlgmXuJSP5+18B4faNQEKILDuzYRh
kOKbLguchDuzLt2Pt7o4binqNU9iTZl7IXJL0f68WjdIZNPLyT+x92GQXI2HhXl8S8xZ2pdLbqGE
8H0sL3c2R3WPRu0z8bUEsxsXhmoWJn5bIvhFV+4gHqoI+tD4bJyDpO9t/GOxS1W7a9ceKu5EIkpf
ob2/Nx86+UTnssryj2v4jgzM2VAw1J0rzZoNHfkv+NzH/yF60PSsXeboskUFBrzuiC/MIl6Hq4fu
oK8D+s5mhf4dpNypFk3rJkdpxuR7Y7O0oXe6S7edLrDBTYnDtoBYxxuRShw+DTVTaJsD0CEhZhRk
jgK7EedQD72loxwY7YSksVv/CfJFEnim3peEOeVeokT9ztC1PQzNNNJi57vtcdEGvbWANwT0n6d+
fed6rU3pNOYhpWdpKQZhXIIcQtmj2TxpRZz5BM+1JZWRXa2VtWWJt+E+sIGtnHQrgBji907YrtM2
2zF0zhqeaxLFTpIQpwNW+Fo4Hi2PhukumhJffV8QdH3O1IKViI0ZQpvetz7U91MuOpQtqThspo1u
HOG4Bw158Sq7yQ1YmJp9kagH8lktFXE01cII9oY8HK0yzmqFTBGERWwIbZsent5ppJb0mBEkyjdK
i4QErouugn26RXkBKRh6Ea+V1jm2uoZ4RV47eEM1P+Mo92+gGADV2MEGsAcZJIkDd9sIUTrpOZfU
FjvzAnjP1xnPt37hk8vo2mqRewozV1PKZ2gumD2CG3lFcqhTxfCmd3Mzu4jCer41UzFn3SylLFHM
b2rvi5ji4nD1U63qTdzC35aG/tSaUkU9sqLzODKm53Pq90Cwsq511/UPhuomdxh/ZtyvQQceaBcN
2WFbnhuJDI5F07u/kwkFsdL4DcRf4cqtroKOZnr/G/B/Chq5iAxPrN3vMll5WKb8hIs983tXJu0g
Q6asWvUZSt31XHi/voKu70J5gN4hBwuIstb9zAFrvg+nLkeKc7x+Ue06LbWARyAWZTTOXYmvLLWz
B7z0CSwOYfu9MkijIuYm62naPHG5bpNLRXuUfGNiXazP8vdZlGQ2KG76mrc9MkHYzw0LlC9vns6y
Cw4vMlSluThfVcDpZbly9Nwrm7PBB8ix0TbuDNJerQGB8KyEVYhheRGpXqXV4rboLokMTBRX8ng9
Kjv4EuWBmOeII/M0QaPTD+UYcS6a50n1lEdBE53qt823zRZC8VZxSn/8JFmB8opuin6j0eKvWnzE
SgJMW71C6p5yCVX2nTpYpd9ychaygJFPNDm0BluyNkKY4cN7pEBjykdjIe9v/nOlbnhaBAxG87Do
LHm+0hI+PE78wI1O83C0KhFikU08sTVpbADDyg8hHd/27yCW1zXUjhkcATZ6mpWVYhDQDXu/Fe5D
iAWdqY6hYMiCozZ4fC+Go0ManZNzJqrCLF11eTwLcF4VhZNOwP9JLkR9+ysk3FWco4naRv3Rtedj
t449rhxK5KjWRPiBdcozY41o6ukra4JHfI1fs75rn1m20C/R+dQQNeK7taYntB0LCu64U+pZjkVt
Y9YRRgeWnRwo0t3Rfilex8GbynEi5jpiMQENNlkWeH3+CiaSGjFhV42UFC7MyQ99JUx6yz2Iv4CA
5wypitl56o9wzopdly0bonsNRdWMtzoCcqKq+Te3JhC9EJffXUbxYsm9FJ0bEuGq3gr0aa8zvAJS
1br794iKo3x3NBITzp93dKZhNzgtCWocQehdPp17sRXrYUkDurZ21W63wqxH3RpXrAGykTfmGTFZ
gc7F8xvszrW2vjjAH5MwAPUYHYXRFGbMcdpc3yS0MtzQ0YgxN+e4HZVvSXufVsHogy3otxKd1u8M
I8XVV7VEOzhqpEBMlsNu3iBtCRHHzR4xLyHEBCjM1zBHG3KqpJfOAytFf0dxHIydN232doIBmhbG
RugvXml4kh0xPIeXyzf5kX5PioY/SeJogm1b8l7AoD0qfUfNvCZMZ8Qtm2XvrhqaDy32kWsA2ThL
kko6Ut9I+Qi+pPdSwDdqQPRaSgG3zlkGfMJW57oHTfL3ZaL/IWsNTd98+2O1HYg/wjbW8GkMQAGA
SYIIH4EAbSMf4XiKUkbS7pBN6T7LMcJpWxoqL+FaJ8a/yVs06e3cCWYjMFfw+dF8/EKwdw+ekDMp
6JBejcKJlbuglAEzZMK4qtfjKBuZhruMjJeUHXXYeWglO4kZKa/Tg1f1oFeywnWrGybtznEXqxkR
o/+C6W3O6ZA+J3Er1t/m5m7SbzruFMIK66ZbetiqCngGppsGcsUb/zxBuDEZHRdIy02h/D/t7uXK
6s0JYY6yr5Nlop+DL47kho4NgsWnysY3AB67wsPbqV5u/Ep2SbWDebCumomHNRx6EKuNgKiSv/Xp
3wwhM+nXzfi0RXXzdbq7I15uOyv4y3n2PNutlmSEtgo+ibix7ZwRaFA15iUS6VE9H1BfTEtxiHY1
wmx8oeeGNzlm/YT1m3+kaSndkyRLINnOv09Ghx5Q32SVpCnJbVZ5QQp3/MtqMFlSOZ2+ghRU6ukU
cBUaL+/k0iHbntsjC9uBOEo5JEDtsA8dFamx/Z8juPp9skxoOj3vZXz1uZQEAGdmwDD38F5py4Z6
qxu2pJRbzktkzbpbRl636k/8soQLr9aI/RIx2XeLLweczqYH289v7wkWvIyRIWz3KI8BXVd2ce2M
lCxf4ydVH4cGNaRW0+Awyy18FLYCoGPDen4ZcTtx6cKUnwD4ek3sY22SUPiOo7J9U1vBoo/7mZ9f
tPAoa3RUg3QsEiPZyMuZw/rl5RcdgLzVfr6WLxvb66jYyrMvt4JyZgtYQhsllhGzhp7QVQ9TMcsC
Q5dt+11HN7PfO7kA3GNNdGIMnV02jNOj2zYdYrJ2oXdkbL//NhDjnmKnUie3CfNHiE66kHJEAcmn
DCdd6/GuXcGXOVpNRbKXRBB6VUgHvfnBhS9OjeNVe0Mf6xDvJr1qTWpq1wfHtvuQDiwQnSVb+3zH
LzL0/EMRplG/zDz/T8K8gbSAfyOrXd0VsEcQe5PWqANL1074l63mNK1ZDqcotXDBWjkNJpMuFLBg
SHrdWiCO2Fg2lZ33/4r4QG4gVSpJJYLGCK3MYl3m8HS3p20lxvVrYGpWtlGs9nqf7vLx/PBmWfNt
pGRqGOeZSr4nthTudMxdKvOk3CEQ5nZ155T0nSli8gv67XZIi3LR28siaTKyeWL2yk93URpJflJy
u1TVBYD/C1dzT62Gobu6T+3s3VfmWZ7pmBuogi0IIdxuvEA3n/99CaQmTwx5KAWjAgBhMn/9zU0s
dKEehtu+k0fp3uP4xkAyeimbnM+C9ePqBFIqD+xgB3fJwVr4x2yBVUEbwb2vx2J+8/BfG1iZ9C0F
oTKTIMHJk32S+SRar4L63NE+LCa4qCnV3Tgk2zyryCLMS+Le+4MeYlZdxZXmzGKTyKVz/9Ofiai1
j5Dc5V+dVSmJph6FReacwQEPhZRpZKE4rrlZjnuB3S9pfAJQID+TpOkQE8IfoZoh5yu8ANoPJ6I3
DHpdXka8SYl0psEazQUZLzz6WmBKeFCDaYmohNXnY2etFmq/VYrlWzCluhsIUNqGvyIGeTBKYlB0
A+h8pj0hRLXao2ZIZZjF4rsbeKoWYZoMKmNBdT5UMroUTfAWbADSc+t7one5M2F+Jdtt/9nsP+sc
vmiCuboL2qyUg7lmb8dHGImYZftwQaxFP2mFRATNaU9fyPLxND5Wvlx3NgnpRWMTppgPTDRafxw8
W/E2bHPikwrGs7Q2YPXloA1DIS9AlIhc+Ae51AOPw1CbCVP+GlbBEik08mUdlc57rY/TgUdyoSwT
25al9zZYvkkFUW6Haj31VqzQbTb6F9boDdnhtJdCvDNQAJ0fR59Fr1gDRqMPZW2fMeIHHA+P/2jy
44FArwJX2htI1b9g/FNgK4FRG8fizuuMdijRktLxiJyLadX/iRPB9dZRKQg7Qd2HzczAHO1IU5WR
gabP5FuJs2XpBhbh4NIJYazSDXFAjPLSh6Onl6l8wLQHtvxMEBaTl4m1+G+c+LOGHY8+YBn0BIuR
BOfhctmsXPT8Ia6UQ2oJ0w5Nm4GGReaLAqDriNvKq2wdS2oKDC5H6HjJ7b6n/Mk1RxZIbT0LmwB6
o1vZMx0BKt5TZN04/izynsJB2+ZQEMChzaPB5rfdGx33CP2V3PGjSoHv1yMeWIjjjmc/ZKITb/l3
6h5lp8sZae6KiKmCSl3LHdhK13giAij83GKbwa73O0vLJNsQaUuMVbMjuUvTfb0biso+vUBnTpKL
d6us/KMBV0b1KchQLTc1HMPJktxxdL3tDzF8EgXfIwCRVHwLcYgee4ZRbDfm3Uej+Xl/fHmABe7K
KSI0eYnik+3XNxXejvAIpe9XzIzGma8rWFfmdOU/L4LW0dm6LYiSAr1/OAG46o85zrjsIvN7NkHQ
fb5TN5K7hfmxfQc1RcQPRi06RH6NJKV25uteIYJaKLBivZQrm/aUjB+SDoGHBbv61OcODVI6W3J3
fCwg2aKoiBPoiscyyR6os/WW6jKfjSaTwyFV4KtxpQdmROS4dQWVbj7tSa7QwS9QnXJPxgAOnnBY
hkqWSCCxCqU/aHil3qIilpCplJML4BXFevLl1qJrgTagxnUPj9/CQk9hPeISlv1CgXxnvDTHO+74
vwAnEnGU/bOA8R7vsHt4JZ8c2G30Y/tqUgulYeFlDOYDAyoioWWH6HfgJZBBevO9QshsmWSvexlq
rSez0pdhrr0vJXBv0qjKiBdwQWMM+GWkl5GAFpcrxGDnctEsBpkwxx1rFH4CR65H4qiI+nk+lk8m
whZR7tLNrIV69eM+fgl3XIFhCbV4mRb4AmuU2HU3zC07+yJGCeH7954YnIOP4t7s6xVrtHnarQLx
0v5M3GKyti9/Vi+ZtPUvQWDmlhv4ZbaHuxWxQo9yAQC2p6airEtITcZvfgLOHrs9zIS6rInl4D2R
T2uecMPecGJif1MCfdX+u+qYQLl2gKsYUAsCky/dpNHB32LquWbDhtRJgo4lFvqh54ZsBRWfzzlH
HuS/nGf7CneXbQzeRGTmqM/9JcIWpLhct3n6ekxzTsZXCisOBmJM6lszpcAdMBGzoqDtQEG2MwXO
xS3tU9201UmpVbaUYnDyIZDTV0rxsCFkQ4y728NZgL4wmwCb0/c5kjI7P4ILA2zRIohtCCEG9EtI
Pj6RFkwSTzk8ijWcp7aWuZeR8dB2AR/F3VG+mEoj2SYcLNeHxw0uTJdKfACTCwQk4QpbZonP+3KD
whzLfOkDserwrSOCKRJHavQ/8BbS1i59eWWGot9pvyUqZMT/rOsD8VsuKAVMXH8Ny4Ilan6qNgql
PXuGwRZiB3gNpUf/SOtDiUCUpSz6a2bQspGY6HHELGjAqaxgqetICLWtFPf8bEUdCeLi8Ujv8GVW
mkPfraEZ9nvgRZdTF0WZ1J2/EhQBx9XRbgf6iztq4rlfVNuv1lplIC+NG2YxkuXRH6dFW48zTzXz
d4F2X5N3/L57h2nZkIyXgD7AbcYpeHFdqZ42Ai68NNgNMFdEf8MSkWsEcBm0fX8NVxnUY5U7HqGn
PNSAkjAnj6VJ4NRdaYZVNp9ll2g4x3qM8J4Hk7bC1l+E5BGtVIIe8iHCLeZMsmWXb21jdDUDSAcu
3eLFuskZve0bfP9gnFBSZUvjGfQmKV+74VbRDMGx2YtRviT0KLJmCzboToSdy3N0EwUqpTT3ASIy
S3/MsYOqHmXNBk2+sk2+z+uwhXO1/rw+eBHyIZZfEQmsS09i46X5DThJdtJrkZmXrwKL1xkOrKxW
QbFep/GfyMmslPgVNydowEbVh0fWJq8lKO0YNiUXHhNwc1rhHfKXbJNJFFUOArXgLJTM9i4c/iD0
vgUfZvpJcNxS8IWHmVexujI8+nsc3+go6jprcwJ9hYuqA9hlF+Mloim8lxQMvVkANgoz1h3DtApK
NMrlA9zpgSoXN9ULe9P5dgPmxH+JLgemIkPA4vU3tcMOK5q31NN07g+Ek7DahPYbL8vZcr7RjMBh
T27u4Wa54e98TRZcvwoyRWKBbTqMRGKHVyQNQl+12/7UULgL4AL0O0MOdXfVWP+vq7nrQHKs4Cnj
rVNFl/o1Z6SMx9drhzRnktQgeZq5kLd2qBYSgKqs68fOX+0XdFQQ8gZQT2Q3SLFnmK9/DOoDhDlN
xRZanpNbH6svPc6lC18s5W1zmQbNCEeIl77huPEc9mB9KQIO5rrjSNMJpykmJmLU772L92D9Y21o
OwqzWcOOfaFTSAc7oe4g4cd85eIH2YFmhsopHe2OAag2XWb6M0yS03Jti7Bu2eEaXx7YuVAj6KEc
uDZnuwYSxb+MSIQWpYlEUuvHd9SdkZw/x/JxHW5UBMgvBHcIM8Xq2X9fOBnK/OVCHmxuG4v2Jr09
GJLTrcXQSKexW7tzRb7BlnD8ScJgC4aVGuF2jeTp6Xr4GvRqgfD0faXWqEhJP2aXeLdasdU0h3sL
Qk+actdqq5pMQADDKB6Pofc2DuSgS3zN9Oxy1gAsvW4B+nQaEObcgxw/2shLvrTMCSttmpZ6uII4
XKP1qzxhW4FQUn0uVAKg0Eu92SbBpzTa+xTMgGvOYHFrZqMAjV6VQAhsWT8Wl2kWTPZHjzwIsOIs
3i3wD5W1qlH/T9UU5sFEnXJb8HEgGemceiplFVCE/5JWDNfA6LMJNSB+c4WnqgalCB9gm/3QScWd
RB8pQOEChXgoKYn8/TkAgYHOC2yo/IkCPoa8Unb8s/ipGNqj7vwscRPLdt7JJbs+jCF0jLVDviiN
L/Y4PVjuLYH2c4j79D4QOEMnWoulMjN1uuGhcroC0gF1Q8aB/ucWL7w6a/pBhv1fqMZ+cbEUUbC8
jfapytkIoP2vFgAVslAxjb3lAZaQzzjCCvcfCutr4xE3fU+jvZ7z/tDfwMrU/+yvTqepT7k5brJh
e9mtVLSf1hWIj9pvKxbTt7zQE3WZWUoi2FgrphLW1mJMJ64WpPWTG1vuKuoaNAiEm6dN8YNWZj/5
7FwoE1uMiTzHpHaszp9VvhedgxG/fbx+D6qRpDcYUgYwaxdspiYkXD99IA8MzvijBSTbuSMmUEjg
ZOImqQ2aY18BsdYaed7i1HHr7+77728h1Ahs68P8EujFxlSn9ecPnsxRnx6IZiwEeF4L+bhJuKUD
kNIqXdIyOF1xBLyuwxdHjrHEv7+CmnZPTZxZT3rvXfJjnaU+/Og94thrdpzAtZaV5tJpTabHzUXE
WK665rwWtW46Vfqrslqe4UlAeXHeN0mexU1O9hl0MXY/SXEPx05xncGavmF/ED28rpjqgz24dLJ2
x+62djLJ0/ZXMxcdh0SGCSc/wkrIW1cXa2/xSYRVvl7dpeBGD3hF9dVHTDKSoX25h7R+AAspTHSZ
Za4oEqR2URTFk71yIN7rWuwNT1W840he9AtLnB76DXya6X5QXKedhRMR2qRmlZXZsba5y8ijI22j
mh2cA8hwmU0OcpnGpZH33FDdxhPmpfuloiRca7xWZN/gdX43WlYGEhjBNbkUI3Kc90ogq6KyhEo2
cn01ZwxlygtGtiWnsuT84Z903vooGyNBamg83GaCRbmJzhg38pHuGep3xVLEJmWQB72JIBIdu1xi
f4x5PIgWtSrc0xTQsNOAZnMeUtgZWsop8CsLhBZ5VqMBZPENZ+FZAf47zJnjG/DZkM58ig8w82hj
BpufrHVgNZMzG9gZZvUrMUb2/ouWUbHycj++Kufth3p3FDlnLFS2WRWZTeGQUABj/58vsnEn3WGL
QMBEYXOGUaLeCbA4qYQwI9zJLPUzJ0DuGxwtRc9i5IRCqTXsSyPKoJSdaixlaDHXzPkso+fOz71P
PJa8LcZyDeQTO0vuutSSL75aNs3teV6TKYQu/pQdDAlPGnFnWt/AFUyTrCIdgjGyo6TMdA0wScAJ
3GDyxOxw/LgodcWdjaVbfEo8w4m3E+XO2y4wKoCPwtpH/fVyDh69Fh2hh7ll15dIfmZOUOg6kiT8
x0k5oKdiR/MwoOvLJB9KSE4/mZhSq3+l9S3hMiBYjIlM99gi+AHeS6IZ7bvkZtSvloYBlMyq33D/
yq9etUqwtKGX1sYJeXSgxurupwNk3ZRq8QqC/SLwbLwhGnlPc6N9qeSip5KwGm+4i3jnrSx7opSk
iNwXmhoBhtWIR4LBmjP8+hKqe03PudTD6BQIabRtMo94jQUQssgiLLhzrakJ5+G8GTTEaa13sheM
iwQbzPn55UP92TfK3vAMWzc28IvZ8KfaA7IFvhpe/yPn45DEJuYvesrUSj1NJND7UnS2N6jJTkpS
n1gSXxRSVjVlbPbGQXabFWVu1iHBlaAjGwtP3XA33J3bs92OuxlUZPhuWCxgyfTNkVwrhTVxeW8L
fDSgi0wzuiyU5xbUU2vM2Bdurk3qGHN0aPoprhFefF5B7N9O1bEtVZJVH77rYmo3SS/VmcD4Eqi5
d12hfmI98AGa7XMziLo9IrouY5CEqQGgDn8nQVzxw44f7XtwaHllzw0QXPUH5sy4vMXXjwip2sxe
IunfQXEIlQFiiwKlPFSab81EbDXffUPwbbM/PvF4qT+41aidNgcQxsDleO3EBa8YhkECNRi2VN5t
6PV1A0KxrALyXjTUvvmbM47YjICvHDEkETOnGcRB3RjMZCfjn2pFH2XOp5h/Cr4yiZ9qduDjLkQu
GEpRT5kyraUSLgQkW6LN9j8cveg//zyCgUestpylNCMJkWoHZ3jeFWhDygODyxmHjba3/VeC/t2h
gL/sk4MyXWWFRJ69lDldtiu3CP32WTBW6BuYwaIpSzBcfQ+XTNiY9ACmpfY7iamVFvK6OcFfoR+P
xz2MC+Qti+2y70QtpXKUMyKTBVdh7zLpLMcLQOwvoH1dL/aaLMN4vEbkZ/PoylROl2vZ3hv6tT90
lS4XRi3dWy9YbbrsDKAYB9cBkN1V537zyMFzTCtU6r8y5K4879Ng4ufDzxbho8iPJdJyBfefhaSo
nA0VWjLfFh1wciAhyd93b0pPCSqA60qDRqyw0HEnVibrORiS8X4VlrQpNKbmZcpKcgw6utF3nTu3
Yo7xJZW1ydDgWj+ZS//8yGbT3vxR5MjB4hrUJBC3MBpMf64t4/hDo+DlEGn2sF8aCt8B5ve34GQq
DvIoAIyLpo0wtI/Naf+UwNmLHMnfas3B9Q4nB+eybxfm+xeKwMa8bEim/oh80pbEdUrmgydEmquh
P7NuL2etE+YfyLORQVxQdYa3RIYA565LGzsIYcJmb+FMjjxI3IWqMBLZfBOB11+ofHo/Gz4teM/D
QdTV6pQPs3xmFIR6tZHRnOrOFP1lamE+4hiMniJqNp3pzEPAWhN/z8ZZcXY4Ab5Mi6jSRU+6w8K9
dreB3b5RPll/fJtuCpeNcQDc22bK6/CeEsFNp6V3XIx+0f3ZALyeT9UX+YgmqaUpraF6VRk9eR3F
VtgJciGN2aFC4HudNpXytoN8Vvxr9L2vGx2RyiwP026YzLsYDHA9Xelz6KUJvd55tudEIWyd3mVm
2gPl/FJAiRjdFH1In7RAoK+RFJZtfevtDiBR+S/X+RNOf07VEQ/iFnePhuIUergBGUm0x/Gb4hJ5
fnxE99wsLu12qpQY4Re+vPsCqgnE8NT+gHF6/fEZbHaVysL0fadmMV28I5e4qXe5+WGQSjREfNL2
YjiC+q95XLrF5TUg/VcOtlTIkIz1AaRAMahjdaxj7aFNda068XPtpw04OHbAuSpT8r5OPhFYvQ2w
8pdn+7NC+QFEENxIOdV9NjieGz5sQhvRsdzAc3EP6X+yKwAOD9v3OTogC9Q26FN4Nqe7Qf38+ufz
tbPUb3q3271l2rIVj7oAoCv1XuDPw+8kGPcPFAEk65w3dBkv75UKedJdWp/UyBBcytpTWgOOgE6w
wePVPYYxKeTc67XvmmRdDTVaiswHRg4Dir5si5OqWiTBP8XW0V8+GkFjnlELWA==
`protect end_protected

