

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
nwVS2CJXupErGPDoD8Ku4o1Zi+AYJi9tsbcPZPL/xRo6X8XC10paKNinYKLQl13EAkPXE6QL6ydM
lbzHjNTU2w==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
FkhL+cK0BtU+W+i3t7Ytk7Op0uCvIYyj8H/bRZnnNtxqo5u8IS/D9K5RShx7R7YRWNheaHMn6Ygv
fDj070P5zgsj8a1IJ5dI5LDna9WXkeMYzmuMalHydMJ1kudEmdOLJKq5WxEG1BRQsQ8k0lvVBfgM
yAAoO1x2DHNTgSLvZLM=


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
nLzdtZ3REDuTjhApuaykPnq3M52YDJo3801ryWYezzWQ1ygkRNQtz5E8uPdI0FLOp++xKvtemVgi
fpsd1/BGm2yq1zzsODcsA0zWeOEVUe7Kva8zwt3+QlNFRV985vvD4PADEGD+1Pg1mYbNGhKEz+Wr
J6fh1jXqY/tdPQg8ybk=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
SXLI3j9g38Qcx+QksDW8F+Y5+N+HgVxbkWGUtbeEa4XpHk0wAY4iMFbTv+HcN+rLS1JoEudk3H2C
21mMje1B3NXO8DeAIBW8MdVNYvUin4DNeufylRor7+Q9+T8l0TKYEjLntggmcDF9aBwMxPgXcYku
RdSlG0f0o+mSc4/alN4xOpAWw1p6czfQ7Bnq35E9wIclYfqCrWOKBuAljScCce4lHAkGi88+FzjK
g01jPDvOfPqK7J7gDmOV4VSR8BZsg4pBqTLQbnfmYGUwhsGr3Nj9GemdhadU5MmfYmDY3imY7ZeI
kPUIS3pjESpw9iA0OuTKr5fKJhJZ2cJ5CvwuzQ==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ftcg2N48NqCHefTwhpYrUPaMvMzpmuLqgqd3DtpYFLSd6DcixuBjwhWRln1WKGqWTyAm0n0iCabV
JiPhKbQAnTvEOylyW8uLjd6IH7B3qhSAy/BYI/1Bgnqd48An4sDXFIT9ou/WloM/6gVc+wY0BSk3
tSt3jTcfvZ5JIi1GjRXAUPYZjCQRrC1e1saS55grMZETTHa/hgk7xaDBhgmHlBHqrJeGKkNc7Tpj
OXQFfzDow7U3v49Kr2+5nFPJgGSKRUkg1X9xMzj2m0BoyzUNgYP7wZ92wQODUCegN8HM3JzCt4+V
1LvHyqIFm8cgkJZknu/d1XRyxL1tOTHlqvDQng==


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
UwEUSIba05kuRZ9C3VePFeG4phawLRcMXZ/OiI2pQEyda5H3pdyOO5c4P6VMWnOQK6zVjMlLJHME
a3HoxAS3EjReH2f/s9l+uJN1GOCXQFIX5mDFVCm9sBuDewxIsFZlz8PoKwVAXTjVVqKQJ7MZrTZv
CVU2unSpN7KHWfuHsfJJHMR7qoMfVxRHgpGUZmrnkbejh0Fx3rGZB53oWe81C0QkicrQDjK1MsQg
jug+MjAYVrdnlj07wJtTfleJYMiM6cBAjv8hDLe4hNRdVn8tG2btAMW12tt5GFrJEJqwWB7Ia7Eb
VxTM3bbsE2y8nRoy1mFThD95xJ9/8OzaVhSAAA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 204624)
`protect data_block
ZGrNTTGRptVpbMLQOCuO3x1UX7VvRqu/ez6mOppHWcnqeD748UokB/JOku2Alr26qzfyn/ssGT8w
OcUhgnIiT5uFWy7Gp7u5BVBzs+GxLRV6cmlzZeH4pzM4JVWsPPg4Yv/B6u2gx4+Jy26crAg01nsN
qwfSpLiXEC1NoBcOHzihfUvsf/MR1tZVLe39GHpqJyt6MYsvxfbL+cMT6gynev69s6Ro0BPvdWnW
fCyt81A71tTAIhK0F9B9itGQiaAegav3wc4EDZXu3UyqFdZwKWeqXq5lQR9B7Gc6cXJ2FfzjTsra
tnAMUcHKgQFbBR7Yd0yNpBJEurVEBisQhPdGDy2ePmgN2An0JeB/jhvtayuO8peu3Ju9ERxTu9U9
2biMYypcVvCJcJQmfinb0KqpfvmCYpD4gclHuK+WeT8pwRK/uv8Zgy0AXpaxVY0U/QRqY32dvUlv
/ik83mVV3Z4AnjHp7bBrH2cEEQtQTxnvjr4Dz0aKfAYsuYOtdq8xfm1KO/qnfkVn5/knzN3OfH7j
A/asLUWoL5mWvViUkyDzYcfQItWVZ7ABlakToTuFTKw0xVjM87zuZ+I8c1rZpGKTIXbKaqCFBoUA
3KOfJudcXttqpCTEA4A/LGkVsAAZpo6aWUhjv57tRd6+tlhMHRK9rWFRSZZJczKsjfQKeP0bXt9g
IoDRcKn2Cn0ScxUJuqlaOTr+rzlaolizRh6i+2BcmrWSpEBbd9VPb1aQDxNXAdl4L4wEdX7kDc8v
h2qNMU9mftXh3EPWREhH1R6XR18uz/I89z21YpDcuWUcUAzDJ/mVWbV1jrHpB8y7tTclbdU4epg8
Mp1q9oYyYEir3tBlg8eBLGlpbEjd55WxYds56BbXKHrTN0rLfhpp8Ybrdfdyc2/RDVtSaG/wQB0a
TuEluPP3/E9EeLVMk51n6yjwYJwjG1lFUMVwnIkfauwFmS/3gxNdX0HkyQSyQ2OAar4ErtvfzPhH
pYjM+qmiSsy9X6SYe0u1igZkJD6KQwzguz8lHNJicT4+91AVyJX1N51MabYawDaH4ti0VJ8wetzr
d95W4p4n5SyoDhfSK4/MZQ3LsjtN8dUeanebKAHiqUOiwq2wdDZa1znLL38WoWBN7/f54VlJNTP9
Ai1pxCw7e644xzeGlQ6ZnuP+QsF4NJrDr2zXZ10eCwXQh8VA0vrefYxBMDF5gRmJr4MUXJepBcUU
d2Ux1V5P/rx5KceeBerl9Q2pddXLDRVLAqphuGmOWb56zBXeutKnPI/od2GC7T5ZQvr8F3zepQwC
AotVHBJsbAzj+uHqzL/LSig2cN5E2PrhsecQBbB8ygksp4Ng5E+yMrx/RU0ggnvxHm1Bei1WvHXy
qSUQ52MXEh9ZVGiDwdRSjDr3lk66UBLJJFTvxXG9Yw4UwvP+S9X8340YI1h1pIdQd9dvQeMx0eoY
awp0UeM2od/ni2hLDV2iTOeo9URBnJSgdisnoagREaUFH4Y+SQaaj8al927zlowDdVFxxs+4+JOd
ZOWfZMzj4KVhWQd4rAf/b4VUfzyaB8Lqv75kssY3IAS0lhItua9FM1U3aCxGphu/MILLyMho4DMr
LWtXqdAOQ+2pfD809HYiC4OBvE5FH3ztZtjidTpLCKPle0vkAYhOwDJKywwSOLVUQsCDxB05IPp5
1o832A9tKley5sMJk7s+B8VCscVDTb6LBSA1+57GS/dySwFqWV/qR/k8xHiijfWGYUNEVpPQhoHv
Zyu/FHYGr3agdk2CbwdtB8taJEIVenKNOHDt+JQpfNQlhZA9atWE9VxdvxlP000P58uMwMxu4L7r
nHbQbqVgOMOm/UO3QEc8r7AuRKUTBM6L09BEmd89vS9mCHUW3wTGuKSQyTyvO61+W5UGs0Lmq3s1
rPLmthLGDGwJJw8dcaWJ/eIhPM1YdPszWQ+kjPuo0tpxHIw4Rh7KO/tOxo0rDzL4R+Ei1sIQNusk
okXL4t3TzHSV5I3uhwMpfYJ2zbTr3moVpx8jyDBUZs6ElV6R7aGJauO/6Tnkxhn+lMqYD21PMqC1
Dm3iWaDSsFQ2QARXrZqW0sIUHCoZT1gdUggnps6e3LSoUDugupkuAD/8vL3QPRU5Zk68rgbnLmFM
Deo+M/XDEmkcnBZeUw+639i1EGI3tvZnu3ir+EMgZ5VxJcgdUMcdLIsMmKi8snVBw6SuDxUpvHBC
qXEzmtFpiORETWw3o4Ly5v2Kq0c5Il4qVRp7hnWdLiebZvkbSszoiE6NxPYgcxGO6vssGDL7YBwo
EXpfb2oyjg6geB3oqQqd41jgsi6FP++wsMeWHm7mXMXvUgX0TRAsIOEWFGuutDbm8mjdO+7C0X4A
Dn6Hwx87I6WRz9FI/tdq4QihvaI0g2W0FBOaTctkmQ5qseGNkpPYrt7RXmONU4JXbe2ilnrYzHsX
a4As9o9+FZcKkxX5mGIiTjt9CJ86Eoxp3+hDxqA/O5/dp4YVvv9rXh6HcvjijalcxyrwiHM3tUB4
ef9KDyq4c4JbcpkkeAYMCAfU7Nsj+l2sSTlsoFAX4pjiFtUbpjNocYdr89qt4GX6TvjSIOEEUHbs
yUFmEmgaiFyLDbPXGTH9U1gtWdWwJ5VS4Cf+9dADoyILDr8xW0BgpnZpVPka2LrCEM13iZ50dJxX
c3WD8VhgDuxxWuJeJRgUFjT2FgTseLbNMcl9QItrlah/B8iAxZ3sD9aRaXB+7fY/S9LHCGIS+ADz
Sk6ZsfPSH3OSNWiGLj2okIvs4L4IsQBH96eKfwwd4oXhltkVgcwXWUgQTGELdycNvRWFRAFaxsmL
hHX8uEuMmyYHwzXqRh5su05KK6TdkGEZloDeZa1bRUWnFvz/LnN1+c6P6jckSY9A7GrasF77lJFk
ieZSlWO1nsodwXpD074Kyru+cepjN7ddbTx8P3hfxoP0JA0+n2ztHs67BV5O6H31s5k7v9K3dvwU
AJ9emE4HMSu1WLjjrd3EvRx+bc/YU1ydeERRG8mKZR+7mZdZ6vx1v5S4zl7zgZqZNg492LPYW2dg
cYaOlREgSWd8lAf1F/iLqLi4Td7C/fJ1y3gtYXscK8ZLpuF4Cb+2B+4b1QK++7iE8A6kxKUwAazs
w0h9tXiaexZ+VyVSbKXF8RI1YTiixw7C9iPAjMX0EN2sPVc/RVBsyxrStY/Q02l4VssYN4Tp6ANZ
UKUkV6dkwed6Rb13bY56hh0NL0HO8H1VQsw5bAxj0fgkg4s21KvsdN0CZIiDgWk3oaIvNFR7PaEt
4fbg3hOWmBZu5m1GltWlAUs8KBr1icqA5REmm6Uj6I7K4YFE6MAl+WXjhNY80cs0qlJZ//ukDYOd
XWIO59FLT8QYuRo/ROPw/92nG4lcFsJgnuuOla9JBIn03Npmojoe540a6tu9OUqf6Tyix/0Z+go3
CIEzG30JspO+m+1MZUI6TmhuwVqXGKdnmqgos+SBVno2j7vyJ6jRBWNR0bmgW3gSMWaiWdKVmIEu
vRW5P1TQlWsSpbMS/MkouU3Ch8qHifGfZz70TGCchBb3I5xytyhwJugjteP//EbwTcpTxtF20YA7
6wk+BQBNhphgvLL66CNpiaYyTy6XvthKPdKUAs1Mcc+vOJW8cGaUueXYV2uWVsprFbgByEM+AVv+
JdOzS7vZWX/PqOWYeOURaW++k7JmBu27pR75TayvgMLZwpY5nz1cQfGjUCpbpnLTh6mCrKfDng97
pk3qiTUBTRqyhVaicfB3r0Y569/SO3KmATd8M2PvVARkO0d84t5RwY5RNGRn7MB/9qMPva0oVorJ
KjbTkj8g0u9jHDLOvBjbQx38BCseNyJ7l7buPmnepnndvM9Wono1mM9gxgu81vQ9M80UOoW2XLJk
K7akmXFsfLLtAjBnhDZyInTPjkQXQCcfI5xzcHCjUfmFBf8gsGE6ZzPwBqb/vb0ll1V2jP+q+SMp
gD/6kqLayiYbbxLi6k48VK/9nqSqoRhMuskq3VI8I/l0YsSbOVNQ1Mt5lSTpMlDGaB6DN/6Wk4bR
H+JshQ9lYL9sKENOyTfchcKjL1UYYHs6MJYiQslajo4+QsjQqBbgixU2NO446tF4zpGHl2nKo/i0
9wiQytTfc+G3B00WAYN7+hv1sp0p/+77IrcHvaI3WIk3FDVdW/eR/NsHZMBZ1+7o7tx2YzhdAnbq
AKlxgh0JTUKQFnGNEDfyoPNYnOz9QZ9IMk46obo5MevzbHqjXi8UHytlPDcEYfElduO5v8eZ8O6j
7XV3LJpJXVM3OTaKMdJ6HZj4n7tSdW7XbEfPK/1sQwTZSqa1YZcoMXMmZraEnxC9fSy67Ynlz8Ni
5OtFWKW4QVeMZaic3aLQ1fvz/l2L+we6qsoBnNJIoxaPwUz0lj2T4fKl3xgOQlbJdqIi6WdtTY4/
k7QpEgeFQlOwmgwP1ae7NcEdkCpYEDrKDoprq45rPxC+HbXEpcEB6IM0eIHFF60HOgaenR720H4f
j85ezMRfO0YKBwEjZJCcjb+uBoJW7YO3i7zyOzv9b+jvUvGuFiWpuKWyDdIXA8/vzpwn/P5TPHJA
e3BVCmtq06AA5yHURA4w/WwYW1QJrjRK5P1rmQtqiFZ2UdCIhkcbP32GvNNF4mNUNBTiSrtTfkEQ
NeSrjIur2R63myTlPA7BZbhcbTs19IG4aCApyq1XpLvA5eIs8Ueol8VtvdAA6ekbFC1YOCyAekzK
kcUEQR5bYBjNi6HkImt+NfvtP2gPCFTKfouZVZsw12AAUCh0RLrNR5Z28gJhWTE29ZstMQUvWsFn
ULzhvgP/pY4xlZBO7YKJXJmPZdFz7/QaViDc0O/4myAOWjidRxBDSOMmC9hn1JSKWswQ3n9OJ4Ie
7fGH+a4I9hiiLSYv07m4rF6Ekzqdl+boPd5Ae3/rWGQbK/B0BlAQyav2sMgf5AO8UV0znr0mNyJd
q08E8FlQ/F94V+lrkfBzOeW43TI0lWV16FXpBmbXcXGsjscI7oX8PML2Ux2oRlvPQosFszQ7NCu7
iwg1iaHUTUWEdU26I8err/tUbSjuZx9+TqNo3Jcw2p+V+0aFepw7Iyh7RANga70Y29cBEpT9rIVy
PhPyXYv5ZHLgFrv3YmIVk65V3zjrRdoeqQvhg8KNcnWq078gdrUryWdSuuGXOWF0ziIFPFhTIvar
iQEVxJjGnN4Kmwf1z+4mQPV2IyDviazxlWqTZ9M87vf3ioOlUnpDYvH8y4ujKE031yzvqR4gfC71
WTbmsSrwYIM8+P+TUNIEVMMQpRaMM2NrYwjUkiKIRErX72EApwUrPgOggOCgcfwfggCiMfAPtjJx
WeXxe6Ne4K8E9DCx9UqGg23E2dBmTP1tcGJm4FcKdXh4PVWp7nCr9eriNdUVjQAJgDfCt8WbhFqZ
+qOCviJSaxEJdfYHqVEq9PL6G5E4ZhAEd52KBlARri62BEMuuD15xV4s1bu31E/K3zcAMb0zrpS8
ViGnF7Bv/2nNAlM3Y2KZ860C/QwU99Y3H2WTs/vspnWOEDqJEXjCpJtWZGW73o+vdofutwZ7yKJ1
Q0y6rzL7AC2q4DwOTtHNVPiP9y9iDlAcIE+GHNevCfnIjPJ1wxnznKtYcqjGfCwkIqG9MaaMa9pZ
6f2PZjSgE1naHg38GCp+vvnREIg6Z6FErS8PkyLXH86X07TIfjnv9GnkVn8YCTU3FiMK1BcjfPLN
Q//DuaVDK/1sJtBzP0Fd3Fica30D7Jv3I3AJsjJKNNTbN0GC2M2vy5gee9Y6NP3nh4/2O+FTLBW3
5fRYCxB1em3rmc4xPieJM//q0/Lh+MJC+uoiLaG8HAZ720xO0ti76FoN34St5jsPaAGEMgQr3xfN
Zbn7ZbLf/Vhv3TF55/PEuRWD5a1ozyoFTEjGsBN4Ug0wbDOdm+wP3tqXvwuTFQvxmb2BqrNc1Fp0
ZATeghzihA8W+8NHP+oTNv/f2iiv0M5Vl0OBslHgy47VfhWU3aXDgD5vx6mqtZdF2PaxU35Fmn0J
5elrdT4jUm8CQq/OW3RfpnIgG7uGHFM8EHhGU/aiVRmfaT1qhYSXEMM+KvyFd22seOKW+KnEy3HS
W9wzVEa0aEwT8zVZniaPZxmujh+/7wOmiYVtE8hVvOimrj6MwpmuqJyx1FCPo01M8a+0kOPHz5FY
3EPM0g84RDGMuYyCGALRn3NtUJRMBUsDZdVDH4uoZ7XwMnvQ0OC/Tsu3pFM6TRmrcl0ueeG3DPbM
yuwWXJFmLnHPYyD7GZhVhCr/Rpw/d+ie0QspVUVcesnBb36uZFshXYn5xUyAbXzZd/6gJUp/DI52
RprYpfMMqlt1q8iifO6RHaKFIOErRXD3hzOS/1QFs8hWT+l5X8vrpbzZhi/5VAhlBHsCUQisXXB7
q8kqj9XuiHGbP88Uq5QA8R0XSmpd0gjDDcRRQMtUp+gYAoCmVwar0LpNSdl0STQcuna/+S10+6XR
Vq9Ui6EGURPcdILwqr0GmsVRPwfkj1Vn1U82gPqsQtuOlJ74VgraMYJQkVbnFncweIHCieEiO+Yw
T3hb5XE5PcmxP1/+H8EVwzL6ZXUi1X1vdDSzxwp6+G9ud+u4fws8EjM02LWJc2+L47jTD9Rowr9n
+ecJzKijLyRjTVhfhV0Bkwaef/y8iXaWEW4G//lISsb7ruNIz0MYoznT7ljkDIH4gy4fo/TXazD0
Y0jVL2J/t70DPS6YN1464rH5GApCYJcY/LRr+MrjsROPFksDMFzvlehqtEv7D7X+WUMINWlDaT4n
b/bIIRHMLXodtTwBZvY3RpYKAqY5z5ImF60H0lAlok0ZmNmlSowKn+c3t4foSLuwufTxqh1VSDms
Lzt2fBef/d/2dtX8+5V8jNkiwMK2VWPjYQ3KEPUViuSL+WZ5k4PqOQUzOjU1tWKZKlEqZihRaBRl
2qkcy4Ul9/d52UBYj1nbjPXsHcgjDA2MgIaJnEKJEOZ6ncye0LO4sN8ep2iuawa6f01L4oQWBtP0
Q7onshoYvtPJZCeELCpa7cA0qNDR1klN/Ap36JJlsHT4NnOBjmNSN+w0Zj8f5te1WhUwT05V5L+F
PIlt3bMeySoTduwvMciYMcfoE55Z85TuiMBnMwMGPKTRhBzsZc2xPmVoPkM9kLEOQr/kOIz7ZWZK
z696UjN2wz/HUYaHMCoogoGMcXpLkBEXlf2Xgrv7JrPsOqkaFWdnG4V0HgQ1YlqsQMnpECseDfY6
nncE7r6LE16YCBBUqt3PrtDaNMn5QTkFgLnKjBwWu8pnxd/O5DY0pJzMrAJKi32lzYjDhsgfVvgy
9ScblPTkDv80XCPxOvGbEtQGR4jMfnQJH9pGbowAEVBN20qa/TwyBqRAUogNdoXy5CXeweFubmp0
cbXS4g4GMFz/aorbZUKRdRNSltwZk0iYuM2LtfPS4jCMmbbtWegHfeRk/o16OOM2oU22ku5k0/FJ
VIjK88+beUYdbxCS40kgROuLBO4oH6ekj8Kuf17Rr4olzz0IujTJ5RPpW/k1/uTyWM331g+HhtEt
mz205kgMm/ii/WrOU8RZURSV1tjtJA0GGOQWjyFeLGI4KCPUrzW4KxRxAXRV+nRLQDm7gFeSwn7E
05Sy1+WWQ/CNRqNdi1y1gbYbHVsGVGUtFoGCkxzTDk6qNJRAUfDZP3XtLcVsQjuBTQ4HFA3/zpB4
LW5LSG4EY+LxcB43aQNh33Y50Bx6s40CnAgic3uHBXOQ6k4ukTzijgOwAfogZP2361bpsoPdwgD7
jn4WrpoWcMcqUUqdfh70GqJAJ4woKGLs+xwwpfcULRSyisGEvAovvxhtD50NA8XHXA+zjNTTMmrA
BPD2L1f8sPUK+tfMTKGWPUzxGThzuKaCSyJsBbWxlL+eKawntCqQo2IB9Q8tRPOraSfEHk36TOIC
C3edbXpwfWUUkD7QuyosJIkYFDkwun/CHfZypmBcxQVeH08TSuLFr1/IVwkuWZQ+Ur/NUnmH8Xpm
jXlI8QtZs8Zhdn54yO8r4i3eMBCKcliH1ADdIaoG80Xp45UA4d7qtWS8wl5jpr5stiINIvLIRFPk
PZ4gi/X9NYyuk9U23Y8ET3PfB9rb2SphmIaiNAP5pnVYAe0qyWepn2yR5E70at1Y5VuN82LLClmv
kTVo0Yg5a1Fa1wsM3jUd4iJyuMZwGD7rE3LRa3oGGxk4dSmPDlkP+Sm/q5qTlaTsewJFH1J0W12w
UK19UrAHFoh1HGhSIgCcxUYzeFHXHGYuEUYzUJl7OR0ZZCh2TLfmZqPpe/UWGEnQmy3E6ETiEnFD
0IMAPjlMGkEwOlAB0xYk2LAjChkPXqSHlN4HqUF9P8ROAt5xua81/i4BoggtA9nWuT3f0w9JSW+H
ENYYFe4CyRfLzEz3iYy84BJZa3mMwi+LdbGyTCrMQeXXRG1rL1o+kGny0Tnk8IBxirMwCRT8Srkl
2lxZjnYmtV2eGeyQlqVVW5GDar/m7hbIv01vWelT4bcbWKtsrWIWAy0zOaMGLWD9oX/u2tKSfT7C
zKCQ/yRDrEYBwLQEScTV607vjRCUwKx+ZAfi1qAE86J8nzJfrOMaGOhsvUZkyhUigeSqeQqFkRye
e7w0Q00XJBSvtYscpIR0reZOmt2dJ5OH5QgC7p3mYbzAeHtsVMg5iTlQeq8CFTnFeDuz5fxlYG7d
G0caDFkp3mQgFxb42accef+brPsg2SGJ0GuRaen3RWw/VE4X+dZIauvoCK/b65b3ipGD9T534HSg
3ni3tkWU4vPxL11knbH872v/vSl2EzEO6t9lGFPKxmTnkMfl3X/e/7SEI0pI57zzNgdkX8LFOFjE
gDfr7/GKmDQx4Cp+lf+Ss5vJk3IMCFb1yXtTf5woinsdYgOozD58vQ/Te9fp5UeFY/2xU0/TRM8w
cOIFLnvb78OGND4TGYzLTQ2nkaYWtVpr1zehrciFwFPW73Lb2Q0LkDJbUGcfeJIRbWgqoR4XseTD
ZOd2r21hgtXvNigyTVu2Od5sTh5F3Bn0OLEvVoz2Z3vEpb6kFqpmGQ9BFUXfuumINkjmXVkSyMAr
RTS6i3ivxLnlJeB26bId1BNArtRKkNOmql/xKT9p2sU8pUMgqfMdXYs/voKb9O3gglYimp0eElYp
JOch302L/wew3HtUIDtYkgInPqRoFMi/X6TC4kCPISmdLhuLkaHDV/hDFTGVxKV6G+mJFfjkdCSF
0YqqZRASgq6CqM8NXtQnyyD8dfH1pwQoo5cF0nm7xp/C4wdYWWXgT6dIcxWieRYz/AFeE1gSGj5/
2KkYHaaP7rqjpWgMJ4ZC4nxtXzwYb4vugBg8VqgmFe7uyAY+8dOPdQhtnrDchox2mS5KIIdfu93x
Wz7Jy7akTE/XQDY8sHCfTgnFZEOP2cDistVmyopgU9ipSq+j1yZQToLHUN7bVzaQZ/a0ZVcgS1P1
dcqjb6918xHp2gJ3BRaksE5pbqIkuHaAA1EqeiH2HVm51GwEsZv+3Rom+0cDoX1oTASPQH9aBmZ1
NbxZByNAs9fK3M/ZK+yD2wHlmrOZSFr5PS6OAA+7mj9pOBCGhwJo/ZgfE3K8SBn/0xN2+c6gb0t7
im6x/CVYsxpt329P1boG1YpqcjsTbq4Yb5oheVl9ZYo7k1HvI/sNhTmmLuM9tVQRItzxa2B5KnIO
9ody0GRbrAj+/ZeI7elaeg0tt8+siyWvWZTOYCicFO+CG7K0pheS+m+h32jc891ctfZpGCey1vAN
fgjfbzJKSWtg2NxRXZoWEbLnY6hqkpaxIOmVimiTyky38e0qDI9rfIphg+mVkFwbwLiFVYJq+DU0
OYcfMklkwS+jCZ1CEw6N3W3jOn8tTfKtl8AIsbRTx66FbZDKtBpiH7iVmSz7eOctnwlWqz3gayP4
Qp7Nk4XI8+aYdHRT1Bs4ixzvcZvhExDssJHeZLqzAaycZZ2tYOa8geComOFRNQO3sxlJmzMX008N
X9oeYH2qy3qpBo8vhV6zedwBJ+cYgb9srt+7W9zmOwYa8gwIr4dMSLOdPWhUHPN9ZSA3v+lxJr+N
TV1CNTwZ+9/f6qWGlFZN6Y6wCQpm9TVHzZXz3PdaGMjQubTKRlC5IsiiT3dm8Em2PhY1Pc+NJ+Tu
6jg+YaHfKvOwk74sL59cOG8dD0xAyC1m7qNEAQOnmYY56CxBxeyPBz11cRj9RIPQrM7yAmulB3vm
j1Yz1LlC0xInMLkNuJ6eWG1WNbB5S4lsbEhjzccuitEu0/mjRR8yxOIH6q/5AnamtEPIwsaKVFVN
fiCgTTXvIct54A5BA98oeHZjfhfw6FD/eTimbONe/JzZu0XN0fneRP/+e9rNyc0FEP3RXmsN8cpH
+mX0eiTYy4zoJlqQCpWUyWyvmfH9FYf8Y3B+qPfifd9zEg/j4YNTqmE4yFpn9ItCvlTDgDLEjtKe
MDo17H2t7sKlSxU2E1EjDfZZCWw2Ntf1IzFVNysqJ+jlJYbYP+AWGxds6dz+uIAjsU9py+ebAUpS
m/C2mFeIci7FLNE1i2fxqasSdOY38BylnrLqD5j9lXvoXsqyAI9bwiPSQsNJ/BpnWboYl/zTesR2
dDwzqUGaFRJEUzGYh3p2REPOBad/kdf/T7U2v6rutjVWnoPa7hIRUkeioORgnToM0Q/v7bY+WjRm
rMXzBxbpLtEHEZtwWkQKvWo/vSTbHoZSo2GXGGg8zw+iWAg5TlFAoexBJgZvWKLOvw5rRpWc/qpN
C4D2sb8X++fFrLClfopMxY1jfb/LQ18mH4DigEfgjXMcDjKM3R2XjUh6aFCB0YEvYhndyLnZiIwc
Rler126h768R21q1ea+Scueo3kI+2tGRsxgKd/QmSJWw2j7wibQwNmBYHobqsUArQrIuDJ3AtZC/
v9cD24fsGruZCyZ4KHpPj3o7Rsc1n9GkTEhKQnx3pcxllY/Y4EMf/KyRsnaooNBbFdaIQCuRe8th
MRcP+WTPnf3newAHeRtxsS3O9I43rYnoZj3D6TB22HJphlyUagUJIW0aT3g3p9wBJIX1bk9TaDu1
l4GYaXOEp8Yg8cqu2r0aamzyRtHTrscUmb2lKHQ3U35FTpc1vo9evVNom2shXce58RzdDLUDYTxC
SmpMSIjQtz/OVFM86vLaqUQguYNR7MEUFjPxkDcgIKEpNe0voQiW9ZC7TV91kQNsBXS7bWS6hwNi
ZxdlYiMt9x2MoYhyS8kDYbBpY/mtt94QKogLlY5viLWEue/ixakJibyPkPvN92Ku35tQuo5lbjKE
u6ZRHuUy58LcT+ZKltgboUVymB+Qh3qXmVHQe9WK1KKSk/Pfdxj3hO4e0ahbsidKjh1sT9MWErK5
mtENJ/29o7OVDsXEo0G8xNtL+OfXu5O0x/DAM4kPlLCzDJ+TnqSj3iGKr5hbPbjLKG0iFd6W4H3b
Xu9y6dimCbjE2DbmrjtKrfE/KG7fMUuhiesCL7fpuQDwRWTI5XiJcZ8ybSBqV4UAkYg/x/gYjJvQ
3LjX58MIrfOyQWh3dxsT4SLyLEhM98GTl6XadC8UT2qk04HW8Tghxruw0LpzrpfKdngXVGujMU7u
FaU5ZNjK0cLf+Gq1RDI5WxpPMGhD34FlTQB97/9ogUQRlcw3C+dZzDYc6egMyn0OKW5PyJfYbilh
NTSvtmMA/sPpuBeF9AZeoDDXR5uE7v7X+rfAhvM7KC11KD2/LOxUbBjddh3F6lo//0jwcSfFsRd5
mKVd1PLloCbhoDvUqG3v9NNOtQWbEkcT6sgIGuKNcMbnHKZFQeV9OUrsPAAVZnml0djgd0+3GCTs
7Xqw0qqOFXp86i1tzuvZmKw5H7j1FzcmGI35Dvsn1j5oKOSOXcPSpFpRBkYY30T/3Y0sStGyWJQ3
rs/HmplMEduGMBS81sCENssf8aJ/AEaIfAfgV8wz+PZAIYyzrmHtvfSCyC1e6KaFRXYr9aVW8dMe
AkUsqAdkFtMhYqrIm9A+uoA9TyUqkC2OKYZai8RJmIZXX75uHPTk3lBxB2VAovz3KFlWd3OS+E+Q
LmSixPkma7Q3vpbroaqv1tNPs7al37VE0dXDDbbI/MpmlKl7Iv6+gkWavUX+5Y1D6l7hdTezeVLP
xC5E49vpoF1ve2DChUpKd5bjx8dZWG17XquqvW0E2mMcdCWeC2n1NUp3SUY8/diBpeU4/GX1dx0B
KAYTd9PP/N3IUlfsIu+cMnL9mgvb31fHViHuR7L4YcPTegTtHwXEVJrlIPzjlxmZuaP5Q0y4mxot
VOqBzB0k9OqQ4HBXJ6pu8sZZUJ3mxhkOjRkfgpZGqvZqbKi4kMns0ColbBeuNfd74y+CQNBh72eE
vRULcUK15zkJzgOmiNySoIkjZ3DbPG6csYmJyaFPEHJze1OvHLsQz+ucqvDfO73sdtVLjByeqtZ2
O4ZNa2PR8wN1fdhDd4rWOADHtRVSTUGmuy90ubXRXl8PBxrO9fl0LRVNhNwSgo5KjxD/xTM5jvqS
EmYUQpFb50HPUemth3+wVW6ZtPHqcrIDgcw2b01mPSKWwIVfM3V8BXG2nXvNmnuR8niPSLSrzsKU
9/E/jqBzfXxEsDabopTQg7t2shG0Tx4fcNz/tMCdkcUOO7Xt8pqpYgEHlIZLPQGWfxZ7a8JhgHxX
j5e9g3HfWSSquFoiny5bxnfNV2z+dFuS6Oje+oouxus/d8xN3e9RnhwgdNa5FYHgBTGyiZXv4Ktn
u2J0oCt2gTz5fAsrSHc3D04xRTMKY23xnY3/dkmx7fw5srKfdLoKKT8yU/l9NyZCVUfSdlYQyLXP
yLoXNtXkA1JAbbvFVH+DH1rJzZmLUF3ACcDs09F93AxveKhIZSPIDGJu+NLsU2v+W+5GhAxsPUTY
EAiMB2/Q173YBSDlrAYG4Ak72jZr1g4p1Xic+C5NGx9v92+peiRwjAGOxinh9J3MI9U0GVhLJ7Xd
CCkX2lct59EqyoZUQBwLGidycLDrIU++9UYXN9oSvHDnEQMTMstFjIHnBnsR8GZftw3Q0GjYQjNR
ktjNzBdZ0+lgAkpNLKeH+Ve0p26xWW9vTVcAlRP11390hXVyr5hfuGopFMT+RXfhAAYoinof90HN
Jst1tWpFdnNki1ABDHFz9Q/+LZtieIDU134EGSeEIeh5ha9Qlae3/9cI/6zqGyKHvj0UeXYmqL0n
rHLrfohSCY+M2s3WMkyj+wLSoYp1QN8JPz8P5fRTzZb8pfwg2DNk7v6bl4sVir6lG633YZbJJNud
wnLB5cn7cVYeYSAIijrLFx5ksVlebUMWOVkn/PykV+xScMIOZsXBP4/2AQbHAkG4NiSHvLltIN3g
F+MToyQTynxckRoKv2YNi3JngqbQieJzMHBRKCw7QHvX/tKJjHf1LzJgfr9XP24GhPMl1KUvZObX
du0/NeYl/rd6MXz3V/0mGkBg9+mfx/JBrQJJHcEtnWX4AKay2Hdebq6WSTnwfm7mXYatYm1kVgIa
1Qv2gbEBiMs6hoEfQpXv4H4IQxHqClXOLXUQh3d2PDBAREu9b3ciHZvk+gSg/gy39t/4kVIH4BGm
levYqufAziVaeaRZ8++bTMg/2A000PJLhmtUO6XBV9CYPFB5KRSFTO8uhj2+/f2Oitq4P9NedK0d
3ABmPyecXuAEqNqkFLLLkXZv2Aip1M22v2aONgE222whSpDfpMs628uTo66GaGTOK913tKSvfcdh
prSay/6Ut+dMcJSIKeLUA1x7fBHt+dSFuPmwwYNYFqUUVeDDvYyiZ2ps8OAo9PpdwAWZdndsom1T
Judi0VhQX2AWPhMKhSsgCNjLkS3ZIHHVh9/qJpWK3GLKFv+091rb6mTb/dnXieDoWEby/OKsphyz
l/1LgZAXD66aBNgB4bTIzLY9i6nk38cSp+s/AacZd/Ay7aRtT88xJe0ZSl6d4SH1ib8ZfmDA4Lx9
3xN9ZIsrBIDK+e+vXOSCZ0+rFpNXwhpwwH9bNtNIXsMFWKIdCAm0hQPT7WCaDH4f6+fBL90+qGeD
OGXFX4RFdp0q7hJ9iu3IGhND8gcz38fOOkT7Yrk++x0AUB+0Anj4qwA1CkA7Ux3hpwXBVLORyqtI
lOMV+GOtOT16rv/vqKDGKTAfNSz0sxOV3CwD7R0GAJ/nEuK7feeCGQ117jc+cQvaHMez/JsSYlv4
njTPFceWIeWKg8Wsil96knj3qJp6umbUxRaNLUelmYFnbrPINJbrGEsqwRcA4bnQbbxc5lnPq0lv
pzVBSUQX7PYtLhG7BiRymzLfq4GN7EoSDS9p7scbXOhe3Fe8OKiYw4ykkA8SqmR+/CYAcG0FZWQy
xa2lfqO+6Tn2tY4KThrcjLaF43hmPZatN9j7xEdmG8WwG1PcNtJU/fnDpMMKH/mYaLAJotZaQz9U
tk5d8o2dsDlwcFQ+cHwh40JhZ0KuBWnfbgu6anZ3vv3RzzWL6RQY9AwMDw5sZs/LKe1QbrgX/Awm
OeG+rHr0OXQvMSYymXxr/8Dzbn4oa4CwacxSX71QsZfF76cjh+J+k/Ylso4LHRF4I52KtYp9RDAx
mBPc4JB/ci0I5LyWoqsuB5GK2wPuykYG6zVshVkHpFtR5lke/aC8gTtveZJVq1/LxFnWITXUhYyT
HDyEUmV7QxpArnBEtZwhp6AVjpELUtgQfPhfSzwDI254LX0VVmzfd2Cw0AZrM8lBKA3gnmTGThSw
gP8HAIXrUNMBbNWpYXdzbVdjmxhQZ/+mJ4BlGDMbfXu8WHjaQFHvMo/YRirgnr4yeF8WMi3O2mvI
HlDuQIRS5N9F4XKFGLJjOp64GOcQgOTviUgNLCEDmuRpgQDz0RG12hN+DFhreEEMSanK0euzChbC
j67BbDydmV3HMPnEohemrOCsJgXYD0U8OLvDWcx5W+EZWR333/yiVCzx6VYLk2ipiyClu6mV7+ZO
9j30cMBKhi0Nvq8KR1rIBhN/Rg4S23vTc4Hf1vK5Fd4/05I/E8243LY1TBostS3lkwRbwaSY327j
DDniLI+XjFo+LKtepBJ2ST61cmcHAcXaYn2rswckeMTwmx83mARrCxV1HDIC/J6R+RIulOSedqQO
4Eo3aXLgmL0rhG/1odLvNFNlJyu/0Pulit5Qco5CgMUH3WhNx6Wrm9eyESaC2UKGEN8Bvkuw7mBZ
HLDYWD5PYDH3xCvXP0XMkev1Oi8napgnFEQdAfuFJkMn6WGCfla7KsI81sBsh5Viww6luOvMFOCv
n2J0sRBpjjDW7rCukvhTL1HfNcLVQC/roIcTxp/gSKUbns/FirhquxhVPKU7qNh1ty8JBH0Ng8pI
O/kMuLsG+iEJxLBlvAwB74FtdynGIEHal3hUtt08SSK97VVEMWEgiuXpXGC3T73y2zRiELAaD6Kp
opeYya53F8vBKICNjJ8beSkl76W149aqKDFfphNcNjsKZqIcO2ZMTOD0FnKCdy5PD/N5kdAJVaXS
9pg+0YwPgdiJiogq+OVxJ8zrC4TG0nOwcrUwa+c2cO6X9QSGvweWuxXZLYXiwweV6/hO/13OLyt1
a5R21ue7XMmZJhLnDpsNmWJWWBeZ3uv5bl8bEkg5IuujpRQr+oUde9Ss9H+KFMp5ensjNsxVAzfb
deKlN3z78wi5oDb6boZzEjfbCukwPBRAl1OHF3zJY4/THSo2FuSl6QVWbqATjCNMtyyKzZYuccGA
TxfSJFh9gZ3x8Hme5ccpja2osW165QO8omxOL1Dmd3DYV2O8Iqr2CSzXnybjoVfg3vNnDVkzv4OI
lZ15wpwT7ksXHu3vEm/OKLE01eHgHqra4f+EQ8R/5jGrQx1kmgDey9pliz8PuXPb3GyozE86a0r3
bRTOlTsf9iUbnWqMAmAllhPwt9EILWTpMp6BaB9WL1XMRD4o9eRE0dg2sT9RRdYC10emBIKBpcNs
WfeWsAijyA83hLlGPS6JXL/cuVsReIJK1lYNnCKNuxkzxpzk2DuhEX7hXjkaUcCjoyW953exMckW
vFExg4TF1ofzKF9IA3MeCEvLfAhb6jsBoci7m4c6VQL8BIsj/dZfx+sTui75Ls4tANS03A4PLkPt
nzkLArK+dUHMd9EVJd0hryzwY6RDzHuVUgNsAs5LSw9EvXEnUq8lG5fktsiWbTVj0vhx1nUx64H+
u2x//IuzbMVOP0C72iKH2zh+HOZWeADHjcV+V/+KYdyEpwd139iO6RogGBrbiUEvcmwVFRJynBAf
EMmDhR7B+7YaEiGsRsYWttdwrrbO8mYHilR/KLBDssO3pVnF4QtEPwA9BfJfcWhwn61fSluIPcvi
y++Wbjv/rPtE3mBbIpVGQnzxeFznFYM6Gl6IBx77WMA9uVH6TB3Hof28d7GNcC7dhY/wCKNVHkqx
Kg+sCRNSIW/mzvqz9rIvo9snINt+0wC1JEzmrrCDwnoJYjMKgil3hlmrvuHh0WesejJe9KrJ5djJ
i5QEZLl8MS9l5G/Q/9uoZmH1x44onOstOMGTT2IJJzBeIyUQwExcf/DHqi2Qg0aYjjwJxzypUZVa
Gf3d+fqZwUwPCiw0AGdSGFrYEoQ1KP7q5zS1VC/pwsEUHnd9pQFInRR06nfyddgFuaqRsy949EcT
P2bUperJ62Js1RR5L3jMXhtQQGXtppJIUHxN3kdT+clSZm3WF68phdIyepJjP9mQRA6//FwNMQH3
CDfIDn/Qnh3gA6t5w2lwZWdDub2VJaDD0z0ATmFfm56RLU1qyqUzEsM2sVT62/qZNDzxjD5KoXxV
bnsaUkSBA29w/Cm/DpeAW26YtCT74ECULjPMB7aCG0O9ieJaZSTUv+Fv+YKYChHes+UuZQ+el0U2
LFU//3OB5+aU+7MheQODQfKYH6qhTdqp+WIU3NYeEbG5jjzOP3VQfaxgiNpIUUQdTfskAU9oL06P
Dmz7wwj/Jm3m7VOUnjko/ZQSv+QLqKe6g9Nbx4PcJzdPzeuPXwqibSqmEYgeFNmD75SuGus2HLd7
0xH5ggI8zLJ0xtejDwryUf0WVfyPGBkSX2RL4fFvhQKlnd4IA/JLLC3HqqTfg+g80Q3MNL6IjAgf
aXalLMBQc2HPw27EniohhEhxPjPDDQnia9D1Q6Rf3NPZIsdFo+8saq8/9armsQdO8Ulhw9u+DNly
G8h+N5lKmmD+Rw/8/pfeSBPZ8TENT33ql655StqBoT6sParujNt3wimlfDzA2ZK0oeN8xd0U5tyG
MdQvSTtNZN490RUhiwcqSeGVCqfuHxG8a7wDU+M/pFoaEUdG2G25VQ5n5nJiXYPzXX+i+4bVGWd0
vhHE43PZA1DZvzTQs/ArtBxtfD6+6TNUueQ12sliTNNQeZFTZ+XfvR1bem4rWdzlc+grbXsB976X
s5rph2z/OXXD6I+Vw4Xu8TcgWhFq3dD1YBxSRwoWXJx5GL12x4l+dFduQAN5NxfDperF1FCVVYYL
6qJjRNCg+iUqTh88oyB1kqNRHPKYlcAWQvUJqMNZ5BkCZDGthNfYFfDYZtnH743+0gv2Nm/a+xV7
UMTb8mEEmMfrabmqDpLH3JVN77zb7uBB6rPoDTOlVVlASkaoz0NlPrl5iMG8rd5hE+SeZ/k0seLa
c2WM3zxXboch+nR9eAaD6M23zL5Na8FVePZW0YMkYA6iq1VjcURNdMlnjv2/yeLxmaJIFWK0PQCB
vGwBE1rDf/ofAsTBsU96VRGY/4U9CTeF2rAQzDTgFOHU4o7NWTbOyA2tfw1kE7PqSjZO1zl2TX7i
CBFxk5keJlsFZ+d91SgkbzxfFdz+1SoviR14Kv+gAC3raL5cv7AaB4HHFHHgySITqY+gdDfOtLlQ
SgQzsB55heG0ATaIiAUZA40nynNUhQ+lb3pOucDW/7HjyaT37CA0TRrs+fk6017c56neZPX6MYTb
whT8LfP9H1doRR9fDTrCAtSErhNHLlHc1+AKE2X3AClgAehFRrt2GARCeAUjSJKOHvhgfmGS6JjS
7SbNd12jmqXhsHbPl6+yEh8ldCWbN/Danj292OaG42CtJsEf7fduRhfrawQf57Edj2DBDECnmJ5p
DOGC2kyRrpOJ85UYOtr04poLLB9fVk7c3jWEuUCrhtU2J2kPkInkJ5NLfLtBHf1z5YD8xPvznUNb
HzObHUZ0025TklVWdmMS5cIXt5THOScNQpgWKI2xnd+M4VKFUP+n2zBatIsI1zEtaGW4j0oMSMW/
mTml+AOiNttyzy+xqAkIWJK4DAzvGFe/e2I5bKiV4hyPMPlXZBn5VgMeEsVeDU6KsbQ0obE/EUTT
JrzpKT2xJ2luAZltpXLLgkZ03pF67izBUp0fMSdYgeVaWc8CSOwl2Ee00LPK5IiLtaerQGx8lwsw
fVgbmwSv1dc8VRCJ2la8HaBq5o0th3k74gDuYUfub+nQ1PX/fPKvNBrVvaUOnF/4tOTZSmZuhGYF
Q7yAapdIE7zuHMp5ihzshP7PG708658X0H6kVkiZO2CCEfKqiI7Rr7sIezYU7j3VQyrDLhrjeHWG
HbwFqUHI4/DxZ44WwWXD+YmnvUnZ7qKfcocl9MAJmSQyguVYkwO44j/xRp2ACPPtjAprbELSZR4h
gHNoy1l5foNTkI42/667myHCzMWPfzJiu9nZrdvSIzi8w4N0MD4SrS+dScdduko3GT4TtaEmV71J
Qa/mGLkUyvp0TD8CH7m1LYE2iWVqqS72vy3DyPMGrhN/crMYW7FioOyQ20IEvAoYZiiwgqP7AJZs
GRQru+OYuc7ejV/pAh92mMdsZ1rQ40PWxFKAeEiyFalW89skAUgPlBqZyBTsGsPX06JiTLwltx9U
HavJBN3y9lpcDdAQR4zYiZ1xY4MgG6LNtFyQVDVvpQ2rsXaW1MIjCmCyOYJ3hGe8BDrygd96ABtm
QKpucmxwWlO47rzD+WqCFRwo2seuc797Z2UWfDVvQQGJrk6ABUBygRayieu9fJPDOStnwK9hi88u
gYjn+hRWd//4+DaYsp1XhsZO/9olHq81kKsVYsUQY9f3Q+8otQs5fPA7dEymm+gfYDbVQIBdwcFa
mUSep7gPMouPG7iVGnxIdcYG2k5U2VN1M07rNB5La+kg2nN7z+HgIuVIUTKquhjHS9K86MqAu+pQ
n4JR/UtUqbKGxP3kfrpQ0qKWTMuTRP7IfbgNURDrUlrO+H7W682M6/gPdsE0oisGEd0S3oisCYug
pgk+daLjjCefYtPDU3p9h3GYQl/s1BUsd8W7gHQYV4of4gNxvWVvXYJs6hfePMMuSNO/j/GiYfOP
BXL4cqTeBtloOGAR4ms8Npte1Jxls+9qEyiV1PjNKuv94CL2YRwuUSOkjQDeRtHnEaMR7FQexnXK
M+k2Maee3u3iCIDWbM6Kn11fW9YKqRuk/WuC/ZvFTo97re3MeJnWPJugg6ZW4KXHO6IwxCscfWmW
8hVW9LBJUWKymqMaZ55u8k55j1U8KDJYX2gDrD/SaigpLOLQdLzOIMN/5gb5ln9lxzAJOjqkQ4s1
aGJVjuEiSH8a5b04JelLdgTEy5cMtheUdLFG6Hq3TitcKKvhBKVPYSogUPNWOslKvSjYdvW37p43
n9bUUETA8JALIV3DNbRvdlF2gHI4hG5eW9iDc4cCQJHt+yK4PgegTfSVkcHoTn1yCGl+UWd2LADL
ot09hG0O+gz04wtq5fjR3I7vEAddKyb+4Zxz4RD2XEyw5KRTjpf3VEp6o3DVJBCccc83ESxoSgzp
aUumynmiDq6anc86CW/wgyOCK1m0WiY4CX0ATgTVg/Kt/OM2vhrPHEgzXx4jIyt7lU+cvcswxfm1
Y6+Yr386kYdWV0GVSkRpxvF9Is12cb7YboNqW9upR7AK/pSx1Cl668TUQsusWmp90pfXeN+UlUS9
Ro/FfYzcecuTu6iJ0Njs86p2RJLUFc1hwfgQaOipMkQUG82Z2qb9jTyXBojUfeEvcJnvYzaw9IGr
CprnYJo3z3/Y38dLUdvabEFke2f+caYR5yhXH1GXwBp06/MU0If8rnFCliLc6JQ2uh6sBNJxMR6d
mVjW9UOUp+h5WHK4yNqJnePXtWRvbDpuYELNTlhBU/3D14R2851f5dsffQttl/TeikLTTzCBCkuD
66tr9/8Uy3u4gp0d70Hwefjdjw1Nc4iJ13EIafWN1C3jfKWVGLlZZylDVgt1QxR5n15pHeDLQrhj
G330LZekA4NETvsyrDF6US1FoT/so8uLLZL64WJD95KQ34zPcDJRazPUV+y0a1nYdymPsnjwOno+
3JuTuKWaUDPxLsv8cAYrkWMSkdxq50pXCQrj9MF1dJysDT4La8OOfzJEsUgK+SNHb/0COfiiARGm
PR/3uukJHdN9sMfs/9ZF2IYDq+JVXNJqYtz0vTngAhhrRdSd3OAgAT8wEZoWcxo0L1kZrDLGil3Y
wg+1T/OqMMZNhywn5m6znvD3ft44NYxD0N4lLxO1SFjI7Ps+P1Eygd+Mi5NbgBkhWQg7M/dCCrxS
mAEmE4W9VF32tQgto3WV8+7pbU6htsTsrbkLkyPJYPLwtecFQP2iIpgLST9Fjnlnlf6F4jnSDFrz
p9tgIspLDJ595RB24u/Pp3LcWm37yca5cUFKMy6zE6oM8oZfCAg4mhGIpuO3Lja3aA4wY4Y0YKQe
aq6GVtK0H65rTkk9R0/0rXZkI90C0hvMeY9F36+2D8vRagv9Sgob7aVO6XqEzS2/WeZ7+cKwMHTc
WLHweiGqHuD5OhUbctxMvWToXQTr4e2Iqo8O1p5b2GoEtMBu7CHE+3SPLXNm6sDcUcLgC5snOeSa
kWm2DZE+3fpxon4dx3s4L1ww/fTfozdAhwSQgup0HwN6xIBt7DNXz26ZnRGR2T2QlEm73CJ+c5D8
2rTZN6YPlZDKBBoeKqlO5xFcGgR5VfCuEZ2KC5JpTYlRmd37/xQb8az0kGlJrMf4QUao2SJg8XS8
MiO91IisYbLaL+ogsuOMDbDWpiw0SDwOXMua/lWu7DwIvOXkZBHve20XVqtX5MJ0zkr3yNFi8C29
jdj8jU35qksbcShZpKrc1K7yyOccyfmyu3ZDqr46+U3yeXG/tTgmVT2++2Hw5UJF/3s+MSKzshr/
ITiQt/UzYywtb3w3zIuscFWVu2AdG4Oa+X9o/wB2Jwgt+E71zFXO0V+aUXrTA0NITdvHIj1V8wy3
u0EA7rZL2uR7Sph7V8HqWFf6GodZQhw87SQ4fni+5zVs6mX2XMvP2g7a+gQPlUIwovdo35T+DkVq
gfZFnDx9qLbAF0pWtEc4Sv1xxdUwJhht+UFgv4VP9LyOAxnpBQ85rtQeoz64ire/8jdKpyqBvLms
DaLcvDlN57VHjUUiHS6C2sJkBZxwQ48ru3FJQ3hgFDVfwZ8xte5MCPOwocM+P81/18BWuBqhEazB
B4F2ZOhDtChgDsElbnCEeEvbwOQwQVHPBNI0UZPAtXco5Y2mejUbM5sRdovtJSTch1BD40cIHPpO
MnmRwf4R2RMR7tloABDyn5UPEoL2B0+XdHN1Ma8d7qnLrkCj5SRrnkLKqPQx1QN2B1inBdFXnKRW
x6VvDi/sMs6uCDUGwEm0sAaAPKz3XUhU0HMUFQd27k8ZjxIiF8kLmAMqb+G1uRMHTajPVrkYiwwh
Fl1681e3biVhb07qhZFrBXxs4stf6qQQXWXJDz6QrRRcQmC/50b8LKjc8gXWk7D7VI5OyVaVBRpR
MwtumysrHKuN28tZlC8G/HZQsJjNyx4NAkD+nh0wLeAj4IBIxlR1igPmbeGx5UgYte+igBOe9Awq
7d1D9ecmtwNV4uctCMQIEyIlfnhhleWuYaJquKpVJVv9uJOfgphHvlrwvVLVCqhCR0eeABbi1CFP
2LDrz9Jxd+VNtkhAs9H3apZUZ0ItlQGKus4QHsU2wXNAqoKPHf1K6SsNbElPUtJsHGj7I1FFIAOW
TBKuKIPuyC32ZW2l4NGhOI4j0+gLy6CBfH84z2bk8QtAjLxwYVCclcZh15NpHOwcC9IhIT8HJ0Cj
DeA0KlmnzNz/Mrg9pggWvl6/smTrSOkaD0EUrKVU38cWOAnLUYmSMSkvKJmH5y+K5SJzTWEryOVG
2fQ7aARp6gDyAhtS3PMkycPOWe02sRt9/zf6eTG+J+Vbkq7ZSlOCEbJkr+a9pYHA+7v7xRiYVPnW
IIckSevuLt1Dr93yLU8/f1LXWB7RUAqEy9EezHj69c52pmKN+r/izriTLzx48pbzorEZj6LYO6Va
B3v8xFsJ1ySme/p1ac9w2NQKnGQjEnmMmNAUY2yRrRsUNliF7yYrFw4NsDS4wHRkV8omoM8eSGmf
UnbJoXda0Y4hqtwhJzJBmu6n79tLmhVnFCansz/R6++QsA5jQgh2ChgwFHfzIxluUArum9VIU+tC
8wIHl6xlQG3ulKkR8qYcMmajLn6GdZ0qDYE8BJeulghKhS/X5GtWIvME3mFMlg69w3/Ilbi+PKDs
VXefhf7iq1sOyPUFozRtXPsGkWPgIdnhuMf6rMZFJIPB5L3eIB7UufKryZP9pStXEbfHRdByCtNK
h2yMWsSicgWoeRvUjafF/5PK/eeN033ReLhrqyBayTK6SLTtfWNER1PZEOYeNu2Dtu3aF76NfHyc
qj5q2fw/YRsehfAjDLDd4qEY1qbLxb8xav87NfbGHSVFozlDJQd/GAVaiMdBw+sAlOmjLoAkUXsG
j7iravNU6wJ+NTUnsTx1CK59UxO6QUR7By8POp2ftvOkGIQBfZTJFe3d3mOt3sOYJfH0Q4PKu2FV
gGwn02WoI/m/Hen1gZ47ZLF+WJ/8BXCY6sBCecdA61dxEOi92kn1e99xx4rfu+JwWIK1jsL9C3/r
RVEMo/X+TnB3hdesX57p0Uc0xlkzcKmWSjYkZu6AnK+RoLhhdxWndZJ6PYerhdRrNn6w+eHuHfYo
XUS9ETCe8Rse8WLu4lvTyhoUvSUZpJHenwr9+zGzD+P6B4WEOUX2esQVr4NfVo0HOuIv7XYf+qA+
e54b1lhtShknug/AKlocWxHeEF7ugkHbfsYBMyMCtlaPrgK8VjZKtkfFV5vAKu6/9p0wMio0A5BZ
OCwmbfeaataFyRZDIVGdl/OOZtbil46qujP5cUikXI+2rb9yAZXdNRqNPyJEQE2lNjGaqovKnovl
vN6SqVMmo1pda/vjKZy0by4X41HHFLyfsvFX4c8KlVCqri9tyC+hFIggCfRVAXzq96jMiGxgxIfM
gO7A6s7Thv3zjdfcZY+onmf1fPtyN8OJPfPYtFmu+C5wUUgttde9io3SOx5HRBLd4V8TKivMgHJR
Qs9MOWcBnqM60U3TlYlD/1nT4L0/ZfGscelCpIUSK6fJggEeDVA7V9xSIKHEy/sGPiVjxr+HjPGT
svO5urD4kMYk8tYhGB6+v/mprchsBs1z6lggaK8pFGysrZGYw1yrWjInAlY09d4Ce6eVPWDH3Use
dtMKwzy3OjkUwlyVr5w5cmuczrEipHApitC9CGeHLd6S5GFykDGdpeVjrEieFpJREItar3L/H3Vr
1YbgVjowPBVMf3LXIA5G15Qz79ow8KFlhsK5AJIUSq+oKMFXuVuBkaEAJPWwu67O6tfjXFwJ0ZPT
6B7z5Nujx0QBIkMqGHaO1rhcQrPmfFgDQozcMsWyB9tHzUOVSsnu9emr3QfaxUlg4avjRX4xmJ1h
s7nZ5VlURBf4PZ6yt4wcwBmppNOvgANAn/T7azG68eAghLSbMYiCWK/ZpjkI3aK4CFfBKPXYG3Yn
x1MR+QMOs0jvD8/ZoiWe/lpspDY3FG3UBdg+hsWCArpzQPNrbHBW/FvpMN0nYx54CWfBCu+7uz0q
DWwmo0NPXrDHN9ykmcLBDVVSAJcfZW8UFZh4jrRKG9qiu97VwTmKSOf57kGyDEJmtiNxV7oqGuOt
7a8gDEC0MJCkJsGIL7ESUninRAW7aFYtekNnkZJHd2SEAqyWat4ZtVMWNFDo4jA8pKqeFzlTD0kM
0xrgByvHi2/ZTGd4hxKi+rCIdc4uif4rgiI+Bmz/a5NVKRobMdvLJmCXWIt0Tsx/5O0Agir6qQGk
sEeJoYRROLh1AAcEJMj/I0+z3sfgZxp6B2bURUuniQIeQ7L+AjUwOHTtTlU7Ixkhqgcxyr7Z3gg/
RV5/8L9ZhRQVhoCqhqaY4ppQ93Idorcsj3/EaYIu2L/73lK+IBSS2+IGr65cvBOOzheQEj2PX/iU
9irBK3uQjRkS5Rpnp7cteothkajsLqO+GsZ0uzZ9NdLfdX7TZKCI308jb1CWJsl7aIvHO2qyTsCN
8umGpkVcyRrQHZ231GuhfkRFlVd2w/AtnaJ6nTttr8UGgCgEx+1rx0QIhYNBNlpBnB71vThLJK5Z
24pExW5s4d0So8n+/WcYDGD4UnhQ/Z2UyKuhpXhnIZqExmkv0rNnmR4fn0EiW+vklWytQGuQ4tuj
QYLuFd0dhTWMyFPKLSPR1DXwJacIxW2izUzaZYBfEik459lXEtyeKxoEpyWDa+gW0zDtaQR5r0o2
/lnX2R6+IeSrFVuchSw8zAr/zFGoC1RjSVgX0R2xw8Fl3onw6BGGgiOhG+ApRr2ZJ2N04eWOPkzk
OUocO3ZgNmgjrPP1D73+5jtja3LIX4RrjXMdx74uQPAT4XQ+HK7E0QL6L9qGt/36FYtqhuIhdQ0X
awQgV0msreUZEoRU6j8PWIcVr7tskehr4WrYhCLB4UWLFZgWoVe3SqeJMJidnvEiZKxWQu1fOzBL
vLGNMHbBQwTDTJIZRQAJ0eqrKxQChUOC0lfDqQcWhhRH3rN2ybrJq4bHqUhQXBHHu4oooc8tG4i7
J+IrKICjm5w3AGRViVljXtDLnNzf2EQ1XQpA/UzD0/2AcPJetBKdD+HM1LW/qHpopkPfmeaj0g2F
WTbken6FwQa29GzR9HjZw8zh9SO4/lkZGn970MXxpj9SZsC8pf/2TsNR6a3xKHbsZodLT0bXA8F7
FAwp2tCnXCIB1L9Z5lXcblKdag2C+AGAVgr0V+ukzViS4w7n07qnjdPjHXTTYPnlWeC6wD+xIVu8
M8EdlDCgaLMOKDX2HzNChD6beVXh+3R4sKHloyw4G247x2Rp7+NAPdo2eEcviUlq3/mF1vMEUoBd
AmKofuMDU8TYKdZFqmaSGBNSL32nQoRK1iJfflCKfw/fSrYIpEm2ManrVYkkWU8jsKeDH2xfHya/
fOyvPHW40t1sv8KdV5ZSylMvEQprvoCImT2SdrdthSEO1yA2JLl8r/Ab+FDMgyidre3p7Q3GWDHK
x3bP6gOTj/KPUxY01QyP+8dQjBc/nSs4lWzDXlOE5PrmsSXGmg/zuTOrGPJf4iyi+suBhwTEzD7h
6/EC8W2jYU9xgOKNK9MT9tcxm8ZXDO5/FKjhWcFwF+o5h+svAearUSGxT41CibQbVGlyeL3saj8s
2t1SV12y/S05upBs7STZYEEQVNQ4nEbvm05ADDYRplRdLvoJ6LyTsXfXfFnBD3CM7ZrL3GN498V/
gn9WPkPTlap2IwonjwT0+nVZlSPB0glFEAgXpe4MXPdEVQhhq3tEXCVgailgsxQmVF+QCLS5yYna
4t84kg8TrsdLT/yoLZ//rrwviC/N+udSa/N1Zhts1EuNDpOnDdNfAiC6ygigTiW01kSVI7zD8nwv
EReu4Z8wg82RDjSNmodvSkuRWc3oH9mt5+1LmMYFQSc9e1HYjVlOXBgwQ3iS488L0tgr+18KaSF/
x7TerbxyQ88sVNkx1SeRcIjrFxGnzu6iC992pDWJDSQjpOfzX5q3p43DCBsU9ydpKFWE1BxJTUH9
b2A0hvF1jePMsPtk3XMnhV0lIg0j5OQ7imbDGwHdmfLVqngag96DIRhhyTwtPqnX1MC9syGa61vP
0gQFM7PP5J/4nUNeBogLbFWt/txwKs0FxuTLGNKyBNZi97AHWq1uEh+mtFFd7Kk2xOFYqd0bUI7m
OZT8TG6rRxGn+QLnoqLhs3+10eoPLSSasGzK75shRp0CVxakN6dZyg43HkZ6Lkm10hoKn8R/vZhD
rMcy4VBkmkLPMyftXIntxnPiwHwak97S7PtreG8isLe7FxdNScF6P5wp3SCgldMLq/HZ3kAMAp4o
iB9ObLLDLDs/47m47flrvsMtoM87dGgZM9cXdWEKRwVIm9lYh+x+kZkr2FJ8pVwLle4Az6lI9MP1
GVaj81GUs3jN04hF//1Vx0V39vkrdQBb66efcUEHlOVQqfj976U90nRvyHFvKoEDBVcoKFMQV3q5
scoUYc7BWfzPT9LvZjCyno0X+FvFGV0cDRNgTlg3mstYaMuSDlJ++iN6SESmpHNmc9DkhImfto3f
ROcIkHjcQ87t1enfli+/6QJxtJbE5Hqv39/buIRIWVSGQ481ICelXbATWVpYAnH51S35CMPYOiD0
/EeylgtkR4KniTWo6VNPGggUBWlG9I2svySi9lZCrrH+RNywZbHMttenQ2RwUa+ZHL3AYT7dHLYQ
94zvL5IZ9lOMrZcd23HZIqcCVHtYPwou7tPjPKuLCVB/3NXqimB19brJxFoxDM8jJkjZB89fjxI8
FTfo21Oa7c7DgAMO6l9WZhKMqAf8LDrXu6L2oZHVkGncgVQ/ItLyex5ZCMBRN/bc17nAojYW3/Sz
bEPKNOfmXP40ScJx9jQIYsKgXOqS8t89YiFGFNKlN+C4AFjPAekjthumvT5fTKohmlNIm/UDWExK
dYYjjPpJtyA4HoclQRCODYVEy0Qa85rFwTSJZgYAITXdKFKWqGLEA5kNWBtYgKqZ6ANWhaIDEkXH
7KheVBZpjvzTyM2Thgp4BQxsGnZQSYkskG/0Bg7MGpqoGP9KzW/Sio37Ibz6K5YHoeQ/zJbYv+aA
kIg8Z6rltZh219VuEsC4+t8MjdIaNsIl6iz/cV3k5S7LS+KKW+SWcqgwn2/3cuxhadXwmOuZizs8
+ODxmhsyBzcnYkP5DAYfR4omjbNkmdvlgfRgxCJVA6zVIgTCTqzIxrpnYHpx40kVbwdPpK8D8Y6g
EvcuIPqQ76HnY+rrvehgdRMHpfUwepyEroOvkWV7YL6vot1htI0LT3sRR7g61FgtNg5yNhgPpxcH
qVpvjYuHqsV5cgPPelH3xCkGXgbCLDRyk7P/chB9PM2UPH5yHcsO6NcGmaH9X3H1UhdynX57Z5ak
Wo4l/Yq0Tckk9NR1Zls01okaioOWvAYe2kTrjYDnqlfglQQBb5F8m/I+ZD7b3N+n8fsypFm9WTFc
OB4nK/yqZrdlIaqDjJaxdUBT9Lu/SlSxGlEtFlyeaxj8xWMDuVZnpT6fIFXZFW7ncYMwvTvIFBsz
Si7Soy53peRHemDenile6NiU8xarAOfii9W5LPclGn+zBUaot3N2ww49qF0r4Whwl+y04F5zQLMH
nS0JJILBhq2Zp0ednC36RIBNOjPiVPqXUV7wv9ljzGjebJgXpKHB6189DGKRwiU4joiI6Zt7QEJU
8+qQDSdGBahobyIjmF/nsUNLpRPkwXndmVJis9TNqKNFSVuLoUsj71bB2VQ5mne7UX4dbeQBvD9O
956BjS9GzOiOgHcnim+hi3GTdPLopCoKytA7Q/Wo68Jw6ZHr7XfvyhM9EvE5wYdnqs2AIgE85k0t
I6JpR/QvzQTHWoytQqob6jBJ+6Wl5Jty7sAL7DUUGNiZm2T/FFcUkuwqDaIyDb9epxBNA/8Ot6IL
3o12W0g8/1C536D1nJyy7E3xFZPFlP4s4rYZJ2zGcLex6AEg4rC3MmTYOfTtIufYCDjv2uRCkN4A
OITD0vDqjZtXMtn8XUnqSKR+UaK/WEpqu/m5teZeFCcRi+r7DhjMTpVth4rQpa229EigatjxyZ8c
ADwC3/dEVjRYrpY3q7TYE17FIZvlBhi84MuVLPCs2qlI0Zx898+2pyIbe5aVGQJea5jg5Rufgxqo
X1ycdZsHxHJrhQDosZhzwnL/FojdlJZzYMiccjz759fIUHdSGyKkilxbSXezqGb4PEb+48392oL0
yYmtlORptcRo+udXc7cwAeXDh5Fc7XgiDLx3CD7Z2A36QoWygIudxC0FjhKpW6n1MfpgCodlE44M
VQGI3JoIyLDN7Q5xluGFwOdzK5akF5DHiGvBOsxJRt5Bi4tHcR0tV1/+Wp/3y1uhvkj0xizSqydt
IpWAhDkIBINJkIOezqNoygG+ySpjz6jfGhTOKkKb4CPXLs1xv0Iu3n/qx4Zm56/jIs6vPKAZ/lu9
W8rxjm7gO7nsg4T0pEsChHVK4B1/2N9vSmnfH6dtCd+ayDdZVQZANfaAUFGOu7nt+K6n7SLk/1x2
u2n5wmwcQiWni/xz3Hmnk5rRE97aHZrEHkvt5L5UpcJZ4NYAM7gJQ/8nh+EPhrBxE8HYe2zCYIQ9
umJZwBNUyp38AZHoTcFGiQ0kd2rUK7+JaGAapyYQkvWdjmSl5COl/RuMH305OlCsw27mFsMwyxFn
POFMBmbkf0wDKreGxEMt6BV7gdGS895p8OM7wr04JjQrNYEUCBlQvyL0dyTOW6Ht1PeP+WkHv2eQ
jyfeWmEB+vHo1Oo3mKXmCQYBp8W4SlGYQjzKxC0Rqxn7To7V5XS/r7eB/r6un+UoNzlXATnCZQyA
Fn9mTC8R7Y5lG9fN70Xw/eA4sO0DGvvFvJf0ZGfHEvMd58bt2acjutySXx2uyuaxteSA/gMvpkxo
GwOT+MEuB1yUiSfY3lIXUpLrRC1vVnzNdye8DngO0VRgmk2H5cau2EilqDQJtgAl5kqeZhtAp7Ha
tbZNMmJPx6T39YeUR6scjIg1b+0W8aUpDlRd+eSLgNMW28rxzlDluM3YKxO+fLvpvp96DQzeQ/lh
CzfRzuicbEZX5hmy1dqI8b4itWJKZ8BCWnY0fJGs2Wtk6MXK7G0cWA9OXBPFc/TLjlmIAp+9gNcp
Dav3FKISoSKZ9+BZBLDIHtiAlregy9lCSqP6RoRLeD3+MCtKi4jdUivV+Ozlj8DvLfoDD+lbuHPz
HFIN6+EYNDmBow6Nvm1b43WHeRuDpMpYWRObiz7231FRH6IOTkvYwiyKyWiwhuBzLfpWU6753WoP
Yvmrp8UL2uZFUUXB6jMj8AlxXJlAELp54sX58FGhcIfJFNyJHeiWGNvw/CHdTwDeQ6rrnBiVF/1j
vOX3gX4M/AcM4z0qtxrv9cr3bFeRasX0PR8s8d7GzqF37x486ip/MBd7xFZdGz+3cZa9IviJCP/n
trh8Hc4mxon6wcZLj+D6J5Wnk250H7PxtjP5dLDs/e32E73pLj4pgZdb9hgJfavw9/UNZbEUsIkh
IA5t/KEUIyXhy0y12B//PAy6robtBgLBdhITKwzDgRUHZI/A9yjXtj3B7mJbFDuJ9viZ0oDBUhqX
BeI5sZ7rnOCDfYet8hX2zgMGZ00lVhC4F8A896NcT6BGYRSPzfD5KfsJ1T4vX8D8NLCV1V2tN17E
IhJPm2tNcP68R0zQeJxiN2JGN6Jw5Zwy8OPFPamWZgzuZOdDS0NNW86OnAroWwnHgNVYV7bsvTom
feCTAjyJc6Z/fwpWAMl7wdm2E4YwHsb7kW9HA3cunPrWbnpRGoZggAGFIC5vT9F3GnzsuE69GLTt
ufWs+ATwRldCi/115Fl1CeWEhF/i2zqY2eo0kpdm+501kQ6CO0ea5iwGyTWYkIjelYwzTKqrqKoL
JsHYSflwYPKpO4JSBzzAbk/qKBZWnLhpEmai3vhw6shql0BskTk8+kDM7NKBJ+PFKbKaBwoHKtmy
UOwGYM0Vb26WfEDo7XMAno5Wlnw4mXPLM3kedxQkvySQLb0xVEHn+QIJNuqAFWzzJunxClDjOL8t
AFmpQUUW3jy8LjK/7UNy7AiK0AS598k73ssrAIqZh3W+NEkFHyydu6Ff1SdAYWd4BfILf87g4FF+
Al6glWt04ee8ImrcYn/UGZjrnHLaR31JNbvWQAlo0yZLjkyZeekRHzvXzFqGxtpBEVwj4Jyyt7L9
oSnNiaPmV9pbJrAq+dzDIgmef1nVnY4C4E1jEIKBKUdVwpijdM34sAdHsHsMUWm2KUsoVA4y8f45
Uhd66Ua+ZrcjbaZ8lGVQfE44mpXSEM4/pQoX4wOXGusnrxhYaJr4p+e2Fgs8nmOjrBKZuvbGeFmm
5bykP0M9Qrt7j/mJBvERvIUGz/BwKv3D/azZ8B9aL3a48ZkJlULOzd3+Q7vYeUYyAOqGvDgKOHu1
zjbyPZE3s1aapqncjvk+lPJF0KR8+OLAsdewdDNTV+YseJKV37ZYwYeE0fV89rhXUKimaI4tXlft
aBWbCMON7lsoztrs7ty1HMB3biCjrf4G56gF0D13iwMYmcsqXkN2HHLMLdvIQPS+8mXMl0ueGhxw
sYckb9d/GoU+kn2eJJQJ8yu2FTY8fcGFH2g/TzYldao8L4v8jnVkhk0549taJulmrvHQkMShDSmP
OroQ40yhEnXoNpTxUSP3y1pcjl1gsnE0jymvReDB3Dm+oPl9uDhQ8FZQydYRkbIy6fPG1TRkkn1G
KEbaKQSM9E9Devia52eFapPl7BqxzFnJZ2QzmDPw4+aGlMAMcbB+CLqy5toVzbUEye+UliksJxYb
JWQRRxy63NJauKQYSwTQYtSvvKjbGRddUC6g/7PWG1VNVwL/45r8KWdStysP9S+c9c2zJ4OPUPO5
P8xpKf63JKrnLbJ41QwOP9C5n0+nbeba3UI/XPeWboeJceQ5wm8hYhU8trQwUNVeH6GvC4/zi1X+
o05zGIwSdg6lXCN/0xamszV3IZasQUvLmPwVUa1ON/8s/2/nDF5sSGJa+G7xBFqgYRpuKDo4lFp0
Q4LK43pAZJ8L5afTpWRp87xcYGM4YIiZB26AsysY2nionajOyzTeWFHvQbG2oknk8unf0eD+/aW5
bzcdmQYpA7ohUkVKNjSnKM1JxlyNdisc0gySfvJFOwwEqobcfMU/Xe2whtl2ZY7TqrUVEL4AoU+d
v9wQDGCZ2rZf49wgzOsGWPXHWXZEhUTo2DKdJeZy0aCL/R+fii6vVGGcheLoPzvYXY9rbAZVGTwQ
Y0AWrTbSw6jn02D/b9M3Pt4/Ci2YY3oLDmNaM/KtbQN1OGDPeBmBC8Tb/SmBp7UfpHzxPzAijCYs
5bdegvT90ICokLjw0c6kAMll3gGfpHJdhrzrWJPCOqhKUC2Fa+uY4V/npKXttAGdqASEywb/DMK9
QjxEOEfQs0XXRB/IXnCq3KTTLOqDoZdB3hgQxiQneT0quvURzahcL6vY3RO5o44sBr4jglG4o8oc
tUHDjImJn7FfAYWmrOjdDUXMk4FNpO28xavUeBT/m5Id7TYCgMrmuN07bFY4XTvfCEnOfn4oO9+m
3aqBpELIITIcdGAEBDny8M5uk+TIL0UgZu+CklCWqjVi6T1B4HTc7L5SJbvAESwfZCfkjjDcmROT
5yudST3kjEC4NnQNMnEAprYXGI91XNu49z2ryzjLSCLrHe/i8qdLw9KlWTYfJk83kY3o/np/L9NF
n0O8nYwhzLvcg74DT8oy+gskxkhhgie5GygeHjUHNBXMx83XMzAx5rXg76oHjEs2+iiMLfdO6GD+
1qfne+iEQDUuNm+o7jZwZyl1+4svrq1t5EvKxlvbgSotztBSK0xsX4+jm8IB9f0Opd++z7QYkr8I
9D5vjG5SdDRhutS4i8u8pzvQLRprIgk1cr30YKbXaGBocOQm64jf/77ieUBmsWSsPm1a48xUxetU
mINhysXaJiCdGxe6a6s5OO+YcbxPpS+RPdLNel9XysxMDEeqDMkwSM+NK4u54RFq08A04XXD6KaL
L6tWzFvFivKqD/vxP1oi0ldc2DWD9jGvFmqtofk298vkgUTQGp+XD3fhc6UW02cXu75Wfc/u4Xv3
krBaFwC2jqsquPzqvaM9vV5ZEkCxMnF6WnDCkwuY7QIhgwCuUEdhwSEXuXbloj6Q1xK60gpiEYPN
QITnKgkNMD8115AuLg0zbCSpZMcEF+TFZTvCRrd9jX8Ecp2G4RUkcfAhix6Jg6Oemp0IrHAapB6q
1XFy6zKpTKh4IS1BQcwbW4vpb8YfkPaSPKlJS4M9LcHVBZjvfNDEyGp+eMqiUk/cOWKAj9W2DEkL
7d4CP/ii2geW5VQzMccrSsiN4s5yNYmZBMDlXjmKpLL4QE5WFtLiXb57NylopFSYy2ITpBr+lXY0
YpTsX0uyDOilG1svFhxXHcE7U15gPF8vNi9DcAdAKSJVF+5pQrU3xWE0Iz9f+OE/Mnw2OYricHeR
po74wgUW0OX6y0zzE+gq1XbrkeRDCTZH+iUqeC0b171o7wdxeD0ohwm9TE/WnU26rOuWOeGd/SeT
Q0G7f9K8CZq6P1aYBZViFiBoE9c8cSuERUR/VtKQms8r+dHxQrzUebIDo9jA0JZjlMoeNc/LvnaF
paqzYf5s8nfrZLwvXB+axoxLNLHG+GGhDkF9ItWv43kQ2gkak7uLHmsojD9L/puOG2R5NJsAUvBS
Rjg1sFJZ2NpDKStmgftIhGsy4MXpX+fbYCy+t1uC5giEsSK8/YCQmBvEmnBsFyOBl7/zC3Dn4zQZ
+z2Mixc8nl4bUxVcK4TJLfFjK4vEg1eaMSE7DfQPXxF7hme1UEAmRm4G5nCSxZ3l5bTL3GNVTzPy
tdVECCR43YeDABpcmeJj/EzbvYGzG8hBjMvaWM2YGnDpZHHEKNZ48UcOudYtRJNI9wqz71oTEHBe
m/UD0Y5vxfHnPJK3TDhI/BHbaXu9jgAZEwUapnm/g1SfPAc1oOcKMToPS9GygyLZg0jjZzlh0yc5
h1Q2L1b6RoFEpNMgmygGOBLNp6jCh8/o9gGELy7Z2K0H5tQGu94rGcZl88K6e7fXn1Q/VwdtCcDE
ifrw25MoA7KsJcDJIJPhhKFVnNlvwPUFQW8GA4Kjed+9j3ar1qkg50dnVWvbsag8K3i/pjoZ8CVW
GNBfF1hi1/jYi3smrMy5qMwBWszBlNKFAtZruo37TXNrovWDorTPu6UOmU2EF0cO2KEFOh/T6J9T
q4OWoitM8AOhdNlH1CjPo3Kk99SURC7u8YUAu/q2lG6SgnaVGoU2b40e+hYQcIdRLNECYtva4ils
MtByzuUKl3gvSplQAGmxX5JmYhHseGhKPwmRogO/KRcde528Sd+55kPzC920paxbWUXmNwOmOfNd
AXvJWGwMROzh496qOEIGJ3iwJ5IqpjqqvV7wYrtbcETb6ZHA68SxZq56L/fNxeihl/Ri82zRpxx1
mXEhbpCqbec2rkuIpE8GiL/Cy/dz1XvRmUhpXKdYJJMJVGyuBOICqmrfe8Ww+VBI7c7+zHmoJj4t
wMc8k87mibFQBHUPeq0+jJkhSbhRgJDuu7n/tJCvahBbdyxB8Gz9EKX2hRLG+l/N8Gxc57A1adqG
IVRcavbxJk4iJpoKQAfMZKy4Nu7MU9gki8tkx8ocUEPDoXr/i5u+zfQkRx+hFQNmqvsOMVmVmFcp
x+2zpOsTAvXhly8uhyxtDVwSG2EU41DbJsEjL/eULUaWH8IPbemyx+q2f3byGjk9Nd6tbIYkDwZ7
HdcgvJTWvXWUu53f+wYAQNt0gDytzcxnuY0q+YKMSTRYY/g4ggUSdqeREp1VCLUzxQG6oLbb1H7I
g7Uty1zbt71S1aa25dxaYRKQ8+3wgocBvMZWQTdeHEo9wkfqEgj0EsROFDUeDLlBedOSI4uygs38
Xy6ainZHuCOfsgANqwAdH7vDBe9KTOwXesSa/bulXlKG3jHE30OBCx17pYH3inuH+ygeDriL7XHp
aDgDFEf7OyANsGo39eevCaHIJ+eairdC7YBSu2qBPyT2yRd4y94yen5Df0iuf0maZ9rnyxrvD+WR
azKdeiN4l6nKIGsCEPR4rR46d1rXCgc7S5OZedS55qRelTG+lfIOWd7548S6oAhpI6RHTDVQsye1
55IMCexY/Vy+z4Gsk03baeRplsC/+cAciFpNlXPQzDhnEkAE/5Ko8+ZtKitR/mDfPXIRFAyqlZG8
YC6Aj+FA971XFChtm5ZUGMj5ALSYhQVCTLJf8vGSceGaRsndJifcU72C6a9Z0V4CkpHAL6tQEm0a
NwtMOrLssbUDidO8kQkK4mRWhLIknQsNtjSl0ap/7Jpb2mfL3klr9jTqyzTNLP2wMKfrHgsul+AC
a+SlSdsK9Ryka7r9gK5tRKMYyBXwzG23p1Iv8taxXi98h1bXomCCd6GyItgjIKpY83QMkUTeDwS0
ue8fgsbCn1dAS3ZJ4mwa0wMSyDzeVOucdYO41+DKXwLYflqoMTtYOFDUzbQbynULkn0f28bEb7lz
FZCA/XuWd52H7I5Hve2vSCFm+RMzyXW4KVHwp36u4rtym8k9gi0LwA3CEYuM88gFk1Gf0l/Gysl1
WUES60XC2PGX8vpfc8fZcK2WZ6kbiRj/M1ANHTu9tVjwfvGK6oMGLvRlOvLO08/etPKnj4aEAbLO
A668bArY5Egf60bIaMHpio9OZupJjKnnhamHyukTudsYID+jdDygSSg08WjPGAYqJtCfvaKjvV15
31Vdij7S2HNCF0siEpOgePsHtRMHGoXnqdVOZxCukX03cmMUxp0v7ppukhYdZuR6LYBwxcJsl4Q/
pZBXcJPvrDbryPDIdQt9twYtqHx76JzbY63y4EAoCSJ+6WndfThMwX7h5rSFqInD6F3UsZ/THYQY
qfRkmfGI5fVafYzTGci3p8BTlgzLJr6YF5/L14SuMGDDhualVBGTX8uwvcmsgfcPp8l1tI/d14EK
hyhot4MZxj03s63NEx7NQyrAHO/RQ4b8sVIte8epre/FbG4rMDpxfHPZxZW5uQXFDyoQDwJ7PL36
p2Zvs0VvqQwaSJp2+L1o6WKx6t0Jod8xz9WAfW2F5q57dlcJ0IEIoEFxITGqSzUTUaz4XHaW1Bpz
drsWwh9JoGmK5L0bjP14Kgk1B91lv7YMPXI1dHRxsV0YzfueLVkDCjI/eEEGq0X1Q4oxbQqInGAP
iAxlkQZtDuhugTT14r7hqOqPl2djAGlOLmSqNIY4NGfKeW/1nNffd2ixdu9FDNDZEc7B8YJH3S2R
CsHTdPNoEzXqn7TKcH5MGnz4eOtXEUld2fQTecbD7baiOsHpH03mFwOTlamijYxxrV8brRM2lbjV
MTMaMEsQShrDdXI6TrXHTcOaIx6hBX78q5rzd37keeiaFSX/t1sAkg07DHt9hn3a/dV6utN6VkbY
Ojo9YLn5OXc7fg5v7Et0QEdXpBK5zAmhUJsFtdrLVw1BmoGbX8oWVAWEqI6uzxXbIHTwdWtPi6TZ
S0sKmLTdWTLXWey7bcvbNLzUyAlI/QKZ2uPQyoVkabovh6yGiylHKPgowO7OZloNUISg6nAjUqVF
or/TWC/QIQUgAGfPvI6kz+USPB4BO1V+7zDBJwUUsimvZdSVlJyux5Dz3UmAuR2bJd256CRF9000
oB7dBVHJ2BeAw29VeKKva/6qs51J55Wp5lyhar/tKYfvG/BsW7jxRZ58DzWxjwMB+OKaBSTlj2kh
vK0gYtCfHEwGFogtdC2H6wc1ByiNahuMsvvuG7nVzI7/yxlZBw7xGl0vA15ozgDQcPm0Q3mm0yA0
I1IgCPef3sgYD7nfxDxGJRvKSHGw83t0S5QUcYB4gLWjtT1XKU7aId53bslbod1jBx8zvw/Cu9rZ
GgyXCEOK0QcKqPBAYCrd21GnyVL+uzKMO/SsHWQjXoeq0ohQCCICkF3iXl6pz+a+4UHO5URp1Bg/
VvC+sf7wWBALN9aMYTM3Eo2+2gMq5rd01gvEoTAiZ/nGJHtiVJw8QTfn3w9Q426FV6rrK7H7qVG/
Pqjbdo7wvxTSW5wX711vRbc9xwlQsZ50LGvXhYfJHhsqPfzwhXSj79Ywd3OUaDzMGtIvYnP4X5bX
CROKW94/C2H6OVnxkg+MVnSnuc4H3ZJ9YYuqJzMcUtZ2ukbxGBthLL+B6UqBiztnaK8XpkW7Zxx8
1Nl/QKK2BnmJQnDvAfbztwHehKXx/Y+3rnnqHxspclXC4chWPV6LXgkWOlRaV2NHYzL0eo3LTq+Y
dlE+Kp03ww0WnbOTiC72mxkfmkFx9+UwoxG6NuATv9RM9tir6XiATEvAvOa1g/XPFaTRzwYvZQK9
+5HW8i0HGUrOcWl9hzRMMS7UMvIcaW+Oci5O/pBF6he/I+Xb32SnZVf3VOmefzoiy5mCnKO/OH04
DuFB6hZ1OYGCHVsdc9OrCazbE3e9kDuqKZpbTdYkNNt0zpTeF2piTHbGn9+8uiYEX3OVJz2rmutM
Ll9y341lALnUXOvI70KBPuaLwCcknFRTSkBHjGion6yNfVxF9vfCQhjSBNjPGRqWmG8Ivq/sAPQw
LP+rAawMgBJufHx4JcA/ntaYMWOlXiFwm7WjvQy+oWALuDNoO5JBoXDVLmfwvYunZu2I0PbZ/q/d
DrQvfNKLmLIdyakbPtmJ/nJQteIUsb4wdQ4T69nMcRf1yy8KtyaNfU24gG5955NgC5fV0SSBJGj/
kLK+S1ykyqTgCXpiiYrGs3ubw0Aw3PqfN3FhEW27SLgTRNs0aBKOy+5pXD9ybqu8eZN+/fT4wqfV
XVLzC7GKxz2dRRfc00Gt9AkCFqzfWro6xi5IM6qK6wq+pD3nam8gB/nR6OZU1Y4LpFoxsLKfZi7p
xmRCHvaL7zMqx0Op8u4mXlhHeC3cPWeQTuQDkbUCDTHSII/vIbCSQoB5XCIbNmUprfR+Az/FN4Oh
NnnN8Wq6AzGLTtmyC8otNpFhrJy9f8dSE1EA9d+RXMgJ9GBILMpLZgxhMgyu/gwdd6QKNB1/RlCI
u7NoO+XUxvZFInZrlEHvKm/94bl3Z/s8HOC/iUOiZsITqCB3kAReiuxEZJjxRaRTVKuniuj/Ce9h
UoTQXnxLur6fccSgIkuxa1z9wUcX/ALCfIdvtwQdS1fDDH1rimLpekKG0xJAGpYa3hlGPzvoTCJ+
F3+VgR1MDpnDrGBYWQQSgtik7Me+PNJV6KwNQxJKKSmjCKTIlB/YA7XWh32xzdMZyDDZBI4/zdAQ
iU1wdRVShqarEijrw1oenBM6TMmwwAa/BbUXsaCoTAjM3qNHUTR0BGYfE8JIVcp5gp6nJwFLdrBR
lpJivBgruhqdPgecuvBLMGeutHsQ3YK2/oiqkE4ozj60VaONAkDmbBSrrxMUGs9l56ga2RLb8n55
qKpXafRpGu8qvDQfFS+oRqQB8XawbD84nY4DyihTzfXodRncrtuCoUvcFgTeicGBG5mvEwmjMktB
qBftmDTTlQkDu/oSPxBP9HdncWnWPAmGw7iyUTZZs9QrGR+tXdqUcfzAEtQxnj/R0hVuZbMHt6Qd
vzjTkglqzJeCXxRwowU4lz7L2zfsIzqmZGW8dgMANQ8TXcRWCrhAv0xNrRY7blenbDH/IFAxedk9
TshaNPDOvbPAr9wVUAjI0tLPzH46Op57sTbTSfYxPzcfr3HSH2svh6QK6PswM/e+0eFhbi1pij0j
QU7SPEwHtjQQhmln3oiO0mFJvFsDbN+crY2kBpBD09BtVNt3Dn+O/UPDKoZdG/hYS4nX1TJRy4Lg
5bEeYR/vT6Ll0y6jYPY+m3NDXyxMQexqqTX0V4Z+xnDQYH82Dv7+b187TxYrwyl5voVVZUnBcMpI
LITjG703Mp9Tr+rnavZXiUshrQELKhzWjyDOVOOXWKyEef+DclHovCnxnQfFg2Zpoe9+gcAVLNsE
8b93pqK8hOfhuAgwsYxZ05jKNAbZq+yFOBgHSgaRszPXoUVDn7WNXaXC/cM81jobXw+3xCO+wRQI
Uj4xqP3N7F4mJcIEZnfGCk764FrsTXZ/gwFmGPJpzTUknfuAWxSfypbzEOunfMOCa4alBlpW3FcR
IxHUHw0efWKLXvJG64xUOyYnhB8+h8tDq9HuElBsQzA97iHh1bVthalvoe170o211hWdMZiAORgL
rvuNiXBSY27ANr2Xubahn9iWnKiMejtAEfXImlrpBmYl/LimvQGk1GLxRfbH9fH/Xd5nvVsFkZoI
lie8sgcJarDGbGco5kv/zdYtbec/3FfPRQr/q1ryeIKkZPHXOtVo0+S3cT1/xwcpf4BZ/pDgRy6r
9d7KegCItbQ3A2GnLi7istH7GT0YK/hJEiCsqiWnpijQt0ts87/VjXrNG4zzmMc+uP6Qy5IENnTz
uYYuW8qRrCIA1zQVc444snWYTNvAUcYU0Zz/LCWGd88NpXLA/dnncr05Hunp6R8gB1SeKmcuGqPI
95kFH3k9q0ewFlcSX88OLL8a+3zJEXhxGh5BGbYNjf57Wj/vxr07cQIm/p2jQPcvEuuq0Od5AhRw
ADc1rssjOZzSRTqeYIT+xwxzMG2VMgAhCSwxL90y6HJA4RgOqnyEdePiEe9tIBD+cs1H4Dd8188W
C3bpBC6A1cxK8qyTziuakWJ/9/Y2nrH+LiUgS5F0AwoFBpqVDCD7/V7jDxT2g9pXPH2w0wIzYikd
+s2M+L1aAHAjx+diOT97aeT8x4QgZy28x7tC04pNdanRrdL+YU3DX8TDW4CQPEoWozTg2BVPWgxl
+yU3nHgEOOW/hDeZ+YaftvMxZ5RiF/2ds0Lx9ca2KtuRgh9q73zCQl4qj9QBj7UGn9FIIB7F5mGi
XQvOjoaDyuYl16rRJb2Do2upDGx3EZPqa4V6xtBvccSsa5SWhHlQKNpCcMjmt1/abjMkvPf4J0xr
FnIyOduN2bws+u0Mjf0H4vILR/khYvRisVHN6+al/LZ/vSNReAz5LgldEiSDsJxNDO1td8B5wfXQ
ZCD3DbXPwkvIkOBFiAUAgTiNzQrPzPoR1HqDWpZrCK3/uDus0FGDSwKj61SAVHsBz9ftkyLKM4HS
RkEnG5GtpxJbUbFlyEi6lONedwAM95t79UqRvaD4U8k6rW+aBxj/BRSEaBlMIzXoLX4BXEZHBzwQ
BJeHTAv7ZjPDBA6Pe4EvilhMegX1er40H/Jp/vPvtOnOIs2iZGX/oaNjQaXCtTEtVGeI2AwzXDT1
yJe9BwHO15710auFzUmHmWPvFYT3Mb3CcErNoLqN8a3aGOR9U7gDL34aIyavEcHd9ON1dP/PJ7Tc
o5uX7anlRGzq+Y08aMJthZaoIZSUCsimzHnHJ21mI3GQxQeFTczyNx5dyo9doSAgOtc399/PD6EV
2axpd1mn1lVI9q3HsKbB1Zvop7MKcrMm7aZgJ8ooz6hBSSkqXd+zq/s3HGOd2c42iw3lw5QeAmjB
W+H2TXkmCis5m9lUGlpkq/EfkbhU+5C1lMsqVCxVH6y3jO8LprzD0UMw/rQCVZunlYnDp0iHEWPV
qv0IeBlNXQFm1dsqztwA+1Q837ZkSHY4WykJqUjNEUF/LU5A50ZAYDyAvMKkN3tf49I7L5xovqE8
yhvaS31EFxGaIIq6StPtGEW2HjhnaCbO345QOmpzA6G+nIoM04zrI7SbtvBE+0R21w1PUs6SzTdX
Y+k4+k8m+qu4ElHxfWwjnRR72CC6LT5hNSnWwpxYkyUQtkzxgb4S6WSwAH0Z2fwdUNgeLbDCmXmC
K94mZ5HSZteD+RNyCFN8ikt1mpSmxuahv/+w3SgY45XXqxP2/iJO0ZsrobhUHgB1+qYlSnh1y+ZQ
TL2NurMsNO+/mz2NeYc/RycSHK9sIXDxfcx5LRo8HL/mUOjlcmkfTCcjcmoYmMBRb7UafU8xMZag
7Jf+wKVWPFY/MMiE6vj9S0wJPFpvDo2ZWMpp66/IiK8bRgOrAAC+FhbaeWHsUsSTlblcaFk6yOBk
W0QcymOE8jYoJv+D//PShn6V3z0uuy6XJDENSJLOmveE+U0GjKeoTG9yehQMYZm+6E7gn02OFHd1
QxEx9nBwFBheUCbfkIMZHm7S4reCLQUfenpMTlqRXz3P7y9OQ5qgfZIE05URnFsJuATT1sWEPKg0
5kMMEButXAijN8TezcS552sFshh0anVmKtqXWk+naJIHOwrX6qIHU+eOQ57Vuz7Gb1rzTAAcKKFK
yr6vejjOyDnweGkLYrbNxHgdOD71LB0i4jqls3+5bi91aUXGt1GxBtDJRth3MsxrGVEU5K8tLYX9
V2/6/c4CjPBsKXKsdj8MAifQyyZW532/s51k+znuySzqUyDhApnF/r5LjjaHHnglq4K281SixiFT
EyXypCxPbsDWKlLrFYN6Aer/ky/61BMXUDcBsZZW3BVx8JDGjQ3Mis86eWP4cGG+s93Jd5weJbAC
Ja5r6Y/jazer/6ZSzvqeFmo5LQfcDAmxd0gYKKHvjm5AhPy9KEweAaBi8JQeOcEOmijVBd+p39/b
2G4GIejMfT+yTXWdOw79xkmQYmNLDYt8KomlIDY0c35KgKw6+TM5W0FEuJy81X4hOnn27x7OKPnO
V1JOcYYvjLXw0sAixk/QyrN3jxJjkV/wlf8QCyc2k2nrWQgr+sB5mze5/Xo7yaedjvl2zSfr0n72
E5TNWkY0QTlTjyV7smCAyyiN5lc5ekbKe2/8ZA0Pa6uCR0+qEjG/QaZZe83OjT/S7oJMVARypyeU
Zjp5G8CldqrZNVsrYeY09tjIIU5xTi0SMVSFAKfyGWncmEJUq3fEhCg6hbQt1AiCdmnEnf6Tq8WV
fqt4dW07zC6DyBc/EdkeQL4ePQgJHYm2Kwq2CGLDFXfpu25CJNrgNN0Zc0YzqybWd+XbmFamQMWF
DEuU3nfGc+29ZKxc4p9I9botWwV+PNI6AFIGYLlhCdVdS2f+dyAlMeVX69V2mNPsMWaPQ9e0clP8
sQ4BRMfhPLTJFLGzfCAyAcrgz5zjoaHFXIrxWtvw58yY6GD3IJ9IcMo5d2SNgurOTID/MVtod3oR
3mgondC16jUZthU9Vo6Iew1NsWBTV6ap/ft+Owzc/dDLJanNGR9ArTSna4lqyLOfnRaG50GmTWJz
dAo/kxJLjiW2waSQ1iLQYaANBUlXU3BOPwGy8HOOmeWKRiqNVD87MpwCnbZNNEbt5ohzGQTBZXCx
WfVepY4x22p4s1rQ+nhh7MpBlfZHl5FlqJleV69UZEItv8p/yAbzSyYi3zGakwQ4w6KKvQnIh+u0
pRoFu9j7RoKIKvE1oev0DWmgfMy+15XMx+Uh6Qi73gFDf8ACJDY56WSTuWLUf7b7H7BWCxA+/k4f
KkhxZs3ptVjtN8lmVFO8aTuybGMHWWjtVjsg9Rp8orraNaAa+5y6qNtf96/7obh4RoD6p6sVxYYG
2E8/hQ2cCeGr6VEPTHGgwlXrhjUYJcqDZlqyno0WrMPhfHSjEoz9RDFgMo1KnbBtr+vJXw0MTPfU
GenxcO50ASKTCVsOqoNjF4X2fMK7KumPn8crbe1YnTdknOHy2eZcgJPvB2ie7N3i56kH9ekjxwlb
ZbS59/kojcO/ohFEDAx3Ot54y0lgXJYca2SojO4JV92qW2XWE0BAIhwI6ygyWVgKbmAdYBI82Gp8
wYsAtNto0t3Epw5RMcKR2qQfkqo+W3JaUwfbPm25mAZpODG+YXKhslRe0XMembyxEWFki8rA2u1W
OfbhhhSYM86LgdH2JSaAhYdJLGtt8unhAdL1P4u3sG6hJy+puUsHbuOuYnORJKxs9Yz0oaOdXeee
lKehHzl7vpF6HxTI5Fh+kJHnCyuooGWl1I/NIsFz/JIy7bXlRPanQH0IMd/LAi4xzPDaI/yopAna
6rM0O8akO/qp3EdCvvlwlIGBPyDCd+nqsSRhd4IPYYL2XdyPY7gZOUxS7Vsnwsr39sMT4xHdho27
Cy6CW/sveMIS7GdyKVik7vAJ92JZMlVJv5tsMI5m1GGHgwiyUUUPLxw3bBo6riUCToP+Sh5FNLxY
4NRGe3KXJT4hYTrkAOCrZ5BcANBEa83wqQvWkEsM/wb9xX615h+NSSOMapp5xOaZt9f7s1y9canD
fNjwMtCOUXh6F9PHmtoPvuwlJhR5pJArYLKDulffDsUY2QHaWg250qprx7+rjP8/o/tuuk/dxZ1U
3J+92///bOtDcf8PnbOwHQZ/RAXexM2Dx1y9NC0sZS4OknaS0jnb4+wzEFgR0Eh4Lt95Hg1G//Zr
H/VZxDVT0rhstDcwXfQETdupEivS445dVm68dxfIjxioKVTBo4oF342sehfKIrwJfJmkd+r8rFBa
aagZYXv4eteq/8vDrA9wsOFfVtaKyUB0prd+85PmCvL3XRWrcrKc4HXlfJ7BhDq2t6Cp0fLkukru
InpPunrQz6i0CQm4ZutV0PyUeF9h/eDWbTKxCgUTW8jWJSkqWTlKl1ENHB/MNkqgfFH+d04SWCys
fWJCBWZnM2Urpz0b2X2szbkWuB8TZsqxbfGwkITQK1Bq7msL9tT8X+IyYaPgGyhRypZOw6/iNnyH
54XxCxcu8UcfVEEJzZhb2F9vAavil3uTDpt2mc02heiNzsQjVULC116hlx1TicQeiHJVGje4q5Ta
XzVWGbKeLf8bpgbaHkwbf7ZaXiU8e5NBP0bsvDFMBYMtIteIUqrakZqL3E8j4imwkgbK32P6XryL
d2ha0vLtIGTC9YJ68AAX5lOTF/meP5NLosP0jPRonvHv4g/YBrqnO1BpnBCO1Wdmc/qemy8rF9Qs
a/OC980s3g9qvV3sazoVItgNzovro+27XUN+0Oqt+Ici3v5n6G2nlsLsl5cJOmnQlAnlKGfZQpcI
RobnlJ7ILk7NFfpHuO2R6uvJq0ApGH7AAfXeRtwpiuGHerhbKsAnW9m2sQasFA1YvIzvChaEHSqi
p1J8HVHxeTQDFodC2LVpPDCpg+8Qab1IcBJwaUWEiv1TGtQe0px0MlvP/LQNWfET7qsyXKKRVyc0
2dGvFMgmE4+Bs90J0LaRNmR/UIlfKs+nRR8zP3dUNuPc30nh4PuxFVXGxI5I48q00UPZmiRhUMx1
DrTaeatXHO1SSH67npHIf4hNRPSb3Rv9nRl/kfN787OG85AN+HjCITZh0NzH27a/AM2c2Li3QH9Z
UMi6z8ZJYtGnFTxOkRl0uKL2nrCbLtjtCTzUwEP+kXQzomTLzKLFV5zRindGP67eFqVP/ryZ5X6G
/quMPibwdqeEMPXyGZ2PkHfU3iakT7zwfTbJca5T4AeNkb7dRVMg6uVyxDvjpUsdk0p+YLbRGPTG
rWieDD9Sto4sUFv6zl02YZ6TA+hgC1y9FsDMeiB75ro0ZvVH0yxn+hxIOTS4fsDLqRvbg0GZ1rQQ
coZ0NvSIczHVrRG/6AYDKWu0qpQeOCXr0d9ClV0NZ5PbRXDG/0n1VlfPNLYV65T481tSGS125hQC
NVTsO5gX2Hc7VavpTGmmD274zRFoWWoCS9t7GueeHC1oaGwhxTr2wbnuj8QOHmUx6WsPXHxckfQ/
JRks8semeC22On/56LkxNc9xbcLChRKJyc/iWXDLPKZOJJEONn77VQeySsAiYH/0dBlpUYIE2/hk
uVvR3NWyLh0W7DB1VpGeCgR30UAB//eIEL4aEMvJqBQZ9ElokxZq1/h7VJN9lxLT/mcTul2yf3aX
GfB+VrKrC7p5+sT7qpWyRmSb78TDfe8FjoLQI1Igrr+8KHvJ9+XeUKSk3f7SDnVYKdYZAhFOfEHd
KC1Jkahh30Rm9VBDQRmSlqQKndMu/SG1B/Ucwjz0SPXen1BK/d0AiHsw5Wpu5cCYIwervtmTJx5D
aOiW1+zpXeTFMbh82zkBluwpnKPLvR+SRQ3Hz/ZFEbJZpa4h+JBo/PJpn5rjn4j0j1cPn515pPWD
q1D3PfBj+FiN5T2q5XJ4mvfRwZRVClWJY5PD/9EcQER5KBWQiq4xtHjN9s0e5KMC2tjwqayqNwhR
9pk1M6sc0m5KYdeZpMcXoPXDeknR+YSinTxxw5/AdMbiCM307kXDDHXXBuSlfRbMbx7/eRR35dld
Hrw/jMx8ieSUVdHaMsDhbhSGJaiuky9dQsnHzef8W3JuC4urUP+bwraolmCT3rNs/GkXdFMJcak+
FC2xbik0LZNCKgrhZazTiSy9r8WfNbAuIIo6ZK9y/G6Lr/lhF70L+D0tnjLYhNyhOCMsXhOLPmpz
w+bU487hC7/bxqm6S+TaevR/YYutZKoY7rKLkr/NtXobcZ9sHERPJO1r4nVa/vRlEUk/AgEGtGN5
pesgDwcKTdzGw6UWnaJaa+TEV6e4BfzQXvvtQsHeDr1SaziHm2tR9a/x4Iwg8ZU6bgFxyKdwHHin
fM3m1KbUZO9rwVyKOFNQ/0zRmBbHt58lE1a5uScjEmAlurvN6z66DxT1vNhVVqrrw1iXwVfZUJhY
gInWrzhON6q5/z3BB9lQD/Y2d6QN3N7KE6cgRcQMVgwFhwl5j3ZpoOIHijEhDH2eLwqojTUKjPD8
x3F+2k0ye145sAas3BoG9QNtNiCwgJ70uws7iqf+wXdsZ54P7yV9MVsnwV/kYuykMlKgQdH/iECM
1Knq2VFFS0dPXJVZBr7sMfwd6yGpYuiXAhYq6JJd0vo03N6XFU6aST2F86E6CiEHOqss/A16cUGN
JJ56GIt5vKS68tRot5KHF+BGxkyHzfJUokUcJOx/1t43AxJAZ27Va1N5SUU6/XGaHW+kkVIQM+O7
bKFtzklhvuT+j2ozF1KMVg/TVGXlxoO9aBU3htJo+/uv6FBGoAFDa3PkUqBaZumVHA48MyP51nl/
BdJmGvI8mdJosdAj1R2rTfC54aaTfsSGJ6gG+hXfPQlwmHj5C55XrGKwe+wq7vpeO3BiwPHqX8sY
mWqR/RilLt/AJGQb5+R/AEehBTpOoYW5wOchub/eV43EIbnsC3xXYgEXuecZpAE+lLM6Y0KMDHnt
9iyrzstR6myWS/3n1u/Q6oAZPl13R8AopQ8RtRSbGndVosRoq1+ALL/YddzcZFL/nf7/oaNzV0cI
IYOBuMw6et5PkHerUeW1pneH/DhavCXbnqi8pNfk0WHlWT26XWDQjBDTnEMVfN0G6bLF+2pnDdIx
AaIx7BpAmopVPFjUUhUuuzB84nMwQi4OwUUzUccytkX7U1EQZ1rKoQYaxr7N3wf2H9UOik5b50Tf
9k4IHig9Ii+0SZXSKB2qtVeUC6o9V+gvgdTB325jUnhJuU7fjcVeWHoxbz5ibQIpuxKxxboQzckt
ra/9B32nGdZdtcuqOakmSdETzWhSyv10cZK0cPAqWNqMUq+8Y4iWY6AOpMWxn4cWhR4c1qQgc3YA
61kZQhAtjuMZpTES+QRwsFgYCDM46SzpCUrNQCel6MnI9brliI7oHK352jnXA0JqI/f96x7EaZwd
V3XMEa0No2PuzTRBOBrKUG474nULc2l4aUUUiUjwH2p2PC9SRSFDD+UYtx75o6j9NF397UWxeOpQ
9r264xV/jZi0S6OkduxHVY9wHlQbsu9rC2dhgnyoNAfJOcCcLI/jznxrDzFqk/fmjSj0MHK90QVr
9vWInLTo0k2G37Fb0sI96W7fpEB5KYZwGPkATn8NDwPYAFmVVVY3IMwuAzkhlUo5bzusASvvnkKt
T+MHQ7ErQKrfvrW6FFO3az6IxnC5FrjBkLUrbemm6JaF79usb3D4t8QiXxiqO2XvZjMWKgi4b3GQ
dVf1Aqj0xdg2H6bLD8xXR/a5OOL9QC6oPbw2hgvrkZex/BSgEtM6dVcp4Sn4X4l9yCB+Dg5JnN39
7tUUemcrMNl/NiEbzRe2QsHaxto9eLiuMRAKU9RBjiP5RlAbq6TZyRD60UBhhrcfVm7YLJ8nE1wR
nuywroxe1oBXEhbH+H8tos+6FcWGi+oHCiC0TxiY6khCl/9gP8ScoyO/QztqGgEWh1FjLUHsFGe/
BN3LHU8xNhJ1deFkoSSF+3o6X8EK8DcTIFMEoVG/qExHM1ECR6JMXzCLY6q66ZtPMjBbHROwY6xk
j2NoZMID8zWruhUW11B4RDu/xeKa7bdXCNR5Yf9zreZX4HEMRvcNlR/zg2VIS99FhYZ9yPXrszTb
m9Q6LV2aVR/qomn/JDXVTNR0UpyfPs17RlaSEbq3VBacTkGYyVJIHstibfB53yUlkoMih+3X5Jzw
/p6xGKwfFejHfjDS+vfOLSJBmahKgXrQiFsj7rScHMD5mNspYuUiUWUMU6xBk0LDK5jHZI4cTWab
n+OQgew2duN2a7R4JBXCbVUj6fvvyaXnLnISQnb6xaXghpH0eLrlYdUPoqN0vWfnzYZxzaf+NJmx
OSyNT7Hc7nWI3eIAf4TJY8h+fQn7ndLD+Qmq8T38Xcjf7ZC3hZjCfggtJ7qV5fD2K6PZ7W7JtCU6
mLW+y4/5u0RApSNx22PuwP8ntrz21m8WpsWmrgFhWsi8LgY04cWehZc2WBXXj4ffRezP3+iJogwF
PNzMBRVs6Lu0ZqSU8/xBMSTSCOrb4WM4NptD2lo3OUxiobIyxCZrSKEUhCMOBbQe9zbQ6yUZGJGt
WGuTzQXNVgAOjcp6h9/MsAnMTDYNVmPboh6BZ25qTpjVjMIfUlPz0ZKXi/OU8QdePv8YhK85F4Q1
er1zQQMvoG3XPWBnhr3AZuHatKhw93qpK8GJtl8z2LPveBs/78GKn5SY97Pe3kG4jN1P4Q6XidoA
bOWjy/wtP/29IdndvVgCjs7A4hq1kOkeEdZrAPm4NCISlv1CzCzEJdW06TSM/B45CHGY9NWFAqCq
4pl26PO5Dbg1gmuRUjTcQqvoxriyBnr1lvg/CIULlnQHLIhKgJIMm0ZYX/12+iI9yY0UOEKx+cb0
Ic1vxI0stQwrrfHPt10IWTSjr2OJmdOmo+2+veYYldiic7pFapX5/mV3DxVJZyziehlNgDv8eviP
Muzs+zGs6UWrDNuMbc74kAlb/eij1LwGOZk8Sye+iYnHtiUYUeQ6XbDuCvOShDUx5fWx6xO0qRJl
aIgyjfLRvkZJA07OKHBCJJK3rf13WL9J1/g2p8Dx+gElwbzNvLkBgVaAoxDLUJOKsgb9R3tlzMvo
TZXg+RPV8ao8OMsWvTablpqlM/2G+3Ns3FEuHdCJU3C2ywERkO/dpnI6kHteWzkKK1eEBhzO7ig0
yGSzp4miFFAiB9974BwugIcrSIJ4m4gYleFsz/2XrNm28ed+6hIac3klbMgdFkzIR1lROKsSRz0z
LmuocHwKkC+NrVuOLCJgsN6Z4oBE/ptnVS+Ma6O+YZwuHDgt+kMc4d/qOme2wVWUyXVYlZuLEmOQ
duOqmyODrbNbBpmARK5HSC0HYwl8UHuAQbPoAYSInKep5tHuTko8UTrQLouJiw6ozZSDKIiy79bm
p7Z26IaCSlrbTupANSc76L6CI4yQXLJ5HSE/xu92yXbEPo1L0RgJjnmJBLleLO7nKXVM5isrM6CL
RGxtIcL9k4/xcpv3GO6PUIh5jIr/6thmx0mPM8VmCS6C0GCip6Pi8WAN7XayfHzR1Z5dAPn29C9S
vmbNb9aZLq0JGecVXPAf8I+oiGejQFlT8MuWRQQjwJIWlFmVMrk+7p/Jzs1wWU+87APXj7yn7h4q
gwajG48mEmSocTdsWLIBcwvwTkkOKJ8lXad7P5sc/e2OD+L66Rddlw9OVmPxLSGrPjKteowi1k4e
WE+QPUizoQuUI887VgIcY4pKDBMlwQCl6xRtgi1JUfzW1uX8EhP0moIgqnKr6TEx3SGLIlxHawaO
/JT7tgTZk82S2OLh4PhKMAEcXFiBGQECfs0EvNY5EinZPOS/Z6jcSA7b6B25FZj/U3CGA539sM7n
6AbMTF/amWg/aPQgpSG/MKss5I185iRvGkxYVSq62GRlDVqvys+p05hvR3zjmN86/b8acESV9fn2
ggFoCBrcIwnwaaB/u63Z6NzFs4FWHPkOTcwCk6KHaBvkT3D1C/dXSYGCNOfA+I8xuOAwB/CCiVtM
BJW9VqoauxuvQ4RBLG37LYpvIxIM0BcbDZ9YxtFtIV3QlleXlBj8tltmSyVOuLgxrDLZUVmiv3VR
YRDIdeR5lRURuS8X1pXtt1gSPK3Rmhd/hw380CynC45siLTBSumLLT6NpcJw+jyKwLdW9NRbkcrr
IMQTgV9RVKAmXgiURwPkzGxdekCRGC9ngtDFoSg797KtSZBf1rG2IOiFAB+2wQKNlC3Etrrl8BuP
5lrdKxmFW9wakkA1+zucSilbGjnQqkqEwcNf2bllqHxSN/GHTkSVkOZafg4ZcsEF7aIB0v9kiUWL
/ZCd1Bu4obAIXeAG+FGfaY4cYcfEYEjF7LPA0Pwu8aaicuNdRE7f9fi+1QbqnQlPLZXiYLHzDeQB
R0Tf5aZZfW2ZAAm7R0rchjJ6aPzRxw3TsmhCu0fO5e3mnPH8FkiHj8NisRJ+TN9Ih/gdRBH0VN3R
sdDyXfNSuh8lbeFoNA0lio5SqXUwuEvsQHS3DaKgABTCcc8wcWHYNRBwEMVMlF/3i3lRXXgz5tdd
gf91URII1pjCZCKysF1o4nsaDANtr3jhKnRdpSHYlN8U0DQ97c8pmJb6qfmThfeQ+culSuYB5nrX
AH4mxNFbNiNljoI3H1CFcyevnmkvpHy3l+Xfi0EFLSISK4YTaXmQVmpFwOKXvLGyQIASTam/ZjW+
8EVxNG54ySgU1wOPw82ejw+0er/FbnEq0SGVYIN8ax4X/nKDV7659uKlmBqwkDm3zf2Sa4rhZFs6
OsES+4E2QC/oQBcZWwk1ASfJ2qxLz0hXRTpOMwLwvAt2so6yYmjCS4C8tdNgT5Lf0aEk/Vk8s9Rb
sI4qDtqXGUPlCpHZs2VTC0zolkeVyscI6cZ685lLN1/x6cEUFX1gE6RH7tdDBtuYHHWTOr+xRR1Y
yOu3EOP/Iq9BPWVrT4LSBmiOqKSsrAS+OBe9j25F9rkAnFs4qF5iEsi3mTSlZEE1FJKVAErHZPIi
t99oj++eLat4VWHDBOIBBN5eM2TsSN8DYDpI1B8t5BEfCiAPKAYfYapFmJ5Jfil4ilOY4BCLT7La
57hc//3PJVG/i7VvydZMiuAMYHrgO0aiWW8rXy59Oe13MmZ99sb17Z5RHidWDfS1huu4JvPNwdqY
O+dDD16E1je9pXiVxWSPYGcYf95J4zdyjF6UWOibrmk17BfRn6ruzuBjD+kEcTDuRXlOV26xfTrh
NC3CYZRtFWHZEMjdmA8FjIUvfWlxCxogek5knlWV0cCJNkTqimDpnL9Ct3nrDhX8CKbTdZ8vt5sm
cDKY3Yz/XczS/hvoGy0nFK+Y5LfRklXmeUULLOpnpafvklQMrj4gEi0disVu0XJMU9cg1xIfoBDG
GhNlFjUnzWxpWU+6lZrnJnDhwd93fnNLvt8XeyKUJ3EGso+Qk0xkgFjMpNHg7aI+ot7IRapQuWpk
ItHQ4JTjiolf3dYmTqfoQscLawmhRdYUFMC1p0mFLX9hRYkk/Ir8fsAslZgpRW87YI1Owixsik3A
mTY3wU8f3908IjJfwp5JSYg1hxNCFfAxLk+mwQdnUnMHWqJUYF1YnDVkTjH2fbz/9HvYAso0UCzL
7m+bO28aTxl1v6s12hN1IiCAwm+el3sU1WhewyQrpmdSe2b7sG3J7p9tGGGjyMfRzoF8Nh1vmysD
fpdEJHEND5W3dwTGMjVVRjYRyq4+CnK1iUST61oqM1mJSjeU1ssb9mbx+UKu9Se7X0EZORNuqNx7
zCU9P6gFnQDGynFZAEqmACAdIq9HJhc4MbBav1v7aZBBL2CBRmhgSCOKUeTv93adh4QlSDWL/07c
XlF4/NGrMkW8K/+3po3UDQy0d69irkjPtPDOKjBjBiBld4zwTZPFU6LfBVJPKxzXurj+2ujebFu5
L4uqrhlRC8swo74OdNc5qNrXMWdWk1rav4VEnKNTND4QIpefSK9pK4f/2mp58VaiIyypSqpj1+kc
3kj7mOAZ9x8+XWOrQpPCg0Uq5YfIZaQMvPwQGdWEJYUxa2YNdP8IzmNfV4nTr2S+AZ7VdW5bXMK5
RCX87HaozljCXp8vV3+rtqgMLiXnPOYODF1sjockPNhslhhUC9TkPG3+KQ7Mxgds6/mjNMQxzOCj
N79K0UMVqxXe1vxiMpJLpujFEERFi3XH6+2+3Yby2kjigMmG4E6Bd+MaldZWdIwF6U0UYNWdj029
pqPTAp+S1mgFtOz3/KOyrBCGJozSrpq4O8lUf4ohA5+5U6O990kICdW7mCZg4hDTDs7U5tsm9/cD
ItysxSvm+Vp9C458/A7ZQeU0neneqdKWPuH9JYfoFj6gYzfq6+a1l88ImGwHFg/Yc1Vmh6ziTDo5
ehsVIlboFxwIWhYhGSy8sIOoX6EcuMi6oFYkw6WBr9Gn3tsUQd9JEnzFazvo6fcuKgzUrPTL5Lnt
qOSRLQ1PoyU1uOD/66sBiPfJfBSHWJlYhWu8GZLlyxKUA9xWbjIqCx4L5z7psIXqiSPlHD1DkZB1
JnNEZDJoW1VWJqGlbOQLW/Gtj8KIei76rmGB1oiWWprGK5z0s+Jj9dWDxi4KDtLae4pMjngJf3NZ
UU6eEi7qkVbYMs7TDUBQ5xmP8nqpdEUkX5QgaTEpyf78xZpaKtPwooPneO09lxvhJUdVQmLWWs54
RV/tnTkzdpGouSCxh2UfsEIRJ2hENKuLG4U5KAlScMzzpAM70R/M7haBahMjmNBHw9SBYEsE+RaM
T5AxQUkPQDnKJhdrHLV2m9f5yZV5dqcdQ6f0x9fU1NpNJIRAgX59p5pmVcdpR+CHNEoL8xVc77Fl
jZGEfapf2TbXyEmbjeaEm8fI8QbzgZVpgkcQhXec5Qb/aEtMzx58P7xYqYKQZXTP9GN42iQOMffp
odFOk9GILQdLzxSqosUyHvX/isjfKcaoOhQOhuqqUsC5Ffj/n0ppLlodeD4Aaei9zh/Gq84JvAlO
gFkbqhV/XQyaOBpo725XSxDYEdu9h6lMCS61nRyaWKw3HhXhETHaGypW3goxY7C8y6pToBF1AVSE
gEpQxMw4oipgCgZPxhbDp/dwqYqbYuktyfnD4v4+8jey3JMGI5lJyPndCw6W7IBTlxB386Jojoe/
3+bPRSMYez5k+UY+yYIQoDrsXZ5uLoLVTJlVVdTGY56mdpbkAM3U1xbcbEOyez9eo6u+5hWQKKl0
8+I1m/5n6J3iUUQfA68iieINkTAaNiEL8grcSCrlSOQU9wKLZjHXdmRjd1admcZI8zBVb2HdalLf
Cp03GOQ78qQX9syUW5w0msiTLncaDaP+Kz4hiqnuUrEciiuWzW/MntcOsLWh0gfsKPvmQMAdnpjx
wKktEH7QjdkzcSEGMSh4446D/Q8A3uhOIhSpMayf/nG3TNb++Rv/j5o8aZziVPX6r/LYwHn8Lkbq
cEPXbA1Ms8mp1Kw8cEVLP9dV5U4+hqB0cYapeujgGRbPrgxSxtS4oBHrZ9y01/PbixTaCDDh7voL
4JoumAjJSW3wAo4EPpJWm+YHhWrLGACBfoeHZs4HLTrM/vos706NRCX50d//c53+CUOYLpNWbfHT
oqnZX565Mh5gft+/p7WvbWh5YPtcHS1Q4OnlTTvHHJ7ux7O8cA94UYfAELHmxD20IRAaFmAKiG+M
1yLiPh+Mznhtb1K7an2Ia/4EOwhJ3RO6EW7v/i25vlgNnohHwsPPoA7DjyYV9utpI+nSOKTGdx58
0x/NzRzlLVltjN8DWYzLIHB0On03qb1+JOGOdmWhOhJtxEbfYByLoJnGu/FFrxmJn9gPBSj5Bv7W
kwgpsxzv+EMrSW48y0HFsdqAJJYyb9ic0ChGVU2Wa/mGM17qRQtwcsdOe1BtWTHtsXngJJBiz0Bw
aiBeLP7nJVSRj1bVHCxXLC/+T1LOeBJWzafIlOSxFB9RzboYs6YNLkPcx/RT5j4UmkBOqJbs0PKT
p8y3EAfJbhwkdSpR47plgf0Uw3KlHohLnSF2keu+oatDhLTEsg9WndgfrnyDjoG2lg0+lZCD3A+2
gcRnLpiWPPXlp3mmtSu5aq6prXysmLWzCgn7VIftzedr6pBeCuDJMPeUq1BN6cVHo87xRB0RVf4Z
n5TYqU7c24JX/qkWregu5CSOVTuq5606pao2PVgNDgTYBLVnw7meXNbURpvicbklPBB+GkFfMOJ3
aCzikz5OhE9Egb6W22T/yBLELYMjLNNHLY6MTwcBMVnqEfrGd/d7Hl6KJ+B5ZdN3YvMJ63xZP00W
xijqeZmPcR3B0foWkXf6IjnAwg2yaqsv6IFDW9xyK/uNaXQu810+yNB1ySvbpiH/MUSAKcfi/r+7
JnIniBNSYNdwu8AXnvCglMRNUNTsR1DcN75++1fbOK26RF9+LHV4jzSOWyeRHUW+DnymrXS/cHZy
CKU9YkegoaUiTNkr4zHib971EareHoeDH11AZKULQuIYLTpJzD5Zomk43Vy15py4Wmf8mR2WQFMY
e+kf/JV0yBTEdxsuQDyRExtHxrQbZ7LtOJlvi0J9x4eN/mX4V0S8Wkvt49n0BZJ/drOZQkgZAlWl
eRuM7Rs/JTTeaard2EuNBEJzXxiXd0atbYWmbSru6rcfqpmYK/jQTXTWxYlspckt4YJ04Hyj2kRB
CkTIRuLpjvXnu6cOSdt0VeqK4xQox2hZGqf9p28KkA5EOOpG1CxneVnwFsnlM6NE7RwTMp3ufKYV
jQTtfV/YpVeqdUPxQGU9T6dkLCL+uzuHVrcwLgchuRQDnZ1gvBEh5Eo72Jm3kJdFWJQQfWceQYAW
lWe38oM6xmBEAz8n422rTWATl7YfraEXjHU5Dgr0NYGG3h8ZC98qGypikFSzKtXzwp7R93zD3ybn
6y8U1mucirDnH5z7Y+2ZauW6/BboIDuKwSvf35kpSahoTZLChCxBx3hDMWRO0BH7+NzNlWcNPbN5
tWTs7sU8OH/8F+mkhtWSDrHqQclbH1gWYZf6cr7WGkVaN58oDPWBTkk0XsbWdv2UdYTuva9cDolc
E/wXH/pbMWJWhZ4vw5mVDIQYqVrnu9nkMwGzWf1ov5R8iTm8FNGHxNIQbXM5Uaz7JXEfhJpzaaTB
7nHguOUpItHIASHfjrPtHTWFThAlvQ64PILFxXkwyk+rjoYnJHYevrpGdXnCIcH+kH5ChS2CWAf8
MN6guk0cBixAELMH0NWJzTq6Voe+iao0FgUZkytEH557LgFlROGvDigs4ro9F+2xjBlYgAPolwAX
nGb70n4+OxDES3VcGgPiAQ9UJfk98h7Jw/OcD6lS3mAQpvQEhQAVM0yk3WNiYFQ06Jxab6CL43LD
Yei0kfm2rkyQ8UEfWpUIPKiFNcMiCn9j1t23TkgQ9W+tOqCzAx2r6FVfU6IGigg79b7h9cUx47bG
zcdFFzZdl5y6yjptum4LSaL9E/HLPEHdAnpaG4hZuy5QCqcrBwU4lSCkA9BcSvdoRGdwkaUb00mq
VbeY6J31DP35WYRTPG5gSOpKK8SgPjF/0JJcOBFDSG3/nWM5fswdDcgm1IAnenOPkCEaLnIf1YNw
mHomugH/gAUda3lDNlqiDJ/0BBCpLEyEsv4ufg5YZcGb+1UJNCvNTihtbUTkTIA6dXxgQTyOPLfU
u7CS/cwtmJpwucJ0vZuETeyGNm+8+mKjyX0rgt+dWvg1ToRWLkIgurwSPlBiLKnTViqD2iHuJOfo
lF1W1DZL+nMyY+wKcBXiJUAWjNB1K6Oym4w9gGXGnqRlM8IApmZHVRD1GyfLkc3ggdVkqSzH4m+b
NMyg/e2GpT0nYtBG1Sy5cMJ5VuqGkKhHKgW4yl0GW8UsUhDjwF08Qr9otdXZG9mQNaajum9ZYfMt
Tk0PjCuSRydwhjMEJVBXnxf4XAfe1YFm1X5VFTsBE+AVcf6FlMgnRBlmqYLeOsaTCiAyAJzMwx1K
YsPKFZkU+0DFbqTP1LC8cwDeNO7F11Gve0yMgaun88HNKx7eIjgRoK9Lh1gbGp71JQJnhAuCBEq/
j1bzk4IUtmPf2FdDgeExPYnMhz8UGH1NkyjopiyEwKnenciw4/3H4/sPws4T9SMO5QlJ5VXnOd4v
UWpFBF4CTtDRde6nlgXPDLsvuOvWB0DMlt4RIJ4fezfJy2YO8ybSzzSY91d2koISC+fCwime2phr
QqU9D47hPBR9WvATfJ8gQvFdIDSMkcefCslLm3mDbv1cXOzqwmT8smshBy93svyh0JxLzXZwJmj7
GqfLWAR9SNtlisW00SHxjV7B6S3nQbGxS3uBLwbdcvLf+lMhK55Z1HhIsq9A2RV1h0yYGosHXybx
vvhw6OKx1GoISOB+c3S9lt5D8BFgABfUaX7Om7OevAm390WxErirSvovU+zis/D6zjrNlra18X9X
GZ46f41qJEFfecJRX0emhmRGHJZ6Ev93D5VU09aZ7669NRdPhgmIdPEHvoL+Qy4yPcJCSYVvAmn+
arL79snHZ7MeK6v1/0+DjkzOK1ZH/kfnNWguDuAd7FYzlQpgCgKHkNY0vs+taGRrGEtlsC7EuJ86
Iottzk3p5s6fh4AAj8Axif+2R+Q4BaAweaYHUE45z1EcytEWmXSN8EDlTSz7EEWpEcrBEEz4amFq
FvBh2qrHALnykYXGU0H79ucOLFrrHDBuyMvkqg0cMSdnzv8pLyYzUwBIc6KZkDStFKiwDbmeuW6+
vxZOz9XvgzGw2QizhYN2XzRkivSNOEXTWdLnNynJo5JqRGkMZ11X8oLeq5goxZi38MkFu6UtThAy
AV6bSaijEkI0Yg+4aTlwKzjyxUAbYdyAglT/OKGgiH8ur1aa6Qg7FWV70bSzimZ9SvIyUFAT2MQQ
rV5ea6Ags3IZ9YjXc4YVpPtj9PMwfDUc+pTr2jDVXFYJhtD9Ryb2St7u80DfR3wgEBW6HuYlA1nO
6gnCYMNspJkkfGLeTa2dd+vCXQNVlhr710r2d1Ecrj/0FXIfQjmostaGKKsj6/edRaV4sQuGCy+e
LX+wBs91qzvMhh41O1hL9HORjKJPXbpbTQ7NdEgW0PU/de0Ji0GX/TFjutjlLYi6YTqWyAgsZgnQ
Rsnkizged4KaODmc/LTv//CUiwwqUfdbVlS1euzNLMczdEuL2HkJQlxYIzH/534b/wtLza3dA3h0
W9VrDAuAZDXD/LgzVRyekKZ+uMPTfboAvQ5gyInEfcg+AxUQzPqSBI7bZaX4IKg/msmYS0yf70iz
DzFdeQRaHgQPwF3HdZ/UHIj/k5nPM8VX5q1ElGg0Dthb5slIqjR7Xw0PDBZQQ/kSPCHyQIw4NGE8
SLcnA5qFDwzzTi7+Wg5BkHd2wPHtv063qadQnJKkk6FFBLtnB0PjkQoRoyHoDzutIV8Vk+V/uUgM
BYqpPtjmHJdD1pZgTxnvBZ5H5Fpn0ONb/rJauf41Jv9Qrw2Ds5MegxbSkaHVwBJ1VFPHaXrCEyg7
Gr+ZC/oyIPDFPj0gV/j4New3LluxpYFTkRzVpuc/wwZSTlF22hmyTyiaA2aGaDu23PwbHrokiY+G
4LI5eR4+b9aye3BBGKpNFaqy3CD9eCOXJwOZ/+tX6FFpb5nbotxHDo7HGhbIxq1jE8zDqs2eeFDW
OBR2aNi0fiTSklrFnGyKEe0/O63iDafNwYZJHAi7rS+7GMl2Ig2Tvj/taUFYyqRT27ARYGF6U4mW
lucRqKAIAvM1/5jj9TWEX5x8UQo6zVAP97z7ZEk971POatXdPU7iymWsVPHR70UphicRFNbhfgNH
9SrK/gIa4Skbji0GKGHknprlGGjG07pSD0iNb3uV1uyholypgAja7Wa2gFbrF46nLZzFol6I0YWr
P8jye6vagxdGmHNewhbDFFHasFxBDiEGkyv37VjWIrwG8Fcobzo+MbmAVfMBu/Jw92dfCxdxY2aJ
zDcgrH6Xqi+szFO/Q+WlWV1KEj76Sfj8nc18lePpilrC2WaVAxGfxMwcfyZUkpqom8LvE2C3zWh8
B58Ff3QlH5nImBkq+goLddF4fEz2ejRYOaFUFazHw3lOFrB/VBVMzTT0C0LQIZmE3vPwCQoJgZrL
vxi8EGQIAh0EKGBWuQuupH8n6Bxxn1lfdCmTrI4xrvdXxqoLm18s4kQQnNW3AcWDWgG43APQ3YGM
Euy9D+ctGDXHvxqSkp4m82nDuwDU4/me/4ORfJYoHcvYBEU8HkSOONsaYzrsv0AiT0rp916PpTPo
+RWxOdG+FLH21rKPbM3E9myXM3PQgCs6GjCnWWhUXlGjSKDURaRI8CMJD8623uOYcKlykuELb2c1
1y7HS+AQrAh2XT26c+pw5viXpEyvOtNZvXQAezrwk4omZqBzm1v0jI8tBd0nNPESvrw5AQgO5CDz
9a6aUaOSj6iKSn6UCZ5zmkJTskJ0ARnWtWvXb1vkkKDWswFxmGzUPSql29pnhQJgR640fdrLk5Vs
EOgXH4uPkGukn3WwtshLRsotInpiXIDg9z0BaDMVg/diTbtOVSwaU/1VRPE7WeOiQ3GooXAz04ht
NGmOwomxT+MtoZU/Z4h4zbUbdrq1S7n70tyg88q3j1tmji3w8lSfnCUaNg7TtrIXr6RFTkM/9ZRu
5p8HTJJdeZybU9X8CcfaeFpOgPuNmj30z6g6FqVk/ORpi4TctQbcxGzebIOj7NyDKGsFj9pT0dX0
FVXO26KE47/u050H22fQ4NonJXG4b8cqO8Gn8abEQ3wpxFw2W134tF39vwLYY+EgKD1y6RujOaYQ
h8p3mRc4zT7EjS/bSQcsYYxqrWrvx1aGqmZEjTzpL6plgtLES4juVvXa6M1qS4A0RwMQFIhA0AUP
KCXJ301d1MwWNPXe7Kgk/GzTWG84hWQhp1W7OQdUAPQ0jdXIolST07e802zOk3Niy7hukkeF2ROH
1xU3KTxUQzVAicYhJ9Rht1Jrs71HzVkLVfhaBbsXY+QhxV1pIlJBO3Yza9ZyM47GaXNLEMqTw4sI
WT/5oMz4Y8Iw60VNNLjjlfMx3noSc6bN4/AnXlgb+IkTQq+umWoxBtNN9wcXMxqmFZeuD2JudeGh
05xeztnklov88ReUFSbzhnoYtmrPeCapjkQBzYHP1qsVcpY0W0wTawNhvFeAwvK6dGw1Tp+OS8Ms
51AACmQyC4S0Dkxh8QP2KfUoeyB2RA6opexN2QQI0xGmAiXu8zlvKxt1ImEOUJRRv8S13rWu78ev
fowxGSCGuDOlKt70v9zlLD4i6p0vbtiWyzTIriT70O2mqKRlFm+6wlB0rqt58VdKb3KLvkAxONe8
JCDq8582vNgN5Fvbe1Hk+zmHDP7LYP6RX5/xzBSfJ3AN5Nxp/lJ5UKIMZzfPzgBRVpFd5yiRdMNY
Ggn0zuCUWRFVXVIxZ930zdNT30FcZjt00Ya0j7xck7DzMPg8pXfo2rnqqE+nm3hn295Lo9I4+8vP
70M/pyWSMdKPAMb+9A4Ox585duNeuqDlQ++ROeF46zJRImpot5zcUifES+zoE6pfOvolbsrYM0mD
JDaUfj/jRVfY+nVHq/Qo7B5OXbmvyYHBy/aQ6mYK0/ZRs9CpSRU4OVRJCgEotiq66jCV7W7SIj3P
3L5NEnorg5tyLrwzaG5IlvSPi1CkQRApdSb88EYEs3mXGYqmexqttbZsVh8jP/oK8sk92gRvtsip
YlOdGZ1x6HYPnc02/jP8HKIXHcgK/Pdk+ooRw5UeR5KTmDsQPxbGb8cH31R5HkEfV/oziwJaT3fk
Nz9pinBOnQ75xf9KZkK7JVThxJtiMzpw5EmxW7ViB/DzTVhqQ9Rx9NmSaV0MfLsXvF4nfJVIJZQM
BAY8+oEqkkr/XEo4BXL0Y/SkLf+d38m1S/mzgSPUv8jQf2ccB79X+5ZGxtPh5K8aXxgoRA4f3fhs
9QRQLVQlawXB79C58e+WNKzgHnZk8qIsLmvUk06ATVU5EcFkxu2AVcLESr/ehomhaqdjcx9i97I0
BNi1OLpwgvoJGG39oENZrMjTHa4N7CZYHkOfbfnvUID0J+alLICCOAI8fBxgPXHJw4p4DM69MwTm
7fc7bpqHKHhTkJ5Eckj7ikloAyAWK/Ec3DwPpwVhhxOIPuXKdwnl2Y691+iWmSuZsEXkSJlOE6OZ
SZrAiJ3bFmRzybrOzlE10TCT6+C3b7XaZfi2ggGqmRQ5DMR/QAHJZlVeWJhJNScgpaA6rGvi70/L
AU5LSEQHBd+TFmQMFRuhHQOPYlnDcgChqOMPh8OMAgvly0uvgIa5QfBqpW7zlab/F/iH/r4DNUBk
7vqlPOLy0/hZAT3D7NQ07vnmG0X0uohocblDd6FtwgDMM3+IMYY34dnVI6qtNSJUmpAnTtdY3QO+
fZrTfpXkA4E+JGfirkB7sL/kKb5XGjCt71vx9NeFBswqK/4QbJUOgb7o4z28mL/Ud2TUWr1GwwWQ
4LxDAI6IA/rTNK3iJpcv9dfDUYEoZoO3Mqt9TPTrRWfZBvnQW2azXF0EcHF2yZ2PDsSUeZEoVJkj
WW+WC8vhMEV53m1ooe2F4gsHr27YiIOroD86y2ClammKN/tkuu/wocKKAjdfOtNcL+PCJHDs5nSD
toHE4/47vUPzYyY3+zHTniSnaRng77892gye//pdqm5uFziJeiayxy8BjAoKYjMOMlpETQfcUMdP
FxvAlLixRqDebg9EHKgvcB42Dci/SX3EeBqninHGRukSxLazSrOOOSqLL/5xyAgRSUqvv3MwYUXt
asYDg48oect9ufSSGEDtQ8p4dJiWtRN8fBY7GcP8hxFUsmBab1sJSDizrz+xPqBdmIkYmZMTkHR7
2e7+k6PYemMtkfTjFiOscoW6/hGKodhD+BchOPzppOdAQqMPQ9DHC6GZwcvcrYfUUWN/yD2pSB7Z
f7wbkXaMIZPd+KIO2kR5B6bQxMW7qZZzrJR6b2RhZA1AzIrhUWBKjkMnnqWQzr47Y9wN1LL+OvrW
yZCMdeirFGvnb3dleXM2RlmQr/Eo3x3pE3MFn3UHzCj+TdU7DaCtkqAG6rUvzZSzWOjX709Lr07T
Hd84O+O1KdMhn009HQp9XhR2AnwhUB0TCmawDpAcGqhlRnqIPyt/dS17P4i9BbLIq21WcDDE0cF4
XAdZLaI1eYJ2co2t/DWyLPRk8beKcyiegCgf6ny14GA97NCKgxkkhxPBRTT5ipZ1HsJQLGzqCm56
eyqCCPVlY1EVHNsIN5bm0ijgq391BON9ad+zNV0ErL9AM0sZx1GiLYJeBkjjiZyVa5sbpxM07TwN
P+TrKsStRPjwICwGu26gk+TBcCkUkyCNTPxPi0OOkBLCXLqmsovPIiRmRr+Ld5SCAkAoGIq4E1sD
ealdmP1EVlV2v3RK4psQwtJX/drqMO2jd/FP+K8oFq/JeSrITZt+D7dbXZgEw8ZdNY18vId0PNih
hquuwVJNInkZOTtWkzjJY2+KtNRd6e1DFMPIUCZgglY3OHWLjUBpMHUYmffCSErYYbS0XSwKkZPO
P5CmFBnhVkp0+Q1DfXf1v5ouUOsfB6dKWbFnvYVaLc+MzztustSOMQdEz5gUHOA61tFixh8uCGzS
lMSHBbWeztnpPYKEOBSAORN9p+V2rYPKUsBAVuoFPxWvsoMbe0oIlqV4jUflR+qHbXnLBd2y0I9J
2ySFm61v5kaF3M+i1tIZNmWF93hDS5joWMtklvAEtTfpjJmm9N2lv4I3c9cdOsDPI00RM2uNemBY
d2HeZMpa96SfiYY6WWYhL/EEoyNkJNxL0jySab7iwXSusdIwTBdGkLWSzJCcZQsM4hQ0EcB2w2kT
myS/29y0Ltfi6tXMSUnRM6hUV21lBJM7EKP+xxhQ5btQvjYjKlNq47cKlTq+GdObNU2eGok7UpHK
t8nhT4ND23kvqAYrdZDxZ1CC1kbg+/y2bpnAt/tNQU/Z3CXWo6acrBiRyjG9uGXkFm88H4uCaLCP
Nrz+WQf2kh0uy2Wt5WoqmfpfD+pLBxusFCChUs57BQTTBTpveZL4tyw0LpyKo2s0l1GDpRTc5idK
hvx7p9U0/THJIGILxRkoDgfb8+7RO/pYiRcddmcLPsPwDWr2aThErOXEYlF/TUTOz8TPxpQIgXkX
RHqJ4Y4cpS8GqOPqzytop1M4JawzpOoYXIG9dsyhJeWJpWviKVu2ZtDMkgCGdvyfXkK1ePV2GVHk
+4S3eWbh3G8+NdFQu7TWwWBn+wxFjAlHkJ+e91+1ihuzMzj2bvSQ6ibyOG0TOW7Z1NukV5R/J7yq
TdP22/4mN331OSJkFIE/LwBrBbz5LQJcx0QLQDYUeJRGHkldZ05L8oOS234uYMzMVo4zVV57xn47
zM//hB1jh2hLqvR2L4/0g2XXFvSpaUR9M5PY7ldLF520MysUf+qBAKHLD23C7dzYLR3OqszGv+2I
3OHOC3bHoetFp5f9D8FlWdLztuz/gAq3HH8OV6dQqddqa9NSykT3Wa6I7HzkB79EWw0lJTd9JPOT
CB9YJqLdFWpITBJdiiOpZ/Poi8thne4oxxDRXoTtLHEbKVUJBn+dvNtMF1LWi1RO7IZvDf3lmJiF
W08Ueuzc06SKNzhaWJprezxa9esiy5UPdru6I2jhxQ+NwAaIRTQCSCNtD6hmDYQU349txlf90Sek
2PLtJfeZMRXkCn61Qc5dQbeiDV9QP+K25/KWRmdaJtA1+7KLR8El9ouGYYrXFxXo4pfqR3uURBux
Zi+XxOoZL2HD18gtoB/zdnCAlYbqkybiEaBcAN+T3pzJkFaqbJs1Qfz9xOzPwCoKI+mA/aCowx3c
CZk2GRNGHYSjkQ3J8oOeAfbxNh9epZtHw6bojtyHzHMceMbjzISZSORCf6iUdkX/UFfMzXxyDxDB
4XnyLIfTegENlldZz4HYcV+nitftvdp/KFuooWQyCkg6vo9viRHjEndGV+4+aguLzW8GyUJCVuD3
Ti9L1hr1iXftUobkOU3tV5Hmvi+7zr2rJM1SiUWTliy1pUwhoZHS5miqbnRG3sYvSKdmFodT3jV4
BNUM6w5r7+4zQVPTXvMUxL1x1cilc+zmUjloc2TdeT5BKBW2k5aDtuXlcBCJbyC2aSLdWvPZ5T1D
vALV2qEzpnjowojl5TSomYV2qqeFqNDi4bSWHN7LFCiqK+8/eLH3ggU3kJFDlbHzbFsHSiYLe529
LGJ0+f9BshLWt0YovDyI2VZlRozf9yCGUzUSYFRKFFlaggbhCwsY2XNLqDCgpbYRaEVHzAidJzRZ
HifNS93sg6rAZ8tiUx+vaa0tfE7SvU4xm+s8PbbsDBP836nse5Hhqj7bS2Hhi0CLxhEZN1tfCFp0
c8nqGTbDTAmb2NcFUvGFpqDpaiXmdgExoJgkaQHTzYV9LhpF0cnO9vYtHkms4B7uFqNHbxGsdoue
GJ6Wtr1h5eVzx9jMOhv6QOZIDD4nccxH0xkqCdX39AxiYZHMEx7Hz+ysa/m1h+95XWU51dUQUwnY
fsB2Guzlk84ZNJoe5VL9IB3hf0090dRmII8w9Ueepa9XUfG9QifQF4abRN7Ln44+jzHjjX0pYXrm
wl1cXgtlH2hY20m1Dx9p1SJjUzxC6yBZcW9ycrgeHcZaT4CCuMAZ67a+t3QwgYKO+/disDR88NEh
X2c33tYyii7Hhk5oT8U3hsh2D5EAIgXCRrAbwB8fkhlXfsUvvdzZ1dYf0NIsJ0WvOC+Y2hdiTwbr
G2MwqL8I15HLgyzd91935pSeE5PXZbNof1opb3giezzG+vCQEEMVV4blHc4FKewUYaawgKvZZYni
5OUCSvNbOwrb775qWmA0SKp0xh0HVefgnuEeukCWL2ziobX7WAlH7ZLCLNLbNeDz7X+e0lXglkbb
ISXh8wx8tsBqx+sVBRvxJ2+3AhzQdja03mFf0LApXDie0YDoo8Iy9cz3ZFq8wYbIvpEnU217FE8b
hs+zQiWvOUab4O7zfKxKZmU7hu6P22dYrbhu/E56hHtMBjRm9KYthEXAAYA1qmJpfa7DDouMVPkr
RF3rE3sJmp604ILMlQQ79o/oQsac2ZfW1u1zSPnPwejrk4L2Dw2G2YQvuYrEESfnlCzJBXn6p0ld
zfBHAV3lp68ImVjFd/vVl5tatjjI+45zaHHtyrnapKWDfZzjElsA3/6PcJHp7L/4ITAJYA7ifPcO
SHTzUTn46gDbaweem3CGvr83qu1gpEwTDaVQRzLKcHzOjd2zm8eruRw8XuLOK/BV+kyUHOgo0//M
ZPb8bz9GiNs0XpZJFcMvKEKoTQCobbDHUuRQ0DPhITnAnfV4bwfP7K9P0T4y+FSGUFtJ3m/B2EuZ
c9Yii9z10xnMroXEn4QojVCfxSUyxGBVwlZr7tE9xFGbwVYqmhMraxi3Rk2i+r5vveAUhzA3EZUh
rjgpsQbQxwt8zX4gnAHnuqOf49FOW+Z9w4Hduac4EnS3tWHOg0PVBwEt1eP/AmeDlkattLbT7RWO
gU/Oc5106fxPKNJewZGkugccWaiPWYvpOJbaHcwhSX0FBZXJ1Yox5qdq6ILp05uARCmcCpBQGvj5
xmo8uNiFtfm3EuJAINOLwhLTX4V4Qx1kwVzh2XCCqQmbvUoluH24mq1OJI2swIUN0TqLsjUkcMhY
ST/TqucMJdIYdnY+z9wUOTQBtyXgAyBjMlAe7rBjNOMU3ZStdP4x7l5mkt7mm33RAqcxqvNpITj2
GWj0fdYMnqa7Lfd+N6HLk7duEYPHLeI17OnBp7TW/Hf4WBertDCU+EAJz0sEmjdF/U/YkCg2XZca
8socVFzsdyNt5eBv5mF+rKWJ+uU1PwSuYA0Q8zmfjoMX1k7PGYpclSpNbHFSgFGAb977sspS7V+g
Kek2rIKv6p34uQAC7IXxudxEdcP/Zf4YuUy50dlrwhDu+g9Kpt6kyklVhCA8MJNgQtBto76smN1S
Wy4qrh+H8cPn2fLyzdKftDWzwslAx/H/4OWtIOZP00aXBisGbqQq13PTgkROlJ6uyKVTXBmeQNcu
RHOirPWfpfiZEJ2d3cz5sbxXDXRkr6S/jZ7f9c8IdWNfVQqho4WaFRoBLhC89PSZ7Lr/6yyMirWi
2WoDdPHrfQDspIpuLjTg321S2Bf8DmAzhf/F/aHbaCw+9rH88uOzcAmJ8JIUDBlBwWITTOaRLzH0
4IJh8njJGeQJOIgP1/VuvzoYyh3Rnas+SuYsh9bBmE9WKITJd4856gbk24JwNjvHTmL2JKuWpJP3
pOpNXTXmszAKr/8w9+ozUOmF+ER3YVHgnh1D/ayMuV6VqILunfLJY9XI8loNhIHM7NRU8CYjL/FI
fvUduPjPNM9+RoU/CLoQCVriIj8VIn3n1+HVajIXbU1YHuN6BH6TOUJ3CT53U5fEUWhphhluTLwU
2kygKmcAAjryrhJk+sOe+In0iESsR22z0K6k0utVlilTGZnGXWB1wauB1eKjdTsUS2gqv2Cmsr3f
O3xqe0IY5ytwXUCwkBU3hHusg9ank0Yt45hOmQe1CaVc2YN8PswVq1Nv61uiffde1AbyFZ2hGoZm
e/Bn7fnO/YeHEovzIQVMl6X88LKiG/i18J8bctBaOvXVA6JoyS3oMzde4CZEV7D2m5WYdwymB/ow
up0Wuc43LRuFzlqralSny+MG6TeRifyQCaEChnxUk9G8QY08MkmAIk9UqWO/L76LAkoRWmbHO1uA
PtSsEHapl0IL8YOD7tF7bALdAIVdLOg2MsjZqeQ7+HtUfN2x6SumLMoN0dehjlmzLC0gA3ctgkc8
Ex5L9RxaNxuCe+3FdPFz3sbJ1SI6eiJB8MObeKyRJlRUW//oGCF/UFsWuy9zeGrv6mbMPzY5jERd
pcGBgPVtl0/f+psThVJrE155FWnnNyxf0TaGVHkDvWAPZH2WPsve3Xx6Hnva4eHGr4jKAQ6wlQdq
zjTaFEc7bMtvdfTGbkJPh2dnHhK/7Iok1tSO6o3ugZ2q2O6N4415bPT0kwqZO6BkG++K4GnFFprU
FTXo4j3cS4+/NGM7YcLbPZXS9Skw4aekCNYebGVfhbw2r6W1R8I2S64AQmqT1S0yx6B2Ad+Xtnll
kTtzUO/q4Ot5EFw3QUrEdFMkcrdTS/NZbVx8Fx6FsHzaIFDybpBysfCdy8lliXJApqTnQEj6Rn9Z
Zu0ZXYKDDzpL8dj32EekG+6Z2ycsfMGKixa6XWsJJ0x481AP4fAgI0j3Qc/HgHjrYe0YvMiuyREs
NkBPKvnYmL/SqfBjelV86JuLtiOhpWApPwyBSgQU+o0u9xEaYioLhtQev88vWkT2r6hnOXq3AGyx
YvdH8Rigfhn15T0gpXRdFN9Xr+B2cqi2rJXtty+RbCqgCIctWOn2DEb2uFKIk5UK3sK7sYBt3s5R
u3SJpf9Eo/m0RRI6THaYc5Cp5n2AxkqtXmkRDgMH1vcMOmJbXi00LeoIM7maR+O2PODeo42rCkAD
cKIDxxy8WZVnEI2jiHrl6cZxph7zj+Zo7yO6c7LFE/xnZ1xMQbHzXMLgrLtHvw3VIl5G8a/2J4NU
4J6aoF75fvmB5p2VPEFU+/rcEMdd5wHztoBQRo4+ZkkeK1jlZfejP7DezjfA8jkzIVKeNyvMpkG5
XzMS5Lzvh6HEz3Yklu/8mdWtInyHwid3KPa6OkBVHtEm3AxAFqQbqLIVOBWXAB3PZxMGAYgGLfel
MpV40Vr1eSXIsMNJ1p2OnSnAOw7EV0AitnT6SXrY4xznyhK8deZycoC507D2AsKd2FYwObpWv5HQ
PKNEjzyMPJY8wl1CUP1XAqrC+Utran6VZ5qvsAdOlfkuhA45tKgUJAOMKs+JfmbAhl3N/MrC9ENo
LQR3lj/rkSPmWwFqcwC1Tk5lXnAJa4q/xkiE9s07lzUGwrEx+sTe5DpiyQ5bdIoyn8bvutyp0l1B
TwARi751CpBfz8XzyQRHIDzj8C2q3grimU4nWiydwJa8pLRgwjLTtiYSMuCW4ygxsoFGA1S79g1B
8l9wyymfXNuIGP4T848iokZrns7PFpuQaXETHeJNC7dtyQ4MkHPH130umtt9NwzFCuG5jCRbzE1D
esFYGHIjPa5Bcp61NijfkDNPUqLQPzlk+Ag+pZlW64YYJF/WxmutvdtaQOSB4e8CNEJTzvMiQR92
4VeKBLvtY/CGmj2RBb8WpSGYsjy5casFhpvAPuYRwQJfbCXpV8wZtbYysbKx8v++QZIaVVRFfisu
nMfz6qYVbm4vCgwqTW4dMcxseVjyXCsahO5Gu/iMwR8Ezg4PFvgJP2nXHXUOaLlaUXEKg1Bs3Mlr
jV5oAbr3wSAyIduobbAQiEo3vDmHU0MY9SrBNLs5Xbu6ZuJjJta2l9mbvFgarWPc2QW1MxizkEfs
n+u9GemDrSRVc0b02yBeebNoUjnnVix2VOyYONVI9ZBbYgQ0uqoX8njxxgJUNe7JNPzFYE5+n24U
Koy8v7WEjMd3DHNGQB+Ehhu4xeejWWzk1Oj07so9IpKw1S1UApD7ba0/hIQ6/ivU6Flid3RNcEHW
FDB2CorN8uFeUH9XcbtmLTQ7N+BP7UGhM4LjtDFL578g6AcnNq+0R1tBbwp3oIfSAcnDUBRzUAp+
/M3+dpVr7jqt13v6lv07tFnRfFdFYnFk7WujF/q2wf0l8XkRvHeG8WLNqH0sje/iLvkGGDFIAZwG
gX86MxjtS/ZsMMMf9LHrNY9c/jRfPUPq3xw5nlcE+4UG2Fz/6IflQrsughgSJLY86y5uZdr2z9md
jaiCgaSjhls9s0d6PFfq8J3DDR8yX7SM/LpRXtkWUCoSU5AaNpWvfLstNNgX+eHFhj34UWiTGUQQ
gL6aKLZ4zsoLwwtZRZ03UKvfL2/qkrNFhhDcR0BeqenKqsRDPzO2NZleJND9Ucmb40wKJed7dl+G
0Wo4EnYh2mX9qO4w0pWWvy5uiCEfDhbEY2036BD5x3LbPpXnBcpnQapIQuY6t2GibFwYwTesZanP
ufD7e2TPH0zIQyd2nAE7leyVqUtukMlTYcVuaYa8SYY1aNRvela/3iWEsej2yE9mA7aRkdYgaOwR
TpKNhRICRBp8XTuI7lHLE4UlQpyhg1gKh/OUiXtAiaaqVXiA+3RDGSBDauT9bGtMmJKsvjBkE2iQ
ZPI0ZwFmUv/UtHJIgrEk7oP5Rr1yu4ZTVU9n7ZkFMehw86srZ3GfY/ssLFxak3+/w/wc9+ldOeti
60vi4VojwIwwXw4/vkfaeubGdd5aI3tUHhsxqugWfsE7T4Pd2HwQV0mcqfDxfOsRX0Hu3PQOItFP
EEleOdJp+8D5TuQnLkY+RW0ieCkNSJFl6Ni+3ikzItH4skCnFAIhmv3G6Ly9ezkMIIa9n7G22g7h
xV+9ssttBArfl6s31ca3eCZmtR2W62Ao0Dlnf7XAD7EGb2koq4r1R8PQqk87ATrdITzFxmmbRAk8
8RyXYbcTWQrZ7XtskSWegsDgYoQNSuRjlCT8mGJIfhc9MDd89Osc1eQKtMoWTjgkSo5hEANXw4f1
PArcFFyvZx6rXS6cCqGWafkakKosQJUlZ/F/ylD+E++74JWnI+95EI/Zbocqj1pjBYxoOZsAIPhP
sIcZdLIflL96eeRt9KnqjjON072BoySYmt0yn2TIlJggCmO1ynU6rDUa2LPXr3+0UhZKoX/HdikH
ZqnQsY5g9El5NioR9WIsGGhufhbCDnBV0i7nMOCw1ZyxlMbh7PFxRo7aFw+yVuxX6cskzEd12nNA
yAEpvsC854mYOokAR+dFqDWgZASoIph2lVrzAtMUeb2wIGurgT+mZtDpFANKK1A/JyGt2WLJc1Os
KhTeufaiS0O9k955WAyP2v1A/xRC5btGDUVRIsp/Waktj0Zv67HFbDVt1xc14RqLqWyiJ8ygriUR
3obK0M6vCiiUOZLe3kRcOIoPFbITCu+q0hSu3Mt+bAyzo/BDoQ6lX1MOCYt5csawWMylz3aL6suL
Cb/KTfgenBzd19MXWF6EhgsD4s9ybzU4doZqmFRmO4Xig3vwT527FOMk0/dJfOCGp93fLbHT9aku
VT0RKtivZsC7fEnUu7/qL27bFMqadqKdTWPYkEi9y+joDX8LUHi/GRnLvuUxTAPP6OqEis1oWAzq
yls5rIOGqMwRkwOpVz2ORJGUtNXKjWmboF1Y0NYWsgQiY5Dq41UFO8v1km3Yi7v6pSvzCVBu+Zxo
TOYeZH67koqHyK8N5+My1oZsTBjZtfCDq5lsGIvPxtKZlSVL+8RmxxDvktqe/XpOpL3oYPVktlLK
4e40EiocIIwycHuE+SZWmvLjXTsGdXF4EgVCzkrmXd8/sSwU7KUdvnSy/TOD3eydOWIt47umzm45
L5CHiIOGokTBVAVxw4uRqy0PPSHJyLgJr/ODHGSyHNxvkNPnCOe1pTIjmh4mUPAXcMSV4V3BNUjj
jqZQBuyymbOp4hrnZaS35b3tqODRHOCvsN39tLKXE3J0RPkoZwyHFmTAyO6fnO5jkMSxt9PwCtp5
YliYvTHgMj9hX7tdPIYnbLuoQSx00zkUe9vSxanGB5kryatOljuWQTEDMovuA2WQFddZqgLYuOOY
s5pi7rs9zOyU/tyBSTxeOONk/xDCB3we7eNIudfGx/tInrANOhHCy68Ci1MMAS4Vt24xdJfodbjq
Yvha9DezCNXsbn45GfqjCOyPZhxRE9yLJDuB8peDVyFOJrl9gdv6GATwGIWVpspWeUjdMqBvgdok
kecys7t2bwM5/70Cz2Qe9YzdKDX685cIFz0fMNOXyk/GbCTPcGW9mE2rxnwEz+5A0D07vE+EsBb4
6K0ZTjngaxF/1OBMCYW0OjfnCHI0IPReOIv+a7iI/MKxMt2mZZo3dWcLAFRBodzE9x6UURRLIQwf
kYq9TtjAy3cEzLn4j63qqHUt/mOWghATBS90Z8UDXOw3ZA2llVGu3CIT3Hi/87jr0XiEqjkMTLcg
odnBgHDatlDISDw7KmY+d4gXfyxD+KMhHoSRuBE5zAYOp17pKBhpa4K+HZWGEc9gYqSH0+24LYw7
gKvhNuR7JzWDreXok6aqq1YNUW8E9EW4AtkUYE2JSMPctEgfzcIyZd4aJkzElVm9rxoF6RLjcZQG
ajGQFVO18mfuvz4m8OH74cyWyCYZpBHVM3GSjdP0kzfxrS59AzmGDs6qGepM+9eSiUWGDZTICNkI
ZbhMip2D1mmiIb8mWd8LiGC6jLs0Y7IS7Nq9siD5fLfV7mrwrhaTjJ9KS2RZVoajc4gFF2dUDdsv
HTlZDBTQn96ShSmFZ9MxuMjrKKifTVVlOQAZGTaDPuzG/RIQDV8OO/wdGwDXkridHTUE38oF/rM9
XJ5o56y8KLzDuAZHfy2tRqdshcnYwWLocJERI3CLkOXOgEJ+oZ4aQ8jIZd//Zu1efXoaFZ1JITJD
f7d48AdBD1pODQMpWyh/Gp6Vhy4tzu1UIlFxB/u2BtRav7mux+r9v60sE2UhYhej6gmwVkuy4mop
ls8qLzZ968tzLO+nMnhCNLfrYIPusgnB41I4MdWAXGu0LXaPk8AGKeuMaQ+gpo7f4Yr514lsc21/
RIBL/eDGe+/wQH4Lx9YkpNaiThIWlKFRLVUsX6V9+6gy9npskSU0pOu7xseGvIIMsx4nK71ziLU0
ltDpCitPmt3epFbsSBD8lP1xhOTdWuZ+cE4WBGp911snkaeJ50ciVTB+dLAfkkYczvEn6cze6KJs
+YUnjTVh+/osCAD69/50GohSkr15XqYz2qidUfA0ZB45xNO4dp7xZ8loXYq0u4g/xC1Wqz+KxsT1
sUuqAy8b11H8yjTSNcDNsKh7VFhIHLzsE+nytdmTnTbgGn4FjhIlzgWEwp/QIP9naJSTworSmy1b
83SiQ5u9Ukx2FKgqSlYm0Vh5AoZZomx9bb5HE8EiE9NlTbWPEgN9Sa5AH65hU/ZUsn0KWssw2AmB
QsSPbBN7K20z2nG64Dk+1vvXSWH8BGr6I0lUvnJyYIWZUjDXO3NnmZ55ZQ+UfmlHUtiV5hI2Xbb3
J1UsGdsWWnzS/He0C9C7FyR/kQ2hitkowbW4SY0UhsZLZlj9SebPheeAhfzmQDzH9jpXaZWGYqIQ
mx4SWZCiOs5kU1K4xOPZDLGFrT19ezWJCjDqk8hA2XltMKTpwLBBk1NOfrVJu7wloatsWXj5HmdP
tFPoJ1D7D8tiUFRGxuW/lVodTuamh90lk4sBhFWSjfw6W5HyQ7kLjMPlWameJV0CLJbxMAX8BdHx
d29KZIO3pULKCOcDJgDq0GVExN3FWdU9rHnGXiIXFLiMMWuKIJ2oEoAl4MEVumHv8vmJ78xatT0X
PswuLnSqyr3HdCx2aP7hatplDpTUbmDrDgLsrioLoOqzG6kFXBaZQ0r5VkFvOwbuAEHgMRPb9LFB
+eMh+xei/ooYyNmuiia+6RMRIybOEAdt4Ss4e/lQP9an+U/ODS5XMOn9m4wR72qhtJjIyvbSh8YC
5csS2MjQ4jFTL52C0UfSJM7Uwfd3bVS+/NRLG1ffMVkMj7j8aZUhpPD6Ss3cE/xZYn6WJhFKPo+K
GKckILfeAWZidkcA61zSdoVjobe8I/jo9ygTdkDeDi6oLeozWDtA88EST3yVlWnX7iWAJ2fHflo8
4Ge3qdRIyMV49OuNTOupjMQZThNPKlQ/GjgBcgTZkBdv/7i1t/Lu9daRuFd/5UdFwHN/w/R5Or5H
xUSjuZv0ARHoKR6jqYW3brgV+95iZoh6EKz0uExHK+a0TGILvU1Z4ENWEEACBZDh0W4t5qCxROQO
nt40MYMCTnsAcoqVStwL9uXUSSEW9JemjgGzEwcSUgX9cujErw6Nksg+TodA8msBAik1pBlcW/lh
ggg+GGH4x5V9+y9JWd8qID79NgL1FPANeOuPoE7GZsK4jdDXXAkYgrqhfzHL6Xul+zdoJDboMbM9
sQbHksxzT/X0zJtUJ3KNqPcEAbmcM8U/G4HQ/gp0jD3aXcZJhi2Ri102l6LXPZCAB4gdndXJY6vx
X4R4T9IdTSiU4N5CBOiRuv9X6dy21YYZh57C7nOr6eXl0JqKjNvRGRCmEyyVSTTb2tN4dbZN0p14
m86GPC7sR1a2miHJYIn05YgkLHonOCoPjf1e5q+o7K8tsH44VSuC8rEPAIZUh+mPDXrtg3cImShS
AtsgYUADAofRQFtc2ZrT8VuZD4gWSSHg7zBv20KdGGBulq30bBpkoGdPE5LR+H3EmGZHVW2SZ+cr
nVz4XkCJFs7cpivCpe7+DKFTKEg9sreAfAoSHcRD57ToI4fJQnl20C9Qpn2bV0XaezJS/c5DdVvB
shUceCVKqOYxKhfI1BJVQ4/tdxUKJVKuLx3dDdWk04hwt7vo8GnJjYeKzumkx6TNJglA/GrrAg3L
pVJiNfelTJyXrHlIzyJuz5FbpQwcFPmO/+n4SV7IDwSzHjl14o39UhOoqfcYIZM5XT7M8FTRljBd
XD+t81QapWBketftO7QcJg6I7Z74wAdK3sxTu7/PgGdO/RAIdYhXRhJcUSaEiK2gjKdkYp55D076
5OEyrkFak/KbXMihezNmMYvwI+5kO90ABMST6R6FR4Jitbaw5Psxrl2NRTo6sCLUwcSQ2TvvV/2u
7+VdxGZ6Mh17/AG95UQNqHk3MoS8dI/NtS2La6eR9vxQm3Pl0gZq1/EmZ2wISVu3xKCIA/Ij+Zep
lE4IQI0WncXGNKPxv7FuZfaYS7WihmXhH8CxTLviPaA7hh5QXf77s7C8HtX2L/Wx6EeOx26kR+am
hqIsBCEpAzggbqU7Msq5GurvioJXgZPhaTFBWHGbtkdD/Wb7FVESBZFdUlLrTWaO4r2i/Dya4kBi
6H4Pf6EkKwDrSN55KTYd8eiCbElv5Wa7uPqRkNbWKTeZ28TcSVeNBShzd8t4BCgwDMrMHyRuvFJh
grFhmXQwwIw3nAzp3UQ8KBGqhelHe9fT5+n5qjlZGuZV6BOK/+cvyzi6Be5cNIjH/CF0z4aKm7jB
yFMT1CW0A7KvebgEYtqLqXe5hJTnAERx7HkwpOun4C4iJUJRciGfPzRDy1/t+XHa6UFHr/UZnhnH
LRENoKDBU7qViFILnQkSN+zzHSA9IlRoPDsS8zG+fEXwloZq3giYeqZN77Ka44FUuTsFenl5sxkn
M8ahaKTUS+NMfIF52s3W5Ujfa4Yg4uOItAJYh/hUdALmsBpyxcyNsP4UynmKer2d2V+jj4Qvw9gY
Wr9n+gFU7LGsJxBwq85CNTK/JOKa+bU1xNyClKqQBTq2AJ3u7m/d82h7PIH2sju7q9YUQh56KyAH
RAWlTC8X1JLfWvrFNM4fn9LdZ39P+iySXp7LGY6pjLaPNmV/6KBwj7S0WfocTiv/hmKMkWnlvbpg
veLPcg/sQndx4I4pDb4kKh26wxCyUmayCcunnSjY/hEU0LNkeZ/zF784CxEjK1Xv9y+hucZpVrN8
mRZGh3ujUJjlMQebkewa1RBz/z96qDqZMHbL4pDcP+osWRdEX75XgVR2yrOzTCQC0HWHdHXfV7gO
8rwdGCzAwMdGuN8mLEzSEyQFPkDQwmSgtaV34yanHInp2AZ4IjNkbEarQ7jSs//Y3LlSbASpi/sU
xbt5QTbqIwjseh/jrVd7tzh4LxE+nU5PK8ZW7g3AiTOi++gIyfSXRncctzxsQTTLEMnI2xkrt6Cm
qVbeQVLuepY4kdJl5N+oGPMvRrZ6mVBp2M7gedlWiers3FE/NVVnEv74MINOId1PVQBuBZYPEtPB
FBq4AOV/BW2p05ou/++aZPpxbzPm0UpmZmdLF9ZgUNWLwOCvpGgchcQJXOq1t67q0kLj+uryy5K6
eOzC/iD1UtWUT5YcPcrYj/vu/Tvy9lWp7xt4Q3u+P59LZUhnidpn37bIDdRkbxFjU4+PxVJUnMt7
0IteCp2+Vlgn0HBACVTgk58iwZvPCBrLtmERrb62AFRxcXiQI0eldOg/yVSrVPJ+jIJOuW3C+Y4T
QcOJcKMgb7JWhM2K5KZck5LdZ0SHBEhjZCBQQV+ZFKlI5cpKp9vccCH1f7+oJY6yb+6Je6zopaIj
c9wCvbN3UM7rNZAP7sZcsLGKGx6XPO3Ci1WUWXcUU9L94cfOZ4d/1305UxPTUZ87RcDkGy7QHy2N
rHGKHkUnryORU/Ol4oJpp16Jef4BzZHXBRa4aAlU1ehPRNfjoyUhxpbpjBNKcFIkT2GP00021hwz
TiGzqwT/uufOl5SmNmKlz/DPXnP6SyZKIb60jRPeOUuIUbqxI+FUYvBKN8apFF87sqmcAR974iB0
2GoJxK00FLiDY7HK9mGL66CqADMhffYA0L82ES/8Nze6/ubVni2NG/uhrdvoAnnN9FCz1y7k8WuR
QzNArrr9oqhqVhQ/qhVMrv/MdruAqoPW7jhRzrkfoM24Sa8RacCZNTQ2DqZ2n5QFXjEPJ0Vj/ThW
yg12NNtutXoeL0IYTwVUI3HSRjQS86w9C2clvlswGJUVhJjKLFS6SI/rbYHopsQBcWTLdx9AtzGg
kvuxxYGkFYwvkNp8VG9jxTYUCtqLrPzh1k8p/IfifcPtbN45+ucD+AgRRveHw4092Lw4d3Ow3hqf
N/pVPrjLdmlD/PMp/bJYjqyWxYud//CbAoK6PoCD3uOQ1sa14DICX6R1WXmAk2RUjIyTc8uPz+W7
sChSSO+nklCE4anJIpogn+TlEowOEQqnxUQGW8JYqa5vZTXgTf8smSTRFuuZxdpcuoPFo8cfjdLm
mOxvpTkDMEfb75orOcMk+opqCm2flx0Uu2I79qZSmbIjcHNAhjq6FqrURu/gQ0zhboZgGINEA3d+
mM1h5WpSttV+rlFfRrAT3DQE8abV710x5dpZhu9ud/uh1o1r1Coy0BfZiHLEbVk8A9O1dkN4Ql4J
zk88SsmsIN1mCygk58QyC6IdvUGxbwW8KgrA6EOgDnzBM77SmdGArFKKT6pJQr/75h1jKQRtdxTS
6rYqtNA1WplZvuJWA3zGnImvvKy5jRUQb0m/+qOVeMkPgEjKuFx6vAMVC47Im3JDITXABhJYSjCB
Dim7Mskiy46nk4wamoHC/N+P8Nj+cSGoZ4Ef19cE5/c8L2oteQ7N5ZU1+yCKQ1iO38pA8iEYHpfZ
9UF+BPiWfBOF1h/79NNKKEW61BUwyyGAfQzOl0qN8fxzXT0Yv5iCZEXbtOQlocdho5Lc77TZwPgO
NSFiFAkKJQSsRqlxsuvyHa6BSnhwAjBwI6JMsdL/3l2c60zV7mMeNHRQmrJpLoKXlMFVrn3BxJDV
dJ9oZwf5qUxKUnTsxq7FmQPh5RTvoVDHDFmGTxrwJNjcVmw2IFyWTS0dtMuLKBSRZ57mm4yHR8cx
+GUgg7/KKXpnOtCmO6Cua9Pi/SuNBRU31nDEO0jr+nnXmWhluF32o5BYrTfs1KvXGQiLrO2FtVxz
TWPRf8Gwkoyp8rl8Ev+nA3lRGFgKO/guZP8MU9LocpeJnEkkDVPC1EYU6H1hdKVhhSg0WDOehr7S
MyPf5eogjiSGd1RRVS+iN5dcRKsD7piQdMubLjYJ11sMzu064ANKboa4bNjijnimgqqCyf4fK6GV
DX2I+GZr6mLbJOXLy0a+sMUSJN+r+xw1TErA9P2vpIL0UjV78V3CgqgdgBDNGKK9Oqeyv20mGFxG
qFInw76Rvs5uib+PHnHdHpySKAfiIh8bKYTlWmpfjgp0iVpqMOOze5AE+mboaqVAaSGkozQ7092I
kGsVnPlhZXl+stCMhRrnbeJkDbEvuCkGFhieF0TSFUmEBzqcENQPysI6JxbedqXgnWu100n/l4eG
UTVzat+bmDv5Nx2KHfG9XWe6A1AjV9sPVOIuGcsM2KZwr/0Z7r04ax9KzJWEYQsI3XgqvCCyTHDG
eN2AqdmXqupWhuWozNn9aJ+oWFQVmqdVAFoce3qGZNvmDQIOaIFVz8LMMYDaqvuY9Ht16VVav3XC
KYNeZa+XSSCoJ3CAyEmCJgAzXemSkkTMNU1ON8GIEsEx13VNsFcuTYpla+eOnr04TvX1h+10/6l7
oVvoecQOSTAFfe6lXVIzc8llXdxu6CA1HQgcM2k81Zmb/js0HPGhoub1mOKkTi1+iUcoDPbELNXq
zKdbI4VKVtOCoXBtXtY2b0ERp7EKnfT/ejGqiwMauqKA1O/GaH4LEwc3Klj3O5KF+uZmoeagzIV9
IFDncnjM1mBHoFEGV3epVb3fpGjIvGBQ0kLPAxmg+T0GhHnVApSSEsAikzM81Ghq4cxSGYrnTbML
v7ZFPuIyxi8YGGf3Q7fZf97jvcR/FpRQmxojY0ZvbX0N5mU0L8nEhvA9YFKTH9y65v4Pwx/fm1Vv
mgz0h09OJ7pDfolN7w4djdYdgkze5aOM+WdTuhrV4wbLM0mW0JlHdUOKEs4ViVdowlabJ1pPMLCZ
QdtCqrzsZJA7ID1XzMxmBKrJ5C0/ydZyqoFYBOI2VSX6/nbHASmgnveLAFQw8BNafLxPJKw4iKBq
SIAMm6Zl5X7xuUsl/BOVet4UkJvKVDUWumdC+pL3wbempb69WtR/LRtd5hiRrH0auSPD8KFPlFox
IxeimKeRWVforkwnnJM6Nizo2PjFyBfUQhVeRA9hFvP8LXYUCLxG46+7qvx2JuOIml2EXi3HcWUO
s93Ib0WyrTC7rk62FGjoIpOEfWxUKVEkuJNCO0+F8guFU7wb7MaXkRMik/ykDJrpGzpL/3zP4ALx
MyX9npsghP7sb+6tGtKTKL/9Q6tQIucFmVTyEJJcRSQlZ/h7hRopOBVUaeYn8D/1KG7AjZ8eszEz
N7Vgc/p+63PgTY58UIfMHaPGnUf+QRQeVgnI3hd0EotCjPWVqRlEx62MYXiMHF6Qc/ZEYBioJ0G2
WwOBH7Auf+Xu8KXnn+yLLkC/T0FpsPITCyLZojXB1le8bqc1YRc/sqjNSIIwhMq9/xohhxRtNzm8
QNl6GC1Zz4SC0XZy+dGZ2YkXJ3qKVnmq0SwackvJwL8nEDNTT/LxNmV5F5l5z68QcQxH2ZdkhpGr
nmmJQvlSpqjbk/GuzDacMZhZOvqGIW4p1tpFWrUTaI0FjQRwE576Bt+fHHOt809cRa7gJc2Q8VWt
EKwWv47+B/89NseQ1BS7avwrXtVKVipmy6yFIX3CvX75qOZYdNshgZjfqBw3ynP/WA0iWHmkpaKD
KQdde9A+AoQeutuMyzMMHNQ7Wm9Sjs0LuRPvKqVrPilF+15neSgil9uxhcmrT7KDfnxnFu86SOAr
DmWsRVMEhcRv6elQcHwoVmzS5irIcHWJ9xOmLcyuTluxOOgkErBxtzs3CiUSGlIRorOtTH2TWRtb
wrhuPHYIRZ3XJIw/ksQ5EXmmHbYzu/ViJv6SSZL6Xz5b1/eC6k4ZSwc4QQh/Sb6lJ2gmQkXIpOCx
h2E6gIjvdJMCgCosm7H0eeKYVHmzHcZpOdXG7Pb6zZAmaHP/VBmQV7M5unUJJTJnCrBD/W6pRk4w
7OGPlr+XEoJG23D3m9Ia+GcfBl4w0bMgLMaOWWxIoQBw11yZpU+/hLJ1KfCgKD1KJDqqimSHz7K0
gE68Sy4v29ybSnddyWDAsppqSJbg/GmEAbm0nS59u2ilZNUGFHHnGjGuoB0g8PFMIimJxrBqJtcs
HKYqlXsYigPT9jSQ6cdgOjdPi7/04g1CaDTNGVm3LvQ/sxp0pCzD8n187lhju45Ze722dlQ2whyk
6FA8ZM7CViHySFhLL38Qsn4LA/nfYbLZj0OmfyoDybirkK/q6Ay6Z8gZeUMA9ySSSTVJkLmkc9vN
RJU1jkaEe38f1FLeToLLLeXxGYu+RHj+D0zK1XYaIaQ6Nv6OxqoNwg0Hh/SFvHRdo47Gy++gkLl2
5FUELexcfGNnP6Du5VTFz6gdnGQsDf7bRIepKdsSsQZ9la3RAt1r7OwfYsxnsjLxVlk7GcYw/F+y
nbBFMSYCnod+sngtAF84XS2KqLIZ2BlJ15EVfTl3DCtMD5+aEF3kNDdqXAqGe1H/JgdLyaYEj40P
Yntt8bQZCYBWDkqKOJCmfmh4V9ccexXtbGV21bzGkxaNAVmW7vKsXpyJSt5SHXiskJLXiA4IBxI9
vHqFSQg0RtxfI2ICupMTBZypTXy2q4j2XJbx4C7mNblj8XIJO/5Th0Spuw9SF7O1VLumXZkivaAZ
JGPgb5dv5t8iOZQJk6m2i7fWzmT/UEKbGF4uqYuTmbAqfoSbbl9yXC/+KyfQB57hqbQuk85/Kgt8
r0QNb1AintOpAqdGQUqT/jPX5LsoCnmV2Kwb4iVmeSNkMbyvQjJcFHQi3PU19U6kYCe94Y3mX94O
4idfYN0YTCvYTE1PQ3NYHKryCNFYpmB7K48PW9YkJelPOnxUcTNUywHaQy5SaojbQXzyerCoEyXj
12sDR6UwAtOKIJbbY48b3Tyx09lhLSBOp1YjUMF1Pp8rSlNcI2y5D1lXP2RoMvk3pfHt8f3o9QMT
yDu/V6DoEcdv5TGB0NgSPmkhbNzPDG8gH+8I4NVN0G2Lv9QcDOS459U0x0g6L4kTZ4rAq6+J+nL/
WbMBmaX7mUB050yit4FpswG9Nf7p8ClC12exloL2koTawtvvPxSCe1zYXWBT39OH5/BfqVFhw9xY
ATPY8eo2MmALTlFM82UOBQ31MBDy/no0JS4rYfxkuy6tKm0BXF6Ioh16UXA0Vi030inlCP8mlSXM
zKa5GabenBTcf9gb7/mHkTUZKfD8kkyF201OfXjY8W5DVgnDzDW0WjCWNqODGXr/Vrq2DaGGrNfE
WRpvAWcb80Y2xEzKUa+z3Efw25CVQMEwrXJ6Q435dcv9tDsfAeWEpZrzkZZCscUigW6zVlIqGDYb
ZYURCMHo9y7cDFRljqMECKMMVL5b60IIrm13F20cmGeLbe9U+eqxNkOAeJ3WElzZ/XUwH8olxSo2
HnzPI7vmXU/X2yk5Wqj22yILImUywkzgMNHut+bZzfOweyyFedSqDMz0HfsVnLNkTkLdJrBEcUy7
N6IS+qsYdUUVoQK7BUO2gi2je1YHm+WnBk3flPcyY6IK2H7lagCkJzPb3Z25e6Z9Iu2GWozB0Z1U
6/87Ne0rp6qpax5IDFP6lW3nQDetH6/7hlDwDnCwGbVY4YtqBLs9QgZUcaBkB+SzxgwaImPV/PJL
l8B5u9IX0rre6zsA/zwdAd6OrP1NlBH/vJl3dXeBrM2grLKyHznzt17BmXgzck/H5lt5LMwVVrSB
5XV6G91Xn0EyrW+wL7WcZFqNl3wamjfbQ7hHq65t2Hq9WzgZVBPIWJ1OYzS9ZsnEs+KwVkc/ngzx
ebmBhd+xcPXOm5wpAjSMUrm1aPDMeOlsHo7s/WgCmOCYRiG2z9AdEL0rEcwkWg59hj6/AeMgugrR
fPBPj/PWNWvBBbk7JNIvplLyLmDjYzfEZp9/Onc/xIQCuejx54+QrCVg/f6YxyM9J3FxzAhR5jmQ
DGwFOr+1+5bl2hoqH9OTUqaFhZ6l8LBva5tWLD9ldcXKhBu3K5eI1ABlCXGBtSLBtTpHC6606je7
8+WKoS/53ovgqIRdV4mQOUDoSTjbcLwEmGG2YPFum5qH7jWhqcpd/JadJNWnLBT7c66mHQepxhlp
8ijcJnykxoI1UUiwxqbA3R6KGnDpgy3EJC47kb2CYrSZzXPO8d1GR2WcoCbvnldw2J1ke54aByXj
dFXOzvLMFk4OIC08fvfltKmtc9+tBKHTokA3NktZ9553qfISxhSDFnpTF7VIMGCn7EN0yqpFaogL
G5Zy8F5cjowBU7SgiYcW6vzlco8UYilZU2NXhPX6qGkMSi2y430YrvTAJX0XPiVsMQGfywn07JiT
K9cBuHa3DEMMsMq/ge4fvryRTKuWuJBqZvnH7wYcaZmq1Yfqp11aadbAKkgFFRBZ7J4UKrQkIlnG
N8+SfEVDOjEitPb82N/hmp6MdCw0qjxpH1yGk2q/LbG4DaL8I5A37w8gpkmy5y10WdaFSyz7fnVq
UnEtVWVIYpzBSdZqGbq8Y/cDyE9LD+YN30oXgxPxK2PyWlLcm5ZFqPEPOCao6XenxUK7qzT+OUMR
THazSnWwh0cKpDQc53vpLBmqHFDg4kHhRj0zmoAgjI/9uOhw7NSZ77xbPEtVweLJcPfCbNsQkMJo
evitwfuhRzCNWR9m55HIkThddh3vzvojS53Hy1nQChsv/zmhzVMK7+D5Y3w/g6JM/dJv/xmUYqjs
OJ0B3vtDB0LFybu0U6K3/fzQt+Mo11WNVKK6NFq585OqgK/q1y3zJufNQOIEaEr8etufeq1VT1Yo
Edr5dTZE91/df4L6fEbuR5yJ4eLxUmFNhKKSncpZws4LIhGZEx+F1oR+/eB2evrsW2TBjdi2bt3P
JFmKxn3If9Xd6HMK2UIrrjhDKhHXDjq3hOH/rkpRQxNjchaHTsvCF57wZQxuBIIPrO5h3BOqCE6D
ejPAz+Ax5z0rQWyEGkc5UIFuKVchj7eImM1Rhzom8xBeooM++E2+yisjROlvycfTbBRgOxGNkYzJ
ToB5g6yWviNczEAv5278goLLZGPka62LqNmeGIqhkIWpQvCFKL5lNwdzFEi4z31MlygQ+kaHAl3m
gKplBrW0poG30CJr5XaoFGYoDvu2jXh3rZ1w94moJBK+zLqFJqAMVKKFLs83QKs+bxN4EMNfU7T2
nEEVmF9JUcu6QfwvI1LzTIf6u4CYX1KYb4TXqavg6Bi+s7IHTQoH+orm3DlU6Ldn+TaA1ckMHePW
kFYI1fZtlZQt24qTTohFr1X/ZBlBsiyUfOuzFfjox/NdJ7FmSCCc6tttxEuq++dz4EYYWHSjtaTW
gDifKJvqIA1kJ93cYdnQ3imCSsBsPqYB53IvSxLtm+NtwFugHP5oyCmTkdUSOne+3CA0UMpjQ7yj
9rsFM57nJWFslTRC06GDReJAOFS4/5yZzlB3R774xohQL+DAu3HQBShGNVyVW4SVEsIU8ZsA3o94
WS5IbfIQ5a06Dbns3DJnKFb9p1GuqcmiGHO5Ejtq7OCcHnmDWyyu2jxYaf8yrD4R/Tzwdl8nyLDI
rVhpBdaEN/hIukOj75u3nTKtEBzG0czWKVYjGysPJehxnHSnV1nDDFmOjZZrpe4Rl4rfUIBl0us5
pWoInnxia+5t4o+HH9Cn/v/kxpYMM8JO7/m+gWkQKWBynVbCZnIJDZk7+1IIkC1AypyQeFyaSFpo
w0CKjav3sTfywfl5XH+l0uXTnJqsGkJI3UvvwE7Pt6hu1haZFnNeibFnlqj6PJ/RDNtWtj0bJblj
RVM9rUydPxGIQDJ0EP4KxrFpmgxqexT4sT0c8ZZ9k1GR9XIv8zZG3EX2EXhuRrlrpeuv7R7a1yzT
+auXoFPmvPTB24ixuYzurc5+XZQyTvDIo6Yj96Si+yI+1RPUe+ARCVQq8IbNb6iWTn5T/AR0Qnyq
rVfXTNfGYz5GoSvSmtdvmnHKuPKTnAdr9SdzqdrXmXoEnclishPo9opFXdqAeP+0YkPZk78Ai3t6
QyT/1i7VeizaTMdBGfL7Awhra1/dufz2wYlySL7praTUgyjI+F/htqu8eJfrdTkwXys5LL3MlPjt
gIOKmfJkJvJ/kKxxZyuf6asU2ZEexXbant6eU0yuoy7Xq89nfhkOku84d7ZXbk2SdcGle/3rZB+U
5+X0FT4hWuqt3dvpXDpgllaNHtfu0+pL6t8bBOTxGhixp7yaP1NuXhemUhLLE86zl31G+LSZxD6h
gCOocXkVEZ3P1pju8QVYgBpaF5x5FNH+bJnnY4AOzEX6TV2V9wsgjRnXjW8lIpuNPkVrCbjGvPCv
5Ib/arhqxlvsFFnoq+72v6qdIvbvDQRKBVoihd7720YdivRYNdJSLtfgRIR/7NcMPc0RToezgJTX
hx0qFDFAJlutppUu7dumNzBspt2po0ZEVh1dms0XekoPmNpdB0SsECqPZsAfC5cWKgjvWXnx9W3b
Bz453GzIAsegJWfe2XQ+xo4Iz2JdaJK8UD8sv0HGFOTKVHaZDHtsOMtYK8VGEW6/DJggTqIwTAqL
WJAG/D2ySBHc4IGNNKJW0MakKf6smJnMl1Jfk0mz5XUDA4Q/S9Vmd4rjSL4UtwSJf9Uj9SyqshUb
Kug5cj1kF2uwn1lgexE6a4++wjnuq+60xRSUTQWEAT6l0ghhrni6j3JZDmoUfroLCv13Tcvd2zAc
5UPv6tRd0Sqbv5AIsPipj/6BSuEPwfMgeXjLfplwdPNoCfLdRNxBE49pDgoI94rsoHV7xNnbwcs6
BsjSwz4k7oJQVT475XU2hxcxGJ9CgDEYb2KmJpIr3iIoJ4JgjU39n7lpCu4Bj9XyCiYeobQq5ryF
xce7Sya/PSSDAodaDJhEGt77XcekEGlWf2MeOo8ODAjOqqcm/X3dGOnkR7n+6HSbNIpyWnWasfGf
b0W6GS2JOnRMHUPMuz38HPApyOVAGH3wA8+xud7eRb4GWbRAkqJBlUOjE4kxVN7PhkV0WFKz2fHa
/heFcIOM9moXhCCXPcc0OrEP86te36GrlVD0iK/s3CNIBCPT90lJc7rWRBHRnU72qF9tmzsu/eMa
izl2eUMwCjzyE86JReK8GQDAwjadFtoyLhh6qP5GtFSMETQlGoHOEJpY25nvk6CcuMDbDLS0LjUC
gSciXaCO2OvJUBdN13ALHedAiWp/QGQMYc7lKlZO9fpBofLwEaJz52D+r+3SDTxqGd5eDcEnxXvh
bgA1aKenUxKGHOH/mSKqDODxfZbO50oYfci4TbobJjMf2et7mo+I1XR2zISz0HXu4k9yfCMyfbio
l2paQeHjAWueSZpVm/FS8te8pC0HWouTgQjbol1PfOhOV056Buyvlj0hGw3jl6zvq/yRjALF653j
QIA9PUvYUk1UUgrB2Gti2wR+A3LmXwvqbfnmnXZhIzo2fbESQQpnGVBMAgjSm83pPK0wrGwQP5B+
t2QcWjX5Sc/yRbXXaxHW60PCf9Sx3USWN4oRw75oPhOQ+bLFx1VsIqpHBFY6dXKtKTdw36cSjuhG
T/2y865RUOKDxIzgw4xn9Z9P0S3FZzxGPvwl+sWOYtsHG38G/Wqd+gEAd9wlh871bhjdiEpejkHt
yGTlyt80wPzbbDYf1QC82Dx/nQogx0HfhVeKKYFohp22w5VTfE+i87IrQHQsnQjB31cq4prOlMPS
K50hFgdxEmaEZ3IOGEgyf78TS7+wXzHN6V5zwGRjB/E3gJj+g22yNUep4j/fe3F+Y+v31kNYRVC2
9KQWfpACyBnuMZHjck8vVyV4cwbjbXabwmjzutNpf8lzY78glfEOlkUrWj1u+3hS2GJV8BtBqbJm
kTLrTpVEYzRl+HBbJqXIfIPAi6F/JqPX/5+5Kqc9Pf1RjAny//7jI0NcfLWkbhWWXhyGYf3OuMn8
wT8wFCTKxFvVt01iyc18zz80SSB4XWkLAShMeQQWpAK+bK0lHGOG+5nUvlxYJNKQ65NSOihW2Ip6
ooUrVzuhXx/LOIrlzvL1TA8PhbQAcKLaN+hf5hdYhR+c9gjxO9jfpXTQZzSVJsKbWa7xal1mfDS6
/5oyNQuHyN1uj5PvLWHgYhGWL54K4pjxCYwUjdN+IbdTbCHj0K8CJOACiNKj1SckiLFnbEeBdGTx
JXfyDD9ntUA1hxz6foOaSLqqLT5hDyHr+zhWKWV3VpEtESxPArkHJE8IB+0EUqCL6XM8dF/Pbjjm
1QPEkqbBnbWk73rSbidSdgAcTIAu18gb6YDb5Twh8ltJ+/Mmk6qhME9rhpaTygDhjnhvcBOtVbfI
aDoXOgNk01gcOdG/TrTohJvRzVVTXUgCQtYFX1bY9w7TTdeTWHLHIOccwkZZvI6+2gqto7rkRNHA
NwlR6oaLzR9stc7AaMtTrZcsHGsuXTRb2m1C2vAENmydOk7OxC2aOhnWBOLaRg6bWK005550Misa
1tmIXjRFmT2eUsHuR0RWIC8udhDtN2jA5z5Ib6VfoIp5UWbxNst7ODD2WjEalI0orADhsZmc1Zgo
FbefQpBapm88CXh3ONG101YIeYhDHFItzt8WFQJfJkY2f4AEqYoPRuacTbcJtlJMULQreVVao3YT
Q/pdfuOnpU38v0hRQyWngo0lmROIWsy9IQLBrvN+z9ChWehuk612E4Osm6dXcfsPlI5HDyvT50Ly
3/IseclUK/l6HAOSfw35kEdr7SvVrrkMZ58cA14cPVzoZU81X/3qW1cSJGobprZr4BuHu4tBX7TA
e1Y0aWRhyfpyzsEEj0PleePL+IYOp4Lxn0mdK9nkzhAl41po6V7fbCMTfgHkKAxZepWjpY2xshb+
bWMiYxGSnClxQR5fotn69KezYtlCoxodLp+lLGYjcDFKVIBtqDfVBsYCwS/JNJv1/tUZoOYqAUez
9a/V1n95ziu/9FfLN2mzb99G1jDLi/VvmIV4+2qkX3wC+4dseqcQouLBcn7dA0yJRk51M13VHG5V
QIF3EDMExhKuryKVwnae+5UHk9WJJhm0RtD8V2fY0i5mgu5wnii2H4U0H5gSZyydI2L8+HVaqlBW
l9+wHhiERaR382Fjpckc8mM9NTHjI5/4uZS/6nizmpEoBLS8iME9w0ya1z2zCtFpzbMXLwElzJd4
36eNkCrX/gZqko2ToeeTg0HFVxdS616hj+yUqby6+XnHE/9gOSKb6n+D58j8Y5KOs+eS1liiSjFn
f1GS390X5H+5oaFgbcYfjzlGK8+Lp6nmGsvMQ+Jw9c2LS6lFzA3SptJNPdVNkmRx/41hbhZ/rSwS
mMIydHUpcOAgXJjL1wGdileyi9enake5CKWkCFqmWKxVfQPljVStuTDWGNGO8x52vZdwrEWU86zo
/bS433YIpDLfuLSemlYlJgcpGIjjrvnInGO6q+/AFmiieQ6igtgInmXgGGkJ4SBfvHmnrZKq5r8c
kPmaT0PWCa2Y2SmOHPxgU5dsmQ3eDg+AgeibbZuBSe9kJDZ28VcSf2E5NxNuuj/hWxBFez90vKC8
VOTuhk5sUlY63M3bx23gwJFxncUeRhSDzH+yJmeUf8u96fMg9Ne1O8ekWl5kISZkP+zxs33yCIbR
xJ07aE7ugESIr8J7HUZoQ7twagmxjQdk/hdyL7XkckfaBbFwkNFIFMgIFB0aRPnvOA4Uibct6FCW
dYcTvL/T6IhpJ3O/05CwORMf6kzuUyogwl8+q6tI69QFd0Zwz2LGPClc4FK7wou9q1USCP6Tz2t1
/jlCi+BiP8SxkMXKo7/ErHceJlyJrKt7YyEV3rT3+SQkZ52DZl05O/OL+XsToeyVIfHrVEzdcVcq
19IhSOfFvZs+Xw443KWMKBPHGFZKVbbR/OzRwuxY9eX4pmMybGLpJqu1/IxBpI7/0pzz4/og/1DP
Wfa2j04aODqsMcojJMFwWVC0tobtDNgtbYSASro1PoRIWOSj4ymZxnqHf5BPVcd3W3tLpQSzwdtA
LdUrX0QNNcyjmTGhc+aZWhw7UyVxMAfFoujB8gA09A1oLUOQVb1eIaBRRg9ZGh6ufulQvFBlNXm7
odoP8YbMZMFjXbyTjF6v7vmifhR0upPhspvu1lftpxFqKliPJGmM66svbzALLJ0ihnUhwdIHpVn0
uGLAmSZBB31ZLBljceVsHR52UwczfIYE26ogovcy0wiMQeor0PrzMZ3Ucay+7L69T4w9NnJePxun
oGeQRhVTi4nO6PUglIyue9bI7dIWBs+lQysDzYe7K0ttckktpXhYMyYMHNC3GsL3W8mWkJQwO1Jl
lN/pNdWmNxGjPcHF3gTeobWQ/1k0wI3A96W/UURMDHWNvCvNKwd/ugUX0eq8zz82S3HrlZDDUNAI
pxMxXCItqwwOrsjMnow05zrZCKWjpYl/pMfYldo8J9u/BVa/Ihvy9YV7scS53VTUmn6KWo4peibm
oOUEize3d44zyYbIjq9auugomj7LXNsUbQ1OGuvxawiz2z+MTgjsWpnpV3hZpId0Q7LmgwPnNyDu
4FSyEiJOXQtc6w9Ip5Eb3bANHd45hapQEgWx1+dFg1ssdP32YBBpjQCfLzxvIPvchvz0AVFUsLVQ
gycs5aIEapoRCezOt95mWv1p2N2uoJ6XmJ3idz09B2Ce3Ozyg2rkSfpneog6Xh2v9Fy51xLZWQzN
+ZfNAnpUrQ5Ts4bYPBFLRink5auRRlBfXL9/+MbF2ECeYj46RWDsqDqtbdUKpXKBb3nJ3iM9YvyP
wVtZHt5IP7cTTACBSYczi2vsverAg14EEKNNr1AOwba2AvLDhPyZLklOTrxCEWUzPJDmONnQFuip
bsIdWKGh6+yC2pX9MJc/C8SoHiK9p/t0xBG3nbaaxlpM0VY7HQebbcd2xW+v+/uWq+7X/iW9tHWQ
jpE9ZoJwryVxvXAxri5Kfbx9Aw9818zyonogcM0wX+GAvpfJUmWlyN3tZ4She849wlssL0ZqByQ8
xp7Bl5b/5d+U1TkTO34bkjlFMZNzsBXaPXHt/JYPwDWX14zsCkVdPzWP+oB9HdWn8PmxRtf5esyb
doKf9FfhqS1joUEjA97PmoLJTDLgsOg+mCwclWjEg14/luztUgd5G2vy/LmqgOhLla7pqz2CGhPe
IMByIFh6zF3ndjSMAiNuFo8EBHuex7eEIHfYE9DVEuXbPBD5wQH9Fjr/Rxk52BunlkwH1IX3IoqK
r5QAixArLxp0L6FkGMEizdq+u1hWJDfXmb6oaiSCDsncTeySm8S2+UMKoTmOhWGkl0tjqUZ0lqoG
7FLUTbxg88dX3iiWSKYrElnKf9RRDAQywXKiguSuPZcsKkXAT9/HkqUlO1KB5eTJpz8oC/R5NSxi
X+OHkSF5LdAwZ2L2Tq52gmZp5ghDrcrz2em3bvxmPYATr0DUAvuu6g3+pDEImOZ8LUvAl69/JFja
wYRGqeeepOyYwW9itds334zdfJd3oX3f8ABlIDcae6alblFBsfuUlIdIgToY8NFO9xDfGYmwOXr+
jw4z7415Vcc47/aYYrqlfwg1tAECGnMtyYnhH0j4MLq7k2EV6cLbsX3KFyzbU1Kuw2YjdUFoUNHN
c43mhFD2/qdVxSPEyDCmw4UbyBxEcVPC3b93aYRX7c3smKKGhvG6mmXFpyWMNZkpLiV8wCy/KZVX
TObwMz/+F2HZW3zS29oU7IdvA//yFIYR1uPe1fvIn7ZwPjaInZbV9CLZ8NM/P4Rtgawl6b0kakHM
9cO6pkoN+8MANaXltxSTeDoh3YJ5vGIuiH8H8tBgxIXFv2bDoflpl+Muk98thLiMH56N7whhQuET
7IoAODZSra2TnlCs2QmqPricNgQiyUruPIXi1jlQwHVJIrF/9Ln0uPgc3NCx2V4GDnHXhavQDgpr
JxxnAvKxOF8p+decpfytaCfNlBJt0kRGG71ljz0mx9BpVSr7w2ku67ZbDcHV/kHMFGiwqMTaoCME
B+hezmOCdR1u92IwZMUUqs9vo81FdnW/p8qj69RrIFX0Q4t1ex+BsBgrkJTDKwaAH9P+4H321WMA
gBHdUgJPdEm1XErJyxAQN2AbRhPdwge7w3k1lAfziCQPB3RP+zdxVMvKMPruyNliQq2WSgeiQ7wI
vhM/60nN11acC40Gu7ExtgG4yBAhE1okwRyEf07vhy/jqILnlpIes7G7s5Sz1Be22tgea+CZYoa+
qUqXFrx5+mMxyNosTqUA6qqUe/8pSMdJFVNZVCpBrx94fqXxnFURjQNm8E2m5L2Qsd4uiFZpnK6E
xt+rO8YwofHEjo6geNEEL85oycMivo/jaNeHr3rHcNXTEEc7PX1uMxIytpoY/hUCZ9P177bRf2Cx
PqdSRP7bS/nT5gazfO1SXb9y/HbSoXvYgi7gQSLWcAdrO03VCQL7FqiFOEQORpzQ0TEcUhkWgg2H
Byoli7qMVMuasQAYAt/brLVyP9rKP/8fuDW/egQwxe8TKPnPf13b3gcYZIV47BTQtNvEpppZp4dx
JbF15ILucmz3PSG9r7yfDRHfnbqpeZaYTjV0nGniqFefPofNV5zd7U+FYgKiUs20Q4eogVAYT/yl
3A0bBcuB2eP9e9zHKN9amiRsWE1uXEaP+r3NbnAa31rQfCEJbDJLq8SlL4GOAIbwumcvnCNOMW1M
rLyfufbARCRg5YRuW6lVFwcGHRrjUuandC3oPQlSMTHWtNhadyFWJbuFIrW77XHdczyrH1CxHPvs
clCLbFME9x9nudOg2eFQLdGRiHOFJX57L0Omhdq154lutQ64+OIeYt6pFRdo2LIMYzSuuUg59X1m
Wiqz//Ex9dnjBwq0i5D+upHfXK8wpMxm3DNWkmpWz7yjFTv788ogctKZmBAOO2S7WpQTwSv1H3NR
nhtV/TIIBbpnqThwGJ5QjePKKrNO5PIQ3o6HLsPAbr5PbVFWf7Ghk0wUSTu0Z98xtrb7GS1iHOyp
1y2JMOWSbmL4QOE/P00BN+3N+jpGUWkOXbreaeNNmtClLlYjA5/2bO5Q7AEWhF9U+O9LNsxXInSa
iOS/LtI+XK5uMtQbz6DOxQgqawj+VmT+krbl1fATxsfkyfC5Jtq+psc5uWewARpS8tSnI4TCo4M+
BVCfiwU1CGqYSDWSR/xYi66MPAtGMhpsj/L5/Ywwddi0e5eK26fu7LoHXJIbWnRv/LVGM5sd3gA3
CQYR0B0THIkwirppZMa34AfvwsrmcubMKpFJlide/enWApEx1BRKiSaoa1yelbCz2bn0s666rkd4
tmbua1Ge5WOkZvwNjJyB0aJqTTeiyH6oKGWtQB1FsnmCqybzikyvbxGtIEBWI9giuC2hQ6kyUkhH
gRRmqIpR2QL2qA8C6EglgBIO6eh5GztQMIA2kL+LX3GOQPGfSJU1S4CAvmMsq15tyoxX5/qcUG2A
iWUy1SIjYZZG+CegI2H1bOC7hG+pMTmNDpfIhLEjPIR0BNQKi3yTJK1pi5v9lceSpgDNeJTedL5k
P4sUzw9JBoc1Ph/v9Vi7BmC6ERrM6o2zmuaNvOmqPMAmfgS5au/CIfoqpzKBhb3orX5yaX1omzw6
BJWtDuW8aJmr/GTLcCeLTKYwWwmEEJdtv1j3copbbpdAsr2iLx2Vs8Sz4cFyFQ2AoVbVDMK9F1Jv
4pCVizQe3+xyGKmYAKEqQkuW6hGek29SEWH2hmkeavNgegTpW4Hr/8i9GoMSmXzDLPSjdq4U9Eqf
6k06+yACElnwVEWYKOqcexcVdKcWxruTSLhfTGYdUCXYk9A53fub2C33TJAVwPo6Ot0FlMSGzrp4
cYD06tXSYSJfMiOk8rc3nQvfluwrWgF1CWZPQ4+eMGtuTGuptXz1/9h5VDxvfHffy40+DPVNxzT8
O1BESzIou5IVjK7yFsNxsPPE0GgU1dcTiF4VKEmhTuGk2S+AVVx02AKrI/WUrKGfNPob4pavsvY8
eMvqRDHibpSwGmTFr0kkTx+S/foVw2txwKIhE+Uo6idrUSn6G3zYS7jw615815mgNfeGECUTM3AX
U0Ny8VgKoc2ExE/3y1KYd/gLTmYXO3r8Ca2Unat3I8gHj8L24A/PVY6sy/fTn27833RsGahqMuYk
DFG5cF11xVix4+p7ccKa0yLcO0/UcqZ2hQlm0MHrLWSUqRT0OFfA+9RwyQsJQVW+1UM8iPmnULZ0
Qu6+u9T9aJ78Mvw1qNhK5VW/cRjIPNlOo9uNwnpODJ7aPpQjMDzqfdn9737PU8lZPJ5+DhyXloGQ
+wdSdyv03f1soj9XSi1jx6SMNoNLjl/pxlmw+Tn5ZXO+KexDg9WenOLWGLfXdHxJ+70Zu9avEjAo
rmpd3Twd62k7LTM5Sszs92JinaSIeqCFvvkI/vr3FXFyphjCt3EvpPIMHzKvereIKzx6tlNOOLqn
JPtMc4yeZzm0OUgW0XfR/M7wPn7n0EIdPMEISh8gH9pQbYUYnb0086IAWeqiL7322wu2qiDwCJ5v
wAsvglPSQr9keIqP95pAbibD5aFOcRj0auxf0oiKrPP9bDF/gKyPZR6pMDwfohnKwQrXfIdHmcJ+
vLCLrU+v5pjLNCh+TDXLjgy7yetdO73QZRVOYdm7zx6Q/h5HXnDNlvsoOuLpv+6b48rxLzWaSQgF
jOOGwyCzC71SG2/dRWe49rZedSzymcN1TuYXUKfuZR0NFfFfTuNM+F6jBKgpbOuFqT1uA0bnBcY6
Wa3eqDNyZ8ukHgtT5JqDxTftb5sk3JmLnMY1fFhizpvMi9EQIbaBiGlZA09VC7p36sYASiHDNZ/p
ECtAqhtjtwxpycDC2qqddcarZvcDlYID6g+eXsJbEQB1rgnIdAjfemX7Fa9mpk/K4+wYfkX5oXxA
Rs9PaaEzzao7Qh7UWf0hlxqBi2xeV0TzHX7BBiMXhl6NwVi1SeidThaxyk6/UgRWhwDtRCxzX+JK
dlG+1kGc0JkzMDND9kW+2p1QBYd+O02GlEkGo1qQ7pL8Qa+hgrLdnTzAclr57YQpAEzS5T3A+SSp
+pzGUAF6d1YJpElhn8/CzgjEaQcnMOqbopLvy2HwkR/IRnLFx9e2Y8ZjowJQGcmGkQWTKBnw8jG+
vpFzUYqfRC1vjcoaIZjwdvh44FVvPtqJGV140q+/z166guZHqRfbHodFFb5WQQVeUit8QLOn21kl
xj+GpR5pSeJTT4K9evooJ5OOXgZ9Yo181GxE/gTrzWGunh0evtCFnOzRKY1O6vkQKNTpeFXNMZ21
VnFwPPPzFrlihuyyzkVK5T19D7AsteDgR6fIc7hXPRk+zzHUmZyw12VoDjGuvGUO3P5ePVw8L0x+
ySpXQ/yeqS8rRYusS0oyICE3TT+OujzrYUq91wTgx752wcxOwRZZApXnhK+dRooww/qJvDjYABvE
kKjc6c64qgZfRuRLLChE0W3Ob40OKb8HJPWGYKjtXzWS7A++v5BWsB162nTIDTFcXGlF+2tzY3yE
9NVyOTCfMV9QkqNIikDMKYBIeAretAyy0pEJOcvZ+imE5MgkzXIhUpfPc9/xjE5KrCa9gAPAXLQU
bnLQs9PgMw4QYF6hIKEl4ufVTZKcTWSd93a1ADluFKd6a6c3oAnGVoZ0zjqHgrlPx44xSYjT0jNt
uwG1MYUggDhIBROb+4EXnT7VWhfnpe//sKXsqggMqug5VY4V9EW9DG39lcmRrBrl0YaegnKUsvHP
fnHqAzeZ46bkwTpNSKQL2nIjxavhFnd87W8A+89kCRC7H+q0SGvCZwE1e5Iuqk6sv8jIrTg48xC+
0ehmgI91vvJpzzYGo1FeUanzHehC4/sgCaAZQUiPULySF6KQ9sww/edg+i53iqBK+OyXXcNLGL3W
406Bz7xFTbUaT1a57yciwm9XCaRdTrnI97qfOTscYrayiZ+e4Bb0MZ9QAKikeFw3/6mdcr5eXRru
QxuJfa4EVzUapliomvvVLhD+txgc1URpv9vizVnRIhXDjOPybPiIAY9pOfuW2NJGUqaJI18VQEhr
LjBS2+fBG3+bEc4T+7A0o9eP/AhmZh9RtSFV1xhTlNPHe2pNu3tkgBSBEB/qoE0SaT7jpttI0RnJ
g475LR+CC2LJYsfufFEIbUm3iA6ebwYbMD0vJpAfgZQv0mqb6IG1MO8TzcfoT/Qq37+y86U/G3uT
8tTFhnBfi8yTXOLIZpOONjussYVHWFW/dCdyfZ6l5CcSJZZlmLrGUDe8p4gMymHH+oZLZ/wOYCsc
SvU7xvZ9MtJx62+wIZhdQ16rYZTNvZX/Bgy7FV1CBQbGZqwoscOyc3jw6E8M9/+NX8JkE+vA2YZD
z90JuWg/zY52144iiE1/YsEYaklYiOvQ6/1COgf/yBE1qLsaIMSTFq0VnknDJbJAu9vUbk4O6Q2t
fVqvuncnar/kGv7EDITQjBIrdpc1D1ARyOdTCOBXdB7TMlwkfUD74q0gJxOdFh3S7pqv43XR5Wqt
cU8BA5AgRrYxihE2WiHFhbagQpQq97zw8M97Jv7MUHA4QB9TTmLiMSC5hmwW/lOALfCGDTiDtH4e
pF8segx3UKaiPNrJ7IjFaJM7BaHfY2t2A8GJvWK4cYzfDfbnW96IBrLNpRUROsr/CRoTUqgsQmkQ
7mnb4+g/07xw38jVtpe8CnBgw9YMlzNUmeKIOlAMMZ7hR5OQ3pOXq9olTBAWCbnR8biBuJPTGY3n
Bqjg1HnsZ5K5vPRWxCsQHzbS9e9rKw4jCC1HUSuh3PNYZYBdXmobkyFXv5oX49SSTJFYHBSHVm4T
5/ps8HyXB+wrQ8VhpuwjQUPBEL6tXtTLRM6Sjvu7j/043Du1elE1+3CP9900IOd4k7PpKfYjKuVp
KYS/TVVJOOSfav1kYzWUIWWgnlIgk3war/NnWzBnrq7i4VfgjK9nApImF+pTezeNLJyaOFEEUzq7
eXoFspBZ0v5VzO3VtLShoMRqzdcvcAleoH7J7n6Ra+aJGfDfLyynLGWAhKztCE+ASYsD5l2pcdR7
928YWYbv9QwI9v+fcANfsBa7CIs/T2kDkT2dRy3G8NtiQKMK8gWkPFvoKyUCNOwNna/sq0J+nVVV
YYcArcss6z631srzH7h96EP81XtV2lzhKUAQhLqJMr9mQPexT+oGTGLvWaDZvQpNYkIGcNFi56z/
K6/n69YI7UX5Wr+GfVf2GVeymILBB1wRy3QbHXkfQ7qsISBVxt6ljAYpKJjBQ00rW+QxF5CA29st
1gJ7NDurVENx0fmpZQhFfFbhz/jIr0AYNxURTPAGJocxMgu14Wh0PYON1V7wPAIXIRofjcW0MP0/
Ch9juKFEvFAwyYiirrywH+wQNfas/Oqw6YGLIH08cdrxdcx0b9sbQ16mk5YZ8awxQQcUfCWtvQ/e
HTkAb4m6lEESG87YkZMuhT1eJXzHXnHRM/3BYUwp4YHQeWknDMohRQtF68hjcv4JH5zib/A1GADa
fvpdVpLobly2vaX5tXrv1SYTVSi/ACQwjCHOhJmSYzssfP31HisCZsmb0ACQoLYGh04dbLMpESlb
jqXEFI11VvLnhNdhReCUbYTSusJjwHtf2Uw3kZ/NsI7CW/ekLgkKfn7W5KSRpVwk8CLiAId9sDVf
w+aZUCPsJKAGG4sXx+S0fcDozfUEAHhKYIofFJgqt+MsE/pMGqSG484aizBdvfsu1Z7oPD9P6j6E
y0QLfWeHKOcH+AnWtGArm2wzU52sUnBZD/orW9rzQnS/JYK7u7k+OcmfLiHH0VvdzDA80fYIqW4S
xRIdZY/WJeE2LIrjHLAM6x790bTsmHkjVVifB+Wxs8Qw62ZRMewlc39G7qObISx6r3cjWJw3c5t0
/vuoQFP/7hXhFL7DXux3xRnzM786/qRVbFoX72DC3nMkY8KHGKYrGoujhckOvzbtLEJmBxyeOwKy
Fg1QJNoP8svU6yYhOMnBeBZ2lQgSo9UAHPCFgSMMz08I86nF9uslluIfMBhYG3PkddL9DyP8N3ml
9zQUA7UFoAVRu2JEXW+lLnQ44XPE03mNKeuoB3x3INCAlm2wXd5eI9as9KNMi6MDgL23N5JvizqH
7hqG8fFMfKbqwVxQTWsdnH0bp4iIPioxwVsLiFwGf0LWFysiytu4nBdcrZImHVxtMPvOUB7Ixrvg
ldw9tZ3REY5m/SNZxeiIVHRrbh4cIatmwmgiSmXe1cmYleOpNSL+m+uniJCZXE9ImtudRLA3oxOx
Rgma99MuXN7zlo33LZVnENsPOoWA8j/OGkehG2QQMUsI7Q1iycFunehab0WsGqPtui5v4YjSQ9xW
1N/agYIHfgN5Uf/QokkhLfnMprmezkk/Z30kzTFuRztHGEhNtTrWeKuUG3QRrxcaGD9OGCPOk4J5
lhWn7DrmMTiv+4FiYTvOMAYzYcY493bkrt3PtLSdQ+3FwU4nZsGb3rN9IbzbC3gemBYCW3LYXhDj
/2/iBCBZUYV3Suhor+Dp9eMWIqwgy05tQYSL9oeRTRY0ayLlM5doFnxgtGKaJSS47f/8OksJj6zi
O+u8thVaVKcH7C+i1KByhI3SYH792K170JzwnFRnEiMLQpJ/NSnoKTLsIa+SXz7RPwdr9b+btJub
6NfLGNpKv24BR9jZ45AK5KgwKSotDU9G4Q7DPsVHEcWMLw5+A1n8JVVAXIfHua20BV09TB9cGO6p
8SWd0pwZupcEXUdVMiTuWwsHQORyWVkky8xoSm/ZeOALaKCD9r8q07m+Bd1bP5XkuBHqjIfY6ybp
f7dydmeHjpoAgDlk3phPmtOi7KdyXOQmn7jVcH9nYsp8suVwXTnTNUk+AA5dd40noxiO2ZFngz7K
9dM02XHEdXbkdf4xn/8TXcmn7Gx3SeYeap0bg15z6FdK7wyLY/68Xrs2rQo8ZFs+p7EJvK/nX9Zs
4IFOTGjNzAQe4GdLQBv0duyChJVBCJW6SRKBHtbWCR+70IIJ9c3VvKHVxw5upoq73mTi0I9WNwzW
+sPkSCblNU2qBayWGZLFK3on1hyKiuYJjiJhx8Ln78AwzScMyyEkMxGFUB+bXQuP3qffNhi2CI6x
fEMOl5Y7WWfkJZKCqpLZbC6nsDhvKy7ikfs3183Bx6sSNmJGtek5ZlzyoNI7x/xBJiDrC4MS56wR
uzXGHI5MIphlmafHam+PIjpRudkvcdkDaSzW6wnJ2oHK92S/PjhrvM6y/Vux80ZLr2xoGItvk5hv
6HxddPeYiguEMOQzgV5EHas/dIztNyOwuMPnNuqAW8YzWr8l2/lBJZBhfoWtIdq/li6QmYnjduaX
TvUW4hPt4SFfEiUhv/G2rB1AsccRDps+ftVtCtTcHfgQb52a7bEqF7BDBpISXCoxOu/2BueWW4xf
F0/SnoDaMihYd1IJL6xsYXpppT1R7XCMYuZo+t7aeR82TZrb7Dy3icg81PGvDFurOjSATjI/wm1a
6xjP8WzvnGOTi1j6IuOSK0YPMnJX0WG/IF16e1iu8Ied0MFJH9xfCK31mvHV7AQB7UpC8YreCFrJ
GACdThl7JXG2VvVa4NxXpFLInd8aJdwMR5SB/MvAfSUtxRT/rvFpFj+QsjkrKbpG5FD2SbXF6MtG
5eQFx81Y1+dcwKNnqZ2lW3jN4lTnMxMuSNr9k2UmJMMtvl21S9n4Eacxk3v8Hn9KWLzmhjhDm6wY
D/8RyKvee2/TLHm+Ga5IDf24eZWryZGvsJSnAKvRMHnNV8zmiua+q4JXb2YgJpdoSQgpRHMnDagc
cs41FyJxqMnQlI45VsoWZgj9bSRZxUglRvL7PgJG4yKUgdJ+Odc2AAGzw/tpXm4dorisa2tUOnGz
hm5JDF+CK1DBDEgsFdRWmCeHT3ZceXr0xW81m1m2saCbcquL73n2wboyfOptJ9jeLijMoYWOdL+L
MwZl15I+/y86Q2NAXF9WTyTzNqGhz0VAnLX3CELRGd9PhZeIQws02sEBzJ3qFtDMLSvsCAed1+5H
7czfxn3iWuEfkKvhnMGzm6I83tAzKqS4y0POCdKXuKVba7Fmt+oxBePxtUfrCnuAAP7NHO73cJwt
xhe07iNTbyZRPMaoq+Ur9CtM9AFMwWhvLD8x+xIhOtFsCJFNPNmh5vgq0zH19cghj6Ka7uGMAUIe
VZISZ2inggrzkn3AoQpzXtXnfeOBRmaYCydsJrQI1/+kp5DbsgjpUIJ1DH2/vDl0XmfLjIcAM/dX
bMRKijUbOka7h14wDLHSxTiDPeZdaol/LJ54fOSOr/58gXxFYHVAZayA++l9gAoQHf49LLCTazKA
1AklDzjQse47AYcbsbzxENx82XVFpG1gTz1WqGjeiSWmYey9Ag7rg4lW6YxcPHv8b0WHiBeHXS6T
g6JVqyTqsHpl5faVQAFjwaoz1Z/zBvCufYahJYdZ27hCGHWB6FVBnignwnf0MPy/Vv/73jTLkbZL
vtU009AmKT7D65/Jrdql8Pp/2llzBlhDmEV3lEBu98XRKeWMxc8Jr8Y7bSphjDf0ofpv3RPF0vnz
mc07JINTw/v0AZ1mR3R7M+PsAr9hYCFc0HIxRzz0uvR1fy8p2dltJyFtKikK3dcP+8b9W7rIXf69
B88wdF+OAZLuFIUbtG/OqfPnQZqIheG5XCwzjq9BM2Pr7T1nobareVw3BQAGmFk9/hUpGtPi1CBd
xVP43i7uoew9va/zUXTT32PlO+tbo/VAW0ljckvKlv3AqtyNMhPuec1wzXs39b8XdkBVqAmuysmb
Z5C5O1ry8Bv9FP9i0xy/Nt9H52HQ6yydfXXZfaVSRJKClEbTp45WvTy79cYW+p8qyw5YgXBwBXXn
j77nrQWQAj0N3ax8TBgvWLQmeN1X0BwUXTAe/oWlI/vv2EqfGZZBkQ02Y7lN85eBMyAFKZI8qTyX
0MJBPSBOnCVc0IhDUR/S6EU5aRqHCZ0w8jqRs7vBoG7GuRa+/THd/dsqZYlb79gXV8Kn4qWlMSBs
LFuZzTeLhhMap3QdZ7XSQOm6AUgk/94aW+86H0zGs7neI7/rX3FHIGJAoYyMLnge82tUiv/hgJFs
UXEUncHDSI7FMH3MZBfwtMgDHI0o0SnfTz0GebfH0WAdGx8LJwsguF8kvXyPjUlRVu+ETYNjzSGg
2FZVrFmDSSKMpuQFN5kb5vSdyLtz6urmyoUh19I3bH9OYgjbCmGi+WO+V0bzZKxrl8MESm24ooWU
tA3iFmY9Nsb/bmeD4CVyEGSf6ILWykXB9zi+9duAYeoMklzjYE+iEjIN72KQX3uG3Wh3PoebB8iC
TrR02JKagvTimA86TBc1kT90FMqNLKiiINisEOh/YhoqLYI/oUaN3uJIbAJYB4YGXU+Ui9vLSYOj
mVAAZwdGr+PTjzxU5Y9qJoHK0nuf/VQIqcMGjpfXlCartIIv082flu4g1VzeJB+tES/GMp3IN+RV
T1ecres6tgGHAi9sZfGzeW8yD0poLLIQ0h6XA0zlOChyZNS3pmkY6Uwv5OQcD3a+eMslitlLlSQ6
5LH92pyVuLdLTa6dOpLo0g6hhDycQe1dJnhLPcybtc6pNDu2vae22+uG1INV4Jeo/KdZyrmDDrVq
o1reXIDzjmamZ2431ksmrWFfdNbcrPcx4u9G/ZS2Wu/WDhOFvdabZansmk0yFoBTpCtDe3zecizF
xteD882J7HxesBLC4deg3DrsM+rfLv32uxBdBz3fBQHAoSTPEsTBn51Uyp2F6F10KRqE06tMeeE2
o8lxBKE1KiOkyiqKn73NRGQ0R49md3DePbJY35egQctlXNH3kBPocpUdF7DzND3yPoaErqRMpKZb
rngL7u6sjxZA7tFD/gMEo+v2L2nqCsujimTwBIuvFHK1txWHmk4SGhThhqDNKvCO3zOYZM2QERhL
RaS6Ixx7p3dOJttfXSidlFGuJZu0u8GwJB8QnMGuzHBepZHOmbzGLIDCkNPZmlgX3JcaDS09enbz
TpjzYAgyrs6o6ygKO7M4eJOe/ZXWpCim3kChxlki7DLfPAOOJ3/RdVI6/rZDjsB2EUaF2n1JvYD3
aTRO78c45Rbk1M+lky+fXnH+lUAXjLQaP/a3NttWnfMQZmIUsW48uZ36yeZTc4uBzv2PWbyY+IvX
UM/LZE1pMltlU4++R55SHXaqtZpLMgkxC4UyI8zr8uHD2BbK4SlqDAG6QfQLMHQS7NGbN/9k8zIf
E9pMEOuqBZB1TyAjoHnhud/ywSl62ghEfMMfWZvwGVMhUM6drByEuoZG0Ue4+ZwXW4UCDJb8edaL
dLAcOTYOwUkac03e6ck3+rdnFb3wdDMYZpAFTXwqBEblg4dlff1OEpJb+mPUZwLbJaOb0pu+nUb4
khMBdUm7F64r9ceGsxmTw260wYpTOYVcrD76/2DFKcHuSr6H5FvCf6D7AQinBhpo21blQcg137Yh
2vUwDJCItjs0K1GAqBkZA9S7cphTHZvapFWO2lGOie9zQH7EFH5K1QI8bng6k7G5DBgqMGKpXSHu
ch8yU7N6MqOeWU6+/N2izzklQ6R8KIeUO+zH4OrMHgN0v/rtFqXAfhBTc56v9ZrbEyVKW8vA9K2b
QiP3aoGrE+1g7tp8wZvlrYl8b+s9bOJiP0DTpjI+kev5d44VSitOHKs5JmOhSNpWZM2l11KOAIUq
yu4uXHdrV6m/y7nIECIZ2Aau88wDnzWT3YzhcRpkxfLes31/u7R8qfb7hwPsnDU3p5ErlxcFZV/6
T+t1t4vuCNTg6O2Em2Rl5HHv3YuyLXaX9lL5EM7N2zwJ8hVF+9xk8hwJPC4CFecZsrpaql3rRCMe
GFR6RX1UdSY4wptFc/YRT9Z2l+RGSgbg6VmvBttWt3huX0DO2AlaNVfzTzYEuXWDvOJZLw3/Mycp
2m4e383BvrQlOdoTGCi3T8lQhPZNKvXje8wwkBo6vhxZvRrhtX00azqpjoWcUd3yf02fq0cfbpfJ
VfiS1qzSOVD6q0NWI70nsGTLRl8LXTCBf9BXXbibpEq9sKg8te1n3KTalSZhhtQXqSDG4SerR0Kz
G0aa14amFNQ/W0FTQ1Q9GmTaLpN8fzYNA0RfYkWW6qhrvWs3hIL7LkH2WcYZ6+cx6P1sqo4rKWEV
fSPjqCVdLgyLJPlL0jwv5oe3u5uQZTmJDfWf29gYtKvoC0uqFXJfoTPkPfpjkRgRFH+eEKlaylgB
aZbrOnLIdQWhGqu1xVHyFCrzJq565t9wq5peX9bezHKLsuooGYgrb/M4h4ENShD7+xddqg+LniGB
/nFV3a/Tx5NBr1ECGhCpUbkPGo7fn5gOLK5yDVXgXStUYoF4j7zDS7I2n6rpPSfplbE0xKtgR3HV
lhlyRaA4AaAbgNvMdyoGpVhbEEUi0MDCdEQ4qiFmQONwnFdg9neqMrV1ZpQT0ofhqA/XRii+QsDR
TBro1ef+5m+yhZZFvIq1B8jSUrmFeMrqyG7hFqjMcPMkZEXNpTHn7jX5r7Q33ONpVocnq1AVlL2k
mNXQ2StgJSkG1G71Ce75dUlVI4yDi0L6SDS2752HrXPjuxg9dTGTCOMq9PnECze8CjWFjuOYiyQ7
trVfhIjEH4Vr6cx95vhrlFdnWyzEqT9F42WSa7RDW6zxQNEHn1cKUVo4l/81JQOjxYjf8wF46iRc
EsosDa9Md7eDeCZMvSedf7oeAvBD+MyoUvLkBbj0gKPVru3PGJx8v7tDeHSL1t6aH1nfILCbTBI9
eIHRcvWnq9f4KFBFXzb6CeYHaANh5zrhdNr+jAE6K9bs6JAFA73OlW+ifD2mYbtSQT/OGVR/nBhT
8GO4aNxI2RUFhq3k7EYcx0q52+lfV9jYxtUGbLZZMOXZCgq/mvRS9OUNF3chndf90aLNRvGe+93T
2a67ZCISFcUqTV4mIJgux67WIN9Xf761xiS2GTNF9DwnoQ9aqRdNCODayJpd0k5bbHd05p6OiQ1h
AuICxvdUeCmRW3jQ6YyFu/O98YLiGkHDeSEfOeMJlUMq1Aey0xvMM8qY/WNV1Dz7GvOJqoTxZcw/
d11/AEmOjn/Kxfd+oz9akzLYJZlfOW/gBpT4eH+SbePCdGfsb77+7CUayjCW+afQH4euyXN9U2ja
M9iYaFltskCALPsmiJcl5gYFv3T3w590J0ghZHeiGHPI5DjKxTK2Cpn6Gmhj+ii5EushUFb9XVnm
sgAwVrAESxFCqIW1oz0LRXNg293ASuy+4IQ4l11UUACpALkw6FHBezzcMu91oV/1Ozr8yxTlW3lf
t5Y1gS01k6S81x5NLhZH86cu3nG1IYCi9h8Z4aqFMH9ebSGDZuNPsTFowHdyHTEVxqt1jvKWRQZr
A0f5ffbZ5t3VMUVJyqTaSBRTdBhXJIPHAylmBhIseO++6oHKJjxglVmNlga1/QHirqMNJf4KMvqx
WR7TWedoVMY2u7p1F0Fj22cQnu6MqVi/IcP8XtmPc1kFxksp/El9V1/LLjs7MqNJw3otOBzI3ccj
4EDY4SaJOBIKW+gFy80l9gRkp4wPhUD3Ggniv5RjCx+7PUIFO+sR/5QqBm0OYuyc/n6RmAFt7/Et
hSL1T1XLFMDlAh6QrjJAMUrATgnKoxycR4V7VYyvPIbekhKjdEgW2yMnIu2QRENFN2Me1VxLJwEu
KBh/xeGCOS7DNvuTcmFkAflveGMqUpYBgPXN2Xy4cGAM8Ehb1/QHVwRPu7pqFKDVCNrGFql+RFOA
Wu3baVW5nwTul8sMaY3s1bR+othWgNO5OodoCZRg6Rtga95kz9hvO1yStTeh2TCRHc8/p0E8dzwu
rkCJms9U5tR/vToBVRmDm3K8t8gHxhqA+oA+gCNby2gRp3hR65LsNksz4Kqun0bfsSWGUGKB/Lqs
VsfXq4n/4oy/x8lB4at35S5oAuAmZvi4XMHH30jwJNpnJxxihTXWv82sRfG0++dJ6MCep1/PtT2G
j/WSMFoATW0Jaek3DkARKGLyvwje0Wv/xrRCiuYUfunTF7cXeleA+DOvbY04nf4bJLNDvvmtAkbA
UjOWjB6Q0RtbVT+AvOvvfHvVNCr96HOLIw7874hyD7nMSHIlZzzZaN2KG2ganXReprlAnDtzgFEu
YeRFkNKR+tbhIsv7biuszFpA/By720hF+WJMSglosqo1R3l7IW0r0yKlaMtEaaEJG8qPavb6PLNg
X1lJFq75iwvx9wvcGSHFGw1ZfYyJU1qtm5+SH27Ff2cweahgfVMU8WGxNEF2FQuClSgn3rv9TC+g
PHHNO5hPLjbIWnB0PVvia0c6hlNnA4Z86E6Fpb+JLaHOSR5OQpbPYlRzD0VPFTOHdU+9DquHcrMU
FaIjydm9zvdX/fdzQ2DtAlae71EQYhOQu1pNYHERd04ru3kRy0HXDtm2ssoAN83UGL090YlP5bUQ
3m5d41Rin2ossCPsQzpq+ZOP8ZhqM7uUDdgQoUAY0cC/OZ6yVzN+NOvHG7QV7dVruoJCWVsG9034
ZkkUN9UO5pqWJg9jQmPRSi1XLDVv13q2XNuaCRbNrw+scZqBeRCsri3TGXa3qIWmRHvCbqHUTO2q
4kNjvg6Hfn75CcHZj9XTcVbwbasc2d0+fLmouwmibK6EISRlxshQ6fvzE/dhRWQ+bgIfqoLsROk/
OamIaxCkju3jcGToFw64AzjD/l61N4WOyLrNtl83j52HnBrpXnlXTIjscWyxgXzCQbsH+uIV2Z8D
R3l64eYejDlq53SpJWLK9bCtVkCatpjiHhIjJJxqxyH2d6aKhnNzV6qYwySE00xiwYHdqYbwqMf3
2Z8DUFR80C0nybq8WEPNfr9tWMqLiJ65011A//RW0OcaiQiWQCx890OHS+CUFp/xjCG2F3+Bcjy0
gJDrR4Ds+e+ahaNvUO0rSXHFeTaTx2E1uIgkXeTOiM0jdV8WXaahzYLV0NiV5z7NEormefWcGgEj
oznYcOLT5q/HAnYYWB7be6roNzBOrs9xJOjHMA2B4Sg5Mqx/fEaC7v4YFQudiVDkj+4pOcVMsoom
SeakOwY8GWTsClgEirzjZnViL/wV1DSkJf+oOTc979y8VNV3A/cLKbpRcM6tDORPuvz7C0lo1Ej2
fj4nhSUq87Us4tpE2IdjcV+SQlqgwfxfsDi94fU68C7gSuMorcTUu26A/hGArsNPPSnMleIFQ5nq
w/z/iQhjfUhaZx/EnxVNtG0i8qxH8zUI7wk6NPofwRCb84YZ8rdqXTgcVQujQLySSr/Tbhc6iZ9d
WctQPak0pkYuUKE2G0bylfszrkNSXvpCwykmYAGaMccA9QVL9KwnvBjrL5qHj+FrKfvDaw6H2R8F
rw0T+MXShEZ4ryJEPOx5wlWhpGszIXs/mxOdKrwF016OA55f81IkMbo1u3S/ceeJGJln9B1Tf/Q7
qCbHwkMeEPuHSkG3zSliNTMUKED/Gbp8ZsUVGJE3ft9CwPgYI7Xdsi4MU/9sGXx24ounf0G7zSx1
yXlqR8A4LYa91ReQtTmmwnXP27/DO/sIk9IX9wijuEp4/QCZq+hfyIw0zXItHXn+MRbPuAQW9Zu1
6OoMUpn+CxW7eVHPt4lvMZAEeWf+dvpdn3CxrNFtb9gmdQKnonad5a6ubsoR3wPHYlB9J9ZHELgr
zb1eR20w+p35uBtfX7fufk28lZ/H1u4XpkGlzGGu7IDT71Rg4IJuMn2epieX34Ve3F5wkkaqNrWv
wEVSfN1WCdWa+qkUCID3EEsCbEpW80lEahIs8yvQCEQSDq48yQ5nqXMkN0Ciqje6qeXC8TFv4eJm
xMRS8bAvpyD3EAj8AFPPmrLxDpqHivUd3M+1Laa9Kbel/ABOIUzijlXLSzuOrVu+JcSPNVvrOlO4
aqilm7NsGRG+hkyl53Tgj2KIlaaFtUrpqP6kSxrFocW+KzeqkR+sX16OiV+pmeCh1P9A1Strh72E
zmDfQ0EUt30r3pmqiziJQ//Q7h8txVQpYZCfQ7LzcKXXAn4lvhHRw5+wjntajQDOs+6YGdfos+T3
jrNadZT8rDXSh3IgtOe560WqYmX/jw++iqgARwjrGf2wxfqNwfHPFeCmPFUKpAFCC7TfVxbaGdJe
Y+CZws31V2QeJ7I5CKmA9k0YZ1sKX5DvhD8tmY/gK+fozHcN7itagyn3mDyD5oKdeFByhTo+/RvF
+JbYnpq27AxNnJNK0zjAohWwjX8uoVRF0L1JjJt0sDFgUgF5hphNSgTuKa0TYecMKPXWQ3p0DFub
PHWWdLGy0htug+0yINLVwfZBqawMONZ3hKUZZhoBSVrbexqd1VgW4EW84iKrJWsfiQY+9nCiQb9D
K9n+JjSriyz71TmyzPAa2f2LbXOuI2N8w1XkX3UHVDgI57k52YR3oWlTsAOfuEr1mxHjEz+d05cj
VAx6Amqepe8XuewdQ/R7rcSm/Rq7I5wjLkoLoCB4I9EYLTUTSAbGofCh09VhytpqUzXVXzVLCcxT
DTa6OcJFIsL9S5KII0cep1KcLHpWs/dvwW4wbZxT5D/3bbLt0z4Chn31PwbOZjDosJa6ksQuVmZ9
KDS3afxZTsRriNrKDPj7rj/EvnnhSzGlzF2P7RqITxMFpxEL47pWtoOkQAdzmu3NBwveOAtxhoHA
W3KoJMZClwPA8yvQiUXacgeiOlFVYL+xz6GBi1PFX5stYa/IBDkhCWEKfMLFS16qU8hP79N5F5Lf
LGjwdIMIeHE2ghqoIMcTkM8eSDohBoOgM5h0rWcqmWsb39UfkDxgiadQyLQ+qV3dcPzQIINMru87
ret9JevXd1YwkHvkLWI7ZaV1ztUWvqy43kMVOVEj4TN5MTlBjGvuSZP7zo0rlCYPx+zlTsxvY745
9RYZriKM3hPAkTj7vXwW/+1wkgcRxHza4DLeOR23aZ4pFd8JA/nEZX/lzOpFod/MQcQqzgqHfOYv
sy9gfHRuON4E7CcUbwuMHx/06fhACMOrQfxFwSKIrB8y0Gvr0cd4c7y3f+gOKAAK4NsypGLNIZ7f
O0/W/OnkDCxzJVjvvrnVLTqrsB2qei0nKc4Rgs7gIHc1/ly5WDusEXU58nobN+QCWZrxGQsedvxM
f/qyPCd4mUjS3fykZUTdGGH2/lLfrx4z5Vl5uohUXq1Mgfkaoql0onJgCHiSYYHUgFmjPBO3vPze
VJBlHmeATJN7o8U/8fVfutjZ0r459CWv4TfqVgZJTQYDA8UYaWwF06inRCiW63X6nrX2+w0Utdo/
tZ5KbUeo7Zh/h3O6ZlYP0C2JFx1lemGAUgMuemKjUAx6YVXZvFin7zn0dkECXrIq3ZRhpfqRB/EQ
ZRWzFoP2XUjtYoUHypFeNTOjMLWWKXj5JBHKGZKIepIinfJhGwP47GQq9211HxoUMJRBMHZ1bd8p
rFGpZGnTNzEllets63Qh2p4uwMxvWbmCkU+FXtbIxN5flCLxEASkTbPtVTti7JdG1mXT4x5uc8Vb
+sYJ8SETGPp1Ko4sx749PNpJNipmkTmpDWnYfHzvnBmZR8XHagnGIO3ltMEqV3Jk2kBRJCBn3cjJ
D60xoYnLUJVaIeeyLBB+lThp4KMXKtSaW6Bv1SMKEgEwOlr1NyIYaB/ZurdMlROCSzaH0Draf/Yx
9i5BeytYE8KSpDpHgW2DkG49HU5XBXb3V+EUeJAuSzRBhDpEMC8LBSMwE/t106k22UsWgOjBN2PA
AA3K8c23ZyOP3r+I5AXPD3rbYd6vWpgIxkkrd3KA0H+VA1hszulyfrm7l/hBzHiPM6drfBB3ifVJ
fbW8oF7AwM5R5EzzJSbZcjNe8Jb5BSDxwTEQ4Yfrh6Djvz1xO7F12tuEBVXL1oZrsOgu9YlSszh4
iipBPZB6CrhVgdANhDRWts6JrIAYkXjVerrLi/jZ5dSfsv4akTbGGcL8vTyOx6Drn96kMrUc96UT
dqiPWA0CL1U1aXvy03MmUx0Yqjfag2CQ6VL3bSMV/Sc6p3EZbp4XHCe1ktDSDix63keS6aosxWz4
JZfJNheq3j62igoo8NWBEPNrJwTO5QT6SxZ8m5rWCO3u11SYznk2XBePdVspM73dwa5lyIHf57ZO
DP7h6T21COTluDaT608dKrDPscX+T7fAPyN3UMXpxn/r3jDf71ye5f6xkZKL9KRNNMMDq+Sn8ZIf
yxWsQ3F5BIzUEABlA3gvgJjn1C84aBggtwBhnIUy4YoqL/+dBg02SPeNGkz1pTnY9d0+9NyHXWs5
IAI58XiG9gWtPyt+dkeG8DlihEoFWnioaFz7kS4lGkduS+8KvIT0Z0+X0jMBAaB8dE3x/oTNpvC2
Gz9RHlFFFJ1JLCpT3EPzyKfZJDKJnn2drtN4BrpaTtp93Tsx27IU7qD/FxY4s4eRfoX25oqJQYJc
6H78dyLNn6h4ANLxUTRwSCievcjf3xyaGHmZPq1P4A9G4e3ZAm8/uCoD3un/ZJIFeL0Bp49Bpz4x
e8f2GMRarq05fVv7YGV79g1E2yeJmSppz+hTiskHJKVKBNHcPlUKpC+Y5hdSHInXELvDE3cvyCVY
KVGjqGHPBq9aghHedtmUMC/wCJFC3eVYwuuoENPGrZgIEiidpVRZMEbRwwo7BFo8CxufaHx+yuGh
5ANKAvgf67aFAq1NSpm+MxJ7RuGgW6udrh2rastszBErutpAD3LYLcbWpgNI91dVwTnz6zh0yzyj
B6CU35n7TBXafaA5C7uuYLZk3HAfnSGA2EW8LwCzdXsCYxJbAU6BNN5M+uU1wbJYa96PTAeAhh76
1x758c0zhaFJWDC+gGBGurnIOiA4GzVWzp05a/y+sdzWf7laBddq/R0XLzSixHTkEsRS2dw4qfVV
b4brwfc7OD/MBkmmOZ+WNCrl6RrKAsinyIn/x9ZxpLaT0nc7fLEpeZxzf6QLM6/PACqESia3hFAS
kQ1m69g/GLcBzsoUiZI2JtOTsKNTyfNK0oYuj4PAuW58WjXnd2YK6v+RFNp/19ZqVC3foI7M9WsZ
b43uGW2XAF2+ijB3Kqy9giXECspgLRmi0CyOBUEeFhuqiOI0mQhH/L6x7BUxg9BdTDTi9hPEHY1a
NHqDPMxuOg6WwE81jx0gGcWsUms63NZaHQ/1eXfOX9QtgzVm2ZbPn9ABVVAZtKZm1Zcge7IcelV2
zL/h/kI74zinYFqe4gfu+4dG23UzF8tKtVB9IsrOvTRGrtLCPfSOgpK4INsFZYKFHjXGJFyuup/w
jiuOfYFTr+KgKpwnVoftQ9Vk/Xx3oCPBli8ZqHz4XqR0RsEhVCprd4vTwQHUCGg11W2xLzTH1iqI
g+i5IJ8XTT9SV5knJooI9ozy9PxNPyxoJbW3DS8C3HQWsFalR2sCLieTuLqNCi5yUMdzR/jC+I1a
LY5R17wb85ynvie6A/UehefntSwfzuVVtW4kdsry/2tTA1Zjn4jn2Eu9lm20si/LVcKYMocXVamq
mjPWpMJtkKFWb+PAfeTW1ddWLL9xKrf2VLcywKFzzBrk3f8Iu5+4l6FGp5wb4VRDK/Jz0044i0Qd
khQQN0uGq/zB8EQmK1Nc4IosJysmeFenLxJd1oPcLMN9LGu5qutxrdnangniWchLmwcaAi5wA0iB
BeLiIpq3qKv3xGcdfHe0ouIR9toInLroK0lswNjUgmt1rEJ7MwbL714EfWikEEa3B7K1eDZDy/vl
pJYw+KS6OqyJjUrRoDmNJ+fQGVjLzBpq/DXaYWo+GPsc7JoucsJdaZ5iP78nqwakX1rd+pUHd1Is
cHmlx144l9NsaO1VNF9PT2ZKWPuPUhhWEW4w29NUzV1PCqxhm2KmHChD0IhXiBWB2P1qPl8JmQS1
KSrQMjU2ZPuyEu/dnzlVUvNiG3iGcN3tGyV/HKODulDELZ2456zxMHYz19XVDkcq+ohwBrd6jtNJ
bhE50JKAI+ItYX42ctY6frVIxfWubJtJSxvR5aD2mmhK83snY/fpqk7d6eqXWaEf4CMp+Jp0DoWY
OE2SspprhKezhmS3edR7LyWkR1XUMX/FK6Hod7qmYU2y0MvZEEWcOZPkOmXjcTUzpDL2I9EXikwM
SgMt1VZJC4OcqvmS1A4qUGGJN12j9y8HaT0P4zvUI20PoCe1TbQAWQoZPyVDKiNwN/NmLlaooJ3Q
V+1e1nGlXUGsjdQDA0vEFNTN5AzV22zdD+fhhaFFNn4ANmWW0IEw5YtA4FfVmUNkr7Jv+vFUs/5q
VfWyE7mFkumPXiC/YpFv2PWvFW/X98+zZXr9eEhQjLQJ5jIi3CG6ZCnaHjkKjwllxHmyYUEIkT8Q
IAZ6YK8nqQBz2zmBW1WS7fSUGjZl6XphU8DLR3wcZ7qIcHd3DnI/MrQTXOritvXMeTyrRiVJKi2M
nln8zTEcceccf9P1SxNTZJl5nbVeeqdWxf/WfDEbssfHs5i9TQTg1MoTNVYRNmEOnqGtqXgmlXI6
OXoet/EHjRfcwMrilvDsdV4zM9/2P7UUFt82sJZOOqSnD8hnf7lzjFZsr6twEJEYyNYES9xKO45a
oXvuNIIOgNSd6mNbHh1gUbKLho614E0I23pDnBXl0ZM+HfL6MtY3OE5f9TxfG7Bo0ZqyRnGa+bRq
Bw5T5QHWmkhQF0Pev2/DxghHgpdnfVg48r6ZWHMEEjA8uP5h3DO4I14eNkodGKr1fpqcXo8OZ30q
JL3nQ+Un+ohT3TM13SAh4G/3xkcPT+tBoXFdkANuZCjSLJXYT6yc6WS2BHqS155Ww976TTJtppFM
4snoP2H/1oh5dmfaMqSZSSj0HZ8JpiquRuuwcnGmzMKZi5SFCsgzX+wtpGulc4Ix9kIvs701+1v8
lxX2fCqzRy1deucoXtFbAdvNtfz+5CSEvFsXqbtb1u91J5QEoh2KQndaRuz3g3kGbO5vPsh7sbUP
yTaEvihjYq38NYVItRlfSL1mO227ID8EaAJwZCckbxq/otNwtmo0A7210hfAGxeoWnA7StUextMZ
DJziYU3AtQROrTaG/85wZkzOvaFNaPDo20hrjRZuzE5kETB/wU0ofGoXNxT4OqV3AMI1GyuWCE5R
mgM5PC8/VCzZ92jxZQVm2GI4Mtt0pZvxayhp5EaUqAQjbtDLxsnzR4kDvmoVIuqwg6tuwFFw3FgQ
lqKZnsn61k5EgWkdsYWAA4MsyYKewIbFq1GyXlGD8yIdJT53bQyoTvJlFQDLCV3xl3p2uwaqpcJL
vEUO+5VxiseQTOzik1rfpvOy4mszuXtHLIHgzKJy/5dtEUIwyyIXgLbGjGOJqUKLKtos9gXx2rZr
KziCY203pW58gamTTp1K37UA1UrxfjdE6zJE4YCWPd0JLpNSiOgDgr9arFACJHkQapI0QXYq5nyK
xbIRcYRQfgapFv+XgOoeI6KzZYlJABioN09SoUquVT7B12iRkacWZHZDZF8tjyjNu7iJl36OYR/4
nigYtCAC9DtRRsbvCy4r/AjiUNVYu7nCzCNYR1zvPXPdtU9Uw+5vgZrGYmVQ18dFO8+DNgpiGOPX
yV/YaYV4XVk5wrhNGlM5FmXw+JKkElvlQZ3GUYk00QvpkXT0w1B/tklRwD26K8bb9lgATNW4/PVm
gwB0q1+DwBuzT+Ac+j01krLkXRFicJWZCRPFNfj5rMv3CHP5aUhBKredK/FsWEqYBS0vMF7yFJOi
XroyFhJ8Ym4Pajy3RVqOaVWOGquswxjbhZoHW3ayZHpLvAalKaxp5BM+SQXlCpahZxwWNscJzkWv
bf5yUpe+9Kj9QUUoYunHyjs7x7HkridrsDmlnSK/ZgAZMFqaPHRwp5iTykEAKpzoQuLWu16vorMq
zejug7vlXdHflgTvX3ZsNvMovCCkOAAT7Ncbw2FNeo6hk9oH4Cf6l+uWonwnV+RFnffZthep68zE
OjUMNBEN9ko06ZJgTHhSaNgATDh6Gsy71VWgDX77VIuRdgiegIJ8wwuPZSYpO+5W9kyEqCxv5q3d
p3oz7VqMlTRKfN+aM1iBf19T7uEM/YNMg3cSEgUtFznH6P7fRNE7D1ADsk9BE5aImiaIfatPmZoN
jjTopVK0W+xNjFWXcu2Latw2IjGGAKpBL4C5OiOT/GFY7FLq7N+f723ZvTyKO71zlMn+64EIHNzy
3ff6Q91qYzf9ORHkle9RpYPYNxIB/SoxffcxDFqBN0sGclufQpUXN5MrwG2WTOMKa1Z2zfadwCs1
i+9WS7fd5HUeX7mS6qMaVH7HxLUOqhnUlfBlfzwOiENctLFgG5BPDg1VayD+iDxOL8QtfXfhQNBY
3ZH4z2ufLy+uf8jmH8H2E79Jlvr0LnRz10p5mugZqGuy0fjjZEVfXY+o3nWY3TYu9hFNYGBapkh3
exqPdIhC3dff5xEV9nGJYsDN9tC1aq9XL703zV5LNkTkqcD38tDfdMXCYqFHjJagvLUOFwWVvA50
gte8PzROMEEGVZqckhjU+xXDknPSVeehjZQoihP5l1aWNzbamM22LGpqwq70rKh+5KHcPYNm8K/E
YiUEOMJn7s1rjJiLOrmQwi09t1osfW4NQ5aBDuVgklVzT0W5hyTMY/SnzwWP5RLLEYhaztTQz4br
7hwZMiZCBJhSzCcy71um0tzTdKwYpov0IlEIbFiUA5DIZOTFHUYNblu1dWPtSUOZyKHwl6UzlEiA
l+yZC6jvNBRwqVeTU4kTr/ioEI0ogpfurpMyFcWbvakusP7yhRe8AGVy+8kXLCpgJv5F/cS+n7wm
lgtw3wf2ZWZAsr5qDFnZADPcQ9r2JzDv/MuxjYh9+JPBwSgJIxRvberX5RfxvGG55DY4N9Iffjq9
16brNt0ozAusEhAi4KGqWeI16oB8B76y/4LgDvZoLzW4TxI8NlbdP/MhK7527fm/G5ZVS98fmGkO
ND94Hj17f1wiSk7gN9wSPc1CPBEm4buFcxGTqxBeK/EBCJWQRQT/2E020lg2X0UkdJ5A4shL65IT
d38vett2x+lYqiaLeCFPkdosgpoqSjmR8VDrIpq52UYmhh+AZTWMt94kH4QdktdZdqISnzgXpSf0
YqgJtfvAQSYtbAinS6sMB6O6j/ghaOuPPYp4BtQYGrQzI5JKVwxtqVSx+51TYUXwL0OeumEjFWOE
THTIBmAksrnkLHLPkClG/+PpGlFahjzPq9sm6EwXDyfHsSXtOLzQ5d2ywMEldfcw+hxxtt8K+pKX
e2ehOygLssgRK4kEPdfywMTa9oIRgwxIDBR/LE4Lp8ttpEBCI2yaGpvEVfsi4RRV+r886PKI8cIo
CwtwmzJ/sK3FRdRWGA66VmzGAm2vF5E7940jMDyVG4tKR0+Cr0DkmdBjEIBR9Yan0faDvAKYNryd
B/tE+otVJ1UumrxNjaOXk2dEXoNSWhUA9oVI1a5dG9G2J7UaRpCyvMlM1oykub0x+Sc72sG0Mb3z
vbyC4UrGQlGLD/paDJoKb41HfEdYt9JZ27aC1Swa7r1AKEjPgwqekuPfHu45z4IWhMIEaLv3sSKA
iF+3x3AI/RLeDTn3xWhsiiLARBVrTF5FcBQ+dAs2r8+f33droxtlSenKb05HE0xQkFBDpymogrMa
4mV1DQD3UhsmCG5yd2uFOxyalyFnHLrYt2WpJc3dY8eUbTN034Nn0ymrns5YDlVRkGFps+2vGDd0
KmwAsOXVhf3MVnxWVp47RU1Pr1Vb+rozdSJoviHFenTDLbPDvgjSbRhuwqX7XmOo2fMfHK3TyNWu
e5ao2kI0edQ3U+Q4/VtixHlCYNP57tA7ecHPjpaQhLE2wI3QjZEuOOx1BB7U4+H1bdk3KNt09u2G
PhzNq3JbREbMYVqm81i1DH1+kH8I6UEPplnNn2d8zjnaNcsn02Em75euUwhU+7uQPjrGgDRpAe8U
8ZrPftphUfXUmrXUh5FGOk5BLvwT2ZNSHYDGq0Zf43H5FWFYJFSyMSjjk/CMFVdG2hYe6lErr0E8
0q9ldrK2dTHjT/sXEKW/CB2x06PFcjRJEGTr59crOwK5haj/l+ysSw8dcrY85LWZNLa5oHtjXvG0
/j7qGiX2xtpCX+cQz03dSjnpyrSejQkEnNH5E5dj5xDlZR5hvmia0poWh2CHyVGBL0eOXAtflWL8
6iJ+pOYKOsY8gGL/SizHAm+0Rds4MMVYEajiW/TVkC4c7LrDeVmqcy8Ydnqv6wa2kdoSS/QWTwgg
HH6hIVVDLEVasj8pAazZ3cjxBKoqXgbgIt/ZKGeuxW8VyBkoz/rHQq3r/V/sLoo4ST3GLfMFTfSl
Q6ZTD/F4WOt0D6+ArlF6Eg832xzItd9/KnuqtpP5IXpQDuHjeoublEXhVDSedv452qtjAU8PbDcM
toyyoHjhlAclYVCpyB/ZwGGd15MtyIiZ1i0A5ePfzPgjDwMMV1+QMRBNeTe8YWhxczciJ5cYD7JH
aKIDfUXWPWem3yzfzUquhyXQIq/fMF5q1nL68Jee+Gau+kVu1DWWVXPOR9qPIY6ohZkUfu+Jlu9a
SjFXBMTV98Ul+62mW/6803rlFZ6hrp7Pdbb50XHbtdbEQ2MuaXqQTrY5ikj47Fbva2AWVTt1qMRE
jGtyJpdtQmOtZmLP3RtOnufag3uRa15L2v4c6kKnu9cddtCvE5FsLPpH9x4IKZJF1BDMaitUUbIT
6UiRGZquvF64Eod5QcZL94/VPG+58TP+BRLnPExjNA50U2viC3+f1Lk7h9Pjk+c+8pZ/QfUsUf8Z
Cxjt+YKIYntzW1p9rXDOH5d3GrGBYhmMXPi8MHNKil/yn59kGXMk/O6E2xWh0oQG6kLnQS7l6OWO
JQB5O/slPlVgCiog066rG/tA3QTqLnlNdyV3H7fQ0yv4O0mFGBXjaDxzbwgzaTYDDyHLtiwfMZ7v
j5jFplP8ESqH4l8pbH0hXMBhnAh08GgapkM2+u8AR3Ij5MYZlyt1nqwcWV/h3j1V/tFZ9GhXdKVA
ZCpPO+ZT3/4Z23ZgHY0ZDECUIFFGad5R9kgMddKkj3Q5S1Z/UvjPEDq317tvmjo8kbn4AbaBBcY1
qw3WclLJpmKbx6cI4w0O7DaPk2cYPXNYuc5RSk5L1SC9ZH5BHgRVs3K+gAnoKJtFjdtHkQWoRSgb
cnLzbVcs8wSButGTqPRbv5T+0zsruBrZGj22y8NAhwn2350w0MoRk+lpDf62EvUkucmWDYoONOug
wdCoXCUEoPPGK8KPGTqnHrx6QCt6dKkB0OPLuyQj4YZ7wMIVn11ZP23NFeuK6DNjuvGbA907Zbed
xTmlgJJGSPBr6FqlFD3ipjLgUTyQWY+u6/+yzysfa861bJdRs7Ors98vSypP2bZ0nkLuqjb0VwCj
/XqokviFfxOtWdYz+lUiks6uhYcJytHJrrxabM+VtJ44wLCOUwXJHGqWoA/dxirwCGt36HiePG9u
Yy+d2CxsVnvk0Fg0EJgahbFyTTSRSEST5YCwIZnwqQDoeTAHT6FpYVFrqOUtTsReQ304CsYcF9Rs
PdlezfvxXK82QCTd2bsEW7vP1QYeX/2eUhG3naxC13MRvMfvSW9bS5opPI4OY/UVC+GcFZp7i+AG
GvFjlp5/ZK9+MGcukXpBPZG3swvIPbL+VZvjeAAqLzH4kdus4lS6iHzcJbjp6jJOdrUinT+USYBD
XqNB+WQxuNgY+rBb5z7Xb/d950lJgbVAe3G6clr4nPi/+tr8Z5GHdQP459QS0AESLvGDE5KGWBsf
Z2+cFmDMt6ujIOfJ5zX24Abk2T45VwGgKGKRyqhlFHycQUva/DD216bz+E0DxnbWmyieqL9K1XH7
WxjOH66xpiqSOfTWckYO2Ho1C5eQhDQshrXSEznT0Bi+C7/coBYwcficR1T0RleFvnj5hdCjJWQ+
KNTzCbqFtcIBVzZ1aspP338YysrFvA5g8j/IZzVjr+PUfzHb7reFsRIXIolKyhQONBIzgoH9oUhY
lVV+NgskV/7nCHenV5MUbrcxWVu/XH4g9yIARGKz1ZvYN6TZe2IdgIzwOJghDDEE/Jl5EMvYtfl0
ypzY5gpk5iWdB35fZAZc0GMSYv/mEh13/5tYAkgc6GaT5Mx0mlQREe43GcI9zog/AXAOznb4exx7
glfewu/PzgNKMkYwzzShytbxDUeqruXVBr+E/a/D6dRl5/pVZzZ4wMuhYdRt7ZNWgyKj7Zq/yq7P
yhgCtxsUWB+f85kivqV6bt+GpW7GSxbfnyGp0tnbLfo7jnxWlnH/7wkDd+xJEKkGVUimO3SrQxs+
UeIOj6TvCUElCxpOHnuaD8z3YNm+TtRLH4xJ5Y0ZjpvhhhlIXJbHrYR8M6oLQ8wRLEYGd+NogA+A
D+LbyQUZGqIen7du2ptk8NMg+DlPD4oiEQa6nGl3lg3fw9gZjqVVWkVZ22NhI2WzUIU1J/2iQpUy
zN3Ni2NksnVwBZW42EOn+kZH6RRnr2oCS/o+SwxqNBcvE4cMXMeGqnoLm6biu9bcT15/d7v8/zdq
DZ4LVDJz7d6jLuT3uYBLHmYdAMakoYXb3Mn8OOP2Oyryib7GB6uCKQQTY02GvYsZ1baHUv1Pnp72
jL42ZOq5nuZDQveG6lvNhzLpv+n9jbRIjTZZoGCYoMcGrlJ5OizT3CgNSHdvh7Q8LMJB8JAK65HY
+q/Fu+5Z5PeFz9BXOOvN9W5IZ2ru1K/TZSUt980d8BtmoygMOQcXESO6n+71J01Pr/5OSy1j4epf
xHjPZr3uE+SwpY8dzVlMz4XxuHFqLpy1pZVblTFQJc0JRWxKBt7AWGXmOpkTHIY8jUnsKDrsobYe
OSamDybDJzNpj4NVS1E1ZF77CCR8XAXcEzmeIwdKKRZ4Kpos8GaVKGkT2/wf8h4qH+Dyp2A3jYqq
mANySnq7GyQ6QcNEVI6l09GArKB1fvyg4wE6YCM1f3KzKmobsMghEyoFJ94pEXqOaE2xj3nSiihw
GNrHKhL8+CGaYT9ZezC2px3NptZDTflBHT4qC+YytHJ3ErtcCKNMxMkpO0XOAL+6/GXJ0fMI7+bH
SPAW/nIS5FxzXbmRhtftzCwgb790GOM80qcP30CfgPMspNWTekHRmnGYmFtqTZDoIp86UU6oURW+
h7gBpYJv4e1+7wG5qn0xpNexNPGI1sZGZKqy5Lh8gRc2Q++3722G6olHdkGhWmj3MHepnMMST0LE
Oe9SOIcnFmRK+lX5g2/w102ruTqtuGtuMJvELmOc3n4an+bOCzLPXr5G0DOiFqJgE49FaaZQVKDs
rn0JZVOYOD6a+0+ZZmOciTnquloJ18qjU4GAC+nFjfUKPQXIOnPi9zswyho21TpGcgRg2uwXNOQg
96rfAC8fK4syP8GYr49Rn+ylpVsaPXd4iOdxWZoeP26UbRIbiykpyBop2I7sUmo9sh8j9p1ifuzR
7JlmbaT5xNpQkZf2FFHmMAy1kqkAZCyLPwNNlZcK+y2jFtcsuwUKYdyzcmuHJQS2n2KWuzNlIpf4
XbIneYaZiNQ9Nvo86vjUG+gl5myZ5P5S7ExbiID87SmPm4fl08C43cQmXJYebRRMBY5qCid8bE0h
8h1fo/jdQXmIERKOuXUMNRy2xgJ7hUmtJ463JPbRvUCOUyJf7OWyYj/Q9iQEumHCRsbMxgksuDRh
9Ty39nD2lKvl9CiypKS/cAkJLIs+wncoPuGORpCVRycgIIxeIQ8EV3YvNUtKhuJGeJ8ypl/WbaRC
S3W7nLo4uTSie3CYFiPB9KJhMLl9t2ZN0U3rNBkCVDrkIx7BRH2si52BIwFNAany8JA/E0UtOuPD
ogT1A5A+QP5E0cN7t4cj0YgezMUL8qzbdP6Z6Z83oD9HmqKS7cBfOhjQX/r52lg6zuB36s++/8do
BVz2bjvgXugud4vYYjpSOUi/cLraF4BDfiYOYZ5pz+4MkCOnvDnlsxC7lstPuQvb3vDtdAW/F9ne
5HYl3+YxswxkdIhKDkRJBVnq4YuNk1b72gt9Ympf/JvaaecH7RPC/PsspbZyRisTeb8fYgFKWpft
J+f3jHOvc4WX7cMFxUPFwdx8hOdI46K2dAhTLkqa4HC8O4q6JAzJJmTdBFlKVNDIoRf+1vb+kE3o
VXyVQrVxU7if5X24tXmWqOgJv0FPHvMB5g8zNV+QuQEpab2pkB1smozu/x1YiruDlx7FG/2wWbC8
vr0iBrDIBskWIzeldkNWDjNQ1ZRukQjGoufbPTGFAfe4dkfS0ks8xY4Ycj4t1hoovIqxX34Pk8lz
lU+ZhUIeeCJYwSG71ZvWaV8Kr0TkTi8NxSoU6UCLywdwseXZtK/xH5FNNmwQiWSF8Tsfnof3wS8i
2Bo83zhaqJVlDaTIRBAIALk9Uf7va0nCEdWXJnNEWrjQ5KCoK30u4JnAvKcwBU8DRgW90qSyhCbV
R+/3lrArqTAu5AWqsO7jOQwfRQprGT7KBEVA/G+UBmH8uBKS72jQNfvj+DDRp3dAuBKRPwk95LtG
NR1hPc5ySMrulcGUuvhEtJJTQ37gyXMKvxnaswYLYDTFsuASGFUUBjniqRki2DLSqgJvTdfWbtcy
CEo8HNZ7PGDKoxUoly5j5V19n7V4KytwGpekADzmMtVlb5SvyljYcwMFflImP0u5WCUVeubyDEl+
9fbKg61n/bQIpnbfmHPcjhCs9pUTBMh98dbR/sIJ4oITJyuvTcy7ffvfsP8fdP+snm2CgaJ0qFd4
tKb9M4VDux9pjXIIBaOMHs1fFrMffjo+NBNubrApf4mo/UiGo9Q+//N5dkct2Ky/JSbOnbCRZzNB
mhQGrc12OrdKz4Nh/cgCUskpZ1kyRT8pAKwgxC4TemoRReuhUhb6n54qtzslG4NDC/PDEvctHKNp
zfkmkRkimO8c9VmmukhvuJKwZ9s3Ht2Nk0DFVjZTdM0WfpkKL9AmUxniyMkP5KS6MDjOgjZEZoUv
42PnmBKtfzEezNLaAFOG9jlEIkZx5NK+5zHc4P3/sDlm1mKcvSJ3FvkHK5YiT/BItR1Rq5NlE4KF
ryuxvcqcc2SQyvkM24jpnE57N94Xg/NUAdDY+G3NMJB+kwijFbq0wbGX+cMkUIMbo/7mObmaT0sp
vaFcDZ2v930eM/ZU9CXhpwt7riQdmd1ENpw8bM5quYHSsew1edGeMXr2mC4ychL6z+cMEj+x77y1
bVCUerY2a0Hkug/pWVYGKMGL9O9XrD/zSkMcpbrbT7b4IOGaweOlDh4RTXcqHCNj0d+g5fVAGTY6
qyDOYsnQJJ+8tAfqlTzcH3bQBB+sKiy06lr8/5wnagANzFFUSLgLOjhb+GM7An8+rEA8EC3sXhzg
ElIAGqNejfEqU5AyfS90JcIg/jPszJzaUJuNej8FXgjFseBaKCoW12yCKH3hcPChFw+p7umWfKjq
uATo+ufMP4HZ/NUjZWzbYNNYm2HvAF7NZsfH7gVjR4OGYX2KxAQkgDW+3TNmDkYCBl9Hjj9/HMTV
rnfwjLLvk8ycMtsEVz8QrrzDfKPZWOM9o5DYswIAYEUG2bJS3Xg+QswEJOQgqpDKoP/fKblczeW9
vM3jBGohGQ2bSncWlATbkh7hWSNUoK2pS8cLi0oRsU7Tc9ElIhCFIGZi1ROeXR5a22N76zKR6UCB
ZPyE/DAhkSHfJ/Z4HjV7ZZHeZKzrLtv7UQWQ16DLJoux9k3fhWJFhUoer2ajl8oP4/YbFWWABPRE
LBm+XOqZZCyAEyChVM2bRdLRF1UIEqAnQ52GeG8k/QFEDZDnaLzLSA4awLWQnoZvAtNM2ItB2ZNL
+vr4CBtqzfLSCmJIOWICHwpRU2LZ1afaN0YD/6XKmX+l3BVAUxO+nfGqs4XUBTpNr4mrPQ50wWfT
SS+YKEo9QZDDUHUm+oQNfjBe8byBo2/z4oDinB5HJIZQz5r9lUtDJOBznLBdF+rjsj8for3XVUVv
pbqJIi1y19OLDW2LAGEuc9XJioiI2roIr7ViP3wCKS86IPTfQfOTKn5pAKl14njUckp+pI0AbfUM
1XeFbW1n2NNRWcdBvswM8UqtbLgmlNvSR+471MkeBWNwid7zzaJZYJn/2MY7bJ54eNNjrEjrxyGK
uaxo9D33823iaIo78ZryMqV4KzsLtdpmnqN+ZCgoVDfA+U75nQ4I0Y2q97Q3VpWTqR/bCtRwPDv6
8cPfJiDqlIfHPTQP7lAw6mx0V6YhpYlVMaFe+XbZ8gOm75tqueCNGRGdExYz78nRfdnKY/jz1P8J
OkG3eYjVbPgGA13RL4mt2LsVpuIpFFV56VtnzjDkzLwhQcA6kwNsqXHIBdlQNQ+zeJ/E7f7Sg//P
CjpAICILBaTCq59rSgCYbUeyW1QXxTk4Y/xB7hdFZRI/+XeBHWhjCWh7jUP18ZIXurTx8NCuKhm4
dAZldRUyyqKxiwBDkP6m7gKUhBAKAM26gerxcJCIjinPTNBUtCfORdZkvyRNuXYr85qFQISsbgtl
CKz4BRNPNhGf97p+uTpuGq48BeGpmzBlVe7n0HqmPUCx/2m9reTORlxbWk+M+yEjcNoDJUSN68Sv
tQ4yeXrotbgIPlo2pEa5pzke1TuRGSkvSjH/2UzO+rP8gnOLR33y/DCAt4C0dlt5k+BBcoO0UjeO
piyDXqpp/p6kPf57WMyFoHoq5M9fBX7osOegJnr862Mxs1HLLln9LbLksmJ803Gk7kk7VlviusZw
/WAcjMcTGxOg/fsy0aOPUwlx9kRSEi87wlpSMb8ISug4+ekPW0cf5OjlTrZi7qrrFkOhbnk6HPp/
/MWK+nkXbvZEgrsSK8rDwvE3UlxNa3li+0QshutqGTDrBNXaCgNauu6PZz8Em0UkWrzAgGtuIUGn
LABiQwuSR2yIVzMiORN5n33t3iyGbkv31PVv/S0cJDfeQa2wW40XjcCk17Wy+8g8O/VkjRRvkK93
538biHWyC7SQww6l7k0Wmx1xccQV4BV0ME5c8nrbJUap3SSssOf/ITq/7laXwAiHW/VJUQ6J58mN
kRjxw12lx1t58KZakHaNrc+OKOCBrAxKg4AMyk6qK2mldWivhb929Bgv+yL0yMVOr3eq3aFMwwGs
cfycyWV8lYYRwhRed6QpG4Y5mh7Q14XVR/s1JaSQZJLfpXzIMQ6h6H0Ge9ojH07mCsV9iy8N8bkj
QGK3WVta32N1VMEKJGjpIsQ2YHId6XKSTWQ7geZ/aBVcAt0zghWQ3NISV6fKW+t4LeBK9TZbj/Bu
b3Hiz7cttpjCJDkQV3HaiGVE8F9d6SCB0zgmcaXVPATiBjc8QnJrVhPQQIqjDMOnKVjgjP67tyS6
x5d0ncelhcwxqkC2vqkGsE9cxsU5rvxs4fhmLfw1q5XvkyrIR7NoD7k3YT3sC2/C+qZNTf8+irZQ
D2sQ1jV+cJZb5Z6HtpAlW6XIekP4Q5bp9V8HGsBioHwmAfgi8nbNswNCcANC9GJCSlB8k/ReuDlD
4U5Fa73w5Hx/tYa96vw0DMPsILw889k1U4cygqPMUOMI41f80qdJbB75N2mY0+TH3HOHcxF5Ol/U
OtezDWZjB3rKDHA+Q3McoiLyB2EF6zEC6bRd8zsMiwXaJwqOiO4EWBoZ1wxt7cZiwwKTGA3j8gjb
LKDGnUyWLKJ3yDNVN9o92ZN35giA/Q7qrwy3qbN60Wa3wWgWmfRJ6gq5dPZXbBnLHtWU1bHWh8Bc
BcgHip5szvkiQsMUgqyq5H9PtU7rGjHJuIl3c+/h7kRaMYdyBgF9y25kJibfFTE+jDfhOtAX2Pix
7amVGgVAT59sScNvSxdKcwhzocpNACQIl2esfoKr3ISKX5i0MWH9u9d2ZoJGaoY8PT1qX/XlYBsb
b1rJWsI5zHNZagRccGLVVeL2IafgVyvAJ2F7d9tcIun2uSGFHvr7fxklzg20Qk6QUQzs70Sv/f9y
VTISln/8UEAkY49m/3fiNLWlu3WbdsCzfc+6U0oP8psFn+u6+9Xb+MkZHYaaxsA6aCiZbCD7GtEq
OJstzxsvjgtfwS7QeD4m5dNTuSEzPUHGV0I4uGoeW1tTnr7wpxP9GxDT9j681cXLbbO0TASoKWW8
bNmbi/GdXJQtG+0hmsNjz3FcuNAEgXEudbrsY5wPlG9UHV2VmA8u1S7wHU/vrKuKNufVZYDDwgaH
yXlUJf3XRyx/MT5e9bk9UqZvFMmOWuZCqoJ6DIyrWDPsbBrgPqKKYPcXvBUdXW8KRXlcaXj9rSd5
rDt+ddN3cyEnjU5bRDWmwnFdho1BCapHn7AfWPQI9tTxC5rhp21kEnol0GvKdv5+PuGRTghd8klF
fTz36B9ZMNX94JzLduKe2DwbLjki3Lw297zl2/pvwNPToMAZ2504lJ3vYDmnirWhUFjCtjxWO62Q
xxN1lpuOPuM5rI8gvbze5Ba8v8YUOJzS0jKTMYoyqsqz+eDT+H5UZoKj2BAfULohVj1sBdjdxrA4
aaKkOaCIiILmUk9K1kH/799mmfo/ycjWAjs9UWVOQmDWM3M2VTwYEKmd4JlbzlOmaMs7YmRNo3aZ
24IEgF0hd+tr2jbd4b2XN6+c3Q4kg81RsECu1jZMbc5oDz6+mr46o/3hcuF+NDvTBF18xw9BGn98
TJxqW6Flhzy9ouQiL3Xxq17BoFARhUoaS3x+hnMxXF0EKUXNk6jmvVEOv+6rpE2yO7eAKRRCHoAU
BHWOmESV5NsFEMiQ62h6FtfdIfVwKKP9MdpGY15pg3FtcEls/vzjsoHz1rtx2GZ65ja6E3svttP7
P3qixXrg4amxJI03dzxRW8WXqt2Zotyii2Sgqosij2WLHe5dmckFE6SqHqF1vNa+XXId+Edj/LBN
GR2gF7CLKW1KhMx9ve0jGbHRf/qRUiD0bVweCaQXUQp3HBn7T2/G3CIWfHK0HZoUAkdQax09ggyU
YF7X+fo0YtwTX8H8M2HqWKYt/GdRT7EFhRFU1w5YKX3PDXItfJOOmFMLcpUE1qn4hODbtHyYDZfr
FLX5emLulZ2AcbPNSKZMY7J2+QcP+ws0Q9QliPjOe7amnTeFpuvEE6Hy+Lx76QqQrYleaOX7XE7i
RqvHpO84RXLNGX8p8x/Pz/yGM892GkyLIPM19GuFb939zeS3pZPxX8bOiSzEa5xEYl3NElBEoPQg
etDN5whHjqMI9cCj1k6YJKK0uK01TvboAkRDEboT7nDNyzj6pshwIK90PvczQxeh/+J/P4cklTF1
sg4Yml+y5zVKdQcjwUi3YmyQHKmL8DFP3rskl3Bc3zbJ6AcIsTnW9XK7YtFrC6+MT75rF3RYqg3g
V1rg1jy2AumOm7kGjbnpRzYq0t9GNb1udifhMdNh6h9XbRtCE+k9VenhwnVJd4n9HGwJ+iDhQIvl
ld+jcGXtExONt4YNThK6AIbHcE3bnc/2dnPmSQGLNSMe+jVXgQnopXiEIS8wgQXpNGgubqn9U+ju
709Qzi4Xt4Eb7GeYUvrX0DajctVU9/6jFDdyLwGqck++wnzesoEvhVUAWMJo3hBNyqM+nNx6tgOO
kppmcjjQE4HyNbzF7DCOlgEpyfZPXKXVWWwgvB5Ie0DPy+P9hRNm5IToZzVnF90MzeGUiKNAIxxk
f6VgdQ5be40ZrvCERGMfPoePY5IQWm8iF0qWHyVn4JcJhRH7Ek+hi7fzofVGJS6UHQk1C5OBUEIH
yFF+TYIzkcJZ7TZpE0/lNLYkEcTKgpw8cCNnyhMSdJoR3q+2K3bBMpQX1oIr9iUPDo4G2vgBExvx
duBMQ6f2MXLZMvAPgFhJzoALsjwdqi2eubTCJ59VDkmi3t7bMKz0i6o6oNpCQaSxP9526FFZKbkT
B/jJu7lwK5d+o+lIY/GDLr5I0rHGjKXzdLttf8MphOUz5hC39q7/qo64U9oD2Zd7OSXJk1LB1T8W
cTVSoV+YdOoljXO0ixe0t3QYZNN8k7joZgfCSbuEORMOopkaIaWv+kbXC46TFnN7/LslfF+WJmUH
Hd5ENeJ4Z/vF+2H3Pr/78uQ1dOKN6xPDj8lEMb81jzFIKfK5iK8/l997omHXI02MAQv7fvrQPxPB
vPeyIGojOxviN7KiXcBKeOYDh8Q1WLzBDnnV7k+kg1diMjoowXVAOyceZy6gxzFq9Z37fQlEeOF9
ULa9gjI0HQvonH2GUwgtKMgKFeRs5Y6cNO5BJEw00dx0k9dYc87O5QiPb+NZw/sBR2MwAHwQORbS
lrI3hiX9QdG+X4Kj3daTD7NqPIQXsQGOjbxQVp00MPTh3TetDBbeHv6602gX1cMcaZeuNjotnVnR
CuwA2jR96ZX2mJ9YgZ9FXVqup9cT9jYtiva840PyqMxfvRYdrLqyp0AXbOyd7Vrm1PyZCsyVv/Z2
cEFbrqDh2mah5KnLGpobNgnQ2C3GxDDLsYbUcJLZx4Y8L4Qr3FUtZGER5xfSy7vgKrAplqXEGAQt
5DQZbA981dMzWr9z6aMd9NcPr+WulTL3MAmVHNAPQo4E6w8n5hkXzrEZ+t7zZkjFpyI+k+8uI8ag
zTEsLHWg+gFu1fBmrhRK5tYURFEDiRn7h+wQDdhwcmuUJ48K8YoNxoUNuPymMyYml0XooWzzgHbn
3+3ldsg5G611XaQtxHk8pafOE0R+xl99O5xPG+c0Yu1Y2VbEh+hSeTXcRn8XCaZVQZqG9rbITWGF
98kzCkD1VeMXgmrxLb98Q9qSL1/ZX+Fy2SjxoaiZmBMIcZRhJhmQlFXQa1g3UZbvewuZRdrl+i9i
F8uGdCFvHDX+MXujP9F/5FyP3XJmx5YFeGzf0YrJcnlfbYBo/ovT5Og4zVdr2g0NxKrz9Ztt+o0X
4ZlwVupbnAW7Sx8B2BW7S8TqAmgnmGPwWZBdSelSBb2RVoSiy+YxKT9EgEPQ9Yf7TMOAD5GeYoPF
fpViqxr/gcS3TiLi/TWc7HQ4CvwA7q2zTSva+xnMX5q2pPhUvveu1t0RZAmHDdxmWPmpfUuxp00W
2Zf7AvVMgf0tCnfGeoNFEVubxIReCM7dEuy7J/Sxeso/F3zIxUPZDFuiFHImmeUb8QdDtIf5+nlk
S4Xvr5/NIHtKq1qcqr47gN6384wRgeYp97Mc5VjR3fVVaPQ/btcqZpUJFsiKe0knFWJIIbTPkbCZ
l9xSeqJ1htxrjK+o6wg9o82f9juzbiqXXCfiyg8UL0jbF89O6vVexs2iM3SwlYHvUPvHQD+QFPW/
Cfk1Ki8mB+i35YOgyCrgQpUuxkzCa5hlza/S6K/Fshqxmw5/gX0cGsb9WQG8ephWv81rUkQuVbsx
mPmeN2lKhyHBCt4utgLI0elAiozJEzIJF8yNxkpc4dZmbxVi9nhANSLe/+xxWZdo9WN7Q+jL/d2m
B4bcTqjab6qI5IQQvjnpuses8ZutqmSplajetHiAqaWau+8FE0FZk/ZLyoJMkDIozOGjF2cLa43n
cGnldYYu6nvVZPrIq9uJm59AdBwmBBSq9D9loWI8hIvAb5rdhMU41fboIX1c+IYjLTozL7pZSUIQ
jWN/YPOFKvXTbibDD9CzvJUaW9BZiMAANGdpQiXUK4HGEUJjJzST/TBfQ1P7QIhvU90jkz+mr620
l6gvoqYcRVn0aqtLUnwjxudDgv0ULzdMFBA6G8u1RzYhOgZmkJS8skEjl8TyGz21ZVwkUf1mDh/w
imMlUVPX9E+Qv69kGHMG00Y+aOD6BYts8yyhGGY0/skQnK/DQRGBUQpdMYbIQ9kUUh90qNQg1Rbd
t8qWjFqKmwv639GGEk4pJe2clvQfG4TU4dTKoL335tgE7MbX1c8gFAIc9YCdGfZywmpDMEPoNzmJ
fMg9RsaTu1y0Xr39PRNOpuxWqHV0cz/zruJ/93P3/ROsXcnBnPS9lpl4hfcLXjXbdM6kDZ23ruKs
0lpiKfZ/a1Vk2wIOkjCracKQvtSkjXb8T2uFlj482awmBuazzvnrCpnMViaS5C8LPX4fQpiKzfiI
qOh9kBhlFTztixgVWbVhnCjLukL5twN/J+sTRABXwPfOSIMsJSxDD+wLSJJ3WCuiltf0UOUq5Yoy
fLnNNTalfHaatN59HeuqdUxmFvvfGFXHAwowU9ogY7tZKclHSV5/0WiAxgvwTvcGlRxlJBX4pZD/
Q120wbZINQgaj2lma4ZQ3ylvZbhHf/dx4YmbgaEy0rPlWI+vfOq29oayZQ+QX2UeCra5jicgemoR
1Wd+e/BidkmjMc2kP2r0Kup+p3pfYQCA5OtyOXL6cgSvHwsK2oOoBUbufkkqWSwCd1yGTJIqqW4J
29JrYGzEY5a9UMhNQNUfxF7Mm/NjFAFVXtH5QA4v+NsC2VBw+d+Uzx/SgTxNIu+C3TLjFjPdF1Yz
Stg9RncXBtzIGCkzDrr+ZR8Cm1uvuHf8C8yftJdA7CuT8amSa0NQ4KglGvwTtnAhDHE31wiSJmLO
cnDknw4LqHY2haUDdsl89nBdqI4MkFXq/tFnO4Wzi2pXns3pTF5DecgiAWipU8fDUQzoZIIpTm2v
YitwG4KZBfmQbAfILHgutCTpOC6KocmQMAT1mIFgwPclcBTy4uIsiXIY9022bWRUBpvvOY0vLw0L
M7TUn3ADIae30qvEJ0JCtt/CPw7TG9BV5dtih11c1zr6ZEmm/DAp1UIGj5fhzPOoJH1/HsQBIt77
Ef4hAZlxNBmqJrgh3lHMkyp7Mb9cpq2oJUmiH6PdWAd7lj9pu7CexjVqnroJbK9TyflJUa+Qc9Ww
Zc2RKBLIyNL5w96WOldwVdMV1dyoHwgchsq3VQkOkFeViN91Rzf/iYc5IezgOR+SneIOHAP40n5m
O7iGKhv+pApmMQbPl7g8b9uc5+vS+baeDywDd05Yl0owRcrrNB59bUUj5aa94rRjMmWyZo3fYVYI
0s8f4KGez6vIuGnzXh2hEh2/WGX57lPcvN5cBB3x7jbo4vryLAHP6E2Z7+YKyxcLUsChM874kRbo
V1q47IY2oG3LZzIR354RVReqzkuDZmd+xdmCmYwSZtf9wTjO/BHy2utezQdogdwrQsGSrhQUWXQ6
BSYGT1SZxyOIGI8Er717uGXtfK2/EoeAKO22ZoY9xA3rNGCWsjksIlKql0N8PMIbQl6vLVjB4vuB
z0ztDHwByJLvv/Nbzpe8BjxTplQKFqA8yUTAufn5Cgfp3D3AAhUHsdRvbR4UpbjlTsp7B3CULVAV
uNX8xuqY08O6AGI29PMqKz/fgbBgQI5LSyQ/5n0Sltt6Tk2I6GqwJXxmDFWcuovGAXqczCUP1dxK
lm8MqLhAqviSxBJ70bXv4D2Eba4EiPXrUJj6ob0mapyaFHV8tTLjEcy+92MSsdRjs1Ho8ht6j3dR
b2KGh7ha+v8kxitK/J3gpQpZbUR1d06TZmvJa0oh+Efj8uMLMHY9Bk17xefSksFSbWmLBz8thmOi
BW+AK/51pLfuIPMlG5Stlw3KmhKKNNfqFGChn8jqlJp772lR5z2NCqF9J0i6PDw8lBepO9mXlfaD
qvDcGx5m8AOh5KfAwVl/rdAnXQrWWkj0xnHsgj6dpSQuyWKgIULx7RQOUwsYImjwyCT/IDbxXYJP
sIwtUshxBCJ5uLoZHJIKyNsugAMlDkGAH1gTz2Ifofb81sPqh5AdGXI8k5m6ffNIv2UeajCDFRsQ
2Pb7/CP5HQToFL7JZtfQ4o4Fq4kruwFocwf0Pzp5oU9VIPLnlApSq/JNdy/lNKfwE2qOnseio1A6
jXAc6FBLB+Vj+EHazMizi4mexcw9TmCWhaJ3KHdqtCEigF7WUstJUEs3slpg/8um9UzoSljU3Alh
+L4hI/YCl3yqe6qwz3+ewtXBTT26aBopzZ9Mp5MD1bm6KbM5jYlwY8+svSnlJD5FxjRNoAXNpyIw
a4TGo3qipl8LYYgJ7qQM23vwL2s3u6k527o30tcsx0TaUuiAFrE7h5HosKlWLRtQx/M0AWdp5vjN
VWxDoXGOo+ig+rl80yT8/2KGHiV6rS2+ltkOHOpcvxBj6hoidv7pOruHQhPBSLVuIuiMH/ynPGqI
IJs90/kEvCyHOJ+zjbJaRS4d/imkcel6YgbBEqD7F4AsoZDzmWcRn464pXLLVv51uBX/f6B+rFll
1qhnDyYEjH9QRwszKhk3pPcQza5PTqgxOCIfx9dbOa1NOGscxHZGUKkuOH4sEGXGuCoDOe6S0ns1
AGvvPl+vW8fe/YHR42bwXRV3C79sMyadeRZD1T3g5T/f4Zpba1J8XrIYReQ9/M1lkJC3pcEXqcK4
Jji0zukFNlrMyU4+S7eNqTJUkGFcBe/59YZpixOi1rzEbzAss/a3jxf+v4IDuHBMHacEQKaBxH+M
0zlW5Rd2YLxa8nh93FWEgeIFp4bZyDc19e/LvAsbiNKLcf/1QE5Qd0sHAt81pjLNZwIKHXiiY4ts
80p6amjv8JwP9pii57r2UPEqKeRvT5D0r5XJISaessCwWEB4RJvgfjTVhpv00HuoF9DiGvUDprkW
2MGMNCpiLKb073TivRLpZDlXn4DZ7C8qydJdGIIdDhbxDD3RgVuQ29IU/DOEVkyqcQjA/gB7xJC9
kgTYckkBnIVIywCKjwswowKN3M97jswQbwdpXbTHo+luOxOx6c/uA20CZ3q0qVfjqTtjPlVZWOBP
W9Ma75KmplR0hGhXrQ3lmtyGJhs9LpGgYSmzNLmifN2upE821o1bUFstGpRyL7CaZrdKbE7aapUg
wB+he4IHDITWVRJuGLvEo6Qh8cFkAASdvRR4QkB0bruVhGpQJU1cVT6H8yUyhW6joMqT7pNRygUu
jj9yHHABWou141WptVTiwvyZnVTD1X0LFXi7VXPtkZ6zSFX3IypsfQWmmCh+RT+NBtcHQiE7GwXt
OvmTxhfZYrBXK1oVJLyS57D009NwSYRLqodLURuECZ1eDW8wdC07p9FR6c4WIaaVaTz/YKXMuH3g
iTaYGx03oFzYssAfFgV/u/LeboHIydKOi5+2KlYrgis2xJobewrdK+ovn60CBs7VUQfeBVV3dqF7
hnnEvolQHADP5bvzCMORZkRtKBEMR1+cOKRRtof9EJfyAhezA1+C0sHzrcPTFDOzZN8EUyNaeSpZ
wPbJ61CgjxueM92IGzmtvHdkALtOxC+Rd4b9TV6LAbQvK/k6O8NhXTrpnLHtXmYJ9iLBALxMeJbK
P+1DH8V5rIGz2copbfsqxsm3ETgDTDEf41MpkKVsTmNfdPNVhr09nNvHWORroH/E/jk8DKPcJfk3
Lgg9hkDBnU9FXhAxHilO+6H+AHitGjiI1rsmHXHCi2So2XSDEkKszBCkDL+CRLaVUrlDKoWEq+Ci
NE7wBjP+wwHbZsJbcBXVtldCdkF5dAts6KEHvTgKiElZrPkXQi+yOG4Zv60KgVVypBE8nSUIp4yb
6BFAxFIo98eABn6MPsqOJePJFVjcck+Lvt0uLLARrVFEdriFhyEG5ewtDDpSUnDyEXI88ZckSil7
yukWWJB7obihr0u0ttJ/gz1F1Rfwhr8jSITIUvcogcr7sCIOdstzK25dmvBztyWFbCO9RCWnDnOB
QBx5UHskm0KjPeP9dKZcIxhS6+NF79ZrnNCrxBrC4Fuy2rlbXJ8jbXywMXyhr3pEPt62c+Rh0PNC
4zqk6u1P9MTItYCrxlcNzHXbc67w818Rs4vJu3nDTMUGs57coieI0kShOo/RiOSLFaa6CnATKQUw
R9IqA6COlzrRDG0WyhQ6FrYJKNn6ckljnm1ncK0jQ+5Ug715bDXmvlwvLzyqJtFtTJM5thuoFCvz
ltYrdo9d4JzA8n1TJcFENqCMjx5xfeKlcVp7iWbT7pl7qNNIETNfIwe6yzvSBsa329j3pB8oUzPi
EOZmIBpkQVP+6BHtB+B4KcZ7x/9a0ZGqwq3ivYT1gYBTnReRcb+tBc0Muyq42YLlRuvMpz2+fy75
q5x4HBcnx58co7JN3tXqcfuULH2ryb5Ky/GWU85NoD2dkGe2eOE/OQEBrXYyv4WflVODnYp7rwe4
Mt4bvP+3RgXtSWooGuQNBG9u97WohvJXk/6lqfxVgf3vUFNjaigbWGFvsh1xlbZMoGjW7oAEw/QK
soZ+BuNvf+85VVPwpCtNqMg+lXCksuca4wIofilIo29ECJFrt5pH9oDrAHp4W5wssVEj8zCXDcEB
svyeYCiESiQAGiww9tJb4saMALcjIwGPIZiqZpCgrQRnFw9RAIQ2iQoOyIEke1NKNLPmS7yeXryL
V11tZp5r446GLdXy3NXc06YhfvKAMCHtxL8LEKWnUOflPvJTPm7m5FY3pjcDFSbQAcDjgPfqEb+T
KMlL6WE/t5qZoGED7FGhLSeGuGwUgwkCIz+5gQz33N7U1qdrHSZUwseiiP58BVe602CaDBvkP21D
IhjLEmAdQLWeW9dGL26d7aiMWx5p9hwGdDjKhO969pBIxxQf5XxnWNzuWAtQPiLQaupWgcneERwG
Zb5o19/jwUI/FsUfVgGeg3hgnNBqlyuHRI0zNx5/549Lc6vsA3bUtk1yYBOE5KVCtwIm9h9S4r9A
CE/egE1EvDbdwOWrMOM7+kCxDPuFyoIquEyPCyi0uELf3s1DWucLjAXlJjl0g9tkNS6AAsRMkJfQ
qL47ZS+U351n3hBXyQ8RQ4/Bs9IepXpXzw7DHRCWIMIW552bN9MuaS6PtxlRJwDFMvQamZsC0YGx
M+xKIDkNN3gMdnklPwj4sBfuVJQolflKiTUvKID8lZxU1SlWj9GlTbWoS1uyaifTYY8eRJS1deRj
iFY0wjptZfaGezCT18oP2ZF7X1KUWTOv1jcdZPmrRmZJHQhTDMkCF3JAyZJ853Dxp87Q9CoXDabl
+fGtvJThUcrlS93F1oAXIi8H+c51M9aT+pmhCBYujcFzGt6NPP2WIw3jFVEOoGPdMSy5odTW4WuR
GtwIYuMDDFAcAqRkZpbwxAYgNrbPgh53Rl8xfXbE7tofERrEOkdtCuNQr3HFlqDoYHxXMpsACpsI
fLBU69093bhe3yPdPBkcUOpSrMlUH0Sw1YBLbS2zrhPC1WNBq4AMee08aINAE6qddY/sD4p4pmcv
KZnUKmM6mj8OjODn6TGPiQxVWPPWMWN2RM0LML3c5Ak9K3Jj3jU08fThqUtEg9hHOEAo5vxJyW4c
KJls3/kxM06Q6TOoteUya2X53BA6JAxaZNypeKdRduqVVudV08F6I0sixonfpcAxEAMdOD31dJ41
suhOkIST8HreQs01Tqb0uCWlmFRCMlfjOJuXQd11prvUO5Rko62P+oJeiIgJIZahB+m04JlIFfne
krn8r66pmz399FyBldx7mYPkXK4fPoNfZYnSEJEkH1CkSFP0CKJILrphPy0u89NRWz06qG/ithKT
MrNG52rxDfa3cKuzr/9/plCeARnR9VDkpD1VdL4rPJUU6fZVwRSqowWX5hnYZVq/EAFfj08lDENE
xuetvlvty3SBVwaJTU27Wm1tVT+SLJA/rCKsD5gJVbRFfeLFC/AnO1i97zYyHYAoxHuIPj13LRNI
DcgMbhHF6IJW+rzlXZr6nqEyWiplfiBaq/CxOw2ECgjtkDN61Inx/uIVBVWj1xa4r4x8YQnNIP3/
br4Up9XdPKQU60F+7f/oX673WlIKxr2F6SF7qlYMOimgFtq22NW3LCQKQNI3lJ9s3ydHVIxlcNzj
2UPfb41/s0cgYf4otJi/b1ZGw/+mZzGVAWQW6moJdSFl748RTNGy7UKW9bYsWg6Lkh/dLA8ZxMQl
KQTx5PYkG94BWU5nJXmDobONDxpOs3gNl+xlIbKLB1NJArtTQIjLTjpZ7VUGMWQrv2fVvCM7p1xe
0RcH/EQ8grvCjvVfHUYiAga8Alqcy8RV8FMtzZ0iGiOB8FlyrW1cHD8CqVIVicFPMLymE2x0dKTf
N4ifJ14v1sbJl9TXEw5EScGdXM9CtyriAAbU/I3XT5xrhyhsMKKGFkhZy3brRWMPxwe2buZINQE1
jZ5EmHrqUpQp53ZdHokTAt0D7Qxwc9aTKVH41S0eK/f5CyI/pq6+Tx6U5tDZ60Kg98YeGAIrdFt2
lW8p3P5nqpO7yB4T65YfXBGHVg0tpG6bUeV3XGRgcb75EzZgz6fx0WL3E5f/dJqx/tPC7so3zHzF
DW/UONj5tqosvbRosAtrHvMYQL1Qd2IF4D6aWsYvI3JcTMVJXp0Zyb+Kk3ByfluXnMaSaqI012J3
zNS3bjGhPtZKZ5wTix2UaoQCw6aGrRwrc+h/lPhoTlcGufkn98pqYI3uxtdQB8/BAJ9yrNM6bRLs
DqiBzC7/d+hIo+jZNsaiVBoyXJ5OYjzF43EuWDj7k2wKIjZd+AV5DLb/FQA5twt8WpD5WqK9lJkG
bUwfsT+FqYyK0by9CsfQiaB8qzpLPdO/fV0Ol6o/0udyFg5ce0t66wY0V8MML/m2kfFmH1dm3HGu
8DvM/tl+fdkeinhye1AHg7g3eA7ZUUXhsS7xeJ4ahz1gglO9W7cfFdV71W4z2vg+OVu8+Mu1JHb7
uQXC/LEJo5utGY8Oz4KrjYGYcTMdus5ZOzl78tSDhYzM6W+nFDsXKoRZ947xTA0zmD+zZ0BkdWI/
Hl3liGWBs5L1dgp0LXdysmWSCDqonGi9lCxr7l39c3ihkLzkthehO78d3FetdlkqVWMypgV2cXtf
Waq9Bp4pTGXaDvkjRk5MDlFvyRDKAZFVXNM+sqYsys0eLfEwhN7bTUWWQ5NdJsl3F1bzaqvLh43+
BB6/A2JsQ5QD5UHazcYAarymHmlybhpxuPIqKl/QJiFoRACidKCkUIhRTkbMl+qzkFN3BHVaHRGU
wDzRmd1mp7252+xnYdthgosU/lVBNoJQZhpfSzqp5P/FO6fk4f0b4T+MeJF66s0pD2keZvofHGmF
FV5nXA5EE1amPUJVAUFdrmr51KNAoVyNhuq3hGfYmfOCfdJspJi8Rck8IpE7xk8a1Q8PGw7efLC9
DxarDncIjbDEmL/Pe/FTMhOqGoM/OwjVDh9LHOT6smQKfKzcMwzL/43JuGqXd82n+M2rqzQF8C+1
nrlUvlBMGfAz92og3cp9V33+vbM+wKl4K3FaYYqAXs4AfUMEWPBC9xHmWRI15yo0QvudEDGIl4Bq
F/PnaXECQN2vRCfP7sj0U7b68683qzTLfD+YHbA3xbw9G73ZTtn3e1prCcwb3nmvwveNwA1wQOVv
O3g+zE/ZBXI3w6sRrAU1CHk5VXaF6VJMJjwTgNDWdoChaUSeqV6WrD43wPODBE/MSR2YBx8ip6is
1Gk/okCgslV+Qp90vVMMhaOC9uBgdKU4LJzC3xWON4EzYeJVUw9zmfVy1P+5OO4fGP41wxDdIAKD
w/BkMDEOEWm5sz0VGhA3CnFZw+vyk3UjRmSteKzvKQk0KvPEEtZZriu6SfeRQlwjT/aqbQX+bkRS
s692Viv9r6HbQtY5WiWly21hYYf0c0g3NYH/8ojk9tzuuIkMP+zj/WZWDlU5Q+XPhoCVAroQy9PM
okuDHBPE5AAHbr58oFuuuaAjz/p0SgDol5n3USHdcgJlYKmIg8wWM9P7dy9XeGUXIEZLoo6UeUvi
Y67MhRQX/5YuP0P1bumLodA+UrwY9doUB7EkqSxH5ti5TV6OMzPD3TLZxtTc5gURb5t4hk5TVosP
5wssR4r0met+krhglrwTfoIp+BKz6C6W14ehjJrneIpQ8RwQVszaCH6Dnk/UTwsKGFILjOk0pLKx
WIAx4ERYQPc9Q7qbskItdAvP3RV2+3h5BI1ZfXPm8vFPgaNpjXyxhca5gJUeCPMteZdVAojTtmFT
Lit+kNS+xhQC2C0FHWUe03308RuyajsYa3DmLBTB2VWFXxVN1D8NAuMtVljc+cr0QdXrCvrYtxD+
1hSzZI2AHiLE/ZYNDk/P2G13RtHUv35xFYehSWXrd8Qy6nfl2ZSqoNki/mUZFvH7/ZaStRi6CAPO
ZmPgaj1MXFV36UNdhS4ArUpm1ibHxmVsLlPaVQFMCJA+yhpAF0vxXkZSZTTg1An13WhxQgtn+OGo
vThd5u0BA8gZff+xdQDi0DV6iXNO19H2uRSviCk77W34tx1ASvSzw8oJUEsnmA6taR3ZzXwmo/3T
TkX61JGGHnp4SBhWPwh/bRwss6G5dJ1cObeVXKfooemUOKuz821bvTqvewksAWL3R6R5FmSDCIYu
vlP5DPRyhzbTiYcvVZGDTTB3pJXZ2KQ8tv6FzA7wWT4PDXtFlEI6KPSg1ds1xaFLhPeSoPDN/eZ9
4Btg5II7csdBNbsoYxMFqPtuj/CsETGU6+Fy4TjelVZOOQSfVBCV1l/prDFXHyLoxi3NsT2TFW2P
GFCXHeSo3cU+Ai02Uu8HPM8lDrCRfKQHN3QzocOJXMkyZpjH3T6Wzm/jVWj4W9NRZ3l14FQ82lRH
OAiDoQGkKCXWtYexyPb0n0whnWYQ+PcegakmfY5lgFR/bbsl7IMbc7kNFbBgGYh/ndXWCWXJkV4h
ndEP83FJvjzQsKdt6YMOpZrJVlsK0MiLJAdjnzinnT5CiU6gzRjnQ7KYnR26uU4aQwAH36UUZLE8
50kSqm9g9IhdHcnTP8KPLW83OvfDRf+CM309xKkL4uQy7JwVnGsIixcnB7Fwleg+M2JG7Xh7HCaD
MFlZVHzpM8KzGRH8cDDU8W622hXZJx0NtaXyMuP77f5DB5fPxOnF/pV+Ezvh2enzxFRso0wLoucj
pN4YVYt184JXKJEm4cWnyxGhqRLHis2QGQLpebRyzgfX8abGxuaAXPxO3YisX8sN+cOKQ9OnQymc
ukDwA4ZRu04EsYAIvdq1CfbAyoJ7jABB6qN0aBRpkca+J4J7vPOwlbPX60TmQfWV1X6Xc8qocQEf
mEZDoS6YgVJGm+l9/YmTRVNCSUyFZKeRUAxs5t8gVYeIEa/0U4oZnXd6dC1r+OIQkCiaY5P9mTTF
e0eueAA6htTagTk7qzt6Cm4MhiFEKXp4pNrN+GBaJJfwFjeuRLMp8UaAI3vxVYAR2HvoZlQhFthH
7rit742kETZ+gqesgIwmDRnpSh9S9A3u398fXzODMcxx+zUZsXcLjlH47LWZprdI7lsC1FuWpPek
WAHH/ZXJzZNfdz1k9bAed014lrmBaWFsNL4kZGiZrY+Jg+EAQ9oP0A2SbxrYVY7e2CRmkdXf4+Ed
b8gyxVzF34lvSnQHjjo/+UwqIHUVTfJ89VkjeT1tORSLrRPzflmwEuixIyrIPnqysLUjR+ai3obq
H9RZvJG5jLnIPc7AQ8501U8t1+RDSdK/0k20qsLLNdJJoVM9hHWtVl0hE5SW0YDIRr8IOm7hEwFN
BmTb6xHfjFmB4iTzhO+rW9xI5HIZznvdobo70cgG+NTObkaIj37LirzKTX8uRIVdyzEFslIN+POT
WNL/DmK8waeVZ3iYWHt3xuEn3nMaA/JA1Z6z/tqkW53Dx3kHMXzCRRTH0fInFOFKQaS5Lg7VoKSz
IdgKj/YbiL05dmnTa3yFlYLIBzVtWJriT0m6ot8r8lu1p9jiuBC/Q+jqQjWg9P3BVwTwJwbtsUs9
bSjhRbTtEi/dZ27cyZSBgfLiUiz2B09q8vK3odsA8BVqpCDDJ0C1TSGBvoMkE/Nivm7GAbsiW5UO
PXi1mnfT02m4CHlCxAsMjVuY9thxDVVcejTNFYpXamaFhzSIrXxfVObv18kG23LoQPnHiGL4xjS+
XatrnPy5ErBBf32BXIKEo5AEt2LcEfX9qvOM4gMpu13HJSJw61QLQcz3mqYNeKAZS2YMJSB2GAwC
99wt49Rq1jZwlnIdAT5xXRqCPvuG56cKhRW2lcD9GoziW2J8e0ZFt8VtQ9UJWX9NEj3eDTumBNyW
WwKKXqlWg55uq77jFKbgIwTrWpC0z0Lb6MQC8DQmMIAOsfTWGzX9IkkJQeJtxjp3D1hHI/l0DU5K
Z1v33jhY52KI+0biMRKmyrCWQoKA0Z33sJtV/8uhX8l0COYi9hB83rIWozca4ZbdkrHcSGhojehD
4xePfwPXTI5iKMdu6Xe6THwqeuA5Usj+MfCjktvRgH8uc/KsKWHLpD4UZiOJRtmUljk3vKlTNzB5
J5rzn9kwqgwg4i93qzXuubXHU1TxzMkAs4sEEl7rWVWOdQ05SOjRaAAK7rnob4Ner7/37garQFYa
ri2/nyG7Ll8Axg4OcVLH8x9iOQYRaY9P4Tbl4Hrb/GjnQip5Eos9eVhs+PDfQh4W/CMJvPRZwt8U
ORpvLmfana7OOhAQAYvz2dyQmx1lAxvFGVntoiQv5Uq5ky7OqK6S//SwJgAvLzcg3vuryK2VMUGC
GTVc1oV/pv99+KhXwgaXeu5TAmIVlv1PyU9KE8zQykPc7XBPUFQgDq85DfjiRWN/gUDSn3jWhOP0
krY+I07BGXiTss+Fy61CwwAKb9EXb93vIT6XLDx94rTYb+F1uL5t1W4h5oYV+02T9bkE2MX+7gf7
9LHXaca10zG4Z1WYAzSrDHFIiP2lXDIcfTiv27botJas8ORIwdOKOcFHRSExRMelU0MUNfRprO1Q
gBvBippWG/AgDbsBQqYGUiijV+ZChHANL2qWxdYgWVultYlJ8aFF6nULm/jvvUafZFklnd127oQT
BeHstMzg7nJo2mLwImi/W0txQTZvu4n4jnjvNVJ0gya2qK2LNCWJ7jgjDHvRaneyBclcgHTI9ket
D/c3DKHWtdntD7q8pfcWYhpOLoFRvQF/Zn8NmdzJX6/p3f/SodFnWmpCWPB3APaSzoK0VYcLpmjy
Jny7PKKrkAwnuMgT7gzRD7nndVP/GA0dDOo5KyOQMqt1eyla7BQvSQ56evi+Fkvq3G14Xp6QwH8z
3tEB4gEg+mk+FFTIsgl5TGTWzqD4wqvM0dLWybi3d/ZJjK/dtwTmoo0L5digF4iw/duL5/Ab2PlN
bU8IpuSMQ80WNReSskABrF6SGGuOmWqtRtIf1ksx3Kw4MkGmdv+8P7aZnLAFMwByJY9jSy7VqYlj
Z7iWSV9417f9nnL9Ua+ERSGMDSWGW+Wh2XxTKncW+5GcPn9swx+2cAsV/oNN5heFLoV1fALzX1wW
1sTDmTOvm9HF34MtFDTo+0yKNbu3wDynOIJslVGVvP3Pe+bslMBdZGgF2YMZjP+ylIRuGnJ2VNBf
6OL8QPpP4lIDRazhYmw2zOAkOKxYhDgvvh4PVS1aLAkYEkKF/ArKrcOv7rkODMD+S7Yxd7raqE2y
juvTG9qbnwfDKcZG/EMQmUy8Hj4zLshnh0VFLSmnBnJG0I+Ie4WMzI5IIfCEbr2T6jX7LoJih2AJ
cNA7MDv+Ox5jpu9U52EHPA65fHsYeRojuXLwcMOhVPzwUe/asE94CyDatpV22fLRFqL4pu03VcHQ
zRi84umb1Hu4tH/5IvTLlrfJRFUb5Fe6K2NOgVe282mxTM400Vn0OelokNmqQDxJX1Y1GtSvcjmU
tUXbIZ+P/m5issYll3ezqfJhGl66gHfNBaoXkWkeELJe3PTlyC7mv0eQBM7VyYDEiqxT0EsCwEqs
iyHw246GqW+uOPkfKskYXt7LofeXuVgLvVX0XX1QbX69tJR6G8NOIlr3lJ6IerH5Wv686OdKIdD9
3LF/hlLrjrJld+G2r6ikJC54FMjABhGQIc2ERidZbiYoe0oe+gLwPDAod3Aygra4Df1JCLeMZ8ye
dU/YUUd1eXelRTEHm47SXFpU5cT4XZ0mfjgSvdeEzkqta1WVlRsjm2zXUQr0gCUDk/WYWkilFdr2
L/ZjyOCSZAnGixZiywsL7Ux1Qq4ufgH2RciTQwCMEssFmOEVS/qwQJDl9IxzoBkR4NWmpOsfY/i0
OlcbAsHD2BcTXhdk2TQvDoA4x6mSHKnd5u7rMzu/vtbq6eF/OGzfAAkEmqu7elCkT2b4TTnCvufm
5D0jvhoT/NdtXTAIYh+dsU9DF/+PFLziJPtSHwZ7LHSwK5PLLdLhkIdqXK1nlvoouOciga5MUBuA
vetLvi17jXbZXVO6/0sp/nZdGu3rr0ogOQhl4bYNax2Kf/yHcmP0E6Wn5WYQGdX0eH6UAPvDKzPu
ey9xTUQBXic/WGZq73zwtMw1dIwVRNSMcLUYws4sRy0Ex3MM5cBP9Ol4ClbYpI+CJCttVt0ezU96
NCQsUK8bWtD4R5kqWEl3eynWyijVIkKH8iW6MZzneepDzDWM6jSezjLj7qSlczMJ/0DksWOxftwK
zgJNZqnRldJY/OHr+y8tHSHDOAEUywtWmBT6vMHY0rbtIN2Ws+IxKKRHJmRK5JHSJn88PTgIHRwV
4Ihy0LUA+DfbEdmv/1pc2a30xsApnI4SKwZxd8MSHNa06agIiuHxOUU8XNEN3Nq8tnLUDge8z6ZD
PmXgDI8HBIpc+DzaGLnO63fUTWK6cXjkRJ9WR6vZZXDyUZJG9OO2GBAW0n51Lhp50udQyT3UoBeU
Ku/rQn6ZnYw1YjI2FSr/N5IWbzPTJQS89xIs8uS2ZQAwsxW4f+v6SKQjcl95Uh/PWCNXqQ2mzv15
o9Y6har2UM9pNtDQ4hWoDufPnxFIPSZNi4RNr+Iv86aBm/u1HBOzV1jK9ZrMfGCMkkakxvZmHDyD
+7PU50xsFReNePITCKDH1+PfafLfilgUZ0guH3pvnsCO+9NO/E74Hi/cSc+lkInfhLD8+vf5YJub
SXT8+r305Jnd34nprtL/E7RYCPrZZA8HF2Ebh1MRFM3gUukdQQR1geO3F8OBsK7BFR8uA3Lk8W5C
Bx047JDsQ9j3pbVRlzWUt2YhkBwOz1E6rHDq8nydGJlHKRuZmf7QKuAHo7sTjVqtB09E/5yuqQQm
cpgulqNay6MOlDJnf4OErfzvlOaXXiB5OD0t4oUOW0ccJvU61UbML3W0BlB3pbEeRM/EuN6eRZew
foyO30hIyyZqSbw0C0O57Vs4Oe6aNpLWNWOtvsATPggZx1TxSFWzO7ApyFZuq5ZjqD2581I2OAwO
i5ZTB8BP4DdU9lGLhbYRrEoamZss8dRBOkFCJD3MO4aggT+Ttq1vrLUsm7y7nKMag5jTfTx4mr8f
p1NtOfXzUSLhyznmVEcjRx9DiK4uuUd/XfFou0LtdmuJ0Dk/Xd11XgXb+6tPLhZlX99M6w3KyOF8
BolOf8wWEaLcS1uUnGsXIia0ZjwsOOJhA7bmZ8Wwfrs0Uw+8jak7nckm9G7scFtVNKk07XrFMZ52
7TEiguJP/igKrd6nVCW/9cDVGVCvAfpR6NlxXqBo3YXeJaTbfCg7NL65B68S9DDdG7YikiGPikiE
C9WhB5ca2K30HCW9bx/1BDHZGfGCsilUhWyM5N0tXF6VFXGNaF71SvZeBDM0n30mL3RmCTYJnETn
z86gqShtxp5BMBf9BSHiFteAknDwD2bX9gU7VSl1VZrJ5exqxDTNXaQLwpzvnoWNHhaBDQEsnng1
Cwx8YQbw/5LVOOFiWma4Hv50m5F/r/kHsqSIR82N5qwIavsc/xcfaxGzhHtGqqLJCvIqKB4MiLL/
zjjzt7dcpO3ovWYwzU1qxTzcxltIhBzYGFr1bSOArKFjWVf+KweVtQ3vi5S+sWuk5JN4r55FFL6S
7K/fNx1mm3dnyi6dTDeEtPGmjjgYtCvNeU8FthgIZyNp1203uncUuVsB5W68RDfqHfudhzuOik40
T6WiTnzfcEeWcFBWDn/EjescRreh5OtRhYmp7xYyC9/jFj/LyiZ3qU6LWaPgJfn8jTAkhcq71pq9
RZRpbX0LGsUceO7VN2j7RIXiPB8Xp7i7Z7UWFQywlsJRqNDi2H9S08aDXeOpxGtDyJi06o6krtke
UYnmO5mTFM7R4acxsd1APbqAZkh2x6Fl/8dAIA+ktPjVXCXU54eLxLgqrN6o1oMYj/1z5Y3kXjQE
3qdIUG/GRFYUcFLzB5682vWGXHeOF1KwweewdhZWfmDeafKzcZSMmKZFuWrw2hjPHAyFK+GHQL7c
g+ZxFXnhxBnqMlTKn+yZ6CKSrFtGDqXR9mZsyJ/TJ9zkEGwX4IpAdG6Hqu4ZaupgzHD4BKrJR4LN
kDPzN32UNgRK0JwOaToj162LLJJ0JFL79DIVaQ8dgyRfPENpKbdr2aR9p9H6JUGqkWPo2mVbT0eD
xZh7+c/bhTlmFsuN1gaLPNec7QttRalZ5PA7MbvsJn03Xdyvf40/ONZh6/Pm93t+10KFiOKJr3ad
riPOImHdiyoFkALcU9zZEotkcYQUJN3mM1ZVTB9E4z9NAXVe5qgSvencFmuOp8wyA3LPL0NvCuRA
/Bfikj9BpRC5p/MpBJ3uiR2RrF7U/JCEWhHbtA1BysKJkcDY0lor6mQJwMyKNsMDa5O2lAXcQLRX
qMFB/q+Hj6eTdgnGeAIe5VHeW2vcAoI4i/5n9Fvyw860bV9vGd7uexTpxEwj1LzNXl5TIlMwJHkd
MxBx4wYD/E+vIyrFCZHL5y1xTFiYNNO+59rp8PESOMRmdGL0J4LJLLz7x+9kowRe0wFwzqUMR/BV
c0MozOo8A53yqL5bBJeEzMsgbuop+S4Eq0moBG/t1E26eVXQBSKHvff5xjy34FDfF2AZsAFZci29
GbjYLkZUw4LKqzC7di/7rdVhltxfeNMYcI5mF5oTBqANYyTBnJV5rO1liptGn/HWAWlGw8qzv1Av
3YcbR2tI4xcktNaw9tpmySIGosFQ7PiLo7Z1LedWXmsBCL04yfDkKwbMdiko9zeV6N1ixTQyZ++Z
f5qMy7/zfIJ4pziQxQbRL1v6uMyEgnBx0oSKGnwWnUBtBAGH4xDui4gpevDKlCyQBBLa8DxXGO5y
njXLKx4iRHIVy2HmVjKroc2238Y2t2QMbvhhflR7bDQ2TVyidfqxXgkAUnE2BeII97KFcMZq4Ltk
HL/Cmu918zm+hM018uf0PmdwC5atIF2fDiSESe8gXd9nf9Jwg/QB/3ZUfKswmFRFfJ16vKTyHgxO
12avmrg38+lLNO5fYNqcjKDEFRSEjHo5mhPw7MGYl79J0k4OGDHxsyuMLzIITUbtzbBACxU/X3J9
wI32SXF+Q8eMc8Z/wrSSxJAzWOj/3D0RiZtZVScKs8jeOLzw72Sa1uMBkFq0/JFfsGGy8uOEhcZC
r/fQsxrWeDPgObHpyBcBw3bGcJzSAUWjpC67eQn0B6m0q7xG4kJPgQHs1Jbcl+yOGaA3cs7Vi4f9
OYxfjVRRMjrxG43qh5lTJ2BsHSykt6ZHcYJ4BfP+/6NxzT0GsmYsYI9lV7EdPwsaqO3eD9S6mZe1
adzKRa1w8Ijw0bPkEpPwCYQ1e0GEEPpqSzHm1SVg4brLugAQ9s7oN52XMlFclMAKYx7Gj0xaTJCg
jL57/+BN7awDWiqkjsQOnuHl4yekcAhUkKL2a/WgPTttlEgTMXqwojB46jwR6iN5WIMVopwtSamC
m29Col4f90CCafcrgTChVJt7i3GgRfGJ2kO6WvAPjvBXLUmAE0GfWy5fIYrBNKVJ4A12NadK1sKO
0x4CwfQlQw6CIBWI1MNPx8DwbXOVVXzc+nlTuu4PDhbDmux8aOjFQmZoFBrrVTpTffJblhI9cjUs
6IPq9J/SCnHTeFShuX6D1k4Yfa8RZgYx5gpYhwyKb+KzKA6nWrVH6FulYS500nVTJ58PusBNSVHl
J1hrNvp9lUb+i4tPMvkeDv/FQyv+XaEuoyzg97vDijaNO1U/7Yh+RRtb+GrcaeJCgOgBd9QpmXcd
GiKc+O3hdYmth3lhkdchAW868DJBTKz48eb5YXpoNtpu69f2n87v9u9H8O0RGpPKiVIUqg61oJRh
ZMfpRQT1ytmg9zzYrpvYVKLLF7XjhZ5C/A3so/tXThtPWW06pnij+scP8+HVZtJwG8VidFPkuB6F
wdvLtEYlXlmdzSU4fhhNiM/LkO7ACEf9iLDKOeqKF8GjS4s+AjrQbDuFgoWuf5gkG72egPPxrt2Q
5A86121ma8T6z2ERjh9Z7FMmYl1HMmVjkmfFONfR+HlodIXxxIHLyL9z0zowNjzN1PjOUeEa44E+
glYn0Q0zanAKEgkmazBCuuiKIJPyBllRSalHpUh95Qp3GOncVD/OpHLKCGG6O1DAx8+CkJi4o0r8
Qr1DfIHuT8OmZGy+Wn7v2aKQia9QAuXAjB9FUexVGMsCQgMkRnmFZSyqZqQNa9bjzzlOnBCYUq0y
HRgY25QBga54VXbvmIbhpMeyD8xRAoneAien4d5AcU0TdwgAb/BGGVJuf+VqM9ChVas7jJ0AlFo/
HRq8kj893R7As2RLOHVB8P4U3awj1Xi3p0eTfo0x64LF/q4tcpPjsXqahEoOcf9P4YS4KCUXaP2J
xocz6+04ML6VGU4t/XVqF75a+cOBhTKeY1MyYeCpKZsckFgG8tSyd3RE8by5ua/kV4d7nwKM4dC3
KedeNGTii7m7xkAZpeh/SFsjAaAkQ0Mhu5jcIx08kXLX75QbIUDM5I0qnaM2DiXGQNp1X0wVA7F/
FXgYeqNOQ6jujgLXk9IZOUcQnMtKmUl26F66nAXSRRZ906KzAknPJX/YUvahHpt4H0e8zzCTQQjO
R/pej2vWNIYp/DDYnxDLcrcXS2EDQVI5/CAMOC0GaD0S2KFOUCRJ3V0LdhPDu21vCsPQBFQRBJvT
ZaM1hiiL7sAXpkC3p8URrBMGFnOyeNPooVvHkeLyIBxNzOTolur+tdnWwbzm3eyxpx8Gyq0/GzzU
/GpeYDZfkbK+g2zJSyNWSSmRwZvZI76vwlhPUQOG28DvsgDH4lfrytcDg1Cvm49w3HbT+jWPg4bO
xOmXYCs7ogLrVtgKjjY24laJf/9rxoqVXgds1J1D5s6KPyT1XuQo8PCMDzOeQpBrK65o5IVIAX+E
R+jnO6Y4oXi29mcJygy3AYagY6pgQ76lr9Gdz7aDA1wyHGNZYT/LzVCydPQktjvhPjCVZiyDiuhy
LSBxgbOud9ys8dq6Jg+C4cp7fgbJJNKQDOGr95NN1jpHyTAcvKmZ0ncrKMhe9SoveUK3gxU/iyEC
SiBAejIypBA99R2SbJoGPRFvBkhcn4vNidz7AMXBS8FC7zjtUKbSegCq6OMlc/qUn5/viKxkRVzc
s8KnIRvywhEf5A3OYtZlJ3emX+BWE06KOTMq5pG35URMCf+a6TIoWRrtQOKvryxYjZR7J7ynjuDA
16gqCKaAHinwGyaZSijiXDFCbJOomeMdgnGC55bdYA75Xh8tyJXkFmsogHRv4Apkcv1/ceZh9gvD
ZMkx+/VX5JCVJ8xX1F00gLIynuxxPwAuOLPb6HdXfH/CZpsUBqWKy9qqHpPj0d0lL/w9Y24d3Xty
/WIv6lAyQ12K2rCslL134OzsSS5qCguu8uGAaf4X2GtUdi/ZyJbTqmTA/j/3puyjG1CZO7gPPVt9
giKdaOXIRY5BCPbRBVsIXzs4wsxkFFJ/kHKadPqcpZmg+FVfZ3Cc2mc9IFMrmeYzFNSsNEDU3ocL
eX5L3XtMb1mehsxhVtWKWu8rLr7IQaFAfjZ4bR6IjBukhlZ2czZdPMJvnvX//ULL6trmC968spSw
HzCWdyex5JwERonwnZ/vFB529Z/QqcxBoQoFkkblKJn/Rl0CohAbmI8aHHek0bIIOiJYlcebfX2s
MuW4Z4ZYwTN0UwmooIByi7nPtWouKgvJgJz7jKQb+O10JWCg3RFP5nymuSIFb/4SzYsqGqd4A2df
bGbZ+CnnTWT8YgakNxHouXrqwh2+7Ae/86hQn/fXikmSMy3CJUl4rh03VhTQsOX+e/ZVpDGTu1Mc
v+dmjXD0TA3NT5XzT4HvYXTITe4ryhzniTt42UzDV3c0r2i7NhiVdxrZ5THfwLyvGepfkGAcSVnB
RORTVIKMFaJn/TeJOsVziK8gin3f0ksmo2kuiHzYFXionZG8G2Ybgqdzqx911tBKgKuM5UHj6i9S
jwVI76sv+Mht0wc0ovYghOhQUT/liEO8/AeFMhrPeiIpXBk4+HX6KEh0C4praaWdG8Y8Fq+hEcjm
FbRek1NXAaWea1BQ6bU7pL7dIncXld7Xetrgnb7tTEu70o2iuuLUzmgfVBxbsU6SBTizyRVKTdWP
E/WVB4njIQ7jEAyqCxzR++/6gx7uVSSseWWrnClsMEflOO4GDd3I18G1CFNpq/2Gw5P2bwGciWf+
6+SS5+2iRfUS5EIQsOaFMXdxYDvk2MALw762qpS5uvVp9bDN25uq21Pyh3XlU4tLu9C+z7cIJRTl
+2XTnkpVwDNXwCRrkX/jPwx6UYYHMBZRYOe9dm41CAJW1AnFWMqhF+GW9DJgweY1nvxKBMp3YfJn
ObUmjia6vYoYqoqcajQbpvYg9fuXcmK0l7f8YBmUMkXxo4NGFraHkG3/b0qhObpwWB7E4IPp/Y7x
cwJAeEeI93s17IrfM+nOwepLgNX6zyULUrIS1s/HVnvY1Wdsu2+gyhqGE8dC13yUGbt4fog5l2Na
G8O4+2ByXIS7ekzW5BVat5Siy8RkJ/WVbuLDjZ0J3F9x2ObohJO5Qb7bM5wcxKPmt/mlEBSfYsjK
ZaoDidhZpZT1KCXY8AQqos4o3RHhLKlC8J/zaX+6zc914hz5ecFtWYBhRtPOCyuZReyEB/h6ozRU
XuhfwiuC2Kib+FWmLK+G5doPdKj47S8Fp+D69kzsEzmVeuFjK+iTQJyNFZeyanStg8DifxqNm/Mj
JCjLMNprobgDfuizfkiQWXgpDG6Y7t5K/WsLDfrRhsvJwTWOn47pXBVAt0fIc1z55vbnYt3/mX85
oqU2r1rihAINq9x3YxOwqPAQFzQCZ7cImcw3j2PTE9R3RBwFN1abZUbNJ/+Sm+LabTkx4dlykfuw
C1UGlDndjCpY2rxvo5pkU0k+azg3KMb6yVvZN15U2LQCAocrAiotKAE37+VxYRMrsaVnMKO6GXyP
3Ik4os1UVppnd/NX33lyN1ULOvYf5pWkVfK/1V49pundYPbJk6xtBvOMLaQMzOKurj+mC/DkxUXz
2Qxn+jTyw7V5zjO3BL8/RUd8IUGfGAtvDYJJIpfMIOX7T0YFYLgLpe0Gef9oPc+bgqi3hLwQdpPW
E2L5QgCjradoBnpmGun/0HNfYLjuMpCkyUpUrwSihcdShtqiEHJwzP6/CYIlrlI9UiRJjt+V+U7p
BphyN1WBVWtER6VF6JmbWcP4WBlbt4ddZ/nlH4NSpD0xctIKVhqucTXZeOW94Qilge1+DgVIse5O
weWiO4g9TOaMW5rwJlVmrRPJmlFec0iL8QAokVDGz+qLew5IrM9dHb2mGbX1BULuGy0bp2et/k7f
oLVLrWlbm6GZu2oyF3eukLRnAGYpYOnNkBEZ0iBgfWXeaMSdGjbc1R26RcPyI3rBEF8KDAslQPdo
/Rcfawhg4eKv3AsKR3eDPLeH43N6nxSmxqG/2Mfk9AzUYVG89z3mzW9iK6o9uForDrKcGgqQLwA5
qIHm/b8oyXHBsHnfXQHyrVcd1WO9tnHZvVX1V4AUIABgnwSVJhUF02X2SVKcFLd4ii0r55biQnAb
MJBaTbpYu65sBstSS2u0/CfXvgzbqNkyiizfxSqfZSmjPapNDwLqZ4sK3RRaaDrAscrcGORxiFdq
SqJ6NT6VhH58BE6QkZNt2MA9jG+lLsH9OqOx37YSPDs6XDf9g3tP4PxGbfKg92vZjwEs1Lzc9+Rh
78RHcpe/QBN9eVSTrYV1f06AhsHjuGyLOEjC8h/ir0yYfa5om/J8qFHSWXDmeDorcAj6xr2a5A9q
y4LV50HYguSEHcNh8OeeCsVDEC/UMj+CX90cNFvLFbRYXtrjUAF+g1jmjLjCYfR1f2lBDJyG2UFe
HoW/jZDU64XFv0QQOqIwRdM5SiEKBGyPJ1iarbuXtgIoTCO4DY+i0oNZmbiMrYL24AZhrAthVxei
Vyn/XobsocpMQrVtgbtcyxYrHIExrWXmQ8QQDu5tZlTgVi/FDE/F7+Zno3ertDtnTLzgeXp0a/j5
7x0YyybtpfDTbQTuBXy3PGxlIa/+/BGPReXTHSSpaFG349u1NL0SO/mmEzPWUd6x1+aTHSRUtQDX
n4P50K9ri7H6oH2JXqNMWLDOlcanrD724PjCVLUW7l7w3Z14SUiYIIJQ+QbFzWUJdOg43RbLfV6O
p0T51TGZWoQwBYIfyW2pimZZZq/EbqZlqdX9KGGraf1xQLgojFS9f6L0ODSOXA5ksW43kTE6wXr6
nwRwj8Jq1wX0isaj3wiGlBLB7F9uz/NOZCDz9I6QReew4yvuOe7kIPoEoOTxSYzIK3nu2zaRGNyo
59IPFt6Folz19B6XOLiIu+mznAGKRZoA8BZlM80yGAPrLNrwhoUUSuM0TBH/kIf8WKDGj+AHGJEA
cn6mCaxbfsyayeJFJhi+0JXi+Jkhg7PJ8cBBUJ3ElEBVTX1uPjfX8t2EHZ4YRQtMx7MAA63XnCyT
oePXtTtup004DqbCfKmYByHlm5PhS6mS719WgqeazNxH1TasLVVJ8eZVEF3PtwP5w2iq/j4I7LY2
vyVRFX7+KCLrT/ufyIm1RCpL4/vKB6tE5K12halywEYdUM60MpfiwQDZq0+zS/3b9Qi5IUDYXVE5
DygnYRY1Hzg/xLk/ItgWci3VsQB37b8qE1GQgNccZWKKxKNdf8qZ+F0JrbR4JUSnISH/pMzkcBkw
/X92GU9GDwuEMa7YN60nVg0AHjPPs3NW4q/Y4Ev1j3m+p6dm969lbBsEuNPRVyUOPgO/+BwtG1KT
JsJLAljy+UnhkigeAHcY2pJuQKcMwA1d+vBGy4kuDlDLwrlw4JeJm+qPl64BN2CwYumY0EP2Cc3b
5tJVPVnHpXPvKvrM8O1Bbgo56QtBxfgYYGxAVpKlXM3naKM1K8s/YTiL7xeh0pGnBcr131bO/Pp/
NpyPMLD0Wgl+J3DuwNwy86b2SFNBFsSxV1x27pLfZMYFVphG1pZdlffDoHCLbXArW8tcivBgkBY6
Ci9ZoT9vtU/rtoJGokqdan79J408/WqLXoX7MhFk4UmvnuMIUPLXrbkmOV+KBcvaLGe8BBY04WT6
qF/u+zdAw63Eo36SKmTy970hCIlvfSsdBZaOMG6zcIzNtD95B6agkjj87OusH7xzJ/+d4QCqa8O7
7u8ADlSRH17HMKbKs/cD0Y4CpmMjkdzMCHZfqEQWY8hJezp0jazSe2Up8eNi9+Bny7xv5RXKnCEp
jSa448Rf9xxrOXK42eLIcGljfE440s3B8J5I+cfLgMQTiUvjDVBj8kTgapocuLaXqMqyXRurn32l
xCgb/fZWFdvWHqFVPJiK3TXdKF54RqOeP6qnqLdaAC42N0YO5L6f2DLhGWGrfDee+btFLpG5ZjO5
mDxHKpc9Op36MmM566FLVKoG5Etz2MQzkaDllLRn/C1XauGZwiepQ/JSM8ujiS4JaKlZwtLcmI86
3vLZdgvjc3JQKvWa2NsFknIjVRNIS011ov/k9H+afVD4ZvyGtnvrey1l7J9Zt8SITVQQ9AQLqa3M
y3AI/V4PyEU/CgOguurKsMjbktKv/Oh45xwGEuZBC/UcyN2R+Rgr9akrFPgPL/F4nB0jrcVNVjyQ
Zsqm4c6gydrKDS1JjCY0MQMj7hDjMnzh2tpAHR81wyh6KAyQfv0MhZc/29OaJrZ8/gD2tV2XpKzh
CC9eVdxEkDXTEWxtqPRhx4GjBe4WzY3AsO/vhztlESHxsAijQZys+Xi/R/pRlprKLAMa4qKvTf6i
/PIquy2lJCrvPXvcZkRlyuexr9Ft3yqfxoUGVU1dTKTLSz8eMGZPid1E9UAu4mududFFC2z4CyD+
MrfQe+Z0SEaF5bgSX3O9WjMxOuoFA5ClVh0XaHQcIDqlLmfZqFZNaf7rEFcV8ZVRKfJkc7zZELt0
0LzM5Z4tqstCPWhsGUOIN9xJv0lG/GcITVG8nzzQ6KJ0fdxG4U/6YTgQzbn9rBAXJQNSJIgctnIJ
qloIOrE8LREJUvL/zOJMFj+zm+siqGGlXNO5+daA4Ib7ZYyhMB69zBcKbdqiEc2k0SNSd5vQo71E
TljNO23PmNEx4ZMxfFgb6hQBLbY0NNeDd3TRmhK1t85jXOlFryEK//T4tzFTbn8q1lPMThcE8Xff
3SXm4PBH/dE0vG7WcwRMNBXwdoGPK8bHXm1ijVlaPNOGmMLkZpiN6o8ZDcz+vzmjEdAzX58PHybE
ywlgFvR32TykTdUpAz7NHTaq7aCbpsTnpf//UpmJq4v6kV2HIIVDgTGsUDSZKpARJG5cb8i4viYx
N26ZEqHBSherbL+36YrpM1uTgnNaz8bS6xQfCprKDr6ZGhXCcpXQwj682qUTlxC3eItoxmu1PR7z
/9ca9RvSDEgkFZ554WQU5kjU65MGZbg8PN8oQbP3OWz/Zo2lS60JHqEybE3/oZ37isk8MOvpRqZj
pZDEIz2IaWiJ+RmLNYVzKb0sHqOVWLOmCx3+PiuvSpfpQcUZiL7E9bfa+X+kYtwE0zw1+h65yfRh
nEhmo7TwgyM5RSw5bb0jSjk95fOH3u6ziNO/3gV0ZYqX81dJA6gcdN7bNw8cG2YBmtJJ0ydYALNy
O7t31OYzMZOkPk3MCAsotQBT3TTxVY2tONyQFfeKcAeKO/d2u9pvAY32K45M5Uz9GswuaofybwEJ
ATYJehS/7B6Xpb9Ql4zOC9PW15axcBHNJAF0q231TYA2xBMEdKfshqQ1U2DNjTKeGrOCvgqRNoNs
I9S8gJ84XCDao6uLJpDzNbIBL6htw6hbiuBHgDH0wHxox+Leri3DQ///+o5R96AQt0L2qaqklwRC
jooW1tIN3A6mwd4S6wlPI1GT/5GwR7xki/DkjCo7tQQi+ctoFtZBzOCNu/5HWL4R13MAestiNVSq
zHhjY+X3pNVK3LUbXhOsdbnRpaEZjX4u18Fu2mla7fQfoLJ0ClPIGlDfyWyYAvmsWl7vBArihBRL
O5sPWakL3jQeP69xTMmICWgTprbvwyUae32/QGsQ+azSNhD/X410+MWU7uO1E+AhspMMLIjE7iZD
N89q3ouKGeV3hbbrA/lDHXadXsK/M6L7y4GwhnOUnmL+7Bf2b7orLelMk7x4Au/LNhIkGCGKVhLE
4ASoIxucGeMfiHtUlmSOYvfdlj5uexyi99AiUaYRuAXyZmJTtxOkJZKInyd5Syqt6fW1aM82+QM+
8OHfA7l0WxarPNMAcMZqxgzPFLGJVVdtjP0z5jFacb39vhiss0R5RdPh4XDnVzeWSWZPmRnNXTIz
Sbiebzpaf065QAhkTHucJgCSHIKUqlsFRQW1g9trjdUQCl4cKPwTfH/r0AbpA28kCmvY9sd2kJ7s
Okjz97ewTDn42bfSCN/emMYqJMCgmT8AXspEe02Qd2W3KRMlq2dKabb9PzURZ2RH+AlN1JmtulCb
MejQ+ERUP1VxKYkB/X4mN32E2W/Qp5ox9+N0uUwl3+cQPZXIfS11xd59lFAnVSrPq/q0w57KP7mb
B0AeuO7Sq5odXx7MSYgjs48c8MVdYBmXcyeGc0O9+8RyhLqvqoilQTLYFv10+HTcTFNXHe+oE56g
BjEP2xb4RckhZLcJVWzBtMOECWfmOZRXCq48A4fcRUkHOlDGnphdxyVfN479QCq9AhsEWvxgTgMS
ufhTRl37yjSbSa+Ub3C8+IKazqsQcmfgqySWQ9gWUOJddTaf7zopcCIgvoWS2Pklkf2in7gVhXc4
iFbqc8tBMAqJapL4P+RWrSlDB7jMA1lhX+5Ox9X7U3EYdFTPHcDFz0M/c9Ypzw3BVNlriOr44Iq5
5eisngJhA9vopqWDFZjrxK0EY5h4kxyNF07YF52uG/cMoNUj+Z/S96sBWQ6PUtHBoTd2Bs7E7fQL
kWqGhg0pPJLS+02Yh3N3Df/1vmI486wIsqSJF8c/mMMoxonpuNLx7LK55TvUFogCZaZkv4Wp/zuY
0zAJATZ/TJmnzIJ+sIL5MS8E79Gk6tvG5kVzXtUIoWs2FWl5zZorveU2a7hS3sPVFeVq4MBWiPm+
YjXyjVoj3swUCzvNYGld5KX+2xfOTaKCo5PD8LFCt2YTVrAZZnghrjk8wAjdrMakZ1BYIgO0ryrs
OufLUUNe0fdDC/U5iQyjYfE3w/8kW/PXWeXUV2tJ4zDnCR8x9NDmJiNBfOvhLrpMl60yJcThCDlc
5RfaNhw4mcja7pfl7TqADpsFnFFJG3uJKRFYBh015V/73VHR62/wIpQhep6RPBmOWZbDyJ00f0aN
B5bYjJebG/1QwBhex4FKWesebV3JylpBFIyv1tCqHVqsJmaYi5db2Hekl5Q5owHbUxhpQw/qraqN
1HrjCt4slCWheyDc5yn+UojilRxqhUKw1jtv/XUI62EdEgTaqx1FAqn2MVtX7tId0B42IuVjsk1B
VRogQKGKhgqyztLL9svoD8p3OHH1g2BaNNPtBkPrRX/zEshHZQ4oIUlOqngobc7HimOXeKSxr6EV
Zt3OT0cjcsIUJQ2uPmSCDRkgfb+A9KEgEiFmsWvx+FoQh2YDAituWcgDR1+X0RM2T1ubL9c0IkP/
lPMVKXMfcfpUw8cPVEV1jmgcXRxCUWVplA6YEC8fZPzah6ITrOqQMjyrrLS4HLraZAkfXWY4IBp8
8vQwt3z/rvaDRvjVgs/TqUIKLRzteG9sVNFo0AugVfh5HuQ+4pk6Q4c9JGG2mYTPjGlV8/js7y9D
aQjvy6MHY61QXhhGiLyZwOEpHf1pUHO5DyYDMAqW1vfTzynV7N13Lg7d+/vP4w64bSleBOpBJ1t+
KvhvTpGLerr7Z/r5vTZxJCOQbJNwsawlPkEBFgA724Y6xd7Oc5EGT3Fg+Hf3LF0A3KKR/Lv2YKtM
XfgTidbxIzQHs7GIJYPM72fEKzE6O6ISZWPqbwlQpt4AZUuTEwhHhmYgvXKfmTVArVUPCZaxkYRL
KGC7A3/y32mbUnpdUf0CaqubEhvAhvl79/YvBDgBm65zVWgukokasdCaZWG+a1qPDl8JWQZXQQ9I
ZviJgno7U/VkpgS20gr6L4WJWozmc0Jfc2gSF15W3pTRk0apUG04KNo3CfCQGS0yCFpSg5fV/mnq
8w9UQspjkMt1lNLkFQLcrNmVRN6K25Pz3yzP+S29LrVKKojQcUVGGnUcNWBhIJe0G2Bti3N+0/8+
JUA3St5kXw1JyZsCUTzbCSsZVlvsG97xx2Zm/+D+sHNiD6kZnP7iTLyjn+UHHB4bCHGLJIYTFiJC
sFH0zOFGrGSPPsd89DO7Hk4N5GxSXBteocnvxXEbOqzFkorEMZ5OBzAUvZgg5+rTe5lgZ+QG25JX
0XmrAytz/0FIndr2zwJOGkiJD5w+Z4f9Fuwz46SN7OnYtMOphmGl+m2GydzA8CBX65C2DcXFXEC3
KGftnrcOb070OHUpL2Rq4Q2D9TPSCsjp4QbnXFaLfrCmFFbDSgsNaLOz5hVUz0116DIYKyRZRylv
Bpg+DnW1hetYnOYnn7o44vc8byr9oztA/wC3hRz+XyHvECXq/5s1efm3OjoG9mcyTXIAH42xg1RL
QyZ7rohwGTlbL/sE3yqwqOgjDZNp5GerRNCJ0iBvExSzg0h0Lg5oYi8w9GCTVQ+zcEv62Ett2xwq
Q+VqCms08bIgrDhznb0yfFICkgFUTxYGf1rPW6xTcRwE5vMZpo91TGrUMuDH+yjVNVDR0LcwTGYw
GsaSQoVva8Z5sToVjpn+Kj4mcCfKxIzuAaAGsbM0gXrFJbIo4a/Ur53Opjq/3bHMhJvMggB0YwOE
UevJwJn7Yn0kmaiwsiSlsDgSwrD3chDwtRypvnsOWpS6Dw1sRnDel6qQYxLrkS5Spt/vJ2XObcf0
kj9kbO1b3dKSfwOq4+HK2xjo8/5Kdy9vcJl+yyc38ATFS9FR14LvyDPjFYbCTMi1Ao3w6YqTdU35
MLS9wE+oVKAHR1vzsS6SFpnZuVdwS2QdmKgYESDcL9v7k4UtHuXYwLH52J5VbaLjsJDg5k77rB4n
/R+ryHoUWhrMSeuXzj5sPMSGv7qx4U5QdF8hY4CEVYl7uWdsGdUZI9fppPVokRGNAXsU0OvZbTVQ
oLm+mJRPfjwluxlEy3drHVEbIAGRpIkOKKrJd4/x5tqA3XO0sZzOOdh3QDhv5VtWZzyDItDTyWpE
oOmlw/sGTNKN4dq4s3HUdjL6MstjntRR47x6GrpROxGCKBcEO4kMAk6zJtQj1ConH0VgM5YTCh1x
4qxXx8o8Ue3ryISxFex8k/WreZTlVPvULmABAg1jqKmIjSrxQDyqZBmd141Ue325zVRd91uwDuuX
HyHfnZhpHjHW0nVc3la6RfPwTYS79ju1cF+OXUMVMThL/wEWOlt7sB4H0cvUncZhEpLoZ7iHPTvz
CTXMdVKzWGWFytV/+oXqjgOR3KQ1fh0tMV9zzhIt3TjZYhQNNlWkZ8W/sokJ96P+rruOi+6Ge74C
/+Fhkv6ozP67Z6/lhV/2AtCMkbRJwmFvS/XdfrIlkHxQsEZieX68j0Tl9l1F/dyZtK5olm7s9mTS
dfHyYcbC2Bpja+CXqNbzLe9dHq+BwmpKEvYrEx+AC48EULFeubJQzmgD/v26NL3Z662JLf+c1bbx
dxoD/zfr9qScHuQF84RJ/2WIMGsU7NjIJoZW6VT9t4wdewTy1bG5HuJQGDCgZG8ekDkBwXoHTnLW
vW9fRNwLwR2wNl02iG70pIeSWWNAgXY1buwZDWTLnRdAssTtXL+TVqC4yk7usCGKXTcVuIxvXVlL
GZ7SSocVtrpHymur+/ht/6p72gRqO9jwj/dbd9jIojtAOvz9Syvb9zbmfpSfC3Z5FeCx6XGFgUb2
TVR/mFq7ZpBFRGiZYvQXXZMajgX1Zs4buhICD42vfCx3lKuIPneTP8OixczoG/U27LROfgmxeGQJ
JAfZSdVphVut5tyeL/qBW/HXlzlcp1bS2aK4JDNDyOBooLeKChihAThTSnsm45T/hvsrHmR0jKqp
6/wYDn4VQL6GP0/04HNuxApQYvOCP+SpEvDjQ4YL7COzpQtZJ4eve7IkWuftPMjRfYUKuU3a6WKf
C+0lM1fFIxL61bE+Zf2L/R62K80aiJxoxdsv7qk5umqeS/8Hzr0ci56PQpPwFFvnxFXa4iRNnsYj
ppzp85X3G3Lu2M1rn/63O4sEUi73V+K42D0VjnYeeQcXK6rB+4tTkwXNXhm0Tlm5FrWbNUP/b8+c
amBkKlUrBVIkgxEr8gcXvFYWblI6gypNhz1vySdUI33Cw7RV1bPqum1rzTQUHolBO5ijDyX29o6J
JSCm/tI4AYDqw+J+1c+YQldMnwaXbfLzxrULs8GZBVqA1dno6O1gUxjA8RF4RsYTjdqwIhOlDOvt
Sv6LXA/TCKFbsJyEfn3Gad8i+iKe0lZ593mL2VAvuMMyCgpU3Wo2wxFGpvwhFE8C8fMiSKi1T5H0
xG2W5nX4rptvAJhXBVhdR3Io2c+0sDwaE4wbA5dWViB3/eDpTItqaKkJoLSGGb5CnMbbv+CBOv8f
KR55Xcb16ViqQlS+NGGTTbcyg7L+qQr/8YLpWLfINtJ6AeC5kbezrIPKJxlnf8ryS+glsF2WsqbY
3CSUW2OweYHhtsonkQI7iO6q9jMJvOHX6Sm9/EIqrg77NqFRLeuQdpNDNO09dlzQerGgVNEMZcXa
V3t//QMZorrwHpwapPat6MhClYkStNRGM/yjqU/Xhk8LdKsk/vMy3ZIAfaXXTe11Vt4vD2IBEdf+
IU8vNi5UmKOvguYRU78O3QJ2Rf2iLLgHAh4pCfXzjm+5mlv/xToOWtOkArr3uYrzlf39hCCGz+H/
7zzQL6WI9imMlFRFVSN7ZNcptwONLWxnLrwCDhUvRO1Xs5bQjXfrzntWx098kxEXhih42MNs7FjK
ARmW2gUVb6LWntPQJCwVnLEMjHY+YXFrbbbRAqb2PCCKeRneSqJ5/fmRMP4xIOUkiGzD0XC/yYkc
ad9hpJ8lRHYv2zw30LuH1FexBKQHMtZ76uG956aQ97nQfodSO9K/XR1TYVinHyC5IFrB9XSkaGg4
T/AAIRazxoAYn4j/wSLgSRpxYACRE/QI24N3Opi7IyEE7V0PXVGLnAbVvK/u3oU2WCnSepYML3l6
6VnY58KD74482k2FXSR3g4CzgZxZzsb2rGVaGmsZfk7i0x3xbdLJweOF34UseLCItqaUAbz5zZza
4lFHW27Pe6Ae/KZWCvK/c5hnPCeCpx138vjbqeqTAPCwviGbi1K8geom5gHk3ixPkC63bRvsATka
PNtpQHrIBXNlizz4TsexhrG0jrvfL29BcN/FeXrc+vOg4aeqOBymzy2HQAL69F8+ancS09N4vA17
7y/cqM8hAHQRoavPfSk9Ws9KPG/5JglRsHr4x5eXKRs2G3Nnl/TtHjLlOG86RBNO39VI3nhAonij
JqUfTb2hl/gCGhEB7UEx1kMIkx9u2C765jg/9UZPtw7b/Cjvvdm103VSHGhpNgY/82oTa/RsDG8Q
M6LU+lz+ySW9BFyMcbjqYnz7N3BrmH0VBfXQeWoo+N7qJrKTZWElzE5d1A7imyk9RIZOj9m+hw/s
3nEgsR+KHy0GLXzpOL+LjzPODWcJmSFm2Dqxo37TZ2Kto/faMoTOFC62hA74OKLu5mt33e4Uqcar
rMYooFg3YAL/pQq2enWdVFXmqaUwLv8K0cqfN+ERYIHUGoU1hOFFXA43OVAQCkn+qyyV/Da1T5/d
PA4O04o06DxshZpbyrXlnwOgi87uTp8rSYv15nvIfKNbq53RaMHiNhKX4tYT3ksDL8NNz4hepIxH
UFPedjHXKWUTyFlw0q0tTZC0i6FjBr/+b1f/mIucnZtmVVLIkphgMrPfF8FPrBJ3WcdSYeNEb4WL
Wsh7xIpia7a3Ktr+7DyQtv7gdht74MQQsuayKeKONsl37gVpmLA8S/W4q7WgKjcy2fKKw3Jlw/TB
/kkosh9Son7bK4lNncz0TzGUw6e2Pfr3B//5Nn4L2v/OVpox2YeiHt32su74xWW6V4P0WRruWUrF
SiiTopp6OkvjcP6bC8MuiundHEtXj4J+60oUdq+m2pkH/dwCEaTkfuardQrmJRg3zqXJrHgJPYy9
CK8kajJf1mp2ACGxQtoYIkd5Of1mYuq5iEnUdqrDU19j0VdAmFOfS8JtL3/4vpYRS+psck44aDP9
4h7QQAlmhmkDkXqCcD2NfcNzee5ZKAnKcNFnp0XhY81Akydgc172niJmKoJ1T5lQn/Az3z0MbyBI
Jh0Qqyc2OVx//BxC8byWY9LX2/HaLrgP9IV2QxK/Kr2Uc4TsG6TV2OunvB9eRmWRDF88NZn+ycXS
KGJgYhWIqRtAovhZhlM/1vWAJLoK4jlVmrYjymV5UjbguhgsF0lINOglv+QJ+cYzyubaehw+CJG/
/2Qj6RBMVBLaetLhgFKTwZblHR3WBptITtvmaWx24aMY26066QJM/V/uXE9ZhqC0t9cB20MofAw1
9K1wV7kJ8Bvzx1trvgzJS5U+gcRzDhkys6Lyh4uGW54JWJDigu8wLkO1PlIKk+sjutFlMx43XDrC
cw8kzmdUGXVG5ppQCswOd7oItmi91T/tOyg6mL/NwluMGaDU6nq7DR+5eZhACOrZx4itB9tDBzj0
ElIR1AutFCI8Z3LwfBbVSxPCEI0FxHsBMMNZ3AFDsPMVFtNZu9nTLahFRO3fQDaA1Qm0o8LgRuZP
8cRYCbDDmaZzXPPZd/5N1gO1NH++n9u7LiMhjMbp8ejUmZJixMDazK8FwDSUdXmd4yoGEXCvUp6T
g6KxCrgi7cbZqq0myc+DE3ZFItJtSP1SEKK8RSn+rgO/rg4pxpoDjFMQtkw1WQdisVI3i+FAP3Ab
QbZTswTqUVNG8UO8kWN1VD+SzNsNm6vc973WAkw2Q2aVeYoBJyuAP70IVKPkLc02ZdulCwjG/uB5
AlfKGbMvcasSQsPejg+jt/q9WyHnD4OcAWqhs4hs22YkoufuqVhse4z1IpNb8hfi/mf69YS/FyT4
QWTKgeb0Pfpz2+hdfNELBiNuaIOa/E2TB+WLKWZguzpe8ALLzuh0+qMqP8wbsA+XFKaYSk2A9Vn/
/Z8egJH0vOTdhzS0TrNedadfue1PMNhq+ZF0rP7GBGSpqA59w25xMif1Mr3nE+PskcP7yfOQok9m
rOJsB3vQ5JYsRbYQ1l1kdKX32cpIjyOU+OePwsV/MEH8jHCurq5otYrA2fRrs1tEQ7u35Eb5mgAi
AfOm7QDwlcXaTMzlniavcl6T+nULjOqVSo4iSqH/XTCrpKAT6W7sLMhmbTeWEkER7xu1eFVwvTaY
mblUU02Oe2uM0dERQpldtqtOMntZuKKEbuNQw6Syfw76bdnozjDFUsIdEp1DGfBGbYJmvfMvdKI6
q4nX0cverW8CK1tFnfno/ZCJdZ/qonnAq1a7NjEklDHptDpYHSYNrLlo/JWf7pEuED0LgRKc6lvn
Jfljv+Qf6EVKvNk0HRFqvMMLUBNWfb/SD2g3vZNo1QiXfFfPjwz0VS/Ayfxgq/c8rer1hz/t6yrC
qFDneMzbTQzy7TB0ZqwmeRc9UObbsCQD1+vYElxWyga1kd9szPWTpY4n2wDrJwSgj0qGvazwxePf
MBovObXHscB+JFXA4p17BM1PKTxswtb+rKxtVo+kY7iRV+zuQ8igPUI8cgUMzgS3p/lewJZHCQFK
IxmhFyioWX6ZBFOWVTRRPzNU1oej7/ztKIsjGV7QFZfPLoUS/4wt0vBAbnQYhB9h6A06ohEAmNCS
pH4coqTDz1vbazVMKPCfLyC8pBrf6ZCghPNvb4kfcF36p3FEF0uj6l53rM8j7SoZcA6VP1P0dFHD
RroqWAVL1AeAoGI5BOjlvn7VgH6Eonj0EVjQcDRgqdZyFsnh67xoKEbElBYs7jc/pPfVxFnZcAk8
i8cx96Vi/g0cIu/peL7KUqOLa89ZmZucNdU9pSKyIR0UJR++2qwnIrbIhVPKh9ACkSomgCJms1VW
ov+z7ksrT1jmK688pDvNXvme9Py/fQu27ZDYHmPTdoJqdetg2YIFfYjaB63muM0uhhoT+KQXxjOH
/iOym3RB4AikPZpUz2I63VZihJViUMn7zHMQQsw50jnQ16VvSnxkKm9I3cLPp1xJeHvceR9nytUb
DZZvG2yFBpk3sJAi5Jb74QuCpXFqTHKInYq9B8FUAyQbtPLkSqg85HXEjFKFwIzBKLyHEQDU9eFq
BEENqBdUTEw77bGDMJ3reOPpOK5ewVlX3EGBV4ghoQVWEf5IPqU/b582atldGqLO+5qIwBg7433E
Rv18YHqr2tU9NiaF0UJoGm4Uyy0wQ+SVcBzk5rW6l6+0dxNKUw3qL10vLmx697wOCUJdZ+PY3C46
49Rx9RXTGKODsnEu0Crjfz1xRxCEl8FDD43uaT6GMo62ZO23EALcBmC0iG0tr1jewqbUx1PNpjsC
MWpxWAvdTiyJ0Q1kEazaN62k7GtZg3Q5LY3QGscFQ1H2YCUfCk1NrzTdsfU3yO8AaOFCKg77QSTQ
XBBV+7jBDNl1rx49mXOxhDFi7/hLHfnhkrNNR7YJWzawgyGkvZun5cSKiiCTQoHzeVculo9s//Oq
Rf4enAf516XQBX1GOgop6x+1+7qAkbyfSfX+Ys2EtD7UCzZ1py8AALYEqml9BRN2VDo+OdQ2w/0Z
/LN8KH0OmLjNAZXACV/C68Z/dRWpODTFf0apfc2b5DiGjNCW7OyF4gb4xcqhUNB/g1v2NUTWjYfB
hdL/KpXPXDJSU3tydjgWOTJSd7B9LqtdVkSmgp1ykgCtsiPs8Q/oUQPj7mpLegXG2MQeNm+QsN95
w7K102D6FisCszlcqNQCuaf33gFgiQjj19jaPSGc2yf1C1TkGP03Iqfut6uhhTC3uhD4xLJ+2/UD
w8uzEavZothvNkHE/uyhR7Gd6OKkRHwmunzDfauRREVI6VDCRmhFbHJDGE11/FGzTM5M+wNcCb6w
KiQcNJORHn/crbuBjLeo27LH4DH3ElM7gC7En6d8c7f4sxqsAkL7CHieeba/M86kCTSx8Z4eyU+/
ZouYA9xGXI1aLZPVYiUwFQQsOMvMHTL4gQSSpG9Y/gfQ1Sf2GCcT+1nMwQQ/TajqQlHK9fIuBQir
cSUx4coW/WiuqvMX6NkRgEzHwf7LkVpwvlkbb4BqQAQ0fZWrFKXLO9dE8fePCzjmAVONfPsXGJtJ
FKiQ+wybVv9im9afLV0kfbgprl8oLDkxv42UooijYjC40Yndrugw8knncdBA5AOgzQusSyMatopN
fgbeZZAh5kvpWwvo8TGhS+lrsveMle+O5A6ljojdbCl2A3A/eBoik7xboc5npmUX32w36LUEWdP8
NHAkiHau5QJts/3Ftyqgh537jNUDpDipTWUhr/pONOpTeEOOIxy8ZtkX/gFmCfqnJUPgPeoPndfI
qIVsdRIjZZcJQgz/u4kRISdhN+3mTtDxzy0Iy+Yu734CqIxBf2Ee0aQ5eYgrCBVLcBogvZL5Lxmx
KsH7qJb3dhfpZWw25YNpnHEmf43UOa83p+dN3JaHv5FN/wZp94HjBfNkl8mTB2kCAwh+VQpNbCZt
vJGMjdOkf8uZxEEZDdht65Bh2PjKy0i8cJVTH00D3lc39M6hKWrPSGWviFK4mg4MIfko1bfUhPFm
yqtwPbJP2ixG4BNF/6VUlkwS0wgpycI3k9llIewXXaJpt2oG6UUsPLe/0OUWBJJ88XWBXR9+GMZE
1E/WsiEnbfpp3ppRpiDQhVpENn5v1p2rwV594yzwOjX4tYv6hO0IeCtU0MKJ3XgR26+7wWWAymoN
hKbm8Tu3nOiwTF7F7ySDzWOBDSl+Hor6oG9AQmQG306MaJAJwK0pcQLzzug/0lEouQEPOh9gLC4z
+RDRUA569/MTVpOfJ6rf4587AgAaCBwRw9PRELIMXqZkrdEKbLgH4x86ZO4zekxMZ2QDXwZDzg4L
ylL9QBNH8RN3Zb4ghR0MIjSkMCybswM9no03O1XhPC9d6racDjd/SCT7dz0av38gNX0nZE9gjOn8
C6/40BEBA0ItAdaBDSGAblZqnUcAp9Y8TB2FqDDm73H8OnSbHF6K3jmavWW48GGPcsU78L3OcSb6
Rq0LWMD6L+KD8wTEWLALFXFn9STHckww//7q9OfGgGh6kG1/myhE/9YjnsSPUd+vZ6nNDjYphKc6
smrTy4ymlizWde2z0D+whNGNQ79Q1MYzNniukUpOio8dP1AGyiDWrq6EFO+aQJIDGwWH8AsrqZp3
ItIwGW+K4YzAlk/ddHURkHIPvpjbavYcO83RNbjrbfAsdE+GW6uCooLvEfpUf95HaYKLnI/YBTz5
Fbt51PCGpLgGYcEMEa3GuQmV20p2sKsKI2/MkWOfV1HjoBDNk0TN228jbqIknJeK0WGqdMYMRdHf
ovS9Ex0DnK07ZZYZ4yYLkT10F19EvsVYEcqZ5GlzcQiuvijKk5S/MgrhEYM3u8B4kQDJ3WWQY5qv
XjrPJyRsonbAvzmVwI9NtqAwBH7TbNKgG790xXISOSjNYKgsFuWqi3XCIZ3gneh8XC0kVV/tKUK2
r52HtWBY5mlJPFiSK84T30eiMrPXlP9QRD50x+OUS0coadn0Qp9Ct236jEnG0DJOMqL+PWcDfV+i
XtfL6sq0UYvUjTJEKdwsYTfpgxkjVvtGpWHnLS0uLJ8MOVtxnsBYztgdF5K7aboiV9INY2HBwiWR
mVAq9L0XAxvZC3Ntf4f9l8VhE8htqvda4cOD8G2sl0KkL37knVvAwOkI1yoQAhKCg76JBYoZ+K/j
e+1XjFUtFZMyS9Z4BrOdL6sUr9R5kFKWeqbTOJWgTROIW0XsPOTatTFJn4ABO/5G0k3fu16IKY5F
y+mRN6w1QltOFgGmpvVKkSkbak0yNdxTkpw/McuW941CafPOMbOOe3WqwmoMt35g322F5YczH/kr
8PqZXCZCM6a0/ZuGxLhYOnsBxEqCSUsbKClSz9SEs/gHsl0Q0ZJ334PeiI9bYP6wYb9SHgXWINK4
Pn5QJu/65M7qpaCsXwmSg9ECsbhTNy9vz83Y/ltwSf8L6VORNRefGoiKYaI706P1AFS/RCos91H3
awqA3tx5MiCAfhfy/O7mgvax9cuOXj0FagtG8xlND1tIfXdE0G1JufKBijfdQiVUrGsbbKNMpaO3
uLX/UZPMf1JRZUn3ZukII2JmEwp+dbI34glfKAqysPtaj7F9T6nqYdm+cQSeCRN4ZZI5voUid6DO
vA8Pt/vLZmuW07ZcIhf30d9OzSZW/8XjKNxCfA1r5G53LIi8iM6BHGKtt4qhXjWaXwwW2LaP9nTe
vxxmejQju336a48D0wq2adW2Fwd85SDrL+LbCSve1J62K1Glbxq9I4YwMMX/YxL0LpCEWWJWrfHr
BU94SjC9WDS51ZvEaDSUajJua+7wIPg4oRYXsORayusNt8pBmE3r9UvjH5uZauICUviV9YwU1pMw
IbwCMGmHJfL5gefSN+oksXH6D7mnI0ITlO52qs1NEtP/yPeJfuOwu7aXapRccXso/1Ib0//45RrO
P1Nuc1lejx2hf5wRL1nDYPV8p8b4+SH9GquAZBWRt/+KQQ+iXSkM65GjmNN1XVmw0IziPgyEuXMY
HsEU3wtJ1L3XVabKIRy2sDOJy2c0IRKvRfQkStEIhVwEXOCWyBA/i7JX4oMPywZorrLVZ7d6685Q
10vawnlX9E7UKY1VMIiYjeoWOAL0BD2qTnNMYi9xE7asisymlBdVQTllifGtPRe97aNqtrreTXRa
JxCjEXFgx37qQJ3glezLzYKQXSviL7MPowiwYpD8BK/pUzu7iSyU45vUCUgiH2pAtIqfZSRuWvsg
9aN/RJcukP1TgJwmPlwaAQvf9luxxKRX/Jgzes6eCimb+SRj5VGdfp4eQSJWFGForWaYBVFpJ58a
0nfrDjFXS8gcq1SSXI4o3efmN+qe5VFJFi8lZouqXAU89t1nGOaERk66/C6P7QPdWWoypvK4tpo3
ED9D+xMQsOSJeER/QOIHZfcEEZ6B7XOAR0M6YSYrhXtAn5hJy8vVTaxT30RGcL854Jji7LjF23S1
eE0rRqjgMmQ7Y1LF7xBzDhS/o7wN6Yb3VAVZz36GSg53WGluTLCiBQ1u8oz+9+ypDMlUcMeiuxNo
1p7ghlJwjdz0kbmDfUCjfhYBLBjcFSCwYckU763wkx76l5B7j+h5rcYeZWCwPCFDU3smXnvAUJIc
MxF4itumviehNAnDYkdbB8h5s9jNQNQQNcXDrTs9iSOKrn6YqOHmdA3cdfS5uDmKGseus9psaqXA
jZXc3G3AxTEqIgrlOqROKqS9iQ8vsl4gPURM3rFPPW2clYkr32EyM3jdXxwYsS80dlzsFH0AO5XD
GhcuIEjypqUBiEA4RhcXJkgjn78+e7AyopHdcc/Xm+qXMz/HS+k3TcwqE2LXts1mKfHKfr+Yx4vh
WLRly8q2KamQi4LDRpLL4BvVchxmbq7ECI4T32csHHPvQ0gIoemBDX8fQ7UR6yQ8iLVIlfz8kjv9
oHA/5iA179zZhJRKeGmHtkV66algAPYgk+KZUetWoI0dwJHNunw9sYJGTIaUcawIitBbsSIk9uGH
KNYo1GFSGwLcRl9lhtxLvUszOJO6c6bRlskJS/q0PRc4ZdbE2vhei8G59HuXsrcnh32Ah6tuotyH
j5Ffj5mtRWGIKjsIhfhMQwQ3zZJyXaEjHSHGiTyGgN3xqjjyZ9UjaEAIyWn/tcviRpjUnKnzBzfV
hUK0cY80XtSIrdlqgrkE2+HMPLVOIq+1LdrpZ77XeK4t7B3X70ZnbYf23PPCaWmJWwXGmuy3LmNy
C+pBfEH87ycd/NjYrGlSqXLCSPC5IeI+X7XuiYRYW6fVmBja09VIHdqSeOyLDmiup4c+0+9LYHyo
XDAkj+xlzW0pQop5WPrR2NDEdH7Z6+dC9J5X9ustNgATkjn0wEfSvFFTiQI1DtOITJPsY363xgku
qb5QTEW2iT1kIYgVolkeFDe+zYRMBRNEECz0GTgUlWZO9sPgZFE0kiCAcKwXvrZajmSkvGkBWORr
1BK9jjfKgDhzeZuX7eSZ6huyOp/V7vYbb9badXwZgH2YIOf65m4R1GnUhSXX8gT68JLna5J82DTf
UKDiu0B2U15CyPboEfqsKfr8Z/GNy6N/78BbQIdZ9XLcYfDzo6FxKP7t/ah8iVm1gb9msvlVRaIC
mNOesH+wkYdY39Rjg8kMc7fsC9kwIecj+mZkKewtDElS4dnZff5UjJD/KsuOrmKfIMpVYQAvbwsN
Y+eWHFui1xDvmASJSVx25574Mt1Y29l2coeP4kmO/dKJzrMg6w/Z2qULye7TIKCGw2EyuQW5SdcW
fP8MYyy59lonel4dD8vKsEETrIbmffDjnRrWdzO1bTTY+I/Xw64m7yu0SxVwSa3OL6F+vQmMplm/
PribAOD1FlW0CMVm5+XMnA0T3INSEtr2eeVWI0lM0YfFW/Elc8zSurw2dm3ODGclK4fj8aJxISs+
I2sMuRYqtKuG1DXZRoPu9WJNxzTeKXKqekNvSKmA7gMxtYK7DcY3UuMfsL52QYw6E5RJwJ6PMQ4F
mhrueeEJq6w5MASaavsHYV325A8aCd+Qk955ZsKNCUN6vnsCbd+G5pdoApgqZiXWHnZq0b5NyZmw
mH/16VWy9398mVZz6F/kGNzqCELYC6k+Csvm9sUHD9YVtRGuyMb82TedEg3Ee4eTfJyEKuBC66NX
vkTd5iutTuSIMC1vcyUG03pceDs7Pw0On3JEc85TP9+kdmiICScd6scNwzaaDiIYeQhigYEROVs2
9dehgu0CFeLCGdKJtez+89xO1xfjhpnzH5BzVudEgS7zEAea4JnvvlJ7avI8PG7iySfTwLx6Qwsb
3z3NCyKROENITWTKpekFpuiuRYUc5M/WajtiTKUWh1qDrkXD41HL87IOgrQNaHVLzFJSWNeBHpDa
czThNSd1NNkd2E2rI2TJETM+fa/TP72MdibYg5m/s1uSlwLfivaj/XMD9D4I7f9bLGWvOCEuSHZo
uFS3tld+lKkzMqicA9V85NhxKGOCWt851XsgRNuhKxLE8G+QAt4Rw758a0cIuxYvCIN+6BMQnxDm
gfo8JHp5dJmppDAe9oP+A1Tk+0oTmvohdkg4p2Ze6qCN6ccCAWLc3z2gi8D3motraFGNTdV4rPVO
daawupPgu/VF+/ymaS4l9F9o0dWfDLfHo/Mqt5D6js+LygQ/S0s6ySYsQQyF/61lR3kpLuSFn0Fx
Zyn0SyHXY/kNC9mbRbvM7E5UwenW1cVoNnxkMpFn9b5glbGso/20gY7aXKb0J88EtJU7oNvvqrwi
s2CKZMHWgv3ww3fBtZuJaj2hyZCchEsiEjUjOXMB9OLII6bcHvUrYWLEDdCRaM+T4O77LuLBHf0w
gYCY456BX3caSuDK7mxFd/hg9CYzpHRZglP9dNh8zjRI2rg96ZzDCg0AaIAah8iF8qRDsLBoIiLN
MoqxWBj4dFOllIG4lR7JLZNtZWjia9O2bF2mRwyfZlGGirALOveSU96sfqWH0q3t5xlsx3aapYjx
it3J5asgV9nNFkXlnYXd+1y/aCGteA1jH3SyzZVV2kAkyN6+8HKvl4kxW04u4+8VcZkGpRBlmgYk
UNa5TorW98dN0XGWcTFfxUfmw/8xlkvtOv1LexHOA6apL6lli1ThVU5RxGFi8Odi25i1HbnC69Ac
8XuZchibpzOtBjbZob81GowBuze9NlASTPu+DrDy2z84F20KzwIv+BvwPGCVT8zJaDfInUWqgGAS
SD8so+MWU4dL3+wd+/xCY3f+PfJ3t0pSEEU1h4ssTJ17+8OvsaaljuGPW+NWfpbKLNtvRNZnfIny
Q0T+b0g0I6iU7+21tgZys/6hT9j99DYzW1bP7GWfAgR648fr8PkiloMM7nRhfenlUsWLYywDJ6+Q
89Mh1pHMaRD7Ym9ReCalswp3nQNkSqvKPAH3ydGHXNI6n+ZDyJJWyVLF2/tMOIbLWeFHcI+bVGh5
R+IrwHkYPD1hRbXpu0T7oU+moKsTgSrO5M90XQhncGzodN+Rs4DwNgOEZtZ9PoGyyWSQNvME12DL
37daY/6cjxSxE8oGjJKmoxnzS8P8wvLi20seDoooYnRm2epYaHit7Q+O8+MGvGdEJcWAhfx06KM8
13MHzjtnNpaySCmhAVO0AMaqexksnQfICb7gcRlzDloOhDRsJWQsuHFM7shkhpAc4C5N4Q+WS7hV
JYrlnDfFnqU07lNzd80H3ea6kgQt+TwrxAADnDIWL2uwoycUcEX1KFa2uAncay4JllMgixHYi7cY
GNByGUYqiXqeZfRNwrvHULUw+FgQxhQjxXiQ4bm4SWdnB7nyontsQpElF8rQTcyDP2WKjGsIK6gN
dEj7e7XWF09gJTGsxjukmmasQkH65XHKgR36GfzY1zTfvrTaV/dmGlbqGMJgGg2DxOi/fEI72SwA
Jxn0LJff8iveFM4pz+3+Qyq/lVHwKMwpZul5+dUfpkB1lVLnZc7Gl3ygMfGwDvv/VdGRLZjXRthr
NkqtjADFELZ92tM49K4qRLukd7GqN+4CMjvN/e497DPd8xC+GokV6G/VWhw0zNQFTvEgrpDB58Bt
Qxid6aQ3voi0oA/QLm8zHTUsChFwc6Tvv6BPPLbH8GUOY4k0c40Q1EedXlvkhS88S4zPQlxqB3fi
3Lk/KMkuvCgAsNoVRWNcI0oMGRh/H/C2ZdACL8H9edbqEkZNCkpbC2JODarn8se8GRjnIIkGmbtt
R99HYX29z/5VNpxjx/ewnhT/ZTNivvPWvGAMZrLaJKqBFbIN3nJ2tWRMizryOconEVUaLhNrsacr
YU0SRhmnWJqlDSF9NOziBRdpStuCenaNTQHs72L6v9CqSj6JIX+t8q8D+0oLVC+/iv3YI2mjPQDu
6pqEDUItxWmOzqV3+yb8R+EbW1HUK2ZWiSmuTdz+IVJqo/P7gbMlvbtHaJNtu5QrmFX4Er7OhYr3
4DRj6ewgYGJSY7LHvjLSP+5Y+iYC9w0vtX1dlNjzWq1ycdbmsQMUOzkAHIMOB12YA94LYry+atNt
bmUY81FAkrDuDFBDLhfdhnl/yhxqG5I1NCerxtM445w+HVkxjq7AOZXuqSB/z8U0R7PcKFDEgm9b
c0cuqsT8TSrwdkBjnE4xfQUERrfZxIlvlHvQJMpCzkMm/qKVnHqzxk0shtpaCG1xOhjN6eVbOMC5
fG2zI6XnmuG9PV3tpdlfhT6V1MOWk23CKjzQN4u4OePo1ASq394H8Z6YZxDW2E9qZPjEUgYr3weZ
CLzidBz9Ox+bUYAd4oorWpk8W/JwjxB7EILD6jmkE4pkNhSrsDh/7602J9SQCzlzroG71qloew79
M7nKq3TyUFhkfPGMzbpe9qQ+os51tYVs7eA0IrIRe1wfyk38p8C77fqXSSOX0Ma77YglEz6jXT0I
AE4u+HEz1sEjA47aTF0PgeOZFTKXesBUvXQJ0fK7Zn5Oh1EUl9u1wg3usvTNSovvkHrRZLnNWWLu
c4zA7Yu0AWSDldG/C5grAOQP/k1VzLoq/crl5A8oHPfEr37h2QWRpfkuGiiK03DMPweHvwlo6jda
fZTDhxt0dH22RyvdM4/0g4UU7T9KRX5JuEPcjAtEymV9PnNmoi2b2WBS2D/jx5SKr15BEoQhYuMZ
tXYPI+lSSy/AoOwIbHPS9J/k9x6afYQHP9kU7rLAaDa1rryDt4BG2+s7igvzy3Kxp1zXNpU3pY+V
rxuC5s/Pdo03th7wx1YXDxfU5ExyZcEZ7JoMtFIVTqmPRHkWDY/80MjOr/HZGYjVGjuniciRDb0n
iPs9XKLeMlg8seR+Vx+OeqC+hPnADr7X4Jkr9YLj7IGB99jfAF/vodnEePmxEvmwzDYNeA1QfE4q
oZgcHeOPh5+5M5UCqvr7knk0CjE9AmoC0SKb17MQEy/fqOVd7uu4tbtgtKafgw/1m9b0yvJuLMm7
3xsBAQ4AuQ/kgajDwjvDFeTWh1JmnG/THtpbQZVCbu3DhlkPJ8VWIark+5Xe8CD9wpPXFpNQlbiO
e4zBihQfQG6s1yXDpVmdnXcwqs71pVCDW2uYNcleleW/a8HW9Mj+sqeS2PnFsMWfGxC4aKX21cFC
+dRPe5o2mz9Vsddgi8IlzTe94236/oUV6XtoY2QNg/11pIoyMu1gT53E0UKg5z4dwGRy2V/ozxTX
s/KCJKPVqfs8CCJl/EA4e8WKSmwxIplUvQzkUbKKhnX+4ER9ytLdPOBgn9LvO4u//w54dq7eerjm
8rUSsgH9ad6argkQ/lMSqjFtndSbwiqbSuLSo8uHzi69KrftK2keib+hHPjYLMMlCUGZ1arYUdNL
HE99DONE0WJJ7nRrNLF7IrEtWdK0Zxaj2lq1YIABOX7fFideEdNPXwdhBFUuiRJPjwuiND0Uo1Hw
su6mlyvkkZvsq/wjZtyXpCVWfbJITDtVPpqnimF/B9Hl3CQI9fuqGvo6RO4sHuaA/132Fg9KpnUw
5m5K+9d0iLdJsF2UysRh1lTtRJggbiWgtRZBsPwkz1Vn1HsekwD5odw5GkUvNk/lhnNDRnMmeQ14
lO1NzNGEaBRTZchVY464CXzC2NdysSF5WzHWwQMEQdUrdVq6r3fychX6WSiUPAXvX7YEiFWM/Wiw
uy5datymRahAQI2dqAWmZgyfR46raf2qPcgVS8+EoWFa+VUYvH5uIjTbGirrQc3C8GF9Hcw5NanR
Ekl8ODWjX7wy/I3ibhYtdWzU/r/cD08mH3m4bYTP1DR81wYjq2dS0S90pdvttL89JvXTXjkn3OQF
i7hENG3wSHdzElfQcY0/GzeShcBE/mh/dCyJATQ0fMDZoQV3EZ4X5eDu9UAfJdV3MX9wSFqzLwBt
hwlI2htdxqJ44vkvzRa80W/ApL49orJ1tqHOe13w/47/KS98Tcci1sCK9d6j1t6+inGG4uwn8Aae
cpcCgPwQl7k1NxF5GL8yY+D+6nXv2WuwqWaAX3pcorx6wbHhyuLjBy6us6m+nPmDCIxPu74OGsym
zYqWpLIUBgtna2LFF5o4tZGGXH1/F+kdJSeW9iTsxzOWpjAsdGhj7+koSuKJWIbjpyyIiStGWwEO
amW4L1T0BYvDa9XGJYbtbWUqQthIRW2JLvoktscFUCgkISFQyKkhGEAxJlu7x8yqVkxD1N6nfrmq
/f8thmtsT2rXBXEl0BRQkP3chNE8vQm+T9SyJexmQhcIWYLoniij2nH1qsJjenzWYeyk7vBgb2rz
ellyps+NjomDASAxMs5gBl+N2SxiTICO5Lxuq36l8lpNd1pHfRVmnkRI27mABQqJetM3KSr4ht/9
rf1D/52QSQul61XF7smgfNVsB0xf2HcS8Ch0rLuvXT/3KAGLII2HRaeDp0niBCqZyny2ue3QoUpB
SHITul5AlrcB8UwDHFKNf5IjCDVYpPUtit1tCC76oX8iWc/t5JeSMOU8xi4RGrRqEhZgWipRV2ba
zLQ0HMG7ez36GtpOL3qtASmJdTtRiEQtyc8fsE6QnCQjj6zEvBSWTmAnqnZ+TfHj5hCWTqrtPYLa
Ebbvn6RS6O2GyGUN5mDTksG6TWumhGRoPMMgFGHw8Yi+SpqwRRf3aKxp/Q0UC5cO8+vuZ0tk9TDr
JGpXlgzHUx+k3BLq3va+I+3pKZ2Ddbax/1wEkczH4r0Y7FcVwS8EP5ikLGMF/WibcEg3qzaiCXbl
DbgpMqWqbSk9YKPCfQlreNjRZjQgMGeCneho9ebnXbY4Q0ioUku5HL7/AnFtnp3nyEXpkIMOVIDa
jvBRtp21FGYnOSR6gFgyUUU62OADTMH/LUot5LGZ3qlWOSy/VjNLjdrXkRxi6Zx0nSutt4PL2VJK
657GPdWbbJixCIjb0iV4VZGKVH3v1LGz9HFSfKpbVB4ldMik8ijfcbaZh0sX0eihRIgriTpaacCM
TbbBxBbotN5qsQV0GjIdQ4nABWbp1Of1AR7rAb64CHU/Z8/1Upcz6iksizSIPKzSWOA6pcMfcTM3
hv9XDYDh73NsRsIGEpZ48g4hTLDiPPljXhNeBvQHbC9Y/4YpW4TkuTKhS4ToyjnV5aQBaIgNov1h
nhsse4uWDzva4/YTm+giKsJFBzylKh54SRWTs2Fqp4rFbdJz83XFyI2M5g3lzM+OgCOPOElC++vo
m74O8O9vq6vcsvEZhAGIbWSQXTwRTOiOxztbPTcEhNDmAzclFUDp33GGin+h1LAY/n9G8f+O57SE
JicKc6WKSW6ftNe9OTMbYb+XPXeHRiHLpLDDPXFprgTzTZXcQbdaDT3N0hAtXK7xpn2MTvBUO4Tj
s35jGoNSP4SIl6xVZALeM1qfS2hzfyMkvquGTXSbW8gEC9XXh5inJEKOPT1K7uvUOxS4fSDfgsFu
WF7VqMaCN8FzdeSQ1GdGzqlfYgclcXUM0VJak1suPpgoHq+mWwijFTZsV8y6bLovR7+/7ACMwrQ1
MprI1Gw44baZWWRt64mA/LxCX/reDSpBsS5CRKSadDsNxLCC2OX/eB+6KsRiB9g726E1AB2lNf2w
bZmSCbWTHsWqegdTUrv48QRv1wfzSJt7t62KJ3onkK7X5ElZDeyiUexEFf/91bR1iTtosUSgat2h
tdKUIKskQzC5H/8V/YeJgwr8kMCnc2wjQ8ptx0i5YAbl/OKYQKjEmrCPhlxrK4ju4q3+oxIMaQWW
G5wMGYq9VGNmUzi1mApYfragOg1kXb5XTUNzkIFt8qxJE+jHPdzA9FmYYcni9jrc1cXkrxvGYnJs
JaJHhqhYPp98ldty/NGbR7tPVPHXngQtIDNPPIrHgN3SC6pGKhitw0/niibWP7bw4UyLo2rUPvvR
lfB4M29gUdYEMV5x6Nx0g7ybhvM394YQuYqeZSIYAaPGQWjZzJTIeIS+EuS+NBoUihsQb3OLsEBg
UJHuqQkYg2J/4UM7l0UN1HkpG7aV7M/m8exxxo+44h044FlZXL5AiHGYDd3vSShiujHMpMRCyl+i
gu5He9PP+5h76MZIdGoj6xFMqsnXT98Rrh9LuEt1NPK6Vg9PWNe+fwRfoqgDwsTJBP/1+skrFu5v
Piz1wN6D5sHEvQ1SeMNxLD8ri0UhXFHuY7ChJyds9UC9/TLRpnHXgq+HIgnTWyk0Ynz66VU7ds5m
OdSsE1YvWajbhJlw/gQFWvHPqbrxaVsLK+wWX8CyoSsOQ4QHB4kTM+HqcJYCvgXujTkpnpDXjfq+
xdIxZ2+hP0hqCLFPqS87jo+Rv1mkcPP2uDN3twlviqhwnDyejEXKGiTAznDeyFeLqbYFV12GWSS2
fjxNXuOlLfbCpqhwmHw5OASyjxRQqFW3iz5m5LrjJCnqtvLEComvjM30Xa/gCOkotVRLuTLfvEZq
qSYjGBQ3iUHY0/pRg3Wrc/X3LNdpxwh9kkBC3GPc/H+wwZTRhy09h88J+HZH8q2Eh8iS9cAfqH7v
FQoSL8I5WqnqPPZZCNzzTkoJJRD1YMzWXSdPy2t/76rfcw0h9G3I6xE4GBovDsrE/Tm9NE+06dgB
w4PwofAt6nmK9HhDVAekl7Xzw0pweXxP0vbTfGEhtlLshifmTh8GYnYbITryUfk2SltS7mamFRKC
v6P0imGoo3jMMBKzCOFhnVw2Kw5G0YdAMwVfRLqFiOm1fSTopXHwnxVU2Iuo4FxfN+IaPQUf+cqO
KkzvWhtEVB7dPmKmMMmMPc2b3qN4YR3dxHO8dzurDmuJE4zp7jcvYjfwNcuG/WvaiwZveYbcWIS5
EkA1rI48yvU+zJ+S5lT67ozbmQ5pcLeEMDE/+PzSnwHHpPVC9nTE3DnvehADpOMcDLNz3KIlO60b
Xiojos9YEwFEz37pIz321aU1w5XOznpclAc+o0OelK5ofBysAgqbb9eKAn0LqN6onBz3xB3L9LvG
mkN5F8zpc4Gcx4/F3FWVafPfvsmLCpugJgl/KQs4XEDNeu61kc13V0P7txJnJlboIaJZaqJyrATz
l3337CDMcj0lQf/SqjA3iOJzk3xuurCpEdg86VvjgqIcN7jXiO7G+3RwERMDXHzigW3Ggqy9GEnd
cGktozV0I5nknO5R8hno7xiKeLBFXph/C0Q3+/rK4jf9/Q8iaKax85FY4NEj+rbyYQdThqp5Cnb3
dt+Dg6bMtDLfSUUmMovCpXRxQ9J4RFWdLa9qiFcCG6+1GeJaoTWBAaZl7ImwI5+cMlSB6EG2HqFk
YH4MLbxiiZd4Fe/zOYNG6A9d9igdijBgKfuW66TrWcd+92rF6n27sdPpoeE7HuAiZpUQzHnVw+nC
9NPwU/702v3jb3PU0evTXSky2teCiF1ywEcPvqZOu4s9jptPqd1gNLtmWa2LfrEOT8TpFZMc/xNf
jGoZrd4SU2hz5aXd75Rp4oWUMwnx9nlGvZmnzYv4liWRcOQcIA9hu6+d7YAAnP12qY8NgFdL0d67
DTGBQEWYXZPmiUXw8IZ8uDpPEWszyOGDt2BvCsl6q6APd1mdtKdnD9bWcJpiwqR/t4442KyTEsyu
laB7ut6jV2yBQ3EJDoEY60pxpTLQiBVXGlK3gdU49YwVcRsXD4tGzWVZ3l1wLm7t1EvKTA5Rg6VF
Ee0884jxLAUONOZ5WDr9ow4ihIIDOCxatEuub37uoXWgKFQykGNcZxuyipfgnNdozCveY3fMaF+4
jLgmYueiBbvFPANCeSP+WpoGNc2c7z4hdI5AKoPM2VndZxS87oQ8/63+8Dl8T2CXijegrWF10tK8
cm1X/7E6Cpq4IJR90E7TATh2MyHMexqihks0+6San0zb+QS5IlqvZ60hpRXam24xpgZsp0fqrX0N
UFMJ3hYCIgaXpbThbxYXZUsaEY1/ZZg1qKIRcwM5tv0QLON2pDfVZKzvY4hzkY29Bm2Wu+spe7YH
q1EXRQF5KrkqjyTP1j1qAQR9ObcCK3mcLmXSJFszWh543gVhZ62W4LjWuBlqwcmitYQ0BN1tyvHn
pYLV9uhFmfZ2hw53iD6+QhmTLFtr7hV2gnxTJGVHffDYevSqdZFkxraM9Y7UnEfYCYaEtd6uEDCx
oyW/hc1AEnKEw63/U8WBYcxbGSboLDriiM8bSnvGI3gMTpQSRgzedsmm3tGabPe0gqPULLuhst9S
2n2B2kzBmx/2VMn1eyyzzRjkgKuOQ+lJNomdA73Kjt+HU4PwAdDB/Q0sCTmfmeTUqtoQTK3j+fDS
v8eL+0VW5JapLhJmBI0JFlGWAe/ea606cqVmxrbhwIsiVCvM/ool4uoOrEVUI8udrP1kpyyR+Oou
EpMn8B5OJDW3kkgxkIecQZMKh9an94PAQbTJWLRLE4HYwjnLfmdKovAgq/k3Z3/rkjNb+0moPUVH
EJmE1FhYkX8YVWBTkuaczK30HuJXmnNW7yr+lEfRusEu7etW7K98eBOfw6n9elgQndLOk+WXds93
WMj/CIp9YMsJJ70wWyQnf51ftpmvcwtNGZ4YId5KgMC03/l1Ung0zO0so1Fvctmx3YKfa5p8b0L1
AXqZR4flg4AkcW+tMOJ6WJw3g1EgofMHKd0UAFIzctyuq5VOw3vbttuysn3r+d63l39lrYi6QHC1
XF9DXmPjo4FmeUv2YaM3d00x4mTvRwkiiTqgWl93pJKxEOyC8f9zl2/Yqo4utJeKIcw5UvEKYIMI
BkqHHEqEZt5vhKyAVuwrcU2BmIFMFmJ1uPi/P2nO9ipjYK2wMM0kyue/1i9+ZxheEhs6wUlrYmhy
pFc6dGgRpHY47hRCYgZCP8Tc8q9BsDRQqFXBmTt29m4O4soKHUosEGFM3EuteoPX0/c9BKa0P8hR
fAczCbtlf/ZABl1hIsnS+KLjywyti6GpQE9U21Bik9abNc0drpGsgFtih3LKUcATPVSva/vTPhlZ
A4q2GAA9yl1VVrLS0y2VnEFmpsIhqMclNpzLqxoqacCMCmY/EEz25UrhOZ86k1dqc0qSehHfy8It
clf7N1AIef5I6HVxhcrLuOCcdP/FW8/n2h+w5BMti2lQpH0emj59DyPKQaJW6bxXXhKttgi5yv0M
jVCyrqph+lyg/lhzXs5C4mnv4whuJ39Getw1BWCenNoeO9jHAEun0iBjmTohwpOfDDVNBEVsCA4v
7m9aZKvTiEDMubv7mIG9HPOTh4G8jDjGQWJV8n7mfYfLAL2lXz8SgGU/rDPs+tGuxa6mFCx/tuuz
KRM0KI5DV6jN5mdyLG1oLQuR+GDU7ZFj7XSwjZcs3abHfGSjK9AAzCGSI+/NewvwktHPKCoq+/o3
IW3HH7qgsOZbExj+njD/zsgM5JVes30ERlolvouMPsu0H65aPMEBrF/3WWkM0H2aX14wk7FC9CbX
wMsWkjGsRRa0qB9fyNQ6jrkbcGbwBVwqrWEVNA5ZKuhq7kDUANuoFMxKbbUJy5cKxoMeGfiRduw8
4rUiNwgHixElcEhMTTR4vfMUCqf4agsRWF8uFjDeoLDrWP+B28ExV+MG8IqwaBGVKEaQhuHzzFOu
TKuGmL0imOyACWFpAkALgoqtlrU/yT9xOaRRZZzQ7ekdY5trAl3RSIgDTjWe3j0jVDljT5aQgxYR
vkW3D50Li67xPSnbUIAVR74h0DogkP3XoAbHMZ7Xca7ojgRqAgCUOY/N2MpuPkokhc3cttqLL/hK
liNEctbcZyvfLNc5ynnpHkwKYuCUa+lWGpUS49IVZbtJWRwUbuqo/8n+IWDTIi841P1qfvzxx6Zd
QIb/D03DEH4JM9FJ5FbR1wrZPLU9mQLW2RlpTu8WE/N5w/NoTGRDoxhP+w3+HPnWVhmaqp4Fx+Bo
76bIszAJ4P7xFDRjWQSGcYsQHh0U+YtHNs6IyM42k6Rkz9j08PZ6lk2hHdqZCvX7oVW3KxOV5HCX
7M93PIX4YIJVbfOP8tNwT0evB56U76cslUoRuoNxaSRT3+XTamIv6PF0N+zWJSjyJFgjqgC8PASF
javRjG0vDvl+seifUNyfx0ftCtWux8ENLajGo8EqTPxLXSPCaIuSwfWsaXQlGuRRBjZQ1OvS/Wr0
aS941Pup2Onn0kxST3qRoruPc9LdDWycx2xd5kBdH+BUxvOHw4EiDwfjSg75aWvPDzEj7KsVNc+j
DyOrjPOnlGWtVo93rViMmuwVV0Dh9u7Bd5YhuIC34G4VVCvtHqtOIlt+qLMvJTHVYwOZE09pvHDG
ew1hWAGtJFWpMo3tZoKLAWgk466elKnU/ma3BQh34BHk7+skEv1P0GsEG4D6dQ7SFqj60KZ+4sDD
M21vKt+CPgetZUh5m2eOFXluSLONuMO4yYaKO4vFAg9/2kF1t7a3/RQ2PmyBg2Vo050MT1BGtkAt
K5ZUH3aMs7GuudjvyHZ8Ebas9MIR3UqtvpzEiYm5Y0RusLDcBtpJREfGJtUwNUr0+KTKuoqnycRb
rRsiXJpzsU8aFECMSK6UcLGAiVHfPi5Kil9dIDUyiwHbpiZFlyK0QPjmrkngz39FIkPOQRS95Zp7
nKHMkFlShe4ZrUu5SUdfXf3VyBw/pgIpJe1uHQMRTE+4gSdGMnDqpPFctcWpunYiPQg9THe14fag
gm9e6IowgydXcx6lKtKdkCmESqKRld8IvZ2vbGvrB9B0TMYpbqJoj6F7YPYWqmKT9lXu06bp8QMy
I4BiW3z9Ty86aCD6pWpQnZUTorhZAgybQL7ewpVOc75I6mSnzuPuiuWeRClO9t1TWGIp8Bnq1saK
cAdzqw5Su+wy9S/EOjFzGOsyEMHfRRhD2X0AdbsAGMsi2LucOlYwjfIsS8TDfmJZbB318/TIGtJX
zGqfUuYnNxxWk+VPfNGfiXH9zjZK4MG2G7X12kkUMLRJKFdpD/iT5Obq9Ox5fIwbTVAz1GYex2zB
RkpH8QOiVBqPBHYUfA4zBVeLMH3pCTdm4rZ+i2omiouwStRKBteLvE046vpP52lmNwPZq2MA83dy
LEwpcmrAaks48IMYhwo8mKNEDobtS8zzd7lF6mZJn3MDpdj/TOldJnwhISrbp+UvkCQ0+++laoC8
4MOwzZRkHAtaerZe6iDVbs/L0sjS7KpeSsEeFgvJd9AJDuAagMoLPhE4DriBSkG1RRelI8PlL878
7VcoQFBv1lNgc9XunmJ5jTzz77V2xdzsuHZrz02Ym6YPFrwQZbA5RjAPDtdUU1O2Vi6yEM3xhj+Q
TcKMIwhB0Y5Fbz0jJkmL5ya5eLu4JNB1t3NkqrvlaBJrEEiX1r2AK2RZU0Ic3PybH/FYnRdUuT5o
ZpytV4RcBG+fB96MEiSDJ3cP7TujInAidFX60E0qECjyosj5Wi0zFQDnj58fGY2pHipFrtYvQd4Q
5lydt+gGbRCKgVY5udLUQb1k5QolterzlWWLzYy90FNFazTl5LSCeHWyQnatsrHJqmDn5KA90byF
ZVAvz1NRIspNe1sfaX+YqegXhjM1ND/xDWufX/qT94zGR/M76Iy6w3i8oZjDkRG8xlI7jo4zsOg7
nJBkhbQH2ue/TtOZf3qAPBLtFlTOJmrlrAKaOuqtOYWhmZTr4B+WGuoSdCCZqNoEkcheJxaZf4Kf
+CKJ6PO5WcBQ4TwBT/i1YkTbqwTDpJr6uoIbUWSkSL2Jga5YUIwsIHOeIo6xeE6WdKvwEh3EqCo6
vQjs6i5eSys8eKHqy4XPWujXf/WEgbKZXy5V3PuR5oqCtz9FYN2iw7ZqkFGQiGGmF5VIipjlxoVd
SJNKYYYadPotrc2LwxjyHkipRgngas2cvkINCerQtHqOPyj71e8PEXE0Vq2orVO5YKE8d2+L/Coa
Dz+R/Bmvibakn84xeR5pH+AQxKTk/dU7kpalfLTYssdcWXr8Do5tl85jvhLCHOF4DItwxLb1nZ6Y
lelQ1Bjt6zQq6/ugKrTwZXW6cPkCQAcXPkLOcc52q7dUiK9/Kd5GRO0K8KctqnnzDmkCsox0T/Fq
ObPdiwCodUzVCeqlPxLIVxJvBTTZ+9xiFiJtaRZcTrI7beCGoXdPf4HbxA8G/IjzMCuKH47zQrUH
pByXgJ5BlfxdukHf07S9hxSC8wW5Hm56OKHUs0OLQzZOO9cUL5ouuSxo9sWdrvO6Wo1xacodv3BW
JSW7LnHc5o0Pw5bVSMYxIsIcKFnfIFKkU/0WE2XzpipCnJIwO2TA5ZfLnXdTI/IyAWiT6IhCB/Ro
SjThiaUC4tf7h51klBWUxrP4dFfQ/35Qz0qsHMUIUWH0jeZf4C8yBJmqiu2Lv5kqr8JSCIMozbCL
fuIxqfagqZUikSFGTtnK4IyBU75gPU521ohYG3/+KtZLY563va0kuOus5W/Et5SO5K3C2H+S9sjm
OPd+I5H1hkDIlgmAxlvCs2wvPqjJ2cPNXZO/tdP4ej9GhPxr0zafgsMfNqRvFaPg+afiauXqhtf9
Pi66xbt9Q4zSUMh1X99BudT96iDjdV2SMUqF+d22OhGJxQJfuHszHQIpq1ZqlWaJLxf/h2cThSdR
eAmR8YPF1GcVoia9Jtum7LwgnvVMALb6mTX52uVM/lMCAS3sZ0bHKBg29/t0j8dzNxeo3FxCpC+3
bKK7GAzwIcv1TOS69WnGW861aAq2+i+ftmrrQ5RX23qdt1vVuK+jlR/Hi1edOykNrtd1oxCKeF63
6+IKc1xeAqo3UqwEGzi9FTuhVZe+Q1hVBe8e8tEgx2cIZ74ItvPKYVrCZJgnUB6MzXiygAYgrxUb
dOpfTqmSc8J0ob9slWgeLZVz84uChpr9MLyt0gwPuMZmepLBVkJz1VMf6NyephNE6+8aJwb7HaB/
0n3RiqGMxXIlxoPntI4ro5JYBpXzny9Z4WXBWhBiGkEST6usk2pM06sCJrzpMPz6IjXPSjnH61QK
jVBSz/fbaXR1Izq/T/klAuz0SGnhBRPQeyOWLxmj6qpWupzZH2xZwIHp1MaFHKBfKUIxA5Sixm6x
ZwMjDLM5YA0HYW7L6wDQT6l9J+Ny3MIgkwKy/rxlsFzeY2IM1PvCpB6ED6Gr30uvSVxXgRZCjwC3
dAG6BFlm5ejkb2nY0597beTvEAKxOKZ8R4QwwVPIEDIFyyEyyWmzlh+kHDtJJfKXnwAyOg4wdzyd
deOugUhR8OE6T/9FXiI+O55qZ7XRyF4XWD9XKVkryXrz9QgNhLGg55piYeSDM6rN+w033DiUEO9b
4GBxPf2lnBUsbpoRU4aufbL9uoFyZ5a4atBd6vGNyGZySYrjaS3xt1BRMLhQGmNP+7XvmAy0F+Ca
CuelG4zi+HSpdLFml4BLzVP2/dH1jBBsQwQwjoCt7ul9yIePpyeeVOq/E00Tu1GtfTF1pv1E9Rkb
/Fow34hzXnpXeP4huKlYkA/xrmv5rK7le/SqFCL3r0WL3kUhVewvY3xvtf6SAWPwVAr0+khj3u5S
mZLud7auiUC/uGwryi0I1EHjFu+DEepDlMmY8yHIMD/LzwuwyhHQTM2JDW7wP/iZYEHXZ8s2Ia/z
lRQbWWcP1ze5Cw1cHeGqIYtoYJuQ87n/WDQVpNkXs1QX1zBn4dUp1el+BU+KUWUntM+w6kNVRx0p
JoXMzGZ0MNdEQXk40SiOCwPy9B7Dv3G1s0f2kRjyhpUFXlwSA2jhFfWDQ7HFX5POtU1EfVq2MS2/
YAck9AzKIynf4q5nlv6+98GY35rUkikzasMlCWyf81Ht683/m95ZNHwrH8dlGV67eVTTrij/WGkb
zVaFTed7jOuQgEKoyMi+LIipvTMZ6ZIsJJNiTc3SRRc1GKvCuN3IaNuipz3bJd66A7DVKJ/FEeDB
gUX3VnfLAOYk3BvNpSKmX/Ge326kJ4Ne476sdfBRuWSugqD5YtaoCPrMca9aAjh+zD6xvbT60QXb
BYq7qiT3NIQQmGDE2HM0M4120+IK/sWledjCMPR50HUjn5ECMF6PEf8ej+ScjUyXHQF/KoXrgsh5
4phpLIyvOjI84NRrpcGQyZsy+cckpntgAJaL77/GTumV5+wAXiDctdwaCdRmb2qzHclx66waG9cB
MJavJqcRFWgf7+oKaFhu8NCY99xqx9qD9hOGDqOgHxvblz/38ld5LW7CjQK1e0FrbGvDqZ6OCZQG
hevwHS0XYBs1WqqqgIPPd5vlSSLtnUQkaIoQy06pR44WKLOetiy4d7rnKSmt70+X/G0+Af/4uZUO
5L2aa0t8VUY+7malF8MoOq7qYrLOBJxyocSqEUu0Gn5VaknP67JbMTdUCYBbIEz0GObzWGd54kGW
bKIaTMlK0qiPH83/bPdI9QSt4h0z3W5hthH6lePu2Gud1aRbBNFKakOfbxDCTLW9UE00znUWbR1z
xfa9bAp1+daeOrCZVrKpBf9Hu1493LG12LY2TXFqvsx6ccyI1FTlEGWaqbHCkvmrQwSKcdwxCmG6
LhRAEXzTg6WGSTls7eBteD8LaL/4Bx5xaHbYMRsJiHJFqA/pF4WXJhCD4o4RuVnWI5xzFe00ML1w
lwdMDMUKXglu5b2lVPAGNvuvctMZL/VuWS3S7mlNeb4iA4+k8yjuz2wbffwV3jimeKghHZmYGQa5
yVAHPC5Y6GcHuEjlvZK7dAO36ZwggpALXNLxKD1s7/QPDoaQX4y1tnYxKvINFrVc1ENCTHIQsqHp
mZx60Z6/wLvBbGMYpa0SgVwP2uFOkCrpzrRPoHPxUkiFyFAcy0vMmjpQD8uZV3HF4TQyuc/KkJtQ
wLNxRyj6SwGEMcMoYZLUxaDyZf9A0+GHd511CWebXG7D6LZ2QJymQIZviEspQUlkgW8TbIkWQEb+
6xcEeOmC6t7MrqO1u6izCriSKFpxGj5tKOwu/Nea2I4ZFybGnffxNTamZMeEz+yXduBwbEE456H/
h4+y7sgV/oqzDCbkj4tg23vCv7kzrvoxNaCN3mTax53I4bMWxQoa+kiCgD3eHJg/vX9mZahtkZGQ
FVv6EOXFckupAXV+y28S7QDv8T302JFUW0oq7z1SkX+0LlYKcCR7XpKEcdbkMcMe90rsyvd0YOgo
gFwCGWJz+xbpqSTF7FXGBFA0mJ6fq8IN6mT5RLcxMt8pTsys9aB6Is/lBDARsa7+MSTB9DIS11No
+pWzSQ2Yv3pX9lm5o6NWm3iusmh0SJxQyRMwJtYP2O1jNOi3L07uurtTpMzVqShsRUyxZtThsIi1
eosePnN5ZNMCKqmPH7yrEnUlmBg3Da72FDl0/hzkz2svlfAwJUqIPV9jcfJ4ulbesxQm6j7317Fg
czstdTELR5Y0+AxHulL2Ea3Dul9M50hxhxoZUfq+SlZUbUbt28ZJDuzja9CNM6vt+k0RE0tz16Uh
2HrlarAlrAtD8/WhqhU6K3Kz0cMGijAwpFCGStlGI/QjmG7xusoCZGJpQFnHUckM/Yee+pIsQVax
PlNYt7QbO5dDpDKklpWBB1hUNN9qpn7m6ZOTNmBWjpp6F/Lv15FCXdmPki04XqWvD2bfo1BQZhOM
kOrq+c/DGBHx+ZRlg+JAxegV3UvsR5cAikIefAu1xlMHPjoDBpZ+bKW1W+KB4e4O05mdPd3ahrG4
zaSXpxLaKQKuVOe9cZCxUYw0I07tbt/mIJy9IYU7BVBZp/N/JWt8NmPyJFQgkTmhS4jfMsxeP2i3
TrPGhFBM0YsQRgCfBEXuSuKLMPSYga+JdSlu9ryBt7pl3exGxcPAsdc8lPHapph3R1XPucaxT2mp
rq9jSYOokemTbiXgIx5uebBlYZQ7jma303KVSze2sxktvYytAMAJK3xbBXNzcGYYlisDDjoBQdrd
we1B9a2jgLqD+p85OgLTZRYXe/ZSDDA9+dVOcBcHmmabaJpyMU3UjEgR+pAvJG90h+I62+Jg/x00
6fZxB5Qj44YhwHGCBYCjmU5MBa8P0JZgO0g1uSpMpraS0c7OeX7e7UpuhHq/3XhB+GRNUh+N/Jc9
RrvszLFkDkye+VZ9D/qEtSGImp6loq+RqrfkivuwrWu4j9hJc7vXencJsHZY+d4cra9VKtllyvJh
W0sYDGqXBMSqzlTKXNLv4+XEyIRH9+0mdUPmR0Qru5nZUsEx0I5ygHyWaCJ/boKgDIAW7QcDJcqa
VuRu4GNMohwPFL5Q4QXOwB9wSAj6kfMDQP0VmONEJiK74/kVxcDm+zKPZYm0XjPHN8Dd0rNlTM3G
21mMEp1nYnI+uFLsQvkCm02mkMJd2huxVIUBcIq/VlIwBjJ3WU27AMikGtuuVtKYQQjfBHH0dFRg
R17V8dlI8jdpD5RxaReXWV3ZX84SDmMJKeNx+Katfxbidzq8DCMQBEf3qBAYtx27s03CJNcB3hBW
iqoZP4Brb3ojOJAf1+u92ZyC4Ue/+hN3Ur5CXVA9urKxFk5IthOpB/FbC2MECvvoDpI1A4tQhG7F
r11ZmTC6Exqn0wX9vt0ANXTB3YotCyUKk94sgycT7eJLHh4n42aYUWDyJ6rRlNPhBfft9MULfLOx
p7ND433xlvfKg8d1+dcqAcixbxOVUsxCZSTr9/gtXQuC/iz/hqlbo2VLRrtBCv/u9u3ROjdOAAeW
6BBwHd9alOEsZZr5SN0eXsHmwJEaP2ZRg5S/hbyWmHC9QNfWlEv9D5ZMRKBsvMojPif1vezDZ7bN
AqSM+1VyiW2MXeGHhSZu+8dfP/i1nu8XaXyCc6K9hIkKHFfmh6rNcTER/PgQNK7j4IubkENIEk9i
X4pVlwka8Q0/QMehGyxXCk/IS8QwkO+wplyzcq5ESlVOIIeZoOfEmMAbFjUtSbU0zLh9Tbe9kw0w
jjbuAEn3Gr+xOFWOaLk0gas1ntredIAU+QoNWTKydmLhmN+iI4L4Q1rYcB2gNE1n7kGSfr7GPmTR
w8MtgT0hyyH7bYij1lnuH0NR7M7FTgGcNBCG+PhJag6nj60PAKbPx9ADjHt/WAj27xwzc5JrYMma
nrSUIy0mabEJ/IX2f1syBit2hWZeRe228mWKNIGHzKQ3r0cvwoKuZyad6/3tVDi2ShFmOE5TYsRU
nGe13v9aoVzLcuP9CDepqTaiTXDPVQTD0xC84i/mV+EsK04LwwxWG+QwlPYZhIm5sza497dypwPv
S4CVDJCXo63Py5c2QGHUIZ7BzU9sJNW/f1yWUsRozNaivNqyY7+WuQwDf0NrWxQdjRKbmHXR7Pnr
qrXgRoc3cKJJGfq5iJtEpFF0umuE95xuaOJccO72SVHUTV/xVy5NGZoLTd8FED22ty2zn1eArXPA
DJRpOcVzZZohAItJYBxuhk6qO0XGITnkpBkZjHqZjfg5OsxMMTlXipQqPFk3taXUKvwJnVIykAZo
S3gCBv2xkPfh65fIVb9mJG5XtwCgMp/sK3QN1eoGjf94NMNCwPceiLx+JLxRPL1H//7WpO40KwYs
GF+HMCtvyV2L7onxPIiLlzhGv4VBdNu0AVCdfBrXIMKreZG0LVoZdRTsnvv2vIOxMyoGeIMLT9/R
J5t2LDXDhxBYPDSfxtv3X9+OOJ3cg3mRza+8kSQ3b9MsWO5kVYITc+ro67kwrqhR1Y8wFPLOdoCD
MuU1V03oijdI1tdkUIsQK78tH3N1sMgPheeTqe1gUoVPgvz+4omT/VPTzH+77ezwEUbQl26z1rIj
ZFXp1aye+00aoABbWCByU8fA67xcvFeJ+4uZv77H95IP+nhglyAVWhPB6LI+CFTc7yaFw1EPiWbc
7Wgdl5mViK6fc+5JX2eGubrt7a7YMqWQqLICx/OCp4Nz9HVT49zJ4V9v6zFjbaXOZzXkd1LDti5N
d+NsnkhB9PT3B2/pmTYWRjnDyZsccL1Dhv09AqW+Y5HuzMHUk2dWGbA+LSXZVH8jEPPJi0UTULoW
eUdCfdw2oZtO8EfwKEl6Q/dWD5WQSG6v1egEUyCiGsVLztnrvLbSR1D4J/+QrBJhkb91qV1RKQsX
ZbtZEUR1gPBprj8EfSIG3XtoZrDjOrfUMUQybjt33sArqOnfJlrOJXqAns36f3db1arlxlQwIhsR
OwAoeVEgAwbNLWwRBrhPuNN2v971KFyt3uVnv9BU/Px3jLs8uW0cAZW6gQInqSdZ+LEP4JrCLE8y
PQ9RTAv75cnVqax1wkPyjsJIF3CeO1WYvBMX/e2oazUGCcFTrM5R6gaHL73EbziT9a4eelqBC+SV
tylzijNqdhSA7UGrynvSHyx4h8pOs3f3P5H+L8MDKAsD4/lmpRHjlRoiH9YH/rWD19zAOt+TG452
1QpD/ClJdJAuywP7ZDHgB/KY3FaBnIhFFvvdqpTPKyxpfWZcRrIPfmfcX0xzQaDlgHgaxga0DTd1
9O+ooWGDidngLP+v5UQ1458JTlmunsAV/kGwNa9PiArzpkQ1BWCQGAnooiGljayZbuXo7QcVvTc6
OffSRDm62FK5lBPl8GZ8uf2Hi4pM0z9h8+0UElNfXyLipDKaKJOTqZRIxlkEGfGTiAqH1QRzMOeS
iwqoBgunm7R3WoijzyZhFErb9vy2byMPeh5kZXXpYVrNgqEVMcf3s91im26qVKOoY/b7mYVKsbao
KJdLrZJW6LfRWJMIsVXF1JvqbGDbaOIECFsUW1J7zCy7ownPHXrnI5q/Zq1cmCGy59bVX87Hunob
g0Xq1wCLyFXTEI5i1jLdSFcOKvnRQvYnYQH3Y7P2O0dkq4IqyMvi1KTRUWCQUUnzOCujRZ5gQxCy
UZ17bwxzO801ArXsKkGfa6OG+Z2hLJO4EFFEjLzDFPfWXzcVqwWdGIc7ymTGWkJHcxurLYS0xM3g
iK5vhj5NQKo+xauSQUVWrLgHO7V6gYiBTrl+2Q0tCQwU4/rwAgg+ntPd1WK0bMaIvx1uorrtuea9
LyL51KqZvK9uE23OeWBpimg4rQRH9scNt+yp+6MlUf5cXrx67zKuCasyFf9F2EX3jrxOuInndqjR
W5/++mF46U2hOZgwM4qniTK9DRlPhLALrBgK+ecdr4BWBj8hhW1RP2LvBI1fkoB7t7oH+ub4F8Uq
jD6tHgbcLEdgl9ALKToaw/6GpQ0cV567mESBFPJ6MEf9u2gKyvjIyRMm+lk69voXIQqWw3PTwl3D
ZvuRBU74AbPMQeXnTPoWROuSeVl/A6Kr9YRaoWK0bpMy9NghLlr2oOUzwICSrJ2sflVwsNsoC+0H
C0jJnZPNlWuor+0i0Z2EAkyEY3uxjQgNGbYorRH8hQMUGtHMd77XIurNf2qva0cJHZbGz+OnQJZ7
XgAS7Tz3DycytKj1bj/OCBlf1SlZZPqbqocv52Bjogj7O/kI/RqX0UQ8cd5NrGcjQL3vqK3kFZMb
BuNlJAMtLiKD30vqTHlHT5ZXonQN8IXu9tHO6AFnKyeFI2erkTfOD4fUjcu+jpwCy7sqQsq4iCpQ
lWB96AS/2Sg1mm49x88oa/afZY1vLvb6DD/r9d4UkDKfkwMd+8fa/So/8Dg4jyb8iVyEyL+yHrPk
bmCqtwBWbqWKBAPXT9egLMWbCmgOh+zxF54GHievRLqi+spj8Xk+G3gR3IQgljCc2t//uY0GlPoZ
lUfy7v3oz31hSvgJG5sxMHwgJwF7xNrhKygZow5EWbF1YVg1++vJjFnDfMzdXEueKtpJvhzKF9ei
TfryH3bXEpxehiwCttOA+ya/HI/HcxKgwPgzVsAPDN1Ocv+OOMN/FUKi5BQHZ4wau99w7h02N20N
YzN9KMUWGGakntSlpkYjBu8EKWkj036OGJvuJcc0LySTtOVfg++B6X0sQ0r33CdTjkhnD7DF4iPm
84vHIlNchDgYX0zl7fFDLUf8eaYk6VocDlOAFRgQCGukmdgilDvU07Rx5I16yY7E+/rdtwigGXb3
3dIssuj+nJWpUqnOweeAEMUpsdF73z29RHZQqfrG2jn5z+f8Z7PXJ8uzf/F0YG6e2+o/IHgs6lUh
K7lws/UzUSba9+hfwveoYtEITd+MGOZ3eRmXYkwcbAljirClHUW/Dpf5yGESBwd8D/kLBoMQ5ihy
2t/BMsW7uZcf5M+sNr1TrkO0okANIdk0qk4EQUIsc7bdQcLeUVSZCXa5/6jOck3rFQkOKQn9Ck0T
z1afjRsgh4RJvBRVUyVymUWq09d+2TbM3MPWB1oVaDLh+s+lY1LSl8Eg0+6RbPg/X9nQKlrWbMxJ
SFrE+DAEbnE6fXXLYyCegp8B1DShNfZiAgaMeavJ0YDm+EEJawlgD3wRsm051aRNohzgGijq2nc6
tC+h3r6G2P2aPo8cg8K+1YImtMcWiYLD4EmE4T6rK8CiZJ0oE39VBkwirnGOXJJQSPOEFkOdm/ru
XSgH/l5oyixMQ00Zac/HFYBecIKQLPSIyZ8Ap7HlWThKl8tO1DHSy0axOlJFd0C10DsjJHPX0Sn5
C9G135+ADAeH1HywpVQbT0E+gAZtSRxN7SuZwH7pzKliWaWU5SeYnhugKa6AX6J7aH/3Qfbcn7+u
RBjjLYhwXJETaK1hRa+BwI+wEB97D68z1q6KWPhlQMdkrBuPhCiBJZEGk/aa0eqZJoDOM7p1iOQH
6uHLKXXhtriiPSwADXdWi4ByP095zTwdLzlaLJbEU/GRDrbta3//j5X1dYsjiFIfxbdSXBdN+qbO
ZHixAHp5b53qJ8Zphs1yCrnN715EKJNeKTgHTnew4nntQSm9gj9Wxshm5/L2XvXS3FtG8GLcw4w6
/uyKTR1hTsrvvLl7seA/lFERBQ6VTpmqP0IwGMcW32qO+cL1v9CmwY4irBfuSF56q26jiL3FNQ7Y
MdsnTT6b6RSEIfrqOJQkF7hvb98nHe77aC4DLRA9qKCaG1h16bi/ZhTOGqXGGJM03Be5PlaEdTz8
y9LCRt5R7FURAXdhAj6znvnPORkaPbDdZ2n0OM3d7HCh4dzmLGbDewxKELDwpMc+L48QW1iteyeJ
+U+xvI+7FiGB7V5gE+QTmrFbvZ8c5eRcrWIm/djm+saOAuWXLXUhl9EsWDtH4F71Fm/RyTs6spDf
UEaUdVJ3ILO/glvlZFfHdeOZX5tnonfgQ+GL9qQMAeofdJPkQHAlcUT0pH9w0lGtPgMm7UBqtf7H
8xoGyWK0eEtJ9nRG+mHLj4s2s3uKFkqKP24NJteWfL7zdvR8ew8LNNzPfKAxkBNu0OId7+bMfYUB
Uva7bZXKJWXg/JQMnONwXB2AzTv4mQEqGJS2YRh+31PvabxA75NeyAFbGmYo9ajf4HTvvxiyR8Hb
FdQXaaSVKgFIkmIUeaAUgUm0PnVhLUV3JuGi+AhS6K8R7B5CgOzhqlD1DkAJ4ltFKN8xx+5bnVGt
myntkr4BKqfhWxZy1DpUaMw45ZR+gFQsPVYbvfUefz57lckz1xwCf0nggCJcdQQlmD0uhxuSNVeg
8QV4UBd7KsGmBPrOPoZJHScjCOd12e3K0xbt3DG7vymc8jfKX2pUbPP8j5n27xqDVyo4NLVIEjp0
IFlnZ3ZM8hAiUW8Ru5rzTHZ6aueGoTJhhCkEMIloosrAwZb/YSc34K66612a/3/6Y+Dso3MSBbK6
aLT7wcZQ8hmMKA1jhNJ9ttV7UBHOxOeipGVAQIUG2iG40OnuHgvTa1RnoK1xKTiTvQltsakC3F2z
CAS98M2htE00ES2zWXXbYh8NKf8D5pGKTfVwePbSYPB3kL+NDLXrMGPEjZy/KTmadzk9geW9LgkR
e45QLM6Cl6ra9X62oiu5NxeZRD3n0Lt+Q0qFExxg5S5+4g/9G8Jvd4KzebwsLcO+GVwPC79nc9s2
lGH4oW5eWNzSBFTiFF7oDIyN/lqymKqb8B4TVzqpdybSA1cot3xjU07g8XFgOb2HrVqW5/nGVhn8
IwC6vU8ZlHnT+zXo6HFz1CigUxJyMFwVDMXFcPjZKoaGWaEtoze4vzCi8dvANigyN3xtbGr8+APN
hOi3QVllWfu0xOE2r8PUJTkIGqniBWB+gdbNToMHYWJiVbHe6T37PSzeWfN8Ynp4ZscECCAvY7nw
1K6n9mwSo2jFYdb4nIn1uQH66/SJUEo0elbE5ruXnyywXcgAj5wAkZZVIPR8pFdocqb0e4UgL2aJ
/sDWC+O5WtKKZvujxJ/Kt+yHRDTdVan9HD8u8QxsP2gTmqEWKNxCmb7B7cF5i7TjzvQeStZMKczp
yIRooJVAhaA481+f3QJfqJpXy+LVjQiUL1qip7DwUBTMOfwH/5XPsTfOf6/l3C1TRrL9BHsy1c1T
pyxDF46yIi7Ylhd9R89+rWUG8xUtf7jD6NUQ1ohgNc7h6MOPz2FVtrbqGu/+TBFYLGQWl3qJEh0C
28wWmmMfDyYkU4kyJwkfqUUCEnkgJ82LofhWK7XAivDBkwo47Id8mPAjloT6V32yr874lgEj1lC/
lGUClLdrgC59Hdnjmefl+kQVQz+9pp/EX2A40KUYStD5hFgATwzIrny9abnxvaLSRguYIzaMAnbN
JwFt+HtsR3Q9/OmZ6ZS1cbUNM8BgLg9lLrePgZSx4YQHUddEV5yyD2UrJvPVJ9re2XGnompQlXhG
irO7dh0XvsYUnCjnlh77/HiTUHpNRlwoFXJUlJb3wdmqHmAl5BM3DmKcWAFqbVvs/SlTUF0Yti3e
0R16+UXPFkN5bYV5XlCVJlRm36JkkLEseDNJo7fdm2uwtpEuItfVOEAd7BCU0JO0V7FQ6rKodXzA
Lc/jvRQabNCD+P4I+wlFwRDq9JFjyZ/q4nZXuPGI2xgwglnV4cDWJmR1LqHO0Qs64A6yXhXikDoy
cbIeYiAcuMpgtaK0yRtVn4/0R4xWJQTVZZrfMYtFmlqCzWlknXbwd4PnS+1YwjMCe6rrPy2/h/Tz
4HoAPjKuHASIXTKgQ4OHuJWNo5HLoaCU2r9tUju/SthZF1MYCTmy189I2yCphCCnvi6X1yaKF9ln
T/dJNLcNiqQgCcOWW0fZ0I3uq4/MMoAa3XszBsEzLKLpEetZ+3OaCeXQkAWf+9lTd4f9ffFOweCg
xAqDt5GViQbMjp+vlEDKWQWyvtNXfZFFwQ0Oy5GFY1kjE4ZQ/mCPgbHTGIiIEI9dYIhwiycWmYHt
N4wY+hMg8cWJxbOgcG4w2Z9/ViNUZsp06yHxFvxkoIRhpMRjW550h0Dv2oTdhRSptmm1nYUNZVVr
BuvYWWK7CFqWIFqegY+Z6K5d0gXznGRXsZTuBgmqdIS0rdd9mMUqCsglnyNG2nUEPhgAswCg99r6
8J9vWRSTBLL06uHo/xgoxfy+cTgDWgnN5HdH0j01jInMrR/2XMz7JDP1uwWvEXbMFj0NghnFfBIM
8CKvr2sqw+JWCnBVyOhuKa5pX0c3uRSBj5+bNUDtVb1I7LXHO/kKw6UIV+rCwD+vRYZTusmce54k
UHKvULCneq7wWHIe5JI1weokBZOpUp6fuSZcvIbE6+whQfBSXSCkiYjqvXHWAPFU8DBW76pYBGgD
gWdlXZoUdvG3oPyO1t+Me3Y7fz6BXi57aT+M8NpquOiW63QrSfhyazduI1u7pZNAS//hauA5pXo7
3+KsS9AkVsr1SksGIVneS7zUgvZu+bT2j5DtP79uz126jJJ9xp3Ij3FNlAOFcVAZywghGWbXxMzd
Kw1irdD6xZa1GmI8olEizV2QVWcIXGZ2j7LeRGXfIPW/yfTyuqR3NxJF0Q0XsCvs2emirNSfYcQf
IUGuhbdKW67v0+XscnXiDueAbOb7dQ9f202a0c1owpe6xxzdaW2LOccHslVHoaAKvVVWPYQM3O1k
dbtbuaij5mnImg6x1QmQJl8/F75eHhcWXo/kOa8HJWO5U/n7JCQfV4guhv0X2T5SByXVd6ZcE6Yj
NG4DbU3uyW+TB5w0QzXlYAlQilhFUsbPQuJO+luEjhIlSn7/INZsiQ18MR2V4ruvf/ZuNJkoRkc7
YthXh1OmdVoCzAmwqZswIfmSXuSWUfzuA3HAeVPcwJrzRAIAquO0FiXeBCUjxtE7bYIXnQ8NKFpV
F7KbWg5OLducVYDv5Wp6DyChE8H6vSLJyITNV1W8Et+3r5tCd8QloEYh/qRMjNbkj4FtjuiTinuS
QItMsWiYoyOspFU6jYK+XTRLElN9bB8S4IyZeCSJEnQ9neLuRsMbpwLU02oYml9Dg2JHNRozyCwL
alozOaFvUuyJNQgYFEAOncZSJ3OmDy+g/tzohaneyIqn65b22kePnEKjxbaE7+WMFviTSP7Z9uyL
KGsI3YU9R5hUjfGZ9x0MbyLYaCnyCnDknPEpN+LsFtcoGJMiAVozOBRYlq1Wd/ZslCupqz2zkngx
glNqaeV9cbxqmh0OjzN4qdbCVpsbYlRaN1S0zbBS08cT6dkyPChyl99IS+/pe/37FDfMtS8YyjOQ
sOlPflLeId9M+nmHyw+rTk63owvY84OERd9En1s/4fV31UVHCexMb+Yfv5MWSU1b3IPIeshKSF0E
tqX3Yjfh5Tj594gbv5/74MZF3HY4nBP5axnf17Kcra6iuqTVDotVkbH2Aby6kiAM0s4US6D/jv7e
efJzHneLgfHuTy07DDY5JwNTHxoP3MACDVoODEHdamxrEtWZCqngEzC8545AyMAOuBNewa09C3cm
29UM16iNGn45nBEPdZXd5bn2i7ibYo3/l3B7kehUgnsMxbrwMiwO2bF4MxxrfkDwCRr9UoldP28t
0xVftHZdN71PP0x6PgkPkKcW4ZW7qAU8SgnOp8zJa1Iy2IaisSfYZET+CGiqiaxTJ7Z7equrdPNV
0pxF4wymwgofrZWPgAUtae/cNkiw168nmx262I7Hha76V07V+QdFeuhLXuGCiYEUKjoLGDDhcUyS
1EwMe3PqIiCr8dqtsDndCjnuHGvQepEajHEVFMu5LkF/hW5Q+I7z32eMJ86uvYuozDjTz1x8rI43
WY67IE1/t6AyujUb785ciyhrbaVoZlw4Zl5e0iZixdXn+ZfQDKMJN/ZocUkjzFlDfn/Eb3EDwSDW
mPlB7UqAMmjMnceCOVcJCCuc6zY3yXwGUUCASD6Ih8V+7l4MhsOQ/sWyERLrcMrF8A6ciqX/0tvw
CXcLny0qGKylqWSTuND2tGQRVDa+IZeG33+D925arkdbRqhb/x6BTb8Vcaq8nxR66jwuvv7e6MIL
MaRPX2/q6p3Kq7f4iDji3BiDr6Q5wfE4wCyQmNCjh9bEc8vKEK41UCbqgsfCFapEDGEU+2NpGtdF
DW5xqOYHJm5mDmSXRkquQNR9hIsKiLG4+VFNkBGeQ7oGIq6j00KDCSemtbeASUaYN7uGPHGSAcET
BP3Z43NvLgl8J0B7IhD31BXP9qPgjJc1XWydYovEoO5xehathBd6roenNHMKeXDHI6ThRNe7ZNkZ
F2yzpePUtlMoBqaekMzOKup6LvmxdMCC9m/arR1KLYqhxdM8+70PxKCcixTfJ5R4pYs+LN+ZLI3S
/dVJfXucYmFggkXpNE6fcdqMuioDmZ9mgfF27eXkI4HxzV0JvkEUkbrdRthUSxSnfV4QV9IC5F0C
kdOEFLHV0RrffmvEt+cgQ7FqEKg0E3Yd87QsbD3h7MLLh6nDmzWAZSVoIXa8EkhKK1NhXpRLrdKP
eU17at2c2fqGnRqR4W30NjbgmbmWUPa4elCLYj1F91/DlTBaVJJZM/0/KLY7l+8UgGsY6b4cmVqP
2vLUxzl7G8lkt5dwiqfTd2K3o8WrykOLMhdqBexb2lVvNW+GpJ4vf/NO8e7u8mypb0tHKfxJllZ7
5ypRbBH6xwbfgCtvDBuVK6ejZhUrptLjodzcUXrx2oTA6jLfAcopi5d+eXPTewhvyeuekDl1TIbw
WMDjprYpjetqEVwGlHYGOXjcYITj5xMFU67BtbjRL9IAjZc4ruW1jnjw6bzcKgNhCF7zq+4dZgmd
1ZFm3pEkWKcx84adRQmF4d3T7u5/5DpPa0MLl7LNKmajxoBa7zJlNvw9JANUGs+hXLVtgAJ0TE/T
igfAGEDMILk3Sye/520br0bs1A2W7WsMz1KBIG+YHu9R/yfnRZQoC6J9KTZbxNJHFjphuDP8QXrc
hnqeuxjPlLiNE1k1/9bovGXMSZ2gAiNWShiDE1NCYKFURipJVNCVZEymCgERDwxPuaejEoSORb36
EK5VywkzbmEX7k9fHDYHwe39L9Yh8i/zifVaBP4r6Dve5IoyHklmUE/hJjhDXuLgIrUHkh5POneH
ibA/Xmhofa9qoFi8O5RET5vorPZFCLBD0/WgSoHOARIJgHwIVh+ToNl6h0cFA+77LZ8e6GwWDqi4
i6q/EllwJEsZx8KUqbL/7qC5KolRmKHm/NaJi2W1F7ZKRiTxNzzPaC90+29TZhKFENIkX0Si9C9r
V1JSDju036WAk0zAggRB8rccHCyQsQ98pTt4MSToU/AVSBWkYQABbdzRRcbANAqViDiOAfMSeNFs
+65snTLhB369wIaP8vlfY7AwkdWvqS/aXr+WoB/EJWHfpUwSTjceVrdnmdt+Z7Cfo+rlYw+VBOBB
SDszkBXFj0gSHF8nM1bKiGE969H7bF4duaT6WNzHnudCOwwJpC8PPyuSDK7FMlqyWP8uQCizSA07
uHNVOJxS54eTaLVq4NEJ3soEBHlkHzPDK4i1UoSfOYeU2N0GBYVMnrbTJXShoKcYDtqLygKxn94j
81lYSCKDc2ILIavrhnHVusc60H2FJJ9CbD95ct4x3TzYztJbhWAkYGmeJ5IqBcVxJLdD1/IYxKEU
dcdLO4/tP0glgzr1YtWeGlrGe62Mfvs1Ld89S0JohWWQJId6B5QOWtQ/rQVa5sefS1+PNr2dTs5/
NJjM7GdU9wzkltmTvPpgoR6Cdk6nDvKIcyEs74uqIyL8+wINqNeINDuUvSG8fixY/kPbr5RtnU83
B7SDhfTUJykZ3Nkh6En6Ow+bYQkHe8sWjaV38x+bsTnL6hlTW05vra/Q9jedAPb2llZx3JtIq+SL
3Ojjd2Y1yKG2hjKySM+OvIC5fgsgs3SYYuqYhN6kMVjnK1YvgdI+U6KbIeVgYitNkkERpnShu5Hi
wSxIj77vbbcL8ywwP4MYhivFDuNC1dzt2gkSRxSe6t2oy2cdUMiROZIuNGL+S/PMkw0i2VmTdjwH
sCz32oetM+nysfFrN+KrbaggC/t3pGTV4npk8wXIxo53zaaP4RcaHoacqZklSAeAsvmz/Uo033PX
eKnQYAjt0fylKQX1CA/SPI3rxfMaf4YeAuRolCFyuyc7J8ibpPZannXTY0F/chGrAzWLXoXTMP97
yyutNkUnhqYIMuMKzhzOuk75JbwKe0wRa/iyHhjcMlQvyh6A2x8+irw8ys66HVdbtOXVgFzMHDR/
fEhYOlP++F7gHJmv5rK4W+WD7gr0PMZXyIzBU+C/3Y10//svL5zSaVpn/RyLreQH4vQNIQM4SsyX
tdJfrur2MVxk3cnMCkUOjMZgiUDgCiozAODQ9em6IajyyQOTtkUc/iXNz6rlEvu9MRSBz1ltOAwQ
ocQcHMlfSriWefmh1y/xpqISyV3UtVrypBoUwM9iwoS54DsR/aeIodXgpLfe++PPXDhU4wCv3yT/
BGlV9DgrPpE9rhwklP3OXX9ahsyLfvvJ8dlldJNZimiIU1spc1XP4gLGMsYstPj9LaKZ5KxPHJN6
yXBWMDJ03ymg2RPcNLajBxwaIjdn+at5V1WW6i8x384Q2dpmNkdAXhjcwL3K70ed3w09EJ/WJVBm
6sg87aumQlH+ESRWz3V0lD0RjPVf0cOeVwukLOGnCPd1dBZvwTKF7nfBGPWRCF2rlNlGjvkJHpPB
3+HTQmXOi4JCPRFhOIWIc5jnzIuSVZ0PY5C+nwwMJAO4fA42MfYokIvZbchTuqzk7i11PrBtO9nu
2c1R4KLJCdqN2VdXZSbEMDLyAUbr6Oa6qvqTxJ2hSATz9b+Ru3NGnXB4hurvDFNEDW6MsLRMGacp
Aei5HI3gAZ34AZpaj6++R+8TKmzdVkWVrlaRGnX9p5iR2g3CSWKVyvTTmDJWsA2jnwHkEco0q0Qj
5M22N0pLwBRbKWDgPpi8QiA/aTJZhNYoqfOhX26uY1s8Afs09QsyxutIlNwgiEJPkuu73Aiha7aA
5W3Y7SLTlFdgs9nYKfCwsz0W3MPKicpbQ8nd1NF1JVQ+6bdl2TvwNxZdQVP9G+XNjZ3rNbGukjh5
oWsMrPx18SZNaJXU8v0UKiaklwFsghinDUBq1UUA/dssJlj+qOxi9MppGZtAcNZV+lHJGPMfsGaz
n9+febNdzwiqvQyLQaWAmx8ucwbTh2FIIpd/stTf7WSlWq+13yFhK587ElRxz1KQ4FHUZv1SOnF3
bwD4VDGOn+3QzSrSw4fGuQr/JZXFakFWu8KwT9kl46WI+d+zwFEhYAG4kF+pMtxGIls1a56/tbGF
ZCRE+27bx7cx1Vy7nxy+DxPqDc4O3iG8e6VtoTJjwCPCv8n+DnVwZyCbnkE9E5sd02XmxVB0iObn
RC2E4y/YXlgwc3rJQRPRcoZ6lBkvnrSwZJlvb24pFPXi/TXctA5bdgqhmzLObxNVDkq2a1GzOR/m
wH1BWX2TUnQ+ghOnbH0GOh7SrIvz0XS+VGGXB6rdSgrP79Orw147xWhvOkQ9Caej4VgndD9CZFAe
k5TotKycWSkT2URXoc3Huc3AQaqpxiOHzilWnQHvyEMBS0y/L01yEjUFKjh1cigDD/qyAPIhRLPs
CFtMMJ6rozzU3RPHqlwzZcWDM6u0enGcnrNGg/7rOd+QjifwL1AdE987lHmGFyvx7cNLrhr70r6B
ErnkUB0XG560ZG4DR1cIhl5d6J04IrDoFn5oYNH3eWKmYq0i4dBXI+UmL55IUUhlttALZNlApJFM
gAMCHn/RbK8xU0Fndbp+I/203nKmMIOsSMDLaWFUXJtqyFUZt3dNNw0P31P01y3OXxM3GCf4Y5/v
JixlsSEvcKsdfd5YaNzQLRZMYbRrr1pUxxLynQ1VUimFaXM1F8AxM3D0ELdmXUkEB8wa/8AFsTai
MdcFF5P2BtD9ijCSOHtHXWWzke/zz0IGTctjWgSIjJoMEpoV3MtWYo2FYW0Tb70lKnb4eNMRNq1k
pR6hV3QUAhwGgAgjvRKfLt0siYwkj8o2ldFinA9/uPeSw+cErvTLBD0ai9tklhazfot8da1ALINt
2nxmHptyXh5j21dAmmIqUBKGubGAZuJebJx7Bn1ZHBmoRRR2Yxcg1ds2bgMnI1Og8xNuQk2V5BfB
9zuv+t51kydp8oXpobEXEQZ7enltw56vpOCHAAfIWvqEPvguIRXlox9Sbsv3YExHqXVTvJeGB1vg
MP3t3PynLrw5adsIv7HyHDQuCKzOjLgnNsNObMNEKuAHdrgC5KL0bcms7tdyPCNWOqP3Qw7bsGNg
LeG5xybvf2N78MZzfYmMAhKrHfNPF/wZDR2H9vamYsT+LNyvWzVueRyYxMKjKALz+Z3EZvbWTtLu
6GrgrAPrME3nzPvNKsJq0B3byckQCsJBtntxy/OE8Y/gMcTb91phQ1d5LkNhmYqwpNbM07VNR5BT
4mWzCNgq1jnWZZAVN4qaLXcDc5MI5Oobk3ucPPtEDUhBukBSlkbuzjcg0NAsiyADL5eHUnK2O9qX
u9ihFjlErnXjWZqlofhn1O3fIAajnoRkEXBWDkr1ZZry8/lzF/njwm+Gz2EZiviHoU/xm8LJ2jqI
hlxmAGDKJXhKf0eSidNj3rzEppiSXTQPiqM1RbwnW3XlWij1KRCI5VU4Y+97ZL48aW46DGHveuBM
abnKKC3VHCjSsZyR77HprO+O8elwwfA99U0u2Zvnc3aQ1ofh6eqyBFacVL5FhJP3i3OgnN6rbb3K
LAQFplA6a0CY1wW7HUg2XGxattbxVu7qO2mMp0Nxn89Rv/Z+0Gt/UJSrwKHMU0WkViL3hH5tL15e
f33YIXz2e4SPL24ZvDtBygEsfbV1xqfCKxuHLMM5R39n9MfSEP/SOW4x4OaWoV0esYMJGhZ159WR
MbCJ8tYO75L/BJw4m+JHaIxxtpp0tPC6g0DoZDpLwhCfRHg4aDvfdM8MSPc1bsTlmOYvEd5/il4/
S90vMH8y6QEo/JoXL7Y2YHN7eoA15vojL/tBJajeBEYQY9UwT4qYrYRbmMit/GSpAyokMznYdNtb
WNSnNBPXZylc9MRU09pFlpVekxd3oCONFPwfD+tlQwZPW+y1si4o4NV3gpOCg4Hxfai7/jQKw7Ay
jSEbWzRwHm3ghZaoaTY7XX1El2gUTXYLXpy2S6isEZRAX2OjF6LzGdbRmNs9kvGnDHU70beBehj8
Wyry114BjS+XAEKWuRKYjUa+Ky66FajtBkQQiTk1e8RYfFzqQqMBLj7UiMbyzrCRpyFWLPksfTkI
EizxP+ECk6MytEs/K9zkGAJzNLR3sTlzU/uZtA20DZ2pFH6IlRXc4mlQJ2g4d7NtDOlxbhXjgXSD
42nanQQKxu5Vzg4nWnq5+K9/d3NVSsz1DABuEdZDxgwsl+6HsOF1UkSREN84MYMMnatSNJu43EY2
HFq0bzV+WhgKTxtOTWDvg+uzeG3+zJvKst/Mi90LFEXE6O9K8H/jvHrmvijRZLC5jQzYpE2fiSdz
OZZHn3I88YrkRwoYBde7z1VKWqTcxw5iZou3/HjnqlSOASiSSDa3p4kq4RMhr8+kOisxOsMMBmPM
KmGwwDIik2fZQgHWP4BfMWoIOnUeWZmOPtlxEM9ngRXStU1rLN90YSZGyIT+wKCjtjlm0cbgmHI8
X/CV3MFVLgydKxQClq6UsUh8+PDygEY1cKPVjiB1IYnfkRr6gde51Mcm16XEb+/9l2rFuCvlTnTx
cIEzOMkOT0s67DjXaBWYVi/hbu3cBD172WT/aderRLR2NXPClo7ZZ5GIwCbVHH4+rwAb0M/APJmX
GaLsvVwGXy04R8Qil4vug4xQYQzFuEumDGAGpmn3LPBA4F4F++ewdaalzBPpMb0Q/sylbo+gxREY
bNi4RFhsvdtZOgoSaIAnnaNWKSDHW2HGqE43FEM+U9WRI5uwL41vvXJIYfwlit4pLFLISQUSlW5V
t4AbyUy0KML+gkTNhYd0qf4qYRdwM1g+0DZZly2S4Sk+U4itNyQALKOwD5rN130fkxxmBaDhxA++
BCkoyINrWPMtj6/s//A6lfgWX+T0xolSKLgdktG0iuQ4XPCroD5I9+YaMp4qgb0Yh6yerTAcGwco
7wgLuS/4nLcvNi/ix8eu2TFV1y+MWFpCWVPP7okW5sv/NZqznPZATVHau4GZ11LHYdR0BJ9B3aLT
HXhbzLYM8yLgY8E7o/w9TIYbfcPYgEvFiq4Ug0MzacZlvKVFjmksbqfHwKSsPowU6uDDILzOMVTX
YGz79gvTg0Q6UwwuekTnf77kuPGNZoscYuJ+s8NnSYgNLUdiobJ03FLnOMyd2vhuGgpP5UbwRpEo
fff/cwVc3g12wDcx+v40HsDtEVh7ttCUtrr2+BkbLQWgqLmdr4KEUORiQcO66geGJDA/aA6I3ii9
fGOlN/K+LBa52U+wQctBBlhDmki3DxUhFm11l+mrDsgrgZ++WURG6YiV+ozK++zXeWkBDO5gTMTh
DBhgwgvIU9ghmS5wylfPpBmoNoFtWZTPx5a99+kAZNxUzOn3zdLVIAP6DYxN2j2+GDg0dJAgwxxM
yvbkKF5GxU/oLCaaoEYr2DYXyBvFt4MdNcMFkAWrdhIqB5eAcmM3t6w3wpXPozAaYkHF/CkYOoim
PwAKWZ9ycX+70tqaAKi0+897Oh6rZVb08sRaZdlNpeZuAwbnNsWbz7jBMqdNAYdg9rzdGSq8MpEW
QRSpr2pDaf7c/bbuzU9zCYUduI4BAvjIJtOOqfosRfH2JLRyH6Fpc5xw3atfN0FklLfGJOftS3jj
JdUNAJFFkk0TUBpuFKQarU2H12QFBUgdnAT1GaNSB7RcyC9ltj/1fOq9QmzhJpkRVaSJmrBJAWCD
T1XxashnfG3o9Q4rOWhvXIMMTeA496pM7hLkzrCGOgZcbMyeKHOiZSHHpJ0zEgKkMRGkc7AXb2JE
sTzAqKh4CUYIs7JzSJDx2jKJIuJ6RGiJvF8BkqCZKdoslpJzfDXUQCpmNaOwKGyNCTV9tbkvthy/
4toAY85bsHY1JPjIJeMLuhDqke9NZIVnQcypHnejlCrQyLqVfivsiFpVw3U85klCU+k52nD20Hsx
z5WOyXm1MRU2/BZRjBk09jWQ1sXOclu4nli2wHZh40eYHDI+nIAmjBtpaGRhP3GNunhvhnvFjofc
JvZWrnjFu0UbLZCr7KhMzRe9FiK3U3Ma9iampOWyGOqcYFVJaWo1ud/RsFz6AeSEqnK3KLq8vIRs
d2CtF2Q/XIIrNQ9wz0OW0ReYYbudz4v3Vd4yOEwfFNQgz6QoYm2J+Xsw4rrRXv60oGEhhfXzkjQh
IQ+6AoO0vCrkER2qgsoHTHY+xUpW7XcVIPMCERV3ieELZhp7V2cruIT8UtRku9AlNLX4Dqqor+gB
8tzrSQYQlEpg0R3sQLpIBRUw936dcfeBL7igIAILga2a0jkXsc6O6WYIY5aEdWbN9ITg3mYK4Rey
HvkbN7Nwpicq914n75U0sflKQwvtliFxKMfmVQ8wP6U8cQeyCungHRAFZJLAE42VelClaR8af3xa
pBAjXR19kpPbqM1ao8iXYioyYOxgCxkGKJ964mrrqOjQ1j6WyJhrFCQEPR7Hs8SQBhiIGEfNVclj
s+1kSqCrxV4AiCpmHA0LaUdi1sgNJwZ4E34lZapMm25ZmUi8iee5EN+FiNEogy8vCEv7OBivCYip
kx1SfYuErSLW9fU+d0ysz6Bi4enZg54JdUQeMNCAH2wJ5C7admaoslwyegTSrKbqGWOMvpM8mzQi
MjFFqcV1sDbC/4kEDLl3EdstNXxt0HEa2KLKCus0iWlmCEB7RJnKg7doVxDJpDKiLGZjqZljL16a
UsptpZhnfcXYha5xtIPR/+kbnGsX/sumeiJfdiBoT5AoS7vmqJstJ3qmR4OBZ49c+5PYNwyFLkyh
UH49Lspjzg5157cLATnB3sz1YUX49/DpRc3ISkCMXTZhzV905RkN8vCaQtqiqoKb2ZI68bkBqlEx
wiN+Tx7sRIDBvNpg86XWEGNn7zy9YbDQK8s6WAhzZvKmEKbv8FSsOQIA+lry7NSDP0Y7rQzpHksj
Zm+/T4lw20Ja1X66pE7a/A3eTBUPyYKvUAdjXBOb4lpfuNezWCOZVLTvchbihoQQQRcAI0acVlGY
OhHfczmA7YM9iTFZKe2qVzEhd2wBdUe/BsAT2zQ1B/Olug0fXf6shrtDh8OwfscVnMoEKItSKI6R
nRemQAct6cUTTjBEsCE+WVnZK/yKBJilQmmHLA9zo2OaZzODzmCC+9UDt5JmkdJhxKsAdZXA2JKe
5VW9NW/ocggpuMqWPkBiRyMc1O8c8flUwYQPrM0UdtFfwIEcCLfZsbpI3012tkOHG4d2PtC/8l13
5cjvz9MOrux2+Zj8Ow5zygoquSGRDNOfe87rEyUPu6gMvJC1G4t4SLOXVSMJS4MqSWObCh+BLtl6
99e17qEo8+Bjpu6ttE2nJJ5lOq4hcckUv79Ot84Zmu4h+dtgmVpS4LtUrDi3GXLR48krZkCdTR/e
VKgfbC0Qv99OAw6jWQPMdTVvWIRMqdLfQ8IeAwY9+KA0ZIXnKMh8WDZ6pFWmPUDWOb+v7NQj9PIA
Z8QkUiXDrIBHDa7GYda6suqL7jo4Xn/W5XsZ23/1XBpy7DuvwGAZvDlv7NIuOkmN0p94JJqPKuBK
Lj39oe0nbENQMfjM91F+NYjaias9y9IKBTwPQpdo3318OZPXDjLzN+umczaWDBsX4PhTKUTLzHGs
UDrYO9rduv0gO00E6BwNLzJOLo4nYC6Dfpo91RRzHzOckSWHVR/ZWc0Hxoc/kabXbpZE147eecrF
qbY80quStlhtIaE3FAioUQGHywnwUkcR0mv6gCjpApEFpWLor7QDbpXiBPjHsP1/cQ6tFG2b+myy
/Idvon6GwtEyp0VTgUIRgebLKLUiFAxdaL9uOrg/CPrKCkKy6JNIzUsdvDugPKXr3Xu5lwMARuXk
VuPsGjMXrUJA7ESBXuApxKUhJhj6E39FNPZPNGYjS8XeMUL5MFkg9UcXEc66gazwk2lcqBJJNgDb
Lm6EWrAAAl+ItJCo/Fy6bgm6UlUUquQTDo6qoAmsfoUBU/0QOg16y29f5rJekuXUvDQ92G9lqhxs
joSo7r+fZPFgENJNCjkQPBnIdgXljeGuYsSbKYDwCRE+le6fNQgR5nI91J6VbmevQOSxe8uK173P
F5o5rwWiI9v+uFv5wP/1Rp9T1EYgWvsf3hMetvGJwQilHyOmrBAVy77CVj6FUWIH/kHXhgw85hH3
H9CYUskB+E+enwMBMlNb0dhFEoXBv5ytVqxHFltOvRYkVASec4m9D7rTmbC0v9jzLYyiGmta6JcP
9oQ7QN7ZCgpJuf+wqjZAvpp7AFW2zwKjHpQd3SPkGgBmheLcN3frrd2zymQlT7ODyk/K9rqyrNSV
sI3nTwCOjc6QdO2fGwg2YpJ/cpYX3IZ2E+8lphcb3UZ2upjEZg7S4ESnoyYj8PmuDozYYsibVNom
47AgI45osqsZ3I+slGTYJrvpZpvq8SsRW8R0ej7pOajNcge8VuS8FZVqux1DjiaKy19gHm1MTUn0
zXjGDqZQGyxDBlew3NNLIGAwFx3a0lFghPBgdwFiHoHy5q4YdGv6ljzC6bY2nWl3+zVXlH/mBOPq
XWQd0N2bFpPsHEV4EGeU2qjsJKqf/wPICD1lrIx6nOHu5j78pg3dcKpNUhyeZ0LmBpgSLOaroAEJ
3CwW5goLcLRb2dL02+wCZjHbvZE+Y3JNIMvOArxqutg1yVJqd71SJ/16hFGcha3LftKlPROs0n+f
Y99ZD+hEgCkmEEmnemwgKHORX60kK7ZJE9BSq/UqfBRHq2Q8L+iR5ZTdPLGR6JG406Ka8jv4sFaY
rQhAshIbQdtk0wWkYOvv76vd4Yo9zZVCABk6BaLNe7oE7wAWmW8FqEB1pLLqkSteco+y2uSI0OD5
2l3qPEPa+Wf0I4urfHsJKaqnxaYt4hZyhKntPPhGPLkvoIUj3146kDlVmwRBpWDXqk1lIvrBs/q2
Mk3Gx/AV8w0l40fxWWCabf40x3LZhvukAKbJlK/wXuHyA8e7kW78qD8gQO1Hb1sJOaiMxW6Q3Njd
kIxJo8p9viAWxpcTBlUybrCNdxO9OgMxtjrz0adB6R73MYPBYF8U4qQtb92fEB//9+CNFQ0YPfwy
xfZrj140qND7UOHChrBSzmDTOZjnieKTD30xD/7Jw+8r/hdOoN9jnLOvEIMnDysf2rpY9seaT0pe
ftHpwxXMI8LerM3YdXWk41D8PQl32P8fS7BycTiMU9UVZK71Fo9tSfX6G7r6xXXONFwuIfzOFXf2
1hgpWV38PebnBk4RCkJE8STN8d/rpxaALMFBTIxEA+5XYj3lRucaCCIJ5tLHA7KH9D+03jS0e4pq
hW4C3ktPV5H+YCQvDHYHfgQ5VicdOmpAjy275bJB1BqY9Ghr27CtHRI43uhr3Q4n/TLWB2FTjS3O
pyxS4ZaK2hS51jO+dLWQBeMs1pgxVbiyaMgCHnaCVoUjrIcOKQKgCWh10b2ehvFibikWKWRMJS3p
FOs32yRHWUY5aMZYDFDVk58gm8gDoGiqLwNE7UFlrS0ZOSY0obTx+V32LErZpiwFPd0Rkyx534nA
+GmQQMDiF+pYLGhoUI1T5Lvq0MnQvjQE5nb8je7sampDSpEzREjNRB2CRVZwXxMsXi4xtc5pi+WT
Qne1+kLuwPzwhsRe+UYBL1ZViVyM5wnu32mR7/fA0VEdrxzmiUP05N7mfcrh/BLwHp7kG0PD0Emr
gwDX0kdl+k9o/BC3hRdTYPeB/mtNvYNCBLgYVOOpl3NYy0U4JqZNoXXyK/+qyRt+7hcFUyEmmoq+
BNoGeWznC6ml/nRQ17hSf8X2MNcIgZUvHbr3NLZSuCYYnlsaWP5SXan+JTDGP3y5KBXbvkZVPOvK
GGv+zS5HDnWAjU+iW6D0+vUMqqoGsWv8Sf2uEW7PnpUGBmgrczLo/i/h4LqP0AJDN3NEvJt8yde+
GZSIx3JunqkIYTZKvx7ZsvAmGPmNIr7qinlJI55ELSCtSJxGcxRoMLbizZdrU3jJYv26dsaPJeBg
QB7/uMyqxjE6PQzVOZfIu3u4TXGEdKeLW0slZ1wC7ALIh/vHgzloNIFldo5qcmgDAW2Ro0H3UHAr
0izq/Hihg7fD0ZLv90Oj6CAY1TXiRhgM28Ct46EyNmtp36lxex65Q8duPD3ynUBTVSvp4uZY5quA
2U5c8p46UJwP3niY+mbHpNagGpVJCZitVSFXkbcHKpbgEYseP/LpkPaRQEqP1tpQreU0w0Cb3uqL
IV0Bvo6Qv858XcURq56cOW8ROJCxTpoYHSq/PdvOrQZTVyFUM0M7NmDERS1NZjqmxeakzHlQ33Fp
mKsyUIpcPe8rTooaatDOAsHAj/5cFX93okGw8blqfi9YKDAnZQ9gH02skwUBQHuy+KSg5F6CWBHc
BR2zI/AanC3Na/HwpZdSM+j9MGfOToyCJUvi7gMOjezQmviO8T7dHUz/vBi6diZ787qAu1c1aX/S
3Ltdqs9b7/l+Dpxv5IwxgOTpoXWRVasHdMcXB6lUM47AbVP4MIZf7B+aF3Hb+MRD9CzdLJvfZvRY
v93WamtitMRWCfzy/xbYraqKbr4pK/U0apl2NrvzzuT/MdL5O5WL29UtSff6s+N6gcXe6w3k1ogX
RaJUtfQNDEvSioNJ6IJB1O7dlrTT+1wyJDLxr3dbCY5eUcxzQnqwcjrDdMtWG+KIXXykuzulSsgX
aFc2syZbRXQjx+VmCz8u/dqQENsuYUfQ0xCe48F1Hkic65wmd1+XDKiMFuA1kF7VrXgTnOknMYP5
1hJS0vB+t3BLH4BcTI2Wwl9w8IkoCoPqnhncABwdUIxOIp91K3O/xh1OwSPiKxm8vpwT9V6JWgxA
hG1xlVnfvHd1cKtPmGVQSb/pDlsQvs85o6Z55C8Jo6OYmS32l0geKFb4/tidGy+XW1aNRB+pSwiz
RHwxLbp3LjKwH61MbqTtsap2EsL7nP7MAEz9GIRGOCyKLcnjz98hhjn9byH4fCUcKx7FFb18Pgcn
t+k6uIeRzjzgURj8VAfLvVD37j4FGrTjGx8q6JP1wgloieF5Ovpq8JzMbHBO+uQ/c+gufAwLp95H
LSPQl5wxWO8wv8Pr3xNmN5DUR29h3MUUgATvsVkBtVTnt5gT98xXEc0HroyY4NG9UOca3C6Czppo
LaTlrk7G7bx9sYaYEdb4kNcRRq5f05Dmv8cYsms0sxMj+6SjMym7TajvdikWdUVlDQxnL+p+LuLK
OzqClPxbi9XsZO03QVvPaUctaT1FZSawA8glgvYkUIk7TEDK7AK/vx0A7ahmQ8JRqW4EAGP0iv+N
8vGzM27Yhwb/d8mFjIESqSNxMHUoNiD9yytGyyYAubyUDKr3OLxE9ijhzS24QRRIsSLC3JfzO8bE
gv6Iq7Mkhx13LskiGf/LcKsH0vBs19SgeH8wat+rNtKyY9NOjqbw9AEj4H2rH0hI9N/XWWt3/gEq
8SCnEdCU0OhamwlVtvdKGTYqVrZzUxhbyHo0dlgQcK89UfQyJXxh+yYxtO/CfWa69X0UpCxG5mVQ
V/NCYG4Xdvd4X6E0iAzIRgwpcxv9FQxyAeoJupgFVK2LUSFB7vHarAMYI7bXg40sxKwdVHpU5u8J
nJ/FKJ5FN+mIDKCuKrEiqTa8YAQT3qFJ28y38Exidhd9Z27vVBHEoqgDd3nIeMTMNu7IIK3dv7OE
BH3gIjq3jBkfRQBJOyCa245UNsXYcJSLeuVmTP3wq76BW+McPax87Q8rcQrAUXwvLkt6WzpWXOft
VPpe5Z7pz8KfKdEg3p7OHgfeMAlUabVdeYo+u3MIvVgh73aSQSsgbtq2JafD7XHnxg1Fn7CcXksC
YltmoaG2G8D3L+nytMm6efiTwXvGKqb7KFPRzTCYpp27gSjzhk1Xj6fygwCa8zJw3+otd8ebvwd5
h+j5gYqrvAU+bY74uuo38yALriPFdYs8SYJ21IFYr9Oqk6vBgaLeNTgtg93fsnCF3hBH6/jEd34m
XRao2uk+EUMIJShXFR7QmsfmBzDLfyxiiLtoKvffvrVz1iyGB9scos6X9Z1dckWHrEdIypURy/2T
URiqGv2WJNDFaP+U18+v6XDobJ+kGAnIyRhxHYytIhQVmAUr639ded/EPGQM42jW9C7Y7hO3dp9j
e+NxOpOEZiT0IXjITr0PwlytGl1FlsuxEjRCwZDR8KwkZgETA+kzjhdOLizue7x/QBdLP3fi1+sq
A9jTsA7/F+H0TGvocL+nc0itkl4+KPIt5dCfCcU43huo5aFTf9KsaXpB0/74BKUE4Ezjyb0oSRzi
vu9fQ0sVK5vedVbtUUA+qIoIijuyJlbmoAuYFi1FDaLFZe9Nlr73cRsj50JJzu5F+4oyvCPXRNDe
DnxBjf5cr3Tjf62O/UHP2ycbIBvSaThk0Scn8OJOfdKJ9QTGG81GA4ZpHmGHOwbPHyfLx4wNU1Lr
PNMFbCvw3HXu5qTS74AbHQiS7k8w+YEOtyKmU03FqNuhbhFEX2Q4BRAPj1u3L6EcU3DjHbUowsyD
6LJgja2pbPl/JPBb+qqpAjFwEOnkyMuC4NPTL39TFfKK4auXH70RLPDHZs8wqByvQ+BIlgjmDgyt
eLlNU9kLtdukuXq62xuThxTMP3d4giZ51jndji/SZRHm6hmDZQTLmf3oRGbOFVfzinF8/UfGYK5S
f/iT9ognsdi1x61q85hawKMV43KrQ76ha7RYufI9G0IPJloYvGMwUIR5Q29+s817w/PtM76tF7dW
xrKtwHjdRzc7fcWvpkmvvttzSd7KywIJPQRTeFPYNomO6xmL1mgEnZR9S2IrcKRCqCeE5B3JhYo1
AhQOyd89R1IScWcxK7pMRjzzxyPZS7Gm6/40dKYkHd9tv+MyCOoaLJy8BDJQyX+wN52xqLtKlcS9
+eGsWZ6Fo2WpDAECdsZR0+PgF6I4FUoJ/HKwsaBfsAW7p5K6uzLnZiKtWEetqfQjMVZv1KcW2YBP
H5ai3PuflYk3zxtW7VGDzAA2YbJBeLTl1rdqGnj3HZgK6NtvdfDdkxPjMcMy+Cs9EWoYJGYZOKCU
bH25AyrvfUM0B0pPcM7YrWtlQFACS94fxYmB5mGNxxRWbKX3L5XZJoAVCaEd3gjVweSqpb4CJVjS
XuniiFGI14Ot29PF7vwmZeMEFGF+28/IHGNUY6Tb1uGifBVJ31spwnrRf/1DgsSVaEZcT8Di0BIp
YI3+2IEwrOg5kuutyjg4jFiBK6zDGaSYVcQXxu7pTiphgJZdRgRiZ8A/65Csxjz5nT9JBiwpvW+g
93U05NYXFpq8vGZD8iDej41MPD12AGJHkcV3uVPxm9/lKsqQwBXw9SwMniCT7hdphC6lPrMKg8TJ
gTVk2ZGlVh1NIXsv0yVY0+wXbjfls8PUiZ9im7YHOH3WWbGcs9xFrGIBB5J1vUp9EbWlvcWuyP9r
+sZ4icGpW9pGMJA07MaUmEJxJWDw2z3KtEHawOMbAhDtizEmJxGmc3HzALW+ZVP5sdHe3rqfxBeg
3G7Cdlt+bvZjBOd2oD+Pymc56Z+zGb+2dmZx5xnE6+VfxsWO+SLwN2I4R3DycRdHJBVQ+KI3nlTJ
msxgFCFEvy7A9izwfhH/tjw0GdqymIynZYqr0bOzvbMSM9mQgOp+dpJyo5SzELT634+FjND6gcWj
5sNINXUS6jtC2Hrr5Z1b3TJfd4JaXl97MoL72YWXKUBesJ7qJdkCEp38sKnWN72U6EuCG/UCvwRP
O3k3NPaam+lQDLj/H7k5FGZeYM6UDozOLCfWtPF+Fr7ck/6NyQABvcFy0I396E6PYCDq8iaDmy8L
Fsr7Ut3rzf3kyWFAtxwO38k4GMCE7odU8ShrZ7Qxwi48OfGNsv5aJo77bM1uZT7AxSutur1mZ/cd
OI17gUWwHTblpjstwgVbtf/r5Y+cmRsEUzjbUfEEoLvFi4L0A4Bok1mXllJ10ulqbv1g8Xu6m6x/
lb8NZLEwwvayxd4Rw+bp3qsb0s20/5IhLi6xafaCqd3V+mi71Zj1aI9cIXUmH0M9H9AZcU02te04
DkVMC9tIeqlEHb1ZBQ1rFNbvMfQWz3CScfAU4kmbbmAONebuGK0WIiZMSEJayc9OPfKMWv/f1sb5
/EP+RqIwqZaY7aX40l0TIUGgHhGnneQotCm8KjuqAtRsdk6YowfWK/PV3tt430HC+WXCSax8/0dA
hf0bjm/gnkmxo6NH5qQzAmvayRfHZoqn/dgUB1eo+dmB8H7ETHVEq8HRNoFmz/rnK8Z1+VEcIHvD
Sji72TnUFKao19eI2nr0tDLNXS7Mzv5gKEz2Lnc6HJMgaAnNEIBh4ysHmBWgpUGWpxTHUc6Y8SjX
v9muiI+6Vd9gv/e2bXbqIS5s2d3FGKmYM67sKX5rFeZ6hE1PGHo9voUgAfBuHIVPE9x6LUfjncXu
u5RsUG46PgCvVmlMHwx36Z0VkgwMHszoKI37uDVXwnnLWm09/iZ2Ld979VC9eRVSzzSb0dS9jNrc
iKTyrYs84P8B8VMXj/1DGhoc0Z3OW4ZT8wHc0TO/7BzN8GcqNHsIKlEqt3sRF98t2jq0Oeca7M0T
O36xupS6aH5/Y68XRNLFsROIykO3PvNStwza9jB7t88tC1A328Zv1Qb0Rm+/BNsl/b/7qXKM2MI1
ielXHZnzZ57amUwmT0f8b0cD4ZFmWE6rKjLJh1393C8/7n5vWnp0ZUj0lBu5bKOLkVACLoB7YFuJ
g0CCx/xm36kiHnyTbDNQEdMEG+09+vkz0nuaq54uFRKtTarb4SzzIlK36BkBOE9S6oe0q86jolhD
2eYHj6P3X6iGUKOCpWGfk7KgGEJDx5v1T16yxbnrZHLdEjbRBPydRS9Bt5hC4tzd27/EJO+XE3hK
MdpQTeCGRHiDqwSWZM14z/pr3Iqpz+v5lRUtGtDPzB1YQkddAKY2KyKXUMi3sxe/4AKAadCtRUmn
VWzNKX5vbdTZfOrsl5mzsPAfZ12IYIGsrJrjerRlDk/H6BwyZu10L+kWYIalp9p0TecRSzWpB2FD
sH2Cl7rruAvdtk7NZ8ybl2YvYl1awTKl6D7XkuvbuT7okrA+2Gdu578A947S4DkLRyZjK9mCISZH
zdX5V0bidOZtOd/OzfT7gcBB9Ua+C9AlpDO2bvxKxfsZhMNaaOh/oFpcSWk1ZzVIkKK6lOiphl9g
iIpvpAys4jzmBdrWfqV7ezPo1SYnt4+BlFN4T7CcQbc+hOMguVOvxloOGA4LZwe2+CpglOtA1wSR
eIhaL9Frqs9QsPn8y61gVSbpHBl7Sa880JRhumyuTa+wmZxFuQJN2vi1Key5vH9G0tswklOLhjSv
+rrl4KDWdZeLd4tFVcJvJ9AqSjGI1SBbrBBAy8Yt8XA/tTUWFM0vusoirvUbQ4Z9KDyWvADI628r
EwhUK17t++G5DsoN2aQ1wwT12oEtc3JJyEI1csyI7eO+epp7shclaxxVlSeMZrPT1Uc6DZ27YRs1
/7z0yeMZVkCZo1PBh/bcvRVrAlT1ZsStHNl/4E+rTeifKT44yBS9FH5x0LNbngrmhqFU23LOh+/O
DkVMdLfDgISzbzhnpuJKaHMc1MtRqYh9yH6TLnBA5lO3Hv2YIbkulFosHGTqBBrwAtxwQn3F1Em7
Oyj8djlw4asYiP5WgRYavvufsLlsQXIqqV+8RYWRzVRKTA/YSea4C0OzHiLu8h0W7QAP1ToBDY1V
xPYyQ8v4JL9rZPWPNc4FMElVmma2b2VReqPJ2bMk3HvhLgVWTHGDT5IGHpad4laEUz25n44j6V0z
W1G+84JBfjxpNVvv+67f7qzmraIoRtTOEBToWgww8Iim7ZInXIydOeZQvpoTql7y967zikRo08RU
CBsl4t4YDpO+ZwXPSRaHlt/Hqat8iR5M8fP5p765xtCD0pd9Owr/hpU8ct4PQryGlpzew3oZZhTd
uSkTKljb+4Ig+FCcxm2m1oX0c0DluJVWIgJCC79ubVC50v8/PmrmarZpxvTOoMHLg68LMOC5GlPe
GMDFtWwSj/NtKg0v8lk5/7Rde3UqrHY1NAZ8i59U/kNnGpTmCBHn0VFz+WFmtVODomA9/f0SZ8WK
rmYNovu1aZNr8VFnpSJzUGwwSJMEYhdYz3UY/yEjA1hq4Dj1GB+DfplGNOob3mKLaLzSc1ayAJA5
qtql8nUSXdTVvDLf+tydIt6WY6iEuvo5BtXjLfPcF1zfh+036ee6t+t8lO1BsqfQJoVODQXpwfzY
eH+E4MZCi2IPXYrHOgPygWm7/Vj/QGlVWsCdK6HheYJtVZoFKAk+G2fTac0sw4WkhgnA7hwtbvYY
gWqRBhBPGnPmo6CafAyid6ykjWOEuHD18w3PQBcPc+h38rRyLUrNaE4J8p8AxNB9b13HJ/0+SunH
Wew4lIOhX4ovYhDnONsMhwrnjNm7cVgVnxa60LjuvGcxt/3iZLT9Z9dohoHfXTPXA5taLkOF9yo5
dqv9yfJgdOWfBGkK7lsgRa08LOfVRD8Xor2ezqu8wEBu38sABxcHbiSATVMXHn9dC6SK5a6ZTYAQ
Bc/XVNaSBXToumQeBU/rMjYP8Eu6LXnFWMwtwsMfYFS90KgKzz1CPObIH3HeFQnUtHKZSEurULj1
f39Fq7khvx4r/mnAk12hZAEchQCKzOeiAHcFTAZPYDXwotA4GIhdEFgGTdRFgiSe3XcRKvfNhHe5
rcRX36exSmOube4RM0+g1IocyBdU7QzSUtAagQtw92ouogLsI9cAorNHbwlCvEm62j4XmB/USwHT
D/95QV+gkuKZHCWyCqM5waq8Dk8sPggiqNbjhOqo3JR3K69IIIgpkAoVJyB7jw9kWdK8Tl+poXy7
njwZqiGrH5kUDxKM9xJFGX+vuvF6ay97Y8Qo1ApRWOxgfy7UXeKzojPXZmgOLBWqMnJtcaGe0oL9
YmjcVhijr/6Q+qOdV5FrVVUjZkvbfrdIGFkm/ScqxnyJxDTaE4ueKUX3fpL7J/bEfyi7f6DEEhFZ
ilP73JAEvTbYESgB8TNGid7j+a1pBS3tpK/Z+3++XifL6oVqcok0qbiDMo0hEB9EtXGD2ZTsBcPY
v53OH+0ZEiZ6tGb/RHuIYrS7JetZVHu49P9O6OexfUNvL/CV0nyFW67Ohap4jylwEz31X9TFcGEm
5d4WogmNTwkMvT1JKNqkkoODwUturWl3bNzYicGSVcsKpVbsX6vqJqFq/5k2zsf/ZuLzgpPStsbk
IdSqNAQkaOLVcfghKv+n8NRc2q9S/TG8XODqtFJYDA3KxVE0iT56HKB9BMOfTMoJ2UqvrejiHHOD
QjI5gyJ2v+bMt6RhTFJELs2nwYa1i6PtaBya3ZfrqDeGvSoQeJlH+OoYGnvJQZl2843hoy4ee3PX
APOxjToYGaM112w7rBNS599uO3xW+PN5Omhbys8W4bYS86pFig45Qkgp4NcqGHzCGOjQ9BG2c0fz
U+6f5FeGYtrNu6HZflf31L/fmTKbDn4T+BV1JeI5d7OGquFINja1FBOn64U0Za7lCvA7x0Zq3ovV
KFEUrNTcKo4OvuK/jxrCHipDjcYXIHy9k8wUIf4QgdMaA2PpdYUF8iayPoPGFNeEmvlk/OhzeCA6
mQBHTS2PwMRS2/5Vb5BJqaEVSElytTiXZx7JMMoeJFYu4o2JHAYy7bA4MjP85ouV4cWHBVx+l6Of
CO9fhtHzmLbfiJwej+y7/DenNxSJAekdcjWU9AI+766zZ9QRHzanslisva7/+no9Vi5imlZizhBg
ZJyOvD39/x5Z6ALQp7I563g5XSgScIMNJVd5d8hu5uxlheIEGcRIZU3qmTxZ/rNgaobXsbpbYzXO
ZCpwaPnMp7n0AfcijZb47P4cXhuQ9Qok1PB1rUy9v7+IowOSUhiPyn9mAxnhqJF79HVm1IWvJuXL
DJEKfHkaPogWUtBhAOWPmfcjoQSJGHyMDZbdAM6MtMGj4K3NoEbEYze3dtHnAHqGCvFFtu39y/T5
s4F5IsbLAUZeuXk10Kun3a9MboTtjJJ5u2ZPMy4AJ2HP9kPJtsM3SPDZZ8iEovt/OgboXT8bOGEx
9HHaRVZOKxa19oJkyyTC1TdOHFSCoH6L3WkKPazYj1s32xME+2/jK0ROSNU/yPRijG9cTuxoNXRD
R+V97vP4W9PIyZioSWJMGlQwxN/CZK5ove0/2sMfRUF1DqBi5RhLRVLH1M33LrFLsDo0iim/5Xm5
svf3DGhIQs9W1OMPnFDq4brL53HYEcxge7R31f4YpX5KBiitjyormPjajCWnAKpkCHhGNg1f3FEw
bWhaBKpJtmrWCXEVyd3Xtlk3KKj7m8NP2TtvbYELMcJPBINVfEGOyrQ1B9erEKnmVdJiTk8h5VpX
xinkfHN7ltLAgpbL+P0yJxWXLXuLKbxmXhGkvy+4PBF4F0ckPeS/9RKzW6ejT/4uft/5hvFfoP/f
QU2isMe8WkqH+vDspLlOssanjwljLIOikvMH/J0P4206teDnUOd3CEFil8uVqvs8uPb89Gpb7ZL9
n3RlPHTU2C8s2nA7g4WMLACpKhfiH3xcW3u1u4FlgvWCvaqV3dGeajvlBuNt2pIO9p3606wvw4se
oA4OoJ4Ok9kudSygLolWMvWgbZA87WRmQ/VxEyEJL4yiVw13/MeJjIn/kP1AoHo5GH9tNjVRwPXn
IOxFYN2Aiue0ysXwS4io86r2m+fH5ri9+jJNAiOXA+2xyIg1HKSrRUzw4IndnNDoj1eNZ5q+a2Vm
b8TwiBbtQCARD/w/JUHJx/ehYeMtjlRwwn4LqEXISfFNTLiNQ+Or7WIigTY5g1iRerIyNKu1P2Bt
F4cAzN6WQab/iCQHWfUKlhz13ydMs1LRkI8G1Miua1UJ9g9ClLT4sraK+2IlzjtCYcJ/FrGfMM0g
GYm3bJo4Y8F0FCSVa9p7nRAapogLiJwYCAE6HjEE1HjhDGhV+rEv88XAafc/eoXYXfPxTqAC2kmU
6t/M1yz8GtFFxjcFDj+QXovKojiASdXHF4b0JIiwBmDt3fNQRv45s0GTINvaSu/f1ajVx7cEpkFg
D3RptaEb/r1ieSjzzytayKuuF0jSYchdFKeZMuvQmRkMFt5/YCcRQABmzLpLqxFm8pJrcFxqN9Mo
iXG/oFQaBnmAip5azNvFNCKJ80ovmbwUWvdZSx4r6D9exeA1WTjb1vyGygwn1dHYxCKkKYdouv47
h5kQpNP0pVMKqV8vnJax0INCGent/TOdcdyNv4N5oM6LwLkSnsWsIp00gK+Zk3QluKTXoI8PGTrK
z0ITfleIImd1AZ5XLCcchX9LDSLDhyzg7AtuYzN5KEupq+GvN8MDCFa8fnG9th0lWxpRIISNE5Ap
BDRQKcgh1RBelXLArRcQBlmHoDcWMOLgGngK7yqZ5aiSMFHD746pxuV+cJ2qrSutVjTsi2MOO40L
Z8d7lWVbKHhyKFJvT/9HBP0E1ZoDS/YJ/JVEU2yWi7z8RV6UqoUMOfNawJy6i30z6cynntNQk7CS
530E0Z6Oi6IhAlzpesGpPEIj3sZnNzaYHX7UaVHuknlv1s7TxPASuKC+G9MQorZ16a3mIpPqv+o3
k3xhcE3isaKZ8ziZaLyGxaUExlNlPEKYKFb5fjV1n2VYzJZr/jsCmZhc6IjN1JZ0MzLurnAvQPk+
Li2CcTtqoLThreYq6isrHvcIiqBZ36DcNhN8zdCiDR85KkQpkGaLD8/0BRgjGkLOb/wTiTxAJ/TU
wUo5qgExQL58Jtzv4nMHWoL5ZM7IwWdFG62lqin40WSiC3b5oVaKOoOPIeLNt2I//02JGbTx3pWF
6RVDudWIIvkrJREVjEf5Kr/P+bHPbvgkpIePqTBD14rhcJvjpi6fumzZ9/rIgICRlhFU/ljAZEY8
wGqPqbifFTE9l7hqJUCdggiHyyMYKzMGZ/leFcvV7jgnf1FXZj4mkLHjc/1M4kDNdGlC0bm+vEBe
KvoL3LTpvWAVOpfvY7aMZBw1A3AVRMY4QlZOERpYy2z/vF4V/Fq93IGdEsbRSsuqBpENV3y/uNCw
mr57np7i5T3c7N6DueOiXKIAjSWD+gRWRH9qfu63r3dEElpRp6ACijXWVebNjYNqmuD2e8MSDAQE
k4rg16PXI3YFA3h6lwpTy6VfHDZztteUf5GltL7Ck6aY9g++KfjRFvb8SoZoSswrPrBWC74CXQ33
yaHVDyOTNUpspu6mwgFODtGA9xihP+wR5l2ItfgvrGCGXR7S4UlNEGTnALaZ9qkKZ57Xdo5cB1Et
jMkIfUNqrHTxdM0zDxv7aOCeZuMuJDFyd9W2JNN+iRkdQKyfJKXXTGjbw1KSMzvDFUSFM9e7ROOl
sZgbzaXgyrlEb3Omlv+kzhA6qtewcM5qd8QUeDCGFcVno5MMovc35ZQ0oDq0Xhz6Eqxp0SELlk+h
h5LMrCulWP0TwDWo80kLKSXLIOCq881BL2f7X2/uZ3pZctY2mEHhqozkRqCmcuYk8mY6MozSdkce
MRc4NEU94PohJlL6m5FkiSToxwYdCNh0wK31OdcjbGEsBFCKDSgE33MOrOqbGO+6NmOqCnJ0TYMN
F2FXXocJtu12VPZRhaE2SXZXyL7nvUUZh8BbFtHXcAqTGaRi+Wq72xYWcpAcOC7HxGM11IPg8kl1
Bdmu2poTCZgxlJbMWpwM4Icrl+Cx0e6h6kduQ5xVg7XtZsumFoaramN9chf+/QXx3eXz0xx9HqJm
vMKW3ucM1qTHP9v8LFzpE+b3dJ53mSh/eyh14WYfqwwJ1R+KiluZCL+WgDPErswGJlr0HeTRkXy4
Dc3ZpzcA88u8yw6lb5eEW3B0ius4A1RLu4EZWYLnirp3QAB0D6xV2aPSPeGNVYI1JtjMbFmW8gcz
T3vyeNjP7kWmVhCgi4D+z3CnWtOxg89lce1IGJPmVfvOgi1ssxVWYPTiclHUcYtuqw5yvIm/lasl
NZNtc/7Pkmj9wbVRT2yQWjINEjg581FNczB7WS5gtFF2HVkNj6gxuk77S3XT3eoVRD+hEZxAJcRF
ivevH21gkcB88qK1b1tn7WmAWb7RtWQ7eiwxRyivc3V3K1lzSikbqvyDL/Qq0hze3RBRZ9ESNwAI
TEUJYIBq6P/FWb7Shi5uCpGE/KE3PRUfdoqAAso+RQAXHMp3k7hSvWUevpEDEC92GXtdTc+Tp1J8
xSxuHFR849++8Cn6zkNRIh+chatXff7rhhgRth++Sz7GzLA4ATGHRRy0xQG3MKB0PMLskWRRAXuM
tq7zvNa2XcJwk1JWkF64mcOsg4qa+V0Y0H2+5acdbAVcdKknA7BQQdLZri7HJFinsdwiv3uhcD2+
TtFEaBFxU12yAnZkcPnuQtAAQlAhF6NucXmn5jqXcYLKgXNZelkdu8qvk/QadNqgdXT6RXJFSY7s
8SJmZwLIuu5AzfGeh88yQpE/Z1kw3qRB/NN79g/470+rpNgN8j7nAKIRmrh6jyKbRM3s/ZwuKkdL
0HVLBIdmRtrNtyVaaDVvnzShrpPvK5yc7eAEAoroF3wt8DbT/EmeMb6EsXFawM2MDa+7aJEC2W03
+f+zq5u9woVLL2z49jd705Irx/T8otI+R1t7/zqgMyArsENBhWkA2DJPJS0GixkQrGKhzT1TQDgo
+JC1NtMNTzq/dxSf22Q3jCHBP1DiqqdwlNQH5CIAti386K/5BDURAWKs1Im0YhvRrs9DeDXRkBA3
Slhdg9NPSIlJ12rchgU8BLartGpw4e5dwQT3y+iqSh0L1rmkynCbGmOM2iCL/2GtuJBP1xDu8D+u
TvKxp4cFjphsCMXlD98j0e7+eNgLDYlMItzSy6TguAlMqfe1Is5/5y/PcOFWiG0k/lmwjCU5Jt3q
yE3rVZSnv462ZupnNa0PI2rm1aiULjr/vLEVkzXBkbmFtqvyZCezEehsMwYy59kYxPu2d7pZt/KP
3rqHLR4PUod6RFUia6I+AJe3SscGyxWWPHTpbktzmfHqcW0pdk8l4tRk8oUT7IldVnA2MxzajbTX
+VV3+FgtCbr4nEG7lf4eyQE0v8nOWJ9m0D3Hd6/qBqTpyuNl9KVzx7k1bhjj/vz6QT9cVIuPVl/N
LA5XmZHGHImBBMOKbC/dwMo1I774J2fO0H4mZBAC6tjBWDIuuNO/PaqbzVkd6y1tezlmTVd92O1+
Emj/SQm7yhNuYcXjvQUJJM92PeXntJ3fgcyuZ1WjVKW+csy5hy8gkIYVc4LifXG1A/bcKTbkWeS5
4tKaVJiJDBssb8lj30Ed8xAYOauuiMo99e8RFXJLgA1lKmMaiDZhg1HhN1Ol1smkIAouc4xT4EYV
GSTPfNEi8wwu3ig+mJGQ6umLHgN2l5Zg+Ic2wktkvuu1fZAL5p2tgdxqKwIQAhUcauocUMvSPb8P
lnOtOZWzvnR5LOX4d2rfR5oTUxOsWt4J1Ak/XEGPQMDci5AJ9TRfFzTB+QMY4gsw5ZgXCxj0fwNx
yHYme0ph7kEDrosqdap0W35oSMGlvAoNdSA5WmjANON1YxdWihyiZTrwmVfb2UzJTiCn9HwgjmTT
8YAvqmoTcuyk20tp8rtp7q3tFcTjYfR15OrYGrK7CQVLoSP3nLTYQOTftyZL+EvbB1/XTI7LfDNF
PHGvfVrbsPjMQmPNoCb1LucIL1w2K/K+ERcAHY1kIsWUvL4mrXeQyp4iYH3UNzggvv0lzUyjVRZ5
5Px9cHvyCkWaSccJ614vxCzCp7n7QVkPF/AS3+o2+uMJ3bCW3wNApowZPHRDtFTQXz3Y/QDg/mGx
5w9mSm7htmy3Y75ry9BaAYcNYcuf5KJPn39Zo28NzgKm1v+M6sKguQAf9Ktae4g5Hv1MOTnKcslG
+38u/f84Y9WIiE4OQ05TOdKBG31GdWsy3ssQV1ALWW1eZH3+vptNuw6OvjbBc4WxYITRuJS2cwjG
2VIVPAK6i0XPvJvkRB64RZ4dJ3rdgwuh81GLbTCBhEFkAQXaqxVZQ6eCvrOrOnMH/h1aF1FTExEg
59KWRti3K+msic2lJaFEbO93Yu5XWsoZgWsJEp3roJAjLlQpJHvDf7/zFZY9STeFjc/PelFNqFug
yTzx93i4i0cfuKlXFNhrwAugr0QcysAGewCkOmftDN/E9yzWwFPipLJi1eIB7dFAyfiQkGCCcDUY
9SGPm6fMYfc5Ij9Jjyo0wT3iPxsi2KkliV9zPT5mmKThZg22IvDRfgWyMbHM/FG4GbCp25fbnN9z
q7VC19KJaN49BpSMJHuhFI6ziLf+HrS95J6oC4bq4U2AsPO1HPGFMiHPBkrlmZOVGn2PKEa+/PU6
cuK8s0EEXUigEOrfrQtBVy+0IdPuhXDItspG5W+xaLe6B5ndp1K/bt2egYXnDdMYPDxsWH0Za6rM
o0L5/GW4NAUGKeQnUEsQCRRoqC77mtzmQlOsNxICCLG/lH6ZcT2hgY8gTUonQ9WcMmkgLwU0uHcA
gPTy8FNK7zFfc7cEYrbGSGabQPpc/YnxYqvuARdnw95oOtoX6vkFA7sid8klXNwvRc9Ehn05sFPf
icDmGB7rO1+iX0UYv5IqwaA4/Z/jRAnko0ZBXzu+CYgkrb8oX8oDx2hXPEww+Dvntrd9qE7yAtxi
5F7ADSMc/V3ZzyyzE0Or3JPNnnhHYMTVz2WcaXkGmE22ShplXPCYfrt1XoO0OLs1Xz+TU/GTF7In
QAROEsNlPztYBx6ksA2KsVsALcwTU34ablnePN3T6nZvlq7p2eesPIHCpsjIkmwq0QpvFUBUX8cL
2oE/K1eDwtMyBcud9Pq7kI35Z0h4QQUMKCZQHWrycoC0EYw5cRPLN08H49RMeM+0uk510YLR7Wqi
Gupx2XFKrNlYOpNc5ukDq3fdHqLuu4mHUdoMlxxilthBSAQbyWQJvPQU0khEWsRgHEXWKAWKJok5
55ov2uo4GBu5pzEN8WnNmw/Q+d2YPNsVpMKMlpSStThC2ZePtLw0L/MMu9INlPfLt4ONcVE7fODm
mpLwr+g6+FRKcO8gb3z09LqFQwG0BTkOnXTye2kePB1H3vkW5kk26nXJ7vYA0i6t/C8QDPubTRdH
H4Ci5ODmZzJwKthwbulSJXdYUSv6WXesSw0tUGL57ifQe5/NTBbzRDeMxyH2e6ZO7YMAgB+iexTi
wZ9/JMgUh2wwSCSIlQrQD5xKh6VLTbgk+ygVfibkelE77wWCtWu64I9+gj609YKG1qTgscP9aObG
53dbq87a1sJMLrPEGyLjjWPi3SgUPZgb8qq0/SLcE9hwHCbCJuByyY4drNFxzPTqnjdIFkIxB5T0
amAe78Nhd+OPHnJVUHYhah9YugGtu73OcPGH+2TmWa5bYgzePOLjLrf8dSgp83HyGXYEpD1Y+RT9
2zf0mXDMl1sFQT7e+k68wRJqMfu8J6ge1hcggiJv53eNWgM+SnXW2G6UCjrsFR/liXIk9aIDBa3Z
uUkqLGIr1VLl1noF9IrIygjc4nxvo1txgn/f+KyJqNECQy6rnUSnj7sFksnDRpQGbBySYbVYmcDL
hSpxqYVrqGQbNKm/c0A3pzE5znS7dAbsSsF56xgeGsqC9y0AEAYcPa19HrKJ58tOFJDniqvxEaQz
Hi4kUpodaxpLkLZRRUsNxig4kj1H17fYCa+8JLYsI1d71kDuFVtE5f1N26vLqGyt8Sz/SHo363dH
gBQwsmWFcYHaDiVtK1awLHKnr4DOUPz9q9xbXFIKobindkCR5UGtzhU/mYN/BZmdAogfdXGDLThP
aYaY55PSZvqHW2SAbo83Lny23+sOsYpoZeaZBIbCw2QL6xyme5QCyos5XRG/LTQPzplQXWQXgTyK
N4fXDXTBInl8vo03t+KsTmb2w+M0SKDAOETP4ImCHDw+KxwztiHYJmMdn9yPo0Dr4kEpxRs8Mmmk
w+my+n6OyNTG9yLiSSAeYvDVAVhieC3f8I9oX3isXO5+psnuXT++wk1E1Uv2E1E1+jv+YH9XodZ4
ftclYuQ+uiQxJbrkiJ1mdIvPN0yHnvSUnkEoqps5REw6fQFUiLia/v2yeNMWBKsYNe7hZ7tWwQn7
dP+8+QBll+cdkv/psNOvaN7KiSmARF/CR+eCLOdScR1xuFSZX5qy1g5/e7v7kTQbgoCZGnaWZ88E
lGJksXBNk7aY4oXXGpNgwFVwIhaCNz8/AMCe0d6Cvh8729S/smhUJgfnVBmMumldRKMUtzEgN9Zb
UvUfyWQz1VR+Zya7kSeHNDWyV1rcspljsETZDXdMsUrieQaw/9qjLuXhnFnM7utvgk6iHOJxXuNj
RMhjLlK8lWxQfwujlBkKrZh9zvNauoMoht/CFJkxxJSoH4bJwTwjvwCHJibeTR7lRLWI7SnT6j+5
dfgIzKusVYn5NmSBClByvd7tTsaVPIu8M42kIzE4+daQSfZNcFGYI5ecpKss8fW66tLix3JXt2PW
CJ9fuRMVQHOCVsXcmi4r50axUut29YM4EZNu9bchgLPiu2yi3096IdchP9YYW+odCeUSUH44xaax
BQJqgm0tLG819sk25sGB8jHvEjzIyNY8kTsaQfTL2jP6UWW1e3rIzAIpdM7kjRhW9BZnTQ1ApaVI
E3qO9/MQYPDt0Hi8pE2GKrLqHFrjKaPkZKp/KcSLk4OBgOoqxWv492K8xb+rUly3ktIOJXO7yjok
QFyeiC87UY/aCf00Cbcb1tpwGJ9YyLssfGka2r44G+7AoW5W0q8iI387U7Cl7we4ioIBZoVVIBcc
mTZcQ+H/N50XryKZ8mp9Ezd+6ef+LTEsD/sXV5LqMHykdw41EnZrl0Dfcakxv7hthVdwgS7m040+
296FFoNPfXRA8z+Tk+xHZ4wqL8PKXZIEtPA63rhO/QiS9+ipC2ueV/kclLTSxT6GPwNGozwdA0n2
OmDIY2jAlzU1sQILq820406pzE1SB8Pq6tYtZRmU/PUf13J7WIV5y52qJl+T+CbCyU0NgytYxlQw
pnqhlXMCqBNJr0Ymgs3Z+RbruBhNonQccYJWc07LHqZ+weXSWj2TsCCSLmRiFKix3ur5WQJ4YkCl
RrEEGwS/RSve0wV4kh/Km8ud7DS+mhWs/aw1wwojW8YYa63mCR5SVZnmHuDy0P1cZ4Da525fjxg6
HckQhk/JnYHkta3syUH/ZLqfvPwtmJtxLWwsJIaBFe7xLUfLHDIRcRLXpSUVF9M7WvLE48o2jyQz
SgiUmhUS2+R10HHzQTcDYKhfGCJ8AiRnoU+HdznJ5KMYxMw3rjM0AsQu/Ek3aNuHkrTJyLVPoXbw
+NJPKi/YcVAE/NYvROTTP3GVkDgPgWyOMZ6QeRzlEE/vyRZrNkpjHSqiyi8SXjK6aE+YyhSldLe3
RKXkb7RwP2bcBft07K2/Vyt7B9RM2XtNy2G5+NF0oEvojImTc7PaLYNmqwgeOg31x+XlmueOGuj+
s6YEqjK8Sq96hU48arlmPyRt5yovvlDM7AkxEn5tmDlrIffV/f+T3dXp0s8VoF757UFy35P6aFrw
xyCXenjThISJ0JO1AHKcqSpKB9CS2CuHZYIhwbvRWNtrYzGFkrnsEu6tVRXnon7YjEd0B+RwRRjk
hu4fGUraZFb5Z1opkyhMu3nFqwyKHj40O/t56e1x0Kvyh+hcvz1+16i4jTIuQry55gH8vSSrp5Xb
zZOKPlwZ1tnbTZEm8RpHMJdLQvinGNrrX9mg5qYruyN8EVxt5NyJholovhF1Sltru8zNeSQDNLIl
EBqQaHk5INJLpCgETPFa/CvplUBZ5f4i4uhLUvZzpYM648I+QNGsIAtQ4jyTJIA0/iUpj0RWtyHy
Xac0JKwGxQtw4dgItGIfvNbKHLBKIfj9vas2eU96dQhdPDs+WNqXvRRMwmjAa8cIGWFk/+9VyTD5
oHj3gaBZdPUtPPD2/iHa2FPBL5snctTVvJoAn4Y5osaTmsYZfBTdLgLIOtXMFLdXVvYeJEi+lfTL
BxyV0hGDOZS4wx37dX5fCW45Fml7vtBoC88HTd3glsXVi5EdWtEnIA4GhlAAHf1oY0kuFK+V8CgX
4BJ1rW3U9LvXzcSa3/9y4Wu6YdHQgowsYf1VqEt16xg+L8NdN2VfgH3BWP5zotpFarm+eVtCvXVK
NUHStYzdFSUktUU3U5Pka+dXQW7m6Q98BMb5qVojxYgdOFogaS7LgYmAjAkdxDImmkfqh0GIpSbp
D0+VUl5CiwRtNR6Il3bcuI8qAPW4Xj12/7CGtwuNyrH52t2EA/V37SXTUkyWqQm8vU0ZPZCH49VF
KirdAZgtP5SEWAxKbAPZIUTBmWEiVWXoheJilzZYS2EPDka+rzPVLvv50kMPDD4WiT1JS/wR9Yk3
Et9nYA7VFORdFjLW8GpLPpVpPQzUa0ruutX+MXRXV4OM8aSFlcqyKLoCrtBf1oQIMP3tawz0n7iU
u1I1jlrLr6GLsl+x1U5f/PUVgAbRzQ+C47Q9kJe/RCPbFZlYR58AuXcVXNnQIqxfjuk6uUITmIu/
YpMwxYl8m+NznB8lKN3aG1aPGS87TC1H8gdOpr6Fvg+XDQeYMjwB/enpn4+A+ogGTMXMTcavZTgY
bQAPt8I8DKGM+93K/2TGWXa9go14STqv50sQU1T5wgAsA3MgzSlQsovuFbfZaeMawY0XBGgPGdMt
spoRzgxdouQgViFa+Ii0cXEv+GTTWz50CS4suGZzRqHkXs0E3ifP7ljPGL9MiSZdC7FZz9N+QpBG
JhAPCmJN3LAidQmiuCikk0JdIC4rUEDnkXEmXSAi4b/0RFwjuYo9JLw4EzX4WsUdhpxo42taT7sv
gJ8n//Rv9Y7ChCY2EpCf/BVFU1bQCAkyNGDE6bUAGcv7I2JgD5N61al3Rfkjraqm5+G5EfRpjubk
6XeF/OS2QKC9HT9pfEXyPYZGGWsI860U1FRryQADfZj6TF5S4QceH0zyzgLUfj7L+3Ob6juncLX7
FNMjXX6siHu7jK95w29b94e0rRScvVZEFZa2hlf9qj1CCKgt/kI9fCQEf/SbMfA93EInRDQgQQDm
M0rrLscSxCDBItYO+FvUpgOjrdVCM8rTMGQrlX17/omN5ltmtFgTy6Gk24NMrj0rNPCPKN4+ICjF
rfnq6i6vtqBoTEQ/Kbr04fzUrtn5op/oDFsLa+OldlPLpxVIlzuzC8xIQ0yxZx9kVsJv90b9+BT1
RTPAJ8oYr3WvsD7BfXOwJAF8wE+0BUjnRIFXp1DJJZflonGvcEXktjvIUv7GeX7nVrE4R9wiSxRx
laFGV+cXsS69sg3A5Oi8fB5Mp4MGHD/qmNYuHfL2R7/R4Vufk002l+CV9uowukzlycniCz6nQq28
gHKq/TizXW4xNuIztiumGC7rofYx40rqn2a3yKNNUiEecotDy5d8Q9KcB6eB8joJRNRDw71bAaNT
N2BALHBnCP9Fl2YBPj1S+eoAHSFUqVyjQfmKqax0amk7JgZvy4QCp+dcpGGxwenf2IPp4Ahm0qer
j1X8tAXOFGiOKdx/fYEb02wNI/0NmupfdW4hQJW4HFDvaeb2/h3w8NNhsu35WSqcvMyeJ+iA2ClH
EcR3cW4gh+892JREkM5+Yaa4ddF8yjy7u2A4MFqfwmUm6ZYVVgv5X1fRfOMxULICgqeoT7nssj0G
Ejo6AZ9s2Rzz607eiWZa10EjmoiyAn6OqaXjTo75sfKKl20pvtwYmpceqYNXRrb4W/yFwAVz0mTu
eBC3i1MWrx3hF0jIvsfJKZz+aRZpHUJ5Vy4SOSZksJdmIS2Lw79HQAFY0NHYMnGNL1JTxnDyAQ4k
ThQnOIxFgkO1esdsi2ypW5dtWd54CGlZ6GZCHwdEF1KYhfcWe5+6C6F/0EG/MSJ2fOihhKdiFXIS
KzMTNQTtMKbaZln83p4v0Xr9F9AwklEAMkU+Z7Vv5W1BSAIoB3hukMLRWjXaeViA+mO+bP8gO5xR
dh1Iwt9rvmCLtRNWfxA/sH6XH4tIxDU7qxccMPIXLHF/jntFP0K2ap8cFZShUhsK6Sg48Y1mVWgj
dM//MBCbNDiGyccyEX0bMlBW635pEwYoOKF+muvN4CNJQdR+8znqLwHuIHrO1XvFccQ9g0Vyc1js
K4Sp1J8mZHDLk+tTnFhaA8kVuUOGxaYHKSktfjRLRxTW2QX7f2pUQMBgXpdIgM9yqqJqQF9vcQhy
upC+z0ZYVwGX5c7Wyzsv4tLxU47Mvrn6Q/LZmSNmclI+wVnK21wwC0Fm9LT7KMguqi9Xsly31aZ2
84J4f1HJJTfqWPkbwODc/mTJJWdZkKmM+yFUNDQaDk5vmgg2Lpmj+k3/hxaEEXFzsMzcwWIeO/ef
JReUVLi49BvsJvc0EqqzMExAShMHbqGW11msfZuJx3k8QlOT8LuFL9wQfvJyDNPzJ9vhSmbChjIv
TANilum5ND1kaOMFOhKfG532eIkKFmwzgTXivqtusPIOscXDxF3l8PKD26rVW3KPGztZo4PZI200
Dh/9g+65l3PlCnC0fXWrs31jb8YXET09zXXr6HPWPS0Pck2h7TTY3GXauf1e0NirymARBdcNUWnJ
bUW01L6tIEdrYG3Umxpi2S/aFaaT3qZ6Osj9PGYsV4z2HczTo/bPeGZ4CFoqSpLyIclmNMkEDDmd
OBgKv+PCNrommmVP7ejXfOx8Nhibsh57h74wzu21YFfeYcCnsPOfRS+K/Xz/8sWMQ43l/lon/3BF
FplIF+7F0LnItCPpEFbHtVNMlevQ/kckPPrLtpXv6n/hAl6aK/cXTQisGJTmREZV2iw3M475sWuV
pYq1l5Ykw/MdjnSFZNF3MMuiR0s4a03VhUXI0att8FbeElS9hC13dq9rBXwz3JRAqh5bKMj+I1M4
cC0l4ynPti8dYPmFIUzKTU5ExzS6uhFbuhYUKTY2ra9O0+RY8q0ojyZmJDyE97vVtVHy+xPsHV0I
cij92VRt2X+HrNz6/6Wco+2jF92Tfpig/gJwoDqMvQoGi5EqmvGt9Gf6Y2FR2jlO7QBr1KjYvNkd
613+B76hk85wmOncAPlrQlZWu8UCcmv+LXTNZUcKqNXoL6vJUG/R+3QTABFLxGshsTqwQKwzVhCz
7yz5jmOlrvThhxfYr7FkcwBCpFdGmWSW9WbXelvXQkdWDGtYGJrodkSthqoyL0ne7anumtnnoaei
NbwcWhU/3VxAAuqgpmObaxbw91WId2uqYOEJUVh6DPrnnVveleieC1rnbBFzAa6EYi+jA2U82HBA
DVv2fVuerRJCsl2jsd6oqsWYRvDLmUVc+SjwNrbDvZJKQWQkCTTlj1Tr7TdZfCoBE2Y2ZXbOgNc+
g3Dyl0Ls45erBJf29I3dxAl+T4pg5qrb1TisW4dTnp9zK2aUPlxmcd/jhSZAeWttE/9jEoO1HGXs
HDc5chJBCdoZqL9PgKFDI7Yc2mBQRzKtKdlS2B0EaQ8r7x1nlekYHCLMq3mdEGb0/hZ/O/ToPmvU
Rrcd0p1L9bTgcPPzXSwY2bliNwjGmjIvjC6JYJRvCExkqnLZCmRpqoa0w+Vv9jxO3+kGg0KB3+Dm
aIrDVzp6t5O6/iq0SYwcpl4IvLDnpM9o1YBfjhztoLNMAD+9N815ckFHZ5nmNW1pN1IAG56Srfeq
3GeK0o8Yz+QuCSWx27/BpnLLxHEnp9SA+YUB0THWoGK0OLTpfnRK+0nenaK6wc84MNg2X0KTWnYQ
6WIpGBFP92DKyhNXkxlofcyFZgdhMGWo8gXVS4dPM2ZvdxanHeZHuwI51JN/JiGWNzpaHH16Nbls
VpNM8R77oeiVu09VYnIlO8rm4H8ALmYWBj8S+Rao+asfLy+9vU2RWbep6Vcjq+4uIemPxjg4Fm//
cK4/oRQxYIWasljgl7jgv1ebUuHdmUGMVE+RDlu9RjiGRDVOiscwv4faWSzgWnp76mBAlzdRhXKf
gZ/NovDqs6r9gfBGsIxf7X5c2eYMMKt2Ke4ePpWSTXj68FAmLj/WUre8RwVQHdS/VunXhf6yQBne
lMjBZ9Q05oRw75YouUeocPP7dErd7h+uhdn4bfhjY09BfyLihZlthMN6L3h+1YpTKdXFv0jrJp3S
1mFM1Hv5LiCDY+afk8c6iR6PMpgU+0+/O2NtnX9qWtnkY/Fdnh8yc0PLWoVaDpWN48fWOOgIeSKk
l+qPI+MbmlpSD3Vnr6xoWr0bPBO4g+L/NgOsCJk/uTxVRmuYWNquseZFGmnwUwTDheaJvu9n3VWU
GBKwccWSXXOoUrH3YnxrzfyZAVpe7jCfJI1xiJhExpYQ+oNZAi2YOgOoNti2BazOffNVv8Ov/Cq3
7wrknkrdQHWxJUx6UFKJgv3OzL/uoYSN/0hbGzYJ55PZphIrqDUAUWI2m8hfML/kpVGpgDWrTziZ
fAJn8h7m0UL5jNhfDUk/LBI5zvDH6B0RKUa3x2DTN4FaIZASQA5/ZFbKijON/zMSOfQsPw+mBMLd
tyAKPoqZFrIdajTaDojbxbc5lCg3Gixz7V01cT6/wRXS10LTcbhw3dA5Ih7jqWlH2FUsZ/lNyY+u
PbTWx4dNE5BzgiX4V268M6l8r9XBindIt6KywjzexRUZxg82N3IOhzLR43BEoEXu+G8mAXtsgM1L
XJFNV+fhtKqtiAsl6hyrk2ffM4gY60F2u7aHNmWx2vdZokJcp/5LYohkfALbD0aO1ZxEFu9CE+57
1ZWaZF4/nQdNOULPfJ6QqOVkWyGqb5Ebmu87OYTfW/lvD+SbP+iq2OudlieSa/1iHstYPVXAcLqD
tQS+gF5hoQHJoMdj6BvFO23EIr1TqnDorm86OS4YvwYgADfcRDuUiiRAL5DhqFqBDRfsK9iO97yi
NxPcyWOrvfUV/LP1NLneEjLi0OYE5vxhHFeIfTclOpP5F4u0PrcFXzhVz1lrRh7pPoYBzS8DrkLL
s34du0jAkMf4ox4DA7wUQhng2hKA6R63bTaO4yXlFoU3taKFRKZOkx2A0vg/LfHl7ubrTZTplKbp
BacFMsHC8wai7jwQOsJR3vC1NF8a+U0o8RgyPnsANZE5v1DSCFEO4J++hhtcq5H3poA4Fo+Rn2zd
LrvJiuA7ftGgdflw3cPBburTwURvn+ROitUFNrIwX7yFQ/XQrkb0csiPAciN8U1ETIF73BD82puQ
xk/sKMkMR0PK1ReWKb4u2386XkzhYd+vg+2/hwlg0PY7Tnhx50RrgBDcHpBDwdV+wMu0SPjJBIqp
VeMBrNR4HDXq1c03gv7GrEQ6bXainjI711aaiUoY1f9vWnvu01R7XSbAsxyGXH7bQwP5PH0GMCcg
U8xpyDIk66GH82QYYzhWEPme3hx8hARHEqYp0V1yyP+pl7YanPDSfARe5P2733zAc29OjUjPqgXf
FaogjECkdB+hcK4U7hGFV/CCgsSkH5k9x1TymQx0mgtbpudDK5Nb3TySbLKj1IkT+xWWVa6dPkOm
BT0ZnsyN73ngdvcrwhw2jwEF0zxFgT51MGmQY094iobQfFKdsoVAK8kzWgGRack7sVK2Jwipc6Fd
m/6KAT2hwy4K60Pwwv2+BLk9c7FsLKfkakDK6Sm5pDNrwnhMjlZpyXRJXExkOY+cz08I35cy1o1z
0mhaWJcDLfrPmnAaBIV3OzrG/jiNaiizoESl9Dt4v7wNWCsApE2Q+ZXtx4RvTWSUWdnFnpADycAi
1o/14pm92iAIlrBh6zyuCji3e5bJxATG1Bc4Wy0r+LxufCdNcdPCSWow8cJQ8kwUo6GOMLtFD5df
0i5AGjnG+eQbYYTD959lZ2RIf3adVAp0MxHrH9mtvTP478e4CRd/2AkFFj1ZMFPUr+c72Iwjnl8A
+SwS3Gd563sdIiRwfYGpaYqqcbO1lYl+7nNiOJcrzJc0wVlndeAuf5Uukq3FU/Kvh95K8M56itgq
u8+xlvaGCi09O4G/A/rCRVc7qTUcuyigTL189E7rXPsdgtGL9ViqOMMKeoz5ojBH3ea0AoUXr8wW
m+ZzYn+Y3egDyzgN1EZc80yNKHxB7fYrPcO/NU2h1IKDQnOPtSUXHMlZltj5VCEnEpg6+m+JMQ0p
fXnkpWBo/JE2EbuuFReMglYvx4cBr6tf+qmWfjoQHItA7wv/MFTdWlB9pWsVy8zyDVnHIVIR3+17
nykucvv2Klkz1FyHpSqX9kLVR/rb1angQVvB7BhJznUUaMfxJP3ZtU/osTrNAGrOap08tLdZkYyg
Fr0jo1U7ZXlP68AFKv/gjhZMOrg1Beo4iq/8MfVPnmhtzzid2LtLY9gHUDvWP44J79lHAWqowhuk
QM52E8jt80ykU8n8KhOXdIG75hj+EAFWGmMmHYCQLqDLZZHEt9sGWU1bcgrqkSXpdBFBBcojTKZH
Lbo3ES01jw1lxA46+dNaQVMLFIs8UJNlpBGgiSiKEKV3/9HtBdqIrQSgVre5lTfA3MuIAy3Ml9Mg
J72kBlxsCtXXG5RmRIonQkL7zLg1XPazfirdnQ7cnyHNR3oeYq3KBm24g/NLGvtNbYM7IPMhYQMg
9JQLGK46blkDcl2Uuo/O0bZkhnlvjYttbAKktgOwFIGD9bbyN5tEBsmmIjqln/CdE2l3xRd3r9VX
cubPHtQdLjhqMQ3yFX4UgESEgcdTaKYtCAVvhbNYVJ71yl71AcU02+sM5tNNaKbnbiPhtwOxr+JW
ukBdVblAw9zTPrPy3rbeVQ8HNwEup+zCjlLeB4AN2YqDtm966ec4Y+B1KZITqPTdIK36xx3tYuSh
pL6OBgrKI7DYtg6TL0lnxUryx9/huZKJDDU2JHPs9fcEsy847VIcIsQBUvPyuhclyjAD9ECBgAeN
qdVbyLfE6kv/qEwEu3jeLqB877Uh2gaXCBuyEP1ZU6uT7cZBy/KTZVKgOapdkgD8wYkwDg7fgatN
dmvzdf4k59golVA87vZfFMmARk9LUc7Wis8gSRFNulqaPZqP0t32Vl0T3b6P92aZ//SSHQiQ2ef5
VjQLe5yUMV16+85fsoX8yy+d8C3chTazTgJM5U0TRlIG5lRdSvLd5DUARu/cJGpLsLoDSj2w3vQL
3aNQVoNqTVllFmwsziH4JRdvZesmFUO870rMywHc2Qi4yagkpc1l1yqinOROJKqZtbIEcZJ3kfUg
mqKy1Bua9XLLHQnxxHhCbZAT+tupQaVpV90Y6QBeklNt5DvIaVEKgq5NMo9PCD4ePLQbcAeaLLGK
0221XecqjENn943suVBIcK71HWLgJRj3rLLdbjev+76CH36FQ0VLuC7UbJV++SpEzCxtjxxc0YlB
yblCk1hGSYYKrTrjTFuU27f3pLoAT4Uw7nzAq+lI6hqlsb1Zisb1iO6YBrTa0vyeuaVPJq6z178i
MK9OQSMNUjfXN7kKr7evpgNnbXbUxT6uQLmgbf4cSO10sK/JzWKx1HaxPpUUaLl/frERDz6gHVkf
uR3TJeEIMGgZkaupnUcwRt1Q7wQPeG6u50py93SFJE90dNSkZuOHSyX27SQxSIlTTBdviWtaw3Gx
F+MDYC/EOOX/UZGOrOnbk3O8O9lY9fYPgd30fvhWJgjswykPz3qzL9z0z+K7RHr//hnZHW2flYyn
23YTL+4Qc9UR7ehxMlCfQnzXLYo4kkaPfdS0ezwyrwYzHgcT1MUdTJZ0x0pnDWs80SmS1qTzgPfS
CERrCYOgUVB8jkyc49J73VxKz7uLThZYiKR30RWCVVR3Qdz9D/M4Kw3+5+NQS4pU5lqp1GDj7xCI
bNH2+mwAWfieG1P7yUjN5WpFJ5buQybj6m3zVR7NR3erxjOiRYEF8bHiGQIjV4T1Rk6wEknRbZKK
FHdLd9N59xmDQ8rMCx/YiJFHIEBIBf7sbBZNX4vYQt8DGFiR5lqa4ZUyFfAoVkLTncBl11nlh6/9
h45BrOdi/rZmXThD5orkmp1zNPRsQaRJLQPy7a2sAujC1dA7idkp9P8tC99g8t9UBT1HYTKX5enH
807rtwXzdx7Vyc8dKjc2l0YLI1L9F+9fhTFPcZiy02D0zLoAc4FoJFZfBT3WB4voXOrWM8VCv4QM
22y6MgY1Kr1n6VxTOsso9n0q3XiG7/58psXCpHQrovddByi1UnICUrLsITEXrMeVurImBtgjRBQ7
1hph6pChe05Z5DZnsGxTF7DiEk7DcSP0cj/ITOgFxsfdx6kR3xJyp/xXeDdxz1DEuSY/tiydAbrl
0d6Af2LP2gdeIC/jTFEtUk+aagxO3C3gRtYcCma5nFxwjhitcY02ZP2MJoMA7R7b1SSt4dX6CeuN
eBy7pZWkwaQMChELEMd1els2hPLAO+u4ZG7Qv78Gxv/kRva+HIZF41HukI1CvzoI6qwbgjJO7aU9
5MbXjlmDpOLxaZNPyJM5E0avhcfLbp46uR0Tdr6ybkb8KzuwFJgLNAuaN924ztoY2Pelkk9ovDei
hQqL4RS3WR7bYP1Ma1pWA7JCAitIGdb9gktLXjyDViX3QmUJOxh1zjEXPvyBQOH9iMhI4bVQiEkW
3B1Bj2xVCDv/lw2MsAw9EU0J1jBYdyG2Py/S9aarVziDmhWTSy5o89VAq9yf/ykNOCo8YfFOPLR3
rrEobHudS1wfDKoTE2eGo0co32/zePcla+AVJZZFzS8xLKAzMXYo1HMhfxnCqcWXaqiFCIbZDBH8
iiN1/H8G/BcKJtTQk9rXX7hlxKXBaYDMcCW1TvixWzYbmek+S+chDI5kiJenO6SJC6cHvk1KH64s
kRDUPblKoQ2dlvrKU5wTYJfYJYJaIhROSnyH/dnFUn11Awbpq87NmzyqwrPy18+T0T5eyQw8l8Ma
H5XNkGxCOr42y4EqBBHp7sfT05AjfoTYR/gbndrSvXsahOhuPBAv4fWK6ts4+ej5gfkHsn1QYUO3
RMU1IdTBulomZGs/7EFNCSWOknfMTUOFEX6WDVt/i5itsdtoMK64YR9IOFAUTt6+wkIsP+rm5EUy
tmn6Y1qvKVa3hJcHtkWN9+EmL9TawEytdFza46xufAQnsIPQaMvHwmDGtN5Mq9h3YEqkNS7F0Ghj
H083iTsdkQZhy03FHFzeI+/V/vxmzlEWBCDgBRjbC9oC7unL5y/OasXjJMMeVeyuhLLF3kZJi5R4
g6ENLos8i1DIZH50oDkIavOUCjQMa/6UG3501YoHddg2P9pGL6Ydohi9UlG3R29HXVeGk4jjOkeF
dZ6WkzIempwjBu8MM/9TCMkoljk4FZl+OuzfSEz+2PFzcbM3nC/3dqihMvpf2j4QZRxdUDq9VeuX
hWheFOGxaC+eyQdgdJq9hnYN94CmnZZxE2APoHWQpvkBbXWSlQi+Ja5KyxYb/wPV93bhX4dwAuSX
wIMchIj+1z/Bc34M1DsRJ4b4bdaKN8MjVDqcd8D+JYnkITs9EdHgfwaW239zHHyyCTWx1C/AbE8n
L4DqxFW4rEOSOQxWJ5DPHe73Qlh10mAcqyCXUrBvPE5N0fHDNxh4wPnJCtQ4PeiDiXAVt9V9cybc
TNPDnPBVdpFdunBtpS/k1+ZKhazs2YdBEYQS1AYEf1a1On3hNpz78c9A0o7pk6mDLa8e2oAn4uDg
L1UnJ/imFksgDhF3sd09lSz72h3+wPDX09R4AbTMY10U6v+i5tAFRSxVdJ5vFMlLcjgFdX4fJRB6
uWlegMLhRBV+L8tfRBaQEEqy4MeDir9cNff0Ee23I3B0BkeN0hRNKeRsXz9NBRdTHivfkH7KWxlZ
spkZwC1xYFRvdV/a1SdAqD9K5YlzBuj6h8bwm93N7tVtmZDm0mplmtJbn5l1XRmdH+QHInRhvQ/Z
Y1lMWO7j93us+m2KQeAfyeRvNqeCZzKn3yIyWjdsVIZyikFI6uPx8NMW/a4i+iKDfyDlvhU3yE+r
dmFw8/ZJ6JpDm5qxiRxD8DrptXQRccnzQUcUYeJsfSd0Kxmw44eHjuz1jcOXQ879WzYC0ppYqJYg
2sqKDhzeHbKVMV/ckDKfaA4dE5aVETbR4OcPEa3ANabN36Gv5yxC5SFlpm2GOemTg7PxNLKV20XK
C9RixTTFd8yZwx2Z1OVqRJV+oNTqLjs/k8E1yYNavrd3z9MUTrzI8nMYPrj5JhSyGQrsBijmwyjv
l58g2tgpJBz0RCYKxO6luwEkkv7A6kuwbQS1qavtsDxdzOsLAcHRKtO6AsxY9KH5QR0AJ90ry8+F
7zP1FBEQWAejnRE8PBP7cvp9/qNexTL5Ej8cDPx1domnlnjcqvUbHzl+wZH2RfQEqBnfFhgam06m
aBCcO4I3kN1FCHeDApdBS5It1NK8IZ3Zzh0hHCr8H3bJq0L+RIUMWpx6t68YhD1/NHlF3Z5mFewy
/eBNNvb+AHATgSt3SHnrTVfBodWuIZ2O8Bkbm8ipkuxvAtJisDjq0hQnrzoGRT9Xu3YdFl+Wh3nC
ELoeIg3Ru/VUS74pT7LlI5oqzOWppE/VgRFQfSufNwKtWUTmMk/chvWuoRVebbNUXZcpgxpV9qPO
9mRwxGto8w2mjm8U4GtfVU94mwf2TCp3Rgq4bkwHuwCRF8f2a/LssuPTAayK7tHiHWCggL0QOKru
poXFt51yZ7aY7WVBmTvgCXbyT6kSxTGckcxYH1vO6GbEO4kV6GlEpU53WiAFGvpt2mHDkcwfr7HA
w5ebppwhDOP7bTB18dvveQ4e8XhHC2iXJpwtYO9KyCPN6wDEUIbKINhXSd0chidMzwe0FstjzCQ4
xOnVgmzF4++N2xduBdsKbvZKBuJBbHUJIlNEIJs1bX6G5RRnPIEu4WoqpBUOpmJtBNKvMLTuBC9B
Rbf8gwPpU+SqGfdAZSgYuOPtMh/8uGl/ow936vtsixD5HQoLlUxEDtI5ysIkPoeHMueZQfxGXwsP
rhLIDHg1fLfbCGPke+ghdN0WwQxiAcYY73R9RswQeo20mNaSfjvfSdP8dAKVttW5wTE1VUY4FLV1
kLsXNFFNUCkoDcnkpm13k7m0nmvl22MjoO34AOmdoDR7IOcI/wsT/NL/axQwH68wBCq0vDmj4hT7
7FugnVr5oMmgKZckrlcZW1H08+c2MPE/ugqwisFaRgDSrJss5dxPw+nwYI+IamG5HEyDZo/aW3V+
QVaOfz4kYn0IId/8l+L1ecWKpXTeFBoHpWka6qiFpykprA2RYV9Nh9WtL3LyQVBkiaHfI1Vb+EWt
MQ9kSR1A4439tJkdQyGWqPoxx/RwIYaXB6RyURrOFGhSCMkXOgYsCUP1UWTlbhuMBxROEgne5Vfy
U3k7TH1QZJ7w1aFmi/yev5rQzWHav3UYJZqppFYrs2Mw7tc9aaznKdPOxQMBHD4anYfIv+iN8uMd
9sGRp1GDb9s1p1zvJgezAy9d52XihZfmcb1pVlP5By2MihizeUBRIyaRjl1hJOopyyo9K0O1qTkZ
ztelQjyniT+PtC9sgrfXEu6FRD84DdxNI/lY6IJ0aXQ7SZ9gfAbbiSEA87rOTLvNe3CCHDHcKley
mlqnIoZPzIuf0EIH+r5D34RwcMyTDhSH29zRHpcCS4uCamMD6D0TucNNitfjgpyOWnwsE2XRcZx1
VQL+vSYwgNM5Z/6KHGOeEEUZhqkZ8uSWN6oNV5pDIzA6jICdTlP30odMJrLh+DpcwbGn4ViuG7w3
p4e6WgGPGqYqqTHUUUk0SCKRjo4o0s9uyqVoaUfmvi1cxNecDESZmroyNe+nE7BxsMzp7qMFB6WA
Jw3GnkGilmDDE993uHAas9KlIdjq4+saMVBEfCosaQ1Fz+EPZRHqhr8hAikV55+k1xEz9BY2AukT
ZzhT1F6hoPGuHAvCdKkXL+xTcJ1xaaCGSC6BwM56RGv2LH5O0eN0HhriJBxFzNj3z+MODxnNP7C6
GVHUNsrMJe3L4wd9jaZ5QolqROC0fkvxMF/WAEKpiGF1t8Pz0mKsWSE8yiMlWnfJBaeAlxLqxQSp
nNACURIU5T/tRp3iPdbSmOOSbgvFfRBoF4+be/OSKQPUXJFfj8sgd4L/i1fVmealvYHbKPjAWvsh
s1FQd05QJjIkzMCBSEr38wrZzowC920DG1bp6KZsugqxw28Eg4Ne+B1qg/3xLbYkrijzt+mHU9wr
80G3yn5CQRl8h7M9L9ZU11uBugGgJWygFGuHtxPzBIGzkAeBirL258L4ikqaQStdQAMjhkhBqf7V
GbVKWUM5CVzQ1ZjTVcuUexKfIn0ycoeGdibi3C5pSW5ela3RXKixnnnkz46aCxBE5g/IhsBQ6j3V
/SM6NgQo2wbY1/S5Lg9D7WmTk+/NYcBCnJdyYRgbJf5Yma9JAWAK6FLx4jgReJABwsCy2V0/3+Rq
JzpPdvxvwAX+9ApZiF3GDzgcA9KfizmgiX/OtL44iNv3BkYxixsf011QpcZW+K4otozpypwsk3K3
Ifn5UszWxAz8QECQcJevxYHIWRTkqak8v99hMGDe+QaIne9ccx8NSyScJaAoPggjqVuI41GDAAEJ
WVDNC1M/uKs5yM3YklIWiL4rUSDjJB/FxSkAUz8tVA8FTS2YB4OwiFyPaBQkFtRvuOv6z5zhlxXc
m1R6PtTKKkA7MfHCJxGNvYn9AzFatMpFuqs1ZaO930mMU5KlQz2EQxNwqdnlUK2x/pB+cEGgZUTa
MiGb7WaOpmvhiATjGFHdWCzNM+OGND/vo2uX/9Org3WM+YT/FA1QGXJzP0Z6TcdGeY+g+P0QwcKP
1fn7P9a6cfGggPQSP4i5Dh98+pZgLK0P4j4PyFRgNm6zsbN3YgsL2SAS8BFuiLl52CNoc/odXEhr
/NsiKk8ZfttyFYMwxK73eBcU7rc0OK8K2ha2EIFwcAmV0wJ4TJ6lAUmDLFYxYf0rzpHoNR06Wocq
5hoK3kedQZuwZwb30uDBlZ+C5bw4Qx2SKonnI0GUaFMJril7uvwNPKPd/DThr6G2ktZdxcY+3hGk
1ZAP9V+lffOl/2bMZDz0EGhutR7xvlKbp++A4PfUxocXVLwxyDzShN7WwmZVdohtbNNdrBVqPzrn
25eN65vTQP/1SfPXQscC3GT1/dHLp7lGd3H5Njxuj3te5TpGaphLykHiJd0DRZ303AVMfkQU0aSv
VYGCt920TGXtLS9KFopLlN9ePMnLPSvj4y+FwSj+l2XKFYg4CX5lN4m4ZFw1uZhyVJnKjh/y4ZCz
GZoKm7gwP77ZhQmCsmG6D+YEUZr82qUHNL0ek0b6SRrpt/A7uEG5sr7cMxZ6qvfzY+Opwfx2SnUf
5patK8m61WzGFhp/tylPoq/aZfRV6MaIYgDDWGLrr6EIHSu9wmYXgCusVUJUHsoV3rto5ghALvCP
MXOQjr7mxF7Bkp5jqcNo1bjWaKVvLU+Qefpr+pBfTTWZ+RXTuBxkZXsODh0fVQrx9Ck3fGZgJAei
dUmc0pIc4QRMa0Pc3R3Mg+JFiS40whcL43FK+e9z8PkTLBjw6hM8zDSx4lGuMvt/dBBiuJqyM5aO
R155r/ugtTnc2vpZqI1LC/3IyAqp8QAId3Yg5IE0EW+fZxl/gduaE/WKQ+6Ut257gT1sixjdYhxS
smFJO36qanYp3FcQeBd8tflvJPusg3eRtCDoJagXLwHXrolCiMX+2CL2h0WmQSjh9b5jqyGAnxlK
ipqLODeyTE1CCWsLuGySQIIDcP8AUOCrDaChpAw6AT2+Go/nG8mMfrtoCz/GGLAHm3cKLC3/4VX7
o5gtfnO4Wh9UYf5kbUKRgLGpNO/i66qmBg1lqjDjZyZh6Ip7734FS0w4nXZNYG/5IqcxfRhH+8bZ
c3SOC/93pcB0xUlO60u9t3CGzfxSp3EFeoJj/1upgMWveweyo01liV3OcVzlViWwJKMaf707cjpj
kNoYXWj/ku6JiSqHXYPSBUa7Gwg9NwJNGqqTK/nEr0yRqiPzqk2zYoHEGwxd/EAhRlCvYILFJ7rI
az3X3C8I7MDXV+vMFqL2daAtzRU1fRuy8e+52JWxPBWMYjPOFMkTKJdjjyzTJJCGM2YSazlwRAdE
UTghyCJQz0tWotDyiX15w8oZVPzoyDkIj/YWGJPTeYZjLzAZ0Ycy8t20di8Hg3Ee3ot5MzmyrcBc
trNhAj9Fx5Flk5GXwzmqXtwQMjEFipIRI1KDCQqpfgOpeMMqA3upY4VL9xeEqSjQMysbcY5ebAD3
b1wgJxBUeS6W4FHsFy1InJT5sH9NxBlPBGKWRg5Ym5QkiIJwISfrc1msPAZa/BCkjyPySP8u3Yui
bnYOpyRHFDxT/bY++iIv5c4ZKwUSShE3tnZWNnK3ofGH1dLvDBNL5NhUOTXU88sWpDIWPybWZ11l
TBI7UkIT6s0HHWuFcj4Y+/KfE3ffMRGnWif+xf1B+IhOxgRsboe/GHVfXvcMgdEw0JUsIm2AB6rj
hQuVWfcwstkDIMJtSVrbs1Ub4iKKxBtsMm7KYtSuaVkDkVWfg5u17YxITg19RqIYETL/nxbUAFBg
gopFLDbSQdKa/BTu8SNfRp9tZ6iylz8i8HPzP4O3glHSQBJMh075JYzY7I85BL/fXQzylkR6SiOf
hzHf4zAFC70SGie+tqSAnI/OGiDtL4kcW7n4gqd6Up3lqk4vlU5ZezFPvlDX5pvYupOVkjs0hFKj
JVzLZfx3wwUZnc6KwL+Anp+nVbNnzhJPQJrr0d3ulCWiCpO6VEyzP3uyG+jSWdsOCGGmQcx9x8ze
nFEXrnG7C4n2tCiBVDvWawCUDwrQ1tJ2YQMt4RNVcg+dBh09XGvAOPF0fTzSG1Jh6DONdLGuhWdc
VUbhJK+VDNz8128kzlOE9lW0loKmhFvEIgQ0heaGVfnd6PWrUUxN8uc5CM1ljSDHuUmf6jMAX8U3
B6PygJqwhm/faCK/9C79ShyJKhdMuyEa3zM7NeW48NHy5DG5qggQIgxptyl7lrU9brsv8Cu5Loxl
bGA3yHHp9VYkq6HCw6pDKjWFJWpnrGpBQsmd0FiCG6bB2jvl/U182BkheatRTwzv2QCtU617SjUS
eTmX9i3sS6PVXQkinAUxBg4+sq8h1SW5KmUGzI/m+OOHN/O+qPbwOP6nkvpXuY/yqF11xI9lAWCz
Wc1ZiK15Dg47BZk/sVr6ChCZu07fONqa55iJZZfruiFsJPLvLd7UiNmeiuyyJUK8Jw+JLTwfYLXZ
7RW4cv3Lq03OXjawI7TE9U+foU4n6uVktv1rRZo6KK88TJNUPxfd5iiNspLHMayWAtXFVkKQugBq
4fNy/VkasqvEzeQ5xfx4k08x1r3rZFdMlhddq/yFUlfIQMzxuF3W2LHrClSEMqw//Htw2erq08fX
Monhm5kfAguTATTHImYIH9x7FFyRCA6PW5sEEAGFgqsUSEu443n+ukDayNRXH3zuRiZo2hpL7WvB
ppmpNDrpxQgZ5Xbejg9OXsJ6fGTQFC1T5Ur/qGVV8q6Lsn2KBZSKXxlTFnfe0szvVH/cksOrW51j
ccEBXtmDdS99HJDYNcK7kwX8koLeIPGvHOHDtlopy+4tdKPn6x9aRGNrLwW4SawF0LkQFDrhhwf0
IjtKxZjnoBiSCwjElsnl0F0z7heXyVZ8XfMQT0bUioziOanONODnl8PscXd+PHB06ZVomeN0vepg
8SBceuYUKiinxqL4EDz/R5wSxigg6gVYIThue7k3eYQn4GflK1WPVB1eCkp0io67WzjvrAZg3r2c
mEt82SeywV46kpIF9FVhNI9CC1Rbo3c6zjk/2vUF2D0XSgwqpH0qHlmqlz5hxqCYBDn3FzI89w9u
C8edYRYvwRplNEAT0IAHZ8TCCnES2wj4xs3kI+ZuUv2Dp4Qj8CQVQqt/kjO76n/cG9ht79efOj2u
4CkG4+YUC7Oboihhq9JcsBZho6uT+mW+IGNdCUW6z3mzNf6zTfWRha5pMbpZXuUpq3c2pchBRp4G
81gTcMuzRj8ox6TjLI8ockZa8+Euys4DxXd+1Uw1oCLjArNyc2aE+bogdO4c+OwbMSBbaC2L+TKM
I/QzDJKyjyKXImr+6ZEyCvDC96neB/tWKWjLZgRuA9Hu75vnG2b7v+poFN7GVfzPZwZZLuPjGf7j
v7dEYkdO+MkHvwtWL7VtVScq86idBdgN+2EEU1vRjCUBZ+Gr+hpoF+PT34N0si2fcFwHZHt0NG/F
TwF7dpU4nmOn58LKCkT03/bAbpPmdKc9dAHbW33QoYacAr+Twzdwp/e0y3BkiOCN3Wy7ngjnrAuD
cqyGjgWvo4gt34rNhS3D/n58VHjzl9qEWhVb8KKr09r927xrDkYzo4Y3pC4eQSr6EmhsI0A87yA6
wwsi4lsFKdM/KqLaspiW/BORKOKKaKyR998cXOmcpyCb5+LM6olt4D+Rl1uG4U76t4BL3EEumrzK
SSSgEgWmG1F9gH+jGF74PzrpMBRozLTd6gsd9koaKiT2fdN5WVkgQkrq+XbZZVbU7BBAu+FiH+Nw
pzK3QqivSMl1LDt0ds/lEBCMg3RZ1FeBBhEC7/Eg2tdaqny2L/9z+Ibu2okGEQ8Rsv2baykw5b1k
YNpJHDmyHfiizLnvqs07jl2I7q7NnMpAXw10Gq5vu/BWGa8b3wl9ZpgO+Sqh8x3MY6x7X0q7LweA
ZXwW2OWiAxMePKUlR50xcqlG7RY9XzbHYinBCz0ApGALMWZuUAZQ+GAuoiE9brPgLr1IO1AagmwX
Zcut0aXawKLAn8zE6DDsxIL+vU824LxKWc7M5+LVL3efUKJUGInENdOFWPFhsAgHm8+EzjWgCT6T
Wo60c0lJPAnAyqZqgGhYWb9CoP3FWbixg12MxUeKUmvmCMu5Vf+awkQQRczBX3DtsHnqqu5+Za/T
NmK6NWMy88Ws/AYYLXDwnJH/fo36VWj08swRrZwRg0GJwdnYCstQ0Htks9QUNknR8Ri2u1Nth/vc
GiouLORRwIkHcDDeBqAx1tYxG/7cQLPc3DEtAmv2EGkf8uB2b2uqbpGi1yoldi1nTqzGqnEtYEbK
WUzDdbRB6UDzc5mpB4pCO1OwZTum/8ayu4i/5lS2JrBlk9XisDSEO0lbIs+uVHMziq1xAZx2QUPS
nkpoVshroaFraTW6C/0GcqxISikOuvRdBXP9nTIvNYuy65YM0pxlPR5Xv8bibi+i5HafmEALfIQ1
QzX0VnPu2Kpl29fbdobfzcA4Vg/ptMwjRxj332IOq19Li19LfVaWm7Ga+sQaiJwFjLO5xQpixFTJ
JLNA4KNvhMjU0DaUbOLgUMb509mr7ExCSzPreccugLB06MMdBEJWVwQJaQKLC6Ned4BMHflMMMyi
1+sXYnvYJVK/2vqCykdTiRhn9jelZNPzYZeDOfZ2VSGbWuv4rMMzpuQOZ4acaOJBtS61mj/U2W/y
J5PcNkTHJcwI+uouRflBeOWMCz7FlXTvCLGnvuxqofzIrwTPHbXZyy0Rszndwwgh7L7Tf6CyCTW2
O/K87ihOQuhkMOLVny4XOCBe1Pkm9vCkD2/81bspMltl1Mci6ud1VAGDc12A6Du1bmP/dpLIYs93
+Y6m69P994HrYHIMqMdIFYDJIfaOfDIUBVNN0EKySB0oXW0Jy5QwMZnklyr56ymvnJey53E9VyEu
q/BqQGVc+30knzDnzWEIvU66qV/rLC8hC3TCStH+5q4F2rndRMrdpPa59JycpHEy1nmqFn6CXz0g
6D3k7XPtA5TYfqnRL/n6V5hacBky5f9FM4w8w4r4sm/bwXxNNFjJI884IG0lcKTZ2dDffwfUn27V
Bc9P1EcNoLBDbivc3pdhBHOuRcja9+GUpbWsMYrv+hlGe1h5fD0a3uHIRxQiGbp+4FqvhNYHKRIg
UYrqsafTcsBxdE0sv7zrzG07fETIgCeDK8shZOKRdspuRo8MTMdwvJbLoBg3Z8qleWke0OM0xMLn
quM7kXOOjY6ERTbfA3Aw/BmbQpVeO1rnwJ+bqQddAUMJ8A9evEkixBOlQ4d7Qgc4ITVrNqVbZ7KX
wbTrncPRAObT1V2CSMl0qJv4wSu0nReZRv8Gnoyx52mFo4IxCBz085Jhpt5xnE9KPzKzMMN6yChD
27S7YjD4Be/tcgDEf/a3DhCZpdGhf9NUN9UZJAwbFTCkAa4oHRCYyQoVEv6K3jQrrZCAYGa9mlVi
2HrlxiNlEuKZCWz5ZwInc7/h8mbRvlghYmKbYmLzM7BhjKNYgJrn87mwSnNetfg+B579UX9UkcZ5
ofvodiU446JKMP/Bd0WK8grl8D4SO4RZlvbUS8Q8Y52aFfZhS0cuHcDtBcWNjoXUzttPiEgfHp8q
YGrzanqAmLLkSySmo1zAhdyzrFiGvNd2Xos5XVByPaFjtjdRhcZNKYCoLqBnvot86dzUihAFu1Ki
Cvfo2V7YU2U9Qw8bFkgNbJ51UyfSnJww1fwdS0splAxyiDBFG2BV9G3D855vpfGIXVNFA2rz+58F
AIGxKO0nskjKkvyNXVMIGB0HTBTkv/atUzrkYlP2R0Frbzv8jSnrttdSsnXmcOa9xkMI/0a0O2xI
xm8gVmouA+NqDDV6kAYL/uPwqW2S3nnbZ3dJMFtLl3wJdmrSaC9W9LrJMFY2OGbFtSjkN0JfIz9j
YmVd9GW8y/Q5D89MnlCZROSo6BdQ/uO3y18wJ1MBkcymj5LXR+reefQqc8k4zopFIYg1BmV843l9
7HoQos71kX/3wPyK5pkf2NKKCidBk2tDS3SEdrRk4+kFJFCvDO3VgHlVIYuS6FY6BkCxMZwlFf0x
6kOBHGBoJmn6pqqyU8b7D9CuJB5QqZgQ9ETLJ/0mdScR/pBYOCa4rcoXlZIHQHYePm8g9HS7nZPw
26B3j4c3WhekFIuCq4OwmRjMbhE1VXm3BjAUQTg5nvPL12nfYMLlMfzWfwnk2jDAXolqveoZ+0vU
wQ5G3kfNyMImQU56y/oLePLjaotoPyirXNGscvz0eYyBXmL35iYsCYTtL0AjuI7+Ej45RRg7ZDqK
LY0pFsRgdYIcW4pm2q+Hq5jB+Npd5/dTDyZ1U1b7EephhL+mtAElSzZKCZXzJwXCJmmlk2pA6LRz
o9ecOAZncZDp8yflzSxaFdZDbQ4lX31iTgv1eKd4ay3gd0mV5W4Jwz7YCnQN3H4eLvoXbe1U7hSO
z7a3hFIaSlN6PPiw44L0yIUO1mV0rVv6y68n3l2qq5tfSXS48TG31yuG6OEmeWDApK4yc9AAS/mn
QTGmdHUBBtIhpybliVbKYScwG9yPY71foM9QNl5BtvsJGui9WMoVy57CUNYzieqE8ObMzomOzJhJ
XV8Wx+PzbyO9AZEkA579rCKzIxK9f9by40E60hGzTLiil5ioUnlS5lyclPjWHON4adwLLehSqFNV
4CF9JPixOlYxTykIUPfoTs+WazrZjjzVQOCckQ3HmUT5RZ0zzuedkTztULt8C5ICdqegl15zw6l4
u9Bz92+AosmR6Fx8FI2LTTf/I7xmcPOqJrb0MeGR5M53MwsLTM6e4Br2DskquibcdZJ+11k8HD7O
woVrO+cnVEAjivsqunGQR6sQYRExeV9E34UappA8RIIMYcoHTVK4qmXBUO8wOlUtULRyoZUif462
9Y4rqePvSroD+f474DV7wmFFDn4J7oq7+yvBidaPpKwgy6jn8EE3mhC/X3g8iBwvp3EGkCD/EEid
chaxVdkzoRi0/S3rSDJpitmA5J3dZjE492zPOPEE1BLFKeywWN6SjQfVzWnoUgVGX0quL0S+Er+7
e7d6kJSZ1JZN4Rr7phmK8f2d4gQhef1SMiFYj+pjy4sgoeaiKgFWAAcxRtH9Qb3krILrhzzIE3X/
RrPYiQk0xnZvjJ2cD2iHlCjwKMkDIoxwLSYSR7zPV5lt5JjxyOV8DwlFi8ItxOwV5V+/Thm/pSAh
ycfycS5epxHzACtX0R9k7T4aolqdR151OBA9q9sNlaQdRcjsBmXS908G+QfxB5NXT41HnIMOEqgG
ZAwuN2JwVWGnw6eHLGxa77hTtdUoU7DBSJLnvR3ABD/I/uLfS+OsGZm50BsMboV7Oshs9VUlYcaA
Ou7m8k06b8xEKUIQsAB/VbPtg3UozlTIwWb9VpeM3wMPhgeJNlyHfNkQhGQCzHLQRuLqTYSGxKoH
EVS+1KiUzK2mA6BC4J5e6BJeNN+P33tlypRUx5lhVHjYqiy6Cn0SCElGXaWsh62BLzkJabH9B+Ol
qiimNlr4zD4L3uJL0NjxWfj8E8SF8heuYUMOTkTnkCUu7xwL/v6s6R0WC06+A6NFuHZsFeAq6X95
IJKNjHJ3MUe8o9WMPmsxH1EZEsh/selJEssqwbqwZTrFfBb/GmxIwD0iUoMz4SIhKK5Q5zp8oTvW
DzyDA7qdEU6AdirzkLJhnq5/jKRHhPjfiyA1IxtuZAg/Hj+WJraaAA1ZQfZSlvIBsYHg03GaWPjH
DYXKHpi7ouqPysrMWj0SHCyKHZdPhxRKjFiS5xRQ7ywdmEsVQvjdn0Jk/0AOTA+YRj5+DRr3ahXF
BezqGLcIN2G7nWWqixiB44csAfkBIXvoZO/ORePBIUoWDIWcoDn67XZ1tbDagP+1jRyjtewC1U9I
ltTcHcLVrY6JqJVdSj7+zvM2AKj36NZGckuKcBostVihaHRAP5S5oRBiyAmuazFGM7iT9vVOIvaD
lp0mQiyx8hftE6MxhtUxqJzye+wcduEV/N5WB3no5BS3jw0/XwZmNHz61yAdw6LjjyWyrpSLCu7h
czgXmfViOYCLqWKbXdCmP7XOvqTQhGAr8YIV0+QBDZCaK5sN02JJvXeNK+adMUxzHYbp9t3jhZEQ
8f77qBvyQD6Iv92LeQy6yyeCi4RBmDNxnkT32H2JEAba5cOkQQk1+WdeT4AuZWwDRw0cs2/ZZg5C
7qIwbWsohnnexIgXv8TMFaagiPfMQX23FG5eyppd3M01awaq6Qpqxl0ktKh9kxgz3M/ndwb64myr
s4WEeYC2dYa4aFfI6k0Yu2mJFm+OlTikVaO9p6mx96livQ+uxeSUJgTkOXbyCrHY71w2Hnq4Rp2z
Z6JA1Aj0Trw2epstDsdJFF7s/mCK0EfO42AEeC8KEgh4T455Yt/yxv8jEK8EMauUJXRNYuW7pVSg
64v0Sytqbic39qbs12G1qvjdvlxjlIr4UwfpaWvTJOHkC906JcGIiyD3hCGNV+2/PZira2eoPHWT
Mzz/06HXYr44XCuUVUhhkbGCYkPbBbf9dbFYUdLkY1/ppF4Enhn8yWKvFAfNdJH4Cn/EkSFjY2fb
1MESqrsoc3RVKcGZCYZK2Mvw87l+oO0xe43uaciNX29wSQDr+hz8loXdS6OxiYKuzY48HnqDrlhw
MEnjST39xWefcrLY6eAyMJu7/jB2C9dQ7F3wNRrBFvHylvqUX49WkoDm8jBIWZ//l2OiJAzBwVd3
lpbF4KLKouerK/pxL/cH7Ui88gcpsPmaybqMWegiclLu0iRiR0DEdL7mFMDXFNFYqyLDuJpSYgSS
3hWElMORpc1qOrPzJmM3SSnXE2mbAokwEwTjaKLfKonuzr8J+X2uWKn/qu4+pe9Zo0WY4NtJm0jW
xXLK975WzYZo+Le/uBp71MugFrjPl32T+jEIFxOI+4aTbWc2p3YwmQsFlGkN6nTQyvjrn76pglyp
sEGhodnrPYqVjKuWO6CEkpa4vxx5s6dDUL3fT2OcP056YKag9/W0BCc5/CoLp+YYCdDKBismspXI
4yZKFmlzhIjPBj/WnUztmQunjvVQQ4foTd9Y7nm+jpkLOGBuPis5LOzoMKI1nrDXZhirLzd3Z+KV
66fDINfXCAdEh5zay9/Bs2FQFS/Ggg9+Sgm3hHutAoEGzzKZWicscBHkPxmrVWYKzJ+a98faT1lA
m16AaktJmTT/pwSHjxFEFn6rvn6AJgGobNMXLluPz03Tuoag2VFLx2c0TKrLW+BAeM7Qz0j3731z
2i25uh/6rXhcd7jgOYVQ0KH1Hcp1kM5seIb9P8QGzvkX3P/Tc/0lp8ANmW1ko7rXt3SKJnnvoj1U
Ah1P2/k6MUe/lJNGh2+VRUuix7CCEvUC74Ddt8qlX0A3OZL8stiSc33JRNRC5qg2ngboVogvcStV
sdqnRXFkQSaXEZpjLEnbLR+EEAYI9IO12xZWWpAC2HmQkZdT/DlGEJAUT3mfZ2R9FNULcU6HctjE
8iPZmiKAGvxMrqyQP/SwIhHzroMO8fDBFk7hKbz5RsS2adra6vb1004eXQcu8H50toxqpWJfjai/
vNWR+cYMAy+kTI1bYY4PHJ6IPEJ9lxubLowevo7zXuZuqhKhX8JABMCdV9u9+8hy4AtSFDsT8hWH
RvmBdANYUhVk3rRtUA2Tl5Dsy2aYDzoVVMTy3dlbXZ4AV0HvR2SivHKNiCcwIKPeeCpT631BmqJF
APmCw+8JW562EKkfSQ5Dla0YJCIAATY+3uZOfpOlCZtRXM695k8k7XzvxplbTCltE0+UqvwWzbmZ
MidyVLeojlOTC573FkFbhf5F1ZuDMNRIYNDKP9eRwDrmw4pTivuJMdDMygozawjW7oKJx7+Bhii/
usup87ZPMU37BvZOZADSzgZxF0c3XETpFUTs8oHU1121rb+KVto47Y/Kv+QkMtzlaJMwm4uV+3M9
EgdriZ2OmEWyib6L2PTb44ACTfUAvIm429MepY9ggguvkrSuwN6krHidZ8N8PHwsGD2NJej/o/6j
nEugSWfsYbnw1zM2P17bmlNrE8VMVgboIfM0ScbI6iog4B6ksUnGk8X7CVo6R4l6GabjJmgmH+jF
3RHAzhhzZ2Q2NeRfRNdFYW5owwb00qk8xX8rWEi0+nMFq2GAfoAwNxhKQJuo3Mhd0mpGmKhzJaQ+
JxJKvZt3yYTPX+GZXcjddot9AbLgU2ayY8ZCo5jJhv1oksYAYQVGQ1z62Ou47aiSeh8wvLstHUTg
Tg6M1QCxhR/+ELxqTDLNH/dO2ipOXID9i3QhAn5ve/BH3uizIAJDHefbb85zuEkxNNP5695EyZNG
CoIBkdVCWNl5gcl6vdz30y7/g3Vx4Tu5rPfdiEvOpKIz00dxlETsHTU/uDD7O8SCdi0YMxgoA3hZ
t+Bdp+aSnGqfwT3ou9ht6JDvdi+e24saSMUGlJSkdChn1ZNx+ROb9rsPiboT+CS+d+FJStlDLw2y
lfMha5F0FQ6xNwIQoZ29FU176f5kRwfqWVQ5JNlwtjwQxKNnUJ4g9IXg3qmhLSedxmVS44D8mvUi
agqwVlu5ZtKnbB3p6a0eiAdBpQuexA0JXZG0DsovWRr/EKxfHQ0qtnn1iGz/HIsZYTyjk+l7jKM6
PeY3NPAmShAPbUavhiC63bG3Qj9DiCzb6QtTD6SrLL+KG606DMX5zV0FV/kFSouQlTJcJjeA80ZS
OA5hRRCnj/QQqz/yyMsUs0h2M0ByFz2nAj8WA4rO/YQlW0sqy30TVY9v093xXNuUBMZ+mOyAt2Ix
fyp+ENn2MSnZdzMtJHE5xBKrOEMXv0meBPrhgypZT6V64UDM6wc4N/hElwlW7RB7aM4IcdaGXW+H
6EpEOa8a/Vr0JgZztFxZa1VVUZtGPIeAYxKzvfIcV1O+nBJcbdtxnwagh5qIFgP/X7BprhRfpcVG
kY9FySyG0qi7S5/WxT9dPSZeYa948q3yxLFgZe8vl3ZSlb4q9E8ohqqSynCfgzXwE2p78n0OUbN6
YTkqVitoo/ORsL3/IIrR4/0LVVQA9QQJNT1NQA7rsf4BQr8R6fk6WIzDA9w0tYl9W7aqS8D56Dqm
ColnNfyafR9t5AXNe4w+AqqLY45xglVWy/e+MLk4PT5jyO4u2rU7Yl1BBzisQGe/feW1mLXdhCLW
DtRqWQYm9d0iSVgrtWl1tLtmPs783e8kbyzCHdhYio9cAdBtCyewiolreIrad5wZB+7pMGqULG/H
WMuMNsMw62arqDfl00t2CCHCA12PjEzhYR/l+TOflPTTQiTqznlJJ37h8yVfx1gdvHMhKVTrXCMR
zCkGdCLTivW9axTrsR9syNmdJ32AsGz5W1fQjxxohgA/cGOaSpmJ9ucOxvCOQdSocPhURSrKVcZ/
zAsa5YwUaNG4DMQYSm/ZiwbsOzZAHlpdB6ZbH+2D7BT7zJbddT/JTswxSmze+5Bb4IH1Yisu8ABt
SPV5yR+/q4iW4hvwoMJwtGlOTcnTALUwlb7t+ME7mLtjGZLLWiaE4z15nKNLd9l67Snh1LalZMCu
Wj2L2gmNEcPIeSM0jNDGMoq9+catIopu1BZyb9rN6DLB9rrLOfo/CEL3pL0OSFy2MeRVovkW9NuV
9dWGbJg+GYOQK5+ZeH1H3dQrzx0UN5tBb0KgthAPSk1wfTi734Afu6ixHibfCnIONQoKo6uaUkEP
GR67ok+IvPjK9FdsV/tdmaRDi15bV4vvJVlEQH3VInLJhwZoMekwB5Qn3nFHCa8OrL+fOimfEOvC
ixoALFTqoW3KQK+TVswqs0gRSaVgJvRpgGZJ5086/SHHPo/HnmMBYrb7HsAa8VU95jRyDRJdXJSR
/mCoB62lyQwY7TuKmEFvb4tzSyaDyFVOQRzHS6r0FuVf/YX+gFKnLmt3IScxYrS7cy0JsWiwIoov
deCuHB31ZYAAqKfTs6DcxZZ0pA46t8efzkgWH4pjS04TBGTJByLbUsSEdzOzUTKtMNAKz9Ssu23l
0eUyPnK8HwtgTRIAxfMQeBTfW/hDrNZAUvafdHfQPgyi/1gkFPIVqrpyXc6Cc5mhLiNf1LIfKcrw
dDB4BtqT3bbjipoEXBf9JqlfvyJy2hUuS8GOSYn8TbKjaq/Gbvz45nTaNuFVoAs5nLfH2SU17Yi+
dvrMHRFVxLmU5KQyCzOCA6sRrPrWb+jdANdayC1qUNt6aj/8Xg8L2YmH4rqdsnwas38/2gCENkrU
YYfpbhCqTvFwiClG0LyYcqh5fvQjxc4YjUCbYWWxAO2sQm7HLEZnZekxrvvsAS7Nc/BXiwXQweaX
QDw1qMqby3ZjVhMF5wsv1WHzHzaxAHsr636HqxmUShB1UKyz2n8KkeNsSzi5pt8E8V+ZCS455K9B
wxjt0NTjwhqLuSb0Ek36KkAsDb8K5KTyG39JOX9w4ulkU62jV/sSXAK+lxUx4S7L4r6KsWZuiTxd
AGv0smd2hCy7tAHgedMetbBsWxrLdXvJYJfmje4xGmm5mwCuNzo4mOykyUr7EcNienu7oTrUbGfj
/RiclxsixO+63LNTn3Exx0J3Cx2IbWDk5tM8sUWakkG3aw/B/2BZR5/udMcluhUrIRXD32QiOMUY
oV3u32gUNWaJpcW5yuXKnhbzdQ2Z4qakVGmqjdsCdSIXhko7SOLLsR9oCgsiiY5Ydt2Gx13iw+4v
C+zeI6FNz7nQ+Ztz/gZR0HoZGiP5H9vw2QitHJt1QD44FcyNFVm32oD6j0SzRbCUbWjKzcXUNkQ3
ICcwP3eqORIW2215qhm8IKZGzJ/l0hj1GHzSP+KUFvJgVy6wF1mkRtPBu/KLDcHxzQsYCYSVJsWY
BtCIOKL99UzQbylfDeIn6zn1gpmwy/nGRZsmFo+T44SwgEvWTCKO4mcjf4NVdLi7ZGyLJZBqRmxr
8h+MYoDo6TnVVU8jrws02AKSmn6Q8lfy7TEkGcqz4Jlmrg7klsxaS+tPfUdk7OfXqWiN/dHjQGPS
4xE+v3iHg+KjgY4p5DDKy5MPIpO9h1AwB4FOB6PKDQlYs+rMMyFMmIZTbc2DNs1+GS1r24JHGDiq
Zwr+KSSaxbSgZQv9X2WmzbHZH+OgOChRJCEtn3SFgQAgDbsqsdzQrjn9KivXCVY80ZCt7QF8giSw
w8lfKmshpUXITT6/2IFksnpgMYNDb5w4GRY27JSwfvlSMEOkMO+Ns6nh3QkKhX3Js7WjRldrl9xG
ZOhCftR3C2zcfuVQnAfm8PRtfDQ3b7NMnsL/0Cjard+lHkMR0FsLi5UIpCyv1u+yZFspaDRmcK/L
11fzg5WLue1nGQFgGx5lxqaWg93UpKUylC+sRsgticlXO287KB6/BPCEWfRPBLfLKxnk7TOB2yJ1
VS8aeW22U6OyoAtEYxFCLDJUJb8X9Sxniq36+2b+NWLm7GYTVcOZcZgdv6HPtqaPL6xJ2nZvYBDO
qkNz+JPe0De40ubeUA/IruR2jJqBSdWAcy8YVwdKEqILWn2aErylEiFm6EYMXTq51sQcwcop04vG
3mT/1K9ljcDO2ehXiKsaIXZ9rXurK56YoSoWBZ0nrCv0EdMOat6MwBc64SQCod4NAsMQhpOWy8de
vUuaVRac9Bldp6bqno4Ki3gtMN8KfcyMhzt5jVLUI4gkY9zAqszJcY5XlT4pMjtZU8KNAp1fX8Cl
rb5OCVYh31rW3qPPXmZTurVeCc+SY1qxUOr52u7x2sXDeUwahzOkXkUyZCrAWFeZ5ruF6yaf/U2J
5bDbefoaWOiableqM5zYXFRRigJ8Yi8kUoxIddJid634AjoOChJzkgViaCY7PIDIm9WyRheU16WR
sOh3KbYzzy0qMk9uzyT97WHjGL3VdYqBIR43kyILOyHf1WIQsPuWs/TuJ1u0oUmdpg9KrqK8ddYl
D4NWgtXxSmPDCsYEKHrLsiGqfLz2jrd8OX/qtZID6AIFQxDZnGEOpixyQMWcu+mrPTOTEaKxRbvt
1WOZ+WCk8ZtFEesNvGjPEF48+TuMDujahs7mbYUlRgbd8RXrWba2GWT8zfQLwiB7Q4lD1g1h2/TP
OUf38opOY0Y5UWl/ujwbURbKhfp78+KQeVq0xIcttzGFeVtIn9IbyPf0Mxe6D1C+LhQ6oLoUhbGG
Dk2gBqchpTQdHjmZXbyb4HYzLfLE0HzCpwDA7JXltL3Zx+550pKr63wGH/e+OseVB4bo5jfJkzxR
nUW7sKf1jF/WghHcCRz+m0Yu2G00+Z1KUEfOGofcy68UZIuYLKSFYQUZ20FVpz8fjCTpSirP0SRM
hIgQZNe3f9pJChIrO6H7sEZ5eHqfVcCWDa8Qb7rSXy2HP13aubj1Ckvz0insIuET6pGL8GVxu+fu
/uQ3njRT8q+MsckloktIjrSMYDHnnLbuWEFuyW0H7flfaPIiucp3/EIbS0ecwGBfbd4mF7ZC0e7U
HX5+Qwp+kCOs2gAkncG4LZWYrnCAvTA+ZKIELiILH0jCow7p/rpz3oRO+vrZPCgEoro7L+4en2+Q
AOp13LO6sBOHwLUvd0Lh46NvnjQB39pkrnlYbJdRM348wjZYN8Ip1MfGkOQPQ2wg9dS9wTNbmG6e
M74ayP+b86Kn0Ox70nnDm+FhVw9ZniwyuOozLZQPbtiGpVFesqIr8il1HR+jregKFAzQmYAd1nRa
wGKIJOH7yFYync7VHodP1feX8aQZxnD7xFGFP/8oadPdiGLG6wGHns5gqsL9h4doZA13rfJkdTzF
4oexsfSWl65J4vYeojboBbL4Ls9DZcvgg+Lwbo+IyK0IDSAeg5tSA9Ns6kvkyG94QnSnRkUKBrNk
fB8ZgXZ3+BOhg0QDfWiEr6tMsTDVCKke3Fmjvypl0s8n3238MLaQ1DF/YbOyG8uKSVTXPJ6m8qIw
sySDJUxnz7LHCEXHWFjaB/uFzeWsT9xKQhqUS5jNMAwAQj7rOJNmqU6ZbGSQtEzs1Te8I9NTgk6Q
C66v0omOpqDglJbEKhjhu2UFppqonnon6hrnstA6GRwvec9HGzf+Yrx1q0GWIIDadGAKC/TwHaIB
p49zscYkh39CMqAWUmSvBqRAppnXlaz792nChfs4KdVIpV6cKhRAvWimJZHOWndmTAkpHsjLLmmC
D/ZY9x6ZjQfSL6+aETNixo3lZ6YOl/rTqpyUDWsJZwXE+gctJu+IG82Q+pP+34X+R/jPjCpXl5rC
veKBC5wIgpf8BK6rV0SQpnGJnTWln+lbCiOQS0SahPfB9h1HMSsIY/tAobfDd7mSC3XOwfWm7YGY
+3ZBZ6sRQYdRESXrbCqvAWLD/0EgUxXWExmkeRU+cTgzhddQ3IeoSLr3RA5NJSf9kO2PlZt8h8sw
WTmNRDaYkUoCXQYmxHkk1JEgFkkyX0s/dNiiSsjhkh0kIu12RfeJ/krf5cMFq4k1kyUGFmEHr9e2
oiq7iGxBgzV+FQKvJJRoACxDfYC+UDxA0ZysqEzSQgRQ5tjgvq/cx891w7TT3ucwXjxjPFF8puP+
8dk41MGbPn0vvdhJ2MfQ2HxVDd3cOHVC9uPdB+vtzTNcFFJZ+vFZIIR70hKT6Hw70ddZHis0AY2u
Ml6IAH05FUWQsoGXM3mrFlgwEmxQT6htx7q6R20iQesIE3t+wu4FF1i0dbUEOgrzI2/AJugv0noU
bonmGOO65Mvpoiyintvdk7NrfCHq/JqFJinmHXTcmsUkv7H2IEdtCSYQW2q9mhINq4X41A5FijcC
M3j5sNFJR3Z9213eDLLyPqwWbyR/qJvdveV1go9vlgFLi3a2da14j50hcgGtWllqUJOxduIxX7cb
akl3FxPeaJ5XmBd0+tmuMo8JfYa12Gqx8IUM7akCtp+O0o8V6YZukkxXFZFMXyVxVTaMRsAGi9yC
+54hAFbQAfL8DxulY3rE0tOdWdPJHdcP7GCMJ0Q6FALte6+wVIr84O2zEfx2zAGVODRv9fv+Otcg
25/f+4hkFWJqQ1t73cIgEYAAOKrz4ANoXuRyDpcJLHpuT59DXuVg1oto2JwOcKMpdrlOzrIXckKa
YiTd0FDIh6revMpD0E9XcQO1OoKWsmUznlOzReGYmaNchLCPKuUJ6IQ8oWAYgwHuzQk2Q2kUdawx
q1sEOOwpMAD20oIJ8YHRGEQaZtv0dFPlKreTlVZSsOlvl7ZqpXtzvbM16BPTiWcoSBknFgWq8pFm
RAM/jJ/DsKhmpvf7DhxKxxJ6yJaU3Qndg6NF5EcqfQaY82sufSlg5IizjCHqrFL3kMdh208RRNha
NY2mtHmRlu0FxbupCMRcvZ3GqnP3P0O6wWYUcasT9GUIPssL/WXw/As+RuT5lWwT/bTswFIu+gKs
ekT5X+CjmYr42tBAiMFVqCBM1yCgHUNuoW2/xCst418jSm2dz2Gvr4xUdoDO2ZTT+XexmIi8wPpN
M5kbZl56u+lN/VhO4sZgRDZjSGZfKGwt1EBWSIwjgEVQ75K5gGPzgCfKl+u4pIc0fAFXDUA3mLZE
bfOWx4jqPg6f6p7bFAav9HcY41c3BF4tRyce1YEocuu+pGRgFoz2L1xr0yuMWh7p9AK5chHqzCTh
OAl7V1+4GXbIhWTZfz1V9m8cxJG3ewOFISRyZ+SHlbPcK+NdYBI8Oq0OIQg0+X3LBCIyAhvooji8
ZuVKfudG7yTRQXM0h1cYjo8fjWQTrVXl9+i7YwxppMSEJVDWahu1Ulp+eVUFz51YUEuZ/vKFrrjq
qMTmJ46p9y2NvpMH88I37a9OX/cebrN8B3ZNdAGx7eOeJ91ckYs+cN3QySCY4MEY2gsKCTIRG27s
VnAzxOevOyZ/o3w9ks7yzV7vIKAtjdRubmVTb2stCfssTW9ClfRplGW/REP+0wvdOXpRyqwIXzg2
uY2Rib+eCNtHJIP1vr9KMH5h7G8mz4Psz26hY+PMn9O/GsnJ7d1gmU/viMpkB/87hcCIyxh+lZaN
YThZbQSfQxoMkT+Bkk85xlTuiQdmx9yBJjenXPrkSs7zg0Nw16heh2kOE9noT9hcm+pTG46B7Ujz
nafoqkUJp3P/0i9ET0qmfB4p6g0hERY/vyfRjSKGbsMU7X8KHVUEh/Ij06jxQjrT8kymjml01eIn
5HFDQ1UfOBsFGv7zY7oFQVjXIENinAOkkM4YjQzRVEpg7B1jNRvOqh4x6DnLb9Su/vr5dJXY2rY3
wWpsaDzDh5wFocPyeek1fDnmZKXp0ELcsf11LOdtxbAYXPSwiJzte8JIEjNatSkph5n9RFndXSCZ
bM8BCPC0Un967dFFKGPQ/dM+L64/NdYGIbPnx+E/LlZFIK+q61nA4ilvMmIjVJuyQ/epgQywmj0I
fmA3zuqE9nXrqOi6GSNsg/BG7B5UUmR+SHivrE+736Nb1hl2mBsISyLB/OF+9Tn6CSrrs/5zwEHl
mkws6xLVgkx+cHwXro0ybqdvXk1lKxVrCYyNr72wwNsVK+6ShbwxV6N3VaVt2/9kRHkv9AUak7HZ
0ds/4zbNLvJwnIt1zTlANMyhdmQiey+LJCnaBRu7DqvoGm73R9X/vMhc2XiZx2y+rhlQRoGR1+Gf
p/MLVMxatEoeaj9qTlwvSMsjz4KHOY28IikiYJLsbel3GIwaPbz8Tle85xzrsOPtzw5r/16jWwQ7
zxAuMbIRz3lhQ8gOFuu9xMPTWJsTjeBg9RiSbhx2OBdH0G4AjuhLeMHA0pKVT/nFXFBOyJJCd1/q
ArlxByxP2pR34rkn51vEp94oinvZ4lvlflC6kB4XTHv7ael2hROl9lmY0Pm2Fz3CLGgQX9jsGDox
YGY9/U7yzvQRC6fF6+vkZOAxutpWHcB9kTuUves2Xp9fQfT2Pxd5h5qFntRA2JS8QmN3myUGkQ9b
SEoZqlLcBKUKPdgYU9SCl+7N5z6fqNhpddV1x3z48yLalq9dQYdrNgSazP9cEcj/zgck3lhPLeI8
yQHn5ebLMrpg907P292oYrnNbgrqLP2hSrteQokaFdeq1X8+ddl2iMEZnGdtHQq0ZZJ5ekj2JR/O
FRjPejVcgnGsaGOg5n5NnkN3vHotC5DgifrwyKSWScIkmgr+vQLCMiy7j+eE9tFaVQPLzwjQLf+J
G2TMSlnnZMCs9tqnNDi0nlhEUrJgcQiYD5LijR2JnspiT+Gy+z9c12QAcqxRvKoP2gVYR/ocnLGO
6nAPSGySgRTTnaqqRPDNjwhMBD/3na6fDxnIDyYwNSAeQ+TbJqoT5hKVcCeIoBqYVT6JRYh26eGq
c+yVnQt3INgrP/JWi2F6fEscvJtUCS5cuNW0sVpFxO3gaCrKOePzE/j47BM+H1ThSX/98sH4hqg0
1oujjF+Dx7XqXmhTIXlmas5o2diQZM8OcvSCTdnw1BcWTd3bWvgTKFtyFz2n7Pygz8IEhJHpDsVW
eajcWpTZTDuBP/7Fs4AE8VS3reM+dkXNR7Ke7SSg542P3ZFlR4Ncx+pc7qGZS1TXnGOmRVxyQ5RA
qtgbWi6W6sXl23fJZ6vBIcK74sptPYLEH+Ibc1TeG3s8MkIheNJMNQnUIRdVzAcLiZImz67Wx920
gtWgsRn1a+7HfJ/25L5c5YB8JMqzTNaDkih6Q2IwTAAGbgKcUwssbGAkLFaWD1PNtGD01LGqMPeH
tm2vABjQqKBcCUnSXYUaBCVm+2kbIFKcabFituqzyn8VwDsS3ih5VST2rqYngQnwdJOG1E8qR6PR
Y5SYTD4TxGTN8QAb8G9IOEfUetGJuru+qUDH/IX2/HbreGgnq6wwFX3nlIJGCt2IJy8Thd+5x1lV
j4aNbuLEZEnDqKyggaQY+SjVYrNH3jhGDsiUj18tuoY3H47O3Nhis4cHj+w+ieO23e+NuNKhbNlf
aZc/XNL8s4TshF/lDx/vuxk9JNh16vpIzYQboHQJ/EAq61Yk1g805ccRYRKxQPAyxTfnTYrDJyeC
livc111zApbi8H8CDTyl0ym5lwHcgy68zWNl182tj0BIiYzdifZhfxeEjwHq2m9KxajBBKxnKfMG
3MFvUVZ+stXUeFO8DxjlAa45pAt0fX4sqCg9wxWJOmPx0AeZSY4O1m45p3ZEfdbqRARIuJVscf9c
ICGWX6gqF/so0fmPqA/dRHirB5d8IlowGOSPWjPAR/OQNOp7Ft9m9DXmAGoHM5Xe7t42cAiBwLl2
vnS8DaPTdc3UBCk6a3hLO7P857CSMNJKbgeQ8cEhsmbIwcdSiktNtMP30QtBO7H7GEOtXPQ5KJLq
VRF55gpkofhC6Xql83hR0P5cJk6730/C84tPzi8bdUgUYit8mR0WjMnTfvQn+vx4FDZuBF5hgjWl
NUBNYgzsa1VmSfmQ8Gi0XJHssvqNizj4tWkAFrFnhcZpyLq5dPaTal1XywNS1tWbiGnKpDZ16dsV
yzNnTzKtd39J4uvwdP32bV/vgiB7jrK7nKRWSdr69Z/pyYukv4iCkGEj6Ymko7Honcs/vXgXEZ2U
nVIBEkNgtTRkKbFhwYegC2O+1Ke1v9MUnO5LhcLuksh8ZummRcRLZkKxoM01mUmuKC/HyWC63Z75
wrdItBcEvsm1rIpYTRyCitAdNHD8TT7LFtreFXckZeM51K9NNujUd5wGz90hQ8+W7L8TyI6f5dGJ
rIURVBrGetBsfc4kMV3M8emAfZ7olz/NMuXNO0pAV5edmERmPNKcCLMjlNfZjroQIBkNButjWe5I
0G+ngqkZ/2CcRagnnoHW3J6y48ibZg+TS0mpWt6xWC/pm7cVCaEdtsO12etGINslHIdugELBwjT7
t1dLGDYc+cMWwvz+v42RizfFayah3lcid8eROAkXCpbg5sctx8mWSAo/eU0fEzemjtw1GjECe3wl
ejygHiC6FzQEc3pCNKt1o53Jo0gPfLJuJv2gWqd1Zsfq1wS40cDjxhoY9+e7W2LkijhjA3q6Cr0U
B5WrkYBJjGET5Aw6aDcAtTneDy8v4BatePeC0MFwR0HLHNGOuCge/+8VL+WtWK+SSnRMorjJAkGU
WW+LgxaWMRvBwVDdZl9qQdmfLyLQxb2VgmCs1Ml1+rkKuPGdhQMZx84UWTj2aDBBwvVZnKYDNm9v
TFcOSQPnywzRyGH1AFDUWhzjCowfkVfDxvXFizAV5DlHZksmXOQeY8uNCTco4GKYk7F34fuFsP52
ng5bm+tB78Ru0DXbIU/jIrzK6OjwR7beF8iOfY5Pox7Cv7qWF4hw/+SaadpGCtrTIG+cbRWa8dNt
KbrzsvHK6jPXAa5IM0RKMF5G+xtru48aBxmGofZFMoirg1taoRg8vtq8I5Eeh5n89/UQUiYIbret
YKGGFrFlPOdh9MN3iX0WmUqad7csMxBOfOp5d6fsfkBAexecQkGMg7Joq4RR8y1qLE+hmHOseV2A
agOrj9aucPFSEDutETxMKM77eBMFz50CXOzzq9urWb0t7Ys50du9T10RC78+cGU1rcftKarfAU4F
vhhIVuOhc9pN3ByettFN1pwJ+8yB63cxx3SeSYZ9FBCcMzrTgYw3b3pVy6MNINUqamMgNWlyub1e
7sZ1m/b4g/XSFvgSuy95rQ1inWHBkV5HnDc7mCOeTaHIlJsoI+8ZFUJRwoHrPnySEd4z6m3X3YXw
zvWQIgbCYcNOuUE6XOPV2tBLOVRy19QEEuwkAYkDoXWEHtASKOmUnRrz1X+6KPD7GhuECyKlJulO
H2ViR5+jXlbz4EDfRN6rAEkVHgzfe8dR1FcLZRMgLjpSJBgCDLOKjZYn7pbHwcFbTcujE58cTeVd
cMM3oNokSjalFcw7/vWF8OuZSwEt57+rw3AzPZcIWVX+4WgfRMsdDjR23MX78nDKuSYNzlYnyBe0
5FGeGFexZEdnsvWPPLip/uIO3QlQYkcZt1tnNcthoxCBZ9UxqdJX40ZOGwcq20JTC700K+08uj+z
GR7HawB2eZCD6PgxBgG5JjdJW/VHY+IHOGFygwRKyrSjlDGHwxRcZuFauEHSuFCoDrswoMIyjCnI
N89PM94LJm+tVxjYfgRCs5Tq/QL83pkBXuYUbHgNkawi1fyRXwubrkxZ1/z6CzLKOrbi3fdxSp5h
jpqHFIm/64CTXeW7CoJm00YI5XB1Z2205aVYg+ue/5bomXOzH7gmbip5Iorsl2ax+CPt7JBdu5NI
h0gdhWllzeHR17qqQ/F2JpUwsGbHNULXoeIivc0ElNtNjgefIAu69wmC1Xgbx6qHW3CrIbPBH3jp
/yk8YyUhUoCjtM6+tNw7ACuTfuzFnN5srUtpDH2cvXBmhyW6PLKBxJ+hmeHkZpsTBWf+td0Oiv9s
Ka/nmOnW7QW72NXtZK/xN6ciQJctlZCpqZLpexEl2olvVb3yLD+5SR40cjnFRrLZADiPYlAc5yCx
t3lo8urlJCAGfcnCLxo2MItR9+9uY6c7vcZ6/XG46AGDcAT2KleHz6vedB2otO58pfEw3gEn1vIg
SHZTxaWojbz9nEdgwmkIZRpPyv3VpeRbUurXOxyb/lkcAG+ivGHuujoZ7ewkSwHe6zphxBhKFLJ/
p676AzXfMrGQIsTxWn9ae4hGXL0/nHYta/NMmn5UIyoP6xj4w95qU6O5s4IuFAFN7gcxJ+rsY98r
IT4SC9UrXyKB4kEMTiyJ+iScUbProCFlsNwSWEX7lX7VRE4ukrXLwBV3WqN6A62gnIaG7ivEChQp
K3TcgEwr3g84NoOghcKU8e3WymNTpO+4Fv+MwzXTHa2jETM9fhfyEHIcN2g05MbuHHYN/YsR/xyE
uJoWEar3GXkRNU7Y5xcT5OPON2O0DgmnniooMQYVmwJrYRhfy83ZSxXkuLFsY/+XGjho2G+sgG7H
W/xVYWoLWcjua9x91X9CoKYLYd6Zzfp0K3Xxrl94JR1uN5L87IdqZFMprcBtalgXhdaYCvsiMvIb
FqA7OtuecDqtxV4WUBERGvjdN9LROnZ2to/FyPtXM2ODueYG/FJ9nH9xRMQ6+oSX/o2Lsrw8p4oT
YdxeEd/c31jnW+JY39ywj6kOad7s9+rRzWyEGo2uYlTkmq0TowZboWLHE/lYsjXTdIK+oU2UfvNK
x/x5eb5ENoQqgc64rIwa3J/JTBbh11fV0oUk8CEH/RMa91gzwTom/sCX6dm56ig/p791cRWu8DPv
mvX3Oi9wxNijQgX1G7fPJmLOEZuVMiGNHHh1GebZaz87E0p2Unwi60jSLpMGe8TPueZJIva1Zf8m
/e1nFcOq+P0zDPdXYiX6AHfjiHz/dk+erfqgog74JS7N1yu7GERTV/KvRdbbzJVI/IcpXepkkML0
Ae3FK+EgsIKktVpCHuIu6CEWzW4QcxKY88st+//xvjO35enyr54G2V5cAZlX6eH8MJgIBI+d1iGx
XjXbZzHazDN+zq6Y1UDHMC5NqdUgutw0yFBPXcVgdtM5e28rj4kZ9BFKI+IOhE3t38p1czcQPnbf
Z2CMd+lAEj37T5lsONVTi6CDrqUF21yAcuYeuM/Ra829DbZb8X1bcwnP9EGvhBIIsuEX8a8Q76eF
620gy2foOCF0jAsSgaRZncOO5GDeChPCqrFRmnmTkk5xWkfe5xKRLs5bGb+BhfIqTO2xiD2IBNGN
w8f3fdUu/H7MzDdc8xl9s7MC1VojG24CVTNaRb+tn58V3eeYrXoZbCuCCLU9vIi9EiodKqVCwrEI
jODUZqSz4kB6fdnQIw7CTGSrmDegZxWMbjyckFTqFLJpa8O8P9HExUPesB882H9LXkMmp5KpvvMP
UZXVhJASlbMaIy9ff8XiKZra78lmy2wnW3wXJac9meIdIuJe4oYJxNzr/4NnjUpck9cYLLCM6Vic
hudmzmYvtZSXInGGnMreuJpo9g+1rNHX2pUgGfcvlq/eWDRK+OdTIgxpogqYzBPbRiqpWDShUpgp
r4XTsj06YQ7UGcsQWkUs/OlLtkKWPkUSHNuWMXhK+coCTYjzIrWf1m0BUlva+P4a3ZgK6DsxrqjS
aLCCMdpjpOSX3M6f0ZssUkG0or8OjKXYl0p2oGxgLbPU+qSMG3VyUSHEcs89k++iqMCq0ZxvWIL9
JIruDX1hh9cFaCPagnOWr8eM/kc7UqzJeLHcPVOjwyywuuEJPtCPHwiR7g5ncyDQglVy24SaE7OU
d0RUhjasKBunoWZsXKOU9iN1fU1lJi/RjAi8iWul7rMyMsGtdM5ygi0cw0Thll9govITOa1Mq1D3
LvrqbtkepctlQTTAJwhldPbqtvjrPTndu0+JZSS2bt9QrWr1ddCH7PF2kILd5WWXgTVGenNYwlXK
cXi3Wg57W3Lg/fW37j1SOazEom8Ps1p19ztRqXmrOH6Afpj6ME7iAD+HivMvTJonaWrAdyXodKdi
iE2rW+wHn7070pUeWzM0cXolk7suZQ10MnveaHB+DSXxZMRYEZIcSlcstrFS6RWcFmFXrszcYh51
RskSFTaFR5oWHxvz3BigRixoR/OtfGgHQvXjOv1fE9zLKiohhsyKRMj7qRC62qt/xQs9q63wVVZe
U5c5KW+btaPzkJC5/zeI0hrktzJZJfIztp2CiZirS/J3dtlOuT44ROEr0MbAFchhfSyxP+Jp5lPN
IpbAF3uGPPXDVeAP6p2AGfJ4tucRoXJoC9X4y9uXd4ZFrww7BCLZQJGN7ESpG8WVp9HP5EFlLkAF
Uaao9fGKKGx7CTrvy9a3ho2JHKNnDj+djJ3lxxbFfAgs3yhKae6HDGyLimhiir1j/GQFBZyulRND
4ZSsLLTRh+kNjgYMR6ZxxeoqfQI5XkmTKghMZCI1YDCP2y/qOmA6Hfo4uiN/IQqWNWTG9auPKgnF
xt1DlUIM7jGOcVqunEXeyXV8fcVCo7qeXZ1YvggwCUHcf75tjbjESAeXRV6RxI+u/9ZdZSuaLdeO
RHL16MawmkQDIN0cbe4OHDu9IHA3YPn4O9YEKRy2VcjRsFvWwxUOBFRm+8XeCkQR4r9PyYp9hfLG
IpEES3XUPc0zCd2FzNHKSJTdNSPdNNBXE5tGXAF4RZu+sJVDOAjbnwB7hRg5+KUuvIrmNHnsLEhp
a2god4rewvBmiyKPNi4OLK+EL4FMczHE0D2rYoRKzhz62cxdHw6PVqReWkXGyP4crPnhoDLjbaOy
0HQoK0HuX08kDiXivDPWo4K9vvsO9wFaZHQf3muWJg5Fz+MuLsYPm5IyBVwATrkTLgZBUuVKeCSW
qT1dlZCupT4Je4o5TKTkRTzqctLPMr2pMYX2Ddzg1ZVlwOaf9kseLNGpTmuNohdr41iG6ey3XJZW
TATsI5vStBLXECwQbnHqU7en78BEwLms86l45VIeT2izmIzWctM6fHydgZCr5uSsp47vaEm70if+
1222s6GQww6MvIAPnPiVHpzGIr+KcVFqd2gzoNMZdqBLvMBJ/WerZgNCu4vwyNIvQNlAgRhkvBZo
vLIOjuUexfwg0nM7mk/P8EOYndqGH+vtYZYlzk0uJ8s4zoOOVzrF5qfqNKoIiujYxyNAmw79+LJy
KDE10rAvCGIrmnPQgWB7KCktl/rD8NAwlyeJANvz3D7tFALcPtb6CVGae9qW3lNzfzyC8yWCN48U
hT/hvYrQThxjsN+0LLte+qLvRMNLrWhA0w89m4FqDNw1rMc3UIUHSX/1ZjPmELJhGmamHH3/lQmk
fQm9pYaqu7bos0bs3c4x+EmaoHhX5u9C4Kpd4YNquOGCfloetYpkIpiIK77owo6RhfX/LoeAIz6K
5q4xkVfvuijIrDR9ktXVa0q5fOudj4CNK9QFiBNIpMe7t0jXcBRN/4itAx0wcWPjHSTUspUhNEsu
h0OO0uABw1z9NZTC6cSmshZ3xe1XPXRsb072iWk1N51rJK8P5s+nRO9ZXDTSqaDToF9jAv5wuRR0
rvKEolXOVEmbT6mcxkl9C//m4M9hBzojnFt4KzFfuNzQqHFQaE1DYJsr+wvTPf5S19+sZz1oKXsy
6qkwk+Aj2lYElx8nvxZVqz/SpAQ/e93KcFdnO5Bl373Py1uaulgoTasSEqNz+VaXZaq45tjTlJLI
MvKwpkLWvn3NXHIVbHe71dHPG5f0BMoiqqmk2wNkn6RTwcAzl9umfNO4OdIRpACfqAEs1dXRsurG
sHQ20IIlCq7YAkyatCf8fOqHJ4qYwd7v6OM/Noc9vQm1uqo5JNAQzJmaFnDV1UUgYA20PGEq4WN0
Fz4VXKONx4RMa4YN60PsAmanKEJiUqQ6CXPDLUvbY+c+tYppypU++zlffQ0fwF/smXFG9IiS/2wY
IH3Upn0u/JupMHAQau3E8emwSOXXOHiUj7uAmukj0QgOa69buSh9hTABpsiR3qGwWzp4+Tm0allT
YnFt5PmBKHk9hBfFiP6qILSExdndB3OViqaNJH0OOAheYD0xvKDAICNm6xGkCpnm5cYRgY0ykbq5
JyyDLYzrRgFHX+RrSlprOTVnLF7XUJjrn0aCMXrkIUA+Q7RJB46e2SQsXPmjYNpErMpJbRFrzBM/
mwAA9C717b0HZDPKdtvBDjvBp/Qn81hzFpxvduopX++Z9GoNn6E56M62wR4KECIMc9OcS1SzyaeY
iJlr/LAtHRISutb98hDTAW2CkxvOu6ywKYka4M7L/LSdu+fXT933ems/JzpI619uo7GoqYLrWh2h
MwDUQOqup/zeYrxgaH1jVPwnMv+oErvlZr11pH9TGhOvAhwigfdKoYeeBSBlBgzA/gNPhQurHbih
3qbJcWvA/eTjKfk7OcwYZfftJmR/bqui6nfwq5lAThXJwPe4ztpn5YewwSbUhhRTxwr09LjVlT7n
e97uKPCAS/5KU+R6I818thAds05+tqXfx74KpaNu4gPuJ7ySszEGKu5xSvIiUsrOcGkHiGhv8Zl7
eys/+ioS//soe8xEbhRSmZ+tCfdRyywHrcdej1u5rqCVGL/AG6qJSxLwmOlDJVuFPSJDDVD+CvI+
Xqtg7Je1btUKAX/+Lm4APlLFIi5JqVe7mPAjpy2Uqh/3gSJfxhHJX5NjAAna/Q9ZkYflsI8xKgyq
YIWqveP5fZ5vTkupl+/4WRFB0iCXRh+Z9Fo38LYFBIc29PW2cDYI98+g/dWnhDiz2W5xbiXob5Y6
dJlZghUzhaWddMWyyZGjXPFBdLqp8jTyjeTaACoekT9x1PiIs/b+0kuDs2LmJdShGLmhEUGigtVz
OJ3iLYAkwkX4HGeOq3rQOxEKh/YsUQt9+mBRsa/qZUhEVelLb2mCufPnrJ0IuIT/v13kC508Bs6C
aYJ6/N1CpVnM3vE23gfFtFubpvtSBCkvH4Fk1lqC3Gv1wleb4cU2CbvtiFQoodvzyXeGO8z7MHYP
rWGvWyTjw7BqtguISut/iWemQHEbAM4luTX73abF18qjvmeFBnTQN+qeqrg1uhjIQ9H6zPMo+a1s
kPpoclqiD6tohfvsVsW+baV3B3kcYThatPyIyWKlWLfrQ4s9CgD1vHAuljlSeSEyRW2mC7iAQHQl
/pgGz2iU3FWDQcRGPCh4Fc+pPJx65BvWNT+mW7YR1g/IoJ63G01oGsNA/tq8sqQAHYe2xb/G2Z1R
lGJPMBpKE8WxfrvjvFt887T2sLy7xZ1KZN7rCSOOxp7WQtzIkOCbNZBXAhitmpFvGYIe88d4YHNl
VYDrosc4eOlWivwkGMD31zViH7Oh3ZIIiRxUIGZlPUgw5bxQliayRLBpfVykZ2NXXxgMZgfEfwJ1
xQAPIROfR2DQWFjhSDB5HqJry7zu73nY1GyoWKH8r5r5p+XPY+JsoX+yJEFf67LJbY8dv4uS1A8a
vGKIX0Dgwdbshxl57v2ypqgOQh7JPL2kLW1YvMNihAQBTfaH/jaI0I9EuSv+DJ6eHFyzJR5l8L5J
2TcG2nEbAPfGqVcuOuPLN6jbASR92A0m/uwPs6VkWflMYurF1oYuLrwVZy3/fFH6OS0sI12WyVYR
XG7Qt7sGq+zxHdbckDK7k0edHdldUXmpacmwpmIPSybzh6vFSGTZOpccfSL2k2ib9NrLf3DgChFJ
u6cRY9RffDFzBXrHzeZY39MdaZH2KugJWtx1aEhWnIB0EPoN93p2objFvKc+OcHPIOhUE1Dz3gVH
iBmHaGWe/PlQ9M4MKk2U/kz3c2+nChkcQZil9HLFkDIyzJ8PadgDMq+JgKzkCPneHIsclYuqlnBh
f5RYuHvApDc4Jh/wlQ95fGeZ0yO/e1MeDhel02Sv1fhK1rtWZmObd3pcjHntLKT/pUPNunqBLgkh
3yzuvsXQKwpPpQ/WTYq7ahBgvr7j7mrKu4HoXmq8aeA9oV63/MK0te7ssEWr4/Bi9aTDSOJIxf6k
K2l6KmQdTG+tBn48Zgaj2TYeCFmJlsHoRp/iqzc2LPPKox/o43V04VCbXKZWdrXEyhi4jCEIYrnS
LwXTSqfyWElviAIC6c5C7EzqIcbMWUPipoBgKvp1wZvkWyEkLHQQCPg51lCFqRb8mn9lBF5W/y81
lCPKdOf64c8T7TOyaN7DOlI4druxH6RqB5QQyJJcL9Nb+sfKQXvm4heVWGzhwYMmVXvkxI8dDzib
XSOw29I75DkIwar6Sb3B6NnBuutFpKLXNwAdYNhi4UHzsbR6CZOEWs8FycPq+93lc5wrf2dJbQxT
f9u6am8O7EzMKGmfdT9hxnO0kSSJoutqyavBlndU1FJJ8GY6yqOXuV887/yteCGEEbtuyQomX2ix
28E3qineL0UrLaGMgsbmz4ssk/gzW8Rrnf4MGCJNMH4Df5EhONzso+m1vrAVvg8cHsXwM1YNmowl
3Fvk7Se4lOfLLIEI0HS2pqGCDxttIzjhPlgsB9/yhLNhl/S2Uwy7WW6aQmZrVMvZDDWelpeGcYsb
JzD/Rh0m+4ptdy157sNrVUDS2m+7Osa9nh+yCcP0hvb1FTwuQsoPlQU8ruPQo0fhhEfFqDis32hQ
xFaVHTmwKQMJ8TAyUzlyX9qnptabPGFvQMaz1T+FT05JavDjJtjCaP2AA+DjQ9pUpO+z0ZYy05OU
TPpMUa4mJxSJxhUFk/cno43s4oj3ombCKlk0pkgHtjdlcx9RoZUEByMCXW1bjOXw6Spo8fYtU0AS
2u+ZSMgDFdzYAiJGmOeKUAQkyAF65irH2Lsekr6mjKKMBrPmVTE8ws8MTcEOsCOnG2NkfkpSZT53
MYqST+NGTfxXmZa58zU1itaRBG7VRGU7IVuq2HmLYu5Lw8OrUQZOyFmKOALGbRemiqWruIO5RBHN
TD0tnPDTJxAIR1vhOrbYug1TzXZ9KLW18RXpropjQR3x180FUzvqabKYkSKQAJC5uMmjUnrTxIbd
t5wUjAkrboCz6no2dUOz1PCT5s20dmZs8RkRxtdSaRABzvm9YnsywIHzNblXh1e5fL2RTv7dY4X2
C+JF5DLD6zpUDJX1FtouRR6aOfsGxc8reHp+rtJ0UwDORd/RISnvLfo8IWN7mE4XNek01Ws6GFN6
wicrjSncQZcq+IEA9/jk782YJHR+FtOg0S+GINrZh4hsJ5bo8VNmMW4h/fEN3P5qPs4cesPtsZCc
e6nCGSdmSXvFppmQu6UQhMZuPzJcxFE7vZm2vOh/kyxS8xRQCjX8UWkYrzSWI7M9dQ3mw0mWGJDh
U93Ue0nZHM5dP5CxkVUtkq8+XTos9tH0u5M30zZtIgdl+8ddLq0SZsE9lWT0nqhljrZ0pqgxgunn
N2VJ9FV0lXrbXhlD99xjd4WsD1nZS1joMQkD8oHrv4RZhmqx4yGoJw8RMg5OnVKWxMB2BTsjRIH6
hgmLbHyhYEQyr0SVGEAzRld0sCwfsnJ4jPdZGwZNjd8dsVuLdOrucPaQcM4i2KCsjc0r4T7Ao0QJ
TRy6iDgmTlVgvUlwTHGozTTjEaEQLj3a+CFOS1ZE8zUpu8a2+SLcc5CuO0fY/a6GB/YHEvtlYi07
r9EAfocsdfcn+Z0fDYgi7vl6SyORdmJvkwntUgwsQB2HOhpVKkWQsKFcuor/Xru3QJcqXGkzNmyD
/IYl1PYczhjtq3veci1gYwG7/S3nwrwkMmaEwvuIm9qXclrg29n/SkV6uvehsLDp6aiehryJa+A1
Q5Ld2Atz2OWI/w1ODq/xo43pQ5ccTbXLSoO8xvFari6NAh1lW+O6P3uBNQ8gabOnfDwShsKXS9PH
902eyghrspZ4uHSEz1qEMRQcgjWX5rVEO6pXMgenCBEsFhAbpHoP/BIeuuMcrKnFvL7JjujZVgBz
GaCCqhe+PoOWIrQ6EazetNI31BFWi9AAdnENY919SEMhhxV270ubo+4U0SQbpDHayPw+XWtm1TPS
k6PFgPu49QfQH51bch7rrBENQ+/W48agrfr+U8sOa30i432ov6Jm/SryRqd5CREXFVU2a0MW5K6e
kSmZdALF2zAwVfG+8EwNo8KBbCqFp0la3qTgpJm/M+Ng5HN3AoZ5P6cYQGIEL/FNexPXTxAWtR/a
vJ/jH6x9PcK0CLiG8VPDrFzU7qCfguHkjKmIHD5RA6lrFLJcuPRYFhNuX/Sd89LUpA5kO7Sn0VLi
F90HKdHViQGm2bhvXyiMvnTpA+W4PvJR6pHbclTzfxh9RcqtJhaqwPFjeC1/1+2NCSq/Dw0pZt44
SvP80Im4QOaTwo3QDzOxUQzXQJLE5+1ZgzwZN/In+J/W/NsooXmxI9VlnTNO42GhTD7lRBdbrWUV
PEbGq9d/opvh+tLmVTGlCpWufZ0TbUDzDGAblNdAnsEBAIx7dyfp125Wui0cEfaE0363HNFVVtIM
E/bs2iTs0UipW5YRzUXY/yHxWw/eBI8zWIVIl9nmD2lAZMJ/T7z6U3BIBy41uy1Hp/d3DTrBGEqJ
bdIbZ5s5JKxaVE0+yppqTVie6AFem8WgL8jYWhqvs1i2IIAIjtPvs1Gc9kn21OyQAZiBAjOPvktB
uyLNilsCpxAuydrWdf295DOG9QiYgHIDWxZGtODvoycgFaArFq1bsHPmGe+rOpCdGm5XVFxgs1XU
bC984/ai/VuNdbHpcohp7yzGoXo7JNHT5nvrETaPYrZ9npCryfHPoxVGdJttVspWo6koNEbY5UV/
poAc6r12ekBKXoCDFDQcu0areTbmbBphlp8R+Zle9APQ4kUZoHus8ag2R7wdIrRPDyv3on7apJA6
68/y6WiiAfY6ogefXzR7s5hQ2+8pLYgeE8crndkKry6KEIFd+jMCkE0JX/Bvgcvu6PXj/K/AQMFe
T2aseLgvYuwWxoDem0rQGeW0Wsb2/cIXojbSJu7imA5wNjSADNgLcpQGsCCghuWhWENjt0RhQD6L
Ar50Fa/G+mVXWM6JA9dHpwRVepVYJkSJXBTc7Ld8FrYUJ75/srFyg7flK7Yj2tWaSKvnlil2ITpQ
zIBAQ6dXfOd4y7wi8m6n4gTWQFp/6ayxsmzHNygJ7aQc2jWjmjtpbA06r1pDtSwPPg83l75cAHkF
wbbNqY03+8/EReJVAbsb7q5pW0/nF0abcxIxerFpblfOKcZ+dB7XvEunx274LTp7Mr+qsUOcZRfq
lbiHtZSfsrAldrEgPjAL1E3KuZFDs6PdvDnXT/B0t2YdJT3XeVEyYksSxNzjRo+huZF6ofcaNfRV
WtQ7ogWUk+NC073opOz08XnqYCsXbHf+GCeJJbXUiDQPb3cgkx20MmHgvjcT6woDTnYHvLE09/sY
rTl7pO9xz22RGBfw1eXPVOghWNvbstf3ZEctiKFPmZu3Bwacbs+n1bHuHEDrS4G0D+3K4nNpYs3Z
aR8BpqHtVpe5z+7QiCK0+mgz/KMY/Y1uYb8aFeFAe0BzshH/LAhZ1wQt8zRO9lzjr3BpF+iFDqKC
j3O1mvUmfx4YN2vZ7FpvhjZixbFTF2urF/XKpUANyNzMt9E/Pf8e5FWdy6iodFvGYVfGJA9RL30t
5sGjsVXVI0DVPGjtNarG7ukVSAhTr4ZjIEmBzBS/LlJm5YMoE/X0SHs8wk1c+uwfv2b6sUwNO48v
SBecbRg6oS4veK+817B1waLWgnUYOiSYcv/nCWpA19RPZPYiLDr5It/jMNVNp3b/QU1osGCeggOT
gJmeBYk8R/GU83OXWq4kMyLsVnWTE+juLvNhYNRRSZK5AA5Bc0S3slDk3MnrmuoCpOZPhH91Z4Qq
eA32bUeuiiLOkw3Jfa5/64WunknhVXNhm6pdS5Fq9Fzr01CaRzyVUXDgPFtGL71f2VTRxKs2WklB
OzFuVr/iPhzDm4StijkZDaURdJWnkjuVPcmxWlZBtubA0iHB2+stZPZxO7A/kEcDF/qzbwej8vZm
J3P/Y8Z9jDreKkIi9PZbdz410v2LG0zux2grR5Jg2KUj8+3KmmMbB+T6+OBq+i+5WyEYawBsX9JR
34dMU1eDty7Rl6+ZtRFqSkiiFdxmMlmooQqsSAAKDd440kw7tKfw8iQ7DnhglvT/mCISSnli/CXR
cv9Zhx7W2s6xWOfnnmSVNxhk0LINWGpY4yKbdnbv019w4mpjSI5iSL4OgWE7i4dJ094DWNiW5TiX
kAU2PnfFGMyQ1d8dk54bmoguwGNFXRIGky3jNnfoi2cFlxH1iO/Im8zUu3tBKNARMb4w+OGk+TbS
XQDJLy1z3SIsG6JUe6jt/lKU1oS+nU2a7pYkibhnDnn38CoBNhN08H1QJbKczDymN/Ge6NAONSHc
kMwuAPcFZnGeO9IcAd/siQpkNlap6KF/Dte9rvmDRkc9+1/ahx2kdIVLxMgQrPdWLqw+42S3WVA6
QZoPzOsb15oxWzQ1ol1uv+2tfe4H5XmxIANskaWW1v3EnO4J1R7hBJl223THrV+xb5RP7dxTkhWJ
32+gYGo8noI61ws4pUOtxB6T/ca1hZ9E2Gj7bEGbHLBW2zL66dHBpotJK7JfOqc1YZFTL7arfMJI
jDFaKIgfqkvgDKbk9q6PUduWPdiXwYpYk0/9Nt3jqKCPbP4s3QSvgG6NZeyyBkGys/UDFs7dpzfC
8+UXKhOFjmaFAodoIe3BGHmEprYcA2d/qwhJviB0/dfdSi3dlZX22Vzo531oDcjfvfLEbDGpVWDe
W/i0DJ64dkQjdBOeFWfPsSvMANLUdpjr7dVOPR5ndw9ta5Y0w9SwBXW9yrdNKccWSDdJsS3GmmUp
1MAfi8Cg/McFbC/m+Cy35KZmfLqeJl3zw5vCki0mYYHHyeXfD6yx5KigWQ594sw714lkGBXLXCkl
5NbN6VAR6WNyibSlzcBy6l2/r1jGm6hzIu0yR5USxrtLIUgtN8zuIRKh5Mco52D/327Bwn/MggQW
JLWp5gWsAelb6p/OZ9OdT5a1/0weRv17bIurv7lrSXA5TWJncIWhvBt6tv//wqKP4bRzfQeZcj4M
O3VJQKjS3KnyxY0QDFxo48J9ZyTHMuf4j92f/WzLj0Tk2wAh/mSqYrfIXIOX2NHP7s1nEt8TngWG
JSYGizuErVctXlXcDOUMQetB9GkwrYItx6Tcxcxa0mPbxKGGkpxfIcF9H6UCpalTDMpODZmlKyYj
cHy2dLQ0ghLHNpk4sLZnxkNw8qM95JE+nuiWfrnGeI+s2cAE1CX8MsIvyT7Fhy2KJayF1MG92Jyc
G3KH1gn+SXIGtns/i9BJAd8grm0G+EuqVSJpoAF5m6PLIUGTjUpCIGUkTb+mRkbZeeoiT6x1H27z
EJSlVgFU07cUWW7zxNfVmBEUKEoxV7D2XC1H6ybx5EsAnYoOFJU4MUBmZDL/hlAVhjASPlsa8/xX
luBPLmAql2197VkdIZVGh7lgj2I9042LxED9hstW3x8pSXUVhclEr8jknKgTNa/JCsEr4EGPA1f6
06F73tBBbdZruXhvFyR+4xtD+V9zrtAPLbrdhomQCskWPyfq1jgwFQK0S++qyabIvGyZZU6KwZTo
QGMWX6Lexc2FbjoiolV4SBnRZZhOpbdWF+Na2YhKKkDKWb8hJuc7GmXLW2vX5r4sr4cZqRzwUqIx
J2C0JmV9UR4WtAAS4NkCx8cxRmY9WWtDR0w8r+qBb7schEyD2UxB9a2/7mX7+q44THNBidIPr07M
9A67McJ67JV0DaUkZOFfHIdCtuZLh5n4scJSfFvgJhEoUZif9cnpwJr/ilxatspYGbMGCvUA6p09
ZN1GlJFlw2ac+Pcvu7cWATzeLx8MqrHzzUDlc2bBSh0Z8HKlmTTDgYczQxWyqjM59Xi4SV5pAXhR
9F5iPn/tVscSRSUC9nEBai1DuVQKj3yS1AUJm/XxrEjmwY/HEI2kYrxCkIUM/Lg3XMpyXPAj2oEg
uTvqXW/bEwztDS+jrAcweU9Z9e5wd+pAtN4egSJJh/3qLkHFuLgMgr3WMxmXnvzXk8PUfMTHINRk
TqcelEyBSg/yoScjOXDBA1pQDGlIVTow2PNx0b/kTbgDOnWib6l/Ik46BOGDmYl0hWMh+OqIh+tY
PoODt0OCzuHBqr7Izm72YkqpvcQt3D7+pfG76nxuNWwy4XFi+mjGC4jUe9nDM3yhuQPWZlq0oB3n
lspKrfB9JhoRrBAzS1ykwaBWL39TZFW0oV5lAMmxEmcfuv9TA9vRlQwukyx6EeFXMyLy2YPjMqkJ
8VQ3t3RRR0zkeSPDtEv4+zml5Qv1V2V1rId8JRJMyxKgEGv1tUoUaF//83NOFP9aiRroK8kRl6lN
/Wl+U/SaO4N79sXb+GkXq66WaJln0wnVpyrDH9ZTAPZmeqt9QHLWxLwAaHZc1SgjqmGSgknAauhr
f6we2jD56fEUpANwfKqeOHtBBmHRAghN2s8DmYCdWhGDiuLvYnpxwrcySPHBDdomZ3rR/lxyc6/r
zskjqY5cQ73JB0Uc6hY3Kzmpaicf+DavaklDX1qYjj3wzRKKIL9nx6WCS96N59WaWgim3ktkfq2a
TAJD5lPvTSfG9N9W/EC5LUbDjuybMoGHQbCXU5W5pMh3RERFAytyvOzsdmZ3K0HXWFVy3YEhDoKi
DMDKH8wAntZ3ktbUPcGIqjlEJcQIXQH78A01ira52xMT51zjxrW2ickyEo8LBZCHm7DGpKDA5qJs
2ehJMGmSbACiNd1kQj/O8NDs/iNaBu1wd8LBd2AS13lcyMBxc+KxZjEW304hyuENU9f9JjiXQPp6
wN/k0JjcE7OsAiJVUlseo5pehmwQYRovRpDyXUQahoD1FldnbzGE6Z60FAM4Y1zJZRWraLIgh3Qi
4sQFuwAQCu7HU6WTMqQLmt952M3jw/W1ByXLoptJPOA2KHXCW3yfPHPRoyrNkjtXh/3gBGyVnYfe
6qPcJiP2YiW8FA0lnnRsDEyzP1fDaFKCq51K1ZtShgaHMUfXsfQTAqhSNDuoTjbEyjie/l9R7Z1H
hxQcNEGKqrlnp48kqngt3OMbtLS57c+GspUMs6XQSgySl+cXpSUjcUIap3VLFJ81Hr32swV6mM30
U+y/OugsHnULQi0rocuJcFWCQhES0Tw2eVW6kEX/Y3lNg2lClQRo5y93MQREnCxIVvSUqSdHymUi
MTwQZCK/tB+QJFk5s8peYqbyDKxq4sCtMB9bPjBG0HVgLhHTS/xsjjHPdnoNSKxQv0lfCVcReSqm
Z4Jw4sd3yzEf1U+9Qny/rakoAbcm2luZmEXzYzHqZhGpIFPIpm7LUgujPpf9p8y9+vZ9zs7lIImk
lEDFHD+QDgTWTxsIa6rB/LDXUgAHtlO+mgoBW7ArVtuB9wf2jHk+tai/+bQMWg3MwRzwJgA+4Jb3
eXbYtr7aj8Lq2w53JNm4SBDDkYGUItLEzQRWIaEVS2VP1sGvtTbwezuQUusjc6ET3i+X9XYHGPDz
7HqawMVDKxUxmySK2SmMYJoRtIos9uxEGYdx1Gu0DBsh5o1Z/R9jeA2OnyYJHfKSs+187VSGaSf4
W6TXiic6hpxpRhzgsxDev0AA+341ezusbyXDXdtLh8a6hd240etCxRt2g7Y0W/ew5UuDxfYQduck
QbqtjK7lKQQqVtqIXFj8dFQHnEpqEuGbpqqFbvUo15FXCoGR5/FdB2zuoZLr/9rMZZfjw8BeYTWz
u5v91PM3ITK8JhTdoge9nJA1AgvYDreacpoxejSGOGIqwHU1yjfBPPqECGuqaPnq6s8yDIZ/ByrR
wk8k589YI03hVbPqXQGWEiTNnTXgsGV2VbrTPREIaXvm+vEUNN6AQZcwq/VEjd8rR5l4Kch8nEyb
n4Rhlos3mD858QSqMu0xim1mJBiOGrqGfmcs8jdDljCf74NGNFrJiHp7rCyRpwf0DwCHYGNoTq7X
Nz0s2IlrCWxMZS3SpEwzCABcL61eP4jr/efg1Vyw3MvNIg/bVFeoLK0lMQBw0J2Tcu6OKC11wjxO
/KKoegzn6RzDXZc08yxE5j/ZOQnw7oSJOsPNDCPHhOe7Fgqg1AxV6fLrNTdKdFE6LpjvpLVcKPF5
Las7br8wzW+VxBAm5HIUg1w5UmeOtLl3QvM+c3p3cfW6gnw7SP2W/2rt6SDMgpspxcwCfnwOtZlA
Fb2WbHgQd4j8X/BlJh4jGiEvm3KMSwnO70H5/oueJG+yIFur1ItefrhjhOJTftlwfhlmcNofIN+X
0EQzCrl91xxoQ5sNJ61TSJmpeDjHrSq1hZTCfmcEwBWz8MLLxPRvFdzyk8Gpx03pDtx50m5siX0u
W5VZbiigzRCq+FoXa0huULMf8ZuplRePulLid1SzU8QFsr/l/jdqNFcsqG1A5AvBPrhZLclyMGZu
FGFYivBix2hMISjkSaTrFP1iR2Pg7UeDiDnaUpHE3UZ8kb7bBcv30Me+rys4tyQRg5IcNdCMfSEq
Y5YK/dyedcO+RUu+1xnIMmRS1Rxobc/9orkgG6EjvQDrqDTbnJhUg8sUt8cV4PNJSkQrHYXm1Z8/
BsrA/ONRw5skxujN/RY3xoL+P1JoLIKHHiQFDSCyyqGmYyENS0h7FKQ1DaCbBOesuPJWgzqMRyT9
rvCN6EO/1/C3MkMjuc/DOD5J9JTuE3bebsQZCINv7XffzrLZ8Ra9mFqSctCcDbMG19lsky39Gv9W
1kLSsrXIwrX/F8Xn55pB0TVHgEXOCBZb+iUKIJsFWgtNHGYRyoKAmt35oYpJws40OgFi6/A94SGA
9Ex+ebWw1RuAL6wDAPY9KOO25J0jgT3LRSYzjIGrqzEiIsk2pDlPY32pcwQ/hVqQk6osbBhDbgiZ
i/cnZZobCIHbmvz02pBEFNp55gBNryNzS90mSlsTKk1LvRFf68G985yjODDvxqVWeBoahKc84qXW
ltIRpLBeUfweKCyK/GNpXl78R4k58+gkR6SwvlRFXMrkkC7ubObQDhqFDm1A+l48Qe3Lo8gZdkgW
WdGloAVyeQQfwzTSg8MhvNPbP3DRG8PZa0nWXn4cb+qYeUbSmUvV8VD3v07LCTlsEFymcOJDWR1o
5c3C00rFk93whOPXMYpxwwf6cY5xnE+4dKBYlZ+jXh2oR3SDV9eGgVx/jP/g9EGCUOwJTNC29BMx
VCx97uLtuz2BhgbuOtgmsj+l5vdEBSRsVfktWjou8CKPTIw+rba0RLe9L+baSJwSEbtFY0NR3RwC
6j1pfESIJfIi2f3ZPM2gO3PgrGsWrDgA94BLBdjbxfWtNnWbtq/AWdc89oYmzy1FeKHAdv2/ycNu
Y2atuOQG97vvLi0AHYo/zT3/A6zMqYruPTAI+p9vd4xYmn9J4ksBh4fJjNHjJ9LYlUvfxFVct3Fj
Ao2dnpPYJ+aMDa5yWMt6I8Wa4cULUCJENO0/yQdKXCUGgcMZZkfZ239gHHyk82nYk0FY8qMQWh3L
M1FSI2gCAvn/YdjvbSXgFtQoE41eHpGn21Bl6msr3ZJ3jznMiD022LHR3enYYggl2EeBUmISgms9
G7ugQZTguoAxWSlzo56ta7XaDc5g65OsrqFfN5WPHUgB22qF80u9gMy8koHaCu+YZU59eNVmS1DP
MdqRJUa9xvaLWx+/xQO79y9E1ENGRcoDy04vcirdg1jFnnNuM5ticYEjLVRiUg7fIo0InSai14Xl
NB2ldsg2m6HYR3P/F5/x0lxjw3ShMzfdsCGihF/rMBK6ZnxSxG5Ht+1ZcNEAnu43J5X8H4faD5Ex
DDkLWxy4bFsP64MM1Spr9vWxJSVj+P3JKS3oVOhCIXBsed6JKQoSVhAGUTLRlkXm54ANeEfZtnCM
fwqZoRN2rMBveynB2VsqpPz0fk8luBekFZYGb8056fieSPSdl92rmZ/eY03e94P6HfBWIZ/pGTXB
HgfGcb5tvsbRt2SDbIc8KM+81M1qXAgdk7ynM9tXGAK6PriyWgMfjcdXCnHNbCdahpf1xD+rcVEn
MGdFvntrOoRTq5RspdXiUIFzyBZaSaMJFCBzQ+IEOKAD7Xskyg2R/HmryGGR5/DMXwCvHBv/qJxQ
2XmGavHgnsxJYFQ9oRI/Dfn2KGzSaxYb5Q/wywoGSH6bvVvMdl3p2Usd6AiYDg5Kxu3JnbpFHq/U
zk7X4TvKDXRX/MmeUsZOE4Wokgm2e6LdMPOxiOFU+GC3O+gj/yvnAWCofxsq/LGqtgItpULj/qSZ
wqJEdjrmbYKuHLlZQftl0I3ZmN8Jnw727oSe4weH5bmnutlRl2UKQRlTaGOsf8u/cb+RtHopZs69
YFc6Nx6BHicMRk/AU9hFTgaU4bZHUTBWJpPMl1n69/SoVKWcmIAwl3DYwbusNh/HycVNBZVpTUci
I+zpbTxBXeLDogyoZzp/rXJhBBrSpEs0PFtoD2aTCnlXLg5hTLTUGjhe6HAfq2hl6ETlwB67DfL6
7cEk0s2dwomSC6pLcAG5JlCnm6eJSpGuQQ2jXbNITw7T8Nos79q24OwRg8rxv8tyXSrmMIGe3uXx
evf+bgYiFHUOSC9p0Vnd1kLwwBW8f85PWz8MsCu1bgZQBQsm0ObZSOHnDTkRlxpWYZ08/fe4u6n5
IfLsErliwJ/M72tsm+62JLmyEWOOf2oZFYEYV2bc9mI1OKqKbG7nR2+lig38oPoVQJYOZxNRnIvP
OYLLQK7w7qU2hCx0IwbK6783Iq1uUWs91VcA2dhgrRctBJkgvVVM7ONtkiYiT39a1reWijMTENyp
b9meoMnC5tsmdng506Lye9tdjTFwvnALGvN+buvQKYnnZEKtAt0cPHqNXI5yb2gs/jc6ruChpURC
+3G2UgH5fK0P83RNwqiaisBpDEtOvUUnkyj2vVg6Asas3zp3YOHopTojXrggxPrZSVBCxTe9dy/c
awVasdZepRnWw77xC7L0rCxVFerHOK2xqyybnvlgIN8hgyjPFVRENzq/YAAJf4tg/ZlmZtCL5Ov2
0vOyNSlSykzFG+R1M8sbq/+zC7Tz0pHy2WdKGxzJ+K8pDXk7nC8IobP5vaRm/uVFgqkqicaKR2Fi
pyPIm0QcG/I++GQcNYNNVuYez3Am4VtBijJLDrQrghMLQNziw0N7m+SO2pdpsFedS+YvGwmqfqld
Q4fRQqykl5/NwitNbr/c4oWjV53lt91Kh5ZRhEFMtX7cAXR8rdZv2Hr5bfoW8ynP0S3neKONEJjP
DE2Ux69uTN7dlsD8XXjUqZx/Z/lhX9ew3m4hKIBAeIF9OsFRLl1ZHv8lEInxsorf5IkRTFbvwlvp
1/ZTmuR7vQG1dgp+zxamC0Rn5tLx/bgZO+VGMGlPTTO0tb8G7V9qOYNpM3Vvh7iOo2pnsGmC/EKD
6mNDZZPv5P6F7nPCz5cV0+eTDCsFXcksVvXimFH6jRkK1OHm7CKwU8rWrDx9aqj7x1vOHdMFlt3k
6ZxLUwj0WiuyEhK7YG09RmBAhI4s8kaP06FLvaPP9OdUtdm836gqaFov+byf8gwZJJE69OmuPGXG
WtjjaHH6lwwE4xI6qO8fJaF5wFfA7iagyhlazhjy6+kZ4cHD/WjO9D2i4LVYDMJtem6IGKyONP1E
PzuNSHyK2oB/07jJZ/l/T8UL1coFwQPZGoYE498kJyy6Azu3RN0Pbv7I9iBFTx9V4TmZ6oPXvvix
bAQqeIRbNCCuyUYNguYN8r1iqYzSfqqiBKPV9CH42yxVR7iJoQD0wM1ptFtSxycgYlx5CR1So+Qb
3uRwTPWsHzY9ULAsvR6PmDFNWMcFDYCuFfZeOz/9mlmPspt6hAm4nd810f3qra1v4BjGky67JPQV
DW9KL0O6x5TuWGJJTDBmHt/YyHlxa+Kg1CcS0O1ObQyLXfUlOcC9Ue3yC/m5LgTEFiZZuJSJtre5
IVM6MBOznrTnCjseyjtXci/c+wjJ/jHhsr4NU0ktXl7Ve8oWkh1GKcjM4qi9SpA57vT+SvByE0Tj
jX9oN0Guv6b3cDWHjDhMMZ6iiC3GFPWvvp5dl9Hc+KyAyf9VVnoBvjx+qK/3DhyTGnJgYfojAaRI
Yl03hWRO9QbPA2pgdSCnwYBfNDrJ1nZpEYAZMemA8f+cM8fgdWjb2ZaaqbrR/5gcyipnmdsiue4T
eCJdgLHd2h/lqWKac3wcSNT4w7OWBU/JVxbx1I3iW0V19hSwLteLow4jbbo/uZapvCyZ2AsrnzNd
r7uciw7W+M/MTWwU410IrsSQFzG4qK8EeKRRPHk55F5r8TBFV8JhBEIwi6bWKZvaKJ7v/uvP1KH9
0w4WPaJWhE17zT+TKZ0lRxDDoIX5w1Gn2qyDy/JKFGAKFs52kpElUMGRbJuVG1jDFdZ/Jxp4728A
XMB2I3IMHwuSbgPtg2skAdZxK/6qBVIIv8juJfNnSRh8IAVclbTet+aapTHeQJM53KQT4PEjrcYP
4xaKsxzslQBL3ed769rGaDPxC2db08h4eF34W6zrbCV05PiZDgBqCo5m7JJQoc5FDKEx3ZyeD7/l
UcG+Buedma9aK8t+ALPvoiSIFQh188bAQZnogq5HDunC0/nrQb9PRcFMMfxn9Sdt6gC9CGceMRHw
C3rZlvWCQ9jEl2e61oI2Og5v2+Tfl8BhcW49gAjIHzJ5GenBkioKGbmxyD/priRYZVWFLK4kpYPN
TpMwsFaCxSYLyiorzbjlzHQbHtYG5r1JnucJMHXrjqlE+BkNwzmXTHBJnHNSFJjnToZEvZwEeOiP
u+MTQDLaSu7O9+x3/8DjwILT+CPW2xRWtBSBsFTE6JFSJ9vxSWNlPBPRgENRt8N7oJc+Ecg7n816
jYbAlS7Mt8jTdjYnYJfXCofIMEeXi/SceS2XkdfFErEL8LEFrhjUywDlF+TfcZJS4JLGLbrZCrWR
/N8TlCsOjx0EQjhPdzinnjVnhhL7sPfEdm4rtLo4ORzbgmP03P/hzNYg2H5s2c71t03MgHmtIm6y
ygEu/IDqsoTqq0D8aYfDa9qTqBs6YGcr0ryRq4fpT5W77BAYf++Q5XKnqDZ6UqM1WTavxZ3iDf2R
wo5xl3S+qLnur4ihoYIZYiMDp1deq21t2+WW1BIYO4YpAc9bnuSH2KgBSMrvfR5Pzraeft5ehXfT
LXLv6dFeKwztRBo0gFhg4dbaS/hoJRpf/TKdVF6DhBu30IeeGughWI3OUVCj9vYvtLS0/ZNwC3R+
PcDqHkQj4obVjI44EssOI6kVaLsff57wk8em+eZRDlY/9H+DeOu3noCeVMk18BazM5Il1uW4TSej
v5lv1S1nLvH14GywGD8l41w8LaOoMv6yvHxiQCdwzdx3gmCftSodpqWvsP316/2v4716QQbBWunY
T+7MNa6vVzYxC85tRWbRXCyr/r1ZTcifv8QIywt/MmzwVJZx6HRNMWMmJKo1wZIVXRYwrk0pBcgB
ZC0G7oKMSpo2XoGeZlDCI2LPP0FocpT1HvAfUUDNPcToBnURX2rH8UjbhCwQpDNYQGrzy/OgH61e
Lh5aGqhEf0JTga5mqdQfDgyI0pV/n3Qd6BE8WZCILMPlRqEY5dpop5G42kIZUFSuFP0tFNi6gehh
ZKYTp1oE/pRYIWfCAmP4EuFZ9n2795dTvFPIxUlhA6xp28JEMRLp9p8Riqv8De2hXfIpoQlHpXei
EiGnEde7xjk1CCv6Vr0ZRl+C5m2LaJ/RXZ9RqXvK4+FpO6xMr9JkIClMMl8yoqIvcZzRIUHHZKoK
Y6HNBjMqBfiG5tg3AD1Z0NZtYY3/CUX1iWsbZ6+Fg6DNnPdvdICdcElkw+axqeNxKfCHr1hJMUra
YamPLb9cBfww2fWKoKWky57fAmtp8NoMIeNIjsZ3WxHmHK7TRfzLzS8lzCsobE90tsdVSC9Zs3Z0
Vz/ApVRrqauHtOlpkpooz6mbVNTGtNbTbdK/K0y4m50UE5qbiemSKHmUJP2k7MzA6EaiVCW91Rcy
RhZdQtHv6qIaHBIlY242BhjCZjzcgODkJJ/a3AHAh0FgTIZRH/OAgm4sZwbid4A7625BDCHyT1zL
pjXwI0gUeFHbSXD8+PhT5reyOznk3avz+3nugBLLMPuANlri3/yuQCEbCJNW9eMen+MFt2AKYfj4
jU6jCAyiNyulwHbfS+VH7PYbQdPiWboDsl9D/MaSlWeQ+y56ISb1CsRbLPtES7J3/3xUqzSKGV8y
Y5cVOmS8Tpkx9Nl2mKzJ7GVv2mFYN1djcmOWGwuzBD2WRB4tc3ODXOEza3Zu93eQ76mcG3M0JTus
0EU216Uwfjp4a6kuJAFDRjq1dSP5SKIThiN7KCWATBWrYHb21f1j6QisZX4pkvvS6oWE6kEqwCj6
dj+7Qz9HONIpNdEdAEUj2Fp9WWbmLARZcA8tXdXxPG2+G3Lqt7USALH35SgHgSMu3AmKJJ1tTTDL
THR2cCD7KaFD/VFo6dJJ9ql/hmKuFEw9KXrv6dg3OlFxCwbW9JScWb3Jl022SKHOU6GjPpWKoARQ
7uuADNV5fGjVRWgORUmhEpFfG2/IuSr3ZWWh9BzCpieQoAnEQXd80N3iDscTakvPrIEGNui5J4Om
jEGrBwsqRthnc6pRt0kVla/aMrqwqcoIJs8WNNPck6zVDVDN1L+2ApXtVP8+UABP2CeRNha0t5hn
O+qmRPJRQxqGmZ5bks4tnvxfSmUWt2HQWF9Rr+U05snAb3Xa1UV0E9ULIxecBox1hPWJmuf3NwaW
29enWtuT0KkR3aHPdbw2inXixkqWIyNsEVvNNiy0mLkhqFRi5su0SNFtToOe0j4/4StutUkuvN3l
f6Jpu3hfd3X4byX9vfLmKnFQM8Dc3IrdjCx0MplvQH5UuEEPKMtLdTu9Mc8LgZsavHeaZpfJPR6R
YapWzL39AaSFfZ05DxiYT2E5uI7BHrPM4KFlpovHZQolMSZiebTLXp6dr43+SP+UyyEboFiKrZGI
ebHMFxHz1XOJk6Kj1adGhhJSnrNqx0oajfpB/kShwVLoW2vjW+3oviE39OKKfz9ez2qFi1U+peGc
/40yxXfTvG4RQai33ceTXGgUu555xEXnSb9NgGqTKFwtzvMpPMomNhsFlN8PGVo+uMWdV6w5mv93
ABsHFhyXSKx+VtCUWaxEdtsI/QBM6AhZ74HXGjJAszRndiaFrmNlNnHOl6sZFMaZUXKIk4XodyTq
COht6t+IrR9zz/imP67k8C9rq/RjI3h19BkRnrke/nbM/fbZn2M7WF7IwdtlQ5ENRNOnKOEwTjzc
jSj1YKb0dxCZ7CwMJBqY7uesC0HHVihBG/l8BRZTTJltPJYgw5sY/Y/KJC7+lTxiv3386XrYPA1e
gIZiTeZ5DG9Vd0OocEEBMdOs7w1bk7gBH1EsC5FQNFXpQMulRg7k0mMFZEh1jc/9LAtsQZnrWg5/
TdVTPODWcXGs79OF3nt7BODAyTppoy9WS5v9vc96CVqE84c+44dqPAAyxlAJayz6IC3d7yezOnAG
jFqz3FEPs8OYeHguuDqap5GpqJ6z3wakCTUoJS8Y3AoioAIsUGqR0WRgkSjHVJi6hc5D2benI6Ld
hiat6e039Q1C18OomxK6u9dYcRScJLeZj0VWy1LGjSbjKjQwLVFSaiNDc1Nq38HOffnA1IrZKEq2
fqoIchjsWZWlOR3ee6yl4V88WIYO5SWKDoPywOhd/g5z7DLN5fAcFOyZQNvOVbZVHp/4TbsPUfOO
eJIDLWJcr265SdDhf3/mgnO7s85D0/VmpJwQTAwCYgRPXSypXRyw2Z7nJ2dvpwaRLyDo8XAembl8
9Fb65eZHC41hWSZdNXaholbFsc1xD2RoNj0gafqYVnufpjuLH+cPO/R0Pv2CTWwrrQOjIzUwzBVP
nG1ik4sPrc/Unty4gP+BR3xlGu7k+mZJWcjvD70V0b7jDB2dPnYvo9B/zGAUzbvwUFWzU53+ZISV
3joIoTrE/DNXjaitOgiZhCcVGnqqM91SNE0AwWrIvLcXNViR1jkeFdie24Ypm2+PE3oKrx6KbZJx
sA2+2FQZxBcFxRmAzexa4QO/lyWVbtBr2DSOwUerMGhZ6QeJPQNVYD8X4qsHTRTiIPXApZoH9SQX
Bwtpd5FZ07H6O1SONEOpCqLyn7glVoYkG9mNMYulCTxdo/0VWIZcOSps2BIT+mCL1CIT+f9Hv6O0
/BNyBwWQ33VMR5U0ag1VKw1/gwTw9R3OZlz6H9kSlWLzMU3LDvGwduifgod81CRwVzT3MzAZMc+H
t66V8aLB+qxkp1T/irCnQ36qFoYeDhlw+8++bj+yVEF/aKH3me+/khNR83jwFwFXoJwRlAa8PtaL
7FEGeKLlWn9atmZzDB1k4XxWYK7FVfAqQ50NP4P6NAtucXSXWYuUTCYVPnHLpFu37fJngpittFgJ
9UPtVpu2SIYdFf+6LN+57tRZrPn+MlTFP0pndd7GrguDAssqPx0MTPH+edxGeNQdp+wdbWfDGOYZ
ob2bWOufDnAXB1mPU+5G0PVh/Bc4nLCoExoKpNfbtnXaIwPHTvxdnYDxlh9DS6KGMQj9IdjNufba
mPkUyd4DsgxVOv32kw1f/FSnXfhmsPgHDubTibMaO1+mmc/+DuXvhqVWSFLkuolZGq2zlAYIYPXB
Zy5aJnokz/A8aAOF91gYDVkgwFFDsMdyCUFTL6ERnsjCUZG1Gt8a68ir3qzB7TMa5zv3dHD23Lpm
QhjaXst51N5+HVpV0Jxo3zXJILCwZoybhaTjS+8+gSbgweEiv8/NDJLwoxawMYPv1418gL3TgrLh
JvKl2Izck90rR1ALXMPHS9jywpgO1yABSPlQy2AL87E8BnY5WoSN+ZM6VlXQX3Gbeidtd/m34siN
6ip7iISu/1BRS/ULn33A1wj7tG1fjSlfENj1LuhKpdu182C6QVqVterqsQvBjUR3uGoGaWH110JB
xVz144N1oj2l3qYgDIX4RS2l4/GD1rqkHVUJZro+P/daUFeHmDrUpHiFeIdTcfgbQ56xDn8w8Ngu
WtGeDPWZJOT78lG0Sa1m/bpyH6SoYesukmdH6SrNH9rN+2Ug33GyR/hv5D08bENRgohtTovsKHuP
4iZ3JCd8V4iNpYodiVCFG5X/wnoMv2pG8FlPtZzIdKcVn5tEjOTqGVQ6IM20OaXfSxZVo8HvQgHc
mGgGt7gi2TJ/yndYzussSp9jZWn7NhbHYUXV/ou6S4IGVHvIVRpDcAuTWXxsaMJdhBDccsedSfO2
gCjeq3Sh3ICIQ9hhGoRxPVGPjcAjX6ax5AHiWUqvCTIlg3wR65AWPtllUdWvgis0oi9OOrbDLF1K
7uB98cH0VwdSqUWPrObHTT7P2A6R0ymoDhqlggI5KNQEXErhizKiRV6lK/5JMEWYwxu2TMiWgPyK
awPqbVon3JsvyPZdRps0NJSUahjSruZMiJns1o8vje30k5cjHJdtjdgzWsIDipnT+AtJ+xzVyweh
o7GQFqZYzoN8tQLJwhQkqYe2h8MczN9e/Ndnd0u8j2L65gk8uoyZL1CyUs3tBsRC+5YtYA5tT5ft
UB+ZBBIHx73QvUImVMhlck9GI/EBc+ioAYi4L/OZeAnUIr10KL/GtBXME/MQdz+xnenU4coiH4Hj
KfyJCKjPPsEcCI41ER/13aG0qjjZXC3UikQdSHxHwCWe3RNVDtUQfaw3NGclUcjPP3n1u2LlDvAr
UMon2WES0QelUReRsOemovubAfPg7H5/PUDnXVHBzg4GiM9+pPELF5Mvhrp9VuhI2RGVulZSoNUD
KNLHOGX5LZ0NVncAHVqfGDWFdav3Vyeabn39QW5/BKIgiZoqNzFcH2g9vEMXnN2MKPi1bO6wpmCk
MAPuEDuLIWBiGvyo5l/AR8R87GIHdNRvUL/Yo3KQMPnOcSZ7ZPMRZWAdoHxFl1tdi3ComlNwTZWb
rfZ2vaEVWHf91v4ovrPT2JZ6BARirT3gSFMtZcZVFMSgT5yeC+LeyvuVXcdqAnFC7ACTpTPLgLr+
2EVBLjevdC6tNJT/ZX7/61r6rhWnsUygWIJondZI7fvsJe5Xs/OnZMVeR28r/RpwSgyH5vuO7z9f
N+V4q9XAEG2j5u0nEut7wjRTA2f8RfwmH4z2yz5VsAP/rC+O2xnw1Cj/vKY+UFROSpKgy7vHbS94
v7I1jkBxyNEbPFa3OrnUI8d1z/UfsTr6FPuRVVqU1xLJhSnlRtpaM0jzjl/ljs4WsDjctorVCHih
xT/W8ApLuSeerb6UrVOUNsSCJncPnIsB0Ol+y/VbJBRECEwRE6OW/j4leE26nAfhWc2YMeBuexE/
WYHorNgJOTmma1qBOKEcofI0ppZ3JHASuCPuKpwLQyABfnseIEURURJrER7oZlG++V/qkBc5nRJo
5uHh44zV03RUHwvw3JuMQVCp7P+df57ttPbnIsSp+RLoXamD1mjSTzo3F3Hx52Vh7aHkFn0A9yxK
i2HwhJfpUXmRSfSnJCcOC9MB/l0EgaVODYD7udAplL59XHKprOVq79+RnIZ/ctJ4GQDfT8DA7sYI
wiwnA6L0jWh7Fjljkpblx5Q6HpN7hBveRMkawbbUICfDdYubK754hlWDoN5eu+xLqLJ8J8THskpA
k7YJJ0FX0xwYSs8NJjLmCoxHMO+S0Pg5A7HMAjSB+tnCfFBb8DvtTClsZuOSF5ix34Gi1rHh0rfS
gQ3tyfTyiSJCu+Noyluc1Rch8bxGdC0iVIhygn2Nwaq8JGDEfJE/Q4xo1AnUgzajRGedS/cTWC9a
LVOpZS/yVNWXIHEfSeP+4qpK4L0xYOw3OxCGcSdDabgTu6Rz0IYI1zQFqmSfibcnzVSEFtjQgT2T
rw55ovB8FEMS+ppE8mFjg4KHpMdKNpwx1lgIzwsxJZxBhKXir/DZfkgULsQWyFJkjT1aMfKaqTNh
i+fMlSDFRXIvWZ65egrLXrnx0avhb6uiQLr+1SI4m1i9LN2ILO8Oiazai9hDTZ5FTkWplzqVH04f
v543j3Z091vUQNcKyFFXNYISo1f4ZqK3TdnQh+dmUeV2Ytx5sJZbIzdMxOgMj8jy5UoteBgZBu9z
Uo9BL81B3hzhYrXaYb4pr8MlFQKuvkrYAYyLT1/ap/K1/DxeKkIHIGr9LUNHBCYEkFPV5TMMWVlr
hVCgBCJiANThS0VtyGTVZ7z7rOJAAswcevPA9L7VilUfSeL1Kmh6l4afbjRowpQJdY8ussM7Hy7H
+U127Vz/xOTVUB5++6X9ly3ekEKZemCCKwXgiCkDZMhaHYAh2WyVo/OmohF1WXVns2HRsSFNGEpM
XzY6QYZUyhVczvKf12avwYg5rca4/lxafDmLeUFNIoeTURL7bYA4GH9Tyzq2AxuTW/w4suo6BHRx
ba8G3nSP//pPYpWyckcLcofo/FTy4tSXvvWcMAH5BkV+sFcMopyeD25fc+KoyFdLUjBBD59M4iW1
KzK2ybgpkQ6X+OD+Bc1BB7JwfCM0aw0f02wAZu30BUyADMq+Vf5J2ZQ4mWa2KpnXQFv29L6Y2JZv
/rq6Vl6ZPbXI2ETdGlXAAs108FiDTN0gquChGQCEjv8HG3TJx7IQETIKQT0n74TeJZCu9PpI07KM
856Hn+avwNy7/Gbk/NvRHHpPofHfeSKC2lBOOUTBZltsxI2QOp0EuMrOAOvUPL4tzq+9XTFRlBAB
QGUQ2ojIMrhWfoskrppkR+YaRK7nweRS9yFIOx9D4B/i3Hbqvt5+0SUA+W3gC59xaBEMUkCxU/9H
yu0zwiiIPNYmuUnCNK4ex96dBltdhD7+ijrP6dZ9FH2Z7br1epM93wpAWvq8F1nxJePbjERQd9JM
ut++qmQg13IaCZ4+xhRFE7fGKVKyPPEGghw9m1y8vSWka/5CSRdn8wuWoy8uG6/cbtPrN2zAsf9w
swcpGK6qAYAatpGU1AYwP+7wlDJEbLGlIEh5dqnNGOhfyrJWlrQl9ZG2aLQ4FuXxGWswHyjBf0s7
JkmH375mSs2IQWj+q4I9mD1EtN1i2MIg2PQiZfohzbhNbyTv6DDrBlQwZ1tqN9et6j39nlwX5Fwe
Dix3F6UeSJkxiLL73tpnCoFjCxNwJPJDLZ8JZSgt8EnhZjJamFj53rQpC68NWiWuKevadHEInqeR
OKGG+Y1AN+J6pgYgpO/tgDF41RT38lOICqFADF7aR/GZEx1c5+Sjp8Pc2r6wytIIbzz8AutNjvkT
3wBiLqNqpLUyessa8YzsObnEAYsuWxQXbDg6/mZdOSu/uFvvzdZUwV+xm66W9lQzFVAm0bb8BUNI
+xFT1s5beoAuRs+xWFr0LGYp79+np/TVWbHnrJU17mNvgkotEWpwrJH/OmkCEBMluYITMg/jZrZW
mZlQN6uhn/Qhl4DTtIJTDVK/nlj+WmIspUL+9VnqpVwJBDJXRCopFyeAGjGDyaKIIddO4aa1YgLG
dC3QNjTeuw4gq2NEp9p8uFfoi/ygC/8qRJJonmfTdBNTxbyRTCvpHQiO87RSGJ9hBmvPr71D3Ju+
jx1mvNYqUiD7e6gwd9ZQJ2c89ADRsfC4yTxntlX+Exa+Swf8N26lsiPMaQDUarprp4q1TUrxzLAP
uxPnncNkJvQm2wAbLMOCsB0JeneJyNmk9+QTk52z5yW+COztyHK4CECj+BEkk8wB1wRtQIkDQcMi
3HycRAF7TgtwhP+7ZmrOH0AQHwWVGnSdPWXVqKpA32hTxPFa9g7s4EBcWTdxK7md0DXUISPIojr6
5QUFJCPCrcTu0bjxyzW/U3sDL1WKLWAEzC7cEXiAsifJF+nGwwFjkOrMyMOFQ/6mKQYmF/nm+rdD
UKXq4G71Pgx9/3zbDVPOJ6WFEem6vXrEu6GfLy+XiNJuYGDJPUDWcpJ+WU/29ej76eL0+8Wjud1O
yFvlxQdWCTdLaGoVydcDxlRurDnyfYIFuSMq5u8SVQYT7RXO9dghtwEmH4reSiRKQrHkw/SKkXEc
EFU6eVmTXpGzooD3mJA1aZZJuylBKqHZ/vrTPKfgy6H3JTwnmYGcJs0sC9H1gjhihoJQrM5xTfOY
lUX0S+fCJxzzK+536fioC5PKHaZMGofQpbi10i/a02/bX4IX7hFkcOlDSQ87LoaIpz9NqgJy5oJA
hOaBszWkZVT28RlgSFkQCXfjAH4J9HyX+kZoqeLTHo8hfp8yfNMEAgAw57atO93PyZoxcv0Zq5Oj
cpRmlQLR2vZz9pA3xkAiIRjIxApbLf8CKQUVgSUrGew5T2VYyCDQadtgE6d1NKuLJbyyO9BtjKoK
b3AZaYyTIt6lOtL1AZMGBsvjpEsXd88ET+/ZeA0MddNNhTHFmdIF22/++b6IeNb1y5wSTBsM61XY
/ausovfrNfRrh8FKhOOrHJP26LmQ+1OxgcsIx/KQlqQBurYrPMcjPcGlPphI971wGeDlbfo+esnn
KouzR/fF1L8fb0DaBuZX2mVvpcmh1T6rZcAYdTz/yps8Z1Asc2aHw3oETsRoSkoy+1oXkd0MNI1r
kUCvsJrC/HnUZItByYvD201glJ/cZ00P3A7lsDbkzBsYvQ9eZBaHgcYbLPuc+jk6V4BVepWVwiHu
FXffGVWOLPafW7mb0NgyI6hItRGHtNUEvX31iU4HRAPhhd4BiOCzSbtj0cMd81w4fb7jnIFwkTkq
OgbjCidbJ3yq6jnOom6rw6r+7m6FvER3Oo52X2iDotilaFVoiFEH6egsN4BmUvc+LORDcsxwQpir
D7SXoMk7pPukiKEpGWFRJBxizTj5GwqxJxGiDQDT4VLiJ134ZHyr9r+TT0DQE9TPHkURwDsjLY1D
tIcpAOrDMWqRtGPOV/QbGMkaRUZsR5NjBlvsHJDHlqe3HFfq7JxgTpfNRNVyF0gUOjvcqpUWmY/E
glyiLKgI9x3mFsdUA5P/i7/7SnnL9J3QnnOQSJkEO3D3O1/Ssty2ABwXOfHwY0vNu14cdZ1O9gAV
gWMVPxS093+UIR9ysKcvnaRrcohe3wGpzfNTCQqIQAZ0NwX9gi4efxEdFtLErTw14wIUl7R0vi1B
ltjaXnDuqx0kMIrYW9uOz+cSk5+MLIWQsy0+gmyGeDjz3nNHDPlLwUAXwx7jjxEkHVIa4IXGHfj4
B5gd7jNLk1dNFN0tO3rub4OSoLqdLN6wI+dlD+TACWbdF7337WA1xU893uvBCUYNEPjOSt28lecA
xEUWOa6T8nv7pSgmps7WOhpqnIy1/hWfo2+SgQxdmf4xL6JAuqlOsGB3Ia4dc/9fBkWw5EP4bDn8
vmyy8XwFJ9jqcHM+7BsUJ+X9p+F3pVS7AspvWCTOFcsEY4sl3+1KQJ/KumnFFg/ebHBB7a6kqGKp
Igh+K/JAWnDoc1x6Q3ox3tlm9FXdyqZM6pZe8mpAXPOtQCLubdpXBA6Z8OwoPr7Ir+p1NXSJahMD
2c4LI6v1NKo/6d9WrlxrgiE1O7Z8QXjpEA19Xk8MzknTUdvaOc2eVrGjJSotNTHrHOD7Hp15q0XF
hAIQvZuE4SFbfNGYwlPhBJg4PG2PzfXgArJjIKZzxLwTU0vr8OquMcwVnjt5K1AfCMuEwhc+cjGo
2Cnk4k2w/6Dv2crkc84a1BOr33VhhCR+RePorA/Jt7S0PKkhH8gQ0RX7v0I+0gemCrWmr+bATqEF
px/oS7dIYJg12GKTvX/RZBIg1j5RAel+n79Tfok+sjYjXtKmZkZqXNnHjCRm7soT7ZZcwVKHPREN
F24CjUU2u1UXAHoV/vibUFPmjH5uyULc8mV1vDF282FbIA+JCXx9JgRy1tqiSmRhiH+Ofm9seyck
PZtKWZCvteu0EJBXBQstYT9sQ/aB0cX/K8eL2G5ez+2m/1zSArS0DqWNfwS3T0QyP89/
`protect end_protected

