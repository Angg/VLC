`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 11/18/2017 08:34:39 PM
// Design Name: 
// Module Name: TimeSync_sim
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module TimeSync_sim();

reg clk;
reg [7:0]din;
reg din_last;
reg din_valid;
wire [7:0]dout;
wire dout_last;
wire dout_valid;
reg rdout;
reg resetn;

reg [7:0] ofdm_preamb_rom [0:479] = 
{8'b11001000,  8'b11111011,  8'b00001001,  8'b11111011,  8'b00001001,  8'b11111100,  8'b00000111,  8'b11111110,  
8'b00000100,  8'b00000010,  8'b00000000,  8'b00000110,  8'b11111100,  8'b00001010,  8'b11111001,  8'b00001100,  
8'b00111000,  8'b00001100,  8'b11111001,  8'b00001010,  8'b11111100,  8'b00000110,  8'b00000000,  8'b00000010,  
8'b00000100,  8'b11111110,  8'b00000111,  8'b11111100,  8'b00001001,  8'b11111011,  8'b00001001,  8'b11111011,  
8'b11001000,  8'b11111101,  8'b00000110,  8'b11111111,  8'b00000101,  8'b00000000,  8'b00000100,  8'b00000000,  
8'b00000100,  8'b00000000,  8'b00000101,  8'b11111110,  8'b00000110,  8'b11111101,  8'b00001000,  8'b11111100,  
8'b11001000,  8'b11111100,  8'b00001000,  8'b11111101,  8'b00000110,  8'b11111110,  8'b00000101,  8'b00000000,  
8'b00000100,  8'b00000000,  8'b00000100,  8'b00000000,  8'b00000101,  8'b11111111,  8'b00000110,  8'b11111101,  
8'b11001000,  8'b11111011,  8'b00001001,  8'b11111011,  8'b00001001,  8'b11111100,  8'b00000111,  8'b11111110,  
8'b00000100,  8'b00000010,  8'b00000000,  8'b00000110,  8'b11111100,  8'b00001010,  8'b11111001,  8'b00001100,  
8'b11001000,  8'b11111011,  8'b00001001,  8'b11111011,  8'b00001001,  8'b11111100,  8'b00000111,  8'b11111110,  
8'b00000100,  8'b00000010,  8'b00000000,  8'b00000110,  8'b11111100,  8'b00001010,  8'b11111001,  8'b00001100,  
8'b00111000,  8'b00001100,  8'b11111001,  8'b00001010,  8'b11111100,  8'b00000110,  8'b00000000,  8'b00000010,  
8'b00000100,  8'b11111110,  8'b00000111,  8'b11111100,  8'b00001001,  8'b11111011,  8'b00001001,  8'b11111011,  
8'b11001000,  8'b11111101,  8'b00000110,  8'b11111111,  8'b00000101,  8'b00000000,  8'b00000100,  8'b00000000,  
8'b00000100,  8'b00000000,  8'b00000101,  8'b11111110,  8'b00000110,  8'b11111101,  8'b00001000,  8'b11111100,  
8'b11001000,  8'b11111100,  8'b00001000,  8'b11111101,  8'b00000110,  8'b11111110,  8'b00000101,  8'b00000000,  
8'b00000100,  8'b00000000,  8'b00000100,  8'b00000000,  8'b00000101,  8'b11111111,  8'b00000110,  8'b11111101,  
8'b11001000,  8'b11111011,  8'b00001001,  8'b11111011,  8'b00001001,  8'b11111100,  8'b00000111,  8'b11111110,  
8'b00000100,  8'b00000010,  8'b00000000,  8'b00000110,  8'b11111100,  8'b00001010,  8'b11111001,  8'b00001100,  
8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  
8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  
8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  
8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  
8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  
8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  
8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  
8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  
8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  
8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  
8'b11001000,  8'b11111011,  8'b00001001,  8'b11111011,  8'b00001001,  8'b11111100,  8'b00000111,  8'b11111110,  
8'b00000100,  8'b00000010,  8'b00000000,  8'b00000110,  8'b11111100,  8'b00001010,  8'b11111001,  8'b00001100,  
8'b00111000,  8'b00001100,  8'b11111001,  8'b00001010,  8'b11111100,  8'b00000110,  8'b00000000,  8'b00000010,  
8'b00000100,  8'b11111110,  8'b00000111,  8'b11111100,  8'b00001001,  8'b11111011,  8'b00001001,  8'b11111011,  
8'b11001000,  8'b11111101,  8'b00000110,  8'b11111111,  8'b00000101,  8'b00000000,  8'b00000100,  8'b00000000,  
8'b00000100,  8'b00000000,  8'b00000101,  8'b11111110,  8'b00000110,  8'b11111101,  8'b00001000,  8'b11111100,  
8'b11001000,  8'b11111100,  8'b00001000,  8'b11111101,  8'b00000110,  8'b11111110,  8'b00000101,  8'b00000000,  
8'b00000100,  8'b00000000,  8'b00000100,  8'b00000000,  8'b00000101,  8'b11111111,  8'b00000110,  8'b11111101,  
8'b11001000,  8'b11111011,  8'b00001001,  8'b11111011,  8'b00001001,  8'b11111100,  8'b00000111,  8'b11111110,  
8'b00000100,  8'b00000010,  8'b00000000,  8'b00000110,  8'b11111100,  8'b00001010,  8'b11111001,  8'b00001100,  
8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  
8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  
8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  
8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  
8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  
8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  
8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  
8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  
8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  
8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  8'b00001101,  
8'b11001000,  8'b11111011,  8'b00001001,  8'b11111011,  8'b00001001,  8'b11111100,  8'b00000111,  8'b11111110,  
8'b00000100,  8'b00000010,  8'b00000000,  8'b00000110,  8'b11111100,  8'b00001010,  8'b11111001,  8'b00001100,  
8'b00111000,  8'b00001100,  8'b11111001,  8'b00001010,  8'b11111100,  8'b00000110,  8'b00000000,  8'b00000010,  
8'b00000100,  8'b11111110,  8'b00000111,  8'b11111100,  8'b00001001,  8'b11111011,  8'b00001001,  8'b11111011,  
8'b11001000,  8'b11111101,  8'b00000110,  8'b11111111,  8'b00000101,  8'b00000000,  8'b00000100,  8'b00000000,  
8'b00000100,  8'b00000000,  8'b00000101,  8'b11111110,  8'b00000110,  8'b11111101,  8'b00001000,  8'b11111100,  
8'b11001000,  8'b11111100,  8'b00001000,  8'b11111101,  8'b00000110,  8'b11111110,  8'b00000101,  8'b00000000,  
8'b00000100,  8'b00000000,  8'b00000100,  8'b00000000,  8'b00000101,  8'b11111111,  8'b00000110,  8'b11111101,  
8'b11001000,  8'b11111011,  8'b00001001,  8'b11111011,  8'b00001001,  8'b11111100,  8'b00000111,  8'b11111110,  
8'b00000100,  8'b00000010,  8'b00000000,  8'b00000110,  8'b11111100,  8'b00001010,  8'b11111001,  8'b00001100};

reg [7:0] data_dmt [0:639] =
{8'b11110000,  8'b00001100,  8'b11101100,  8'b00010010,  8'b11110011,  8'b11111100,  8'b00100110,  8'b11001100,  
8'b11101010,  8'b00011100,  8'b00001010,  8'b00001110,  8'b00010000,  8'b00010100,  8'b00001111,  8'b00010010,  
8'b00000000,  8'b11100010,  8'b11100000,  8'b00001011,  8'b00010001,  8'b00010101,  8'b00000101,  8'b11011100,  
8'b00001001,  8'b11111011,  8'b11101110,  8'b11110100,  8'b00000011,  8'b00001000,  8'b11110101,  8'b00101100,  
8'b00100000,  8'b00010001,  8'b00010001,  8'b00010000,  8'b00000101,  8'b00000001,  8'b00010111,  8'b11011100,  
8'b11110110,  8'b00001111,  8'b00001100,  8'b11110011,  8'b11011101,  8'b00011011,  8'b00000000,  8'b00000111,  
8'b00000000,  8'b11101101,  8'b11111100,  8'b11010100,  8'b11100111,  8'b11110111,  8'b00000101,  8'b00001101,  
8'b11100111,  8'b11100000,  8'b00000010,  8'b00010111,  8'b00000000,  8'b00001101,  8'b00010110,  8'b11011100,  
8'b11110000,  8'b00001100,  8'b11101100,  8'b00010010,  8'b11110011,  8'b11111100,  8'b00100110,  8'b11001100,  
8'b11101010,  8'b00011100,  8'b00001010,  8'b00001110,  8'b00010000,  8'b00010100,  8'b00001111,  8'b00010010,  
8'b11111000,  8'b00100110,  8'b00001010,  8'b11101111,  8'b11110111,  8'b00100010,  8'b00001100,  8'b00000001,  
8'b00010011,  8'b00010000,  8'b00001010,  8'b11101011,  8'b11101110,  8'b11100101,  8'b00010001,  8'b00010110,  
8'b11110000,  8'b11111010,  8'b11110011,  8'b00000000,  8'b00001001,  8'b00011110,  8'b11100110,  8'b11101011,  
8'b00011011,  8'b00000100,  8'b00010011,  8'b11111011,  8'b00101001,  8'b00000010,  8'b11101000,  8'b00111101,  
8'b00001000,  8'b11111100,  8'b11100011,  8'b11100100,  8'b00010111,  8'b11101011,  8'b11111110,  8'b00011010,  
8'b11111101,  8'b00011011,  8'b00011111,  8'b11110111,  8'b00001001,  8'b00000100,  8'b11101101,  8'b11111000,  
8'b00000000,  8'b11111010,  8'b00000011,  8'b11110101,  8'b11011001,  8'b11111000,  8'b11100000,  8'b11010110,  
8'b00000101,  8'b00001001,  8'b00000010,  8'b00001110,  8'b00010001,  8'b11100101,  8'b11101001,  8'b11100110,  
8'b11111000,  8'b00100110,  8'b00001010,  8'b11101111,  8'b11110111,  8'b00100010,  8'b00001100,  8'b00000001,  
8'b00010011,  8'b00010000,  8'b00001010,  8'b11101011,  8'b11101110,  8'b11100101,  8'b00010001,  8'b00010110,  
8'b00001000,  8'b00010111,  8'b00010001,  8'b11100000,  8'b11011011,  8'b11101010,  8'b00011110,  8'b00000110,  
8'b11101111,  8'b00000001,  8'b11111000,  8'b11111110,  8'b11011001,  8'b11100101,  8'b11011001,  8'b11101011,  
8'b00001000,  8'b00000101,  8'b00010100,  8'b11101011,  8'b00011100,  8'b00001111,  8'b00000111,  8'b00011100,  
8'b11100010,  8'b00000010,  8'b11111111,  8'b00001100,  8'b00001001,  8'b11111000,  8'b00001001,  8'b11100001,  
8'b00001000,  8'b00011011,  8'b11101111,  8'b00001010,  8'b00010110,  8'b00000000,  8'b00011010,  8'b00010101,  
8'b00010001,  8'b00000010,  8'b11101000,  8'b00010010,  8'b11101101,  8'b11101011,  8'b00011011,  8'b11111001,  
8'b11111000,  8'b00000111,  8'b11111100,  8'b00000011,  8'b00000011,  8'b11101001,  8'b11111110,  8'b11110011,  
8'b11101110,  8'b00111001,  8'b00110001,  8'b11101101,  8'b00000001,  8'b00011010,  8'b11100111,  8'b11110000,  
8'b00001000,  8'b00010111,  8'b00010001,  8'b11100000,  8'b11011011,  8'b11101010,  8'b00011110,  8'b00000110,  
8'b11101111,  8'b00000001,  8'b11111000,  8'b11111110,  8'b11011001,  8'b11100101,  8'b11011001,  8'b11101011,  
8'b00010000,  8'b11101101,  8'b11111110,  8'b11111100,  8'b00001100,  8'b00011000,  8'b11101100,  8'b00011000,  
8'b00001100,  8'b00010001,  8'b00011010,  8'b00001010,  8'b00011001,  8'b11101000,  8'b11101100,  8'b11110101,  
8'b11110000,  8'b11100001,  8'b11100100,  8'b11111000,  8'b11110011,  8'b11111111,  8'b11100101,  8'b11111001,  
8'b00000111,  8'b11110011,  8'b11110110,  8'b00000111,  8'b00010101,  8'b11110001,  8'b11111111,  8'b11110110,  
8'b11100000,  8'b00100001,  8'b00010010,  8'b00001000,  8'b00101001,  8'b11011011,  8'b11101010,  8'b00001110,  
8'b11010100,  8'b11110110,  8'b00010110,  8'b00011100,  8'b00000100,  8'b00010001,  8'b00011101,  8'b11100010,  
8'b11110000,  8'b00000000,  8'b00011100,  8'b11111011,  8'b11100111,  8'b11111110,  8'b11101000,  8'b00101100,  
8'b00101001,  8'b11110110,  8'b11101010,  8'b11111011,  8'b00011110,  8'b00000110,  8'b11110101,  8'b00001000,  
8'b00010000,  8'b11101101,  8'b11111110,  8'b11111100,  8'b00001100,  8'b00011000,  8'b11101100,  8'b00011000,  
8'b00001100,  8'b00010001,  8'b00011010,  8'b00001010,  8'b00011001,  8'b11101000,  8'b11101100,  8'b11110101,  
8'b11111000,  8'b00000110,  8'b11110010,  8'b11110101,  8'b11101111,  8'b11101110,  8'b11100111,  8'b00010001,  
8'b00010000,  8'b11101110,  8'b11111001,  8'b00000011,  8'b11110111,  8'b11110111,  8'b00001000,  8'b11100000,  
8'b11101000,  8'b00001001,  8'b11110100,  8'b11110010,  8'b00001110,  8'b00100000,  8'b00000010,  8'b00000001,  
8'b00100001,  8'b00001000,  8'b00000111,  8'b00011000,  8'b11101110,  8'b11111111,  8'b11111100,  8'b11110010,  
8'b00001000,  8'b11111011,  8'b00011011,  8'b11011001,  8'b11100011,  8'b00011010,  8'b00000101,  8'b00011011,  
8'b11000000,  8'b11100011,  8'b00101101,  8'b00001001,  8'b00011101,  8'b00100101,  8'b00011111,  8'b00001110,  
8'b00001000,  8'b11100101,  8'b11111000,  8'b11111001,  8'b11110001,  8'b00110011,  8'b00001011,  8'b11110010,  
8'b11111111,  8'b11111110,  8'b11111001,  8'b00000011,  8'b00001111,  8'b00000100,  8'b00000100,  8'b11100001,  
8'b11111000,  8'b00000110,  8'b11110010,  8'b11110101,  8'b11101111,  8'b11101110,  8'b11100111,  8'b00010001,  
8'b00010000,  8'b11101110,  8'b11111001,  8'b00000011,  8'b11110111,  8'b11110111,  8'b00001000,  8'b11100000,  
8'b00011000,  8'b00001010,  8'b00100010,  8'b11110100,  8'b00000000,  8'b11111110,  8'b11101101,  8'b11111110,  
8'b11100100,  8'b11101111,  8'b00000011,  8'b11110100,  8'b00000010,  8'b00000011,  8'b00001001,  8'b00001000,  
8'b11101000,  8'b00001001,  8'b00001101,  8'b11110100,  8'b11110010,  8'b00000111,  8'b00101110,  8'b00010010,  
8'b11110000,  8'b11110100,  8'b00000010,  8'b11110010,  8'b11110110,  8'b11111010,  8'b11101011,  8'b11100001,  
8'b11011000,  8'b00010100,  8'b00001000,  8'b11110011,  8'b11111000,  8'b11101001,  8'b11111101,  8'b11110101,  
8'b00011100,  8'b00110001,  8'b00001001,  8'b11110011,  8'b00000010,  8'b11100010,  8'b11110100,  8'b00100111,  
8'b11011000,  8'b11111111,  8'b00100110,  8'b11111110,  8'b00000110,  8'b00001011,  8'b00000110,  8'b00000011,  
8'b01000000,  8'b00010010,  8'b11110100,  8'b00000000,  8'b11110110,  8'b00011011,  8'b11011010,  8'b11110110,  
8'b00011000,  8'b00001010,  8'b00100010,  8'b11110100,  8'b00000000,  8'b11111110,  8'b11101101,  8'b11111110,  
8'b11100100,  8'b11101111,  8'b00000011,  8'b11110100,  8'b00000010,  8'b00000011,  8'b00001001,  8'b00001000,  
8'b11111000,  8'b11111111,  8'b00000100,  8'b00011000,  8'b11011101,  8'b11110101,  8'b00010000,  8'b00000110,  
8'b00010000,  8'b11110110,  8'b11110011,  8'b00011001,  8'b00010011,  8'b11110001,  8'b00001011,  8'b00000011,  
8'b11100000,  8'b11100100,  8'b11100101,  8'b11100100,  8'b11101001,  8'b11101010,  8'b00000010,  8'b00000011,  
8'b00001000,  8'b00010100,  8'b11111100,  8'b00011001,  8'b00000010,  8'b00000011,  8'b00010110,  8'b11101011,  
8'b00001000,  8'b11110111,  8'b00001010,  8'b00110001,  8'b00010110,  8'b11101000,  8'b11100111,  8'b00100100,  
8'b00010000,  8'b00100001,  8'b11111110,  8'b11100011,  8'b00010101,  8'b11101100,  8'b11110100,  8'b00001111,  
8'b00010000,  8'b00100101,  8'b00010100,  8'b11010111,  8'b11110100,  8'b00001000,  8'b11100000,  8'b00000000,  
8'b00001000,  8'b00010000,  8'b11101101,  8'b00001000,  8'b00100110,  8'b11010110,  8'b11110010,  8'b11110101,  
8'b11111000,  8'b11111111,  8'b00000100,  8'b00011000,  8'b11011101,  8'b11110101,  8'b00010000,  8'b00000110,  
8'b00010000,  8'b11110110,  8'b11110011,  8'b00011001,  8'b00010011,  8'b11110001,  8'b00001011,  8'b00000011,  
8'b11111000,  8'b00001100,  8'b00010001,  8'b00100011,  8'b00011111,  8'b11111100,  8'b00000110,  8'b11110001,  
8'b00001011,  8'b11110101,  8'b11111100,  8'b00001111,  8'b11111100,  8'b00101101,  8'b00010011,  8'b11100001,  
8'b11100000,  8'b11111101,  8'b00010010,  8'b00010010,  8'b11111110,  8'b00001010,  8'b00001101,  8'b11100010,  
8'b00000001,  8'b11111110,  8'b00011001,  8'b11111010,  8'b11001001,  8'b00010000,  8'b11111001,  8'b11111101,  
8'b11111000,  8'b11101001,  8'b11111100,  8'b11110011,  8'b00010000,  8'b00001000,  8'b00011011,  8'b00011010,  
8'b11110101,  8'b11111111,  8'b00000010,  8'b00000000,  8'b11111110,  8'b11110111,  8'b11110111,  8'b11110111,  
8'b11100000,  8'b11110001,  8'b11110010,  8'b11001000,  8'b00000100,  8'b00101111,  8'b11100010,  8'b00000010,  
8'b00101111,  8'b11110000,  8'b11111001,  8'b11101000,  8'b11101101,  8'b00001001,  8'b00001101,  8'b00011011,  
8'b11111000,  8'b00001100,  8'b00010001,  8'b00100011,  8'b00011111,  8'b11111100,  8'b00000110,  8'b11110001,  
8'b00001011,  8'b11110101,  8'b11111100,  8'b00001111,  8'b11111100,  8'b00101101,  8'b00010011,  8'b11100001};

reg [7:0] time_offset [0:9] = {10{8'b00001101}};
reg [7:0] data_sampled [0:2239] = {ofdm_preamb_rom, data_dmt};

reg [7:0] din_rom [0:2240+10-1] = {time_offset, data_sampled};

integer i = 0;

always begin
    #5  clk = ~clk;
end

always begin
    #10 din = din_rom[i];
        i = i+1;
end

initial begin
        clk = 1;
        rdout = 1;
        resetn = 0;
        din = 0; 
        din_valid = 0; 
        din_last = 0;
    #10 din_valid = 1;
        resetn = 1;
end    

design_1_wrapper design_1_wrapper_inst
   (.clk(clk),
    .din(din),
    .din_last(din_last),
    .din_valid(din_valid),
    .dout(dout),
    .dout_last(dout_last),
    .dout_valid(dout_valid),
    .rdout(rdout),
    .resetn(resetn)
    );

endmodule
